`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfrxFY91sDZmzh0NPvTPqIq4QBMKcUMzQO7WgOnTpB9cshvBrWOWV94se
wKXZ32OAl1u83kmfCVN4NGiU/SwV236AWMoRED0jWMM81Gzpb5qU6TwNnf2NTE9k/rnDZB5KN1rO
+71xZOdMUpzw6RwjgdiktsiI5xqJwEz+6dehMImCby9s7TPH5Imq4l1zFF2B3M97CojbSJJLnrPb
2nUDNzp4IAnRIgw/IGtHgh7sFdgYRUALa5cHzm5dc1gH+ZE2nWz1Fo2zFeQymwW9RKeTmDNwH1oU
K0h0GBI6n4jrDpBc575cou5JC5TqAoVGq/9wzX4c2hAMiT/tu0RLgRQruMxKkEiukxHozeNr4NPK
0QBvokOFNceGWU/x3w+77UOAPIImuhrFoVnq5YUt64GF+Qd7SqhuLNORt9sH251SBzIaFchv93nY
7xtdAfkiygjJllmE0Q5PG48awXL/GFqGMI2q4lZHqRKrhgIe+qIPD+YToHnPgEOMWsMniaTNsPvr
GleghE41Q22sp4TFhgGmmZTNv9QyZPTv2eDgi9cN1DUBNN93g8Z9PF+3a31xOAh9eKbZ7/AyPD1N
1u/WA09sPia2IFkis2Qxm4dJToQ00jT1lL4fr2C5cYssnifmzdpui/gx1ygQ0mU8VGAe4KQssmzH
w8vJ7HgLsAcw9xSEZad9w23u7v8QogPc2WQESb8yWJylA5KwhkEhHCLs5XmLCg24JR2Yt6pclt7p
iILhbvJJE9+DGqp6vwRPgnsmUjdGWDrOrKeIndIMoyCnVz64GsBLPsKTlsGcHWRUYEz8Phb4yMJv
848ifMcWnFDBMu94MutOQzqUe6pqL0UyWnuauTVHZ9o6KqR5HR/zWL4YsPml+gA3+vus6MMLg6s7
f9U8AYNNwDh06mrgAJpD3BZsCGOUHpRg97dpbU9qG1w/qye/KoHCSMSCv/Dm39Siyy9uAwrbkn/a
ZH/++o5RP8jR3+A+r+tcpUjcAaKlTuD0MuTeFdCUikHyXeLindW/Mxz5N9oCne0DknR95OyLKF1g
xvxTMwzaMSncQDexcVyJbNFBacsk0STO0gmZgXHhKQhbBymvgZCjVwAcxAJNFv53Slrs+XTFu5V+
LepjtdmpDSCTi1GD1QmeqcNy3NAkr1JtYQ7WylKzs5e3HadHI34JVGCxoe0yw6dsWnAn2r5nDf2p
YJAWtFEFv0uf8rFimXy5B5JOKrv2fuu7Jb3Xc+Jnft1ikYe3zRYRWSOCMkmt8ZrGCHuqJBLF7xkh
AGD/DfMyTmBgB38EgsXcSsKNG3rUNPswYA9GdrvF9rPGcvoCCecj3EqG+sN5c+XeyUvd/AlRyMNb
TydL50pECwrmupv+oW7sLMwN66/4DtGlI7HnTpF+uom/vZ8ibalX9GZUDUtLozQPbopHgzu1kJER
8YG9T79Rk0RoZTN93c/YkbGfB1RynPb5tz2g+v6ZzLrrPdXUMEb9u9Wi4NaQ4gy73tnfcRw7P6rW
Rkmb6SUCtyijZJ3wYcz5Jb2kneyY167ZDtEY2JUl58mbyp32rnxrNDw2jUkI8ZArQupDIOY8/faP
8d/cBlf9Jj+4Bzwlbj5Lj1Rmb4C/64RSAr+e+MXUD5Zx7f5OFn6Ej3mXWm84uX25QnLY82yBBIOh
fMrgGvsYqu4v3FMYpi6VjBBz5cXhsPT3hAEB5x5sAWBSeP1l3tYTtCxLuhCo79CtQR+4ISKKV4NX
afz8QMLTcvh1GwKDZMhfEmf41GNmS1idqOYtzSt/cPqipd+dUc1N36Hnx0P+I7HOZ12VY0WoMAOu
1Dp/KhSoHUgumwtTla8F5mM+7Jt9weG+Wj4y7LJuV/7Rvp0XYU8CdL3a2paIW6270fkdlIy/bF5h
24iMR22xs64h6k7Dk8+Vhf8QDykomqb29OcTx38m+p7zuZh2Kx+3JpZfErPID199lAXwddrHOiOA
atZYdG6zp4dvK94cZs5fn7Z8nR3UrFFh8rXSkQEybxrQEKhbIh4nWu5H9PA98Wi5z1si4DaJoU6G
h/4h2COgJQ6wE0n8QwH0CyI/oxyb4kEfmF0+8Xo7VnoE+4zYxaAySKlGAExNVBF2ddT/Y7yKJpqF
7a9hdWXMnog66dgU5Xq3Z0RaW+CelWqvI+3A5NqsOasPYsRq+eaB9oPyNIXN0vCvlaqrYioQ3zq2
vux6Fr5NHS4715PWvJFUIhMqYbQJNmxV50aMTHZubB4LCd2K8jH4rYJ/TTJUSYxn+tM6ERVAGJEn
v39dm+E2R0zE30P5Pg1xxZiBPIis0Jblw429uwonUEXR1cYZ5ZqagTu8z0hEVJl6xqOCwbJQyWq8
rA9RBC5RnwA8tyg7iqQgr9wrRpCw2F4Ix6ERo8UxoxJPP9Z4nJcVhyJFcAn2LtTm/4liXvBqa85+
WpMH27iMJkZ1MyLXEORxZRKQ1CPyIXsL3Bbmc9r1L0YcdWuA4bKCt3E7UcmKIePVzMlNPejhd4YN
OEt/JzTprdISKgL0SYi6OUpxiycHhVtEyKE6SD+HXgp9x962SOnsTXxglvtTGvDTRrb3qoOIz7cn
wN651IkMxVrKjiXQd2g2noDr3LSLdTP3y2aZ/u7rodnbF3GT8GmW8c3nImGEn7ZoLJf7dD03q0QQ
Ngri0k4BXWP9i+9CERUYMeV566ruWlQkGjvICumTwAfL+O5SwI9/DY51QjNBn2kGzPZd66iypsE7
jHgfX24orUghssT3s+SlvpUCjQ+zkl7WK3EnR0K+4jp/aWZ3JExTgM3pEw8MjydM++ImI4uHQt2C
0cvlfNBLwlQylyMT9mB/Sd8ood+eMnYMSJ8O6tHHaVhB5lqWVbEj+5FkHuO3glTFMCdcxnTCnNko
7b9gL/rWZZvQUVDT6bp6LdJ83iiUbSmg3D0wgGdOqaDbrBWymekP92/qr8ggnictH5rFiDCaWoEF
sDptxBH5rX67oVleZss/N53PRxXEk5FeGfH0+OD2y7DeEOuG98XUTlorycoUR221kfGomNDvpS8w
oMh6s24bvjzimxq7mIPw2O9MLEBcmGRqLpaDx2wB/7y934sQ6MQ2x0nuF3VJk/JFXuM3IhxRoXtv
BhLGE6MV6U5qdjng2pHU80xrPT/zx+4JIzABJeQ0K4Ib1FGyroavmw221yyNWkc5/c9QBvB5OkUw
Vdg+tCbrPAROgSA7Oz3VDane0XiEWajG0zLF596bfjHeNPnpLavFXZ6MZOp2QG18+WX2pqsJ2YAP
3ytZzQZ97Zmb829RA5zmn8oJUos8tpMBdc5tY6+l+81kzAuQFpU2kJ6scs/dS7RLMYMO06pOq49G
mILqx2PXn8l5qvMlGq9JUjXD+ZhUQcdGkc1QnRuGh8cekV4wGDvO/D66LtB4UAhXqxozGh0edoYU
IbR7YsDUGXNcHjp9+clG1Ys3GdUucjtjTf6SVaDa4t+s7Cu1brQSyYIbXGsRcyglcJ0rrInI3J+p
h23rsbgYBtkdY0+uYPI/f9FDbo58YKPIS6TzKIeVMLlXpjAmw7JbXfS4LfI5gff6pZWiX1S1Ihw5
m+VZccEfNC2p/xeaF2Fqfs9DAr/Gi6VutrLphKsp8CT3ljl9l249Q5emJRmXqJDbHP2ONQt2GD02
2r1Krks+N+nS2sO/j3pNQ2nU/dClTK8LpF2jwsQ3dvRARrfSsCrnxBxWvCVh5A4nnb45t6kM4+TK
iQZpntNsczAJoaSkP1V3akZ2xa0hRKB3KU9M1Zab+LJH4sMaeR9jtdCyX4zM4NOtOIDpEGyVwcY9
S/gSatkQOKEfWC+g1aJU0hpgQA7lmvoXgW65Cvrb0j1Ud/uvCc60Aq7E620Grx5+HL8UIPV53Gwf
7B6SFaAtbxqedpIE/FajffFxykanVRztC35FN+b5KXki1nRtFgqT9VM7SmbMI6eTF0mmHm8QiYLH
2WjNSQs/GF/624qeUiLfVbkDAcqTZSvaHVgUz5nrM3RFFYbL1voAaFPF5OFqkRAybV8kf+4FFudk
z+Cyv4kpZh0JlzYGVeglqsllnOYWq/fKGFW8XRyMNdonM42l54D7ruPLf69MRFPOTAzl1FpziTxZ
vblawg2qZ5v/dBZNvKvu583issnp7Nr9ckjfEGqJgT4DI5OuWQMLx/TW6z9hJn5aFfH1tOnlncw9
YSOjaJGsnMdrocTvjqD7j3kJRGoxT3MvnXYx1vVKAExt2boLvy/wJyyNcEUtAVpEttSFA7CeAjJz
/V/gPFVnuxOgcJLJk5Nu2wqkUaHHfEx3EJITWPjHW0qah1YcTsopwiWmLuiO3kKlr/t0nPZ7jujX
gGE6zndU5JaJ7V7ruEROM0OHLhPVq+sv89P7380bO8Dwlx0lEm7upJAL1UQpp5O8xFclQjRlBs3s
LnsKqYZuiF9UJ6teEn7eCMPj9DuUWtMKC9b8KfllfvEti3EDYYsil2G5sm8YdyQdYYRbnOATaRoT
L8BmkhjBhS+I2dlFpcN6hXXZk++avBe4wTiNnJENk+0T6tei8B8buA1KLKx1ccTSQ/aarZpzyiYW
xna1cLGqa7lMePhMOOcxOMGmJXQuDBs/xOTf0jpkwX7oNAOPowJ3kz/ifV1RFo0DcdpHjXadNSGH
PqPdxnT5l4miDZux1hTrOVg00W7eFHHaCOe1EhsQYvQ/4nMZntqGiEEQalaeLuLk4cyalKKTrPu8
1j//KfpvcPcdJsriAAQGv6LYFarn47fZgAghlGMyX2Dxkk05xF9pe82pRPS0qTjQnJK6EbuDFKuJ
E1t9E3EdM8KB1sfmmw7uBrN2G5YrvOdyqLDsYsdZdB4xuyzbJyC+F3gB0e+Ev+Cwtc/+dn1uFNmg
92cYYlA8kb5kSPgdhqpKp4pEQdti/0IhRufavKnboxlIBops8K/NP+QVitcObxKRlIwQUiB3ca97
syU1XKqeDTyy5mMNeeb9Cp4mPofYnRzBVCRUslDeUy0VM5Q+ZOaMo0A/S/modZ5KlkB7DX0bP+6p
Gp3MkYrGjMQy8O+9Cgl1WB4bXHAWfhRUdyPO6/IFgZVH7j22vZXktebkoMRnkD+XcN3feRSyEqrJ
Fo0h/nM=
`pragma protect end_protected
