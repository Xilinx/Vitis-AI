/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B63nwYNmpv8yBwKbUwS4fI4tfq215bC12H/jWr2ITyUZ8bAhhKHHHuhmu
tLCjwYGpDxkCHQepQDnKydxXZ+u8n0NK2oKtr10IfAiGPs1GEVU4X6CMfa9L2zpk0JVzHC5Bo/de
6dYVxPEiGoS4Et5JvRneSxRhIGjS4akX3jji60Uc2gvudl1djOpcmHExyOQ2l/nWRYCZgpE29GIS
OfqlRo5ExyY/Ltap4EEAJo/b60kOVOBBV/T1Dlz3s+KFTfaZ7tPK+9yliTGKRkjwtOqwLvuEM/kz
W0yKexy/u+0I3pDNj1c/zkFrVENkrY2oeapWLSno9RtMglUrAfhsbsv4fC0QhUKBH/D0iCj9QkaR
8Ug3CFhIKM9399Im5aMqL4ASxlivE4EtW3CQ140kldvkuddyOJfkgZi01YMGG3qFi0W39zYvxKmj
oxeqD/kzr+SlUc02U/WbsNWfHjg/UoRJtVgmN0TnJFIwUNeYFSjTD9z3ngCnSrIzqCdvX5GTZNzQ
EXRLZIG45VgpysY8MLgOHwXtmlEjcv5Uvnn71nnYe70nwPwoBBGWU77QSXGLW0Y2g3dCdwuUqiXh
kxADCjw3X3RpRb8hjAdIlyxEFG0dguSiB5J4QvbB1ajXmKNvzqdCQPWGmupLJYL7sJYm+fAJrkBL
IRN/vaZt1pIyRdReHVOOUzv3XC31S1x76u0vY7rYTN46QBpZC5lgEnJ/GgGXrUp6BuVOCbLAG8SI
HFxuvx/dgwW52K24Kvky69/P+jILlvWRtmVJp8+EgvifnQBJU8SlW3PQtZVvgFa8yoWn78APn9AV
XU9COKaXQG3uVHzZjvUd+FzUH5LhxclV3sqeeuiJCy9x3MNrgUcu7DVOls5iBbya/fZIxZOKikl/
HaAJfmJz6ZlGAfWoQCnY1KFoTooSr4z1e/P1L2Wv9QV2D5J+hDkY2Emkp+9J2pxTA04Qq5R1OKTg
FxEOJrdow8QItlxnVWMacJp3B0qX/+cFvzxP94BFLHzwafElsQw9Dyn7wcEmB1zLSUG5AGXU5J6g
Tq/4jJU7iNcATYOn3OX3CuD9Xul7j7FrmRhexYVdILb4KOgw0Gvsz+fBEOhV0qjl4/EnpmydSq2v
fBJWr2LKYvRvrFmdTGcUJdSy/v/H9xl5VcSqyJpJrA6uyA6YInD5g+AlE733ZImC9an8Jueuxh6Y
lyzvfPwjbZO4B40z9BDkmXtuZD4DusC+aComnxmxvWNXNWkdo2bY46iQNiOAEEqqw4wAKmm+6Ei8
THC8mSXSjd3gjp5eo+qooF5GPtTyViheVOb2j6oTCvh0hFnRrRsEICC8ZlQMtDaACKxOyWcIhE3H
2XudkpHqBC3TT55ArrD0VrgjZRaV3xNZdxfHzl/Aeq2N4q0yWf4GS9Ade14EsaqSjQfmNaujp2F3
HnCEwxUnrvNnZywYaULVB8JfRR6kRa6ulUenLuoqigNORhiOx9nD9ae9FVfEKca6pwizponRXOZr
W9QyFz18zdbkHKJwEotFIifnxx6bVtOUrM6aB+rURXhHFtfe8UD3m5nQ/Vpa+TMSGhnPq5C4HtFk
yvjw4qYul5DstA8XBdyYER7YMrLJDMVlZrT4oICP/6c9ZnrkpGC6eLRJfUlOWF/Yl94ATZ1RndLB
f8oil8V1GFyaE+8B9oK3Z1LxpdNetwnTcBTZqrfHmhZZMYO08/3rG73u4JGD5M1dwVvTsCxN02oQ
9hcS1isJrTWCWyCotqYxgd+sTorQvgvdSfpY1jFvohoAW4REeWvM9Zj+h62//bS3apYYgfqs5m1k
wdeuNkofvzi6oF+zNwPZ/NNyQvOJQwqNFg3nPsZyvZSXIoQG4wqtYsNsoxzYykGeBA0wHtzwH7P1
hynUeFg0NgSxIQBhPxfdbeWTVsd53yEHqh3LnrTLXyQkOujn9CKR/+89gG2VMKTUjMuwMhmR5bkv
ag+stt3m1r5wOnSPv9RJ9RsncigPJvLH91rwnhYVTvFRcRZHSvoQ9L8A9PIzB2gDLxvV4FR0HA3K
wbD+l5/8QE1wUy3Q+IdRNfiuqHBkMSgaAqM7FNYr+K0a6+6q5rws6efLg4GpgOYLlsmWN71DGpBR
Io/+NKpNh8JEh+5ChDRrtz/aRLCM2VGfin84Z2n6McJ9Te5iKBu/7RfWQCLr4Ua9TGPr/jU3tXDs
VIEIY7L4zcbxxdJVeqgGhzw+cyCbJnlOraqRB9T+Z2uDlGJKtrofeLL6Yw2r+yXXsM4eA6XDrhrA
6pjqclnb4vSmAF53mrbml9P7/WOXHIPpyX7Sqeq87vms7t1Q8p+p3HL3ZfpABSVN1TxaT48wLFPm
jeMAUu1f852nQEBdDhcYtLQ501EJnRXBFb0Vzcz8VoPCp3PSsm0ZLolsSNl/iIXtAaor2FRJbKb/
waC+w1Ne3UCMze9OUJ7sJCsCfUIUJEHAB6vgCccL0WudQAvqzF7FShX8zEThTSLwUK/pcKC28W2a
qtcfN4FrTdJHOaZcf/OAKBJEQg0qyx/CImj5rCF5M4VLLfLOvnbDqnJ1Wg3wX3h5dgSVujc8bPPx
tjViX7rT+cwdLIzCRtoruQ9TXbcEFLX/ywWyiAqxOVAB9BYx3UFhu+oG458kN0/SGpjRxvCFZNJP
NpPe+GpbjorvzLXxzoi+y6E+xE959CJbTuGvinZZ6nv8zHEiWxTAMxgUCwdJyaiD/OLC8bk1QBv6
h3FPy7MaMphKA87qtD1Szdum/FMh46Lc8mTryH1xQONzI8Qq6v96JTcd/1d1Pj0ivvM6S00aYR3k
LFUEcQp7z/upFaQrzLlIJ0Sv++SPhai2Ff9/iHsaMn6K3tRQilna+ETeBS0BxVQUUCf67Am5hak9
st5AGRph3y8FLMPPYBQ4FAzuIAUTFYxq/9jax0yEIJlmvnGZFU5j+N5g/ItmKIDD/jJwlT4QROIR
aaPbtzTrOlZsLwJoop5rVfAoVrHoun+6PeE4qSbT537yBFbFO+9rSq8msCidsLtm039v1sopG6pc
sc8orQmH07kKaSdO9PJ3QZ0j30NNFtBaeFv9W3ttZMNvrzkHCCTnKxaTSR9MJpq3DdipnSCOFoUw
ao1YO3KbiSR1BVzuBTo5AwCUCuvFzQB9RvuJOoduFHU5cybRPhP509XduzhMLfJVzGU6K6tJ1ajw
8eQxbKHwESJHLYgntjt6UEOAi4P+zDpprXrhWffET+cW/n6I8Z8BTQ5U3ocULMtmDXel3RC15shN
b111Asef8FEdb/tWytN3TSj+wZyE4STVcdrjDWMdeph6ZpV8Cxn0XcecG3qt7ITPpb5VkY7MjTw/
5rW8eM4Z64W9MhkXWOf825nLefrdFruc5lnQ+GQVFu13ooUgBJK40/Ole+NWv/q/Qoil5FXbPkkK
R3pkcsGap3BMbfycGPS6D2a5Pe+VvyEuO7EM+6H74QOuHsu+t3gzxTZ4MZ2Nk1uUD8+1xtl6HHJ5
kYcnimyQNbU6Z2ROGsUHrs999ESngYixv8ZwInHANrtuKMOrLFJ+aJN+eZ4hHg1eUQ+W8Q6lH3xo
AkZSj0Wxo8EPH4KNpFAlAOR/pi1+mbZ2HvYQ+8fU15GdyaBdo0DViQWs4kRtCAwp6rhja2FhJfHe
1r1PHKCQO2HT5p2YrZlNQz6w6RdLdzoFed8Gn4rHruk+st6/Qt+WUahl36v4Fh6HRHX6hc2YEy5i
/yZYFPzKJ/Iwn5VOov8eSmGyWieKLwLrlQUDcYy6LX4jAGVBCcVVx/FsU+GoS1zLUIVXz+XobPCH
3KEwIMiZ+8aOjNk+tjbEEd/lGek8P4pClsuFGcKSQ2pDXDez5nIlL3wOfVuS1PjFntfVIxdjSM0+
YkHHW2d1oh7ClEQXfeE7Xb05M2mMXPqGKsnQF9EpHv7VK/3tt3P9PApcUARA7FHnc3B7qFctgeKp
t34SUSkMSkufBTftt1M+Tb35aSrGAANHK/KiSXU/A1QctlEmOQLLWa8lU4cVCN4qSY9KaZri63HX
CtSnAv5l+XIRBmcjjOYDrHcY9dvpEn1vKlF8PT15A6/ChqCiryof0QplW7YMO4+Iht5qKkfoz3nT
zNT2/5WVTfgYW0u/ljnSSIlm9B7ZtRB1FiA8HYG4y792/MYh+75mQVYt060NxE3dNsuFcfa45chs
3IfsMAM9lX981c2KHMSgjgUjX83C4T2e9uew14/zIe+NiMMGEuTO1Z4zieB/2/3mpmD7RyzeaDDw
yWgxnYP2foBPuAigTNtRnzZTYfvgXS21/A/jpQI16oJlc/kvtjIBAqh5MZ0k6+aFI5Ht2/MZt36/
1Cw08BnFidRa2DJsALjqxb6yqM4Gb4v9ifz2c4MRgHgcPyNpiOovfyhNJD8cwcbkrNz3G5xfzOiG
1g4wnHRmXEDZ16qxXMv+5bjJogpEIBZONR8IVjz6RkEBOnZkMltvtPl1mHYB9xWV+cIWQ+xMQtuT
SMW4zjkRi2QEXx92duzJMEgQdL8/0rYyQ6ttyg8JDDRzREC2R7spLKtECm8/QlVFwhPn3RO80MPC
40kZfi+0Wopdr1EafBSao5Suw6RROLcNdxLAuFL++zTTss0Wyuui1rbLXBX6V8M9vBz8yZkV37/z
0RgOo9qKXWOqgfYo39MCs/NPnx5mfl1x43qbJNumNzdQgaV1xAta508scn2gjiAtI5W+dk1YKzFs
ElatbXtVDhyXXNvJrhHCpABEaXsjIAXiQgG3Ye1VpXi1zN9viPQEYp1YwQvL8hd1AXCs0SRClo++
+8XdW4Zebo2C0F7Ezes9QF7CGZmeFQbc/trEK0JaXUQAzAheJvXkJY/zX87S4NEGHjQG65Z4OScO
NG/zOsoPG3Yeo3OIY+dtEbVuG0IhdujglAMl+mwq5z0zBC+DCAMvxCaK3/thNyPevhTwaUSQ+rZn
yirPUkJ7joRJbaMt53eR1inlSbMoepRYf7H4Ash1BtMV8Nmv4qkVNBM36WaEP2vvpL0rSG+hj+Rz
aDXAJJGkGIx0Ah0q38fOya6GAqcnExInJ5LzUjexcbMx9GAbPphhJxDgoJ4XJ50kFVvp/pgymplq
WYnR0WdmBSBsp1ek5ud8Ysny0shyLfX/MuXshCj+ZyUTWrqly9l24rkAleXe92cS07TJeHIbysVZ
rHqZjbM/DhOnDaf+B0JoPya+fZns+fSZk3Cq3TtTztgcCJkhubQMe5GjzwEzE768/+m4GOvuyuH7
mNwDfqc0y0GdTrYZhdIs9zGKLKoMgnio0+LjmvlvEbo8G8E2f+nOk49CkhaHfbznpBHk++gRyPGw
S+qWk5B0Sj7Umm44B02ytLJmyX3CAwO/6t59ENOyXQpbs0SCz7PnYzfuRu3qBPNUwiOjPJVEehL0
Iqm4EQgunbbdYqISKRx42JfseknKtIMwxFEZ4mMj0qLY0eAoaLzK2Dp9v8V96fIrX2KWF/BEVMWy
Oigw9aVf3fcMHG5PlQSm75Z0Il5v5sfkq2Anp4hHvuM/eSWxvOWrsVq3kFHSpnI6PM9k48edwdjB
eaP6sq717hkSprpFprKxtq0pd+LFHuukZ6BZAmBaU/dUGJPcSsMbUBT1TUTDhzBVJA+XlKfhql/Y
Dnl4zY8nNxn5HU9xuxLS7+D/TzInfNZzR3gOEaiYsTwQdAtp/ypDlKo6/vwVsn/fjgjHU26DYwr/
bO/GHptHWNJXSQpUtah7CoV4EMgUKiUfCDj2O/+L+2FsT+s0tnjHihba/13LBglBD7CSyDnzayrN
hFIWWDIfWEbqn24iwaknbWZAmfmf17sgeTosArMq269kggJY4KVNYMaqtegGbb3k0gJMbisEfsBp
r8pGwAUYwQ0pl22bogaNYN8gl3ct0aOp4fhNkdnLY6hpBI63dQ1SoQh05F4Rd5952voSUAOazjgC
akCv05f6s++P3efNu77316mhXbESgHxg0omXIacbHciGPBHOm5pUuammcKwd/cJk2dD16dH9B7TK
MxlUuzp0JhbKcOCJezovHrq2+uqJTEixvg4jiPhQF5cQlLmpr6unqLRAFpkylONsFOkb6kXmTqol
O9kuNhN/SxulkEHlk+lxkk8KaEjp9XXm8wKBYq/KnkLS25hrBf72M+VEmst8t9CbR7tF+2OjkFGg
XO5vORUU/3onTLHhBre9T5oABRkAogi0E1dTz/n9EMHSSgwCVgN+WaSoOiRnpiF75uXbRQ7aCJ/X
kePE67D6qVhGi009dILpZy3pxD1sNj2cpfu3+Mk4Octz9wVs0qrs+exuWbqXNKgP8w4ygmIRiAnC
+Kxm8lta6y1ExdQN2baIo1/8IM0ZOtYFPyAVylEDE/HPkMnfp7LBuHcmAmiXeqLs/GQtn2qCtxdr
agxaiEUVH8FXibSq1li03JrxvoWsJeyff0EUW6Hb0giI7e5Y0SNLUqpq6W2p37Cetbo01JaI7oaY
5fyEX6lxXUZgGZGtVAi69srZklOFKnmefKxTvZ3UsS9Gv2ZTtD8eIFcgMX+QuCNH+//BWQf5cvfe
LkG2GieZj9m53Tob5pMQ4Z0S0To6ny7Xav+GdjFWaFzL/U1weRuYb5YdCva0QA8q5UlPhtmE4Utx
ZTHtdl2sEB6nrHlJ1Usk0ROU7qe5AVi85anHWsSYtgOJ+hfc3oMnK109RndI5EItbORNKH6MGI/x
N4JRv9RaxAcRZjct/GfH+a+u3SeZwz02dDoLQuD+1UGlOuyMKMnBuQoIbTg1xcdQSZnuAf6/ykZl
cF1cypxRgAd8qAQH33oIUecD9P1GtnK+HKqaZPQz9WdH6Wxpz8Dcqrx9RUFsVH6dCSblFe7KkML+
PB97PlQImS388sPGRFFOGoCt0vi5CKndP5EQpbvoFzGC1pM2az31KPxOW5pnYnYjDz0MHBunE2G5
LA/yf9l0EZxEa21lXNgypMW+MaJMq/0TpHwARGpWq4hDKcRXsrMUYGgx8cY3GYyq9HlUOy+ZGS44
DdtnZFx2fPkrmxlLJvBipeoPyvxCX68hv1hwCrZpFOtv/cw2XNJVYpN05rHcxPaVmK0t65yY2Nrw
GGXVZE+6AHTb9uxyfZwIJdQxVVwL0mwRdGExEccKPb72eGD+LmkeTLACc6h+d47K/BwFbxBLQv+i
n5kTdl7lumT5AD1EW02f2WGX3HpTt3Sng3TTU+sladq8oBiXJm4KOn0/9GVNMDr+QiApQyWvPz64
n6PlI/JRKuJVbEybMDD7ulq4k+F6Px1FNFKU1Mm9b1CX0LaS+zjaZQ5AoTuv9RZxtoIogE/2hGKX
Ed7EoVcDI0jptcTIMpTy9e+AEa3vCte3S2z1TYKZtz4jUkXRq9hFf5edVljv75dcbVwJd4p3W9Nh
qy5hGbneKUAv+XATBooxMZsBdnQ7HqxuUBzEfsYvuE49QTWyhua6ELOuUbQXGVTnRMj7Y1ZjGf+e
gcC06pC8uJVpms3Q/K3+EJuBVe3qhd9z7/0N0M7WUjv0P7lWtyNgdByG0RV30ppM6CEbwQ5taFkC
0pvPXh2p9TMlylM3qwuDwgIY0S5YV005oPJ0BEl4BJCXML3B0e119yRymnHu2bENBuiwU2e+Vc9/
Go4Afu6WCUWsp40a3GIlNB4wLNpDavNiXJiM34xlbc2ZTQWKBDW9Aub3uV3RiwQsRsQuKmC7G9kP
1SWOy9A/cqrW7kNFhSMTCUSdAFx1qJWhArxUBctTTSwO4N4JgvvmQtV5O3PJZssBeUZWUOw/BGVv
Nq1zfJiKk+tgNA/bn0osHo5vhNSkxUYiUSX/YR3gtC8K5xzzk0qjV0hSLbMBwAa1MoABCnMV+V1t
4T7CfmbdoQiHbowQwOPJ9jyDifD0XMvUxU2XgxqDqFYwT9obgaAHKyYEQOR7De8ZHBEuas7SUdFE
X8et4f0717NBrSy6koqCzn2rQCnHKbkRhxlDQG4HAIMgvfLcW0eoArYJ7LSjb+jc4JjKjcS+6Pw4
C3CGYaPhP1yOET7peNsnDZmiXA67g++RkfA3JMY5E9EB+KlLRYiFEWKjRd6enFUGRJwAt1A7JFax
o4LRGlUz/9kgUGGTPoeUL5pSI20abqhdDAQea6Zwje3AA+jCi/53yCo2chnVG1nzC+Wejml6ozD6
kEJYnBVT8acHfB2s9Cxrqdnf3+I/KYGmoCOuCKYaVHhrj+4fmM26HgedhYPM6pN8nEZcQRyKBbEr
sqsM0icrnbEU/EngYNIW1ovLr2xlgkNyNom33hrlVrDbpD+iWZ20DbtBHE8SoIFWI2yrILxQR7/M
JdD9w1cAl1Ybo+eFEdZCfTQV7E40MJoOgAy6AJ4uJTc0Zx7krhFCQ8VDcdYXZLwJxd7iyYosOxUH
H7R6N1uYErRCiHlzb8AsveN6VPCOiYptWEVxVLNvx9yevrkvuQPfHGWIFeZmBt/gw83VxCce+C1q
EQ7aw+TqoWdew1nZoVhYUnNAL41ylkH4zOpy7IRk0C/n8ZAA9Usyg8gKAS4CQHk5Egra5xsSHruQ
06GaNYstw5CgjerGr9ww7q424Wk9IGcea9VEOBSeIJcZYFfr/WgRMi2N4wkVwlKHP1GVKmNTuCUj
KnABSbY1ctsKTSVbvMXuM9KopmxKtzaC0F75A5VXk4mZhTR9pfahc2UItL+n1pBF444lMCYOHmEr
c7ZYKNF80cat+rNpqQieEs0as7GlgRx5L7sivMH19jGzWh2/jroOPBDhMXqgHSXzyAorGVZDtLU7
AnChTr/9L3uUU1vdfu0buJkKsrwz1aLmHGrip9jv4Mm0jpMoVuyV99mD0inLgP0y2KIzl+NndbBI
1/60FXYkLSk+UxbXVXtknbakbFR1qxvjRqf+OBJhp4BSuyuu3Tsqry4J4nrcqh6BmgZ+w1dSn1Gz
ngAzCG1uy2I6uJ5ZdpfyiiWeSv5ukQZRr9WwJvtPkWNng3ugtY+llfZ71TYFijd6TQJUYWWVuW4S
HOfPN1Pv7tA/r8bZc6B5Hb59fuS9WxPyvY/UNL3RXd/Sdske3BFgfp9K+A2KVEVoU3MlYn2Vh/BK
oXc5M7RJ8/+fPjTqdnT5/ivqokjrNnO/VMX1fQUOksofaiOVS1IZ+dd4D+L20JPSINS9unGolGdF
PrEaxpQI4xdd9WOttFiem+v8FqL1JOJwAHX9F3vkxFhxTO5SYDO2dlQwrjr2W4wAgCu0HuZ24csm
CVanl+Aff1TGJ/7UoZYaeB4gKB3JQ9/TZUiUYedL29B0m/KAtzXakfBn0KKGNHHM5mJScD+dbMuC
Ot/vh7GH4D0VUqcfDA6vlMBK7cd8By+ZdUVH/GAxWC9v48BIPTWELqRpLd+9Hgj9GAJo4+pixsDZ
NB9voK3ugspsyu+xyQpGgfeOKZzMgksKFwfg8ogK9sBJEExkdfMqHN38bXQWMj1MjNRGe3Mo6qFO
poQ90hztDy9wWRbbX5JhHTOowhMGgevxX0NWbSCRisX7oFlCWRQQtRNbgtyTZx62buW122BEN3WZ
NxB1IQ3WhGXhiRFgdSDOkX5BzNIW6UoskzGQMCmreUzhc7W79iAhx3BUH/0uYL7ti3qIYar0JzDY
H1PBF3zlnJsn0SKbOOfyI1T9IUzeZdedM/Ww8747uZ+cfy32QQegMdsAC+qJtAgjrB5bt3+ABvVU
X1O82wHl+cqQslMzcS/sEF13HJ4y5lcd64Dds4zeT7ZbptbfJXOi+K4UaPia7e9cvtkpO3ZA0AQi
AWVovAqpRJzIH0q/bdUPHQA1ovi0LU8Z2u79bJW3jlbShADzj8ulkqNbvjQusyHYMg6OTyNjoe03
3DKySA9ljOoBcfyhamB9OJ0wbbBxkK8fjNYg7X02fZSLFLLnAKd204551Lt9KM98C9gNpLiKr8VS
8prE8H6CMhk/NwL6FoL6ctBv6S5qSBP5HcGt17J2xPI1KHOqgVoiiyaGHVhsiwZN1dOInsWeLGr9
D3KPnZO1oCiIjQGPObELSa13piGrrLoGRiLSCLFoHPK1fOr5hOKYx2v72qYbUIkQWacWI3h8mkZY
P9AM5GDsQIkc+SoHdPML7D8wfehtSxA+AhcNXQDbsPMc3RvwjzjZgqVVDFCyE0++t4UBfywxneIB
qVRHqsrtpLAmiOYAMG+YAUYCNd+bitUEUvXOTdYq5u6b9wEC+UDnuHGCuN9PhiGbVZ0uhoX93jsX
4QTxvx9491EXZ7OXU1xXmmG71aNfUruvOEAWvE1ThbzrWTPSjpoPLonTJCxP9svqJeG0HgnxjuEV
2j8Vs/02Q9EKk47mYlHHwFgEAOpxkVbHLOxaBfbrWc6Y5Xy5eclI4MBlwVol2HF4/s8DmMUShUXj
7dObUYy/wTveXh7itThxnq3rV//d6gOAgTmurcU6nqZEafw2DLZDHrr6DvXZ7wJcOE457AZiXNV4
ykn+RnT3xR6U+DaFv6Rc5HDTEn37DvZfsaT9dCCfX5zw724veB+ZHA9RrMqzsSDQXaYTROnQs1Sc
dIwAJ2X+b2u8B+OSoQhxki2GMmIVIKHPRCFIDb6D5LwC2tAJp6claqNxZkI/c1tSJGA1yO4+bIDC
75hgRVLdpehauh0QAOBgKN88cXvrJaGnYpiPspAbi2jOZ0UWpYVSYOoPhHt+GG3WBduvdX8Tc9k/
+ev6xAvGB0DpOiLn9qtoretUrlizkajhe1u3PW3t8B3YYrzRLevUIzUSVuzcQsueCRkeUOJOJdwe
Pwhb340fpuLlY6DbNRxT94Q2ImXFhCeaIOudnZkBDw5VSRACTzQujM5Uhkp8Y5Gv2o0qWWxYj9qb
7bH3PtvS0ar6cDRrEYJw4608+Iyvv0U9YFB1/I5Ga4WOTqWDdsL+52xMMkKdHpdpirqpf8NneNrG
/xdqteiUaAb6ykfn0bET9vNX86ANNEEQd/d7Aqb0wg9ECxji5N9HbBwvgvS/vByH+FAE1fH47Ytb
aowb7c9sOl3zGySz6GDP7UVWY5AjlUbEvnIdLjCIRZnCTVZKtWZpPPhDOIKE+74AugPl7TADRMyW
r12ZsZhlxi+cs16ofEan3OlRYnc2FgbbeXQ3OP+gJi0bIucamfX7t6yZ1ewI+q6YOl1NVpGcKqQq
zeKZg36Za4MWKWpXPbNlBC5/jpRefW624oZW9alF90djXwWCXJwvv1rgRSOCrTVv/fpSTbFqyDNG
nGxApi//fkCj5FgBoKpvNklVk3WY2f8g1mPUKkhYKkJOXBdaOHEbWxIH60LVdTk1nkkSdvBOakaS
kJMrJ4yZfYT1us+16qcOqIK9WhLlkRsvHogD5ATfRCrE6qNTyK/JtQLZk/QgpLXJevfSqxbbjxuM
Tny8tZrFhAJATMUPOpb8KaqukPgE9YTVrYmo8Bpl0mvw+1lFBFpl6Q+GzLTR5zqfY3eppp1Hkcpb
16+DeLnZ94C8zTePQ508GCl/MSwQhyS/S659RN5zK1kKaNvFZ036x9/1UFd+RQtIFG5NPimD7AgW
tJM4sqbTjuTGUBSNC80zmcWWJLbZOoc63CsfEFd9raQcsZ8eb/pLfqZYCGsR33CZgYEx/OtR98iY
1Rk5Z1HvruBb90oXhPJBdqg6NU/dkql7LB8S5sgOPJzu67G+sGyx/KU4oKggEZSfaW6B+EAhmQg7
XvJSxnbl0mBTmvtsuPxCUw2lcBAApRUe6a6Dddlh9l6aFi9yw7NGLDqLExjuBaclgCKvA5xKHGUX
fPiwxBO1JT2pNErSTSuvs5mznOGu4H/OP+qUCtu/sscaF2pxkOGV8YjRaWPkhBbiY0ppPd1Lx7Tz
PpQ9rSOnbRlCLXbrmNSakRfcubl6p12YPJHdMOE2IAlLVSzg+yoBfKh0CGTW6DFav5oeUPuxEoxU
hywdu9LlQCCN5QvtcGUtiqKh4OeMg4UqrlulbmeN1p8yE6EjYuN98VSeSg7GVC3cL1d33thubb+A
/XwKSw5IdvCbjUlhdArYempRM1E+nie4OdlT5jkjmSt8QjflLY32fUOdoZSE5MUTLF3CQsS7ZdHs
NxMwJ3ZGzrVAamuFLUAxRFKWXHUr5MfNu3Q2HBNFhCXMisRokRrOVZqaKlnHtuj0mX3ONqpt0XQI
1FHH9wf9mTJ4zUBydq/zlpz2UJoaR14aUTS7noESegjia7Y6b5ztGUpYP5wm+irCmLucnbtoej/a
/xunxyT1NUR+pZJhlhGa5f6x3gsEkt9H9yufSVqf0MzgBsXP0w5Ixaq0aKU81IJbeI6KzaiM1fqZ
hZaELDwYCkfB66SaHvVHWj2zu/CAZSA2YmFCYUCXqpS1v8QMEntmA8YI5HwlckVkOGFzE/kMLpk+
TMOMUKMoNE+9BN6fejd0WBNWJW7SJ+RbUY+HzdZWVCcOeMaOY2DB2iCrnmltT0K5GxaooJEthJVM
8DSblpmVlcQU+/bPm/3EGWufy8avtkakw8HbAk3JOWRwCpbHmyH+H7YXc35OMRxfZRZQEhs1g3Yn
G+hYcDPRMqmqyyweL62LSpJgb/PPinp8cfn+bXod869QNXahUEumG4i4zWk/zW3Dcfd3s+aZConb
eR0xzT7WFdfy+kr+x67pzFMxzbqSqun7dbpBhVyp4+QN7RQSrTf6Cszjkws+1TB/ut/cpG+KR8oO
XwoFAdVWEsjw6PghlS003y/d2Lg2VKPDOVGINxL33DFq0BO40Z/Ujjvccoj8n1Z4+G/9ArTYPpAj
W7RsaQ9Vik9I3dbrIlCtVfwxJ6BtC7mg2RGLZTyA9HsKZtZm4wDwyrDnitYg7wbRrQEBSW/aTMUx
ISl6IDEOY3MKnZYwAT1CUGNPIipccFY5dayecWJFONliXP6fHz3wBRg5dwZXaJQIDkbN48wVQV5O
VLzwaVpvD6BOiBaQF68RuASYPFVoQbYofG1S0FeL4k9CBykWvkRuHVPnjN618C8qyevKxLohvnk+
4xcK/JwGbITB9AqlTbkZI3CTVgEOavSki7EuW0JjJcB29ZPvIGAydecCJ3bbhxxFkop4JqcK+wfy
ZIa8MwcQpPNljEN5in1CfBgXkMJ5I2WmNCygoojkePbcmgPKuv+nsqLldPwrLc1pbPIZ6mhBd5IW
6hzYvqxXH8j+90rFZHb8CuDJXU/4ioI8hWZYJZHvIdGt/RqBLbhGtnvUUC5jLtb7ylE1157lmxfl
Eliu2LBdpegryimllOBq8UdYqW+eDGQjG7yt610202C9j1WrtsS9rsevs05/8p0QolhVeKp5vs1+
Y9I9OAKUqdWg+avNZlZ/2hDKAQeL/EHFbfox7T4hUjUeikwFTgKtAjuDzRrs4jeITHjseqzzn2z2
gZaKNvgeHVl4a7iTB+L2mIIalErDxDRzY1OxR4CoJegsYIpo8A+JM7tOij6bea7KHa9kDn2DkRvC
ZkNfAqB2fA9ti8Fot1mtIlAebIxKvdzrP5dHo+qYHqRdj6KFeGc0FTd82XzMAZW7l3t4LBou5kpP
1YEaISd8WcObuXimwrewEWoti0NxEOEHsOz5nexgMbT9GotCy/BJ5t/mfFkqMzxeA4mcfKU+3Q76
feDZh1rJW2Ep3xQerRj7Szy/E6i4BXLn9YYhWppXT8HEAs1KxSZ0mRoXQocXfJ2pA134aYVmmlCP
l+nM8oF/2GPYPWOEfXqUWT28ZiO3mkzmBRE8QMO+geCst9V9NzDNQwf2JVWm3o6KQToDmONDX5wW
22//zAKnbkhLVpSGpz40AtoykPXx+RpBvgZm7d6LFTkSRBqdLfrhd/qxyVVoP/UPiY94IF/0+X05
paf9IMvD2RgkH8fKsy01PhvUZqQ2d3W4Zn2tYsgiyJjaLkf8KRI5pfdhuXPjqDMoKxQ+YnkbOtFg
wd36Gzy9uGSFDx3r6PmhuY/umkawUMJH6D+R6UXalRheVrB3VYv1vfpImCciO5X2gMRDeJ3HHfcs
LoUr24UQjoRBxFWUzCyZXm0IORfMdyEvp9PgJFh7OjUAIzc3Lxz26rxEaZhNG3o42sBEYkOU2WiR
6y/ilJMkhGANfvQFeqfBDdVjQVZOfO29q0Cs6qNY8n5zRZwDjEnA+LtoM+WKbHv8r9KfrhklqTxD
x2nYHG/6z6Uca6c/yANKG2EBy2omABIlh88lnsl+S295emQtFbrOA7RxrEmDMFGdJY0IQLAf1zjy
ezDlPNifEYAzEXT7y07VKrtCXMhxwAMFkiOOmOOCJQ60+1BwsgawHv76lhpWrJs2Sw6zqdyJGyy1
I27/Fp4mY/gK/rho0/V381Wp7NTHREYdFzToVxCPnW7QKlqNpFrZRlNT5q0xp36lEN/rHE2WoVn1
gz08F4lpohQl4afvqE+w3NCn1h8E4glhuYYBNQTHOLds1+rEnuAes3raNF56eRSpn+DvKRVovn+I
szuhDaNvp9PgvXNdRTKZgEOtuEG8xfz1xAHqsKO7xViSypVzh3Y4r0pvIWp6gY0b+3p1qIdOjZAj
q662Iym3SK2m+ahmPD+dkg21MvCPrSVutsCqcroay6xKQwKNOD1OehP7p+EE8kEuRJD+Jo7EXL92
C9RMdCDKXb6Ko1HlOWxrlzMFj7DczkrA3DSLwWXI308SzrItm+JfnTsOYNHmkQxaWOaGDHN0F/f3
hHmwO6D54n4lVr/gfymw1ZX+kD4e2lUFcMsBrsV80j81aI5g4MXfQh3TZeUIDzaX8Y64Mod3Fd5s
q8oj4Ft7Yr1iRiLCQG6u7U84Z27hkz7UpQ2JEcal/ZYLtodVFMaLYNbx78Fe1VA7DXDrwHi6X56H
QkNiQls015JKTj94WZBM+fjJcTqZBG/qu3oSiEuq/WQKj+R2vYiJJjScX3dfmrqJ/U8MlgtGIroR
OKmmY0m1kCrn6BZSk8V3RpAoSj0yOose8yjrbPe+a8hwcDx9PV26fQecHm7Z54B/PzsE9g7d6BBT
eU7RSkj1O4treu9pc40NgIM709whrgi3scrYHFu2jlPL5f1PRt9uZHXsEQRmzx0dewVgGpzWuSja
wGxiCxz7brlUfTHr6ve+B01Z9pzSg0nUxNwD0S4VFpcKnsYFO34aGVz7j9bbq/I7+wscaEiNWJhT
//fLIQ7vq5vCAPTjiF9fLc0WhRpP8PUaD0fZpUt06Ik5T08x9S4aGvRajEcTQWWIXhYVltXMR54f
buXnZ3Nuc5JRDTvAp96g3uihWvmbCuAbw1Lempslh0HWNPgNhVOQH/IETubMtDcaRsC3NKM2dmgd
0K9oXwAkp6+UI5Hd2ya63BOcW64eEBNKmaauR0XprH6sVjfrZDz20HqEoGOhTtmHKrAMVhRcTWIG
q7ynZFnrc8SHv3urlflK7i3sG1BTqFodttJ7xOtVt15cAX4R5R8naK7w/lw9ru9U5vaz2oDaZyPT
uHRz1rqL93Xcwfsm3n5IGnwkVrFkdy0g54fsQm9rc2UhnZjL9rEo6lolLK37pL5KEfNQZjNKNRyC
+RJHYj/qKVZZNUddVzGVfqtEv8dWDBMmqJm/WGOdVjbQPqtFZhv3T6KN49v2lu7RCNsxeeqi2qm3
ZX4XNKDrJspIGaLPAu8DIUxWfek8XtkhlIpB9lYEC8HtSwe5h94z057AVnN+fJ54R3WypRDoqXDV
OMfTAA4NujTeMeGfYjABkfYpsIQonmjE0vYl1pGoKZYUYVTvsAy/4yabb2iqka22EEa04TvaHb/z
QfWaQNldX7/RNKyr6XH+o6X06+dXT5op6ZK8BoWVyTG3jon0zBHXM6WLVAnEFOqQZwsjzvk0fL2b
F6KPBxw83QLZNwmfk7GBG8W3rbvOu3c10XzDDk1BSGM8He96NvVCRAap9eEa4r7/4e0326Bpo5O6
CmRzjna13yukCFHcdjl7ZO9Qc99ZTRGwkwmXq6Pj7Ax+Ne4La5fQGs21ODtQhfadlhpboZOjBGT6
tDbCkOpdq1J+TKEqn3n1u4dSCODbeTPf69Bcq+xJbYO7Zg4sRgX6mU+HvAYyQmRxHPv+O6Yj9dgl
24j9eoUvzlYeXk/yNAEsAO7fSDtpvrVT/gbXqiBMnkitzbMdzMY9yJUOfGuW7Dc4qK9wjZ2m5igY
jA5foKSsCvm3gPw+FgTttCo2Hd/rqaar1VgGMNfAhHfYE2PVBqcFlvkD04NaWwETMM6ggntKXXVc
B2CvEDj7XbMjJO7l7nRO8qNdfcdb2V3PxWmdYJC2QKQq9IhzJlTYYI2a6Xsex74+3bEW3ny505s4
VR6f+VJinbkYStdDzybihbQsThdZiTLRcwk36UigLpud1h4qvaNQLEDd+n1iblKeO2OzrZSf5yYx
oQHPahUvT3OlFzZ+hS0edK4dQc3xZAI5bCcL6RThXilghMSCzo0JtJF3W8dgzu7TGBE85s3H1qZi
qIDvBzTcyQMNBZZh0RJ4ILHVXk/4q+Ah5YbRZsHhP8j6dalsKS7dEGHSj0rRkpetfCOFi9aQYKxB
Npay/55i8fnucfMb3uTSsyv8MwW/RFzlJUk0nP9zXW56Bj3G80cxQG7bQbCM3MFvGH/ccp3TKYTY
ngLa4kCDvIMicH9bpjvowY/5NjzCfwxw/IyfdUUEo86xi7xgiv39LkxZr+WMpH4pnXIY9uyLukno
+QEWQdNa9+RNKdcqheXT5cPfYLpk/RPiePaM76CRaP7mgSp+oe+FvuMPvEnonlM+9Qpgv1EDXh3N
ZSg44Gbp7R+buVhb86vGo+i8Bgc8fmOkm3OObSyuG6rnvvVYvSpopwrf6aVuMJUjXiRcbm9eCiJ8
oTt89NOGgjM3eY+O9Se2dTlA2hWmMju2DQEGXulG+hHPfJv5cx2n27tWgoN2XeHjECiTGRVRnvqN
3B3N4bMPk+OhnxbIh2CfdXEUHWgx5YVIwFtsukcbSoKUSTsDKFu9DmpQfwCHlwzt8AoaMyQBvtpn
iQuyJikNHEHAWAP7eWb/gLp6HRsf9fBSBtSmSjgyFgD82UdFW0xvbmnHdvKuOFhJg5dU5hqR5Cac
8LCunuy3xgnFrJGOTUF50qRY2ESDGfAmn/CXR5hsq1qpFfS3XRvx/glfwy91uGa5StKR2MYPekxt
CiEjcddpsREQr7gHFvBxiaBPn5guX4rzMsrOC2s2XbYGD6EXcHpd2fn2WTWqFcShe3sNf7K7kYNR
6jqOPn8noHmOMSAlfoxZtQI/AO2x/2RkXKHBn0kEl8J2pLc+54LPmL9GpeY6VdAbHcQ1Pami5Iet
QZtRZ0pt63guuC3xOVEpUTCvudZb9169rAUFk7IWKQ974wK9vW4LvU3YJrPmGrgsWJiTIx3c5YHR
6zqLFYzhuCterAT6yxz95zXSEnUM2n/yxMxiCKRL+3vLpcaU818VzzVDR5evMqheTwRELK5JRMTJ
dbrJajjumWIZtz8I1tNDoPAfbl91iNjCOHsWyVyjvVeHfDn5M0datRWAgjy+L5PvsuxeDYvxPJNX
8HTeBUO+aUdvN6dKKhAZUuEJiP+SgCyLuC5RrXy2/l7Yx+x3xNMmcHrYJiOCIfhtm72N6c9ZuBSP
79uD3I40gfLy0ebweVavM/7khWTQMDzDoYnyeXSIqZh7EmRoh2/aSFtU0+J+Gcqqppy+vrU1EAoO
+2qmGWZZlrLecNNZFdVphxtKGvw+fCxJZFl6EtBBiCPm1BzKpahiL2Adq7OfLs4P2jAp4Dw6kKPr
JecycfBBAHKmsx3qRpGjCvYdsZpHxxsmNRu+rjWBjC3Ps6d74ACtrrCL6RKvWHH3HZkVlnES1X/x
ry9Iv3UTEp0GiNCYh4WPcdkwojl12ZiQ2crWmtWK4S111lz+WMJOQINL/ONkMWnIoG2SnCvieIRe
PvXMLloxUqfClBxHEVvgMJeGvidgGJnHc7iPBdIw1hEENQdFhPmVDEepJ9OLYlR/6RjmnwNeAGH9
Rt0hTK9zAkd6++hlksuo3lqQ0OY7SQlAZJBY3iMfNbDjSp6A2DbX+gOJTMgSvCMQ+pgUDVDtLOqV
jBN5Esky4du42YS0cAjeglfl/tAbhyCwcjOT4JSj4eumCy/VNnRIs6S7iyYhdBNnkVEM3jvFoY12
BrcmtLbv0sVSWEFCBgOp0hDxBp+UfMAY4HKtdBwFvksk4Z1enu2x9CmFxgFk7VWCrKfZ+/ALREKk
RWvTN3S3cTXluEmL/ztVXCLOLoEmLTxoTsZv5lAeDNPHIvIokjrYmzMHWb/AFujaaiKMQf5UWRhE
qS0n2jxamh6xuFw6+i2xkfUD5PfKEgc4exMlSpzVDHUFEVRPKdyN5asCJ/N85gqCCitoh1F7E91d
gHcTd844kxx6RxVoSCYc654Eit60qFu/owvttE73YLoUaUxktGuV8XBLIRYiyEfpeCsO8wjCGKWW
uOeHE0R72tSmE22USytcVyyzpGZaSS+pXxSXF6bUSBg76AbgZEj09L5diCh9W3E7bvB1rdmIezVY
MxRUfFtVm5CG7Jxw6cJAUX2XtKJUcSOu89E0G9YNcXYgadNI7CYtSWG2b0Lr2mqNYBxQkYpOiF1+
EoiHXzwBtRZcEjE4RlQClvGc0mJxqTqbGQO5KNpOegngwzy9zTPv5R2ijCVnYY4H4mmycGKq3lqH
tOEIv41BU8yE3zea1br7uB5FY1lFcyJ4OfWHCg7UC9Iw4HErut9c/sm7/Mnkm+2jay4XiVU2GJ02
jPhZWL2WuTyzBUGZMua/+vNQp/ErO+Sffkbe+zc6Prh60k/lLVr3zBM4LzFer+tBKv6+hyUCzcEr
n1bh9ro/x7Lng/NXtJYuqRQX7a0paO/lJGUGruvghRprB/DRi0/RdwQC2vRjYfpudKc0gGZgCyes
tccSY3vFI4qDRNDgn8nZlnE5rFkpegCsL50HY692SEZ8NSfO8VjbbK7Nn8bDaJSH1+8bsitfQfNf
8/TKIhDyK3hA99yspkoAhxh/uwjrD9iKJW+l105SwX3G1Tgf2Uh2CtbKYyYLmtUH67sf6zYAwihm
wOv3QSWbBq8qJbKI5TPD9PUI/d2H2mGS9imIlFxKB01gfyx9Yi+DZEfeJtD2bTaG/L627ex9Rk9N
gf5wOPdIwwh2OMVi+boif/PtJLWK15f9yf9R3Xe3m3EF4uN3YPUq33hYLAEIBc3pzB1EW25vwpxx
hQ/LJg6FP1ETunl8h4HG7iGKjBw9B4oKonP0DUEEiHXPEn6Kc0rcA7IRl1QKhnVdIm6FnT3YhUwz
gkOHCxCBaiqpBTE2TVfcOPe66DFyryK6uq14TISt9+jw9aD+Zaf5X00jAPOk6NpWyUEOeQir8jK7
O1iECp02Yr42UW9JSAXjbt/9N5Dl/RaMio956JNupomQ+wPA8VS6WLRPS9KBSKjSgpd2H06bjpzE
TwBUxnLOx4sVagEv/UjdVkEKHeihaEj5cI8wOTTdpengK7NAWjH+ReDIiRVI2tYH+WqJj7h3JRR7
AkTpPS1GU3PLuQZqk6BD1Zgd17FTGnIaaEidX2nm2lqJ8/02y6zO5RBiOIn9ZJNbn4OWBk9dHSSK
xF/kKd56ryhb+xWYuEdZPAZZGkcdBlLpDEoX9sqUBDmNkDJUZIWIU0nQ70p0qBojzhzfRBil4TpO
AAYdwYcp3Hl5MjhgAmBkzV7f9BcqmwTcry2WbVpK/vRKgzjehZqCSDEZMn3KyehkyVMHA+KK8E3c
iiV5CXBt6cW9Ng9Ol6CO7rZ5r7cRAKyIi6klGAQtNfMxI6SDbrP/9azNKG+Kkcy7CBd7BaO6IhLT
HhAsXvKl5dtHP2ZDQLJMFhVZN3rLCOutMfJ2fsYmxw5ZqU8qiTWhS20+j6PyE7DuJGExyRkWebpg
G+6CAB83mY5NBzJNfoiygnJWqyZO4GxBdSyxyAfEvvCKXp4vnDGt6LNVOKVTQU8IKPTUxSdL1X+A
Sw4T5XIl7eJU72La4RN0BspMaOiZqtcbbu38FfmVW6Co3yK3UMAaiHJe4j7bg0SIrnFfaBaojTIV
EJrrBA+DGrDNHtFjqT7N+/805Pcs/2G0JjqkGHoHmr2ubTC9ainalCAFdkTVGGjiYJSPNBT5DZfQ
6SgKU8ItyDL6RShuYplhZXG6sySEwr2pH+39vEDTbX0qyxURlcpKiSHT/jnank40DNICT/0Cb81Z
wDFuCAyAE36QKXC+c9DRQOlqVYWZZC99wkAMmGC6RXuVXVNHEuBPYWzZmwAYMyeG3NMbdVH6t4gg
n7zHr6TYRlACGt2v8yvWPdvqOA+m/X+VBEJji/dscQ2eOHnxhkpCElwN2lqsamYtzUJ5AtE5PgJW
/2yJA0GM6xeAtFIg1TRutjQwbUBSvWAsekPrmscsxPo0oXvBdSu9PgTRcOD0Lq67/Ic1ELDvd/Km
g6TprZGkBFl9at0BjCIJlJMK/JfKsBFpFXbqmV7FdEefkM1fRRIzuj6ftKtc97FDncyFecEpmGbl
NmLVn4m6eOTssmBdnZHA15SSgmhUjl3HbzU6LRsZ2gMHBogtWe18za0hziA/sOPF3/nT/VDYUm8I
xuDDGbKv975w2+5JZ88F1+sDXIe1MdE/FAhhiF+iWeKgXxoWxB0Nh2pLGJge0hivZ7Jeh3fofn8y
eADtBrUudm3yPpZKfdNLQNZrlxvH1qQAYEzU5ie4E/qaOmTFpA6ccBIysCI5GAsW7lLxsX9qQ6+B
mqUWzF6yrMyCDiZKxA8f7dTM1mJMGvuzYhXw5WcO4Y4I4S+shFUc/XvIGKpi3aC4p8I4kP831Tsx
rwh6dTQcvyDTsX9hBZ8jwWkP8zrj/fluH/Hv7EymNAGXAJw//a1/CAyF7YQB7olotsPWSLEKVF1y
p90K2uDHUjL7421zuvs5sD7tZ0f2F3Kl06q1NuuUzt5vGsLpFB3kjBfq+lletNMjfGUDnE7BmL7P
hq//AA4EJUY8Yb22DAedu7Chs0IQsvGj6fLZ1EJr0r+u1OD72lINQV7bZ8XZXEYwlfC4kND3+RhS
zD18uWnRqqUXfIRSeks60K1TurQj8JnEQf/5VSCffUT7Qa8EUhlaxsGMNJBHZ+NCyze3EZaASne3
q130WZwpKxaZ0idyuIzDGulhzNBj83easBf38DtVv8COD3pwLyb6zwiPd4TZSUZps9TxEqIRGjFA
hjOwG4VuLWRpLl2uiQLc0vQiq2ONJmgZoLzNtXSspHYcBy10SwXrASfd7OJF5VpqBqwRwxkWEuuv
7rWmqUvjosiJgMsOudGP38yQD5UvkcBZJyJLix7W8VTOkCzbRZJQwLLf07hZ5/wfDHntscgvxAou
vif7A689MSpyf+xI/3N6THkwg0xxCqM4bxF0/Fs8bTUeivtOYjwjZMvLNvDEKrskxR+u1W78AtgG
lZ50VRpAef+M2hTi4MEAxo9XItcWUAu93rtxHCBO3lprjhk8Qedv1zux+rA7UZzxptfKzpvGjfgm
LQ2p3aanm5W7b35giU7DFO3NABr6XBjES9MyUYnjDmyFKyzR2QGo7NVYJ2wouvR89gQ+68mW5s6+
41L0iS1txKI38UmDbIvSS1eG1a3fWuw2WCv0eacPxsYrPgEHJ7Qzzd71YmvjSmyxsEKuXQqhsu4h
Nxtpj1ISiIMb/AV7zcDJMKkhggpHu4ecVzLhnhDnf0lfLCzMiuz37g6wigWWC6rDuVtga2Ln/19z
HuCF3/ceZXzEY5fmpUR6uidSYy3S3PHuoSNwaWFIIS7qaT1t5ASKpLPR63Z1AxTHG85h7J9Nm8Nj
GuUxlGEa3/aS2J0KtmArp8108TOV1Fse30bl05ds74rjvMwXMEiKH5Ng5cmmjbaOmh/SU0tWz9Mh
GjSGfamzHCqVU+1X+6CEv4C47exSaO281hSpBO2cu3C9YmYprzrHIYSlIn2lM8HwqdVdwFG+rJUv
/Yx1RMvtBGbUEyu40cQ6gs1prOzoJC5ivtgD0m5XNQnzogoOJ7sGmHWRYYLHPMef76qrf5nVxSOi
j5yJJ6Q2Sgus3KhexMxcWua+vmwW7dVViv5tC7/cZWcYc6pmvoLqtM/Uzy1rHVKe9pm8HeFAPfSA
V+uNguHi++jpLI0cSNHfjNTU7/45yM4jUt3VkISEiIrzmfmWSbMPrNBgnE4iTJcQ5qhEUMGrEJwf
3sGxOOi3uJ+nSMi0/eksPnUsLJBtqQBeBE7LsddTvKYFhMWGfOUKt+f/Tmi75aD8MfHSSupSOImA
EczPE1MwwYz2vRkiTqdZq4Z8Wu9c9fqINk0bpqS7C0QGl8fKs6Ng3EOa4YGmUmW/NxNuxnQHmWQ+
GiRh5x0NnZ2vzkzp0h5JGzXUKG/hbjZWB1CgxyootD7k32lViSU4iTY/4YWxBZ4jDMUw1iwvlMp/
iozuwDWrSxS6DeMK6dQiEoiqUIGzzbuXRB8w0aJ+cvJRVZxHiWs3gpNTM0GsMtPI1RhuWnuJJJOR
gT+Ku5cOBRFS3/wJpR/sFoYv+UTgnnhX7nyzWOZHhD2sha5bIh7x6Jw6bDgjw6lVSL5zpmcdSDLB
DMBsBpzY2uO/bnFgKRPdcWOhOlqimS5DL4yV4D3ufK4H+rxaNdkLYfMcNJr/QPRiF++iCYjxQyry
3zs8+9gbm+V4COjAqk6DYkW6zTYATb6gQnOPf6kTdRcyVr/UuHZbm8Fow/+sJ5Wolq3WDEMZZdTn
KvT0sRLvDwU9ZDKV3hxDIMIBamtDjErblf5c2MjTjRt6MpejI2KZs0L4k1DRDO6zgelwRBfZ3eLd
jjSp7Ndtk278kZJiMztVfrXC31C/n1NWceBo0MSTcWC+sBHgREQkagJHtPyMFKy69jjdlFePLXVf
wNBfQzY1hU/FTTcCV0UI8EtaLxK28BdkncQYfwf19YCy3DwDB295eOwkFbdpbIlqeZOiC2VYq0Oa
2GhSJK7ovb7dN14jb/QyX8r7YMya9ysgkdDiaKyZUPSPjhAS1oFdfiyfODcjxb6mF5cBwhPHNrYU
+J0weRKXE8nEi6ONf6Qc0OdmDAIP7N5P32piJoGa6KRAU2picBmUwiJGxzNr6jTz1ZYvpKo+htzd
GPXpMIqhfi3aMMHclztNG6BRE05P6og+9k3hhYEhsn/OjIuh5Ny/sS69a18ch/Z9/zA1T4IS30rG
FIRBg54ZM9jQdsGFNdRPLCNzb8RJf29+gw6y+Xps8B8azxbhSd/lKLm9Zm+DtixplWGBn2GyLeEg
PUzWoerBztW+u7J6/h7Vdq/lZPF/EoLT6elGgyBEIA5rLCswic5jfG0E/IJC/Icxs902qFJduYh4
0vdLffnXOWQyZAsPIQZfIU9G1pyqx9z9UHZn5W/fc8z5Q+8l0Nham+2DlngFgNHKxsveAL5TjRA4
WWcQTGJ9c8SuQEkzQ2ROaE5TzePuDDt0/uzmtLLalvrJoX9DiMg5ehDvk1xM5PD4HF5MdlDMOdiq
nNPuog1Ku04L3qLexxmOBwbknkQH4suLqzApBQU+AokvXaeFnCkr6clvUNNWPA5fYgXM/l9Z+ca3
wEcbACAVaVrk/WCP2JRkMx1cRHxpDWsGiouNh6m6K7x0K8p8+3fr/kaD91/YLeiWcF8BaFLc1qUX
I49STVf62SBVzo+KRKJRCZNSNwnAp7Zu10RMy2Pvzldd67IX2+BqsJANr80AtnT9DQJIGFh1sqKc
tdb+HBbQZzMTanOePNW9dXsqwlI9f7OHUsZOCnBJEuy8m4FwcApFJuj6hj67qy0zDyjonRpfycBP
jHh0jkWNxztgbOpOBs+7De9Y7nVRvwlXAYI0Mkkj77W8uvYpCyfbli+mYI05O234C3iwvkQ8O+Z1
Xm1X/qEuhaKj2f67qkAaK1tACm5wbcv29ikESNLFxylpa1BRgL0K9IYFILIGCzN7tvGwTzyDafhL
z9ryH1tg1p4YBLO/7or4lU3/iDWl7TViPMz/qgQVxnGLGdCnHkf9JUXwvdhajexixgqdQXhy31CU
ab6HXBU7edVk+KnGartdID/a72SCH3sX6S2QBFjNjbV1nI9+BRK7v4tvXzine7o3GoPkwodINUV4
E7oHXmOmju2NO7HWMWOAO0EXi0fEueu72kQvJXrEO9LkEqdD1rLkqJd2pfPArSSyNFExN/4HEe46
fQNmw7eEo4CJ8LB8p0WEmQ7lebrbe834jRFVDoYCcTMSJKluuCpVqPpRZ6PPP0W54Y9b6HCEBHe2
TcSg60a+qxB4ezICho+GMGEJIQJ/OL04/1utiLorhMSHYxLdQ8t/EtoFtPnzpwjVfCpEfmdC50kD
0yTz0Q79o7t6HuMm1/0SOQMkE+tt8E0JmNlzc0mvEvXzjTxVnfyK65XE4DXri7L4oay9GF5mjCov
o1wkWvKC9Mv2/EaYN877FKzHfRdV8y6lVqtCUJZha2KbE/biYHJ1PWjNXZX68s+VoiMf4611qK/+
Y9SXeICMUJhAwmFlwba+V21x4LPum7mlWT4jmUWNjlG7Rh0j+m1IbMnVpdttroV/UqPZxHLEkN79
q8O4un7EjT8qqchx3u7ijKDLHvZmafI7L7oOeuDl/KuXmpKCwAPGVEpCRjNqCaGEOfX62DR2TrGI
hdcb2BR28wgfsorGD6I1TO69p7UIcofsZwhO89Z78gHDNeV0rLrTpD+05nUFUjwTbUQZ3frZUpIc
jH/+YyfbbEGoF6EK9En58OiABi6zwJGrDHXQDyY/LiZG4k2Q5awwPScavQ/IJHDcq3HXkCYfFM7F
lNTUbiL9uidcMqAOYBwXk3dhQd+GWEMDT66BauP4ATbHYp9ar3X+c2swCuw7bitmPW+DimInOOqZ
7jhvCCprJw8fHArT2Xf9zIsITUl401xWDTtX22UVayxLnitSzbir4hZicjGKbcLg0QXJlympu8OY
UtAnXyqiqvuxc72hFEf3lHsp3hqxY3ePdHqXYccYTfk0TxbXFwGmKG/z9IlZTdpd4+ZybWQDLIIL
lXSH8g3OMZ8k5UWmOaifELIKpbR3MnfwcyL0WNl6Tq4xUOqHWTJQ3xxB/sYNsA17zVaTQ5m33xZj
D3QhvkTx09QMMJdqD51hhiGpnnGa2Qejf+IFW/+fFwHinnU2CtZftn22Q465sWt8vddCTEE/taSE
8HqzBGdyIIr2PfS8Vs+kwu0b6n8pxCm8ZdOznYLa9swFF1mEdygn7tTaZRJJtTdcW1JJBqXHwx+2
50Mi6IUGT55PPC8O72actjBIrwrd/3HNf1g/YYqogmRGn3ferGqBNkV5yxGiLXCSBh6quf6e2ehn
hJT5NeNlRjL7Z+QRNf035H6UmHLVnHanevr7MryPtPDGWfAPwwuOBy8zZrG9oFpNPhprVTyA/tRg
4MPSyP3xFH+8Kpi20sIekh06KdYi1TmO8CdYk5YDrz4XwUsm9QCg1RGQUoehK6JwZK3ddCy+OLhH
x395JuSVceLJ96QWmJoOKSXCoHoLHxQt+fY77JXu12Lya9DZ9pxpOQSCoEWVQopyNneRnevEcaSb
0b2J2vIbNnwwxxXE8rHM2l2Bxna4023k2lY3pw9M2j1/JUcisEk/Rstcc4x+HHt3x4/oVWrzQUne
50D8xzwOy3HkHOKJqohLhw0n+0V5nM2szedo0OVf8BEyhXkk01oXQ0LNDNRGInDabp6LjkdeLLq/
sP+mx5n/V1zFPealSciWgCT0Gj5891Z0yiYhy24ahu+yQBl1BZ35lTAci9liP7can3IGQDpFYs1g
hkhywsnUP2uij+9DbgbJmi+hCv1LvPdoCjbmKHZx0q6MmX6LCaEKgjHU6O9mqX527ULpX7N3o4G2
T8rbAuYdWagwKriILH929dggDufNXmebqh7gbijF8Bh+XyKZX2YGyBfq8cZ0bvQtsXQPli28A+4L
l1pTsD+VtTD/9i1uvFQnHhSzXLsUdajtKxU/JcRKGFJqjoRba3NzFrKqd1Wv3xEHP2FXhxq3R2dQ
wG3itkou5LQe4oByhspWRBTyPTt3SvNkwOJHvOQvCFC5Z5VN3l4RKwPHqvLM8S5d8FTkzMtw0nAB
VfibSKAO/+tmUy5dc9WptYSRquJ6ao+g+beH8m0mmVmxkbNL+Y86QdSU15d2oySQYvxpHeKuNzgK
IwnHUwXkIWhNn4MljiZSRup/UQtCJy4h6MePBj/+tIbnHhW5pWw21P91JpA5BrO4do6HqzJz/AxR
JJMqQeqaY/1UOzFPhWMl/msm2Cr1D7Qz/HuM+iTSuAt9Dh5u5bCt9sES8G1LIvw9UrBNLd0CDNgc
wW89l3Xk4hPAq0siK/uz3bAgRV4U8EbeZn4RJefCRK89GWN3DIfzTKle1ZLijcbU1oFfK5nWkGpb
K3kkkVqUVXTEPKoHN77JGxtvVveBiaXtkc+Fto44sL57//mb63JNUDRENNaAvtEbQyPtFqHQbbop
5r8208ZqrfDNs5lnzOLQ4+TEp3K2teHSX1KK/7AhvmS/VevN1a11pEweoJiQ/epfx7XEJDyFi1G1
TIpPp3pSH42VgBw7yf4AzFW1DqBWYKOQWZfNJW3cjoYaVDxE68A/s/aDguaQFxix9N6sDQobKStQ
NHgAPnVqg8D6W3cbyNGctV/814T8Yq0ESZSVlBXNqOT2qawhN7RTNEAW2Ff5oInQXD0lu80Z7qBy
k8970iRUzb5GvKU5HVCt/j4j2lBWuaC3sR9suyYwjVRZ0VtEKGLhB5qPD3FVh9vHetzOAkKRwiUm
RGPG1Ic2YW0wnfXmKSKV815a8mp2X+8ibSTWeoKaDG64mMhouYthqOko2fTKXZteL/7Yb8BtWX+5
icE1wMQpOnSeSrJFM2AvAkxtrH4Jx2o9WZOq5pYdBNgFZeyKr4KeU8XX1G7QXCh5EQW26tExX+Am
o0VeKnWlsbWAAmISjHn8q5xb62xnDuahlTnBEsr2wCLGQfp+UhfD8Ym/QsmBHgQDRUQ3s+cvXC7E
uz4VXBiwoA5HYIvxqh76r2R7n+JFGgCHCRsDkDUIiSj1m9t3ytx3S6R69xSTD610ZBNQ5XBgIpBH
rOYaOxDvj8TrvJWk6ZmOdcu/nv5TTcYYCiokavoxO4ce5sPGlJOXH7Nbl7BxCPdsgAgBiFFyTCmY
dMq5Zly6oxT2Ub5RjFcgS+765xVHKepy9szaID0PXAx89wCl8JVp8fdv53Bz9t+RwlL9LoRIB+uz
xn2ISYxhXoDx0ZZlq/TpC6/Uze+R7kDWRB6oIs598BYJb6jiFqpiasdmVvMvivbLEvdba856G/Gq
JmcbHXqzB/ZPdrHaEiroNMrx3zNDYmPCt7JRBlc/Vli5ZVNF6iVERpv3lyG+GZ2BMOc7mh938MaE
VsneaHRPracY49CRsmp+hvrbHe+LinQIxCiOnKjOD7NG/odvTCdEOn5yMEzslAKIjNMLrbSn9mLD
riUo6Zq0VyNLwXBzSKx+HOFTBcy4NDsCZaXI8lOstbpUMzv16wY19Lr22uQpfty7xpLSGwJg+DM6
viWN+nzIuqpjCufSgRBmTTdOM4nseEzDxy7CJGnmA3N94grrSEGVma/xsBYkYjeLZm2uNoo+sh07
OTKupNf+W4o5P6FTJdtgT70lGL/SYYqUIIXZvvYBnRjq8KoJFJ9Bg93zWavy0tTYp99jqMglXpgT
3BlO/FtpeThUeuPu3qmimus73HOr9mjUaWcht5bv7nmONT6aPF2aBWEVSGYUOfw0SM+QPkotm15E
1U5yoNFJU0XS3nGFqmD0dQtdgXEvqfw8jFQbcIKXYnsMw4Q0erJpwIfvm/9seO2++xsxGGDBhqH9
SwxMKzRfjixd560fFhQRq+ESj5rlSwyd8PbtzhC0T5juplorlgwPo8oen/T9meB3PunEQ2ZcdFGy
l4sbRt0TBeUOZ70RIrwZCxryp4ykdleI4LKQTvdL6+55JxPSFuSN4qyEEx2I8nSlogr1XJWB2jUr
hOTnb0CSjZj9ZyEpdJp9djSx5N1pNNvRVD+rPK5KrNTmdut3FKatHPISVmJgo0IL6NIAARAmQtie
x0h1q2K4xLAeLPQ1CxvCmzwLLFZc+031pCqgwYmd/DcSaD5NHW2TzP3HrYEa9EVvTQqevQ5BmsvC
QCT30sZ76epdzjaOvqDAn7S0ntjHcWZNWieczqlLMasW0JKNTOtuLEPGmZGiiJV+c7G1OUzgQFfr
g/mPJ5fitOb/oJf+w2FRta9X4r+fjWanVa7tMfMruzSCxnMDAxlhz0hYRtvcE0zgKYu6961KPyXQ
rd537hbUyfhvsE+ZRo4VFALky+rX7G7Ue70wNfzAGxq7dsLXBHPfOidAeLWqjweHqteukJXCxsvz
yevHtOEKagubkFqVnITrzrLpsA4Vxs3DtAq73tCIUFuBNqHuz2OlgQNVgRcHmb1Y4WeSGw9RVhyd
jDc6MnSaRHv8O1wrelnBoDl0nhbTmsmHgpNexmr7eAfNLT0exNH3X0YcWCqtGGiK3Z3o6/UtAJ4D
gEYA8VczMG3lPw/c3tCulrxv/7GO7nONbz8JAfURxkLajh6klFTS5wwSMoh8gmmIZrN2lPo4UIOJ
D0nqMPo3JB9hrNHs3QfHbz6GeAZZVsBABR6Il8v0HRHD7LA+soKd0G8kYtRgNv7/3dBiTVwDWucT
TA2yx3EN8arzb+cfnKMZVFlEI+X+M8iFIgvj15TtxeQx+NOCKdlM8U7WQKMIcHYODlZl/4rxV+Tk
Ty0XPrBdwX5n/7nkyD4QGFFrxo6iAUMY6da9y/DiVlN1iCrIZx28hq2FP2+slafgre9zfYsUegJ1
BmGyyNhX1sGFWwzHaBG+gum+kkYAJTiB3Tv14Gm9d9kNNPwdFQ5DNwUs6l5pjVK0TgfAjegVrPse
o+CIxtHjiqRnWZfUySrfLUkACXkUZCiZJEAhwQxcnjglI32Zp+OhLyYAa6WEy/T6eqLHrheORbWN
RG4jfCX8FFsbat0qr4ogJ4bwqWCm1itTXkFiDDed4vLz4OjKqU7Pgungtn7C3MDenNc+TvdBt4Q5
CxtKKQDLiveKBpRvVZ/XYFadZJLPM6Yc0ZTprYk4ziEqrW27eUi5CGuew1Eym0b2YWEmmmbUmB3L
xMUocG6T994UHg5Ey2N/zx1+DGE477qpqtmE6sZMtpvu9l66tjNC0xawGDh+Sje/4GMg6K/CJg42
p8Vvpunug6TaNKc2Dsu+B5S+067kyRX2OdDyyZo9NPwNVm0L7dmXwXcacWSXV9zsiGPe4ok5z5VA
3zjnwWvMq7fF6uuEPpOSyn382lIwjIMzQXPmErmkzfW7wYs0cp0qmmGGR9y4yv0mKsuw+ZeCaXP7
WF96dl4VFE0tUUhVfNMWJ4A6g7NTpwTjswqCaRgywCk9FxnBsM8oN0R+00zjhj0QS4lOX//5qdoZ
NhpvvCu7VLw6STmQmYG/vXkGItPPValUEIYJn7HOMBLs8Au8CJfWpZbWAYHjF5/rA192DpiezKO9
9aqM9cy51obDKz0dOxPQ5EWHM4z73Sa9V0JuWttTFxTKX9GM+mbezQ1hNjOReR8UxgSGPKnZUR6/
2RYNHoK9VKj9JppbUSMAWBI7Vcmv+F8deqeMaGjJ5KJt1yA7nA3UAj6shxTnB5ZzTNtaPfABh0rF
F2VArC53Vm5bOSct8wOiHyoLFxzbLhVNnkd+VfSltWn0Xe2HqRJRGgYQbGlMn42MeEyXb7hhvLbo
2fJluu8j6nXhrMMGDpf0DDqTVFpD6OdzMncAw1VrpuVLzls6KhzG8cYGyLbmjLYBBHeTZN4/Z8Qo
lEEFp2IUBsFpPgfwF7woPsc7bEq+dX5R53KWzWHV71dxsz3rnuA82VPE9YEtc45nPgxB1Y/rAO4E
31lDuThtQk0NBbdhHnCcAa4ZP071Nr9ZKcGtkAwJf6cH7LURtxrYgoFbOPiwP/aI9p2htzNGYGpk
DnKkTwSit8jK8cJiYFDUDGb105yzTkC0Jv6Ia6dFdMb1ZuoNyw3zwv9nOI6ZIPZOB+1WZMvhiWhk
LxyklYYsqeZqxLiseS6ZiR+3Ev0rZhHgFMsEdvM22ivtmBJQToELGgwqCi+/sNIgYuXDlbAqPkjN
8cAS94D2ivCHiP+X+7QSdchmz44r0RtV22zBhKBpFMCpBKZb+SMIdpwRh4IPZCV9H+I9Nz7/mqgN
+G607rNST5/MH7DQS0/YXxlFUpIfo/cHVuX6+Q/dkhO7OjlBmpd5ARx2SoUCabjGfYyBQ3BIxjKo
jh7N0rC2TOTcaJSLylJs6IRA/5izoxPtRvXiZncSi5a2W/S+fVhN5KrtNlrwlS1skQSQCOgaExeq
1yEeHpp1R+fewxgyYw9xvnhiJd/B8s4FgPhKmuo9fkCtlJH8y3rFnBFBH8499X9xVvsNjYKjKYHO
GJxOy3yjSsoSv28gTuHHhRKCjePwxUs9WrdCOi6iiHmbK4jX+tFLGW4m+2SCpIWU05yKVHkwXR7J
js00U3IqxeUbKaJwEopLd3AD70hu1Dh6kcAtmF3+j7ppvsValUL+AgCbP7vQLjmvMAe9iGlmXgv8
kY4nyAeLdJBbjWMP1KO+/xjHvP1Pi1Q8uGZRgLi/gxqrA83RrOlJAzYh1B46rwi9M6ctsqDqgG1f
0mOlNHHronKridex5LM+E95fvMcXdJLyzQOaMDtCUBYzXCO7o3hoItID0b3YVyBFTkDEQjvmazRF
5Ms58MTv9aqXwK6ETOoU1HxLCLeLHJO276Lijc+vRq1g5v2wmP/bEVJHLAH9wi8i0IJ3EKSlwMS/
Ie7OnxxHLYLxnPR/d0NjF0uSA7Vyh23R49sy3I4xX0wLCS5i0gzI3Psb6fjEFPXEbABwl4j6HBIB
qFSss+OeX8rANnBtoOvho+wp37pQAC92k5DZ/eTCxp51rdqw+VAABlPQjhVzmXJk8WOrXpVqa25g
qYbY7JNllT9q/pY5hcvsOfKvkzSD8DyKzWsfqFeX1HhZLPgMHKo4CkVBWU1ggUvYF94dIS9BXpZS
6ozrnkZWPR6O8Md0o+C7eWm4Gnv0OaYDj1IhxdhYZJbxz6n0fU1yW+xec5IqgyzAwd9Cvj+JgT4q
JUImwz1+R2iE+GeDm5D1wfegi+qbvMDqBBLCWe/9QzSnyaHJU/wckwfkhg/ivZ1/iTqVQ+j6jOAQ
SBjeIP3Zu263w+hFkkt7Lre7ybEu/kF9V+76j4H0y8hLcMHtV5WMIuANTeo8f1BJOKH48/sfNpPH
dQQllP78eVMSDLNE4+xdWbZokpYLztj4NwTs31UB77Sa3VrB/4wL2OKLsn9DD9JvnkICRYx+8ys0
e7VU9NYaihMnU36ssp7VdCyyAhwQ2lPL++Hwh3l+o+ZAOZe/sf4YNPGHmTLH7Ac6GSC0BA5lpJgX
mL9WOmgxDwnRgOey0tz/slzOPKHFG6RJgbZmrFGfQO/Pw5hGoMcoAnXezIL9wmmK4JR9EVWpdU5+
tzIQL8LgnWXslk//AfjkD4hrxAzA5+3NVyxKamMHj8slcNoA0FpCWxy0hYAbIHQzHjDxMkPmFLpa
EOZjeJJ9eKjNx4SNNl8XSAJSBpYXeLwpd2oqqdUftnc6qCzzKgL6Wrm8rOgdw4jWmQb461LmJbzX
1JEQzovJRJf90douBseg5rCtEHV6h3htSEuZouPZ+UzCWfV1bqxQYbi8g5e6wbNKceFtFRFFpFkq
9xGNzaAXsjfBszKoDz2xFC2AId1LkX+wB/MvtZR1gtaIUNnaaSenzl6EfHHytOH8aOHJ16eDCElu
zn8gXBKEOnM1CUG4l7o1Zilcm7JJLPpkQhtTplpVRFKzRv7S/iKpQ76QzUUxmeCKrXWU4P5yhk5p
yuggnqguoPOwRWmsy01CnIp2OGFmB+JlXMLOKfhPfK8P1SopwZd+FzC1R3B7cIAHbUHKEhLyt/Hp
3+PhtBvRzNcQuhwN6XB/ykn1Lz33uOBJ533kqpCiz8saUgX4rfz+yFPKqlG1a6J1GbEIMwABk0W6
eSudcUHFQUWq/V13HekTeGxt3V61BSAffshDUbFEpPq+zxEIMzpkrBtmthqjEe6hLGZ9GdnF1y6T
WdlN3t1cdUmWMPEE/RFSWi7mYb8MS1RuNEDCnlO5W7Bk3Dn6PI0ldhDXt7AR8qP43JdeffT8v2VA
Gr/57w3qNEISgXYWsCuhtTgl3bqjiy8SaExX2JHXTubQ/pfTx5OIS0yCf3X539knfF/zQk9EOylc
jeJ2VlWKMVuRPa99PIMEvsfvmO9acBnUT379JgJtggDh5hutem7P9WV0q9d8wl1LoHCuEOqrIw0S
dk4bXUPt07zyKDuuqzWGTwbJs/o+oFDUFaBrY0N1FklPItpk16FD8/2L3pZpvCMwXY5XhpSI+EWQ
91CDlqF7QUgg+gYluQRjZeeD+ez9Zckk7GNlv2ImFkEoZpff8BBZcJhuHU0NsLOZwTZJNZikVAer
0fWPjfpc3cZbQhLpRYewfDMOPrp/+W9Caw9xNKLYNA6NrzJAHOjGIyG5LDJbPVzm4v4qrzBPPrla
8C83YWO9smbaFJvA6nVymUXhj8WRunvT0u3qtvydIRmCK1Hn9u6efHhU3b5g1zPOFw8Gk205SdIP
k1t2RvLfXOTcGiiVnIwOLBirjY/nEQel8HLEcNw7d80pwjwjH/BuAkSknfRTlOYX/fIIi1zPIwwb
MBx99pl0iOctX0fMXkXUODNNQdl0eGB0K0OkehGMPxE67lWJKBqFCp0dfC3TpOfZmZDImTM9o0H9
F4KfZESZ4G7whzC602wWn/9dCMr9dmFgoIkh27KVqUWstaZ3wOeVmrq5zj/yr06pxwARB4FQHCtl
oeHKTbalkvlvTPH3Fb6vaU6LBVvqhCCGq6xTKCoBbM5I2fYFusNIcb3pTz/JCiHNjH33J/8fDHJN
kreyLkqE4FEkq7Uy2RDguA/IlV7tE+9T/cRFs+HLE5OotL/yrOG8pcTEII6exKJ0U4QHqK4hzoFr
6ShHOiO0KC6JKKoyzANdDWHPK3sLgBNPuCPv7o9++KQYA3ZHMnlzKNk0/CCAFkOSa77kOCzsmNwF
Sl9vWdF6C1XWLWAflFVOJDSGA4pWudAJ6F3qqc0AKpe1QDdLNLfR+yfTWGTQNB/mDyFoLzsXRli/
U5JOoUI6OGIt0azhPLgt7Qrp4Xh4+J1yYXBCTn8ql2QYlmTuITxLb5rwmYEmCI+sH6udv8VkLOVe
gBS0+XuLIiEy6sw4i9UFZzVYPDwqMFHAd6B5/mTn2X65tm3FXFp2tsOcSoUnNq+wfQCBJKs4C+3t
ZTLBsDB/yrLbzvUC7wFml0eE82npMbjYYplvMXCGUkj8wtJcyUbn60it5RO5HKHIqAUfNwwZ8ZqC
odPNuv+7iFUqIEdwl9gEEuvkLAds8PE8g/tSzov5KzEJkdtMNki2KDssEewgjv7Hagpcl9aU/B97
e1UkB4Y/zHGp/fUR911folzGVWf22Xt4rZ+GCGrrJxPNXejga0gHf6Hy5RBu8nU+ZOSO1+g+NGNR
JZVCCN5X8Bv4W9lecLkWqSLKs096DTrcNaVPlT7lWdThyihobXdr0xe6jLR48h4w0cKyDO0rBq4K
u/Bqebq7mTZqlQ9KPG5wd6/sYBggnsD2hw0HCVVCn7qpAjA2kFO15APN+GCgy1aIM7HePXASKZTC
+ao7zNAhuT1I5EtJkBHsHl+FCuNK+i8ohpjOIesQCf3rzeBtIMyelkPQW1C5e+/J889SPgTaCsKy
QMnqHjqb9mFLjgsDX5FZz2WynNDOUlta9buIoqsKG/t/OZ+6XXTV3yav59/BWT83Pqq9oiDy2Ipf
2TYL4CikwQ/2Z4IofIDNHLSmPg0B5Pqywx5E0NITKXSqBA5J1gRiPovpWbAq5y/4NS+oMwUAr+VT
QMLD2oKtDNjL/YUQxzS6CHnVetqk5+61j/rxzQfMtbZlF3j40xYXE9DKYqWB1PS3MsYWiaWRm1tB
Z6H/R7KsMakPu+uXI5emVIYAt1s5GlZvuL43SPka8qZ8HM8Sja781UNmw6pLWSAJLKhKdPh8CaQX
NPI9BcUgc5W6blaSxVFkLv8T74QKMJQ8gRKmIpmCLaswHV9dS92jyxBER/KNQhx5oiNnB6pHT/yh
t/auwiNkOTrDqa8PbzMNl0B9fk3obRCBaEBCx7dGWZOcgmHoylBst3gVYjwZQqOPTxn+79QJy2FO
9mMfadLwxcFYblE0Kd4GHcatKU5XlA3Hf9baNu+CXDIKVDAXWfu13PrLLKGWoSq0LOtdp1PB7RYq
OzxVp0JXYySr2ypMCZZ+CYpyIrTaP5Z2dDZXQeacF21BoMhr7u/tR0BqW+rJUnIv6R65IgMRl4Rl
+xSoaf/Da322AQ37B+YFu6yjua0nfYm8kL3rn7KQzjCRkAdivMQ5cAIHhzkoJZX4DSr0G97Qnu6Z
Zgy+5mQ9OyQZ7J37xySBUL24zUX33itObsWFc8ge41FJa26tkN73azT044+f+35EPkB4tobjZi1q
TgdqJ/jAyCiYRWgjz+2SEekAPyarEWdZ8SjRaOwTNsiy1lcORtcqAFxuT4H6tt6qzfiZ9MCFVdjh
ohRRIsv1iOYL4GdLOxcYwFS7vqi1lDWDgzu6K1e6raQ3Gsi1xVffLXhsVID1yzRf/CCShMSPbkwo
RgITiLbBHXfcUqUnyDh9S2jRUKoWrTAeQ627t9vCn7hWAieO/XWie9QIiTqY2x8JTYhn2YCLtCFY
8wrthXnFU6hr7qU/Vu7CapI8RZJHKiz2V18EF2esdAHNELAKHXgcJwSgFrIB0J+pE0pWmrcq4+HX
8CFgubc4B6Ar+uFkR8C5rHraXWeykkVRyohnsRROFL1gtcCPjeN8gkWFcOfJdi5iPnCqOI5HwAYt
mNFotFPKderNC55rx2hQTlgwuYSiMkv5Fd3q19WnynX5O1jGKs5W9QR/voImifuDz5U/eUccd5TK
etMpKGw+IYQGwzDKQCPNKk8b7ZL9WMdLflbMolBkVu7GFxaqZkIdLltgKf7QDpzjlMnSw5Ph+sZg
eXmm4vfjx1Z7JVM6TmWTVaSW6NFMOoEt80geDWm/Jiqk7MTuz2wpmHenlQe2cZWp1S6oAH+nn67V
4kwLknWOw+ijg2nmOM/onJLfbBLMeRR2Fns9SLbg40BLux/HdCT1VvuUqE+i/WEQPtf7KU8Yimde
5fZoEqG/Lg4US3ExbCeGdgPBGqIc6hYm1Z+vLIAkEWW7pHBsiCPfmJBTNQx+pCHdlQ4RGHnX1i6W
W6sCwEiIJhGqfqQB3RHYjsnnsrX6SJcqCr7adnWsPwGqsfcgfNWApJ6rllXWLhlAZFXHdHADAxgR
HS54MwUpX2UI2Oh4kQpVEuMfOYJ1Fc7xDSmjhPedJoBb10DeDS/itiK9u9Qs11IekNbdt8MM03xD
qqhNKmX/ae1u4r476E7xeZ76epq/jVaf3KGUQIogUGQ6rTG7RW3vxT50yxu7yktMskq8fuJyK7O3
qBdk8o2QAPmF3sgBQqXOKh3/z6P5zDMcs0G3JOfRTblV61p1XIZuB5SqRCwcIUMIf/lawbxvmLaz
ciqhNu8gzR4Tpt0k8xOv6wgLy+SXSBSqcDW9CjyIb8NO9lqxXER9RWedgt6DWZjpUxHBSDshWqUn
roCmCTaOuR9Tz/Ggk0db2g1HDvUm0qCjWYBhDcEe7K59A4/NxUswqPIiRcg1E/kzDsmbMJnzbvUs
MoZbJoVamqsKGC2ouFwnCL5/hiYVkTeL39ds5yRdyZR4idBOOXM8+FG9EyfXt40OUbUP6NRZb0tL
viOxJ7XdQs3IBks1rRbRqP0o6tu//eNjU6HSbz/Zn/kX78hdw2u1BRdwuMvWZh8Asd2h5tN2uj78
nXLWs+GtHATevAC8UsaXS1Jz5IljgJYRJXIigLlArZ0vuxohv9vWafuPsYMR86O4uX2EmSIoyrli
IPHoyHve0hOKMf0Sf+TBMNmY4YJ4F4YCltjdkttvRo4m5Cvw/mVB+TAbH3aJGL+DSRo3KylRs+qH
hLB59wZ3fqOePwjgcJnEuZFnSwZ0WTL5eK+4bpID2h3V/XsXODeZFD3/2TlonKGjlsFXTmHK/avT
x8mb2twJHtENyLy5uS7ydIEBbsL5palmtpYYcF6hxxt8xKlQhpvskNfesI7duP2poGc5IEed7S5o
AdfCFpmnEtgGneT3LMx5FB9T8L35A4z43MYg+AMlEGOgbroUn6szqJRxUaX3zJ39wm17hMEwCGjt
bM+7hAKXFmxxIzta4LRzA3HzIL1CEpsfT0shgbHbr91e0Gm4DWn6ZXGYqMVd+Zg1cGT3pVVdoPJ+
Rf2+NsLu64HiklY0TTAI0SXxQjuoQoRS5AWg4EyM1hMgEjI065z1THcWxaP2Ctqwp4z8Aj0yz/KT
1TZIxjqtSRxIhOl8cCZtDIp+aspoQwq0fyJOE6Zki6xg+GdpMvyMSm/fr2pOL+1VcRBrcvLm+q7A
vSGy6IUglQN+psuJgQFxGY9OoKbqDVGOk/rdNGQ87IXOhGB/4TiuByPDEqsWYUsRLRW/159w0rGk
DVTU+h4AvySzbOJWSGJs6gQsfbX/I/EXcdl2EhLHfCZ08Q0GC409FjDLR5HyEl6CCiWege5d3IKA
u4yVlLv1+L/bFEz0dH1iHfH5MddalUnDRK9A7wlpWeDVgrOuY6r7bGV6+RthDtpM4AjpDAmAEgnc
u21Z0dMmzPZ03vOISJeKicvRuklEdvVCvyUo/IHq6yyNUOGa/6Al81yQC4xt55RQmJwHURNsKfQu
isTC1sU5lOKTXWGP8SihrJzINU4hehi22G7aXeiBHQ5NAG+9z8r01SGtjv+PnFhx9ZDF5Lh4k32c
t/n9EU6yZy2UPdxhfpT2+EqrQ+gWM9ymFU+EBUwjDnkinK84FLOKNCEPDEqRvn9L5/+YbGYvp1rl
qkdeVH6oO3d8zYFphX4744x9zfBtB/AA9nU3pOMbIbiTmXMGCQU2L8N5MJ29YlQN3DESF++G1UBh
d2nKGkFmAHZDWzEDMV9sdD0dtZNe7fuEfMUfDxlS3sKrTN3G4oSRSgYcUSk9qbPUwOND70+1UbOA
3KzKNZ24mtoAFdzd56BCYOFjiitDOBEWCULR9fJUF69wjw4BpP+sYa43gGLTGwBWet6z2DGo2AMs
SOR8qkPsiQGHQ+fk3Tmn4SOwE+UKnnWVWnEv7W2UzIQmf2k5j8SuaKsH6RkWjmKe9hnwn99VOrgF
eD34c7z7f/9R0tCjHyllPFcXuMtd3k3/PT07Qoim36kaL1vt08oE31K0qHAD+87N3FHrcOMCFyoa
v34n8Y/FzlLh0syLm0hQIncwXak9lWWoH7vR3Uu/Ho5SIW/sgfJgKh9hAvbaIVm90QuJU/+bRDG1
BMkYQuMwIQD33QJaUhNoKFYadi674H/Y1DoVNzJwZ2Dep8B5KkCfjk6KS1Gk6e5+PZ8g0LaZD199
NW6R4IFcea0ek13jBUQFY3toGC/4EwU2iONbwRhlEzT4e9RMZoJgT5x8FvtT+aT2yEeSri+i1o5n
V7vo3SoKY88Q8P+k2ToBzhsNK71vrlZpQKIEadaPEdCEjarONXdDNSUfe/I4inlueaPRBLxyrgUx
VHVTgx8Tb4HTcMBMDaAt7+edt85Em0m7jRUrlQwIFFAna1iZSxBi/U6MdesoAL7dPjR7pn+VTa/N
Ej+9x7LKzUVnTeTYqlXR7hAVrKSz9hRKm/rjP8ZJmDMaN9W0hMKtwZKo9GkQycjdyjgYORzXB+if
SUVjoHU62YVkq1v1Sq8rzt7i2aUvgO7Ya/c8O3qyPt8WlogzHxLj3ZgJg1N+AuYS3LR3Go14TfOE
cWRf6kTE4RP3BH7TP9Ag1yg9yRrXm9QjaN7Qr2jZdtYF8YlX5niEvG6lui97p41up9Vg1RRB9zJm
x/qVfFgitrExy1dnMtCCXhdVAmeU9fbigd/g29NZ0YrHUFF8y0SDpTHopAUqSJ6CZRUqeTaV70RW
icq5BtTXPU2VWr5AloSWkXCi4YKJkQzoHzi0lvqMP3ZpGrZ78+a7rY3RRv3zhlBFOHb0rCE3kTti
u9hCZuXtuTDd2izs/QO/oSe1dibz6unT8JYMTZ5UMV0LkUEVXAkc396eADafIlj1HInV1NYAYTzz
NjtrFn6QN5UncKCewt6mglVSO7N8+f/30VX57Sv+808ucEsoyOeKGaNmbPCcmTO46iTDEMXveTHG
+m1eOu5yTWnn3pHgHBjrAaQ4YB1CVJ8eq2Ur1Z4ZVtt0GnR7FAmAHKC2+tWOpgDajylqe3X9c5Rn
altsTCdlUT0teLvZN6/zXmGk8bmmu0CjLXHxoUjupd44CrvThJKAs1+VAds8F1sJBLxg/O8fN4Kv
H+To91dFbAcCOpn0v07UpAQiFmcN9g2y8a9kZ0oGHBu+G3wmC67F+8JaYwgYBo1mcof0rmCQ2rx+
sk5r/w+cOpvKJwFQe1u+u462lVDrg5Xd79ddo9ebVZ7dbak/zfmR+kb0H2tSRaQ+MCIwDoxf7utN
cNfdTH/HQgwAB7QBPadpe3+KMzkKypzfhddcK7MJ7zDi6GWxQdyetTHqtQu5zx8pd3+XnGoW4fG1
dKxgRZMOoM4P2ExAFV9RUj69Imk4bwD15mmzcjuwbs180FqILAoed5ZopRZ5iVipVEQvDE4ic0Tq
2hitinMaNizO8nht/pl5wlaEkRVwWj0veYa0Moxx+1xcstqYfj6xTtQPuNj2sXwK4PzPsrOmVqaa
b0yD7R62+QZZ9rgz5eE4x2e8q3z3j4kLiHbimjZSvcxaMVeKQE6Muqy6GehO47O06gL+LSbUVq7q
Ko7X8oqjIva/Ov0m5k4sJVuh1HERGnEcbiq5bO20965uMKyr7Z34fvLrdpvPJXX/6FTkzo+Dpy6F
yt/0DnxD1C8mZYM1+WUzYvsKytFgaNfAVm7iBuvqjMudbpEPvyihX1jgSaHenL4m4JkEPeJeuRdW
GDMBlgM5q6xeywvjnNzjmceQGav14cT4Afl1MdX2wq3/uQtdKkJCxlB582et3IDsQkKs9T6zUNmE
szV9cFNLsca1uy798Tw4PeK9FeNOFXGQOZIvGb+ZEudxNFI++O3BSs+015Xbf4N5IYl8hPqxi/MT
8wEXglkoLrDGQOIoEQ3T75IFK72/HadNjeYL0NGNlj/Lh0Y5BMB95WKBNi4GbIg2/z6G6L+0oufR
FLXutr3ya8maX9igrA5CilPOhnSnH2gHAmhye/uZCpbXix5m4NO8zNad8MnXMLGRebfLTJLp9OrV
9joXwiPzI5Fmp0cJXZqwn72z9HQ9wUDFysUVT+O76S0tOZX3gxs5cNSbOjcf3xUwOdBGz5BFa5Ym
i9zgRQg6WYdXqEB9ytOjjo0c+AykOTn5+ANJwFtlsNjGJZEdnLN5bnPk+aMZ/Ye1XQzufNgbOvZP
gFeBUVx/cFHCxOJR9JK65+MYWcP8fDPxvVJCqc2u0tVt6PbHAna+iBSp/ZmwEfSzJkszEmD3tAua
gUx4JWhxxLCB/1Zr4mhPfjE0n7F/SYpXcbSuETCag2M76Q7/bc/axxXT2r42bVDXLc5JMXOW425G
QTTB7lihjad5VEQcEUHN9zxl1Z+mFjM5U0uviUddwX1q1nqsNR1bAWAis9Qe/dFOs9/cbckEGCrw
07z468zOyi2AuF/ueH8ggTEKdNC9Y6T00DHanaCLOQ+7hxWrPZr0QWKYzaX/pfsZ6dWF2/TTkzL4
2YhIXDa22EYrGhBuw79z8koaqhsI5Q8nz98ffonkev9scGXgb/RrmgU1I9AuY+XgtLkk21FowT4R
h7mJZP0tNWpTmzgbxwTKwPT9wFEasngf0me5yTsGXxVCPBUmP24MtdiaM7mUi/reYVvPvQ26Jpxe
YBqFEI/oYLT7nTO95q2S0na4L+QqSj5SdSWLF+7MZIokLIqNs7gs9HpGfI5jJK3W2VXZky5Rixa8
Z66oYn5GiSjsLP/i4qxJpqFqKYDCKQ/4pobXu8bAjg0T845hnoaIBYc7KsfYnPF5mX4DSLNr2Atm
BjkieMb/AVD3QyYIEXjWiwK1tXEeX6yy5kL+t6IX6jRPVyeeLNBWRg1abFTtDRYHoNHJwBTnZCAs
uIlbcuL0aeLtjt4XZ+NeVU/9atKbueSis7uc1JOx7OO58Rk+PUEgysP0jl3wfXRWLivqjObcsGmb
NwfjNU7+UnbpXMDZICT0rMVppJBR/6CuLwvgVnilLYJ/XYlUBPDz2JzSyg8GQzZDPJ+pLjz0Xl31
EmPKfLb9J1GneeptPz1PXVs92s17Ocjj0Q/0qgBJ3lzKJDZGuaDGPsl2/oRjVJ0dkyBgpk8zmYT/
BHs0wYb3EWuoBO7ySEPRlOYjg8CNv/kcsFhzy7VV+X/8EELChdzoAO50RydGT7veKVzaXq8gZrIO
nFcv8ZhrO40NuY8WGKKkosDp5tTAU6+/56pNNDr4TmpUCLGDHIRJBgbjxWC4eKCczQpqrn8ggPyb
QiINEh54KOucsCnYZZvKL2dk5X5RHOKJFaelRpYSvtme4qRmu2iHBfdbzzdGP6vos+IT+qLrLKIJ
wVzlp5ZNGN4O6pmzMkIKMfA5cKjZQ06JnyU/LWJxNAq/SnQInXKIrjFKK9F9y6l1/QCDOrKWNq0p
K+oQ1XBwt3y1aq3rix++cw1JvLA5dt5+vRp3wa8XyOtcFWRnGi+EB3mgojp0UioZLOO6X+R5Wp8n
uRmarNHERN2RCkWYDBjfEyTdzL6HQRrHT4VXazWNWTrlDFXS1tGw/bElOUSehSxfXyL7qYRz5JYp
RabZLKsp4l2czAg7iaN60BiiwzRggVCUJVmdCyukFLdfvciGe8BAwoIQKs66QGDU4ENE4RaQTCX+
ZYfFgOAx9jVidxEtLEJI3MR+ruOMGl9zIzBA2xTj/wQ4TkZ1u6yug9Fcs8vTLdE/UPNkBMUHT2ZB
ac+tYLOWD8RvW+LDdcVzhMlfYmpDn13RYO8RarokD7zNwHypMbvpzOrmCojPkf7GS0lZh561OFGU
Xr5U9DcjEi9uUKF1SAh6HQA7Qub1qyVffi30v7MDzMwfU+OaL9eU/zTjvuYMonc1hxyCONvUKtI0
M+n9KERPfgja8kea7yVKDhbi175rVaJhBeDjWVp+yxS84hVsy6hl8hm0YOq1t/BMg3QT/BrjaFn/
+PFc53bu2bUIQcPlMd5VSER4xSb9B3bLxCfPSQuOxcULBrzniKuXEGTIecT8IeSIyKQ8SMHQhxQa
8LkGI9YVTr3jThnCAWobitCftoGMNrYPWYQFyVHwR7PbEbIPBDGd7VVQo5St3k5MU4CgHfo7xgpz
59NsZSyI6zDIiOqDOyHkEgBdxqs4sp5DQbR3nYes/j4hV+xyM2lWneB/qTCW5ocq6j03so8/PLVZ
aTEl7WFxEF8OJAPrfluI1KzInQuPHHdlGShtZMCJz5mZUpUEAQvVu3jABAdfxHJ1ki/6i9KOpfSK
0LWjzbJQHPT3CrkNb4ucZYGam3+SusWo+vZPghA32rI12wxJ1ms2OwOA5a9lc1cJ3SFvCC90O3zP
yfi04NIw1X3ERQUpyj75pgnDZ89OjfvMwOveTxFdhXqjKmvnCQk6oCyu/lbmgLpcJHQdXW3EhUVs
M/WNEC8GMQE5V+8RpCJW9Nq2Xd+mVuH0CaYkUbYULHPXaynuw52d7cdr+vqFcoq4z5jMFqqbkVko
FWum+tMAtWAAhTQDOlQUgJcY82Py4vrZQptcXNrOH89Tad9YIvH0w64nMkxrWv2ILZHpOvlqHMrr
S43QgfkWs9Y1jy5NUNg2CY+jhUE+JSsHALl2C7BcekP9OzVZnq5wqunfGvoZoGTmXunf1STlD/8M
nOKV5afpQLsFfYCxVPnaMjI+34q0zMp39Squ7RkdRjAnAaegCVPfl3f/AAPolx2kuR89hbPaO6BL
Phou2TPIxjVNKrgMBL2iM8rTXMe0mOjJzGa+qgJwP1ryyUe9sTNYUaCGD+8B8KPslcR2BqW2sVLA
1NCijfmIUbTPtrGzN+Qsyr4IhWJyL7mJILCTKUjisY3YVe8TYpRwh9qSWYDbh8XM8oAQil6WUI/6
yVnRlLfZid91YpmATXLDEEH2vBJicRkjfzHvVvmqBlPxT7y8P29hz2aUkarsYjytoC+eAJ/0fWod
7I/MiTPWl40U9ICRWWGwRITCZAIWy+6hEJLAX3aBCQi4HM8wwhGtqAD2AzATaAXHXP9vVJkA5GCH
v/Gg/xYJ65dfc1AHdEOgBB0oePDDfm6RSdJlwuGCWU+jEfKFAkvTZEyUywrOCj+AKw2kfGXHm51L
Zys0OqWX06o4MTeJHlCptsIGQ8/9JyfVFIwBUKJm/bxxHJn6LaABHLfpumlLjU5yzobV4x7ekyKy
0qOEeiqg4iC+bH5tK8NFJJBwXMhnA6CBjfhM9fWV3+yqFtrD8IiZcQOIIqE7avjFqs7DofQ8xtxN
vrd1kHRCLwrJz7qxAdX1AXqfEJJ10PJApX5GuSaHfFZ2H2z1sxOS+vNQccem4X+J/zYCrAgsqp3h
o5/M7/uPevvE0UNlNF9c9668m/eCRfWSaAddj6RpznoAlM5RJwYUkYa6sWD+8mB7uLZdv37o0fuP
Tqd97Vft0OGX1FlAuNrcxvgywGsm2rz9QuuLcyttkU0I2uPYB0lalOZK5ZyG5vt4OUiJRuLJTGKT
QwouadgakH5P5MknC4EBrjTRoIDWTxb9INWTm5PjqAjmuB6VBRN/6O49EwDUUxmAyQeQycOAlXyx
bvtA8ZifDQeqHwM5QNaVKc68zI5yRG1rvtLiqXj1R23ItPrPYhQ/kS4BGJeXd2SURms+GXwEAbSp
86JWmUGqcOU0vJMSCdgQe0fTqQvSWQXJDySDDec2ZuXLpG8UZblngokNqgyps/YSiF1qh9IZEwFx
BtLPGcjLdWYPfuQ79w209p6Xn2fnaTk0bPQyDktpxNfRTQrW4/VPKwyVb6AJtK/KzjyF/w/PvIic
99LrrsW6yB1bY4K6l6s9GuJS47JXtlloYa63wfIys/IUUzfne88wBXrK76eVpldh1ymTIh7Pezg7
K4m7mXz+uE874V/X/XHRDhJwbCIqMrI+gqzhvP7FTF7dF0/7++c96vGK3KDFZ8+XMnYphFqgud4n
H0OWubqiHO2T9C76hg+20RoHzbsa/QP4nRKGHkF7p92vUL2+Q1HInjYd+uIOZv7T3ZwH+n1oB2u8
97WkVjaRK+hFyOQY6lNsLJU6J9+JFsZO2Fno7vfXAcCy/ME/psYXLvtozNP9V3WGIV6EX46XUuHS
07PfMMwJk2bktlUba0COPqMpkl9JceJ+EZISovbn2g3D4oE9tRpx7P1wYfLfJ61tiwCzUsrRWc1b
+5Vn2XTo9jDZpW51QzMPnwmTeMWHhdrZkrUTaRlT0keejpbr4Oxx5ig4iIBkGT8EC04D8UCl4Rlj
lTUmWKjsSrNGj94QQOjW5RrPcWf88ZSeE+EaLT8sa5SWc/AmPdMVoPFgEbN/NlLxYtPjn1G3pKk+
61M5Lgl6tUQpRvg9cXAxv3HIDQRC6o8klvwGvtfdNILATFhm0gbmppkE/n4cZcN1fhJgK056yXBk
OoM7C9Z/mIN5JMEhHtmvcXDpoZxf8CuZBIV84llbl1pmqts4O3+6JHdIgCQiy9MWOBk0b/WDditH
RoEaQxIS/Opwktf/JLlTa40u9a6JDoH8XKg9e3NWSchkz8GqlIT7moqON1SEEvC3vpzsrH3jTQP1
9Rqb/vtCo0Sl1gnI9kBdKyRcSZbuFfGP4TZdeWyosXbtIxrFw/cqo5/gz9mgooHuSY+wbDAEDHRW
RNwHBkQ5/KOwpBgdSmHJimTRXEODGRa6xxBdQUZ34UzWuKVxp1z5dbYofhabQMOZ6LVHbdR+2Ksh
GrnxXmAahWwDqg9NwjgmZrv+IXRFIC5PO6DEiT8hfmpquUfBuH+rVS65UqirWtHHxLI7tIjD7XRX
xtTYPFPWVz1e3fQLz83FSRvchDM8g5dEIikQNTsy8/uLQfeBhG69HuzSsjDmc2PWkZWAp2MRKdGr
4ZcVo4ijl9HmUwAEx914fSksZXMgVzhyth1OIJ5LmaZ6ifR04NZJBJGRZCQVqHHJOwY2De8o0ZN1
mIg9JOuQy7+3sPXQVTRRgZNORo4B0SPhIstAMvwGB0auGkyVVEkv6hBmLNJegvKjHKlC8iS8OizV
RaRS+lgCdeVJl808KawmqHbH0e/xjQvbDr4k3/L2pLY5L9aM9SFfWKjKh1HSDbjfRw9lYleUutDt
NCxQfDl+NT08tf8QNKzw1Ekzp0fOC4mBasO0LnZ3Ul9K4GGd+TDfPsz6+BoDSWfovHY5EwUmYso/
tUy2dbpNGztwwfqucG8ThWOAM+CvtkLNL+x+jIwdMAATcpJnVGtf+CEWYxZAB/3JUM78e0FSkec7
YRu85yQo+s7Txz0lQByER0m1vHgfgl8AIEuU33NiUKKoMRrnqRDSN7y32emnZjtzr+lZMZFsoqeW
BmCNMim16tXf0/mxaqmQ9veTEfMHsXCRcMhxG+E2QXgdfaHgPyGEJqvg2qXo7KQPM3dizSsVYPkV
wRQ7WHnB8tdvqWB9vqV/rRivkK86EM/WZwOlF1bu2KLrZcZQZldEj5QnuN6thIpWdTnxYZqW0C2a
UCixZuhRHxCGQ1ywLADq4mwCaNoFG/VZvWeLAb6tXWPY2EJ/c36CKNeXcPoyxa1hcrjVIH5EZVau
TrdnnrkpmhIaoE/TW0/yZ6ihg1+YAaZ4ph7SMBRxcY8gVIx/WUq987CKh4wcFyB37FFmuYgjo3hC
wQGcj8yVUnJOIuVArLStPuOnViE4+pXPiazs7rKjHa+vA5eJpAL4mFqulV9zmRJCMR4E56DWPRq8
S/grxrumSziE+uEv0coh30WCKMctr7Tut9e6wY7ApOQWnnSen94oTzeG0QDv/NpVDur5qfUBmJf3
t+00A0y92vDIUydw66H1lJiJ3icbXnqBVFfCby1OdOBNcjV3oEc0c5OsIzD0e+YeEb0qrMhJjqNY
4lpu1ZMwJKav9IlIPfGgw0lfPCjCyMA626hFIQUuJhYFuNAAchdDqFXdeSZS04cMZqkFxrizhcji
XVdbt4rjBr3oMHO7w8UvU6LvadkH6MWknN896TFtudsBUoXkk4EneTO+mKwgIcscRWP+ElBF7McD
KiV05AMty7Xraww0qQhi81p95PVwdlNnRfZpXWYoV7DvNbfsLnnCxLFiNz8VcO5FzQEFJfaop69s
kxqP0+YTpnOqgtLsDEXkJTIs2IEjgVwRtKXHXme/Pg+L9UFrmTik5r183ROptBDc2yL01zJEt0G7
RbnJiNkOXPT+FoMejug0jhPhCpzLvrTsGkWQggAoOOERlsLSfBe494nMYSpY8z1JUqUHB/cDTJ48
TjORQpptpCCuU1VQinDhN/qutznvL6Uq1r0bGp19eL+qM06qD6ftHnZuPliHs0rt47YdyD9kvh6l
a3+jSqQ8XiUDS8NDeyODFsjJiDjF3cUOjf8PUwuk71IiFQHp3J5KlVNx1feOf0XUOk79CX0/W0Ip
+feUVFTL+8iIZr9nlqndNrK1QJZ6/lFfirGnwYKu73fO8tu2JKNrKk9apM6QKJ7uNvBpOlLKLiiH
59jBSLwkcEU9+kBfcgY2jlOqwpaIjmAne511B4BuOys3B3HWRF0B3l3ucPKQk3hZCuugTRKbIvp+
AENoiyvcwgx8ixtRW3F/agzs6AhcsSwoHEVEryTTvtfXyT9dHOd266xXbZgW8lHIMc4H2zrdEabf
dIstkNhpT4Z1ONB3ejQMQ7rICd8U0p/rjaBrB7Yl2ubwl7HfRyCs3tw0CMuEt3h0rv3nYqdKg2dC
+19Xgs7T3VUeRb3T/hy00ngHMbk7263htPhrxv2OCY4SOT/m9AX4W/9OLhOpREqt7M6eCou7XThy
0PnP1mGgFIgZPChtsIT8T5oO5kH0KOXHQTxGMF/uZbhl6g0RBDgnkx7DoTG+bZaidSFpgnmhhduw
2RYY7Wdh74pyieLt6QpdC4qBvOo5xq59G98PjmKZDiCdyJN1pg+q9+NHMWIJyzIhPXXMHinnEJ7G
zU9+ls7XLQlHMs8jCN9LQxT2S/XrstK3Y0b82FnWVSeubIXf/Ol84+neQd7eRpPC0xZ3PAfLCAri
tQq/buEq4im2nOq6mMsk3G/D4Bcz8kR0el5rp3eIKr5owCZqKlqG51AZW1QeuRzh4Cu7BpYkCcMu
mGYWsqL1shvZB9G+axVcWvO5kgl4gufvA9u+3DCz1lMTYtb0Q0xOqNG0ooIPcb81+LHcNygjFcL5
S8n1qxoKOFsuBl/vO1gUQay7r774vTxuc1B9oV4B9zNdCqPhm1psjh8qSxpArENeOWLEzj6P+hCc
W4UctG8mCGwZR80+H+M5RHC4gGWCbIy9qzCjuvERDBGhaK62xLvZrS7qM8wiYAAepr8oX75Wyozw
m4u26VES24XxDbyTNOuIElpyPYtgZ9MxLdZ2ToZcCqIWyguhnXx1b8jYC3ojtuDnoRWtmDf7KjC6
U56Fx0UmDwxXNLcU7il+pSUE3ye5awHZsi2ZIQ4daOy8Ljr9MEQG2cack1Jw6x111H6zHtIR22UN
cKz+Lm9AtFCOSmfkUQx0/noZVgZ3/uHGhZ8MQ0i4BjE42SpEPJQ99tNQlEi4/bfHIYYDIgZRI/FF
lWEaHKaenh5g6VZaDL5qh47b03et1w1Y7xWP9gryt6yD+UFunfQY8MAHsaYGxJJuE7AZhq1DcDWK
KCg3cMF1IpjaJ0C6SRyJNdGBM6a/bJYtE17333AAdXGOR+3UWcSqgPFBf78tvQXX6ZhRPRR+NXq9
qNjXJc1piFyIv/F4b8+J5k/G7TpSLtGjyAD2wgR0Vt5+mK6pKsaMoI4nu08vV6DaWOJykrdnmOYH
jWsvEMzkVIGe1rOCYwWuLjUPQ+I/iHXi5/H8BppeYRwbxRDu/OLdFgIG3vertmBvoP/OLcmq8GGW
boqpKFZTlXT14DGRsXaprhCASZ29AfRdSW4+SnG687oNDY0HN6UwpNgeAo1tdWkZSOzGuI4lszq5
9jPqbsiVv2v5j0lmheiuybpcIaFsnmhefHXmgkN38oH3rAEDtyTXUd5LHToQlMOJq15/iGCHE1cG
VkigcMuUc82gkgRKf6425YsLxlP6vho9jFK1gOrXN5+aLW00pKSfsN3Tllhe2q9kqSCRy36F+wBM
/9Q2oNRe66oHLttAQAE28i5MCksHL9hjq2POMwNbnphupADg+tG9dbhHMlXdMTzj/ljBFbyzgpzJ
+Hl1E6GPtIENMdrRLHwhYKsKT+ySjOsRAtdyNG1sXUQYqW6gAdKaddGMVPpFHnEiSSdiPWT7Ko8t
IzmmQ7t1PJ8jwDRPT+kZuegadqef7wyO2DrS/QGLz9jHs0rcNe8L+Dk53u3lUjSuOGU0sFFDPIwI
NukiiWdajIJK1SCj2Ss+WgPo4VIh/vjOaNJi9EmXrVgNidrH5Q1SqxK36Mx9CXHmPV0n05A8bXgJ
tvgVfCnvc4rM1hoJB6+ZCkWzKujNoWHVYbwN48rk2v/tP1RHvGaJYlSz4GYkQjBuob1t3r3nu6qR
bd/Yu/LPeW7wsCy6iiKOIPsKbUnVAPXKiv8zWmTKPipPnNkd+3Pa6vsyfEnQhvwQCNbsd54lZT7d
5wsem39cJ115L5IY40QY89sQw68QQ4oA2saf4cd8fYhaRNQLCuiuDCyEmhHonN/cHZUK8qumZSZ5
+RBK2Vc4OAOta6ZXrLHQ29l+ptkmUDoiBUIT2ZyiJsz4DvfpeeFt2pP52nrHwUhahdN/BPOpUTI2
ZQphNvHqI3MoGb6sPIBNHPdJokHohmLdfmL7DbNdAIb8Eqd0EVsoDeRVQ4vAQBe9dOk24rUIXITA
nvKiNf3TcxuZz3d9jGmbcIzfBvx6ukMjMB5fVfRzepFuUX25vI0tXF90ml9plkZLGnAHuq8+FHfv
THZXT86bcnswRYifrHwNPOAHW3iXAubZPOnrEIQbb4aUzTvPxncIOACB8ct1D6JT72rB7e8cg4rD
5QDRg/bfxwz5l3UP/DcHpPdJtZjmj6XhV6q5AkyvnC1v9po/o9s0zedyguD8pJPCZnj7XD7zA8p7
Z5iO5BkFuZvkx8Bj4lcc8NU777V/Pxy6upbpxAflezZ1M+NCwQ+6Mej6cY062/TgkzmHs7HBLU4v
Bp0XMswiXbuOpGKamdIS9nnCm2U3j8Q9nITOBfHvJ/5+qmk+hnlsfcBQE+gGDZ2NCBuFgVwe1v4y
4DVHtYyDrgdRQp0E+u9UvfRxC80wGcCOFkoJxlFNdPfboeo6R0AvSomsVMPuj7C3L36bY0tDpX5D
tImFehEunMF94yr9WkTu3y8P6x+DIl4ktMbQADyvLPT3Kwxn3DTJm+43yPzPJVjJfqcGw67cyz6s
3fJIqesKo014FoLADw2DtY76WyrXjP7yRKFR73/+/w0rfLISMDq9BfSF3I2ALJ4OZslizZfgXQBl
mnPlMRml97zJGkbyYg/KEwJyo2IOsEglKtcWejDWbrUdR0gxtW8QBUluDrM14ZKe3vT94Fcub9bh
H/7Xk4XtjIeNEbZva7ApDcQMsfyQ1Nkl9rlUON4+g4omPpiwLOjEX29ar0vVu8cLi/X9BhfoFT0b
4wGGtl3lbpAQOUD3aJJKXs7IYQ94RL3zhaIvPgAvcBCT+zhnxKnvkecsqIkkPQ/gYiBD18Y84VUK
Ld3ArWEK5MqBoXNU5GD/72r1bZXkw5iFvq923Ss/+PigvcxcF8KSZIZZzOVDnkPLGLvbxdoT3Uz2
5foNMOJ4sVljRBP0p4GzSqSr0pafr8sQ6r8RbAWLsu4TDurnkHNFjJqCtXES1XKAoQ6ZrHzxxdVV
4YZT8JnLDJPO5fZY+d2JM9dECafOl18RV0OS5rOvP300YkgPw9HDvXwoFORY5t54hG7rKjMRNIJO
+ZGyDaLZG7Va97j6bTW9ypL9ddT4UJsTac2r1wpeizBlL/3EhsUo/PuHIc0W+d7f9FVeuQfcCTTa
hLCT20Z8uVsPP5KLF0n+f1SIt3sytEs2w4ZUa2hseAt9DVT0SZx5fxqCckd1Hjn9Sim65AZehM82
1CZbh8+VRwGQ17duQ297n8c0DwnevCIjzY3+Cow1mxS5iN+23XJ/SM9guzXnrfWe22tqx+62gOkY
vHv0CURK9vfhzlNoiM1isojyU99R391KSeUw8Acze/uucjJmGzpsnrP3q7FcXloXxoF62M7HE7FL
JY3lxuSs6EXxnyrwIG9mkrbrRVYDfK6qPxYEqIH2GQKRri8eMm6cswpv1iul1D8joODwr+gDbn1o
r+4LuDEWdTdOJkUUWq2ZGVjUnTFeT6irTa4iVz9N6AR1bietLuSr6DW/IxqWIHWvhtl3OgZwuaH7
umyvYcG25hETZZMc5pM/QaUyhKxlCsjcsNvd0AiyKaxwzUVoy8cK7HG7S20kJTc8kZ+pnUKrSH5r
npg7U5qW/zDbIXM8G26aHMdZ0zXDdNWVlVWQ/5DJaU2cF6AXvbrZBO6oFTi2wqL00LsnXBkSENlq
pc+ie3TuMoLkp0ljW28/BP4BpXYQF06lFUCTEnJe22/8GLYUUCUViNSWc22BYoO+KGX+gMEV66y6
NijRqQM+AfT0p7n65T0PkJ1q2etRO0mC3XHOHtfh6iWwPr+OSWfgGrE/udbwlcscaeeO+K/TOw5I
eWXGO6airNkL215bHDW3h03dO/hTTwghStmJKC8nj33UZccZ5Z4k30edw27k9j1z8VOXbcy3joku
fwrnZqFHjCv++EBUppzK9sVtOOzyiV2qqJfTwaVj1MqLIfbVz6xiwHYMgj7bKIKLga/vOlOFMI4J
L+49Dnl9u/9lpB8f5gITfHWcoS0Cuk1K9zOxA82MjTRW+IAcMucRunszqNy56GAb3s16Ahh3z9MQ
B05yQHM3sidRncuk6T+HcRtCUOsgTjMhlcGFc5/cV7U4NmZ5gCQAuZcN7oLAC0coFofC/QYiADRz
p62zFpSt2SjVeMC5vwkQUxqWcJrGW1Ua/MbTvBo5fWK5gpSEy4uf1MpFEgts5cCcoLoJolg7fuNe
DEEvWHe29GMk4Wt5M9TxNf5eYdHWfPAxYC9JFrXjdd/EOeE8auL3KphHSaqz8ecUxxnaYuQqPd+v
fcKrbIavwshJqND7Dn310fYQaa1u7KkJTOL6B9nu3VAeRyKeAP+3S95sTtf55kg+nwjF+HDmeXYI
GzqKSz8iLJ92qP0Nrcde25DUSyU0WPVvvt4tkPEbPLWMRDIFGJdeb3+ZezOa/Ibt6cywVN4eoa4B
Vmm1E2MG4ln6RWBKI7ZRmhG64kTtVvgyyebAd/kcFkaAY32/BGDuxQ2AHQ9tG0KbgNgPcaiRkRj6
QL1VgUvbawzLGXjOXRzsa9kj2BeSAXFnxhkDJkOi8AG76Eycu1svsRqtSQ/fS2FAHICf+wUCO0en
Gc+7A951gP5NDNlLBy+6IvICh4fNdELENNWiAD4Xj4YZnFhV0jxfzb2JNryKNYOJXLWQaM6cG9bt
1YRwKZ5h7DvZ0kdxnHuLOzc4+LcVI5X4bhldG3dxzb0/EjCzHPuQVDL3d5axIpJlcMYPkmUU4TQ/
ldrwc2Kd2cazFPE5vynHpDqbb9lm479Mnbc8s1B6OMkFj7QMa9FXwzTNO5LdSPLrA/AkVLUynKw6
bev+pjMy0b/KcuHxRR+tOFp3YwMHrtjtCD03sav3zPMzsHcc+IWFBcO3128SUMzjJQ3fdRS0y6zi
BSJU3rQUR8aT9ofzaHTF8uY6PNGhOLqiYkHEyBuVRfun3unS3gnf+Iw48E19Tdanvfootdyrovo0
MZCVPW+Tn7RqL+uEz0UfFOiCMaJuqEqo0pHRkpSSpctQ0XQRKyXfitWVXNjNeW8BmJolvq7TU1IZ
nRDB8mYy5HTnQl1YDnlJUseoGssUJ9tu4/b6Fi0HG2jAt27D2cWQ1THJFbmf0bI6j+Ud/iE5euJN
VMOGsuPZiMOPBHG0Ag9XeKnOvm4wM9yQMomhm5dxeflfcS9sy23eI3DkDfODESyvjp432Heswf4a
1J9dUYAUju0XkiP0/LVPW1B0UEo20YnxzVprU45e145db6w5IHVYAFwhHr/E9QXhxpo1ZYKuU0bJ
gzmBIENSeSC8PPJywzTdp/y6ah0tTPyPK86Jckpz3vgvBuzqZoENJ6sE+ws49I43G97nni6048Um
VQbRNkfKiUXuVvge8mh6PnGtxGAUSFZBZzXGnaA3jIE4ITNfub0ahEEA3epcfUaVrq0mmmHoUvjZ
p43RQJQ+bKyfwnuirTqwEtYNltygPW2CH486+t08/57Div3btbRDQGfuC/N+nHzZVJV1MrUpkFGa
7PJKAR6V6iJ7ainLmvQwkVRxEj+RSO68cHM6yajDTIts38IAEt9b8sfrXwEoiLr9UN+OMiiUd/Go
7BZD0Se/KZ4VZWYO334TufCEVlW7T9qA/I9JrgIDxWOeNEoZnyViWcHl8Mi524DbrZYKQqjdjNUD
oMXro09mZ0SH/nUFUBPJYnZLNS4A56G7HlSIxrsXy9E9wvswI93pVrFVnlglCKYzMgg/utdjfH1p
4dB6aFUXHxljIY7fpD5U17m+A+cr3tSglQI+Fo9F+ce+6zVB2pSp5n/q45oVDVCqdtcu8wE/b0Xq
LPx5eyqofP8Cqjh+g/18N9cPNVsX17Qp0zvFTMDyGCtuODSfx5JzMKKWOhOz9ahO2fUt30xZ2TMY
S9ERPOHi1KRFl3+qJZGqOzTsTi4OFwPD1jBAnc4ukBrpO4b4iaJv4Yt7fR/3lazLVkqB7AwAxDlw
GOgVoeMwvoQq3xhgLuklr2UIdRJhq+WUn8HLliduPQvaca+2f5w7C/EP3a1k8sdKiBhn+XE9zJKl
Ag5OPBWIZqqa2k3r8H2+0HOY3nfqBcnLEqOqrveiJMJVP+WgWjZ7XgVTJ1fmTzUZSzcOv0P8bz3w
wo08vcJq5CfSYhmFSRkK7e42hw9UJP9zNLRIg3Qf6zlAClvlQeU6luN6RE4JjopXCdCuKj83Itvl
R6eu90CrRGVm3eJQSrnZ+8v8lEyuoJpe5vWwYHuRwSEe+iTZvdqjq5N/6R7YH5kqHPKiiNvJeQSx
eT789N88ude+vkibogaMiic9PAe/FXCkgx1DaHooIRVV+Kcb+AQJpNlkoxY+JOQcqPOyLnTMqztr
7KZzCbBWiIa1v9bUp51jXO6uI9Tc232gl84K3C1VUsVY/1S6vAY2UIXSTfK/yIfFY+wR5KPNvj87
y2JlkMobeUAjnimPN/wJbijUiPzMxtSKzGXRQgzmeRg6HZ2OJPLYcrl/9zgG/m0DLBSqr+16VoJP
ODJUbkycm5ljYWYzzWPSFKzlXV0LQ0gdi36VVNddtl3SRuM0nGuthcquUITCUl1GHTb5NvgyqX52
gmAvezj4/Jtp39QjZ8WOTilJxXbRhXj29kEcNpg9BOtgUFlfrxlclMNQDEH/cB058RuRXKY5INny
Tpyc4oEpeifXcRFm8Z594mldTRAEtYSHebyXgoJHUg9XQhYz+mzBz6fqTi8tjejxmhuMFgXLOB3h
KqRvqW6jmznmr+xURbWomovi7TZpEK1OH+Rpj/DvTYK8FBnM0HxAZJW0fqEHqyUryZxIyQbVgI+z
Z9cUM6b5O2/m8aGF8pR4NrpLfmzoHc9I6yzZXRB5XFXGYxXs5nNoKf2eYjYC4wSs9n4Zxd7g2yM/
AY8ghr4nZZ/kSlTTvw4HFR0/luOTGuBy8kBj7bAqVjVKRLZltBYRXiorxRF1Bl9h2DogS+3iv7OD
0LyEG45gTt5Fw0eaQNXLOhqFB0zIcKYdAU6ebX957AgkpHNexcEPB1mB8XlAzGEXMAzY0kf2ceT/
OvUE1Aa7bEvKpN+PDDb4RjKSXCU6dUuseVSegmuNttxZIO6QoGQz9fUiDB8GWb4idp5++k5HcWCt
g1QNxpvmfn9DqBIEuv80tOz1wQlSEywoJBD29f/SPpwIwg6jb6z3VsNntigaHsdKMJApE0c0+t7U
/fSajoAF/8m3AIzjpKr9EeIho6q/WqHCSSG8FcJGXJeQsJRs2i3aosRXF4PNqRFdmWM6y6BmLhGB
eEk6F7eIpy2ypQxpbbRk3k14O55DUfLDcOMVeRSR03Jf6lHmmh8k6LeMQxdoK+Vx+6ccucfFbwVv
Thq6h5VfaWkZjsj8CHz93CpPHRa3gYmxnbjgtcj2Czhasq6+/e5nBB2Vqv1xP5ugPMDT8LhOwz0F
0h9gzjiLLQ7KxOaMe1CyymlQWD6G3YTKil2bOu46i0dpjaj3Xqr7PGVjAHZB+Y9Ob2epdcwyHqTr
Z3bQuEgzYQ/ucTMh2k+qzp5nUPmWyQZ9sItQdiwGoL/rtOGdmZrY+8n8mQb+Noq63mNa8eTUeE4m
ct6YeBRJuOc36S9D5/mScKFkjUhsKOslDVjCuGDbe7vTK1idIYDjqNnau8LkwzvbPcs+eG81oLAI
NcV0pV3C6xe31ep2dJoI/itwUOfTdVzuCmZ0FhqBguhFvxla3gGgOkW7bshPKZXFvX4E5wzQaMM3
6XdhiIHsZaWA+urk1JZ9c0j0zOoqz/P0KVw1YD4yDBhndGtNXTXOqUHeqJ1z57oMR8IbSFf5q21j
xbzPOstrkIWw/nvg1nuI+bK+50gMmPZE5EQPycxlVHtuMvwTjaG3zjcZ6a5qCT331x6TNFKSOEn5
+QWEaNzFH/Xq1CyKcjmUtLqZ2DhiCi7POpOpydVHlMsoDUnO34+mmKRRWDbHcZkq9PfUQUgbTkFw
2lOMZBsQua27Fp6Jurlemm0aPMXwi/Z5TOtKzh39AiNQkC09aafkCUZsON1Kdgd1Ppb+PGTGL+KJ
sz9LGudJAoJkdZrqe5vUZhcpITtJ0rUmAC1a/luKuk9uQJ7PiW/3mo/cabueq/4jmOTAsbCsjEO5
pkJM/cdCUpKylvhBYaMrBaHymp6Dod8u7BhqWB1ROslseWqzW6hGj3fYhz7lt3y2TCcVVdhVQbEO
NXOrwwA6EB8UxfuM1y6D78TnKZArqVKG2Izt6Hk9ad2t9sxuZ1EH8HNh0WyrnTw5UqnrAVATWPB7
AiFfWUeDTO3IA+YX+5T4Ydj7mWjausiY3az8FlYYiePdJQb5loXLbxvGnZBkzcyYsnCooqEeFecK
DfyybnFmhDGaLCQ+w5ZTEUOqLhDG/aXlMW+yaxaQx9fy+eRktFSLFgwtn7620cDVBuJciuO7BDLR
aSEqPL0MfTMaNtjKfoIEaDJKeWlb6wTK4zgQNRE2a+kjdWVRcStdQnL6bFtsY4vm6SRYCSu9OUhH
zOSVAZwWumJ6n7P/hlfooh5fmR0F4FwyXZAX3/ERjBCOmUAT/ON8tfQFMf7/LgCH52BWZu6kl/4C
enP0MKjl9IpYsXVdYWzl0JM4HCtWqSaoMsdO83do6TjC3mX/3OXANjK+Yxqr/okUO4Pe+pHSAGjY
MMsvyQL69Gnyg5pg8K4aXY4Q1AxvFvgEcQcUMSMNkwQs7jO7pRZIwMK0MhuK/3yZee+DkdghFS00
7QdJ1UWPB7x2yafRs+r3yLTe558su6u7vT/t7Ln/nWYLD+JmMPkWX2mGQRy0yVZieyz+U23BM3vk
eX5/kD+KUWMg4hYY6Vk1YhEXdq9A8ecoF4/hpvLUmhIvXbTaKCgkt1G5ABU9ZpkdMteYXGTU6cX8
6S6fXU3XjYJvtditwyMsLmcK0VAf/WO/dg8amnaLg6QU6Rg96/akO3hx5OarOnQzpHZcGJB3arCZ
d23cBKCSM3iY9OLAejUIGZP+5BSvvwiZJU18uePqM75zBPw1M+AsPWtinXFCF8ZzGf6kD1576uwy
ZmAl0eFDmjSRNyK43/2q0Gx8QUUqOGREYa2LC6LCWTbSn6gRi7OguKLgg0Qfxiy06XR7PIihQgEV
25KId0mBwbzB9CUPN44chLve/vGH6yjw2Z9T2HjlBcT4AhHerMGM4DpRJZW00s11bwVvD90U5SVB
Ly/qLAjry9j8bEXy+VeDZZiTAH/oGnMtAEf6in4y6K/Fw+4xIYrKpZF+0AU4cfdemp3nhIQp8mME
NXeeZnUwumSmeqeCHwG1yPV/eSxjTIklijyKfUtofDmqRQeSHMmnT8cz2NHx43lBL6ffm1cp2XSf
h9H5jq2zIwbIEgbXLTRbCf1QIrY0PCJDfxEqWRHnSkEte2ZLTS9aEiPMTVj6AXbxyweISHtM0OOJ
qon3jxoiuBku5jVLtnIc/jQiIKMgocSEIx/gEFPd6/OWjgoOn4ZMboF1rg07YBmcXqCjxTKEhdJ3
85D5U8vbC17rb3VVrZPxMiSDQY8Q0V2myHhQv4sj7g2vOseGGiIYD2U+IDcxJ6wDFR7ZdFdFggEB
JZCduqFouSwaL4v3QwwbALeBvYsGnAVqLv92ivBmbJ8kjun1d/XuyyxVcG4vqDb2VZzNmVy+UbJG
wpPL9F6A/M4JExu5h2xaiiybNgIvb0EBMVf9bVR139yVSNm+sMpW2sMS7BvytYmEHhUKZ8pi81I0
3YEXEevuJBZCniwCOQbJ8nF1rioJFzMWi35O9t8d9ZVj4M02yJlRST4Hpvj/lNeYst4OXlhyeADy
xTXK0FnosldlEBmfrmdOUYM2I4O7OGfRENeUEy/zlUd1w7YzZg1uNWoY9ixiHN7Jgfh1lFh/hgAJ
Md9ahGPX6BO818y72YHmbPlYIKCQbkHaViHarWEviLzB6xgfRkYNM+6FlrNTm7uiQUG6Dy3/HHjA
U6OmBPwD9vyiFuXyyYykjFwtdy0XbqNoXJvUFcTtWbCPjDkWjd5yMhZQCqwGdejCLj20gWiJTQfl
3poo95WJHfbghm9jtXtVxP3dLEkDuhUJY8wdo8tIlNnjiLWpyNUgHCLhfnGZt3j5WQ1Wu/GOEZYQ
uAxHYXRrgJ6Mcn0QDpoXozXI/axqwtVD2a3+Yf1B1w652XWXpxp6+4zzFsAQmBeKysKFQtSAtg3J
KLMOXUbk+GaPJULroBGsEvDnLs2tqbKYdzDgy2npLGr6vByh7SZxtOFZU+JA972Fi+nVKx+xjNXG
CMC5FH1COaJmwU4jMWAVLHUlS9oMeKNuoIqEqqVcyzxRa7wcaeWbrIiQLA6jUarG3iKYmRKLFTs1
a7aimWFoOJYvGTwrTWDu+3HDUb8BD/gS7vbsub5hWv7kp+bCoNOYtfxMWZA8eHO6MvuXKmsUjNks
JQ5KJk1tuZOcNt9quhlQ75K3c6+rwqJcAGDOISSfG4v3ikBz7XRPH2rpI6GEbpiAzjRPg6oeP/iL
ltiswzsCVv8Pze5xarAmfZIJ53rMt9hIv1aFby6cWO8jyuWvLlkhVyFEdhxVjhBImgUh/cW9OCuv
C7KH1TaPP2tz3uotMetOAsbmkPj89guzuv4JAS9VqsM7+zIAI57jQ6Py5X60V0PcEVO6+gsqB45l
CdbGDaum6EUaTOrLU7ZPQdE1fEbhgmxebEHU72T2pdYrnhMorhQbT3K04sdVeY5StM2tjEs2quBI
c7L/NXaaQ2T2a+/Q/vKea1LZWdQaaoOt8pBleYJ3Ok4fheHWsOKjnD3RnPAyw7HZ7OaKMu8p8V0x
pTGrVqzf09K8VPtUVp2MocTpQwoFjw5KS1dEXjM0RKOnLsOQRxy42lcuKSRD8o9uVwAAW/Bmh+5z
8K9KdkdHU/vU+RpzK0XVlJe+dKLEyh596hq2xnKC4qWWVAK21m5w0A8+nAxSE8uumlYNXukG8Gzr
QxT032GndImWpgbOKIRhcypBnpmk/xzRCiHC9ntw1Ovu2gHa+IVBAAZHhPNkt/wNSUsXTp4DcWme
cBU6BwZQ3S4MO99l5/705CLc76PpdF5OHiH9kdla40nBgIwalxYnazg9Bh4i5BrW4czEQXyBlP/6
/ExFcjinK8dZeC+/tHdzFrCSR3TY0lNgZevbKdTkmI2vM2nW+xLV9uA55I9kI+yY1RH6cZf5yJHz
ZMerRvuYtUjoCyDvW9F8JGqU9iyp7Zm7F+5RErtyqqvHlnZ03kaH55Z7qZ+vQoT8W88E+IxKU7fn
lvkVK3Yb1iVu2nuC37SpOlYk4K8rXdLXZCjX/0qpTuImdACa8vY0pvPE0nFGcRIaIKU3YdiGgRHC
3e9ltcSnghxfNzS1hToG9PgcCN2pYOtnPADoHTh7/qdfTMJsFOni/mu1PaOdApjnGtcegK6W3ZxC
YUgLEe5yVs6wpXNxlfPjHf1v8scepqnMMK/bDaGNu2zI33AH3mMonFIN84TC0h7yPg9VGRHUWePA
2yTAZdO3FbNcdpfVRdKxBLthVbLuINBBLxbOmu0NgxXPsqoNtkgRh56kbVNv4FLP7pH0YUgSIA4j
41KYhpe/pGiTv98Be/7ICpGNN91dBhPRg8m4P4ePO2LsYUxbsnm0v9ETspvpHEyyiGpIAzczymmf
+xgvVJ0yRWY7buR2nIaT3/a9PfE0jNtYWnxmYw3BLNVsHXEmSNlT2Dt9qWVdfQuRIZIJszf8bWdR
F0VSpcJ8AOVKTPk3HwkRjmuKwshBADYD7u0B2L3FMl9DDUMnWMWd7EbpRhCi9qH647Dw/OQynydI
MTRJyB3Trr6B6RzMpXKoG0aLzLV/sxPSOXTfuiwDtSkQhIlBdbKqeAOhDAXFoLoaQqshtF2zFp2V
C1M9efMX4f6UYPfq4yQfmVAs7tXs405n402E8n5m2tE5m5NMR8xMLfBrySCOqBS7LrtEQMNRAcsm
EAYPViupcjYSjHRmxV78mEjZ+hxArCoJXr6jG94j81cHHGnD5n7hz8ab+bMTs8tFfdlc1J/gqu0V
HLSp5tJbdEjchLpRx1jErvSxPFNENhIJe+jCR9kmNlILXGjo3PKXkF+3iqlZvZiD/LyNuJi0EAwu
5tHiP8pBrA9Pnl4mGLC+iLxVaj+Fc5RR41wpo8xwytYNRfcJQooZxy+Vh3tvPUDXqzu3hRqrm47B
Wlu5iCdgs9gFtzzEpizuC++3PgdAmEHfsq/faVKP3r5/2RY5ctwg9pVF1Qp3M9qibGDcqjsiF5Lf
HYQvFJec62CriGhik4SvIdtScj18MD3BHrWdPy7145etP3lLTnpKacWkTmkZxrAerAfOGa4ppNPz
idpE9IVSaaKhSCfdT2+Qdd9oQ/cb55R6c5gKZs+sMUArk0Gk4No75GZQ2PnRnmg97Dy+4mSEYi7o
vrAWCRHfNW0H5atQM72S+KpoDEF/QBugOyGawp5LdnZlzzNTxBxswfMmdI7o1wlWncNm+vNDdye7
176pdkwikzjKqrcbb6mlezki3ZawKd6y63uOS5H0W0nTzgdKFjPCBX1wtPPBoZ0ynt4a/qz+/au0
aG50rLVrjtI/p2N1VsoGsjrD66Oml+yZg7Eev47gIKTU9W2TqKofu5cY5iJjV+VevW3l4Ru2e8Yj
i6NpM+lXPoy2hOlnKFBgkc4zGW/poZaSWQVaNrfLOXfvpNJyhtLA8xl3Pfjh+mEDPpLuvUh8T7K8
wNKv8ZaRKF6jCXQPIzHx9dwbnZrXMYtbH1VdapGWyoBD9wjP4/6yy98bT0ipyvHPA2iePE7W0N4J
mfxhcu7XQ2b9W1JiRN6CxTxbL37dRQwuPGF1CixcV180gnY+LOFKrPDzmmHiAxsJwXEExl5j7TlP
fRYwsqwzSiEN43pBlwKcPeVi5mG4QLEX9dETQu2XPzU9spkN8Sz1G6LGc5/hcRJB8QL9DUxqgvfG
2FeDMl0nhlevl2esKNQk32dr60dMMyeQiYufypDh4AI2Dg5rUMvtpUgB6x4HZCKSpjmNMzRg/UB7
wfL7RrOu2/1rva0u4J8QoNyMpjcSSEJehOhIslaonWyiV/nHPRiGp5jnCC+s5aBAtypKY3GnBiIO
8hB0gHB0Kog/Q1q5cdCHseL+DnChszHK7F6IKW9++D+Jr194k1NK6wXK/KL+Xi97xu4pgKHdktIK
6nOEqBYfK005TTdX7U9vp0ptCFqh+ndbHpJKcNMzf80YBBDcS2sM4idJHcnJ4Mga4zJD2O4SuUQb
FHZtr7Op0mbO3boak/LXrzVazdwq62DszseYarDqXby5da3EhN0KnvH2A5tkAkqhFXdlofpeRaxq
kXco7ERo6lneTzo9XBsTobQyC7C2/KrkAaRME5K8pFYuTvjbtGi8etai/61EppyncXrMwMq6P8ta
Iqv6Yk8+EvcLCn/25Wlk7l1YX8vAdNFDgrfwbGhxUU/anMmkxoqwUCucB+tvboti8RPAiTa+uZ8F
qA46Wr/u4qRYZzaPqT9+qlPqDQEwuWoBGdJOoa0e7pg/V/re9TEft8QSvak4p/OYtUVpbSoYboDj
gl0i4rCPaQmqZGaagHQwvvpN6ycL50EhfZu34xhLVkKT3DxEdSpDvOhzdNzl7T+IOYl3lUDMzfoO
UOCDV/q9g1eN5iD3qmyqGfJz1T4BqGPfRnk/Fvgsq/teJwVT177362X3vaZLcvh0jqAlDI6Pi9wd
0hiUBtLgJox/O7jh2L5kouXSQiRE3CoQ41bwxmTJpj+4v0Sg0UwiwNBt92FmyZFKRhKVS+V74LOj
18befCfvo2XIKwPOxdAkcS+xBMgZenFtklqT84IWoFhijX3+NUFJw7VxEi3Oy2sHNZAqFZk3aBAa
RBWZS4GW6N4wkGc5lRdwTxWGufzmILY3XL29BEXhbfX3FOU+2dEYRqeN4uQrOSYjbBR30H9o89s7
GJaAZsm57kQaxgHPlRw9pN6J/LF9hKWJ2NzK3ErEGsjnRyA7AHe7W/cX1GU3IIq6uQHs6G1Kg+wm
ry7lfZouGMdOAXTfSN2Z4rBoquOkJeL9KXGQovsA89V1ffYpRGg5RqnmqjZ1u71Rl+l6W1XQaHJo
oK6m0Tx1M1JDx/eoy31igviHRlDdqqAEmUF2D++aNqThHrveOjbPTuYClLey3EkOLXw0q1hyn12M
yRnxtaTdu0Iaw+RLNmEmxTm0D/VSgC8faQ1f9KtyLWMN4Vhh2m2SeOyPNqtHEdLlCW2a5WkJkNUc
ybUh8/868AhAYNKKsjygYpYUJSdlolqAOpnby/lkmX1ATyRvpSUcWBDxhtH16onCm4EQsfIPWqWM
J1wIrFOg7Dgip9H+xUyec3mv8sieh8wkjdHdZy1R1DdpW1esLQSSxBJJODIOu0XjUVkgD5WjUOqe
4Z+BP7TFhgvyIeYugny/aHQyXbEbXV23DwCQibzkzN3H7OV+qUCMgPgb7vT5UWl3OhnOBLtXADHj
CC+Q2lSeJB9g7JK1QGr+pDjKEJbOSPkCei55CdSu4D0iATUnFA+R1BWuozYDJirinxZawAW6YiuJ
N7YhvMXPRWRZ3gxz0qg/Gk2Jm/bLI5K0d8G0RyfaR0yCBHw/igjB/+UQVyCe+Gi3gvsRV8whJHQG
Aj99xLnaKwGyjYuv3pUy/Xps59GwfX62w1gXQH9mWHRUmo1SlNa+zGkDaKmWSJlupqzD0CE7qBpQ
yrzkhQ3qW+y01CVFLPEkpsFAZGHszhRgjhzwTkDg9l5czLMaKKWHknnFo0Ny/a+eOxgGb5/YmFV+
369dWLYkOuRBI7P2xIxQAsrVjPx013OY08zB6m4I5FcBKZQLc2TOpp4/hmhB8pJ65b9rVAcRQRRX
PwcyrdYJIbkfYCAf2OfCTrGJfWOyL4nxG2FTfvsz5Btf+wbVoocz8e/32ixpWrz+I3lTWsJqjjO1
V/Ywy9V+Oh1gRjg4Anha6eh31+C//1B2lsshBSih2YxP9bNWpeoGokvFTnTPa2fjwj/c0QrDJq64
/5gLoEpnurT1VDrfy4W01LYONhcnXQedBP/SkXrUmeNVvi17dzVVs3tqzuPbCMkMVxdkr9sWAYIn
KNMnaWrIf4L/808d5DFb70RFY+nPT3nE0eFlSPUbjBR9s/fELmQ511aQr8tzSRYJd6440JLd4M/n
YR2Tpd9i1qXV9o9NnoFzR8d/zQTNXDDfArvtFr5K9oVADbx6zPYUjLpRE8EoliF69OQyNT4J2Oqa
7VS7oxGg9mn00fwlfUfLwNSATkVIG6Yo9vmCB7ZfYlsJU65mEQtUUj4pSmNcwTSxbenYBXvpytIQ
1FAthfSiZxjjygn2/OmzOY/MSUBGCGADLr/FTZzU797bSBbg48NEJtHjfo7Zjiqnim0PMEN+Samj
hipXqy5GKi8Y/4nmdYhWAwy+Xk6p/NZxz+9hgWy7r0UBbD/a3lqzuUEnbgSPaPqr8NZuNScRRnKX
1zlAO04PQiEoMWKt/eLN/KHUkYpK8+KWMbWDhNvzHE11fZyZJgqgUf8aY2ElxwqwcIJsSOUHgJSe
pW/cLrZstNfgHXBioHE6yPInRtLZv0xjKXcJwLOoqshGjYQCus524XI/78eAsEjtCnGMau2dX8m3
hPN+yoQzUxf3WN6MKyuAt+F7htisKACJbcXewcGEIXe8j1w33Qf1apfbwPh8YargEdRm9IPtNEjB
8ADlKxj22SnRV6S2iwiTEi7/JPZ3Zq0UTD95QZ/m1rK/dBd0sFg8RxzNSEGZ0IfHV1ZjT7GOKQbe
n29sJyuiuNjSk0N3iIOUNyuYQGQvbVR/VM83zNvlN9uy501JxX7H8CDJCv6gyhTOag1XhHJypM60
NmDfDlLl6Bn3u4n6O0lLTeQDyasSVRxRz5KFl6mH7MY0Gfe0X3UjNvlBLq7LiGSGkW/ofDP5FIZ7
1EkIID9VSRloy0r0Zahd8m2wRV10wami/VYQgz45OfrtuuyibRH0O106HK62qru7ZnbdobEEwMiB
PtQq+fFmVtuwo58u8UmLsuUN2nfugeV4Q2GAExPv2E4JwGwNCqNQtgF9cVoioXUJyHBWfd8fVer8
kte9CCB3VYoUUzDUQ5R/w1Ip33zvc7KKQ5cEaetUdoflnynw8a1xO35ZvADiNHBGE+UZEJuUfFrt
PUpYJnH6TlEVOa2PUJ8XeiCbfVhV0VdYOSkoh4aWRYF1QSf9PtlvF3x+kJQqM1rj2Cpa1/k09h2H
UyMupGwNdgq8NSt4SCy3iznG5BNXhtvmdb90C8tx4PmVmATXUpm1D2/MUqsw26WSjkN4mJxVswC4
GQ3Bhwqxq+tb/yQ/8+0lizYMJLzTpCLp15ohOI0UpxRD+JfKJ1GRBcgnhhrKDYnKXWWAELRE7pf3
M0/jPoe1J9qCk8SuHQP0vItm8KnrnKfchXJsTtNywhjHVjOzmmjRKg+/dqQujlbHgjrTfbkhpcuJ
jwNkHkYDZRekoq/VwEb0KjqIqRn5XchKLmVilImEg6sUbyIxAgmTVcaOi3stpYJlVMyyL5v0emeQ
a1GIimgOsJgiPO5TkaIlUEKiUZp9v4jgltp3wAWY65hqedfIrYnrUOmyJPI9OP55hPPrKcJv5vzT
j5eWUKmP3wLRFtXTsEihLXKtVigWCwOhrweyIyosMy9wg4XOlwgZguZhtx4KkanmBv2HmXrRElTn
LbO+SHuWZmdNcv0She8vcD8CXJxpjXjsy0Zmn2jWNXGABaNItAMdIBksDJ4M9TWYcZ/IJZTuS2vO
P170rWsCE1Idnf44NVDfAlGce/QE2JSzIA6GvN5EqVcDqkQMK5NJRU7OfdoTEMBzuEdFQ6r5Nf4X
ECXWWkqDKQV0QC3PbsTQj31shrgNe+4zMkyuBAKaUPZ7XqP4MHUzhupz8nVnY3RSq9clSsWrldNp
V9PC/TpHQBvx+bHf2nd8DauLfiX6/iU7QPonoAXcEgjoIVpFan8oI/51MjTGedW5E4huY+ORwFX1
/QlSoIx/AsTYPOR98UAUDazvSMH2jUqXRs2BWL92AczD8Qrk0ik2dGjlbyzHI8ZD4Eg21HkwnJ7i
bzLGn4XtHau12OesqmRfi0JehSbVejFLqrB8hatW9V+l76lZJHst8cnnGd+GWGMIJ6Rm1TFBAGLo
XzE26oAbUkY9ni5P9Jik1NSPScMlvY/Davk0aTGOZufeVBRFpEtV4fyaO1YNscsG/vi9O9mvHfzW
mlvjvnTuAvDRZAEbIdC5tF5P4oVeGI+wj1H9aV922FYsrDVzsbE6TJ/lsa+SXKyI+6sqcJDQ7Rpg
gLFLrHenvfnT2w+Uh3PBSNV52FcFMbWP1WDwmkYsOndmTdPebDgeH5sfqnijp5rlAtFL0uU2nJiz
Cx68JP8VEvxVLcs3XkOchlGuxRKGV2QUUcwxvPGljMtREb20Qx4UbcceHzPJuKQcg8oxtUAvNwE+
7xdC+Sm9o48CZwXl2ySZ9fzNoxdq5sG5xPrZI6cL1wCLs64mh94NkvSeI8CKLAvcjzqcFHpLY22P
rn2Bnx82CUFd0jmH9HQRwpYfiVZX/wtIefbb1S7zbkk/4jFr3jY21Xmv8hsNrLUVLzvDhKs2oZ0x
arK3dJIqsV1Ihv0NnhIoe0g2Tbxf5ng7X2gJSipTfZf1QliOJT77PZEzp67Rnc3Nu9nbelVmLvII
ZoVmfHotXhBK3EAfsm2KkPaRKbJUv7SQDmziw+vsveOUCUr7ubCdYRUcSqiCtK++B4UoomAmp60q
kTY8Nna3sDyO+//KEl4DFrlo/SYh+jaOFfXvN+gRc5sBvOToCh4qqraxK6sRix5pra52htHbQH7/
6LBYlKYTzH4ZIPvz2vlvcJPCAhELPVmeudwt78qODBmm+clD9RpTfKrFaHzMDqn+/dqFK7DUwekl
Rw6ENzsbDpWE/ah0cyllT+igYErVSfOv/NMvu7jUNeyD1N8QxNvV7b5tRr/SU9WkZK8LOmwq19CK
yY2smH46nDPSmWHWwAC3Lf9Up3VAhra53C1e383LWLGl1ksPrHip5jNYYNG5ut/JZKOirTxCTv+e
7C7i4zTuXF6NrDUY7Nnt2LLT+byNVHaIogjbAfmWUSsP0el5AgivHqdC6komi0aNQitBE9Uv5mU1
bPupdmTQcIOZMVGVLtpX6/AhgKs1YkuagCLwpdmuiyyGzZ7jxh2zmnO8zueDVjsFDaQlW/d3QhN+
D6TeEgLKr+si+ypnYY4hpGl/YYqhY/cbf3FdGc+RSYVNllTbWmyhifFCQIii5QLwuBOpmH22EOk4
uByCT7Hlbn8BktMwFafJ3mgEtLpuQ4NDd9vikHSfaA1UDooijx2hfaAs4c3Bjy38Sac4J2Gbk6Xx
Yr0veBykA4P1PZdwAV9WspsSn4nznO/f8nghmGfQKLfeDe4RQMQodnPfms7STyrLgencaHIrhgeK
phsDW20DYOGvVaosRF9kLp2SPcNiBO3FEt2WfUnqfUEmLKJrRvff7VbVxlV222INnBz6WoxAZpQt
3yJ8uusBFvfY/S7piYHMIADl39atI+1YuACNjeQ+7eqadCpDOyJaMgyQDyumzKg6Grh+qXM/tptY
qDnNG5McVL+mWeBJDyWLRIdMphUeKIjWam7jd8cyQti8hg3dkJ2f54eTxO3t7VgHeV0Hvk5nMLW9
IO1jKs9niZwcT0rwWA6XZvWh0+fPqRc8GpuhfZeioW+Myc4wqf8eTqfwQKYmsGnVcJjAOzDxtgnG
TBe9SF/dWm1I6QtZzXTvjCWTjNCW3fhxgIe1ADRSwR9ammBY/SlyN0IgqA3Sq9GaCp/atNamHoW7
kxyc8yWe4fEil6wUYqRInQRju95DAznYUITihb+A5I1Py78zu5PgJIxNZuXNcT5mm18zpJNRTqXx
Z1ZqUPyk9oXzITg+6g9Rl8H97Rl/FnUF7K/Pe+3bQN+4R2Rtla7ZHIq1GVaHmzL1t1k2BRcV/TYC
dTCX3tYgsyFQd95auzuqukOmDO2kEsuALoekRLI2RUcgQ7ucHQVQ+VFqbxym1c3cThUPqyyfLTp5
7Zfl/rDrKACK4y5EzNDkIAU5SmC0kXg2K7Ipu2Sjkpb037U82h4sU+cHUbphGaGIxmyGmcnVgO9f
dG1yW2BKMeWatq3umQIOhl/2sjCukZi+QMeJ24ozKQgdaJ+Bw9DXQ8xdO7bbo5E6ShCvqOlKnpV0
Tq0mqbWgNHAvUxlP5+S6C/ZTizyfuYXMYM05eNLPqAUSri3I3rc8OeGR4iDCIjGLXO95r25nYOCx
9PTCTBJhPFw5EXi5GxLSMmgJo5z75HXleEMBxlr8tTSrfXbbmtmCYKL5nKCaSyH8kL8HnT7+J+vf
SGXJvJRw6Cg4bg91mNiEECqPlvWN7Qc+sGW4DxrWnBQH3jWQDrWp9I7dx2WkWtPspClKPrDoChyf
aXKPGhZfFALY7ebBJ6JcpOo4dS1LGgofQTxMDcHxkhI4HkBGgrx3G8TBtri9Luiypme1dYf38Onj
Me5zuT0aeALWPjhYm96b9R2f6L4hYmqXxqrg6VcwRJSWROYEaYOstOfXM6sOFbzBH0HQeqDtDYlv
09mdSYvGaPpwG/Y7zApzC4yQ/iuRS0YVBYlJicjY2YDMAwmh8xjNZBLVjSYW7a3MNh6xPWK3kPYy
NVCi2QLSDktV28FpVMHtoVfc5B6vb7xdpjnf4hlGCX8zVPF2QS56MMw0suSsSeRPd4pHJPrzDjaw
+OY/cbE3KdB6+Gy+i6DqCD4usemAI/xmUBldrkg4oM4Dv2/A6NBxxItUV0A4e3GfvzLlKvP1CyMP
3JeWXYdOLwc2G0n6AePPUdnM2updXq3895gskzA1nxupgE5JaNsTLzl4E9C3Rt9YR/H4pmhr4VkL
dmynkjZT6H28/i5SAfCQ8u0gIBEm7G8vyRzWgUVKwjONm+lWVCvL2+ErzoUgO82zL/VrxVPlPUGA
hqcdDHKmI5J5pAZMOYW/fQ6YZGqnKtGnQ2DzUPuj1AZcNsFNN+FvZfsuTpo1WkzeiOSsARovnv+e
SuNhfCLM9nm7NVqrynL1Zea0CHnxwkHLM5AfAO/jo2/39Y4rjg8WfiXg9klK1B7q1OX0pgunJn8K
0BiLgZ8OLOZjc0pp39xtjqYOYTvcF4UjhbHgHzfVVoE6IklWIl/w0DTf32h7QrTtC+V1Cpxzh3Xo
9JXmCxm60PqJhLtvSRQ35mGtjRX5X6N0UutuUjLdDSVBI5P9vUo+6354WnzSENfwRK5OYuyp07aT
n5wBYohRElXIslnKiKHNTqjY9sdyUL6FcFUKhmW/qJI4LCYZwl2kws6hhGtTABwy2lm8AGBrKki1
w/R0+KfXWmZPKBOReH2E3ER8rdQQeqYIRFm5HTirFyBHAjmDd+ExfQmmd5WrLXOk19g8U5v7ajRR
e3GM1/g7gQ209RgU7K/mKWX7IiXu+1+2xS9IkS1Z2vCP1PRHubzRqpiMbE098amCMtqb0zSK5K+A
1f+iVKLTehCOK2CvusNUsnImQ+XTGBliQaLAvmwmXsK1pavv5WDtvjR1Sa6lEbIc555/pg/ZYJdQ
Qt88N725Q/uuo6wzBz9xh+08w8KnUdjAmOD+McZTlJe9OlxpDX0GYAzGjXDPmANfO2+ovbz1aWvD
nYx853KBWqIV8fJUVSvEdHE/u4NGwUAtflBw4bGB3oSz/LePHVOYzdPfVAqzzjxI9YeQOYOt1Xgg
JpAzwLbYaaT4j1SrVT17Dv+4qGycvP/JJV7HF564mJYEdtJabg4bDWioNZ4+Yq5US6HSpsa696BS
wv4KnbCAdm9/PAeI1MDh9DAkzSanHJ36MNyPZoSUETQUsJhUEU2jyembUnTrLRshJ5AklJfWOvun
le4ctjZH6dkjfGaEcXV6UcXO5P6ZC7cQ42p8CMnt8LjMed3+ge4MZqYlZ1+vcuzLe2qKxeVYFglA
89MyK+skk3H905AQfpxETPM0U7r4Z3Yq0oLKQhhYsO66EwinNLK7OlKhB+DJYv0NInW+oOSgpU5D
/apTAf4OWrKBftNp4Gpg6vTaPeFe6cumTVSXRB+zk4bia0wBirB7Rp273S97Neu/NF3dZ7PIDKVZ
VJdD5hPhSx/q9diQyRs0x2TWArI7W5/q4rvDQwAiMHQErGGHYHqUbiw6O/Id6odgWxVHLvSlgkOV
JGJ5cyFn1TLkhTE3tOviZ0PoXqt4KTa8LhAMYcPl1q6aynfClVKM/zjTapNyqtG1ZCBRlbl3oHcd
2dgCPPZNV2VOjbP9PSXESTR98iNufPZ39iw5G9Jkmb81/P78HI/2KZdzZ4wPDDd5ERcBF3wYh7EH
vRc6Xx8N1euAli6ZpWPpUd2SguoTc34VN53eGsayreSKHcFA4tH/8Ifpy7Lcl7kap/6Q+uiFVIzw
HjPQFYPS6L2nsZL75nzzLILiS6Fa6rm8qLYq3hNUtpqFrxmxcvDsufS6W2di8EnaPtCmt8wE47MJ
50aJgvLONPgrleG41+u6+xEvCm1QugXGYXnR5WWBpaFJERxDeBRoGRGfmnbU02XRCzP/tXXI19QT
Tz563uPVMA5qfNVYR3upO1eVeSF8+6c/ZCjrSqv0NMXq/QQw0BmhyDO4VvZo4f2ZInzCFm9fRgCF
aK8ysVlb9uJT1FCKKv3noFmsxuI1vzy2zXtVPXStGGzaZf/B5uh7vH3loVqvBbTyR8LFcmcELjml
XMFO637ag9g2LB0Cym9eFUs4FTTskMMoD5GWkIDZL8sPrUiuD/43iJdRrJSlClJPfLBiL7REsHM4
gXwGkwksrPZSvhcGxR9GudwPUsIARokK4Y/fBn+U0pL4ObYSJl50xsHO/JrCI2BX3bSbFOjj985l
Bdz5wKO4FhZqzJiTO/dz4YH/ErlO8DtkV/JrkYbPojJOnQxcvipkK9FGEvtqMFLgdyfNUDL4ufcd
R+Pcl1OmnCOntYxabVPnlQzkh6ZJ7iwzzcSNZih3lmRdDndXlHqYDeS0KjeGObJW9J/Y9prO68p1
mNmEzRQJpYmmwvlPAlazmr7IISWGEz5cqtL4rCxE9mK5ZG511BgN/tonXi4aCZsAXKhOSzzRBQgT
0RwiMIE5ltz2GeHPbAEvph29MdTqOiIyyArejTa9H/mWSTLmFZP6aEQUIYfQbq035JZfO6mkAgF0
+W0Gg3c7TNEoutzmcIjJXwYXB2MXOW2kuoF0++IjHaXPnWV18TdZ2ywmh6HONO7G7p+7Vgn+rMN8
UJBp/8rx9dKNFN1ZmRbyvfweb3+uLDk8aIT6S/MNZTWvOlbxBbR6HhTUEUK7T4aJNU9DSMlWjRrc
RTE0G0LiDEg7G/uM8A1H/p2TmSFEO6OVexbgEWUWLRlcWI6NW20l0Zl6q+l12HrTA0FSxfyFHP58
N/HIbRaR4RNnfiU7EwgjOKCJZ3JisYz/d5rvLokdtoeO4d5OzAyejoK9cJXKrDrUgC5vaNB8LOfW
EfCP05YpefZpB7s+moC9r/JA8Z+1CYqeO7VosaX95Te0gEECNwMDTUY5Y3tYNsRRHNuc9adn1kQb
FRk1vhL2jkstEdEFOix0eLVPdPClNPN0LGG2LTRkkg5udH0WfmpQgap9ZKPsHHATxWpIUgqcQVH9
99OXpDjogsy6mb/Ee67ZUc3g6Zozpgy/t20V4Z0paOrvjn3Iw8NCbd0iU8c1cHOXwbulUvivJk7I
zI7vh3BaNlp7JWOnUJMUEP9JjZbYK+CaOeu05i6HER1l9q2Aj3IPdQGQNsYbPb4TJswURnDwZVcY
WUQFT2H9QT+Y0s0BmxQc/Zy3yqdg0BgEo39Hkra7tmjF/6FAPyEdHDPk9IE4Afh9rFyoXp44dIJp
jZWTtC8Vh1iGhRpUVPk8xuysoxYXl8SlcCSMdDnOO+6A9L/fehCPgVBdlp+y33YioPpu5l2vdoEv
bC54E/QtW7VV6jjAxcCsaxBrcf5cJ5OVTt5OEzEfZUW0t2RInNOXHE5Dhvfgiry8GpQKIGuEFFC0
2nE0XABh5DTsw0yj0vNa7SAkWBH951P3LGEcj/ktDLfCYNjQrTp8R1hcUMLYCt14/7i9c2u/fucX
9pSZ5Twp00mxT0bJSi0h5wGfsSTN6SihZURGdRQKA6R+xq+11H5EXBQcCfHsLPqEbseLZqzOt3Lp
oE0/4lQImplUmMy0eZVc8li6J5vA/ffNLuj82jHnTlTPsn3pZX/a0MU56OvFPP92lm88INmiP04N
BuUboFSUwYwhAm1yK4XGYVfhtZaMZGqxVSK7o1EwYgPacjenY/kft6jknvU76GM31Dy63yUYmrLk
weUu8RBaikKPv2i7zJxaug7QLbJgxY8N4/YRQ/MsQNiwyAwkMM8jyoHHwAlEHVZLr7Ar09S56H6a
41NWh7BDbPTlTnh0Qcs1nnH79zonsZSLb6XVgA5WvT9WooiXkCVNrjB6KlmiL8MoZEYxas+rYbXL
ctNJvK5Xvzv7o93gIWpIRwEVtXBotGoookIODBgSlPeSy30eUK4oM7uhGtOKqj2JXX/xjGhNQ1Id
hQ6PVGpHBR0qkmcHMfoR0W4sYx4e9RBNScae3EeQKHZBM920wyoDexuvqzrFgpAp9i7t4/bCrItd
1vIF0l6jacf7RBdk4rnmbX7BB9a5aRpY7uYhPfZsSdMKlvzKKBt8WNUn1x7IIHZXo7cOTkZcfB3h
XGBtw34rrbIiKARpWggvu2JRTN1fL/wldIN2WRCZ0bqEy9qHl8ukMpaH6GOpeMnqwZmNhI98gBuz
0FWKMjVc7nsi6hHXCqrMuxF68eDCBRK9nqmrdhMnNtnjUPxLwROITSxVHnlqVE03BLmEftIqCWTF
zHw0Cbnv++u91w6qgf2ARUFNI0LNcCil8pJyZY2jmX0K2Fdwc0zeevAVBOzqdLYSsbVgq5ojFWRY
Lpj3Esni5qXwh5poY+V4WH49wTfoPJ2KRsZH2OX/Mc5soeV3N3i7chcpQE7LEfe5jQ2uXaTor7th
BkAGtGihlRY6RyDG4Ckh/cwOfVdqzfTc2pGgvU2K5KR7XZKqmMcY8LT2dVPDgPozwUn601u9nk4m
r5k1fnquJqqH57gaQ17aFrlENa2UQDM9jKG0BqoECUHL+0WttJhttX3IDEzHOcWVLolthSCthTmz
yieKk8fEccEM95iDzSyUFd18SfhneKGsfho+Y4QSfHEnIKQq/3tuc8c6IbNBS0ek/oZTNaYWpATP
+LtmAAgTJD1RI+HkvQIaY+Flrj49biA5JH9k2pz00hr4W+m+qQgc6f76sGjyozdKdHKR08FHJa4R
aeuyxAk3Nu256Zgh0g+QEU9zkWws74RpATI7N9n7I6a2jt0czM4D8S3a5IxS/y3EkQUuiQBns7HO
Sce2ox8Srb+FvbMQOnTndlqe2Zm9ri/HP5wHU9Vgi/px+ZT1icRFzd2sNOqc+nAARN+8z8xgtsdA
uGDeGoh7vMR9Dev5fE+96W1R/sT8+m5eiGhUWhWFdOCB9NmxSYOEHNhXfJS52NgtCbj6HfzYn6cM
cFlo4FAyujFuw0qD5+gvC4J0VSMtq5F1vAa+b3ZjRtAtjfJT2UTapXCX8IZ0np68yRRfW3nABvQ8
2OGI221mDJaHV57RH+fP3kxxV1swr5OPcLnY+TIstpDQ9dhkq79hHgOU1jFAXhywx+Ui5NhNwA1x
OLfqa8V6+tbLMf6mWtljLAdFV/MAIZ1rOXb27vKYizR44r/zKCgbcTIU1Go8B1YCxb25WUNqGjc+
MsA3stPDTttBH8+7LUP7wk6xRpiwkYJx8l6CnTBJEPJu5f9eLKwLthS2FQEjXBmkHOwqKq16ccjD
IG2hVl6q+SCFYAjjlDIF8GKipkw4MKc5QU7sNfbkxkKmRh2vrvdjTD3VTqnSDZnq0Wa53hSypUjE
PZte39WO3XP/wXSxzU7YYcibpn3nYpKJLg2R2wRuCPi1b4G7DoR12C1xIInsYcyXSpXOO71O2hJ7
ihu9w/Pr4hbiHQXK5QtYJLbi2i86UNGPILsZnCLW+tnAssO3JJpmRD6TsKkbibKJjhEIrmRp7E52
a8Oo4AD1bhnhcpoBhjzBuBJZIJmORwPY8zP3EwpE/0LO5TDAOdQ8TxP3h2Z3kMWWQmFgZ+8YJo3B
lKMrME2l5BnuSbNgYHcTSrNOT5JtObBWpTZD/yf7rMk32TCKsGx9Z4QpUYAUROZG7qM7fXHBp0bf
1lZgJylmbbtPwf/tppORe0cNkhxjiRkz9p/rHMK/TQSytxyrk/kXDBiTZ5kFjXetCjEvh4HtybRD
fFykRquHO6XspbCRI+HROPW1OC/V0vWSWusSUBv5j6Zk8Styx2vwkRKq6xfXEHbhqVkz1/1+qde6
YaUqPo9D6kPXF4kR14bLVADYBwPfp9TJRv3Ad7ar0TorAb5pEAV9wjiTnTkYKEbKtJkFkbBOoivj
fAOcYzwHtWy8yinbBKKTV08EXDoXQRqIBx0cxwK6Mu2mn20FTQjR5iMFqyV5CrUYQi6b7a2BCILZ
shgd3z2NEsLsnExoKtL0+V4hvEXVyvyWKFjL6R5Q74dNJsQIcFb0zhRSp9DnKinXGdUVu3okmRLT
JRDA7gTY6yUdfqmlHy4j9aypEf76Yl5pyIHJL7CjmDUCxT/cEIryCNAzUcycuGi4Ch/bm/YB/qUt
hWwsab+g4E6QyEB7vY5GKZLg8T2ROkS9XDmMIrNZ6KEMf9pJZecFW+0YacUa7Qz5y5utPhpFQC5y
/y1MVzLxM88/8nBQLalaSdIOgbqaw66LPYDyInNwzHZePhKBi9+qMNoGQhoja/twtqUn0xF877nR
vauaAG2By+DSyGrX3bvSr9Po1BqAR2bV2gSk1OuTSbbw3yThyxWIkr65Gw3t4UJPdzrNPjrD2vGQ
0veT5fQVm7YjrwYg7qgLi9p3olPed4+KgQ8kESIMOMz06B1UQ2m3+xy8d+g6Qpgzm5uxUbDzu8Kn
EZfHJY+Lnv3KZea8WoUoJx4crpdGw2JHktat8slKHs+FiJTkqPu71KPN1narhe2T7/X3LafkdFjh
4zJPcXYnyfR4smHOIm4nAqNBrruTQJvm4g1xqUwjvWj91fsVWZSJH9K2440hmaFGvv8H4S220/PW
f05q/cyNPHdfEDStePvOiLh3TVcuRijqq9EbaDn311cptweP5hutgJIqhFW6TWIrpi2yuOswJs7d
3kWbYwhQ5ARxAQ7Cb4PDWFAXD/a/lnZd/ZiSJPqxe+7MtwEV55ShwxwmZjMkC1uOMXZQ31+RZ9/R
Pn5Lig3W27opwB2aftryzbi++fDaOWbaRu+T9KzSv5LPS2EclnXgBbgBUcGAOPy/c3AlZx6dgsKU
5SBMMGnNfGUTlD/93uTUVbZmSugz+rqUixCc+W9EVuHmI6NhDnv36EIrlHMHhBy1xp21MrLrlChO
gBhIluGpQsld25k5/jdM/5UF9D3/VhkueffUUHKGxzD+jpkoyw4VaLdpH5fIsslYQNr9pXSkI/zx
VVx3FSJnnry/uoa5Ef85fUr91FwlM7LSBICwpm/abUylPvlKKnbz0hzTeT6il7R9Bf9N00VaeXGb
9oT+OwlxRQFH3fe0U1VBiO0SSCEKi2zcbk+ssyIjYwizQxLew1FNW0LUJtSz4hqR7cKQ8UYgboyO
pw0vJsvmWab2q51X9+I+3QxDnQNvLHPoGXQ2cm3nV+1EQYichqBLCqCmJsd/0Z280QD0i55oT41q
KiFw6bYu7nLlh3XrGBxw4t110cFwoEgQvDnqYN99b6O8BD31TA2f/2keFnxYF6S2qAs7ZIDvUInv
DwS6bcD+Ur2/I+XFBome71HITB9U2uKWnyJNmvux283Je4W/AVBfqHKJEjSHI9NjKSocog691b6D
m11Tk8pIdEekk1RBvUbptf1Ylc+p3yHjcir+jHU5JbJtJY0hXfNizR+YfCjmhX2urdSQXbXq1g2D
YJrHqmr1lMMZbR6540qToN9TtqZ2L0tp+hCpEBeS4WFnCCSY7ftEkr83mae9+1v2lKejJh2TdWVY
5J+K8AfCzsOd8o367ON4dlbIR4JbfqGor59wDHM2QQIhVX6EtPblogVrtnP4phw64Oa7kfzOuyCg
7tXl9MPRjzyU9uN+cAdyKHbLOYMMs73fjMc+BywMgmE/FWOLP0xUgVJZsbW+FQHzpVmZnCyGnFzS
d5zU1JhUH8cN2QVsPnO7Kxam1nVXW0Y0nb6azKBvuiojjGOhdT49gePQwddi6Yz+SU0KI4y8Oqo4
9coTlNNST+QSGPRFiiBbx9liK6cPRFPxX38CBMZF25Xo9/kPgYnnHvetmvcbm5BTXskOTvxq4OiD
i5qOwag8RivEGm64Vb8cyHPzQfw0NDmAj9O+i+/bfcgSBnVewR6cQfAZirtG9J4nuq6FtPeilUth
rinBnlHgJQyQt9zM/eC2UWSQbIBkJ1P0zBNMuUPAcTjNizokRyPZ47yShfzR34EUoyjZWjP1Hk6A
0H59C6FJjpXa/nYDWIlc6Zf0W0BcPVRf5CrkynP8euQev0vu7ur35I2kyOb8feBR58qVFBqvTUqF
bBwIklw/rHHH1ootig3q36EoPdxHekokFJWSelBdHgN1FrsPzv/nqtezB4gDjpqb3asL9ddGSeod
6OwHFrE2ei59tYjejwUKqKHj9duikBAnoOMWGs3YKzGD92nt9NOw8lKZ84jnO8YZJxoZfSk15MRO
GVRNkIoAKm80koCbMnKMHrIGT3+uMgCRyt56bhiYcRou7jYjF54CMCh1wdUKhUoYYxLYfBVTmLW/
+EeqnTPx1zno5Yc6InYXOoen0vTU0hsGMwR71wqfmQpughZCI8CCvhVmNqOzzg8EP4RCQtya3/zB
IhG7zE4sSZCPp9w8drlWppRqOrJUc3L5VOii6brRwj+EUep42LPJoDJzyWeW41O/nzNNOUz01HI5
mjQTdu/7t8HqJ5wieaMYqSTryyn8XTmEdd/uGCN5igJ2lMKUOo1CbCcBGLXeHneZennV4nb5BMz7
ubTxWIWVTjJiC7AsILXkoMQWbL1qa5iK17FaQQaPvLOzrK3WV5seIgbG6Id8sLAfS0VDIoKhSZwY
rXd+jktd6o1YtzGEyAk41SseLJ/Im1WKVgomPhuDl9xpU5rYjyxJASgX7qZ6kD5mECR4Qx4QSlT3
LdpqSOooDIJBgRR54ONCoOuiMn2AGt68pafPMbDYMliYTxdLyuRD9sN96MVgtNvx7Xv1ppui2qjw
W7R5rVv7hf0DJQhlomQYWppAcaaAOCU1kMhsxKypyx3FIoUy3DTZvT9E9RI5+2JFQOVGlegpTGd1
ooQRtJjEmTj9t8tF7XmT2FL3UiYaVjfFMI5WA3jeWkLp/ToZj7jAZi/olwQaIMBedAc0l/qQ69/2
G7LWFaaDa8HcC34vApgfTjMxaWWYxaXAp01Y9SQbSl7ewgGi68m9N3r4C4HmuTobkEYsUv5npvyq
GX68By8+f0+wCYb7liH7577gpcrgOp6yhMoIr/VvydZ9/ANev6p8NC3IMDcer0Hv2rL0yDtE9ygV
zxtWPaTbEiDJG4Tv4d3fhlQP7hJlhYNZcpHz93Owu1x0oKcsCp3PBlVHRdC9R6FC42xYDzfDEvui
nkDZbqvWGVzPcsj9v8XxsNuwmArlvB2mkd+EP7l1JUEG6fJ7crBhgeVxCrAT2/5dYhNyN9SrSMti
r6vrM9YEH0NR10ccf6j8Jc6xW07UD5ZmdY7lzCnnDTk40t1tCkRVqrWpRhOQEjWeUP31JUzlfvtH
4oCgDTM0bvOjqms6ba0qhQe0vHwQIruOIoDHXOm3PsfOrhLpiAhBfv8AL4g157pJ81UFimykCorQ
V7fID/WKtWhOT77Bbj5hn6uzf33Qv8cxmkbWdURYLH0ewWQZacVAEcyLvQEuVvpzcdP/pJL4fMPd
z4bz/JcBFJsrEe3B03FiFwYAkEtAV/Y9/knCEJiNMYUefGGFu06CNJ4EGr7AtwI0avJWB9nzOuX0
foL12jov5PWWnWwVYxA9F8EtpkvTGecRqH89caeOVsfOepOjJKjk7ua67HMOI7C92Y5517lHFXfV
fOIuzqFOHkfzZ6pc2X0KbwIcu/WwlK2V+98qZBS4hecLD8JTRByOttL3VFi2jn6DVQRNpJZsHwgI
+yme+DWmD5PG9wIgf/hmHZEvMtQ1BYHNRyUtTYNbNJE1ePTFNhlbGE60KnantiUXVzuo44m9515A
SDEJqBO+qk8x9kStGR8F4yYI6JSDVXkgnjCaoZd9dO+FMeIqzu4JJybpCipWz7LZjyhWG8oBoWXO
lshC1vzC8QuNtPOO/KPWl7QcOAkI9n1X2vAs3CSQ/suUAz33lnEWU9eZdk8cSJe9KXHTFl4qM6s5
1jkd/Dbfnu1TM1zedEKUVGKJ/FfZNvl5+vL0kjeeUkz7/7XuGhpajVMCXcymtsmRvLHdaIjtwDya
qOLtm5RCrTUDO9RpNh5Kan2uI+1EQZ8JYQ5ST0PX5vmlM13Z/iw04v/zvPhdnSM7dmp+BE7EzGG7
3G98m78vQyaFO7PYC8NEUGaRO/YOCUMIQVNpL/XZDyRgo9YHRSZ0QEyQ60SIq92yy0EFYIiDtcIa
+NyBpdhbQ+Gqfx+P0K6hAdqWY2AzIw4DhqTcb8RLx2zFtBiO8JN7WIf6O3aFHmm5g+2L+xU/Wz4w
gD1Xyn7K+LWsrMCqNyGBhS4mCaYZyXky9XGFz83ktBCKFoJ45tuKGwZyNPtLIQYQ962lBEfaYFtP
S4rBfNQlBPuB6h/vim2WSgHZn7O7/Jvj8LK7cn50U9yI8IIgTCoBrh5pWzNQLTUp2EkLQDR6uIMu
e1lNJqAolC46oIIbFsfvZD3HsotP1zx2FEhkvFucK2vSbWiFIbz0XkfmnBEIIfnD+EMY8GT/u5AO
Rc99k8Twz6vQra6qKOWYinDuRUPxNTNppNZ60G3T27nrRMgsg8vRXIsRW2P/oMGsGaSfolMzbySF
ldblzonVVHHWJ4/im6wqptYoJ1lHZAwpk88YiWDo0Ab27H1JiFk4deHOrNSRkB00H2LFcWwIrArM
lR1JSpW2dC5fF6qi84EwZfEeSEtMyGcoeoTgvGw0vwFE2liN8NoqFxnfJ6DbWiIuvZpwa3cTsjk1
aSsbjifCNeMW5if3w7EZ1+sOCTz2QEgpFYPubSVzpl9FKFLAKQ1R8t8aS6yGaf5kGZ5r/b2uy+7z
vZZ3CdAYAg05yPkfGuxUmx8=
`pragma protect end_protected

// 
