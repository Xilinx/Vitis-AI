/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/zpj67Ydd8itZy7DZCIJV1iy0ouFbsLUJAdk7SoOY9+L2vYOXk/Fmw1e
l/921URodTiSUKKab7gocTrrV9ZM/XWPllI4/WDR3HvULRVFWaZARDohl9/sGPL3hwR0qZKlDov/
8UFvL2U5Nvq7dpd76dWbYI+LVN46hvKH4MTEigyFhBd3QVYaIKPmzXhk/ya6Lec6fxt1uSeq7Zso
xhFPvPBr4vPd+V2fpHv9vif0KpyqQwkVtEbF5wwSvSJnMBfwr/whEXiGwUIYKb1N5bhhDgPIJYPV
Ocaso1T8k2Ca7xghXtG8CDy/08heWfUrBOWkf0OJ8nARADbfQZthcN3f6+R5w6aIlpWQ+m2EauYA
P57T6rbq9sTk67PSY1F6jz+QJBPKXhz/koShurLswsaWy+TftENSWrrSHRnG6nhNpEfV8AK0rXb0
t5afRIRyBcKb/3co4LZZ6mn+HzRiAUXbq352XcYvBNr236BJkK31NEWCTF/IrkvvuAGeS4l1WPPp
ZO6U8mq7tLzAgsqTOtrm+IRfFs3DDmTUtynivI8nxGxE7nJHaJS7C4wuzeGEi0UuDuLmCXdEbFpt
Lur/2d+nLhjTTJLb/bHUZAtS9v//mKXTGWa4xK5zyAcPtpje5QekXwefT3vc131msMulCNosXr0b
wwdPOHoU61I5wFXPO6K05gboz0lg89fhtq3KoNsFtLCNmxkiwzB77qgD73mHHgf0qZQkF6yrlwRQ
NqasGtKP6IZrQ12PIMWh0GpqL6dnK4FOflDbNLHGRJvREaPe8NuoK91o8jMUzivNetOTpYB6b++Q
VtB/SMN2FesY7RAYvS57adUB9RtdzVQ3pE1PHdSpdISJscPS7socYaNzkvgOe6daEOMtkpnZaHhV
qh28QhwU2NmOCtYTzaALrQUsTjm5M3lV8oarU9OJqRTL005KTpJ3WeZJ4qPvAhOq6azf/+ajZo1m
fbJODUNcket51rUW4Xa/FnNasyNPTc8IaduldR+88pZ2SpkStyLQXfVBXer/znq3/iHnJyqrfAGB
OjlSvbgXwHH8xU5P5YtvLXtIw9obp5vKQhYJePOiyrIhZbJmoYM5Mo8CASCgwC2ZBVFysR5WBxUL
/fipPYeqYNiNxgX+Wz3/8VGeGTFjtJIxDvZdLYRghHD1La6hygl0j6WvtbnfnPSaWDjR8AIX1Zn3
vHTVwXgaYxWpT12gN07SWnSPMPQXkOiXhHihBdSzKGGCFVOjv4p0QHyoNDv0Ym2hpkV9IfDc7YIN
TnFeFpRSFqWdwbPucSzT0h2c20EaaH4fGJTqRYbr5quDga743F89x9T8dgaxCAhYMrwNYRbgnBty
6MUTEFkFxUEp/SeSFitScbvUl/a2tOJTEv3b7bjp2k4RnUREWpABKltHYCDcQW1ZqyTJN70IklvE
yjmroYvf5Ctb8zBDa0RyONPnvU2hFDx23ghNBxT3+8nm9v/3golEh2sshzC04jlppxEgrjKFAJkq
xz7bZWwuAozljrTmdmAk9nKc8LmW8tldgIXcymgB4byDmB3IwnAryIa77RXzbuctantlGX6QsqDF
R4LKNdKyCPdmjHCMSOiErKxJuftV3nnAZHI9Cvt4zUajzPuCbTh9O0K4E1BGlbXORto2t78N8Abk
9tTgdMgu/J1spOGMeSG2SzEm0VEOLadivLaT8kCEddLhYxPLNXy8MHtEZwuO6Il7mbJr6lXVLB3z
CQZD1F8ELgk6tCztksrD6MN05u8l8gxhiSdjt99JCaqUr4v+8sCKCgoqJbYn9Y6XjQZcpFlnyK/h
5+pvS+bxTRaE6uR9ayudKg+vNCJdTD873ndKOo9Sz5gLKduoUI0UAOcBaa4s2RRrZsNTJtplOt/g
m5fNq7OeZJdV30JMf7RXXIz7DsBltSGAI1kGcjE3Wfoyeaqw09yEV1BZn5NUxHqFYoxqN1WGGP0W
947TBZyJ+nsiiIeK6tMjrw4J9ybxdOWKc3RKaUWyjNn2i3JdTtb51EYg1lY+zZcM36gtt1VLbP/l
Qly/k4x8DAhoU1HHhj6RwjeecptmxaMoZy57Cn7PqDBJk7TnXo9Q6dR6gzn1YYkLUaPmDjx5E9sn
6iU0FpUflXyAgl0sD6wPWRTxLpGUguOn5L2lm3nxnjfSDdGNF9RUimt84XYpAcvFIV/SMuSTlZAR
rDLyzh6GBZKcqS0ZUuUzY7MSfTqr4iERPZvkK8VxfkXZbnlIFa1yjztMMc53NOmAuQEg6JQcK8Zl
FalHwnF4Yj3UbZJ8Uk8hJAV/Zx/OwNI3zNw+m/hpKq0uFTEZO12KZ1I0Y13ip5L+47Mj4zIoAGNa
bUnF57kYG5PvfdlS5HCGGeUND3aQ6HYEI24++x6VtZ61wEHbFU3+1IbmWwTB/0GinBHpXJM0g94F
jujqoQMUs5URYoLwna4xOEf3oS1KqymxMt61BglFfUKoNprofJOzHzgrTTFJOlrIBRugq2VxaQyE
mF45Nj0ViD7idHkwKCrOq820Hf1e1hgrD1zLBIDUXAH1xZqxi28ensh+FSAihe+hIe40Fupn/BZt
ZaoHqvcQvZPKbZHbmtWYmtFcUlP2rzgOPsxshc55BxQjLhZoCFe9L56HaX5ZJL3U6RzNiEZ3chSW
1iNaOxNiF1YFM+68S0SmWF8T+NRC8MVfXrb30TJL6iTz7VoxDjIiRCYH/CNuKnJcxxn8/Esj8ztD
9W7OQo+CAm7tYKmjJMiREgTlKqZRChRiEtSCzCYAplaand4XSxCOnJtHvw67pURcteXAT/3rGLts
MUbW+nnhuL0Iw41krywQSlw7+v+WVo7XKIqKJm3mGLeIAGnHpQ6mrpCIRJUQAOLcylcdpaonST+5
Yd1IC/qBc+npBSgsQfDgTf1COsRmwFEzVy6MXoQNOW2cJpEYu9ahP8YBNdkcODLv/fbl+TI78kLx
+7+C/MrjscXa8e4VkcR26FnxUNB1AlLS0KsNktq6cbB0b/t3fugLM/zTge1e/bv95az5fOTIIA/A
wuz4E7lfs8lf4CoNeBtYDRSm3+P0J0LiihP7fXGi0I9yZhXXolRjPqVgXxWEQcQL3poUB5TOqA/v
R6vK9PiPTnA0YepNcJqt
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
