`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43936)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT+NqHfB87+1HuXsgYQv0nkUQvLDACYxUbl0ZQX1BE6qLhTpR/2VvYV5qx1BWMGK8/AhrHGd
1rn1FQYpnRM7Cs6xtdYBqGcxtxh2ANfFdAvElxunmSoAxnQ0ilqmpLBCBoc8NBB6O7Z1vb4EOk6p
qadlGpuqAvGDHDdYn7EGOJAOWgsRi3K330KPfXvIGFhvDItu95kUJyFMA4qs63RtGQAZYZHP2o1W
RECi4RQJi1iWfRvvMpI9PvRU2GyoAnft8DY08d4mMUu1cCDYkTHg8mdNBOIZV5sDoh1Gnzw4wMpF
ioNIEsmDzkM86AnA+bZvtceuxotodxNdvgn7LeBpNEzoOOqSwshDVHkWTGMYU7XlNxNBei/gi4wQ
wGMF1tH4hiB6+EW+fQZxcyRLnSYwp4B2EGmNPAt5xr3KSijggLo/SxWVFLRW248ROMvQSiOqITjW
JoPsVjEp1K9UbUz0qN9jB4IZsYt5RFHE+jeJkNCAeUN8ntzQGBzhqaKuuVwmS02vFdPX1S2hhWoY
GC4KG3YJEW/FydF913CY1h1iYpwjPgLftKYgEZyqG+TmK3Wf8YG8jxyPFmLzRxNT3NKXJJFzVE5O
0NZejqOTaA9TcQYmXw9G7wXbIBMcY4UxJdJo5MN0WSFaReOCOlJVH65HcNRzHKd2tvwdPwh/19JD
srZi0VSu7MoJALw9ya3aRxc0QjnJdWqGBUYzi2u9LD1KxhG3H7FizXfRVPXDe5WUoDfBiVgd72n8
vSIMOxJYPxdI5p4HQi5D8hKryh1bhNJl8MpnHOt3zW58E22iA2VeU4nUyO+A0vJvFRIg7GqroLdv
VdODF7Yn2TjzmT2WS4Adl7Vkw7XVYj5IQqLzyahi4AYhALvh2MlaOHiNp8orrRLCArIttpKy8m/x
VIqrfd9EdbckW7Kj/mdlXyc248Lksf7WUSww0sjMAVtnd7P8WM1Z/ptwqQrYvSoTkhA7y+qsp+NA
emdB7z2FYLQ17BtnLcNolNy8pq3Scg7NCkMakhIOO82yr0tUAbdVM2z9Jtc97nX2oOaS6wKn0NMj
Tv2OLzJbvzNoWlasFttSHmVI0akYsu69CmGgWpu9bKNOudg03dPcDv/KYhJ9eJo8foZe8jYte1e5
1LEmZY4YkbeSFlHJg42zESZG8YrOdujONwPemUKXptTEgQLeuznx2Zwv6AljphBWt/4dKV4/9Gql
4y14rPBJNCaqzu2Nlw+UGWEn7oTovPWULQW6SoY39d8ghM0MNgq13p7HowpS9gZ+asXjj+yRZz7v
KLoiR/KC6swfiz13VfB6d64GfonP9aEKpsC4wypVi5QRAHrTFN6k4WQoO5EXSIfIbgGqPX9vFytH
JD3A6CcAE8E0KQHk9pZrMljLjH4VAfza81IeRt5zzI+1WqLOUYSK4GU6XzUir+yHiMFF89W2VrV8
muyJIRLfZ3s4W9XYPl+iQjubsTRotwpFZpwhtV8QaII6UktyXS/Qn4oUbfEgGVt6F4EHSytZ+79x
o/I0phjM4+KnTvdHhJnvPnStUZ+TiRiYE06vK/VDjKizFnGDFrz7RJgNytJmZD2ibeWy/pzrGLiP
ZJa7ak7SKgfukZZFM58f7sd0+D4v4MOsbrVcD5VOZ+grAGLwBZTBueiaNTDDB7rK7RuzSCyyLdQd
3xafduqD6Z3qDml9US//CVS85FFWMmSYJW+MtllNv+geYkQWAfFhZNwdX9eU7A21Gtoh+NP4ywVy
NabWU2aCtQeWGFmwtyPdQv/8LLYvazGZtXepOatyxniMkonOXrqljSGs2XLUOmGRmVd99eVtvDjN
RWbYNkGpq2ONEa6nwjXq3Spc3jK8RF3CchXFq7HX9gMS3nzsHgoAzo4MGsCzr8oGf3sTG9q0hb5O
9om9rX9+naTEoauyAY7ntxNrQeTi+B1DqsVZkgHezogYixc08QXKNUiREu+IZJcf1oD6Ot6fec/C
uUYqACbKuNlEm8MDo9xswxO8krpNHWmuvYrl2iHL9cGGBKldM1uVUoHqecFX2hYTXxe88AgxGg2d
rhSbBpXHm2fHNp+wq+8SyDpj6G1LbPmtRpvSw939mhK7CKoWsOKr0T7XXpdlpSaJ81PvMjKHoYRT
TwYZNN2CtLnrNUiDo+HDJ7gDDU/vHjWc2aC9DPEysOUSXDxEysI1tvL6wzaVU7afx1mtU+NtsYP0
HKWufrDO7FE1gko6nbix2/NIll1jeJMtT5fJ6lqKAzTzbNJwau0xb0knFT3x1cufNxk6MLnlDFk9
7YGvERLcxVAxHPUYgC0+3LrDCrbrtnL7GETs83dFXMskVH8Nhvmo0e//a0yNjF26zzJhXxavOeLI
9HEXsS6vbvetHdfFZp5/U8rm+VGgkbCJpr/K/IyQIzHQuNBTTwtPHuMp6ZmTtb7TeIntrn+d9KD6
rzkyJ3bqfm7AxTAD0Fzl6n07bYkDRnFrjJ8q/HkAKjQnN/xJxoAwSnVR/yrHenUJVSmFy7SPYw1c
1C4Ix0TZeuYOlpX479OdGMUMwNJudVnwekuyJt3bLBLGY7gr8Ucv3SfSwVyE6vHCe6JPvKjcDJHu
y7ks/7hXfmAEnMPjls16qt/tNnG9VNr6kE6Rx33LsU0QxBYhHJRo4uotJZTGATSXTNP2+oY37c4B
LuPsoCfkgPReSQ4XBb8kfQqRpURE1ByoMFJn6u+WERQk83EmzbLhAeDU0NYf8ZKrOxKE0G8+MgmQ
fE2gj4ykG7nZaexe7kfLE7IEmfpGUm9PgfpcH1uHtwtRX8Q+2KsFzSqdRE8eizS3etMpvRSZzNsM
692FenIWkZ/88bGkQDrTapTZyM9tSY64dLf1Y4g9N6egcCXpWG2en2tnCsIs8m+QLaQHyw9UXckg
T5mYha4aEkrSXuIHo8MSrshOTWKn6lmfIEYPJftcH+6Ue8+sG1d4ipA2luDK/IkP4vMqrKzWDLGp
NnkTWTJFImwxcywTkvuGIhydRD2rjUsC7Ur8zKL8LhArNLQjy92Q+1z4o/i0KZa9fyOaIJX/mtSG
oB3HMR05FdZ8DTDmeADHfxm0AOGkL4qJ/e9NVevnsYYf7JZR6JRqcuMpDkqzHH/iN5B5j60sEVvb
CS5rKPEHIxGflFP9lrFx0GqbZzj4lXQDD1ySJfxU+Ggy/0AViw0o1+EWUsTiiprAHnvy9kSO5Xz9
0zl8Ye50wlnUTVTmLu/ol26fu2i3VLPi78tIHUNK/Fk+UQMWZW8GLnw0aXCokT3Dcg4D/6QKd9i/
OeFmpH/NLLiTq/7+kDlJQtf3yfJBUI2STSUmffvtThxOgCncjIcMH4XDvnHqjpkyYIO53UeZK2VP
+kW8jLMM4+86m/uV/vm6qqzJiw7dkDx7zcaKFn1jN7HxrmuhxF8AwDlTsOU0xrWzKqhdP6nk6ie+
rZjInENVFRBw6XlCmG6ELel9aeAUoj16aocmlXm50k87Jf/Riccc+tCE/BYmWe3oQMnHJx/8xAg8
8x1LtjCEmceOnrwJpS0yasLobf6b4UzldmjFXolZissj+mAewzElyKX0E0wCzZzYmiePXtRF/OAn
LYR1cnao9F6hAke7QNxIDJ+7zIxk9zBEtQKWjWN8FaVkLFG72AVmdIFD9g7HY/sCr6jzgAP+sHkT
TlEOApM/FIAxBXr5YkwzGZgbfPwk9xjkp7awRyD+ezcPbmsZo3LUWZsvEohtuEnXXPQBNfPRaJWn
gqTdhvr5d/H6OGXv8ATDGDK6jXYogRQPAyniQLvVrTYq9Ct+gMBR+kjk5q7ID2/IrJgSHJvb5MF4
qRMuFohtM7Y1MI0mtpR5BW4LvBymFzCv/kIjTQajniQ1wyvUgxG0TjyIL2WQC17CdB9YlXtVbb5N
jkVVir2WGU8c9gdKmSQ0wGD02L+q/T4iSIZqnIZmo9LzfrG5gaFIMXaca6inrj1AJM8yHrJcbotk
45ajoBymO9F7VqBDnhSHkpIyl74sPdJuL1Jmf74WSr+lkVC7tpX/L8eAgSpbGbfdj0+uNeDpGHyz
I33kfgY9fkTtnNhcxK2/SEzQDOwRd1jDuivjPDpGyrOB9Hya8PV1pI3lTvl2Sujb6Jcr4qNLHYcx
jyqq7YN4Z0nVxZ3K1EJR7NCj44zdgxCokqi85QyooxVTMazsBLKxYOkDpcaJPhH5/uY15Ko4p0v1
Nuwp4DSbq+yzmGDo5EY6vtcRfiLsN281bieJ2ZQ8ux72iTwQAWjdCf9sdjQhOlgICk2Wg1UKyDQy
Ulg6IG+StyLl6MjW4JMWd9N1Wt0DFNws4q4mPeEMcGJpCifmrJgRsQ5Ecll67E7KVkMWdRspJNny
/rslR+6NIFi1jNzaDQIbxHexkezu7r48TKHOiouv/uhMrsAQQKs90HMQYW8LD1ms0HjFJpL0W6TP
wyBGNSDz6eufO/9SiYHb19AE+yzoomp3LDJHFWpiD2zRV3E32dFwtkx125TPpq7KFYi9CQU2hp+Q
NCpBF+sIun1++iWfMBljJBLAazZru/++aQ/xduxKF9Rqm61kXfytXsuS719qoCBI0h0xamMkC5nl
lZVmZS0Mk5MsTd0xktesOayvK/aLiTzF/+3b7NecxCnHWHus19IBrG+OE5ErWtWCPwhk2CyQ3NxR
QE62VpF5uC4tfiXwx0+MM8/UK4eNk9XfT40GG9cBoXUngBPHkgtLkYG23RcdrFOIROgOXTqaKXBm
7WDF6jFV2HmOI8CBE0ptQP6PGKP8F+IrbHaZWLedAaODtupN9S0/df5Wj6cwgWVYGH0XHz+TvfS/
3stwyOHzUIOYUOxLb1Ugoy9slppQNSKZxrjAnUYuBVisqv3FC8k/pyZNGxZjKYcaMFCWR4yopLXx
+5whvUBjTYMJVymwSyO4fvk41OA2DllKNGa7C266Y74f2E4ICLMoqAdURVIG3l2UhKDbL/1g4x8l
WUhRaBp/P+j4fB2vCm/ZwJkA9Egb6usjeKybp6qW6Uw7U3RGZZdfkDhHmwhRLtFVXbQOiPaC/8d0
vCj0j/rPyf/inuONgVPZNPtp6Dvkfapr9DK9wyAVT4e+JqIhdQlvXssD6wJWx9afcDpkXlhc40YG
go4w1aHrWch6XRshBpIqdPpDPi6OmqRf59q8t13KL/KvL0Q6Fg89X1OLH3BKcSiJJ5nr/r+DvhjB
pLN9s3RC2PJD2Fxek+BPAKqN70GMAmoV0QkrN7uRQNhG6zmloSkrJieke6ECSCzSe4p7msuh015t
hTZiM+ubAu8NtggX2db3tIavXs6H/Gg6XoVkkkVieQck9+iscthc52eFnxkQwiZ0BqHgjU/6Vy/B
SHcqxYyE7bIO5glYNvNrQBH21L6nwabePuclfIvwFfmQn80RNFZzfyWtvYcQvtQ87nZvlHUD8E6H
SKwmU3eAPgkYH6phJIeNGr6LscFgNnY+bwEpnA888VvDHoHUMDHxJdwKG51UnHrJcD9XhQ7qLjFi
+w/+rNg1u3c//7eRQ/B48NqFB2bB6P14RTm6HiSuju3ndZNvkhMKqyfuS0F4tY6Lv7X++8vZ/DVB
RHWVI32U7sxGN1kC1zOFMy7+ZEvHY5j950GH7lSIgf8tnEif8qxe7dcGDmLPijFvQTMN4DwQvTy3
/ACDOdKUA5f535TDptIt7R1/cp5b4Thn3C3dk2VRLessYrfjRbPHlFhWUUeEc4W0jHRSBtUockFV
mVfpGajR8bPMll/JmxpM/Utgh5Va2WwdJ3yImrG/byjeqxnGW7koWw0q6dnF6o1Tl77iqLW1ojs3
/e8ab2WB+pCURxSlzPeZmNY/X2FViGcM3PdbFhGYx/dzxhAS8IDVDzORax48k45jYtLGcMWGN+D/
Zkq2EGKUZgb7SHIN8CzaD3dAL1j2yyhDqz79qeibZxChL9G2eE3FjaKOv8HNWJHxy3jzLzXSxdpm
U6FRLmZn2qUoldBmIW1TzftDqC8dXMcB0c5EMXJHJTWuKSpqzSfMZBn/Fvv7+lDRZLnfQRrUTSGz
jVu/HyZgxSr24vhWhy7JBOh6pdx2TlP/Z7vCqzFe6ijKrgk0iwE6n0vPpGjJvbMrz6EDXsb4iybv
9u0XJIS9gAmnFJTIwBqXE+PgiLVLLD339XBJd7giL8df3SdZHkE67uTXrbB7E9M7rgCTxf66FdaV
O7uDdQHxztKoRaSmWvJPiBnZYegXHVYWr/NQC1NdJqGuC80CEpIFuuYfe7FQYw0fEYd7hRX3jvUP
fh1wD5BucQGIEvM2StdcjSbkLzQJmq88qOvRJ8Au1+/3f4bgysix9TzZfoe/TwN3d7Fsc51dIOO6
oYf354S12M3ooObjPw5iWVuFJt88KJXjz6BJ0pmzMypftwqNWNiUcjF7q7qAWiBBnVEMJOPZimXn
2Ake2Tm4hxQQvKgaUlSw7PPU5KKRnjPTZK+3Q8aVoK8QzpA+kd9VKEqsdVEWYSER23Y7YwOsUtxo
XoKyEYu5IOwwpYEr3G++JckQ7X/ozyHus8ohH65BhxG21OAE1eu7AnJbdL5pGKvm4F4B+jpk9Gvs
hBV0UMp6bxKWP3BYHuGrFaaRjvK1tb/lPXkpRoaQV0NE7I3cPggg1PLpztg+sb9OYc9+tFH1nNrc
23PKOJTIc/GqrcHh3z2hMOwXOjnpZQsEvgV0qlJOf9JQ4F5Mn4fLwN9gQdgoSL3jqKzghx0psrYo
2DP1UTp4MXRfnzVbrXcgIeIje6krjVev9SesXOxQyJfqoo2iNYtrWYOEGCZ7GXAukyjSLt52mkBu
KCl69GQnoTaWgfjktTJ7D12jGzl7ITsvdpCIr+/UNzVptLgr3OANJHe394ty9jzb4g3XBWws/gMr
70w2v82uoOHrnjL+ssLAGeJv26x0crnihFz7U3YZVNM5VCUHnheFG4MV9og4g1hPND2bka9LyNWI
IMDEao3uF0Sp0bf0TbVCqcJ4Gr3yWQyJJmMg9bjE2HujNJ9TUXE15KA81HMZBFZi0AZWF8lKcrP9
GWWTto2mJCbfjRIoeagc4epWGbZfcOJthddx8K6LPXbinyK907lXWBcAAK8TviYhCcN4VdUwTAop
Vlroiiy1HoZlKafmcEtW+txH6FPmqDovsylT2epks0MUB2LeqgrUTJl73+BEr3eaJ9itiJrcaCRj
+ChqD5VouwzAeWWpFUcNk+Bq7dsvM5E0x0SEFE2RjQpv/TKM+u10j2I7OoG6AaSo5+NSofQYRbCQ
ZLIGIGh8kgL1prnvmbDIaVROWxK9s5zQYwB/OlkWE0zHz8wlw4kL7i2fz1eFeBFh9EkU89Jyd8xj
05ahRkI3ngIpzLQsz/5WTcpd5mw62NqN2WCu9A28KjnGELVUasHz721xEtJHt97oxXjTq04UPvHU
H3x/GtoRcaksOq2TnLO06mUuUQ7/46aMPfOlCvXSTs8aqpcUw7ByktZecajdSOBJov0gH3heOSBv
nsxSYfLKzgyYnT5xsEfJ+hH7Nsbt678bngEMUBehj3xWYpK0CYdXB+q3cMwkEtYbH3FSQoqtlGVd
QQr7rpeJ3oN2X9uzXpsYy6qZOiMvChv3wsy63Qc0fVi+0miMatbNsgTrepBdTd7/PGLO/shacG3n
5MtU4yCmk17+Dccqeg6KXzluIp/woYHNQCUJWAWSgQh/NVyiTq2KZ1uvjB/SeIcEDIVKBHQrVveH
DiIEr3t1zj3AwyuUWT4Q0azrW1+J90E0sSA3lc7U0IFqJIa2kv0f4Shh/55BOOgGAF/dVzNm9zqA
0pEXioAkCC8O3Ps60JrmabKE78Pl50DJYvC5C5tuVmZBNXQhyqaaj7LfvmpV3BzJjSHc7nC14mD8
KstR0jozvcRn2MjC9vPlZ9GGK3MY0w6S7UWAK7uVvmD5B1tT9Qnf9JELHYRwL/9q/JiyPQM9Y3Ns
SDL2MdZiBmJswoQ3l+MATgBNK/iiSKIu5zfMBYCBBGj0AFtZP8VW4HBTon0oVtHco3I/DqyxnupI
+Pp5ZQfQZ2tEyhIsXyGW9KDfiFiBzmEGH6EAxSuDKp8p7FbbFS7yyq1YfrnkRpwbNPiJjBFVvVN1
O8TvgumERGqlyqKUoLBDNscujCripdpgs936Wcv0+YD7POFdIDTEoEF9DX7y7tbAArP1Kv/LaWIl
mBh2ICzMg+Ff/jeIDSZ/3he3aWDJI6BRH9OEJzDh6t20TuMqkbUhKsEFp/i+owFQAMTtpEAIROtK
erpYjM8N/Xl47WoETSP9BVoLtjKuBB2AiXaznEsusDglZ6hoElkA7xCZw5fSe7bVfjZYz7ApDauJ
37y7VuT2mNnmqPHaMD3OHQsKQDPzKxHJIeiqUT3QUTvmYzL719V/oZoUhw8eomLHRtzXlJ+j7azL
j4lDKax9/XUCdljV1Rv8sCZkPnLHNIPl2eGbsCJ+LZunWn8WzpbISEPY4GrrHmuSV4oYulM7s2o7
4RAu8gddHZO/oLArSWn2/Fk+YndlqrIvXbyjJ03bZUYiuwHBTRJsBR+pU6imroxxDe2pIQzZLack
Y26gnZHJqS6sy0ut9OOjfNruL7ibml1A/0e3GhKUbomIPmZssAzfNw8oOe7hYc7T/1aPT2weXlQK
N0xVSL8diYhPB+zZXZiOZtpEy9HL06UHW6eToXLmUdWw1h8yyaQfnB3xYYt/LzmA34bNk25n8czz
YzQH7xKYp2/uM8er0wPe3oyJaociEHO1f687oULoSJJpBJVinEfyFydl4x6iBIl5+aQHavJ1V4NP
KEIijZWbl/gywMeboZZt0Ql+A867ec0933hLfHDqiTUNTmR2l7ZZqcHjfD/zZlfZZTtjEwsBMlKa
u5dnH/R/MKp8d8h372S3jw/0nI2OZPuTooC1e0fUPE4ZtPCdX2IbW3piT/JQbg2rzLTynXYJTJlq
XBbtB/wksWPsZXDXywK2B6PB6uIvWeOfZjghSTCOHezy2pZMAB5pjIly8tHUpYqstIfrdLWVNsVm
Yn5xLOJONIHg3dFj5G32neB8jBZ33EG/mBMhQBbfK0TOVFKkMEbjEtTrqieUYBfSwRGxZcJfhDdV
FDrhLF4pEK9KC0FygQ1kJFj9pSwLBuLztGLt95RLZ4m3V9gEgi1OWkY8IR1+xoIExv9DPWawF3wu
DinTA29hmdE65t9Nvt9pc94OYU0FnRmybAFWEFlo+CyUvajOOxh4QghrVmJzAyjxm2l3CIVW3hMV
1HAc2cTmsCaTVjmvGXq0mtnJNYD0OZWIJCH650PocN60EFQAa/p3q1eoRFP8kmP0t6mkQh2koN+Y
Z8FCysD9b7V7O/Ipygr/JJ3rkB9igREvHPijWNHxW+QW8Va5q70+0cViJDGWv4YTivtNt/iiB+Fz
Wpg9gyAqEmu76q+OZQdpu6WfmwkanVIVyXn4PwhmdECzC/EES6vZ23ESwNu+Af3xyeGLjGbT9X3l
6agrf6vOsrpT9JP+yMQL8fmXYAtVPaHt9jMZNZTwFXmQpoxEHOOrMsX+/a6DFy3SSZgqtZlNHRXH
e7GTpoknTZq7D65r6qII+pKiHiBkIpId6iB2Q29ugnO1mbc3pUA4+sKDmpMYqamJcaLCcmt5OmMH
mqY4WWmp1lCav9UjCFm6xoO7dX6b/L/K+BlNmiph5M3nzOlGZXE4gl5B0m4fVA84UwxgJ7MHmsFS
CmBzdUpjkWP9tsexqJO5gfPbWyCY3TpongMGsiiIw2UD8igcU+wKeuBa5WF6IRds6emycMX6X+Ks
T/1pp6W55N1AwTknTgzmpvkJffvh5ODzO/J/d2b3VoB6wYKOndT3C3OTQppOhWPdHnz4QoJYQAna
VhP8oStx7cKSAQkQYWW1ZkVJE/ZmxtXUbcI7jyXYhtpQF0Op/Yahj42OOH/plIFW0/gchai69YfG
iSnU91+beVuhhAoXl+vewKbsreAJhF9wbODQbfnBxOkjUU7QB72E3GvYTfyNu9X4PFYs87BgpIqz
cGJn4HR8fUDrsuFg6ydxbdzW4QlcgtogkGquglwluz6xcoals5u5oLig4tN+H1tjLLswVGUSrLA3
zXhBEI+o5+c/xUGW6DK3VzQShc+DoeptaqVXbtkFSmULG3JtKCXWjVYPEV6r6F1mtffuMLOajIiN
cmzisgbgQt2s5+ecvyzts+3MIiFOhHMrAOKLLngHcS7TXlPfg+F5Rty5d5PuMSevRaJFGOK/43Ly
FGV1PNQohbIvJxV/jkZcBCBRtoWcU0uvt4/D+y9F/sjj2nQmWmanN1YLK/M5wOunX3fztF2EBYqI
swKDTxmOwx+ZPKESh3vvtNsl7CcLhvpb3nVRsBey8r7NLq2Npbqhoj0bSLV9Xg98HWQQn6XRLLUi
ZIo4sSLIOCRqN3HBE7CP5VJu0IzaZmP7zs20DETWKzbRaHcz/SBj/T/Wy1Kl4N51RjKxnHXmQ/mm
vsYjrj8c+5OLk2LhLqNlCvzowuvsOwCufVZgXFK2f7bO+jzxCBZj9hYNB5F48GEoJhAgUU0edFsx
4ivyOYQtPj2eRI+bXFKyfVRnNyDpFa8cjUYAu8aPT8H+RGKHr4fIL2gyWUKjT+q+pn4WrjPj1hab
rkkJjENhz0C9ap9XaOkczf/1uhiLlK64mF3pc/zjkRxXaoXZ5sb3Uxz4sStD2umft49alxiyQj/F
9lBmvRj1l6xp4TMKhEopskOMYZi5w9qRk2zCO3CpgaCfrLU8r22l6surdl2D9nEzL7gYNJcPrNx0
sTvQp3BYSL3CuR8TPqfjFBil39kVnxnybWUxjWBVdOVROEmfWZ1gzhP16Hfx1PLWME5ESt1J11PO
Q6oeGakWMVkBAiQPZvHWdgucD9v93czaUnfvOvtxqP7bziekmVNmli6azgHFQBHF7hNKLz/eZCbk
ztHZv9L8crQw1kjGh0sm0z/5CNC5sT7K4NNcO5WNFVP1AdIMIRyZcMcaPKbzSwjb4rxRydiOjHod
t6WaqdTzXL7INTj7D2dhSi86bq6UaEZ5oXvYgh+CHpwJVHt21XEnV5FmBiYQtmnARuyxmM4x2AQA
L0MTBJTQYSjE0E8RczPakurXYMKkucY2qJwqdW1zNk3OGrjQsGkT8L7fSymUY2FwmZt6BD3xWJDr
MdYbaQk39vrYxU4piQ0zGwKPegbf8XY4XiZB+q1VAkZWehrEt3umLuTD6BI0Mc/r2GbdVCwoktkh
HiKXP1lWaimwP7HMv3Es3RAGGsHRnDuO2zvo8HY3LKt2NaYAky9UmRtjdz3T7H7quzkaMHBxCg7c
QyGtj6ch8dG0yyXuGYigkko7zar20HUIz4KEjc4gLcxmZ3mnHB6EOUJPOHPTFyQMatJfP4+0tCxz
RLa9/vVio+1y+m4QhyjBNOKl04j8KKZ+wi+unaX+aBIHurPC7oUI5ABYUR8O31rnmFXZO50/ZvTe
WA2TJYlM61d15olaZM1ViGapyxxIt7RS7gcPrExRk3/TLAZ4x/THbbFtAaAPIOzdFtY217GIqUT4
8h6GVAD9xIBWskHyKlkmkrhtvUWTMfwk75YBw+xK7QtJnHxG9RkzMYmc0knLtVJ20AW/yHyqNJc9
TVkA7eg2RKZtgsT0N/dlR8RCXqksvqjlMz8GGzSTfitCKjntC+l1nOcUMkzuVlGGUlPQLiMhlNpB
0v4G4RimWmMWhJns3NDRO4ccitQybJ5lR4VW2+hy/XLmj8mDutotkM4gTcipkwaqmrH9r5sqGba5
IU8BlvFB2/M0apyN7OP1lRJ6zGfYWYSxUKYe3ob6Qk+nX/iIDM53KcxGwxRcne9vw8lWYKqDCSdn
tqbt0DG0raGAvlxM5hhpGFtcTkmAjL1D9qXeaZWH+wkAxeyuxbQ0flyn9rlXb+rhUt3Nq5I5JUFc
NvdpyLCLWEPIFFJMsb6bNN6gFWQHWpr0EaaLqV9969GOQwfYFGS1HD1M+ikHtTmqqz4ZK0sTa4+Z
8KIF1XjmOQOje1hV2om6eNPv4PXbZPVbwIvY99CVTr6AqmTUr/KdxWpJBG9cC3hm9a7hakPZi2nU
S5uIReTBNwRNz7ZAZZ7k9vTEQi2RT6zAL1T6nKE/hfY7uK8ajLMbp1B0oNWCCAiDA4wk6KZ32bkM
DgtVoAt9uizjGPj9wHjUWQbKBJc8eF7YDMT18r5v9mJpyL+E0BsIjftoA8BEN1EQ+I4unYrBwf+g
vi+vbqf/3aDjH/m4MGx8VRmAd9bFSTlKSde0OzfmZxtynN65IEKZMa1c+D4kd1Hr9ALQCzDlksSx
ss8k0ynpwtKPoEmZMo4NczbrDlVCoy9D4xt4T05PMEaBOckfM4Q5izhEx6mRQ1C57ApaCzX4GpSN
VyjJtQIe7GihRsggmZmO6AHYPJq5aiqRXqFEmZjt7z1k6zFDJVY3d+DFUzUTMXOxA78g8K5eTy06
D1Js4DxJVC6TCgLA/ljfBJIZrox05EIJs+17qV+GJraTbOHU/XhZ2lpslkkIev0ocO1KWXRDsQkC
xjc9NC1eg8T5RAMRC7YRNd+nTsqYnojcwLptrwJ7mk9PRuYwjjiD/mvkZQZXtDukmSVkwAtnt4Qv
Tro5IsU0oAQXkQdMJc1u0JfXvBQ4ixjATO948Y2gn/fb4Z04FgrySu9AnEAWyVCy3U84hT6a83FH
ZQh084VAC5eKE+nrxt66P91Z8poH/aYkdwDVxCbNs1pN+dhiRwO5YWCL3AgVT/2OXZSjxbKwzeq/
t2zqo6vReoZH3PzED5SzNTApwv7eQcDeqwllqnEvao0V+j37ch0mORX42geWKxuEOMYg5fE6nwDq
EInHqQhvFyB+7jZSPTzsM2kmn9v4NAi7IVvKsqtcSOQpvL/Wr5q9UaWKLj2uCQlBBHznHYo91FNf
vRk2LVXE+jtkutl8tInIofmfyjmFqec8s/BZ/+od2jbWVB1vLoYsLVdnZs814Y/NxgAXxnX9kcFc
nlqCLcowW9CxeQU1kY9xc4/oqTkpmdqVUDDORJOio2MPrgisd/hyBHrqSB6uw0DIbJ+au6c7uROo
kf+sB0ziVZema1RluSqL1gv1VPFbgRrQCA2JWVFjNLklONPemOUzH6lebUs64Hd460aP82axPjl1
HlUS6TQ3irgbY1UgpReO39RlsMASOFFNGuHL122BHelFQG2HPOTPKRkvd9yVjlFePYTMsJ8IM3ov
9UF3w1wGta2Ma229n6SiY/u2CC4PvLih3No6bFfgxQZPj013Kh1WVu1h3QUpcQoniE+8iwY/Wu9F
LFZMLXwF2b2dWmOSlLyKD5FMCva60iasu3GO7TmmHj46aqby/ufXpwRdY6r/OSs+OwxF6rj+VYD2
qmCvtYhB3Us8UbXpnI6hrzdx4QPx/tu9RZTQAD/nYnspV2BW3kdUm5K3+QdfgrSzVHh7tnt0Jh/E
Y3RAjcCkbPOGtzHL7c00/4m0Y8yVBYWbYZ1lStgyEkwe1GyXA9+KgOCSbhL7QCUZfbwWtkjh82/e
Y320iyi1lfTLsRj3JxYps9r5Kb1rXLSMFooEqaDdHLaw9pBX+c2Rkja5IbV5keElbZHLsIL1mmSd
tucYJ0CFDZfFKsbe6CP0/stjok3e/gtvyGlNQfkk97YEOrA+VBueQk0wLlFaiC1kFfHHL+jogGmk
sE8rBNHmrD/uLGx1Q11IW//8JGlbAayCciu7m1onfG+h/J4l5Z6TRcAutgf50Wa74+UIeY3VL6CK
w0sOfnhuyDGf6WOLLm3ckkgww9WDzq883CXSnGH8zCS18bm1SLgQZ+os4KGCNZDLkSc5wykAER+L
ROh82hg9T3f3Gm0B01RRt8pBCI4jKT91aIJTrLM78zuZjq5KSF76RWOUVPXRDJ1hwv3zTpfepriM
cONqoRAKbjBB7ezhS6oizha5ouc0YOBLr1WaazH+YLEXUR+nkNBEPI9bs++6gUOFH7Rh8Him5HZ5
ZTjGzazPMkm7WMn6Pw8RUrvEX0+enx3ap5vUBUWDfdiLM5TWQvr5rWMT3Wn9V3IxYHAiQ7M5cVRm
T9DIGdus2DegxJWMCeWzj/D7gD6NFANbz1urVDgBGtck1TJt/UtKy2A7cgfZUv6JRt+28sUsbMwH
HvKjhMiWyEI3dtxuwUD6mQXFFhjKGnvidy/lYqWoOyy51jvWRATovhjwDnUC+xb2T9dfsdrd3v4x
UOWBeibwi6jtBrjNE7Ig28H/OrLdZFeN0vEL8Nf3/KW2Gwb5rQ75xyS1vAX9O9teNuqsTxENB54c
BEyfKRs6BfWn+SokK5DaAY5sk9jMwARK+0CLvCLIQ7kwNtPTRQX5uzeX+fQQJHNZsLj15Yk+CsB2
hj8MAx8u++MwblTDWooWdaZW4jc5A1T06vh/+e5Mzpd9s6/cS+2bPKZ7Sm9oKzyepOLbpgAqy+nU
laJT4N1pxDR+8IRESxjNx4IAWfbu5z+uIkBmTF6aINDd5fiDgaXN3eJx+IivZsR9eezBzTbR8YYN
GEMiTgpiO8B/IbU/xnqRZL3g87GPtHjUQhEJtM5egDHLaZqKqPIeLUxOC+VAxTbLu1UOH23gjpNv
q776KCNu6zjcaa7g0slFrkSQ8qzsxCP4sg+P/Xu/yg0Ei5MW27ijMTPsXj7DHIPNdASAg5X+OVLT
GIy/lPJj4xgiy4HpwztRLZVtAHo6kfBLc2qGCFhWYdZyWIIBfiy+fAYnEnFN0eiWTqU685ucndg8
JlX2tDuZGwPviu4wn8Q4oo5fbydBkSjSq7xoSJ3jaaPUcw1wW5WvtyGEqj6lAX/XQfSfOLUx34rI
31Edx7Cjmukr1Tel28eAaKeS1PS2rv8jbmTF96Af/TEXutMHUJbvWVDJ2Jp9I3hv/+BVP4seM+/4
BU8LbhsjO8SagZjqgeQfqisNVlCM5gMXFZhtV24cf+gxvs8IFxEi57K/sSikgwcwNfwrAJjP97D/
PedBoGiIitUr+cSeHEcVtwEsiB2C+LlJwHCTFpQ+OuLnn+79n0LsRa7Hdpn0qNUqE6S7Z9UPEALV
pbGeQwsjrQKo8Pj1YvrMCzLVD9YoE3YY4/qv2NCTi+mg6T8QeoC8kL6Ibmj3/lBoo9dFg9Bu2dyT
5o9f/hPAMOFN5vRA1RCl3y5NGp0rGiUIgD+/KHMQJ0G0Vj4LPRe6qSi2CwA4DvTXFjsje1xfAxyE
p9Vs5y1QhRMfISCAjX5btvSxG9OmnTDOlas7ZyehE+u4taHliAQcLbTjWj//Idw2a7VPWzgg63rZ
yzVLaCWc2qhZnez79hnpAsd5jl6sofdwUyT4zKiahQ45/hj8TSZumqbO5PaTj5h/X+1P35ujMqSI
9M+fvxB4tlXYH+TFLrMxTZ4pmuwCa5828v5Gm/lxiMj+P820JrimoGQQpZlA8A/gUjFCZrIp0i3q
byI3px2FROWnHl3xZBzncJve58xfI9tOqaI1b5Gpo7nkw1M6UL2z4mdj1kbYTGQ1Sr/JskrmT8tF
MUcUjJgrjKWr3tEMPqCSrVp21ZVG5Qhda20Qr8HF0aMIgQobizrISekJJiHNMDpxM4yj0nHCcaJ6
7fK0HDRJQh4TcWBKB6Gtg/h8fOtlw3QW0L7wfZNzR6TuoSREBkM9Ltw7lUQZUT6lLPNXzh2W5Ms5
MOQFYCQ4/dPuJbz5n4gzYLu0x/FzPX2cCrjmqf8pD3b1cxUl2oagLclGWxa+rg8MuaKe175X0isB
+mDD5b9bt6jSGFFd5Yu5ZUL9ODCx0acEmxR0qZlzfTgIHhQQYKDZDAy7qjIHWXd5LCAyDCuwML7c
6Jjk8HZFcPQud6c/oYRDkiPlQBwt9Lo3KiPtnCsDXgHxXFOBS/SczUNE4zvGEfMGN4BJe0Vu2zwM
txqM5RJnZNvJR/jqMia+Ju4mQohx1SNB5eFoQqwT0BYBwiQ6ftzzragzDEbkWtp5NzpL1t9NFiyu
7FFTrmXpxULNcMipJQL/Z24agwsD8KM5AbahOLEqrcDveKnOI3NeiY2GWsHaD8JE3MqC6yz5j9hT
0xn42KlR5dnV6pVr7NwokpMo4BNjtmsT9JJC0D8TKpvbBaA2XBJ8AVK0oEhTU6fXnbxgv9r1YLUO
34yDlpuswnqlO2FCtN+su2R7oWzg9Tgop2oZX//a+kIK1podF+y0QKahrw1RAme9i79FdQF/YFou
0DhkDI5aXWbb1DuD2sl67KS912ha2sIFFLg6bER7zRA8ExmW+5FNhi1wwPUefQlmA7Z3dfzETAWL
dPGwVexer553nQJnJHnIZtul8ztTIIcUA76vHdIg2c7s4T5JFmQX9HCu32qgk8IfuUdDg7zZhrdn
B62PUftHfWvebuDvMEQiECQq3FKUanCOSqW/R6b5YMBINnK0NkVc+WdJl2sgxqFHU/YC4Bxf7IZ/
T2OuTQ+p9H7nFzeApHRcj/aR8UKsFSBySJwXFFMWzuU3tSeNNus1jzrFveI3BlbU7QAwMh4tRGJZ
LHa6c1+dESLhAvxYdiz6bxoDxBpb4CTZmFxKnQfD38hwr/DbZ9+j4ovJLyKDKGus7y2E9NN0seQ9
P99P/tv90GVGwH4znV3hflNWSLxHUFFylGbvFEAAXJ47PPu2HtfBbt4Iv/v5PgyxT7T6EiVVMVIM
4tzEnGCJV1mLkpg4ZJ+kioV6eEKn1YNm4Wn1C7yjLocnoyr5p3g4d4CiolvCjmpCoPczUOobt1Kx
ZUoLECEC4My1bJbOhP/9tKtanDxduwhv9luE1BB3U+fP6+c6jkn8Z5a72HVd3DL1IKzUWLY67oXW
Q4FCq1g2uhgvAnnl3qd97ngLKXfvpFTbWOGCYfxoZ8M2y/id8r2arMJP6t5YMfgv86iQIGuT+lTQ
X1uTtOE4Xta0ObarYE8/KpJSXDHD+bbKkahj55OZUL+3A3TfJ7psOgW7H62DfgSXIiqPURuCR3rG
Nbv8Eu4XKllyMutDDeqJEjlPIx25WYkftkZTx7vziQagQK6yDxcDAILpaIq7njMkbBaPMhbUGHG/
/+hxdeTrGA0ipSv6Fl+A/jM78d4pTFIG1FaWdg5hTnN+tpOyJ2YKKFsz2Kk6FgxgJi5igzMtWYyX
qvJ310i1QEoLe1oTrJeaanIDI3E52trMrKGoSbW2btWYed6PUMQg3vgpER/3ivnmcT/VX01q6Mpg
1ikNw51NRrOJnGX4RZIvLep3Z1aZxhLyxYgqxO+dM3SphM7p8VHkRQExaKJFAjvoXesHeVs6/RWv
gaIHYQV4bXppRNfuzVOCOSZJCISIf1GFKwUk4W+oNcp4A9TY97fM0MoiRvyz9ASQyIMaw5WRoLyF
Z6q0udDhrGb0ciSkdCN1DRCwZzH2pCtjr+MnUEOnYAsagZZx3/fxDoFfXZBiV6ee1oeCaf3vUMHr
ABqCGhFaMjPQe7pAAym9Ic/OLoFNzCSGAnpuYM6mU67DeXniBe6ZuUmBo6Js0kGyOOCBHLn7uwKW
RDxd+u6VPvW1l1vgdGpxgM+IV46f/L8nMIbZl+mEc235q15NmQCI6VcF7ObG89pBNY1Md8OgjRqR
1D6p6Se7tju9XtG81CIavEY7uQbBrvnmefipetUUy0hPPQd2rv3d1F/eMy4g9x7k9Bo2kB3ED7fO
MSlLElWypSNKNzC0agERszR/BIZylt1ajgZfPHGHlcW57as8cVkZIHjf9iDC6/uHElTPrPlJfwb6
XLWms3e5+R9w7WBIke8sJJ1k6BztPMUv/Ptszw8Lv1vmBMaamgnwueBEgwnGiVLwDNz2Gh/Ghizq
MCFddmwnkmohoxKz+H2t91rOdLoZx1rsdhjdSu9OAV/BmHoaL+ZG7nTolC71rtrzWXp/SLn3f9MN
EK8UuRjynl/n0m7hEOmhHQpim08FRvUZ5o5bnqdVFjbZUoW+yoxUCVZluiDSPlpoZY3u9POQ14c/
M6+hYhjwSbLzzT6u4TlAoOL3MPr1EMfaGLkc+7hMDJGPKAS776XSqBiiHmNZQkYsVnbi4mEwrRtB
Jqs12/IMFUPNPhKaS3MgSxh7h59KjMq+iDgFaQN+2EyBn5gT/p2Ihk4eXTuT8iKRK/cSb5ilxP5A
0cnEXsyIdAZ1CYpfAZRkWWhT+5iD+Gb/bav0RkezZMbUrgHx9VjzN6tvnO5WM7Q4W1t2U3+UVc66
L2ZkfdhTuZlkTRLPv0H9RLu7hjFHzV8p2HsUiJjHF3QjOjtC3mG3MD4/3cUdBd/jVvzeu7b84k75
YnoPyYco2CISjrPacP9SGVoqRouMthqfCPVDIHdeVavJ170idWxGA11u6LC6mleMn0uK8bnBEmkc
RziBtSe/ureCdzv5F/SqpBDRTuoaApqVrMVGHOv3iiCeN4Dx1pkMbJmc1L9PE38QL3p/e32COFvQ
/KlskyOsYrSTFqSYtdWNerwU0yhCURLUIt4eXfqcs+1dYUyHifs3epbhtUFUH7UgQFa5IrfVrl45
uEiPcBjSjDK01qVPpCHwx8htdAHxC+uT8CzX9u0kIVHj7rNTru8jpcvQ0x2hfOjaxKd/pnAAQsld
2BI0e1qJX30zOb4xiP/WdWcX3mbeBrtZxTApyAkCyQvL111+ObR9tPpBG59bGzAr8rNyTW+gThaG
yUtRYrUGTgWHNw0MQ6E7/IOHtyC8jpYyBWgHh5ZAFu8GxL7mZbrX0gJj5h+7p+IteoK5HpcoqJGm
rHW86LNmZbCB36yVjziGbyEujCYG0HQOv/9dkLi3qinOojnz/eBz2TQOOZ2ESxMPKYZXstgsfJfN
sMH+yxB4GIGInphNa/UqiyyDYEbEwGnLpQn3l3mWcaWLrOfVaHK/+gO6D3DUmneZNRZ6klr2t9pT
LYZOVuROvut2+mSs0X9UhTzGkn0Y1sCykujnvv40sNptXtWce4o17TCPxcDPA56AGWkxTY9/Y+am
ZiTO4kIfgHeWze9wUyuMsyxR+nf6zYDvABj2wLzOTfEMIy37jxSdb7I3EThavfjfPFQJBhUmzT0T
h1LjafTCin84xoAw87mmfHMwT3LhpAq+xht9bs03g+bc9MuYQc6suxjcG7I7+nAeWiios0VjaG3n
2OBiHoy6EcnzNWaUCRbZdhNirqQGpV5+rTdkf7wCgtbvkBoGaRSTVyqP0MtZ6ABaN2lRwTKZU0G6
88G4UurXIvUHxRwCRW71Qo6FcfZbhKBS9fohPi9QtzhWmRDAD+fPRBgr5GEnU3z6oDdbAp5zj/oX
rhTDnAYdhzU19t5NxnP0hgO6Qc+xr8PK2vu+q5dGxzJpLQNXIWcV6jI0wpAWsw8YW/3/Hvgq5RiP
8dWIn/cGyDFXuKLr+mnqqAAaB+MZpFgYNNk0L9qAbW6hzar28/fG0yoWv5zF+vskTkf82thhnnEb
2rDgNpRVQVhhOh26dhabRyxr3SOyfXK/kLEQtX7LA6Kzx163MvfqU3Qh9zjD1Yw17jkFijnSlTaV
NdH5OwpbXj3nBIQxXRXh6ZndXrQdTMqN8kf9vOC4p41mjs3XgWn6VHrYMXzAMvijeynuS2aApLIv
J68izn2Ccw4e7gbZgV3URTSU1r3oThH94rYKYo3bk8KZigycP5krwltCBvYgdwvsVnxR0xN/+S0l
+V9kWOCz4+xQJ2PJW2A9Lt+1NtyB4UkDa1CN3/H3Xv+mJhM0ff3KR4oWDB6rXRYJZRZUBSM03nvi
2FbkMBoGe6kBw+kHu2WKZDFrRUATaV70c4Mz2PM/xwv2Ub7ihEJWkWyjyuH7iUdv5Yk2UgSKXCUF
1j9q+9Wq2/7wB3oPQBosqxP6rnV94AGLGLCKR/wT39aO+AO3gA7caQkwR2QQcRcahidLcEm2xILj
+W7qEBinnedJ1L8w2g4f9JZi7om5QV6Advk82l0NMRwLEcy9veMJMyov9YkFHdaGPP6Z6MuTIfnQ
Ap6IGB0HyPpDCJTnAzytPXAiew/VKFzlg1KA9UTudLu+U9/vkNqwMFmWgjrRgpFmRWpBB3O+ZOqp
5AR07xT13HaK67DaR1/t2LRykjWWB70JEhsIK3i6VwRDigjFBvSFQ0mDkUBaft5WWCKkGnbbxGY/
JNGHNYYzylmTVq2rca2100Fr4Qf50hvmx6b9bBO/KJs1/1b94dOUSkDPCR3Po35L1I7WqtvXvh+V
nx1OG2P0+GwOXggnLEOKxkN2ksrCxTjc4dhEgw+BUaKUPYwMGly09AWkPKk7HCHDPGRRJ9CgOJ3Z
SoPnwykjcDBr4l39242/8YOqGKGvNBa8E/jirJwIRxdi0tmYUj7ojMh8atXAAYn3Q1NfMwmEzkE8
EPDBQR9yCFPY7RbszMEnr2057fPIldtSs9XYEr8XFHK/58rb1FAQAvhod/YB8U/PTc+fP+K/+7vY
ZP5+WVq23EmtLeD3Hzv0QPh04Bb58dGNz1DPXOz+xD3tC9Hc01MupyLyu7xH3BaysLPZnN5zW+7m
292yA0yQcn+E0OYO0uf4wkP+dD2B7q5QKbtf03b+Buh5bDqSKLFA8TXTDmDiUh1oMRmFPLm+RAAV
zKIA3y1Q1MpDFQessW5Vi38T1l54/fRVCY8UVs2TJ4s8MjTLG7c690FXQNtp68LVcYga9EwmQDe1
+neLMVblv/Z2skEOzPIaDSkp1nHaRu5ZtyhLB0EeWCf+k7b+StflvN+98HD4yp4DLeaQOUQK4T0J
lIyIUbIvasznlyNNA74Sf1TGypcGXyPqmdePGWQCX4BohyiQHPoRClwzy1N6miwDhbFF3ybyCQv5
+tQI04D82ohnoX7DgrkFsiQ8ek4hy7eE2fzDlbZIObJlRFMsIRO9cRbNsxHL1ww2f98Rx0sADsKN
Dj061BjO+1XHIucWk9QcjYNODnB42EiEgeVS9OfbA7r5CGjff74D736Y+G6/2K8C2NuujP5g6JPw
LXVdBB20/9qaje8GdJ+DbfpIgzgGn5HwJdCKp7bJMDAYprqqGQJkVZWwZBTIGp8/hWO2YECySki/
4bW1zRWzKa7ZKeNyWRrLboTtmRQ3EKIGcYVip7SSCkRKJ2Xf0S6It3OJdNOa75CP36D6QdulHI4u
s/GY0uz+uTIFSPCq9Nd2B4fDdWjkqMGK09arG7CgM9Pm/sGYrx1TDqjSoqHF8nM+25yg2wzWAz8h
9T2g071lIvHrCjgjZ6xWF6Z9AJwPEzRgrmeuSGodguGapdOvBELpQ4/9PpQn1mnNbxLA/MFlaxhl
RqIxWa8kQvWUY+VEtoJImY5rCv/QrsS04iSbgdyYtPSoHrSiGqlZDuyWZTqsbxzDWGkslOKh4xI+
3wnQJBYD11Xz3oci70L8pLySb7Hvo7Ziltejyb3/w7GONiCyx9C50wkMJwjxvSoQO4RiaqbKJUmf
D4Pr01NmbSukanVCGQJFvQnfloW9Eb9ReOdzA7QhiF/OYj4szzA1uSKErfI1voigwKYyheCbZmNg
733nkN6AE9hHp7RTiREQ4KG7qyn8R3PU/rRFY2gAjv40EGVDWQSQwIWEy1zVVxp4OsV18JSWJnlQ
ufDVyn+Y9DdaoGDYvpluyANGbhlj+2aNjGv/ZzJih5O8LY2LXQo/UXX72bNyutwRoe8HZmmgsNvO
zhDmyoc8BltV3mmn1/37+X7rbwo4gU6wH+3axTOOCGwxRxl9YibqWaTgZwObbeVpEwTRQ+weZ8fA
YeOHO8X/NyXxqiYT1dy2GORUL0TM2p5jd4GXPMjqg/5dd4ooiMwSZ/HpQzqWJQo4vUdPhYICC5Yu
Hs/PprMEne+uO+ZFsnn9tykPlcsbwGlnawv3/VDFsG9nxcSHbKc7AYXZi40MO6QD6qAyb9OvIdg3
d8XN+ypWMxyr9SxmTL17DZg2vSCGGDTt+UF9jqucL13wD82ymEERYnBxaTN68tusgpsg6zCgNZJE
183E2qzz4V/pUtyQI5oH9LckrqT6EFRyvbJdLvmlZv2aOZNpWUk2fhjozm8WqO/rSKTpOcuUib19
gINaZWzIA1wMWYTLES4GJ2ThVllgrwW4gwoTQEH2X2uWlidX5Ild6fv0bggJHljxSb+1ADRyM3LL
coE+NZCtIjYJ5QHR2jcsbkx1eiv6Pp4j5qZHeOBeBEWJNpVNJ/EZ5BRiR1X9Kpf2QE3zBsg+m/WZ
D27104Pm+SQ/ln9i3Rm3kagzVRSlkhOs6lVnmc70Z1qKHGt3Uo1KsPk1H5hvLodxrot7OsotGAH0
Akbf8ibM30alJSJbBDhJNkP8+MNrCG/YmWdw8SSUdZbJhMa9IMunkiP1LwZcc+kPjJDH0fR62dBM
JbZUDwm4cY2Z56d6BUvGSPWiPAM0y9/pgGLTsWsnmv22vc1fvLyivXY6KS8/TImgZHt4SPgEYJ3l
WMQrJ5zAhaoUeoPhF4R/8Jz9b5lTbebIG/vt/ZnTsIFsC2nDl9K2Q+d4SBou4R7g/OVy3SwF5G35
KVrHxoAvKUjTjwHZC4G2Cns3qpIXuy2uLAsBmvQt9I75Cvd5lC7fknCMQtWktqh1uVZzDx7nv/mj
CyTTlBfOZoP1XCZjjY8Z3Garv3jJQ8QXNJ9y5vsCbOfFA0zDe9XZ2kVmvZonaq7+YMA5AwYcxO3c
uMNBD47pcY9nzmfGjNtKlibDmjZvS/HYe7nVYZWZZXomv4yv+a+h4wZlmim9fS1yOHQ8NIKutHuP
Cw1sTHYTFTfmREn6DDgk5toEhqT0OJtkPJBlbFGCxd5pW9w/mUisufGOb8lbo9Q0yAu17bt7XxCz
gPTT48EUc+WwE6bomadHRfdpUmFyjuoZ6hXJxaTE+nPRQKcji3AbagUOjrVCxnETrMAtbFY6Bf7y
JMuHqWe5e8b2HR5w7FLlr8sOmIm3beC3bniLvtRT9XnyrsbulKadjarP90eWPw8YMMJcEvVnSvE9
HjgFcm6kd2XaUZpjYVwH1ZKT0vKUwvNQUWH/4vLNeshLZEuxHnZHtPdsDgBNHf9cPEFbHpis3I6c
NWy6FGPctoqR4aKGMUFiQGm/5Oc8r8NJq+l7ksN5im5BpLX9QAvdNNJ0bzmhIyQxSz0laSvaRNJB
hy17lNrmFimbm9V15r69Yzq7Sn5LwbNDTShHBuVXZf/ZfRYAqTW+QyM17ZS6M/gfg6LPBRfbDGYP
QHDpN7beankDWzxaM/CNPJs4ZUBR2jhDkVEyeerZksHYMOSbBjP3m2c8tlbtNnrEww4FFHlaaacf
aVXPmxwutf1Lm/W+zVtRsTpj8iv+QDGqkbe4p4pxS7UWCveRwTX6aBkksZ0xmsKuWaTVy5CdsKmM
6m9j5umDJ6EG3yV2wpNiVXQY0lhDcYuBRrbwO6r3zj2yneqeUv8vRHMDnKlx3ve1mE2c8yckFwkQ
2WccXFJmuly5DLycQptjk+Mbw0WkbFkJJ4S0xV35avy9DuAspQ+e37FfZrH47KsYDZF+vuvtI1Md
JVKnLoLStjxIe7upS7w4sG1dZv6uqf66zKMVoKnSFyholLcVNapmYls0QrCe7iy8YJm8ILm1U796
g+E9WK17gx6t4lrZ1hTvyDv70T2Po//bGrvXJBX4c6uMMR18WQAtEJp9j6O3rpmF049p1XdOkG2p
CYsUO2K2ESR07JFNWFBBdQY9s9X7ySAHgxQD9lAHWBLe7yWSvtQZp7OZksYOj6dSPehou/7vFmA1
2GOBMuDYsNgKtZ1OpTbnVZq6pTB7GieLa1TSfkyyCt94ltaKyv7XUyWrsZoF2FZaMsubeNfFK/Os
0n2uzZhyMvnOwYMMI51zpfZDbm0DNRidkXnaroO122YuK87aMcra1jJT+JcrLWNFaAihmse7imfJ
626TV5QmdBeI0cZ2sfBo+EB0hk/9tMmMtdO3Tv6sCmAPwr4Qx2CWx9AD+LudNZsssYXbuLJBza9L
8igqHF1EkP5jv+qj8Ckexy7FwlYRetmzFLo3hPN721tzULFnn9CDNV0dLn5XuUv11shfLyuEPFgv
rdTdMRpOQf0v5ynPTot6Nz8+w/gFsByvSJtkg1spbf1XYYgeSHxRqEUCq0VV2ACuhunadSuseM2w
ScK0/ewZQSMV7i5/tshhOvFv9oEKVJQU7EmN285XTVwV3dZMhKBwVs3dA73YLU37kOzZEuQU6dpJ
rY2zqxxYWuQMKL5vV3Ed8tkYieLERoObq5Ak8Bwc369BUtKmqYOkoCZcmq10TZH7kmXJ/ps7H1v7
HTKIm9FMwLQ+MPZvvlNd+JZJ9wWKSdpHSUsURPMwKi43QuFLFQR869ExE5MDiMj6BLLKxe1AG0Cn
gtKxvLuHI//U0g0YhJ9r6FKW9DUunAbXMdIzNdCVXPoeBrCpafUZMtEtTcHxTNejOA0gKZnteNuE
pZ2D/AEpWFtKR3UqQxVe5AsoBbx+GAgtyo/5DLeKD8dYqIAuUWtzlSWtQcO+skRqsXXWUrKKKmgQ
Gz6WUqfOAEwsHqYgpUuzdM009YmQeCX9oiSMAmBcjAcrYqX7CJi5NidTvA8liB3ID6sC9MpdtZmt
hTH2OEpAcAQ2xwrwpOjJpQG6200KNg67zQjAIptdTY73pTi6GSPr9hdUs90pbi/T6WT9zjh7FarM
xFRcNgAs5f4mo2rJS146ChphndXF5UHwQfUrwo8PuMVEZuJUf38ok5fn4urIBnCJZ2WjtNlRi3qf
nXO2ZuLCYqR9kT835Ui+EB9lCu9VkG3HuSdzg+FYBMcVJl605B1j9FueB6M7LR8v0tuywm7Uebl5
XkMIu65iiliq+c3ncaqlbYDs7lSALxDsej9akXxjBeVINIjaTibBB2Q38kWOQlwHk7Q14IEMcGzU
ePGpIg9gRrpob9b90UpQYT2wK9ODXOf6jDrMze4PcLczldnV3IjGh37H8vqifAoypBy/EvHZg8Pj
3wRS4/oBFsaqFLeayw+aKONxHlFyxMqHUv/cXeTd7/BGyP48iPKe8ycKArfL4A7OJV0HNANFp7Y7
5y66eQoJ+NOKJ1+YsP6dwfXc6BTiUb4LnO4dTRECaeyIILvsZCxypQUbEmRlB73uJtXRxGdzOgM+
G2S/BmJWlBZf7ngyHBqKE2Yd87ScDDPCFXE1uukZIsIB8cEMzdR7tOGFDEe1kM+9ACga/2mXnnmW
klVS4tGcMC1PqL0IoUN2SACpN2q3EFWlIdz63nFSa6bEb0lta1+vREQSuJuuyRaniIXcgrmzSiY2
UJf2OpxXHMZBhEwMB1kL5m0L2gy7EDKn2cWcx657y99hAMzUlFUM1mIXu6uicDUAH2W1Jlv+VoUm
5gmefTZZ1pTqKseOJDCdgzy06JO96oi8CKoTz7WbJyaK2a1siQEShEVRJ9klR2OZCFeBvyMarbqL
zI+sUHF5lIX+4z/iYHcD/zzsUKdA4QqoGU4pdU3xzORaawYHIZRopfitbl7N/2cfCCUv1PU0EFjZ
8MC/Xk5z4B7WaWDc81elpmMvtQSOT9au09VWktBCVoZZmJ+do2yWYpkGS5aJhMKwZaCzeb9l9di6
SWCA87OBoY+WC1sQtOwrFjQXr97lS4md6YrADCa9CoWhBWgSzSVFTLDLG1sabFi3oFp+VWYEPSbF
SJl+jVCCshNZ4LqdPQbSG7MjeRgYR2swJiFGy2DgUerlFGGkt3BZMbhTpQ6f8DfLdvqyTO+h2aAm
n+JIgF/uBg4wD25HTdl9rJeqxl7q5De0/DGDJ1ucS5gCYJaeQNQygaWyaGc/lpKvn7yCCH3qALo0
wyLOhwYTBdcskWS6u1rF4PKecEgPudJNxgSrGL69p1BCBvlytlvZi9ug05GzBdtkZCdI7FoPBcTX
9GC84a9/l0ZveCoeeLlTyi7VinzmVI6ge/bTCPUMwaiq3Dd45xwf01JJR9lR6EaxRQ2HlRMWDqfj
UlkTuUyQ1ALcKJepAAKyWC0keRg3jRRKdk7oCRh0kaUID3YOuOFlOnmAQgNB3BylkGAJ1C3VYcq5
K+5pS4TD8HfeONM+5n4co+dyn4N/mCc3710a9xiPWyZ14lLjcLtbr8ZhFy1fRx4wU5F0umOg4ckj
oUHMX0j2AMvoaEhLt5iFNpZKgQnt5zl9J56qo+XA0iI7ON4u+IVaJb7XTNv//fNa19/BcwBKK9bJ
X7X5O+g5qFyef1uJp1V8ZjDNDBJ++y6ejGo5d+LRQR18LdFIgG5MSjW8B+xPuzEAXTyNTxbVpaYn
6X6gDZr0wJAe1C4iOz8xMOwNr+e8Yx4q9A8+3AmpHLnbyQcdxjFcXpCvaVn5PqIMddOf131g7D1f
+H25u+QH0bJBVx8qj8gY7yRs8FSSuVt5ptSUIpeQtSb8DYW4zYmC7d5U1GPlncUXkPU836RXDCZj
sOu3f+pTz6TohmKyXJLGWmQshXIXkueAe8t8oS8TuRuahz3meKdwuX2MEUW8pNKAjSn6tAXkZefF
MOxR31RiFU+SQagqTBpzGxZIk9uKp2Ezt+/09gudXmsZIRVRCOgOkdn/7bueKks6/IctL+HKFKVa
xAauxDntm6ByolHnQaElyMQbo9zx9nwCvO1vAW7QFR7CyM+y2l0XmaPal1GmuR8DfJzh2gTFH4nt
Prs7E2p1b/9Ibe4pWrDQAuosC9QeOsxRQUCXYRTYa/bck94LyG0j95cdZ4o/DHrVgF253yWlKdCb
ddgpdFaCqvOcaA58kxwlBtVNUFm5QZkwVEK9TUU8sEmTzxRaFu2W1+/O9rEX1pXD3ryB8bE5IWBO
GzXTTz52UCx11tpSJOoMXRmOe1lhxKxDNtvIvoQJKhE0O3Jtc7mF+FkAJdztQbyJ9i2j6KumVMcq
NKTCF5k+Sr3p3QiBP51rqd3PCrK0UZEiU85SM81Ga+Zyqw/qgin60XboYKL7FGofGStWhTUS4vRI
v8f73Mr4Bs+7pIxhXjAQB2fJ8WvmgvRZ9ASGjsyAce1zru7xKnkQcCS0UJqytI0yhwjtg22XDLkd
ZoJabo7vTQpfZOIq98o5p+StbXKOe+KpOJ9Ty/VgXEIciJRHW6fLgPb88PqUI8S3vOXfEkEtiQur
OYEmKBCOvkMgISjHMijJTJ10vv+1u9zqAmmlRAGW9UjyV+QqEULyLOymxYtAm/aeg4fJIYdRL0BG
UxVf9Yl3dT8Iv3cgXlCr/5f/P+eNqykv/CkJgwcMqDSNP1IB4Y7spknR2TbdRCMSHI2ccdWY4SPL
ws3Zo6ODdVwyraKWLtGhiE/LPHEp6Zs/LUZEvki/HCn540P0WSfRjZ/2BDF1ki9RIU+RYvOWYvf2
mcFZnLhwFNyNKcjN7Y/jeJRsM7hePOyoFDhRSTFI8xlRL5H9nvNPAtfpATMFA+9jqGzu31KZkRE7
M39wC3Xnyn9wJKpkFdDfTZPxow0j1hTl2X9v5ASSge7UCsHRWZsCEX3T/Yb86mbm1POP1CXL8NC+
6GUZ1yLtT+5mzZZkI01T9G7E54Wd+ZvHOwdbMhj/gafK1gTZU7fpx8bWMNbhfMkgUXSoLue32hcZ
jvCboUw6Ec8dhMyl61bCM1/V78fsbg/uVOA/fNpWVpP0Bo8PGZqGBwzPZEz5bocChTlIrPT73XLA
jjHP2yCesSZa1LoIHloVyI8HgnFWZ2+DeuVGW6oHYljua654OzFo8v99oNpN+sHnBdZQRo5OVJk8
kv1uxsBE8pDJ5pIm7a+kf5ddPCWf1XahnAF1cORSdSuiEE4XJh82h442C3bvnMqDcrfmY8fdZr5u
xxEVwSqLNp0neF2bg6YGQ67sAiOqjUdsFzpCXF1EGi7d4b0Uph694zwn6i8SB67WwLZQWtrXrSia
YHOIh1f+nbrAQ0DyUcHn2AF3AtfQvlqVkMerj4bgFZyBAoAMDBV17CFR2nAnvEEjjjjpEGvHr2qQ
tp0cMeHNu8ya7VZrC1RnvZ4ERY2lKOyKXcwWyqNzEeddgB32fJkR0afcdQx1LYhgcdYkscOx3KlX
XEN52S0IOHgEMwN8KLvSxfUcYrRh/8in8+5c5cS8iy2x6etVvVvdsN75UB8KH658Tna3nQQP1jIZ
DfWxuEgpILX3Cwtk0S2NRYyop9KmLuRIkbQRKKuJn7ghIcVSUJEKTBCAJEmzkMa+yRNQVw+/xDXe
o9VfleyO+NXc9ow8sI1TYqjZTA2Y5d88nArHfV9Gs7VS+rAr0BkRporRxO3VCUdhU1V07h11PQpQ
i6UyxXqQlToOXtLz1sM91c7qloZ9lgpektgE6ZsA1ojhlCMjoFThafprFSXeunmk8K3nTxfHjxpd
Vm9olUFyebJPa6z575B/15jciTVi+0Sh7sBF7uUILEpTgKRUNdqqPgyv/RHq/vP+VTfr2xWquN1h
leO72GeAukIz3I9FhGpuSVguWN2r3JE6jBSSKppkh3UFKS7lLBLGmcKbXnJSncjqPmV6BkkhYf6W
AEhQvpI3utt877BO/Y7zOeSt1Sd01hY74vxgIKg9+j9cCGsdL/BSYuMfVHepQt+ry4NcuD2OLA+4
KC5kdPjzyWtP9dMdzS09Oi9HEZyi6SGEIzGBBJFRZv1GsIjTNgc5kTrAZNahhQgClgV5RoX2rY2M
vj/EiIP3u2LhTVFGTFrS+hhRK0rfkCLuNgiRbdlApuQ6eMaX9nf9/viGJcu65M3N2p8INt7HUcbu
Ek4eUtNDMN+dr7EGqocE129nGXdbMeuoykKPnKmWsUxF9eRtXPKb4EdSZ5LEqA4Rkna4TZhw5Qg0
sM90M0O4/tw/qZVb434nHAT5F70OrDh5Ns3nVmMxsMUD7Yjf5orVjOy1slxrqMJTwR006dlv6LIZ
KliZjOIWzh1FM5OtqVKro/eMjRDFZg2cfjsbF4z2iz/PUOGlaebBTdbiu9gTOUorUGtPYmqvoxAs
lRHOOodY5grzTZJKHTbuDFC54Om5jI5GZpxFyZcK8KORgxPT4Z20YrMQn9HoPt9y/4Totlobdf8+
Q5GOSj3+DO6JXHvsR386hHXGzZPNDMbUQ69FIfFbwb8Yqqzte3N/0DdcbastZ1R1zARYNupLXTkJ
x3wSeaebNz3R91uJ7U6MaWIfKKcNeqh+72BI7N9QwAIzVqqYtkC/HVdJHz2vjplNBJrJ7gSgwMr4
g95BGwKl47PP2wcBGaeofRwo33g15Og+600WM8o4JW+gexlDceQxHheSXbY8w6ZuyZEnNGxDl+JO
93RIKm99RzgsSKtK7amrAEwqRPYhoGDX7SpKz9BWLz5MQ8W91/ZKg8Lqa5AhPtoCBBhyp6Dsurqi
oLl+wv0qXGW9TXZv9o87FUVzMV1S0iQqDL2a1y7MhlW2VjEA45PlmgYmgESOsUsYpwUJM5JilcPS
/HGd1ePSnDO3HWR+k4/kVXGzCHEn0MenjdmkX+evNYmE/JyyPkj0czhOkusBYf4r2CtZ1QEajBLj
ER26beusnmeRmqxvOEq1ZQQxujSKtr1oZKJlRKr0A4J+BcJV8HNo9UmFPyqGWR+x7XAu4Humy7oF
1ZJc5/GSvRsts9aQhqYnwyVnLyatoRhQMVFVmcWCkpsgPUOtXhnGq7u5eUyhPCrTGGO1lRswbckt
Gl2COirZoAXurYpqAGUSAQmzJFHyz+QZF4PBiOQtPQfHbuWxRf27Wffo1QG37CPkrb7dMCvsKBNJ
doJhZFoY3G5kSdfBwcBTtIWUOkwj2Sil/iPhvDLWcEZnu8mnDgkjmzJTlOj55eQ73+CNJ8waLJuB
3kG0Mzza0QDMmzxPyNu6NeE7IoTKVnQGsZx/w2+TcKedBo7j5pnZNTWPG3sUNqJTK0EDJ9/vKCaI
9uvLRwAS/eOeX76FyhKG9M7RDLWzLgtoKbszUSdnWSVCIvbOakgcA7fKTFqWzidzW8EQjmo/eNaP
KcwactrnJL7dZOgb+rR4IqwqId5Kdm4VacvlEhXM0qCqhJiYX8VJs5Lh4CWWfVL6nuQkirjcG0zK
t2KfJ2pKsQNxK9cLvn+EMkb2cmejGJjNovcHNMqXwZxGUW9kf2+5ZkK9c/LHHc5hGCELWqSW7o0T
D9OjjJhIBrZYRFU6DxmJ/FGD12gCiuxQcxodrmwp0xzUPPt4Ot03gc/TFZjLnK9rf60xPS5nFYST
WWjKMWxtAgZ2RGpx2w/OcgDNPXxmkeXhkq+AUipNURYO/wi5OWIxkbyy/Sjo7whE/MJySJQHbw0k
ErQP9/pKIuR7DdDwaYedkavvq1NtkGgURF0kacEHbCMHJYbGe7FDfaB8kegzIuNA6/krWXfYWGYi
4c4e0jLC4pCiV4fqS8SZeP2W5/RYLTFCLpiyZZap1nJjHMQMz+gwKcyrdpvpoxm7XGx12bjPyUeV
kwJJg410niI3X5hkt16+Sj3skMu8d7LKM2ODus5+GmW1AoFIK9iR4FqrSLd6l6Exlk+Op3w7/Dfk
Okc/yXkiZ6zR9CZ1YDEekCvoRfo6Fnvpi8gpewgELN5c7BPTzQEOuuCSzHHDfNN/1LJKE4R6Ocir
IxrSSjNcXg6ptdO2whM+oPyNwjY4kkTw2CkkLfgX+5d77mj3p6oc+7cQXulps+s+A5F2aMj2BRI7
X9aivf1toiHv+y/m30Eno9cc826KRIRYYWPO38bCkHT7ZrbcZO6Y4Zy6WfTVowz62/1Cvf2t5iei
K0PhSChYthlhtc1clNsG8M6nfc7ZDil4I2lAXBng9KXDeaSsr8kKzbAX249Kd/9WSgG1G5bwaZkr
k3XnLH6IcVN53FJ9q3t92hdbtChnz615Bgl+xy4eMJEngBtbmDI5YkBB9sjxKgfEnDZ/JkEO7BKo
HNWE8MDkEcQXFo1YnO5/StBuMCMEDYss88mrjkkpBFTlwsVRq07gSiPzKVmoUwi2GgiV5oXu2zXK
b+yvrDezxLk7dZPT1WPCcQNXNQX9BUXsaTwB+chNDEFvGDT1bl9h84EZxEiNVEogbQZmzsPHipdN
rVoHFjQ7McNCjJnFhryUihzc88ItxMif03xzB3o7Ft+R7fCRru504OqB9ICkEOBA05Tvu4bG/VtU
BxJSPEGBijG/iA8AkzdoEh8iO3fPjqpVBTA6ZRCO30zqc9T8SEKNK6adYZgiQQwlIrjbOP2ds/J9
GPbdowrVbaZ8lvb9syLlEJ5IqD6QZtPQZk35kBuT/4QC4lg84l9fRRP/K4Td9x25tCCrlF/nTYzX
y6uUK08pFwH4IeHdaMSKjoB9eC13LEpL/CVxX8hyJ+LB8LrylNXc18JQeC4STStgwhhZTQUDWrY9
zWwlpjuNIzw5zfiE0bzcM7z0yKxXz0UJUdcpqEbpZ14dJREDFEGN9KGOs2MJaGi3NCX/678Mnu+z
smiD7iAQbW/ky8N9CFN0RDKKR3WIhtK4lSiJdoXeSXu3GF+4S5l5ZVF0UgkuKAT6FfKIDOKChFik
w0orwBWwkbeSEq1cs3HNWkL8RalNRiZakhvpAgdisIYXzaHJTIvIWleYczuf1yonxeBTkSy5PgUJ
/dGZ0xsQqOV3dazNVHlkBIWuajkcULoqrub/+su1F+9wR6c/ilBJ5H6ID7q65Yg7FYtM5AUCMQQ7
EZeJjD98UIkxohv7/IXm7gQ9gM1M3OJdldlV1Iec+4asDDbQkBQUPrbzl2vcleOy3CmqJCuRrTHy
+BIY2Yixn6BEEXNGh6d/trTxiBSn0JHSOrZCK9uflOFrvSofhANbc4lbPpOSh0NPDa/9a4THjBsI
+vSxXAK01gzSq4BSxU7VIgT+Ffas7B7FEjzIIfnwN850PdroOrrFj0uU24pxT8rYSDyM4YKpkjkS
/rUkXl1a8i5Qw4lY6soxHXv/PJ3ueEHXW2bobSKaB2SSSkGQgBlO+tPPeEuu1rGSQBVXnhmlB2hF
bRZO+nQEwFw3csjkCDPJlqDFqlSgHEaXdy3XeVuUnc0y0gEOWDpbQ+hJMN3M3LSbkHgzoze0IG8E
B5DhaIJOY5gmNaqCJJbKV04M2mL/Xq7AFtK4clvpiZus8BsynzhPopATnG5zAPLNUK/uaDIhRBAb
w40Jnk5Q2qI7cJBP4QqWJcdp0Qepno+jiJzt/oHvkYApITSUIfqNqaBiKdX1QHqzsTSWNNrY1LpL
vkM/3YhlhP9rBJyN6L4unvSny2t2SaVqHdAeHUI7gnUaKDj60rj6JUDxaGaJmCZ2R/RG0p1gy2IM
JES61OkC6WgQuT5nFVsmAHAJLNDGziLS4k3exiDt5BGNTIrHaf3yUhk+nsP8zQlKy9l7timnfUey
lWdKD2d1/GdCfkPHWj9SAdKPDKW1fXqzWfgFSC6XQsZLorcPyI+KmA3u9rOlVVHOuXpXzurbka0L
Qg2VRtE+5fNG4nL54TCqxYmIJHCkulkZg06CY8KWrkFTTv5unqLOGLa4satOBNORUkOy1svw/a7j
QWScBF/NT5gSkNSs0wynt//KKPty+Us+AOc7PCozPldSAy2bHy125gAHsw6ppQbA3zNpi64isbHG
tPq9ADuWavAbQ5YgormftBCqTkIIAs4f7kowDROXxCwsV760m4ChmTbOQiDe0zmZPIQMFg5TW0ll
EgeN8BSDPWNtsMuy6Wb/Hhr2dHmZvxHyUvaLfhzxlr26ixnZ6ega/MSl7aP9anbMW9KbRfTFnrcw
luqGFSiUiNjwbrKsYMA1tGU1Gn8eaNKMWC4f2azwVKuz4etYvuei6QJ9Xyc66t4nQ230yl1CbamF
lEpCM78abokXvJXCoJooOESh102CCYJsE4FY6KvfnSN7z7bBVgsq8JC+wiEB0WD+RWVPo/p6bAIv
32hodUNIe8FbSE3XRXSsyfrDDA2ztCIs944l9us8pwZgXCu4s9jDmMhXYC4INcme6Tz1yYVOjJlz
t9S1SGOk15b7+Iyz3cUk+VYRNnfE4hIZaCRLu919Aqy8Sx+4R5UzQlUHXds15AtlIDc6enzUAgRi
nveVr5h+ht7MRY/VNsyV8U2Jh48kLkhLG1UtSKRz9PVbjsiAWiddpgesyXcmXUCyTVouCeVDkUjX
CAAO8rGhpZNhMUC2NTRfPljUzEQlJe6y05cRsitd9hH3XrTU6GsZ1SGK9CmfQim8sUgXsGgJvqhi
0VYdhvoErHZTvg1DbCQXRyXIcI4sRqWlDtoUp6N19Te+lZk/etLFZzDEcKQKDJxmy1fcd2GORu0m
PLJP3jsY4lAdc5wR0gsmxoai6Dfc5LgIT46eM4KcI43uRGhjsQMsRX3sfAPgIwVEU9iVkNf6NTpO
lce+HyOU+dySRquX7L665IrmiuQK7LX58jDmlpFFl/0wkKEhuYRd2hoUwAs8Agjoe0MCiMmu5MU+
pnKgCEavREK1Btn+nPwG/DJzA+TptFtf65p/WT42eeIoN9G49YnJkaW5EvMi+1SaBGJfhELP1ZlC
8vGixiuf2oDVEfZgTPh6whBVLEgbND2+aC9WoB/rxZYBZ2A4hfdl3wbDCFbUmz38As6hAi0w9M6B
hSAS1LQ+4qRPTZoC2tx+6vvfsgJ8jQk0hcg2kGVfsNhpWh6Mt8ulpg4YMdjulx5ztzkohfx7jYdo
OcHC7a5/RDw18cFtJWuhk7+FuKmDgw10OzLKX0ZZvCh4eUSvnQAzhO8LU17bXfL6031fuSjBnVJ1
NQ5oq152cVmCQ0q7Sfw0ukvfXEpDNS3j/t2QjfybLpyp5Y659MZcCjDiizyHXlXaejZGQsconGc8
rbZhKA/zhOrEsMakb/HW7Ez1lr42j19oSk7WK59vajG3aVlhcpZ7GIBdHva3jQx1rHblfgL90dAh
5PO2xG4zeBRwEypZZ9Boz8t46WurfpaTfPweYabgGkylKd1nq8uuolfbSdG0bz+TqDjgYAptygSu
wuC0UtaoK1VRYgogy8rqRnrBJfI46/ySMK7nOctADMVJns+0BuyAMGTW/yY4ZnzMp19whRt+ALnQ
MHxk/0XYEoW2YnMrazhZAyNb+1B2CJGPF9Y5TPXFX13XNadhDlBfJDlDk4eA3KspxbWVxy+ybqCu
8GyYAAJ85r0/fpqwTX8cr85VpvivhZhsvSVK2H7Nw2usSRGumkEz2kCFEeddH6ifKasmKx2BpYNA
YTgFs1AC3Deq1CmfsA/xgB68OBJz7LQ/5wV91JpTd9LJ6p0FMmUX2ac3VJaDiSVuD/bB6/+9Naou
S7quoilqD/90mZkisc9O/bRspEtU8RcKqrwCYGCKT4U2kUs+HF1/+jx/eItCr1I5F6OyvzGj8dLW
olqpVOeyTgTSCSbVL6LEfiFubvy+qQZkWZBIKk4NtS7p1TEvr2nidVpRh8Q4WFckqUUw8oQpGCb+
56E2UtR+p8v6OMQdUngUkpUqqYMxtTQaPxWiBOkKCV8AG8lRpdZnWrFjkzsA5/w6wm94uu2gncl/
qt0uUntTC1LeSgI5erb0DfQ37gSuSXOSWby3CJNUoLHuqK1+9pgBqYCKnRUAV8DcpKJtqgpE04wT
98jebPtuilpdw7o+BMwZiL26ocB42fNK10DFpS/7Gk8DHoPlINKl2CSh3s7+IOhN/e7FWZNqFMvd
4lHHgRklaGYleGyIM52oBqPoxj8Huo0lWHD+qDjSq25Gw6RLjadljA1CCGBTYtIL89qQf27DBNvz
lajnu1iNAOSWC2yJnXMhbhdFqTltjRBk5JHMkt+VlNjHHgVtyUtv3oAVGhIhIE9vgC9QmejqKKdp
COb0P+1CoCyNOEJuCIvsOTguia6xYerh8a4soKszua0VcrTfXiJezUuwP61lb1Ea7ejGg0M7HpKA
lcRiglY9GzTKudK1kNBeGsHJJ715za2qUGcrJ6Q8WWNoJXclXazyA4aOQhK5P21f+3hgJmBVj4NF
g2L/Jn8/RD3XwvAowkIfFkD2Ivd/ykAm5xYJAJVmA6jwOVPZVHQ6u5EBEsiS5olTzeL2+2DhrBRk
wF4okQdTLbgYTDP26Ztqo0C7WeEAKD5Qyhx4TumwOMh1U5I72tCZJgANucyY1m6+S3HY8TT6H2e5
M1F/BOwLgiIEO/uf/n28KCfcDqn3SzEVTZdPwTVwmfbwahdh4OMAmg0ZaYkHtdQudtmOVVpUqJE2
hHML3iyb6cUgVUS/XhucY50aXTpt5s4LafMEXgcXxWVnKs9bmiCJLUHojPC1pEqmTReG9jZasAim
riOFcAaSFM8sGpHoogRbmHQUUqTd4v9Dc0wnqwj2iSatlEDqOsfoR2VC9C2iFmVRCoaW+GqLi3MS
h8VYU0TNqZ0gz8Nahxa+Pmvikd9cJAgvq/Hc4YdG+4zuGkmrD/b3rB16RvBEFpaZ8Nim7LHyBbI+
pmDRQDMFIuu+shhiep6Omron/L4T78H7kgC7bfDKkbEQWoAt1vOn88g2OBjc4NvX3sjQzHOql53r
5W5iAClAxRXxt/VZgQyCo5Gtwxe5HvQD6ZXLjL/Hm2ZPrjGCkR/rCJQpsKwo3Bh0pAkBli/dM9h8
xFwmpctEaxHY1RfVb/mh8sYjwafknbyu6jwpqDRYSUT6yzhUgF8wlbxS/LO5FMK5WQL2ylVSj7F4
XxGG2UQW13qcqGOw+UhBWX5WxJZRvrvdpegiaI57RwHtQI2skWpuSmhKq3imrRWoSClKi4DIhp6k
MWgcCHYwHd6TzvrpORXYNtq4xAF3F5/NU3r5sSDvX+qGxlfqXuO9rtgJRNqkJf3Pga9oCN8hrJvB
BhQy5gyOy+D24cASGZfouf9e5O3QOum0v0WpXz8t9CIklyciq7otRdHXLkbaW78DahOrrTUg5LwN
+mDMCztOEZOORxJsVK70dvssKHAd4c9q9wn2MOBcze05A4GYqTLFqgiHcfw85lMpD5Ug0FRx+0Zk
h7sIsKd9UEQ33Yc4Vj+7paJG2OTDO0RRrXlPdiIVdMLqRw3roYs1fYg4njYdb6bYfbWjdAU2tcXR
sXYb7BRrYDjpad7RGhpD1vBoZvIen7bJK2ecEGmUXBWLWd0RmPLQPbgqiZ2PkkzdqRDz/HvEIViZ
vazX/AzCV0CfwxVipRTn4Zg9KSklRrC1OUvA6+VNV098yVt4NmDW3Cb3RMSw0SnnR9teXGa3JFe1
liPn8JaFGsNWyN5NuWLVp5AXq3FwxvuDsB9oKslD2rfoTV8Cm3+uA0qngHgQKb2en7QEXQRjoqVg
91p1a64+rx9BCSfrWTN0tm6I7qmwxebAB8ESb/6azGT021D7iqTdURvQstH9LvyAeQHrx4wI4DrA
d1eHWkPfZ5Jrxbzp0Olw1MpPVUZclbi8U14+w+/DK/JC+CXCkefpT9/skMh+g+EpqaVmU6+J+ii/
4QXINl5eAcQqM8GAJz1Kyf2aoUmmbY6SSrgaMgo24V7MfEuEEs+6JeLE/7jcxD925EfEqVmDecnR
pHLp2+60y7/4/NLVtCQowyZ/MG8fZ5qUH+QNhoMJb86b2IK2+gkXRqAXoohOiUfR/KaVOzvHSf5V
x7K4b/xhA7zHcMD+eyt7laqo+XVRCtXf/4qXf/YN3fNSAkDQZigroOBrETrKJK4ohjPRcfVi9Wkj
aMhVBNeHjAyE9oAghQxBRa08oq00y5QdfNua7YP/8RCu/UrP+zO+d1x9LQkKr9RboexPqrOSHNI5
4IKAn23ZqyAVS0DKH+1j5x31I8I2VRk8EEI72Z1oSzA+Y+3FwwGEfqX6HW7DNmcCRtFfddyJGaMV
sijJaCOBGXEueF8S7s6QbxVfTcAD+BoVrm6kSRyH1eXIBxEn6/8Zu5xniPlAUocpm0Dr5hha2SR9
kJTiGsZroiu0fIew4I6zc51VUwD+SJlFox+SrQljPCrKFnuPHkZuAOQxQV2ShuljQgV7D7aNxDyz
7FeI9FrSQSz7yut2fsfW9aHgWUvyun3ko8sBbnSs/bklF6WjeIiyCgZWCnRbWDwFwDqWRy2YkblD
HXyESx77kuqAROh75DvDQQ05EstjmmAq2icUuJiYTsQRWwFghsuJzFT/lyAw/hdiSDKfbJv4Cju+
YaO9IIT/V12O3xOIdweF5v2C0vnpYzFzuPe2LVc7e8GmJ2UVAnMW8gKMsHsye3z91GSJrOAJZduR
iIkAxYriBidL6a98Z60pL9LtQJUcesyxMnt6QcLZOMa3mPf2hBqjsAqXl9aAhQXmREfXmQQDgjmj
/aXdGAy5qe3VBNB76r8sh4oAQ5oosvBlbh5QEJY9rKSXyeloloa2h4LBsTDZyySVqyPRyPWzJNjn
DyPw9RdLYAKQLyNx1JOYe1SLt/LY6HsyVLkx5G2+xYntTIixmcyVprk2HFsZS6iBxJNeFk9mN6yk
t0hkRv9iHbnhKtZ6LaJ1/0ryyUymVtGvD/KEGmlBTEJ6KVCiu7gVcx6XxfOfcDE0HpibJY/gsVJO
UOdRJtsPuCWyKRNzAYFMQomyz+BDjvjUg8d14wb480yDqVeOckynWG2IfDYWBOxn5f2yq868sHQy
L+3rohq4PsAQiWjJ49s1YMmgKO0bOTg5U1gO3n7PAguV/bCchLZMpBMHBmKdD/IrQKiUc9XAyCwU
ELbS3lXdPY6G3lM8lTxJwu4YsOqIOY37sIGzl5TAjnc6TccmLImK6s72VN1ApSfJcCWcRz1zlik8
mEq/6Y0jVk6oa8dxRqZLbxmrqiQx2k8NITmoAAV0H9bZLwg6sK+Jwajejj96ngxUoLa7aYLmxJXz
RpGZF6SWefrlneDhFxDLlbV5vA4ZQiVL22pQ0Eg+SlLR2XuHCGmnjYdtMFlXwE/BYhTNr0vqHe82
Du7gzRZLCOje/XnbCY8DJZ6IX+2HtN1R4KnorYiwQ01keKqROWD1IMGKK7rI9JIuOaRkYEa9zvL3
NlYFcBTk+//mtV7B2jRikyGoWO+k51cqq9B7prByjFw3KyQjZYLoFHaGymKp7GWJiJvMgHKgFe9J
R5zlJ1XbIYtRxhObXoouqM9psNXAXAl+l9yux+W7YeKYcATpJ6YA+dwy9s0X4jGcmhNgOv6NKidx
sHNjTApVTG07zIX9IpKI5j56pO0cyvWdJ0zSKvCDr265M0+lFgQiGFMnlEFfJ+BgB423uF8yRVl+
7A+w4ghxJJb4GmPuD4QS/6ZDUgbd90Rwom+mu4pIgVVLsupJF2T3UKpM0snddXsud+oF1qVAB3SU
thpcKGmS2c0IwAnfoWEkDVveKENCtddxGtliridScdq4s489zxjSlUgjtrqoQSbjCUkGWx2iljiM
Igo4+N+gMa0twJekiK92Ihb2GfMbiK4tBZ+/vN++6LckYEzOPhCmBg+jmKbfPK7zipwdvtYbUQg7
tUFtqtXx81c/3BqX4o6G7vzXOXAw7eqq90dNXU/n0CyiBfXT5k6ZEvnN9OxCsvk/0/gA2eTDiNGn
Q3Ri9IHyrBqMK3RQX4NBzG05DhgWuB9WjG5y8maU2LcTPH4pns927zzerBFCULpH62F5QhmwYdSy
pVR10kQBCxMclaOpl9GBGZ9Kdnndk6ge5mD9trX5KUxPrenK/yp6NrbdfpYnb+98kl0GBnI56b+O
P1eLZDV6zH41jyneSAUc3U5cURiuTJZQ6Wy4G8Hdq0ZOBj1zmC/Jpt15krgd2zbPNpNQJZKV7rcl
x+BFp1mxpZItR7sv7MDWKxow/qt1lxDS12QMmtleyLEqda6GBTrD1WAaCU7HWbe2FH7Q06YyXNHu
S2zTopZD3N8fN9FpLKVm6UVaj8ojwQlcldsX75bWubm5unsZ55UJ3Vq6wDWhUuf7xFndH1KkMDw5
hphhSI6Ha7SUbLGLXqdSPqGTszgGZmuDnwhpC2ZmlvtcCzE6MoLOlythDlpqmS6EqU/W9zXzz2uh
+AjIq5lKMVR3hw40WMUsWeB/jqIDfs2rPOtDtTVDyxyjdJoMqzvgipC0WXmXM9AaWbPkOjl46gUB
udtsYxpdhltYXmF9eu8aPjfbV/TOGQiNah98cGETihPEMhr/QKAw2/MnR0ZNmXE68cZNBwMTwvaI
dSx8zoo5cozFNIKdYXf38sMRkSXbRZjy4mlzgd1qWLM+etzaHJXjbw+GfOiIT7lTWr9QH+FSBXS9
CPJvr9sV9tb7OqLG1iOpb4NdWl7aBNNP1/wxGZgVEM3ZwsGB7Am+p9+Cole0ZIc+wynW7eq0lSXx
WkegMBxaHHkbZO5GJNyTaNI7c2hedAf5NyvUSuqkdGDv1w0M/WacWj6L1gav7FW+7Vrp0KBID5ws
IFm6VobphELabrd/a1e8/Nkt+A9mvTer+Jfb+V+5ZO+y0qLJQAOay/hln3+GJH8klPRwTYLjVsfW
nWEa5ydlh1ncxUIyOALlQp6rQKnNiUWDBTJw2zWLFanx2xU3Opy/1cE0IrzF69lw6ctxCZdiHlm+
FJz9/UEqtvwsvXCgdvHgTd3fS0zh4Yf2ip1dk5HF8WWBPqHGaOxJdzQbK6cANUmRZzaT7T7TUs3x
KP8sX050St4l80BxM7HtFMuLH5ReaSFKVX6JPvs8XIsr16VTRbklxYXifQKpYiTbWl1bONd7quNY
A82OqQ5QMXwBkYN1miBW8zSxj5VuMbdPf36tnjQ0qjZc2k3wMommyGvcnPGp7WnTww9XnFybpoA8
FlTWoWEwtG94w9lSEUmZYsGWw8cWsIUeLyopAPU6VyHTn5/6IQpLkgqwVQtO26SGdedGcJKRyopY
h76rKnheb3KQZCEc7GXVFOd1krkZEMeE8a8ZskyhWmVgs0cu4R8vBLV849oqvb1VYKnTmXQwxLDZ
DFz76d0KKdvqQM/+bvACyHLiVVIxWIzYHkWXtXdFWaYfwJLvci8AUVwVWJK65q0VLyeyaH4PukjI
+bm3Ali/mzukVed+rMwhhuQFrp0Rd5u7/LYSRxSXn+kN3fwxquFGqeNMLftOVYQrkmyXrzYbNzFu
VWkEOAj/QwwkxGCH/V7DaPggBJXCvcWLimO4cL71q/fI4UI0xGi+k92wUNCvTqflNAfmFktdyXSz
IfFOSijvX+PPwdxHf3+GEWhw0AsfkdBJ3b5KUZFDW33E3cL8r9W/uBb6Pml1yjxZgdYMpWXd6ul4
Z7Erg+j22EwFPXkyhH/ESVtmjX3JsxJjmDrrdgUzDKmTBn05o/PuCJoI6cgT/sEo8zyhBvPw2TlK
iVETaGlXwue2flGfaypdS1IQ+KZAGWeccWRJ67NXrCHAY81yMG5EHLvcZCJjaSm16F3CqENMVwEb
p6bwBxc0uqrozj2mS8yJmSC9EF3sgYLC1ujazb1Vm8/LcbmFvfUQb1nQbu0IqsWkApB6ydvuJVLP
jLXhBLuVXK1av0hd3lA80+2vWUQCgC6oqdvo393M8JBJmxcwrs2tzgzYKDOmFPTfv2SaOdTtOOd0
oCpKSXJ3E7X2LnIdtwAM8oMgEUnLdxJFd4dYsn3S6pinHja07mGMHXilHJ7PTH8HuZLfPXOK5OMB
TJUxp7BOWgg3CWoa3qrC/vQ+OofSrEKME7WmoFlHMYkgmRVs4yBGIoU2C674JfQ4bS1NrujwLnkE
4ZzLMM0kSF3lFSYPjqvaXh86fdlvW0Aj/DWJ63O/SbCVGkjYm4yjy1LDbAYFg13fVx/L8hwQAAxL
5PKdY/XBwwRMu9uJ4IUMr2fciSqAFv7eXDi7bYxZQ8h6nn4tbUVxDG2NXdmq4G6Lt1Q01zxJWSsD
pyyvBCt/1hCSb8FC41xQ65FVt6o47qVImfwGBUjPKcOzFNgDDfk+l+PfHhWXBwP5gUv9/1wYt3pG
QWkwXpORtV6gGv0wpn7ReSxUhA7jJWhVZXH1kLTrnco9AO6uybsqC8gC0DwElm6qsGrPUZ9il3wd
6VdfLaQ0kU9U41XDfdGrjJK/aL7rp4/pRjM2OjH5HCTP0uvCa++WFMCv3mP683P75jiNek7NiEwL
CTsdrg6oVtmq0tYo1NayMo8RLwJPRlGq9VqMG/y7A9bt5+u0y3l1H9+qnMvMkhb7yS1makTTYIm6
c0FNmGwIX57ITmvoNDrQbSkLtc5JaGCXa5DPG2C1yOg6SwkgW24MyWnKMWEdZBG4SGdZooT/K9Dy
ukjuYetpNUg+d/f07fzshr73tMbQ6uVK76d1slM/ibpoJH3alPVRREcbOg/lUgbtzhKEXxWXrWSL
oKRHSlHLxgTAFWoQqQu2zaZfEiUcoCm/50mb/e6nLJVL4ybPZyjgeP5vgZT2aG0Bnx96464Uf85g
sQEh5Mnm9YYiIBUQH9K+Bsal1ZqMvDCKXoFqEl/F3iiRLV8gnkinra+QYHDxbrpQulFIo4/Eu+dk
UKoyv1CoitkeplMOs7c6stDe1KnFjch4AzSJIC3fKJaBRApmTTRBBiwy7Mv3o1DTcjGnn+ikX0hw
BrEMY25jp/4GkKLKkUrBJDonjEhiCoJY8Ljt3jdNSh87by8Bkm2GV7PUxbI30d611Jbh0HCa1+Nx
5aEA+QjZoNH6ibLLOMeZe6NKqoXnYheLwHlamWF7iv9enyo7OrJLFsNcjxYfStA8yiGC3Et/jxFU
8muqm+5oF4Ck9QSHetD23hwz+ueLwaJjQZ6xpIZNl+7qFiMR/3lanii/9CRJk+i1EX03eO+c9IYk
k28BkNypozHLKndIioX9It7JxAMDKLB6SP1rA6N+lHmy4rZxjF1oF+FV76RJyl0AoWqkuaFbT6g0
b+D+i2qp15FOVYiTS9d8CnpTTejxnfdBNwDMY5ON3fVdKKubo39NQIvaLDT2VmMy2lnA3QSoucSU
gYhcApQs6qJBtYzk4c/LBwxcEN3nY10+Yc9vAGr2i5hnPRO1aRM6JHaFBUet4L4jHP9ZNnwcYMAK
yuwVeMq3dJEh6NAX2JOiF4vQNjC7AZH8N4QnX5yJQYcRcPy89VxddtELfqgHAEoFrTvnBoeeZrX1
f1NgSduqTm8dVuqfZH6BeRNh5hqWyvEOIFeGarUpk+n9djw0nzwHvOqWtndgnSi1CA9+g59Y7xHA
dJ51OmmKk7aTBGaRRDXdwFmjZyjmz+XbFyB6ekwgomrdQnIsZ7XRqIZSYULR+Z9WRZd7MHx7Dig2
7r/7q+2+bNvvfjP+v+UrPoO3qV89EjUqmpVvVGg4d3HbNstkcwGcewWV1LhqEZ8mEFOrIxdTPNVy
l7YOn7+xMFnDESiONo6IpkGk2gDMlseZR+LQjgJj9o/lBrWyun/yMnuW3SUrrZHtqSWnfhh23TGX
95cQMDhJ/cFMRz4EEJ0iW9FFAixNKGNaWU/hM1RVCPZbzDiaFl6dNIJms7Ah67UWfMiypmI02EWa
bOY8vG18ichTXk6nbsFuIgOaeU+TkjUxlFDnXqNsbvJ6/PDTd24c3qz+JmhdsOwMjO6vy8scUenl
w3m5D8/YwwDHE2lsOi/EgaX61xjuyo8Z0cURJbhMmXALUDVaLvPGsjyVFIXb3to1aaI/GYEr0OpI
LT2BSBVowhuvXF6XJxlkp/UEXgwbl861i9tvsNHjLIX9fjJDhaaltvvJfoTyR502Oo2580qqQduC
+ffTwKbHdw7QHfLN2PhFg3rdj0cTUKnR+IIeTQMlYWeYn6IiCWzvq4CQ5xlxILYRyGQAgdtw/i+F
AKC0vrBovCLbgfR3Z6oyxcy0wONevJvRElte64VbbLug4adwsLmb1sh3E4NVpLheGvckUPD9jX08
ZTz9QjGOs2uNlFU9mzN8CEagDEhKA3R5vb2rIEbDGFSw0ybCGaw7j/cA4PVIVXESgupgXgWzO+DL
HHK+bqmXmFiYKe+OxKPoXVhw9gnXbU7HGpMwiuoED7KUP2/ss5EkpdntMjneuMJrNaPIZe6F5u6p
K2CfIm0MOkgs+k/jaWeJ3tWnd7JHl5A0YGoCGc4RgwvB7qi5O5802YNWDYoHLvQYyQdJL7tU0T42
evCSO94mB3N5CNI+QAX7kGogd39+XkRQNbrTVBuLu8ur4MBWqziP8zwDBxIuiHjNR1rsrZOO+jfq
W9AnZniKpNi1UP4qdWRp2vz+pH7xmQzoAsR6xuT+48l3jgDseFb6T2hGjWhJlhdz/1UeGFdyfb30
8f/KKt5J9Pgx4DQaiIYeO7MHHJzZPvN91im/qDtu1FsMGQGetnzK9X81xmh5FFqg9l8SgrTQhBn2
Y2CbrjE/R7wnsnG2n+MU2vnnB9DBRHcN0bYIg3CmOhQJ/czTJSZyO6hTawvRnQH2IBFiwfqZk107
zQ+9RHK9wV4vQ8cKU1HXb1W9nfxXVepf9u0/0ptwvLgABASR8nfbHWiNTqQZJKSczlrljyW4egGQ
+rcPyiMHT9KR9AP1fGOImEofkVrx4W40ukpqhPt+1dHwo/vggEcg8KLlJzi/mugEKpFtvlBLSvmA
oVTs/eDHdZLpOhVp8NBbYEiyKgUYjQqCwnIr50wm6bCSTqbehPZBhraUIuP/N6hVPuMkrD7Q4Tt+
ryCvB7hgWx7ZxvlI1DP8zHiMJngyl4N1ToCWf7sg6zwe93xilhMT+7SK9DIczQDrorpC+INV65R3
6qhH+tmzDOOk7oc6IJURI4ScjRJPNPNF9Wb7mAdJjGxYdMEQIyIMUgit522vsALCj4NUA50BVUkj
w1iqiuL1FsBYGsuIC7Rvqce8/ZkU1T3PBfOTkV7ypigvVfkV4XV/L0AUMzGP/WS+KMa9ItuJyJBV
vt+ABGG9crTwmw0JvEM+vQNuVkpx/CRsscfGe3RgOu1Yg0YXqd6zBM2w93H7Ay49XCIOpt1G2DHm
JKXGUIU+7jxPwtYNF4u+2Xw58wbdu0Vv1dIPJ7LCutDU5U38xucEBUcPVPb9j1lcncX6++aFl4Im
tG+3xwBPXYInajqEKtjgmYN7uh/VdzOzL/3jfXcttDmz/KTstUpgSxgExH+TPJCMkoRrN9f7ONvz
Q3REJipjIwLZsY9Gqy/M9SLIRGA3544VakKDLv6PKqS1er7hWjlyH8tBW1hy/75KfcCYZBCbOtoS
EMX+/GtOOL9JpdvTgb5JMOsHgZLQ+EOd6eUrYQgPGuXUnWks53jpMHcPnMSTdEcfM0xg+VXqVp3H
s5VL2rFBXMzX3v8gkglVCNEIsa+VgRM2EyLvp+8ctjpKHN8ZZqeQm/wW3kUC/zdR2D0Hi3s2P6FB
8ROSleoyHs1g9v+dbfKVkH6CVKqXXiy43xgIQs1uuJ+dE/cpupLIRTwqe7bOeonRLJ3H+OXIIf6A
GThI3cwONhzi3lsY8a1bmVyMkGI8corwaHY/BLliL1wMM3ko1RJ/zCmKEdBkgYleEfoob3VhB8QU
cMrivx9ETM8EZO8U9Py2Bzrsuwxel5Iz8kbViE53jG40jd9QS83a7sNcDQNfoJc0MOn2cmct7hx3
9cuEsJan1IBhHKIk5oA3myNXHDkKXaLFDlWQCAx9HjhAgRRGvJiakz9yNZ14OIeL5ujYekjBm8Qg
2AvVj6jO6yIVXa41jkBU2lxGE6VRlQs/GYdRMgWr8/yiVcwTi6DWDxCcKtwwoSQAjDiFuWc0h71F
Z27DfSXz6MSVlxht8MjGxAAtNHu4HRnhzfRnij3/Y7hSUrGCSeUkqhZ7mZ/8c9QMHXCfNi/4B2E1
Pt+ETu9TOjpeXUMHcpsw9DSoBmtkByJBGgKnzxMVl4YyBzcUrp7f3jJMAm/WXKUcN2VsdPGlRaWm
gsdX+hHWcIHR1Npj2wLv6+YmVByBADrZLeXNINh53YSJbvgYyepRH/68lTrW4XZdQQm6pg++u2S2
DH3+Sdt9SNqH8N3WXKnnVSqs1Hx10S/ht2y4KLqxwLCUWRJ8RYmQwVOteBOsR1HWq+sP68umn2VB
UQZw8l5K7KRrMk/tgotATc5PDSCNuRSu5vJ4pxU+fDvwZLq0dDqKJMKCznqmuekcSYzaZ2q7zHd4
EQikyhHni64cQFKXQsJrpfcFvdbXoem9CJa3sAhACcgCr4bzJXBANyx4lhWwC3EmhCmwvoUB3KX8
ssMbBzpnQ2/lK4V5lMJIlXu89yRJr+x0m5Fh7F5MmriVwtIC+hTvFyMqJ0tl6jMmMY7lVbL6R+Bu
DcFtspzMg+SkikK/2InsM0VmJFj9dh+7V41lLWZEAh+uxe//5x0/2RvzXIvF46s/95fhQTuF7EFx
sUSSGLby1ZuEqYxGBZErjZUv2XB842YCAtv7oItnZc6BUZf7/FZOEg1uxocgJpno/VpesYVh+MT0
hyACOOD7QN+2vawzb1w1d9WcbxhOlsLKp0BmhlB4qyYjzdQHXyp4CkD9M7EmWwTM6CUdLnt7jqoh
raK0EfAua+0jWI44YASw/VtoMaYPpWUS0W6czQ7kXbcMcZxy93co4Yx/eOg2B945/Eou9hEo/XCt
Tj2opLKLUn7bqPvbk4ZPW3qXc2PL03lj+3SLDP7UFhkUMB8tBAPqBEjLWhz6PlTsDLhRuELOwQo1
bD3Z3wOcVS6ihEiuZB7tPmQnGtL0fuY9GCg2Bh3XBG3YPs/qpy891UThKBjakw7qRmDU9JsDYvJn
muRuWEMfVrgFwi97m4f3mODL2z+plMI7e6ntN1etcsrWks6pXxsGp89oc1nwsU44wQ7rrZZYcbWt
Fagti+sFgKWEcdkPqzm/548dAAbD2kyYwiZYt3aYkgDTVY8XiAAXjllgOl7SpKK5u3NyHYIaU7Cd
aB2p19H7TlrUh6Y0NkdGEZGfmz1nfNstKM7qupVjQrv78l9oEbRdF2zX7syJah6KVeC5uudhVM3a
mCzrpQBtomxzjsXz6VfWsIG6BaYfj1ZojMzx4pxFNFPRLCRYwbrYgcdKtNae+LYuq98PlTmB+xbS
cs6kWyaPt6O2LGQELvPDsAu6Jm6yNEQHxiwE6pMO+a+5K/A/5uY3r1SGVH9vlL8FXvNHIO23xF4M
gkS2GGrZHRu5QaTvOkrbkkZyZx0t6txcJUkPPr1sSCRIF6Y2lmCcVfK2FxZwQh1XXZtorzjDhBYX
L/JwCor+yvxTAmd1aCKE2vINagWF71DCr47S5rfNRbF38JVh1eUQIX3sHTA4UIhr9XlqH90FsqWf
1RAlnIx3Q+DCjjoOdJFMVqFasWpQAE9E0zDPE6XQBqOc8fFVf/5l90L6OKEnGde485WsiAUW7Lnp
VRIaipJ618DDI9gzYQa8bTH2aoqL3glYMp6VWrd0u8lhfAuIRQZlNp2vz1PBJ3ThXSDX6JATCN0w
fjFLnIoYsbrNhZ8rwV4lpppHBcwpH3YgEInIUmCwAByaZQuWENhr06PVN7dryL8pk6pXI43KnSLi
7iCrJ3zA7j4uofQvjCX5YJTKkThMvOErBJ6EWr2fMaH+0l7ZSJpsigbO5vOb2LmBhRmQzttE7Pdy
Jfr9SfqcGYYe5WPRrC03UaXgPDhlrRtgimjrYGtCQxRzknWERMB1pQPJvgX4TVXCn3rJZNSIPPqU
Qp61/U5BM3FieZWFSEZRsBQBvelQjcq58AwEUnd7g60oE8IN5tDeTJ2BQvgvwNy/LZnz3+OqkhNS
oCb+pMXR1LgMB8OT2+ZheIk/WqCP2cmZiONzYtnMlOD1IyyqXiW3gNo3kGGJtRRQXQ9jTXvod7q4
IcfPQm7BCkpLVP0mozBNCHVoAp36Bqn56ycXIPxOZItkTBRWXHZNFL6yHoLOV1vFer9hLFpZgnV/
v+G0iCG1nApJT2OuE5plnuXl2ddDGCKxSufU1K7jp0AW5DfOcMf+t2otbk7RgqpxOt7F4el9tC1g
VkuFRSVk4pELd6295l1ZuXqyhzcKqKNycLSCCut/DFZAOLGWijCFOpiKXm42vNYOBzCl0QEwyl5J
f4R0npIuIZqBFhAhkRk30V6prUqbE/E8NLHMN6aaBKt+wxubSygsGNnnzzIK7k99NzHGlKKA2m7j
qrKduCUsE9Y++yxu4L7a8Ktti3a4isR2lGe7gF7IqneJhbM1wq7Yg/HT8uQ1/udgEvLO+Mm2JWQ7
D5Xf7lzcyb+/o0sfgeB6PPjyNJblC0FM/Mf+VyYfHFnIchDWYCWPGMg9hbooLZ2uzRjoHPh60SJk
MRNGaxFoOvoIaJURWTUjStwoihub+BJ2h6DUclvvOMPb0SNrZwduMlDNHjuJvH6dJYw9qTDW8xZV
re/0skSXwrVMPIfHLBFlK/TEhtSsGkg05eGQ0xPHdTvbrG6bhcI+P0lUw2H5FCr15vD3AzGTOce0
e2rvXEtwL9D9W9OnDQUKtHtVuHLAK0flRnVfIJnlhjiHAxyZDvKuJA+q1XOXFGQoUWqd6/HdyLxT
FgGNpKyAAm/p4YKvIMYmMLst6K5PrsLd5+RiELA7KHySwBehkWFUH6A70mwgEa2JOyrQRFXVQ1yi
K27I+ssyHjgm7qWuHgGPT2L0aoSRuERNw7/AGe7im/D0OPXVK2Odoo85Vf3No51aoDNwobe+oWj4
ZmxILetEVYPhWyaPuZ8YevCTBAmevRIaYLjpfEDy5cabtQ2lxveVWh7mbk1xJU9jYg2JeKVUX38t
ikQdrygTKvRysPwzS1xAM3ZTjUAbWGDGx09qx8N+DsEKsjk+uoJJYkp1tuJEQDCl5NT1aH/+fkyV
DWgmV/BTtbhR/JNF441yjupqlGXJOdXt136XM23Kn4h/+5sU0ozx+eOuoNuDTYbeDFyh5AqLtnc1
PX6xHIQEV5o7FTEh0Gbtcs54Q07pXMN0djU+0csQTPk0MK6tKQCupKu+/8GOeoDE/b6A3vJGH7fI
CDcalLfFSp7/tfJdE2qrQjsGnoutoRopTwGGjfcMQeaeV2EJSMBx+RV1w+X3tSsCSXYxsEu1UQWZ
OXxAS+3W8MEldzZI0R1E93rL1CgX+6Bg4sYBtzUnFZSiGkllCEXbA6ciLNGUTg9guqn3PaZSoKv3
nLm0hB3yhRJKAO8fgR+m4og4it/KwBhHqtQr18ara01VJJy0UQ/hzpIymUaZhVadSnfF1QyBSY5i
pTN3NT/agLR2IUzp3ynynqmuoXRornTwEMVh63hyhuzkGdj1GDzyHYAdh4EC7lSDujbqa2bHRwCx
oBFrAkVBZjr50EKmx3YolpPo4Nj9eEoLGYfMCMMx4MyN8DPuLHyrfHJ8aekYdyX1G7KEImF9lutD
IY3S919M+uDHsgsjN5VFx84kLZWdmzX8r+U5kZQYvP9/5fQsLeIF9oKat3dEKt0qAYP6p6FlYqge
SO91/Sr2FEc+rNv4HEFYukFWGJmkW1n9Kx+Xv1mvMgYpaUn7RjD4EYa4ovwxHmBHWODE2wUWTs7l
ZZFOc0NIyFDxiUnHBevNPV6ejf8YNqCRE+m0yY0m8ewpH6WC4zuhA1CKWBXeWMbtAg8JgVIrY2OR
pNZKt58j+NCERI4DbcZllGKPdJRt4AyfGCH2Y53gGadg/N2GYdjG00/uOjHq0LUYQEex97Y9Vbeh
B1vFyhHtx6BVf5hmQRWH9Mw+Huf1yRnO06RmEZea+xoLJA5LF/XXbTq+oJMhT+izjNW/IYy7rqdX
21rOv/LryfQOUI+RCno7iLU4JnzUcxVi/58bhmHgK9rlWy+68Bim8bwwuDDdWoK197JT5Dba2Zib
rkjaaxIINWyF8llGxHXKKpyi+Ciwvss/aM8tb3iZZElMOGrbV+tL7WZ6XH6HV9w1pFYlLcvoZyr8
W90DkPs5CM+dGVhRKxwa3lyOHrysLa9CzjTetzcdF7xfMGfjp9beMHdO8ONhsjGb2tanQ+l/Qsl6
lvy419GSgVAMqMgycmCl41bgZeJbYy98MPouu1ouGHis53+HnOASvlkN+Vbq05SA+PEiM+vsFaOQ
TEjTaH8w1he9YYtWWM0p24vyDv+9nDusIZoQ0NYhCLoj+3CSiwZ12NgVQQpAijKwSY2kY/2BgbH9
QiDt3O500Fjx9/p6iSvADdkoaj9tmbNGrHCiCotnpHEpw+HzU2O9tqGtBqqDBXoj/2djmJz7FPNE
hFnZJSGYhBkVIB3Q+QB57i9hbQcslXtzqR6NB0vvHfUkPo21tqM2JjrGs1txy8xjmbrya33gDrZO
Q5/Pz7n47hfxmuVjh2NdCE+nL1o2KFunurjQ/H5NR1WiqRi8tvycSdd7Y+Tn4E6UT1s5q+R7+7V0
q6OVesj0RSrsYPJlgarJP+GwGbkcJWiw5Pp8reZgS9RKo15lKkhBAn3lIf1GLkMPukLISei+vZh8
Q4w0M48ylgUEiOyI4uuUAAp8y/8XAN0czKK79R7xFQC9x9H5Hc3qjXIZGsXONCZKyiksvYZV1p+u
sr27FQjUUmrLKf9oBbrIxINzN+s9iPDMVDCSsVwAt8e2WDa7bXjUoeS1+XKGyuB+nxuHb9rOp9pQ
pWVvplO6z4oOks6nvyZnzzUkrc2XH0z6JW3B6mxwM1OwIJVVL5t5x2g1tyvnzwikdphEv+RMyL2L
dXMBvd+RHoaBOO1ykIZEJSwz66YA1Ek74EKFHVnMduGJGI9baxXwX/GgxUrvsyCGELIp6/Z9Av8e
9O3RPjS8qEDX7yyLvUq/pbs78UUvtF24oYzwYjIW3c2upcQ+fmY5zlrWS+lX6nlM4jnkb4wHUqSx
TmD9iil/AzcRTTEg6s93BEhm3gcR+n4App5e3Is3+jOIbvCaiaiPABYcWxy8eHVAgrX9EqTXiiT9
YYv75MVpCNWpUdQ3eHArrnqdCdC/v8IrwKa0HeWQ2shNK9kaFs8JzFghS1iLGRIQM1+a90hT/Mvc
hzeoIQ3uV0axQiDDtJ7eMH92gQYtrIKE38BN84Kd0xnpkMKHJHAds9hasJnI+11KQr8cE4bjMeXx
pwL17z1TqvT0LGvZuYfYUdVqY3UX5b8LNMnO5ja8yQzAXfY+7X7DHvCQVyUp93knAUyPTFqToRyZ
uriOVaLIC6KWepNoz+5RMWGYapu4oGzrnveHC2HZWT8GqBBQXFzag9kuxl2+ZaaKg5Vraymf2JUH
xGDNHYxtKxArjUiMMKFkdHx0zwfTCZ4R7IF0DQO1CcGOSgemyiS3xb7mO858aRDOGv3MDZOhYlp7
RnETYNl45BruWWfOUO8jmvS1WBDz55ZKBnzdKpizYAyMZLcywMBFs2ceMCIZyA76wjARw2053yZx
cvkbIqPpaOn3LKglpOecGm1aHTMMTU0aCnOsVsoHZjO22QAdTRfef4uxFPXz+nHLrp+4F8NoOLz+
Nz0amV9V4MCQYqXDuENosnlFheXMthc8iD/FN4UQ3i9XdM0u3GgS+56uNsSr1cB1w0bsXcHnfJXE
L8NeRVYsGY7hYDuada5g/NgYFHYQqdljPr/EECR7nz6BVoXTLC6E/XPEbzdReEW8VP+ktcy0QmQx
v5GNj73j531K/rwXVmCUtei8udCEOQZ6zn67CeBcEQIjqwBDKjOX+qlrg2T88LBTTdYceXTJg2YS
3O85NlHaw2ruQfIJ0V2y3sb1xh7OgpPNQmJR3HibYlJ13aJ/iSPYcziJ09kXzQslOTsY8bEDxagl
QZlJuWUrfynnWndZ+tXXWapZxJle4Nmv2Mn/UKHN5b7uJabf3zBJvyHY9BtVGc6e2fuyyYX9+1Tv
44w1MauH+rbg/LLf/FMtaPwPtyipzKe0QScRj1Ro9nvEl9ofsSqJnRXuTTR1CjwDI3uz+9N+qiLb
tKvnaC8S/mL2HiFjanHy1eTkPCqnlbzkvtRlpNsWSMavoPTSEKwG3OoN6EsW0odDAfAt4jWVMPX2
R3Ox6Ro57LWyWBcxisUyB0nBAOgqf6k+XlEUwdopz4xmssQvlsSVP+310nyP4qc9t8dEJ2V3kUUw
ngt7nTVURPJJvcRkdYKkak5S98F/ji6klDcDGfTB3MzD4/U5leQfepxAPxPX/60rlMheidSMlSD8
QlMVDbl5Dqy3D5WjkznWiWdbS5QjJvzWwQIEycrnRH2LDTHoT0STi54gOQAzKTG/Mc4By2MxuFqH
L+2JBApkrtG0BKbOZM5z8XcFECJ594MUnEIZ3yah9jJ9epr3Airdovw0Eu/y0QXb7+bbrTRXNHBG
bqfK9xAdDT/XjqIGgqCc+aiFeiFlzpa9bh6DmliFvKwKHhwRhU6eGC3mSEZbNvT0CCUn5kWLebF1
WKARTdTH6U69xsrrMyqVDABWQUJR+LgGWqSy1PnphTDY/YjUBhGbP4R9rFSEHERm/FfoDykcDfzC
XIZM5XeYdqfDpRSlGGeBHo6dDDUvs8l8jKeeNPFz7zVEqpN9oggN/zoz45kJ+QfXfUwDAjfc+N2w
T8IaaYlaCW58+139uXDvBHzHA7fiyXtMCAMFh6QwN1ejRiM10xP6Av2gtvVfIxpGKHLUFT2fcudk
cIDt+DKNWjau9K8xybYDOIaH4BvkqLWLZg7a+iAxoVhcBcEFT3cmwHzXBllHRtdMc5ESWVgRdWu5
N9Ein7i4jWcudjojHqV8qrIBuQ1C1ib/uO56oBOBDwth13uA5BU58AlLlZLtGbLhLGIO0CJFdw6o
Zmn9SCz5JpJXRPDxzOtzk4fTvgG75EbSMgFeeHiCyeX98RSLhW6CjhX3fr79JwXuv4I9n/fwV7Xn
wKh4tdTZOLah7rZ61FMYLOlPbeVCscRBurV619I2dLJChEi+vS0Q8vz+b+VonL8vwor30eTgx+0w
eQjDn/e75iGCoYg4Nd/KzQBDGtFgoAgqlWyAm6T+TDQUcnbJnTXSIrk3h6M/ebgSZkC4L3PD06B+
0E28yIhP4VI1ieU2RBh9uG2fjX6PQoCjkmR8R8J9a9v75I4svH7BuFkRwa5ppVQuIVnQ+yUVN5PS
gQB3N7plKiMv01KJxleeMdGRMSDDdxJw9Y3u0JnhG/gCyMmQaE6kk3wx5vLIS+AHcFuI4KyyNlFp
5JZJRb6Ks6WRLRjBndyAHWChVnFmR5E7Eu5LnnaPS+qvWBh8PxvpXQFGhollQ23+YbdGKBzeOuiR
gY900FtlCKafFG9iP7qCjphWXFylpj/pzYyp4xF+DY0ptin6cStovjd2guFFwLPPSlWdKzXZDEoK
LwzVb4r1uoEF8mK9MXnhJBif94r35oud5pKMK1/PL+BjkIeMPNOAQUBfwVQvawYJQkJJdGipQONe
KRFPSI88J4eYpPfo/qnzu3ToMa9j8Iy9jZyfCrXZ5atdw7R+9JLol98q+BkLWpfAfUcRO837wWRF
qHEsJBekoSuFCjMbWaDZ70wQX/27/SwDJg+NGtkTpy8Ce2VXyZjrVoLgOlvGOnkZENMrU8SzXacH
pQEk6yHXq2J0GK9zD/RBcGP3X5FuxBJct8fs8g+hXakqMNdoVWaQrJhaqbvOsTIUJ4AXQK8CzP3T
w0oM8cb5iN1tWoP6qckmX78yHelyKVcHHTCcFCeX0hzPB9o3C/zWE7Hpx367akU9H7bUOo45M8oE
aVOdlrANZDBoG5Fl/XOVFPsZQwg6v4yko9BLwTjC/+hlIcYCSSJEqVvE0PwKM0lPZmbgkIQetsSJ
OifN033MWnF80HsyuioQCb3HS65QpV4FauiJ8IoOWdHC5Ba3EgVrskfvTLbNq5vlKh/TmM7mepYP
mvqKO7MiGtHtlPpvb1jUUUG1kiYyRZzDnLafpgJHIbWwlV93dC5BEpP6Bu89CxA7QOHkwqegC6lI
MPpYzdQ6yycxCyAKX5imOIWwDoTiwV0VmIEGZiiTV9f4lwAch6jJyDHcVXeNVhfk3xTb39jTB8QP
XmVN5M1+vB/IQ8ta/3Vt0AFCz39BG8MrWEA5HSvAo9KL1VDyjdSxMtz/c5TdcmlectBNfgy8rl7b
EuymX07s+2h18eJXDYKBpzExU9IbyfPVExkbOC5eK3tIx5pUL38uux6hjVTidnU5W6qavsznlWrP
KMVxPTcQfXq8MKbEXMidiA1A/PGsIdnwnaQVqKDR/tQtrqbXjf2Dgf4OvkZApSvJS9WD/+foB3UH
CGgdutCmDh5ld3l/o8s+GBQ9l8Nofrx769nGcPeF7jK9zp8qkoGK7jc0wkgU0PygCli5H1wDmDFs
7Bxn3LieFuqJuGM5JLtNsSdw2gkCx1fcndLm8ter7lrN9CYlLD8c8u0V1j/bIn7Rvpr67Nogy4Iv
w4OhMrYHvjJhlrXsSGpxixb3lex5A2YzG6BUj3J32WOYtPH9Wid2UO4IbbgCbIWDNNIqdiP8dQHK
x7MPjIGm6PnZGJjpbPMTyUCAWiwQH960kcOvcaviJQrMWRsY/NzI9hf/doGIbIG+DCiOK9JFvN1j
iG7VgOFgw12obvhCTksKRPzEOuR0+1440+HUrYndbOm9LQtyXtWtxvb7G/rx/qUDIoASimFl6REr
gFM9Y3EkCXMjkxs9aW9PzlInxj5wv6Fvac85GF6TIv14f+xP8dbZZj/0v+8x8z5gn5TW4Om6H8Gg
aoVOO2niXBNHl9etxukXMeho7bHqv3cYV0TLoy68qF7kT1fdaFToJiXoEWcN4+EVj1r/Cq0zz2aq
pBJZ30/b3JBxqap2HiyWaZ841MYnqcIXNQFcFq7te6Fpm0ekAa7+e1PoA+JmIYA7BOd34+996GgG
xmtGg57ywv7FWsHwIWptXDJFLfQtl5XOpdHn+dsccy2BgXTrLSrVFNcGyuApH9P6Fa1emG7Fkqn1
np+BnLOS3+aXBI7B+72EggsUBPyby7RcUjR8fDaQ71wG2vl9AJHMV6z/be++e9GdUWqeDFhb405/
Q3ZXwvyZQ/GubtsO71FLvXt5BGJL19hkNbLLSJ9hTZ3B/JJmmz76ML+BjO1M5SKTlJfTrwNaCeAH
qb0D2PZ+GBAXSJuYZ8He3hHrwTcMmT2cMYFnSe4qNeCzPL0PztxCU/DUOhhJB4E8OwSYN4PAjohj
+uuVg8sEPiqYxqmUBaGEJZQ4qml+LWQND0LFWWqJlK65qVWBtfJWuD/sbO6ckPGouzjnPWewysWT
ewpkMpWISjFcE9SFJ/ouqlflp+SIGdXtvP5XarvS/OcT3ypLAs5hKbzMMdIa13pUyvRPL4nc5/Og
gLo2+2CgVZJnUUT9RU4bXryXkF2eUGNPlNMk1oSAyM4uRKkT8bQvCaGPWPpDitPZZXFJO5ngof3U
/T/Vrq0ACpIgPf+pyyKc37jc3bwk+GqhO9clIV2mymMOL4IbAqO/jGFSGKjfHbyfMMt7FcI9vuPq
d8+ZTV0Zm8pmFObOZu5yiFO/LQOSp06J+HKid5Qnl+xOpKVnOQQu6SFkM79KweJeeeYoQa1gQ/u8
bD+BOE7EM8kOUG7J8VZ/04ouF28V/DfhFpNQKUd0S9cYm6ixYdM0/QIm4CvyLbzHsa7aCwJawqoe
FiQ6mJ7C/+gOAzLFxlVuJc8vG2jKcGZOlVY2haQSwPsgsNOvUWxeiVugLoLPKm60amZ+BlFdiEsC
wqeOvIB3qpJhyxP0E9GP1bX6E6d/1uH6RYh57ukcRqVZ8l5C+IVyb9CnWcyh+2gi3GVQSno4Z8U3
LoaIpe41yBqvu0BdkN96x8CMMHGhzOPHZzUuOPhpLMAbHZOl8jF8VPQzXakvXERwlxzbndPuxZkU
CtdhML6FmjBdF3pslEqbrCcoImHVwTOqpZU02gB+TiByWwZWRGbSG8qRBQJ5dwvDoTw90DMIOsqz
QLioGw2wVAccvmF2l0e3Ox9O3PIN7pNvOlSArfos/57iSGMjPC9CtxCnZG4YYlTnpUhQVqCdHGQN
eBobgl0/QbwUrhaRI8l/2s66roZd4kmO/MDKJe/PSaIowWQA0YfbSolC1PloBr9QJg6iCtA/cqcM
y4uVqvNWRChZCmUZrFfsjHfQLowPvG2P1Bq8DnlyzpaIBsd4ymj1o2sa/otIgjgCbKhhseqp9ULi
XRBBF7uZXSmmAdFoIWmAJU+/2de4OlQUsu+PJWEtjdCzoBvyMobtsUGex7hmeSmhXedFd20JLGsv
ivV2FdpANEXgwnLcmEroy4PcvQU/8XdsjhUM5wBSW+ZHW5q5z+m9xdUcMzI6A0gsFiusAomOSLU7
9FIZ+dWTv6voPgYPBphHry20EGtxHtgE64gow+GCsLmQ1m6R3oW6pGbtAGeK3dAWPxp0j9WR9BTz
doKvN9TRoiVPgAKiTvjzY+N2VFb1Y+Jpd3J0mTB1daFiDGgYqeqEcW/65/whmLFV3Oh3gB1ZwNCc
xFS6XZ7+642AniFfyBhla9Z13jq5kSL6Wkmbl6znVSoCLbfJHan85bZB0uNudRdLEyLEBa/q4ImY
9Pv6LZptD6pKklN7Ns11iOv/lIr8YkEFux1TXvVTDn6PerKUBLzrtcvzhUTT7q8//DDKorhhm/ac
UAADInmW6rcmTh+BZCedVRFzg4qVmjDy7eLGmU4bX+Dy0Y8xZrzBOTLte77xir/GbWBpgUpeGhzD
bevMXzI4Kz8TSFoP1Cgqo395eb7s6C+NtQZ/7eNCu1HSKNGweuj3G5LDyNtPY0P5gW/5v/u/17sJ
nZxpPIeONTVCCzayyvnIDJY4xAfkpoRF9sluAknrG7aGKGDzfzrN/cLphPGNF3ZPqrMcFyyw894N
70v/zte4MJS8SfHs7MDNOAtZG4DfaU1EO1o2dKJoBDs/sBzPKLLcuK6V6vbJ3Dx2XRxH8wnTF9nE
X6Becbt0EQfdvvLQAOYlMPid/AtVFV6V2Eny538zEkXQzIV4S+pAGCb8XbZaHjWK5t9eCxiRXxct
oKJZMCPeGFvqBMBz61Pq1IOX6k//QAr7i7tLK1rZ+xfqF1K2uX+q+gFP/yhh5TNMslpvE60ZJ0jv
3vJTm/uyuCDgujMm9EOtDO7VLWMqjcCyWCVJXc4ZKH8WcbfVxggxk1bkN8qHrhHmQ1XSC8bUp07b
lbCrilw6j9TindgX0CCY2NjsaXfI7zr2TeOdZVtepNTTNrleRDTexyLma84TLSFPwtnzmoiSAjTu
OaSiMpXDm207u0g9fjnMSXc2AMuBLShTi5lLWel05T79anjvSda2Zoouh0Ghov6JI0iOSSoXY9yl
z4ZBCeRDcacssvHxRZvXrnEuNXTBDbK46MZlF1qQzaTN7f16RpGCeU+5iozMUKHoijVYhNXNofea
bXU1aNnbjtOCVJfVfalxoJMvaR+JHeOw4KWUG5tx9bg59OVuiXgcYoycaF7O3asj1/A4JTXF7ZRC
Dsm5VOV8oBBUaR/cX7lViwpNRy/bXkYVZ+EmoIQWMBoDBK+8N9JAOaSfOCRqASauojrBgxNFxKYa
rSGGNNvqD9vJQg0JQPXuBHrPjQyiw7vhIlRFTozn70pIKh5hV1JdFMe9b7NLADkSOX58fOmHZLYg
qeINkZR56gGA6Q5oIaxfLobGZ2IQtC3rXnbj8+gffzl43QWtNZpWE4uu3SdQK1KCS7W4Ho+rtCfh
l3LwPwgW7hdlG37xJVC68LdopSonKpChq0rL5I6rvlJueGFDQl7f8mBtm2qJZ0F+6guoeAlkyA55
8qvCYUEoc/fUn9MMx8v0wmTZwZF5WndpeqhO6lMym+b2k/5rNri9nHbgucssA1T/UsZBSYG4xRth
99jCgL6wjgadF6xWqWg1nEozibGrV5DNEYijy4DIi2wKJlHb4PL6OYA6PBpsRme6etQRqoRcFwXQ
9AErdYNZUFE7170SrzyoWoEThHzfKBL87SwTFYhTvUR2cay4glVHq2896b6I5pIXBduo26xK9iXQ
g4JqGK8kEs8P5vmlBc4rhsh+/tGzhErgvJIsflwON0zCOQaI4tnpQaX1NcLIjRFxk8ygW+R2rFYn
x/jqMkwvOHcIPYQ3AxRrxSxb8asH0d2/1JHXKcIY0ydv3rQAXXJrJY0xIwzSb6XPQpMJ5HyA7SFl
Pwi65uKN7XTlCmUjnCMpWu6ToLqAyeVTFFA9eGMtfrYc4OZO+shalhrlHb29U22XOiesg+n+L/Ly
olkPfcEpYbTp7uvHrk+6fra+cDbumRxir+fMK10UZoLSFjR40sg5fyEIVgmlMBe/vPTocKzfxmzY
c86xgUpmCYPpA6XGneC2rsLZ/gVc8loV/RV+DyZ/b9t9HG/64X5PSfwrD4kPJBsoVskyJm0WujnW
zRubNEgYELosP+Kogca/KkQ8LKqO63hVTifQ4IhZhyJjzyg2VsTHFnLu+e72tSsCvHTEe9bymdim
HUOL3HHNZFge7Yc781CxaNpr5ULCUGf7cejp9QfdikA/7BBWqToh1lTHLhdLDuByDn7SlMHZnJOe
QCbL1C37qb8y2bog2nD21Z5cSa/Come3LsmlLDUImFhSptvfknn4hsbRqAcM+MP7XbGibo2I73L3
tt2JvxZ9zdb+LjmBM0Wp1XhdO0aSHspPnNp3fWhTuNGeKz6BXrDgXuY5JI4GXbueT4K/3z9nFany
PIg2cCQf2TTVZOcbBNO+6NSl8ODf+aoYcnKhG326N4E+b5vUfNz/aQtS8dI7rVLQrfS0XSmHWXVG
npR+NSJ3FmCIy4J3OYURtrXQ76PV2kxEWdxdZTgrHc01cH+mzUF3uwwY3uXNrOF+YJMDqhsaHwYE
LeqrwUsvOh+n3et5JwUxMwtZviEV3DdNkhHIyMHqz+viQ3EqKsfctg2nJFawYLfttnZZmOQNUk0d
sn/4pQgO8oNFuNOVJ6gTVRLSa1sUP1O45c+efNf/Nm+vDc32TBj84ArvlxIVP9K9/B4pCpCn+QC3
OupylNAdPNFUKQjYEB2GHOn2kXfXKDKXjJmzFeuS4YO3BxKjVmMF37oEhhW0cq//HFUPaPBfOSpw
FbiiwF2FeEvAAkF2KkxFBcGmFKqC0OQmjOkluYK8W+wWKebUZWPmIcG+Mz/yYX80FcjiH/qg9aSc
boydVtinbyV0C12vus6auBXgaUgIvWQw5knRWDqAssIhcQaoJrabhdBcvnC56UnO5d6Ri4jwjTp5
our3PAVSAK/ox93oG6pAjLXrvQDLh1LZXp1W36o1vQHc/Pi38po1QHHD6G1it9N4MB3TXpuXJ3rZ
EmRLeW/pO7gjKqgrcdaux6YvRZ7TiZWFIHOGJLABk7u1OKTC3GYmmaqtnHSHdxffs/t5d7dBE4KD
MqCL2pqnu5qgt/w4s4pDlWSPhaCSArpp12DXYksXlDHy+mxal0bNrmL4xsHjYkJg/GQHDkKL0yaC
nYcSg0VFsV2WrSthjnLDHRrGPy835/sySMRYES4Tv9/1ZiiSbZc9W7MU+IvtyFpv8zHHmRm7i6c+
z6RdJqDyGLKCb6AYUi86wL53tD8LK9lqzdXaGzlOFBTNCsDagmEj8XeIyC6b5w1wFqdpwqzznpRD
/wN5l7GWBTmjnu64p8UQvMABpu2Kcksq4HiV3sZ86Y2wcESRZmikRWzhxAbnR45yRbEeecQFARGk
On4dWj5yo63IbecH5ZfbBHHpE3xX2Edps9TmPMtvFezqAJTiRP8J5/zjPlJKjr+ouMomA0S0wO9z
SMOAgflhoFSjoyo0nmCxAh44YtarHaVhC4eDurbHW7D+APeseVXKTBp2ncMSPyvc+uORzgt6Mphh
xxh2T51hRoWAS8JtbJE6Vn/YnGq3kA3O7ihdJhSYkEXiXOmYTy00SUWVk/bMRG8mA9NELNiPfEZR
NW1Z8tbpsHvVSurtcp2RQOpq9yVNHxj1XA0SwDHfCvjr83Dy2qyCx+B98UuqOnOQSod5OHObkfYn
ssrMAV7sHgMcnHqIDLKGpbhf1YiXtarJyjhSKUv76fislMm4fSN44eRKDK3cuw==
`pragma protect end_protected
