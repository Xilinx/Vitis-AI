`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47024)
`pragma protect data_block
giGA109OWTgnmloyaK8oODsiRC9RZVQFcgf9mR/obyjke8kkfwHUD0rFD2w6Qg5sKJtvAY8b/b0q
V+Sa+ZX24LFU4BuS1vxLWFGohu1WaQVSB9HQcsOWHML849yQr1UuXHS1H7VUn17v0E61+/PqUzk1
X19/pJmyYW1BM5ZHOhJulHdCd99vhdUA5znwgIeL+qkiU0sf11eCHljau90FYmDoD5m6woWzKvoP
6gHK4sf+uEu6z5A+3PvW9Z9m55mkt2a/UNoD0i4Gx2DEeOPjpkTsAXgRZkx7tNzlh61RWJtrXYVN
OimA5sPsUhnXl84NhviFAZiJ68QVQc+mO8WTYdtz61QdOU24xeJmT6K808rqFNEukbnTDDa9xHQN
c0tszEm2Xc4zLuPeXd/rqCdBdQrCbzr0uAWFMuZdt8znSrhBcCud8z5SlV8eGaZ/fQZq+9J8QHdw
zfgghBOi8mkbih/txS0fcFOe6RVKekMC6nemH5a5c+L/vqjCe03VXizNCtkeV6d03dlgJg6LFmsP
JczSfXQ7L9v3qr8VELRYRI7xz6TfWc3ECICBJA7ZaWnKDXUpClwkiGe5bocF/eZFyAAsvDhs9df7
YbSe2UM4N8jlVPXOkuxPtYzscpObgWvjyJuxNSOKna2th/8KghAi6IxRS0ijGNJVyQOCnT4Tzo5v
8qXI3Ydhf4/tCYDGni+CElqhQnYrxb4F3JgfmwVCxd3LVaVPBhyprdBRYnClefpGIwHYSiAKMEFL
hAqggBpcfNWZ3E4+ai4/HdovVk2gJPnm1drMm6BWBX2tm3QI0U4haI8SoQ8vLtWBKgUQepDLcC40
511oGQZtsyszFf4Pnne2vpiYO4q/+gInA1DaQkbdBCItiM23AgA3hgM9xq/0h4u3JVpSmUhACcXQ
EtfNsAXR16ekjbfW+X7KC+jhPgZJNl2MsvvNxyfm9MG2/FH4nnsvbuRFpeda5N4Jn1TbA3iYrHVl
sXnUl2VnaFoJA/P4cyBV5H1mQTdL2ojZC2rxQV3Qpurm9p1bgOQpa1gVEdnJp4UXfqHl7c5dCHjM
ksQVxVzTWL6Qvx2o2j8VYYOyoHcUO8iqIIL3hx57e+weSwRwN2EoOj/9EK4AjvZqb37oqRMQ4OwF
cWusLHXS6fzYvlDnrwX7PSUuPUoNEm0orUn10Lcr2oy5O+j67x+QkQPqx07Ttc7KGwZVagnwLZHT
ThzVEc1xpCBU0iS93QFt9kEMg3Oe2JkgpyO9NPdz0EQn71qbSwP3UpFCQYGQawxK4WWD5NDBJ6eg
Nyhs9zXY7CUD78WTe/uId6aX8jlxHrLjZyE4ZwS8XFsHRds7DlVli9z4X5Opah7TS77sxg/SlxcC
PNVReee7HCBcEdcuqgARSVA4k+pDJntGDLyr4oyCwjOtBvGtH/b58Xx/je+KXScNA/NnwSDVF+p1
JqPh6rTfTSbHOvtjM9AtFadjGx/2OHB67ZeMF80ZPIQ4fk+J9xcpkDK3BnP1tETc77nplBDkarSW
DoqZe4aTgWxkKZFJ4EmRh+sKya6VLEEywek4UIRR12LlCWRERKqDerqveJ98kcUkCFhE3p4I1ZPT
P4RLihfshD414EXw+8jUCJjNujVN0secfcVCVKKekLoakP7w4mH0Ynb3fDIHGyWWTJrrPjPZ+f07
FkrM20qbJq3LM1p6pl9vI1nG2tkzCGaMkdZjMO30Tr6qqxgWRRVUoZG7nG460BJqKv5TjU+QteF4
39BvKT74kNT5Et7EDY3zYQSCZuHMn0W/AEeUMdXxFEUvT9czkf5dPkIfRJByHARMDHZm02Ypndcv
0nM57c4Nt9ILvwQQ33AdEmU4ClkpI9KAFWjhVzDoysrgO36CWvlJSWDRZWJQslz6MQEfPlFfm0VF
91PArFgh/zPbA9fV2mx1clsymMeFIU9o7NYJmKLsnYO5Du6nDoAjgJrZiyUxyH2T0DIcJWB4h/1h
saoLN4j9NmMT2PMs4ebrabAe28n4q6f9SEyJdUfYnhCfIU2mKgaDGLU6Y8kNcchxspcBvAC10zr7
DYat1k31C4eeIBsTQBgptWzZthd2PkXzTPobfk1L+vAjVzTZGY34Z7WS6wAvZpzRHAbYfgk7JvBI
KtOXv+AkWNgPBP9DGXbSCCLmDwqaoG1nMPorpZLRS2NzswqeKwdd5vxpM9He/3Rk6w4YeIvmcGvE
ql9Sa6thlly4HfGRkT+rYH9ilj1NVhIFjXiMK2TAEA0dUYwInXK0hTnYGznhkGCXYR7F5Eb9ZeOI
lnsHedYNKhTNSMeNrocwtBaCptyZ9VWmS64QYq9amyj32+RVusCmkV89GF4LdspvmLkAwoIZUm3B
a4jvq3VkOM4mDPg8zOwEK1J9DUt9eDmsqGApuwPLTlSkb+6552VnINezK0d2JR42j12UDZh/OxeE
20ihRCBi8yxDm19u7NR6MoNG+4RBRUhwD09Uj+xmV6I1N0pBqiFOMgZfCylrU+PDPWaDwJSIYu8P
+KNYPtOGFn67hnRW9E6U0qRV9NilaZre8KZjgfITAxXaycSIFabSEVYkfyzIk/gZt+BhzIOg+NaL
RN0AZgMAxkLSG0IAeIOfdzT0IdjZ9f4tJRbnQlIIatiIyCH0BAf5NYbW03oEcCIAoBjKllTMcRFa
uV+Br7zYyAIXeU5MvODZzn6Yy42UrXvjbHW1F/alF8z0uBdyyGVcZRGOckAuDGWVE4Kv4h6bNTn5
SHe+Q8CLUM2451Rh0koGTYSXOZCD818AC+DOSTNCEs7kdl8QSGlYfv5mINZt1RJGTEDe4psgnC4J
DxSyipZgO/4z7lrNLJBiynKSE5GKj+7hWQi8VbkF6/OGLLQOI/UefGrhYRkFSUD+orbnsj1aDfTk
pnNR+ZUy9FwN35kM8wEkW5wz4AmLwbeNh0kiZeUQ2bwWz5cNT/wHgW6iRk79Cw2XLCn7XjN8qGUf
LW3pzXvVn18OC8k9qqF+DBNm5sKQKuZTNPb8193IWYLQEul6E7IJAL1Uz4YE5Oa8zncCJn4gNzFZ
RJM0ZCrzxLDEOPbhDDLYm+7qgOMNW9bSEe6zDLuKrVeBm7E0qkJfymCgpC+Z0Y28SUcDOxmG6gTz
IaBfTO+eYTZmxvK97qXMk1+NXKMzoqtsa3jMrIJVbZlGAwzt9aGpp7EXfXb48gxOhelvTFI7xDZa
nacGf7ybAbs0OBR4LtUmhC8ApJJE0lowqTK/RGFUegjNDG3MOs3nvYBunMCo/cZAlLGroFJpsEP0
wmvrbu4w1/c2Of9otpIZUHiqTriiKM0qJlNQHK2BsQUtCXAXePSnskukThYBALPr4uHjyRAd+U+t
iGPCw2Q9qN6eQutcsIbtCvc4t/RJhG4Lxx90A2Edi49v8n9zhBV+KeC+hgHq7j3uqDooNKMm8BQb
mM5ZCYBlKLaEqGcdxGOSKe+h2oMy0llmtHdJnhIfrDw8bPsoqMeA90Ycybq3xQdU4XmjuLedsZEq
eN3aXKPZsqRiol3SfVxFcApS10zH08uKEHwn0tBT9LB2rB+o6AersBcysZOvbHBqudFyGWUleRQE
nuys134N0exkISqKrJuw1tbX5+a9+z18GCJJD3800EdP9Nk3ywiyEIelBTTa4Vdz108lXr82Y7xs
nmkmJRv60CcSXk+4rED/Ot992d+h6o7NSzGtzh98uwwa8ejR/Ggpzb4iBtIzaJFjWsQIP7D5iBB9
lESHWSM7EFAV5Tj9otlWRvBjkWelKVGfbJgVuQVy//voHeLpFM06d3Ml1jChldUpiO1eFFysKPN8
zxuKbX0XKMGSQ39Fa5atfPxRNsWCH5iRNEWLp3ogyEtqgxAWH0hQqqhxh8O2Gde3Hl2bLwY+9neW
Vc9qBGioEJN9KNnjoGNbSArgezbJ+pEVIUHFTS22vNQrfQ2mtmNEtuPzFUoCV+C1i7AtTBu4xNKK
9neEVC0vNa39GKnzqtGFklCYxs6aGygXcnhRa6cbdaaXV5A3xWC+lN7k89hwjczpBArrUVSbUSgn
/R5XsRLHGCMO5qsiNw7V2OCxSZVTmUUUrUc2u0gFnbpPIi9yW6mPBL+nURN3viZCO2fFBU2kFHJK
n9IqosOB422UdnYJcOO54U7gi73jgY24252rvurZ4xsMzDJD8cE4AKG+WILoqASLE8vYABMffK3Q
2of2YgDhMLKFdVjKWKka8OcSBOjWn3Yftv7/Txz991pOVfxDw4/z2cvC53gc5fVQpQbKnOXQMEnG
H4LyWYypJ0f28LAoFX9tNIVOllXkgR+z9YzIMUFegjTQx3h/NMeWjlrY/70zsdOUEw0Cx0SYZ4Vi
VnwSw29ULJywI4z8dJuPrlM8pxzG4tcwMm8QthW7R/hFM3FaULf9QRYIHFsOOVwoJUUf7LsUuPVy
7mwrWKgKRaHKZ/8wUdJaP4QnF0l6i2FOgZIdCjb87Q0QLYhc5LMWDF4ZSHdKuopgP4Y30Ap+b/Ba
vRf1k3uDdfEAcQwWLaG1N6J5h0W/lzzQ3Fq8A0Y/HHxBnV3cL5Ey7fGkrtwlmasvRvCx01E1MoOk
xqgxHZvv7UikVVhrvmcNN/n8t8q1cOmbAQuvQP/njD2Fm0ZaHjXWImhdzJWWHJwErTnh/YknM7bJ
SNOmxadZOmAVSHH2I8+oMxCTe/i+oTDOYRh+GIQa0K13dDCOMcbhxheCIcEUV00Rncag4F9aLk7o
przH4+7Z2lwpJ3mlz2Z9A4vfodwiAmHibi/XcFYt+Y5pBFj2PtJLGdqHGa4u6s0Jt6z3z7oovRRl
utb89EK8MQt8vcFCKCbePWc1NkMONRCV9bwPnvyDR2j9fu5lCKYqSIN454IrESUEOixWBW1B/i+/
GiGcL4HAll/qxrrmlDwduFf/QjUuau2fcDX5evanqeOKHv+C/J6cdRmO5Os+8OzO+h4J4665Mb/S
DMY35t3MCPaHcy/BdNdbZUyk4MV0z053FXpPFaTIfwniq2UF1TqvGFVdkyOojYRNTawKILxQcyxl
jPb6hRYDfTw4X3wizMbFBFsZxJrzGhX2eSC3XPSSyn4LscFZMk/kWEkBuKNS0bJg0cliPk7fjCMk
cF5dbf/KHuF2jxvO4o5c07BTixF9cmkhHLgoYF/Uj2azZ0XzE2w3RxaWa2x38oNF6tl56cJLgZOS
vs4Rz/gzLhxaNVXYMIBhMdIIUPlSKyd+1w5YYEbVFDUsQSROFG9w7hFLvrqm8dHINRfloyzHjREb
pP7ER+G7OM6rvy9OpgOHugJw5teuQK+MdnbbH5l6XropGTd672BD6QcGMep68cafZUCGfVmD1eSY
xtMkJBolFF18quCpSq03ijkLZ+lsBLNVIn2Bjts01vJjNXg1rtdRmNC/0ujTJdA7smgP07ebC7q4
0IRn+yzdsksoM7MV8Vd5cHs/QOjylTfANxTzI7xZKtEvVCMyeAipk0fA5mDDreQJP6nxSBohIvkl
a9wtj2KyuoqTUm7ucib3SYOOhPIODBsxyS+L64fgQ0n0GemFUKmEHrQZNqc9L5eS7DMaNGA+tlBk
f+20JVlr/EVI/p53U5VvqFOL6i5UeRuKdsMxdcdxyaGcoPIzmnfOmqHlQ+dWgnkg0pDgeYcTX/Wv
2cQ3rquvy64eCOuVvR9ecy4oqQf+tqbg4KZHILiBRZ4vwxO7YSWj5UWYk2sL72WPpBtsS/QG1/fF
SZONOR61EMaMzY4n2GfuZdiTBOhuaDlOAMDFSONVPj31ePOXg9R3A/10buNXhuVsvj/8cxFVP5c8
mO6+pp0HB5BqXFF2weT+HAnCwt8kvbem1xYhlvgN56EHGzX67UVf3VdmwyAVl1kcFRXyrqetq8C2
mZ603EKfqNinqEJW0OU+9TAqL93G/TgubZF++afqU4/Y4A5jRikUKHLMoqMyJLdkb5WGykFlqa/M
0oIoOFO8loA2cF0BodBT3ZFIqeG5w0/mDrd0oJALtbF2isjlaybnSqHlbZ4hxSWNvwWc4TtnMdIV
8vpTYM5XMd1glpecJQgdw9ptFRKitHCIt1/YXhL8NGfS/DhqUbvajd0oeCwcWL4sP/r4f+0zd7Mu
D2qjwx6aG3+NOwgDPrxngiZ9wOmRXWkVlFSuBRFx9qd6lSaxnfYS2KsLigbZ0HsoOQ4iR4eu699E
2s6yHImBzT2vZRSizXlOqTqGBwyog0g3pM9y0uPNq53GIBAfVU1hJE6w3QWRYO4GwurvxgvnTK+a
18JR/NzeXCPA9mobJsEO6peML3e/6b1vBY2kbPb3/k+LfisLTNl0XEwQIJsGLSs6xlBVqFztVh0h
6rS45RGH8YNidx9qLZ3KccrYDfUAZ0D5R/o8vqDFc7xEimpVeuTpJKzgdlm5Fup62qVYwpCy6C2J
yGT1oDnNaaxDEan5d0hshPlrC/CWuoNCdaptcRJSQEzHgWl7UbGNCM8dcvZd68S38rCECDpAvJvd
EW6DolH4uH4JosChdzfLtCFrt5lx/O/b1hdMpNzQLpOp3m8+cTeEzz529+Z8bpWPjmWP1ZF1pNFL
ee/67UgGULE7+l3kN1thN+vhsGQFc1oMK7IRXKlqZwpVA1oGmcam5hw7qAN5e2kROpcHSf6FX10P
22/BvF6dcgrXkZ2QUerR4ENGph6g1jbMtv8gDxCa9GjtKxAFCp8iqbzoLPjklNw9cNYSN0jyWd4S
x4wpEFNDcIKxnaUxgCKMDk+nnwkBuF+ULc5ZFogw4HpCOTM0Cw0qw/llmRGvkJpKi2PfwZZpeFzW
bVEbXiBpipuDYiVM7dhfDSFEviBNhEUva9o6TnNqRIG6dYkkc+6ibpynh5COPU0cR/Bk6ry2QQCu
PA3xFD7zP+NLxvOXVit2WxpIW1n56/qKUwT93IyATho0oGYo0tIy0v/7iytZmKpuifhj4Fm0OQOq
8m+YchMaEfPYGt2aF+V4MmUjFlEZCB9/YjFvCTJ9BLJZ8lDbEtxd0Itag45KHgn97SUxkCrRfN+s
0X5icutEEhfmF9SOEP6kFJL2vpv2WSyIqifKS0VTI4fFNtTvEwiZ+kHrXD4cMSnOuuyEftZZEwbF
YQ8lPkMlSCRjDhJCpUwtY6oH3yLoX7vmy+EvYPNZmp2fKciDjBUWQan4ivGvx9SllVkq+aBNMIxg
Fv1AGp7X2yZdlZ96Qg01ajhU8PXSxNYXnvYzEfzlR7t5J/vjIka7+rBSBqtTt1pHU0Gvgb0wFDhj
Ae/v9Q/63wn2grdKADkmzYftN7Ag+1Ao2yKIF6RTJesuH0h8NVQG28jDlhWQDvOxt6N7n7iNRKKw
mV0A2w48tPEUe57hHTTDQK62YtV2tUjZUYxbkzv63dN636WiORWizI/y0Ic24Gy/pXj1nP821LOc
ysYJfDzZcycBR+M4enWkl7j0DnSO3gNdR8PG1KVj0S/3lcoGFQsBcGxNvP20u4zb07JnUdljGFP+
ym4T5H/mZgsL55y74PCrSw+8GUeToqTgo2GNfce9dDuBbwc0s98+28Bc4YXx6CH9J+eWu/Ff8rc/
F7URHWzUD6is+MZYrMr/kQl1MjinkpiBgKEnCQk9Im1oW4/+318MLB8losJQsO3jrKyX1EYxV9/N
VnZgyeMmBOvUR6gVOmU8C0ZuEfJnwvhIubJreqEUb9fzl+6GiTknhDcAA4u75vxBiCNaNGgmAG6t
tF0YvJY1XcfvgIhpGyMISXKV34hfc2b5/VjFSPXEfDXyb+Wcnatom0SOybGj74+WaHOny/Ffq/U0
0m4N4Muogc3+6gTSePPBYS6Ck6dRdXaQLQq9BiXteBmytypSp+Cxw5BsuZH+g/pAoXFUG3paz5jV
Ci2AXH60slqE8aPiHSb+hRYXmBpZnKWOustkbOON7eRrl55k9GmfQE2VDCYCP2tC5XAU7GCLi6WR
TV03KTfpR0Ieq5ikh6IMzA/ZsXukHjP9ZcdCk+g7fpL8gMg5kOQJ2ApaBxEiUocOJrv4jku7TNUQ
jj65uLtL467RwphC+A2wuF2xKQMktdJOsGmTALn4imFtq6QJdO8sgqyirQt2l/XHQW4fS3RDSxlE
jeFog6mFf33g8Oq9JGg91VSAQVSsrLLdzTIx8hy+GQo6pbykVeoAwme/nGIRAdrAzWLMo0XN6ESZ
nYlNmiKFt4EXHPefwHQR3YBxgaAB6XZHhDGwbMa/H/z+r9kkWmw+P4mJnsQZ3t0SosU0MEdIYYw8
tx6/b+fHpJz1kTv2uAqk8ShqLAWVcLQY8uabPVOKi94KG9h6r9TjSLmmXGBkHmyW1ZcqtDrgo0xP
LbeLuwaY2fF26vEQwgJ+aCLucoUZNtEEYidFmVwptWsqSO9tsGhppsJg4prk0fLW6Vo/5ak8xwp0
urYmaSRFpJD542VW0qLyothlAZAMiEe2TkFp6RScmwneCtx1xutKOueyXOMIzXjmz4pIPvAK/ub6
8+u7kGAqCqlgNwNh23waH9SkxoZP0UoBhmHmtsoPHn9tzHTOebMXpzHFFZcKKIcG4W30Q85cEUdf
HArMYHXT/SL1qyEqdDuJLewNWkUglUfo28g8hfPDiOtCnummc1Gml/vlDZF6k1BqX0SQ4duCHmRn
5bzUKNSY079U/NKp7/a42JAo+R5yTiVu+P+qweCUWK2OEZNeKi8j3i6xj4aGdVaH9XLA8N4h0yWa
WKR1DZkTWyGZdPuVE20VVi7va98g5NxHGXyVlsmh6fQ0OS4JnWWlThDsnevTAwW+OoWCOGjhuds3
oPBdMaz2WKh88A8ioXK8c0NQYYX11fnwsub6lS+qwZSrlFt+IXzzo4XV2NeRPvU3S0Be4M0ShoaL
dR8UIWhhx3NTMLO0v5olCbyP5MS8ubcAJ4gIJ8iGCM9OItykR1Y3abwS0dZ0n5oWSWLUPzl434gD
LCIb8tM3rE4cxHW5B6MQ5LZrTapM8P0QEeApcFsvcdrS1nXzmU6O2VpnpWrJf5mOmTwKI0hNCuiK
V/gytjdjFoMMHb9uuVrFHXT8hGcPi9eQA61E0dSDTqluZXW3M2U84xDkZySbI4jUYjFLSLzehtrA
nMoonoYRY5GCFClMakfCjTqjJew0ZmHdGf/Rsom7YMruJRdLR/UtQqYsIf1rnTeem7NoW8dZTlax
mLBgJxX7f0Ga4BlkvJHjxmjYnJ6p0YkT7aF89iqP6o/XK1wy8utD6/JbKv5TRA0vQD2R+5YWS5E0
gM+EaqLpTTAXgjicZGRdWWplYRsJiHdoD2I5sUge4Ny3SY7wMLH6kk6n6Bss0Pqsze9246EjheyV
+hu4L9UBl26MKa3PpJb6Fss8E7oj6fpufB548v96fgH0KX5bUQ/9Vk2urnF9jCJ4lT03cIYqKXWl
vg+DU6bqS4Ijw+FW4kFndcM65FOSnOO1vMbGzkf2KVlEUVgLp0fK8rMYoi0e/o3scx+romBFqFmy
6HBahCYapmXhQB3xs+XqpCp/a7wusFGYByiVzzOpJzEUcWF/Y2ettGMl9QYvTHwZpVKF0Mvp8H4M
J/J2kJp4Hp6E7fJUMQdOJ1bIlT4PElZAWGthcqGHEjO/Vw49mJVa3uWuXLACxzn6A9anA51j+uOQ
e4ryqGqeuyCFQxW9YpF8iFTzgdCmqNjipJ6F6DirC0gRwq9YlJm/N9dLDtwryJkf8k289MhJpPms
qg1Uf1fircnsWiwE7DtgHW4B3eYeKW6EsvXcEBG3cETPEM2RJtWHkTHXVmFD5N6Jy9lxjScXAnVJ
u+HsFvFHdgpja2WNEmodwRC47ZE/yUiIo+gQfytPVSNAGb6vRoOAQtZWfqi+quC2XHmsajTHcjQy
q7JopGTffQhJVTBBieZXkpbkwMcqyOyI5NNw6W6QrOxmJep/yn6TFmwtkpfLkVAflhrdPBseOnFk
DMK9fHB9fo4sJrtUc9sS43ZA7kmBoJT5BFv8+Ggp3s3GfZsnnHv5BHM33diLBn6iDDZeSyBqLHeB
1pI8sJ3Daop/CVsNKR/aFVU5Gj2QrRhNy5bqPmppDMZ+wlbirCtTro2usx22l92BH7DZo0sUAayz
xswVMd9OmCWJm+9+Pl2BXQ1RDSY9EByt0OXGD639x1uw7gKNe5BH1BLixXO2FCYokUDOiFt6cDAB
8ZDtOpcjkiIz5Q6b/Mbw1ADJN7UNYVo0yNO+swocyP17NWyNFccZNjvoOeQM29OtTLZ996hYqV+Q
mNuu85COil7KSURMJXA9mM51cgErtH8Ob1cDRK9MnR5zJTnBUAsWMrsn3HBoV2vikpKLs4PYG5BI
gnZNCZERFwuL2Cts2bbOTiRoi4aC3DllHbaNVQ8CTDH7Y1MIqaUR1OSGr+fqyC1Uhm+/pZmSxFHO
Dz+vHBjdBiTFE9c9pWw2HBbI0kgNH8z0CLsJ3Whzs3k6IQ/Imp360A567WepHw62UgYNVkzZV1Tf
z1WsnlZlFvIv6FqYGzNDxdGYOSMkWg1TnVnvi7+stjo62zs/e89xClJBGIChmICgvG1l4xNnxJMC
cvTKzn/xX0W5OSEsGP0Y+fdF0XldxCs67jxbI2ZcUhHYdHrxh11e/MmBqigDjRLOl+xq8fO7Qt1j
+w9P11eBXl/OffR/PfakJw2DWdq3JQkt5/hfd0rIuW67/siCKaYtWfnTxeB8O2DHuEqpPmVPeHSL
jgSaYRFX3B+JE8nvZR45kl3YT9MWxlnQmRdrBsHwaRTKxgFkPW6ThUeFUh3fOxCpRHtCxl11pT4w
/ErUaoq7rFC0HmFe7dTHbyMrUaq9Fy0XB82wNc85BgmqtjScRVaKTYoM0vyzG6uVFtawPGLbcJ7U
f5ZFYNolB//SgIHkQHh+uD63yocoXDI8pGWeZ3v0dUcEOgBIBMZVeDMJno6oI2HekERnUJuGxF9y
qVnN6hmL9iT6sSjx0lkddS+f3CmyQLJrL1OS/UT28bPYW4N83Ch14oz6Eq4UEl1be+9hb4scE4X/
moHB2LDeKkYbiI5FwleF7EypTlA6VrLy5H3NPLK/WgFPJs6b6g84bzd7bz2VSF54LLJ8psP+JfIT
9tkEjz+urjMgmx5atrC4VuIKI5pwtM7WcMAO0gm3jxAbj3D3M+88C5iQCqM8/piID0GVyZwzz550
ytiLzqGFs6YVK7GUISom7rLtOiAhkSHT0joppeKvdL4q7T8q0mCx6VF4aIRic0VEqaQvAz+ec8C3
QnnHiYXHyx5NHjhSKDSaX7rBZugTF//+kp5Y+uFym8xBj0q6WxLdkE1j/+YV31+9txY4RyKc2yU4
rWeIUB0s0peAqqSCxYi5aNn9hWS75UcpnG1zKy97xeffbLEKVVY0RF4BN1V5usSl+ufF98sGVXHN
hm3CbPTghdh3giBvrCP/d0Sa+koEsUK8s7mOsldMtiVOPDCvT6Ef2e5DXw3/EDLyYe49P1GUS1Uy
LqcbZAieE1pTUV8sKYW1rwNZyf3iPMaIYrbnLixjmWYj219K0NmNOAItCuVKMEY30znqEq+4G+wX
r+/2tCidqqGakxCWtam/Ywk3alp75OcWG9K1f1COAJMl+/6ZD8vNfvbzG9uWrfBPHuCUsz+o9lBm
ln+TYu3HE0FXKQ+kdeqN14hcoYwa7Zr9ElUalCPAKEQNqhymR/zpvGG7QyijuQdk0RRpMc2NoQAV
eETLUSpd7kSw8b3P5G60+ij1+tXdZ91AvZMHCY/ckNZdaCmiBKLTXm0541rq4MSH2zM26uNiFslO
G8rrmRzZ+oepyT3N+qfhKtEW3lii+DOi3MZrSjYMCTyZfcFBg8GPVufhmdkyY1UpTirahPqxfewB
8ZzyByMRAmqFb2oeZhVAwg98+NastORls9/nIsNG71E6qiA4AZAnhAPSNSIxjqrg/xpCmjOw7p8o
qAw9TQrZNaZBGctS8Pd4iMDoB7dhWUQIT/mR70Opnw7ubb1szXbeWkX1kyguSPcYB49kMVK8tfZb
FCWuQUiQ9dpK4RWazLP1lXIy5ZxrssdWTX08q1mKIoR6YfdS5TaLjnZQmi71TgDXX6v7OcOIHOXI
lzNb/WOV8+zb0rYCcO+euFZOc5O7BL9Th0yno17Wq8EqyBSwQdSlbob3ljmR0ZIfxocoyg7pka/9
NduBp2qeGOxtemAuL5OghiPUcYHZGVrlYVHcQIfQLBGDMSWBhn1VYKQSuEVql34Pkty1bi9JGXO6
jmhKlv3Ho1U5cB+YeJm4ecKxdTAYDNNEusdwmjTjQJml16EBQXIAmuzUD60fT9/979fXcFZwohDq
oRac5+4QONz8QFuOEjnGMokmXy4Q5ciel2I8/7Vx8meXwP3iSOfbMFlllIpiAgSDKPwk/fTXCUNB
/y237JH8BxVhmFG3DaASIR8gNhPE/9n4ZmI7tc+eG43DLIVX+aItJyXGNH3M97fk3Pvsoj7QS4CE
lkrC6vBJ1V2/4E3qBEs9EmCLNYtd2l0Clo1RfICzQbN3CuUoOv71oXY5F3a3tsaRpoK15VplLmtL
gmSufDKJOUAnJULh+jaciXT2+10uFHFSRLhNBhg/o+QeeJSMV09rhJXnNoC2eaOaZVrfJSTfxVW0
o1B7i+fs2B17WcTx+zk7QMyYurXSQN4QA+VGWTLZ2+bI4wet46aFEXE4lnHzCNF/+70dushpcG5M
cRXelKBAh+oftS8K/FjJg/4LfvbDADQXvR7FK2jUGtpOIHRNKLjPQzdPXa9BRvUsVOGkIaHb8iSR
ydRlWA1xozv/tKnwdTkSXaB3VYEYofylk17Bgh595l4L+SUT6HYqU6piBR4SVF1/xYuI1pPdRoIZ
fZBT5xdcbSk5zpTuIVNzQ3lr+h7rYHe3dlxOMkPojG6G4jsl9mz8qdwQZjMqKADWFHsJofmJhPS8
cbpSkrhvA7p/tjCvc07fGq9KynnNT6w/tk4tqhYdnmFkEUFzrJfO+C8vE6N2NSt0ySolYuz814s5
WcusXKxqmzDS8Jg9ES7WU6A9k/SaRFTD6mz76NaGEXARo/TEzdqdZ82IvVhZkkbbjh0c+CoUjYTI
Le7xppRUmRSUgSxdXsPmw3iAghawrsenqO8qKFREnMxIXEzS4gOYetgu6fHYWmmFLMdYThiRCWeP
4tSDvr38deiKRaglrEkh5PETcTrXLL9HEC6OitCLirqvYHTT+R/Br99IRtvvJx8MTaaXbwFBxwJf
Fr60A4vsd0Zz/5MaWIicsOIFrkOUKHju7fZNtf4xPoiKkZp7xQonBQ5KClN5vQSHFKXIXzX2tkzR
/5knm7wfsFmZ1qpwUTO0jnyNbWN8eevhbNTO7hqqWmLDqx5a03bOk1P5bm37VWOlfsLNwp7i1T8R
EkfnSVGVvV/77YvgDyBYWDINyMJHS6eACcuj3cwRjnZi7Qy/0BvDn2iZ7WGwyPhugiJZ4yRMJZbD
FC4rNWVs0XeM22821ZahniM2kt6SCV9HkF7n7bJUvz776WmbgMFsGsu+QSWvXX2HaIojMqH8HCqc
V2Lz33qaF7TRwHUzFRQgf/hX0txk8ZibWYc7ZYiJ3rc4oNDThsMAonE+4V0Y2/UANlGajPa4MSn6
Hr7hBXbvy0y768nEt3tFSMZ5iBsOOSCnrY1ORN2LXSvi6cb37c2Ui6/BXo0d8T3Mte5yxP84KZ3J
+XHbLpko8EvNZAEUIOa9NUz0n6+5Yc2HkCQkri0TecBZvQoDvUQ5Z1E+HQtcAwbPOZIxuTvC9n3H
cMkngW/ye2o5WUnlP6ZDtpbmUN+FcLLqTLAHG9yx/J9Jfum8WBG/upZS1dYzjHo6AIFRThdzL/aM
81r3eGwFKapFMy8giSVE1SqpFMCvPISWfaT2V9KEn9iXPEvecqXSh5VCTCxHh20tENp2G8NIVWZm
jsMGHw/x4cAemXHHOiCU/0DM0WfXm5eyxzbtIKa+3adAn2yutEoZoJIwOEq6vk7q/oyaAX8HWOQM
zfOYrV9cUs+B4nd/KMm4QPABk8SmDY6tkInCOvkma8pmrX/aKwO9QzxaR+Ssx2OZNPNhmBXid6wZ
oCDiAlX85akPZHRMD5jEhDRjqVvgieT0RtP3LcvvjWX3rVcvNlE77TmQpbjrzPnibV/xb97o/xLn
aQwDorTIcGHU8ai+5Q3IZLmJ/rNSegAxFO2xpe10TKoR7tHTLFyarld5H1cumqYOEPvaJoIZm3VX
ukukmh6f/l8KrjRFtc8DlsrIfU/bVKgNg6p0Lu/wpllUXt1ZwAxiEhI0wMEnQwBP5Kjfy+f5l8ue
wRBlDrcZB2TeQ6xS0ftT55SPDLM1ftQUfp3fRhz1OKYIenzeS3PHXwFjTIEpGwrpTG/vc53ZaFfc
84fD74Q4pVqjI2tuozvOuMimE7qkO/j7HxZgvgpAt82K4twJvRbgVkKote4pHeb8u/h07xDEF7b7
xrX+UkzpeIHytQD6V9cl1kCntRWV74wqgk1DCaz+vxppZtB8Jk/i7Eg55MwD4Mok7HkcC0xtShmd
NMxt0ZULCHG2EYsUJyYhlG6lj6qgmErhPCwmCFHuMIxQTYykEvXp/hW/kB/CsKhKY69qzh0aektL
ksovCynuaBBEDi+w+2cG2etqeQKYKnOUvnKDs0/KfSArDDNGdQw3Bq6NE5MZ5sjiyGhFeTjHN5UN
x3H5bIMswOxXKejrnilPniRKbujOu0tl8jmHnYlW1feMfGrdlN4mY6CEACvjIahtUiS1E7F/LjR9
rbQhUn6n3DEjvsFrJLVwVpiS6iy0v55O3HV5LwvsfpuHOzStPI3BSbs491BfYzinz0ulzyeLUY9r
ubJR9Iu1M5caIOeSof5v6EqNwKLEMVXctS5tj5qtqWqAwJIXzdLV1QA9Yc4yMld8rsFgEjMJV+Hs
2p/OFvfOrkVoUHBossaqXqrdYV5T7oYjPTNTFHcJpDx5FEZDa1mlzKbFurlA4PWpFiCZI5NprGg9
QAG9K9QzxF3nQKWdjOob+Ne6w6z60LXy2hL7s6GizIPfEM4cf85AcwyjaznATp0tf9p1renIq+4B
D0C32tB22yz61Z/V457MSf7mnYYMPgVNmb7uinUrCnfpYlsAFHVLFWwTsTgJEuKQr+zfHI6gDySl
mwYETkHuCHGuKs4Ak5qiRCgfqBwBnTBi2Xtg6Ye3A9s+D5izwdXn8LC8D1vOnEVS/TUImbLlo1EJ
YWucjenCe4Pjch8ZBMZi8XiL2IM8sY9VCmw2kqCSx/uHWW1voGOyv4jtCwdl6ZUXwE+CfUTpOaJ8
mUuiMM91PPe7c08oRZRp6H/2oPrsvkV4vksM8ZlksJGC+uZw10jeUhoqFYcB1pG74yc6FP5XnS4F
2Wybs5E4E1liQTlESy9T5t3ca0HUndSGC0D5E1Y8Rr+Ta8gcvPsDzELEacaQxmtj6clr22FfwyRs
tDZ0ZTZg1nxkXMCjk02kfTeRQN2ybDIB9dofr6Luev9zoIFE9UmLGWemH1kj8UwSKWToDuqVp7EM
ix2EyZfi/h4xgHQKdNUkkF9B8Gzpaa69zSAPhLeaokaGkm6lHjeG/zFugXeee9uAN/RUSIgh6cKf
+z75S9g/X4wY+4pNQr//1o42Pv2uQDqVS9kx8yNDPaTOmwk96F0n2be/d7JM9mtWA/W9rL610EBL
omWAZt2AV37GomwLgMNKnmeOqXkTkH/HVTgGM4VW3CVscWf7CXhc3nyx/U96eUzo9s8JdYUu2WQd
nOwHxg693as1QrE9COI6L+78vhmLJ9dmwO4CIhs7xl8z9LOwKiBUcepbRDP8Duct4wxEJ+2VKvYl
waLY8HeOyapY/3Al0Mq8FsrMI7PaJw/Joa6BfMfSgdD7WSckur7FVrt0KqEjRiRHBu+mJsN5MXBC
d65L5MuzEOzVHUpUV6i0sA+XxSWmnq0uTnHYq/obGp23PrAz14rkL7vJm8WS1Th3DNF5v/tNsOpf
fuqIxYmMtSXjE45oHRds0wn1s3BE5PqsJl0IHgOcTmE3SwaFU/UxVlC/5HQm27bTCaHL11xGOstF
4RrSY6GAgFtHb7Tngkv158WvPzQmyMsXmR120rkAP/a7ZMQtXZlyHDTpxkOuyBOrpJfQP8/IFGwj
9GFzngEo5SM5zdSAsshthfaVLywBy7cth0FGMzkXxGN/Cy+/nSzRw68/xX6UCnm51539EbxT0ggJ
ss0VWVv6xXWvMRMV7RHa3Q7KzVUlq44DSZ/XAhxZtdYI1SjmagyRFim/FdVb7T8+MYjV2FOaBRIa
kK3A6Wb+50o5OoK5adcVg+RcNVG9RVyo5Kt7rbiAJ0i53DoUapbIXio4sD9d9Bbr1JkUz6A1CPXx
dVxKl9vw9MToHSYmJ11Dh/08nmeoSwEOz9aOs8+HCHJIeiVOjy1SHTQftWEaWOKlWkVzZcwTwLvH
vL9UwG6rceNzuiOZkLj9QtRjZb45WiuuBf881fmAEi/SwBZy8CVHemESpLNQgDRsy+Gel3ue3hwt
IzJehpzAYwAEHabwTPWzwPyY+NvqT6YJVZjoVJ0MV3y25iVrHzk1/h7Rr1aHQr9wTiLsdYH0S3BL
CoVEq768iU43o8PRYmDp/gKkB8ES2abWrhK1c3hN+JNkJ6E04XXniw65gSrC0EXCfM1jb7PD49Vn
NIiXG2XVQ8XoL7+qQcwuT0D0xGV+iQZgiPnPJM36BEz4M6sr92r3eDXJ4E+9GpF8CCv9LcBabaln
S7/ffJgZXVO4fA7HTShaCW277f0S5/iRM8gqtAQdO3P6lAkteq7VCYhZ7Rfctn5KpquhPf/7rlqo
C/+MzfNZehc9s0jin0j84I7TL3bFxTKozdZxKmgxb00qibckpM1MamLk+7F0tX5lUsEeBxh2Q9yK
KKQqDR4qgrSSESATUuuvSHZQTB1HhA5dRj1t//l/Ow6bY7q4HS9V873tIKE06iKNHZNa2+GcCalC
g1rpuM9WMnANO6U4WcCTqw+U8SueoYBnYbpEmIbIUDd60PBTYAv9wd9bjwIWpjUf7mA+LJnywCxH
HxaWC4PBSsub/1cx0ffFRgc+HYTDOQbjxTdes3WvnikalnzcWDvpQOcKmevY4fJLZCjBtnI4Ooka
f3S4MTq0vetIjyNnDtA5p37o5+/HFgt0vcEGJufEDfrlvAeeXHy7keLx/ZP0JpVq1y4ljgpKV37H
eLeqeHhVEKmod5/bs961o6I3mZhaQcwHBcdpBOdLs36i8uR42FkzFEna3zKNP8LalXPcOQNoISGM
7qljGNhdbdN4VfypcOcs8xK4NMaBSGscnQ8M9rokB+v/9rdtC3RUQxwXUhuR6r13Q8BsO/E3djRa
5/AnXFULGU7AhbpxEP9e7MJff55/Y34RtQrBzBdOzeuKchv1/rvIf+QHZCaNfZJSF+QvH/achiVo
YOdGjFOpD+USNh0RoTapRsXWHO1ACRKHPSwAC15Tiz6FCHgJGWJws+2LISUB14M46KNj6fFqS2oY
jV3RCKmWrXewOmay2Ej6go0uTOXsa59J6dyuZoQmgGp4DpJHhTLCtBGY1t8kM5QoBCpY8ElUDOiK
M8Sjfi+HKZrZRL6YORziyYKD9rIsL08rhZzafc82vBCPOkAxBVQoA7CdgsIPO2FCBU0ekhcD4Elj
IIB/YmKyD3sPCB4u9M7q7GpO0t7JhWk9IB8qfK8OfhIaPrYa1jvKOxLuh3ZWO2OH3FnY2ILLHGw9
RR7CaCeca44vmpXIXXYBITUv3woXoCnhj1ARWPlkic9QidIxdA2zG/wD6D7qJdcu4NeV7Sr3H99X
nCOGeZIaIDP+/kdiZg51xzHLnmdKO0YEc1cdSIbrSDWurapggJi6jdVlETZs3RXfYQ0NLNoJ83db
nsZmpP1i34oR8V6y6xJXLEhigF9t9gqIS9FRWm00XZMMKk+7kseyAqJsV/3FMgtglqXhyv7HvKGP
zkt3d5bPRwad0ZBDUbZpcI0qznOasElHHnVf/7o2Bq/rSBRENw0FG4IgH3rUD9mBpY6Lg0Q6a/a8
oF3P5H16+uqIQFtXfCXO0tS9bKBdm1XN5Pgqeofk675dOP36ZBVp5Q8jfEopppV/3P20VhAesL/X
0+yvzsDBsAYMSf2xhWcMS11JZUbkzCdsf++UGwXTbsIWY9ozOoVcIOcZDLfOOuUB3D0pjcO3Q0Ea
g6j7sCupO4Vmg6OLC4i2dGMn0vwKpHomePfoABFx8+F45KFxh/0uGtMy3K2V0mwz+JNs3tfofJLA
LoSojH1G49IiAwvcSfsVeBqH4CyVilLK+POi2TB1YZieaYUDB1dXw0Z7TqBkdlG6nhSWaB345RaM
Qkq2XC6lDEtVGp4qpMkCsNXaJVZqfLb/yqBp5sOIZpfbYdd7ma3a0uyio5C2DYpE6rL7O5AyoFgr
AT9dpNyytw+hkDuHmVT6auZcviUraPyUTTZwwWWscn+tPYMrXOqE6CsNnn1PE7hmg1NJjr4PAVaK
mMA1C05tj7sIz6hyP/AJs4VSFIi0sRCCOD6v5dQUlunOCRn90YhKnOl7zv6vQnbMAcceUSDTcHHJ
Ur/TJhVPcBHzXKFvF07AZMgRkhfhdMvvM+aDnlBTr8O2ZtCJrWRisn2B597jBYO4uROYw2/hJ6ET
uMk76x9Cgoqaw9rglFdclsNhFc7e1cg3z9N46hyn6GBRuwQQShgQXV/1KptgFopyBVcCmiXuKUBR
AW65BHBAtJOiAVE+z0YZ81e+8IwrG9jgqDcJ7IovGeUZmlrPvj6LEbEMvX5mr7QA/RsiBxq1bQfx
kpZbGTKSTwv6SycZMuta5e4yONlKFPG/yyzj4WhFXf63bHs9L3cZfMIAQhbjw7BcEdxcp+c7TAfx
wdFEDatIanG8tAvbgZK6Dls149nw8BhFpSzRI/vMeDEEspSe9ft9FoCFCm3niEh8fcid5h3vQBjE
bVdCI78yVCXCdWy6UYsFhZ9PsQcL1swZuBrfEVLJhmtwJhsDg77ecCXXTSE4ldsygyxYiMdY45gS
msOOAJcrgrn33CqILqVHDstnqNBqpzm5oluqwMR/5IHUrLij6m8vtH1hiDg1IEeVnOCil5LVdLvl
IzfvpgzB0f8TiGR+J01tvcVOPJmhvt2PgzaY603WuoaqcoosX8RQJGPQD8fvXlxeNIiNXhDHuRz7
oSv3njh5Na/SgZX+sCYHXlGqEgXVf4xwzgiYd7F7X56PfYt7Ut8ESL9oshcUblGZ296hkIa7O/1Z
Vy7fD57TT0NVp8H9pzs6QnehtIObwQVUFqkJ4+UJlwYsFvZZEvzzFTBAP9royQcPKQYLDoWYumUY
W3G+xPJ+WV3id2+tNlFCxvmtlyq2EUVmnLMsYdjllqAXIgiINiLIUTlPlRFNZOW3GnwrmT/ulZvC
wUzSuXAupXgfiCJ69cuk/p/q2+uQ1h02Mntdewkqn4Pktob+c18oUR57HJboFHSiTGVP5LfcKHEF
NaF6ElWeTUeQhMmIJpgzVIHei42VyrLnPpeYSh9iQL9TgAVmk8v7mTrhiTy/P1Z89pb21HAVVuR5
gSPMslPRYHumqjtEbK4qUxjSmSil9NGUcNMm8uZflboCC6uVfaufV0M0lC3m6YHrnFF18IISu9UY
FJJbUDbmzSRrHEfS+h4pEpRnQ8ZjZvvCGVbHPUfaCP3TFFZcU7++/sVBusQr9kKgXreQnMNo3oIy
PBbi/q2Ej4vb4hfji8E5qolOj2e7jUEDUR90dPgDJTj/1W7+OaYUQVnwrpb+hQrIt+efEYyzV7IL
exDFj1AvlJA0l9gch7IZ2Z+q7wpyWRJ1qSzv1Bg9N4D4qQewwMN7HfAl4tukK14Whv5z7qvwQ1BU
xh7k6PZ8tVkm3GQ5NJ0g1KrBEedeeypACISBx4vMtX3WKbVqIZO0LCmze8hb2OZnIsEC6+0P2Oli
sXn1tz2GWaLzk/shx56OcKhMqast/iR2JD9E5lOSH4RfUBqPn02032KbtMdmpbdJRU0ihu/2tqOG
eVhV4W+EwHE8tD3JuW3a0aiUs6ldmUrUsv8QpGnSwAuJXEn3k9TGOcWhp1xS4DNGLomQ7la+2ZQN
YPUlTRIflXtauY2UclDyceVhbYhSO4SY8HXm/HhpQomZXlFlOxJTRodxwylz2CMWSietAn6NL7Uz
vZd4tvXTZPJHyNG5aT4cualSZcFSBco4VmA01eSBABYmAffuGaw95x4SOdqHKho59MSk+tG6FQr1
7+dS2f7t/DAL37VPDvxA2bYiNkGi80E4bYuIm3La8S58NlG9yXGbjZG8XxVB2G+RhKb2lWStIzYY
Z54Ur5XeRd7rqCKVlFlZKS7e64Rm9xyIfC9UkHbhQidThrJqYbCcdN1cBCDUjNStKAopGcA8Hgz7
CaYK4BTIjyi7Wl+eKiFKRCzrwRteGFpZIVJ+2SzssbdWW12Rc5xLTDWgSa7NrEgWqKr2M6ySb+lN
Of4bK7gmRQNEEeQVUK7ik2yFyZYsKSVYmZIdFmBg7nLJ0Sj7V5q9+o7CjgyE4hnW9W4NyXa8OOmm
I9PBUhlGne0akwFHcesG76qJgq2vTCnU6eLJMfhWAmUdsleBr9/VKQNzr3ukz/adxsetwPYI8cvd
kkITwlH6bkMuvOfPkSSSHkhs90cDsuAQCGmiC2FpItFqwBoJT3RzkT5mbXEZq4CEM3j9He3d281t
DUppHP+YH0L9oL7nMOA/cTkC+yojXkfnMknnRU3YYzyl+Rks+W4Qv8qCioP9P7k1RbJOi5pLT7b3
LH2TghgOWq/z8r31bGTCoYHrr9diMLqzS7Y38lHn6LfWAE+q/6rDr/McQYg1z2C1hR94guX9yHsu
iD09g/Eumr4wfhfMqLTy/vGGdtELMniA/Ez1X7CxwvAKnU/E/68A7IFW4KxFNDmdxXOuABEI4Gbb
vHTnLlzn2CfULdtX4J4Z8McD6RU4CRrW/+YL6Qh1iGo8PxW4zEd8K5Gb0Pq7NhG+RqVNWOo3nzGt
R7lYViPaQurAzYNjw4rmUFUFM1gWAtNiz9SxKMsndd1eHJQ5JmR9O5Bu8CZowXaGaKmuW80OZYXt
EcvBUWVVVO83mk5vPXCTremUTWzQymqEBpT4SdhYKxcAU0HpoboyxbCM1D82YBTVAT9TttAAnNN6
32sh/jLmvD1GKc3WdPFefULqm7YsF2o7Gqg30AfoOfERfwC+KCd1x8NrpYkljHQV2+bLsPNYyBNi
KRekNDnSbLZxNOM/26DrXuv97H9tazQh61Rio3+riOeKkw3EGZZe469bpq9fKk1q9HWVdBXULOfm
g+3Thrz0ZVQbC7KcsfnIMf8l9uye7uMyvkmSlPiJIuEjSGLieT9y+GOKKQbFkxiQ+16wtycJ2dJO
3d1cTCKioYrA1uzz9uIaB2LwRslH0moqtfu3ng8vH+jHkfYzm+eL66rOglVTEwUXRDXxB8zWWhXJ
M3P/qlKnkZWCK4k90HanNuvrGr4XXK3i6ZVL5kLsfe12xmfqLf9r6MB8Fho5uhcRnCG7SC5Y9M7Z
2T0GAXNJdW2CCRlIEZeCmubDaZJTau9v3ZotcNE9/vzj4VotKdCkkeUvKhrimREAu1R292V/BlZM
73UbxznHLCMQfHbdq+4+Yug7eIeWRVwVVBiG9ubPml5DD++W9ZTymed4HNs1oyYAcQgZOjC1UNnS
WM7yZYEIKYu4ZwbEMACnRGlo/1+ShbyPRZXybZOHeE+i5tpewiRXr9fKaBNy1Rjys5QtWNL1BzSm
vJNFM9BgO7FYLZj4Jf6evaQMn+MCnuQ5artvpxrwWTI+3XZAwHanxhYH61Iycr9TIwGBqDkupLFj
fyDb62env2JxMCQcXQVWe6J4LiFYkDw7MZhLQtvGlVgGC8jnAMzMRlSQGS5iJzcWZp6wi+bLk6gf
VeGsb4Vslp5TmEq5NMiC1scEt+hluBwaUH/cyxf62g4oIQy1222XHJC7VEK5gEAaVoqnSVbyPA/9
8gkM2Vk0l93DRHwcBuNylzMeWrECo6x0dFu1jncR1OjTLwYa0mv30M2gFL9a6mCWssGUc/AJM6Y/
RsD6Sbh/GI7/VM0td63iDcXhRSx/18MUxHmH7Q7IVPEMUpDAs7POyeBsioRIkQe9S6v1ddyZARFg
ES+cVvYCN5DhIG2pDpOQ2cU6hO2JavzfG7C6qFHRlwdbQjE3xpTFQETTxtlPy6EXLDs/uQ/zBmNv
bzaVdzfxTZh/o59EAwnlBrTC25bzoXSLGgRIXgWFs96cU9EZj4b0hH1WgCB+3VgBfPCWLshSOvIm
bS+MYP7cLGOs0mWzvvmO54DFqp594bLOfdU0OHm5RF1isAaGAmCq/eYBGwhA0QNcALMcgFIX8s2I
s7ZEa+xUM15pVs2Y1YPBIVYtJC+HXR4fz/IeN70PTgcnri7a0yKcwxomHKG6gZmVi6ohgBgMaeD4
MnTCQDKZNkMqf/+STybTdFTLAOku8UvbWmwTK8tl/tb0ARhGygZRgpcy3uk7cOJDqCCaTvy1PxCV
nP0ZiXL7u3u3AF50fvh0BWCRy8TFP6+7V3bGcaoG95M1ENjJH7GMJA5ZwDJQAlG3ei3dydSYSD/C
gk0YTus0vA2VM8bRv6z4COW9NKlBp7MT9VLjHsPbOMYAzfumCpQLX0SKra/6cWvg7vdLCYSVDIIK
Gyn+SUvORgWyXS3LCHcC99o36cjX4HBDKN5gwe1/63Fp6j/SeUNnDLwU2EdiNQIbGZ6PuM6YYriS
nePQw6dyJcZQloEVqbfRvDaeBH0PXKcplqSz+xN2DsmaY4J5cCgyn03FVHURGtqnK3m4T/3ZJN52
YrXmu6P215LPDnKOATEdqGfe5e0VWvRh7ACLywJFBSBlUmPiNtVTh/XPcmD1Hbt3R+DybfDrNruV
8++edumnHbbyMAQB1BE108/QUnE0+mC6Dc5Q+/LbOcmqxYmp5pdruw0Tjx3m03N30Iptr5tQx5Wq
AC/4I/JJ2nYpIKKv6AKL3q+J2/ce3tdR0dkLwyqc81hJqtP/0NtRCXXJicYIsCYhsF1Egir8F8vS
rS+ZMksl9TBIs27Hl93/fm2qkJUF9E3rr3SrSwdbSoNCkpSbyRNWd4ICGLfuBL/SCXTU+4A+W1bC
BGDtsd0PEu1U3eaABPLKtXCr3ZsE14nioithRStyh+blIpPG3nj/FV8QZY6s0siQkxalWs57vsdu
qC8O32FaWktz9t2U286m63sNh3L6eVeQXOa9eXsXd3vAI1O936nWx8j0x7FO7KrhEmKnGpWqi3WQ
Kj+2PFb90pjfKQIB9nzu05ee6Q/pw2Fede4Kxf9Bf5iX8DRkAzyl6/etyKwCN6UZEBiI2e+2ayLi
aIu6mZdZoTV8yKUfnmwmzpPoyOPKR7A3up18hyaemWKw2oD2W9Z+fDRbMFR+i2HXJeV2E9hWF1PW
IjkG/oVsfmXcnboqiuN4g7ZvRZPHrkzE9ihUlgYdyI0c59/Ffq8DB+NdfuUG294oqU0tdBDa5FRz
zj6TLH3BvHoTUw/UKC0XEey4sYhmZdi+aV4JirRwBtFAGegLOukJXv55gxMvpL4WyTKuHorc35aV
DGpcbe6X28TENvOOzmBuhkv49qKNDNQFWjtyE93kcEEylEVia0i9vlCNW2IMzSGvD+45QY8nsVPD
DrK4UhbIqpFso8nlZB0rivR/RzjFRaKPmQ6bO9CWgyQnaTpvw74t7XF4nrecbmppGnUXZrmvAHNv
qLGrDQI0+kpl1acw/OkBNkqMrJxyMVzlUnFzVS3tlvezyQiqEeudV0R62wafb3tkv5SuK2X9GBEq
8wk0cOojWvl5BWGldWIehYAD51TioRSvs7nfAxDQlOIGzQaUIIIK1WaYEwX3EkaLFw/vT92Shf8x
cC4t6TVz9z74KA15UVaVnXaKVevnbidUvXCkfCJME7WCKYHA972tzKG20YpT+88xsaCC7ihDxa+4
9x1T3z9uKGEgRZcu+XMUhvFPiciS2Itc1MB+vEbrvluBQWH4XzVZd0Zju+5OMHpHmt7n8BqKwJTb
yXOC4N4dblgJwjkYRSwaKtCsq/QEELK6vYM3vRjkKnpDXdLqMYllOC7XzN5UWN9p2P+yKXLVV8Ax
l/xkvd++aKVDM36PIe5wHkUPxeJ9LOt7b6aUY1qhnqwiy391/aoY2MZ4q2rOKNwodCmOLhI+Ig3F
WClKckOlYXOujtCyhOn4+VwgXpVQOQTDGw4Xi0cJR+yuJvk1lJ9qNavG0fQgU5I2Xn+/yHu/t5gD
tZOZa3cHBL/h7AjXXbCZiL1pyRZVGh7I4azUJTTTVmznhVd5f4R7lKZtDaVPhQZGgpi1jPSuj9Oc
8ZxfWy/KtKO0R+/Yb2xIu1TUOcwPnZQ9gXnyDKbxwh0VtrcGEWA/Qfx3BYN3p1vIJZMHIzwXl+5g
0Wt9zH6rw6+eyyY/AhOEyMra1fUDgz2HWaBL4Mo6xSvu6avxyog32Ro7wTq6WvYfdg4n1y+UWNhs
Zk6SUsCJdF5vLF1oqtIxwTycvY+HK3RHjXWn0N5YyQmfI1bB4NaYLGw97LNrbAEeF1rQCcp1Fdmx
+2zedkO01PgKiZWq1IiyNRV2pyTSCb7CH2w9YkLLa/MfHHYzCrKwEw/h/dscbqAEqCaZYZu2i46Y
Z4MK0UGH12CsNTGdACGWbSN5WV4TiCDPxj95gXnSu5eiHF7IkE0y1ueMpqyy4RFWgBfynzYUwgoD
vOvoXlI3jyMUfJKcYoIQjFZLdOza37cbJuJcEPP6zzTzvBASwKv4HYBAHRBlYJZN9i1SYTHYVrb4
fpI3z5CXFNCxdR2qKj9w8QfPtGMdt7m8fh7zN24ppOKi6KD/qfOwaB35ITLGIdour5agUyRkaqfp
8211yE0RCul2giUjDIDARkebnSk9TTmHUrzHnWMawW8byOmy/XuEcDfZ88Zz3gB5UcJlaMDyyR+T
sysTsrEwJd7LNV03fZwZ6+5ucMSX50C0UCDg4cXv6GCR5brDYDGmIhcTSdh5/lPxUDOq+qWBDLtq
VnpENgUlecRkqgDW88ZqvVL6UbOjxWOXpQmDwozPiwMIUeOXsJz1akiMJvdG5kfXl2ESHc+nqV75
xsbCpWJ8ySE02PZ+q4rMcd+k1Ca56l1oo68dWz9nsbWxpjAUL/faWVeQ01kHZchQjdJROghuPwYA
TJt1FmuYdaSDO4wdAxQ/5s8GOuUZ8BO4teh7yT64Uk/fs3eYIQjDs8MYyoBYdBScXpgm/kAgv/nR
T117bq97opggXFiGKWb7RVntiHeh6ZzBDTqUXSHKLkd7bqCZ+hegobdTVhWv0ub7GfA5aVoWEh/o
dyCVUo6f8K3wgZHDfxirFH88r21tno4VCjLGxkJZecaKbIlzritCPc/vWDCi/lSIg9rIThp3Kl5Z
UrYZmgOrm15tUtleSMxStC1IMZOFfIg2ONhBkF2G9ww9c+8TqztQmZZ0i4glbv/czk45S82sp6IM
VB4wDW9kHCRHIzc/8ZNpnmJ2gKUR43N3jXK0dHc6GvioXLBQraB7WVvxTFmANpGdEC0dAgJ+3dAy
Kjeukio1dX/Ic6iBwxyHhvngV9onKay4/Ufn7YbfoAZTB+LSAXbZRm8h5Qq5EaTI0dd2WkXpl05x
qc99ix2j1qqXvJdmK2DtiascxkiWL5tryaFAcdzCjKihGD5w3P5YfgTCBFVFG2f4j4CVhQvbRBpp
P+I5DiIEp5HHQdCqwrZPD5RJQc4uXcOaGZFyxvmsSZIk1xPvB1qVDUyWEXANrkE0Z5fRkSLjSCTR
xTFiN0wlJJ1LIa/T7kkTBGL6quL5UY1eOmwPwOf5klWVdL9jJjX2JyTfC/kQS8eelnPtx8ERMAu4
rEMo+jpdNQsRQ8SjSdRxlHUdaB5xMloGS43nvTAd2Zi966BZXW5dcV0XlgZn/J3yg3eSxLM8dJ0J
AbX4J57kGXLHpCQcgW2f0nUuFG7PhTVZKWBQ7QKdIQf9/GGzuISJ4XTPQ9mS6N6lcOjymuizjeKV
4neOD+1yEvkuELDXHYoz8tE9lWvLspds21M80JyDcv1eN0spN0tmYew3b42dp5OMC8rNXg9uxpAw
vRlvDrAOROsk038Qvg87jasNn1bqjB3nQgYF3O29WCEYtZ9ZSLgbcsqQlu0smIferpbZy+CD4iYW
SLl1KDdeZWdaK43tCwOiQFyUFeqf2NQWVJTUIWK3ggmplxQyNZnDD1foPCNGTc0ricDzXJmYE0O3
KLNSVW3OT3rypJq79Y/xaOo8GH15U7gJQzLae4oulx4WoFcqIn7Vr44eJcUlLE9QzEO+M6jCjIGq
VKXrVqQy8JwZG35ulIJ/5wMspSIqDXT+K+W4S4eH49cQYvuDVfjwxIXr5DKS/e5IKvyZoQiJL4gu
kcIiCX4p+eX1L6aIZvp2m/Xd0roz8wJ/H/FX3dQRwWAgITs/fMACZoif/9lU/UYqPBYnkychblpd
8M4wLA3ngR/RZpG5sYUpuZOhZBmc8biIr+AX/f/tNDUe06oA4fPjm96d5lj6kJ2yQ04kxyAw4X36
eLwD6E0tgq7XGDP71mzjZnH4LYmG4F/cfC1qhsNM/psWVARU+nO3L40UoauS0YE1TaGGVjY/nSLH
V3xkCasMufIb/UyBV1gfUyq9ON8upPrkgnde2AZjICiUEpM4OoQczzBBlvFTPQ2RD148U6Wt6k8b
ydgxVx7ZkjjlgmrLOo28nmdgFbBbNziJGbdM7h8s6MR8o7ZoXOQ6nghx5oJFhKo5XoUbx0GqoGoi
klzSC/2mLxQIu2QojttoYsFob9y/g3sZ1jdpVl68LL/66uHNQXdRLAPx4Gtw/HQtvNPHGgyzgN32
lvVNDDxwaGsr7LkoMpeIJ79ArFK87QHL7ARYE3jakNnvhWxBr7vOeioJutVITHVn9qB5ApVeNGIC
WCoNyU9YoqI4mzHcD5cGgb8QMREh21M0rwyKT/bf7fcEUhwUXwglqSjUBxfpHsQpIS0Rs3FY8wjS
HjseY8JU77GwhH3NNI5C4fWiBL9M4qmeDXBic8sm470z+hHGx+BEFb0k/4PIae6ezJ3Np7wTE9Pl
kIh0dklyYT8y713UwOIBM4mw1JpzVHKGvXfdfdKaJS4RWbjrqr5r2flVg1xhhdHswObKq4pnwvT8
ybUJiXhrR4UR2uEXBBVsvEHIMjIikTdeS0ZrTd9ej0uHbabDAjJM6V7O3DmNYnWFMBmQ8E9j4b/q
wOMWXH+RzzE4jru5JMxEOp8pCBQpkTw2cT13dAl1WdmP5wut04Md9L/GJPaEtf0E8MhQZ45bDMI5
CCbp4AevpJ5HSgaF9VIrKhTvyhOzLtvCJW7WJZDNtWB1OcpHSCL9kLT8oAcBhZpWYkC024W2xUQG
YSzNAa4D5KOYB9xNNvLl8RceO+HORE07rjZe1DyZuCTra+Qo2LgdMIx9f57II0nnIxvqlU6Ew53r
9O6IIcS2/eIvUMgegyIZuE7IdPGOuPEaaYcAwlIPf3q9pz+22ZfKi3YysAedl/ap7P9aM27k/h46
KZiRu1kKRZUmhygB4/rjoyDv9BLtqLsvMHtnwOYtYl18x/WNprIn5ANXkCoAUNffjDBasQEY58va
ivIRa54I+1U9reh1pm5mvn/kM6BPJvv4UW9sAdgGdNZwWT7+yHln7zQ8OJhQrjHtJu401t+DDeVI
pBcacxzVugPshJgEfiU6HV3LQfRTLvEIGVcFsF87mbHAw+3BESykjjqIMIivKKlad+gug2l8W8CC
ePz8W7vI0Gly7TWb6Xl0XsqH6qau9CtE9jj63GBblgOiIiGczDqLivnnrume+aYy8doPcfDfCOzR
ionqD1GpGfOGKZO1LmmF42Yqt8KB1gDq8aHQ2ohlZO1FslIpIWC+JHij7GCSsZsh92ctNQPPxOCR
IWU6u4Le4oqb7PF+Zj7OTSFwxhw6YPLy2Zd5dEguqikM6pRDxdFPaOisY1TvftkJdyF/FWIO8sXM
Z4tQNHwl97o0zgTwxhTUWttfqNcp3sImm3CbiOy8OihBslrSINOQvjPkT2HwwnFQNmRQsB3ru3nS
XJ5N/Wr60w2s5ODtlWAV8KT0Yywg0AiD6T9AcVVLJTdpugV110SjsglhWhItSIe8syiKtYpCv+jH
pdNZ3Z1ecjDdeULfd2VPFMcaSPUs1nzECfBJSgiqj6/FtD/lI5CEK5A2yt3TWZScuYZOtce8qGi0
dZG2mZD23EMaE7F/q8ijDaI6Nhf2Tds3faHDySTpH3SeWH9zUwHhTnVA3g1nhAsmVnzEeqI02GOM
I8o4/nzMc8dcqOwp1ZV2ypT332NAXCJy3HfnJ8LgNY+Dvb5x1e9h6khvtwDSGzblFPQIceJm6oLM
AoZyBCbTVvFdX6F9OqwPqTh9Un31e34I/58RLvsmTOFIRxje3kD1FSmZk8C5eeoz0YnkwTlI8wDo
MFul7lkoValq0ZlEGsshcrpUX//UZRIT6oocvIZHQMfDfvEGbQuln746WBKWemyvmtR1nFCe8gBo
eree8YtmcYAf3KM1A3vRF3dr87oY9vFkIgzyqR2pAlA9+Hs+9FpiUaLCOmYQ7ZCWfnSrE8/tVnuj
niw0cbjUPO7VU4pEsOzDFIQpWZH5ECZdGZTtZ+OgJ1YRaH8nxdkrGcOXiw6uFRd26d5OEaM+2d4b
EREcUDKPRBD0+8rohPLv676Agfgnq2/4bch3tfV6MAP7WshTfSHk6bagnyYTTP1whMoWLxJ8h4bb
igDCxRLtmDEwYmbnAWsaxuZKskXKHbEJpzv3uJKGlE0yNMjQToyuHd1YhUHz3JXN18lMhvxZ2iQP
tr9/pT+XrsbNvk52QcQb9B42idLIbO5Xqy+BRr6obJ+7pETWClp5lIRPrXTq8Dg04R5VkZ4PvUQ2
86bs89Sn74RJq6L9bcnE7orMo67228j9HkTU/OO/NGH03aQrVqwzk2uPDSsEkpGLexszyEDVhYWV
YsI86wLD6QSvlK8C9pXB8HPky2zLuszePqkUPMZPEK5QTDKP64hkQExBIE9BS9qTL3ZpREFHJcNl
Ywo5MO1jqdrAyytk+7lwGaaz+O0CnSWU4kVG+umBRYwxDdghyyVZkrsnPiOUojW0IM+sv6vkTadD
vK0FgCNn3by8BOrJ1xCkyej4UuNLhsa59Ra5JmhQ09Q8S6Jfy+sQWVBng3vNoUxKk0+saXgojjVv
Ra7cHVZED48tETYlIf6i2tHefIUnszGp2jKxUdog/Lb6NPRWB90KXTeCLHa8g7Q6DbA61Slh5wIW
4rm+yV9F+mcd7kj+tmgwnWPhyOrr1rvY3M2x+ZvS0lZDBesb7gjDEZBRNdwFsZD6NTG85Bvy+suT
x9O6m4FXmAzOU6fPgVmWkbrQ3LXN4UGimM3iVC3VXObm3UDpr6c5gIKXrpPUFZBhJqisDzeuqT43
GdAw0B6E5bQrmAWtUHSfdEHnhUBYa6COeLLpNtBrGJbp4Yej9YFT21T4cSSZjdoxzgagfyVWkrao
/MQOfPRkYta0zh1C4YlHlT8bNiLAqxUVFmN0UHBEnM9S7A9/5fiNKGsDvyFSWo968o+C2WsR6DN5
+tIpO8BnCLHZfn6x60mF+zfdbOW3GKpGEfNAIeWezAJhFo8dhmlDXH0N4BNdS8oF7N/0pY1aiWEN
H89VTyszLz1xfttanuNVpuAv/17N+/Dj7byvah3uVc/NJ7vSkurw7k/SB1+8SJAyHHb0wPT9dSQr
R5RdsQyZ4vtQT44aU2XMcWIAGRbK0PmNwhp+kUa0YtRKK3q0IX13BujQN6pjVAJWf22Zb1tolquS
ifQN+MxdOLxRP7gUvZ63jx4zqL+YXpanr82Rr5z0lMWCpJyZGMvbUdx6YBJidhupDejmqkxqOyCO
1B3kCjeDXaFtpcCby1eRPjZbCj5VQKbiP/tdVqcJjtaell2H5IBTJqj9p4lVKTntitEjrCLUMBTu
+1F1nATfV6vC+dK2j4FIiJCiDqfuomOunI3J6rpx7djgOS76KSRXRIPXi7QSDtqnOaeSxWQVoPg0
f0ljO+KgxxtMd0WgLF5/FrX11flxCCUVqQK7Y26vFPkBF5j1mc8sdHXjkXm1xZ9OI7rbJupPN5l/
+Y8wQSsi14vnoz2ydOnnzveNM5tZU0XBdAO9v+noDku7K0gH2QhlKgIJoa150ahhPAs+ywsBGsdY
apTpDIrjtjhQzudCwzhV9hm85OxFdOOTzJi6APScpwXBlL1FU3Etwgn5XALiu2o7AtyNTceekiWa
pRT4dY04lNydSaHdObQf6p9IaqdxzrblsQOkPQrOqR8SAIY+8AyB/glZHWGAc5eFwI6EZTnpnCm5
bffa9kdnyG1Y5jGYeQgsWicAUItCXs3lgcx10fV3h5oIwFRXKJdhrwREYKHCWd3EPHRxqASAQNdy
KWJO+edMreIHG1rHsQfhW67rASivh609kMzteWPDoJ/w/qL/YxNqNelURMuXkQz06p2zQLA+O4MI
NqXUFHCBsheW6/Dj1e4gnibIomibr6hoCfm/GeJaB9TsqgTf2pX43uwdMsNyzNF8bg0RoahkcbHN
BDurrXaLDUCKzXLQKrQLkXyvp2HoKtOi1hDnuMmEtPuQ3wlELy6kxGhwbVllGgMPqqgpozZJFfTB
sHujp3eimJ0zQxBMOSHNxdwMTW9c33S7e8Ch5qzrgeT6At9P/T94EyQtkyQaMcngNPkAd+1nc4pm
UGlAMWw4cspuLSX54wQsgSxydBOMRfmnmui0T7C6/pxOrPiqTZcBM0RZT4FFnzS4rY5fB2AJgpn0
geyrYusM6gOnjOD+TqNEHqYcPfzd/zNk6tM9spvmgKQoGep/blfC0eYkO+B3R7CzlwdOBPjjLjoC
AvC+NGTiCM25fd0j6+T11B2jXUpQ/Y0tvcWMT/2e+oPZocooDYAJtt5vtPcuoRN+b2unzfKHyEcz
YwsU81NTThWOyW5cP92ctrho9R/lZORzxd6k+KHNhTDi17+JkPzBwwHbust5VgiDHK3ipvJRzZmA
V6sGGRg/wccgoLoqr47s/YXWfX6+Ws/twENGNFCgSnV6QEWiP+jb75c5/cUhHMiu1qUg6e2CjDT7
++QN4ZjnfHP4z10nnAX0CRPMr/f8cH3wWCwMez4igC/L87+AvXYVOtamqmdteAjAYRnpxoGpgIyU
ziUzLBVGyZ8pQozsdUMvdhqdLMLt9tbtMrp+oJ5vFKOxULacR/f0bczcN/8rBuxOZ11mW1ReE5mD
/mSaApK+DDjDHqUFf1YdAs9ci8h3RaAwxLECX2DuH64k9ZB85k/tiFO4X+5/pq+F3MN8LNxZFDl1
4tKOR+WkBxBoMJSOEbLJo5U0vlC7ODgA6zbCNej3de6iljVTMs4SmqRduLW7eSslwe7HIlSAwZ2h
6vnUiiKfcwWFwBT1zUeZZBQq3qPiHbK0GTnTiQMCwIE1yY9RHaKPv4y6AW+/21YR1uaDpnCTXyRZ
RL3NY7oT2Ni8NaS4qvmWKJd387CHsk1D39DnqEmuYb8fy6Gse0PGWRxUrd0jMd3zVQ/eoZDY0KjS
75JIE6AFESRqM89CIoWUdIWWAne+/IwwbmP9HizH02ZVHzCrODAHRHIhNoRoL8WU4s74l5rnSBDQ
JdgLqMIAERl4fT5EP67eUgV6T4rzoguGQr81D85akoTgu6NtL9xu0MWpxJn/HBNcCEHdvow8Rl8c
i0BrfMDdPhXab1uzlN7opcnIgKe+7WOiLy+JMN1Nbqt1XvQcgB+kSEauSHivAl3JUaCkxP9CmBMJ
w9N6be2rmgrDeeBmg3C/Jud9QBF47n1jqetpNGiNvfUegOcJllr+FVf48GWKG8PhS6DLKNITcErD
fEpHvr35271y8OIeMXGbsUyioDn9FCbFkX8yr2k98nE+Eu1lPJc4Iq/E1h9nYaxxRW0FFOxor4d6
lvj0wMH8vi1D1paCVJvGzyV/XB0VgFANcqk2E76wX4nCkF+dPSR9VqZN8Wa5bVG5CgTpdw7NmCQL
omkvwWclE8f5xg3zEC28gvU3rM5gx6qoEuINw62A5kzfbr0gNIzGUAePZkgvyXFe5nzK4vkv225a
kJAY1OIKNoB0QDUlc7GmLWIGhttSIjVjrov4ozs35dmFEXWYJ1EzbM5sic8yvIBFyZO34/g7Hjns
Tetalgoi+NwUTpnrK0jlCrQhsfynJCAzhhSuRSiUfvRafDZAgCNhl22PRkBDWG3yisqFbKFVK/Bo
2LnIcjdd4xwQ3rjp5ekUuCNLbEPvcjtegpfCKfk6hM2rVKDHwLxcNH/vOwtcUvAvWFOEfj7i6tkX
Dde3phfHpjWtkAvmmVeF090LmzlP67mdix6ZsDi+s52ay5tGJA60ALyubvYf/6SdyZvhj/U0x4oS
xIoK6q1HzJVv9eo5C2lYHjQBMZYWg2yD1Ofa0GO6Gx8/jj2heVwdEAORX5Rhc/Zy9KaCaClzgwbO
DQ8ckAPudfLZf6lIptUGwDr2CudKjkJ5CTdztDbkv+a0Y493VP5MwCClo/4yRTLzFnIuVt4cCkW9
48D0af9IJYDG6MIx6pyneQoGiKdIIS5UfRWsbFx9YKHZjPcYR9+x/qeFf+UIaS2KKiSnZ2MORbAe
89RGQjL/UdXGGQzgcjvdxp5hMjtofLwhc7EdICEgczRB9g9lt7GmcY14w0H7q/bIyTykPngb5/07
cV41zSLbS+S1Be4GphYcg7dPWVKztV8QYs5/PznH8azjlYAIVjJkuB8Br3FPZhpwcWjkeTkensty
LOMkUxtkKrd6h5VzCZKWs3hU5p9DfLe5ILWKPWlO/IwwUVplYutqOY5mhwZPIwM5CvHMQcxEE6Ua
mlEwt9yOQ4C5p7c0DnHkQKqmckXLhKluJhZ+f2t/r60iuSsVIzjHEsqdqBXnTmJmupyCXeD6R7pi
+bBOG9i3npEHaeE/Ma4ApF79K/WWMmN68DV57Wbhc63U4iFnQOVv+3DXN6TWXA4GHcvBYPFREZs0
ncgdVr8K1z+sH1JJwFgi+EdB1H2LO6gIfMFMzqETAymnP16USVaKSWeFgv83beEwebWb2iQevJzg
rWdGJhgaUgqLM8onMLcxYJ3Lk1JbFsSX1zJGBoR5BHSQ6V6C03vjm09Y0ktOBFdqfNkBDLFRJCWH
W/BCDBYPHGbQlsi+YrPhliOOtzs1w4LFtguDJ3qPnFLh3vdN75cse1hqoYO7H0TBzmctzOgtf2jy
7Bc5kS3Zh8JQPk/0ApZqA7GdqMAQ/pswXt+r7BoARU8srehJx0CugknxZO050u97SHkb4UmaVtRJ
hxEEwiZo1iHBO6y0xp8YZIUa+0DzcbhElGUZoDVG+gt828V/7H6DwkvXSvtcKZFVBq86nsmGaY90
NUMoEuhcgc5fOR6syzkASm/o718y8ecWNv5HQlFbODCl7qsg7+MoHJe8bWr8b05duSeLLoXucbLs
BDzOBsQR5u0nqDQwyuBcm98mWbkZiSEAalzEXj4iXMQBaRfNf/7OJj6W4sBnHAyQQpcPAQ6l/uRv
PkEyb6QYrt1AEjqD4WaUySMGQDnqCfyUB71/knIwm3WfgZgJkI0Ib/Y30CpJySLeG/Uw8jPzLPIu
TNCPuzwdchbdpgdNcWh7CGmUtolBOr5Fu4il3MgVwDR0RdAe2q0/CWlFswDvtIgRp7fi676tqR50
1IPnrpyJL9eKJ+MK68FAWrtEAZ1gIMD/c1xr9O7ptFEugNkcfs1Z8xTwGDSpdDILkxylHSYOfXMF
Xe+tksZqwrBj0kItaGnNpSEtfx4f5+2LCrFaQrMpl7/5c3nQsg3XwZ2eFK9ivC3vsQilnMXekKZq
oHHCOgsGLpmtTMHKDg75RTiMrjcaz9qikJWk4RxHHnSUgLTa5FaMCxjvNwyMZE3pzMfikpNcWlDI
oP4ump4PQhfYKv9JpPx3lezsbN3wq4nYNMPniP2dp1Hoxas1IZIkcRkqeBsa6x+iTRsaegWweSI3
rB+gkvxd8XRbWk2GCdaMeBhhQP4/VW8Hm2ZQMoqymmLzx2KahmLr0C3pEGZ96AmQuenAeau3NNSb
KWxevSx4pgHDcpX8YwSsfSMP4XJv3AeKndqbOZ0X+IgvSdGXdL9Jq0tq5tDVSIvJ1/SsQMD9goJe
pTxuIUxh/ZgGcQUx1soyTENtJq//RnXemWxf9PcFBSt3hdIunPVFdJGUr/cIm6k44qkE1WmKDm4S
N+0ZTC3Lq53d3FW7BOQK3q+ROmlFSHehWwdk84x/fr9d7Om/aI+hcmq9UTzNE4U+9ODPmlO89ms4
H2WDMFMOUJI1fjaqHrHg41RdkFujrGo64BiF2fyOMizTKaja53v+nh8yZVxOnXWMm+h6bvGLDBzP
LyB+YJGQhEn7veSrXS+i8opqwxac1B3QeiNosQMi5hW35DOgWtvW4sbkhCh5Ppop3s0e99GK7F38
VN9dDKy5/7UUqd64IKDR//QhaUPzyftgSkcp7vBILLWxj8FR+4mN6s/Jx2fZ5mQdF+ekjWGxFDCk
nJogWv0DbzP4WYu+JAINtFy3ibgcFvwPL7KhzWAmcKo2mPCLUwXbFS10M6nhRNXtqVfXhDPkv80/
gPAp9+SugK97jf6X1xQvbL6kSjB4murOWWykIf8WMKqcn5w/J0UhC9e9do0W54PW0xo+/yv6KIZI
HHZSqQkUur49r9QQnIwTTJAP3eVfn5sJCNZaqAgWjqROgaVgkKoGc/ohpQmRvNYWJv5DevHMNV/s
JgVmjHti4FoQa2ESgG5KQCPzekQxNWQ84Qr5cT9INx2HpJ474Bz+NxUCzxQBXVMqxBVsIbG7+03L
4dtjZTKxzVUF83A0nS0tg3F6X4091hXEAHZvWwCGBbN6zUJfN2suV85YWpC1jemqG/wztKZlMUol
fE1bKQxT3YPIg6bW4fB6gDadMHQCiudJvf4gIxor78IjQ0a9IbwbuovQU6M/NmNxx+A9tyNUe35+
MelfAGPDflEEwAdaFIZQspNA0C2t+9DhXgtm5+VdHWwrJmGCTRb0yki56wZ61cJx2jyFgqssmCej
SmTPqSkG37oVOHJAUNWKNGXKPAdIat1YaQb00kbRLomiO+Orwh2pCyBkQlMTBN3+2OZcLHULvG6z
XeS6PMwtlT7CNYf2t2aX8Um8t6QrTjtos92NK8LymfffAsOzzOA0pAg4fvQb364JjF0VMdWjAgxs
QGGFkry7u3OvG/U7KNH3ozgL6u1emLnfUc9lSFk58th5yQHJ0rSOxAcr6Zy9sOY+wxq8GSLXYdDo
ci3twV0HORps+5D4syB4Lk34CJ4E0wvF37+dn9SZ/DSjyBDyPc86+vnDNk1O4ub3OWE0kBgJX/D3
rmXxi/mCXc6QqfPGHhhAe+7nktBVxUwqtyn+zoZ6e2ZFzsiErHz8w10ZRbxJKVZFqHsKMXViCGv7
ok70XfA/WML6Z83Ps18X8+WMhKz/FuoYedwGlZ9lan/5eodX/k1YP+bLYzws5zCTjhWYdWs7+cKy
hn1AgzjEefZV4hTwLSxewingoHA8o72JjFbdXcBRgRLsLbc3Sx8EFWGbeUHR19NqTTdnm18CHi9r
zU1HJqCoQxoSCkJcE8f+iBFofD++5J4xjgy2ZPsBdHKtfh1nE3/BWLdSNdPds8Vqbbyrs1CoZ6M+
kl4wJkDVmgLy3uptVx1ld7v/FQlMh4/3IzuiL2TmcRhV54pVM0qYBmvgF6g5aZfz/yz4Euf24FAo
jLXSGej/DZW1UOr+x68HZmlXAFgnt669ZiadT3ndrL66Pbz/REuMvXtj6yFi3FIy11+55R2Va9/V
HpxCx6yUi+A89mTAOO3qcxib2QDTKT7sOGjEvciEx5i+ZxvnBzInJpNosVkecpiARPbMpPz3/9s4
Kz6uXWpps76vEpNM4HRz2CWf0b2dAoBafP7P/UKVTjdSu3ioC0RORtBLEidNNHboGdAasyotmIyh
K+mCCp5yXF3EIGRE0Jb8AKCHWxbP+/BHYJWpxMtNLX32esnhBlOlUrALEB48/3LBMb7q++uheAlh
4JCyWG4u8w0Nb32yOAGwa7eJJbJZ8uILaCU8rNXMZFUPprwfj78U17XJelEK0NP5BfG63r4r7vnu
g6z8yICJzLh31YaKNsSRknFZCitNFq/TQ0T3r54zaZl2Tf2CqmNB+Dl853oopkLnr7iVHG7HqQp4
XGRD/oPaJlWgMEzQfM0TchR/Nxu/QhUnOdrULColADoeurhxwsB5aAZ3PvsZ+vvJPY9155Fv2iqs
fj4kaTKNFJj7Z5EkmRUXiz/41eT+NrfmjCqEoZ00qdCj1m1+g80GwZvlBgndTJgUtr4hQXenbhoB
0peb1hMbiVg8UGvlDGsHekXPopQvzlU7XDAtsSbBcBdZUCsEqWCae90syqY7JDdRU8WX97bbG40i
EGhlNUqnkpppf12NiHpkJBWB3t3SwKvtLdiDHbHo2C4fe/c9rcDT/UDa27MieiOn1PDyQHScy7sT
pAHV8vD4fOwycPnE7b5MA7mWPOFftR2YPffrJ5TPfk0ECLX2Rp2k4IL30Nj3ZcQk6yDUCRqZBFAN
wGHvyvJWGflbtxZpMgsDbbIWu2fhVS6hdjnQRrbEZiZ10GVgQ50XhP5d8Y7RqYpo8QIJLN2SsQeU
bBBEGfbNVZcpBVbcCXiV5yWK1nmMgk6qlShDBoKAG1i+GbtKaqHAd33l2isk9ETgvMMF9LRYG01Y
RRiwtH1XVbMnkuHPnUaC8Zj6fBZwi+oYxm+xjsgxur+MXcGML8qDDa3OczfbzJEisQx1tDzUTBHe
UdBOdgZp8XdWG+vLDDOZUFJTmBSn6ztq3CruXqfhucBpMJ7QlyEBTeCmVke0sfgAs6YOFbM7Zbhr
FwXSO0C8dcZaf19sE0H8f16Cp4WFGiac8fC65/HwGnI7nGHYUgg52kgfWSIvAerJxRH24QEY7yhR
p79HkxbzJ+czkLFnu0xpv0zPrRpYFcBFT07ZKaKTIOxqtSF8aaBHbPysrqYeRbsvnVWAK7uj09/B
rVL6BinVnauuSMQIPiHd7x4ZYzs1Woag1zusTwoD/BzCGm1vt0uDUvz/0u62R3RnooxbNhc8fwly
yG6geKSRaC0JTwgr++Nhf0ZUF4ZeoRIOJBWK4+nSKxpFfWkFNx9MmohE+uUqZQsPwzgU2TClkH2D
7E9MTXbukvmRtNBfTsL4XARiEet39RLoQ8lv/2t/lrP36WPTu7/b7xfMt7w/Obe4l6bLVr0ZuBjU
ywKfYRQIBv76LzqPkXmUya1mvaf/ERm/uLEKZqluxutnSDZG20miRjTuw53fszuRyMzoIfKKq5EH
4kCzYg+UAShRO0bnqN7JYq+zYzGTXvIMeziIsYDsm0nDaRCHRSZUwqBu6eeHC7oaLv8u0sWJO0AZ
UPWXI75cL8A5gor1o6Taa3GPgyg4Q4cRaueNzT8bpm4dd+qXs9o+s+hb6Ov+tLJG/o6nxwO7UtvJ
PEZaRvv3zj5MU7H6U6iI5spLabwGrpaHI1zSQtpSonbH061nFwCA+HRzXOcI8fB32zN1O7M/V18a
u9BF0L1qvhtGwAmLIMYmte8FYsfGf9Fkr6qLZ4UxNU9gf6S4um+VvXcAa+DxYIOzQOHNmoJU+VJQ
Bj1LwaFvLl72+BzRN05EUL5E8OrmKSPqXJ5IPrO3SeQTIuxD9zSb2H3ScNt8iKWnKyhYDJzgh35n
E9EoDBMW5cErFImY2K0tScd7IhzThyyWh3QShnA+SHBGX8hnznDhpTIv4ue5BfibqeWToOQBMulf
2sAy0wHyaxclJkUMXbxrgt8whPym49b7rpX7VsGrD9rEjpYXBuUB7ElvtWsPfhlFrQETmYVz2eiJ
CX/X/DS2yd9XrY+LrvwjTzjWolREKzFtsJ+SgSRUFsq2y6Gzc5qXeaFKH1/IC/TCMt+SyTzwhGb8
Rr97F26GlBDNkAoOJUuu1zNfVSvU5AdgIFd3q55rmuNTx1Ehxvhulec0bHR/HKZwubeWoO/NLWoi
uUbWC/T5aubmMfMiGvaj0zT5rIrlG2yi8Rxs5zEl3KH7fELH+LrrJbvW40r4JTHWA2D+YjlyHZbr
o1y3BXrdkvZsJlr5aRJtbDz140vYjZ46qDvgAdX6i4e9HsbLXvtWK/PRMXlfi2BZzLyUxFMtwPQy
7In+4rzizhCxr9/ug9qD0PkFKrLxpHpHXW8Klasr91LJIdWupstQWrj2sErsahfsCXfqZc6Tv/kb
PlpXsxADPor5o3Go1v0mzkQHc3npXM0qyeCTPGCsAto7ms15KM/b6dfOTMnY+5/L1zYZiDuonKNL
/KhuJZz/uuP3EW8z4j1QLAZXduK72S0Y/CxqenKlnjudvLLoiUOQagWnGvheeclUX3uM/rk2I1Xe
7oX+nGDA4w+dwE4oO7wRJON4Mk1k5lfA8acVEIwdPXmm8ryyHfldzSueecOMtRco2ALV71/RJ2n4
b+5DxribweEKFNdTYVf1uAzLuRPCbFHfuSRM3/5X3IfQXCpZmqlXM5QQxLxWY0h5IrCTQIsBXnDE
WQXsKA/lzCPAdHKAyx5IUMZ79U41cWf/U4DEorgAn0Vw2IJmqQx0pcpj9t/qnsLYgk6klB184bFX
V5rP4XlYibgyH1dtZFvDfrxREKroOXK7eB1fr5juAaDI6/b4LLDioslq89PHD7y1O2EeYJgHZrmL
Sw4lguexbMbbRoJcRKtxoU3WGWcegtQSDWBf6zEbjayHT/i1iFhI5MzksWzC04LZtqY6hVL+1Hy/
fPfE47n49DWSfQdOmNif91Ye1HwRrE56wp6XH0t7gQZV/LHl90I1KfN5ZBavv/bJF3a1Wr/bTcm6
8i50IWJQm0/0o48yZHuYXELRJLxDe6gc7PNBkGcx9JBQXgcbydjz3BVveJHDoMrEdI7JyOInyPhT
fepAIMW+czD+gUvx211T9KkWXVOzhwExUMsvtnYm6gq5S/p/vGk1iqIDTTT1oBtbWJy+ugp5jyPC
4/TRNWaO4k02fyiw21IY3WUSgdqfvHkNQAnJn9W4xyOXC+0FhsHbNXjA/3Q2+HnhMyNq+A8chO37
z2yMEeovokQG7PQq8ZfgLB8LPFpO0nIcA9QZZNh3Xs0FwORxQOGwUxaUZU7H/U7pB4Q7op1lDql3
r5GvnH0YLhSOGR+yq5OL/s+dPwRd76akPapsPiXrnJ27KxtjJL6GdM/e8vWaQbZ64vCBbEEzL0e2
NCKWTzN6evKk40gCAkGH/FSRWor9cydP0RUum5fpU9pkl07179kdynoAmWGRYZG33PrY/qKD0cEO
AMUkpAZKep1NYpek4uu/M8KmlqhK0kOptmJ2E5hOOFo85zEtL5+xAOqRaeQG5FiKH28tb7kwWdbB
/oE1hpau9uT08fJxHEJKQlfqgDkqU0rQtHb077Wf9gbLwpmCiUXY4LqXPInqa3OWUw51zk8u08B3
U7yKZHQ3fhkuDuf3m7wzKM5ag+WfoTVSKLAJZBpO+jZ13pM7jQq1Vdb0Z7oPKUsXl7s/Tx9albHd
k41XisPvaPZM3h0hwIfAciVtJSWuwTN62EQdits+435PLD2Lk2ZNdpmM1ixcHfd6XcInnd/07Nxg
oMGIzkKm0JxBVdM8bG4ZbUp/Jb614G9FI/EHMiAT2kEw2vY8fRr4VAd3z93xKPdPzdhZ1gFA/LdK
HYk7JzF/OOgn1UvEWdW/vz48WIfEui+g6XyxO8OiLJsUiRbHC/PVamm8IKyDqWsP9Oo3JW7Z/dyS
ceFPVPbl6lmSHwDEGX0UecCjHomaRh9uiDhncX+ATV77/JzrSBNlpeL8UGCSLrkKoarnj9/G7iRv
AZGTrM5CRxeLsaLzu55KmMeS0v8UkZ+EwBUw//FV0jmwKoU8XkxIvgWOzphxi3sudGXJx1zFX6Bq
E4hVurrBHC9zm4IFncoUI4DLHOJFWT6y0CYZ0Q5cVCJboWendVTF6ThjKFwev2FyiDlmfadge0Jn
gUoXUSN8wiY+fLySjSiocNrVFxRtlqu7jECMZRmxYZC/9BrsV4jRToyaD7ZQ+L4hoyZlZeylS1l9
oFhBSIdj0GYVhRiSf5klo4ma4GdmB7On2/HHYFd8ronq5wF77kksaTbU/PiQsxUjSaEKlXFu1/LX
HpX7yrAberEzAQYVMVM3t+iABC4Rtwd5LIEAODtwj83irKwOy/H94Hk4jEqV07I8KgkvdNTLPuKc
oNUOUy0NVzBaEpL/2tuz0sPs/Wuw6sBND6hhxYR7bZCQrpBz1PbAIePtINKJLfQxn4vJ7XGpjiQL
ej9V0qxxZwKYkehXkUAwJkaYRVPPBotCF48au6ZG6didluPCJ7aDPxU8MS5kKHniKEe/W4Hwp0Z0
eL1k10qgNZ2LypW3e4PuvSqqmHK+C4svOa04T8tgplO/Hdq2JiZGBIEcYcBVJhykr/Zso8TOoLLr
DRSe0UtGhw/SgcA6t543X4I7uaCK4SixpEqQ+FD3t+/Yexspm3mSHC+VOU01GZOuMXdyvCotJY3M
2MDGsgaB3SsInmTW/VwK/xRyN4l88tmGjoMwnkMqoD8Ij+k8tfQqX9gvzWymoyY/x7sowFSRVu1J
/k0g2jb4PEvVMUjdj1jB+xFyiFk8ifasdX9yyAxL5+ARslyLCWqglF6tp/Hpu5bd/JWvKqKFSdKs
OVTceq7kYdoz0pnQ9Zzuoy0HfFrDkl532+LpbQ32kbgPtKQWUDjWNzTin3qsBodiWebfY/vpjCQF
GdYUEdqqmv6mYRCzFy2cZkWh3a/WWqmYrTM94G7eQFSlMy8PVmJc09OC9JU5Tv7iYWvBfDu4fo5h
iYVSF+GeMPynWTFIs59bmL6LQvQV0+nqWZ57mNl5Y5TjPEgmN1IVvSYj/8oJOsGhwoHHGJ2gI8es
8p4Co3g3zZu0nL9PbWzUcEpV8zE/kKvVHBxp/oF83i0EgX6O9r3C69ToXEMrksL2GOP6FhdHFqdI
svNdSXzBdfPBPbfe4VhIOBxVPdNJUXXrJ2Ojzp2zgGijra9l2JgCkfJH5QDTutUqOtDGF6e4n1NP
571rrdRwLZyfCWIquyOKKa6xv16NWF8buFtrmf3/aY93//n38M0P/xD/8W91AypwK8D6IypN6g6D
5rFiUmsSDL7DbiaGSItds/z9vXTyekhytxOOsbpmU8RKY3EBmk0K/riLGcD5Zk4Yh2hHeKnEhWpB
dgH/68jYp2qmgfqTS1FM8Eqc+1xsaGAdxzddMijaE/k4oDYh7VhQ5ioq6EZQwAyPCqqjhb8NwG6w
0FaJvG5TUIU+AG2JOVJfTLEU+sdV8nQkXOfBxbJLJEQh2qlV4a2qDBf1YJKeauKcYiNtQmOtYCYO
ioPv81wxo4J1nfrKCdnWHDHIYPDZ6AGA1Xatg1/9WA4MvktRiYJgU/5THqvXECG9Pb5MB/Ks/bkp
1jM6urcq07sx9otaf3YkBND0buwS6KvQE0oPC49N9O2pbGc82DVSCunnJ38RxsNnbLeTgoY8C5St
DixSPTbKVKdoVAx+EyrPDGZsnewXy0Ze+sdFyC9eJ6PQPxM/R9DccMNbvtiwXKSGTHGdX/lrZ6wm
eb2sgRtZ8dzomsTbMBIk0DjyPE7nZk/3KjyXvw0o1NLWMZE6F+Rk5ieM3WWTQX2xP4pWJP0DE/9K
DBF2B0zWixB7tYiol3O3ZRiCTJuUTIAgosx7eeGNevIs8XJt/5Eb/WrvXvJD1HD8GJDxIpwqeWsD
qLmLTzSW+t4FX9o3ZB1EhuXJbXjnEmApvprlzqIfW5UMbysZlpjLHZ+1Rkdxe3Jsr2Xaw2eb8XKz
4skPMhBVi9fzgb5ul4boYMV6DNuQ8Wipfxmq/1YoR+JUt0AX7iaCd3EQjxUMqHezdgbXTG1f8nu/
Kq/UFPJdMEnpnDWYNu0eHDqfs3+7uMgB2o9D2BGRJz/Y3eMwLvUQd20NtI2XjDADes0tKdAYiPhi
da/9aqObe3gfrF1VpZZC2ssG+7ogkxwbcp9Iey7Blhhxy4DgG5PPjJ01KSQCEMa40JOG5xK82ZCK
KjFasoV3TQsrLD3liwBhBm4cPrUtJg5ntGWh84e7K/qAyXyp1FDufR0mJGdbqN2BX0tBwSlhgoaN
ZelUw9Ko/qNvGhMpJvjmohFE3LHatjBcfM1LGalTN2BxfL6hwb9RwNBHhMEZCUAiVfvpuyjiL4gM
vaQGUSuEwjIQLZZxS/zrrV8jngGHx+Rcbofc1Qgt05RiLF8uALjwBR8HkONI76jRuVLE/YHMEYON
+Pj2QC8qhC3yWngM5mSe4Ytegrp+EPU7bfDf1blt3zWb3E+n01t89DV8/JdhvJhecT0Y2IkVySs3
FyOee90MmC7elyU2mRoVofEMVuezevZfLGL/t/nvmNXIEknw/73EglJEuXTbgv1Aie9Yd6QmSqld
Y0lKsebirkRfrWl2SMn/6k5HS2TfO1nuzCrqZzqpnxbkvEznIFnekEjYKqupnPl08omtqR5CyywM
cApyLc1OYx4SoFRZtMq35ym5u30rQyT3a6Nz9O5PRxtEISbJmbS7ZKJ66U3Vc3td3ZZT+pSY8SWP
BHo2pS52T+rttF6LH9cgvJKeM0JWQifc2vvRRVBA/RZKW6EnnpTha92f0tXg2fszcWljeoYgqjxK
dGb1GLWtE/dzoAYKKYUX2WzTU7YjctMHoNxRZZq4F9+gWSitFEY0NZWAeuqQ0LUszcUvTufJ6aH2
InJUgPho4MlaV2tC3mB9VEakuMxHCudmH1QfgQw/dMvQMxMvnZUK3YdCMbdtenOoUopSQ4q9PUhs
eJw++ASIZYnWDKIzIzkX7qm1NjDEYOuz1IkIurQ3zWO2w5hjzk6hbTK0yLCGH40Kp40gsQT3pAw8
RkTGafD9H+qkF1k3auweTEKWyPzEeWmvrXmPPmLTTv1neNd9NEkntYQuGxVu0gJPEL3fU4gXMmvN
2vz/yXi66mv2H0GopE7fZ6MIJURTLB3pLfjK0XG2d8g5LR5wb9Rvuewf1KrpEvYF/7AfwvMCHGsP
wtU+pEqz3CSyhg6NjvAar9wsJt9wAt/JO+TFbNS67EuJlNURXzE3Lz4p8SCLOJ/8Kj96/yjM384m
PjY+2EqiivCoiNZtZT1LebU6x43kiQ7pMRYRDaKPViJh5Xc337vyArznFpQyMLTv/FUwrhnemuYd
Zjao1nhNCptwywRDWRqv2DgPVP/OEBVeZ9UxPHQwcOLgZf2XTV2cXJIDWItuyLJp9f6iWtbyQXlW
LqPFEc/OAYqRdxARwuqRR6/eo9WYsNMKaQTORNhuSsWEpCGDOGoPGvlDizGccTXgsTSP+EftsmQP
JCqfRkJY1HC4bla00XtrOt0S83TtI2uqi6fM5Z7tgx+9iAlw3hhFQnEWdJzWRYb9fq0irOpKmoNX
Fc9sXVpXQhCwYgNe7TQfiAJdQZWwQ0eqJMW/EdLXTIbhDGA8cXGswxCD8+fkpZUYgOvgL1ODMul+
K6cQ8FsJX7CneaZG2HRhAv4RodiYK+hj6mPq9rpYEuAaLFhpChoRGU0bQ/ifCOKgUCRu1f6lIs5S
/Uey72jh04rLk05u5MhjxafD2XiqQuKqDB3zHw6m81NCcPWHr6OmzCxyBMOOe+jKHqj7ChRBCyUV
GmdDoOkjHuh4guThapGdwuQZGaBfGXkTb6mTfYaoJ4CXVq3k5axz3UX+EqQW2E1axiuNWxtSltOR
ltzRGXW4UjBn5Z6XwxGI4pzGV4r1maZGhRkwAduEd0Smzao8LSJSUkcA5/0/dKmzCL06mQ6qKvkJ
w5hylMGbpiaaq434Q3dYn3xbQ/JIYVf8UVEcEgYrikc+FvTos12RnSXa4/pIqFxatXdDE3t4ubDh
wpO0AkBzJvxLCUWpCoRjKEvF6o9NcOIMVSCD3MARXLYIxWMAZtVS2PbgKKWG4fZV7ReacvMvP4Nn
YCYtCnFTJwaS6awo1K0c3Frau+9N5lDwCNlxE8YiDXiJBABwRtflZw0XUzQyFNhgXHR6m8etMzi8
5NfxZG7uzz89kFNnsrVV4X00a+40m9XtEAL1Nm0fsCSZrfO5n4Jbmz0+u0EUAOO/CJH2dQs9g/Hn
Be87E9yLXYbrZ0uIS+n10k7IMXGudxA29jznRS4o9mjJNuFHDG3R3nvUNnjpHJBicd1bz1yafDcK
EKB8WX75NFr2nb+cpwo1sPmUWXpm5kAsm4PaN3USfy27pT+9kSmS3nLkileODnkz5IAKSgvDYeio
3fX1dFxXh0htw9SDoxL85IkzQ1jYedl/gpF5jg+MUP5HjzW1nNDAAE4LLh72m0VmOiPrUOvaG7Wh
WHqixyvddf3LqlwPINcY/8hEx0RxKoqVsay6ampom3aFYkEZwebOKAZamgsH0TUR5yjIC9ychxjC
AGUdgk4Z4sIAizhKgLCFRq/wMYNtvrOP3LPhuvCOqrCr6buIWJ3hLcO87GO+dxVVUlmkmP/5jrY2
Brevgaz1mf/fkVt1gDelmn8vz3qU7M6GfPqYv7iZPatNnO4PlQ5Dsu183rbuu1O6ikXhSQ0Anc6J
kIxe+i4nC6k5U15K+wIj3DVhOFrDr9LlwkIMkpOBZZad14QNmhYxkAgDTyg2ghlinTRGcqiKQWZW
f3PDm6fItQn/S4DF3B8M3FDcWoMRz3+7N+aYlrlhi/Jssu5PW1SRLpmDyFyXfZFM56BSgCebBWsJ
U40QHZZj3pNbt+G80bFZmzaWCTYGnR6+t7oQOidX/AyQznh+g1w554+/gsv+y9IUblh3MtuKzxoP
Qw28Z+QfdLdQgZkqvZYgMOilS/ia3rmRgs39klqzYBs4TcCFQTzjOXZ9sYlR4uPzYUFBjzk4kmne
jMzhWy3JODbOvfgdQc4uW3D+CQa9emryaRIliTYLMgoNtWWDFgQh+A8hyZYEn8BWGRNxv0CfWzan
Zdztk6U454ayt913q2b1g3+otmgZ5/xGyFppSenkgHpg/x377JptyBsJi8Pa5iKkmR85RgE5Zzgy
227n5NRNVwYH3DlNG8AdBzFJRTN2hysbPPb2/exqEByBNdZhBxstxjfphkBGcZPp+hbIWbFtf6Jf
WMowuWS7wHbzFZPqpec7iSucZdXgQmgOczwVJDPejUbTwVlBwfDs12K7ywd1EfnPocd7tdw+aGTb
siZG3FQ1RgGc85cUYLK9jMn6qdlGwUZsN5Aj/2BFv1U+U5cJje+0zsP4U/2gtUMzCmecT1CViTyn
2EPiM5qgrf5/LOvDfP6hhdBgSNS6zf7PP4i+DGNQuQlgmuAGss6OmjIl8DNXOztJHafh5Ew3fKYC
y15KHW2ugxlC0HCOUbsmyrB8TDxmt8C7TEC0qeSArvzOXfTZgGRd39zgZussK/5xNqtKn6iwBZnm
PWw6HCqaSKyXAiHtgNxOH4ijCngUOm/JZ/Y/Q8Qy7MiX3wcJp7eISWg8YuONpW9Mk+x+QpFquceV
IoIIufW73EUAp2af2m8Q12zIEwwCVlmzIXN/viEw2yGlepFzmKwiH2NVLkL7B38/MYHHYlmc2fh0
rvfbSRMlK+Iz6huskGG86NqrDmjAUz31K4sDvyb+zfIgTeG4SxllACs6urCCctPRNgwIX0QtgplR
ikZDSSHEO8Rd+6G2Ktyz5qbosBOm4Lhnr/es2z2bY+wJtBwU8wHE6pvwq6SCa/cX4pA9iyyniHJJ
ZNvBTnX/l6x92XCF8/zaIIm8yyEtOhLoxUG0K8+9gdBc3U49KJAr9rX18MS+rdd1uT2JWX85+5Kp
/9i68HhvXIAKUHvBvtILZ+f/Dt7YNrnwsNu03R2arwdLjtuZCjkZfanIWQaACF4HLpYEW4vNSBUR
f3vc0T07hqZlFNug9qXoribvI0YXwXRbFMKMfAxPMaidz1vSdIxKSttrmNzx9W2GoTJtGhnPI7y9
K+W0O8jBwFTy12w075DfvCqwQCHPV0dBp1rHlw6+f4xzc+r/lYQagADne1dIPGOSdz9fB3bQdAHv
5Ouopa9zJorTb8VOmIWoQrbwuMjAkEO4sq+a3Auvt4SAfzIgp+nkQGSPGKdIWbXXJ8jrsFehGfh7
OtQt/F2yUUBh7gl66ZBMnc+WI4/04nqvsY4l969LckLlX2eeYyPP2qOeMf5SvbS+uFaPhANdiEjp
Q9t1F2OM1+p5H4kwbFtGx+xVW3XbAye07TxqUje7g0LiMhjfR0jVlo7cELZFzm8+6hbs/+4EZAiz
PQadwb108F86rX/6SaolAdCHDtgprCryKjCHXY8012RJRLSiitJUelWklxtDotvzz6mUHKuasWBD
go2oCrL7hKBjCV6YT1jOxCqOQc/SVljs07bPoMcP0ST8cFR4we9f2QpnDpUyfNBRutYh6RZX2tHW
nDV35y3bUaogKK3wSjQchwgg3uH/USFQPI/d8a8HRMfCRR8mMTX5VzwQ7iyQwNXf2ZxM2Rlx9SrR
Y5IbNxTrS7ir16arQ4IktZaNhh+OmFvIPkXis0HstZh8pKe5vo8NYxEKmTAthDXlxHfTd3JBgq7z
g7Zf6H3VRS7kPKcIgifZCrF+g7HUeytEdOV+TEy3iXWiNX0JGv5kG7PPLoZdnS6YDYYBrdP3BdcW
WcSztb0Bki5PEJX8A4uKsDIlwklm1U9rpMBNmDpJ64N8OS56fDz0MixSgQWsWStpVheR3K1+e+bH
GG6uLyEVQuLyteXcX0Ez/SkYGypfIfMa4Os9Ozqa5OW8Lkf+mebRMcTJJwyfwy6xQ9BEFK02G2jM
orqSPOyxwOT7TYpbiYvXVxKpkp/up273WBPFjVMwgN5Bd3BJBEAyUpVYumOzgoTOrScOfS+/S7ln
iKmNgVZqbbBZY7M1pKzGGdX0NIjBtKFj/BLEkFz4PdE46YjOuPBu9Vg3beZRltF1Xb9ZvvIougbS
AuH2vVCJ0OfLPNgBAypZs6CVsIR2EzHgElhDkozBQnj7fBWfmGMKuZriDvnj76XIKyDoy9aC3ZWg
sxG7y7zmqJgiSVS0/0g1Vac9FKizqxwxS/YDEko1J93jh+vxL71agV1XduhZDnjSZ3kmF4ffuD+y
0Vn9auut4ayKBbK1AjJNJaxfZ1TxWVLW8T0vJtolAyPcTszoTC5TKxVM8PAUW7goOlSDxm1b9EOY
EIYt7fVmeQiz4SS0QwqxCvBE2AS3T3pqOylISM8txkAxibeLfxYD06sGxEwz8TV/FfJmSRXcAfxP
pvYfZVGcFebyQXUieZeJbCJt92hW29nT+HFWo7RBpSSJW9XqFNYfxx+k2TBtcDkDFKHrr5k+aWkF
RMyaNyCgaYt+R7pVzkn0THz/VVaZyIKA0JS+DoK+H2FXddz7eO6dMyVaILk7ARCNk3U7oAMRfIkE
/P8cI6tjwBmKSdEhdGa9eWXDFDhPyBeKESoX7habmO5QwFo03iFuWRVx53i2nAKIS0hRac7cusB1
cXtEVGjZ4mPq09+KmRCHgrOCwk2F88ke1kEn02t31JSHXuDisWOu5iVK+L4OWiBXcsv6SacKIeSV
kwjDY/sHSIfJxcd1/oDs730yMcrXn9ZS6qx6AiIcHLzogh1t2iV6pbNO5B5Kf1uuTKhFDO5g0uM/
hlWbE6cUlfLwWaQGtsGaDr8NLt8WAvrs9zueqzdAQrNSlYirzYBsIDearSo6FGleY8OLKvrJynvQ
9/Zi+GhJG9YC59YwtNhhX1wFX/hOBzyGgSgCUC2wmgykRpo9e0T3huCTy6XjAsdaUgsKnieveajD
Ca9fvxzTYqJxXTDoF0UjCrssLFOOLpa6ufb2tCqX9y2gfATHRuYb3KSpAXnGUHJNOWDlb+vzSjHO
pUzxOZUwJQKWtnVRgWlHLH0vCf5cAWwOrjiah+fbeRWgE4thBsKFAvu7jfJfeIiDk7oqcIpvAn3Z
8UQhRcRAkcGosBbTKGjcK1OqlacS/05i1XcA0cLNLu7Tunjs1oEh2gh6kx2yDx3b6zdL0CNfxDWQ
V5xQbbnkig+2z3TfxL8NwJWkUf2T8rq1LPbBJOuRJB89I1RLxsP5KKX2G6/BinFGQUv/unB3dIJL
YNpIffxw3KM6nvPvL+YzzAWH/fF1nbV+3bqwZGX68CikWZn/MI4JLxX/QExAk4q0gvDlx+uYNOw5
BUfu4Vaft+7HwXuwjJoeDJ/OTAWzzu4GmhfrOqStWsHfPucxWW16Daxpw9hvCFvTejj/UA0xXVKy
KQtdUjXuTSAiNaTHduyYspMF6cjM+Lx4wX1HQUGM7itKZNJL/LPlQJFVCRCU/YAw6+hAErhBU/il
J8yj9hObKWfbVWyJ24tKdEdL+qm/3F74VIIACuUPIy+EQQ/2c0sbsfAcX0xa4iSl6lChJfmhk8hz
2v5rbflnXWvjAAA+wMarBbF/nVA2FxOWJabBK4ugfQnWsIHCwDUDFDEu9MAq9Fpb07OzwKAs/R6C
aLR71bCHaxVrqt1PIagX4UBbrMMmd779KeudpCMYkTlU8M5Yylz/5ymjMi4ZtDKWK81RzKN0WZwz
g+IAmDg0TQzYelR8C7bQsPoJbHdeoP64ULXqnTHIU0SZ2gkPadY0ea+eL0J8N/bH2CRzeOJDDHSL
Ov+C7wh7aXCiCTqeoEC3ICDuJnrrdf5XWZQmgfqdkNDH8DHPCCgj54ovfx4BhFtyXUByzNhthTfL
O3L3EgH6ADMIP7lvzPXKfi1jzTt0t9/RejXqiN/nPLy8439VgX/KCf8pZPYH+Zz894HbG4irGHpP
TXSkRRWPXvmpH0FPvZsn+FiNULZvr1qOLtrUR9Zek1zdeB4vzVfzs1kk7RWWY6F26eo9jEt3Ah/8
s3o/0SIBOaagMhA5VrXMvdOflICvRBVru8alfU8NUmkCSdzLdljJYng93iBhI/r9dTp+Jg2ZdRpN
dGo43ZlzOCqFD3I72uNOiXg7PQeS+gtLMpRzf4iWx29+RAi6+njcFcKilHXRmnQ20kclOoP3atfs
nR4T7mwAQWinShJ0KTAESiEkGWaRN7IPi4C5LX9Fv93/itfHxR8khjRr954HWeDjmOU/aWflf0kt
M5Uy04NxwJQPzEni0+UPx5aG/X6/3YuJAnt5GElp5Woba4TT0TnrJDLXtFkSI5IUakOlza3pMmfH
CEulsjeM7kFi9zeE5lTpAyvecPIRK1LWehZ2yUXnByuj46hlDEjdkm5kchF3nOOMrHb+RI5uZYdE
G+aEqiMWqmz9FxQl3oHxv/1Q4ncwmGVfjZkN1aIUXXt6FIaDYfJkf7c15fI+mcaZI2lJ/28+wCHN
t/qYQLHYVbFrxg588F3kX2FYbtBhz2MfYKZB9g0DaR/lbo5iiFpLH9Bx7w4HoZNWqnvt90UL+Epu
fiTjt/jWzyPJGi4Af1w48hqROhwoG0fwFJKcCFWP/y0iek3BiIu2SAaFaqNRJ7qf2m3HMTVoW2yI
F0k0JWwdlhzpEGhO42cxVcfjNIWQxeYfybYYz5ZxcM5ZvF1WlWSA2f00Z5NloCFf64o+uuEPBPsi
81m5qfTI2UqWRZgUA6eunSSJdInzPZXLuovkKEdv7BWI3dzAYw3pwPG1kyi/802i8K2eBVZcgaze
phSAtovd0R1odI80HxQG2W/l8R3MqKjGLqNzer9rl84w3Dr1lqn/hVexRxwDE81BGUCn4wJg0ium
1lh0PEY2kot0TZxbA2sEKoWzNGnZL16ASt5nWBNIk6hcCZwxE4g80o+qLMxZ5sNv7vKosEianZzc
5Vk4j0xYayepiYo3pCQFmkhQfoOF4IGCjK+POuZO2uhlI3KRDnxmDRc7C1GXujxKqxrp0w1ihglT
ZHLQNcVZZOarv4Yc6AiLiAWUia5CwyO4Ak5VsoQW5DkWgxnzAZAa7h8Y511aMsojNG7r35jjOFul
vtpEwTpzpLpmSYVfZVeTsBhCC5z/BDnLjXeHGDSAArdRbU3HVszUBFuQkYyomvOxsDREfzhH2aNF
P7pnXEd/MtaXhDlD3LHtVcA9883EOBfkKqoJy4cBFSxAQwA39xvVAWO87MGVLxBhhx2JN2yxz0zz
hGR/hURjpvRkjAOyoWsN5fwRxW/syKpTxmcO2ezRrdRCyikM9l9L7r8t4FXUNEmpXz+uFLrRuMyf
GESouCb1gGiktdtaM1zXWnHWW18dK+qcJn51DPPmAsY/2i592eM6HRQKJ7tAN0SLcJbudXGObV73
GyZ9VQH1puaHxcpVd6zqtdbI7MnoghfW0GdlE0Nak4sD/pJbRDEMyNSuMK5JYGXQElCM4WdmCOYx
iZB/54bLXMClQPnuVGjPUhZEv3gXUnPnu7l8qOg6Xa/fUr385+QrE8KLY6LImYbbrm+2z+/VE3qx
8kr7CDmcrxRhj+2UEBBXzmOeWCdP/Hn4LD6mhzkNdtzLXYumbUQfXaqYKC410E1gf2wNP/UstOlK
+fnyXs0cJTfwi5owCZnM/xncynnLJi/Xny98smMAYKsjwZ77UG93TD6PNX5eq7xoseWUm+viDP7E
QDLnn4NdciScsuWbQQNzwjT16an4ak1u4GL/WKYyZazniGL6K0eogFnv3iAcH7v+/WMHxlzxvzeM
d6WJUImU1488yktBgTpe47Wuz6qJNm4EpJbhkId7EG2t8he+qZE51E4S9XQGiot3sTtWTe3Rczt+
kgZJ0wFZ/Hh1myCtUyjRPyk2cbe3RUE/kFf83bbwoI69dWKO1OQOheSkcxtR2gOxh7HystcIN57V
vxh9TiTckEv7Em8umo8/xnO+n0l4/C3BH3UTsffj8ZbYx4CW1weDXt7z+e7nbvC48ftP+NexcYe/
wkZxju1Zy7ib3gpfUvbLOzj9DVz2Ay8H9ynVRSeG7JTT9e3FpQtm9Y6dtvSvwtCMwVI0zVwfTcPk
M1zPPQ+FMrIZ1GNGJwmp6paUV0ZadkaXhC5f6mqkQHuvZ/+6CJNxYspw4iEoKpJ+aBYM07gAjt30
Zey3a6VX2ph2fMZyfEH7Uc5ZFxPL0YnagFEwbMGiQUqu4ZQ6V0/eEVRDrE6JpcAtT5RxYvHI5paD
L4NIK9azKIt8AGVnjmNNQzE2UuHgLL3Ukl0xWJKCKXekCRw/qXq5+kU7nyklrwL8bOSxSPiXx58Z
wla17+whwpc4gbG/G8FgcV2I0gVIiF3J0FJPBHft2S8HY5ucTTZ863CbB4FzHspJQiAI+KmPWHeW
GLE4m95zzlNexhXlld78OMoWZWQwmc7fltZZpZEEwU4Ma+66j8R7fSdJwsvJp2d1un2N3KPqVGAT
UA5ie8gZzhq+nUiT/jDUb/FQelSGfoHmlYzvWVAhpDCfXrL3X2EiyZOJx9RGhF425QneRSzSgkU9
emueOhNStO6ga9pquMgBbudWI7Ly5o8Kf+z1FUnqT1hi1Lb33gkpgmy+55wqcsVxpaW3EFefvhqR
//WHwe3G054sy95XhI2bSr871C0bK9A5p2tUvzlLGLs4+C6Gw7mIsMr8vDWy4qUmnEX0hwLKflyJ
414epAuuytUiYq7URF1hAxtnPPH4lzV/xyDSD7SmExoAMp9FOLcm8pCQ8l8/+LOq1y3rgipDT4oQ
3KTBAW97XhLQeMYAXBMb5Z3P1V8iA7N9T/3NbeSJXwVYN+bp5arANVXY+ehQhuGcLUey9OO0UF7z
zyJjOioBCTjwWRtQnSpfm3+OEU2NU8al0ZQmo+qzosx56r68Jk5PTCq3J0O0E7KEAxoIib0CxNKF
/URgXZQFCPtEykN0WPCQX7v/ULH/V4+k6Y962cCIyboxjwmcXXA+a1PupSQTiHAKOHsmWSx0PKjK
6XeEr9eecJAPAna1/6kAMwEnXhHwZ3BqD8PynzeBXZxCD021+l0JDWOwyKFt4t3tYkiiVI+1YOep
HEFRuPNr+Qrh90hdOnIb75LpBJvBSZdG7wkeESwuPFcJHgy/YyHiPbiRb+vHm6XimS6NcuQ/DF1J
MRwjEWtaa4dmMKi/T4CJurw0fbqKP/K5ACCFYDlSWCKmvl+i/39UEIrYRaw6EybHt/XuWFHFGiVz
q2reXuYwwWnqY+69ZVFdTg7/wtySvWhC83Ik55zegvJBRFLloo8PE2lWoPJVklGclneehUAJedJ/
3BrH96J+PMZGa7dlgTa4LbOVbTKVYAFFt3OO/69EjhWEGg7Qq12u/VNgZNq9LjQqzUoL3U15tW3l
1MYhCqN2bIVAkEQr66th0REazqBzCeFh0YV53PJqgb0S5z1PomD96aREHNJa1EyVI6Vze8PqAmAC
dkHJFExhgSML4ClJgxStkmjYL79ZjCcpu/NVyi0nQVERO/xkRaIJL3WUivI/cZ5BJzDVDzSduuk0
shXxJ/Qxuqmrkw8ANqCa7CnVASbyxIGBJ0j02h4AIdW9mY/6F/MW1T2pQ9tyer7ThFeev1Hk4O2y
wW7ae2/iUdCLzNZ6NZXDjHnbwVUsZbc4vbj4dfCMCoy03BKzCHJB3A+nEo3dXClQ2UQSf02I6oBT
W0FWbWumved/OGLRanwdU0FnnymLJXo1RmKNRqjYUOnU8mbfpsf1jD2S8Z5MI7roTgmWhn/AwFAY
Ec4EMwcJlkIRa7St/mL7Utt7HajR4ivtrmzOEYx90l15MQti7GN97iU/peTJ7ahGDA6kWpVvhdn4
Xa07/+R+GOgFRukC7id+fPfwDWDINJ6hW5LIHBBn3r7cr4aFV3D3M0zNtmKM1IfXUXLBTjR1TEKF
r3CGFxzu1HXQ8vcTTKayEx+uc/2V+u7HHFBGQa64oOvIC4cmQiHrz9av2flmMfy759WmAcaJM0JC
BYEWRLUK80yE8tZf28IXlh3V6UvAXeU4w8mZWjW7XedkDC6tcl+ZIay43hYNv3G8wCaeXmdrvJo6
k9TDk85HC99W5rCLycrD/j9/tgtTVW8VaUpA/8xuRAjhSxYVvwrL42u0hSdFF6O2M1f7N5vrvki7
puQ+XrSdzBw5xdwfSj4GI2T35ru3qL7/3DNeWxPlEzVmAs5V0sj0lMUlrMKnSbfd5ECcF8x0vP1/
NWRBSx/x5C4eHT/Jxe61oSwMhYF0SxUlCwWfXz2wzZpuZyvbO0nqNM3g8pZa8QWUpyiK9XCTcNjt
sP94snvU9/DPpSdCdW0qccPWCeycv2jZvSMQ5DTSuSUpjkG1UVLxvb744qGl4P9GwlzqHoEbpzfn
kpejZ8UFUBaI/Zih5UVYIJ/Hu9cB+z1Ya+wHlo/yJTF4pb8JuN+HYSVSW0hlDnvTz/bSs82eFuKe
reJZcFNulv3jaHukyDD8cZSCxQa9xROc4GZ1KtmRvNPsMdJmqNZIYjyFSvnWGJXyOXWKJ/jPIjRE
0CQJb2k7kAhnmhF5jFaRZx8Nbbjt4kQJQazpCaE+i5ln0TdLTn2ABb37E+UuEMSZJsLUBbyNdKvB
21QGBfpd6nu17JZM+mZEgGd0CrV46saeK0IPx4YvSfuHsO2ylcOfUNZntD7uStkVNbgwO5U6UAcQ
QIAGSZlWvuJqaQAucpkWCRiYL6ZAfASiDfkp8guMIB4KgC/aLQlCjE4pokMZulpDN1heKu6PobIk
X4x+KMPajUwRgXq5LAQRNHMmKtbCKcF3F04yyNT6VHtBIqLzrVCM6K9CKowy0CejLK1ehhFaSGU9
v/wB5xiSchDKLlSZn/whQfVg+Tt87LwtifWf9ESDy834dWdka3ybpbY9Hg0y92ycAPTOrIvnD367
cQ3hjnSTjW2NV9v++8AgVWMo6bm1YO0baDCn22VPID4qWpzXmtSGVBdl6VMO+l1fe5WGnhzxROI3
xpMrd2QUbRoT1Tf7IGb0iRx8/PNxkojICRYwej6PGiQfm8t4ADxmLUFrgeQgcGdhixzdnrJvnjDP
h6VaJ7nOhIM4r4SpC7jskVT+dVCkEgdqFUvRudMT8srsAsH47KrD5MMLQA4wQwO5TRnh+egK4Tal
TAe3vzNAaTQTJvrXRcsABEZina50U2udCkMPxeNEh8/LiPXr+zNtDqJTTovlHcElxs2EpmfSFqR1
lle3T2eOCVGx4pg5q2F0YKXNN/aRP85YJyy9zBoTxl29Kk6yKE9jARPzvqpWDdHwTuOxCo9569ID
z7/c7y/9HWgXS2GDNQYlKskqEUnBa6geBWEc1H5KuBGC+is4ndhcMxzBOVOcVmk2QaHCRpLTG/mC
FH8HPAw0rAAYdUc+cz4H6NOqVZ24kEtxm77HAZTovCthScAnpcnzZsfxoh94O0FmyTbHyH+uwCWG
RsEt0cUL4Rc6cCh9MUSe+tsQmKLDttJL/VCUY4AlQ4bxTxywaQ8xIuC/d0DSuGSmL8sTP5jl5OCq
6MxnI0k76tnTtR+bQ7EJA2DDbjYk4fPcq7wKydeg87+E5k+p77YMTmRL/uJr0/jsiuD5ckJcTrGv
hxT96m1Xm7r/SJRtwYC3CRl2YnZbTNG4HlwsoocY2M91k9z1OuEAoy7az6ffEg/LLBiiTiCNUw+R
HuZCGNHSSBl99KHkTXoCjXijSaGu0PoBzNgifKLBRHA4+vCbE0Tm50ef9whfVzl1/lxEZ74+Sud/
RCO73ND1kllQoH6YSplQt32o9tuKY834tHSxHYtb7DwB9aU+uXlzm93QKIXIWZJ9qNbq61zGcT32
wqAZLKeQ/Ut3Gxg82dDt+oaNhFTdune+8+MjCaRUe4iGGGs2BA3vP/aCmyDLkV5OBsT2NKk6Riy1
+7sZMUlD6nTc+vZNOmjzgmw/LHSllnoKv0pFakgokvowlgbAwKmX4GHiW2KDUfM0U/MJwDDHvuJw
5k1xDWKHBalyROIjlToQTFc85ryoYGWHbF78N+9mchAtN//31vsn9yT5c84rAXTi7hGDBVOq7kSA
SovB8tsJAklN7Khd+ouxoWfgbBts9wuq8tm9z6t2zCgnwZuqixMuI2yufG9gQjLm8oY4W8Q0sCh7
fiOeBfSunEdfO3aLJrCQgBVPtXIefOYN2F+R5CsIt+PS9U6akAJMmgPXLxHWPYpWuzPKxIM3C2zE
g2JWbJtGaJy7TL5ttks9B4PUN6cy9wqD7wKyKlQYcMasvDlwOaggXE371Vq8wdkYCXqAR39wyarh
vPUio31gWb8JVVm13XbMAxR3/5A6XA5c8Yy3jg4Z5EfxYkytC2tmTx9DCQHAgvzGjhLerHj6aqBS
nV++f1TUvPdwYCBGwzfu8fUExg1irIKDfmT2caXo2s0LHVfQRL4R0udQFQ1aDpZ5OQ5BavfgOWyP
HLQuCSnUKhHi6wWYOIQoY6MhS71dmmBYPnDJohGoKu8J2xtApFc/HpaA06+5KcB0LvbC5lSXNRXm
xdq1YCJZrzNUhOBMhkv8+5KSvdWQdKhs0DLA/AGdYdywOMBqhKY+7kKz6BTtSJjSsZFea63hDxBI
W6lqt0b9hQsHSgqboViA3ynpCfSPSUWpbyLR0mOYaKzalq88YxVtw1tXpP3F4GAh3ZSXE+Hbityt
3oOwNGEnv1S7EvhMraC0YZVmeAfeuZI1/cEMrtn7BgJkPjA/1Qy56SwHrGm0nF7vVMF27C0AglYU
UX1iOT1q0fXr7krBc73eTL1mbdOPU4A5lVSSbq7DyBEJHoNiYVnnaD1c6Mtw8NEgvE0PH+CraArF
fMkQNK72EWJE3jCF5RrV7CCJKJWj/lsUKUcM/faB0Au5KwUBZmtaXWjXh1R8WfmVdxLEX68cMkKP
sDp+0fTFpGJfquHwmJe87uLRyVMPH7kKo0rBBLAeUoQDwFvf+cBCYiJXXU3FEH2ofODp9IJHft5c
0m4jpAg+Vm/wKp0bLKfOkZketieC1a5NEKJ5ZtZaYAQA1eQTwrV5Nuxhiy9UNrPem4h39T0Xz29N
c/dEL70TXceTfI+Ibu65hu4WP7BqcXXJvqa17izpAOuNVvHam7cQ3ymAiCqORyRuXdZs8jSXc9LV
2hz5XEtVOltWMtYjQXIOMFhVvDX06/kEmiPE5zNkwQQpZpsN3QiNlYU7UywHDYTe0g/Rvv7Ciuh1
5P93NWPxgCZmRVXDqmxMx/OcQi9tO+gh+pfis3bfjhm4UCaZjk6PWrwK4f4itCdosuNcwLpIix05
DDefpwUfLid1+BAt60G/sAK+9egoNNvoUrztXdmJVIoiLap6KoF8qIAQXKakGMeUAe/KExlD9rLR
44clWEJix+xbLApkOSGI+QjpvH2VzthLYPN/5brhizFqnnUZEFxtIzW3uTqLxv4YDRcSd9+cuXD+
j6xYl23IQcixLbeJ5wFxWAttR7l7BqK66Af6ewOTnMHT/SbRAYppgsLszYcNR1liOXttY81xBuAH
XGmRxXn1eiRGt2LwSx0qj6Qb1669gxYSSNrnRgOT5J2d8WiD83mggEmMoSD0QWg1B46Jq1vby5Pd
D02BIkmNcDLtb+Bb6dD+CmvffEXXXljZbpbNo17CjpwibUwSGIqPY9k981pMT7vKB3OaAvsW3Kll
ouK8Zr7GmoJGCPEFCK3YEQ046OKIuF/unrfjwQ8dkC26dLxV0gxzu3zDfVG6FRqLeLhF5qcmOWhi
Zk3WRa1mMPxKcyY2BA5MUHIbiKuZfGVkVAkPAKy+Q3QE6eBAkT9SC4wIwkcHSfp5BWkWFh3J8CXI
/Ytf/xE0/DiQSXfGuFfSx5fEnCRYew4mgOqR17Qw3gvXjMvbwWsknOjRPimVb/7aE9VCUngPMubW
d3J827jXUX0KJULGgj9a59j9lpKiHJjMzt4oe+abAQV14XCarki8P3jyeGutnNd2qHNrXs9vz4hg
t9GPELA7wzzxv3xIxeBIsKZ/Ct06pyPcQcNDm0zpjl+ckloZOyxl6Q252fHuyQafSrJB0XLM4AsX
Wrhx0F/G8+yxTBzJEZ5aYPhBq/YhX90X48lYci5gEUBeTcVGQLWs3cclEAJM41s3Gdwq5YrjeilV
RRmyehDyTFeM93I+lTbfLNa4u8vGLaSB9/iK3JmVaqglqnNHchb+gJDxWoXLYfkmQ+n5VWgBDh3t
ih13hT1kPBq92JDlXiycEnP4z6EOnQkEMczicxrhAJp52vLqTXnWsDurqOV4Oijr82kIMvnp2TJl
w2JeXlgtJ0tnD6q5xWOgQYmwu0GhGCwNwsv9kOGWhXDJ8O2dcRRtPNxpsbDBmhwTgyFoXqdY4Zi9
RSly2bc/3vhhi4QCTGktQRmx5BV7ABhk1dHvqctvIueUkKy8AfPLfZVnjcIiQUkPfY1la0FPuwuC
GADDKDJkn0Elf4OQ6veBLHGXlmpEyx4ZFD7REhjgLsqBu3wXGDHmtKfYe7mO6QvEolXOWNuQ9dE8
gSxKP1XvZblTEyQ1gDfeQbkDNpSuecxTo6aiS0uHi6gsq8lqMT3Ou+jUonyxQZmosUET3kFEiBcZ
0ooGGuF6pQ6S8sjaExVg9ygTcUqo2SBPcTWDWFHyphKzM4sIpw0oHQg1pPfwqymwSVWtif0ambwx
99yV455JdOPwMISueRf8M9dItLplSrO3mPSehtF/kyJdH98YEIy5ok1uQVrNbH90m7pOBoueRhp2
wBWia16vuLVURs3ZbGdKeyOMl2SiElHt98UvPA+G+NVU9TeSCLlJbQ0G9+p89JaRcho6+0Wy48Gz
elHrXKl0NRMbbVK9KT1TRzN3nw63uijYQ9h3cDUNmLejztzRMcNBCaqF2E66d8QYrpDatl+LCrxd
bbRemaW3eopitIKvaSiVbUbnkLZRmf0lF9muIbMlL2nX+RzxvLJ0Smbdg86Mp7/dxWYynEBpCjvo
/k20urnXxbgsT7oLMztKttmFrD3n8ukaaB2xcwnJBZ4jFTZ5tGEZHcxYtqgQaEjScu2O5kr8qtSd
nHPfNHiP6ZuuLf4pVCxIaTMH4h60CrWJzwoFx82bVm3hh63NDf9+orIR42iRmgsCmusrMtZ7dgR6
GUWSKAXPEZzywL99APAeYhTfrQU/Bx1DLYJ8zawUlr3QQht2paGlk134vL0wuhiMwpwrdjweL4jF
uet2Bo4BNGoaC0FSJUK0XStbrxB0Azt3zTnRnZ+JAAHzvFy5LM9QKsJ5bYREKO6XTcGvrFQs30us
vpNF0uLBIdoCVzqRJqQaLx0N8sLBXx+0nVdjt9O2Hu11VV+w9O7vvZ8OQ2wB5gHHEAnJs70W5XIP
Wo30QW6wVHK1a1w6WURVA/dl8PzmE6c7KURa92sltjUS2cvpWjBhGKFCd8cYBZlcia/aD4ngI0Wn
qrfB3rAiH/LC2mVd8uLuFnPETfTgkRUtJaWFvJQjTSlQsdx0uy70pBwFgJp9A12/VLQcheeYKwhB
B8YBd++Qlm1q2TPeotWrLbsFm6tg2sI+iDEHQwhlwt9O6kjH9VEDQhgPrUvvi+jCeIhUeC7fZksE
c9zhHOd4Yhv1Ux8IMxSNQWlu97ODR+4DmBEY55m6Y8f5AskzmGcdgl39GSmxPTAdUlmow7656p3a
ODp7BrxzXs5iIithPBCrwdaPprHrJIFv7NJj9mEScTJPCWQG6M1m0DobPZRMbe3VKr2OsgRDc2Es
XbMbeBoIdhsjo+tVx0dTgW6MO0T1/TZ7Ka6WB36nCajaWZJZeXAt70/4F7h7AmviH/9ZYPHsxNjm
z23+gkoPxznVUhUovr1fHUVEwN/j0sBSnadHanNU0RuWw1PaWnmJ4dcR6AkylZ2mMo+UOshNd4+7
nx2ap2QPLDgwpTgHr9QqbgfLRR4CfQnbbZBu6f0MirnRTu7WzgPG6/UToD/cvJyc7+cIDlipivyQ
yem7bCQFW6b4qv6AOaPm/azpOexYA3hD4klCqFl9n/YgHsoN8P7Oi9STTGAPKlxACMAJ9bupQeX9
TljhmsPHNcgVgzzHCaxAcNmM/8oTwLW/kwZTiPGolPfJYBoOI4NkM6l/v4bhZw0GvIM+oOwX6uBf
N8Jm0PrrWLE4YQAk4v2GtJGTetztMNC19L+GtDb5ij/mJc+VG7hiYNw2IS98lkxM+Jzm0zeQ35xr
mZhrq41yi1X7UKfj2KvYKo5UQAzOfMdox8f91x0qlePLik/yKB5NxYrydQ4MPn6J+1LRtEobozJU
5W7h+arb1fAQbMoJ0HOxzn+5aj7jKzYkki/OmksNEmZtyDlBuzHc0C9WDojrDWPccwMyXfWEQwfl
kpgb2wZ16NO9SR4hMpm5ToYFHCZKRJEK3sQBUk+aQ3VhOily/jNDbHcBDvV/PswsOeG5KN2XdLUW
+Ew8u7z4v9dO3KvNv7x2JOSzn3I7BeL0xKIe57dBGiq2sXuH7ktSs4LW9+4toIuY0wrWM00R7LgG
YtWM8ZWHOl2hHcit88HwbTRNJvas1t9katfNVHiyQdeK2BjEn2yLVHD9SRW0dIDLc+Lkj6D/ABLP
xoRmWsVpdCtaHRkAJIVOFrisORwnMCODyy+IkVJzetNztj9rEeBReDqmcrUCR8yJl1dEUqD4G8bZ
GdpWhbaYCyqyNwPKPVxm+M6CrphJuaHJL9LaHm9tVO7DHtTtkpo9re7ySS6PMRI64cSHtdmUn5c3
sklG5dVpw22m5BXCMUVGAmfof6N+MNdkmankSmwvOOlmpm+BDYuk5ihbniCGEazLzR/FMF2ce/to
T0rQQ0C0wDysA2xMeWdhAhq7GJmgw8vTOZyyKfmP7211hQjHQnBAHDgO+dJzhhEt0X1w1xhVTskB
g/N324bmWTbqAOsjHZe6db578KHXTpwNwt9fnAjOntY6g6K3koDPnixWLy6i6/43HMVmGqSNbPFF
6C0tvVnW/dIEQqkkaiKfFDMh8jDqo8AWE9kKC6FdOgKhOKnxBadr6/Pc/8EDWcTPrm5eitl8eKxD
faTBXKgFHnPy4Q7PKeRF7N6bFM2ajNsQC218d0a/IxbCpz5M8OxqIoLRbZRlNpGP152UR0BBa+98
z0iqVnCzn0cqBcUXbM7cKWivDarR2RCulJxtZr7bEGyw5ayO6Psv7bitdkZ6+M1Brw5+PBRT2LLr
nR/z/uAocEuIuTKw2T6ibNTUaNPmm6PWZkDfWS87T/HYm3Mh+bKkovgow+rd6n29lNOxbntgNZoX
a8bni3+v7PwvfYD9Z0VqBSE+dRBZBwL6Zx9VEudZ/SZVX5va9D6e1XPs9VPb4luc2L0Nh0PpmhgM
ghrOVTiVJN+wN4lGKVMRSiriWzG0elZ4obUfjZR8Bf+7HMGI8cQ4yC+KkXGrF3UXKIMsfF7gTLan
2lcJY8ts/PQm/VC9KYyJtXxNUeZ1KaWccViqRFBYEjN/ElVBx//DBiduk8GJnUULcHiZRSTKauwK
PTpiwU94bmjfXKJsDsVa+5ojdYrqeNKzNb0wropM3NKYwyk2BkR6bD/r/uFxON3lKlfhQVqMzxRk
w/uWPrr0AdLILAcIOQUg/HBrsfz8xiJs6EaL05dlYErVuy3ds0euKnQd7t/7sD2ONLp6l++gosos
zG5dlhK/8quQnFVoNrlVu+q4m9nA2OVwsnRoy82CLV8yKsjyL04Ijw8boS26vsKgReljsb5f5oNv
OzxF+zebJ9JzkWHyPg2xgZqQkmOagc2tdNyGy5Lo5x9Y6hBSz5FNrBOduHn86npSVoHzukdCwBIP
i3Akoeg4bW+qRHTOq80JDlJl2MBAW/Csi8GfNQ9xRd4gwBaGlCImbLTiOh+mYGDKataCSOtBJX5/
yezwg5xvUUgoUS0pMKjZMBlnqjEN8KwP+1E4a2KUblUWZp/koldR/IEnv78AXBx+o6eBtqXD6bL/
kduyf/QX48vk2tC/Q57z2l05YkrDvJbxiwQD8QDXXfSUuOFm5gAoe4hIc9PUupSf8QE2W4J8vFiq
2kQQvFqrnQYl6F3jfk7eeGDfot9jcJ874QJWPbi+54TuPI5KLYoblxp595sB7y4Z94NGUtJS12Fs
yihqWhexhlCFkivgUpW+h25EMSTeOF91Y1jMt8l98oTOsQFwX9eZ9fCQhg5QMc6zfPvk9kit5wVJ
crr34LI11AP2SdKiHzQVBX4G9hkeAA2jqTWOggsPeAACM9hj5HwRA3Y0rdaLzsnbkIHNsPPuEOOg
xj04mcLpQWM8/HjU93Ph6kLVIwIXAYzCaXh2bEj1qJj63CC429aHNzuJAFSwdACRCpqPIG8f4tUw
cm/v8uS/SxRO/TB7QLIaoq57rv3mwTfbWHCUziyzWR7yg+VBRaeqzJxSbcS94m5GzX/m1HVNGFP4
/tAj7EOY3bhBXiJI9n6gKPVQoMT4b2V3xAcelkx9admpWDGqwEdQV5VdZqy1XF+CqHCarllZKJbO
7T4w3nnemyK20fLWEOmrRiUkS2PnepWgiLV+XkHEGBuFkqlwdRYzm9Yz1qhVH1AzFAJJ+kR6cVWG
Wwibo7ybv/gZ3lpKY65abbwtIDU+7d6465AQ0jYdvMGjvHaYBmw9LG60NF1E2+/KWwxb0lL6aXV9
mygca6l9YnYYxV1inQb3/a9V2ZLYtpqCauIZPPTu+WSsXNBrjlu8S2PNqPIb6b+cDQPJZdP2GzZH
h6MuStwjDwmhU8hqCMOzTGhB7Pnxh27HPAOrnEKEr04nsZ6bql+EAP8CSSAIszYEIFP8/CZTNuFO
v6upiJY5g/FtPzv/A6tgk10ZZEeXCuI81l3RZJ70q9DucEXKIn1DfGfQlhgVInxZCMx/0n7nf9Mt
wbQ+XHUIVRMiL61CLySNdmsi4kYY10sKR31Qib/urXbgTUPkvWWv/9o2vtPLfCxV0bXlHGSWKrkR
GoWuE6bQjYK6X2vquUtOwD3HlRMctPzu11ePa1iF3PNiheG10RNqxV/oMDy4eItINYYCJQahMUv/
QWzqYM52NocE9qQCFH4j8kFlwDC/2rE9RWapHgqHTIrAFAJi2SQRy2qK69cazfYCiNVvevxotzV4
aVhtwpQPNKTY4/bh/OJGCo3E9TgPVE5+AvFdql8WsQOOyv0QA2uPBSl5sW+rvVpy1Bq03kShO0em
MxZaO7xdDyAGymbeOgCDwEvjyNGTiXh7ld2eOsOP/+4/yN3D2EA94Kui7jRsQjTwIP8lp+8y/JSJ
Ttsi+OJfcPmqdGCDsIgBOWy2SqSlWoiwtdKdF7pt9t2/tXmsQCbafT/mOPADGrl0mk2XDr6xl7eF
1gKG1oOeTLHnD4uLYIoplrfz4xFw7nWFK2dUdxHcsHXM4ohQPMn0LM1xW7c4Zmk5ODM/iuFAsIE2
oGx8UYGVk/mYgL6SxSmcKOf7/LNv7xtokMftLAyBOS8f5TwLurnl0EIftaPlqEyz3MdRDmjNP7+S
NSDD7kSBEFxlmHDpfx8BO57tbao6P8yo9Hxvi08x6nnAB7613txz2mGOA9mGYvj3Nh2aFRD5J2tj
c1pJjnsVVN+7rTI+pRErPBSSyl3dTmguMqBfBnXbAzvlPcIhwwZE2qBgxBU+07j7CZwhYh9bq4dC
8VF3AJkHSxY9grMMuRYfgQ1GTLvdy65qcs5Y8i/mk0PKwMWuaZvnz2W+bsFhANobw15wwqYed8xF
r9J/T2zoDGz37L0dJALLwHBvd+d7TSXkxX7ecA4WqEzIFiAlZTcSXB1xG8Y6iUB7fr1IUyJx+XfG
faLFZxB9rSJNBs+2V1kN96uKVEfG/vtbL21e/AYnHyww4uvwMvTB5tu3qov18qOBEd8b+WC95ZpT
87c98mkgXsa9GUjZWpv9Xp29C972pjnRTptBnR3X7aXm3JDJn0j8mhEyttq3+BgkPIgJVYGnUdun
mGecYvMhgfOSNcfKuSnMtkbvVJWntuUzdnlRFJdrzSNgvOdCH40CoM54m04lThEHHggZiNOx78oq
pOJH0dF4s8qMG8TdEIvTPcIfAql60V3GUa58QQxYV0NGmxdIpOxbslCpNoUlOHnxB12OTMe53gQ=
`pragma protect end_protected
