/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzJUk8dcFq4JCoxWnokPnSd2U1Jluni2r14o2YwE5S6O5boAJnTFHCzAB
yrQDYD6Fxy9yYLBzBImTfh/t4DTvBbPxVs0TBLDM3Vr6lsFl7av5eWjMPuHiG2n05bmOsfr38I0G
U6E1KfNiu5r8Cq9lOdzvwpOcG2I5d64kvRhpQ/iyg0xDdRTuK2DPfkDbpfmgCnLRCYUSaLQ4Ttoc
8Lt7Wbr+s+OC/zt8gqFA4TaF/4nyEyq+L9K/xs6ZJzHJpKAg739ol83sOY4d2YXYaJ2RlHWVC37F
izdPWaJew8Kd7MlpCcKNpoKfi7HgjgJ0lrYQYRHBYL6jDNXyV4qiq+a80TX8wTqW3Ef9PcHrFi33
KndTr+EfvDbWrDQKRl1+Wu67x//LaqU7jzpTXC4hmmtSAE1eSfkLs57M6PTyVjdXx5evZUOvXdDd
aDjktQFtU2wnSsIZLhyxJ6IcHWI3ytZnfz48St9L7D5eTy+wahYH2y5ddiX8vMgwSvvcSyCyf6+U
ltt2dXObXHwjffUmyAX+YWWmbNDD0zsu23NeKxwYGpkqmCtJE8BM4nfQ/gLfc8AKBjMa6MyZop7r
YevBt9smCuVN65UshQBwivJKv8LZiuTN7br2dBakh/FgGBZDgRQYhRI7FHCxUXPg5HnlwDElWf40
pWF0y8ni1DEqQcJju4NXEXBsvKPqTmJjDTK7MUZtUnjfL5z5CZMY8Dl0Fyn/oiMoUzQaOwpUqByy
I3C84PT0+5m88e7GPz18QiwL0guBuxPZTZhK57YzutNsAblCt6piKogZdIrQ9E2yUinntIpcHzab
81LMhcxxnfO9OhtRzfw84YbMJRvg0LeBofDGbSvn8fZg6DdCrPmENWo3mAnDb99EDJ9ujHGTKzAe
EwOeZhA12wvU4ABM1XJrfkHnCEjsiE4J2GSAf1+8OqudJTAYV/hOEh39pk7V9tEfE+tnTGdO81PY
29/o88QrH4bmQiZbR9krH0n0ggi3iOHeWQQTWYyN2lj5lSl8Mj2chCh0xCpPuXlyRi9D0sF5cFJg
lboxc4xT33u1xsbiKKZ338Q5l02x5YBvN3vx5bgvXl9sLG9CKo4mPKm/wMhk0G0EbtxT6RalFtT+
+VY87ybHuz4nTMnuM6iU45/ME6T4/WMmi8N9tbm9iAwMKTCckK1aqvzKZF1gv0bRm2IHTsjjn8jz
irevxOYxO8UKdCQyGiZyt9O/gG8rlSRtBYaCigFmFEmwL2W9mBLIktXzMLXXqnOWOd3xd537t0WJ
IOpnYge1e3xRvfAi7KL9u8IKxhNe3yk7g1+Ubb4NSBAcNoK/zh6jb2Okn8kSvJp/ylpvTpxRNjnD
50uvErGYOkN5A9xZbZ8n05puVdG84mr/ilLatpaCz1IS1CjBe17kpVNWiMcCZ0hmke1e3jzgIh/8
5ai+P1/riEGaJlZUiOhMJ+xjTRIz6+gMdUc54kKOEvQ6XmOlfbptxsf8O3JNxCr2zmVH6sbhIGoT
tOX8Oz0QCxl+iWP2UP3w9ONbcvVUSNzG4315cvNLxY2TaUMQz2GYWpKqcGp7qGhwh2VfrKeHGsi3
wUV7l0lD4E8j9OtoPpJTK6PaKNjuZaBtzjr0R1VyhdoPzsv4tcnakMZ7VYxmOpcz6hkB4FVxP7yb
DeVbSMd/MIc0ObxiBVLjWwaHEAx98dclMCMjSj625hLJTG9TGgvgRAI0NtwZYJf7DibyfixMvMZ7
55JzS8FHanK7P0nD+ENIziukyg70IqBeMeu2AJjlWbWrAMAlSc5Te5bHJlQkt7vADsR0yuqAQEFO
tHcqUAz/VDMimvYGwlgvbXEsIvWU+O8bbm6Cn6FMqqHM8VJUu/OBZb87YYTVuVY6rCfLpw1a+cTS
zh3qsmv5PVwpOYkGxlBFiJyE9s/GFxmY+CixAuWYlGigUCOmHCWAOTR4FNhoByV1SBaVYlSmOoUT
WgHSrviXuDTyRjIqyZ3OI347zFr3rbgf/0ppqy6/KlIPeNc8T8XgswIbDWZyaCNYTJKF7awFz+11
1gCO8uUUiycoYKtdm2PjF5i/GyMzK29uW2Wga/s=
`pragma protect end_protected

// 
