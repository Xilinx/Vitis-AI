`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk7nu4IBtpiMabox1TehXznQ76DC4pemdJM9Tf10zTf5Sn/SFKsrXBtfH
CcVrpC20hVsjxwGcrMh8wnUfKs8eoCkWE7e7oPOaOt1gwxMP48zN4Y5QeHRSSwG5jZIA8+tfii8L
ANMDj0Ei7U+hnPukXWVKZhxzmDOtZmVuR6DNchcWQwQoGX12xuk+6Iak+kuS2vULAneSk/zoH7Sa
9LI8YCEcWkF45GttWRNzcZ7nXLlcY8c+JCtAtvwRolBPpo0nTTCjMqM0k3FiJ/sVN3BD040ikPxl
WpZVk2OQkYyilUT/sTos3s8NKh3nNoHFA1nvZXVYtimGoO0rNZbmxGPW+8k7JlgA2685tbjYksf2
MejTCpSvQPu2qN2ldnCCUBjlFAIGi4XLE6re38mSVk0aAq0u/kBVUT/nM2HXqh4N8GjdvLmMwqp1
Z5vSX0iEPsb42sUQUy1BFYrCJprBifex7Veu1XFkm2EaUMhVR+g4Pn1Rc7gFuvCApTrXA3INdRn2
LDuxm7p1DLxfMwPfTkEYe7vA7TZeE5w5QtiC5hLFWW+1oy7mrlgKF26R4m8hCNFRVHsq5BL7EGZU
BbSFzEDA0C2xfM23sEjrRff0KgnoHLn7ggQeO2sNk3XyCJ0ZEvMVKY+o2yAP8tyMZ08fJrwbS4TZ
VGAgTQ1+eQlzY04lcHTlBpXR+ZLbYDOHX9849dvrJhLnftajghptznnf7rGaTUo+3Dzndoddqooz
/RBkz6syOqupUKIZ1sx7QoWQcZIk00NZZEl2mNbGj0oX1fkmJhPvogxDnkp/DcALjK0RlhzX9y1f
8kmbXmDQUsJIQr1iR6lNc23tgE/VfE3xXeNTyMh6pROx4fR1MwkpwpYcmJKydvMxHnoAeNZVUCPg
nt/UXWbqG70OXVTI0mqTPNP5M2DFIGVY6No0YT/Do9QE6NRipe3ufnyoeQPh5srbuAjDhvxhFcRp
MSipv5UhpALgE3MdZWR05AHGTZbnIvuXAaC7Mjq8B4+vF1L45ws4I9z0FQEXht47DfiN7jcM/Wvs
dEBGoKL+6M0YXHNkLbhQg68htmRxOUK0AT74RjXbuyDXjGa7+v95LW/v5Wd+MnGtRAQvPFBxTTR8
takNXPIspEJFF1r8CZZj/0XvwtKlN1+KRpZ6+TQVhs3DPs3RO9e8fISU01ZdIRvFkQh68KiAcPXm
kvC4E9TbksaCpGoTOZbag9F9/SSHWAAjwrHCAG5E5arJbGRtAwV16YcbXsJJe6MQZBtdGBkdrT6R
uQUqhEsoVKsQP1+2atNTh3Dvrfc9Kehty/CmBJq0828ELW+zuL2LYTHPwhtTJogUaiXMx6+zDhzI
D/+0OIsboNUCbttIcBCQFJBaViOjP++vFXf38dyx1NZxU44s5uwMbYMZgMZ/7iLMkjTr5+fYurf4
UOU45RUYBr7Vkd42rXCEC4kIVEWmRHxVqaPs4DW4Z05u7hLRi224T4Fjz8aO7xSI65vL4nmHtIcV
+rAwEehNTTA320lnbuN593JAM3e+SEKMecxyFbAhz4J/orEBrkqCEMcNNHLktf7k7KwxUuGImdUW
Es5QarmwLPur3B27V8/Byv99LGxw6ds0dWkGZRHNhfPEK5Vi24WAlJyxec6ZW0a6I8an/pjaa5jh
4f1faJj8WzQb6BEAlrg3HHS4HvV+8JnRSfs2iyXmNaDAdNY7QgWZ3jzj7IOG0Q6Hlonuo33HwKD3
9KtKADxbNVV+MTdGrbLuQwrPOvRe9pEyhF21MqJxhN1wn5VbIkCI/bijJi+gRma+zrprJa+NQwUz
HPcvFoJuw8kcM12i+/I0lAzXJtxT1M7F/cfzzdBZGbvOlyfoPVmzURB0YDSIV7JsbjNOiaXg3y0b
hK1npHQqEufhKW12/9qPB5eg3X9YZ5jeCjr15tGiBgQmjysLMRzTOivGQedlb9oICxvYmmkbEpHO
I91G6bD3+HasVf0X+/hiRpbToyzERoBSjwTxU+O9eWQd80KeW2JsuUoCNxaSPVM26qu0oApQMjIp
wR746jqNEsY8+R5zWz865i4Ow2PDQ1NbwpeWRxrOi19xskZoAuiFikrm/nwOj+35bTeqpE57B/KC
grfEgltP+L2WV8I3r5lkC1Iy3uQK0PKu2h497bIF/8d99gSYdi3lMdjR+mLNvW3l4pMoOMt8PGHw
yKGHrqRMXWrIkCyamK/kka6jsL6285EvgHCYYEIBW+N4sPXSoRMIU1bOrREdfEOvIqa5L5Wl06Zf
cLiyFMIftCgdYYkiLuJtJk+10vMxgtwF5a/DkbuqMfjSSIFkdVgDxwzJXj4a2ahWyzDwU18zFVlg
S0JWSy3qXLsut9Ln4laRodJSHkca7ZbatM2+/3NafwQLUEy12L/gpqirxRctMSqzshtPQQSgBLjf
wWAO4HtHnqmccQqLyo/W4kz9mox4DcZVKjkHyXhbXWzG1wi2fyySLzYFfIue0qfidGWL2/RKTOqs
rkujff8Ti6YQr/V2a4P/kpowDg5PswTxJ+GwFk5kVeG2McZcQx/ISBHqP6FqeJXzrNWO/epownnH
ywlmpLeiNW7qFxDm4zXcfzCqfEyqS+GqJAr4VRncUWyw5F41KlxGuYrRw8kbUDLgNEIUPaZNjPF9
P5VUhEzvSCa3vxpKZ7/k53ExN+zlkb2F2mtTeD0a9vCO3uvjWwJsqpLx3BIsNY2zes6AngE0qkLl
iUIpGAiKhc2u0rYmFvo7kaS640mmidiLNMWwa3dSaJnUCihhX9CNemNcvVVL5XL9mn1/awlec7dO
s6tSvdl2+xgre33P9Q/NlY3ekgZlKtou9JJjtXSCa7I8XeqUvhNPZ5cH9gY9W8bGlQ0Ag17kmu23
vILZqznQj7AAJZyIl7/zh5ADSMe6kYHzeMdYapT5PgteziMaOMeuGwiFuH7B7eX0j1yy+INa03o0
gCIcPPlaBqpzEmOIp4639gSeBiwRu+hnLIokl4N7hiMIztiiCBgacup9s+uQi1sUWwt3JNPiYwpS
QHnmt8tjboOyGDpkmIIl8Lwa3X26LWJQUMEPibjITawOX0S22wTwrnCT3qKxVgCjSOBd/yBLV0dE
d01DG+/FxNJb5H07UA61szkYCjnXNGHMP0RFGqQSCMlnxh7QmqgbBXzCmBjcuogl3y2uiV1edOtf
nMvoK821vWSj6JvVlojw73MdZ8otKkQFIK1MpczH8NCfQAiWi63xtnHHkA3RNtb+2z69Ur5TjyFx
xGAXzG/pyoKZs9DXEuqBcrXXqfb9qmx3AqbY7MAnQJsLNXCvBc9ruGZ5WsQvfKtZuoO2t+rPaVkr
xJ+vJn2dXwK7PbToHU+oHzYKyOhUl4L1yWQAiHeIhQYB/o0zGg31917F4dYBsPxChnUSuY6TQnPb
tBzrClCs165twEqFuwp4zBjcPxg58/+x4Gtm+cRUwI9yYDmSWNjR5SmOeAJi3SoIahX3TqLYJ/iq
3u9LFn7o8Q8KMYSieinoUTzdwiOBobwv/ZnucpCHqHfU1LDOgS3+h1CiEma9gwEoWRnxhaZgphpq
68kmVpeEsrw6/jeh3Je0eunMTvxbzEUmCkkQ5I7dm0c0NLh3zpKIQnUrCUX5aRcajkjcj5Jv6Nd7
48akGrffgoa1GQYLnRWvtaiWO3a+30A6zv7JQ9Clnhi7dCFRctcm43qvgYtfys3SdHNji+S6kvdQ
5AIk1jcJ9Uut3T9RJTbliFXoCu4sXtcKzZaZIdBQQWETmDlk1MhHm+Bx9LjvvUOorDcaQiK0UBiH
re+bLY0/7WB/uqCQQnuvNutiZ2CqFArDkOlK6V4HSV/kB8ZYBU//Ya+RNhyEdqzuEaOaf/Ah+EyG
OSau3JQu3KtRlAeqyKo9LWpxOsDWchCgCDAuk/THRcgL9RfXWq4EUKD01lLXfHV+pjG+w7S6/p3Z
8X4TIc1vIAE9nvAy36aaevGj8k971kBGXR6ygaH85YUyCN7LMmcMnd1sRpStJQc5J/zPJjVYuZXD
/2Z7mvelEne/mX3ENBFChyF+YsTwYIPwk/OMwyQmlvq4pdvbcD+zPny6ks517NeFNokVcnTJEJ18
p1J3GQm8Uhm0kUyIQOTYO4kOfY7pj58YYpMBXVDsNHBybvXyhPkN9Ub35dsBGf0Jdh7F/3v6jqbr
31C4C8ttarAhwz6lhdcBpbplLePkLLyzSjmBKJ86yJHAC3TzoNSLA7KDjQCPrK8igYsQktmvSLT0
/zPtJLUmaH5bCFPAMdfTiluJ02+Ub+0w0S/srRAGPvuZHHttPBzYCLmq1SDdj2RJ/dyTPrFbq9VX
2onj4vf5kuoZxGSpybRtyXSmwzcHc9Vj1pEdzAS8jOHZLuTqVoFhh+x4BkPKKhLbB+FptXrNWy/o
b966mnsMkEeFBnD0hCgfz3hQ1pMxbKy317EQ15KEabVYzEVxOzKQUVTBqmt11HSsg+lkr9NptmsY
fA54K3TwUqLpXpA+7oRzBcqMKfPGH/BeaPObrxI+baD/pAABzkRiZV0s/5S3mvk2PvlL94JBFrXv
GA3lrvkoQm0gjiOhMv5px4cZ/eVCMkb7QJmT+MXJrzW+2g4vxIcrK95a9kHJfgR+1vV5NXt4V8bl
ZGFA+ESMVJgTiw2Jf2/Ez5coDx5ultCeYmr7F1nZlUBnaakBh5lWaoavrKfaGUlginaLmN50VciS
LDshUrEmsT12ZOj3C1XuInm16tKsRh0Vdto7zd3imEmsqcTEjzY77YA/YvDxPDyrWtMmENu7ps3z
0vK9fwDukLOzgiT2Jh2iRBCBdMVgvxJ6AvSlcF8LKhd7AXdOpcym5w/llM1gLuZOLTc3yO387LE8
4XvcjbJcv1Dod6bdgJRUfKLRJaHZNZ+TaMA4HgnOpSUwZVxKG4b+3/y49cE5L+krsSZ3i6859Bva
clnDx/aewsFpu9gjwld4FhyvTrDBkx3lSXfY5r73gprXdz7R3c6cjN58kry5AJFTy7eBAosgA9wP
uuGrLFl+/tghXTs91Oaewp3nFfDjLpfJZhAqDg+CZgEGCu2pLRltP4VqAMV9tTr02oupD7P4c1ZS
nQNyBbH61jXlMWdxDSo0NJdwF55ylgAWyvXjU4nCfWuAilwyJ3l8KLK1Lyi4P0qXH1MJ1ehh4//x
C9PRVS5DgOmPl69uTG6YC0qFCnojWRZRKsU3qjUICBUwLmPThF2m7C2JrRXWyGyXixgyqDY3u32t
un5N6TQCOYm5NTeFiCCxhhze/ltB1pWf7WrCV7Orc6SW8oj/QUogruoEhvmSEW+Uajos5KtZQRDM
6tD+syUcezkxZ0UotaIWxerQe7EXLyWQpRJ9EZqg0xxHA2Kxh2YXY5up1uWl+jDrLp9RhiLm5r70
Kr84dgdi2SPD6R1+OInnFBDWAHAZF09O3WXD1dYTwVvykq2esMvTzQgrgs2cU11n15g/4KTMDYCB
K8xK/Bjn/qiy6YEtyr0z6fYolZe/WTGrwrMnyRV9ZRsOvD7fdObQP2IzGAa/LEazcElA1eOPzbjq
I+CY5FESzmxbvyp4SUBQH3gdh4ubwnNFEeh05m1WCsfW4P6nLHaCs2BhyKvWjRCBA38XmzzW1hRp
VvU+jCyhaKlULZKUBbAa6VSfZT3WQm9B5qlYOvkajv93s6bClo1nTMtPnSrPG4AwUfBMlycvSpm+
l5Plj7DFEmOL9sGLnc+lBhbpARADbFoPNBfMtf0DvSzcvRsdD+HGlbBJd3yFW7suhVQaTDS/qEFd
qpN0ugThhxCA9yVYU0EK6qmFxL4OGaZKUoFODki0LImDnhjdUCdMw2LCf9Y2ncYdhtY6ABszwWIW
PmtGvLYxw0GI2RUgktBTrj6TMjIi+DCH8o6Mh6gREAb+bywg7zlVRdGEZdv68ghK5hjKENEms/AP
+WTDkTb1h0+5SnMtwhem4vl38SoSTNSVRrUoZk6+WVlk0Yg1uF8GpKly9ZmCtfR2KcAr0ZQFyAIc
ZhLODDbP5l64/CeebrCsbYFUtualg6nkoZKSCFMeUQA7Ta16XZ1x0cytohoqvhJos+CwHWgRnhIq
Uoj4aTVFdQxTQ0uM2FvG04Qg10LgPiv6IlLu6g5TYgS8i22A8Y6U2Bn32m2FiN+yjVlmQuXzYzDU
Jpv81g+YQ8n2FGdAUy7V17mP/VkWoEqhyRfkoYxE9b7XSsfw4Lyj/PGqLih3MrCDUsO1KoKF9aEo
OXWcYE/rAEZ7gHIhOxLaZe39nwm9mezLu0tlt6WxI9d8zJuxYDK2Ip7Vt51Mro0FHJ1+uNy73KeG
tsiTfApIIdMMZhV4WqyGsfQ3eGoSfgkiOBfrMNzamM0NezpDJyva2JDWXZTqJ8FKH2ELj5/mzqaC
Idra524dSCnZprphLT9wv/DpM9+8nQSH4oFrrFdeSmvJPVeMVwuC779en/xkgdIeS+fU6B8BxQAQ
ABWrif4HaxFlHgN3JGE4NtxLamhaiVAPBAFpxGI2JtXECqAAbPXBBcwlaBbmHmeGQir2cubAVAlX
jKzDmSNltBCC1d0GED1+v27aDzFXKalc59MvM1UBQl+Ma3q9lcDZj1dM9Y+EZyA8rCQndM0PHQuE
3MrR5W+x73qFWLSrAqk1Zz8HoH+3Yyd0pz6GukImE+92hnIQlO2fXhu4LynoZZiZJNmzhwHOmSfO
SYl5UoaGp+hAiG6Gbt22lqPSUezCVl+zvLIO5QV9u2W7Ma+scaeeY3nkxgaeRjwa8Iom9afoUeDn
K8lTmDks/eYgvUXq4XFA9x1+cIMyNtrBYP+qoSUsG1VFFJ11GnDf1EHk7du8IpsvlLMJ3CsxuFa4
zOaHyCjRFd5Fy55A65Er819cHzsIafEjQ4UewPB63s5jeX8ljd2BBQKS0ylXqfu1sQPcTzNhYXde
OR0LOuXjTwP8+Pioo9NDaSJoB5A/Ji2PQIJgsCR/5f0tOUP+PAfw9MQp/r33XnMymqKOmzieJmU6
Dwx88WlV88ZvPHBP4s9i8QF+eV0RnSUa8KOBr21yHzAGod2+h522vurQxfUemNAUkfTJ7v3veIDf
UmQ7OOQxB+Udv71skVXiU5iz15caXauEy3ce9aDJww6SHnYw+WgQ2prjSKz8lq+6zLdS2ve3+09v
RR1yd+8nsgkoOHPWlrTl68pIQ4UalxU+Dv6/oPYhx2e6NLemV35xymDnJmYBT2y975YHSE407TbF
MXoesv9tAjKcDfG9wxqonuw84AAylGH4AMNxJxNSADo0Dh9a/2Re4Fs8AUtrP677Y8Ogk8XP2pXU
Clj/10v6nnVcYNQNOX7J8sXG8/U1PD2laxq6jjxL2zpeqDATufN/bKncC9hb3nOoKtKeQyp7CsZC
tL6Z+2GebTgbekt0v19vaRqL2tztu3v2iTrF6uVLrkhE8YGBHL/EYgzzVOQ+yAS9wMrG+80s0ncd
Ca+LYUUtXDlW5C+eo2lX7K1s2W/EFf3uIXcSKds2XPK1VuE6tpbaapoGjW4BivZj9oNmLPFm5G/t
a9IdjgU=
`pragma protect end_protected
