/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1472032)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzOKyePDhxa+ALY+EYM3kanMi8kbBo+vLXijB4yiHLBya0SfbcMB/mv/7
CgThiRtFD5azOX806b+Mc36kAoNzqN5RX26FH2X66LgX43HisqzEmvN886iO31ABKv6A9DUeXsGe
cGl6/9ng9RpxiEjEtajWzkERImNW67lCGjFIPsOFeuCzHevHcOrfxr3Vow4gZyvOt3QiAv4LujL4
rPTXw0tv1kMl60ByYF3jzWYTY6JxpaCP5ZrYLFCz4BjjekgVr4Omczde5IoCf6QEwX08l9NyUpic
Eabdmsw4NSHm9X+XLRh9Akphx1EcQSgY+yRHg6dx/2hGZ7e/TBckvz7473vr/3ccGR+HSNxvOMW7
A2UL8QtRl/hGCUCe/oTYk1U/TpFiWw8KiDavxZuREPcSTUWq4Je1fseHq6xNZufXThiqLPoORpBL
bfOAMYxnezzr1xg19d+CjY9ncJYi/kI97U3fiCnHzxLbcwFOXZ1eBPYCipgaNuvfROWGrGci1kpT
1yuMdRIMqHpEPo4vt4oyNFg+XFrXQymq4xIqrxzjj4dQnJ2QqgFIp65C58swFLtOmeLCUQA7TLXu
uW27M6c5m8g3GJSXQy9mYQiHTwl8xZ0MRlDn7eOW5ZMafusarcraD9U7IHV0r3CcnJYvsfuns2gO
Tx2zFjOOjKxZwk10eROjJ1PR1zsebYc+meqaNPbe7HsJsjyDJaNOvv+sHr38DuBV7a8sMBwrJbQn
j929waX3oysge5GZIcIt78+TJaUYISqr0jwlQsQbDTPKoCItD3uztC5/ErQA/Q/uG39nc3KkKBhS
cqWNE106WhHYseXp6jytzsoodKSqtI42B6aveCU++//FLwwcYX3Bg/TNx5/DaQzYEcJwQvL11C34
ObqldpyhRwzH8Ry7WjqXMcTvBy5dSIbHV78mxrBgP4znDX6cPx0Em4BOHFDKQmjAe4WDDdBlG6Z9
vuWnndbNh9C5FiQOwjbtCi256b8NqWRCkurHPT691NNZwjW8bdUDX9xgeTHdFJ92eZ2X2URzqNGx
I5LsmBSBrpXypEuu6/G2AL8XhNNYBAcfdkvCrv6K3GoJG+1xMm8jz6BzNNnRhGdt/M9hZ0G+49cS
jCrwLjv33SALEpzsTusT2pB139Mx8ACvz/mUf1TYqz342yrdtaM/lEeevnkf3lxUTVTpDnfjMihc
QFy+rWlNAxm9tdfLC6hqAxDUslpbA9RyAqgsdEyJN13B2ZrCF1GZcPFL05NP4ee+P5KcsalSsh9X
7kpAUX+vAK4Zj/aNg+HwqCILkKzyx7OFB1Ee+fvfMkfgPLl5l7JvbP72L83qHzeEnn+QYqR5FPtI
mpZ8AwOzH2fJUCoPYSRzv2IrF27gpMvIgKK5MieBEMraPitf/YgSOkD1Pvaax8HM/FMefVxiaZ0v
MQgST8JbBH9T/8xVo4w6UYzgJChx/85xD7YjPEwtmauHNZneQLdQdVtpyO9t4fzg+f2s2g13v3EI
AxfFIWtPSFl37esJ+b1eCY1mLKrb7Wd7r1B94AmMHoSKJM6DyDiz2g7yBvUDPMfsVLrsciNHrEUL
iDR7k5R+8OAys6WQNlx1QB0IVckLqDrmwKR+l3XenCHIgFmNYUL+hirltYOL7mtstqhoTzHCswTI
jQqukjvwZJVr0+0HCPTbq3tKcGv3W4CEFzO7UmewjbulS4Wr1liJ6T00tRonqpFZpPbjNwWIyFV8
8QG/f38Jlk4wY3/bNDJopEXQKjfHgIjYNQBRG3j0mXT1tUA2xyU1Cj7Tw86yb4KTnM5quqwoFL4E
cBY8fRPQtq2Pi92Bv5cs2Em768bZrM67Gu2qEA3UrmprKwi3kpoEudIO8kEe053fvbBLO/VYs8jb
u+S0i6VM9uL9k23NyE733P9VkEEWVC8YbIOC3VFAxBd+s0CKzsuWp2KP4CJHWiC1PJuRzu1OhHQL
H2iFTeXW2n3SpiItYcFVI7zw7AJpXg9eG9WsLfMDRnSCK8SIUXrnwWXHoml/JaRWWZDFX5fYpMRi
E8iYZvJfbTjtDrQe8J8ViRzyCVBorHHVvzPMpwCPn7QZ47rnuWfh/e32PAr+gyarAA1xqrqUwult
Gh5/gAnyGQqiRy/x1+kh788kUZEBDLkiRrO0CiA7HwO1f2mYXI2m+umChUmnrzFavxIeMdG9mRir
9JAIpjsp2VAcpxKaX2AIM5yew53l3OOwfmE10YTsR01bGGaL0CoD0LlQ607bJsQzsP5Jpv6mOnZb
7hOUwBrnjZhtbNJF12NqFhf/E6yDqNx6+ywkEqTHV42EK1H8DWmvUTHTPkHHQud1fJqOuRmpMxYq
ER9WRvv3yZLl0dkt95/HSft2YiyHcpJBDcnE8rd70Mn9HUNxDKg7H0IC2M/G3qcUCzvlOIVQrlhZ
WHj6UAU9XxfxJmLbPUJVa5Qod0wYtg4BVyg1BOLIb4BxHqLnwwaNJ/jbJ0HhbEzkOMls7OgfNLkb
SHSX9B+9w9Xh79pgCHXTJ3S1NjoRAbm9RJ98o5By8BANdVN+87a2VFGv9Z1FkqV/UJpJfGJwgna1
EmcY/CO3Rkf4KVaAl0WTWDXGfesJqPsCJ8YgATDPkJj2a+xB8T9TfeTDa3Bg7731tnFjbf5KB8yc
tdaWFPi46lPKNs6g7fv7oK5Av+HgO17MS8kguY8b0yrdJPbTjPmOVALyUPPD/MG1tnp/4RzlcFF7
kX9P5KvKMCr6lTjbU++v7oW3S7LYm6tszS4Y0MgzryDRk9O8/MThzs+oZLOhNioZ0FuFX31UkMxX
38Z5rhzdUmu/gXVErKSnGHxLp2s+m0W3IBnVjcG2Orgiwl2Lea8j68WbDD0sehwRA1HAXnu9dpDd
+FcjhUn+uqNvprqrb3006+f+D5rN9mUAtmQnGSfPixu5DxX9c0OqaK3QphBrC+dkkj1B3P3xFD01
yaViLjoFZwF8Dmxa9MSFYdeFxe8nM24SM+v0NW5IdsuH5MmzP+Ufyw45PhxSf4hAm3Xs1x3tBcjv
QiHwnhqkR+xO0pVoh5rHGBL79sOUVSYHMDDOYuSRFqy1pgtID9G3u0+fOEo1BlfIxEWRlnWJNd6D
xdMT3WXJPmBk4J1xccn5Zp0LjMfaW0TkU/coYrD/0l415tN3rA2CFc4/xujphATjekqzvHKAPsaj
9Lw0TXRBgq+baqWSigOIVhvImOkdjZYjSC0SPiDmx0VVw0teJxrWrBHGNbg8NwMxlkNDE9bclPY6
bN5BBXUfdcXuSqZ3K4AV6k5bcAGDfYoGwiCyBJAYoPOeINnwHnnPPLW7z+CaZt+wsuHN4Ui5OfOx
9kxmJy1CVYJ/sJu0M3pmXw+CNTsbmaqljipUhjeQLm1ooOosN4Frh01y00xoKhfJ1I3sW3bKSuj3
QVEdJXmRjB52dq31t/EYdzrM1lAztYP4he0A0uJGdRTtq16wy6CCLmvczuNPDQKS8BYtmhNneCJr
J+5oz2wzpeUANIVzcZaFCt+KjcOo6KgYA5Ews/+xMWdNXxwnaVUB7sL/VnMFRaYXOguLbDApGBLM
EVTIH4EIDv/2ujxOhx7CI0faxPbGAK2Z+qVCZBkmAuS85RNA18EkAPSnlKeJ8ZNiNiPj9mVsXlaO
FmwtEvYyLU01+elSDaA6geC8XVYaO/Zv+niwalUSN7YEsU3JzRIFR+WWZRMGSu3A0hUOeIVHh9Lz
Ffxg7qNBG39l/5BFIWvJmGT3kcdSNBPCxsZs7IZgv33Ht0KzX1k0a2EY+vTzVEiK+RIojKLirT6C
j2OhSG8EnbxU9CwNhO+KbgDuM5v+u2l/7aUN809Z2X4GK4b4vu6WC5jJbS9uKxzEjtP5bo5+BsXs
4CCC7R2YMNf+BM3Jdx4GCfDBO8yqcTNwcsadV5KlnDLBywMqwmv1TmO+Ib0octmjTEqmlr1h8oyH
X5NaDIQ5m+qWtNgjKNrh8MlmSASugja0V9Ag+OsNu7sOw9cfn/veEYs+ctvwU70EaYWxb2vpyAJK
zOVC+Ka+eIVYlsuASru4JpWU9YziSMwerhhUUNaElFzCr4ZaFvZzc93VMFAymhgtXBDyMsR61u2B
KpzCN9nyPr4ZCnJk7rA+ynvJ8hIfxjMTLER89J+/ZmJzM3BHhjRj6Aer9h1EW4QKEkIcD50nugb2
tDfCG/RJpTMo/NK+oVEgBuSayyfyN/mCqmqVkDP+WwkoJgcVu1EPVK5Fx3oouyBhi1QcRPaYp+eE
KwZZg7ry55uQg9/gzNAE/vTx4avyK7StAnrtwSc8tS4PlaAy9cymBw+JLetygyPZWLEQjeWGIeBu
M6L+JBajOdtAxAPtjBydqFfLwqe9UkTQcUo5d4FvfhA+7sKfHHghn+asUmBF/EeFwOAZTJG+fL76
3V2l40HUpe9KCCnr4xUVtwvqf/YK+h6BduIVYT0XRE9dlRsuYwE5fFxuHeoRm40oDBZYEzmsA7On
Zk5rBGR+awc2CsOF1H+3JPYHfWcies3JgtDKgGaIOOlq0kPsHbMHI+fcPaKjlaKzgg2Fzzb7Y6kd
5BHV+2IJEX8h/+x/EtZBHu6vnPK2M22iksFHKAznfAMk5uC/HF9lPc/6zT0oqSxM8hMWohJeVttG
2qiZf0mrj0qSFrIkwAAzQcz90E9gTiDlT74ygwRpYAxgU8y2HGaW0JbUfGeBjibM86Cul/eX25LF
uIiLmwyvElxPZ9u420z2dIp7MgaDfBEJScYQ9zEQmAWXlf5xk0O5M6VzW4Or3EcvrlejO4wILXBc
C8FW5VCnFctRSeit5KbSqF2MIq8/WoMrpPN4kxoHNpfZPeJIlmYUO8MvEJyIIXXgYOCNCpvsF8/H
2/EBa8oKUdK6hTRCJRpgXSyaNheHC+nCnpQLU0aQWqZfxOCw9jXjbDIesNYl8ejv5aOciN8EVoHZ
ZvBO4XTvpsEkbpVGphpgM2squKQd8ohrd2eJz9ERaSK3dj7dlaZmxuOUr+UoYCB+K5HXAqbi6AKG
IXVPojHSTpnmpNLmVIH37pG39y/woq415wrCdKTSZiChp2zhXVxKxAkdkp2Lt9b7elWcXl+n/x3A
m2uIocBdEKxb9nPs8ucmawJ8faKQb7/5PM0M9lnfFX6L77K+ZKei20gxGW3z2okSYb+OpqdDHSUR
9vQvHJBUTUB4c3QgXHorVY0AS59DkWAA04p/WZEIqOXZSLUIadKWg300/t5SnRS82PCr6ibCpdLu
QWJtG2FFByngUgqKiot10l3NunTf4U6PTYWiSrt5NmzNqFlit1Q6+L1e7T6bKHYzlXqwszSZl1lB
Vn2WImWRcjghUV+lQsKmo5VR7W2wKYg/JhWJZqxCgUowoUbmWYXpPaUuVQzmc+j65MNO/KwKvddH
vyXGWjhy0sThkCzfms8hC0o+gaa/S0J2JCGgV+hpXT/DtgPKmYVGq5FgU/DdG9pPtGgGYE+cfVFS
SAE87PMcM83nFqcIe5kzDylt7RQfJLJeZEQNEb0b/swSsvw556KDIYrmjTm7wlPqbn2U5A+xRj06
d+2r4QfJDD16HvtHTCvRwSEPGZSkzR7nLGe0Et/7ZMWX6h60RNXgV91r/jwfRZK1Ony99sqpI5kR
6cqGKewVW70AxV7WFqTTLPTJSeu72nMeXHKMMbVlFIBKWWNVtIMb+jPbSYqy6CKrA5ev0CI1S1gq
+fPqEpS4YCAMVSL9VCHq1+7lcbWdDICbJFjsPSofvM58NC/HA3kJnQ1TPoCw16bYEPRcIMe/ktx5
IKNJaVSUZHSULstnWs+iJt4LXKrhBJ9jAw+ibZ47WTa0KJ3vTfB+8pxjBR9blOMjfZr1394fAa40
iVu+9h5VnYlWCwFba3NJncFVNWOMWLRbFi/UBvC0Ba8dEhzLHcKyeYqObAtzdi7ZSJDqQKJAg2OW
8n5uf/lv1A5Wnh2BAjtwzc07E/a6K4j7xuy28NFq9fQOF9Iai+uVED851/fHKFTAH0lCW+p+4sIY
5Z2rMGrPXRaBOdPI/FgB0uqvl8O8bBL58gZrMHwRnE2x2alobA0aakrGq1kMQAiBLrrLMjJNEa6G
YxBqdasr1s0X1nF1nCMhljpFTciNo0DpCNmEtpD5qDIgkm0P5EcohCFtvwm7+mMxYoe5tM4RuBhy
i2belYhoiMbdSJmR3iBF0jEH3GGjWgQRGoxyWFLoWDtfbMPXxrIINYriC1ZEqm51YnDzHenGFLyC
5q0lgLfkQHZpMs4sSWKD1zx6eERu/MMqXO8icuMTITeDn1SR7SGgklRM0hlY9ENz6O25pb8iXoCK
sfzQ+S0oOaCwb6A7A0XyfUhWVkxFVC42fgDMzheEHdsbSqTZCTAH9ZeoUKjHVubxjKHk2bBsPfXc
+mJcp5lOtSsraOVsiexzZLhMO2oi++cixMWed7aqKoks7uxB7QbWd4lgI/6DwTXaSsO1RsmkFXWP
4wVJnfYMmPAXwWUccm4Bn5vARY6KH++Q9AaHhONPd5D0m0uz3TdTMf631xgAtAASee8b3k513FzC
8OFqEDsRcEWfhauYH4jFLeCAPZENuGvNPQxdv1cv6Acln2gxTI3FS8JjW3idpGTmGfMb+FQY35NB
KU7k0GFJ5O/hXO+ooIFLSPDZ9NDaZBvS4cFOX51Ct4mYMEs7dGz0teeCNd7m4MWFCNdfBUqAt5FH
ssUCwqoxK55a1oDcWDUsxuTLxUnLCc03IQR0lIPaam/t/pVeg+W0PykfLJFW/4f32KThqWGHwgPo
py+EYBfZgMUedq2eb0BvTW0zjEFNMACrqJXDwXioO3jX2sTa7i0jqo8FHwuSphcptppdEt6llOY9
aG5WCtvL4qEy71Uj+YJBnI8DVfVxci/O0NCc0busSm3rpDZwNX8mViG9tamK67BHqnAGi5TeqjX+
Av+Pa3r16YH1WrQQgYnvAGw6QAAlb7looYl6zocg/MBlCbQDfQ3syccjw2eLPcSz9bqaHYc0RXiI
A7lIrrWse++J2ke7sm5iv+/WQNdChIggTzzSh5XRIn8nXgtNfE5eX+jb4Czgw/m8pEEQYjTsjAk4
07bbymsbmnmD9jZF5v2FZ4ocsgIP1IVKMjhY1da3cH7MjqcD6KepM7q3RwqbO6g47lMqxvMJ+gwW
Hn09buSoUFvtd77PuZO2HRE9AUq+KW9+wCyaPVBE6YLSS/BcXGpKnrVnJU5vhICnLw1YQSpQjYRg
inYTbleAq9dJhPBAJbwWkbefP7Yb8TviprBKmfNRhMAQazzhzHh/F5hrRzbYenN+3hR+jOsSgD4m
L3rdfIrBT1vbdpJ3eyvGTjxVU/StyEy8a2wrd6rP5L5EjaFH4jQYSJh54WiRWywvckPc6bfQtO8b
1osyGnXPz4i6OdmBWdVrqsLZqK7ctRSqGEBPQNhygjKktoib8Q5FRancG+lbBaSdBnB10wcBUBOs
LqmZAWxctylqvZpg6xtCtwACEf/Z2YyYYZ1/Qaf8SBqzEjZ9o0P5Yzm5nKHwFv054K41UfFwx7NH
QuNsRuHaX81GMLnVh4ACdl5OB8cOnQNwPTQD09Z1+7cBdXjI8/kkVmCxTbH7NcmSeIKUwQoBZOJR
TTwk6T8RT4IbudvJNmPOANb5vojo+pxE4yFavBOmdr1N9U3qmLsrZwPZhBp2c0AJaU7IsUEjLoMY
1wo6X6Nt5P5jdEro2ErfSPUtnFdyJxTK4oAqTbiZ4h7eeQlRU2kfC3iu86tQW91UJczggiqduV4W
yV9XaGR+cXc5LmDYG9+M0OfcAtFMUZeQjiX5QLby903ikFnKDnDRR27IbyHJ/WGIB2vj19vKssMP
OrbeCN1+NTlZd0RhtbPzKn9ByZarge81UfGAgrpvwji3guOeDSoF79j+OHag0D4JsOCreDgaSqlo
8UJPt8LbKZ/xJHhEnNVS+UezVcnaQBLLKaOFkng5Ws93EGaFgFHlaY00HUrCxCCx0+aZH9PLi+Tc
ozrb1Qu5KIHooZosL/7vzJGNnToxuK4ZuxOu36zqUnOKHURRlDvWnZvev8fKuEqO6RnMf6l5GWkl
YIA43LkfHlZqkycSFvH1jlZ/fI22/Leb4awI96om2cffghZqVTKtN3QWrkesWrbVwlOkqkFgekMv
Os3HC67cn/xQd0IA6q/uVakkUqy6cX/iLPqzw/z7v7iYMSJBhHtJli6mzBXL2wGYbvUxaAqIJCeo
7wZqObYyCXD/g3n98ZtwSU4sAzPr84Aneh4dWTg9KLG0wf1RSjgGVuYuV0SQbABphK+QMKMT6wnJ
eAKxS1+4paE9JQNVkbDcRNqReGWkqJV1d6j0jo9KDOtCPoWe74JJ8HndEk0lzbzd0lVthCrmd3Dz
YEYyhs+9yYHr1okOC9fDnRKVAjDbdVNcd1Zz6Vv9lJ5CE/LUNvJtltjQSsuXEHGr16pUsXD3NG1t
pPq8Ubok6S4kX/cRUiquKMkLqhpRannHJ8yLEeTAeAU3nZQRqPPnhDozTlDFJIushGYW3oRduXeA
cqXTnhhbfA46QIXd3WYSUDIsLaCZI+Yc3pNshewYD/7Q4eQ/+lVbykbbLovO52+i+LUOGtm5FAw9
sdfgru3dUbaXZurXp/NsAGlBok14vWF0bAP1myUSnVCyIJW3i8Rzp5oeNtSVQLeFsCn9ouVPYFfE
ix2cfAtPjvsz6G9i3G6Z8bpAGkCBf9KI5leZ41cM1fdECRl1YI2BG0ppzelN0K9FAlEtKqJyEvkn
TyjCLC3wb4NVaj2Kznej0+uuOhSwpFyphnW3Og7Wm9vJ9+H4pYQV/HokM8ZBMSJu2+v4g9qib5dO
CtAegYnTmKlGFcIrjVGo1TV2nahU60YCoQKusSuEGfuDENMaL+ToXGjoo6xEzD4mQGesz9PLlAzB
feIcndq+U0uxZ6UIARp7P8X+meiwmJJv65JIIVQT1DLGuTWsfRhWDSvheLQoyN/txK2OPDhqSaqU
wiyVWSW1Zx0ySf+ANJz3QZi+8/5VarLGE4eGxXmobt1JGKpjDYwihR/vf48WpBliInJI2LuDlrCG
84Jjo6GsFcWqOmBzkILop5tLVkEsJ5sj0JnAP4wjOSomqdHuPuzzd3iEsiBvkZk0bXOwOu2atelh
QpjhrqiIUXfxayCTAL/PYLvrr3tE3MZ3UbnOsgCBmiPmhlt9IuUfscPtT3BEQf28rCkVTvsjKtnF
vcDx+23jG/UV5htg03zBWZrxXGAqV++q4+xDX/nRCj2v01zu2rR/uXpYlyCm+Ucim6GrRApOYjcS
XDCfofaH8udcBZ5L69szdADCUCVVUUZ2QyehHwMFkeHw1a4Dm8jJd5uu47tPfcLLPyyVPnTnskLe
J+CaNkmFj93qV5AnaTqadgj9pvj918Plx/pLrf9wJ0WKQXbleLCHi+tmmipYKEsDxMQNC6cEl9Cl
GUaQTrSN9kQa2FiI0NWcEh/mvvUWqcBlgCr4ubL0sRAFQMrO7fCS+P9vuaNppNTwKJgssRncPTO7
FELMXXdG01n+cx46VNV8aNJebc/mhBV2tnSLOOxlHkX+7+PKdZW6UUlx1fNuu9PYz6jrBsJCL9UX
zHTUPEOISzu5Yyrlf3iUPkFfVf/Y3GkvaKXl9GlTpIZzMPWzv2ZhmOWqmmgl6ELyZpiq5M88s9Ii
wT1fPl8XhuijfOX8w85PeRWeRIVWlV3UqkEFsKwbIjd70P8gxxwkXiZDQiXqR7xhatfVipqwYjo1
oDWuFWAIIDvcxTEYdGMGiSbPwZE54YmODEC7BL4txH3Ak1ybWg/dinu43Ps9ScQoEDvaTOtyBPuq
Vvdc8/vJVqA4AVBCX2haOzn7oZcUuf8acKCNmY18z0/IyyTcpjeBf/AjjGe+AEqe+5FzRxIA9NYD
aE65ykK90Fcb9/Cu6RpQULm7xPDc4pDtgDWvsGNLhBV4lQjTDN7s2tZFtC6liz7zidi38mW12Kqd
fOzJM1iIh2uA2usv7eQNWyvkLKM5eecpqKZ9PoGBRyWj/s/srPI+ocZNM0UfMkwz407cGgox+rD/
R4fnpQ8IN4cefywcNc1E/HeVxLDvVVvZY6E/koWs8oLNsJhOz1h1N3GNAe9z474Uw1iR9X7bUF25
wGt3zZTBI/CDRBTVoFyzpf3dxi+QnlcappZzSkcqryvGwnLOSLAiAx0aFTRjuKWaBk+pd5W5s149
VK3ALOo2GHkWxCg9Y6F/5GOJYXWW+DYVNMqGRM6y6m9j82hcedc6TrQyggdMUIm33hNgyFdyHfmm
0Rn8QMayw+bYX+oUT8ooEKKEQCzSCt2v3CNpZCqVKdsubfmHIWObK9yjeKACDM96yub3tfyXXCr3
7vMZOCWQXEpmwA0ivnZZZihS0j/v1GmwABl38UoH/pojZUX4qHrtWQfLkjZfKp95BWuecpzmBTtT
q8kA7ycuNiFoECof9fS7v0YRHVeGD418NozBx94yDtNzqiZdSEDkz+/qG+eNO1azTWYwlpDK3WBI
g5u6lwbey0AfqSOcvbxutu5PcJaIapWqPIzkuHbRwscZF7fL0uSC/zlFTH9eQox9WwdhZ6mL8e/P
JpwgJDTHzBqW0orlrAyQKmue6+gbnGS+JC3xQHtnLWmUBJQT0AldChMGZ54n3hgXAKYXZVWC8DI7
nZoxTMtioaV2/qIiUr91U7HZ05h06pguJX1apgNad1S3KDcalPEZylCt2JB+dIbDgVHWKv28sp8o
CmDvgqFv4qf10tkkAI0uYG2NFEofOmfuoDxSAYQpq71rwitseYUmobvLtQ5saoTFFhXbydXpmx03
4KAU203123WKoBmgBjkkkRdJulYueSFd8Wu4rplEkDwTmh5+6SeAqvjQTB1nA33AddN7qK1yzFBP
OHNZX+pPHWd1tj/SRtjHhsyXDN/NNr2lBqNNyFqebGzPG65JH1GQct90WEcHbqMeQ3rWmgUsqrtq
GvQNFgx6dKyia+HLubJJCaXrXXm1qNLVFxQn7V8dRJOfdhICbUI0QQV/kUDJ4gj0VHdbjE93oKKD
WqNWlQUAqkUYLgifENfmNkpyV2Ah39ioGkJlcZkplffgJOmI6c6rOoFAx6Byhnv4wCLyVVXD6hOQ
R0lUls7Ss3LXbmD+2tEuVJPeEeF+gaEq1NAx12dnTeu1S1+/0pqK8TTqG0IFCDHCvkkrrIhOnZOk
yXP46ffkfUK54gnjnNuMV4lR9qBW+MztDZ+zMWmz6cEG8+FfJFBb3GImAQ1b0eDYBrEOABZFZLbw
LMgEa2cgQOTBZjg1pwJXbIHnyh1hqichklVRz+oUdAj+8XqrqtBWY0H+MXGu4sFPSsLEE8YJO82/
ddY21LfM16ElvPHoNaJTnE7DxskSOXG4a7Ljsi8Y5kZlG2wdZr1w1CvWp5Sb4TXNNQg+aIyoKbIR
Axuu30sC1vKaXcCcC52nds25q9Oh7pIQSftRzNUYLsKj4iC2FMMsUPSbeWcXaO5IBjGKt/+A8XEY
Tif/qzwG9WRVriCR6nZAWLTJ0jj57grxez0YnKZi5PBBdJVmLPV4Cc7PhPrw24NYAlM4x5480P8k
fUjHxV6p/yOYM4qXROXvK0bO/1hw11wfsZVijlh87x6Gj4f1P3RN2HtACO9dyKhM+rAGuZgpj3Ar
t/9F0JYIOTnsqd5CanQ2N4uwNEeA+Ud2T/rXDSXmTNPHATIdw7D4xoXl1e3a4Bc8lH9gpDcm1/QL
SiEnUf5Y3T1JQkA5OgdeDxYAnV7MNMi5h8UoU6RUR7KKWWUV/GmYXXLbaPiumr4IbueUyUp07jfN
8y/CGzAneOpXqr13I0ECRYpw0fUXzu94+O+lfTar+9qT7Ci3F28+l8FPGlHQJNkaxsbe7gWehgcp
q1wWIVnMH1k7YltVfxW+64tJs1XFt5vBTQvmfbA7EZvllp13Eficw3s7hObxjMwQMmgE4caoSu6L
yrhvxghMgTA2FAeNAg4mh2nt5o38qw6fcoGjODgOc5+Z7hkK8EUOCEYhssZz8EDUXAwJg2188iHg
o41mQr4LZ8jEhoVV2UPyqVUNEowd2KgaoIbzRRE65PUhhaM4qNgcgLKYbCFoAD0lVA6nwdZat+LB
KAEZL/58GMaiQCDeH94FuE6k+QJQR1BJivC6aLeUV2BTU/3OQBTdZXfC5CpROv1SJtD2mubcuXL6
rayKKLVup7avyW8WCNht/X6S8i/nbW88IqI4p7El4sxue93pQzJkfPrVhHKU/Myiy/CoG9NN47i6
ObyKwzjcR8gxYCggfs+NbVrnepN5X7cP8r/zmX3eRB3SRJvh9UpbiX26RrTqy7YxJdk9/AHI9885
P2uFRKYO3ButqUEw5hqsBuAJFsKn77YgmtdNoBEIhVWiXVJ2F45icewfieguprWMEWtGWcCIbBGp
DqJLMm89dMwWeB5gk35mpzfaKRq/ff4ajTKnqxuJaDr4GsuD8Ef6DgOF15HnvwFc+0nwkVTXXk7h
usTC586xmWv92yFb5SAzPZG0Q/YyoKwjROaDpAWeOUpsxMSLiyp2cb3/hcwMHv9c/C3WlKhegPGy
khQu/U2owJ3S3GlN0SYU2BWMteFNs15oGTeQZCa0jxLZaQ0Uj5OYk3lr5cMjklyRBnkqtUb77bUF
TwkfyWTKUKiA5MbQrAsvhc0AQOKQCf+xBXjaync7niKWR+1+K8pmC2ZDp9HnOR4wGw2oxQIz54GX
ZRbCNIW5HZzFEfWfGk839cj3ColGY8TjBnOB7UswwvhaJn8H9yvA5TkiBdes5yf/MCnOOqnLhtao
/BDa/u/55bV+qmNjN3SPUg4S0BuJfCTb3eKhHHnnjT8UIJ6iFsiWSNFD34+Sla5B1eH6FWwxvpSO
+6vHcWXBn0DX2H/Lros2lomyop5NhFYjrBmge3e58I6MWtsouz8jz7JLguBTDH8VU3Y+2iMUGHlc
RINONIi3zkasomPimAXlqMDqKg2oKy3xju8tbQj2/2eFw7ndQ9hDNM7NxMOWZj6DXy7aCJKziWmd
5aVGlgd1eOZPhQ8OXcRNGysQUG5uLezi4H/KLvmzncZZixYX8nRszZ46RZ2zgoWB6sckYtQVIhcq
cSkpmqbPR5goZEoN6EiQJm34NaIG/uwyZPsSveF/5+NX+qtyj5nQ01t3IdMMgeDEYc7OWFbZ4FIy
/g93/NI9ZQevBLz9OK8CYfSpyJRHUWMA6TEyg/FMl8pbGH8HSUE8BijZOoFikx5uUR1W2RfjaAH9
cDkSR6tEGhSTkAi1u6272c5wO1D0TgdTo8RCBiowDUqOj/XFzO0dW30JhYKQVxrfu3k2hvSowAP+
+mjkwphgj1JYYhBtjdnj8xXmbzne9Q9aiI5JAIaMOStYo3sdR34q2Ch0VQzjZjYb+sSuRyXs+/sH
ANzcO8bGzlgvd3qlsHEMGL0sy/HyqkPv+fC61MdgXbqxL1acQp1hd+F0ve/D9Ofxvwe7Z6zYD1ZG
M5QCgp/fo3NzPQzDe2vPzfictHSHVb9N/lvrdudrRCQnxyrumecbT4S+b1d2mjuVdGZTVvt0Xe9f
LNE5+yJtMpys7juq+5Cw5hj1WAmVAWPGmSshbuVdMTlTexeL8Wdc5huwGADZwgi93heWyePExxMa
iLsaGiTaQSSRMCpiqM3X2P2Ey5zzNQxUCh4hJsrFAhWk1Ysa3c5JBjs/ryf/Prtt6XaSPkItl5OF
RD5FhmuSpLiMgDeYHfaNgcSFtjiVFTmco99TqkhqClmZ6DnOIx0TeW60j6poid3L6jyEug98dPco
BhZ+osTvxzV36LbtZtbWOyGZ5m+fS6TfhGaka4xdf4iLPuNc7SsfsH7/JhrYC93Ag0IA5SIqlhmW
KtZxHyxnq8tm27uWS/EbWLbQ8tTnvgb2rqNpUBtdfPRM6p/V3fgNz7vUBHfhtycsPhsL3wz2/bbS
bQPMpYb3SNnaRa5+tE0Ylnie1fdHpPPUnXE28tzDskc6x4Pe1C6PWisqJbVz87FM0v7OLLfgvtb4
DBjQF9aIvH9AjEwUWIa9hX2I+baQM3BVlA6inB6dRskUPvZK7l93AVq/FdpBCuu0WqSGCKv+rRsQ
6VUeFg3SbFQqX9/qS7MXqMSeywIcNBhJN5sQX4bmi4LIsuYkPPxIiOJoLaYIYtL38pWIOp8JJBgO
QQqwcFffQp2GbuU9xlnfLSLHg3ezCzh9KZ2iiu/KPXRnrdzf/sd7ZVXRr6ngcxOZUF9p0MklVc9h
Xnq+fLTrcyMjj/JRJUE69mUtMgticgiVtGqchvnfEJpZ2Iu/HWCEi3NSBgFBGm8ma1w0VRhFTDnV
4Y1t0ItHmL0TgjQ+lPheCWtNJzSw7wCwNIJa9yEK/WTsby5EvIRxd+PYN3+rlLXDIC9FekdG0aAg
qdA84KAZ/KRHamlcj+WbB6Ouztquo3oOO3QWdFeRbq6BhJzM9U1KQbdACmJflIvgLVRLrSAmtbmC
ktVaWEuMJNcqwbkHL7x50R6PXzeS/TNbS1P/8reV/Yf3AAkO+SQZyrGRgteKWiA1wCRTMO2x0heh
UlEUoxF3oih3++OwIQf/q+dMRdoylUSTkHSag/Bre+iF66aup6jKWg5oHf6745uf3gOrJiOCgeeD
Oamdqxar741ffbHBpgm8syQpz5Wc1jk8oiFXmtQAXCnqTLcx6OTlLELfJM7hc6zXD1U+IgeZa7Mh
psbbPBoeaEDQ7yeex/WLNX5tCkbMgyhqhXECV8Zdu3pLC3Myf4T5dJVDxITa3zBXzn5vQrZRpsuB
2uujyRHsuAIAR3mx8jGUtX2DMVoti8taRPEZLv+NlR6it+yCi8GSPVfJ7UB44FWj3D9Pu3c8jfAY
4HrzrHbpR8y1N1JdukQXDvNxiasdVYMh85pLr32nyDZNHvIHjvcLVkMO92ns5fuw9r+FtdoMV9ke
+CgR0MLii/zFeVQ09sPJ33eLK/28vnXnxGj3v5iPioNa7HLkEkbK5ub+sSA5RN3NBeuG0SIIroZZ
dZED/A8vW0dxLbO77mJ1tyMYxeSPLLQqJQ9YDyRn0LfotY/Eq+Ab9hQA09BzMs1cfIZUdTo0H2La
tCI8+NN7o1OLfJBNWbYl7Q0R0QDH5YIa/Ws+JRUaQ4nVMuKQfUVqTWthi8rv7Jl34iilqP3pdVnH
QowQGDacm48IfvWCKD/TvymPYLJ/MR5nT9VtGcyBDnnko+eTDLNtR27MBkj0aMD8K6atqulduWiU
XOz6/rClBhOT/CzQg94TEnoPmmRQusbnsHj/y0elTd2A0rZ4LP4spPBfpp3pZp1Hzb41s1e9cMXt
UbmmDc9CBnNQn60jp9iXPagqlx+S6m9o/rWdL7wBeMPVpPHtThbVr5n/4zDdtGN/ftiCxpDHfBV3
RIlIV17hmqP0scfLDSVLFkVrOGcTn/5umStXSSo2u26s3BKP2Xxr4orIo2UPN3b4mnl3bkKHa0fF
ujmVctDsJfc1IuY7NS5QaooqSOQi1ETyA5Im4GwL4LTCqTUcuNahAGbXx21mufjQ7bwIcSliM1qO
MmPc6hs1+Kpt8/hl5Nc8fkP+KgqFMm4I3uppk1qsNzURnlrmds/NwdNpofARc6hu76Iz5aDcnJnO
Z3Rxa5fEfTZjO5Hp7tK7lLofgqqa4lWpSNLoGvyUv0JepS1DXTCkBIyOd1P0d+lsagO986Md2BNp
kp3zxS/E9UMJJMFrJPvJP6XGvGlyHGnVsH+pXXeOqOzSF7pyhtDs3/wDcNTZmw/lO7BbTWy9Z2zm
9zDh14kGo0Wjtnc1oJNlCuI2bscJwFupuIpsGR6UzF5EoP6pGrAG2ftAXTbC8w1SDllt4jS5z2Tf
VlLecDTNEmGn6+m444Jf7MvZLUtOZjxpqvlhzIDkHm1vKoghOZdDxNkYsBX29CcrOK2hMqQqgqez
NdtgotAiCf4dkX8/f/ICXGKgvkv9wqaJOlbq7A/HQAb4Y2IlLqUT2/DLqSQjiBKmLCx1yAEXcFgk
UAoQZwd+kWyQf2T78qcQ4EVQquhrSmR4A/xiet4QklrJkNXTJ6eNmGQHNrGwxr9xRrqOCxD4EqJx
FnX0bOve8kLUsEr5bXpfW7Uvv7Nt38u3merBp5KmBoHlUEExnlq8si5upoDIBwT5pAvXkHEScach
vSc7XmTWZsbhv+wj07ezc96q2UcH8ai4J+IkZyWurBJmSegIk2TewoJ6w+J7Dev2yaufJRUI/sv1
VS2x+rzEkLtFiXkoIve5U8PJ3XZMT4gBB4Dom05DqBmAQ+ACXAkowwUt8Qc8YYD/SMm8O2cJqkS8
9JLCAtfFDg69XI4qlK7RDkof4qUlfpQ3DNJqvNugvOi95M0Wv7SY+1+OYY1iUvkkUMFkbWTWO1J3
+7J0Rs23T7SGIDQMWqlWdpeikjR2lr3nWNegTwxX12BkSlY0k+NwyrXNRibEtW55bPNU6CV3+VzE
WxBu+gE6rMFnb9gUxMUiLYpOowauBvkN4p5F2n+B0f3+wxv4oJi5hGr3LxJjateQ1Zmi5/bPROvU
LKCWixkdhr4tpfWHwIIpJ3QBaGXr40UYHO41r46T+nuGfNim5//ZK6G03nWAOsVKWXvPJR2mXNZu
IxTjQjuCf9q4e5f/bfjbL4UPZIFLjtbP5O5+0bo9ul5SHg9MYmPMa+aChQikkXI5LYtlAsqsAtXa
Mj6wy675fxK4cfAglWnKwDvITOha645EtQCotnkGtz7HT+FqYOxNUPD0a/428vKsVXwxKmSz62ek
dTe/GyjM/lpFfog7ntX26dnvx+a2gTp7BC/3vfPj0uOSQnCFwpo5tdL9lf5e2ETPDuTtJ2/uK4xW
wFr4+QW5Lk1b6vho30rIvMDretgpfXpN24QtxFr0/ZDusK3YkAyqdPuCiPmedWh6j2vPUebUYXw+
jUxYLGkYuQQrhRPB8d/3SbNBoBALUYHnqdfNEfhg/IyAueoSeZnkag44roVsWCOPa49qlrdrgX+Q
7h/1xjtjs262KDWSuOo7GcSmVjh6vROqjI5XClSy9/tV6YPd39fb3FmFkew8xZIsDLN0BXbHZVHY
bhRnh+9ViKPs75OWtizMIxOXUghAC3loC52w9JT4SkcKq95y0CKQJ2XM7tDI/G85YAc1N/eMlKOS
Mj4DHQ36qoOM3eorEvWzAdjIp95OZqDVkGwTVzUgfc3zOHSzvg4Y3zgp7hfMtLCIr+FLG1rekoyX
ExOAhmc7Ns4qrOYIyI0/ACRYF2CHQAjD87kTFlIhf/cbxcjp6Qt1Ig7f8J+TFwcT4Dbhm2rYXHzM
eipR2Tr/Uq0y3N8zCfeV94d3S/rIhtT+WsOkE1QJPWxfLZrXa3jKhZZ8eei1GGkqIGqpaaDoXLIH
t/1o9NzEBncZkDFBNVdjMieyYwOydH7GqH2LyL30x613XUlHsNSAupI1CvY1EXc8rVFU9Wz0lNIH
RGTUi3UGJ6IFMwNJPwpm3uLxp1uIfEL1p5FtTuQyS/LGYPcyeV+b5t+Riy8rdNvc6a745he/8VmI
n2aS7D9wOU9mQONWUHU70dC+8nLWNgA+1vJBaoeMq0NMFOGvsFcaT1x3ZW+8EhHN0SMgecbixlXK
r2dY9PqrbDUqeEvQJBvm6MT5dUQkdQuILUQD5aQV/nhmethGHVjv32DBHNFksdGa4C/MAotUES1J
/tQ+XrhyUMnR5IDH+wrdEIpRDmSBWpkYEe9zGS0oZOm9xySy9NvrWpfJTGQX9RmfL6wJeEJ8J5bk
s64dm8EJxMImxoSyj45E2kRFQbfjtmQj9bgilOZnCv/RsDH0zOInykkf7ojI99uZCWlsP0Jldvvj
elE6ZbULx3GIxT7qJwarnLjfzEQPw7nSar2ZKoDeNaLp8RuZOI2Av2/ewiUCLyv77oXQjxnloZwq
LJ9VYfHl9YuPPJqpnzWgT2B9QDKp4b2GRTxfIjPQp0dujPB4uw17r6ZewqQkJOqKc4mfPh3zsvlq
eBSmCSoIub+WGJJfMLNwzzm8GpK1WoMEMrhbumwiL/GAcUxe1eHrAckSUSlHsJxDjPK0d0RKBREN
RMH81PCdi754eZ3PXDVWPyOltCzC2369sV4eFZoERDPcA9YNb5ZqLbngjT7BhKnweIGxPuK2NUkG
M3TFw0anuZZQ10xqlUvVVKVsnwR8Hoh3CuiGja71IhOE6RQ0NBtuOSvSV4fsKdp1yXarEpgFlu1Y
la5z7cjxnSUorYGpKoKofxg7HTsSa4upGl18pjVce6o/pfyJpoV1swOr9PMRSCKFTnLhsVfBvXie
nGdPj2OUwoyTC6alNUFx7UuXs/DFaIV95R87KxIBbU6GRInhrusF4pbeLyzqZyB0pzAXSW7RhxAO
eUVbGcMwfuF177ungwHk3FHokJMQESVbfZN174oYFbk76VjPcXLi8ek/PqaczdOh+52B+WU8li/0
UaqtgzhrWZQBJh+MarvTSyxwYux044qOaFueEpnBEPMHy+ozqJOU6ZroXY/cMikqjYmeTp4R8QFy
8fjjDc1ZXYlGGEVg0/GWYNSCYuB0cJ29IEF2Qxhs4RrKfCdaGTMZJdcWXLpsX6ij2PvVmufXcsLA
WzmdzoLeVsSxhwUZF/HmvTCn+C2HMq6ozMRBa5iU/fERaToiOKj08QMPbvtDd+7mSQ/5iK0JX00F
vaKYpfe/oejf1uEPyd5UxzDUKQaFysdGgUjJh5hP8Bp0r6Gh/l1EHoxrEAwEEtTjT4OdScjQ0oNQ
TdUGm6R66X5Qprs968z5K2Sl4N5RTHuf4zXXmz4RxTRf1cZLA+noypEUfirjeE3TbsOgvUwdWuPm
QfyCN9H3TjTj0qa0AWFzy3iKokQVo2MGAQ5nX4VO4hz1rxRSA5q824V3DbXTFbbECyfXpJGWU+0Z
Q4pkUyDpUI+n8CQ0H7EAk0Gn5wbokA91ugc8BRLjfiH/pLCv9EYgYXcrZ5L23f34yf0PnsJe4sU/
JrW5F4VOyhyZWMTO9UnBsPYiUtCWGDfmzgLyM3/Z0vhgvT/dYF6hdCTBwHdWEt3EZooC7D5IVqDJ
sencCwOvtp+8JYvgdaxu6AKZtjY9lai2JlLTdoeGqVzex1H+YNGY3zN7fl3F0gxTUjGAYlCW20BJ
i4wNrlanWV2Ob2b+MKQPJ1vuPPqFoHnG9+14FGqUTEzoqO4H5OM3NPQFyno16yHm6VyDL2iHMfza
NmIodliGShlrBU/84q180d/UhD+nSgHt/QHGtr6pz3asMdeBkOeq8vE7z5TNUFsyQllr1PqVIYs5
VHRltjnmrBG9pyQ1B7eTCyz7Bb3OVI/pmpZPrwiJd5Q3LaULwkEm8239Pb57K+ATcVzuqEeSqj4A
Jlx3X9uaRnFn3hY/lE4pbIKwJqCr2GdtAyhY41r393GlkvycLvuIHxFLHHmbVdB2o4V0/sZX5q+c
U7ftXaKItBVYbqyTgGV42v0YYWG/xDd2+IQ1duVKEMYRNinzGe94HMH58mmCt20JSBGj8pzkwI75
9lfG0ncTrwl7Eb61r2cvPGuCZsifgLXnc+eAt9rLTYw7gBK7saT+V80sZrHk0ZYT5LicUstrug4W
N8lGR16UR7Cn5Jf1uoHNftPVETG/3lhHdjhR2Uj8D63X188iLWHGxyX9cnBRkScqi7KRc255SZnz
5nX+6WCwOhr3zx6A0cEj7Eld5Gv5QcTOjLmEuao7zNB2yhlzpSV6ymBLVGt2Smq2kJfKXXx58l3u
NLb9BJ/xOrHWy5l9DxRDoQaZe6H/Waf34TD6TQJAwVtRBbxJn8s1uS7Gz4D28/dlOJjxd9F4rTbL
RweO3I44WHHHiFP3cgDVAJlYIxoh/Sric8I6CHgrw/DBvBD1t8dVuD/cOs+OmbRm357SkuhBmT+5
ZA99Acj7SxQTPjdtOzeggH4crYTpJYppkmoFW7ZRZi+FJw04BWwU50pFBRVkeiJU8+PwUCDB7H3U
iDTEQP/N1l7YyPIZAj3FqOmpdgoJb8OlgLWhhtN7hpAoNJ8osPm4dGkhi5nXaeJJTjxkR/BaoVMI
dYwUQc/eOpBtgdYFp71WuhhcGxdQAFa5Mexnnrt6sRKvgaI6jVso08daNTsVsm7gjS48CYQLi4dB
5ogA0GHRCdegKmd2Q4Km7aA44Wp8JaePD3q/ALoqeMcRdGR7yuFBH7zHvezK1x3jHaFO795mOCY8
KoFoSpTs4m70+0EnOgLBsZwim6wvQDaOVReS5ZAY0DEAA6s9LnYCSqjyQmV9lUKr4Cb5wfePGqQF
W3XbvmXPAhaZZsEK/V+gdd+7E0CteOb4G6ECQpV5SPJm1j88WMsms640n5KYZBV17fmuoCCaj8Z2
M9F+nVUVxUrfcIKiJ040EQfZR7H2J1N1Rt+Tkm9u1+wQNnm/LjBc8pg0ZFhpAkgRCQzaET1Haw56
wARp/h7dM5PdlwXORx8nVE471LA1OYavgP1CyeqahxZTuzUZM3bqisZdWwgULbQ6JXC8K61kaOma
NjXJLzgG1pAHYi15xChFNJY6Pa5cPWgMPKlHvsH5yPFTzgbeSeXWDCv8yI3um1RL7ghOzP+w5qcb
VGrZujGEdn+DIhgS7uQXKFXtEaSJZMpKyu5FJ5d/apAwRlmTZxk7I/olH3TfLwVQWHyTtpH/O4X4
9S5nedJMW4PlQuhlqJU88IS+yJNHK8aiT0lObxXjIcT6ByOQLq3ZPd3dspAS7WnPH3DNSmDscNLp
3e7RvH479nnedtxf+qOoJ8lQSJLVedHaNB8YzQoQdQ20il5D2yuuZsTK6V4/F4ihn9G4UoJCjJn6
c28kKqmnAOruXVJ0Auxxdo5Ww8I1Xr9u6SvJDH15jZZ2FLpIELinXnur77jKR17VOV+YBx4YwyuS
rNBK4+hHiQ5Co4gBQKqhgf2UTHfHuc1FsF6iLm0lxsGFIicckBKmErtpUpQy7uZ8YRJbYKavQtY6
l+fYvkFxoOljH+JICbRqgXRpzESkbQ00P+SMxsTc8MqtHlQrirv7hAFZ++eam1ByMzUUD0+8uM/C
H6kaq9LSmh4HpC7LyGRPa/EyaoR3TLNTOEP0nVhhX1ZIetSHcfQOKS/JPmvFx0QIG5UdxBpGJfQN
s2W6NgKSp6CxboYKvH8xbVvJMI7MPrMqzMUr6GZDBwbQnGjd5mWCS/0/XJuulS8ctwMxTYAa8tIV
fG87HOFENHDDuh/qRcok+NufE8+YaMQRUwOg9Au0NPGwvqGfODBbvrLp0be8VsDaTA84xB9H3E3h
Bbout9nkI9//6wGz4FgvuAIF30dACm/acN2RneMD4XKakwO7DiqbXE00xA4JLPyyfvf5vxvDDftm
WxxU9KraNBTSLxOxubjeC2pH7oM8CcJSW/CAo0GAHQM+7+PIfalEIfr35jR2uAAacMFEWNBtjyRa
I35ILOkAiud9nMZ0CthXwf3SbDuMb2eFdGgmI4SHaayXluFKUw1Ul61T7JvHkTPCmGPgcjYkFPO4
O064rKGW0RMOwfIjhMknZwruMRmvQmrnZ4rWMwmqjNvFpRmhf5TYX7u3OH6pVMfUr09w05rA6u67
QvLbuNGI2tdAOT3VLJhFv7Z7sdrvmsS32IifjBOOknwuIlp+ghQXPFmkSZi7VhcOQBVWP/3l3u/H
2bWDdvHxsIvJXphEnvH1SgMKgmi+HlU8nSRT2F61t52k8vU94zHv4bNExCe8NoA0b2pUeJli0SmT
p7Ithno4DHIZkxIMD9OPfGgAqwd0rhM+Oaf4OnbiNC7Vt1BuNsB6HLWqSAK/l0oukOoWUwpJuyWb
AqlxCNIlmzvespRnXFdz0DG1ahyx9Vc49iOp2K3wa8X4XBz8hSuvZyQskDjA+9BM7ewk3sD+CujY
n6wRb1OwiGqUTWjyXwuDBxyBYO4ICD+lVgLrDGoHcr97db9acn00moa6mZI4ZOMTVaovWK9BYSxg
r2r8H/Lmp6oNS035ILUfsOjXwDQRinCE6OAAh5qsVin1FONk8SNYBW24+iLZ+K/vx2qj2m+oK7mM
tSJsJE91JP7uxEDvFT1gN+jHle+o54FmrIis4EqZddYC7IY3+7YRFcoyt5mc0dR+QzQg1nkRlNZ6
Kd3VXtRCkk4ki1qBPI7nTHCcnuWx0BdDssBs7oC4g5vG9/MSvpld8c7+NXCsd7xc6yyENWv54Svt
+ZwFHUVqckzuuTM/ydbXaEvETiRMSktFfz6XaS7FY2lBgGQgEWAUNp4G50xoUXz3/vvedyoeBrlh
5xfAnJhDd0sO64R67/a/N1hWqNpxzFj/YCT+WHav4l3ycFNrys77JaI2PZlkF2PGxqRgr0sCVHP1
dYPn2REfJcqtHIc/ZWZAqb/Qob248bPWNGA0ea8KJf7hMvwyZVFjq8zFwRnOWiaF79RkuCGSRseB
9urRdLiBOqBsqNM1fzXNbJvy1Ys43zCdWMOLkxm1peY+FFlFOhnx6LDwRR3jy5SpxGm+41OGAn3Q
5S6agXa3dIk7rIs84S4G4HMOjziiNGXiwmZ8GxthFbXSOiDbymClRo/JD/tFFOFuuEFcWvdYyfAb
k9ewyf9B5g7HtBGKcG9/TIu+UFAaI4U2YQmthXAQl/G0LxjFOuFErCVLUEQ7UOhCeBNt+K+LRLrL
2k1qaKuRqr4/SaX1dXjvzoC8SC13XviufP6U7O1M6Rl31yqEGofsDksqTqq200z7FbMSRcYaOmfR
4Rf2hFlwYI16XL/Yr7HOMbTy+3EcCHyRqAXbFUFaYi4Wq59pCwwNzBJZAb+La9JMuj0t12V3VzJy
tksmHuYYbHKETJDRjlkXAj0pHKTY1G6n58P9wYZ9HKgyXvUyNei59cSUOpobfv1PfmP7awbXfOx3
hfkne3rYgfr7Pcwya/7W3uwdiUW2KiJO1sV7wy/EeySjgJZZrgJP3IxY3qJgORk8EkWvr4qcQGgG
HeURKtxZym9mmiDuJnvtOggAWHFgxq4qk1ZF4z8He4cF3W5O+5xtLEt2OVKz2sQFIOBH+PoejM2/
Hz7EAtdwUfTqqVDDxztY+kousSp4oIkyY78g3lmJJ1O0T6b/MIH2SXQluVgp75kr2j7/1yGnMibn
uKmuW3CoHoLdftjHgblokKIm5fvsqpgswhwLFqKAc50uOKfe+ao/Qrx1tWG9y00MLJ5TU4gE3bwm
e/WTmWMFxAGuAvNYHunz/pqMhClIXZXjhpKr7A14/XTBg2qhtlxxFWqZL13anB+Nd/nA4EVn8ZHW
NMWzS9LnDePQastE8vMB0zHgviZuv8eIew/WNbuPyW4mx65GJrZnMOcVnFItwInYMmQHQzMS5igc
+qZNHtZ+E5TKvzdkOM5xMhOBo4GA7EPpQlhqv0pvDNJ+g75YlS+YsW72idJ+6Y50wGS2tEpV+EwN
qG2K9pXs16Oa2rY1ueo9+lvUGiRuPH17HQLztuFbrmC/EZC0p2Oz22cuQfEURcXGnFFq8Mf45vyg
o2R4peo0dY4aXsqXHLvUWFrTr4agxk+4mRme1gf0oeZ1W8N6/GgA+h1R4zQCK4XQGlQeIe46qemC
/Hx+6li75lLoQRcx4BVA26wT5GAO0yBYaRnqSCdEENwcoILqQX8xZwZSysMPsubDhNZyo8xp7drL
wZf/yZlaS5xFaKWb0pphebhw5PyVnhGexUGfkYdODEsVhTPGVyiVbB+GqGgjLZ2j30g9X9NgdP+y
PJ+NjC+qjLYhJtPGstx/8E3HNcnX3rwR0UUDe2pvR5kKy0KYZdlj41xelmtIgC982WAHyHd8LGLk
NK/t9RXPpSdyRP2Ivs0pRRg082MmWSjDWqNPH8e2bpAOBW/PA9xq0I2t8KeO+Aj3ZnehSVbiOXj1
pnaQM7uRBUeIqZiL2/gbQ7kLnu3q8HfPrEC92DiUWHSNIauMkG0bdITM8RXokJfdoLSR/kF5RAvC
tzIU74EpjQJkaVrt09wFDynQso1nLT/q7AwldDlK0iSLO2EV7DZMo8eEX11G2DHXpvynFiIs+YVK
krfr92FoTskwuiv2AzCNnDljE5LmoMTwNDme7r7gJ5WyXRFQf+NA2YYXUF4TOkkb3cej/y4s5rah
/EfLPedbhoBGaHl6iRsO5y1C/aZ0YQ5YVdzhS408BRAdAXyVoE2/Qb1W16Nheejdf08o/BglLuOG
BXJ8sp2dHilBdqve/dCsak67HiTpkIhpPTV1sZQc4WRiakmJ+uFNmz73NDu4i75gswCyE0RsyKTH
VMuyR6m+nUyH+BCIb8UkVlQ53dGrZQbG4izZcKB03HRf0247t5mjbg4zi2FVU2u7AjFKkmZNS6S3
/QiVzL2wKO8o/faXtSBoyme8i19FTXjjAiGqN89zwSLDwfmdLasH8ygp36H4LuGFKo09KKwKTCzx
nKLLwoOt7NaZf+Pl4y5R87NVHSID+wHapDjWShYNw9hKAniAXbqxt0T6PGm06i9fO52pMInYbTbz
DcGgW06id5TjuXwTnaR5L1plH8A+m6E33hOBB+OWa5Nn1SFnjI7g/eixudjPDhkWd8xKgh4/rCsr
amMimqEt2a64R0L24vYE2ttMEtcLHIzngVxtp0z4mPaLQKqXvC8Qv3QJkOFLfJA1CWP1cOWWiPdM
8fPbt4b2B3qGO8JcMVMCDKovqzu3zs7XymV65WvZlrM5GUadvyCVVc1OR/5UzJPz0BsidZDda8SE
dp/3C0CHC0lw2QNWjFYw+f6hr5Tnb9WuD6sky9uUR6lPzYYY55co8+HcwzRx9sHYSkVDLimsLj7v
eozJIdrXQsYfZG4fCIjiUw8lfpcen6/MFQK4eo9Tz5xJGj93aM6w04M20C8sliIlZN7FCn4T/85q
TxUE1nxb99UC7uNF8XfWmfSviEJRYJnwTnqohJ8trOqkWh7GsRkXZYb1mqBhTJZiQPwHUCojpFSu
5jWK3BXI/e2sTg0XH1SHuTvUECHh46pPFLCFKdJX9qRUZH0sv5U8XCzoyssWtGV5vfvrQ1hpwsa/
0po4jiZUe+M5XZrMxjjhLFBsV1WcqnBrVjgXjm3mBCtoJSG0X6yeRG9lHu9U3scXrv9lSqZ09GTN
SdqHwwGrR6NS9gWQ9m290NK209x7F7+Jps5SUJxcqj/BFiU65zk+BMriSp4CDWCsKHK/yMAHS6b/
pNsQEil1sosbJi8IYX+YAHyC6odnpNcdfArCe8vNMV4AFJ3G9OiP2vgChCqJh2H7v149+nJj/Q8T
6O7QrjKYqc3y/nkn3iAZ6mUL/duxZe5ihxVLC8RwQUKFI4yc/eX1Kd7Qs8+pal5AX1HC4rlJE2lJ
PprT+caXnas5gWCCbYzJ1qUtYc/8EgbJMgWoHNFu5ovzaGlWe1vOrKS27H0UuQ1JbSZXVuXc2eYN
jklghjOpObG8AuiLfuJNF7lZkUW/9Dgi9QlMF875P/R5ewCioCI+qPd30DJirQBBMbdA4KQV6c0f
ceSfoMP645XXWWtDib2UwgM82ZPYkjTK2F8irGEGrudZvu3xJYAtMLZc2zXHMQLj0sJABEpVL7ev
aVQXhny0iot0CqzPmsdZo5Tl89F5hCabw2r8w669JnV8O2wmbqmy3E3fPjnKT/RYpZcUZYRrFQ/X
n2Y8JDsqzDmTR4wlD1bfsWFGwH0AIbnd9qP/g6gDo51NTPdtDcU+i2YQjF66bkOQWdnYKSEqylvg
avc9mktXmjA0ktekmNzcDjXJfTAhgG9yNC4n00laMiliZOkphLPlDELMeufwJrMs4oWrV/znteM3
fYwf51zGNw9MBKW+o4YKh0elfWCmlAq56Jafm5cV5wGXb6/PJpT1JVDIqqLmxgUsYAV160dFyErF
99ajqhViUDB1IuQjTrSto9Mf6y1eSVi2dzOz4QV+DDvvMjDRHESdh43CI0M9rIYZC62dG/r89Aoj
GFm3NJbzQVqGcwxW4ey8OjN7YOlnFHxBP66ldP9YFlJE8+CiWIB2hDOtNeThsvv1ZVZEg8IFcAYv
TeAHFzwDVRYiH8grL0SGP4nkk3LAVV90gh/WCKySSXuqeLEw8ehJ0zvMG8k88Y+wWe8tpYvT+i8p
0pNDvnuAm2b02HulEjwtapMlggkI7gj4GOPdT3ZMihx0mqSPnvF3Znj9QN/j5s1Xg+eupS97MDG2
Ph1VukNmZaagPKOnPaC+2kCTEKy9E+4i66s9421k4jAyW8FxwkfspZllS5s0hmhSgiTcnz02gfUN
5FxYb9xP7W523cvZKwm8yvoKJVndHCl3rXFZIO7Ne8HyBUVLcrfHmXTctwGjTqPfukDmweLkS0X0
m/a5adO6HCRT7WwhjenqkNyy9BJrVl2GdZB6oWTYjWBx9X1uEZwFAXEimtnnADF0aaY7FuKQuBXg
uKVQbr4IRyAzwfYmlsohBQnkfO/Fpv2oEYqh0wWvkukXqqzgcNH+0BY3QHRrsXCP5fVMqwF3Zqfu
DXvSwxaDccd2b9IGQ87j5MxOeeXb1Q5jLv0yt3SEfUPK+4iczdGBguV0TQGjNM5VHNL6TYoOOzKk
1/p1RC90JBJ6J5MYpNoihEnLn1I/q5vubXoLdfP0lSz7SDjJ3Qo0f8Za6xwLLLIuqzvHF8XkkF/p
8jN2Plt/MdsU1c670y1KVcexQHufIIaHZgSU4bUY9e2NxMHIPseNDSmV+9tByWPGXERFlm3ki8u1
usaK6Ik3yoXJOqsOToujKSq0kaf5UJDQvGrKgSnUaiCLo+UAYFXr2L0JBIVW06iVBo2HFA0a99/e
FKWSNjmzrCzhEqrn5VoRSkfm6Nu0e1FPEcA4mUS1ulMvsJAlRd0VcBatgwN31gbGBHKwQp/2YCaz
yezDZ4BiNsgcXln73hUEwV8IqevFc8MukLwIpVsk+dVNUAFmTdvoMVJU4uiEu4yI1bt/CXQBQsia
L0RZSZuUP05JgzjsUK4F2iNKw7fy8BffBb57WLfcdbrGkmcOfw1Eo2rCEw4IcrO+S9mNM0rPm9cR
PKo3cr7SgRE8u7cFBZ6G93VDBALyoEQ+Nkd5ER6GPOCJAbYevUeVThWrASrrhg+o/gxG7enzZxkF
SPolpwLMypdag7rKWZBZUuvwrX1WfxLV/rrU/k6HX4deXcqbbyr8fkzl/O1eQE93ZIwXE3iWHJP0
1tHHT5UZDugL0HH1mse/lCmN/tqwluvmHe6sz3GH9L1qcueG7aB3DyWCFYz/dt6T0Ki0/j5iUPfI
1o3ZZ8qupSzYtIJCpiwF7PxFcA4u9/YUW2P5846t3ghBeIDLMqye4+kg3RWai2hH9KQeMJbtIEbT
ibIe2FOGonN1yxmjqHeSY+GlRA1NA3t6vzr4r//EUxEzcjgTXhKl/AsNadfJsWjlxaKQS6SqwBvB
jJG+t8acHG7+TyR/bbqX457zzKvQWILMoT9OcfEJkSfDBSmm5/EPulRNsBoNx/qla/8qx/pdDWQ1
jvXDwVSZJrW2vD04Gb3NlEMrKk7IebK85k/gmH9hfJtpJvImdfEf5lE+3XjeFVt3kzYWVsKyxiYk
0BzKi/Wr+YZlfJP4lm7Av4iDHrqgmCcz9GPI1PT+aKbd8shjTZkZ097TFybz+dpFa+NJe+62hH0X
e4zL4ZP9344KUCiWrsmXs7kQY1gRYudYJ82uSq35hrKqqmK8uSZcQPsdt4z5gP9bGIwjNCNpqCFM
KznLZIROFg7bVgNSjUOVeZ2Eb1CET09HXeCo0lZvggdz5sR6OUTBo8KS3T3OK4RXM1aj+hizNtR9
Avvz/u9IPrldxWZqTOll6bkqhb1sdBHcw1ZoG1LUimCkx64L0L7SxpdL1XtZ6+sQWMfNuKNBjq7u
KusWyNyMQRHIaBPmPN8/qvJeFWY53OBLFmjS47C9kzrjG4T5nL1d/WLeiV6urbEyCPRNp7nz+qM1
SIQB71Lu1FmVnTpBr3C5etXPs0LRy/SZrZ/Q/pHo7PF355EWVGvDTWQxKwITrwCIEYAhn2kBWuz3
nEMdC7tu8r+3KJNIAbr72fXfmyZQXTkiSUx4+P7J43pF/thYm0QHfG2HvCmV86LQH19eg325mlWe
jYjGU5FmCLyMm//lOz25XWf/cP30aYzV5oAD/t2DPSW0Bo+3w9Rv+b4ivkXefFXAi3NvQs/g6fRn
lIiJX5sgKw6MThJoQaxq2ig92jYJq+DXmXtswY1nA5FiZdzntCmiAkZNvcewB8wDBNvxbNVJLif/
XscIn7c+6iMJA0y2G5ZrH8CH3eW6JcN1dHmVl2wNxNH40ikTS7qPZ3K4ODHzbci+W+rPNCFRuoiw
Ayrd6xBvvVaAGqWM0qp+Dtr1EA/79LnC3VB99ED644x65SRjgLN91c7bi5ssUySoawLR384SnHLs
ly5Rp7ZxHBitAjHHbv9XuQO0Sz7ZwH7C5zyiiRPjCzC57VEPHsABlUpKV58dmTabAUPP+dOwp7q/
gTf5Reaf0MflfDq+1BFADph2sJ5DEh0RG5KmJiPYxLk8mJaBTjUI4q6l5LxXWVfErigBfN7NU8XS
azDC2d/wxMVLXQnMi/4t/SywAwHBMRczSwkFh5s3RvSeMLcCbQV5auqqkLWmLhQjkiTqaGiM77FA
E1+5KmHXEhPWTR49aBP/5iCDIJJa/jN4j/0Kt3jHvtDKlXeBQ9M9ruEv8cvtGzEJz6MQvUG8TJJX
VVcfr5AVB4Mfk3kBXCy8+i+QnQ9Gh3N4QbjXRLYjs+xjLjqQ1YB5/xq+5nD3bORjhtNNVjVBC/Zb
9dup0GIwvFv+c4gjanzfFW169dwruuMqcxkgJX9YtU0nFQVRW14waX53MXAMxVdldaEohuhsUW72
1kqGCPZONZbajpalcUyxtNzk4i6HUzyYqLdq6hEpkWKX4M9NMXAymWItTIn46qMjTeromhBB38yv
UwoQlmnOtDKDhVfvwdeLua7LNeYGPFaQKP7EJFzMoaYOHKKU3BxE54kFx6EgTBkfnhZ+LkKztGel
+Pq1kw+4qQOt+ZTTcUJPNSS0vjrKtWyy9WapsKT1o78vEwC/oriw79SKanP2T7SlfzabC8w05BMP
ii4hucNdtLpyGjPKrZqpMyF/aYg/z4rSEYkewn6qH4ReZVbJymD5zW+b/HvekQjNQeqHFugVP93A
l7UNcrfxLZW8thV7k8bGDUatjBK83i0Q8+h7ejnQDerkRlMLLgBQWwkylVHbSlheqmtWHq6fszk5
xP1gr3m77tF9H86bF+ZMMW6hqxbU6Gv8kRxWYEfInFph4bjvxeJjNGWdmgHI3NUsbgobAyjvBIsz
+WphaADUMC0nHRQrE4cAFfLjgFhfRHh9J1YpaodaLOIcKxyY3DIBxLBGPuQV5OR91wxkJg7lFFBT
R/AP9umloWoGQp5j9weYmV6Hvk4O0jT86k7nXtBDwkMBLJ8FbL0XkN9KisuIWfWX3AWj4yIAlqbe
xUZa6TDr2oJEh/rilEXC3DqLxFfSuXQDxoL7uQdqI99t7T3w8NnRC6OocIRE0S0EbnONPGf/f3LG
emOhnoaR3Wk7dWMyvwfRG+ujIBRTv/jvn+jZhLHu5Vyyd6PptsMDlLqhjI7YO3grsotES8Gs8R1G
blrDnAdPfFs5s/+e1uOgn4hCgUP8vwKKafH1Funs48JnwxkVDtAxsWfP6/nF9d/EJjJIY/VQxbQ0
wXBFiAPB7nUjfsRUAwTu6WPqE+VNwJFyNVDcnLzcN3TrFyPGv15DYuJxw4padMLyjwEv5MD2NpMn
QZTP57qgd1hpCOQcnn+yDUPWWoiGTWpNO2HCSCQAZQwRL0UW9guxQ+V9rDGxa73Dxq5o8AwaAKlC
HYupuznbFD389qZr+Skjh5a1iUpIeHKcUc8+9miNXkItmSxM6icjENg9CXCh1TqaUhzNB6D+04G0
FoYLpZimzPgEk8KYfZ+WrmYvsprliuG312oKs/DMhP94/n1GZGgyBWY8DNHtjEpqTf+gtx6UjHd8
b3cEsmq2K4GNWFbLNHmdlyzs6NWHKevZBpJgjN2U+v7XiEkh7tejwiMdGOARAOrQyyuABRUh9XCR
8pIUQquE2HGrii9IgFk1/cSPv1niPOwjofPd/IdLahow1cG3Dh2Wft7GGjFjp6SWEKQP9iUish6j
VX0CS4H/dABSAy/KiCyBX0B2uRCQX1mP0Qw2izBGtyALlu0gPJsUHc1mF6fmMmKkyQIVl0gMfJ8i
LsOAGK2KqDld3VskeD5ZSxexMIIdlby5OmWb3JOvPmuBcpUR5a+fTwIvGRNzL7bTFptkwld0/8H7
KfH/nAbWSRIXmrBw3c4iWQpY1iKFZkIrQTPUfbJaFx8SyHsFSptbLtisruXVKpa70MvwMQm8ykMR
6vcYWa1NXQe2MnBpzHOqSc8Qzc7cFd08wkVsBae0oZnC4O3V2Hf1KOO/bFFvd/8Nc30N0uO3f7I8
veJKWlc+XwXQKyvcOYfQeS7z2yfKLKO3FFUvYlIN75BPFlu1WE20GJ6hcOOWOwVEwi40MCYJDDBh
GTatHjQk04EudmCyykFYLJDPug00JXkEdr8yCTGLMzHg5Da+2glCeWaN7xWaivrYQakC4wyUvXUk
2vQ6WlqtRY37Mg+gVsdmNGKb82WIt/ubwHIkr3Nm8Vk9cyPfIj8yaeXsehzU3GD8UxAZQQE0t6Cv
qbWSMYlqJvqjHCuBmtyscmfbyVG7IHAgE4CkdEk+RU2zRBGUaZ0StPrwUtxFEacF2LD/y9bAhqCr
XA+03VuvxOwYz5aPwfVZFEHDEy+Axe/jrOSRtuRtaUQhWhxF1EDUBG7mPdYQ71EpNkpK8U2cAf4n
w5FpQgG6N3rvaYSzEWJjuxQ1cvoFnPBhN3DHGTC4s25FK2vu4wlTBLi0rAkAmoxTLfkfcK0BmOCJ
3HPt6kWREhEPMjrU8D9wvMVq1CEpnm3EbGLvxtSeO3LYocaT60jA3HrbVi1hZSfv7q0yFGW7A0ZA
s7xf9A68ZB6jsnzIasQO84/8WfV47ysHYqId1MMILhu4JRb8MOvfpcwr5xk6KzPAJoAonop3cMGX
XN7xeUayjy7DfbW5DYxYuMCybBy8do+vKFl9wI9W8fEkQw9ED2EDjgm4XmrZAXFBrqT8GJzn1Ars
8pXy7hywqOCB3RpIpWATfuSzuz4OtF+qGu8uZ9niVk5qzuFlgyIAPvS1/keNtibSdM9aiPk8GYj3
W6h5VqlB3wYPq2GV2IaRriaAHpo8dCvCNTWhOSSNXlmpaSx5UXetcp8RZU4PsK7U5XWVPTTEtKYJ
t+AWuQRRbpP166UqSzfTcusUMzKMM0uMsusFXVSFGTgiOU1JMBjZCqCLl8xc3gRuR/t7q8yWPJ30
x+kC6HmZZMjS9OGiwNjhTy1DKgXw2zObUV544ginJ/EBaypu3zXEL08Arg1C0XtKYsgsy+oTCKIm
StyYfRICN2VlxY3iCeErpCP0ktdb1xl5hgi/qUfSkiRUSX88WYV28P7KJ/MVuS3WYcLjbg1Otr3N
+EqdekhjZezWRLr9nfBepa13wlgcffn8xm79z61a5cMl+ARg/VSaTiDBokRNk7l4aNaI42UbroFV
B9UpsFvFFOt5rMwCUNgQ5c3djhQs65sz9YwyFqFJdjQ9j5JroQ4uQCVr5XCDjiUACQvVccHnk5ci
Ee2yz8bSGdlk9N0waZdFx/3RwRbj3ZL/Xg5YxfeLIJs7zZIShwkhMDV271CB+Qp6bfndsT2f1Kod
wIAym7zH6l+QRLGg8hRI222F12hSiNQyDt8RCvQV7lEfjklLYTDCnO7AiazT9UQKmGdwAO6Iv/7E
TVFphvPhPTYnU/ObpkvDHjGwpFtKTwwDcLtykvxMjx1blK3sUG/AP+xV0vodROkeP3c+ibv0woUT
JjPZdTAyGDo5JGgXb+PaGCohNRXq5UoQs//fwsINRJkOFSNx50isVzJiNaugGdQKDyHaZiq/8Lp1
8uyX+AEwVVkRk7fyo/j4des/Mt4FJadhXk/f/cLGrdpgSYhO1Olh/4HmY/9IgFnTypJP91coJv4H
1NZ4OeyMNCjTexPa30F+4xbpF/cYkOmDBL+02yQEhp/4uATea0fqKL1dlrF+b5E71YN6eUJ9VSUT
8vzidOZ+UsWYLOEAfJsAHwmQfNkgfoPznowumIqWF3yrdaiIPXOTCooH2l6RN9BwrctX5zIdTKhX
4uHNAu0Y777nEuUyY+v7gmrMTjlT8lGBDoFAZczUqiQniC4OmBnoIxqsfUuHEctPlvzP3mEQJSm5
ALGn7PTQMGpqk66A/yULx0T3vTDO8JchIWVugV7xorEFk+9WWMnxMj+aI3WcrtW8UHSSqEkT7+77
lxr9sj0eKMk6w7T1allBjg1wlonhsouG0GSmvIUMdzQB0IqZqE8RMViXJvigcSbvTFi4hFqGLZst
KQKfn2qRDO9/VG2rQx7IzNh5M7GnEEuKAbdgn+IGZj7XnrjfMGlbnCDWmthKpYZsBj45JC7OJ3K8
prHCeJPPlRiE860f5wT7GzEg9Oae2uxVR8Zxmfktv0SqPNjjVp9h8QOJrBxNdrP2hhbRK++NAahz
lBtVJgMvL/2XSXUKZ6g229nZEfLGpSz/vGpGIsYdv5+bJDJ17Wzq3up8c+oXg8K08IyLJgD8Eymy
aJ8AYbyG17kaz4xYmy6p5HhXo2eiGJE135aeSi2eEia3Z76VADybT5OmKp0T13xveMgXMyB0k5sg
qjoMcPkVjwTokjKMdEowRqxPXoRsDsLTJDKk8G1s92T3+tgos+iG2GP6CrjxHVK1sTJoUI1YLiFe
D3qFGyHGW63JM0Lz5X3tO6vAiXBX8FMCpz8x+Xz9t5e1KslodqX07qouzn/ybN/wevRrP+DVx/of
H6+xA0jXEkGdGfZqfFeGbOJk48ReQB7GZ8ar91IY3P1FhrweG6q3Gd1ZISOwssJ+Ty2RSl8KNh7h
XYWaQ0vF9qfH2AYZ0gnSm2dYsL1bs2Fh2M2RTdliNfV1bopavwBrYyFGO8kSllz1ssAKzKmQ2oyN
kERpyDkbsPboZwOYYgFJOZ44i9zq7yRPyYdOnxc9/Axlk2+jLwS2gcB0iL+3cgjv8IMcUhVYuWeU
S+BrlV8CyI2vlwAKxMKwAA0QdJPN8HtuLWHXTVuOtsI55/A0HHIzMsaPmyXRapyMVvZQJpJz//JY
E/1/f2D8I2o6hk90xKcFjLd3BQyAtJ7AfTiAXTlQmPAOvXVxHTenn5WQYyDN6VyX5Bp987iBHRtW
SkO6vAefSNz7XaEL8XYwu09qnqTL8NQFIYaykUV3bhsbMQldfmZWNKzpp3yvqgNEN0uP1bS5u7pk
HPGHTibqxxlGdkRAdJtS8YoaMf83qj0Ga3jAKETC6HbZ2nK06fkKNfYpuIbIBEOA7kpMITNabIeT
hj6Ul2aObVD95nvqMUmH0GiGdShyfVSamxGSDVHPEY3N9kyPQD+Yj5LI9deGIBfH/u8FD6zRihMJ
WF0pG0sGI2H8jl2laGxkR8kU8VUEci3pz9vTQYJ7MMQpAy7UuA0+d8EPUwIHvGCHgvKDLdcQDyaM
ke3B2i3MTcDNucIEf2BOiFoVEK+1pj3JTtTIyTFUGMtB2VqlJ9fQ7VC/+XT52X6Ffhm8EmRJCf9d
sdQ1Ebtx0EJfYX0/vfZtASNeT7FJrNlp6b9+W1sRQ6zwCPn99GiVOYDjc+opaLKOr3MOQT9dqChc
KYcTSAyHAfO6JZ/qCGVivucA5C7LJB467JDTgugYrAv/S3EMxabcfYxYEAD77JcAJ34o4DEgf6Ce
wBg+fUfM3kDYtdPVfJ0MUkLTZq7PUGkQz9EdY+LeYB28v/qRFZHgC58K8rjN6veHobD6OJTU84t4
jycaaEWb3ZJAD2JQTB8EBumr61lHv2UgpOToX1PdVJuBzjsHohhv5Nf3uMkRJg2NeruE34fhcDwB
vZ4Vyzx5DGUU3RYliEv1FW7WTcww0vO+3dF7wChdY0yIu5LcmAAHn5PrxcEqtw+ZX12cUFjee3UC
vDNJorS/rRQVrAfAQVCCLgZG6iqz+rca/o4KMQ/62CVT4NxksxV97TdZyUWpHJydU0+n+hFq1P7l
heYY2eDgPxbeXN+AGk5xyf22Yq7gXzUJya8QaI/UhOL+xlIoOfqS/uYGYGfgt73gc53aHcTu22TV
yakWU6OKgd7cFihHOQrKnm/mDgo2hGC2DxXt6dIN+eWLKIb+pSGj+wuylWarZ9n5rAxM3JyxlelT
QnTk0JYQTACo5xUgKXbme6OvlJDvZM5R/+lA3PRXVq4Zew/6mVhGX0EGnMTuPsYjr6bie01HMx6B
PX/ebVHTFBJD+buYOXCun88zFP243YLYsB7rMVNowjX8G7AQBJiD/G5YnN5uMWuneLfIbzjVTpyS
tGThtY5++VG1FrHb3wKlL0MTTnhqr6cGZQM8YgY5XtiFftmjgt+GD+aWWbbbpc3efRAllBUkf1Pg
NpkUNmJqbqIgqEL0x+nlg6ugsw/rgqbD6eS5LVlm3dVQXyQMsk/CYwvyQ6+d/S2NVkggU17o/jVA
WwupTTRORTTN697amlRE+fk4UYhfeynIdW9TslJYTTtQNRoBLoIlTAkAIb7vIc12mu+zjVcn/gxc
fya7PFCIIqZ3XT2ViO/h/j1I82V6LOLIc8U87+zB2xeCZRHXg+GIoeoWXU4vkKoEKd5y8/ynrG+Q
GIwXkAgN3KvO+avWfL3bPOkanhI+NFMIrI0LQTTueEvm70bYlyE7PexiGPPld3rzzGlfYRg9fGUj
mLS0C5d3YjmbhHwFRi56w8G7YsXwxw9HtI6pW+8BgC7BTq4+7bg7GeiZfxKIkK8EwgEhEGUZZeBZ
kLaP8AlpG7JMEjwYidz7viPgM2366hK/2WRrh1uderKVJcSzQUsUgBJzYl+3319qeKaKgWk4DMoi
oDbvK/Ek/T5SW55W4DhNucWaCdtLbcVvwDSaySlouh2V0GZVmMGOTur+j1QC/6Y5a7OBF4oBxU6h
4bX5GEf585EptYVVX1THd9zQpxz9LdlAyuurSm1rxlcB9I0iFZkEbJLLAfinsJ3mGBmFwPyp07L/
ARNWFVn3aZFLaGeKwLEdN/p+4Iusiz6Jtkj5I866FSzM9NewJ5chAwoJJj0K/Kpd9J0EDjthxyJ+
RO/qDCkN4B1Y928TVlZs6uTn0/kSkb/6n+HvZ/vEI4pxGWxUmvuLekJmKqDCvVhdRJ5G5HczZmwZ
xXjoEpOFRFKXLJBT+QkE6u/ZkttW22b5GijHZ49nUkbaHGzw5amLAErwXkWnExebWpo0/3cjdNyN
zgG2MGGS6egzT5NSpFSb176giB6bpx3kz9sl1H8qKoPabScoGjJmtNQfKNVV7rtU5kgDIogHrCJV
1aIRMUgwLmK36295Vm9tGs0aSOPL0koRdTU8yaq8mqgiEdK0fa0DWeGIEjin1SK/E8iGkyrAhwY2
cmRnqBUIkiDDRw9fzrQxd3wSsUqhb2c0RELm7I+ZOSpW2WF85cr8TDN2K6WnbVAklcdAMlMn3SDp
2+7DAaqLe7SY1/jf8JLbdcgMmbv56uulJtXxWiYZOWXgv1gjGXnHQ3f3Kq6Eay8/SeSdIusjc1/d
CKE3+v3i6Ih9MypHNpHdWNk1+bxsn/ghIgU/eB+YJP5/QwWxjZRyPwz6VDFrATpSvnXBnJLhoiPO
vtgbw3F/J0SEn3M1HVB7goPBZUBVcqosxFdpj0ke38+drwcXpWn+YsHsIzjq06iCScrL28VedNX1
NG7XJLNzpF5NhoJQzZLty6fx9YNVHxKlGnuViB4u95s5f3uBsoiZx7D7bC47nRbzPTpTuI7a6IBr
XWejnrYI44DyyZoqlVSc4qBkXt4k05IzvTUuTfkn/7Ie2jiSoYyrmn6j0aSsrcC7o5BKjgMcDVeU
DsENijLrz7iyI5Ud7iDxXqa+1rPaJFhov7x5T5TKgc+bYDG/exyQ3rXSGd23qjKYeR49y+b4Orfp
aHzL6dqcpmFS+vkRK4ux75ih/seG/jAx0Hno5SngjsspDVftwvfaB5vMOxeU9IKZJF1jsNQg91RI
Hg+JablSgXnUzhrRsYfHqbFbQ0AW/3CQ/iZf+/W9/2WtYX/Q5JZf7UxgJJw3AEfupV3lS9Z7UFwF
dtW0YKKwZN7AJirC4hBCTcWUoQc5jYFcMV3WfCom28m0KGEOO7j4JYObhRxM5/LgpJiwYAZG3cXA
LgkeCi2CTEMLVwgXOXpXya7WxHSPN03crRGFsgPjmH9I3l73Z86qss1K1K1LCJ97aHCNMIJ85jou
Ie08moss5vCCqeKNspSW63kWmwaBmrkBK6FuI4sLiw3M0DULpsEieB5KxM53YlvR3Hnn7j8pUr6n
x0dFpU6vOStak9xXNcHUIfb0DQf2cA27QAiOxnIkQm/fnjt5tXUluQvGqjKRoerj8BCx3TQ7CDSI
pN54bbeYalrv5HEMTAxvLWJ7umRNzVE3NzYdBVfz1vVrvc8vNVP9rE6fU2P31lVY1OT6p51cJ9j+
LT/B3m0zilk7WJ1PO7Uuewgnlg+Rq0WS4xU3PW1CuEwIjb+XgS4lwtiKbaxuU6HQKhS8f+C0rSZA
TRO09aqPmU9MnhMtdzYH0bs2Rk+Y4EGFOjM8Oy37GyFNiTbwdaqLqET/ZMgVTXtehwnD1coR3YuR
kHgRVj2MuxN3XyaGGTFFoYfIK4F6OMfDje3PTAymmQb3VL5hdmheSCEMbV8O5vT2KURvp6faaOIn
f0mF9KqIkN/vYiKfY6RrOexfvjrRJ6+xZzwCoeTYqs66xADMd+jkDjSkY2W7K7+PCGn+zFhkYIlf
1vEjCpf85FGbTOYCNvpxABmINfC8HQ1qPzh97+oVgI8MlWGRcUA/Ed2RMpVh/47+9sVg2Yhd3iCI
22OXV2pGlvR7lJdtzb+mUoAnmAeuiPr1nwcSfYOb0A5pttJp0b1MVhLCmE1pBfmb7NQKYUAz8fK3
f4KK86fULwBUBPxuWKWTE+GHmdxA96KtJEANUprC5zA0PeCfMXeGWwilq6cD8pFFF8A5uyKF2umy
DcCVtVbWfAykpYgtQM9aRw4DkpqvFy1ZlW/1445SjbiDlqbji45snaCHybG921TNeIoJeD3noihP
sqDUGqfAPq5G9bbUcUw0OhwRo41QSeV/e0Lihl8vfM45cc2ee/WWj2R9o98NdUGwY1gtujmnFzg2
/b/0aqt5NBTiCEi1VwqVtKZ10lkXGOoOV5NIUi1e6Evun/9Y2W6Kzt+AaUuCPq4p++9O7pHujOwf
tmLfJLsp3/nAPmJNCPLQRBPDVPC0vB8+1BOJT1CZU2yj7bTJljw5dkhPid0dZKOzw+tjAKeO+2PW
Si4YmvAMNGk1WtBpSp8Lrk0ZgIAtn53nw8ZR3psyxdT3F8Re6EaQ8Li9G2brJXFF/2NnBn/gs3Om
u26LpPBbuTf4mAoZfXCG0FNzqXnHdD/iPh7xzteP9NPkXcIn9BGe0QzKGL13AxXUCgr9MBUuv37S
jnneOUkL59PSmCb1UzTJuNIc+BJrWEfTj3eCy0tn8+YYSbHNbmUJx2+dKxUnsCNdPCYkmNUbdlk3
G7CFEkpNqnV2iDyp7xO13kqtlRFBSyRkZr7VKwOyhBWPu79B72yZWVJ6P+JB33+2ucXxfJLet2WT
+/ZOWQOQs8eAf4jOtXa6JnZlgQcBXbZMs9HLYw4R1O4CEe/j+rbAmZBedPI+vFIAg4AA6LzRc7aE
JwodWiPg2IRO27lY2W43a5dwp3/rJz8ZKQfTVTAxhbhDrwYjxbGyycqMKLkYnl+dL/drEp9FP2yZ
wuRr7mlJ75A9sDfCHzT6FTdFAhoTClmekUGuZ1REy1DPs43CeQWQOkbOeGjSVZkQaejFchhyJK9J
Nf7YZhd80+Ubf5J3j3cFGMIv4jGUFKPSiEh4qu2Bfmv/1TY2HeVa4pDl5VXkLOSixs64FgwZ11yd
l9UYcgCF8FJ0jKnKJNh5CjBxbNChsA7qnmbmbFok+AKfUjreClQDpSPGQBbRMl2UqrhdxAyT6gjv
jg9bbQenIsJdglHUzq3ieLCEnVDzkPUIIdtbU/dbnoK2RZLFlSQJ12rouCi6KkUBuGpyXvQ2cZqM
ajjBUbqXA+zA5MWwnNknaNv96joSmOVBUSejqg0Hn6nEbIMhpTmebsQVNjO2Tc8jwWt9Js8wMvvU
vQwcrQvzTd6qshX620IYYqtHsT+iSvjLTN5wpILv40QTAVfb0s14M/uJfeB+ASw7R0h6L4TwvVhj
9gIdK9YeNTUHZDVBsSy40J7OowW7ea1qRy2HKPsr+AtLIPwAVAmaiN9F0tZdlTlRqmM705Boy1Hy
8o9q4cuK3qm7LDLO5I5c+qHy2TXxKZGebFdIs29iG5WkZwUW78cfjLP93tkXWSnu5W2tcxn8R4tr
FmY6rEz9vYzzmYVEs1XzJliecP+jKWwXalWRocJXQO/UwEssXjqD8DFodIXhuJNc+du2fEKH5Jgt
CjSPtW0JHqdltqVBR5EvgHPyPNq9SdCMY2tQefU36BAhmzcdSPPV+TKDIClBoeR63/8tZgqw98oC
GMV8GyT3HU7b4fzNOu1P5H0fR6ekGbPIzRJ4s3iYyhNcFn1WUWgknOpn+2mO2pup0V8i6q4Upqb+
0ZMYl2lCb5SjyCWQtCjfD+r6PIWDZdcIHcwAhkWUfGC/PqNF5MqaE+EoEqYuZSXTlq6FtL9cRbkP
FIyFfmwP3iMYyJFvFk+FqOiRXDyOGgjJkFMDmVI7bkxE+tH6q7ro31fKsoSgRiqDY8adBU51yt0U
+DrRj/Hiqrwb8MDg3wksdw2ZYM2qXg0GQi9nu5sZilJPSPq/QwtA1MVjEIxpsNHccqOE1o+bSESf
VHFJXPvEmqBo2IGs55U9UJRVyNh1soMgS8tUIMawnplADoT3s8C8aoHLXupnH5pFiAV8Cq17tOdx
ty2U3tI1IOYF2ZhOb2/Q80w1wFd9U6ht0Rb921OxNDLt2f25bmXCMmOSGUex3yaJlPiCLyrc07G7
h07TS3+ZAQFGWewr7FWeg0vF8Eb9H84EoECXUYjD+pWMQ+4sTEhfAx1mk5aWDJK6X+koZwIuFx2H
2Awa3HXDfLvZ5piw4tabGkEJngoQPnaOaZV5oWfI1zXjB+rsYiUyxVlZ+dQ59cS04PbgFX2+1CtQ
tMevBHm/GqrmZ/alwbXognhSFAzRNpL71S5daQauou8LgYSgOwE+X23POCHtYY4puhuM80XhGJtX
vkVZqc/IheW6lmdzc4KCX6nSisrqPpNI/lpjl9p+RadUMTrA80/nM3OuS+pgQRcbKMEJMWu9n64g
oUPdfzOwx1y4kM6FoQK6zsG1ylxlNJ9HMsyrAkBGUthH8PpCiNF7Zckmjndcwkp826dSGrAg9IEg
gwkAx8dVU4JVb2F/9Vm9cJVX/HfRVbToIJ1bjkiK+OkoGN2umpTHwaskzUMx85qB2azak319/e58
1p6G5csB2wRYhuYaSxQnmHCPsko5l+TAZd9xb+5isMFQjx6YtliHNMcqLKuSpipVeIayz/Ir5yDI
aKKLjcdyH2DeDiWt1OwXbD4ER4r9EWPrIAN/qjNzwFBq3uFoxpfUY550GchwBwKw1ONYQcFLtj4s
LlZPVPGHqB7aJ2re+SdClknr2j71mx9H/ighxq9AqRSY8FTDRQmn6frmq892DAhAMmnkZtvkDoC9
CnXJSSZA4mvVba1N1lkCePtAWiDp45Q2Zg5gmttQNMrYnOlkbHNlrneAOKoOU1dxOFsDHrZp9+11
R6baEF4mWAzZpmFCKov1+0uaOIMC9Ub4JVNjtZdCSeEMvTQC4cN+6f698p6DKQEvUztpJSaciWCd
5zZnITye8swklM4y03/l6YSwlU/EYrtqux8qjbBTNAs4FNlmYW/0KFFC4sOdy4NYIyH/YZaPEMqk
6EoKidnk6hzoZcDxOpY/Yr0vFvSm/v5VMtnL6PVu30ZJ7tcLIbzu1PNX6/6BHaNXEo7C0rqIoD1n
jDMnb/YxHrYjUTsUg0iaDHoC1suDwiW0UkTWZ9qEcq+piZ00iK5cxyO985JACVw9pjk9gYvOjmvL
36NtxbP4HMXb1r4nqDUX0cWmvQg38JiE6PbUh1vxszOZzSy0rgD8dH/MTcRGZM9g9YclKKtGqY8L
e1r3YTH63lu8y0bxirCzcz4mdrpJDbyigQdrEezssOowQTCRl9S6P8dXQ/qha97g4MHPI3vmiTv8
YfY4HnHBx3H0S9tHyexoudNi7XOY+voZNHSZniaZbs2meRROKRfc0aSCKu0sgQn6ogGmp5p8Uhfm
S1j9xub3hpnq4E7oCLd1NuPJ4C5pST9h0hUYVfVtu6sBgIHdOwewoO+AJkoajku046sPDIvLoRkV
hWpaMj5QydWNmOoUav6620vWZP9eqfZ2mOgs9o/zQ2ESlf3Qx2zXeFeHf8e5Zvn4X5dLycbehojY
9/5hiwMxHl9f1elWacm9ADT9ODxzXrr5+MGAVBn/rbgR1ENmXnFQW9xE8kAMOTrzkArWhVJeMKvH
uKmrgbYqG/DBJFXR6gW6m3H1RPuV7Cezg7Zk5viuixOeLuNB59m05xac6FseFf+6TcBIqfhr2YTo
iVDXhKQQubDA9ogP2otbIQT3LR0HU8EaJTkXZTcgEVC8OB6fhPcpcvsOF1osuXbiK7IMyg4/Q9D0
x4AT+ytOUX3po7mrWIKjiqAVwxwsdoeEzVA4SzoSD/sQqsnOjDPInxQEQWQhRGkUajX8+L4Gs1wh
eSxwmXCoV4t3FzmQaxraqd3tj4mP5pkrHSou9Kw4bhXua+XE5YvEs2PE+qdtbzwoZqJl8DjTGLQh
jSqauA3M67gYqg/aqN9e6fyUi9rv7ouD6t/QVApooF8H9kMBmSNYtbCl5aVCEACShQQ4XkCTtVbk
lJEaGovu0z+ZJis+ZzPIYdsstz2DR3VcWNq+w2w3shDMKn+imMXp4UrM10D7VUlovNaCE7uQbs/3
YcqbaOOSWVJsTmgXBYgxDGH16CA/EIU+YDXr6snwVFyJP9N1sOFp7rCl9ZCFKBJrmrBQGscDUIen
6+IpAOmGbOj9F6ZPhvMFUZZ0agm9pe9WI8OtjEnCZxwIVxd63KGKq7Uyj4ilL5v9sYTwyIg3GocL
2xWhzeHGQpxAJXQ6Hn+7QO7Nvjbr4GalboOtMmwWp1F76eiDE8zpJF/qU53ttsanUwuA3bRC4fgS
V6gCzFDcfo8zP2StrkovEbLzPlbnnYAfLgqO5wT1lYsB6Y/zWfl+bsWH20hdv3zNbFUDVrIuredh
2hIVERjQ90XtttAZ4nnxKiSNJuZC/Tno4eqWKTLaPqlGarbSjTO5EfOcNELCZdbsNr0aFF1/Qe7m
7kzljZ82agbHuc/SBuoY5Rc4YDzI12eAd4IG/hmP4gEB+wDgvGMejy8JjWds5UYOYeaJHIBQwXmq
MWiejzcAktC/BPL+mXFFGDA5SqgBFSQmKI9+WGxVzX9hUHJEv6VWUgQpe1Q+iLQZRuSX1Zt/KdLy
NkC8p6e0AGkZ+U10VOogXgFLNsvJYIAnp7WujqY1/TUpwrdXtMKnsWMaazFvG5Q6Z+gAywpGT7K4
L31erqVF/IPSYGimn+vMafmSaEl8wyzgh2XLCIY1ECKpXAVAVwRTzU1AHHvBcRNkZiQRbEpTaWf6
0TdTJPvey/IC9Dw0EVGsXPTbv6MiVC/Lqa5Br1EgYZndCfYg9tYu8dCT/p8uZx4bqz+o+y6HsYnY
PToBdsATNucJV6JVHEge3sASUPXa87WHVrOD+34WzSCUL4I8ufl07HO/QCRKvOiLp8TxEV/2yE4h
L2p4FIe3UTIJzbEJxU4na65FVCwvFiF4YHDEZM4nHhmWyPox1MtipxV2PIXD0g9uHX48Czf1AwOe
ejjY+igwUAJseOKLIOpzECTfBqtVwsa7erXN1ae9gMxPWnB20BK7aYozqbhVSYEUrt7bj4/a9F3s
QW7IxjtMrbqZMrU1IKQiu2pnnfjutMceFzZLk5bjPCZ5tvkZPE2N3zlZfSJ7j8GGquYAVGYSTjCC
wyoAV/FljLHYTfwgYz9s1agfQ0di4w1HmnL8Al3S8QnmGjk6B0Xdnyc2E9jeVBCm5OcGsF41SfCg
yuIXLWLoxNgvFNupXG4lXKn97LsIEZK2nZzUEL8cw8hkfbOkwxiM5n/I6LViJ+Wi/AweauznYjuy
tqxnujDl2nIBbGKIMRRT9Ekz70EXZztKcKLkahbf2FwIRL/I9cs8EpEpuuCBESbZGGdisfao64by
Z0vNT21DcI1Cs2y5kVOXZQE52EhBphhTPJIH6NiX0/zNOsLGYhaQHM3WVPcEfxsudFgzs/URviyI
X+HJgkOeUhHcGxi1swh5I3zUJDB34Na852pA9k+zaP2ue/pJ2mPj9nDvJtQKodbrQOApFOdpLrpd
/4YUgHBBdKkMKJeF/MOxaa+7FTmF8xMRLZKTJRg2me+6NkDUNGo0Vu68Sn3Sth9zUTVUyuKsJ98p
UUuU5TcNlfjGOikyKZ0RoLAqzkqbhDdh8isWCREbdakilWXhQwwMwE+2c23l7MIygzC0pCn5ug3r
nLD0RYRGeUUhRJeK55SNw6NY/y6ikSjvszfi9+XR01WSPXYvHNd3ugv8e3FxkU8rOucTeGEHngv+
rVUna8xiJm5lNUr7af4NlhL4U3vST0+OcK5XvdooPdUy+B5QGtfvN91D/ukZEsvsiwLcfwT9IjoT
Cb9gz0YkRq/1NZZAtGwBtTlYIXAW+FJRGzUfhIDmaARLI7QkHKPVHaHlRXvqKZPk5+JP3Cjd8EQM
obvi+p0a5fuWvvg0Fm3NAi8ImXdVEUlsNFYVKaaPei9LX2Z08SdqUSUJDtbKPo8PPHrqjXBl1x96
4O9Pj9NlEfjg7zPcRfXYMBcGEC9l/C7zbwGjfR7ecUPbkp5XPRB6PXgVwktwys/ovTySEmgMk6sS
ISebQQFUxqJG3+Lnr72pFolJg6e3UIrFFQsHBlcr9Mq4n4sRHiM/JhKiqcaQWbJqYei1TtfKvtby
s7apzzKMD5bA9ea0apKZ++yXcYnVL74m7skjc4oSuFPS9VqUKFDD6JySiokGhj4R4sluvLa4EmHi
qef6d3ecXUZ9+OtYc3RTjTdkPTWL4zj3m7e8CHHp5VMWUJj1RrQCjCudpYmv+om1AhMxelaOKCIe
QSl7uhDQ4/EfQ+ceGCXk8w/GwM0qkHLr7ukk4+G0gBNxq3Ks2bXGouVeIcjShPd+UPUIOspisBaJ
cO2Xnhcc6DtRi5+hzAdno1B7U4+xQgnc2WKcE/jFyyV+rtZoZcHOqeTjdR1lKJo2Zatws6hFx0GU
5yj2+hNWW5LKOGEuNJ5gxfqGJKnV/X0exttQqf2q8/gEkm1po0HLXRZBVbp3XC1bVgm8mYpZj+y4
rtyNoDHT+Z6DHdtfdHPykVmRLfmuMTvnNg/f/x1Vmm53xpY2SN4FghTFpf9JXHQUXnKsOFNuadGq
Wg2Yha7BEDgkddceONVLMeJJIVSdbxPGF+/Zwok/ieyIdklRdkit8wYkgcOLoW/+AoVQ23k6xuub
ZBql0EMaM1G6qkmNsFjR2UYL3LdD/EFBJpfPRZaHY+e8vwPzxjh+8UJZtdccO4WAEIKOmIOx/VM6
rqScqun0l7Dc+ndGr+m8BE5u+clTC0Ui1r+vRpJMv3+w4uGUVmB/ssklVW7ahJtF+jJpyTWncXFG
q1h7S5hC0hraMv/sfVmB2rVNzDlZ+HIqlnIB4a9WmWR1aSPCVa4fcF1pwoYirEPc9xw6gNpdc4pw
HJpR21OsPo8oR8SxtAMs8va9DSRpHqSUQQDVzHsQL1sUvnZ6kqxOCotKqEJ52k+V6y8meq1zWlUP
r6C6QSGLAXRrjqyv7mCKJesJ23uDKrliPYswv5Gc1A6bUB8T8uTjrnjocDYd+9EF47Q/s2J83AJQ
MdMB8HrRX7LXhqN1A5S24qWvFG8SqVBrkEld3WshSkuBwD+S1NzOWuW1chU2hukZIOkQ/R0KP6Uu
Ea2M0EuP6TYum8a1ZQhaj3V10iJ0XkruJ8LJIkg9xSzYPDZ31P1gEuCPRDTpje6Vp9ofhUo1pwvR
6SoWZsInlC7KctfncufM53af3jW++/RmPkDtMh1DgGkNozwHzFnCZ52E9kO5sh2jFsJoF3AOA+E2
iZrmTqREBw0hTz8XGPuX6RUZ6bXnrbWl2wsD/Kqo080WcYMgRRY0lNXwyWo+Xbs4lCiOx6RH/x20
0s6uqdFCEfAYVqUIUZJTshv9Yw0F2p4lr5nqDePRbApfY5d702ecEUHOM2MkKsXjnw095hbHGZon
0cawsXwG9AgoN6+b5IvV/yIOgNzmZZVkc6Fpcx8bijwZfgZO3bc6M7XnH3X/jKr/w0wZqpN8hvXP
+dV/MpxifK8N++u8mM73MkGZ5HUujmdn+z0Squ4FSGfkhGraYJc+/CAq/UFnyMzGyUDweU3vZ3kA
s187rsCYyp8QZ5ld8lhsPlxJvhifJ+91aoHW7I1MVJYyQO7oUEox6g1gFIOC8bcp4M2UR4vOZGt9
ByOmxJWbFGtu91jPvj0osi/ldvYxqgFrFNqmGZ7gto10NTyirvkxuZ5xhVTm6zBEnb4q6evm817n
0WVlflJKPT16+advwHFCI01RIZ0m14lVQVoAGFk3U3kKD+gj3itlsDo30CFdkAuMBLv5JoOE/pRJ
8E1iUcY+v5mGd0tEKUOEqZAT4aZ3o6mDuS9/zqM+x/mBC+PVvIQgI7dBSdfwM1RGMWe/h8z+yMb/
aOWeYSwp4ASwAq8nyjHgjzqPkC0N7cr4O6B7Uo3RCeP+6uYUsIqDLxP6WXXemDxvrTUBRjFpVL+N
YsXQbKWtxVatd7wGfY7JwteHxZUByFDGbBL7h62YbIpJhCWM9oP/xZ1mUmuyof9jT6cN0iVDaWYb
kxpeFOt7IMwQFHprzDza6h+431vhzyNVAdPkTbz4JLhbqUATkRUjG5t/DQyehfjbph0xtFNaH3JN
i8FN5IQZfrc1GarlabEUc3BObhYoxGjw3LrFdGyklvH/Jc/fspuydjvx96tp6DgN/gbGRVa92ruj
rmm74PGh3lIwPC6AVG0IC+Q35BHp7j30IJuYvQ3DMzGrKCR+ysjNLoAwXrmwHuvaYBs2v+oYPE/c
50fVRkh7CfUiMdA7p33VCU302zBhw4O4PgZrM3tyGWUBAwhpRmbopduhQAivB5VVEWPkQNDZDQXI
P2+R4bFiQfc0P+3IOAUDcnHrAzvtquCBh2wwLOdVUpxsxWKoU/DaBfNgNVofsGUBwaMwiOp14k9J
0/aE9WcCAeO1SrnvICQpkZs1QDxlSshcQYS8moqE3f5dGv8LcaukKZVxp8HxGJlu2qa1IwBL/cvD
KFNuAVxAi3T8K/BWK7s6pwY0+6AtrlwIJxqI61vb+Oczn27F7rqLmw2GEOjVSwKzZugU8zxLA1fb
qhVC29KB0sZ1lqFIQs75USL4bfBNOMkkIc+PyljPardK5lKrUkBhwSfTfT3V6LS+4UbzY8qCFHzH
qyf7EfIezkTAsxWciakXOYkCYfiLKdU61DqMGO2mA7fyUEMGJVbfLvkK/FXT9r/w6NsG60L1I+b4
r5LlCeZ/8dYrpC97BKjf6+txlZnwQx1iXXtg5GswjhL8gwkonQPKuD/bmv8FRgT7dmdDbwPISrx6
4miPCn2vwnciUc8l/CDpvtUhVqilLUySHES2YRyA7AmcPOLt4ZG/h4nnSOGftniIJs2sM7VzSMM0
Fwa0lzCMcq6C3jv8ufXb8SzdroRS9txgyZNzah5zHYxevUohKX9526PGGjNeY0tGPlmrIx5ENvZ8
d4tIpCRjVDf6+4zfbHKSFWo04ryz0rLwTX2plgz6+bYUe+BDOg2y4lTVNd/TRW3dphMp43qK6iM3
77TiiCINRUZJOChEiZA0/1jkt/FLu8HCaLAwMu9Z9o7dV74xdA9Py6lMvqflWhGq03BN6oBGx5zu
vaInH+lxgezsFn5Dw/YagGAkTKHwKWnMzQgEdhcsKO2AeHXOoS2pj3KDLCfrPsRRXWMqHt0uXeNC
beSN55zzEU6nBmTK2tdw9oGNVzxoDToeYSt/C8KONCFXEC9gfMoE0mKpbJTebjDGpKN+Hno3GpwY
6aJRNLjq7x6YiMK1exubJplPSWGozdLLjDyrPAzdokSDdTC4X/G5v2lF5Mnye7uWaxAzMaW1Ou2M
oMuShLoHrGRJ0N31GhZthJLm6RA4c1/80HbsE34mRnKFvWdVUm9fQVb+9wspjy/RDOWw9XYbLyM4
BEh8KBrIoW4ypUZwVNLw+wFKkrUoF3L2UPZL60Ei3HkQPmmGNS5BJcvph1vLqxz01hSVcdtRDJsQ
Udy3X8o4wqbc5SmED8rpxAur9H9RvD6aan64pEaqT0Uc1cubRYN9ah+uCDjdj/TeynZ8qmQQ83qi
Fy8U0ckzvjMf2Tvkae/Met+5Rpmgmgc6i33yRyDeouATuOH9c46DPw7b/uoon2gZt20TRRC6/wUq
b8z/XSpBMVV29rDElfOp4vMnq/BDRJtf/xUD5NuYQWTClph/02HyoCK8ChW1B7bPmgKspHKeX0ji
j1FxIDjy773mUA78vNI9J5A8578dRBMYpnJHQJwS2i2E406QFjRHtLVu6ZqKHFWmACGvJR2KZYcL
xyMGlUYiYN9ufCDq6pleorle2Fle/ZvKr/tZPue9Jy8G7K7waQQrG52IDF4W0L7Ih1K7J8TOCUHo
suVyESiRHiIoQxunKyJX5oktgj/49kot16jRchALM7mM0xSxUt26CkYsDho/P9cmsvwOqjsQfcPe
CssCt/i0lzqKSsm2oPy3LQoYrJKk1urny+wAt28I5xYPofMpMaNBa5SeQbR3grr6hW6ugo0rUxJA
/BIs94bp/H04X3ZADf6MmnjgumAf8PisGfoGkCr7PZPTN107s82dHeNYOmrcIitTWtUOr4UnuVjN
z0V8vx74qzt+i9/w36yKrpj10PAxb7edidXqb4TTGWHCY9wp3VUW04CnctDXa0eG0o60csosQ5cG
XuvYxSLeiSz0udkaue9SDOI4o+F2r5JIfvXUqaCLF7jdw+hyUr0lsFobKhqGuYfsxeLyKkaDA2tN
qBRHz4GpxVwaHEAvMd96Tk4m9gLXOCkDTBjGIghHPq5qKBcaXMNkMzCewCFjuiv5Ucubltu57AGX
BVClENtNxoyxetYsEKvLtK+6r61ZFYha26UXkoQjsEMbWMvB6niSe+BVvSvg9AzFgc0dlEftViVe
nVzCGJj+PAk0e55NCfIhDgbiUkAxpZuOS/MfxETHvk2icyu1pD9czTaEWYuOn089E/DCDEE+5DC4
gE/ChUJQajSpG2bkJ/AFsrcdBUdqBEbZRo5lSaNYKOvsvSmkseGwp92XMuBMD1EcKs3gDe8/Rt4D
HYIiXhG1cKhHqA3kBIVzjRzip2KNPcNXdSR8JQyN5mg6K5AMyJdcUugHMso9P9QtxG2amT+YTtEh
YP9sGaB4oZPTElgv2IWNqrSXDsvaANN9AT85eugLWO4aHFzL26C2PjHYI1gocVe4TJjja54rz/Uk
oOUxgKKY6XrGfHxTAEhceNn0LnenIa1urcY1T7DcclM+0rY6T7NjWetN1coqfmaWKkv4whwVm0E7
6j3DIY3AVvSS6Ia364MK8QdkkkuVWuOUpS8BKfQpmKdWVLMMlJuXPqgbEEdY3h3dvr8AbtE7UhPQ
JhCeeFaVoYOAHP3njFAqlpkR4OYLVcsRSlTDqLcVIE0XgX/RG5C9hDmVgjUs41lFPeFp+e/rGyN2
lMgyYZ+lTS1XyNMPpRJqh+pi8DFWsmM9e5RX9P8qiFl163+uFMHKOI46Qbw948GpXdKuPFKI6PSU
VYthMqdOj5SEB6RPofxqGdGKyDoiurGyu+LUr/RFCZGc0Fx4a6tG+3UuCljyG7ch0p7QsELmFZBm
I4B3KKc0X7y/Qp7idzXTVFEen8buvIrE63+IBnYtbgN1Slm4rIuOO9VBxF6+EnvPC6hIoJbq6JKw
kAB0wOhw2M0YYWR/7fCgYhvuZBeDqBSPb74cfGyJ+DhM5hhSfHK3+DImG5QWIh44pGM7v9K1NFLv
gg1yIfLJWxDZKb807wcMx3b+GEQTsb9mwGXOJWgBggJFQMPB7fKtpN+R8F8aEj1bXRdLXhTiMAuZ
edS1gO3YuEXevXmzEwCbgjBhx4j4Wzhgi1s27mqcDcP1FQy98+6gZ75ISK0/OwJ9j3rZ5WSQ6kmL
eNvmMy0C7pjuD8RUS2kOMS4Y7qBrRoDpcxGQp/RsoA2d2u8FfT63TmF1V5BZ3hsWLlZqOzRkBz/y
Uymicwi6Ad6cG9JyzdkH146NPtQ8DHf0l8g4Y7g2QjJoi5JJdD3Rn1DC/uQXfyElF1bYAAVqMnFh
uPFa5YcGRyXTlOTm40MvqdaT61bgbpQIP92+vuUgOfTPOIrXY0agCsf70T3g1FLFHNsSLETC+OfL
yALwK+Wv11UsiwnRYB6vVngORDUaY9j05k/GI6sAOwh/9Xnh1c/6O814mjWc3ZL9HOC7eHHJ2yQ2
XJvhKtIRjrQv34K3i4inUiKFCwmIamtJbQfSDBiarnjOtGb8A+LPUFr9ivaKO2N4ZRXC7HnClPzB
uA8LCP9CZksgdSQncR4W2rbY7dGOofQfKimDB+2TJxkAajXPjn5RZNNgYjCJjbdIA6KVcXt0bfX2
FlI45JWNfCAo+vU+mZ+uQgWB7RmLR4mv2Mc1OnIiV76qjeJbmqLjBo7bTn9krBDzLfO4j/UHGf2g
HgiTRwIQ1wH/V3Zh32/Ag5hSy1wGDLdLJ1MtyqNZWC7ZstiMSJxLubQ1Ydrny/a6eIsgzvcmldeB
ydk27TZUHv5vX6TA1fVSb7tj+M0LXIietsxP9sdR6Pc5mvNsfSWUE+gGonwPXphEnrmWJTrQP5ur
b1dMN0euJf6uz7LfDhvDiUcw/yEWzdHeQ5iJU7Q+6qz3Iyn074dav1KYYc8VU2/LXarundd8qZE+
aB/T0bxnvTlQ6lTQhy7iAjDFb6fwzkuW0wSx24wodjBeFVHB61TcO4V3lgzDOfDGgcRC/sDD3bXo
51bICPqwt0mpKVHLpNrVwwp1zj+N7yW47JY61Tcr8TX6FGGMw7cZuAH5YtWSj1BIOEE2FQcwceO+
kvy0p0jviItWE3XXf5G91UOCXhjyUAEP/OyTJ9dLsMbIVr44G6cJV7CS5JENrsWvASLf2ThTGUMr
4x61TKM5B1M/PFV6Eetokew8pa5pc4uVkEIxEuX7KZsj7iK2gC4r7tOMigr0BBJTE9nojNIi1czL
OpQymuN640KSdkBPrqOXMDW6u+IHRFDBRemqUDVvj4yQ51wzv5DMzWqLcx/qgvSkRv93qwU3aHLG
yHQy1RYD7bwODtPILQLb5iZN+sqi7iF3mihj6ue57Mp4HGQAajqvVRKKNuvpa6bQky4c8WoEvECZ
SQah3Jczc8+pblv5wPpbiOkdFMC/60uu1j6DSrTKpRSdwUCnDjwn4vgU5mmWId7zUA7eoPdZ/A7t
CQcCZ2tnNSWpKMd1WkVDaKKr9EgFWbi391kete/6emFGsCAG98fS5ETbhgsrgPiKwDYK1KEji1RY
o4/YHUwQ1GI+pDZDYvvsGazrSLaMzPAj75JjnfN25DxTj1Qnz3nGDLqne5jGjXrcZDYNexS2hReq
fI2iW0gPccAMDmoIvxJfHfes1ZPOPNR8/mSvd3D/OvK6CJx4ngPvFJ6nNGYBDP9tDYWCyQIEOXuj
pwWURQNa1gRRdlqeLnVs/tb4cwMHAbrTf0e0gV33b/DGLQx6S2lMcUT+CHfvEMeiFEIb2+FUUSKk
0/cotf9096NRRj3rM7qs4xYib1JCHc7PH95ZxxjDLFYF+PNscfwOnL4gKqE4xWVnHviDjryJ5Drw
L6bje3rWP21oEkvpqbwD1IXWI2kKAJh2iFVzUtA59BTkEy6I7v4ehrwTY+YF/L7eWKuEw3+vIOVA
B/8r3TpBiQYLvvHPeQPc046ORLX8joWhdaNj/bMLkIg7HwjaXBpRfztTPPLtTgtv1SRx/enKH53f
Sqjyd999Xy4XV4XkpQABhpd3skn23iSWf39ZmNLb6NIxG/rWgdxaucnK3XHB8g/kFaU4ZI2B+rj8
2fXwTdiXvaOq8Vj+CF0Iu6QZwHV090grZruvwV7pNyWxJzRzuDXZnOs1TxgcXREZ3n4ygFjDLlg0
jeyp92bAyhzgbYWUb8Z6yyqhwPDgF959BFl19SNdBEPW3B7u9X98SpdVoZ+vwCbO+yA71EB+49Xc
LiHNiyqmGpcxzaQosQYoPzbgq1S5wJEPoJ3gRZz9zIoI94ZtclOaCIzZA7HwKZGgTjLhW6E20L6l
Pbdmxq+edEXU/Fn3Op7H/lg1lctqqKtIXHv5HxUf1IAndWclRiI+bn4lzXtVUQf8fjh90gf23NW4
2yNclLQ0R99RcywgKxukAhY2U9nxDj3kon/7oF2xVPtwNL/SsqZ0aMrz07PCYaa4kxnJ1O0qP6RB
/PM0YzukwtMLVH+kVd6+EnXWVbF68Xg4psZ4rjxWVnp6hvPBtnzS8o7d6HuiHvCKYaAeo3R9L18F
miMEjnQGB3K8t55j43d91nAO8XgK8xmMuTJVM6fIZkmGlq0cVZ8Atdh8iuacl4KKshuChXGSGWrD
PtDnS+V86Wu93GGbU2qdoOg/z40q21JKvIF+REQx5Ce3CPoQe0eVzmoP0W4jvfPiYjUMDmwv49Rd
sChXgIY3XPb26li8p7qF/dxWcH088eHLKezkTqnzzZ0TRBU1Zq59aLS6ZgMANT/y8wkLY7Dd7r2u
iWYWjY+Zorj51TZXGzzVbI9Wqg9WgaT/YAm/Tx1IS3kAfyweAtxiVHbDWbXPB3znlzAfefxF3i0L
pCjAmF1YycaQqul1PeiSqNOs77FFp1PP3G3DgDVoXgV5YtO2npbBKsq8fjeY6PQWLNnU6/SnH8iv
qfDDJW4mV0YmZAYcrKO4S7LQYbLSW0BZhBx/XzdD6v9RDahUpzht7Xrqq7gUay8i7iGMrjTYCgJ3
Xl80hCwYthYmvVyiXofJ2H9b4TJFy4BWCShvqv3tujiAH6fErRAb1ODsbhtm+7Qq0R3xWK4uKHGX
YLNTlbJ74l0H7SpaGUoByUQrArRU3XoXilX7GJMpgByAjUeGC9Vs5/+NM6gSbDLlwsdnUNk3GAey
85ByhkyDNiwf7ozHCglurtcyK/rkiwtLYYehvL+PgdExr7QDCTIECCjBHeX7+O4DHO4WNQxqGtCF
X8RgcjeMJBHhhmyqGiJnjFZI6gtxf3iLzIyxAMCaAhIU10PMYJ27dt5q1DhtK6iFOevRRJuVdXFj
zyhkboe0FwjrWIOmp1bSs11Xkn3oKtcg+L0drkFyjQRDpzTJlkt1O204slPA5jtugjdr7c/LVNUB
jDRmSzPGGL0j/9WG3DVlvqMXfmlqDJdKoL+nBYLhLEfPXWpy0YJRb2vk/SO8FFwGIyVrxy9nbZSu
yqr/E8qJQq4Hr9S4UNVfpaCs5x/zgVlQ5kVGWAfME8sql+P6r0BK5lS4shnoS31rs8UYyYWsUqr+
/EjmF4JxAWZ+Oaar9G9tUSYwOOw3pxD/2yJtD2njqJybizNoLAYU29Uf7pC2wR8Fdp9A2VEofI5P
goajzdL5zCxkDzPTQr+cqyjYNItdigcuq0JjzjP5xJBeKXnnU/S9hCdI6ravMjdUmJK2k48mrLuk
1slG/e0aWK41Zkx/8h8RcboezoQaBo4nH3cY/gJes1J97S3Se4vlAFrWpjjwtlnZ4bv+0GwjT+P2
/7Akbcb+WdIKOG2c15Q67ZLH+drC2OomMaBNjk/x6CvkIhEhDRWtm88v0BQc77vT5iQ/1Eyc3R40
UDQycgY2tnO+zUvwiRo3cBPMfGp/pAJRzM/TXHVmS92fE4rXOeV1o/Jan3htlDgoKmgkIsFTPj2f
zr7/Tr6+oAeZU0Mq95U9vQw8dNUVTxmUbG7TZ0aijCKLEidNzYv/N9a1A0BDbBMubdDkMyZVK8D4
cPciFcmN1RJfQen2c+z9xaIDnSP6vRZdYIZfgiSgTrO/hF5x0A9T6MaLdX0+rTA2dTOtoOI7VLNs
ZI/zotrApT149jbVWJ0bw448f4pKR4YmAhCjXZTuCzx+8ju8MIgRwuHG1hbWZsxi3N97g9rsEoMP
hRGsnj/JanRJXvxsyn7eMhi2G4xmPxxml/pLJ2uLdHS1m4WPs1Ox7SIK6G7kvFag/MPaRmVAhAzI
NnIJ0Cv+RWA4Knd23xkYVw5PNj6h0VVVYZvSw7KaoXHd08cwWVZlJrwigyqXnlml8XsITf0LvS9W
3YqPHbcpxSYMFsEEZQERM99Kky1IX3SDYHxr9DTBtf/VDjQ1x7n0HFJy3KnexGDwEVysbAxGWry1
Ha9+QBWfyINtnh/eNa6MQMeVjmzA9je4x1l59FdxwsJgUwFDbPxzBYxU5OM0sO0OkuqxhVDWosFH
7rXGHEgRueDW8xz9VVSFMc+XWbWit4EF6A/gFvLlFUE1vZdIXT7R08BuJ77LucA9KKtZe2HNiETv
Rj4XfdGzXn3G+Bz8W6d01SXaDo1Qzp2hVY51kRhDZhRWI11BpP4fmqB0DZm1dTpdhcj3Ar2SqnTE
y7t7TfXz7LNTwK+Hi9wwRx2a00msGCt1W+V3pMDkFoEC+XkbyVrYe127HmqNqZIHPvqCA+hUUUhJ
XehbWXibBjkiQz/kMiSfKtAyZYGtA3q4vS876hIOEfXdpdJK/Wd04kMaH9SjGaVIjESjNIGVeDzC
oa0SBfsauhnsI4c8c8zKI2n40WenBezCvMaBBv+BFa9XQEaZTri+iMJR1fa1ju9Io4pzeI1PoPtY
2GOy5uPeErz1wxHx4eSR8ZSSicBOcj3EmeldGsRE+Tl6vZRl2w2fYNNaMTm4gyh1p5hIIxO1T0Qk
SLOi55PW/qBxRN9Pxf4Dt/JnG0Iuwz6knvtE+ElbIMVNoAIGhizKjXSkaFEUTROuDj4eEgsqeRHq
3yGg1DztdjNeABvaNh892dm5XKaozjBQApyGqUEkD4DIW1ND6vTD6X5hm0JuJftz96PBHIPqj/jt
oXwHwRxVlyDEfzW8WilLYx/OlECtlIJdjELuJcp84+x0FJ3F/oQsuKjbaEI+JNUzC9/0hQyneb1O
QD/uixvx1nOCFMz5mHn94Id9XskvZ5hlElgy+DHvn3n/Y4if8pvvKxz+Bj6FQ3dshiGxoB8xpyzq
rVjLvfGloA0wNxaUWor0QDbnu1gQL8xHPtJW4osdN+9ruwtKBgRjPL/Nkrx9fY6tuPHnozefeoZn
vDuVhsXIAf320U7mQAEKN6Hh9IgCCHm1No8HuDv3V1eA5EdXWpQreYkUp0+dd1qfynwDoDCTIVQG
g6kLoBzdkUhyhNBQiHr12AyAB9oLpiMu8/DyGL0JiC+RntjHWEWCeS9Z+jaOiEu9FJJG1Wu7NolQ
VDU03bsSVJPMV1mbLi4m0HHA8alF8ldZMEzxylZZKx6/oWqYZnhKdfTcgYAAR/lC7k/ZqvKTZx86
sZAGfPlPAfPU8OCVLXTRT5KRC+vNP+JbWzBT/x5ruAp76Zfy3OdH3pbk/RdSjTH9EM/Acu5DTHtx
LKaUNSuHOl0vMK3o9vzB7g3J1g3CZQ3wL24IV7TcKYXNwNwbPScK4FqXHd5JVIfCKU6Wjz4bZDEl
Zgl4ChBcy9/PNxeLW4uCKOyxdwC88GLZ1hsGKlfgL9Jq+u04TCYoiz+mY7rGInNeaOO6sgooMzQX
pAAfxxtCOsM5DJ/PMKtNPRbGA8yuRnx8WMGbLTuHw31+W/1QBTLH1UEIY5ROKBtQDuKrIx9WFECB
1DGmGZVnQxK/krEt1pCvDmbgZbJwN7J/StX3e7f7OXJOey2nACHP8txHv/g+RM2pot6RMAhw8T6J
KjSI3opwZj7JtOWJe2+TzSlT6wxtGEpoBhmuAd/tvxlWPNvzXUjKvVJqwbB7iCHOcjI/s1lSklu4
qulb4hqJG8K2WQujOs43EmL5Wka3U/h44B0v9Ky3Ay3HnufkjxhFzLzZv8iZ0Bm3j7fghurm0xem
QkNpp12Ue5NZagWa/exOWZGzkRfC7jP3IVsMTo3nsKMKuD2yrEiuukCi3gNNKK9XGZ2yVxR/zhEQ
mX4+BNQ2lV52uSpvzRZbUWKAw7iDH3pTUYqfDg0YHe7pYT+Gh9Yp9pBjepuYnBOLyJ49sSx0eztt
16nIwec20MamMNuBmUnUWm9s07aJv+BReR7A4DJe7qMGUZpFGbQZp/QOdcbcWLoBnl+JIC4iSOnF
vhoZxq/s9BagCbtUISBMgW/6N3TgBxgpOvj9is09gDY1Ck01RcN9ngJSDKoByvPfniw4IA03ZnCu
HpaXpfKpS7mg8AZL+8E2lMw3qO2UEjjAwQFalbkUOel1Ze5asMJx1vQmhkw38LhKXkNvv634I+KC
lRrpGpkuNJId8yfZpBXI0D7QPLFy8k2oreAduvNS9M6wSmXKwWbev8k8Jl7nrj6JNshmgineI3IM
xfogE9SKi0M6+dunNSUZJhEKdPtzxCeumBuOYkpBdogNeHTgE9YRF/kXZQt/VCMs0fS/WYAWQOqh
xcOUkkYlfYMpYPk094LI57EGyHXvfQTjPnugCndXBdZvOxZjvkbBgQ4CfOTsDDe0VEj/bX7PDUJc
Z31ZoPzcQiBbmVrHHy7P07b3v/0Fs0t/hrh0v6qhIVMRAgG4X5IGW53+6HN+aKUxPkHjEn4oLM+7
miruSqCRp2OITBDlCpzOFiSwaw8pugFsWN4iwckzK4hGLvmfJ2gIV+XmZugbJzyGW88+b7umy3tG
0Tt4x0IDtFNrZjooz5E7LCPy3lgg0Hlc56Qj+SWQXP/vZcXJaID+DW5U2OLgjyd51zT+tcRwqL1X
XBwDMBLF8WgumFQ16noLzbFNEzSJJa5WPxWgWFUiYZdwZx2FHKhxhKlWfcr7uN2fvXsuq6J8p/5Q
cxIYHEqKpZG5YJBlXCVviTURWpwQjTZy81F9aiQR5dvJUyii+DZZEGG30jnFJhMXo/v+QuqWMvuA
8fGuBdWbKrg83X+JuCaLRTdXxbaAl4UKSuFx8Z2am65fOI+mjRdrkXClx947oA/N2w1IFiUZaL9I
cQ2VrS3bX8hNbYekff3M3cUldg6uoUOOplSyensg7JKX53Qie1HMv6ZoXiOpr8Rgl4707dtC/oSj
dsDdL70dU5YBjCxe7ztnSxpCdTQeFCnCNCD81p4Q6+EGVXJG3VBQ81gsOyafnpF6qfaJp0Ebzmu3
0rJaotwQyksjtrJnF45KsFJtUsZu8D3lLx5fXSHLfn+xYTBDpeC8E/oEW6hxK/6ojJpi6UnFU29v
csBJcLob3s4rAoJ7NSdNU+g7piXjMqfTPu2+WJE1W2wA0AzAQJafcI8lW+7/6MWYEnSupya0Ighf
UYQ0iHnmfq4Nqh7gaUuFSISCR+USEpSpPV45Qur6GOy6NGAGaBvVv9ar3HPz31y/A8jHDj2B1gIR
gvNl/LGKBnu031yUY7QfrK7XnXbPYRmcalLPj/N8Pu4R/XJAmeO+EP3S/S9wafGVc6dgbV8TTPeZ
DDHUiN6HJOkZPzfv/Px/xWIZHnSFS6odwHPtp35YqdQLWepC77T/6bCs9k7X2CxKdCxepO1S9UEn
wv4RXj+W76/rZHqAEmXL67hOgcbuC10Z0FWgQILdg3FaT0wYa9WA37UTespx/iknlVmu4B4cFYlF
NsKKJVYnrGJnLgdHUwW1wOn8qdtWl0NKLqHTvm/L2wXSn4xzkUTzo40yJz8Ug8Y9JMyTjP5phwMm
vyafYQk4f5cgZYMqo0I3ZwNMWHJVK+rfPIj2E7Mf9dnkXu6YwYoheUVZ8C7llUUPZ+WTsFqqc5/J
epmB4qwC44H88/EoZwpJ4gkCm6uX7IPTr0GqJ4derdvGSFPUm7ahRZege89iSnvt211VgNzKO8YJ
2VFZA4IZSEH+2AlxoGB8TRRC9NZNNmivLPh93k5R4H1CemMhwwy0/05blERW8plGXepAxNy6jo0g
5SIHMWAa39/DGweQBNyHhiqlxmv98pexGe7WxCbWmroF5B749y4PsSlZ00t6n4V5aRzc+Ehs4UeS
IMZ1zGL2+f/w2U5R4zsoJm0HtXISJwmVArF2b5m7PdWymJP8/aOGe7ms7jD2j9kubycCdPy8x0R5
OYQuf59b2KhOqDa9cVloKxIaf1TDCsEAG8a13m7QMp79ZwKwhDZmdGJtRFNnU5fLd4cvxxn4hXoc
6sd8KONQjwojXhfA0lzH+sUVDK69w0+dpZB+diMuLm4j2gbbHyn/Xm1Z/kAfSTLjJthtVPGEepD4
xYMUUDk3by4GhuEuya+JfIRazYNd2PBpCUHhHJ6Tod2WvKoxf4377BAp/04f9xCdcDIASs8/P3ob
1bfvDmoMi7JZQN+4O07nq3eQnr97bIDReEWLzC2DGOORU7VvKJsBbHKmk7+BD2VCUPZE3e5o97SQ
iFnC1cvxphnah678B32lBgTc83LxfGQbS4T4SyII/Tnp4yUM+CYcATk51eJcbWY4nO/fwZYGc0wJ
xqHagWn7JtznvpVTGkSe2KwZVdgdKZxIoQIXoX/GwYjhTPwYJ88Fr7pxUhKIFTUhYyo+DtDTsyhT
YdX2Vdl2Zd1eqZXmeRhHCxd5HaBrFNrPnA+A/ya4I40dH2NMooqaQxwhHPrfNGuPoFo9Qvl49oI6
M6gBP/i5tQNt9hjBKtvJ6m6WQnzevTXkbUVC1vMvj7bBmHuo9cy7TVCbLH3cLsYAy03r6YrUpOrf
FQcVp+hmIouApliL+SRLyvTYpIRoUejwD+0qICaYBv4TGHVRc733zEPJryV30Jt5dayKVDWgmIEe
M0Z7YkNZseXhKlgMLJEd28PYRnsZtyWdxvcOddwcq6zIKFZRmPpJpd6v4CjtzOtJzwYedV1LfERk
c+LNEtBCEori87goig6TvwlRMEfj39yV5rLaKIZeynCXC61gcFbP7ALoXPsr/BKJqvOz3i+jYAjU
SfU0WrxXBR9IZPUX5/NzONRCTl9RlHe3TKu1D0fvQ0HcENYlA1hztdFZDqGsgH7TLiWnwRivXHzQ
EIQoRPLG8Mc/lLgitORF1c9fMs7FSTG6cPRd5cgZgDKVMSllenFFS93E2m5CfPYTIs9jx1u6ZTJf
0jMjDsaME4q1n+3a+YaUVyovBq0m1BQequJTlInPQnZgQn0hhzTbx9WarmjCVJMbU5HY02WVNlCv
ukva8Svsp7CQqXaoKXFF8SQ53fnFIhFKGdBCMTM9IEMqQaQB4L7d1NmsLjFPERjut5FDp9Y/uThn
crNeUDQOmALOrpeSfp5VKGzDkBli5UjC8d3nCO6OudrVkAWR22MX0v/CoSovn1jZ+IM3xSgkj5Lo
ZBQpEaNQFmH4n9czQdAUHpAf3OXuBurJd33rRtt4r18TlkjRPZZM9BxfkqTV8k9EcyZPczrH7HyL
ty24ekRmLTk+kohc4GVitbt86Yaya4qUfL3zu25TI/EleOvI+Z9KhYEmvqDGGkOxJ/gdoEGIOib3
ejY7yEhh1ITpyU7QnpuRThpoWGY6l05pjtMPcNzow/axjeQqualljhlEwtdKVrLWRmuUVc3JSZfb
SYT2XKm82sxjMZkl9fWZliZPhNHmWe9gN2FdUWqykXEvmVg40cQvzKk7veZNxPIyJuQ5hL1t3inP
Z+UUvVNzsaLes/RHk2lDupPb9/coiS6ZlcWXPn1KBKeVHsJxfiycDQqem8M/TXJqP1T+HOM6tdZd
z/tbry4H7Vum5jSUcPimhkG+qSvRGnCoHTo94l5o+V0kb3jUuZyaqJILW/CadUEMHP7GSSIPRglf
TEx324fAcf4W9gWQJRxvmWnh/xEPg7jZF9CoBc2nZF6xWDJBMXv/ADeZdCvt5TzkzKLIOCtH1j2a
n2PShvdFeJkRAddANXxgObD1ydSmcae1ZDy4qkDnfHPNgNCX9OkEtspwGn+E2IH3pek/trhzMaKv
5ERhBeSg/lnmFsmshUpG3b97RgmnmKkSwIumYffWZqR/ov8vkUT83xy2WMVb8mA88IhknWAH8Ux7
C7f7NM4X8+sxPSUTtFyEm+3AA8CLAQD59xZjCXHv9zlHuoGWDNyfQF7HFn0urBiLcl19BiRHfe34
8cvVZ2Yca+9vo115aK4xB9u92wWhchJJerHai24F9gyiawTi/8iN6fLfdFEi/jYghzQCmwk96e39
IQ/ynDi9znxQnEJbyCNAZFSYGFdp8BZ8lFdogPeH43sDnzn3SnlmitrMQsdXQZC3W1UUG6vvEW0b
eYg47maIel3No+8Yv3bkD+v8L7UKBwGe/VXrjf/H+x7mFBGzeM9dP0Innub2buD7wgmtlVG5qAN4
/bxzY8AkU+3gyAY4/xhXdd0kFi7qmW6CEJdvFQJCrJ9SeQnFwH0EPEhFq4G+C5epfnawz6WAj8Bg
SP1kjEfEVH5XHKubmnNmyFJtFGwwV67GAgUY9JTWUR8j2vU2veA1vTtOwMT1QN7AQRUwdejGyXAw
J3qp8A/QYLULAJBSwp4CFqicvrnOyPOMkUy9cW1o9Rmx0ze3mZLJGPwieog8xtNGK7WpJoykVuxZ
BDQTLjGn3Brfz3dVkW64I5g5O4aZOnylGuWEg2Ud7nn75NhlZrYGLDG4Ut44G7DToZDFizZ5nI+R
ADMRVFkRUnypM2zl+dq7j46IOslqZlGY0Uds9dwyvqeQcW8rAArLPd/1XPdKIIkutmtT1+gGxwBr
Qh27Jwfi50lh5j3sB9h6jpeKRXqm9bRiRhDi1DgvlSPKDVL9oSbEOuD3MAjk5KgH/PFmvd+eMtsf
qSBZ5h4vTlQrhhVBQAciR9pQMi1KKQpR1VQJiuBKC537PPfSkbX10H8nn9XG4IaoMbEkTo0+eODe
vBa2ZLPN3lhlihcfjvxjyYBHn73UgGczODghhylbAsemWAtSu9wA3yD4YemHddipgx6jKYt+7mDI
oTAAOuk9EWxRYhA/4wSoKohvgfU9zdz5K8hZEoZz8whArt9tgAnQ435JGtYuakdtB0MbtKzaS2QL
+/sitDNgLjWxh5T8c/92xgQ77fosmI7lkfOvojtI4s4jki2u+Aq0lJ5Rvf1ExcLpdntY0T5RtDLn
9xlFq9TKDPeKVPckUwfiN0sbDo9lJPnq2xgeBQ+QYWtTpLnZXz8Damq3rL4gLd0UtSclCY0o0cEy
DidDwjPlha9Hf50vgFDkoAJuhAiq2DVpl0SkMD7eGpJ4A70Wi3iXSij7RrVW503utdIS6cw484yI
J2vSTMKzGwVMj4hKjApRPN1lo/4wijMYUt9dRlXAHujSlm80I85foA2EE/7E2JQZbnsLpvHNscZ+
e54oO9hFje0h1bAY7vzwPvKnpUTJXPHLU1gAfrDAMHIBcpQQJoaQyvDBpO7/zL6IBC6HsREbADwb
dJAHhADyxKZxmbLO8izGqlYzcdtcy9zO3p/tagh3yrVcWom1njtVCza/Y7FkH8B3oN1qqWgHQprk
Q3X+tGpBwHNKgxLjpKes51DY2pW3dKoFqgzEdr5GyDdjcvUpYd9xC/acWGiV4fuwHfTQmR/eLUV1
XLPftTxcOrp6KyjIclgUf3VM2cBZuPAKGEYr0TR2rTrF3aeSc9O1spj3yKZngx3gQUZvUIiCbarg
DtQN4XFaoqITMGA3TFUqLbr3Qi+hOLYGBDaMj/sWdLVdV4pFKZCK72fpJPFcJ8V8oPjXTZguM8/f
RUbjrbTCwFDNXFAfsIEz4wQFC/1YO8dRPN6jZTa+vdTuSaMFCZg7CXAwOXzl5XwF4RYyRqjboalW
OD8kb7KnGanCfX82Na6hq/eKDWR8sMt1AMEhxrOKymquqfYq2O1dquON7p29/Kfe7+Fz3vp+znwF
+MiCtKr+agPJMk/HtGgw703F5KfX2fBQU/u4Y0x1Q1ZXpLpiIfwgXw3fjhqBJbHXRjzVGeof7hsj
XEFiD5IGV2r0/RNkXnaHpgop/5N8+pOJZmew+1F5QJrKj3QQUis9bVCMIM6Njyf0p96gfCvM1TG1
EuPGXLsYlvtyeonN+k2RnNadmM5I2TMtlX2JGh+LfBQHNpfOAJwnO6meCj1QaSaCo32RpvHpC9MX
UZdyyNDRAKjjaSLFfDRsIfWv/EZywj2Zgy6AyH/ctmNG2XXbU8rpwsEMNgGlRepCiCCwyIUjPHHk
gs4wo7p4UAD1QaclDDPqXMC3/yIGRKI4YwUcABYBBurL8u20iC2wEBw5cxs/bkE8+aUd36/61+IJ
Mup6tybEvpNS3Djg6z28wbNQ5c6+vEP3toQKDOT6IpDC2yJBSBU51qcFu2ot8QK+jUhFTYEoC5PG
douQSjqyQ45rCwtkLPdryG3FrrhDiRQxW5wk9+4GVq/30HrL9DyFSX2tMa3WAXw5tXKeL7QtgB3K
z5oVKwccKhnbAche1hAGDz5PxyEWj4er1a0ioZ0xp7FK5Qw2Br7V5uuKeIPtbBrpp/FFaY5N0pKl
5IbgizF8Uug94jhRG1+Jkgc2gsV9nJJDNcL9wxN+CSMvya5k2mmytTFoTl3P5Kid63sRAaRu7/Js
b6I/GCpVNPbupJFQ4OIiOtbH8q8Fcj9oa6XgYnuZgNCJzls7thoMPhZvK7fD8vlK5L8jA6iKiyZQ
Sl4v2NNdE2kfhz7SxPM6avEGfxx3+3n/bfGv/ms+BSMDnZJApAl7A3SHNARpHarwbG67r9SGhmlI
nHqpfbPMGbVtZeZzKqhONj/pAZBERF+2F569v7VZkyH1j7+C8s5aQ7A/cQhYoi/YUMIHz92jPP61
K9JYTiCwv2vuyALrWHvj3HTJwJGUeWeF5KsvRAk5s8j+vA/2LuLmqqo5nmFcVbS8hokA8jsk5l9S
aELoo5Yhxs2HSjrXqCo8ykLqV+kRQbqYRrHV4tOi+wcaFWhaMDbKUSnmx36wHrY5369s7eSONjPn
1MadoTziWF+KNgy2pcnoSZ7wtXwFt8fli4FbMyMv5NbMlOt6q6ckkv7yag9eGmMQ1BTL63zFBFdn
j6GuCFTefDWjn+R1g7/UdmA6oEsCAabIePz7b063B8eLyA1j12eLqAordFiXUo0A3sdBu6ux7WWI
TUYmu8p7Tte9i1lsc9im/J6wSD7tUlIh+aloLAF/lb1EvNrSkjDlA+gT5sEDhQrn6rrexTQsXY24
uTQuOLVTLDHPIVqY5ItBqrye/mZ8Y+0Q5LDYK+xFx+uXsiAmMS7KhBgQpmETgLtXFp5ZKRGSCUFh
XMzAJbpLezyQQfx9602OXeyEweQ3JMtOhnbxYZD6ozoeLHzMbKvdCcFY14SYxaRmdqJ7+z7qpXwo
dj9iVawgCtLzvCQagRPVnY+BFVVHiYMobdtaycEolYgMAMDjmAwYI3cYwjPyA0ePR0ljnZADFpiz
NR0i2Kvur4bAo3goTol6waQQik/3bBV8TzYWmFObuGsGPfkW/Rzgg9jSw9Rfv9ntLgUG7PtGwtDY
25xlclxX5Njdoq8nN9BVRANZHHCd1rPe/0QM5YivYo3Z/V+VLWrGsXxqk+cTL4Ttlks1lIlW5Yxi
FRzcdIx5jEfXt9pDOFlwAGgr/W00paifo22A04s9iA74TOOP4xPmmLDNZEkEY/3UaweRlvtPWByK
uHqUZiSAx+sbU/gX3AsOnpqgNKVe2pSIixNQ74Nsz6pqae5u7RuvtqJWMSzxdHPdwG53ZaodJlCN
tT9zQgJdcniTb/BOwoZrUue5+xRHGADjYHxz0f4PKHx0jc2cxEYevyEhiGibtwzX30leRn2j9dlm
ad13N1mcfzXMCdWYl1eYuJM03oWtvzBYfGXEYKvQwLHOB9f5Or7bGNdZMw6L/zC6nmwKtWH7k5z2
MyvxlmIJZD82+IdEHaHX6/D43tWxoEr+P6kxi9FL8NeUvPhmbHBs8wa4lYOqLBmUyQrbNqjTLzG9
d4gl1oUUPDpaz87kQgW1zrBpJKU1ReRt0vxb0H8mq/35rn5Ez27gu18+zCrnz0OnaAodDBZ+YZth
LhVGjA/8NKmKbN4oQVOcK6SE1zcDoDkAsuDeBc+a6s3REZCdESi8NUmHlccEzzjZ/B5H2aPPTJ81
2v46I0v7LMhBD6Kzy8XQjLmRf8Y6hjIRfCRQT5yjniLWUFsPQt5J7iSFOYhKHzprMY2KC3M32MiM
WbJyFgQ10vmBcAwYc1qX5kV5SSXGrBAKMhOmK23ZPHJ4gFOnZFnEtPYNMLAjfj3o0QXG6n6TAfEk
HI6WGKcS5ZgxngLUNPQDtOFPN0HhRkKv2PXftp8QxLx8kT3KJ66CqgdvnCUt9qAuXg39aS+VRdu/
ROYXsoa0ZB+SQQNljXePWmg/ZO97L/xDskECgtWkB4NolSkfABOOTANcZJcqSVO0iyd8sy19LKHc
IJKLUdB+3VvmBB9D1O6i1/kGHzVCN4DlwyMO0sm3KEscr9f47WQBI241zidZo+CaKH4Ww2tZQwSA
htSTHrZZ14IV9qYgVgeUa0h1hZe/8zUPPsYAXxsIsob8O3tW+qjmMF9NjVtAcmwTcmE/ejWl+Mxz
w0pWftu2xKjyMQg4wJ+Q+QnSeEn3p1X2GWOffxe4VDpbgCrihBB3RyEcsQ80cEhzdz3uT1Vfc3aq
by2XNxCXh1oEkIKcyIkJQhl4KuWVGiMC9Tg49c3n9R/uv1LL9NUpwSlhw4DSo3M8XiA9itSyxmo9
ksnsJ90V74xWjHBxPAQtGNeXZ+VOHXny+l/Y5E6jpJGo76u0/a3pVc4Ge/YN8Un7YD3TUdV6Mope
7U4GWF/0j3CaUfffSoifbXhWBQSoLnNgl6fgqtHI+wrX9z4aLBBZUft0Mq2KpHQgzW7WbKusMlpm
qx7VtTvm+HUOc304bBm2avV2QvgfXkKPBwZcl1y00N6kiflz7W6Hy4o/Dh3pzoC+vsXUTFOcXb8m
RdWqEqT5DXFMwzqdPBTgvtAVwMjcH1ig0WORi23eiELodqPGTsfDVZQHKjSHijCAnolDXPgP2UND
qdT94nDyQ26D3QdwWulewEh8Q16Ysm4lrYIJXKK3cP4isOJoixcdmt1n9RgtdnPb7iMujJkwHSSQ
xQKC/rWXJT6Dha34H9kt5iYJekB0/wdL8T8i+dha5qIJpRXu87G/GpwSv85SJXKJYweAokA+d6jW
ZBywOSman4eGDJWoLh6+a1w299eTWbQw8vLa0B5tN3/bUQOom5/2ajMykBfKF14AqR3LC0wJ6IWu
ziZ+ck/URHt4ovrdZt6VXNgZ61O+PaejT+Cla1F31TsCj8NGCohI8hYNBwtzsnv5LI9DSOs/zqPW
/Kon7RT7/hnkQrndUgvP7S5fpjqylT0qDeTzTwHyPCXCLU1D1p2b0VPGtUJvVaXc4EDyQZt4ncS0
HOjqaLQA65ZpN8RiMWMQiVh/I7rDLHkupCURaHOP6aTh3ET+TW9IBkDxkQxtvj0VoYzA/JfwxBv1
UfkxCfO8x+E2rJ2BAxjrnh8k4BC9sW19QtUPU4sAx9ZPxcMd8ETjejhXHMl+iDhl+mAUCrGpdHxL
updPIjlyXYtfUVsnfHfo2I6pbT22CjTVTgX+00NsKJtEGMocKo6wNEykXdGHBKpcrRFcxCiv8G0d
vdFlSSmFTUcfUb0K1jU3ToHwA+h2+rEx0c46yCWZvpQnkdCAWYOaPIJetBJVkk3gCr+YAfv1AKip
TG+c04E3id+c1FDL1OBhDB2RaOzE4GBKoA8opFTLzVlUIzaB85H8WZwu6dVY/IFtffB7TpH5Aw8e
R1YBRAAwqtBab94x90yCpZNwun1SbKebvXe+ZPTMG0iwXuGFYhwxI5hyeoDs4YtTZzhxhCL+7bqx
f0zjA7u7Nve9Kv75dywnCjk5NQvae04cpBuXqiwZg6ya1gh8osozX0Xz/0ApJZSZbGKRwpBmG3Ob
np1796Ivq+P4YGeAMNh8ATsaaVU4q8X184iXMRNj0YVnHQwLxm4IBxeW6AyrLQJeCcJ2WTpUfmyu
vGQIBjTOy8a8Dbhdkskljp/uYnx4/V4IepROrj88FXnl0Dwv1RmGFefZlWUEWJdP0/7pMMNm48Ed
ORiIHWLcVbwTiTXqEs0XN7581Obl6aohzJBtAuZEPGEzQ8Qm+w9X05wg7kQ2aRPF8r/tdyq+XSHZ
HpD3aA4Zz6VQ4HxBCS2vQShz3LXp+vHn3u1xiadZ2kxWFBHtq57MRlEIASkO7ZlHp+GgwXih/0fy
N/3WbYwYZG9lG9J2EM+2PcAQllbuJ4HCZk4114hQ6PmV8QcEMigHn+yhs5FGIZ84EgHEtzuaYBjm
M/6B9APFsHMnoXyhdQPHRsdR8PFOzql5UBe8o1n9wuvD7ZnmhMZiESMynho8NClReOYcV20HThru
SHH+1EnxkPR63JAb9ARfDANPvIPDEOx3lPtj4s6f049NXpLXLfbgfJlBjF0u3jtHkb/f/nJtgjE1
BqNN1ijnSDuvERSd7oPc5HECihvH94bT0uTmJvIIfo27c6MPUkaVHkOfc9OZhl9F76IkZkaVzCPq
8zMRva5WZIVxqZdWl/lxhmiDPQ7Qelrlz5lWviGesWMWj0armgVHrNQ7apyDPwsjhkWCxWPBy014
qotIv7u+GoLaH5IliDkgZ21Q3e3BAGQw+RiBrNc9Z/hq/47Tc7JO5LaN2PmQG7W2aqmBDKIHseeq
eaV00YRguHe8VnRR5l6FIXHXWj3646rthjLyCkpinClsVF2MKTkQ02jQUEzinjpqQFozo7IHvs5c
LozbD9NF1l2sgh0fSJvV2yULJm16JJnA0eTPnLA/6vqBwAOFEUe9E/Gk8plSBf7baNoeN73/kkFN
TDetN+hh8RhpxKSh+mq9dS1HN07MV1JvYu8yO41FALvYlUxHOuAxRO/tUrt7xqsFObq41Hv2sMpA
ZVZyR/WgMHLfLJ7ibANzrbITReLLfcESaZ+9B/dtocI/rtJZNcudx2/b23r1BbR2EZgd1Kzi145N
GufGDBnOHYvucwdg9S2LoSUdFRADFsA/590c6CJ8wdg8sXNz4v47O12V/TYH1/MTDjP0x1AlZkY5
N/XqwygxSE8axOdLEwohwncdeDXZNbnIvt3M+RsSfL2YpzMCyei349YHRYDSIQ07gMH4BVKFlSfY
dNVYlOzICoYmSnq0UTIbg7RK3ZdA4lG8FNUt0PT33p5tG3vjAaNwKb6bVbHiV8I70P6Ff6B2I8C6
JBeO2P7ev8pZWc4sa6iUKinbymtyAXKhYTN6KTLqktazs41i9cWbqbfAXtzt4U/kA7mIkeiKFf0F
4gNL7kxDYOzZUvFQ9pGE8WfgaZ/7InwkcVyxIZfSt/lAu6qj1UtDclOgn6ioNW0YCGRo9CF/PK7J
GK0ij3a8GMT4VCObLZZWrI9t4Hm/RGcRcHqvBZRw/tRav+4Hdvj/SI+b9GPZQAkdj8BDGSPxv+A0
uBksWviAVVpm+9MAK86PxC8V2faX3swsZLZ6EDJxkPus6kWELuN39fARUoqZySXmwwzTzks4koYR
SlZOL++RL3ii8T48yAvkzVi1fRia2R+/PqbqkwBEa2h9x/1YEDtNkiHjhIVmdu3Rp8QJATvTfhCG
2rfe4571GVnd1nMetXy5wAaw9wSl5Ae23cExzOQW8osmoUFUIt8+uaiUU7Qb93Gmj6fOnYr4VLsU
08fMkFKK122loeYgrF04fh0SAZMtiloUOnrXZoHwZiStPAU8rI8IZCzOaZJ/jULEET3SgLK4GI6p
ATjVwiBhVd2rFEnVH+wx4pnKYCraC+vtjW/4e6iO6SYG5fT9U0O2J2nZA0nc+dD43CJHV+Ac6gsj
Mq9MIHRCW1b3NY9au00VmWyc1AIJMxLUh0HsCz1rzRBigvQmAHIJRbT5akprjE8/hpAfPmwFwuKt
FmWn9DSCxlZYKc05Pcl7gUAVGNeGZuk48dfvYWryPG8ixc49KxLv9gTEimtTx9xMC398dMMdjvQ+
A8Ys7TAfoaJzdRMJmArX98CqmPu27bduwfcINPzeaIULvPzaQJoEPAkwnGy46L1ja+ZtO6+0qE4n
kFZG9e7ttR8HIMn9GXt2lOvP/4Wq/dg5MrEbt7NfXoSpuTSq3zKv3OQ0wDJkSVuVBRV2aE1R3fum
yahep5WcuJdqjjIduJoQDTce72oyaRqotyyxD7pEp+6JTY64PCEZJt7s0oZwYM0XKKp25/noRtNT
+1qZ4FGwoMiEKe0tFYD7cKnN8zREfSDZKc6ucnwzv9utCc2ewgeYOM5WdMbv5+WGuWOOtlRlRWij
/uCZMtF2vWo58eXcei9C5ju7xhuBTW9qIjNjmW/qBE6T0TVvQw9+rzxfUMz3w/BTUmdqNWpuhPDZ
YS6Y8VYSvXI3yMZm3gvapuarU2hhYYOr1WCZJ3dS3F97GXuufI6O5V8gQJ+EmDjDk0jysVHssSDC
8yNeqhzNwWeYBjd5bp4nDJT+CAGLRtNlxy3bho5jSa3IYa9zt6Wf7ljq3Xc2U/MULSNvicAndor2
Rl+gd3iHbo7UbNqYSBuGL+rQGxWJkf+19Fv+A2nH+PF1peM3Nqz/pcKFTRFlWOO7WEUjs1JLjcyH
x8Ir/f09egv+aMXnka0UBr50g8scTdPG0wKaMBgr+FaOv3ro3GbjTtSs5sbpNuiHyCt7GNRDabcX
rVl/ikH1hh7yGVLdBfWG+5sdmr1hBBmjEbWrBZE8qyV1mKm2KliDh4nLl6gAe8VPORI1zyfpUdrR
3vzTCCw+m6zw3kwFgbkzgdbyMJCiG83BPBXcR3ssiAPdlhkKQKYZ6oEl6HTd2phgJlNUv+tA3IfA
gCUkKaVGw/HcQx5LjJ8uxIwAvmRlThD2PQLCNZ9moJkGa0CKE6HhY8MENkrs5BOxa7SREXwt5aCY
jWz+wIVw3MPQiSbmgguo9XndzMt8INQugG7ODl5G/F8OUBdwvpGcudLMKLIz3v2xBDTDUN/26Hnh
tGHBJ6CaG96cEU5q6bE4i6HyqpXyDpPQZVRWjvf53G/Y3bhCbm5XBgyLusyxzRW/ZhRW84QXFGUE
H8kGTpfaKUCX5k5Maw3dhSroE/jiMBeU0YYFuLKfo9HDLrdU5Uq71SFc7Y/ti3HHarFxUYxIFgH9
j8xL16R4ociK7SHG9sKdHPowH8YBtSIObI+Httc1gpyJJI4dsCWskvUotUUazaRh0kZuCSgF0L2x
7k9l3473XHaNq3LFIr9khp3gq8VsOBtk7LNfsH6WIjVwNiBnA0NDhrKdApVyvlAqjKKnd58wsi1K
QgP5ZmQpaAqEqu+8QQ25DQA6LVUmzgSg86HJe9eVsE7iErodic9abphfjMdqjwB+9lwhyw69HZkm
/6uMPQdQE7MmokQZ9ezLyeTGYdPRdzF7YmI9oQvXNJ+TnXCs5Wc9C2h4ruoetNuyRHECc/wZijGw
xQOj2oK27oViFoKkF/0qiRr626orpxAZO1Fc0SoglO/In1MGnubVDPIJ+a7Zz0JbAA5uVP4qOI7O
b+trde/wisXzpKxIz/h8/LpD0Sxp6gLCWrVhSTQQOkSVCxVdXQQLt4G+ATHbn1/VJvQJ28Cq9loH
yxGNPtZty/+vtU2MTx46KEw6h+6XlDya5XG9iorGxT5eUvtnFVGcZCAbfgvLvIvWQXiLHs9s6Gwf
YZzp1ao0HmgFJyLuARW708CRkOOldbrsIbPzW/kRM7UxZAtGNsZFfOMRlP+xYpGtJizaqZwctJTN
2OncN4r2/bJPYR/MXUxSsOYzCkU6iGx4F5fbQR4ptujOlWv6AgZpeLKNSQ+IqEYrr2sJvpZd13Th
BuSVPvTna1auwJk9u2nwr74IXDSVgcFCJqA0pPp4vmrtItka0Cl1OBYqQ0EXUCOJniA1FQ8VCTDF
e305VliCImQdo1yTJZsm/xYx0cwvhtJMikUph02b1LTLmOgp58JLoEfDd+/JnFsVst3ZuD8O7av3
5VQRzLe3Xj6eVoBqoMaER/GFP+gLsukLCOYl38ScX6CrJBE1pySB73f0CPreNgrSk2T2RrCEyG7v
Qf3np/kIz5xmk8oIY6Wz3Vd47Jbia/ba8P+uaZHkiwNoCC89O7gGSVsrTrRj8fV+/BqtYpf8duT/
TjqTKqm7ZE82tks4am5FwdCArcTIKb+t4DdGdqa36PF8kJeNjX4iPtzfylrDM98JZrq1IkKD+mlS
0KbymY4jvIeiaY4V93rpTvDzQXEOCv2B6jcZAfXM6lptitSuv6YLYkADK2xLac4GvRKhH5HVR4R9
vC52FL++ZT/HiPjbXULJsYW2LvA5dt3UK/Ww3FPILMU+hhMbjZDHt053zzUN/gOrbZq4tPj51OnD
6NgUTtk1mjg5kEE2SgNW1WPfIKc7trx86yKtflWfdYQ+IMy6nch+NjD1N4bbE2zB8grRhqMoU+Li
8AyJyaauu50Yk21Ib9ZR6nblfJN5RKi0SGP1u+uC6hdzF34b+qQbq/nflMRA+haKIBefsV80k2ml
aA9Qp4pjtvjD40acj7DThuFwmyLpPddWe2q3npwxxrODdhZy6mEzxBz9/qwKk0gVeYuvW2F+EtEL
b9/quMlINw4EWkdqLn1+4FpY/Tzfa3hwYUA1cAYfpnuIG/BapFrGryLP94nVJDAXQ0R1sBJlfPh6
0qP814KxkckXM7VkBlKgHp+4Yvp0t8yVdi9ae36nI1LCU+saEfCoXwBB86SjlDl+HRQLUe49ODPy
OnnkVI/Unm+9pne5idQLPAz7eHFC0V/4LhXoJOEmVgso1+1J09dt15W/zgpeBzAzc7NZ7iLARFDn
/POoDvC6ySiuA4QLEBqodgjXEEi7VHKjGcFqfFQDMA0tcSRfVYcGzmNJ8fziHgfL9HsehvrJszqP
s3cnfrLhuy6mX81I9nS0/vZEMeF+0bqOVU2JKhf6kYfhemO51gMN47cLLLBqPGOXKfb0neFwNxv1
O/3FkXIljqUaD/M/bLL9ksCZ5rvZv4YH/RaCSINxntPgJ0aKo80mCao7UI8+LCu7fpTaaSb8hiSK
iSyAbmts029W7arHcn1vwbXgP2EWLkDUzTnbcIGCmtN6NixHNtkEsM4M/PL9cO3GHfpchOQ2AaKJ
Zq5XTqEzvBMOUkbPAfQgtl43OcvBKAlMC8J7hQW3R9i6X477a2wyspvKewqG/NEgMU8+pWM+INdr
eROxsJDYj4UkHLbZvwtYqPORhPbCoCs6wOLOCcjfxmenDGrrLN5RmagcOm709+YzcbQViUAu0Fl8
VwLrxsaoqV6iz3yI3pX3zEpyMWSwecWW8ghv2tXYl8eWTzUTQFtBaLA6FAZq1zlH7DB6AyYWQ/o5
iv63NuRxneOdoNfBxXKhWHwC1jZ54ltJC3sjZoERNA2kn5DafP/f5YUYpSPoFuSrdxcayP1OdIJl
wlhcU2mm/HO+N+i6i5IPN9YSIQrqthdb4YbJ2oHN+hck+dOXyBrEwICXGaGB6NWVn8DlKZWHdy0J
WqSlKZOXFOgyiO6Ra890b9u46HETRFPQuPlbYDlY2qvrpK2BDYFNjA2VbN6JfRKnZjiYozhXa6uX
8CCd8QEy+CYGPBR1eMPw3mqL1BolZb+jFG3xYSeF4UtCsndd/B9sELZCOPE6BA/mdp+E3Y9BdGYR
copjyt3NihpRqHnn3U5AOWigHWpsEoBiEBeOFpAVg842W50DuZSxlKQtOv/Nc8nzL/cev29aTkdY
ZlJsUcuJvP7jYRrt4KIAzEpTUo4wLgDjb/H+Rr5uw/wiowoU8o8WyaJnsY2gzkBM7ikQcrQoWGCZ
HQzUoSF5YRvGaUJFvBeB8R9USikgOsBGmV29PlX9vdhc1WZy+A+BKxvoJF22AC7Vh6Yg52vntJnl
Qm65eka+c5vJGaTxydFE0M9mgV9ND9EDV1U7XPwWinyWpGRvdhjwGwn6G83IsFLBIPXH0wcrxkqm
Rti03pIoKp8QO6z5DWcnQOcrtTEZDsCHeyU6athhhNBOGo+HhFNP04wdy7zSGa3aISlI3lrFkT+0
Nno6miLRUNWM+I7ebxLNmcvjizpXe3ysPX1ahXhLUU7qBXXU7ilTiaAVD+HRbfxe/jaDerZJZpEp
uzPiJ6DiJwnoPkDlOrB1U/H1oTDXZ/n56jJ5wDQkBx1v7XbtT9cWh3IU0PuvI9yB41UEMQ/vdpD+
kDkq5CCdfhJn5SNBiYN9gJhww3IpYmFu3aiV0wKkqCDqTn+DHObugxbOCIHW/9HFIFgDUqsbpdnd
8C/daxQ+oBPX1eI5KLXPjaO7ZAAHAKq++d1ICCYQNjApyBya9Xk2jJdAIdk3aiPvQ914VuGMOhWF
GDCQ5kZhvy1C19b5BYmrTC20VUok5cQi6sUlTffoXAUgJrVE8O+IIyuPKHoeOQzFuYwjizb29UYR
hsjTaBlrnPL+CMP2O8jZlIPeyVxJq/WFeZmDXJLcq3ozCe4U+gxSRvpdqQmkyKE/LsePcmCcWEci
ZcICCeHoliBSf34w6S1HdFMZthvHAJSG+72yRYm/anUJgJjFr1IqPNux9VCwwlAVenVpJyzm1nP1
XZ45G/G0VeyaIgSyYxrqaOQYylXfqzf9PbwZhTpqkJCWsNa4tXu+U/dkQAPQv2CJY586m6+ieaUj
afHqKXz9cri38KwIaH4DoH+afjMej5v36XdCVb+7DpJGSeNvdqM/aSInUoJgsYgbsz2Mn8m0z514
GYyLRovySj9P1AjKI0AXFCfl2Lxw5JvoddPdrvSx/FDr17UEKHudUigYEYgk1eh4CeHj9LzUKYYN
mcjSU5rJTpp/spgOwgkmkt+WosbPs5R8lJO86eH4RSNlKwwXt0b3bA6rB2Tty074lWtldy40/An8
YRmIbv230ZMkKZe4iUogRQF6PmZmYxKB2UXBvMEMQ2A7Fh5tcLlnDdG5kse9niM+7cMTqHM0Qg8H
MsqP8Or9ZEdmDLaZk/G1kc6rwHPdLtftcbIUiyqGmRNib0SvuDCQKsRm1uTXohUkwX3rfXz6HMLG
fAeUkx58wA7hxMrGj5XLjS0BOhyHiG0ppGYy+d1g+9IY5Za3x20mOqaP7RRZJ+qsaMPX32gSqly4
M79x1gAkFRkyrQZrV6cU+YjYBcPbEFxwGALjeNIYveSBY2eVpoWB+KURiC8vN46HHPpv28smNSh7
pI7hDWc0sTxlTzIJyea5nJiM5AYcJvnaFjnHgzIXzc34120K5hSvWZ7z9RCqywL6HYqtOxjSLGXx
MAmAxE6AiKLVjDw1jsEiDbN3ulE3lOOndUGCIFMPTzX92gaU84qCskPBK/+vZR1I4R5swHgbOlAc
zIgj4caAnrv1rp7Q/f1d3mMpSf7EzQBOd63bJA2fVlIJAzz/jY65boPZfjk4dDH7S6S0lMSP1Ftc
NigGiT66MYoZgFR8528PzjIhDN1dj2pJCYTdhLQKGyOZYLCZjpZjGtzkTFCMOJn7VT/6SZHHAI40
XXqkQ2Fig0QkWAZ2JY01g4oYe+LOmrT85aVp6ZRW1WrEamTW2NfpB7dAtdHOPkxGg6QOaxSLEuqi
8YaI+5R1UpnD/NrorPEH0KaoErejv0OS6l5r84mrZj1KApWcM+vYydnZsxRrpQlFK0MlCZCJKoM6
+Kzzo99lNnUwU0NznilBXdB2I4I/Bs1OgqilNftNqUNFeSExfYiKy8/NbqZXEzg7+OgRpNN47f5E
G0cV6+HVwljcBrjvoAfcMt0F467j9HYAEVuKv6f2Os2AzSvYmfxPacEPec4i54YJ+7Ujci941FT3
FB8JWhMQpokRKBTFlcAqJLqxLKApj3ad0Tgdwt8RlmtCQQCb6nStt710xYcoovAOvpyOJ/DW42KO
VyN5FUnyyuZ7QFDiNkfh2Z0WlV0JeS9cX4iWzFh+llPdadYj10+KTibPg0/02ZiO9Ph8He1aQHOm
MA14Kf5qBzCQKPrpHz5gBfeG+iPeaan5OYB28KFKlrZdf7IXKnzvC63N1iUOHU5VdKuhtui2Ylbb
lW6r1g7mTPH8u9B/1eiKu8iukuUEOPjYvLIewmPvv7lEK6acKlZ8MeO9R2wou2fF5sCLq7COXYZo
u/X73RNPE7HXDUE+ne2aJz1p6F/CdB4bxLfToiAQ1i+xqN61h10tx4q4ND1ZY5Ox95657qZc45Ij
pLWbnUqFONnNHZ0Lx+xJbkUZxeI7ng2HZVISBuUJ4gHLyXT1JAas0kPqp88AORpvQ5n09nHSrRWP
KvyGjWZl7A9SFs+bL1lj1mGotdKMWKPi2mH68bHrw6uKKAHwYtq09kuYq6Ch3b8mz+MN9AsQdyAQ
I27ttKdYXOWte9J33ylakC6N71/VlEAQ3IloNk09x9eo2HQ4R6/x9lwDA1TWEfoolXwlAjAQ6jOV
Tujd9B22CkK5+G9IMc9OYxwZOcqB+hZ35KgEATZU5LoOb2V/Xcmydvsxn46koYQ2s072b454Ix6J
KUGPA/k3fuIExgCZUGfQ0k0jKS/kcLmJAMMZDYg+ZzUDaYYq75KJSsttF8DIW4eM+CL46rB+D2mP
GYbVQp2oSZTlMZnQIoNMUTCbK/bFxkcN00J0Rs/gSYhjklZOzlyPDodTELE212ezThiBX7OiodK/
gmFfvyjlVwtE6lwC5AzuOIxBS6x9+OlV83LMOLOhCkDvmPgC+waNcuz+M6Cuc3gIb8Ex+yitfx3f
FqBI4kTe5xcsqrM1mByXr/9Ev2HnaEED+SaNnyyN7IgRDRbudcvl9galJKl2D6hj2LXSHu+FtOG2
XThLHTUo1110CdY/oERbPLpnKCPemCHvdlBjvjNoFeN4A0YRJhYzVH2Zi4lxO90rbX5pzlkCkSE5
R9V5KIQHZ45e7wkd25d3e1xFkowWDB37JIbuYiAgaLaUUpeNrJ/2pNT46Un3qWS20PB/pmHubH23
8nAM4Tpxpv1OqTS7kfkM90vK8HTr5PZZy/IOtSUaErNf4nZ+MvyPzyCqrKixdAQmEaD8QM7jAYUG
JW1nnGLYnK0IKecrj61qjgPscdLzP6ZvjecWKRp21iGvCBnGAhmQXKe27drvyPRPSldERtJd91lV
FtahN+ME4VIH7R7I+avVc/W3unYUP60ChLyEZqGRh3u1qU21d6RGtZcQWf50ti7z0SxhTi1MOnOe
zx8EMLKbIe98RM30jxb5d7iqiZTK6Q8qMz65FFhkUrNZlGskotiy2Rpi0Vyx1QunXK/Qp9Gi5Y7O
hvuUMPwiXeVoT1U/HjIpkDNEVmC7lP1iByPTB/X5S4KeocSlWIxcuiCmGNIyx/A/SrZeXJ9WqTmV
ZBLULndDzPPCaqAKf23xND1t87mb8IGJO8GLIHtpyeT5KWJoApGvR2Jc1r4OPUIclz2kghVb0+xb
apcZ94OPdQcMg1G0ExqHlg612Wzk5p1mupMylHJvCaRqCMRHs49hehHiv3oRUukiqygsv9bP/hEk
6E4Vq4IUH55ia5pRw62eqFKso+2GLajvPu4tziMOJDDtu0da5CEj4pX1YRfHAtrxWnO+u60g44O3
FJHmvK3+GZZLQA+1Ng2F07tzjWKpZGE4zF72rgxe9lcmPM+LBuhdqTjcMHaUG+UHM9pJHSjCKXJW
Lsvac3alMC8Xg/rAe1xXz10QbqMQapYje0CGad+xU4ieDh4F53qqseMJby/tUNMs6Q2MBEO0UyT1
flwvpPDZKMbSmNuA7pnCPTkljq5eOlvdmngUnCzm70Zh0SEHi9+fXyTyhuq3eUXezhV71vIs6Zr9
j72eYIfcZkJYT9/Z4bn/RRDS+XsTkSV/NDivpoDcSHfsiiSurUhlnqZthU+FbLC6ijXTZk/PpM0Z
cn8HJKgbWaBDZtvypch8KJ5qBew4gsTXjjYQquj6Hcnxxi7I6abuXutfCvs4EQEhK+1D1yaLUPCr
JDa8xdD3PXSuxbQNh2AEixfPotxh4oAnqgw4AGxt787cC1rbeo9lQeZevJIPJXM2HLP74e7a9/l6
pOWjK5r1MG3A4KGg0MWhRrOap4L790LlsnbE+ZCVVhxN525dORmqlJYM4AEK4FWC0cLfQljOJWvs
PyuIIb5nNcypYuO7/C/KH6rlQhims8/9kx3TycBUFJdNFt7gIema0jUHpB54AVFVG7M6WmFOL+6l
chnPFX3/gtoJVZAaP/eO5GgIDHA0WUpLA7QJIjujAgCKKkK3u02BaSNUf2tzToALxLFCCpuNTRPE
C9uxl2UQ3m5EXjDqxl305MYLUxcVRDvxKZDqG9XG8buLzHBivyauKsB93H6q8jqgzWxiEof/umpX
uujuR0Ntk/taC90TrBowwE0lVIgGN9ckfRZ+hdRRVdP8BX08bCRW9mDsYoiYBSADxzijiYkBROSP
NMbRYvzCWgGuFmSd2tgLO2rqjWgLrnHCYsEeTMzlCSFnQriU4g/8owiMywT5uccqj1BsFnNz9TfM
zKKnAyrwYtFKlCp0H73TAyA8ujuZGeSQ4tT1iCSeiH2e/W8aSvIc+sNBXMbq/2FG3qELc95oE0fA
0DLsykSSBVCvFKrOgl7P2bnjwEDLMFtIR8J/OxSm46UXolybFsHPIREUpkarj0Gkg/2ZydJFac+H
M0X0FKagyxIYCrmLl6Im8fXyDDmNaeYNNfA8A8gOGpe4zaQYovRS5fx3BFTTQTceMC2Taye6P8jp
Hu92lcmQtTH88KhX5MEB8xFOdfayDF3GqGSpLjjURDbsbQ9Go+/PYP36IPD02FsrjEgtlxMVuSVT
f7p22nr4ADqOFQuIPonjPUdpnqMXciJEJhaEHeGyJzij8Qjdgh0xYSrPuK0RiZkg0x3XsumTYdGX
4HgimdXO89dE13rWVuynlr8C9b7Dto/3VNDnuy7yr0Q72zQc29ZDcVcOn5jq4y9KSdsS6v+HU490
8B5nQTp4fctA0pejDi7mKnmCIww4K83pKLZPbZSkTCpwFffJ5iBWDkT7dnuJl+4Ls1olenTDVAMu
NPPzDmqi2Sfv/25AlZffKafaRNqkGZ8EnngE0hzSaiZN6no6C6HwqSFVSf8bZn6f1Ovb+Sox35IK
uM+yH/h1Tt36CtT+JEhVYNxWhvjqs4xROLwx1cd93fezGcj72UzS7RJXu9f2SyDPOeIpkABDS6pk
sNcFQPmahA6FHs/v/I8H+ecPxM8q+WisrMm51S/ziuYYaQwFKZyRO40DjHg1lbRob3NzF3j4klWB
2XNlT/7kI8F6SXnac71xgRPXaJceDLeiM0nCMI6vRnKclDgf/iHYv2JOlUavg+Z+59fin9D3upJV
UsDxFnZmWc/4YZ70WvwRYknBAdQ4H5jZ3u6TZt5YMKrjmr+V9CI9K1jDRDGZ74NxeM3LkbzxUZJK
trOU6KlXX1iL2RpnrVq88zZknHOzxIYTDtUOqOEscR2OXfB4/07YYF3uB3OvogQzBrZQJtS4MTpC
LT8Yzz5zMN5xCqJwYd7meXd1mznXHbvIa5EpV5Bmvxo9u8yaa5m4cJYNps64RQObY6dlilxtUVci
bF59dBvEgRd0ZjVk0FX0XaxpJNKfqCOQPKkjq+K/TZnnWQlmDTw8Foi96zm5NoDr5vOopbrqmYGj
08vQIVzK7fw//b5eHeTuBPygwDDspr9c7g340lEJDTEpV8LcJFUzbI+IiJL1Yw1snDgSe0cyYH1y
wrAHOgporTVZ1wxlFpSB5/0RbBtWFiq6IS3lfatdHMNyBZFJ9p+TQCyuiQ20uttdvHHcESHNv66M
P/9Fv+V1F9j9n4tTqa5As2SDy8H6TKM7VRVjlIyGUBcIr2MKqs8VLZUoVll5OVtcT4kkh72FhNYD
uiifvZgf+FNMHnY/5KarBOSC2cUiWkSHIIk8euqKhrMkHODMhI+gFcGOD13lzFEa8Yn6bY2m/CW3
5Y9grZXDPlhPJzBbNrVJag4uPAkV4EYcd7ObH2YgQ1c8YLnPZXLe8t+cT+WeM38BGAsByLju/Cxu
kcHUYFcZ/Gwe6MhfmaXfyFKiF7FW8V3sZ8l0QHKZWM9CGCpvOkftlu4b8h4qEkN9YpWiFZKUu1qr
IdB4YF0sDTaAJJi6Tcqos3Ov4piB3UJxWfSlVQcMsfpI9CmJDTnZddxmQncJayS9bzBUIR5zTq5b
2nUfsr2T9WeYBQj5ShjoL4vCKm57pMPrf6GaQ8iD50bt73EhwB4i6RsgTw3p7ETw7+o2l/vn4E+X
jNoViQ4SbVWOB5HUbLob+lr1BOjWopjKUHEwAbrVRM+A+dwd8U+jUXAKb4+2a2ckG5RCiGh/su3Y
P5ftL6NOEMaASai07VLx3Z5RXOkGOW5k89Mpp2LomINrIr5pO5iRp19eM9OdQyzUSttdXHBMYjjP
nMZIyj4GpuZd6VHmMBXd+ba48Aika60OjGAObJurgt8xphE/dC876fRvCMRRwvEidV4HhWjMEnzC
Pu+kVqmx+/zH3ihsMkGHhjU0/EQ967c6h0ydqSTc9vztk95xNuiYTpn6FPipSzj4hRJlIYxIf2iF
4iL7wYSS53Ivn4GC/D48sfpaH86UlWrmDEKo84KEaIZu8DYSRs/5Efhb6Kw1Ctv2srAoxTbVALR6
10e7rx0BlKXCyMhFqG4P328c6rM9/ijxLNCs6xFbYBXrOJA0H3jBoGHcX1lFLjgDVLsKrcFL+d8C
PncZfhTbs0OwM+hlFgM5sxebv+jWla/uMndHhsXZngEMMPYXnflfbpYiWRMMvvPP8ukMb57K7WGt
TIT9I8CdKyOlp+bbSV3dLneU6rHRhO6X/Cx6TBxUslKyDzjF5oj4ByhOraXaMhlD7LPbg3DMInFf
WAku1vNA7sg+0Yk/FiSdQrZ7cL8O9Z9MVJXOTc/J3XEHFAnUWypffez6GkT6116FAXyEYvHBLwUZ
URQoB+fqOpzNIIClZEGDHuWe8URuH+Mw0sPm50YsQN0U82OWdpA2ScsglVKYyjkpNNt12Z7m8CXY
DO49I137LxLpVb9fnrPWDC0aRPQ4/tHxsVZGOqIQQ6b9H28Pw1ToleFs2EtFFQtVpMIX/5d56Dtf
O+ZhrcBvoDuU4SaiQgYA6yUcE5Ij1/cQLEIAu4/W5d91q4u0UafkxjT70/YhRMHKsmn4JTO47VMo
hRWlVslIT3etbWJZD4cvJlr5tAmy6bAi3Bn448b8aRSrlqMkvQH4VfI6yRojj7fZ9CVIpvia2rIJ
NPzTeUHxG5djdJ0SiiBStdEID0599+G2lyIDClpMQINpOHiWA0NY45g1QRRKeKDxPIuOb4OZjV3e
phYQrj3TCJnWCjF7g6r/Zc8JNm1aAM1EqaPv3QcS+zxydiQNhG7d0fh62thYgne/m7xrEPBitdlt
LJqG/xi3ILMzvLPSMG+MJXv/r0OOUEDXZqqTT7eum7kR0bh2aV1aGQDWe+khL4U3pddel08Xt4yw
rlXO/aiRsa1inZ4vqbfPzME/zrEePDmXXi2CdQ69VQtpwj5fByijn1FlMToU40k2rfK7aS9jRGpq
6HtG+v9q9GUf+v25DGnd8wXEtniUc2y46AIyTjRk4YT9i58zOlBF6kMdU3ERrtPVUSpjLQe/8KvO
iGJjtEHsDj6r0z3Z0pdFLUz9RqYykKGdd85xfuzlrZCc3xZckQn7vFANBJzFiEHS6SzhFuupw47Y
jKQnvaJa/y3wtl7mhuQY0n+b+K/MX1p+XzMstdgN4zAofmyKDKyCPQNv4siuU7P+2spoVcT1gcrY
4TB5IEo30JXkROroxMWvWLCMOdzM6PDOYk4ufZm9eo976aXCr+F/J7nDqPCNNEb4q4jfpqWoTZSf
70UWPx2QcGOQiW4gKT/mD/3B5ciZo7FkPNhXXngfFxiGlK5qyX3We+pEemz3FPvUhPkRekllIFxm
+W869PFSjoH1CIoSGZCLA75Md9FjIlgyB6L6RNb4q6vsOe+aYrfZh3eWM9dPWKIk89VkMrCly9Sw
dP/3LyC0N1LHnY9KmNxaT0WsyM9KrpCLz3MTt5Ebtct4jGo7t2L2kowA1AI+mqbE9N9Fn0rGufVI
Y6o3kr6F3doFzQRNEAO6VepfyROd2Q/8gdRa8ISFG9FJdpllANjbrcDdN3tW5oDh6dFXyw/lohBa
/l2jnnHbvjT17tfkF/u2Ycz3sNoFuojS1s8t3NpZrz38OeIdPevPSokiajKNHw1JTBSeetmcb+eU
MLtS2xt+csTVQwM66sEvGNi8Wzq+dC7drh5nLsb17tbkSIUOChbV4zAv2vBo5xynoHzSkk1aHFHq
XsWFT6XQcgKiqx+DGmJEHaoQrZyPJcReNmJ3G7pUBVE5v9FhdE++CRlWfcpgN9JIE/lgFTpy+NE4
nFmqn6dSwQONB+C3hJqFXVwtAFtqJOnHLBXnoemZDtbaD9X0R8AuDgp0unMQxCUaC/A4mezUWY+h
2dN7Nx818yojiGHwcDLFe/JLttRenvUCfVA+0O24BMmLxLk//LB1rlyTRNxaMkTzhgmJbRHje60v
xCs+UjzUjiyOqBIek32U4t83BDhV+kF1h51NmKoPblS9yi3JlrRkgm16h7sF99LDiB6Y2UTOG8Nd
S3b+qI6SCvVQnIfmU+5bGC+QZGUSIiFxw8qh/1L9x9S5B/7Nd1z3dor/rq9YaPHKROcxOKlxiVFE
N54zTXgtXFGYaGm3YAVP8NOY4FP7yWu3eiiP0sUcL86OrS+trrpmoKvpzrx3PLRKeMaxKu2FFGcU
xKgicKZBthgeBDe1wS5Qq7w7GVn9N21Na9XcW1a1ud8AcuH1a6bLukfnVjBn68ID5T0hD6guvekh
bZBBOhIVE6VUNILv3xn6Bb6pxrP25ieoUv6wBZP1yjZLTEGiFoz2Jq0Uwl9VIsotWewjkPNvo2kX
EmNoJ7M+/o5NBNU3kPHfcqa/5BXzjRAxR49Na2dtnCS/sfcVxVaJvoUmVXvFy+GB9LDvFbGCblZc
Uq3WIfmAJ/e+24e0lUwapQsSipBeSEBE3ykeUZ0Zg0keGFkVfwT0QC01QHJ/VSocg4NM9+Veq8k/
JyaOLlHePs2btLMQjTgR2dm0V5DpXgRWSKRcFyrx2COSELeyu8lRXMkwVCR/1DPsLDwt98VA6jwz
tFBcW0nK7N4W7ao0cZLqeOvDu7u2H1Jq68jsF6cc+S+YqcrfaUpj5nBzuM/zK/uayoUlCre+tDdg
JK/jOKqyBLWkwoSKNDvFsFZsah+G9GDHAGPKQaS3AW0ECiDuG2Utyw3l6JjU+83e23m14UoAlzhm
gusyMkasWizsOwrQ3kYALpt3y4Y4l5WEAaP/LoV93d/vicvD4o5P4osoCIxyZuEcN2dyTaDlGWuy
XpMeo4v8fgsWEF9QZcjFuS/3N4+wQVeaTZOsFqf+G+wBezOJ2C5kxgHmP7EocIhWyZ8W7txkAFm+
rJBvzSi6TkhliDBeBO6s00B+6S/V1Hmc9kWqJX0jT7nsnXGWKOj8IcG4bIAiFhhz8eexfqqjt6eU
ZInPqQxD9TA4tkU4KSoshGmkOwLMPqTMAzDvAyLyfmlQyNZSqX9QnQr2e60MGF3DrKXMS0Yoa6Q9
LU3UdeUhBn86DJKB0zMJ6W8gqbefplDgcWeUSahZpIZkTqatniNWfdwjg0Yu2gxQUQPeFX4mzzpw
WSbG9oa22bkTIgbDcC0AhkMOQmwjootcjNcbVZZ5odBjssv+PCmgFUGQFN4rrpIGhqgktgw4PBSg
26TJ2FeOaUaIn+P+zhUtSsdUlS7eibNGJOFfUz9uo0GY+u6BOUnHaKr0Fd70mDdEn6WcRy9cMcqU
bYLEzAklFcV6XBaA85W3THcwnkaPzs8QkPZURUkWdZPqMzyrf7jWhrCjnmPjPcwtxN3o9zTZZsjy
q1P2M7sCRwEJcVjFM29KxWpb/iD7Bkhh/wMWNfwcueP6uyCMsuIdHDTKQSE+T2RNMbOQQgQEIP9T
/xmcWlYe23lDGn8TSSZ4mzGm5FMTxz6YT41HPZBIa07yGNSnTg8hBJvgkY66jSuKCS8pKbrUEvlu
hk3cJT356XoBIB9txZZqsYWKVfsWU0ujKOaNj2dShcxd/QKc3haMZwHpIhOWZRb6RjMcXzOi/qt6
fBfDLB4vkeamm3IYEjcOo4zNO3ZelSiMxBf+GDJte39StREcyD6e5hJ8E3IXp8GGEg4kzBgoWdSV
VFZUTPtrxzQAw3N44knb42NqOO0gdXu4ytgK7OY850i8ttmOZ23jOwc692xCfwJNWoaLV+RLrQxS
JMEDiLgJF6uLjRs01/uqcYc4okYPQp/UHV85wyPDZSQIelldf8/mbFLnAPp3aec5Crir7lY/uUKX
qv5q7OvytoU3sG511spdsS32yU2EbAYdgEje17CriulaoQIOmggaeTMrdETg0cPP8ZZHebC7Dxxx
qekKUujiWnc1HSFojRbdKca4wXryVQJL0bbplESdi/hRtarbKGAPCqJPknSFM22oQhhD49b496tc
yYkuuSItESUFtmwhvI4ce12vI+epWwD95oJ4/ldKWYn6PuidkB+Ccc6PTj0FRqxx4I0FHzNrS9lF
T7tNHBaYLlKp16nDOK4arZzBAHerJXJo0WGYfO8KFP2miBmAYyD07ahmST85VZKUFCl8AMBGmnuC
949FAnWo6snTS5S/6y4P0EUMB98mvnzgyV/yZzYyrqTOKm0RJodaHc6eVt99M9nP3siZxdU8diuK
8v3j1idQ2MdyU6JjSepYtc58JytRUioWGFnuODeBKGxKgMJ2AxPNJPeFm38KtXuO+niCp/bNE4wy
NV569LQFT8L/4sSCSiPlwT928KeRVm1YF57+8m24nZ+pQMqmTAuFLdjCXqpmYqg7VkIodNwvzes1
ELZG2hCxP24v0Lg9hkEWCqVXJ1SIEvwxOXFNU7jbTI0Fv8x5DF2ysbmFs+GiIDlEK3Xdi1T4Ng10
I+Pg6DY0Z/NNFLJdyeJH+d1mFvMtCwOMJlSEwpyyN1Ebx5sysmJLFzNY8B1QWTexKTjo5vcj+O1N
02mcaVasX/gQcT8vUrF3qzWTrdTp6GI7XX5+MSxK17cpBETOxDZ8ZDL1qdeA86HLYVW5/Iz4Tu3M
yXkIPlkMVJq1VoikeQX+iehn+syAZe5zM/420rQHKoT/e4ui6vIOFbbJrgOkclsYS2HJ9abXviAW
O7sx+Z4GSbKyk/gGFnLBp3nt/+hmREsfBcrgDxbDnZAfZhb0ST2eOgt9wmDX470y/6r/XGxeV4C6
/cOa2k/ZItfSlb/jm4Ai0zzsHpKj0op5Xs58WOQzdVOkxtU3Ea2De3mFt/PQA629QvMqCyFPKE0U
OBrA4KpI+Tm1zTX0TvXGoe8clIVXAvtIA6XRwAyoL/k/W2s7mVXON9W1v7AAx5chJqIAU9Rqnw7m
eieNUP5sAFg9bX3XgqZafQ2gC165mz46U7IsOTaEUQDiYnra/oHOPbLY2EGdLAinrVsckGJjDxqq
jAPRz3yhcOGtdrPow4Pmk8YN38jSEeWHtYvQEIjV3nNzyXxrrKpwyV2ybCjfUzzcdNLyLeuSO9Sg
jlOFZKmeEmXKt2pvDI9duMCPJPuyq+HUGapb+30b9euz0L2y5uQG08VFSjRFOh4caO5/wiWm+aps
QnJ9s5jHuaJHNa7QBrQoanV+HjCERTmBBwVISXwRVbuvNHcTdbGBnqzw3mROdNJjWxbBBs3TkvWe
Gc1MtaUrfXCFYS4htAnmoAYASpGyHw1NRLuYoFCu+jfmfLpzv66a2Sdp8iyvS7YU3SOiAYZuraik
hD66aIRS12zRKefxBnM0+xKJo4/b8z7X0ciazqSbrZITiSUa1u/NUreQQ/ZpV9wY65qK8iXgkiml
0+vt6HKszsBtuXOt1gLhsjFDNuVEQpWUI6J5Lp71lpoXVGXevhVFYyIn2JVN5KAOhRYYlEAjedzL
PVCEWnhADInlg/2ElcB31I19Yf62G8+B5Jfz6K480rzhE/DLA5wFWEagl6iktY3gGnFdwyv4bW1t
nY8zVtz0axxzgXRMiwezPZzTm405mPnP5gL/80HXHS6//rs56takB8Qcxx+X7FKar8zNk8FAPLYi
H3LFTvJKBOwqiFICrHO9cezys+DPJN2b4Fk/JGk+XUwxZZ87PQ5TWkDglt7AvC52lS7A6eBB5JPJ
MC+DbnDrStEALhcRk+teKJNfPMtSGlctQFgYIf7Bfx0kO4QA0nK+03XYmHsngBcOHtftlgixnqiK
RnTlJZwalvttJ1Bf1nyjij4yN6ohufNUFqQu+gch9pquN8PP/6UKqGKHL8O8ExG8ZJJo8mJMR7fA
0j7bmZV1QeXgDBDOpRZUgWysnIME2izuKmFMOiwv9bBAK8twVO4PTrse6vUXE1k2WA4N4vylFq+P
HaFx3ubPkwZopZf2A8SWfnixOkJCJfN8fJaN87VvfOlIHgHpkHU9Gq5K97wExeLxQe2WYDRyUVpD
xvnpUSYVyde+o6sgfdtEDKtiZUzfz8u7hA4RdZEAU+mngLgbMJhRZAa5s3xj6F9vy+gr1cvhOfWM
nr7xKEEJG2hw8hZW8msjOpZzNcOmLyzot1tFACot1tqrqUSYcF6FX4L46K+utE/AzOATvtwzf7ju
UHHi0d/5nAGS15xhxFtrluCnleHUI6dh/NVSPWUPxJiG7O04YIpxfvKbWat2N+G792Y4tC8nmGSK
CB67mC8xJPVjAIfvXyMyn1m1MyJ2u1j+MZR2+fV1m0bZZRjBRGA7FZdNmVu8SVQeBDnq+OMgAWE7
lcPuwDMgjRBsylcDtV6bfZ7xxUujopYeBwBoZytxPB6UI18ic0zOPAq9IUc43b1odraXWTqhczz/
qvR0ieSw//zz7icZkppRjEZnv/K/8ey8jz+WWrR8oZ42V7vJAM7vQ8qWREmMdvPruLtF4P3WAD0+
GTB2kiGiKpgHYMLrl5Ou0WmjLqu6000NvWqYHz1iCaDQ4OKGTY29+iGLzkMTVlZQMxKr9txxgCbY
biCK1/AKdA2URfIATYx0AcH0KKdZTYdBlytK5/R22ZwJs9mc2sEkRWrDvZmwNvKdnX1Px+orPvnh
Rn462m9lQur/73Xp8qIGYb2BR6A9H+2n+mI516t3zrYwKW80/X3Wb9i56yQu5cmFj5X+PIHpkUI9
mJcd509gVqHjJg0uoZpCt3G6aY6WzsyaonjmFuC6VKxzpFRPUUXTlw71i9Tr4ktRWtGzomUBIujb
gsCzHdAyDz269tiR0GIAFzfYpXZ2Z0UZtxgGeeE5RQ3RRd5bj/NxX1zLdtBUFa14re79egdqZniw
d5qZyLQUkfGRKJcIBesCE/xOI6PJkGAsi2mAnBdHvCdhrDwyJmDFX5KPekRJsyJsORt7ZfCDkv+V
SxHmkJbbI01FaSjbaODSSJgZL2qxl1hEWgyV/GswetvAYPhlY8bCUh/IDGm0x3qfzPtpdkWgxeDO
fLOsDOj6zWy0JiEKZeSAGXT+gHSbANnt76jg1htNcZYtcWv+2WUphtaDGTwysYiuVY46v8Kb+b/x
6zAiw3wdxCDrBNG8nFygOh+X687BZkjAoafDbe8bol2GV8FxopaWu5QjepozdjHStKNMD8+WtvJf
QHlvCMyIjWkCrveQscHeu1ARsA8SDI9OP21ax9c/Rr9pMyT/IpZcGwH8TJUeCyUAOpbaepGN5Q20
jrHY5vpyC7FXvZ8OID+tRkjVqyQI8NgLEP7MCXrqX/ZtVmpTCtX+n91ZuaXknr7cbCWlEuHxW6s6
Z+Xu+3t1h1xTnad30GEkfv2n3Jrs9G3RK/uBX6SqOySvmgxbfgMEYRNwak7nReTDVBC5I4vixvy4
LqTEDztki2GS7I/PctPN+b1+N7yCWqnzs3Nr6Blnr3J/glT0IFpcXhApCZYxXxOczvC12836c+Qo
jGzAkNBQdRyr0IUC/evrPPfOZ98R19lMt5lR+HIkjj0yITjeW2Q3qCi3hmCc8lrhdywzDqkCp6o1
gfEJQbwt+Iw3tpf45+Hn/iRxmcfBZyfXXdlDFX+H9o4n6zgeyt9RZ7IU3CkzJpwcZiv4v9K+SzC/
aM5yISoRb9J5YsxiKN/wKC2tCg/bMMYLk6yPvW2NE0olCpBVPQ/DeC8vnHUj8ffSPEA6k4XVvWDT
BKTXsW3PaJeP0NadxNQILvFUxwBA8U+3qk8yveY06U24PU6riZAtRPg7YPMYh36pEt7adX8HKCBR
WcZ81+b85Pop0dai/3xCTUVp0om9SAAh2H+JlHZxio//eCnH1kUTdKSWXGif2kcwClost1HPWaQQ
YGEMZ1rYFQo2Ew9pa+Q5CJNbrgy/sRkjIWulQSTO0Nu/fz3pkp7Ky3UkJ4pHWOXsopEpWwL4biJA
5h8sff6XPg3bqGbHfPFlOjWBUkR3hTJoCcagQK3ahF6H7+c9sFHzB/s94vOPYrXM2xr6S2ALFj2L
2OUh88DkuHUwGgXBov+TAGQQhkjVIoRojGxj8OXYuqMo/jVWbIg795I9n5UwBENSwA95FV3EczEh
bxnL8v8uAwLtwRzUWyJHwCPnYc2u+JbRLA6NI7qjCqeO5xz0xeoiulPc0UZkwhi9v9WHb1bn5w9k
UA40a97tjAzGIeW1u5AVJto8+v552Hik/IKlV0PB2N6Hz0U+7gVg0nBCxo81fzRHgPjJ8/6TmUAm
ZTVq1TAawfiI2aeqgYpUOz137ndzQmDUCtkx/lYPRHM4+cHoayvNjwxCkecKfgb0ypEdz5XJEL+P
G8z4MWUxCXGVN4r49Zre4i0qdN3/wHLVQhTul6EcI/KySb6HX0qlFeQjeGV3Sh3fD/vT5ykuSzj1
A0oGOfNc1yu2xl8zCZFy/lESOK4mJLWln2XuBW6AhhkQDOvAm8yxjXxWlm6T1Xwj2zyFs7GOKo9A
ioWifJo8LBecYwevGQ7Wi57dYyuHRQ5AJ6ryfyD1uiETuiWrR+mVmldIfjMavo8HWFozfrh4QbTz
nBADFEZnGGqtGV44tYQWxMvAmPOpUvl1xwe4aHV3OZsavtYZMf5Gx/hVErAdwjAaotOLv/dd179w
0mSi+vdVhpBpAIDSWQRur+ZncwsNyRxJ8VGEpAxtDFbWjhyiD3fQEka/z+3iRC6GiUHUxoUFPwb7
81JgqE0mOmkSsF/0o3c24Y/FWpEJfDaj2gwx87En1GdBvDMLEraUDXyyh7kNQ9AIXuAFIZOD1WBN
alCM39VzaX1Ubg/vF4mfyJuPD+fDRpwAfRSoFdNzGahW1zubyhzmQBLDwte66qxUPClpAKp+0g2x
6hrCce/vYUl2tXsyc24xY5fozk5BbqKaxr1VjOODEvbCQrkPbDslB+lfGp0bSOZ0ZuM0QK5lpChb
OsTlnFFkKD+uDq00mw+OuqRp1HU4UnuUFG/JBIhB656rFRJGJVAhH4GOk3fb105JQF3f8RAhwFzi
M5PxRwoKED+KtZRU3mTaQHJusNnh3/6KZQdVrdjG43idGCquK/WVNwNqdcBanS5HqTbcNdspAD8A
hMrjho7m4d8mHmbeF9MljsiDOM33qHTPNNnT1knf+Cgbe7Mny8Dp3SeZdpWhwILmA17LOAgkq17B
WYLkgK2yegFglaZxQ28Sh+m2BJQwiMffj3OcARW1tYT5d8+ztNq0MMqHzpnR4vnb/eZblJtODO2d
6f7nV0cbKu3PCe0GpgAIRxrYkUrmqwInGyL0A8AxNs9SiHoFN/6BinTvxMRLAs6wCKsaici6fibW
XwFJ6+Qe180z7pP02cNersQ5x72XO1JmWZcWt1fxesXfCjns0LAROPnfObYhd0RFhzWVNshMhWOP
iKlXmSXV8EZ94Gvp96DebijP5h4165BlCzQ8O067xPcvyCbAzIjl9L39GTv/Ng+irNS+0SY0XJMM
1yUIThP+HkBv8GIrDbZfj6a6tN+AEuBedj7IMaYSpifxDligocaLewuNGYFW7WwG6qeiTZkrp/29
XHkEvpagHA7wnKWylOvkxW2yGNYBy/xlmeF9UpKM2yGhTK2NLdHLMIn3PiO1xwT3Y4mndbM8MXGN
+C/kCbhyQgq06bgA8vbNRIwBY9nECLRRyBYadgMpQtpCkDssyzDD4iDLUPEcvriP4QxSJz8PG/4p
VhFXO0kVTnA0P35mkalIMNShK96baXLSXOAWIAFzhB/JE5bROv4uAyHXWInbHFGMjktq+1Bv9KRJ
8i60wgwjlw8tvpj695Nk2UorjrYjmf5WV+CSle21KVIKJhbDjXmneRjeBulY6Foyey5aZ9eFfPH2
9VaLS9b6jA4HuMLVVmrF0BJYtWZ0mOEvGB/5GX8K5fxzmYP4bhxQrGQDAbwY3hFts9OmlQGn9VQw
jKImPaFYjvWOne0u63+Ty+6kjHD32P43Jdh4oiZCS3SXcwfDl8xvJRv7m7ngbzfg4IO9TDu/ssfQ
mXO2ZfIn23xEtIs9xYY+FXmk9rkMmdFfy79zYigd/VddJGJ1MjwGlKfug74TkpogMnaenPYApi6R
+PcbD88C++LDPD3ZYp97x3jtjJ5aJ60Pbjyai1WNS9OBJLL56QyF9rluHaCzusl0j2x/s2cvH7wY
3Q/E8GfTjwkrKFHEnx6lltUwDt5nuxi5g54y4KEw10XD2DKMClYZ0mWzxZKdgDP1YylVglRtH4R5
VJ4d5xZFEffLyI9WCtfDMxW6otGsQkeY4WqsJ+jWPP081dxZyQxCAqULFchdc5DegwNvA3skK8zV
36USVxNsYYftVybKjwVQe4LGYPmYjbOQ0rKCLK2t1dhy1pUGWLe6UWG0Fn3RVKff/N4XqAHOpIK8
esweXdTP5BQeI80c2rlgmXSJQgNELBoGDD/sP4wOVi4uPgqDAy9ygq3z2kjkayVy5+g6hp8lutw0
KCjgIvt0H4XGhaogcWqcEgLlCZHAMb/vV0aDurn0Lyex/VqtlKkalodvtkI2aY5+GXRXlIEwuv7l
qebdWrJckfLRuOvp4gcMIf8VYhWmbJje5iS4jmG3zh06o92FSIg0Ub6ZTRLw7TZWxX4Z2ro2lU56
nQ9EE9DkLzD1UcK7Ow8L/ICogsIC4eRq31Uw1cYOrDK+i19N9J8Mwuwi2Au51U8k70q686/mKtFJ
o9cCnSmRsee1sWtOYnMRsIbZKWomPmLuJasuOx+0mOQ6oPLUW6GzpRVJor23F7dsSA6+ZxMrolQI
AEcrsFuyN10xYMtdIFI2FvXQUeUtzP7eY7lvkUo+OMXIpL+z38EX21u3kAw2s52DYKwOVInfTXBC
sY3em6BTDlIBejeEc/KIzw+yBst3JaLG7E5HlmSycfHsSYjpIF0APhnBXJ+ixG1Rty+WKIYEwYDX
Fz7MSN8Xvnf7kRSjeD7NNsDnBYyGq06+1NpVK1mGfj+ZDrCrDXIfHIPwApho0xF/ThqTQWeEpdg6
zO+nP34kolBKLn1gnCfhMr1luTY9+f/F8iXGR8d79jpzLsiFgHMooUpuJFTg/hS15Z/Es4NbEB90
3hEtjQyEVnPdUpBEHyB6Cg0IOhEJMTQdvnlz4nncUxpCg41XdO9maB/ytnopIu6up9HnhVtURGD9
zPcKo2O1pmwjv/xXvKsPXFpOil3I7/zzk37B0/euuCE1tasE4kLu+ACyC5fUrDh0maSoWmkYATGJ
aQfF7vhIMwC4JQnzMQIKKhrx67DUgbMPRmBFfr4xzgxaXpn579vZfNrN15uAjE/jqyl5iYnGmMB5
Eiq/9Qf+z4B0bpHpx79DlRK/ZAl9B5UjhcG8653KzIipoXTzYbdH7kkWrA5g2J5xcFXeuRPuqtaB
Rm/QkxaxANRfT4jNGXeCAS9FXrLDVpfPxl3siFsgzuXbp2Io1XdVOWuyyoJtd3ocN6q+LpM72VCf
PHNj+02mAJ4+aVatnS8cXOUJ8jvfkkb7Reo5p3lz9mqvBg7xjpTioNpGE6uACdcOsB9CwILWxV4h
O+pIfeRQJHowPeRcEwTr3asXY7O5ryTL/qo8ndgAH/qTFPFo767ti9wk2mUKqqpARTQP14CechtU
iRVOstXHn4FpG8J0qWV7FA7ZjeSi8U8AlRfOxNxvESGi/4aEfn461WoOlhMQL4HJzH2La53qdN/h
hbH5gFK+as616N0NKbxUnEv/0R6141C+SSgerZDv59U2Lx2h3WJw0z5r0g2XbtwdeZcQvOWU5LiI
PhrwiOBHA2WlKlInEijS7uKH57biVgcuOcnVJDX0UUKQWXs9ozbzochvSFb+HGoNOF53ItC+v0pM
qtbwFQlBA4HJ8IQZtc6Vw+rULZQDQkesuk45FvgIeLlujN7H0re/nmz6zz8lC5rH2NENERztGW09
sSTujSmC3VrLDqKatOe5lCjSSnwcy0WmE+9L/UMeeGzFoISxXm1ucgm41/qiDNwhKMdQKLuBkEhh
pB8tBBpTJTVxIGa6Ws1mQsdqjbGcRgoNHEyDIJBUa6NBGnkjaeG1/t2yiw7CEBWdKJsfchkPt1/Y
XocLYOgcGHNJfjBtNNvmjizKGAeZYkbdJ73XpETj1rMXvq8oQLtLPU47z3421buW0O3jseHa74yc
XfbaHE0KJyQVnMUtdxMzqJtOUyzAyNVSNBgXyYEJdmIbwKN/YrYHeqb9C6qHgeETwBTG1YZCZkEz
gAJh64eDq0nlZxfpPkiiTHebgHBOy9P+2SytEHLq0BPRfEL6KzSWk4j48iwwUNhyOWJioiFQRfhI
twHA3QgR8EYDEDgbQtYHLrJrurQyl+E09B4BZjcbYwGny7pGZwX+X6/9mUssxWmqv/ALgrCsj/nh
lPuF7CbFwK4fb3lslUPBjbRGgFSwPbU028LjnHKBk2HI5ha9HOQUx37qPBpuH5Xpkju6/6DEMMpq
Z59qfivjx2hCgbXIOGkjwj+uP+OgS4n5DhLQaq6Uz8/0tfEdPImGZ0gOm+jPcebXk8/6JKiV/uld
UZ66MT4IF77gf1OTDokbhwr0Lam6Z7xSdQSSiNOXp3Qn/r0BdZSzHhw/6q7zpRYUc1Hy54JpTFOp
OW6vQR76L6i/poDfCm6NF+qfZkNUX8gjKMS6qvAIiVJi5TAa2KEKesr3R+fGqRB75Uc9pr+zMI3u
HQJJBIx+CLxNZFXPwpRucUNf3HN5p8LF5vz3hx9NeZz9f351M8Jdky1JiFpXZ5LDoNOozpBAhIUf
CQaBLwOeM43t7dE8nVxrlMDtZcRNnRDuoZRN96ca8yXw0wba8z+70cn9+ksjroFlrtPhlAWWhk1Q
0xu1jbNPhqYrrlWis+Dy2iS+gm9gGf51e5c2iwMKBgDllafVlI9mmvBITNSYGKbZ9KpNq3o1LqBw
pycx2yUxZD7D0fyBu3+wROeDD+qhHhsh38jLNjJoEZ6BBnpP7qO/swlBMnO7YQW9CIna1qpFR1vl
Z4OfJCZZ2rEQ8c624a1WSe0gf1rciuEdzLsnb1kQ7avA5gey27lcKz6ztanSd2RCo5cz6VwXWakC
ryyKbxYVT/+3i4yNu1+OwQEnZieSUP7U4O+03M7C/5NBKr5JxyP6zeOXM7n2FeKyHHso0qqTs+lw
8i1ZtbIOkIE+URntC2F+qrzoCZYK0XhMyk/U1mm7h8KAKDC5XRW/ODiLBb10zQIGhkEo14TGvWAm
zsdFGwAP5BaJgAlGlG0ILSl6ylJ/kLE2REVcWVJGbK9z+0U/qJaPbsb+D7t6+UNzRoe/NHxcLxeE
q5Cs5kxw1qON43/zuu8Fu2x+7SCVv0RTro9rsYfVhJy/9yRszC6LEHbHs2SDEafMAjy9nOYwcHF9
i868dFw71Rmeno26IyeTJNc3ZMW5eRN8Vle3RjpuFFEJSoYP0FHmN0mPGguxDfJ/+R/SXqtenKcf
OJSxSMPnYD3Hp59LpyseLUS/W/js0STxbm3WAPjOLO0LjknUgVxERt0LnMCDX4xydvnQSMQ7FGn/
gnOgH8zyjx2nRIxpE8iH0GCsmHK2JwaJUkCfgLSA8Askkc5P4RaKiEeC1iDHaYXXyNv4c4xi7QFK
1U8x46iOqPJorW10ctXWeYDAX0G1gUOfDDePAd1g5eXzi8DY3Ub8AwFyjk9tqjSvkeBTw0RXPML7
wndypJfUv0MgE+wGZHxiuP883TSNnfMszYsMyXk/1oatsTowR0Y/irvBfP4BGCHH5MsNFsE835F2
raCCl/8fO22+ZaXcZV6TOUgCI+DgQZOAPu/RkV2eDVYYEtZ78JAlSwj8zMRDklPEpaq2cL+K0rP2
mFqx27DjlQTnq20PKUtNQ9nIbqtAV9X+fnTEMCZMWfcVuuXXzbRbjyJFWY1pDfc+86n/DjRRWcxt
QdNzHquR5XbpE8A3FoTsHNvSaW7OJgVGccOXYnMGwlC/rHIhVEVd3nlqJnzPsxFSzE0t+kaR9TZ0
zFGQHeDf6shZ4G170j5qjrYf3gW55wdopyy6bBu1QFlgYFvaqqb+ugc4GxzZ6zZZant6y/aSL+jf
+r3sU4DhcCJ05zFF2Wbkj252IEzCeFklGYWyiunMKB9tCAZv8/cnzbCJER9W/gClmeyKzcbXTM8E
WEK9ece9U/XnheQitm68NeP8f02hhaOKHqotv0tTkpZjCchcU1MT9kxW5yWo+MAMuLn6VpfqX+4w
SUV7jP8YaEbnSRjnUagwVJJTHvVEQfRFaYk0nwDvVDlcAbxWggsag4NOe+o156sGM8tx8rboavbL
6xefjGmhchzNrrbdvsrpJdG/TPVZoAAx600sf8N6AThdI+sytoaB3slCrxcgfQGWYnC/sEzBejdM
6VujIbF9DO1zBA3lDhV/NCBZdwHIYcNnn9EoftNxB1ji/fnLs8H/b5J3uIeVdaHsA7GrwRGOFuw7
2/IotJVGYNzP+WfVChKDq/LnN3WYSrz65xhUHICg9OIemcqQ62+oXZ5seD6c8GlUcEYGCnNkPfQP
OOl8i0p7kfGHqj/o3rCO6M2QIzjeu9frn65t7PF+MjmZNHX3sgUnF/zPxGkbPn2GHyIPb4GLnB07
zpntNjZuq6KlqNg7HWtgq/AizmzYjlLU1jOi0EjvSTj+XTxFjdVpe6kui7hQGnqLXnV8svTEAR4V
AbYEa3g8z8skt4yHIemUAahQ+m4ikj8ZyT0EFqlAxM3COMGgneSAhmRS25cvK/XDW/RNde2MQK0B
cOIVrG5Bf4p2T8xFP0078NZ8Xn45nTqsg8O2J8uX9xjzYaXcLl0JMDewxOMGaBD5qtD7QWkvmlvp
/ujq2tGpFoNdYLGJ3p3blNJ6PBBcnU/c9uSMPDZt4s5WjBjnNxigv6dPPLabp1pUOFEIH8cTWUVo
DCkhhfkzAdq3JnZ4Q9ys6nnciy3AoIBO5ANP885WkCgBv1BP089gO/HCvzUw210bUQDx9bFBpjNW
tljI59Q3Hy0ReOxybmjnWEh5PsICXJsd559TCIFz64eaHvyT16J1ZRje4Hxw9Tzp6sYMS2VT9AMr
S+fvOH9ldhu4lE6eQyjIU0SRg/nxzdofpU/qju5QD7ADpRKv/esls2crq2uFXl+JY3PelTlSpV6s
LsSoVWsrEe6uSPHmOFws4YVixuw/rmchlqbXiIbVcDhVnBqlDQg1yNMXVmxFrc93qIi4gM209ndk
8iKe/PE9ku6o2AkSe2g8sYdo2qA+qSh3mOjNncStvWH44q1N37MIQoWDCdSSFmVM+mXp39Gc9inT
qZ6TAZ9i1+u2WZi+Rr6i/QfSKYxe8AQMk0UGOAXqewG2wtWuAx/YBOcXgE7TduGrfRlOGjrIOrvl
MvMrta9C2FWZ1zh9nAQFl6VcLGevUk+eaXo3M3g/cGAKcyePZUXvR8VnJAKswkVfO6beDDOrvNZz
DAEpYG30bXSEx5X/7Y3M7IQqqY0TFIaEqy84L2tOFxdxwewmHWK+yd5mA8gT9h9cxkaSSzjwX/HB
9S8krQvbvzQmc4pw6WMIkumbqjQD3fC1z1DpDgiVxuChfUCn9fHpHr3eRs9Egi8TfU7B1b19Gl3B
wNQ9/tfURGSR5644z2eeZTrhrK8EeK5gHzYeEx05dOxefJ0YgnFID5cMuakLQ7i6yksp1D8oFgxb
tyrh1NsU7QKqq1C2WR2YcW/r7fxmZExx6JqkCnCIvCmaXPUuG2FJtbEFeGH20ewIcGeOSs3Bb81B
ng++oz3PenuTnFufvL01/fUP88kQI0gFpH22Arwqg58RxuLz6b5WIdkEAhzUAm7ktLYZTT7HqdXX
GNMhFOWlpadTRUi0YkKqZN67hPpYcNeUcb2FtnsqROHbHu1TDyFDpwWj8bg9VrEBZJSKrEcb2Sw8
D5GTd4TkdY45KYM1doqNffw5tAS+A0qmu0AFw7XL+NnkD3P/W4G7aiX3w9+r2cLHk4qmW4VWlPU+
o5r5fR90+JZaILhOxuBBEF2vtZHCkxoKkX/6LM3J2EIv/n/N0574msSxI5gu6FCwanWADm0oDSf+
80O8HbVfLmhkM3SUUhBw22zKgRIPVSRCWQcw6KGsz/igwwg7/VJKBaUNyFEEYj5xfqQ0CJpb63PW
Q/okGFccihCC0KqXQBm4JkQjs231hUVhUFnHQvrHzdoOjbQ5QZ7XRjhuwzQXsmClDLOVX5r4Zato
0rtKS7RoyEwd4EGjGwpKlpA3IpM4gevUiPQKkrjvoLzewb9ea8NFlqYJ3cYuezL/1ckg1K678HmT
UerBriLHcmG3u+GGxlV169k/k/AJgmDnY2oun1nGJ4SC4oo6hyJfraIQIZWQHgb9T+5736tU7FAV
ud57Lgl1cEVLPm17hbxphNkXmw14BgIS1KzMbyDY1oGxw94E0a71D7PVAzbLWJEqxvlZhmFA3Z09
hi9RTQcN4nkHEz8MHslEX4vmMRiwZiaslzuhXZFXYfi/ueVdjnyhIyjvVto7k3E0OaLmiDYRvyuT
ZC2ISyCxXeJBkLK+TxqXJ5X5mjfZlRKkw2bU0Ygbt8aBAu7FYQxG6WN4PlZ8Q1r/HK5KeMnwA0Ua
w6uG3MS7S3gZiMlojfx90uDuZciLCvJVzVx3gLW3ugRHXPfjz/a8pAJrNH3/tkzJjnPlo8NwPMf2
XG9+JzGe+OJrc9hZ5fuyDEpD/aO9+01wmsc7cJYLucbbA+P5OfizDx58ak+t3aTZNApUNwp6KqDp
ia56cOO8MkSFivLaoC+pEHkNv+Uc1xWE85OmMPqH6PdTWgGbj1sXVgsy5RgK8S5foRO/OOAGOjf8
NH1BjNCy5gIf/YYBbz8sDRW56h+Kv2tPAHFlT/dLAUt3OJE4DgNuTRoKM2K+3+RUlifh1f/HMQWx
Qg9R8SFPHe7dKK8l1waDaAOD0DPoyyw9RqiMhrbd6g1RiZkjzkYXvoyOiJd67TN1H7c+9s7diKfa
CMqZ7LgwbmNy6qoZjeX0NZDAdz51u3IuiJrrG4rFSS+m1B3/jGP5c2ZCNSwLy0ct1SF65ZoYy/nd
S43dm1ox+3XSQi4HUkNxcJe7SugC27wv3xZz/2uWktPMSjcwY6CqWd2IIYL0EUKwDESNJXbYTbt9
FeLHbmk16KtMMSqx+034PYFS8xN5E2pDkXCkW99OeUlnUXGNk503QjYS77jDZUU4Km5CVbfotgSc
pPqIepV0hOG4LVCu0IIwrpQP4rQhKCYfEMxFPbKbwntTtQFX0O1RMyIXdCHuDUHULBz1UXXRLf60
aHejwPC/EIT2Q0mKPxenyXmZH77XkD1+syk0T8oJeWB9erFJCNE6Ge/gnJyHWJzdRuiidxrK/60U
7iC2TA0aho1LJ2pta58+FFKvrpQ3hMnnD55EPl89jeZlNbC1i1uJF4ahf7T5zCkoDvonPF5sSzqb
35l7Q+G4cXaTcCH7K09iT3vWUzMjk2XuyZFBYhUlqocs4SBcC44XRxYVsISq7RhWfvv9QgR+Kwy8
aZ7lqJYFRGj8Aj/1VeMJj/e45ExZtJzqFo9kT35zWgBfr+xBaHfei/zGy+y6+JedkzoM7a2Putlr
QqdrOW6BYYelUDbqSCqFJx/+mBW4vRnBZT50fW+Vlh/N+kp26TQNGkWhi3gk054JnnTg4zfJMLUO
q3qPeFFSFq5tSjVjLUg1uhj27uWZpA9Xkn2K/0P0Szl8Xs9ocWAfayRbUvjYdUZB/31Gv61IxYA4
IjWKj/3GgaTbF8F0Aw5Y3GCBSCoWnOUG983u/hyPIvX+wh2nBqE5irkBhOD/xjvnUO6Kso1CKHYa
OHu46YJ1g28F8Wnu6GK904UhbkVKsXOoB1EJdoZj6z3PBPXp/SXVAPvroeCjhfxtQYuGGbD/13Bm
GGi4JU0e/c4LOxGGhqHUSa91rmXB0MdefYTG/KMAgMyB3q3Imh2PPWTA3sP47NOll7gkkuHphksA
/NvvuJlg1c2EasjJAydJ4QcKOD1edYdJ+Zk7qKxHPRr2CWQpDKo5R8AVrZcNpFwRVagit+obmPpS
cfOLe4J1djsjxs20XJb8ZLbxBWTtOLSMBxO122sQ9JX2eKT1q8qE3YRzvY0nIvlf9WA8Cdqw2ruJ
p0tAltGMz+rPqOcBixcgHkyVYmh/2X+KF6FJii9ENJ1CkFQiMoY7UULl7rr26gbf4Ptw3k1RDv7s
KrP4oRtJertKsRuT1KetTSD4G0h0IKcCDL7Lbl6nqqULTL24PN3Me38ktAqpNYawLxHquHeNj15N
rGJfnlNccBeaecAs6purD+tHnh2GEP702i/b7jN2TQ2qdtF8utGs+7aDmrbJ0OWCLUnyZP5djSQx
LdS1uiqc0odhOhJ5VKYMAIqO4mN1F0KCwSukv62OUhaQ86kSxlt1CEcVgJCcYbb8Ddyea2cOW35N
ICvfIs4WqOJlOvgfIQu3JtwXua6ylqi5ix7MbataU0TCZaSD2xiQlVjqClq5JJnuTBv2I8jAja56
Mp8qjWhb2N/2Km11Bj4xtc1I6LLb0L6Hs2aQ2+ZCZ4WnCA/lEVjqtiV0tbJblAkPuKJ1Dahm2QwJ
n1vw408GEneEhEsr1QBz1kzPEU6dwgt3GzEhrjy6nJycLZvfSVjtvgmiLTXCHzaj0N3tb1FEyvYD
8fLVoFlFOGp4/XtL1kH2851ZN5y8D3XP4jI3drFVjozT6yVUJ3pU25SH2XN6+THly7h2NQr/sqTK
iHODiLaYXhIDYvht5Nk7tqiFlsy4EsgytHBu+0sjXlalZE6kHfkjLlNwVyZlrS6Fr5tJTUOZpuD0
0pN2o9/xmOFamhBkwYy4B477VF4jgHstUZcMlgeaGnTaxgjo4v+sEi4psyWOYBzov+mYZUUHGe6x
OKJgUHv4/Tw4+fTCNwJW3rkbM/LuMQ7UVvYN+KAKmWoH23p9BePqq06EoqAoAJytrwEF73s6XofC
DRhhRKNmfj21+uf9pAGa9T7lPkKT0oK25sIi10fJvQ0tTzFrR+IDDpH3eKPrxLfJvMbmf1UFUuJA
9a0LCpdQxrdnZKfL0JQKJZ8yKVH92atXIeP58NDuhU2d/afrFxufYgVTkqkTkpepbKAGH8TK0vTZ
u9A9GNLNL0+QwlXUBxBzvdCCvDf3foaHmAEg6iwNPB1GjE1XVdhvBtrNvG55HCBLWWbN3S0365iN
CEaY34qqWNDhc5QJlbO1E7k2LgKz8kN/SYc0Tz93K+JWSkRdeN5VG4ez5/bbuoMDU/gt7xpTg+VS
uM3Q7/nbviNatKanffF7E+3BRLUO0FpJnnj3MReypSCXMVhXNQWsts00C6gVIAd8o04rKbvtg8ko
1EWGbRQarXPUi291fy4wq4Zix4ytYvU4rcrpzsKXJOMOXkpIxZt11nkWKaDLCo9We7ndP9fO7vdk
J0FgkWQ7huC/0IWzt5NcJXaHDSECvAXY68AqTd7h43cFe28c2X8qJbf/nYXwFJgvWdtVY3iUQJEP
6u5cE5Ic5DlLEE9R9+cZOwS15QdUKE+xX6728nD054ezbupsxT83yFXBi9iJW8Mzc3UcbQRF71Xt
0W9xhrmOslT3KZPbdWrNKduxkUEfXQsX5YbiSyDVT1HCb5qHGLU2ognK76BTX4T2rUgeTNgt0QSj
hGVxgySr4awGbZ6Ub9FvnnFhFKttyqzxxGZ8sog/Ondi6i3SZci7PPTb38h5jraw29YZ6AQkAraU
EMPoH8krmX+T+kH1W/yWyQ2Jc/Ga7EprgeA14/yla1lpl8nqa0JG0a4gf1yLXieR42lU1X6l3d0K
j4C7Hic7P76GWJkKpVZxRfnUHrjsDXeE/aRmJRzfBSSfw8jOUYwfRa/2Hc3o2MbBG/6EDFPpdTkd
ewep+PxLZg2i9VQkNesPMJL21ur65ie+ewXMDHrQnaIIO0oLam8mvgAvLK0j4jvBvrj9/bLl44vo
OEecwQlcNaIG6yYR7fen5p7Pn/DS7E1135pYtBGS6z/WE3eGI0IqLx/r63thLzRuYuP2QXqH7EXc
WL8XnFBFcoCdMXCH3Zhnu3F9Oy6R/guSCXeNBoW4AVuXW/I0UCuaP4kh/VDoyzSUF0EKYialQFzT
U752UwZWirRZwb52HaRbwG51iXVCXH3uR2YGGyNnYfZVgb57odyA0+N6Cmd4WOxNme8vy9oGHCYK
pjDH5V0EnsOQkT/OUr3lg0K0Gm1F8giRc5omRaYkjgB9S/8Iw4QSEiRzMTcLTbphV6n4YtmKdXzP
DmDFdjY6c+b+4UQl3PgY5i/wHUt4YAjwGVKBczaNPff/gsoXv0h9LOUP8moMzk1bMYoleFOobqIc
11EX+50D/qUOu70l8qIKaQKaEWs9CydY3XO7AkEK8hPzzS43r4VT8r1hat5AuTXqV+PxONtDYihM
RC0anfTssIvaA4QFtpQNUUL1VTVQorJ+mptcs4s7O1JBhdcnLJypqveLeNXxzMENv75jZhLK2vd5
x3+3PV6gYvokm8S+1dtCHndan2MeoSz7uP94cRJkhpQVgq8U6VjQPWB/6Y/uKO8y8tsBmNFY5en7
4EhncqIOGhqD2+fH5u0/9qOxitAz62Ru6vytFdytqAENtUbPPq+TK5Q6U/QOLcIMcR9N2xuqWMk1
rx9YxjJf7i1Gq7gUKlAyf5JmL046HRhMQDOcpaeF5p0uqq9J0MChCATkOu/++MK7Z6N5USM4jlzc
rdIU+9xNoU5cM0rziT9+vS0wRjqoVYDxfvLFVWp9R7EXsMfaxdybb5qXIVdD/kPoqtxrjd3C4e29
RWj08mJKEwU1ojp/5s3aT/CZNP7MXaooyaKLyQsAJ4xNkqdR1uUxgz/7xR5eeI9EjjrOIDJHtLK9
rjPOFsKvNoTcMcyHDW5NrBCgaX7jpCWr0T5A9Tf60mQxRZ5KB56nNPP/cQs01NNi/ryscRA5I51j
0rnWgZfR3e2FWSqI0qo1iFqi1StLGI6tpJlkSjqMPVBsA6amnGJVcB3NurMjqsKrXuJL8X2Wi73F
iANepGRXcONeu0y+PCIjCB78KKgCpSfCJDjt3KLCcSSSl6jDIvp3avg6vz6QAi0v+ARmEUH/YGyY
+1PHH+5wsqViL0XpiKFjcE7CH0M4bW6VPVRChhuByKaw5bKaqoQXxLuAT5ulq3/UM7KPu82bRlzF
j8QsQiC4PVMhV0X5bfSmVduiBu9qM7NJigmyntV+UWrQpgmOYY6ocNS/thqVffw7vCeQzawS01/L
kFP4dEiOKPx17qKwJWGQ8OsahMor2Z2Zvfii+GNbwgCVvhUyiaOUcM2i6mBQNoUQiJGzs68DmX7g
EdshEwNA1TWJsaFUNUTwjztdcAqJ2cSRIZbfvpXzTa2uRKwB67G0IPZpHgv/G+7sVKJH1KTesfeH
Q0aahj/rJFDSphL2mBuc8HrT26GJlck71yc1cq3cZTT5cEN0t5FI110lMQb0c1Y4V4AbtaPc4wH8
UQg1qCkN0XUUovey2Ja6Mz/KFynHmNGPs+ktDwynDHdGzyjq3GyTYByA6dS+y6ktWFB8wGZQKVga
wLYPeZIpSFbsDaUQNpU/xC/0289rNe7wTUL8xjQKkkPcIjPmQ8Zbp8bqa22pLjBWGM8OCAw0ggcQ
bDK6yp8ZaDIpByHsDr4i7R7+e+ckrr0jZwXcsxMsrqJoT90ts5eXyedlOVIXhfMuj2rV6rvzzAun
lN1GytyFS+Iy1AI9ceruvToi6nGtC3Jqq5Wuh/pFMPYhMqAfYsRLyb8y7OkhqTuaQ9jJqY8FxDgx
bcsQUL0tPyFoJrHSWPYEPUX8bMyAlau8zSW/v6eos9U3A1lmkLA7WHjhN7tH1oFRuFmz5K6yAuVU
5KIA9c6Eu6TklWyixGy1GHEfMSsFhT2IPZZPOybwdzTSHj1qaXWhnbMMmTDZesKnLCdro69W/dEN
5auO6jmeQU9eWfcIgvjI5YlGyGkkeVUs1JP8fJqMeTwHBNc4eIwLX31ZfxsLn++BGDTF6S0LDbrl
NrAndWw4C8U0DycEW0N+957x1vj9bImrd2kwVnNyNagFPI0oiO/PvrLrDkH39hcUR1USlKozyhwm
Clu1T/gNu04fJv00Wv1aUvFDpE7yWgNXeHjAcPu+VYtRqIErMLQgpgbddenW202aLdSiDH598qAP
XPaUUitHSHGuVWSci/DdNpHpN+394CU3xErWv29C+DhtatQJ4BN9MZxR53pYDZcdUyMkODW7+vdR
pLMRbNAqt4/grQiau6e5PrCIQ7Ye6YB9O+KVRmPsJ/P4QEM03E0G6QhQLY/LKCIb8yE1uW20tlnV
TvZ2JGj90CEKCyRrI3Lhzyd4uAS+uMDJGCQ8tD7XCdNrA/9WwppYKtInd3PUr4Jlz2rKTspHPehl
v6JmwmgrCJbvaNiaDkM0KMj62IU2a1G/nXxEhK89xVJb8X1WZmIjzlkvRu1o6ZCTwrpnekGxKWbT
14v/w3qhRDBfcgoQ7xomtJIrq6AclfXEpExM9FSbS0Os/Lx751J5pWTLDHUXEoJ4uvQCVpMC1AqL
3+YlcBePYKZeju9FipwyxE3XTKU8D81R4JPO6J0nUfmo2N3XmElY3zaK/RIyzZ7677sU72f5LPPg
i0LeTngpBMdpK83Gq5s5xI5fguNwAxnPIT7WVETUZJMyGF5TX/I6NgT7YlbQC9gGYy/1YSOoylVv
c+SCTNE+cGHuJap4Mhh7fh4Sjluqy8al5V8WMTYU9zzerOZWIdjXcTisuISwiEXjf6w9q3DkMMOB
v2ZVDdoJzWxWbT8lxcvY1y3QLCPDLkmA2SmVRMvG5eH9CRsjb5EflMghRhtSaUCBIUz5T5ZRA1g0
2m2k72vqIlXRz9jJKFFHb/82ObVTSHuAXmzleAQFnoRGPpBH1ol3F97ELjzfGfBC34r1m8JDoecp
GkzD9RaznFcFa8eb+UR6cFQfSkGTQO3DTJhzanoprBJ/ZxvNaHai1zE3xVyfGkboVCiiRTvNgkCF
3JCIF7G7GWF6A2fb7EMYgmfkuakM7PUYFbASgXlqfYCjYgvlsI+zDCJ5r2UKH9peSyfURzxhXJpy
L4JudWn6ORsNSzd79SCRDNk1/fDWmBJ86ZpSJlKKtLURFiBwMo5DoNjkwZwzqh8yQh5Fyr0SfPw2
NVW6vMUxvWR0g23COhQMvVGIfv8ezGpZiitSS2AN7pTtQzi6q6zS+1RGKDEQY7nlTwDmDbpW+Cf2
R021okrBk57qrbl5pCCKk6jhkZVDLXUpHeC9vIQI4BiXHMi8fGvM/UCIs2iHgxWp2dmE3QpRMqRg
pfB0VtiuzHoGo/tIA6bvCKTD6fV0aTytOfvP7aM/Mcls1jM7AOiQUqjxpvuRF+cHN34HDa9LOsri
bvZ19ToDNq9SPBom64GDUZU5oIDPafLwlhUxMmriK+KdVK0Q0ImNqldxvv25HBD8E7W6NirgqeQB
Vc8R1zcmiII6ve3SNF9va+ZDGmC+UdNN9MGLMZBfI4wrCkYHrfA8gh9+SMT7KfKugu2Emq3SiWvu
NzmutAH9MW5AcczhWuuMwxlNydHQLYSNJNlgBK6JIzGE5BJGSH8K77RPQ7xSyS4fDVcCn3j1k/vO
io6gSIhhCgfRfNSKaV64ne0eN314pWiaLDOnOJXkUKVi8I+mOZXphBTETY6I5W+Az4syFmN0HRcq
HY/gwm0txjmcdgvdETCnpLcowuKoaPS+QOhXBh8GoO3/ht6+2QayEcxuygEHglewCCjkH1H/j0YP
PKS+EzHc3pDK99R+J4GR2YualnD8OeM1rnnWVSRVArytsW6qmMJduuKhuIr9hd6dW5P4dS5xC40I
Iu+QS8sYI/NbgpErrlxTHpQIZ47/DWXQH+qFj3V/0L7J/e9jEb7iPVpEu1LDwo6r9P0ZZoIomXGt
JRNM7WuuG0+S2t/Pbt7lc3VZ4F42+K1maoIdCL6k6Idcr6K/iDd0+Jzjt0UdWn7p+vCpZEdKUgDC
kXI1MO+xfnBd5dvP51qel6vzwyS+WxBm7LLbxBy/EjYw/yjiiGVKirOgEc27dlXz5oPMcPGRoBxC
1z+CWm2yfMhK4kyXLJn9xOtWC47jB9OLwcr17anZG8UXXGzsObBc2BlB6F+0/aDonO9ZzNmaWdQv
djiWH1swJ2n/d5K/wsVNRAzwXo7u5pVjJXoUSKtadlglZN7aUNr8yrW0hhuV2Pe/d2fGNmvQQLco
78Zcom+7cqTwnZN1wxZkYZTUp7Vt4lNGJnhTR368xkCEhaPnit0LdHST4R4Xe+wCoehR0s3WzGHO
lp5xkxwjBkMNjYPcevAEayPKHorUlEjDW9hPGLTPGvKuyE6nlfD0oqcObduSfp2nM29m5HXrw4XW
QqZDcpFEJLWuaGu4z+puQqrXypPnjxahYqFIrtoeKPW7zeGSXhR1wY19EWquLKJxb4dxSVe27Mlz
3GeoPJAkpQdtbNUxWtAl54WGia99f9p/574AD8Np+gxOsipTfFeeqFpFidvZ6D6c3JdFo3z/uNBr
gzh9kIkOeFwGv4Qg9Jz06Tn1lXxLrbcDQLsGiHJMfxqPbvrj0uas/kEer/14VUG3Scj42YLbcCNO
kzDLLNh2u13HuIRi7spvLxh4D+NdDFOg+FeelfMO5jchGWYeAhl2RwD5TZMU6g2bOqDXrXfhuW3n
QkmeDutzqvVWgVx7p3Ea3DtbsPlqgoQ8lTOyN5u/E4zITe5AvEp8IdE7LFOUx7apcmEtaPWcE++B
faCGVJDkRo+4+WlBE4GF8mTHxM1fYrJRsIjftGZi85Y7p5fVmAnDwOaTdY7TaOn3tYRNTLzHEA2K
mPvs4KsQ3lXKlzA/0lGeQfON+AxX8vUqB4v4U7wXfrFxMQtn/Gk3stdAlrJul/DpQT30PehSve7y
AjDTmm7K7aDNHF/zio11SwJYKrdT9nDBZcROLj4LzepzYknHWD/asqiAUR+nnFiym/M48GLLT4kc
cBrYlmoFpspc0hCzQdrKLuGgHjt3NlAG4kfcOvq9Q+GtUG8WWz2/KpJd8ZD8ksy4YQAxsI3izH6y
TWTkNGewA27slo7q+3ObX2npUEzBW076kCQm84aCrwDvF6Pxj/1WWuh8lY1SKQEZFhnZFLbHIm2a
wWon7q2rr8oyV5DtXVc8LGb//QG9pi/1mhb+pa71ijHeLR5/lvmYIKI481EGQADk+ln+miiZ0NrF
Nmk0fBtN8NaYVwXYYvK7sL3Adr8L8rZDjn7QQw9l09AE/rQtB7aureVUYYXUwVJF9hsltKPhx044
QSg5/udu2BEWaCwKSDcUU5Hw3VDf/JqjQHCciDdwpr4wLy/X+NeR9C+tNlC+fP7CeWq1SroOQSTy
19C+i5QDB0zQY3WL2Ia1p8j3pm96GqT+D4gwIZRuLz8sMvAKuj7VHoMNGIn7X+9O6+IrNZiYnyAz
BmuKkk1Gb0MFY7fqnyfkn58z5n+YJmTZxRs2Nfw7mSpPYGJhcizNAt2CYx2H5Amm4Ecm9oxHkGai
gRA2Z01iMGdsXnGheM3eZrvfQLpZ2uxo798xC4ahplTtQ13hglLaiInYwHear/fN1pwFxMPBpnmN
emAjiKi0iZYWsDGooin5+4bZnj3zrBARsSR44ZkjBgPJ19+Pygy4DFRLLB3Zky5uJ7jy6qGu9iPl
6TpUHHEG4ISB4sCudNaX62FTxckBLW6e61m2iQJ2UXztHr+/9GRCtRQXjeoyQGqcQKEmSSlQz0VK
+gqCQejwt3jExlxHsz+s15SGCbBpJgM+RfeCcdqUsxK2CGxmAdK1824K/aPK8BurIfix7jT5a4ZO
9987VlweROXxtIhZeBEiH3rHCg+zKNs3KdD2bfSm/HnZSVyszMHm4KAKjGQCh8qo238n+A91Ci3R
o1qtJjXIGblT4MLuqYBVYeyiQwoHTimJSaL8v5o8tMr4oHZUriSko4s3gqGccbCBTHovZQlcnwRz
E0PkwkAtqYlT5yirgvRmz3qmUtGgsMt+cgB8Yd6zExSRbxyjMzo4Zwn0B5Eraf+3qDfKkQB3Sb4m
oRuhDz015hYXKttWCG40Oudp4qb5PjkRU8I2Q2dnyNYHzpkYm8UQf1BErvYu59BvLwiHFKVCpq/g
PxE/IzV4091Xf6MFiMpTawkxvyHpE4KPhCscyEXzX1CSaVpY2hypGT1M9iA/V5/fu4zbuK4GFrxQ
cOQF/qgVqmR/WlNWNs/pEtaHwv0AcvokCTK6YnbLNP8mtS3H+1GZTw3O/scO4EVVXyXkYdjiJ1ln
Zr61oarpMEHv2kgVl3V15Wl2IXZPHI2v9f7/DBrhLyNuDr8pcehqoTHYVYHg2+0x7ID2Q+N/KZq/
neU75f7pWRbPJ3ennYDVuIJYJhHQ7f8UJXeY41LzCYsrRua47u6IN6fxp5nFPnR9qiqQRo+/aEmI
eb6lu9810RwvUAgGW1Kgk7Pfja3KBPvmRcVOxVmGykEF98z/1x+hsJsLKHK80BIHS3JG1b9GokIf
Cu075Grt3EFon4D/76nGslnZVYes8NvyoCU9/8I2rBcjdHRCxdHlwxGdDke7DJKuvFGxRtx4SLy9
S56foYpFz7bm24YHGDFZWHrpLbqABb4bwCjAYcZrgtZCbbXF9WMvgyzhoir5XmskYLSiQIDezgXM
wxngd9gSjhyVsud+M21WDa+SZS+xKfwJfXV48TERtre0bTawPTMMuMZoIq99xeSp7F6dTbUq0bkq
r8haGJByNNUpldiKi2WZX5q5Q79VXtvNxz04QUD3yvinjcxljkbyLgWaGbuuJtxrhcE+fY1aAxc/
lxChrd1+IXWPdxCIoDEzY+tnJa5nbrBLjYPWjon+wJinJtdHFMJCZ0XjMlx5nxWgrcqfae23ieoM
oSwQp432TrbDe/WpONvyXPtQfFBWbhIagKJwBQw3UF6XfTZKfx8NuKACAI1+KjwzH29nEcqvSEQt
YLPSWO5/i3wEgmpVc1b4b+FaBV8PMnt/NgtvQljJPBcu49GdAfGdZ5C8Z59LNe6RmsCWhpuFSoOp
Lrw97Q8hy9BTEig7Wy946amimJUSkH/ZqSsdbQ+k5qCOgDd3Py8PMWaSD2nLX9w9ie74In9VsShz
7i2oJGagC2UubXZFeZAxyAw5T92izHAORdouDjQdhPyTcnFUCqnhl7RoN4PZKw/IUrhSP4+upxf1
oGTTdLmadZN3eOyvW0p5BJOtlB+qaI2r66qR6KWgBrG4wCPhBFui7EGOffC7RehHATNuUtKbJOi9
q4EX665pi5bIkPvGz6zZKOtGiYbnNszeVCgFVWqtyRQb15C/9lEMq2VxIW18ZJHWGKWCvjYk0srB
adpG/1Kjgoqe0fQ9yCnR5BwMKkR0xc5ZkIBrJF8JDrs8sOql0IVGWQUJjtV6mggU/mR4I+PTdM2y
V1yAqNIvgOoH+/ibse74bL+504Z31heJomyfLVKwbSlFedwrfRSJ1+WGEpznBI88Acv2YJg7DrXY
9D4aCy+sGJlPfXeloA+f1DkmsldlVFkKwUQMEg1XCbQ4Lh8sfoKJwRoSg3nYQp738JbSri6sMTkY
hnIRUYQpBuBIyut8TonPH+dXZhXTYhLLhk5LSNhDy5dFJycdkFJs9ZyErmQ51STdZvg3NVkK9D9m
0qVk5hXjTEbH4I+fSLO7WWRtbivsVvEb7P7lpd1nyODUXDNpdJetao8kkNrv5Uft/O8K78h3h0De
GlABDC88dnkJVlTONlN/DeiFKcr3SeqQDoQ7FYILMKiUhfHbRtL/M8B3Hs8eE2rM3UigngEW06gY
mldGDEW86+mZLtPwwDMuAMF97Qf9I4d/KH+ZRgZFfsu1elHuYJ+ItIk2scZJasejA2S7TP/FxOZ2
Ise6ajbVGm9NrAlMb19nkuAgLk95OXEjmLDEgh+DBEpQO7nRmUJzoohqUtvietmlqltuu+gC5aDT
XNmeN4w5hS5UIoaA3vrtA1/vCi3NLWXje4QAqLkzLe1Y7dLCJAjuIE1aS+TeCADm6Yl6KyV8526E
5H87HiVepOXNYbnPB46a6jOu176/nSMPiO8YRiDoI21mL6bPkEHa8YGinMhc50X2JJ+7DcMVtTq9
9E/l439wMf0bFwsUtkib3wshh80pjESKKwckNzSuQ9dsefGXnFhQVBdw3ae0KjrChh6vS0jmJ5aR
4WaEeq+QvyAWhz7Y1wJ2wK6q2/N3QZIZJUUkPAyjF9qS8d7GcRcEJnotdq5bj2xOZ9/sMvq/J873
gKkLzh2S+rK8l9ZJeIQRwmxUflHBEMjBYMGdRHE/+UJUZDrf29MbSFrGRHh3z3mkUZCUJ4JV//au
E/znztjfj/lmNhHgPtIv0d4Q09f7gdMWfX+G/WbCAKP1K3nASDuLaVqeOK902YPm4itpiVnjsee8
Qd8ycO2jPUkDZ480z+5us8wZpvy7vbJqIvYqcKqvPv47nZrW1pZdsZVmH7Dj3r7EYmgw919FUKXJ
Tb4A564cQmutUgaOQ4qv1rfd+HFh1/IJqt5mdA5QFddLxWXR0UvVDq4u0aau201/8vnmF+iNgCzS
luijH1DNPZ2YXfgfBv2DvXFlDFNnzGWwe0oBD7y3noHA2F0QTbiBuvWtwixsdVuKaO2N6PZUr51L
gx8+hd5fz/7zSt/dNSy4gAjeTYbmEAW4Yzo3jWtvrQ6YQm0PscKf+pjJ17WL6SMGjyV3eshFYCUC
DefXqqxcIPSlPtlttfU4hIuZWeqsmQnZP36RE96+Z+Faxtz+S19urkPYCeOyswmDF2U2JChfEse/
qmbe/h/9WEBN0LbfPliGFQwBsxZTTgoRteWH05NUohpVpyasAwyAKSxlP9SWPScvY7m4dno6tuUg
LxL9yPHOg0d7jNndhfEKQ0wuuz5ZhUnMkjSuIzfG5nPjmgFQeHyXpm7rmWiwyoYLu+d181FFAGWJ
Olst3z1VePquENbgjfHoP44/cPzOG0F2IoyGybN4y6Hn4XEaPmGHFFQNF9M8FJ1NwOTJNJmpT05w
jmGFtAH9DnVqgvRB/5BsjwaTzpPO0k+k0DVOcyyuBQGGA9Q/5er3+p12tMgAAmCuDlDhh/aZOJCw
4+npi8fp4jJ3ziUUvdKLNo4AdnweCrBisFIdzYwHzNQaLBovTHcJAWAtrqjdnZfkSPCinpOKEx05
Qz0sTYtTF0YznTOpP/mGvb4FfZJKJXLutYg5c/aQmX9SzKw2PAGfQKXYQ+ug7+ZZp/WHcUN3rfUS
V26QbLHOknryW54ArzXnlPlxunNBv0m8Fuq8nl0QYfwwIyXR9tqQpZe4hC3D3gqNywJyJ0dVU+b6
YOQJbjt5bnnVmpWupo3KzZNy9gGaiauEe4b3nZ0qv2bWhdxXJGTKVNxIPJ9Y/+2/+7jOVh1Ade1P
xQRfIFa20g+5ZtxVDitiCmMSlE6YPaAMQKyZfbfWxFwNOKgJt9kGNM8gHkDYkS7zV6m6EZxpfsWd
0lHjGurXpkRslldYRREeG2AT5l+3suFitJhjeWrbA93D6QY4Gw3AKU9MWmCeqvJptykrNOGqB++G
Wrfh+ZmUe/iEwcHZPpZ73+siVTnZ3wpJWlnzdN/rEjEe02vBUvvhJjrrh+OB8+lQR+ccaAYVweIm
+9dk/fl4kdshspXqrqw6GHkd/hrjWPD+w2XnCPVO20bloJPUh/tptsNnVlcCLP7CYpRGxOwE2mQ1
CNoRqdcDQHkUDYqc5wH29UD9g2Osk6QnqfyZNkwuI8dN1yvQsjITDkJYb0TN1fBGgV/uM1htIoTO
go9YwNE6FU6RNCJetcKekkLtrh3Z4jhpb53AdHRzAnwSKIRX/EenSi2Cvf3PFtVA3Q+wo18pdNza
zM8rjeG8s7cDAHmwa8MUYOxCsXXIqbgHGjf1S/eBb+O0jVBRFqbE8nDEJTaKwY8e8uQnqTZSM5IX
83PaiXhMai8yMQF6E76cnMl7JF59tIk0DeoDgY0dUw7UGruRrwyN5g7jUsXeeBUVe6sdu+kVsmcQ
OdojRXmQx3sE+O3FzXcgAfHzmjXbrZSTIqTW7asXML0Toyu8N6Lzs+SpFc6MmAZcBtQ0SVvhVcUM
akgrsNNbPswha+YcmItBhDKJJD1/gQ8DEHFEKKyUq7z03NoUCsYh5O2Hhd/PFTu1zPs9f9bOd8c3
ZJf9xJOxKFsfS79HP880xrtjPwT4DV3Vjs8EB87Zx2tszndcD4EqxqmG/hoc704110c/7iNfD6Z1
X8UGQLxICG3ihpXcV4R+qit6ld4IbmO4pq3wZe11RQGpTfWvN/GgZAQFdAVkxC+JY/7k8wPaIkR2
k4jUS/FnI3IVMSTszgJ0yqkVyzVJV7wO+gg+VPzm4GHWndIlXO1BV2phQ5mLCJOISUwci3Iyi8pR
Ge2Ofkc9/l0sRdWwfP/JOOC4m1LDmthju4JUvwbzNMka6JK98qjRKLZfdorScrZAunCCQvmMAsX8
UdOawV4VcBUaKr7gSD22MoX7Dn9svb//F5pVr5g/qva0CxU7eSxOyX0lrgIuRFWUMjyZgDoOWISH
zrdcN4gpWBZLM73UgzjYjbjPdpV26b/yaYcr0+vC+m2v+xPRLYxPPLp+TFqzGXk4e8CQnOTxyHcg
VVsjm5qjq08kju/+XsyDDZif6jn1OBF/uJXLSvo6wq0SSpp4dlgI+OpQgEExdCLs3gAcFiQ3OzSw
o7nt8KDaHDQ+xGqeAfUbPJD5MPF+fE4dGu5xixuYQCOp0Mvdi7MihjJ8nltDMyJhS7i14h69rDaJ
goRl8thpNRHc0h1Jdq0HJejcADmtW807cRyvrZWUtoOgLYyZfDEszuW6FA7GKWwnIFJnFw7ezalL
8Tury/gBDlN3xSEqFsfcfAREPtwyVwfE7CeokQQWkcD9LTArrZ90CQ8g+bhIfv4xehGzwyFKoZ1/
+GDfy3ABCPeb2Nxppv0GP/Wb8KK+IQYmMrJUCUdkK1nxuI3Jg7ZjIpY6zDQdqVA+RFfpwOSLHihw
V6pl9tthlBf8yYuLXa1g82BmOFLloRnNOAbveEHxV/Xl9/agjO8yaWhDcGRaqD8xoGAvQvy7BUn0
n9+amlMXY0Is1hI324JXR1z89e0vlGJtGIGLABD9KHy1Ip0gcA5TMvxt2hMH+iDl0gJ0bCAXHi8x
4yuHnMPo36bKwaWl2S5lgxPdI+8riOTxMVm23/j38saXsQYJq0I8FmQBe3rh+rOOalIo5vzHmyDt
CC9JOpxNmVI5lLpGGwIVNdZhB0FjKCYqhyDj9dVfHDHkuXIP/yzC59AfKAuTCzS/9CzUNtv6/SUy
aTurX5XYR7BcmWrGuc2Q+MjgZgF5tJw9M619I4S/6zQ/O8Gu/ly9W+FPJasFQw9FxFCqJAAvuKMN
FOkvJwYPF+oVXEOgNOAfdSMYtIaG3fXzhfeQBL17nLAEnGu1QZxWjwYjBU8kNd4ngctz41t5AoDY
pDr99eo+0jdkP/HylU6uTA3QFJSu5vkZzIACSwtweyBmGE6XLu6hN3Syin+SlgjGeHpYz5l0ph3R
C9GZ+ZqX868EuyGpA3vnut7ttLU2ieYzYsdR2xi6PWAHysI9i6ddDLgD7rHjUEXEHX2myV45wANn
/DLfCqMx4bLXaZGci7mJCqW6/lwiCpHpUFCKEhURqCljenhjYdajwMHdFu8iNrWlJYlUS/ye6Qhl
AEYN2Doy+V5rwurMTR4BqdwX53fgyAdHcfW2GoFRh8855y3D4tK5cDJ2RRNNa2YYOOtTzhnXEl1M
scEijMraDRzTL2g9itYGa7tN1GvTmi63Hpv5IBvLn9TxM4tyrZY/6ZD9ZEArEGBFnxV8Lo6hNgj/
RvFvIv76QZWM43jfj/lChUsRHORZB95HIeF4TlMFygt4azVwseAQ6kzbeRu5VwRaxgBLXq1JdWQ/
W8XM0pQYUo1H/CA4ecOjAKG+1vi0qHBpvGS4VTQ51InoovZE8uc5kwjeH2YiGZYAcGQOTxC8BNm2
mm2RBhdNxkG17KpykLQRx36C9AkzaaC4hYBTT17FUng//3yeWUWHGcXtOnN2M2irRZpHntOAJ8AC
Rmbs+94snONoXiV8+C7/9jRsK0StUbE2VT1Kq5j0tyqj82xYUmckyDrLtcoScX/2/REjM28tIS+X
Iiafi6Z41zGJOYshmV/4y/D/u5/SCuvSTc9SaEg0SZ/yl/aTSt6r8PXAWrmRWXM8m/LhkWBohqmm
rLF/0mfBhMFRmEhaneXdoEhvXRBef5tdPwxwf9qxiYwyyZ+0oyADLfUOfUQvUAN8jGHRcDa3O/fr
641JAfuO7GYz5Syaz2+/auzLt8wRsvlbpduEClmZo/gTiwUm5m6FTK5YVlTl7Nf4h+sOv6IZZojW
ndCyqWSpVvsud3qRkgzs5ynAtOuQs6fQuyF0K+bFdJVwnh+3kKXeSMQ7tvWz2Uvz7/OwRobFCjZX
SBJ9zBqYVMSknYhrPtJbzqsB3wbV8rEzqbNarS+CESveYjpLVyYpVI1L/coTRMYd4hXaZOpaj25G
tGaRovBsmrsapMaPbAyE7IfLeNGwfQdE4vIOwuAVjSvt31uwW3G3tv/lj7OdC04ClOiO7jvao80f
1xcixsZbuBVp6T89PCy6eHh2DfKi2CCjVm0Ewac/O9U3Gpw+XZocFhxt/aloG1B9hAqEOkB/OYkr
n5p5+3SymfrYoiXUWDJExH6mMOkgP6DlldrSHjHiepZ8DAZPw/KlvzXm8DfYM2cPS6vaiF58/G/C
wS99u9b/ty97cDPOziUkedZw9b5d2ZocQm3ff/euyLYuSjvgL8kPy5inuCW73520YNxt5vSUq09P
Sl/hPvb3LezNWXAmD9bIBSIr6tSKXx2qJ2GCxkIZZcTGaNWlo8feXxx5rVx6v6xSH5bvubxpLikl
n3UwdcF/j0dC384RJy0vD0Txde6etxlj6T53mzKtscBwXuI0Sy0DTXsst8JYX6zixswSVlxBSomL
R8IAZiAaeyUkvFgtpm8eJ/5ee8a3QC9aY0EUizNedSLgEO6wp61Ms2tvX8wm1d8Ho99+xOq2pDkB
atd4ZDyoBf1sM6RmnIVJlERSHY/V8LOelw2OhDdztTq+0N+kQiurEJvfHZPQ0YUN3RbbutRBsXjm
sUPG6NyhwJfLZze7husBgFdSEtV1+Y7c781O0qG6TpB9quaG8ASd78NvNbflq43XnM/eWTXZhbO4
7qjMXYH/o9x5Mc+h5tZaTIUTtXwFAExDkEQ6jvFcPvBER+iQutDqsXHWYFE0HS9HwF82LqgTWgJR
5mcIEXUOUOgghN2xaTmZ6oVTs2K1HUSSfY7JI/42YSXf0OQAa6GaN2anDUhvR16mYPT+8aiVmyh2
9JGIsBMnffdkiJIFCGhzxuutDRzj30eWC3baEXRwG49sokNl1qwsWNkoh6i+XyQRHKunRzgv6ISf
OgxiIya2dyrlaX9R5dw7BMw7pW6/WdfY2D5UUgzX1V//IZq+Ra7H5JfyLYjcN/k3NUSKqNM6GrIE
QoqtiI2Pb2RgdZHGssVWVJzc9pPgZQ+dmYFkqOIL8Hri1Pxt1GWKbh+P7NFuwl1CdTOYUmSFMXv7
7JF3wOa+qnpEUGHFJ1PAZAzluENh2O/yk1RbxJsVSE7Uw79f5xg7Ls9+Zfj42SgXirtvuMaeq5nB
BZIyWYKV0UrFV8B9ZDJIJYml0fFBSRnJo+oXJdcO/AwhVdAPyY0cxRYitaSSffEP74RPpcv4B3iA
+M3S2ZHVHPQk/yAv87NpGh0Mn0TSLghlxWNGw2mrTyjuRxDdnXwD5sUr71Vr5ROBbiFVSRT+caqH
NgNtdhtVXjnjOHAK8oPjnvOy71RF+WyrTXERa2ZrnSNSk5rhXzp/mMzRZrZ/yVQnm7tM+yrlODqe
DF9SX8yvZZcev12gYMKynWuSe8XlP9B0r9Bt8Yp317j1WLTabCaS65EByr4qIa1fnwMar1nW30qu
i1iLlr/vchDiEC2u+87hfJ9cD5VO4kvcrVuZT9OTHuEzzWJibhG3T2Q2MH8SSY8yxBFg+4rlLJnd
ExV10xoEDK/9rP9Pg56CsZglKJMar52rtcNl5JCYNVxY6R8dqdLLow14Ds9LecaDOKLKZxV6EDMQ
ap9tBRssq0RozBp3nSbpK8yGAIHag6Vi2K7u724991GwPdjoMsbXeuP3BxFb2bNyZfzsry/YLNv7
sjujyKo1nAJfGUNI+vNgrA4r9Mh0wibBzf+LV3Ex/J4c2PO7abJAXuQRK2WUnvYRis1d6GMUbbYZ
1Kx14M1Sm+F6eRPzg5bz+9oWVgh8YZHK9CRaFRH/dGriHL4xQabVahD68WXlxGeJMUlyMGaDPDPt
p3/Ze9I8ujyzq+3Xi3N/NqOVKo7yt2OuQk3eF68yGKZOlpE06Ca/wQILD0u/ccGgiKZjpNotEIdh
iUCYm0k+h4ei/Lcc33ON4mLWrCa2tJpAi0elgL3/OCFsAdySuS15D9z1vZ5A90K/DUMqF05TlPlZ
MtAt5W9ByTjGZUager71lPA2csr8kA2IoUEG9OypzkW/dEDVbla/vVhtPGxF+x5B5SPLIuYOOS73
3pa3/Yq7WJQg4sxGELFN8P9y35Th0OvrP/nhHvLZhHwYEAQ+R+SIwGqfh8mujR6WuM+Ba+Op5nJX
eLZcGSq+ANiI9bhebj5giyIAIMs45z7zaEGIXdAnhcHwtcEamVLZaLmWg8eVdnx8SA8Au+IPWtdu
znCrUb2/fIkpbWu92Lp/DF9fiF23UUIZmurR1kbweswVRr/ndX40rMf/nFqBQlQoL2NtAEmvgghC
ElDx6hq5nokfpfk/6GT35Voe7cmK+NxmPZkLBfDbZtQOkq97GtbwfWdHo9cW0gJudVkwsff9WHgL
LzcQXdYK/I9F8aSI8negBlj4rV2oq8QN1gyzzwRL8Gz/d/HUfG3o0JQtTPicKkcib7aPUJYD4q2J
N1Ej+zFbmyCBNIJMyfX6KGYdBw96JyMnKtpxH7MgNTXxiOVs7AqlylM8kZp/VT8E/1u+p6os1ZGG
rZaXudCGhm3ulWlDwwq+S1F+dQjuhog5zqUimT7qH5BaEUAKKDeH2LviQO+lIPMEcL6Lno5bhez4
SIN94P1tl7qg/tPh/hWNpLlfx5IKb6GCQs8avr2o3gtne5Y+UrTt4CbcWK9JZxMOmdnK/VxBbFpv
Jx2oFlxfz7hOGojhtim832pwjE0uMQBQ+f2gnfbRVwh0dSf7Hkp98FqM62n3yCqD6sPyOd1NsRb3
mdy0/a48Z7QpYsYe6mvTLBVmfv+8/PRnXhZrHlcZGZj0c0ZalCnC35ZO7iyhb+Y+nJ+ULeiYscjU
BVu5quiFKEjjAMD95cd9E9jehHsXHKzmTvyJL6Q78ff8Vlwl5KhHQ9Y7Bhw8iviAfCX4yBK+ET66
NZ81ETp/QZWCATeyC99tvBLX59YNWc2BufuCdZJPHQhbgfTRLq/OY1aJl2Se6c+mkyyyyOI3jdBQ
FcEEBr9WFJoCniUdLlLsthdMJNisr6XTA56FcM5KlgqknVbG90TRATG9Cx7lyErAWIzqIHyhsBmy
M6H9YXDQyxh49E9qZkNL0U4S8WS7LGpiM0vjXBj0Tf9Rd4QXFzRKdpprRcVIbDe4F9XpLwKbOm57
uOPf/9Zs0BDabgIFTLpx07G8DOj7BAWlb6S0wJNzv9HM9VKnB6sVeCy3ebfyTP9L7o6PM32JSIbf
xu9naqgbrumm2JBhpDp1zuof1Co8pwE1FQ/eaI3awkhe6vjINY3lSMIxnK/6ufbvPxNiZtMkNfCz
noR0UzZ6yZtgfztVR9Hn3Zkfdui8He1QVmL0mLiLtZcGBMsdgeCvCmdTaWd9fLWTOPHDE1V3WaZ+
RAkt0vygI3K8cc+O7x+IyV0GbyU7IWnF3cLsitU7uNjtb65N7SMB2uk8vThnoMDcfCku+a5gcT5w
CEYzaeC0STkP90gtNYdQnjyt5vDps72t9ZLoXN4C5AfNulXBLoND/hNNkbuygz3NbqHF5ZVEOnq2
9I9y0IuHsvF0LWJsrv5Fwmq9ax7NtY1o8XZ7PwZiZU2heDhYeD4B2s0bPS85fB+RPR2NGNYYFvnJ
2/xgsG5P0/yrxZL60waGHJQyujXhUB6D3PHFMBTUMILHcAQk64GNhcRCDE/JbFKsvvnV3yZU29uH
KZoP+KNbja3IYj/ltIcPvQ7vntOxHET4Po95MBaYtXX066iJGgltDlUklKyw4dZT+k6RjDIJQ7yC
Km6QLCo7r53PMJ1fcjsvnTcLMddk+OM63gbeNewdtSKm4gVxN3/7MW8qW+zlmkw5Qt3If2TjSXnq
CfParxTuJK8+hh4riJs2YjAwFYMPGooXtbHrzNfrwNX0KqXlI6fgc74vwSB9inreywnRyglHN6XJ
2VOY7QTizv5hX1oUJeB+fCt+iINzR3ukZd2BU0QyiArG4HR6QF8Hgljc3w4IJ7pBJ4+hr3GfIOt7
iXUJWTasvOwyCAHFMMUJdknMQP7kOcZN4T82r5FowhvCF6rB9S3LxqCflO35hmeoVkRJn370LwhQ
KdctbV5gzh3b3AD/EkkJMCOwrgu51SQ9/VLEuMpWfRzNI6cnfdxzUtFCR8tSBnAf7cYTqkv6dEep
gLRR9Qu5WOW++8GJ+iIn0CkxEltip2wdyVu3csIT4/xJTqIyTbPZ9tIn5J/EveR/nWr1OrM4n2lS
OiuniyZGX3ZCWlIBBuSGmQs0xCUhWSI6veObiWrK7k0T/j1UymDwF9QBzSCKgv9TloMUR2q0Sk/A
CbpJ9aokpnazWrZNr7Pkgp1Kxlz/YDoUaLruWNpechQKq56fdcSZL/NsWbLa7Qn+G7GCT/pu2UCS
gABv8LthMOenitQfbEq3muoZUpsfFH25hgRb1XMP3eehJY3Du0e+zdtE05z/5z3mBoICiCAOeZOk
WIgiyZIlQu8KGJvmi3Z0ahCXKROH6cFyjgi+KR+HAsgzepE4iJSlG1dUV9acPxNugk8fv92JAZT0
z7BRzKZFG5Xus7+gRiXoYMW2VDIxXKWaSmD3nNtiNT+U5/AOkUJ8Tf47LigSSvtbH01yUMOhy+NO
11+UCKl+iPUaxnQQhZnhiYfBG4J72kmxkP5eSA1yrUhcQhgNKrvh7iWyDNK2FVC0hkvk0ncRQ/Tl
zOY8ADf23l4r46gxKGxUDgn5pr7sN6p/6WGWCR8pnPs4nnXOs1acEMQlJ7nc0+B03GGTIJ6WFRr2
LFJv85LoIQLVw9k2IfHL3hp9gHh4E8bbeaXZ9p6zSq1v4eR0vdLDXjMFWV6zAPYdw/LwVYgbp6q7
9TfnpqXJHZZf9cZHqgK5iB2o2VH/rGGjZRfBVa8aZRmgE63JtN98/1P2ipdAO/WjFLsv65hWTIPm
qd8u7OKwhSBAxubq0ll3G57Q9k51VgjHW7aoL3h4rBepmGcBdUXj2WkwOYk6J7CxyrMRme3tpERZ
zgsM+VITu7vxhoxNb2UY3JvFtNsWNTZaLZhLY6rmJ0+9sqJnDSgX6oWULhW25o4c4cPXxL72cJC+
TFBMA6GoOs9oHLUOevE0ty8eHxdISM77c9X44gVM/cjuZ3Rpa1LW77HGYVLL9/edQPO+yE0sclas
TaLszncmpgb73nn0WO8TicyZ7/vCiROI4IoFIyXOMaDE6/Tuwy12ubmvfMsBVnV/YAMZvU810Gmu
frqKBZN1Lca/PzPnLfPMF0rDN3/E5iQr+1LdSnuercodokq4bTcEVSSMwt6cNEDsSYPEJPEoOeK5
Gn+m1ebEYDFEtNOgRkINXgIGXMNont8NolP9GE/8+0f3O1JiQA3nnb1ekQhwbJc/AF79CRKOHBVH
sN2sHWL2kuV4SBp5a5Fe+fKn5Qq6lkjJ+QJy/UOHqnqsl1HDJo2KKLo9BhgUTCC9xZuCBUkZVTdX
ssYk86KcU+axikSkHNMndGHGdh9US4GAgwqWp+XdVQtX7+rFLmjUVhpBYW1c20ccca3ta0n+TYZx
edNkxJ5Ub7MLM6wIBfWdAIkEvEuxToKJxIAl21x5c6DRC601XE4qb7oEHJ4kR0kg/ItxL7LJfzNC
IKqISSrSrcI2bbr6G4wxxtbY8yrHDWdG8379g3ElNcLOH+9cnhTPfqZDEVLWSiGummnh8mGLQun2
vytP+xW94RhNRAEIw5OiD2/Yn/jatODrpZmY/lDsyS7lqkTIpuidK02M/S38VJRgymzrDJHKgxDi
Rt3vBpUu3nAMRA3osp1G115FHdahInPHMi5qMh/6LYorNGKGv3gD0cUOduPMEEAWixFKo9snz71c
YcwbpprGsteaBgFdzM4uf7hiWly8rypNiBPfNFo5sOntdZNaMEpszhODasgyruPQhksZghZGbggX
zsycK7GGYWkvN3fke2jPjkoQ9S0HBGapZ6LAcG7anOm8hpVzMw+6351BYYDH9ahWmmZ/mOWbLrZt
dB4lCnbP6X6aoQlDsfLJJk1EsGTszD+UprZkL0mbRJt2cwNXSXBVSCxHKPNhGFiW+nLOrwdMt61u
T+GZSGkbhwJItPY5GdFlRS4qzUhcNPvfbxYOo9J7ZAPT3EMPgp5V3alF0Mv/ZAe0eRTgO43L0Sk5
XX7CLeh5sUH4dWxmboioqD6BefRPygvLq6FMsMIF0Oi/OvHEc5TO5tyr1cfuxpGQZl2lzKH0Y5gG
evs83lGcBOHlDxeTEGY4JMb4t91oVLfmcuAml2fy0Bsu7aP7sspvw8KJPmT5ERj5m4rgxgRi+MjF
PYSq/+vWnSiWOFOqqOUyM/suVJeNyPpflN7gFVfFOpaooTJVghJHwbV4nr9ruDqqAvZAeSrri3DO
zoY/GQjsJ/nj/esO/jWYyjQ097CEVP2PjJVT6UBPHvQtcWcvaZfDPGQsr+SIyvWO1/elYNgxS104
vfRXYmLQilCS2FXl44t09SEHX54VWbC0ndVYwTovXymPQZhZlTI8AgLiVEKM9Yhg7uglLfVaYoPr
+ABFn5/3uFAFTdbi7CCoZgERupU75+uJsQEPPGUyBkXs7qRFFettRN9dxxRloOQXZeK7+85gAuMq
moou86i2u1PFgFpyaUDYkh2udNH2fuV5xVGrhJ3fwcqfHkSNthpdyDOg67McmDsDwLdtkif2EGtg
n93AAdnj65cf2rdguoiFu/DicjuyosU764FmN48rd0xNuC48E15vF4KFunvppSKcHqRmDGviug44
WkDd3Zza9bMuD49+fw4Sn230tr4nceQs5EWkEjcP5M/qoQnV/5dlFwoT2pkmTSfrbrjtyWxweEvA
jaoPHis8rCcvjJmyoniakTpIi3osTN4tOYwYtR0cvdJ8atg6p0F99lZvjYVJ4A0cZIocB5qHSrKv
BneVRD4cqaWPjpln+JbLhpjZi7aXoXG7jCuFqadyLhk65J5SJxK/ZDsHxQBei88hVjoOCpBleEhk
YB+j2+zKLBm96kTw4qw4oJTfl4J2Hh6mZgCsZtOkDb+E1Kb8gvYQZxSeXmTNp6bGqh54n4//7Epn
rOXud6W0ZDwZmHNjsxcPlTif0jVICKqjYl3xYluNuJ1v1iARfxW3nYy8K8tcx53KL+BiybLh/vex
JF8ELjKvM0uFBdkoxhrtBHsrJLUM65KwYCYpz+MpjVkM3sQU76gq4WDWNKRHC/7DLxtpfC6UsRfQ
N7lqb5+GuP2YHroxOryj7nHAEXgblFh8QcZ0RAkL0yrSKngETfUtpH6n2B6g5BUH5hchpEaW0PBc
+uY6p7jfYte2RUhAQWd/sCNP5E0zK2bpXaoKSUFkLygUK23/PyM4sSE8H14Q/IpSWlga4cOgso57
oAK2eK6VWb12AU4vJG9hrb2mZhcQU8Mw18EuzjvJEwk1u7jWRDzi4ldNmT9FxtdgxXP329FFPJGr
LGwZNraaiumFfQ84oF8J6pL1j4KynO5I/wwmHtz8E2+G1enTSOZ8iBW+uEyy2YkjdH8sjeMSDBNg
k++nup+hDxok4peeOuN4V72iLHRQjwvyKNjf9SuC8DAomD17EDZ32pXeL4YLSo/X729HD9yRkvcq
/AMtli4nxtIhqkDVIB03sqPH+ft8Y+FZInseEGnGHtw0yN1HegMc1ZmQx6s64KCCLhpV+Ft7SOS7
aYDF2+ptgpZhDf1UzBbeOcYoeRUCb28ktaCcVuRR8eeU8+qZ0vM2kn3tIE+aqvlAFxKnVCtg36RH
gtVL1fEQjsL4158TKrpQff8V1bK1QzELvyGoAcCMR6EuRXMx/ZQVmOaShl3S/bkiZkX9V7avetIS
2GilvMRimBO4pFrGzBrdTquBTR435h5ZC1ROEqgetngs/R05dpvCPpPn1IISxJCiWkRy6oPc3KXF
SohHUI7l3gkVmmRLTpBGhA1QLF1DYurWvYRRd6EvaWpadhDO0EMiB9Ev2+c8X/pyVRhcc1C3TPC3
NNt6Xjw0TiGDNNkPcGDmqM4Kyxr0pxBhQ6eP19e3Jkp2O/jAvv0qLsWhbAPdapnDwGjLpSfBjt9M
wVYQpsurTbTX4z4kW4vMO34BGrE/dbrd5dRFwvdefrkCHvrJbtaBXy8vuoxp9iaKYod8voYUDAAI
Ajl8hUeGuX6/bxA46XCNojZP7VGA5xmJDXiICq18XW+zDAnq47rQR9UaiIHcDzhKa/7OXm8Gjsqx
Z7nM/eTkbcAqmNjfwmdMa3yzpfLY4O9i2dP4wm5VchG1pL7vXx1NZhegaDSY+5GroNaknnRW0+D9
zseCN5xqrXRn38ywvp8aOYFX9v9nLiutjskQsQ3eLSWson9U+YP0jUe5vO04cqu3TqciS9/Me3OU
SD5ijSKM2/NTahGkjT0Z4wMj4iClPHa32GKc7uQmkVgfFJBTVm+jDV+/hNy3BvFs20dEMMKnUraX
1bAhZS6BUpVMDq18EQjyV9uQceCqYfiHlw1oLO+DzBGfXHX5iRRA02X8LznwKFJan7D9ZPsBrE+e
CnuKuiDSsvNKU1cABKIeDyssHmfJwZQ34uZw00eOIBEp8trF21wOgz+SBq8F0Ph/FfalM8d+R8Fs
7YCalBSMhmKkD5l3GHtaw0Y4jzOG6+I0Mzxf1pppudYSVsBHSOoqwdD/aFgnjZIagx3DVEXRJm2i
4VC3LXJsS1s65etFcuAnVo+dEQVP0l/I2VorgwCRneUe6F1WAfd+p/679RHjYk0B0lsakhotQ6LT
ng7ueeJdUxwFe3vyrgyjfrh7GwPinq2DjeITYExBqkp5F5IWrtL8rLVcYcNYzIaPL/2rncwYQvn8
SKVD4rB7A+60u30gCTNXl7ugNFrM6TkYWgCwMuhJxaHqaKMBQki09n+03RpTYPaKmfhYK3MIP4w9
G7CNbIP5eDFzgEvaOYLz9yB/2t3lbXZjlKdfirq+HxLtBJoar4k45Ep/0huxtoYOZ+HsUlUwGCFA
/8NIWb9zBAelYYKKwHIbr0TdF4NaVPsxULiK4TVQqZI240rQpd2b8IAg836aQ+GcpQ7r/NvIqz1p
NZrQvAvpU91zvEZHlNCkMQ0BRfZasFHZPJpK4+jGuDITP2ZXNv/nX4kL3nJmxEZY9HurIB4vDD6Y
oNBHjsoF1EYap55Z4885WpIIrmK622X74A3Ah2laEIVVYDu2e8roHGmSlYskSdGpuoS13XAfNaF0
y7VNIqQbQWq0r8mtOZPuf7TFDsDcd+l6VOgYaVGxcbS61bL5FqIUz8EzJRenYN/Voxy8yq/bfvpS
YO5CwI2waYsAScgvukLxGFvfpq9bovUZpOQVO/G2dXmv3OUDoKOoKeREkEypJguQ8pY1aA+Lh518
JKx3t6txdYMHR//PsRzlNFrkD3pOaID0W03Rxco4umJy0tW2IdSNDAvNvYUrpEaXNe4Mr4veOe6G
wG4CN34iugwF1hVaUTeEsHtziypEtP/LEcYUheh9XkqgrPPnHC0LVrXEyPVTT/rc5NapG76RZVbP
Zcn0GNlh6gxH+jgeSqzK5Ai935FaTwdM702x8ClQ76N3r9Q34fcKgcOn8jy8RL6WaOKU1gIH5a3N
Zj39hcImEPZ1PZs+9CzkrTbysDlbFfit57lW9yXKH7UfpC7w2cRi13rs/ZosRsWsG5DxLd2CHlK6
+gjys96/t62dJiHgZlVD2sMat6LZWN3stAvcN1XUgWk9H/PrftM5c6OZeYlaegjlJ6L9c/6Ue18a
24su3dU/DW8zW8k30HoL6Jxmc0ZGAa66OzlKWy+h/b5z0ZrY0DhJPW/51DadH+/9Ko/ui0R3w9gV
JAHHV8VFr7SlCRpYtZpMxN52cd7t0kTcim1c6SAYk2SBWmOMO9v7Ozn1qeAyua2XmttWcP6U7OzZ
6EeAJYqy8CtoCl1SqvgrjQNVprj4v5CC/dMd4hR6kLl36wgWY3eWZmiICW6dONhcG4/pMHJwZ7of
8bKJ02GWkxXNSlSHVI/Z38j0ASP7eIHf0WXfUbex9WC05ZqDl11LfBL+5pp3byMnv9tyQQC+qese
ciduQaULHnHTF95sOftL3cwWrC3ua+4djBv9Z2Hs6Wavd2ZSbnFNSbdl6ZvaFKV5MH6TV/PtXlWy
Eu35pwwJMb+FdSuEKE/tfHAEMt9Cdgh4nukFD6y4XtQy500sYaZbDoS0N4uYMix2adHIq8wYOowB
eq1TxYMbEaAHzFPupfJfxtnzXhUH7RXSKc8I/fuvP2d1QWjLrMyXnFFhhiRSjk6o17/0ilb1pIqP
aQ3D/ehbnwyQ+4SISYpgUaoRnlPk7ekBIYOelQRvM367tFEwRwGlYkUKDIQ+FCnXIEnFOQXSe9xM
VrdrFobDhfH9OeqWenxhlG2C78EKfisRDs5jA3rTGipMWj98BNws/nCzda6xXb6j2eNVPRti1oyU
bKxscyeNdBP1mRPGOiyTwR7YTuxgjJbkSj8SNmwbNOl/512yDKZeylAWBvlA2GQXOdDKR5CKuqWz
p7TXsXlpFj+8B6isBRpd/NIbkh/fcjovMnO6qF6d9gh5U6Czc3xVqzgS2EYJnkecRSmMPL8bdo8y
Le0l+RZLO6iE51Wdds65w2eMBMUA5F6jn5L1/d8oH8Y57oOBs3qehV2ILBBJE+znMjExvgVFFPGX
pEUhvFHEKVlK628rHbLLSEqqVtv0zE4rIV5vkr/Xdc//+mv3qtxMpWYMsDnvrJ7auUWgFNbLwpXy
IezE61k15biANUbNDyOKKUzqAU6XSLWKHk01gbTAGHTLqvlw9KLIHNh0dqYrII+yBm8nDJ1pqQsF
EbqJUZ+wiAv9eC1oryw59kali2QN6A0Hp02Yz2ywJAFYYX0luVF0a3VZKLLFi4hx+IkAxT0eHGQP
uOCbwG1FWwOsOMve3J/ttEjHQpHFoz/bES2vr+UOWiAqCsXdEWtIkoJRUoGgbs8zLi/5faI8sLuo
QvFPuep2hcBIAlRDcSRNB06zIljYWOR6x32vGkAkyWyeBm3fVAnKQARooXItDCuqp4WUGEXNB1eh
5P/If3aqZpAj0rnsntU1boTKODtU23AQK7kvc0jzKQLi9iqpl3bTBpk7Z20KDJrPAXSeOwNZ/fvq
Ie399cEZdxy3d/zbjk++rLQ33HJx9XDZgxIwmPjdccOYa+7Dulga7xfVTz/mLjX86kjudhPuhRpa
GsaY5yt2eSXiQe4Zjicz316wTx9vDAvsQnkZrYmTbS9UEpPjnIPMlwqTmfU+sldJtOQ0TLqBqP2V
GeOprpC8gX9TGwuzCUaq4epTezw1kQXqZsTUMFYacxfwhPme6jz7n2jAQJDoeb3o9RurA1xDJtLu
yX5x8/tlAiHfwpkFwZb26YVqca47okOEhe+HToyIo1Ta7sxfsqkMiyDRf0NFQ9C7P4q02jdonoFD
2UoBdvzHi+RrYJ74+imCFzKIru52sJ+EGwfpzZTyCrhqo1uZIx3gle61Y4DUC5d9SBrTuhp5U2Af
PwPYCrDAaNK+PYQIife8wlwA1KB2vjRtMzQOdh9px2knZwisuimG68YcnNsF1/GNi8fzJHIpy9cj
xs72wA3AUnJ8tnG9QaXjMB6UHpeAxmjD1AMry59Jiz0B139gBo2GUjDvbfSTyQIRMdksLzP7cFDF
IgeEQpkkrLJN+mR64Uekf4Kb5ngWKVJAkCXXXHJEtoXFfvlE6RUQppSM7Ais3SwJqdDBeDWCfRuc
6PzvhvhSZ/g+yPuvNasUQYNmDbkPWmxWXf3u9IH9VJH0c/IxX23bQ+eqxwYEKnmxu/PEpiXsuQ6P
xbtd7C+mzDEGViZ+6n1Vk/xeDZoR66Br0R/UYilWq69LZnDVr3LNPRJrCOfPQFn2UqSUSfAJJ4JH
0dlv9kxmaRwCDiTxxEdGCt4OduD6S3UA+by56QyVMdh+O+z72jFaaFBYrZLcVZqUxpV4GXme2GXf
WVEe4w06QXbeoVSN4brU9i8fsXZvJ/tZmFi6LJleUUpQ6TB3a4+e6PzoPNizxxOe82E/sHPLdovx
BnRq/MzYXpbzCmEaSc+fGWAoAz6atmB5+QjxK1TCl+QAxz9kU41LDV89rNuwRE9vu+QizXeVML7g
wnCFnKHyd2tfGAXYc1r+47miAgFgn+1G0ZEszdtQrV+EfZBIUGVvYSOH52w1BfkwQHbBC/6knZAS
ixrNww513PeL8oQYXiR3Pnwcf2CD5nRX07EAIJsAkLm+HKBy3QoiHJUDEDo/tAdtqTGEHHC2/G9a
fzvLRA71siUHl860mkbUhGAqdu2owHSB9vPmJBfk397il2l2Xl8Lc0eHKE1uddzqXjpL1HSkAeCZ
hZLBatdKfBmUlW9PhxISzHcWphNL2Qix4pvNwyp16UZtja9sE47OTojnjGQyhZYjeMU2hTwCoMOR
I6i47/yzpzYzTbqMG5dyW8ktC2PUBMi/DUjfDrH+ayP0ThbgqLKMDQJcSOPHTaRFTsFJ9i/0+UUq
I4jHjeL/x2iDAOhwObfBT+2UzkjNyhYdGttSaCMSKcuKnMwWTyEp2b3ae0mdSRICU6KiCIxU9wYd
+EsQsB2LWt6F+JGnfNaDO6rjhlmYDi6/oTZ1EFLYmqFclNFiDm+UZkOZ6suu1rmeQExn4gWi7a3C
AxsoAZRSRfFrVXoDetAD9PHhyyRjlDiV/DaxX+ijL7V3k3H4hwMdEk6UP7VZJFkEk0qXKgMlIDkY
fZKUSNMz/x5x6hW4IRWYbDv5b6tWJiBTopEFuTswjc+iMKOEuHh3qjJ5quOPvS2vDLFduiJlcvaM
zz/712imXhPduPhxpNnMTB4j0QW1JRgO4t3w4B7nAZB52bm7ls25j0fpiE3TUzVB4pRlK5vhx2Q/
NQ8mxnEgkV/t11XOVPpFS/8pKzhh29ffqLaEPPH+huv7mPAGKJJo+bHBAbis7lfnBpeEaKpMKt8S
xgYJ0XBeGXD5nRGPff64BzwVu+n3DqsStfcpWFKEIupLwNQDO6p/IYKqjy0ve9CcKg0DLXTTVqdg
ItzNLgk09ls0Vx/SIAMgpC8h5vBIMxsIVT+L7KFKfVHGHbzGYZDd15TRYRRB2ZVftW7sii6aSmEI
XuAkIksfL86+hhP7ZmwJRRuyCHK6O47PtKera6wfcf5qyXGoJ49L6xZpa1CdRS2rQ4M1U8XVhnq9
IPwdkcWCdoH5qJQcHgM/umebNXI7pSo/R28Q4HyqVDhyg0/k4h81iO2kzn6as1ldNjwchbIcmKWK
ZYiQNSyoCqWqizF+HxrUGjBrJo1O/7oO9/N1HEC8+BqXI7XJJ/5hF1On9gQ5YIGKMe5g/Tu0qoWF
+3JY9Al/ooTA/h2MX6sonnPnyEJLfYTVd/hr4OkStj/RGe1DOghzLRPqN6IiMshniBbN6HziFVm6
p5UodCZeJW8huNy1ZJBEuKiYohTAPU6F9LcDkoERnu8ZSK8p/EBLTNYc1Wwb9ItbOXxVsB9uNayE
1BWWUKAWL0vQbKk57kf6HyNCSsKq1Jg8BLr2R2yr4zQ3Cu9fbR5dC2rnuczJnebrFAlvC6ZGl2nm
VSeB4EsfinIqJJWJ1Mivl0a2GcklPBoa6l+Vd+voNgDRDPWLaYs9zFRf5NWWCjzzMdAyXD9iefkj
nFvYkM5TVOYM/lW2JYkFcGZXZXRYrKgqlsl3NNdZulV2iZnvDevUMKwgB7dz+/eGysZnm7VBV+c/
gAWke0X3ttEKyoTK8vhpKLFi3VtwAoZQX7x0TWGdJPjjoD5uJ/V5oR1i+6WUFOdCnTwkLK6e0x/k
NSiej3PzW2wL4A9gAJ4iW0AuEOVmMYOREdLM4OZr5lkAC48cuoLuPCbCGK8PDF8xCiyTRGPNplEu
IJYF3Pm55FxF53+PitVltekJK7lAE9M32vEoz1M29zP8yC67WBqHlQA36bSLlmBWsrOEgfC8IyGb
uxiakjqOUqVGotTvgdmV2CwqQco6V/tf5nV2OwVUDOi5bQwKsz0Q6Pr5JuCPeY01MhhOiXEFsNbm
k022F6e3041lss/GrgVpk33wn3cowMkVXBFSByctFpc7ZSBmuiJMCZhWzMr/xMdMhixHTkdlXvZ2
xE9XJnbbYhFxMHAV2zAknGoeE9v7tw2QevEBcZwS5LjEkD75fNVnZEVOsoufn9NE+4auJVdrevOi
MkJAWOTMetpNDyymWNndR/mEUYfTdvImE+pTAuuii1DXzMMsTCJjDTdpYlX7pigNRNh7kICdt7VO
4K5EfKP913PKr6rCwHkAtc+Z3UdLD1b/0ICwy9V3SPcBAPo/fcUnGhYLBegGL2lXyPdqhmUoRz2S
wQFLr8gzPhMUnJFwGpZMpUr0AQ5kcsYDq2gFMx1vWtVL/kXB3ncSPhlzqq9Dj3FQcgySIhaHHhHR
KsvadFvJ+qFvkRWxQKfqLBxQ00xlE4uOVyZT4mqAVuZ5CzpuvHasF7sbU4H4YGSffKtHulBV5wz2
VLbesrYIp/7OWIOqXBdfrDQcch/N/egCoHUEXSgFfJ6t5StY6c9YU5tcsLINCrrbCJAuyMZI8Eeb
SZw5ob8FsrXjQ8+xURr3yb0LmvnbQlCfUGbSXFNFHax1RwoxMusnt0UhmAm41yej6zxzMJ3KS+mB
dNQYn7XjhRJ09u8WCI2MtKTD8iz0AS86ry+fxBlkmjt6z7yRN6lFg4AERnooHuvO8Uf/tm5ie/81
1PDaCALAtM4NjBcYbgkjBCATxsfZKsa1ylN76bRrJCN8RgIng32NfXyakdcXnY5+A1Xw/kMk9ibD
m5vLaQylasy8LXiX665+MDWSkOg6Ebp5g9jMOJayip2j/l/mP6SozrWNjRISYGOqdunGOvT62TK5
25oHz6MkQDFckJpJvWGHK8Z0B1x7IRzPIx0fS3Y8+V6ifmF9eoQsBAeM4H6WKHxEcbHvmFUHRN66
vMBR2/Ir01gfsnymoid4tkrCrT6iWYQQFjehLEIMzw8StNzyHYDRk6QCLeSysQbBERpjWToEMjeH
YLIZ7botzcfQDtO+6+jnT0RndlZWsm8JK1zBVDPsaXORrmPQo9FJSuKayV30c6YkEL98jQKvEfgM
HT1lcaC6a9zLB3lJ/s2SygaovOYfw0c4ly9lY1QhjaS+Uk3dWQVQJCjfahezOO2dJtS72AaxW81D
N1WhU+cPO1p6cd8wfuLnlf+8Rg1w6CNrkvhd7Nkn2noEUNEzSPMoKzVbfzgPJQU5o4MoOx8DHIcI
N8G8zGFEoSV4wJTjGEVeIQ/ZDeX0MpgkaadoNf4IuLwSFSXbHx99QfwlcU4I1Ls+ygOCrXtgP8e9
2UlvW840EPxE0pSCnv+3gCCQKnQGQktudO10YIv/fjYTAvIpEV5r9hTNx8pxD5zfvg3g/cNVgxdM
DVP1FD8tAIcd1dzCVs0gaanasD+d4m7uzpYrO3+F5mOrUKH412WERHtHgVLsoIGFFsjyKKj7q2ec
v1mVW29/rkK/P8WJF2N4Q/JevgrcelZp32HpdRxDIUd6Ks6x/TMUAT2tibuik6BTfR6fKoHqEwzu
0YwlGL/Ctw+OWI2BlvNKOYLwv2+ENJ/Os/njjGg/nQmFFzLFsU+aTDHPKVHGkrzs2fzcIiCJc746
t5m+YbIdFCIa6gKsQ91NO+Oje1fcn6ToL2iK7UvKvhtnUSo7YuWASACvGH1RX0K8X+ih2YzvnZNx
uFaS43vbPkOQyRULx2JegJSkfrW0KFP+OqK9BJNrItTEnBYGAa0XgQ3UQnhGtIIFe4zK8BmUxeDR
d37Ggg8UkPRcxM6vNqWKN8cLTJqi2dzpFkdEAXQqw5Dg9EeBmz3iXvhZL1EbHwBJ36hIm9dHN2cA
6SRx3Eaa4DuBtbjNIVm8teOdQ8HsaX2Xk3jwY0QjgrVQVe9U3mWZvsOXtb+AIaBYvDB9gsndHEDE
JKUuKISyTrWPgQwlCUhjDMPWKH85zh13m3RsebXW/hpuhpJ1ka8D7Lgv/WUpUo/jLG831QmPP4hi
41elMeJgubMrW8jUgdm4EnpLNSMdGtbBFQgHFQI34lr75U4FRmvEhRkq4Tcm/B0/POWgqK6hxaV2
U0mBTnnVZ3F4Z74COz6Kg4RNp/2XdVVBodMRwxqGubZTJfP0DI70H3ewZns1PA12P9OQ+hSv81w7
rYuRDot7DFW0C0lfTNuXDSLyHIj0ouJkvSUz52dBKA+wtw2krHrIb4MMKhO5qlPGGDO3sAbKiMGq
DmwlloSCx7Jg14WM8ElDfS8eclqleiWi+sZmMGzBnq4T+IoK0/9/6hAJD1BW+rIqCrisImih+pPB
vZC0sOT4RCq/sPbbGKYbrFdlcrnmxrVHWdbaU068KKdopcGo+cfW6azTqtKwNg/qwprrm3EIMW6a
4718K+3LVxUmB+QwwGs2QopVAWOUQnBf6ckAoQL/XaLSpxnUG/VPp+oFra3dFXXeFBM7aBA32gcm
Rj+3B5XRwZZzg+zDT7XGMJsQq0lzBzVnfrcfEYvxsz1/G5UIyx7z9wWlsJRxEp0ppLWDAI+QO1fF
7FLryINdNnOOQC7sqSA2pgJqSXMDGCXhmEsPE+OAMsZXl30fBzbotHWY4RSsDwwxk6vuTxH3kU10
vSCIhmLMBsoLMrt9q71/M7v6A+bUFBL9QaVp1qQx3vaZTMnuMcEZJCwAgGvarUPOb9MOGvcmCTmo
01eMS9q50g1r1m9Ci4l/tCfgtJES0/4GZlrTM4onZzgLsBYjOeEkrmKeWvCfpDHZisjBSRmGe3kr
ZpXUQhdZQn+178jovFby4nguQPC1CeP54OLcdIlf0hhJ/I7wkSTgi6xWeDiLMCLYqxPTr37rbNSy
Bf8Pr0rsBajNN0DXx5/tdYMLe63O5xRn4FqJj0v+9p7V8hQuDALFlyl60HB/EOYYdKabo7c/jndg
1LwrmvGruLmthkH742hhrryHlXTQMwPp5hFUKWPkTWJryViqsvFvDcXiokJxrt3CzJ0LgAbnY+6y
1HL8YFDsknigDQpkKhYPxYWgx0eJmVL/KBT4tDnvJkQBXhfTK16dmXi5Xs43U7gv4/rtkWqWczNd
5oZYpJ78LfiAuYsqynyglcsK7WUDVAUoNb7NE11Sdeaf8qWJ/xp3josaLEdbr/1nQvgF/wvy/OXQ
CRT2bwy/YcRlzcbdb3aX/DaNmzWtqDJwlQnenOUcZ5CE+4r8V8MMythv2sKIk40xmrsylYsX9tFl
qTr57FX0dN7wxzGObMWET/kGm8Zmo8UpLwJ18Gqc5qD/M6n1ng+e0u/UtxvFciwsOsBI/QWmm0JY
v4zmB8hOdSJGWifux4R2FbEW5tFJ0N1mAAQNv+cbZId1e9GNYKN2DBfk8+fXLsDleiMeCRwuFb4S
xW1mRKyfmdNLBsrK4E6RcI2kqNZkwkJlCbt+skJyp9K6rmfD5A2uYCFGxOtnYSDpUXLx/aRQoOSq
tmupoR2AJ+hNrtvWrPkn1f9Dilx5cVtGcQ6QM2U7UqXcyXodxDI8xeT0LOJsA0ykhty9fEWyS0t0
LIhWbwg5WdG2bhzgiuKpY5f2MiQ3kto4YolDRhkj8V9hnJeyEXc4Y5RAozMnPPPy07pAXNQnKokn
Aeb8IsrmwyP1LR4uULxRuplo5LuQzMKAbyZR3FLH5JouGSQTIu8WvnZmTZ41IowrwMwaWROQYAZr
SxHRInuFk9OaDIkmF9y/zJnsMUaTcCUuFFpFDY5gaN13LMgzhJPOFXAi9BapiVp1o2UR4KeJCr5y
ndVymrjamQmhwsUnMfWJen1jjSnpxfv8Rup+LaE6Pr1HwjfZvrrVrMZ03Y2mpf0mgB8lWoQr6wEI
T2/2Rye0yP2rtWXXqcN8p12rEa5lew4nzgczeUSXo16948jZGl0O8aQidAkUGOhIBpkMltkWns18
OGfPm4ZadcBe8FuPYNBYGY3Dtz0+4f7kYJGk3DMrS96kTlVT5JzJm6rJ4VFyaL31w0F68dJur6EZ
OfB9a8icNc0TJ6z6JmRIjVslRL/g4yo818PrsmUKH5+Hf8vBoLEaBTPEMkuSFaB09hbPF2HbF2Pu
zv67e8uamDKrJqpZ1CeK7iEggf9xQ8z4v/6TUJNlDTX/uD7WiuZRPddVfaXHwLK/qzvbTR6opzKd
TozO9OBndvVvLxvyma3uTTBGtrXJDAnZ7Dtaa1/QntvWPHPOZOAP6f6L8xade0jfUvs6wwu7F8Jl
btOjcOAL9ysxVjEM+cDhBfUMYXTcC6vw/ZwbImDosQQL02ElSKAFbFBlc8I9xo9PaucvAMw/xvi5
12oAlcNE7+mF3gunw/FUqcy2teVY7gE/gGkZyqa3zpcsgmsO7YirNAHNyj1xkVUPasR2T6UlWjrU
ESraKEqrNx9PpBMzGE1h6U+3WTSdGd35HoZVSajH476oOQ7R2C8Luhi3aq5235mp5EAhdzvhr/6j
Em3yTAChX+It5cK+c+ILk93m7Au5EDKgFC75/YdvR73t1zwskENRJkuUkE2Knlh9LKVTXG6ofn2r
F1GV/cfMclDP4z6RnKZdug5m/n2gQXIAmzGS4AX9zPdhIn0kcVbuc9Hz3SwFYLx7SOdy+aK3d48n
NVJgWs2N7br/i/N+piooElXGESOE9oA420+zK2usB8mf7yUjjBs0d8e8MzFblMQIAbefnxtiE5cL
mEFMno2XWzml1G57ZFGrpmar67Kt57v5wPPz/Fyod1QlhuaEBaU+pgewdvZ1+37foY8jYaAQK5be
W0Z03BK0Hn9zuCXp8+z2CRQRab77QWtGcWBL3on1SqK/HjNnZxB7xFd83ZrTnjvlhzndXtEVbpLZ
5kCuSu6MJKgxZHmOdiPPqHCeppKa3mOukzm8VwxNCYEti3yndp98FGWHL/2+pk/GAIHIuEKepyMW
lmhjKtyXyITLVG07St2t4mNWnd7gm8IRPx3GgKjNbJAbipoa1P6LTplRvgIak5SXR5YrqNN0uMg5
0nTE6F2CuQPuW4LNKRngV9gEMRnU6ZsRA/ZmbZP9ShTTPUoxL4zntRNAGE/z9HoGsHYmHWgS8e9n
o4F0JpJ9fzqCOPHlj9OB72OrVQUXO3O79ZVDBVIuH36/817jvHygIxCiWeSz015oa3Su+OGq1ono
7aEK4mmiDejQ27sfeXZHOZ6TwLCO2HJmzYc3A3Ef5wVpW/YrrGSABuMADkJ3viwzv1slUz667f5k
l/oUcK9f5sFRw5QSjkNkbyYXKeKEuhzOchiytEjosAXZ/w3PVowJoJnCUJLf5mKyO52gMw9txCff
/iB4aGFXmtlgjrhM9bdmGQB2TuIGZjrdZtKC3174XG84d6ZbyloaHmF7ZYX+TjqkD8b20kUjGxcM
UV2oSuYu4ULgPtzTQbLKHLqScs33d886i75c22aJhKHXmeSQMO187lWhPiHYcMNNj91a5HgJJ3wu
TlH7ZiajzibQo9vBC0MM1Tvil1IxPT+YmYR4RHkv46RrtdMJyG1kjYTCGqrTZu2gqL4QhkyeIgAG
xzqU+Xfvs0W2fysYOTLVC/D00ZPsOHeLalzpBPn+0o6S3BZEzjCogqUkF1KoBVtjoqLA6SuEyDkP
aGuwk6VRvzB+xngJXXWMLtf7CvEy3NllLIkoMM/DiA3SjHsECSEdCSLzKBOZT/qraoI4eA1/lkCM
iFiAJFadBRoBRE23CN+gPawR8XsEcBKdYnbYQtFooKWkneBlr33dqq9sD2s18A9Ha8Bm1z126mVR
xnY7bEf9HkUggxx8qqOwbfxK6AbysVtWfdabULSIkHWE2DUAKs6KaTlCdzJxPJWdXY2EEhoUtiRs
mXaj4tMUR86cOfEMVHAsmnPtUJCnJvonj66u6mGJHzM1IVXTN7tPK0KAKqsCug3PEmakuxyFfSSz
FpP9Uu+ZV9JrV3VAV+i3xuRrNOCfdCurEYCs3YmAo2GwW1dGszUhmrjjSEzx/X7qGW+DQiNSJej5
DIpHVrrLoNJz5rLgraEoQPlpqYjL1d73ebgsj0EKJyCLD37C7oh6x2nze78AZXw3qkNM9RQ/a/Ag
xK0kKHtYy/0UKiZAzl63A+XNC3x5xqqkOiFnU8JeDNSNhdseFhLdBJ0lw2K1n26U7oLjGdgoQ3Ju
fAhMLYklZnkctv4TCo4tSGnYaor74ePdkqYSpY5hf536D2GHGQXEoFDVncbUmxZXzScjomv5Y3su
4AK2IpDOlDKX2juDR7qaoK3106ZUh1szgjVtwtvC7PXUGNn1zv1p9zjhCiBy6xQHsIOZxoNpfVZM
QVgB33pzwfJs6FxzB/JkZZyR7ZiBhzOx8DyfhzpyxqIPuGT6DtmEJUq1JXUxyemmGjIMY9yOHFKf
ImLC65sMaknGSqsd4g+5qnCQbQuFt1nPHt7mZkmGA3GzB/Ff6tP6ouKkoVqfStshOFqfChoAcvIX
q0d1eLtrd7XMJaTCVtEKoKQWjKC1sLIWBxHCvCkougJCEFsk1sCIC9EJ2xk3MlFQgRtdNSvN2q2/
Qf6yNB3TtNmoPHkzLn2/AhhJyFhzEGnT3w/jLvkh+ov0HKR5nhDOgFuRjqR/Lng4hjEk6XJmedbD
WrVY5okPC0yK/991QmRlK5Gs9uEelemvBhU+xs93ZbAn/T1u6Xcn+ELlQZmPaGpabRfHWO8gQGmz
pTKgsTjS7wqorCSW6mud7uc7pkNYpceHd3nC9r4iH/EbbOXGuE9U4A36qaFrtWGyoSKqhmmnRcQS
V8uOZw9zZQV+avdjDxiPN0pmJtF1KiGqbOrklZE36rj9HpVsZkGTZ7xVcgzHwbVXQ8z9sexQI47k
vuFnpYGRiOGBUgp83Lb85Ne2rsVzy5Pj1scLJ14TqgHtNys1xjWtp5wXDydTxJj4lCY3WAoUU3wC
tzKOTSFBcdrmzS4ATNghbxcJYNi0saqIeaJ24kI7FvmqM9KbYfZ7nlaOqxFgZN2XVyK/qpBMGIWh
ta0T7p+/7FviU9pJXrUjL936617TFYQ24L/RO6h/HsD4scUASiC3f8gUUOGn0RS8FweAfbaP5Z+w
e3KEva+NGL5+jImPQJhydbgXIZGJWdXzX8RHR/Mmudce6JvyRq4oWtEHDPyQPqMo6N7A5IT00rWm
HZ5KiAsELfnBJnO3TF4NZfL6/WZBOORl8FvH6ZUqkDSuEKkU8OqLk9xzb+qzRDHu2yWq8c2qKoe4
0Ts4Am6wnyTUAb8DHD284Y2dD0nXIInqo1YXbi2qPKe+W7AwVvYIiXBH2xpMTWOXd7TFOLC+hntK
CwoK07WsFF/BsrPjdXwIvK4PtMUQ1c7j3X8b+CTmOxxQT5dj8WHOapDLYFbuiJKtW8WDWHJWDEeM
SnIi3qa8PyXXG6dOv//InpeXG7UwaqaapdMcdxtaokcFUNvcSfVRGAYZS4usWV4Kis8a3gD1tC6B
v/Nhg1iHCkxm9EGA6+FMtYyIEUHzNr4gt5XaGHtcuKk8FF6mk7vXwqsHUqeArcGxON6wTrbIP228
pUGa8xQg4qiaAhU7Qa/ezu1VyzqwlTEb0yPgq1koZa6XiT8etqPYFjnSJNNwJKDPSI1NzmmfD9C8
SKdfw9/U9f7umdJz9RfQ4W/NsZe17Hg5UniMgAx4wADZ515cWr3EtpL1KXbQrAGg62L4o0kxUN35
4dyvqgfgt5Cg+BQci99QvT1RtxLJ3MZ9OmClyLOqZq0kqtWCDoSvBxCXGTVmHN13ajZJj0rCHALf
QNoULRwSaNqQaWl4JUhEE9MqX/v4sS9lSjNrcsQLhzeVql/KfCq7ia5igqeWT6MdGg/3RJlwcv/B
jBolGHSIzh9OH1B8FVJ/JgcA2UwOOFszjNKS8E9q6icokNB7ttbdijtnSeclQM4ByTCL44yDlReU
4Zrr0pweO9pDYOMynrHObP62sXIca7vmpW4AzstEfXw8RfuOI5KmEtCgFy4BdzRv35nPhXSJO3dr
gW241vdoRPnFAaHzq2yVPTqJmZzgpglKlX8V2wfjK6OgDgyzrtRaMzRqNiwu/NejnqJ/I6C/eOV7
u6X3fHK0+y1+/4fL7XKjzsIiLtUHjgf0RwxXIdiiHUP4d0tmh4OZiRiu0Ifw8KxdkJXhX8NRxtPD
tNgFNYjcPiwd6dL1dNJhvt5T9j+qnp/Ig0DW2Dl1BGwCQalZaqqDj/rnpPkGw7eB4osl6Gc9YpPm
93oqPBAYBJ3xNCENZWGbNw0HmY0j4+a7mNhlIYV1BliZ1wTz7pKnyeazfu6RXhp22NNhrFp5nPnD
7eQ4gfntI4s07Im3TPhqY3R6VzRuf8lP7MAfc3mLl0kH8it6ykDGrHfPHE5OfGswZDydiPx+pL6r
U9DZVFEp3GS5f0YOpG61GZp4UVkDsOATsgRrgel7GdcEPPhWXR06fTPdwOS1w+2wEXjft64kqWo/
Etp92f0G6xT39/JUsZMJkuNKaSLlbgxvDeUcwf7eZDKGvECpKnCkmOw6uzSpXaVbzvPtb5rolnUI
66fprztAeaEFTlyRdUhl7WfOZU/Sv6wZT3XExnFTWIhd7wP2DmS+z6kam09RYFs7YTYM1EXNeb8l
t39ckl7/D7nqdzndVzBkqOhbK1PPToE0XkhAeI+55guxnR0iDj+BiehukCVTUQfPJb1BwyV6Yp7t
Dj5RQwDBJoH4bw3UEmDkQBZ/zvwdDIMOgQKHsKKHKq3Lp2DevNp2K36UTtlP4FBs7qXCjQaqwEQE
rrgzoo1VkrQnWEBJZhE3Id+E0nRfw8itsn7oprWGokhAPPX7g1v8ffyeXumtUeQP40CH/Iln5wT0
FhfmyHboLfOkqNYyuYj3XpukOzFsDbB2opfJ9SzmWbkj/aiq6sB7TpFZm8VWeWzLHuqqpsY4AN4T
KhHhKe081vgin+5PSaBvioAabgJv+bQC1Z/T5mTbmynqt7TBmhAF4JLYYvSmwcUX6F+8Y6rJpSiv
IYcoFikXLApPF92p0zIvJZj7bivP51HeCHebIBDGWqypznsir1nD6WGy2mk2xoH0GuGvX1w8hujw
HOBSxAupKZxxOyfQRFAsLL35pys0lHbcLdZ2zyqeJAdCizQ8MW34Ud9nSONlp2QNTyzC0jEhE63N
7K6lLoeqD4ax5jbNy3I8hJmdUJ5B4LjFYlssdyVPcsvHVnXPt1/VQhU+lpRdR2nEJDPgzPKgGkEt
hF1GyjoaKnJAmbgAvhhWjMgWyhVuKT18fFokloov6bHJoml5iXGRrzCYaiylfgxNAVVOEa8B9+dE
7v1vLIN3IWudjWQU1L9cxyvdGDq+STkJAouIctu8RHk4OxV/qlaBYw3Z0cQrk79MlUgSGSnTyAIa
0Y4X2sEqUqndQROezdJCohNngKcPTx/OpE69yj0ynm48SVlKAKdskFwRgf7TrsQzGuvr3gEQp0jw
GuIBTR6kdNZTfRk45yzUx2c/JCXDXzI4G33FXVx5z7AUy5LI8oO1F8ly2llKtI10Jq32LgLT9OIq
H5JIU8+lGkjG1dpRdCeUU+4jNTmr4m4EvWLHmgEPK5yoBH3kPs4XaNPV6mNVDYrdbGezSnVOz3Hg
5lpu0BV/FL89T5gxauE63qYbq7bCjyMDiTBiOEgJ/sECTzJqZSB2biZD5oWpWZPsw2OO9tokoQlP
2KBSop/2WWZVx+a4j1Z3f7xPvxXIxNjLahaeTVlf5LR1PHNEXUhNyHI0IdRYnVuTUsnbXEP7Qn5f
V/1pLZI3n9/FUoPhcOzJVFB/DDbUqh4zL3p5hh94DBitx5ow56SO32+6xWkw8cFcKWF5KSTiLii8
tIhXyvKbKKyAizq4VFCQ/VxM42g7zgEo10t+Brap70WIpTLgVeWklAy0H4VFC9bOJRpQV4HsG4B6
QtElPQ+d70thVeM3eu7Hx7SRc0w/fb9qlGssR/mAO5SONIwNmWgrNLO13V2U/pLZ5kUnrPAWHR+D
4xrwtrG+hnD7iw2xDWt6Z6P1UtL4M2N8tcGW6gY+s6fUI7dNswUmlwfbEKJSDoKyHeJZJ8/mejNi
GgS49ImfhCe+4CMx6Fc3fscjuarzz2VkeB2ehTpHjzglFsjKqvRAbRV8njIst5ZDL9S4kYYthHHc
fjp+A8LyHHPAVutBF4J0Mnfv90wWbe9OW6Eu6KHwBjY7s1PLsnXOKijWV8cyrRv4ICyxRR4elGhe
oaCN/rV0oyybBjtgZYC77WiqGWskh0EwQuBXdQ6BBFUOrgdlnwEk3b0AMwNQZ5jTtLvIjHb+bfZv
1VGbX23U+sv+n6yREovwh4TNwcZ8Vgkn5CUAol1iq9d/NxapyungpjHHZG2rb4yg+/7HPjj7Uaaw
MEyDBYd97T5AlAa2rhn+xivxblv91znE/NSkesrD1VqQpI31yBIHTmB0Y867ZKJLFI4MwxxGVNFM
i+HnA4LQzC5YJzy3BlscHQ4QMY0DsyopPUlK0jkQmZiCoQ2Id6vLwIKljGrWjQGiffuUvfjgGW+Q
WAJFL/UpEa/ZINBR+HhA3HW5Xh6PIEE238QZYI8Bw16fzU7rtYaIffm3wRIXyfZ/qJiKVO2QGhke
qqWCkf9/cQ8GT+AKQy5bpCPmpH+ohEPaK/4AaNiOv/nb2FJBUtKXt4mWRMbIV1Sm1q549uqDhgqI
KsxdoO06KqkZatnSoGTDJdjR1+ddVEoJ1ZAeCsC/YlvQVmV0xiMPQm407ZEEV5QbxZxn1OYfvvPo
V2jJpr6R6u9aX4yKEY0fDwFLOE+dwJWVNQNil569Wm4l6DdDMHDQbRYuGQ+DorQZ9B7ykqGn52us
WywHyaw13aIGW/fNIpjh1Ze5M2dtzEeNJe4fLiG8SHB6PH4TIkcKnSeh2wxhx8aMyX0Zl8Z0Sst4
OqtnPV2n2bES1MzH7V1vLmuCQ5A3VpENZz67tv3kqP/SgLRDEUOcgaLjKJZz6TnYVwqb2bLoZVW8
+Zum6J3WV2Lhp2OE+FJiDnRWiM9MaQWKKOv9TKqxWYPwu99NkQOrhTYD/FDXer5I9X0C4nTFytYM
ZDnT2436aFHpE1pdtwPZSKZEcOsGSfsedpaj41pnvifaOOkiI2G4stFUCt1Yj0TsHaff5HOcAigl
te5pmr1pvqltrt1e99ThftYciaVfYaka8RyL0xBMHS6L0lFSFles7JyTn8uID1TtJ82rgdjaMZ8m
vvCe9GVD3rz1H/x8aUQ6iN4qsX++CTUiNwifZnJEYX2aRjIJGfmTjYVXR+MBZJl44A7cAMGC64dj
LZXXvki4EB1cnIBZ2v0N2TollNV2AOfPIiFqsdcKgBbt2S0eJYc5oehftkl56nICcSc3FKhazBt2
G2/LBfbHj+TVjY6sqvKOAdyHNQrmYnvHZcPgcP1gzKWQGAID7xiFxCgcOGaJyXY5LCrfyzEnxsEN
dSafhmpwjTuQZjIxSsma4i9yAFLSb+uWLfm9uT9bq1BJEd8Brmfo+ArV0XFpE5mNRqPXqhDS3Mki
/2FP19YPdaTTA3DzJQ5gMqGJgcxTHd5OI2W5OaqrOGGHnrp9hrX9H+HMx08X2D0iVjQmA8hmweMu
3VPWogUPkzUTxmq211Ehrx1vrUK5qMUq0xqU8xFITDYPbINsLDmOlxnLXL3OlH81l3XI1qHucGA4
6V6w8TyT+JfwDQoUHzFqhTLyPejaIiFhcrdEednDp5zH3XnAaZXAs75X5hzkAyy+7uM6EiTB2JFh
21/yDJ2DBxdpl4CAYmyBKruIrKqJKM34b619KMRP8cWoUV245+4qN7Z2xDAAiGjFtx7co2LRN4z4
901tV3wpHfY/ZxTy+Mq6h9BmutOrlG1LmbwTWos7vIPjnPd+pYJkpGV3Eg8B49dOMCPqVWfnGnGe
00EmC/6G2g13pc0sRcNQ/QhI/PaLPm8yQKkz9fifdNn1f7orz0/bR5owQa4svthcnTDkOferf8Cn
QoqAIZIcwDq2W+OwSpM4EMuQ0u/1KygpZ6aXxWSH9Fdyr9xTu3DIPwIyzsMBg6s+BFJ83iSNGQ4q
PccmTd/LWBtWjd1QhUavca3QUpir5x5vpMnvz4tbKFUxRKq2bEuYGnr+FFS4t9yFUWI7EZlTO2Mc
M0oNUyKqTAbQp86ouEZlW3HP9JM+Azp1mBH3uIuhT4xL7ylQHDLBncJBuAUYLcqE7hLxwGo/W7Je
w+Hl6bf+pIRSHW7I3/gMMNdhA2m1g1pytqC9X1jIAA1sTbRA+F8m9ngYrGMcCWLv7nfqmaoSPpe8
aQupyvpCfR7mpVF9qzXN0QrSBENEcQNKZjN69e5+uiHGNiUIf/PcCbc1ccQhwtlWIfmKbxcO3WOs
B/A4ixh4jlW/1PF1LuVG+kKnsXtpzAbMHTvQG1VuqJwax14QI1nutDZ86No3FU0fYEdkwd9jlEWa
Am/CeC89pMEdQ1zsNzNGoz75tcJQkWNOOT6YjTnHn+GnnXpd7FrumjA0FzAKQq3myHR7M4GWWjyt
f55XHJ65lVgai9WLTXKyO3yGKd+FQJ8s1JuY98h5XPAGZH10sp8SuFtLWdz9OBYuBGhqqWgD1vMm
1PkjJNfzjA0k2TfW0xHx47kYvnoaR75leDec9R+YwOh6jTtPcPlO5t76p820BQ+eVsPOabF9FO2O
7ek/p13JsB7gLLrqglNq6PCsa9+Z1xIVoz3R4V5TdH6fMhBKcPWPsBHuVS8wOUpZ7tEs5ulNa4YX
QRjLveokfNUGLWTo7rBH0ZrrjMcpaoZGLXF59eQdZxWofl4ljCfq8cdLIH36pIaSYVXZWdOCc5yx
lulVNecj4Qicu9rv390fNVgzQ1N1ngrTaHNyilK7EladwigCfGg1jS5C1YXwcVTPeY6z5Uz0pB6j
hKQYT2Lv7Ou/B7MqLe9jmc0j8URub9s5E79FZmcmKB4WPeshIcQXlcHqc8OE6+quQ8ljB4Ghj2tj
PNc9sRQQUZi3Gldbg0WTghGZW1d4HJ2by5SIOrIY11y0vJyh0A3+V8hkXWnzLFRavMmdl97WdrwG
Yb2hjRV5BZcYjUZgUA2H6PJocES74RlkJLSQU/3L/e0dTZX9oBFCzaMdjgU/fkM078x52hxMM2Uw
+Zl06LUdC0uXzydq73cv6hN/j1T+oMFqKfQyFWeaf8r3ffaQ15/ASUXS19+obhb4nGZyrYpuVIfA
xhw+h6FlugyXX4I4nCH7rQ+jda0ydmfGILUeLw8s2WRMqxwxmPAMuvrwu9fPyKwH9IEJ6fQBwffK
i9UpmneKXYVyqugObLVc93MknV7aDLDOTcFJqjyUGOTw7IhnwgGvT3MQkuoD/nZ6knGm5qIfUXmt
EkYv/6My5g/U1HdxKX8yUkK0ly9WTExSMrLimaAxqIru+5WyEFmfglmpFV9tOeCZq11/nBd9sKnM
yv/phg7149hW16uPtSpZd9Hq3Vu0XQzcQpsdcqncBpGRCiHNY0PO+A8rdN9Tn+uyGAulNfzbEsZK
eb3kHJj0+uQ96G5ZujSt7BKq6+nC6lcuMdxDvzAzPc5FASxdC9nIDZ7ADJDzJWBQTBU/DrmcdZyS
gMOnbzTWIB0YADBp++kYWogEB9AOKxefWIgPM3dZnTkdyV4opL5kkTE0bVyWnnWMAe0b4ULqgMU6
PTt39dK7EG862MmVyQAG3ttt3po1K0hOViR8okr47mvKblgglmScfTxA2s1Ld0fcUlajNFCh7hTJ
Aso4FbcazyBbEcIlM28dv5aYdmEYvNc08AE5Q2wcFuc011rZagOkapagk3NBNpnM4wRwFBaiPFy1
i64EAzkmMcmx/a10hFfl0+FURPClgM7uNE6hB29JsbDSyQoGlB45LkUDySknP8INfYL2tFKgC/Om
xLDYUElT70fosBPSgeb0+ywdikvAX+M0rH440dkkRbcdT3cSXnxAreO24yzpB65PQ6/R7/uhlMmv
07PonwUH9+79j+UZhhm4PTE4U7TFUPBxgPb0wAAUjAVpUbjFjmqMwA6n0/Mz6QozO+l9NKkoSpxk
lOahOGKXMm0oKRvuksdCOn/Ztlg7s/+zEDVvUTKgdhZxV75vxX9mI0hq/DFbBR4sH9aGduo4OsuY
Lt6bGWkxMXBtjB22o6ZCh0jLZ4ARHNmGnttbcAuweYqGiMdbiCdVUXV1n7zNv+N0cXr2cMIK/i1k
AmEFogVrW70W8wcHgMO0asdHULAOaukhi1KmFiSxxZd7Cp+LeWY77k5yVB9WbNtdgmMy3MtQs/hc
cdL9FwEevgtuMWAndx+HN7E+yAbBi2cVwm8C6/QoCjTYld6hZxy9Z1J+xJWCtR+virKUleq8BDAC
kfoa2WFu74Xb3H+im7MtQjY/Jo9QVd+5YHEDdJ8trKxCsigEt/1ftiGZFnQylna0RwJ7hMhzrAR9
nQZ+XdwwAsNLeLBUvbKRjuIBZumJI4Zne/dLQ8++3zDu9YIiSpmcQ+5mum5wDbIdZOtCEThiozMG
Sb7D28H7uYmfYOXOTyQZLdkuI65WD4usYrSVg9Yr43Af9ltP7T6i/ci6+J4Uv4XwwwHtV5Ck7l4C
UfFz/Lf9IEOW9pz5XnWTUqUQWoePXFPJq61Rent9oOt0irTdL+OAe19Z9Jlgx1+nTS2O7fate6dc
Mbb9d/HRDW5xRz3XuYbLHPIIPj7wXIn49/II/jQp5pr94FRbb51nYCm5kkd/UwKvHQinBnIzs46X
hkC7qOXAZvE3SU9O0HC3HfumcWotAACZ1/zA8aXPvMNfU3oJZvxMPjPkyp23p4N5yWLOqgYyhpAh
/CjeEWHMogcpLx6MleQKj63FH4zaSY32QzgpWUziqmsyKxVMel15jmQspf4rNNBEKhZ2YuYIzgvT
A9lno+g1NzjDgvpMCBUseTL863PZc8rBd2KMTL5VF7uOSbwSq27lb1+urHN8SaKL7nJWf3hb3b5x
93SzHmFvDH5/cfHdzrMxSxL+pGz9Iwz6zFSLzDYMNu3eBgNkgbDzEHodMVqyspJOworlXnknlVjM
KzBPTEQEHno7KwtKsGru5hG3FeOiAuDCQKUdo8uZb9fzU6R9CV/H7BeJR/VoykLcU2kjx2zBCXew
R0AUZZyrL3+CKcWw2JqJ3j1CMRCOsrhzVjfScK2I56Da+8pBondurvV1ooGHbal9FFExHUqxQhj3
fioDW09i0mvse5zfBSK9ySbEFiAWXZY47h3axszL2dpippcQz4sKx5ZKO5m1ZM64FzlsNjzWlUvD
NhISk9SHXv/xMTJ8uyl1e0QydUO8sJUFnCLF7FmT3mf1UvoJprTkleuWhb5R+Vma9D4Cj36HncVx
SZt6PRRqlI8jqXrv3BhVTaYHgOIZpenm2FMrc2y5WoKqCUbrc2Cgc4tz6vUtECYjIIjEY3RozOmd
IC33gYuMwGA3n1FiuYcfGGOr0lrPQM2x8qKwjDlgIbIqUwRsBQQqHvP+k779op5OP3rE3IwdWVId
i4+cj5H4Fy6L3aLTRis1mACS/j62cnmc0iXfXXQguffK4F7Jp8Q8b8C/OBLzzmwjlcUzdFNpTIF/
MbYFweXNh4mb3NiYwiEmQDZuWqxSOd05wiMmgRFaV4tcYcLfmoiBOrw9arOLLbNBw5zwednp1vw8
TcL8bkuwsmMDvtGWZorGD3G74HR53CD1VMnTM4JNDiG+0ACEbO+LRPGUlaFXusBvtq+KWm96Oe81
8p8xEd1103U/LJNAT4sTNNRK7fPpPWM4IfhNscg451NDYHD2mQsKUkvX4rotda41ysfe0G6fw5VK
fFykson26jQSRFias+tRJe4mesaOieYbA0kXJ8FrsOQZtzbZF6ni/It6uGst8HFurBAqmySZ4/uO
UZxUAJszfi+WDRVnRDRyZs1djRN3+TREl+BaFunmyiq9MYN0sj8+S/wJf2k9VeZ0jnYKAau2RxK/
3MOEI0XbTI4kcAzHIiKjglUY9N+SxKcnROHebdoH5AfT8yYuwEVHsZRY1MQh35yvtcS9ad8MiVIl
5XsgkgC8G3GxFH7M2GU4i1CbRazS5s4d8vklA4cTXbEz8WxwLJQ5gsO7xa67tHaPXJc/vsXNvveH
3DfAMS+rbbbN7eSM9drUDkhRGqzos/nB7adgid8/UzIr/JINCqn5RpZMd70sPLiClTAnvtkEE3VB
zDHVi44yKPcErgG6c/6V8ryW7VA7Vzylf6zC6+x3F63OQIpdhpNao1JD1sZhJttM+nKv5FizdMJo
QVBcfkTD0jkpWH/w6+RAsHviVSECGe4TMjcvt+TgcWaYzHT3HQpbZ6gCGAAt2sKF3/ilbpH6su7L
tK97+yEuSGk7TyyhM8TVcIgcUXEyGGRD4HFBKNz7/T2ze+pNO/8rGYAZEIEPIrBiaeQOEWkf6eKy
eQgxdT0jLCVfgOnYqQsESW3sviqtztcfFmoGyMRneLHx+MjxD8Zvc7EX1MzB9LDgDU7yBUxDxx69
ZssPxxmWAelbLYyhDoFd0K/xiERbNwziemf5CsGfle+7wf9d9t6LUoiwXTNAl7dGVMoGe+tzSIyo
B7oEw574jx2EnkHjcBq+nNmZG+tmurRZreJ7PuVOi+TpimBPd3hch36oE0vn/qrnP2YgnK65vA++
kTdMBN8ZKncG+dqnJ4/cfeWGdLBH4cn2rX/F+Np1JCTZkQUa0uuALDUDK/yEfAjbXhanNUPoQVs1
C4CJhx5F09GsFNaF+G08ed/6szYi9Q3iNbQAzuznjB1rBZXOFZvd4lopL93e7mZfVEgP2XyQCLnz
C4xOsDgOrFwNnIkkysvm5tQaIh3txxcHcHQgjBEFQiext77UxlZurhBKhABjdmVsWV01ggZnGBVs
/0A2WqroVlMsB65g7fxthr0yRdDH6mzqksWGPNolmCSBAJM1Bj4d/RfqL8vO5nAVqKFDfpuE2gC3
TD91FY9R5j8yK6VFVPk7Ix2Ld3vEZ03fPmpcpYzNchP461gqC9Ven8hvTCUlLHUi/1K0Rzp257pv
dUvm4ST9mcKtKLr0htHT7ZhfdoOs2MbyEk7V0ANYg1jYlKJ+WQBOJu+EkipUlM2wGcfeX1jwxZff
hNt86qxlFeoIT9sNSj0yTmftykQYFOljEFb+nQR4fUwdVOXGEK0g7Mv4lc7icZnHMkOv3IUVE8nl
yltvkO1x3EGub6MtPsmJo2PIlSuCG45YO9GeitaRy3EqIpKZ1D2asNOYuNtgQCQJQTDmhw8cg8yQ
uPPnNHdjBVqmECg1o4amVEz6IPmSck0LpLYHQ9vtBWDQ6Y6syWHLyKYhSQSciANT2KA20r7aIkU9
AyqR3CbiFBPVBovSXDlWV2qiEtZVMI4OskpT/GYLNo2ikIgb7Q4sA1ARCReAt9sUpTDut6SrWeRf
aokXR7SYCjOmAg9eZ/UAAiAkXbRVBESLj+lt6wzBBB5ESqwQF2oBUQ+gVhLNoSq7mMZ1TPeJvHbm
xbeBkyhRNcMVAFeTt00mMmImjD3pwdNqyLLd5E3rXgl/ggpoaEmI1G+vmSPO1fetviMWM03zWcDJ
FB1k2Z5GH3Wr2XCVMBcb0FQIJ2aJUYDpyimLYjQLafk5C9tn849aduoB8NYrQDa4tX6SFOldmaDy
oDyILCNQvWATy6WmxmHxw5FGvCk9fmOO1kjVAKttZDHJsfWoZtnPgfHYGxYlMFoo4aeA7lYvwIuo
m6dQ1c/ssVBo+J2+eEPVZzJYp+meuutUS9IwQ5Wh/o2mz+nvJuqlfHnXDhcIfKI+moAlJQlskf7R
yID3kNf3eZTQ+UDeGpMAUz74WUh2AZacFG19bI0cOKDSe0wYj20WmjOad/iC8wBlPw4UfY27auAy
cb9B5nIyQrihitZ9fO/mCe+3Rxya+K1LwfAYshc8eanMANnFozLLgGwN5+LDXGs8NPPU39/Di8Ii
CM+gwWi5vhnmVkB962/WJxj8HJDARN0PpPD4YEy/C9SikCTucSTcomRT/HoGGkZyQIxr+qFll6LW
F4gagPkU9Ihc3k2pNnsVfNAHkIipu0AFZZ1AM8Wj8yXvNtLJc55jWVe0KW7hJd9KClaFUeAIwzDG
u9uZcGMUczRdMSKwgrDTLTlTmG/rAnDJbGc7BU8T/1YdzwiH9a42f/ed0b9JWwpPQTcFxjXuT0pk
PWtcxc+/RPQVNvGcTE/NBrKaPOwalgXiXtBX8fL3MT/rJ9nQVy4VRdKDYlpD3M64dwssaCsuP/mb
R+Cd8yD/yNuhIkUvvaxCamTlnMX3kFJ6YZDOfQ0U48L9PKM8Ky1+HJTVKNL9NFDRTtvKHUuz60k2
+i0tSOQ2j7m1Y8nISJwBoA0ZPU5qqdCtipNe11p50SEX8G27dFoIZGPofSChF77VN+bLj4fxCn8x
YRBnhb3mLW2UDgtn+2T5KBVziLZHhE4oLDwIbn3VVupvvXeGvSwbZi9qhjiJ4EQ+TTotaOcmCuRV
B5nzB6f2Ej3pC2caCWbqdYxpk3QwKfFIEa7180QmpYna3UtacMTEPEL9IZQW5VO6XS2AmL6bZUUS
JlVLYFRB0cG2eaAuMHDsb1taWcXGoJxhFWNymbW3r3LlexfJw/KYdrVsTMYd2Y0sDKDHnnUx37U9
lSwf5wCpmvR9PL6Sma/AVwCX4EDP8S2sFs6UK0t+5W3Mc432UnKGlM+uVV6beFq4LrSzR35U+hOW
iU3wurLC7I6Bb4uybpugQ4d8Zwmxd1GTSD/zu/F4A9m57h2rzqY8KjcE1O2GaH0X2zZu/RD58E3w
JCFsA4zRmscy6BDyFs7NTAUWri6hiONDjYkQIXcDd0NGksBJrNtwd1W2/tzdjSyg+MLocOm0rSt0
mt4LIASaLZrBcesOBw2D7JOcLpkGivM5RpgWKaMTR8orDX8S6qOolFfNe3mA0RHtvrVrs5zUOY0t
dvUAzh83nAFwjyUvi8a+5gj7SPQxJysEG7lDZ9ZMYvI2FqbuBs1gjUg6AGtxudY+kjlGeEkZ8FWW
qDxgkOxlx2O6yElVl4hT6XSqh4FVGkjXFVOFGECBDIUXsiEZCTcDZOkJ2EZg9ZZCsVemENxirTKK
Dt0NM317mGcumt1LbwqVHwH6jv5hrTzdz4OP0BeNyMfShNCD3f7IM9ztuGQU53MWQ6ZwbwwWCu7t
sCFGSKRXpAUmPEFGYPlwA24MNCEw/xMpCFqAKyLWJ72toItgwmr38LdDfZIcp/ufPvHHu2ULN0WR
JCpi9JVFIN0xdL+PcaFYJ8X4K+8FuUjY7Qpz9RPGO33UHSa84yH9hAUnB7xrfJoLA+8RMVrjg7ta
YKoq7GCt4ei+DzqPkmflKJEF5g1XA5QZc31PJgRDWEDFNrmQMxgl6Kjc+KV+uXjDK76ksRADuorz
iai8BVuIe24FpLpHvfPi7bcFxLLhwcXNncR2BG79aNqT9WeVrBZECPTMEMiQWmyTJ8nCS2IDOhjS
DJj5nqfWgirszrUFHNW+7oE/tCgyxN2vyZuV/g/Mt5KDywK9XCzInprH/m9NOIuLzqrkdN/woAZ2
dYCAfLR1kpfM3MqWhH4z67bSTZ0KxEEWzF+YAADZo0ggq33bbGt/LF3Q7YcqGnfH4LMH2Vpduf+y
Qk/uUGZqHHbR/oXrRkM0zvDspasQbQR7jGqNISbPq7kt2NYahgyl1tGCUejwYF5cyKJlBw4d6a3a
fEYkoiRLCyJV91E6d0n6DyuU+wb8vWpoYWgti57FiTl9NpFun1pn8sNCZPjlC4Ct4oAmWzyhJTaB
yizGWExJBsLRhWHsg0h4ngU2KQ2ebby1vkuU9H1dolmCJ6oLHDPsmbYVn3JI48dszGRW8VM5BPxG
q07LimQBS183/gGg+9ABM/mJ68CRexeAjdQsDlH1djRVuyRpiVJ29AcJLP55avpoYT/dDc5GrsaM
tk0hmLuA++XX5oM4Dv8rXrDHJqA72ezBgGd7hUruGGu42aMfylIomE4+wYVH3Bq98Zf+XL0g8vja
KQH520OzPBs2kC0/I7r1XlOZD3cMNzNcIkmV3E1U2ga9dP+/Z1ihnqmyKit9nLvbjuvFtR7FYRlp
+j6zFEq/S/NMdOmO75dh2/B7PdDZN7re84iIMv3xZ6eVe0KvqqqpIPJkb/nmH+gnZ1T6srHjPwZT
454a4BKUTxPUK8hJjd0V6ISV45JsAmB6k4kpqnG+JD1ds4CNt3R74l6aE2mS5qFKN4GAdkfmrhBR
AZWaYw0kgiNLwiDGpWb+nRE74RNHJU1eLB8lfbV6X3QslO7MoMKNxRKHF96iYes7FslDWySKax/2
ADUAswfWBypTsxo+ljlLPh/Kzh+v1pUCdgQrLVhKt4dZgObZ4pKKfbafNUUvf2wa63UcyHEx+aiB
b+qwYXboZ91F87W2r+c6vdxZ7BRjE1Rcd+UVVhjdiko1drinbeTSTJu89ZswpZ/zC+4+h+fiIyj7
5bEkHwL9shpfDlqCPMhINKbMjszXh8gEvhuIE80qDc9Rl1mIXyyixpyTgHH3NmkN3klvE6/FJhIm
jfD/7Kzi94fbv5ApJ0hr7kmgSYXxkD4H2j1kDpzIRi9DiBbYNW1VtvPdx66n/VZyRn4DQOsi8hub
vHLiDKJuF3L+AtlksHpfDGg505yU+BJZVFz+Zt/mjWWPNsbbPuGjAl1CunkzvmscPwY+UdORH/mc
6RiIMKZlNd02/I3auPAkM0U/Nfbnaqn19qFHwG2NtSsLIuQ9qqnjzN1zjRec+WSdmoNFUdWqR1ez
NEvIgwMaZmqJnxMUQ8Dwutnk9hmEgLgvra/DVNSGSx/Hw0sbF+0kBG4Cg6ZbC14G9Dw7esrIqPrX
sXWx+ceqHA12TGJ5U2XYvHaEpra2BvdnvhIGn2+fhDbufpi6UYUzoI50DzMwDrJDxOjGMnluunXi
bmSP4zWFVvpzEIYNsIBvh230nlHhLBFW6qt3llOKLq5sKMYOqlpApzx/kQft6uY63Pmyr1CRO9sM
eGdyMvsnEcx83c3THiOCuGVfRUwWjj37E+LMIPhsdnJAuNyyMa13XA/X04QYvTg94E6vS7XRUqYV
TYUu7C0WOudis0KLv321SFDyjrNKJxRbsY2Jj0EvUhq++uehH0aYeCMa0Um9SfW7hnlhMp+Q/pe9
IyAMgODXL/LXJ8nXY6zAHYFaZSzkmk1gB2dE8c3de4FFYzGeYwneHcB7g7hnbJbNfX+gf9VLOSw6
b5CUtetEYcnsaGX44CWh2+jYJ2psYeKorq/ILBdJV0DNJZ8Cm6rlQtemM0pjDVTJlxwcIP3Zz8C4
dBhExSmhNL5jKfycJbwzPzQcGnkGAM3v5vG3J6Fx5XplB4VdUZU9H3Wm2xy6a5uFSE0BM0/PEy6Z
ech69ZGF70/5tIUezG3P8NNHekQ1wMyLHM8JEsAWUnI/Rrrpi8Pd11zdXnvkcyl3Q8Am2EM0OroA
h/SF+8pvMhpot6bECMbdfm7X4jdRyAqs+FWo5pgxE3CilclBP1WTL1bXn9PhuzPsd8MuxkZLGKfX
BH1funyHj1basYF5LMxNBxKKqHKIpnsTUoab98lYNBovlnZw+6ADVWA3P6d8jN33eyRKlWX3K+s/
mIWYCNyrgIY/LXKVNn1G9NIJ2+ifvfJ+MJlSW5gSGDJaet4kH1TtBB1FTaciMy665GSj24S4PyOv
XUxKa1I/UJ/oPH08lP09QI9uhhDoeCRaP8mMKlh26XoqwunmmJrVQzYAC49ur0n0mshj9M2p84Ys
78qpbcHVXcoHPQfFdxaA9z56pnjGQ80rpN2r/w14NMXNT95zgzidfOyiT2ne7SlD2Ev6V1nXX87y
965hPTbJ6azmbdP0nQ5fmV8NqBQZZ1l87INSAXiXHJEHnYeWQfC3S/1O8AqjE/wKNDEw2oKofdvR
LVOS9zgpBM1gz1ODMIQtoAyf236z/TXQa4GNIirOYOfZntAgaYV8TTYbVFd5VJyQAZQmwAhETsOs
qhJ+Dg8pIHLeBoXsA0qO1/ZKTtIjT1fvQzTXihT/3o9YNP0uwurAw/SKgqt94CVJwn9JMDtLfqGa
0M7c5o2LpB393S60S6eKYLz2Mr96AESmM2zACJRHAEZMidwnvUkQzJDyXBrNsdJ02h4X7I1risEX
5KWtYGRDNZO0d/NtR7i/fOKoY9uP4UuYbseSDdEX3IS7+gsQRReA9bnCQ0W5mDNeIV0uIVUwY324
9uhFyh6UO0ILpGt7+pJqPhev0MMiO5uhUv/E2X1O9SuixZp8MeDp2zlULLwPrOVkZ5e/KLCphwYO
ylWqgKKSS3aiwzUwZgLbQwCZAzcjxbzufHzWGP9bGyAGjiG6Rv2UBVX/sz4XAcVr4HWUhWFVUZ0Q
i0JFFKVNhPTyqgObeq5KHa9PzUP/hkaKuIVqvL/sNkuC1e0fSIQxg0uUP8nZFtKFdmImZ3AmBA4L
iFaKN9/UFuConYPzJI7XVIVX3g3Kz7S12C6CWcOBgsIFfmrx5GPjnTqeyBqT0s+ap3YLpqrO9gT8
9k5+Hjt7CDulI4K+R5QgB2b5Y6JwcBaGjgk7XZceRg0oyBHSHWws99+lyBx21+llcPs7QHcvFoNF
Sxjkjp8um8lwgNcXpkh2wHDO2HLlzY0s/K7k9cQeSN58I5ruiRWf/XHA4Pxn/tmQ10BT/lHy2X5c
bFtvSjYmyZMlThjNx/MieNg/LoqjTiI8KZALiE6vDFE2y1yTxmf8h4cASn8yvBQPJWogoUq4AiX5
CCt4mEMQtteHmQxi0S7TPvLvYbp4cq8eqxmeKngLEJpvX6ACUj3ddAywmmc7/3drrWu6pfCpZHk4
52ICTTf+lxATm/Q0bEBG0hiNjHG7SwSZ0Tp12rLTM7vjjHnFwijnq574Owg3cvZbmJzU6nYmEtmp
zM2syJ1f/ZRWFOJ8SyEyHTIDVWRjpDaPGA4XvZn5wfB7QmrqDTMwHxQIMruWwf+gQp79GEM3iT+o
MdWXYIbyS3lVZf/5VZIJw4U2YlDFAFqRiyJeEX+CCuqIOQc5F//Bbi6pfgrOHRRSe5iqJ3aXsuz3
2BJVqUQ2RfhoPMriGjkuu9j943vYraJ75Y8GcIw2Efc5gV2tZMDk+RV4VlA3r9S5pYN/czxMI1E+
jo/Sslyka3XCkdQoTscy/wmnNfXT6J9W44jVcadhCZkHKpKKUlRbJVKnKT5DEp/fwjuBq473wzYM
K4+cHBXAtZeZ6E1SV/iftDdR+7DJSbwR3GYoCOsWDXRKy+iifzP/paozv/9xzcdUJ+n/aejmEDJm
yke4kcNFXILvphqrGvCfeL4npxNy78aAfohpsZOCPC3EIjE4WgwgDiyRiwIJp3qr6dYXwcQ0X7zF
5XA/BGmikHTRysuF0AAp/3sQuv4kTcLAqlxFa5dnK0+VCKTS6M0xjt9TNrPPPSAcxNYzbqUuHlVm
0+RbpYP61NA/ykAD/4thREYKl1mzT8SCcVGNqDQ0BJNh342OZ/Lvxxw2LvfV/IADrotzqtZM51wb
lW7bGchSumL1u6G0QsrqSYTaEZ0hL53faSSdYaOHjaviRLND6t6AQCjfPiRKRQ0SLn7yqbO429qv
PigDpaBgFXPItPnNqtjvxz1ut707+kBAR6LOTh4KwSJC3TmJmkmKL6ipdivGIF5WHNp87fI43/oJ
7X1ySk/O75FjKVJZA6pdCMGz8jNFs/mTqxppusyAuj5TsxeJAADmYuMgcQCYche7c/oDw3CuI/3z
kO/MIG2i6UzWKmB8aCrq9GZ21+JvjB2tVJ++EXKerd/YJRKnpaFywgP3nR6pSWcOJwk9OpVqJsAl
DS3Yt7wXLwE3SunaoV2zNN9LrMg7dOWAs6dFBaJ/XXsZSFaEQSDJVcyOdnbajA6ZJcefMo4JKL6U
wKcwEanu6zEtFn9cIZ1R2BzPp3t41tMLEGnwr+H2lCC0kpNimElQq1VklsPpKP6kGqonzTgF89sx
JivdVYq1baSYKYuHQIRim/hNbSXSLpl0JLbf0QEghQ2w0D/1/5DfPgt/GuIwyAx27NUT+nc74KP4
762yrqCvr+8rg1KbZ5o7wrlhpmyNe1kAHZxQezU2ITEFZpLPna+y+apHoHrQU0iX8YBAwD7+j0pm
ycagxndFs/fzk/d+S4BLXV3U+17jms2iyYQ0d6WS0QU/c5/OtnPGCWWowXM359PCDaRJNkXFLXUU
vZwPty35Tf3ZMhr4jVRX9AzfFF+/chvegj1anRcHw8vOW0Z8ZnorZGWKLAKPKIeR00HdTdS6PRwY
0mQrlkGMLPigeFKzcfYVXa1Gma2gOBxbfgzmBr4845S7/3K086E5WraKxrGRrCY0hFHPAS19UbeE
hlQkfbiq3Z9C8CKO/y7iyNWYRIVHblFyBRlGQ0M00uBQXpY5E0cxGP0OG2afFPbn0N6u4yFvOrVj
vC0enDKt60KmjbgfELnH7GAsgR4OFEQmbJI/YQlAJY93x1MfXyCUzUJ9O7HQYenTGI6pEP65y+ws
WXiIuHL6QkC4awnwVS7WVhtyzqA9ZyKpia/aNR65xlOWy0pkLYb32W6+3pufaArdqzWeYUZ42bBx
bbb5265mdUriVbMXrePiK/dPeIzbCtx0uncE1gjUIPCj2LbOEazzUzFYs2y8U1FiOJeVh/V3pCYk
yf7LxcUcBD3BL+HDeWal+iOJMGAVY6wXYJaMB40RB/hzxkJPLJrQPR9/E7nLxBuBT2MSoWZTrmOZ
FsqYLDQyu9TwHQ7RCUHgao/UCX4+X+ZiMArR+4Os0rjHTd0hnmUgS+/omrwqCel0Hru8rLFhYJBB
oSz0PhQtK65qDOZ4/qzCl5Y3+cMtSkHJ4yXGS91ewe2iUQdENBPRTuzIDScWmM/4jtUt6QLg2QCs
MM/j6T0k8fAOx5fDystafuKkkj1su4t9iukqQbLIlwDXOPenV9JBm0/HHcAIOn/hxyeaxZG8NVbH
nKXWOVNpEL7N+7pFgqX/Z/U5SYo9MlF+VLgljbHRxQvlkZrKLAGF+XzV++a5tgzPDIHeBDW90/IL
Ol4YLANlmx3WPtA2u2GajuTD0O39YBrEg/RrlzV9eaKer6ufFuOp0YVtSTiGqsRKLZW5rhPAfmRz
I7FxRB0fsbj76G6Wjx4kSRxONhQJVnclLt1XI9gzVPFh04PBB2jmaCggUezwYGgVlFZrAFK6dqta
OPXleoZQKPqKWj1Y5d6PhpUALeOOvBrwkIjsZKaib7yApNt6VAo8ha4trNx3R+yr3nNuA/JvVvnU
+j4ZvGHV57IP1RUpuBB32ml/jD6eLF88tlIjq9o9ibEUuw85JuHcOMjwkjcQQFu2SVmLQBF5hsjZ
PGgp+b/OxD6HOmMb/I26ZBEfhU8Psr3X9xaIVvZGnFxuUaniWvnoLnrBBvcxSvliAH5/Hi3mTewQ
P442Dano+2awWbAYHBM3Tslartm+AHvP2UT/LUp1kb4jAe+hflbq4TBSP7BD6rEOxnti1gkClPk+
AknJKpf/wvvhwVFovYda1jvpYxOgm0i7WNcILnSUBlSfW1wQ8lmVdduWoJ+I/Z/fTG5zAcBEjEMw
xBn9WTj1KxXNSr1OdDpD9btzo7JWm10VoZx/M+v3k0gZWETW49Auklb4pCOFOXa4zPVcqofqN0Zi
xsYpwQ8ngD3OlmAvdXg3JN16xAE2Qdf047msXRhrkjpiCrENYiZRHF8dB1c/+mN0z3H71Wz8XCcE
uUMNhuBQ4YPVcBlI+pUUNGeq9hmxPXnSrFu4XKz5aOK+y7gA06/PBtAYRJOQsuHiH+XWMztQmQqK
TyFkIgxj6ZBpliSpXmSXCY0ntYElhfTzlcnW1q0P7HCMI6D6tqxehNgb+VCZa9HN1yDgzyBkSEQU
0lzT6SENMRAcxqJdOISALxv1/65/Mel/VIcyheOlZrpvlPl6VTLgjHs+TEcA+TYMHLa5g4bIDiby
aDqyqv/Au9j1WLyms85yF+gtICoUpvejozLGykqtdxKoeQ7ipF1RN4OQyFprdlyYhN9jnCsG/wgc
fuqFH1nM5vwIvxmjaZ0ZZEL12X69HnmKbMb2K1jv+TzPUAbdRTEhdcgql3kYlA9yWzf6sY+77PJo
V+TXcfZIm03uDHaBfmPUBb1DyCz+nbGPwyYxRU+mk9nkWP9W3zlNgVHCd6HH9YUxLj1mPjkf1wT1
D+71tZ2Sbs9joIcOXBZtpkd2RLR/VJIUTTnpYwUdoZLrpaSPT7ZBSr8D7Ig+ky9lscZf7WT44gme
mRi5P2ePSW1VQIPLxz1SaH2Csyy/oNbtYWvsy2seKmUYYrlA9IX24c5cnMDiaOyUI73gpxqfGbNN
mSv7k+bLdC9u7W8iyhhHNew5QoUWKKojcdVeRdd681YvrhH+IZwskoQktHXbJuqN6uT4T8hCtJ4S
8IVPEL1gIHvVJCl9K9W7vSiuBydAGzdQBfK2KMpCEL44/zruQcAnYwCAHFxEs/2u7ZfLG3MAJk7y
Ss+lUM3LU3h76DtmI+EtVhe2tSKfVfvIGCNg0loxnK8piS66hl92iEaSAUgNU9ymOlvBs0uFayOT
H8izzzy9iFLiEqEmcvXbLsdfTXUKgCiH4lA/0NYrbpJdigND5/KIRe9em7OanxTqcEtN/zVfgyKO
GllYXKGZYIi3UvyfzadjayXf2XmI7ry2WpYSPUf+9PLjjyZp/Vpo1H8tpcsgYKDd2nZBIHy/28kb
oNOILf2jVyBSHmDhHAokU46BloP9Ppr7FPg2KRiLMcn1w34KMRM0peSGBMIJSQpPPulANNtS0Vsm
7dYUXPpXTSzVfF30Q3m/2gbn3CznFGe6U6iDYJl4uAh1z4OHSDSw2/iQESXd49iHP4KR6KAZ+xCt
XSzD8ZEs6cH/RRFkMRDxM1oVw6DDKLmBjYFvKwDSJWrEv6UJytlL0jSRa8EAdyevRpPeB/f7bZHj
GlEN8SvwTme8CtIdw09oZ8ASoIdjyTwrDPUbt5RbryDdYh0TF0UnoHVpCHoFZYtRIAJFARa7ZJhT
NDb9j+l9ZXZwBo9uwYzsAaCFDsE3Rh7vDiQ5LiaQVrSeNZ0XTtelTUUZUdYknNO2NktkiwQA1X5l
mthhPFtWUFzDCrByg2Cr7jTtaE3/dkh2Vz4HaM2jZ50huewxxzE121w9jbESnV4+JlWfKxuvdRfv
/Y7nBxIg8Fi6/tlvSBObwFKW0VYmZQQrqnVdOZpMFl3yIMXM4O2kySIqOt7Bml3op0P//CPpzMUI
a0VzKp2Hoi7axhvvEmbGjBHR5cTQEkRehQKtvo3wg9WkORfvPPgIodTH6NtikbizMDZqFQE2IZe1
+LNE//MVPtyOyxOj+qxsXRoeSx9jraJBSBjPkD8UbfThkqgEgNKpV5Db5hHVq8iISNKzpfECD1fw
l0kcSaJkhJI+7iQJ0m/fu9zzwrFET+3OaPuXemqfI962F/5XsfnVWFEW3DoZs1UhUotPMwFQYI43
XNaii9fhbGXoIqcDtEdeJHquZacH5S7r/OEVG45Cr+G+P9uzOmE/6robRFFhf1zUn8yxdwxsQssh
c6EDsqNVzMkCtHY1vFOlx71JxHpNo0L4crxAxvO/iMnljXM2KTG/GIrQJoTAmgU9GnFvR5UFKAq1
PIGS8jBC7XVjxuR8d/GiJuJmrRmWmuUyJCcaGuY5xcPuQN3RA26rvbLLn84iTf9h2A1jURnxT2Vm
isAfAnuXUSVNqE5FqLrTThgjO0qQXiV3svH7CxVirEc7L3e3oHxqR6bMw6MnI5iNGIn/y6fTN1Fw
iQzSMmYy99qcA/st3lTB/+7X/9DA24IPcD2bIfNEYrN/zpshNkzHq0ab8cTIdPW3Pfosd1gHIYSn
+74vSKBGUyMZND1Ujo8cU62azor6siOp4e76UNiCwI+FOMwS/JJlcZKSewtly/r6eU2WgLanXRyw
L+y8j4/8roRCz3VCUSCU+M0G4yHuiCPD99vsXtCrLFqJQ1nZtQuzMKxiq+ElQGaOQtGo5YhOX81P
FdLOcsC8Gw2aN0BV1uGzylmQdO8q2OPf3dPtXO4zTeq0J74cUkzR13nm9MGaUF72e0VbElD2Tu2Z
+OjSyKZWYvvReKuhE9XHJhSesKfloyFvf28rhnAdxdoZVbcfgsNKAvtOWiOcUBUXRc9cuEZNQsbT
onS8krK4E1YDdsJE8lW4kTKpG3UHKjNDRJB4dyRe5PWdf9KXXX245kX0btYjbY66H0paUJxHXc6H
lCI+iSm5mHUS9c69v9avsozxb/YvBAwsrP/sz2MjplYbQnrAX/rgU8hxyDVLFjm5W3Scx4m5awyd
cvkTUai7ez4DKhZ4e1l/gtFvJ00mtvjB6+D2XHHtqISyDk9Y4E60VvN5sSofy6fNGahynEb9QhNM
UB/cy4nYdUS8cWeoK8zOAQQqQ2eRo2uDht+MCoQdHnpanj2vN6WDiqhiv6NBhhfomzgyfQSxIvm3
MMdpzK95/BihvGC0k2h9BcdzzAJvSf5HMZLXlCVmd/uhcgFF7I8OAIMuTc5QS4QP/uH4wTgCq+T2
f6BdEoBvW6gW+pMdYgqVAlfT/NzkWhKk9/Y39YtT4dt2FrKrptniNZDCsOElavw0llvQrFIdAsVl
o4iPAIqaRyrzOeuZQjLnTZUrNvXpzkyGcYps89wFEgU8b3ciM2k4SBq7NQpR7+rU7Gkh0Jnn54Z0
Tr45S6irmeTFo6QD9m595NIJhN5MQXQuJKEVucIuBnxf5oX9Ih0KjzGtPXlNGOUaeJ6qrIPBSqDo
9e8yXb9zAsk5GdpXVp2CLFtRHh76rMCS/sTsmt8t1PXYpKQr5/qQq6Y4TD3j5IX7n57qDTog4tAW
BUMsxtZkdUGtrObbuUGdCcE0szvs5maz22HogGu4nFNVpLoxzc7b307n2sb2UphqHWPctOPGrkk3
ygHlsMXYKhbWvEQwuD6ooQIQuDfgnRyUOYcHWBzKGna0IAPxm3GRS6/ef1CyM5cjz3zZJmgqxRkK
+zAePlX+30jFJzpsPkStJvkMp/8y1ky0x6TFlUS5fdL6beozYybMxUDT5KWmZXkDy7kkHwEOqIzr
OY5s6+2XsE6dOTMAeHB79PN153yfvxb2x/DAd8nov9/1V4c6KO6IMidPtKVNItnkqks1MwocnadH
ptggUyDAo2oQjjpYdULBL1tgEcivPwUhRWu6lU3lS4kHay1yvbCdBrxIMraHHgvmQqPoTD32aFd6
3dAQPiG4u3FGdhQz+HILducd8xAjSn9ZyClmNRetSaq2NPSDBbcOeiXJcu4vYrW9KWUolWzqUHqN
pAg1SR2wRRlZOEr7Y03hLtfCJHJNL4isrETBXsvsxD6k1MYCN5Yhe78B4XNoEL3rY2ynJb7SkOFJ
EDQkK6iCJQtitQpug0bMh0MyOMvP7iGHS02Jbkgs/xOiwAje57J+NFfX5meaQzQgfXUmFHI8FHuL
JO1qkz1h7mnVT58SpaUwsAh8DGMPW6wGb5Nc/n55LviXolufVP6MYgdhRcTN8r6YLjOibDh9osEb
W1HyUqe5eUDdq7h/7OjvZp9BvlbRXhRqqvW3YjkxV1ybfDr8GwWgPPmzDGzblRjXju9eGTW/M+2l
too4nPoNqykdiRAzBqMQfbxjw6YHg5CShHr2ZVq1m3sFUNheulIA6UR+451eFSuZ+5rGGHkOV3WZ
tDpbC2zWmPPtAF6v+HTB7PiOWL3NvB+NdNrshd1pNVo07455SGmjxmsUgKIuCyLiOxk0h+2PRbgn
woAP0z2K16okCAdG8OUAtx4lVdvxHw6CfDilXgfXdZDnx0em0EK5hYmsmKJJRVg7YtE+SkVdOG7z
cfbIeEFJogexq1Hc100gTu/IvcVjUphVek87NdmnKFzd5ghA3km9h1GQDQLgFU1KEcLgW/EC+Pwy
NZgYsut8lrInta0BYI8lYjTBPRQGV/A0SLXQM1EYm5mFXNgqmy/NH88y3dennKsXJLskLYzoS4sB
w2GsyGBK5BEqT80MqyZPL5OH7mKZFysKWZDpzBk5U0eGm5N4waMAoJB42MV8p8WEwduxuPddFK1/
vuXUqVbsB5CnQqdVlKz4jQ+jEz5cMjjmM/yddM6zc2Znd12oHW+gagjoeysYjaTJsfSbgqJs3s9T
2/pG8yaodHj5bbLB8BFXaHxpF0/+eUbaiKu9eaTd2wvKARPZmjwDhz9EI9kuJ+QOgW2/v2kIdBQo
93S3SGDmHkEvKUPwN1EbC9vbXLYosV4OidygLjy6t4CylkYd//B/+31z2tLhUVhZnSNzWOpsm9Th
sSbzgZkUBVlDqt/rlGHpukoKxfzYRF+2j3PeB+0T7Rgpk+NFz7urqNkfy05oDUH0uAEU7uZAwzqt
MTpNJcB39hOf3DglRUAZulGFOe7Iey75salFm2/5yLx1pZT/ggUVaJSoexi+/f50LIZeMgGSooPe
WSs9IDHqyEfEDiMi42spTHdLEwphr7by9ip08vHWsJ+dMOP8aeZ9THwJy2ybZGDjJZqMB+7MjgoQ
L5JCajG6Z99rAD0SrDCRfJr7URlOSz2hXBN9k+1OHobDQMg2CmD4y87VD8x9G2Ob5C6mQ8R80y5Y
BWAsasezP3CBa6AgJJeLyQ7XbpPtvVsqPYHGFvjHALa69JWnYuQGinwdWopIkSFxz9re8vXBqD6I
BQZHkyTYSZqwYqcfvY18Y3i+aJj9H15zS5IaUXlq+hhwe1zAHSYtqvd7qRqopHl76dHh+gCXj05H
QxoSkv0wPxUUC3i4zbslQmoyZaAXoaTYortrFX0wfeuI8iztZf/TRWQfWYVwXDZb2iluIKFBBOby
50A29M9WAsSc4rJHyDPJxJXK0E34i4YLxOmTHV+JizhfeGVw8nnIgQVThYrA1le08tYCUJE6G7Dm
I1LTisP8TQkuAq6a9vKQzOKD/ZTZsBFlmSBTFvf1ELO9YekcZ5nbU1bxdipVvoBeTXmPg+fUgjq0
Z1YHXt3rBoGqrlbTjNux0Scy6s98iLtfSlN3yPLtNXuNSVuK94/tWzIuLPd8R+b6dB749Bpkl5+p
du1vOX7R6Eyjjo93E3Bj2TZqxuvxLeJpmgwn8hG9t8GOZDNoC8RXOGl0jNT1y1iiQ3H5pOy5Ag6g
0MDPdw0V7RFiWSnRFvk+62+Y1EBmt2WA0qJ9Uf9A8dxpqNIvxpWej2/OUosj7Y1XtaFAIw9rZ1Xp
/OfSSmN0WLo6LcHSrTexDfk1Rix+m+iZE7OywPm0xly4Fk3sNtlEFR1kYIStvfUPTrsCPXNch0dt
3CW8FT8gdW7el5qbc6gp0uLf+DihjEWeb95h2zg2GIpB6zeoaEBmwGECpfJoO52iaBX4VkE6ZYGS
NOv5+59wC5PEHju/tTcjyv99Oljo2fS0Gf3YlVNENFO2tWwwNBuGiDJfEG6afkdnaS/etwX2VY1k
+GD+rDa161GQqUFDat3K3ISskZiKykcIv5td63Ue1ckOxobjDB4tbNkHNLHQaTQsFZ7DL5ugIB+T
0R8cXkJSgiZffUOzMR0zDzURDcuxV0O6yPziGqUle3pXkKfTrYefBDdN5M1z52/zgwp0/jXCY02k
Sz3u4B87Dsra8pueAQetAQFtLAFfBm3tYnJ41t4uxuoU8hFcTYu2xzO4uw2LLV1+udM6fujWyfmY
XM5LUoKIXR4PZdEwEDNDJZx8jwiJ95rUkZBtsHanbddT26qW6QI5RoUFg/XfWd4n9u2QiHYlFnL8
h2DsUfAvguOFdGGjSNnRx3MTgTP5p/d3xEYpnhJdo9s40ul9zjAtQIL678mR1walWqS5mnhHtiuR
00rjJV32nY5F9Wn3EU9dXuPXjLJY5LgkjaDumOLMvYj8g2EqcLi920weoiOsjR72mTM8aezVgGmw
JpudS+ymnfCMCqfjIHLUaBQPEI0USb/aGfBv+DCNUkfMcgv1u0ajXV5b7XQI+gEnre3HUiDjl7Im
IXR1QiTalgrF8c9vrGFf1Yyz3YlpliGqFl4Qov3tawqlrTCc5ob4smtCkEpx4FaWDyinJevCXrrB
7Wz8wmNuRP6eXioCsMZEjpSrKuiVF88szF1YL3E27bt7pIZKQ53F+5BLsRG5yWwNU26wG5+XNRY6
ydHq8cjzfQUo+2CcNrxNbRLeOJ2/4Tb5ja8hXVNHXESdj0V56mzeaejZEMrZizsNffhxxCZpAmCt
515k2iA5ElI0oWkul2oJaUx19d7XCZ6AWZvn5vyith3/jeRzbOoeo4DvryWYFpngRcclEFDr5IsN
3CzdCLl13zS1U/l7TgwJ4fMaoSkOaE8pbTe5k5Rq4/f+zXKvLdce3nHGt2HibtlJWuhaxRLLzuID
8VfRx6SIYFH36oWB+nVUX0w/iyXFWfsVbi5kQkPsnCI8bohpSI0xkrw6NUeydPLpeeu+UyfZ/5te
E9+sH8vw3P0rHiEWNSFZoyxejL2zL7W64FDpdtd0ou36oVBBbFAjZiHBNcnnqy+j0ZNZYJNMUeIE
fLvXLOtY8CxM3KnfGOI0u8hEVx1aDTA+XJWi7KP6vqo8xGedombJMaVetD7JcpP+9HV08R3HuD/2
i4SUvy5WWnJ5YMqo3qk0mknsFdBXJwV3NTkLRLEnCmyAUIlY/IENVPo9RAxqzp79GU3iwwW/dYlC
Cpk+z+dcnLt8K84QyK0Ui3nJQwrlNMhwgr0atgV3AsYztYV4V5AlxXf5B0rsn3mebnItpjMEd+PB
kMag6KcxdGfdkRKe2HJEz/aoZGgt0ICJTe7lP1HeBkXtH14IGVZGJw8+33TzU0lxKZDmzTBKJBZP
FOP9kqI3/+j/nqwdTYXj3zsCvtoKHviDFswpv7BUnB3c5mREBtrPB/POTcuh66Gbpq1ttOCEZtHu
135+AVs9EID+hS/8cMz52HH2eXDDyda2+xna7YTmEbwykxJO1YYQchaGWTDrF0RGhDYqjziUY2Xg
JDXgAmZ1T/DrRvXNPzpqcrqwu3Ot6pYa9FYjSivQLIseh6BR9B3jPWTpkE2x57MsmEGtK+pu738y
R65nMR0+OyPKeeNBWd/OtChIk1Ggo5KDby+TEFRmQxPVAsUBv7rplbztqR2QeWVXkl3I1gSeMuVw
GXI/WmUqC1YbJ41BDVYXoMXUnY5+Wh2vqCVGHPZWag2UUaCnTYgIifVG7FJd0l7AAWN7KbzuwWyF
hZ+AWG6rs4lesyg6pp0NayJqlZ4f/mLligwCmgQwAIzveqZLsMIz77gjJ76zp+5y+NpxMdksviNf
b9Ym7qRx+utD0y3c8rl4hAV//+hm/ohJX0JEOSrJtMls2AtEWKReTEU5pzMdsl4uiymTHy1fsVFv
iugKZCqjZKQdNPxgvFex9B7VO7SvHzpEiJwnMTR5UfglwjF+ux+2GUdrMugKIaPWAInXD1xAlgyQ
lZwBjb8HZtWGO+RosAVXYx7E0NmVnmRDh+lCPgjl5LRsPQ0NaAF+/ocQEc2DE5CK55preqUDWWa/
jqaeXA2y+IkNFGvenweUNbijlmfwjdlWFArkDvc5h63MOe+DCrz9EIqGh+R+YRFM89kXzhkiiV3I
0IoTgOtjRinXejsdc4XfPA7IjUq0KT6X4+pAgb1LJ39AvKMt3Rk+R/1Imah9+g+qVVMSYUFUv/SS
QJJ+oL6tqS3S9P1LLQ6LyznVlHS5VsR8jwq4Ua2LtNEmPPAc57mKGR6NkY0ApZZTSS42e47Wiz5f
2mGzChGAvWmRqndRWx/GEuIhOr6p6Gk05Z/lsu9TGQb8rNSHpy1sDxnzQNBpFJtLH3Il2R1OIN0I
xnWUCAHl9Z54fU5zCkNJhy3JXtmCak7tn3O/WypFRJZMOhFLD+sf+WkyB7tWf4H7OUTU8lWk8NwM
ZSJbw0gC0UpmpIrmrJSxKPYwXyyDaaZSfDyoOqXaoQr/t7fG3qtCJ5a3n9AGGDZMVT8DNIFPkv+s
3Iy1xGZ6BaHrcOtIKwxDazzBIuxH3EZVOVp+Mez0c2ebgEwTXepjYNMVv7ifSjYBlDrSpPPDhvU6
L2ovDQKYIixIUwz130hmfoI22+3s1sZn86XzCu2eenLB+62rKMfBvF/RGcxw2/V0BWtotsXIAeA+
INquT7tOG5nUeVIoxGeEVkOVfJox655uxKN3d/5HNQUPJ47xgZDLEwwj5yrzPHtA+VPI8Wbyv1/b
dT81J4j5U+FNiEh3qq78VndfV3KaDXqbzULKQAGYx8jCksXzc9AMeJ1ls43Mmw2B2V1h6O/VkHlR
q42wVT/HYfYGCyGKUyKbv4X52OcJ+D3lgcEF7XEY5etIv29vBwnHQXUvwXcuEOJpt/1PsgvE9Loh
x4mry3uHadDSqUNGoLljhGIn1IMkedmUyWnnh/eMuPLUUoDxERwymWfd3VycWBxR7GzX0XRksZWy
NtVNtMRIENqxAJlUw2YP/SdS/3KF1fpC22lB8MUn8euRMtd4NfUBo4o3THnJH/mnA7+jUPZskxby
UZnNIGpe/FVS/1Le68DqcYO9MykRW1XL3WNv9m6AHbqn6ugrRzJTJWOTl8vnEcGzeA6WICIIBw/3
xEaxjBictBkhEZynpuEnATL8kBZogKvn70j5MuEoBloJ7d7xz+wkQyG4f97BBi0YBHqZ3vBR/nXk
+Ns7RskKST/YA6ugPpfGAEnBLcf4RhdLlT0tG/UIb/YjbIyjrc5ZOBrCGTvkO7pl/jzPucFDVDUY
kMRwY5HZAJwu96cM3UQY+PpYjhB6QfYxGPggnP9ojP2PteQQNvGBGoYJaaULGLkTVi7Mt7Vk0dw3
uWd4weyQjT5ASLW4Jr3h+ZKpvvctWlqqcN666X1lRCE7PbTaIoCECPpNl6OjKbxNk+QTCcC9Jbo1
Xbq1X92LUSpccP8uDOsB5akwvBdhxsT5cTfxfPuMohi1IfEKOVrF+L/mQoET6+W7iH9D7wDO3oc6
IjZawSUoKHmtusMCYLT0YtBiyt5aHwf2STZOR0I1VGiGNCQj67/tom8BA1+rL43X7fs5cYU/rJFh
QnEqa+YN3j0AkX/fEkxBGAuy9ow/K+VqWv01fmqbyqWZjZU2O+As7cP28pauWIZrc37lypZjH6uO
sw/nkPazCGE1VkjWZIcF0JXcia5tU8XnCrDwATUL2JRGANEJzIhi7rm/TbKPH/svujWX6eT6s8gs
s7Y+tMDNMIX8AGvwihnpuYFzsIxEtqPAf/GQmBbopW2/ZocbpGGsb1uNtuJS7eAvPnxq5Sh16ccZ
9c3GZ4LOXyeRFytVTubUTSyn5LUDPwsReCkbtB8vIYYDAHZiR1jeyvXWNYSr9XFHH3O9/D67sFst
h4gzJMuBaWDXCu/cVmf+uYQzMjeF6mWebYqetEQLX65jAobQafArMR8Ykl+Vpp9QnCPCED+FxPjk
p70UWuDD/n11kdSZB4GTNu0YuHCAADvJR+49D3Z4mqmZkaWq/0JbjYV7Q72oewhaAWZ/13UntBOZ
GYckeg7NFcEZ38H+8e6iBkMFgUyDZEb7EUYOkw44IXqbh9ofIyVU9R2zokKqnXI7AJnorhjrQoUo
XgXrEeuFM887q/pbrCw5LEFYaJuI25E8A2myzfedyi1jb4/JGmWQhMuS6tY9NuDSCsZRCQtPejOV
bhgXgrB9JAZ4wrIAkIaHEbjPdNgKo2i9Q7bmN2IyrfAuzM2vJ4VTIrYOB0CZ0HADb0NmNVgWSybV
I7r2irbwuoSB/BCI3ppfQx/lx2W7oiynTK1ayQNNw0sQ58isDJ2Ct5w4OvrvBgNBk/EqVbOax6JS
y0iW7V5f78U01bGLPb0lJ7G4xVFfJOV1auS8czY5gY/fXhOM2aXRWRXTXunp55Lxl+KwUo9bZmwa
xfJ0Tb5bag+pH1ZjtDNi18cOYCDTHtIfhcD35WwZHikN0Ryw9QGDyjqOjrLQVAWRS1w2mPtjHfiM
YVMLHGNgOYQfXItwHDPdBVunZNaZnoEWHbzzbNPk3hkzDhBsBoR2JIPBkimkZQ5Y69yKhggUdWWD
hA5sj1iK6xadOrQEyvugsWiXn0H/FWiYtaQiWe8+NV0UnG0bskxQWq2ne9Tv5O5hhohEbUFU4Z/y
MFM74JlUwrHUJBCerTdBTSv7B4OZmkyQ4VQvrcjIe0vEKcZGLgN9gTxURUMFMh/23W/CBY2eVeA8
mwGZwvX9gcprJpScHmI7TKIUHd5zWvn5BUQgnE2v5foI2M/PSpbM7jM9c01PekS9P5NZPiFEzYUs
9789CQt2uk0SKEHeHdoREo9SVZWf296JzDqI7yERgMzzjZUP+Y8jd62Kp68Ai7pnuktMztHjQEhp
9liqjmzaPwaS71DNekDH6AEm8knsqTz25ovaLYwQcwqnjwH8L6vgcjnFYskRMEcqfhR/4LQHAAjU
QD6uDkzOrZficZNXBj7fbCxEoFWf7K30zz2yjobojmN+N36WDk/nrjHbyO9174DtAVyZiLB2OOou
foWDPuukKuo3BwBUcgFXEw9tcFMpFSw4H+RkLt20zsGGR1n5+2qvr+EGr0oEJ9l/WlNDEamQnlO2
r+DuRNcfZ4HvOkNnO9ENzsZPqceHiohYqu5c2ZUP9PnAJpamGSfrbhiokhTT+ddxRFzNUPAltyXJ
IdkzRiGlCXNuphqs9a5GBDzSrKWAT8TQb/mIQ2Qw399P7feXj9F9F3CizzkNN6SW/HC+48uiqbbe
WOPP3UkzYaezpGDM7kgKgd8NtaDeWIoa428Qg+2/CvEZ0kx1ikgejxI1sjb+IQYNhTPC3yGA8DYz
+TGCvE2Twtdhd67qdiCjLGC1MAnxi8WbsIVgUFSxGDjrG3YNCo5gkQJ+fHfayQ9GgE9DS4414Nbt
roZX66p5idzjkvEXPn9iMjLJwjq+zqugpmJqwpE1HkmjIiUD3RpjxSiiNIY3hfg5Azsy6I/hIP3D
QhPq4S6LDaNx2FB5TfuoLeE8+c6I9SsI7uHLT18aVeZRIhX4OvkrzuiMMOcU5TbCNIsPGDm3iTSL
OenGLjXleYo2mzEXeSPIxQkO8m9jUG8JEbTvLGAfi6CCRrKjqnSCH/56fZNJ72dU5zV3MOheAyA5
LvciLSxezPlhbFCGrkZztuolnaWkI85r/OUChU2HfoDkuVdNdlE8Jeu580yGaFjXNVFS/S7mETa/
eimnxsH+VK5u8m+lsDu2LH2dH1YjmRdcqi7zl7rAgHaxW9VJrHo+Y92DcNArWOxZ/XlHJb2mToz/
tWgabtZ7QLKZNOzoXyejyNSPEcWrmFlmZtUDEtrTZflevmCXnr75/0VJ718gd3jcUnM5RayUEWB0
9wpmGXx3I7fGZzxGGgu/xcdufC8rj4sY8gWfNCKrvqO3AJA1IgtyomGaAi3TOk0GnDVVBE3g8tIQ
syiDj4wSRjXp/fQ0fKpH9vmZrE42CGDZmHWeQ1VWADhziD50bvERXPJt8OJHTSyACyCPy48vj8C7
39hEKmk8Ct29BPapBpOrH0lwk+hztF5yxYUGcwnlTFJMS0ipwuEO8W31ASv2n8/t9J8pKBchC6Sc
tttELxbM09PlizB53K0zmAhVfuBFbXNw+wuJiPLhitcMxkU9py3i2mBz1E4UXSBg5vUGQfUugfk8
8ob86nYKBRC3bEJlTi9yet1jxGsYR7YLirui8fhTTHcel0HnLcPvhlDoczAvT5o+6RVuAs70xQ+g
H+CU+8hZ3/LOHiI08gKO0ezyRnARvpo/uguShujA/8WlGpkl0dKrrAUE6tSyfHvgoRZYvcCOivB9
rrMXfZZXNbppRRYc0Gjajt0bIasselLDouPz88cOihLldfp3DK+59aTb0x44prWwhIu0ygI4NmRR
L/U8AUAugVlXDnN85NtEtZ+k3i2x8XL8ceL9uMx1ONIYEo8OMJ8Iijzp6lTtdcME7QMAoE47wdX1
c2JT22CJAK6EHqzZ+Q1SqE38hyrm4fEtT0TKEZdktcJP6iwYRjNZv2qXPGd7SwemAUjSjxWa6p8F
aNO8neZIQEYBnIIvYXqKbZ//jhcrgWZm4BjhDOGueYd49uBQA3O9xPuNaFR8cokvnX4X+ImovqCM
/EMPsd6A7aU5qrgFbjayryPbiRUSmaf+Yi6kXmgQxOCdRuAS/oplGpaZ9nUBIrD2x6Bde5ReokTS
n0ebU01UGZ+o5eowBsFLd0RozFH+pcwxXHjdqBPw1OAxmyO3c99Aff1oZ8elX/f5/U3VYmHJ1Wfo
8l/PDq5JCFg36NSTugQfRNO2nXTeM0saV+o9Cq909cuyHWJDENMUM3GFKY9PK7tFmk2tAomWHMXl
KMAcSZuJW7QbhEeTXou6lPCLl0G+pI8RZLcZ0BHaXX3USjK79flGfMuoCydQtaQfvUhnUgC4nigV
GwMmAE20OdOj2nSjUXQX+LmHVfk5hFfNmqPijPShXf6U8pE/HvfMsx6KrmdN4c+/IAodv1sTjJak
fSW9es+/af17mMIJW8w7IYhcKG4kt7PRZLu+hz3CQhphj/6IlBqMHeWtH1EwndAgzNfaoyXa186i
sRY8bh0cXflelLmVrgL2nKyS1EPnPTj8hMJfHtI17QxHz/p+viT1Y/BqX4POokMAL/jp3i1UCnaa
+eaTFUORybNQO8h16bnU6DM8fJpX0SDFccFRJ/fKCoqv6J0FUp9H37skyu5NrLef6esV+5WnBqRs
ZuKYwIk72C6iFDr+PSTy4oASEiSdn0knLZN86AYmkFRp56bltx5D78nbf910wI11RsDy8w2TsCRx
lKSFv+4CyM+Q8fvPViJmi1xlpWdPyU65SI9PHRA+JHLrXbwDWsNg/yvGF2LsVIhgHL+fvn7ZxLRX
fmMtAzCXP2qU+K9e/OZC3VKBvTOTBFxWoC5pOxcNv1ZEYLbDD+6ZprzxolHV1HWDGnnSK5Rz0VK4
WHYwnFTTrrzqWqYXqEFpc+UBbM9CCX3GdhB0aiMPFKq3pIKrhRv7pSKTttbSz+kQJqHPntrMJWa3
3uq3MbwG03YH7/P1klPF+E3JAavio3tYgF47c73g+uK3zo6TKni6Vs+Y1U/VkF8vkmHZXeuZ8EsS
jabJoCwvdrJpHcoXwrvacHKHRgztRUxpOWulaKrlFc5/pd7x+Gn2yvaNbB1nngBx4rQGU3z1V2ls
bhkpaRw0NhcB7zSo8eHVAv1zq3zuE7B6zbyIR59DxdEEMPuYzEa6RcUhLkkadbkm9/gmItK61tFq
59gmGwA+o4NBrnXjPdgbxTwmrwV7DxL5aAXKnoMjDrLfFu8VLCV9fRC7KsVaKZVwCZlHRZSDQcZ3
LiUrLoXIsq3ngdHmCVt/DV3i+j2H0ssVXr4D8Ukheowci+SVxqwTS9NfR8Das4Tlrlxyt1SX69aj
6pUuZgAb54mooE2lYChNsT0QtNHq2mnqP9D/79Ut33kclIkSsKfAKYBMeugHBVeCLNVleq1yRS0p
xCiFK4KmWnUA3XNDgXZyNBj+jCLanbiw7aRGaMeHGXRNtTsX4s0sYD+3ka2dhhcQLCKY5KINFHBm
f/RZFDjNmOZdo0bfXpeyElRS64ZggtNYLxwxua0A8nN5bPlElgvd25t0Wqb96xoBLOHiPIDBCYrj
EpwvNhxagfBpYGEmxVSJf+Rq/GUrfBH0VGrv2AqVLVDUJcuuKuoBrCwUuuWqBr7mFL6QbJp5ZLFx
4+ADTAU2kLsanVCE3ieTGZFStj9eojGIvpNmc/jAlu3U6DcjWo4EDwCqrB5auixznmheNm7vJhaO
gk9DDKU0FyerWEZAxD9e+ac4DThHnZvBp9vk6drLQv2eAzKUZ5WMG+t6ZTFkDhy92SeIlgIwJYes
P9jRGn6cs3l19CPx23w8qEX6qQtxVoegJjJBRPzy3TeHNPSYDJk03KU/B5nmMSPicL6gXk97qd49
nc1dt/RCkXZr8/Tk8m1vypiol8RVsIPg0yGnUvR7uuz2M5rUVTbXAIQ0q7gn1mJNrdlgs1zyP2Kq
EEqsntwWDWlwPBSi9nmzNcW6u9AuBzd6piE49hDCQBfZueSovXsNtgLN7SJzpnd3JdX1YNHJmNvF
xbf5WW+g4w6lPMM2vlIVstis7/12AUvQF2xSsfvSyfbeO/ksgtZTSAmzQpoPOzpGPJXb87pwR7Rv
B6aioR8ZnIUjJycOGQka10hCIhMYlxEr/xSvUbPugWvCus8kB+wi1tveoHYd05vGdPJMzjbuBIGS
mQ7yRbzFq8CuLxZDRdjUP+zkEtAQ4tF8hbN1iFbwI0vMqtzyTEmFo8lCINDOILd/9uPhSAr57iFO
qATfptdH3hap/q4jx6xqdDUazEVzMOcpKfIss3Hnltp4BksUrhapFwITkedCQEYBhacaP5hpzqVy
eExL2w9Gq1SVBTQvw0oe3H88oIguVykGZPPZouPyyCum7GQ8VNUnAf7ZtFGHzyTF51w3INvOLbcJ
1EGuizEw6RhHIPvvCzgIVrPn5remDbTXb9MJxAxCtrZrgnLLiEpR4FdEgidbQFwXAaZGdPGgYBl9
8vBE6kRdLPF6VuiW8lLxQCYQIpdDLSP0lhMqm/lufdnlQuVWDuQMIXqSyewl503PzSNUJDWME1jT
jG5Ov/hv9kZEACZi7d66dEOm4rK78uobBlqKceJQ+m0ZG9bgmVk2m49SxUeE5UWyXra7hLuxlJkp
cNfrlHNis773DRbqBlni547ym9JKYcX0sXn37LhynbeCoI15279VwQvi8xrWd8Xv+1J7lpWNg6GP
CJSNugejpDn8nWkFXiLqRxyxPwVg2m0YtUNoTDiXKeORuRyG0PqXd3e9vUemEwQ11h925lKTz1O/
JJLJRt+IhogR+2jz3IYIkNChQYv+cYhaBt8+6BTJ6bsoAMgHK5yDPfAk+MS/NtRTwuamKLvVCHnC
G2CeYhuLHmYKD0Jn+WTWY1ne6NJrcD0Heg2/wPq6DpG+/BEeAoc6o4QLRlo0IsgbTRFcRRdf6WOS
Rf3uZhMhiXcDac1YrY0RBVsLUnVx7KIKlVfcMa2ZY7dHjN70518Hm667V1FqOMCP75d4u7/8pEPG
/GGYWJ/mr1JeAniZfkRrAh3Dj0KIRxdeIgqWc1JyswdPuN6tLl2mdPcst6HO4iZtcDwLQ7/7qHd2
tLBY5rD5BICRl8o4k6ns+296E0UQca5nZ8KXprRrO6UCLGI85Y6VUx/mxvTGgOgsXTQGZJL00V+h
pyHi7tGQbQTFTCzv05UWaUmSpFDltq97f0GnpiVcUI0DPFi4dojFOQjS4aGC/I0A4u+eke0C/o+0
fICAaiBdxZu0FeVtpm/fLJ46+8PvC1ZmBIgqnXjJB3CXDpZ848Tj9VfjLUV2FJN+c/tr7oflU3aJ
/rgY74+u0tLLqd3DN0uFarg2sJCUmKNK3t62w/1JDgbuJDMt+c3PDfd2mJgUBcuvMR7fDnHCbwSb
bGKFpx6REQFfmTHeHMJOdxhxtbp58ZcfoB6oDELbFFhd0yDvkZRC391pl8XjRbOWEov9Vo/nPEVQ
T5IvWYi3SJOPrortX6T7fRTCBEHRnuoi/WyxkCnl8z63DuOmbwG6nDmkqXIgkrabR8fa+la8+q/U
z7rjNIpEwSAw798kbdADfSbb/u05jkLZAY0SyR6SCQLZwEBiI5z1icsRqwR0kUGmHZZjt+I2PrJ6
b7KprXTGtmBmv5b0lTR+rM+Dx49W6KVcv9z8hngdey3DQgvXDQ5Ue1sxTDdE3aRCBEEHCElQAhMg
oOKas31zIm8go1ynJwy3nuI2zhtst0b5iwmD5vkbQJB4e2tgL1JqRNH/FQ5U0h6qj+GXZY+rXKrG
TEYCbkz1dKHughJmR/YK7O2ux+aq/aJg6dMDAJX09dhiC/I9XyEpFjFLQJ0qlMRfOj8cwYyeBTuM
y6Sl6ef50qtIDhYhE/v+MrmFrNQPj0z23yjje9svI+AbfITFprR8vU/bo5AhGueBun0zrciNpC+Z
RUckPP6bIMTtARHfY2EBgLsPKpcPW2tOhBKTypIbSRNGjALT/QXtQl439OniC6fUPLunNeChlNSl
vhH22pf5XMMaxBfhbqTXkx6BseRTjhQCmjaZJmivjnSlPy+TPipz1/LCk0eeb8JaBJRYkprXNy0f
wGoCqO/r3Hlv4GlP9G+mGMGgWli9Y6YhZKFcuKWE7QL8fGPF70pJX7vvuwjahgW+mEq9dcio6IhA
iLZKNsSTdvdPSnZNlOZBxQwLDctointfbc37o7sdSYd0QFrIPGlIjnESuXY0+C8du9RldYaV7Hw2
U9uDcVVr/yqd8Ah6q69bQmp2rayNZm+OezGpod8q50hxUbQHup8wogNH8MTOqfvpY/0AgzVqVrZC
+eheZqY0OYe2EfFYynIdNMLNpiC6znDttuvMABdkH4iSvn66NCBjwSjpZqg6yTYBp+D+xD0nKtqh
i6qTV7m7aL7mrBQRPUoTBXSVXXWsBoadyJ4a/dR7YxGQrIIOl0T0qfon43Xvc+bx3QNDWnkYiwJy
eUMm2JAsYCwvP81CHaOOCbzc7hCYp7ZHZtEbNrVHk8vugB3VxCQwFb0P7kbJzxnKUKzKSYE/wCLp
U4dcszATBhwoq9ZcA4i+pGXLtnQ/CLGW+fbHtmYa1Axn890Wx0C+D0RRYvYZOk+T7ZInBaH6fMpY
0gXvNBQEuTeCs0zgkIBz/s5lcHJch5/uOt/0C2r+Jd3CUi3KkIcQ24P89gQBrt/FY6Ubt9boeexp
FhXlK7vDJAtVlUrddGJtQXobwKLmnfou8FGPpkUB2NQBk2woMhIpBwIv/INNI/8eRlsZQbHpYdgN
2/a6H70CE0OIRpA9olXFJFF1/bDQI1nkXAzmgals/n28YVSwvXEUBThN/9ToBjLEu+RnxFGD5hhy
felvnIgUUfR0RYxb5Y2hbEf2ipS7KYvgtyUEzY9NSz3ot7zOsJadbDE1V2Y2Tl+0qwdQrqsdw1LG
Ms7qFD+kibvwjpTSwLrJuSPJyzoVGFtVZIvO4F2tO8gbug5Yo4J0KTHD8MEeBIm3tFmJTuIaxAgj
v+o/mPDjjpCbIfL62FSWZAPh0WfCtDnZEPDK2QFC2NdfUqNsn5FdAeVOP54tuZpaXEnFSgbM5TiF
bD3JCgrDL7mPbfLqTyW1owQKbeCUkPSUqdJlaVLqtr+rihDp6lZqSnjHTx5EU+cEwb7Rj0UFMDmj
7qUQNcWRiPdEUanfC19wF9FGDFdIdG906XVpojhFsy4lbHnwzMd79bcP3iqFbbgi5vY5PByPTtR5
3QIqWAO/s43TsXxcXIoaQ/+vx/DZUtqU1PhVONvq6NqsjFiSB56G85kOTZgs71AOu8MpjoZOdDyh
FTKp7IzOtj+UNTGZIFrRkNfmRb9FcXO3X0Z+pQ5dJ8YM7p3erJlsMZLVFKXw2cSQFFQ2vyH4ozCX
08s1nRR5u8iVnt+Pt3slhc8wZ9cyox8h0VzUVyl3Oki2GUz5y0ISN65V1/8dc3W11X5mX+/ry0SL
0nBFSw9QuKcBXiRY7rtazje4xO6QzXvRNjbd6Kq2YO0BOSVGcy0lKKBq/jApNAKCXOpIlxVPL+X7
y1GlaXDxC4xWqrw+/y4d6p6cOOgH3kkvkPJupcyj8jx9pyVxemG2wlRkR2o+2zPJF853A54SR+Uj
WhlcfZ80vQmNN0QGvr3yeVVaDC0dtNSLPHZRlck5qwCPdZScelXEqhfcG3G3MHNZtaxPXEEpVd/d
C0jIUMpw1n5PkIfXcNoJd0BR8nG26H1ZUwQF/PITXwoj6c86jDCKxxKfkgVfJnLZO+ysy3JAKm9j
eFC3h6ZYdBIkvqzgDyIbDrODWmXjNv40VlSF19BlA4KO0tlfeJqFhjrjMWYywFZ+Y8ij3OjWlpgM
DaPKlk5RUPIUeevehWLxyya90TusGOHHiKy1aY4saMM9NfSeYOcatSEi4VxyMGU6dhrn4xcblZAG
iQVnmszyzVZbUGtm+pUcPbyI37t+2fVZs70fGegjzveNattHi7rbLOk2j/m6VgRM5zLpskcnnR9O
WhH7d9T0j9TCVl2nmdLOvsb5wrtoxfIyMGIgGb5AEl79BVtKjMzGHSJKVXab0yMUAoemlJWsfRwJ
Xk4WA+9pEPzAkNOI/eR5cbTXQcDhMgSNJeVtcyLErQMEwWuROvV3iJcXN00GFgtBKlLOr5tu8DKl
rJGgZmTL8sy6O+Ff6tCMEuQvoFrr8hvFD3Re+UsNny/axE+FWzz3zC4IScRT3IZW7rsr3uXNVeeS
UVWBP9M/G4gEbu3bS/+HOJAJFnvN+SobgSWyDJYBHaM2vL/sqONOLBHcBevcfzIbT0/+8tY5lPGd
vzb8DoWvgRAwX7TOrSB1AEaR63OCoI/fxK6EMRv+z6RNbTUM2gLvcYZtKaaoZ6Wiosp+Qyknh0HZ
0904xW3/1sXplgmtkN0jCjbrjTvCgScnMIT3VXdhMaG6kC12icdtlbzcJYVRL4C7DrQvaaiejAum
DMBLn+DdyRCQNRogvn+C4LYaGmJgLYjD6Uz7V7Keap1grGMuIJIfy0Gc4qehGAyAhclv+MN6ncmc
2vGNY2TeanI+HGS4xkUAEEe2pkTFoPWElMrOElEdnrbAvzEwCYXPIyIBu0xH016Jquuie2Cef8Re
W7njfoM/0quqvYYAUAeDoImU8bdNNd9Vcxha38v1LKqL1DWSrnYYK+uWB7oORtYtbloxdCaVqiOS
ZbzWAzUu9rrZaNAKoE8GP/GQgdSiU1VQtjcatYWDniRbEB8Uz1uojJEy1qUtcBTUD3ag0pQUkz66
GgIs4WcevVhbsW7hXz0U0/cs07yyaw+Dl4A87hlIvtfmfidleYOXDVk3MD4A7ZFLb3Ec65nKzkXj
rMJiYOycT9aTxkt/9VuD5Btcpd39Qmil27CTgzVrLMZgMhlyKAjNwb5oUJmC4QYUauVWVGhOZIQn
b8Ook2Xd/KPjFBeUKR0jmjuuwvFfCBF37nNwvDosyZCWv81MU86GXeQWMS2lNSVtWQxYTkTkV/40
iEf1KDKFul9y5Mn21igvikF2dehCcUU0/d5IpQczgwCWabG2nAn37fmODAw6hAC7L1RWmFfn/I9W
bnETHLRqEu91ogO6+RiyptaKTEx1OEVthEWydQgZdvsQZSFVrstTl23SV88Q0z4yJp755TXk1mEI
d+bJHq5L+vzgmmImQlOV2YXC3105B4ZfiMDvy9NAR+hmXeVbxaOpG1ptHUTJ7zcBc5Ho9uE3RDUb
eGsG1OMlc94hoJ2G5tDVjVWmuXPHLtQZBDeSxmMf2+TgUUcdCgItjkdi1lIDLMkkue+r4I004j76
i+yqNr9HwHiSawecK7cl3HnxpgYVRxpWcoi3xMDy0F32tAgje5DZBAUmzps9oyvo+YlmbooDVcf6
Pdn4VoeD3q/kJmUOVIOR0IJx/V8o31BnwzJ8be6DMRIDj7kSYYk4dvvPrG8vkB5gQU9sZqMfQ2y9
03nmv2FW+oe+dNg9ReJs6QQR8oj5clQhaAJ/h5LcZdtjvvABV9LmezMcupGgKSEsnL1sfzj+/m5u
3YRF9DwzRSsqTcBJTyV+FTdS4ShcsGLGdEe81m/n0VMbwg5ZYteP+CIuk1c13XKOifWrGj77661f
6PeaJEwWQcsEhvfMa4G/eDRsr+pXZ+vbWfnLR90VWd4fwVeKXghC4iOYstPGJXJkRvsQJR/QL588
FdmLHMpaL4K6qSUHFVWeg6jH18kCqg22/Xs5YtuDKhZYkd6lmfUD/HRMeVU3C2rUGdj/c0yqESI9
WdepamxFnpJy6xaVED/laA688E8/BErHabndfra3aUz59EHi9sHhcNonfmqPBen8ngI9SkCFkBfE
tI5CgEGatttMnqHU49kkclujX8urwI2/rBmQf6GhQRvpXH5rb1lYsZvVthQnwiRHha4V1wjThFZW
opclUrCqvyLOldgfpy5xAETg/p11UxkQ8r6KbGU7njVlVuNpY60vttFUyerd8qKQbCpyKjM8TXyU
8NCcEJxMoye3pZkfQCQn1QEkLzx7/z8kLtW9aFLyz+mqKSRCyyM8Mmnjupm5sYZKSHI5JsiUCuD/
vA8aX6zH3gS4S+cOZ2tH+mj5C3h6bC7xKUeZAhxcNUNOvzudl3Zqh9jcRVm+iLlE47ghODcb5kR5
uJ9upFTn5MW1ZfhKl3gkRdDmO1gmVufk4HWSuAegK1e/kTdfgsDm4sSiZT3W5I+ZGuK4FVnXhjXP
VrBAqCoHYsvLQH1vLMWi3kZzN24CV6Ft7MfcGh66p4QdUdf6dmasXuXRsFyOCpX+5tl3/0Az5ro6
tM62MI9e/XPufYcUpZnI1osiSNcSFFclQnOzZxHBSsZN8fV6GDq4RqYzjWyGwXqvznib0gjAMEgN
jGU7NFx+27F6yrkRnHnosg+VetBgxu8XuM7LCWL6Bk8KhXKlolP1eX4WHTR1HbDz1pgd2CpgCFhM
/C85BFyHyvZXvbRYo4qEmxqkCCQqya8kTyT8YhI8Mg3CjuSu5cYXhHxIUM/TjeayGsEfEVNbZQdY
dcPQo0tGWNV+zBD00S/E5TKc1NebVvMBtleoqK9hC0BKsK23nkuC2oOF8kSutPnsKhPYvjQLVd+H
6sGRtgwPvlkruDqqrBx4rIOjZUiTSq4M6jFLNH5xsX7JX6nw7zqcYmzU9Mi4muVrdy+sfu0VPpQt
g1zxhfaW0R9Ok/uZx6VTFNJD2t5vtfRMi0q1RxYm24N+/FNEPLSPY2QUudjNN5xNzRI3eMywOxFo
Qugo3qoeswzspMPypsWHqIOfCqRbOu+w0GdsqcwoU1sc2xbD8mlQbqqMf+x5TEMZfX0FtWbdB20f
dmT1eFX0T3ZhWDsknspwZZXxO0JFBGzqcAP/cA49iiWETKxKh+BVTeEvKCIH16LB1TcEKRKBE7HB
8YbYZ+AXo5yYVqfzgEzh4L7N6eqjwbrqi38rsdGfeSbQo/wxWviP6j93yMrEaEDBJYLS7dAZmwuC
In6uEXcU6HmMYAFtHSIy4YmrjpFgaO2Ahi684L8z+H4qct6pUYwT0Kr7lU0trtgYZwaP3tjD/xZ4
DnCM8X6L/A7ev1nxdK6ASKMKowFS5p6t4sIs/sZlIjo5sVtQo7T7g71aNDmY9IU8YUQe7U/Tpn4M
vOIAHzJOzVmwj3V7G5KxcHvMgF9u06q1T2yqMuYmd22QmbA0jbuFLVnflnmJd2BBRKBgGT97VB4C
q6K8ePpVJt57+fg/HyY75lLxcW0KOIEZI6KyyIRpSfTd7vRjVJM61nqm5ccM+FExy3du1npq1DcE
HaGgwcqBsm/Hhlx8JGEVDkDI4ispSGkl22nGhAOrJWWlqBBgKSgqt2wbmJSOscAUwMLeW4PxmAVo
gJRj9ji2WtH6pvi6Z9V8YYVjiUbfJt7/iz1Z2e75nm/pRNTgn+x0JS1z7Uoezl9degNNAk44eaQV
Qt7VspiPS1GvPnwsyHGpWh7y7uErU7Ar04ar8u+7ouRJdBtQP9QIdMwBzaIRDwhGrvQrGzAJulW3
VkyrpfwM4tCZyT1QtxwDzl1mQPkO3h+j8wRd+ngzsTLf0/mx3+2p5yPtgi1Rglh2/JbpckbsJq+E
9p40bz0W6mGhInlYTG6RtSAd0VRfVi5AwsCsi7tyqf/CaoEiGnzNttyz0OFt4uK+CGYuDAkvnTYS
II5OM6JUWAASXbFO52kggX4wHi4xd1/cKZBa3pvWeBSIOfye1tiuOWmQlbR8N0cGT4KEs+wf4LOz
b0wSv7vbgM/gkb/E+u8RoIwFSSoglecSmkWaWZp25TmudZdbZds5GFaCKPYgq8lf4x94p9ZualtU
TtbOGNGKpoiYSpOvsvpRAhdo7mz1y7g6C7eTjo1bVoszEiWYQXftb5gcrvmC1KpULJ5bIgBAJ7S9
lchnP7kSvRl21Rm4wnrpa7U+ofrH8i+CDDJqMeMILjhnId2elP9jvQoaAYpRVjySidnZiKw0AF/u
npt1HOE7PCo/aGFjQR6pPmbZuPTY0oDbrYcpL6jHVCbCVMM6NzkrRpKdGdoEOLNsI0EfT/w9+0Ff
Hhc2DO6uK3ILFC5QFnnbSI5+iU96CbFILSo1q6OwLRJ2zi65rRIfkGcBdWwASl0LD+R40cQC7UBl
Jm3OCGiTU1f8Xq16NbbOkirc/ebZ69pocPt17Gx+WDiaJcDNm1S4FCps4U0sU94IqKS11g+XoP/v
vQ1ojzaTvnURlolR0uCPp67cjXzTI8cUsVkncbZGhls53Ph1bSKAHytoZX6XmP+C5QukLgWzWo9t
KmzgOUbjUSFGhJsVPqAeKP+1Uw4dRX4/ymju+cI4qd4AgHOwpNPapD4WQu5HmGIKswPsma2toPmz
b6Eq9NURU01bUa+FLCyoM20YXI+wiK9ns/lJzvAXVexmmZ61iKQSEz2pJI87UsxNlW1GGaGXYS01
YhmIkpNxlIVrtLpygcmmQPRT+VXo1QkQ3ciZ4WgW46RMkr161/3hCrsCTO9nDm2jSXd2qw8Q/Y9B
PbxEaz2K7k1ZTGwhVqIAe6dSVNWp7RAWxBGLIV7v/6Os4nRAV60o+fMCExn/gB3C8l//tdnb8DeR
2CeDxIQuR5yo5Gn71h3J5D2kzKPkXh+Qgcactz1dbAaTpZLWBNcdOxSnbKsap0kn0B+O/++83dtd
zMPRWJJMKo+CuKsVCMuzgQM/N2ISSaq3VvDD3geJmrSoRNMgtlG/P9C8KLoEXmfnB5Q39jqqXlgi
0pMdJw1DTMEz4P+YfeKgSB0q8uXWJTKi3Hyih9OISORIXXpkWxUyIzhL2jlYilv0smNzVEDEp11x
IPvEhgQvvet0D3tQ2h44yd1aCMAfGCKjBBBgkjOTsYfEcB0DQ37flBzsY0mW6mHnJLTsO6oGsXzP
DdnulL4a7HTFd97EmrBgqmwdwfRvrqqfxKqJoMcQGWocx+stIFrQ8txjM4KYACPwBro4SljCSKRc
eaU1INdKkL85UtiVL5z/D4dnBVqnaK2rVK95+bpO1Pa78HS078KsMz1qfag0WdDQaAt0v6Dl5wGT
i0spZsa/eVlFuFJs6D5uXci1mlMYbS069y1321S25RqM+OOl6N5ksBlGWYdcu991X1ra6ysUgC/J
j6e8gYLuFh3o7nGmcbftTGYP0ThwxENLhGoaPgf6B/5ZdbQeTDZEm7ulA5TeRLfUP4fdKMjW546K
o6BNSVrB/V6/k47qd+b+pX45c0oD88zX2yJRRIYwdlrmLnr/mNUzIqKLBOtzI1PbJflfLikxe4W7
mw9x9RNg9YseC5Z5u90V+PVNBxviY3+cTNbJVJXGkglU5UPDYfVmyN3e7sTuX9btVigEJVNnnEHv
KMfe28g3JWhGGmRXe1GsMMRBnJG6PowZ/lzX+HuP9yHRE/D/l8WrqAD/rRTh7ZhmM98GqrZP5NKN
usX5OXCUwEr0gkpwWq+I0h3SWlTNC6iHotFjLyrkkQCCldRtuRH/EYIPj5xf3J/tfzcE434cHsnV
I+jg7IUvYl+b4qZ/fdKb8uqYTD6mtz8bxGONpXkniIagZFVXUrs8OyRO0JjKnGV9EZOvfzv2iCc1
xL/7jPNDPd2/LctQQghGBtaC2af3qZHeAQtEFbanDyxws1MMg55zynnqIgHxSLsjqFwg+nwoOxtP
XwY0xcAK9zNKQI0jlewW4ZuyB1TAV1B2eatqqC7SbuZVB8YyP+Y4R5F/6RjOf+jVVsB0JzgcyHop
KnRaBnlIbSssE+q/UHZqa6pD3NrVXebzDR4ZO1kuXKngz9Am7OO/4FI8edfXBfsPU3yMXg8vgB5A
2rzjltQi0uptu+w1suBDTNNO/xPYAvr/MKVk26UGzXDyLudBNIJGspHWR1dX08yNIy0ckJawred7
iYEf1IaoiK24sn+NsKDeeiZhHVFiN8LCGJEmOG7gTTp1uIN3NkuMnjRwWzWePKVO+aAT0wfNayif
G/A2gtBNTaLnmUaK7ChMDlozIYQUTrY+68JuVnhbf1fH97CGrCANdp/x5Yw4wxLHVTDMwMWD/pzf
k0fdpYP8ol49DlbR7esG78QkguPcRYrxdNYw2IVjDWtM3+f45wJXy06iUbE139q4vyvPtHo7xFPG
NW+pS4MWY9AAtzmVG5bwJDIyh9R4WRGS84kdbhWa2N/PCP0vV0wPoZJyRNM3Oq/QOKflCQQWwLFB
O1e6NAEXiwD3+Vb6aDFb+eB1rGZN0SBxmmP1Bpr6vksFRXuow+VX8ik5OTFv2Ecf7EbumGw9bMsF
NooABOjMwxsQiZW4+Jece4AQK9ZbEt98USyO++VdW9d4A5vYamPLAdzoPHV4dbT6+Hm3iCaWXWsB
lhtzcoo7adDbK6OnNKAP6xwqsa8mBWWojM0ofFmobJ22OTzoGEBfpUkC2yvnnHhJkEaGHnX8+V0a
kkl6cVD/N8EDDew/efDW5L4nW7lFVPAFQU0Ke5YL8NVLvbGUwN+LbtmxfyrAbRGrdQ8oT/hEYClI
9BjKytC+QuCbOsSsi1DikQNTLTbSQLGD1M93QvTGhrh45+5Ut9PAhsqi/IAVjd+eqU0QtF8wApR+
m6OtLr5aiWpJfDUAC5ij+5AqWKuK5ng0NXplH78Z7owMh9DLijh69Q1g6quY+6zK+DkflGc9TPDA
FiyQwz+bWM3rE4r5ikPFdb4lDvfqCyk7eMZkmmw8jnFObxtWP1yBmkK9+6vqScia/a73ea2h644P
5+vaKCIRYEnoJqAqtBomVIOJ28ulkHtD9Qw5Nm7nZUWV6Tt9yLbe4p47zPSgJr3j1yay63ndHQeJ
Qr8aIHO+6gwzmSuDYS57j7o1mKwdsMCykSXKLJG4XYp7JCSGtmVLOMMWoifLZ7nXydiNoehngehH
0MNjESaNIWlsHbHjif2QBmFbgMxhpMtoCmHsrhVSKXiKCUKxrpAjoqAR0aXD2cfHQmj4FaBsN0+R
GxxsN3orM85rLkNNpkabMr+4Xz383C9+UrakqbbxdNWE7n8PEFk367kz/gmhoy0e3FJhOCT5tDDB
fCWha0A8oUPGzBXloulq6R4H7+/F+Y69EmtX/Aga/2NuhWSY+Fo1HnHElfyPpCcNooXVDvdsBDNU
839mBprM72nZFrCOx2pqFf2kmw0n3ddXDdDy9YHzKfKTYG2W2i/4pikiu2kcF9aiDR4xLcbW9jVU
T7y9f/HaU+lnwAVAmgRA29VA1cA4ApVFVrmOyXEvzYvSkx2vsAjviWeNMn0eSEyj9T/zRcL4cYhZ
7W8XwfrqFDifYIQ8JJjoJiim/JTMEBcaMm3HbObNJgM1VJuYsNS2/KB2RoAkcIvT4eX4vcg2Cq7V
DY0nWBtmdC0A/Rhbj6u7MXycjJAQQ89vYN9eLjyy8X52l8L+InknhgfMQFsNI6R18qZsH1JxaTnD
ErEuO+bQxlSO1/qnHwK9Z8yFNpCTRxFN4IBFhnFf3ck42wAvDrQ9rvygawH1beiAiQXDpC26ZpIg
tYG3JcFtp2OpPd1Bb9cIYJlyH+idQPBKnDC4sRpsrttFvaReKH2dutDMnBR6vj08DxYBL+pYNqiD
SRxr+D5ltbsqlrVUSggqbkV5nusokcsyIpAFoz3mZA6weEBG/WOE/hzgbPSeT4Xl1VWUrBl2cVPu
GieYuoRjeNb3Y7bP2DtzZlv/IItJ1ixcWSF734sismiuPP3fpCMi60EN2OKKrfXB4g7LE0xP2nYP
P3NJZlYYC63HTi5pctnG4QX7d98Hg8NQBw+Ifyn+Ryw20pM0uTbR2sufhAIILWHD7B1MGr62jHwj
3q5MKJ3430yj9fIlQ6AMpONRZywM0+DyRdgtqof4MKD137bqCnZ6YCxrKkMvRqFV8T13tvd+K7Ht
0CnqLqhsq+ephS+ThmgMISXqZaeJd7e9yPqUv0+d/4iMoYy7pWVY6up9U2PrlUlm3LYbvXumKZdY
cleQKuMwNu9sqIZYEoMKdjGjotzN+EBpkJLYaZMdxFslFElfkW/DqY/o3zCtFPhqbW1j8g8yhSuS
Qq8+iVZBmXNq8n0dfgtQQe5jFYpC49gtSpE42gkXIHkI4KfJ1GOrM4790pMRpKxTPVTUHUB+Skhu
lIxy4V+Je0BW2ATN1mrdfmsZ+cWTdCtqQmpkyd0VyDDYXN0GaFngCxpGknquDXhN9xzkU4v8k4Fb
bNdDMQ7xRWgt/VupN/yNb36wWQsHSu1tgQjMvJ802Hq/AahRdsG5RNpoPakP4EOHQQdjA+xjNuJK
EfpgAsUw4Kl+69VfeMLBr09Jh5QY39POq61XdBNME8V0BZFK7VfWecNbVKAk9I7fXxvWDj43W6Sb
qZVfeGYEzqlX0uKdVW3Hqj96JR6J634mVhTnAAu4BUYpLbe6P6cSxaPOS+b6iMvfNL+eHqtom+yI
r66wXxnnoJfHvU/K6hcYrUJ2gNRvK1wYpYYtCwCAE0kb0/82QTdu1qK7Q5qbbR4ImIFhUSW/Ph7Z
vZSbHftefumPq2D5u+/xq5FbwmI4u8UozriAXJjqXyziCu7jEAnk3XxEIX/Npms4m4m0VSWyEgWl
L35raRI2Pmxi2rvz3O2zSdWNIKzmwlxnt5+IG2KyHIdXJNsrT+1eq0jRVoBVm8Mk+zNVYYh833m4
UIRvfubvxE5ts5kM3AXIR1quXwi613dbGEePJnuKH/t9ru/Onfpc0qyff7l4YW+7N77lIG+wdwb9
S4B+SWsKVoMb1YrZKjdUJ0WKChmrrbx2Sl/yuzrD3W1rz295kOEho1rRB7zznaQqvcQtY6UKKcVh
ILiQbxAGNzBuGiveYPtOgeHh4RZkEwxByCuIeh14tEObo8dQkT7x5em8Cp+t1u58KCbLnbZIyGo+
nsOHAOjwcHl4L8k0N+sb5SCWYJJajs1APcciYXZZ9pd2uyy9LHwJPcCY1GVu69hp2dv7POKBuYY3
XTgbpupDPjr0GCs1WQ3Za0+cC8F/vnLuMJhFZNf1SxoTMnu7dxZ/gS8+WtB23H40lKwGcH0gqTXe
oUxRV70B9avLJuxh08+6g9KKw8Yg3AHFuyZmq9j2DclBCL5dkXeG7I1WOuZOp96N/6MxE7jZiwN1
fG8oe04onjRH/8IoSGH1suZZ4YxyVqIFhu04GKIA+9JyKk3fldKT04vA6AO6SBfYNqc76K9bHKYU
nQJOSLIGDbmk2gbCn1fkp5PsL6m7FzFOY8Io+ET/nb4L8w9olgaSZlbjzyxmmvOF/rBqvPR9zIML
LLIZfQ/iLF2dyQfMJ51h06zvtVdb3QZjPbuJc4acCs2+dGv4UGI5ijusfOZg8nDw02Um13Dsi/5U
kqyNOqgfPa92KwX+eWf4rEnJkk3OGMcZ60R+/qUjilSKjrSJHnK9H4LjAkgwUh1qe9u43KlQ9n44
hFm152LKkThEQp6ORCJVV64kBVQFMDb/ZeSlJh7/LDeDMVUow99+KKHyc1VcvO8k+5haoV0uDX3W
Brl4oEhO+d6MzGVw3PTJKSznjpFlBZhdP6bXd+nXZaU++Gg/MDSaMiOTOFCzYZMgK4J/PsWZSbKn
mHx2Ic/CfyQcx9fSKYJJNoLZy98Ii/H0WwUmX0vhltfJ40mKaU2TwPrEMx6A5OwjnVYdYHwqkEbF
iBVGvqAaG7CuurZmI2v0JwwLIV5Nz5wXvoQ/ev4NJ4uphw/NXDTAKv+6RTwNe/ts9txB5pN3/gq2
ZczvgwDMwjAtWjDHDzFkLIVRMROlwT2pr1wTtKq+tyUwLWHbTgzhLIfQxNjM0EI44mT2CpEIcqDM
ZMMeEkfPtEzC7NM7Vqwu3NtSezDuvwTgNisnEjOuPKCLCyfWkjU4Qya1JDCcVDwByyH0JHM6+8J5
26PE1+nqoakr3oHVqT8HMiY8ekl0sZUCWZOFgSuVdWujiu8B2AAq4Mdny6CBpQ2ksRm18YMrQ1bh
ZI2vV01GGuqBipGrcUll1S4R1pEVmgu4AQLY0SrMypBPOjXPgV4xQ/3gRKuuGsgiaqqyBvi7orSK
Uw1jDtlkEwfRz6Jt0rVq3K+enyT/pbRMFgXUnSYr6eLYPdJ5nVPuWPtqLeD9WYqZAo+oSqoRlzHp
b015GJMzdXEfIjJ0BWy8MolPhSRcWx5dKT3ppzWtGi+GvgNUAfo/TPfiaDhNAjh8SKUQS8qvgblr
G+ikrPFdBd41aRuR2IppdeW8rW2qETLuqd1eBtg7sKVG7a7X0nZ/gQCk/ybQlhBlFm32zzAeUHuY
WxNN0RvTwhxrKGPazR/0jUbvBDzJgzxh2zthhjIYxHb2hAMCL8XcnmQ7kOnTfXHJJ+ncPf0UhOpb
y3S1hnyZTPKbpCxMPfWUacmhMEtKl6IitZwjBr+TJlbjQPY5N0+d+NUDJ0iaf5iNs+mEfe4qVRsI
BxkPxXz/dm9gyXrSZzdpVdGCI0H+CEXiIf85AplkwitWPLshUML+D+zV1KO8wuEjUzvDbIVNLz75
FeKzydP/VnAe9UqTzJQYq4b9eP4fbMoBi9Uyu1WxsK9DZgkiSdaR+tSlqq6oT8NXpg9jT7Eq7+I3
6KX2ldjuZqJnQ2dpDJn6Yg4wKASH8FfIkSsatD1JAtXmt9VAZXjZ79hRK+x19B7m2WS11at+ICRv
buNLuweKZo8+zIlfxNWV+nCXsp61Hs08o0cwS50+sTalv0SBAOoclYcTp3bQ6rkrEHAngNLlHQ8L
P3m6n8QKXZwFjtxCKTdMQljngIY3n2xF8GKrL4FbZX1ahWJQPhY5Mb4I0IAZ3j9kC0rnPBT9h9un
LsJrsc2GhzfwFCgUWjwl1/EGzSd6Zc1rSd1rhILnuiHtJK7oujxTy9+PxVnF4rQ6uCy+AEnIHrjf
/53sy7+fRyHbFK7fMPqgGIfMoKhOPIb6w9z3rCQH9njBRmI5iWA6FcIyAwCyK4O+Ecw8TnYWjWi/
nuESo/KJIV9ryxvdMfVOMV0yBgQkbMp3OXOSpf3q+IlT1OdZhvGTaIqXISkHjzDvzgYnvcYGl5hR
LWfTGi/4LqPpBE45cYV5wbA/z/X9BZE/xUWQpXvpXKnGWXNW6BWYOFgNV4qM3RFdeIrBvxFQYIL7
tQlQRsFe2EKRPlvR97ejiOPEu3+Kbb9hOpj1VhlhTpOvSBAqLjYGxFLZwHElOyYWjpOnEGS+VyDM
AinKZ+vbI10ZZsJ6GFvGf1+0p45taz5ZLck2vMsDfnHKCHEEZPZMjjSdi27Q0lA8MGPUYWSU2c3+
bHqr3hwOKELpR6/HNFkpukBcuGFiDekzeeKesyY+D/xZ//MkJNcXVS1kY+iS0Vq6JjtcxtP1tfpC
advQSRWbvJZwlhNyNFS4H3ZytW7nqMtP6hFmEBVKlqmixiNQk5AAgV4OkK9edk164BcJeCo3sKFi
/4sGYTDEgXnKgEsFyrY0eZgfrVBF4RLSdOBXXCbuLXeDZ5nO1VgKNJwD7mrSbxkjPMBS7EgUKFGd
tEfT4sZIj64UoSfFo0p21Z4HgtIIP2xpF74vlJihOY98z0MrQ2XlKk/OwjsKF2g/3i0ooCRW9Cqq
u1zvXzmj0Z5/gAvot6soiceI4UW4MZ3lWWx0TCwjSwJHhH2Y9ZU1vZ0TXTBj4N7ZIW5MzyFMDXNY
mrcG7LoVh8/2ptF4Gc37/I+PB9A+JvDWzVPL/cx4Sri/P3Jj5xc+wzGu0mv5rZd62/IfBw2gaqZ1
8vBPizZ0x45FEETt1Hr/RusOECJsqMxBhZIP6uT05vKsw8+XUK9YnSZeRwGoEZNalp+1kFmokHB3
1H42pqtJ9Yt2RVgZh2kjI/QVt2kmLgp8xBMjiht8LFp8eJSubTdHNNE7k5yPcKWmA2ZAtPGXlwu+
Nhxgr14BiasIViW2ocTtujp8dmSc7sjnatLQYRJoTxL2Q1YvOa/mr1DS9dbrUsr0mAylhDyBBVAx
K4rfsNr3L9PIz7PcjsLvhNDNi1CIKVKoInAx2Ur8rGIpspyl5j/5KJv7AEu/z06aUgqfkjQJlyRz
FFLfb5TAAWXCMY78bb7mxfbYqCj6UXtU1p+c+o6wmsANkVIyn7xm2AK+NojWLheyd21zOYu44/X+
+SsVUpU5kylU5QRgUKIXeHeg75lnxKiGSLwIidbzgSK/u9TyLa1qKKqSybarAzil7DM+SStGiSG7
jMrkIPRWvvoWLFKhu0Jvdb9H9p0bcAPisa57AgsPL+MhEY39JPXRr8NenU3K0wvaALEDC2jVaZbx
bvKIVFORVvaZzNUapqQOl4QxIAFfA1FnzC6tmEWoctkJfxIy8qEMgYEUSA4iHV9Zdm82BmjN3bxl
1whTbc3i+00tiQ7LuTfoBdhG6cfGJVA14XUxHdectfb2kca/d+qm9CA8zl9MZx6DFGJ4458gCarl
qLUTfMyMZWOedS4CFfUg7qe6ghmimh4dkLu21iEKPx1Gs1KKGwEjEp0VIt8aL5PX1ARyTlbFCZAP
fjZXjckdMWZRCgq5ODli0TlW2dQA6ji1MgH/6cLQ/7TQinmvPDVvxHIzHeKBvFGu6Hhl6/PrNhrU
ZY+i1PZJD56WjrjuSNzOz8IlWv8N/KynV0g16w5TDzUD6NHVZOFzT/ep+PB8NCqY3S9zEzt1xjZ3
cam9yY7eBJ9+EeyARr0uVlQ33KFxE7p709XSrewgpbFe+JFAIcplXY316HJ0KG9v30bWRjlttZTk
H2bcTSq+QbUYxNV+OZmNWRRkSKdC+iB5NpG0sPyqBNADlzJNjU3806MxBx3CejagJ7Eq4a1g/i4V
Bt8yKJbCnvlY4Tj3uWBpMQUk9JAUxTK6gnUS+POMSqeuXYg/kf5sFP9Yv6yyLW9+nER/knR0S5bG
ABcfNXBW7by7we91CnNwBQUjvbOSBxuyjTPFfHX25kBwBxyvvD9ngyDKWEcx5/bNbOCc5rgNljzC
pjXOe3mdKIr6PslTuU7FpMDuq6VieoV4FlFMVgpU5fTdF/49NkuoP3xXSlSzj+U2TpeEi92yGT3L
Otm4EemLyceDTfgI8o5okvyAfsq/TeY6XtJSbnKsLPJLiNKtRMCac7vHKAEQ2Iip3wIhVS9+kFFp
0XoNUTUhbpKa/nzGE5cUx8ot4pBQTdu9G8hf9WOZpe99i9kmqrrU6iapA11NjiGvACjn6j+RZ4VX
f8WRpAr0aLW9ubqi4KNzycrmqSzIwMPileDNww1yagd2qihrhEAI3RSLVBEiWGfgGOFdXCo1PtiQ
45BHbwrYFckUNI3So48HrqPUnCM/TSkkjLLz67uVAsf9wowuGKTat2LiVGQKm4hlWJpN+IQqnC7m
Qjqhnk00ckmZsNyeYIPAsuahQxEtcGWlgfKU6qEXZw1uyi02LjAGzho7qoqgy0CZ8Wtlkq/eps1Y
keRXGy33s9mrU1aOS0Nys4IOb2G678Q7NxxJHF5v7Z0J8xAVkaBStMITehxlAKobby9cMAajl4p3
06wa0p1QTjLdaHvJUENrbLjMyGeAAm99f71NPIzRBvP46DpvuVKn5KzULFw3azbNstCvak6itFPV
SkTfZzuFbNXr1iELIZs6v6U9ILl8vRqXXxtbnwbtrl1Mdk3YsP8ZCNfgAFiivkj660XCDhELdXUN
nN/GauSNxyRkM8zmRotnJ37MFGznjfztoF0wzemxCMDhu2Ntxb4wWvpLsNPscccTW/V33aVjW1kJ
PLx7ouxJRQi2QtkrghWIvOrfz32aY2gy8k7z6QWX7RHOYPDWgtz5kRS8qRJlhFPPhPrlGIRDN9Ar
Pwi2HYTwPxKNJLni/a0d/uijvWBOjX2rk19otK//SfnibodG0SAT4cQ5eavW79M0ulYqvQpRiMS0
zOmNT+6B96BkvKl478KE3wYyfq5m2oJxPtFPwBVyoX24WDHFk+jB4S1zLrjIDqZyK49cTAbFTwQc
ZvNf/ThBU0B0fq5MsqPBtvUYEzAPzmxGy/C04prDCArkv6DEMecCkRpdPjYAuuhFzfw4nFPEmN0/
TWKYizORuPXdqcEgpKfZO/TuURF8kprfubckoKBl4pIWVS75emEJOEir0KHYNZX7Mxdqg73dqMbz
sf3DnUCeZF4tnfSkbxLN6h3+t13hjVpXiZ0G+DSAHNczgc0UAt197kLd3nWcBsoQIyqmLYZZymYl
JcHZ8/7ZStBF+Fb11gwbUahKFLuSInyYnez1BYCOCz+eKVkC2s9H5xh8uJpiCmgtJcpsUObqZnOj
7zozSOf6aSayZw7uvPsn3ioWtaBKZfcUItHq4SPf2kXOzbI6YAbovpNwCx+zBPuIAkAEA6C23mEV
CWBomhVgJqu53KcOzsjjUc2gzdWatx8Fn+JLfBVQ3DAiSqLdv2evaoWveJilKy4EYzSALag25eeO
QdJBpmEj7mvcAcQYyHLq4E4NoWx8a8cwCdRyI8557sNx7zey0qXZ4AB+mfqYpzj9a6aWOYwGUoCk
BwnrGcYCuLZqDAYgZJKMY20fhWPU2NchxQ1mEIf09OMzLbdfu+PKl7P20wxWz+u5rkjMWaV/qqmi
en2cI2jJkROyRB4XI0N0GdubWbUz6wJZOQIxC0y8otX6rLDbgDZGMBgNNqDJZRgxYDUNGt2yeuD2
P3mfgm0cHNnBwEbGhzcYHcrLGtV1cFKqS/3hg29uZ/wNsxHGatbkyqIP+Gd2LKf44qnudxApE4ir
9Ew+qSe5qfju5krL64q7D0Y1f+hQE5iflKsx+1JVbq2XQAXlk572IDZOKus80sqwVjeh+jnGVK3l
eR3y3r2NvC10/cCcVemuUmGfBZMMTvQgJc2oP6oenziSiUpgvkC7PyWTdLNv4Q6TFhvy4FHicN5n
NUsiZwkwArWMdRawskc+8q0yzUiXrHemOpJ+jpwH6LM+k7ld86B8wZCbyNBneKyRy2TFzj0BzN44
EMhHCvOgFAX4XQ4VYwfsIobE1udoeMTUnxj+7nBkd0BdByGvACH6n9zFjxsWECVptmYVRJb8naNz
0jNyVm3I4O1ET6BdZ2BiwmVmHG4oCDH6D4AKrc/SxPgx4u1lnRipnOzZGBxdyzG2SzrqzS6EDH3Z
9izw1LnQcbMcBVOSkOJiDAt8nnXF26aIcQFIF3oB65tCdSQW8lUCEKFZpwqP4w3jkPtSLZueJz2b
pvlOYDLAyVxTUTIvJfK+mQCnYLxEk9RAs2dhW1k1mJI8G8HomURyH0OkJrwNZiyCrAPs9puJzsix
PtkdEb7+fe2WR8MTsQiUbLupyarU8jJNF1nZ9TPkoUPU3Jm2RQURkUwTBE00Ca3V54hUh6GRcs0v
Wyjo/O1/WXHtulp7Qspx3AOJdh+xUTePiqhTeAwDSMhG+liIBgvx924YvaFuQY6l6oOq7rnMI/6j
jYTL6OerMqWxsmAQLur+FdJuzJ04l4L6M7Vze2hoZYCBbWGlOSJEc3/qTRN5BLEIebZyZd9YBqTx
GKB6xO0t4ST/mRYCDUy4Yo3NlvbT09A0tFPBUBAmP7cezhE93Xlubw1wkHbA76OzNvbfo0yPQi5F
Eb1VWi9SRmqt5QK7R3aFKytm1iYj4T81yuJ/rBxa7sKmqhy7jyx0gzb1Oyw0PDYTywwFZWlf06b0
LfoMRbK1i0LjW5qbAGNLNJa4Ft0ijHRFZxngI0kc4Fa9RyJMG7++DjubxVoluYD9n/QfGUOOC0a8
433ZqjvHex5oFCj+CDBIaRUF7GId4UXshJ8V3Rk72ZMCrCY1vjAQvkloIdgThmh2ZYlRhs1MY/YR
kSeKe1SblPraTjLqTQEAfjwRSurAsVShoTi30tytEDBCUgCrNT4sJXnQxpw4Im3JnlDp++w64mx2
KdsazG6JrZFwGqAXlj8F/nMGDwABv6z0PLO2WFq4acXIL6KfJrDememfr6Dj6RIB8/8NTLKyqORC
P1vj6mCikfWzCg2sEWQs8ZC4k2u5qW43s22rjAPZrRrVx1Bkbwwm8zoyas651IYcb5vwO6CNm665
AhHl6FuQaGrf2ktVWq68kRQ0j3+CkKAmct/Fs3xAyzZa/h0kt7WUJDTBUzoCgoYJ2xYpTYfOL69j
rfrF3AqBSuvUtj2guD/3D+ZIiwik3ihFi+j3Xg4UuHw1eX/eHb+HZzuppMax/opIZJRjEtr5EuVy
m6/1qmOYOheqgxRwln7r0e2ZI4ljjOhVq/uW3PjBjHFfAwlKs82XKFADSUQVwDHf505UOVqnHftj
jDLjBWUXuEcoB29Bobz//OAk3r2PDDiVkAvGKVrFcPZVVcP8rAirRPyGpmix8I0tY5T86llqqHWg
zxB332Zvkmz/AfRC2LPS22OyqlFEq8qlCPZBFcW/xQk3ABW4bI3FuIJJiyuLA3K+ft4Qs2fnR7gu
A7AXdYwvEKETIc8gg5EUJ0m+YTLINAwzjnyqy9TiWu0ZC+fSOvt+5eO55Opzv4iBKF2CweynZYbn
NKAHrtDJVtOx6x2xiwpASomRClKLAHs97FhTQu2q6pZP6YtRWzW0+tRtUtzksQtRKnv6gaEzAbJ3
NT+jsJh/cBR2NEzJIRNvCO/RdoF6pLLfgQ/qvU9rK0fqL2HLMC7lbCRkELmnUnESR3TqA1yCI6qU
oW4HTaJkxHLBUsXa7iXqRmqUqsPc2TBd8EMH++KUmztUk1CXqz6pK5NFWhHrTyYe5XHukTDvO5Bh
4HSc0qwPnPAv5qn6mD29CC40fHFtqyqDUE3HTF66dAR1vLBdghUIXeLyLgNH2drF1mR+RmqzQTj6
0DmmJlUpBlRsJWgGYVGleL5cvy8KiI9+8PEIEHULIMep3/Ig8J/hDcYTqkQChv08TQtCcKgCCQ7a
4e2n21rwU6uf6Dk9dH1zeNGKDxcy4TJuFOkTY6IkVxlZQVgSrmUn6MVl4stn0QFi+LSLxsVkMtZX
zjLjaE4rtnQVT3xVxmOur4Pu1Jzgf/C9wFd6GN47ihqxqfEibIKczep+oAXB5SBxKjEwkNDv28q2
dEuKf6rGXsCGN/G7F1jjOn3bHAluYUco9kbiKSC5QbhGjbfZdzEZdke1ZTRR9FHW83pgaW+nc8vM
mVah4D1OcdaLG1o3EnS6w4uIE+Z0z2vfj7I+KWWZmarpPpE3YGYOz/mEM0wYLLRJfbinW3SUp3cb
aQrSqOTLExepT4ed4dZ7rLWYK9LiuyronkSAytzCU4R5t3ZznneEcGIYlo8LXDfEXzEq6twvpodm
aaZ5g9isJrOGnHqb34MRtANZb7KPnMPIKk5sE44EH7DRcRI8hCE27W/fJZaWEI9jFdfhg1xgn43f
zRKKpPaor5KFH8Kwb/XeQETuqEapXKloPSGjH03aFUKL/M/WmvDzZVLh/tbPdst1CcyyEpYyjTno
UfpntWT+h6gZexHBriltpT8r4j8sc1kKQHnxFFc62nEfjVB3Z0Tq63ny3788ogzKCRXdDPnrfPZB
gKw/KI/+jAUG0xjyDd/fJSy2a312QiOUozXTBJJwLQsBT1rgvS8P+NAWQSp/Nyye6ZpTJtF4tp6Q
qhb17NbLAdIERgttnV2cGDSfgoDvA34vfbNiyI5Rn/wnvKPA7XgIrbTjNfd1zo7dKDnXleDEQott
61qnUf4VSGtO3NeKZK6iKmT1IjvFOrS9exIP57sta/JKpRVEbG5ZgUwt0z1/eylkG3YhtZxwSeoH
IPvmQ+TQCjiu2zFnE86G4Z5RejW70pIILZOUKoaFtULqEMbgtYIcg6y4KcWi3fBaplErFV+kdcdA
3Md7mBzRijDT7L7w3zUqoYzvL/sBf4f8HpbFEdR9V3ZHzdHwUqsaR8NQRa9RNHIF+gDTnP/PPgnK
GjCICsn84OMtZuU2zuiyXmdD8P4F9eD2xEJBdjjPkVWtV2SrmRtORbmvlxgCqvue5ua9f8NMK6ZC
23P9TDmKm0nHPYctyQ4zTX+90HPQWH+GZnmBRhUWrjJIY1WZZAN6lo/tEMvLzpGP7VYzvOSe+Cyn
r5wFcqD+psENIaqY+fJPX+abuRoSBvyF3QQG4W95Of0dyzKmgs0YBLjywUSFlOr+NPR2JTdnmQQV
AQARmQAuJI5iuPDJXSkS+w4xN6d85D2JLkk0InWDCVF3jmS86vUTOKnPVO6uP3db/GMmA5HK+6Ym
MT0lO1ybZ0HQ0IPLys900MAC4frbEFb8/ypFYgVRXLbTSecE315H9YBSGyP9sWYxEb0rhKrjNaIV
gCKCbPvr0a13TbAoeU8cxHAesL4Htts/hUz8IWQ0MIRSFpfnPT1btkE7uFNMZi6XtUfMZrFQ11uv
5pmnBjZu4+BFlVmbxlR/3L3p2XU3YhGFXZTmhX7jR/VCPz++h8VEu5BRSfk4thJw7Eo83kMvsQ9I
H/P7ZNCCX2ryouZsweHCfOWj9Azh9gOQYwKPP8ANomZpn4MNc3FQ+tmp6ELGMXJ2o9A0dE4Qtc61
oMZH4t28P5DAHiWmFj6tVLRQX4a5nF6hNSNtabr7cgudkiOZSdYVtmECmG+xEK+hWFHpv1rP1nkd
AIRtmyaEzq1Fib1RgQ+qmS77pS+S3WW0W5Xgk+7CDjHpIIBK+iSdSbYFID6fAN5tjjajqyXnTpeX
/uDsTk3xL5Gmg6Mdb3fK9Aa773atHVZyDRR3kV0Km5VqTI0Cp1Ds0vE3uikO7ziX4TszC3AQq4RL
Cj9VxlQ0S+NIKWx/VF8oUMlVodGXatexUSozEKKHRguhw0I4H+x+zJiE/HULG/HcAJFIIx99z0F2
+aIVQy+0vEIuheP/crEAffUnyhufL+Pr0eFqyODY3aAIJb+5RBwWJe9wpj58BDj+C5vheA1ItB4n
ZHfqoQlu8H6L5LJ4+yLxbxmJO7Z+972Ur4YKbq3bq9zOFXrDUWV4OQJWCKEpXvRiQr3Jfa62ULZc
0AVEE7B2EYiql+9BghD8pkm1UjZexLCozNfE+zC9JpzPbjg0sm0yns0fStj6GvP+/ZRPtQm1mb2X
RcNyiNbkxxzBm9VRab7XakCCnVREzscxvuQdE/UNFaCvCKNINPL7xiUoTjhTlKvDlwV70jRZfjNJ
edHJosScWx/v5OcMArx/J304HgcBJkhJJsshYU6C7u01Z1lCF4Q/K8z9eluWquJCFGfr5kfhV17y
biv3ZBUF/1pkSIp3ow9nAKyv6sJcr0A4mAQk13awhKSzgyO7/7qHaUKCOPfQ9OZh/Y6JCNo00FOB
JgDzSzaiQ6JFs43VSZtM9vGqf3eHTh8tj9fzN950IsFprGqlIAKQD30XXPkmQ1kQonDuKK8c7dwL
AfHqjN2vITqg4Pi3Sb42TOkcgAgOkdP0hC8ImAWpcQpGKyBOaYjWrg4l83t2qj73jNe09ezgTDpP
tj37HqgI6ZrkNLy3DTp/V6J1V/+3dj5886chVRb/Bh8EQNWZuvGXsY6gXAbAOXKOtymN0psoBfBh
Kvj+dtv++lz+inrihe8cfV6nyJOLuaHqQPQ6qvbefgb67L/xmMeTHCRDAdJaA3mfYMp7PU/0vpqB
Xlr+SVIFTCmucmZI+elZm+9Y3GpZdeQJDvnHfF8AZfRLM6GKnc7IK5KYe69jBA3zGlVnqpe//Em/
L5zuAXflbwj+GSD4j10t24WtNh4tAX3Jd7GwiNBe0M/ryGkUyglyHAhTHHfAd1gGFcMh3ji1/lDr
w3UUN8EyL3WwsIswdhl9UsMyDgcKNG/e3KQydAknUoyx5IVIN/0PvHCa6kd1kQlVn+P4W8T37kLO
5gooM8AByuWy7Fmd7M5Bh2C0ivOAdC8pXDuqGhRHxDrooQGSYb80c/XbdDQC7czKpSGUQZoqDreC
aY+Z7ytc/TJXTkxXEx3fpA6JECcqOBY+lPCsvwCCXHebXRK1Wy7MCBDyjUkwBBYl5cPaSatr3FsR
xVQiTkofcYS8pQZ6AXq9hx78pxUKSPjX9rMa0RHZ9EbDCedswiocM8suMgMtx8o12ffaO4ImMdJW
8Eps9pmR5H3vHCEMHUO1YLzgxbUR1lVqKQ2QiGqq+B5H2lp/Fm4Ygn0NUwHOHOe/uAKfgXaF2eHr
2HcYS6lQfGW4MqwT8kBZ+gzqbbWPuecQ9d4MB/9SKxBzM1XrMheRkRloC3WVERrN2+6TesvnkIfX
K3l5Fe3Fx/Y86AuDfGKEd10EQ8eXFsFBIN8cvECzWzqfotSFfVyH4SjMQwPU7JhKlo4ggmTj0m5s
FtCK63yDVXMJSnkoHIAOMRCUYgHx4pcLYp1RIx9iamnadJ8QjRo8ElOuwxxiuutDKUyEuyqWnIEA
0Q2xwpZXe5KYpPDz8Rg89EROqsrSF8sL+w8qcdhISJH847/h4rqg+eHZdzkt6+TErkevcgaAcJUV
NeoQ+gQBlARSu9ugA5yoxWGZ8UxJ/bnIhYhk7HUKZy5lk1nF5AjdnsRii/pMN3c3aqnTBPzXAORI
hQb3OQk4sMvH9OQCWXnUK63LXz8Ult3V88faWfD5y3fJFOfOtHXtmHv8lxIarFCyRRwF6GEHY3SA
unSkTSGJ9i0/r0m0x4Q/WaGu4UGBnC9jbcpS9Qg+qaXsQfRoL+Bkh9vn0Wmm3HR2hTj2fIv0TuT7
xFUFVxRmNwAJrwwBD0G9Ax2EmKRBKlAx1XVoGNDkMdHUxOYwezUBp6i3hU+uKfItWPAZqvCy8CXY
DLfAcRJvaS07Upz02EU9XjU74plH72rY/NJ7XvETwl9XXI+kg6lUrhcJrT9x28vQBHdSTJ3ZVAxF
XfZy6urbX8FNSmCI1uqm+H6tLjiX3pdSpBQjhzeN2k189i4sUoqVep/6/2h7J6UdcE1NaKIYdmjj
2dNKKr/fqh5FVpsUuLhV4vNT+2WSsShbfGsu3Q3bRyryuxQZzuikKuRs4/v6AVtBClusB1SbbXQY
PGEMb7fFaGxhkeDtDvHG9yH6GEXKg418d1uRsfvlLpCBRPBnpVcCJSsNbyi14pANW4tyrrGTBNMM
e+iabTJ9LnWj/Fyk4jkFILvFDcGdG67Y+/Lsjb0Lt8Xago8T1/MPcpUmvLMWTfSkgfHUTmalkG/2
kSWLQHvgBkHzzW26iHgnnugRszKJcQRWU0iOMeyjcEsmQ1YTCjkjjgQE/LSIbMsk3goy6S2NSEDp
+veoz7TwW4rWNSUVRSY3YWW1yChiYGIzBxacruMFJ9a7AzmF6tIlKYxdOYQmEr3htO8gPql+U3IN
aFo0FojHTnCH5+WlHqe4Lda6RrNyIgTti8O0M9JU5z7H72xCGFQAx9gTj9QDOKIeilyrOppE6Gv2
yMQVO/PmWyoTBSOw7T/03qv5LSp+8B+CkGgTi69nqtN0P/MR/B8+qdoVLacXd+Yh01aecuewWLXq
9AtVyQAHFo5PHJaKGY3RoMO1HPAdeXoinKWb4PVhz4kzJ6bpeoWFmVJAkEpQ6IgDl34yQXKZBmGv
YSuaP70TRjWgJ8jKOvgkH5grblmcEDRGxUwIUOGxyYVZ7R6fIiH8esfvJyB4BxcdJucq9cAKCox9
wy5HLq668EMDldnVcz+keWnxw0ReMgu19ahkiGeZNfJ//q4BbIbyvB5fSr4fyalPHSO0YBCu6zF3
8SCBdoCtxb2kCqMiAvQjmJ0NzCP5VtDsJMBeUnS5P6vgAHM3+QhJork31I0xr/FQNKa98ceBZEl0
KLD1V8G29hrlHwv1ET7MMDkLTq2l8MW5W70LVFC769UBh78et1hnNIk/GRbXjoqkJG8TilaLf3DJ
06nkJ2ilv8XvFLirbK6MxgD5y9HWCFJZ13tOsrYjo7tBX+aGvYZJIsvrlyDoPGFe+UDlUTY16Sv+
b0RmtRc+QqqFHZlKumfapSRbmjG0triMtQMGQVHlHETd5zHSRq3BpQiBSNvetHli5KIAPXDa310G
fQ2Ds7hAgZhXZgclzPShUrxsOAzoZtLIehLLTjwGRputWLPNCyYHtuYwhuMf3NSw9vZV84xigoV1
qdSB1meNHppamjmWrJCkyQVkxe/PhKEXaxlyN7gmxLSOwPmtmAVchKLrpIys3wwPSEMt63gs3fnz
riDqBacTbhr8zOgVRe7P7ixg92OwKtTzHmUg7QMVsR5uhhQxyMxwLYfr9xGtdG1XuzxhmmNa9fT6
vNAcJGvPyCO79welzVnu4spf5+tGSzAtJIJbt06s459u6s8nvjtF4ex+66KAALoltT8ICne1wjNe
9YImW/vMso0bL7kwx8ntb4MaSsKMoZ2L5sObGkeZAxqVyxAUlGXu1nAY0u6jF672so4/d9k9MVJs
GqzHY1asx0b/52eeJfI9Aku7LpcmDA8yB++8cCzQWwH8lrZdkauzYHTWyrKon+IcUYC7m+oEd61A
FC4MyERaJ5wYcPDh9cMyReagnoSkjGc04WGjb/EicVq5ivhoj06HlV14EUyG09Z0XpbJop7+aFQv
GTR2ep5T86slKR/pkgvGaJDJDKERLgFK5EfcIcl+TIvajlG/OMPym8m7DHrHtwudfFEPx1iedRSB
mjiLnM7UjnFWslxvx7ykLK3xpY5GX56qDXAdAIDaalVNwNrhRx24I6eZMOME/WqCFLIYMNYnXnI9
OOg3+jJhi/pPx/8gwNiTWU1y9fiaA39WKoz1D/dsJl46DbJUlUFWldBzfCK2S5p6Lqk210aXBhxT
dYkevKNFx3jtc9hTBOtAzVvPK+kynUMOyLz0mxmcGI5dsQz7dHIxgI7mzqevWUOooKhJpLK9aB6o
UUgF1WfOFLEbUVoHq6CslzH/ACJZ+mCzXDp4eb4N30FgUl0qe7bggzkXF8mgWvRu1jHjrNa7aB5A
b+77EgRHdtgbNGoib7oP1Xd3Jg4XGBhxq5IXSV+HUtMH+l47Xymnp/+pU+iH6GevAIdeBZphuMit
tqZ1n4Nub9ZWOgW9+1HJBuP1VAtKrTC3RYCJ9ESkd6nAgznOSdaRSn+X5xN2JC3p/n8bnCwo0K2h
4lKvUENPoMNsTjD3FbB8x+OgqzBFoxNuw0iNalumrkIWkfmcbeVDEKm8x/gS6RfYV/gxs/AbxAh9
9dIlBzJNauyPHA8L2pg2HEZTdQLrFFl+oAuuezFcqg5Ec46ptjwOleOJ00gtxZ9oihXBSGF9bJ3L
lxMF0BRehHlaV5yeZ6fnduo+IHKEdkXr79l+hHVbisbUqXiF/TzeQPJY8HQYCECpGH7EeJCOyFfd
jMrp1SxfLOFExCLEW8+fUAXiuib+ydNATaz4gJGlZ838PEKPy3kG6tUbEPDyz1x9VoqHuE/IQPxc
yA2NWxFoUxKKpYuEs5G7bMnmWS3VQLhf78/nV4AsUxh1MlguAZnyMTiLD4o9TzeF5csa5KTXkznk
AquRTTIxCoI2MEiJfZx7noVUXxh1KAr1YLAh/igyMSAVC41BeETqQohTwkivgM24Uix4sllySF7M
yXDIB19f1Zk4bamDwoJxTy84PBAyl6h5c/XzQKz6MMF1TzRzThHJFpP2DcK29PZQUthYFm0rXREF
6XbyLEb+y53wMfEc/ofXSkhY5nE7/IXWalLkSEOkHFvEMghOFds8sVDPkpw990SSLqkkIrnjrmk2
rnMVJv7hLJPWefM/hVuv0kKwf9qbsq3xtFFdq6EghIezMwIsEU4W/Kg2gXkt44N/2NSWr2ZoxM+e
LyFTkf4TbY0wsPp85FS1z/eNhjE50dl+0sy/WGwxhWDJw+xrKku50U33+MqvhOhjBol53AVhF4AZ
firbgDKrYt+2FGvCsTE1kq7wJ+2P9Ixn759sx2fXLb/4SBJVNFeIYCx1bg5DsFesjPA7cQBJ2+PF
dbVhC3acS3t5w7dFWhtJoK3Mp2aMq1o928/p1qHZptnkBVfk2gTK6AhUSUvWBHy7U3YSfQJjOq04
OBvdEivQIvYYOxU0XT8WxhCw5ueBHasG+EmuhYXkBOIlmVI75FqoV0yz0Uk/1ODo+NSc0RkbQOlh
/pM7pe09MJV/I80xjy9fK5zdVXvrqRf5AiJLL4BON5Cy/LrguSxlRvo9NxLb9JTtt7JIWuyTpZF2
XfTTTm4lVsUOQVlloGYNkTDi5m72kGoWufcixtpSba7pxigH6a583ZqV/vpG/3ZemaLvZ6S9VrPC
lvM2qyb1dydc1rZlg83O9jEWoqcDWBSSF3KjhbajIq+MdoCJGJW2iYHcMPZSgSipTxyYCHFS+EA0
KHxfyBmN+7L0jm/vwk4QJV2AJWmdYfWMTBdUxoTGGBYu8hBye9IMjKh7GUCPewNGCXNZQ4sjwZFa
9Rqc2AKLAriyDBepnrw+b2ogNJ3eNaTkU7ZcIjz/yY6c7xEYSC+drJf78e5RNYaTGu4v0qLxwaMm
fLPaPvy4y7Mkh3F0Zk7ockhEiob0v/2b5WHyoLxgl6dBMnR/D6qxoJ14Iul9Tcd6FtVpDr9Vss1I
PG1xdMqY6SLI0pRdSixuWm5nomcHwjWA19OWZtao6KFDGWhLlDp18VRVMWIx1hgZ7piV6n/SWskN
u7jAyOo5kZpJbTQHSaE6LBfQM1mcQtxmbVBQypMlKvnXVNTYxdnAyE6y59a6+6OxRZuhTqCMqMXq
M4csAeOVRTe+ZxnioU9wCSvdCmD0TJ8USaC1lQdPMEtMD55kGO0gKuFCZyFFxdaRfpk2/tv67kT1
k1hVfJjVUolaMpobZmRIvOL4rEUDhX9Gnr9P79xXyZ7Pl+bKcqInWmwFIcWJ5RK4bR+7ZUyppdl1
qWTk//CUTkXpPGk/c+8MToUpeLBkNr/HQcJF/cnZfgRnXAzPcCySe9AzhuRCL6GU+GT6ma9Rsio8
HOJ+SsGYzN9NkTc4o4J2GVhSwtSXlJ68AdKt2LhWJ4w3jma7TJhhseqxq4VabEGRl1pMir+9c+cJ
dIv4rLhvKNKHEBqIQGKWxspKoiD7wzvsgLIwcLqAotnJWJeQ/wscCf7JdROwRNkBbBQBXg4PyJm7
3tNWs5l3gKDkiwqr4OkU9MhnzTSEgtSU5Re0my+qevXIH+U1DyB22A/CWYFOxJdZCL8AyXCarZsV
E3d52SD0XMCjpWbtIxAMqQ42CBc7f9Vi4OuwuAX8YYiFzhHa6++WbnzbDdR56L/gEcyToBshX6Tf
Jp9RkvItd2/+Flz/E8mEnSc3UlCbeC2U9D1klJ9yis3ikv//XincC7vjkPm4BSoqv0yTAxvJxQgD
jSwJcpvurKu7Xi6RC6e6CG5O08uw2UGO/GxbakhuoB068p4G4coS1zS/y1cVbo1MiELxWGe8kWF9
sbdTJAJNgVGRNPiVECBNQguZKrTNgge0IaNp9HQ6rs7hOmCMxSg97OPUE36ZZ2wZslofjxN5618V
5qxGDwQ4J9ujvhgMzo2BkD0O+/ONC1hm0tTlun6ol2DK5aghb2btBgmPDS6tlcYab3l+ksQ5WLtx
7TFdL3RRAhi3vBHMGvp52ZUY5z3fv3b3aEvUVnBtVjZqAHIQ7sP4B0inJrTTxmI80F6oDRm+v3MP
FiuGM54ocOQMiCMymeBg6hnB4PlfLEfHNPq0P43b3O/nNWhnnaWl2PguPaB/Z9NoZ42VVQ3TkAZx
id/mYc6EPJaMId2Wi4ihlSBtfsBKHLdTOB01Z/qIXpn4eAj8yshANH/5/pWmX/jDX2ZcxIWUKT20
4iDv2DazkV6utNdYj4IRW0dIqhmGQ/kcvhm/d58jeTxhWYAJIJ9j3SvYsgONgYe7GOU1pcIDFaDF
/4iLGESsNnjYiCoVp5D/dCiYtal5dZKBj+6tHkRL/+v6eiv0Z7Nm16ZXEK3/vQXqihDUb2Wpg3L/
BVryxHBFpUbc8uX9yMZwiLtIIPukXwqwXN5dmovPvtYZGnDsBlv17rcui6wNXe594DKKE5YTaX7K
yWzUPSQscPqtgUp3Pg1wCCHis2pVQMfVpl3QYmJhGSMwENIfqmLvoydxmtowdhm6rrO0wnqjrKGT
VOMB8R327sEjF1ifzCEg9mXNNk8DfVM997UYnz7y65E3IRysU+w5Ul8wrR59NULMyVfIkc6eMtiQ
1h+5rFY2s6qoIGchjJoASXDvNpRmR2lpKNtbcxYUhIoA4wyhKR4Z6TePKw6LVJZZnfN/Jf0wKGLJ
VFhwj4nrMuryTO7MSwjz3RKbdAquQcNCzk2DvJF2Mph/7wbY6KFAWIzAMUXN4iYGLj3MhXwS3Dt6
IvSySjnxfzcyALw60sQoCwr2TvMJam4LDVNgYNBZJt1ZUAnkYfZJeAGPMRUkDWRI4iz7YzCfLSIu
k4Rf52VKWSHmsN+nWCz1WC6WzqiqRGt7Aj5ezoe9wHoE04MnxU1/xQOZMdayit2oqQ6X9vzk5M1h
wP2nxhlneAB4eNCuj+Bz378lckJJWTdW0PV6obvlT9WaoEYjtHhtDSBtE++tCoYRAyXh6BU2mi2l
+UP5V1AO708HVqWWRLMGw8gPOceiWil/sdpKk52WGCLzyrjMKdEhLHs0dccJ3CdoyoH/Ba7DUX0u
yCQ++pxpTKTLkCwABVZS4sPHN10gLhYkDqE8qtHj/tb9FiOlVXWmlK6J3cf2GmWE78OUOgWatZD9
+A4XvtiOyidCgomq8g9uopgwFRfHq+p0TEGKtaKWv258544C3tzijnru3zHQ6kNQimVIZe8k1Df7
xxZP3q/xWmk/SYvNizPy32V0SP4CFHToSUHw4fKQoyUnwPh754HmAKO1Tk1Hm8k/K/EgSfJGSE9W
LsGmjqIrxup/I60xRB1BTcVf9qVgoCYOxj0tgicx9N7eH+YZpX+YD+4JrLFPwQQBmsVELbS7p6dU
CC1OreMGQbmle0cVPj/2sekw30K9db6vFhrmWE9aOQVt1M52xBq2hUaKP6dJr0lJLACqmNSbJ9d5
SaJEDLNBPzhgDmQqf3mm7xZu2rU6zVp4F70OULGmf/PpiOa7IJnZWThQg5K9sNbuH+cf/Ct/7aGM
NjzjqeFjHYQTcXDP/8mHKDdi9AkMj2f8FcIaJ4YPK9K8SXzewiBW4mJrTw7vOwhqX24e6T6wVMl4
vV7bUhRhhG7Y9iZ1v1VaX+qknM2XAfqO4S+S2GpPPA9iZ9umdjiqCqL7PlcM9+F7dKw5MFb8W0r8
pB18nlJZojxejSvCUTypAwCftNF9eUF00bqjbKdTACH3TvDzGt3sca89sEDEdtCsb72x4qxI6W48
pikfxEUh3pZLWtilKTKkcnXg+0xOsykQNCCXraO6Mp4zvOHyl2rnkff0VWoj/ftfa1jfegDVTY7i
8yCPWD46NXroorQgN7qjrrPChixRNUsls9OpQgEDbxJeFPcwzC4QId49oUtduy/o1hUYYtU43JnX
mrVyo9lu3mfhQL7sDAO5f1Rdhogya9pwM1Z4dVywN8TsI7hCLjDi1QatyIivX2Cm2UxEAhdi6qPn
xKu7gLWD9bDzETu/4+u304isrsN5+ynDndOu3qAmDVQzbgjjUMqCEXgV1tGQRM3gvRkxn5zJyNAy
BceaWaL97rRqX1xnSqhEuahULuv4vxcvKnKsXwck2+PybmNJAGwH/ixKCa+Y4WWFn0SzUZaLxEaC
qoP57gVR0eVENvtuofX8f72lgbWwjnoKvjuSEIsA2zg+80L7t+rhANscSPu/BY4nkA08X+7Fl0vK
uNTSbmAGXsg7PRkj0UNrnZTmdNU9sZgHxppYG7cvyXOpBe3ZzBMWofixPl1W93hUOcnGUyTmbkOz
/lPS7UjB7MAh0YmPxeYAFuQQIzMA5KK4nGXq17CDWZknSbCe/ntkrPJjqKj5s29wfVOdtA07ubNU
Ke37ksdMjmhrB1ljD2roBwufXHPDHP7XztJzdHhJjC9mwTtOEiEx5S/tvf+l3XcX2MAq7S1CNNyA
lBoI6hX2CsEs7TU/g7wj+Rq9V61O69yduNja/CBW6E50n5fStywxQ1W3yXNXgwPshGc0P7ewdW8M
6MSkocOo+CZPi5fqkXeButVogh0mu1njkAEG+YHjSMWuZq5XGUL0sA+P/2jcPB7e/mCIXqWx/m7K
TA2YAymaKtERszI1UWvnTX2+mofW10kGgz1rwDAj12IUtoJseLd3hLqSFGZfHEZMyPJIHobwqg/N
4au+gJHRzHtkJ/c+V1xRmTEiLuRqtD32NhjS4Lhp/5JM+UjGHDZM8zQU2kw0HRc58qgE+QPwoX1Z
OU4I0zyOwxpDkrrN6Q/DrjBDqldg+PBCKwAJ4FRQGg0DOkazYchZpeYYOQxBDTYTzFeU/s2ANOG+
u/0yIS8n8IblAXWUSg/rU7txd4ZosYGMwul1FNyJbDhrpwh8IRM4l4AMx62CRXuhEz1yAh6/psu2
Q6qvfwdR/ayWGnOX6x9Cbe8hAxHg5B9uJvpJcBxzdJ+nad1VIxhzv3q7ue1TAELp58Ebia4dLjDm
SKBYzpC1l7rEK9RNNfe5RRQ7AVAVRQmado+eeYTIK39R1ydDAbe2O7uDmDFd+a4eK4fQ3k+N7Vz9
Z9fUlDIY8qsRdJkcn2i19be25AugoTCVB7lfh7W5Jo1bsNacOF+FsOkgE2rYYz9c+0YivTqTFOgx
FMxWLcBBOVGTpU6fPzNhoYfpUk8PmPmnMB+2aqmONbwO3rRZ0Ah1j1f7lca51CkrFvU1HatbzSFj
OQlCaQE/W84MaLRAKvR92hhSrnHjmGLb9CqGG29H1ynXC0WHA8RL8w5kJWzyOLrRnnWNbWcLOAIa
03EkgsBhi3sqtLrOUSSfhG86TzET0RbUPB09SZspeKcCJLNAR+3HYHGipSO43nklL4HvnITrNVmF
bIQC0wTTvmUsi9qMuP/x1sm50f7U11y7uvP+EmylSxYvfKvZ0qn8d68mBuiqkrP0ihKEyjqDLkz2
lpx+ZfaDktNZJumxMjQeopRM3q2PraZ9+eNaptq5pE4N53kLXzkqoPl7kvTYytQQgvJRSIx+hURJ
c+bIhPOBIhnJFwr8Gt05ni7QH3RnemeIokuvyQzVFEcjJL1qR2DkqXiQywi7aP+9slReBJd9rtkd
/V+QGWaBaA+WdMQLMgSkYwCb0qCNsNGps1mhqw7HhX0paGXEVRW4yg3zmiBYVT26Ewqyrw32fclc
F/kplvFLdvV1Xfnr4opRbnmLDsDhYSIfAGWABKsO3cIiokkRa8jX7+INRojHGY0s9FoYmxz7FYHJ
7wUx47BuFQJzmUDr5Hlb16OF3fpwRdG0iWgCqyB4axmPNhEpKyu9PGmiiyzy7pVvScdvWjkibCy5
rU/WodtOtZZi94gNb4WIdtpIVUYT88dx/O+rha1QBxdhbGjq+eVAzluvdRLvfErsCg4y0/pJlcHE
RX4ApSLr1mf5ODj8gwksQL22biLdhVq0N82f8hVZLZJm8cEM5Tbx0N5KoE0lLHRV+LS49hM9gV4W
lOzltu3DGrkoIGB9mlCsKJTMA1h04zHAosWJB3O2VEQZP7+G+jv2AGu7mjLqyuMiywXbbwlTpllB
1VGauQpqih2JcjYlEHONtOZjJctwrNQiVR58corrO/5DVxVKNT3l1Z/Ce8PNrXKsyWgyx6OLqlNh
ak8oxjkAAlSj581Yp0sghrUkSCZ5T8EZlq/19BJt8QodlzdLoom2CkMEOqkv89q58aMBHxoCuNE5
2wvvpbChhAWCE+pP2Gq63O4n5emhU8U8Mz/ChXCfC5TCBbQEWXCH6Gy9N38SJQnH6qjsKselNz0e
vAEqvERavaZrO5OczNAKpnHNgV9ly669spkyuD1yRidqhtfXYLb80N7pRGJR2XWbXLjvklUbeDh7
KlmrjSup5loK6VNvatt658mtSv/eH8ACgYb/F1M2uyu5S3SfPFkIB5OjI8A6alhe4gAQMtPrC5Ds
rfNzAE5+jzFpEHLhmQki0Yc8SFgpA2wkg9+Xlq96ObUS5F36ocjYAAk4KAQKRoRy4NmNga5gKkcc
g8+Z1YqEALmYkaYau5Yzg8Kb0G8Bc7Af3denp3gCTC3fJ4/1kWOcEr9l1YzNQqQhc4GSVQWc090W
MXfkyHrl4RSf0rXlc69rZkUJm2DdPuP+QtbZ2myu20YgSzDEXXQSAomIuQlwjNT/ujT0NOdezxCI
O4sEQuueuSrnfa+rjxcezmRe/MTaaqiGPcLGWELHX1eqNsox4lH4Mu/j40+t5U2o3/k4anlW61T4
ebV0hfBOychYE1wdCDek3vKiW9Z55fWVw7s40xco9ZVnKq+ZXDWGt96dZ+Bpze6f/jWPsWEOhxXe
wHxKkp47XnqhdmqQRaNXYUAoIrmbjBqVrzPdRCc+rHH1cY69JyLWKynNF3KHWF01tR6KYKn2ERPZ
6Qv3kNKpDowo6NWCdkEOAQdNBtfydJl90Ckt3wWzhbycwVTFYg+P8fBKTruDWRNKxI2eBeYvA4D/
Qb1lzpbncjeqbjdyTRtgNY4XxqUn+mMIaTQzfy0WBsD70Ry3DPt42KsKDBwYdM9cnqUg5ZWMW0tv
FNmEiMPaHvXH3uyEsmvPnr/T2aSHCxHvli5TgMIbMZWb5UPh1R8FdK6Vk5SNbhQs/sF1ACES0ngx
gxihYGY7VLunqeHNQyqe2SxAPrbLFVBosVhMg0IO0Oc7GUmKSXx/iIVHGPOEVADG48AWrMFsbNIh
JH1gqAwqn5jFwbImAb6Y5V5fL2cufkmsEPgjkS3z0qzAZ41ODB1zNCqKQ7PTc/v6lJouV1ljDV+L
ZxYK9oGr7D/2pkVacF78pSSSZNy0VRulBYWA1ZMhFyLLnetE7tK/gUMM/76K6ZkzFEjIjuPrKV3u
gTK3l/ZlEWh9YnlmpdXWA561hzZTIvsm98Mq6rtmpllN64z4SZi4Re9JMFsua+Vor7R/Mc4vhGx6
p2Bv5usfzKJY8ZrKsG4XzEsyesRmYzZWDMgw7WR+jQEuZjzJx68utb/mSzNF19T3iPPLJz127sF6
EruWDRP9CWrKlCWlu4IxtAOsjsPH9egQu0kDpv/TJhBoatWNcKdDtXsI3fz4JkRGRLXO0YEWmZLw
pPJj2eiITsZnVv/01WJ7KriXVjtsA3GfaaTjTdw8kVLgMA/dFE/5Ks/QccXEkWpS8x9fr/7r92kX
aOOylwvwLWIiJNlgZ9uLTtNJpsqztTIu5Pnk+8JzbktXWEUNLvyp8EpQpJJBX00BYD7QxHL18MNu
AYkcH3L8fwDE2nvlbY/W4gbttRWUCBsCaueFvAyO7MxTYMVlT9PQGsFXSpkMksiRbfjTTc7GCOtG
gEWt3xrMOCCCpB7SQRWcq6BTpG9oHRgXgmrVc+DSrSsWPrHfrLLF6D0VoaVT9BRsOEO53uacszbh
1PO8nsMKJ+FriCw3f0/rvKifZEpotm4lViprA/Juqhq2aUkGVWubdalW8C/rDeC+O0ERmPLCm7jN
qmmK2cp18DxlnFfvjozo2hfglF7I2rmRmt7Z/+hzb/S9yYDNf9tXVWDxmJ32pHdW3LU2dT8a5AIC
pzfjbkmeeYahTMJ/4HO9Wqxbe+yy8UjomeDNT052zr3c/HMXYelA3+Z85Na5GnWJ54+EdVFAt5dI
HlPGokO7IbbfYCXkSf8eH0+Zrp0AnVJPnCVRYrlD7AurZ2FBZc00rdNi3/gKyEfI8tmY2CFWjIRC
odBfOjLaxN7eLL+NwEn+A958WkAMeh1LwGX56I237p4knil0JkpkISFpgGeXdqpu/ipZW6sXt2PO
vDMHkuZuHqAckAwNho2T95DUMwozRo084VBkB7YF2trayKuwGbm3NKgrpHemr5yAb2ef8sUw15SF
c8VAzyxiypP3Yd/9iHbROaWqUcId4BiwVp41D2LtH/TuS3ILyAlCKXF1VE0lfqi/5aQtUNWAL24U
S8UJnBOySr6+N6WuwZRUlkFIyHeoZJLAmpEX4BR0eKi1Wy3g7SdLBMHCMpeS81AW8jJNL8X43+BN
YbOxtiJu2BHkhPlqxbfkq4f67dsfVQp0Ebmw0vOS9P8jq6St4YQvhgOgXA12pSB6oRL4FsUa5cS4
7XPE/M0L96murJ+dpcafCU4R6gigsxk8OVpb4t6cbJzOMjUQXXaVqrf6vBJaDpzscOgvqJ7kdoHy
jvClwY/hWW6LuaXMiCEd6oqNeRL1exfXe8nHQs4wb6Ux1zXRQcxCSCxWt3+BxR/f5PvNa/BuzJka
SaGneR2gMI33uF8JOAeSjZCiGmCJ5NoG4IYMqjfdZlfytffgcRJ4LDNHEuAmvt/SRo60wAd9Ao8c
bBAIlrxk8PAyC3gShAwNXATkc0KKONrJ+yerTv3TnuX9qvD2ZVMSrowoLoCHVoBCe5oYhdejTe2i
VSHsqbpGqPKwNRJ3zNkC6AZnYd3HQnV21BnQ+AzoNdwgqbDhthSnj+nbtVPiWyxi1yz8LM+X2lfw
aRfcxUcYjFWaB8HQSDODHnA21L6y8nDbMPu5+aDkxy8x3zd8v7beXU8SQ6i4OTDfVHo6LlLPWLdx
U2+okt3EdBdujjUNCJTkf7FOS92CLa+OdeL1xyg3ElnyzIaNHrcR5mQjWTrVX+fIPjRPYOzD4V/B
yFXOtrMspefOe1imvaq+UZmob0o7LnDFxsj16asNIej8aXkwdHNCWqQZxXX7p8e0Qbbc8IYd3gm3
igHFqSc8JUUZKz2jyIaCB1K2z73Endh8EnrpoEAWV6poRo29SAmHDRZT5HavRRnH2BnJBhqZNXFP
tKnVrTfNogApYyobOrBIqE3XNnI2Sy2LF+Ip6zAPV3pG7jV+oxa9HFuzufy6oi7mEKmQtAu2UJW0
drfslovdAwMGm9knKV0XSw5aQsfvDfhPHoTwB5ReSoGlxBisXZAoV7xdlZY/8ElBDZGPZlts6/+R
qhpenx2hCaxuSfX9vWsIAjkO17NIa2iSICqXpVTdA1wMPoEZ7fBYcveO6Ht3Kl5i6bWDn9qylRzc
M5zXcy2GuN4Mh2hmuamDdDOy+i2g5xCs31W4SabjYGoNB9DDI0j9DpaePWSWEtFAI64n5tC+YLHH
3oGyNJJzc7sUF+2xaMrQNd88FG3iCQuRKYH8Mr5EyEKpeN2Rm3N1qyMfaPx/sUzuga/pgNZOqGDz
P82LRneG0pQiU4cab/RZejSJd7xgRGOTqBzank7yG46vN8vOSTFpZUVoCpIxkiGbWUZOUHNKYRly
51rTUtGVCrhgpwqFweIxSqoM4vYKKQRvwxovPycmZYZdd9yCHUCP0VTMZtXEXTpPtvGDXBu33680
rWRwHESlEUIBcyH2ZSf+tbFcw+D/sTLSFxXp8iD6XBkMQoDbIhBONbU71d9w73gkyJubhNw4oQ+2
aHaxxfRghce8LnvG2PnWAh4yB0sF3V4jcRPlusGZN7Z9V0J9bIZZJHwJKacYAQQUnTtlTjgKjWAD
E4kChAwUY4J+VyGuQGMnvI1E7dGLeMYz6KzC2TJEYUcouD0rkJ0a3Uc06hZE5OyJjshrV+2hOdqY
WTYfm8lZZFHm3Qsiz8WewIejY9ULLcQP8iszi+Y9t/aYybzJUnumvEvEHVKVdHDt6Mt+ixN/raDS
XOljF85GkER+HGhECbch20enTtgcRJip8duawjjgvwhrnewWt6oAmBMj2zl6b7REVhrjKX7YCKjF
KGQwblGUobj3yyK8YfZp3x9WXyRY1Jcp/NpsBHdDMnKYaSxGSLN2ZnJsRLU1GtZBIhQhHGzY9z5w
KnlVXz1UFblTyFTvacqbVmSJmYR4Cnd5AtV/n1+f3piwon0L8myEkNX7nsJ2n+p5i4G/k7tJ1rwE
Dom3ts6DrZvFAoYjrvTGAOPix6LM8b+ps8VnbmeB/5K/8yxmDFF9650aRtSQWtKiw0lktxnMm/7a
1yyTlRWgdtyYYpiU3rbSuqYwc4blzbH7j2oH43S6Y27eaLbqxrkMffxdkLe/ehf1IWI7R54h06Ir
yTPRT/YNdYW6nTOfX7pLHBVIsBpZ3qMI0DX+4FaqESIa7vAa9F19hWFBo3AoCajeH1HwuQFUaj1h
8FYC8q0GKHDBSQ6RisFSgdQRvQVXZul6vaDLWxFs0iuR5o8m2c8Ksv1Dqp1pqan7r3QbpvQ5eSnl
CtiuBPbUvAcHAdwr57vgSexN8zY/eKKi9Dalt6gBrloYR3Kzga8ImXwpZklNgVSkOGtPey3eyovz
pAR2WN52VkiFglquPC1xoWiwa+Lr17FMJcJ8WFVtVUoFgbp0P35zT54DvWVE95nIdx36b/6i62Lo
Mf8zS506eYJNp7F/bFrHa221VQr+fxQTUzMDN7W3+Jd+yGNHPWECuK92drkSRtjOj9MKd3oK3ENn
GtQLHVSvX8DusUrSipLp9fUhlrjTnKAG1iaCcfpceHSQlo0So8lvj/edAV6JF+9KMqFq0wWOLi7R
PuCMSuXu/DZ6/b+x+f4hgiitx+De20A7x2vcOFv8p+GpHn8Ta35/BL4BWuiH4z/4wJHJlCkS9Hqp
2n94kIk4jMfN+98YPN7GUj8mzJIpdsoHfjIwGDjBYnpD5VzfPvxfEpn1U8hO9jPKP2Kdyk4jFmGl
LZlgbICJfirgz+262CGyGSBvhChoYJqwrOlcfhYD13jzrFgRZt0YSeDbxOI3wnwOxl41GD9pg8Lc
DVUqCHmcErBaG1NXYOZsSYbDuDF4e32+QANuaJGokh8yO3VDPUb39WGVEY0tlddo6Mv++lSJ9eLX
rS2i6OY7YTZsQ9KGCiYudCmNTyaD1jj6xQpCUJmDPvYTBzJZr1EE3gInL0Z/T4MTZD9cDHYutDoX
kkhF1FGUaWUoJYI3ISUiBUCMXzA1xyxJwdWoc9caDUHj0tLNogE+dxLLkspgmf5AzO+wswjcXalq
5R67fQDtoJmJ2lR+MQaKWmLvnlAIaZi+GRY/vyrHpvngfwXiJNjtCDzA6RTO9qy0u8nyxm97u/9/
TBU1pKilL/1X+tqR6MFjg+4hFqSBRzkjZNuX1RXYvjqS8emSrDRSK7dM3L3S42Con48dWcCEKX8O
Samzt4+K3GOrTkdKY0iSg+zICrPBX0kFoI5JSuj8NXkKEKcdOoQrTpAqZllvZhhVDKzb2/MrSYQi
0WjeDHA/B4uJHM+B/BRnqIfjJ4UvP28W618yNOj2fxJdleUD70RI5t8X1Ye3vU6kGbgKHx2edoAF
bXTliu7Xv+QdPwjrnFfAuLtMNB19pz5HdkOjG2JvPCODdKgJ2Sz3b0vj+PqIlTaSIGekN2PVy2Xc
ECYz74/hdLdkh44wSCBzRn50Yae7hSaKzE93FH5remUg1iOnGU7ViWhqR0Eyu8k4KIGMQc4KlcU/
8GMZiuNEIEP0qZPG56momYTWsF9VSU8tAdNivLDw8HGD9i5mr/9YBnXgxBAhJSUBZMzOcoKcB+/+
AtCxUa9XxU237kDFh/gdyBaKTmNMwJo2eMAjJId80whlEvHwKbPXIoX3mzespbLItooMxxvzWkRG
trdYNota1VFeqjk43TshnmN0BDPiAlK4zEB2fs20VIBTBUwuCJqO9XFHzR1JBHRBUCpp9N2Jb85y
VxsumhWA8Ir0mQ6krzDlBMtWf6xL117FuFBaOSLlfXZaAlrQAed9yo+sv+OlI/zhFZKipO5IgCfy
JV/MUzfv9wEdV3ppCo3KOighV6+L9pZqB6LOw0XQgW3p5pN962BFihJUAfWnOF6GUHCjy61O31LD
eCrT9vRKY6UP/6i5OKjiRdYNr25rZb2bEcgZbSJg0dFvBxAi1LDz2u7KCj5ewlKnXmxD2Xl4hbgS
rNYiKsZKNQHDKPEJRJsJOew+mO1hY3dvfTXM+t1ayTc/XN/YTTrpiWyy3yJT83Dttnrw3Km8xOfK
aNoSQP5jf7ooICkCtkZYeZivJFoNKb+7r+mSkvYULeoW5SkWqJ5zpJncW0cZ8PaoTIIgIyX9cbGG
dcSOu/VJhU+2wQOVp3SnBaB3yFkepbwxbtXGpzGiQwZBSeLkLss85duWQA1X3wSQdLly2ymh7pkp
n6/dUaq12iHr7xSJC1n7+v5JvjtZJfwKSFqOA4EJ3Ufs/4mvVJohLyYIqvPe3LnoL+X+oBFn5o59
tv9/tE7UwXrqRpTdzq6Lw4kr4eQHo7/HQXS3xOulDqCDX0uv00tctkJ0zyP8EzjCmI6viPidSzjQ
7jxraPhQtgAEa60bj1Ngq0jvJ8vmH+iAccEfTzREUsdjIIxLi/sOYhWAZi9BRZCS6a+5t3Km1WY2
vUh6KP9qGJoyqBnLvd1xA100XCdF4jQLI/juXfaxrWbBKoTUnpctK20jjXrVC6oCse6VWB1n1WKg
NzsgKDZaJUpnsJjdAsGMK8OgrDNONHAUXgbBVipJjFKWsIw44Oh6uoxfoNWp7Id/2DgNACSGmGGL
NoK+vbbkZLvmxLZMXmyV8Pw3np1c4/Kyoc5imUSHyXo9KpTllWwQuQCHwUBNUOwlh7xEMtxFU88o
y4O0CZGN2qbVKFDXNm32wP3kOjOJkGGrESsJdiJFnGasjfoyg+cPEas0ezX/YncbVKuAsmxvlZ/+
Z65GXSTkSxWHGw+9I7shEOVu6P0Znn2Jq6KxKeb8XJFMndfAPtBHapA1x16d3Lt0p+A1huU8gLH4
DiTeTXmw+dWY2xuB7MZrkqOBW5t5Wc+7X29XAyQO+xCgQ+K9SQ22iz//orDWF/2BpQlPduALPU5O
I4WnZQQ/O+dp108X+cgZtgva33wJ/8JahSqF37guwMlcKvfWQzlCnUaEwYqGvT/dMSaY94l/5NMh
O+0pjqyA9UCkbQtr6bn0y4BP1nFN+1zJ8LZU3MetTjgUo0L1PVyBT/QG1K0fja38z3yUfNRp7agW
QifiI4UhP4dac3EixYO670SBAL82XjnW4/JGGkrGy4GvR6QscBcNikdZYUA1taQwUuYy2ShmII2L
rHXxTVRSqCmxem/1zyyWvGYWxT/nbL3Jb2l5cVpsCMsOunym+e/rWxt8xunzTJpzCQ6419rFWm8j
oDj1mS18n7wbS9vELCKLoYDiYh2WUxWBLZSal58cvb2Hj2GD7x7N1iVXGVbsXVz6emU7Kpg1D0lI
2blhkKJONE/HhKcMfeh+7apaYIBjvwFI3vGlSgi4gTdJ4DqSXuDxwG4FPWuN0b+pIWopf1uajbTt
Xrd2HiFupNdK1l/FgbO5bTqpLwi77mCewEMiHRtoqJ/iRBKKklbkMHF2YDyHlFksbykZG0oAi7Qp
j6LEpH4i97LVnsVkb83u+TNvpR5ehFHh8M0AIioaBj8gaQ19xr9m4nU+UNHsJ++4nnGT0l/7Ajjp
C5Sppm7KZsnQbkqJqK0K6ubNJxmw6SHH0gzIGGG+XXZ5Tc44g8tQBuSFS9j095HKlNVZm0UHSN2p
LL5GBEHswpJ5uDNVlf+cjYZlTOuf9nOQ1GpboksJy6pnBkGmK1CgXyn8btagc+ZHf8wxhmuRk34I
lINYWJP1RYATGIT4jSPWoos5qtGvfaP/pF+bpZl43SPXeINvbfVV2QwVpEVQtys/EW6q5Oij4w41
UJq+DGCbGQOXB+GA1bhQW5AB0GUAZxMOecZue5y6fNkqz/NzPl6JfF4Hh6FAAMHwtaiyirkvd4un
skmZa/q4/+I6UCghpAi8rJBUYC729IWLOG/BH78uWC1D3xBAf/l8gUfjk5O4QTQTmx9C/aZIGKH7
vzIW7Obrsp36FnXarhKgkPcXjDi9lYgnT1J4ygEudof3oXBM4BpJGHsdNeWAfDNZ0jCc9hnLUiif
DEMuvcS0Y7mywwf5pyrfo2DPA8+4/q0MV87b7pGdB/cnRJwEthCyST/cZZkoFbF//Fh17tzDYXE1
JM6tP2grAoHzBEYr7Cp/xIy9HQ+dZc/hEZ7KBknIHBUC0ogUX5BmKuoreFZxazDMNMfkr8XjuRmz
fdIBXIDGT1TedpJSi7uGqTdV+jSZ5OOm4W1cgj7WUbKGdTdi2NgYI3igl0dDRz51lK5M4bJWxfHS
nGr89jVM5KumNGCI6OaMbdxCvBntWhi1kK46ldvMInsndXqi9aavtGCvsFJBXI2DUW7zgoJKqLv2
Y4sioIirquovCPuYd9ErM6B4wkO5Ep6YpZ5ax5jFZY7i+jHO6FNKQc1TVQgEAr1UI2ePL7ZYtROd
fk6AIi7ABu0xKJPpnhBOR9M4lA5rcfhgKfT548pCr92Pj/Pv/BLPoQc6wQblAaVQjYcVmau+7iE0
IKLE0haGhWw4WVCMkDbNoiHsrfp7RCHyAsSmcnfZt2VazfnoWQ5eJmL+tRHvMq3K2IVMTwnm7Fs5
e7EOvziokzOUC5GRsPwvYXgn4u9kVAXKoG93tVL3R8eD5OLby9Q39AnEWnaANJBU1kiEitjnyHp6
jeYJvg6zPtTBOpfWPH/lPyfTUUWRC+aKfDl1BYfPHHSUE2O75G88/Leyygk0fNOcHL/4hAeiGU0K
F0KyLtGGN0AOyJZ+4J2IAZOXAp9t0Gb7KfLtBV3HNNCF/6rfLt3S67KTJ/ZJw/I1gLEH5VaqI69r
AowJN5nTEyouDdzFa+9hG7PVyySgS7AyhWr7E24om6X0JPteQOknZwBplhlvxSk7wlYVWZQf9Gn2
JTqJYqyGv3duigv4zPxGf435l38YOR9bk5uqmuBIQGjVtrnN9zKLCnodBmqqZ+o5Ex+ADKavieHS
W7oreAujGK0CgslIBywL1pVRAgctHqsZy9g80uPkOmKQE91Z2kfc3osJV8z0q6AzjcFALgShL3+w
1tU5u9Z6hwAAaeJPV6YjuVXi3hPHowsTmQzVfl1OQ22yqkYRq/3hZ0AGR59TgT/R2SgF7wgD9Mxf
Osv1vGHX46LU+fjyB7SkL3QYme2J1XVZjozzj3RnwenHu93zLUuOuypRQaEGLyI2AtI//Y4YaNwf
3I4B5TrSCRD06KVuh28rzl28SEDvJHk28WYsTUniuey4R995ZEvjQhUqEi0p5k5s4es4YHAgKcqz
Fc3AMs9vIPxzQMjeuC3h7QLkI44zqX5WdjhSs5lNZ9p6gcKzB391K6MDTnBS0oyhUf7ni4lT/t20
GVhYuxXbtIwiXPE+h7sJ0oZmV4rWiRRLBhif2f6h0x5twnR9auvWcokpBtR6WXm640IJvSlHBkwo
yKuN/R6/N2JyVcLlcZWQoKvZvpVWZuGo51VO6t5tyk85AH0iTrlxnoJGLWblrOvfm2cylOZKue1A
7goYRaYQz4txpLZHiD70i7VP54n/3TT/Qx6yaAUNubmQ0uJl3+/+UwDIFuTG3Bu9dR+rnO8K+Igv
bSPoxcsO5TP0Mc33IH6RjYCVJEmBON0fgpA7CYqbcAENoJ0UULLwSEAnFL647yKeCK9iHezw+p5Q
1Brgz3lMIrTpQGJm+yc3NtQf9U80Z69Q05iBJRdTgX9Ss6vpNSD+pga+6bX+MPOqV6MtgtQzd10y
UNaq84ryNFRoaSAhsvtjxCK7w19IFHHmQaTk/+cPV15cokRqwJepMeTqfKaSNotDDj2VUCJFextU
nzLCiA4pqnGtLECJp0GVk2Q2qHp77AHfYjNXeXd1ZSAFOj+0fgA1ioUUS3Q6g1dcOnmMzY0D/evJ
maKFpQ0ix7AIb37JcZFo6m5JmXtOp7larutXgeOT1/GClF+uROoEOYCRm/cQtcR3U2y0TYXKC20Y
LHkKQP+Bp7p/jZ+4+199l8q4fnUvCdUB1C+X6PKTjIHLP0ThMM/iozcbBCDpFcRaCNBCEQBvsnfV
PgqKITAm5qmjtP2d6PA1JPouod5ZbmPLJZGqu2mAN1F4qndJJdke5S8w/ruGU3aQrNn+rDL+FSW/
3lLJCgrtAyYcBVtq2xx8h4bHaj9BXXv+OuyZZrVtsyhkINItblDon+hHJYgZMjrG5oqVgh3FIf1I
XHIWaQIf7C+6779ax5nHBK/cAvD8R+7+AWtCVq/wHjk6lT7SCuyuXpDzp/jA0jO8qHYGDW1ua1t+
lN/8dWxfp5OCvVLYJQLLJiTLvXSXppQevIgGzAXTIFwrd8+UpF+0slGMKIQqZqdAH1UG3QWs7hol
YlSehharxPyloh38AeZ14GkPYqHuE8ojNGoPtm5ScpQ20516aptyEdCKXelksmwRkH6e6Kmw+VEH
LwRbuviyjltms6liiv3NoRYGDi3BVwacKDBSC5S21BiRmaS4k0DvaEl1mr0e+yS61m9lHHptCbxg
Mee/sOeaB4CQTpIc/Of4QoIcZc6rbf9NC9EJrnJ7Y684sdNk+U3PcUm0KMERWBvJChNuBzJqdb3V
wqfSuDikJ3QxTmR5pVw96N59zK0HMCZgH5LTLsqk6HtfzXpDtjH33/r0+T5IEtStdqKscNdH15U8
v3sHrEAwMPw7hRtWuAobQxOKLqEY9A5DGWwx7yMXiemtparEbkOctiOrqBj4xgpTFTQ5HxTb7svX
DRNji8jIAmJMA8FdYwIqAeOIBQaClt8PQ7WyA95ibDyYVNYU0XwqXZwgwvRaSq/kqzjYTzu+vzlC
oCka475W9bwaZ9Ff+W2bqKAtJsiaRIl6m3MIK1Vpn9NwkUQaJ+O86oW54FM9Mx2gdHHIsVhp9dW4
1iKZHF1Kei7AcLP1yJYLUh4olVEto9nG/uVDPaOph7efRUdtDDGokp2ApudRUnLoWQofThyxAqor
m9zp9wsaOXB/JYjDc3lR5kvsHmumL0ty6JRDTduv95Dg0AH4c32rM178DJrVsLFFyGhnd/JZOxTn
jYidZs3Q+m9/2WOw+eJVSf0U4hia+zAFYfXyZ0w9acIu+ZXsfTZl3a1JwZL/KKD6d2/2W2rclqKB
t4x6s3uRir50lCmO/lXeZyc66vOPLliQfxau+Zuvq1nHuauNIeWQwfirMZpcc8tvAg9OAlHKQ9Eu
Oa0VBbVcjvmTBSJ9RGmOz/75Um8hwmD8yRqDj/R5842uyp0BfxkRN6zAYa2aGL6iwSqpPlOgp10v
E+fCb0AmTMqGqfuDDIOSyiFVJX57BFgl8O+HMDPn0xbWh5qbyWG4tWE4nsRPN0ycAmxnMA2T/UBg
YaVWSiADsYIHuVyVAPstZUR+N2+PzL4qcueNc6I0MS6Y2HSZVj+qOiZQn8IRQpMCrGnzHICcOV7L
M2eD67Mdd1X68czs6MoobipO9gV2qgSBhIbXDgizZCj3rLERa6Pcqx6pu04AzISJ394wE7OHGpjp
HyAIscExzgMmk/kI2UmkbLGjpesIt4hH+oh0FTCWF6L/0g3xLcqFTlnZmhG62bASivqPJEVby64U
xuEW6xEoSicOzt8G8VnGRo5qIKrGjK8LZBlfVYIFfEMnunF1vPQnDnK3obbblITaD6ILB3IJ59cQ
e0CcB7qrh+v09IVhr15BJESL0m4HrgrelHa7yoAjq5CtuH8q/qqs29k8AarxHQRzzJTq//lzhz2R
UdRNyzMA6Rf9C21KTupyfvz0/enkXwG1kDFdYINNJcVkKdJ1MUQTMdv/b6H5kMhXQAOraLnC3FK0
t0scNIyal/9rhZ/aoFE17hc0lNrMNcz5T8L+0G9r9QxA3of75s7+OLfYBHHZPQsveHNU7CCLwmD2
erjYft1UVr2zquTs1P+pyrQ+/rfhSAITY+de8DiVn2TpYl4gwxp4p4+CJGJVvYR9630LgWXttRl2
e0jXRB8sPb+yVUQvypO4DN6nA37ZqKrM1VLNLxJo/4ltXv2tEOkgZ/tjtu6nxpoP+imhy6OeuSso
FjszrNoLWk9LaCD9xRaDuuO8ByC6KI27T84gY8zalULOzgTD55V0meSX3eevdkwZY3ZJjQO9b2kd
n/cuy4SEsEofw086y9qPODO/S05o9zWnR9FJKSq2aRPM1Onfzzoaav5Tkuk+h/Oitmv8qppQLFK1
F56M2qIVtCaxd6K+iKexiDRIEz1/yD9i5ITN55JUvsh1C7DHblKyxA9TEdECZLAMyBXdiyVijuxC
JcwoR+gRF9RfIGzbiaVCVTcWroJsjq4IpI/LSdCOqL++Y/H5k9LGRU+huEx82KTgmWkv5zIgK0Ts
6FGoPwVKW36GtcbCnPXgULT0x/rQN8q1KJQlDW8/bhpC15qM7XJnauAmH2tytpNtmDzdWIPrqUhq
tzuHOMlVtzaVGrt5Px6i+Q0lahPyPSySvDdh75Vfs25+OOoX3tZmlvRs8cbff5Yf19uVI7ndfhJC
nRmVxXqG/a8FJhQArFGAM3V1RY/cEDCFVQxLOsql+GqZPF0dQnzvzU5LQ/Z1wbBOZZgzgghwxNqD
sejWGnJj+By/3QWhxZDm5LX+dE8E+XKxoBCl/pSsRYKiHN8BijsKIrxVKAaxq/GJk+uWgNHRSMv6
Hyl/ZtukdiO5ovtcUaVPhALOjLWtgrh+8yfQpTa3eZnmwqxDfs46+Uqcr7dCboFcqpDuZzyLihiC
Sc5kfa4BK/MW1q05lgU8/jzsiT0sB9bMT998kI2egswxb5/UVX8o1kI4uRLXhW2hcJZKWXtIfJxK
PkT1GISJUBfb08Swl9ppQnf8MzOn61vVYMBJgLyjzNcZJsxhGZTy5RrgTBJjo9J9Io2VySoKmjqM
5O0n5Do9WsLUdzRmuA2kVJiq8KYMozqc96fvZ4dFmb/K2zqZZyfV+OvgpPa+YxbsFbJhotTZptWY
WQdMxCL+DeupocTKi/SrstYDdj7xByIMfanLNwUN5kg/BGA57MtD7Wi4toKsyqOpTj9cM/nYqs0o
DxQDvr5hhGqekE8QJpMhpxYzM0X6NOKxQ/iLJBKfVFkAUTZZLdgMK6Wp3fgcD1OMmeTQjknKh5cW
x7UclE3R+LWAJ54owF70ughOR4a4NDVMDdmN32oTFYnyurMfjOwLOmWo+ED8NM5WAZvGPbFyYYaW
fQPAppMUGU16opWC64sq5RoANtpne31V0ha0epyscgjnh7DZCE5GnQXWOUcb53EvzXEUtEk4yEtx
FZTYXW7quATjoYVyKJT7+/rtUk/yJQnE8wHQ8N0mOvNNSjnfyD/CeNu1S9jGvRQQ2VL6pmw1AyVf
KWFlJTLvPxOjy2VXfhwt+X3LdsU3me3hRtsvlKaho6WOrEDWzlDG9rYhB8I2YfdBOl/LzS4uMkiz
dTPuvEFtDY/FEBfKYvENNJglfTjpb75IgBK8gklZCKdchPcdxgch18aW0vUwjIWBVlZmEyCRxcqR
/qR94wr/KQhgM8mVKwdeVwCJerUjaOouc5kJGjz8edn2FSKDf/SNI1WkJ5E+6eg2NR9fKrHfXG9b
qEU31yxdC1HNEb4gIvHcMjyXz10n04lHyG7GSBd+QbXdtbZ1AT7r//FFqlBRF3rB5IZ6bzTL9pqc
PBuG4nPfG6yD0JUMRLFp8aR7vpTimfQqzrOVKwNrkktAg4z43Op0NQPVnlPEGHao0ld68OFDdQgc
ngaKntSdiwVVh8EzAPeDSAyeyrng0jiWwOvWl/1DtXB8MSAQvYBLe6TZl0SeFpg6O3XF1WvtIFLO
gVvTEOxmwBqZXM0e1zODgndjfBO0jDqpVYnNDKCaiTQ+eyQ5rzZwIPtVnu2oIXptML4paT0xja+F
wkDkhMPHYlbawhnBYhOn2iZP7FJpq7arimOlzqy0nQ/+n09Nh42p+z/kdVH3aOOW0PNbg3bPOJES
OkrEupYZfbjUgKYwwJBTI1iFNi0nNSo6e20FwShSKMaAY7WcN2ZSQn5a2OTdVok73QGFbaIHOSdh
Nf7XMxDTsuB7ithWoE88ik0LDHzwLpdlJSL4EhB3p226OjA+Bo1z4GdU9g48T1D2ED34VQEk8lzM
l/f2wC6i3hRmxqmi9V4SjYlb/MiMnfo9ErpG4Jq5z6Pw5FBgFOEpkADxdRH/1xVWpT1Yvm/Nm0do
WIn2JJdZT1jNhcgN31a8qWZ320GrNYu5hB8eyiLUxe4QyHDNMxmB7Rel23FgH/saCLKVGM3j/CBc
W/oEGLNMqw1pavqysFG0lQqSKoZGka6cF+xUwRXDsBpzjw+gyzcXqahv5GzijxJcJw8PE0wq1iac
HpgIxR+AfSH7wOHA93mY15TqBtSUYBojs/H3w3DvZkiCddkGBTwOj9my+uqAMKZXRAIzhn5gMQvf
ajIPkSLdhsIUn+vymJkDBw0G5imwfX0wY73vsoo5844Ttq+QXpIz2RM+4xTxhbWNAf2ABH6g1Om7
mtAolQy0W539Vk838nLA2gBhszA3J4FCphFUBx2bI54999z5p/vdakORUY2mdpwiH3PixiNNzlgj
z/tpf8p/g3PaApPNlj6rCrSOteyTuSBa2CoGA9R1IIpBdMLIMQOx+Qwd2jcHvzdxxVYVTVOz5eeI
AS7bF7+xofBGqqylTCsonpUdDRviDcF5fxpphSyZU6/gX9hAKrJHSlTeIh2ppQtDoPmo6cYtvHn4
lpCLsSB+quYvl3ypaUxM2hFAaYfYL+fs1frxkoYa9+vWnngjR7hXhNk8kE31edWUlRg1DaP2oBu0
Tr0TFG9mF2PkD5gs2ujSH1xtZBpQfcj5uA9TsiWrWHn+I7vdkP+L8iovBPuKaixrqMrxNASxj6nh
eK4erBdolKZcLLDYQMHuO3/cHolFlQ3a4nkOu7sBw9Knjrz/lOk5Bc7SKB8GhnHGMNuqiHikzMd4
Oq/8UlHBdJcv+mVbnIZjKnGtifUQVT9i5e3XHbALOfTBa7YGC1zttKVl/YOaSB3cx2v4Uw0EHasg
/PYv6F4J5/0TGmEQiv3pLatiUjOggRQzOqTBqbglFReCm7F/92fK0xxp8u0SUr86LFLH1pmVrnaE
GBuLxbE1xCo8lAjgB2Ea5dWcqyJk2JJaAzIt3ewAEojJ3cwtw8D1v7CfzSAwA4RpbxpWOkD3BW1n
KOTh8zI+SgyQZpr+W9n4RQz1+81OA/HDQliCAUmDccj2LlVXD7YFhflGtAr+LScN+SjlQQipQlzh
9fsa6TIvPoix8uPk8FnelLxqlzno1plIJWwJ+yp4k672yO0zjgZJF5G5FcSmO417efH/MNF+mOgN
uaa/RpGp9QMkVmNX7Q/AiJu2ZVcmfw7m4zG+yag30bVI+x3MYwMK8fAkbw7qAwF/U45jShPizF4n
zRjp7i4yARmpLpOvIYgvjC2uAHtAIk7KjQsWGdezCTfaNRMc+iUFhs3yrue1EWEInam4T/66OQkD
qs53lVl9psXI9HT443UFo9/dENcaadSKvgvBL/R3xUuPQO399wtA/BPgU7JGTiyeZKpyQWly2AAr
wTgIywiunzgrB5iSO4VUFRfwAZ/QJJLwq4dIy2OqSoCcfQCYLQdXvIIQvf6dLIhxTETMMvo6WNn/
dclxpLXqk61I5MMU7++j49OqZW9Wlt8X7pw/v75Me1P3/XYOl6ih0HsZA3wgLyWMaY5J6HP8hHnL
a79GBRiIE7XpMh5l9Gob9s6XlJoQxvJmymTAlt/nbQCpCNP5h5fkSfy6V/YqqQIpp0AIkJlxdNGq
baLnBU5iHbJHxiZm++h1umkvbM8C9lDlWf3uLtkYxqGvX+uxLyzIq/wXIS7x44xIxbnnBV+d2KP0
esucCsVopyYADFHAu2x3H94GyLPVyEgsk/dbtHIhP1zsGB7x42FuFQ/8yhRKccH09LP00BN2UEhJ
/5rx36MRnNYd1yLS1m2LtIPVwe8/QdV2Fc1n66oYh8tgCB3mKPScS5fQqoZXF6Hq6VwISllANJkq
cORiGa7ARyrNaZYafcSCByyg2AU+YGLig5iTR8aiHW/4f24tdLhyjiFSxSy8Rl8TplilKbv9b+FF
VevNm5bC1LtEc/vAE6J2AvHBqjpDKHCwkZpRSVHy1sgadyQMMsqMabYfOpMRwO8xB1/HEFhf7gfm
J70GL1gD/hg/JblLNfxQ3u9FM5SI61x31STki3ZOjuKaVyc+iMq1uMRbGWiWqgZxH0O++HD78tPR
1c/23ufjXQ+xud6aEBLr/vE6eXj1Y3RnFQhscvgHv089nLKNBd4g5vC/8CpfFvko6HItUQefEyUl
7GtF4EDGHPk5TK2qGPEsoUS+CtBSO8x0xs0I5z3vphbhbiFTtvasFmp1iwiDe9TQIW3i3AryHhVD
itrCDx9f7PMgkDKITcCFm95Fvtu8stJBGqoOWemPGOUF//NNcgGpCuEYduoycBDW4Atd+MkDqAVE
TNzGzh7P/CREVDWhR0VG6B2DmAEff67iCSzdZ3iYYCE91+xANZPc1c5pStHXaSbRCA89HQ32QE1T
YCmJa15L3MMwSlQ7hK0Yue3x5wJu6dmSP5cQvyYY/UjQSOltZjGiU63mJzCcA+I7hSZCXs9+5KgD
r3Ng4taLjCt73MAWHhSeA4YybfsL8Bcn8mY4Iu/YnbJ5mYJ+0aRhggQcA4EV56K7YCSDmorRjHA1
xkFUEWlJw1sFX/AX0D965z4u49hyM4R3r6rSUXNDnmBwiUWonBqZhQblsvqizc60uUfmv0JiJ+75
5AkFd59ivD/wI2v6WnNsnWTM2NBWtvZKnn33oJ0V9DLD3OHWi+BHW0p7mINwJcp6sfMCyhX7f4kG
LfEWo25mf2Tuwy8cA8++t6Eilp3N0KM+FKMlKM231qw6eKDHpqYgMAC7oSCr/Y2JQhlhIdUEs3hX
oU7ofubnE2UMIdbYaUhd1Da07nfKOnJ4CrXh+2Zh0FmPpE0N3NkdKiHg2eyQHVgchgIPNJWBM/M3
aKcZpgy/88ajH4XUp33W41egyUq+boRii0md1f43HL0OGQmoC9YPaxfFUtZ7LCw/ikby+z2/98ZK
jBmPB+1qthpuHfUK5IWHm0V2YVRZskt3mW0Gk/+6+1EZGZRoNkntWJI/zE8F7lsy00w0vcE25v8r
13hVf1GbwwIgleHI8pWBlt+Gx/nzmxExOtLVqI93vX8KpuhFtBiGh+kg72QnDM4w/dbedwkzkUbM
w5fcapuWkUPJoVVRkaGSmGG/8VxbH/MGSMlzGRoz4Qaf5R6mA8FpsGUXCR3A19e8N2zmWzjnqjFn
NamMVJkL7IWtv0oU3cu1UBQb8Maho2l8PrT+SN8a5T6kQBW2rnnJca+aCGkX76gcl0E+D0bDGLeD
g3xI4F6Aq4NnYfc8Kux5Cyw3ZFxNimMxVagOspo+vR3+YFopc+8R+AdOak3b2U3sQ0HuxEPowrou
Ir5V9ca65FZPLMTDJo3jpWiDEZLgreVRnMFZuBqGMFPWECUu0U1ZX7SRKySCidRrTM13HuBf9rEU
ih6FMltpIIogM8a2nWHtUG2ZEBWGwS+Rfu3U10bumTMUNndEAkl/1Haudt7jXHjzNxojmfr4efoh
YmWNMy+f1CW3ai+7TjBggqxQRo1rEidzGfMHHvr48XJPn8fSUXLOqPgksUJeObmeTFLPIfGxvEH7
VYfJ8mF/iToIuzQIb55zjQ8Lz0BCkhKfvbzgntjMyl6BpD1obi2bOzsEJBo6IIboQ/twVW5rHLkT
GLtsLeMpCnBh9KN3gO8VUT6cFJRQdU4++8sTrt+FoPlfTr/JoawHU8b7yeUiC0/EW3K3sw1WW/2C
PMT/4XjByUgcJWA/OcVig3XIaPbNKoyPRtFjFZfSPKf3Zx34gvwV69LfjHobJ/z6eZ17C2vwuZn1
XT28QF23XExxMSX6LZebNgT+hYmud9T8audwcjcaJt/bmEZdn+RxLnYZUZvvkZoxopf6+eQf4lZJ
mCOXz/OIX3qmhIIdiA//iOLIZSe3sHg38po6MutAeVFAlIQU75IMJRIZIq1m5O2UNNV9ntCrubSe
rmn10IPGPwTxS6ytvnxLX5uV9mFNe7bUgXc0Z/pRoo3yCCcpDcH22jGGTtAktISwtpmvKwmJiD4J
7a38AnBqX3R5TLYBm+l4OD2b3RR4JfyZi2BEre9CnC+B+rm5MlgLQnwGPSjlvrYfFL75OBb3ZLqw
F+K7nu6xVQQEEkYxfAp0UmA1liRhEwY67eLXkPTBUGtE7fcGS05ui8DynZxayZFflk+Jpv9X+jX2
NiIZAbmjo6PRNmter+N69+Ov/ucF6isOOD0wDUXS+vQ9v2I4UuKQMdo/PX21U35+RfUCdrz0r0gX
9X94v+74dmW/32uoV1dG2Fm0+RiGptybIKAsWuYVDpbq6tMByizfR+AINZcP2gtSSDH6Rtga4YHg
VqABLZmLiqRYkDhiDXtRPN2IWlF73EMU6iLVNWYXNVodYa5JPOVI8igo7FWcpbgf5sTa8vhcw3eu
gK5U0mPVzXPVpDEig/bmPB1q0tgFR1kF8l15hOddhQqB+v/FyY4fYPbjp223u7SO8nSA38ueggWT
ZLHQprUBlvP6bueGHOPc3vNrETWDgoe9j6BS9BslB2HuOGgbxoPXSWsZNZAON/VJUUOyYUmvnYfI
80gEHuqWvKN9ZCC1FKfdKOYUH9YiQ8TrqIfjDl98YVDFsa5CtKPTn+qBcBNn9MaqEyAsmK4kpVPw
OaJmykz/32J8Rjjj4Nh5YdOljKSTTf7FdJ8UzRCIL5e5Z5i5qNX5dtFL4P4U59ZclwqMVqnAeh12
/cjMJM55rQMztRtHOsCxUkPRZmQqAjfSXHdsnIIhaj+nfHw+WU+yNWvYp0R7cFUZcLRmEOo1RXkP
VqS8U0xuAKgs/fMmMRIKjo9A1s59WnwrT0ODOTtimESVNLQkUkE4tuNjPSEggHyR2Q65/BUdmAsN
v4LyYWtoShR4AxKH8jyKFz0zjBkWulr+7lFws5s70yQ4r4OtIxIJOwtnGRrQrwwIoBic+mkWc4mL
9CIeWdbE7JR9icmvPt/LUTi9osm/GTcO9vSWoU1OqFuW4e4Od52L98iTBGPlmBZMsPtFGdlcQoWr
gXkkclY8a8Wvt8XFMa0wJwNkI4odKe2ErM/KO7CwkcC79di6qWkrEPRM/27djYTeLcmUV4XJADny
FCbV3559AsYv+LF2vxq7ofePd8ExCQoRlzcQaS/CF+m1pifWu6ZQI5s7pf4UYF42FbpXgn4WBKBb
4Avv6MuPOSdgbvBgx8GMwZOdpEZHr1Szh55LexfKsy6xV6huXSlZ54fSF21T/dItm4ptKTPXObv3
uu2JKmZGB2fSGvUek77j6QqaJRUgzC5jR9HZE1QC7ILcDlhIgpEMkRCJHP5z209p+sHLU9sF++t3
FTZJbthqBfnCWsVrHYk4DmB3SqcAOrGNaiJp2GtbE7CMGDQ3HZEpMgdwl+2UR+JoZzMjVKw/UMkM
oJDsYOZqVy1HUo+VreNsl1DsnWmlMfvCsegEdwl/6tv2Shvk1bTZZq3S5cwZGKJ9wM8lSyQI1uEl
p+Po1xcELR/Rsyrt8O17H/5ort3VUc1cU/HCectWLSuXvm6RP64BWacIhrxg6NaxnU+UTqPc/D+P
TnTa1QVGpjaomscWvQfdGuLhJK3UEyt/dLHAtb+XeFQwhbjg3M+u9LKITcSuncgF50xYhF65CIkr
6eVJLouqePHPTjZcw8lAnhyjXrzMOU6PWV/9CaHlLcwN/DYRuojL13+YuJw6ZlbSPCka4LsjA8cN
34a1PX5IAgaZpsbRCG0xR2RSgsas2i2ZxnrdEPuH+eZB9tuutTKIk1YupbyPf9cviDPu8ren+ke0
ns4U3gIjm7wAxE7L8u1Si311TcmEGyGrFSoGAERj7nJ2Ejy9qSb0mmJlnatphBBMQxw/BwqHSZN6
cOpsJ4x+xnhrjrz9EOkXkoMvqmB0Q6DaQ907A+BzIE1d/oPnVcvv2+jRrEKaOwRTJW6zOBe+CdoU
54HPe4iL89RPF+NQx7anWER/Y9RGhES8btBgvconJ7XkSduYqr+//+6jGZLNJOZ2w7f9hpCYYxGi
7zBHiER1O/+Zlcq1tkjkuYxkymg3+wc3LBSd4G57vH+UuprtYO9QRUBydyT2KC1soZHC9a/17VCd
PxRZsbtIUf2rUbeY7+z7Np//ToA3tFBrpmBY/EL75XjsDM3p/kypJSSgdiDRDpxPceEf+6P64E1B
3rgnsNQkqvZahS0ZcaZSvb4y2Qr8ZlC+t6WSNsWUG13MG5bC+2ubfa933bz+3cstg/2Jlajr1u03
SNRcg9u96wEnDdk7vxU40JPpt58ilbeacuOKLg52kZ8gGDKqWRQH/l8vQyfbxgLKjoFZUzsG7QFj
6v1kupAWi7hSga+lTyI2vH/7zRrjhL7IuCHAbiM9H9LfKgsxu0K2W6IaA9jhtVyxaGRkFsWmkgOc
5aDAqYC4CdX1YxAwV7Vj8GvrZFpp80KzeyxgXopmc33FrkcCJHKKVlhqAWwkzpAd5tIrqywdHfQn
P9bkUUhFnOBvyrPtXZWXFVTQ3SmvEwSa+2HQPYJz1ZTFIuikZ3vylcgWQyfrhONN1JEJAXe/ucQ3
DbDGJNYPNofRgsJFYGTTHw3da5jbNPKMHlR9Vi38M3c+oAQeQPw81WWgNSVMaTfK+rr7HNWmHqwb
XhNSrUOmy8KHs/AzF0r0MTQY3dWOxNMtyU0oXMrl2TR2tdHqGJWOW3wqJEDgk1s2GrSC8dyBxQVd
LtGXJyc9bwuysyOtgWllAL9/eYzlf97SV6ml1fQ5wBA8Og9QNIPoOtfHhiogCVPu2TD8pqYo3eZR
WG0U+AHkZ1s+kHmoGKGkdttQUDBpGOCA0iXLatlmPm4UuA5IkKNFHilGtE32nIyc5ks67d8TfdL6
kj8U/3Ceh2KtZ0uD8cN6xLJY0vK4bCf8VETJhBPIuZoUCn8RE+6zvcUqmRgHVDlqVx3fPv3bn5lg
83O3a/qMA60W8x5RbulKr6bF5Hkc9gssM4Rh6+A0CqbBgme0N/2lkySAU4jcO5cCl+WoJMkxEMQL
Av9eM6ET4fWL6U0wJBgKKJkP/fphZWiHMAvfzUxKbZ00sQq5S2LCEMNvxvuZ3xy+tv1+56+/tSrM
A9b6B4ev0NLklgI0j4S/6R10OmjWSBrAhlaHssy6hA37YM/7Zywy551iYB+UXgYuPoZBTUAVWFQX
k6Mxj0TQ05M8DLr0nXQOQG+9dlFzGH6HejCyLXyRiza+LAPhSeJiPE5KL0fgA7RZGE7+9Evbj51n
+VL3Xlw2uDWvpMrjt6MinV24/pA9vyah6hWmt4699Eey5VISUmmCGdcAN6xwxRRApt/exiBfvHwY
lPQWodjB/xWIQwHbp/d1L4DVrDT6q+YjeyD2swpS6U/mNbCHy28wovHT9gEExj70PkXAOiMy2t7E
auCUAk6rLGb23qF8C/ATOcFwyIiVvcr48TH+W2Jj7AgfeL1A0xnX6izq79Whmxc/UcQtHsSqpWUs
9Yr5DWC7FUkYDeQjHB0i7a+dpa6f4ZIqjPAG1FQYCFq7OQS/BTbPINDtPVzYKT+/GF1MucEyxFxx
X87doPb7/1Bvm1FeRFEA+K9KMcZx6/xIYGBoIigDjQGA/T+RqtmThg417v2iSPwRwMgoxwkq5tri
Y6/Ai4/HZELCmYjww9ebeYVhk5AO+B6xNe1Fx3ashydFgK145kAEW9LOkkPNnlzGDz8QWqYdBV1W
J7tObzAwzeGwHbWgbChoZVAI0e1kyyjSmuw2lz6gvbaHsJrRquPs4G9qtG6Q30Mg/c3lh7qPMWld
CdigVz+e5CTxmP2inA+laLMYjXYuIMOBddpoxqh9iGEoFqh7l2Ss/Diyo8zjsCoIVc2RN56ZlaDA
B28EUj2suj3/Fq7QFK1/fIgJziAn1Pyl5UBv15R3OAuSuPPbPXHGM7xd1e0DWvQPf96aKSxrnsMr
+Ipcxp63wMWmY03GTYCTbm6DweUUzP568dk4qh5QBB1JKHPnnNVTDnQ+/X3aQqkmW9b3p9dSgDfy
nMjTTeiDXG8zEBrRXtexkq2SKhlUZGDf9nN0qyN3qairFNgy9/7i8TYzO3H2b3ZpiZcnJrEZ16cu
01Aldt8xABmLCjEKtL42sVPCdJkj9qilyYYh6UBvseOS5wDxuPSd0ilGbVrIDnwB/bMgfzE83EzA
IuP67NlHwfZFE3vqkYm9dqMrvso/Mkpl+S91LD0pzpDeg21aUUUyqfzT/p3YAwmp0YdCrDOmhM70
o5TpzhDjiuuXyFvW/K92XO5fpcxtA1IGK6Qr8pbZC3ULfhsvyJFRx3fxtLCvuLxDC1mQHKS5qTe/
/4tX6pm6khyPY03Z3PbADo77c1+iGwzZRlDFuH2rJqX1Rfoh53WoCDTsXUaXKknPC51K+buNkIth
PgZ8p9sHFRUXp1+XriqauvG5KyXXouTNbMSamYeTjD6uoUL8owO34xD7WqOKrSPiIIlu6xkq2hWG
Fc5JiW9hPREozWRVyhyY4EcXwOWdKJeG3Zpi/3KV9mcGcft1DGfAuDqKi+TI4h1FzWB6rOivuYE8
eFeSsIaABUwiLFrPMx/jbEQgjWcssthBkmiKECnmNt/gx664KPVEoDjiySyRHvW7cCDo4JktpwBJ
4MbyuXsNfQCjgpi/zS77m6+gOWw47psfOb8ilL5w1EBeWkIxBg60L7mGI5AjWwXD5xKZnkdmvJcZ
C/+EtJrcchWcT5ILocEP14sVAD9nGRF6a+jndwTYY1oyYQ2mfVOL3xiIWzdkJT9WOPtpK+TXECIb
NvdMyR6iW/e/HC26YQ44v8Qi9Up3t0YScjzGGtCLFrGktPGU16X8efXRfZs4nT335SO2tZQasoUk
UoRukJtBAtzOilMtvltt6496U2RihjlTEZ5nDpa6INGiLrM/aWz1ervZwGzw2TY33ymzYVG2NHgT
bPamu2YlunGwKtfsswQ7z0H4XMkXcxzgpkErpdj5JiO867/YIFYKsZDcwskYq1BIKQ9CbWUmfC8X
IgkBZJqVLGy5YiPAcGpEeA0gjjaSuivIIxcWJcducTIDpBRlx9l7El/pRtcnWjJ7+8IrahU+6aur
npxLDUjwtPISo3N6Mk7jheehZNHA5iRbsB2233+PlE5gWabZc+777a1NsKp7lwISS3stBPMLSpou
OrVJYblzkB56mMf7SDLKWJmMIpiTMMmUPWqf88YweFFxTpZWPYYA3l+OCQ+O2EKYntr8g2jHBZBF
YT3CiDLGKqsk01F39ETCj3zgqhyB/P3DGsPliQIZzpWu5y5T8/GeG9edmeDefiGMYu/ilgFS8HgM
hNri3h/gjNVlxgaZPvqxV9KyhKVpljy61RqgeGNRp7EWA6VkbDPMzLm5kj7Se3tek9qlQFZH0hVN
rOmcHJbgXkkYN8ZNlGSy4J6JWzG7VNlQS70vgwBxqNGQx+z1SAejd4v3bDqjbBIspSxpSWhMSWnW
uDvAOxcGCs+Ur7lqgP1Ji4Cafkqld8890Tpr1ZJxgUGvuj3LfFaItUJjz8urzSkei7K+Xn/KKnKH
bqlh3PKEZjsm80snsF7WFXvk3/CdXYSEXHwQDF3tCrL7PET0hIpCjENoOIknvOs4pkimNFGq4dVL
Qbr5kgdNwMexaWgjNEzx0Bsh8LsOdKLJMsMw2kMm2zJ/K5HLC8A/DyvIYJ8fzqkh93yWaykWDsq9
wrfbqmkG37eGH53xpZY8GgN4EEi+ACH54yctarsRZqUL87q7AaHPL6DJVEWT/kUtyu6bNb564DWy
Qe2dlDhV9V6I2zhaq4QMXg/eNRCk5E3PuwFR9Pm4tb/hsoewpaIcQ5Hxp7YAGLwnMLHDYi85EhLA
2U983PhTzgu7XiYmU9Xkj8C8US78JatJ/rypbn5FKQKulKglVsQvVUCGNmg7IcyYcEN6K4kB9/br
3anyhb25eglXUhG3pkcdSsq505B+Hbj79jT0zlrV+iw05OO6y6wyY+rPYukNDdZMDb6UAKRFO0MA
MDlKr/ltkDLN4mozh7aUqeTXlK4LD9WpeAZhuiLBpxHBt6GyLrmprzTaTfgrdoNbDKSCcWBjf9vE
O4usUOvpRyNttyyD8uOL0ysvLhyeztuyvKY75Y62ssKZBtBSFUdEzs8cfuCFjWp3TLtymb+1tpjQ
IPdtRsHcOb3riUodMH/ZSyIhCB1uCJ3crcFIZ6bD19EOuUOyFYh2tIde1IQvXz4TYapRVtS12aCo
6rYpfoUqgsT/Kg9WTfk2sJFW2+3HN11f/Vs2wfbl+DUgJje6Oc32CAiwQDP3A3QjlUmKysWF09aC
UhY2iqf3NrnViudAHH1qJIJAyo5idfw6O+pPDPui77fzZ8PM7oaZQ5SzlHednRjNsLX5Y4D8CRbu
v7S2DU8uPBnhm7cs5Xyg+lvowvU0bj3wo4jI43nkJbV1cG/2c/WdS55zimgToRynR7eCBtRqvJZP
i5dMGx2nf/LSF52hE/3DnewpxBVDyAQRCsqYiKvJd6sWnunf5HpjLchEP7HEFmSx04Iryp6i0KQ0
73Y3oOuFxH0yvHH44/HcROnhVb7E71ydzB8jlyMZB9qzZQpmqOuipoxSgJdtOGSi61JrVSlaEYuC
5OP0Ezr5hf1fgruEBD/pRzpT17pTELzlSy1QRz6cc2zNVaneNs5KOsqLpECcPWlox5zH2O0H3in0
AOr9CZCvjazsWYZZDZFXYasV0GvDeiJM0u+D32+vLhUj6Q7SUOF4MOy2WEq9akvdXe6byB7AxiEr
2mMpOeSbbAgHamU5Ww2eg/nX2HrxrV/en2gNuw43dSjPwJGXeFMxCSNL6b27Eyie8Fi7zpIj7r6y
qctQZBZMOGpQ0EhBNEv/0rXjAlSjJT7z7yODWJ4lpPHN7ZH852v0szm/l/coDV5wLKjelzg54iBj
1rvCqsw1umlLzgi4HxnoMn14rmc7nbgpKkvarRTs+e4dMpRyreyS6hb6EOgGbVUN7zVwKguevwRB
zotruJyV0Zs/NkLacPQkAhGkZOOBUvyi5erWrSiVrOBWZ8S3ebNia57pI4eN+3Fblfsi0cDFsAMT
rM1rklSMqnyn5XNsWnC+j/Pctc/EvGYXLjIINzOFAmAOMpVqDmiyoOaGKetkF6XE5JvyhvyCT+N+
gEi5La6cU0pH7HHYcwpsB6tOGwlRkMy8auT3X06neyjeZXVTBj9H+lLBpHX3DckYU7iJRSilVFGW
oz0dU4iGaN+ku3JVWOUwwXkH3zzQLCzeombUHhjbKHY0UFNpygWlzlx6824lZmWren8dKB7A+IhF
EYpUO4QN5/7YvDnJl9vUmVapVHVWNzii3aX6qFCT+ecOy2xptufh3DnqEMSqvPYtvJpZSxNL2JxH
r/JrMpTCI3t0OmtTyqwGicvzB3R4Wwrmow2hWR2ORJ3D8og82lpSlybhbTxSkkN95E/Y9oqwqKU4
vwvSdL9qvg1gcc1rZWRm36Uy2YhRjJb4dzSKu3B7diY21pOspFveTRYLn9K+5fH7VBBtttHJ9Wya
tM/laqHjmd+2hXGE9HmZm9/j8BQZuOGzvJ/fXmvXufNIDAJfp/9hBCl1k/VCd8CuuoodAs1KrdXv
WuuWypJp2mJPci5EVpIHrKQhkkI4fBbBVB66nNhxijgCD40PN8gsSSnTxcdC/bS1G7aRTkFDiwZK
Okxt3GghKTRTdTp61nYdlbSrndUvk+CSY7AMcjnO5f2G5kIuOpxou0GtdTipdeyslj1uy6cVFHo7
nZdY3vFPOtE+iXqAJ9ZwBbhM9mDO9svJ1/Xo2fHQO/aK8rQO4Ib7YwN8cw7FChLBkRCXBW/W22qy
+trv7d4WjfxUtC7IT1M0XG26eWL3LY/9DtWQRlIyVIXy1iDu/qQsZlnctB71ZvD+sTqlx612pGJR
Xkjy3/4PVfTMJO+uJOknFKhO+w9+txrcSOZkUTh4KJWN31C4Z0Lj5BPg5QJRAfUP4lpcPWSLZJ/9
hD1jAzP1CQxONADBMI8RIxvZ6B6KZYgRn2h1wHfD98n1ggyMIDEnMyE4JmMSQNZ1H0blAC9mUfXK
EJ+ixscdjj/S1E8PfYUf01uiV7VhM8GtZlQbxn9uWMKY4q/sMxY8j0H9nc1uRil5TiK9H1RjOkyI
RF7pvo5lw8ixgafJcLsgKPhgtst6jU6WfAcxiU24XDjD/CdAPYrOn4DU243XLgPTU+XeqSgut1sf
w49eKrZFf2tMdVDlxjocLS9CiATI1XDE6GIoEwuvGrf4k4smEhrIhmYm/YDQPKZcKB7Zt27qNY1k
YWos3g2FQHRwMdLs1009zLA/GVBlqBervJRbuX6yyYwK7N0uw75NoeoaF62N3vapMRbkd6nqUAjA
x9149XHR3M7NcwNrVlMa+nm1dth1PgGT/aeuhzYKNX6m9cJFP6kDLVuAeF0QA7FI1zrVPk997ySq
2zyisaG0W/QJk9aByqGZJ4ri7VnGO9P5xbipyQDQBOsotfg5w2qHFDWOW4xmcs9JuH9nBtXCODer
irSO7ipBdMRuVQJxjggTklM3D9E8BE5ZelvL+Bwx8G/BhNLPJ2VOz+IvkwAWTVtDBXZHm4+mtozp
ZVQ6O2uYynMSnLlYPmlvLyqxomEQjuvBmiCzlpiJlQjIiw/MIfqmdDoU0qKRGMLSraQjAWZEG6xj
d08E8cz07XcJNGr8xjyOwIJ2NaqzrD6RVVysCAlWXxmAUbyRYoLQnBDl/df491MQLfdngbx4NuVi
2n2889t99lPfgkooR85O5GoxOCOeSuicvjJZt/cjvku0VIbArfsSxq8bpW30JUxyU9H2KrQy/+24
ovzEVAgPHHMaGPrKU5U1FFP78m2cI71anSuPG/bWZShS7nwnynD9BL3tI3e3OlbBNshXNkIre0MS
h8jYO3B2whMFmtglPXpVYpzYcP+EVn/7yvPUa+AWfiGYd+Sr8D7/1+LNsfnALU0e5lkilviQxrUK
YkwiogcTAdFxEnIcm+p/UlXIq2Nji7z/+PIbU20IBvuwkVXNPLEcGvYjFRqcC6zuHx1U4TD5SJ7U
OYQB8lX6y2UuiLIkSo6Bgeth9tZAXuhTe7KexiWp3WdzKbmn5Ey0lr9BBjq/xy8t+C/n2pAS8OqG
17N8jkRFnLabfxNVy8DC9u0IO25wQpyeze8MvCbjVudCvlAUWQbehJYRwaxjEenw5sbj9xPuvFXB
BfJncyxSEJbcWil3FpKWxdjlEdt9mVIBkQR53VTG6q5dmm3eENeSgclVsefSrBQ3V4PfV1rnEDba
1QRzeRr8oV9Ng2oWr1c3iWt6V5ToEmew791MKEm8IG5ZOGyzc9jpj2iKrtGNDWweKLScxFouGie1
tHx2Dj5yubCpG5kKWh5ft80nj/fF2XWf2bGZp2YIPqJTeaBH2CtHQL2Y5DVLH7IlGwQaB4FcPnZF
q96Z5Ng+l4/nP21czCQeyc5OnHv32ZDlCG5Hgzg9kRGfIpBoFgOsjPOJMZFu6sQPlaSDHjEGJwnQ
+YP+CK/1UeZhv+SEB2CkjuTTWO0tQdJCQqmCYXq/uBHVuEQ4QN1dklLSaVhF+9hlqOCfIAHSM+wD
8eq4Z+bgCKL03OgmMA76TGX45wYAAMXd8IvrCZmxOGflYIMfBqKV852pBS//S8WR3YS/TUhyF+eq
MLj2/usk0Bjwii5pC8hBeKqsq7qPMpzuJTho7ZIkfwgaBTu9vo601Ktf2eppesHMhKBqLqealCAQ
LX+pTwJCdHQSo5J1Zqn/YcickKET8IBhMTvkGMAPkIGXMnT/rFHlc+79xSxC6dYjZt9+SEotMCNl
Jxc00PHfqfylvvAEV+XBzv1yDT+A/jjx8FTsLm11ElYA6n1aiCqKhao0kFksaqW2T3nQfgVKouGA
ixat+y2edGAt8zMzUzYNyT9Ufs1JQH4cVooHmIwqk0X9SormhqMwxQ4t0JGq3srWhaR+x77SgvQ7
KjVyk5yzx1S/Q6YLP3px81r/nbOi60oK5Yd44jyRgsGEWZVr6NaoRGw9WZxCTVjhv8XqfwceP6U9
0AhPZq4rP5DKGHt77nOaadxu5s6qKALe5ZPjr32JCoBJDUJaYv76McASprHtul/AJcdlmIKNRB0M
3IyRnfNVazvxQV4KJh2Ugf6nz5ozGb1hWXgC7NlNDSZexuZ0hIVRMfDzYnWGHq6rUlMqoLGGe9fx
B79kUXYe/XuYaxnRHlFBdP/pzUjP2KwnDfhfalqeYe3LBu5nJniFCazre1+MIGKnkWxGY6DYOdgx
WDYPrSs4b/T5UvmoyVgjKW/A8WHEChUlJBKSVvcBtIMFfhgTu37RjFpsOs5y6O7L4dmUNA5YlsfD
/BZ8XiQ2Wbz+VPqzbaoGzIhc/VGkMlY7lPgIMlDwFry+wO+/HWBKPQPECkTg65At01bIXTagAyWL
b97rZcM5BwgYOrHjfBa7zaI+tLVTpkS8rEbJNHmPvVzSlOjlAy9UFj6UHSQ1sxFJMBUPStSPwMkf
YrSCGFtLwiNKn6syfyGerxUP544NKwEpjrrnIhxkiVS/RGjfCP+R6zMBghP7Sh4n0/QvxeqPnqPD
kOLdsVCygRczjXPDZZLE7gz75vEclknTU1B0V6wBs31C8jt2vjH7Yd+DrWoUV2Q1BNxGYh+RfFZq
bpiPggFB/ETGOXaoUUDPds6AYEBYS9rhsLGdEmA2unn3gflooSqaLXRz89bmTMwyRa73QT1KSqg/
1tFsR2Wy2uZZx95k8Bj94yPOo7sKkasw5EprSwnaM4ZPPGpYtRZdSH9HH6WwA4PFLPkoEWWlzv78
iC1+zGHRymT+K2O+Xut5OYXMt6h3yw1rsJc2/79tlG/iCs8sjY89k6AbVcrXCj5Sd3xiADhk/tS2
DHrTFBb4vhppHzwSqH2crJxpR2xXHHKyl4sPK8qsQJJdZzO/bR6VyJsprPgRDloWvWDEiRneDuNu
i1mZpSSM4YzWILvFBLJJRn3Lgox0M2D8cbmGTDzJkApqj1AdBynLK+Ee5+p1vtJQStkCsYhJO+SL
1iBQYggt3JMClRonQIMEk6hjG3M25/iLEsCGKJtP6Ljb5lVfU6E8AkdC5asWTaDuiz6U3hB/eoCN
LkhNfEAx2XC6ZKc80aUctYdjzbbEUbZ9yZHr4N7qKVt3A0PERorFRTNcubgxQF1jhAdQq5nI9SsF
y6yYofepKlzfzeV9JNdtNxyj/al76W7665gvLXUMQYao8RlVqjXtZgemgdbJbcZkU8S8rfT3RBLC
rbcPPLciHviXXuofnMMIrrDrR/JYyKMuBV5wkPHZbVh12L+/sFk9HJXYG1iOIGnYNeRxtlhQxnD5
fIKugM3jhi1uvI2nTvbuqD58WPuIbsBw/H8Ip+vwiLQFY3Ih3o4wIyrGIcay0UE+YaIp4+2tcEms
PGu+Z/5JjuoNb90/t9nhamIhNPkZ9ptXh36VBj2VOrb9gDMOe8/T2NmdLHAc5v+FqypKVgY3an5g
mQzzX+XIXf3cms7I3+hcdhKTcgoXyMChCrUdcg2q1CiVrZWTYVL7ye8MBKrm2/2O/+cFErD1JRnc
prr5uYMdtTwS0FLpTwwvLOdwGvFORHMwMCEBqWzpI+Bt6nusJhIyWjiL0tRSXhgz9jIChEhiO/nD
VPtcJF+MrW2qcFlEzqQC5HZ3FvaktNwi56ztqs7GWMCWjFEQxDh4lH5Do+xeiAVyW5EoiqNx0x52
oJCyCDPmTVLUH7rgKe2pdqYkk4hpZjlA1tR2RHUJQa5gmAYcmO2m8SgU190rT9C2CoqsWbDJcbRN
gn5cIIsrbvnos9bpeUPqqELDtQnS4OzDvMLIBGrWqOnYNsj2Dg9wRNC9usH+IF1kmuAANZNNGStZ
sRc4gnaj26iGKQzOETDpZ1fknO7FSaIK2BlMFTVgdFAIntX+JvW9h0bcAaopCh6gCHJWFyEKys0d
wrW+j4Yv173a+rPxN3FerPrJ83xGtBHJgTyiW+rBQ+ZyFzJmpb0pF1q79fS475ZgBfj+g3DOd/p+
/d5TEgJGxk7mqK4Y3tMFVbW1bW4yfD0ncl7ghzBzdU3DLRli5fRP26cVOH3ehNLNUCz5EBbgdUz+
bg7IEm0n0wPFM4eR3g4MXs3MM/leU0xh6hynbotROSsHqO04f+YxJAKcu58dORDbbUy04A0ScYo+
4KZ603EbPR3OFKBEjr5WOsIejEsh+aZXnyQ5ChQicq7lwcdknkXwjEFSyqrLGCJVH8R78gBWmAT6
9oUB+7SPUfA++WOuljq19+iAMI9yYsglzUSwsaBfVymuG1dZZ44BadbHt0Jhh2I3+a6C+QCDthof
0XVOChd0vHf7vd4ujB1Itrqpk297JcN9LfPfd+4IOGFSevDCZgTMaIO669xb+Kv4wbrbKZ8My1SQ
fZUFEYcERY0ph5IpFOL1aMZGap57I/OIAWbPsnCrDT7uZMsKoqAVHiMFjEz94+uIl3q82JK8qbUh
GnjqWsovkGM86xaw3EDf+eJIz0/SUCfqtjzvSqRyb4WUtCAcmVUT83t804bLlJ7HsobAxQoC9pdM
MSBMlJ2JPJMhwIl1FwP1NIoJyI3qnFk9ohhtymkHLBcz2Izgwivx5lzaOYQCFJUKDv6fvEAIMIfr
LILVuig5o8RF9Pr+2j9UlX7S9yw51CXQzbXx47dQmWoNVr3xQbGw7AmAQ5uc8xo0mgD+CY1Bi09Q
NXyPcB3ZhEvK4YODzBNFMbAVuZiz8kVaibAuNsFDdnf0/l03d7OUeMmRRJ3P8KpkbqI1rRMkGveE
leLcAWB3NqtrasXeRihl4h8OTxaSZLa16p17Fnn1bCS+D1XMvN0KMmrajsocGUW9A9R6nwtz2jxX
zPtk5h9Xrj+YEkDyH42ppNeDqZXNoZ1omxdPeDhntEEbUsy9VjZD3AkrVU1jMLeEh6/aR58Ua4be
1cGr+pKxzRTf1DyRIGLl+8z/JuSk8ns1F+k+3lmCkL38ZFRD7AvPvBVp73TT4PMEOcmLvZd3X6mL
gJvwG373lP0M/ktZQuPoxaOZC416nGdnsVj3pgHDDSe3WfZWkte4S6KA7+KhXVayenu7tR1A7nOq
UNcyWjiTSFuhBKslSdShXBTx6r0mzzZGS/WMHydPg7K7/mTInjfPov8Q//4YwVKJUFLN391xfwOM
OSOpABG6R29YBUDyTNkD7RouIL/APMa5UrHTr2tNF5Hcgm32wa3m3SROw1CKu8+jdubVcpPhLt8S
g6E2ns3bXVkUNJ0j4Tb38U/YCwy1ZXGHVnp5vS03md1g3rO+H8r01hZA7byOQ9SIRCfs1rWuIsjY
+Tgeuj8x8om5mtKU9VKErolU1tZQlj1JrfvA9YxO7pTYrYjFSbrJmlIyOScLLeGu5LHkSCDsbP65
Q4t9reBs3oKCXwEALHOuQhlg7V8aarLJbhJLlW4/DEVNdvm12BTfIcJBIA2o5+5+V7gN1oP41M5c
Qqd1/XpiE7qxQq2eX1yjLeHns9ubLy/oIMUjrdSuuFRbXF6sa+KQDFpcIWY0F2uoUj1Ux/AsVmuq
paQ5aPpb6SlBZhPRpZbXcw3bvqr251BQ6r4LyRhyNfhBgMStcYVnH9d4j9jT6O7Wz3ZwSqlgvUxD
qaP4FbIkSITmz3a3XpR5Xoe9mGchQIA3K2iQB+vacv35KaFWaTJPoxMlzSLhtd6CdWcpM8FWRFXf
5WHYzK5Zjr8BnXBnLwu2nMMMwp/Uk6YtQwPyDo8DtVOarzZeAm59y3WbyqMNa3pqulDkXaWZirVl
fWbuU3T6y/K5fAHPl2a9kODVZVc0bFofwpJAk0Gaa5pEaEt1YZohCDbHRlH2HP62CS3J7IOrr/X9
eWEunEMFGLRFpnrp5XCyizq2hVs3DlJAQF9GdnBYO4YbV3QqPoIWjuqZRXWoSVBzYGrL/VfGLJbJ
N/Jt0Fyfw/O64aCmCDWwSBLWx+LW2iMZLyF9lvxAUG61xKwsOVCSLODbBnPntqxblknK3eAi8eDm
0aRAARhaRvmhXv0UOkkBOkhj1NhXrS8+ztNKZEtxbsM1bH4M1e+J7W5+eM26+PMxMIsoBHjMGBFV
AwazMw10oaRu74rv2YGdEHWqpuMyitgv+O0CMHnXXl4E8ktL5gXxhwERRHtIGxNDQPhqMA4SQYJJ
SGdkbAStpDZnuGt9cHQJpIIL0hCwtMZQjU9cWIlYAb2yEmLU9DfzFQ60vSv3Snnd2+rXyV6b+iIY
AHbP2u3KJJ8VFWcvmTfMb/MZp7BMCTZlu+OAEd+eekT4PkPzKmy6I6jBhgEWrgBnnPlxVLh9s+cm
Py2RnUFTs7f1k/0+P7JIoVBIoFPQBf5uG9NgxfqaCZiEljzFBIgtgrlPXiPC7mjeM3by+pQXU5Vh
ntz0vOhiCCnOld2kmC4bKDJIOQJi5jsXvHzWtYs3II0QlmPrnbba9HoLrMuqZsrpwB86HklIs7qJ
X38wqlm1w3KUwvCaYske/xjDBlKccWR1OVW9CWlb7UGYjVWSEsqtQBdovrpAfAvfrdM3+t4h4a2q
AQJiajk2QUa1C1ytiB3bkmlqEhbyJd04pkwkxEXaN6mhIhWuNbXk2DP5yz19tbvFBS7Kk94huJeQ
3r8Qj12fuEBpnQ/uX10dO4AiyNnWeHQkiop5eYVum1JghTGOmkjcT9/hVaLDo0QbL57xoEnix/hg
EZMbMSCWGpHZP1+7Ka1bnhzqlCNu0Q9p2CPUOlA3SUcZiuLDz3gEtjeB6iWP2P1diXCxq+ILsoFO
hRD/0m6y9DamoMZy+DbCP2A9JHAUiKJD31Dr5ZxT2ZVgpBDf0WeYaTnI9VzpxlQXb5vTosmZsaOh
jMqRMRczMfXQCe7QbSx0/dlO31Pn2Hwq11liJrH3p2umiPdptY+iJZ16PXvucnNhuybi+UXl6kjZ
zpL6KzKM51MDn2iMgNQqIyuNNyjbWv2JOPhUhXVKesd9HwwaX7al8LuqfJao5saCZLE5V5SsjU+Z
nMe6B5BENbPEzwEwk/ktB4XiWxD22tDIjjRTu3bhGZYL+4wTy5t3dN8Qej/GEzkXVpRhr88j0MvA
Oo7pjCx19EZ+jz49j1Bl6lfbDyjOV2ElaT8ixZgoNBvmpLtX279KIWwJgNb573ZBtw5n5fHgPTPy
M6EEKo8O5KGRuT86DndiSgpQ3C4/r97ChfJow3fcFeBCAc/f9MVbQVxPiuYwTYlexR3GVZJZexQL
NMH/t6UUtl0EfY5+qRhsjBk8a/gt5orPv0hD8zQDxsIO2EuanobkOCkGt/1IQJwiEct1HVil6MgI
3eraMzwnF/r67jw2rGZx6VGjkFVI37tTGR7TbQIdOZQdiq+T8wnfz4BK3zvsIjx+GdPhFwEvvuh2
bsGCVNiig90tNFjYiKCiPCyUkcEKEdbrFrlHAd7pTWFjEfYpAGxZ13yYot6mVDQV29wUZQNN79hr
N15NzceLqDelGN7Nyht/bxqdF/d3vwOf7g3pqaRK1CFl4M7gaDAbRz2c3eyRfn05bJVm2hD1qx0q
x2b+kkkCqFVkS4YMjH2qJdUwaQ9dGPJ0ia+Ltq7Vug0z7vLsSss5jC8V70YiSi6osdhbhpcBlYn5
5YCcSlPQ7E3hiRcMAK3//wHiMn/IEcRc9iV86vnv/twOVYBKO5YNZATLOlsvmEEzo2NzRYJRFrAm
Ix/Vr5m4ZHP+kBtSAeTbcfq+OgBbopkHlUTmVtcLkshxqc87r9zYqn8YxpBKl6SRHOz9BlrPNxl+
xj4bMm7m0FjhXikcX2fUkz6hKZrjajOrk6qZHtNNPuoAbFTiyirXOp6/jiv5+cWvFHY2kF3NlibZ
KfcITzCPEkp1mTDBZHDuLcb3XEQ7ZI8LMVelwtAgC4I7vuSagjlLsHjrQBkhNvnr8TE8pTODnDDG
kehVKfApZbCbAtzDlB3WO/78wyH5zI0QhHHgcwviZ85RJsxuOmmtOm2fjsokTVezwWvzTTc3ROba
A9pYI4KaTrplMrWcYpVzgLof5TAyW4MUy2HAGMQr6NFIIJGRD2rgN4x3x5lzh/VXuoe4hDjV56iV
L4I6CkJuTmfO1tAUs7HCDEXuf1jt0WGZSL/+zZycnuYV1LGhgX+yCK0DI34Y3nFM9h7TVXIQ2Ny4
8w09R4t2HXl2Cxi1W5ou3GPEQnLHMnwkSwFw2WNed3HNfW3zEfN4J35sBEKJLv5F2SkbL1ymQULm
Wpf8Rw3Gi0+MCKyNgVhdeKhlMFW9woXHGZ0Sb64WBzORRi27WH6YGMm4Fa1vFtcW0B3UXfRBx2aN
bW5rbQUYlAMhrY04mP1M2O76RjWKtDZwyyW4BNt4Je/qy1OsKx0ATDpTBi5oqEwXnetSF0K7oZRV
5tf7a+xFqHtA5Ibot8hvI4PSOVk6Bfqzfp6FAUznh0xVnNXgnuc021yhy6HDKlB40Q+MyKhQukhZ
Y2Kpt47X+/w2EgbfoynRlR2pXlsdjl9hgjpivNQJLY41iG9a5S1M/e1B6SYivJ+IA35gwbNtw5b1
Az3/OMC3T5PFl/djIVnKVaR65LkomEx6NeTNqAdvamewDfhUvq4UmPJmwnOhSbnqN0zdgjdWGld+
tbvLofgrI28cUkAgBBpU7QBZHHCigAeICg+uh3Ww6nXNHKGKLOqE+ytr8oHjL4XNMeg6bz9wN/YA
Wl+dm104JrDsArgt0TJiw3narUyh4oyxoPuLAMMEelTtZeOujyFEYPlPoJUiCoLnCDD+AI28rATh
IqKCnHYxlY2lcNShOQCaQY68y+vD1v55R4RNRx/xjRyJw6MbN9taG9aqlB+zwHB5W4Tmk3Jke+5j
UvkEsud1HX/AG8zEk4/PP2W2aR5JQ/CtazaP2G5Lpe0QIozMRyDzXI9zzrdHKLNdueamomQFhU95
kQY0fIWW+Z5Mp7ql26J41kyAUYzvQejGs/DfgI4BIyiQfePTUifzOFpde6lc6XiS4++Ds9sHpj1C
BHhPLrQqomg6ogV4ryoWOCo5bAaPBeTUR39CBmVR55RtB9TJrWSeagASwWi2YZ/Mg1ukT34IqGX1
cVN0NS/8/BKp9UxInqQbynOd+vpcrwrBGSgA1czcuQZEEF2XxKxn1OsbvbxjYo5fROnD2kUaSR8w
N4GcLoj9zNaKSsYvf2V0JAIscJx8vQfu1MqPkNTpdD6hceKw9DGLsLcw+JrjZZeSW0vq3QqnQry0
PHJ3SDZI4EfIsXt1683kjrlJfN6k/X1B8Zn9EINq8w+vvTV1llO9TH0eP1cxWohSPi2PaB+GfJmG
ZZfvgNjTd055PoHu1mYmUMXJi6ZaRNa3AmWZHtM3UqW9pKAzY0n/lcd2bUPal80HXVAXwEFSMw9x
UHq9qp3hgCKg9Jlyriuoa/5X7gF+YKe2Ta90MlsubnVn3DOjVRKo+wmR1JXqZwkhJTPO5v6cwzAq
LKx1JrXFtr/opwr2N0TqoxFhi8MT9iEzyKq2x/3W+a7Z+iR6HvIHRHXO2ZDY7FJWvUdS7TISNKSf
r+9tI5vXIYTcCTrUFTkFPZ3ctRS/z0aJlXi+hECQ+2YCnuN0h+9bd5yNOkFNsF6V97g6Z3CEqGak
xK1gVWpAxZvKLy2ghEx+Vhg8Oo7DpXm/r3tZ30YjF2OeiXWHjmgnkdrrfeHuGB5yO6IcYRMFYPDl
IPq3/VcBaGOQoc1c8126WFlNnFJFd9lwMaBSY1tJfjIZc0N8nXaxhjN6wWeqssgNwJW1AqbqKrby
9jX5HvKihY9E5ct+A+B/kRXQInxAYicx/O8JuckxWcKrXvNat1dr1ivlSo2L/MWYyxtwQTCk1qQo
SBr8ucXYq5tfXQPLSm1DGVBEI+byzCPZhBXUvMd7jODb1Sn86YJqTz5Fx5EOdD3/YDMuP/YrUpp7
xLIVW3FOrxsAwbySdUqt4hSJkhVW+eX/4ujjblumjt5SiMvdoxvq1qVq/IxD3a57Pa+ocBtvQtyB
tZmne1JW3BcFXHBCZA3njgzhMa4dTvVo9bRUJJpaoMqMEksRfMy6tStbVqYyKFvDrxKHYl3Z/hc2
pe1IV5xVwdAIwu7LA+mkI1VxC9biZC1ekz2eMo9S/xJ+RbUszCpew7v72PRsI67M45VHUSY77VQg
Tqpmsh+asquQKHHFjEFUWplkouebcly96s7d1w84NYFPR0N+klXHLKf7W1xeCyaTI7LPaVgEYRx+
mPqNSLenRunsDbqc7FbgRIVIrEOwGMRANeEfYxoMJSZsnhvya1eWFxr5jiJ8OG34Ph4YAONW+mna
Xi3+q3e/nWBI5UikDpTt/QG0FFpRIPeVuhlNN2LYXhH5m7j89WmyzPCA9rREWDJPNoykB7/I/bb7
RVbupHpcHQZf7DSY1sDttPIldJ3qN+mmYG8lNI5s8b3ufJYd89LveqgTEBvnIavV7Ado4mFlBiuj
4XSvn+MaJeapnFoXU9fnUH2wDCafmSboYEsu1SmloCuCyyUlTq168vtl41Y1arwUr6ADAJ1+qQHt
PzUfSX/uJiZo2JT3iPhV1OeljrkowvjLPhgn9MTEHmBawWUQKkejzV5A6sNQOGBdrBcREweKMAZw
fv35EKsd19wCU9yc4t+8/2spUbiTcWxRJER6fSL920TKYbjUd5wfi5AD3PaaXONcBnjm9GjY1Fq8
S2Qm/+ooIOPpfpaatOTeRpBTm1PpcB46TRuxLOBR0prFQ4l1wYVYg7cs4Xup7awCDLZyfdYiTqbj
QQ0F7lN8fxJHSA4++Vkwtkdizc2daz6yEK5NWhulAA7z/kVTd3d7pmqxMh710Uft273+esbRKEWU
vlPj2gvpws2Q0C4twfyWbETxZEoYrmPxKrb9uCp6eoH7B0+Ak+YyOxF30cACizSO2dxfdcoMwJoC
zV7CiYFC2vEXOkIo9cUwzewgjinaXwhD0nA9SGxKJ2d/PmNHl9iIwFIgn6432S9L169qBkQ4JSTY
BD9eRDB3PH5/zIGQUxPw6UPx/Oxt5qUlMGHbCb6yXRtgo38qqCQU546OmpBFfEQzM67TGupQEpsL
a5ufg09fOmdzq1EeaAr/t87TlrkPUzB13BaxDM6lpmuIb38DRZQSyhNmULcnYDYRvw1vbp08mv1d
NQaE1nYztc64o5JAter722GZOUOWm3T7Iwer/8dghGExnI/7t6qWFAVkZH2SDDVbiv8WDGjEp6GK
nleXvhgrQW3PF98DC7iKeeswfuKhBOPKPiMGWv3S81QaCm2GeCcusmCEVTnAvUd3pr1kkAbO8Rec
m/m8LHaoQr+6YJPkvUFV0/UZWKqi4NgxQWfDJAYIlhmU5ug5zqEjwI+lASoGAhxafpoYBbYEqpaK
wF6gXNp5+ivAiEHv0QU2lKDVHqKHuBfJ5W03xDKb8RSlCW8LcDjFcBwCfTclgQH9ukwYCqzZK1jj
V5iNkFmZBMrWyd5VH1TbYt0NUFVgeBHX8sv0OWBp+3NJWP6Jj5l79DXBY1ivJfIeJvCbRJs6Wij4
5E7wN+9t5YHy+Z7gN88QZmACOWOG/UyORe92r1KMI33CUruVSRSdA0DQQwZbOxEIaEO/BtoEKH5v
Zrxhakw0chJ45xr8dfqiOLekkgyp3J1yh+YwU+GZ/O31uvVnttL9jJDF/mMRpV+s7CSX6hYZkkXb
DnBGZ+eHgHsqICIQKWqqLqX4R/hQznz40+U1JTuS40tl0TXRWNMuLbGlvQJzgEja7Nx1Qj0VdoSQ
Tdaxp8qf2P5WbhfxaJga1xg7no+96FaeTLDv4p46zc6/1Ksr3KlZPMWTe6DwG4J0tdi2EYafKgT1
OVAGSJ8wDP3gqyK4IKzVMi29trPy/Pg2ikOMAcUnj0lhUEyi1BRYuR3Qu22CKDgSfnU8vsDgeb70
L6adZ1KeS3TECLymTIfBAk9nFOM8Wc8CsZGKkllQOhNVqP6SmA2DT4eieteVziH8WBi9MJdVChiK
GvspU1kZ+CGNryE0qYGlkQblUjuatb903m3Q/XC/YAPQ+o6yoNiJAIBXOpsrgVOPylE3UYorMnBz
zM7omNsFz18F5VjhDIgG7bZ8dIQk+phIhnxj7CDqR49/eyIUeHhdqu6Yg7AnaHiCwmE7fkJ7yT4V
qwWzza1kw5C9TwBSuYXXrjqv/9Y5p0Kb5y7fT11U4Pw4v7FmgQ/sxhUjEE3cuZsU8QOKhaRAXGmW
QJOvdrfUIBKMZYAo5ygIdFFbMzPsAf8kZJb6+ijmbDytgNN4icGK+kbDr7yz6ZraCADpPlgWlkWa
vn+EBL0vyli4C92FtEpQYcg3J86aOHk9mL1AyNIl7mAMljBU5v3H4vVFGdHkZ4vKh3zctDIrsxEG
gie1uGb2qcQax5sPwVeHsJ1dfSCugPL/FacmC7cfDQNUHO6PWuaKHg45+6GLgB7v5Y5DUZdc0LhF
IdZVsA6Epno/cYrfkh5bFx1IQhS4QK+2mmH4Y/VJsxOtEBegp+CqJgDcBTv523nA9XUOEwS+HP3G
l7HR7ZLXR6XAa3/kN8ld5khLZn4e3RZxEEzNyrL2Q27D2n4vLI0GJV/BMBDDpJzcAKAflheckqK0
LDraRaqDnXaOEZEElbOoSHQEk0FSQ/ok4f7+c0Il9FxUddaFpXXa8GCrhUGkpVtIZ/xVpwkCoPA+
O9lIQwF/xsj42bknCSa5MCaRw18v8+ev1odptlp7gNXh4YARjCE78ZJlT8TeFoPD0ccxz+X7ypOv
xaQ0q5ul/3rXNP5IYGowPwdEbKUGDJocaT5Tify8JsiYuDcAykslz1hwZe/fLpik3E7Ko/7xvqaU
t3NvmtRzjOnCSbovI2Iw6Vk6k++DnCxQsdvsayPC5oFnPGrjMbFILOXeWfk2QsfjEAbFEHYB51yD
vWha1Hm44cWZ5u2QMQOUsSnVBSEnPDjKtfULE/QjmxDbWu4LjU9719M1ZhOcsU4lV0v5eiT9lUvr
YoHVSM+glQW8jP/ttx1uEshOefBkdLmee2pC7TR1LAiu7d6QpOYiIYMf7X2Xe9hNc1u4ZjZholSN
m5bDqMPTrxQSXbcOdGq81kDgnOXzmqQalRRoVBJV0wBp5QNNSYbNODuxqgipiN78oPSZXqUAne6w
eSo+TJnQqw5L9SRuhxIY3TwbVKlDaOmgytWr1fdLkfgw0NXCEvvHXVBuBodiL568tKPh/ETW02+E
E/mhDmQRLvTZqDBjmp132wP4/M3djJD8v33hiqW0GoQxmGKSzEIINXUI/hHxNXTbaPGJf33z35Vz
FsXRvM2TshZwD96aUBd1yEPTg4fleOv2bgNhbpmn+WYCJ5YkiB8m/Ky/t4YvvYh3Rn2RpyKE8q0E
ZDq466YqcrnRBRnMujVSvIIVoH97oSwg5xVbWIfgzkFPyv4jG0hdbUHp2S9FYh3nagpKVeSosUN9
2oTMhddtZW/+eWUTQpqIZQ9N6nWfeIFGHItuhcRtXfR+twXCtZU6bDBs2k+YejiR5Y/BcxzEPHgE
Cuggcwp9qUTf5j+aNxcF5HW3TVPNhcIAKceGCbdqRzBEoMJ6YP80sOyXch2pi7lUMBEf+fkhKGkj
2AmlE2k8QJO98f+rqBo8vYxjxw5s+K08Kf4f0oKuOfNdSTIUvFu/HkDvxg+gD3RMVZgXM7DkICTQ
UX09CsLoojnmwLyaPIQKjMiXfAISyBBFzLeVh6VteXnqbQo1sJHxtXqUlTl9kcu1BwgMHpLQPzx5
2aOIwxwe0qutqLCl5J0qMovE9i2MNk87G0+sKgWOQKRLufPlWPcd66G+MG+ZGwdNcpiPQAmDLeAY
qxvLhbfkNg72ejrOAOHuc85U/P0g0gt8U1wEIRGcBGuhhXVpAmqRHYuqYkojyWJNfBhT9/GTeVO+
x5DKs1dP+y3Q3ZdjvweK1i74pX8+N13Tl4ybUvuSJhmNsqkQy1QA67Hm6MmrUESldBiBYmdj8bwT
wPcqAcCPjcc0/YQOQ1eO9J7zYuEwX8IYkPzE2xwjYmE3VNkByh/rKhgQaoKbtzeqOloYhbHX1t5z
BaIzKEIdXZZ7fyWxXP0Ax1AnSYQI6iLiEcuZKGKx1syhq3PHFlgc+xYdf/WI2aHQWFok5XcKC6Mz
o/Iyzcx7hPH0ZvgFz7PzJOoZ/6A0oQB/GTg7puqM88xgqWmbI2D8F1JIdszhTMsWYV/4D+nP4NDJ
Le2Uj+5zvL9it9Dz/5wFSwI18mjP1oLXb+bMU2eiB8tZFCYvepDfHV8U5PIO9H+ZIt7DrXiZ8N5o
5Ii/AFh79P+zBBRm3WYFUH/d0j71680ePVb28ExigtnRa/2zGmO3r9J8M2OX3tiVZ2QPeFPm3nfA
FNX4Mou/MbGqE8X5zDZT+9g6whdgHw/BrR0Os6kjeOk5f+WLcd4wgLZm04Hd2AG0gecw+Xvc/Qqk
XJeRm1YdFIwghxdX433GFnNa5BgyTKMQ+9FUmfFqsSWBePN0BaxCtFCGsOwWlZlJqqM5JbyMfZne
ZQ72MBztKK39gQo05LO6Sj5rEB/4xjLQcPVU8foXJPfMWtxQI1402egWjQW84SOmsq2HXaOtC+67
tqdVsO0IVcphffNBcS3Eb2h4BvB7/VRmLwQnmUWZ8mlTfIzfy7NhKYoE4AkBKzFPDUeiSuzmrU5P
0n/3qIdAPkgKNFfnupldfCH7S41YAX8xT+e4XD9rY+iblcgP/Nj4/vI1m1/2hpBfA0iAoh8qTr/O
04v6BBZLvbEsfIeRqfpyH8cq+gN3R8U4ejtwu6Mh5PJPnJOmFV/X6Fq/h0Daru8VoLS0O5p+x71w
ZZvnrFssEX8cHrIV8p/doTZoH6XvJvD7K2clCWZNJhP51iCIGA9d2WdEI4jsmlqg6T7L7ZIGUrTg
0M84Vgtt6ig6zLoMOkln+lMvmb7NUQlCNCmYbqSD7vAhWtpM7rj5we7HkTH2gRCGZnWGK+BGe2CJ
3q+58OVttQtPt2sla7h/I3sBzydRxtR7KZ4d9fAo4OGttd2gWIsiGL9DulRvbKATPSfoaWV2o67f
JV8JXIxYE9TWXFGCwdxoVcmXlVw5gqebCiVl5F7/yBxdDDnDpjbI8nSTpzq2OVmKd7NnIcwY4GB2
PeHh3frob0LYzXKYUXA4265uvlQ6K98bxMY6p+9yWZjTUTUiD8/GrF96roohxMQz7n6jsqI5YwCM
POuAjq47i37cZg0hW3rFwsF+yjkMJwikgh0/5qhzGORzFqh4J31awBFxLwiUXjFX+caGMSXiEe46
GKABgdfAHlNV9N2wjvPnz95ZT56meluvWF/6XSzZK9gAtFkEwJnVqpgG1RuuYdFokSK9vUER09vS
AWxho7jqEOdZAYpDFmkwOtlxX3H8Sxd+Ld8LVHLsZuyanP7Un5YYB5cWRG4wmbaR5zEdrhN1LTWC
EP7wd/yTkinMQk2kH9OaaNwqkWPtzj+qi61/SnEM8w2INDWcx4usYBFioiRRzVv6yxJRsqPXta3h
LRHI4pAWxX0bhzg4vParySfVisyo3gpdoDn5oeLGtgtJzLKatvsH3jTrZgQNzAXAsodWw0Cy+Cem
3SMKIazk7W12SY1ND5UXLBpbRTx8WIz6XS/Lg5nnt9d5WW9OrgJLf/Kuh8N7XBMLfIQigEcvQpXh
BulIau7Ep3rFGwgMBsJEWtOhlCkmHt4pwwORFL7FzyvT3ImWD+jMN4tYnlo/5AAC0RkgEjbEX6we
+nZyBk4YO7RSr5hYUmWMMRzX7d1hp5i1a0NUqxNe9ifphRbnJswpQvkSe2/XYcoDjj/ElpaDhp2y
FqH132834Dix1AJbO9IUyfU2Q0mGYXhSHNN3KlkFphltb8CaXsWzL2FvDwcBpfvgwGbUGkI4iGn2
yb2H5UsxcagXTQF+tTRJr/JT2IYiUrlxw6B5KXH5MRhAuTkSjIUQG4vsnqYzCXAOUAat48+JKU2e
umwdKd1izzqeam45NOIXNiTcoZn1z04hXO86V3TSF8JRw/MTnezv6nBL/rcciOGc5IRtuZFKCue4
JAVZgaTt3PURJS3nTf4u2F0XqQCn82pfjsf8ZST+sLX5OzdBuRVwwVOYoZXJGgFvgQRrwJMLODWJ
nwyD8k8mllkj+iZGCps0xt69AnGHTGh3b13DmBiADGcM7hmDIIwcrR7uK/G7vQpoJH0Q6pazzTIK
VDW09OiPpuNFLhObEK/ouig4lKtag08RV6XhefWTuvUYksSotMsgpFdXhKep9pUiWypGkzt0HWf2
ITRcfOPrv+i9MW/cD1+9Hnxfg2nhvukOoAuND52otiRxMBBzKq1lffwA32dV7gESm4Fcxe4edma/
TTQ0YdqsanPp+fuG3wqk6YQpyOoRdwzKWzaxuOEfWmBvgUY9fu7ayRPp04Cd20VWqSQstKmgaIIf
pIhk8IVBH8+A48G5r5B4wy7+EE7aHtIqGSvQHeUEnYwhEEQr9b7vB+OB393rFExMBfQNzaA85MPF
6IGcX/p+t05c0HIvrmn13S0BmBm8xNwZYxO8QViiyYsMyvEMh36uq0osEel4LjQGW332eCfbdV++
qnO2I9s2ORgszeIfkxtGopbI1ALvOOdGOj7Nirn4pT5WNTdfz9UjF1MrydwbUONR4rKactOOCpSz
LwzZR2NWivV0HHDdMAiAdullb50zEWDi5ngViWhi7Eua5IgKEnvVAB3F8MVAAcP+IdBIHb2/xd+H
n10WQe11AmCGMUObt+lVTn6fE3mjvSVfiDqUzREhy9rmrrJueZsC38UOUQLNxnF2v0+WAoXGSm+2
WtVgvlTL9Okn5xfOCx2Pb2wmMzwKE/T+L/fJKsreUHINqZH61kRnGRZQT9iGLuOgz/1WFjsuMmHR
KUMzkD8Odm9WtFw7Pxb/TcBGdKplMI66D0MVef3qO2MbNSVDahtjzw9TXUDvQ0mELyH0/tBQ+oLA
JE9eMK3qfoR2cgy+AIG27d5Sb3MKndi3Y01UFnY6kh0JDP0QGQjFyBFq0th2g/Aycev6laxfE7As
u8Td0z+Cumq2vKBTHhQnahGXPDsC0sfr51dXHGBTh9QTuZMhU6xt39MkmM6rJ/EDsHJiNEEz0xam
C1xn8O8EMD7mAkEjtTYS9QORo3QFRh5ZD4Nnl7eaqALWFlILkk/6L8FQHgijEqnlb4tKlhVNtRwE
9/zzGnem8I8kijB1IU0/Ov8kpIgTCoql9VPRuiBhNKst9k1JdEttntbB6KC3/MdcyMLtdEtxJ7vb
E6Is2HiT+JBLl26qSUVW5gJZcLcrI5CM0W97zD24VakMNezlKTZU1qUQGaxmA7Ibdx/AQf4aBGED
I09Cv5VeZgSMzCP3blZEUNPM7ZxfS3TBqoY6fGm5JLTGFtAI0nu8PANCx3tQVUSk10gA/EwuNtK7
BbXpjEcG7G0RNFc/Ri6sJKTgkaHnZTfvhAcT2OvctiQL0+Oc5kn6x//6QXH2w53P9cM52WJN93RZ
fSKmskrnGNWdN8anDgxIN/328dX35Smio0+5Xf0HhbLIkq9fUCi+IW2MaAZBKEicdFyiXcuAmmgb
0TnINwAo618Rwx+aTSJm9ovfZ1WaYIiVk3kyXR8+iVO3UQHA6ZL8FjibKonpTckt5cPnSGjtLpqR
boO2SI2H80Qf1er5xa77kbhdWalJMciJZ++YP4y5E2zYfQeXQeNzER6KOg5CbyuPdy9yjfiHDRma
uZS9B2y9BFmKMTQN3KVsDQoaO1+7uJKONiVUwrKTk5RlbRw3iz7iTJqS27BnlqOx5L31OOIgAh1f
ezkQOIS9dz+yCp+DiBXyMoxJ9JeoXQvc8Uy7ajEf1+9xQpbaT6jGSl3r0V4s7ZWhVzuQYdhDHSZN
eCmzsjl6NNTrg86uk8cR3D5QnyE587qpYhH+mdUCZtwUhjVIa8xKXxE18IcDF6LVjp0TZVPklD03
9Qqtt/c9NQ8FJhnk40zqBGGe6C+TOk7+fSwtgRDzE6t7db8sJHTay5OSo9BnpC/K7MA5BLNjMWmS
V9WRK6at4bt2i/x1ZVho9BKRGWJ0ShlPPJEQPRXXXEfuDirOOQ7AqCN50Ilvs5vgPV8drQlH7OYI
d0GTWR2xLwpGsTjMtP+Et8K0xQSf8mtLO8NkbHGvI1V7bH61Dp9D7W/pTcihrL/LCURjG/rWHLKJ
5KvWWP9K1kSwxtl68l0djLbaPj8uRqymSiekQyWRVpGg0nudWXwR0zMM0RdQ/Qqeg2iqhsl5hmkM
Vg1T5imseVTMSXjrmlmKXF2KTvE1wXjqptOq/atLr2tQlN4HgP5m2RyCLVCyi6tfK+C03ApEGfKp
ASTAaNyIUoAl3ZGx1QHWQxzzlQQmJa1inExQj0bOGPfY4p9oijmczcpsu375JdAAL4xKhH5HUnLL
h6Cho+5BR0l1PzaIz5nSgUpbMSNNOx4C282oSjBJzU9I0R0JjUAC4xEnfYXWZXfC7z+Vr7O1pkJO
TrTHY34c+Lymbe9Xb4K85DJjQPdqde291o8gN49BKfBKq/3BkCYJup3tSB7viJ0nMZ4lgv0YjOHW
v43BXp7lL/RpMTKuTsGtOlhhadR1OPfKRHs+xloUuO0iMrKjFgPOfDvoc9axK5WROR2khkzTOfpa
QgkvE5r/uf9Fls8eYfBa1MGpULRPbfiuFImBOiegZC493mlcfBupTAEU0Vi+s8uxU/jTwSAGpcK2
+Jf3t+EeYc4ILdtC6fp9O5LJOKKhhq+Y1hAls1kxmcG2MYhZgunP8PtOJvK/JY6kbZf6xuBNSg49
+4x4w7fLalW9yvdvq019RiL6tT6Oe1MI/kDYDdij9qwsido6I57WZMqZAKAayQ3XmGjMvgryYAFs
VhErnvw4C+RE5dXuZZE4TJJ9Y23OD+PMaX+fS4zVG0EK0xY0+MdPXPB/97rAQJWRp9GAoFrbju1f
ye9mMStPHHQGzoNhqVMUBkxOF4st6A3ii/PM3aAAwTGo6X059OMtP4lCqzw8kqzZ5RrdW+CGcA2z
dWMUMx21DjkAD0uVGXUgggfDoFTzNXq0s7dbQ/YTzkUA4hzfx4xMErUGuNeFU9b96Ag1odkLRVzh
Q/neOr0V70fsDsGawXZJfsA2vRmXSLqanVhiw48eJNuUkZw/XnTmem0TV+FMcSwKnNL0ErsJcU6n
HQVzc990giC1cOzShxEGtAfzNWMv4fS1ZYKjIo4yRfiivRPiBz5XOQgBKNPii1Vk+bCfgEnUaJKb
r19S5rwU5b17VPkhzC48moPpOrkI3VyGVdbWpN0157XivvP4lEekXDO6UEOUSHsL1UEp/LREBFfG
Qyy0Tq5CElAnzlJFHMpDhdQNUXR3XkgEUcSFeCMV1WcHnveqsf6ViMPtJJD1bmaHhuToOo0GJKyJ
b1jgXmA59MODMYxc6PH1y1SJALRJvETQ7Tf5E0cNZJj1H1ZjQWG+LxAUR97Oo3zTE8XfhKcKYiwJ
olX7PoA0lF5PA+PIKbQMRcTQ6uDSHP7vDNMoGBzeopAoiaRHo3Vba99bIYeLPDFG0iwKxbOUNrDL
B7XfdsqcWPguBqOrdqehjzDhfxNjEbRkO35YpAbB5QToej+ef/M2ampofbaabCw8MdGDu6uNKFAt
5t5wDJ+SRCzx+bJyRyS7Dezy3ESLanyr/JaNsPtb7dHIgnCFF0mhCpo7qcyyFZ+Rs7OavYYVmeRn
xpUYlABni/NCaGUpE/bRZkFxbbahEVb2jOSZpYrYdcUi6ARWp2ID7TRM8/hfxz6uVxRQaTTGwndz
BuQ8bh3yYlDjgLhDbzgfLdMwYKPuhvT8DlR/S1xpVJR/ZZ/BSHk2uPTDSnEcYZ1QlieHXmbZ4bB9
HyhVz4lYxV4OPtZYwR70T386+e/YgJeViHYjYiqbpKTcsbctJOW0Hv5ar/03gBivRCa0i6YWBCQb
MhSxekkT8l65iKjz5U5667GG6ewbLy2+fzHsVaN1KrT+G9Wz0RXeNu96cRPsbCgbrfRCbeALDoir
SJn4aZgERZ/0ZOilAaiN9242ag2cGE/1stinmdhHD7X6K243mb6IyzTgu18DC0bMw8zZWhpcJaRP
Y5+GjcIEMt0iQaiLOeQJbUFL1Pmq17PElSz5Q6PWcSKILK9wFhFo54QQAWi3vASJyljHURKogWzm
y3TMXBJKZGaDZLoPZFPslPrhLZsleaxslMcNl53y1IRRgEgyYAbxIgTe21oc5L8O3FSWZCv3jLQq
AvCPnnMIBNbVEpuuViiTInLKkswOg79aXNheD447zw+L1B6MDfhm3cIzR11lkLLAnG4bGz1SvPfF
asrwmnl6s9IxmlS9rfjg1i6p8ZpsXLplzMOHtbkJb9CavbyC82vnZ6rZa2YFWqjMtfc4l3PTYnZ6
7SxxUMzleaEGh23+YwVk3V6N6gajy9rZ7GkHZNM4lunopYZQslYEUOdVGzE2/hORvSNnQpRFdzHR
FznPpXDmrOEgMa5MgH+YslOJ0RMUlfhanfn6j766uC3ABHzxuVUZLKmb2mHyafNMc1B+Xcz1TyBH
nhkZGtj6Cys0A9HF7+PUhkVFL02CTGEsQsQnUew4UGE/T+RKIVGZxvY6IaY+87qU/2iYyJwkQ8JY
9toUAa2J4BLAOBV+IK0vsprRu+OJqmdFs0iteC1s2CrlvpjPfzIgXMgGGaoh/jqG3dZAqJarOV6E
ghQHg0OEB+tj1VBP/btbU8+GM+Qbw+EHhZK7GnBvbCcU8H3aD3SdQg9mcaeRcvWE/BYZZrZTQqRF
6RSwqRSyI92wrgg9JtwvhxqOtZreUEu4/fRsaLLG0Bez0SfaMao29r2jhjK9ba6SFGZxXa32dUrz
n1EOt2K9uHvKnb1/Dzle8a+Bab9Nw+vIrKllI9DcHfbFHUAUC7nzE3MVVA0yCc8b4JTqRTJDGqTp
jllgM9PDk7QI4pjgKDTfnXgBjqdKnNuGDaqMqR/gY3aTFwjQh/NOFyG4WUxwP0oYEHp98TVB93Z5
VUCaia3+ixN/zoHCZRtSyaa97Tg/gcz+F8yDPowtWB9iS8m0p/iu+C2ops1AwJ6v/V2rBnThHDQ1
Szj+H8cERmQ60HordFeJtsqy4m4uEY/fC6vqkIcPvE86kKGoTv0Rm4USPm367ilVp6mo44RpaLyp
EG4JsiUbefkP8RRgkS+lFY6HJUKyqy6aQmXeaC2YdT85qwcV2a483AI6DthsZRpVQa9sULZbtaME
3TbhNTYWEfuAGCVh8dVatTke5WqrYBKrYweh+2qgbrJxo7w/dQAOLAwfqBpO8+8rnMXuEGIDSn8M
wTKbWNFI1OpCjVFj4JznB6r6sXbbCaRd/d1pE8Q+1PicbBIGvtCd1O0jKuYEtRwZf2EgasXmtiC6
DPSCjDL2qnIbOzZOKNRerRLt3qezq9WIj9Mn88ZDUkmUEsQJXlt+qBKpWbrrc6E8KS3EwnushpzW
YjCmnw6PvcxaIvTxAUAKcs2XtbKb358z6uThXCjW40f/9mNbIag2vwzQdyPpDFGAHJkP+PvzD0dn
I5H107uUo2Gyz8hq//BENNGIlR3LWVQOffY4IbtAgyG0ymf+d02CtalArm2TAF5t/ve0LQx7B8YY
Mo/9F2RCfBGhXoTBMq+auvNhTVy80sIgg9jyR9IW86P147UgmfCPtGdYA+UIQp8WpEmK812QbT+k
tNZkTHmvL9UjeWSQ0mfnzSmg3q8H9ED2c1Ii54JAmoys7OMtL+6G0siQDU1Cm1ssYhLqULH5r2Dv
3yrkSCXyDQP7cXcMqjHKxJkIP7YxkgRWxgloXbqE1SqMRrlA5/AI5sAdFQPUjfYOzGAGbQ/1Ehom
zsuFN/U5cyzXfcUI2tXnJAIFmoLGDVMy4t6UxVUu0T5DPZzhSZ40acs7DXDa6dPORrXYHOPL+THl
zt6ayGClVVDzUse6IpQM2pbn/XE+pxNprLc0BCBhQ9GcFcnGcNskyQS4iWB6Lmf9QrSb2+Ckf6bA
zqzQdSilJx4VFa1AvTmTFIg4S0rtk9Hck8GAOLLSzbk0rAa0R0ySBp5InPQVQeQUynGss1RCRxM1
1PHj9A+Opx2vpE9I0tbTPjFaw39gc4miFf9+MVQ1r66e8Sm7NXGuz3+lDu6MmxTCSFH7PYQ1KZvC
ZMCtH5aj2Q7m5U+MN1V5WSZ9ZPeVJahPOlCePC41yMs9uF/DY0lvgLkAPNeiGpNs1IAdgosUgU/3
L2eQBroyu/x3sxskzBvK5kPnqH1YgY4BSeNi0ozxh4pueKzP1T4m0hdFmwxyd4kasNzUZRWLHLLB
kQtI/HYq41zWpsAUOP8jH8LqG2gaGX4L6U6Yl/KFEzpJtge2cvwSec4nxMaS7XcOAazfBqDx0rr8
mHqLYeaUx7QcHH6qMU2LEUL5I6AxlMcup6SjCNGZucde6VfgZ8afJSYu9wi9Nxtn5ksH4CnGap+s
wOxMBYvUMbBv8Y2Gg9O1Lalr8nLkDdB+qUHVpeaHJFKH9F8DrbBkgSJF6d3tYxbRQabKG6/uVvHU
Yvyoco7VXyiAhFaW1rb0/3zXhQiB0M/qghVIwNjCEX9OC8Ky6W4yFbWd1JFymVGy7o7RolEDKzBA
+BITzcanZk42vmqLS0pUzo7VNDyiDEUCfRtA6hG5pBdOjhnHl4NzQWZqCoi09bkAj4m8HAANubKN
dqHMv7MvWtLdLWosWCaMYme3/8ED0qaPnbYv3gt2q0PMyTPqpYCvbf5Gce/zvACM4lCvwVFWxR0W
krzFI3Epe4udVRv4bRIWF7U+tJ7E7TINZFq7pEReZYf5D3oO1hDD3UOrCZDp/zjaGiviPAcC4kQM
FQBib/wwggLSjPxnX7IxqX7YoFFud6zFZ5LHlDE0ZCgmsDW+/n6mUi27hcgiSSmE8UQATQqw8gSZ
bzKGF2FAF5lhwNXlqj8S/jUzLE1Yplm8T9q9DGgPhVzRwzGSzXFMvdxNqW/OjBsnDFe9Dxj7cx2w
q1bG8bzd99bhZRaFqGH3xvlgha0tXlpRS70zqpjSKMA5YvHn3kb6V7V/Qvz9iVTpssu39uvJXxx1
A/PBdx20D4tTOxCRXkX92NeUwrwu/s5L05JMtN7CCZW9HgnLGlKudW2ZRuDVN2l2+BvoEyeLMHiq
ZHJNXt8nN77h77g87InYD2gpHab4IHrdS8Jy7r92D+pU+t302IfhFKCseHEt3HGvGKnIpBnir4te
k618rngMw3pRxbrkLbg+/4XUK45Ylgm4gFy3vwmK88YojqxVLSTIZxousJvzg57NHXm1nbiP6was
s0Xfn/v3YCohvHRz/1BjTPA5bOP861t+CKe0ZbGf2RlQ/uZxGOcg3i1hwaLdPghgVoMOIzv160wl
pNw9m8e/ljd+WnEU0cW2b4r+a7b+9S43gsskiFX5xkOPiTUtKjdeB/SmlAGwK6dLwI6+aZp1MKQx
SpT2SpDrKeXWr3qo6VgvFUCvl1pr8qoSN1Ea38K6tPg90paN3nCQp2FMJIDqZIF2g98TLZzauJCW
jmX6tCQza/vFGST3cyctgVACviau5UjS4G4+Sel7gnVwpRtR30sychd9D5sHEyywg5Zb0qVgIqSW
YkwXfscnM+ep41XzDB+PO2bnhkKaBF9tDiZ38T83vTyXYuqH8B6sHWa8xyMjx9K1JFTYJ2ihe1Tv
/t3q4f/RhpnUGcG+tDGJoiEOXxjimRIhNdx/r1HyQF6UFczwnGgKOsAb7ODYY8UspFN4QZwCq8LW
iPuiTiH7d6LOQIA2erOXigu4sYiQUxrSAi8C6ARKRZ0uPs+OSd0AatVfmSscz6iTlUBjYZLH66MM
VPUoWbFz3QNckB5SinwSOlY/xb4+/b2kIev7l0Vj2Bwzb5YG6OaCHd2i1bhwAyHKp/UsF213h8ku
qTOdbShk7vLqdtHVFg+AmQOCgl8AYLPERYL8t9uD3kfGjm/VJaUClyunJjGXJUtznRvSIE2IjsVY
qxbkm7pIdN0yUh6w2pQ609MKULdEaGgw5PJHfGdGPMY+h0T57sfYCJOKT6aD2wPuyqZTY55V4ASW
NIZYnBwKKhjt+xCxRVpnxeIlDIWuaWZ6wTTGgiE7el2I/c/XWsN8OQ0Y5aBLVTgN3E7DIG5AWohd
UuhbxFOqN8SXor4xKm4FBwlesEi14fN6Mcgn2JL/0xHRP/5HIQdoB2SnRaEcv/eZO518yB5vXSbC
NWkdKE/kKBTTx9nVBvpECZ/lu2EAEPGv9dsAVujLvx2FhiZG3YlI2SK6ncjsVMb15FeB79s47cyF
YSlt9eyKDI/wL6clsG26Qkbb0LYiiC5oHgNvHB+CxTOr1dNt4QbYy1LemFHC6AC3HDOpwairJlcQ
H7FiYyGVmUoq142BXN1PfNeqR6aMM2nI/QZg5LBPYWWZr3MjWw1gBrR3gJNganh20qUIsZSHwUsN
AYJEqxfr3Cmk8424Ev0dtBGJZv8aJr9iApshKwSIsRxXrEZA11W8KZhBc57dlHumGn+ZXG5b+Jmb
eLy+6EPNe8cr1QxRVmZdYw/TBjy3pVOSxCqKE/E1qoZ8AS9lmjK+D+W/aKEXXZQPHNZwKfp6cXGI
xU3btlZqsoKQofHXqbTterStSR34l2rIZaQdc6mNIm6NSStqFmKRB7gge5rzQi78UNZrTa1Wb4Pv
MEkvvNQX+tupD8nol+rX5D3toYSKE82hl+qFKcOCJlyx/q3VEHOA45TLg/JLmbuIM/KZh0yQKY0H
U0floMZsLgjpfhNG8InTSD8XB2Ln2U/bE5j2yGcRVKDyz17oiYPjIXsiaPbzXJ3kWFMeah8Lt6gK
wBpmr6mP8j7oXzv2E2czVdPAOA0NzHst0Er3uV+I9fgvuF51bh+lWLifsLIjuOD6OYMyV7kmf9ik
Hg2pyTsKAE/2NLzcfWPOkLqDBnq11ScqYZ2bdrT8z40iHbhyOiNLIj7gy2kHuoU2UMPG2aqvawbD
Hi94LXi0fqHm+8LwsTVObd5GXOe67taqGUNmR/uG+4aQ39m6Lfv+5EodHCCgR8L/YND/kPyoL2J2
chbKVtV0vmcQ4t3yErO8nR2s7DKwaf/wY3NA0RrO8K4vUbQ6eaJ0tJ5A+hQQnLilv10xUaGuP3zk
S1Z8dRqGuZq9mz9NiJgGbvZ01DpdBVs11XufF1jvvkiuSIb2cotRK46tVZ4WZfwoFRUh0YQsYbi6
2IxfEiSGs1vT2NavAALLS0AnjV+E0rcgxC98r4E2VzORTfrjW+Y0NjlM/zfEtgwYy7QjNHNAc7Tt
P2Yeu0Q61EBIDo5T9k5zZqou8YZ//AoIldFYwDwIy8HR5rnryNMxjgb7cJ2EgwunFgWE3AIG+mgr
nJNJ/SMujm/tYlLuPgnWbfTRn1nqeZwFzg4kwYigUMPLKcI9Egykwo/cXD+8tpfNOc+n+24J3Nal
CoGB9S2R2gai2lEvHJLs2eXQ/10psyz8HhZOjl17B3Qq9qTqVaMivl77mYbMr/mUpwYwWxn5TSok
pgDBfnSiuJB6Z4MUgAFcEPObpyhWR4+WIWNhz8AZ5w2xfP+2IWv3wEv4exTazU2qYALv25cnVJga
nbYokNOH2cL587jt/gLq+pIPiQbmXhGEklVAyphyZhYosscRGdpKzIb9nxLrsW6smG+CZqkO9/sw
cLuLiTigbJCFZldKQWMyIMnc5f4+1x8cgER+S7IjAP/Q2ejg4dJwCjOKgcFZ3IphL3rhGDs45Dke
SUgfRsDvwvKACzlOwXQhu173WEiUT2aAJnZR1fx+5IWIRuu9We+LzaDElE05DbjcGj4zziHgayN4
ojrUEKSlkqhTZ3XsoSFvIaX1pGe9opqFif498KnIeFM3LYxyTosXEWGKR/DZgvE0xnQHIOrDprR2
RrRT7JxQzMvkeFWGu3aRpU6rQDkSLaJSc8HhJOuyU7vokt0vHOQvBQgBbGRexqeK1n9kpQ7fuR7U
7s2ZvL8O+GdPbvJd7xsUhGhIYbQYyR1pj/Tw4LIuI1LIeFgSq0o6Wb2jsAbDU3b93dLYn/zMcjnL
/N1YcQy4sTsk3gVAK1aGUhh+WhLUPzvOvD6s/bBnpNn/MojVbXVdZ7VoSJjcXOlVAkqlsyy6JHMx
HXSA129wGgN/VGYKd0k11/5aS/C/vXmiT4fiX0wT7OmSxoctptYQSl85GvLS5+62wR3oKb55Onw5
jZMNso1+89DbiqUYWi6QIuY6gr/UKXiWYTcLkPuJ6oPgszPTt+SNSrZnPLnhf151mw97JYm9wcEB
H85CgDt+NVsHK1ZsPDKy7dQfAzeYfcm66CmjZLrO/tVHqLuwFrkqPIYfeJ5jaZ4WUQMxUZfVZy9e
4UJ93BIRKq3mXR/Vvg7WPMUUyyhe6VZyEvyqPMV6gVKvudWL/A3+7l6fAkUu2/sYeDtUoc9B5bQa
IJ230s4/ztKojqHi2MPR+Mz4I/eIa8rKNFYgdAQEaAaStojpjK2NCKfu+PTYBSbh4kGB9KseOfM6
RI8DJa6vtcEQ4d3UMWAHZRtgePf+i1hM3Q/oIy+HyYEJwPPGBoZSuRlolIOhmzMC5CPcqRNOBK5G
73Uy19U9QnodMDS+GrI2HnRYtq41hMXqBReA5zhr+yZlGL1fqNtmwHK6SsyBzlzT112deBZHMwYJ
wSV8jxEG/WUVqP5r4jbchFeNEDWsJkgO9Q/rUBuZjhob6TUjYI3v3UQH7I9S3iJCRXLMD2PyZ9vR
G2x+4dFzasianYkAxASMuHgSdP8DhCccxGTYZTIyK+chbaJTkhMlYE20y8ktgttG0lKhEAMxuVT9
zTfMIAfO34yNtwu8amYwxjR7xtow35eCKeehB4rDAXJdhPHAhmWCZUZGdGOZF9YqysNuba2rSRTS
v4plgoyc9T2BmZTk+vMAHgzp7WYQPKZ1EosFDVjYOnIiOQ2Ysgab183UN2dOrrFs0uWkX6nGhxGj
eb4EcrKoDsk0KXoQXp83XqEw95M87hcUPZGadBHCC5StegBgQLxzLRfjqxWPXDa3gl86kgtByliu
jqSOP4PtPzGuob/UIH+8ofoKhFrYR7ZW+MdCX/uP3VghkZCBETZr1j/WGuWtby20ehUsdPYf/fsG
VyzpWwc2d0Wm0GKu/t4ddGusCfYWp3dittK56YKRYk/1Fh7gDD5aN/l/HA0XP3cUx++cRjeGJS7y
nqcQa/RGwQVq70m9s/31XO9qof5xz0kTLlcbJ8BhbUwfYP5xTmbwcSngabdUfNSOnMx7FYQ5KPJj
iFv0Y17+GE7AIPIXvBU6ScCthdaUk8KUVOCd/FE8tyrEAN6Sw3Wawy8LdRccaYJrIZnXLNHnUaJq
308XrEm08OeZL7/3iVKVtahuUY87xGZwBKpvjv2jevI2/cHAf0cSXpnmm7kcsOGSFGptiSBkpX2g
9TKM6OL/aUdK0BeR2MUiY6HNyt7Zx2zFbE50zWc7Ho49b8kQP5NgMHiKlwg0dvLv6Qh5ff8QXzpX
kUuLitQAf5Zik7hlBRanxMpn86x7mvbz8+WHUmzU5SGVU4+sLNT6uhvdsQ/VvCQITLaB65Wprnal
dqvSb6ocLfcfo02k3+u+ViHt/LL4QmapCGtudtpsdsoipbtEjkFVYbGdIfesqSvojvFf1xkye5D6
Dkp0LL3Z71ixGosm8P5fJh8L/FVmaeHZbo7/ahDb7eqFig1DPbmvaTqY7orTqi+IjeAVqCB5o0cV
Mv1PeZSxBJcr1egBOm8fCsbD2ZI0zxiq7M95A/6Zs87LW7fs1Uj0/bbSQbrsBD15wzua9QjzqPb1
SqXFSl4McI2wEWoIn1HcV2ISiitD3BVMisq2OSXSWjh3Sm8dWS8IdVTMQRyXG737SRweEot0XoFV
ntA5+sq0+XToA6uzT12ezh8huh49zAWdrOTzW7dZda2E3Zdo8bR9YMcDws4lWdYDZz6mBdysg3eQ
TGH18/Fi2g4F3lOfUWiY2r6XpJLDszrLAJS4GLwVaAvpQ1AvZZvpfBXaIgrpfVjZS0W04L90Vhy/
v434qiFiKNtmG0kmLLKbiF1QDBO1IjRvZttgJpQJeYkKzAm3LsXOua8HgcNRfSf330OhJi8Dgdng
pUisdsmXiSPBE7ca7YGTIYyb5zj6NlkFLb7gpSMNhLrbaxlAPvUtxpVSdw7aJhD9u1MhTesuXK0q
jfNmr7nvAiHbzvjSnaLNgekNoNiyABEHmNlv86Bw/QDOeq88lddv79ynfDSweGPj9ThNJvT6rlmW
PU52Z7EPD4vK5eQPUzTnyQrQEibG+d56jccGU5LQnBLnLMljkfg2TmcC7K4/C0RP1/pZiXqnjU6s
J0RKv3Uomonb+Iq0KJIKnxGAPA++VORfBcUkXE36UHwLg0MpOAsOOWe2OMD51DDKyzeYF0h6Kytf
hBenab/YD5g26ymgQ0ZWdMG0CCVenVY54PZdTBJ2dNNaTEj2ytoLbhX8N8Uh/XkoYrrzpwWAd0U6
5DY8JetdBAq896k1w/lIj3UbWFF3TOxB/ImX5DIGd9lF+kPb6G5iYs+Z6RKueyCurfC/RSJmHrH5
rFguN/S0WOQy2HIwJkvf3xBbceTVaSpmqajd3Ggn3Xzfh0Fl//iSODGgynaDlBmFDgdizytW7tpS
ZETLokF5+1v0cIGOvvf4YbyOMIQIQpmN2Z2/wlHovDbrqjyu3H6df4HICb/oiN10srb7XrwHnqj9
sAjF8zBNp2V+xg5IIXe+u9YduZgZbz/Z7+OggByngf4kMB+lJ0U4f8Ox9QxT+lY1WY/Fpz94Oos2
psClhY4ZDcQh8x92RfLqUYnv4nowPXTGQTSeKCDaog+8/Eug62kJxWq3XG+qMVGjSKG5F1vpg43F
hAgC3xn9MxV6qiyyq+ZgzLdobOX5nSCuarSCxvksqm0+FUwbsSIoj59wu3/mO0eoDT3LvXsu0xt9
KK+5bP4GId6H8RokEUWFBs70iAeFYe7/5899bkhIB2+Lq3xNnpzDxQ/gIj0WetNw2OIH9t45xYqt
dYpLMcG5FAXLpzHGXRnW9heMuW25ygYt2Pk0AmiqHmQ8hVNqTXK3kamjje1p9vuzCTFlKFuSRZU/
NmBP+PL+mzoaPOH+O4JD/9iRGbbo4+o9x4reft3662c9JCZkXThl0RV3jLhn9q19Bnb1Myfzark8
BP6PeUp23xWVOeZXYg6qMFteB6tjErsnGBxpnYfob7JKOOTH4R7r0hM1V4AygGM5m7dN5ehqKlUR
DZaFmVio1lhMnpRreoJRoR2HTHVI/mhOd2eC0JoCq0Bm83O+FsPU+RttNfQaDOzHcS7bAdF/G2P0
D9MqEj+H7JXHm8qOXQXLf5ARlPdGT0p+JHSOHrgLvcdy0zOP3opSt8LBBOinhe7c8biFXXGo+8FF
UK1AWAqeJg2OSImpeqGJO2G/PBpufGNCU7V13DiUxAVSTSYw3Jp9e9PplLzY2r+PE6eC3EkztOHA
Ckbl5eS7rhhaqyIkl5g/iKPnzPsFHemMtQbX36sFPebjPKFyX9mAiGrYrMk9zE9T/4PvPykLn1tv
po9yIm0CP7WcAfz/2ACKUyfy4IYS7PvBWPLXari91Q9+mnlPheVilvvNKTb4ex6VLuQOaN9Qmeg6
DB8AFmMWT2A33I4vSMPLix+LcW1LMuuVpLqq/KuSj8Clamr70f00caU04qFkB+A9+4qCc6MljTMj
S/SfR/hhKKSyxswQdpZtZh0/hRRTIdqR+ogvtVQ4+IqXeGONEZwbRsr6Dmo74k5b9oKIWNj/1Yr6
glWMy4jmhm6/2WjvecvmS0NlGLQDFIIl3UIgKxns5JeICqXLcOlBbLQYbey8vVhTTvE0R7cEw4CG
fkq7U7+O1zn/3I6GFQZqec7qXHkbeMYeKcdDdO/IGMiR8rbi6AgdiBSiut+Wmd9e6rN3g/xVtU48
Kny9Sl1lz3pSuIu52qLd3yIYfRjWdBzD9y+ArH+NJPA6puVV51LRK4YfIVcA7W87hTK3UhVO6PCv
TqaywcCHitPiWJDma2vDLeTSS6OxM4grWsgZzx+0pI1dO9fBkZjm6GKtOR0n2YJJiFwjWekHoqiU
9Kf1c2Ja1rwBypa69wsOG1noF9rDqMu9uQjfnjdKH9pQpNVnlftv2BlIp35SQtoafVtd/fBpOSJL
e1aYj7Ozk6vkViHDoi5e/SbONj80lN1E4KjZsNJ9DdHx0neGnwvjTUythjsX0hD3Iyf+UN2J5U+O
KnakwadzO+jPyRilOzeffI0zvaY1jQwhqV390i5R2dpYU9VXh44OHHS9HoGUky7O8MI1R9n8gTHx
tuXL3S+Og7SfvBr4s4tEG/OxTV1a0E5BUefrR0H8WPVP9DBFe5lvAA73hrSu/UcN0C4XnSiVBpWo
/Q1Qk1fNQDlFGNE+ERWvENQLGKEeTFyR90Czo00L9e1nFxjXwyjbAL/GxbiWK3csrm7edX99EfDd
nJ1Qn7/AKRGjW//URJrVqcuhNUCjjCrntlMUl1mX2ZjhhhWsmNmgm5c5RiWAYHLTRO97C7/hXdTc
Ss5E+/VyjI/iTJYRbnplHTmH7sEVIxrxPPLj5NqxnNnIIcZt66pGBZj7Vw+CkLZ+k6UBHXd74axZ
6tLc8L5VZOXcqks05mOKOhIKUcdyLmsUA0hABME/oS8ZH8pLu4hu3fQrT7C1tP9MVsclL+v1eT5l
Sjo1+9nwQQVbnA0i9pN3WzhGO5Mg1WU8Kn28RvIiq9mOnLO5DU3la8x4CeejTUE4s5Dj/e9c3KLL
iK9igsbFY630SjwzrSUnWJ8gTpcBTFnplDUm3mkt1CVFm56lcrB4QtCFofSQPnqGz5ic9OBUjNXx
C6zXHy71EIZQHcUCr46769WUZen6oDy0PqdxzX+dO+QttjQ/qSxV9EvJWfhHqcAB5uNPmComvblp
xTazlPgAAUTEBX8TevOpvlKKj20/OZQC1IL6Q56/pVRDUO5u96F5xslpwVGCNsgeQ/0In28F7Tny
BNzhb3yNNWhNOrbYfW2YcPN5qG38pooN/F3Fy7cWjd3ugppBtI1kJkI9VyNeQBXl8DXxpo2eD3i3
PzHAjha8aH854LJ0B905I2Jnb9JESgkSPraC2Ouv2Co0aaVOscfwzUg/r1nCvQlW7x9TBpIS3nvw
UAvqPS1lLy56xX24feLe29lEAC2TtAE1KK2ThlNKV5BfEqyYxtoQAq/pAurlXpq+71cQcJlyMJM4
GE+foYZcc++/I6bjM7mRyjjfV8mYyMdumvUYgf7IZ4mVZawr+XakBG5G1FyRbKBn0BsUyWc5V90b
6cj874VYc5fo0iMgLxLM/9CE112qeYkNTaRGcj94RokrE0CY2aCp61VUsr951YMJdfIMfdKvaFEh
drOFULmChXNh72PrVVgxpih3R1kKO4qbQWIzIXBeLgs0hg84MqE91Pkz1uWCEg6sQPwLVCwFA3oF
8fHtHWBqGo88nCZTeo1RRqoyOPePbaFxojITw8ec+jrY8p/CuXp/bylYBZ47cj61FjFi51fOo/ap
gVa7K8LwGXPRCFUSvDkX+z/4a0dx/fvX77uKg26Y/ZzoN9g19H+/yMOzdE0vNwfhOQnSov13uAFZ
aZzO3n3ZmGvq4cioK+a6OhfTLg0acbmN+8krznUiVNAcc7ErKTHC1DQPvHiwWBXS8yMZ3vJvQypf
/ooyLbWTHBObz9tkMKRlR/CzRPnr3eKj8MeGdEl1PziqeOGzFM9vi5oYvxEcsqQ9be15AmPeZluJ
stYEXsOjgUos6iSNGL+NAGVsF5nKMHNNnQaHXwK5arbpbNEZMWy10P8WMohc7rCVplwqX6hFXuD7
/EJPm3Ys80Uw0gntAFj1vn0Qcc2+A7BNFNAMuCe9f0MnNd7qnWg9rf1o+FlN92NyEZy0Eq1YhCrZ
eCaTeYuWrBL5y8WWlrCJ+RRLfxT8BYADtK/EEX//YCCpfrCqHmxKT6EwK68UluhxFDEdrW3Okld7
Flrxv3J7nNX1JfVPCwEvndFxuAxQnOTFYsznnXWTM/84wL0vS5r6C3Z1DkLzF6cUxCmvj2p1M+1x
YHDeWIp0BtPXbr+XAEtbnD9d3xq2ZpluGfSJVk7z5CWccJlmbFprI7UTEm54/AjnMppHmFGResuI
mzq37jSCQt81nUdHSgvWBj2avCusDWgThsLpWD1hDoMFR02OPVdP4p3lvYN5+Voq6QF1VgfPoutF
rNOA8r7Se9PfxKcSA/svg2IRDtKkmOXa7fJ1zEdGZPTEpJRpIINWlPq419RHOKqw7Pjt0vyE6/ev
mP3MmQ8is5Y7yt3EAfWphGCx5j7TkaMZ32dP/11zrgBnKQrPyGDuSlS7rf7VbTEr/dvZbLNZCkWw
obMHI4GTxZs10Q3hIWi9llq9HHSqq97oJPKMZBw4qmzuzWkTcF9t7QNtF7Z+zZni4uA0a3TmdMrF
nfLmshJw5fUGcyUMD6ohuNj8KwFlcLh66FuyXL/qmb4/gqHy0HBXGzg61XkP/gTfOaUy176KNbdK
XHnztzjsTBcAg18S7w78w2WFZdMDADt8PMsyIoZUjZssv7VRhA2UtsBSTQLWjXe0npMHRP/ZBigY
TicojCUNmRO3CIVTZZ8IrNDPKpwcJSODcAU/lWxTkxlGt+98WriDEpGiPnE3EhMXPw9SdtN9ne+v
LYLg3S5TG2+CABX3XkT1bDc0Eo8sUBV4Nt6clCsUfD9F/BhX7OXhRWaaWWCXyR3wQ/92TwLXb15c
GFvK+h1sx1eo2y3eWTmRMnyciF3tK7tsB/cwLMrj2t9UGnj0v1fCDi24Fv8d41mORJiR6pJNUOZV
0G6L+/w3SaIbrPKbSSGFTYGuxLJHnR1pLp3raQ9tjHMcv+xig7R3epvNsLa7HqKnomAaqOad9PYA
f+zkFE/+XB0C0VDgc8FQtrmFjfsdKBLf7hDA2Hk2eoS1eHp5auausVYhhvr9eD1BheGuJJVDfuze
kfVFpVhb9YwGHyct7B5u4skvewlKjVwijAYQ8dolnnh+if947rea6rOWtVwB1cbJeoRApkwi808P
zkaFFlyAKPjlvChFiRvjzuj1zPfu9h5uVbP0nqtvdQqXiMVYdLbul5QbWbQSyBSaD1hRC1e9Y/7+
CzWfjb0oZomy5Yp+bxiieKSse593ZGbSo5NgSg69HZOFokYCbQyRhHAkwSQlZeZmL0Jhv4boNuEh
LYnq7fUVn0LjksLn97NNzISuhZ9qbje6gWAwLLRq0yrnyYmQZKQPJjTdX0bcH9kmp9FouXGiQ50r
JpjBGQZis6zAagXubM1RBvfN1d0PccYIMJ3ePF7HD2Li4ShVpIQGIUb7kbZHDE3oGXHSrUKV55lG
N4gnJYYqx0PVm6+rfYZZlMfXb07NGQoEcCYhulTq6jC8TpHlTkhZ9RfcTTo6EC8Z/t5PyG/4SWXs
XUAJThERSkmtAIWodUmxMw32vq+uJY/IRR+BKW4yCoVvAiSNyABsdsKTRnX3JYzokx/h4HyVYMzI
9QvQXJolzKm3G6ZDzHdyA44lIAvJ9aslVIruOTJs+W0aHx7rAXP6B6K6tnpQEIBNoVyM9yjLyQno
8KrfzjAK1OIUlidGUYZOzp3C7m6PzCOmq4SkMarOZOH91qb6DTQnZYgHN5qbX7b/dFijF4fnDD3a
B1SssKVflBZ7W2EPQS827vAO8NHjHRK4DV29KI+z3+WEy7LRiu8TFVAHJUcXqR9tHNxkaKaiaVCR
LsBR4ocYKdwbBh6zRJOoGF7zvtrJeex3WlLlBK3yz/uCFLZ8UyDgGag88PEmYgidjnwbRAm1/EbY
X0Ao3yp2yPlKwDOdrt8ONepGy2fjQFdzlokfah8KKlPpMw2CYmrpjYqkrfa5IAk++j/LBzAYDG3Y
Rm8qLJgXjARWZ233oUZQhlpQywwsUYu0c07X/cJur9ma1GGQvDhrziYmG6PjkzxDhRQUAUQoe4Nm
okZX3ZGZyV4T/M7AKgb+7uhC/3okvzV+DVOZ6KSJCPtEW1Wfj6wGVTgIcMVsUFzlJydrYfdMYl+F
KD4NCl25g2xTxjxjlQRKawTCskREKDXj6wjOZWyrEuTruY2cWClmKD/CfFf8VmBdaH5QkUvV5zxZ
VemALZWRlvRGeDz6aad5DKHiyb4GrHX4HsUskwTPjhgBRWECJJr3Aj9gkevOKVXYFsPYsImuuuyd
0XVHmMDdxCSV/eCyHxvjXwkiu5U2mTdjb/Nw7XgLCXt8t9M7QQ1F5h23u2CKv3zzCdjUlaJKAK/Q
K2InsEnjx5hM/sQbWTDeXHtP9/6J2WfSKxak4LfPUHCbZHMhLsC9XUKgjo6kf9P3BVdXk3tEvOZK
REKRspC4sWftc2SsjWuioS95R2Ug3Zw92jQ9Iu7m1chBmLxoavEnSiPenwul8ZM9RX2LO9rPk3ou
fGYqwKc/s7IxROY+Eey4g3pNLFQZjYq8/rxq+Af8ExaqkCdtwY8arwG/VN0E8FftVuEcUzS9XGjn
ih3CZvNqxL8h7jSdLOcYxhpe6FTRKe8I0HRKanaC1bvlzRthxibI7DvVkcD3ShiBPUHyiR8zHqqz
RkPlTzgic+1Ki/A2cihLmWMLoT0L5+Xp/JFc6ns8HuG+Byb/7x6svcdq5yVcd+ibi6sKj4BEW9Uu
9/26SlwnlEcneZH94PlujKponSrWxZNtYWpfUv1oiDdbnQfMZeUfN9mP0u0NuW3Naa7aTAS/8rDU
utAsgvigujBUDtOrbfSJfPYPBwTJjfoEhimbF/2pHoRZEwNtMUkhZPBp7WPMyUcWy4GCyNDgrE1H
88qhwvUFycVEWmuZKL17zJTVdO3nFjvzKXcdYZxSAAdd/R6oMQxR3jbGBIw+/5OzEEG6VsIrnoH5
6/oIaQxcW9egZTBxABpHcVjgkMBAEpXfKjSJTJdW1UvC6fpltW9iZuvTcy83PeQjdFOrpUIRfj+6
OjvmD8vylv3rCoz6oGMmey5gDk0PsCkwGDFVG4FfZDvgEJSQk5AN6p3qxDpm/X/aJ3e/WhbEie1e
a6q1N7ftQhilBEWoXEYeQGn+7uuR6rqH/PILNW2BCw8xmqCxLmfE8f+rWX4WKetTJd6dRiFFtpN/
vLo7zukY7nEQH4MhQ3i+rgeYSasPdl75ucu9pE6f0MnLSIRRqSOaBoqGZDgkJyhcKrBcB9PI8Cm3
KjsuGBx6BljAycVq1ZPZ9smYQGckFYWHFuUeItSdvAWkAPvoUvYKP1pVRrI7cWHnulLOtbifdjn7
i4BPj4ClHr4rHSWlEiRNPenK7iAe2GUM/Hr8dCSs2TkaJHUXlYLQKIT75j1vwtusJZcpN6NOm5I3
ob/UqJWUAWGXka/kAVt7zGup3+mZivaXkknHWt4GWto+f8kTfFDE9it9oKBXAwI1s+IdPbEvVeCB
v8zbc94AqI1E99ymDc3sxWImy9XvrI8ICXL2+nbUwokQ2tt8/KzO2yPRIjfNooAhnVN3acAGOo2c
qVuNwwxr+jxGBQrdgEn18HN3Z6oPq/++I9wEW7MWXEVraIYRmtgtf49GkPx7nPzH0FCh7TKLxlPP
p7nz/eQBP5rClqFy5vFaJ3L/LWq4xzXE/wiqE0zWiKERqwtw2vF9//sNZJaYaK2vt8sDNOV7kbQt
vJqOQCh5LXoXKksZVzv/WInS91KDuWJ4HLFuneAVOPa4z/CbAUSyahoEFms2AVhYDYoMKYqAm0BN
Dc6TvBC0ukwiq7+bDqdErxOrtZ2bgI6YOLzVnysC/gFemjgnYWSJzX9wQiBzFhsIYRaxt7cLF0Vf
WtoFLmcEcF4Lgg/UN9/kiXjc1fOZcuG9iP3FATvZ4zFLbxJ+gQ5+6GRlFWTYwEdx395SgcRGjQXg
2y731PIxz+azh8HBDD1ROaO+3QvCjs/LvvULa4ZgqGH6tfUxJYi1upZsdvUD3act6e521CIqY42D
KW1m3H4gY5KIhwKT3Gl+c1CpYR/NfvmJ1uPgsGeUTYAVjiGm0aX2nXfyLya4e4lP89zvaFmvaubb
WLpRpYiuxB92m9Fdosyk5W5pspiDiQBS7t0B548t9DmINsYVYKg1+90kpTrHwpvLazPCQm97myGO
QaPNVVnMdFX7Hjes/madOeNu5x6iIcGpXkBPHqZhV9GJNJs1vhZG9rZSSLsv1zEtJAhed/9eQ8kP
BWfBf7xVECKSo7NJMqj5U2Lnggc2MZHDIu7K7KJa4VO5nhzpyu3Gsy0JK3khdhaJHO24psvwVkMw
W6KLp71b+UdbN588NxNIzO2eHzg9V3oTITGp+1dsl+PkuQZcRqaMQYgSoq7ONsQc5l86qARQ2CwF
ajUQOMVYydE9EDMAlLyLHgfAHn9spcwfDFoY1ZnCvy6DgCg44w+Sf+dmsJ1NMMRW0cKWeKhvu5Rl
/P7fMaWuOBra8GfW4zlpUIHa1V4SSAUqcvIOFJOXgWZeaEfhx5w7OfR+ctYVn1fWR8z+qmX1fT0k
D2ADSkpHWQvebOMjbZf2P+uXagi1NIlu8Ihe6LhMgp3WF5N4lQhFE3uJec9MfHm45yrLTPg/2ial
qzVcK2ECSO1HIWuGfaxTiaNWIHrLIo6qfSqD1DURaWeo5OMhfUec28dVTnagNJ0pADlx7ieu1DDu
GTQbewxdZ+KjjsYVyCIsE2zm3PliVlSQCpbi4xVtAQCRtvm4M9v/FRVNPiJ7F8C5rD2Te/vwBcz1
nJUmtI9PZaMHeAwIgLBmg2VT2tSGcAI4Kz3gQn+nBt3rmCEuB/qq6W/Z8YuDzFMS6iHy0ltYCM2M
BjhY6uu044n0QEadl2Hcbw4S5euIKZk/9Hz8frC6GyNRRdE1bO4cMKsV3g6aP9zf7P/aa6LCpc+L
tmzxgrT0B9pFEaD6F4cfRUdbT1TxPaGkrsxOSVwdHnzRMhj04gd60UG14D5omc3wkTTf7ipbW3uO
UV7WisVnAKlacoqzXSUIjVAGtUEhhHwKBHe/ScKLwKkPS6Cfpp1e0pszFCRYCbdbquA9lDxJRdi8
1hON5E+4GccXCtUaXN1rAW3zLL5W7v90tAAUhf2g53eJccFZ1IxHUglN3qvpGSivSWRdBnBhrkk6
ydJIMbE+JWozA0LF6t222DxVMt4Rs/9PkjPt7szbY7MrbH4W189asuRNb+xFxmJm6rMOmGhvAPuA
AwBVJnyDDNPwlSZ1Gt/hamp8c83qdBp8AU/OYfF1oTdiT4fku3rpa53D2Ayyz2j2G6LHtOQOqdpO
UHNWi73cYfDmXMNnEquzhFLoPqcp/ZQEmKkpohZ6BXg3Bw/jyU9YPw04ubGS+aOmIbN5qfEO6k6j
QkeRRX3tkWCykWG6PDoNdSR5NSg+Rp/CTZAN+jia/gpb9g8o5jrfIvQgHM9bZtXYKLdnohclmubw
bwVGKuuFhWz15eL8XVBFG/g42QSC1iatvObDrb5aWULa4zp8LwhPNLhUhn71e5b4FMLUASGXv6F1
Ey6SqdClwdyaI3g8ztHZopMs72OaG/qMmpsH4oGciaM39b+u3H4ratX5vMklOw7TpXCl5yKew4ga
B3Tls9FWkWK3BY9knxp6VyCa0ut3zsLIDVk18SztFJISF7pDmxadgCG03nB5x/X23F0h+y2g+IOM
OKdn8jue+hKmAqmEw3xPte0jiumAvoh9xnyygaZ//4uGXGs3UXPyGY4abt5++dgWTPXKyj7T9LkQ
iF3TuJqVv9j3h4XoJZK4EfAQciUBik/v3q9sw9raP40jyb1RVY0UO1dVLN81BBCJkk5Ki2qDX9vJ
UDxMghfPm6fV3Qup+4i/SRZvH7sBAvUfUxGR0XzkLLw2fjlzsk3p7JuyH6zWTlrF1VRrVjKzRVnl
YxNc9Et7qD8N9+nCZh4H0O6WN239SYhkl79CUBGV3JRaS6UyeRtV0/JsxoRWBORVIEnOzafdMpZ7
zrhMKWkaEmZGVAg5aInASEh1fYYGlmcU00oSFqxyIkH6xO5DRp6P3PViz4bwqtzodhXBQqv20old
PaB1FVlx5mRI8J7FJ/+JzNMiOu1lbbEr5k//ADzE486vUipDbty7dx9UNMqA6cVxh2W9G14nNcFZ
rNemmyv/ErWdVFsmUVJpWlFS3Kb3sqTgGA1skzmu1MN5ELrACwBsrtWxB1Y6LT2VIKS8+LaIEv52
Dox0f2A6F5LtVBGD2EbCB4n2mSQ5h/IbkA7gd8rf1v1WbThrTpZpmF8PTs/cRjKdkUHGen0/YjNV
ripw3E8bWB1dAm0vm54f0cglZSZJu5UJkRK0yaOe4OXd1vBpRULXEhpdcymzuoaHOoGnbVc+eO7y
RBC7ZIBeGatRYdapK2eIAFSdvGBPOdXG2ANgVVCT/W2S6ZBtbeTuxx5gZir/m9ubU13ahbuKRSMG
j+Q1rsFTHyXV3uX8P/Zd7sEvc0dSG09Hdgynf7XfNj4W4SG642nsJuHL0za+Zp3hL4cYPOb14++X
WTqYwuqxAbg16lItMXM95sy7TlC0hObfwNiTaYRFkdCNvWA+oGsAIuoWxcnSfB4lyDRuvkKyTi3P
J1vSmM/jKqr70ojMncrHK7NVejg86fQaswkY/mFM4aMf1xDUznUU+DOwUt/LWZ5gGF5s1mzhVCWw
D1O9msdbkiZyYEhK2A08x0kOFfCWJABnUgofZpOieayeZC7ZgFT2FFFOJCwmIoC4U95RHy8XG850
vqZJyYByJz30+aFq4DPM3SMwXhLBJutqlhBCpgE03EZmVw/bSaqor1gjS1C7F/NCpjdjUV668owi
VD2Aed8U4BXtq0BflVUM68NiWg/2Lb7B3yOoEgpeiF9D9HeXtQsv87h8eQ0HGAg2AUsAjpRaLa4I
dvYnJ0dbJtwqoeaiJl2vK9aRzJ5U/Cz8a5Wy/6DkG8140UxV5IQoUYozuxFxoxmil53Uw/oCfxTE
Ix/jtJ7GGZVGTXMeElOe/sxgPVRKO1XAJIgehqbgJ4zTD0ryQZ2IOJom2rbB65t6il5fEs5DfLl4
FVVw4OKOctLZHI3luSU7NZu51wyfaDDmyk60E8kbklBj5ZAgL/76ApmloIvlgKSCGU68wnPvt2Mt
CGT9BJQiKV1zQZFPpidAnSQhNdDW9R+eWJ6qspRqy07h7+FBRyRuxNxUEoXwh9vmjTLiOJa1j1z/
rnfQFO5RpV3I5utc3Xp+LNgj2t+3sKOknU38bITsaLmlN5gbYv9zHfPH953K3WfTRk+Y6Gyze5sk
YVS43vZrAi+tOP3ragB/NJPuzKwC9t9Mj3WxmAumGLLMEbrwE/px2Iyrt6p53G5ZSB3U99bAWdbU
CMXaH+vh7m3J4+I51Q9VIzTCEI6Y0elTkoIsrSEGydee/tUxOiKB6TWkXcQGBoTDbzCZW4opwK7J
Gn//eyQVbQQFvUMg9Z/PxzhtY4YdFYE1Q9r24csRfjYLA4dWsjLaomgjUu9nKwHAQWZMcjFyFYxK
0Yw62hCQeAOU9yzse110r4wZK/f9bog0VzLWwe/1/B3M/2dLohXIK/rp5tkNtyoGra0tOsFEujYi
CE31OaSG80BDMKZBrTq7lk1kjOvZpMLSA9U/zSRgPFhQd0JB7uJcp0I7wiQWcjQKwCxJRNIIy+ix
Mba+gvK4+r3nUrcAjAClvxiZJRta2sE8dqgk1GxA4jHr95JP3JJMSJpwRtUl50J8Ty9AU/zlLBqx
MgQkmCkoiZMpmd5uX26sUD98QRUG22fxeL5V5/S8KRNyPfG9gKVk3dn4QJEbe/zsfasNnMyEbRL9
vMzwPhA5TH7VYa6Wb5GyvS+LLBEmYzIsmo6Ee5ArRVXY1p3mQhYkIrYsSzledfQdbhiEWcko8LpS
FEuN1IQBCzPO0fIMpqBuQIS3WAWIwWx/oz1scYJ5lu5/gyQGL1DvenUlrwNDbSFPRb62uEmvBi54
ki6Mb8pnRA9eE4yfTOHqNiQ9gwijwNtTGO6eAYSkavf8dFvDO4Pt1/M/HlUgZayfKGfj3ZlvTE3l
4/7NIrgdlO6HNepNqa0pX3em6JsAc8Thxv6qSBnfu7kXmY0f1Aziqytz9sE4LeJomTfHykUt910K
Snp6x4274OLEPTK2270hibu7rMYpCCLDe7cj70aO+2hRlzCLM5FxAvdP+R1D00j8FhNroAZBf0Y+
Jq7FdtJb50mHmn9PqgU8GdCUL3ch+AwgULQTKqUiMyfvtCLDwD4q4zSwrf7R9yxAOL2tw/rZ9Er7
ZB9aeetXS748x768fPnfnMmvmo8goPgRj9slHVBtt41SG2mgE3LKOfh4Jk3XnVZxlYvRCulBWYm4
KEhcpcrMIzxxGYiBljl/Ng7D/79uewch5DMcflHGeoUhxndIxxxr0bEken7o2XHjd02KQoHJQ/B9
ps3/7NIzhwYu+5S1paL0zmI061bbbnye1DxuOdLckl6H2AntljLJct0AQfMHbnC8Hcfk9vYDZKxk
C8Ms15SbZmczHUHzKIfyaesGGsccMv/1Mie0ZZFGA9apdHiW8K1xVZ/VXsPFk9FH6zVbF70b9FDl
LiDYKa3KrKCm4R25c6at9NjoKPR7VOrtYBKD5rAGGOCbTYjpypOktDXxHG8/QO+4ZfD0ZL7hPsL1
oWlrIz1GebymriNS0QSRbZmHldbJqqaxfq8fSTqOS0eBeYzYrYvv4eOT2Z2ytnKGBEMKep3mUcqa
rBn5hVyMy5wdNe/+PmbgEmsSnTL+q9BSj4n3Q36jQBj+/BcnL7a2FCxEl/It8VmZZTiQ/HEu4V2y
aoHUOtAhlm5ZBhR++FSFvuocE8CQn+/TQdIR5pq8nZiPLRIV9dTuRzkR5JVIz5Gqqx+qWXaglGjN
ii7L6M/HbETsgCDkf5IDDBNVhxyCHrYRQJkY7jVSSFOfS/HW7OX5SgsETNC4+E4cpHsjjo3wXtOE
4ICRg/HCSWQRFAnp5BqNRppjej+4j8zDKIrJQw+uT7kOHkfd1p8aCJZG0UDNLcnoPBLxuw1I5wo3
fElygDbk7eop4ztd9OM11rYJvIJRhunbe41XAFOBZYhGwYKegCPpMBP3a4Z3odvOdWy3saqSZhck
ICAMmQ8JdO/FRD1nYOSLrLpkcjXm0roeKpzFY0wf6Zt745+rMNYItixDCHAPzGaSo3P9EVNFs+zJ
2TfFvzLUBAdN4h0jvMxnmmwrRJosm4MEZB/xpFySGkfjZQ1Nv8QnOYH7nKL7vVMVxEQmP+Kaf8k1
ZaTsHU9yv5RWqJAWyT5KCTPEKv/TBzoQNYjksC2Btcw9qVAfO/3KQWH+4wuiS8Ob3Ufjgl51lcqc
yyqvS9dVVIMnQuteqaTbTwr91+d7YTNBj381J9SWMYLory9sHy+fN+iqHe7aYro4KLWk2lF5f5eY
99morCi9h7j8c71KQAQo+zwgS8HH58LXj41YfQarFZK+7Oksn53oJvplfqCp4pDnI4GaPmtYvN6C
12gHCwdpH09o8mIGLAlMGK3osoKV1uFWyi0fIiNrsAokwKq0Ly6ebW5QGAJDPQxG2DXDtYXc5xyx
JsiEm74rZt1ju4IrcZkkB1491Yz0qS+MgASeCBvR7p8k5swCHDguS1cQpldzupXTl+Px9Yl3fNRL
L/xs3cvL5dfLTuU07PxsZ8hYTBW7tFiKdhj0Fx+/HIobpjy/g43rZdr2AV2/uQqbozU0lX5Ey4Cx
coFZNmcxp7ng8qDpYnAeOlmf4tSh/o9NUayq1XxLbzXyAd9KJYJ4i2BZTDkdbW6NyY7aF9N/zMEs
wECh0h8UDMmqrIAZ8wWmSl7Kcb44CLSB5d7Rg3ay7EkQtnt/0TL1wKHPRVPh8imz2O5K2YlfSY2s
U9nH6tDkNv3EY4YQXLk3g9p1pH9Ja02Ie1ukHg6hH9zm4MIGWvxpIO9SgpBbPcBLlUNl6FWrWrNM
PkWTv8X8FmJ9GryI+8D2HaTAPqiF6IH5COJucGulZoMUbmiMSU1kDaUAYq6luQ6JAlOkWwli4tHB
zmx1btvb1vqLVz+BuxDMfcVpRiix6K1kAfTYyGu3sTf/O8m8JH5nLRd5cDZiGCJ1AO+b30wkutwK
/y9Q0mj62IUKIeXjQExSruHVC3LQtGmgdt5MlcMoOhcHDsrmRNfUmmPh+V0tPTuXu8kFHQwnqK4w
0GRtlLLnwJs5rg8SEKzH5Y2Z7ERG02fuJsiNHbwx3Ca0uYv7wWqBHpJFfkNuMX2FmP1+j2jHG4sE
qRy1tX7w/Z81rfxlP9H6jP9gicePd5jT9SgjVNN7dGq1F/0RSTC9ZhY9NXtDkC3wID1B9IM1dOYu
f3hp1DHhjcsUjnHpYJR4lWys2lC4mxjaEWA7a/+U1uyh+7H/Rhgsbih49EEZ/5aeN3gqlMwbesNM
tX4axED1+XxSgQy2cSIaihKhKqlBfIq0P3ABCyAslbuoDSxRf4WZ+vYgekpCzTevz+DhwXoaSc7h
4OuRZYKcK4bwhzBv677a7lac5rZ7P9p8YxNIksfg2s5oUbdrzCVySF5+20X2e91biB/iS7zBpeHU
1JHWoZFVt9OiPFx//N6pS9K60LS4O/WE9eEVaswcAfy8PV58/5DNjSKDvWBwI+CJPK1wSo/2BwhO
jg8RyHspgTDSBKy3QOFefTmhq94VADHzY0j3+a0uilTgsNeSuz+0AF2K/rsdhl6TIGWh6/KHdS8I
BZqVxUsFKok5IwVTjVOXPtm3aIONLOEXcxSG6nllS0UVv0ZL+Folo4mjiVuDwdnxDIhEHby2konF
oFXaX8BqrRXSzyknA5oWP3wT1DUnDTVnvruLS8QZM6UJnV1FYT7KzXo4FsB9cPtwa9hETGldY430
fkHO4h/5w9Fz0XrTWgIVzKePyD1DnUKf8+8hBjnTV0QTX+XaL9UnNIgVVtDWCNSsOHvMPceeRv+f
PH6SHWQTWPNTJP7MoPQUf3EPffYwAwopXLPdLaxzX0/xN8sSWatyBSqQv+qWqhhKj0LYTP5G2yhV
Zo1cE4MF52fdSuig7uvZvpZYnk/I09EJAFe49mwAcXfNML9Ch9lS8kuLAGwOM+ktN94e80xVQHSx
38mvsjXOjk1Y84hGKztWaFVWYItRZSkqGH7HurOPNlyRQr5QkYTgNcj8aL/EkqPSHS+OPBx03e3X
MNKwESEt+zwGBOjUk7+Lj3G5+Ni79B4Zxz6Dz8EGgexj2uGTLIquX5YAz1uubUwFX/RGsff/qbAf
hkaCCJXmK7OMmR7SPRgOjZ166U8kXka2B2HdtaJhFuyz8UANRnOXzcwGxCruCf1aRLDdlet5rXhB
cKBkFzFUGUluJszTWg0Z5mmBTekxj+intVC0F+HXGc5yx0KARPR5Lo6gNDxnkdB1u3HznoLXaFnN
HGXpvM8ZDBQRJuyW3DLzzya5qQdIO1yeCq2WK1euUTIrcNcWwQifk2//xl9zFQ9JHnFcB6C0Lkmg
lzZc+FuIwts4HbmQoSSG6K5gmllix6GKOmjq7+e62Q5L9KaZ6Ii+qpHFdyy8HbrBO9rFSTyx/Fod
Okxgx+p9XSVPNyEAJWPpCzFhYeFOzCqI+H0Stg64NOFGi5cQsgB99ow5X4WXhIp90260h/Sj+EiF
maKD2ZnDJHBFzC264HAgcYZbO15S4whhosfQ9bt5qxfwiGP1Gh7lguK3wJerrHK1FVhxmAtNMDEJ
x87oz7xV5+nLv5/CqYKUOAGLtU8d58wiZII3r01NnB0W8mAFCmKnSMp23xsRY8qCsk1YeynJAc9V
Kpi33X6SRpV04jlp5xAzMXJCkn4CAReTliPWtLU4KOWSTN1MjLgDLbuE9yvFV0XqeYmfBtKG2j+n
8zbjeFKGKuFqXUsPV66LGMQHPYGc/S3HoeLVYPo6N6FQJP34PiLKEel3Cm4br2oyI6lh6wwraThY
kejsVuldjQcmGl/SAKMmaZ0uL4bh7weE/jiDdqisS5ieWPVSTpkPkps2TGvj3P+q1el/M+CeKQzC
z9WWIhGL0gkJtToegBtPZD50rIAWn+D1kV9iolWJHCicMIDENLjFlugaX3o/2XVwMH4gLUxMdmWV
X5Oj24FnFZgftAQYuf5/+WuizcuLZiAWT9M8kb+muidBPPF+doYUpkJ4AkYB8I8YGw/nLc9JiLGz
R/vkvFy8XFr0CUy+5BwxzHHeie5Q3XVBzwyEmINe7eXiIfLMDShfP6QNSx03KI/iJ+SSYoajD8IH
l+FunR0dSOZX9BResD6oArbzIjpqGSvdVJLHSh3lQ7L8ve2/z+nzRF6B/h7r2edL/QBisi2eB/3v
3vZTeqM9Uc/YYdy2xNOisiBtEiITaaQxAF00u7619Q8Go1U9I2x8SnjaY9UGotNtUlLHq494gOAi
OU+C9d/eSJ7RCsRPEQJSkyr13AY893q05Hs34+S7cE2hEACmWOpB5stbYVHcaxC7U4k/zj0FaPv3
960pMF5IvG1MGa1dqvXQwleVr2XPJlrjd+UF5xAaRB7YCxvRarwpvaWWIgD/z5rg5dbosT4BmON0
V5ho6/MSSLYNm4p5/aUSkfkXLeQJ4HGPIILGxB7rPrfBDTThSwAMC0NX45zVrU7CZMJn6O2vovr+
oHo+enqjbbYIoeSu+rGHSrcpKWvexZWbVU1rMrNCjCN8l0dYeGxcan1BEh0aCE/FeLnGtDz+BYoj
KiMUSvU+9E9n8G9f7DiGgmMJrrADVF4w5P0kd2MVgk+v/ybuV3utS7kz6t1r6JR3IQ8nCOn8rZpW
7Ecta2KdfnH0UAl4wZpr3XOHLnA+TD33AkFyGa9zvQHAABWmwqRr9Kk1mtiz/kepSi5MSbxRlbRx
5nrMjir8js22YsKFvB+5Uz/XmqLlMptbjCKriuWsWfBnL1SQle+SGdi3VKy36BADQkltlivpva6A
WSn9r/aNAmBAmMiDv/jtBuGe3osl8Cmb+wHJ1BTgUVazEBzLLHl1NbO/Mx3zKlJaRod0VDWe6Idr
JL1vFxAp3OhEmfVec76OltRcXix4Jn5If0a1t5Ndw5mQsz94e4yEcRLzc37VdmLBTzIsVJKnAJwM
GZEg8eE/hwmyHGKyDuJxunseq59OFf6IF+YAtXfCFVGFqftKzK+4GbVIFrhrtp8HQQGITJ1AEWLF
gcr/+twLFora9XGaSkVT92OMhiRnLmwePhgEcQ6SLjbX6Hd6zwe8p+O64kTz1onbTFUcQb0WkYZl
7tvq+w07lFntuP1FRJOXTwUfag8igaIr2yRvcPrGhq7TnTECrfN29bm7GDiLM+/LSVPW48Ptvzn7
dLBkHwDfUCdkIW3IbD/WmsanHrT4LzmA51jaEYcyrNp5ZLpk3pk0KmpYZNgswBL4qHyHLOrE5Ebr
y3Yw8YavFvZ5qKmBZ+BkNyAJxDzCQR0VnQDmXQXEk/fDlE+nC7xujw0EryDVCOTwUKUr8mCqisEK
u1Ec/wcQL2XaO/5VljACxwb6ZmHgKIIfYbLzr3DdE3wpalV9BEDys3WnBdbLR7q3m/shWDRuVr5q
wzUJNcfAPex4HCvNEIhS4m64k5kqWRE1SAbxxg611Wck6Fk/Qh+zBowRLIj4IBDr2642U3FrhPc/
jfth6dB7xvJUV5EMb2623nJPYmCXnSnxizO+L5mo/mDqKHaKMrBf5na9PVnxFktZRCMuYcd7kRW3
+/JHjLbwu+2srdh22o3TEl3l3+5xwnfu1TDmD/KWnaob6tZoz4a0I4rWOwCA/NnFFOH+bL0P9q8a
I9TFknnu+S+p8b0c+YwWKLY3EDswA3Z1CMDaLCJ2HszWwWcBasleDEfbK08yUSsx/j9cNqinaeAJ
Ea+310tBhCt+1250K1QGbwov17b2T+l/bGls5vST16dFBo8oyhfPdC89oRE6VJbYT9a0uS73HOQ6
YhwUKlkwUgjAxYR5bM0xh7WLvkXSLN2hZ6gGsyX+8aiaOwxJvKjFvQL3/NgAcgxW8i5N8GRRhFQk
tP5R6YmYgtQEP9Ld7gUcKE8ouJ1wFwLQSc+OafJt/aOsyZH20hnL32fco3H6jjNla03gtWUGxVZl
sVr7+Ve4THdZN1HW38Kqp2eVhzNy5guT4b3xN9+O1lRIpjyRvfxFme9j1u0zP7pIUNw1395v899s
p7KsKYinoYEyTaIah9VgN1IyY5FikzgWOGuIb1DOvMmO0vCx765YyzNoKdMkjLk9A8nl4X1zrmU3
YkdjITcRY2OTKrc1cudtIYWCPnOpvgJpTbRiFV0vWuokeCKm5tGMTtSrwxpcpA00wXn3cyAxvQU2
VgPkpdoKbI0zmTyy/l/inywjgNtTdGeZJUU99uPXLuYIcIP6O6bkUv0rPw+mXoKecD8QCuscwQmB
LoOwbr/Bj4OAtZpZiLrI7qbF86h56eyze3PaU45VKO9h8dRNiEIl+W56naNlIlBrMhnEYa5CGoDn
u+38IZE9YQnZD6cTPDKNZNfVkAs+JtuGm6vWjPdmuSSiqarVCBMeWFi2oKJpihlKiP/JwGHMRLrG
oYZ2vPRA+y3H0nCKjhXo6gu83qqV1JjltV5JwdVtZjj6dWr9PDrVucEl0prXdgwgojL38MUBllYt
3L0B4HbxqGpbp9WhSeV2ANBepkzrKiDS2TmXLJlNTByYpY0P23J9Ah/1Z64QzQepjsyDJL2jn/yg
+56hkDwYeEt0/mv0Du2zfgQKXqYJl/PUH1TlphG14iwU2CesSYO9eHznZN9eMJkNvr2f4N8aRQGc
bzGVM8jOyvUfl7HJAwLK0G2fyblwHZGa4V3QfY/45pM0rqPLF08whZtGYNkvbT+FwIK+TcBcdyr3
IvcucL4NHsLXjoyYk0se4r8aMwsoXZAgCl4VcLB+/BSAieT44R3JEp99pUdZ3lMLaZhDASQ6ug23
OtJuwYP4uuFvr7tr9FE5+IwKYQa9h9RxxQbiuzRAkyAOM69HrmRqZmU0A/cqhJWhn0Q0cgwpJ5e/
7xKKt0DfM4u8WCWs6xAM6Z1NAuwgpjSwcRVpJ5ZOIjs/s8nOXh0Eg4qDa5FdpOp+Rn6IyhdOySsR
eRcUdNplNsca6kh9CByOHnQIh0zfRIZqVMxGsY673P/ahTuECd7i3Pw0vLSAe24Kw7M3/4yrDO5/
eYmIZgRB1dpP0mJYRrxjhcQ5t/gRdax2CX0fCzKwHV/j+aLVW/YbUY+jW++NAYUQF+NsGn24p71Q
yieOfEpOH2WvmRLhmTqBOOmCLqzjmnsCFFrf5+qj8gp+ZtpfUN/kmDQSSa7injz9U79o759OJysd
rxbhsUVFradNrjENekX75YpXGoXLIFBXv+4fIdFt6KSJIcDZzKDDJ5hMzY1mFd7D40nsIXdmXy7N
okm8CUm/2JT8ClMjmj1X/eUDSE26WeqDKMTNhz5hGzXensuJ2ayLBbw4oPjXoKma/S/ZLZYyo2Dq
zPQZ6sMAYThFAhDJ7jjCqKGYUY5OHz0o/YHX0Z28F2BPWdxWD1UEIaJi6327bfkUg2bzSBJO66Ox
pI5O907k5WlsmrEIQmwgG5Ojl2yDJtK01fddK028jEbUwCxch7MhWGQs4Br50l/9cMcIpXyZZSzu
Gpz/xWIU/3ifD2gURKjL3g5TxIsfckUgohMppIS7Fmyck6t+os9IjpupudmHT1wi0jJnHQIVMrIX
zupayHQ1zVkgGgAp5cmgxEZ25cg/cxJm2alvs+9USgmyCcwZ/Fs+WcW0zKEfpGslqYHDku5gABlS
sSkogLHPWfxzdQFb6ZTeYPPNGJH6T4DQIo06JwHO09cYorXlvG+bSrXAe1heel+xAekeKBm3Fk+a
IgP6WzU6fUc7wylNhbm//ZPK6CnMhR3CZoG5DlNwNd1DBJi4qfUikV0/MinnW47Ow927AMWTpZQS
o7hc55LIcFljckS/pvplSSWsW8mJmIxn+6d53BiNmUWiQGmCGsoD1pUiAf4TDZ18IBC1ImI/OkuI
Aa9ylFtuo3zl8IA1l0aM0qQxHuMRCwGPvNYgAiIGYicMjuSKrv+4kMjP5YY7b1lSWI2U7yGjnPCA
4RQzVQuAgRlwxE3KB03M+3Ok80jGTG115OPMpJlyejKJVewc4Ucg8wE9jqLcSt+h9qYCYMm15318
u4jWH4/ZKQBjuw8QRjjZDLnhR0Tilheg1SLxryhxXHoFR2W+nSFCmtktVkq28b595zbOA8LavMr7
A77Z5zIs57atLUs+6a6t38KCSBYvqwqYz6dn6Smfnq2R2VFNEB6ux1O/lx0O/iXRGKfg4NLgIAb3
nBTU15TEvP7URG6lyfZoZCbasJHfQX/IIOm7ZK0iMoOHKDLbnAVxLo2FOBvp1z7bs7EBOEMaVSGG
kVInrhXBDQnCvzCMXLsk3AmNXwGlVMdzshP9RQDLuZDa4iGOaIuo/MNB2AnPnguJjIzeVXBl2o8+
e/YI83GojYChlHwEpeb/ht/5XOro5lGR1OX5vnYJmDwsQrN9Srn6tGU6e4HyhYF26VhtLZRLJoC5
8n9enOp0K2NKoWMfEyWXJmDEUzAiCadxQDotMXMU+MmtjfdRiTojNtdUxg9WheO9eqq8FaawnlPA
JOpHxirBLBPy7fjuLr/rKgH1CGEWIG1iu8whD9RDYsVGTItZXpDMA2jcAUrvpYySlscoAvN12xv3
ZUh6sFJ7mnk9PfX+vno5jNWTYHieLmvUY98GMgG7NiW2XdxtHMdhht2B/sqOwESRtE9dckOOzq0o
Rag9VJ8QnMGo+K+dLqdcIoHw7DxSclIvkXVEgDiRNWboCl3pXcKsgsynxDS9Lrk1ljXS1GsjEi0G
5Yxfhi3btIRB9UrKYgnZOah6OlsZgh3Y1E1FvzdHg78WifdafrKGOPhgsg6LjhvN3R4lmjyqOp4M
VuOMBkJiJ+81agE72+A6z50zM/GbrNTvgk6J7UZ8vVAmKxgeUtaRsBeWsd2grMcV5Q4dKDEdXCet
kHwWIrkKcOIgcumdyf0a6KDsV7WHGnmTAfltaw7+PSrjXJDlyMHES7wCVremzlmvlkPpXcAJf+hT
PR45jpNjRr6b+3Ez7pLDb3I2hAtlGrn2dUuOnzbrLFcYQplcZKYfKLKc0ykZxhhypCh88Z7DCugy
3IWbzVnrfRB3eNomFwQQe0W0ZfTKlGBo3zCQyoBLELCWfMEwg2Sh5afE2h+6/Eqh/dhg7Jxr7zaC
Y1twH2SHcDiExuN9aHq968CGnrwJrOQVfV0pp3MMn2t6/+FzF11wAZkr3Z3g9CObFCudDZNdCW1A
/7zVRWheeo9R0QVca07M/PyrBQ4e+x3Bso1whQ4A3e0F1s9VGFGe+Ajs8GFlNHCh1/wpdG8hbH2h
6xN/ySGyc8g9krZHe6hLGE+9iW87O3pJWgto8zUSF+/2uEs0NWojEn3Q4GLcD8jwIACillCT1HY7
BYlw5Yx04QdItGiakol3alw58SFTmtP84CEDxkGIEhXfXINU8KKxqypkOusEUJq8anxny1uo5PT9
ZQT+zDsZaI4alK+4z/pzKax5ypiPUwQUdOUaEX0vVtJTqppsE40Yx4x1L0LwuUhwhwxsH5fLUMOM
8IPstu9na/HNfYwbuAlqDiYuFUaFPCDdlJ+lmaqmHOIhkev86ypFS36cftEqRlxIOaQy5+kE1T58
JN6bMO2XkDj7hklweLDbdHjB1sYu4uCYMwil9g6mC420IHM5xuD8tgrQm8+V5uc1WiE4aJp2uZTU
y6VtqpWY31o8M0czXRc8fu8AzRhh79z6Ckyb57Xl6HCS2UQ9b6Iw+Maq7RVbPIHaDWrz/1+BDi8n
DmAudAhtzQUWWcJA4WP5mYWu1GsIBC6+w88YRKLqkL/5tpOth8R683qUrJU6G8t+Ul/8ch/l3KiS
9SfJxOauz9EInQHGdKUzvXIaosTekL/cneICI7J3fISuO96xJr0lbkBBX/GVANVxDC3CB5ZhPBYc
ANpKt1hpEol7QLT4vAIKS1leYQAhNKg1ZmXNyVqxaHxNCCXokAM7FV1lsgGxVDSeCna5BYPwyPP7
Hx8Ys02V5UNUhY+9TyM9XOD1RNzohX4yKziJ8gICwk6k2TEunphswbHsMR18JNjlMIwh/gnEkIAw
2orlwuXW7v19JVmKM89Ukjl8rQiyLkMgkuXNLRt1BtPKGB2el4TslPWXft92DMo/zLixmaXhynGI
dkjkocuz5jdzDIxokpH4RU/TbCl9ySA5lmmROM/dl2LSmss06DLZpBssVrdMMqfsOYlcTHvwYOoj
1SaqwUWZOIBeJjfgUrD9SxQB+SGlGooy7dsvMZPiPcLCzYpmPAOyZD4rtrG7me7EDRO2/v7n1tFY
KYEE6dqzkJxzwJjl08m+k0O46CzGzU1u1bhj1CbNpV4VlIHNF1DpnHW+m++OBkWX5Zfe4sS02ICt
ORIgsYFgjbrvM7qe/hWTf3ozx0DLcwlReiez3Vh0cAdstkFUu8Notc+e9E4cI0/oMCvSUq36VMG9
PBEpJHcE84KyduCdIAXKKcvSjSxP/ZTfc7tEEqyjYKEywSi8vnXpxxkShPoywVbCzULDFFDaq++o
Ztt6Kkri0RhCL+FF+1/E90jZ41SQv87Tz2A5oYK8ORBAeTdM3VteGvy353mLIEs1i9I/8jqT+eX9
7hjta5m6QB4nc+QIlMi9oUIe59F+p8rHNvCOcaXiVO+CPqcjKnQ1BXJYhy2sloLuAppJMU5D/jmj
KwHCti/4CDhBm93mUuAXRsTMs9BmJc8Y4v/vFG6YcppSxJBT6OLSejBcIedcHDmZK3EfBxZyB/XL
EUuFb5IS+70zV2Np+rEErhDR7FgGOO+fOGzBw0bdIeUB7IWu+6FrUmkCRw7qp4V6anLd5iBsn1/T
soQLEBtkAo/Y5PTN4IgCGxYQD2xl/tClUKmG5uLd2Hg/6DdyufOKho9Ghp9nERDvOakCLEz3+/YX
JMjG5Gdl+RET+M6upf6xbrmwycEo3xGITSqbu52xR1ixABmK0cCdhj496Mh8MhKXc6ctQ4ifhGgV
PeynsuyPSNG+4qQ6gwkpEJtp+g1PpzJejbOQM9BqW+n1A7JTrd8y6egQgolTaXQQLh8sk/x5ZVUx
Mi7W9wcAAv3l46QW/0lj3Qgg1nDK7aaIAB/e0Vlq35/aP/ZxvM6QH/nOJ0n+otd4Y4zD/f+B5SI/
qVVdtgc/51AOUyirJ4wOgNSGNUYKNi7W5QF+Fw6X5+y8bXLW4GXneplsR1/ikhlfCYVlAYedM3e6
5pLRZEvtc7UFFmiVrZKITQ4D1yqCdtBMaYOvSMPrmsH3BEJ4Ybu5PY5yOiTkIzP/+1U9vl3aingE
Xu9ZYb5fH9EobrITJigQfWRA95tbxqkFSgCmYPPxyPX3ZpJOEeTJ1sRaeTyot4QombAGpMXI6+bC
kHqZU7FB0WccfxbugXeycBRMQYWDcNas9OaPvf1YyMJEJqiJpQDgcpQolvL/S57yedJDf0+PLhdX
/51etmXubnSYH/2Nt82Iyg6GIMu64LiE6fckPrDsJmnoVBuxLcPscx51FY1HAMetmpKBIBZ/yEDf
tDi8k9QsNNBk5X9NMhytFeOkevTpUkewAqXBVHLosDFwBhSWGWUjdf0TnVfE/jZyLTcJr1uaRWd0
to2Gy/Pjs4Hs1fYrg7E8/9eQHBu2Fmw8ofkY3e8gRlFW+hdQjoDL9ieg0NVXj+KT4g1e8niV/j9I
y4RqXmrpZjy2f3BxKdXo0JJ62buhozd3EhYlOEKeRs/2hmzvKQa7DA4ACdZ58dqMSnQgFJVvSJgN
FWcnYtDctkQci8hspDOEHmL/msSq9ZBlWu1MVrXzUG2S/qoqJgUcOjRwKS7IxVjWIQC/aFFNsN7z
TWLB0KtapfrSdE0bP8xaNRlB2TSYmhzXmPuIJZSUrRGIZ8MZkQo0GmvG4KL58p1kfEv9fw2D5IVx
ohdqD2ns0QoiV/0NfoKw8JvXJhJHd6cnneCY0mRHxLW72Sd1cZliDMqaYg60h6Ow9OY6bcGPrVOA
lXpPhanCHKn473VfSaAJg98t9kzWDykHjzgoRRv1T4wBL2WK0je61UhaDrmbGkZT1NvM/DY8jNIH
oPSMCrYp3REUdU/VvpXFW6Zv7fukVP1V6Ypi+ihCYnI70A3vltjtjGdn0CrDAVDY08RPK8nNgl5d
GJNLPGl3uke5WmZaOZx+Ks75uqZw4Z64IXTSUFlpj0nTO8/u89tW21ZMb49CdVVfvKkf6kVW7+kp
cOC2Jqg6l+Id3XFKgwS3qzep/P6W9kTM4aHv8xtCkAnUzaNWO3l3AQIwSH+ESsSQ1W1B+1EohtxT
UsiUGVrGgRiqTZl4FrvDzFTZm6XmtIpObGqxijATjxbAyOcpbbSP/+G2S6aq5WXyYw+LZh2eIbPW
aw9TcVp0wBBbOjyKhdf4RBFlIrsnyy1scTY30tb592Jw8gzPRSdWyq5ThXCFUst5TjX5qwlIrdkj
SNojG7aAyW3jAniPEYlDGTBn6KN0A4U0fHf6FD8IlB9D6HK0y5/fRl+gPoyLUAq+jcuENdZnXTfg
nlp4G0qooBw/sCvbZrZqj+azh6/x87VNDv7xJXviBW7M0L7ELCq4v7ZYICysbKg1IzPF07IdGZ3o
c7GbBI1kfxFO3m5o0raS5lc3Iefgh3kJWpmGkj9wlWVaD44BQBU0HCE1bJXQ72pnCzs0bnuWxreY
24s2cIcQnEUGWBWPVZjhBn6PlgtexOCX+GpRb8UX1q1TTnD1Z27ou6tk+jSAOrATw9t8XXTUJxUI
gaUVwdKvcyAOQL7TxpWVSpJ7Jl0QTpvdLm+KolOVqFJ4F2WjgwxixV/jKznxB5w+yhnDZXARrfau
edi+zyCwVXDa4koha0sfkn8wQ3NqIf+BmX+sGlnqS+/IrMFDVgeIFryDrvxuCY3dtOrpQ5W3rKKk
vwnEdCsL14dIbKW8tLL97UBRkeL2PSaJkBddQdppQ9Boc8nxg2URdAIWs3zK0F5xDipaHX2f55gB
W5TOOmrF8MZketgcKAZ0q2U/w5PHd4KLcZXsrErsxgiKXSx1bEMKb7twQvjMlQILvtLNer3CC/1A
XcMEPd+hwtryLI/zzbI5uKJcnnLe3zLxTgMJGuU5a4G1LdQMqI4fiiM3gOx0nSO7CjOSEOWs0A2g
oSIj9V9knZiOts1KCZpNuQATJXD47hBbl1kxjn5uKrkJ2O3U88Za2Z3xxv0a/M9fupphKKNkeEgg
GA2M9JrOfIcHICmGMblPthYvt6NTXT3wILqikqsNYcaQKQoXM7wjpMCx6/LPTIuS2Y4wOQ6Cbslu
7uMuyaXlEpTawtSmBQGlSBUo79NphnSI1fwTPLmytViH3fywNbkBNFHfpeQI2TpJEYmdRdUGvcwQ
O40M0ISq2pONAgrRKK46k1ZBsSl7bMs83dH+87zAIpRVGqToEyn4IXqQkBvlkTvyGqo4uPN77ZAU
nvhbhgqqZTkJ/EL2f311pXRrqtW5TAEq9iUwlKmcqw9jth73lcQdGoyXyOl/lBgKMs6LrvyZCWHN
hmBk0DQxjC/qN9OTkpTBKE8ZU05n80uMKHyj6L9OST8nPbPt/XzH7O+CTVy0Rf37ZltwengIdQkx
Hx1KKyg8wlU00lEpFZy5m2769VC6f/C+1DTUiBiOrrWqbSWf1itZcdc95Q2pvhXyn0w/UPHZMyP1
MubEe2519pcqmsOPWfABQPx9xLzwjb/Av3b8cTc2w3IqSvVbWsqWjxlpq6RYow7oqtLtwBitMhAk
joVcA1aLVZkGnpqvl6GKKkfEhg8Pmgme4TZwNM7csDkBT9eE195kNedGf1mXq1jMsYJXSU86bccX
MNu2EPWRVLZzOYiKSwiDCkQ/sYBvk1B68f5om0ZVGuOYzzldy4HQY91I5/90QOml83YPnASLqqyh
VjTvld+ubZ/nCzk0Am/EE2JzEKot9/taBN4scaxsiJW/LOTPukiQEoDRaeDQCt9avUNFx1edBXlh
LT1CxMtU23S7PIX1fl6BbZIql5wfLSb1zjy6tGLpNiZCOaBpsj52PTC9fGpDF+cqGFQnwqTKrpHU
vhvgOugeQcm/HqMoKRB43Apo39wH6YUw4LKNMqFpYOwVAUx+VS0pqO34nOtnv8uyvEBmuF2Jrw1i
gJ1LZH2jHOknzit0W2u1LL16ENfE16sdNLKJBd7Gy/eZ1Vp217ftRGxKEGThRF7hjmON41iKDhSo
FJe/dHTv6usu3kqzAAEpLOWjUiGsxPuF9iMuRq+tjAn4EWgHtjKvNXzCOb062kmI7G4BqHsx1IQi
jd/hvCbZfDP5zWHc6fkHwxLgqpYCMDwnt4o127qZTC7jX/i+r+aCt6GCEXp+W/uQBoeLfFzPHqeD
FnyXyTuyxEqPwze8fEE8RLJXxkIJhvdABpXUWz8nl0rNonm3FF6FPrjzJrd7KrWk4TIAdxXsNvha
IEwO6zJ6DxGlAv9fKd3oORl8IQ80Irau16ACSrZ78VzXVKwrR+0UzxPZOI084IFaNNUKwL/nYRUE
1MzACSLDM70ixIZz1Ojtfq5fS1PsC+rm8tbZR9W7O92wFYZTXb7fnkD3VCPBgjfFvBjtdmN3stPB
pBeRL7RN4Uum533YCDvmJckCJ9ACcBwn0rjfhvv24WkBCTl7Ok7C8AYFJcwBCSTa46X2FwmKNIfL
xLo3Iu0qkTyLvfnOyTrirStXGyjeKBr6/y8SJvIXMZAhXzba2uhw1ZCX7u1GVeekl02BdaFZuSwa
2nMPt5/Vv92XjcMsSWvKISO0kTtdRwophvKwD9vmmiQWAZR3lvexfeQtrrXV051kJXsVuc1adUsI
faspBT+lECXKGDRocSSj9Wq7zsIH6jQR3HrdezdPjfES/GwgtyVr8XSxCYnKzZvmc3b9zqdnPXZa
TB1hBXegWs9Y/iaV0nmiFaP+yeqoo8C3gedyh+d5YISq9nprCjxjvkN4GhyABLr7uammGLjhhiA8
aXV123KXbcO9eqrqlWRL4gt7l2wzmnwpDDcieDALwfpsH/KsK9qXjXVU46903sVJLeSbSNh09mMD
4Z56f7iD9l31VKuCyOKTT4cq3pp4WIEW8R/MWYa27ktxqLLOZpqt8f+Rvj99Sg1xQ75HalmdZAqf
F7wemXtGzxmV5P16N7jMBueOgYHYZG4xB4loGvxPdgpwr9BMj3U2Yp5r7e2vIFgPHO7fAXtUrjUq
oODZpKlPuenNgt4l6hFlxBkmvK3DlWoBDzkt3v8nutmpprGRzxcE0YrbkH2+8OW8SKByLZkhegmB
09qOrwMtBiQm8308MTXHyO6pTL8+TLr5TyREIqfNPJGAvhaSqkFQ+TEkNieP2k3lI4YhuEX1l7do
+vJiKX62lg0jUjL168Ao4B998S+m7yvnALO+00P5+CxplO436ebtOXAwm3LBQQXaFPueUvaFq2af
evzgzu95+mPMoKRNNlaKYOQH+a0AvjvBTxdyhjsexl2hU7E6CY5EIyr4QPH+Tplz/z/nUW/VAO03
gHTuDnsTdTo/PRL3D23wLhgF5+N9FqmMDO553UoiUCLZez+/I90pAR/Lh6wmSF43YmdxRsOWyskJ
Qe0GPre8QwDmYV2SWngKHp3oKmnkum20Vg77+JREVkAvRuVSo+bw2D4aFKt8kYPxmLS4+QRrztF4
SCw20T4FhJRTDGZDk/ELkK2KVXt+g/sOKVcluhB19IqU8KhrVzkLDrjUlrSkvHfCqzbFLOscfLgk
s/4n+F+XSUvQqtTjS1H2BLV44obmVylWMn0bWgTSt9COVHEtF3Mf6x19VexF/eenE2P9F86kIajx
uS4nXbmWnPfat8rpu33n9ueP8F2SnBSRNRUWHnFrry560nYh1vnI7+CesTQvxGPccCLHK1nksVMO
rEJzJpRtxi9NdeXBbZZqv05XdXJpghfF08/NyPzzRLkUjb618zpTjM7LO5EjtwJn9TGCGNwBwvr7
NAib59SNunJHBhnAf4T2vnWi9fhnoyv49hOT0Zugcvarw3kgBVdQ/NL9LWvLmY1OC8juPvsWLedb
Zt0pUT7lhjKv0pqlYb7d1kE4tlnDXTORrthiJyuR4dzof/7fOciHJM2KWkUc9bWUI8X6LsG1H+XK
HpXf4o890UpTAxUqqB8Utgo/GVG5Ixnzlru6t5endyUAAhSqaK76Xt1l5K6DqTWUpGe5bT72/BGT
V278v9qQVRXCrfUW869CHvmfv88qH9rHwN/X8/ggYlABdz23VHbns2bVAaKsRD6yr+F+z/f1W4m7
cqtchD5pVbPFDYyuVqTDREHd7d4stbwBrkf5OAxIokGq8zkpYI21M9zX5+J57ab8SEfvhAfriAns
fKxWCWCy7cYxL8VKNGiuZoFbqM6Q9xbUSUeLBKqGYvZkxdtSAHHix7yJxdmfVt2iq3orx0qMcwy0
iAVohDpv4uqh9vOppmWwhzwglRrIeC7HPeOMb+lK3ROH9U7RFqtwx3M6LrbgLpxwv8bFhG8Esimt
geHywB1AIPzCfatnXEdNkEZarn3GNJTdtONp6Xt5TBx5GY6iCandpXTYeDbIiAaF2fvc9cE5fnoY
ceF0yFQLi4irR6RI1bb1ayRqheRhDvZBUaAE0hctAHtKGqiLK/DeVu9Fk1q9lkGVgGRW3azvml4H
n5mO/SKc5lCWMzX15huGbP7xYr2hT7D6nPKOfO7RZpeA/4mKm294vLqfSgPS+e56gO5SrPTP6pmC
wuuEMNxXxMBnWXKUcEx+SYcK1m3buCGHm7sfsRnQgB0FEi46sgyjezKPD1hQx/3zQ2VI/r2sPb2X
4DKf2dJZUFaCpk0po7XdLZwulcCYTFDC5P3+xXuTghT2itJqBLScPpUmrq1PgrVq9OacInzKaUES
9q6gUjWxZv55TbOYqy3aeyD0hnyxkK723/XFMY56y3tgK0Mt63VoI+L2+jElyu8Yh6ctuG/yw5be
zU9VGdFfQZtGTQPlaz0VLqCmAsfJ49IBWRjqrBThvmUskzZr55jzFbD2GM5tASJV7FMlDW9C/Szb
KARCThy+MyVcg7h6hIVpypxIozHI8y+FhHANRBdUkRy2KJIz8UWjCC6N8COQ4qic+CYpJuRHLHaE
yoJ+6iqLMDtZDaa8yr7j0aBzA2xRwMRDndSiGiSOBuhmfE47+ue3VRcxa3eaAPHCk4ClnLh9auwL
mgv6ycNL6U/hl5EipMVYK0QY8KfHURtEaDAIq8opaJesZadF2Tpc5Aid5YCQlM1okmZMTXegFhkv
6vcnytEJXXI+9MyoNQKru+gk4HPKYwFXzMBVNMob20I0+bjzLwGseLn5VHJ42xgRk8lV7mchwm0V
rkn86pO9eGGptq8N9oyhs2VP+GQk9YPBmqPtgtN88InXmpSaJmhLsvy+Bi6220C0X2HwmENT3z6l
SY7DA/u2L3bRgO88lEVpJwIuUngTDXrOxB428SSfogACkTlcydhprmsfRCdC+yjkgIay4ENdKBnX
d3cjo/Ozq6kOr6YglRzs4HG/Ml563ggVG+zT5VZraZQ8byfjt1s30UUSlbcZpqc9dfaVAq1L9Znj
UyROdymeNaVFFOvquuKTQVfacpFeQnsiQRxDBazWjjZPKdH2v+lqrXR/S/b/VscuCpE9YYEQHbHt
6o/+0jLGPuLcA7EutqvifMuoUnifCvn+fO3MD8IUbsRCnK/Dec3ml2eLrUEGrxVDvaXeTm4LG0jl
6209lIgTkrvdOD/emgmKNg5fDqGE6x5CGVZYDcpzjYq1f74N6MAeqlLLOGyjGZQxP2lxM84580SF
8648R2IYJtN7961xXeZmXeBjTguR+0xK6hNvuFaRZkAGU0jfxUb2oAUSvQwVCUEv5P4FixZYFjKb
MQnLH1w4FOE9KM27eZ0PmYxB7gxTMrb63b8PsePKs5csQKTPLFK3Awf3DsGIS9lCdxU3W+H4R6kP
2Wt2Y18K0NcXZACIH9IWuevkb2YFb/ITfGNK4bKGLoHJ0dyOFIDziNMSzeDTbEEGI94OlUYpNNkG
c0iOjv9IDZCOAv+q8+RpUreQHMPtZaEvqr5TvEeyfyUXC3VZScTFZxEZ4pTNu4N15T8OmLwiDxq1
ljN4mjhaMii7pCyqHmEqu9MVZmlmYLD1AoaK+UJLE4SNARP9/quN5A6rLBxczjVbGMbwoaydQTRc
cBknOdv4JQaMdft2G/xgh2ZqCqqXcw+7S4H0C/H55Xk45kVD8+nIGbWs0vCuDFOXGB9rPib+J4ri
LruLm6vb8C2u6Rzk8sFDXy6Z/VzBIq2IzRUtqSWYBeJyX6vbu/jpAVPpu00Hgo08H32iw4mT6mcM
sxFXhNDX227lyPCSIUcyalGYj3I3ltPTqWPuHLxdMCqvR5stz4lBJP5OYM4Ljui6ZT1a5V+jQ+nl
s9e2Er5cCfE8noo5FLebZCt1v/06JHndT3MzTCyV5GSkZVzJMJjH/E8S/UncLGkyoqQFjh9tAwmw
S1Hy16Z7L62MDc7F4OHIlH50llwmIhxXe2vxWO0iCKhhrc2/fHXNV1JiwYowQYPkzhOEw4xkM3AI
mD066gyJteG4S+BXI/mitR46xMhtnNT97DMMzldq/vIfduZTdu5x1Zap0Tm2O8gnKbTF3CZXaiQ3
Juw1Wky6Xcsu2fCVF6YrixSjvYqUQpmtzGHM8omYwbY5iN22+IBewsvhkeRv7ysxUzC89XYYTl+M
eLlo/5/lwCvy8ID9Lwvo5Q851FdUErEs8slcxFLYjKa5slLqtZc+w9Mk6aNOoN6cg3MW8x4Pbiin
yO3qGP5nOtfiOgHMq6sx2RYft4e4ebprCWyIpblgBPjfpmQnovUCdWZ3hhAfqTxcomUyN7Tmaj/D
MIBYvbukzjMZJHSTAfnjBXqzGCSHOCbqa0WyqW1FZsUIVyDpgrLQoArHmP7J7jzhacPtk5+CA7go
XfEHy+EUec7rvve+eP2NVgBeJtQak+qv2blIc46K4Xd3/bykqn69yWaJ+Ps07qHjLSbk+poaxdus
gmFyvm+W/9X5y7gnmatUUgQjajDMbzJ9o7hJ1unAO97v1j/zGtVjQbXgxdD0YQopiQV0tdRdsSis
ZGhqzjoImiY1MDkZRpzuU5qTGx7NAXESsBhiN9PZLPYiW9rCPI20oV5hH0W+ia6Yxrn9uweKHXnW
22gQptDTM9b1ZgxIm1BlYMUWoNR7dGT76aY2IKDto3l9XVrg8Efi6HwCsyT/WS8UMLxSU0gpcIIX
et+/6+NvaP8rpBlN7bkBvrlJTlvqsMOImvRec+RyNMWSfjjDGzkqUAn6+Zko3oDnXgMBkZYttYW1
6s9xjc44JDY1PpmU2gCOu/GdjuQN1h2ZXp3mU3iqeKXyNPAmVuywcV8BwJQAByTwGfnQbvshMkjP
qAZVKzLRHy10A8Epb8t4onMmyVrSKsQNIKnfa1Xdc0A2qf7byPUYSOBxETku1GRUDajgiJ6VB5NR
WlV7lJHhcQIStB1I3JZJjjM1pmCvoYsY9HAhFevZBmCGbl22XLhO4YYyCkHE1Sh+VFaWiYOTSti/
yL8hgtQdAi78veAlpd32g3VKB8bwgPgePnOdHx61zLcIJXp8g8kZulebsFenta4I0lKFLFda7SWa
4XBk7TLKQdULv3HRM8qG6gYpdVUKq9Kb2EMeJWzy9cRTvtOT2SZUv7Z27LdgKjNjFwYNINF374K2
gB6q9ejhEZkP0nUjhwIbBMV/k9lc7AXIkn5J8l4HeJZE6qqv+TPvvMzMMvDxlMwtQRyec6rqWQWM
yzlr52AEexvSmwJMzq5V6HDVOnu0QaFaa92P9kdG4WipoKNH/7xaWaKsQA8/om8ukklPiy9j+XO6
iMfO8bOtY2z3Dl36u072S+u8k6tHjZSdE2sqmzSV7ruZcFSs4Wu7MdJFkpyxVacSTADnTAj+ebGM
ZHmlVnvvSXB3LmnlYtAU9z8Q2Ph4J0LSiB3aaWHaNiQQNu/koP5EbfmRZqngqCHjSI2akoTGsVfa
TGRe5krR1dr7eDcXG6KVMBZbkeczae56xy42KEqd3eyI/+1s4XzcwSWUe0IfH12VgkbQcvFp5/bl
D3rXlOmLrYoQg5Oa+IpLa6SO0FWpJZT4Kf4K+N6Qtzm+r/FwXJ+V9k13cN+vqxVM5sLEH4DD+Hh5
xCGFI1c/21bV+i/vxmqTTNWBA0TDxLRyZa3Uw+FBchgeb6jh62in4+EApVnq9i4u6fKmyF0rnjhT
iFWNHFaDOba3CQt9Pm9VMIHLkmaBj2bb4tQYk2p/VvxoyQrCSK9T2TrCN/0DQ0PZxvYB90vx25ZC
OpI+wdHuwHfT+on+FgC968mgqbp96ixZGna3nAFjaRd39qNg7opxYM6m7eRPuvL1A+9ITAaVii2s
d04xmNkq1KjOlvYBFxorkde4TBb+CRkVPKx1LtezIXm3tIBbOPqc9fKnY8HYzCYDUZOAfHl468uL
5pFG8IBokQqFb8okq97cj6zb42tY8FeYj0nvwOZate7cmefKG8ftfoI5Lio7+u4v+ycmtQMBJ+r3
i79UdCZtAii5t62XIu8Mov04P+vmJmLHdsPRhBhvPThFtXCwxBO1S+JadWU+ObpLxdDxGSXIcse8
Tp8qtor0SgfwTUA/YYyTS1xdrVGsNVAxtrkV2TOM6LTiRgsiIpsBr9SJTSwu78Wqa5kVTBCfsnNP
oaa/Zq+e+c/LMm6e1e69fx/l+3MJTs/vrzD+p7RBAma4duvfpYHJQvo1Gar7JnEEmEhUMJgUx+ZL
BlM8kiWgqyoGIdBXakgFUNBV4rN74T7YK5NBw4++zk8TTOvuAErk9gr2mLRGIaPmVo0dkpQYNOOX
pgMCAPY8EBDhbnXUBcufd+bWNLnz/UMW8S3+guubL9Vs83dSlLVLd4VO+/mgvzTFmaDYSR4s1Lv4
wZzJ0IHzO/qTYdAKzpwLXo6LdBWQ/jZmgz6SKQ2nKVgwi2oTEfcy9TxbdSBDrzQjoBONQKztZt75
bLs/BPRIK5Yiod81zdMVBH+FWMO0sEnQcsOoY86CnCTYFsGPxZqx/9Ksj6YGocWsJBf5AfeOFlKG
93YLjdYoB8CHbfQDzcV4+sI2q65lyFYmxqMHOyYBRY+o1hdVT9EK9IiSswb7fTn8YpwtRFL6KmZg
KXViby/fwhzy0IQXk8lKkHSOZG7rZ7M2jHUcN5URa+U22aT4BAH/cc6K2EzrgAdmXsg6wHPPT2GN
UJjdrloY/VTkExTLSwBZkVuPROq9DLCd9aIjesXJBy6bM01E/xFxG05/DuGWLzYhiklH8WqKGi8z
fM7L3Fx4n34YcnS8r7fx8/F+J9wASMkLd95TEvEmKfCmDVRy9e/HWA/pU8YQwluBt/uFKxLmKV6C
OpRI0oPTzq4aF5slM7HORPFjv5ipFp3LWNgiSsOe/6hWbnzAy+wu3I5QsY996uXSHlYBV3Gh+1Nt
16PI+PS0wX1b/iK6BROMQnmsGS+rKyozyX/RSzXh2bvYpRPcgCx9oCSKDFQZeqVFNFa5I/M2qSdS
2Mv/kpG+UafQc32+fUpdGuv/uWGQVaSPNbgDx/3T8TF2ymZ3tKCLIlNOlaLT9lvWKeIGPogYjx3p
jCIvQgUX4hGgzdLgx7LgV48gdgVtQHw8VO3f2mR8Z4EOrtn88B+cYEa0koKodXt/T30M4ysGtVV9
FWv0VfYaGR7hFg+ry/6gsHx8AwPF0ytAgRGTGdG3gehhLBGaALSSLA8NpgFr8x40VFZY3iEnyCSs
USDiUGI/u4wXbPqkIwyC1jr9BFhpYn0qFc4qArforDcl6URfbPiLV+vJuiFwCgQRzHJwrE1tpc/A
9jmWQ9/tSGxHZ0MGV3S+RLlVIFLzRuDzThgihrySrwuhRvAAT/UyJz1wxLVwTnaBEmbG1wekS1vy
2C1Q3FXU+86wIa7ItXmDp8N8vuRfYAcY2JwWAiD8CdsweZ7wfTqrAPjw9HWmDqou9KLlcE6FPrAs
tsPpwtIJ8l5fEdmvawkjujAm5XHnv6Xnp9aLCckGW0dJy8GrNWxF/HDlx9E7xddwNAKEzS7yhPRM
e9IywYefq81Og8wx8yMd6NafZJ4/8l54Fa3ONsjdPAFjE5dDAI3mO/F1FX1mFcC7gTxo/0C7OReh
HfUXLpRE+gfFhhQSHBoKMjHsbc/Vbtk2siqxKK/7enMvT/F5NFZqVGB1WVLisHTZRwO6KRl56BFO
KnpTAC5+NGadWqPs7hggdw+/QA14qu9X/K9wc3GHJsGGV0Z6MWNP81tFpkAdHcp2aSK4hYQ9erJv
UYaijz5JKnrCHheEfW2MiIaNqc5J6zgRnsYZHBl7pcgfggP9PVNjrj1vh4sD4K8hV6kSJUGsbPa4
yYata6A3KqxVFEgnplGMbDGNbfR8cB+Kle/UqftR841+8v4RMSlXCUnBB59zjf9Xy5V3xa7/BzEu
b4bVxbFaxZtBlfVEdCPSBarCOWYtGcYvuuflPJ+Rr5GR+vAfKH5C1hfZW97abR3BrB6APy0W92Ni
Y4nrPOIZ9KP7ogmlCJSQhrbQ992Oq3b6/ZDfQaUZG2i7jxpbBn3+87znnvedzdNRni1cAh9tISZW
cNvFvNAV78/H0KO7RjSMyQwMnJAg16s9WZgR7/MZ4H8PpDfxXMCHZYWtQ09LDPBpxm41u5k7qf2u
dw0cNJ82H7HL7VjteUBZmSgkhaVROCO/8WcK6d3A4T2wWDqRBQFMDE10KpEVdKswvlszMYE1F5CZ
pQ1PH9iQObLkI75ecwwvMZhUp1Ul7ofD0S1X4HKZcUWYe5VxbTDv3wTVG3sHzlScyJkZaAgHD+io
3fXsCFhmLJKa9XmUDslSaFt405WWiqYixZNbKkEtMFxJQ01xUMnW1jek4j6ckMlBKSO5QNgSnn/Z
yZIcBGJI0xREkHhEU8qOQH7XlYi8CBwkAmssINXKy4BatvcHUGQ1Y88+sN9vzMoPYs81Ll38Utjq
41CmLBPFxen8rkrNci97UlfYLMIVUKrTL69UeS5lmGqlS4ftmDMHS0QwS+yUje95ZmKwP1W25N4h
YMgb8rclAhe/9aT2NbGWxkbzZynSBI4i70/xolgszx2SBkk09/AKVJxJbJLH4c0VyKTVmnQr9HM2
tC0QwYLTyVV5cxRJx9fdf+/u1p7611TYSReIFYSjE9FBMXd8oPtNNwtz3xUv9UV42Ssl6V0Gv9ry
iF1dymeg3K5k3K+pQGu00G+8ahcJQRpm3lhyMIVdADcoOrLANbZyzAS7xAJAcKw+cBQ4wFTJxSjk
i/gCnd6Ce9Xc0GllIS6IvaugFhd5jlJ8299pfGz7NEsdnSZ5wxJS27/ToEedJ8Fwo3UsUD7Yidow
ULqV0jOtfazIQd68eLb8h48mu50cM+F9RuuGwy7PbyAPjM8Kg6/urNcn+VwMjoNT0Y4bOzCWWjyR
bX932P3XKyVgC9PumKcAzSvS/QqaN4PCUwAOP3TwxxYwP6o+zzFkyP5JAOaEnRBG858bJUNL4lxs
3gpteoa3+3fQ1N1mVqlXLfpHKc+/1mxTP9YnpvFA30XGAU7X3s67WrRr2iapd/H5YoymooCTfVa5
f9ber/d1lIwKRYVBW3qgND7CcyE/ud+/AIezMfMBVoAZoFJPbl8WEYnPAI62tdAEqaz0U8AnkYcB
nukads/5VFbEFqOslIvD1lA0d3QtZono3XVnn5gHBZZ8dzgqg42NMwgz8XsZcczIOHp65FwSt8ZO
xgw6Js1EODPdI2o/R65NCBiyY0VoaEVvB1I6PdkFhxDhg3HfMnTQ3BoVO/mhiVtuHAb4Y/ZONy3Y
xJTJoyqpY1lTmd491CDkwH6+flYazIJK1BfJKpjFKJXWT8oTVAmyUheqsY+5v3wWJFgtDczbgIPF
1hZ4UX4OYj1drGdN8Y93/4zcWInAO0mC3gHQC5IUocis4Dma9JEq6/rgGz6voTnkNDZFlM24Ck41
WeOmRX9mMDWtXeuleN09NXGwFJD0jrRTwnwWA4JHPoNSH3NU9z2J7iXh5lMPuiJ9BQTQMGaA/eRF
lnxzur/UlHkr7dV4l1QYLikoDxZgVo6uj3fMPgQgM4k9dusypXzU58RQ2FftXgI1ofio+0m3jIjr
LmuoCaiWW/3BUC7dX4g8UuFmW/52RIE+gNgyQBs7DQdEKDXTYbNT2CUA+iZCU5/N4WcSexZCCZHJ
QayW+rYP4fYKZIzaOTJlCaT/C1ntagzoWA+JLhRp2BgjD5rV0ROvTFLtPAb25LzFcJmDFUrFuFpE
jMTU6jZOEBXt7qF+3lgeiOq7I2E5u5kPZWxURp5TnLpPSfoI7sTYWJJaSNgI9GN1aOY1Np9THooI
0X+/ynkKc5DNF6W34T7Ewma/lsWHfAZt756TbOijnItdBajSBv+TIjH4vvidAjYcpZZVfjSdEejS
F17m8qlFB/J84e89Kx9VVreVFSIJCepzoCtllEGACjNRkBE5qa3yCwYY6FFaNqjcF5dKM87ocOLz
/ifV3K5Puw2oQlvkYNXVaTi/AlDgnY4E2mOEZ9KnLPO78aEF3xGm0J6HNxC0lnKa89n7QcbQkEQ0
a9laWE2qCYM3PCuIQzovY7yF9umAWsh0YoErEhTQPIZiFiG/ANBopt9GUiMimeX9mhRMom+T6Hmr
ilk+aw+vqeq3xDIRUnHX76yW8sXT1xfsOP+t6oM/1T2yW5Bs2opLc9WZArx8SQD5NVM70/SQm0/M
SXiOYoCUhf1vQUyzoYMtprNNRUx/4sTrGJK1OHUi8N5mz1BroT9JXsM8FIhWQeTdXGuZ27ongyf6
5uT4z7weHwrzhyywJIxjXa49f/Vo1DCwkdRIWUVolvberZDfgaQyGxtQtb62EL1M4Hl2OQn5BxBN
FKW4BQuMHHO257y60xMv9ZtSfbZoznSHuxWlJyma/zIFlpU4ar6ST5UWZ/cRq7LI1KGmeKAnrUtz
5JfAWu+/q4PqVHjSJCIkanCaYf+HNftvd32GzqT/Nypn4J56g678tjdM2do7u54pVIDszXHbsaii
bWHHiBMgQEzGSmTIW7Xp8ieD7shlqEqvHQUAeY6NfpvWI1HMrBnN+lnCj3WzUKFHIj/GPqpnVWJo
0N6FLJvdIEWi9Xip3K/1feWXr16ZO48O5AdllpY+Ryfl+3p7q4hj1NDC0TkFj9X5vIfgAd8h2Biy
dnmwiikc8tFcjdZoNSXDKEMI/5U/KOtluGPKCaQl27G4DxeiBbSqHi1rCQNFLgKJxwzJBFzRUfsd
fLtbczUKRlthpuoESVS7PZgL/HXYB8KS1YfiAOJxFiZSqKFEctA9Ry/1PUgqkw8wUcUbdgkD5T3A
QHuc6Nvru/dU9MBodYGmdOTwjp9q8bCCdHmjaZQNjSx0RhwGRD0teof6R/AXKXnGlVPo8GTDs4nQ
vc9O33nrEtbN0JBcx1JNHvMV8O0gR7THwtsCKQsSRxcAw/IAjqyyEnjAKMi4gdT8opHQOI+EEmvd
WuC32c19DqXT8u05S1RbOSSZuBGCTm4dfJvIAe62YD/zqW32BbTQqE2e+ngMnKKVHKDtHOia0M7r
yHSTBN4JZMzO68N4NCXWac4Zy0NeLau+I+/qYEtpEOkIGthDkWzXQeW8YM2zKyTAxFAJo2Iq2GUU
esWULjj299/nLMJOA+SZG8mEcjh9O8RvqhbVUkQQq7jVDyfxZk4wAvyJoTeQqa3dCMo24cBUGRlD
n7LwzfjkE6xGJdSuxBSsybMdz+b6dmTALGavllsV/XtG2v9kYQwd3S1MOGshk/hEFYAeNrTOxVxm
mMeSAqxFaauQNMYU7qTk0iQIlPKN4s1fjq8eITwyvDgIeZgJHVIDLcK3PbS5ZYgPbP3PBHAyG8jX
rOnrLowSDg9DPjQL8clBeENiLLv5n9F36E9fU0zdCd4vTvwijVyJeHnLGrFDaOBM4HXxqXbvMT49
IglJZTV6/V7s+k05BIx0yEa28aLFIpo7OqzPyhzwJQ1NxOzFWXBxdiGy+W/kZ0dt6Dq4q/HQAi1d
atSNs+K0/SKoOs0SZs+mGx6Q4jp0MLVZ6vKx6cH7jEzjYjXEWKLu2P4vG0otgwptTodpatDQyT4G
GYgeuknGDGDb6MTC1Xo4aBoo79pDThc76njOwwWjZqVv+nzGcFL7ebFpGHuRpwCSZBbVfAjyAlXd
1j60vfrvXGasMutzqynPLGm+KdQxnu1MyGnArjVESoyRbHz+gFT59bAafVSrgUUG40xoib87pGlH
ssxzIWVtw0T4++CS1EeNUnpoWq6shS9X24yIUNYUw4OrvhD9yw6lpOA4fScpIQA1WRXh3Nu2XBl3
IB03nzmNWRC4dyJJYbIxtOoMzr1RrnXou75oCFgtDF66NlDKJxwtJQZKhKIXz4796pMCetc0pECu
5r9qxYZJvU7kxY1ijHDXKO8w0BBvpgxlE5gZRUsfQN9orJNVdxac8XjCmYZCIw+7gQ8L9Q6cBVvz
Umtw1JDhtzrCm66+7XiBdyVbofPs2Fjq/T0dru3iyTu82EXNXFGI5Ts/sR/SYz3rh0L+tSdIDZ0o
VAVZeUaiF9866B37pxa6uYddOzFSApsY2aUbE6NtG3U4EZSZfr8g2RoFR4l+VQYdlDslZ8p6wqea
HTtnYms2cutyygCVpYS4Bw1aCt9G642mIjB2a58MqqTw8jW5yTHzemFpTn+Pi8BahNsteM0lJDiR
0aJiRQTxtyNOfAgTN0lSvlEQFGt2YGAr2dYgoAtWj3tQ4zhiG1qvKE7UOjQ8CYaZ6pSz+osFq8GR
SHHwSOZEqOIbbOV60KThe7nKIVRHWeBgilm8Q6fO5Umi0wWddFTyHN3OJA6UkOQGDe0AiYKgt2yg
TbX5qibP5G1eN9PgVYlCfHPsJHOwc6LL2wmJP7ApeEup3yCX9AMza/cQfW2z1qU2S6VnsODlQ+UM
S5EsVMO718JGIQ/8arJU4MxbMfSOBk9SdE9fKLDpnqiU5dJRMS9XJ7sEPZGmgRdRQ3Z1f5/AyFm/
tocxlmHfMtpw7L0yAcmV8TLYkVRlgS4W7TjoqPxOdulKxkRx39l2CpPAuN3xqrBWihBspi123lgT
dsYGd4+P2EPAEyUutIO1W95+eouGu+Whw+YlDJ+2fsd8wtmoAP6tRnwbdsptjNM47qf0nekhe0Zg
iCZa1mFUPh4Ho99SV1awuwT8+6nm4wE4T5blf+Bd8jdwSPNtenv3Srg9wB1guEzmylXJrtlMxfXu
YSBElN+a/dgLachUtOi5tdomvV4wRNNo0N1/uCdgt+5fTQ5fmdWNLNcR9qzBIbKCfgzSqmndfp5N
TOw+uBBUtiXVaLzGzCYVXblb2y1KgdkaQKnkknmXsFDlGmLKVIoVnLFrsvhdJ2w8C7atNC5tfzOr
eWHc7DiC2Div3TNQ/9RyI+p61ozpgQy3wsxIlVL7ll1CSTmCLL04I8wJZ06MV63D5gJi2ZUD9rxQ
LyKfV0m75MrP9DND9cFaSAItxNYnSZy2V6ON3L7jLVin++jN8/MXmqiVWAeVO6mepOdBAMh6Y38q
UweMtSZ8ptN4thHQSVxSyjiWYu1xe83c1/cbAi3wXxwpAFcZqxrTMfV5Zy5swkvcMXSf10Idxfm/
wky+Q6rpgR979Xgr+FggmyG6RFF9iMuVbQP0s/4sgCramPWiEJHgUlkdeeG5+CKeknYAYVtstD9d
jXWIbwdkoUXiMwVGlL5OZhhvaSp/XOV08yTrjRsovtLOA9woB5CZlx4PuCq2X+z8DbdPmWOcrybK
htBYFOBUBW7hdD9tU4lNPlJxD+Hmv4AT8egDKuoGIIyLdhjY8EnyKy8sOj+rwrfmh3SlwSbKHhvE
ZsOEs6ZZTmjZm1BNmNo7472G5QN8nxOsaVKjQhbacC3ZEV2tb/kTys/2c/mu1JUbDekI15wOBDuk
1r57Z2V7qBbuFtbVptHXt1Wnxh5nKXEcx2GsTHbgtEonhHVhymv/swvzIrUpXcIdxMxQxtZH2ddB
RZ702zX/R8PGD/SDztCmgP7P5qSUoZZ2Vkc8Md88KE0BdnY/VrKKE9bX7vWDUzFS1ld8BPjn7Qsx
xlLlV51UlBG9ShXqlI0jbKJImd1PB/VqSgq+3UvjXtg1PhvFm8LqyGHZVw7mGnRAgc1FIz/+aQxy
CRvDUE/q5ZE/cgvNsBpFfLJiNIZguTfwzDbeLgDRvcmTXluT8oXwQINUlo76mHUHAOamjV0unWjS
/0j8Dd+xyiXuYQK3ZA+sK9G4fptnafeVVG7tezSQZGQjCTDSDHfDQkUY6afQ+bPOu/nHkHdk6SqO
wbl7H0lHPFDUOcRiZCfDUexeXQopfnVewp8vzIC8TrnUallawxjdn6+nTAsj4cPURJm6MkMWbtP8
uCTgarhAIVanOeJ2MjRZmBSJCdNDBmwADjD6phhOrmP7ni7+BKtY7H6UNMfdAUIfBmSPSUK6iCtp
JybCM6s+hRyzv6scxjLH4r2jRXDf41HWv2J/jeNl5aPVuSVH0Kdq4lDjHjOmXEGOEacvfYnqW2Jf
08SrB6sF7e0O7Ml1xD2wkQLU0QHBW1GVPTZXDdcHcD3vPbKx9Yys9gsIma16wM0si2lsCv74TxEc
uW+N5Z3UF4yWRTrJXcqhwfUr/DWrzb+dQIrd68HMlJAKmNkH/dcQrxH3GYVn4vM+ZLg82eguOppJ
dVRhO9FlYfEQmL1zZllfexYiXYYkpqsjUrXxC8naK82U3qpb+Na/tI6JQ4qztfeDezTUPwoOH6//
I7bmU1kfrkl/RPdQpRaCwrKAU/z9C7EmBDPUrpUGIXAgDicm+F43zkCz8/zkNU0FEwtn5FqN9mSY
ap+d4pIlznMf5pn8/AusPD2zFPUHSE2QeBm+2aWbmHggTlbzC0LdpmP2KmrptlGzghD/9fD3YBfA
chYHfmmubUiMe08QkzCgL72UEb77M01MPH0O1MzApj4qNNqAMF87K6p1uvhEqcR0FuP6OFxnd4h3
grBUA2sAx/9Ne5smAW19MRZu0U2nl/WAXdLGtdAx30R3plDGdm/iicaL0CsTNNq6roOKmIiDhkxO
GRTpyeoGCggpFgVlMP3ESms0AMUTzS0sHey9m7Cnjkhw/NYdkP1Qm4fhnzpWuhLCaeASmlpibmIT
1CEuDmW28+OXWSNbMe0uKjGG8grlewDOoWI9FlOSOgvSbJEukfwfgnlC94yLtoRIKHIzsKv0cbJH
dV7+poXl9rj0g3Ow6f3QxkLDteKW8AzQAg0aeqxOlvMbywUC4LkuwkwgoYAbDpK5hoi6DhTmEIme
ueHnDrPYkwzBTnyWfamq0usEyIYLGRpio7vhf63wQcAaQY0ifEH5FXWOKOvdp7h/Oc+VP6EsWrO1
G/YPtbgOeN9ivVhHXJYAKIoHI4A1SC3lR+0ggGE2HImN9TbaBpGBpp1ThgpqWK9sRnyeJ2xWExNk
ZAUvVeydKH838Dvm3FPWEdS+/tZ4ZDlet68GxOgNXW5fK0MyWR0G67nBj+/7bWcCYOO9Mc46tQGy
M9E4kY6TRGJOysUsCF45uWxgwcOeOb1do+VqGkiGFQ0LqvKFNVy1axmtSVJyKyDUkT0DNju8hF+5
QkA2E3k3KdAGYMQlY6sDPp2ynwjZZkXt027yl+4uOWOa8ay5mTSoiKydrYvtiOi8mcnCpQSJXCID
SSAHSCGfTZsb73J7nDHgBm9mZrAxnWsn/cBrtADyWPsegNP2YRNwnpjl0OEIpvvyy13W44FwY6EY
uM1swhdV/8GCPmkG5/aHWQ9ZT74bXMiFA0rLKV2bBUnXUxZOKScmzazGyhfk5rMsKiWre4MMXdHp
NXpRMGb4JokLW6+q4V1t8poEaOXEOU59kmlxkc0tzhGhv6Dw65K/VtER5ZxDLJrYFsUnk/8pp56H
+1zjGQX5IZZjCnKLjt9cRNqvFLxcB2XkEvs0FQvG/+d6igjPkKeVhEkiamZRiu/BGdUwkEDonTAa
r2q9bj4vuDsU0izl5yXZPorM473iHR/e/hD/M1rGAYfWOIAXBkYH4y9C1w3dYAjOWkSKh0hbqlOK
bO2iXAzgLfp+wH2zcqTomJwpFDkySMDg3l9QrFsr5lumy8ubOpODRN13IfITlGfW39d4+8IVhOyF
57pbJl+rdDgolMT4lKrM20YA3iUSe8cxT/4V1uxwStSq4z3L7KMzf845XpGWXFd+0hD9XJRKpsKf
5Iqm/qci5MeVOUrEEo994Y3wgOstsBhOSHHhHBnAo4hAr4V2BnGCrNfMU11PQiH70YWto34RBrvT
GW0CuCIV4SKdDCYvrlLf01BEze2V2RqSNRD7vxpT8Osge5TUDJN8grz3m5VTNk5M1AU6679KmObg
G+Kih0EVtkE+MXuhnBNH/WeGu8CacqNNuwWDjV5rKKbMc7KfjzsLIqBWCKPYnX8x37Kll0oBvt9G
FWhU0iJUvYeiaA9SpnmQxBqA3C9Dk3Wivbxakvq2cGPj9ASF2K2/pInpk2+aMLwOUoHnUoTwBcVl
SjCtsVGhTJzFW4hLR306IY+m2WoBcBuVcXeLCXdRnkzaheZFk4J/v6QoRfQNBLG274L2l1rqA++X
cqYpzFEioqa2PnNp263Izi06oduO/28J0HJI0QNp1ijgD3qJdnyD8Gj59y9OIXzuqyMUdppjhyFI
tU1re1RYE7PSBF5mzEqB00JUMn8LRMx3pth4tkstIyqTC94ifWjF93rcMB6I7id7kfNuPvA4sB2W
SYIrg4vGJvCoWtqrL/o3V0fN+jMKddIarrKrs6+aVqaLQwllc5CQni1Yh+tuaolRUVFQQ7qBUKgM
TI5Y0s5iJ1HurqgLMUVTGdoj5jpwJsfTi5kMVXugCf/yVtQSwiQDO0F9l/+MtfBGRSCqQdtZo25K
+z846zfVFS7BQoythk2seKCi/gW44MwkuOLYBWK+k0+8Jbt2n9Up31HtzgXuaEVFiGNhx6vuXQoz
5BRx9ZrCUEEjT6t6aHmkN72YiSMm9IKnFB75MOL8cI6tefQK/yABQK0RFuoNESK90liEo88RMpOo
q+g57tdvshWz9X8spVZALbVN7ViNmJHJ/emCF695t0f6XeC/6s4mWzL/Z0i2zsvln4w66OElp1F7
twNvOthW75SpZ8nlT56XoT/HZCLSSKvk6ke1cYpjiF26GJxJbuMo7bzCNrqmQGgqlnuwsjHxHtYy
q10HNrkLtZlj92UAR+RXv9hi6gve27JxQ8cFdHqPd3CkO8JI3ek6r6Kflz7laI+aif6NEf394/dV
CeDS6Qh2lqQ0G4zpXznyNioQ5TlUP6DwUT+EOstY1eTcDAs1neUDrvHFmYn4Cnqd6ER0YEDaYWvs
7x1VuTYWWd117o6Pnnp/Bv60aeOp1uHnJ3oCJf+ZZwdnhSUSrsLpBfEFbSSymDHsizhS3A9L2O2l
ksvF8HZJhtQWvdk9N5xbFjUbZSSWpUHZBLN7TRZEgZHRhB66/3PxYK4sT+DuaiGwLrAv9DW8/aTf
SC9JOpqtg89z7C4OGmwraGF1pKDM/ym1/84tA5GxV6Wg3P2hveWvQgQ+vX3qdCvOrKRYVRE4mTwc
NMnet3UeEYnwng/zdbD53ye7+Vlim+e7/k5najVaXc4eaAg8wHp3sCa6dAchbk8FzGiNQma7ZNMY
2t9zy9aLE409wJwZbyvtdsHmMeq1xJDdrv6hUw9ag8Em0e/vySajiT6KCGLYBu6JSG00ZZPZ1GO2
yh6c99+UPhhRiXIWHmXN6vMILStQIgqAkdTKqobS+0pjAclMAQYQqqxo4WvB3wRFGeHLXkW10IG1
0kfveQ1wDdgEQ/VVFLyepC5XkZwBVi9tl318LWcNpSMrU9YRljsw5dEr4AOoYH+bsrsHVIxrpIeB
kq1AzDnx/w6x8ke+rOKp+MlkMNnQ50tqHFD6DOQtXYyXoejDZUF2Np8cOm8awpez/0VUq6w5jNGs
FmXs7PCq6qNfTqZNt0bjeRKsEu24uZD8oiltfdMbMfFSM1zeNchnX6F/dKCe6d/8HU+iZ9pq2BMg
ZNp6dvWgYTFbhz5/30w/xCtpY1ulNyDm8QGqv0J1N+qKM4xSv2iHnU4japMggyFkS22XLYBeUuX3
mqITqzR2+8tzBbt63arEs7J1MbvDEdVyJVfe9m+XLZPBJCGuIJwZQ2Rywpg8QBw/00GZqiPkViPc
Mke4Na0Raprc1e2TxtSVJbx4XpkYxYMj69GuIaTzecObu+FlTk7erBMn1vnM3fxrAktUiE7xd0zc
Ri5LMR/DBll5D9wFhcpaR8ElFGq5rreXqKhH04Eqh0KVQb5XNmcjnTHX+6JDeMrPtpRMQw48muC6
E8binFZ7W6/8HP1Gi1GV020mjYmXHUL4q2PaVWz5JRFyJfBuQ91rUBKviZHYaC1epBAQAhvo9k5T
OjVymxjjlgMbphnYC3SGbp/ilzPWJWfeqEClUq22qVNHUu0CUofQbMnw6ZOLyX3w5lV7otFUfbII
MY/jQ4JeiA7CedxWx8Z6qZPQrE6j23yWW8VBPSqV9rFsi0u6apOQjqMpJ1jaiaRZo1InJaHi4R7P
oh8Nb7SNLCXJflQ4TYL+rJai1irmYvdQSE/8yGSNiaa3swbvfbvgF+UMXmaIfa7EipEggPQDrLHs
FumyXmhyPBSC9W0E2eZPBlSlhS/MCvVmJSvhah+6ZF+HIrtVv3bUdGNqXQldfXecLX1+HYNx0Ek5
8TZKlcStV7YElWoMCeaWGGuoQrzGPzV/Aw1v1eoyANhVhcphnwoS+DP3yVtw0eASPQdk1GM3e5SH
gi1Ov5mjYyD3+usvtgXdQ+XJX0n03ph2afkM4kXlIaSFKQeEbyWHERD3Fch+HfkFxJ6JV+fufvG9
qEO6FCP62/KiW2ayf9iDzTEsYJekqCEF1U3k+G268nVUiU1g/cgL3KhPqWdVsnboYZj4dPvUr9Pn
z+9Cq3BsTL0rdvynNa9aMQLsnc70BqLnhBkBtUrF8gRHpjqj2LDu+8eN0ZZEbsT/zi7dajThCDjK
mjZSoSMdMt9Px6H19GNElpxhfQAna1eO22bl1HEvpPJa2WUZLPFxxibj4iDSydOGRrrLnzxf+q5C
7uSsGVpcHq1f/6tzuwH2fMeissqJJ0ye6PPq8ixRpEmik7pfkufNSjxGdHyZX3nG77y4pYEDd+GY
fNojapcpGYgsj1H42UrWYBKecvXw7aonYOuIm+aVEaZIzldD2ilwzR+qMaO28kXX1HQoZveSp3/X
OOMnPFm7XWtEBnVAOKsLT1Z0aw1nc+UMHsuUmwMFP33OEvi40JRfl3u9eRssZ9/KQyBGFiy/EK2r
TDqzwuYC8J/lYwXFLYWd1zhfbXXXegby7zOZdXVMrAc2SiWqOYy1pXSiP5vbKmSNHlQGO/reL2C+
cWATYhLKA1drcevpSIZ/AhSprdszYdI/ujcwpPKtNCsZQ1agEVynqqeH35s0HH77WRGuRJTWM6aQ
36YtAEKhtBa7gYk2SFOc9m8LQujE5S3XAGVrFdubFEysUlgIISHk5vVHuw6jiIxIu8KyTT0XB9+l
9y++ONKxWCNpw0+ZiEw6jT5/TcsGRZu+t+infSbAtUZRjljHpF7E3mv8RXn7OO8QPvFZi+A6Xij5
ENrHd2ETwUMrloRke1ygfJooRfvx+H9hT5T2bZRH7kpNOwd+z5uLWAa7SWuJj+/+h/kDM5O5YE+U
VSZ6sgpucKDOIzP9UH0Zrwqem/5WXCU1w9BEVTCqf8l+yw4GHmAkV+59YQWCFyJRL8QBLDrlPS5Y
lrSr2ISlsRWiRerH/nNRwNKCWziejQMbKMye02mBnpYAE++8wjx3nn/RTMvqbT7UIDd76Hz87M6y
gXBcuCKW1xXx6/ecAPKvq7yFyyBwLKM+5RioGRGcU3XrlK0Beqfm3Pkq+RMkbJOYo5ABxELEEWi3
RG5TNBJ68y0+ThSKqciomrvsjMReRqwwhB07vjHQxzy1I+ZBLSyioCrz2gETTG3dVKwJ7HL2JjLx
DACpzLdkL8wmSLh3kcSJ0rXbSXMSqJu/CaOLliQK9w+RngGoP7gLW4iEmsCkI8rkK90usrSYz+V7
rB8Y2NxSZVVUYtLuq7Rb7a1bazu8oNyvvOW4VmjTKd3EehR0GfDsfVIV2IVmIHhsx69l4F/mbSAx
YycldEiyglITqbL3ZUW3mvBQLqwepo1afeZOzwTW7jUoY5EAggm+Jc82IIlwSi258u53iA6Qbcu2
TxwgljrQ+t0o4SB8/An2JHO2tvsQpqg4TXMzsPEuYdkOBqSq+AqVG1YpDflENlmIn+yFLAxtutuI
aVq6KAe3kK7QKJTt2zy/Qakql8Yyu6Hm0Pmn24UP35ay4NNcxgKA5tAwDX7QBqnTNWNyhBcSty6M
fPgEUopUtdl+hIsQcA5/hqrbmSuQeLsI7D8yhZuVZ7xRsuZhnTH5btZcV8rhyic4iGuy9HPPkc+t
NLUv7WiNZD7JbeDU0g7sqyYu5WVpYYlvibbBYFbhqYMaRLCzKZ+K5bqxkyf45PDfajEdNoI8bQG4
KUVeFxqslc7DqZU0QpwyARhhv++FcG9eII/1bhGY2oDHLMWks3YzV2LLiHYQbPgJIJ7lEzclphxq
CBTsX80L5sB/KrjtkR4kyhJA1tBdOJyNA0YpIqNqfZSSmGLpHeZ8UHFQbZ6Hektf9T7RZk/ViX7X
z/YkL2GuYn67I6AzFNudu2vzS8uOTStGDCrJExOfv3s0F/kLg6d4ev9yUmW5Enu7ePWxH/GnXNiZ
s7YchdjKavHQJD25RUXast7x5V+6/ipADCTr2mFvuFOztKJ9tCVahkUhjr0vuAvBP7AdxDubsHIw
4MlHh6vKZ5vxfOl8RtNZbUiqqrNdLauO5Ov7r1s81BVstoy0hFNiyDxlR+UWarcxdiNjdw0xlHET
MM8YXG9lmaXrgyFPR8I63rWL52CzunkdU7dAa7TtutZ9DzukghJct85Gf6hCUrrhLbGH+2iG4ZqI
Znltd44S04P3dzQkKAdNNig5SKXHQQqZwluANBxd7G6vs2xOqY8GtbmBauAVI/pLvLc7UC8Z3+uX
MZsZlwmRFOGthi+upafHOcwrAguNMiwjRPa63/gXFpBT4eYlTwT4fYFxMniBD4deaM+Dr60tjy8e
VJ6ZhdYcVfPgE0En14G6gpMw3THPy1OIei7KqLjd592rOMWTZbASHIUJ1zfoFTD1DfL+myMXF/Ma
SH9+Rh0Q1Rev4475gAx0k0PPrDie9Kl1OO12MhZR8MTFavsnQLxG6u5/7T1Psu/40QKACB1h44uc
UaOQqfRhBHJTB6EMUhuR66oB90X0muv1h9H4oWYkCa5xbHDM9npFnKkxkZZ+OTazSPM89fg7/WPa
581jUGKWKZKnmCmOlLx22/ri22UwFyWjriaXSyl6PXVS3/bJIi5LeZSPX1ZN15v5Z1ht+2gEzHu5
gubzns0DRNIneu9wOFyOIRoSTq2aPpelp1q35jE0RkilQKhFwkPu1lEOTQPx8ByFIV2yf/vOrpJ6
eKoKTM61sp8+sblebPwV2hHQYMKSf6tq+vBjLBUvvEuYZqAeVbrNC3y8nW3iCdiftbkR02nkS5Wn
H6meEq+CuTlUCoaA4+qeP43SewIN3bOwa3BFX6RgOLlswESXSKZIWbYMZmypmoFjWMwU1Xw2NRVc
3vBq9FUQ/N4vtoHQrAoOkYn+NKyKYtF82cbZTJffEYh1EnKRtgedf/OWBBnwz/hv4jbJhs8ckzuY
DjVHrWbQtQaLDtK/hEEP5N3JeT05LIi71F4FT8cIyd4OwrHp74O+k9vezJBUzZywy15jPJ2gxFOW
0W6MEUmHLq/G4u1jfaIlMzqZgDixVNB5fEfN7O6RlxYhdwUeyapSuWzi0J8BOhmvbiffTh5m1qBr
GUqp/RWbJoV1SPL6eu8OTD4Bt0BYi7o/hVYsDCg2sdCQxzj/mM3H4WsxF0WuhSXQLbsJVm6cJpvP
eGj0K+v0O7RFB04f1rMzKtTknaZOk5zQxNUYnP23ulCGV8+DrHu1YCD6hC1aiA4mjrCwFHM1A2Sa
PAVY3fokZgVqbMKm+hE+gfp3RhBF/T/6H220t3KnfLjpSlp1u942hp/2IHKSWnn7iv9XINgBXcbL
gwfINrEzkXKRyacqBdnN6yHip5D1znOP/ULAhAkLSAC5AouryteDvqzoQDgJSV0Lw03ROjkuOFNA
E70MhA3Hla3AUxIOvKat8C2aV8Wz7Fe624yoNesaRtz3uGEB/rcZpBq0AtRLmrXKvwPdxP+mDBS4
XoW00E2tNNqCY7tM3hK+heZFpZMW2Gkf5/Sgky5f085HkR8i7O9tM5/r+4ml4FddvJ+Nz1vYs0ND
q3cxnDUAo1E27AKCTT02UhBhB5GU4fE3G9FQ8I0Q+lvPGlpSzduyJu/KggAAEM/BHPgOlnFrNzS0
gCmIbwVYoN7FiyIBqok1J7ePFFuBnJuFsylyCsl3sy/3uAFHdOus+vEhgEWU53379M1zAoukFj73
9sMTqXljACnm5C2y4tKvSZtNwVCnU6c3Sza8kAy+/OgxJwNcs3+NV1NklBKEoj2srg6G35NdpxMn
DFKfUk0utzI6TBslW0+OE0W8/ZZFd+HzvvG60GOr0lCOIl91mXiMOJ0kOlNrHqqPUZ5xmtUtywUN
8MJ1Zex3RaAL+Pq2Pa7sfRtaKC+wxlkY1KeYwd0wuQzkbAw/Qui7B4rzRhkEy/NstYP0Pg0x4hx8
7HN31uVi8Qc4nnvplbM6nCi1YAPACzZNPE6LKHnbr37mCpCQ5D6E//sxXeGIcg0wyxMe/ce6Nrcr
KjOXR8IOLUyKUUO4FKzN+lY8iUEYup4L98Cs+93BUXpgwGW3d8+jb+QMOTpwb2Y6R3oreSzHar5t
GL7B3kUjl5LvLf5Oo8hlj8RQ6/t2rzfayihZtSf+eweKHiNhT8haxyiCQxAUJFpjGIe/vG7egAi4
Jw11lHNc1y6Nv91FLocLyLCi3NVHEnwa4eaZpsI4U+6mtGgaBTa3seN8b2nqJDfoR315uJR+Vrux
xmYfAcuuT+afa4Tkn2pep6e5fVKGeVU559jEc+S6i6x6uvuctTZmX4K27JVvP3EDcmyEzyKM97g/
2Vl6H4N1O/MIqi+ssk6IV5UwdGFW4wqCpK2/HjloQhRPmPh5O48S5KFRjh7TMf0/ZKccf4QTC8Jo
hybezN6HqtYxDaPdIWwEv6d95VJEgpk8kdT90SAgxRYqvEUPkeC5fWMqxv3HTbWDz2ZxY4dL/Fx6
mddB6wiTyHUkzEmdSDp5xHKt9s/IxituxAfEVZA+uGarFQ/1u+VoDCfxyuosx1IsWz68ucl4BAzg
0yiVkpCET8/K1W6Odx1VE4UM1JI4KrhDMNCUHAvSBc1z4VjCqkGDL79r+s/QU+oS7tau1gjWULiy
Mrl6NC9aYltu4uCoecSznyt8PfsSVFjg7Za3HVL3K7L2AfalKvv+gNPI7f1W2tEoeRnpc2ydkU9e
ayAJl8O/4pFmBG0DfUnTnMVUXyj+JwoWAJLOeoqB0a8f0UmNZ9rPMrviSd9odFD2+gKIKgpBv9wa
PTEEhRXehT6x2kl7OrNRS+Qjf128VKVtqpgbdUzEogXRjAemkJ0YM6P2597Y/4Wyg4K0D3YuzdAQ
c6GurA+4mGK5kMp9Kg+i33kT0erm777WQ1pdLxo90N2fCPWFRYcNB2KM6kB65HQZGjv0XXD4rqnd
Ei013UTS3WopnjQYr1bGMqaPf2cEUKwSOr4nkClFog6Wg9WQxw5a6ozplsVNlZk21d8J1Rg2ioPT
DxsEDTUhEwvo9P+lunpge6T7DvcJVa6Ou9bG4kY+GUuPDl+v21dTEmq2lGvWLlMazQRn06v0GNP7
Q3mMR+NiBDMjnzUqZLwlwbm81O/UmSh+w3JnPzxgQzXyPWbIL7pcPJ7ZLg8ftCn443Ed0NsQCyIS
Y/o9+f1b1Pbkx7mxFYhKSzh+okrqecmz7KAGhi0VQT6jk0HHLyNz+eVYY7Ji8wT16EvTC0OCWvwE
/26b8finteBRAJY3cSlVZISvnzpB1FEE3xKHOn9Q92emyNoZonQpfWvW/eUV5t5C+cjcGPi+N1kv
UcWix6r07NYPrbPvt78jFogJCBP1wLe5oNttmEj9d5TU+RBtDZtt+s2nFjov24V/R1ln9CL1bm6/
BSgIOCvxRwZNMUjJYs2nJ4exvgymwjHIFmV1/KOjvlLg1Xzo3UKCPjcBrA9EDL5eu2DxvLcmtsGK
ViyFr6H+cIXjtWPihVZf8ESAvHvNMUAgtS4aOKArm+wB3R2Ux+6myXUV6KK4tpsZbKWAehplg6pl
xzIBmB0nu1rCXGu9OOwGgWMJUtp29i4BzPAks47CuD0bDewM+vp8kCiXKNlfj7dRmI6yBmNcS11A
Lx5Zax33UDyFzWAPdpOQsxMX8dOZRFT81ldUypF/uiE+uUjOmYOXPE86VeTe6/g32qhowGPXf5Px
4UuQLgo4gFTLU6duV8CxMutigF3fl/XrZLfSnNc87HsDRIDkoOUsa7oJN8BGiPAGO2rLC0U3bsgT
ZAct44ieHQcfeEYmnQgEoVE1eGCGmMLSdFfAb4qqpoUq8R1HyBepb9N1pHd9EFwSZABRoZm1nV1d
2Mu2Fy7jPRGtU++T9Ycvd1Bnji+WTVHW3x5L2/aEKXxd/HioYfsZPeDOkKVmQh6YS+K0E8DH85bK
qFasku/wksNr7v1uxIodPqL+y2tF4Ac4VPIMjG3BLmzd4aMhxzNRecaUYRIokhGraeiVm1IZKDPm
xD5/EbTkdt2YDRLfbI6LEYOo8nF0w53n3Zn/VX8N375upxUnuKw8P4XhrCUOetHu09JLJ1wKdaWW
4nHfKUVSS2jN24OsOpflBmUowLNWr6MmPdMHL3MSMzDGqAPneE66ReAodXc8g3OaRmRQkMhQY70q
u5XCQS6UaDr2BA11b8Hkiq5VSvMpGd3jRnAicZGhc4jcjOKd7OlVaB3Mz8KJ1WisOLngGFb53TTz
7KrlZnL0yqp1lRGeROSzyCVns02uFW1twzhyi0WjU9Z1k1BpkN0iPYRY/uLh961JgQm5VOgaPmL/
/Ft9PaL974PbpnEN+pe8MHybfCZJvqKPaNm2fussK43z7OwqMusAzRXEO+PSPN1qMA1+kq6x8NW4
/03DaM5hBqrWuyxeUrOk4vcIlS6geRUXIIqJhRj6oRs2Z39gBo7Kt+IIelxcZ64TU3mYSeGZJXYp
8/wWgZv1Yy9wLnfMvCY5suP/1r87u7IDZTDERu6e4KVOg0M1P9RGHfLtfgzYS3hGOFkXlHyTCP/r
J5UtpLP09vbC9U921Nlzf7yyO5BlQMEX3fsNrsNbBOwQ1x611MRKzoIJUBXtD9jCCiEDF/vV0pby
7aCyvFsEo54j4JWcmdEHcbGTvJTqe9r/SM88sgO6ANkJEJGNob0RsJ1WDyznYr5VoDP7n32uji6t
gaP2Ko/M2QdpQX3cEVzqxGEGly7yCDsD9VEeP7vLiVug0kytYJ3KJScqE0DnHDrw8tc/hxZB55/Q
7WiNgP9n/jZbr99GsB3UDqwk/8z+yDQlpALFjWDy1wIHaj8VCabmOYQ/JARKFBeNEn63PXKnX0qP
86ioDJgeYM2gQ22RSLdKadbJiVIS/xUr6PAQZ4xD3xeUgIK2YAMoKm01nihMJzRGOy4D3nwLC71c
qv16Q3KLwAsO7eg1r5/Q+tWgKpFq95uIqfjKhZg5vccNr31+eUM4jwiYA9OOIlFIFQej+uyGRqz8
dY2J7pdEYBTQA+NQwwPIOHsW/5ca8B3IqPuPe82/aufPgAYkNX7GMCYmTTCDCnp9tzc5ryANPfGS
mCmyhFYRgyq3WPhcaU627LoRRSf59Ty6XmAMMPy9XfLzTl5fpZghbkASbBnKXCpqf5/bCEXlJOqO
NzTWT5SFiJ2ApHgyVbzZU5xXoxa/Sau3CSXKWhxWCIiAvih156FrIqHKKVKcn/BJn99c5jh8XcEF
KBgcLm/1ZqRH0pKONv/H6zOMr50+5pU/qzwlZA9okFIIu1C/okc4Q/oYf1JiNvzGTXw7jv2sC2U9
4EKmnvemTuptLCkfwek/yf7aRiLakq0FPMnI4j4HARNf/8urMgPuMgZ71Bjq4oVpGLwbwEFk4FyK
VuEQ/6iWQp9SmV3lg+yfrjgeBNnUTiiVtfUCh0fBZ7BEkkYAaIyuwZ66/beCZdrsNZ946YMcjDZQ
gcTVIQXfcgXs3qOA/QaAhrz7VqWZTq9itHvsTowpD2IS/55wLjAmJduQ+lx9arqYUXAvvIClgSc5
bHi5gQK1I1gtOqbpppuUV7PjVhUDT0sS3t/eUonmJM5No8KHOOWEfjuBmjBRpVoDWuo9eB3AlfPC
UDyuM6ADKiYOKClc/FSPNlgmlSmxX+Xaj7Aj59hLpz7hhC0NFbRO68/8oK2hkGkBJKNOPDAi42t2
UGgqoLuOSmeeJ/fl90M0/8VWQaE4fBQNFbSda7v4rkwSjpx4mE3ALg6/Nf2yFxE59/treiLJlBne
UeGHMyUgnhta2ctH2uvChavM/xBp5tIPelSyOzQYzDjFu9kCzGt6W9yvMm8H8FXERWoCiabP5rah
rGvqrz/VkIqAM7IOavcvVD7cnycN37Ipapaup27wv2BwKszg6h5vr8OitjmFzsk5MlZTnF0FawiU
JRTdz8gc9laDX1KKCOaxeDMQm1vu0qh2XzN8fLTV0/ZQG78P3/ii5qqZWVPwMvtX/ZC+mV9QQI3F
6Q6UJL0+rJF3Bq1sPKflIMJLkwYJqPq+kO+zwAnWecmL1JuDbf9jRTq6A/rSsAsjmO8fhhhzHyGH
/tZHMHSpnbFxHLnSk+3tEjT374re+QvCkDWFCrHngZQZQAN2Wf2ZGvc6RbA1ajs+XRrldLtARkRu
xAYICPqLVCbRolu0+IFWg2tvKYgmu6XZ0tg+LYmFBXBtxBWvn2tCgQz1ddyYfmHfbcAEuiQW6m4k
4Vh8/MU2z5wInVewaGe//5yhHn3lWtXm77NxYHWLgPoPbZftI3tK73HXkYJmOOcR1QG8kdN/w5dJ
ZE415rSw4aaiUE69ZY79kvzZG5l8w2IY7kIJvwyPGGOXDzeDZGwl4BqJEgzIAIMfEoCr7VNJqppD
ZIWiXtOI8CU7aLNCOB/A3VQMYmsYcZwLA0V4gloTTTlDjEPozrn8bOkErogvqSk2TCjpvx1EJNFZ
GbJ1MLnfAY2cKl7X4doOPsIn3jjFBc1BNDhMI/Tg8HTJFPvu72x/KsMbCtUqmVtPWwmRciCEDhuK
o4jrQpTUoFElQS76k9J5foqXhfhuOlXk8Rkb9SN/Q7ASN83FTfBDn2NGaDcZmflzDfCzHYxuzJWr
5lDkrTUlTX/ijVDTNNnAV6UkcDF8JXSrZQCBSb2FH4bBgxfn1BcMQQNXzh03TDxY90ULyTtBnQZJ
vPoTsgBJ4F+VTrGrrPlenbWEB0J8Jwded3ZDUjw/c/l29vjx+TVBDTcwj/kaX99JJ+cP7z9f3AQf
uide/27otDrOPVEzOqUgFpb8BPDmWf35mqs5AKf6eYi/XP9LkpQ6YjDkZa2kDA/ybdxOG7X0NZxH
apzBhSqaX5NCm36hgUSrCZWmTISkJ9xM4xjEuVmSpai1C7VzH0TiQ66EfoNEyEeYT+iiLPwOyHKM
pV6uYkrSb1GaRuFOJkzgwkdLYXLvIkoq+MFsfMIg1SQgj0XP3+NWqdOEsObwMfVaPvXhy6sMK0tg
Z+glBCEA6cpsLF/Tm8qXKr+ZyIkzbJxJGEjgbdn96kBTW2O/an+Pz9R3fM1e5+4Bq4pVB6ArDhVe
Lew6xH1PsSrJfyqA6OMY990qGd+alMNusvpVnHd/O+Y9jF3abZX1dWyXCKGHxk2bu1Zie1qRoQvc
RN3jGkSNX1X/ph3atiNJ1ItkTX3P/Toi+aaEPRABukz5nIH6+gkXE2InMhScC/4kRVr8JT6/qZvj
WM3DeZQ8ZSpWucSirDSDAL7BHFrSNaIe1zhFlNom6JmNLfmLXxpOxwnIEZmfEYZ0Jg//nhArssVH
lv6sqd5M/I3ctZY6lvXtjKlrY/7zwLKQR9+Q3ke4wYQMmh2NJE7NKQ8Ua9t4sMNOFXSbAzg42wNB
Zua9ZxCoQtOYfOL54svdM78uovGFXdHWQ5aR0f2nXyRMU7p6AyqmlBHgxbk+tLrxtl/zc4mvauyw
TNqgd6Gfyw2O2yIjyXSQGTpbzh/oXKX4f6LfEYV7ndtp0MPbjgKg5Htsv1rCcEL8vucBzIxl4uy1
YRS1+h0JgTnv3LjXT3lQn9YKK9223e+cEvkLCSVt5X9Fl9P2opVcAQwXXlenY/5DjmiqlosO1/5j
jUWGp0Yod8fv/gvFCeNjH5YhnWEYWLysYY4OAmScuyYR6gAeHlS8F7hYzo1v1F0cHrStsAcjKrEk
lxTPy+CAB+65TvrwzqR1o7TLDy//YO/fjBjPlqtEU+F8jOgZcphkJHuoaZ2RTJ4i5G6ltDmNFvOD
BPss98eZ/PYY2TWSCE3NJ/rBLEktQspqb5Y0YYPS9JAF69m5SagRiLEi64nGxOhUYhvn9w+r+7Gr
0IT6Vww26D7kCQHrcqXY1L88Qq/BE5WUd4kW9mavpsTLPONZEOcGSJdRa2eXCsIj4t/5MTx+IxSE
49I12ydAx5/JOl0r/Xxbocej5caUKCAKgm9CIG49FGz/Ak71x3f7moVxAMBSRg9w+ZyOlKthJNvB
ZxQdMlIP+L4CD9uJ+cISZvuuQ3R1hw6T9L8M5JGPwnFweZMMklk6HJALA2eJ+XU+pW37amWXSuOM
gBlTvoGvPawiPNjLV8Y5PQsb2cJ0ipgenDglAkqRM83seGn0PNx53H9J20m4/0cG+EHiK91uxXir
4fPJwArNsyXBZIlfMHU4Vn7mc7tB83z4fgz3DtHiniOy1/XeFyhkP6Uh1po2RAiMPVdAp6xNo1iC
gEcNX5W+D8MLXfpwmbLjw53tXh4UlQfvrSa/LcAtlhgxW8kAWsa5hwmAoqxBCH1VT4lTrf/1hBxt
ncgAVXQknIcgsfyM/HgmoWcxk4Y3E+b682AMZT/zINyRkgdFxUZUCN7Y/pMrY62s4aDG78UctZo0
SAE13rbq+TdyvLx+pFCA2BprXbQeqdgBawYT6iv2Wpo5ZdzYmx+lnBkyOaj6LenbZUK6mffkzeda
WBEzX/V7V7u2FUHWt9N9OaS3UDlt1Rewwnsg/KU6z3zDmLthHxD5Jq3Q7aE9qBiyleUQiWS5xVIL
idgZso6yzgxqa1nZRCzhwN5ajpHbQWBT+CLxyfYg9pAr0Mz025UOtiSgFvncBL5qjUaPztu795yb
q2NRQ+DKnXUTWLZkCKMbsLd3CJKZNXFQo9xLwmMkyNHeNvHktgr53kWLsDSpv/hqZvLqa3rH7CHs
JGVrWTODIL+MLZ/8wiAOzpnJGmbigJ+SlQjfvunSvByAVAVp5Girt+lZ8osb4y3WdmqDJkhEuAz5
TWwON7hbayxftxn3byPqjHayRznXYfs5q/NvD5aOlOtoWQefqvDpTKuFmFkDlCKC+vfWKDqpZyh6
OiA3VEjQxyrEz4BYLpHhnhd/o0hwCxJYlfR/nB5z6dSzMc3rjrw8yWspH7+F3cgWaoCgPiTnxWI1
dz8V/SYSeL17hQBlozOkmSUCnJAxnqw1LzUy4SQ5TZPg8NbQVGZYqzA6x/ch2kzvKl5gWefQsFmm
m5Bxt1aY96XDL6TJepzk/qUDTD2FupLskkTEks5pqPJvGv50AwTyJp756R2NMN0+nfTdEP4MGaHa
EDxsVJ24Rd1txPcpJYf9WcXWTqYIuGUzWZS13r8QnbY26xRVONO2R1nKHOIFiEXBUShN0uzeBlCs
jxJDVLDX3O48mDs+/rjYk6h0/Eug9sII9scrdeVybeOOsQGmvcoYYFASRwKO8xCzh+FvnWYcM86o
mO60eSOqqOiGVnJ/Xf+Ixzm//yhxusQQnG7zxLPQPwvHP3+rEuXpFNDeBdHxdsQa49vF9kW8pHwL
7IF7D/Ycxw0lWVONDnNXbICBJK5rwCJkBQlFNvAjNn3Tlbg+9If5ucx4c4ri9CdOfV1rYZDtLX8/
82d0nuTmOLAuMRzvjCAj1zQQMuQCnlnjoeBdBHVvvRrqgK6URQa23IW2QUVk7k1zapx9wFrW9Yt7
5MuEqQJcAwOzXRiw+Jrl3A2gj9mx3tJNmVaFAvivwnAHhfW27TQD+n+1Z2di0E1yjxg8vs9rww93
tYM8dbonG9RICyUp6pd3GqMCxBLDHB9fosrS0QGnpdI4awpMz8SxNi1df+Qfs4s+PZFAiYHWkkXh
tc8jOSMmPmp3P4iPNVUyZjWkhflD/6ittTYTwPbBVf46WycQ0DBouNVL4PJ6vYwPp8cVbMnb/MHs
g1RbBPeZs30iZqJeafBYVqCFrYsD3Cf9OFRvu21LJ3J10RGZjQXb+TvOmjv9x67tG78RsNVOKWTN
mda6t9+iVpMA7M8005SD3c6OZNkHulHqPHFMCuXT4eo7GjD6ZPmSA9Ksu4GRNYmF+QY/8aXg9cxC
E7oDgGZOP2aJexzo8KRhns7V2x4EYtKRBMH/+mngQoV7tzlM5+iSZO0NaxPzT9iLPHexbPynwJkc
mxlkVYhqcCJFxoxAMAwCmGX9+JKO43AXHZKDPpNw8DO/wgR2c+JEkmuZyRm6pGPCXidifhPQHyBw
vVrEd+GTNfZbCQc4y1/HcdEdqtcV6SuYLY1hJZYZmgE1ekc7dfuzkEypytqM4me6XqTnSnXQWz+m
VPKazOiBo4oq2v9pQSgAVQWlyevXIRsLKVGKNBcqbY6CMva3pDnxkzyG4lEB7MUIH2gmFXQQgsgI
uagd8tVCc1JOypsRuSU8zsw/NucIT9Un6a/0Jz5Ox6QQ3og32Z25xB/eiefcEA/zr+Ptc1YcoiQy
0koL/sa+pz3CmW/nVPWAs1pBiyjxUhJuk0Tthuyg4OZbyCI7wQ74AQ9xleOWbSxo/UxrDQU7l3Uv
43G4OHo1YTsRJO6+8QVMShvsLs9pXHsH9+XGgBXydqMzaeYnVhDB/GUmqSs9ul8gGyEgjQRMDSg6
otzZZoYUPRCh1sDJ31NFDcZ6ZogzroCxLkZiyrqyN3C79hI2L71kCIlOJPGXjXU/E0MP9u6/Qtuj
3zrX68cV1LQ6cx5FILqvyIf7tjbwTPiKPEmYa4OqaACLgXjb0mt9x3nmp/eHonz91lG8V+P539A/
bvn6ZZvPluiwfFU2TRVzMNQX9+dSpN/E922Fsc/xq4t9LNoMfKFBn7VaqZchwb+fU98mBhOeQvZB
FdlGD1Qj/BHkDoNrFEFejBxiv3CxdJ58V+x6PnfoxIfGZ3zb4HId44lLQMFQkEb1zFBR8ypIg9+h
G/hFOztbc7FX/Pgldl76PggO1cEP+fjupd32HDsDMdfB/7dwKw93+eipeUQYNR2nHI0M4Qz36Glq
Jc3bSUcDGQj/bl5eCRh2NAUq8kHbG7ify7Zc69Ji3Y+H6PN5Uwmk+26equDy4814J8fK9dqW80DS
LdiMR5jsmwwBFObnLvVPz0Tex9pXw4OTL2UGnlwyBN2N3me1kbWDWyBLVUf5g4lTh+TESl2CufcQ
F1PJEzAuq8BpgF3gb5TAnr9IqsT/nq3Stb79BieTw4rNbJxT4Yh48/mxMagzeDWdcP6D2IqppnO+
B6+jgKhRuPNX9fdYdCOyJhXqs+9iJI9QNnWVFO6zrEYHDEcaf6nZo5pMwL4FZnVslxSuSFkcaL38
v0xAczMzxmqtycTlf1K9diPQMsYC9TJC0aCdEZ/kHyzCGq19BvPZEpksgL66QW/YI78XWBwJF+EF
yO/SW6mXJo4UlMSVqKvTysSBa+hzzMlu2mrME5Fc086rGtX5EK/4J6LV8tU+vQFzcPJBi6kFeaVY
IUQbGjReE3x41n5q3dpKXNybEVelF8CimLpcPw+dGFnGqJSJhPRasT1apA9nEkRfKIVpsMsnP7OG
5whZCBKUaQ91C+YKRZqc4QeCX7aVd1XgjeVnrnzVm5zp95mYyXn/IYkl8l48+VseNHGqlEZ3N5yw
JpobdsVT/JOqoekfA2Td/qtu2vATS7+npQr0HEBx3U8gPqDN8SkNKtB5Z9/DEh/LH2yZeoNVhchf
p3kugJR61Mze96txbx5QbmtoIUsOdCMJpv1J4oPkHKnLqyYvzTPmvaVl7zO6RnmJfH51KXNRPx0d
tOxGeB2RjoQVx3FLyVFbzPdZuZYLMRYB148PewbrKA4aiB8arCYIfMYw6hpoQt37trZ7F8zFEirS
7WYpsN0hWjwaD2urx1bsBerBs49ZcopBnJbgFpNn+G8+E97z/hh+yLoL4xsJL/+k+e7+2v7lJGrp
x+VXzROABbP2TzgwKjfaeul1oLjcsC7Z5mi42FtfrBxx2pm/KauytBaNN1IRvDJzrlXdYUu3m5vb
wy7jQBZnG5ALTEbc9It6fJntqnDfWfj6cvZYqTq0Lfk4LP9+pYw9O9KYJHnKBvuukJPdm+1qKOMP
/FmJsiQvacGwPdYNUSzIiCh8sB5JjsGXSw56zDg/pRTLpFCDtYrwBgDRuUJHA7TD+JicTLl7FE3H
I9ABN1hSHYDaB1XL3ASO+lU2TOdyWKnN+t+/h9qNO3ku93T4c27T4u7cLZ4Xo6MumiHOavamULOa
fRDODBDmrnv0HSFQXIzfD6Vy5+H9ubcJXJ/g2w33losn2sj4OsVRHFwBTmOKQZ/SPrVKB15ZHl3A
7tvib/gl7mBaJt8Z8slDg8icRgs61TQ/598xyIfbjHG9tOiDof6jTiXx/tZk0QoiwlDh4ZK+/MxB
uW9Yfcsu9M0RBqG5nlLobsNix/ZgUpLRn9u5xfRiXJYdq26pErcPKf2boAJfbAfKe/5q9NXqqM84
SAjX3CFcePmxQRcz4HDL4mzH4btGyIxRmuUxppX86hdCwyrRC4mCNZUji15htq1t7bhfe6RwdXlK
3DQe3hssH9B1A0Izf3RblRWhHlYlFZZPADDSWNkCxZyNntT9natxWuLnUneUR19nOYXzchwylYUF
eqkBFtvZfgeFfReen769PEg7BGZ1KS6GBUdleXDPOYuPim1AFNcNZrcNvVB/BLFPYhkX/sdtBiOQ
Um4uaTYbscmS37YY6Ucb3dWvUlCQ6r1kqqSGA2XJn2cAkX4BbCGf/G6FwJqR8cm4iez1J+OUcRIn
eGj5cQWmBv5hzUlcZtM4CIwwaIY7BFyo3P1TnofUlCVIm1WOEGPSA/A0xZm9fFTbCilnaMbAeOyp
abf+fC8+YQOvhldRnqQ93b1JkKa3QHWiR/HzhJkXZJM77ZRbPK5Y8+nMb83yxFNU/AAZ47AE3Kfx
pLae7oluDlyaEn9nasy7/wjEGnT0chj6Nnj3MBMKe26f1iiQ6X8XlTlq7pOTDPvwyTcgcMKjXSCu
VPlyp5sv5iwuelPSbi1unoFyv0GIuzxFkiL0L0PxDs41n4JKkGvNZN/sEIgjpwAB30YwC54IkQmn
aoO3+qWFUVUtFDr8dF0rw6opLXAbqr5S4/ItPS8eEN/Wg9auSxTKTIur5xxE2QsYZmkdmVWNsHpe
Tl7KQgi4YFmFEi/JX6qaGeJ8Ij3qDC5H5rWEVoeEa0FjGzEXZxnBO2kBUagd8Riz5n8x6ZR3K9tW
xRASIR4rOlEjG5smHZB3CbLEGhH/ICp2ZIYPnQrNa5tDkuUhcJTPb97cQbEryr+Hnwwe8x0CD3ao
o2I/wSWA0OKPMx6KofqL4Q56V/RrL+rvkUhrdnGHmdROMVP8fK9mv0KVFq4Hui0UmZeKpKQquMUK
LaAgZe8bxwO+QghIP9uhDNlZaBmtZEaJ+QdWb8FpnRehbjeMc5TS6OWqX+XYl/XNIzzd5oaPHllX
9loX59k8tRUMffeHCFoeL0hVJMRCoFsKkmbyDby7pS5bSyGqT8r7NiLtJaeRxf+IexxSDWD3UN5R
aFpQa8GNDLdzSw8PsR5Xp017mrJ6IEnN0hLEFL/mCgR7l8Qir4sxTD1BJNqbhD1fmRkTYpQlVQZe
/3CbsuQwbMxHpRZ1RhuHAQRqAl0kZT1wXdJD49+rKggi/j1CaBLYOAWpV2EVu8Bp0pw7+oAgjbuK
RkwYXBFuqTVWz1j0OCm6/E9RVSoB23ilAZstqkhQAEHxz3vetB8XRbeJhN1V7/au8z6xW+HAbFqQ
d6xZiC1fbvaAC0aXc5cuEVjk3llg9UDdDLaHgdT8e0v0juVOowxFt7+WNgSQxcX0YNXSiW/FrxcZ
PrrqLeA1CHYuAI+5bewOxMg6hGXTjKKrp1BJszkE9gpsFVHEoRcaOe42lVDUvjxv68l8jFBp9+Nn
p76SuG5ae2+SfPiqViGMYOWtg+btcMevDW0eo8zZZGxsePJdGsiuO41Md7IFOfhRTTT4YxpvyipF
DSwi0iq53ck1/+m7c0w/2x9wSHnnDalHHqPbkyAAr1fCTegfUX6md53zWfhCtOZG+eAD+LanFVn6
z/86T/8wBQm+ysfYbxdZ3KGxBsYOiI4cuv/VZ/hKm46hTjnvy+9JQz/A9Kgsjj7h4KQ577oWuzRY
fkt1enNrvujGw4XCYfozKHvqAcWBxTQGSehd0cbRNVaghIrg7/PAKzZYnBsAVxXGabSsA7r6szxJ
/xHG/9P2RsN2ys+pC8OvdcuqK/mSjY1B0LkHBKJD25O+xE3TGrwEsyI/e9d7FzF7m0Huo++HadXy
VIk5Qc2lgCKu17GUx67+ge6Wd23Nxs6hSgAMcnxmD4xoq/VYrsL4pjZJF7fAcopJQzRo2yrTV2qV
UAVhdu7LWoH5np7eJnuxyHBJhuLAMSPyGupK4HeZVcupWXUjMKDPc/nQcBnyvc3QMNFkQ+/fzbfx
yXJ0MixHFaC/lmzm5VMHpn/Yvd1MegxIYAYXsLgOYlrnJn0Jd8c/kNHOP4lAaZ2gaWa8sf09pWp2
weQ4hO/X1pq5pRJfD7Kk+KjL/0SYJjb0yvp4EIMcWGdLc6koPqrfgOmJDunxkurDky80N81B3X04
WygXg+oLKY9WjIHGdO/W4/qkwLO8xbO6OhSKxksIP6WT6YMRM831NwDn30mT4iKHo+DFG8GOMliD
DA43PlKwaUAXh2QyfQJYqta0nSiE0n/JTKz2Idnzp8SBWugqCWkaz7DjrA0yF/xgM7rOdXLacYAh
fSFW4TTET5eUNtMAlz+eAxx8wWTbNux1OiJqOGhtJERqsdamxbPzJNB7ycF0MIBvdC2Bj65yOVof
pbc5mHQr4dWAV/DzATawTzbeOs72oHAJOBa7jl6jaK8cbp+YwZ6Sm3OCeSV08DaSm7rMZetmk0Gj
1oump5E2KAJT7puLOzJ3ZMQ2oPYY1ElErf0swvhZ2o4KfM2Un/wR1toZK2pakReREJFWhl7QaxCi
Wvk7JIxKdRaJoHudIRHSJ/WK1sGUx10OXCOJe0mvOt2wTcc9pD3ilPQuORoAarIuu6BDAc0jpdHs
Pj/a47FI69M3bwAE/ckhYBR3TpUe4Jl1s8qhAOKvi7cjrndSfkwmowiUmpYsftiTOn6kevWa/hwA
umfKNVapfv1Q4SwKuJBsJqdE7xuLXN+bSxhuPivknwZmHCXovA03YKNl8KDWvO8wp14tIyMi8x/V
HV4dzFG02ofQRxAMzudcuVEo5I3OIT5jt9Sf53zDt5DF2gm9k75Wei2FbL46xCrpRJ+UC1vH618V
Ccmsm9vLRJclNqvYC900zr5VT+XbuYyNSAumoLJvlMUJrhbqoLsccxBQ6C9p8SXIRaOC0UJZ6rN8
zODhJCDZJUlmCp2e4dW3LE9djEfV839Emzpaghc6XkMsQYbIjYxsv9yChtGspYf3+nkYOPRMyhke
9sxSRpMFXdmfTJSVuKCyg4ASP3te60mTioKmjS+ZdCUtc43+bZNAXlOPbPG/P5j5EIOC0DQMlkZp
ADofel0IY0GPc/aa5ys6kjEoC5wLKj2hNA67ZGKQ4Aa8K7ctMOtvLb1mYlT0QuCFnRyhntnWRZiA
3aoFB7QBtn40Mlx50vsLDT2P0L2QC3S19r8cfZuaY1j6q21pvXWgBUTamUWXGyr+M0SIKMd8jfhp
YF43eEwQDwCYbEOQHGWMcsmHU5Uaea9cKefLAYMHMRYC+39zwllWL6B7/KZDlcptCMqv59BFjop7
hb3Z2AdSszsU8fVt2PraMdSCu8vyaMoil3EVA4qWtcOrmqws2zeGPg0EF+GK/aa6TCLQaL7Zbviy
u2QtS6tOJUpke8mViH42wHikH3g+aob6VZhT40Cccgy8QwKnmd9NJFd5ykvTOCmwhO87NymfB76c
WeWwEnbQvNN8yxWCBJh9C04MwErWU99DLaNtGiOTOgbUWMqnS5YrIDXhmTkO1SXO3g0vWcQWUXHR
WEQ8Lst5cT91hEUV8mdROxBRwFya3QNY6bFL4/k4BtbNssvvOeNFy41FWi+DY6GV0OxfqvfJ8ln0
P4mv4Lg6j7qdvkAG2H4kuATGU2Nlp+egpDJwbZiRpSUejhD3OLVdjQr1V34VQbuEQaY9bhPojDMP
wtMnHvOvrIQwlP6qFXLKK1X0WotY6iv5wgJvcYZqqvNveAFv47Ikg8o1CHolbfRI2tqhR0LHjSx6
JnXgbz2d1yWZa8/GriKS+ojRZH9LaqGqJlh/EHS1DROyg0ELzV7LOzc3calF+7WoA6aujtanK39D
RW6g2Uov0VDQb8LS6v6iHQaI+UG6vKN0ViLhO68fhi0cxp5Xwq2zbhQrn7BQvR8DQMU5+3AWXVdY
mYU7IjOtdnIsTnDO64Rp9EF+iwI1KXGJL3m404UdaW+YtIDPuO21IXVSLuPwM2o4f+Uc/4WrAXLW
OjsNoedk9VdQhgrhbwDdLQ3b/8cz5uAgFWYAvN784e1wkkLLYdsb5u2y5WdTQCkV6K545tgkHUc7
pGnEMPeGXfIGLg6D0akGiD+f0FULm8+D1L1MQaVypMq5hUA9F3p1TaBebUuMzotbyKZnpDBTPzRz
jCaTESZsA2CvMyTqUaIMuvOs/FQzN+B5h9IUHqQzmEVjUlkxCZWgMNOP7dE5Vse0vfs3n2pc9MUe
KxRQuIz1C49uG/0x2wQkQDE51wHVnnOm2c4YNLYAizisbxYnxRggg+HO0T8TqNX9n0/4OqNy8SEZ
JSnV7caSvY1mxYntjmiSJMovxLabIPKwmAKWgZlKbJENNcQRIdr6SdRZ5Cx6nPqI5h6o03YcSGjr
OCyN0JKqO0a4IRU2UpkqTfWEwIzk9+xjENX8cDatpk5IxadVTTkSMzj4b+pJq6jCEUsLAX828PBB
qIK5lA5SjgwNmHUsaY5ss27+Yq5rJ9XhArpc2vTYB7//LHE5NZXHouLUJ/Cv6e4ZkrDGf2WJVc7L
uC3LJkGF/cD2yQuITC90SkFiHwXYgJTAbsN+fykSLgYnWo8dgAWeb1FsARBgnoftEmuHnK0VJz1P
JdowxWfMmbzLUoI5O0QHTX2s4lX+JnsEDji5MV+z2FlcrfkBp4iGEJ6+dlc3KXOledR3GI3iloUE
WqM0KgGIxTPrIUD6/TjSrURxL/nRnovwEc4IsP+2YQ4yaWxptZO2riXpdytQaGkj4xB9QvM0/LUk
F5PAT3+T9ARi1CqjO/24ErVP92BkLlvGvOud/QMJmiFbNqKU2vf4d1SWg/ByHm3qyx8+4MYwsdj4
98zsAHFEctBlNqS/Iwi71x03/n3ymnxvW8fE9mTIe4wCPi3L7FQ7USDK3JtbJQTZBcu6iT1XwJIr
vynxKy8sCFkSTyyELUgynkPZUtaz2QcXQXVX6U7iUSoUfigsM8PP4nkhquOATeunPknYYRUy6eHe
4oO9RTkmC7mLXro0sougTJ6nTyupiT5lHzaNQEO+r1MEdgBqH2CjGVWknXL995fFXkhxikB/dwQA
q/0g0deO+D28bg0uD6ipCJbRPXEnmhXw/d91l4Osrd3QJt1VDmE6hTNLp+8O1CvGWiUXjWYDO/oU
rJXORWJ8RAZGcTYYXKHq3TrtLGazXqAFC5msuFbNligdHRIMPm/PoNN4Bo5mX+Jju7KdY5pYwdUs
POloJU9WK76D66MKX42uTPdJ1OR2QObL5UqHQ4PHx2bWGDR/pcAC87KJmzQWf4crHyg/d3wkwoeP
87HWONBNOObiALyC2tvVd+TBu8cePnaLBc7h6kJEPTAeYcMmFOuGb253jc3hM+tL/YmocE1lZJCS
b1ZMr50SXhrRjHjvkq5jy07APxaVMjFgUo17819G8VFR5yAHn03/jXpyg7EjSCjPO6QOUi6+wurp
oDLWQ3/m94XeVyifhtRFPl7ifYZKlmg1fE9WJEhMN0C8Jjs0zpMAEofWWlj9A1suSruv3Z9jh4ES
Lu7+rIuEdoow6v0bpW9RvcHKsd2Y7SNenIQD4XyssGI9KxIEXXxpRw4eVOyLwCCQOyYVFYd19T+Q
YXFWoF6z1WqHU/cAOw4jVi/8Lz65AY8R1Khyed50VRR6C8hVdscj5v4njSE5ewPfesVDV5uPY3qQ
Otx8nhi774LWXI+CnXxLIBloYBW7u++mqzWUQiI+h+Hz3PQyWCrmOCGcczyTwh6K6wN/TWk9E0E/
Ti25XNDZgk9fuk16eCQCXtq16Q6m55EtnDQA5T98P7shz1cjHrLUfaWVkIrAleN6nw83MeDNhAXO
Smhc5j2xvmLZnDbmmfNgzUH4fGuy/RjwYEeRYgETb1sMeD0pz5tsdiMegF+V/Sj06B+T7LEshS3K
2SxmKAfpyfhiSHqTRc4l6+IkskK0J2KOL+yh0EP901ZSAOutN9K1u/43rzUWdwFdXzivUwbvw4WA
7GgohzCyWs423iqlXZBCbTZ/xmOCFeh5UQbIyEeaFqE+L5lQMfNHCZngaPT7DzrOUPP0nseN67UV
xgPqz2MhnslJdrS1n65PYGNQ/SDa0WmWbkmosYumEi6jyPZTrHMQKF+b+JXM/Dy7/ftnllT1GXoc
Uy3AQyWSC27CyO8yVplxDzM8+ywHzAP7+wt13yytllCzdsIautubwZ0Hgr6eM+LHB3pXsBINQ+Mt
D86cczTk/EGYkbdsd7u5iX0qX+eNCAUQyANlMGzf8aU7JeISCRcCASlaSGsN+NnybVbfwbOmUI6I
225rpk6KMj+0muKhhFVnxvafX17eGjmUo3qCuIO875Pgz0Qp8rTtn3OfasrDs44bY92uluFHCbQJ
GMRjhE9SI3xjErf7hhQ5ZAu81pD/hPI6gx1oJV/N2m+WSJbbK/yg0ZziLE3fbiWA6nVJIQK051FV
5J8HzMQlhT4uYkw6H6yoVUyXgOH7KijFz0KSQp0u7pI8l6BEYpB7Nu9fDDyzPSBWfj2rzsB0ZeVR
menIrUZgG4/jOdLYBLO9Yd2Mv0lKajfUWwHmSWasad8IpNBbKrnIBFlN55vl0Tddlbr9RYB3jzMk
h/SKOoP5A5EURnu8RP42F9wXJrEbcLRCXyTfQfxWOOqRoBqOIhjC3qViWhpnXYgyQ2VsKo6s107O
pojVPSJBwbQ382O3yXNXVB9jd/c0s0PGQCjwLNsnk5SApeXYNQNJCWKy3IvQoDYgoFfcMj2kC5OL
iquB4ZOH2nliLi3sks8lYEqVx5RzSFBnamEPFAab8X33OGL2jF9MLduG2WZTHSJ5cYoKszuOOpd6
0Pkf5SIGHAkPoHWxm99VNpqf/33n6T8qzauLmDkd1jgbwmgkjU/zOjoZC2KDELaf4zTZK7/cD7S/
ufrmMqcaj3SyW9zp6sNTuHDuzIXuHQyQN6xzYa4aOFq2b/dqtDRkQ64J9F+XcNdaTuPj9yY0MUi6
YHHvCyUD6GDaYw6c9GoxgzKoXvLEluLm6RBjiSDbhGRUBSyMWdynTLGEkYNW9eXWfmBKvKuW0hGB
I8L++vtivKuVwH5DwxOszYRgEiJPTj0eDbS8hRopo5pXZbn4Z46cJsqq2VOIPNiRyq4+nIrmJnK8
s+88iEnLZaGrT4g7t/vVmDQQcxsq7YIgA1gyGn/V/ZTIQHR9GIlSIeaHgySxbj3ClceGK81aTrq5
4zkE8tQYj9hHzlP6/ZLG+zUkxt3zD1DY81QsMLkeuZeP9wFZiCAvDGK8n4EUDCzFj3MTUBnhCrhA
lC81XAI5wCGV4xfeEy9Tl9zzgHgQAzM45La9nsonUNBxVAvzLV5dIdrC7f39bdRdS8jZ8qEofMon
0Q90o84ifxV2RzLcQqaGr6FUyboXQyyiQu9QZEi4YTH7UZIooeSFJfKE3fIlamnMZ5h6MRSyWFDR
ZbSD3BntsT03rUk94ASXSaeqThCZ7309pveUy4ILXKNztp4KR/5bxUI2eoUkRoV7RgitF2IxUksn
qMQSutlHSXnMBck3mSrFE9kgZ/HGkdfd/Cbvwpqt5qFFcBBOUp31qccblZVtI7gXe4HlLvk8/2ya
Hb+YsxX+QGJJ5aACUMu+hSlOq1zOA75KxJ4AG0+jYcAgZblxbDi42sabYrWLhA+0GUlfNaaf0dL+
3p3pUwnBTH4NEn8jfRdItGNvU3nfodtATzlj46AbFflUzATz8alZ/+Ag6WSWJf6JtD9WgBgt5w0q
4s2biU8qeYuLNs8360C/q6J5HDREfug/RxiM1BRx+U8MEDgUZFwrYwxrnM354N0jlD1lqTLnSJg4
MPbtVibmTW44kTfoyZZT71tuz+HMeBc6sJVJYJig86sQnK2NUth3HKPBzuHEY6QZZTpGqkamzJ8i
S2d+h2hSl37Rsi/6HeEyGuoaBfe7r4MeuxrDcKMDmpJHXw5kCI/q37x/ZVpmIinm3I16sJCyWYG6
iZZABVP3IQiMIQkJ8QPA0IIKGrZgDICireEu3g/Q55r2d+qeE+wlOMQEF05SksUpodKvJxnTj05S
muu409AvVKDnKiDJc+vDqc5ZJHDompUZhdmMjKzxDDsrBoSXapr/NJMo63VyvWHAXsMxBdDnALIm
AYs/Lu3tUIpyAiZ37iGqZrpF6OyfFTDcZ9yMeeVGwJMihoTSX/XVoj9HJNQc0VzhxhchGiJiJdQ4
ZrICmlZVgCdsFF9PL0A8B+GhWmEAsRvz7CBk0KAkpLKM+L6o2E+hv/uHXWin/pSNsUbxOqkHnLt3
v4NYR6pNoroqgSDAISDKS6xrpenxF8A046eYZ2lWBd/KHS8VOUV2RsUISLbqwyJTYXUECRc7HAFJ
ZuLRJY8x8k0v4ooeo57Rer/3inwByWR4pjOSl42XpcIkpRkiivuk5WqtYGtJXiqtl92mZuRAzzTa
891yihIDLPWS0d7EgJ6CJW9r7HF3jR3hYPC57lIro+NuiSslrUfFXXSuai8mW5m6xW3Cn2I4p7mN
Rxv6HSM7PitEhUOTPxwLDMd/EUNkWdwD2yrnEm/d70gcASBkjFkTrMZaKKGLUaQNkXd1cPWDgZ9R
2U5ZFyXbYy41zLizw5tp9Syz/aBFRHhQCoNeZQ2POfNeGFaIiN0RkND+Oo1Y2Oj6psSSjGSU+Rvj
wZyo9k+a7wgZbqTl/tJWogGDdmPnQj1kAKu++ht7N1o6J+kGZxhVkvLWVO+soHhTxa4qrpdeAeHA
3QxGobGdRPHXXstQX8ETdUHgelRFveaVFAmGFjfzyZeQKlcuzkRFK0OodZeFjRKn8T1ElcfXqA3E
M7CJ9RHSSLbBexDS+AbGEAqKT1CSYS5INIbLODVTYbZSt599WvGGH6tfGGJAseVXfbNCBzx0dP/i
T/GONaiz9HZIXh6q/aRHEmATYdra7iDuas8Hu7PRqXj9KluMcHmE8gvVlmkv+6x2i4PUxteH/G3+
pXxUxHtsOb8aomz5dkB69nUPXpovj0pmt6rA2Y3+zT16z+WrUcEp0n/X6HsYw7wKShKG2cojjonU
rfB0jKu+F9zaC0XQzNOqPSFlobbsDIgjQILmv+Q2zIDkl0nMHO5J7S1PK73engUUhLQZWbv/NRJv
nspBMYCscNajqN/IJXyBhe3qlSxdlJoqpC18BZhv3XKVGuL2+VaWHnURmkGbWzmmQ7NirmaFbzfO
MZ6lLqmz55hkcg0PuZWBhCSuzgCXlMEm+XslncUzRW1toxF34H0+PS6TEMGDAeSl4/F4tge0y4wP
WwcHm/9EMmDUe92aZs5T3AJbDRTGvkcF3nw+EhP1B8N8AnWMpNkz3mTkS0FoFBBHK0oCxNDpPXar
N9OQsus6vJy9bOW32BYscwIW8DRH7LehwlbUoPusw40DIIttNHAIobob+mgrkVb9UhIjocvyZzlw
c7hljZjBC/WU0nKqQB6Vqeu2z1tQVOMDTehqcIZI03hOSC8JTedaF9nVj1Hcqfyyw9GRmcM4LJgV
ZoVsZ3V1SG+HAvscKoodtb6abLbrw6djp16Bm9N0cynhkbbrSJNwnzkNEvVWJtLDQ1AKdRPXFL5C
+bwlMqkxLyzqEv0x37GUWhBsEYMkIy+jO6h5BacBoP8ORxwTeoSrjfR/I0XOif7OnZ2kIv8yzeBf
CBhgFI5snKVGOOPuEZ9wDy0Hj1K13rT0YlyMlfWDDGh/Oy7ek+zei2wJtpnLEs9lzPYLqjnUXWVZ
j6yM8QoFWigPtzpQp+8oZFOQsCH+PKExiEhy6MCFjht4hcQjQ3dEBVbNW8nVL+R5EvRFcn9HVx5P
G4EP6KKaShQ8AivtDKQfe59d4xidxF7k4804xo6P2XARv4IeADvH5Fo0WAi+TWTtnVxGQe6f4Gd8
5nu/ubY38CdsgJq0FFUl6jK9Pmo8JoO6Hk+ZlixQfp5VSWJu/MGI20HScxUOh+pDFc9hx3ce7C3n
Idwa1HPjm+OuunGv7l3q24yJYoUcwq1cqojvQmdN161Cow/niQthgb+Cbneh9XlFg+yJHDqIU7bF
kN6piSbaJz6A56AzzVmtCoD9XuKQCf0mdHreudTWMWcRz1T04YofRKLquyanJlXlM89+cgNvXGTg
pz/uN6TjfHvh8KUioRpnsrDGmm3LFmBiCpY5nJQ6HxYCgmbw+Shh+1Z7Bem38WgPJXQStsBBh3ic
Gr4eTTzRNG2nKbpRWDiMntJc97scTY9a1qOMQ2jdGinWn3fN8kgFsqHqqcgVSB1fHuXF5XMYd96/
NwvhDjzgM2upQO1ZrJDbbi/H2Xb/J/1VKZq/jQQpfrGjnl7ugJoZjH0ksHTCsQ0Aq4f955bSZAjV
R5GWkFf/gvblOYic4RUbPFzeBn4BWtlV67EoO4c9LRyG9F6XM2urjW3i1qYxqUdf4NfnT+Y0n9Ey
+DKsWzPu3dC2P2UEE25za0f4aBjnkl7M7tuHqaf91r1KvKwDIk+PLdG39UG77o6kH31QE7sqp1tN
DtbSvLYsIERhMOz+UAc7czLMMSz7T6BnSro3nLKs4Z8dVgtgYPJxjVV0cL40qKcyzvQHjCZTt4Uv
IUTRyRqXn10066pgNjs/6A+YFPzXcsA8pRB0Ha9ehhdJ2/evl17sYEoyxCogEqUaL+aioybeMv3n
eadsdQ9gEo4scwzF0vlmZ8LTC7OjLauqcmkBq7vKuTx7iLOV3OfGfOwX4mDZzGgqH7ksWnLweW9z
dvvNvWRk4nfVveZzR7A18LD3dqI4/KJov/JcYv+VGzwZrT3ywuvmy1JKJk6rrrQDCX+oVDmM0lMD
sGYSZCQ35/NL8ewtyCHZ5nlpSf43avUIKMFUfLDIq1EyzvsL09r1uV1yPZKhta/UyWbjSy4PUEpI
eu5HCpSwgm96AUvjrrG8vD+SSlmWHcdeoAk1HpmpSPBz1efI7FhBcscxKQynnPvd4EsbGBDJKoZb
3+v3aAbrQUx6Qk/0E86HXsvespkwYhP+O4KH8VuuiN+QM4XSglbqaHKysXA4kuDBM8bKGysIQ6kH
zlqUyo9VZuncEZXS5nfunIgkzzlK0WNc+GvShx+dRThO/Wy4NJFfRhQ8uarxVVsbng1NzjU/Ne6u
rME4BupiJzvpyFgBnq6LvAfqTvsqCqIoOnEC2e6ppUilwuQHLNl4Vdu8EP5ojlG0mPqtCMOdGlL0
ttymaNl1mtA+TtFplHSUOFA7IP0Ug+hU8YuJctvZ9aAbclZwbPzIxzGQCkEYPQgSMCbu+KkPBzsR
CPgJHuiTTa0Wo9plNO0pBFxekEFntZOKVKkdzod0WPDP1yU6+YSaNt4RTwZ3I5JnQMu9C9koL3X/
qQv+/w2Qzg7SAXC1ivf3j6Zn4J7sOUUTt/R9Dnw/wXARVM6Y3AznPXZsWpZuLbTl87BtGJe4jNmN
v0u5XP6UL6BuX/eD5dGK+AI3L1mR9/INcA5GNfVmwtK3yljMN4FKiXMRtCIPjmIcPWfO7wymQBjA
z3KPVnJJ7wJzM2qLeugu4JehQlGcUdwASilqMoHCrGsqo2lOYY/OLY4O3c7j0mitlHsaEUqtRUVX
WwgFTh9PnAPK77XX06VWtobEuzcO9FUXnZ22XCpG8vG7V+hpwvHqmIT6xta06E/n42e/tLDXvurj
GEpOoRUTG/v7Ci4vro0bXllZBOLxQ0cQvsu16JZ6F907o0iaf8p/TgQo4q+mPjEWtSt8Mh1++qG8
1nkhhiDPgwHH/kra3GcrnPXYr3bCxQ5aNCKIZuCtgO7Q72cse6H9+Rie7uo6B/Yw7AmY7M8JT5Dg
LV+GX6pCvWJ5otAVuqm74pzue4avwEAt0ROL0BXtlLpBcvwujPNuRZ0FDZxCEa0hnJJ7X+7+qoxz
YdE9gfC9o+wtKKSInAiw1WPVe9dcOXN67u2lPO+qtQ9/m91Lyl1H8upAMr+hEoqSTkm3Ik5oWosO
36jetrQRSinNukilQ4UZXQ61TBOtCFiWD48f3LjmEiqyWVST5zZGxN8HVnh2A5yShy9jrlvJJ1+c
xM8uOU0kAJZ3xEdxs2iz+tAcDWSjuxrgTxE0UYbQ++g+yCc+OuCd6tkRW3fdq1Ryrd/V6yvrcHSk
TEsosE6OcLkmAQDKJkES5JcOZwmDkugD6ywtoYXrdnPaCSfnoOCRR/LAOY12KIOtq31QDsYMQKzy
Cg7IUDBcX2TvDZM69hlSsncCR3KTcURv/DG2M6FWO5MVhtXGwATdZ2lXeKxYYTbZFK+xjPpLgOpr
Oae3yKLZezFGNm/OCV+RIMGr859CcVQC+kczGjiDrBHxl+F8Coy2TLySBi35cyTXLaf90vx2ohrb
GW1Hu1UUOV1yGTa5FTQPYlZfSKVx2eHvNAOFlYMm8ButN5SC4+vriMfvtiX/yEPi+kNf/rw0xwXk
ObCZWE1CyRzDH48z1pn1gtZDzEseweW9rQz5uIemRB9ycVS2ymuJeEbp1j+WuAJHOJJj+p+S/3GA
iCCItj3t+bI9ckLtbNksquZIF9oYFPkVwuRQvrCsvHoesl/Cb8vyYIkd+oqxjj5TQg/GEIQNslOZ
VIdp4o/etWrUp0t8ONrd4ysnCrYGzoglr8NmcPg6kb8C2WUy9AqM6c+1k6pBovdVbAX9m6InkaFS
Tevqi9dwvvRxdqgGUvT5zdmvC4gavWhyF/kHhq5MwohwkTEIoZg5teHp6VWvEC0YXB6Uv8pF1o8Y
EmpQ/U95RHYGKfVuBUjQBDA3GJjMQN+/XRv0vonMIJ55kO2x5Q7of3QjRySGVfAnDXQ79glX/Ko1
FjScClvilx8ku6ZHlafNFjdLCsZxKlVZDug97DQRkliSl9lMphsaVBCBh4LXf5Ea872U8S23KBRG
t5YkCzHWSdnbfm7rslzMoFEcYkiF+JU7L39foUXJ2WFO25ptFVdNRUgo7NQG6BOPFXsckVVurDZ1
sIROvkUB/qE1WmkkyV+c0H9B8t3nCH88iFzHpnxfQ8AhLik/ueIpV8Zk7G0naZoSUaLJT5jTLOrW
CAi4T8mjuamVdUTzPd2CHyzQLlHONCdjeMs6TR0vtSgwj9HjHr0Rjr8mMdyHqa0uXpjQJIZ8NOsN
JVXxOvO/ob1GOcPsBtTS0xkg3qgRvDr5xF2CBdyMerOQrI8cnUqs0+/KmkpxM6vVbNtyapuak5V6
/JElmxveqIozhUy9eHeNmPRbzWZNVl0ILju1IgZkbdsEZID08b9jXeGM8tZU8J5R/NYR/KN3O+Hn
s48ujYlxV84mQxG88tlwZ4fAAxLMPpxr2RGnNoVjG3uNgxe6c1+FlEIiJ4jqgkZBawOl+y4yjifd
+ejTd/JYTTw99NKjL9PmQJhhFdWWD9N2Xa4Hj2SBd7mnuXWWU7jkin5shxst8zLJFgHVDoqEI+33
+e1ZufYBBbXNb4O/FDhNeR/PAVR37zaCRweEru19+cxrDqw3B6gBSSXof45YHwGfoPmRiVDQscIV
pHZ7euU5GRoFpIFvY+3yIpb4YiVtQdC2P16c9YrBXruccdwtEfyzoruwfTOFgRIk0hP5vjcrhXDp
sI8igQq/jJpewphDT3vhRaquRn/aKh6FSKJhS1cxjdeMeGmrnjBkenRO0jEwTUafoXJDT5d6tNfz
/W6WhWc3HnNeWqsgZSFsJcpdJdCdsPsJHXfrSkjT3Yx+UsQ1JuXjCQ6xpoxyZ0LoCrnszRLZ7kEF
KZ764z2uh+HP0vqrbWjxlNrHieUjijIIDNf3IW+9taSmraQV9Qudb/1nmm0Ffu5+LFCWesxvcGlo
iTEO2sapnZdzZK/zw39HWbRELrR1CSNePiXRljLmKWqeEjxPqr5p4979pwwNBGbBvJWn3+5+6pmi
KuZTc+2XuLoKrN9xb9WQ1gPdZ1/FtaTaMP3z91Mx86NeHwLmBD8S5C+qNB8haP81dtu2mepkUojY
fQQScM4VtLN/2mp+quyZZJsUAVcgFmeKBJA411bnnGCtlfls0zFIfh+/wbL/tsJl8/LroRgJ/sNB
gjB4G6P0RY6uOz7zj2G9XtVUoaGxvT66dzJNnOvSChcsQhOOQKfXxNBtW8ZtruyQFxr0/+kIf2gy
zdyCowp0UcYbqOO8zoTJyS3Iq0EWLeexWgKQXl4Ioge99MZ+vIxLPlHtCkmvvq4n4y5dHzj27TBM
Yi5HnCJnOg9cCcDvUQ2emxJEJeP3fSK2Vr/kezvmVlZo4buYxECoHnfBamssEpzCZ7HphZZ6ce3a
AR4DsFUwPXrL0fT9QuLpn8V+4kn/uk8dWSQegkqtdNnPs4JDOJwogETCwEsEu4LD3K0q0lnv9+nk
W3FqKQwgLvqNrbdxt5ztB0ArwDWuxfmI/DwNUp4E+/ztbkyQkfb309DD68ev1hkWpUDgQD/joQDt
pr29I6K9IDE9ExILEY9MLwgrHJDayNe/GhE5JubQOQj1hZBmXCoEY+cmdbfauqjhGhOYp/vysJpr
X3FDlhBK9p+QjSNYMvZNDTQB+WjJZGI4zLKBrmSsQt83jhY6EGlrgg1bCLYmBgAmhtSB6NZYFLUZ
FxhJdR3BnTgOi7SFgZ5OY1xWzDGZf0ySc86G3y/7fJmzZg7bHAQaO3s3zFpJv7SXWzbQfWwIeC6w
Sq3dsbZawrYy/JyAOdD3BumUigHcb/R58WwMv2+dbCCF7Y1Dorp/sHijxX2j/KCbZtjEjNkjeSOu
dUJ9Qh/ZEu1Xmrx23R2gBh106uGovpsuxfzVSB99I6A/0jCz0HwbgEz3ywQvVTYOreDYR3bD0ozl
IYC0McmnsFSfsiSGMQ0lqs52rzRWLqW4OkGxRRb/K0/DOqI5FlKEoYxgauPwOv3tjhhTiuQi2G2s
IrY41HTDxLydmdrv8wbDMogtjXQ43MB/vBz4ejX/FRuT3TTjMv5nb3+0o2OzXOvlJa2tgdH5PD4K
fwhwE23L806//CJfG0idt5Vx43J8/kZ5pP2s7l/bUN0iY7iNP5ozrB8LIrU4CR5iuqGuMJs75xaw
z0OS2zeXk9BxWhJNrPbqh0m7YzDUgOPQI6nkSHql/6kqzXqiUDi69IS1Fd4rrmZKi+L/xpXNakfF
ECBJqw2YROqrNMsoS9ysTI1iEwySJtgY9w4PQG68ubnESXWuEaw+hmX5ZtfXH1Ywqnnnb8VR1djq
r6v+rHLrMsVFLuAk6/FUyIFy8urmRFqX6A/SgQZ0XqZCRdDBweY9vzyeRYNgR/+v4B11x6LIhufc
nF3VjeCiLLDWY+lKKOvmDKc627/QLZ/om3CYSU5RpN1oCnsqIK8JohcDB44ubVcK9cG3JHn2zZsW
vfqdqWgjyrEdttaATpEKABHwnqulcggWs01v24Kc1ZgVFs9kStJYS09bhTb4E6LhkAuhn7k9CA4N
kvlRa6fj1I3yYUesnKJkbWMo/ZAgrN2ltjt/BrWuhkr6Qf7pJdWqxp8po72Mt5bcEQp7kZSAyEuE
vxS1xDOttq6yNJLQSmwcUlbb2KTf98KE1PkARaaJosGXT2SB4qRVhWLdiqkr1QbN5UuO1Kyw6bMB
EYwcbVmm5JjO8/pg2AuzRLpOBA7DmGXLptsPfGW4iPgVi5N56ruAJ1kAVG3Bm4iTz4K5BUX706Fo
M7WYLQcubmjBuwBaRPrhkwXzdfdpJri9SDih7f73wvqKEKpbythmAk7rfyxB01KMCoYXhr6bduxm
camFHD8xYehRRR95DVqi5Nd12Vp8D+TZPt37f72xHfutAFZkyVAOBlYrIW6g/+dZkNlt0iOvOjS/
QvhZVn9w5DnTHmsuJK+VpPh0K3Ucu0pZJ3dxVA5H95a3rhKURqmrynhXfOl2VfK9leRPoGMr9Bst
DNaDzM5SpdI/3gSjXggivgKG1k1gbWURSMFil4nEYvOUMq+ZIapNV2REnxCELLpQnnAlY6BcWC7l
+xOlOvcOw+3SKE70cKWz4haCvBm6AK8faosuuis1A0OjIYDbKShPpBN2q15UwnRx+Cpc2K7IvYb3
7KkaPbv7YkDYTT6dhudwkP3cDUhIKAT9Kc5wiJP+PWUatph5CHohMVbIgFh+oSAA125YERrg4rFu
286wQIjaZ5eu0GFR4AAEDXchL9iPg3fC1u54bMbRz3eG0lzzhc9VTp4j6D8S7ggjm5qZ0gJPMF2W
1qxCxItIzXwOPniCehpKeG3Q5+DQ7XARCSoeF+SSLdQlKq3kCgOZ2zKRZalrAdnd+F4NgcgEhFew
F0Z9GUef8UFhYUlQ70+THjZEQvTxl5mnyU7wPNEzyBuuXb94LJFqqfFNfkZK2zSGKORz2KoCfHS5
lP1VREctoUdqolTj/3YMQoYbQ1YIxnrdQpSN60bO26K2jhQ7d3OgXqC9CinK8lkjv5J8OOoy7j2W
JVZG+0C+6q+WFSWArP46UT05yh56P6BtpGqWeKvgMQgKyC7g36eMYmUHUen2jbqSPU8NXyrZeuCH
XIKzgOJ6Xs8uvcjtzH108EJDg/xGs5ahRcw6DAPqa1IePlrle72D/FVHiTHReJuS9pVW8OSLcU4S
YQAIe8THL1xeJUhCW1TzrVXy5/U5I5YYB4/vKPR4bfkKeI1ksk3USAO0UNnwxCDe4x/XLtimnj8L
6wS0+g1sgofPHF6VqMNRLMxUfHe5RvZPr0QZdjdJ/pLL8SgCZsSCEbW0T+apGPcItMgmx2eajRZt
Bu9EglashDNSUfgqvlGXZqbfysl3PjiHFsGXs6MPnxSYFfNKinXNYwPZ5sKAS2HPhjWQzde6QTql
oLYS7imaRaYqNIlSl1hGVVygkhpicZx6ugfN3S6q6w0hqojA2kvohVwJFrYzuFZMpqtxYGDotjFd
yJU5HwBUn1pIpCpf7apz5ph1Y84+HwYzGnfp8ofsijXdF305LOgMdG23lcJFvjR6dddRQtUdi2Mt
d+lJc6KAJ7X70w7aMQ4Dj8xM/fp3VIPsqauO3/H91aycruomgPVp3V6TZ7wDxPmScoafIVr4iM7E
zRNpygQA6S/m5Tq5+Twu4lt3p0/0lzdx3NWEWgLtrgXpz/Lhgs6xg1auc3gRmMhWhrZYlvtbWB23
g5Pa4Jft0ZJNZvltp5j6uUoNv7YSOStu8SZVcIauJVhyKJhsJY5wVDlJDBSLyn3oBrioeNzGRUt5
cmwQBLiJIc+WPbS7yi2CAabt3ySq/JtFxS7HzySBu01/w80FkU1y307sCAFL5jZlDAoUCfyMRtHs
iZoTTgBRXGyCVcKsRAMISVMOrzxiZ7wH3u23XD9wzW8BHJChZ+U2Y9I82efCVGEt5EnjK42ZJ3jl
CRhMHyMXQrIMr1bCL/7wXpMpKuH2UgpPRgfi6UlW31r/K59LOa3RIuFMf3v3KhHFv9gGHSknOWzR
r4Y2kMEbSMWkrGgnckzbgpwLXTCyPupI5U8Ow4wym9fat8fvmqT4QVMWXJilri+91nDCSlJmF8ic
7eQ27qDsvM3uyhyGmA26TCWSkP4LnQc7F+UNymLxuzFQeKvNxDKfAfqwMnp3Ujn2aQR7IvQXsl0w
wLwMGd88E2xAdmOnBnuW2NrcK0KrRDTGOrLwJeq6wWpwaw04vz4EWbfbDKC6uq7aYQVvXcwMuJCx
NlpaLy78RyetXwYsVdO/ftxchs7fJSXUYRpqZePgo9Bq9RhmSYwDCXssgdLiCAV6hoEVY+Iw9LSw
fRICNDg23UpzDhTPNgBKLloMNQ47TjCrco9DWu6gNxRFQW49nshTPUpHPHbO3hfDWAnLGrrY85d4
oE8oZbE5SHu+fbT0hKv6wPkT0Q2dYSz6sXqw2dmVpkKv8s6pENeYmgCoiodlpTjVTHNvwXCweWeo
BRJHVQfXCj6F7830spN7Vm0t4qv4cmLy01yT4iT44PURBcmcyjqlBxMm87AqT/9ezVbduLFk8+R2
Lv5QX1LaTrbIPZHWhQocu00pymThB7w8yoG5SbCYUKsGAJdgJdMIXssIOIKnhbK+j5h6FfgBAdxz
dEF7TbljCPdox7fO0cRC3eOwBIJE/0KGiIOVkkjn/PAuCOUMIeNK3BduGfx4FjNamCpx7tpbuhaw
nP+xvkufSN+h9LwAWJyWZmKB2RTJnv1rS4bHCEy0CgyZhM7iwJC8pmob+derijjHXuLRNIKl5ntx
LloXc8w/Ob7YvM0WRwOYZwGHIk3b4Yvo1eWvwXrHZLinoB8CXNiCzS9np05ZPYcjMfkvtn9twzSe
4wDfQXKA0/XHGpHB0Q84Z+ME3pTYuOC1waF/hpyTI3YV4Y+OdH5H46fR4M3+UCnir1Qb+YGDye2p
g7LJ6ddmsXzAUCsE3n/U617TY1oNyILoL/tB6/jixRkDRMtlhOI+FVolKsUFK0RKXmLvnlFtG2TY
1fPV0EoImozAmOHvUUFa+sLJWW9cmxbCMVRLbmsEL6UsGnbT7epF9JoGz8xmeQ1YtZYBejg4G4mF
QWyhmC09ahI/75LaFM5zqUekKOdzztBKrbL3Rr+9f1fv0JiKii3QOS4RN/BSfqksk2T6TJHXGSmD
LuVTnUeBqbxiMwfc6Po9xoPG5RDkVCQahACLW6hu9BshQn/5J++fQu4O//OOiBQKYldfxsiy2vmo
s91FJSHMqZdCj5zJ5gFmG47qICR2C5EfrkDktlyrnZgEnFHWJKhVJynPaatbAcMeBprCWrAaOUfm
3eKpPcjtNkIg/C2LGx4CuF6c1PJ9GNPuw/9dpjnMAW42QuWYB/g71B+yznnryAdkCcUm6YTi106s
BgKYqS4P2n7FDvgnkxvsZgR8uSD9wcrAff1A0D4AbygfNe+CXEzGTMZVynsVHek8bVxu+nOcniaH
qUGWuOj43Jwtk0pEQynTCr25PxZR9ghEsqWcxeufgLkM0ZpEvl0d+Dimf7kUZSB86Z4qR+SDC91p
gAXIBDzK3TcafO6I5Bek+/hf1xxA/ZeUEWjJB1hQ8MlfGdhPDo7aTwqGT8c1CD8AqJVE2PTdiD33
YGyx1nrnmtdYf+B9vOW1IyhC49FQOPbUqyy+Pr/OOO9K/TruXOZuri0WXoHth45sYMZNYnpSrZd/
TsOF2TaRinwI3x1KxUE6dFcWiId3UquufbCVkGM5iGJAo9sWa0o0TCWw0Qg4VASeyRDG05XbNlgj
912fiMKUbtX7pyqHs/6sYK9dYuQarhWQPTGv71xE4RctzjJg02s8p6Au7dmTDTpUW6/YS/DA0vpm
/rl32yARXoaxnnKheASjT3kowSRW7TWDGGoYmzlKFwwOJPkHoIHUIdZSJK+anfAM0HFXLLtsox2N
CSpOm+Es6azP6hhTHg3kWrSnNVKVubTden/MP77NBvY847/bToSS6ZRWL80zOvFi6pEVU1bYv+Id
Bliex8IWNE58DERMiASLp13Q3vUyE/eWs4hW9v1o2XTws9PwH+AtM+McyADcYYlNJ/9zkB9dTXwd
Pve8Jxffl55l4QpPPeVtAS1rqfVr2N7IojBZJQeBq77ncylcX5nRg7/WQ66CxWAfNy16K9tTxe3n
uzXct/RVBBPIhNqv355jajnTWG8YBD3jXUp92ot94I/WD/tFiczx0TKnwefuVH4sIQW6xtACXyaB
r54fMsU4db5ioqyukLXGjD70VBs1KTqCsZJQk1sFvJreGRaZKVwvvEC1484yXvvGXAi78heq+ni9
D/iM1gmnCT/EL1OgLOBEiTdbB3X7u+5CFlwP3ZdnSKkndwF56iiveSOBasgjZoY1ZPhTB9gt5lBE
lj/GJQWNfIEiXHiZiPeQ0Hnyc9Vgy1DKtGppY/ttA9y/5xvl0EBc3eENDrpkdl0c+GOidb4d2j82
PZvXHXVZqlDvhDI64mRXqXfpoPv8F1vgTI+05N6olp7Obj4QVpfNmqv1RXiNhMFrbjRpGyV8cQ4n
bPigRuA6HGZdiz0V4dj77lZ5IlW9SyeG0lNp7WdO1xQK/8ruiYARy3qz2W7OhgcxaELt52CzRJy1
2HDtuVHek0pqWKOYFWr7nKDDTrtY2qfoTZdUXivCDWEIV8vk6NGAl7LZaEZjsc+PwhKyBhTeU6Ct
3lWI4Ayls8DDJ4+aoe5kX3YCNilcOpyJwuqMu4Ea2RLOHKbdAeCkJ4YAakqcIrYDIa6QfvEZiwmz
g64h9S+dFNxI8FX68FpShsI65/9LxMuDz6CMalK8SLHo3Z69vynrK3JXY1f1wFbGlKKzs4yyJSH9
Hoo+SFdXW4G/OxTzmVoh6z1b3XzuMU+OJyWWV/mW4i8tV8ltmtX2n69bCNPgwNOcBRV6Wg8mRczc
wTZYEVgY0zLKy7nSVS0TGxVkkcqIIab9iCkM8kyiFucVz6Yf2gVvG3fSDh/NyV9SqXbYOJaICYx4
AlloNcwAGbh72NOzPtNBxG5ZU1Kfum1mrF+ZiJzD1neXa1Z/bZNcqG9QDFkFjmnMkPdA9Um70psw
RlGDHc5CwajlfKsm3F3R2qAwQohdwmCt7zEbuylX9ViJ5LAm0Cih9h1kSziGRu88OhZgkRchwzFj
Sbn12e0JWCpe//yaPlQi/nMlB/tXI/YCt1ECkYb4PRN2lTkG5qsNF7UmJCrM6O0OfPrRsUx5yowR
ur/0FUQr2na3UOm6vqegMlXeIERMkF/UhEQ7Aeja7nCmiUV7WAqAgIoMhRx+AwK617QMPUgqskza
lQlY2XwQwibKyB124qFzKObHSURah/Nu5dsA0z64hbuLh4WWBhcG/MoP9Ww/NCqrP2QqiIHh6yxG
VQTtZ6DRn/QRDkHQKD61j8MLki+c/VeRauOcpdQviqeQwLD7eftCSHAfCKtc0iXodcPgaVNdNwD6
B2+A4PINli9eWcsfEizgxREXwADRFtnRmE4AEu7CEfVPzjSJbLJL/AS+klJ/XI/f0NUW5gHHf46o
LIJJfG6BRPTWVDsO0MVAWjjT32hgUI8m6Dpurl8UTwhQ9Gnrs8PgYhsWQc7d+duac9IOAM8taOr7
pIlDdH76Cny8aldpt4FVTQYMwAUrBdtPTYplXF4vuTKSi1hjlsKvp8WOWkkGBockmlbC+cWKhn6r
qvJrM1H2ZuFPkNXoRZb85y/Z/FSQNYtMWgu+x4lWWNiDb9uEM/bmeaKkV5LI3+hh3Ni/izoFteTb
RQyVlMmN/5DBvCy0ks+ONByFPCKmu7OIBgs0er8Cq57i4WaTDuYkF4yD717Mbo9lKLVJH5uqysjV
Vcb55TgEsnMmmiEt/0T3atiM25KHhC+2Zz0qslWEZlxcu8lJSTdvwzdZ/ltU6ij9+LdmJKynIfce
+t683i+5MPxbVYpVf+01Z3kpdalOjYmxvrSDhTCszmJx64xJMwGv2cZ9H4p9Mkf5xuqkWYWYC88U
w9kqjA7yni1g25HIbw4DgBhSjEPjmY1cONhn688EAAhKQHQGVVfOebR3v8q86YI2TCj/iEOT/GA7
VJR+XxTzgj9KFvVaIpMVRxdHOa/yzlugHCZD9jv6tgT1/6UHtcuFNPHGa1kduqe7lYTpFNOtDA8G
FYI9a4TjRg7jaqq2dW8t1Fz/84CwPbkinpp5ohV8ZMStyUUNm/acesExmgOzGy6QPE/FzHoe8Gsy
GQOFGk14QUKaytF7aW6zDzfT9iWRdIKLU1bL+jxhU/KaP5jp8Gr62toM5Ec02O0R3xQIwqTcKprN
/uj2P5epqwYalh0kGDpLRFSlZaaEtRwKCjxZX6jYHmkM2PIJzPNjeMjVpM2bp2+LIY4K7DdSirbY
X8yPHb/RR/NxOwLDf+SxM88fXXGs+wWU84jJrk1Fe/yxChtswl3mukstZLtMNgCLhsvjdaNCVzST
8paa8qsGQ6Pv7eEgnxXh+R1UMbw5LJZ1bgDBTdB0lXKX4bRV0BhUrUaKjJIeQtUzwNBX9WmOroOT
uKCWTT5BIg8+SzVYI9SWjfAXwTPxDbDY43IN9bSSL11qeh3aJmPA1CF+80SKOxJJZZRU0PgUetFy
T5+kwuFq2tRaFrPIfpkvzIE/KtbGFoIknZDQMpsz/zEGIViG7rpXWAZ0nntU1GQJisbgc25zClQG
j30VhU6oj983f9SSnKckBlA62FNepAAqxWCb+ZlHKortn02wh8PHdEmPK5CsIZt87WygONuVLRZt
kwoAqZdzkqYZ/c7RX3Ej9a4dfG/u8eKALfpHoJ4Glu1WQpQK6aESGAWE4yCMWHBaoNAIILK+qajJ
JQUoX3zcRv4hxlCvK7FhzmLiDFimv47iUMCo0PRYBmMCvhjhazKwqauCHOggt+Fb+Or2Int5oDRx
FH9GZ2mQpMtOTOIZqWQ15GETZ1Yq4S06GY4YYp+Afn3fqRhcTzXWWseSplpFbHEOKLwU3v1TU15h
5SdNkNqmRfRefHFx0ASqnHv/GS+Z9h+v6kMLgUeyU7pB+mXj5tSX7P4VXvnEGDiLPDKPbAPwa3VF
AVGv2jPDn7weQAit7Kdxs7ZPsfVz+ke68fDc1vn6xl9w4KhQ//ch9Vst57YkLuJylMXMi04eaPoV
53PycJZBTT+EuA5U1KH3Z8xZcqJl4Z1nbjnj4HdZ9djMAgw2ZTh9ZkqZA24hCx5LlO7/0THnMrno
z7IQza8Q65m/t7Io2kZa5CAfrM9jw9yCvk/pcDEHI63CWXi6fltMWn2N4e68ylip+Nvwj0r17+7n
fuE170Wy1xTUjb3UwuXTz+Qn9u3djjFx4ba11BIeK5phPfUOBHZcxz67EUDJn5AqCvg2HBf7dUR8
Vusj9sCGpKSC8nMhABMkoasRsyU1aN2J7X9ug94bRTZQvEKskdkPCGs4ZAWDmX4F4uffmq2ovpNU
2wMkqlEIH6LTPVcydMuuGcDqKdSeCgLEQZ9Y2mUSUvJJ7c459PrznqmSrCKbORRyVAFxF6UWtvqK
rqeH/tp57jNO9Uufx1uSEhE9kaQHrq+QndpGymuPflvdiV0oOomcVm0KRRhyTKv74TVUhN7CuVwN
r0M6GyfdkaprHjVCd1Wcs02uH1ZrSpVgfKAdAJO96MnxLvTS0uUGafc3gucADtn4zKr4sdYdnSqe
2NlXtwD67JkZtcHkHcUYoUGZrswhwE6tbNJoGeNKwAXnpjx/QvGsj1xoqzQxyV/ATVwjsSCp0o2N
aCRI4kIzB9mBmEYvLah5iQER/kyg3uL6uTyIRg1QDoXp/GFfRRAs4YYz/6xDYpGYZPtWu/yLMK0c
4F29WQrhd9lW9c/0D0+Yy1zcDDhRmN6GoWAnjniEiSW2TePqqbU+nRpMfvIX4xA2a6U2aBVl6jHu
kyz94qrbJdgT/ocqnhqnLuBLt8/5v7QG4cv+lmwDbhWBT7iROkZQXZXW/6NJnztY5fSqQHMjdQgX
eWUS4X5mvCFZDViOE/4lav5RT/5+4QzYW2hN+m9fnjeSCfiF+j7yYzPuqgcrgznqE43qM3Mksxcy
yT0dpOxm3cSRGBUgYYyEhYImHFGZ22w1pL562TuO+JUCAkDhRJPZkdMclWw0+WXMUUiK0FMOUbRt
1d1t9A0ZzWpBiMlD3wnvK98DS+jLzE4FXCY/tudzwQ5pNRy11AU9PT7dA2RJcb2Clo2uan7Ygi7o
Koa3l7rCyN7pwI9wjDDCVnxAKDTcMwcA1S2QhULGVgET5Us0S/P8/wCk/f5+qgKnUJJrBiLUPlCl
NI+qWL0vq3+ey/nW81PybGKXf0hTpmF1yO+AIfpP8a1koYjHgTv7Ds1v+amVnzid16GKAIDc8mTu
k2Hi9RZH8g0oyj+koVyo1d7EC0n0hjSS8MU6/x7k6yJeZNnx2o8dsJYJdmdqyckrNxMKcmW0fhGg
uR2elJtSji7i0HaV1UIwA8yvoeMKIqkNDbEE6xdcgOzmM9P8hLDU8BPYo6z1304ivGpjNkHxMWri
Dfa8WswBEW5+aZ4+NSe1ss3dhCPOPU7fipFm+SZ09mNL1JPVzhgw7cCNrX12Rmv2Jj4ZgSbmJvNa
/iNz6PPl7PnpZy2fgd/jozkkS1/B6BmsSJLBC9VJus/pJVr21Cww/bwXn8+afNNQMDAJNhdQxtAv
thBeG9eS5Bdk5ukzJNxdnlJCbtWPGs8LjrCv29idfJeWEziZ8DFluTE8OaNHb9rCLEPgx79nwRKm
BW82ZUSWHtgpwx3Yof7+pAzSFZb0PURTLV9DO/D3u41RQVDEIHncfciHKV4kMVLEo3JFXE6BZuIe
dLfA6rYolE1x+hFnxsAvH3KVJxqb8tnBni8QCgpq38vQV56gz/j/xFINAdY6ncCzAa6eiLn+ghgF
eHstahCvFRB1NB6b9meY+IC7bSFlPyA+32wWLzBHIsDgZccJzs+qviZ5gV+YRrbAND/0NevQJ0UW
pEuXpMZeYNpFaeAg89CduysPSV8epSUEW1xPN2WpZJYHc5UVulde6UBJExkMtGEDcYY1tfPO85YS
koywjNg5j3URyPEKviGXGEG3aDoc0AXTWnrKBWizg6I9wDOQUlHGt+zK0eb5BxtCRlKDMxJMSVY7
SDO+X9rRU91lUr0OVi551qgzDS0qiKsEQguaWxHnV5BlL0VeU66zyWKrKIbQAiNbDSADmtOdcBrE
9wPq1mfbakM2pS4DZD7AdWeYVcKxW7xnRT7e88SJeJ7vicuLP9EZHn1kRYomFgmmG1KUqOtkpB94
hdUWSwIlF7rf6uvvGeadO+JmsJMtLny7vUeFmiInwFtqEVQt2ox386MkmYUpMm67e7DkP4Cw0kWD
tBMd8UPwfCYUGgGn0ad/SDpKnsC6SN69Y9Pdi0dARh5AorriP8wPUtIcDnPs2C7FV4B3Vrv9BUll
5qlpMO+GOUDsLwNmbtXgBB8rtfxKQqzpHcxfsdQn3hAysuHvCCYAdalu3ZKFAi45vL+W44AulbSx
SMJps8DaIcshcBLxRjr4Y7kXs+NoBmkQ8N0AHrn5/EHfXhLgRqGW26bjT+XVCnpQQ6rCcJ/5YgRd
niVubgkz5wNWiYNYEXjnpILK1Zn2omfHdGodAcMlhq1utGHh8Th2LNHdwmk9D0rmzPbFgE56fkL4
4yyJTmZMhl8Z459ejZTnhOTsyPM8rBiludF1pKpygKpDFK9V7srcWnU1m8NaNEJD8TtxeQ9aBd9z
N/LNcfeXxQEFPqp4jevyDBg08jk/gmuuZibDwmXi3nMEODVYBHtIjUsKDTbBpvp2QqwVHVRk1kTO
GoB1vIJgIhK3emP2+W612MxZyvA6WVwx2CxJxCVPLtUkXyYBqGXoSGK20d5DykhJXfOTKdHG8Et6
XUKy1hoE8VzbjGifp22tR3cN0UG5Q6n3cEcejM2/H5BsOXzlSzOXZJSo/lrrozv2DHrXRjJIhytY
QmjIDN8VPYh/deJ74s8geyVih6Xpj91cV8gIi4BsxvqNxgYUtfZkwNPMIdfPMlF3OgF8Nd6p0RzO
G/NiLLH3YucZ+w8wHbdK4zZ4Omtjjqesw/Ul255Ni7ut+FBPKudwIazoEDRPUcQs1Kckj1wr1NqG
/UjtUCmVsQy42pHr+GimcW2ng13scp/SIh4SSvzMUZmVmhmbdv8a5EAFFlQfBF9SIY80mzHemSjG
qb1579Se9tKumdIQSW5mlx2RGAuzYGIoZ5CwDpnNG4Y59vWVVHhYjTV3B9kEa8z6AU1MMoU+hEXQ
I5A2IUqr/l/f56J1iL6XjlAoFi13t72Ts8p3Q6x7pHHinEcxy5U5q+sqoHGOFxn63+W7S80zAsTK
0jlsfncEw+xoQ13o5IxqDN3wmLjjXEfvnDamgu5tDagVxQIQESiJ6a1BmWh6hLWt2GlwI6DqWbrb
wdEB7f+Ep/QtXRDIAbXXLX6FF4nmzN3XENdc5ySNZDKDuygkYOwtNDd0lX6zItcPzgSSjbiJtB+9
J7VH57M5iUAYzrpWhykEEuXg5yEINOi2SsbjQrFZez8KwrkOZnqx6yvkHjZdG/VBlkMAnxsD8zm5
WCPKZmysj9M4u/bJU7kK5A6mvlcnrQ+UjLieswo9XMTKRdLzXzqioMKm+ZGH9K/ZXsLE5Ld4OcCE
SCVhb/EfPppsbLYPFthqWncvOcUfLV6SIGk1Jw1R9ooYDUTAhW0Od1pdGJvG088y50R5txnWUwwX
/OjY6mUSHEO9c6WBI8Syjfyk4FzxoRQJfs1EB57nN+rB/Kd3qxSrTZXtuuOgSGZG2sHhkRAGnJrb
kca3SYlIq5U7BQbdUeBuqdpQh/QyXHnkQ4ZPIWqP+Z3OuN2Nuo51KlsHsRUl6hIjMRknjhya1S4Z
djWaih0O09XAgSXsrLldZh+ExViYAQLjtDt6W4fMEiQOvEZiwgwB+4QdHwYPVydy/xaRRTi7JZTK
UhDuqQC0ocpwb52tF7HKU2khC40f4hIM0hWeOKG2orGqb/K8YmhrpQyTvFV1RGmi7dsl5WQJeZ8G
NLMm8EnI7R0LD0iYhEUibIB/Uk5C1EsiC6RKWhQ4LMel6TVSV3fTQgGdDneD1CKxgLUwBiFubpoN
xu0RdIq3xFETLL+I/dDsIxyUeFbSa+I6mYGeftwsaJvEFjqsMPx5tiWelic/wo28sCG1OGM25Vng
40y0EVM2pBXHPGeJTXUdgqtrpeEK8xHgC8B+/y+2+JUGPrlYndk87PboN0Rrb/LG1Q8jD9KLr8Zf
EK3m7220i57F0JnpkiCh6kcaTOc2GSZ7S+AaF/7miuI1+frk2vu1WlL5zyyUkuy9uWV4tUrUvKRA
mbrylHL4fVeAWKbdTVLju2wk56h55jMQzc7rbk7wV+9x3LBZ9vXjAfNQQ2VicELQ/TUFlEsTX3DA
LihMMnFR7SmxfzjuA+VpxspCMb7ehJHQY6KFWPqbtdBYKzRzUt2Oue+h8dnbd/iyR9Qoqh2jblXW
gCbnv4Nyn5+IzqE+wJiRrwsKNzqTK3vd/w+MjPhVwZrwF+UmnnfPYgP/yO9Xajn+d17TchXtKCkp
ZDajf4Aw4/vw62lRr3D0Wy3Imucy8I/O6Hfx+sMM9AsUUiqtsC4eZvsZs0Mzej4OlvvHLprOssHx
HkSlB/bHdJBROh0QsKs9KD83NhWQJAamNvu0IKkLLF56mp69G8PSWny/B6Ghq9X7weFujGFvJWG6
ee9qZYWELveYC17rptltiO5AhEO2O2ngiPgg7s398OT0RNAdPVPiOL6yDCTsXz12+E7c1WDVvrwO
s+wWxM72fzZQyT1CyX5prZMPELY95hS6JA93JeXj5cjQ5gjOBeUsorTGzHy9jpLufwwrfae6GPTk
QnxtDk+SJxbzrHeeRR2hg5e5ht6wwvd9G1BdCw6YIxHJDjXXauP4r2ojhurfCe/eYeD+M3soPE3R
IjGkzzdA7cZ3Jwp8tPQTHMkHmbyQF8n5Gemugf1BwPHtUI3b5Bm3Y/m83/DgSjmJP03ndBhoOh+c
2yXtccr61mnDv/ob8QuoPX+xHHtI+sq+7fJ8zjmUMHeLZKZUmhLPGQN+NoT57XYhP0JnOjh81OiN
FrOWkSrJxkCHHheRSCviUbVkOjf3uTqDbFsSh1r/xpyQ6bkLU8jlGJYhsQNvy0odIiNRLV1sO6hp
AmVUouNWPG8T1YeRL7MOSi/DYLjEHOSII/h9g/ajE/10EGNG1Rtx3O/bRcA6bGcPVUpVJT6+J9eZ
sJEI8KC7ovlOS0NRgqvN5HujBgdDH9UEDiqFtXSVwOaEzn/XgpEEk5Vr2ROpSMSt34ERbVz1g4TV
fFYFonn0mgf73xKJj0jG1gVVTJXPhw7xRmB8gLN2JH5KTUcC1Y/PntKpTFaxBxxcGiVYEVEVBlXy
IKIRYd8OLb/oUhDPOJz+Jzh2NVhPAPjuTznG9saNcLqtfE+0xVwWVxOh619aOL0t12Z8hix38ga8
Qp8g0oPRF+xoC/UWZNASv2A8IyPyjMJwXyxL7af06Lpas1yDVSY4+FgV8UrcQM9YrFmzCeisRhYp
Fo3EdKMFcHCxmaCG5zG5ktq/aOL/+DCWHwPm6b0lIHyY4V2gmn5boreg0MDXwxU3q00ryagxJAhm
nXTF9It9ZJP3lu2Dk5F1LebIa/N5QDZF7FTxxwln2noPExUIYUnY+skCOP2N2njoq1ZZtZ0Y6GGM
F3I3b6GxQcm2WVq2tYtQKmlQRfn5pQahExJcmimdDnKCl/NRZIRspE9pTR6iEQFw49xELmQ+Xda0
cYkKdeaGXDvf7zNcxXZ2A/Pq5RfBtFWG3kmdp5bJGDlglNqLFLOAVWLR9Yy8evlgPFycU5J7XV8l
juRWWqkVTO7NtvBFg4u9N2kf8V65wJX4HgKX+p8CCAZFsJOaeIYD6IltYHQiKNqetWx9uUH/lsuc
q/tgfYyJGVhj3O3xCZas/ojXMzDTTCcOjWskDYRph4FUhldhSP58UXhT721iJeEhOICkbKZaXRtP
QYotbRRdqkh74slqBRVEs1b16SdQ3vfg8F4hAPTB4vmcgNogRA0mFGlP/g3HPU9juMrUFMunqdsl
HASVUbjswA44P/mvsiEpA+iiYfxmbtf4jxzE7Wd6V/1RJj+47I9o+hCgh69uqR0ycOBT/bXRPmTA
qYSXYulSNZRhATZVi12STDYcuXvmp0V+phmrUbtCp36B76gP0/0roQ6z1j2alIoIs3uNTLFY6Ve4
JpCDAHTSf+N0jB3UctWhsuh7CvIfK/3UhHZG+eGkPjs9zm+GOIHPXexWIM8/PYxLgy3m1lpappjl
sAFp0Mee5vSouoffX2ufgLo09wRSvD2LnD3XB6L3AgRhnxtuG/ODiRaoEFOcULXX9MAEFM9543en
DAqtHW+mwLKJ1XZlFEgUwLuAW0kdxO2d1ecYYDI3POlk14NPvMZ5X/EyQ36VIydisYp6i7n9ZNHa
7vSEX5c4MDYYCITpyUeSmROLBX851VT3MXm1TMvykU8thsKUD/pFEAp6HjV/qJIRTgUscSJXFFLG
aTUneEChKZ2f273aHR5YIk+u2ij+FQWJYf/pI5WAR+RPKfrPh+2IG7bYFHtdJT6cXYh8EV0AEGMK
m+mZv6WO3+0Isssa5nELd8iPZ2dc/LEqDVa/sPX4EXh0LNp2qKrsIQsDcy9DeFArvUEcSzib/iF8
272VsIkojN3BygxpTgXIOV/DFwOIo0flPRfFwKFbL9wLl55G9v9Lgd3OsNEoMkCYhD0x7F8RFCTD
K+kTFqmBhLe6FrBmgjXj94eG7kk+X/2lHweeqp/lfcr6YnBdzQ29+PrlJ57d87srEaMCzTUQGGXN
LvMFE+3K15uGX1mAm92z9jiDePhuB2hDwjfHhITNu5wvkEHITnhc7dqazkNOM3JOlVfxVSX6hKGr
6v/hGCKan96YvdvE7AqkhKzxyuHLQTUFP8XLXTE+TAE2K/tDxT7I4/+MCkC7W20ymGfhaw+2yDjc
Sy1SQwslk5fezArD96Aopreb1aKRe4SgdV1khlZ20gzjbzww63tlsDrJI3jYmJavwILVeudB06H9
BOET09rwTRXW9K74+P3+ygXWozH2zedycf386jkp/6TdpCrGkvI2K6qbQOmJZvWeTNzjXoX35r7+
VMFbXSpoVB3lp7tZI64+kgfavwTWOj233F3Q/0KMsoN21yEip3pIReL5ysf/eCwIpmOEY0/Btg8l
sjVw9/tkia0kCw03WfcnoZtLFOFvRDwFcjO1rS3HuY272QtmEAOqEAYBLhrkwS1r6I47B7Y6575F
T9jWNHrfjbKGn9GBs2GMRP+VkJKLffZ4QrVC8Qyo+m3Amm/aw9CrHvWmIDqEloJKTIXWwbYEndRr
DJ0BIfPSyiYPBN+GmtrKlY6i9sGxpcA2H9koie4cKJsPJ9NECi56urxVH8FvIysiwqo51ZtY0nip
LansVkhZjKcGRsk4G0DPNfpKN2sayXytscIlqufL+uSX7oKEsJ9G9sj3N0FixUpMJRo+LREg3veL
JxBBijzadUXya10MKHi21/Kttkodg9iALO7dlnnVZGJHucjDe1SGxojBjbB8iRezgrAd87saH4ZD
/nyuDDwjCEnz9ESYGwavRaGn0A5SMQZat52jKlvqi6V7Cw7YuxJydRdZsiJ0WsJbLxcEwWJdvQvI
26TLPI/Wvuw8dccfw5rWedArOHG5kBebMoHu9DsRtsKzvBQwsPvciMYt2noo4fw6mSktZ/zcVEIF
g4JHNrPxtdeUbwPrTK61g7ty4qRLit/YKTgKFb2itwBcTM4Rpv4U7k+Lpyns5fVKXRBPU5wXstlE
B7j7+RyDn2m+220fZVdiZSH4bWe6b+iiIz5bWeyMwwQkQmvpLsaHiiS9qo/A5WD6G2UWKLudqKjA
lQjgyn4EU7spR+2VtYVycchVzcvDymtGuCzeDYIo9UC06OIftHzJRvqypkShcqcYORJNVZUlyGnB
yTWWQAlks7b3LP4PiIYOkeZgBm/P5Pb6wd2eGBWYf4gCsVGd/eyRkBybtfj1BK91YUZQGIPj1mJ9
zroyJ0Bh/zaXXsMvlCLVWr+FhPiVsYYE56x5iFiFreZjiqG1bJUURw/CUNSUJH4LRTV/xt+shUdP
IGxjfkSplbzDfSPG6IXaIIXzkhuWOLZ9/X8WK44J0bEfE0KtjtPPLVsnNT1gtO3GHix+yDKGx+/S
FHdBADDFkwB4ptTuftZSMIPMu8ULX8xC1KXQeEpOYIXLGLzjIaKZ4edAasELr5jNnH5LYdDg8a3T
6Qxp270xD0Owfp6wdRjW7GcvMVQp8Jc0Qv4qfMtxABRhsiIRn1O2dEWZO6T/rzX/TFBtsh76smzN
2XcnODDiLarl9Tbru2e3k/AE6khZ3QAFXQsydE/AwWFn6MOa42qM2osH3B0hqY3uQfvGjxUjmQyI
nex3bYPDA0OC4MOAqX5OsvdwfAU3N8iiwWTTIYgPuoKvZN+LsnkYj/r5rvdWhQTlT36H4zfhQMC7
/IzOShwkyvkxUqUxJLlgZYBCH9kjPH3Kdf2jkuTESs4zkKycytY4zd7xnPvgbWp6rNKnmOOuXTWm
9CSwm6/NP5WDSpcXNnf5bV7fYq0xzoAl/lTFFTn2ZxgGSM2otjZ/4fkuVNFuF2Z1WQnKim2+dXqN
hPx8o6IbiJWMqKeTZfoy7D0Lu11SrLQhpRBlVeiC2CvLSCEuxomTdMPA7yHZaksdB5F+E25W7TK4
LmTovXnp8320fXkMYSGQa/tkMuuS587AxOOX/oujU/YpEdvovnD4S8x0+ic+AYj0XaPH2UocvNbk
qQIBaEtM64JgkW+sH6af8N0CR7u65Y7bArUYdXg734M9jBVjlS2zD7hame7GMGVZSpH4XXrPMyoA
xur2rtIGZSmZ97DO56GZQn/Z48dcHCphAhk6WfPedGubb/DHiDQCTHGM4lW2Y6ACJ7R5BJuNNd7/
dg78hcXfv2XP5dF3loUySExZ/OGbTBAeU8G0aMLJm0f2cEmlAvHf8IsvU3at/EHDEaZkxJ29vzRX
S1Mok34RQcGq7iso8jjd6Hfkilwm+6sIE2BOSdKY0Pe9ELtcmhbWhO5Ii5BKLmECwi+3LGkvjyLq
3CEYkv1sVtmdTmqG3L+Lpm6D8GKwCPHUzZSz7Q21hfd5VXEbbfgJlwnPIccz3iXcURe5Bkful6RZ
Mve5AfxCiUNeckuU8Lekqb7kR2ZSS3pY6nQ2jpFmVK33tVEnTZC8f5DmHCXwi7MPXyq42ba3CIEw
zjVt9wMgQczA+r5b5Jq09rV77dD/BnA12QeEruUn4g9kdWV/5VV49RMgrYwcMSpIWNIjm2t+d/+u
h0LM9Og6qZyhhHqP5G2ZuXYFJ7twBnaBxbwm86gJGHEQ29Ug2NSWHyiwZ77582QGn4T4taBW9/lw
aEsmYvTsBgCT6t9InomTAmtzkJvaNt6XV04nFAZhadXRtEZMf618U9eDnTKWEOo/CEOdMz0dpktg
7ETG83VCSsO+9beZPzUsNZ1t4Pa6PabG3Gh0GurhzCVLfOjR0noj8W0rvr6MCKGmVyBAbmf7c2lo
nqpMDqFFqqIzV/yT2mcFCyI6tD5EkEy+SUkotD1SQq7zN50TA062Nz+XK2x95BrPNbebY+VT4uHg
8ebskuIfhHgf0TgKorW7DInqQn3NBYP6rShhGq2GaISLJp92QOwziwRrEtPu16nL52kjUKB5VDA1
EH4DiAjisPLmiPpRF6p51XM0An6bihDGCYoGzL93YI1s4+I4dmavqcbJVG4UDlQQBe2D7A9/ACbi
CtP+m1xiDfN15kTw52lfLk0MXkehpew9zKFuxLpN2qgjrr/21h+Qw3ZPgGC57D4+rPFjLIrvtgf+
mVqMQKAdXghwyBKqzu4X58kVdTfUtpVcTqp0OCAtbmokFuwYa39cgOsQWu937szWDGqRvbIQf+Mv
+AIJE2svKEhJIcDu6KlS+e1AUMd8H80gmIWnQm3ZOgoEPH4j/q0GE9yiFOObW4wipbS26e5IYL2r
P4cwdyc/qjjQfyJksYL9bCUsSXoJCCf4PS5g07/PM77xdCntqBXlXPA+tqtGMlW8+nua9Oohgf93
8HBKPmN/qBM0THm7JUD9qAYIlZIYrKpgttUJH8TDH3FObZAm55PNj2LI4flhMf8OMt2p0JdmHIUg
ZPtrxAWAV4rL9cDcmkSo+H1aiaAzc9nLudzisuGoaFOEkrw9lpOPq4lSsLoqpCKYqvcm2LN0MrhG
G0uwSM+u3m+9DvjleMmClrrgoMQ99WD7YRnNvYA1Es8sH2bGY/0wEn/o0WWE/YrAsqAWdc3oZi1Z
JPnBptFMG5sgf144E0j3AXx3m3muMbUM8fhzYrGj12FnckQPCixTuKF/9BNFcuc81ZQmw1GmKG0o
QKUb8M8zP2TBfQMLMC5IctUZv5sNILd/rIBbSMgs72+mlBdgqaPWx9AddlD8BPoAPH2QRBq0Yi2j
LnsFKpW6hKmkJOQtVT2v08cCh00cd/Tpa6YNl7tfLRVE9RV6n4wW2fGCNZRA/I46S5kuAlyVw5pD
rjUfYwVjBhHEiug8vreKlMnhsHAFDakGBa3ZxtpC1Jvku3ytn8w7evIIqFd6qdwuJmyz3fOR746v
Ege1/syQeoazvhNGF61bfsI2rgaR5piDKy402dY2/CVTlT/UuWnyoAojqFjHYjiFlBzvnGc5O0xO
G8qnnPXAf4j2sdA79M6g8QMwkGigTx9bR/cCgdrQLNcULgssNmaF5ikkeln4xvk2fJ216syBezO4
ipmXaKZRh7PWTlJ5PAN8HDTjVJD8hn0QleeRt6PEaBtix9K16TQmiUAgQs25D7Vz5lyWUHGQW+AF
iwg9/EvMN0ZZ7+tQC/CXR8Ph7nF1LfDAsdR7q/gakuDgJEuZwgawej4rDbUeTHZLFo6bNfNpJebu
mU90SEmvtefsQZiOCCk3mRoaHqBYxVwLFtyi4+iiGAG3N/qmdjytSwrLGKxlPaI7qkT9SDybtWQr
qaXdmuGQZh4QJrFZlKDUQXi4x+XB2vvH3exuuzY1yvD8pn9mezBzeuE1Qf+AYWMu9Q1qJ8y+1QqB
7cpT6id7gM/W0XuQg6Xb65OZjFGe3Kl7RwgA/F0drRTILy4chcVCqEqqqVhBwiz7GrMa1/fHUETa
oCFZ16dM8OWftCQ1uxvu6MUFj48eoorkFvjIbsQawHHlnGCuN55Zhn5UYGVTbupvGqgrj3GbpxPY
qTgbiZlrTf43m9dfUo9U3Dn1surQZkyPHZVTd+K1jobhKyP7seaFhfWXDgy+xgX6z6wNJPnEYFbA
Y12AnbMzxzDW647n+lxZIJXxslCl8RHHNypRtsEX2mhHY0EzqN7rTfwd/tQdJwnYRHzhxvwCr1kE
ZHPv1Zhofl5J7Rzo4Z2KDuEwOh+LcJyPyfq1IXYU1Ws9tZbbNwEy1q/JX7R6AZ75PGj9HbUhOii4
MDUqFa9BNO0pr/KnJDicpBC7JjJX42NRV47S7SrX2zSnQdYm5EajcevlRk76F4xmDGr0rQqIkVZk
u4tvftaHWUMdR7OnPvauHR8fufWnp5Ron02oo89NO3xBIU4m+5pvCWTF8XTO4yRr5upPtDbUnLJa
evym2SruR7+EShEVHFzlUKThxYc7LEmj5XdrgPXMQlTvU6S1vHEbDR5lJtL0lGC8YZkhWgjolKKI
LEnAqWu4Y1g3VHi7u1DelQp2IW942kZyln7r69oWOf8CRc5IaKDwwtP1lfzZ2FEx6lg99/imqDOX
lCkzHXNfFcGyCqlsqjDyvJIWn/4GzGstjKLHj/y5c8Q56bPSXj6k5tXrb7Hj7mOt2eTizuvvsOzE
qgO6lWQT7FjqRzeHju0z9lITGdOxYxAtc572G5tRxt8VRP87A2LqYWkiNbQHYm4sH/S2ayZYJnFL
P8uGVm8XDKLjYdglPxfn+6/HtLN8HLs7UTnPhIEGHrGIBCJjFLzV4cn8UssROqJ7f0unVD8C6u6U
Q0Te86hwTMS0cxBS9Yd8hhtPr4OegEb2dpzw5V6R2IdMJthg4c/ZL1bCJ3UXJnZf9wYp+TnrWls5
lUsMybvyoihmAKY3zHHmVdnLGjOBOU+DNvfV0Pq8MjKUXiKzX9lFadF/+4XKG5lBNCs9TGvbelEC
x5sEYkkOD6PWHgRfT291rP07OmagMgvlTgWM6rPtT0aE5oLu2vhw2E0lV6XTU9S/BRl4jHH/UWQV
95d2f1+Zz5m/WUGAOHWm1stctu+Vva7e4KDo408QAQ2/UO1S3K621ufgE7hewncKcOf24ueOp8c0
SiXt1wFkYOVDxT1lryK5e1TqXmseULtpE/+pUsejGXebNUHHVMvnvCxqtkzJVFWuljgROHmr26Kt
EPvnrqSpoXUcfiY0C1xl/9tXWa2syIkaCcucw6w7gh8qsWcfAs68aQUhOISF6UsAA4kSbwlSqkXo
cEli0vzmyrN8PfYUrKWknwgzJjnuMT720URxPVKJqSGZH5KnAWkNu9V9Dl+yFy0tgEGRysF8TXyj
yGb18+fYHZOxvFG9QJYcJMbWWK5pzTesMyQX5cPVW8K8Jqnnp8FKZQYwVzCQ5ZZaKMI83lSfY4nb
TJrPJ26I+grXg3uuYOtmT0FAsQWY+GC4qLQe9IHotEQtskdD+kijAtPXq+lHuewFpMJexyxYyETQ
EJcLZ+UhErkXwRqUJZkHnymAy2lFIz73r8bjzOseW8c8vnhjGPvzyCQZAJfanZFw4asMmSBt/8pt
U81Rydm/NTC1Fx+LV+27MU4qdnurpoaSQACbUyk6D4Xc78rttbhLTyM8BDIY+l+kehNAIUlNELrN
KazL4cfGtWBdN1bxd99r5FtJ+vIuIg5PPGERaHjlngT4aYvhcIcpLaFGdzW2JAmEsUBgtRE3eDGZ
50MxQKaoyRY+dDlQJZEI1HmhQ87qRkV7BsDbnd7Yp/oCm42ImW2IF84SM5dFJiRgFworZ+qoAuJt
gIPsERy46OQtWJ+eShJOLhPj9FtAz3c+g3fPHzrYylV2UVR/a4uum5FPTzvQ4h23ylm5TfKye8Hk
QABZHZeLKCvAAsx7nNklaFbYEbiFecwuxeQ9myo4vhoChnSZlVLT7e7dq9bBHfsXBBPJL1QWzEoA
AjFbUcXbnYeVwAP7WsyryrsSqvDsXtiJUgzc8uhv3TR4Jd2Img5SO17UCmDaGN7gJs3lUSaPOpgN
T/nEr6+IHtqbmET3uATtkoY9hwPp/+ZUwHZ5KKsOwHpHEB74Mmqz6ZvZqkE3AsWXKsIR4GDiuZCO
TArVZ22zq3EP6wbVV/b9EsHkA/AZ3T2wnm7qUg8Zzr3pSy0xP0jHN7wFKp4tPQkZZs65rCGXbMpe
632WR4034LX62GYvf8eNTvac8IfXN6EHeantmCxmvM5/yjowMG/kuXO8HfMN8p3p1qzHAtUtOSUy
XB0ZmMOZKcCDnbuDtAJ6K2b3bru1WtXDs1PHRUzkbELds1AcUmP38R0xH7XrMyiDpkbS0OXP0yct
Atf36TA2t3Js9++I3pTtdfPfSQf//b+y9E++cgPKCZhM3Q5j22ep/XPmhvVdOpy7gDkoC2QBuvHL
P7dRvs2a9OYhjN2xA2xxc0NjW2Dtp4UJZSm8yJvzZM/KPq3gvEbwfInG+n1wdhOU8tlNFE32IuCA
LCLcfEdd+Wm6bRx4jDFp/2V6UZDq8lCE/5uNfEeTE10D/GrRDkYRdqjAm8pUNpsDkg37Qe8a/v5B
fNOVKvuPtc8VzgH6OwT19ApIUAC3jdjbzWjM8WK6tJpE2et2L5LYPgvckqI/Jq+Fu/UiKWfCNc3i
8ahyX+OtwZJ6LI/NMOpJlJor55CajSEg0GblehE66ILma2kDklcP9i434EZHtJO9chq8ZC+eUpmS
Ak8ru+GpmO79LJLZla8Po0Pck74dLpzNnPzybotXti0S3aYI75GMXlbVLcdMHlfSdftu7EU2mgy/
UBuA+4jF6GvHOxge279OBuobKp2xkZptsh9qnMQwsV+lSwri3trbojgVSTNGMLJpxELvJYMqUlXB
wSI4S4sk9/5YgePepuVJ72J8tk4jnvmzZk1VDsqlpmyXHkZ4zgNXzxqr0B74D2ma46nMCIaolOQT
pdNl+k/Z4BC8/DeAwIhujypSAk95Uq2KgcqTcdQVrGzMMx8u6QkhZquPy39d/itSlwSFli50hvqg
TSUUBsXyNt7GRFr3wY4HU7KQBkySfWi0T8syp45L3Nr9+2T7Sf37AQxxt37ZwIdHUuKKJiLeHK3Q
XESGWjc9x8WLnJDyHfPpukvWseZTl8XvDTCnQnePYbwBT+T6+O9yu0axGpP7/FebSRbah1Dz+c8J
NaV/fLc9Lk+DdZ3zs50TILvl47EKkdY0TQ8T1883hf8xSamjVyc6IKwVdXBneXEMi8KVegFqvRuV
UzZU67prdQD3FColPa4MGmni4dYCgbs1BpfYhhOmwASE3mz+wMLqZbBRCOZ/+lsW7EU5RRmkI7cx
DP2ZFkIuz7hXazN9gamiohLGbpRfM19AEzwPIo1A2I0rjmxEG+DqOxiGbZo3BZHnuXe3diovrx27
PA72ngOkGanU0TYgD+qPqlzANRu//12e7TC5g0tZFqh6FVdVuYVsX2yuylSHNAOaK1udpZQrOwBx
3FMNLBwJy/Ip0eFaBKc5mYGO10nI54AwicwtUUCgKmydC9BU4N6HnKp/Oooe7MIvJUYWL2Uvf8de
+51kT0pSoMB0htsGe0jYQeB3tJQfgnBTKoSBbCmjcYjBQ955J3Hi2OJZg0c4r3haqAlFr+wKcnmk
wYhQmmB/b3SSoNdNFaYdzzRjHvjPd25HD6ky8zz4jnTJtQpDoC2mQ5cvP3IPHsuGU1U0cLg2nC2Y
mW4JEdIebYOMfexzb3mwyf2o4o7GWyt451RTVjmF8IjyGtBLapYDuhEZhp8aP0vKLjq8XISQW5rq
NsgD4VYHYFHXKTVZ0uqT1MZjWAsPDm47YX6I48grHSScMXdBuVxcNsZXlGj0HMkK7+MB03g100zJ
c0NTz7/i6TIULdS0LEldJEYRJVZzo4lCOjOnM3lZw1s7WuHOpiySLtnpY/jGUl4RCacNzA7P73r6
xCRT9H9pDhzp7Tb3sz0Zbb6GWtAX2ChO02Ri2dUguh7xuf1xmqX3xLZPZTB2PfqF1dk6Ukc2I9Zy
xyNskIYdVFGhuqOLVj+kjf9OywFvxVtJH+bTDvbFqalgP54OuFHLWMHNt9Nz67iX9P/Q+MxehJSa
/Oi3DPKQ4ovt36+1E291YsZS9zcshQl8Q+PpK2TdH8H4O1WmPxhWOKiGW3/vhLIuQUqpGxtcN4TZ
VbhhFhexDcId6TKXeR3vZ+uhq7eVbOsrj4bqUwfZm0FiNb/ZCaowh8aqOUbiYonQ+JGEEb2vRUwk
zDoshsKLS2hVI3bExiBMSIjKKzaHyLQakSEhIdBRUPTxs36BwZkNSjVKdj2Ai0etsWkWQF4Za5u6
kyIEHUM/eQyWJG4PJU5GTtF+jBFvT75YE6JgUPsMYC8IAx6cPHgxMO8yIIqy6Kr47DFqpZugBm4K
olq3Cunp44ss1qzCfV2G2Q+av4Dhqwj1J+RuY2UAKIDm9SGwpTSFkzq2J9Qhycrvrer+8VkG4Hng
jA+VKX9scp6eFNQTfJGGWXEA6dnlniVMMVqmoywZZlGREn/lWf9T7Kvfc+71bCYD/P/q1Jq9Pag9
dMj/OaSW/mnWcHohNk9XepfKIJQhs8avQGlAgzmy3PfnfrfUGV5wTIbtZmIOLMijCNhSwMdR1k6z
euq3uIYdpS/qnaBX7uu8hl8PjRyYUwZ441SBX1ygmgO6YJ97+duwiSyEijHLBMCN9f1YBwuOSS0n
8Vh6HWZhCmkLeVylDY95t0jyFkuKIQZoQzAucZUYdWxv5Ai8YIE9+zrb+YFVx95BlQlAKNZCukPe
wvLDozG9D8Vwnx9eXRgHQ/2US/5nTTfqJxqIaXyQVizFzPJimxUkTrMMmr8LEZss1kYaWtnf+7vI
IC5Ovde+LNtVXT7Vzama0L7NHzKv4KBhQDYyDRKk+A6Ku15wGltBMwfrTI+FUaswh1uoSnT4LQWv
KzdQASVVukuZ3hLw0T5kUoE7ecyH5pwaiQg/wZUf4JrpJuS3F9YRTCa8a9fS+nZgUpGRdqQMMbTf
WhDTctvw5xnWtXcyqfz2ET3iWslMP/gZwtJX1RiyiBY8XypYla3lUA3vAz/5Q5K/AXzpY1dQ9UsJ
lwcgB8g+cAzKBwjXcR+wEb4O31MBnOq15Ct7jc6eBlJHqn8cmMs9+TRdkn5a/HXHr2mKOSil16ud
WBvGrRgrnfoC/QtNqycenfBhd+qhpmk1RyH3XdV4oQ6PyJMzToel4bsT6Co6qdoPFo3kQatHVRlR
mdSqvZPhF55ndvpsM+E3UukGSH/1GrCNIoJ6IXQuqKenlqAtne+rK0v4HmqVvc5inpNLjgJRPR3G
NiQRzLJocu0WsBSmbkr/pIhKFmyLMHCH4F9Z4SAvD0hhAMnFleXKeB/czh3nmNSBiPcKJWAbwjpT
ZYxTqu0dzS6ltOarCyU3RhypaAgD8VevfAall7bpe0iUfbzR2QhX7gcUhTNGJX9UzrzH6MXcWy83
fsiHiCQ0Ozx4B1IqhdbexoKbAukDDZwt/VPuyK8QcWpCimWIvkOo72sPWy/8BOnWexojortc8cfT
IkZkoVgPM+TOhsIF/ccH0EPG11GmVBhSKMI0mPybxT8D/3n8fPJ0LoU8yG59Uh28cBalXfU0RWfQ
PAlovEoi6Nyzn7UkYyIPtvzHq+a4ecfCiPKjcAd0j4u2Ybv+SXlz8Tz4AAUvVo/nDIN25ZI3ggWX
f6Kpqu9afOlIJG6HRQzm9tgbA/Mk9IB0tZRhSEfv2NSTVDzS3OhTMBg2QnzCvDAgr3VW4kyo0uUe
xuAhIGboSKOx2gSPPWEg8zunZV5CyGNez7raZwALiSuNPuT91MIk1/tkw0T4jlRm6difGHCHPwH/
SyQa0uFfkAtWR8r0uPIq27dBMR1boson6agWuXR5aCiRnm8Jq0vYjz+FLWtRi8IRo0VHnQjJzxPF
20Hscu5yX6JtVEAErFrYbYKnfI4gKC7fmGh6oyRdbuwUDm2JY23oM+tjNHWszraknIZkQ/f+DzTa
pWkbDoExcjp5QFJbWXXmonJQezF/dFuMqhWHzGt393jArfJ+AtOVbh1kSi9FtXQ9oNLTvgWib/DI
sjEN11KQ1UEkAWMGDRZrFS3EAFPSfTBQwNj4msgRu4fHU3nBQAwLmP01JRyzHIWpWBsSyO+LOBZ3
af7iNzxjYsBvz/MBxUnDXSjLcyw2p/aRw5FJjWWmAFMX4i+jx0dvmn/1ITmqOvQjMPnE7f2XCVfS
xu4pJbwlFQlksmFUrzj5RV+bhmirNCNDRljNrpBcFykA+nA2Jpkv/vJOUPm1rrhwG3hbJuV1QcpE
OXiHwdSRDB4cB7k0UCsESyZW3uo6LsgTqNQEY66PHEQ1aK2WBYPcaSk8vmmic2DgXCMU422dFISs
l4sc/l/+CXQzx3/Wy7FeilW7n1qBfsKAHJIA9jh1D6iPLDuI708025Vk7OYXct9vWCVtkQihASz3
QNZ2KG8v+L3++nw/eaLLpnffCq+X8mMo+WT4nEnjGGjRB85b1F5wOJK5T6fPNbW6/CuDCwzLnXcB
Ncf6GUNsP8YJ/rvBYAUzpBdIT88SISmxs4vxT8RV/zWN8L78/wD/5e5jrMLwhu8HuKWJLfsux1+P
0PjBgZs6qegixw2/dpuKyET5TqH0/CC0zLp0/o1bjPUoDcvAO2CGDJ6tBJoFJ/GZajkxaPfV61Zo
i07iuVKFvrVIBjR5fi94JVOE3+FT8qW3FSIRi6iOT809dnYUZYfW2ZHGEl2AClUupWj8v1yH1u/Y
vqdKe+9aZHQc3MVuKsemBh9jJLmlVvAKg46ohSNH/qs4QaTQ7Wx20T45EBa1DxFFODrLndF4lnQZ
DuSTzqZaxL7tcZNICuMdTCuiteRvQFQKGRxkSR/2HjJLdIFIMmdpuFYBokWevNm0B1HrpfQKFUDc
MCjnBEZKMkkpejmGI1lUnmyR+rOByxKDhqtaXCURFWINiz61uWGr47cKHUGWOWjzXGPmJgJOxNcX
l4wIY/KUCaItiI7PfKVGk3LGofqideWcN6MGQYzbv/18qK9QsmROyJP45kyXpm9u0jTx50Jf30+H
nIlK2lwjb6B7VKshW5vNzkLjdjmLDV5YJwtCjbGbWYs+kHmWtuqzzpGRFKnHtNipVF0F98xjrcmd
5K/gDk9uly0mjTFHhx6JorjkoeHj3ILu2IyTsFzYtQA/eq8K3AHPE5UtmAMIiPQl+GThzWsF4h1P
nrwJuSVroXwT+bS6rpK62RSX7HCT2rhXStIuG0w3d3AVXelFPkrcVY7+dhAZjrGlBRApf05oQNA+
GPVLOOFnRV+AWgH57zF0jSLvmIRXrEDGuZ3NnOQcATx0PGOsPGERXNrjvu1a/ty79ghlWR+PRE6+
HRjqegZr0sMC6wnuWxdae2RyNBxM8vEhemKGqN0SFfTTNIfe8IlJGspkhTeX8FXI3gorrWQKz4QC
Z3RWWp1YLt09dRellWz55+rzwAxxLClD5ZtcAuU/gQmq0LXeO9FpWHwAWZbga0AuIHxVOC4hB/HP
haKfbQK4XtpX7t6+Tdrb7ApjUe0QXUPCcVIJnl51cU8hw5Jou1g+TrR8xQeuifKuQMp6+ZNgd2SP
jfMz0jOfw1FcJyetQHpNb4dqeITgddgh7fQt2JtJcAO3JolF4DkmhMPxqFwB8ifM5wjq618vp/Xc
dRvYu4lZ8wOZ2N0VZeup6b43NbAWVFvf45b4cDCG4tF6n52lI8+vIHQRVSTsQPnrGG3e1I2uTxTy
znKa5jBqGIuMQhdhSpAVWCPfnC1nd9GVwiCUsAbXh/0t0wHRgzT3t2C38pGMV5ecbVNhC2fEQLJu
KrsPn2LQYDsxcU6BqkCe85joFIpGDd/Wrdm9cLSEDoDxCxLcW139+7hbZjkJifoGFK7eBUStPcFL
3rkplyBAhkOwoEuFDOkth6AhCTRq/TLR9g1JhO6/G2ZDd4VuthddglSe1/k+paolSCng12gpaSkB
R7n/9h0i81bbE/NX6KlLb+Juwl0ZBCr9/VRItabpy7Oey68QqWlBcZrMNuLgCBTNoIzWGFm58Jy9
kbHQOLqgB4nqhtqcw/qDrCZYLDu/RvV4X24w7Hib7PvzYwVXklH+hc0sVKNAiXyetTboESHEFHRm
Kzws0DDxRZl1cualTqR6NK3IPehtg3N37z6NqSZ2BOCNHmHpICFXHyx7CwAgtg4CAeIfyg2hu0F3
sj7fDxxeIoaoM3ykcRUSi8Wt/R2FEvlEZ3/y1mta+XQZ95rSHKIvgNJCqc46DVLxeBrtM3gHvrQV
zvOpLUeP1CeOqEX6WY5EUWpn+f4r8oOXd1hjuff7T4aNHKCPHYB3NhUbJzeVL5wZMvktpfm6ZvZS
wvcw6jlatsduXL2I4kNkeSI8VonSkIqRU5vYtRT+tpkc8LO/Mu8UMXt+WmP+IX6Ypd/u8P2SuS7R
QBHET62St1zn0aCTUs1gwpW+9wz2NmKQN0hB/uKyR75pvV1ucgBfn+HBz/jEept+/dMnmf1qhqm1
87PXOFNXo3FLo3VrVHS+qOK79dMjPOL6VRQR9frXPumzyBVL7WE0BOuQe/XIIasbez8GfzrsQD42
tnZPucSkCXbymhqgbSdSWeRdRasFihw2AXywGlh2IJcELNemS+P8JiW+dT5jCoggD0eEAV7Yf+KB
X7PPJj385u099DmxqVgRTOBMswi7CRbp+7aVHv5TmIse5Wq4MRjrDKxJGSZURQlGrRLn0OkRnVwl
rlNPFTkc71p2DIrPFX2NOTLea5JKCCgXTzo3REU2iak5e4w+8eNrdnUkjrx7LUuhTNnUhB8GkMXK
D0BhzaKOBwqa3SPLdpG1gM0M1iev6PmzGyZiuWcm5feqZ19vXosqq2vLXbF//eD0GArvAgqkGKaE
tTIWdllk9CWSXs5+JpcD9bm+1/cwzlGFVP5mVdmsHWyuR9MHdErT2xy4An7Rtf7imWUmoaPE48rj
0T0pgRpl90LrzfEK+UZjtEK5P8Mz/zpyrcPKm5N3/hI99CU7RQyM9wqj1y/N1ecz1S5T473Ycjq1
VLCzHRpmUB/LtpDgEAT2qRX+sdCB5NOzFEZpYF69F5ZwjxTNW666fm1qaYg+pQwitOxMd6aU8Lle
fn7Pfhz8XgbGuViSq5Tpv6RmL9BUiF3XLufnxEY9ZEZymX/CCpDNlpbinwxeh2rPHInBUGbencY0
WBpnXp7xWsd04mbab9zp7NkddW71p55bxZQOIp53KZbT2Z1X1LHCt939PbbJAe5NHG+noVRsh7XV
l5BLqYkWvlMuUXhX5jm1uVlvjSosfq/QzxF6Xvbv3punnGa6g7yCxdCQYGMJuJ6Hb8Ah8tw1UOx/
T0k+jzEW6Db/GgrDNMWAJh1NPDJsnYAUCRxTxpqMwSrSHRo8h8DJKo6dE3mrclOVzG7FTm5Drz+y
gh0kSpnX4xrInDJt607J4zlnVChNtFmRaPaYYewzSBkVkSAzEM2KskteHdag+wkzw3SuijfmhU97
I183QOxziazvnsDlP5peVdm18orSD9+jullJuFjgBGpqVjVQjLqSkLLCIZA/Z/0tHPSRaZM+tzmN
uBSwo50mD3t6xyFFS9Sj0L1u1zF4I5avYCmYcc9/oHWQy9H4iT0shvDXkrAx1XLQ73/VXc5AKmPW
MIERsplnkCSbWbFPQZEMdiYH+Zgyo8LPtyJMKz1l+HfI2C18IiA8ymGzQrWe8BaF4fYfFPCgf6s3
FZuMZKAODZv+nEOmqdcKpAyW4pGGCQvnSBGlDwM5OVNwRRsF/tAb4VIys7i2SBOQl895u7xVGE9w
alJ99KzwVVs7KO2CKO9ArNOxd584GyJXrNZeyewjZfQWDenYHiKOwbAYMOE5u5dL9bIF1SHSRqTv
Agj37YTZfRu+n2LAKyx2Zx1FfVVYNrfA4givT/yiv8TbNcitDkAo5uxeplKiOR+2smmuR52NkDBd
Hi4kjC8KNmEqZtoYluDv+op+by5UtL2sdaLtGputkMY4OvlE2tZbA6D69todww1GftN0irP9BFe9
H6h54HPBVQOET3eMCl+0AToBsd58LKS/XQEOMgLNZdqPOLzEgiHTvj8ZO4e/egkZlSoMcVS4FsmJ
54mOlYVEI8+/nsiRWjzrBDiRyr8M63Imvxb6+1BgdhEAZ3RraIfvRGurDzLdu7NhU1M5nnDR37H9
ULjbsjOIn9P64zuAXvjoy1LqkSPP0EDL9Ty4XE/Vsj+UXaaN134K/pyENFITfqcgjv+CJT4damKY
TaugSjtSwIQnaAEGAZ4Nec+jVlJ1See/xt3WwkMQrYRYfMOBtY91adMg5EO3ZoaeD52MrC69pxw0
YFWpF4gGyveGgkJgVAKny//6kJbnls3enzSI9Hq5jrkdbAKvCYDCb/GNaxy357G7jl6dHAFK7gbE
S/tingm3OYGskxPlz6HhJ+RmfN9hIUAb+MVBGivi90nhD/81SBL0AIucAw3uVgXu3F6Pqkwxp2rz
x+M0XXAk5e10Rq3FSboAct/q7BozZQFnJ2apMd2LowZpA1Arb5jrqEsyW+fFehMpS0R7vi/R9dDC
f7QIl2k2ebXKGU9lu2bBcH+b39CfCSe1d4v51nc4Zxrvg2UnKUJ7TvUXQsoZO6+ZpWBJ2x2IruMH
CRsgZR+GnMuWSrXUSwVi0SSfESt2QknY8qNTROJn+UVGPtHvb3r1TjMvGdA1RMxlUExD9REhauX8
ar0P2oDcN0Rb3CutJyAt6yO2JgREDSCfmh1sZr32TFAi4AQT1vuLgMFsiQPNx21/tYODQRew4eoG
bH8s1oKeNisNK3v03d/5ljMkZT64rl5uR3irR1Fa0k5SP65yfij+wwYgrU9moOab8TEgoeOiUaRe
RJ3dvVjWY+33xdTWFw10EKdY4T2fHx+A0eXINeaJKIFFjgnpfSMzZ1YV8wjF8uecm0EQY1LQYgYP
xnUP48gIOLjAXeKe7dH/jK6fC3SZ1dWCGRwawneepGFBDI2dR7z4irNBuwRHhvRlmkzez+Z2g23b
0FUmGKNXq1auZGAlOSRmZlJ18e+GKsjRhRX6Q4o1whwH8JqQxp06fPs2UpJLYN5Zz950bRwtY/nq
3IP8qsowFuGoL3wotEbQFBCJ8qBI39j0Sb8MfleHBMgyt2HaiLKrIyLb9xHjG7xwMzgV5mKMq1I5
g0qRPvWMtCmIHuOje2nd2QJFnJeX0jYlsLr7TImDJcoMHIx8t0WjfheKVUU+5el98xAsvRE9Kn7B
aDqjO+Hz/LuNstqdcNjx5x4XxdpYaOvdM+cCtVJ8coIO/nwavwvwDMP2I54JgX9I9r6PJJzLEj4U
+KByHRS2aQng1nE3c9CoKmRckLY/xnwZs+QQ1gAULuZ7Yx7iMC/dgr3xZPPi6ExvbQDrVOuIhx3U
E5rC4nMXR0AabObZI6rvjt9ZBH1l9i1bLeqZ/KEv6ulHtdb2yt37lS10qIlGoQSpQhXSIUumwUyq
WY7ENjKPA/r2oAboCByn/6gY4tPj67KQtoPyV4+WM0k0OBCFaGuBV9D0OugiggzEZDRml79/LG4z
vgyrvRrxgZ8iv1Zk1+2ukIbVx8+GHCmNmaXZxX2TJiAFO896gtUlAQvavxZKEtykW4OsqCWF1sxD
FWx2F5vTEBA9Z4GzX0pg3F2uXPdPmlGO464pMwJXywcz3LS64ObaAradMOKvqn1RWy2lsK6f4JCx
M/26moDvsTGM0XX4Nat3PN0XDJFYKH9SRGOYqP3Amz850jBPKu8HHFc1KYPvnWmzpOy4VL4I4E4+
M7/5HN5B3btnQjJpbAQqYzZ5Noj7H/3Dgid9d8LSNvEoqlinBiTHma5B9oGYbfIcZ2MTscfgcal0
x7ayRleG/OwHiyu4mbgLk9ZPgSGfn2Xwm+L0j8vuOsR24e/uinfvv53guN3MGaWML9mc6K9icfXg
rrfsysI5Ft73MmN8+bfsMTUeZyvN8ddQQJy5uN6iQoCCUgvRbzdQwUmb71AOxnwcQSeFpDkKKzQm
wvyf64/ZTKwKmcLYdqVxIOuD6zsTMg3RxJO9Nlo0TapJYgThu3OVAgZCOEvIzikEviSOtjYBzHF7
9tqGDRzchZMMvqOKRpJnjAQ8yu7uLkkjAmw9XMCVsFpIx8gXXlnlhU0VufZAxqW/h/Z4bx+IEOXE
RezkffgeZ8K+r1ktHQ4J6VmmE82+4P2KpR9i3zSp+t2zbzXnJvOfXsbhacBhuQlXYwWPIjXlv4cO
/h0vL3jUSsMEqd0lMG4NLe9jVlvZIcH6gqllYRoC16TkAL+W4z6fDNmEYY2Fy7HUmMJPzm2gA0/k
CZJrZxWGU6DXFJBQRQ2sdbZ2+muotJ4EwXWc3XFkoQEan/4+YLzZocVl5UYRnpQioVCVnn9/O7lm
+yZvjFlFOfsy/TgEmwZVDQ1vY4uvei4N1xGeKsrmWcIrljRGXqK2FBfmXnxYJLGHs64zdwzQdzo5
+YaWu5S84IXOCfb6JBuTzWyOVH5wiv5nMF/G76OOb4Dlw6jXq/m8KM7gXBD2vZkvPdMy4d+fdK9R
c8oUBvOvkHl+Xee0Duxosg9oEk94pTE0rwQ5BOV3dzUe0pXVogyLFuiebhmIIpWEYCu5luVW3q9t
GNpubzs/GSa/74lGctRu2G9DxOU8m4ZikhbVRErzNUPypltUIHXr/KcxhiRv0xjFNwKqgSgoEGQb
1Xi0vEfLjm0Nj5mvOhViXvmR8Yn8LbUWjAcw28Ik3RXXH+IZsAfrsB1QrWrrhc1zR5VNck8ktMnc
C9uKoEbQ6jKxibbSSIKnku8XQVqAny990VG96b4O3ihnxguAcz7HEJGxV4eK8WGM9Mdq5QFsOipd
Q3JbppGJXSdAkWFoMXipAG6Xr5eiudgx+kZinIs+rpRXVx44jIVlAL9Uac/6IG6GXUae0/WGnhvz
p+RjukJqtuPP1N82y21WvzrduuiWxAvCLwH7aTb/49ph1eq/P2tKSsW3KmUn1m6oaGl1aHzCwVt0
ehACOsnrv5RTGgxg1wIabzS0P1PB5ksoJj5DmmAlN2kVfpUDU/65XZ4pwbkCmWZL5cTlonVlaWKh
SSMz7aliF/INYE1qruUf/VkJvrDcv8l5entwwrVSSizORMorNRrsakmByc9g0e46WF/pkH5FSJ6X
6Wg552mF4rjyDYX1KamoVoQr2XJ7Hr4Z49BI6HJwUM3kYQep7+YBC30cMjuYs+LCqGTCZuW0COQl
fZfgGPslHcJQVZp3gcbqbYBDl0BzQHtComKMx2uIdq7G4Ofk2vkN5NQopjxk5no+12HX8ZohgNvm
78njfBFArWFFWTRRyHpCpiH6/zHqQWxf9SagTCP7Bfzxp9bPkgldfaPjCiihpdiHbX96da9rb5lQ
W3jGoLBEy6K8zmj9oxy6gDzmRNjzypxWL/tVu46IcRB7yiKjTDh/2l5n9WPc7r3DVEXfcDVh/fiN
X3i+Omkt23YjV+U3XdFSTnQrpWUIuuiJiJEb+WNScMdjO9ZRc9yYehHaMZU3nMFhMjmuwvcUfH7I
I3JRqt1A6FVrSPcXMmlE5RNCGeKuFqeNiSwYgrHH+ORZEgyruO1h1CT9OwfUx/fTTq8OjwsDJcCp
9PTc6OUrtzF+fOyS4ktbRFhqIXDETLis7dFtuf7WLPU9K6dYahpLddbmngXxmjSHdSS60U67y6HM
dZypchBoEma8/IGUC50WOx9SoxwCr9GcR2MCVPKvLwDQV/GWLK5FMZTlp1g9k53mSC/WcMw82qgV
QU9a1UN/UWg2nzJBCiPz1pfJ00n/G0Sw+ROceLE63dG9h6/OiOKk0Gx8h7DsaN3z9TDVrvSa/whD
lqGqlQAn9GCrzCm5lt3kTJMaOjWNkcV1c7yKC/yad8L9PaRzU083n9H85n4e5s7w5WA15U2PtPxz
QDokwrobyIFnYL8nHkjpjfggaZhKP+uIvDPpyBEd/k4gHPiQ2YDpC54PoAGqRk3HiZ9Iii6j1yfZ
OWj+acIILFOoj76Rqdt1JMIaMdHwFJRQ6/u++eatLQ9Khxpg/g1xbeYw3vXz4LLPUOxr8+j1vcOH
SWh47Oc253j1JRDQyD686piyBci9aJQYtqWZXSSJkUCZrOA/L6VX15KvLHJfNP41LdQB8lmr0LYC
xZs2DSGDChLOrJbMjerrgQsmqufDjTIpecrhwPPcI/Q5AwXBoPx8tGP6zSg3MYEp8snAeEK02FLS
RB5gUtuB72TfguESWqi1FrW21GGpM4nucEZ/vUufTrygdrYDrZKEMIyXhU4B1qSZNtNdbJpGeNZn
h2bOGGcqnJ7eejjxA9RIo3lcnL6GzPjMv+MvAOYBVtnDmNgjK5J4p6bJZYtLDMY7YlIAR2hLLEsC
LTXZkNYnbtEcrgOhZ5ng+O0JhGM5k6Lq63uper+zbFRZB4FSafPZfsZylIYc2AQSyYf/SL0X1qbM
PCU9P/kq5HCCnNB2hmdIaSa3TPHoesTATOhABLrrqOPPTa5DcK395RsGJ48CCDSNnNIx+cyj3Z/p
fwJe2oQzCuDbTpTp6FusXjCHxWH4IgOfbPhi3MbYPAkunfvDxd97GxiA6beDj6fJhYTttJNaVq00
vdNjS+/dSw1VmX1y9pbbjJkJGITumCFnmKcvqGsIwiBRx7dp+uWP4PLitiANudY/suBf5p6hSCRl
b/ZKzkMXa+mF+iNsRg8mXhxi1v30JFRssxS8kbRd1ll6cXoeC+c68MvVEQPK6HsIzVmhDMuHvqgZ
dOgHvluy+1h1/pxfSVqtRSUAx107WaeMkiXdzf40yoQvg9y11YH4AdyvP/If2rswX/gMhsvLLeAK
hahjR5SkRjC7wnE62mCQdfV+cHPUATnINg3skn0dqQmJ+m82sY5XHyxTTYvX65SHeI23VdthpjHa
qyRYt9r8muPU0JIebnUgrV8vypzWp4wa9wTV3d/O4C2PfolALZxvxnixr5pJ6BroGzPENNvJ7rk6
8BQNrDjq8EbatRPGhz6FHHy7rF7J1OFINk2LQuGMB5KyxSjdwGorG1Cg2LMQYZ0fAjiKK79rWhxw
xZ5PlMUtIz1qVyY2cAun7vnGXxZQLLarQwRG0GRN52fVIq0X7EjjJ854PU98jW5QJwNxDqZfGmh4
3Lea72vjIbIOFHbQMZ2LVW74jBTiyCGKBTcPXrtAItFV8GDISlkjasu5Ne2QFmoX+OE5y7tUXnHI
3ws+imMgIQxT1JGm2klqTmh5QNiTpzo0HBmlf8Dq3jWnt4YdbeLt53+wrJQriKXmnQE7NfihYZkh
qaM0+dkdKc15vcN+dsHFDazpcSZKA9K2uzSkKo1AplIxFqiV+aRuU/RnyNuqCxwmG8Y4VBnLTS7t
/34G7NFELddEBPdUrRjHfIiaKpFqDw2HSXDUFUQs4ftSr1SAHX7l3gld6ZHFHYN6tbx2Cnpn2EK+
rTlEy+10IrGjVSLHK93A5kiP33sswl9cpMlrRqTzRmXZboRQAYXPHly2H3Pq4m3AgzxvgA5fX3bu
ZqelJgsHHtkGm7ZQWKLyJswr5OX8QhAjlCYBf00xiBm1TKxnKnmMUpbYYOeyWl4+NcUY76hNI/IL
rBiC1bz8fl/rlAVtfD8/ixgI3fwW0xIgDpmpbTuupE+TDBVpQ9qUigJyJRsH7MPBSfmBgyZd94/R
852Vz4R8y8yw4h/oQKxi4k1iVawewkbRz0Sh9H3ACKv0iaqK5iNjOSTCF/Gud2PmuT1X7jqsamNi
SHmX0lm7ROE7axbbi2whgqDFp1UcxUt6LXaqjTUlxUcpZH37/uqNOhlwy/l6wdbvET9KdGOFPGpl
3rQqEqpPa+Iq4ptcN6suR/X/xuJXNvvN2FnWnF37qdHopP13kJN222PxF1KhFgRxrJvQKVNEE4vB
fXdPQNCPJNrbSHRmEZ1W0aqWj/6T4Ivq9e0EY6uguT3e+RPe4lqTZcJ1yESKmaaqNSGSmK6nG0VZ
wM9n1lRbpHIpgMX3aePK2M4QyfF7u/u5m8upvu8RhbOHo8pK08L7ZU0uCLP2tyi7e9az1Vp4hmGE
fWzYkeIucjLWtbt4i3AP/U7MmEuSKLLzUYMpMeIoPMbej3ew4B68fMMAseKG/U+dlipeUITZlnUW
R1U7XY1TKcFHXw8DPqIsoylXXq98W1BmCvh0f8Hu+R8HofqP89UXZXIpRYN8g0lvXmSnh72eaARe
UrAumNS+gNfiHLL29FdcFuDzJShDw63f/+UGIDjVPV9J0pJaJBrypUWvqsHVy9CLp6OS2BMNAx7v
cbSg6/Fk0i867N3MjGImkLhfGp0xhckVf5BigwntUzxvYbTieZgaVdm3sOdJ/a4kY9vM3fNUBXn9
14p/cCpbS7i8wB9M5h2SYb/k9/JDl/8PWab9yUsNQEOk19S77FeZe3jZKXy2MfPc8jJ6f/tipVd6
LaLQAmFVa/M27nMs2iO5x0ZCOcnqu9UBuP3TaCpudooVcTzUoLQD1VkFQcWtZyNHF/Y0WaRW36mA
pcM/3Icv3n5DDEjymxFdy5PxD5rrFTPmOEsxqZBMaDP4mBXIwPCUHloJWsk8iSv62v+smgO5bFAj
zR+3ilQXHlZZyX59VEykZUL/cGD6PvH5Jjek5XxlMTmd108YaSOJRJlPj0sOMw1Q2HZo/aEwlUY6
rPTiwKIDEFl9kW774hlolppYv+uvXba6+oq/RfZqdNejc5uQkvEyqOgew30VDdMuHn0q/YiltOw9
kLYiTWQ49IMtn4w9U2LWCFcypinkFmNKJ7ODnPsdCsG7dNjwlT6sqhKEu6OFlyvHC64e0AiDMRq0
dvEtikdOtROFQNrOW1Fl77cvQvCAz6JluaApQvwOSMDb58V9nRZ1NwOwpBMTsAeX6vWVSKLPfdNo
ZwNU0YQE8ClGwoB7cLl8gImg0nt/rnXvnqw2rNQEcdtFIOzK1IzS6OiSI0ohWkroN13/5NJBg7Jk
gElG5v0lIokv5e1efTbx7REJsuOQnVK1IqzCVr/FLVnuZFq4jXJ1iX8kqBOolWSkL6mzjBFi+XjY
NmD5BX+d1pXAYujOXA6hAT4w4lFXdgRAea5uBfu6ucTTvvF0OSgwbgvU0BmLzo9bqyDguexN54mM
9kMpAM2vnRzrk0Tmi6wFO5KpufaEp2fHWmlmtUIVjL5yYTb+oPVgyQxhWLui/zQmgO1zwUQliq5W
frTJpxmynRY3nsx17xRYv+tu+yUSgHt/S23vQBLUa/VXfi6a1MHGCu0EnGNIn9nBc08CHjfZYcor
mBwQH+CBUhmtxnmCR5i+lpkOHv/tiQgz3JfwGgH+l0PlCHe0EZr0Gga1P4+xDgmAtuPmHrcq55mX
Uy4AZIYVkyROvuCDuF+/56vaf8I6B4Jy50UE/uLiG6fHZGJ8Hqa3y5bg0r32pEGsQZXCZOxgYa9S
blhsQqzMddERP4lFhTbxu8r18QMKoVybfMSRK2vTVDx0TaxoEG7eXSTSiKE+pw53Iq0+1LEbBP62
T2qPzTTHlW/GC/VW7cHqCF+stmQPQbQvnFpI0h6HW6imEiLsyftSJ6w8Lff2OGaWuLQdiWWvE7mu
supMtXikR+otbmDMluQCe0Rd+FIa67Xd+7+SnWHYQUlER2UhYgSzw4qu4SZtAKVcrG8X7+XX/qwj
Id67EUQVeY/D+LfhlVLf0DZMazQDjOjZNsdSIVjATpHgwSkl4ci27YF08MOWuP68EbZoWrmsDTG/
5RN6iuYtkhLWe2tqLOkObakKLmoDbcqbY9A5HxNTvoDXURdhLmG2Mqam4Y76/YTCBM9VoQV7iu5W
Xju6O5rCkxaK+TDirogLRU4ilZavH1O/ScBVixLpvIccb6CMVPq3HR4hd1BrL5s/kC3EonUOTWm8
zh4JbO2vc3bsTRiuE0RullP+7GrM7Jb5J16K7pDPv4Zosiz0WnTPDzlJtEhf/gHAwOn9DLkPRAhM
rhm45m+kBsPYCx/0xUis95bNkePJ4MU25op8mVSp3OnyHAEakajcayBVGUyRKUl5nfHlITogKxs3
8LIg+hv9uRruhOL9/Qhz/7cAMr+bP4gvKPyH5cdyqJgbAkjkP44E3vQhgyY/hd3ggw0x2ynlfBkz
Dsaarv+lg3wHCNdFfKmCz26Z8HWIcS3HSCE5Hq2BmsjfIuTiFVPW6BRfMXlkvTfx1BgExUQ2mAoh
3Rrd62myTF44gbGAOezSINz+viJanLlg1hU81eZVdZAmyUB62Wp3J1NDNSb1rwizOp54SXCx7Hpy
CoS/72tM0yf7DfBHkqnPh8obMZl7QmLqoQbOVR4T4lg07PTwloWR91nmCnUDoi9OWR9txSXWcMt3
fauSoYlYQDO8AELf+cevNnbOLRYgVXQrMZlo2t2UIvU0dhNlWZHKVucEO2Ernl6O000yp8aiOUId
2bNui1Tn46M+kM1+qnFOs5bdZkxYq/meZHqVUnxuEidjWaX0HKgaKGFeJmusKj5ikTkKOimBnwOY
DspN1ElZx4S2B8exO7SDJZl/kqbH+8Z4E5dN4vuRFhXn9uZLiFWuZshEm9moivak55FqXAFqFYW/
Y7k2cYSGSb0BkUPwqNI9Pc2WAeHtkWpfPcZwJ/0ucJusTwvciUld4SYAvcAue4mbgEztD57M6b2b
vOoSnqjACZ8c6YYDFwYIUekmSHuM7sRnDeLe5T6bpZGF6rryz4VHE2r77k+8F4wOd9nZtMVUy8aM
2OKy57S5t1EIHVQW738g17Rsfw8aqG4O9u/08fZByAaXP3ApT2D+it3LQGeBVbjE92hcD0+k86qv
tFFRkv5VkOoI/SUzRPQDIg1EDnQZlXyav5NdrN6bfmKsgD14i6cFsAbq/iYOUGYDkeZBUsBrr5b4
ISgCk9P0hdyIdrGfMefuAQmWFOG8LhOcjZWdsWxdmm/VPO0a8MjMHYtDB4iYW1NbFoAYETX0ic0Q
LvYOeDH+B8V5dJbQ4wjuz2W/XKIvyPb3JEHOjMAs77s/8xMSzYXFQG0RHrrV9wj/SryzyfcMEUGV
q4ClD8ufilI3G3ADer4J4j1Le6/KlZL2GsDDV/PHC9LBjAHS4+uT77tjdFALmwyJX5aw+cIoR5bw
aCm15SKn0vQIsbSjRdJhSb+0+qUN2BgyAwX3y+ya5GTDQAf7BC5HobIQNRtGZKphN24fGPCNg+4N
0DTy9bYtD81qLAlCACZjKSLP6Yw6NPUWTs5bURn9KYvUSwkPnO4HE5YnSEgAyLY99GKMFNCFM/B8
FYe/LUMl1OyK9aPdVQNr9N8AaOk7QR7X9b5CzMKWP8HxGbu0se3tN4qTCc9Z20ToQVC3hKfKMlB6
XhD0XXxRRhtzt/ayyXVA/Scf08mBFnG6qyn4NIadcRUsjtJoQsrEPjQ3xWZVkTYbjdhRNZXwuDX2
wvwX05LtJQS/qgSBWomQTr7wuceiDegYKu4dBl8ld7N4XrQ1+33UIYPzelJzgm3UQZt6zs/BR76E
7YlU9hbLIJTmSOPjgNUOOPQFtyw2wPcIKIajHe5zvJAIlTZJIHCXqGF42beNFHRsxTPDJumWIGr9
VI0XER5WML2E/yYGArYPvG7mZmmKXGkhroraNINqJsudm/AdH68yOAbey4/m5sknaHxtpwcKyTX9
6Y2ILlPWwiLoYbF/eRSNBsnE8KBUGyzOsZgJOtL9fHrMNcessVhEbEU8XFdrRjvttNiA1RS8VOyA
j2DWmnLQdje75p7IvaBZhOAT1y0m+UvZVN5x3XJzxhSR5aHHxWIh7OteqDEbIDOge3Phs/ijk3Rw
VhtkkqJk2FC7q/FO+5lWIg+GmmaPo/vYS4k6EOynDHLWgTpdsB0TSu+X77fotXtWRZqGTrURk1Tj
iO7pXnq0H21VZ0FRGWO+82S80vavuy8MtAi/PlCyP8m4ttLkhTC7YegeQoGQN2/FqPmAaEzRjHX1
BHN4u+Sz1HsHQfbw55XrBN5qGWwYjnCJ6U12sd1mAAUM9BrQH3QyywzBVPBO72pUTESbPRVntRnv
vYXxEwD+EtZvvde1nx4eAMNQ87vMbqJQOLRnje//Sm/auuD0LkM3vzypXsyhQkFPDzSKZ4I27Xds
VT2F0dG3s6v+AkHgGrvlpUCvmyd3sX8Eb4cggKkEJu5qG+GH+VtlsMb1MpLK603LIecvkOuGNF7R
zUlLEEKfVbbynl9LkSsFS2/+63whM1IHlv5ZISPlJbXEZ8rtcDGYEtk3vyIlf6uKwJ7GjE6xpDV1
wl6hp00gcj3WnSW81F24OgdetkNDl6ByoQMwPcyEPZKkniVY3fMULC0JHt8O3pWPOk1Rfutnp65v
ETuxUuivMFFjLQwTb26GnNwh9E1t8/CAlghKva3Rnnd6PTodH33iajF3aDAnfcYQS26pBE5tWsfV
73LnP5RjTfhAAJ/FR5V+lWPzqzUI7T3Ud2utBc9H6ObFTCNTkiQSEPQKfipP5BQk1UZJMqUBt/x5
kq+xjC9wAWBXS+ZNrRBl7Nefn/F8rt80PeS1K6GkM/PEP3xbtx1Dp62BxJyetbL/FGxZH086MgpD
HG6pGld0swUd88SpjMTEVnOyQddSwy9D8skrY3ldDaVVj2qXx9iXe5HhIx7JXhA4+HQrN0uK/dGJ
fqTG2NmgCdwGTRgMGjTnl/P1tS8rjj1/BMhE1Vijw7Ze3OFskQyp3yZ8FUXSC/cMUzxGgfNmmP5L
u866BLJvdgAmCQ/JolmFjIpMIC1U/ShPrFkzREzZWiVrwn9UuAhQK4l5PS+0QG1QyLK/F7wBh5Rx
UmIDWG3poirFWLGVLsfb3+DDvutG+AR7lA0jNlLsakn1q8Rr4XLLtDZ+9Ko4C59LjNkxdDSQyYxt
A6I6PCWngC943knr4eA9c7Yrgk7bPbwlBAD09CBSFOwHXN1A3p6jOY5txwaNgJ25BdSVbvjLCV9/
fPDV2CR3515oHuqkVsjBjyhjS7uucNKj7LD3JtnncXqE2hWUhvPI7idiVOre5KALljniQct5Hiki
/GMX94KkyGbg0y8o9GOEgz5vYbe0Lg7IH3AziEK4IfatAPMVVTGxaaCN3MeB2GlXTZREAtbUZ9Ly
T72EGgpFNmaH8PAsLl96otVsxWZUucSvYTorq3TqcFQZgtywfO2YoWELTdw4/+ZwFoVH5I6GxGXi
tNJwJ47nY6oChIRer+jkmnFsmBxI7ytNah3Q1GdK8SHFDdwkWAHtiSmBGc0YOSkl0qM3kgtU7AKq
U11ng0/vXrjfGDF8dkEMYiO5+nZ89vDkiIsgP6+Ci69O4w/LLp8a4M2Bf1usaS8PufhhXAfUH13z
pFmBnMf1mGTYoByamWAd/fHZfggvPylHD97hNOximbgvHCRK82hYCHVsuUitiW+F2Ufp7/J1eXX+
Jk0hR3uyTTEcF8C9p7gie5xZAXa2SGutkl+teFRyLWku3S4hEVEq+LGw37f06XF0RzLfWl4+GbyJ
TT46pO57KXEYkkhUbHYulsZtjTotcZqIA3J7nmp3gkS5m39QLRp+UR5K2J8GuOiCoVgsLhzgZApQ
g4M8nAtdx+FU5XmxRZ97RZyBVZrskwIReYF3jqC8fgCtiYThj1bsVB6D7MTfJoWFZ+0PZJ1R/3oB
RA0CnAymy7rj5DFANGcaAwUedIUpVTlPY4voGYUpwnADjieINlqTeqTyH4T8Mb+CB8g+5oHCZCp1
zMh377XgkDk5VoTxMYVR0djrvY09vVkOXHOXTRnGr22PNyXhsV3x7dYStP2Wf3PtRROINBOjnIlx
hlxusFIlmL2I8vCwqor/VopkasxBg2HzElSGaoNzo8hDmtuEjdlr190+96wZFAMTKjCu5c/nWIjn
KrYCW7gLfeCNb6WC3oIpmmqi3jafZcwWT75sbpoiVoJzt36b7xlVVxBKpPY4r/ZyNkibjmleXgXI
y4gTWR9WuuBe7ihSyUXFrkzMK+u7mm2I0CI2pim8ZvMxFHInoPF56KnXTKD6whwsZaUeHI7IJMye
n1Ic3w3DudayzAsd6ZhmR0sBSqHOSTf9VrXi0JoMisBtCV4udGOW7i9kOX3hluXDQhYIzW+zn+CT
vgkh2ZMVs27N9RYNrwy2enK+/kCYjW6os1vQS+AgU8UxeTVe73FGTZ0idMGrXyNClyP7Ew1xLY29
VdDjE7uaHbCMHf8xv61l8dUU8seIR501RWSXo9fY3xP7JRTcG2RKR6Khj2vlzvVKj8mlkYsf0cN7
hh9C+AWHKavKUDWlDqH7HgbOvpC5xqsQa/dfy60EfZM6kYFAcm+/YZ9XZN0fCmniglXvbUus7n88
t4Qg4HExhKPiw4XWmNPjQxM/mnJJmsYZoNq03m9lDq3KngRkq1/17SGac3u+qV/fC/CoeAblIbZU
PMKJKqBdZVD5h0jUdu+TM7W2qljjoW2d1BcYsl4RPhi1QDvdlGA5op4DojEP4/63PW6F0hhODGNM
3fZOyUbqLN0Udmqwo62JOqSs/4Ngklrv08Qyd19KME/XjL2qftlKmlpET6U3473Q/p7Wu4HQcbo9
nICkgYZn6KYk/q72px7Vj5w7V9uD6EXszCDDE5IZBIjJs4VEC/rfDL0l7NPzua9eBDswNfHITmrt
xDRv7RwD/PcZiIvMDFwUuApQMv4T9cHjR0UoycHfHaF5r00KrAezvOmSabKYYFz44r1q5dKyY2mI
h1Zr/CILlFwq5qI7p3Fz25yUYoj0oCDo5FKHphMlDvz2gbOjwRaXf8Z11gKxuiNKXOSwNcg7HOjs
yumdytOBBULwVR8gFS53Vl1R36uW/IjoqiBI4+alP7zKanC0yWmQ7Y77FQ/zmarnj9zdlkdYNMYu
plXCxC5vAaY5aV+LAUO+0/eoK8AYvWuDEgC5XNYvPGQIG5E+VB1nFZnG40q47xTUA1NNSVPWQA/6
yQmabMpkyNGcKk+OM6DNeMHcyD4zD3BP+y8EBDBUSCQPEVlENTBQaSL3upRWu6DO9NGOtACbE8FN
kpMPMVE55R75GSaOMfjyZ7cD4pvxe4KOhg3wuZEhC0Qg7gsZUqd/f2WcxYi+SZqP8vYrXNRDbNo9
N+ORsIuWutaZ0G3SwcJY5dr8Wf+nWA4BuZZeehv4PhDyj7UfM0pcPea2h/XFURo+2VtuOQPkk+vE
24tmdkxgegQ7PdHO8a5Bve68HHLZLunJGrWrYK10gvECTGRsajNU299oX13ft2I5j5A42IWY7+at
voo68Gw316Y67Ze1Fhw+5BDTMv5qJfl1vK6pVnqMauEzDmZqrwM8xOYx6lZVRYA6AMUgxAyM76j0
DTZmS3JNZeXAr7kTfGblnZJzbBLjwqs2fS+6lQv1V/eI8NujQqsW64S1DT1KRI+eICjuUaokv0xf
qMjXTbP433OZEwhfXHmTmHOYSgCMazESLESHrLshpApfWXOX3C8M7Xsa8L8VC4eaHLKx80MB4tL4
IwzoZH1oau8GzF7B/PuHGVZQb2tWVwp3bq23LOJh/ztsVPskPc2lfsAykUXPCAYQIfIPqfR6LktN
XR1fsLB2DUoiPGyyyB+ECKaKxl0gthAyGptrKfw4dIqbGSIluTuNDk0Dtr68ipQD2IIgjmFqXJvK
7EgGewiT2E3ItZq6NcFNq+PmDXMcrKWI72xQO6ZrxPggRwm5UO+1magTwIRezZO1SygYxfQhF+q1
ShHGmGw62c5py8kxaOT8gAVnWjcnvmaAkiVWxTTcaEzMFrKS8AgsaClsECs9wPkkyzBf8yaZzXNH
H+OIegiR04e63TqBUAzyOF2mTbVsZJybs/GjWqr0a7WzKsTaVmNYSEM+y/Qem/zaG7LLqREi2opi
FDkIJgtLGtYlMsKrE8iFE40eHIdKquBLtElXwsNUeKYe8N1axVmg+3d+KdrMudLIKyZWE84BOBLw
VwKdbaf44GBznJzEYGMcNEDOtolLmyPV+WkDYeF0XKVR8139QYthIbDDiWDn2UincWyUv6z0vkkX
W9PAyWmfSeYjXzRsIGclN2dmOm5Tovqpka8d8/x2TyvD/B3Ycdx4Wh30u5ZZsFkTb8lgdibSgBi5
C5688nm1t6cVsTC1kcnLbQQZ562g1jwtrAYXjUUixdN1PPRzZeLALbr3IxjC0TcRjWsFd1gDhX8N
tBEbngF74VU8EZ46XBXJKttlYtmlFdQ79+BZ0+wyxjoY1/FNHaP3tAJHytRGSyIBxQvd9D/jAWBs
JGq5q5Mb9rQ1BWVG24yDKUebOnV0X1MGA7oA128cyCOdBjdw2ihHBKFzck1qkKfCTeGrJghe0z2v
2HKqY1P7Y9H73uu6AqvE6Mik90x9h9Iyuu9x0wyt4rwjmcZ6brGQH4osJlR9sQpYWCLlRwlfUdsG
j8Ggaqo822iR0FzK8Rf/Goew7+aGwxO+h9jjYsDUGN8TC3o8e8NkL4ji9MHVTtyWxEFQ4QaYfRzv
Edxu3kvMEIEmE3ANLGoMVmEP2K/6QhUQpuQyJk3S0CrE49NoXIgXYmm2sYGh6WRsxofb5OC3QgPb
ZvuObcpsaW457HdWDX1CQJ5GbZOLIY+f/rThB7B7bpNeXyAUDc1fgahKQcWGSZgBQLV87dxBTM11
14zrEMkrr1YKbbEkpTrTal7gVsA97KlgO7a7AB4+vmxMCguLQZ7LHzuD5gwR1gvhkH+Ui+rVxVZX
L6bZ/0mBenj7GQzm2YNMbokWWnYX9rzjf2hWoiB7wjL3G9eLbIJfD0Sr5cYD51syBV79gg67XNtB
jibuF5Twi+KcrQZGqB9C5Xouy0x09KP7mkTAPlc1MVP2UZhDi3DsA4tIl9dUXbV0wdfrdxmghX/9
7CWd1Zzm7m3nmnN9I4dUAUutalY8VbmMCwPpsv4HSgGkNB9/xpugqNu4rAWd9ueqz4TfddlzX4pU
WbgrDYxk1zAzjRXuxqHEuza69l188FbLZmuzevK21SSNH/O8EAnhfU0Ka0uqQah+V44hzkAdHjXb
mbbKHWyrF6H8cxvBN7B+lazM6fZ9SuzTs1PGF9OyJaLDdu3JN6wehET7nfxASDgSEDTOYVRi/eLx
NiO1Vo1wOnwTQbV5RaqZQXGz7kQ8IkG+qsjcPSsnFRZ8OCHgHRS2ZrMt7rQ0lZI4L0+cF1sXShYB
io6pavuZdY+SpxWyxEAA70Tr68g0/k1JhfjVeJnKxAwfEMxakoC7vbPaTaola/V7SA1xsiHqZTcZ
jUiUmewR8RyUEo4JBUTObfHQgeJKJ6F0aKkfisN7qauyNgVhqxZ3QYyExMqbu8H0yD3xASp7DmSE
bDzlJVRyz7JZzvAWvRiTBJ+ZYRkE6jXGNtoa0DI9oI4c1B3fg+YuVedu0xi0L6/RSgFaN9go7zn1
ZQsJY9opLfdz9ihdAfsKYTW0BFpuzVmj7sSVNAa2Xfm/BhgM1oPi6Qz6feZnaTUdL/Gv1hQzJn/X
wiAxWLPcpiYEs9IH0RjVdQfE0HzarXT3cUoHAJrF94kvaltLNfWy2UHocE5teQ6r1MemZT38IIg0
vq2+v4UBy9VcYcUwCA+CTnf2/Am8WbEjsLNIkhz+cUR1aug9nZ9BZmX5y/vwfmTgMATaJ3VjIwp8
7Tc43diJTr5/iToOQAJpvs2dzVRsTy8QZ2E1h7Fiyctwyd8oWfjjB8A19brXr6tUO6FAOhEGKvTn
OKY/3assBrfK01AoQPBxOfj9ePLc16G14d30wrSqBpQyrndDUA8wcLkz7bW4BkaBza5MVf14JM6H
SG5n72LU1AM3SCVMoXys27WoRu8V9s9+GMgJPBdG/EWz8jJjGx8m8QL0ueR1I4GLN/iJdKI3dNpg
q9eJSpcS19KsFMp0o9HLrvHDcFnOHWVQdVVl6vN/RjEJ0JEtZD2lnOkUwvfsA3hKXkjcFBkQLQfn
ZNC7tWN+5k5636Ru/A0Tw/h4wmv6hBMNG37jqJ/59JuSqzvB1woFW7gXBMhlKeOkETraaDczYQBr
5HZKYW8Bqo5UEVAK14BWqoOV05yBwMxRIMThKUvsQrtogEogxA/7MI+65C8ZYnP+ifm8X0ciV4Z0
5TACGX4jZ9jJYyu5vG/vveETseoT7oFUPlnWKiH802U3nvDertAmff2MpnspN1pVXMQMtNS7VKLn
zCfA1Mq3fXXZUPWP9AjBt/zCdCTUMjwm7M+2I4oDt5Qr0yhlAhLIBv4q47T9Gzh+ZgMZ2SOEmvuA
lDUaJpIhLvah6lvvY0hXi5gLk+HrnETB+eW5gfEnSEOKjiVQbFQizX9xc6E/bVP2n+w35S4vjvx+
zc4FB3/7zwoAg1pbbinlpVYt7oQo06YUj9Xjm4Y3PcPrHlrke7ctVjk6Hs4Z1cfUfqyhgm9Z2dk5
RRHsmfHNyskFIaL2IELpvtMd5Z/QzTWZjybmnhs0h9QdHN7ftJGzMWpRxmKo/SKPiOejV2LkNU03
Uj2pOtHcUV0yCxoup/+TYGeOXqraqhg5aQFTm2ZW9hLHzIBrSIFZDtm4q2GODYGpB5ukJlc+5dzt
fETJ6zW3Ij2JQIgOEw13XfexD0QaZYH27xSuL3k+C0lfkqbTtXhArikPtFCR7KcOHYmky4j5aKax
npI/W66I/zlwrR/wK6OIH5qR4KxSaSJLooqxZnUrzZzWfkxS9RDmHKPl70uc9KXO+NFqc1EBpqFG
/ttTSzO+Y6zHpsVCPpC5qComexPsFXb6LZlkWztHFvG++PZSqbzKeSIwQhV3xZFnpEYh3fSZvHR/
hckd+4bnpaNmFdbQ2wrUri+tuGn0YWDH7xLlvfEBSMNgLfBN28lO7TQxDGcXIi53K1GxuLgUrS3Z
Iarxx0QQ8uxxUdFwGbayp8OLv4lRkkWogycdXDanV8+Ic2xgdzZdTQoYt2rsobqrxszPpU6SkG/E
tbsvj9bRrEd8oGOkCe69aRCp5RwtWF1J2DN8j6vm0N1MlsQAzfy0+4ezQ/16SvkOogKOFETQMbrH
reYy6KQ4sfPfsnPBlG9j/07ByYJLDqDz0TaWwU5KLJEw5l69GRugXTUBS/ERB0y+DkwuCxzcUBLo
lZkuyZSHgtP5ne/UtfCgKPPi9qWdQc75UAn/MuiQHGXN1EhmnPhPHGQEax1uvQFYp+knrQQWBAHf
NlldsDyqppMSqykAprxn4GUZ4Bxn2m9mQi23LgI4sUjrCDhD4/zkVHBoR7vzT7Xz3kvOC7ieCecf
fTiGHS0J3duC+98UOxltAngx0RPBFm+05zL3g0m5BT+ki0Gq877q5JR+wF2IpE6Qg1e/5GANpwv9
XpJ1ZqKmlBNCsoE7oKn7MuyjD1Ku0lu/Jk6/OIPhYDhf0zvf+lYenmz0j7tLnQV2R9VCtDrb7JG2
XR9kZ3tuYCbmL38JoVky5cVVeLHJ/5dZSmKbpIpCMXGxlNHg+5G3NfOMuvhKoPUv284FYiQnwEN7
gxuRHlOU9hOCjSfXHyY1+bchCI19kC4H/sQQPkp944r92jdDzLtsXto6nLNaQupFKEkehVg8tJS5
sxnWHDusQwFpxkvybfkX+6HXvjCSvbLoQqKkSwOSjOkNLPiSMsctqdSa8VQPy65G+R5kavqYqlcb
zxlPfYEEUGtuwhZBlaoFxeB3MkOMtGii67HfOaSzYoS83F0Xzd6sbHuWd9vBZU5Am6BJPpsARU6i
pbwFnj9PxjPXuwFlbU4V9EoaVDcBiVQwhzYQszVqVuGJxgwfjynOUE3uXXiEhN1KoExx8+WQQMLm
oWY501D6poYG52Spm2JYn82CM8tGjzq2yyfYdMQX/AKkb1ZY3zjhgsTJNvqXKem21dtlE0xkI7v9
8oDN4pwDpVCu+QWcqTiS9hOc4YefLmsawQfk7bTArloDhyngD5lMl+2bjv1eP/OLBmLuJ+dzHm4A
fLEvtuc+/iQMPJrsg2YTgRDK7+1Tri+CeOdpHvEjfTjK29eQK5l/Q6gRlZN6nTbBYy/8+u27pJjz
OyLMHL4+fXfCcG0k8Av9XonsX0KQf9H4U1veE/5QanAGV4ITgG4vzOSZfP58c6lSjUVIPig2h3mA
aH2VYTwuqs1mnmzoLOSZsjruTfIDEpk44phzegU06f4phKNB9W3GqbasCK4Zu62gCOHHHDYmyGYO
AaYLwBPeku59OOJ3dgT3sB1seo2s7Mn7auOBoUlGH2Jv8qvvvj6jJ6cl7TyYo/zsxCZ8n4hdcxjl
wAha3onNOfNfHS7dkrSOsCuj7zxscz6pmN77oLdmmeEy7bXdMH1SsRJ22oNgvMRyAiOX/OxbJ46n
lQowp6rKXDUS+xlMYhtIE91Cyap2/YzzyIdgEOUWInJB4eIIlw8XzEHApxgVsLHOla6E5fvzBLE5
ndz8hgKdOsDNGdMudvaCJrunNKZAiFvwVcj7Tn2sYFfARoYwK5hvsudq0sGpTkhG/p/4AsIk3POv
o5FIOTbgs+mgld96QwtKD17u5UDd29ieiTrHBgyY0QUzphzN3g/zn9ZeysUG6e/qYYVio6Jlf9bm
zHWEwZ4iQpAkaB2noAMRnLr5+uePV0FZPwxB5/H7sW0jdOp0kcL63BCym33cS/MRaz2Hw6fTr6Xz
uKzTTQ3PQPRjz5FjfodRikuh53j9z95rD4bfKvPLsnKjmBgdeotDMYoUtM+dc7EWSt55wMOfkl9l
Tt4qZ6QFPVKxSIEyPKhuHpebRiUSc9BLiH3lx9VBSwWMRERJfmIdE9qljwJ4zeyiduQIoRBxRf7J
YK8GLYeUMOQHMGzkTnBdA175xaw7MRMuRGTdZuR1wT5zbVwJcpZXYJiesL2cLB/y7CZCAdRuGwIx
BM/Q6sBAG7bY8opg0UcQxqlYHj+SaxMvc20m2o9M3UEjsA2MfVZrjrjLv4hVnF6ztm8UxdMq0yNn
vJwPIm7uvGLIS5iOcafrcITJD8UGP9/y5F0xDTIi2wjGLo4AIMjq4rfgtyWIHq5LYn6zAaGw2CnB
nxXgw+6WkeRJ1unVkaYrnXdvrc8fVSmwpXz2f2/qaGd66cN57cHsApRdESXZZhWMEuQucP+EBwYl
kI3axN37R0lIfIUmtSLf+xUfliSkJcWS4qp0rwZywgGn2GklR6gkI68z8A8iAhI2Q2kXlLhqeRyT
hM3GC3cr2zMYYaShDGha6eZPjYK9om8pLe4qJfOt1Z37RzVJLHWB0uRHF5gzw6h3aAh0ZTVRoqAM
6JsZ0SpI1uwFojJ7mO/gBxR7RHPBdDf4Yb+LpocfbdY1CWtJMzrqcQUzOqUpZzkfkq+WMtVa33lb
+CvKllowY6nHNz29JrRlefg+GFc1wQ4bibha9hqs555HfBbdZxgd+hL+USgoELlt/HzppyLmAgrS
+pTE5Fx8Q4IswZhIkFa2mG3ix+n/PAgzTjd0RIPmWUgceqrH19KWGLA6oIPYQpShKMCoCAuF2WVm
mGmAgCEPmmURQuC5Y7iDJ4JqXjf50sBGpziVWtJgYgQoN2O+6ek6yvu4eX45PVn3yVmbYw0Yc8li
XunsLnkyKrWg2v2TIb+/qZFh0rec7qo3V0H8zBn7zNIN5VxYpwv9bbUGebbMOEmQ9CL0Fn5eAhvH
tWJMJRt3lHJljOszy2L9I5LAP2EmExyZgOCD1tmt/e2SnYcyZsps3C/Fv8qXE649nYHUdeSP1Ywh
eh8WqRDS3wKTI7aZmLbKaU1xL8uppkzOV9iHQo5y91cMXXlTco3o1rJMbR/ZWHVoe5IXDQizglxz
dILing25QPhjYkxW0BhaPIFlD3lFgXFUc66VhyJfCSefGHg/ozym5agNQSync9xxzdeh5mNcLhMR
Skkh45zF3I06rOi8KFABN55pVDfzhQGiLQOGUjQXOFf70hdWc+xRicJcqqmpmoKmByYvPVvXsxu7
pLj8VGkJRp8wpaLf4Q8rZ8rtes3a7lYIQIUFM390B3BkudQFtaNIuNPyD+zCNFK78aVWvVhjrnTZ
Mrsrl3Q+5EumXfWkbcTwNn1v9qy6/GV5zBX7Yl+Mc7HuWwnUO/resm4s0VhinEDI39RafuBZz+9a
l5Ret5RJWR8j8VISBhHWiB0d7eTycV9PEB/ggSIdfEkS8Whv0nH8HgUy0DaSoeUZCYKFTRvd4kdc
QUblylRXQrUDfYrpHpu4ru0zwFRVfFPgIKy+Pco2CBGPkk2o/c4mnoPmdvhplrF8RbSgKikQ2w8A
DY2tD6S3sfph+y0LEGA8THUd+VDAZiUYEEAIg36sD1MPOSNc8VqpEaQTMXNI1hP93r/Ob+OsSYrv
HGzu1t5yM20zDOFEhWLPywyOFYj+FnxzbG6sVX1Jpvfu3MMBWZmaAvYmn3h8c5ewkarQlSzCplOK
qM1M3z/m968qiktcdkWWVCpsT7ALr35wKilJPqdNHjwDo8cEhhQvSLi/UiKOyEhvYW3ugQdAfPKN
uWdJZJfJx5EsLP/BKOUzEa8touvQThhy0gTFPYa10ZPEASx5zHf2p1n6k0uRbbg5g4jcsa61KvRB
wQJeTto/rtztxlTit/UD8tg+9/3ejJBJd94VcL87PxL5L4OP2eQrcmt93hPaJE9AQblGLT9mQgcq
EtgiVmu+4+v7NFEIm8YspU0cPdJabj1QQjdiXRv96WXDhLe2fpqOR/NDKKETaCqHRFZiL62RMFYD
8p+bbbdrCzOfndEbBDdLwj1hC1MFw4k9GYRc3SMh/HRJR/SUZBlx/VJXPA5RicZ/p+E7rD/ANxfX
6TuJ4pWiiqKC0qWUXHxk7X/22uWp8/f1NqCtsySxL/V08oholDAAr6i7Lmz5aqRx5Kjyf61pn1eG
GOvfdYCk5cRHNAT6M+3GH0r2ArX22IKqWsHZ5tBp3d/iIJG4B69fRVbBj9pqMBzDpv0QPIbB0ebj
EnUSc67jLxz+kQeDbtfcQhFrDY7ZmJ7ny0LwykKZ7A17Kt7C0nF3zM5Tx+0VVw/21CiWwHCCTYTu
dKndEPnI9QyZZNY7ZR2qm7gJTiFk8aZBAl4zPuGLi9TbMaH4H2j6hoajo+7mjD0rHrUUdwrYdGvK
3l+DU1UNrrP/oEsjv3M4IFNViDgUQoUA0givKm9cLDc/YUt8SCIT/914B51YcF+EF7ZxzK2XEemv
J/Ty6QKKoKl/VTWSA6wyKpeOPn3QBVwbx+IsRrVUA3yhIxkgyEKQiE+0p3bqVoAKPKvNbL5N+w2k
2sFwuINtiXLST809q3ffxOlUyKnzsYadVBo2u81CqZ3fq9PUN+ukj+7KmWW2GYwj+JJ5019391NT
K3jJAXaMj7FlzSsXoFwKboA5i1uszWnLsP45lTipY/D3UXHoCDgcqRSY4xqISRFFVu52+WMhEzKs
SsvW3EE19FgG/5HbQ00jaYjt25PfKycR1EmWIDvQimqpCBHBspixWreniMGhRvQKQZqmZNE9xCzR
yiqLsiz2kbOoIFXnxRhmQ6X3JI4BYgoU9sJAFOXiBtahU4wKSKwmr92EDPXvtqG5cI1qVi64/1I0
RSuuU691sd5ok13cbjODliRd0pJSNtLgzgs8LFQCabkx1IF9erkBMkxf6vDJJjmEf3C0U6fFqT2+
CuJrL055zWrWZNapP0SHQB1F8TcMPU2mxpRbSc3PYWiXFq8iZIpVTCRttyZXWi+FFexGA5/+1fwC
LeYhSlMUVfMYEtXg8rv8TWcW5Fn4Yfs+I8OdqxuEnfAI4Cx1T1go140Rcx3q8DzcNIOdaIpO2Tuu
4YqvEKvzishehJnm3RjNf9X+rK2X1FT9J3Pg0+Ka5UtE29jYih4Hpvd43T6njOkTy+lFaPUefPcF
tiRFSziq0MF5N+28OVpyzST8oc3oHSw5fvZ2+RVoJudnW5amm1B34KfNOnLnegHkMilyObcWdGVo
afQTmaiFvHsVQ7tcNYCcmebdhse9YXesptEPMA/OSOIOIPqYXCj1ajafH9eiPW00pksMAVjaJicf
4npUN0kZwWSh9ekM8jMRzsnRaiCB7yEmXPc6GPlzIHwHRzPogLuE7d3usaT2aivXXxFv742RoKMQ
X0LY4vGNqVkwxmpZyzo12CiIegABnUJYCrHyY6OyHE3sRD7ZEw6tFMxtln+rahncqbB7qWjaailp
rWWgqVcuziopJxgfFTHDW33QMzJKWxc+HRf79mMSp3fgEmYBFPiuOYYArW9XOfsmw24z1CmES/zL
I9DjUwa5Sk5hHCbIjYUV1nA59hMS6xnLABBYcHRgDi5m1X8tBnPrAGw7l8HFGvTumifevWSxCIWd
91ySHyJumTtylhPwUuRX4sY4XpT22uQa0tl5MLTDSLm/As3LPvDcgerSLnxiPVoUNuN7JiEMS44s
pB/UfvIjJavm5tkYhcxTSdzSLqf2O8EdA2CXbYn93Uxw8b3rdGJv+JCcHrcHoJiu2nba/Tq8E2vN
pBeoxBIAxWEXxDMs9tU8OuGw7aS+hCcKpR57r94Anug2zM0zjQoocRspO5tTqbA9RSFnx/YD0+hA
3GlpsZoXyd44jXGelcovDPsv6d5hv+Lhgf9TNKX04Q5Hu/KUKRTVVBb0DJXTFWSZybz174/q3sGm
gkGyRlZE/xoR911QC/H9Ho/0hmQY5h/ln4Fr20dg6UmAyYADx0AqFIrAIvN4AaLyj8fzfZXlM7OS
HZuuEYEwhX3mViSN24EF/0Vt0W+UjYNIchZ+oIOM1RHp9Rpo1LJs+FC6qD0WAqTOVVopZ5CiMvJK
iqTLoVq+K+G8cCG69IUOptQRxljBEvpRvJvhgvrbSwjBseXTMmjcu4TE8uQJDrK7X29s7YmPB4E3
T4DBzJv3ovOrNtfnVnS0Sysnl0QqM8POn04PPuzsOHUv8HRA7WuI3NW9KWBekRzhWeWkOJZF+WrO
UtlZ0r0gxvtYNMgHM4mmcI7ARcC5L8bctLtJMiL8eEovZGGXQjjnd+vyPLlUJ4DUbjTVGCq3KQz7
oxzmE4mOGe1QJJZbuxMjhJcMT5BjTBRQ1Q/E+ru90/NU6p+a00Qixm6ZI+42U+6O2SlklBhn8gBQ
xzgA3Y0Lm35sMTntuB0RoXa23ON005rrPtHZxCusHp40hwbNi93sZqwRAfBEajSOP1y796ew+tXK
8esUwvChuVrFic2HSNkyCA3875Xxre8wMClzJZ253dOqLibSJa/DnKkcm/Zpwg0sSxkRdvFkubBw
x1Amvk/4mb3MTdDrq0YU5PJM3ZsQ2KNFzPsGcuFt7yY4yYxEuQDCvTA9QwkmZ8JMB62A3FpWP6Pw
j8uv6f0eN+zn3aVTHGHNB0ot55y0ZNcvRUvPCabZsYSdPO+osTKCb87WdN5/nZyNF/I+U3ZHJVVK
qyAxhAqT/8BAy/oiW+rQ+ImUD2xmzKNo3VyXqSxryKCAkSaGn7VYQGcXXZMw/Bzos4JInHSQ5dOU
DmYskwPRHiXE4VcvcnEiVd0hHtmWJGTAf+l1+WY8kgEhlo12bd55/tERyo7NHL4nq1o+Cb5OVsag
vETxmLMSR1JW+HeQjnUWCLUkqSwPywh0ZfhINUjgRQGfPfza7JYFtmVEeJSJvlCka8GUZ9DWnOJP
FEUR2r9n8BBlCU3fAg2M4yIeUrjj0Ay9GWnpV/36xAmObBE1+h5vQ3amw6M8QXCP8dlHf2pgo6uC
4adWPSR/FynSKuFFSHoDU3I/APbv/poDIMOkfDh5VHlum2dNH6oD/dYcKax9PIVSTrarLwwg0NPT
PTV2MRniVguZxrmgG2Yrn06+6zSw6pxcyKf/f6PsJOTPIzViLnDbnadEowLmCWgbHRWHzF6NblOg
nRqFUb7Dv8W/1RehSUJquKlKbfnhRegPQeAfnabScO5O13T3AaLqnJHLR1UNVMFQiZD9/o/IFIdt
7QSyX3LmyDnYr3Jm6qkXMjgnBn9BEUY/KmtoUO80iWPPoBsQEyte9v5xkekk/aFps/ENKsCj3P+M
KJQwia418acDHHL5LqC6L8VV/5n7QvSEi6hX/afDr18aL4WVJ7FBLVIpO/q6eY5K6/pAI/cBlnb8
3XKBWITvBhWZipxQ9SkGjdswk5jE5H0oElcS/hkhoXKabwU0EkRhyli+XvHrEXZmU3CpBECQUuYs
F6wiORbhXty0HNMBWaMKTEHUz41U9ycoDGNx81MN1TeY8akWR8VhHIY9m1aD4tHwlNQfSYWcpG1e
1JJsrHcMc3VTLwBfWXQTez/4Tv0Bz23eUxZyi6SBZflLt3FBIqPt0PPuuFhFnlzNI+U5so/wUjbE
xhI8HZx6kNK7xmIJ6IONFFbMFpnSEe4nM2rzk2stOGnaLMm8mATO/yyvpAh+scj737BzWjOu9Dr6
0YRWKbwaAISstMNsd5o8iE+ZQJFVeEJaxeFLnVfAx5UjIR+xhB4n3kvl7NfgTSDAgMrGPoPpynDU
uhuU8VNycjKxN1t925zAGr01CACCEb3bYmGpw2eRjPWwsdb5wU8CQudh1Rm13R9V88g1xkI4eHTA
BRbbTjjwLBRP6GquHpsUbR7W43Y6aZIbkzNSP/Pf9Ui3tP2kYSr88GjAMQ3Y5yjswLEzZRh+ah8l
89hj7E7R6HCsMNfV4vvMIi7RTXSdQRPOP3URSqNR7iMBvACAXeSUsN/Hd4VkqdaOIIj4OZm6LvbN
z3eUhCmv1Z60cJna4uW3Btzo+/kzJFG0PMOD4XUTypTYtDSrICnaNffZvwIkKB/IEk+hr5xJozys
nPOMTwMWAz13oxG2kwGwS73qePX31YpWtzmuV2n2GWmYZQf2BrF8T4M8cHHMZSlEoa7kYa1D3Lls
SZ3QK+oa4+wtMPX/wVBqmeqNZ4PufOEW6haeZrmHgLXRA2X8sAT/iErZrQbs5KQ8GOGiDiZaGqVx
e97PaslsUsgOjlA16sK29P9D2lfL6o88I6QUCR3pSqJUqsmeU778c6RPGFHKC1uslNF9wk03Nyw9
fCNptwJ3Q10j+7n+5LGeQ+vJ9vgKH4XaKoshQhW5AeXa2RY7LXJS4AKKWcetUmyKx98iGoQzAZYp
0zTMSwvk/dEQpT08voqLsZs/tZnBsgYJBL3IJDxQO3R9P/7aSw28FCpKwgz4otfhC35lXSxPsLO1
z5eIWZ2n3S7cXwoQy24dF/DbpUPthEDfPbWnh24/Z7LcDB8UmS9m4+tSP3bpHqiFeM3ccVPUoRNK
X3qgTr2XSQ44JI2lR5aGY9fbT4svhECnGh1fc2wlmIpYxAN/j19HZ6G7gXiry8mKvT/06dgq+t90
7RFkgrTCAJYt3Z8yGhvX94DX6vCsv2/Xqfw9pKTfhSWehnB1Ac+sbA795eoYVqozy4+Zh2XjZdCP
yDaV8ic6dTCFZ/oDTw2+/9NlOEtsnfADmqM4WCnny5vZmLr9xrt8ujxX2yecIGY0SbRXktHyaJdn
bqSdyiNf1rWQCYC9aBZcez/9TdLf4IA28fC+x/YJQGCiFGfkCm0xj8fQrarwfEVdJUr6PgmzhpJh
Dg3dLl6GjBqoGgVNmsU1oowXgLiV6KoM1XhBNZ7ypg0yAUQjLd3Nwm+Dqe8AvlJBo600AzalVA8g
m62oozANBq7HIYlfFrn41xgFgSv0fGTm2DyfBNFJaPiRu+dB/uAC6NQpogaYop1Y8jUNdZw6PIS3
TG6cw/UNw0sHCakq35UOqsF2+AzM9kxcgUo+FWatjb9QgJR7RLH4Z0To26yWCxXva463ZmUBomHW
ifed5T7rixprbB6X8nXGBiIERDP+Vms1Zwd7aN0+7hTWCtQ5U+z6382nhZQ96/34XuvLuIEFIOUq
/j8Q6NWPmaNSH5O56c2VsaqseRT6PACTMwRtM9m1LM0KJWnp7AVZezYOg9ZbujaBTOILyaXDkaUW
6NBUHzMpUUQa1d2YsusoxIaQq3DgwiMlTMBn0v/TddkcmW0N1pkT4RYylS3drIQ9F77z42IKFDkh
/+kJ9VRjLB9wDL/5Du/Zy23Oieysx8vUqOwNktZSeaKr+bxFByTbxJa7jZsvzKz2LgAQU4GWQEai
xBfqJ73qsvEQxKHNLzlBvD5Y18h4auscvLe+Iaj2OY+NfSdPSW01m5E3Eg4/sbuZCSNKZR3TOmdx
a7W8MjZeThe9g96MrUY2aVW8xXHnCgK+1vxK6exzF6G7M0SEXmHLYeVrTt8etfG2rYqm0QqCaBO5
wT6KjZUSDbAWLi+S2AWy53kir2VYOdTuTQyF6+juae1E4k0K9fudaGmoBiBUuTX2+I3QsINjTUiE
XoNl2hIRenPPx7BdNsg87FzWGcIibFfjrxdgkqT044zTxfi5EcPBI//pXk0kg5TaWK8dhOEY1hr5
8DuHyBx4GCi8PVRTIT9LuRInGWigHZN9janMmd17op9VdYkJrQlMgRhpNKjWsueYE5QAsA81FQgb
0qIZ7Tlahj1GK99TJQMKTasJ1BxlPK4xsNH0EB+hncPhVo2EVmTDvSgPdedMSqDvGD+NWeqqHFTn
3srQxvUZ2H/EnCRmPx6rfersLPaGALVTa7QPoxokTgjGxg9RYaNcRmdYs97fRX0usY7tqLMGwBxr
mQhUtHg6zvlVRXdRQpyupoGpzQp2zGBFlFvPqXQ/xSjFcGro6YHz9tiVJw5Z2xcPuwDPq86bVoBc
uo7ZEqNxk0HR4BPspVNql/lVlARHlxz840rziC6PY5NvNJWjEem53hs3S9UW1Tt3uxEuTy+U3XFT
1MlYMm0rg+Nm5A8m93sovFkAB3CC73OFxJSENpIcXwSA9VEWv/rMug6j/V9SkdjauT2w2ioc0bnB
bM79Vwdof3AxNzpOYIqqjM9f5GTocM/XFN+Uf5DN6202b8mzNfnCVKxUwjFWwZIyeqbXvuMTq+E+
YqSp+Gsg7UgHBOoTSPfNHL5SHtTPmuaNBZ81ws6eDUrQAinlnIBIbuudYrJa30LcijcucoK8RFw8
xyOxtTqxOzqnWeXqRgHy2NmWDH8FVNYHaECkXaMcgQlrUULZ8p0KytNnocfttW2OFScD1HjToQsn
5uACv+74TeAnHPY2bGeAs4WwHoNdazIyXR5xKkzbh6VCNDu1qyWO9jGjJzCZxriuRcv2vqVeU+CD
chWV5ytIvwuA3QOZAOpMAbrzPcZW/RpZxJTzAsFb6MoGe6HC+GgPS0xjTGHy9F3ZkrYFkzetyFyU
/16kn9X3oF2kNzUXmxWcZPUT5UM3Hle38s/1fn/lusrf6MZ9mykRM/KioxBDmwMwpEQ7jp/JAQQw
69iegl6atwujgEBI0nNGc17C6jHucYM12JGGSbqLffMNxlf9/a85ZtR4CEXIJ2jp/6tRf7g8ojzr
GIo830QHsdPM8xNlze/YaeW28LP+hzTABDI7NRqehwLuWO3aL3MrXJWVItg1MdaMCbzLlDfRe4yh
sqTC79BkH/IdkEKu4BIQ/mIv4mtzX90HKnF+E/oQIqlIt3+oVclA+5Sy4nImjPQObJOxj/y/pRcC
OrVKNIl5qP4VVe3yOtr7AOSpL5NXLuIVp1RKoRVYNosAh5bNJz0abMroYp2j0cfj7pB9LGRvbQ9e
oO/XicPpd/2GumrfeLdAByP27Q8HbUv6Rs6TfmBZgyE2T4R2c2yxWhbCn8z2AqGfxLcTayshbHMZ
oXW/FPBB9fZJrbQhl896CL5z2VaR2jGG5roa5Tq1vNX0D3uNbcRntfgHT5bGA7SuV0sKGvS6shnW
rep/p+xf9hb5ElxNo1tqU5/nJvoJ8CLtJDt8B8r4iSoSiE4Ev2Mr0PN29N8LGIlBfvS2lvFLwi+y
oEhAQd6zi0PPhsafgKxY4oO/y8hGK3+KOB7BArKtgDTC6F7T2NUmomGA3D63/EkiSw/88nIxEZsK
oDuwtzpi7+LBHaXVxx1x1m85SHI4bkdAfMdwmIbZXRw9kLdtsJ3FX4CKw+IYpZnGCCqpP8v9rzRF
cYM/7/F9fGZCstcFYiZ9JQCqB7yZS2tJBu2/g336h/tOk11pc8Kg0Wf1dFk5zGC+o035uMAHS8O4
vZ5LET01sf37U8YUTIcR/5JLQLH5glE+mT+EtxodDxhbGsySYhqdckhfnWykV3PJ9ljKTU+GC/0Z
7yH+tqYwLXu9nEn0ju6Z27sITAtxM9lxP0NkloMgkYRhIy2l+BxvnlzFBXMXw6VUyM8fh7Tiseoi
TWvc+Xt4XKShm/GmqoSL/nn3KlrHBv2vSCyV6zz23tU+sRXn4DzsaD3Ivydy0itokDWQaf7ZadQG
9b98a6fy2J3qIfSlNS+9Ndx4dnU9MH3CXa3BuJT8EZxQcWOuzRanXzIVxb4Aw5YZNOIEun/UKikr
CxFHzU0xTX7IWtenfHHFasG9605QcNTydw4CodBqkHfmCYahU0XkBY2nA3mvDzq6THzvVa1SXXL/
p1zuSqqzZv0CIFflcbbLn5fcJytGRQjoyre9EWBSNxsrrWb16p+T82ReU94HZCC/fQ5eloMvFChm
7i8HZv/P6Jv8J8IWFqUzX5nA4FnNtdaomiahV23AgQ5ePwAcrG6SnDRh4uPj9NL8mgycZUfuJHI2
P9MoCHGMkksM/ZdXb54VZF4XuOsQyaxwbKzUe0nJPAhC0VsyULhf6r6TUkagA4S9HmoK8NRI7qVT
YqX9tQ+ex2z7pNvbeDm0bMpOB8Pfpa+j4EmBDjLdiv8jDGJatr/5qKmtQ/0HhjoV/efkq2WaVYik
BQnSSBvAfGfTyDTa2rmE/aao0JRxjdP8la4/ycPzQjcuV0hlWTC8cv8orawvl9pVkxMTdrr0fL4r
lEp8rUiZ8T9egzpbuxye2jHFqkLXB/6N6OJtcQ7SFgrqwf8PZX21WFL2ZctRfG75yviPlnlBrByH
9HGrrcLDQawwY95uZwTtLqOFetJNQjGIBu2Gk9j13ymqYFmxUpwubH654ei5f9qnk7LSolN1xlLt
FwDYRHMGCgcd4LvL6IZ1vrNGZvMrpf2zjUGGeHj7Qs4Mx2yBLPminiHt3uXdfl66c4ofgETcicqS
4DOSf7sA2bRQ+BsUIxi9qeD827QACnK6W4z40XE98f0wayIGcErSz1CBhuItEnHEyCKboFydQEgy
BfCCxCjiQX84eql4Zr27ZMG9NIYaDXkA77bAgEUut/gTwz0enJtyJJfi1TUYMRP+9F1xwn0h7k2C
qZR7/6PAI5eYQfrsvG8BR0QYm1nsHI6HdSS2tt0MvTN3yMMJWhoAAF/odWT0Wi3WVpRl7P8Fz0o5
IFoku5xykZ59wo3ZjSAPsqZ/WggXxxRik4Zt4kucwqVcLzQyWBF6YCpUKW/BWKd/nRxMtNwaw1/q
t/3HGpGdLSfY6IpWZgEGPlzaI6srXydSl1OttOk56u/qvUOwE/VW6wIHxRIZ7z/LOHULbSGqrE0c
/raq0HYwjOJqC5CG+mpTUS9bdO6iFtV3inhW1jaiKK1gn3c3ANaF/a3Bb63gxtAI/bj7TURnnZtl
Zw7Qu0ybsBe033dav7Fr1SVxkK/A/EQ7vXie39BXGXJMYk7RT0HUp2upsYL8IFlpPRnt4pzpWOm4
xaMKmBuY6Kiqj0SRYNhLprcpJy4V9F0t+c/DGM7e4ipweHztrA6Uxw9jF0GGQImMvb5ejz8LE6pl
5ZtlFZ02bylTgUcm9VCouACwHoaoZINh3ACp2M0f14+2hQnqYGQ+sQ/DJoTBJRchJkh4dQPNcDM5
+xQ9Xns4xNVAuIiVnLw9eAEzsBPqneY874W5i6WQlZdtkE95zPAwnpzTnrc3hCK+FZKto86cxFJ1
FMKwhTHB9lc54xSLEPLGfuBkHhmHAOQcA0oCwQcuUo4eitipM+N/ISdbkvx/kkvRFQfSJO3Xkxmk
d5jtZ5lgmsT2kG7SJnTTHzONt+Ms2jVAdYC3vp1fuivyOb/niwIBdBTSTOKyP2IYYD6Ps2lP6Q3p
DT50KD7yFkKvZSc+uHD7jLIzQDYULfeoJYZCXdIAVgycyg5qgZfW9kwvspKT3NqPnVyVoyHwfXOF
QhSPASl0BkQpsml8EmLGJ7NxXevfR6FABn+SFtA3K+iI1lNVvhh1hjBBlHINqOqNdgxxdeYIFAOu
BrwSjDXE86IftaSlKng1W23kSW5mtHc4ZZoEfxvNZ8rRTzGooKzVI77mAAqXEQ7tY+WzmxXnB4J4
Z/8o806m55fTZ87pprau9jYQRQ0TFqTi2Ql4ZLoljI1pBOKLPr44EzyzgJ4e7Tu0ff2hjqzZFsmm
JPSlEhlNtJnpa2qPBM2sQNAPf9bBV0jrrsXgi3XU4u/tqhKoOfX+8PZbtSKq8CMoBQYjy+0KrHKv
IIk+heuSc8TCN5cTDAio3FeypO5WOmuX6NTgrZZEr++yESB/HzPVYw08p7vJTjdnhg8Lv/iuU3YS
MuZgeuKkTTGrIOVFpe4ciFjO4DoRZEZVFgiO2DfN+Cev9rW83FmlPa0aMNFINEUriz3SKTouzxZC
DNBeDGopQwaDOFivwOANW+9SloJr1rp+bZCy6H7F7xiJvcat3W/tSATiaew6lH+FDMwIW7Xo/ous
81qt8rHI0P0Ouxr4PjY0GsUTXtUl+XVAAJE4mmLbY9BPHtgNE9kqVSs2r9VxzpTpP4XJ3yDowN9a
kJCciqEBi8lvPaC+H577y2N59SRWU7STjY9RdMCuHYmy/X6ma3WHpEcHR7Dk6/OSWIhnfSSSZw9N
Hdrcp6orzqBxrP+ZyXMRE2uaAY22YZ3I6DpN61NitTDc4WmZVIR7j8+JwYwbuMr/ghcml1WmIdwC
I2ocXcnLsKcUSSGMOhy0J1Q5L8ucVzCuNDRKmVA6L2kNykrVc4i1gSsmrTco9MWEu7sMU+57lveK
dRefl3e2lkTjsYAVd1dnRDg2j5jya7aY+sJyPEsENmf2DWGGTW9poYJ0HH+5Vh3dUBPNqWsHoVxC
CxxSBIWze8pJHlM980O4IaV7AhNjKMj9tvDadblQYh3zhdeR2Xu54EYareyaCHdbKJnNfVA7mTMh
NDsNw2tSmCsspCR9Fv8avn5ENcWBZ+zQ9NwaVDtFGhFIRZ9ck4FsOx7toVdAnC14qO8jBZ/4IV6Y
51EUuxfUs5WnxQ2TRnwL3nzquJLl9BUym5dvz07NXIENiHSyt2jLueJDToxJmcAhboaq9gdaiMAO
/ceo37l2HLzpjTR0+vntzeBKGgc68Xt3jIkigoxnqhZd5Mq37O5yDUDsAs37iHnZz7tir9HSMDnV
kYwsVcku8s/b6VsiqLl0KyJ+F82zdRgRBKqzl8mIg1s9dl6gO3kuYBAi+4OB6ZCwrHt7MzBdTjTI
JpXlMWIslRG3Z8ySevJBPKhVRGkz1xYSTODrGA1Lcg99EIRRGsr2qP/zJhpPKe5zouS472Ong7ye
mNahQBCmlwWDRvyM8HLbfh+T+U0hgcjGWmWmciL20ULRqtCIsXkcVqjtrHfPdunF2+lmjubQmbZk
vBpzHpBKtCqAYO5Xsxbo9YdNk2Dq9FpIZlGBXwmyalMdbyhBjT79UfmB1WtGgKwx2wBbeV1u+uqE
r+X7pYo/yE1PxBJMq3kTyOiRB4ZbCfr75HZ4YHoaxUQuOrO01e3kPFUxLiiwOhMQfWglrG42aIE3
Yed/+c1efj34mIjuflstPYIzkUYHt+FcKZ5X6jvX2QwckD6gD0ciX922M7rC5DNHzt0RM5hphqn4
MInR+ch5oNRjq991ccFRzQqmDvrAX30PaB0uxau/f7D0jRTYdkxfC7w1MUpjfLNuFsC95tsp9YM7
dvc/M9+k5Vh11Ktqqr1RTxqBeMU5chiP366CBdoON+bgtZy/Aw0Px9/w7X6H7/dig2s5W3c732az
ZFWjmdg1ht7obdXjf56hTLkKnbQ+4RCkM90zWYenZNrLTTZNO7VYumuTSJAb1A5aMOzWG3iSWnTG
4jI1w/7hDwo7y4lN6RPKybl1QTBW03AOMr4QCoItT7f+bMoFk2mlQyBy+NVDteyhJuPaqRdAJtHV
ttNUxpZnERh9f/rUPHC4jDMn19t2oLdW1014SFoJHU77+XnwRvGdWikAdfIrEeZQ4dZaTWfRjZ5/
I6SRXpHq/aqJcZmSu5ASU9f7OeVjMruS3RDTdZGmvbEdJaTweCCplSA+KgMeDQS5t5xp0Lk/wr1Z
aSD8d07iVoPrKHrgasbl99pXU6bhN8YVI0Vj8I5pXhQaGkTMhsVNOOjFYxCtkIMFRcn3569RDvVz
Uk3k9paaaah8nfPyK4Yhlh1l5Am9xJDwoDSFIr27sYdipeM9EO582IWtDW76Ush879LYtf1Ijjsw
LG+ZXht8fxBLs/vG6bMSOd1ItQMbxnbwoTH3/u0dpczFOw5YJgRs7tFtHDbNksA9aJg4vvr6j3Cq
82P/W4cKcolFxE8EwgjWYZA8HRCeJwMZmuxDEtp7kxCUOr0kMitKG5vCbEq4wrVEAh25LolU1q3V
9bTbPBk+RzDdewNmyzmOQCjr6KGYTCzYBWzAZEUA2RvsfTyCAqDrSucGivVANgg7D82mubtbe7qF
CbHiY6WxcbLz/j7qHHK6Q/aCXPzBQERlCMBqVl2g06ViOyawBS++LbMVefUBQ3DIal4BK3/mA12O
RC0rCVJTuHNoQRtzSLGeYaMdvP5fZQl4nYXZJ6DwZvr1sHVTEm8M9dFYyPwOsSIr//E1q+ClJ2vL
DUNMuHYWGBa+HhIXEaX3boIU+4+8vzvpMKM7wh9jrO+vad6GRpgyNLcgdBmstk633hZqQJWDBXen
WExNwVxGpapbxO/kdhWBhRFGsgu37S+kAwca/zmCYylnMwnaAwsLjh4ujgseQ5c+i64JaVxeD+1U
sLyFbi/HTos9dPZLHd+SEHQwcXE88E0IQoxlluJSXWXntd7EU8EQ0qYpGo6oK3+SUHquYOElf7Jx
V+gVOPalxg4nMILXZ7kDZdH6dxuWBqAOnxoG5maM+unUnskrAkaVLqPZqyLZMxwN0qpqDFgzuT93
iiWnGMKmJxDVPKr2EiqcUM+PmPbcunHX3/Wvj1sCQYwv5J3CgN6x2EWkm4ludUuEYShRoG37BXHO
ySD4QQjDk5PzpdwUPQEwBPiQK6UXUs3G1LTckPjP1lYuzgaNgZJpXjzSP4pQh+dsXABu7tERdNr8
fBFuFhbo/LspEA9J+D6nvVoi7rSVdBSDIkt1CtPWJ1FdD+HZpzx5QfUInhz/N0gy18DK5usQMHyY
lO7xb0ELFqscOC57cKFbrs/DNl1K1V51PtFKZRSmSjVsN2DaPq5Tm14eW0Op4WbwOQuInZZYLbhM
hWv/n+isSZRU4t71QViAyI0m5iftrqE7hEeaut9trRa7WTuuvriyhvyeV6KQYaFjONMPxUG9MpS8
LTazChV6rpF1PFa0eAugQPUUWaaQUK9TYVK749wnIpMTMGJ3BZGIdyJaGt/6MmXSl+BmlluEVU2L
QMGfqK4fac5QVrG1bF7DKm8eHi8qfsPNfvFKrylAxBX8ClyetQjj3kHMpN3FUMWzd6SYlrYGKJVr
d8AcWqYasG+Fxjk1oN7pk0ZYpI58y0MuMSTpyCKvBzhXVnNduYnkDpXhJsjtFonfJkFw9peE/2Si
2pe8FVlIYESVWBSE+Toj7EI1zotdrfG2LV+ianRGW/2Kx5YyPlbVuJ6xikbCHKKUt7FxKMsOlRV8
d35SRXaclaUY/iMuW2PoYSVrmuIi71VdK+OqD1Lg6JLHuNPuKTfGgV5QBHx0XXcI5grXJTf72QTS
vDEgJNcFdm7hX+FCJS0/tK+U2HD5XN0Bbeu56yodvK/U+CByDwDxNKiNUbyZRkFFol8X83e/m0iF
ei2IyhJSm1dz9qanAZTLvSHCGc7KdE354BrLnKua3tmsxx1Zdp1BXGPtka12KR6iVye8VsiqqOpp
2t5+9lWbwq3fZE0pnQeG6DIXvKZEHQp8211iY0YYsJVIg0h7zko8g+VzPPbWfTDRJhTALwnt5bMK
Qi6njopzjSlW4rvTyYjNZ5+ChSgdLVx4vN6tZ11PSytQZ2a9/ddfNJaG+kTQAkRWRaryj4CbHxTr
nVU7CmraVmCQ2g38xUREe5gckVmRloVBa6zt7Dsixa0oq+j/kUwE0dEhl65Bf7N0TDssp7REbngY
S43+6vyPOeF4HDwRaCZZKxC3DXIer6dK59R9+3ctuxm+WC7fqQhTeKPEAZmiWgp0tcsV4sZKBfah
zhmHs14n6Qe5WAd0NK6/st44JMkHuRfjf8rp9/iSvFaWXIYCQdqnbqpFnmuuUerFoLK4Mk+Iz4WN
Y/2MLkgJb4TwyT/wczu+5kxw3ciiznbUhOoiBpL8UaKWP1TSHSGGhQ1PySCyydM/lwkzDuJmmIyc
lDOTMiXPfMTJSG3Xgl9qpIZyPJ3EN1uiT6E8jONTo3BvemEfC1vsg6xnzXuRxDBKgmWSOTxF9v5U
B0/eOmQKvf4puvUshfEBNk8YRk3pFHPi3DyV7/qf5MBRWcPR6XK9OFZFdrZFCJ2ZyGTEXRLtvbE+
xw3aCtHykNP/Hy8sOEhfrDOz35xKwRIfLOxcrvukNYxOloOjHDU/pG875qaQRwso4mHxQMcSdqb2
+Eo7hhhd+lTYjnsHriDobvJw3VS/PNgq6MxzWSy52MEZA/mH3Z8BODF8FsoUwgWrwW/hK6LnKCpa
j2GxqzbP14muy9XAY9Rx03QR+wfPufgjzNHDPavxFx0tX6d66SonN3xOzmviwSjt2kuRt70WXwYD
t1laIRdiW7yarLFcuXMLTbGiFCBOelimAWlCXUcdam/scknZyZOAViy7pJpVUMdrvxnkKs4H/ile
oVuJxvDVntYR60Ahv9pwJlWTkcUvMSgtQjDV4eEeSY6NChRmKda1MxiM3dKUt3HioPXva/0W/I7b
QEleyiEATkz0CLISxWKHnD3DuCPaNip7TeMHPpOoxo+MLMVIa6Iqdk9f9WWXHolQxsyGVYJ4tFt2
dduKdZFhw6L1pcr+oFl62KfrtxaL/+ZU+c7qfBSV9sfW+1dGIGYqsqJJKYww6SHQN7ikiOXa+/G9
jovJiUvJCXqJ2jLCfX/DwaoCg0N/+m2wEA/wTvRTeY6pW8pVvmKLqWMwWpdW1b3T/TReaN47lAJx
Ns0D6+aS/zD5W8/JsYK1r8IWLYC29pJf40Pu/ets1CFu2DUcHRhOJluEUT+UyXLqyhdRHQUF4jlW
QuBb8cnXHRAedkF+eSTsDqu/xUmSbKN+qhbFt+fsFtN78Cz9EDj588IGti4b2MO8fEslZl4gBbNP
lwGS/W8zC2jadmZ1EJpgz+hoRi+od+cAsbBaXhbSR6ebpSujTR2E3eE7Jl+jWL50S9e1/B+r4XHJ
BLDI4jjxa4QAfxtxUrL+ngAWS7ff3dz/IiYqi40fJWpfDMXoeHynWul2CGQLx+cmpfdEuN8CRw8d
8KT+ebkrGEfwXJ9Gb32JJLGRq+wCiV6SDKlrqpG/r4cvGi7ShNRXCQZQXuwHj40jd4C2VVywzZCp
irm7Xc3vPyfWbsfSFP9NhVEcVRTfAAF83viifj+0ctZDGicPZ4BzFZ66a02+SzeYrzZylJU8Gdzp
5Y//1dKDFe4JXE8GAjELOyGTv/zNol4gz1Ip4z8gOZMlz/rWHdv42ue/0hL1RwwPwSfbjyabekS7
tQ/zK7CI9J3QBqOPRMMO7sT+QCCzX1oUZH/fje3GffT5x8RXjv+N1QAtjdMFejOtb9JA8RsaP06d
Qk570inYozPbBu6hmk5EMRDxt2LlXW/jQpTXm+VSyfRjajrNmzgYrQ1LNUWFbGJlPf/O3k6Rx+q9
/ui1+Uq9FI/ofVyn4SUA9iwJ5Vh2yO07GpFkSjJvyn4p3o7npMOe3kpLvmbGIaSmUkTSn5RmUv+7
HeVhYLwcoff4gCLZi+2gJIdOZtK+nNLO6ckQDcvwrmtnSdrwSJSFRD9sHfyUif3EgLJsaTj0I6o9
CvbFemRyxm6TznlSz0cdIWFW1oS4XVhj1rxtW6sSzgfO9i6KP0yQQsyH8zYWD9bk/PMQZwMSuJMO
WHO9RDUlDUTdmF2VFcWH+PEHf/7qB/V7dFBPjyUqRbfBml//AlYiDIaNVoTeFG1MymAOGNDeOS61
kzt6l9/sUPp0SLpN9Lvve4+k0oDuW92hUIx0NvB/lC43H508lzdjQRXGRpvsPHo2xpUb4f16pfOr
0hQvMmQYPA8JGmok4xhb59IYDmihEvj5Hov+nb3SRlSBbKd+EkIaC2e5xmxy+ioXhn5jVJB1t4Aq
nKWj/8nspesxGvR8GEBy0IUAYw81UnHO1SMeaQwMQ3DMdnD9mT7X30PF/zFlXadRHv6y/beDta9W
l2XUUnjExnwVudxC9YYd4Q0+LsbVXBtWH3cCeJwGwrBKPMCYLdaJoywQfQ7ZIG7YOP7KriQkgsGO
CT27wpO6aeDZjf07rd6o1qjraSK1j4ubvaNBmsvO/sBTXbGyB+YX26feOKFBOSAY6q90t+My4neJ
enXiRtvxWblAvc69v7pwVNrM14jWkUjs1IT0A3+C+FNZ+mBG8m3YM/ypd/2oq7WLLmZj+Xg7Pbk6
I74pOn2ZprUmnskQDUuax3rNqR4AuTMmb0nruKNAuDaSW2qfI+TvkOErBoJFTRZ/rN0IsK1Vu4vv
ejnI8AMEz6bGbfVzEsNrDVWs/scMjsq/qvcpLYyLbBzbdQ4r4mEpVRIhsY+Py0TwvlJZ53Mm07te
8i/O2kpBQNr2/a36OTOIF1vHPQX6sL0g+4YWqNOdjEx7agqIGmUwrRXBiy84kK6xMhdV4c5xMXWh
by5i5pR76eqxCU5F5ipmwKhJTEk4YuNFcr7BmX5rvzME4ZthCOtF1HfIwdfeV+Pd3inh5wIs8WCk
RtotKqqqRMRSaFxomnWgboCmSiBJy8xsvQYi/A5eMwpXmIPKffi3XLzQvEFoX5NHkIbyscLMZuH+
/KO77GxUZg8q/3WuNT/IpU/n+uSVaINQiTQzMnqADSvhPrtfHzYKtRYryeDIjVO4uNpzxcr2F3xL
WfOSBsbo9RUkhe6H87HycNPqjB7evonWxJHhadXviMlzZSNUKhN6jJu4E+HnoSbqD9x6H2Qz32ty
Fmzekcb7fjfJMD9EMOg/T7pyhqUKXE1EnPQvvQsvswhBFvT9iWap+a9b2+IhqBP3TWeK9CdB4t6+
dey1t+oylsA/LOZky6QJFvxssEoJLDidepEGkqYxIsfSiVIrCzgiURxhI33FSubllLO0MLC+q3UT
5nIp/8viLo6irmLTwBloLMRyAg2P4bJzO8QsOVifxYRglq1cjyb3Ccim9tFyvQ4s6lZU6odOwlTJ
g+j37a42E6+jawHaSfbxeM+bIKrSLwsKV8NuCBirc3bG4lEC6X3c4CPeYAGYT35PR8TLu7pbzGb/
++MIE/Bqiqaf9WYD41jpgQklM/sNg1A4AvSK8lwKA9gohpyir4BvDn+W2nrmVz68BqBJldvWj+vr
3zHjYSk1Z8CC0fYDUsQ97b+6IOZR7PzeU9oNe0CdIv/e8pwSpy0FbRCVjyP0Kkx6JotZnXgr2kyk
NysVuYdCeuTThPXxLAHCX1BMaVG2Gq+vQvPxuSdKJfCsH84dcAhNhdzYf74SV7DwH9Py2fo7pOnW
oXnOXyavqFP/nWrdu3rLB9FGlcC0OidL8m16HZ7oZPWXMBZRS9/Dx07ImbCSeA7dP8TX+SR/wife
eDVAuhGjn8E6YVb6iLoE06A83HXgmcLaqUyX8qZ2n8Y5zPRpVtUEz6nCmHUBIv3wyGbV7CrZs/Xn
m541CnXZFuCcgp60szjvYKr+AeF3fqMnn0VeIVAlbDYg5BHnHccqRTAYkO/ahunGlNtCjXCFiOpU
uAe1X9HO9AYDg7X4ErYnMApIe/OqW8OAMLS2PDE0am/I9YO/qz0suarQcy0eD1RMmBl3tYTsoRUO
SCEXIY9BY0RJxpagqmtE17LxLg3zIOB6hzZRvrqX6MTiOD7xeUdEB/sTYh4h/+lJAHqexX79CAuC
ehJsWdVozcPzVmTmWIOzOcpbde3ChSDaK1X1rdZ+Dq5I58vm+lXnIaFIJIyNtg2kTid2raTdx7CC
t2pYuwjsOxbMGGnWAWXmng9sNXQUsl3j00Ox1HNPiD3Go4PHyGvaYj/0lD4M3CAf7v8cUV1s1U9U
BmKCeHo2/eVqeQ2fA7GiQFvzOx0bXsTysyLuEQ4wFnjH2KVnz7N+ObG8hCpGpkyphWlw7mB3JGDq
i7kcoyoe7Xq0fyAyn6RnLHmNPdGLF3MDvImjDAhioq2db70iEuj4ztuQvWaJPJaarsH6ytvp3lnf
uBm6QzVJba+jukIYaGzEEtlNexM12oNDwa0fUV+OuQQQRZoOifkk/Q2VXKCb2Yox9yjpifjEHpyf
fem0KBkSBX++ulw9P4rpJGE5F0m2J4QqALIZIi7tNBxEYIcXeHdj6m28ElVCgaH1MzgSF/78hxLQ
tNlg1KMn+C1IRb0v5n3Dp5QKZV1j8+IKh01KKxBSO0NkvC9xfqcNfZmj8eYbpEzTV8L1Z70MFiVH
lSXplM7NdKevijNJxdj71TsQUzcXukRfDc9MYUoxiSeeFs/f95gROZ8Z1akWbcwrBASIfY8rSYab
bexCPdiq/kLD4/O42En41UWxjToeabXs1nUImVZWyc9RKI8moeC6vCM29n/fcbHSqUhPKhZlUMh5
2zb8Px3SZHfqXJxfGNLY1BT4w8xxKxSGqW5rdkr1c/A0+pBzsgiQRqEsujrUH5AIf/OdUZ+OufOU
fmO8uOr4hwLdr8BMggI2/1iXc7eNy6LARnxKGT5rjftHj+W1LuSZ916dn2ZwdBX6YRpQQ3tuHIgI
oRdkqJc4k0H2OJgQVAZzekLbmdUrAht9Ae6UfI46gq4ucLBenDITn/ER/kmR56uLAu580kSl/NYJ
pP2X23L7/GMpy3abLnBhGjIZCIJghUNOvyZpM/etCFEsjGKGOUoKQcPlG5ecIha+hkVAn4fOWu5G
oZAAcoKULj4b00M19HNfX4Z8S2lLQ+JmEYbLJ6IUhy44VXrI7dfd6PJ6MzPl/vEWyj9ftlOD0zYI
tm96wW9w/5qrwfnhRxrfRgS4u5XSPpgvIcuZz3X6mbyrlS3WUqJgGjRU10EAG2LUOqhDR/N3LIto
bjbV5cdGcLK4gFBZTAX7qivsSieLcZMr+eZmMuKHB6SxWPGZfdjejSYfDtb7bpfa+hTFeeBlaggk
dm6YMI/5Snt4gNrxsW/mBpsoxJtE0ytyaYXfHCMYbYXDvsqcXseD5isTAT+lkNnkl/hFLqPIy0jO
UCdxQwUTc8wfs2LXNxN/Rg5oWetUdVW9COqqb4Pr46YMJZtdvimMi6SsmsHSblLdTHxX1cDcVUBO
btpRddRpdzA67eVwfwUJDW+3QNvh/Oqdg24h5V/cTUVTsEb45WbOkALvbHaAOk3E6eFaKgfECSRn
Y/T9/xB0Tm4vEYKJA+BSbi/G+71cDz8fpkhj48FEXOOIprYq2V0js1mYjhbw+6BhTdn9qJDBh7em
abygLniCOt2Bx/IURqxcTsTJol9LxZzR6TFPCbJ3jmxf7Kvoi9WmLEFzi+n5PgRY56c7rsStqvl+
ywZWfo9jas8+tohXh3vuXvxcmv4ckD4Kmkx3JyDLIK0IAPMbmi18+wY+h1pfC7EXInP6SmhPdk00
6wR4/mMegKuoD9SImuBaj1U+7ji13lzpSJwxzF1vTC1RiUTWClOVl2r6fUg9kTB2r6kPMvKNnbnC
Xgwns5KXERhMdZGEL/vc95x9RWslcoTTMHe1FU3nS/ma1MLJyC3ye3DblxYJ9Nyb5bcQKIhc3xau
IirfliJcuMSJrIGNlT+UDMG/eowKS695lNiqHbss1xyTyc5ddhXgYeEhLfbPn0WUnfBLYF/5F52Z
OHIz7uRYJ6KKkcsYk5PZrjooy4EXnS4Srysuy58dITSTf6v9kvSQxeywNTDwrGryeCZRmpbZ0bQ+
lfm0ZZTk4P/AO1jliYRr7/7gQWpWrxCXGa+X1KvC8J6acMYFD5Ve4WuaPgFcdha+QUoXBu0qC/OQ
iknTs/rkSTxMZ9i5e4Bmefj9dqEqk4tX1yF4wWVRB9lDfaDm+mDSM4NYmbDWJpqfmdNs5p0Fnd10
jST2cHXanmyyT3+k0P1RWHMjpY80D+xdHY0OKo/OUuNlRZr4SJKeEUqEf1Jy7/6EmTMDR284X58B
84iFX/zJs5V8MF1o6b1DUIHhrMgH5juTB8skwZ7bmGUg6AXIFH4ur1wSQYWPT49bz7hemPxBaANE
kvMfqkmUq+cWwMKkm/b2td7A577g3fagxdQ1ilLUHYTd+LFVFGaLZhPbjHvyocC2NtpmVnrhHTBu
vJRkaEP6rUXDA7PhqYp/+G+EB/dHu+TXvjDYV4kA/qfE6SllcnYX0q5rMpDqgad/tQwV7qZKOv79
LTRBcYOPqMDbEsiBfU/ussC1YP0i87ad8GHnb2UJgIFfzoPmh6XXHU0lM/PpxRX9ClG4gGQy/WBe
VVZ/O0i4lpHB5B/1NQ1Y3BXH1QIWWgjko/VmJBEs7aXjoQ7+jftxetW48JKaNzg54V9XWPdEKZ1W
H51WfJGOL+IeXzP+B+diNEca45gBe5llgGmYo6u7fu61LPo4rm0KIH+i/sue12I9unV4/9M8bDS1
iygRAeGkPfV4nwIMh5h2QAmKDbyHVGK7engYZa+0dT3sn5WMFsH3wVzdLE05ibNDGzL9cAsW3Mec
fR1n/k4Xy3xAP/wpW/yWlMAr5NiQCaULlW1fpm5nAdx1Vn3jiYXxivQH6sqsqs+AE7O+gMno4lii
ZqVvpIhmwFvd36mdholCLFQcak4K0p9BcIoTglHK6S9WZnGXBIvvqV5geZ08e+kllC4g+/Em3aD5
mFn0Y1f8jUQbbL17jB03umUuu8x+dMm5kHmJOoDqzey08L5YR9w7/c7aeplFgkEgle2hg/lQiE9d
TtuH0JdQmJlUsJuF9Mw0vZIJnmb3W4BqzAkPdxlq2Q3i0XRQtqQycJKGTosomgb6xVXvyYFgRRTr
xMso6/GKgmHJrg53t8ttpYUZBlZTEpT373T0RaQwQKs18V284n1abACSWjtbIQRmytRO+PsMNThX
haE15oiENInlb827+CDoClneYmC8nIqpI/J0cl9HaO1VSNj2Ekq7Wj8XyN5XjY1TMhhvPdbiIBE2
kczp7mthqY2qeiiDzlmQ64bEoR4HQ20GFAQlBdx5vMg4u6LRqz4e6mMggpcgQiKErQ5C8zScsTq7
Ou4N2E0iA1ZopgQcJR5vmVkmf6noesLLBvWKUaGr4FJSMf2C8Mter8j7c3LztiCxI2v+MbOisSYD
hc7U8C1Be8Xa/8NcZ3J5Z+n1vio0baZmGPiB3wJOSpky8LMGGClz4wXXX2Go8CZruscmE4jqPrcs
BnVrSTaeNUgozDBp7OT9yuDpnO0cIOvhNTMjMqKpnL8pI1C1QI/eI1yDgPN4+YGRs1znNeq3TZxP
tH4tKlrBT6nWbRcwUzWol/uhpuJYx2ya1PeI70Ug1ThJF+Lijy+FWCSbctRNf5H6x3Udx4fWgX1g
kOR8+5Z17YxoCAdDXOoZxUtgnE0kHpMmX8iLfOR1jbzWvY6HrbBcCQ+Szr4+JigXiZ1S21Wsef4h
qMt+lmtwpPjiCuyhMX0Ij8w/GjtKDUxByGxnmN6NG16/78TNkRAEzKBNj4h7PV0M0V2Qu7c3djZV
XzbLHTVxYr+YJdIyy01I6T5+IwjYx5tJFs1epewzF7J3DoZ6+9mxU1+DCpuGcWx6OcjBdvhAZRfu
J0dnnBEqiK6xIRrSqmG6pKKbsfFQ0bPPKlNUyGbWsQbJ3OUxIQF7h8uloqcdzCA/laR0CaDAhcd2
bTa/P6QNx/Z4zx27ZD3TuCWuRo/Zc+W8Uk/pJazmL7saMOOfhe9FLyNLXwa+JhOBSM5Ndlh97iOO
hEEu66vUvrnKeAmo641Ux7LYe2qg1pxjuYQePOSC6KMq1URyuv/Uh2O+tJcr3DGMzKWEE2oLRLKw
4e0zgCmDXHvXBlKegA/iC+SP+rD2oF6wDmxSYaNdDN88FwvhBcl7M+Cuajf6KVfjW6pY5B8Yqhht
yb6M38NSy7MMTGOy29PbHvDWBzJtTVmukI+EBAB2rAguPkVPvLPk+zJSQOUvBSy4fOZ2s+ZjndsU
gluz/0HMWS0n8aLuZGQYGBM6CxY75nQaXXTmqcSCgSALl+wUnc5AJnIRdO/9gN8P19uovz030XZ+
WvbVjUg4xc1/ny/4fPEJ0k+q8/E87yyd0J9S7OgJHiR1r900JxUJQdp48k/et5DV9qaCQq2rWJgl
YEouV3IX3lgj6EWCotP62rYK7SrGOep8Z8UtKlQ8oJXOEcgExNRHv9fJn5n1KqQUBeUISVeUDEQO
CpX7k2hn8IvJcdGQGnLtSuDLH7cRsmd6yTZkJUNR/wZ9ptSQnlpVYuirndJgf/VVooIKDeBGtplS
mayWRMJBEs/5r0cDBdBaqtSDLoVLN8WzOOG4aWthdK4imlXZKxnddjmnqDazVtu12ifJsAsIC6v9
/Y0jfT9Pok7T8zZw4bzh24yLD6byNRIaqHMyIYkqtGPinu5tnrmHpBECqLsN6VdvjKlWEVBsOcaJ
dPfgnM0jY1KaJFpUekmOQfZTZss9PyusuS3xOxWPe22yE3N4cUY5XpKM9DHp8BMP4jZ7lgbKxytZ
d5SQW2SC8d48hcMp96giAb0urXai/j9T1GjVlYDi7i/eD2JLSWZQZ5qLSKuHhcyZ0Foct89ZFFyn
aXTdSCSI6741MZRnCYo9ZJdM+qi/k0s1UzYx4dI3rxDZkA2mQiPousfrrA496oABJ2+ouVenx94u
gwor9JDKOlpWsxVgLWwYv8JAFNpfbpI9LCqxCGxHgljJTeIPKCflwvV1rtP80blS7AHjAYB6PLhA
Udwk0B2afMD3/ACoJk0M+hl1jD+bz9dO1LujEYaTnzmWV35/PO26t8OkkflPoS9O8Uy1a0ylStnb
wxx8vuVoaUP0EAhH40MdLWfT6Rfz+CPuzaEBY7+R+Kl95OxgPkQJ9zXDjVGfcJsK1dNSJfLbudES
emDiVnLWzCeZNkbynAKc/JVPIJ+ko/hlYIOzDqsUK2W1k1k06tH39Qa+6q3YoRx2XoVEexNrgjTi
TLRcPnLsv4e0OuLlBQC9mM43qQZQoAuXE4pIi0W/gkuwN9rXI5J3s/z7andIuR49iwpjR2xigjlZ
AoHEBivz3BrUtmE8j+aF7SJmgmbezov5RZdm/Cu7LJ3k3TNWIEMNJwfzjBk/Rh5LjOqZyVgGUYn2
2kuP4FGXF5I7wAlNmODknVs85AKWuJz/9BFbVo7suAmxNgs/3zzna6IvFHzGudtgdx/5SME0KqPx
ik8AsZ+sEEPAbfMHRyc3yrJkoJAuMTjr+pRXH6m6U+VkgRcBz8Z5o+i7QhkWxKgZPR1eBY/smcSq
RpySZrwTZp6Nw1fjrLoXLvVUF6XG0miak1VQWt+xsvDigb+ZerebtoA9sqo/yit+UesWPHuhtLUr
3b62Rov6qtP2tB+95vH85wsZiD/UgtFcGE/3kL+/5sEx3CAM6I6fCRu0V3CZYcr2hstb9bM5JYnC
Fk6QSsiZj4WaPRSlj5cdIuLlBufaTaQBZ91kbJid6kQV1X1hKqP/8b+FwFt3lEu1jNTQHrB3a9HU
LL0O9SHLMI6XqZDIxyXWgu5CK7sKvYkSuoa2JrH0KVx6et+d+kfp0UFVxBd9y4Tpk798OsmtZFbe
RU9BdDxc/MZSTZP34Y3oqwRWdR/El+yTcSWUeDIwIU57jo091ByG0O6twGeyy+WZTqCBg5kmLqtS
9Tp3pwu+ZYXJv4d6P3iIu4tvlMQSNs0IO0Jcurgkmkg/wrL/Bfwrx6LHMwCHk1agYkC3zUbrm0FF
ReNsFnUC4CUtrJHY3h7MqnCdoT6NXp8lk2IVg9h7lsExXzM/ump7Gk8ITa0aA7ZG4do7h4WM9HSI
R3j8i2UKcdkPVrx6iU39/MK9E8vz5TQmRhRjSPpdTEYFrOQ/cY2TWEKAYnm/8btg0xADln/t/bHV
tuQG8bIW5TFvluezZw8Fk1TPc3Xr+gQKoD7dW5mglftDqbTJXMFNt/+jXMuSGO+/fdBuKW+3TNMY
zAGE7qtGxAWf4xTb6ZHesfxRbULTjDtLlR28Ka363LVRBOVkrXVzuRgf4Xl5bT3Bz2WqgsMMTtH1
B3kYt0aJ5kBM8ky+7idg+TDkOx6a0BxgT9V69O1upsw/ZYImkftsjCl5bswmBloY7s07F2ucEokl
tXJd7oYqxh87VgPQDoSdYSZMIEG5axulkxGqgyePJO55khdbAvVCHD0qBLr526oXIF/HiuUr75rz
ZbMBca8sOoUDPaqN9FWLq4fYdgtpw0v5EKa8PJaf+luzKwdHZonLXl6dEe+1pXSihmtesUgTDNRc
5v08ltZGTb/l42/l1ncatgv4ALOQSGdvthzIhRHplODLAZjPx03j4BnTwegdIW23lywd53C9ZEw/
GcE2ItJ+KTCgQ+OBMp78hC03s1ZLK2Vv/SyzxMszjOCpnPbSuYVFVzeUWnby19+SMOugzpYTe+cI
vdVQdiDox/rJqx4HmEdBc54YzqhyvmykcYMXSePBL94N6sNk8AXsP+f7FVcjJNXHJd4soQQYiTwJ
F4SEjIN1L47AihIqYx12CN0GOtAB53Sqn4BqA2EeVYu3ErEOmPTVtgENXFMUMyrukBUCD2HNinlu
c8c+kgZPakf7Exb33VOWWyRIA+yrAbDIyDwFop2ibiiJChNoDsHBwfrFu5xB7U/Xv1mCfeoDtQSd
IYjZZPgHBxbphnbZgTbQ1jymBKx5tpQShMQUlWEZgTEqA4GSZ19aozwyeacSEnjYQuaSyweh0MRn
iWEOQBT7Pe0FT8r5kHzyTNvXxiZXp7pAACroxK+e82hTI1JirDErwbQXnDoMOP/RA37ixGOVaTmV
zGeC3nNCBJdSclFECHWHtg/BShRUh+iI99vkLfg39QKm0J2XSGFfPxONAfk2s5LkQR3e2IL2G0Mi
7hbkMvln3Ck6WiO+Dkle0XI8irYIYO5TvWV+rhgF1Kxydsj8m6U8go6dfBm9Cv9tDPJn8NW1/0AR
lmfbzTnVYN+wYmSVQW8uEFdz8cV1xHWo8TKVCv7Y21G2J7cgOt9Vo7XWDuPAf4UEgxIdpwrLWRig
zSIrWzkeGcWoB+fvA/W9JMnhQQst1+4Fsw42hkzu4iA8s1Bqka0Tw/EbC7Tz3gqIMe1sd59esex2
dZ3n6eQnmBvQGBJQlwZw972DvDW2sEeQPHaEtNd39FOyeCUohovF/ero6oz3zK8Xp9j81jzOSC2+
LPGXTE+iK8VVvHOwrlhsIVtsFIvnt/K4RqnVKlpfaSfFmAqEN2pZiGilqgXqDLg5RRabTlpz/LH8
IU6GY0p8Huym3kdL8/zNDudVrVWi/Nso3S2CmIIAZKG+Jz5KAbVRL/jQqo6+d+QdIl94vt6aOxSG
o018bcG7KDLGenOmyFR40xsxBZNK0KGOcw7+PfowX0qksDqMZcM0eiI0WzIphr+llhvVnezlo4Ae
RzWAHkQ/zPa5P1L5VevbbbYsiYdPbXyJBUig+zMgFFyOJCqZdyjKn6TBZKSv75658PG37I/RhkMp
5gYGHL6W0pWEl6lhG3zyV46CXacDBT1sRxJaBqXcXymQyrk1FdQcXy9Set0jfGivJiBcBmzWpfB4
RbWEu4pvvgwDwjxBhl3HVHs5wq4T+2o9Yb+wDisBNTFdFkwxR5YuSSQUNoufIJrelTnVZn69LqGt
7P5Rvh9Lo7mGZ0qk7sBOkOcKDDt775J2nYj9eKcN6TnJ3gl5DtudkOau40oUsUGUxqwoA+T1+ug6
xUksmg31FBqkIegF24aFhJ+ENu4iNXfPPaAUOx3VJBrhpjejzSM37EIlt3AGxAiDw149gIlSBqtn
kgdUyvzwsEU7IP4haQ+mSXN+9pyfMloRaNIaChVG/hkLQg9PC6txx0qSgUrbomStexBgYFNNMW0U
FH5AeQMZmMRLQKg5prTAIfXUnIx+u/+vOnWoP8qE/+PM/yRoQmAjmtEv0arB0brCuD9x/+1jYEW/
tovFwV5oxtmSnXcRqWFX+Q+e/I1mYSgWJOqNF9zEoErWqs16uc4Zbi1zYTKEItZjDEK3TPIJ3iCP
aDDaI7xhC3SzZugEkssgNJkG3FDpo7urN6V8GwHxnHiDxybq2dJ090MvN0lQQqnODHrMl+kyE+eo
Xmo36TVzwRmwnrbGFDQoa2hBIgoBDc97MgxV6TkOJJCXnPu5nVpIhzbZuk82AkaGUF+T5uAQMMqq
ZPtaSvdOHuc5jzMICTmbz2b1/vg18aOPHZ+WdrNWo/Lwjorw3DhfyjDBb+6sjeW+bnJ72fCiId4O
pDJIbI1JAxcimr+x0comUwhkfsJk0UwAMZCgponXD4xFBpdGC1BqBQeh8gH+SNgOJVrHBHc+Tn3+
fwPLQPlJBOUtngDgUsKihHfNTkgCqIeWqDzwoZIdnnc5nzfAan/NCZsJRBzYo9GF/NWeMet9d4wK
O1bDdmTR+99miCGvZUbm6vSpmWzlAugmzsA7gSom1cuOCUm/mK9/wAXFebgyVCYaDTBRYONw9JiJ
bePLgcr+XxXMY64KeUSgg52zaaq/0vvRq+GHyfnsIS2PFE3aG40GhBFRtIr4u6rPBS89fUes5M+x
r+BfBY6O7nMxW3Nh9rp4bOgKeGVqSbU015pfom1RlXA+BfHjcl6TTL82wnJfyRZLdovoqeuNE/S5
EmC3o0iJuGx7Yf/hvBCR4pSZwHmqFTTzCUBDYAX8q+lHPpwk0Saov8b1cSuafX1ggB4zMIFqh41e
Y73AuRrJEu7LZp5v1Ywd+qOOrCu6eLLxdlauDWveA4TYs6XUPnliZQ1Gk95JCrICs2Tcmcl9jNO0
0rVP2DDFSyexc43wCConBrH+KDhzFv/v+q6hM7ZmR+xbdnJyIxaiiokMhhfliqWO3bz1sZ1rhq81
S+fqAWwJ8sh7f9UGuSK0OkYnEd1ja4Nr5JVYhpO9IRFYjWONzcdE7guKF0aZNlDeCRkcKWiYkil+
ykZAgfFqBRgTIpmuUwnYBBe834yzvEwEcy5i0kmJTsgAo7OgkGa/9LscKN6+CF70RqfyC7mgVtMX
eKhRpOnmd9DNbx2IHbOxFw8WnPmSvee50GHFmgOjx9cK84EWqsI3EQn2qeq8QPzOupaousTb+eKA
OAZi4yTsRIsYLYvbkmnmnO67679jZ8UdPVa9f1eGQzrgohKORiG3tf/ISLW/4QATzGIDLnF2tmZ/
071GRLXXNd7SfCukyxrA8ZN+h949dv6hAA9eH9pIJRdoQapx+HVLGW2Bxvv77tgHgHBduM/dfH1I
RxI6xDRY/DRxx2DuGJ6FnU4lppW9qHdPOGe3wWwA9zyxReVYDrNXOHqrBP5DQiwbiBMiIRojg6Tq
j4YSPA8DIGTp131oeZs9aQOhL3GYuPtMfgrh9rgdtub3ILcYKZXzkC56FS4ceIvzRjRrAz6ehFjy
Ut5ebdJNQn1vfnN0C2mGVukJK1AhvFj++MjFHYoV5IVsgb0DJdvz/Md4BHL/cgg4JpIIpDfC48iJ
rj3iAdYLjH8nppwtGFeTmk12VhN9TPQKND1zGGWK1mVaZ3LW5OcvYnSoSdP5+dBr5D0rH27WEeVa
H7IvaDE4kxESB8U5v7SqKhPiXNqQkz5ltWFOivJUC3Vgun91p+/MkYG/CYJe9Uh2QYRK+SGApL/8
7TzP4jIQvQA7poqTZpiydH2ufmPzZ7vdPz247cVSUfojrWsa9UVS3I9qyHRnIRfwQDxCeangAd//
D+QoRgMd16MCAyjLepf6vRHklpr+j6SWipMZUqjfSCEfw6pxVa+j8DgI72oGfZbILTu8X+aTSycl
fcVtAJVnsEgR6RIszVVLzlwOs1Y2aXk9qIp5/WGe3ZoOo9Ozr/Cg164IDgXIC8SH76XEq3AXSejF
kq0kUDst4OvRwF88CiE87lNZ81w4oDveJzwZM80AoY6BfU0v6mtH3H/aIxf002Nk9zuIvAjF2mln
5l7OJZl3dlCIQDyQKmCaQSHCdejO3nUAheQzETDvIsSggCGR6LGO/M1uTDT5EyZnBy6cAB93pjXZ
P7gR5tO63saQnIxXJ9u/2rkl+dovWfo6aNrfc2PJCOjHA+BxfJ4Nwp8S+/Vhc1qHmhxVB0KPZLSv
psPn8kM239fGexoy8AHwASUZ8vrmEoGS+S4LVZlwISe2VYp3exLi1SAn6pYJ2THqWWKzjhE/OnyY
IaE2gu85atlGgRQxpwlai9n8YBDyG3OErEzsGt/fywlkryFLnOdgEPY/3jvypPb5iLc6kwrhZiMp
E5ESqrqg3WBI7SrIgIRR8yujACE5dkAvVPip7zG9yYPOUzZg6G40DyfgbI3qmSewTUMBj6PfXIq5
3xwAsLFLM6QLIT0ol80ASQO9wYXEhsiL9at/FwawCgT29JSPS44wG2TZkqdfPmId1/Yu1rj9Undq
J0nruLBsx42xbwdsowZPSkudSQ8aFADQKSUElRZ0Qm9zXUp8g0zhgWJ2CWDS8eVoncszB1J+vxwZ
MEjIH3cDWL6jBhlGOPy5bVRXqlD5dWTFm1Cwck2iUujV9sfW3fDWF5q2QIpvreiX145l0u95hp0x
UdV2HO07ipKVeXf9X+bthOJtlsBB4hHAV6mgTlbBrEUrX4JapygcCqfiJ2ADUikx9aZKXHIbRiHv
SQIjkEzlOHkfoHG6wKOdFc38rnXE9kQG8ajs387lGqT/CEKo8ZGu5a6vy8/9W7IQaECLkyq41WXf
XDmxbT/sZkNs4hC6GCKintu8ayrXcfZoRNhNXlwYVfh9c8fUL8n70DByK6pWFRs4hFebnFUQmXe4
0iLYRJ4B1BASZOnCd2AFDPagyeyXy8oOBST2JgkOsQijxYNeADnQ4OvNYFOGomsv3+KorBVUuwVm
zYiIA7pLpgQGN95Ngc9+idYUNgEQ0LRRfk2ypgqQlEzNPqsQgQi3XZ+eTkXBuBOApRNl6/F4PQqg
AhECeHZXJ7yCsfmjBTI3d5BSFEKGI+/+p6D4eiqehS1fs+iKx3NjkSNw89cTf3+YwgkvU8yOYfLG
8vovU+eEB7XCAloEnWYEdI6RsZHNrwDSb0gUVyw0363HXSEjV7K7sfV/d2ebrOw3P6yH1n/VCyA8
hqpnEmznk/VgjzOfLKtpUOEUprmnw7o+degRsGdEFGPWJ2qDEewCUMVAeIwiJvbMEM22F9QB3OsS
LuyZMvpUQsm9ofPZh+0lCF2KuqBunSt88us9wcFPQD1CjiCYrJj3RSPA/QRYWVrqAM9yVjKJV+Hp
isUnVRPoqY/UA75L2jHztheWY1k3jIdocV0qbOooNN9+3kv/e/A8z/8wJJKyYfgdSl90GDnAkzDK
KrcRL7Pd7NoCQCtQvqlAd2XtveaMsLhxs7pJDlecfkYKY6y8qwA+7M2n3dqezIfTb8K7LNob9xyW
jbrBDUN1Z+q5WnhXOapVb8UCd10oB8ovDSMLs93FHw7aRQvexqWaConOeeJmi3BHXaEisLaZ+rNC
OTXCMLptvY3E87IERApY4dW2WaIRTEtTPPwicRTxH2V3kpCBzO/M6/3zKoca/RQYOk3NF2cErqx2
XpfnGiL1BJK1HEuAGnIoaTJ2cjmI5gpjsb5O8mtZ0y+Re2o1dLWvWHyWIypMejelPTeONHhRz+z0
q8U3HQItbk9fye3lepf44nMzZAQMm43D/FeB5i1VHdQ7t94cDsgITJ6xUfnig+fo4HGtnrw0eeal
n/1rS8mI0t6446j7ZwOgV8bfvctfH3kxKcXzgC0pDFMzAX72ADmHQ24gctM7iPYRNuXWMKZEBFk7
LQsfLODmxy30ETflpQjTtInnxPImU1cPsjpGtd4o2VAy3A3NmbvRNte8kPTZeGMjF90eeg5mAyNr
yyMjEpEkhfVhuGY5pb0HPCL4WTzgqMMob8OhDWXpX9dsvkW5FEn3sYnXypbqeawjd4GBcP3Y9ZZH
79jkhi4U3Q70a3TaYXYS9RXFpOvzbVHdCwg7p/jI71f9FzM+F9PY/fuQFcsx2VRRs47GISG+kiM8
qc3ZiTP7YXOu9mlN/4C00xtsUH17gz8F+hubgZz1L5HtQ5rANr0HOe8rzDlUgieg0LuKd5A0Sw0g
lGr6GGXEJXb0mCPyfcgEdhi4Xfl9uo849QiWHQMiVnNvEDhVCNKn9V3tbMD2g3y3BfWdlomZhWPZ
jh4GtrXTyh/i7oLXrGv15IHh3oK4VxIQRDoUPaMdtVGHIyV1TuQfTYqTBu4EM6ZNkhu8V6Daad8t
RZ+jqnPuPftitxxwD0SlPuTsdD/KxdRsOxax7goF2vnLbNh8+w7STPpQSBL9DZMtSQtMivWsPdAa
kqQ0qOTznWrr7Q63/lNhNppk0RYp/KO6F9kyso7OuarbFeLjoX2u4+ZYoBCQvwNbO+B/0T1DKiHA
E1pj0/8wRlTbu1OrKcbq8v6++0l6rG69UJlK11b1cXxykxYzc1tSbusGJi28aqOLhbAJrLZSIgAf
DvbsOcLcCzg95f7qvZJPVJG2jN3BYdRRCoqs/Hon4ar7iYJJvlrBJupdSM0KRO7bpkckgn4dho8s
+5J+H74xFr6d85bAr43D6d+yHr038WLXKoV47lQnXcGxbGzaNUfjQ3hoZh3jaTnnbgIWUyIqbcvm
9nMN1J4NjPm6sdsIxhbYWRWquMd+M33mSCdITOF/pRvFLngk8TVa0Om3qvra2eOGAeQ03XuEj2Vr
hNWXAw3kh/WvlsrRwQkdk2m3uHGn30GPXPAc9v5rCZrhDShlYvmwbl4S/L92zuAQdL3t7MVem2EO
YF+VdrNt4jhpNAJ+TraGH7VsrH2mHj9XrwQyrMeTuf6Bqt8CCfeMhbyamH2AmCRIxOmPZclpav/i
4m5GNJKF9ZnC2zSOJ7HrY+xLQXtoaJh2W9MmTfNQsTznu6hrUiyP33uKBCBxAjfB36YaHpeAywkl
rb6rE3sFKTn0FJ+gbd1wjN4Tn63f1k/LjLHf2+xbw9W/5qNpy8hl3HI9DAQC9tlDEixW79If6pyM
vtqr6+c8qZPqLo9DfxSqJc7D02fdTR9NPuYuMG8L6gTTar38V7uGgjNe1jBTb77kh+WXT23BA4iq
0FKII8Gd4BTUm7N6mbC7qa1ZK6rDbUEPrT+RNwoOWkXig1iU9OtVD0MEdHJoSBKDT9fOQAit6NNw
48U1vAsLcmkLVhAy68xIT9QJxEg0XC1kmVHu4WQ3ihPresZyNTka4M3obdhBLUEJEN/GxS/PIm3z
VsnJYA1MkZUEdGpodeR0mld8izOT7lqC9FmMCevjlfv3U4ICP7KAhOyfGjMUWAwmouthC1pKUMIH
yzQKLE2WobRsNpIkvO9nerSzK6A2iW4QL5HkvoMhXvifD4/3YYGropEgMmnuL13KghVGq3QGku1S
nyX0iq6joYqxGB2Vaqcdk/jrTXMGMzg+rQ9eKQUCvOwfaN/dUY0iAUPEQctaYcuiMcSshuD1+ntV
ajiZdl5KBf2tJDozVtUQQFWvtGMXsRIJYhgaFI8b4wkzdSahlDbe0c+brwiN6mAJZLtptlQQq5kU
3xrYMrCw0PGLM+aWVnmRwCwcvBuCp05FIqWD091ZzSW2RQT88k+rZ5bwBx18x2DUYEuvbtrpSZtd
bH9mX5gjwsLSqENS/W0QV7djuZ6HEiA7kFph9FQ8D5G4ZqcA6RqYYEzDfywHxC/KY0ikOi8HBtho
76Il75iSxSqiQiC6EGDWuHpQk6CPbfcBxHFpsfvanemJkS8dxCd/XE1BXTtq8Cf2wG9Uz8KfuCxc
tmbcs3LOrs58UUESWrVIzy1N0oROsgMdWlE5WsyDPJJYArmaecpFgysihNDDUs0INCL+PLNPEKvY
3aqV5cZi+X61iyXEx3tTEt2pJ5RmwkMZ7v78ApJclmfSTd0MQC3Je4Y93Xq6cZTdxJvdLQXM/E8s
fpsnqfugTAwOUMLiN7U/nN3fGxrsvPZS2Bo6bpcgYmeOeigoTr/ehqyTb0POaCt1Awk/hW9pL/Oi
XMznkjl6Wv8NN9cT0Q2Fe76dktghMJgkurGf+N38bnrb4Cju+Jr67SZHysIT6z8ht4yL2wQvJ5Xw
2WUuCT27gKEsNysExlkg1ovarz1lYN1WQglzaDaUPFsun1bfsMkFEOtE0t5hRmO9TqPvaC0G8jbP
9lUXYtHnrmpBjYCh64/GWYuFYA5BAhAOf5/lY4t97gMgZTE6cWXiDM0fUYtrDtyKkBfhe30wFR/H
89FdV2q4bFM7hWEktDlgPk3D10HYLs/coQ5dYTwREexlgBMZtwVGgyiIak57TEOyRyTnS5/vwWqn
KvyaILoOL4Sx77Sy7CqUz8/Wcn6Ag/ZXKGhaSdeI7ojJ5LhU0aHz07fBSaP7wWCVlrnC+WrBQRBl
7GjHMMFkD0ayJ44GlsHbBdI8Ic4amlHEnBEVtveunOIybx9mftP9H7/Cb3DGYEHJstu71M8AtUAX
HZV016ak2DC/BmHDMEpO8IviEAq/4JvHrVQ5ssN3qVXkNL9nzi26VYUS7S7COkn4+2YFSJp2L0QC
SdEjAi7asc2A7Q4Jd23QKCYYem0A1S0G1P3evbuisYu/kPF+W2bdjdUm7wZCsoJcbZ64sOB+o5p2
pUgORRUe/zHEeLRZfKTu+H/vJOyu6AUlT05K+iJ+yKTiwEphmEXiXeoOndiyfiBABk467r/+pr9d
DBoXYZxPM7yAF3XUdjRJ3lQXRM6IcLg3PKxqpGVkHu67vQ8neoSq190Tz+ooISnVM48uZnvxNlB8
f1VEITE2b9TjLU9ywCBLoe5hiMdQW9bYTtqCGaTJRmWmL8sslOLkOL5p+RQTBgjfZK/ODSCnfIpL
vyqJYlMDiE/5WsjCa8eOd7OGi564l2XQ9hGDldf5vWN8GYj9vgObzfTNT5cNdns+I1ihi6HDvm5z
idg/1aZdDEysRfSw1HkO7a2Vn9fSNUPRaNjIdaw3tXnqGjN/7eia6YUiG7M3pj74bpSNXKq1Qt0G
TFap1tKFWoYDtGLQceo7t4P4LLERwNoNdehjfNWcEXZcJaZYDV+LWQKQb+oHd0LjLKffIb6l04Gz
LvYOifikQ799vHo2fwYn1GC+dh55oC4Q7ikx8peGU3htHgYJbf2VYarc2cwLlehlVY7r6d+/BXZM
Bnof/GegtolHorQVJRX6BIJAK+eqivj1WDwyv6/GpXs2H659V5JnGLlwUrDN0Vmfdn23oncj9/RZ
i7/cG0xI56ls3Q89q6iNxGijFeCkuE3kYyGz5JQcGf7GyoVhx6/sEJcVvVI9qra0aYZuKdRlVZD6
V1DVRESdSjmhVx+b+6h7XnyN6kf95Vd5MFMm6Uf1SoYfMOm1m9CZHry2C8x9Uu9ZeW5UA53mhRYm
Oi4ll35Sfn6HooBuQSfyg+PNjsDt4vrsRDIurlaLm38pbKG/6CWn60fMohOfmiV6TykbPgu+vHG2
m1DqgR0aq5QFsf8b2dBROdHNdjO/imd8+XH+BY0sIXx5fOLxfg/KrzkhrCON90GqZNF97UyuG8nj
8gfWb4RTt6YKJITdX6ajezf8/tESDOIK4GrLeWkK4ROyHhNiE9hReGbP6JZFKlxPYwQA40B+Xk5f
y0CGi+CfbPUyXoOjziBDbckYDXDkhU4embNIt3YCQwdnbojcmnvTjfl+/Rwu01AYVRt4GcUvzxeG
0cp4zzzYL2d/Sf7KnnXT1zMDn0/SuMntAtDPiA+2HLfg2MKPMEHti7FQ7D0SeMApj9M9rX/uVxvw
MbvLiknAqpmm2xw4fgRerQku6/dUt2RMLIbFNYOAtN4oyoqdos7pJ323Za5w4HPNZCtmgqhB4l3Z
a2Aji0wLiSKPvMV0K2dTlHovlhtSZuiH0B7yiXMKTLWwlMAHsOJXWGKvz/4It2b8A4dyfg4PkWvt
QbFkSP22ODcrKbt9hf1nm/FphLX0gpkxxRV7ffKUs7i2ifPx2uAfvM1leupBihZGWTMyYvKgQCQx
27cEszz9DxCZqJa+WHOvBoNUtZHioU5eb0T98h+qSRieiqyQwieldhiPVMTJzWOMzhtwfnrCzr9R
43t/rZZeTPSlGCMoBu5Kgg5HADuRtC4J6qPRmUuwfwFaGB3Wtha1RnY0sGWaak6ojRdUQlanSWyp
uzTLJeet4vlGewDPBned/ouLuVzKCXSerp96R+1vxIE3vA5AevOQcblyhxEn/Sz1FiksgFCMkd4S
ACacgi/d1kdL0EGjkmnLS22t5x7G5wL6zG3Yys/WM7Ecjsux9XBaugEbQX3FxH21fFStvCpIQa4L
Gqvl+e/OtDoxwlb9v7v+7D3N+deOEsQxn/YAmDFPzQetFm4NeBxbWZcF9IDXYQQlHqC5TPKa4KCc
2k0ejrSBYgiTD7MZokDrxdRk5zSNtn8vUKsFXGAEpS5H3pRq3a/WRI9SY7cs0aLKda2/5vbUP8ZH
e384+jBUnEGYss5ywI3Ghb2SjgVXzWF76G/33EUssuZ5zmwT7XllvyIJLPWq2yqq5Ea/B8oKyYYs
yF86J6dKoe4D5tLuNkhzh0b0+YcyQyN83W8ko0DNvlPJNDx4dEhhW5zVweBvBLqC9sMIXFnee9JJ
m3Zry2P1g87BM5aUvhxHXhZcFoZaKoMY9ii59lTcKj5mSkU09nIjXr7qa1kQUxB36WP+kUiNb25F
ZUHJmjOrk88jOpP25UbxnpZJu6cDdMA5MgMUTz81adlj7gd+Cqq1/OP0h5uQUThXXCZgF7RXGsI4
l/0Ak3N84AH2lRUm3FgIcxQB3zn5FgaM2iqNrS/qKklB1Svtdpd2Z2+eQxtipmZLIvC3/whaIv78
ugJmp5TeNjn9vpRlfkbcjd+6ru4r4DXXQkQgBlohA0PIolE5cPJLSH16XL1lNMQiMBDzdAAcI1iX
wHFn6mOlOs41OCQzKwExA96SZfgIV4/9ilmE41gq99qF4dOUHkb5TZOSYhmvi7PPmYbCeLZSCIAD
H5EQdtrq1VHLBYal3aa0P93E4GS5P5Ikl3dIN2NVX2ESrAiWD1hKv5n5P3ietyOv8WQA5SkutshS
sf9XdRV6IMRZAVlpYRS9+GLafUmwnK4NJJh++ruKeLnd3Bghfy9U5Hopg/ee10L09iVyRJl6Wzk3
8oNlI2QdvgHOGvXzqg4JVuePhvGtw9Pgik8mfoS51vDBPZwLWemrDZo1Zwxg5XDxXkwiQH6foYgO
6Vt6Qxl2hRTeyg2V0wHDbxaLAeT2EbDhFUF5E8l8emLk5eXwGQkeHEItmntRYNXe7opdNCEBtppn
TsMfLDjb9JC22q3/B3K4235hOT3BvGXchxeztRhYtncZO/4HeqAYvayEiIt126UegrX9aYzSt8xf
5aviLmx7O8FY/X4gKaAgnkblC222cMzNHgRFU4pP/Dje2GI7ayx+RN7643cGUFaHp56vWVrL7t3B
vfMOdIh7oS9YeHwgb267d8l47bpHi20mi9N3pcsti/IdUtX1naHe/Ylt4PU9EKvBZd5/8+M607eZ
srRRagKxpSzpHdtSsqxlVjaf1a/RgruU9gGwgvX+99fxQWdLqwKML31x8bADaBGss8vW3n8gOipW
W4REQlbpd9uYthpFOm8VfDhDCf8Q1yGI7iDF0xSWHnhrbvy9ImNAK8//u8FOpSDCRnO5tN/ZaRST
u16CCyuwRlsfzJD7yFUwwz0uPeS/TR7IgBijq+i8RtjzOa56NYE7XSvmuzIorEiqYLp4xteyWNQ8
5kIyxgbOITxmQEEdKTdWLwpWiqNebUFoARhuU7/q3Ts87WD0Q1xun/lEPDKK2Y6v3fsCr4JzW38W
F8cnEP6FHQJElIKfoXsbK528bEMveOxahSbSWhwPZqlMekwe6+Z3XGb+9ogiz1+1MTimJyKl/q2S
OzHFWHCqlagmftmxC66eec7DMzeSdRTo6rTI8Eg32ptJyuwGykp3KDsgwUbR+oe9dBRBajrMvRNd
pktcqkhb2ye77TDTjo6WHA5Dk320FK29FThUKcgzIkNrrY6xaOSFLt4u4EHGRp4M4M+L7iH4jLkl
tGU5tvgRJBFDpPAVmpIejqgmpf09/Fu71RBQnWYVMkauv+HBQKcBrHmTFkqJ4E73P0UO2mI9K6+p
OEJRq7/UzQlGz3prWCHTj7eFO1aBM5/zWVdsM+rAf1uMenNOYIb6z5/QEl1UPG0wHxov0Zw+ro+z
f3rH6jW1SKiBunqjvJRWwy7hNJW0BZ4jOhVFbJjJ5qKq5QPRZ7YeEVAqlm96Itggd4iKZaW0UwiG
4RBTbX306UwToj2sI/P9x+EYblMDQI5HAqE3GvjcUrWzxHSfIeliqq38ixRGxec0ByEEo6MYtKW/
5nlQsHTSEtEIcpZbEzSk+s1U87qn5vc5yLHxLgzan2BRqr6MPINMp2Qd+epqfil7syx5kK/AjwXE
EU6wMS3johZ8cCOiNPqUkSxmYVtu4A4jbPfxAZUZA6mjSmu8v1jN8IvU/n/CS+nmyNQihJB84PmZ
5YYjGVdbg0HvGlOSyhUlqLnZiSjLcn9Eads14FXA/fg6jyAyHTzhR2uQT/e9nUVQogdSVtah/oPb
CmP2NdVjr6cArOSLxD7A9nDlRkYjgm8WSiqlyUM4HMAz6muDmKROd842k/xEdTPBqAc2C60i281o
61/H/hRqsPI9/eIMKIdtEfYJ2vJZqEh2pG33lb6hk+2EseY29AcW36WPh6mabuW2uIar618rKKv3
zi5e3Zv1dgets8492qQpzyzwpPWUJ3wFVJn/5lCDdPWfnoPgDoKMIVaY3hr71bh3OBNfHb+qYe6s
GR7yriQl8rXeUDbHPrkPuGxUt5QxpFjg1BhVHmOKzl+jrLSqsiBQHsE4jSKKY71IirSUKc2r0F+W
VGUQHwmsooUUhJL8MTJ6XkNJhV2tYsxhlpiaW1OxQEqmp5p0VqnsE6bk6YdNHQKI5ZiBeD5I20TE
oB1WXRFjVDHVSbPcxj4c2W8o64ox765Oo67qL/FkaR8vjAz7fFxBZWW2Xv0rBUL839UNptZfn6Ak
G9Jg5TYkyyKtB0xlDHJf2bY+00DIZZleCxVeVVTzRiCEMT49GN2e/ZWjCL3OH4bUAEookyGo82es
/FzKOybX15QAi12M7I0aKjLwqEzYZdQ47jua4dpFuyMyztaPjAPTVKHVSvtgrrdXxJc00gMyo4EU
PJGLwWvutoI53rQ5cx2U6f9fvEo/GKKKR78QPmiiVl1T0Bqjv+LKN2f6fpTeVfTWp9QsDpS9GeX/
R5pdnWRxino35GbPdQT//Gw8cUENT1bv1I7wrDOdKsVGFBwb9wgLxOBQVhzMnNDN1iulnuo8ooEu
cSEAy7j24YNQWQ9kv3DFkErIujqVtF6+G+rudPQdp06dncjZyKWj69ectNSTTBx1XFsmNC4BUt6I
iqzwSH5WvsEvCQsJQ1qfZhN8zbu3UEWE2KuqbTx9f0vzBy5NpbBVuDscu5GvSk7DxzPOhwFuGBcP
TVGlIcrpHLIzFHb6qefyZc/ncx6h97safN+UnofW55h2pycsn/oOlH9He6Ov8gblfEI6y7vZbRNZ
+ZmMsajlV6r8+xoxWwgCN5JDJ7KuCh0Oe6l+NyXCfXdAIovrI1yZeppHYP2AvaeBBoo3fAxe0HFy
lq+jtZErDq4Kj/ra8OKVohisp6MAN0DYKMNcCfXYUsbhtiE+sVNB/PFsGsyqjLHBGbrCnk46jxA7
BlJF+HQuqMhuJXt4WcJ60z+4zE88H3LKpdwzM2SSQnRGi8U6PfbKpB7lI3lcMSyszBDquwXnpn8q
dbB7A/cl6OzorX+ja2q/71z42YXgFptKQ6ZVf7f/OyCZranqhSVu4Eb3N6phgXiZiWoTVSVJUaVi
45C0ZqFWimMIvV4PX7HRtUcb2G7c6MlJKhLfH6JObFI6aIy/hJWidyOzOtIOBkSD8cBbyvT4qCGc
YrDW8MHDKMg2sfaHjW3UGAGuiaVsRpTvTqXLQh0OUurfHOVO6j+4aUFi86unc2ZlLtJd8xpQBrAF
iHLeC0cH2MB7EL0aOwlYrnFRBWaUAMHxaAbrZry8ihnybebv47hyM+aLqL4dRTp1hjzmghW5BmMF
lcXAKTAvwAJzvSi/r7E8yV2s5iCYFZ/lc10rfTYtLOW82uY+drVLcHhmIsTIGJyre7K+SSsijQZ4
Xi36CKkU5hJ6HKa11+ya3w4+B5HkYsL8WxcFcgens5GJQ9kHKiTti+n5bIVllO+DKlfnEx9Dip13
romCphyH/CEb6+evgsXw2YKd+fMatnklCC1SIgId15LkzWVMfRbQCcIcbUHxwSRo7cI0tapwqy2w
EOFFSIv7h1V7Vb+vVx1f5MggNyojBEF5rneBCYdZmG6zjwrZ30tRj+3jYP0GHSbHIqKcBLEJrbac
IVZI75hE1rclBW6UgPJbeP9nWm5EQYwHmQ/4zfMmiERKy6WrT2O7PWAbQPpoV9ZvLJtqjRGdWEgZ
GMJBAskl4Ij9Rt4bOjPfsdPA6x0fDYV2ZF3ZHHJn46YNvFTH8Hz/Q6/JMj+Uti4FXFW63/B+k626
O1cAQ+ZTcNAT53dGcC6qNPINRhAyNluzkN/01L+/AUjwy+W7BfR42JPl7sspu6S3jmoHKfHIpuMP
Acxe74TeGWqUo+KEbbQ0kODrZT22vHwpM+ZcC1yB17mbcR9modIrqk3QX9WbpBS4cahFmcUTr5gU
9TJc1Wvlz38MG/MgAAKdDw7gNqO33U/b0cnldoDt6nyTaxssG+lqRhuYFL+JWHaHhutEIHRgicMx
qFGGCle5Ta13JbeTMlFJAELepxkbjo+6CCj0w+/rHi0vQuCKjIwg5kDN9Ey0EOG6kRl2t3veCPE3
PUqX1Z0eaIIFyiq0Mc68zzFF5nW7fFaLCum5GRwtv2AliO56DJhaUYuXkOLvFw2d55p1MxqlZGyP
UD7hYUC1I7R8joUbrCLt4WFtmNdq8gZNYbKzW1jsjmABZohQkpBZKZVVag0PVN3WfJCjscSOht1+
Ej3kmNtoNwHAvLlAFVocia7ZMyLWatc2KensdJ7pS5FGQS2u72rMarMrqSNdpN1JN175CADU5k61
0tCqB1SktHF79JsAKW1Sl5cpt9mQV4yuwki+H8w1gSxadUOPjYmB7rBUoexIe9XjChMuQCzpUgWr
+srhZF1twdEzVx5maht0Dl1pAXox4WXUh8bob2n4dFRdEFep8QPv9c678NQIFbQC7rf2sk9BRrDo
CFh7iTFScHXOoZ5w1W0d/BgATSl05QHOgClNwA/lKt9cp9SScdTib+lURvpyFw0AGMA+iVhdvbP8
72aKa7twJUGQ0ZdQ6BUphKX/BOeFFLxewQMtjBf7KwJlVTZZq34ugjA5x0U6qi05zE3cQjh1iiMO
zlY6GTndsmv8jFsMlz/iqAPrRMzpQC7JWZjkzlx1lpHwkTrr2tq1crqdhbFeHzaoFblmGsogtRxm
QuF3xmpM+wuTNr/K6TTJ+F+zaIZvuWkJIsO0PE/WvC1bhIhbQmWWP8WhnO1rclA4a3GaleK7v8wd
gsEtwqnnbMh9LITm9h22/Axzg1xvyLrUz4o6RVuEEV8cOe6ELpi5eyaCxA/nXgxgkgdW3mdgSlYP
WGRIDssIPWdzOVIG81IbH/5sBdlFPhD1OnNdj4/Ydbgoca/Tgp/IZSiB2GWLXn3qWuLxSL+sjNEP
hd8vKiobrDQhnEKiPmnhh2PvjMabG2qMnEBVZbQvI2kqRvofpIDIireLzZoun3K6weUClvPMH5U3
8wKhiP5FxSHP6cxiuwj+VMHgMUknRurNiTDHutixepgoUtTXGCKpzgQChdcmDg64/I9xYD4GlRlS
tN3+1KB+vJ00sUtIh5GVS1nh4oO5eOLaXrzcNk5gQf4F18JLYRLeZy3fn18UC3RjmXgLrWpJPfb1
3AWwZWr2qAGDu8eLymtdyRwKYfgmvCEIUzYSUJgLj75dYvwtxzj8pQ2qNdih4yrtTNPkOGWJRS44
Mmh1dBda7c5ya4MJ/zej3PrkmtxRzpgGsEGbNzmWFunuxD0uCnwLcJxLLERCU0PQRmCpbJOrQvKu
vSTNsUgwfmvM5t4YT9MnvjO3CxPyAY4tpsKvy1Li5pA2A23hCiRsMVTY2KDVvlmYxMTKtsvfqDii
i3D183xSFiSfxY2Z8IO8GPLvcGbe1V2+0yRRE3GCs9KhKBQTapAHqfao0PP52P9ZFFK/ONrrRene
VnxJ8XIYK8o7mprRGTRkA5YVDGCLmAm/XSb6zGjBXll72DKwSLXkrr98F7ihY6mFMhqzUxGIDL8q
mHMqNaGqwN/slVdCjO5KrvSbqTmX61x+yZvUh3RGPW39ps/wRSKB4YxgI5G5YBbCR95JZxDd9J+D
fu+uXug81Zx8T5ekMn81fYywelk7QTV15EZrBtlDTnVO2x3rZuUi6aRb7JYtLuc9SugO8PcmeDOd
Xs3Cxrd8x0qFs3jqJVOf85+bfZPkXp08TEhk08nzK2WP7DzqGALZjpBwmDl40iukvCgy/CjAIrfL
SL9uDivNBBp6EZh9HpvfQ6sMvewpa3mlSIn9v/YcPM2Yp0pHRrQIV653uSpxeqZXxc4QhWwErqR7
dOdQM870mKepMsaFzAWa/3/ZnYjcdTgL8xw7OOIP7NZnsAAqe6sRGHSEIuqFGvHOxSAzjWMTgkMW
ccumdXZrsqb4ZywGU7FgTKyfe2jvovBr+UhTyH9xajvtzDLO67jJTiVdHnQeiTFC+AGEDBazrWgQ
ZpIjucKE7VV48BIgoCPyvEAU4m1YSSsKv43eopi8bZGdj8thuiE4qLk/EZ26Qm2xJljlA+9VZS+K
QGcP2MmFi51l705HFAtchaEzWfJTCMTIC9vso08+BkokiWEFpcddtf7TQSy9Jp0ke87de4GY+5np
QD9aSrjHlDIQ63nuKQpT6pjwLmosvfUwFL9HQ3DpW4piLofV8sjV+XEsFF9ntul1Izr751+bLLGr
sT3CODUkkrsvU+zS+6pS0boqe3P0vL9MQLwPNKEBLZvr/KTTHKOY18ZXaH5GxmrHHhoGsgKeo8ld
8HpcFNH/POyKIdDXkJeIbchsRbRLdS0MFDjMtRDgLrktS5ggW0kFAwqblMJ90DHGbcvKRPtVkcSv
udmgQUKAfMjkTkolAjMBdiBSeXP56OVY5oHxWmQCzMJeMU48q5K2eA8bBuaHB0C8TDLySXvpW4vK
zU3F3cH91DSCHoOLNuBjrye4Fm0eBSGlSvh5w6B0gWQqXJ1PTdPOQ+zIRLcU6Uh5ep4y5EC6kKkz
RSnAS92ng2kNbV8Lj0Gk7rU4S6UgNCVZ0DlfZjJQ5J/3pkEjtv6iez2jsJYfpRtQl/pUOyFaZLJz
hdhl7jsgl/8QzVIvDSqPyrN3h6sCP5PYOlMfcVJqLzmq/JGb4/Ly303XHNTxCgmO7/KAh4iM5bCv
1u+Cmb4NqPtYlAZjGhQ0B7NW+35SP04y87FNzkAMvvNj7r4wm89oRTIngycufEdtOhIfTxKEnrA9
U9loQTua36FCsA3CpWpW/UXU3TrtxlFdseNYGKJcoL02li9+9L1Zxtr0EwpucZ98pxIEMssbrBKd
wz3XH3Iad8FGPbuUhZY1bLOFCfUIgnpB4GytvTbBxqvckUKe5oDkuUmK5KHhdajopZBOfuCpCR6H
8tG3KtTASNqlsYkZwL0SdzkKOBsfkyl9c5li43WpsMYns4ndsh373032ktlHE+r5J6Kde1VM9IVd
IQkNp+DPvcAlSTQ17AnAByfojkknJ3dWZSJl9tZCmBQGlGSnHkwEgnRFE2fm3RG1LZBDN/GsX93X
LMrrvM58mw1fqVhBiJA9364a7hfjpJ5b2P8SLTL/YDpt8CQrxVoiZJ8pmx3/iBTj0+soJSoUB51I
S/MPvMJ4Vsmg5r1HCkzrbN5drgmzAWPH0I9dJ2FuNaWzmg0h/ECiFQZN/fplNkObdAPzSr5dVtDa
FH+FyZKhrPL2eH2k4tTvBkWZRX4MAfXyzi2P957mM9Aoc9QT1GajoRhNwilGF+Dj5/sMP/KXaRr/
OZWHmj4xMW9tuvDOfZtXeKYJZeanKtk9tovsjAuROuRhYywLyXz3EC3suzbBP3kE3dYocp6UzoZ4
7g0Fc9/oYQHsFxx/oBtvUFgBJKxEVZJWgQc2yzah8Xwb2inUKEztwJTbr9ltt/lZ6+W+dLPB2YkB
YawJ7qoGoTY0hiekpe4XgzD1Ga+cd8Yl8qKG7H4GikZlnR7X1wDACFSK/vK7+qcvD03usOXOWSzn
iAwUeKIOaj4RAZzI5ehRinlKv5zVhPi6WMfSRqYbULGUeXko0J1LJ6NqiBfc90/XvsoAczUDSmzO
0QQzZDeLdM7xcQfbtiiFWxGCOoiMyuQnox+jCX8LsaL3wUM8rYwDlqv2C1ZM2lUAzA3eaeUVPdEK
gGJNiLIhDWyUkfUovjn37K4j5NgTkNIjmELBZJhejB7AhsFAD7AR62ngS6td6zFALjtm/wq7HGGC
6kXYbRKFBeCqfHmcaDR4O6kpv/DRXUxswAez/B9+Vw6mLPQjOpV7srhK7ksGvvlg0ywh6dzYH0BX
9AtdGS6pXU5xFAQ9BmRVHIAcj+11/80DwZiVr5rjyn1pghJMs//ow6MU85jGKbBzAJemTaIFt4A+
k67gv8ClAe3FdrkgnNN8/WOMxUDKyP5wMCsA6Jzr8FX+6dOroNF+bJ/HejlhGDPQOg4qX980eY/6
+Zplc0cvMmZjUpzT+T9zuwIalLiFJouayY9HVFD370W2UT+Vzm5ruI9W5+apW//gFxAcrKvS6Prs
MwSR60cX+z5Bs3BrVy1Ym434KQcLytS/xYOdgTXfZ+uH7Vj31/caXDwXV/8LAuussFJtiw6p52IL
cUWIYiGorJAiNI4Ua3jMpFKQE1ba51TLeW/nD1ANIQw6/MJYwx/9ImnT1j98zCFFV86/r3veO9X5
tYNak+lx+LpOD+iFBSUuxK71b23XfR5qFgtH9m5UReZ7WYn80rVB5KHrIYZ69UO5Ruhj0jAV07xh
nLNW3BTZBURUIo8y7dpvsTW1IeFqngfyXz8EqdTgFZMhhgheyh89s3iit2w483sLrxtjDSs9IlVR
+ZUXccAJm1ea7oRrMzFdnnYpBAsbazVCO1s57PP8YcNiIP2jZ7W/+3Y2tGzOGf26NKaISE2nF23C
BzcGZpb8VvuPIvRSOLf9GCghvTTfZPyjrDwMIgaeKwXhIDVo/n4oG99fecWDRNvJQZnKOhjy9I9R
K1ODANpA+6hIsc5bHPTjjcfmu5lOIJer/2+fH1YwiSpl7CgyytX30qeTf1CB735TtU6oxT7IDZWT
jHHzWOMXOPF0GQfZY9sg2bzElzJoxAm31R7J1DyhS5AK/wS7XpxVMF2O6lxV5ZcgGymjfUZVYBUx
p3I7QGprn0tNikuekV2ZBoEIo9sl8jfEgicb+eG36sYT/4gB7n+Xqw4ax2r2qfFfCJ7dtvTN4E3G
gJ2HStZfuifTt8nkw1LfLFnFkQZjRNYPi4u143XmV2vnaLNJdp+zrxUlOAvsdFVE81jh6lW4chR4
Hm40OnChOaYjXydpkFEvZrUFSHUCDtf8frqKofPHlwKeuQcWf0cEAGQEJSr5NK2TFNLvPWt4fCDs
Eec8p1BRhhApaqvauvu3fWJHpa631OjYyuSXtzZrM4TeD91nk/BvK4BN2w7nGJzd7rHuPXSsSVVT
KvIgkF/+lS/Wwo8wJ8apMu2Rn4ZTgWLVMn1cpPk58/tr371UBjQfsCLe6cpBhvsxTksLPseHkeco
rav5hukxJ5RBSe6D9P0wrZR4Z0qHgAUVw1Rqks/l8RmPn80Rk8/aTxwJ260dD1BuFFFHJQJNRUiH
v2toi6cODn8P31SDRHAY1G6ibygAzEnOXqpWVVRXtEq31M0fQJy8zh0BDMyjybw71HM/dLBk6mMB
BR+nDjbSITIiYXO0dRM5FXmU0bBapxpch+q5KqvkXOgYa/ky/dpHTGfkO4mEXf3PYsp9u0tYtZow
qhaRIbNPC6k4cYx2sVBFlMWY5FUEalZWe02i0PP9IXVFJ+q2Q6PRXvOAn7Kjwgo+1Hsygnj5FLls
FqkgnSPcPLziD46ZNHbKFqkY9cg/q7x7UywjkekQTqpdcYxyxgOAwYKmozF+pLNRiJHfz0PmBRBi
izj1hoHkZxjqjMEZ7DD1b7ATVs3qntzRZli0tm1L9O4mOrwFK8eAeiiLgKlWOIPMYOjdrQm+RpDC
+R46v5FIiWJSvLJG4Sr/dac2bk0d/RKsFQb5fUu5A54z/cdZwIOVxjE62w0UeVaQzAV5hyf9ja/O
jj2xrxHXJAjVHFzCRpaaG0ZM869K/8QMAYxpMZVSXB1YULvGuIWx1+LLF0Ipgurgv0Q0ZddfJQQX
Iz/zWAl1lGFvZZRUTv1I9VQ8tWyzd+lr0EC1QyLxPWaEkOLOFc58gN0jrDOEsvDUiw/yWnIoR2ZL
mqGi4goYk1ZeedL9zKAuPTAnTz2WYX5pD5YyfrjAbHYyu1qQJcHzJgpVo9c/tGPazjnnCMc/ywMs
4Bx3zy4pl5WuW7B7j0fOpR1GiUb+e4c3Wc0Y8v/1k0ZWhFPY+bhbakGwxk24VvC5PUceF2xGe2dD
wwO11QMiqrzIhgL+U3aelgsXPqi3nPQBDlBGQtclRN54sT87xEFKS0HlyN4y2hBQocNLpI9tATzQ
CY1ZnUNcwGe8IcBBcbh1Mdb3mq9S2kZNy1egJvGQEXoQIHzBG7Gn+sycPGuFxlMQwowA/psEv9I5
OfMCRQJds923iyGRCUgqnOXEblFI1z28AV9UWPsZc4xoNzBjcPkfpiShyD2j44Gw94ZiZHUTJ9dJ
QWzAVwImd2Ic9FEN4Xl4JBk4O+9xMuXTiVnMaSlPzKH4BY5bBI39MrNgxUiWutglKNDvEKh/AQPG
njdc0XdTaBU6/HLS+sIgwXxEug9DCFBtJHzq492mtYdR3E/FyrUT+KeO9wqIE8zHkZYP2VqjOtHW
C+qvSTiM3rd78hEFq76jSP4L7hAMmEOupr4wbz93/DqMFt6JKY4iq9S9ymwCpnKsIsVlxO0WsuFv
H28MVguAqRWkQ9/uaynfUMmn3pfpM4r0qxc1kqPku/i44kb/dFQ7NoIceCUXkitOH1siXPHsRMPL
aHg9+68zux7/vyP41v8Wq0hVYsEQTr9IWHean9XbO9Hl8xEXyB4CXc+by1lrKWXGDdJlLyF7z1FT
V9N+i+8YMp+3BNOa4OAz4h+VZr/3jaUNQNxjE8cBJgGTfoIJQzjTn0ivZkjKBXJYiHbvgQMk+j3t
XbYJ8vihjU/04J67Lt9W3bDqkVE/UNrBdgMpSSbZw1YEH/+SHH/vGYdQsdfVAdjoQ2IwFznfvNZB
L3KiMp+iD+GGLd4WizzFl1ec8Kcg/bzBAPA/l4SiNce65B5OJxhDsYLAzABadt9DCbTk7VmAuR+p
GPMVyO5MSpXOhAllTGW5nRFY8BXeI21Jy6RMqjUC4LmuSNpbOSckblPRy7wU9kFpn4Kj8UG9mx2v
+4FxAa5qSuQ6J2N/FOIKnnMsDXoD3Odkm+haTLFgn8t2U2Ilq2gh9loQgDZ3Jl1q0Eip1YwbGDtM
QWUjvVzKtr38T92z9L/uLRfLCpv9YJAA5Dq7jOySgVAdM1kF/1qcII5ObQ79AOH1/bi3Ne8PfT27
xx7LbThZ6JNi+2gcWM3DKxmrBj3HfdR1tFlHswLtP/PBUBztU0SZDNUjQgnkypoPNjgU6ZxB+nq7
NELLkYZehGoGZFtcl9JMlpqzemtv7Xwpeh10LvD3s7YH2MoKLc3xBAMHaGlyEkW86M0FG2JSnbj8
eh5l0HligpmUvgJ/lKOpPig53ux8t25TMO0FFoMLk267PSXCveDwsHGEjSjo/Uqu3CmpDdCHqSl4
7utWiAo8x4jzzTRaVN+4zVLiVrTBzj/d+OIsjNtFBq2YJ3HS7+AtrJyK5aeoa3NvAlh+BKuZjjuA
RjurNYCQPWJwxh+zMur7UBTJOAbPhUScu7UL3MjJ41fadtEUddSpHrUVDPrGRt8m6bZIoXLeyqtS
m5B1aePyo0bmU0mAkmvRVJuR2dZ/PCPM/GxVzuEg3lrRo21tfrkdW3bLGFGhfj5ZeKrKmQGMYDl5
WIglhRhnSL/Kd3rNCA1K+F1higO4MF4nUNIU4sq5O3Puvu08sBV9Hv8aZSclM94EbgbevmX/RpgV
N9Dn69LfpyicIhh1HSL3Y9jZZr8ustczDxuousNnESQELtS3aTANQH8Rqz+qas/vNsD73EDDQWDU
8+FiYn7XU+tDcRaN+rj2FPHHO+SRyoLC7rj41cRy6FpjVoKbAhMDgYjrGK8lPf+0SDKFMOJ6NejR
/rDoR7/Y5MnySrhY5kj40duWcQZxqgiujaUfu8/uo4ImyKKH6HUnOOGfx8VdyDIkD69/4/mc1rdh
BfkVcF/eGT/f4+8rHuGmd5kk32OE3saqfZiwUUbgTN3V2SV+8+ytksJ3XXHte0g2RfDi6/0/l0QW
VJiJ9FA67h24akkTzdVaaBnFKCotfwx5GV8e49yezk06zT2yyNsRbI60f7lBul/Y7poV7GvNQIlb
eLpbMMZ7Q0n06D9n0U61wJbos9JF6G892slZt/hkl8sQM1mYZqQ3fzMjbufr1FXphyip9GIAmPTl
YH3KWthgWa7+JgeHvtokq8sISztB14/7KGtyw8MAdvJKn4fvEtazMSgawCgso/Q8lari489aukwD
JYLnEr5UVOHAgYg9ZiRNx2Ax6R3xwOjVhI8rixpo0g4w1O0lYR2MIb1XFqu/YTQmZ9FBixDHnFcK
q+6ymK9uJF1VP+VYllICdStt+B4ujfoaELUU2cL1zi86bYs5UNu5Gpk0McPnwRIyxECvb4yB3vkz
3A9aYmFje2OEKnk7yu0lEcGPjEtfAQktDO7a5uyClvtA8a2vR48YvEIUST5rPUwy24uwUVxqhVwk
5Itlwq5R5ny3E+9ihUZmquX9vcgTFLVuQSOulLEs+HkvS3glriJi/Bj5xXFXO7s0B4P2Dda1S7F3
JOvWF1a9U+PCdiU4v7V3hQEzPKNpjJEqSwLGArYWrJ4DWokPwGB3G+wnZjFGXgGcjtcscCMZ8B2z
PfSbUP2APCpfdmJi9743MFNmkIb3kw19ny1HR3ERfC3W6NjDsnA8B+y72Wv275z8XJ3kC5ibUwN/
DcaRyy7KlI9PCt0D713sNNDgBEdfBKtp9x3gfcvysKNOmFaz+O29hdcZ8Gnf1ASm46cxqOgLr5ca
BbbXduBM2xnFDCrJqvdRJMqJ5PRH7rqRcsCan4INAYdMjbtsOFGoP2pwtK/EMjO00aUFX4UaoCYd
pTkakCvRuyusVb03EQEA4BkcJ82deoSNereWSUW/Naslw6wKyrqVbCth3JTWGFG0ioQNDZ4kJFQg
vgHY6FbJxgaVAD1bYAVFh4+ckd8B8j8rMMzlExE6FH0Hwizj1SQYbSvYuzUctimUgHL4fKbmeqQ9
OVCdyqweyWnQzC1J8R2I30Qdm8gkUKuWVzG1NnfIs3YSc6fpkYYY+kFGbo91FgdpgPnIICZnU7Rh
Z5V1qi8myHvXLFHnu3TA8k7qsoUulbfO/eyoq0hN8wsiTeFeYLPV2jlaJid9rb8qs94clZ+hLhBg
GLs61geTRho887gXM3cbRboELr0+mM9QjTQDPYhBfjI/xztFhqOkbU4RCJ0z8Srmf5609P7xYKMs
jHfymqkbCc/LlHit2eQjkLJ99I8GHY8loUMudpVrCAwcCAbrW8vK2MNGToZFIq/ndPLTeOI+R53i
ad/E6UbYnKvsrcE2b9kKFy5gI0Nd+Zmdvg7hWGMIVkRwxa0CsAE5FAh+CgDA+FIbFiTPvXuBBn04
52qZ7FIQsPvw+KpbuKJVj26rwJupmmRMeZ+7yQHWwC8uFRV6V1FwmHjECYqKWVrWGqRfBJFFrjI0
jMOIOOgKy1mFhxDfofbZ19jUj+UHEwgVJz+smbGk51F1qWKFyNhKSyOhV9dWdSnEnpzeWlXRKb67
xqAt1vaWMeZprWhay3zVUZ0lKGHEP4euMlXDJ2zxuYHTI0Bpko+4O/WJZ918wWYmn5uTTHbNc7dG
09L7bENhuFeZ57xYz7maGFto+9vp8r6tt9FxRZMpkFPhe8X5SVtz3U8z6sABm6vgoyugaKBUFPvB
FXkJEYIGLj8cADOuUSwPxXRmm+MRPa9GjYOP5HxyhTlPeDoUkDMsg3IMAdkXJb1Sq7AptEsPwMgs
fcVOL3X/K2srUUcVTltrkU956usVYt4YI31TEujUd2PU9crhBq/wLBx2VSbFFZlMyprlkqxWcLuu
VuTliaTmuyGfvofZwztqwzJU5EaUM37UURJjS18RGy869o45eg5HcqyCIgjvd0GU9x63t5g+I+OJ
a6LGVIuYPJZz7nzlBfCbG+f4GQobsL/Z4zRl/vLSkyEnoBvndyrlYCQK9g/nQ9AZkJ7Hd9ydmQWU
8VCVi4zVZ5jHq5mhIpkCtgutbHpXLn9ltxi4iSpxDiuz69O2wYieaSFsspNSgg0JaxDJFbWa1umB
mjRfNEFcoYFAf+yLBRW5J+9HL0AeMRy8dNvkj55hCnhpHZsTOi5XEKh96UCGsSgXtERVkWksMJjJ
viMuYK+TeQ66G7HUnHEE3NiHyw7MZ/urW3hTllKFuwab8MDdI45N/NXNm0GqZDfUL9WfFzJUyuN5
YlZReeoRi5QSOZ2xuu1zGjePNdHVvDmQfWrZIpCyxIXjoO4XqirRVPN39a8Sj5TeLFAFKZymeOuz
Gnl/ai2d6Ci++LTjRqm7rmi+jrA8VisWTjvrKJcLwu74YCxdVDr/5Man00Q1F5HepdOpoiC5ctMo
bthEsVZBAY4lQ9EDeFwJDajQfVeFl9GNQDkUhEjHJ3xoqpJafwojZhH5LpnyjSUtT2n5m7UtI2q6
h/3n1SNTne2WOZqyPbwvPTsGZghB5V8YoAyZ1CcLzH30w0gBDd3dSoVzyp6ujz6KhDiYbLCf9TSS
WZsjJfTzNn+vtT6kbqWnRqx1pvn5fqghn9TeczCnQvr8NhgMOVeItMO+Gu7XoSE7tvPyC+8NVwoa
OjTF8JyTbVC/sY92pTZ56HTb5J1Y+6S+pg985EZ5+FGXtYlMvSUuRmHI1Hu+SK7Cj4DC8zlT/+Wn
oeGrtpb/GO2j3DwF0BA/XcVOGieKvXexnWKyFNV9Krcsz245YvN2atX1SdiOmC13ODv5quA7R24r
s7GRZzkbmosk/XUqV5UzphQ3gT0NMHxIWM341th72fQZZw+7fB6hHGPREoY6P9NcbM92ahWUNN2R
THDDsJLxaeiP0SyjO0e1ziHzjsEdrYbHHne3tPnZNJIBG840cmd8f0EFUhHgL769EAnIUu9P8JQz
qipxrQBCTgwIAr5iDXLJ5fZO/WtspapW9PR0gldv2vNiH7RG07reCAOef0RSj52P/vtKTQH1yLAX
xhqdmiBAOOESdrTr9cI26E6BxtM74j0+KLRaaI/W41cfih1Xyz9ofyTR7Ztt6D5sxld/9NUjPwCs
nfdICB0U4k+6Jb/XH8lVnZcnnprEicl8wV2EysgjcOwc7BPmrBIkxvJdSKUSvu/N1QG3Jr9ellAh
+wpIiyKMpe1ssfbGQ6ZZj9U0azD9f44l8zpMUUf+MRm6Ls8U3X5UgYxfB5T0De2pNs5a0ldOYrl6
aBYvGCONv+ob80BTUfudMuFAkhtW1LLJkaMl5U7s6u5kXxSbJ4LVfJYoYqOJNO4fEukqznc6hXBo
RTj0nZLqyLCaHmTdtZa1QeOtkRI/qXMYHlyMkmjYI9vHCJ+TlOTs9qt/3CF5ruxTTvf8svjpii8K
P5uQHJCThUXcgbPsIXjn9cu3scmM7cJuFEi4i3KBZeUJdNHQYXOqdJmRXawPAbFs/AwCW9Z4PBwu
u3PjbY5AILlPI6IZssTG8ucFScULYJnEmaohv5vdtZwL3ieGyxwnnhwccbA0v9sgZE5Q7H/6jfse
p/3145NVCi750VjaHXYFcOeb1aze505zkvPYdNGR6QDdc65TqNqjugmcK7aT+SSJ6i2F+0F9ci/0
qsHsY2CzH49+ospu6HW9A7wqpgj8Zt0uFzZ43NRBrHBu9DF4ct/yiBSG0dVLow4PBJp6ZM6+ITaO
Yv0J15I/1nahez4LU/ohzNHaf9NNPa3gowA+6ICCw0YhL6kkMzOij1X8oAPQsCzvSMX43Z5Uy55N
yqY76SuP8tUfgOyrSgtyPRXeit5bDj/FPmknWOt/htJ6A09cDQllJ+w819OA2sKzhiBUahdRjFcL
BmIwDiMYd6hKNfvFAiX7MdKkBTCR1IbVSOIPTE73Ic1GkJPpG1iHphm83jTeL0gOxsFT9TorIpjN
AEF1sY/B8Hl30HMwVgx4A8AV8rqnXM0Upha9ckkGRlo+m4GwK79kVSSTdFlsqtXc1vyyciKP/UZ/
3GVZ/StTYdQK7bPcMUGNS1lrIy+ci86Xznioq8RLD54hRckyoar+T5+1D+f+GuYGQ1BSCXXzST3t
J4sgeRhkGBtugsn5Q4fu2JVOHrSMoJ0sGswz9QoBAPyvpMLhy75+MWOoU1WNuZK6MNcLVABuyfnN
vROLEGAwzXEmlIEmB/voYUKvChvRexuZ+Z5drmdRrcmkR2kXHTGNHoRpsklEByGMQ2q9vC7MtKZ+
L6pYeVaPXnvZbe8Y8U8QjO2ipyY5C22p8swrDApja0HrYQSut7frIt0eyT/V3Gy90/7x/KVrgn+l
LFdmxcqvPaCRHX69apmtioVVkB7PtK61B/GD6L3ui1iVTwbOyhGlEi7xQISWi1dlZ8dkjZrSgQuB
eaiolZpIqV7e3AeVG15CWvaHGMf1XtGNXq/5lA3bgb47zBuSICPvi0SctqUV3Eq3PYbWd5M5hntI
VDFGmvqGG1eLxMHfW2DAf8B/z3X26iaqZuuA0czepRRo5GyW/i0hujO5CrD56ZfBT71SEzxNMjp/
ovaQf8ncjMCnFZTuzZhDkXch9P73Mu15sP0A9TLITXzAGp9NzOiinM/jSWfq1Baj+JahhJeN0QPK
NxLK1oavfT44h77lDi1TokMo9cbiFWhwU1ZOL91hmNN7THcZhGRpD6Gq4/J/lRA2SRW2zD6V592q
eADgKx5jPNIkeeOeByWLLsMKkZMF7EEwm/1dPvWcWSYI71CELeQOEeL6oY1EHDHwDGGY3z0TNlL9
FOvqQoBDUZBcKN69hG5e86CQNeqsZyvEbnNhIHvlF9dqO8f+/B7T9kmMRu/rCLh6D5TaX3SIw+NR
M7Hf6JfT/Abn6/x3nMasUg+pvA4C3KA2bfGsiZ3K92x3LvKMuXlv5xHa67p2qnOZnf+BdvA6eaH9
EB5Hm2NQyNQ6a1WPrjkLaWWPjniFFG6HmNckWqcxdzTeJeRRZdw9kavFDnW9n9EpRmKixyE/08yg
j7jV+xRa1mQ7Z6P3t4JGhd0R91/bTikJIzr+PbiN97sUNeJSE4xy8pXQk3/HHpY+Ch7X609f/UEx
rCtUj7lQBCOFls13F51jHGaZftWcIEVBxbXycPNeDkxo55Drp0otmWLNy7AH5L/ySh8vTs3qWH0B
9wnH1abb1YscMtogDKg1z9vFZBMaZS98FyoYevQ3mfKqlL7LGPknEJwRmRSAh1v4tG5eRN2tA7nl
/mZZLu93MikvWg9b5mq419H1pkAofw6PgZ13o0XjjNK8FrcEev2ImrP3S5dkOulBg8S48PwbfePA
qz0qO2zgxOcNI6j5DUkEVH4lFWydRjwmaCu+s0KA7me0X+j1Owod+NA2ks4hz6IlXhm9MsvoJYPP
eKz4SX3R3t2+RVDY4cYhRzaYvGnp2rhHyCPHGwn5Qb+7C9vz3xYWxtnfVWrzKRh26nN+vXW7YTjk
o4DlNqm1GDXfLBSI5hYF+pMwSF1wjnNcJhc55R3iC77iEia1+zh6qY0gOL4YB45+60aC9lN2/5ao
ccDXR9S2BsbjEl/oxzypJFsVEFWmAg+v3f2i1qtofnZUHrjhMRQ3z9VQqs2Zw0GMOj8HZh8bOU72
rLywMYJQIMSQyHUhFVi5bYkAxoVTR8s+dw3389vD/IW56meMuTYg98vJqPHhlZGSwFsYDgk7QZ1r
1tRqF8ZMdae/lRNF05RI7eRX1lu9NJGc3JmO4BesEl+4VPrUs7TrDb7hMQ7AhR7pm4Eob5V9ks0L
v2t/tjb8PusYpiFnyTBWrWirBBxvHJZah8sR+4S89tMaWrDTreOnrS34aPgMEIurZEUgm0p9vZcz
jqKNLowUUX35gkzLhzdGy/D//qgvsbMDafFGbj1NOsd0ItttaLwLZo0VF2zXcECTBlAoudCZAcOt
+NXh429Xde01BDh24lqaTbybgwenCwN6n12XY2gzJe9Dzj3U2xGVlmPM6glWHG9rlejNrJv2008w
bC/Q9gTwGBBLS6BkQbHJ9fu1qrylWmlT6BcrvPlTv1vVZQXvQTuOq2XRwXWBHDP8/BKmI/qbQbB5
gDWmyjcIDRmDXZ8r6OlWJYydOOQt1u8z97Cw/O9VOQx//MsbKZ2jI/Yu60Mu06J4IWkSooGNTg3d
PXme4o4xdq/rCP908jgQCjhECrUaCWmV/S/YUW4wIOwz3wkcgJAbrpbVRTnczLu/ArXyj4aPPLsJ
ow+YJDmgH4FnACk6YXe6WJ0iZSlMDVXG7cYYUg1Z9wKmb1ROaUQ7AjPG0PAlqaIrJAysx8ju5pe/
P6OFSBox/Jynx95CXkZO7drIDgup8XWLSxqPUhc8q8gxiPLw42kf3IpguPsgdXyIDy5o0puQ+2TL
ASEAo20g3NFTj8Mu5j66yPqIMCKIfj5qia0fhzEo0WO1BFtf4xKzROVLEMYG+BW1DELvtYX9zQza
/ufn71yI1fkVfVjhnS+yVu1AaGAjmEiXK5ZDmeolVHfS/c3EvnWQMqK1uZ61Zy9Izt1MX1iVbie1
rzZSVpCX8l/8hZSU25snbKeaxSNsG3wo1b/PV2hfYaM3sAEEw4JdvQULv73ZGaEvjWFE6yBbEN0R
CHP59Sj5MNkvy0HidJUtvl1zAoRwzmb1WaWW37Ha2pjWUvL/iAjsIVhXywPdjtAA9V2kmicZkiuU
CSbqb6jHTymt15Rl8gQK8wsirWVxnsiY6ieOIpzVgcu5dabNyzkimV6YTFy2LKtC1hIEImuyfTrX
YXSviGmiLTfmw4rmc1OSep9yDwjtdb1jwczWxiojys3sbs2L3Ky4ssPeZihNtp/VXlyya4Nzaimw
2y2NSkKh69VZKYi2eUNO8lQEKB/9DxR52iCOgTKRrioAoMHy+qLnemjTHQlbUsa69grRylVkbFbk
gNlxjTe7MbmSuEJVGnPdg0LlwzQgdGR/N8I1ePC/QMbh9BKsJz+iZa8EF+vzDJYGn6LpO9E5RdaJ
yUwO7PYiEPVu5G8Ign5leeUxJ2Q04dnTQqccZKK8fJIg7NxPeYQ5UeMLB2iXCY5k1vus5eaPWjE2
cZaerrf4/hwBTL52qx7UCHsUPVGy7V8WpawatrHgoCoZ6iF4rla9Vh3LoAXfWTgkpzSCJ0KU8gFN
fTUeSxzhqsMBh+VJMG8l1ZK7yBBxJs/Fs4bgfseI3cCRQ+GGpDs1owLfUeGQSUS7t408dfQjJ6jq
wz3hJV0/l/peD//Ux9Pi6H7Mh5k+9hD6dwpTxT0Va6eiSH4U8VpnKnWJ8qDMXlV4cSbok7xJZvei
c5bRre4X+m3s4+4uI9XqA86toIU0JXbFg25+ijeROXq/MDzPu/B946ekspRQgqAkjve97MC/WF/p
+awMYfgq5SgyxuhxdirEf7C1Van0L/SLXs1JmtYEHOWx8yO/j0Zm9/qatbIxT8gxhVW6Z1S0dB8m
22Q2WVbE0zWCbW8TM4wlQHmT7uawCfojL4geleeIIK6MTRmdbkYM4/o/g0NqEVMnvK5IIvzmWESU
HVbgR71Gi6tPEOkRJKlTGsvGEPrmkBeDWYhIH+rwSNdHe/7VPtcCu9u0Hwu/KlUDJoISLqADjXY/
omX35XVur5hRGIAn3Iwigbn+jRO9AsYGWOK8UkVshfAcMzQnQT4/mCwpfqvb5Cr/WnkhDHKa6SMs
WRTvU4vNefPaVbYNKUUwJV6hxbHC5H5g0q+q2J8Esh475E3pKWZL/TmUQU0xWkKyahnb2qtB7Jcv
szrcvBFz3qSW8X6yikKLryCHjiuXH14zF5KDhwMTV6ViwRjCaqmrBCt2z0qw5d3h33TISzCeHod9
fsMfXyoCuRFS63myQGJICCswBJYi6JDtLHkpxHnbN5pUtrvA0aAa/mB58S5i8+WbgdvhdvUXgnTv
mykjZPnObwrnjACZ2gFgEtNQGrpqbXvrdv7JWf9OL2qlEidn62ZrAg/EuUaDlWIKuxQ0ZWbpfu2A
u3vCG64PavKQu4ceVGG+YfZ0aUGsSavKyiwocK2mEpq1Dvf965cNLKRifRTGuFaD+78kYloRg8Bw
z1Tp73YLXPTvADOHWpiU/3+gXewp7cWhgzel3mCM2kNzf3hiAyUnODyloInRA9wVyaSC4+EJ+sne
YbE831bG1V/ONFWeRJYW/PQttSOj3V4tKOmPKqzWbIgFILT7XB6PxWpqqLvIWw/6juSW5s4ljVyP
YYFEmCdIXKBKTklLACmFVA5/9YwNPipTh9o8TRj4oDCzHF5qKQutla6ShMUSJIcQrM94dt0qJkwk
8SOUaodgxnZlWReqId3K2E07OGr6gIdcR69hEaMLBB5M2kdt+oxx4+nAZO2EhbwSZ3ryQMA78GgO
OKBuG/246IeX5ezAzqp2F1r0G+xMkCrYOj8ZuGGUCF/70mnJgSLjcBkbISMj6ckRnLFm5EoNCm5x
LF3xddy6e6AIhuCwMN9AwHKeFHJsblpmKY6gtss8D9uvLTJvLoRtM7yYmYQdgVtEtdDpOlaIgz4g
khUjX3x0FwcTFEZ0rnfM2kqzVnNDZcX/eu/TmLB7O/T2gKjCQVBfmMdbsqXeE5s56C9i3mWx8MWn
1XUZzb0/btjWhKhdGoyRujeIf6Hit5aMXo0DnSbJ+4gNyJ7+vQ3IaIuf51uKmWzXm8lnQtbRoWtj
BTBbZeBIBoE/rYPaHC26vca+8WxnagbWhbqqsM9UsWOArsX694KnYCA0sJ+bWAWpXLUULbJWCm1c
UGuL1nDEiVfifecOWJt9vXkUyjFph3l4CT5Lo2z5/UP2oHJC2q+MYpG3X6SUu4+sZCom3ncY8xZ8
rsTjYrV5wNDTMvhsaYLadNCYKdVYzrmhh7aMkfNFh1UR//l5AzUUZlnE5yRwIugJtyPgKoHWn47o
hQO8JZPTie7oKJP2cC3Yao+4rBjbpM641n6pH+sIDnLfeJT59JTAbuG7TkGBttFh8iVt1qvegvDv
ZeqeVip2tJAS9FCbq6L8C4xLLGaa0rmbqN3r64fwxiVGyKLxUkfNHn7v58iOBLsyROnoDldlKemO
CO0gBadF3S2D8naXWxWHJFR5F2qjmPZxN2K4g5hzEBkR7VNMiQG5NRhx4xguLMEmCTUvVXvN8Rx8
IF95V0zxdW6/k9Rl41g9WWvg3XpT579tiVzlwKprNa2k20X1vUnL6v1pGvugxG0hze/8gzmuL53F
yJkO2hi+ZLlmyK96Hv1ML+ehBQACmqEjQ1dHCnPM+slIPS90aT5mDy1gNU0N7ppI2HROXU+elYuW
QNwweLd6+S95yYS4sk67X+GO3Euh1DMUxgFGabxY6ue730NUM+3Rr1gfXHiExaG0FQcidLwiJGj+
LAFQoAv7YmFRaHJnTRfX76vWQVyS6v3mJJHphqFYCBdJak/zoq+AwuJ3M4dSQ8Q6eBoGeAdX/lbO
22tvDtBILPDiAGwdkQmWfsXe5B8JVMbwCK2zkqjyXNFggutHPzMh3FhAG8goIdG6uS01p4jon3xH
4Yz1zAwxVI2vsvAQAM64PVgZ1u64PixQiINad9O0YzvJ9JE8f8mSibOY8Rl2p3G69RTnjNrgzQZL
ngHf73+sW17T0YAvnyVjlWiXr/6nv3U8xoD9ZGtg6aVf2mAQ3vO5qO8wI2R/zi8Sb00GU2bYwUEP
2ksXcgcxpBVhCETqURTOH/CFpE2hmBsqyc1l+YiKMrQQup6U3CxaW7+02B8d19riw/q4+jQGnyIW
BS/pcr18solmfGpw9jml4zzwX6Sqtsw+fu0P8kUmOVv73qqV9Nk6UuGjUVXtMZqAMFjJaoh+uLe9
bGzSAd1jl1OmyMlYPu8IBVdnQvXWNLs7Yw9lNMQHcNWOsR/7g97NmYPo/AhCX/J7W5fQp8nY9LrY
/P1raC6a8qD01+w7Sm15wibAPUJueTVbgikR/qfMYytz/umuj3Qo0hbbN1LpMesl+srnY9Fo6Gzf
i36RmVYjb/Pm9HIgCI7qfMwgqqOkOEww4aS1PLyZ3nJfkFmJV4nrxcyJb8+09uuyo+Jsft5J+3O9
z9q9CQ4Wam7d7p1PQPSx5LQDx1CPZz/p1KUYOr5w8ASAc3HkUbSrcC57XzltjvAWmyOD9fh1Z01x
DWoFG6noJ/90x7njwDkjuGsPo1hpIKKj7yy+vRb/vFW7/WHUjyP63Eq+8HwppC44mrzldrLLvKeM
bxdu0QKpcLXMY9+Jrk0qWes5ckqJLSHSWCwagIpU2aCRHGNUHow12dh88Uf/cF09LOacaOhzjWhk
KzyndElzDFMzd2F6OZywpoCroyM53mzoQ7u57HXsn+KJ2mP12ElMP+MuX6x1DuzGOQEJOVJSRUOD
Z9QXUNHNET6HwJlZ6j1sQ3RyRW8RXeFJb8Lpv0gNkAcuxpWo74/cWJXRS78yf84+Vqm0nZT6RIUB
FNnaTlwm+QdbhrgGNU9diUtmjHI7t8IUTiju/EipE4wyeAr3J34WacPT0QGbJHZrhu6dcrmGIwlO
1mp8BK6GUHQknP/ywPDAlQdanf2djvNEb6ovXhENgI4zGBzlMorVJRhWtzVQA6EeNx05lFjPJb1Y
zWzCaFKchf4nG7+b3yDEoF0ZnYN42mCoZtG46uBFCv3gfSJldtgAOSOuyKrZhFPK9zAh16V1cDT7
PLeW4+YcfXkBFhQcyydfDlInMmRo3L3DX7LJqnEC95EfbTn3xae2ZkHFU1mJyFL4QidAuVxIzreB
7Atehtb6sWgIOLBYJon19PGNUHZzVhk081IPlVOS5Qs2ogVpIZEv59EB12AKawV4F/Q9xm0GRb5S
8ZoMd3pJ2X612Dd5+/hnqLxUIP4a/J6Ty+t212+6PqfG5c1Lp5FEl51s8tBMKNlH9ltL2Z5EPCY0
bdz+Bxo2O5EpjRTQzU8gAHiMdr6NpWlwtzWaLG89fRxwggUqWiQsJIBIPvMeG5MDZLgTf+3WgKpG
mglMMpr33OfJ0nD0JaARVkVuK/ZZAqnlMmy37kaWwi8GUcenFRfBHTylDxIz22WVYgzofoFzybOj
YSpcmuyj08RPIYukgzJo+C+OHmrHy0/enjlVi0uIhjHM5ViJoGyyG9w9QjpGlmlAxUN7xMnmGfRk
PvJbzmCN6qiF9VlXoYTP1VUsOE3OovZvnK+ccisD1GnZppnQPplBgdDreMticZhvAS/4PkxaosTg
L5+3cnB/Ua35olbb0DRphPfYbEQt5mWkPTRemgQEWd1/GyHhu11VMMo65y+0lP2Hghe7m20cgs+V
Gbv4d8QlEMrREb5Y0ZQ4hML/Tg9NbchI3cmjv7RlBpobW91uOPewBQ/b+DFCfc+I1Gs0GYVKjI0T
07W7kjrKP8aAN4A6Ui83nVkLzUrL0UfvU8u9DeBRfxGATgCkDCJsA3lycK/tABvPvA7qNdMt9QSl
jft4iy7YEMgOY0YyCXPmkogh0toS11U8ZVc64bIaYEtwLpx49s971ioRfvqNa+/0XH4Q85WiIS00
TfeQWDhqnrHUIS0ilxnVa0ELMOGnan0+5C1D3Ptq11cNl73HuUSNopNTBhCAj7bgp2sq2r/r3jBq
dAtNN4v0KN1IM+ftdyTcwf4Bw/UxI2/374qS5r4crL1AC2Aoic7H0O2y+Sli7iNeTmlHEtc9hozn
vBaRTqsM8e8ilYPKuwb5yv19RNIaKYFujWpA1t2Dlq1pmdZUGLidjFTarZczNwtt+4psUFTTPIVl
QhO7z+GosnZzpYbQEyR96//WspIh5uzviQaQLHRNy0ozS0LEnlbkaOGJ6zj5IW9R8a3naPlnr0iE
Avc0HkyUsZNmL3QWRcIku7rVEB/V88XIruzjNrd9Qmddo1pyxMdQSk3hR0WkHgJ5UCjBEIzv6G0U
+ji+xVukoRp3TzNlB45eXhERHTvthBEqp99aTCmsxB4zutXj7eLAHOPP2pEoz1uQ6pwCYUsqayn5
DPaevlg4CJR1kBUz+c3LWLAgTbPc3CFhQo3IAO54cLponChJxTAsaISNsYXsrVoKc/k1bD4tiulX
YsjB718ETad5U3Ghk0TazFSXp64RmGLiNn39GwRvt1yUj0dOgEztlWeE3Kd9J4pzfZxeN+wLcgUZ
s1q9LSO6fWwJ94z5v1VRFiLC+mwljgUEF83Wiu9EHrVED6CUFIIPodD0a15WY/JduU34iO7RbtfQ
fvuDeZGmyXnlIfg3wfH50GGk6oZFuEmrjzmNLfPm/51054glXEAILsGRnBWq0RGr3n7EZlI6fxSP
6s+MiIP1L3SStNp23JLJm2+wDSB1d6rzZbP84GSolQvZz/ufc3+cT31l+pnYIPC0s/tmpHGjbFNi
TwJzJNLSekQOsKliSGskCV6VO8XT/coZZJgb/Me8aNzUC19Wx3kpLRzoAeQCS5+4PKynsBjjd91+
2GRZ+nLvvufyC25nHiutKvZJYCFs6O7hoYbxmL/fJRlL3Kk5RpoUQ7465g3XfZL6UkGwkpr61sv0
fjs34FQWmKq066S66tdYUZNYlWQqFpFKcegYyFWObk7ZwscxY13w3JL2iFUWnu5Fqz/yMFTry1vS
WWkhJKK/7TeUNEjo1aIW0iZSy5PxPLT3ZV2EEWVOB1JjjlMbNjR0YCDJt8JWrcEwVnbiKYWex4zh
p/6sZx7j7+x16JjfYwye1S40LINCFSd5l4xCjcTWOZ/ymqcBXO3ZA+F/k9LlTxr4Q6XeB6QRkzec
bc39LwciDOPCNiqaY/A2KpuQzQuUiAepOthICn67a5FZbQ6deASZ3nuUgRYFUCrj4h3vsuFkvHnb
1CMI2QcObxqRnpm/17eJrkAodV/M76VOh+K/oSrqyIi85taaDBupckTW1NUssESX4KTLiEHPsjkv
VSl4iPfCxCCGfBWQgcS2C5C/V0bfI/612cB3Evc9x7HF06+sB9ONiIYJn9EfR0yuPvlYfT+OBG1f
UW/DzCv+EOBe8FQ1xTAwBkEqCGqclStAU+EW3O/8O3kfrRnZYmFao4/vvJCqn2ymVCBNnzZuYhR2
9A6YKUzbZoyNfRYWpEel7jB638p623dK4ZFmID+xOLmv/1/jxSP8cZ1H5niSW6Pryc+q36GaVA6q
FfLAQTMCcu5h5QfDI4KS4JgbMo5oTjL0FfZAKPNUiw2JQhN91vI2KdSIJ369SbY1DIMkXf9f9Blo
9L2cohiBNUzGI3X6XDHPuijiCeE0rtLEOvS5+W0hGjokjARLl94KK1JGD1oqseMA3rzLcsjh1R1e
Fxz85QLlgJlvvUL35Y+BsIiMsViEAFX1Kj/dvYZ+7QOyyeS/USO4+CfrYjVsvfM14GCWz6V2FRD7
HduPXtPo4n7cACowUwhSMrUAVdAdn+45iWi4FfyPegF89tRm/XjPSV6GPdSpqstXla83PyT7g96X
AH6KkWX2d0HAx5O3w+V+E1lSaGNTxrUtf/RyvOXIBxjSoO04url2l8Oa+zcOuNgsL6W6rxYXXMkE
S0ePrYsDSbeIXq8uMbM4b/l2GWI9p8/kMwDk4VlVojHWSHvUc7VT6EzzN3aw1fejiKUqCZjKXgJD
EaPtpA0+QWdBTSYLhf+6Ysf9voYi6QeEOvNU8vKOXcgd+2UnMJtR9tVVxssnH34l/dD4GKF/01P3
e+bW0HodFhCLHw84DFOgtDWd5rdkPvVXhADOi9wvijHZxioUefjVh1bWlUZe0RQZRx66c/g/tdnp
uLc3SyBVJOSBnMUOZdwrCu4lr+330bdyXknWX5QbLdPlHl5r9ufIbeT9GhFDM5mTP60jOmtFClm8
rddgbqKA4dtarFHEzFWEkY8RHHz6cirRc0IlAtBiwRCbVyz2n5b//1K2g3/BGEgdZawu2FrXr5vD
/piO3fC6e/UYvsMDAfusttxjTO3nH2ZWRbTexvq0K9ugVHXB3D3mRIFYQ9e2CG7AIkTmoog2sBRP
04+voNoE4Ji58+1RBNlSH+zElT52sjnAcVErnM+3XhLmvhgzeOUEbA9qle4ueknAo6oD2F/R8dnQ
YfEBCXMS0L9Aq55Vr2eqPhtSTCUcgVCvcumjj9Vk0HmRf0wF1vk0vsZgaLxAVfeDd4Z+pQbmKM/h
ytUcFF8rexQopNrbalWsn7EeNjo02gUm/dTO6Sow1LxQbXhJWgyhKaQywtgMTIZ7veEWd+luminT
Y+YCzlzokWKYIuI9j6kZzYX4S2DCoAFCorgx/LFHiN5GdIg4jIa60zi+U0g8zs4qRmBCiRFumMre
zdbxmRnjtX/1ghdi7xmAGq5NKsGvG+0A1KhxGTQb3hn6z0IygcVxHvc6q8hK5UGFM40DJdXO5WAV
ZPw2BsfgiLHS24bxYvJ4sjKuytwuitS/0sqt9sfLyfyxKeWFBw/gV2WlLWvSEHhOc7Bi2i8Lll5Z
qxSJpjgeYGFcCNjc3sg9CBNcKH/xPnAkR4wZJRRvu5QGSfaJmfy/0kHSwdK1OC1Sr/DZxzqMO7dG
UxXZoSCS4oFjLs6oAG4r+w1rgc59rzIAWOBwJSsyCC0qFjncbWiKT2wqmv9kVcRBnEF14tSPcpqr
O9V1KqcSxPrGKrAaXywHn6y3ppG+igbPvqB58uA6kRAPxSgR4M1VdDXXAl0sxTRARvC1mbQd3YtW
BgpvS9pRRDCVVQ2LdiPILvJDhT1nDwJNbTlAP4VkUYo97WI0Fo2Cx7KYa1u0XaD3f+QZjVJnDsDB
rzQKDmfPnV3SSWum3nrGHZAG2NW0hb32fckK+V+VZSLqlmE7EIgK1ESxpRl24yhthv7gGpdnBmyk
99CNi80ea1LYn86QsP5tg/vD8bczB/SL8pEiWFZ/b7jTVxHnfjRrOTB8yuj0Y6C8qULr9um6Ik8A
Lcz1vhycO4hhXeSvSfk9YjBsFmEc7HHkirEDVcj9DxIEIxyM4Ep7ILAm2qANgDoLmtEG4DBoR4p/
KZIFNad9wDaz28+RJv5a5hu9ok+/iPsKT+K4AMLRMDh2praBfa/uAvbhvmk6OJDyTYBYolylnegZ
MGcKYRG6rwxpzyuo5hkPi+cjhSzvZEC3DxRhZACytQR+NZHd50KVR4ecSP7cO6EtDyiqo8ED5fIu
1aP5NRqOxrCmxCC8Wh3zaO+8VCBmAlZW01nS39tQ+9soWSU4G1vtlAl/5VOCKX0e+8qg0/VjQufO
BRUHxvwatX8pr8BsBSAdfZpKqBNwJlpYxhtROe13eyt+DwJidm3Wcmxe3pIPhF+7TXGTylr9YoJy
H+Ov8XPPkQwL2baRTdSd8QOn9+C7gIOeZE6TcU4IYA6oKoGJVTXSKiWXtu5PyypjE6ic06n3BfW7
86YYbNSVLR5gIxXZ4+Jl0Px69lp9iZDG4Va1f2G3LK/8+98uwGnItHHXJhx8uoGqW88AzDtyI7Z+
CWuiugFYwk+Lpwzh5GQdj1TqVxY7Nmtp5RbqCIAVmQy0Q3nNC66KtG12SkPvV8gQ1NaBIZp2Yk5K
2jFtphG1QTutyDkovzmWXdAyy7it1+ZDAvztwl0MYaE/8CEKfXwGxgxMRE1E0JEQa7ER9lHSA4LD
lSftIlseKbdAkhiNmqCzTxs9fF9C0M5J+UrscMKHFCmvsOk43GJHA8vGez8AIE8HcSjeXuiGQfuf
WBp1U5zCln/e2VdXJc4s05BR3oxRbsKCjlAvOcex6hg3LjpA+IrWPkMp6VGOtmiHtwTlJPpmCG9b
ffN6vq7iN1UPcXHXrPIt8GfJLrxKN9K1UsBTDzDC3hMqT/1rKUVqfweOuJ5UUL3Hc3popiCjB6n/
737PPOroiAHwuS2Qkv4xd4ITRtLzvg3Z3iNgMNFG81RKf6Q6A+AWrXemHj1krFpzSu6BN100W2FM
JLrZOz+QeFaHhlErgZl1IPacbFHzcstWCuTjv1KMkHTvzOcmQcFgojiXA0zeT5C+k1vw3f564BLH
HQ3pzRK2v8yQ1o9c84UPpvAQCz5mVlF1iccYpu/qY4RWG0+jpwAcjLMXIfDUiD4r3inHnHEMznSN
qjwP3bX99xHHPGLIYVfIcg4txt3Qs+WfYTSUFbytnfqCOR1EU0Rt1uzMr+3/y8IVaCps6dEeLjev
fuNvc0DN/8eOFFwxxjq9nID3z/fNkssIX54jGeeJkFQBLo0mYU4xulMpO/UnslhLMZfJ0qFFXDCp
ei9HqQdxaT0E4gdFmkmRJMRKGXQHjwr+aTFI1IMImcyf2s1bTRx1Xdld75TmkwqKRHAyCR2rQluT
4bOem1kE/5k8Ye9hHGIjbe4LeAadWqFo1ArTOjUtEj2QLvjRsnfZpHE1TxwYfINpkEik85vU+eis
uUxzQi8CmMwP7ZBiOrGzX/jeD8cTdtUv4lv/Nj8r9mbw/wW2lL0SrVkwjo1Mm5Ediyr5yzrzpKN1
O4Gtyb2PusxEuY3RlXjqdGvoR3nbQ3GQz95RiF9CmvRyWtslS2JXFiXPm4HTDV6UxNeLemhZdtAW
cleE1M13ZSuhfeNE80jDuN2diHSO7n97P4t5m4ZgoSf0b2zUz6wMZO9FIxM8rZwLCI52ZUNbx2s9
/C36sLLDdrHz2ARbVHJwxUms0HcLuSafIDlxYtZQiKwXeaWKS1EfYHi0A53XKH8xJFGATqQ8h681
ZlMlU2ndAAdLyRlZUBgn+3c4J4ZrGVDnAmMdoEEi9vLHACALmWjyJaBG+pimU0fXes31ANOl4TB+
zABaB9tMCHIlczCCMJC/ZFIlzI6N/Ub6ASgxyADmMF0kvLgal8oj2tEB0rmJsfiXP/4AZfvvXqk6
VdvrDOWhWE7OVNlnZd/RbnawBGUJNHfkJg1BWGzuKD6AYxzyAGTj/eOkxJDZEYPkynct7GpTbm8j
ylUPLZSv9yXlgzz5lht/WKLNyFQd6nRZuXUcA3/+aJKEbJ/7cxGdy1N2ZygpcbDPmtIIsqOd9Qaq
LibgyFUtItIZ/26BaurZMNfhtfjBjcNQVcKG+VOwcBMpjonZkov+TpUB/iUgz+kuVJlwVmJdFCJ/
e5TA5TFdmPk/g/dug9e1b7JsFNzXqwAh/OVY+u8BSxuHVyW0iZ84TD9wPRxOjkawrt+U+foJm51o
6pwrVHuot5HS3fyL1CZhOXvQOFyubRb3UzNtIo04KJotHEpEu82P47i+pyUA/R2lDF4ozXoCvlvI
Pphgwc0j0MVOsvBMZEyJQzQjdVS8xfAZL6QOqP9bmju/pToFv6tXZAmeR8qwO+zj/kn+1qJMhBTq
ExanFIn9dv22ZNbkyyJdVlUPM1deoO8E8w2k1lHfWLSWK0ZXoRXHGVziplLDGa7d9jleQgjvn9k1
z1Z0Z1496J+qmq4jvA1ySjkbVpUunYX19yBblvugaFnJbfOOyhU8vtOc+dtKEk8JxDC0tOhnCIUW
GunGuSIdF690CelFDjNZnBTw4VpEe22iBUbd4VF7sPKwGujKzN6dW0qpTmnIOOS5cL1MJfxQHf/8
AOYgNvnnPsIZInAl+WzxKiy+R0r1P2eKaEmGa8eiEDRjFSKjxkr2ANv0va+k+GqVpl8o6/wTyU1X
BqVqtpVKPT0Azbz50JXKsy8qtPVUiscT8qmbuWclq0sfbWLNDHm/kwW7vSyHhM500SFyRYs/Xjk0
/B3vM+MSp95uBqqac34591pYAgDt6I06t67vf5II1hF1VUPv3ABjYhtd0uoAq7xVL6BUAv2QeFnO
IVoJUoeSNFus2yM04jeQAHyvCoIvPAKzVYEl3IkCLCYMUMnJEFOWMwo7VcqIJi/RIz0nnrDF77aC
bMavCxNRcnOfvhQT70KnvS6xJXaz3km4gVSVMxpz42SNp2PLinnkLN09wZT4RZXlMkuk7Fgw1r+F
eNt02KzRf07J1YHPctJR8lluXJcOd/gyjDbBNIBfyO6VhSaTMee/nwbBHEwOcFIltLtWc5/hzQWH
zA0LlXXL/Tb5Y8OtbUBDLpTrXVSb9nXcgAbRvsisIC5aSrJQsKRQlwVHbMJ2DFsvpAjDz6FQOmU+
mkYlkvO997uAh37Dq1iwOHJF8I3HAfaO30DUjrWEcDaZbE37ExcR1Ifptn8DFsRldD91iuoOUASi
y7LCijZhLZzrX+mGktvKtgAqbjWNzlDqJIVkQ4Dv/Wwe1OMHGN0I7aqMAyceBbeb4NgEl8lcZNly
11sTDngALxBVNEiB0+O2EeS3DH8euits0oeWEF4UVHqf+qb0f+psLcZkBmwEZSroPDQvIwAESoyh
OQCXnVaSgkceO/M5eXL0QyHkHckrmoJ1OxPXUum37kQEHaHReIsUX49mBguhQGc+akc0Xzmj34VV
adDsk6S5hc3j1IcKOA6GJwtPQwukdhWxrlOlxqcynROZr3+rV93Iw6JoA2Zo15YI1CFy4Up8idQc
yMFjnyCoB6CMRSsFT1Nen6HdpUx/J3FEDbKud/KcVgMApFiKVIKtVHhEcLV/cIXsJ4ghl6Hh53d0
9GjyDxwoUk0hT/6YNQbLcP+yid6QslQNRxRwBTFkWez+9aVmUiJ0YmqHE3M5HDp8VLc9gEg1znIz
F+9GcyXZ97sAQ3V77rIsgVev8hIc65wIbIO1hQ2kavfwYkxu9r+fERI1bVZVzuPI8uFHVOBo//E7
4f/NMK7EwZRjuyecFGBNmTOyDPBKpf4VsMbux7IcnuDJnYESahCZ1poHj2E0aapZhz1MTYutoj5p
MitgAzX9dJe9PwlowyG7xzUvLRSNp8QcezpQL4jtBzB42ePM6tFolCfPvNaeoMh3z56AeVurWxZP
SMWKHzztW8kHGq0dHYFh5ZCmwAZpWKYGi4oRUOSn5HapLnghDyG37ow7poy6XENTA73vzzibDQv2
Z2Q3Eh6fpoNQ8GyULXEpNb0Xpbqt0JkEDEUWQSjKllj6nd/FUfvSzyS0/NciTvmRqapOrD7VVXp2
ygmunXrg/KBPXstJ3MkhYxyg11Qcm7axYRNIuIk5grQ8ZRJgpbbB7ZVi0jUhSiUAeo+sFx+3s+6v
E+ScSmJrJt2cvS3bGOeT0ICtqOxA9mGonpmgo1wWXilB2rGl4VNQF7vBASq8IGdSGSXIKleP/zab
2T/zxjVFoQJReLhj/UFWHy6uXxToKtlPmkIeKNbjLbj6tQlNz4WH1vJBeu54ZHuAlP0DmCnGdhjf
b9u36icWVASXpVHxtuDHFFwcCfl6gg/OAl8anzaVLfHJBhSTNBW66dOvTNmlWPTmPxBCM5GxGd2E
9HUNqbDkFtXUY/cs7Hv4xE9v9d4ZC2ydvcsp8IIv4yZDCjAE7QfP7IYBBWzO5dc6ebIBOaMKTo/E
nLomQE2kj1arEnn3u8x9VNgU9dM4i4wD00xqt0fmffR7tlA5q4fBb5AVvX93O54MQgYKKBsSYCj3
J6ioYTRWlOdL7T3Qi8Kj1KXQVX8uRMHs0Ls/espXuWh6YIunEmD+OHkNvED/9os0Y1ANkfHsxMSQ
pVQp14RWEak4d2h+YPbtolV0z5y4p2bejgVoYzL++QKygRS8lzC+cztp6MOgshtXKK4J8wATtzjm
dxkKnjizs81h22Rxy+T3UqIMZDS7d/gdb31dNyEIhQn7j3P8ALsU7yYgKpM8Q0WZu97iFiSDxKSj
UGJCO/RGFLakSTa2uJQP00spPlcsRgj36++2STthZ2HD3j+xVDegKX8Ifd0usQxrWcX9kg7lYytu
eTrTHhzdaljQuG1XFaJNK8vBK5B1nf1jbJ5YDz6HZ8ODbJZIXMmPoJGTqmt/jOtxk6sqRQuOTbRg
VExd61QHRlV6nuBrWUprR26eTmfIM8qU1JyW//UFVa5YoNCPKcYGrIY3OAbWVhYogWfVa5spzeFF
IAmx7rn47xDz0pD4OFMkLa5TEpmubX29qZ6yOkl9GANV0vkPUOy2I/hvde+MM0eta/sQUs1vDc9B
9OF3INmN+/btgaLAfqPG0T/srLm7DmTWfWN52DdHJOvTMofdLupvrnxlLf6JiOk73QSEaVb7x3z6
efKSqYeQnadV5b0TcSlHjQ1RufOdwbeAcouMLsFXVcXR2r9960XVVLB6Ab+hwr5wtferTHdCiF8I
OtUQ90mmziYdKfgWsMdmVq/S2JJAd0hzgPNZwN9p2N4EFNPvigLQhw3QPcQg2WUyyZTJ1sQ2Ja2q
OB3yrmRjBwpsrItpYE3kU5QYudJGFOUisqVeiqKk/GBwgh2zQOUXBD6ZBroeQrmrZTB3qX4Tym7I
rfUoWHup/17y6DCPyPHmfoBKzvpNUmcf1Pz2y2A8hmd8MLT/OAkKs/DIzFK2dqudTA2RqxP5j8XU
10723ZH1tp0JI60i/xEwJ+cTToOEsV2VYNscnL+RCNV3ybWZ5/nBJqRW6PugCkr2XxfDUTgBK5Gl
bxHnHkkvRkNFeIMOmo9+kXB9mA0Y4r4QXc8uSF0WoF5Hrp2pVdkfg6rY7SzlCAiudjBJfvH9z2xV
tyv9d46X22OSBH13lXC9ieOwa8gIwRUCpCtNpC80fIhbZyajLAJMW6hxjjjOGoQZi6CAffhZsxlD
kborJMEHtpUORdP5znI7VQVu16dHtvmdHBIHpm9Jb//NiEe/fT3VTH1kjUv8JBrzUSFrkSuNyvGq
7t7dM+D9N+RGO/IQtZYCqzKTzqf1jeBFwN4mi01i27qIdzSIPcVNyvGbxESB26Hlb6epnBDXPiEY
Xx1HWjbO+TGQX+Qy9HRQGeYoUsszwNgd59haCXjhRU4wdXUV+rcwNhBOSZn8id7IDleGMjuTl2Fc
472XoMN1juzsHGS5Sqw8+4DsZKCvlWM29/PdOumqTLoDJFg+sVp3CChp1yT0sa2W3NDGZz42+PBp
xVfYnbmCqIoxso4noAWqYjx2a8Ej/poMzy4cfUcHu+gkge0cBc7Y+d4tE9PD6gZ7CwUg7O/zv/SN
Hyp8A8BCgHaGo7I4+dsl84sVqZYv2dvO4t1b7scyHTHEol2t20T2ALH5UUfe1o6o2RmBCfSKjPE2
jj3G5z/nbKUjS95MBQdT7Th9sgOEMu8vlw7z/h20VfcjUl31IWffg3fCAUKAf5bTgUeKBmpwbcep
+KOkt6b/WI6M0i0uHK229thIXxYmidEkNz5J3qJCz8d/YZDVZBMxcabiIg89RrjrdKU5mX19U3wU
/J/xgnmdMe217ga++qXFRMTVTeQFrguzeDOwT/izhs+i7E8bj8Vv45KIF/p1krENL0U2vKyDNxx0
6oKTU255HESYoWvP/F7hP0iyqxPj9qv4wxeiX0Jli+se93k/Sa3gkhlEy0gmAnZAoTHPZGjXMPWv
1EXk7qFqoQlIe+aPW6UdOYoXaog0YP+N5Ym5XPusylRpAaKXovEGWtsEkwD4kHjWFQkFpQd6Ec/n
vaowXLGyIs2Km1uIMEP8bNnttFdtGja15ERFP3auzvERLGAnSe20S16tXyRtdPPbKGkGV5AeIRYK
lXLmSpwMHk0yn3SzsAVFEKRuorwlyerDEFgbQij+G1DvEcgKzohrKfhosaKebTCTXk46CfOQ8JGb
MGNONT6xc+Vi+bAOINGw3CmjgN2gE35MAR+Bosj0Dc+xFNKaf8j08fKTyfgsWcgqWhOjnnigCcr+
g6VMZwz+jDGsKpVSIircFh4O5UI0lrbADNQZZtuC/M5C19kWYkk0m8PMLvHyG32zal4XEWD1X2+n
4IAQl1ceX/HTIPO+8r3+NyC4uDY/VPRb0ya4dNmzS0uykFGRdmPAPyaAX8FT+viLKmKC+datbRyC
AmbS8NwInXL2Pe1vxFPoV1wX/MGwDjq1GSPz491xf4YmypkTQkJnNdPvyy1t4vnFalfOxDOURW3b
TKMMKifhLF5ZW0TMHD63Z7kTc/K6BNx1VL+tMbS9j0a7MIws2oc+OAUHgeYOV02/F+68EaC2XYH7
G7qUIvzDS4GpX+bwQeqfwmpNcPydSUXHRHz+SPeqX3LPT9qLE+MQpc3xod108lPtZsaRssYOlgsX
fa4dOfRVnc0rGLM/JAV/DXLXA5bsLGMeL4IACu9keR87ODnj1gyFKKHqNewK9tCot8D3vvQjW+hW
KFAm7Ch6t9gAwdi572wVqDIIyb+5gtb5QGFrjYe+hV0frzys77qIhWbd9aeYePY1FBaZyOnxh5UX
36lHVohsVstC/UuNb4aanUWtBfgW8x6fVS0OWNclymiGV4BZgTQ47YZXY3tyqBhNPvYCNbuqtVYa
lu50spKfTtQFQwWihANBIHoXjDX/Q4rDnl1/0vG64oFiOMAKExqa11aNjVotPx0TIG1tFFUXx2do
llYfGSN75384AcwS1+/rxk7DK2pro1CX7LROnGMaquh3q0Zw+3fmY85VwAp9EonDnHg6NUKX4nIg
N8EwGCjOtE9ht3tvrdqB2wzfTbB6WWBnV96o11hHz/X6QcGAsSEgvgxKDZPvmMaKE73FYFZNhsM/
raSIrlDeOjIKiFKfMviUXkMLvlNzdkeKweubDeAQiu/MwaVd6Dme2KfUycmUYRTr7ucV1CnkyRoV
IVxGAzQt/DbFRpNzkbMdezHizkEaNJVopv3MUWU+AZzY6Q2oBy2UV8wm08PWcN4F/dr2MRcMxybq
h1w+pnBo2/0iYfBUxpKmoLeBrIabitbdqLf+gZTN9MgWKvp2hNxF1b1QW8M7YQcrPqSVF108TdjW
MUHAFTcf2vTh6oMGGUpWERHVsa8aAE34gbD7QvgQWQKXG+OCMYBrVms4SLMy9vYXulFUrQA3jG4l
uQ6Ut/8Pvw+NFbCxEax1ylz4gcR+PD+CcN8vPP7X/xH805F+fTlbXTwXYj4oCXAx18gX19Q+SaRN
0vK69L9iYm6ZzL+8emcaoaYK3fH3ec0jL6j0HMuOf5tXIUA5kt4V0F7OptmAgdSjztzNE5yXFwmN
NsSzfPZcNQJLvbfD8/T+J9wVosFpaanTIt+lFgZoForMqTKoU5u9AUlVhhfiGG9Tq2Own6VRhcvc
XEez9AyEsI36brHYUBOaVnKpMoqx0DTBCufBurPVw08ShYnaZhz61W2wVg1L16u0a2UPv2hwY1ZY
gIhH8UZnJMev5b/+x9XJlxSFWHPebPIujyOTK7/Vcbg/P2sNnf12tnIg/dOn0CBDAKEhNouM7Tw5
sGgpGUgLE2rDYDDLKZGTsNaQtoJO6Ztt/NXQLtfKcgEU4npMat5mpjZeH2A5x+3m1+PU3nb/lcuG
Ky7HXcLGifd0qAtHT/QNaDexOx/mXRd1vykYTSMeZwgAHMeF1IICg0Au3/7yBhI8k7nfn6UAaakg
C9OaH4nc9BQRIjIhOQSKR9SieVwi/9w/3hpFdNjDElplVNLcRcxFmVj+7ULN/tmDAiGMjgbX0pt4
z6tOqnclAIAT+ZGIWxwtwqOCmXHZDD/CgnMRg6HbSNF94PLPFy1N9vunvZJcMfqV5H1w4nMp/OCa
aUyyFWA2ZnR9Zc7oCcZsVMOk4U64g0Oky0iN6OCvRBdiM5EaoCT0+2M6SqdnCiz0023IJtmVBTgp
HXMdZ+UYOvuJmWZ7XqsK8LhXCZynjN6ogZdfdN+upybikYwnBWWxms6qlfhi7nErZkxixtuu36YI
e2yRBe0tS+tYnmLcEqSWVwLmyOI1fqSDbp8O5dQ/4TzIoj3BcmGWat443IfDodPipALlsS9nBkvv
adr/h1g2dnCpuU3mxGoxpKB0tMgXiW1tvKBYiI0BY8zyfi1LYb86jZxyV68QAY22JVf/RFngN8Cx
QK4ZYR4u8AjhdeCdKU76KRVW3j9fWVY7P9ONO8WrtqJDqgFe/8L2sqfY2Blejd5Uo859QYWrvc8U
6i3mYPxvxl6f5pqZtMH9GK1naViq7AuYdwtmjfPwaNvCPvq2hL4FwjGVoukVIKhD0GxU/Gpahdtp
FvpdgpSPLNDAHqw9kwxWK6t9OZSIVWtotFcUEnSg0lVoWx8qdHGZ6eC4su6eiZrI1ySxU17Ieduw
ePtBHbexO93j4z+hQHt4KFtuRtKMGWJkx/K60OawN/Wpp49XLTcg16eRh5zxtCY1mHIheluFGWiK
xAaSDdZKf1Z6NGj25afrGhXGb7BG0sard0tUa12K7ml2o5Tb+5pE3x9bYxCBQ2f+QZeaAFryzzmy
N3BXGMCqkbEDaYfG+yVwUCcm06AYI7nFrAfJ4VhGWX3Xoz9QhcJ2M1sI7dVtVu/zBGyKXBpXdvXB
Gbt26/kXydLl//QYB5k57Nw0CUrtt35QfOWIr1gA8ahLWkG+znuMNTs8VdGfiejvBEJ9C6y/4e0q
vsXbSlMVyefXOlmDqvy02Gx987xcHJ+fsQn67rTxVC5ldObnoCmG41D5xaTmGGAhBeTaNbx9m2dn
OBQ5KdW62yRtzldD9Gxov7ULDe+SJrerqjWCG1jYco1RNbq09vecnSDKErmsslRMvEslsWpCGcoF
Q8vJKXHwHjFIs3/eF9Uea/QIW1nx2GtgAjNUjtrVijiRrPZxcRMhiTrs+aC0P/FKbIONg7gPi+XV
qQF1Zm9rDMF1Er1BJ8bzeBM9OI/hctY+3Up94RekfbGqm6kX2i8AUHNQssUe0u4N6YN3CDST+YyW
ZJnoj6oE6Ng8ej1HkKB/1ZFFars4DfS/pWZ7iQPDjB5/TJCW8xnoQ4cXAI3TtCmUXeXWqayi++du
VFZ4oSrCep/AZV6X4csLJ50HoWOPCrxGylRcYKgIUh/CtOQ9u73OOqvb5HkK0yOqGl3fzGXh+lSo
Dk7dtsjgas9uzlyELS9ZzvaB2MDzWUCwouul0ZgJv8CR8r76kjEGzm/b12AMOIG9c6Hx8LojWwgz
1mQ70LIEla2qhBgsLurIgaw4urkyhMoNOXxnssdphCJ6JV403YLjNVlineD9pzvI/vkWOB29f/mQ
GCgG83V/ackXmHIT2v3/Iy9hMtkz0GX4VHGi4BVXYLz54dBLjoSI/bMfjtqYzdCeVCda/WuA1Zq4
bNr/I8wMcsBOv1HeLUDYMxPTw6S8G4qPVsUQVSCS5eYnk3pYHZN4+k5cOl+PaiPg3jQ2tEr15yLD
er/v29nE3HEGToEyymVSzSJxmJGdgoziu3YW1lZ3Mfc5mI7eu0+LZNIk1Lq+GfdtISvNUaz6bDto
A44hVreeDd9sYIlbzRni5Gq8nDUethzFvAFA2g7i7NAyznsU0hsDclhqZIYJCmSoyMUam5xsd+ms
dWUGEDRt2cGOndMVuOJSVLEeSeRfjOGWeeKLTGt4YwWaCDZyVDZd92Fg0Y+IyajJBCr+BekXAZOy
uB9mhvWy0Xs8/oG8JNTASSJBOHH/GjKnGxe7jsfNJw2B0TXHps9zULGXh5NngxZ5r1GiAGtk9eUd
oaME2ixSBQVvgyrJWFI6UMOIFUO4ufF8Aiu6FuANSO51rRH2ISiw4ITpW3AISIAYL1Ocljhk/afr
QNCoi75EdZIJ7ck5kyQclSlQV7Xnnd8TpUXhFZ2qwUDSE6DJ8Xg1d5GFPgYYcMKzrWckCdWUGlxf
6Zea2JJ7kzpEAcKUCn8reT5EJVj6cXJxxIpA0dLO7BPFE42L+T4YGtohUWm0PPheGJcESqQhCg6e
81JX+/ZzTkMROtUKaaa9taROE6foxupHVMXzbcElZ2Zf/9s+20eUq4N617tigp1AVoWDdeKLX2ax
+f8bs/T+bfIhCI3E3yD/r6a4NXjTVzw/RDpXquwlQfxAKWKJRnLOHz2zuDEtmBdcuuqZtloUgniM
V6xLmGerv/HrKnK3yaKuakNo5x4QV6R7XwHl7hc0P2yFllbgtaiYQ1kRbISiLp9Wtk2m3uc98ZX0
d7SIE/UH0W2tM3Z0Thogk3ImuwYaxkSRzb8DswBlx4IN+PR/PrEnDVkiqjaLsiyiid37OQbIOwqS
PKIBf1w3anC/FabRvqjt9qZ3ukedNwc7lueQBIu02FWIYBuStw2Bxgu7oYEKOeBu9SDSR3dnrqH6
YDoYS33SIY2DzMk32Qm5ihSVlljzWAwiFGNIm4DfRh/JM12byWWNE640Hm8mMSTp4wFQn/+mWklT
hxcat4+vNyss8tJZoupNxa4vinXwUPsXj/eSuXaKITVJGQn//blOMKpYTIBHT8QuyhPh/134oZDk
Rxp9swkQPflkbEnC2OWCLSLK71h7VLrMbQ3+kcUPpEZGDjA33VjpX4ngHDOzz+PMCGVngzumWO3I
1oEUxIymWGmWNlfEoZsjGrI47tsjfN8Y2IXVfgEqYlQyi6elsOObqGavxEEB+5UXsAOoDIskwoUA
v8b9T1ZzzFbMNq9YLyfw7YzPvsbfE5lxWU4DlXLklBH1RqaT4YzYvSGJwhmYZsG67qhnBUT3l8J+
6fyVdkPlD20uGCJHA+AnH7kYr7qhBosKk3IU5ZdTyf3wCkWXFRzdDLOrDuxRZdPNZu/TgsPcFXBx
IGiUxPsISidsuWtL7C0e8MMlBnRF2C4Jt7A/ONqzG6GeB56/E4xZ+lwZQ9wAB+tH68FqH0vdn2FD
J4GNYnYdj+Y5gI6uV85cQuea6VbpkzlK8i+fm4P7KRRwooVs3IE+tmnecAVE5/bBQKfonmsYjELX
jchF42Vecrwmili/V9dfoWh8GJmz2k/ktJRFWe89or/Y/LwXRFsNJe23DFO295FoeWPxjXZW+TTY
WlAPDtQH6exXe5xvv0xg7s7oNIMG/7p5E3Nr+2XYlhXRWrIzCxQUZ9cqR2EyERaCDnQs9wbSJb1m
b7Gq+8SlAX826lHkwVZTn9o91ZCMxlAyqKJEhcwOSbaOHUUp+aI90vbI4fMh9d6tt6xDJ6dbo/Hb
aPydQFxwpl8k3K1rKVgwtqYF113GBzAcJ3fPz7Bqw/oP02vPp1iIjpvsObruoFLPTHdaGMyzpowB
rF3xRgGWyKd44Os0jN/QW+9fOpC985z4lLLYnRwd+87Otz+qFuFk0OZHdKf4ACgR1869v9Iqf+0A
xeqZcIh1W/XXv6LYmf+MYfPUu9IKIAPQ/FunmLxMp462eFsHfUkVh5OiEtXCeAaKyyIH49pPtxdb
a296K3ZIG63fcD6vvyU8UtfHg+624X1bj4Mqtdf5pkIo8Y9vC0A8qfa22fwrrPYwPTN+qxwmTzc6
vF10NqZQkH7CW982Ndu7lyObWBdb8aiBW2MrKfquCbuvQt0M2UGQw97DScDZz1eIhuWk0stSUigS
HiwvEHDaKnz4eFje5Z+cvGYcg3y2OTT9M4IlGgJhn/Zw5K/M3QeFIimuRKY3qrBaa3Irz38pfDGg
W79CTXDkEZXGJBdnd8V4RqEGDREnHXzPy+dnFwlwVqfjMDuhlA+iYYgUb1Zrr4WzpcDA0oj/IuR6
TQe38934XGB1XQx3pIL3vDpEjg2Q6mfMKFLOTQ0N39gwaV+idu3XW0gCGwDUFrZgqAxNBfs2SJPm
68hmyyPYP4ItPK5W1ctVdO1skHEseNMhwgKOEkrB7veYSBs7sbJArHDMmNXV1hozR8Gxhtwo4ulg
tVjACqIXZYFoh3pPvn2lMD3hrsBNqgKbL7ZetTbksKcL0eYtX1IibLPNnxMeO9RmtGEXDUUxlDv7
P0kdqIDkaOsQgfGrAa96rnL0dLJHbiWtxMzGGdn+q0QBQqAgr/VJX4MY9Ef1SC5Diw+rnLyfibQz
41PTjZrt6GpouiLeXzA04mBq2b4/RrJ/yHk3te4zI+3iUPOHm2O2iiZBPWwRMC1md5nIuXFyWyvN
oURt8ZIy670FTT5qbmI10QCSdMpVMpPfKH66lLenmGFAzO2OlVbTMa2SanuOjmxr4E9KvlUdD9k/
DZ9Ud0ZWeu6/9hgLk8U/haKsrHfd8E0vSbgcOX5ARULGKHZd2lbyQXUeMaTOtX2fCCFur7L6KgRa
0iUNgODTuea3KQJyMj64NGtQ0VMVG3tv4S9DrjzV4W7g+iPWg4BthcDYaQ/HpK5W5lwiK87bdmkm
E0EE5kNcraulMFjkiIh5B66y/RJXCsHYJg5Y0gzY8YTkQGM/J0SkT1AEsyNj6BaF/K3bzKxhOlTX
UXf7Go8tXfUWM+J94J0DejC4SgqyVpZ610Y8VpCD2ik6vylFZYvRZ/24ZBtzHbsEbyf1vHcoewnD
n9towdS+P6hCgJECge9HXrFsFYGsW9FwDB91pt3K/999RWmSemMAArfvkwC3s3cc1ExwGSHKJS2n
cxeFDNeEbn0eAuW6YXf4L6zbCoCPBiXxsJZ45hEYJf0PkvXjCzpsVwwol8/ZPMdtjvGIMU5S/BuC
GA0OWg1U+euRlfwbGz7pDfJu66If0I9b32WTc+/MBTvgvMhvdJSO1l18/aSP/FizjtqjdK6teucl
GqdZeMgm3GV5g8+cVVru5INm8supoKXs0xGnvQxwvW6TjjmF9Yfd6mIXSavwHA16e3+fuQhsQq3d
UloGsT6B4WZOmy39WeKkl+qW00ijngny87IDVAA3xHitloDkvOEs+Yy/UGEaNFSwRHyfWUmRT/wX
Ppxw0SuD0mZX3CuPMELt3DVP8/vz1A0OVZiLGLRsDQZZsWRJH/HVd6u8qSdo/8nXQD5Ca7RJObHR
g8VaCRCBpuc9eqmdLAGUFaTyhbi8N+Me7iqpdMqG/fF13V7qE+2kIohB1az8wMNvXgXxwzgk+m99
vPd4BJ6GKWjAr48sytBwPGIiWUHOHN+OzCFXX8QlfKTvJ7SNsTQ5xG35vcfYSAae2vKmsm2lztzW
Ip/xQ85KR0OA0NSh2vGcKN9d1gl9IF+pEnSY0bUvxl4pAFVRlYerw7DmuyMKzkmwYUeJNre5JPTC
miEf+w1PZD8vnIkbSKNhk/8PxqQC8cb8v9QCWnYsBiiG4y/3YGY52nzyhiCbd56XXUqsj3fzar4W
603iDmLdDfE8Zv4VoH9p0M1VkbuQOui+F/JK2HQiDjxnIkzps4KHR6X4YyNu8ITJ2hX1T1kWVM0d
ZcxZlzzZpv3nIkn+LJErZz9VqzfGNrIYtAoBZASQ+6us1OcvP4dUvc+IK8HzgmCUzGVS68pVBgF2
yqTTiRfgqi/wsihouA/dPPfex+yakSv05VuQsap4Yh5GMJenkHBnG3pJXTSs/atjY5FjbVD//jPH
PqxLrZ+CrsP3gTCSYrmyOT1SIQV2i11GKp55ieYZOqVoMV9PfVK2c4FppnPQp8QqZMfY0kzkZHxw
ED6HKeE5fIGJsLy3RCCi9dqBkQ7HJ740Wda7K3i00++4SiZRR1GrXe7HsumWkmP26hsIruxUQn4B
R66FdTM94CzXwoRSutwI+kVC567yT99kvk7SD/PJdws5d6rSnQPwzmbZAEAagRiRnu+hlanumQ4P
0Y1QYj33O51S/w7Lae9DLlWvvb2F727nX1d12jDDmbg8esFlY3Pf9wHUD/FjhWvP12vO3yE0U1Cu
r5/SG1rfKc974Lwoxc7z0LZFrRv2weGQQogiq+4lWhxtuybF52zrCsC1yAovbSARe3JJAjTeLqFl
iCV2Mn3sLfAcQgz0/to8dNMvZj8ZxU8Hhj7b1IzXdD1AWhI6uH0vDhmKS0FFVpnHVnVRwlV7W7hX
1A8JP756V7yMpuIdFAPrlKE/igTejnZGr/kLlU8ixSzY2I+MXZqJuQAb6vwI2AXGbwwGfzXQztrP
dkd+cjFRm+n22q0CpxDyOAlh8d2WuRNKnwMLhuhrbZU4DwRR6it1PD5didYkf/ODOSvlu+K94XP6
fTwNFr9m4+CqNJj0p2zlHVkDGQozfXs86sQB/OK5CVbtp/5ZgF+NeoDiJk8U/FB4z5FhD06Y0nHU
VG3/hZBA0ud35Veaz4BMBby8WHVdNZRKeHRrornhNK83GvObTdMNXo0OuakKIZxt8vrErBzqZCzS
8wJeCj59ueEKkr0XBm5rwTPjD7MevrmnbNxgTyPHJCkFO2ZDsKzsp+gligrCsRoGRPDZsTOF4AL6
McnVx/UxsyfqCn1uCY0JBIXbNoCOnTn7Mh7LCIFfxarcumwHTzj3+2jPmUuNPNcCOrZBm+6rAfwL
1rmj8Mxk1LPfSHznwMJcGkA10lm/Dqq4r2VO7ztoaSLyhIyFPDdbBGVsB/kv6ng1iHaSV5kolLIr
kPMAM1mZqYiMrpxWEarKqirSqWcFRtbXD1EmOf2+8Y/NP+BGk1TWxMfSY0Zf/u3rHWd0CSJujJhg
5VBcYeIkR7a1fV8XyYKQhZJp9XKdeeXcVm6HVQZe7dkBoNeU4ddNxRWGimcngJPdbR9BZd/9Ig6s
tA0NI+uDPa+YjTBjWOGto2IhY4Dz5lqMB4cstgBnak3GOtEvh69zD0+Qp4Q88KlFo4r3z5rRRNNZ
1Wur6QWgwCrRUbDCRrWVF3BnJaXstKJmUQAkDuWuvyrkE1++l6nhCC8l+MnLdjE7EIyUvC8fOaLd
IQJVVzd3By8E0eWjOPvg/Gn7rUhh4iorZSKj9C+S5H5k/BPoDfZUYOZzCbqkFO/0nY7XG2xOEKUD
QffDq1yt385zDfBIHkpsRacvJiH5xI8b3/X3tWpY14UGjLZUFE/NuQbW2eIwL9JBGKNzkYET12uB
PyFBGpFynWlNsMnoVp+4QUwY3OLZ6FjY89AvSfIbQrZzFkoL5M7bCo3p08FYwsGzBwsFJAtE8B2N
qM1gaREGSbhPjBEuNmdj6uK4JCy3ILdF30wEtiwDPjfx1OVsovcweR42eqXGcWqEB3sOYvGFgq3Y
fJKpYPpPCQ/wOc4D0Mb0h2r+oF64bX7PiU60oZvnrp1NtxJ+rQAsNhJQysEJDDkAuChSVFCaSxRZ
rgGPZGiW08GrmS0NkRXTxWGVxxjdA4dqjgYI01loFxRjAhb2Fa+D7MoSYsP78QPQ7YfnNfOPweWI
36ofYMRCc7BtEYlE6cl2i/iL6/8jqMEqwsX0A2eeN5lrsxxhFAtDoTzV7+vbCH0FjN+DdQ+v4KRo
vSfa84794n0ujyh1UGxTQbWhqzdKV5DC4c9iM4UlTirH+oadiGsI0Ml/bWbtFEKygrJ2k3hnkcG3
GrYjuaH4sYdxqTO8sbq9cqrcSpYHvO/dNpEVRYbEhUTMN27ttxlJeb2PZsZNu8V0BFTtS/3zwc9L
eN2lhzsytkxIjQ+WYWEsQpDLMAhhUXXtp5qLj8rTNE7wJMU/H7EedOSBkWhtwWNcKTWOfp8bC8W1
Izz5SVqPaxWhxKTFqgAYlJvILk2vnj/en8TApO5ureRevVcL1MZlYPv4rRwA70KfvuUWNDLS10WA
06Tj7pLxNZ9lrvYaGie8343pK2gy81vF/1Boib5vv2DJdzDNQXuumhYdIWN35cF9QU9OFIz90ny3
w8TRzbeFJO79BEXDszULhNJw7J9y5l9Het3Nl70F6a9+2A6TVY0riIEScWnheMItJfCi0fpKf3Gh
ppm5D43beKDJMqIE/FOG/VcIQxmL//dhL60DIczii5dP0l+LnXORMB6z7657Y+j/89nbWXudOKIW
oOyWHFsVfebcuHT+GRKP3VIWcKguXwlyeoZd55xTkLOKXxGncJyM9jquQTBHMlBDuLj1wZ34gxIm
B9oiwYEga4NwpPKROl3OCQVteYoMxPtqYPnfb/m2UGtEl3V/nplktNsm/FY5XiNccpn/nmqa/21/
8+6RlzT+kQSRz2PoOMly1f5GfoSd1UBE9kWu6Nd0WWKOCM69Rci1hqD4NnAIhq6lu34jBZl7wUHu
pQcgv7Nggy4u+8DO+VjxPX+asI2xMfl8y3+Mc25NMvF6CwLIJoVmtwPjxblNdjmK5KQ4r6NlgJBq
cvsgqLK5qrT+2DkKXeA4lS5xDUaYv4Lz8Cxgtpb2fzXfcJX0SazP2/7YV5S/bLvTUi2h54Ry0kY3
aMA79OFB7Ynh4+NIsbSYv9d2SeflwEk3T4bQDBL110G1o02PE0TOlCS8qKaBveOjSRZQQCWay8B6
yNwBHczbb1gKx+ALa9VmimgylukwolgxIieu5oHRAFxekF9DdiL5enIATQYodiGpckBPy3n4r7xa
mYc2KbGLeZWcseGhBe/xCdyOg5Q6mGivbwOXzeMmMJGmpnpXMv5pNWdusF6UOU7ARyOupLiWrSVC
s15w1yHjTTndrAqrSwI5mwIMODIDdZBjZJJKrY6taPu9+EUoCRbpft2OYQZ/OPCP17i0B/wPSorI
ngFGCWBPzxaVEwfYuGxRQFtorPGWm38aYPwMWUcr+dnk9yh8fAaiZ+z+0ns2opp3GqhXQ8NA2vHI
KFUu+8Ft3k2EwBIAXSSAAGiYdTJq/L/zurJjS7VIMLZdJYADzfFegRHEwqz1+hpPAUVqF0GCPPqn
jLT2zUa/xET7o5balrE7QYRAAICAxMLdmE5zKzBN6LVXoF6MdVgctYOUn9n4BnaJxFwnMIQDnqkp
QIRCycDtX2d1pKZfdFd+squX7gYNVMnAAVgOwEXSSPSRVfTw0ywNzjt16VZtcbtpnmQL/EZ1CCAN
mAbjExlW36Aao+bydiTl6zX2ffqxGlDrC3zZnZeD3M/kERuzOh6zgQuWet47a2G/743rX5XBDS3i
LPDrywGcfXLkcCokKrIfphItgtkgnniQrGlJpmSWukw8EnauyVClovsYSx4nnOvoHwU1ZulCzFnQ
28omZvAxO/K7XM5T8Z6+IJhyfJUQqS86wuZq5X8aSDS46Qi5XXSSMFZw8K6QjCR29S5wKYumKjBu
pp9WYuGK8I+yxpnjjdtipywJLjpgNeWfkheH/gcpng0aSnec6SPa7tOYaMH5hin6jF5vgkgSQM0J
k5Ywm4Kidv4ZmSiV56CGiBSLVABf3WFmvg3JcMx+BIJmTDMrGBwAtEdwEgmQTOmHTc1WTqLEpVEC
11HBAfYk4gfn/wmF99CNEhjiVmgwvHM1gXPBKXduvcyse9CuxRUmQHPqoQY2dHHDNCpc83HL/1DK
5fA+kF+YH+HN8MU1pT6+d3COibuHydmyNNVlK/Ylo2GCrwHSPPwmHRQSLMR6e5IH5Etgb1Y1+Q2k
CZNaHUfcuVI+KG/FwMnsoOwWMM1Bj/9q/ojsNQKV7A3McqyfjFkA7ABWR6tf/p5/RnrDWhhlS8ec
z5FxUKSiCnhxkcqS7LRI722QKqMDUGhRBBXJk+vg2sKzrVzd2uyBInVzXkx+moCosg/dLtOwC2Mr
aHloU8XGk8q+pIePe0bcQrn9s7rQLjZRApKUPkDJmOqEr3jMfQKv13yBMvd5Co0sBW9NrepKZ86Z
/XbxCMW8be0CPbrn3bKgTCAL/Zoqtg/aV34BTfPKEER8hytqs+UW2j+mGTKLurQ8m4Kr6L3orNh8
3UhtwM8Q+VBWbwS1it4R+ed6D7dseTMWPOq7EqUkJcrSN/+53wWa3qkcEmMUEv5IBao/tmybpAIy
ikV9sl7wuEE6vpvdI6TmWzmkOX3/mHAqPNFwCjHHC8hSUBYBpsC3aSfXKyisymLOQo+NdGqVC7/m
dUrWGNSysgb313CC5Rg+B2OKk355D+3l7cjYY8qIxzyvTusJ3VMKWpsgiYo/xssDXQocA9LSN/xn
yZ0TjX5+weUSD+pgHxXwRNjb+Y4BBwldC6ImYs83pVo8GzvUkicYJLeK1tvtYm87Db3gl+2CRjH5
tqPRNnokJDUDJreUVhotuVMjdLVC27oeTcHYLhmc6Oad0jjylVBjHy62lHVlYX6XHT7AR5CnIcSs
IwtRmfseXLW6K+Eb+0hGoZshsh0R+9Bxh02GUp2HzvOuVtxNuKG/CvjGiWDOAjZtudg+mqtk74hN
+y/qrVzWEr6uOLFsGysElLWqaRdIUVyzvWeicYwbQN5hDg6TWbUNn2bt5D52UywG4ygH03ZhEdxY
k+CIEl1xWOnh4d3nFKtx/kmgTN4Z7KkK7JA0S/ctEK2AgS8C7eL3LGUQoW2gwY1yLbSLluAMO8tO
LO2TZ0wIDIiQpRaRTE9BB5lffgZJts8ELAA0QUGXJrywxApp40R+21plsaKb7hUVHwXsr6tJaUOr
O/9N5qbbpNeh5Ag9GUx1QW80KVD16pFbNJ5eDAth6xhdcrdlbZ1xnd/CwZwqDxTRnGhtN/dto6eF
/Vj4XqfragSZHqJgFhnRAMs2u/chJqjVPP1AJhLQfIWzcF0A0qBmsgRntNcszGKuMuQkt4E7kLw1
jtS5ClA7KggVuhzWn4og4h4g/iNlDH9AO2/TX/8sDzUCnb4vr2pjnK90z6z6F3LsCcvI7b0CTDRY
VWgQ3dJSfW5q0Wjp6QfAKvwBaKDqzY0XDkj+cTp6IGl1Y8EqeaENqIV92ybvkEkGrVtui6WLXVPx
2ni+iIsGgyhGMKNG0o4W7S61eJ1jSrEYPZkgsOOaHeIyR0PabP7HrkpWGvocGCbHFseeWx3xjcjq
sw2ekAMoVScT0zahrQRD3+vcKNi8s4GnjCZXEVYqdNIs9A2Hb+q9/7qZVui5RZ8a7jJ+XJyCrEBN
bOm6OJ7DHP8vsi4ywU49OGAVLYFSolI2/TcU5/OSRm/DAiSfrWQJllzDoV22FHJ83uAL2KTxyl61
yDgAPdlYsq6qMpQwh5pl5ORDWESrUkWErI2VcHjwn1gtfHmQS67NVwqatBWMv9HekgE15O9kt9ot
Bvar9fxHE1kZXOQsWL3oS7tq7gNUDmcFGpy4RN/18GqgXEF3gE1F6eWDxKtFL/RtsLnV6A+Y6bi3
Nnbms2RlYwuzlaZVAQ2chYwOpkyYJyat54swWryws49B+hoLh2dgnAy8NftHGZQXlnKoj3vhgBiC
+W+lzWlHBCIpZnAMcweY/PQuTXS85voO6c035LK6VYOqAbm6UbU1TtCK10plZFXeUJwaD2844Kyr
OanGrr5BCQYL3gAZrdTaNkeizURkCQP7mcHinn3i0v+RnS/K/hsW5m6hoxRPScb+sUAai1q4Dqn9
6ZWLFxavJKRM/i7hVnP5kuHbeRwy+wT3ZOepSXHCcM1eXkjAK6lsVnqezoKzIjmOgA6YAg4UntW3
fRfH+MoDtrSxxh0k7+QfYgKCsbXnNGo53hc4M0FPdAbDCyF1cyOvfirZf9pOY3wAWzhMOV6py+IN
eSakT8as7xTtQFAipUdxBHa0S+2dghWTuW6uEi/hobe8qrZ7sjApwM3mo6+jmhyNhfxP5Ng+dusr
vm2cfsM8DtOpCJDvR/Meqc9ffkZ2OIaM40SqH+SkddIH4UMLCb/J06rdJqSHh0b+RG1YcueivC82
6VCTPvXB/IX/0vf2U70q1PWDL3qhBbXAGzly2oF75F99xl/1iYZybg5RleyPK7jsdBS2OUoKdPGR
nwq/6mW1k+57ME4ea7Q0jy7bmvQyAbI7H8/5MKx2oZBy7ml+aFWT88Gj5Jz6PiQUNizAOnprvqIl
1vUMjHUy+9De4cnjYycdXoAAfdxtWNfrDva+DZuFBP5rsffsCqdgjF+hsMOl3gSKiiIGvwnNlwb0
Mdt379wKGiCJtTUMaEzaed0D03ehJ3i9bbQG/5cmHYUXBq1Ky1KROo6pRRBnafmHAO7yG+3MjDfZ
UNeg7bYSPXtuXRk1SORwLGgtQYZBNtx1A9L60DZbUNeBpS97d8h9UybhcLZYJvWs7fE44WX+KNO6
qaYU31V1IlJx6zYehQfW3vBATDeLWUZ30fR7KXJU5PVGmSYGtWNtRvIku+0Y2XJMGyOsIwcOZOwo
m5B3tkxZxlnRl50NfFWfxv7VD8DszlvSZ3H0sOYEHuDO/MpNwEC8+3bKD07fu6INWQ5KpD8J7ZCZ
CWMmiHRnKyxhVF+gvQmNWqVQbDO6MfZB4DAxj0wDEZOtkfFEOS9J1q3IiRJisg+pPTCHjPoTVd4y
hwZSBmgrDE1xxNqRPuQZihJjDXLLmdYewO3UvBfMJ+wtO1AcpX3zMcD95URGuIV39vhLAN2uIWMR
TYRS7ZGPCsUZfqUHmiFN0c8y1RhBw8ishAOsHKstK2rdqqZLsxSbPjNsk7aZVm7xQGka7IGDCAxf
V6zc5otH6UZom6qjCo0Ba5kiNypy8i8s0MWA6maRszuXjWVeM4FTdLC/+hzpuVAVLI6lM8QtFr9v
qVRBEvuwJ1RYYWJyVzZvTdxDtiRVamE77A6g6BZ2br0r452uP5robeYCTU2aMDzz7qHdn7tf5Q47
ygbz8x0JcSuqlV7MZTRV2QBgTBPzqwZ1qjcJmdsbwlMzU99pYmf7w3/xxt9xWuRBXwkIhJF1zhUw
SttxQeJOp1JCHi65K9k6dHOh/Zg6P51oxbOk/VCJjM9jWtnTkl+SQPMf1irxMUfGirj7iDnQT+OD
3s/sAw4EWw4Mzm+VzbJGLqF55BaR+P6XbMkM5qJbwiV2iYGNIL7U23A6f1bLW4yMqp8f5f61N4GK
31w1182SZRNvkFTUN2o9rpy3S+AVr7rZnXTV39djNQSNyd1KaDU27UxvUHgFwyi7uQ8gpIDNzBux
vCI/kUstaw8Mgw05mmTD1nHbQvE0CJScYPEUvMpS7BmFxbxNFJ18BrxfIjMM1eyB3oG/0ok+IQ4l
F2XVwzlTAToZDuM8U28Gct7vEGw2o3SVpTx3AzX9ewcfZSv9IyxUjkOda9XB3bOsWPIgbwRbFez4
jk9bEJWxFyz+K9O9t4kw9RxjwjS/C0Uwq+yS4iKJsigZ5lHHmUqwkrQY04UXHCRu4sQIROn77t5E
11IXxFMmTEDtELQQbMoqY7LUTY9Sgd30kUCW5NmNDGkCzF+3YGkKOS1Z+/aEhAn6kESW+y3DIOi0
s3NGXUU8Er2mqjy0YSyczXVB2d8fgZI5w3Kdm2wZHbA9Zh4LS2WZthPGmqa+wcwCoOVFhfF6f47P
bYj9YZbtas8gK/zQW6F8biFrDgv/AwsSBNo2QbvST8/DVUT6soSEsMo5WTV+0ljmxIoSsAOmE2JM
bRKgPURmRFnFRVa/rmC2gjoqCky0xd2hEB0o1JMANBqqwW/gHpkCBODXYqZS9Sqs0tcmWlgw/vXx
dHhrfY0SpdJUESxlJZ+/gos5IohiMcacC/r9Hv2iRSLJ/aM0lzxua91sm9b2cXCKvKFUFOhR7hD4
PPfdDzxao6xaOQanBrqPF+StcioB91ENVn7D/ID7fLtBLNSIW27N7iPWPFSW8DEOyGLgvaXpAkHV
BY4kvz/Oxs2HjRu+0qrJDfO4gSktkouAbhKEZUe8xLWEWsgE4757uPUM+PgQX2dMl6I4OxYB5IcU
yPUy4nD82fhDdeCuPsRJ8yOpFl/ExyJmJIQhGPMvCn1Ax8cjXua5wKaumTEVRSJ+zKyjeTAZ4lqv
Le7XTqqG2Rb2LMSdmYj2/pB/MjadeErJ3tu9uRxuzRiifTAxvXhwmbCqYgqZGDOhEuem0I4JKSZ1
hMJUjsMR3UGc+bUlAGs6eUZscWKENzU+36RMqHhKTOyVmc7NIm/AQ+I3nLky7CJT6nfQjHS2AVHy
qtWuTOyoK0KmqEPzSSBkY83xQvsEI55LmdO49D3tb4+WoV4tC0vP4CfxQfPyJwR+sczmth7P8Wbu
JGNwyol6m0r3j2CE2ACN+eWrfNlC+55F+eJuhrzAq9b0FxrRc5spZSvciK4Ib3KFZ0d8fwlDCvDx
DL/b3H7N0jSh342hLYoZdpcI04CPsYkXqTuocneIdKq26KmkZEQyKHaKZv2DkAU5qZsOxEms0ffq
Vw+dPhJVbG5wFhylLKLaN2MrgL3bCptgKxO9e26jOUsWWKicfAI19rYsIkTuRNKwN9EDQBTu7G+w
8KZEHzA/8FAfzxLkvQg6Ir8/vXI3cakuYHxFzKs9OvdIKYBHnty+4BVfPbZNx2CvyfNZeAoBc1fx
yNlmOvC56r83kEHiskziX8FNHgXkoIWn2MyrAJ+++YHr0tUFI4vH8YG4bmNx0BW3vlDcpLhEwDpL
qUAViVZ52v2GsZMsyeEUjsjVDYl/s64lSqbBhSHgUuZ1dfTTN+YNNB6KlGRhBSo/DoNoi6Li4fI3
QzstdwiM6cEsL2156pDFmo2EZaMQyPqcv6I22opZV88dbU/ZbOvRoJxTPXn5td1EfXYn2njXlHAC
b1IkyPjaO19rUOzrDgq75N5auvTh+tmZe8G8i2m0WuNuOfazp3U2O1pzrnoLyFG5+U/DX9eNX4cE
lbvteY3K74NgUJQQM/brPo4pgMiNBMeAU9ANSVMEIIDDPg/AJGqxQRPplDGKagyQDc6a3jiLW2i2
PSX7KKPWkQ0TQG8FjbEf8aHGEbFLQ3P7ygeB/x7cfnS8b94asI03T7YqUF9TctnD5d+1OBSGFpxD
04Ew0Apbyeg7UHbpMyzWxW5Xnl+9FT/FcwcGAVwNYf+SRVIR/AH1u6HOu1a9kauIYkkR5GlZtzR9
N+jQSBdvCODq/rqP+hkXRIF/yysVbih+1MUSw00MWobPYSCy+IbiAWuyp2ECPlC3XdDcp8gBCUn/
e5lMrk9UwhyQEtcylkE89g5axlg4Kyq0HqoFY5Rr+ojFlwCHUwNMH5mhyxgUSPLb5mJe7SWmHLcM
a5QACgkmOAW6WKxeiStVpKZNTInjitwflYhVrDAW2YoBkM+K/7nMNAVCo1qoUDCIGmfVpZbDGEf9
IQHdknejwYVd6L0B3MEGs8S44qNoPExnfjXtIMRfSuhRSQe8sLmbpbr/tpXWny7nrwlod3+gwV8P
NfSO/9jhAEsHrVB8twav0SDQ0d+CX+6kocYVpDpuWb0ElY+r2QWclwFCrN2qrt4fDYm8iW2Zx+Cv
YfszkmDzeMmeyw2VSjB6pyXbPH2QcJdwpTGWyFcRuXa47KFG8TvOn9GYmDxMVjNFYDyqWO9+B9Cd
mc75GjW44Oiabj029y9EehKoPUVu0rFuazjYEojn2ilwgoqoHRQm/fLYJX2cIraP5Qz+s8beBjFU
mnCeGEDRIKreMma74hWF1FMXow6e/fz5GR4+QwL9Onq4hijecbkOHZUa7nC0EwPo0wUBoyhNtKyf
OptQpA/DkwjYgT+ZX4/mzQ54FQBZUh9vVdvipztr/aijPq/2lHWwyNPnNQ8qtzhLk6EDyyA4w3B2
qgUjROCRlMz0XBB4q9f/4rTlAVxlSjpCIEcWckz5gdscsqfVOJOURWyX4eEpk1tlIfJ6gLn4HMuK
QiNodC0mjOSdAKZEvMkLBBAipPvvwBZ+sa47VEtLHc3FyZm+VT4OwzJU2HJz7f21oTsx/Ro2VrCj
cItuCh3S+es1kut80gUvbs1Pr6y+lBHAjDucIJDoegH8w54UJmqZ5rE/8vAOjzakgGz6YKYzrZKg
qw4/mIoiKS0phRQmPnaF9vp1uG1pV2kflvNglRAd0beH6qNAnCRKzaVzM6zAhm4i5KWSX+A65jMh
VX7f1+RfBCrwby0O9+FSGAxJMae/1Sns6p4w15NKwyY7+FL9S7ngo7q3d8SP0Pmv14NoWXsTODnM
JgURhGrsGlweulA22QfvcSNObFQoQRcxmyV6XRuL4xSCQBHgG14CTBEUzFipbj3i2dbD1Pkqk5r9
cD13qwH/gdcadtBdWz3cU4FDkba1YmcOXa2Baa4a3VfbzARZheqyCX/inG3ZqYAcXM6tkTINCASV
7TJv8CczEwRPA2zPmflaTf55gcI8cb4yLHusWTwb/E3d9rMY9H5uMQ1SgRt+9vlnNDAHFMuZ2q5a
6BmbJMHkkjbCUxlNiMzPqfqNEBnBoedPC1RGi9xW5TNNRFlIhGHUN4bvDzbgLMtXooeAg2UJxAo2
zdi+MJW0/9Cmym99kExvdiiWuOlJShfb7jPCycqqB39fbRNfpLGxkhG3WOUo+I3hf29p2aPtvyW3
GgSr/0e2I5f2Fr4ACzT1g9SJzqO+VlcKUM0uvqf6Pwuq5vO9RIJrJA4OHi61bPSVMOsjOKZpLpoi
S/CGHKPmGNNYkBjkASfZy3sgkVqrK+8lBB2zQmqulJ0FNDFSQL0CnUBqQUZpUD0gZY5rOYUbJgdU
F9HjIoQDKXkYrLtIdHsEMd+ZakXgq6XBIagcOOpGVcB442AEsvh3FGMSt3vUX/8e9KMQf7/4GV5i
3mbtw0OsFaVYphBTZL6MH9ogsxTwDG6SEI97rcR2bjC2xgqYYCZ7NR3VvayTNUdGk8ljmaWI6+Hx
MqivYv3K5htB6cdD8U5TggUEHxXAxGIgPg5mQgm9kXqYNuSQG/PkQP+1UBf3J/JcFTo+RYw7K018
g6v9W2DCeMLT7KSBx1b8wD54vG1Ino8DHMMjVWAMdJqSwNcAgwrG7VKs8/94dI1lbNpgtMCRBuxg
+omCeNDDWG3cYtfwaEYksO/X6jxS9v5EOuCL0oiRUUgoVIPCfp4z0U9LADjyB49UdapX4Npvc3Xl
pXw6aIrydvtTRfrz99UlrThp7wYhCzYA/Q1MgEI7rJIDJ2PxVDAKpXVUWpiDtubUesZNyRGloO/z
0GGZZxmekDN4g+aUMCPNKNx4NnwVTr64K+Iq8Q1kGSyjYpDToNiymW+XMu/9526u+MHaGye/CMR+
rRIJOC7Dx6GkcHmJGq0QFWV0x8bqjXukKMRfmoDsZRC2jpmW+LsnVAV7nxPJ4xpDm2L5Z7X07vPD
EnlMI/cfwUU/rPT/oh8hgiYFEjPHVzCW/cNOSSuI9KRQQ4Umz2ZMfzfnSgrykCxguU//39fksaf8
OKuaYvDNwcZn1tXMT27cIGtfD/pjIrBR1+z4N7ZjqGQ1zfEK6M9nNGp7Pe2GlBz+Zfb+TuoH6TPx
D8sBIgqDrVTgx0O+sE6eHcKYAcmD1HEDJ9qzfONw8s0H2Nzs9rhTYkNuOIUGjIIFrGywz3LEm16D
QClJZfxUBnNJYzgzPh+WC/CQ/AKl475faFBtQ+sayyNcQx7F8cjX+GK53rdxsEZXUib00CNb1dYg
3S5jabLxwYkK6jQf+pg87nCie3fcJ1C7fILMNd6BpgBDokB/moAQu38S401hmzbIPJgLWWb4/o1o
Dllnui1YmWP6uu2172ongAnEFUhIvt07TzhhFvycZMfc5yJS9MvGjM+arCEJ3UVkhonSl1YlFv3r
E5fj9KC7nTg64dYXgRN7+eiTaQrzEp9K0iGHZMpgkRxBonAjQFRc4bBS7pFELtly26Rz+uwlSTa2
iM7pmqE0FDzGdqVu4iSCjcH9Ceiy3lfuTeJxxsUGz4YMZ+ieuypfnSUXydPhd0zYMT3Te6xzl+45
cYlAhFJMMeATJTZEQKen347S65qJzoaPnXESWXhVI/6GfrZXuGA426HptKocC0+vnkn1WfwfBMRt
quEbx7U6FKh6Ecsbr4EMkRlBAaV0ZRB2TTjbxUNvmsvc8LiwEII8wGK14RCXr6H/jEo81j0t4pgx
CAynuv1wm6+cLT5H13e4lKLXpfcTZ8hVhavBjRUs+zs2V5uKDevKHXYwKF1/8ltkk21QBU9qNO4P
VhVrSAht30qhuoWtHd6DLCq8x1n4weBzQVUtiM7Ia08ayBRGzThU8RxM79OR7T1Vbld72qHNIzrf
s47qApkB+EDI5F/WWhrzxPNSoCUBWpxt6/aKPibqO3yhSWRuNeH/GYqURXPx0JfOy7XWXFsqdapk
M0QGGmr4Otj1e3qg7twBMI6KZmDzfhf+loSIKehu5km52q/o8NqSckSYiHFApGQNsQxGDq3kVavM
/eM5dCjKgq1fs0QYdHrfCAFNyX57PpVg5orA1anRgjKeBMAVJx6AyD8h1dFlML6SrJzY3i9DFZi0
azaeDLUwkyNoPR6TPXBjQtmbgJj2wSpr262VU0/7FG++jVYpk80WKxC/rJPlCsxAKY4osTq2YbZi
TCuzaZNasWZSyDLf/OkxIEUnWpvXBBpDFhkOpAdlE+8jkWGKivlNtdcZhtCJJZBg/T7GYi705aKl
UpDsLfa4DuS2NObl4/zLEfyHaeReZCKB2HNMMrYIvV39AebL5j60fUJm4jR47RlYsThXgHWHarlc
TpinL8e9LMuLum5LPrjsbxyJrfAom4F2L74UHf1ArP8H+ngFP+hqmkUTNrX5MtpGi1AY1GA+oHi1
7eH8cAaI57vq4ARtazmAj2dIreCKgdvk3pNDdHxnkcU/FQ03lxH79Fd2GjHuXNgsW5qDXkUofjuk
ieFBBF1RZu241teaFJKc3CimG5swigqSLO7ZKiCRWVpHN/vYoTpQp1JGxfqACelUPIBfrT0+tSS/
fZeDOHo1NvvAuaRInVihqsxPB1thi04HqHE+0yMxYDcRs/g7+x+P7dr5jY9JCKxk5ZN9hPpWNmz3
DhNivvfiy3jHvM7gI0rkFNdtio5v62cufaOgvD8l1IpDnkfmySy1zRwJ4Suol0V5tvZnQhXzIZo2
G51FYmAKsYlKbwHE/tFQzHupSmMM76da1mIge2I5QbQAIMDmWkDL/XJka+4HvLAAcu2qoqwhPIIv
2khqVdytLv8DBf0cJKescsQVcyWzG0saKlgpaUYrky9oo+ST4zJEjokl8YKwNT6eUrV6w9rpM+gF
PIHA29CUbDdktiWHuFqrHgT9hc0qQw1Xg59eOwC1fxKhvRMIHNOvAvbYjJNGbjVM7dxnE0nb79ib
dDHQ69cn9gccfu3ZouwOYsQ0B5QS2WPcLipJT1pAPpWNjpFI9W3/JJ25Kp8v+SpKrRx5sd9CVQfV
lS6C+OHktTq3or/Zi5DL6m4ACR8nJf6p5wixbduaqLeQIcYrpDXYFjGV70TeclmYPUaH+THPZyGP
d1f7exDl6Gi7jThuvJ4RspaTd9OI8ruGs8AhJDeyAlFhAGDvZEZNDNE12IKsrrBCO/3oeV+6sNau
8TNKdMm1CcOZdwgxj4QqlJBIMLtlEjdtPw7LIXzbQcbXTsthD0E5GVBibr/44I8AQNMAZkhMRbPP
7d7dVh2/PkdB1+p9VAjP8Mo2oXM76v+YpUjJJTr+qcexs19rAI8uLT4yy97Ptmbgiayqa/Zhtyvh
eFwy0nzZIGwsXCSVhpQbILPyGzNk1TqCiFKz75vICKaWfRmtzJ4dF3673rrM6TXG2C62TDgLoXfl
rhEWIr07cKaejtVecAW6IgaXsUjZfDur9hjE8zmPaZJBy4XVBv0JE46z+4gQHD29XPO74TO3pEec
Sm1PglAFshrSVUwOwrz0DfGNe/td6VgnkBx/QQalGlnASAgJggvIn0ihqlRwMpylMar67tGN4lWp
CYO1zJL6Qj8BE8nC2zuHWaffDITZxds4W2Jv7fROONbnGWlSo6FCERN14A8ekgXh/8ZSdTMM4VZL
CQqYRBvhXicE4IDFrNS/Mb15VKbQVusnjudnwV2fecIWF3ZTrAdV1huoDm4qESDohawRD/p2LQk6
5USP66bHQNygmbnm4AVdQFvUcC2MHEgnYfewVcZ4XWSDnpanNn7fCGXr57HNaJBBF8LbYzWv7te6
UdhHeQiE+9SwU6V6afjDP+g+CvW9J1gxGqM5WvWc8JS/FQm1lrT9SQDP6Zf+TFJVmx3MdNAVvIBk
NvI4b13/RlL9MczDuBeamX/hXHRJLn91L16lgnT4x7NBMEPdaD2mmMR5I0kQqVH4gyLVD92vMuZ1
e5PdOeL/qbNfe8EGwnmsMPTtXCdJhSpll14izS95UagZqOd83rvTY5U/Kjhn2WSrQ9zOxKuItVl2
ESk6TRcNhjdK9Y0o6l91R8XzprXufFAPHlsJ3rOi8LFwtWuicoJyPiVWZSuqq6PLOAsES4kt6tiS
3tlERiZ2g0PzuNcqgdD8jcXi20LukmfYHXINyGGoYn2h1zgExsvWhgaQPDbZM3pivYhunQx4MOdP
D1ZgcNrAhwGUOGH5Se8d4GUClZtEN224+PMz+ci+e2O32tX+domcmgB3FMpb4VB1NRZU2uxfQQck
EhW0xze4QE3Y4lmdzTsIzfCnqixodjjlmkXnoQ6zNor4vIo5n4rnjJ5vgpWvuEsQS29xadlz0CfU
6qqASRno0PnqlmndL0rFjeSG9VwFfpYUibP/ffspcXMCkxeomu/kJKo4LoVQe+y5CEdnVpLcR14O
6njJ+3k6cr8yxDhPjPB8308bEOOXcR/nsWGG33UwAdk2q1g2eKyqevrm17UA6jcaM9auDtR0xvl9
BTiBo+iDcbg7eIkfOpl6CGLHIde1CCvGhRvOetJExd+tiQVr9pymbzKKHjeqmrr4flZE0C8ph7Bg
4nQC8D+4JJW6L14auMBSSIJa+6OC7FHFVbgb6nR/Dm21HM32eBYx9ydbGeo6iwcGEXgicPpAEr+c
vZRxZZ4xYt2tQWWTnMC16+5O2JRifyfE4cRcgkj1rEwCeM74h3f2/P+xuD3IY4Lm+ZS11KIdKw2q
0NxBbzY2Fn+9YgdGFmeEOD5peq3UyqmQ4GGHJB+Z8pcqhgVXQAMv0od9O2znm6ivldg4SJqwL0Ft
MRATuSy13kJqAuK8Z9dQI6tzNK+MFBBRJrAyQxgGEp0k2+VErx12pf8oCpWXHg+vc+6mhLQoF9ee
4J4peIc1w0AWiuYbkzex7IfPYNkWwSUW2rKElXP8N3pXs1rJ7isEaKs8Azm1C98mU7d41cqkDPtc
Ca349cQN7Gpu9pyx3gC52Mh1+AMPsqqDIN+yntY13f7HjGwWT1ZcMqgJstEf2MLQG/bT67cjvnyH
AF+QpcZmF5D4ONhhbIBCem28zsrZJ3RhutUODEKaXgznzN+A28/UeZP2W7bXSMT64VprlIe2NudO
QEUOmrvRtLTEi9rRlXQs7j7mkfkSuXD0n4YblSPvwj7FwWx3DJIWwAMwstRKhZLwhutRRmW06v4N
lfJuKJkoWwLn6Q5clASysb6JhsQPIF50eB82gLNgaOjQpT3Ubtu2FbxnS4WPcGghA9MFhm4WnLj7
SEShSt4dD/Gbf6DrFOvzIpxAPRGR5+fxnsKXjiKZLUlAm1uO+8l/qJ8MR4poDA82O0apusKnPrVY
BcuD4pv5HZRH6vi9ifh4XHTlTpXZWCIWGqHTCG45xLiDLLn8ABaCClPO7o1qXWFlnRfkHXMW/ZIW
a/pyP36lm/MS4ZBE6XgOh2b7zNMqKP3Enz/5EISOzKq80lEJfRFryGp/S44W0fFUzQxaKdtXInqY
HwQvaTbYmgb/SSMMshcsp+cZy4P1bOTUEitsjH8JLTjYRbK7XCYC9U8/l/ZPN4x6zokC0j6OPVis
kbUYkEiX0VcVfocC9Gi6X3Rrr2HkBmZssT6G1qcLMt8oPgzYhUSYU9U7WPaTG9b6qCeEJ4k7GBcQ
YgBihss5sDWsc+8VKvAp22Tbwm4TPDcTrjUt7X0uy4syaiXdMYF/sIG+HDg25WZ26NC+S+09CYlg
KBKmwvVv2ncC+wmxxVGIogt3aLwn7np5mN7SZS/M0ub79+hTx/cEgKfqVTTsIyMKS9+AiQDt5f3k
CyIjnKPPc2j10mQlze6W/NU+Szj+9TmFQ6/cAHzsUuFpeuxHQXNyQHgjDB8W4C+WFyi/f7I3kUbD
9R0lSqCemVfcKGIpphE7BPaZLfDDjPunnLMB6ivEWbO4I1XB/aJMNBP6IiLFAATH+lm35/Vp6ssM
bWlZB6AysvFmtBQTdjCEBPMXEhRl+h5p77EB9mzgT25Dhgizy9PHoxBLe2CZg5Dc7D1XvENWD1QD
TbXpJ1x7dJfQDYDbaXprY2b3R6kXQiSM+nlb+9FvKHC1Ppzor1pPNp3DhWX1WmmEs1qjX2CMPKmI
k4vauY9C1VVky1miRnh7ksi0zCVNAkfWXzR4mmcRmidXczarsRMDFp70y0enSJMhSxCbk1dTF7xk
yuZs86KqlGG4KAFCs3cZ2kq7t4bGMhI8qFvE0yRU+HQQpkXDYV3rfIraW3DHHJcJQGAjXZJpCT9S
03TmXgZ9rk6eG7p/pfuhP7U/1NmPmLB0iZ6o34+QKamfNT/C6da0V8262zzQtQYhF/QRECF4qtUs
aVhYonLd+bNQGsafiMkDeYQ2kSPW4YBc7QuNecCQludEP5/W2vKdB3YBV5ZCRWkDz/DUIbb8pIYr
dQqTxTP4bXUw7fEqdQkUQHwgbCgCmyzD+AwTiQAHl0WkM0kIKjggiRw0qG6R/UhS4rUvoDbyWD+G
Pm+ZeeCl+Nifmxs1EAN0s0n1+P5rh3JK6HvojTg+cZiRD64j8gQalzVyvTvV2nbSB7Uc5l1LPAMR
/PCHnZoj/WzossHQz6WwyEe4ZGJSp0k++aeIo0eiOKs+l9ydY4nhIIkmzbXiNYn0rMWDZ6KYlORR
mjvRT2tOuQ6i2B4cuwejgprIggJImZs9v1vj70Ojr/PPst1wJ2wvzLfuUq9jTej19sSKk1NxMt7G
fH7Wns0P3Sw6gWy8moRItn6mSZXekgf3tXXUFM7oNnpaylDrF9tRFn1tsaNl4u/c2HvjJSuBnj3m
hwN1YWpmD9Wt6Rtqr162WHxh+PmH4/Cnpm52enGpwZB2YCi1OhGPmt7+eEw9+B+pWo0MYElCQs/F
1RQbhOyq491/4P6TJy/aRZJiwdaURNxir107JIixpcYcMCGSqOlAF0dSj1IrG7Mhiv3bEYPpmjFw
VrXTgiond25geR7VgtiIIuuJ0qLSfb4REtVtlpubLxSos9NU6EDyPn45My3Ez6tt8jPr0M+oUm6/
Sm+1SmhBJYcR78s/WMOgznzuIcVgfBVXo4AXFzwhoM3s5IGRn2akxJrcyDJjt31Y0IOtM36ZKpqF
RBuUQAxOGQ05BprefoB4PH8al85imT07PrTK0kyuwwalZTUxkKL6j4pxPJoDkEkV/XETfSIUBdvi
60aEvssDY7MUvWNuvfuq/25JcHieNG1ByBuqALIUfqB2SG8Nu+jrWD9KZcs8cfzICsptxplmxmex
gB+p0HNnkFcq4WqJQjn9JQQlxIH3NekoTX1Q98PEVgeaMjbWxSuXQT6SWXLntD/wefYNpvBivlYE
vYP0Xeb6XPZpMex65n9bkPi/3XXz69j41RPuNELCQZbWRyIh9HGfTHytaix9svmN1wV/PCN6pVVq
fTw4EBFlQ0BK0R6yLFJKTTCwDZhAyPUOTCLSYjRby5tNqdv8cgYIlV8mlAiR3YcM69frFWDxJy4S
anK98wNuRXFXxirFZPWdPRQakrmA5XKX80/3RkdYiPf7rIB5OeP9AlwGDfydKKXNM9Hk9nC0O80N
2thkVACiAYVNJwhLWGjkoX1wxgw322EfDIdZn6C858RWX5dT3sxLopcjA2c3G6fl75gs4gDZf8R/
ZvgOlM1K8TGsRmOwco7OR1Xaos1IJYxaDARyOaLodJlhkS2I7P3QsVG2BUwsWF5L8ubQR8At1Rks
xioKVe/53cTIbdsB0+OCIsfJ7CWnlVrEFMBGSB8VprAgBb7LDSUXEgup3iT4BujBh24+M2RdPF4k
ech13HIRJojT0RvX6uL8+/dsp3Ihm2UtCghIWPzZ7rM+0rz4vZ61L5PGHImU0zrsC8icaiyNBqZD
njR0aGUFlQ6G6LZ67W8niytcmG8WOzu5zZIOhYWkC/g1e8iQJd+Mn1cn8Xkp9kO7A5s6PIYrE9z6
zpCOGXw2vL7olrHjrfgn9DFBPFMhBuoZ5dq7yeWvXYkyISEF/BDe1KspVRkirYAjIDdNkvIjRb9x
hxmiLlLMJIQOYK4TM5fzgMtB4Np+czwdxmK74EzT06iybn4aD0EYpBl3SXJzfRFRP151jGEQgWwe
qWD7lVG5KyZnydw44847pL2r0SlbCio46JstQujGuyu4yVxZ/2JGMj7JMOwiSkREr/eeYwewm38x
2nfXIJzcS+ueuQe8C7R175cvjxU3zxd4a217vDBUrYj68gCi4jVSv5fvKr8pmJgKnCt9jDw7Yjwz
pZ2w/YLtt2YFKirruj52NyHaowmJa09YiBkNu0S4O9h55VYrhyquplFSiGCGcVlmBSbRKmtCjaRy
5eZa7CKicWgWmWt6y0OMru39sV4G8Ro0eu1+YIuxnTeghFGyCY3cZ/pXsMuh7aTM6IfJqQJrjMLx
50bZAOPDbju4bgXNvT4AVBe+PSiMwKCPpkAP0Xc0GL6GZqKzRxYUlJaJalCeBk+ff75j+QWT36+T
3BjtaOTMLOWnrQIj/Jx1zz+H+h3Dk72GJ1l9a1BaNjVvN7w9xofMxHMuGTsUU2IYKe1tzxg/16lC
aABVbhlLNsXL/Z2pkt9Q/me3b3BQowaMQstH8pgnIZlbnHxsbbwTP/3gu87la7oYED6UXL5REr4G
YqIfJugzw1FweY/W5EGzMDFv8jjjg8jDjNowkbk3UXBwEj0Du/B90g7S5Xxswel3vhwBDEvSQOSB
IdKZeM+u/ocn41qPl2wsYZg+ht0ZH5AdGiJYgEJ3uYxCUNZpSbG2bZkh83EOc6opIpiEyNfSybdv
VGp2I/uQttp0Y+Ixi4utCkEH7DExbTrsUzC/7J+Fv4/Vqg1GbbCvzKEcROIKjMlaYgWXjD81lXHf
4/qM2Qzrw1NE/YiIKwL+zMMjCLXhz5cMFjRVce/MVkRWTYW/anmYhT8GPjuEl/wrZ51YBwQBLJTn
2kxe4o4M9o/GkHyhuh4jSobYP4KDViUXdW9ifpZtkpLl9Qah8RhF6vjoYmgfd9P3qI8fg5egwCJL
zbD7M8vSbqbzcjXCvG0G5tO2+uZptnmgso1Uq4vzYeZQLir7cYftdV1ZDwce7hp+U8TulDw0vv0L
WT+yEsIwb9XXHVgAgKTGWxVXGPcfRujOEED+RVStG1RIAFNslYQdvnhaJZmvEO0vw/e9QoM3wCRg
esXoEWAaZYkIVElw/JlEP4z8t8cuBwaP99wQJt53/J2CKbcR7w8TJ43B3+5SppskDALYX73CfRBW
AiQaG7Qjxf34el0JSvhare9aBFT3aqpVQSRwpz7roANvJG90AMYMQst2DET9VSKI/KcuGRXfVa4B
FlIJKfA4hq4b7o70XNoB7iDty9JN7XDOrtEX/enTu7JH1gwUmwafP+sB3PU8iUb0pn9Je8r01Z0L
7cFcrjuidoYAXWjaQKyoTj6Omh8tIRPqa9n2+vKm8A1RHkhWObHYhGxl4ZjaQijUzElQWa8RzOJL
uMBPCT6HOn4nB/0SXCCwIA7V4IhLwm9oVaY9290saxx+t0kXKmFklArv7pMZItPAzAPCfJ9nON1D
8oZJj2ZJJ8/u8djPTmlFAQUhsSd5BxBQj+8kknjAwU5IHosUR8jLg+5FqH5mLnR1RrEKjqUatGrO
UxRBHCFH3okxwbEoVtw3Ih9mlPsOFXfwpN6j90Xz8P6vdAcTCK8A+ygNqm+TL7jgGIhN5oSnngRr
ZYWa90r5GBxOrlX32o7XfFyanoyhS9CMBOKxUT53PS8XFLt4SWrWtWw/o/varNKF1iZsw4h3Xjyp
/pww02J0ofuXoMnfCTpPDHHkzLGUMP12OzD95HsL/Ajq1UelSb6PVMK7kW3WmtHPMEvXpJTeYwgB
EuAsVR2BUoj71s5eHHjil/ORctHtDB9VLePlZifugM6MDojwB+AGNvIjA/b8dYsnrvCXc4Rb4rkG
WBy5xGTO8PwFvHjswYw2x4lg3/gW+kB/X7RIoWmbhpfNgy8AvkY4zm2C/rPlk/1hXSwlhv5Z+d++
7rJVcvOCO4rdbzZi1xCt7njJZ9YVBAqhWe5pUbMMx9p/VeeNz8gouTVho6m95v+RrOrWw4J/fCE0
cJ+UpoQy3ZAhbtnzTHOXDEJaa4d5N8/yni0V0Dfvkfva+aG2cpFxSls0mV1rpdEJHnlD3ta4vJ3s
tttj57o3EhxdggZAliBJlkIvPVWNX3ZXlkXtiZ13nT+rwTpXzQCiro7hGKL0+ssN8bCzRZRHEGw+
wEaNNbS4VlvojKCGJvDP7sK3Mn0mDH6YYYQQijDXVpBMmEro3NCVrHL3sSNU4oVPigZXrzS+ED9G
8/4Gsvxu7IJhyySyvKP1BYgR++spgasOAcKJzL1ZBnCdVqfd/JyPKGnpE3N5Ok94ctaJHqBgYFYJ
qiwxtWzb8+4V4dITrHn3Qpk8NnIqIZ6ZEbV7xieAGX1AThj/Igqwk6JSxx0mbSE7EGOXi3HhGh7O
h6Zvm6a2dg163uQw1YXHQha2Jr1Usk4lSArqJqHZKIDErVgtNsgaQ/fdrLnh3ODHqT3/+lhXVQOG
N509wvozu/qv5bcI7LhHhYNren0WGVt7Bu4gm3A68VXd9PDji3j7bov+frPcr3BNzGh8d+4o9d5s
1/sXCeMu05jnd3CDVGlD2h+9gdH1LHyPGzrwZPYSEbBRJTP4ET4KkGnMSF9TKbVN8YM/EbuVD8c/
ObHNHfLmnoXSQkXXbQtGfQWBGhftFIW5SBNSr8DGzDe/KGzV1JeplRwsFV8t7tlrluOrdXVjRtWO
I7mLNBXsXutlEwkfwPJmPoPeUHFSJDVbCiia7pHeK7QYMe5UDQY6c0kEIT4UUfOx3jvvoXyuXsnK
5YjWHGIkCvjVk6jZCpSNumX6DNqOa1Bg1vYFokr5Fb2J/k0+N41qc7iO2w24k3H3c6dtC1ugHnM5
Pi/hOPAFtp5plkRrM1oBuDxyyl5Pm9mlp5Rfpmc9yPcZ7nXKXze8Zbp/WNxcyW7xZgaOSphDqmBF
oae2E2YQASxIrkJlT2QjGriZsDlC1ANlMwJDsu6PQl60aiCQjFmsaw8p2YLIQ7YMpc2Btn+JVlhh
76pbwmVLEWKpJYwptpdJLlFbpHOmm456Jk2M+Vk8eFBjMCqPrgMWMpbqb18sD4ZxXsYa1RjQM16C
Csp4mU8mRsClaFW1PiIpXkq7XX+B2TvZ+yA87IyBuAI9TaEK7SpL5sFtvmpRPaJ/XyUy5Q+pYzki
DbsMOqtQcWPGEcV1sZeGw+uj63w3ugnl4m64Oy7dhdyelrIkEpGa5uo4aAog4LmQ8iBUSuM3sboZ
1DiusZ/l3v2K4Lrwx8F0/l468LD+kSf8aIZ3//xnJTbHGbzP4EYtXHMf+Rxg3GaGu3wAlxnoPb9q
+n0EB4ioEKGpNerDT/5PIbkHLE04gxgeSQ+cgUZynv41zD+A7YAP61FrubifoOYYyAJaNQpV3BM7
bycJbNb6i++ju/yfjZNUVN3Zf+spn3L4FpVFS/IkqlxYwKuJhb2Axo/1OSXUA/sZDweTU9R4GQmX
obD+8a+/2KS0AViXHdSk7QHTuev9w9fVo0BG+lG8ppGNBIlaymc5/AVnHQDjvLy2mBPexdQdFfa2
JDZcaE+Ji/3aSs3hHQGe1x1J0iEeFIPnFJhwHTDFCVq0Z6/FE6+hwiLW749SUVxT2FFPA2U7Zp+F
BCT3jEWceqv3PPK86zNZPYm0jMgCnbxsIiiKIoR0Qm+ybsPFjmzvH0vLYGAtzpKAYxutCpDi72CI
R6VrpyAuNc5Ek8GlnTaM1muC/W4FzQQxd7dq6gsQXufRvQQuZ4LRu/Guj0MUR4fDIJy1b6DiL/9d
YpSzgIb4sDGGjuTa2LfWsge9rFUyU5sjQ2XS8ogPdtKvSzENzYm+kXclhWmRy2DnYG5HZlOp09nc
cFZ7PiCQLE0CEtgKnPoIvDubrLKgY1/F4d1jPGYumKa1CjjHZr8l+pK5PKscxjIz/9F8ePRx/tsz
DvepWWfCEG5ASmWPKGAsBhVKfPnRNER8GSd8dh4vJwiqW1up2iZLTN3tW85rCR2YIt3WN1MHBztP
sLPvMrx/0IUKVslSYj3912laUT+S/xHUJGA1NljX9+++73hMARxFxX26ZdJ56UoJvM222d8wdzgJ
hQyTLoszm8kTnOT/dZxFdxHFYC8yIEaSVu+pqCVwzIinY7KnmngIUQc/1R8elZJRXywffV9hH2FT
fUOIy/pLnaGNoGlPUFaVlhxaLOPeasls7Ti8RXxSc7L4HxcRkF/YTjppvs9I+aTyaa+VQAyy07tE
ILKRTWiD9MZ5xYslDa7GZpI91TubqnyKfRdhFRqfSHvfiHsMjXhcZwzlGU72WjkX/hHr4bnxpRGo
RCNbrEE3hVM58OYCEwlLJ2XpdTAb6duxxev+5kwtwibLeVK0z35sKpUS17yNqtgvk5T16tVeVzWW
Lb1xQuy+m4t5IT7q7Lkz2S9kmsNQ2Sk4zuCaQ95KyudoUIDlkWbaoQmzJPha+AX78diK7xXusHI7
97K7UI9WDLOeXEm3gStcQj9LUODGQFIf0M8VR59hJ6Hk1rRfvYPzqMdPhEd/moCdTfnvKZPBmjya
IzRDPxvOiexaGVHpeXA8yobK6B1S/FXNz8haqkn6y2uuZHPVtZG56/fMHrcGyd3BNJVVxDemwuL/
88ZE8R98SThKKDMAucd+9++nZpTWHiw+ZvHXqFQgGT8znowmI6znlb0iGyuMWnkL8GSqNn6AG/4o
8YuqigQQzToUX8Hl6tB6qUzgwbM+XRcSi08rOlGfr+1YHsRc22032nxOJOPsRMCMsoNjb84QZ4Eb
LE4cka+pcRjTdgreBX1SfZVJYK9Nqu2KZLXbT5BJwgZr6rVgqGvsdwNdg7hPeaKGXdB9kGiSXq3j
nr0ZNpVbepyu4CcetkxpPGBp1TpdcQTjelk/AowCjsHOhCLTQ+OYUTbGYxgFZUhr3Px2U/y9Dis4
w8clDcVVersjxr0x3pRQ3J93j4S4JPL1puPQlTLKqaepd/OayT4UH3QzxC3Wg5jw4RMYEzkw0JCr
YHuuT49y1DvJruwnNbJR1yU+3u/+M/ATfH/d+2N9L8/Gw9f5D3rSl/8sw090+ov5rfAXIJU/pQma
jGHUFog1i/3PHzey1HOkmWSc30Efw4FIQMOsYiR+bqSEgIOsmoKkLz+PDm9PVRHP7yv6OXfQibCg
Jbk51nTv4QIHmqCp60jtPrsx9YaCuUphmWccBRLbehnMAcKrb12HVDR6qt13khSxn34foxNbWOHh
F269i3XOrK7LXZ3CHf8popgADiXjJ8SitOwMTFAqis4cO4oCwjH1JEB1GfdJm6H7xejig0PXZWOo
86RG4cDlqMW8WWszFavU+0DIO6HJEKzCB+tUxYiR9EepZ73bdT4s6J34yOmtXp7GBMQ7VALR4CXE
hqpkTy1PJp7kqO9fM+MDIyCOJItqLb2d4dQA/jrLT21Pvu9B7CjOUG+UnY1DYaEqvhQpmQQAuhUT
euWG/YkOyULBD6eMFkc5m0BopvbwV0PjIUW328xjktvE0lWMDmG3y/4GqbapZeMgcUKQv/+q6bo7
CMRFhVDOqHcmag9j7I82mj27hnPjV3K7W/kmOZsjy++t49vpFrrz/ghCj4ZRXjzPp5nrkKOmZRyn
oG4OFFrrEYqvtR3FCBWvxWJYvJbbQd0jTP0XHAQ8+3zLRFQ6bK3dt0AJNrzfUFs4i8szqu9geFqa
d8nFF8VpEAmXTG764jCPEn/XHaslfb5Ziubqz5jaFAsHdXi4M+oyKEakHq71XkSSYHh0EPjMz9U0
2H52wgieCzprt5qGHAPdarrdHFnpT+WdOeWsdq7r2hh0mwkDkLT3vQiHzl4uu6L9qnIlMw5K52AC
4mqzXf9BHhBKe7x9oCe1WSQYpY8YFveR4K86NsOkmnQDry6yuu0HMgNWUy2ee97rfmdwWPTle7Vk
05zyPN8ZivQ0nCx8hUlowrYt0De7CyTF8f1FkCIxvjUpBSf97H1pGxuaA/1/R2uDz8wzv+gksFf9
SCl549+FrfC1f1DNXstfXutJ5ayXgqsQuwqYdDx7msed4pR5UApVmfUvPMl3Yq1LjQxtwbgk3VKz
3qJMOb/eczA+31zEcsDen7Fn3X7TmgVynEvKxLCswTw5uGzNCnl1BzyaFFP6xprP/YC5zp6M6CUJ
zvv8KLU9ZF2KX7rYBmLQ8c1rbjfxteI1I0mqPnk7DzgusyrtgWCQMfv2rAa6oipfyCs4LLt27AUN
8ytaYqVVgQ/a7rI73CkYQmCkm9/6tF0Nf5CXW9NVcxEMIaP7KxJHxcjohy5myoNrxXWvLNNsYaEi
AAzhR6rfdPaz1zyz87FTYTQSr/jth3LGL5W1LPa8vyvq8pnrQh7P9NVnfRWRb4lNNq1F+2vA9Nzv
g5lPIfOA/eeY+Hb+7NQMd5O9594xn3wNJ/ERuy14HSUPqgF1jxok5V7r8U5pIY69+F6C0sIXupO7
5gP+SJc4yn0psUxHZYUhVcB1BuVEKPtEZIraZku4MqA2cah8jJpJEL0LVfHwmIBhgbkZTjM2r8iE
UvZGZhKsx/bLDMCJ9Rm+BlmZFh/w2SnwWNYJ5pOwTHUPO67yiHd3X7F+iPlDCKbK4BKahWuaziq3
8bcyBCwdXkLs2rIBaCWixS4A9qs6tm2ZUM3kLpLIBk2hWMP76rJjvWFQkiefC4KQiUx5sVOkok8r
W+sd4exFWuCqfGGElUYG/kI+Wp29UZVoBHjbOmRTrQwtfFvY3bHtsApSf56xAl81VJ23qtlWDx5B
nkUoVwAVJkJ2oG+BHEcenKzx4H7BNJj51Wd+C0r1fTSpDuGsv/wvplHt1QtcxHImtdqSmFQxA9TJ
7DZsvBiisBUq3VG+FZBuxdYilhvWW0IZx1Oqwx8dP+Gk8VKF9tcn2zSPQv57eAvHNIucDnG2C5/U
vS6amDKoV78oj7EZ7qZCflLXF9XaXB2lZrnR2bw9MZc/jwfk+8AooL7dfIoVjeRZnT+1toAcvVde
iE2D9otAPGRMIukkXwQJjSuDtYZ06d5K4Up7SSW/srzCY8LMXv4PbJVvdpvqmRgCB5bpmkOb5Mkx
SYhP3RaiR241pb7+er3XaWWExZxivq6vZhXa0kaF7zyiigMVwhRFd0DrRQNxR1klS+ANOh6xCJ8Y
zWJ9AMMWLJdjVzPdIO5h3WQf5r0/WBaaOs7+QjVjsQ2rHeRkPuPeBy4pS7rnC/EftWnk/ZM2QmGy
YXGY3mdpWR7U+P7cA0HuTUdzQ3hwu7NYVRPXPiXno/DLzJbNw5dratcGeMj3XQNmF3lpBtM2wICm
ZNTNEM82Nq2kEaDQOkv6sJXq3sJTCDs6GA8CZCx5W7mU2Y7ZjQ34VQWIGOfYIpVAfdqZCStwBPqv
UVBAyOnVgzRCp6slowcaI/pgedzaY/kPf2jIeBd19bOuSmoKdBOiUMwphYU6O7w8RCWPlYnSFV8U
ilgMZWXMkB/Br4ki8nexYxxxR0i9+8A80xxyHGobtqm2CwX/erWnw9oS7dYqZ2IJpRctHpgpQBV5
qiJ3Q/5ymOtEeSKl+vA76JWlU3L2pTkWvVEf+gQLZjj52JaihLjZJmZjY1dpbLB/HpJRVmnwahEo
nEiZC5shD0Mkjgmi8HcvUvurGICTcclPRWvTnrPfghurXs4DnXcbEcT0e1lGpptHnYoH/Df4ND5M
RBfl/eNSaag05YgVb/lpTnkLUkG9AatmseIsRl/xoOJrx+1MH6PISPk5nvvRnEEIG8xc37pdNqVf
TObBBGhkgxmjmns2Dsl1vDsiyC1KSdnmTHLRgx1huSI0UBnDnZtI9UWdh34EmyuIRBaRujPvAeS6
LG1PbUXoxxz/Z9J+9qE0RwEMz2bLyvMR18gHUeozdWc+sdTOjizridluW5LQCBBRTW9xwvMIp29R
LPEt+o+9plR7zrbFc9r6yAPOfL4s1WHDNWWLizlxTzAMrnjY84fNAtE4k/lVxTiAyG3SSccbfnsb
ESAt45PmSGY5gvCNao/3qEqHQ9Pmj1Q6/miwNd1A02LdBTC0Pb9ONhNswKt4lAyjKBlgED3ZyV0C
aesqWxQL0X+hatjcMgc/vIsXWPzH+CKwCAW+N6KCFX/GfRMmqgpoiq7/KWnCsksCD41Q5ihkUppn
+oT7L0nxeZ67k8RzVDkvwZFYNF8DcdoXVBUNBIB5EL0iQZaLBksJSVextwPVtJAOitWDks6fVuNF
MYnnRn6pZOvKkidcgVt/FQsPfamcmTimwI3CvwSxYF4c6DM34VCoT5xihsZ2Lm/fbKb8TyOm9NGg
PN2E/yMhgKulPidE3bkhzS4RaNe06wzegeTDI8sbkat9XRpM0csdFNwOlFhbF/31F+ZaRi0z8lM7
TbnvYQoBGCMuu1cOvvmHFDRP7GkAV7icaUCTLIuHhr7kBvv6X1g24sz6J1O7Yy2RaH82iCek4rhg
qUKIO1fB1+NBoR/xHP+GG9/4iIbnKMfP0qODYdJZnFslOkGMeAEtN/pwd4vtqxDfEKxjOn8YSjGi
X5MAJWjVV9q4QBzNrL6fQP2hi+rnrUSOv1cIryd7n0yGkRJhij4rABK1HohCLl56sMCadOKygVvd
TSbiphwPIrwAUVDq9LKgKmiXcwIBy9/E5l7gTiBV6fY0Hy2TGLT5yYworkQN8uZh5XCddg+CMsMg
Jg4hIiT+dOhRxUI/qLAvFwSywdZT9j6/3+L/Oukxc8NpJhv+zpGe1aI5wCB79zw7FxrPqLDBdrS3
Pzo2gaJNwURPXSqMnQbJRu3M9cLfYawrKmn1okmhw3nCvmGjQHJJsQfFu5JSXJABpruGjsCHtCCe
wOY2riNQpGvYVoHwT2QPf6+ymkBS34H62rO5O94/WxEl+RcqqxTMIWxZyn5dgV4DoXeIZr9YdJFO
MGOaENQlUcX+FX0T/oTeT1HpoedBeUYvuM/MX/LTaec8fvbXtNbVV0HDlXKRY4sZXDr0Lz04lgYS
O9rEhgWqnC69QYNizuilNnq3rtIXbg+keXuUUm5vKQfe0tbAa/Hgx4Nt90/0lUhb7LbdJNUgHEwQ
HtQ97EG9Gvgff+/S9tFtM1bCC1M9kKjBjcD3BpcQlZftEHygjSvcm9RRiwtAw9rV2NfDaesaAiEM
QEcGkMmcAinzAYlVT8TsbNNsRqAVhCkKYI0/3O163J0spZJRtOvrmGWarCZFJmWqSF0/trZMXsjk
WeJHWhccbvgqPFaUhXe1x4nSOhdAxuHsgTC7n+nXqgsXp1r+5zSuXYZRcXS0ZdyChVZx+ZIEgmLM
x6zFYbiWoeaU9Evi6Jb6miZLz7FKVXAlMXfgs5qJ+NrW8ezp9AbS3ffreootrlMHrZRWRREOkC7g
ioQV/MDHxq1+dbj35us70++Dh06cm4AUNEDDCmjvtwGiOdiCbpHt869zU5FMrWpdWrMMSocTnEWy
1uJODhp+mxeh21/8juASqrtdUrbCYu6/eM6ya1PRFibk7rO7l7fCBZIsjYi1V085pP+EECkp0EuS
aEAzoC2cj+QcPnd0tKp0DCqsE+ZZyzIHCjljtK8iOgGVBGffM4ZTG1lrYBhF1sEsOy76r777T0nd
hyzfFUx9AuOLFj/3753he1ppxBB4cNppKiB1LKFCaydVTzFBJGo7pjiSmsGFvg+lCQJgSKzLAO6w
KVNdsqCLQCmo2c77/KgcpXrhfzl8uMjyWuXPqUhlBxsscfVVg0yVw8/eCK7ux7XnSLKu6sFJUaKW
3hvTSCByXRF228TZbf5NIsSJtXadut5IS3KqY/3nnOAuBnm768BpusP0IbhTqYurMUs3DNuaVU9G
wxMIXnNzqwVCHpgGSNX9ACsIzrkfHS2LU84frW8Tg4IY0t/sEezbJuH01oxO3hINgm/o9f1o8j6o
4oSQycmgj2Xg8Mb5mMT6B8AOondSfqaMhJtqbVyU80C1tWWQ1tCwF6PmGGLnV5erMse+LpLnQC4z
5MYAzzY7DtSFU0tT0LpKkW3WsOdiOj7Nvj64GbEXkgs5mF5/POcUgie41nZOSbWSXA7G0dT7Squ6
rOsna71YDqvlodnEcKMJG6nlWgmJIoH6sQB920Zq5fcp0tViUkz/HgibvttsRyTgJU8ixNUlK7j1
8AuhOCy9x33ZsAM/590IQq31VJyukBjteWs3RjwVVqipFnOwRGrsXHruXkmcHMfQVzxrpQXB1ka6
UFq7fEyT3dXTlGCvbY5yA+qkq/hETSp+wi07AfxkCU47RC97wvsH8phO0ijtiDGj5P1R/L0gt5EE
Szno+zW7SAM1UPNHiaTcyUA/N59sofx/C26I6Dkw68s/OWZ3rLMLh0d50tkGZo3LKRbUvdRgCr3J
NUaHHgdkZVEt210JYzI8dIGvFr+XzKkYijI9WvvTPHGPqKAMNtsVxpXRV/s+NBpB3Z26ByB0KzU0
PRHe69pcz9pbZJOP5akaAsB0SUK49+utx2JFLgqsbbPfJbpyqMkq9nvrVKzTIjGryYFtfLia1T+0
/HnQjvsIF7EeKL7YTUlwsP6HVfVeC4hwk3m+IdNZEW+UBrkoiBiL4ep+4UA54whxGVdgOat3IzNU
i3QNZXI3u1YM5tmQfk5X5XoHH/vNj07SWkLCgihTjv+QNqtPYph9ecXnFziodk1dYADZ8+VAOaX2
7/tT2O5WXIdFWbnRmQvy92ZRU9w5JfaAWt6ll79eivcVBo1uicXYprSXxxLbr3wmMvjmY87ovAxQ
Sgwv23PzlU2DlrOPxErHKvOnLdYfpjUl2mAAN0v7slT21FlYxEuT/oiIrbZXBjiTTuSuL1MiAiyh
UY1P+OI88kXyfO6Wqq2zMUUtRdsh8IvnlQfS3sg9Is7+8VNAzDddRYrrIgAZqo6MquuWe30vnbqK
utpI0Vh79J3phnBOlOa1fETZe2FP8PacKn/NlFJbpmzrulITtzPzivvCeyGVOgoEI9S+TqO0vICN
AEY3ZuoDjyV2WYVv9Uouhl6lm9q9a9/57b9jp9obuWJEABuOk5uwn3h2gP/P6jMaYjBxSMNQKNLd
isaVZVc0UAN/sSjVa//1e/kz8bf34f7lSYSJysMeBjZPUNRq9WlLcgWvULOPq0GDxNSkUrs7Jzzq
E2+eKRubS+uJUuIKB4qescGu5E9GXqiVedf1HiJXmkUsUqM89LZOZpnBbQrF4vqZezhLPzx+MWP2
nIpmyhb65VCeu/MKDYivfIryDyZU60EaJLGZwaGEuOrcsf6ajE6yWolA8lsIykjhWrN9prBHl34C
5TrU0iWFFDt13Yr3u3GvD4RqSuTrnxdoITBO+efvm7gTzB2P76M4RP6wBDADNymadtcZsuW4GFta
eRCiYjf4pTNDiFlTz+OQHuvd3bdHRTVTM6Wx8bkQ6vsQLCAWRmjQ4buid/TDp57N3lDXUNFMxT3U
zVZzDYvxbtktsKNyfmebm8zmDLd9G7XgOUn5s9vA/JXocl/IpfZplPiI/eTXdvSutuCieZoHNuOE
8WFPIDOEe9OySGDyoJQ09AWOrxrpoFRpB292M2O52sPqhl24C3ZxeWOXfPAUyukhWgvaLIUG3F50
KVmUSGO6Oq/TGajhY1Wp4dQnySILIVUlarABi61MaPWCuteTCkZk329u/9Ftl+5oph62nXxvsc9z
BgRXiPKq2RXMRFydV0Ndz4jk8gnhMtoeVHkq7zwSPUw0D5zQezte0OzifKtRVLN6wnVYSPJn2BY+
NaSAvG5FpKpBlXl3eKcyxCXdmRwlilYBpxgXtFzUJtE2roL/DHDRAJGfeY8j3iPbRWwqsm83rVhL
IAdiqj4jsR6Bp4rm5RpxO3hl5UDpyQlbDa5K1C0efTmXww+pbqCXVVD0l2ZGnhX9vdKNqxCx1PIy
WxTFU/1qYTfz69uqSroXPXdA1NHc/yPULvzBC6x66Hv1SxbC8Kt65/tIyuOsEoKIpYEBGx6zSOwZ
KrYK3yGUJVdGoViwhdpn1xPiOdjAUI9EK552i88POPPr4zzA7I0AsC29a/932kLnyEGkUZHw00bK
KxMb/qMFkVEVVjysTPcvxSPPCWS65oXCTIqAPQpwNuo1A11MjRjWwoQ/VSPz4EVDxbKl8ewgnyuS
29p3OIUKoo00lNeLmV/72EnzSd+Bx64U/2t5n9fwk+z44AILkZldm6XqJI+yIKDLOHTvHeq4XG+L
LnHEeqyhZ1TFX3PnixxQiD6VXxe7CEwabc4Q5VnNzEAOHgbV0gL6L2SPD/j+ZOzCYeGMqAK0faUw
fYtp6Cqs/O0Vo7HNzTCQ1hB/mkmYw8VzNWQQeO3oHy9lC/hOi8NZ5dTwyPPOZIDg9nTgby+LsCYk
lS+YnWnfRQNxakJDTvklQawlyS14Tk4IKucm/B11fK39gbYTZNk4QW67pU7NTZ/FwIxHEOBxXTP4
6aoJML4y+V8A7aL+dmVkua5CcCY8EoAiYqSuTF7iVpaURTkqINaIR4YVm8PkfwDXK13c4qS2VNbL
MX/sZqjv4K3mzYUKCLRK/VMHSQTyyCHc/3Oe5oLqyZo2E7uHi6+A1pEU9tZmNPjOH82Ib+F/wJS7
mHI6ScqvrqRS0ey+8oMv2+y88A3RncLrN4l2T0gHTYwUi5WLi77wXeCsghFg4aTfW1FgzkXrhQgV
4SRfpPzAeIz97wbqQxWMVcQ0DmPfc2XYqatkeTyLGAsFJC2DacXUvdR+Xj6G6PmZpighAPMV/qn5
yPS2X+7u2UJtYfBHPPdYtt7Gfqqw/kqUUF/fGeWpETwAyfhZA0ayKBWe79yo2JPG6m0nQU+fZZHA
YvaojhQ6zBJtwLTgDqq0zuUYeAuyvJBl9i5/fCNkCClvV82X2OvexkREwLPYlplz6LpRFlu3CguE
ah4kEpujAdj/ez/CSuMLg8T1/QPwYfM2n/wFxU1tgWacAZfX/GfzL0mFSPGSNr6J1iVEGJCNIGkL
K+0xeWZTscM37lXJ8FUzb8wjYZBuNO+s1PRFA2Ia4YhYvVbNWTycUiYlCS4rrllUdYdBmhmqEoct
tTQIU8rTa3P5PMmOHFscXpA9FlDlAU94Tp9mCGsSNeWuWJx4blWVKg4o0wA324EK5Foklg4fGKoK
ISlVf6i0wvex7K+QqhYrocVM+DfH3mpYHOdhjsP5pxX0YC9cf/RDz4NHz4t1GZsYlbGykZ/Kmm5c
00gwBd8bJlT4PAA6yAg0NVPKK4qSEZME5nVhBBFij6b/8tZhMqANFAVxcWj71hscRAqrn+J3Yc+0
F0Yjx4YCgnCYtlOupIUT+6rnSe8y/RvICMqdtHievdUtPhbKtm00v0+BvTXLEwbCCS/JMEDP4lWr
T9M+kcNSXVU6P5iUFg6wPzCuUYgdifi9bx/8JjHD1sHBHfKMtDVIJBpGTZwqWYZUD1P66hpBjdnv
BcXv7YMrS2HdezW6Iy5dvPLa+CIZmcb7LLp2UmsF1n18rfbazwy93IHsNxBVOxyMItuk28itctWR
eX5KM46Q423cR2oTbT3kDoB/Cd5AQcWrt9QB3o1Y033O1uBrx4O1zQ7Jm65JJy7A0b4M/IjLluls
G5zZ75TtUVq2KUde55thz0p9TowO3AgyNq41EpeKXWglMstORAkAGwabDGexqmjl7X2wLr+jgXOX
thV++t/n5kIiSc8+jj6AXoozG6eELmqfV7pu0ZJjb++vV3/m9kkqs7zqZnzeJLXurIX20kLK1hro
5zkADkfxbkjXDcjmKaoyfLnudyWkRVct3ztsRt7WVOqYETkyjjRkDytJ8wRux6++4rRwFEjvnMcT
kqnhOOGQfw8eeIbslaEHS8/qSdmIKa9dcu6mdH++fWvNxOf13RylhJTmJVPUBAwqJyq16LFG9dNh
5XOqsoTd4PNGsy9Vt2RCH7i4VzJYi/lS+KuHvMY5sn8hbEr0dABXZeYSKkqPBiBvjqAtnefDvUHK
1SbOSYKAbG/ulyhtjQcKZ71ObzSKjVQuAJP1W3zHPOBLV2T141ukuYc4U+QCpZAMCoLGITEY+yEE
6hjb1KunelcdtOM9lieJ8t1NnodlS3li7FZIEaVRghpakv6XI7iRuu/h1ANbfzFqSPD3v+aWmXUk
4Rn0VmdhfRS5asld/NjGEiuhUrDhXp+v9opkBqlGsF6+bkqeeOJlm94zemRjYI4EKRMi2C+XxicI
8EzcUxX2PfuDXCJyD2OVGPz1CY7u8goedb4olKo7IKkqQ3iVnJYps06s+do3xAG0TQKhDe8GFGaP
+WNAgM5DfP2MNrdIoCugt4pF7uiIyF365g/DaRVtL+KAKUuLDafVGNAypxc9T9nb2PHWdJIO86Mu
cFVtcnyUykMsLKYIXvdBDSbvchkyb8M6K3PLa5Qj1J+Gr3iziXDyVgpTngMT3vBX3aWaDFie2hXQ
Y3Ga6xlmXDrAmczSGAjfVcIQp/cqAD1P0SMtx9XiC3kRYLPkNYD8/1SnVtbqZKX3SXXHy7Vlk3YG
73VM6jrdhv2HjAxoXs12g0LsLWOeckZDsBK70j+q3hmRz08n7EJKpUbfJ9I9eQTdVKNSHes3FGbt
HoN1XSmt+ZBMvxxlMl5bV/Bozx8Q7AoYLSwexyHfByxCpJwJigo3kOtrWCWNWGTypTm/ClJQN5TL
2lWIRb4cT8U27+A9DCk4/oAy9hysbVPjfo0I578OfNs1heo23pB3S2DyjsNkdK22lJVzijEVz4yv
faCYatUjZR1bqrNr3r1XW1Mao0ou7EFdmPQ1bl4Jd98Jjmmp1t+9IHwSwZ0F5KQJZgzkMigyNEac
Mu1R4A0genbc1ahxBSrdvr3MmsN4l1WZHQxdNkgNYKQl3E1+zDqQ12SwNavI9OJTy8AQidLc7Q9p
pXdXUhJIE2zNRMdyYmMOsddXaQMKStnwqgy9wk9/ea9dmq1GZiXvEKSVLm8axLjsB7bBTKGUphH4
utEOksmFFCkJ5WjzPhp02u+7vaNqoMRSSfLUr9aW+gw9R3+PNrFZOIhiQtmk7sHLmDuVh0vG5uhT
AaTxhvOaPWSTEdqOOVHSCI82oQalx0zcwfQrDva6DUmjpnz42KlfmNTRiX/B+BAo7EtR11xWC6Tt
BGrJEVaFsJeA+ZyCZj240M1Bt/eXdiK6hOxuk3MaV/0myFdmVNsQBPD8AdBtEKcii2Q0vcE18bFA
B3t6trCwMPPt7Bi0pa7wjmljac0YuZ+ZvHP35D96lzAXu9S16K4vVRXAJw4aj7L6YbnfBaLKcBYL
NOdEtB1f3Cwbm44Fhhh4senhqtyB0Th3GxI6bb62pUp6xfZ6QgzsorHiAh8t7pF6Zxr9z/WQjx9q
6tUc5G0IxrkPcMT9oT+3BUYuAmBKAkYO6JuAw74B4GJPHrDngsoUYIGkmeAFz0SBiCYS1uILmMUs
Ake6RskLiR+gdo91RiKoMhj8R7b1fbHWJowE+NUUpYQ8OLM6u5DXvxmy7onn+PPtGRLrCBHwc0K1
UXIyPuLRLW7PqiZzyWHGbmbhI+PZaePAmPLBDDB3J+QnxLJZieKooCBp/RN+HZDGpXHklkuFP3ed
xAsjNX4+Om8/mSjtZCuXhjzQjPf73zRD+JpCkMaLvlvCWxEdlbIGhKW7dhOxSS7YGRwV2ubsEX6S
Pmzubm1lsWSTX76K1GKgJi9/0Tu0ZCp5KU9UqQivEtJWkwAeynskSyos8ThzFXLnfxljIntv8Z6r
jhpDZfAu+ByEwR3uV2Nrk4gmQzqTYD+SZ9SbQdeqri1qZ5csFKUY63jdGe4ziM17+yihnrG96SEE
ymHAtonyCnSCbXuXGK6x9zxGpdhmsTDcH02iTZHYjOVgnrnMwG+bUmpGr8b6W6vNsUrH506jA3cK
6PzIT+RRPtVr+2wUaPgTB8Nh+Hw02HmKhvy/ZCh78wE396NEnpgEMyRzvj5Cs6yJ0NXgNxZjiA2T
bmuvlN5EIGxF4wTIlbWdDoe82VAMQVSUagAxunbmeKWORjg7hoISVXCJBNS0aCVvcgu3pd8U0HaW
dGIT2lNCWl7xIB9xfh4jR9N8C4fxG2n6OTJbbuIBgxnhMPbolQeDWWKZFj8TcpRXiV/D0YkY7Jev
p5YuilJ6RI373uD//vUJ1i1epgGBSwJrEXg6yogBqz96bAFn56hpxdN33bgU+RpYoXqJzqYkCx0u
THEM8uQuK6fYsuxFL7w74W73l3lwg710+Ll9CKSszQtpqdDZi/JZx7AAtw8ep0X+eSNE0S+TEEaT
GrVLZHrH27LRhhVKyhbwcut6kXoXXKeNZsHruHTffEM+xBLMCMdT6LK83BW1vT1/g9XGPGTIZn2X
eEXgsQRsHijj9Mn7RgYIXfyiCUrTjHKyt8GUd5ryFkZpo7PpQ3iKtZ9ZJUMIH3xsNPo92XNGljlS
Y2HVQkWvH4V7B6zQDSGrJd83bR6mw7hZYo95YWsJfQ/dc7ey7FfadqDIBwO2fjRNZ8lm60brkjEz
pMXYQCYrqWHKauXp4HcTvuCJH1uN2B0Q0nWJGAaJmKNOUnp+FOLBrHVpE6/6tnxbRnASoVR28Odc
tlfPhqh+arH+A5b4yx44kvIaAT8i68p+TQKJuML83SrEjkBsqGG73gd4Vz+VZF5fqttpY5lGK3Qm
oLZl4BpZB9S9GBmzpCoSMbUJv/vKVLUHjDYlRxUEuv2KzGB4dfEIkpSb8FM9ZWvZO2IPg+QWqgEW
PAPOMQrh5WAj+E1B7YWIWGqKNsARQt1EIiU2pzZ67AwL/Il57pHk3XjpPBLe6C7BK8oxfeW6exIl
+Gc1EAw4IIDY1bYLHWutLOEdm2l/cRs1q/he+yfrQFP6CQSfTsJRFSbUzPoY6JrAcyKNSxTt+zEC
PAZgTaNbgp7KqBfRgzockA+jzdq6rue9qBQDDptovfGJnpGi3irmndoYmkjYG66nzWvH7jFAgyzl
rORzpMXvLVCg0fzS7YsNFniExCpR9ekAF4MOK8eLFxjBuy0ouYB7ittw/3RX6LB+hXXaEcbY35c0
qciHQiPPmJvQ2WPIJnIFCZPQyznk6DckDx/kG8+z6qIQ+9D9SOYOVsEyc1mVdkTwB1F6kEwLjN4Y
dQKIum8hk9G6nO54fosxEfNLwxEmicUC1cC3OPnZ06nILKBVXQEqG4V428bWuaFsCl3KQ38QXnTs
yrBooMS62EOwWsDj14XHzWustq1szTdGCHSMq1093NV6zs8KEY0DJu/qpt+ngx8VHkZSq641gZbr
WjH8pI6jJi/zaEQjKJ/bdgSb142ZGCSXSQ5gBD1cr1nGkqncIOkj6/yDQACoU/4uNGqy7YJkgvjz
EI5ZJ4f89VPB0vpwXMU2H0zJRoaSJWRSPwg0Jp3jYcMzUw6QuK/kIE34Xh0sqllLqWKJX+NxTEWn
+cWRI3c/to6cbxLS44aclj+bkCkNRws1fYvK7WVeOXdTheZ6k3N/IzHAVDx+GCrSoDfGJuFTSdk8
tf1d4F5R/xx3ZtjyDaWGreYbStn7MZaOAk8yD834VnTNzW9tG/8QFc5RV7DNvR8kPjTWCNk7NWSd
xtHhSfqoXa58gCc9L9iHxReUa0w+Rw3kJfVoRX31AhMxK6HDOv9sU8RktOTPVRNbx1N/SGnbSEQP
eq1B2ue5/8ZUTUoZi8vlbesFqIJT+dhqwegDrnuhjJBgD9iK455Xt72UGAju+4dbH2wWpxd37lfm
jBCV/p/GMCKBvq7eIqxnXJ8hbvUCcHM/2KjO65uuMP0iaGwH29i+0nORKcxnntaFetR6i8qr/nCL
APnn+6ua+RYWooWWf5ySmr0fjxpyc/7bzqcZXg/5IcmrcmWxF2Cvd9AfS2vijdwNff90R0jn8L5e
tKMEGW4/SL3KeyvWT9e4GSXoCCP2aCpB9R8VohKtEDYsDn2WfTSzzTV+pNErott7rL3aMcRD200f
sZomU7qGPinl2wjw50p04Hs9QLRMctMBDzzWm74WrOAziPhaKtTM+6pwehS/idRQQVdxdiGhbiNy
roPfcqOdOTUEjEMB4/sOqCReofiDi4bdJpqsLohQDkUVA4hpW067a3UKLLBMmJB9Lg29juHclX/s
LEksXdrr/gfLD2hJd2fBl/EQUd0SzUCqtXaXA2c6Oa51MYUdrHXU1L27pkNqy5akTamiwnsxz2lh
l186bQKOui9F3IqzxP+QK+OBhg4IghE/Uq/Djlrk2/EuGfQbJF7oGyMhRA6i0264hqGPPMqqyMlL
E/1RzpWc/9rzm+NKBzMBjQHT3kwREPsOorOKA4PDhQo6Qk3bt3tpXcCriL+trZiZMD/r2iYbL52a
C4aW9Nc/yM0hoRpX+v5xP22aAN6n+XUFAT4icXnnPDZzy11HkrgNm3KiB+6lgkkAFCA6i3kd6MGV
yuZ0qMb07FR0tRn8/qITaXYPn53D6BSr6DC1hSbMJYMVEIQfyQ/I/Yur6OJ68SjT/20uDwTyRH94
+e1WejAShDf4O/fx+/Axui1rjb2VT/Qd8YJ68cL2IpbmBqAkHqHNtLmdlcFkVH4XOjzn+VPXZ1WN
aQ1M4UfDJ6QVJOa6b7LWqORixHu68+ZW4ejW6RoqD/N12apwIybavyF9Z/vSVB2wBAPVfX2XTHLe
Xr8/uJ49OnLlzwa1MmbTQdiOCCHKqi2Rqe6qhGTidcvI3Y7/b84qwEUYlxnI5/jzotTNEGL9ueSx
AAlpmEqCRqAOVRgPJoqBVGk9QPWNa77R2QGdSjVk4R8Azwozex4eq0Alxx1ZWM159IB4UmXCe2ab
2QmTsIRuQmoZk3FfMsrg3cGf2buw1eVltB/RwZnpxvJqQc/f182fdGBZ58c2GgKrrfEJNzkTQLCg
Ja2+4QH3CU0esuUP4r1/M0qhHde9rqe7757qjDlmg7Wpd8rDv1c1oysLtGsrVBRe8X+mB8ji2uqn
9Lovz95BhmgzfiqWPP58fbvswoUjySTuekmTRmMYI2A2+39qF5DfnXeloqk12QZIvifnWTIUAeFp
56cmi+RqR50h0KmWyDb3kzDgUjSM6Dkv/qKL+rpNRn6GrpG1nX9cgLjy5uzOmZtOQByY1xADMTlT
kUR+V7RV3Co4ueNpXE3TC0f0AvUM1y8Lm+QZnZFCQMTvNJn/0LDrvWnZ9ViSTsxGn2TO01I8OeOx
+mhlIRmm3e6N/T3zBEkgOd7Ey5y45lLM5pZUcw4UYrjh7CN0wph2fkZFGwKsoOnd2EONC/9yq4RW
OEpZve2dtIzOyD6avFJwlEUIt2NoL3Jdx+umsXiI1SwJWv9FxxhNmzrDuyMTySkNYQUyG7sAxIeE
sOyCHQlGl3rwuTUpbZxWSfmijhxanBJdU4QAbSD2TFpG2nYJedfmZcBbPUz3BpKDshgniCBrtaQO
V61eH6kcc8mnskaT9tmZManYB0lSb7lsIZHkhvO1emlkY2ZfUlkeFNmXu+t/wiNeXKMbgKdzaXwH
w3FvhXv2wv+PO9KQaQxvm9vsqeF0KkGwZh+i0r0J6vOtpbi+JYPNOKpx0rwXA37El/PudsqKZrHq
LPo89gr90EpGLScNx8dBSurCCy1yC+qLZlEAYuZPlNAuG0VI1pKwFmVn84oZKpBdJzmEjpUKWAeW
7NN3jcwk7+vVA7FqEAiklhwRnQB3z/Q50u3eZYkh++oG46l6NsUA0mKsagf3Sbu/BIMzHHqQn3ZV
L7N7e8mpW7S2PKi0i2F6gaSM7wljljrWyiVsnnd9kWiaLTRb/aQANQD7ghP2tqpSd1+cw7igEfi/
HxJVOaqfHYv5hSH3Q/B3HL2z8OcZTnPqo0HWYLa8I2HPdh1Lm9mobycfMhIdMrGO2MRsRru3GkEa
1Z5R8D7TmgbKGa5rfhCxSPQ+74nWytLoKhVF2QXShdhEmtBii3Otyj+MucIrnA4yAtcqZZCGgd+n
tL0Mb38uV5+R4obKEYGdFtsn8tIRnc13xlKniAD1rmdtckpt4Jj0hYaSDoqmxrzXlXEhIwgVx6Dt
+1t4myzW2u6q0jZgQfD746/OxzAW8Xg9hXBS9AeWylAjLkygvA+3WPvdf7qC7eBgL6A2UFxxivnV
NjHkC97bvb7RqD8IDUpyx7K1ttLh0/HaFyuvWdbgSHocJpVX31XWh48mAqL/yWwQfK6p3kHv98SS
q6XPluAFsondHFnWYPj6Z06AsX1+L9lwkg9r88EFUKiDWXTi2SxybsNc77WsqV7ABubBfuOcFsVw
/6/CXHe8HqvGP8MhdGlSvg2ZEf0vq2d1bdptpSXS7l/MIiy7PhfUxVvfXarh1V82DWNJfGvAuBXV
CGSHTRefFS4jpcQI/IvbUpyy+U2ybv7YF3IYCh77nLQ7xa6jMSH5H43tu6/GPneC7ONjxnEfbRB6
BG1D/QWEhE4PF/RpQsVJpe+NLE05fKq0a8W1rNwxEyxZ31MJI1tgEC2PKzlAC5ngcSyQoV/KkpCY
Iw0wGPuO58Wvlam4ZGk4g3mvUaQOHnIncSIO9qQnS/fLtLDl3Nf9Qn/mRM5D1hmQAyZOMh+BHjFf
JU8vvDx2eJtWYHWr1CVMnlLAY5/OK9BIBtDLKVXgazkqRqOpBSS1622762QHxUAd/+so2wG4AS05
ojS+bxsKI3WX1UJvtWBqT8Vjx1PDkBy5cVH7IYJVAxRj0381Jr2Y57EZNWJHaAqcUOxZ/Vg8Zrtp
8/GiR0JgRD2kNPvnwErNot0uUzJjaJxl1vGFd/F7n8bAxWEwaqyQeVk7BvNl9KbCRBz8/IsqpDnf
WJGo3vNyzWDqlYAHBpuFcDiLjRibyQE8vLPxUlQqu2KlA9Fz0NsJX7rq7b3vrCCRs48Yq/vgnmYu
STPaLOY2Xg8LSvsNAI5M9vQzA55yAEj1wcWYwAZKGwAbSSfv0PBwqoi70VNQwmHPyM4o6Nw+e3Wn
V95n1YOfjXzQDOHFBhNXPCwMjexfjy77vDKak6wz4cstHdOofad/0KzREZ/W+xNJiTc5HuSNM/Gg
sfU7Hoxh/eoaKKqsFpVgPN0n76+c9vSbJXIvAg91k9nf/yIGG9QKwZwvrXNAyemZ3Lphlnpkff4P
5kqzIkHO2FSmOiMMbaHG7fQMxFMpsUxvIsk4DSTmkWJVdBQ9DR1ERqODIAdx6JJMkBYds9sYCMPG
m3G1rLQNAwa8k/g2QqQinJDDwK7RhMbpcGOGDTWK7oA24ZdZtoh66JzWu8o8eqdGjlDhjSHAq16Y
mCU/N7vjMoJFxoR+mFXJ9Xt+DVQn+RavVObi979rneuDVcFRs4r4ERI/v4Qv5UFX+cRj6mZGkfwS
lHph6y2EdQ+I4Vto/4ShVjDxR5+I8UyEU7iM5F+d1FCBF+QWuyYnt9D+FO8qmrnlmrthhR2DcxIC
1XPDCktvu4vyw0Qq+t4NYS97GfGCEsbiOYkgsSL+7rRuNtvyxnjS2Uzxd/VHR1Y7EORy85rpkrI4
oK3wQ2i7RbQf7qaSN64P81tpKI6kBSea3P9n4U01snP3VQ9DHq0IjAMjAhjGl8UzI7qRw8A3ZwDe
CUiXG08w/X5EaLmhGgpaxKlEHQljbma+7yH1wS6RrLt4RmUKyWUffGS4QjlpYA3kwLhrNEiKj1V/
ty4SuAE4dUJtoZX+0tUtVhMKLjQs1Z93/CaMrY2wNuf07LWcETFrk1UqUjgVWXffkrx1ARYa3VyN
iBJnoR1i0BUtv5rZbNbLRGtP50LXaLVqkz04pxfclzdnKbcrz804tAzmfPuP1KnrbKZqiUEtsX4m
Fn2zuUS49rU3A08t3T+G5tQaw8zIzzlWIZJmtwn2kzhiHRRY/09fBLAxg3Xu42r3ilRe+Ppn3DtP
mvONANWgxgnGdED1FtiaZxJ+HDDOU7hvMjQHOrn+cOvBYkKVtYahN8lRwOh4p5P0cl19RIbVVU1I
xkKBDRQGMDWMJZ0JohG06Hu6votKH8ES+5FqvYaA/LG/l6THEE5buGK0xH+oIBH7ycfQbpqX6R1A
AANYei6pYieu3F3oNnPsYRJPfnZ5ObD/wjs1p9BD4f9AUeGvbG21B0677neQ0t1BbXnGHB32hPvw
jnMKqxtO5JpyRBHkUoW9DT2ovLDRjEaHRBCvctNQQ32H53cS4W4dQ7izs55ioiL2Elg+1Tt0YF28
Sseuzc9XDGn/Kk+nd0k54ylI9bm2ZuaBpxAZrOk+1bolhTS/am/V5zI+84sWkv/Qw/BfLbYWrNRo
LVoQaVSPyvbQUV6zG8ci/fq7+HcdepyoqarHJbgFMHIT745wktdq5JeGBBgZYAVC/fX2LBZAnSD5
jGRR8pZ9/onIGsydTOluDn6/Swfzbxf9GgacgLa720Z65hUzVAOq4V3dXyedqdk5I29G1uuU+hZc
niYKzj54mKL++G0RUrKq064uz5kEgbHsS85cwGIMqyjMv/8SyAuA3cOSpvR4IHP99ihmb/tL+/9K
z0eNHMnaLBS7V+K0yd0heb6dS8EZ+eqTcWnTPLatN4blbpzk2yuc5G5cASWuxRO57x1hrPOaxjt9
Dtw17to1U4SqiFRbVnAAITnFvMqZrD2oc/A5usvznPxTwTqEnfD7HXmXUKaNmwBq2TAfH+3T5CT7
0IEa2wlkKh5TVQubMLwT7Rupe/SrW24sZCoM4V4wJp5/lY1pkgyWn8lZcZWribVOLnZ7uwuCMIz4
3gzJify/9lQ7hypkZu87HwlCGN1xEB9KpEceSiGSad+DNIsFP5+szpGwCmUbWMZInrFcA9YwzJu+
1wKyjqqobuhDFk3D0n2u9VdfyWm+TP97Xh45qWKxCBhSrdSs8l/x5Kj9Zp26yw/jihFMEn1+m7BC
WbT56MoWXcSA/bCh0Bw3v/9aZfUujQECZLLBZVX0mJ/twFTbOHg27OLx0sd5OFk6t972Qlp1sU1z
FL3aV9zqJDRyZZcvGl56X0yyrV9F89F86SZgTtxivxE1ijR+j69AeSVOVKeAR3YP+QYsHR0aiyjD
3BlVI8xzSMt8vOGChEAwUaCIuh2tjtM8Zy6To/70h5KmN0vASjcctrTjht4A7VCxA6WlzDZ2Z8yw
2pK9BgWrWfIogiqFcz1gkfTdWukgkJ6h4wZGmEkeD9UkEdzR7PSU6ll7YuDfSIOTO3PiqyPHgebi
W9IqkgjVwL2Gss1VDqC80gtTz4E6JGOGPE438l8ntES+TZuyaEkips8jR9JVGIzylXio7/1puKIp
7q9FUVHQAuHO079GVZmKsfiNBcrkBIv/M2Jy6gIWzOIFIM5MWt4Slz2NFMhtcxR0TH9NnNRf+ZDy
QOz18vfsRniAwoz9mdpg2OP11rzQEsiaZVasuaVPfmYUpl2FfFaUbAtgj+A5x1eJJIY1nwJJGb9g
7InYD8ToLpOF8HGkE16pr2ed3GIcPVHPDpsdmfFgQsm2S5GbW3sfXEpvn9yzICtn8GLxIaVQmibZ
1AgD8nATQbbBNiGL9Dyc0cxeAVVASS5X52Zx2ckSORXWoQ1CfFth/iuQUqdrqFxod797fWMl3byk
EuMIgsy9uOzWA/TrqNEjYRfRjgWIqnRI56sGCccLqSmLSTR4zhqYsFcdAVOGFjEqThogmFDCWJgc
GEqLjbXXv1ptTLNbqqE3hfoRs6UQCdxuPRch4lZ007LYcBHd1p7dcvSSeceyBLqlOGafl51nMdSU
h+rHRqaqaol1FNmflEzXTOZwxc2M7RUMqj9h5UY+H7Bz84LrDQBcebnQbsunVeBcwZdNK0ci22wA
p+LJVXmluC+0w38KecYF2H8RhbnWIQpggDlEmlqP8yW8Xbrrq7754XrfHA4PHPDjrc6tOIhkzxsB
PIMZwfiKXaywZqcLosiRqu/Gd7jdVlzF9GVgovZDBNIbw46nJWYzkiBqZN7kgiVAd2HmcEABONV0
6HUU2iY4rjGezqMdLbblcdJLACP5wtsAirA9NjuWfhPeSVyRYrhEBryqZbQagxuUKdO7kwlTY02s
O4BLb1OYTo+vMzc3QO+nEW1Wc30ViVcJPRtGG/zxdtSZC4ImF9xHOtslrV3gXPGLYVzNYEShcWAn
g2d0e+BbAsUWOEaWtEkb0keMx4DhC44o+O4OsvQ5JpYn2/Ho3M+wtNZ0wNWqyWPJxh3AFKZo4jmZ
UimJ+LXsQ9kqlnmfMtnapA/l9W6c+Zr6qoOKMyNayseAyDefWgyRaesM7gOQB5gzgpZUgd/XSOSv
VE63PBjcDEOp2QVm1pXwTSSR1G0KH8wMbi3fwlIvrNSLcuhHTDpyqvKTiv2F4pwoEI84xzS9tibX
zv00MS56OIW+E53nlbH889uKmTMANjvesQuWcQ9xFz7wNbcWQIDFQlZxxASEwCgp+GlII3oCBsR9
e/z2E99TFdCKS1nvP1TR5uPrCLe0WGSvSA7S5DP/ztlPAWgrwGPrj+5eD+9dv7rbVVtA2cDyS2Sx
vdb9dTlaAMmyBUD8LrVdt/S6WnE8goEmpf/FSR+A91MDTngCMfVCg3sbKsJ78c+lO/Nh6eBxDigY
GRp1Wa2bwieYn0QHydqpk4bidveXEAPvHFsoKvXnWN0d7n7h0M3oWpgNaziM4xx/ZdgMnw4imkkL
UkatOGx4uYe32dsBZ+woexk3HZCQcuLzShIXTP9VRSP1PuoOBEq2Nf+FeyJQfFXghG+mEb9chsd7
BtgxG3698FAtfh08D7yz25bS8r9GfgOUpX3mjVuGf5dv4hC3Pv66i1HSCbZDHlRVUD/APTBBQi0X
kqy62d6ufCdxrzwLwVAQReevwSiRIKVjABk4LIyXYjZn0HM0klQ9NZyMHntA6lQORRUu7QOAB9Uj
gNj13ShNXkIDaywX3kAxrejVHsjUuiRVJUQ2tr/38P+V2HRTyFELU76E8m1HRiU+NB2aXhcb77Iy
sG2mKFaEINLCnuAhO27c6U4T5e/gmZFeenr/VIYuh8GlwLicNwOynlV0ka98+EZ4eb5FEOEBCnu9
2IImQqTosanksqwMEVz7jllvjkTX/cmwcXw6DuBNscbCCAc/eZfR27JeM9E87FaKn6bgh+co1kAn
DjMFF/Mr0jap4RnarM2ak1PzghJRThGxqxHoDNrkKPgtZ3vNCgOvzsGRTEgtqGIaMFa/XC+SNqFx
O1P2GPFApOvquMp2FLElP021M5HYJZw4uL3pXGmOV1Z6JaF2186sI0H8+cqb2NTLi676axdOGR6m
UtEbG9b4GhQtoKDLnc650oQapHCpDexbZn0r0VH1bM1TMAcfE+uSqRy6hQTsARIBPwyXPJ/0A5mo
X9Ddu6t5J5X0LcAI3NhpEX0TGEN9S4FFbIhR+ZOTxbIQQ10QASt2F48AK2ZoErjJQOtn6jR48dzt
1dZbpS93mzSqpnnzJ/i5S92Ki8DBOkQLjlQEXy/YoC46/918houKyjTQ9VIEFRaA1aDYWIwmi4er
zck/+ctNO3/xaqXRXOtYmjfItGefXfh/Uox+P4oognyQUiz/zx5BWEMwfCEJPDOnAYWb/APozJpB
YoVynUUMBUTA4V9a0qeaecDKpImudwwV2qTtMQnqU/P7xF98xUrsZN70++Z3w5n2NKKIcONdlD2U
OTINDxP4mwvh31oj1i1ZPj8xWnd+kNWMDbydDmDsQxx0x1iX+xT2rbVpoK34W1S1VugQMyx1lMno
owz66JzL0qCDotslSUHzhs5FMTgEmbrOfU0agUZx+Aouk15r5w2lQ7M9YastYDLEJpnInr+P+BMf
4FLSvL6td6Iswt6qAoz0ogRnD+jBz7YiYqfBNN7sqYPwcuWrE3pAqXV0gd0gJN+LAN7kXFJnFQ6w
P0JlDaoqLdCFx/0auMffzXuk5qaL8ZXGHPtdC9/8Njrbd9fgc2KlZgueDblnw4U4HcSWtCjh5kCf
Z9GFkbQDS9tql7RPdG6Vt8sPbH6ZjI3DWsCZyjvv43xfOQ2UoQMvNkzbcSnTul+CpmoCdgulvHrj
NQUUgkvTGxWUpedBdYngw4pEdnbCH75WOSA6z+he3xV9M2Pw5FLIlbc7GXZkP3tzOmWAI9eFUrTp
2ENoMNvRmPi14dISKqw200BKGIF9FngUHIK5NYxlBkof+YIzmqpvFC1jfnwDX0DvKZhA/xdAOZMf
zKXkQtWK7y6xT7Pf4e2BT36PcHZEaz79P46xYCabYiXPcVt/HxMLSke4OEJU+ojLNE6Q6ve2Hgzr
T9/JpklJyMHnJFaWBbKJ04rlSp38WNYVE8/nxLQo/mtJBdoHEmIOpy/loLMxeor8ajffsj0PU5U3
gytDo5ADI7XqvS9EFg+cHqgDGSZHGlAg+WmNoQIde34rzi5paWdDo0HVLkfv9v3yMd75IgWfgmsL
eiOLFremWlzZ1y6gfiNgVj2Q6wvnA5VZ5Y630PWoaYjCDozd/DfmoA/KwDWYWI/d7K3dR0ACGqSG
7klh/88/Lvm4zt7LQBUCHItQkutLhn4JH0PtKtFybHTWrnUBEri32KLaJ/g3oXzrkWYhvDJ7d7Y2
t+os1K2276Hw/ApW9iaqYeKCY02iwINLJRJemaGEWnGgHwozFnrW2KP4hgpKHohy3UFAoWJI58kI
mLaX4xCOij5fYXyuorze0LlSKkJySK/TEXDoWOIt3jwKQOVCbxg4rJ4IX2zu1lC4i6epkV/AmZYC
VZ130SqpCDQZ/UxkOcQ1pv6xt3A+fCOSBsqLf/a2ALp6z0Qvdvr8DKZrhDjwAPlKDsN7/wZ/0JrS
ucvpgTfDEA0yAJN3M8wxNVD9ULRDcL9rJuh03GDAulFDEtKy4rNT3xYvyz/fMCTCBpMqBJSa0gCv
ALATxFEuDoTIi58usAjRuq9Dsh1JlndoZTUPD3wpNh631CLMTj/KyclcbOW0qfJohgC3PsXH3bG+
q65ZMy9bzQIVgbE18oimF0UWjppTtubrOuGf4wBP0r7Btr/yftUlPK3XyEqbTcyPWzIsjLeyE3Ge
3A+GOkYtXovq3chsHiwYPdoDQL+7kim8b2a6+AGtSRVQnNBeJE5mhJpAZ8zHcz0x5YcBx902B3DM
QI81WpA+mb5FsMIe0TbS41h3LNrTNhCPtCroe/XCAUR1/pyp3QlsTuw7laQflib11wu/LFtbHQNj
985OZH/mpsP2RLBYdB2YwW01Xhzx1UngXBU//KxEr2q+jasDN0YkX4r6Qe3xqdHEN42h6xlUNyG9
KbRjxTZy6livMSS5BQ+Wj6fSPvmOL3Jx9L+gJUgxkOrk6Fz/c48rm1rPTEsbaq1EXfaMdsSbac/w
/kld925MkFC+M1mMqEXDu0STOqMvYL7IcVZuEa0vfyEyIOZ2xwbNETdpWQqARnkUxF1vcJh+fzXk
uStKKumSdfbx1l01RYAImNvRz1K6OtKnQxNDjsRgoaf97jmp/gMcC0x+nJjQXPpTqwOxX1Y0M51J
R2Ywr5Ai9Nlsn292CiF4/BK9tZnYaZxMRAx3mL10IMOJc12p/eNGz9kNVwzMQ8ibhrIVbfBhnGNa
JemvnO9BFfnAnfwAX6E7+GXEM+Ta6ip890sBAOCJqrdRBjgTNkGlJ9UDXf4wN+FzZZ9Id6yk1mCp
2+TGEpKVb/kzShgfGm4uSB7E0xKf/SWqL7eMpdgaL3zpKv5T01N/DUnOijUtDjeLo2PDvJrtYBfO
6ycuRKc3+U857sFLCh8Db3749vJSUZz5qDXDaiIMiIiWmKlQL1TySNUKLvC1so42/O9LpavI+N2j
v+6NXwsWmdWF67qtiXJS0s7J8LncPz1hFZ09Ki8jiuPBSkpuBWLK3TTXmKnydKopoI+jYSeHHdhn
6e67OzSWfA4ftYIrEccuiEg+/Ei4kHos/NnRM6Pcg0RumBdjGgNjtHwckgleLw9DHqQapWkqtvzD
OjXqEcTrr/v4NCfwWWRbMcLDf8Ah2pOPaEIbgCmnQHOELP7s5kF/oJ9p9PTR8ks7g+AoU+glMQhV
zVNN1JJde79735V4lETTVcL2mK5s3MJVyQSP0P91iOmGBaSXa4J+shfKDcUgESND7vuiRn499L3l
+o2Xst+FrqssLywh4yVQPuGgAWTN8bJ76o/PcBwWHCo00SGvyFVhN8PpflGSdaoWRUjOwVjLk8Jq
izd0/FfX86s4RRbCtyC/E4S0keMKsvldNWmzPky7Cvb2vLZluOkj6VxGI6JkIWVHd/WwL6pvSVQ+
1piUS4GI7OyNn1tlFhr8v650Dpk5J0OZXqTX7ra3v/cLKqUpX+08jOuUgVHGLBQg0qVy7Mx0ALI4
FtVmBqJHV78ye/jSVqlb+toEFBmmrNmgGVho+0sTEtXj7RYnQknEnhp8GdKtTHhlQLvaZqgylQI/
BqWyKG2vy9Y2UaWE83840hFQ/2+tws2+isgJ9xe5E4idhzhNk81EqvdGAZK/rZAa3hPWynzYcP62
QQHyL8whNMHuIg3ADR4HancTk1KZu0VJejNX4l4Z4dD2HOBmPg51iD2P/Ao7hv0UJcceMVrWW6mt
2ScPxuMg8hUu/SU+ZwHucPxB350U3vbZC1dHo5I+YeQeauJ+d6eiDCK2CXreXw94UYxkNg9HtsBC
WveUx3ssqdS0eFRESOc1Jo5IEHgHS35wg0y7skV5tdaTD2vR3cQkzoaw7m2HhC0gOPSV2oypkBo4
fAT/vkzLJ+iqvXpIAGzDDGePy+9rTXRVDJBE1aaXJXRiw/8Bu98k13W7h2ov2G4fKxZSj1tg2fdK
Q0obueduH8gmf/PfpsyuSxtt4KALWk0adlY6oA40kS5ssrAsGCDJnQZo/N46TFUNivy3a7iCKyXE
OqJhdtagYZP55LD/V5GUuKjlrFGJWyo3sVNNKijw6V0jmQx5w6rwQRbTjp/PEuY0wsH/aYadr/dM
sofyZA6vQR55V7OOsoVh/Cb48hEhXQLXlhCgaldpJgKtmqjMiplchvJTTDhhZl3a0XnnEkIQFEt8
0GmOlJNvC6yemNgDmLIfzMq6uMLlKNV6HP8HDM8y/0tCDB93I6opH0rQ4Nzd1hVu00J/AQybRsUa
H81yfgpSKO2mvpla2dzrGmd4S+RrJOPpks5UcaFOG8g97KPW8HPUra1spJSxAMMBPdjAOq/j3HK2
zst4mGk3LTxf8kYcbhuTpvip7NUn1Mv1xJXebPmdAXQS2qFzl9RDPzeCh7BTEg+b6VmOfRRgPI1p
ctnG8fgBC5P6vqskud1Yif1us/PHR2dmjS+b3C8r8stZ+gQZ5pRY/g34eaLpk7rlblC+In5BFp8P
D+ZAHw2hrzFN52aoEnaXy6DM4LOPdNOv7EXWIz7Gbose4j9Trhv5gHWGqjHj4HUOrrJZOaarcJ7l
Eg2x9m1WCJxX89sBHCC9ZVJo0rLNRa4qza+/U2wYb9Z0Jdwv+pnf1H0UOJUQyhXhwdJUAlgZx4d6
Z/Uj4Ya1uiZ+++MswOZvcO8kmuQXL3Zj7mzxgzpEOrxeDijfkMNSNzzfFIz38JB7KsFBZprU72M2
vZhWHGyjrQgdxGevqPC+nxnqtD6aSafHiXSZODx7PWAUJsMUkXDnsgu13Li4U81jdDwvXwr0YGz4
cVXj0f8ZzINgJJVb2dX7s9oibhbE7LLfCgrS5VbhoBgH0m9KFto/7EWTd0OxVT58TGyE1g3RKKfn
t9bx/q7xsaxzPLk98I56xcOKh569s67S9xhylckvFOvkQNsytDgFXhJlUBoPX0WUwrSFJcHEcN3w
ZXagKCnsynErM0bLl+Q0dxK4Cd9XU0zf65+oOvK2nubCgqXe8SsEAxgYHouvTix4prNKsaTp7EC7
FNebtGfSqosDWhEd4J1oi0WRmodSxw53XKVh/MAsBzMW1qSX23M8BeDbnV24+kLTw94iOj5lyPi+
2oKn1aC2nLwRjs8IEi0MeaYxf1xEL6tCB/u/VrI+aeLqr5UVz/IWBmkPmRct8fngaefaM1jebzXE
dL809oYNZoexVOqjFhuwomM+ewu9uFkRNb7KVVxuScB387Ix/Ux5FUI+/cJnBiBQViNrO5qXNzzq
6+wFryXZAbmp2D2ggUQPvZ9U6nrX6+7xgglLvjBo0IR0rgjhtETtIGzHgYMX/ziXZOiZfv8KeRET
NfNnfW0YJvq6mjrOEOueVE4BVJ8+5FKl0PANeoyPxCJdfBpOU6B7bjItEwAf5asaIIG/c9SIWFwF
8CEqbCn4jiXEcXh52c2NgAmEoL6deSAJveGAhuQM/Og/xva2Bpa+HVFE8RX37FlfE5itldKmNTze
93KX/IovN3NBN7CH5umNPxhapRcbeIFlgqMP+YzVckWngQ/+YxaPh02legiNtILjUFyn8YEqTHAZ
/VzMUHqU5bjg0UjaHLUxx7bPlkkW8bNAq6Yd/RuKmhh0yDGxNkLtsqcRbCclVAUz6+kq21wTJzzN
KyY4nHM76qgMdcPZVqZ+mCkBBCH44s1j1t1XEKfJZe7UL5Sk/RJZd2FzyN2KdkqOSsM9hT0LXUSr
lcR8msw8J/1dMeBRBKJD5YnoIp+ZXPVGKHmngmd8cGWaHLjCXk+hUjlpnuDfq5MaN+X15ONoLD16
ThTRSdo31R6muKdT49wwloENtyLaE1zQN3fa/ToxoFr1uY686cKWiHq0OzJU6BQfudtFkJMxOiYU
9+Z2Y2I18ahiNNs5FGqbKQjMxn5sexuF5W1wW2qCVj3aR+JhQBTR4FFHk0yk29lZvq8aOyFfkiRM
67w8+9PRQW2KzU0xuqNUtuBIHmSuFTw/9q+4f2kTK3ErP713+1qdk+DMovQHNsME8lrGoQ7lYR5/
2A5+asLGMMHcxVnpOAIdqGxBLfl9pf9bow4VJlKPPpFoEdZELPDwiLUUSjAp56xxB7kGwkFneVBz
MvTSV1ekiMKjBs1QNCDORMECFAdzNMSIQSQsXPKppcWNYI41DSm0hCaj1bPcFTrm3ovMPII07O8K
0J5jPjKOb8doLHdNf8lAz1MxWVmlbdxotK4MEYtUXlOdNEEWZKjeEDpEg+7+EUgJXKU+YrAwDdsJ
SNIu++wmQYrcAG12zRWy9x6iL7HKOMwBae1+YHNbU/rjO8gL29H5mUOwQXbkZHUTeZo7/LygTUs0
eDxqaaOIs9YzRKBT2O9OcQVbcQoK80CRY8yii+vkZR/7LGgUtBiOqe/T94zxyMqCpM4KO82AYSP0
Ue4sxOE9MADT+gdzCt1y8i+zfZA/3PcdpglHB8klNtzH7E8TOS100c/zjYrSXF7Af22RtQuIHG99
3cuJ1IQ5pWkp70leZOmDPOSDfKGOJoXR+JOJ4t7QdlG2KFaQf6+FU/ty+xoJPJWBM58X99Px3sxz
sL64p+WThfm0Jyg13urOkztpjNh+qYilVLPrZ6CsOZwbyddxL5rWC3G1wPxmoOd5yeHa6mVCNSbc
noYz3XUFAOKJY8tLWgUbFwO85h/DNx9JKE5qxkeqiEVTzwPZrbqoEx40bUXhSpyAktwOoAUNl1Xk
46MkT+LHQiSnSVNA3CWIm8zPPQcmgbu2PLOnYs1+d5TUAvSNtCyr9Va1CK0wC2n4fDlar+ETtKge
FMxcaYmoJgjX1eUx6BwSbYicNu1PqSxEscc30wBmv/MsLFwtY0CG8d5PLjTzlr7EcJRS2HK5/1NX
UensBIZ9RWKknL2dMT9yeuzyf81BzM+i6wWWRZdFeXamWn/YQqeyb4jwagupRvV9a5oX6A/KrcRg
JncfUofqtDrQ1I8VEHborJqAXtlwauDrQsb0o/0LsKsOEkE4b4+VObHzNRKf4wjTHWJA1HhhrLAg
H1Iq2Zd3WerXJbVKYbb0tkwrBYE5b7+ICPPP4agKiKtgLJ5FC0fXl5gtjkxaMKRMBcSb3H+8HY5j
V4ObvldCnSrq5bJccoB93ZlvKCfdUi+o+a0E92uS6c+xBZU5rHlEIWIDEXY9sETfTr21jfAjjQ1f
2zkP7aX92ZXYFL8w6smFie/44aenxbKFQJjt3ujXVCCFjPI8zfV/hPHzjagu9UJLH+7s4H32UeXZ
C/5l1HlENr4L0j98ZCoiZg2Wkk8Kpy/NgIPi9Wq/SG9RW1+tAvnycpoAyJ2o9Q5nxo408zJSpfnI
4M9pW+sSFPrrsIkcHzQw3b9uR1RSBfw42MX794rHKy/ngk9B20IVFgApNHlIlnlyQnPlXnQ5ujqV
YJrfsOJi5SIzdcGr09d/5CV256upm5Ne4FELnGkIq3HDdflQ1kTtMKsO3UX0rtKAbc9PpRekN/bq
Eq3QjmpX2KtGY+JD9NHyCHPTrcJJMFv0PMI0waNjKLcrDrGwE/uITPhgEcB9q6a8LXI3P7jsmCnp
KutOLwJO8tOnrdp/+8/hRYNE9+icDWan2Zub1pb1jPDCh9cG1+E+ZTzC6DK8m88nniMqasSFCzBK
YvBtlKzr28EVBn8Z2BbxxJHuCKics2CsVhiI0DYYAA6yAbHqZ+M2EwbsYWuotSZ9rUwEmKTBIKnN
LjB/vI6BK0Aj8G0mmHClTUDWR1RpeS8Jn52qNSGCiKIIS8VHzHtatgkhonMquLBC0+Z2EPnMH3qn
4/Gbv1gy4fHoE+oZTk5T/i8n7nWt9StEXgbm3pyUATZhfnc9nUweShgBIrIkkrNl0uPtuwg3lueR
oNodCJWNYiT7LGGBZ+jU/kyTV6bzvja0IfSh4XqyM1TGQclZe1Qz1rqoFCzFakkjMjTyYwIcWiEO
mFYKN5xsjs54xHyVdOUv1NOOHZi4XgbpESM0CmJHReq+KJQ+i0ArHENCiwFtaUQko7NQ/zUsA3w3
fc9V/fvSReUbeB18MBTVdd2HYcd1Gt9Sx75sLE+kiMBXI6rslo8JAO69fEIqj+SVlPIsvvHHKKCU
a/l4JdMt+kqNaAoh1xhVd76J6ja3xxIwoFxClDoMg54zPOuRpuG1O1ESnOIPQZfsh2whysiOpn5l
BaFMNYPB5R4zRix1C73qj+wPzz1OIGSjCaLC6jbcOKIzlVQUoGQ4ZeyIGpZyF1t2Q03oxHSzQTRj
t1BjKb4KXx73lBCAk0EuVtpes5K2TdNn5k/+vn3Zl2BgI8ut7Zq8RTlbfU92ouEEF1OIlUr3KkAI
OxYgnlpNKKq4PN0e3Y+fSZCai5ZsnknhF5sWpP7u1jaGgU2l4TPyiVigCzIZgcqcLbyKqJrvIPs5
dK/Xyi/7OWICqckhBaiybNUW5nDrEVjoF4eaUOo8Lf3xyLbNC3D+QD5HJ/3XRuaeimE3Nom3HIO0
QKR0jP51/zC/h4QW0nDn+DIKEzeUP34RrjfwFG/4tY2GMVmGTdngRU0vX6Fmt6SaFzF1u6kJuegF
K0DBvrXtRmRkoTae1aFcAfLzWKHYiprpKKN4/oUYIVwCHvM2F1R8DuFet6j5BRHQg2Q/CWRpzxfn
ZLl+EZStduoPsUUSh/m0LXNwmiY82WPj/TK76z1U+arvdIDDh4BVT70G6Pl9h1ei6Ytf9SjzW7NY
kCSbqWwHMqP2JxahlRf6ellWoXBKbU/+DrHCkLkJTo9KqrZSoJ+ENLn9HFbadQHUw6gS3vSGMWe1
CAnMcGqfTD3jgFvd9tE1TdC+9oyaLE8HwlVIckNJ6gwl1lUH2htu0f55w5SV5FveK3brz/Wx1bMn
BbXk8hQ4v9oPNx2HlhIhZ/+L+/Kne+sQraR+X2OmjuH7RKtk/GiL5jDD82SZoeyZshtly2AEbtV5
bT+gqJ9xZX2XVFndrm8pWzry+OP0AmSD24th2oCQr1fPVP+iXScQfLi5+kAs38SfRoHqqhf4h68z
lPiMgJ4U/9ASJ8v2UK9ajJ3PVftnqF4d4w/eXdzFIzEUdyezpQ1dXs5ThHhIYnCYlf02HugFsQjW
o9TH/tozyhVcrUdQRN9+lWOHp7I8j/Z0KVQUysccwHP7kMtWkoGapHnDAc/7h9wwtfKBnV0AZVf8
Y6n06Ks+35mY/Y7z5qp2ARBA0Eo/PrWdZO1beoqZ071BqG4DjdXJ4pxO7lOy4+FesIvurQYNyfAC
n9TR8srxOhOchS8pyDTCouZscbBnul4bFq10VelXStMm4qAQE0Poz38VRXPr+H2YFMI5gL9swjxZ
CiN90g3vY5vIvIEvac3HJPaOZtwK7CADhYb82gNEJy4dxpFpW2170b+dLi4CcVWBfWj4dtykSXfo
JV6ZO16yh1v4iV4LiubUnoU4m2HvzAtkAJgPnJH/qGuEhT//yKtj3uYHVOOOtY+C3sHWm8VeccfF
s++Ngqkr+YAFbMqZwR0e5BWvk1ljp5oZBK31BEPCv9tD1z57ZgrcAFdvvEIJqy7C6E6Mqn2Z4FUm
O1rdI4asPhzzvNtuAq9CSAnBBFCMD9RUkiJ3PIBvapWLPd+KrxKtPY+9oy/c61N9DDrDw2P4qCH6
L3gZfp+ssD4XOWABGH+txsPRoup3wzAY2+KLRARC85MKIV+37DNl4ErExRJ/qWr9ccC6+MNI9SJb
RR1UPfS/jbgNFN4JO6mgZ4t87ij0paRs7sRH5spVh3v3pbUaNwt13BAgE0W7WHsOJ3BtwGody9kI
QTGdMlfz93JiUxsInzRM7VAW4uh4sibX8jmuwYQAK6hApl1TBBZhKgyx8m55NElPbz0ThBoL7VNd
4vpF4fYNuDDpguaWhIz5ZOKP+RPqg+bbSSA95nB4HYGdlV7ZvZy77kH+Sf9Iru7lKRVM5mqer7A+
dIb5o+avpHtIkxtmZK0wJeriK5hiRz87Yv3yu0C6E5ye2ztv7AG/q8mcTxgyXIc6fgRVJEBu8sH1
aSdYZ9x8WJilQvl5N2zYLO81o1Z0ArNDhghIQ+rXCkWJS+s5X+E4zDtpjuu1RIbNuXYZwnzX0jlF
8N5ACGAlzHnie392HF/iGvkU5oC/SnjY29a31uRcLSYBiTT2SmocjDhPd80S+O0ofar4MHU1YRfy
RDblBo80XZmb0a2Qq34LKjgtdzot6IfgayIPDHf9S1G0+3ZR+XRm4s8dBElikpJ0h8DCUGEDbfEH
1jlAmyyn435/brmCBBc3z5xzW1oHO/w+wDCXc+nAVO6p3k58kr9q80Pixr11vBjGWKlWE/01rkyM
FwNt5Y+vPwnCTAl40ql+2esvsaIhKa2Zwzh6A5thQD3a7S3R8vW3lntwAYobREGESXhNzIdMEZ0i
k7fzKZnkk1o1GeGAZpOvM9jwz7DSFLG2sDc/ySWHYWdkD6KvgM2rdL9axtZc6TM67/xIftGyA+In
C9onjosnLQFbb+eWSyCvFBfm9UdD18zCPn7rGBqycvwGuohJDrdlQPW19Kk2NZRVgf0FYv5hA2d/
+9ng3eWw9IXT7XNveQjL3kUbGk0e7d+iGauyZZjfoX/o0Wf6hMVgyDhdAyV8eARcKrlGIFDnSkeE
vsVTvY8NKlzRXSs8ahDnR2qapm+XCtQ2EGKaNpv4Mu2qZpGcASWL+ub0X4IrsqLr/tZub1lldkrd
af1GeaI50EAqxr9wbi7pi14oMEBhcNSQF1vCRzm/C72EWXauKfNyLmYfhjLIpR4RlS6pWAHjQbzq
CCorasedgPH5bmsLLfh618SSngNZxGnLnbJruadyF5VXaaKIUpWtZlV8iudb3jQJkapaEvDQSkpT
qv8JuudpYDHriz9KgaupeNV7CpC4B645lDpn1vQbSy1XFIBcZiTLtRn3GqUczBE2z9Uv58/9IQ0X
TmI6ry3l+FwqCI7pG+eCEoUUIxK5qCa+STbc1mcduherChdqqbwdGD6ajHPsAjO53zu6GE8J0nm+
/NtKL9qIbj1ZtKzaqQiWely4Jt86byJrAB+QvEEYF3B3OOgS2EOdIDHTf7iWfU/ZKOLbuP5VnG6D
WUnsmGqpixeW+WLEUbshV1UX6Q146XLWZbb4R6I7/fufEIKnIM2Nnc0x23OLXFIt8BuQrdU/5T78
2H2pCbyI4jOf0qQH53DLFc3vBDksMCxLuWschhTz/hUhxJV6Kj/DYigO6QCowUDxf89SPXlN4Mj8
U9npOH/6+BkFxskr8pxzyDMWdrh0jSdkpOh4kmITjtw/Y4aIaltcWdqyycHmLsz5/NFCIZAyx0OO
GDL89YefipJ0RoZ7/85SmlPlKR1PMYJ50yKTwg82lao74b9I/+wzPvOiiMhXnBrDvzJeapUUMoCo
cOCqPrDbksy4xzFcMBLK+MktkfGjb77emyMX+Eidz/2knTYlTeDjESu8rfi/5VY4kOAUSiELPWOu
4JcE6ch2oWY0JxJANZrbhj6yvBsvYqz7aMXmeqYKD5RB7uEK3K1Sg2/wmAq20vEeN76C/d9RuEeS
OFrgEUM4EZ+CthSTcB0c2KGPnpiJrDJsQXrKmosmdELOILi72LRYbNKmaeEu76lqlgb35Ncd+Zd2
5hDTG7GKeIgUuXSscDniIJxPGc6qnfFNizg+wYaUgrKqkfdVaHRANrvpl8E29gzzHdqhw6PeCxdn
5IdgiVervS9R+jR1385Zw8LnWneCquofonNpKmYGFoVB41ylYFAlZDFSLhSMQXqE0NnI8ovxXlvW
95prgQb52V6Bq+XiWzuApcIciSgJCT4FZqkjQlKPcW5ll6ajyX9pfwxfrvWKBilVyLi7MBBQ2LfU
Os1O7qVTnZiyYiwAdCQxzGzZYSRm4j/FEFYCPKdgYE/zY9iOyJwA3ndwyVsQ8Z0/DnmnuOqQRfMC
W4BikCCqz3vY1rwZMMeKeWry8txE3wrHJlJBDKpLXLktgK98v+QtMGKQh0ei4ntQL/Xr+4aAWN1q
ukfM91rrkidaNzuiqQDocgUTZwMoo/bZAT2QIAU3mKHvGltZIlFDOEnjbFovejkBsfvzyrnDkBYo
5vZ4bmyh1L+joQZW7g1KMxucRPVXiV4M8iDW2cNRGfYahNsiLoYUMhxEasb+i3H5yPCQWybnRca3
lS1Hd87NlUIxAq4ow3XPBAtird5SeLwSQQRc45DfSZunCtP1G7ddx2283L/V6e3Rd73KOhLQufCM
dvOWnSOYCWMcHQ6qIDYWU2M0vQLZcbjbHvjXHXuCSmM91bK3PQlVLfOTZ5qSXYf0zr/iJ07TMC8k
00mcPlsSbKGbYcGIIqC1YVpKfYu6oTU8KuCECt4sixfQL7x3HazcJgIL3YZDtXwUHaINVyfVrMgp
inIXQ4xnfuo/lb1tkjHk7Hic+YVYCESiaMqyC425xNiwK5lT1mTz8MwxJz2dMSE9dg96v1rYUQB+
MG6rAGqymwwlwjSimtzxjH3pGEQJW/ZVl3Gf/KWZq9pKrPjradn0TC/N2f1jYxqhLXoL9gYCwv/L
RSf+rfradIMk3KvnPm/7EfZq3hxZMadWXbh/9PcLVE7c9ZPwLffaZSd0WDMOXPaxSdhQuxG8H4nd
gUUKjS8I5E5ms4SafwWBCtn4wacBHWYEZ75iiiCXIBlZo0kWHtohURsN+42MOr0NA9ikKkNTN6Sw
B6ycYmDhvkLsZxAylLAnrW3YzxwBKOO2QC6Sa655lGCxeryN9loWOmmEJX/fulLc4QAgOuafvK+o
/IojHNZrpMFxdseS9tlgdYum0qIFKrGDGnTp5ES99WSML/8txyPSZotu6mz7nv5lb6zboEgC4LdM
jzInEjGPEe+mhzeGIi4a8rSFTyNLZkxyb31CmSAFa4vIXoupT5pICfrwxr6Qe0gSxpzVbEdkXYkS
gho1DpTx2Ds85HEAb8mcYXdT25TzWTOWEgzKsDlcQkxYfzQHh+m1WBHgOwtjZWYL8JfjeU0ek+Qj
y7Pb/skoNy4keLXL/sT+qbWjC6EVZI/Rd8x4bmk0TEidO7LDyoFIch/gqxVjYXgHuw/QCH4EXJcC
nZfjQXUuZBcU9pi1gpPfIrmeT54TRvCjDc0S3HUQsdEMMVclOCAaaw5v0qrfqETgGxZmSJmvZBWx
vwapulwEZJ7QnLadz9XzMZH2VgOFJmvX/X5XhskLgkOZngcLsFIth+bHgOYVcjh5IZGRmlLAgFI7
FE78Q8AMKDbdqeVB+n027bzWeH5oWLDcTyTcmhjwqbtxFJ6hwSn/YGwMpEE/n3AMkIr1eYTDBxqM
IS6DGlawCzgstOFs8hwLOBB+I47yQ1TfTAGTBEuSO+LLOsL4l3UdggcvyMQQ4bM7Nit9xXPDmaRV
4SoYO+fIspmBHdLwlihWSp9oYZqUmmobDa//Anxd2AUm5xitr1P8dXQwWkAyB8tQn7L/2IBEqKCi
I4wYW6UwuHNaGo9+elTNgigPqjrFCtbzlOHgnGrA3ytM+Ewgrg0yKcMUUkoDfwqHCP9KzjY1isbm
56cEcCWvI3Qcgb3bmxjJIdrgMiVKZbLtvpBe6TQV3NPrvxl99t3lmGbZiFRc2TczgLURrpdUbE11
/u/nV0VZAYQlIY22IO5S2fhGtDQ1GGnkrW6Lt33VP+JV1AkT/2NnCnY6pWdm4r8Qe5LHKgK0/71i
0xKr5zT2ty68ZWaRkYWtZTJ+q55hH828FIAVlq5B5zwzdJBqad3fS7aA+3e4/3p2n+N3V/XoWE2D
+urY//HHaC8Xv/8kJ9/HJgN5t+gNCneQkx1aAYGc6YTd6t0AhYWeNnWQoIXj8FQ6h21wrQ9DgMQj
ID6hwZodkbDNUYLqjVTvVHCtWykyvKmz75L6eVaH7IeyZgZTX/v3QaqsmFCMeERGAUekRiEhQXqH
4/jW7daJwwEgnyXTatSSoDW0YXnXKqho95KoeuW/3GWkbiZsY5Ekll21cDQ9PPzsigntWqPvMx1B
kfAtZAc/yt/pZrhfhKFJHHgENbHBZwguRIQsulodM+JE9Jw+usQl7TDWkz7FTkyJfsYoBbGmbAX4
A5VZ7gDlj70EdAVUQSL+g24KW4ZIwNfFgp/yn6GMrJHD/aO4R6RFZ+2kMJAWHTym3+5mskjNnlb7
rdsJEEjaKDrtrwUdKAqd11LDPK6e2AqY4E9T3p0EpFHlXnHHedscR4i/uTqSdVxxmsX79Ge71y0e
knPfBYhE0H9akY0A+eN+hX5Bd0FC8/11cLlGyxmPg9CvBNBzxyl3O9gApaA7q0IjZH4i3k/LQvTQ
HmkNCuunsX96GMh8zTu5ObdhZScQcXw/3IUtuqnE/tFhwBnJqPXRZab7pcIFLDRusC2KDEGkovZL
pMVg8WOe0sBEt5+PiB4iyHhujN/yRHt4SBAL1wOmqLSrEogiiuFFY9GO9fRlzXNDw0WnRBldGBU2
kqxbY37D9eKdm2ONKjMEB9PFAHHFc+WrJdtVgKfQF4PT1V4ueQymKEIbDXbTVoVoEGn9iv4RfQv1
R3721fuTm18Hvg5RdJUoCRm82HYsIr+JLqmfOTzDLl55YYtdrqryF94LiwtKMBBUuHQexnKzMLOH
WJPZrTTV33RqY3mXxqr9vexnmZYNKm41pdfEI8VGBiFXlL4E9399NH4R7RDhD7YfuPFJCR6Fjluj
Gdmd94Zw1A43T5GYYObz/aKXtiXCOYp3yqBc5vduDF7AP+/nT1Di6n3es8T4dMV0ToEebUdf5lO4
mOB5T+17Ft/Fe+XDbcERdEo9u5k7/0A4wjtnS5oboY6AkSb/piFE5YgSsFpn8TgtEygA7PQfN/ol
VpKqAyZyoRMMcsA/ygr+wjd7+g4KIZfWGhrk5kHLvwolKM8UWRqS03gZFMLcEIlZoyPwC26Kh9c9
uaOaMUyIy4jL/RtqIfZDBOm0cFrdcp7ZsnPx5dJjg5CxFNTHY2bGYgdGb8yr3TJVLvGTFsXocUVC
IMximXwAYb43UuHnNdF+8D1kklsUYjNBPMe1hLTgdfjtmkL4RTFnJgKquSgurkKrwgkBRLc2RLni
IAr0UPEFwdn91rN77MrsU7KqBC/tSKJ4auTfNULHRuj61N7q1nMl6dJhT/iud+Zk/gPvya8Iui3l
Yi9jVQfZWnfXo2z+2w4w+eRCt8W5le5rP22+yBHtYal8UF7Gr5qRBr5nnfmn7I9UVqG5ig+waRAA
WcDMcgC3SlzKAazuJg6G+0ZtrApL1YKeYyGULbhKYmRaStTtVf4uLhgSZ0xCGEpvaDGRKLWLrnhv
YadHNwdNXHLXgPQISoTqTq9lQgtoH44jvnAOFU+msJL9FUpkSfWa43N4lGydSrzXjDQAMePzNe2G
S9StK0GsLGJ075YCEh6Hr3IumWtm+t38XA7Y+Cpx0B6oQnsgvMK7CVF90t7XAjV8XH8N3/ri5JDN
19yNWNQjyVJmhqzPOJNRmwJDrOBpA/e5sElYhtjHMpvFm2pY+5gxqlBjJlKM+Cf6Fw5ujvdlGKv2
2R4wft9j4mtKs7e1l6pXAtrazR8LE4zkRICrxbG/AO8dCBCudCt91XJCteEr8o+pkzbdn6L0rFss
jM32PL/KvBssLA9kOn8tm6jPNEa366xAGpslUIliKlFpMKcwEt62hUNJ1Fgb/Hkkj4hxFQdbcwy7
wNaLVUIXzUmp0n/mLnJ0GplQ0g6VdV1Z+5u519Wh6fpJP5CrxfRSd7D24tdAVaFCM/GDfzlQnuwg
N8CEMysSUfw0Ec2aZ8my5OR6jC48pNoUw2Ml5c7+n7DF0NEOzUc6Wu7SxWZEpmEBFrkaJJMMmHBI
sRd8utd/YH5bzqCwcxSFppb6C7+Nf6+N78U2sEqEFO7ps7zxntkbB4jwKm/gPvsoGmJlvwkNt3sN
xsvQoiXc5Gva4t3fDaBiJoxXP8XGEfM4s6PuUpGFk2wQbGLDLD09JwYER5eexUQFMMMnGjNVJp/v
zSQbIy4U2bNaZ89RyXD8Oo+1rFzKyD0UeSWUUwbjMCRlAqHENqhSeumFFQ6T11sYxWSmUdm+ks96
uY68RpIhZfbUYxjSXD252Lljz3sYJU6F9xGr/ONXL3cmlJJpwas7xdmhuuUHna1r0v5kZuROWElN
OgbsJSVeY+OIxibk7XHQfFaJauPKklyRh5zHJRzfIl2KNAJTNG0auopGaaU1FiqSJAVxktiGb73e
oB4Uapicg5AtoJblncPaTS/4LV/RfcnV46V1m2n48cqr3ymlKrBuwU5gKkwRr+zL+k4uK3+YiBgR
pVVFcDdnHZmnJNsjLvJvpDWcWesHdWFwCcFzE9Y43Utl16I3bP0O+2TwrIpCb0A9wvSGQwOxKpnD
WkJG0quJ63pljGtSHhezDPf+dZV18lUc+K/9TWHC+1ggvseMW2VUzcPF82USr5jkPVC8tMlZ+Gog
9cLsbY9lXGBQzNv+JZoBmxE1d7lNhtoJU3ZwR6+l5y2gwbxD5UEd/qOmSV+G3PeREEVKvcBstxQA
0J8KMFaaP6Y47lWzMLwfcPcDhZlg0JTwmOVJbjMDcO0Fm4k5U73WBuK3327r+uPKVoiYfPRzH7Iu
608TjDzXNYCof6PJGtJDb23zV1wZuJnBjqmfLWVv2KOH5YqfOHBlVhJIefUVfwrtgmWBrIJsvpQ6
i2PN1IPUln9qs9brQYB1sdnisoqzvvGaPbI9XOgWM4ISe68/5WZZAwjqrhuxjX+29DjFPKbaVCHp
fqaUUXI6lh/YxfCv140XnApYb0GQYj1Fw2kQ1bbpAll+3GfhZWfqzvt6S1pGt1X8MsxTV0qmQoAM
xZ5NOFFB8TggC5RnEwnXuJ6TE0hS7dJCriEm6Kf9T9dQFbec4vPBjnY8gJNrJ6ykLYVZglmv1i7G
ksV5Fmd6CLzeUUpb5VLt6BBzwRugBY1ihKBJqvsZm831Fjo/US5ATfMYl2ve1VXD13y9SKF0NtTv
pyp/W2PpGRScLY9tx+3QJSqiumqMExUzOfZ60j0kHQc8lEG5kdpAqUCSv9jD0AGJhArQ3I/G4J2S
C0cnG15/Gaerx1Spnn3fk+3SdDVtJz6+h9XjvzLJAQjnTyfAObi9b2VMi/zuuq2GN3j3arP3JCTt
AZuAZummrL4VCyIkoF9GNg4w1PPbqWBIcAFr8t3Ifunz6SJBgmEcqEpfGz+TMKc0MCGE05z7H75o
51Ua8dKde1C8HuOV0SkOp8W2nLZcjSpUP5+YZVYM72k9UxM2aRlyPQ+2YEM9WlYbEOV8CXfvnyu1
bOZ5tbOuFW57iiVphDyCxKiR1l58K82UrTEzqfDKqnUyb07aydQajnezoC1y5zV0vM3xDHqi6AiC
1QbJT/IaGWTHX8qvk6sg7/1vNk4WMv/nX05BmmW/skkC9d0fr6OUY1Soi1QqJIj+F7ncQvQcsjCQ
CerWyTk8TUdH0aTGIcLOGPxEEcDyL6cuE29xTNlQhJU7YzwkpY+9xbXmF4bAvzOB8OypwXGhfPrY
DFS4m7y9wHAWzBNCnnwiwvi1dcvbNjVr0lal9r6UWXH510n+UyifM2DUKYGSlb43n2aAGz0980zg
ISjBWrjt/5upB0uODSr/WIExi/1ZmA4gXXgaZcADveb2TmR6F1wnX9E3eaQgKJrl42eufdZTPPYv
wO51G3v5Ekq9eqECVGlDSr1DfWVK+xat12F2q6Cx4tuJK9KyR3chjg2G3IbXpjzvOlMg1iQryxHi
1T5idAndXjaxHk0NEeGPlf4bDuXi7e1J7bVt2LvENOvyxt2SNfE1u8eTg+HABd4OYW64yrNttvVV
AaaNIU30Cr+09lD79iAV0TlEE2sNsbFrXf+PoSMVyC0eBMVhyz9MVXk5fL/mJG1jQVnATwylazQM
kgpK/Prx5h0hESRAj3RoibSGwKPD1U30+lPLEsARLGHW+DcS9XDcZr660mH8J4S3HLA0saZSHzYN
w5daMtjHUfFyPT5TBTqRFSF2f+1sTHaYPK3rLHkM6KEGuO1lU0nypzQMKJ15itUzDwKheZeR2UfR
GxR9gDPQmvYXOtpD4yjLLyQxG3+A7qB4+aAkJgNpEFByDe9iUgeByBlba03OY36cOhqqdyK7tO+M
T7EB5e111CEuuUn9H2d24m8iLNmI/+8/HOle7kHW9sq+gSY3LMWZ/TG9pum86nPnXQsYU9dWAaur
En5+sRAcGplvAAJOqSX/OQvYWCJBHP/VcP942D3T0zbxHJlr5FeF69xIadSnehtZYpq6iEqbjpQA
yJMGAvRB6opcWTiO1fssqt6jLkGqaxhzsrrEyDTBP3ES+8tuqGEwu094E8KSGxKJQ9IChYArl24y
5K/e1SxpE8NElNfIZq82PFrP1mJH9QL6nAO88nTzWVFdNCzSw9nczXNaWp3W4NPvUs37dtwcFdPF
eMrR0pd3ehMfxXGNMUXrUTnFwClZkWjdIC6QZt0LHewfy3xZeWW6qcixqBFagxo/PlTjMpwBAeOp
Bc2kchF2X/pC/XlBlj3AnVZTiCm0DxNdRJrDX/Mx5aau4muUbkF0240Cy3VZn+npc3RYBIVhmKkF
rJkCcRGjv/F3wu4Q2d56Q9ffAvohjCnRfI7O/j/nhNf3J7bjI6lqmNhZ0NS/zbAcmgZDxOKBKtM3
0eNJdhqMC13CxHjc7b75CoQOTVhtWOZyV96T97KTGNY9izjQZ67Ytuaz7Zeo6LIxPPkOli8U7Tb3
Pe4kFSwQ7lgikMn9f+YKLg59UIEcl3GVmIvwGSN4g9lHYD/qCsr/ePxR7ndJdIQIsSpsC7KWmvIU
wwEgzPcMijswTkA7jRNVkPWHaKQF8j5aShJXd3c0q7cc7Fpq25gd1QpgAJPSkuqiBYLo60E7tCxy
8vwTUZ/iLp/QfSpDANmhMraTSmYX8m4N9pAWjX6C40PqI+RB09jw1N0IvxTjBo+7PrfcW51akYA9
2groPQJ1tggAuD3G7bdXJPP3BxKmhRqxk/JjRiXFoE/Tp3HcxSE4TjsuNm78My3qHTklW4VVUTXJ
wM5PSTYdG9F2BoDIh6zTnd2RHrQImyyWz48+bVky8oRjgymuDwAv1EQPXq1nt6EOTxzfk9/sxNoJ
XYPScoHHFQbWOonrVpIY+jVHSya2VGRt0hC/Yqx9DGys9AIm/5CezbnEskWG7i/SRinYpFYn+kuk
KmzrRyjAyuBDWuu1fNam8Cnyi63TsOULEpSF0nW6an3Nmiv2TOb1/owogjd5u+JoUe/L7J19/XG2
4ZUR2/7oZR0mrGkZHX2OPbyVxvHv23igi+iMi4CfL8Ap0hnfSeVH3NrzRNOmbzdnW5kRGJBKkFk1
GLNBbzuxTcqzts19ShJYpFRa8jQrfnqyz8aIKZeOZ1y1bQ8kUhkCiO54CKxNFwZ2zgo905EPxJZX
xD5Nu1YGwZhfOGuMPOUhrXOkp6O/CsGJ1tgvYzLYsLYdprXtILRp8GxxvISGPX2yE8m0Og2kCf9x
iUZF8biOqxlAEsAZ/IPYrAf7zMswISlRW8hVOsML+gqY6jJ+cIp2qTEquRNqh11nFbPkapozpYBe
qTg9uLHwrmxt8MPYjyHyrLO7Va/yXq2dkXP9xJe9lgc0ALR8ic5EtxvaFGuJ8ltyY45zkD9GndOC
QNLvAc8fjsgBZ+A9c4DoB49JrBDHniG9oyvgDhfubOi6fOB83MKPjcidOvsF6fyWc9sHF/h0VhRi
SZnq8vZMvzeFtbzjRTY8T8vJ+MZEIsd9zspQh/H1L8nQAx/3iSR35Q2PQNEykPXEM5ujrYLWkEq+
1r+I2PQqinjhp1yYsrPY37cZNmMdaUNtQldEhYD3eF2h8ee5gXgoivdmqcIyHHkfvxC+xK4cz+ol
uRKsHZy0nIg5gpAX3MV3d+8p27yYfHo3pn3DRaYyuJ/g1kw5/4LKwUWLSFPFql5sfRRlA9lNpahw
RO0w4uMiUM97YB3pvAOxTyewkwRe+dTfL9UXcaQrPf/QDyWVW0eTHzMlC3priXQ10Npu7PbD/bzg
K3/UjH1iBKCdyWnI1V7UdjlvANXWnG4+anE7B98y1zbSISNdk6fbwMmvw01762XUcTjtrtSpm5KJ
TE2rpFdjeXmWoBaOkTuY/q8xr6SheC60aO22QDSe0CrumhtV/bnooDcG7oJ3qzR8m2eQCxg99UOv
hGfNJgm9wbX8HhL/t60zOR4mqzzRZdk7/FOi3Hbo6poNiwe4PFbQp0AxBEZUGDE9zSlsqSbtXj56
FzMdp8+q9Is8KBM0xp5QeSuE5lrQFJdyF7wEP4whjXFoOgRA6BXsEDmzTEG6SuI9MYF2zrO9jUk4
wv3yT0grM7hHNptwsIF7cUbTwzJGYG+4yk8NEd6U1BjN90JplKmqptSkUFya+VfZZP0veoUiX/+n
KxlCg2NgN74QYgi0j7Fe0lN0FolIGANfQof0/WVdRVN0X0fy50NmFgbdqUZalyaT7/YswBNQWK7P
Wyurt7WJn3P6w9z+iFEEC2EK5nHGeZvyiyC5Ns5S+zUIqmO4fZQM0g0GWDfWFX1Xol5LQYCse1YH
D90QilIycRzC95NFFFUO+gy/XdeCUFGtRcZfYWFSdu5DELpDQKQVRX3eRSuBB9j0JWflEzwgNGYr
cDLTUh1WFu6QVzNGTsH4owtpfZQEmX6edBq7bOapb7hT9D3kebZw22Yd66I9uuWQmSAtWTT8sxNh
R9pP1hPngJROz1TuxlF5SOvfghwKrhrQzcaPhNms6HPJYi/7PTOz/WZMinTb8PcWPc9iOUqzoMMf
/EVMXCDefnCKQO3Hlp6YihBwn2sqUmxKx70o7RIRL1RKAtyOWiTZgSSkj4s42Vzagu5zM5ZyPQI4
/nUxQfblnCDxOhbWeU47Plg0xvDy+vA+6aHGXvxktRHgsdg/upfh1fWfY0r1vkT6da4IMgvBYxlK
Uxj3jiw6R+OB7UBKyqj8zVrwBp8wLL+1TJ/MTtxQDTyV/wekoO0p1ChRVAvgLpgDvTAnAzhd8DwA
vVedDkC/YyQ8TBLME1znHappqr5tn4Oqqgx3a9jeaA+3RXJ/QDXh48n/KjftAD3FuFV9fU4QQ0XI
bPdUEfeeDSM6fs5uR/nHe8xOGxRdS1dI7Qx6RuO+VumW3INU/rCZz0iu69ilHccB8nKRa+GDJpCW
ohiiCmrWKI/PMGjZ2yg4oIlzxQq/JUsGEWQURVeae3xomrAFkvfGdhDVZdoDjNigXniHeWkiPKan
l++ZBcIU5IFBq0blo+M4nq3wYO3zDqTKlCgV838lS1DKuUZzfyfYbLu2rZLkhYh5StuxJXNFDuYY
92a6vLwYtEE9y2QbbSUf3agqKsajXel/6jDnlv0ISTd+FZb7RIZTQ0onkC/VkmqJRBpJeWYW2WzB
3VaMSiikAXogoxxSuhPCXWTPTHZyAIaq0qygDJNRpP2ij75ry3uR+N4nsThhgH4iz49YKdrVp2v0
JmbQa0VjfeBDItLms0YrgQVBmrXlYFGSjgh/EchWbeZxkaiUiBiFKGu6iUUO8KDGGjtYBuJOKj3c
4wXVBdSFh9f7FYQSZrwzu5f/T/DeY7mPmCM1jmC8j7UZrn38RXIADzHaYTBhpipHoBDJNFkDsHG9
CLlWNjzTsdjaScsm0RRt+Fq7JXFlkL/pfOh57175y1S64oE8opn15Dx4nFlqWPZTTn9o7BEsAmGs
gsTVVyO9adMZHfoFF90VtPTG4Mcv3SeWxStxRLbqAM8a+uO5TcqeziM2a3/HQp/GBuoy210jNYv/
VOx7Gg7xdgxDSTDouvTp/OLHCP5F8WjRVXAAQBk0BY7vMpcGTHHJU+46OH+C1qgoAj6EV8D4qy3G
feg+DK8+7Pd5oyCpxEbvMcNx2lDWh08KDAAQhbglLfqGYQugIspIx4Jp/T5vBCrUHNwFjCCdAybl
wapG2TrNZ0i7EOcBo9S89J9HEr07cZwLDG9RfkqgVSy2n4gFdNxhtm6rMx0MxJRqAJrmqMDddtuP
KUz6zLLARl+Nw0bSZ1jSTDJp61K2p3mPV7qa1bjZkZnMgW86sAf7tIMOmkdZJdnnd9bjGVEZjGz3
C33z9NO7xIZHsthpDWtjvSl2TWecJya0u8GSxRQ3zSOd1OWeAvn03z6SSzpdMvZIJAibo4EUXIzx
B7E9Qij+LBpd0rFujfqEB1HVbtV5cewqG+19Du6AjA0ynhgQV2FHGzEsg0H2jwd/Y8EEYGj0fhIm
pCwV5a4haLE+ykjURPtNqeg6xoxyaXfOtK3nW6rouWT4Fspa0AHOumnwsLaoFmv2e/AKMpGUx8T7
scBJo6J3U2cqjWMw/JVCzNZ+L0NMEtn6BziK7c5EPCStKJcLuLXy1VsyPtI7B1WOYVG0BAyk2Pqw
7iNdBr8nFl8EpqDEK+6jvBEP8h2nBJzWFlZWORb1lgKiv7GXulYRqvZDZCTOKi0V5056bcUKWpzB
zb4MG2jpGmuSU6gPqrZ2UVHhQ6nofCsTmZ4ryvVn4S0ZlNjfv9cGYzAS0/tuhM4EFfZv2SyQi4sq
IidtnxN55mVqS5r4d2Ov6Mf/7E+4ulSMtaripuvSQcqLIL3hL3UluWOoj4YBp8PcB1tcNi8Kbm2c
oqCYELtwXV3biUyZmBEQu4FAj5JqmOaBBOpMa8ZYOfDKrhk0Fk/W2XZeofIrm8AjaIjcnIrdoUdg
0pEC4AtgTgXsHXe0yP1kG9G0dq3t/xdOGA7VZgM3w0nDG38IxxqSkADtmPunwZgXq1awcZswsNNP
6qGXJ4j8FmvrCHNv5sk/lMhd0ys9/nziCDMl7OpUMNlOSl2ywn9D/dHRRdSdU6Y/IGVL8xCyrvJ0
zBFvodts3EGeVauIiPilen6Bd5GrDojygmncpWjXe9ZtRnPM2mbFf48rMd6jUcSsZYKAm0oVEVM0
ojtLKFWBmarG8LzXAwQkIoK3vUm3Ub1VYLW5MpvjRHPSl5KO0jU1IYwPOLSaC6ZBcLBwmESxzgen
jovU7lPKSv6hR4Mecq2MDnWKyBDE4Q9upcN+KRS0/Y0VQwrtszYe7FntceT+xOG2AZbJHcmd9vNq
C/I2qEMg5FAsvZWXuwIKP7DWrA9psshjNZCX6suqxV90OV3agnqZ7N4bUrXs4LjiZdfl95JvWVgN
tPl9gfra7p+nCTQjpZbjWRvUUA+Ptq7nh2GvSzLS5RPD4g5uZaLsB8cZ3WIOcdSXbCHo7oisyuQh
wCYUQp3LglwvwFZWLDMA4UgkfY1kTZKx24K1y/3R/y9J0LNo3VHA/eERyUbwBzLxjgXEUlGadTJL
4wZm5pl9gV7W/46dfjpct/r1ABSgDxtGosVxWqPKGAnEBPnUCAhnExJV5a6OFpkqz5zLbjvlD+0V
/0teFDoA4sKLKqou07Bun/20f614sVO8ZFFrkUEBBh0amwufMnIGGx/54/cFYNKKbcJiOpf3MIFG
mbTLOP5UDEPIkF318lKvmH8OkrXMKGZcXX4j/OZyNhbnX4LcknJoZcH7SzVNvhdjwyg39EnOvc6y
ih7ZOlpsHdHbKdejLxEDJo47bLk/cYrCN0nZ6O0U/8rlGlz8jaDdmOpj5uJwC7i/wrDMUXwQ7D3A
0Rl8v+nO2mh1bxadGs7qAKLkpzT+hn2D3SyklJ6Z6dsbYMsSBt4xDP+JJ6pYeQdPPsLvRIVZpowQ
/IAsan6LmFyM1XIY4w8/8OyiiMsN1cEJ1/ltpzxmnraxwrVMhI3HfpgpRbu4DGqaDGHyEkwyA/Vs
XIokldR23fsjJcMnTVB/8zVBWGVSbQ/fmXzHFjNYHyJfLqpGO4L3zUZa8G98eHQPgWqdaDM4eCQ5
HSrzYTm3qu8pvJHklPXLYgO4tPJfOXdLDqN7mzB4Dy9obLuLHkjY7EYfl3eIINbOVaaERwR9Y65e
L6+68v9knlm+lRvi45m4/knoF/a7hfFvGIXqunSCOwLd/3F0uipu2nUL75W1+QM+u6domKSegu9K
wRor5m+TK1jrPuxO83CCt+U5+zRomKvpC7z9eYa3tQN6yPCGV45YqEZ0YUT+17TEHcROfH1RWHh6
FOWk3ldWeVBGz3+VgMNj9a2M968Tmjki5MWQcDoxQPU2lkmqABeITtnhCTK4kwZr/JfgxLjlB+DL
d02WG76VmikeUbkmxwp99sHp2TnQjxwoIjaWHTx6lS4e7L/ZajQ5aG/13VLjuWP8HaCH2Q4MIiL1
O7PK7G088RKdn7q+LRKuq0Que29/prQWGOwepmUgiSi+mxMrUH968nfcLYeIyvZ6h7GnHc3QdlsG
IWJ4kmXTVkFS1KS9QUOoLF+reZLst5TpurzaCSrH6L2YYXMv2TQTAIB7TxbbaW7LbEqNyNVt2frt
Fa7mJWinnwA/hjpO/5EFNrpHHtdnAD8LVPMNqMN6uFrY8UknvhPVe7735E651SRdXHdRu5XDl7ys
XvZsGKvFU29/ofolStwSzbvueft68LTwR0+uSMFygMUs7rzi7rt/a4cBoO7lHdZzyVZSJrdsZ8S8
vOkjEzUWBzTz0RKm9j+h+VVkXOJ4VzG/rdo8FNfbxpiCGMvYuBvsCxHzC38u/NDh1dp8pL2wz4/0
qt24DwUXqR0zJRTxnCrvj2eeGsPh/fBZn4jiUtHO8UXaVlZKmQdySoxtl53aKEBh1WdcX8f7vIpJ
bhEg5JfegeHhI2F5KU5VPuNfDdDsRKYSzYiujc22vrE/JjnFaUdMgroPpEePPxIHuSIoi8pEwrg1
bYegN3VaxgkW9ocCrh9hT6ZYOEazNSJNpUDp4Lpe4I7ql1WASfe3KmdYk9SlCX8EMkW10iR6C3gb
g5PBmt5XCfVQxfe3BfUF9MRMpj2SWONuUOiRtvfA9zrvT5OQtb5+EnMdr80IXCoU7Cr3bJAR+q3I
R7MGnAQEjKvgchFXk9OScUzhNlrkNAqio6aHv0rlQGv7o5HqKk6GSjclUy93GJshnTgTCw5cwIwb
1FetV719VJT3R3xCGr0nPsopv2fsZIlyu2FQT/K9d3SoEoK3/XlwBmUrLYjb/9H7VhFCnyjUSmU3
PtgnJJSZVk+wXM0NPh5a2NpDTJ0fqU23PdljTJz20iKs0fXRPLDJNeKDxUFUb/K/eaTXc0FkWH8W
yBH36FQddCjH/mi4s4JE0yXRjibskRvUFU/xiS0VZJAcXf7DV0h/++FF2Q0uWcYcNWotSeQEGBIH
fuR9pBX+7xtmDGnmIytj4qPa7hZXPv7k1K1DjHn0RLmoFmRirWIc32QP7piGy8tfFubtybjQQq8U
skKb6WTMA5adYrLulsvNtzFjAU8gzhCHLE/4SFePsRETHSV+TqjSJ0AhA/09ShTnfu/+k6ZpK3JX
rToAPQPWPPLzGQDVYc5uRrEDDmfRDMjtqMHoYLYPEbdJWTl0JXtgoPSsUHk1A/Jh1WrgPETTA+ai
SapsyOGH92xXMTw3aLtvpeatw5CsZiz9q5fQkhcskZqU2+LxFQ7aQDD8H8DJ2tW0RktXc1FyHv+r
tXU2WwdYsZRshfChhor+FRSrL7jVjlxK1GpV8Tu9ToYjhRrOEG4o3fefkGc2eR+1NlkA+qhSXr3o
O85bzVZyJC/HZzt2z1J3sDxt4Kohf3T/WXT1Y+JJRBUBkGLoLlyEl/TCAVijAM6dlpRTmnd/zpKO
a5K8NtJt6B6WqLvqQ/oNzAtrlWUQtXsVARtzoVdmi8kmrWky92+6dmJJZCPPJhGojwE8CtdHKITj
TKiCpT1yOEVpJx3gzSl4nvXkX6keZGVzeTNjfnEnalQeFqm6LXubT4fYBM+952CoofsXQVYBKV6R
9IP215AvWQh51mki1TyVO89ptLOgPrYHsJsE4D1oAZptcsoWFjw/NQXXSRsGAK2W1VxyNiv1QpDZ
mLGn0ETYwYtua/L3mxZCLXZjKwg9mZ1/2UPPkzt50AKVaMmhVWCrTfNeq3I8ycIqN07D6PquJamF
naO7rOzeuwVau3CnmVS+uOka2BGYUQM4N8ijFJJPVFfNuzrYCT2ypbfUE4pqfbEhecO4Pm3p+IRx
VzfmEbCsNeyLpniuX/qbxQomw9WMqg8tKAoymi88mtBvsDk7IrpL4GK9In47FTXs3+qlFMh/MwwB
TCG4+LO1WQc6zINCTNubw0gtYAjo3TrwY6r2nj/E0zIWDC/A2mDV/XKoAg6WDwL1lgDWzpXjs1HC
bVAjNaz/LB/iC7mnNsSWobT6fUFGadwNNgM55QEcWuj8BE/OHc3hhf4rvy6J9LA0ZE9Y5A1BQloc
LDGMCRu44DU8Vu++8zzDQwHX1okxd1CrTgmLIx1XQ/VROtzjUDcfG3K0wzLUmWQGzeq6Kabpur86
jomxBT8dQ1EJTansUSAaviYnEdJpjY+c47PmJsjKE18uKnpKOL+dYowTyQGfusDPwzgbGRimuWgk
/flUX0t2lkuenwntL452EBvzTv9gA9Xavza7oH7FD7sywo8tlx/DVYdIFEG2pJxMMI93P/zgo7Do
7wBFe0RxXtNj3cawW/LD6t6r+LZ/Pj1Wo1v1Lj2IfyjLpI+cz0bdGAEzrlK03QZEjeg+D8k2zDUF
nrWQOsHrzTlKIMi+Kw0lh7x1b7FayULGf2MKwxRYsNLWjPNVqM1KroUDmhDeec/tQ6pq2Q17wcaZ
tmkXooI/ontT/CNJNV9Bmmwru9dfm7PlY3W+HIZT9pHJdcPp+uojwe5D/Vr8zcYTY2/4+qlCE34H
7Nrz0S7GME0K7v7cqOa0m5tZI+RvjiWVW8YfDYBpjMwTOwdwOveDXd9fUdkVdM9jQzwrC+k1hr7t
tjMGegnAxc9SOQ64hHz4MCsYn9eOjY1Jpg9NlwbQJR4guqjqzQkyzchXKUDWFrsttENOxwr96gx8
4CmgkaCg2+CNqZkGxXxZqkOQCWu8IgPQub49aW3MNoS0or9otPyziE0i9Boky8chKrBdBXHLUpL/
0u5KrYY8gigAqRloF6lnMdKyScDlCUExBu0F0G+3g38cZSDqqdA1zz+FN+qcnv1pxx070iWo4jGs
36TKKQ7DDFiZGai6+u2SbVgFAvH2pWqjVfGkU2KrJMhUf+tViL8nw0Y5mzquICxrkze0yXQ48cDV
JBV7TtHiZAOe8snQ6vXr6Swc3dSPsL/091QZIPMVQtq44V6i/JptnI3yxUzQT93ZORSyCHm+wT31
tsKyo51SUcb/Cvo8BTqm1NGFQO6BCm/72MTPeEV/3g0+V70ooRSReo8mPj/k3NMq5JgN2fNd6fb9
Se/I7njbBD9MEwL7iXDtQfGfi5mBG0Q10mAN+IJx1vxnwCJfCFN/du3JjFniehipF4GUl6+i1Veq
eQk6dQPAo+j3WkwTGbMg5WBbQydiuISpTb6s2R6J3jrhft3FE2Z+wMSCY3inrx/nF2SLZT59Ttaw
sJZNpHLuBKIK0xaNrIh+8SOkC1awqy5xohhzQMo319jq75w8F1fNvOTnPdNacjDkRb4QrGe3dLE8
rxq5AWe+j6gVUbPq+Yow98mUvanY3kLTruq0F7zjXZ5EkWge3qzk151QyebZxSfNhi9TK13Ab510
5fZTeU9Yeur+wxsh0DuJvQ8pHK1XDRyRcIOvPbaGe3jpu3zbMqs52e4sNXse+PBZlY213+bbsLG1
jJO5omyaqh4joNeUTcwsjldtoHd3JKVP5r6DrUsEiN1QSpnSwMvE3w0Y2OJJwR9rSPP/FX8Y/yY4
ABoCb0NxigJ9yv8lgly2qfhHQtXxGuri3K3Jurv+Glq8OngbWqG99llpyhii1ANqAmBSP2Gdm6md
EtghGrWIz8b8qfyVTdDYNQwaSdXMx3nwTCdDT1ymQcNkx2XV379AjR7O0CUkQBYgRC5DoSCTLPra
fx3Oj5TdapWforEEZ+P5zViEKqA3N5nO6j1riU5msJrJZ+ctwmvask7a4o8mear1VRP2iNlNuZaA
9ebY6CntBWUE2aVMU/3GirptH7c93oL31E7eb7Sk9hVXafMQe1+EdJzNueGqBtbv4Q7hNFQZ3A+B
a9jo35rpsLjRDNVxRnvRC4wnCNHK5CUUFPvA8lquwjCHJQ528rKAzcnz6PORNW+uiS0OJOU9gMuI
neVdaXx5hO6M52a7fWDWWIS5vTy6fxXVuinDuu3OQOWqNuUPAHkDUymJWsyhgRmhBmGiXq1MTBPK
iQEY2I5Z/RunXqEUL/i8TWYMO9/msSpbVAvKH/EjY1Tg5ok+Ob7ggnFxpPxoqFXPxHIqvMDWU8zm
xoOoQyMBdEdMjYZAjNpEU4JIQQNiUy31Lk5vXhHA3t8++8Pv1u7UA1uaMCEbpgO6UbNfg0u0/6an
Sb5Mxke01CeTZKCJgFBXf8id/PTNPuyIU5AIb0O6h0STUt0aff7K+apWu8eA5nHEMWS+yWnYR6l/
wnlzuwPJ6nGpV6kY/oa4AYm7QfkPXGyCgjXxYpSLolc4th1uzkC6N7wnhEyz7qtJ4IwD3sBtmQfh
Qpw+Nyb9HmYghUGPtcJz08/gHCDYCeObmlTS9Ne9D9E1T2gki9kYSsid8cz/eG/bQcBNl1ozQFyz
Ksm3HQW8BDVURT+tArNxh/5JnYhzDcLbpxFNuYxZeBYpdaPTfhnL23HJ+6uYHET5Yy1o/hh0A20t
eVZlAZcf/jiZLSm6EjLw4OtZQjsWYCw+aKyDkS+jP3mdK/gVlPWe2LOVK0s9zh2pbAVTw0/gRpJT
61zmojnqsT8pYAwWbXYH7VnM67/pyd9e2ytHJ0/FkS13cFQURoDoWbe9NeHL5ti6KSf08WdVThhD
BoR8uamEKDTLZg7a/V88n6oKJWCmN8vNbUztw0lp2ySXfaGEBxpH7IGMBdBZUM/rKPo3jEXfDKDW
3M7zkD/fiMBgY1wsaSguVhYAECozK1sIgvO5KWN6ceM4pJ+PJTWm1RuhV09fSoEi7SoQI2iSc8ZY
IhtnlqSYo6aOLTfGbR1HHSHaG/xLzDrIcGCI/AUrfUkUS9M3g4PM3fK2p2faODB/DxAGilXeoEhc
K0clMoryzFwRQgzMWEc8Di8G4Rn70Veb0CPP9d0WFMQyXnSoyr0V5ackjJKa1PzTuiXClJV4Vs3m
8Gg5kv2bFxjdkWlRps85toaXlrXSNB2Y3FGDaLRxaubxHYu3SKrNckJw6C+CxW5fQ0Hg7Vmt45nG
Ja5YAM8PL6/MDfcO+oHe/j8vfEuTVGW388+8TIe04CBNhXJuDpwkXqrzoe8DfADXfASQQzXwDFto
LlU35J8KZ/BlvGOWCjBk9U+Mk8CtM+8eS4PnnRDFvgtyK3lKCcMN/B9hoT5r/YGlTe4FPGNqr/mD
3E5RhZPrO19ntHdrbFDQv5v07/ynrK86JkbN27GC8hEkUcQFftXuMXc9RSqV6fSb/zbU36OBP03g
bKzMsVUu7PLBPshvrrUvDH144JCgc1Tss8fyhMZOEgpVu7vRbzBTEWU4pHc0mKW/KnAjCgPZ0WsP
yGYFrWuiPCRUiDF5BgngC7MiONPEjGqJ7aoa8YzgIVwO9J3V4fEq3HJ2PxSTtZ3wjC0wXSAQTRHR
qXJiWJq+F0jiYC7VjYInJnQexg4xa5PxV6U+pBxp/uNXiLoeShAlEyvp4iA+GbtfIEFbdETisCfp
O6E7gdjTuC2r53QcSxawZG8NDEqRv4hwVli/NdqIWQQRqyLFDmDQpV4vxm1a7fU9a1zlUEIR5lN9
Q4ehkRZP+mCuqwPQL9kxQcVzj0XIR17DWVKmvvsa1wk1suwVCg5ip5f9Mo8OxQEmZE/9pJxf9Awa
6VSUXVCxd4vWYW7pdZKtlLeHPzJ4CkzmPk1yynT3j4ZqkTf/SDBKjS+V14Tz+E4HywNbict4zQIb
Z6P2puMqTxzKlT4OjpHTc1DqdjroGkJR3BgwJu7npYxbM5fvfVnki3hQI2aD2xmPSNKY/9XVkzDe
7GS8yAvmLWVDxvUmTwfo8McJ0CAi2txrH6fD5JuH1Vc6xqWbh1G9V64hgnZp5cBU7O2JpvG4+7kz
Ugo0a4QHUCkZjPByT1wwG4dv3DDaJ/jmJX714jKixezuyZt5d4guL8h2dNxoJPWq00NfZncBJ2MD
bphUjrlLsSpqmB1LLtCoOjEeOBkVUG8j0e2JSXC7AnjypycQCQQZ/rBSxLvU2VyGLGft03TkZ4ev
tGenqEgNjNI0TAckuqHUTLzFRDfcrtKUAxhZdgzgw5KoPgy9tawznJXEfjJK2uFhu3y183+oiKm1
1Jq88V2qXPDvDvBwsJTV4G9i1mG2iIoHW+Op5KEfr80Soj6KQ0lwlZPvJlXROKItKgQRx0whmUDq
70jGnDlr4KoxdO3sWKpOE8SWrGhvcMQomix9Z0GTbcMJYkecTiCYagfSASICIFBCDCb9mT4VnVM+
HhLAsCVsnfHfGI4bcjtTSljh3cTXxgvky8+HUAwGCR2L6zcu/xjQGw/hnTE7Yks4ITnxLM4hFpcM
AU5HifoOfg7eOU7WT2VvwCYOUFYwlt2K5oVwK1MAK0I+VOU3urLW9nBlADp7+Dj6rcu4kDdLY5Q1
Pmi3vOQ9r8I66hV9nCGTds3AABKQSrXCUzqlPAW/BiuxCZm5A8sWfM6WNIkMx3c/aSwlRoDpncKc
zCVDQ4hCR/rg3HzcxFswE7x4NOL5xysQPmJ7tKuYts05lvlK4nknvjg1EA6YAkVN2h9bLtKHviUa
U113zkGDVdEuGRvyQZbWIS454Dn63dCr6BgC2yqmUw4ZZZPR2rSUC4EMbasuJpIhbcdXxDBvXxmA
JZ0seULKIWqPf5YCgm/RNtAOJWx/MglsEU1yPy5/9qfvmN8O2r9Ii9p8BMndGDT+F4ixkABFNuMr
hsecW9g360lPfFPl0NOxaAblzwxc6P2B6yNUi8bARPTrR5hhyOMZlmwfoUlaV4Hh18BtbammrNz1
FC9MwEkjPypsrfzIj2Ky6zREbzQwlw/Bo6Ilog66YVnrC6DVLn7EkC4a8ajRtUC9Js4fUCEWPLKh
1aoqWCHJzIAQijd1llay1WknwNswzr9XwXbl8WFQUfSdrhkBF5ecMVCADqKftktftnDizS1hMCxP
LtFhpNmvls9H8G2RjzoM8MHbCvwW8xCPjBE34ywfEbj6Ri7CbGTy8Gs1a5hqIBVsYG/3yUzKco9V
BukypdsdNqv3mi5NvEyN9WC4CPr9JplHsEo2whF1Oj0GywBA5pcCbdJ6bpFkhP7mAyhu0mUdvLuV
zxTdEubozMLD/zBavPrh7k1H4Bj0qBbj658Q9tN+h0sNhrM/3XyO2CarK/YkMNn71Phra78uE161
CGcEXryRsorYT4YO/bOVAUSz8gvp50+YTFNLSKCYw3rIi7FGmS3zyta7+9AZ9EB2HhEVxJvtDALy
kDjDhqYorM/D1RxN4MLEwuSpA422xf0oREPb2DggU23ma/YwVVENsJO98ytkVdVvhiV+bPgi5GqD
UwKyhSzDblCcBnCZfUq+PZl3qeJp3Kkcvv0C0E7sXAcuSqSCt8rNqU3gOGTSUZqBimCi11veYvs5
1FLPhW7eGPiDKTZm2L+p/xbdmmScDVpr+4bhw5hThSTyFuip/lkNNyMhAZMt+puHddoajmz3Pgi0
QcBh8KYxX2VCcifuJ2IVJcVdRlfxDiHDEszqKPi6KjwOVheT6yT4OPRKH+CsGgz28JA6gf9QEp7s
sMnIIdcYkuDsVYL/NG5fXwnFOFGGcR7eFGyZSszDnYUFIH3+C08EPhaifCKR2dSRQLKcsAjCx5Ge
393rHO2GD493OSvUtxDxQH3qvRKRbY2KAsfAsLLSk8gVm/UjG9F25yuSh+qokS1xEcaHyuEHedi8
KdzZ56aWDAoeV8UoTIsYqUs/6g9727M8K3bdJiGLNPJoMV2rVe3JTn0nNAAXDSrZVYa7iOZ7YCJB
IM6EEVMCrHujpDWZ+mtZMWGBNPM4EyBUblATB7ttp9NxNg0Hub8+spOKn8AbEw6foT+WwYs+/JMJ
5yzSx13toGZEQvJSBM80MXNj4p5Ec+zoKqtS+NH/ae3H5lhQJyGIJTagdJ6YmYwQV4OBicGaUwRC
Yj/nbvaZUPrqfgmqWICh7Nm+99a44nO0/vLuzbRBxhA5RRgzUvWHOfRWoGDNGisom0LV5ZiBSSGO
mAc1xYGb0m4gUqACJjSWyi4vCROTM8ZJrDFJHN8XzZFmSqeJ8Ypzg9NI7KJW2uC6hBZ1bmDoOKul
zcQSi7IdCE3XA7l+A8KHNjLJxqWPcuDSiYgdBbZCWXJpsNk6VqZauevoIyVdpL+QNXzk/TiSZXLk
+9QY/mH3L0BqNE5axDicrDpbMcSsRj4HyvEHuFrmNHZeAtvkpL3qF9HmIKoHhNjZAgjiiFJcik5X
5d4hmdgm2hV6DY4naJv6i7spAAEWa/RvIUZEdOouz3qYxCRcFESys/tx1Diso8o6F4duOZ8zVtbb
WAO6wtdb7meWJDawCWa+5uBhrRAoOtqJR0APgsGU3a+CJZGZFdceXW5Oh/kbcXltvOoV8AD0JHHf
iBjtxtFxHeR+lTJn7G67HLOW5GVS9Ry58ViTGWzZeyXwFZOORhSR9wlBebJnJ5o49NDWuY956AKy
/ZILu8Yu1zmsFu7QV/ez+IYb5Xn5TYq09LGqj114EKnvlKzZ4wOP/5GflCuY0y9Kw5L/x9T74PDB
CDWlGG4gKbCWqVOIdeNVVJrDC6lN5oSfDjMFmCYaZViRNrdF+bP6sWyEaNecuOLkT0ks+wW0L2aj
TJQ2JoRrkVo4RF+zJI34UKnD88jaPwYl434pQ2CUjpeczBcFcKQdXhPUHWqH9Wn/SUJXqwYbvCOT
efpMeIYq8fmsYL7anW4ofVRH5HlXKbAsxPLdKb7kLlt1ogs2zJfVzJViiJDna14wKsOSf/CeoEED
NjQYpkgMt47sDo2zstilXpTcjDBu/E5oxrxlZaarXR3owvTx4h5niccPhQsY5wFE2crzQ+c/sAtx
qRhybp6jMLJBnmvkmEBo2DDVSMiGWwbNvg+wti/Qf38KMKj1BOvUfrNBN/svewp8SZCA4YLwuPV0
b7kT0eGobmRn4cCAg4TF69MoGIyudbJHXZgejfbFZ4iKGks5Gf3bZVxIXo0P3mJ0HrfkaafjU1tT
QtAwmQWE0HtrkCamr0PrUJJBr+Af135NjBispY37aSQ+i78QDLUJ7tE1wcXbnWDMMZkcuxHhpiJ+
r+21d8Ct37ODzlpAhqiQgD0JG0Zo97RG50LitAGBptJQuVF6heZMNbfmCmadwmemTtH86ptOtEg2
qR7MMdVcuHLa3brv6oCkaX3rO1mV5a4zBjbnKZXa1DI10cV8F3rw9LLCZ9oNC8aisIPs0xxiLp7O
OC5ZRQ4S245uJ+BMnj4UoX0EcOgoc5EHR502B1p8V4rDutolD7b7w34xOvcJ1650d3UOFQCrB16u
oBerwLvGI9OkgpQrbsvWasib50TrqNXpJ7z1PgH3x4fFI/0WRdS6yca1H0aMrEvZ8PQKQ8oZ0ZIq
vxpn6Hmb4Xz1932Y9DCtXKNh0z0m8IPPziVHflDZvCKec8bYKeuj2baWbhZuwFKk35RPRrbV6AuN
mTNpYGcBy9Kn4YFpH5VGH2drXNIuqNODPiUnEYu9MiFBVwaGFZfdPOHMN3xh0Qkwq30/CYEsTo3E
Tgc5o8/ppEvunRUlA2o5luaoyGy+YYsndYJvRr7XC6SI89Vs9ipJU5WKQM+yGnEPrTCYWNFhgDBZ
8u4h++gjZ+zOtg8mPQVNtOTVjonLEXsle28IMGGPwcaH/ANSC4+BUem7rGd5PBM9/ujw4bYTQqAR
7Iyd9yVNUhsdU5qePPHffaiHplw83JVFQyDiH5+yOAaL8Gwhep1jK+6JxUQFAKPnuVcjYg1ZOpB7
mRACUab3bWpVx/OaXS3KZTLtl7Sghgre/0AQarLXQgmCthZU5J4TfYgSmXDEZZiHGqeUsX2vda9C
zh1ARErBXLS8bjh6OGxooWgKMivj/hPMOwfPpj8jAIjGpyc3oi1YNFvuH+kDaKlsZf8yPPzoYqLR
7ma0xQDqhmTz4SpaEfs+TxMRxrI+TpXZBBWkKZpRNFVda/PB67fTOzKrzNN2jo1SMa8axDa1rVct
641ax+GqiW4J4y5FVIkr9Yso6JsB+hAtSMguwcMYWw3D0cA7AFebDtDuusiy9u6ww7XFWOh/M4nB
nfa0lCgEJE9nzNek8wDzMu6ywTuSS5S7KZDspqd1OCH0rLZoeOg/KspBpDSUy0ehOGMNhsJhhwVE
AfnV8r7eqxYtRL4xdsCtofzDRVc7w3cn23v1MToral+R/VQi0vAnXSFKoxfHYLtjPUBCdilHN87j
LbpHWXTdpsNxpqE+iCZVZyvJ/jv80nsjoeGiSTvDvpgSJehUqR+EUWzds6Por6n4D0amsjp3/Q8K
20IlSCN2NyS9zMTpzDf3gjdNWDuuQXtVLPWyhYoz4SmYOBuY+S0t8KUEqOXwmG85pa/6KIVZ+jY3
/8gFZ2HP7GmopRh3S4JW+sTwPX+FetVSaPOE7OV+haRfG/54PIiVFYiF28nUv9IRotIqsU8e0DVj
5X/WL6PAHtvieWCtEZ+qKwk7LwzmgCOYcNeQjUAZA9iM8Do2/vz2kblQ2Qk3US1jiEpDoSA/uO0X
V601OcIkidJlUbNO/DaIs8QVcsmCifdVpe7ruL2b3sPOJD892LLxosrdkJgyrWE0N9poD8rW6zIW
VIf9Ab0kJP3y61Hvj/2bg2/3hr3iR605xiQKBs/R4uCUVjLbAzb1/ldhOBn53XzxjbbbgCuowP/S
gAJQL8rzmMd/o09dBG9N+sA/y9qQ1DRJndTcNfk938blN5Qf4bxpOIhP7UN+UoL1GWJAll1ZXWiy
628S3KB9ZJFqmdoYq0n32qKsc7TCEo0KsyXhU4tCF+QTGRz/+fM3vOvWAvkYJNJL74xbXn2lKfC9
AfjTaiYB6jSQZOok7aj88BatwiuvNjbSaFtNlzp0f6G41LhqyDA5ngVezTq69RGMdGHf5SAFDMlr
/cM4BKrVEpcbtSCcBj41z6q/EDH8myzpkXXses5ysn3I4nian+Rr3JH4JiP1O9uaZfrVBmcQFlqr
wnmLIq01WX0MxDt+7KGNuEoZP6ti6Dx3NwRp0HEYdu3+ceUykm4ZqP9fkHwwId5hbWbzdVnFbhSX
qpwxpNTqnvXKzqKIHieKq2PQUbjrn9wVZcm/jcAZOik3atT3xnCSDX33ClPCUxM/JNwzXTMrVhvV
yaj9hCy5G2+MnCRQJHpNV7n41TC77PAh/B5Fm+NtR6Oe0xnB5c7jeL2OChKtFm4fF7+dRG1/lEFv
UnkripjE++9bTtJg4mt+CjbhuJIqBQNyAwyIO+E5vYUhu4YaNn9O4nmyG5H9+YdMkkANBAU9JJUy
qYjzOb+nx5NTWejtPtqhXk8GqFp6M2U08HobcTrxXjcnM1Gtcj/UpFkpUqaEiOBwUM7vC+fwm5P4
ZD8y4+6hyw93sz0ti5ioAwYCurQdasJkD5Zc/ANDFeblPGme0hXzFrXWHP127utkrOr+iwDl7un+
Fxv6wa3cwLVbTnS4FMcvsikeLB0okjY+IDvLQdJwJguGDb6qQO1MPgRywlfeSMOCzPPDguGOsstf
BThaXwVxOXx0Op88ZOS3Xxbawdd1gTZ9drb2SpYgmcMmEOO76KbkO8ym6KJmLt5U8Bh6gpgp6Piu
vl364LFdT+p683SEHbmdTwhJjBSWNqhkpT1jY5utWKwKNxNp3/Xuz/Mi6Pc64a++hp7RbkFeY0Qr
sK9MMswgh1nat7XX6pGaA/MYvUdKu9fmzRe65ePRx93rE4BvmecQ0bbijc/AguvtX0otmNslfmmb
VPDhfs0AUqcYkQxQp9/3RauY6FThlCyL3xzi/iooURt7btqHwtzhxvmEMsinetx6UKtaqPmBe/xI
5ELBPr3AmMUX+yF5f27E97U2pEOfJHY8kzOms4UA1V3fEIK4PZlrl6alRbkvj5+jberG80yakBPy
aebmrMZg4AXiPVeGk7IeFHVPBcuJut6b1YxIwGM0IF4dRkpBMqvqOOkgH9OA/HLAQbjGVSnzwt8O
Mys3EWoG4bXhI9YGzK2NkJGNScqfTymXMAejnyPinzO3YZ7zNtEoPcewqiZaB/TYnoCcMJncUVgG
A+CvzHcZtvrU8gA9NM1Cqkceh/eoseCRf4amK66Ha/YrJOAjSDQzcVLXerp+7+Io1GAYSbsn5bpE
nKq2zv+3v3fOf4+BCXdz1TzwMt1u26hKBgSJm4dzisqiV+1GtfzOjlQ9k+KZ8SOMjNzM1wiJrq8e
HaqiZH/hwcNmDQag/yuv+68QFkm+iHPNL1RRMT8y87EZa57YCGFwTZ8RUx5sM9b3SMEvRwgCOHQ/
PHhRhmiOKxkbXBZbZh8IBymIFu6lNaIxXegersxxOgpQBSjR7m5ZW+GzdQZaRdQh+QmqtRwHtOfq
SsnzbC3XG5mxZROMH03NozmQMeEk9Nd9G/pKrN4nTSqan68UVW9Y0TzCWK9QvBra6c6b0+Y7GMsL
2lpq5AczE+8moCKqU6QUFbqlWZjoYb2GYRC3qIg+FXUOL9hW0i/IdcADEc+koWzy6pe5/QeL7Xdy
MXWw8fhBlml9pUPHCqFq2ZSYAFGoIMKVwleOkcOEaf2XnOwP8r8EtBKNWGQtu0mXOzdV30wY+3sT
AqM6EgUrzE+GPbKcllt1gZhQcOQyFd8iLuDl026DfwRQ2pdPCKLPQmX6H6U0MqHtQLhl4K0J8cru
k9nvU+ED3qTH5Jwmn7JqQ23TEgbYXNycADUOIWjcwgEnwQcQzr0WcSe41spMKaK27KzN7rKpqcrJ
Z1Jk65xZICuK/WFpVsJ3HYz/k9pgqd1xVTaf5oXHB5ELAgFluofuQ0IWBzDsOmgY4RM+PojVBhQe
lxom0wHSQ2GIhgN83fhBAtENF5pBifaElDGCwC7x4TfL3Y8meqTSQLZJW2d0/tB17DLXxDC7X2P4
CkZEI+JVjRuva12U+Uvbx1SXZ1254YP49W/Ek5SPOAY24j5PFNYc8E2w35koCNLp/eyWwAAlJPNu
VLsx31hF1wdzb1FNDsUhxlfP/UyC7mKTJ+vc0rVsmnemyhYsaJtFNvafxu+tpaYQMzt2oZLSA0dG
ygSE0M9Pzyk6fquA48vhykCZHQxx/QZvO4tUYxe1OBGOg2SYXtSmHZZ0wdllx2SE1idiymxB9GMi
9bffjGanX+QbuKyWDLDPGvGwL9DqjqNQOLvbDQx9/U8aXk17ePf0XA4R77rnLvZFlhQlI4TlzXKl
0gACde0OUO1kl06BE69ml20UkNSAUNnOicjHTSsxK2H66wFnAu8URU60TxodYwpPZJ++Qmk2XkN9
/NZrtZ7X83qUSN2DwCIEiitrt+lsbeYnbQ9KPA3nEPqIvHhzR2QJur8ictIs+Vh8BhsKuIRyUKb5
9lMOGiBmPj2223U03zqhOEruB5SYsnxuyjsTUajPBPyamMn55qnGFlZNwCDen63cu4XIf6G0py4B
FyDXZr/5wQJYbWOEzNpoy31rmVbBCt2k/WDOyqc69Az0/7UxBcOIXMZkWN40t3ibaH2AkH7VrKEj
ptGxIf3PWwRDyEHJ4d5ddfqQxq2hnEI7zy4WghH5wOPJ2KZbi63XnheTQQg6l/lLbwc6dmf9Vtzq
M8avYFyOl0pWcD8mh0w8AjLJv2m9N1pPiOfJR9lb82UsOqI9VdjeFtKKWfxOShS6gDLgHRaWcj6h
o6WCBTOlrjJ0E3kPRADRSg4bEYYaZgiCHKV4e/Rznv7xCZ3om+SYgvQKLoLuIzngLxn9hba7xM8e
snPAPguIAFo+ghaNSGOb0gPzhSM5bTaCktyuDv5Hhe1u3gzoHX7Ms6Vx/8QW+Q2DbIsoyJRSv9OM
NCP7FtmCPpCbKEeJH9bSdH6TGcciSbQRhWK+TppO+nZgdtg/hDc+sbrQHW9N4yK1WKZqLHx/W4fg
ZRKvqOuxpGm6BxWYYuV89f6JFYLeXgc7dDrV0tMTBXaLQeEULfo6cVoTilTRXt7iFOGxJQOy/RDn
4PFTRo0fdXvMe1qErxxVtSzf21qaG667iRXwJsLdJdMiABqdtN1K/KL1ro+gqMNRClhgCnl5sAwb
RufFrTAuOkOxy6f9Xru7ukKyB2cXZLTWz/Rjrw3UJpaL9H6D7GJL7lDuY56Dbyfqk5GDNIaKmyak
F6xy0OgPVS07ZbwoNc8vM9Nf4am82Lm9GWcZEXaWjtq3f71LGzJ+dDNOs8/UZdWabx7SPtuHMqUL
n+7fwD6car8p1q4p7bdETw3L2OHdj+wSYYM4AEU2d4TrI1tNl8OWOnyjr9fDjid2SuVeomP+5729
Fs/xetfXfOkGRHckHnb2UADNaBDhbfkJDWlqk/leck/Ta4bYjnPjPvB/ZN4IHXTG0tmhyjOfTIn5
XPniDo6nXAE0EhBeF489f03i+TnN8CkTWo7PfUioE3JZjpxJOibjK3JKB9+pqWJRPRPOPU9No5iw
iCQVDDk6p2XWCCLRzN5bYGTpAZpJrLuWY7Ly9qb7OvxWvKBOoBU0MHPDK96TmaHBVDGhuRJgciFu
19CFlsB4LJId730bwvVGm+QaQFTq8QiUBNqXG7qfNSKVyNkBY4i/RFwjjv1c0tr7KsbKRYRzTS0L
HCiqY0hhpNpbqDqm0olGhVKp0yCwUYb+g/VMOM67E7Mj3NzNmuW+32+LpfcZ5Rmi/ZJqrzrfH2Pn
piDCrgNboYUcN8mRfAgciZLLdqt2HMnDpyHWfOR/5S2LEs8GRY4J0qlyCy0f7Sch/4EUOum9b6Wy
FM7wrWo392k2Pg1CVEqguzuYvvkoBd/HQJIkWIsbab+tN5w6pHfMJCsoWbtyeI3BUG4PlZRzM25t
5JmSomDx6DiPevqG0fYHrpvj1nbqREEpaWUdhmWnSPmDK5QQoi+Dl2O3IG01hNeVQssj8NT6pPf3
A7+8xAnlTCNTHPODMM8F6j+4ObBuXOSypRs8nMtK80OesSResRrsdSYbKtR51tUbQQuFSbRRadv4
Sj7fh9yN2s2T6wU9raAhFrFp55uyyduBu4dCFVQJrM5e1T77bhFsc2b3uOKs9UefWYULDj4P09Ji
evXviGex4LjXhPJPlUPd3KdQHJRb7rN4/S9Wizprv4cDqSQx8g2Pjl0qkD5qrfvR1pBdl5B/hc6+
kRqW+VX/HE2SQnc0RS4fSLURrRFKoTV91+uk6j23dhNC0PCzrhAPv8p7Al75nU5gPe+/KqbwpyYf
RE4Qad208SuPWkW2FCPYxlUalRGv6OIm3aqriYf5LSXcimao0aGtkoL0Ic9NEyLYHxNRmFfb5bls
tFQm44V/avTvSUdTINCzAcEI2Hp+42h3PqhKu4Vjbq6z6POZ1pPfftOTu9HM/wQZrJpzJOOuSWsU
GtJIxAVO7wzJ0UwlTcuvCRa9DsCKa1ljBVn0RDg7f7mra/719Ybph3SLIglGiS6m2WkMNfpSrdDl
Rck3djbIp8+G9UG68oUNzz3+CAZdqR14ntz+OatWOP9m/xJWx6M2AacdC2jEgh3E9OW7IP946+VT
Rj4iC6xhAOm3aYUBthKYWuyYaJvZRA+xt0r7wlJ++Q5LTn2U4z2IJfLdRz8nlUyAvJGw2QLB2slP
JNj3N4HXevgAvSKyxYaZK1mv4LEptngPYLUUC+NBgnt/2zd7UiHuo5iJu+xR4nPmrnwXQbqQyeyu
oQfxW8ZbWPif7RDapHYYVaN/Uc7ikRdYlnydzQgDsown1PmS+KBPdCYiOHDQ5F6kcevGSTStdWrz
HcZOrSFNAuaUQemlJ7hkXPs6KNeN8pUcGvkkiCSzbuE9CCwCljxv918/eMMGTmkMu2ussVve3xUv
bp+isUHwP5muHeV5HpoT6IkyfE+LWXMtnABW1s/hmc1/RUsm+2dtrbYeyngxDG7FSgKhV90jVzSv
jZGalHuXkdQXaC8syJrsxc1a8hrG1ey3FgIDCXV7LnTljMKcYlCX9CD/ZERTIXou+P8WDMSfO4g8
l9lR+lzSxkszgBG9XK63O5aOr+SMpOnxSaYyAtQ6gdrUtb4qlX2T8gX90xaIDj+nnjWM4HaytZOP
vlFBjMHlHvHae0z1vJx+/JX7tmGRRxAqDw0ca1TX2n2vGEiPwi+TyWHLG2iOTlGIK3SBDw63nTJ1
hJaAQb5wAZ9HzjKj7EArAtNb4+uEwOylJWBzNTFP3UTg89ccQA0TJz+/BVmhF/RmvBQWk1/Ui5u9
fVxd0k9R9OaTJnHHm2/DBLnDp+327lVJWV1s7B+4aj/PNCQP/u4dEEgxEdKT428dRZDvbMcN6iCK
VqBPpiHNEaSZvfDUTjkeekKmZ9NcPnt2PxKXL3kV6oa5lL7u08+6YSYEFxCqhb15oIJb+WPFCJkE
3uLzgNtLcWefjBeB3A78fzmolpPzM9qvc9mObfx1dzKE2DsTLgkfXLNOW5dHzbmhZzbNk9naeCQO
I0hfXHgB5U10BoSU3IjqMJqEwMaxLmlFyYatWodgB+ce0dCIQqrwSOPTWMoV1aR/7omq8kn5Rjt6
cgwT6vn6ZmYnXoF70oaH1fcv9B3IK+vPobMDTWFvRnTNMKdRxrVZ/jTedDzfH5TR/U6FQpLdEXZU
0CvB5ke6Krw0OBp7tix5mgWU9bY6cDVBhx90KiqSAcGpg5FauComB9tgWEyLvRaRlvuqA2AsUzlB
vysO4L907AIweEvWL20O+S37+Gi34+YKsfyYgmMYFoirnrfEN9MMT3uJn8J6p0VthKMXq16m6e6n
0zS88QlvOWJ/OxNelYBv8djRCTlG5HGgRwpQ8K0nIM0wteCYvAjqDabTinytoFlAB7sgXBmQMPwU
814WJsDoq7lphm+ofFhdhOrlzRXyma/L+xkgowisJGtxlW+asyIhbIgEEsGRpj0mSnhxPqmyD5PN
/OWLrkQks/miWxvDWFxiZkqdos7XVtELyP2SHF12U5k5LtAKuAnMl2qATsQ9f+OTvnC978TP4+t0
SZGJ27fnxZQPh8x8XK5XSKvGeTBHhFYv+B/mZOoAlKasOBJ4bWrU2bsKPA5466hFm8PlSZfWBekB
tbBQ8QsOwStCiIW5PDSrQVWdZmdAGRK3YjaBoLjgCvBwXQy8XSTzR+v/A0pGQXP0T8Ig70SfIFit
LIfoGm702MpbiIQ9/muqKoX9fxhrQVOUFleEP78W52jLTFA1hR1XPJEo2OMhH9zUnGPXQ7fFQURk
VQa21gL5mA89sJLyuJJjPnDIwxHl/n+3E0K+J/xCRiWA1t5if6VRo8h95CCjB1/Cww0pN2t9EXdz
c8BD0E09WhLAa8CIt/lDJVBKSCKZC+8MXlB/cN7EnsshCL4TLNtZXkMHhCd4ghej3olG0R1D7Lxq
LA+OhAjgQ7AgFLDsmunHYK4b3A/nBR9sUYnhbXrEwxVumCVjB6EjKHJiy9eXHCM7rDbAsbxQ9W+i
EXFPchCzChq/0n+3JgVV+iq2IsMsAbBHTIMXWrUP2eaRPsXxrVaW2XPvyr166Xo3NN91WGM9PEiY
MPg2G5fMefiLq3hjx0sPrHS6ssy5FCjN8ZnYnE8A7LIKRyJakzIb8vOiASNWpe/YVvoCgCNJKuPB
BGgKEVWOiLYFgRllo4PdorcIMNSBLojxXuWnTZYv0yUcGtAoBsIuCCvIl/LQEKndOWyDZamrB2Lh
YD6Wa3sPhT+vx/DFeOggOVnOK0gTwrm8YPXRr5Io5W1OIu6GJ64jcRk9HkIqBYHtsCssxaBGGiBK
5t2BwrcVn5dHWhR5PdhRcS9EuRlnzMIrCnN/1mvmQJQsi+AdbXhriPVmOuxE0uk3m2QOBvZRVny2
i5jndEc4HXtnZR8CEYLpZM7nE3EpKyO0K8uJBewGwCK0Lz985f6CF2IAR/opwIDNObleugYqAt0n
em0NlvJSxyOXjcnHdA5M8QolvOxjxW609/Svh9WVJPKy/HrG/laLzFIWEQgJhr8O7uD+k+t+6d5P
WKXFijnl3pfnNvYAM4td+vg5caZX3RMAGvgd+2opO8qRhjThXeEoFeixihcD6tscgPrqSKOJZdmi
tRYDHAshvFpLMa/GXyUAcTv/6D1i2YMX+qd+0ebb7sWtaCCD6a2XY9evSOpSEJDCYVRUdd+4iZ6N
GNDAGsiMgoMFfetYT0EEmSOY2rsv3/vR8IqLDq8hhF9IkZM+TT+hiHrsx1p2UXwWv46Ehd9Qxgpx
ZAkLEN/hZ9S1JoH0LCspYRkhHyuWS5LWL9r2ODoj76FOXsL10Yt/LZdpRFUFzwJUouZf5VcLMGUu
jFUC+hKYwetLsnXYwgShzWk+4a2rkig441A2wxzrbUXQV4WcbuS/dY+y1ezXYfY8oocSL7RpoWIq
DQmU+nwGZI7SJQ3BZY/TWwWw3DO6GP2E7nNmdh8y5T6iMgRnFwg8qd2Fb17tsSIgPQ+IpxIuZY2w
5KHnV0QKTp6lDmmuGgSnUYrf3aX+BR5v6z8uJ5sKyozXD6GeEfXskFsZAbR0kq1boB1zCy3AmH/b
05i5hhjoBxw5hArvaon3u5Rc2SiCo6eKbRRIAJjP2lI8JxoT6zHAOyVjLWVS7V2Ugql/F4Sg1oON
05oqvr9YG0ouZXhuKGTQkEfl1M27+XXexhR1A6QhLy0od8o496qmvBfKW97ahbE0VgH+S2f1poKA
6ZEp4pyDdH7VB81f8l+OKUt7Fnx+gaoA0QLnCUwfCbgZvdFFkI446MSBmZkiQ0sL4nY0ypulmlvd
/e9K3z4U32c0Kp1xSV+J1pOkzg2eRsdzG+9lb+iz3O6Qar6+WhvxdB4oXmmNrWs87CaF63F+/YHf
rikG4OktJzmeFsC8WiMEhOOngyd33/Dr9Isn7frC4GQ9ryd0mrj4muj1Nb3FUV5+IchZmVPKn1E3
pBwCVSCMikY7/U3b20RCD0ttI/OeCIX8XB88atnkjaZ0lwAiIFWmR5s0Sl5L4dibBQlS61B2EDoO
U5M+glTS+/3gUW7m8fZHZAn4Gdkn+sV/tQB3yrz9AlGshW3U7KyQhhYp+ok9sxSnjf5SKcqqZ485
EK0daF4Xq2jRsrVhz7MTm1XUmS2zoa3koqol0vBx4RRcAbdTv9QAKX2ApnIXknbIgZH0LEUJk5qG
eqqK5tPAyeeITPEW0fYkXn/vcxJ2j//q39C6SlM48NeQ1XMH/bYr2CwaVJ1dbl8eoOIk99IAdVOQ
fp4CVT9OYec6ybfdJ0gEumfGoTpgMGI76ckcCI+1+1k0HHrmKHHc7JuTcFDzPdVy7qNhYn5QGYpR
QXPFcEUK50sQC8OwyCQyx8vj7slfSU3UMhhQdA1z6k3Yn6IbApTWO6dZ+T96lJYXkWcjVK/MGmgR
XWb+5k4ef414j6Y1A1aofTI8NotTIYx1PbibYXOhUDL/tzG33Btloi/fnG6ryIQ7jiDTkFh5dUuG
2LORTZNTGr594/N4dTNeZ2lRdqmluaJfBEpbdolUyM37nfbCPV+s0utyMx/hwim3/a15UHZPegpK
GKPCGhiBhKH+gBYNwOP3yZ1b8P3YwqjyuBJiMg90MS+o+m3fRKrTsUGsB4HgV/Z8a/VpCIa1IF76
77UVSUp40+DWsYvhGAgrqop8JS7mFsMmWj/Rziz9e/C/VAqDuvPzWgi9LIuxxDy9otcT8kLbXYaM
HJApAcVi5Zu4k6xLkzGblnUirBn8NQsLVn17oF0NHHZnTBxx57oo9KU2A9xBy7Uai2BQ/Mf24fDU
SvUN197X4xdaPK2Feui3SwFwru2hueZnTSpy+80Qt0jP2lfKDgsSk6r/8k7Il2VUz+B6E+XXVVmH
f5pjGIBmmJ+L7RrYd77tl5Auj4ZHzOouIbhYzWsQjwm4e5qXALL7Pl45XoRnai4RQCysfA68aZTU
V+n/QShV8aiBJXagdmEG3bjdbzxaOHRmXYZ1SIjYgAx208d7yE9OtKWIGNP0lDeG2dBgRleuET99
ATZkoLPJiyCBreHrXy3d0ESbs2W+/YZVEJx/H4HqsgWllyAoM+6cyWpvLyXR22y2veZG76py9QP8
poC4WqxncOvKOXboaJsVOXg5544LCaabr5MG/06p76ly+h5Yo5mgzrM8S5fhRYjsEWwM8OL1Nlot
tdE7VnqUwp95V/qP/bOrDsOi50RVNIrbUnILlVMGU8nOye/x2E5pW4pbdIe6ZN7WVPDbpQ5A+AAE
loHyaXkK5npD3Mb7xFydoBCfadX3WtLLbtvo5qMddk+BRuJdbvavRCWhEC6hNE2IJvXxYjKZmN2K
1B9GFXaOsE1zD6Dg4e1RTRygi1vKGvEkV+jjNn7QiNqBQ5aNVPa3IccWiiGAXZ8qAZCZCp2XWAhZ
6JRajqlvdW/SPfJIm8uiYvJ1ZF46cSbPVWKfncdxLKPwc93WF1kZD/oAYmDEES1FFyl8BNAO0gZu
mX2kPBx96AeDEIRFAq8RIffVwmIBXCIjUJdmSuR0UwR03wgi2VQEyZN4DUmSguGVJObb8x0IdkOm
VCBxl3ctBLF0lQLJYiyVnJV3ypArvI9vDSpJRtVuJGunYqB52SZ0bVuhaNcHsU+oa+dfI3ltmI8k
+Nvqls8ZT9xyN46/4QyrpWYzGU7QSk1VXHTtkNgnE4ZPIYELrj4YvL4A9+kk3wl3jluIfbMdeaRX
DeZRRAv5RlJxJHqRNHR3phqojMIiOtEuO1nf+GZF3DnWcYEpuCooj8X6cfJYBTyVid4qDdV8gR7H
wwiqwIMj1Z/xA5OXtPag8zu3FniaIaYnmjcAO/NoWz1cwlGyAM+hDAzyq/Zlr5Oh7c7pD8JTHcBc
+hLnIk+bpsxgtPSO33lYmiXrOFscMiF7fKpDoh5k7EfwJPI0Od/SHJPzAjEQWl7NuVNSLtUolzPM
eb6/Hhe+FVCBRfUzbOtvjoG8dH9IQ2xgs7APmCNuEeGb9g4Muv7UGAE1sY6GdvtWUIqGFG1lytXO
JWg4W4/L7uDFAfvzx8Mi7JDU1GA8z+rw3M6zbCgxVfpWrnlprxlb2tRb0o3O+9xRsJyfRJQBLOT7
giyp2DiPzYgjzRzmLuoau5alCYgtlOMbOvN2iMIOLFoVFx/LJXm54a6pbYxsOt2IlSou/RhiN0Ug
hGVqib42XRmXR/Uo6c6hdqunZtIvaYIL1wdpQaxLkMDCFPeU3WZorOnM4UvME5hb2d3MIRVz5/Rt
7L96k8r0yos2OsBA6p9KIGCzSCI0T5ybYk4Ruj4pZmk3c5GTzmaOUT5CcDQKv5OFRA9D6LUBjuk1
mm6sgAiTXLZzmqE4gPvK9/IFTHyflyXt13nt/VxdGNZHTVClFCp+H3Ob8GnTfD91MSRFvhxOtWQe
vsM0x3D3Zgc4HYC+k8MGe+DYkdghV2+bNoziJ9zTiiXAVtBp9KNuSF2duxKMIA76pnItXMoY3jJv
+wQ3lPrtG10KkzTeyMaHepy3oVtbl8qM5FiD2Uz6HMPsidqJFuf25TZI3v3hwKyMhP3XWhKI65qF
WNlzthBhoWt4ijOPSA97g2RA24XykbV2mq4Kx0xuGtCHtkedHhBiP1RWafHxrhZ/7E8LQOkw5OCr
F+mYK9zIK8t/ljPta69oGHzvywiF0IlIOvyCTgKoEtFPslXEDsu/vCNghlh+RVTZnm6+vkmAdtI0
cQj0iYAmoblQKfaBypE/6yKMHHGapkS+X/CNu382IhskjeorOSGh5neRTdJfo9OmsmbJ7GXpfghf
L3B9MF41N8lPy/9u7NnK0YUVf/Bwl3LzTEUC/u1KrpunIVdA7uSTTk21nzooVQ8Sskll8u/oEM6J
K0hkhn928Df2bs8wvRtTG5WUUGv4eGQC4gEV15zYitijCOdXRQ6Pspgfx77WUqHasZhvOyh1BiYd
xdDj7+nPHiTH+uvWy7HRqvakmaOh1kIBcsUy5zhrzt/3msYrcbb+39DpUgrXeXTzIQxqajs5COu8
GVypW/9Wr9e2PGR3ZuGf5+W6dzVUZhIBdn/uLgxnhXibkptrtaAksS5zOPKWn1Bs/S2nUF2+wqfZ
j5veLJgymRg2r11B9LquWJKLxUwsXGNop+Q8Khbj+p7kpEKrWlPOPQup91GjhFaEBo5l/PYtJ8fW
pfEic9HTu0FvPxmVsro22dXmiZWCPV+vb6c/u6p5fbFZtdTuoqroJGXKz2a/6T4gq4JBLCA0W+vj
JAmv61Fh2ULHum8yWLr0DM5wBrJn81rLGDRdDu6Z0Aw8rvFF8uOlrFL8/wHgU7zdCCBQATGJv6Px
L7YbquJZLE9RqW1etFe10RG7K/GHH+fKBX1f7B2ATbgwUD9HE7ipZM1PKJATLCxxzUhm5HsyTqQV
Kz9WqjgPRAolUqYQ+FCleCnkrF6enPnMryeHDTaLkvaX/a7aQgnJW8IaHmXWR7BSeZDe9jx7BdPL
urhSw+OxlnYsMlVXGPoumh97TILWVDo9moXtnUjJ2EHzQiYR2+6kHHVvE6VfJ9icECXbXm7VDo9t
0oDeutdaCuCPH/I2CnYngOmCDj6QEXN8DG0hiylgxKrOUennUV2p5YL6BABT6G4j1mtHgOdJtrge
S+fC+2yeAkeCz0gUC4TB6Tk2Op6/q/+3rXr0zEGiAkOdfYX2hus9Wk2ldmLerFMXIqXGvjJokFY7
EKzKf3pfBMMDMM8IfFik3H2uVZT0wjV8VUNOGj+6wvPQPKrf2IfYxovQD9xFiow6eQ0MlQyIn7uc
NJAvnSdscvofCh16nu4Unrapu/MHzIgWR49qFUTFr5LQ1VQZhG9OZmzl1QbkKelPup/tKO+Oj7/O
S4QCkh9VmijwPvPLMLIU8lRkzJa14XAxlNOpLQL7NJhXibApPpkVrMGE87g9KSluEp29LFXKCNHI
pTQenR2XjGgUtt4ZbbCn3+JyP/VSPXKWe8ZBB6X+3J201n72XHQJGKDQBsgz4YQPr7YGRfICGHEj
vMH+RLfG6Gz+ITlXpToWl4ns1uCXDpbNLgyB4Uu5yjVZW/YkmMozS41Bmh2aL+VEBsj0cqla9m1G
rKYx+PP7OPKgUnLWl+5z826YBia53UZOlZWP+UP9Kpvw6HqOS43J6/IGc8fAMxFPLh+V44PP6+bW
32dJ+yrBuDamcH0bNRILiS9yUl1FkckyaQ9AzF10gsQ03QMyoSTkjZo1pKS6TkkWPSzT9403kEUK
j6Y3BBD0rsSnlBJsu1nc+GarOnyFp6cZ2ymm3hmLlUqJK8UX6kLV+bYyijDUqPIFyvxeQRcvnONA
f7ZOY0Y66VBCpnalEOBNVn41I7QupJMCzKDRP2r6WymV2L+QNSjSGIeMA5qIBYCNW1HEOh1ezLrX
eIJl7FIiABSroNcilgjnXEXgwPQIzuOcKWA3rZ/WruWbUJKmEhVS2WlGUHMnDCfVKex07hIlTsHx
JGCeHkJDyF1qiXf/YRNtgAFFoztsG9exJYX3MDh4actgn8oFzGO1Q5+DplYk6XO2GbVZ7KJe30jl
QQmQk9rGY5wXs/BkDkoQ994hUVHSuibJdzDDFOme9Q0/pYPd88T+Y3PSfgG/YtZasRhLIaXmcrkh
HDNpHsO8xVP0hp1Fkvf+Gs7g7AM0OKJlZb4yVtxAKY0BeXAHlEa8lsmdGbz41XFA/cnbxsS+/Nqq
OWWLJeZK/4lXZ/51VQi2mmeMowZNWvuyegK4zvmmnaNck+B0CtQjRhAKLXZZ2eeJXdbWJ5LGM4A6
k9CZrE2kJUpEpWm3OiEwFvibLwU6F/5zE9OmhlfOFu+iOQRH6iNAs6Jj6YB0Pk2l77PPsea/IbNo
6+lmV6S4Hyj/C+nWAhq92lir0H4Xd60xNjPIFi3+7wldle04+jmpvkwPVU22WwWJZllez5PY9UXN
I5JwYn7YqhBouPNy0wO8oadhlhqzkhNC0Pv464pEP6swqA7pRKLzGbEucXiqZT9wB5agPEwiXlC9
vselRv4lwcg0cFFgfENmCwdmr/bxi76zEZ0lABtLsg3nedx6l9BusYGO35luDRBB10LeBtPgrlAl
l+zzINdnWqzDkHQszlR5pJPyieFUUvBcwBgDsY3OZhQjx9VJmr1RRMvX9tL+X0qnEr8FPaX10Zyb
cbAtWp++DQz55RWIs13V8uVMckBQoAmPNRbPDyR4A/VP275HYFnQmTIEypovRYiDtHHthpqSriBA
4IIWBEhr+HFXb9ys2byI7zUsYScqRQNkJKFJDUnCwIAolWKVz9tEryY7zRiaXP23lIno1sanrO9h
/Qa1I11/H5Rtm71SS5nvSl38QAZC15t2YST1jQYoKgHBxlHEyLYLPd+28DcWEANq+4JLn+U4tY3E
RlPIJJ139vm6quVlFDuOy4Zxbd7ixXGLNglA7MK9rVRG6mZVXnmd0O8gWvmnqwHXw3c1Rx7TFssS
5xK5IMppgIavPxYCttOGHupSEmASeEWR1SGlFyndceqYxvAQibB3vQIET/mSEn+KjWtt++hFtt+Y
TeXarYPQ3BSaAMMkd2HS5f3gmtSOCpt7DU2Rr/pQTEUfVFscDMEOhi+kJnJ5kpLbrMK8nwGn1s2g
ueKWefWHSuz0hltihxUK7lPY8K/HwF1T82n7SWATxHuSUaaRJGLfn1cOX4xKmpJGNbh71A9vrCSZ
vy+3QCRK3hpOQY8NZ4qNIT3/gDeQ3Na+0aDQumvimompy5WATpueVulrnNuXlAZe3f/1lBOAh4HU
79XUNH5PGaEgUaUbb7Psj67D3DhrzdaReInrf+E7rtJML6LaX5UwMoJIvb5dYsljPV5msRoPXBQc
ypEHa83PFeJtNhS0dFxGGSQ0JjC9ahVUh9ORRgM03Hq7+HVRaj/4JQBgE6ePG2RDM2OrTpgr8bDz
SzSoBzyeb83aMrm880b6n1O8/Lj05j9RrBcby3KOGYNeJLhKR/aPMsgyXAtna4SSGDOcZvVNIr1r
946pouyPvSLwDZlgTMyQXkqkSVHYYF52zwYiSADHZPC8UXJAL8V4ymRv4GC6hNujDQybedtKaP7V
Zwg8xuq/AepNu1kgdq/ZIOLreWHZujeR9iHFWEblN+2+5GdJPoJWzBzaO0VVMHHWP67iG/wel7uS
X2HYwXOjMNO5/gYhnTdmF/UbCdLbYYCtTLkc0qyU5AfIVzN3sZ1VE05dlKEIpuOACISLjXI3Fu9p
VxecAGyfm3djBhe/KReDBiS0fUa1r1ECsLDYykfbA/+eV0Elggxip8OimaeCWaNEpAsyr98dV5AG
F3wxxFQWx/BTRB1p0ue1y9NmgteUBxkb4PJL1KBjwdK14iwMQU9ttbo5zVGvZoXWVzdZ8gAIj9r1
0vyt/IxYteFAGwkAI3xRXlzMUKOwwS48wY675lzYhWrjWQDdpJeAIfoGsNM9StQ2I6jIFp6ESekT
wYFw62LtVbIwF1Z9wXnZOw4vTjNGfIohVDzY3fjCsf02nIn5HZ/qigXefalRySsahM+evXyYkv4R
Tq/sNlq+/Z0FcgeL8yGEs4MWR8oUdIojzlACbu4y52smfpKKoDavPe14ffxv0LIlkATvs20e5YBr
JAdlP4YUhTiE52h5rgDcxsuVvvAh2kLuc4i+X1apLKRdAPFPB/ZmaE0e5VYKGTGhJy0CiYcnU8cB
CkV8DCwNVBQBlA9vFBEG8KmmneZ6xz2j4f0sQ1VBcrmh91S3hSpSHrWhxB/z0+xGaZZgdyOZbfyH
N+LH825B4Z3E7LJVY7aOA2bqukQLkEomJJLH/sl8yzQYKmUkWc26hK+ZiT1duU9nug2SxAUUOyYC
s54f+sF7W2kx3UQfeaxPyAsuuB0TBhR0IG/7fpysnHM9AqnSnFskUA8i+wng6yptbhOhJCgAVmcM
A5GFcya0i3dtUxLo0RDaoeCOWp/7V78tAu8e7hWrUbj7mfVUmWwGzV32g9jApGuDyvp4rT+m2/AV
p1ht+AaS3NAY0oMgDnrBeXlqtnRCfwGDSpNYRUpJMIni2tlhZGhKudAfeHYhVakEhVLir4yNPulU
iwMRTSLhSppjZGCL5FKxvG9wj1qn/ndtJ6uQMSHPZBRtRI/1nHZKMVwcGX/c6S5Gng0kz0a/7CrC
R9wMTybCkSP8kh6NBDaTMAb7j7+oalid5N10QnuRVDXaztrOojvvN7/PqpQPnZVFalf9Dk5Nb/f2
xi4dxYOtvfLc4VZ8Dsqi0w6uqW7pyy50zQrKGbX1zYYnqizjqUPkckwUVoexqnPdPoe0nYzPLg1Z
8RYpchgy6UvXtgaf1QbmRtHHHo9GPPYlxOD+2mi7y8PVFCToVudPix+upKrnkAM1Ul40G5UscfUj
dOeyJEDKIQM+GcfcHhSPV2UJG9ciaLl1a853HjtBVEHNvMuqmBgEtz7ILNw4eZ+eSEWycXdeW+nh
2xSoK3zFTefyglE3A3zohALjbFsuhKOVJ7Dtdz0caDSZ+pVUVdC5WLLFu4XyjGJRGZfAZAOtOz/0
6dkDTRlwnjm11J9XqHFThaAuAcTKcfjbvuYmZNyRMNrn4sWtx5WQzN5ilUDAcY15U0XZDrXxai3I
/cWXiLoBcgTQPQsIJNZWeGWC2vF7tU+NQSAcJL0gIVjRvvBHTDk2ykoRsQDv2dLtIQ922k9W27vt
cGovH3LH18HBORM3nD9VxFOfhzDDpbbOqxY4Mk2w0HhnGZLPvY0b7FT5ScnCuyo7mfrG/lPBUOCf
CssQF+RoFXPTj8rjZqbRKSrYPzMmaBOtLtkcHHOEZhs06dfns4joLHj05g1UF5YKssMZVgr8I75c
eqVw1JNbUG+xsHVOLRFfJC4Cq7LUVxqhIcTghToq+k0ZtdFReNWf03rdMyXKU4jDXV5MEaE6IQZH
VjZ+CTeI3lLLNCMPdbdv3b8DHwcdR3Ee3VhZptK9dK4nMi1sbzvEI/zrjBMVr1yMiMFEooBPEUWb
iPiRo6OuBFd2wr8ZR4t3IK64wTwiGYi6AYH/qGNVEIdxwmUyaZnBh+FyQk4+hMtGqBsovtDXLWSz
3VbIRfZDc9fwwf/QL+vs1SFOJKizPwPI6agMK6o96UnZnyS3VhMV3u38KNCJuuJ6AKqdxGtZxAbU
vDraRGOsns4ACqlKxcBpZpbZ5z8wo8Aq6XVWgs5Q08pZRjzu1d6KR/02O77gs3qffFaqxF4f5uHq
WbR/cC3QYIhCb8XQuSOIv4tLo94Z816t/mRBM/BKovd22+m6xKiStvw9oDKDtn5ph/6m9JdiV7I8
Nd2CZkN6Bhnst/P6JPJKScrEbFwfJYeJHfe+rS6kNSELyGdriq2uPNfxZMwkxgDzrxHmgCdpBurS
e7ywM1dMSnXq4r/a2avYVQ/qeic3166/SQ50DK9ujpNZHEomJ+ZgdKYyoMMiCBSw5CXBzNcyZJy0
+SUAM+DL91vN70zuIZtQoijgYV3iqpENX+a1eTFFULlO1N6YQ0vQnGTXghs+gboUMxrc3q3MGKA0
cT02n+tQmd074pGfXGOClSLjW00VM4NLdTdthD+aes3QjBmyMJEPyoVDie/C9BXMoiJTMxTN6tvv
AJ36pw6OBIcSyri5bzG0aogtizEWNMoGtAQOHDq4Ite84tkmG0H7BktFK8XWqQ6IkOx4XthlOJHE
udHcnt7lol/F2hobNmNQDS6afG5mOkzwOj1MENgW1AWuBFx6GeAOizGV5YvKVKtlX8+kOJ0/FjvJ
lE1lebNd2xQhakYxbwE0FWVc0PBhCeG2X+KhjBaJVqcZaLeblZctkN+2pss/fI4AtDsPxikZq4Uf
vXNa9uetwgEb+Z4f1GdwCtgU1ARhzm8HO5hbOhv0YZ3WyTMAXttTYfVyLAs5KKZhfKLkTwE8zGFl
Lv0QZpC+PkhUEzPWIxNZlUD+ocPLMq4KyjYwkRtnBpRx6rvBbZdKRPypvwFq0azQS7C7v1GjtRS8
OcuC7eL2WTZJA+H0/3rpT+I0kbgLngqxADj4hUqpXfTqk8XYxEE7G/465p3Zyy8Le753OTeCqPoH
9q+K3YlGl4nhC6DNeHzmBWjD08PK51VGyVQgFpPzg5YvgAOK336XEGr8vVNA9R71qy0r2EfWw4Ks
gJWCQcIvVnC2hWU4txks3RUr28UCCUHBz+RWHql1a1D894d7g5N551Gw9V1N+cCksLsmxblOy++I
CkQChciWWIpJ5XOVHGHysBbQhqzIEo+OLa4HeNYJp+IWqldYAMOopzVkDTyCLBY9J3ekRzpUeo21
2dxhFVK4+cwwSA7K2DVTcbYdGP1IiOo81DrbQiiA3iVQsRJyZ7NNd37JUcQjYTKhN58IAk0qdsGl
9pYPTCiPHU5uL6LrSPDO9xn9Au3jd5zngh/NumazrW/vcuqr4UXcAncy3utZtAI8FgpI1eMZ1GjD
YqWG+NTcuQg6WoROKSPr1h/tFhaSZRkHA/BheA41V5WCNoOyg9sI3CBAghsjDJjC/hM/36bIyTpP
i3BpaqqDcR/bsSXEUxuBQqzzpqnt/ECIPOT/TO2RAMTfchmMmJ1EoCYPszJO1Z2rPfO+VHyc/IEA
LHiSrC1LuUGCWbT3FJaiotgvIdP8sNLFS0e9QTJpglNnKZ2IvLhJyCw8NDVvl4Y6JPilMR7OHzdu
nOWMKiXqUS2PwlPnIOt2Fzi4weGGAzN7WlHkJkoWlVqZ9UhJ8RZcA7P05uChvGAPrSgW7kHUZKLB
WJkBbG+P3I9vogKrVN2XEv7flosjh2CiOGt/u23tKabcpHnwVjtxaUsojvnXUbpO3scMefkTC1s8
mDA0Qz+zsxg8+suxaAxOXWcIZEPE+sgLhVHBSZRolwl1nha7h9HYTtU2LIbYhXp2311PPBG1Xg8t
eXBmYC8Ab61OxW5Y2anfplVcEr45fb+OR1oyoMEvyckbsuZYTtf0i86ObO7Fga8ne1YaohIpu0sy
V1TKZ3bssRaWMo/eiVgUu3vUnfFuZw5dMcDIiYDxdpSEKp/FpGk6dsrllaCVgH3HobE895HDFo07
C20rZZtDkA3f/eSFw1S525cHJKvDvfvwCpQ3v4GL3ZVHaKORtWGPJGnMNfCk79afpCC0b5nFlOe5
nNHUmWhILsDqBhvVdC0YqSv47EJfcMdLFh2NGGe61HgsFJBxhD/mNG5oI6HamFcyqoO7Rz8g8HMD
2+ANQTGxWLEE1OXow4q2j+UXZTGCn0DkQCZcO/MMtjBYYWa5VgpM97obwmmA/gVmBmxBk2c88hpL
ipwA0eGyLdW4L4K7HgH73gE4QEWv9M8b/grKa2smnStPo9c8BX3XY3qoPhfOCjZXq9HbusO0/WBg
PPTxxFdLHmIZCtRT4OibuSAjCo5jtPBTKcDqp1tjheR7DgL9lfntZng0FjIcM+D+DBF0KyLScWfS
csgJ88FT0kVgWywbaegOJqHSFOQ8X3j3QEzOvAT4TjMb9z8gqTY9V0ouwWuDkivfx8VuBY0iLe7w
EfNMB08sSjHKUSwtBj95PprxtQ704yMD6cuDzvZXUH4t8NO0pJ+K7OmOkCm4OcVkHP5jbRINPm9F
grx2o3Kt/WHMTkm5lAX+Ar54q3V+y4EQ/V151RvE2KCdTLBlxItYmQhAQUZWjOfRPUn5Ss2XiUqF
SIkOCPv/z/CCUmF3MqPRLDm1oQ5EwEFzlrI5GGL0PSQnpH8opTlcTBYltpB++1kwOALk+a9oob37
yAFZOCjdS5SCFMASteXMNEGmEXaNryOCX7YqBpFcchtlKYfX2WsoVdU//DA0EmaO1dhgqmqir06U
NIrYg2+Lpx4CbTtNO+ZE8Bxg8uIxPmCU0WCnqqByVtdIS+XPv7LnCCupv2qciv6Lf8rRKPQT6ZAY
PiuKgWxtSyUs3YcEotGC2EdeOmIbtPVvjYFsT5/KyYnRssqXDAplexQbBnvzaRzp93Zd9vo1be3C
248EuwA51ezjVN7uiNDjabceMDnqH2m6pqOtYG+1JY4DIbgqCPzQ3Whbw16HxE6j8nqKt+WUyZzO
ZSWthRBwXSp2pMFRCpZ/JzkfzvngfDX+gxOVH0MS4eMB/ur5Sc33rzTrP2Kmct7Gusr3r5oqVGtd
uxuyUtPtzIPJ81yZk191fL9IkE8HXgHVQMNHehnq3D6L4jgBM8reXk2yTWPSOniNb9bD6hk5l4nV
jIR20JDo8Q+7ipHfh+5seJoQfhyabp/dB6iszby9byYysksKYb4ImOZFudHtuAe57VfCMAGMKRoz
Qz2Ml7SzlkXoE/XqgPGJm4PVOijtHt/7FnHgcD+L8KRWhRnNkkSkXJGSCjZgu2H8Ux6W0zuKfAUV
G480sjtVZ8s2zrma5NnTM59ugap0N6OVMpQMF06iiy3qOIdCqPVGrJ3YBad88449nUVCCwJyB/N8
tSS8powPsTqbPdnXQBghUXjznDyDn9+8Ceokc9CVInpi6MgzHZkG38qu8Mnx2pWOBmDKoZKIclKo
u7WjTCWvkiBRkUDxRpcqzLHgSMrq+RscnhlIph0a35ohTUha7QmxxdD9c6h6HcJ3HQ7PHlp413vT
L/c4ookiRaCO/mcwmhfQq2sSnMwTXJASkNH2y1PHVKPQYCaWv+P1OJW1+IH4YnBzyfycoOTY5B+l
i4GAw33qT3nB0zZf5FDeQDMSoDURvO2r+4MmA21cPZaSgXisvVsmyoA7IyvyNEln1ktgD+3CsseY
RRY4EuM3YEk9kyeSFldvG/gfB2UbVw6taNIFDqAUNkdRTpi6e6itZ/QwTgRgkNvtqeWyql3uKAls
wWwD3dtGVAAPx4HY49Mq2i4SYpJP0jYGskx2HK8IklCV7jH/c3fa0NL7a1AbYSczjr8YR7FudxAf
/0/YDuN3R1MVeATp8OI/xdYgqL7nwvFnJzDaf9vjUqVAyv2FbtEu5Vj1ngvqGVZlht5KHN1jHTXI
k8pi/0CCc3k0lWHy51C2hhJDoo3SW3GJHKdxWAo6Hb+gaIIUZ+XPGNewDrXub7fQumvNZ8h2ox3b
jvscQhAHI8BDdb4U3SGbe2M28uVICLfrRSZhvvZIY4sDo2Nwse2aVi0obz5wPB2Y86yovHxE9A1e
j4FPMinQ+6VOzaM5sNZxO6MwUWAFpX15ATKZu+IHp9ITJmPbqd6xCXemlxpmTOaDdHSvr6CXdb2L
rjVK0Klz3jSc73BYUjXG+bgD8Ndxt7SrvP/AGrri6szyh/bbHsS8r0lRCeGzx+zof85bKHqysiMt
lEcfvwwfBA/7eMbplX9vrv5N+eDbfdqnfTGMhNJE26RlRtnaLXHEd4rf5RMqU1pgq9t1tenTqIZa
pCiPDseMaCgAiedI+SO0T2VRbTWDzFiE78/9uBWWGddFWp08qX0GhHGhBOPwA44VKrM5kHsAUOyk
r8548/B7cLBcHjQ1RjXLHxxfk/PqBfQPEiLwALQ4AgyuuSBZ/Eqt/YwkkNJ4KQXH5pSScc/6+s5L
Ym9W2pJx4TnaaXHkL8/ajfMlgBMPVpeEbDxmxcfruMzSVygtnEWm7IVxs0psGGz7dzOrNWfotwNE
Ukl3Hq9ayHLdgqw4aTcSdZe9c8cx9orOLEp/00m1MUj0Qqb07+vl/RFlbjh3pwIG2yPsuP75dYNp
gXkMTnCfKqKmiV7Dhy9I8v4K/AeaWkq3+pqIa7+MNsgDegQjdxT/I274/oY85Unbig+cdFA53ouc
iOlgViDS1Q1g9DCsK+6ydZ4d0sN3cYXZNNgZBdYPOILwuV1Kh+csghxpDsmkNo5mDXbM3iz2Hnj9
B8PZRzA/SjYq3aAWA4SBQpsQwolA4jCTohSYWTTyWkAd2Nh4eT9GIkVfe8LlWNTbLqc2NSffxpv0
hSKnJOnLc50Edn1qjwbqQCyGQRWRaVYWgF0YPx3E4q/wowe6/gb7e5+4zI9RMm4nMdfU5Sj4U7vF
PtBMcFQ2tt9VByACNJ0coQAH1m2d0NcVpspWCi5iEIK0u4JijF+rq9NTqn922255RZeSErHWL02h
W6vgWw8QyBTChGiPJUWti80t7MXsBxXB8J3DjLXlTSuqDquu79f1edN/7J0MvUhYiV3PMHFkUQCf
+QDJ7/GPRGA6cSAQYZsqjdBTIyEgBkv76OE/AamB+VLpLWq2IHrUoog+HZs+EokMoPhE7PGx+Rhu
bnJO9+3ZGBAxXizY5BcOwjEgVz3KPC7U5HfYKw31q4DLyj8Jjj8NP164NZSEg4lVULygGKx7f0i4
pY/xJf/NLbamyT+U1fqKJnEiRk7A77rUCZSbcugJuAQn7A0/x9LzbjuhHPUYa1KQPVnsLWfr1TQk
VSs8g+PROwJ5ZZohp3sETZ8YRDNtx1SCRUmpDOHjmTLOW6ZE5t5Eu1kcK9Wvsb7DG76ZGxzaydzi
+GgiBMM0YoYDXdN6m23ANYqWF74gs5grryWUmyulyMxWec/0B8iOze7gscLyAekMgo1J6Sf5+GqF
hJmC7Q73/DfGuZ/nKTlR24plp24p9ML+FjoxuesBGtwtVYZdys63hbP8xzq+nEzDX/tcVxGaN10A
QeulA+jYb+7lprD1e8RDTEfXT+jcqnhIGCqQj2nFns5rNi7YdOoF+jDQG/zKpf1G3ZbN+h0w2yab
YCnvaU1GVjOZOaH7emVclcg/+r5fBhi/gihyhP7+Wf9qmN/S3kGpApp62AjLRtpX7QUgwmpPuogu
Aj6lG3OZjAsgO/xiVANkIu1G/1k5KG69eVqaGcdjBdFtHF4o+C901LbW+wly9v43qADBWoIDxzfb
vpM/spzTOMaGJT7drtY7jW3dx1Pstg798dbC+oz0BHjKdUfz8O8ALcyLpD6EWVuU00SnVxdWPYL5
RBucSHyRMEqjrf7cHWML0SRTk8mzqF2BPSfERUQsnGpwkNHmaXM9pBoNrUplrFnIqNzKTeSSgCTu
TZNIWti9pUzsgKo4jsf5WFQdU+kf/KADWCw3MoDQ33btZ9qRl/xMyKxDvJUzhkJPJQ0Uwfvchnjy
MReCD83nBCmFzNaDARWFLbMxVQvXDRhpAttaQNJwa4E0EMVgZ/YVwtgMW/67j9Q8pG5ZqezaYbtW
bMT0MccMT2kE4PfzXueeCD2xvvQ8e29yjjx4S9eapcXStEsGRUlEePtPV+DimGAQesSuh7Q8lkVo
qee9weZzcVduScypZ96pGurCNwttKrYcbbTJAYDFuRLESH116UL/tsij3KlQlgQfAyWYghZwbL+/
hLwr9WI2h+He5ToFerSMjZDE72ViPV7VOQF3xyXEapDdhjOJPM+2fWeTeSZbKMuLzZnv5UCYhCHP
EKJZLGqnyvBKgr3ZtHcL6zDXVLWjKDtAoHVrBYK+ccwFSZP2n9R7v0DPHHhlGJ9yE0D5nVVsw9aq
P1sGu+D+42+EX7H0/fyHxDrcDBgTPOKG5Bn/GbKYtr7ybh62JMww74qreceFCzLVL3YniZaMQmzc
i9cw607XgExLWqz+yR1wP8EI++iJD5criJa4OnuFIT4h3VJ6u75Nim6WZ2dY/we4R4HGXcphjIpK
0tnC7XgyMy38xtAe84uvV1MnzmwFQJ1BEPJi7wzFu1pOI4IHPBe0pLYTR6VKEK9cgo60Q+Jb3p0R
Lp/+tp6gTC3WzuPi44I9qlmFZD0KCgK5d0i/a6dt/oV1VTSs2VFWiL036Rj/H4HSb+T66Y5wL4MH
wwGzP5XYgbPYoLnVXUszcwGUsLH/Zd70dwwq7HzB7XVUnZgZgTLusDNidZ0tqkF/+C4qOSIm0Nac
cyYFsZIgYUiWfsYl8aA/YeWYBnY4TD8ugT7gInkyfc73FlBinLDw94BE1w6xvIg/YK4jiKEDnK16
eDpgDsH8UgSIMlj+OvOu2SbZPOZsG17FTERfz47S/rhLPOmO5Sews2UAd8A1CUHt4XjiHsTyFwWj
A/3QnG/vlUCwOTwKSqh5tk+1B8uqFsW9H6sEEw88iSuFMLow75ZgcH2n6WooNxGMVkR1jYX11Okl
uIgxlZg9igze2yy2uuzudDIspvQC2o/dV0NEVR4GCNAAX5570wz23SKLVa1fCpx5mnN3fq3Cj499
Pw3WT5+4J5txXbDZXdbWkRBVdZJIY+MGzBF6QGjxjblQsSeksh1vTd1sw127cvNUqqQpW6qZq0GY
WU3noObD7XNE+I167CQxvOFg2byiTbnOsUm4+CuXlUHXe0hlwEgTLf+4vrgPp6MEu4j/n6hQwFJT
qvalX9hA03aMfQZUKM37PtByy+VZOvvehclH1SFDopQtJAtSDDLzofMf2SE3ms046uLWz0tlhA/D
8qIEKcT0Sj30wdeX7eyqbt17CL60WldroY5x9nJzlfaP2PFi/fspM9+NLCbnmRK13zUDJqKoOjuJ
bjy4K301fGahecx8Yz4dYMqp8L13/rTaortyN3Mdz/Ys4i7dto0JIYjpfhzT6GKukq7fedrTrFZu
IHGiaWf3ko5sSF2nig+Jwdq/dYfwHdDun8/EsfH/bqWqwtBcPxvWmrHb54B7WN4c6FY3IwDODJYU
aKReTc0ybMpZG52k9/kMEYIvPonP27dnqWXAB1OoEmCaaA/LpPKUjwEjSkKoUn2H0TaRhgXtudya
IF+yHHahv/nrlf+sWFOSvkuOUH2odgF7impEv+7EvyppJmAMnI3KfPd83tojktD/iIElf9W8sp9a
ZasTl8mLgNZoA0FfYoMu/qxe8rwyG1NArI0rIgzf0+GnPKqKFwZhHJVAyIdcRjabNzkm9oPprYdS
y+PqqYrl/ombHxQYkd1Mn4m34uS4Y9qCmDzUKQ7p241r4nyGGB31AJG217gjXCcWUztopLRtG51X
S95XbiOf3PMyk1DXJfEdpcrX3xAMaQHGBxFRSTrD2Ltdvhq4LHuW80+sKgjr65My9+31ugGFswX4
maCqZjvfpaQE6nqAsSKCwm6a4vTFSnZS8EU8n+EORAvc4k4L+tDiQw0MNE8W0ztKltAQ8cK1xqcL
LxdU+wgA/+kFEUT2tTQP9o5Ih643nZyVc5Hq1jwDJuiAAfkWPuhZObYnO/y2L2S7jqA330PhZlJN
TZmsGXDqQRrbkUtnKYLwHhQMGjA/i5uBs2W0mfjDTzVOlX4/3B6HGZzsghxdBlwqW84DuC0Z83fq
2nCrHmMCRWTe1gPP2H7MSvm1kad3to9/1wvyNv+YMGfhb/rSqGW/MRArgs7eTO8TwG7vL04Vyj8G
z9fRNoaajgnlivh+3WUv30J2Pkob9k6UNV6aOk/uGTx0zTiInvxlYqX0WzlOvXgXaLLkeVeTOa8W
7du+vbJ/6uy+m4I9Vc5YUIldQQ6WMWps61OKDIlUmBiYcpby543yXe682HPIdiNhE9wC20hBd+iO
WwIHAuSDblSfDuToa58eZhIUQv2iBqiCC23zovTkxGmQYNINOr7X422taw/6NZVO1KTGDBrzVzca
CyXFCZHUFOegTeC1pfoKYyKrSLHWrkkuHzPKtxc+el8QEyJm2iD02P0Uhcz4J9NDO/BPwsX9XiaL
4gM2Rxfz6ib2P+x/GMJJkhqxkCiz7kLxlNCHy4N4t7yiEIjt5dbsu21weNTt3jiYyzLGGBbteCss
6qMewlrGimkzk+5kK9LCoI6vyIOxZyNXtXeFxpHhN77MFsUJNRn/2j/gATlG8fBQ8zQHbJMem1qB
F8TJ5LO+NO2TD7XUdn/V0y7hSGHRsLuxyD6Dlz+6tGZCFC8j6EMwSDM0M8qBbFJYIZI7/sYcu6pm
6eglUSH0Cfb1E3gLssrZ1TMJUTC058COskN01Pk4XqlL/m8ezVxURfsCckvmGJlf2H5vSxNpYUEh
c+WartgkFF0DofOTbn2lT7pcMlp40DZaTYGE/FTwY0eb7I3y7iZ4BiOrIg71HEWURmeAKpNnldxm
12HFQMXDdneWQrXMiEHJJ/AcDDqDj834D97+WOgQLatnpLy2iu0Jf3e3+mkLgtX0R3vY1rhs9Efl
boGm1iv9PnmLZui1yoCbepfPKF5NhoKyzuaPq85JuobBgC9N0f1TEHA/qy2AWYUNWboAqwv2rV3+
RZo46Ucodl7TBjXIH+PXxM78uZKgOg5SQS6r4uJunxyVWG896TAT1Dsvo7CUy+rFTAvQgNsLwx15
2ASgjdg8/VqsZl1zrRo9YOnaXt8n7WqksrEI+/RPsHLg3bB7wSxuH0eiDkTJwQArScTWOahNOP2S
QsiIByqUR5a3tsRxLWNWO/KGR7qOJ2chZ2w/wLWZ+kaY08DdRWi882IaWfL5W3hFbN+F0XiS5FnD
4p3JH3ceCoZjYzmi0XC1z1/D+fL8qgn9q/W6oCiL6zyALFbHICFUoLq165TXHyCGstyUZsypLDE1
njwkKCt0qh1rIPcZKjRD5Q7Gxdwoei92VrkyjiUrLpEoKGUO7T6zMlepkGv97CZ8K52D6ysYahwt
DGkO4QqslC2gjcpWj2EWc891szbj0aWSrvVi75OoPAS/qxexp4mp4hqyOg9kw4OwR+/Mb1FIH4R0
o18KCBA9f5j/MMFCi7mq2xT3/su72e+MQjmtZ5rDLgXZ6VmYaXx264jyH+X2/R5J/kfwgfNA99Y6
K9EDRS+uQJppKS7oS/cueCc2GOrLPbQrnLfLnRmuql+0I1OyDvuSn4TmP6TajIYaalwHz7J6MOk6
gMGJroQuZTBltz5uSgIe6rCLnGW5A3mzI0nBjmDpL9dQKfvb5odfPmZzty7kb062BPSLXOl1h8Be
QGvbu+D1BFvrlv13js/oYlcyJj1n4gBsRCWhNPDMBsTHKXnMwZ6kionATowWxk00EqQOe9UyPq1g
zXlYqYUgCcFtWw0L5ZUgrZhkzIJFq6nCC8owNAyR0E03ixtb4hH+pNAL8Sc6ANXgXBQWvhFiKw5j
tBJPkZqh57fZ0zrQcfzkJf3KwxH6Yi7srhvvzZLMTBD21VNTI7J2zOT0XL4/ZnlY9op6MV1rxGoC
A20aVefaPYFaN//L1jNa8HW5WcXRCfPNXw5NN8jjbe5ks0TOLo2VBtKLqxgu43jhwbTDJj4mFEkB
pNM+k0Ptk2iaNWviUY9l8i3XC+Vsw9IHMtBzJgK6g3lMpNahso51Djw/Oh0rSF1xn3/BoT9PagPL
kABb27IcXRaDuIDiet7s2/1hMScCaAh2vbfW/qI1RXmsAKoOfKg6Uq4+Lylgg7vuu2Bb//s4OfUV
Yau9a30REYKyZRMuBUCNk1XQtpNsfogvDsJzFYOxYtGZvDsN1yQhr/ajumINwWps6BTw8/JtBFOd
nKZ+aMkLPmVV/AZxQIqgJfWl53H6qPHny5VCHwExoxZJNmtKaOrJXBALLvgqq4mA6y09M+Upa8ho
s9wYh3lNvRajWF1vLBa6mYmRYVhkec1PqutuR1B/oiQMTNWe8P6v9y4UB2V4o52aWOspTpuZP+gV
yAZSY3lWwEdg5G1yqMyJe4Afil9zVcsRQIcpu6eKwg+IDVgL4/A13b+nrJkVa+jj4Q3yqXIH1PsM
UVczZ0tra7pzcen67jCUKv0qvzALyj0gv7nWEXAwrFoxJvSkIWMg2GvuORMFSeeK5rXralwpTyRM
GWfYS4DzCpvRzLe8+uVhiJiucGJ90gRpqidybGmS/JW6BOUQ6cz/szMv5E/IVsyMMYIvgBQXVca9
3OXjVkQIn4zdGlOHiQsWTgnnd2pIv5TqjOxO9phHCpu3PiqQXfCpwl+EoXb/SGocL+3UOm9HwrcZ
wN/crnBhxgt1hxdnrwU4zBc8wD0fJS4vPKssr29884JfSuX2YEbQrFnxGC/uVpGE+jecaCBaq8z/
DDz9ABeWIZQ0bg/isNAngJHrNPo2kSVzFDH4kZNVpgDr+uTPj9ybPZsZLD68qCunhdItFVJ84Tm1
9Xv7dRFM+j2vWca24btCXiEpZy6Nd29YWlu6frlS14YXMv7KgTThMoljz6uecDpSewvpGeEH/m71
+8b4ErlwaHgbvD0eeuZRzxz+KhqTjanY0AZqrfuk7MmLkK+b9RphKMKArV5bn8BDKLUxxlDkc+N8
1BVtst1vRrm8jxr1kxWo4KQd+cdZpBPf+Uy7OHDRdnUA2NnRvRUjKXmZIIUiz7tohEjYlTkfksYn
LsxuKj+jCTfitcsamgegmb6ryOFpTUCe2BwKj/PHSWouvyu+OUO/oTRN1zHBN+VxnA+s64f87BET
dcjr2FD0o41/IvzTnFfSIdE2KWkBnBss7Ye8bvxOs3LbWgxKO4+YAlvlGeteqYd/3dB3BxpMBX2R
gvXnpodY+zcbukzLiJUEecKJWwuSJEd1UKp+gyFFXxLV/gfX/CqcrR5yG9N5lZgogeBENWlrbL4e
eck4G12N0exJ2MiGUSlZv7nfljJXVCNeW/oWnHfUjniQDWVHvugyVt6jag/LJQFzzguvB9GiTJA1
pImPfI15li3jdhf1Fm5445m+WJGUtkDM7nPwQe8Xs9Csk/O6bUaA0eX2Udpx/LoDSiu7ez7Y8Wsd
NBZ2OiQmkUr2z0ws3VlfuUXrzpM8ANkh5TnOhUYHihi2fmIsefLhQgHpr7cctlZyE8Tn/qoJcEkq
3/bdyy+sdMygendeBEyl0H45RZSfvDKjRr1a5wtFk31D/KIqBH4YDN4hEMCqe3e5u+NaIKhpSQcs
DqJGm6a+H+uDPuk2pQiFvuloR3n9pj3ueodNc9ME6cuAMMUAwn8AR7LbgoHT1HHX7rmDYBduKqaM
yAfsS4qNWzxaZ2hlGl/MtUu2EhK7ttJkYVliPToHhIiBkrZdEOE1cifi0Qv44aIELdEpLrgUl1kE
mZxvjOj0nSnwvIznLHOu2hHwQSyMaU9Nfoym6XP4NUSJIoCJ1AOHl+MyQkeEFMyL5DgVVoMm3u9w
65vKb81qX8OuqqV5FL2YnuBqCr6mimKxhEYKqwTqNP3+LRGUMmRlDqDlyF2XW/79JXN8feMlFZ36
gL6hwnLOCe0HVcbliEpTA0uWbunM0UKJPeBn02MhuznBy/nWwZ/jfZ9QK8D9yL0Pz68axDyKl5Ar
XzJpfeJCvYKaCsHHRU7Lj2lZ++Fv6WJzI6fZtZpwD8li0AhbqxzNbIS5AkztU0RDwM3EsDTxaIM5
ulkwA1ZFByJAD57yybXf2SbI6H9tSQXxBrC+l2Czxnwl6X04GOjuT0cu2MfWdrGbEt+HSvG/zCx+
h3Xt+yL3qIEI70ChqwjhrOmTvhlRD1iB1ZVBcw2evOgYWM6MtwJkqK5LkRQ1bxg0h6jZYYM+X6bS
pm09OMLqjRH6OiFAKM4LqIL4Dv4akjxilaPTRa06W/AxcDBvhUI4zyVSxLKLrG0i3+aNt4oZF+sK
i9Osk6pgl5wssjPUf3ZYQBGPn8BPkFDFwhjGc+ZIlTAwE8jlUZkKmGNVtLya2HeJb9prMS6GAoBr
SSIl4mrEoNRg4f1BVqprd88yjpxp0V66Ze5FEL1hXfprxK3ILD4ylAjWtwno9RHK01TDF11a1hYD
bTQ8Pejcit4TNK2ObPqMzcD4AC2kHWIMlqRv/004SdrBZlADC4VvxZJ9/TweFVCwmna5T7JS5yAC
Jloq+GDG/TxBDrnSS8dKp3LLBqdg++oCIEhZXDjpwHsuZmBxf9liFT6bBkE7Lcj8GJYD3DzuL4Zx
2drjZh0ddHMqV79ofUSqgQPEG24rG06PCpspD51foFnlwulde3PCfhswZom19dRGV13b5NP2Phaq
XUKE6E3/lN6RXl4ml5sMQrb6SL9ZzB7suDldqVmWUAetwMnF//3kixs/QgmV6kIfOGSz94ou0/fT
ndnmJTM+gIBS5sDKEtYBFJYUpmDW7iSNdEDZVTPcWKN9SVnl5srKtIsMWJ3BpDg+osvmqIhEk2bc
oGaAsud7CLg2r4oQ17xU8XNiZAVX5lDFHphk/wy4bMRhXOYxpEvualXy4WFj4OGMpzuQ0uFSNTD3
hvDYZSAiJ7NaikAATVLN3uhwmYEisoRekZ+fJl7ZztsDDV5HIMhTLdeNQ3DHMk3GEyntF70GGEeP
4dy3bBgrvS7V7c1TsW4k1MSZIDrE/uL++olUbB649YNI6wsDe5Hfyhi6qJ+3890B57xE2q86AzaS
j6X8ERW1ND67oCJByaFHTULIer9+5ulOR+BS1VcTD/h2aiduBThzifkJgELVUIYvOj3UtMC1aB9y
+SenOUOq8cj/ljbRI7DLFEQLXA8s/aX0QraDW3PKyIpBVXTA9JYjhoLsSOVdpYWmhtdBcUPzP028
ktrzFN13k3HLfsa04QcKCH8cX4ooUbg2E2EfK5vgj6ByZCRVKqI0Fm/jVWjwzEPwRBCKdW12Aiqq
ajcI+ov47jSOxO9U/Ajr3fMtUTa2sPLvpTMyHaUjv9NHivTf55HlbjsXGzRjs25yEt+GLLAwQkp1
h5a/m/FYvEv7S2tlcF8dYTrR+PqN9vDLt0KZUjzu7Hxn+2HyiiWJ8I9TteQ14DEB2/vEJFwu4Zwr
oimJqxGwXekr1F5zSUwUoKH3MMPwHMYu8fVbphJsAtvySlbLEO8uuVoGpyeN7wq5xaKZp+S8OPF9
Q/cEXOMqJVJa+kTfab1o346kY9ZJowsl8gOFUrYfqbuPa6BUGVXdJWtKluAzNG9yMnRmLwYOs2cx
ybwt00FiH7+C8cP23Gik522l9Zjsqgbv2bmbHyfmAlMMj/lsLwle93HfmNeCl0ow9tmmBDfDus8L
+1IbM58mLAp7Bc8s5/UjlwgaWjKNNCVNMUFNIcBe5M2ll6lALPcKEppgPbDm+LkSNs0zyxU1AStM
aJoCQMMVM24gNNTBXJ72b0Qm+4TtLZd5ksazYiSxfl8WITlX29lCh7G076jP2JJ/GZIkPCV70ovA
d0jTdpTNyIGQnyq2gRVu6vzI/fPTAvw9KSTP2SigqKQaJvLbvIRsWhmc9RDZvtFz31mEkh8GAAG1
Lil+58ssi/8Q0KYxcnvWaGMZa8LuGBEkXDG1NOjAncujLSexxAlqMcMzpR3GXs7YDRXFcdtd5FEx
lsmd7LGcG09KwIAM8fgOaaW/74U6RSyVEr8qIFY8U5Q+I1GZdv1bfTFQ0lP1UEKaXB9z8q59UuIq
o6tJ3v0lo8sRUKvKWDQKc36/3VFZ3p0KtunFCsOSlf8PfYgmYaZ8Wy7AAA67edKeRBOo/cqxSQEF
V58E/+fXPmtDq0GlWW3141ED88HuPnRnroiehoEVeSyoZsfhi/G2isjuTgPMljPsDnQNf2ZRFk0a
iH6guQmy2zwHvaGEYkwxhupkigI9ekZkqQt1HunMLHzYm7dM42tzS0zM7SXaMwunVxljc6wp+Yas
J1jxf1vfJqRbkXKFmW1OxpqLapkE/6AjxfsKxQ+21D9DFRO5hoeOG/cIVYtWxJLSz5Xxo9lTs/CX
LC7MT0Gf5rJQhy6xkdYt6PWTt3/OGoDmeHfTgMXv2HIw3RYdSsneeVlmg6gwnn+/9fIjAuwqpJlp
T/ftqB/IPOXYz3dthYicTLhavrkyuP76UKN/n6mc5P1UK8jaqu3euJ60h5gGqERVJWdmi1MwGh6b
/6yX6xhyKTLz9VRj+Optzl1Af0/0LJ0WcCB7NZUNtrfnSt9r3AC0ZgP7p+RdvB5FZ4VWz+b4sh22
sQp5yE/sDrxsO+g1HxigozKDbUA92AuJuUL91tMvI8tFNGhdhxWzxk+LZinM036nGxt0nD9eFPni
AGX5uU9uFj9OTAxXDgzw2rV7pLDPYbW4t6zmSQikeVorgU0mJOONj4+l3p70SnnhcV0A/8n0I6vv
SOgXoI3jz+FH5kAMk0i3jC1EEJiSTJT1K+iFtmogtSfGKMv76so/oNcUAj+XxYivv/T517teDJux
NYLPch2qvMoUd/RE6CuifzIpHxJ1Qbuy5sXFGh3oTPgfexNU2XuBmvyBrvrxxcwgK9OMPL+cdHHe
vZ2UhRqOYBqUqIbK0MO/97uIyfsy7zWVl4KGoL7vKx95l5ZvnpUGmsZtg1CsQJoydyEyS5N6NQS/
1Q50OkSjr+gn55F5H/OmI2RzkyeH+wyWDBQPg0m1q0SH+UMCSfza53sxZMbyprnX/KAZxf3SWzmr
U5JuZqeYMCvZT0xQV7NYY/sRk+GdmBBU8+UARk739hjKj2i+lNSJ1+2uGJcrl8zabyzaZt6galbL
ZrPZvDr3h62m26aUqcfHZy9KNESrJf8sRb+5QvkNIszkNZ7PB7wX/NMCKwdAZLptYBUFC4GkppjT
SIpP36SF9juEuc/nQk5BX2UK1dcGd6oqFkWRNnjbwKKm8NdFxhYu72n1FGtGmx30SRTVmreXkbar
X5+2H8DJnQy/yaqwZv67arMgtlmAjSO6kmWSWn7qm9DnZ0K/z1fGKE5rxGMxyMFCghprkuTrJSCF
kagTb4+j9oe4/DEHme2Fyr53G1Dh84PuflgVI8QxP/UYzBbGCIV+MqsOzS48VnGq8GjhA5YOegaY
c/e3q2N91PGpPaQJhIDxFqNBKWhsJ3aEDQTqFTVpnmgsFYynan8ZkNlWBT+OqJkzYLmwoB4dQq3M
i2S67fcBHo17Yn0ODjxADYaLC0iO56PVWerXpgaZXyRdznhFeevo2Q/34Ma24F7eGbk5Mp4vQW1+
WvD+Pqr+XXd/Pqatlo88wJVbeDYWnoKEEiU/uklWRUw7yt7g0eEycd/Fvg7GoywxLZyVqhBL8FDy
kGTiorfveGOTMoCXeWS/QMN8T5KS9VJLz/IvKKh87Tyd7pOBcLguXdd/EJzN3dqr7wRfv0tbKE6a
M0xBLtMZ0Ymd2zrEEf6pB3Ba7TBFtm2PR7JyKP1oKY8ipRs2YcGKG1dZ3EsEIlB7QfVFo+0UWmg+
Hx0cM3hab9wqnya+PJXiymjWIL9U2V75OVZhhb+6i9sqQ3sVqAgBuRkARAXfalV1h4H/L62yZp8T
8/FeZIEOxOyNo6GsCZZqSiC2qIwBl+0BLB1GZVYZ6ZXaDBgHR09I2dlm5voL0FMu94W/ChjXUwsB
GZa8+1ndxePOl/xKtovbe4/J1AVj9Vnf+iCbfOZJT0W6IwJ5zvuaQO6QRx31SmTEjKjtccAjJywP
/e6QxXJXUYvRT7UU1/ex8MijZTmUpS1rBJLn4aUo9BF/q1nwiY3wqLtycbqYEqkU4pn1HGI1bvrP
lhjmmI4pmbadUYdxtOXSkx7qLAYB2tH5WhDaAbSPD5CK/qtOardXI+pC3TzOvcqAGir69zSfNlQF
ELmVpW54Yxg5KcNoVfy8fMaGkx8XC9FaByNEkStF1c4ZMYvl3QhJC3nKiepZqpBEy/PXyrxIh3I/
0gjNaZyj+PUYKr+gvB2yt42rUpqM3q0E4Z1zkvOQAZTOXaVgdTwKRZSSRDFPOcZCDXkz/16rklAA
uBdqF1Y+5KvZTO2ph/4yH/9Twg/aAr0MfxxnbxB827IFJ5U5seo58yHn4lOri7ALHuRdxPHk7nYq
izVaP0ltozFJ/7zGO5bg3a8O0JV5dcXtU/vqs4ZiNQl9WjckSnF/HSYpkQeMriBItWb/ovpYTWrx
S1s2RFmiMIKhbZCzGPPXMqwQvROQmhL2wFpEwT8O82/uekL+CkC2h+nBzV8J1yVilO1wssrEAc4R
zeUU+KsBE1gvC4x4jxxCbaHIR2ojd7HZX6CC1Ai9uVE53Zqat2A2P1JtQ77YzlBo+l9wlIKP0kTi
HGg6w43iYRI0N8AdHJPSPYbrAP1z3soTkCT+w1vr14/a/16TYOhE6UzGlx0AyA7i9j2KYHguuZgH
SBAtWjE/uNF8f97qeFZtD1yuDxJ8Ep8CKv+cgmbssFOxjvImvRRdyRDMFy4tzEZUG//K19jccXJx
Jlnf6cDm9QmKsd8Yt2bFqMsBnQ8+Cve1bIrGYpFqn2ciro89EUlROHtua0fqbfHxDw4lKl7McYJp
9bvslT2VOFT0LeXEl/RpGiEAVfNH5kKB+d3wVrmQxYyq90uBKc0H3ByKiTZqlnknoto7AMVRiayn
r5NuENZhaUnhjKzeuX66EcAMO+c13QNo9DWboCKlGmeI4Gnvjw6kdYUap8sKnmXKbMX6Hjvx7ZqY
Py2YrOjFWFuSdEobyF5QCmCJa9HAy0dmNDeGP9DlYDccY68BPmSGWz3JWCQVX3c/MDU9XhP8EgEm
vtj2TMyyn7yiwNJzsYQOhElu9/HM79g51DkxZwZkeGS9H8jvCNnsw3ZRww5YHanrNNEPsKTVJXTt
PUCwjBU6kNIECVgBQ5TNajOfI5db79EcWbIXv446FWZZpDo50EnHDICrCXeh6Y0GAfPJKv63OBza
ajR+BKSAfns7ORvfuScGeM5GB7CCvOm3RvelAPzPLUiNZTjs4vkcIWQpFBGk4WojGrPV7Uo/ltfQ
gQROykyfRN1Nt8AlbuphB3oYRa8eNeX3PeGkDRxI4nyMiSyH5TEkIpMo0tVl4ONkIXzWY07juZ02
+TaU1G8xbcm+8tmLIJLa+FpKQwk7RAuPE6Igw3YhrIHckR54RmgoL1BZcdOsISwUsTkA3M5OmrUM
+v09cOUqTlk0jlUygADLfM3vvV0yPcYkR9YgDUwKD9Cf0JWpaIOQC5d1wi82DKiJmRExkA9LFEtF
bPzlybTCK1D9oYrdnTGtaWVP2IF1sjlw3542zosIvhZXKh2lSq7g48Po23EoaQZ73fI5cw3VPn0h
uXlfVNEpnzAatklVrtM5quqEHNqAStivCqokmqITpeTQa0ggqFLZMM553efTloY9dc7Co7JtXWgr
NzMsdukI25+7QVyO9h0PmLdpp69AfGlT7tMWk+Q77clSx2iXjltsRrrdfGI3n4q919N+VLurDhdy
g1f19/Kki+VpJe8H9P0m16waQdmPWBItMW11Gnn4d7Gs8vm4N36ue0604iPM5Ls71e3h0wTEh+5H
Qqjto1r0eDu1dI02I/6XfzhrnhXyfFOUupJ7fW8bLJDdat9aCtYYOzQKXcXHY3ZIqnuJZrNgX+rW
TvE/SgGUhJPgPYXVwq/aqwaxGn9hKzhx9jZqt3L/YjSl62LPIm9C4DDXiN/6N8WleAFv2HmmlAF2
W09DJau0Gcnl4pXICy3xld9F6vrzf3z/jyAgSnP31Wj+LLDhQ4j/Jp6p0oa9B0cy2Y3Gu2uk75su
YsOOCAWgJcYLXDNOj8TwNdJn1/B2IkVxmubi+yiWtuKZvmKuGwNpdq7p2JBnaKbbEZ4GmCY62uUS
+j8oi9zRm792CWhqQ/aLoO/yFy4bNyhDBEBHxwBTMfK/dbRz6SjVCJR5HpsiZ0EQ2HjB1AjTn0wC
ru065Wu1T14CEu9urpfatXAr3pYZfNq/bKmPxgVfoXLGGAD+H7DNFGe7UycHRSUOy5jwZl8dHIsy
+6o3qTf9UMdVGWOhup5jR+ZYnimIvW7MyhvIHRLKFwH6aWL5AKVcdxmyhmL+J56FRciYsDWCXJoI
5Tk/hDOlCfCE+OGMZXNV2B4G7nFFINWA9oSjzoftAxk/lA+NwqnjSg/fGfwtIi2F2KKAqVttYYCO
6NGL+w3xm01bOSUpj9NSqsGT07DWObHIPfICua6V9WvO8RnAPy7zR4apTq4EZfqjEPv3SLOYDDUi
ZsqQy4v1RAtr47Swo9qhc1Aq7Q/lJANhqcBp47ADUqkfS1ZkWCrBQmteWLAL7bZEbG5DPpiEwJ7G
UhlqYh157eQv10hPflFQCIJ3seMqK33SE3bqf1OptDpN8YiTEn3TxsyvDMV002ukRUiN/idK+y7j
AiOBYa7shrHdIqNrD1au3M6MDy/JMeUn0NhdeBKLoQCvcRIvYFvhB/PO0OdHR37UUOnEVPoXXCZR
10f1+MdZoCn+THqIDuVCyqI+tnQaD3ZtEuc5W/g6zPL0wfOzBudniO/qEo1J2qZ9HQze+lxzvSE5
QfuCDO01I8agkglqZOYZhwKfB4IVSX3gQknHedWWUGCWZorJ4xw7tqblWWweJTqZxHCUelIeiNgi
PFlyTbQB28A0NrCxhG1XcFqw+RdUoFtS3yVrgpnJ1nGtuw3/848/xeJxGKhLEkGwhwypzB7TDKvT
l8NJLuenqRWmelmsGHE2vttoofd1M66zCKNeOh19sBRLw8G2hN1SYL1jjg4ttNQs439+5DDLLwih
1q+Lyef3Xyfng7pRbejkIy6I58q0eyjIMErckycYTF38bowg691R/JLcebylLvhTduEJCFGUzh4i
faD3eAa3WaSSJjyGoC03XvEvcULPJXMLH7ZQu5oAtspKIAN1g9QunhRx8uV0TbvUD48zdANkw+qc
eNhmS3QCrqv1bsi6YLtlGp4FvOZ/N5b78Z7S08vD3j0nRy6Dw4Vy5rtxcYaHjnBfpwcbSy+3saKv
p+3xfD6CeqpNR2Te3eczApz6MyP6d0+hd2ie0JQ41Fwd7uAhd/XdoVUPy76epp+U0m0rw3P5f4kG
O/qO8S6LXCELqb8iRqpLcq8pk8sfsNUFHdy4P+cu90k+JkARzA7oFsuhN1CEXkBZ5pXkMz+aL8ur
fIRDWvGIt+52EoxT2ei6G5acugUBXu22HtSFHAKQbgOCTmQYc+goKh/UaNda7WQiHMwUpGD1hn99
9c51OvetTWZfGGHXS0qyxFK2E5iLm2OaxwODRxJH2i/gWltqOU4JLHeSnPSOUVYtgbXVg7KDtUzA
WL0ZYL3iQYC6i2V05IYHCd2HSIdBHUHA/SUz8bnZm9sJ9R0gSliThfFsFJ/MVzdNOZCORVRMtZtW
MJnMck3iV/FwdNHgSP6cgE/bVfD1XDOgMqU2KA/+SwNO0k6aSrDsFJUjyACjeTmOiDVVEiieU1wS
cR1YfO09EFS7cxVBSbtrgMqg3ymYp16m1gzGRofZVDd4DDgkU/ybrQiSUamnDm3ET6rbAKDqPVfL
m0gKNtG/6SEQSLjmhAW3hucRKn7Rp4y7+SLQJ9YVncsIry6POWqcv2lw0nkkEGHllWi8iYfTmZcj
cvAkcz6o6X1UhctoIbtCHgzl1Jar9M8MJiIEfKcSp4uGBHw+wga2WPvZwJ83R6NI4na0Gl8MBQDt
A7ylAk5gpo4ruQLXch5hIde9obnTll/5aJZUQ0kcAufv6SuoZuYmpibR3KbaX2qAsg9LPCu66PBg
i5otPrVMVZvbefH+W3t5g1ROv2yIYSPll6+qmWGXNgQnMJhNH11C7uYneqWQeLZZB2gBxeZl13na
lLowTYL5qcCg+1srjzrQAMVCCiQKey/1Wy53cC2ElxrA03bwcjfNGUO77jC9aEZO32ei4CP1IFoH
jWXnCBC6SGzjxSowTt365lpU9N48tFqaVblLTaESwo4dX+lIb0v900oRWNBMy6Pc4LLG90oz9snV
hsnw6yfip1qEIRapD6nndhLjFZLmx636yvsN6VHvHpZ7cABLa2UGZgRZMXJJfUJAJJbXZyk6qEsE
bRYi9MTyjQuYKNfgQEmZz/yJWwbmPSkxtif/Ws+70D/K3uxt7Y91FNK/itgpnQEZYm66OfMuesgw
y/X49thjy/4ArpwjJm1kFc+YPRPR+ZiSuC48tCmZZgGVRteVTpCHUsA0w1RfsLT34rqWLpVvm26R
e1dfzs9piMKEmZ1CM9zq/Jz0KizZ5BbBzUdS9gmy359MXFt3CDPeFedhc3OqZ7krC8gKnThWz8HV
uBCeHrDoV/Y2OER+6QYWc9XJOZ9Mfn3ZAoaKvOGqzpjABXJCHkWt22x+Qp6LVZsCz+Deb3e0e81r
RgkMkDTkBR7O3DvTN4W7F3CBttmPdBnsPdglYMk0AcsVZ2OIqJbcGebygwLvuHYYQZ9Pxcm4ozTp
wtrjVA0wXmynqqdVteB/8mMluVT+eml50OygbqCCGDezxnqvgzuVVhaI/EavYGDr/43ZYiJ0VqMA
vSiwplawgYTA6ZqR6sjm6a9mD5lKZNc0B6nMqpiLGPrXDO/2sNaKswZlFhJ6TcPIjALKtjByRdnT
PDAQDpzclRrpq4+fwDKCXkvQvNPmrBHwpqdvTv/tJc63ZfpSaHIbX2/e5bWo78VU9bxEbi2jdpEw
mARwATVQLn4HWUsVmDW90Wopi2AReF/DHyOiFvApu09zneniDrpHTZnZM+vxGAjdqZUDSV1jaYGq
/F3RdBahPSZWN02QtqjNp1sT8X4a0lGyVjzr/PaspW4I6Ix4LtzcMqLMvd+XmCpk8UVrAOlWjvG+
qhe5zt/gqS41uhgZ5+6g8iGPcEB2bUeLSl+wN01FdxKlg/kuJoCM42WSpHeerHUMwOJkzlUTdi/9
ka5qLWM0k7ie+SuZMnK3YrZng3LFsNRzfNBViDbWmV3NrzvOePc5SH9TP20+IedfwHZ/uikkChUr
ZPr9N3SrTXukwegxfws0HNl2swqy9qfJ8EF5Mp5/XmNrq5+1MGvhEu+M56fzktt6gcJ4mn3Rsl7l
PCyJ5Evoaq26ZNrNLl+9ZXtuWQP7un5nbX2ac7tWkCrP/dKFu0HQw+wDV2jF6Vk1GfXz1xEVNfKq
fz25Ks5cjd6y6CtalJJ8k3luTPf5gsfrKK+sEODyP66Em6EIethQijlkCsk8HGgaQDLSB7DE6Rx6
lJu1fWAOp4XyomKqj4HJenq++l9wBbcWn6jJg2P5IsRplFQeY9A9ozkTRT+Uy/W/v90+mRCgJiuP
ytA3Yzj/5VzCLMFj2MsESNAtyuYlHZexFqXm8NrC7I/HFpY9QF7cxmnnnndnspfwaI33dlgYeA42
QIYBmd07X/GWH5y9DsqWq7EYBoSVKR4Tv5UUi1QVgU2w0+bIhS16NC3DSKptqBE0t4FpX4cFqkl+
qPBIse1v9IhkDkM/91mFdZeRMbn7fBs/MH6ZNp5H8HYUWeggH1eEWSHd0U+95S7wRHSJUKTVI+um
uKuDau3Y2JBUoA49wGRvhw+foKWhTeXl/XTpNDGcQ8L/NmvqI9lJkea+UJ/kYuL+wtTeS7VkznK/
mwsQePrfE+nHA/LHiPJWp3LN8FaMtf8i9r+Ig1Zrp59a+beCM63IUopnF/v4pTzVsN0EaEYXLRGJ
vcQf9FrgGtuAYjonVUzYYVqQlmGH0hXn3h2rSQ9VcuKGS5Y/VfXE6uvRfO5AQ3UP5fE4JFt4Evfg
aiRkTq/7ffwVwdNcM7AY6kdhRg4Q4Txpsd2z+/68IFYp4w27kJr7s02u9YWxGoz5NDEnvEbNl8Sx
TlQiR1VI2vz50qms27+RcAeNcA68MCbMkn72fzY1+KtUd+u+38LRFyyg0tgOEAK4jP79DQ1JU+Fg
QUqfjb8eI6FqSoK6iCT/xolKSHX8FDI4EP0EIwSx+q1bwITarO9zxdoF9But4LV2qNgG0LnXEnQk
wHr+XKn63uAJn0FFbvfE5KgnBj7rSGiuqmsSQxiP5NDtYldxISv/Gy1LYZL5c2T4lclhi4EXLlo2
gKNljvpSq/sCXAwUsqr5uJVzyFcOEd1ajfbUdqWhNAlkCvwyV2OGPfA95fielAjpfEze4y2Dpa5e
Q8JVkfIgeaP37tpEO6RSsSSluS6mMOYIVA09qI8VG7bigiY6hE5xuOuXEHb/6Isz36SDocyjug9O
H+vSheazdTu9AEV2x2Y66AjWKTQFh4gN40fUkDKg5mZz606PrIYNufEM86kBJU0QmGUVBJWlsRLC
W5bRQhmKBjtuafxzlujNPi3a/SJTdzqc6JuY5DfuAHs5zcWInrBbFPfR2hDAlM/NtRA4VSce6cbC
B5XHpD7rDDSMP7SvhT11eUu6XzV/fGriAqCtROdNI82frRW1qPY8dZwiIVjgsPHH2miNgslMQo6a
LrE6WBFY7FYBoqx4TWlTsLtYK2mIyg8PCF13/5orS3NGRagacrbK+ITN30dgwZYcPvY5gQIggil2
BXcBGXr8kThSkytOsDo780BA5vwu6uceVTHjENYb28zN7rGfjIc5YmuILbggWyrSnBRL7biUl46I
BLUIqfpBObkJJrWHSbQmwdsruEYUCdGYpMj6xv1JBdYBsEsXDHePWj6XAwLcGd+VYmxEywNgeA3k
9xTqgItMsmXSxpYX8n+h/WvuNHLmKe3JK8luLUmoVS9Rdjp7Yc6YGVPzpwkIXjV+wLu0mlIPXZ7l
wQ1KxWa0zG6Z6kFJfbWPX2FtGtEjG2158tQ3D/72ZxSY0ZoD7cI0fwxNjp5aZwqhTgzGlz5JoxIR
s3C+i8WuMSfMMoRBfs9M4JIz5eKUYZ6kvvjeZH4DahHzk9PxIQIVfzRd5lBeLnst8A7HSETdEdDO
NjA5pSugyeOgNsp7xCm+0vTQWDI3HbI2K772WOKONlUWvLqjoApWLL5+Z20NXGGAfovdvqMqnri1
abuI48aLud2iyd6QaO8Na8eDYqIdANNfzAoFM3Lu2QyYazpvhTqT6skKJONW2nw7XGhj0wR4pFPO
Zri23EUAp86FqyDXJBtYO7UPsPuaA0TeqIDUvJa7nU+DDApAUklTLxzsq/J7zlwoWr5vFHUQQxKm
I/Qx8qRx2kJO7Q/TL2rHN3layYGmwa1TmxS+CclWh3IYlZquXIb+kGNke+bLNTAgE+m85us5d9MO
7vG7m4B58xNaDH/7tVGQja35rDnE8/AjDoWDHSqLLfrlX/LAtL++Ajk6n0U6szQdLjisRwpcEzQx
W49Xb38fXZSTmLUrou29YtAr3gffACvvQXG9Z1TfZmHvyjgLIf4yLFbwUxRL75eHt3lQi02hMqXy
BxpR8TA0+L5I+sKe116PLOL3LrBmmfxEMW7jYGydJGNZlCklJs8PnvFwRY8bFLL2MofdroU+lm0Q
cvjdErO3tQx0gGJmogPVrjYdw24MA3sC8d3hup8OvNAo7J5R4Q+U1opG+OcTw/gTNebVWePXFmrs
A4YgDRoEIGqgLFTpY25dENG8T8+Geefx6uEJvE55d6jIbPp4rOFxZYxZ9YFDQ9CO464Gyrme4vCH
4GPVRlzKeBsL8w5JOG5EksA5LliNAgzYFyf+EDgSKbgOY2wtvd6UZh9xVnSZbPYff96dq/eUlVOF
EYAFwb5mYpJYjnR75VE/OYDhj5RjgowWI8m+kdmNPyHdGE6+OSqbKGh9GonWfVq4DWOFd9t1PGb+
AiswSkEv7ReKGWsF9X3rfBburwFIEWmJ1kgQ6E2nGY591LLe08aZXGT2C6s2C3wTLmxBo/Mu5II8
Uqidx2f2Gf2GEuouSVK1VEghKcUK2iLBfb1FTlYfnosYGCZyai1klARrUHIiiRUQCY9Y1oPePWOe
aBS0d2rtei971SbIEUuitrBNg+/hFTCh7YIRffYnMcQ6VaXIzipC6J7cEvoGx3BpSMmRv+VeLUnq
DbgwsPY5L0Tnee3AffTJSOmnzi0lETcykOAdkhCGJQzazvf6dqRPsilTDgoj5Dpv7oArCahpImJO
cWHJQt/ymo8yhr56ueGEuuyyaVd5Ms5IWyg+j93QK7AQP/vhcYXxzxgyUPx/Os46d0DH2Vq+Nu5e
w+qk4RryQY1cWd+j8Eib99QCxjH5//dvGxXDwFIVo+ZkYoBzM8hAWinCxh0ehbkPTIsye1cXYWM1
BRdnoA2QfpXB4nYy9WC25t2Jf9jai4NTL1KKjW7BjWibKJRBl3HIWkwtzYHCGG2ABgAGbPBJ4+wM
/AAbx1AIVgu7n1wSlaacxrim/k6hTI9AxLZHWprM9REWkJahQHXLc1z/ANbTK/h9HuhtNlgswTDo
7XfY/HUa9ym6nmK8LDPegjY/dUKceRFV2TDG5nx+fBjgev6N2ffWBkHsmHw4mRXeWrdGnJJWx5j8
15/QCA8Xi6hJkkjO2XQbWpVV/POPV7xAECHOT5sY2qImZwpeTGqgpqJ0smBlDUDZN41ZeIDocAyE
VEJ9KNyB6PtIT0MSfpzbWti0XwUb4glFB11x4ksRTvazj/z5hWCdRWNcaeHzp7KYf5hx0v7OajN7
pLW4shalqleQYfJq4s5Yn6+6N9Nn1BKvEkdbMODZy9ZtSBw40Fo5KF70ouZtnsmat667BEfSKLKN
ag2bsDLTy0pv09zQAUOhG/a0Kv+ZYYIqG541Ra5nYjJczFiHigUY1cUBmi2i5bzdPcbrhfwFiQP/
N1qryBTU0kN0xMnhJN9NTJWCmiMfTPJUF33az5p8SejQrVEaoNQ5eWChbJawBL84tg2peFo0HHLs
kA7e5xSjG1HmE0xU+71k39CQjuNbqKsZ3HvgLyXPA9sYRnrxXgQ11xXp0KXE4mIaiACVHyDQjHUF
RlSBQIcuz1kkej1RBj9MQch7P4lMZYsVsNucPkcuHIEyuNgkzdaI8/DFhEzwGbCOYgDFl0F15966
4ZTXg2OP1exhpMDaneGcIiEWDhPwKvjVGGl2FEnd2pTOlf8fxE1kK7mqdIK/kg89aMydEwMU9Eql
zmOhiEWGWYEysSlDsZpEaLHCIRdcSM3xrNCW1+Mt7QUQF2pv4PMDG2cZIehQ1DdHLb/jtSPn9G/E
x1iELK6VQrUJiS2Yx4DqbRF1wfrL+anzvE0aaziW+Fdv/TdmE8LYLIKWsuWbC2meINv1Q+O+knpt
TOe0WuCz2D8mSgqsgzu0VMV16FzTQNoBHOO/qMNihiw5X4kVAD3T7ZjOs7nnU+4SzvYSS8PUzxfB
feOH2o9HNtiYPJz0dIvdZOU5yiK5W56t92ByxcC2KxKZng2F9o+RknqluxfP7TD/MgCEpm3ZDhk5
240JCMu8az2SEnbrnO2hlydyDl/cZSB7VAKAipoXAa4P0x+3Rq+8lJzlNBU6U5WmxKTfIgp5j4bI
pv/UDH294MJf/3iWoa4qUhUNK1W9Fes80KZovK3fKFQLNOwJo97NLkVBamxmgxlhurVjFtiB5ML4
4mQSuDm1ycHTufbSdCWJZfGNkdoizynMap6PZw++y/DSTkZ7gzczZ89OR9iwWiUun3I6i8b05LrM
JymbPUz322pAMzdalnm45NZU3AKkuMmpnv6lYXtfI6gGM0b9th282zAmQZI3OEs/VAHxI9gMmJ9B
TT+dg43FbXlsj52yDOjC+gLiQ2LIP/cdp+c60Cbp+pHuN0Dek2ntT+QoDrH3yvqX8bln0IaVE7da
/HDQUIpcGbhKz7sc5wedJTC4K5yg1/2cOnhPtG6Vh9XcKKO7o92d5o7mvUjnfq9At54k1g7ym7as
R4AG9w9zELTVRpTiMk/UKlKegnWccBLd7Iy4sVkce1V1mWsnNMf8SloVJTz/baXUlNdjr44Ozcus
ins4Y7IMpAfrcyJIb57nMiz9kXOurDA4QbOohkZtwDkLCpKd5XBfR9u8oCr4Vk29raINE1PGaglG
0RMCwfox1Spl3DKr4h9tEuMBow9LIKaSF9d4lalLupvlvQ9mV7pheNX+h4TE4saeTgpTfSnJ4XTG
3AL+JF8AI4355FjkmUP+SWOMjRm/MQwRSUkIVtjgt6OJDLTEioJITI0vSFmMlH1eKY57v5nQLDuB
PuMjaUbv/7es9qM+Y/sTDm2iXX0v7ZSeH1ErEsFyrO6smsWKGIhJXjyLd76fXFOoYPjtSOsfTMaS
+iICjfFVKxR4S7GaVWR/LylEAgVJHa9HJRtE7HdMqg9Na8Y8bXQM0cZw5fz+vWVJuSA8Ufak6+rC
iKIOvAFILhPEQrAfBnGEm7/ymKMHugFm90OnqxerM0dxs3F5S4nMh12ZoJWLWXZr+vY7YczDF5uw
YDF5LKlO4qpHOfjdL1Af8XceUaZIVDlo1nWi0pi+gaHeEpM9vKT1BHKWp94Gumkk0bmb0QnwYVzZ
Zfb1LLytHpbM3PMvjJqMKEuFswKfZL2a6O/NKxF4hRuBq0EICfmGY5WFo1O7HSWfAPFBND9rIrKN
X8oWXFdXjxSlxZBIEvselhDLfmyW/LGYlKyJkODFWfdsGbE//uuc9QhB5eHNgHJqLeYoTa9cqWZ+
KKaJ60haYNNjtdL1pqe4xjzfaoTGRdBVvSe67nR+2Y+p2kqZfgAOLIieLjm7XdBVymtHtEoDAcKG
88j4pKKYDBGG0L+DWDSu0sGg2nfBWBLGxM0x6ncu73f4GBfyiXhm+fFJE1V5/VvMXs31l9UJrk5H
hFDbXZT9QPLdl156+q2dOqtuqSn7vRfkRSw9U3/UAO5D0+GXhuy9Om6yjDWOofpKT76vhBU6WNRs
vow8HqoVjWkXO56BFj9dBWKiJm9jVgy2NAX9Z7WppTpIV+XLdexc1ieFlV7HE9cBZYlxLFzmQEqr
ZjBBjW22QZ5IL6h+/gEA+e2E9BvqhuArSRpKeRpNK2AnhR4tfySe9irQMa8RAPik3pD3sVPh1EHe
MojfczFxO9GJOgmdAlHm3TlvAZSMhBD/r1Q2+B+I6RbSmZUZxvnIbmJVqZmILJ2VJn3a//YP3IQf
mD+akc+LGGG/Xcto8ba7EMhQbBuWUq8Suh+qSuNJiTADrp+xOjqAEUoDdRujLkLMszJMfcTAQpRW
/1whs4AA58sDOUxqUNXyynX1mwWKAnSX4ezW9hEGTE+4/XAnwc/K+/QZOImZgWWgXHeNFdSLsWrU
oGxFhf7nlPIK41KcLGLQiHrlzQNUCl/pn1MAog46VwzJabgJATM5HViClqVaqbatHrHs+ieT3aUA
oWGTNhHKkw4w7vKn/Izhfcx+ovJWnju5rHPV2NJi/Q2ZICUlWT55XE1k2rgBG/8OahR3mlnyb2XF
uxvowla5/VdqXxxmoxtiMLi81wB5aJoPwkbBtf+Bv/LxwbK4P+8R5r5arTwJ564yEVVqVb6Rg/zE
GxasJvCx8eGVT/zjr6HPKHp7IBRlQgYJioQ/aSX89SpC2eAewsE0GDrJj1Ncef14RDA1HBRkq748
u7CM0+/j7yOFIxNdavsliq6vbMTKmwblAnCmP6aslDq0bMtf7sLirDV9LzBPNDYi9Cl7zlkXsMpm
bZ1yGHvAikkJqAS9Gu6lgCMl1eurzKWA2dbY/IYjW+IsFlY/G+lSun+75/HMUmCYEDGTng3u6fHq
pWx5aYIMl+R6yPFjy3g3hqMBnA8YgcrxgqVkp4rqq1Q/v9zOBHmS5OrGsSKhRcIYouaeJ1k7Girn
AQiK/faPHHP/LHDx0EImddougj8RcdX7PdrczV6MbrAtA0CQ8dPWdc6xaO2ce3BCqtwt8RbYCLA3
gv1GJr+ltLh9YxB9f9mBpuXS2P8E2jRQoJrW1ltxFSe4RhY3Kl8sLi29TgV7G7fpt89Ya1B1onnq
3L+bz9c31HRpZ7EdEdiI6XZgfnemh95uyBcKGbC6bdKflUTiK6jIOZ477T49G9hN9pyruN5C2HsR
WWmRx8sJ73F6m4FyI7r6wehDLcpeTf/wBYmNQmngq7Fvg8Jsl54yss6y4EkYr2NyE/vyVI19vrk6
lxvdfaopsLCvFWSB6IoXrxPpttISi7Dtk9xhy1iaBCpzeY3fM+T9a3GfRP0bB5rLIFxQhjLL79Yl
iLZiUG/BW4ssS3mgbxA4f+ABN8VapwQDnkjR12r9ZYQm9BiDpI/LxRgCMq4HCLlJUnBMWNWSDSNL
AVsrk1YWTGwUXnxD66t952V0o/P35OgoK0orotOjNM5ed0dXfBFWTnBCgApPqmXiIGzNFosEmqBJ
YR3TH+dWMsee0/kKRJzP2BTfJOON+6CgyfcqI/qzNGxeiqqO7F/jzlSp2AtXDY4qduaBaVcmyDNa
pEEeRSh4D3DjFXKQhxP/eytg/JjUfIVSpkqOvBB73gBuNx+Cn357RRve4hxYQkMbI+YSmTsa6fKc
Pyox8Lt+OAke/odym38koCcLmrWtnlUQWpDk3qPbkI5mzv0JGuESyJHyrjcT3KJVjUtW8LfJjOyt
US1/t4q1O7yUF2ZI2BTcZR57Xc4Tqb58U278RhDpTAVEQvB2LYA966GXBg4iSx3XMJFxpHy23VRC
ZaunNGs6Q8pNYRWDTs5+5/CWanE8xAb4C6NBxs37F70Gw78b1l/FQrPrMEU8uLWtsMyBHKqG5u29
Mf+uB6tzlm5ogr2gYAMOLbd7LFwsEXwZr80J+pzH5UM0adY6x0iSjmvigLncTx8nX6ov7FkIy2pw
lyARdxHJDpeKJ/OruP73lzbhUixh5szBVicIaFwmBChLeEKyXpxX2nAkPMn14zcJ6vaJE9SLLJNr
Z+XWx1e4565lGC5wVVKHNa26mEKW8p1Qhc2o30KxpDE0uohjnxOU5fLnGLCbXyiJfZ58dYiA+ctZ
uqFCmuvG6NfZi2cYhnPE5ZMXxhSD5ebpvvXDPkR9d8QimQ2GNFwAGhwPpv2cOtbQfMpPzs+4NJiY
LQYnMquc6lTwUx27lzPH4ZTIOWNfu5YGPAlDNr7Jqbu9XBqS4O2rd7G4mNcZw8vDqeJ4eM2qs7Ov
BnFXCEMGiNfAZwdaOGInOG7REfB5DeS5TbuOCSp7gypI2frcRfq7yj6U4sV0yclizfbmyDWuRZGr
btcvwh74t0E20aFlJFLZuUUj3YDiusgv7RDtI6UUmeUI7n4zmWTRcfsziQ51jjavsyOy3mgpFAX9
vUYAdTGKAUILB0i6YCGGEJrAOCfvRHSgru1kAzAfnB3m5lfrtY7yqqF/ufhUjQAL95Q3mZC1UQt+
P3X7iNUbD4HUmkYSv2I8HBzHRZ7vmrKGXyqeI+5Tscb/zg9QvxGBV2fv1wZMzK8eINTe9Mie1q98
SUlt39jhqiKiRQQIQwckfrJSCHkDjtQnKw9f1SuxWgffsjVrF4ssZk5bavD2bztjFVEH2TgzUpcz
vTknwW9LVFTkWL7XM0baxNWanpHRV6u5HDwFinn5TUfxuOPhDNdd+qNxv8M3zOkMKXSfq3dceBpL
OikvgVuFwWHb5lf6Pp6cz5jJDQloDZSyOYJI6RWtjbNJ8WrtylopkylStAh+KEkAcjyHdmRdsiL+
VazFVeeFFeW9s0dVUEjFgjYASIsgCmGHhMYE8BvcOj+7D2C9/oaQ84zpW4Mh6/aNku4u5yJGnymA
v/6f1XNKxUVZUJWLu4y3nWusLRDYl8AoYtrCLik3JxZSs0pQ2P9SubqvbgpyXHI1PNZaVB7iVaVV
NW0RScE1ZidF43yXI04XQBBVeu/YoEPXBvJuKoIzrIlSgOdvIzbyMpnA00JZtDOFz8amoohnFLW+
ZNWAG+wGpxdSx/1ZkTpCqeHPbk0K9SjBDvvP8wHdUvSMWCtxrsPixA4G7Sn2t6Anyk/6mESHcPT9
3GdwFX4ICWukCsrtDWKeQj1MmQbULIEBvjwohRUhTTGj0l6cnwgS7lEphxLgYMCTJed4SkeZslVN
GRtm1W+FOSQoaFDLTZd43tXkI5uXXQ+P+1AXvwpnFBh6/VZy4TfDNEDySk4QRd09ljVdjWELgYjy
vH/Ix/Dl6PXKO20AbuF54mYavjHSHxkSVRcc94fY+f+dSndEN5NPuHw9K1FnNpPo1P5WdToO8Qv4
oaAZ2OUE22sGmZ9lteeWf6glThXIMRXSY8R3ye4K7hybskWrU1UPg20AnGdOajmOXIWo5NBdBhxp
QkWNWVyMI54FqZ3kXYQmE0bIS7IDpKteT0192YdOq+tGRGnC8kb08CdQ1djlXwZLTn/rn3nb4kk8
R60U3kM+r2p4t/PQb5ICxxFaQm339iCoyquX0C3eZh8ijHHc9rTesvdDzJIuic4sk1Abmu6pkBCd
Og9nSSZycAD1N09wYKRc/GhbRmI7LW4psARhmjnJZeA9HenXKtVAJ3DLoq780doplpijrxfwyUFy
67LsI77jEiTK553XQJzaR72bjFmU/Pt0UM0cCT+30FVYoShLCu8iDgkg6KUD8u9CvQnqYlKMZK3k
YtyEgoD20wmw/rE/8roP5zj5nTJOrG7ttMin62km3gqTXvsGwtSI9VTE2PdPC5hX85to8nplYoX4
DVFyIQyKDwWCgjOduV/8QMcHeq9Hy56rGZDyF2YhBqbvdeK1EYR2zENutRy80xZjKkd1njShV+Mx
19g/DiDK32vf6fep6LZHURS5F7dXV4E5SbX6yDmQxOBoaz6U0xIsL43w8qGfTIfXO0oW6mSb+F7T
C5TvFFtguwSOPIOtTylzIVBhyPZVDkowRG5+DAMG5mvVYGGlBytRCJGCg+onN4z/fvG8+LiZQeq1
CiknELDPt+Rk9aKHfQu0AyjBvScjj28MwmfZDSPida2YduJBDZHi+L0f9UaA5Z7DFAckhKnLqs7p
Mi/nxdXeQGyNSnazrVPb32f2SgN8ipgzLsthz3mGTaYjbsQvYKkJtds9Jtapydm9h0U937YOD39V
+6ptC0fdbbbZE6OSeI9MEtwgFaNA0zEhLTpC++CzqcA5sQB5QOZUOWBr6K/Hi3ohbIr+MuMJquDb
dWhxtHs5dhGlPR2/UwoCExpTi8Shb9VCfheJchrXx8GULZzBOjO2G9aW6T5o4FnzNmOc/mdI7JWj
Z7+LwQ3845p10bUFg2HutEzX7xC6Yt2heB/mxcZLYqWl0zKDvc9Ab+0LrsDHT8GVc42B7mgtiiNM
C/vg56TQaKzAQHjbK/n+YeS3TZ80ADcjHmnODiF4iO9U0zj9CDv0MqoZ2jAuHxrx0v9Nmw0qT5VI
XoJAWtMK2HhLnzkKpbNUdmTppIw61TqWuEiqWPQ5KQzDsPbO6vvyBR8tbiRGkkKMBLhymWKUOTLN
fTjcH29+GqY1hddCFEs8seIPt43InGCY9u7koWC0OWO2lRFF7FfeLYuWAAWWxd7l+7jTCOX7VQeo
PRPPG+OJjHEjLAHxQF1UDD7uOFFEx/LpIzNIOjUSBYULD5UaKva53zUW/41HJ+U3ghnLEHo0f8E1
XQ3QZrw/CK+k0D2jkjqpErWJTvBjPKNVsfs6kFhUwIFqrKHYWISW8iAfUC/eZWVUj0+q8328jM8C
zXe/VfIBy5HOc3c9WL/KiPQCUl2FqZrG1YQ5QX8EL8VbeptZrBWjn4tK8dxIQT24gZvZWV7a2UK6
EuCsD8oD4r/aP14viZbG44+ZxIpGAXdogc978L86l96Z6W8dAq8mp2YWnmL8dzl8EFtHOb3OCp3h
wWT4evSvZ/oipKYYBcM1HAaLjiErPjsbYqANUlNbMD2+LAy1s63UhuCnO5F6Q9oAsOWRblzgiNuk
MnEemlzqdHaPh+n+RhyNdavofQnh45Qh3aQFcHQ5wLWgzaa0I/2pPrBxxfN3Nm2pvj0Q8Uh6Crro
J73ncCChPZ3mBYOCFYvyS9adXqedY6iMEtLkl/g+ODaGVC9hgkmmT/MWUmg8TEhMzcPmMHbaFn3X
HqV7tJnayYUbjSb8h9yqxeS0JRhnQVQT92DDvoJhfo01o52naeOJqGEmPDy4ffOZw9/sh4fTjEfz
728Shq+MzJehigUXi/2JDOO2+vG79c4wOvjVuVopfv+/K5Wbo0UiEGZD/m9EIddoCILIMA9OWSK4
TqZIfgZAe36RaP3YYhDDcmK59yg4RBoDHGqT57p6YCLPMiWqBBQkCINrk5efJDAacMav6hETQcyx
QdmdsM/tOj2v6a3cAlsTBRHDU8uqjlXxH8fpk65oQquAexhWzWl0hPi6Ts9qzNkQNr68pHzwYKG1
ZzsiGLcrzy+bgd+cVi0vo6huTYHH8GHJNF8tpX+pny8VwFEYYyHjvwLT8xNXQBYpS2acqijLRshs
SPb3E7LbuQEsWEq7cUjm9jResjthOGIlCv3yjWRCU7qWxtFTdMkCKgvTi2yUz+TkacVaesEP5Euc
6t4iVJ+bBPf1Zx0UsC7OYyL1x/FjKJmyiDnNJBiGnuYPyVOAlmWcX1klhT38SKiMfmg9Mq+9uC4U
PzDWLOZmXf74sbQKZSbfbuR7z9RVo0qWKYV99KJGwWHKRB7sfIwV2+LndRpm1YNbhYYWh01+GIaa
lRU0T4HQIYPlpBpVbzRit4Da/8tmDbTusnTEq0ackDvCvoSieYnhMNAss8N2B3yiVkIdNFGFqESt
x90K8N9CpTG/jRmgrZsoJ8MyH4KYRLROy6+Dhm1mxoMcjwAZ4uMcdcTlplm/8pB6CR53OrkvTA/I
Y4HHsgOOh4F1lQ7Sydpk4sFiqRjZVN3015u7QaSDgkJXgNGMUHVi5pIcK9h9c+6vsLfUC8pJMEjo
3Cf4zCXKbhwbVPKUhPZOTZCZnU6SN169fEENAm/jB6Y/LKqW75U6fh4ri0VZA5EjQFVxTswGmRa5
P6Wwu7/n6y3a/qb/cZaWAFM0T83TrlJHA5BZ05VUluIyhOl8HCT5MY+T9aAGoKVmtwcqff0pgzLM
drZJfmkd8djjvxTKsKBa2pT5Me4D8kX0Gms7uRlOzDOYhZUVPdiG9yVmA8ahBMolLs3M8HEkmYqr
Lq9L3BiS1je4kSHfs3OJxhNGFDdRFrYDKxozZdnrr0TC5jtFadO1M9wLTTGVlGMU4TopFWBEz51I
QOExABEckvFh8qw6D1T4D98dIY1HggQes4Gyg+DZT/74Ckx9qqiJ+MEXTdaaiMkjmrv5jVMuUUhV
2LXFOa9VUC3uwrjJzlir79sj25BHWJtnLxNrPcd2NAVNiSfvVOufWY/5XJQaQTZm1a9cgNMEpQWE
MtKL4ksCxWTJT29ZtPvamDM5ssdwdnKPZGPJwtPQNuRngzW1C9DwE0DLdO2OsI62z31Wp6bTQtBd
GVzhuCN/ELthfKN3XIw5QEUx+t0nYXSdmQ42A/yLGhVKQbOYWWrddYmD+H+aK5QXCo97NgnpBj3K
ALeYVNe0Ypgj8VJZG5Yc9V3hprA7TOTcqsf/hHFUNy5UXo/WJFxutsGDUBW24X8zxzGs1aqb2KoQ
oo+VXoUqwyaSNLw8MihTCyApahI1C/uN1y2f/InXIfB6I7pYUjsEsvM/K/r6fsGmW/r665AOPlMj
csnortrmCCehPNX3RPDX88HCkd0eSSvzYIuikz45zZf4WGcdkfiJ8WrlnmNMjG3Q+ZoTWsyc2hTJ
hmOoPrlMrWWjIak7RY1m2fVOTe9ShpxCNdqXyiueAVaobSHIHHCezsIrcbVeZy9Ros2UEtShr3+7
Kd0fSzkoylhuab+md+wTWiMajNpT8tvj4AcQUBTEAtkjgFF+tzfqyQOdKbCWtPU9JFsiPzqfCkpL
DeMndF8r6kQ4TlEt091rU3+Ozmq9eZVWQ/K7j/tq8StCHGYwUxzLOHC3nZQ3XBC95TUhZGvEtsf+
GeQtpB/NGHbiASYNjtd4VtJ16kWKRooDzYKACJ3OrCb2pZUBcr4MFQWhoc2bV3n9IaiyaNyq+9Bt
14vNSqMcOVh09i7pyxKuDpAsq0MG00gBRU/T1N2INIGsNxjElArhbbAzL6yl25JclbVb6ej6T5eO
K8wjGWsVsEatSvBj8Zyf+z/eXitS45QKnEdFoGYDRPuOpCQ4NVCx3VuWErypdqsnVq5GAOvorEsz
FSy/jG1JeQCefwc2tPTFWe0pta6TpLi+OFA9zd/HT5ue1WTkN+WEGBUPSDBuz6jJGuOwaObpUNO6
mfU4pysIjwpnYc/MrZwzl/oFC16St9LvZQVK90Oa7tNo3u4ocoAAELVZii3Cc4DWy+kb8AMPn0Ge
RnnJocPsXdchlztdZIfgJsOhwNi1advxx/CUo40V95TrvifDjw7zrH5+v8LPyg8wpLCRfP2vKaNv
mlIfx+Rw61FsuRWbGNH/XQAUUOk4R7UfjFUmHIIza2lSmTlajkW/nky6oDGvmXGVQYDBYcESKh4/
kxzEIOp4Tg6EwbkBBzvuHVlkGljUJH9YBdhNQgPwi6Sz9r9hbQZLvr2uHEQyk4fsWkqFggFP7R8k
6mf2gotf1old6PvlZCbuJ37w0UYCRSBvHnyM9qB+mC4V5NZIj6vM4AxU4alzTcf+OPmWJ08B1a8I
dHrVdsfXwgPEd2OL3wQKR+qywNL+AlHB6/3UQ8kzSXPHgspV+sS9opx7k3U3SQgWZW5kNUcKCu+G
Jzn93egXgXg972yT9RoTj0MAftpdGsJwoo5G/GOItELqOkgvA2bX8NRp/uIjzM3p9YTzUiW2Dy2/
tlRAgWcicB7gzbC0DFocGMihcrkiqdCM70CFKv7iez/hgezyJRPmGb/xQHX5++0lY7Tj4nrn/naf
nnmnOULviQWNiafvP1kWZ7GCnnpZREi8TzgAgPOXrP/v08dtujCfGM6aDbto7/ee1t3NKpDixjJ0
hDX4oj0iTJBwnwHrajpmyULV39NiIpXl/DzTAvZELmkl/59o5AxpzUp5AqWiZmQrlZGNkU7P1df2
B6kBlQZ1F3u0tNw8GBO+D9L0YInPmSsKE+dLBPEDt1/sXOygt5lYG/R0g4KtT23/MA352c8wT7Zp
ioo4PCFfc1LDZvsbpTd0GHuwkR/S4cNsPs5VbP1kBf/9algVYuDxpgC3tzAKfafYiDFmZRG/8F7n
Z1NHKtxN+DMBsvMFerzBtyjmNr52b4MWLSdHRDJzQa34SO+2gr6TgCmJew2AImF2y4a0oljFMppo
4pQ9MsEcEHwThMQpwpXqgAxoMvSnwi6VZksKfBHV3hxzSOVf5MM++4Fa+Qd6Sa7EKJlTT0TFIQPR
qm+qZPv/GogCEf3k5pHpDaBX7DMLvD2sDCvF2sOcHg7K4UVj8djwDYcsHZk05lmimEVYMrfvsxLf
LN8fIMfQEazi5ADv/uUGBGveK5PN4VSDAQZt9D+HjMZS6r6i7vlL0tSZn7fx8aylJ3OA1Mp8cUVf
nTTk5nAPvJ/DIrB5OFR4TXr4LAYgTIM7UlbIJWE9KZrwnPNUO/QVzVaASDjnRz5W+YqANoILpCEh
Os9WVemZQE7xaLWbnqxXbI0cSop6uB8esXQSAUYhURZo2zuCf1L0UhUfxh5dPEk1HEQvecV+//te
mT2qeVAW6dzcmJoDMKuYKKB7n1UIS8FZ+A+LRy8xtDIjLr/C/Vr9aWiUK+Dd11hQKXlGuJ+aVkwt
sB816IR5I3+G9rYhspBGki298/WiwJFBXut86PiwBkpQMFmz0Rtw53GDK0k7IgtcKxcWNODkOyAQ
4eVOaj4Yop2IWMtS35uf5A9fngXHdMZQ/xHWWq4m+kVfBWBqmeGA1RJoHfTE3R0d29I9QKGqYPRu
Th+k22HHJw3EFf+aXXzHsjN1SpgqzQvw2nPTXIA7ou7dy0Wp+6RacwhiW7ydeneY/nyn8+VXZrLT
JxRIjPx0/dJ5PQMaTq0aRCsEeEQIGA+S8kjSl1+aU78QZRuuDO+R+0gVyXlpLnlkjjrKxaQhbBEK
hcn3gV8RzaHOcn5yGHswEA9X1ZGCDnEN48AYQOai3yMlnrqGUyoMKGaaWgJ+zMsKjcs5nbZaXMjh
te65BbJzXDEj1QKQBKqWmDrwbWEqW1LYRCxh7olByWk92L/CieEbnfVnKLKPSnDW20gxVjVIG4Jl
dpcdBMnDFC3ymc+K6l1q+wxhzorpKwlpR9Y0BT1BgVmY5C0ZvVCrhog+F7JnB7GId5nGQDpOEWBM
aSnGtF9/leo7dSBcUPuaSLYZdmA2hw6TbIVc2IDnvVu0K/0SXR27mxEFgOWBoWjak5KPkm4LArua
3Tov5E32ngBn7Lo7e6xmig0n/TFfAvKQb5aVzE+pTZ1cWXDWcXDImIzQZZ+wmz71JTvgk+MMrhNN
xcqIpjCtRP2Oii1MUZ1vTHLv/BxTBvO8jVP8QUTubz7Ya+FHREoG3y7BqeIMPbAwMOJBT8Yr35MZ
zSYXSNrNccrwmi3S72vF7BmcGxHhfepJ6a6/csc/VsngRoYuEpeEL03U3dilT7HThBNrjC/RSoZo
J1FpgMfNyJZvvYQdQ8JlBBtGlNDCqyBU+9odm7SddMKmxc3CZAXSxhrCg8tXagiLGl6Daw3Je3oL
legFkOgcBkD4BKauwZimYn+fpr/blFfUr6gulHDZAWTiZFb5nGkYf1vm3kvu5MG1g9ncjAMEH8wG
+7pxAbcZfNaW/HCOqGHQg9heR2iT4jUj65EmGyF8hHhLBhJJh1MbGXI9+WDIFzyhb+JP8qc8LDs7
tTKDKx9NNIGA8KQe8SECe/8VVA7ztWIe8vZpOnDd8pYH5DbVURGaXM35IBZJkhinAUvzIIAthb7D
MzhOt0sHN0aZAL4Ta2gs31hQ7SOgAib5ofal5CGt6kKefZ29gBkaIFC6kA9or/LhspamvVDd0tHl
A35BE/sYVdgo8lXedTWdWccRVhNkXj5H3IhqxJ+034DEtRaLkahOqvStbWxsCPDGvUMcxmGoUCfs
zWySF5L8dzm1E2T/3buy1rbOsVj8z5rAz6QO6slJtjb3/0pTdnWWpCcKPViQIr+e9337KbM7Xd+Q
aaKfPjMszID8CUFn7ZYgaGTf4/VhOCs9Fv6PJ56f8Or+fWHJ+f3HqAV8wxzU4QK1JE2C6siRkdk/
f1G3jOJu85BGj8rj0Il+DP4HDk6ajh9+TVjef7Lj199H1Pwv3ZV0hVsGne7E5IvJJmPgPoC3c6es
txRiNMHg+ZNrQVOjqMkanoH4S7w8BuXJKb3mTn2b2QMl2Y/PUAvUu7X6w8Kx+dh/OJ0lEUNlgAzR
AbF/98GVCpjCRzemW08bnYtjWLAV6ED9PTesHby+t507EsTh0vRQZm2tZ7KR+epMEFcFY4TI+Y77
Uligy8rwkVrtt3Ghe8Am28Gao55aJvnPvez0RRIEMuu87PlvW00XS3WPn57KM4eU68N7sgveT8mL
O8DwsXVU+7gGqR5mM12qS7OP9TMTzrAI0JTLOAl3A0CD0M9Us2H8JA4jjPUEV/EzSM5oORoItl+J
lBpLscqEbAeJPH9JdrJ1l/+9jDNUnceW6aYhrtpA//ahhVvSfmoUGvJPEABpw8DN3Dxrmk6MxXrr
Gzx5UrXH9d6CtxN4WjGy+9byR5qnnRKr2TiqjUcH9AF1lbdbUeSpenFgs5Luty8v5wUOgE5lQVlG
Qtl4HR7kxXiewkCpkSuqMDxycRUqAEY8MTLhdk2EBbnyQ6an2nE65fXZARIPN6FrnDcl9pYDQJGv
SK4ydPwm1+XW6M3V1WyhLjpivlLosyeG6yjxHZnNL+2jZGL29+xdxEZCPrgzz1ZwMfuUZEg/7xby
P/fPdGOLVkDq9WGXNv824aK/fqcTI84gHqpfeMCfo5u3Ie7ATHdcxE1rxcy7ReumSBYyGiLjncf5
bSiTkYaRRf3ZunZKWhCzqO1caKmRtOcZdkFNSaur7YQq/qjtMdK1NSWDBaIbkCHnmf4JdZQK643Q
QBbGhNj7frVY4m6TUv99zDIqHzALieZ7WXGkaUOIXvetqSXuVSmc3Dtbp7G8PQQUjedic+TI+Og/
bL1VchovDXTb1tnzBNqHndHNv4TG7JtT/VfXHFg58hz2T2SFTI36xCTa6+uWDCdCTJapv8AVmhhJ
vyM5ZlGa2ZimQoqXGfoaxXfg9yGqwvfx/y8+jCUpqpENhzGNyZPfjN72CwFxlLY+j0KayiDhR5In
FTFMu+jh7oz2gSakuiEmkGkeaUbC/6IgK/343k7Z4aUnPgD4vsuUgz8Pc+IOXIgNM5qpj2BVBaG1
qd03Yemub2lL8iYncE+xJ2L+pvmf9MIcb6v656t6R3Vcs/5xloGNWOi2dTIxPMTem4hKEfmAIqDw
RCR3PzAHKToDzeZXryZSU1Hw4ez5U4BwfvQvr6Yf/8/qME/Kwmw7rzakDc2/QkYvkEE4QrQD5HUi
246Z8IkIQPMsmj30LVpiW+oSUG+On/Im4XOYi3zzWF0WRvjlQFIjuYFMGjId2OEV/FwtYCqkULpC
ZizH/LBUWhOs/rvhu2BU/XOHq4dp8wjSZD4dEzlqBM9TuVH/1gb8hpVWx2TbSYEUsAAuw6XarAz3
UFSNqlRjpjG7yFqx3QXhAZJwDTdkih/FxbCYTNU1NOAOHxWRjTstViuosJcnffzImhMAGnRZkCGU
X3yt8q4thG6i+qY77hjduv7C+LY+L+Y+j8x57WjTLeZWqZx+Xh9113SQ5xUFyMyQIOP/TZFkEwpK
ZrE/U8outLXt54EaSRaDlWm5uLMmcaWMBApwrxZ/QgX42/+YdZiZaH+HeEtd3f14cu/3p10w6kp1
A50PdhEQcX25JT4lN4zgm1B7FAdmSxYLu9vDLbG4gsFvStmWZ+ioYAA3o/1SB0YdCbji8k13IHFM
mCotAvhHHRzhcW/shUOlsdW1pvBrwWy699Gy0NHpb74XIfWqazCOH/APiw5gEp2ngCWJMFqIb0UX
3IxsDiZDi0QWsWSaz1dgaj2tcatzVrKDUMtellwO6OVzK3suWRp3DuhkxxjXgTZb0H0f3qoDcNvN
/2EaZ6Pv+p9t0c53gvKEzwCLjgRM6s4kTNbxi6WEyO8suqr1qNOJ76BLUUdL2YtsKfbSVtXn+Iiw
PwxUe0dRjthyK4gR30Ocn0+4nF/j4Iia1OziugWk/wWVC0fyebP+QEfbLpHudOIUiT2MnlE+0Bg7
lE3SfxF28OsZwAzZvWJopf/v0EC0nRzIs3SAFZtYVCc9NOIMv0V5kzOA1vW5Zr3cecHiuCHXBhUq
7zLLxLBCy/EC06QClAYNN8FbZpKG75ZfvHoELuhAKnxhohIRaE08wwnB/u0yNa9vjAYqgK8epDe6
Q/FuGdxr352BI7Pkvlf8f4U4JRECkCdWOEBaqz7BfRYzVI4bx90wTXrunL0UVHlGI4cWcv/xX1Jh
7Olr0ikIXlGlDzpoTWgMa1FSCCcEyDZ7o+K4SG+4syyXgy9IdNKtWe/VicBp9FImeGYdqwUf/VjY
ZaZl8q3AMllnRgBe+62DRyTkcE76/V9YcL6T+6XIY9Z1M79B/UGkIHU+2ftiPt4LUyTIroLMR7/z
dagJ9dl4wsN6EGlx5pnLsFrma4/+VN10/GWJWefCUS/8tHrcu5H7eouU46vU7m+3yd/PO9rXUj1c
hqr9fPJlXCTVgcS9g0yPoKXJP0xbJIRPDKYFO/kv7vgfmj0orfVEVYgJ5g8/iJ6udmYL7ogbeWLn
B0Ja61tdSNyY18OwuZyMQRb9phWHpRrirsBk8iRPe+CU9ZXqD2540Oh/86rUwbTbYiOEno1Ekowe
RN/tZmkVbdV58G4lbmBDmPL3OZCTli78/IroolXAGCH11eJiMSLfhh7/qToLkZ2wI4h/i0y0m+O4
xVXah+iQ2YDdSMX1+2pm9wHHEpYaSwtu9R2/PX6UccQrVXSDspNKPjBfQm57+oAjDM4nKNt4Eb9K
e3F3nTneQSRFGJE02bkD9ejyTCigwQD3ZG945DzC5GQnAk2l0IK+MQrXL9VWLsp/WKUlyFOG6GW5
LzoEdt7g4uRjf8h5qMLxI8KTP51u0B1nxA0z0YSea7JqIe6Zkbu146rdlyOvIt/16LQII/KfeXhh
wyB7xNNEhZ5xXFoIZoULaj+Kzh55TtZE7Ehu56Ek3ZkYm7dvhs1fdCHKWeYG7v4GVyOOcHFVezJp
iGJfwo+ir1zrMisg4TowDUdSGneqKdFTvjmk80R6UluC65a3vu22LYURE3vSc7dchskvPy5XqsQG
2fh6DWQG8BihsYbxDtm22ngBikjMaaOoLkQpNS5pjDfUloPmrfIy3QWt8o0VxI4hLu/oCAkv902u
Ru0H7UJRNqRYxoKdfdajKAqO+s+T9Oi25V5hblqLiP5zManaaw6R2ppXN45nqom9A0HKDRVn7ZoP
rGnorK6F9YcVHxEKQ9cC4xsvg8NP9hC5nCcK4WIrA6jbFsVlD7oZfnvg1QRBjI2kAX2cTMT1PpcJ
kKqw2G1lgwwy9o88v7nvCOFkJC89fzTWDCncTw1M4yLsGJu8mDBhxm1ipb5zRK58NL8sjnOEW306
rEu4KhaIRfIuUfWg1c9+cAZCbt7K3A+ZfWLKKCouNu5MVNOa55tdc604QJYbP5Pi0j3Q12uOuRM4
yvVpGqdZAnuVTDtxlxfD20IfBOKHCDAuf6+M5C5TlKANCfMoygvvGxCcb2WjHp2hQ55CdUjNlXOT
Emgkv0vZfcg6hBFOSRokQqJUvkjGnYblULr0oBGiuFpwiDwLpfdu/0JKuzKyDP/6zH6i7lmifmuu
YtWUDaJBTXhlz94D70/nAbDXxtaH50h7PIGBDdrq8gO8BKAGOtEZCAMmWP15BotunoOxV+KL/pFa
7sRouspe+jTOxTO6UfsFKJPTT9saHKrQ0L7Nb45itcHZ43ypPJIlSHi6ChHd7osqTA5GnhG24mGM
lAWHJ0nX7Na5DGHSVHZ+ByJdUTCEmgubx/daDq3IK9TSnfAuFp7HoQeJTEk6bLs7JkTB4kQcI3vt
B9DpYNJ/5OGbBoB1kP/6fmOBz5k+eVipk37HI8JUP+w/5LrOg6Ww4/czkY+U1pJc+pabRkXknemt
uWZelXHhB1mwiAH5WibWzh2mYpPIqz8ZkXfyYzse0KEZq/c0s7zwYusJJuth5RBB2bMgVL0SceJ2
WftYGOwwwuTbyyrEvFutjL5v0222s2ogL4AicS4cpDrm+NH9nbHBfvbAdK/dHexrVcQ5mmbfCTcC
9k3qB9SkSaHna/BcEKV2NZEgQAQGkkQE7u6ASj+ZNWlN1mzFxmiP6CJA9xBrqxDPAQLXuTv4JF7m
cvddXN7oETTPK4sga8TU9YjxBFftPD7Gbhi5SMEhBL5GtQeyO5HC6u7IrCK8y0TmUKVCrHh3vvrz
meVw96Ve7FB1EVjMctQsbwtoW4R5GxgF3yELzfLj4HCvIwFX0j+epzy1VSphXMCzCUb/9R7S9rVt
K1SWATPSd5HLUZD2AFcgItYOVLYQyG3y9Cn8pBDSmSVWoTMGbigtGWgqYQvPy2j0yoL6KRtHeFKJ
ps4yZ0S2cW0SeexKcDDWRYWz0LkjpcjbjkI5I7KKqCEtSZNdtpGd4Gf2dEdmlQVA+lpqWw81ZLGF
OEZazM2GBGA7WRBoEcFfiZazTLqTsQx5DpjgPkGyKNMyuONS0ZTlXZPvKgJHJJUfRAhyQHnpMDa0
NFJd4EQygO8lC8o0mhrrBqA4bsvqR+4crq/NVT0vTJ/vQ7/A2J7hNlzkRr+UUCaP17WaIqRzHNsQ
4wG5jFYcCLYl3J9gpIUFJDuF8R2qNA7MfZJl9Hly2DZWd/PXlQj7zp9hUlk/Rj/VfVdZXLbPSA21
ffI0o6z3uwUFhzDywmMuE6okSyKiJdwbgmxheC13Ln6iJHTHQwf/DkxOEOp5Y7i/TDGUsL6quvC0
Njr7ejq6kP4lZoYgog3b9V0RAgBjWMNgijTUwrRg/DjojJZZFyRm/nH4+lbY7mttjMeK0QJ8bk7K
isrN2Ph+VKdHDq1a8Nf19uGX9z/+3jCrFtuXa8i1R/gqjfc1H8/yaS9wl1IDlEbLHmGXPAGy4CdF
i2B1wPNpFXi08czTQF+nVndBcAD/t/tZJC8LXcGodRHRAgv69KawoB3znapHto76GlNMqgFG6MWQ
1WaDDgMW66xIihsWvPsyvWbq4XWMUqKfugJTbiB04OuzjeITEGXD2qa8CwSxm24yf7vyZJL7a+2j
RHYwSpWrEPPazTKNB/cV5Bcpeb5eZGu3O9ujDAIN8pXmHze0ekRWM+nPTYGFUuQDYPvEmPGaGzaO
ehugiQqemyAb5mDlZreGQrAmW0s7NRYaxyQiP/1BwsA6TotJTzIPwhCfdxdtWP4fwMPgpjDloqSu
AjeQWknrQndeam5aWVWYfLmhgNGINm9UxFYk5vUYmNWgEUSJq2s+w9HLB1tZry/+at2X3n7IP081
5Gk3y38g9w4ymGktAFuJ4DPm1H30kUceVjV3WTR+gOcaHxutJvI9knYfCYfMQSQSJsNbi2RyjUyB
ZBfi6MyyFwZHOxWkfeVAHxKpzZ260ZMijwhTefGhxKJc7mkPm/cy4/EqlN5+Ddk/CDhKKPGhWbi8
t92c3HFnGPqSB2tNM0tzhK3ZT7fL4O6xoyjVOa1bC7HJEouKA0YeuDPWiZvYzn7P5NXlxUd/idMg
f54rmQoIEWHJk9D+zETJQdEwMXlmK0PSfUdk51Lo8Ot2XPLNopFL1weNqUanUPw8tsStN1t7HqEx
8O2YeYixLwboR3KV8iHteB8mMtbqY/4p3v4pxB/3jcZaMja4I275Bfyjh812SMw8lL+mxU+0IbQ/
0R4fP2zbTomq721zh2mx05NlqgMtCVDUMwruLh4gnDusYXtCX8ebWvN5vkDPcu3niORturOnAdME
OgsNmODP8jBWl+SaZOh1sKl+TTimDpwQaAVoOZ1PAHntHjtC8NmM4GFaGbpGa1Sh5Yu6kimIRlhW
gpaIF8851qS2hQF7XUSCw/pwJJxjpb2S9T1HsILLEiNPB8F1T6z2n4GZ2Up7Mk+MVwas6MSLISSV
+ZVyj0UD40ALS4TXLBe8jssAWusTIYmP/Ux0dGr1WB0u/8rP9zYQ3B9tkCV8YO7d6JxifK3D3BxK
Ez2yWFo0sIAXt4C0pKb3BJrzZwZeepjJkDHPpaTLCdgtuQcT/oFni/FKn14TtQqQcJpcr0F83Bdl
ktpQZic+Sq/ojJFpKf2TFlsHaAZnG+GIq9fkBFOT93y+oBR3csydV+OkRA+shGL3IjB4wbhClyYs
+nW476v3EUAcLFRnqkpYIn2EKfu1NGJjOY4MHWF2dIn7eKnhHqSJ/cdrQ4YU+T1/c9znUPiDJm3w
74dL2fK7fDoi6cDIT73npvJEQNGTpfbRgG6T5vB9BtWqaL3vNUj/gUk6rFiQEF9ns79md6wLq9zN
18Ur+GMf8ir68dwOUYt5kzQQIgN7MTsbwWtrDF4GwD7dTl6wzhfh/pelWc8U8e9yhmo/P8W8sL3T
Lfl0WKvyC5Fs+soF2iHn/ewU9mJflXnHU3DMcyVpH3HG+XI94KnhX1+ZpraBz1d5Wxvh+HybOkaD
XVmCXhyslkxAWMlJ0nfAW0jp23r+0HfEe5dEMKvO3tNf0BlQfPLqACilAXEKTqIYlzmoEyGRMpBG
IrPMPyTjTT+xC2LSlpt3N/bG57yfbZrOrQlZOmgymItxagBDoairWf13VE6xEppeORnj/AxFomdR
oSA1ug0YdBEXQFasilz7q7nB6ekRpCk8rUVqSc/e1hmYC+p5g6l9iOfTFokaXif4XXQ4pCPtVxKl
8ZT6Ywft+Ob6smh7i2ottQKRO4+OnQhIKGc/7pR/eYYdrlfaGAj0Z+JxJV4uVI+LGtkMsIa6Sc+U
S7/ZocLuK7gSIT07CaxYOAi/T8L/bbunYSyakh1fKqwwtN49YENn1nbRLmqb+wh9jjwumNrtRcpI
JM5g19xjp7zluPiGfvn2078Lz3euLc6HeTJvKDD+bBqCUzqjOj2nXGaX4Cgzv7ypqQ6jrhweqbmn
4lFGXT6TyF60MuVmhE3uE1h5QLqRvlItU3DkEd5DNapXqnrAf1vSaduoPXrz/SSO8zE+K0aj+SBN
wgwxAZGY3ZP++UKCJ3xFBYA5nu68NN/Ih0ugugvJV/CcvzdBvLoRflZ+6z/bmd5wuqRk/1HYDnXq
22eIK9lW6mgPxddQovtUddcXZ0wvTBXrg7jcpbsb4w6nZRdqiNR9Jr1GfCJH/LHBDBLjyhOsdVGJ
Nf50hU4LEaS1+q/IhuVSABEbHfbxV5G4yMieyIjFMSn7r8JfuYhBKaQ//yeTbvx6aHEVBl79muyQ
sGikrl5gMxxtIdPra5Faz5nrd76qk+BpEJzNuj5rDApoASmru44ecbLKHVmrfGTQbL+ryKhUK7lF
rlF05+PGqHJjuTuVIKoV5edQ3SFOLelDS7CihEpRw+SQIQBN5TLHXz6xwun+BvutIfNuZjfRu3yx
U6gpVegsdLHAYSEFINVEJL4bT4fq3zQZyouGsK1RHR5pvpsvniTJCkP6yyWnnPcMuEoUh4yYjMTj
pPBSYQRW3Kn9IjX6+/sqin9Jiq+xm41t9vTNpzNjRXXIO7Upy/jJA8jzhJQqqMnGj2LU096Vlo1V
4uhljFTQTcwcWVPncC+ykRN3Du+lR50V1OkLUzvYxE36i7ESEqVP1dtj/yXUboFjjkQsowrrwwN8
HkYWWUtz0wBZKuCENnB48JseasbawQgxk3Lka9ahid+RF0/msL8kWadNWTV5Xu8UsBYuoyJIbz0M
p1zhFb4eaA4039Srp2kRyIwq9H9fKBCJOodU4GpVztwE7wWJGEp1SGE0iEwzqnLrfw3VYKZoN6Z1
iYKSnguay/oZgIgm08BI6A7VBNlgmrLYHNcPx1dZoxmThO7em+YFy12STn0gkpO9TFztkVTJm20C
xqax4HoQc25nmkLq5exXScteqs93G/LXULAAlJSFS20wk+Ke/NCIktbTz5+wzB0pA3UPyEOT+J4O
lBSWek28Ot0S4cRnorFay0CH6LxcVIE5npIGSp2TFUbxGipY++NBWD1gfNRMtZ3qqUKoGZugHl1E
6o63wwJ+kyw8ZNDLn9N0f9Zj+tyAZGkd516IrnlZ9HJW4TAVOYWL41jShvlDl7yPM9KpE9cneFIp
5RBLffIFapDDNGqXdmQ6rBy4FSj3qZmfAy4k+gEGS0FZA+wIUXNwMtOqUpPXVWWl1487yrl+Gkr4
rDNB1bLP5ALKixzug+lf+0z4NVJro7tdOXKvfBOjQs4LZU6SQjx5tpFKqg2wCoF/M3NYE8o0yl70
bXbAPtipU6qJP9yxQeHRP1KvJqu9IwOMhOzbtWXRKOq/wSatVhtk8atVjVH0SFuLEOYZNnQPk9Vb
jDRBah1NkCLzpppJEwHCxT/0qvOO0U7BJcflX0WyKBJ3WL8IQeR0lTH+H0uvHY9IZ8du5YucU7Us
+qvVAGi7BKf4dO7JnwBRItJ5wOpDVrbZAjjK4FRK4X8mEJQ87QxpV9IN8e3g9ZIg6t5htqhBjv16
3YuNT0w0hDE/nHFFhLeNVozxuLFcTpeVGKNVTLxCIefHoQuI6xXa1IpAnBO9ydceYEYIIlt/++g7
D/3W7ki5P/Oa1Wc/DtBq5a8S0k5GeCZRu1GlEd17BtWd4yU3GxqtLo3jVnMs4rQDton9Qiy7wuGx
wPUJIYSfj9D/5HQrEBdkld8h5i9VO3MVo57uhyDf/4TCxkuMoCNLB0XjYLpw039wlB5ezzNi2g8n
dhr8Im3P/HL3M7cY5LqC3FP5RDEir+9lF5lX+uOvAm2zyJo66j9FU+VefFVxTSXxH43ZtELaNN0Q
KN/ADX7jlLtoelik+Sb01Ysk6501ONrkiTPhRrmLikmeoZOTCf982WvtDJOd2FlHxRf7GHpo82Yj
zuNByxfjHceCANRA+miPZcPcVZD9sebe5p2Z8cUrNihiYNA+WssYgGJNHRBKJ7/uqMpiju5v2cfS
P62rRfTZgmpmErRAWlewANqVx9k7+G/vm+dYM7hmqE0gfAOqWProjWtVB8a+TTEDjXOzJfI5qMXI
2/Gb0WCpruupYKgPJ9qwuvGgROb7ibwo2WZEa1cCAKG4fktsBzJRtq6yT+0wVAvE3k39ujdnmGJR
lwPeP1rHny28reu1Vors1CtpR3S364XYxH5iXOTfbvTfm+txM8cPWLmlgFQcv+ijwkVJ1pFRSLMw
nGbCYqNjL/0vkCCX1A6HCYEUori6b6KOH70P6ilKmUykLsxPRPTfH4Z7dufsWVrlK/jbSK4zfhHQ
ejSVKgO3l0LP0yVXC/9k+s7kJ8Sq9r17Y9hjNVNQtSGzrwNjx8r+7bI2ThbJ3MQaV8ZOD/oQ7l0J
cFR8TpNC6zMwPClXLSI1GzmYYGsUki7sF9M0UhvmIVzblJz0omqBh55TSlCgUV5h8QLdMvD35Nks
um3s6WX4MriuF/E51I7t4w0R6EN2X3W9WnoDDf0mGEPB7rJE3HQelPJoFWNfVmzM5Q2BvfctFbbI
H7tr3TYSGqS4H6pi7Fjvzo7kRdmysjstQgujgJuynYcswo5027uw+A8e2n7RNvUatDoqo3S7Ugbe
ckwHSdhljeEiRUaFR5WaGQFXzIaNQAJE6jxYh8efcjxlf7/c2c68md3gZsyqnFSPwkRcMeNXlDXZ
Qjn6lEHjndGm/P/yq3XU+CvmQpYTQZ2rPsfmMqbNWvjqMJWM2ia88GWzmC+2d/J/wA7UVSe/jRUz
hNIaMV5vFOc5s4ZMERhnPyDGOIG6uhAXUgZ9dLe9cRH7CWK/K/pbe6GA0/qXx9P/TiEE+Tag6Ed/
U4IFVng36w8d17xoLdizjUZF5UaTQg9WQ26zMSpNygzz+ysaXeHnN63fImp3r9Vpo5HWip5C95rI
A81xYndZpgqgUmwP/nCmbkesJ72YzK43NsJFbpIQ55l6C9NkxFgmJdRw+xXSZYhRJr3i+UL28GE5
yXku1dpPvhQA3dqs3KB8cTaTuC6UGIQuTIUIJ2fowy2BZLB8TgCaAxB1oAcg4HUyB97FTk4I55gW
8iAcQTTNtGZiW4J5cFFeU9Qq9KOMytjz9Zp0KDsgs34bcshTTfR5Bv9xNwsJYHdC3JRqdqEiSpjw
JkympEILpRMq4MCVqjjftWTeiq/Snr8WczpTyMgIvSVIa51fgxD3ytjIOyRqszNpoVxXc1GDT79v
OSqy1+8spUs5a1olfGmAdlxq0+POf+ZSTQv3J9q8bKw46tNwNGA/eVC9JNoeAN3ec87EaVtIRYxH
3dW7ZwaT23RjwpONZq5w0bS+BcVBB3UjVucw+neHsqZhCwXeB7jhUlmqSo6qYH3Rsb0iM3Qj27ea
2R8/816kMHrVhQpLMMmrbBtv0SCms+qrhY9DZt5bsnC24Oqgl0BT1shIk/+TRNsx/NdGmPMdqEAT
aUg+KmGSnS4bFL1mL1LvbXXujbqqw05DqlfFXTeptgPwY8tuskh91mEoW34f57vngG34qh9a/Ty9
NAf87kR51X2LTBzA9F7xJ8Yg83XO7oXlFUkUd47iqKeKd6mT3k1iWKuPG2HxXfyapkcsRVO0BC8Y
58k4jSDBoaEyG1hAlt4kQcs3NAsXjH50d3JCCYrQs38j7kwMfJiyNK8XDgp+RsrhmhWelUBtFVoa
JrGYo7UCYVxzkjvl1+RrNyeBeQlsL7cZMiPAqOSqcKFLrpvHj3PLkPspS76RNleta2tzVNBKQmpQ
8MA3H7DdnlwJJgJraMIoRR3+9OWP2i04D/E/VxGa5QlDlqkh0dznPSJqVy0DdOE7TD7ZoZ0ssUVu
BsabClwo+YcFKc52HRNlnpQlbRPlBrA3xzs9VFiQMMRxBijieQMPJSPNKiO2klmyLSdpkvUPO6zP
W36mEA8zj7FisUAF5R9Q2J3uvKM9nHq7Pw1F1U0GflHwUzl6mQvHabD3IY/40VRhDojq5IQn96Mw
1bCP9OX5ZxLhHUK2Y7MowhQpJNu9fnvFu0PZ68TPncvA64UPIRE4fx22lhFVZwJw7Xpt3yIeG9OP
mAhwBdw+D/KP9j4YXgNLHt19MjS6P/opPo4gEJ/GElL1fdvDFmd32Bsl9htHTcGFxjCw/6RS7bxm
RmRrUqA6o/PbiYhRuaCZRCK90SjVU2W5wbCqYsjH1CBW3i/ZBEc5fINLPZeY6zjiOFPg10hMeS/Q
MVB+P38ccXsAPtEfpnIGGZpTBhE02/or3WeiUsDAhKXzwBOpn4+wMXh4mskneQ4HNx8xVuc282Wu
U9+40bvcfQZiGdiUhSuYUPszl15YbJSuuge5hDcQY7pEddDwdcYf63stQmAfeNhfGBorALVd5+4M
cQGHCfAuLlPUsNI+3B/cVJE/RS3Nk2vSQ/HjgOSvsK2EzonFx+ipVi8rfdW3zro8NtI18aYAKON+
eWmc7qYOtqBP6kPRusN/24+3i2emLrgbW8et2Zaq7N/Ebp84arv2sm6YAvJWSew4a/jtlutAFy23
181zThJSlx1qWYFB0iU651pmXF5RRFJXTb38XspjPHB+cwS2xy37im2elBwTNH1CSE9o/MLRozD3
NPirncedmjVzpmkbosejM6ny0GKWGsmSpTcaVzaQgjCHksLej3zXgQ8hdXe08PcGADZyBbEmqB7o
zlIieiBZY+7AYmBR5uXiMlRFUAbwqTkwZtYn+lNRZLdPwIgjoNjM2YIqcNIsRP99gxc/gda5Fzh0
fN272PNYYwMdtvwDKubzfETq+pTci8yYC/vJJ7zkGFwxodIsy3eJQUdZu83LjZijrHbxrcoAj8My
UOlx+Ln6zrrIzzOj0c10i59Wk/wkAl2+UIxEwOsvWOAUGPzFy0JSlDisTIuzZrSdX2lgloyDRh1K
WPtQEzxq5L0EYexXbqsDvx2kwBd6ESEa9ZUQDWjoBLoP3QAe99l/Z7F4FrBy0sHiKpKhig2irJpW
x2p6G8eqmutQNKLJjFRFCi0A9oLiIJMk52lQP5u1NKFfgpbibk/Ap02EjLFmlR3W0gac0respfI8
NYsztgIAnNSSIOKiA7g6/csF2UW+1f/oWWBVvsgm/QMo6hxxJZN8Zddc9LxuCtGMJ7zp+EDHlHNZ
k4i83qkKESDHlkrNaVb0SC366HLDJXGMxXJF0gmbBxUyWfH30yZQvLZ0plkvJIwqS5v2dB4cxQwe
LYvUnSlYlv/gqov5r5vtTMJ5QftMweAoKc84HdVS7kSN4pBf5KgGG6evUmAv6WICYJDzpXU4nmX5
ktXVMaSd60rX1Moc81Lvw2T30WQJ5qPqb1VT8RiY/ONgNb4SQoqZHqFolFNBngr+NVwUKuBs9moy
4y9E+Pv/N43DFRB7MO5JW5LONV7MzzsTn5DAx9cwd+cPQ5OBZusrHTjQ5d0lJ5f/2b3rJOeR/V7p
rvjCB4Lnms1836BKJCU9YjGREt10Iut0eY62G5QxUlAxhyudNtZPE1JF/zTcBICQbaJew6qeIApS
HX3BmnSKgKmjVKv9XFkYvguuq8B+KiKPsdThdNRFe2U8+/yTsIxQMXi3RhaxjEKzm5ejeimKCVou
etxFfCIMyVEKm3p00B1brxKYeng8xC77HXR+Bv9U90Tt7j1IRtPn9Gz111uw9bHFSa7SJXAxmT4C
cwEYANrSCsgD5X0k4BAB3z1hYYm61lTFnuMc9uXhwNSksePi4kFpMreiY2wqI6QXtW9ivG6nOPQ+
+wYSAHEpqDA9RDi6k2GpY0srZPZjJphREaVpjf6kNGJmLn4jIwP0EVG9iRtmfLJ6Nn2lqqRYfk9s
xJa5GnVzVpqEzmgt95Z57frIJpe3nIfRnQB/xW1Md5n20wu5pNswLY1YTPFf7UT626Fm6JDGJ1yU
p54/V+Bgr9TeOSYNpKPdORVUdnLnu2OLisZwoO4i7klSkZHAiqpBUJWZqcUkOS5UckxjrwEjvYT6
FBZrzkoMwnWw8VwV0lY1vIFcZwa9IKArn8oZ7TNKxY+mHjTnLZeZtfJWWLxpJmSkrpQu04DEBjGf
p9dwOuthzo4TQV7Jy8y3fOZlWXWLfOH1Ge0XUFVKK5v1Bh1a0YKAzIJP2Qt8grGpLWd9Fapg1h8c
w8mSedyAuyuxUPetRGb+54EEE17V/XgyuigdTlZpFqAicAuqPd3peF7droNzNSUuPHeQAim+SMh3
koUblNTCLZADkGpWeX+E4Q1gqsJxmakOwWXYOSJuUMqXqegBZVRsmfbHkGFwoA+xgIHd+4ipDfgq
0Y4It0GSjMMoRr2FwrluNH+DdoHy2Z5qoCcgdUAMVpMaVourF/B04Cwm4ebEajeg1vrqx3QnVpx0
adE14wf5f5ULmFi4IOZbmeKj2qRe4YaNt8jOCEQguMx95j5XOO7dOwgkE6Qgeq4Ivfj+B06BbGJQ
6SO8u2oxEDW36q3VjaMoQTo4VcCgiOB6lHwmCqZff7OBIl6DiJ8D05x0k2n9koCfGa9io+bPFIWT
4EJEnGj8ITRRgDiCOElpBU57xS4DeGj6QBhm+Q9pvTZKf1zwg8xUIAohxsIPaWSeeGqT82OC4E/J
Fo2ElAtpSluPH03ilog7FVhL4a9u7DuwwDSizCh9yO7KqYRtz/+GFjEP/hef5f7hSAoXlxFtfGM5
vn9KN8InVyUdhqA7PoVTufKOPA6TWgNwGr2jfZh20oJ6i5RvNQF5u7PBGhd0I9mPue1GWNPaMAl9
qHa6Gj8zMDyi7OCigSj/OG7jpOIt1c0cPf1kH6cEZa+4uFOvb4mHPyCkFEykrBYJHnkJj4G8D8/p
jWso9Ep2kdCP55dzlPZV4HIg1AIjMGwZ+1JjtNt8ccb1Sdmy0SuIsj2tqsmfD2kT/2y43rrzqkMN
jrL+UYE0RthA8v3Ivmjmqw2tXYsW/cT/Q88jXjxeb5Azd/uSKbyMqgJo97FFh6lb3oNVLDKv1sxD
iczCrLAo9VtZ09B1yZOhKQ2Y/bzz3YBoVTJhb5vueK/MbOzpriC023HXQ3jdgdSr8fHoilWpw+ow
P5K/1jAyA+2eALi7j/EZqYLeN7qWco7U5ChNsEVl4AVM/inRwpGmbCRvukqFTtLYnAyuQHQPyceZ
b4PMaXQHzeEKymx0J5zBWeJ4m1fMDAhM4ae/55rPDr4qjz1Y97AYOWsHdR2VBYpkhk7W/M+q030K
r3SHKeq/xCLNZddKdLZecW9Zrt6p7uhJVi/aEstPGsNeLbNndhp0Q/nYfRrzDH/oz9oc+Q/SwxeB
ooee7Evz4bOHgiDQfA8xDTefhLKRY8E3PvHj5k2mGMg8hhV/QyKYaYIbtF/QzL41i6MsQNAsvE/Y
TrzqxMNV4+dPYLqhOJICEtHc0maQbmmNtBoTg/NeCLur3mdFbGf5RZo9Ne35wf+P0p/yBFSmC+FB
3poXFebNXudOK7w9n8mm/6KmvhifLA1+EsSffLY0m1jc8dNxM1eWjnhIpG9I21FMmdnr2Cxavu3x
HUfvGKJ4jxl4FmNEyqr/QTS44/KHaAx2YjlrdKN8j+PJRPWuB3x0quaChdDtfM+LZhsSK/JxehbD
WqDY7FbusKlTmWimtQrQVAfKHQUx3bK/qz0+/MpfFNY75NMwNasJ4rL3Cjvzd/+XsBUaxao0hCZ0
CX9hcPtEWV4SqtTm+uIzrUc/es+tbdjqJcYfGHcv8uY5SzB+MZJDVMWaDUAoZdXbj3+1iFniezt0
p/Q+09txRh5lVxwEkaxf9xmGYC9w1VA7maj7T5aU8/q4euh3Z2iJoV2XqAA3Co0s0n0kC2KAwACJ
VOVKen1yfOhrkZeMOpsWv7QNgVN7OdQOYawT+Y7tYvukth03S/zG9/nnTg4MXYGu87ZqojU5TfOL
6YgP1dyT59EIvqNtGtMTJkQiBwx9AEnW2EKhe6ZoVQwzDs2SI7zSwRKxOqjn+A7QGI8rHa94iJ6B
2MpMyf58Qcd1EMd1Em0V6vTZnXNsQyUQagMZZELE26ili2jcGp7PKBEKBtm/iKH8tzOVlZBfC7I+
gk6rci6qoB/1fJUc6ORmZFFaBfz2rXkCQI0GiY8M9ctwqPolP5921QxsQtTH19PZtxcSa7fL6e/M
0UtVIw7jZg9VWP73YZdXqRdbMzfW+CsB/RMp3VXEm2DRfpBi/xdD4KvttVHHcGzRIOwxxBlx9Zm0
19KDOZLpLlsoFpr30b5DJyHZ0VQS8NQwbikCKA21YP3RNqljRlaCemkpFWU+d1pu3KCoGPdqoSLD
G3oFDxdorooiVXKHQIT5nKPn21yhN1Bh4ri/8xE94PwpQiLucz9zub/Y0wAu8y6rLY2OtS76rQ7o
6nWOjlKfqB5NxM1eQgyiSaMFELNMg1KnqZvw1gxAMXlNmoLVjOtK86JjQWesha77ilNMcDSOcMn+
S9rBDwCvEWQYWIfAeWTX5RVuned2jhHng/3C3ZuMkcKpIP0XayNMrwD09fk8KeLUcuCpiSt1lv9j
xjajC84XTpPMCv1wSKtkPl+p7plAqpqWiRpZ4OQ+GuwRADpULXW5ujjlnjBHmmdbfodIbSPYUeFs
X2h9/EwXsJNf0cLcDOCGocdJk6DqpjJNqDWoZTPBG87nhKP0bilU61WjaIDM9F+FefY1hmxyCWnZ
D08hSq5SAbx/HqCrxw+3E+uN+1agw0A9O6aCs7sF5XRHebMbB1Vu5EUUAocNLU1FPIP/ZJa5w/Rp
6VSiM/QWNK63DkWzfLB8cj3J3xNeQsViAdjGHCaVLl9fAp5I7KWLVVdAkYZZ8sIp69YZNo+rSRj5
oh8aQPlyQK/qpv4bUGFGzZbZG2yGb7NbhVH5sW06AnePFsoQw8HuiXhblFoI6tIgOeAiFaYmNDJX
8m0pPMtQfc4rGsTgbLhLksj/xleLdJlprnzyyWsNCYfXp/qQZkU/z5sKXi2L7YCzb/Ryi/sa5j/b
5nHm0L0USJUv644Kf1znZvpwdOpHUi785JbQL4vv8ORJw7kJ5D0Sv75c/8CIQt620+4IrZ+KqKKo
nW+cwYLvBKLvIAP0iLdqzFp+axM0vHoIuP+vQwogHFTpg9l77Dcu2ri6k87FpwFIgeu1FzsYkS/K
pdoxgGOoJRM9d/ms/c77FJj3ogq3CL7AY+WVI5tQMOGJQI8nex8idS9tsP04NCpbdBM9NO1ybFPr
GCU98DLz32qBvIAW3nfJs/onDLZneLC8XIqDZYUs9uo60LoeVOah51JfmUzvS1DC7o2TBpGnhGmG
jFNC+IteLvMVgbFL9YUmtvMyuLzsdPLVKkA2Zo5wD/U1Pkpm15c8E6b/BhUMGezffI5whOU4sCZu
jU82bH76auNregVsBJmWeGUH8hfwbMMoebLZ4dGzWxNj50LPMpwPQYEeYY23D8FY35AFmAAqAkpc
haIQBIChkLGO1rzaUsqgfsSmzpH47jzVACyN+Gbnq4CULzZUO9VnuQJaOvBxBmsOGzhVTg/76yA7
tyVrW5QpYezDY8ZgVyqjalAytHGUnMJTplpgzUQu42raIMb5D+HIov6RhgJiclTquztCjuwQJqsC
p9C53MjtMXiGGkSnjBWhSvDM+NmXoApih7yTXUx+J20v6fyS97rEQKInr6AKO31E+nE+vEgC+Cvg
bCYO1R01urzukEzmYKzR1rQQco72lhTQPn3IHH744/JbS+zMFG3YQ1iYYnnnhZtaqzBs7K5kHdfC
c5a9e55rvLv04dg3fcDi+INKFnhqREph1LQTM1IJgwiJ6K8GleVrckSdJoxdKhK99i9Ek0sSZblR
DI9l8er78QvnWKnn3HhyBQuaobR8vOjd289VUzBCBgCbmndeznJ21fJ696pHwFA8mczTCPB5it+h
zd+e/WiuoBfO738qvia3fDxT+bP2h9/P1cORMMUXHOVU5eDQQaYbVB44rQZ+jT7Gqgg4UKLQIWUn
g/OJkcqT73o6y45pVi5krC5wQMXp1E2yvVOyvwdW5R0Jkev8gQxBotJLSjtMO0FBQdNEJ31gZP3K
B5NdnEDM8HcRDrTuy2W25k+9wpIzOGbjWNjyFsrjgKaSSFN61uoiuiTX/7WGxgAEm/4g5H+Vo1W6
VtxKZObnsVWmmgYJDz03jzzpmnILXIu/XmnAcPaHWx4TbgrjCC5edacSH2B4Yj9DjGLT7AOe33yJ
0RQv739323YUtJ96h7z4YAGryKycUV0+uRPH0gWl8vlPoWxwJG7zDNHfb9sOd7r96zjf85OS/BxA
/BXjDClpOKCiWqN+RuTAr/GbXagUDUxZ04qXhrDhq7PYa+L3Of3ehLDLS8Lj8pPmjF7L/ria9bMV
U5BjHxDdsTVRGrYJ6riL5avxYyAmGMkmg6/rGbHhgn2sMwLve/OzKNsft8huGbY/US6sH3xRNbVv
7IkCAVeXflajgaZLWpsInQdW8gkqPtIA8SpPgoAhKsUlppBy0im7PI0/7zwNSJvkfdOqnxjCCYEh
A/B2xMTKRl7swRXWf361Ucu2yYi9u8LJI+ZpsXql7Jarrds/vsGAL/YF2bs0TDszeTOTcDLUDA+o
XkM0lNJL8ZtsqQpNkqYB6N7sM+wG/F0OQSbR+bf34HmjK+MM1RxtCsV/K1ubOmT9NC/cGAlAoanR
a8rtNWT8DWxQpujP5dHAV0jxxk0ocPegBbLTk1UsLBFytYIJ7U1SwcBAo34KaUfa8dTMdifPinBV
Tu+tI3JT1xgqi4dbH4xreV90oR2kX86XCqq+iutTj2p4vv1DblvFOdyuP8UpLOPMMv/zKNuUvNVU
7+NuuEt7VGU+hLs86eXAXo1K/4DjeuAPIZHOlIGLQ0rJOnmFoyVZX2b6QyMPyP3oH1JyNJgF1son
ZLHR52bkriXGFBFhnZ73iPSfB0wH/JaifRA//CvSxNK6JlKPnEZzrt/ee7ha8ZH9+K/BS7VJOilS
v9bgYE8g+1rUnask1WxK3Vgrc1iaU3L4mcnF2+Pz+LWLkFMwZhDZYMEkuP/7sTy/SCvafr5oepNj
UXguVSenqJBTKMmO38l5dhXjhUdiZ45kB+JpOjUztPzj0RsHsDcGSf/fNhhR5NY80YnFQlodaxfG
w1RA2QQURDKKxQSipxeI+OI+X+PhF+narkYVhnuVHA3sj2X9ixWcyBinZzjPjk3HwF4xHsvPuJmk
7BlCeHC+mjzolKsyBq10eejDdTbBPLmAb2/kQxapq7JzM4906+E0Q/znIG8d0NCPYjt/41FkylxJ
yXRHJP3s4mVUC3pUNwO57LLPZodRbDCkIbY8qzaGwqowXX1mycCriHOTpkSdjzik6QtMVTAolSaT
vQqVlv9kg+ddev5i59fPpBgO955HGMZP1FW8v+26Zx9i0kZTAoztTKMkvvGrkw2I/CGtpnwgd8mi
PQXRp52/S7DPqBBDwkMMKeUOVC6WexGKHExH7a7a+l6dGfpimu2rrSuAgxnWlrpKO5mkEb/7ZLGw
8IhWo34AWjQrYaR6eR2Xc10NqD5UGJU+f7NT7OXJ+TxSHmnJSm1BLGDX+BLjcpkrmqjybDNOz8Qe
gPFnNEm3+8EuOu5+E+X7AV5cb4cnD1fmCYfvfsjOLfTlsGu+CM4m8PsaBavWVSIEmi9ctrOokL2h
JfjQ+xC45hUPoHLfO7F4DDkgMuDatljTlTGA0Zp8fbyh797uR8oktxvRspHnJiBWq9h0UgGntYTw
F+1k7C08z2DzhHbp0BOCvmLd8au7PfKjXz7GXIg3su/EE4le0MWDbSdCesA8O2TCEybTWHxmuAHN
wD0cSq+kr60D7xAkcxhx0NbYkGB8aAcvE1DZ6aptNhXOY390/prkHDVnNAK9iI0VZgD4zkoHwpxS
d1RuCT1HPiBC4lN1dWwlo7sIrDAwlDLkJ0nBGyInbrI3doVNw7cTbWu7nX8VUn7lA77BTLAUCTk4
kfZf+ITAlDwzc4nBMS7XfbOWHmhuyPXkyAjenInSDnLwEKMYjNoQ+263uGozIknpC6NT7sMb/EPx
3d1161PeLtT/0CvOhBr6uM2tfyGLcpfpEF7IpR1GY3BYIr7i5tvVFdx+dXB/tnQi6WGToPF70iRJ
pv7FLrEKDD5YPAforrF6e+zs2VJSOUa20KlXQXwgueTZx+pu/gJdMW+3p0UCyavoplRBNKjgQJh3
Qmsq0r2tI5AMSgBnwluYtq4yFvWNIykAXJUFp491fXPbZ4vrGflGlLY75Zmgig3dwIuUvqeMvD1R
kap4zMYkiwmsFkctZOISI+ELsLN9rDvyWAhkHkdmDyV5QpOa6WH6Zfgzm2Xu8i637TT1ewO2lv6s
smbfhny5K6SoIOfoYIwVunmT5LPsO9m8N2YSRlTx9e40DWWfRoJhqR7pFvTS9tGVPNezqs/TktLA
RkLCFRsHKaQ8Xkh1KVgjzOCfe1CANUSZpA4ycDQBHM+Z2bg8O4vHmen+Ryq0EP0smH59gu6hSRc4
A7fRqRrnqIwERB0vUbdj2u2hHRnoUgOTszJwP+er+2UK//lTA3Ol57I37GIKZQZBfWWsBk3y8Wik
SinxnNpuB3AxNyAaBe4G32mY+JpqsxgZaoJV1mYtzGFAEmZAg1wgi5gFgSUDVAKtwKdizb1mZA+e
cjZSk0A6kz9Kol621eUtCeImq9GToTHdp3X4YHpjrz5pv5iWE9WSsoqEVYoHiyihyUjjP+SNh2S+
brhZ4Aic7tCiKj6nWX1rmQdHpfSM/Rnkg42uANJaCFAUHXjrkI3kIhds1o/JdoI1fYlM59UK4iBH
VFWgONhjGKGvrCQhz+QzfyCNKt96qs8D4sAo6YoqJLuXATju/33Ca7go12hd6NJYV+AwsNMjmTg8
9B3/lkOucskqqcK798tYhahQigwWblFFquD9R6oFTgOoDWekfsCn0Skc6+39KnD3vyScowanvVkU
Ux6XqVjlgcBBkPEjCKcotyrrEY+mL3FpzwjnCnMPQTQRaZfVQnpHi8xy/zoaZdsHh5xrpR5g/FdJ
ZWNGlaW/pccNxYjuz5Dz5wWKIO0e5JxcYX5usmArNOHYZY07gCFgKe0oGZlB7NprgfpQwAZTWeO2
RsFBn+l1n1WWAYqpoQWxs/7hddSCT11b94ib/LeXV/84wqZP2fJdFNFE3DKHA/75q+eQlS+AyZqW
R5dw6XqzHb7CKWdBTCe5XrdnbfipTPMYhE9+GfTFlA/hwclcYOGguUJaiCvWkUECsVTkwubG+jtO
ihIMM6GjxwgEOOyqhb5EaiTa6SjAyn7hXuQjnVKGBiyvOxcQMrlcWeTfELRhgpHBm4b8nCfYSR4M
HRQB74SiwKsSPqrkWcykmlt7LC7ZB14Xisyi9IgtsxkVlpYU9+ucQkBn6YNbgWDNzOTb5yDuERVq
XRbfcgLdE+Ne5ZE37wSkAo4PtOAnu9lc5f1/vn9e5dTXe45OQu7vGGMC19Kz4LZV8ktdnbrSVl18
GwYf5UUO57zKeJxOG1lT6yq43PIdwztv3wjLyc3lILtV48CjnYSnSLqY4wUFl/ndjCSS5A7Hu8No
XBylwTonSTVSwL+F5aRoVAMQLFRZWmWTmwGkiRKqYyE0UXJtLvacEiOLJbjkjfwiJBMMeEPvaeCS
8gNuWji4dIJNZOfTtuMu74XdP0isICWGVrUVWdmMgOBtoWYI7/mo9HzfNYSyH2+OxydGcvEI1J/U
3uC1rYAHjYvQeLDqT8XZvtHS6GyEqt1y3C/pp+WpNtidupLwL9HeF78mrKps5JevTWucS5K4AqNF
B7M5znSDy7DSju5fXPCdeIQASH6qUuwEyfU95VR/tPmMA9Y7UUWFOArSsgxMHs8ZX8b3drS57C2u
cE0R5DDDyiutV+Txgp6iSo2xfKPyR91CJgMbica1riGQE+SU2pjsJl3USovZ8z1VZdR/FBEDng8/
LFNb9LxxIfCqt4ELsgSZqxaeaFNCt0ZNyhd49TL+9xqUMLhiEbDlg5o/SejLgKWkTQeF/Pzqc5Zo
bbnHVz2Z2bsjZITp5Ke053OYX6ZIs3wf0R8IjHbf+iCseeZuJ6yqC2r1Vnm7sWzjzOei7htWh3i2
93mAmJHwLJOz851a5xTNB71j5l9hQ48jdXtXhJ/Hd/ubomDSfXmhNrobqfeLBuurl2Vn/jtvJ1HD
X8NRQlZ6GDfsg1CaAwi/0Dqcseshrqpt9EckHQyfXehco5Q/h8lQZrVDdOyHoepREl1sZceUw1ST
aCvUIHNUzgXKWre8nXL1cNXTeFhACNwodt+Waim3nIuRpa0Cbvg2L0vCNza22pVTrmarht50+oMs
NNC3EFNbguuZeOnRSLjD6jUlTHx63K1NEitI7wSBmsYr+/bSsdo2bmKv9v32SYZc3/Ijth9YROav
CcHI4OZDwSKl3+rKUCp3Puu8u+JuMv/uyX+OU5pyurpNFQJkOGYpxR5Ny1fXfgqNkuqeTjTHNoEO
U2K4OnC1qHl/g3VAOMioljYPSa+pRrSecyFOL+vnAluQjuWDPjNY+mGqkbk5CkVGCWUbd74/R6rV
5SPKW+4Bo/EbbI01VRX6b3zgHR5VZr+XDiJwaQctnp6EP9l3J7oLJRo7ts6nFGqY+6vI7I15wslI
96/2Dbf6du4m2A6RiaP+WQmD/C50pPU4AWZl0XdfEDCYpwgjWufdsKuD+y/6zacAyTUEFvTJ6zFK
M30aWrBEgoiDtkguewyqU5dQZ2Tz3Kh7NLGmL12T6XQIFGWt7kl2Q7ldBFLDQKkqZSIwi3ZYe4de
pklXQd7LRPxdGDoOqw2J3MqrvE/CQbh0Ec8VXLjUpPFve9T6eir9vMEvk0VgATiifnCp9ke08dJo
KCzD1Zz/fTKt92AVI+4+hVePDaqgzaX0Kz76OLZsC8mU7xHH9MPc+iojtY9Z9ggroExujLEdE077
sPdv4Pj/ntEALOVAfvKT3UsZtAG4aWIS3+FC3RTW0fRLmFn0HjuKQP38IVQFk8iKQEF78QPiEalI
rDKTHdabwa9QAoD0rvMLZvJWG50mXETeRQCoUvQH5gjDnlNyNyYDxZ9TEcTE90SHurYzAQqPRG4z
6/0AYs0HYjG6PJfQEsZbT+7Hpjv40JQDk1LUxHiRfRMUoKsaZn0iX6Dhd1cLbrloG/CX8cT1ijye
nS/jMBeeKKTM7nMiZox+sWZ5zqGmTthuh5HHIl1Do7XDg5MxYtzoGTw5soGC6Joho9dB2jsdcyyZ
SqxAu9tKIHe1vXvqipGzA7yBhOmm9HyjCe937Bf1VC3y44We6LsFi0SxFSi9HFOD1rlQWMyi8r/s
n9JUDdPsDzPLW75UHeQY0QVmWu8uZwsepS4j0u8AwPfyYiFP7nGOycIOm3M7nJjDTXWytJgB7P6d
vQXOn3EmqFuz5VWQPU9P6S13yZ9LeTPGrmpFuuQSnt3hY4v+ilTkVdRDBigmHVwRQC07Htrg5kNC
JXxHtQd/LpSbUaFFaZW5MRDlpMlBPknbzBEvu9ZVjHPNpJYcpLENdRaP6Xj2sCRe7c4HJkSgAecG
0F1jXAXDvN7n9khwBukxRUHVdoos5kI2o1rMOivBKdrR5hx2+O5kdh7Q9sHUIO4MAhUQsSH9RPKX
kcAu/T+pYFYzkxhqZDg/vqby4zb5Sll//PZhcCEWDehBH2OGQ2tjabYE/wtdT4qzrxBloGXgeFTZ
od8fsJht09s1RKOOoLE4O1Xe4b8aC0O+WVZXhisaHyuwvh2aq7sZcp3AEd9dwGWbCKVFg0pLj5Q+
lV7VfrI+lh5TM9Lo4cvuL6RDjGFUxqTomf5FuiVV+A/aS+nOIZHFP+YN+sOuQxcJGQn48P6nV/ev
2Ut8Md8v7QspC2hAQoexTHV7ZkJz8D0V7VNNrFklLY65OjgR9HT7KtJ5/YIALnpwkL0ubD+MJTAe
TL4hoeaqrZ09sc1Rie9Uq8VM4QPa3wUpibJw9cZ2hXp3bJegnXsPY80ONOfUjTj2NjHnprkunQO9
Dpss0AV8Ua9RnEnZafOtUK3Ix53DrTMuQxwGC1HTEIJZOMgnYg8dmSTg8uAVD+6hxnPkc4KtS4IB
ZwRWrbkqhAPl1SDUtV443E2/ocQjQ9ykIDl2t0RTQ785YAQStbGecUkSLS3yO3CH+DybK6hjFZKB
bVixe8HQ+GpOQ25wtL0aNSksfpB8xXzSEdG00glZWtNPPexgNGlIizqjdJfiNNTiHb7iMQEbzYz5
FFmGTcQZ1BAUNQoq7rVw5eMdAwU338x/9y3ceqkP1fr4qKJ9DZIwFBD6hfstgHaMr4RgiWAxfa8M
A+WuQgvbon4LNARvk9zsiUNcfAsbTvp6ZfzxMKWT+K+lXK9wkRk8CoSUf6Yi4ZAedxlp/4RCGtCk
exDwmhyWWilp2AIhnf8tuD1GGSwj9Uuec8hDX6Oy2mOEMdD9lrP8E4TzuSGDUCTJGPxxRR2OJ9Js
cAxsofoHDN0I+oqyn30xZj+nnLVXFQ8c2fBLy4/YrUrUznarTMm/hEDgy6l4d8CBfozTrqW7Kwqt
qEnHhMH6jcWENUWZK23WQd++cRERuDQAeev7zMm0w0E32Xzaje/QXHrXDC3CmXAr62Rp+p5Y/prs
rDYf19KtdDrhtpvn/wboX194kKXjE5nkbY6kCY9IWGrZysjhZ1rR9YDUYL7mJVFdJJtVXjjDvU9l
nyWwLtc3sjUFowQ3AP34m563uzsj2k4mrJGUu16H0tjmODHPlo8xssSwX2O0Dl86oDI4Jp62ko7U
8ty1kyP/QQDfZ6/SFSDqEx1hqaxAy8JWWyWw93bKjtzPBQQNUYHyhSmcgmEIOKl8akXxCraxXwTs
+ca+S+zcNMypZQEsBhQmRDS/ceyVwQarx2Jslit6/T6OY2Y1cA6jCrow+YoysQtJvy3iRUDnqG9d
8Z8tiQenIJo1uniVl2VPxCmS7KR0SWUa3r7w++YNBYOzDmuHP9B03rt8FpTxUymJ9BwQbfu6oDDK
3bKDo5vVCgUBs9eK5WpGJ2NO0AVwXG+SHISsWgOYdiOBADaPk4yOo+XT/Cb8/LK+cWGTJ8L7m2Tt
kIuZJpY8l8fEUjuW2tYLaLX9cxFgq0KP3IONO5X4Y0wb0Ip5/VwHwRXcr33N1b+s09GUf7G29LvO
d+OiUdt3t2t4Nzp1aPHcj+byuqsimLkI0OM8C6HNeH6mMr5h4WdBorOpVKwZAggJXLURIybTrb+p
arRHbGJIYWoOhPlH/9462YNt/vUGu7d9eo9q0d1zUKvxwlLHu1kVfZF6yJK3unoFCfektngl2+Bk
Z3AIk2rBz9ADazUWM6dSLekenhzfDvSVE6yvVPQIrrzyqxdjGujQgrTdEFVQR4AU6Ys69HX7qHCx
yWKa7Llf4Wq/C0JfumiMwem/nlmwIrHNcndyKAcU+eq03g4YZnXCgJexbmWjvyhObyQ9v72xrEdK
Et2yqPK7JTar03QFMP4w2ZnKFROwDzFiPKkOSPn49/3MBJ1PaZkYwODCoslIeAnVsg1RVUbPKiep
00+Wh/uRxRUSZ1lKwa5mSlf1PsojV4m3218swbVudk9ku19tbNx5D4fcj2GTU9d4WkPJcgoZw31o
RVFneHOzEfX1El7HLxlNAZNsPyh/kWoWbLIck9LhTdC1tVX24cAjUkE6QAoHtRlmbsEZm6wO5c7n
QfE7k5JvRnisreWwVh9Ya01UwauBXYIHnFBrGkIW0FVC6WZqQDJRJWYEn08RA5I7g7cgjCzb2Umc
Ycu04WNUWfNfNxjFip59uufODwPW/182ATvS40Wta6nd9w3RHHoOmWjbEHgOT/vLBvfdKrNnZFiZ
KTACPKa/a6rbyG0v0Ofyz9vovHjmOv3jRpz2uJqcteTSaM3zalt/CS4Z92EaPMezV68wCjHa7a86
gQdZt7XerRZpibJOBRKWwmshA1sG24F8PwNdPLKwGZGlck+/ZiOZEJPVd9XLjRXA4DqxWUpUDlyx
Gg/qd/Pu8joNWY64r1ZmC8ZnIggWbu2riBnRIQ5JXHLJg/cAycRU2aPLCG+prn82mpD/5DG6wWHe
a8aUCgBCLf2wKQeIzDgb9E0TVj8ANKM7wkbqmepLOxjPuxCzYAhuhjBXdFNgbVYzfK6Ea9znMvZH
I6xzPn7REcC3KmuzxfhJM3SZ85AS67MogKU0G0SMih9SOILAQxycjBm1m8YCOessEcfo6nhmTxZ4
gfP+kU4ryzE1Bu2Kb6pkaL01WKTcLxoKhj0yDHgyRNSm+kbpr1mT2Nqbbz2GyFpqx3nbWPEjrxn2
ezNRxDg4F+mGo1hgsWPhclTQi0gxRTOj+mCx2UB5NSZgys1rzK7R889bqPyutPvMQJiP0clsWQ4j
oJchsoJE6LQD4bN0wPhQya92epBg9ZAyot4RqCUGA995oJVAFjf9vFHqojtLAzo/u2WfGhrM8ybC
ztypgwKXa4eDhfhyHWV3Sa0kwNBxaoEfN4jQ0LnLPBrLMsFzzbZmI061T4FB7xZjTIqTA4Okdiqc
NC4ZfuWrIISHG2DEcvNxU2ijGvZqMZVtK/eMdphaHZ21OM7i6CMWZSX7xgql1X5uHbgsN8A07uxP
ebh6iRsr32bBH5wWf/AnlssxRNipoGePRHUNQnfTQE/lwVWZBXiBCre83ehP+JmmrmVW6RvhgTgr
OmWR0tY+t8tLgDN8CH6dK3fqM1VxKTwNZny8mZW2iN0N9LgE5JifilKpfaH6FeuCfQefB169pSEP
p45ULIyv6n0nHKx+i1ryyIAwqEdQ62LrbB3HfVkkRbFRC/G8QzroO2ZGNWOeczf1P9IOTG3OCv5p
VCTGiplEMLClmDg0i75fehZbnHgMNC5sI9hjLfvRw3WY+Kp01EfWd2iatfJKtac3A5PWR+/Pfybn
QCcnT3JIM27pjW/Nqqj0YvagCaS63k57JgHyBGyk5awUigbE3shNkZfXi+cVGMLShIdaulBFkTBZ
c06RCRBPq4+qUgw9YZHtha0IGKUlm2sNPcJuebpGjNqncQzMY5DJuQzHMn6ByLJJYKStOLMnUkL6
HiOAszv/3WCn6grFgCp4AqIEQfMpjP+wHUT/Nnionfv9GbXAiq5t6jZ+Vp3ekKHYe/nVdtZSX5zY
dJXrs14UEXiAGPlkcnJ614Jx+GaOiA1tjiLIOWWTG2pqTZjlq+Q/x+TEm9GQbfYjMBVftEzr5JBP
d0b5TJqagBKmqvqFFdaMlRZGVRAse90W6LqlHVO+eatZ5Pqrg70jJ22mPnlKdP5ROuLvZniRONmX
phOO7t/GJn2ICcIhhXNOOASiPHrSCO6iPwQbg/7yQPxcC8nmfauWSK7WgdsG80/vKhcRGI8qyQF4
rhN7LiPNG+nJfhBFIbGAxnDN8van/rm5bb/Mejpp/DgZ4K2xzx3yPD5Ep/c8F9qQCvja2q94B2jj
hmkD27ZPOcan/Hfqzx0/L3oIkOjZrzk8PnG8YTTH/es23CXI1VDxUIuMTjF1BBcGvhPIoBHE8jTR
2lNaEfMPkndVHJZdtnyulAGaXtM9cdCrAYUFDani/BBYUJqQHLILlq6EQEbU9f32rkmHpbccKHSF
w4QtqlqZazamywnxbuqbK/q3zdrDq74ikVHKGx3ub/DIE8NABytCdMF0aozYhgsXJryfZwa7ibDm
eYOyFcT/WK7aWo9sJx6ECLWqLmLu/zGkf5I0vwb5lf+zUjAs96eNsI3er4a2OyDUpxIFv9pEMdGN
PvoljnnuRurhawXBenZWm8G6aHdYcHndT+rmQ6Yipax2Ea1YZGUQByWTsN/iPyxA+EJQzhUFM3A6
4H8sIUQkQFYelN3Z5GqNMvKzUB8iNK6KYI1bLRDF3EJcZi1DQ9qEpLJW5sXpyZAs8dgMdzLLKm+k
Y10L+zgOT8pmEUSY5MBg/Ous/q7q/B3pPutPqdm2jIollHbRfYoUBHsezXzGm9ULAac3rAEyiDP7
pqZDtbEoumvGcsZyCB7y3fy2DN8JS0boyQaU6JV7dPNPimtoS0YbDFSpanM05rw8EPHnkZ9tKHL7
Kllb7w6TgMNDzbVQASbbYv9u/YokBgmbUglRFaT2on6mX/4PnoORSoglqsTgw/Pb34DKidXgu27l
zvzDiwdcHGhLuzw4MnJXOu8KaDViWpiEGwKYR+PcTyhB2A/znskzX5xDw4M9VbUW4l4ydce+p5yT
qXhSILkQuEs7zp8hsqDw1YVbjuEslER4bQryUkqZvOovga2qX1JC42L0Vh8B+rLmJZ4PfDDB2sxO
w13rEzJ0OLY6/rskDQvxY3RpjZdQ5/DFqA3fBc0ZWH0aHOghPHRMXUSq1LnI2ituoQA2kjFzmz/r
e1a5/1Egs8triIAIcGL5E52K5Ak1U0FJrFCS9OSGez+LS1iTbfLEmqYhiGgYLUV7YXyZgWQZzcOc
4Il5ClbtgO/88lrECCU33b47DqDG1x9LvIgNCWjdLOioKP6lRmfSnHrpbGMrSDIxTfTwjg9kFDgt
PAE0pODEndMev/qxPGwFEshTjuppAXJ8vCCD28SP8NN/p7QuC+z9YvfS+l46C9CJsYDd4f1xTteH
XQkha6drZNby5k9/TE/2nwdoX++g4Gulr6T3YTQ9ksB4lQhMgo1DSIPH6VAoho6bSikJUMDOah/1
qJjkGPUIj51DzA/YvQnwrD8p/FblGTYfRVh2HTEFrMy+kNX955KjnogV/Uby1An/SQtxDklnuDw8
oQLQHXFR7eu+WKlzWgJhoJ2ptKRYHkKviNO1BqX+Tv8gvwPvdBB5t9ALqO74oobdy2/aLowOQ+vr
m5m/7PfO48X5vLzd7YbKYnJAdRiwg57/HMIBDmj3pm8lcG4z01K329JX2F4S3O/AjVkr2HZAgly1
KsWq65c7sPi75qK7a7hgDqgBT/qZUYB7/SEab6nVUmtns5z/h/pVp11m/jkOVlr8lNVWF21WhY5Z
AEHFLoJHk68yed4OPm3/Lk2qpJNnzloRgQPkKU2PdXOGlJKiB3lO9n3jz5jvfFVpRaiUQNCRM8IT
PO7aU8vtWBfEeePkAMKWS43KTorgPer25QSEzoveuKeWx7SM7oluvDZ87kqU6kldf317GzijO6Vh
Z6nbJGJ5lUTZ0VRHqIKLgHJ3oDxFg8vr8WXtiiNpQOytXsn+r1S+4SdxRADU+XVqPSjurXTF9ZBq
RplYSTzGZ+RpX9elu1XSL/vQxrgpLPIbNSVgSDoSdWA9rssLq+xLOpLQw3p4OgqqP1uoPBMBHbDr
30y34aOeuazg/TZKplSjkpH2tb2CzoJbDhaiy4/utCvWwUSm3riUCnLKBu59SuKJzlmyzZP9KDY9
o9VsOlPLWcpzhEnLfjBeXIA2B2pSPNVPlhorhFTSlpqeyv2j+L8vlXu97DtcCg0gkVOIbAEyy1vq
7M4axBfDP9Iw4pEnn1QI6mHzNvxA6Ib5fihrpi82jCwoliQ1tvcJeMlp0rDb18NUQ032EN5I9nXh
H2ruLtr8fuLNgjN36NigI9AItpyG21ynn0Hv8wzAyqUJFBrS3tl4IKwJCeuaMFv7SgfiN+xBICo/
cbXuHIq+nhj/arrHUkmMNN1Mxlymp2kNmLIuot0MXqWMdxDPYhyS+U97IBRYe8HEmiJEP/Ij1fjs
K0Z0UE+C7uivDRILwZNwgWwR0TiWt4mSjsUi5G2zzRBsKVFCsovIYoM1F3Y9F2FMcHlc3PWu7Glo
IuZF5Vern8qBk8qWqsrSUezS0LpUx0Am9+MWd0I7aRzrcs0G8Vgj4KxcdGT6xdE4Fh1qZs5ABT1F
7edzY0JcyvNCkJOCaJtjqKNfWdJ8LcoZTIiIrCbUsWy8PwInanVc9Y7XL5/oRWJ3ENlmKsBa/Pnq
13tUTB3fo6srDlrzpIItjqQSXIZnK46JFk19oWUd36tYOpnCNs+Jm31txAO+g6S8tWbwydA61zNA
GRskaAqfE8RRlODUY8w63DecXModXEb+ikzCBGJhc2o0B/xvD9Pc0IczUyI6JT7K1trCtzdPuo9Q
pG7xN9q2/okfY/lVA7DCeeNnNjiezn6OdNtO3m7Zgbb0jGOYY3+h4lp7WohY/pWbSgTEUU88pOEW
ImASH3fXPpssevcWeTrIs/iILj80kH4o5i9cDF/LRwJrG3zXG80ZJIV6c3gikXg55/49E6QXNWp4
XDdGQneHl4LSH1EyRAWBb6MVorUb8LjTwdhJLThVkdlDHC4+uS3l7urlUfqXiMKqYfXG9n/8QbtZ
mX4d/N1IQqZMFjImbpoeelsHnf8PJ7G1HnitWQ53O6AUQxzpjDLIUXqrUoCX8gPL4zeohNRtKqZw
jvX+boWqiIF3XjiNOxQzmZ5QB6p4XKLeCijFSKBSWx5cotiGzSB/IYlNWiN9YNmcnpDZmKd7w1W1
JryiIXZXZsht0s3JADXK6UqnRgp0BrXTnoUpcJgYM1usU9xfV9KeLQLY0XCLblWp37v4lDVnwlCd
RiIXD7UJGYQoSOFzP8MJZetjKFCZ2JH1+8kmO0C9QvqfdoDdcI1I3PELB+5yWQ7hPrjjbd3kFEm2
/o8/D0XWvo+JbzSX/C0CbY2+GaIvf9/EV8fiyUItSzD03F5K9eA/+eJyKvcqo8/ufMaaG9lGx33l
1qJe1NeptzXm+yk077R99f2foGg5qwOSedJKzPZtJeLFnVgZelfLjQr58UeJrEcdXlh+opUj0dKw
QH7ozycsdIsQv1yd/rhKJTyE/8c8SgAvCySTt943ZMqWNLz1A4jNyHAWrzt1vpYnTY+Bhq9Ym/Ow
hT6+byfijsx4IYdVu5b1V5pgxwihDTVz7UA6ZYxT6CJ33H97vbO8xXcbK/kK6YCA88BgLxYhiQYJ
f3SoRU5Kfp+wns58ANxUYoQILORESBP4ym3aZezu4AK+ngJOw2bt8TQfUzH0DC/5f4xoZYVBguXz
P6m0O3i6aJmcIDsooPJCW1TOAtYKiNJZBJrat0H0yUcYNNN1mTQFjiGCfGURB3mzZuu2fxwDk/49
8QIz35YhXMPEB+1ioEVJNUu8n9Nw2MlCoUl2fiR1Tp+2RU32wKUcf4u8JOqb465A8Oa4PdFTW72t
2+F0/wtkZcSjSGHStXNm/ImKFMMi2Tnsor5AbpNr0oinB/PnwSMyqwx2fb3dNtezKGjguTyEUeP2
9JFttxVBoyxWcp+ETzmYO+FggASL6m0ckApyX4fen7DjOHrCT3bm0XL9oZ1BRShNxY6UMbISwn+w
msDXVYtlexGVQ2fPVKgUJ4yJDyz63EFt9ek4uKzNkZsgaEs/hQmAVEOq13q4xcgmG6qB3Qus6ZQ6
3lh0CJu7Y7bpFwmEgL40Huvlh5iqcaKqBofH4XQS3HvTx58/twJ5gcupx9LOFcWf8INobGHfQ3sD
cZHKcQblkqzWz4pCgTR5GuFiHxcN3DwLBeT4keRD6S4tm2CvalXogfqivCczEQuKBqPWOjrL1KD4
nJPup0/14xUcowXOp6Y5qtfFCu5rLcaTDa0K2GM8199OdWEkeWDToM+sJyrtktfDZrpUlSKXp7A+
h98GXdVqPMczJpwTWeLsfG8OH5gpOXhDpjCabTH6W/+cyi9XoaVvL3PobNEZBeY3mCU3LlGYWGt7
y5FW74VMdI5tEWIl21khRItD/Zjf8vyr9kNLasShD7cm/daUunhlG69TCAGKEU5kRIb1oEmpcCIh
y7JR4W3aURu3T8exVKEvpPK/8lZWwTSsgOi/5ioXEpvlf0G/r0FrVlKxpKy2pG86snOHJuAyzKJy
WcGBLHRbpcJJvWWfcdI+K9++WflmNTtzPHW4fjwHVlp1k0aIGjOtvtN6VZrN++TyxNB0eHevMsnM
unHcXG2FhkX4B3mqzHu1f9QkRmmXQIcKXavJQy7AflY/PEBLu52Qr3SaHY0hw3UEUqONnqhY5QyU
mAZWDLuHZxJyxzGO8GdVdKJjwI5DElhs3zkIcr7149Cwp8Svq2/Se8tMW+XTglmIC4o4Y37m6fv9
tyVIpLio4YjF/d3d6k3fyO4QYAd6nkPeDHdNfnaOts7ph9elmAfBoAd113hcBkCzWSWcAvUUNcbx
ZkvaPol6qniQ6I4Jwmuj7YlVhkFXHd7HTI+jehBVV8Hasx+Zz3fKbX/Rv73wl4K8+iPeuaiqKUD3
CNZA1RAtuJi35aMuqFWgWCkfdbowXAIOxC3WCS/v/fuJYh8EzPJoHBJxOcy9m+O6WInTcaHa7GyH
fkZfLhTPkhL8r+CLKlOgAJb9aVEkohKjVtWKW7KZUHDPWKcxYc19StJgmWTSS4ONvAL2zX48N0b6
CBaMQI70GdgAWnhPPUzD6KGA5FSqLHjCyLnM+6ijiEI6l1EgoS87iobRy96i579jcFlW8ptKB4sg
2LibVzCT5AvS89WeMBRbvrYkFsc//+G4Iw3qWLbB6lmsabRPEfX7B3iOBsvRZ7DeG1kHvrn2gJ//
nUFmBm7dib0mhS+Mm6pjt37enQSzhbGlQg70wfRLJePkfe9Oe6DOO9LP+kZ1g2xOtHnXE/B/zvaf
vqLhp6SMahMxH6mD4DQ/qfgUcvTScReCa1QFhaoDXvvaYO8Ted5nOp3EGmLvpcj9fDUwk8JtXkFa
t4Y/mvlABoyUrDmDnAl3IMfc+/0kDwAGdukCm6VRPEnqpPcelouNVR419BcICg59GT/d/lETqfkr
p426iMqsnwOskiGkXvVsKHEtf4zDsrSWOnqWh3lz+h/OGvBy6RDNyHtQtJGdv/JWi6ox+YIYlX9e
cn8Pn0XohcLsZObFcWORwnbrOmcEA2vel2mtXMUhjsLxTq6/wTXLvw2Y0QlLHZtRZh/84RQ9aWXA
qNE+ajIcWubpFTp2NURliYi2B4rww7qaiW4P8QChTQcb/ddeD7i5sxI3LgLWZFA0syCTlJgjU+ma
TT0x5gzpmc0nVDAlu9bEKqnFJxdX64//qxndiE/Tfyg9HZI50doFtv2Achh0D/m5dtXQx9y4aStu
u24qorY/Xd+BH6+GF0tBtvGcDPJz36BP0obXt2O8FvdrYcAPzEoUqzEoGtjDcXalRqxa+HudZgaD
hOnnuvjN9dUom3w2G/QzUhpiOR4gq/fbv9pPQsMxFX5ALVXOlJiOpYsUJ8G47UreBVNU8yh/sW6R
USj3byhK6ferOfuY4Gzx7x19z0SQlYd1x2W7QcG+AFsTY+tO5WeH3ozK4PKzTcejyJxrsoPBV8uU
ciTcRspUJiY+vbFnMW+ObXil7FdKJeq7HyJl035PBO+m+mJC4/507Wc4IUN8yBEVtRJjvBClTATK
P5z3S87Oy2/JDPldMrqzD5OAXaYWHFjQqyYmqAfESZ5AMOM0QPjWorGL1BmyJgIbCG1haLqzHv5A
WUp5++CtKvXjrby1mwy1KnwwywuR88+HToDzoZZNhASKF332a/kNU9zgzrbJ8D3bkupcM13ZMpKi
RPH24BF+5gOqqDrIMeAH4FGf5bePJtBLiS1LFUXuNoyKTJqNvDZeaM3wftMKgptZEnPOMWF/HHuD
u0TgBRE3NH5yRNhN1xyff2si4JWMBNlxAp9C5RDaH5Jev9jwqHe31fBOkEBmVrL8H08Xj8cE0MYk
RBNDBJjQilhSrZ2TxFul+5XYCTozCur2OHKmCBBDtBMfkBNa28jXeTZS3OSOiBfSv4umlYphOcPf
iI4uH/zkW9cGylwVSQhrS4kT1meIo5HmWYVVMWZCOb8vy1VAP73DItOh/1cDk5lJX2/NoXubPcD2
lNAOfuFVMlzOivrCQmdqn2qhWZ365C6uxlpT6ugdJ6QCpkbwVnPBRfQ9eUkdjNisRH1tZSHQSjO9
6vFWza0OQKipOQMkTqt9bLcU8XtBhkIiyqCNMNMITzc4gZIKCSP68/nlzNQmHyanMyrs99AjrMLJ
EybcozdJg1BjCF2J5yRg0dRO/HNq/MEdZP7VbYY49T6f4LvwcWETWpRfJG2dssFcZDf2YFgGM3Lp
m3FewEmtWuIrTjgNSUXKL9MSpoPB3P4B50TzGLA1OwNt7AjLjpCTOyg44i/6mZEsaVua37c3uDj1
9mAFwXNnVBuCPHbFoTcMh1Dz+JDeV94XZdOyrMOXsuRySVNG0gc45kgolRG7I8QfPmPIYjeqbcTI
q9sKbWkfNbBNZPEYs+b7mKYsq2ZDkDkcpPKfyKVBb333OYxsUSFhWDuPPwXfvAZgVdm+SQ7/3I0B
FHFCHg1/x+eXqFvQl8Ze6BEoCMXTxmlKInFCU130eloMy1LcnR9uByLg+kihb6JxUo+Zue5D5rUB
MX9CnVWXCUaE96k0sv146BlZPyeMv2AUYuZ1AoIijIUK1vuzvPveTtwjOLx3LHWNarait6pPJ9hF
3JL2p0b/96+AzYqylCwxpuwAPDMp9oACZ4RBEhoROUS4d55p88my5e2/CgfMnI2vL36qCKkVVY6i
DU8JlzIWlUJ02pchF98KiLeTmkwMB/6VnKSq+GLXR8HSUGhtI3+M1nsytQI3I1TVzbj4bULZRkX7
uQHywZ+KFo/2Lf9wDUEw289PfqpsoZTNrPpZpFO+T49nhbNYjRM+sml4bCw8+aWhqnxnhOr6d0Nk
6r7UAA/LHazQqoZmr0S8vRCNRvwKP/vKhib5SAq/XcpnFuhCHdgFswPicY4Uf2TN8CMX49aj4BVM
JTUqw7RtIsGiPSdtVR7MWP0mP2qUg3ZBFECnN0xJZ1TTfL13oFjFeo2+ZlZxGhmPwMnO6Q3sDkzy
4aFzTIoZl5XwF9sfDhHINXeLS3Hw6ab81+Rn7v93dRz1OqD6QW8W+hjTvJxId8/9MqCrdmHQzn9t
04CF6mU4VZOYZLpyt6yy4/CJlbrhIuLeZayJs5BFcvBCFLkvUu6CXkXR+0Da5U2elZARq/668JCu
CXYrbQa/51/+MHEF7nBRIvkZ0t5e17judfsJbgxl355CUs9TYNkyYQ8G7+Mi+ztTVzRf857h6buy
+noCBQK/H2CqpBWznrCBAETrG9qj7vGD5FL4jwr+HcIxjBTcvsAg+VLRM2/9tb+RfghcEzSAsKWv
Y2XbdTSZxItn+5xWCHcSE/o4FVVc6bzB+q5/vXfbviH/dhUXQ1lGbIGusljddbryHOJTPLZlVb5j
kO/RZFDgF23USmVa8eU5PCyDToXI2WHjdLff9BIAeIfGxgh4tM4+vTGG6NVx8YCEFSRDxjMm+GYM
zjOBvJQ0I6U+KYDplFsVYNrD4uQoPngaAZ8oUAmdPLWh4rEPHIQ8ZBmlapz2PUimWbCty6OvEv/k
n9TTwX5WRB4Fl4qX5E9UnFJ8jlYGRrzVN4WXj4Qf8abWyTeooevioLGd786rRiKTmGiScyYrRL/U
TIriMcFgtXQnNVkgcgkEq4HOXiDG9fq/nAeY9sE6Nn3Ga8o26MRcBE+QDvZYsi6qwtzaMSPPKXy6
QZFWeHzX7qVZ12k9Rg4qKYjCeZ88l0Azzu+9OXbgKkAXIAhAfipDMA82L6CRgRGLvgktomF/PMHg
SPiEpfRzRdrAwhYgX4K8MGj39haLz+ET5nWqKqSvfpVAHbR6tW474+6LvbyhZl1N3kXe8eDzVjqC
j0Y/kHghiAmERvIcFXXH6cCD5vWSIJ8tnHTpc+R0qGIjKhBKTIxNKJVEEzJVEPU8KisYYiD0Kgqx
EkQtluR8vZC1QvyTnjcC09XjLNVypzhBnWPz5xu9duuSTVj40eYZK35nEdoyu3stzYTLYg/ghd4m
Bhag1w7gG4fHh6SPTnOa3nFAM1poPGXU4gptBWNNeNcjcvNS+mhOvvqZBvr7KHrO9rTWnj9OZi8M
n21dCEJWEionymJ3HPVSlpk0MbdW2cxiutVN2XNG7CD34pIltLr2IOmd5OxWVPf9VXNbs4s5ggcW
dRYOXPNGXfe27SUJXwqgRCJ86Uc/A0p5eLLeQOJD5TgZgbKc2bVnmc6XsqszkgbKhVIMsHRq19sG
VE0yaERWxzCzGcEwoqUugAeoggdlhctFfYh42IMXOp2cP83gm5hTcnQoYMLxzw6GA2z1dvx36KUz
ONPGr7ewUdKiZBuSmg6/djcl7GJUKY3gHE2b6nDWinLLi3S2DAag2woMJsrWs642IYGEqSflOxPw
XsBUfBTopxsrLwwblfJarcm4jpemSJ11QNqhaWtUdVclS9Y1tDZ9iGMtXDE+r6Y+ZIlcYQsCZC6S
2iY5lkcuU/Ozrw2mFaQIFEiUh+M7dcbdv19fajEIGl/NWaDfaPRtHSROt2iR7xGzamgvQypqWfIF
fATHl9gOSUy2b0V9QLK2H+S5FTGAKgcP7t1h6tpIeQzbDrgV+M1BAjnLmvFokioRyN1Thc8A4AcO
cFMbzZY3x2DaKD/wX7+HBu2Z6RSNGBTQdeaVU23HgPzURqwZCGoRofwtnCizmhNUGv+6Suf5hl9Y
RTIqTdXTlIBAYUGzwJLOQGYe3rihrHnYrsnDoCmUynW/1toQGU6pYprFbQIrRdeIyiTFlBscS8yQ
pZHdTGClxz8UYaQQ9ACB6V6U7ew8a67/VXc5P4Dh90QP+vcweHmyhiQAmmlrdn2zNf60iy07P1xX
yxGR1UKsCnQcwr1tP3rza3SH43RLalM00G1HxnPhd8ETbORhMa9/EI6fwjt2x+y1y5mqqOuYlccK
hnNfsCRAzI8UxDhDWTXLmT29AQlhZVnzm/YfgY1n+4iNkdOTwkjTOWEpExU8xiqG0PAIskKur868
w6qXxNLUzX0msmDjhlYXbvEm9UJuHoIayc5nUizaIZ8MT83duDxmFpG90UgGifI63zKsDOyHeaDX
tcueykYlkyXqbtkClPmlwhuSgHllrbrHc/eR5Tkb18Xb5EwBJVmbjqMBc/OuB9fByrgsenrROhGo
Kww8zhQ5N/FfDqPPk1QXVfj9I0y2HOtSEQpPAoyfuThK8EVovLoENfgAmsRWXx9CNrA3Y+lbnmD0
oHrrm9yYU5l7Ja7J5j+qsEVKVA/9w8qUgk8Eurby2gXuW/XMOkmVkU94tnLGKYj7ObaczLuxdZVQ
yZSEMfRLljQ2BN/XqrUQhLejJRmW0GAsHnrGUJOyf1w893aoYvd/4yF1GV6w7Ez2INM8udIOaqJd
vCAuRUFOblGuxvxUPT+2dygNV/KzfTy6OU8zrqeCWLZAy9D0p0rdIzCkkedC9tEAaocJAnoJ1fGK
69dVdALrDSYC0/2dWY5mMs6sOItgVpGNTPiX+D29S0jf0kFp42b7I5PoiyIV2NmtbBkIi9Zg1fep
s/NbCs9xNEP3343KFTd+0dXhVlEWpOSHPEsUXJpcdMMDWlm95BlW0mWaRnJkdemb+BmA15Uq+sY9
9/8egHY6bx12Zm1wGP097Hak96g67WPazWilagOjUM78mRUsUfK57CFliaLT+qCZ4QY+XriXmOMR
CIhpUm13VJz0dqW9bQ7kVbljwa9clVe1/r+n9wW5mQpCCBnQ8k144m/jVL+OF/lQi9qIV7Drztd5
cxaeI02NmIAzsyQVmn03ezYuj8NnXCNJAPucLMXr0J5mFaExKdC9z2iXTEa4Oi5CyS4iHkdq3W8g
k7KCezIHFqXxoqyRXNNFktbWgRTRZkjibeIP9luezQTtGCrob26nW08WinEnfJqRCn49vlWUA2IZ
Jpfn8scru/l1t8CGPDY/QjIZS4HJJ+MtlKtnPGhTKjiL3oEO5eKIFGES5iviG84Gofmgy28kD0Ji
ALWTY60e/7tUZru87+vBaDctYKeQbhsDlUVDhGUi526kwh7vqJj3Y/K1CgY2u53NKiO54CumSjhv
Y3c7c5VFOez5W5g62UhpA0HEqunYJPoqOZ1hQ1NkLb8SqYT66jCnf23fGGz5KzvpAD6byaK9EFrj
KTI3cwqDh7ee4oZyQDSvBKc8nvsC3Tx9g/LUiZ1n0JgUn0Zzh9sP9MshYDCkCx19n82lStPU8cXV
7xnH05lRldCs9m+DFFD4R4FmvWgP6x+39a9Too0ySharF/6cy/q5pZDwMSIbED9bOt906Eaoxs+M
96krz2qHrolLLWJQPxULnUePyQep21+oSAWfLHulLRGi57TiGGeY4ujDOKR2d7DHgKW0TMGEkS2v
Bx/75pxnZMMVYZizu3V1rFnqZYcw/UxGJTyckhUMBkiEZ0e+/7WNbTcz1fv/+E0JtC37QxWcGDh4
kZq0dOPLIsr81zBdiAHZKh9JsFwyHBLj57RQ2IV8WW/1TKSuZxW0Fb8EFO16H4PUcsV5NKTuaGZF
kTEgBtIb+SxhxlvpojexI+gR2FoEMasPm4+kMrY+XmMXFIFAALrE4vTTTD1nXa9eSJtPlItOH3ML
3vyIIoT1+aoQXMOl6yzSb9wJYp0rmEoEmjdoDZGyEIPLw2QgXB8hMpYhYPOzeTrGCd+e1o65SWpG
ZEzzMD1dnjFjvoH7gx48oOr0G2bAEb8Vk6788xvP84bKOd0+IRsB3bcn11K8bYs9zyTOWUh1df8M
4ZjwLHktEC+8VvG8h/yvTC6Y1jS1mbcp2S1qIphpnSocaiu2FxNATdQQmf5Fypf29OCJ6GH4e77Q
lFzIOIsT8dJXBzRKVuibJpl8JH31vJWlpao10sNs4hQYoGj2oC6DWKY9Rf+yjr1RDAe2ap81zFgQ
VgyzJZwDrPa+Z6Z4qkKSUx7RW8REiGFcwkFioezBfFfuE8wt12wgbC8RaOEx6DwPxpVLRBxg1MCE
6UHt/AlHyg+mGmXiWyqs/g9npnITspRtyUFT/d7BmNkm+UXvqOmC7cEiuRrx2mqBPUU4YnVlpSen
nFKkFuvD8aFqKEUZaw+JAhW5hPWcv09ekOzDmurK+PXUGCsQNGlLM/C3Qz1mGbk395wm6CO5LOCl
9YQNn7m0TELjaRyywOk4h6nifXAeDJ7tFjYjLNuMa/0+EWehDSUR4/3dYxTNltz1fNBb0bgBvc3b
ddNFtEMo5V2WF0z5QkKBSAYekkBJhQpN0+Itmjo30SKznDmIIl6vNgx8YzZ+AcvC8sb5YWtGcMLD
yfA6To1mo/H2sii63RYWNc0Pqa0df6t5TDMLkHZGneAMY/abNnzHlxdMgDNwuQxflK76relCVMIw
e2livFtd1GafGfCmEJ1AN/pj2jh1yNuwN9ERa5UNVgqZF163fvxhO13qVvlDcUNqjqCz/eXA2bJi
dL3UpNQQCrvUmvjjkU2salr63o2kqMgnSjUPbgc4LsNE7UP9oKHg9+58gsltGISHDm1LA3++BrPK
VgxZH84wZcIGBp54fHFpS1ccjqJ8+PUM2O6Q65ip6wtgebSv/hqYMKPaJVgHuBVq2/Z9ftupGDOs
k8CQ6XG4ogVOSWpyGAVgH9gmW44hlrbuPlH9+RTWvs+xvGmAOFFlz8f9fY+AFXI9qvOWzJxUu1Wm
9G3aLw541DpWqbDFuRn7rr9XyhsZxLkzzp35NItYQB62zMO+lOEjq1zM8AgWz+ooBMAa8fKkDWu5
Zhq1X2Zcs91rtW4f57iBJG9GCg4w48jFgYGwOnyX4gG+EPOBJyMv9p4btgnE4OMGdUDKxjJIZUov
e9ciHGPDJ6FjirjV58GoaAbUULKI0mBXObnvVrDHj6CMIxbhucZJXmxOcov53foGY42y+xueWGEB
IxCZo9N/UvNKvupA9uMvzrevJjWFgX+9GQTffGuLoQ5gZWfaLRjTeEt9zjgJswb1GV9yLlYsbLTY
0AtxN2rq2pQe4bRTIw75vr2K3pdoZn4crAkTekQSRrg/8tBXRs9l+c1dwrjAcX3BBZRaNLLyeKzW
Es7MDfAg1xYeXNaUfK83le5PjdU7U2Ijtp3XGXH0JY5OrBhHPb2BH4bEYo9h6zjNfMCFV9wYP4UG
rU8+J30hUh1rg7mMSjGAa6YmYsqjo/2MVCcg9DKBlnj3tW6lUk9z24/uz5EhatDbiVB94V6lnbgM
a0Hs+4/uQ8FcTNq48hK85N6Q2ursmSziPw3UWE7xIVcbmu870HZoJNZA9Qm2GNy91CwOCtuLI1C3
yT7WQxJYsrDxNT+h6mN7qPCU2fxA99MXPDOxHxC7QHxwhzkDaoSjbdYtZLWAAnozeclAQw787qgC
GhRpBukUIJhhWoTMs7MlQ6wEcmO0eEwdiWbA9U+R63FH3EK0aZAYcfLIXzsF4WaaI3+h+DKssXTt
EWhxUbCYthIRxyDUN7U0qlab/XDsKsGQxJX1zZlmcfyOBXojW1sUW4uyeMDE57xExjE/LHM3j+Ys
/oBgHNSlQscXN5CePjZje22k1eZEURSf2HNX5Hu7G9CVsMDMTBlrPCWHAhltFGUIB5qTDxGLlHAJ
K5PLvQ5eiv6gOLc2jlXi/JhsQzXb4pmZKbpS7LlTtDuE70FxPfsr5y+VPxvY/NJr13F3n6jhXii5
c7idAUoVUNmzze9kz8FoMPlnk0uzTQE4u+XpXi+cIXZFkXbWfxIW43i/TVuiBSJ+qjCYZol66JEh
lv/EaNPGoDj0wOU1LpqbADtXS00hU2T5nCxydgZV6VSgEWM/T7JRIXpJJ4M6aVRhh68oMxKMD4si
I/IXpwEO/g7UhxhFVy8TO0+OnITIBaaPUo586rS5iGEkH6AhGHy94+xhlYhkgGYMUYVHJxvSpnsR
eZhiP1xn0yUKwwgx5laIgWvIdqiyPLedr+9SGTq7O8jDOu2mSV4SKFA/PLSzY2VKi0R/VVSuZ7/0
YCpTf76ZG+HH4RW2bnXJlGIPbxR+lbeS323QFVrt/prey+l85FuOgF9OyINlDhBj91OBUDq81yNs
Ai+snOzuGshXeMAlzgFvIAZRUPLMHZoONpEpDWPXdCg/XgTiM1NvFNSZ5PTLHqo0mbFyGKLludj+
iFZv8LMIUDvQ5vzQb8rKK1O9oaVGK/Y6s35EMVgM4WnzRtOo44VKT5Z0HcCdTjwvVCTfHiNY1mUP
pZEKCjBvfrBfP7kngImLYEOe0DRVa9hY3nIcY3Qa4+0rcylvm8s6QvAOO8YDz9i4siWp5W25P4zj
x+L+k35xyCQbiQVaj+vmmsn9YZtg42eFlc3zeHCgGgvvlYzTuCCBOX3mPphICMXUd9UASec77pmE
4pccZZsLrDr15hx9kZGQ4rQNfSmuNGdmiLcXbe/ULJNR9gbS/sSU7RJrRs/OtqK7LDURw2+8tdXt
mIoHwie4Zvv3VxB3hUgjAUCQUnqznW7Ea1KSMIApm6JKBTH4dcQREcPkoLyDD9u5u0pEaCw9Nmqu
8z5fRsBTr+aQG7YymTR7G9Q0AF6HUgSeVR6Dw/lLzQPnxTt/weIVPMvIe3FjTnwtTPfMo3Z1Uojn
HlvfZdTLuJiM6ihrfQAc5bU03v4wMKzwHgHfWa7Jb9/Py54mtFiBXOYh9FGzPwU7ixaAXfjN2qQU
XejRvrRlpJ0mBbXUCner80WpjNPQV7XTlAOIoueGJJrq2c+ynh4yiuMBl/b6wQnHD6qXXlQwUVtY
M2xB8YqshM5xXkI/v9GdRTEwYK9mE0LM66ifqcSoqRyjqWCBsNl1115Y8jrcLab1d3w5NJb0l6vN
4eG9w/5eiaUubSRVHLU/McGO9qPKgex2H6IpM80UIVnDstWPnRo5DSvxfbsxvQMIkIcETUE/xA6b
1STQrCjqp+3gbdMFYdrfDOkSxHe54OoYzz32COUQB7pY44mhNcaNbj5WOB7C/ndboedWXnpoOrF8
Kcz2rIcuOqPW/4ZK3dVI2VLxF2kbpknfRi1PYVbYRW1dQN1UZIi5A/IZug1SXzYqQUbkN3zbpGeK
PbfcsDTBQAkVwWnRS0M6r3D739Y9AxAOzxCaSuOZ2pKHjrGSs6ePntRDnStwnDyhTWLZrkwDZvP/
LRTjNJe+Bejkhm50bhoKa3vHaz33udS0c8YaaRZzMjBGgrpZLcaTsgF4Kgte0PdjCRGmxI1R0o3W
+hRB+692mWEgJBPcizE7xV+X7MzojTl795j7E1n/pUfyFCLZ6JimO+yeAaSUuYIwMY51EWiTBLDO
5PeJfJEm0Jje0NcfFNeA+bRcDWjbTDLETF2V9TLJeWmxji/JJYJEsqGsAURpQhQZ1I3TKUygqE0T
UDFvVJaZ8C0Mq3RQt3UrzZOmCPeJCNuswEHE8pJEbm3vp4nOXfbOgOg8lTXayuEQvVkzkkAFK4HV
3PXdZ/MADYQftsF7CAZ8nocWwRZgaTGU1At8dpA6Mj6S8//DqJEQnf4J8A22MPbeKO9bOVBUdR7/
5h4JU8K0/wU/vGKG05MkPGHo9D+C2xlAyrraOsoI31L641tEs78fH+C+x5wqgjdZDHuFO56InUWw
WgJ03ILfmuXTzlxhUzL3/WO78cRdatvWnhOX4CGc/B+ne7W1VXy0CJSzq5ME8YD0MhL4Ymz3Lety
puPN2gUKg7bCa+4/8Q14Lx2gD+psSH5Gel4vI/ZeP/JSudG8b7cuxuIGQk9kveK5fpGvGfeeYYHa
6azC0aSBxUtyyalv3QJmIZKcQpl7Eik+1ikgSO6O1nr09Ic2mbALW/lHk8ZC4rquKFQkCXc8fK3z
djcC3yiBKQM8P8pzLX9y2U7FaYzz567JJejoN7zha9rnLlTtftkiQze7IIltLzCe02lhb5qKfPxg
PHJfy3laGX1AicsrDfiFvlzIWXH/SVNQKxh2upbyQD4HEvZ2Kkct7yJ53cyTlnHrMu2ia9XuJB0Z
mWSUY/vv8qTQ0Fp5MSFmP1KIQCmJVSAATj8sKvpT0j+83fEelESR+rKR0ek1xajfsgmpelzAer0a
owW+7P/2TRLlgFQH5FNwOjBmm6rKq/+vvlEEkR2zLQh/ukP+/bRcDQ+APGlsLUmwfagRw9RZiVbl
olJHUFlKB1dvwLkHGmY9sq54GtssuVSF2XvEWEPQ8Nms4kJmaWs4z0tTgWVrbrPaOJsZ8SMxXpt9
ePhRqje5TKgBOqCTUKOFz+aGRg0OSZ1sKXQkKVFZUoNUlOZL1GW7i12r13ClHCb+WZPH75R9G+wU
EJH3x22qzUmSY6AndzHmnGJZobi7Unce9isi+q6XbuFXN0NOh7N6W5AiluBcfpQdJUdoW2n3FrHP
qTC9og8NVNVJDrpEWcq2nx7oFkyj4Z5dfm+1/G+38tfSQYHKjtjmIpC9cnxSFrYtJtCI71oeMBHn
fiwuewfVoOi8lFx56yqPXe/NwRb0AyD2MCjf1s2hxAGIJKbDmYuF2w8g4uOg93NJWZdJIaheyoy9
c6d0yVw0Eqa6Z5yX0PzU5mnXyfOkU0y6jLcq+PwNsqZVreE7fVxe2S3NxgM+ZxF541ggJiQnxfzr
Ykwy9ZYZwnMU/aDTpyQ7cQKLgmaO0wXAysHQd9cIc27jBcaE5hmH6qZ6W+EegsnwDFRZqZnlzLvW
0g6INiUcZwlawmHMItvaByh+0bgSGucEhboKuFtThy/CDe8C0pCDtc0rC9L/fMeCAOv3ocoEdQux
YrUkM/SpAfR07A8rgGmDl6kB31Q70y7PjN2FNN8hthfT8QWBRMsAxpFLgfNUNG8RiIGck0yuaDb0
kM/DefVLydga3r8g/VSqdRXp8WKz1IxkhzlP13XEwr8I6BXVnMyHw7PGoYcY/C+IxZzH4oenYX9Q
HZfm6eGjb9O8KWHXIOSnVNJgN7Cg5Xop+3W3u2QdPXmNHkrzhoGGH22SF4j2hDdsF33Kxp0XMSuo
nQ2+M28s3yC486Rlkb0Mos/Wly3GZtlHFn+5sDWrxAvyZ6i7lZqz42sdD1fe/24bZzpX6ddthNIK
Os+0YQhXhhYohVXlULxAysCwrvFrn9s+YYXyZmvo9NZ1HMWWphUWse+xFpczEM3SXSD/JV84OCff
8nCRGq6TPXcIN+CxYvqp/nKXZroBK1jrNMti1EOehK2DJZrq4bNNwXlg8Wzk4XC6+ITylFBEoPAc
jQkyOI+lL7sx/IK9Lv9XRJ3GrBOSwLex67nekO9LgrQ5CotjutJg97xJ+IuWF5GoQ/2U6O/d/jXY
D9FE5sXsdV64JxFnrZRIh7uwhhEE5G4wxB+icIZGSaRE3mLNRZzSC85gtvPNujmugztSs++VGGMs
6Js+KMRjs33x3SdnQy9VBHmZ1cdz7VaTyrnRUfC24V0S9pFIPfwYOCqcQHMpDqH85fa+TMsc83zG
BRu0t5+wvnUqW04tPYM+F6xCt14Yxqul6Etf9IE5aDFhRCdzE5kDomc28+uVDwe809fedCe0b6CF
7YuhKrSbsFoBXZhVEEjYYb6g7NIyDtQuXdvGkodsY3E7sJtRJh9Gw7bIYVHpT4AQY5L6Bj2WfMkF
FvG4o4tHm+okHahphtPvSPTwkbEDUGY5yZdONXS2tizX8siGxXdZNmGNxjz+Zdg9qzpdZXanfffk
4njRifRSyMShhD9CR+4HzZV4swsM3JoJbZ6THnTJD+q9r1k3thRRh9nzkPVK3ijhaxOP+6q2YmbL
EcAkwiS31Hs6tPLd50oK4G0FIOxH61ys0YhtqFeynw8XPUBg/bKGzaZJEYbswpar9+gbFn3QdIsN
mRyIS/M93l3JY9elABkFrlgMT9gUAe6640zxeOmVpvTm/5vw3HL8M1P2mdqRmwNDK5/Tdmgr3RvX
Gs+JzpLPnNZ6TVbOxomBAiJy9sG6oHtQbiZY372iOP0C9KTfgyD7FpyB+jKFQ2ePnd0dxidxGYwv
fl2jgK/bwln5Jz2j03pxpLmwCAqNWPsXsiJPG3rh/5lhRiJ2DLdBEbjF+nQEj5HdqZcqs8y8ohmj
d8dOlR1b0Drh+T/0zGJbAvu61M6QjC314pC/3AjFlBR8nb8rPhMEMj7DSct6bSfwvHhaEaTviZre
XK1xjlt900teQGtJOyX8IiDmXIknXBNT9vLd2CsKI6y9fth9XxYc5bwbg/Xxdm9AwR+qjCvB17nf
Rak+VmWM0DFOdUm1fXNOBSHhP+KfXkzmH5fdXh2rhhKSIameRDCfnsTrspweszi5aKBzThqnh7fr
/B8fKec+6XYSsKXi6cwO7cl++e2Zb0MxKqBWjYb8YzLzR9jkaYpwDG84l6aZD1lkdUNF1lSltpE5
WwhIlWGz3HlTXIPKtmUGZZ+aRxGKfnLM1V0PTaclrIdMUVDE8hN3zRHefdd3wJm6PGGmCvi91Sgy
EfINrSCD2iuQ3qKWpa4KrZxYIkDUTHv1BpQ46kmju0WabfuzIkcypq8uXykvaK4B/VwQ/FCpOL7G
X1upyFKg/F9veYWyssqso6qf0+UF6/8c/h3i0JPEDdYO0b9khw6/g0fuD3UgK53gdxh58JvRxGVy
DPCNluxyIKCSjSaDVH/UdlgyiOSk2NgvX6bmvIIJfYGdhdSKQeVqOigbUpPP088vXDvFyVgVMmmW
WmVIjutXpNL06UpFZ74zWRCepbruC/G9pJa3KqO4aMj8AAZ4Ree/TVbApxlQMphXDACpnMIbbqWN
JawBGl2ZKQ0F+6sODmCKoZW0ZyVnlCbXBqJw0rxHFf/qtTJsJ2Gy0SgZJpzXK06zaOE2YHFsmXun
cuh8vC7QPpVMOgMa26t9yNYrSG8k782ec3Df6NH+U4gX9jiHfGPIBWxD5VDXMgBRi/Q0necDCU1c
bEoFioqHfZAE/UUnS4nhAszwuhCjkGpC1NAhG+8yTGytBVM8LeGee8FUAZoLBJEozuvsN9hZKH08
zprW5qaJaxTamqcCM1Qf6yLHpfcXzX/VGu2BSBfjSsnNhs00I6RqvW+58czf6C1rqsoK6ZdPiBad
76b4Bm8baVN3L9d5BcH4miiB6HL2s0ANKEZ2bownmZtENMWRdPtv7JjGHiK7PpUtlOyESj0pj0XU
b8pzPDw0IXYXCd53F5qG9xjO6jUxRfrkbl1INixmo5uQhxSQQLj/Cb2v0uKhG140CrC2ipOWBotR
qU/rAVxquzXfNTN2Md10f0D/EsTE0Drx6/3+Mr+S9hrq8mCzYvcVjPnPvYWrRDMKS+7OaO/vQ0Mx
1TOCyYM+ox0VweCVKR+pgPj1nUbszLJAGI9ha5xpFZ1u2YjL7F1DDazu01WQhEnVKCCA6KSN7on/
5HVDwrX7H5cJcEpIpuiC/eTm7bkwV4YnaLOUSqfQ6FhjTQXh2HQ/NUiwjqEE0cNstyGOxzQyk+PP
7pGRJmv9J356WQ1LbhOIbq2iCkB+fjvuJqW0hWEGYgp3vvjzHYQe6esPO9QFaIpjQGEZMe5c6U2k
vsVunWHt44iSMG3x5ZZ2oVvOL0h3soWR+WxfOazehbEpQJqonIEBYKTUeiP8ct2HVWVJNIdZT2Yd
qW0DXfl0SZgnkkGhuuKEdxgIwHaMXCgODjoCpLlgsi0HgMO/2wWmdFMx7I8oBxBSaiWffnIYl+W9
RBlV7uft0Z6iABntVJNUw/qxx5F9PDTR7jJrcwZsjtFwMmc3n5+txKDgz15XJDAYiUxovYOUBLda
946ZSpzlLJi449dPySvWy/eG+AxiMTSkrLy/7cU4FKpSZHevgZKe7+5A9BhiXe52QQQDPytcjL3C
AZXboSU/BqYTa9TFf/11GUAJlaTOHz42mGdYO0Yn6UB5he1MdAA3tzW+KdKQaCm9+LToobZ/xYFu
VNxnOaAhCBmPgeIEiFRmpWT1vqwq6Fv0wxQGDLKDhIstR1y521SNQBDpBV8RdFDHN0COUUHZa/90
CnNXPGGetmdODUMBPB7WuRNwJEGB9qZrJAxMtz6y/voqd7TC+mzI+VxsGZNJqQYiSQU2Aw8N1U/1
pivrMVRsWCkslR9Fh9gdiqUV/Z7VNBIyhNfdfsIBe4qqV0i33wZVBdgBHnWIdX1Mbq7voer1s1rp
83ouzE7JFaC64/gVT8+ZpnKIqXJMVVS58Gpm+gP+TJduAMUIYtPDZtPnjyJkYa2WQ/B1/mXeZEb0
HLbQZDj/PK4peRx0RLEHu+LydXM0JuZ/pgGNJasRN5TRxK//x26aoompWnTJkkY2AuVEU3XUTJlo
QM911PUu3N+AdhFxXQE+Dnq2kZWkCv5qxlujVG3ulx8PyASm6V8TVti1QGW6DM3iXuwp3UgdJBhI
Ril7avDiQyoaWE8UmeKOdlQjzej9S/g+9+B2oyiKCXF0BpCoRIC0r4eq5KE45uBnQWu/fABBRLad
wZvUQ8sUL5FFQdjMCs9ds8Jz5YC2YWEmMA0ZqExLAbCaHStSHe/V0Euf4m7NM90ljNrSQ0IgDryO
f6ZVba3cJ3S+iEvY8eLNyxPf7mh71jb8RKoKQGBdFz/xgFvYCUnytt/XDcoGek6C3r3stQQ+Xs4y
R7bFh0P5ch6EiGp3b2ZFmV21QuHGgnv4BCjMFywdj34irKDMe4zcXL7lhKPE/Akn54FXPDajyKYu
g/9uZtTMhChvfrgUEdtwiuv4or062cdfbTlwwAUNd+1bIWslPlD4S3Fvg7THy6JQ3058oOQ/TFO0
Jv6UKWcEF0OxktwenaeFppl+GYIIbqJpLP3A+ugqi57IGaOsJ+pgn7zkH7qx4hR66GEdFeg9fcIA
b8zvW9u2uj4HNr3y3lrpZhZwXdevmlN6IvRmKRoO/13DH1vlqiEJ5LrpqCwagt7nkiB4TtLwd9pW
Yp4Xgn6XHSdGNGsjTnMb5Aip6dyfmbbFMgvsATNmQb8wV3P1Nyx8Q9acD+sjjguxWtEsquZE5vxU
T83ndBThMl9MbYmHyPLndDSi1iSb6JL7MkBan+vs11hZoI/XcVQVpM38kv4edLH2e2YsCSaD1Sxx
IhJDKXv00hyE9lLXtlXQUtSh2jY/5MM4OLBeE/bGWG6+7zirLyNSJ3XZpSszZ2N/VZPBsoho43ps
jQoudZA/TzvFEh2Ky+tEsL8/Y0ApObW3p9NkzJfZnh7uq2vg904S+dgtN7qsDva4YoaceyKzXDM4
JAeZYprF8vdsGl85vrIfxyqp8VSYVE/w+tUUqXhl8JdYT9cljlTtQRPltQAE7i6lgqXyYktnIzHL
vkjWk0UQ4qvMsfxD5ihvw8uwRLwhqz91fhlYXwDH0pYbi0QCfs9Gikr2919DCkh1JdjjT9HaqCcs
jwa9VUnUYI6GHEI+h7GnC0oHIvDQgG58xnlfQHFLjBJt72hLM3Y3NHaCceN5/Gae/7RwsSLfMZFy
QXmnOIkiU0iblebcjjaviwMKabsKfvEUyr7Mr80KfYr5vAxWWOIHbXWi6dSg2cl2Gr+mZAnchd/r
JCr0UA+Qy0gRfDpQei2NMW44ISgdkS3/B2HZDYNIJug57JmeLWqszUDmggWyDzR2Mx6JQJLw1yEL
N7qXxxv00iqcST9DKbCpGXLU01BqjJ5XZhiRYtMW1Fwik7RWj+gzTXC7Q5X/H0BvI4i1X7Y6mkVe
4lDRRh4sOhUxvV8PdQKWd5psQBJ21FjCowDXRm3GnHoMKQci8potkWXJ1E1wzoTcKHRw162DP5/t
zv/SWbkxsNlw2JV9oaOt5DTtUDeTN8OPhR3Sw+MLidllIIBzjQzvMdpGVeKMOGihg4p5Af2X1J+j
DFweNitsDcwpg7Rqq+K7/Uh8FlvUjYKxJlgwF1HStC2fgaJZ4poFG06Uu0X46nqc+EXY5u5927PK
YF4skCcgZQCG0ITE43IIzR3gZuIL6a6dHDuRuVIPp30cv9keOAtsrqqiu6RWDCcWN3fHtb5lIzvf
zNflwe2d940ijtqYxj7C3nbkJB1grbGr0sPfwZakk9cr2wu0jwJDUSKYU8crb1mibPj3D+J5NPaq
W3RGi4Dt0u0kDrk7CfpFEwvnoOtCAYi9ZknpAP+jiwv/q65llwIefeQXuDnJNdmbOtY4eu/IV4GR
nhrnqXlCc4UAoQSoBbKOwTc5Iqh5BBc+rAV0MhQG944/Goy4JzKOo8ntocKM8cBN+PjFdKnIVkH3
PM8WaXW9Ro/BIZRvBmJeHRHn6YDVmk5fqA/ucEVcihpCXs6bVk7YO08MEubH4/DAfMnFV8AyhLi/
YUZYhthpoiq1XjAO5DCaePCAj/Klz9JbkG9Qt7prOLUW2J0Ru0S0thcYzTnyLxYTEVvhfF0jYdLZ
Ki5IsE9IzaENFI/6HFCMSSbxk2qgRIVtmbHFYsMkhRnL0B013iPYWy39F1EsFfFqZK+CU0RYp318
6X+ZZWotT+1BI7gL6XfteYhIKQku9LH40ZwvJrmMoXqZS0gnOIPd2Z82T10y8RzV3Xt8GrephSPD
cdPakXay+s+71uLrnrZI13pcilWWaMwt8DE+P+Y7KVtO2PY8D/m8iJsr8i81vhlEDykA0k7VT4AD
21js5w32Cax3KI1/SyUETX0P4q/4G+UEp3d2J8Fz12BR2lwKM+lkM4rA7hKtCQjmdCv6e6JF7q2A
cyXzHJ/FaLEHlkabndpXwyRWMDVvwqll4yCfmwWz+wlpisKazyvNmL433cBrmXpP+df71QI/nsnI
k0+im7GzPdZHmmYgdacu5fGRfIslrYRdXhXzyukXvCxBgh4dYkMAlM9vQHxIeFjt+elDK1zyHiHP
giDHRIJIK0EKX4967TTF7fRQxRHj0tQSKhEbr+sPA2sEXYSYuxu2LE/xWpF1em7MoKF+tTGAq3QO
+IoRqR4EcBIC51pXgCuEYw3uzY+qg35AulfcS7tZdB7wmqgiOqzboYczRIrLQ/WczgqEb6cVhmn8
6NPhN5e3pQWNNZdUNld71yJYFqXDzntdghRXSq9pTmkuf2LXJHuWu14x5vcwcA1tsUxHuUL6Yx16
/r5U99jSGCwV8HXFE8/tj8DppowVCYDVlb8M92mG5xMCqJJuDL3eGJh3Iy2xU0hKcgVHOIxfvijj
Ok1DZNN9ZcxZKXIOTU1CVg6P3gJfLp8SGBZtS9Yz04ZZ8rMQDyzEIsB/FEHgXDL1yRwZKILCl8qQ
lidwbriPOPj3fE2YXCWqw9ux5W3G8x0Yn7COm/l4XkNiNTSizdHqW0mXWUOqlS95g0NYbtItjNBQ
woWADlFjnrEv30XQ1ntLT5G/NGycck5nt4M4x+NozM+k9KFTyf0mBSoV0ifUn6wuMTpCs8vfqjYR
yGaQYETLo5jYEPnDA7VtA+O6lq5VNaxsXqN7t2i1Xs8HO0ScPAZzN65Rh3/IRHULLwRiguMY3Nzu
lAd6QCu3fquI1jRI/GK92+sZ3iaUc0nTD9f7KvrOcVbNgEoK5OBfZN98VnwNF5rxSX0X5GB6Alds
dFkLJ9ECwoF4Hb2nhjzuu97A5bcrb4H2lVD/BXauXH6QmmQeslMmLJWulMsKM6ALlkduTRYjwhwv
aRepNkMuZ7MytxtNbZxViEr2l3ISOSIqocBLCGnTjKVNrDrcWzg8XCePNv9z9j93Z4LzT2PJkfix
IVW3s4wcLvwKKnblrfYVT108gWevM55b/ihPO/aJHsnk3LbXHFtpXl312QuvqfnSqRU7l8Osxamv
7SQsr9eR5c+NORZxkf/sWm3trHDvtWwulMLbNBEgYFAacR+phciadoVRbdMQmv3vOt+BMi/nSEjd
fMG0ZWHjZEJSs2dunkFV7znYOgySQfC8+RpeVwC3bCeBqgR36O+O2WP9VWPhTrNUsIw91ho7881a
f9wuh/CvRs6W0M7A0x+/j4FCXuwuzzWjZoaQN98gHhw/FdnfuElMWfminyGta++WZs7aBThX/1in
RUyzAnIDrzCBSlBZr4Pw1/XOofkuQ8cW1jWAIXFOAE1+0b3+1bQRVUIzW0fUk36PsmhSINJj7TLG
XVE3RjKGTL6yLB1pmWdIQj5XcyGqv2+fFTUemDa5z+we9liJW3rB+QEVfhUVa214FfET1CGesEuc
LCjxU30H13vE+dGHpXypEkROj7uOzRilMRVQ6YRbpqr5RiL1cddhqjj+hk2Aw5UVJOr6BAl6nrGz
yZloni67RDiv3/GGS4iZpPqL9jxWS3pi/SkvHuO6DoX7Gc/cL9EEnM0XtJ3wOpkqBVrqpbhhL4yK
5RVaFQD7hT50p1SjMLfN7ZTzXnBjlLxd1dTxHHtzecCnwWPY1mnYguQg1mjqFgaoNz7jziYZYWPe
1sSx4jz0MsxIUxa8r+sJthTKJmWI8dEPhsjDxgFeFAlpcxRI+qyJcIort/qM/VzqHkvktRTjEJFx
OaPQ4INLEiocPwVW1xkLfTIinUHMbouiddC92LF57W8IOBOMf+D103rPzvJIJBKgeMLAy51KQeSI
uy9WcAym267wqt8GtREBrgcve6Kq2k3dYbjZRh9HEJgfqEi9z+1IrA9jGyrnhNfxLtDcjfBaFP7r
nWX96bAxjUnug9KGF+X2czP8khTeQ0d/Ga83CAysiH50MlRV+pYVRoelgBGJkQV/ftClMtuNH6/Z
GGp0b0hARym3eLnrz3aeSFrCQkF90o3kX2ngC5RLpPfH7aSxRw5tluNRpUxisFxQ8unwAuTUTQPH
oXrhDlccFtHpmirnTF9xZ9snnWD0jyD8Tdjq0h9RZzakTz3Ybr52GKrMlzJKIp2GIf3TwY8w+6p5
EgWYzPZbbC+BjsXv2bO+PEpPBgks8PvwrJjsiAlGPMHcVTv3m2iS9NuY8oTwOzllOAti5WgfguY9
pL1XU5iMZgRFdD0FVkp0Tt+yQTc0BAmjwxSol0q4JbwK3kpN2dbFHAB3c8ZqVz8Myaae7debGwXB
MpPibFGVEiC58HenxkE9u04ra3iakHNO3VHRSuxDjQRaETVXcq0ALjE6D9ihiJ/ieldUSsZeJrXW
ZeJ1HZFvNKRW58l4VzdKe6/jbX0eIzl/9IkBxHV0+r0TMyNqDFn3Vk58KAUmfZxVe5RmZE9RUEr/
PIKr5HL/b0PWpR1NlUXTl2oZzKQPAjEkJo/+A2ZGnMwm6QqyEQIKl12D6szV7C1++mu9u/PdBbke
ZFAAF2ZzkSXWTC6k4ATnOI0uLN2wyTbCHrcKOQCM+eP4v0rGqpdYpXkvteUsyYSpOUwWandQbuCA
G/oE5mMgCC6Fy/73SFOVh/8jvH3bWewLcPsB1pT3hC/lUPzFsrRaBx9W27n6c2hqlEBOgQZq+cbN
nliffVT6eXhzmlvPhTGO/OKEkCBotVS5HD2Jh1sGl0dCSW/GQeBN7djCNqL2qNKF+QXzhHmar2ox
/R0pYM3lPcYbfkPFM9UgYmxNTU3n3iObg1vcbcsth8v2Wz2VNL5NTZywmiUoTWxL7O92AfOPcUec
lb+ggMD191P10DDX08Ci/aeRnj2B+b8DCeU8tMoloIW8BnE3Mj6O4m4f6r4JzWND0h8bZbhZI1sl
mrlYGBbjWjhu8HrR8zzuY46QJ8tX4UuGS1hHFUh5CtqT69/o1Gf2bUp9zKCQ/9U3KA0AMuy/iesF
n8qO9eQDuTS1/Qqs70xGbJ112m4+ny7NIlnfBGaB66DpyGAnRNvosYlqcHDbJ65cOo6W3tePPCYR
yOY5+PayA9hCEH4mM/oFsbo5lIU+jX3+7+lg+PAD3R3XHolTeiAtqlsugH1yxhNqlnPP31NnarUc
kWGOpW8fQIe1Hczy/pOn5cBq9rS8oFlVLAgK7Y4NM66FCeAegfgvO/CkcUeZsX4KrIvIkoEKW5yX
GrcTIT0iBCZcxwUtMJKfBjfkPOzYUWP9anrP672Nm1PYMlkE67WZpW+ye1+31Qn4hTrMNwk7DUdP
xqKLpDTwTshKg6Rh5BcMEoCz4OBpBmW0buTGJ3alHcaJMa5ZTgHbqjadY/wN2BZTDfdnz2SJnIcA
mwgvzC+2uS7fb0LTcLqVC+TDdITMEZ6ik6P1BobiiQv+up1xWX2FC1+HOP1c7nbWHsGMJovwZukK
lAmkLOuclfWbPCl41b7qKgnH7PR1iaBUPwDeBvat6wmbqySIhSxDwaLrK65XaC9xbe1lMcwmJoWN
awj7s+UK01Q2n0QduCAlcUJ4cs7Xtdlh40jkgGAywdmj935+ZHkUF03KKyCP8yzHnv3ziYvUUivJ
9AOtFb2wINzzW1owbhvJCY0IKHRPZy9jMAMUJQ7QeH3qQB4CflyqZFsi7ypTdNxC1VtQUiJMJzJw
dpRw8/IHJuMdW1qqjc8UYS0cXNnwwmjZPaPvcCKASGerlUUDkjV8skbsP1dXSvTwR07YCbHYwbaC
SGmhLBIEVDUbwx1yyKtcCXT/QeJztmK+2tZP71/REq9SnNnwvK/pAV8x7stRTJBXmruFXooidwbz
zFgstOy66tW7kGCLAaTPnZBkjKxZw6NDdQIUnUT2eCDx7FCBE8w32I7S09ZUhcXTeJ93gfJ1l3oU
nAmwK5xjOHMK/Zeov1tMhi3P+BXck94MG7686JKO8mjs4kmyf4uD+9WD0EYDKJFr9tZvXLW+lrbD
pwDsobqouEsIPZggk+nhnJk3vcpQirfd3Y0XCSUA2ZacFI/w9TtJq0q+0oWwYqWyenerv/3Ndnk6
zu25R7P9eaw5Te/Q+y+lwgFdHNX3WLNpMvCOBC37x724uWX3OWzAJCFnEmnJ917cGicSFYVAJ1Bo
wWdF1ZVY5tDTW40gCLOgPm35rb3iKSL9dEzBSBz1Q8Q/k5DZpE35/KUGDZF7bAIDYmT3SPAuAB1W
O6h7wg1IvAdEVj5uxXPcr19PPZMlrJky++mXCdqJnyUzwgsoloXWNo/NNVtw9eHmGvWOZoP5rhSe
58ujDdcBZKJ1f9c7BlU8q3ZYRw66Qss+aLDFM/ZBmHqw7G/2X/L6VQ2Rl46rHASOe+XOzG5HqHTG
auI2Pyih3yUMFR/IkXXQcbQXtXzFXDcmtWUWrtVdtEVSyNb89NJntt4enLX+Uh1bSWIRqI0y2PQs
Irjck7LislJxAbSpn19eroSMtm9qFYlo9kpX+leb3S4vzlblqUea+IdUlR9qjjSnRnZt51ZuLDlQ
zBx3WnrI9KbwaEjl8S368YXKVLuI0yBOmdN6AmH9hrhapR/i9i4xGYTfWSLEwh3iTi/yKGa1z+zq
PW3dmgCAIwz2ig7fjezXIt7w+6gAXM95haxSKn31Au8DFvgqaokN23VpZTEpXnoL+2M78nTAjzYb
lueohG7LNWpMWhr95/KahLYUNs7f8KFdS0oSzGuzuN6JjiRAcv5DAuKHdkKHIPTzIK2W9gwJF2hd
8OM8Jz+wp+K2r3hnSTpJQjcJnAoTkHHWbxOSqtk1CR27JPM9Ar0IfMVx8XrmyzvMrpISVGiZ8WDc
9yulDY1cdsimKUMA+CB8xa8v+BL8fU+iwsnn3TrBwGqMsdrTXQBM5vFF2iOjqDKOwMdtHWl9Mcq+
bP7hjofMCH7AfLnHpUNhTNm/ERyTybCYulK1WECnD2By/Rw2CPstFDyXqiWgGp9H5aat6aT+QJsb
MQode3S6wZ7pd4aAMyM686xZsGwbvq7HizFUJuiXdpABlvcRwv7zAAvN0P9cmR9lrq0dKOYmvJlO
4SLMk7+DbAX9diFvNWFEMxrTB6V8NBEFOi4ySphBLj/wFfKdpgnON/tuJdIkV0/RpauPiLf1fE0c
zgDGR0VHE1j4atkYDDocfmRLS6HD+nUDCj28sUS+7vhhC2MgJH3GkqPe5S3T5KDNTkaD+ohba6sA
oaEGu2144xSwqy7I9usoeN4343I8sGHKoPpDcOkgORjygc96xINUYb5pRDL2m79oqPS3vzHoRFes
ZyEBwZdsLTEPhKkEW70RMG5I8RtkKWIis++TU2TIQHRZsZwI6aU1yPFwfWYFFzUGrT0SwHnB5Twg
1RQgd7di6RMfES5Rn8dFsCHVDw0BJRdVft2NT9qewg3Rd8HA9OymmB04U9CUAIF1ISh9X994kt9T
OuUnoUldHROo1X8NY9TtrqdXsFd6FOL/8TzQtp3TCQ3q2MMGH+wFJhUpSJDVRuLohgbOcwY1+zjP
IaAVOb3yYEZtTvUw8m+nonIqwZirLHp+KW9BKzy4E3KYFnhCm7g/IB0PLjuSI4isBn9mZrX0E+MT
PLs1jWUuFzghdXIcTlX+D4xequEdLKRP7sHCY1eWIjLqp/5ghhee1z6cISkPVbdFalSMnnnZ35oS
e+mScddDpf929JakVaG8v4ElBoaBeZqg92ARE76iOK7pkFdXP7APXSNFHh0I1zA7OaAcKGWtUYy9
5APdGJA09/HTY+2dru2MmXOrzo5UJMI050qyRJ3sNlH0lOREruehFk7gJupBf/RXDLbxeAftt6cP
qOzjXs6seJKGo/lij5KPv0gwUln8eALGmcPhLzO4YI+AXyrDiZiPVwkZc/NssAYpGO7Vk3COxV1F
qf5ZriYIuayljEEAXhjZbRQ5RQ89PxSbLqhtN4NUGlzJsTsTladSvPJnqZje6dscxsUmFMpAbxLj
ciMMxTbsPPUvVJc16AAARLVSZ+KzdqWZWmqf71Q9lekMjxc+YNGdz3PYOi2vnZEkVo96sOQYyz0N
qS8QYuNbbMWnGVSfpKL+xvqGLo0MpvgfG+Z5V06EzHeN05+UvXCu5Q6hRMuihGd9qaOWKMngAIxt
gIpf2MlOZ7xavA3V3ZYLu40H8/CJBUb9oDCRBysdsIFfyydXjnUiMYza4ozIaFTWWZrSN1h8lha1
raWDjSUlxlhsGa2xcSvdWTr8A7SLM80z55XcLmIydVbKFj5nJEmJ22SU4kNUgDqtoOurIC7e2RQL
zkr4U0SaZhansC+GqZWL5oZYuxeryub98DrJuYV6upR4CQ/OqNsqhLSQaexf4wgE1GSI36bnpFn0
vg/Xxm/mPgrVE4zSHJ/kvdySBJP0WABk6kFDEOJEWMg9QSUU1e4kAqNbw40ZEVxvLY4Gx8yhn/0B
DDtPNAqShv04OsLABP4+eA5+8yanUszJdhtdKdcy2bl+S3Dm27/nQEOE4upBq2GKeKBYiMQZRfYa
T/V8vFxTVgQqdPAl3zJU4NLCGqimuVcpXci9YQ4RPpad1+cgptooMKUWSIWbh9GeKkYEMJdCQKtl
KgjuNhleHD/gGXiKhc+YidapDGBmmEJDU80CtF8BUQa118/Ogw5xZUDLLAuVsJ2SCk9KECffpP5v
1qKdRFg3uW1U4CjgeAvMKu/mvwl0ixb7DfUBikrA9nesmpQ0ctYpxQuOUYGohhVASi775NwsDnJw
bLpbOl7BrPceXex5RJdXtik1tDLm7HgL8/1cNxipMr7rHZhS1fG1UDAyAwn5Fic5KlcWi2JVR/34
abZa63EJJv2WPahkHsEbfawnBEqJVQbINY5ubLzNt0rE4UdyhdyNthv01cDRKESvaf2E8eU1k0wi
0C37BJtYqhoOsNxVJv3z+8cwGQdJb/ymLRH48U5lwC25Eyrpi2qKQqpFS19Uy+dz7sOBUTLXjhji
Xss05/qFTUgzwM70+9Ciz84zs8Mn991KPXNJlhmX9NNZ+7akK9zt9y/4Hv+09We90HUudgKnU3Jv
5onLCHt4svsJhPAzwfVC51I8L0Xdeegkk2kZxzN5cWHXHCnuT38TcpVh0+Fz4TNMbE/lRXtGSKoB
ul1PiR/VAF4ydDYSZU7vD1E7fg0xus+an2nizo7VcdYF0trulZaQzAZtVq8LPfvF8Sb54x69Rnby
ZZdLO0HzWL2o/C3CHRNtjSvxq7TxRlgZBUhrq7TI6Kz23HALGSJAXSJNUCh1x+XOabKhCbFvXlGR
hySzuZwtnynz+6OxUs59eEubnZ1if+ZbD8CA9oot65NvuUlH9y4yFHyGn2PZV+zY6OFU+Dj6Vxa2
HBVWI4IuGu7LFVPHX8vunfa9FVFlyShACYVCRosAX5yxEFmqczzfbUT831AFEhGZp8nVd+GFI17O
QSvUzTiatcpAHlBLtU2qlKcOFSlFgAQEOLwhtgu7ga8scs4+w6ZbYImRzrh6aqtpzdpTY/u+VZyw
fjGP6KiKyI3W2C5En2BH4Qpm8IH2aJhetjnehueTcEpBtDLH3g5WFMfF1SsrN18s00SUOzVzsAjm
7PNk8kyEWCP52ypw7RFtKVAkxOaYEDRUHeFMnQd9/+UpnPCT3JiCTgXWXfkfMDX8xPUMivyVuh/L
u+IW1qWx7Dz4qJAkUPaVFQzEqSN8xH8BrAp6ZvDgpn4NoYwLjAHnQ226648D4Gb2b8M19XZ9LEh/
KMOYrGavy95uTNOLjAGW7HPkNEQYVLhcH9OlXsA+TzDHV05IIE15LprPLjntehJ41VrbQhk1z7zD
GyI195HIdcJDiOLQt/fwI9O5eZuxJZFB4D6GZIxi1V1H6C193ZPHZKca3zdGEAltEfdUSMEe9GXZ
xJuFAprQutJ4IZVpXXtwFu86iOtV25bxjDBNUEdH4LzZVChx/YeY8p+4Uukn07MlB1VazLItjq70
R7ul0D1BRUG+8XXPDKC5QiEHbbIpgGQbJw9w76GBle1Rh9SUkt/mMUuf8f3qYGUaQhV6xwws5pZf
PEA5vR0WhGOXw9hWgx9le8kYbXCDUkGEI25og5TTYHgxMBtR8VoZBwIBFM7VN5oFJBGLO4nR1upI
n6nJBZuUR7168kePa02g6+S3iAlFnkjxHEb0mPW66v8joNEY8YXvzWV/RFT49ak9FWx2zZLjnrgE
i7biMqqG2VG9HFCLD6qH+XtOFCsbzMd6LwkAI9/tZijckkW93pJ2ARFifS03hmPVSETByB1D+qJG
b+PhyoZi8n8Sfd1V5bKMPkILcF4lQtFazjNY1bqlGNFGG4SlseWm9jeBKjrvZA0RdkaM9NEs1Ygr
EIGKrN5MKqZLSAHoLy1uNaNaGrxfkKUB3UKdhMsJv7T+cG+qpv6qMQj4ak5+uisYTqD/2a6cK8wM
PGLZBzUqO50teeukKm6UGs88kPGuMDjvmErr9FNg+H0L4RO+kkZG7HXDv4HB+FLOYx7WTLanR0Yv
adPKeEIvOHUMycl6KpgFJjCucA/eROmDsksnx2pOokQkA0uvCkUlPnvSDtMCSN1nDIUC/7rIc5QI
J1cid5jEx/Xs/ZHtC75kuwckaAHayoZ15rN6+kVpJkt7in8bCOWiC5BprLd1jjNMVNle/a46c8VN
ideeywJfOOLWA9Kgmvc3MWbu8kzV1P10JLiwRoYhmzJHmndsiu4ipg14+sWZY4q79X22B8Prc0dO
5E5aXaVlVruFWeOGmfSQxYxK2W/3NPaz5Fkn0USwoKeA98sW/jmp7llqfYKwvwMBLMxKf5MMElhH
L/td+3/d7h2QLzpZxjoy41UUdonANEWC5wbvmJDDHVl55mJtVtO+5ShewVjw1LXXB2O3sGerzUbX
HYk9UIAdamXPUFzv4/q5MJdxsx1z8wzRqY82wYF0YP+tvFSYxmCQV7SW989nupK/4S1y/t+K7vz2
cKKrHFgK8/pUrcHkWiUOmtrqz4WOyNt1TouJfXURwLqHxFruk+iwyigylbk5ngQx5ThuAkwlKuZP
tSr569NTwknZrE4Uo7RT9p7wc4sh12azPRrM6F6QlZxG2cDhtabrNMJTaXMkY5d64e9+VnBQBjtT
QVB/n5UYK+/5BD5KrujBtSlrxVxBarMfss++jeTUVmHSehRPVHr5UyQtuSKBwIH1RS7G6CLsL3ns
BYuxnbOIGK6A7mAP0jMnnKeWNNFxKq4+7qBwHhad64WNjdzzt8wW6+/2VWqIackkvDEG/0rAATtx
lvJGekVQgtjAF2VWK1KxLxEr4z2hUfpvVR6CEBl+5sIUI57UTcLUBC6f46NZXc1y4VPEcnrP367+
bxstbOSHw4tgRTfNBbwZRvnBV/2ujoW2WMNCHsUhWKkkIR8PCJR8GYWMop21K5+lWO9s5Ni8Paos
uwVXSvbyzrA+7cgzEXIzoicNJ11kyUVl8lqbh67euVTiRnJcI8JrKu6dHvVQuyA8Vw2uySQQLo+z
jUmMigAee2nq+bsNuWIp1Jt+EtWBU0Lw+ztXBe415d8YhygpFB0ZCF95/3r8V1yY5s94WcTxMjZb
Au75gUUWUeXg+d6co24JS5QAnC53bvKvoV0tI4upqKmpiIfy75I+iHmnW+MVmm1mtSo8h1ELXNHY
EP7MrqJGap4zOEozzH6TKxYP2PPsJm/owTdGKKkUkpdfppAaVEs9v0zGTp1PVCIN1HnSLzQQNT8r
YEe9Do+eAjNFKwrv8a19wezjUCeRPqecsERJLsrmqJye7LRPTNoX04sPBYkHSfa+d0mCM6yoB4mQ
ZvVcPuQ0ZuadVGoS/9jktsGIwGTG4v0QWuwe3Fzt1BW3sr9nfdf2jHyC+h1GcJaaLLDaLEUnF8gE
MhBn8wJDPZSSgYw8+ja4FDfGQGMHuKYvVYQfkoISepKEbR60k9Arww33b6DS7sOL0H5I7Ww6A927
wcn3hR2AS0FnNJWT3kQzgO+7y7+0KGnXFIz08q/2plSk1O0halCKkqbYDLysu730bIxrkCa2PSUb
nBvDBYpxkMR1u7nuwCndtWWz0MwyJBvAjAM9ghnQobA0TsYwPIAj6xOhTyV2+VxsuCxBT7dPtzBf
avE3tHZjFVVvDpfFUmyDVYnJYvXCIL9sm+XPxKn3Kv/hLH14VS5u5sCRfcxJz/86ri1AqIZlLRn5
nQN2J+U+RrS4D8DX85SuNWagY2DUhO4k11pkkYcM/jRjBfDWj9Hx8y1h3bxtLylaL5DghqEo/mBZ
TriWq50o94COilzd7iFU9UbviKG9qg0N9q4BOq4HenmZZum8TGHzcQA9BSO0NcaGghTFo8FnjPnj
BIfq7Lvz8z/LeH7PVhhjALbi1ApWmYJsoV9LZutoMGqDTGacbLicZAgE1A7q6GLaeHarUnXeHUeJ
c1QoqOgd+Ivy5q82bmd/gOBqrTWfp/f4e3m3sW5ARt1UIuxdL0BIRVW0ehQmV4rkLcvayYsBO99B
SHfRvKmPt3xWqiST3Ld/x2EyfkAqxDdTwjMjB2J7Gonf0HjBkGX3MPPvSvUH6P8s/Kj2+DI4JmGO
vVcfkh+GBCIasuK3GV543my1/4QJlO583MWtNKGRKECRZB2UuxzUhQcqHzbwBpnevPyR1PBVes7S
YtgBFvESAZptguV4GJjHZQhpBA0fRyx1bTA0ww/c86PrhaEDP50rtG+aRm7ImHStKd6VOqDB/WM1
8gvRPU1WnyZj4yrFoVhNsmjmFOsFArfARfDLm1CYCD0UYEULE501p9PQW4qSwOC8WfeB6ngCi+Vk
tri13mCDEJmLh18PlSmUUJGpkFs2fLViuSXDcGlLxFTy+QNTxCDAkhEpof/I4aR1fUhwYrtvCNmn
X1cYrQTOg2q19abaqw12uHKSiRrkf+D7G2gGe1G/3FnZRlXEogFS3CgRAEJKH5eKnWPwlpD/z8l9
svotg0zCQAcKU+pw322AOY1vfr2vfXNkMKoel4EpxZ4WFHj+VMGY8lz9hJaEyKa2C0VCJeG2v7G7
rIF7aTyr8i0MJOwFORJ7GpP6SHUyYxJfAOFMG1C4nCwmHd/K2wtrIfcmpY2A4cQtfIVgNzLWo/o1
CttDYjJ7ISaRFR3ZyCBnA1YZhesJVegD73s0yfrg8w+ve27j0VzhM2fdGBtORN6N0/DJDewyQLDM
LR266PbLL/xkhqwrif6ACdd2hZ3AJKg01Bmke9jwtQO1kroOaF6mOtpYyGUdV0d+vDI6YZq5p5qv
4DR3EFm86ahnpz4a6IHcsLPWw2r3jhrWfSybTqPUWJPm26rF6vwX2sj579D8G1gtNsvtYqVRGqv1
DDTLE3oRYuCuqov55lsGEE+kOlrxdCdQcYLvETGMs9VtcQUe4KgKBRyoGHMEjfXFXpUgcG8naTGA
4v8JpguZp4d5EBNpRbrfOOZ3MLEfmBID9kRzFps8Z4FGbnOC2eGoYKrJA0aU26MEUd5/naX5SYxW
Npx0w/zZklEJnJzCMviLHgAM4Fa2EYyG0uTYnthijY5ufPnoGaRhrE7JYuMXnykO7m/hx/Z3eOhr
td+rv0OEonw10UqB4MLj0gu1w9IzEhN17FCCmQsu91stunjpiM+Yf6Ct5Czt8Duyryj8rTZ14x2e
qooCs1AdXsLFCNfVv10Kfx1psIqgX+q5DtZmkK5wZ50cgkU5H0HkUyvVvSdOWEMvlbBQZfUUp8eV
yqk4DbM0CGRJcPL7atW54egzPi4MEiDL3LKeLPxOMXjMcA/eAMHYVtEmyWZCQALJN2FddajmU7n4
9ZfafOkQ9UApzoCyaaIcSX+TWluzrG5gCKs4ZgvEJeW8Uj+48D5JyGEl3DCs9WlleeYzuzOAGFp4
KNbT+LX1h4QaNpLHOwgnw879YtxUZMIniO1ywfzYyEJ6nhM/1LGUcAXZyLSWEnudZSB76xGn74ym
QhDVrQXyGsRJYOuGgDJK81ADSgXbwWO1ASiV5thEAFGiqqb40Ar0o+IRkcYIPVTYKUPpRadJXyzz
UZwQ5NBgb+fuzQrBi9HU9JZXtiGMCENyt4+2hQ72CWvkJEbNc+DjQoQWcFp7/HfxlQywQalOQw32
ShYzGdqwa/fkYohkZlVX/8Olu314akR/TKE1anytC5F9B+DF0vc60xhs9bAtxAOXCBMc8IAQTM0O
9NEfHcpjVVPkevqh+RbtAhK6BEj168DMod/Sa2QsxPlu9AIYvn0ieatKGVyxLSySovg83XS7rZW/
YJ4WrVbmp1hJ0fNJS5lY5POnLNgztujCBaDpky/5yEukoxj6AvvUqrtC15Dx/0OGIC9MzNNQieIL
O8atVc4HNnfg7qjcDx8Bi/tafaep/Dc1gwXXNeRcjaIvHNUucNPvQ2UEQhON0WCU6vMlZ8XDPmHq
8/kzCOqkGcRUSrCXtCInY6r20luoR+z/kvqM2Obxyr9hdnrJIwIW3AMfAIJxYdc1uTidSec/+BRC
/DRUxC4mu+DIE8ltrL+VYWMYAYFyCnd2V5h+HH/XNnH0ew8Z41n9gkAY4zHj6ty9f83IyzV3KrAi
kXVbh/9QJh912WgsrNt5zyTCcZaNvaUmu3b84HXzqmlV+xjFMLp2jwo9DNElcaK060n/lSewbJDU
IqTYk40WFZQVZO1fNnPYPdBJB9MirAJc2VMqwUOh9uw9PNGCtLHovDgcd9p24FBFEXQB9Thzh2Nn
iKVm56hPU/VXgtAuhx4CE/0DRx36p0jxGnMNi4OAghTVzUZt0aDekqvbasL1rMsf/Gw1BX5QtR5Z
OZTi/3+5ra8QUMw4/SdqK0DMo2yefJTAtXqPR7ywtBxS4CAjUyr6oWZhFQVaa1KRVuT7Wo4guK9B
oksY9k7HJprl6Vwme6t9FmdmJXOtNCkViRLeHk0AebpGuOlSnJqlj24mQ222QkIeaaue165zhdYY
gEBoVE4Wyb5Me/rBvlQDt2qZJV1vmfrfZ/dhqlKT/wQxFI8rqRhTr8/+2N4YiIPqJpBzEJ0w4Xw/
OraJ8ayC28iQPSUlYbM+HZIVsJQKr0hI8RehVQ39QTl1IELoxi3K0n8kYZXEp/mER6rne+kWnJtQ
ZE1+zM3BsZ+qgWqV9uoqAUr2s7rzqYe+FnE6DfLEasVJcdvHgy5HHp250Wuj+4vqHPYN8KIlZNha
oFrM3Jm7jWScS5+HMETmAljhSZ+VsaBg6dI+MwQd9fJyjhjRNMVuuCauAmHbQ89ZWP8QurLtBkJ5
n6gqheXOY5/52mIxKlhOUcCSG0WILXWymKiUViRp/AJfPlh95fQ7fsiQco+084SGa6WAaA4dyu7I
PIrnPsn6r79snKK5qz2pa+IW5pHK2JNNn+kX4ww87/euZTpKEAXQMYOkMTa7ey6InsIq+4YDZwiv
WKaXFcqg+sBErAXB7UeLYwHtZeBwQjjQJ75x2y1+zb5SxNaVXao+SaguUiQGYTGS8k6aX0gU1gYX
r5ohXU6U9sc+L3w4kQmOkdt5azKNgkr72La+GKXPE+WyjRaio1ZHCvicKt8JyBvpx+qxRHhqGRZ4
HoWD0BueD6lMoqAM4XEGWKqCAFXhfHLwCJSvbDwpo2fdfWFGUdl7WOmjcQK/Qzp7tpGB32hwrVLT
J5YcrZw52j+7S3bNR3xlEQReeRiPz8Tafwo59t40W9hQu3WztBrhc4DMWY/qBTEKU80oVD8C50w2
PWAUduyR8+o2mQhAPkTGOsu0LYv5q4n1OCKHd3YYspR/z1knz8Y8/mMqSFe62adys1Xe+IgQjAAh
LqhaS38mdb5dBZ6g5DVO1y5tnOPr8w6FKg3BcDaM4r3vA0JfJg3JWEH9wyjbMp/e7WdmVLYlHl0N
VKXJEuo9kvDPG/ADsXCztZamhgjxY3N8apZDyGVBmL05EZgSkRSq8sZvGM3z4z33O7Z3jv0iYvRo
P541zACYTv2FSCETnrWbxoKkXkuM2LNonbpSc+hOp/zTNFWL97yU0FkaZSWXHImLgWwnbnxPRMEf
lHBN0ERe5TsWItex/HLiLPGPnayIzwz0Q3ojxBoM6jARxib8C9JV3aePl3HquHKJ7VED13hdnkYc
tLGGt/yK0gxJ9+KH0JQGyC6Ca/H1pdcA+xHMuxz+p9HgEkdR7Rx/muWn08/0osiOtz5Wu2sayW+y
zSS3Pp6uBaCP7Y0VdiWxCY738vS+yU6d4mG0kTbQSzpxVKlDq4XB8UhopW+SJPVgiwcD0R0c2QBT
z/7KHL06DgItsLJPXykYWI8ZXA2nNpifdhS3rbF7wSf0WAzfr6xGQnukxVbVWRvRqzYXxdgOHP0j
sZDVydOkqVKJOhxuzYpvI01yQJVEiA2BkAsIoDjzlbsph+V+diGIv8om0o5PfM4Jx4r+SdkntGSZ
RO73YarhwMR5ginmcFVbuX6T+a00SVWBcbJSWC/fIzSEewpvGztdLtY3djaERMUp+YRbXGv+8UCx
r0xrja9inL3ObXPBMu21nIpREkZ6YrxE9tWK5s8PWpGJiMUGtt1yDEaw81P1F74x9rzqmsHpjD07
2XXPqNxqCF82e9UEGXD/tAF0PpyRIS+xeACq0teC9r4Xzpj545fPz/smk9HUshYk/lwCqN8rSmZ+
JCplsHxUlqQ1rwkvOalHuVLmUxpkAmz/XjuomVXIvyHMLZA/epWNvXIRJJeI1sfapwls+kkrdaiV
Lx92iwfrsWgv33FM6z35F/iZ0GLn+527SwiTGh7henmTX4byY3lHzVlf2tVRVQZZA4xCgr21x7E+
cVLi3/dB7nZeiessOFvpbYvFdl1BGm52K+rq6yQQIb15ADDVppu5L2axQhki/ME0VF0Bfw50BAL8
SvJU1S+s+JJ22e6i5dCdDyenk1MkEp5Q2/qGpte0/eU8c7SR4lDFG1bZWpYlwagvW49JtHrfsQgr
XJsVZ7+MwPFIqJPTAQes7Ru2RDw+vg4nq4qrvstCZPYbAJHoIlxx1ZPlQlRYWXqBk5DDp9nPZprE
6iAb2orLkFyuQOds41wxCNL63iaLFbGdKGQRak2YMDAYQfhkYSGM5Guxk4+YvAKuAn8xXpaQ7/ym
CPTmx7tXXtVZriiR/mqWRh9gquQomqmK3CzNaQhKM/hq4qkt8NNJlGeCgmncPhuuV59vQYa4XPUq
13QTxg5xgKnJ/fC+iFWZLVpV1G3/THb0UIxXmB2cxbFK8W9DVMEp9zPFhDOvtS2Gt/9n7+cKyPsN
TthQ/IdLo0feA9al/6N6Y+anpsuCSwYIxVLm4+9gjgFdYZ37OtKAjY+hG5HsuP9fwc9fhuKe0bQL
3OAJJ3WER9qD+S9po4mKSE1qba2VektjNoqrlqWjH7Uim+fW1N2j+1x0BXOtU2oQTo4Qsc3xwOFk
dN6bzXAVm9WCMX+LPYvyVPWi7bi5ZZHV4Ho6S8x2grcUm0Iu9WzL2jPpz3gibaLuzdHa0hGuibDw
hHDxSvCDEWDNqHTlkXrR92ne7YMj7ZnzQLeBWjHtB1dRn5Yp4M1+WfGNaVKCJb78uXTBqqCV2te7
B3HkgQg3xaMMpBlBFRULRkmj1tqmeRUF5fPZMSsaBxB3Cf2VRzeoDuPSU/NTC1noGYaaGGa+95Gv
K/3GxeRe1ZYFCV6WyoMp2v7MXwa/a+iCWthY40qIWWtWSbFZhHfH7dkJQyjBoLxmUYZfgKZtNn7J
WbVcIyJcLCIg+VI7CEsLJh3/6QbDNh/HqnyyeZ8LFZh5je2TY/fwS67Jg0HhG5R4hKuOUhz41Vai
tDypzIf9oAbz9dm8guJAI8MLSUq0to11dFZjEDIwwiHrbV/VQKYDqp7Lp55gVNDG/Z8dSAMIwRl0
Eo/IyhAK3kKznLkjEFSoR2sROMzpCW9HyXUd7WWTKi7iK1AJAAdvu34CGpKxDUUoBvCaK4pBGeXA
DNeIlcJi8TD8cBoM3xLgTOw6V2/OUGyVPzYEWwdW5Z7D5bXWnCmg+bLy8WGYaX7qTeSw73ldDx+u
Sr7SjaoBB0nWWw8lM15/nx/AgP16wJpCg0GBRjlYovs4ngW4r/WMsr3Qd7wk1SXXzN/nr7t/TxIs
Tuogpcn8lBl2CZxbYtzIZSRNFBp1pKBST6PqzABSP6aZv2Eo9eKozMs11bvHjgkCt6OV5bNCrUgn
vIxOqphwTuTrXpYAG13p0K12Aao84/EicF78U0mPFLaj+lQh3GgwGUZdyEZARX8nIAwh5Dp5U0sK
/RCWfSgCvs5Vc1xwK5XoP+to7CrjGYDCFFwbczV1qMUxszK+gjmjo1YpHIqQlrbsU6PvFmudCHrK
h85wvRjjBULbiV1o63ahui+hc2Q2YolwePPEiW+RVAFXWVPtln0zv5CMXSXvjbAgcgEmeum5OyzP
KyM8IItvmZQ0X/ZK97k9tErg8IjEQOvZ6mGNsoaVICSNqdtjCVwclM36HvEum8es/u+hfle2lxtw
Ch6tJE7wf4suqeR0EjFKuHTUTOJ7kg7UAwWgCpSgvYZUNT0pQoWoyqPEy0IEdA/wBLWFYcoDz90a
CodMQRRDzRz3V2/XpkHdBnrAYaL7YM8GN6CY16/4/lTx95cgazKlmltQHYAfJIeC5Vama+osxFfT
rnKoiPYr17X54Is/mpr03d5y6oJYO61ky22i3zLzWAeKNdBnTWzHoEFKFR2dcXiZ9svnLcW8LNmj
QIYmKrLE1MhzIKipJyfCu+D1pQW+EOvZ6oVaSLa2ckiBglpCvTq5LnpBDmJdWYAV8lxN82j9w/H2
N0jWOoWZRdNpOnlAskC9oEHx3lpLhmx7w0A0uFyQ3SLdOPwEctQhuralYVVi9xaGCwXDAEjjgTm0
pydzifKL9Jrv+wirzakKekaS0gX2aroNqcoZWKRvATGRPtCdKaJ5HXnbdEFwXOIFtypAf+Ynwedg
7w0u4kxN7YMNz3zlqsiMPg73dottt91NiAMMAehdNb3s4zXTeTkA0zOAIpIkaqsvHNKkAAhdJGC/
srkT5NY6vSZb8mYx12hdmXQ+szGbebKeevgd8xvjvzZC1cvFiZ+I2ZphT+hINhFJxOpVXKczSe2d
zEHhpy2ZORx6PVjrimopqT5wt0thiRxEvIS0uDsnw3pTd+u6SUPUIrquOwm7uYwfdSo5vLAmJva1
ZsAi4HKYVlTMZAuqq/wQaUoLhIEXGovE7YBJVuE2uYaX6oFpuYnBuVCuwiWLN5UWN4T3GquBlb26
fnIwkTQhRWoqPClBFyT65reP/emiyw9gqp4hTXXbQc2uF8ve37KFuxm+ePHtUm3bLjcrDMhAxQE9
jynHOT/Q0C3gRdEGOz4ZzMJyo51TaBpo0bTS3F3zwta7kWUEF0j4hopMjkgOvS9SHMe5Vm9RVDw/
zq+f/A8U/Wmt76S/R3rtA4O9GfNDIY/p9pPMM3+4tiF3dlXXlfEIhC3hao/Uq+IE0C5ke1xcsos1
i1NO1255Slh3FZSSo4E1wgPwm2ggJ4f/SjF0Usrc3T5/bSezKMqV5rVIDAiolAZhiFA+VbfRRqWf
wmZmMGlSYQ6ORGQ8TULMGOHcRx3pme056hesPo2HKs7jXYgX35CIGGrkteJEUzJRmEeLLBK7tw4X
Vdora57/YzVlUe3d+hybvrB8TGNSJ9dSE5SOFlEQv8BqWViit5Wj+veTHAiyGXwUsTFOU4KnGK+I
P6dED6CxvJhfAt5Qcy0XlBdHeERL1NaTrvVRjrKtUeyIM7MgY0HQGhzmZRrfsVsRnnCctX+mgH4W
69b04w+hKlBioahz5RCy+R6gkdUruQb2vWyb5DFUEY+nanBYmIdInL1AFUQ+EcBquNhGxQCQFyhE
lqD6vSG7YOqh4YE3M5tMv8LnJR7+foiG44FXZrx0eq2ISzn0SkAjJoFCkl8XRUJhyjx96rE9w0Zb
TbCcnw3PKOCKFBBQDgiNXj+5qnmDi7w85oYy1w6JD9QU+FSkVUbnJdGnVjV2EYKX3tzp4qpgVrM3
WeOL4q92PcIrS5SRRSIDEhRdleup6bk2Fn+LqMo6tSXn5AoGjxwfdkG7hRQSuL8iSE0QhhBbn59r
WyaXO7kCeFOsdkeFgaHlg2OcKHJj6uTaLfmBQ2M5IZEpKf3dIKQ3gTNnthmOCDk+qPP5if7foxdD
xSJ6NjjBzNodsCON7qcjlHWj9GRjOb92LoCV5V1zGCFizrDQYJZFrquuJuT0tsRebpPQA6W4dM8N
dpvlskD6E5uWKpUmjSyY68BGzzaCYdXw3lcOMIlCOrgpwtVKAIvA2IFPp0S5m8D+kad/4hDGWpRl
qDSJeQnoOeQONUEu20D8OIycXEogDcqLnMXvZzavJVVRelk0l4qBWB1TDBl3lX20sDFYQw9Zl0FZ
/akBZH8Kz2usEjPkgfVrg6V29bRlBdq4ZL5KKR1COPlCXIyzg6pt1BU7rRtrivupE2/kwIgg+RIf
DhOZ8y+Iyr8N+y/51JGFOt6qiyZvGZSbZikoEuPekiLPQ+Sxk3emNfMnyacW1GYDQpRj9ZrvlZcl
VkgNOB9Os8oJ6eFkmgHMw88INM7IzULP1+LqCIz2+n62Z4rdamSdT1t3wgHOdH/dNWPeWXNTkFqt
oy5otTZKQHCfD5N3LLyYvm8IL9wXWkJUjGOEaEMQZkclEpm/n2AEqtpxX7EWHfTFQXaJ/40WQ92r
v21yE+NACLqzfraKPrVI3gxUYdkeBRi3yeHcTQw2EkS35iqWzFhGGg+f/Z1e5YrVN1AJz1vinhaW
QtZwWJesszwgp7rtVHb9sTvodzxqnPxdqz6dkrZdMprm1zcWP6+x5kZbbry4s9ACDf/ZKVN77Jwh
LZtjqAmVSs04HeNun8JNqsQLP7dQ2xmOXpH6DB34IBho12sQBH4lqA2NVD2rBfjDKr6ONn2hPO6z
raIRkulHR/s3VqMlia3EtaBtsApp/YbJ06t94l9q2ISNucP1GvtcpY+Ie01RctPTQIOY+sSwOpn6
5pHEUmJ8HjJ6T69gV6B/KzKdsSWJc3wpStaq3DCMzSuRN2y6dtukkLRr2qNvKcuoS1lZ9QjKRXvU
KUWItV8XjTUQc3fk9TQEqJLYZvkAAiiYh6MhvDT4Dl/sv+GCHyY4mZkYK8fmezAjlj2tcr8YRhNW
lw1KSSnIBva3Ox6g2yKF8bP4+hvpVdK7Mnw0Acl8skPlTbTLVap2Nhei/D4Xtn4GG8hhuaGy4OyM
B8h47E5d2ZGynu6mZ6sJdYQBMXI6RWVNPMucwoVGwi6ohJNlimvM1E2jaInmf51lBMceUxqofpUY
bRWHVywHWTdpwFBU8+zD2X3rjdcd9BCekOkl0OawXC5O5c+dxPbsT2riBjpcWo5P+4/Bw3dMnqkU
Naalq4tufuySB4RN8ceBbKkhYspUeAq8KY5f4JMrMPUGQ9JbPf7Yjo2YECsEgLFj0h8y4bafboHk
XVWM+/yHPH+WObENxSZwiLc03bo+rvhab01R1DAd+BX1WFcRYM7ujviWTd0wWIu+1q8FGDaz+ET1
qSKJbozfRx4SnS4dkRDFsdADFbdhKQP864NekM5dQTXiSrwF8RMPhAJPtbVqTBdB+p24xN1J+WP9
hqkSHy7FKJADnO/HkfisEYtRtAWAqhmXLnDuJqEnnSRcggQq7zkJXeEuuVtQzsT7i2fOlLJNG2r7
Jc9katF7umLuNrQLyBWKEAAWtwulTRf/fLxXlYwZr/BDvY2Oi2fg85k3EiMca35A2Oudke8JWPGn
R9/AZPc4NuV5CYC25fMG0154ydmFruG7Ee/UxnUTNEaHsoOksISGyGchMPpaT83jsLmNPJS7etiz
Pg23UvqniptPCoIEdWiF1w2+vxGMgi78wg8wRNn7o+j45JjTogzi0OW7zfMi3koG59yvj8Ra8Ieb
u1zgaQ8Zy8BCEcmkxZHw222JquDFu3iD49QS218yWSRUR/Rpil0DFX12U5xVEdLxfMCPmOaORWvz
MdzTQESuZ6wFvVmCsNm2bjclTW6RIy78XtF0UwwIu2YAikB+dItkequs8bVWx/QpV8TEQt6bkwuw
Epyr2x9RW03FftFkl7a4GSxI4TlpizpElIvXF5XvUDvxY+wFqK6L+wPsqULXyYHsa+Nk+VZGdhlG
i6Z1ZSazJ5SEMMB/AclVMQZyVUWfhvXROYel6W6Wuexl4WMq6WAbkuiGJ5BQYwzuZOPMi4NQIPR4
gDLPj9kYiItO3ven/I7vb0FKGbeNLZgt4pHWhSkHvYfvxZe5r9uPLmTDSWkZKpB2F50jACzUREUX
5XxIWd9XO0AB2YpNfSIVvr/wmJcfbQHXELeNz01CMnOVZfGSg51RIu4uXB2mqpF+fg35q5pRQFVf
pJRns9bnj6jwsZda+2yzc7V76uZvAsGgzNA8DMCCVN+OT4gCGwyp0mJIgKBOEhOcJjQT24G2TPAF
Pgd/diQrED/BYmhh/IZzlQmPLRWh6RasYu1MKv7Cof2ubHmqgDXlp+WFPykTk+tmX8oQedb4/i6f
Jr39k/xYNS9rhZSTJih+Ji896zxM3SEUrOdsXEaYc+1/WyN6D5gmWfrzV4m79wRnj/zGiahurwbz
uRvl26RuFT890Ll4FCso1jt3HaGunX8s4XsSQocrLytb6hg5LKgBdyjNXo9aMxdD/ZQE2vWLvedl
mhpNFNRLs1BXRy6eipo4wBew7eVUeM5xTqsM7YQ2y3KXScWkGlThFmcOxTqVdEa7mXYWLYgpeWR+
7Ha3jewGtqFq1RwNPWcHyqC2yy968bGYfCVIT+JIMFOHrlYj61OxhTa1EfMg8GpGGCVMKSpcV25j
NnsOcrYztoDMTYh8BrCjjp/6WaNd6HwfYEybym5WF++yxGQZCePlFaoQboWbrcrjMc7kU/wZ4xxz
qToBXDCWlHS5xz84GKVBQT5VwaCM8H1R7k14cUmNmOG0Uy/wLQ3Ns6krR7BnmM1/Xxlz/C+bivnW
0lwVmqeaJQRPbFTFIkIB8/Fpnw516PHqSZFQKBfC55HTjQmZNADwUDi64FQQpmjWtclXZxX2phaO
PENWN6auexn/dwMbuyD+NTRjC6ypwcHQSPh7ErUvsk7FGdFo+Osqeb2dWjQgLW9vHvaY06/Tks6W
Wg3+vCuYsmsHcYHIdpedXkQ7HV9CCn+7wsI4Zve875+X/y8mWbwzXYpieGeMklqjgiFzT6vst6Os
7+CCL+GOcag2F9QXnoTr7JUjBYFxXBiJz2BAhEa/RGkknNVZfAB8JOcEJa+QzyUY5BVYWQTIPL8z
w/M68vlszD8pUBFSIuBBI9PFThXM+EpcekDmj3sgt7PpHHIwYHufRGB5fG5SQVUVOwjd2whaWnkO
ewtZ8nqSdEVMakywE3xlN4Sc6bfHFQLQf/GuAFbD8jL3o9o2OhrFFsLzzPnwn28vhcH4qpD/EDhX
LOeqa2VGaAwQtDx/qwu72dUNugAyNRmM9g6Mj3ojb+jXiOFJYNtyCYSCgg/oc74G/lYFO4Bcc7Wz
tM0+pM5NrLboLDe9ZItOLGguN7FON5JOrpm3pw//9PkWjRNUxFkf5UiPQPOZCFMDtL4zo4tk0u7l
nQnRvgoK8Q9mzzfU7OAssk/0w9jNFuP4gkVkbHiKZ2Q9kb+cX6Xqpvf2fYLpUutjRa0w4qgc7daf
lRIwu6eZ6HBOeMR6hz9M0KsxF0u74TVoP96zX/muP5TUYK+NYTCfPgOyfqG8UZCD67sslzrzld1J
gPVFcQ6MTb6RpwVHcIUQTewF7/fz6TB0+/l/q6rSbHR72b5+XXKfrj/mykxCJ5ZTkCH3AxosJb8w
mykzcXyaEy9VmbJ5qMj3WsqMU3rcxp9eYdguB/RuGx9uEmisgrdkX90lTh/I0XkY05DZzoHsB6Js
OKGXbTQ/tvauKJv/dmqPIvJWIzljhdb4v5QtYdMb1QLZTzX3E/8/Noi7OgAAjMhWmjCfMgt714rP
LTtx4w+WhYD4sGwGNdqySs9240TmCx+cwqbnRHNxhFNXl52G7WOuFXoOQg0KDk51CNlpeiUbJUtY
UafiwLREZSwSnqT2qTW+Q8Nuv0aICFtDMo0+AES3GE0vQLYgFgKAghNONJP/lKdVNlgyEszY4bCi
QvAFpZq5haG369jmZrszIrFyHnmHyLfIswmvI6M1U3GEf2Kk7mRdtcZ0jU/Vs4BW3xRXn59hvRnx
P2mmddI1JskNfduKytH3WmW+aouG7hHPzyrB3pCXXTPWAkDRd3WZYqvE4yDdyG2+H3Ef7xQ1izLf
EV/KnSrcuPuMI/l6eLY/2ibe9vKY183/dEhdoGAFhOkEpNNyVsjfYdmRbOUoKlOCgSk9bMWS2SXr
DJvAckrR64aEw9GUWvkJMJo7JRmSp+8r4iiCAfpvyTi+fYyzHADXIC16J0Nk+cuHDsdnLsFGK3sZ
AUOhNweLgG3IFeK07/nbaJF2OGAP4AkEdrvf5uOkiWuJLCY2BqeoUNdlhByJsBEo/afXrEWMkTFE
mxTkkmyEwqy1kFkVm3kE3IGIebXECy7hvMV+k620356z49nbjz6dmOMiQbrV7p0pQFs4O4hEhE0H
6q64akR4FInjsze3M2gPjkCE0y4FOskGKjUJsF2jTyce9s0B9CxClBnpVEFbX4FbrFca1gPAY9Oi
IM9RybVk4LIBTGidaSsmajzrO7rhOMECUSidSbuuK7/J8cCP+nQlrBgT0mpZZsW8P1TpIlSgU4V7
xHFcWNDm9/0BxGwONlIOTF8ACn3L0sWBCpryImK21oc13mE8KtpAQsp/eCUKnPf0+I+dvAniDWqh
pI9V8RZ00Kx3ABmK0GKdvYi+xy8KmX38YNXs+ikLQwDdcJJPBlI9MqyMiFbXqhMguC/Pr+/2bl1p
zDkMbi3L+wWRYvlOggLCEvZWWrZTKbhgGwbYDIUUhb9qK7rJsJSLmAjNmQ5Qflnt1V2snYw4+NpR
sodbbQfPa1bCQ/Ov/fNJJzNKJe72DlQg3Oq4+PpdQ+v8fi09f/pCjAqRr2xFvrAYxGeiavuLzU1l
g1qNcPf192tFiWk/V4Vz6cROTnHZpbn+8lwCVXlIfdPMTVcJ++ZeVVY70fsrZRMY/C2yhsrwKNED
Z2j49LHznZtuDono1frIJdKJhyt0YDeqMUngE1VaA8ricyTS2P7p2UdnRBneLEQR7FfrLByuW7S+
4d1s4IpQfLUgCkC16Dc0bZMcAE7ydKDc/IBeLk6TaA5Wz5vCpeNH3dd1MZ6cb2x4UT8AauEESgbA
KPjbd2lCZsOmJr8KxWmeVcI2X9k30N9HG/aQzeohMBPXrhSmgqD4c431oUSJIqgEdeRieMMLhcws
GvrKEzQ/TP8pbZYQTARLbwAtesoVLvWWuiUmJ9ExwNXGIexWC85CH+4aN6x98AeoFL0gvNdxB0+V
zDH+SAJa6Iaouzk3Z5dypXIf1NfhtzrSOf2le5pHbL1J9mecgPQl7YHRqTuZU6E419TY0GLn81Ub
6gKJjxi0fI7rS/MO4oedFVfhiuJcTKsjeHb1lhySjtOtmNLOHp1Pkz9QPV5frSeUwk0PAJgt0BH2
USMch+xJuH56FKSqENsDKID/K25/LPXdZlMQrU6+fWz9BJj5T9aAzHuCKfuBrrAJFMBVODTLdsZB
ZO/ynxB5jcVwo1G/NC8CZf0NjOOPFx6pYYbbu8M7VjP6UW0R1GTLj9hNWwQwkLCS42k3y5ySoviP
diM5JbdPNOmnzW/PgZw4H26dUOr59TgzWeGPmmICkV48o7pEfxvvzeHttQEHPFL10iJGC0MyMdF5
2hiQ4W7lNvC7We7KR+hUIo542v4/JmCxyC9r2Q8cHzP5l4z4AOWmlFeGk3CXPA0IFGP/uNb978Xv
5E1I4BfAba7mpJJiMcd4ZG1KVNfp6U2Hv8SWLKfsvZ9xgKnRtdZ/jN5eT9ZGZw92q7IazouZMG3/
28vwfHTvmCOJnqcjAmjN6s8OBr0yfwwH1jDan4UodLBeOkoiJ5mE6uWt7Ymg0SMMu5irEYN0tFWu
dOhQxC9ojM8S6W1gX8w3mpboUtQ2x+urOH+pvUfX7xZIbJo2TgS5dJ84oTW0yTHGevUib8Lh6/kK
GXxgSoEWKhTFx6qFNd4rGSXn9YiOe2hdXxOf9zG0SVz+TgyD4e4vTkcy3iH3T/OEq4kZRADfmGBN
87b3JXsjXJVe7UmVNMYEpulfW8vWzWZBh3xeTt/PSE8XCICzU4EGjRsxDv5HdaN88RH9U+XPh91m
PgC1OUvCsK0mUBZ5NnurpyQAkhHzlpunWJDiXeHTbcAZE6g20QFGBIGJHW+W09RxBB620ljlfIuT
JugnhJJDpkdq4MCJW9h+4KD6OfzNLTo4ZN88gvWQqUF0NQJ1ROjPVefkZBpVRCWl9lBNNPlf8gz8
FPKv7BBqebVgZ2vM+2mfyQJHXOIEpeuMoXF5e9hYElXSs6Z9iTHuiiEEhjSzlI+0auVeMBcQ5QBN
312p7XAPQbLgzEGgR8QlW7jLhsKBNKs6aZUtWwY6GXFaW0iFK2ldYwSU0UWyJfCC9FBnNlTFEjN7
UnUDMM+TXnbfx2QViez0+sRv/EhDBCvVqDhTH2edGczJ2hBIrl6dQEOTYVEw8FPfbZ5/GxEyUvFx
OwDfnehV2bVST1vl4pFuAH1SY1Ov4fnnS9o6u22mNZKcH8ehlA1sahOWKMgNWa8BTDtK492wZodL
OU/7y/lovCcYOGgAmQFCL9scl9uAv7Kq7sHcSrROejjRm2YMdrMF4mEK3peN+xFh+4V4xBMQGexv
WJBzPbEAgbq5lAVvVWyQEWjhFj8ihb2F5P+EKbVYSNcs7W7dpcCPTJoGLS5lDrJ0i6/eVfFaplkD
qnAk5ukAOf+OhyDIQ0bWaEUhYeWMxmKSnX3CKCobO11OL7dOI5wo5NLoe/pz35HjmIAFPn6v/5dr
fmp8Fb728Lpl+s8mNBvml7dSaT3MtTnEE4li4hNkLRvOk2cE8V6A40brTpie3ufIu5D8jLxRhKH7
D8scaHO0QkudYkMhflzZytPGZB1vCXmuI2vMt1xQ54z3M5U7oHEiJM5ozQcxxGY8StxBvtQ47Jp7
mzm9hDAXNJtLSdNU05kHLbJDH//yRjI5kekBDQFYABzlS4nrAzTk/pfAxcO7lnoyqrtEgaVViuoQ
B/8cob5rCrCERIpi5p9/VoNKZ7zSrAduoHAQDo9UYWx+XDJbbY3qv93qNFTgc8+cUf2uZaArWFrA
kbLOMGhew69ZDN5S7CTLgFiVxAdUHxeKNcf3mUzV3pp7GPGxN/sUmnlQMIkxbl0+ia/FQwLi4DgE
2nPwGVpG3tpK8neWh+8cdMjCBO9nZfxPp4JDuC/0DgW7dPwGy7k/MuqI4mv1DOzhwdp+NA/w4ApR
lj06m+fUo6IKNkSyPaxN7s2r1mrw0taTxUV4LWEAVlgFN2r+dI680dEq8nG96GOQzk4U5VnMIotA
wnCeK6PGppelZls41wP28QbMsr7lk5AF7OSCTpIhvyauxCTe19Pkw4mtsLmcRVZflGo8hA4u68/2
pxPgWM1m625+0abvoRNNvYbSfFXgmVRCVZcX8+mD8WD3v1c0JmzApN8bQEYbOfEH1WrLp6Ex/iel
YmcTDTNp0HKOCSGfJac9Sl9YBCXyIzALq5GWUrtb86Wc+PbfG5dGmHZLzHKyChzDH1m6sZR9x9XQ
OUXdv7YCSgdjCP/FS7P4ZA4m4qOlvYvMl/MFnXxiM63yvULJBXwKGkgTDpqFOmkFEwH93jg1xx/V
pZOWKIMeO4L/6RLWsUzMLq4NsuMYxSW4oyXY4svJuHImRKX5hdaAOAzRRxSjRD8OOKW66E4L0D49
xA0pvrgP5Goe+3suP6zewIKD2BsTxZZu2cdhB0bXFdWJmnGwV/3Y/XWOk9drpJdjkW6f82my88eq
XpMgYxlQjg/jVy+SfWgIVKjDhgX1iVqVJS7T6FbrEB5Sg5Jt0AzLpDANEOupsa7JcmYZUrWOmJ8E
cVgIng6zguA6Y6et4QeghHKeAa5x7WTiww18l+aQ7vIrOPhjF0RBucs6IuuIU2l5nJRP//zz3Nhq
S/TClWOqywN1z0odQvwYKHO9XPgamWmmSl8pKHlC+lmzINecmCwQp23A4xIEWSJybKxwl/fXIdUJ
laa1ANbfEFsOCysb/8E+6IcdVBdz8t6ed/scCJke1swEoWvyQYAG2oMoeTyc5AnID2f1XGTWf80u
G/o2iOdWZ3xvfjzFRcxfL7n1RishI257i+iP87YVtg6iE8dGJUZdd+CwNvnbaoTgDh28R5hDI47b
jCQNNZVd9WaQlkPyhcsmlccsYilmgiLSDQtO4yKE8awUhJMXisKUN2zrEhkD+ULNUTNj8xpKt1Jf
kHB1hqllbpyD+JJQTW1PoupFZBh5FBIHnRVVzakOYIGXnAyPFI6plbycp38siThUZCvv5XF9lYpH
Fxe17EaPEtWrpHclLy0oNCGgCWPps1m2pmRNPc/vN7+fDbkuwLOigbMM9NJbDtWsID8vh9Dv5yGp
APXiC5FQbnX8mqZhqABGuAwMDZZMBCggvNIyTTEUAij57hkQsnp+Wp8yvRcy/Zy+lAqqWGUyPLok
OWZBfC1ejzRYUoLWr1Z1NwmV0cawIBc4QYB2AZE7Rg+vqBZbd6NXzjz38Lmz12MEHLQwGx0nZSXY
n++a5C7+yevLZLc11l80K7QAUJm0z5RX1OAZSvCmF+E4rjw5x+RP/OoEpHXL7OpMai5dMlk5683G
AYpdOT+bFF5vYekeqhJkBk/F5cVd3wkQ8w1av3Lt6hXmw4ztEORGe74+hDvHB6x5P0vlOk5yCORM
U9cNuJ/SGX2495X1zjrZC5/9xUctaFUKTFkmh4BcjdJGjvEhobNlPgHkQsMUAFVmYZaRBBFqfkgp
M/3Iibyf0P0vWlXXanK8KO/ORU6RAJgegjOAJ+tqdBFD3NR4UO/ITJH7UWWdk+4yjpKCUU89JXfD
rPiEPG7vtqyEOUUyVyzKefwZAxObaWx9Vwjbx/APC2+9+kb2OJOADLvvpDDUvZrp7PmlIRVGViBx
sI17UuLNsZ8J9EsOXQfybKqh98HaE9YGM3o2w/+LkizVJpBYCcphwHn+VjMrHV+i6AV5QVHSZlVP
nC1CcAMaour4vxSDfXl/Ls5JveNRhZZpsrlNPfSaVEqV2hJPXwFVZRoX7AqFTf3zJptqd8Ij8GX3
vhJTajGINrvSLcVLrapEqrK/aXD28QIy1m6McheDEuHW1sNaNjzbnhKz0m8exQCS7vKmqXsoVI03
Fk3FJFB/wNWmzKx+1MsPYLU4N0PzzvR9vFnjutNbeep7Dvrqd827MQsO2vxCx0SzGvi6KtVcPd/W
vvic4n2euCso65pePc2Eq5vKDGuwcGT36ppur/Xc7e/gVQOxRgQyzphmQIjBZo9dsKVYVK8aHjYN
6pC8sfpiiBD564voHbnAxMwhSc8ddwx7VVjkZcVCWXn4/ausNbI2EqZOx6awH76MR+5vsrBtVVxB
hl+tGD+kKo09/6c6FIjahyU/7uTB6BHALqT9WvppkQ10sRntrbnk06PjkJuVESWCN5oRt1NPHYYH
xWfI/E06peRz6jHYkuS3HBS1C5kcMMrx8rL2w3xaA8rzbX1+Y+TH9kpDGZu2SHFZEzysC33EvRkf
2Nar6M/UDKOCx1zLBsJ7xliXQ47punDZPbqEXcCJXwM/pw2bc/wcHGYr4yKLJquesFJ3xW7rC59W
BmG9AULM48yJQwNxDDU/QfBegfIinIF+Sdg0LY+2s1Ejnwtsecl3EgWmoyRrElNW7TI/IIn4jsej
YyK8CvT9BbRrR6ivY5eeUDMap3Cazj+rozJzZBPNC8/EOpmzSB8s+aHhaYTDafnLqrAhDj6pbJag
U3bZCfPs/khcFQRSAF/MICOWuacxoG07aDaeD3Ky+Jfhe9pFAYxBswdhine5UkljA4b89Dsnq39K
kNVm8+dvi7A+ZObZDFzPUZBznnF2qqR7gcrHASWddm8+7ORXUWeehUgI8EZSYLcRqiYJlVBvM2Di
WlRjTz8bwcARiN9owC9H4/GQ9aA3TffHxB2jcA4+Qy0kEZWE+HVcCuo4AMeWyJKvNehCVwGBlDor
3jovqQ0ZSKlkOhoYV8xmp1uJ6IWO9WI/PZisz5/US4TMO61XC9iIdvoC1+JP9mbrX/eaREgSbD8o
2HeUEDn3oO1bBUgBiVjX24M7nd11wNLExwS6Fbyhpn4XDowxeHLSdo3/ijbZejqbYvJTa9ivBLG8
VkbzU4Qvqyiu4IMl4Ocfb7DiPVtrWEvjOacvf8NQRSDHwGJNXHJevs9PRKyTxn9kB0TfYiBhsKA7
/pNNyb6Ox5GYBxg1fTZoscq94vfx4eVLXLzgvm+fysy52+FYhEUVwyG3kc59PaWFsDDG+mA0c4NP
IAfYiMb2YQf8n1v7B6GH+N584FeKtbOPvk7g6oRpMx1JlKQhpXgVZvbH0HHjKxbmjkKuZTIZ2KiW
1GtG5ynHYuJmlZNP0vdnTLYG/1xLT4Z1tS0wZxMU7IS+0OJcGxQlBdELwPMZb6EDuRiGJ3k+wOjv
PxeF8Zaa7tKCWKP36ZWnS7oLRbCcQIp9nk7VcqBICixjgoQxmhK1WLleSUsLuADGl2WQhuwCk+lv
VscEgKucpjhsw6PWOVCJi7Gyi1MdVSAHRUDEB74GAVW/Op2kgVGsQCNtTSSUBM6ZnTGfTrZmRkj7
f/D67PkhyueTDa12NrjGFKIQ73mMpX/CQ/sKfwjrzsbh5cuVd4uNWW2/a0zzyFO9ZTyGX/93JaOf
EFno0kIH76k5h/w9h4oT0j8+BCuMjCQYrpI3Cad+Rodsc5FBxPncwEBZcViskGh5XWzBer1VNIET
5RGVnZyst8h7p4DrC3/a+zhELs4BXnGUAsoR5ymMJRYJ7juyC+/OAI8+/RiWOGbbftRlZVYLJdyZ
CN3eGtXHb5Em2TWOHCi7T8CXBvEg+KUlTuSt7FoM9OFtpDZqgV150ecZh0huE9EArqMUWaG5Y31H
kFu0nToHcTo+sOQ/ReHZDbfCmP1ukSWK4e+lZW5xS9PIdyZQ3v4DOO5vVpgcSLJvROvMswzCTOuV
x0r6nlAyZ0gUZqnL/CkT9lhEpaAqqM5EcGa6CBPr7FpO/UmtwI6swQ5IJNaZJcvOVTjyMo4V1v8s
MqEYbLlGMZbJP+RSVykUbfjFP2loen6kl42LX/UO7jzdjyAcTD7sc53k3JLkgEC32Y4M22zR13mP
blmEYbyye6yWbMO9Qg7Sd0r6Y3oQv06lU6IfUw5E8o/Ef1U5xE91Gw7VbGewGHxpj/CbjCS8i20i
v5lKQ4rxBfU76OyqmKDJP0qPufRcNvaQZMOGQVw+YHSo79Fegx5B0b+d+38hr1cpqr3+E9R73guY
FFVWwP7+FqD6keEpaSpaBrDoUv725sgWrNjfRpzdD2vXnRfoeC4XfypVnrQNNN8LLYW59+vHYezS
Nc2pAGFviFUr4L53m4EHBLbG4mUBNGpPflU7FmH27pA+SEFFL08yBVw5TRa5a+v3td5kUl7mPqEX
HyMpKTDRDAo3VUVYiNcpeWbW0w3NEsazUjhgIspUAydTJIDlWxmUXncNaAw/nHg79VRouUAKw+xC
YdH8WLQEkk4zySenrM6DI27xslElLGrvF9yBFtWYXcqRNXuYHvjS5zWLxXnVoto/m6FVj+yaLhQn
CVcdMzaMw95wc5m65JdKB1J+W4G20S8Xj3ssP0jhrjKk+zgqMh7WImMi+QK/SnN2PGWzFTdFx6b8
er5vdx3kVeuGvCgwMAUjmjIbFqEtT9el9fokxs2vc1+HspBRMHZm1MBEJkReLaL9FQ3BXSVo8xY3
KL1NZEUU7ZvDkCMLFp/tvQiwwVomWzGbZuzkRCNv99gXMjSnQs2vqWFDOBolngPV4V2lGCOy2sS/
rPoX2n5qEoegCK62ObCvitid8WylFpl8iKCHDgUGWjRAhykDWzgKm9n9tSKeuXm734Yph/MGwpq0
qACPbnp+rgWr+yW6Mnmc2zHH7P8Qjn9op9iuvT5URpAEZvfLiBIpJz9ZtSfqNBF11j+3LwafHhTY
L/EU4BBAGZpRcadTzE9vzD5l3SyYCJgXLmtIoemWwiDyNPMGMHYDM7AsnxMTLn6I7mpv3DkdYvTU
JNEb0mTOLqYeaTqnLdlSyV1bHTQAZmhjTIGiPOWaQyZhd4t3lcXMy3TnQQ92n2PtYJ3E63IPQQx7
iKKIxuJbw5ofHHRZ8Ksg2shjhW7p4ctldDAtefK6JAdr0GOair+05SjSWB+TZ4ZgsLBkBlq+0KUE
tDHDbUv4tfaiMRM14KCl7SZRlc28j5HL8ycE0BektV3fdjQATfMyiTr3mrEmPxWAOaiCoPyQmDSz
wL1qCRVuU5zqWglJkvltTh0QY4x7XCH9ge9/S/iD3mahYp4n4AluYf8D6u7ov3qt/KvytLB7WfeH
VHSVisrmXXsLOaAiZhtubWuIn9QsiKaC8WH2Mb0SAUasBPRN3Ggnu2tXyuKv/ZKl1lifDQmTrKgt
gqjNVoaSry2kuxrLsr+yVnSPOHxp9ED1NOXpfyQAld+KHUrBPZNdyHtJHf7m30kkQr0cAlZsbkr9
LlQ7kPjJSosCTebTw0S3LaRcrjPtyO98ybv21WvYG+Zwma69gdPeKwnPMcKD4tEKVovtvSa0MOwl
NthYb1XPjYSM7szMdA1Y6Z8A/soFaU0CHXWVJWbUMgKM7dAp/ZZ7v498hiU9zvtYLqVD5KRhpLvH
aIN6Cfk3kxcDfL5LwSZT45WJ6vne5qm7cHjZ8vKTq324sYNSljdPdbvvnXGXbtPe92ohkClcSDH7
d0d8S8m1AprAT73H5tVtFyJoxXm1/LJhG7IfvGDEoZr2dvjYzvnQ831EB/EveoNVkwD4N7I+XL6r
gYkDpcre2ur11ELUEFk25cAxIwwsRpn1kj6upfs8eBLkdDcTPAR0eEyscBc6ROkb8dHQVpsgoQ3A
A2VTae2g76NpLQc8SlbQAtWxuJHjchmXyLXomrLtwmIJbDqYDDOmJV2bkSgDVRj0ZnUE+fDNQoYl
KMibxis4/O/qs+l9IelnfZRbq1W90p1A2XtSYHGx28xt7xv/dMn8vbWrLpQY4o9d0eT59BRIRJpK
GXyea/b4PINXiVYzy8nG18ZyJiZxOCtBKoIx7iM+zWP677paXHmj61purXEv9dJiku6eJf8MRZ3w
X8m+DSCg/QY9gqLfLFQ5fjwMi7Ray7iIrSUIPkWe2U7BIB8XXG+ix6D1C0Z+H9OzeUVGccZWVhaO
9jmLh5ZSI81YMf7/LruO7T+Wc4mMDLmIleIi9ZD0YIxYwnDKhAQ4Dt7VfE0jmMkvSKuMCQ8gDQcP
ITTzreSHoXxIv/zFmnRdP2DkykcDkmX4gArh+rQrHK1RuwbpSocG/Nrax09uD2ShfOi+7yTCPBsL
kT8Ujn8b3R5nlKAY+RwO4PfhzQAtv+DoHPkSEBEaXAhDphuzfgwGYpNVNkdkL3bWoDOvLUDexpLv
iLtQ4/TcPw8VTzTRKZ2w9AR/iAZpZUteinV903ilPfBFx4UYR/Ct+LNoYKnVxXh3ljY/FyiclxBN
lSrD45zqftb6fO9ZuCFcOATX33mgq8o83hJIFHGsDgWwkWNVeloAlHf47zevR9BdYvTyGVzavjTD
i2Bf3eMcIKhCDgjcSXQjpfBWHffVtfZ904hFgtHaw/plEm11TEzyaR48bmzo0jZ87uTI+T6gHvAp
7EhlFexwHjfeIjnyJjMt9IXot91YAewlFq9gcULwtZCbkMeo6JFbMsNHfCPvmzRDXEH62L+xtLTT
91v5RG67Y6/L/uzmTzx2699RLXuB6xttdIlxhpiUhadgA6LfmDzMz4CuRC8V/Mgy2+ARMZ97P4kC
BNS/O8aNb2XrsJ+64Gaua98RZFs9OBcU+0viz5X31H/c4GZTqpF46osFYUoJ0fz9rBtjBaliu0/Q
ZKFGG2F2a3+Xzuk7NrghdnKO67IQcgyGAIzpn2g0FR/rslMP0VQVKPSHBOkUJxnwQXaEkD5o/hmq
TIl7s+JXoGxxXliRIekS714qp+JwSm7G+yM1jiEealmchGIgs81H2kbXyJ9X0w8A/8s5+FLTz03P
qSUDiKUqdfhVhwg9v6DSCjNjyZOj75kj6GOF8CFm5mkphdQ8G7yJ322CGJ4l5/hqczgznZ8iDh+c
gHJONIuhZAQ6arN8j8B0sRM7/FUAolTrZVdljYUJQUt3XAWqj2FqfrRSU6TlOWklR7eKQeGNjp0P
8F4eoxXi1PFpDj02KyQP52kRMKaLSTe+Jx7q6gJD8ukd03MxR9rHTHFJGmpyPn13LFs8wVHw/KMl
T+FANW2sbNrqyguW0MWlDEwMsMWDjVtKmr/3QdAf55SS0hk8B8/QJjNLxuYkQDjI4CHr6eqS7tkV
kpMdkLcdMSCU39vkg4wzTirHfdmiLQheIQPQcf3hluL/n1wJeggnoQ9cTF0ys1B5wQV2AXXrdMaY
YuV6L9Asue3521QSPNJ6qvRVk4j8RAsTXpGySJZ0WmsGla9KrQXrXRIUYdEDXeA5qaiQn6qrMtkT
FzcnQCe9vExbY4zYChcFk0Z9dU1ACBGffuQBoZsohef2Ngf3P4bXZRTgwEAu0R+kO8WCunrr1uX5
eJPIsAYmr8tQfThLDRLGB2+92cHd3occe3+WuZdH/MupyAf5pWV6xQNSRb+422xrx+YehjAyMO+C
x4g/vXtRdFNSIrt3K+G2UWR+V6Wj7PTn6zRBOU5i1rccUppqIp9P8S+eN3lKScLKJ5aMyJ+fksVj
HhhrW7jA2vJsRHoNI80o8yfjiwd9Qp9g2s1JaP+O2HV/t4MtMgyJ+S1U2pOa8Y7FW2cj22r+FZ+N
LQVwgtl2Wf7G1dYpdNBbItSFSL+6QkJ268j4757lX0ZUtfU+yxOaAu/9wu8ZwBkNPTbdGs2g+j9c
kEWK6y0U/haOhtnQjEQHx6ML3orBp3nEZh6vIcEwjrYChAzpEXV/RzV8fYDVrnzeHrYo4Tm/fnlM
LOHTPLDQhjUNIwVb9D4cPlVdfKetwDJMOKpdPEx8yLuAneA/KSuxcex7T/IPrqcaJ75AyBLNp4w2
uVs83KXKTtyJLyK5R/g76sLdaRcdDmimnWOj3kN8KIMxV09+4lFB4C+z6OKLggQgR9+fBWlwl0ms
zOMarr0RSZr1duAB9JJ1IWxHE4lfA3RO8wUsZw/0Hm1sXfark9hBXxcW8uuY+JROTU6HZIHbpdpx
Lint0KEAc466VivcwMKEF+ccCfrY7bPEg3YSkfBw6PSFRcI2r4u8wxzGroTMbrwE/PkgloyquItz
xK7hgi/u010NRi+MTBy4OhfcDNSgPkPacUNIIT1nKtN6qdKP1OkItMk6vf60hoVFxyyDLwbrnpy/
ySrkq5Km12o/9cpPrzB+1jy3yygl+MTpeVqANAFqGENzOBqt5WOSRir3z0u5p403Y6Nj+dr5tqIW
WwF+ysxVAUWQdBgYvECjxV1Q7rPEHi4jzdwrM25KP1yIOae4V3Gld79yTC+/UFm7lLYIcOeqoY0V
+KWB/ybhUyspih8BfqKzGy2KrKdBXRUZjQM2sFE9ftX18DQVq2BmOIRTbDZF55Y9rayqzyOUTnfX
DBFoOPXMWk6aEhgz2jcH9JhyZ8IxnFacbYeOukk420TwZiNZTY+/vAo6clAfjL4qkLoebTC9aOwd
aTD3NB1TJrzhbyawXrPhaD9U25FjgMUw6kikQwKo1vDChGrAthBuE+1xwTeB3xG78tC66pgr7hd9
nxo8f1rvHdUqCyfVtyKsdR0gggELS/N2jrWleWG3UmdRXmV2BWx0xjqu7s956Uck6pESrGBpywAl
KKE2FCYKZ/3kOQCNQedeSuqqMQGrdFqkAjEHTX9LyCoojetL5wdilPxRdCOY4jLbn+c/TLWxnFeb
bdCyf5/D81xUr1uLHMDH8YzfgHxp68dAcV+MhoYT/YmoqteBQo4KqOmGaU79Y0IPz0nJbCSLRwdw
6qtC1N9MsrdsXsXZE1zMAgaOHOtK6ea3uG/74qBrE58Ya/7OYjueu+VF430iA92h0S7eroaDPSK2
HL8DaLksRg5bQfauFJVQ2VOx3dnHmiHSgop2Va5rwV6WbJwh+xZxbOJINcf3f1GziRf408G5Beqw
cWRXsBuxcPVHiVrhD6dxbwIfSzZB8+tsTD5Wxnlqjal6N03oUd32NUvy5fQpNsyxHW6aFYJGWOsy
2S6zUrArL+XXpi93JxoTsOnkFFq6j/0/LOLpjhBkNP4VcLILTdlzntb8GZrXcu7i+WVMaVhAfRXE
vnLbqGZz1+cWHyWY1C2reOdVtALLOwy4Qc+GTE/jwDFpEysxbAdvqmKQK0jnIgkDJ8kTi0JWvlNK
yHlpdg0s9tn6NCA+723Oyp31OQ+W82HhP9Mc/i/4yB4o0csQUBZCo18MVsE8eQTGy67rS69NjAza
R7ON/DIauSz+XUCf7Vd97t9e4T3yGtNejKVVXiD++xyJy+oiq0pi6VnBqqWX8bxEYKOXc6xUE1HK
X5OxU5/tUXjknMBV6UlSNPt2yQFGgtAG+M8xAHZYIgFpCWGByXdIGX5s1rOoycn93qdKuYpAgbxA
BwFlwgaFnms2lHRBOFZLubgGnu0dCBtDiGDcuoZTQLiRIi3eTwcF2zMKHrxSmzCok54JRd9IypQk
PcqpsUJCO14tiWU5wQwtLwLaHJbU/Gv3L+EWYOon1patVIygmmapo9F0bRg6XS2vzYhGi9mqkeUU
FyBZvGhfqXBfDGBbTX/WAIfVXCp/HAK/CQB8Scv98zY36WcDNWmqsz/CRSEHKsDSTrBGrUIMiKKq
RQ05ZkgT6cB5S0ai5UtHDO3UHLgO0qkDTu/TTbuYJ8aKmaicnEICDuO3IVKLqK0Yi6JDdsqD+BkW
AuVk7X48mNVy4eTQ8DqRQn3zTeNI5UZ2fJtXFt0uRXyS0OzM43a3Ywd4p7Sxh/oBGXtNF+bYSi5S
Kxx+jURnfGfY12FWvAC/mENBBqExe94EmWBU3RrL+YIFvfUuOXSMjimc8IOSapjYF8ARLu2FS4sb
IXpnfLTZB+qQ2KEhoekVkiGgUEYh4mSdjM6eV1KGYJL1rLzQNk2B94I0vmSl6Ju+qXs0mv0oHLwE
8Ojc4fwQR0nw+/zPRWArxQiAkCpD6V6RQpb1j4iazOtVjWng3WLLbzcOobuX30K5MbWJYBhekPfj
5ij8lcRfUaApwLFA74JkEoI/wyhZcOTHLrkDTJ39zDBZWbrHJOO4q0u2mnnK6wQ+B9fv0lif9kCJ
kRqngwmyWHBkcxN4bAhLWi8gc4wvRa/o8gfF/yORjtActdm8uDpxznMCtZwNaNJ+9dpleoGyzlDW
4zb73wbMZhj3z4+6OBC43DRUWEqwYbAZbB3U7OGN8vdx+iY4kJhA2qGuips0DwpUQj6jyYN/TPxN
4451cnbmGU2VM3bFu44osjeui3z9iwUkH1O/RiK8K9u/Lqy94wMVH6M/klgvBK9bOehZEe+KYZbD
7sZvr6k87p13/8NpT5XJ5AL4qR0DF8iWQFrE5RvrNdz9nASgxXN3TksUyEsNZ6XB3zRrIy+UkNkI
zWyR0pe6TzGYU5u70CXdVLLBycIS7A9AKGCGxg0AQENqLEmLlw1aW6NrGSdt47HCMIJrlyW5MBQ/
0WivtFOjNVhRn3rSr1RaOVIMdywTSvYMX7GiXg2pfLOu4xLQIyqosjpKfKTHxXp8AGYe80iAJ00g
yGID+nDtJsMltVUaUghcjd3+Fajf0gtZdJ9+DnrWHZ8/E1vy90vZ9r4F1zWdCHrtujZVA4aRpm+r
Nw1qfi2FGWzGDzTzNb4MFfugti557ErBCg4JT6ax+iyAAMOSF/XOP4FnAIvc2O+EthSFgE27FL2q
9VOgZW7Tn5qwYXqiAybyBl3oNahJvYIEDlOhHsqP7xqDm/+cgGYhyxB2cQt9xYkuPW9RTX8KnMtj
n7HUhuZWJ+huIepJKo8gmSKQSJvIlQ5DEByGM2kWkwqzWJwqlSz7bSSiKQQUMRPHi5QC5dEJcah2
kA2QSyNWRObt9W3f5W6qiK+XH344rb5agE7mBOuUdSdu2pF9ARF8Bke8Z3m0HgqaRC0bxCCdW20u
PkIrw9xt9iU6rDBSnRzZbMUlx55OQs1wFuud19oGTKVBL7WFmi+Mz5G4RSYW4TLxASQyuAWkSeN6
iV6W3iHqN5Ndo0cSgOZc9roCVPJkyfHAyeaChilGUsX9T1dhYrZh/Kr5IyvCz3si535xcESQ4WyH
UTupzN4xAzeiCWirjFw6h2JNSgDbyrjM4qUfJEaPpFUK6ih3G17rblPi9uP4pHCEZsqzhtZ66Rmt
VCBr5gV16er8JRwsIOW0z41SF76zHIIAHRgtAKzjxBTFGvMiRZGjsdKodrir/wN/Zjo90Hb+Vxcm
dZVwrXNdYuJupowJO/Lb117+3He7zl5oWO9WabpL/tqSv5lBFX7I2y6lVONudVbpn8K/cEl5+EKr
vluurEN8eSRf/7bFtT5fYaQWszUlja8ts/4jb2zDe5iS5DWI0+bwMmX6SFG1s1ZkZnw7uoABPt6L
dld60eOeF9zJoROX30XsNR/47TxCitje0GiJ12F+2L1exuJE58KWhcOBWt6NdbTJaF+5k3AQJ/g9
oZT0oAJSs57sSsUzGOX0PY1/gKwcLomhg6PMRkcctEFQLO1VOBN/W/hKkwWu6S2n69tv8v+5rgCP
1h5XLSrWQmQb8Xp9IkJCzNs8vMo4gJGXLdSgs4/As+kkI/D60jUBW8jBe3IEFHhUbagJuspH4Qa+
zUQXWXLcHx/WjEHuNc75P/SWSpFABmHFPeBBfriQ6+4IiosfPO1K9xb2KYq+jQ55GSlD8To+scM3
arZmcbU7EvyEkQwAV4coQg+kWo2xallsRg4MHq3hsFew6bQ2rVE8M3aGAMqKHGLuO2ui2fqEsSGr
+RyuQPf7onJiOn5mAKIYirNn6hIHnQoOp5xgQfNNS20vAmG4KNQuAnAfaWGvIYFfJpK5cpbPaecy
SlA/BluNMfpW/aXOD96lgOJ6u9Z4oS2+bvTjHu5famPvO7XW+/mJhAUbRc5Y1hnlwWpTXBIlBOIZ
HNK+mOtQfusXw8yNDWi0EeIWfTAv83v+taCJusf3bu8qyc4CWpuwxpAz0CXgEMx9qTqNvYfLN/3e
dzdatmsSxqNPgIeWMwfMP0H+3NDkEO2ksLydq+E4Ft7jzryMfq8y/UPGQmnNMj7Xyw02e+sUHAvW
NttAlnhNeO90uvItxg3uBf6ZVNllj1Dx93U3UjfFgUJAi8LKAmL1lhKjTzQn4HD0vN8ir6Etobp6
sQfcnhMjFKp4VrGmj88ps2Y2yRYGhZTlMSmyfWEv/b7KvPc2UsybAIVBlxzdtWna1O88qxtRKs80
qXqL8SZjrCxsBpyMAiq10E7N3/58OHRcJfJxFL+lWqhxLTzkjK4AXYn1CzAIal8XIlSEfPNB9QVp
x9klKuNK4ep++EYEhH0JBRD8uiDuYM6sU2f6uxzkhn67VKsuPKvPR/udBbkVbZNsL/soETgphTjY
3MpALH/gR/o+mOmM5EKY+Q80KlxbexIT7JTzA8r+Df3ENvcOjlmJb8rdPK1WiMZjtvDFsNjU6PI2
r8QaQtTgw7wbDY/itZhtWwuZt0shIDoRkiXrTDCOArTvTlCIMR7//Pj0gDxgUfLRhCr13GIq2E8+
TBYSgtInpTHfXn+Eld0iUF1SXMouL3KFowWpbqaMJ/q1TOpBetTKA0PFEWNmtaXG+mGqA6oHgmPB
LNMHCHLOAaoStptbkfs2pvv468FWLqm+esF9O6tv1jmxA/7R/BwhonKr3eZzOzZhCQ8X4HnSW/jP
zVFA5Bd9Rsc5kzkflQJwNy4JvT6cX0R85gG+I7+haCYYYjfEoVu0L+4KDi15bgCeGlni7evr8bmR
3hGCF1dE3HmkgyaJqSWNj6PnwbfdTSjmfI08BTmQZoodCrGwcDk9YiFfQzxEOyPGLG41Hbix2THo
hT7gN2MBAeUbpi3nyvhAdw3uy0YDhE9Yz+38XrtTASr2UZlMIYSKRefrOG3PICNYG9JHWrFBbuAO
nDgUs+9Hd55EQ9pjg7J94Q6I9g/cjuRVcI6sbBCnfw9wtv0Eye/Go0jaykDc0yqP/4foaTV6uA8e
C3C34sayUWIjxodeuRX1cVZqVGO/e9VgAvWnm2xsDGzGWfl3Sg5CpMWVXtDHrwQwBlzimahSkPsd
M2X834mR9tRwk017409LkfkwvJg2GxDvt40H9prW/bcjxBoOGnhgkubMVmMcP2Gj6iwd5+6hlKWM
jhdgjiHn0AB0HXRFDUtQxpSe4+TDxVkkGW21BT6p8EU1J3gDrd/laef/Tnu79amOsj7xmBLiWOjm
BovxAcKXip3YqZLH3zKpmDAdVFgikP5P6VbmhntulFWNecodCco5qRQ8W+w4Ujr4MPUtiT9yCGpx
4Ze+mDCMY7meciC/BDfjx/+UE6bTtoBwINaBU2r1N7GblsfPuY5ZqrzJCMRhTIoeHa8yuy/dNdUp
spUYBRfF13pZM4SAUeWaFrMhs8RNwlMr87uojvVNgWyqUdws39htC33oONqz9BlrexAH+/Va0rl3
uGTprO5XUWMT8a0dEocfQDAAUNivTM4EFhy2XH6IKBBs2WTHzXmxHJBD0KGyKRJ4OkXQSGwll8zC
QjYO3Gch0F56Z9Hs20aT1Wy6RLsrFUI4BTuvQXcFVlqya76cLr51kuyyJ//ezfmjKzvD42WULa9u
WuL3cJ2DKxJ5zM4G+lpGXsgqc2amlZfM9AUKIwSIMsJQRVYYF+Wgvk4r07cSvSU4ZLmqTL8gBf3i
wTOR5F2nVJgL9QTMk2invJNozfCa1xWAW6qylw+eeEE+XSFpNpbdu78Pqrz5RTH5f+6qJXBdx50f
89WyUlv9Hw6aM+3xh7wRUUQFXILPz5lzHjqCYnMqywtsX9AQnYwByaJ3BgEm08TkMux5JaPB+LcQ
HnPBb4DVqkxeJ1edj73bfWa9psOXXE2zzJT88vy3wKEGiwO2l0qbbSik19wqs8wVc/XWvn/qYA2l
qAJueiyau8S+TdWxTn2F5Qj4wTL3pC71AaStbyvjltm8Iw/WPe2p7OxiGNNQJGThdTnE1L2ADT/v
fBy4h7CZPW+d/nNgl8GYsh7tjsrOdiPGHbESkjF2IxEDY+TDaOGRviGHNPYsuiJnXS7Qv/e97OGI
gye/BZRpmlDa7wsN2mOWuip2BwAB2Wt7Ya+0G2u3Ze1HYlDIy5zqlG+r8RBb39bky2JP8cOPyJKG
bZigs1xsONNJBjQPkdSdX7rvLIDuiQJgBRQfWk0V0+eerF/9GSXgNp4N502K69/7OgO42SseNci4
/RHiXtD6/HulBAihdVcLi/BzImbQZRYOuc/Sw3wCfOqL8X9/dka3p0V04DN6zpJOwiTdpZ+cURxY
3/u/T68qK3fwRsWg6yoha7/cjAyQW3HG3tW/Mt22lbj4IiK+blETGvYXAMpMaY52uJaHHQE1dl9k
P8a/hfipTZnO+8WMAwI9jkyVqLT7RRJuRfwQUqWc24LvU56cyLj1GFKyvhsZuIgbor8zcK03o3YW
83IR7nABTeGzpA2ap55EwtXjVW3X2eJi97SJY7zZuyi3nlOUNv3GIfOJU+jcMPfHAFRPqs/qWF+S
BQI/4rBYX184i8aGnJaMvsysQgatR6xuOWw9YNQVgif1E6FNqJGeCRN8UvCNvD19M9FJMLcAATss
8bQn+uqXjJqTkimyRwkp8gFFwaBMDAlCo3aO8WBzive4NaXOadTS+MUTGZMsE1ImiQ7PH4QRAAg7
4U92yuSdMuPbyTcZMbqTwKBS+MQu+jt9enwBqXbC23VdZccXnMp1RWYt36YYozaSdEW4zdHK4IkE
FE9gpP56xD3I8UBES3CNMEBNiEm3jWdwbaSQRQfRTs7vn13CGSbeBKYAulVJ8mjP+RC8adRu9qLi
Mkm5Z4EiN/s0ir06GgEo6Fh/S5PjIg90uDNV7dO5xAVM/Ur70DKMHb/grpenusqniyVsfzM3olDE
jkWmy2ilasXcG7Xy4p9QXBr+lnL6cfp8e/pPIL+j60cETLb6Alo19OsWsvy/TbdhUIAO9kgYi2a3
Zi78IUUdRLiJ2gFbX+aCe1O6qxxz9ZtWzxGviYL5DU25ibFaMNvbVp5hDp/QlVmVwdjRGEq/dVZq
+IE7DX4KCexNsnE4w/+/PSi2Y9zdHuJb7arpQHM8yS1S9TILqWTYVkT8ZL7Pt3kc+6Y4r5kHWBxk
rjqwMXZc8iHBojNlH5OI7XshvOnch4k0MBxU9VKV8jCohppwIlfdgczwCUX0ktKvmmYE9gspSo52
576FFnd/5cwpVa7gq9Wk1KazqHiyH4v2eU3Viqo0vwDytjnM7YmRkJGO8XLQ9Rny9NmiQrL7K74L
CrPAWbm+VAeLYYFKcyEyHptYw/MPgsAPV5M17vkIFDeeW/yqEPMb7KidZIlmsladj9iWA0TWvzbF
9RY84XQAruyxrlU4aXX98o6q6eTKOaYStZ77+cvFL2HENXbHNjSVSKCVgzpNTONaq0msiAjsdr23
hWhK+EBO7f8MdiOC/loMZ8x4HS9W2wATboCZ5uH3Sj4vC/So3Q9gX0arQBM/cDGDV4sP/rtjmxke
pF+ruE2MxfxVlndF6CJ5USOSjszFV2khyEcZRqJaDVwAMjwFBqwTqJzyH9fsg4AgWkhsPON9/ZK4
JPj6lGdu7hSt8/NOwWGgsKZ3DpOz3WhlvWeUAiodpjgLGODOW5FeTqHXEYjsJSUWMuIkvfH6Kya0
0SGsevoiJ6K1sim8F9TPKGXKo6OtUVH8aO5SwXjUnGAzxBLwF6dRXZ+666R1Ey1guFUC9WktKZUx
SGdkrQb72xabyEojrn65Lm0MrhdvT0YrQxQfeH/87l5c59bx5okLJhZClnhQGRngTeSmqiuGj7yy
Qgh+fAAEiY8SfpxQEGEe177RNXbpwRRlbo5rdOBrX2v4/0mQn8pi3L/NQNPwsxZhoaraB4TWCDLj
0xgoU7CHvniYqXY/tupMdIWwUc80WtX/iSITeZV81qHEFSv6oehkJtQN6qucxDzY+uH4F/0CPcDh
YSdqUnY6J51Clw7xz6XW1gYZ2leOAYX3faHIEy6iDqjwslCvNaHvzkrQKLVS5Q/WFGfOocy6WfQo
VKL3Mk4EKCWH7xW3UAWoRvMAH9/4x80gJvQo7tTaLx+GFkXXZXl62Iy0YIgg+GTJiioH44sbSC+r
x7KnTuU39qOvhfTnnxHjE9j3OJAvrcLeyRKlrYZkQzftj9LoUm5hyk0V7JVUEUAu/rFfQqsRnQjV
kJyIEPbWGZX8o/2gWOqoxxjiuKN0Qq6q7DHBjlRpWz7ti/gSKuw62UIUplIWgTwec44MSF993ZL+
Fzhz5VO9Wt5ID1hILXdW4RL6eEGDSWmb+AITUC4MjvYCOX6oxmfFlmcBUXvsMD4+hsGWFPJkQmmJ
QzQpV9z/k9NlhG4a8fxaELLBJlyo27XsOo2i0G+rzguV0rgQ4Bvm2Dy0UoVsi4v7rPv0ADJKdMto
H8tfDBSbrEOO8HhGMhXmWEDjf9DIEZw4scEIxDH/IffWs7OJzA3d59ao2ZKwXWROlHMOof/jDnad
BFzBL/p2x8Co2SEgKgregKaoC9Bbt8VHK2X6wKZww3OGadpxn473L4OPYxJNl9nB21H+nXimJyKp
TJS5cuBoI1ANBjOT3+KmqHSf+AIqIzUphrR6Dssi8f6M44ZvHYYL+dgGXlDfQNrtHYnncRVuy+G6
ZDz+0VFzWKnyVewX25MKoyrCeWG//DPAtutUmaShUL+vTi7ovHowKjPn1KWlARG4+SZoHkGJkWUe
sZud6c584Qt7+kZ8UXyYlO58BO3k8+PIDi37EES8bV5wExXuCR+apNFQxq5pf7G43imROk3YvHG5
17I9+s8zhCHdmFMIc0DJIfABKO++aPmLXr3DkCB7/BOeGcEid7L2dvEr4rAkzEAnPhY8yAp437vj
TS/oY/jrgSPeeYRDiI74NnWqbyqabYQHj9SWyC29TaiYbPs5ZkG+j7xA8SrqJ2kEjVIBv4Y34Xy2
az8x+ywB1TeMCShKiefvb9BZ+L524unzYn/xBxF0DlBFTktMznWxXrhdag05IoTgeST4ABS6kKis
TXeKkCaold6ufzCkA2vOitZHt+tyhLazjH7qqa8ymWb3sugCAXoxu9gPVUhm19D3GiN/kLi9sw0f
R3cfnaasgLEDjI5cyd+l3gXtRGzSwfgefcRO56R4ELUaM8XTkwayscqkhZrHWgy4Ev8ZTjLg8JqS
oyTyiiMD2RiqnfO1BT3pGy95h6JmXBN1YYuwXSFqph3+fHPeo0d1Yi+hunSWB5HJ/am08pEa0KOc
o1ys107T6X9Ph8s2c69AKJktnwoRStmDfCoxjNVW0DiGI9uookGDVOFmI8M/NryKigoGFZYZen3g
uyiQBP1pbiu6aRDgppk4zS/I8qCLWFVcvxI3jUcqU89/shuEXRxjcIZarN5XkF1JiYA5GHAezq74
O2YHr2NdPQMhN+vwHvJCsn/oHKGo3CLcH80mpFB4aYSu/zzhBjkerM9odFKBzELQ8EO20HGvKSQk
d9Mmf7NktHVM6L9oVrlbcQrMeIE5rwvx0PswqoC53AqQx+V6rnwscDZNXMwv6tgzxLqx8yysY9xL
7wiArNhhnbJ22vE68eqFh2OYlngdgOXEMo4cD/v6I3bsLBO5rLzMV8V6OXLjx1Y/KxfbRD1Vx2ts
I6rN4R4Xb27PdgfYdbLT9K2ScuHt9oQAkMOyM7O1l+r2odWmwkSR5ZRHcIhD8ixXwHROuRMrWfMu
y/YN9LM0dFQDOFBtr1By2/+g6M6PiupAqMKVT0SpM6L0qJ8l1iHvPSMXwC+FN5Zewap/rcgkRQqt
Yw92IdryiujwZGj7vyJP7PKZbgYIV80ehb78Q4crixA+c3AYX+RLKjvCGGQSZ0hfcJCFiLj3aK02
dzDPZpMKPRE3zq3GoiOL3IJIP0WOtnAzq+IPMB6gifuc72+6k6V/QeClI5teJWzFIJWzUoMUL9Qx
ACHrcCLh15ehFReP36ibQboEsHAXM4RNnfsKNKR/IBQfi9fcgNiSzpFmKbwTGi/kjFVwcr104/VT
4RjgGB3aQFQj23x28RGomJ1lpbYVeUZKiZMIu4mZ2qXzW1BqH7lOtJ37WuAEAra50GmJ+M9b3FSC
zRHhOi1eLLzfCl+b6+k4pUgqdiLyc301feI9RKbOqiipQnkgLWWr3S/HO3XT7hSqOZoGRQi363ac
SkOTcalLlJMBvxhcG0TiThE6iZ3WnGd+KWkbYE+ur5I96PsncJCtPn+I0qvb7PfJeD1b7TZCV+5h
JESCHv4UC8yUcnP9kWLqB2K7mj9yLV0LCHMQMxfZVryRIrFg3twlC65TUT4AjyIPvqUwlcOiY5+a
mue2OAK1Ny5qvahPa7VJPm1M2nQCJ+L/+NFLdK3gHUizwsRGel6DECcprGod2oQ7vN7u/l/WFj4A
YhYi9kydKbzRLjHJO82sTqU/ZBCZ2oZwEtZb0kkPoo/igjjoY+AWhFgjDU40Eq5pf7GSxPPF18da
G5EBkwEcr3hmtBsDZq0HFXhqWed95Zd+2lNIL81P1Zc37UB0Uc+m5rkIdnaobdhv5oJyyZhR2wan
qrAQCm/VoClj0LBtSPCl4LKJrGXYyfKPuF3h4pxH2r4xcyJARHSatc0EvJjDCYN/kus07z98Jsfp
cqLnZCd3ccc5Rz8Zcc6VF4cslSBuP0q/swTS7rTkubFFp3jXk9v5DKb6Q7DXmih3znrsJKXp0zRN
5sDVZVjYPTsKI7V0wD/3deU2Vk7OTNzLZSx2LY7LOyA2TCwgOkxP/H/VzdVgzNAQmMCMyOSKoBkT
mC+NY7L1zBTIZ6x3xlDQfSMJfymtBce2ekbNbOnurdlBmUqMGddGxV6us5/gRSq69lr0Ds8OV+cX
g4xOgKVPxEcE2RtN3hjI+Ji3fubO6KU0oPjMuHt46FGBwc4YYD1oyxaDYBwooLHXmaPaRHKmLJEe
giN/bobiQOX2U/8djeye3B4cs8KFiQQf6Xq5t5NUGsgSYD94QpdGjvHkltNdF6RVt1YcSYSbUdGl
D2+Op3DFJGAfjWAR8b79KqhQZ8eceuV6Mzd7o7YWLtPNSjGypvU3MSaJYUFJUebu/aPyxsiFhelC
RUwj3VOoKsGigSUUEvVhcL9PBZmkyR/myixobQl0JygGH3W+gLQH/lGZjbO8/oM1w5h0wkOWfuMH
GxMLAXksFHvjUV1zUzcv6q7j72G9bwZB0m6RRBZksVYvVf5HkHPg/cXchADmoUNQBTJVoXh9gANE
f0NW42nLgbwwJeUoti/LmfQTCjOhOTULiIRBAIwvhXEKAPQ/YiEeua30SUkXxbIIe1rMAtVpS5h2
HE9B37Tt/0N2jW61HlxX6VW/wyFVgZLpQih5EDFKGRzS3wPWyh1Anbldw1eNJCkk/gk0zsp7OBKy
bb+wqg2DiBPiyrHPX+cWt3NSS+LUff1KvUsH01Okk+9vEBaS//AaSdas0Joq83X4wtmg1sid+bjw
PlFUS6Ol7xvAD0cFJZtUhViKl2ubou0sqcyGr941M4Twg/Zx2rOclDX/8nyn3l7H+CtsGJych+C+
HaQAIH7Ifm358S+AMpvPSkn1k/7IcY332IZZzkWyf+hyucL0C1g4e8TjGP/ffAV2iT/MlCuN1v5a
e2DBD1yLvhIie8RxmSj9c45cxMGBAEjKTPdvRJmADPRtqI8T8s1rkRxr2Y2zSsVP9qpsoK9t+8PT
lx+/22okoWd1r5DOrnb/6rlGOLYwA+YCURGYmw59hZvbPJt33SH7QX7a37rLHsWrblZPBGOvKFw8
8Gp2c6clEx/xyQv2Sn0vGCwyz1jlTdLfJDH4C97I4/gs2sGvkG9k46FbwHsH47yb6f0tDBO06Eg1
Fj9QtBed4dOOwt6Q4h1EvASbkzHuuqlYxOU5rqnZHHE2YNKfDG6+mpFteaoQgWqA/D0hVsdCIQZ1
OxBJZ/LuUAN+HMnXw87DzGU1253qfYWkcIR+cG/NeUxfSOSAHxH/UUnJwj1XEzEiH64AMxwqk/jF
GJ9Ey1yKx4e6rc3PtEgPJCvK8mqOsbaGSOKShhoX3i1m5Av16NVJynHtGdT2nFMCIdH+3EWZFYs7
Wxd6ls1WRwyZQ0wYHIxweg5ekxD5j5BEeGvrxd1MfQYXPsg/lfmq7wXaUXmoxp1mrWRa/CJg8Hdz
vThjOBmDMyIQ6OEawlgY27kGybwfj1iDUptEzvOrX5r59pwkP8iRXs6nRG1JUwbONpEN7/+/3JXr
ocRrkSAGR4kBuRr27zoFx1q65GoR4RfX8BuGpJIQtp+EFZNwtkeMoQIQBBM6mHO/N8fpP2jnRB+o
4x9paKGL3WJYKLSCwlIWclitCkRNqEa2CJHB4SjoTtWEEzkR6JcggXxLyHYrssO0gY5aR0i/1xET
9TA0/ZWPXv8Dl9eN9LfaLF7SwEWCZ06dU14d7xkEzQHAU+bzBeL473SX/NbhsHvidzMj+YY9h7O4
cvpOdaPDf/QDZLDgMcABPYiKT8DgB+3wYFMG6/Y3zWA6m3dhXALk2+/xdpNaR/cTiYDWyzKjKKxq
tQeyFIPrZfye+8IqCQLdGx5uy31AffCSn/2bkDzjDNTV0hq5DlTzQKUSBPS2HpU0g4B2eRIveIv2
XDOaKA99qzfFEv5gg3ot02O6wQCYjIlxTTgzfSQi0OepbNliXnSPj6+iI/lPNRgqnipwKyp96Dzv
C52OwM9ScbBdERN187yONYLCyHM7eZm2KDOhWH/nyIZ+kYkssJo8UagXquCk3jU8m9RvclETBlBL
IlNnYWQlvx+3QhFDVcOO9/tR4ZstUIXWrR2bwgqSo8iCAOcfg1gg95SM63rJoCFo5gKG73qgKAB3
SZYq9HKCmQ3wGK/GbH7uB5r3oP7l5jelOsvGVKW3ZAou6SGMbU3rn1MI1zOI2loDhuieAbwmiB+6
oVphh04IwYyQAiJg7629cgddIvCJoKUVXLlAkkin1EBsCYMuHD8rJcH4SH2nM8j5SuIcqqxDqrEL
Lbf5Pb9Mp76IRmkYmm9zqa9byv5PkUO1q0+GsVNl7SUH8VotyXUq5gXbWlyPFySlu6hKA4uUDZdf
FOQ/g0uRQScm/2qn28G7ihLf+xZVQMXklxS8q7f8iahS/1rfTXKn3fxMxWfV+IihMJjknuFwfw3c
Bk+WUtiCisiFoln4BJ0MkcovQ1+yX3JCTDLud/zdaaZXuUU4vQM5Fh9RarllzI1YIq0SDJKoCmg0
dokMUCjkbLeQwjo6eWv39X547JNpyWr4w1hnVKrK9RHoH/Ec2P9B864p232xUlfWCcHq9lkaNwuZ
iV7EEwowKKBAY/6fG44WoZS4pDXphbs3K3W/WO+tKuoNocQxfD6pmootbYJqmvpzbpNKt9l+F6R+
VgE2OdoLO/0VS/cuGgPgtbjwwpghNafoJ7pioKVV3lCGo7sCJh6fYCqJ+pxHtcAe+mmbDrQZDqVT
3fOtx9NX1EEc5YNWzuWfvz+yK+Ptea9g3UsQI6BsezUaGcVpUilZHnO4dL2AMb4wRqDft4lqneXp
DQO25VcO+0aDec8n3gsEoR19iMWHgwBTZSDiaXYwpZVkYGNceq0Q7Mr6VSIeuHHZ6nFWRZbA+Y01
GLidjnNUeAGMyGwK4X7vRLTj41oAmy/lW9VdKRwzIXpTPLSn/wKNvqNj4QzuRigFcPQAbWScGM14
RqLfO19WK9Ifp5672VljiOaqVhm3YD+jVMP71SrvY4BdU/Et6GLjbvpnJvKkp3sIlWnKuMAJ5pDQ
XhE5vJNDEAquaoQj+okyd0qdpd9egektPra0L/DP+vGAq57umCOoQdCLybCPAxRrAc2wkWMhXHe7
5as7iHFHN0l+0/NGDt7dhqLpl7zl+ok7AL28HCmmMzSGMFHPudmZinm8FbiYC09OXwYds44NsDgl
U6isRJHShVbid4K73TgYCZ8DuPXIVZjB3K50VDCteu40AEWf1c7u1AjmIilPjd34s0GShp34CJ6c
jg2+aDWlmK33IvaZAjYgCxoPtUA6CZ2JU8zJsCBkcEXuxweXo3v4cO9HuioUEVDzyy2Gynl99YeV
313LUSHV8YJJO+c8MwNGLgLGXgVdTMNlSK+NW0KTKDZpMtK2xGUrdxY8IRvcSCtQVLnZBsICOLnc
i95MuhTq/MGN6sRbk0XcjkiK/25cX0wgbO1TirJHttgH85EL5RQHpZ7/qszk1tlA+SsPgtOsTnfM
oUfSypE5qN79ijduFKTjGZX5pVobLzSvpp5sD7fIp1f5jeCC7xCtIzJAwwE203l4/KlgzHYKd6bm
r8HDIOTL0GEBdnQPIOWcEeKssJnuuSrGUhq/77TiUXuS5PcjxbmZfppKCiAyV3tLSXgdWTwTwyzU
2fsbwl3sXyWI6f2zVzYwcJeUl9ViwhU+YFuNVEkhM4yI0VJkRQ6Xj7YmlesThmol4TtU0CB3lBP9
no3svkJJeOV2/F1FQvWn7p/XyA8Rzr0k5ro1Cv2y2qcsrsB1eqiIUFtxlm94NKqh4CgLsV2JtoAZ
GhqUOATUanSh3d04wkXr+rBC/PDmTss9amKcX5D2UVb+UyDDqOzrJGvr7rB+y7px6VaneuhXWtD2
EH0rPPM1khNj9PjYlMvH4KwHHWBmJ9ohx6AxSjRvslx6QK8Lo7DrWhvWer39Yd/1lImboOtyYyZa
MAUD9FIjEtprfuS+lRnPiprhNvAY4GcTC3VfkN4GqdGcI5QQhVPqM9hNIqxEfUPnV9fk03B2pBOS
klMZeCk9xIXJQuZkcEEBLrOx82s0vbR+xM5BIG+9mzczh+tLqtql+FQ21MaYT22hCH2hI7/KDfWB
jcN8yTW3Y+AI1OKKT2cQjWONvHLRmjc1NPqvCiNHDt+PwDQP6L9EVG5Kox8aRfMOXaaeG+N76wX5
rliciRsebjBouZUnJiSAcOEMzqwlE6/C3JqJI0L9EDt1J2aLhb35pYV8W8ulLy9QdwwM8Kj1E2EG
P+SPhcU7h9NnoZ+yA2NCqGpXGQNJeeckGDSnHycRiLyjmpO1ZlBcgBTAbsa9xzzAWVZCCjnqCmFA
CZGMgelQJde88+OAXd/KOWA2hn8ugaA0h44Jxzb8rc7Axpcexx8ve0l/fqJkJE2Jx/tOV+1yIiWb
pNwqtMXBE68dsGhnRPWU2HyX7d6gkTyAcES6sjOl1lA/ipJBO5sVvt9EPqLBEWax3NAp1uWJkCH7
POVhqye3RVhPTjrxziunWyZkDi00mhHej764zCnsctP0EQN71rNB2rwdbf9wNbSO1OdBnoyNBCU4
J2UZ7IOd0j3qmQNQ7lNZm2vRW5jlvRWLNMsSwIHWCWLHfkHx/6i2dLC37qKT7QfRo8UYUnaUkIrY
HJ8Ow+mz6BPJUy07E/t5irYJkGh4uejs+tbk6WqzW/sFFycXG6FvGI7hTRXMhkrtpnVFd9aHNoLP
TClooaVGOnxvLGkCXkP1tjd+H+daE5JXg+nF2lXC8oPy+TkUZUPUFeMjye8BJhiJJ5VM2dau4xsD
DJPqIlAZRKi8RgAr2P3yFiN0mLLGO033C8KJgaiJq62w9AwMPnG5qiKfUJspmTbTMuJlfrElSeHO
ilYNQIuVptHwpFRavO6XZt8IohIXw5mbGW5LdTa4slWVHX/wx8ptHupr1qM/twQApFEGVWWdWqmS
vqaR6V3gkyPqd5hvrmpMXKGOfF4OrQ7/huqPWicV7qUImJ9Mmf1lnNvRMfD6hJMEXaIJuAQZrnxC
H3RrzECet42PNqf+v4796EV54xrLI63YDW7EfyNXjwD5aAytjKxptbWa3Hg3LZpWfiBVo9yCqadc
WC1PRR9N4h3lYphVyTVGf8Ei4w2ePIiuMGfGt8iDcpdj/ES1a+cDOjd/mNqxN0X9xZOiBFhajsl8
9o8paNo6vw27jYuQvDE6g74xDym1IzIDn1mUJDyZTsadG0Ul/25pbwF6auiZUBqbJ9qo1PgWmcV5
b1TD/UlD1zUjnpX9oAgUQY/lpnf3QIF44aZYEmHBy1EAdOemsrqNmjdyQ2HgdkoOA/biwYPlA+Li
AdMVXKrx5q49wrwwSRI6C39KCiwrWbBO9PDKQ5JvhsITZ5YvsNehjY+7b89QV55yr4fvejkeBPdy
XlNS/qe6fY4yHQ1xeqokX7EXyKaLnNZV3rxfzi1EgJMhGvlAKtrqHseEcipsj4b5lDC+Db+MmYQt
dQxsjdFpOl2ixhaZOFn1+hQgtpJL3DPqKUTxtmiudU7CzjqConAdVolLRS6tSA5TOpgYaov1gnYV
Ml5gEYt/jI3CoPPbwfi7azPMH2yv60zC8p9O/7m+ZE53GfQLFgfbmIOD2BhUGfrVj0B4U/6AJ7Zr
krtk6DjLcUO+kUCnq4Hcpv5YToOU1aGQ0cNjZ/D25MNnNu22XyfU3ezPAI/LoSfSVPKwX8gQebGq
Zj+ecvubO1TGCI5PhQAWqElV+YUo7N9XrmppWNnzNPV46Luv5miTS3MBaCJzSo5ECtHtK5+eVreU
nVH2/F51AHhq+7b/3o7ct99d2y9t7Drm7Ew+jG/4lZAgGO5mtGsnFF54sLFVQOpG2R+fRDQBpQel
LTORfWH+rurtPhQDjjz+NKJIe8/gWyjO/yqH1Ubv5gx3HA9lIx4mNkwXzmiAUKPGSTY8F8BQb/Ou
LdPDG2WLQDcrroSMvCJQBxeo8RLJI4TBBYhHeYcdoRMfahxw4hdlpCZtnXtM157rQHFJRJtn+B6Y
LBwqNr4hs9JE6NrBswTfWbao9HgqMX0QNWFEXVurGQqKSxC9UC4AXJXotTxsEY5fM5rGSoXgQKlK
ZNKJJtJ9YlZFwsXALfKw9ZtHBAB4ETjU6M2lgWglKiCbdomM1jX6P2KfXTxxzcVM/ydaSFfSNqN7
VbTnguhqYcVyPg+H+x4zMQdCZpIlRflWsUKuMmm+W0a2vICIq5bFF6iDkTx3ukarVPBsTpFpEynG
3uzJVLqnSlbNMiBEmIKF8upbfqIdXBTCl4CdRQzrS3BSm1or+Nmt+y/8BfqRdXsUGTQN4dqMg2Bz
BI+aozYkeOjn/sW1nHRmKX27gm4hfEiKPpGjF/vlsonHufxYxAFD/iqXeKF51wb27kODn7BiaYbP
Med1FtcLhZ1L4GCOpNBSeFby7qnNUwJ/sLiXz3TCCBRFGrxmD2rUcm//GDgzRHDruWCEAgp+wZER
ViyqVgwMOjb5H7+4rRFuU8C6sNadf/XWkAS+AG4BDUuR3UgUgXDwmpOvu+OXoDyWGZGPss6VtSu7
Vg5oWcUVj4oav10PXo4Cf2pwA7I76eLSMqk8CqzPqSeiEs+2HF8Slgpp6YeCH1QFe1tlxOWZA6+h
d4EXQIaXLBdyVb84jIzTj0lZ6p2A5sZhjE91KcQWjTQPt3V3isrytwTm1tRMqi9wKxNF77V4TTXp
SNLdJnt1tUqNH9OmyBWJ3ggVF54FEkEpehn2b/mgLrzQonnKvyE8eUDOaz8UM7ZdxGpQ3szF7UYy
yYxwIOLAEGEru5nZh12oOd+UO7kugqZipA7X7EX35RsfbRuDB8M9+S89Pn2LUaNHnl6S+aGIhmcx
dHnk7cMYZvBp1GVb4Hf5xMkFJAnUQpW+MKNSMr6mave6KYMPPooGklM8KUILwcIja7t6gRvFLPMB
7EgcM7F7w2R/DUzsU78U95PxZOOnd6zR79YDcGwSkMhY1zLDxFSXSHwvjJnhEpt+jULuLgwUcIU4
zWnUkrdVJlQRnSGMNX/vjwUfxxUB9P9wtSsC/BSAIzoO9CI/HwP2dxo9TNakAvR7NS3C1EtdNxhm
EIliETkNcYG3o3ynfXoBJaX7m6uxWZCFDTC4imHncWDwuwRGZxinovOoMuBq9/3STgG7CYqsUcU0
T8QJD+R1QM2pN0WIwu6YJANeaPSSqxjmJUxxNJtxPPKP19AzUtLXbUMcwLWcViC48gmH69S6kW2x
EMmB/f4Y7aMRb8aG/A9tNh/SVlHK69z3tbxSUjPCwXK2ap+lmawBNI3mZhSim8XJO91+99rJk4q/
spbCbaCwQiYwpBs25RK42tNgjMwuSh6jlgtqmM/GMawuqS/5BYudOhbLscMD9WaKWsgWHzhHLpXt
ub0JYTevLcciIEiFoLlYIsdicI4TG6q+EZq31QMglUinL8qTwGZ0SIJ6n36LBv4KiswcxyUrHMPr
IWF7GBXfRDJm6tJyZDHPwXd/gGNh7mBkNp4A3HmbTO1pjKlxHYQ30CUZJAuQlaMQZHbz2v7Uki2V
zw1xPMrthqigRBBoag81UaV02ffDbedcUhULo/uE/L8rKSjkek9h5r9dJChARpIvIkmYEWoVDEB4
1uSk040QDarsu87J4JN0qHyEySRkuKel8N8jbLdBsC2eY8Yrz0leWaN8Q/cdxBgSJ2vWBlZ6x/y6
bWCX3k58BNizyUIEGS9sxwc3z2+j5S0LvGB8sxyaMKrzvqiqSrDj3GF8RNrIrT+iWAN22HqEC1U+
avHg8iVSpQ0GwB0fTluy0bxbFpV7sDd0PW27usimbN9afuB/kcRF4amPa09Md2c7eUv9NTSVvLf5
+GF0gYDqSZ+VEbCquSlh1F7RN0qxBi5zaonpJbWhbbRPFAkoqx93YgPwdy3nLpnFccYL8dc+AQwG
QPdFcXS9OdumbM4ENUjwpmhIsQlTTYbdV3SAO8ZRHcp/A7NLcut8pgtPF6tiUtlLMR89pesJkk+8
rYrChx0sLMQ5ToyrIL1X0kHb/wDKxp1/IWFaPYl/1AEPJqSAt6uaPK9rkOGfQSfqiK0Qh8l6vvfU
kIvlQX/0A5kykkOkufZVrXyXJ7JpTs253sRsIx22jpMuVrBOC4CxFls6h8bjnW3TxF9H+eAW0nMG
DFh4R01KXVc023WGqWpcIAFC+EGd9pCBAbDx2eNN2ed46ttxoERxEYpZyEV3GGosW8QjLHz7KNtj
2rqulNDult76K5imsD9ttBy6AmPNpV55LkNOjSN3TCCNPkGiVUHNiftdytdnGrCD1AwqY7SjZk0f
EfWhRXot/Fv9f0eWobonQTMtoM2LzI2QjdzHPewYroOF9db310pJ8OToubDB+051Qe9x/GReDMtG
LpJTwXCCvrepL6xoTTiO9VIaD4l4kZy4b8zlhN5jhl4Fj7Uulf2Ahquc1TJr2EkS8qMyYVJ45pgq
H3IJWXCfseL+ygsYNy9mef94t57DqDfCEVIrWOzD1mMZbFT+4kNX6mfoGTMB1JrdzQc0Xn+oY/RT
s7x1alfNwhFPb80Ro/sqqTDS2ltUrBFWipN6ujX3K4nWuWm2iLnCMCc7q5yJcTTDz3TRk9JfJWLC
YNpnz20pbL6BIR0i7hqu6hiU/JJOcGgjUNdiJr2JXOvhcM7jfax/ZhtkIjM1c+4myszAJgW+aKUh
h558sZAQWSk4zKhRRwtWbbboGrVZx3MN56t3LjwpCIRKVzrrmMaPS1QErydESPl5ANmBNi6kmyn1
KfoMtOM723yOtFpYx3liCS7s9aX+QneM38/L/BvJaXNLGm76bWxb1b8ZiFINl+tBvm2DZc1B/1OA
cl6C2Hm9l/3uOFdejgdlKdxhZTXSZvk6lwbxkWqbIJxS305qTAqschV1ktfVerMcdIF6/I4OnLUP
fLTRXQCvfm/c2aFf+pJw8YT3QUwhpNDg1uP7qRePZxMUcHbXMA2gGpp+0TRJ0TbKLpKGkM5E+L1C
XDZtHbP9vk4AIPN8+/aWTj3P3bgQh0zsF1YIJfe/+mCKpqSe/iF0zwXvmwS4IUpixQQaRvodCmEc
AJBpY0bkEH9JlIlDiAXSST7kRBE3WcT1ZYY3bfrw1Agld+dfPUx9vTAd5lCjPxThfb9blHZzekeM
lOK4FH2t5po+OahD67Rn20JZ1TMzaGvhtWZSutKeGkps3HPKRh8nR2dRD7noJ8NhS/jGN6pnc6Fs
uHrpH9356ey5bnaHChQ6D/Ys1wAUWVR5nEXgivhREha3wGJMxKT3bsom2VnYUWT7o4UOMoOhn4gy
G2DG5QpFneqKi+a3/i5/hmUM9PWAwA5AH3aCXB84m41O+V4qWKTXnkSgM44VY+U2aMVifaTC9wM8
6kmu+yLGAZH4T035Zl/vr0e4Yw7XmXezgTb8k3s563j2oBVeTUNWRBcqAo/pO2zuO0nH9yTNfKpP
gpM+tjOL3zSHcZ8+zdXqEdEa3BlfPQ0OxlG8qONKDodx1PI7LBFCALNAhk6ejfqYIDKcYknpxvFX
FRPxuKhEvnLUpaJIcF3YUGAq7NkmwOJ9nhW9fJgZM9+LYPJo7btTnXysM0b285wEWb/+1J2Wt1ww
WTPNBimp5Sl7Q6XUk/lRgeugouHuhCNxphE9F3Gd6RXUkHGp4clxci9rKAfYEQ/Jt64w59ebs7ja
bBQ9aOWeTtVboVEalv9NYdVKNU9ClKrV1ZQ/WebrsNjcFzhvEGFC15MdcBrhU7JE9WS9vXbXBOqe
veSKnih0PIP5mbxxavlqS4NWrw67wAV8aq0F5zu8OfOLmNrBjp3mHo33+N7tIaDbFtIw/0u4+dfm
ekoveNUzAUXH8lYoMWMTIX7sBOG12Xi9jS6opliNTC0DgSOoYdE9mvCX+Hjfrbx1OA/61UhJibb+
+t2lwzRQZEikHY58JewxK2vXi4esrPp1mdgP1te9SMrIMWfY4mrbSa5+L8XTTTGllj3QOoQxBD8S
b/ZKhqeay9i9V2TYHNBVy79g2VbQDfaHzrBaqRu9dvH36jc+0oiIcSE2pFeulUVkQSaVsQfedEAD
897HzQiJVTZo7h2J4tQOudJAVnEMr5vDbJ1Cwxwt92p5jPjMSorJAhuDY1j6f1TOvEDh/3Ym7tVd
u2pyweki6uC5U4fQQcrYY7zT6LOamf+e1ERXtsr9i4CtVKUxRyt6dRCDmfPA3AiRf1IAS3hI/Lyr
fU8dvG+mfG3yGoIAGCSpqPHGB5jpyTHnBwu9dugXfR+hiXVF/AkRgjRXtiOgtZuLx+JC9t8muKHF
87hwaE0c8EUzvQQgE8GTfsbQeKN+/pl1Kxdk+V5fY//NAOHMYmHAajSuMiY+U223Q657TkpFllYc
sF+9g0fwSGGjR9FUgs527FNO8ybd15lvnVWBkgXBAZll59BrNcIqxpcQVCiIlvu9ERF07d89UVoT
o3C01qL1GpMg6BH/dYNPSquINYEYHJwMS5WPtuBq1tIjh7fOkI3HQxF4bW++Lfc68Eq9vZ7/OmOd
LhcfQf0T1+WnYOeMKlGeHzGkfiv+JlCjJ7g4DSs87qKKH7UFNjP1JU9bApqZddhuusbHoDWrJfns
vvsbUXhOol5YpqRGQ9BN6J6KrXJ8fdiP5mn4ysNlzQ+6Y8Y0XzZvjsWlT2A3ySPfYBqk35kqSeyc
7kfuJ/0OpZixFE4n+73Zrw7tpCg+UnosJsOsfkh6fL+2du6MeXfKaW4EKSBve3PGP2t3XbFVpCUN
8Qlk2wPJHbzBBQJtymaJTiEOgFXECcul+0aBk89i2EQPm8fG/b/Ygw2i9TpvA32J9vI6tCiwUWzn
g9F+hM3tCjX0MWkHaHb8BkY+EcS9F83AFL/XQZ5btoWef+SygBnCw3NuUrn7B+1kTvesOIaA+Fpg
ye9yF33v89nnCHIlyUtjKukW+oTvvK4/MNAQf+Jn01CT8P8Ng9J/qBUcRPOMUjNuucMEV37+IXoO
ZQvmNqWep5Vc4hX/ZRschMEstjO0PVbkbKzXO2udPeJ5d5cpZqvsOYxWpMoW/tSQpVn9fIa5J70e
jLA2Ja8JsC33CxQtdaF6YiXpB4PIX5U0/B3RUrZX9ZgOi8mNT2/kLnZymh2+uhqmAqbdvyC9480C
mQ+gUrhQgHwyZMcNO68ycsxU7hjTLx4zXQuiaSbA6DQfnCMwBOLeXeNIsehsOQoTxrhPM57tCA31
BiMqbu3DuH7GqtGuS5Omtf0Hmt8ul905FR0pWea4TcG0mYtZuLqWeQg9ShY5qGV+XgpMLrIWjt2+
dE2oXxWv2MKeen3HdtHbxwV/9lph2cRSaSUe8yl6MeL5xCz0lVyfckr2munbGxfX6ktOkb0JQFiA
d+/fHRT/GURwHXmHRCK0GfKZzHBb63a8MLQAgWWVVfBtooGDKSKAt3Mu7U92WMVGs+2VHO6FI2Lp
j7dNDvrwjKuXoA/igNMOLhYKwWWa3Prd/SYd11BwIwPdr0+HSE/bIST8Exw9pBT5BFopdfPzmkAs
uiURW/sciRtQhFVV0cc9eHkF1uRYpwlPcqutn6EMxzzaDDu2dz2My31l0QACJWiNOzYbcwRntWIY
46MdhcH525E/3UNDPUp9rT1+LLaSBkr9q8osD+ztJZ9g/OgNRPpp68Wdq6hhPhFmB4sHTH/mMlWv
3eJs9todDzQtNovmj9nwmDpk//KuxpQO0+FQI9uTncpNCkhPcfj1hFWQAS+FK7aOMwtgjwYtVZDE
vj5yiZ3gZtwbuv+H75+xVQKpieq/zjYt8KAwRIEYENqfYusVKZiJF+s/BIhlIQCJYkj+am4Nc4Ql
nCl9NP+Q5IfypIZRj+Qd+rG/BLrJelNP+WI4x9xiiRIhXxaAYUgzcsyaRMidYDBEKZRbcPQrUruU
V78sEujEA/YjKzksORZ279KAfv7PiB/VFG3e4oaVbl0tFzt5mWzFdRF1t42bQHZSfVSrpKA1Tmfk
LSSeswTvH7qlbqzoz8C72rInAtTd+GhMVfSAQ0gnxLRq2FLa/ZL8HQytRcq1CyBiLQG18T1LO2NQ
7MPN200YufkG2zdhpA57SDzZhsDmanIJGnrctZOn5YUaurMPToEPV3Er0gr9AzrfiOoLUdqa9zRi
z/ZnlSWr3qJmF3AZP+hdT098ktYiY67Ew+uCfiHOHGQ1S1k5y9KKEZ8kZK3CK3psh3xhTZj7Gk+q
vnY0x7kB+irnMFUSfAdj6sqj86ryW+BWaybyckV5J/LoIqcEFB4NC4Tfq7/jz0rqqQtcSF0I/vnC
8qnvSzIRufUArvvfI6ZoSwwd66TtZ9HBNDQHYSllkL7K7HJwHVCVzaPG7zaXOiDepoHmL75Pmbn9
NuyDF+XyLaq9SilZ7lYHsHsiox7bkGpTGloIyGjoQWugxoEDT5N2LMX1X3rDPbUoacxXlT43lfaW
luGaSBViB4X0QLXoQPHyjVWeE/kjGq92zVr/yxuyP/NIAFsSlLmKLpjQT/JCp66qBy+CelmwotNq
SBxcRJwQLx4jWedMcplR0xDenYFP5p7NDH6I5WGFMvnMm9vM/JFPQFJKVcHDFBd4yrDZKZdUotM2
5fcP5JNFDa1naWSGRBhhkkOfQ0qQyJ1XhXt+K6lC9Y5UijMrQps7PjlkNeZKXI6OWO7KnVsAj9ye
LN4DIgVVzkEohqtstAMkbHW7iIe+wMcQcaHXj6Kb6nHvTbbE7Eu+CTrUA6/mO18az/5Wvs3x5i7O
CxpV7LepD8sYUKEsSzHDZUkAPIRixrHZ9Led7+tb09+k7ArUNTCFYWUNd0Hfz6hj0Dyday7yuelT
mz6JUJW55qsYXOqZbgdN5WDEvEqSi+Kz5qiqEGau9A+T3ic5q6JA6YZG1PJFJjzcIpsDvJcL1Pjr
SDFRozojLMdW6jQzpizcZOIhRdTaZsd+XpZ4uPHnGE15guz7n53hx8GYRMwD1KBE4JvXvJ7WxmpJ
GCN9CeHaidCOwCrAEz619GzUkAj1H0+Zz/A7j88zJaXbg8z9wzVggEwtIQyt4nKCue3N53f0D/Ea
LdDTxVpZunj/GqIGyRucCrEHtnks3fS8dr+pXV1PTlyHCYt0Qm4X07iJYhmmkJuEX/9qYggHLjK6
koclVNlJA9IVS3KhZz+bw7YYiGhUWO7Cb2seiScYmjVIZLcrN1SUpEn0/I/cvMw62SWvMrmRJOOz
1NFMA2Fl9dApHXetIG/vUXMvcUAzO2C71lFnUrvkfU2BcayS0uy2rI+xejSvZx6THtnvxeFTJOt8
BafEddFCz2YpC9bFaEXhBIt/vCRbkyeKgeLtZ6MHzMtozme0nRcqniFnwFOsjRxNLRXQSnDJTDd6
vB2hWggS0Dswg+8IoJwrBo7b/Bh8VJ7s8sdydsvYnSwzj9bmkrj/aWp5EPDM47G7ILZrGmU4XwVE
D3/ZYWqzCq7QYvNgqK9A13ZNzx7fFcd2pzlDVNzzK6ed7fC5KtnBjZvl0n06D1HxzHKPBm9Tq1yu
1a0fAeKrbi6JWwCgwv1UDk2v5sq11GrfIHq2igyerW4qhMFQy+dIdhFDLBqeTpUqvJsEVWRIuC4R
sMxvjKyk5elM5WXwZBLykmemB+BdeEhSMFVXnn9jz3kAck/W/sQxjiZwNn/bY0bkfZbC66o+GqRW
povNMOuVFA4an2FrD5fr0OMhXhj/z/5qgCXQP8CgMlwXFcYCmSBRearxkT36+CxpYJoGgR0FDnCe
hmeRs67ejQsRqnYobG2qwqbo4B4wnu1M3TwFW8JuHtGuC+aV1DK2VwXhjvGeZhqCn6DXvPMuF6xW
uTFDdbLMVp2HPGAg7lJpnoqtiuqBR2eJyPo3dZDEB3eUMydg7ibOH0JTXWp03w848OIg6EMjfLnt
bF6LCjg/Y+1sUPOb3SOCCKJdwQaZUKnNThjUJkwS5enig+kzTC+rIoj4G/0Cr6esngLjGlIcBO1l
YEqxZYijHEUSz5wSEF65OGp9CgaV+1iPniY5fE8jZARABzWW+CsyZ3D8a/zrPmWy1+2h0+wQt0E7
2avjmjGvyT2+mI1pE35QkF+PiwfNQm6iMdWkgJZn9bcxdbhTYQiDO+4xF6Ovg1xHSU86s3bpRi5k
qjxcwLcoMVM32Uhz3rTovPcpHfHz5Gf8v9ADioDCupFuOrS6CCMJlCFl4BxRZxjcg6/cWSJyKVAV
2x/dBVp5F4UsphaxOZRz6O+wu5lLmyGVlgEO5hSG2wg+3czTXT79GV2IuTV+fKa3IX0yAi3g+3OH
50LU902+MXf/ikOM4/opuHRzKSgAMWlg/lqWPf/+GCicqHv8DnguWtex2tUwAGYL27zByubEUdI7
ycqwYpGDoxCWHSvjMskZ0SN60rdMSo3Ce6QfzotwdbuPMTj+CADSMqYX2Kk1Q0ws1vejQDkVFDco
5Iyj4G6mIYD9b5S3Zw20D5xr+2uPKVSFWc6c+hfwCr6yPQCPkB3NGhUc56phA3dHPoBlhBJqD2y/
FJeDZ4Zm4tP8tdUh9KKEIIsLzTVCcYJQNXyZAYtZ9gzEWP/pN9SYCUIqMGpXgw9k7Co+VT2jzox4
fdoGbojSYrbRPT5NetWrTrBLk21BuvaA3El6i7o/mARF5FhB4Ya89tZO0b7AKni8MxPu6TzdnCBf
NVOdnIq7EPfxbQH1EN5J1Skz2A8yt3/RlJLC/vw9HS1x5acqvbtTEb3kmPKg5qsQetyTDgGtIg+c
XP7xf1olzSt6O6E316JQ3VvyzhzvPBZB63XY0KJj/O94b+ixgdCqAgBCM9OcHPV0ZaSiL/xS+Lhw
A1/obNCSvGMwWRBi1db7tgyqF1avfallt2r/volztnx6Vx63X6+z85SkvGCxv1aqDaFdjwwtOGv/
8nFEfPo+FJfWhrJO2Za3Gn6rFpKQRktfizPQEpzg6etX/a900Uz5gAr9YROJYSOCQtLZmcLMYewR
hgwEGEr+Bv6qxNxiO0UrvtXaqEHHEI3J2G0qQfAKJRu80qxLXxaUJF8q1BTiJIXDQppGUfmSNjvi
NNktMoYDtY9Q8T1yo2WB6aUT+xP6UJpM1Rx3EL2QgKbSwrR2oM6qQXqNbmn/bgXhwuRHYMdeWLX/
kIw4xsx/rlLI38vWiDvcilanOKE7lX9IeazpTgBs2aWgyox5uNS6E28NuXusUAsgzYZJQ6OsFZyn
WBzEw4QloMsjIn7zjj1dNG4Uf62rZ8dkhONf0FKo8LRaMzi5XgMhm46mjC79MMORBmsrAzBrko9u
osAEdQArr37UGxcOZPlHMOOUW2MvM03sjX3O4ngL6nwuLMsqWK4idQ1sAzP/fWCK9jx1ebPiDTKx
1mx0/MBh8WQ4YOYIMZYwQEnStIcKSwhaApy/2K3fM2M04Zh9wdvz2Rzuz35ZZRPBWgRhewPwJWnp
YhmbFP76il37E0lcRTL55oKJO8qJ9+5YYdmVUpMahB42I3F8C6XlfAifexii3XULWfyvlliYu+ai
1GZ0yGJyKRp0FDYdqt83Ya17N67ax23IF19SpfwHQFer1uK2j2WuxpVGsu3CiGS6eCkuuxQWzpoZ
GOKLstSC9LerfyX4DPG1VGZu+vIME1HotLTEfwlHLY2o5KHuqcnpVGkNX7uKbr1f1Fc6l4ojPb8X
7Q47B/THD4cJyAQUx/oQEqUScKJOEbatUvU6vVPFa18mtchvAqC5YHD6SGXKE+jGedrLfo0P7BWg
fPpxyiFDAXm7BpEUlyHqFoLhcN0fowsgYtRC56C0wMGqVC9oWmzo6+MEZZgn02ZlzPFqjiHCmo2V
nXuAPTgNB38U162zku7+lLJzCrygsopWNCuCamufRt8BPJXkjNuuhw39lQMHWwpUssKT2Ncp8p2I
4SrE0J77Xf+MgDcDz2BNGBarHFsDhDSlhducPRKx09Jk/fZ71sayVdECvBqrVW3pPn7H4lsvTgkW
9XbZyeW7vUzjRGB0dvmYA5dZHIpHvtEna5Yuf3PjgCgYa5eY4eTjWGPznFuz/OMCOmFN39Ay5362
5yAZP/KFy5vHxOBPX5fjnbdzLCZcB0oNab9Mg+NJbtgLZ9LpXCQrICqKNp3eBsnLR6qTJYHwjovU
e7CvDjWhCHZzIhspBA68YtR5OGqolQf8nvBjhUSSq3yITL6PcjgJ4/vqyrqTGgMqBGy+O5KV+Wo7
+fzrDz/KZiV/bn3a+mcH+077t75HBefx/rLVDXlPBhk0yWp9r4XlFDYfIHZiyHullwZDDiQ/WMzg
kcht/JLzSEYKQKR5wGpR4sQUf7GGK+751AI6KQWqohaySmxmgbMcpjrZ3vgQ2VdaY3IOgT7BQHjf
eQMpPPbnPxUhqOhfSNKN5y8bAoQBC6986gkwDBVJ1+p95GgwC/yrHjejTwCbPRqeIkOzfpkGF3Ho
1nVf0oPB0lZw4pYOUwSSHSnA7ITrpuZbbTgZYamB242z+t4yeMbzDjDU2x347Ip7jLh/1FOigQox
qscMceToko11PDzGGi7wjwVNvAv35DVeFaJeoGM/s2fCPvlM/QQ8MjXusPF5YotKVlnef1pP3Vpv
k+JPDRX5b1zMfysAdas+kTI2jlKEaqB5gj7/ROb41hTFyLMOUCumbLdaA3KGFMfyDDv1ek8y4Po7
X9Dc2vQ5Ce7RP3jbdAv/Pe4Vx+AnZz2Vb7WlvzHfRp4EMxJBMsGMI+9visfAq2ikyf4lXmDzNEmL
pyoN5XKhRaZx/Sh1SzzIPg9pdl7dH2eLQhu1GL22Pp7NtNsW27hE3f+wS8OUrHPjjQhNCZp5J+ZX
JFGaNTnsOxIr05kT0TUb+arLfbjizL0moXyVA2FRSNnu25Cxtp38ov3QmZ6nVDHTuZdDW0HC6ZOB
udzvBhRhrcVie63zuHLq41oRBgNtTyGzr66f8jp27aCE7cXhtJ3zBj9Qui/TW55aTvtl7fPB9f2X
T4QEP/2ZA0M2+1jfjk1w7Hvx85kTpT7m/7yRV9jHE1O4Q8RWBo65oeSBdWlyoc+EoB/9j1a3aeEh
39cae6dLKwyd4Ql2XbLdsWifx5+P/b+koAosIRPEYAxl7BgKbvgv8yxFCxuRRyU/eS7LVj0hJC/x
yQlrYW0e1G7Sc2qP8zSMMo2lhtNFTWSRPF0Qq1ZAS00tlRbn005xlJfcQedA8Y1qjNGgjQaJbSgP
YLQ410CQAxIp9R8ktIkHEW/5BRiXj4edtY9wd/85PeBTZadjB0Y65LWFjLP1hJ72u4KKi6xIA6mE
WDQx0rsd4ISkHfucxp83xCE0T5/cSFsjU74MWZrTvG5zns2BkevR/OUwmTTLm8WQZsvgwI7CE7rd
zqzOvIid9rb0tE0rjaPZVUFIBKawYf46suZvYfIowepB/QSuJ0HRolOUdhZbPk4QPAQKkORyrtHX
uu9+rPMwjgIduplHOZjfR1k8HvDQSIXMpNvvEgOzoqjVaTmkuQVIQmGmNxmLL9ZKMuOIwqNf62o3
YP2heRZ9JUlSpdmsEEZqcIfcHFvMBvhuoIDcixy82odH5DAs3uYtvgrMl2zfWZ3vQppGkG4udhXo
3TtXvFsJRDR9/XK5rNS4XijqkeQEnAmJqDYJwuGhFgIhZ/aeRfCyS+A758KEq+ZMkSZhyS4FQgt2
EwyQilHYR4yuvlxV7PAcUo5ElBM7Nj1IJiBY06IOBWaKhjnSi+GmTmcY0yfNhj3tKop0tDR6uND8
kyw+Sm/vJjBPiWRHemmONix1vo6HtEFHNrHmWvwyuhCarEcsCwtSUrPbBnVl3vQeo4aZdyfahune
D0ZZrxJ5lmkQe6EABL8C0ox/mZqOQOqrdU2F6uf14gjG4s6Zl1wz81r18NETEcFNLuI+rxgjety/
+wojFavpRhHBdKeLn3bWUxp9JetvQy+ro2v8geenk5TNNvbB/KzHaWdzXqG6q4+sdbMLhB4fnKpT
uax5GqVV3zD4vIWEBlI/4AmICI/r3ag+O8Xsuie2NrVveatzLXjvUm+CpXoiD7rTNmO/A8Dc6wJ4
uadAuMd+K8KXm5KunSrmT9PGaZm6NMXCfhKz0a8rvD6jreLuwAgXCNdC1MPWrRuHoE0DbdM8d+Tv
ltqpLUZZIeOG2n04GFYnny3nquEu0Nb0l6bPelbxXH9ELsnmHv1++oMGqNJJjOcfTcR3wjU4LOuf
TLpNGEKStSp+JUQOYHZyjhMNm4zZo65WsSpXh4Oj+evR5qW/4fXVjrR5BU0ZyjFUNi3HMCuoG4pu
xuS+2WMyfpt7t34sI2VrD6AjUS0BoA6U950Sq3zabgRHFP02vfJQbpsOJMXT/9WMTtL4T2TgExH3
6c6jOR3OG6NU3LzuE7uTBW8MNd12wiyN+bZARnVdLQsmUBxDbjEPWsCNyvfss+PGC61lU3ga2BCS
yTVzR1qYg/zmfiTnO/ZAYnhugB5e3glWW/h3IkNlXv2G0n8qbFyUsNRhwhLApm1E/SGeNiJItX+Z
r2ewJpQrLpVUh+ASaifaDbxgf8/LVflgProAUXneTlm4Oft9rkUabh5poixSGm7Fw1iQACJ/PirD
PlMa3AEulNdvxDk4mVdj4YjB3pibgs6yCqRjd3Y+7/blousX9c1huTwnp9nrAFrGMTH3cVKLFvZ7
TpPNhbf9k731riMLize5SWaiQf9jVKYVhIWfJw6iLZ3N7ajMKVc0pqgyG31aHnJZ96Bb+fu+uqRW
uxVzDw9GoF7lENzxluW59Ea6LMUwdwU0F8/m50OyEBFgU1IBtba8C7IK4C8xx1VVHyU5k8wqDsLJ
5PvF2/BVzS0LXmxMukLlTuFGnpsOlVN0ECEoVQ//APcrrqs6Y5m9/CxeQCzjCrBC/sdA8qt4VbNV
fhehPNsySXAV3Ezb6AYT2YBVoaBmHU8R3gXhYtdZDVjkOIZLKclIKZHBcZ/rSsqwLEH76iRuIUEy
v4JImfbNFPBa3EEVLY/H5ZyrHOk3lHeIH6H6psxsxpRGjXc0NSm2ICsznEeAwRgYM0cphbjkLt+2
2i+ZzwJXX3kFL7Fa1yaNUXbyFhma0trDz20i8VRxnKvYSP6ijJz8jwA0dPAHnhzy6pWJJLo30e4A
ABnvKeNfrCR/ZTg/02DCE7rEIi66RPNhfOs3TnNa7WzITX5Gyva74bhU5gTzoYqua4+uiYzVpagd
4kJPGhvVblJqliXtQTu8/h6ggp9JTDUJCJENY/zRiBRjp+34KzZKGmOEcvqBBv0dvASXx2sMXtOW
6atsFaVcebhlUgt1qGEfXZ6/VJjVW3Z4P2YK4Oe+oYoeXRhkUSTP/NPg8phZz14BcczgP0M3dELj
qlkcH8fBWVmI8ZbLtakfHyVFtbQsmP0gVobulAEr62R4NYdWDj8CV3lCqX26YS4VnVRzIbFT/P2Q
ogY3lCNyNBKRIXQJm3nqHPKUWMKMSa1LdDMdLopfX/Kh/wJm4x4sK0fk/pScbqNh10zs8RGoqCpm
n85dEHapi7erb8qn/V9X89Et2L4s6E6c7HQie2GcWWf/gqGAapwFtRuXGvYtTEZ4FYZCdIz+J8j7
NBFcDr+vteVlUkE2Zow6Ww4KGoZ8YDg9+Nhd2UkS8jQoz4d4PU5/1El562iNt8RwF7p8Wjne04YS
wOQpFL5/jFnToC32gSLyUllSFpKVOTnBJOoK4ONCyV5iMwjhtpZDfgLTW9pMTxFW8JOXEgoA6r1/
2H4tto8aKo2LLMk54GYGrHUvNoIHHDmFUnklqCMsTPwMBJAw/vIn4bMH9uCvGWP4LXEU0XmZndSb
G0T9i5i5X2jzVBIqStlbOj9e9NMLahhvvMiFrjYlx5oDqkktTxyx1fzsvZ4G7ThsHHfyXZA3jqo/
tLsfHeVgbyfyYa17YKLP6YkzMyoB0Id4XRKKT3yhFj1FilUZEOP+EAhFJYpFAjo2grR+FyrUKN+g
HFeLkTcBHUK5a+pL5XomJX6YvwrXB/w3to4oWvci4HdRlfR3Go4qabbmSZS//+Tg8wEGDwx2yCzt
wFvoCwKMswmPosTItzExQhqQtLRGCzYYWsstSlguD8JYDrepWuD13FV1nn6Cgt/Y4uUJ63RDZ2Ht
Rn2hjkyXyRrylzHYkoLCOCxQN/RLskjqONOsUtJNhamQDW0/38TQ4h8HuahmQUww5gOJnl9GWRxT
dCb4asJArG9372rqHM5/f0vPo1a7TSXHLLlYSUInZJr1tcJZq+rXa7wMg3oIIf8Dui586XMxuuC3
3HXQVovssqdSvvopmBaD67b3HTEcoZP5C2qu07c0MYMhtEiGHdu9jHmtoj4oN3UgzKMvjYgK1Xc9
e2zBlSLcqSzlCuWLlW/4iOo7beF9zuZbfF6QR5Imdth4iY+qSRgYWepkIHOsfJ5WJDB12LX2FqmD
h6UvX4eNj5lKBlELBhAeJfs1Jyr4I3VV41ZbK654fC8qz3XbXWcNUa05JkkxfNQcYbBWbdhkblMd
AMzAKO1mGrWKcCs0UxlOqb5d3pM61+ut5oU81U8eIIxbelycvdaVokWZqC8r9UqwfEXKSC+zxw0V
TPG6aAXiEsIYBb7WFQzRvjFdA5IOfg7Arf73nAYKVeDDgZxGXGlhH2qfqd1Glk8JWnl51ajkh1Cu
wFzBCwImxigQYSfD/kNIIyt/uAqIDuBepOs+s8kuGQecSJgT+WuAW3aZRVWye36FlqiAfcoK3kLc
zeJCSYbWik3ONwCmsvSlz0+OlVcvy95ExuuGgZyOg7ZvQ9YkqfDYlzcO7xVsxbGtNHXcLY4C7hd+
94V8BNk9lG0d32wRNFAJZf8uyErKQmR8BsYWOoZX51m4Yc5JxQKrNjiLcpkqS7utHocawwRrI2HC
SLjMtoytPU/LyZ9AmWavpYdZBQEWCOHmxy31bjPpnQ0q/GmvFl4boSjb/COgrKsm6HoKWmElauPR
SnWOEV76xRvc6KLEecUids2rMFzsi/njBr5ZU1mWGiwgx+vuPuWNXyiu34V1wvvWqOPGZjiAN5KW
VdCSx2AgbUGO1x4puYUlNnAvALntQpqbVoU+BmtGVVoD66K96b1sJq6govLF1joQ1+RdJY9zLFmR
VCqtixLJXm0CRAMSYlbgkh8AInVdqCCkdGXkRLlYqudYDN2T9kjbe1VooJrUbnqGqSKRXL68aCnQ
SsYSP5/PBAByVs2FhUo9K9UWv6adl+y4mgRwCnXZ3xBOHv2iYIJIq9JjNLE9os24S+eTxCxTKfSE
Z9Lz5YgQ2WPYlexlsliiur+VmMOKbECLg4mHSxFXOCYxdTZtd3Q9MoeIcugdNZw2TQ+Nylmz8Zda
MP1U1Q+VdlPd+TRV534YBNmNgaI29asnSLXOHyyk+qh4CnquCLc+MBorsY8EGCynFm7TR83PyO0I
+9KXghcxzz4oz9Ud+nktJTt2fBRcEOqurOeBhhdH0Rbo2CSGbFZwonBfMq5hgN2xAgpzN6sPSSG7
ziGlZmsgC+3YHrs+01a6Z2KqoZNNiF7PGpEuIYgK7DyQM61pmJj8x/2z7sjscSAUfdrZ1+xsPyvo
aqBDLzDzn822TeV0sC5A4r2k5j8uKkjjo9WbER9ohrBlzLSgBdJyW7M83RnE7q9zG2OzWb9vMmRb
NDg1Y4DigmbZRV0U9aB9vKftuDg/gjrhwv6e40CzU0JROmCJNdzGb4wZKkvT3C6ji+VS+oV8T8Qm
LOp4QPnJtIgL0rpmjtY3WdROOaTShj60MRQjvwwfFJZX0lR4QVt/HecfcWWu+3NJIONLKJK3339Q
YaD0eGzhi4RvFtQTt/U6wq5Th7hIk5SwK4xIN75w0IT1arUEAYoPOuFLnMh5GsNrGvWWwLknoECh
zCy/oa/sIKkuDzxWXJcFbz75oT31h9tcyAWNKvWvKXRUy7/KmlxHNsHRvJSV5ZLmUzTJsgPsPWKT
csft2mtnrLlfhR9FlLOaY34rR+yb//REkBFbf6BPrHomqZPirlcB6m7U0L5OOnIl+1/3fnljtLPa
DMJSP8G0lHaym31Hns0nQCt2dCBiFrFTcDLp+4wCtS9cmEZfHF0cmyHVXNzCQ0gKcFJHXShe1/9r
xzvkjmROu36yirNXjMexWhmprLBYwuaT8H01iq9wcVvIWirp4UP7MCcCsuEkGs4sDMSrdWt2pSmG
z03LURFnFO8kVwmxbffMGUPblFpvvKamlklIhDOnDDtPB9UDUGMPzbJkNBiXQ7b0mksY9kzWqqJf
dEHytOvxMuSjBFWiE9g86keza4uvFgz20iP32qGXiUbk+TJLp020vq3W9/+lIgyiSxfiZ+aTxQCm
uTucTYpousoXi/RZBB4ntzi+Uln6fJNhbl/777/gzFfsMohRojSsOQGnraXfzt6WWVE73byxHeTT
zQX7V7ffPgPiMWh6dz3AKfsYJphsYc169Hf2hRGpnCpG2Zj1DTDxYtySDFgaJclF1mMvf+sroS+q
oH7npiZfrC00BronhT/GZNkuLrnLBA/zWiPEWcz7GbBP8wza3VvM8PHqYPJACjtCcAcjXNw4wbIu
pmFOC74vmVBzndJFuRTJ5qmjYhEsvYaHP87JkTtD5+XxtVQwau3WOW6IpOeC96dVreU6RK3K9rp0
uICZOYaDbACjcl/4dHofJdEXHa9+lZvAmcqkq9p1/PrlUuGXNrFI6zLgdLGTQxokVPeyyoUt/Hbp
1nM+GI1WnzeLdb0AcmSvHqBIwTTNNjPdjIzDQDEd6cx1ET7ZBKWqSdo2HIyVstLTkJd/f4Iq2UtH
hpYYZQaHUNyVukFNmS7I5LIjErQU0aCdoOVoML9M9EcNu5evRckLxatBYeICoizQWz1VOsSrX1Yd
ovKFVmvG3a1QrAUiY86MNzgSGzJUsE1V3kXLxoTBIyzCTuUwSv1bxfnKLH07Pd0z9jse0eUBg6mR
j7MDgaUDNwGfsjE3tsCjsqvkNwycSUUlsr6JDxp3ib3biDCddi/GPbgza74ophEm2wRwNY5Wf+We
5HHiJq6C+a+OLmiTp5ZFhL/En1hbmuZqVj1cAZpNcLqDbju9TOC2OUO+qF8vxxewPB5kvNi5aDsu
1obn/9vuv7yhitX12sNX5sEAklkXqfSEZYohn57/cAGyOFnL7xYj38SbR6VDnYYJv/nTfEesojkR
FbT0dJNmiYMMl2DPlTvru66a+rNJvRHBrJTMxex7fohaaGUZqKiqBoipf1HZ5D8ke7Q3tj0JQehB
quUY+5zIDL7shu/6hMrwLdqablWF0/rQmbojplszyBdprbyP/ncCNWZbYxEeS47TC7iNkjNzwmL9
FBp+S1oeclYbUeUd1YG1KgwWJEdRjqD3ZuwsWWOgxE7teA0qckBiJqisjjVtimTJWQw5tRKMHLH4
//YD6qy8hQACdkbd9SewEA1UC2UspU89+osLKBx1XXWffaybNVmKHA6q66jNDf3Cd506ih6JQ8QI
StKqGhmrg+KdC0RqAeEl3me24XGGDFbtaUSjpXaoI1khkuHKF6yegICmQsLZ5bzARVYFaHxHxfMu
+Dn97S/7mV4vZsjQs6ySJglumevnz5ob5Ky64KbnnCDPq4zDe0rJJAfBG56XDPhBQNcXeCTyCWIx
LfF7NnGEKyv/Cu52g6ACH/Rq2+4mOVkUKwGJ/y7sXHoxkDW04lj0YiOi2jHVaG3bANPqOLEkWkFb
TXd1s55ZMslGaWcEpcQXNrmPGEyDJ3B3BNQzL9EXHOshq/4+5gQUZ3CjlvYWRax47/dT+ZcZ5uli
h2XIbTXrxAfy3mfO5e0roys9CkvczaOLyk+/ynjQkEY0ZXCiiQuKfUl+kctMAxOQnoVqTh5RoiRj
A41GF1ZnR8Evb6dCfCo6s8ItO7hpsNN8Tethm7UWgSX6cOIZkINeNDPfiPeY/j2gwCRZEJHEvmKj
QSTR34BBl1AAe9/7NP2fM/pQzBcmQhToZVmOyrcTWOP6CNWwCDskqxy8tvkVehbkUP5ads7Xddq0
dpTsF0xM5JeetPJdV5DdXRPDfdMQ3o+dVX6ZdlvvXaIJjk9hpc13VL4T1VnuWwEaNJGEi7n4vspy
9R7CLBcp6bJnJZshenJhiPZcJMiu6OHX/1a8l7WCKwc8CdAY+7VLWf2a8tOuWIE/q+RW8CX7A/aB
cBTyk5nM1R2RmDz6+YyQ2VX31ydFeIopRkEycF5p8GWgSaP3ORY1Q0iQGFZW6jS4Wx+Vug5cPCpZ
DENs1CBJH55ebV/d8yvJTyFeVgEnsKCpEo79Os+Fwr/XokE4IRVlTKAeL/NR/r+5norB3y5PYNPm
CC7S25VxKOVRVdqWdWhFZJnN5ccLSfWi++5BqOD5rcj9qDmGdzSdV9lL/2YfqrSz7PfmDdu817Nt
IQzBir6UNpDoJ3sb3F4w/rTYVp/KGwPkr7LMnmBoj4KpBMPk5gvntsSTVZrOMpJGr4QJ3PJVAyS2
uczwo1+ptLtDn46RoJhHiQ1NlzBMJUe0fD/YHwiz3oaqTfz7lmLV1kRsO/Tv9aAYSD5IbnMTjNqN
C2ZBZ6itT0yJOQg5xxHyS9IIsSXQzwK61FlRTnQvQ+F2fSPjmqpE3OM7LT2EDqnWqHTONLBCEGMJ
LIgAbYm/HzQs/gUQkd5UObKbXB5Ho+ADkdYyWvNdT47XiPVTmkmGKQgWNFe7W0/Da7m5NJDyjCpD
5TuzJ7cu75KS71C94N5JGce/3W+mHN0zFQnzvQ59BDlF4ei15KghbkjB9ZWAB43KBSWNOD4QBNjD
+LIkazBqPsEr81Po2KdH0VJIILWJaFtqdtrVKajOaQa/2U0M2/2vLLxCk0dH6aesF1hJqEevUyxK
O4B8rTAPKe+M06sbyl6/tiKWyXzd+uAkaSbCK9JPo6Cnex7pYkd/RaZz6dInRh209MAMrQoqqE0g
T/yztP56Nks2JDVU3htOF9yJzMO3pzpEbi8supfjJ1psdJUVweCg8rw+oNi8Jyg00QM7C8oGa0lM
2hTgPD5jC7Jn6ioW2qiqSEfiVoe46DRxlw7zo4++zkczsNyPjAlGLdGqgk2yYjNZ7yeRbeR9NCyX
Cykrqe7i+3XIl5dKvVWDzTMsvFwnbajAZX1PKxOwtlQuuvoB9EqE6Ac9Sh18lTejNHEgsM1laj51
MbcVjwkTcpQzH46LbF1KL90wLuozOaowznYItf8pe2sCqX+UZC/RVa5WdlpVnUPQ4UFbWZ4wmBdY
4hwW3DVaiWFnxrHHQA9M1wqO4n8iwA8mxD8swrNQ85GCiInj3zcFobuKnB7ok0krCT9oraR4fdSn
S4YahKgoMekBraD8iCgC3cQ5Oq4KO2mA9urGbj62qhKUgLzsHGa3w7wH8SmeB1ygHlxRfbihJl4t
PFQMhCcU21LJAjyx2HP1bXz/e1Iqp/4ZXYLPi2cSnwhqqwODkf+Qq6koj1YrX/cPPVplKChg7Qs1
LeLz0i3Cq+AszUFLPPZ8FdCnrCSqpo9i5MByusbclJKlqMtwthnjjrcXSbGMj93JS1RFLosW0zLl
LTNAKrDVbWD4ifova0fcjODbLhAe2V2YWj9mVylpD/VCvScNcp0C/lGYKFTHlbORxB1P+8X750XX
6DJ5Fi/fTu7LimDZmQ89+pcn2pvpcIFDXGMdc1HXh40gb8XkFcbdZJ3zzyhOO4qTPJvvGTJ1fxQX
R+wZ/cfuAHybVN1RuCPmCoQ9sc+8XpRPxCtKh5bf/Yo2DLXC5vxz08umAMhY7fotpH2UCYsGZTby
nD23kxGsyKa83SGDa9cnBqHBYoysEKNYQ8vUpkzAODQRHz3tu3VfSfnrGdOBsof7Mw4V+Lrfc7JE
ASN4ttwWlXCJ9r9tbwUeiuW6romVRrVM3raDFTvBpr6TNLbVBFdb8Cxd+yGUuzEp43BG0tQcgtWP
pitrP/4Fxd0qVIJJw7WUrTA6mGC6Yu+Ml+cfDxlDfsze4NiN/MLRX5i7nFZ2/2srHIjo5d+XTfhz
VfkOeZbTlskuQMrUUV1vkyfzQuqZIiidiRzCuKvIV+ST17J4bodgYU0BxyV16ScI5B5ljseQ3pw0
Ngg+ACmsRflIJIgRDaC6/O9Dd/BQVSWeVY2gTGl8k55Xj3ddZx9BcmbTcyahJux0NSCkk4GU66a8
84I8M27gWTOCtbgEQGdXZ6ACkrcWtAz4ZNCeZsA4j8aFMRuk4WBoeIIM1QsNu1vYG4UYkZO9gSiQ
ZZyKb4O9sIoOYMs35PuZHvA4voLZBe3XthCD8Cms5Kuq6ZJF0KwnZzYgUJWMgQl5ybeeSpk0Ek6p
PL31UstVfERuSrCLMASXwnXBsz+2MQMu06c8w6dtK2u35S9af5oSglHSuVtGMOcq04I70Bw6oTtT
Dlw5176fAXTQW3AUR7AbNWzzBeKht9S2GdPhqPkQJoFG+OLhu88pcpD8X9CDopM8z4A3Xu8T/mTq
R10qvmbbB5OZkfriUyxWqQaejCr4jY87MpVHR69+u4Yy4d99f3lekyVj0QLq1b5q3X1mBlb6uM/J
prFc+uRJjCVCerjH2z1LjyDH0UeKNRFON23OHVVZ4irkon+eq995ehYetdbhf5OhxDfKjtlHDgnS
feudPWqckuPX0nAqtqHfJCI/DfXjCOPgYizmuLVbiD06Iy5KrYPSyVzRLq9NZDvu6dylT6NQ+QkE
ttaJvDmWUJXZ5KjOqqJOCZstx/Dr2IFRz0FbsemFLNRB/DikYktnQnhK6AtAfy8yzgCGYdiIZnwF
NtZM9z1V1iERVSc2pMFdgEl+mSP5s1g3WDNd1SCJOWnGU9Ejt/PH6D3acZtkq8/j0dGn2P4TXrYP
r0QEnMqK8flBxya/6N3aR0HJ5yzqG4MuEpOsvy6fHNg0U4yMUHrxmOpsdNTcZ7XoZlbWNvB48ZQx
eBqdFLgs0pD0cJ3UNnNenqKOsjwcHCXTbtq5hmiGRW88O2azug2hEOM6t3grRt65yka3rfXClm3r
79VMx85+1xAgOF9jEqBjQypOCc+0uM2Z2VvqGQMZQrchG5pmZ4pxE31BNnhfxBc8QZkPCrtTOXSe
yzDk1+hxs8sSjr5iJettLPHr2zGgOEqK+JDsKYQwTEzbudkRo8SFL3DMPeNkQvVVNAA6qozuhZ9Y
Y9JYOjl0jrTMGZDAqHvVxGByn1aRUu5UCggGSDn43HT0wv+OgnPfEVtef0QvGY2WU5ShJ52aNr29
jt9DyNfjkSs2rZq1dnL4/RqmStkpceDHeqd0BUTSbjkdr0pgo1MTtVtuSuy0hR358yH9VFcsCdDX
qF1pVTkT9S0pZmlKLqSfBeJd0gyXiYtMs4lOmFTlMb8qhr9GOzct4rfppdG8A/bxBo3krXzvBQLy
ikaBVWylWP0yAnxj2fE1fVO1KlLsUdCQZVl9yQWbNyDPw/mB58CtOywzhBAdFKutAx8AGbyFaWvk
BTNzA6OMQRZk70E6b6RRYGPszdWc4LDGjQYn0DDtiU68H/whOHSq2F7GX/QVh7+M9xKhppjuHsoB
NjRqm6PlC3fQunYtH+CBUL9wqZaPCqS6+iVAcIlMOr1JYHyV++HhoIwcmqWW6BaQItF0z10GTHYK
H5p4FuRUk+wgQ9fqoDbFgnMlD+2qsoMsLcq6eBUWS1UxG6tFPKY3u4wGnvEzHQ6EAqOzB1KgS2FV
7mwZiUaWYBeOjbSwm46sApAeo+Ry9ysgEKP92wy2KqZEhODgU5tkCB3qfvF1+3VpR6nS+TkY0Fm3
N5QshWT5BHHkKIB5GKIRpY/xbF27I5wK2pMbi/+1H/3sFPe2SEP0Dt4HGSZVvVW4hqEm1OJGMG6Y
tdklX7V2v8ncJHZKYUm09T3P/ZD6aiyv32YJMBV9woClYtg2CiO12fmNX/SH4VRxDD0B1ePWbXRq
veVoNM3nqzg3L/YLPtLEdLcYbfnhNb2ptkVhVAjzts8T5KhlOafXi/E6qsZCbNoIC+aB2i3SvbDR
f27vvi2cW7x4EmqiDYQP/0cMKBOyjs9T8ZB69q+kLlioh5fVebNJSh/rsNjkDG70nVwsBY9d3HbN
HHYouNypNuR2FYvhDMyzg6DtR21aSjlVY1nzdFoP5w99w6/H6E/r9ytRnnkITSz3KIS8zlcoSPo4
SiFHe3Af5G+GT5j2g7KYpNbKrIRQomYVfRqr2lxj/0mrYxStWWI9PGnHLdcM9zwl2Jl9L++aaXwC
R5xe+TErqBt5wN27O6MwzfAO3RzdozntL9l2qE86p7on5M2e1z3UQC3mjtKbaXChXawnyTAW4EgG
42Z5OWVGttODH6gnis2uz3coSR8sSU/GEVqdH9q7k04Hf3+Rp4i3Mwc8jQwQ9Nxyi5PoEYWTUb09
U3WpFhK6t4egmePvC5Y5iI0gr5PDX7uuHs7aLbggCQG2A+gdkDCoEqD8PiBIFHlPAuzweDsNvzzu
W3ZVpbCVVacLnmf3nwf8ve10UqHyRjCdj3HA6mApF/ReI5GpqmybChlWOC4N1r/frGta7asuq2v1
e3oxHeR+QnnU0uZ65kN8ve/6XsXMKsidGRHBVdoDIXCrv4UeGYGZw0kfywVlMOuCW6uVsLnjTS6C
bIYMQvQF0NYmfwiPhS2YynS457CjgvNmgW5RRQPYavPo6lAf3o7Wy7VhwVhuG1yM9hpNxuJT05ub
07bnubmzzHMqmrfg8Hh0TrMyXYyVE3sNxSdiUx4Sgyus/bqtHL3Hy1Zwhq+lPcV2FZWWyF1AKlJp
k4kHybDHcjbdretdFZ+ET73zwO2bRHnDWkrjooAjg6GwhLEZkCdJqATQVBcP2u9N6c6ockyW3iEO
w8iEqJJmrkJLXpntHhxSG85qN79yln/bWTAr1KzungL04OQ7I42sUbiGwlwQiRkfJhjJXdPfm9qO
TgnMwuwLkUnqLVpz5P6HDK6F49KkDXWFV1lZijbFugxZQIL6uWYOQGj84n6t8uwZtX6u1PcZD3vp
fmem2SqdonoPc4YZnpLebuKKWCVCXbN2C+1Vm5r6RbrpCC1p0olcPxRqi4QjdW3AbysRyg01EVQp
OEMCQRp8RAb1Llp+ETr2hOENhsCCmwjSbkYkuC8du/cBVIabqNBl+jCt6W5Uu3gOkhcxYzFzuqta
PlyOCX1OFxgLicFJaTwWGm1KbZNOZ+H8/u1hV8F6L6OKvAN0k2p15hmnijoWClbPg2hLJssNFtxg
lBpXNKYrKol26ILPy/oJ2EjXbdplGUXf89cZAQkmxYbWFL2qtSB3sAYgQyzY5Sx4ZNFVSpWxDi7M
diDcNnQ0MXn3R656gD7FoCqA8XMXG7R8n7vlLO6snBJpODyONwdJcL+vx492i+xncDOLGtyvablm
BTvkrIsOx8GMdcTmLoWTMU6YRFQ57fR5vKKr6o8VpT1IKrm1Fotg58ZXn7o7Vr0/j6oho8mU7PKZ
+jIo72QF4V23uIMDSEn02p9C6UhE92f1Q4eHobdTLqWgIK5mWF5YRvn0RlcabzQSZvSUa0/LoEXB
xwTFrWtudpSKevaPmH8+PUgy7dMsJYB0qOR75KLa2r6hJqaFNty5/JESMV+D+XMpfVcEYoZGRc1J
nynXZTHyPreXOEwfYLTPhsdvQ0wtNrAicZltlSi4HiYowxYSxbnJ+LS9ojFDTrYDrr0b+1kYAlVs
tpLlk1T+4tegw0u2OUafh4Ll+Lls0zwxnYyZvUjwTiE1k0zO1NmT3VmJ6pttKJWLYPjlCIBFGwNB
8e+hgORGHE9iN4U83mQVvBm2TVNTUQZThppGgVnWx/8oMJLBDMfuApmrOkGCsNnHyx5sOv7XTPHh
cS0Ke4uk5VvDE6G8LDMStVEqI2M3MQJAnj5BHQpuy8iU/JnGRm5Pxvj7tqsreXLWrfQp0Hqyog6o
2tWoEx6dnansWCFD+Nh4t4xQSGnk/7ZDaIDTxFuHQa72h1csFPd8iQfV+4QZmZ9WcdnAz65Yaiqx
O5metpfghdmW24KJiZWfQurK8tfriBLtddlKg8o1qmj5/fRSmy4d1v7WuXLCfrzAvgZUJWWXCf1H
jBLX//IQO7MSUnibCDBRVzjSeGGh4D7rTS2WGzEXl9J70qyRJdbjLs3SeYlcUr1YeZbn9/WzUAUY
xB6sONp9I7L9xaYjguBGdK6HLOFlnemT7fIo1Raj8/B5dHZOsB4e7pP+lQt/z8/hpHsxrPFF9c6g
oEQL4kDzZfyZgEt8ha5uavka7WuX8V9b1MRkuEIlEDAmXwHR5ymuvcUQ04yK6hXR9rdoG4c7QzwD
tWg8DKFjVVZ47B8cEqBhP68r/DdByqpANs82ufD1jJx0MxiYYfs1+YSbzG0RpcUQyAelH1t223cx
FOEoqjwUPwdy61Sa0ubXBoXUH2UGeFpwpn3WoApbOQkGAbFiTZROHfp+kIYDhbj+AtsHauPnmqiH
kNrwS4OL74QDZ85mgaU8Zh9A+BYmn5fBbYxTGcOpmFJSfUKAz7WSM0oKWAzSrzKUOg/F9EFQ1J5D
Y+Hjp6Nm1bvH5RcSALRF7cz/X6q7YKTNyn8/ol/3JyuCfkHoqR1VCgAZOTRFKVW4MptHpPK8Rh8k
bhwneNgJiVNrI0lvTs7g9L6SATdpGTYPui32WQHG1gXInCL4b+Rb4hKXJbn7Ml+48ohwOjcR/5zb
tz+Ametx7SKMAN4b9L1M3gnVtYBNv3BrBNw/q50gInUG3tzWvhxMHFjF4NmawaFFYMEZmV19ZiIN
gG0J7yA2Izv9pPBehhldyQN3duvkciPhfGN+Yuv/kuh7kmy20TxNf/MCoLjwFssTUZG6POhvLhwR
/YYzkBgZ9xYiFaaUaqOg61D4Oi+Dn5wHlDyJ92T7uhjfeNEL0EIMBH7In7Hmxt6M0qPtwi/iIG+6
JasEPsK1+0yX8CNyiP8CYUBWNLKVG1emsu9oj/dKjxNIPbJLSlilNP+/PHwr5lh84pBbh7DyZPbE
f30P8D3Xv4OSK13pfPQCNgvqPTeOrz8POw8uF4lApMN+o/LQeyDi7J+W81E5dvJMW+Hy+/9xuuuV
W6nh/fhSkqCDlnI1Teu5klFDmIc01ZwiquA3FWciKjnhZpSDQjrgxVWmGfjXE/TDigRBvgJHHSgI
a8xFSDdR9VSh1ZfeUuzU5LcAOe72MlFWZdt3ELjSK2QfKKIGFx1AfjROuN693b1O7PQukXg7VJIF
JdFJ5w7oCDdBgqgdpCmcXIk/B5Gmh26xjUyZmO8eUr9V+kMP8gksKM9KbxcX+o1KMNObXbZ47QVv
y8r6bSGy6+yoAzqHg5vmTZb6Za0yN9pVapZL3ApLaEf1TLclXl3BbgcgKoPG2PsJ7JtuPOxRaUeG
PzBQc8RI8sz7XWf+EUPH0kTNWpPDZfd1k0yEVyO7ygoyGHNVxMfKYiskR/WHXEHbm+Y0b8t/Xitp
fB4HiW1QrDpOpX/DPZ2C7DmF535EuyMDDRY2+gwGH+YuQD+ZwMrJNqM6tKU+YN52U/LTGKU1pu3M
pQGW6v9B9h5fAcoKZgRfjvBjd86pGRlV9msUiiL/c1xK6BBXKG+Amc/fCYyqIDVESp78bgAW7lRu
TW3FImKR9P3CpbXBk24Y6P7oj0zq2V51X80nWBYG8H+bJS1PQjMre/wyWf/RQ2J/7OKPl3us88KC
sxDTJFGdo1kjNPV22exd7LM/Z9R6jQqwqR4BeZ8HMXZ56k5Cy3d8Qxmk4T9z7ZtbLtiNivj3teNS
teNpom8PIXv/AxComi9qfOqOgMnaAZG7Spzt2JzHcm2hVDFm1UrMAI80ObylbwHKt3boTexW/18v
1mAKgm6i5h9d9hyio6gF3C9grMioxEbQUyJ+gZZaZDYF1IlmSC4ceheULoHJazj4SgPIrioSBwZN
wGcng19G5e+4WLMFBBE9RyQkXZvSLkNril8/sOmTOpesE/csg9r2yyuyiNr4iEOzYgX+n7HeF4uW
9f4cCsLtbVl+nEv9kSXeVqpMnB5qZmu3UNHhD1x7M2Q3WmeMIAoJIHtnWDcEYxuHnm5UDyNXLsVR
Mwnf3PiJBVUlS0U04nQysN+Kop9t4n7wMLd0SUnATdHD3sArBe8lnFJA3lQOwBkH0Hw+xdy+/Ino
LjhqH1eJg74uLxeSkfR5z195MBgCAX8OwkSBF7u/sAf6mYWe+X6eW3jdM66AA7YMV8GzSBjNAUnl
C8/hu0aIDZ0PBT+ldbIy0BLW0AuLKusfmokyHtODNWL/Pw8LxmIoaPoojZAAVTQbVHaLE3Kv2Yg+
fkSfpF3xsu5u08+Bb9AGTOqEG/PTuVkYteQcCM6JcuE/zZ0eR93tstIKqg1+bZROzbxqheSuAkmz
lG+eKOvpcPjzAev3VXd1xAUDxFhYy3ieCS/VnHIzyUiDx0FHnc85Hlc6sGUCSKiuWNrwGZNW0kZR
VUbpuBHVezMcN7opWjS1MqDmWjm3atmkIOlvA3N7Y5xmc3pSRrTB9V0JC2UWlQcm4a8/8HL2jPF3
hna+T3mnUxYEKdJ2X6TdndAOuRLiDWu48pi0TWwbSjHqqmBnLeroNrWik3NqqAdYL7fJ4JJoVVR+
u/9MRc/irEELY+YAu6Yjh/lhJwEExZHJSWdE7cppkcey7W5GKYdJLiPgm9o2xOcw0uwJcViwLZTl
JkyoJ0N73MGlzbFdrlKebFbA61fml/iw5ucBxmnZqUiUMrnGZYlz17kqmCji+jnkTz3BO55cItxe
9XE5SH8qXLfCPxSsLZKuDhHx5ugTt2yFjarir+JLIGi1VppH0qMXUAnNSbwj1HJl4EeLbq845hAj
7S9OzGnthDGDCLxFBOXB5dBsjQRE9/KIHIsz1KtG8Vl1eBo/2amX3zoXi/oQrAsYvpxuaIr0c13H
l/eaYzWFqj++/UPQaydXEHC5oghwOdWdC7hTz1EaVTKGuh4MoIHFHK/mqwD+nuUys3c9/zTU1Xjs
GedsGvn1KRvAaC7/kmKR6MK4HmXO4egqKUD69kX4CQLy7QPayLibBjoOb0Z9YcZN4Ku/1hCyz3V+
1MPZZsEpYXeaGAvWxoBDc7Zk8hgu0/ydOEpxHYVZcNYY+xRlm1Tqsd1Nsq76aH9+2ISguKFgbSA2
syaCzz17TqhWVjMWFDiqA+Kz+uoWQhzYUkXJKI5LI8HiBu65640k0jdlpY5x/PzviZrLL4exaK5f
dXZgsxYAaZ0u+bEqRusec2AIA1/50G+fid4vBgGkrm6v0RPMz9AIXrcmEKQlcejFUQV0WAGrMN3K
p7vNOUUgi0QdLbZhRqf5jOTDZ3acedYXwh3SaB5OJUQgM239MFOKw4ctBrW1lCTbr9wYjS5Ipvvy
3hFE4EwL3mt8MYYb6LirwoGm09ZvgATkqtfUIR/KuKx7vFEjxyqFbb1iqNM8tenosFdaxv/70ygX
yB85COzScpZKL9dc5gNJaJV2digS68e7B7MEPRkDKhC3PRrg6ow2NVK8cpG9+LAwrFxSqtaEivYN
leICB+ZgRUf8dml5yXzBzXOAUkLBdQIvWWzn4JD6XgC3MOzCm7Ls3VJPkUZQkLId1i0Wu7dPWou7
TLatAL9DdkELRXFRJIFDm7dpWjIJs2LvrU+T+DUFeG/KQFhBRszMVU5CYuRMgUsLhD53Gzt7n76+
2mxHNBKYk5m8qR+k6lc28FBnS2jnHf836u35uH4kuiOEVm6kpNTlFQ2HLIKtuJwg33TWwLR85rXZ
OyVffNleaF4eN/uQQvTpc0HU9nQj8I+YeowiPaPzzpmmTZD9dBMGB46FY3yVmEhMPIzXeT/UTEFk
qC2C78f5Ygy+7PinhyDql8mSvZ2OHPzqOXkUtINbhdSQLtCz16Eu90D16Q+XfCiZef6wdE7SITo+
2DejBSAuZiRsjj14VMxBY2u+R6jT3OpLvYS3eNBLhjil6/bv5yXTzlWF7Mn800daxkoSisrU+Lr5
8rW6Wi6XxpAfTgyaF6vOFVzZmBuyyu4tht4JqF1KSGFIgAlSRsCWgJPCxWORxtb+RXDqujMj6Mvq
4IsTkE7H8M+ATHuG0U8QX7X53LNxgVaovNKBp+loV8TJDLMG+//qDnU5bA75DxjYDub1A9+LOv7Y
nK9PEBYJnmVBwPF3RKCBg8qOoPFTjwhoV4o5nGfLAPLCv9f+a3pU/nCymieMjyWlZ+oROD0ECws2
+pCjlEOoZz/uhWUruV3IcKvvTGeEitNBxgciDxB/HWwYWPJ1Z018bHkv9qhhMzexq+idYsQaMxzS
cpelpHNrevL4U8U1b6eR7dio4N78kVpgk7NSsHTTERoImSirMxBA+19ygL7psmOCk+ki0CZqkqQd
Mbv1hsBOsdAii0guQISyBEhOYIsdG0zTfb7P9ef9iuSCmEp7P0Pyxhe29t0RUYHPD3lQb9rEfqAi
JnqKKquaEqQV5RD8HZnnpeugWvfssZ21hqoS12gdpM7mzcd6mpAzX8ev0Tep8qoZOjj/HUT8R2L2
OE4udcrSdcZi6Wxo4I21FAQoVkPpwd11K8AWbh03k8bXzFtQHXmQj5GJYbRoPd6+lPEVpsZVMUsd
szTraxcCfuGsNyTANV4W1EBdghOCjSAL20n2mgfbcbGeRgLGo2c+XayhSAuTLpzN1YAcUBsEuK55
ziq/xU0yVC956cmov/bllFd89PnmnO3gRg+APfY63sHOQGHA/Uju49Lsz9Ad+jdPaFLh78xRPEfg
Be00YgLPj4xLef2Fh/tS1C3SuASZn8f+PAWh6G07xf/rnAKfzMwXP4lO7doj0tROy2UdypHHX6dc
A/rrqtlsYPHZwOrYDbYa40v32nhSIIGiZMddK8vDNB4p+DZuiJNVzgOlCYn4EXl4mYP7CXE3tmS7
qrvRbHxC3Kmmk7E4INO5mFXFPKEzhM95j1bdxmfNTmGxmn5v0tEo8NuitH/HwrvceqV1IU01MEnR
5BJtF77pp4RyhdMP0FVJgBn33GbJ0n3sqiLZVQW4M4QRAtYPe52odF718ZWUDHoDJvdFPvp5ccIH
GTtdgb5XaeuLXMEN+U0QiuzDp6xfgW61Emik5uc+9amVMVrDc8wudUvdOrpsZLrt1CVJTvGHO7cw
bM0QzGcvFVLAJYnJmiQRy5hEbkrKZL06Usf5XIwZ8Kd4RgMx56mnMo3Kn0I8bh6wRsESwsWYUY9G
5lAJJOHbEJqKJz4qT35DdVFmUP1msSUnZFF6giurptkRm45dGUTRR5RswGE53wIbg0ZxPf/TdB58
wX9wj6E3PdHhzhv+gPa8Tj98wSQghprPUTpP5QhN0cjsHf7n5DpfqbkzOvqCXNMN9fETXjHFSr4N
tH2jTfuryAPelapFElQUna76Lf4dpzCHUtHYZgtYWr2rhYXTF+EMUh2pHLxvNXZANWdIXwbj4brK
k9R58IyRF227C+fL0m7CLUHUtiTn0ZwwyeKu+ygX5qTG2aRSTM2G7DQP0OTWQmX8sKl5fNgvNF5Y
jE2o3bp1pOs0k5MTzyotm2XybqkX2tRiMAfoB2JZiP6djG6ztxAdy4/eyASaCYxPaCO7JpGTCqDv
1e9JFzm1Fc4MVrFAHLY7exucpSfauUbF0tbW7nHRYs9CBzaLXgX3019yvgcrotYk0t6NusZLs6E9
gbRAjE+FnT4bGYIMrI1fSegIgmC+xySFqsWXxBUiLzV0whgy+d/67+Zgr1wQ7rhMshkPhhPQW4u4
wJyAQefzdbqtz10SrWcGNYjWsJcJT6Ks5ADT19d3LIAcrSTqZti4YfrGNMj+9odZp76pVn7uOnhg
Cp+Dn3FdOTqbV8etELJTv3T5IcJdiJkbJtnaa+pW/oJd5P1aW7hUGb5MseIV7nSCHpVsyJd6Dkr2
WLCseChS6CKd7jwQJUWSzBlCW+f1FkxOlPkjfON0JNPoFqe0zhVr+cGzLvK4q3BKk3mmBpYXo8EU
3qiRxzj6C0FNNCmUAwhCWdeQAA3E0RLSyiVv3CPlpmtAswYP7gp9USP+54fKQ739eQiwY4MMQWR/
J6ho3FoP0jmz1d7g3I3Q7sMb+UQZmukB9s/GzSOF8vD4qpb1XYp7uQxau4lAqyUUKIMdE4fL9OZR
1Gl9y86kxYJE8i7QeZOWCvrAF7jL0aNwC9Yw/U/uFBz5AgotZs5yG/mB0F8z5KJlpJbHNW6C4UEt
mSlrkMokhRDwv+gzPDlHqhZxQEAVDugq/+pFfMlB7zIhBWUYTcYDQaSpdUJJ0y83CBYLiyV8yumu
13aE/mTeBskAgwOOdI3HLi/uwGZNl+AdhS2X4EjYHxQ6IFSr2V56noyMdX2H8iGb80RshsmXKDo4
AOfkMszkviFX5MewXZcMMBLU0MJ94ktmRTSNGT+Hiu3NBKG8UbzdIcg49JAalJGY0VZlNM2bKI2i
2oBUBgrQblN7ze7jk3EkQJ+xDJOjWQnB32+hv6y8s4JpxRKxfbzyeyqqcNkcuAJ4QnYVDE8aNd4O
BpLLQ3SQSREiOLir64FpLKQojbfe8I7I/CPxR5Hyf8gE0ZVCrBuAFVxftyvPKTT5xk9Kpufmu/Tn
boLrBVlBo11HKnbRxUiihSKL7DVYTWYj7j6yMKt62teWiMPXG/wjSmO3VmCYMHHjrcXHnMzUdFNv
0TtQZ0OO1CRApj5T2hYpsAhXPeVClkEcyN7kLuwlU/rj7sAhqBt6S7+tAYe21a0jVzUvWwGqrV6f
cu41k7lgf8i8UF018fRuln/C94gRVewGnqSxVbIRjI8Lzi+s80KAQFALmoqGgNVeQ8Uibjc2psyd
YUtYQ6HHJYnfYXE1erVcO9u2n5rknuRGG5jOyPDREUa5AdivprpkJ/Bgw/NPr+vVA0eKvKvY2vnT
u7rGhnBOq4m3c8KW25Y6m9nLMiEofUxZh9I7s+UxaAAYJPjS4S5hR28cajZw43D9ioZYOY/BPfFp
xdCICWbU0O0bFzKYRONtK4LVfOB0h9ClFZWsu+KOymqC5Zxn2AH6CBFFvIH30bsnmtDNbu+aSNhu
kiT/PiMLsdOIfZ0HrgsEFGsyBtlRJ49vdLMG7u3UyIms0l4/Xagc+5doZOPA6eqmOg+YT78kjMX1
Fnk2F4+4bE5sKrz0/ZjRi8TVRdnuPo1eag6iSYmTiUecPp/+mMnii+5lMzWiZs6lI2NDZW2j6C+l
GcTC/1e8Cd5dlFrO5ofv0BAPSPQcmHxr3jQdQKEQHGn3utfF6u1R3sjAV5cn0Pp2lBVtOhJOzrCZ
GHkzpwGj/Y6jK5R+gyHla5fOIYNc5GxVra4Y03HmJH9HmgWAdgG5iY/GY3SgY4TbsBqSh2g4WC8w
horXwYZifhPggiCAiuAflzMFdnelRNSNAPy7/4bC21fgIr8r5nidejJgr7+3yU6/eB51watVxQtn
zGocDXwAt5oAISs9jhyL2wFXgbNuyAxx96ZFzQ8yJknyQgWOdgzMuf7Ega+YHQmHWzv/x9oUPhKW
ZtiK9dp9T4pP7Hlp/PMWsW1x8ioMyNI8JIjXpq16XRdJuwCDy9fLnqoMekJbKQGAVxsVdV7Ucn8D
P37te6CxxTtpxtgYPXoC8ssAXUxjVD6HDPB9a/FVl9nBTd/poQep5hok6KHtPdEAcRY08RiUUGmm
YISHl7bjAwERNv0GCSy6fWYKpYK5Ygcobj14r/xVm8uj2c2gbwmWzEfgGsCjC+IXBf6+OT2oP1Le
Tn65BrMh6cnlpnL+/j4ixwA3NLsnabqX6kNgq6ipoikb7Wr4hqUhrE7fJjd9CICri6T/ymOjuNPx
BJdhBU1bMjGiOXKD0+6tAYNUpVYAi76MI+o5gvbl2MaCOcxn1TsPnLD6eFE8H22w2BOD+8CR1BEq
7nbjilIcUY1xzf0fDJV6783Zyk23cDE1HeGenJ48hpo+6diobO8dOaA5t5QNvx/cehP1+bOLFjw2
+QH4VvTprsEThx2gFEEu0pybHSqBbYNHlgBltGI24wRM6r1NkfmgOTQTkxMx2rUQNcyt6nlCC8p5
s/03YqEcbgue/AXh6+Nv8KJP0M4dzWYz+568iZ1esO5yt4uinv+vAzLNMzyr6kmlIqsyymmYXypI
C7a/Cu1VGabh0khgryWtzMCaMowiLadIxithSDwm8jvduab8X7UxJKlFHYYig9I1AgoBMAGM7NKI
rZNwTpPkYVZeVKZib3015bH4rGYAJ3uvD+UOLYWhIR6zmujgAui8G1/VIfiHaujoUoUaK+kk7DeO
B9BAxfCps3N3XM4MjKMqtVJJiNoqorvrOSUmMQpLnT9/zQfllqPivoIC+uz3DhQFohv/4uGGaSUh
RVSzKmWufIZJGSwvEZYYUEbJGkcaaUzJz3EfqEFrmlwoUHawrLYhjJnU8gWiE6/3is3w/gS6G6XZ
catT6okGUWvVbVdU+njRpVY2GkcTmOuOopXOkqqIl9B0y4OtsYBzbV2vBpXlhqdtvGA8crQ3KGlA
6TcQCwCimX9rz3d8mc4U+aRJa2I5ZKy/vsodUuMjWO7RymTyNX4PHBiofyDA2cc/gQ35VsgjeDpp
xfB1tZMV1tlibINPJUBaNk9UE8/8ladCGkr1jXxTaLxeUBY+lr9ibYtidinUxs1ZDvg/kj89bte0
VbMAgUpl65E3RWmrMSCdHsGYpqlzk5pWKazNUU/bQsZ3mQvHIS58H1tDx9RJ1QQR+GTPDDmbdn8K
3vC5GGhC7uwzLRIVvEsgDKBNaHEAKVPTB9Ek6PgsAPEeWXHOJ3aCdvlYgfn+1yEgDvu2PD0v5E0w
mvxwUOjURDULW/pHN/i0sQkbT3Hh+obIus1aTZmyb4rPU3UGB03q4dz11v74+tX30RG+ZCMGuAtY
hUVhnSLNbwAFhUg3UrQV8nLTt1efCd0gKlhsbogeQnVcvzvtUWCWpT+JHnIMYN3oUdA4CGRYBdJ+
S0bbLVGoyFNBaU3+XDgL6WyxH4H3gc7iLw2lX++KrT5Hf5OtMakCVVc4E1P0O2wPpVA2piCAh/9/
dCc6FG9EN6G/bhLsCqtpPebTsxFPCzgKQK575MzIIDyiu8uBLSNBc6jcu/pGn+rGR+pZ1IgnngsO
f/2EUBbQtnHsPvztci5wqg+tB8Cw+zzjcUqCwargAyQGEWTDCEDNKf1o95DGPWZtZuDYamQQ9L6H
ZQI61dwVLHcivaGZTJsTyTOUiz5Sxj75usvHGCHN1H6IO3vVDNRW4rR5OchcKwltCHD+DdggKRrk
68UkF/WK/KNpP2hFEm5OMz6dhGsDLBEhaj4EdZv/1Z/w9yntsOgrCUcNS98EZUC1nwNbQ4J8vYG7
eJWDNeRACZyepVoSJ4C5YoaCheioCVo9pMjNCpMWFA00Qmi9XOQzwmfW+jU6by4j0u9md2vOoLMm
TJjtLnGaw6z5ZhwIWKiqeUdlRfz4aJGUnix/KeSJAImPNJS7rkur6VAWnvWFUAiv0TJ3vYQIqSaM
6izf0mf/YlSXmpt+qRqfM7RJ9MBB7XEIHTMu6tJNJdj+hzFVv/8f3Z9RuW6wtThAGrcEMX2yCSFp
LBtjaQ4iGlbRAhvpS/tsysiiEs5/vM7OFQDCn92SmqLpU4nCH0CZQ/oFIlLqkBO6tjw9b1lMptkV
uAfkdQ2OhRh50ZT4z0j6X05+Ps20901osGDSNoGDLKg1GyJQyQnGTNCiDOVzzGTxNf93/uHa1yC5
fgDhw4+/ZzG5slInHL4xvCezYQUjrtDOYz/Tz5sQWsTBmzvkN4TmB7FFn4HL0fIExhd/pKXuOo+s
Z9tRK3gpp5LEhx7GGp6MZrc23r2rHuL+2Wxc9RhV0VVwUbO5xoYgKnGe1tsm6ur+rvXZewaFPC/Q
EBn5Qlvs/owlZ6gTl86o9Jq3kVGVpEpGhwc18ql0v/1Bx8yui8b7PFSuiWKzJ1o/tuVAH7wPSoUQ
ing9o9w7yk+WBY1b0GUOAndIeRnprCF1+OJ14PtkU8gTLfGnG8Yd6KaE65vvfDsC0MVp71b5qBez
d00EX2wf5V1qGdblEFhds5O6LYDn6pmvTbZLdlYwl53AjaVoraR/yxoqS0Z0kvcPnFG+4FxlDXbo
bUOy1uDToay0b6eD9UBbTADPNZX6JYfZPflAXO1buXIfIUg5AX/3Ma8V0shlqsjRCOev22w2KYtu
bhQ7Arna+6wMzaMFS/YUZpE1D+olGBuK8/CBt0FncrkEWdWjp7Vr8igXaPqHhHJZ3jn3LEZS5JOE
E2npe/xrd/AV5TN7EJzzZPqcgt3q+o30NTLlYj/OFMLQzus4/gtDTHmrIjQdyvAq+S1vINUPGXbi
O0R8RUjv1xQAqzUKhgEtxR/fI/OCeydnZvRK3bHO2cpVCSiBJQxtiqGBiHz4V854zFqtnFax9Ig3
E32NG50nSN7S24GZ3qT5SnhnJ/yyDHPK5uKGP5WgoSZVsjSlAGDY6Bo0PrwL2MqR2jgK21FAHHrc
OiuzYe9f63vwsOPAGdlsRwwNzrJesU70JU6ZMYSE8JmidO3OGmlkhsPIfyBWbqsFbzIHThKHO0mL
g66i5ChAfrpkjBHmVHTM6FXbZDQd0Ji+S/Id4aFUI3yl0aCHNoXKyuWNpc7DB7VN+lxBKcge4w6S
qCfJolMI3DfEsLQULAREq0AgQfIPMnfUQ1I9Wx6QNI9xxf50pZguGG7uQCLWZ/z3GuXn3eDzn33K
PKOKcnFE6O/R8NK+DuuoNqAdabdGcFnZgmhnM6Qf4xQtRETd5XcpmDljQ3ewWhAx2yBgmcCz2WgF
DtD4n6GJYOrJ1grr5/55DFmTeObRqV+GMFDqmy9r2gZXg6CYusa3LmAnRxtgG4tg5/ho82ofhoJi
7ucUi0+aUNmc3Z0/jd6Rrjhz8sLTjhabiD1Q9iVof5fC6+V/KdWGxX2eBwfwVWelT/ywumBtHp6B
MPFtGtoe4MVqVcOQnSy/3VPGTSs7DswerhjzSqc1XSXYX5VwzdacWcW9oNcxS1KugVOOsampkqZf
0Ccx+9gKmhlWI+YVAhpnogccbR/eT8hYHgHFPzTdvv0xX6k87X7ajZOj/kUZc6n57IDN+DLWHs7O
zZcIPl8GZ2yWnj6wXaTqjIQ+h5fixTawClchMxT4TevLyWbZoYw+OxT15v5v0sqrlZCnElPYsI3e
s8A9qUfUf/TyM6qLuS2ip7xdTHgod3DOhLRgldf0tBPQt8xbPZVTzWFrT73p2WMtBF8r0Wo+Pkg9
YTLsEqXP+bLIG9JuEAaIVeCZgKUK4JhzHRe8RKrGyhtapws79mvamOL4dDE/x8H61NFO+SkkmuFs
muBD1piDD3K+pC19s65YzTpZHE9fz6XRK23pMrkxeuu++ryOp62Zwdo804TpL7l26ePZAOA9Rn0h
KJqDC06Y5b6I+DLMdDHTIaEH/px8cFYPfdjox1DZOXgz4uB1Tq4Vebf5mkYcciPlK8JvB8fWZoYm
ZSqnW2wokW3mFtKdWdnIJhcaRDiEKamrb+6s/whmgmq4z8Gn9mToRXkO0K5pJ01zTqPv/CQp4lwf
1qKRKx76IQptyjOshHFhOXVyzdmgdGKlv1iDn3rRnQ7EKnTAAf+e8MLJu9cvZpbX8aWm4wv3BHfx
MOhmHc0UzQt8NdEyb+LomgirkB20XvcZ0ggRkkdaWU6av6+xZCU6kLKuYH6lni10pU1TwO5EIVZr
Vzvh8ESkqovWKfi/XClPa+LkXOsdn1rhQMSQ6SivhapsWeLB++bfF/mfDmcCTWRSM4+m+oruE0wz
Qzuk1VBINaLKZAl89zWcIYfeLQPbH05O//FCALNgEZQExEglOTyFpf6WetzqvSMrUBySr4Z6h+NU
zLebvQRulXabT1LITC+r3CamoR7HO+aiHZvbpkRMh8PY9gglTRPKglph+DKyeuy5S5vvrOpELqXN
TrG/gfj6rWvgsdnVixjDo/eV8t6/pw+kPUpqnoIpYlJus4M8PkXHKP9VdD9xuD6O58R95e7uqFvX
xD1cbxvS9U2QcggKW4tatDuCGAKPX+a9HXvWVK/3PHedwWkPBo0gAYbksvPveygURqTVwrHfjfOZ
GtV7/gfw4ImqY0T4r5Z6AivSBaymn6Tq68evBBHVf45oeZc1tz/zJOHk3ryzhluHwVekKmrsYgu1
s2xGwWEJSds26ySh5DTBKzj/0lr3RKWVhzsk/zHeTss1ZCm33/wnvazpXG7dyb3FLz4vvQGAM3tb
e3po1D0QS/1rqUiFUqv0WjxyT6hYNxdhCgebLaEJzFuD36XaM5vjXdct1z9HGsQbV+3WOYJlUcfu
9pfFgTZmIDzPE2FDRX+gvxR8vkduAeiRNfkRH59wXaFxB1JT9lKBf/7LPmkKIYBpUrBhFZl7PFCi
mEZH68pzODc2INvBwK3SnLHJQDicVT7MSdKgcyEcbfbWv33m9taZdnlM07iDQALYPEePoO3C8/JY
dOqJFr4tRv0iAC6gJ6UbCFkWyfSDa8Iu3wdKY9Ode/7uYB4f4KrurFf8q/hm1XtsAf54KLp/WcCw
qnYLsulfh6Us5UTF0aimGOcXMujLtHbB6sCA21rqEtqn7YCohHuXI1b51WLKIFcwBrTq/eSupXWg
xsw5SCjANleEvwqvaB5vKB36gvzOEZuEf0vTrm6SjwidGbzf81Frjfn2rz0pNGwe22EiJFxT2MZd
dxpulUwY1AH+qhPrzJ6565ahHVcDn10O9r16gx3bUbk0lvPpHfal5A5iMK7/TyluIlDJxiGbdoT5
eI70FdPxCKhdmK5NGc06cZTkVa86i4Q/l6b71g4pE0p4vCeyxbsZ6kLM0ZUd2CHUh38ZCDt4clVj
GNh6R1MHGbAnBwhm1AfRvud/3Oo/sq/1rs+BUt7qzg1WWOED+PrDuSxzAxG5ab88+xxh0bDGgDFv
c9u56al70JX/w3o98+IuHs1MxnffBl9CCf9TMooYuzA7dWe3wOjKHQkekneASnyu1uhxTebw2SBY
px3oLsbJkofvATu5E3EatPa62qQTirpVMRjc5XL+zZMO0QL37hB19YQSh7Fx4DKnVEdHR8nMKI6b
aNRHwlZkFozVJiVtEzznC50mbSAN5bBgK8/YH7pw/PIoidAn82kF4Dd/Xm+qeEKZZ/hCvPeSe3b2
7H500JrZoBgW5fW2wXAaWqoYrWayNFQ4Ca0OShwJR2AYxvfE9ln+vV9O9HAXsdJYse+9kkewW59h
/dHl2qjDvEElwGOyPFwiSe3Kb/Gb4yzkM9QvpwNztHm3Omr/Zq0du1Ql3pzV8o25qXxhDPwuwJmX
RVH/D+akA1ye/Oq1RVHnGkU3P98i6igKOhnuecUSV+71cl7TsYE1k4tBsqjYXVkCdaAWjalg2TVM
quzAXmOB4wQShi2dU3W9TY/go4h6epTU7FxmhYcx+MImrR1ClWQaiT2jZ/h1D00r0BEG2lwUY3JZ
NoG5BY01r7OPKpd0+3Y5Apfxba/fAtb+LASKbdiVp4xpZte9Qok8F3xKH/mWBp0LqO+QtdrQpGxd
aPfDlLo/cIgZZfHpYgNdWUKbh7fAa/w0/JJjWhNhe+GSTnqFmzMckhNQARDwmenaV/l1Kj9ZsRSY
JLhJCV5FsS5V8XQgCpTIByCrO5iUdtcvndtbiGMq4g/6W25ZQRiHXQwWUmpOFa6Xyy4+TPXUYHLF
I1tKshnIxKX4En2Iv+KTG/WDEtMCWQ1iKT7dclK7JUWxNwWLEig8o6JPox6BiB+nnYEBr7TX8N5y
9MA5VJItbOGOeFcYUadQAKYUqTuLEdyc+KuRkl8F/0Ged34ZQwVxEbldBPEfkb6z2yIL4C1hI5jJ
Bdz0+YB9Q7v//skk3hFiSrjn6fvQxGpby0QTDhJAczcEJgxiN98AC2fdPMhcgBH88i8bu9EDA0YE
R/3w94Kr/DPukTFwkOnTAVb9HonxZ/ktnaFOmYK4orvqZj/mJsAjvp7zxlu+R7t0MnSe8cGYh7ZU
WJwcSEeBrNLi/eokTs3DzVrLjCz5nSoXOKiWnXCLMyFDRVKbmmH7fCN7KrwdiOjxSV+zVgoAnYhL
8mdoLMoEVOKeOQ208R7jiJtKrQD62yfHIV2f0TvWb+y/mweIyFajI2VJHyl+us0NGVLMPw0+dT9d
3jSIggvA+uywK5nuDggFR4jtbl2HfEcq/oWiTET1yp4ZWDbSZ1lHmbS/5EmW1VCDnvxXBJbM15CF
8KAvCP9pUxW2NJcq4AGjXRGrdU3Af3I7vRp331nexFWCsVw1XfYjjxm9w+gXQ5ykopTgc95A16lH
IQ3ZihkwSBtrEivajFg7uozHm8mQ/1MOQxRR8D/v7TKwZxcCpwBt9HxaxCV3dtdMQtaFbea+v0nL
2dHdmfeiw6i9GHKFQTJjipksyhliamLaqGbjSsi7312giCNB0z8kfB2EqgVxV8hePtFmMtbDPji/
jK3WPyIeFoBBs8IFYNDeblgOCZg1qVjqS5WoISjQSI6vkO88UaqWW5yzVZXoBlf8sPLwZ2sP/14r
ZTDQ45VV3lThNYLjUAmNIJsSF/UogdbgD5zDMgWxrK2Q1sQBBBM0cD/Z9rg30nUeG863Dpnny+0+
wRplNchlJ2AcTkaBZEKO58nRI7T9jNhc9FemBuiwSH0WtTkR/v8FRlljVZaNG/w/bR4d11ToX43v
WLorp7FeRR3Ux3QQX+l2E+TIEAYIBvL3U1R1iRa+y7fm1EZ456A9Ik93xbqiDybtREhiOfjYykso
9EjMz7oYC3j0dwqSjEb61ofCg15kfR2BCFnXCOLNY+86Orlgtf7AnHwKB5tEF/s2IPNc66IqFExA
oMrrCTIyE1fTsCnx7R7hZtTn1WCUFGO89590J1h+BzKpXpcU1+a4rrgYpwZSmLbooVsz/OJEo5Qz
Ayyv33GiHCNgQ8YKzn8oiPfQ89gjG1YASd1NXR15rAPv+m5ObFyorSLm3lQvHiz6YYBTYkN51EIM
pk76x6NKTAmcMytSHgffScw+xxY4kM2iTSBhrwy/Xdww2xEM+uUOGwkiGtzwz3VruZyrOQZgVSKS
jg6QK+Tij2aVO/sUz92z/5loy7fS/5003HRkroX/qhYaiWupHFyJzdKNiajPJ8MD/6kmdqTXi5UB
1rsa9EVeMnFyhWCB4s8/FzuRLTk89tzHL5mdzJ5PBAgxoCTM4t8WrF4aaN6++x3yM8qNGieko8Gd
CGGYmYTCV6HviJLWBZPxoUocK2p9wa1nZCP+jA0oqQogOQ60gDhbAaw0P+d6Da7VlfzmacvBYb89
fXrBFdyWbIFI5puIUzCd4QQwpIQZGpprwyAp9i4wnExL6Uu/rOhY5DSncGumuhn24iX4fPRxp1KH
ZkFu+zXuhhcmqSAP8mXt7tcGuvpNr29b6QMH2eY1U8f1oUaO3C5t+aXmYx0QSc77RvEVTMitIjzs
GdiOAbCRTrxwqvMqPetFbWk0vYYXxqE1JIdWZ/Ux+CXRoBiOj9jIfq96KQ2qG6HOGaEjMS2eRacf
kNmkeZvxTn0EWT233R02+C2oKxeE8kyUWb8GUnEIvDBt4hAcpmiaKurfzR+ViznzbziG1Ry30ut2
CE/3PD3K47uDkWceVYg/0afrPySmuJVuao5hutIu36YvUdu95XzAD3E8iRTvX5feidcRL+sF6+bD
hsg0MKp+GKIhCyCRo/wFdRBNRYtzPMIL9UHfX+hf6dsvSGpFNzFggFiHdXHmqJQRkJybEgdLl+yc
yyUQ+QAHV9nGKwMlhgMKQh8x0I+FYZ4jUCETO/qUCGweICrof6SsYnlccGBPtrqTLGy1J3njE+xI
uS4HUZpsHoZTpWE5Hystdgv1Z4IMzLA3oal6Enwy2hpd4bSwDkq51/oiQXTPuYCSRt/qBFh5z/eL
Uke89BCIrJIbrNWzEEoClryv2chX42TjgYNG8yl+Uhl18NUihaHsynFeey2bT5/hjNCTuKveFCrd
GWrgNhwM0+BbcvxEyfMCQFWpKfzj7oB12yO2F7x7G2YdipZ+6IglGgxhbHBOor/xFHBS/LGoFWJ3
u6yZyX+EM7WBP8gZlFk1pdo9GB8K/KbKafNZ9uYmXqPZR+vZ5KzVCbhh4uCnE4DSVbiRiV26euza
8Ed4htOm2tQu3/TiOrf0q8XkNXWN7390jW4JOAaDLBfiCZUypXWJU3R1lMB1nvkTj4CmEGFeAAkF
mBE9A1NdGRaqXLWoSGZieN3gbHjE5IVjQABgOP3eOGN5m/L6HPO5Ol4m/mXwXcVgKgj3KeEoFM/x
k8wEMm9SogrSRf/KtQdt+Dp26IymYPCMCNKUSLU+mPsvt8UJhO9Z2q8skXZb7YndYl7uRoXjc+1N
vGr+zsutzxlV+Y+IeqQyaU77qNj16BxzZtEUz5hxb111hP0XeWXiP9maYMTEtpXW2xxjWKmLl8EE
if7eXpGwV3XBvvhdb08ssl4lFVkNlQZVjcCRRMxeuYN1GC54TuhA0dNhX5w3chrgtUNy0rKn1JIB
91mPjiAti/mQO8eOESncxtvNxbLy7sy3yinZ/EBNJxg1agCNEMRNFRyAgm1ZqezLDFqvLs508yoN
laegYNOXCFoUNv1PzvqW81YSUlY/PBrGnwbmTC06joraW68rOmiV+URnyUzZZCxurhrJ5KBeBS4Y
mm2mFHxQzlMBEZm7/74AX6yCm/4VARyGq9CMLUH/9oYJdrvgJEovf83yF7L5wBLlnvpycYRYhX4w
NFOD2OkTD5oEjPFjPJwX6Lfni9ExPIqwSQBjGjGxlMnHKpGtVxblV14f1P7+S2TWfbHUOMBTQRta
15Bw1hStVUKG3irP0OP2jEeahgtaUbhTNnChzN77GjCErceHcFh9IziCYxQd/64uVMLU3B6JFu/D
eiOC0v4Tah+A4bNcstbjlF65Ji5MhjhImdezCVjmupAYclNaqv+VUVBBhtbNRv2AnZ8JnbWW/4eH
yQkY7lz2u7W6w/x/+S0K2dGUwkus0KDrZ49N1hDaeakKhkZAxvXu0wHrXlbqrxB1QXighRpfPQCG
X74C7jJ6iEKMp5alos8jqROLnysbFoHuCRevMBux+o9z4XtV4Gvx3B0qxzAsoXEGBWATsSeYpHqO
aNTf6USTA5vdOSy4Oe3D29YyIP3UljY4NoW+H8N3wM25D0Oi4JohU7t9Fl3jj5xkb4pcNMXpqCL5
xQ45Rzxp1eCkHCmhrauKSx+bakZ98Ph7DYnhwFuWXp/Oe2nAxyU5BI0GIyKBd8OBuMF4RWiQAzdP
wXENp36KdGr5CF/TjXOIbcwpxA4x5aCxgemFjExuMVqoC6aTZ5ejspk+gzGCtLvvsTwOAHOal8B3
uR+Ed/97LggBBnhgmtOgde0ake53bBXhZ3motdl90CYtG9suXWklT4LtzEHFz3pyfYYWuSLYyh9k
oHIH7x5ihvGMTcBDb19bS+AXSUWw7LoTQ5UQqn6pp8NXk4x+NkZhoZzSNyjFsapxBdjavLpwlsYX
jLD6hkRGWu337gh6M2ArEu2Uqnsb0up4ijvUjDMWRlHUeItyD6DoDBVI0xsi5YrFn8r7vxlRNi5l
fsK0T+hkhC2NMTlqOx9je+d1rXgo3Dy6DBdvrciq9F54WtQthDCySlyGXJvdrTMWsZdUpX0i++qv
ZLFqSV5kS2/AIB5YLKU5WVWSaWoegxgigJ4n/iz0hZb33O3SQCJjtU3RZxN0EveWQSgaFXo4GKYe
S6DztJkdiNPfPhJ/QY8keK7aVIGFobjDYTxg5xbhZE01aKjSzrvCagKTMw/V/hpcvJ4QrxteQy/Q
hpuj86Xm+4SKXUWwxWtfW9kvrwEfAI5z9vXwIhipCUNvtYsa8yGDLiaIW2gWe+01mXehJNuaa9/J
tQbnZFZClRPOJA2JJmWvr8eCpzNmXg9tidt4Ar5CjLJmJ1imoahn+q/HUq8qrJmVUqOoLxk/nzz6
ug+uiCDF+TypwlAEaDGeLTQkYhrXPCQT8eXden/C0EzIO2KZoy2bdhHQWaScRkkMtMYtimBz1+p4
cFiUFEXtsJTRb3Pbw834YKXRTZGEchdcyhqrq4TqVMxPP3mEHRFA8EErOFy6P9UW0qC3xc9xYfzv
dY/AnaDKrIR//+G8TMvBCDm0N/HjqewPSfxiwFXAwsPXvvpuGQQfaP19oDXb+R15ba3NoHJcU7Z7
hLtU+rmHUTZqx7fLkESrp8+fF9MsS5+PxIetJGCn+vfvfHKi1fTOgDhzhem56SJ2u5WUOx6gtzkZ
yLsQ6q3vNhnQZZ1HWNYBOpoQhlnFF4que7ScxTCkxUzKb5tSuBwYzYcnC9/a/7O1MRfp6+fXI6Mk
3E60GPyGd0teB8dT74sSqb7CDyTMchiZjkrNZwbNUkmDJxw29i0jFV4Eqx9+sh+ThZSQr2S4LKAD
tlSlf2+w5Hkwu0K7GYVqUEpKSBnMH2nPF1lskg42ftij5po8uv/PHqXQVzpadvQN1i6haYxyHKde
EeunTmwA6cN95+0bei2K3tuMekAtk7jg91WI4Bcdoa9n6xzIp2WO33E0msWyd0GepkfFdROE+OxD
2UW236sw4Uz9lx5AwdQ3duwy07YcjlSvyIpADsiw339f5I9sDMntIg2VWAppNRfmZW+Nnem66YNv
jzLpqYzw4ZCTjzMwr8AxqCV2cNMrW2M/F3jTLjNDlpPryMf2TR1JANwjxkXayPBDEtEwcXpXCKZW
zdfeqiX4IK10Yk5HUbYPcQnOlawIgb/wfg5WGKELim4TsXHdianWZD35gjn9hmT+RMTfGMJZ82Kt
jLqHRZJl+DvFXbnWoCsODwgANbXASg7zwZkBBYCfjLzH5mC8La7F59FyCjvuy2NHAzZzSkvPcUV6
QEmCX/cmDfmjztx0Sx7W+HloKSYNpDRsBpTZdPAhQBL6Vtg39foEOFOKQQ5s9XXCroSyfaV3a731
W05swfIchXKB7OkB3PDfJ5EbYDC5YEgGeCPnHNRBODeGDGuUpW72jmC7Uhu2RjYCQh6LzfX+Lzuz
Y/ISt12e6NLIxNPH2f+NA3gBxQsJ5BUiB7i/g/8KTbv1n1WG1dCXawFE1P05eb+iyuGZ55gx62ED
ckGOVjk3+JUZICgQFgosyyGv+zcdL9D4J/bwzXXixDnyy6EJe176F4nGqNXjL9H98N1UFOPArYxf
SeWXp1UKcfQmupUpXcRd7fOqsdeY3/Wvsrbp3qigLn8wC0DymfEL+zr+Y1wyQTfdWI7nIqQBoDxF
aFGtXPfJ0tIO5cfcRGXx6Z/jYCeKPGlZ79rYP/Zyj+qx25353ZcpKejMJBe/hCgsdFERNRXyxr/y
m60txvcjszlWXLB3VvuflmGEcKgHKZKZCufMITK5PKLMF3FIGncYDqsB3w2vtW7Ju5QRC0UtKPPS
rWGoIts4DbuQ9rsz0fvon53bMnOiSAI5WpF5InTh+S6X9o33TvdZ4eR4jQaD7oTY8kgAbMl19VMf
Wq3hip4eoZV5MiLqez8LJcu8/07fOCOKV1byxRrkzx6czKwNJ5vqdk7brDXzkQzwagiZRBTQWHXI
AsXFRsBmc/RFAePomtbJpu2ndiGlcntMDWSAUeD+w8UIjfhE5lSry3z9Xd0ztkxhZVqtJd2BzSSG
9zp17yrN5SLrzaMCt8xrLyUI6OOmkM7MqJu0n/L4cfHAExZW3Vb8CiCk4HQAhROa1Dl9P2iPwyKf
ahUbnh8SiXmVazGEKrIx2NX12dBON45yE92CeFFANZVymP7jo/9g37/P+bQ+9MEJP84dZpVgQgy7
vSWXCSEiphlSiINQBW1rqW5UpV/uil7Gz8IVQtFCIb+Ee1rvkegCLiYT/yBW06rOUQeKcvzG1Tv7
6UBvPhLK35jX3E+cM1YNkYVWz8ZbnSqf2y5Nu9RpuOwJfLWgCiS0Uze9eQ8V0IP6sTfXDF9sQeo7
qxM3HNYOnK6+iV8H7gMhrgVN6TZHdqacjYSywIX1JEfl1S/TSN16x61Z2i/m4nD6fp6H85g4IlKF
aLM2/l3hocrE/qnyJSitEJ7nGEwHzkFjPTweZZb7fUC2jN++P3x8UpQc6d3MfzrxIncRDYR9Yn7k
cwF1dYegV7GBRPgSDEyTbQIFwbVdiOZsB+XI+R72d4DoWeG4GWK7UidIqNu3BW6VbGtr+nqVi1sG
lH0fTd1Qfyc6ZQZXs2fMtf4hHAjYDo1UWPn1Cy7hDucUia3bAweWAz0rZEHpZSL/AIvrpFzBXv8s
rbmCutngpsZWjYlls6fMe54gnNdvwPxAxRWKmHtA2ZqFRfiNmTwkg9xirmCmLHJ5lEv0IzRYQk/T
MPXwKNuACt2jcyZk4BrlZsApE+pA7nQGL0AtcbaR04NlG948yC6+T6OgobY2a0F8/ZM4QAhRuHnY
NDn4RS6cLzg/A2hdRjIDIVe5Ymk8BYYHwVZDSYtWXX5i+QUooMzOHn6b6Vh3A03zfADO7D5ssAw3
aiTiMl2ugEeW28p9Ko2k6BRYg+JeLxRTeFSfTAeDuX73zNnBUtrmL7hOPwM38P5PtPiNXTH+v9n+
SN64A1WBN4QgcDxnda7qIzQw5F5V4t0zJjHXQgwbIvN2CmSUH5LrBe0l4G/lk7ApkJsqLqaFSrzu
hRFbZU9qqBdJujHrLOIy8ceFjRcuacj9D7+2KVPIZEqXJxzCqDlvTZAt4tLCDFdtMZe+DRX85oom
pH3JydCIotRkgMEXhWmZ86vh9DCODqjXlP03j5pEGwpNlppPWFtZ0y5y0AAhOvL+iHT74fykzlA6
sGQSqRbfYXTKJMV6yAqQCSJdSrKaV6zo9GY42e55V/KAOJfpYodSpxzI8ninc7W8i82vDsGLnL//
ISVirsbX0Pf7pIN0XpTnfssTKHlPS8WC+1Z5tuiWp0qqvqr0e4mIAcuzpGVFw3zgBGs9LQ5ISm4K
KGZHnvvUR5gPHjkN/Py5JyX1ckScrAPmkkPNFd45nYfZjSoIhWXuGevbRw+B194w0Bntqlz1nvqe
oYDxvR3jcVNCRGnCtmLt8itmLXNWp6D3uH8YZlZg6Tp3ofuGChMwmGCCtYnPxC/+lS83j+O3a7p/
nt+itD41k8RqDwjzYFR896Yx5+qosP4ptXOjbNtJ1jOtEN1VmOYY9aoaREajMYbf4dbX2FYrCLFk
zooMRXI8q6ItbhtskmEkWksWkDQUpqNqMkcw9U+64jRj8dqlWC0ZVEfQd/WHNKHVCHpRjUv6b6HU
opnNlQt7/XhS71OhmBTkxAGuMzXv0Pk4X0Dr1FMp016/hNk6gihn9RIwsbLD1LbOkGERQk41vDd0
c3UOUgn8s0zw26sRXXiniD1sRtkY0W/spKAwbz1V46njyGfUQ6sUkQCsJDJCPQbVANG6JXi9Tb/c
f/uO7RHlezw9LV9jwvBEqL2TjfTotLOVFr32xD2aAw17XrFEJrZYdBeEHQAadZEGpWd1HKEtW607
WjDXTUjtHG2xPiF8gjTJHxsYaQ28cPCIRLLCYBhqpZNlbteU1qiEUQYijHggWgn8YzWAcJSCVvpA
P8vqHyJn4SPHbfZqp6JeB+6dVr9RtL5DOM7hAJ9HV9mfsTZJ1FVO9QVx5BEYIY26WqmwNXiaGVLP
hykh+m5ntcnA9qGu3bFdq7XvX+ETyR4kIm8BT5tgLA6Ydr/R+Km+3fsq1y/XG958gw8Snv6oX8Be
ZNoDI3Hd1h0AByWLnKTNY17cvumfAP8uIJqA1DIKC+/r6NxjLDpyhmUV+D9zc8ozQAcM0hj8G4Xd
zOi+IvvHfjHZK6diPGTFErEf0ZwJGZK6SjdmWgLsHvuCd6h5/E2C15evtE9oTzUS5Qby0xmrJMjz
5+9UOYnkyVoYj9xHz+0DRZzJ47NHvN8VBfeX1s1N4VFE23Ax2pIf+jODHxyG/vk5/M20jyBKm67c
I6QzkBJAEBqrqnsuE/C0PtEP6PtFpbxPyhFgh+sv7jXY3OfjcUtUObzBI9f2ZMemRhZ57nnLGYR+
dBxNyilpYq9qyY0fZG+y/P7ct+dqxETgmx4inomXm3yAO5q8iXibU6XCjJ77AbU2yqGVHsthMNdT
SaYr4kKxB7I402PCFQYZhDFdxMEefty7g9EEBJEvXXGEBJhWEjfVGghPCDH2lKsSh3kGrK10B4BS
gSkVpjGVmRLWQhMxh7e+TZUkfgylylT3fhjGErst11u23R1m8kgrAg9OdUgf8UWllldIiHpk6VCN
YVBDs64tFhq+gGRLcNBtSF9fhIK/B9/663YXejCyWjNDzw0Gr7sfz59DymPoZRE6ig5YmMoz8Z8z
giwLp5Q6DMmHAe2NHKQ8pe1VWPWuTNzJJcLlz1WuZH0PDqmzHQkBrDIr7WW7D5Z+9JM+EuakT46a
NmpU1b6wnxMlxsFrk7a6lhKaMu3oR3wuguQcx+j66myBql7Ta52mwLE919zEr5uR6u/6E49o1Acy
KAZxr6MDDtViZ1fm1sxL9wUmXtCQsshUWUVa84f3F2+g7KOovYhPNUcQR4CaeKSBch1E7NBtZMAb
1hQyIyz++NF6Jwy2MVahgQznyp1B5YTHMuL/Cm0mj2RCW2AoNXBrqqMNIXHUGzEvy6Bhpm3xadwH
knrWMzqA9NUaP9/cGdvfbKes6MzaLk+oAjZ3rlwMWfqo+h2uHZCawIGvOy8jK8b5xwmpLd+L6j0G
XMK+bHGTyKMGiqMWMS6g1KPsgGivQELi24x8JZlcvvOvYXYki3glCMFmDB0OMSBEhj8z6Ox5NTgV
ODo/fIRMwzViB2NkpHCE4kESNexzjgfImNgboO5De+ZYvWtD0HjKRsSQNAj51tJRmM96eEiBvu/n
kujxEcmuRbjSx7UxpUQKJKMp9R2Q5FqujySvZ8jqnmDgRSKlq8sRktJc9/dBXrMUDvpcKzJYqwXr
F8T32N7bAgwALvzDmWLOTpAFlwBw5OKEf/ugWg4ZVi6OFGryzNTK0w9MCTwIuT+I0szokjwoSYbN
0G6n7s9UUhKzOLRTxjOlM4jYy0w4vDXDOrQABi4hpDN3pRAfa0NU3megkQhuH7kOJ+wh7oJzZJ3S
zZF2kQBSgZjzdZRefpdLCO3VXZpP4QqkPdD8iRfwZeGRQR5I9Ec5leDwq59YsEM6UfFJaZLECsMr
yIm/NCt06r4aUe1LxxUvUhKiRwG2ccyQLBgDI+qUiPDUAAiVWsYu3RflNogh7d8U5+wDcg1fo47j
jCuwN4LVB5JxnBVJU15dEy0EuDboEXpHpc9kpDo5OPBFbKKYUln/kjTwlcJsOXIff0yD6IMlBoma
AUGoUJp5/HLMqeOpULV5JytoGA1jI4HAdFzt/v8gX1B9B5Oue8taGeTVNbAo+iv+r7i9WotlZLr3
RXF+i6Z5D4K9dyogoQ6IBM+5l4xSWigmwlX/MB+phNbdopybh2h3FGnZ6TlmK4sHct6phZE37pfc
Yj7IcWrx1HoMFWRXR0ctI6nGJacLhg3iOj+ln4Nsvii4oNQHFVhIIDBelfErg4ed6Dl2eek6jLAa
pPoqb6GkfwWdFN8EahIXF68q/njys/g0cczem5vUaqkVNXa9inHH3eOiXN7mT58OZsYv3HwEMpIZ
dezSLW5m9WVqdYPG+RaQf2tqpT2tU5UvAPfA6d4e/vxia3uoyXPRXmK+uKtFjx1cyH5tC4I3HFcL
az/Z87iftCYGy3pWxYcctCaaEQGRKrm6PFes2fUqLgb02MOyduz/J67eepitOV833S+ZBRDbExzU
zuDd4uR3UvK7Flwb20ZSsfk5Eez5BRT8RaSZY1TOwCzCKDuA/xkEYVXMgnHY+KfOyW5c19ptI4zu
L496FzwoQkDJq3MYOuO/LZWYCLrpp7tKlzK/peSw3nfdop2aU5m+fCQrbVItzq1Gx0H28WMhr9Uk
gTU6QakbA4qEE2vNtAkvOJ5pTgzCTZpVxhk8pBo6lH2jxyEO3Ad+yZ9QmNYXl6fU/VTOXN4QXfvZ
9pe34gnBOxsGqH8jCqOkr2q46Tfn6egrNQsNKlLSwUfz7k6MA/V4muOYjYtruhg1RiQ8HGlmvEJJ
dMWTzEUSFQKOyV/BnhYCRWmdNjf7SMB8djwJ7XrIhJaBHj6KmoSVmyGG9VJ6RKHJy6sVNZMlfCuy
TtRiFv6X/2tW/9EgyGUudCe6mfBKr6H3We7LTbROJgo/+pd0JtjBDyFthp4rZMzdSnfsO9daiy5E
/e6eopy7qmIhGwgZcwV8afcApM2oPpJVRFPWXDMIjo7QHLtbCY4n7tpuQX5xV0Ci8PAk90gfP55R
n+zzI0m1MRiyZ/LwteTnTXL2PKGo8VkYABqANLBL9uTFtRHPa103ZEdJV71yp4UsUySF1KsUq3Xn
So49LfN0h+G3Z5ms0a3a38TxV1b2kP/kC0l6Z2+XctDaxOBv+wLJzyz20XC6qCnjXWtHmjzTef9d
D+JB2H8qLxhNb2bUnlbF+uX/vRJb6VXYID6YVYDf2IvyNxp5NwyRfrBjC+9iwUTG1bk13s+vp9i5
zkMI7Rg4lCKKNXR1WgWAazxw6rQjvXyCmDWNZEPCoopkNSw+lZzNBn9wmO/9Y3bD4Qrra+52yaXs
oe/nf+P9b1KepGaGs6vHbX/smTt0H4TTVY7D2x2LYDtCx4X8uj8yTkEP1xb6lhtqdKLnNXrMmeKY
eb/1e+lWgIKRlsGKjU927pFxlAopFU1RW9Qhh6z/ZkoWbFJe9xvoRrDSk4IpDcwPLwIPOChnX/9z
5x6JFJTbOiuW/vNO+m9fL7CzNWNzkSGWZurFgp1xC5u5RRiglUsXjtU0hpxJN0ZWPJf/zoEqqrBb
gCPrgqTTXIpxJUwFJ6gVBnfv085VZh55BlIIq/U1uQH+8YcTwoi0NFgwt9Sol1T+V0KkYQlf8OCo
LcQNxqexIxl2aWqzMubhWdSdJQR87+B2R9rnFpSYPBqiTeWXvjOaFjziFdGAhnpUqv8tlMqyxols
iwcOov3PWxmt8wfjUTw9B80QDDkhSR7gHENcLl90di3vCJrpyqYi3deU5vC9j5xa4WsWQF0urI4m
/Xs5JeQzo8Lpdl4vrwqA8sk/DkMbTq+Nxb5a3pViHltsrnoN9U86W1TQXc4WrFqqi5SsKqTJYR5+
LVMYQubj3Yvm/x6B4psXtluWhDWUyXkEonpZ9hDoZx3Fd/CpUn6JAFfPSRfk9lO72dqvN8e1pGsj
LlH3OPvT50qyZeNg6qCdK6OQFfdqH/nTTUjdfRaiqrlUPFQCHCBZWZ3xZ4k4L32WbessBTaTqCx/
V4N0RohVFXPIVuVatifCBGuycRV381CZ40Xv89rJ9i7NepWPPYx1FQ8ZGxYPKGbe5Tk8b6+Eq/LD
rIHFiWDqM/breo4hlFHdb+KTEjtTsIAetJNAm5DKgCnSvMtAmGfiSyt/VDq34EA/JZ4Ww9uv6Y+b
FwDAWbnCZCXxXqyMztbSFDI3+j/ZguFzAYNzzhGTsA05D82EYEGrsWFEBPa8+HQAWDb2R1MrBho3
kPmXWafOBFtMSZ3fAckXGd7X85GDwM7DeKEIWZxiFd498nPTB5DxbTO5J7HIOgCKHSkLkoVNWiYL
1DsRlgPHnzh+XkBRBB8OSFlMXxJdamqin6fEoIXPlY1f7i7i5RYLBfJOa9vDZuOSbn1vHpx8vvS1
moGV0nq27gytzcv9dHaYuhJh8XXDjhPBLUbePkySFLa9Yj3uF39Y34eNOKjPGAWkbdzbkk3izdwi
R1Bqg/G0cRyy7zCxFUVCES7gQmDfDyJIQhlLFLTQcIEScMJle+71V4jEqhhC3cm/n1yqj3PAVNas
LNdcHEkCgNjKHPdeKhYqqFIwVkMDH1XDB8EZ6cN/JX0RC4uvcvn8/xpVJncXzmfHWgHyGkUTecxE
EkL4i6Sg0/UzDnwv8sbTpDP9S++G7rvu4Jz2rSaoQr3vJIf5oMf19waSVgu4UeSJL38IJ0orloYC
KYblTaqle4ThA6DE8F3CX9qpK2iBIcEQEa/YAJfr2/fDkZ9PVlR4GtxbG355W1WU8aAaMwf5/Exe
3AZLbR9qea8XWGneLPaPofSvsfPKQr7WnZDqBOCGbnyxW/L/rSPn07qXJUeMZvOliSGc9ef2egG4
Eo0XVxq1b6813zf9thWitAfyVQkHsY2S5EeFWhJItaVc+i+Ipc3NHgnbrhJsBdU8avlS2a9TEbD7
P8IPB0Xp/3BBlOv3nfu7QS8JApaFCCibpPe1utkKkJtSKcQbqh0661i9w3QOL0k11UmG3HRjX0+j
7DHb5nt3MhpBlRZD+ywb+qgEL1Mclt+9Iyt74V9fr0IEYcWXtTrycCw80uP0MSijACBhOqJyelQi
1uda1cTSkfgm0UTC0jo8hWdIL7mblkosWuz8XsSExQqxWQ3LuwC8gMdgJ1rfdL+FmKpoofxl3x/2
ZsEOYP8RxZIqnHozRxH5JGVfQ9807d42m8GmAe/2C7tZZuRhmSSXcWLLLCanmt3qnKR8i6ons2gh
g3rkeOXVedCuYGHEmSqBkkPYN97Fbxt1ivEza0P9DFZER1PJxnL8jSxYbzuBukOjQtcNUupGR7QN
ZNP6ieW90ABKhZPiGsvXIp050QX1jpw7SB2QiRuo9RF4qXNNsByQvnwVldr7gtf1UQ/kdCdV0DXs
sDCW+7ZKV31a2JjT+TeFx3tIP1Z6C4xf0K1+Dp9Z7KuyoTEgnihaBFU8Hp2rDm4VhwGCo8c8pqEJ
joTwvnqhLzQ+tSFDAOSqTY6/FpiXn/7qOTJcJ0URhlcC8gsL3BAXf9wu3lzKE4QAakNqq737ll7e
hSLUoTdux/O9kH62vyQvjBwkRRwDpm1hDU5y0lFJGfn03YRNq1N60Um8/tzUzFHtopCDdRp9LHb8
zlwVNDTwxfodSefBhVdtI+2tSHbOWEs0sCy3PIggSWYDvanO7ZnQso1vYQ61nMfpcdlUzuqKynWg
OTUJK+s/gDebPyw4mtskBSE/mA0gbPH7UTHg2ULoByudipROE3Zw3byUNNUns4d5AAT4uKWiWHt7
2kmYevx4sDJ5EsySsDAlIZ9Er/3o0+8SHU1i78+BYy9EsQDulnd+d8c4k4TFVCc9Mq7zalDQQKju
Lo8pwwiBLowVIjtxya7LAHpsAPunl/gryuPnvcDG+WJ5BCiYcLUhK/gBZIrOpFq2n1iH/nwP5N2R
ymBp3hm5y+DDxS8X0BUt2R2zrRCbuEsRUI7xvKR1n7Ps7CmBP/Dw2YBzM6YThd28HEoKhFENNIjJ
p6ZNwMV6q2JMWoI7d4a8lqOYs8BUyxW+mLOKZmyRPTn8rIKJhq4LeRsHHQb7DCbFHCrco97RYdWf
Tga6z84gQ86iavbyK5Nq+BDpAypUpxnvfurSDhGiVqLKkiWUppZocl1qOzFpoNQsjNgOGhXZLi/u
eTO2tkcf4vJYIiQdyt9RUm9J0IW+sI9TbQqWcFi/fyKQqM+vySw8TP5pKWezal+LujaHsI4vxdJm
b07n+E3XAu9AL2Myu2qe9FPivFQvdt8oO+THLLSDWaPvEScHHJVngXIndCtOGAxii8FtF/wKN80Q
iYgoAAOiS6wMWhSSbPj+BHeb0Ydw4sQKfxaVF5aaCPrqOgJpb13iROCWfmLppEWEdfsQjAlVzygR
N8sLioHMqUYQGJgAJq0BkFXL+Yzyz3rbXLaLL1loB3SgjLMdczffOBbzN2wsKkNGBKSsS/2IlFWu
6pwOeAlYV25rdqiCIircFE3Mv/yGnlvHPt2IBEf7NWgyM2F+e5ftadd2o4OnNmIn3H7UBD4ag+JT
Ram3OV9yEl4J9qC9Ss9gmv6qpvOc/PVl90NRF4oaDJGoYJy34tZEF64/K1zlFz4LTR0jQ3cr1WiI
6w17U/eSqa81TfdCVWgFtAL5tbTgaSeqxjmAK+m5YngZIIPZEidl/Ipt59hG1ecwyWKrvO4qHplI
bSCtGnSQmX45XGD32G1MfM0NZOetW9eFLSUJpiBTk9wLSkZYjTIVMkaRvwEJIiM82csufIVGpZib
UsGwSQ7UtiIqxhOodEZxboR/eGEmLGolsLpdJ+TD73cTIUvWRMdr7fC+pe7N5RebIN3YN5psifrj
bQQibdmvH7KLZdnaze9Z5UAt+VJfExaqQ3ipa7XcM59lkFOTkfuwGjgmF5xWggnQQATJVYmpFsCc
VmxsSLaYAnJXK/k6TAavLty9vCxYPF4zp1vP/HI5MSLXLXeS4WDr1t+UvzpT1aZBvk2pXbQx0K4d
sI7ukfV93B9AfDUboLG7NGJEVM8ddzes6ZnvJBy5w/Nsqi120hou+l/kdeAn9+e/7P1a77EBqR1y
jFwTpPiwkHxoHsHRTwpEsXoVIoP0FURKmKJbIk1T7sQuEYWcfQIWDgVTtCuDlEGsgVYkgqFaJBb7
YtC4WNqKphNGsmDWDDvpJEcn7/K5LnTQ2f6UORgyefDYO5k2JM4qs6f4zO/7CiJd+PdZyuawq5qg
KdVj3mdFmwZPjM/zJONJ9xHY6+LkqYmFyEPTa8NSqDgiR3jInzermpan2LS2H/JWF50hMbtJ/Mc1
C0rzllIXVzUvBhDvxKetE+L1gTy7D2qL/GL5UaVPyjs3VSWu4iu8tuanugUGOX6+8yLO3ij8qgDl
rdLNmj2r6GY1UlPANtCnAM57t+fZ4VEBgEowflRCbtJuEeJScvetIv4ijEm8VQN0OwW2hEGYDRI9
F1V/3Ki+fbeAxDDvMagg8RGkXnnFTsOJx4Z2Nt+bonUsPjAqc5eW3aPWS5kDlvTuajGBryMa0LYW
8/PjIVEbdBRyK+RPEsaqOE27UR/rqS+yM6x8ndk6qc4gSUgYLmDyR9kp/eKs+/2eOxQShEqUHjpd
mTWr1nNcajdRmRhlHgrGTRY250zQLLKupiVJzUCvufLO483Ef+ZabpjJBv8ph86yk0LnziS2+SlF
z1rq6X6sN2PxVnnRH7v94Py+sDcFh40yebkzjXXIIUIFewNhuzXJDKaExNrhuykoVp57NpfLKGF9
bHG/cjn+sOMOQEsrRV9aNV+jRhcjZupil5g7MzDJj7WpYMuSZod9jIEe8nXAW4/PmNWFE0D0/kqu
mwfvxV1vz+0syPWZHxNA8p7Vc8WuicATofl5P3eDMzhaZiQU75br4B+VoRHkenruTJZAKRaG8JuM
SFaRmKpoFeZNMPURCE0yKxZnHaOrDwh6Ghwr9x7baohFPm6VU0OXSePT0SpE+Fo8wcsfWWPrPJHW
a1+V3BUfSJ4GTJUc3GRHcRB5luZGSqt4aowCgsYMGZKxN+yjuDEi8QNcN7Mmefp1FyVyvmYdOODa
jHoyS24/y1DgVkq4RwrvQ/2grCGdlp3lmRI7ZjROcNiEB6IBgfOsYOo49U8sqnn/Kk5AT7P/thQK
HOG1ZYbE6bntiprmdom7M5g11cWwsPbBSHrNUjN6X5VhNXG8/8i5JOdsEEQATeGm2olzdgxq7+kj
wBdTgzzBDfYOObKydAdxspoZgBWpZ1zyMdVpNdWiw9QyL9v8gq2lfhslH/ZfK/i2NiAj1MM43DzK
tu5d1g8SW4avIYprMxt2SeMqZTgLL+gE1Vv5VliGT2id3w0UauwSCyPIq6ZeApADMdyaF6qe9BUO
KxU3b1bNfJEc1WoSVFih8EEHg9bVN8NqEgy5DgvcNmMf0EAHlrzwXl4nR0sPiyxJk55OBNFkCxey
jsvuwQ/jUbSBEQ2S45hxWPqRQHUFLyx3+D8W1iVswub2t6ONe8sUD6fdxuhOrIlieREpj8FZeuKk
xcWi2eFpl3YiomkIWXqmB6N4RgSRBlrhVkO8toVjDq2t41un34qXi9G5vkEaLcFsEO8Yyag4GFnx
j8Vxe99oE0PCo2zbrUfIbjb03FoYAQA0zggHTLYP4Hj6QXJdtAqYxDmsOrXIXHvzGajTPpPnK8Cv
VqOoytS3QY96WOXuf85AH5E83gONcxcWPNnHUb34fKS55r0NrCEyKNCNNRrTuLHhdOJlMN4WKvZq
DAXwb4RhhVYHaQlYdGUen8FzJw9Ab4Cfnwcqk7fqGdNnUQ7aJsCyIMPB/x0qscf5LJaBCQQKJpiN
krMRSwQygxHAf5X0oCbbZ/paH3/jbD3ySwKelsJOpvgjuzNKAYg7VxEUFJhHY0RIh41caZi4hQSH
3+87wksJJWyV7pQS4atbu/S7XNxQ6rzPsmZvfvfsN3K4frh3CnSGVsWwuqZqBvT7abAxANa8hdXR
XTP5iRInU8nYuG9cxKp1cP5PtAOURC9CXzZuCjDmxjK+HPk6QAQeDBP7LRwASTL9pFJAK1nhYfst
qzuONCT5BOY7HwNAX4JAkO77X7tNKaXJyRWgqLFm9BEhs7LHNy1PT2o0kz5gw5tB2HB3Lzusg2tw
gUa+xRYg1gS2e3HZWXp/lnrwmOqpa3maOpb1/KepWeGoQmj5ysS8J+Hmz2shGrdk4zlgcaVWym+T
bdyYWFfKPZ+7a4ti9HILCMc2PUI8ceXq5p6xs8FjHxyV7R1pFyQCvqsMa+WAvhxY2O6ufx9d3NGg
mW2tXTEKdAkzk+u7zj6zfpLL1x0sOR3FdjK69FSFaGH9Sm2ha2f4PsOkbKpdwtSxRUj5djxlvO0x
K8CwkYNTPzBzECMT1tFzpCtCpsyqpgJg+fq3vDQ8W6lgKSyO5gNN5kCJVjUcbmmD0s2Jlp6rGJCv
J9h7EblDrIVZkyuuejF1GJQY7vC9X1E/F2COhSX+llnIXpDe2AWfhd0lbHdivilhTv1ebO/kdJNt
KWb2wEYGTghGTYIZSsNg48QAEXU5T1q9EPZ1Fr396QPruQuqBrrH8i8CPoG9U2c/wvFCoj8qisSf
lQwts3ROV/rTCVPvY4zMgg74lcr49Zl2HtRi8vE8f479fTjOJbnr55gKzpz0epTjSEF5vBNbnv0N
4DM+BX54BViSw8Ad/A1zvdVex6jgiT66WvQhkfe/vnhPAya82nlq8V/K6S+Ls9uIq5/dDiAl10nO
CGF5pa3rB3CLy2xI8OSvnLoUA6GjDt+/nNkoFonrH8Z0zkceMq5PyH0j36FLzHL+oTQtd5hj/xJh
h00Arv4ZHrYzMIn3zFVIGHZPE7nSM0MO+k3vOIfr9c1KDtNRh56Ax6r6r0fFjbMiliM5wUX0s7sx
bMCYcdCV/ey1pjGb1th7fpKE44iPRNikUlFy8KsBO+emzATVL2Les67qz88hTGZHVuJINChG/0tW
E3Edif7pHmZwgt/8Iyih/jACzox7irMTSYbJjuf6ZXFYXvpIx9oluMx4fdKZIFNA0lxZjd1NJEgP
ZuRrlDY+0XXSc9EjI8lOhCRjcOa1ph5QQ4WmwTsP7RMequgRaSjfwZBDJtBIVvirA61stAB9gjvz
KDKo+EFPSZRSfZgnrLDvLN58MY12mPuweTTnZsoclw0gEhipN55cDklygbgPQV5RxUhflmQaas5c
f7RlWNZiaYx8q2j07lWqwjzy5yW7y0daOLWpk+xuLsjS3CNt9W6bDkkHimmzn/SLiVMn2M3SDp+S
g5QGi54DRQS1yrmewIX3WltX//QWV32wDGGrFpYXuCPLCmD5ewUO2dKmXYTGvo2HsQdG4Z2sSAX5
QIiSJsV+Rcy7mWft0Co6QdRnfIdX5M81OWrdwZV8qke7SrOuZVDWnRo0aM6+4vKXqRIuTQ6TuuMw
uL4ogERJc/yL2E1kVimnuD01JPoNNPIVEG3LgTTPkPrnVxe2H3x5QpvE3IRF89JWArg/TeM54tUY
1PKaILH04yco0RumCmremxv7q+sR44GKQSbuGhyU1RU8ThxcgXRVtoba7z2B6iGZSG8r5ulSkQCL
W1byc8igH4kSR6f2X9HCTQ62eQeqjNLAqOrTLyjthP6FjGV9nxUdUIBKIHF3biYFC/R88RNnqqmQ
mIdy92NuizHrM2XowHBkgbLVELIcKS8h4zMcS9h2zyt4QxCSAnr5rLrezMHlg+U4ObiXRcRN4eCR
vrhQKclLT7t7/0oqLOoyAAc9XyX0ENlZCed2/svzmwrDxw1X38KrlZ6g0M/Ly+/GPPfzJhww3Sk6
babh55qP30g9CZ8Hnx/AgNgv7tyWX8owdBWV7PDSsCoR8oaNb+TjKFcbvYFjNLteM73bMNnVSlEH
hU2ihk2PbQ0n20BKlQO/acAU3Bw8j+BhRmYqUopSyd7QCVn2jFfrF6E73MrfDKB0xjpoUFVyuXDy
TJsptppHCM0BAenm8+R711KCecJvzw5qqi2tP8rXNwsUA4joGwczes8cW57x9kFjc6Ji9TJgFstX
Dit37VzPWCFrGOVw8gAtTom6hP7ggry+D6STYXyFAvePfNYwhjyA/PE9Cl3xicH62OGIF5YfyBeV
9BDu5RkSyVsAfsxJHoNI8pyP11z206DzM2SRQtPnzJE48EFS/mc5TtxHn9qcIOCVAl9kjUr9qEVd
lfmHDtsCSwKF7JmlLImebVulaMozKXeUMqu3b4NDeYY2yhV27vKJpDAGVUiHkDdILYDCyd9uYKS6
LIHezyS746JLL271XSMOkUNs1VSyoihP224QGZPHPX2y6ugYMHcyQRGxi+ZcKoHclFAkM8ROQ+4I
vsW9dylx2itn4xQj+pPypeKMKOjtpNoXRhuWT3z/f6MHHCedLOPX/iu4atVhhzssu9RLWY5tHcQ8
Xx+5v1cAxGu8a5Uh2ELw2zgzRHW4SkBHfgfq/jp5Sp4VAXQbf8CmGOc1uY1vxps3fUwTmW5vWvtL
nfmspfTULRNIwvbQTXJDD5vt85/7LXwvaEbbY/HsgchBsYTJ8OjxeRjq9XrwK6IQSZUYxey1mgbI
tksu7A6NyRa6GEiu0wGKizuZ3FyndGCrM5nTTK85tblVjD5qA7JQGbaQc7mJfPKBAwDW41BUl6/x
u57MQMRd7VDkeKLBSxP9PjZN2yOsrwVBTaphzuH075MtwhTsxDuK59YfYPv3b27ILrsauyiSjykU
KjNJi9BuJWMXr5zeq7fEBRIVizZr2XWGf96SKa+bxM+hkX8wfxD8pA20vZ9ZIHQsWIA8HvUguaYM
oxjoUQeAyYRAWJakfHLPB7eYUDBOzLe5VVUsASBcR834rVgn7+cQ1LZWUMSaXqyjeg5dWGGD7AHR
NLvh6Vs7ueotfAfKNCA59hWbPY6hzYDgXoUmYnDlNUjnwEncf4aG6IsmcErNe7c7Ut/svXzymulT
O+wO7kCQqSn28EsTokcFXdgpg0JW0nBbvOSqv8kvL8wpoltp41QwFHVaIhIhTJDz13mOAX6IddGR
Q5Cb3coa2eeRDJXJ1yee2vs+ih82qpCpYUG+9oWTXQENNxVl5HQ+eHcEgCr9J4UBud+UoE8XF5TC
tFR1vz8bD/kF5UH7stSc+b1+vEwn+DvRcTT/8VfLnbmn+MFst2uZZsmTu5tDfAvbFgg/XQGIf9X6
QLD77kyQGbiE0QVN/xka8mscGOxwLqVBf1fMg3n6j834QNTdlWW7Xmz9PsSQcPXwsbTD9JJUAD/e
wUOx9l/XYy0QmdARddrQCM24wt0Mssom95BOulLiLGZcXClyY86C1T4x2DwJaQg4IidiADjrRgEp
c3M7GFgrhM2kI6p5/P88LLSUvgjtd7P39Y5AJwXQmPXV55lSWZ9H21bBSg3ZRM8SUAiwy7gA/tTx
L6dDARf0LDadJyEDsKNcZXKYtevO4vRZYKjH+dxV+fYexL9cBjaE+nokUmDIeucEwOc/dl1fX3qM
75hw38Y2n16RLPL1hIjlw/n+xmtGVHnx4+O9mMC3bDS0IcLcIA5F/sX44YqJTAIaj3qeDGBv9Hi0
BoqGzQg+MQh3pYTlloDGARav85yIC5ZeS6mluCWdjhaFQZY+QfC1+4ymOfwHjUue6RixPLeJKBMB
wK2VQdSmPTLLR3PgOChET4r3ohCWIuOjhq8XE8U2BRi0qBsKM47NYXsl0r2IV1jiEVQW99AFL7rt
oXb82Cv5oI9EQCRHSe/kQsx1R7kbiasse8EdbBglJNGt7t4dVHQ9hSQLFY6lGa0BKk7SkWygywkN
lj/5YVe6FvIY8U80+og2TRVWS5I/i2DCnhM8Vsc7OjI0o3NywRXUMPiX6Ii2cZwyiYz8f5UBCz3c
WLKtbqikzAm2dDcrE25mfEqNCmo+IRQzYsLqP3O2Ipb4L3JITbFvUPdYLM/0hacleFYTFJgBH5us
5xEmLGn2Ms9NP9go/DlfAezadUmjEfICRCccEoh/6SKU0zXIz4rHUP1b/l8o2560m/Ew41cl3f8O
I6JUWph3PUaW/2aYUpo7V0ftXxcPk1/QEltdGK0t50JbvtlmjEt7hnMrP0+NqQAJ8NVd8m+hW1u1
6pGDIfUelp2HM/ziPfTw39FMqfjY835ABG8XkPMkKTvQEPnBV3yHiX6z0bcriI/tPGpqU4tZK021
+06WxGYCIFdhYRMqEojknWxJ8MVPx+wUAXzKmhA9PRIEq0Vso0bg7yiVn0MEJMkkUv235HFRZAs1
YnzjdnpalmeHaTRcbPQi5J2lpmn83qd8wlDi/O8pVafUdrWScVZICyyWtGqNM1vxrezOO0ewGKUR
jFJhkpol4LbZs6HZY5/Rfc+fbCy0qXHvblu+7abz+ulZQHCuhjQhPaKhUVapmk9lUhmHfYT3CVfk
YBos6+/6XMfmiKTIADOzcOtKBaYhX6yv9srDIbz/lfqWLLvzh59lHFV4QwZmXlaAr3/mDYQm1YsW
EhLWNc1hxsey/CtnULrT6yHNxUnQrNAGty3nCBsL0ESwApFDVI5gihF6aO9QUOmXJj0YP214dFPx
egNxbBXIoZnpO7f+QWMOp8TRBuzBgdCCU33yJw6r/vPm7WaWcRi4DfYvNY04GDjyIokDMgN7DeRJ
41hIUDoKeoB2DABrG5WhScKdW0SxPSGy1irW4LSdR/0iqVLNT7tCQrZ7D4yw1LuA6OOaANsm2wnl
zKIwKAhZYvz9JhmunRPC2VJfSiMwDo43ueOjnv+uvJZiE/irvqtzOVVwZ7g9kw3W34YKnC32gazQ
dRoJb21+UqzqxA/QlPmBOby26ozN9mFmk1QO+lH51sqizVfrxgKuZrfNDPpDzDbm7WYIw4qsN19l
fBd1M1p3EeEmi51IvGB+nLJ/IdhCf3mtKGmiJ1mYr8piaSZ9LF3wNu1qvp70ywB4QmvszMtzSLP7
NGfd0iewks5eT8lz7UYL1Zvz7P/M2A017HW6OJlFfkHh5TgaeS8zhTAsg54KEy17PqJs7hKMf5kc
M5b2qKrvxOfHnWawPPBSzGxB4qLN51dq9kminJLjOKVuMd/TIyXjGqS4/xi30spLKaQtoU6BMmyH
iiBojJX0oF4niKDs882roUOz+og+cb1Z/VndCuXMPzGpzakq1Pqaeb0rSEDDDR/OnAfnxTu0MIDn
38HIdmMgXIBmo5IDiaySxtZS3Y5kqX3fOY7NqFHUVKjgknXJk0VpKZATfAUcDlVQYaTa8/rLLY8m
cT+FYfVhEfstXqhwS2el+FGaNPwuY64h/NH4nJfvfGlsK76CjFJlIByxeuq539E38y3dJOJJ8qta
RaO9VkchmuQEHgct2hKU8zq00xsO+kWHTh9aywlmppzAGQgQP2mPjxTLGzlRBzp2kVn/X0Z235/C
aU47kQylnpZ4y6byuQ8snjr7kaZTGLL7uDSuxtlaxkbrMhmijhI1ybyxuWs98fPzxYDrWTr1mQNs
ui35u1UmU/t/BLfem4smir9uCx6AjThwR+vf3jMDgXVZghMUNCurAf9l/XDGCeQrEfQZNNw7RBH1
PTln01FkhEe7SRh38aDpl1ykeN3YLGyf7zCv1DT7uZvuj7XQSV4CAiUFE6A4MkYK5CppqOlevtDi
ow4hvW8s//6XWhNeYlaGiameVAl8y0urdhJkJMbNO5wtBoOKSiPYCgpPNu4lQsiqPkQzPKo06VN5
tkPbi0hWUTqQPPaE/s1rHZSiyEM9IUq0M3+HBH80qP4jncKQiaBSG9JmumsQw7khebBZkyEhJgro
2Qqh36CTCGm0Ronzc2zbFTa7uGp18741CTAlTI/MTVO5P3D7vg3UJLLMke7uWtJXn8PzH5IYtAky
31taRRiiasDvfFLc1rwvzdVpYXQ/+qU3N8hFOiHL5Ju5GiPirns7mx11nSyFWlBHiYMuXsxcd/g4
XLE4YJC1a2IxQhI9VE/inhLsET4UVE9+NaVyB1uavCjcTpi9//t9v6oJ43URnuI1z+iTvOuuXMqI
N5cbCVNSsZv0PbXXDtDMiJDiP6qrScH22KTx6XPSiBqQTLtoxFWzgrvwYqs6YLr/WlG6ev3aTT29
tUf28IYPSlELu4VptmVn62R1qTd0QA6a/V9eBKM0g4pRNMHDievX4fqruz3dZnwQzxybwYYkKcIb
kWRQ3pYJZt4NA5zaAYhUc0NyBpVM31FfIL0Vubeqbz8HywjsOaYYr7wjoSoLqvXs3hSFBgzR1PvP
E6iXN5+Voqi6bVATZdwP1WfPc8up0Y7eIF4/lvNf68RlBENtbvAx71NEVatF6GuSHfHGE3bwyNNe
bj0ma0JMb5PripI2RPcis0yNgIZaio6ZzI22hSiGIJK1lY4SstsG/HZJ3+LEhSLuyrHECqKxjHGZ
DDZRaR4lH+Xe6CpHDAXrnhY9rc+FRVUwvKHhqVOPTLfQK6wcGiIQrjqoVD32KQYEQfRc7o9GgIxy
Szsm44dRPm6JH7QI/D4P/pJ40B4l+O00gC5g2TdfQ/V4ceQs+mpxWrStOHJlEq9Wp41pRy6Utg9e
rgU8NX7rwZJP3XYhuuHO3ZDQA8K6Ua/MALRA668kay6hHc9IgFZRg2xSCiQ1YK+L5JMH3wRNRCyk
GjZE7v6IMSssh+BQbC4rKILMsZhw/EZ+f6JW6N8CRs5nv93pRgeqdCRpeizX1XL150qHSvXEw/Yw
zl6mhFKBiG0iWSuFxXAAq6Ra/1Fqq0JIUt4sT6+w1rfaTiMZsT6vVDpWho8lJAtLdmQLoJqtSbem
o7FlfAQ7CgMqnG8IQcOv68djpiZUmmFQ5T4BTxqtQ9pScF0z45Wdq0XJS5vjgBcnqsisIJ2zsYjF
v3VUdy3YYj+Ak1WqR5LDmdp9L5+WQBilh4oqb2Iyjg3AXuerBVw/lHzp5Lisqb5MrNI8nB2WVKFh
rNCTAA8XvesXUdMb2HKvaSbeqXFucxT2Za3/eagEqVRjoKM8rb0tlxe7HRg9ZGZ5thQUN8CDm0jt
fzGcwDJKGraD6DCIZfLx/GqDsx7DL61VdmmrsB9IbTMgMg24xRIeP8KKwhP1d6Are1cuMlCQGxpv
cpxYFFO8z0DFUxgJCzAiwPn4h5Ok0Ha+Zq4EUXtjXZ/L4sPvL1tBQ41zQvRNbDXGXhls/iYfoYby
Tl3NipKScDXhHTCs2lOcU10oYN05jUp2tz+mLOlXoLiKql3bEizZB2cOijdeGw2nao6b/Kba3BFW
/Ub0k6PF9BLNaZzK4aTtinmQZ9W+WPNk69fyLrMaTDipEberMgiZLXJglkJUd6K+AOIpFGmcvYtT
2OoED2KFYNcyMUhQ9cAsBzozM3qvFoGqWWNXhstw4AnV5ppZ7INdzSN2cEa7QKCmNiIc3wlJW89e
agxyM6t/myxl1iECzt2El/JLN2DoP/mKnZzRa+tBRkKHhJHG+FqQrOpMJjRuewJbXRQmu1uAas2f
1wMXwDOVm6gVgEPBeMTPofs3H7ToSpRG54h++wKibwvwuEDzjb3pcp67pv0vyEEMbxukSuhNa/Cf
TWKv3HqquiGVJd3KXIR21IFwxh+aC5Aqney/6sGXx5yZ303kJ4FEbHGVVDd1Rs1uWqQPg/6v0/RI
58bCkIBJoornjHvEbSRlPiFPmDYsoUlmgGCcq2FP0gcF4bcbONuLPW+5loYKAPL919O2GpqHKQgA
NHY9g51WatM9vV51CPKwTTaJdXO84h2p3pzpdUmgOqWpgM5AdffS/KyBZbW6646xFT/MTcgVLdXY
wReB5eIBDuKIx8/k5u5NiI6qXmzLivxGrXtKA7D8Md27uaUxagwyQQn5u2/EMtkWw+VCz73vrCLb
V7kwc1LllPF+54xXyuVcTOhX2N5T9cClNRrcW+Z37ig5JQTWCXkIevgokhF8rXnRFzOs6/fSeYXw
qur3XBJgGEvdu21lcMQWXjgn0wDWpDFIMp9q8R2vIDwIRQ15oF7zO7QOW6OeLD+APyrEScdVZlxc
ixfKpoDTu3TGnx/RgCD+9VCt3t6i6ZX2L821DPvRWo5A7NF4ZUYDs1Si0+DR2sch0/OLl5mJQV/x
sWeIn/MnNCyPCi93bGa7MTrhW+wsv0Fq0NfVq1UH/y5xTEpjM7vU/FBX8GGfHADkHh11xnpV6s//
asjRM2rLxqf+vtHPTX7cHbX/iypve3625wfDbhIO10R4BPJ/D0FT00UNPNEewWvcJENTSWoezQnu
xG6n2BbU4AwLWl19A0ku3dQcHROaLuJK/la6hHo5TKUCth6Xh5P+ugF5sxFSCxgZT4EdnIA49zDu
xurb9FoId+4OHoKksjBCGMR/qMHFCQJ0YPyYsDG5fFD3/HnCG62OkdfV4FNDNrA+H97LH+YsTB0E
chF+HVIfsTanC5phzvgZuEqS8Gox1+noIgalHd0navXFoejn/A22nP8wmWFz9B55eJZ3m0Xb/N+O
7DNeWyGLt9WKBfxFlyUPob1LmZ+3gcby13NxoNXK7MnQWpdmnBBl1Itr/FLRnbLH1IBQoTl+rw/T
I/5y3WjzloZ4Mmsi1+VTw035mHjvW4antcgLKoe/G9I4j6z941ACqoAyN2Bt8uFtblmJKIchrut2
ktrlmAcAFI+PYX+HBsrt8XruNzZbIlwZECWREDNdU66jrLsNlkU6MkY2LNa7p5qv0/nXYW38iK0u
Yw0EJrZ3eOVnQprb2sN4QD6eOL6iyOu9CAzPEsVs4Z7Hn7rSrPxt0w3toysXSv+5XC+ExL8wk2di
KmfDq59otEndeELN0Lbn1bnlJRnErOnIDo8O9axXi3w2f/UF3k2aQjqYW7gGWMfb1B3yVOUpIlyQ
+XM+5qmTaXMfLxZFc1PNsYh56fGRlBAL20re80VcSGi3t9E0VulCfDwzdFms0QLgAtNnPeu84mTA
Y93rpxvF44/+cSVNVqxM/SOHYhLzOBedcqxzRmgvnGQ5DWFXACEKSUuvKe/MU2Z3yLPmE5IxIm4k
jfPuLZbAgslWDUVyWF+PecmAj/L4M/f3iUIq7P8MnOoC4cilO3qDI6l6O1Sc0Q664Kw/qWlBCkct
t2ZOPArHuynwteGgoPIp78FtTsV9y5dB7cly8FHvRXWSRjsAlaYSN5TIMcssiVQc+PdHFFRmTpuL
bWS8Rf/mf6+QHmFwgseazJvO74ClCWpKLCBZ9izFHSGO+EOHyBYjlnA1K0YmU7eznsUxaeGJp8yu
AoNMiQoGbunxMMY4mry8B+Jf2Yvwx5hby2j/BhUpQzHOdB8hYmGjt+d5L+XRfvWdBdVEGOpxZwKo
mSId80yqZ+5sjvOTqKrBGKwpPzbYcKpSiCbkDNZSVt/+uHzNBFR0MC3g1WmM1mXeFhkSpMSBrW/X
lg9aLbIeDQOvtE9V1wSYXWL7dDKE2oKMqtz47mExvdN+FYXAO8tE4tNgayYAnvLzwnEOIP2YbpYY
+XlEvg9y+bJ6HUTZE57hqU0xdFVovtmJDh24BMH15HfN3VOZeapf9QzaWPeeWSLEqjyZGOgpE8TN
ZnC6isSIQlRZflMD+6V8Y/R6V0xZjBnKt/VeaMevezzX2O7hysMDBQ5qnVnPrdUJ5b4xUjrnNMOA
yPKlPKWKxbjqXDzwb+FnpyHsrq7HL/bbfm+U4RrYyVmGpoQUyDt1QVY4+hbxCp0w+1PukYa7Fzgf
tt3YM0ai8tKPmw8WlX6ktB3fvz4DxLkMXMj6otJWCoDVJm0BJ9hPblchAdZS7lZ4ncRBkNLX4Ku3
3bxgevOLmdntLvYG66obreUpA+SY9mJkQJkp1R7vW5BgVVreWM1g51CrWrY5jREh5ouQzKtBhM1E
7y6cMWtOXJymTTHV92MB0CsEhc38KPJUwoXIikdK1EFjeIMNE9pad3D6wBOVsweE+xQ2MzTrloHg
tISJDjduCtSHczz16TypryGcz6l9UsV8BvoE9sO9SC6q/KIsIvAq7K8qmpIk/hmJ+GZiTCw+FOEh
/m94PhSqPAE/H+ItNRRQyAS+8VHMPWH9mpoLa07/FQSscNbCteYJl3k2rl9Tt1qjfOSbCYJtJ4Gk
BisAEBH4KFuTv7QQlDKt62tUdii6onwd+ma9SX9kuEU8L8BCAzB3RTghKFguR/IaZTZhIjqItGj8
Gb0wQIB1fyHIdV5lcLdV/rwOfX+31i+hoUStn8o6BXzZmWUISvCLEuIOLssExHPgiPGFUI8XN1Q+
j8V6MlvMgCFjRgRNSjOPAUyQ8yxFdEQSPyGINz/fQLkXhgRRVTOYw3VQ1BtLRObJJiYlaP5TGvlW
RjzfoT4BBz61K3rbq07HL1TVyt6VtSBL5bnLwpZkepcD13+HPyQ2UabT+6m0VXAD7N8IHIsOA78c
IvFM0O9Y7sgzWPvZb4SCZ8qbSLr2yYgi5y4zCh3KkrlQ04qBP4Ttwcmz8RjBQU8+DP60qqeObNF+
GWCYSSrB4cP8qF40wTNdkgb6/CByfZr99d9gv2iQAkqcQohJDBOnvX8m1xczs5aC/CF1tuTgLZYe
ptP8E8rnljtPzDVHe0xS3BXEaVnUHFVPM3zOWhBVCoWvuBj5RG5FPVorP3eAydayh9cwFMIwwS9b
qBCLYw0eLY8j9lR4JYVoHNj/GOYOjmx7GFhLkCx+fsMCygXuXSz2KnMZMnrfIkGrv3B6E4/A5zFC
n3+lkvO5+sm8ewlM1aj612VK+PUJLSMn9HNAJW/5sfFjCLh5THlxeHy9wDy5dxSW7tzwk72wPdZe
MorqeV4Fll641/JiZ+/xz+W4GLEyOMaspBPffQEyr653/Rf+F0ZQGNyZ9Th38xgUWhwbtn0wUw0T
ofWPt9aDkqplmbL6cLIm4/4BEAeKcY2DVQ43Zah7qQvulXLsIkWxLeBu6lWIzTapuucuDOjHvdYj
PFTUnpj8dEPu0QsUpGGyP7oycwZ0sSjBVwN61Q3CFF03Jvf63lTLZ2lxbYbp71zf4An55aUl+3gl
V3fGHqFTNelfqXLoTfw2VuT9CAEegtaK9TSDKPwWH0HGMpr/navdupI89rTWUGpFjId2k+JCwr5C
7Hc+P+iTGET0R5ZaTrRDxFkYpfcBr3e8564ZBys6TcDw4jqpjAOGxmXG7hEmdSroJvWBMomXWl9Y
k1mWO+tcFyPHvQj8O+j9GFaOwH1ZDgG0mVDmX3tS42YKBzan5tpLnZJhVsOhMP7Mi/ewfbr+EUt3
FWez1rvyMMaBCcMU/aTSAS20DCAWJiWPftPyhUtJopQK3mWebV/h5gecDqD7XFIKhWeqHE2YRSD4
n2BpvFtfMPdGj0t7uas42rbhqvi55Gex8eQnKkGkiwasD5VFfwAu+U+SF6M535X3J43NcEm1KNrq
GrMhNh8HdmHu4LHubf3jUn0Yy93i1145t7rSPVjvdT8+wu1XFikS6aHQKenYZ+qFLYb0H4pX7zsi
2RfrPLCaMNm6pdLwVGzf2OCtyRdoZO72gcq+A9Q1KaAyUm6PY//0Tq5cx3zwKFrls+J6Z9wrU8jf
+AOKxdX3yP1EZsEayXQ5bAA2kohOIC3bm6EpPFvwPfkhYZI1Ix9lDPJZdkuKj0nGcnOT5Jb5b/Zk
KDzJJL9M59TjTPpSFQMOpE1rqAEiAmwUKow9HAnUYLQ3z9cknnLCEJehSZ6dqL7mUbk3e9tzddZP
+3OvOo8NM9YMiDOC6vMsJ5mu69GH8RY8vsttKItxWv/SDAraSmrPaBaXhjoFp7L6k8R/VHVy2JdG
Y/kry97NiGeR6xYAl8kMWn56uIzjJZeuO52PUNJ8mdTGGMO+IpEg1jxwFWG+zq/MYoLXIjNlHcC2
GIjYriHfTy0DvNN+t8Da2SAK61YvYZ7LQYe7l/PJiOY/7MFYFjd36sc7eMypmdtDVTKqnsJgqiIe
0y57J0rzfv95aVBOifN4B8koqY2YzUb1QbHED/1c5chuOPQUHk5MGxtdsQ6OpWOkZ2IZHH0ST/4i
EBH8fnI0tB0JBD9x60ocZUQ2s2GeKYmypfcBEPjsMfC+G9p2Re3eS+E1tmt79qRDHz6PJASrkwgO
EucNF7F5LzufNEnO/Of0s+4+PaNShxNPp/HONvq+lvXCM248u+BJ0kC0ogOaPODtprEv6zN+GitS
uQW+3Fwa3MdTOraNnF/3FO4n4eCkq8rZQT/Izb8M4+iDU9/GB9rWHNya+oZtWrrL9H7S7pDGFqi0
dIqu3X4t5suTqcFh894Qxc+Bvmlbec4YyykQE9jE2+J2zxIRn5xXBhwidPY5BV8W4e0W3+zizUJa
v/WQp22PZMfyAAotPAmD8AZDSPoEbV0DGtLg8QjaPIptUsU2gTodVOKjRmzcPjHZ/vxmrNYRubkM
SVEcZkh/Kq2iDuqFohgD0VIOYX6OQYfcX+k5XfhTRpL7ob831lD5cJFLeOT3OKOp/77ZOPCnniaZ
/boQMLImDz/bc9wgm7l3/P7xTPC9FLNQ9+dYi+raJzSxAAqdP5ypLeoJQ3vM1CwMELs+PtUcDeY3
LPKoogooK0LBM3auCET2yIjikXzC/dy3pWSDT63utqUXVSXo+djPm26/8XIbv04KSC1KI6qEVWR+
LuysD4kmNXpWhn/OdfmAjQRSPOFlHea+7/Fy/OJIq3w3m69dUN4dBdv/pDm8J4KtmRkSaFBg/8Dn
paIvPZGM73e2QzIkqrO60fZsYy6nyAz1IXzHNnoRDXHJ69JGWKsoC9W4ztQofifo7BJJcETkn11y
aNlA9QwwZZ0lv8sI1WU4PKrYyz9TgASszZUEVtUAiQ5iogqIt+UmIBpudLZ/q0wQZeg1KcEQvlMB
2Ln4Sb+INuduZqXah1OEJazv8jYJO2IBt84dhWJZJEaRLvl9CHv5xj2b9qzh1TdvKB0MaD+EuMDM
SQs5LVoqokAGfS1TT//pxPMc4Uh+tY36gLKUPeQcNePZr3WTIx/5B/MRdryVXgq9BRFscdY8lX8F
q5IxvoalZmh0DPDSyAYVBIkI9CMSt/B6fWvwnO2mzWrC6FENYmt0B0XTN3C1WSKCVFzvUIzEOp/U
TwuzaNcJerKtKaG9Tl3nunKiZ+HxIHz5AQiRD6LtbfKsOyk3trZzsPq+/XXBIBfSXxGJ/Lb3quJ7
vjVbos7TFb4+MEc9OPJ51gihL6X/9KrR1Lg87U6V4/XGcCidb1kAqkxp1FJT6PHbw9VHw1seyFwY
TuwGL0pxihDxBP7ewAAeefimqsFh2YSJQzksVsYFbUuARzoK5zDlqGxghDGWVVZOYsOL3+jVuHs5
iaAJc7vRu66FahdP1hDuhScH1RSZdvXD2MPkFhMXXkOquMOz6r196QiMszLj9Jdl0buPV+5WEZM5
YeT9oesqkYtrG2yWnQgyM7TFoIQlVwZuj0Od+XDUoqkIB/dq4sEoUlTg+m4Nyru2KYsEe8FAGLFb
Mzar+VRWWyogToXYP8BquH1HbeesHKlF4pOp47toKXtXau14KTunf424uf/eB4hHNPXVkx6+lCOl
lEJZtwrB1K2+gkDY1u+VCUMjjnzSBb7X3zjyO5W57SRs2eGFgL4qccaUTS3x6JagilYQfxtOETIm
N6Zp398JnVmUtvBmZnv2+6bE1ABcR7dTN4bQlhahX9UPqfGE+U/zKAuPgBtdVRhNWhDR52i5lxkI
DijM7yAknJwUs2L5PkjIQePTA86hbn8lferMQWYHVgCuJoHtTuOIArF6bog5XMRU1F8PrPoUrNoi
yVIBJTJfk9wvVT2hvUe9iEnxWBwVq6BXwWhlkGP1ifFoji/h0itGPRX/QyU6gWRV+sNctBqBVNVG
QusZGtEghQNi3hcc03WrX2rFlg0AvpdC4pNWHarzm634/MxIccrddVp3aBytUgLdnxo8/gvNIfeh
w5bciA4WeRV2xq6dG6cnTBYBpdeLOLdVzFR0zSdpGSpxQyO3ESApcSeEz8qZJNSvLXDa9tpuhWnF
DPSK8KqvthtQMqPApmz4X/ahwP+hsXo3+WVwlZ9Nyl3GvbMUl3akfWu8kw9SBCz1+KqtepWexD7r
ASi6x8SjmoszmENlFrIUpJXad3Teom8uLvGrJmfzfsFt0gvXKrbWiOqRl3P3p0IjhBdFUVMsaxlc
HOFGAFiA9YaglZ8MOP58TszIXK5jN23/R0G9ZVEB6cQBS67t007E7muwMe0560JAkhGJoXKmRZ18
L3SC7gi/K4FbagBkJul48BkNfgUr1Ga22HbsYQ3EVkKPex+JDRmUPToMXOUkdTyGH+fcxNrU2lJr
/ttgyYwERIWKVODE4R9+qxD+uzx28uk5JutBMcKiswyv/bZ7Pmycp3o5m6Lep9AEmo9pZ2DwW4vB
OO20SLxdRRyW8GrwpSxDBROSAw16XzIv01vFE69YMq5WNiEMsM51VBVVYlcu0XGHWxOIfevpQPbw
5QbJYYmicAxhcUlL3aNcYQUzEO3IcKIFxNUtLGx0Ee1JJmlgnYBJcmQWjwixLQDJRna5UyK1QQDT
ZdnuOX3R6lcrBQbtBr5fIYy1qcLjQLTvdjH53zRzKVSoKqRdFqsJp0tLcWEPIcGhQdfOI3/dOg2w
sfClvyYLSfLbG+Et0AQu9yyj4pbcuH64IHOokEqcbD4P/qEKxx/QsbwPRX0Zv8gn7IjmsZuN6Nh3
D76RkylzQRM6ymFFvesL80S91bOCRoTzHRa4X5G16h5S13YT6C6IQYG0dutkzoIbJ3G26LKrmw0C
oeGIbc3tM9AeCAkrC2PrhBVhaF7DAlEuUTzak5l2geK3L0beLGL1YJqV6944d8FpaMkuX0J5dYKa
84OB2X49/owimYsfjR3UtXxkwPLt3CJKQjzeNGYPCUUraUY2FAxoqBv1iAjM+LPPXxFw2gio7PjB
19hu7YSEzrrXJaC/WhTkL094kzZRSpBmLSXY34f+C9tiNgXC3lv/gy5e71m5BnWWaKJLHtJ/aY/K
Q2hznFjLs9ei8Vkv41dSMRgNl+O7R0+MCkuNU6+OWx+7vaYZ5kZcyaR4NGvN8b325wKj25Ej7BKu
mLIpL9JFpAhN8KZ2APg23aKcosKK3ughNBGdTu9vCaT7ALJO2Vm+o80kLl92dGC5SbBzjjQ5k+yM
6GwuNskI3rzRpo0kZL7zY+AZqXlbWKJG64c7fQMirfv+sUniM+JOfLmJiKmT0u/4lmXdVnN3LFQ6
PHj1Ua86rHjHMDsHtfyQERN4XcqvCZVKOgATt4CwKeQkZOXbJcakJ4zylLvOzECs46OMI2gpTlIk
gS66a6o47qBThNFCozSdm/QRiMo/vGOfdN7R5yvcOm/auyQQBm7wbUM/hFTr4vokg92LfEApG5w3
HQe3FpVHlrFsMTwqBybtCioTxXG86ihKNRGvYulQ0aU5pYheisdAWzVG0K9isdj131AaDQOl0rmP
2NCMiZx8mliciyNza+GYhryJIXR/5DimckKOYVFGmUgV/Lf0SziPl+zYfJR+E36HfKDw8HnkofLI
++js9bKp3Zp0F32sO8MQHYKqoPEjxhHI11vp+fUD9ZVZ6c8DiIKgueoRUQTL42HHtVyULS/dT7rP
MfFuiqKM78Swm+rNCykKQG7nDoT0PRNIQ8Cs7gi+sf1dsfaahuyh5y5Rm80pui90N9pDlvp+Ykno
oaagAs4IX0J8TEQXziMdLTBT9JokC3D6/RBPP/ud7E8or+NBAesvkwJVtgc2G6Wc6/DCYBrY0o8h
rFsz1b0SFkVLq9BC2m44+Cj4hEAG7w/eN5D4cS6Vnha+fzcrjun+1U0O2bH0tVUpqhjCL2xiI16s
f/6Lw3qTN9N9tctLYe6zwSxP43BwElayxSneqT3pIoAweINjmU7JAgg2/8YYjdUBouRhSxTl5Qgw
NaSuI7m+TKOy7UFBXazL6lhneOqkFv8brhU5gTdfrivrhQEAjA9dtnEeKVWxq3J+X/g0HvSDL3fF
cirfjH2q4rteNgITMhwCJyGGG31PWSq2xAwOR9q+Y90AIAR/b7j4fIDWnWy3Pq97pd5dgDqQtazM
5H5K87t43AcnPzRgshu5DCdhKtZMxBqNnJ29kYNFIm9rxuZD5FDrHqmsbiP9wz2LPaRwlbxqfEV6
DA5J+99YvRZfuYeCxkoQVZa6trukj+5AcHjB5v2nHIhg61pWudBNEU/meFmvrl2HgcbPkjLmaRlA
JeJSVRl93Xv7u32bGcl4CPj1qss3RmMIaL2gmiBk0u/1I1aWIqSzFOmXaSMqeoFknr5//g9U1Wd7
UGt7PIERzvsgBLDZyNtKZVuoR7MEN+uuno/HgmY48D8kOQ+ue863hHzLElyqncCH4TTxsobop8sw
BhTR8UYSsQcmIa48sLRsTpVT2eFOmNgjYAsFcPqZuduHXJ0T0Co+7y7gbCBvoVhUDZhXNr8BzEeX
kH4vIEhtI0iQ8uWvinXEKt9Y1s//AXJ2t/t1WT0ah46URYXdUCTVUJZ/TO8tgoBHhtU3lUe6uzsl
irmw+coIxDgcfCo5yUN3/AOtlToBB7Xu4SSO36viBABzuMOcBK2Xg8bhH9+VK0b+IIXiZR8pKnvV
bEsfT2cdfETC486DIvLJzbKGV8VmdQuwIDYG5xcZ+6HjJp+sPPp3LcjGgSLVEsYo1wy4MMRMqtO3
rqmQzAqFD3qYcQkOnxfpz1yng7Ok1dGY8k+5jkKAEIvsuGKHqISccDFbai7TgxVBKnu5seGtqidv
WKHl5RXa5AKOzvL+BR8sYxGwSFiFz3+wt1ulbNlfHoOT1aLCZVR+SZtfsThfIDxRGCYyXBmcsOxO
CETpNh03XOccgjJ20kwg1XJ7F7G2UyeKGBwDkmEF/a4i5wF2gGjI22guLhzRqcU9XRRMX4VQnnq/
G8eYuMpjfn/K3UjXBiL/goW1maZHXRhL6DtiSxOoxogdauy6Qt6QP1qq2fqMTwDFcVro80P7aYYB
k2xkS65x/mTVpZrIMzqrAf5JAsl68dd7i8i1ykfdaeYbvSWBs6zmhuCifVn/X0X/2h9vrCrQ2QVv
Wtsdsv86QvWGagwfV6eSd3MOnFUt0k1VAt3v+tegVHc5eifWU1zFzS6wpCA4pNdvl7rzknG3xJ+w
JtBJIoP010RUV/LMgVcnZrSYb5+Lbkh9wty+SZLu3AUrDHPB61o/zIbQQnmMH5eeKMPQpFikseQC
bYEU/NnuENxIlqG5AzULOlFye4B+XOe4UMYwJt8/F55kRi/Plyd91zKrFtQ2gNJFtmI2pdSUrXSy
ad2oZFZTxYwedC5HUsXsHzkrZN/93bdsvp/o3q+tW8ttKt36aC8uu4PJDMxLV28JN4txjH8Uzu4o
Myq4RU1vJI1nWD0dHyxADoz6ZoqSQs379JpMPvHHS323q/fGCWSFxVLF1wZyMK5prFRL4VuQygjU
MdMxB+jImTt+vOlJJFSblolR/tbkvf3UtE0uN+4NHykg2dySgUqFjGiSTT6sNlHxRaAiAsFTgl3T
GpbCNM8PSGxPe81QRPl/OPBXRHY44CvXzC+DyuySzN+YOcu/F9v3aAaeHx5PIJv8OvUmuCY56Kst
PMa3t0M2fs52tq90eb4Cqcx0S4DwhiD+EcPH3eaKOQpgl03sVWFbZQqJtx/Kokb5Nap2xxjzwa0h
rRKneCLRBArMuPSddXCH1d7Z0y6ubhuylbKhvS+WTxgPoo1zFESyy2EgP1zp0miXbiXD+rG0G5np
pfublfLldTG6z0zYWbPAdnpRSYVm2HKtgzUFFWwarz4ZdeTkw7yKQp/jJLO4uWgzGJB5TpRW+BF4
eKEVvDejuyKOTX6cu5i4jjtJTK9cueAIKKvL+8ZpDTRG/zDkED9x3+LG7+MZo35ungEIKyfNQ+zu
TjJvWK1mSrQHLrBTCMzyWVFP39wNgg0T7zjbxNaj/ejQvy0/JnMNx4oRLtSEsGQR0qim4KAVUgUF
i05rES5D0ZW9o2uKxULg+imZsIgUdADntLNzLYUsdb1Y0dhqxHesI1D7n8rvmpzzTLod4hGJYZ7+
Q0ceByC5R5cPVDQ7oEG6nCsETo4xEYqwIChKAT/zUKOlbB8Y5+oQw/I867fDB32QuEK53sitCLju
avrd0gvD8NP7sxMvu8m3WD2hrV8bYoKPWZetqrI1CU8U+599FUSoXB+FPlCzHCkhbSJ9L1x3VCMD
Qw+immKCXK2iN32tNp715u7cibL68hELObr64YlZWuOF73EuUZqBA/IUt93Yi0bWJVOHB14MYQBk
e3G+6UhECqzP/O2BHNQj8iJeEF0FdPuKk/h9rOn7BzvbUcmZv2yvA11JOSCStky0Lbxv6Z9nIyUQ
nC7dHXD8wjHwJPZziMHt6IMcx2u2uwSVbNoAGNmZNm6EyrxiTFdIdWPC7+AbT9r85QiW1Q65vdR6
/H9aY+uVSX0BgqOQYjfQtRfKj1gbkcExVeAutGh9SWtxdTwnkL0W74vpEn1HTHfrVy7x1Bf/3Eb0
TJPFbPCurcqSDWDnMGlevtyuxLreI/9fznqS3BJJ4OhCjjuFg8m4OGRh/AlX/ZvGeINQX8unu5Oi
n/Ul6ZTyJa4UFGE9NuqQe+wBPg/PhY+/xsGk9x4FAC4A67z7ZLennA+U5GWqfkG8jFcAK2ysawxi
/Fp5gQVLNbDXUr/pm1K7MrI3qEhsuceTlSB+2vlVGqvh2z442H/f1TR9HQaiKfkJQ6JDOHh/lQOx
B+vqmY9XkjdB6+tukU4bOmlHDI5M2CMZ1/WKX59c7t5O5tORy7qbJ4cSDxJVntX2BluTDL+LVUUw
7jwEYATSKwguCYSpliERCz9bBqYYK9nL9ibczS6tn3yZk9B0LGMpvfontlyH8jq1k3IcMyh6LE19
9/Sg/j+Sg3shlCKYGwObQMYwEcqKKSqjUHrAlfgpUNZDZuCnKEiSMcdgFdL3krYdlNofjc7qze41
G6oEP+xBqi4DeOgc73aFpRlC+FrEeY+rlJiHU2V72h4eY2VdueLN97JM30F7zdNWJDHsLpcDPCg0
v4CnGM6P3qiJjRgfguNG3+jdL4d8pO4D2Cqkzo5hMeYXBCEKFucN33wQjnZl7tskvpfLRX+Lrqp+
OwjsJYk9Dr6v9L0EmUvnAJlSSRcHV/rY9r3779q/QCQ7R/JmOJnRbMtVo2BoycVUFbkGL5wKMChN
n+f779GGl8T74OEg2DqPYGN5dT4jzSJHRxsVsStP1RWuBgBrX1oQhMteb7U7Mv4eVFQXAf8aT+Xw
n7Axx5HuCaZqwcSBJlJIEpzNB64Ai+WA77wPleJUVg65UC0iWVai2dCQM1AABuYJ0BjOxPxcyTxJ
V+QlcbYwnXZ73lyP45Fn/PBt/F4sK6Iwu82N+zpFshp2y92k4wo45tWMdU1NHW/rdpoI5ZPOBjKs
a+B1ZYh9KjsTxLVq0cA6Dz+u0WWssTCVoSJmHg15j1MlBVWHgI0agRK7+M0m4Wtgdm+lhgr9dlEy
sk7TCK+G2qDHwNxW9hwSfqnHbjj4gCKrRRhsTdAfCwaXsIBPv3tXMbwr822lKS56O8x5sX/qZWnw
MWPOy/CQcUas2YphpMz10LUcLMt45IjWyx/EQIWhIL7XjELTgtqdr2zE4fstwBWVv+329Uxf/TIy
/zqbYWZThzRZHN0a9LcZgVGcmskkBHrfOmT1FipL28USCKeS/XwXg2dsdpMK7rKt77BTfZUuawl4
MpqzEaHE46uyGMbmby+uEpXr7/f0uMOZL2mIgj79XDUYNCCwwjIXPZjKTSP56TbZmZFaUIvPBa/b
og+P5sfSzxsxbH7wACeMTk/IEHFGdRN3oveHbDvmreb3siKZLB14kHXZxjPxnnwowP0eSJr36+zT
84XVwTv/j0qJhsbxST2ZmYRiJ6fQUw7Ec5hp9Jvi3syB2u7rquelp7MXzRZthAa+95iofgqeuJ03
+BTiF+c7gQ5TE779YgnfxFHMChkVrgANUv0eUfwLveaUq0SDR1Ixffhc4JM1BamMteF2o+LuYIia
YFqBvi66gDikFjxWVGvs7iws/sgAt9XMxXGdcUScn1xvA2jpWsJroPhsSn/EOH1NHZzrsd6T3a4K
z0R0jyYzGjDypLDyFiSF6s+05d9aNq8iXznOXJ5shVDpA18/EbAVJWwb9H2QCKBQWQQS6aAV4vUL
UP1nuKjfLJrECfqcTS8kyEUyS+Ta/0I9hR7A/0Hl9eXuLxiKvbvQormh4OXRNrFwoo/cxMD4lp2v
cxfoAG9bzS51tyDaS7OHdIdEyBSW7fTpeKJfqXc9HP3qTD0y6d+V7KCspVFPO1QyoNC+5w+zbrKo
DfiziJzbbSQ2ZPhfgTS3Yjunf0jQMFi27jh/f/YVZO+D6UFzWklz1OrAU2WFY0ydgVRb4GF/rAln
HMAc96JbBmpYbAn3cetxzhODoLEUIEa4vlCeQzLV/lhQGGjYufFnqoJLsA1XtA1Mo0te283neRNd
gejn8p3fY4m4gEE51Artp8Zlw/72KZGOLtSHoykLjLMCbH4b46T61AVKaawi54o+Vhjv1ujCmdBu
4RJbq9UpoF3xWONUQ2bxbWl4S/K+Ii8LgmIOPj+1I8cq6sKggrRKPzLyZ9cCpv395eK+B+1/1tIh
+YZh7j07W6pQ6BgYoRo20zYt02F0g9A7rlWygRHos2BEQl9h4Wu4pU1355cAh3YvKjlQb+2POCsD
VxTjEfnYUlShsWgVXUFQ5bt5VzVAvIrtTGm/3Oyn95jR7ytIjfTztsOkRUG7xIla7OlBSEvPjULo
v/TrQdCTgyKmG/XGWeJvyrLxg8coHtIe9x7K3clHMzRpwCueGpg0VjSrmO72CbEvpm7Yh/zMM4lm
+/cAgrNIEOgMDbFyW81jz+oD0J/5rkOTdib/qhzN9vmQo30kfeHigUf38RRQU+akMIy06Hqp/THF
Wmk5PF/EgECzYWGYpvkwkYKL06IlmHkCThVxpm38qJIbcybSfjHLQRmR/4BEbySzWxgVTy3vBxD9
e547/E9iSZoJSEOh90lt0jtBa2nsne7ff8xnqr0qTWMMwZjdUrI855slU63Kl1aSvmsADtJPPnjX
CE8tBKwOe5j1gvfdO4uX66gBMydAo3mUzMiP5/9Unm6wE5U/5k2X14YIiKsEM0Qky04LveSs9YAJ
KVxeVSR5KzNg4/jAwoJ+1+HyqqTvZEjHFm976BHdPDdcziBRW9sVkuHl7EDSOugMMdCfPL6GiMf6
n05Huc06EdxOuoG7b/t6fS5X1qogE5ncy/6t32ei2kwofVmEysgQQ6GyyKRM0sjWch3JA+0pTLks
Wkabe+FHWcZMFCoGKLWPGO8H0DQFFiptVfVoMIpby4+UcTANuwkGqyXr9PBA3s2mFMa1pAcejyg7
jRQGFui1YFjHpgmzh+qrAoucpK66NOb/5d35bpYdmPYPz0cuWbcBJ53fxMRGcvGzkH4FOLTceI2l
vGZzoJ3mzYxywkrFS+vb8Pz4cqFNVhmR+STyW4ttokLV4xfgFZ9VbWUimLP6uh8752sNYfpch+Zn
+96GlzPr2gWlipE7fCS03oV3YL/RxNi/fJk4tYhfmWAeOSk9ItOYbdeg8WoiO/dKzMxwmJiy7Ree
7tXijmj3UOpFFkeqfqlU+qikIw9L2CPAmHxj6AkviN5otZbVlXRSc0zj8Juzbhh4InzzaHXJ431z
VAZDvExDQ4IdCugMEaY+RY7Ri5UZTbdKtYPxUZgkOBitd6HwpNGnpxx2y6eHUmis2V+oqBhpShxw
PHmoiEKo1nnepsh1g76v8cJp/558JlbGFJxPERbDXiGo5OJPi+UIW9fcqfAw+l7o33BonlCvG36+
uRcejRDTQJwLqk2yO/SicV8W1DBXg4LMnPdp36CD5BAQDpFPh9CUixrp+DD25pH6bHkocvOMfSPA
DmtwVoJlg9RJwgbihjpZXEg8evQAgFDw325uk4M7WYPijWy6NkntKnnJsIn3mkWQoRGlBwmNDbfy
DBHnBziOQQJnthJQxCrtDZdHG0tNLTDFoXwX6CRvG2PtCDTeHkPNWUaKJnPWbsYd7WTPumnpeCzr
gRR1OmFP1vBwm5Ccq2zf7H/z5Bzrdd3+xY4sWtblcK0gMlzaYqiTZfTIq8h2nwf0EgyTLy0lzLgF
dgDNwi/3hBo1JkQnKYg77ll+H4MlcWU4a84PIBDxOUr/BCud+d0HOq8VZECeAo82bVqXtTb0nqm+
HWzvvK5nrN6jpmA05Yi25FSb8KUTJHbVXtYvIeP1GEa+FGCi6We/Dk72w46x4gtAxWLPqjY3h0ku
hV43YPeB3qVRdpnzDNs1CqUe6765/k/8ZtDEcWhf5oMakmWKxQn/XrmFwYN3cOfPQ6RGGx5abctS
+X8WwMYJDUcPUYzSnBQKC7kdVN4tOJMB9wyjmYsfzpYDq4h928NZhEYIvLDGiQHQ/+QPofqR+oEp
RslpZHlCnymbCR9LJJYYQh8kko3n1RXbd4rjICapDFjgpal5zoqcw3cbvCH7fRcMwEWviZz9tEXf
I3zBKE0GnxGpwH/S/5gJgLtIIO8xhH7PQTFQkEXRMMZXxiQ/K1F9NtvKFH/P4YdiIgBC8g1oZBcU
gf1qmMNAMepw5LkGDYdsccKKwT7MRfdNiWzlDUiV1VrkSYUCTRNG/WtEkqJBgrSjvTmq58LY3e91
wR5rvPT4ldy5QK+NtZm6Vy6+lE2sCfkEpzPO9eZOm7SK5gxgdEriygHyM7hdqvtrJ1hv/ZHW/+FO
QiC8ksHwfjqKB/0LyUQcxN2f8wkHvNj4jsEFosS/0cOTYy8SvHRbdmeT14kKhbjj0zdeAuxbV7fa
cZM4UKW7ayPrhZAw2kreIosoe+B838qaXnAxcIEHhuWnpz4VkQDWoKEmNoGa7UaEwh07GB4EijNx
Pt8Buh+179F1VgI+yNO2kpWGsd/TwpgWdI+6bMBmhZd3IF1b5d7Bp4hKG/kD8i2d15rMwHd2wr06
vi4ynKjeMwx4298tCrLEFpjeWOfmyilXcqR0+/HU+0dxhb7iOMvh3kKCA42CsYKECa2HaXOJYCLP
jRpjbCcjmZZDz/jcrKp0/vooKmMYyOfwjiy8xi4vh7o2SiutbPSmfyC00koWebAD+ECxILpKGWUS
OsabEIUqYPgS6UvCSO6uP3dzprUBSlh5uBgVQvzXCckvN1IGI4EeNQnBltW/wpaWP/mMfaght5EC
WqjborGpNl5uOmfdqsMrzW3z/0rOl1FSbv6KAWUNVlKraY7zCEFy9KEnHxfxgbfi092IHUSETIcC
p1NHEWpP52mdP7Wffba7OoJb9czEVqUnRU2foT0ulgzPSrp7eWRZv8P0YvXSDn7elLIo2qXVpzQ7
uJtplHVj49ZTBLE3Oh3a+vPnrI6WZFsWjVLccYC8yaCe30wsZPrr/C/Q8MH28uHoJotWSoRmfwrY
cwRMgpVIhDBe7hqNl6KSbUH9peNx4YnXJHhgWLdWqRl5HqKZUqimB+O5m78UMbVWiEsOAwdGly3b
AFQweb250dGDn9k4LOsjtfAc70rQhF59zSTOXYSCutJL0wAGLJJGhGvafBfPF2R2vWyB/lJ2Q2Hu
U3w3Wvt2Ff+dCLTU8dvsbZdZnqsRwKeLmMjCfLvZXGn0lIyx45bgYdTET+n0s1PlEYyCgQDEBpET
pFGNIYGxjlj19YLqd2Gm2S2/XoJOPedpXdxM3Ll12sGSpylOh8Zzx1ZnmeuYEx34G5nsur8mp3hW
SavJNwZImmmBU005V7cCzVYgmclkVe5BONRecVZQxy6RI6iFynYMt2F8ofCLPPZRvqK4x/CtLe8S
8o0MH35OMnuNKm6zAXAwDq+Earo2LtquFFm50WIBncxGmDNnTddIuwTBlnUeEm8PWgL7pY+zUrSG
qOpT06DDhqQsD/0G5ZEaP0mYLKubbB98xoU7W+9wbaKpDLNT6RG0PpGQVMmQemr1xjPxKthx6Wzc
EEdBswVHULMALXkFudtb7qfnhFB2E7ZvVud+ISwQ9oXktxo4lHdr7OhE13so1ALJ2ufxShImaXh9
dsF8uVOOu9lNEmqyYCctsAj5zx2fHkoSmckHGSNoO6peJY95zU61JogDPXckg2T7nIQMFxvjcF3c
EPN7HcUuegAqFN0uq9Th0dG8GZ5xh6PAKeCbgLjIhVF846tbmt8/AEMWNI2xLrq3beicJq5a3beE
u8HmlIq65WLjJt9D0HoDpHBvZB37hrV2L9g68IU02tDLkoe9GG3gAoPO+hMXjL5N2LFiwCf3cYxY
BVkGqtuslZZpux2SDr3vTht1TnEGcaFAluJ2bNXEO+2JkrlEUF80ouimP2ALwqjHY/nCQ849NCAJ
NbbJzJrDgGlbd4wIuqxjRbhUz5etKXYkWKfWT2DPe2Fs/EFR8oJ92DAQ1nqLjKBKbxiImb/aAmYC
f9JvpRuxomimmarmt9A73B9jFAc2dowe+DRqvIKmycsTT+2hdxW9VPtV4sJiBIWwuxw9rFNByuDx
OCltmoUUDlwJ2PazXsyrVAvMObX5dQN7maXE/vgkzLuZpBxvBPaCZ+BDcG9+OhjeybhEAyq9oOPD
NaG0u8By3vedVGxXa9YXSN9tR0u6dwWStYpMKqpcDqP6PX7HNI3Hz62Oc2ELXMmx8Bo+Mk4gY7BU
nk3g8bmwV/h9BOpd10CjSpH+9ewqCTSc0Yode++EljBooevxzaxcJv9pXJch7cx7bCE3/day2yES
PaSpLb1IXARgace7hJajV85uJAWbKWkCWQVDj9O7q0GdwVc6on0DHq4pyDv3pUYN5MwwBdOleaZI
e0Hd/55SdMBzdtd6aEoRd69Q8eu2jdFxNTGbiFewltcxM1s4Y9rGoHfUq3zIaK2p6L0y1adckttr
7TFqQJRxPT5163QdQvl3NDxMuNR4vblR8FBejleW7uZ7kcWUvrKuKqE6ssFUvN1slb3xS1FFLom9
cME4mfP3dTh0BKO9RB1c2woyNnCqp5XXQjNZK0n1tI7I+bMHnHTvEGtH7Tw666OOi0FdN59pw+Ii
HnwMZtyPedJwWK/9+/pAZ/B/jpDwMw55FGvEY5AcB1SrRIdu9jZmByubug8v4BqElvkEq4nLFgCp
s6cHx735exb0gky8QWYPn7rg/PQFRbmZG8DLzrxWx9aIdfxnIJVx4Q4k5XDBWc/B9NNjCIh//AqX
6ZS1z23s78O3WjMJmTgwFWOL3RwX+kh/PQdI4zX/z57/61yh2rQFKRP/eLOWkwEJWJVwxhWGviKX
1kbEPkqq4hWsnIAFWpOs2Zr9TCKJd6S/rU+b0j/7sb4a99+Yxf/X21CX3wOOlzdGBGeBDjLhu/0x
h63+vGNamkgwORfrxI2QEpDt8ZlKKMA1OJPJV+HcQQhu7lXRdQkMPr1hHwW8eN6RSGlVbYvxAcje
pM/0b27bwaYbXbHubHv8VzgMyqeqwDU4F2IHOFtKt4elRF59c5/6yXEaBuQlW3HXFlazoOAzxhpt
Tj11WhjjJta06ZOsIgK0EAr6JytLf9pJ6c7RdhPRPqhVnIH5MYJAr77NinDY7OqncGklMYq7lXGX
9736cFGVqfXGm+EFM20L93KWnkQBa/fnm4cOa41MXzIziu+ByIcdBiKZ70iG4a8nNwaqQrruaFN3
DZaZeQ67AeM7dN7ALvjOJRFTFHB9w7/sbbqCLDpGT11IMwg6dqOaM3bHWT/okI/Si6trQt51MTHq
d70k62T0CzeAJOOIQ5qf/INzlFrzTeK5EBcnr3SOv9aF2tqrpj8r7daxoFpSkyp7SMvbWjyQRi2N
WCV5Aw9wfysPLFH3LWkzVG4EFRasF923jQF1T3bWK48mgLsbhV0U73mI4+Wlc8fyBczL+OlgSP4A
KjWbHtTlyIwD9HaqihazFtjGFqxNGDA6H7amlVDGq9AZrUDN8NUv/FHagW7mApCP9Ttu5VdmW8+4
1NANDyEkmFBFmVY0yf3qSiBgh4SvwrrOK0BZpdgRbk6cUeRxjzUzNnA/hrdqb6OK8zWYRUMUCFR9
bhQpJ2Wg0hMP2TFAeBUM0tp8cL7CER1Ffudwsc93zSsPq7rR1rgnGa7R7ekyjYc1360njXU2rTzz
RLY+JFB7Kz+Q6V/KIXa/MfHZp4X6bj2wczX7F9EujAVFMZCRuZf1uzGJMcRTFSvW+/5nuVGntYL5
nynwh/Pba2KgnjqQ31K16jr0eeLAPthGLqtPaeEC/BAdk0KDlVFmy+Ftpr+f/OZcCAmrlhtWNDdM
OhFOqGd6LKF1sRhRsg9Ntw2V+hUa7aaBPwKkqJF1bZRuTDN4DsFNE5kPHguj7UXWzbzYcOXmgoIF
qOAvs61fppbNueUvxX81EDWFTd4xiq1jAkW1G3s2T7UyE5irILoJleC1ZPGJ8dpK+yIAXkoiNd/0
ZoDLYJP3i403Q0VsOx2cP3MDxHNV+wVQGitC58KNzYATQsuq10l9WUaayUrbclVeNj0BCDU5sJs0
qtN9BjJBnE/w8cZWAiT5nHgEPvsfSz8dore8QGTu75keRdAM2EJfByas/3Xi2nMbRTObed0tMU+C
2zkxqBe74qW9abIknHalAsea+pvcVsiYxI607AN8AlgW/awE1mbqtDxwhWyFzGMqY5DANs/6dMnD
z00/7XPjBQAHtqiZBExYmfHWzVw1KGgNEcXhUmzGQximgOzMQKrtjc2RP3S40VvUb9uTtfs2fnfy
MecNaB3JMZ0kYUI9vCLf8ebcosC0kmz2JTbA3bFF2Ywh4Oxze0aM+ZlmBAdNxYI12bb8yyvG+OXb
EEPzVMcvM+Rc/SUMBkyJi4oM3Z3h5k5IqjSGGJ0m/MvtbCRBji16riH1O2H2tdtbRueh+kg9fOzr
YB85k84CVmNFWj1oEXA050SHrUiprZaw3epGwScwA06oEtPCXA3uItjLz2LaUXLlygdrx7qskqq4
oZPINA53qqJ95ej+00IrK5bwZlEV4WCBbCkDKnrwm9bqy0CI8QDGGRGtpJCdJZjhNBN6Lv7lYsay
RkzQXSrvYjBcObi6+JY4ezcF2bynJED+rf68SMIUH64WTERmmMSC/bjiOqxh561eBhRbj3SKDjz7
a0vicWxmtL1oiwRh4LTWse57kJc2joVWYbTPLFn/7KjlJ1JmuKDLDCFsaW9x7MagppXCFfP0MmyU
a+dsH6xRQEVVWYoJ/U4rhYrziP4f0DmfogyV0gTD88AJxW+NdQHiqByi5kf1H0Xc1tV3b+8qxuoG
urr6u3APv9MuJ+Eq2SnntxGbNjgks5X4zMKN+rPCbIiJ0WQ3tNFcdBlk2kooJy4UFEbhuEGoHZRs
nXqRiCqQsyiTqrP7wUREuGau0nMaAeMHVOG8lvM9qD7GR0ktTFXJEKjwvrazAFFh7A/X+2aE1t6I
j1fJrOdOj4ofdxBx35sfv1sAzC2kS61QclBuHtBNZTCtz3rQ3mLQWrCniKJrSJsHvKHoSXYYeSJt
Gwba0+eOcHyvdrFSmtdtoLKwjs8XJUlfWx0yZ6pRqLk8gr2uf8uN2RGfk0RlcrqZAxNYYSEy+tUp
cG6t+dGmK+ZUMgWB7j3cvc5WOMzUKLofHn/7rhKXRjZ0fQbWgsbeWtLdsrsqL0pcCt+OiW+XnS55
Z+GtvMgLWVz6jG2DTJZ6T1sfG9+RI2xaZbO88Rd8Ry2FtN4r8kInL2FRsKD6MKcZ6VUwrVJqYaaN
mb9UIhtDRo4qPC2uts5XzMG6l87sRwRIWEfQ2s5uvva9w0b7jA/KSCClZ/r2q6pNbcNt6Rm40QEs
KI5z1pP7UFYt5ndoml+EeXw2MrIBVK1dpOL6D4lTCStkn4IMbTwL39vnbIQ3uRQScnrhygKLTqiV
8lU7S250bbY7jalFp3dsQdueLrUBhf/Fe4E/3llSM3r38bC+YM1Syh53zB5tPWd4ZsgwJI2I2lgX
T/bOr6payEYYZhGVut7aAVE6wkF68aWrtUWOr7FMfEcITW0Qkx0N+jD/C54OyDXuWzCsKDbjvf3N
sMt4w5bQIZYU0mfa7DYc9krt1Fapwd6H9aj3xgHN+MBPaDxXFjzaYKS3twXbhCsju/NPmJxsukIi
4+iVXiXDxYDcdwUaxpwLrmwOqcwG6sxnewKYKbiWZdyAZsPF7YU+LGNmGz8jf7/6+GgnejiBUXJc
wO9bU85iwL+goIVW9Ju4inTXpqd+KxoFxar43Nop0XUhhUUWLT/ryZLMOsrSzj/5cScKT9DwobFI
5/zWPsnti60/bAofveAwVeo9+3pV5l3alV0Vxn8s+qi2Wmuh1gWd+oZRHxc5/W5sxUdydL6F+erF
RNKbVqUzy1+Jd+ES97PO0uZ7CoWlW6DDVnknQm8UjeV4bBq2HuGg4sshpXELYE5XgSRMrJ9qmiSB
Ym8i1jqAwRN77LD3pdtewjjgDkGf9hPtIm7AUhj5UnWWPtHYX5ownesUgqVkndgAW+Dy67A4KjNc
Rq3ltmFtLMW8WUahH24nWBcMYLPPimLmeIFza937Jbq6QVnvazSYrNHt729lgp8SeaDkT/TEtLqI
MMmmwegyNM4xhWaQpOv360VFP2JQNspgLz85CWJSE0gNZCscdZvonQI9x35eJwDK2pJsPiVFFjLD
WtFy1JCi6qwhIA4QOh9p8vHLIFIm4t9/YY9/00RGLZ83A9y/D6xLUrtr5BIQ9A0oWJcbQ81sX1xB
nYHEjz9q5cWW+lonm4ueucEt/7891mKgApoycSmR5FdCrwNnM0PP3473FeeyCCbfz5uhiAAPYNYD
+KyfrHtVvLJiqwXYEGSoI/XLVOwll+O71xQnJYpUz7XuPw9fd3j7y1O+gQRkmPnU3KD1WD0DlcEf
tRbcvJM+180gUQSh/TLLgMViVJJEsICczhS+HgNcZsU8mQMq5r1tZs7WV2LzfrLIPqdIgYhQBABo
BGduTxACJU6UhGaxbfZJvuDGOfnrVXJrqpG2FWpmkXivuU2XzUTng8nxCNHuAIPxcQyxMgEEZBZh
EnXg0OY4FWV44PL+JxasPvTp86vshOaJFY7kLRYYaQLhhKVHQf8hJzGRGqn1N5csxZ73319L8NNo
b2Pib6f6ljNbsUFIZn2OzSaJkPF+CRoej9kaIZ9m8JmZsDPCvWlvd1iXuz8B4dbtnw0dERuGTkJ5
SBnHHGH7DNsE3UuAfEdF8TURryoCG2JjptKwig2mdI07OGfXKW8hMAtVskwRzW/4WlCMM1aSg3Pq
ubYQ8iw0m5sE4iFQnlqDW+XI3xy9AmSyGSJ8c1ImYUZAPcUGTEshHTYhEs7X2VHZhtySATAPUiPM
bME3zz7H8qYdxy59F3AqRpI66FIuNTpTFsdB33WJsNBFDyGmrQpE0Bdaq1heCszObsSe+v3XzM4+
rIOyMQRu4JUV+NCQGcCCXBE05CrbzEgP/akB/4O7oc2/33zmCsHU7/trQng/OIr13QzxYFWeHyRU
6dPLen5KNOTod67A+yzZa11BvRxbny9iYgY2cuvDb6U5Z6Ka4N1xFLZ3L+Lqkjpz4L4V1QYWJtYt
jPRI88gL5dEe8kbEVC20dKsX6k0g5XVsgd3b8/5MHgF1JLdtNvs9lHnG7R1fwPizWUS27GQcbVqx
egm8xK/+C59dyScMZcoWBvu7yxQz1xZ511BqDq46kJgWqzxwY+Io6tzqKZwLWKnQfScYYNXUXtko
S4fHJhVoIN1+s+xO3ZEI7HESD9AOTOuf9PWItQvliCwQZ2Y6RFHeHIdbAKgBGJcVJ3wxYXyUMh3j
rJLMXg3KZ7+LbxPb35C3hUaRNnmu3EE0n5FQW7KUhbpvtZgXZTwg1Dk4e3cwu/LAXrcX5WIIklOu
gZKIVGx1obTbo3gkkKLYjMP3OJIAUkolYzgtXm6asAoQ9UJq/rAiHyrThL9zIt4vsygX3s25IJlR
ZHE+ECpYNhYrIa6YDaZtJhTBka7A2ZVvYmIP+6wMkrkMykpdnLpU7fJJ4J3mA8agPPgpUZYz9QLy
4uPSQvwyuMz9GgT47emtA1po6yWlpZUbk4sOS78/lWDBc/YrOzVYdyEEqOmS/u84bb2amvvZKd2g
jgy8kaAvUcU/zdOVx0rmInDmmdBOjciXsxbYw4eONZRqMEjvfLFPTof4MA/2WJl7KX0MhVwJ8sZc
6E111shahMZkKbl3pELtEAJP4SPrXlY9o0N09Ltj5Px1jDEn2QR3D0MxgvpLuiSw2AjHJn0zJUod
MjKjcsHIJ7Fk9bQZKHkmBbS/wkx7oQQZQg/1LuT7qO9uma7wA/pCriWGir97hrxoOwWgtr6WBopB
JNPPENHejpHwDP1Gn6ZkxxvvgYHG3LHZKIbGXmnvmAvIz6yqTIHA71Fy8cDHBsaMDtPA6pKkIKEn
hr5vps6quO4/PBMXwGaBcYsX06oLCGk3I9/YbFZVvNSYA2mzWfJmgyHQZEsvSDZrwGy8nPt70rRb
03Sxo4y0ynm32AB0Hq+jB0vfmxP2Gmdr+vCb37FjijddcMmQMnJ1bIedwobcQWGu3Dsvrnvz9ZhQ
+lsH93JSu6JwSt1XfzTGqd0uLDtkPEv6bxPkBnWWWJHZ388pCaqixQXjX0hWgvbMz8dKt2Yyqnge
O7pRLBbaHAB39QxdqTpq2ay4zkILTyuPI6pcKFKSdR5BiY5mNTDJFL5DXFte4+uFruw9VZVEIONS
z2ghnxnfXsFP3Jvtc6zXpDyTMkohAOwpPx17y1wUvmNYf7uZOgJELnMGi6i7ZJTXCD+0yIczkJfR
SpOUwt960IKAKUezF1cWQc3WcW8AkjbyuZayvTGiW2QSD9PcC8ZTHt51REa9dAI99SuL02D+Y7J/
zdHSXCKPmiTqTPA6E+4Ym+yJs7dtaYENm9YLB1KwMt/8fn3tpCJuRfG5GgFRQYwt5aBtehlebNY6
EbsUSonaTVoXngFNMH3NLdv3dhZHTnqWql+Ysb3GrzdxK+i3b06BohCEWXmBSmNnFhXSrSQhPsGR
TwI5VbbyhLLz+mw2h6A0H/ymA4uS976NEdUrukv8g/c54EWUzmoaSIujUonHXuDtiTmzpueQFDce
+bND8diMqJoNSJqXKAmC/ccj2tuKpQF3IETAwn78t7fLvtCI+zIjjmWXpvrHyxKOVyQsS9Hp/8gd
VTAN8m2jA6GeWi+oTEiYNITEIQEDp2pUPWVXsd+EnulqE+y4+q0AAYX6ojRTzgZAm/fDNT+IYGhW
/mqjF8W3i9FBcGkKs0O8080m9R+zuDofJOqbG79HigVnNygXVhNW7ujTZlTrTG3RLMXe0PDUvVxG
F47Iquowv3f6640R0Ej5+SOK5lDbVMBMKr60mc56DnCD4bR2iOGEC2CCNISV+rrCj7q8gLBdXrb3
MBE0e88jIYbWVRU3DNMQfEj+iU1Y5LTDVUBBzIfu+6QB0JquCOPlgdIcMEE0i1/cp470SC+4HCRo
IVAQSMAN3ucF3aDj8N4k2rg6rFdDOtUlV680SFhWve39w35dUSDROxXsRQLKb+Lt8CKafJAW/E9l
q09NqnW0TLG+n1Z5O9mfvghpk/FXJVfgxEhtBT2hXyTAGuECsna2FljWtl/CeInxWWnxE8QRRLvQ
QqfcK0j/JHHDeBQ5VaSImS45YEuyOVFcY/WvOhARVxAH11CPXObbkxtTL9znXucjyd6e6/1ijN9h
N9DlVIcxRrBG8KjzfPk8gC57NBofM6ePl1szPe1cFrVjcLSeecs4RyGul3xwGUgLSsbxXuP9baah
qfoBrk18yA8X+YGS32rODsOqmTKo62nCJbjfK5t22hzNsc/M9OonWMxFcmXZ45XbbRsQfEr41zRe
VbW5JmW7+KRHpuKlFfRhBIczGMqpJ8Qrd/yCy08FuOWtxUxuBjAMQ+Aj/DV780Vm15OvifufcOQy
gn1lRYmYxbNR9KW0mdSTdZmhT5RHd1mpx6PogLfHumuPliDncsEC/GBxeM9AASa0GhRT7+kxlV3B
SHUSLAQ26Nxt/zKxBPOPlnfvAIehd4D3TC298Zkjav0Uf9tNdXhUWPwcXI5oQzJmGs7fJ70vYbBf
iEyGwmBxYSTT6bWUg90Cw8lvMh54LHq11wUTu+eyoMrMD7/EczxiHgNzSphcjoH7RBOiVsNxKQBa
BXiF975ny5jgLDCGPWveUQ44I9s4eRdDAt1fBWc1PKDA0eeEc8gfxjqgD8nq42WNTZwQ+thD95Ha
N3PjPNyUZSDHWmRNeV6glKt22qFJedp2sv1P0FTBj/m1MThtsH3Ym/NEOwwPj0r2i4WGshGiJbRr
PeukFnAVdppN/4YwVcDakjkAUoyI3bZVv9zIq0m7GKg7eIymzfgojbnWBJx5u0pNRc9+5hWMOYU2
KT6Cpq2eLb8PR3q3dFLNuUMlf+KpfTXPHqB0Rq+uB65uqboN5UBZ/Zy4DL0uYY2p+ZO6BqUYj/Oj
56KRq2XS6YlYXrhq7MgAUJkeX2GLOwVDHl6RkKnMiC87e26BAdvMUgwUJe+OJPfuNqCfTR5noV/T
z8L7i+5VeUnhuFv9gRIZeyQcoeyTJoibRrAwWdImZjlHRzaRjn5kbZ0LaqH+9m1SxfOTthbRPxbA
HQb0gADwySTgqni17+SAtybULzshU1+ZDClxRkpSh8neo1kNRUwQcyUN/5yKKCymvLnytL8ShNPW
iQka2kGUpP8wgMQNlTYh5XYnTlooH2VkFXW5bQxRfDJUJI6OY2+J5VW0c979GWQXXmLyya+pmvU6
55r/J8/TcHLaO+3OactfA2GX+RZK+j6/NkKEjYcgpeLNbET0YvROZB1cJDOfMOJBkIdhxr7HfyYi
yWjrvphfWJvfPq6QlVIAAq+CU3x5x04XlfGDeU44NVDf9+YRZZn44M9ajIuVwQlD1x4TzH1t7Wl2
ymYDze36tcp6Ne7HigEVaPnXD+K70mutVfb9kH1T2ZychVwF6wk0hFaGNrcnb9AxnwJbfjQQcodf
rv2J46JTnJpuqMvyvYiyU7xIMoVoAG2ky/N0GPowneo9pSQQ9uzhne20FxqSjH9MEkOmhc09Ats0
J/hyyHpEIGDKrcMsxSQfv8G/5IIXDcBpf3eXXl2qawjOUeBStX1biGJ5KbfX7jMwdy2ba2j8VTz9
YDRkIZDa4DHoySVdJ8hq7FT9A9TNa9s+B/0a2Db85Y3UpdrLybjZp32tRPwCKIsUSFQVLaSEzc42
s2NmDNscri8b06J4d9cdZtZ3nmUG+DwIdlrrJxYzi1YdG8dawOnEgl8J5iHBDAZqisnu984zDLx2
9Iw2hUj+8RZkR7vt9llxTD56CYSKs1+HagwnvztVk11wSAG8eKkyaj6vX/1QMGlw9q0tNbiqVrLM
voFJw6d8FzXPJJtCmBe77sxNw2ZI8Fyz6TE5Xi3m1ghIbBRMNZZ5IeOgLbxKFVf+x+fdi3lorkZy
VAaq9QU4oxY+hzQhtAvRKo9oDVRIwGvudT58iJfYUxue5aaUIH+3ZsZJHx2MFwZ8U0y+tdXnPcDy
Q26zMmfQhtVBusbHMnmaCONoMm5Nb0tbo/aYv610Vi6kFqS61cQ/eoNZ2uuQi21rLDTUqwMstu0h
NGEcoLqbC+OrJgiDgd8q5rfFDy+55goJ13wiz5ytTq6/VCYlWj6f96PPuizUZu4GuzwozxVaeLhQ
5KDw79kxnOCfSWGHWkVOvkBHkrPzrOqRhHmUimjIQ+A+0gSMyJwt6s6Q0gQObG2SaOPsGqBz20Xy
YLGHIKPsEykWSfZXovzEL20X0fPmR/MBEMDseH71Gk4YzUfgc1WsXcZTe9saipfHgoDNZ0PsM9Fh
TcANb4HHiH4MEGDCYwbmikzxDbcsAmhsy43w6dGh79v3E02+KCf2ZpjNGBx8ta0dBTx0x3VtORCD
H9FRGDtf6+ZeNL3S7ICWLa43PwYvwA9Cp3vmxzROL5Fo8xgx+0ehGkCqJL/LPPPcuoheWcmYQgXm
wUKhyh7J3IpgdqpDTKRlyJPw5eGfRS/oapNNKvhLBZChaGOV+LyweApL1hOAwX3/zPqe/73QKVL2
syocEyDN7ll4TEzkjbuX2PVmPJ3ASVjV4yulCyujYP5oZm1Yjf8/Bdb7+7r1qqah3Ml1elIrqpjj
VfO/mjbhW9J3/nK/X0X3xnvIqLccKY30MrPXm4PPL4RW+eXJlBT4UQgCNyEpfCh7MoZtxguVNqd+
0WAg3sqTl5xs0IQURHCIw9aRsJbD2/Ym3bmNRfN/0+myEeZkVgQRn+6JG8cRAMuE4xvHV25W9g41
1ZhCkE2A6VyxzvrTzXvmZ28Iph42T3Q4rF7qlEX1ifQMOZ6b96J+PydXJ2OGpgzYOke4yV9B6WeH
/qRcwvUe7Rcfw9f7HsJGQMHF5dxDCt4FxPGHrh+b4Az31UBpRLSHRUqr2A2fOSgQdBV3bKphX5/A
rDyZZNm+Q+xcpwne1knhebTJztjSqH1vrX2nXWlNH1bGP/IN27TVnQovcpQRACnMltCEvOmopk7j
akVZoDXoEp8cCB1kx6jP+vqrcKg9MxL6FPpEGtFno2+E8YACOtorHZb26xnufme22QmcxK4squCv
x2pPzXdidOMU8I6Zi/n+g8jDCxAY+H+U6SvWDSx2IgVOJDW7v/vvtweHXiNtla2qVdpRpqcSUMTP
LU9RKhkPxoHiyrhhEBIb4ZZRK/WPgm2wZWw0+ceI2+w9unVT3FQecaRcvrA3GN8G6oYQBC/bApsm
50STfVh63XEAqWEQx38uMmAXEoaNnJgDfgpETKOHf5+ecVRczO6FSMO+4WMh49A9XimFak5QHv31
iiSYpq4wuthC1P4jHPjMvfjSaWtEUU6UW2AzW3bhGJsBGTNW43aC+rGMuGELNSTNryhNyI2/Z66v
OhSCKCUyciHEWvxuNU2aSvfv3gnhz4ueXz3fz20k5IvSelTI4JL1x0MXCkEcKeiRBz4i9FOyOwpy
RHSUaFTULuPgrSCEAOVXsZiwLf7I3CUw96LBPCtInFCeve+XDa/E3kMQXLuIH6010hTs4Ub5VJF+
zP1Te5YwSW5mEvhBm9nf8W5kFrANADhpKJx18jVQIOeHdLvjYB6hllMAstpbkhT8FiZ6WIaRiack
pt6K/bDfU8cq5xgpE6y3PrEjJzGjdGJzDPrKFgcQCfwVVh00pr5PwzfCD1/UaRPVE25riJBPvP9k
HJW0CaaxBfj/dHwDsgG+UH/yvm4qLuAv/OrVuEmcullHTHuFr0vXDax/0AYpU7/STmRUUckuCWVt
USp+X5w5NjjJ8opxW8JtlZuuwmyRdMLlAgQoTBErRCEsVLzSssgAVolejTNYmvxv/bYIEde6QZlY
B059oi4kRYFmnzX/mWqs9tyxUbffLUpJ8jSZyVnnpm//ah+rTh5pTluurhSrEiroEchofJw+cCkz
eqxHPJ3s6zRrM9My51ncjtCpijVmfV9kJ4Tn148oeax8MsXkQXGWAQ60BlLrVuuJxjUA2W2//zaC
LuSY2Zal4ctdPVNWO/cZXL3Gkv7YL7DOZny1gpBUNvuVYnXHX6BNYil43QhNl0dFoLrvMrh8M6Wt
wLp/53KMeSELSa+jD+20vZm5+0SCnaJ2F0TrDTPXEr116nwxKHesuUyCsbIcfCV6AJSgjX7q/bcv
HiI1zzMwGL9M4i6GiNCToBV8rg+gHjOGLVpcW+R7yf94NGg6jnWi4JOiw3+Dec+EM22KuAdFI0zB
d3E752iQq4nh7AnYY7gsrZBl82xUtQ+DNkHRflEyoh7atYIjKJZy5qUnNfeDNo6vnynTwZFLWasK
10d5e919bk/db9Ul1ifmmSLSTUUtZKWUiwuLmELZxrOapGEecHAlQ6X0sd7MsBSNbyHuRT1CA7DD
2KOG/m5cpj8Bi0T48Z3xaoN3b4grQscbfJCV4gk0FaLNBwohjXtPvXeSLQRT6ToTy3+L11dgVLbG
w+m6a5B7Vht9iPepr6D7za4lkLPWiZ2A4yf1ovZKKklOuR5ovXF/TV2uLc7c7x6eNxHKx/wnNzZ8
d0vITNKykt9tzsa1PjumCBgtw79ie50D2syalCl9fUA1d8wFafQsAent8bba/28Q5Dpg/B/AsqEv
tiKTq9oH4wYn6i64bBXPz0ucA7kkcm69VrVU6XNoW7N05ZkR7Z2fVL+7jrGvGomX3VRI9OQcrWv2
X/0KbjgvdFfsIE0fQ+nC+Q7BqU26LqZ/xYUyjMR0nhYuYPFglBa4jHjV0Y/EUoXykF3lyinGROQQ
HzZ0l3A/V1ZtP4JnPR66lNnhjr/CWRcrN0ShNiB5VUql/IZy6PyfJOYa/NRFph02g057oaWNRNp7
C8rRM8QhPKadYGTnhSf2sQl/Y7XAwu6ByivHjSv0seyr2FzpOGckiCWHvh4omqo5qw/Ilz2V/tvR
3QNigm6B6QKoN/aHu/qKquxqtGAixa5AzUOUtGs7lJdqsGhQyUZOc+VkmMrs8u20CEOnmZAznM5s
xUT+CsLpx2jbfM3/UzMGWL+08YgUWwD0OuPEP/eofZfcIc11/KliwOBetn/w6BsKTMkgF/pfARZg
TXWKiJKvGFz1e5WbLsv4TRUnY0JM7kecQLG/rozAMplcjADZAayZ0OIZxFjAxGUPtwxZaWwh68B+
kne5pS8eTklKi2jWbOGKl4riNGRiXo3sxl5WwSB3SiJVArVxPJ5MVKaDnNanm0KjdKjBbmEtf29P
gcrJxLU7IDCK/jIY2l5jaLfQOtcsyv8SSND8t7F/V2Aq8nLBrDCyY2X509e3zCtGS+hmxTB5UzTI
Rg7xf+DExu6xbV3U566cXV4oOr8wezcKRZjR2f0GbK5m5ys0Xc990qxjpeS357kmQbrCC+q9JTPm
1lFh6qlUEsJlAisLXv7ZamLm1SUfWHBr+6o9iIrNq3N0bnAksElAiJ6pT0spg35QNEw6XmDO/94N
VjOwtSxRPsFyFEC4IuuMGyvNdK6WnfyBD2WqTpTH0SH5gGM/kfd+GbXn9Mu9r/Kt82U+XKFxS2DC
VwmquqIolvsa9ufx3V8F2qic05i9uV8tuIpxt6sxZ94HRwE9RanOFBeAc4l23mKK2716rgLH0aDv
R9RZaIJFJwAFky4a00Q3gHR1nSGmZWbLGl56K2D7Aukc9/mTQzbTw8dYYz7S+Bxm1BXXAM538iHq
0T7K6jyw3RcxNhj/Vuiq78yzsKk+CSxxjLF6j8haROtC2XHIpZpXpt0XYBNHdTPcQocqXQmUDNeq
KSi6eRR9aBj6YDbHKQXtNygxAlmW3VyhKUTd/gj2yo7xPvU9wyxM70uRd0nRID5EiXJRk51XC1gL
6UTIHNUNFZ/nswm2+pFaVgbBV/mpZw/x3hVx9pqnE+TkoTMU7TbAHttWcAZEolbvAchOswormE8G
JqGT4jG28UxS4ONH+6gphpbFC+BRvePErLFR/rFv5yWPBQrDluHRPoqS7rPFVwkrrneht6dwHoXK
HCCkN8RD7FTgYr1voHtCCyjfMrLjlomczeSQ9ty0CVZmSMsZZ3q2Hsag8BX6q57BT8/TZJhIbyuN
92SxPvEK6Uzul6usuAScNgmiA0YAjKB858OprsQ7fUk+Z9NFck21P3wB3vjZf0Zw00gGZMK/NFHL
4Vk1uuZ9sJD1D/sMzqV7a85ti1FqF6FoLp9BQnL82FzspNRE6lZmBf03dEw4mopJfSW7FGzbqew9
6G/u7WMjiptocsZUBJbLxTy1eXdcy83jtzHNQaAZiTthg6ImnZb9WitAnCV8CBY/fLQIVRcABsIl
A0Yoznatw4oEHC01Rg6xANRJPR+Tty28QDnIqr0ic0qPV5MHXfzO3NtUfIYhpgra4AJvD+lH6GnT
1mkyAqkoTj+pjGif48ZmGSELnGXeKznVL0R0Sh2WLc7X8adOTQgprB2pZluqTxYsAD6h+9J/UgZV
3HFqYWZCXVLNc+v4rPD/UsJR+JPLrUzNo65wYQPoJE7eEb+OIGSE4BPrGQDlhhmka3BCzLxgNCam
Vqr3yy/G+u2F1gmlVe2/RfVN5L5pJQ3UcxjHW7J+sXT1oLcpyWT5MXgbs7u8sDmCd2frDuZ5u8K9
G9uefkpMxaIpHrRj/yIfDB4VEQtwkgUEXmLqgA0iXRu8OhZqu5EaPBfvClfoZ38NNj0UPXqYeaZv
0xr8cwdd9ff9JjzW38Qpo28kB1Z+S9q5Yf7ZGU1A0nXD/YvpkReB/NMDelLY2lWH+fr0N9huwM0C
xNvG9lIQg450iHumYDhZzFJXsZAONXdNbbFJYWsC2iktJ22yThp2vC0fDY6mE+wVxTN+gLZMPNA4
QZO0hSAYNtfX05wwOV5bWij0bayjLv2ntCVM26dnFHZ22nyphmTzmMdadzqb4sGiY4ZjtX+v/z8D
qiOSujz/7T1l68rnsG4GjOCcKRSHONflbMgVMNW8IvfDg0ldIvXetYRois7mN+4pekXeIXF0gbAM
EuCquyvRcuGn01yBVhfLQfRwKRzZxvCFYupEpAbsLEU/XwPHFeY443EBBWJ68FQWoM7jun60lcSj
DWEyaeB5omuUhAkLVJ7FOQdmt413G0EhZsuP8dNTyDd6J7vGdMU0keE+eZ2Vbiry4YsUnz5RC3CC
c3KrQGfUIk3dSUfFqHGnMsD6kLS22WH0brdOjra1/MXEQafclvI1WZ2W0G7fHSetBBkaZL1IzPmw
FTw5AkzDHP2WIOWnI/8mDIQR7UDD8DHNDgA4UHllTOR+SxxiUR99wV8peZXz9mnZKIt7zT8oj2HI
MN3Vh1RYpLUXJnAHsVL6zL4pn+utR+mxc3jbIsHF/kpkBUT9HCLZfleyOutdbEBVrnCrI/wiBTQU
nT85r8ahKWuz1S0KTYgxHkVDh/0f1KnKCEbQ0LnoPFb0GVkN7fCJpFP5pqAura3rus1eczNNUwNF
No0iUMn3rkNixQhBVpE12ozx21zB1TuPWElKJTuqrnO1brMQsT6FVIOiSZ/cIcdgO5kTYTb1gL/P
RmQS6oFA86RlA72IcYB6sHkrlO/HG91F+med4JGzk5/Z1fwRsKHAAZiwB85OBtSX7mDorVmqwwqy
cPz4zD7LAxqHxmhw4D7jJT9yn8wvZp1tFP16Sl5QErzmBcq5XMZBsUY4yDwxAx0mLs65H54I5mRg
Y3Y7N9ZMGW/uuJ/ZGOwijHGKknfykxJCuFGwUdVcCBpr6PV6JZDCmysIdzPfDKv90d+Q2GJ2imFX
R8MEk63uDUyQd85kWuPkmeO5hpwmu6YevLyOUTjvfd5tXgCR+Xi9JZR2xtbRNNy5XY1pc0C09EiZ
yPdgV9gLmWKDC2D7cH+lBtM+n27M+gUoYtbg6Ey8GNHnhvtJx077Md2dDxHxXEBJt0dEzM3gyGgQ
y0EMHCneDpNVwk2bZ5U5YjmdIhE0RDY84eW0ZS/jrotcARkJxDOti76ix9RrTTFKt24YxVvchcRw
uoqdtCsb2TU5nBpsFwCmVnbULm8y0VwARnI37VIx04mQi+vDFpjl6Vwl6VHtBGnTWzYs0ejmuAac
1495bU4c5i2fcJlrnZfHraIvfgh84jKQQw9pmVNqzklcoDgvd7IFre9rMONYqxxrlR5/moQgWPe7
BpdLiZDDU3RQt/exLTbC5BdcngIg4hKXEXc6FsMjuGdzVEArAAx4UBnmiaoY3hjFi1lKYFITIpmY
PLUPjEm1TvE+utzHfq1XWxlZiw1vC7O7t5XJQ0CjcsS0hkZwZ5j20zBdArjtoA+biBoLwIldTiWN
EJ4cIG3DMX8rki1WMENSKrSlkBxUuXXh9xFbnq7azUzSlYSNGQ1qO2mqtDLiVFBjOPeVGDVGkwub
hU7qBwfthmZ1TcJNB0wlpBaIi+UndoXCYmbm4NCDMDzsGeLw+vYrlx4zR652xKo10NGV6Nm87ASw
FvgfZNVqHKp0OOo/wBS/QnVm1YaPQNgkgTwCVtLvZEVuT8dcVnkq9bTU5QZawr32tBCdG9HVsr26
EkuW9YnSxU1flBqLR7jSQQLj32/o6sCY8yotGI47r7hAvfTkWduYHHyTYjQg5RalcbikgISegN/I
DFGASVkxqeCOe48euv3DXvrciY+KKFbRGxcD6vWeu9EvPE8QICFhyP6c3cYuKYmjmnxXGMFvBkwU
BcrxisduleWkll6C6OexfqYMEBZ032DXskDvtwKIlddnbOq30CTzK8vzIVOEriIqazC6kToUfFXj
Zhw4de+rR3GutsGtfZAZFCv6LMIrHOnJleW7FNDLaW4cgH5TTTxxXlibBoo6U4UgTYU+rUEhDriI
64zfE6cs4dklKf3z5YL0BMvLu3oLs3fLszziLAjSbleD3flRvK0oXNdjjzbUGWy+bW8y2Y0ridrf
6xvEGvZxaOmngJI4mpKg0qIXPPGLBwlqIIEQ0KgwJO7um9GC0FFeXDu9zUhSKtbFdQ+Zl7kNXAv5
VkdvA1YiVcexSwnTQ/0HvN5dvVP3YjU2tsuteinIfV4Xsl5jwoqrqWGRoebP55OzJ5096V0b8Ehd
XkUmLkSS0kAuUkxa9uIW9tmZwvIMRCLZUw9B/QSSJhsipNf+mZJhtxx1d/aH9sHD3oTILj5psjrB
Ft2WZVS8Veo8JFuccXq43O4e69FCOwiFK0PFeqqlKG3SyfIsF8CHmlq7m0KC4fU7WKNkcH0xjBXn
I5CG7VRZdQPIiBnRdMD74PDbLUmaq60VLGrbUKIJupJ0Jt9a5fgzF9VCnGnWRSfttL4M8hGTf+D9
uhmXcXMxjEwB9AI+vQrGKNJ33D6DZBI5Jp7J8FAWPEKrn//aCw1laL1IAtpMg/eMoEaGt/0QB6NL
1wbUyr+6vtB7UA7YW9VrOQXTdt9cLwb7Qcof5rDO9EOpY5DYacoOU7GpQEOMbxOmvMHZlJF8oxKX
NDwJLNhS1//jAt7KSx9ImyJaTtIxKiqRa/e7qHbONNomYNTG0qDunEXekZ8vpdW/3slrLt8wImdB
/y92d1JI5x6emnoifSRUmIIxliqmqpiuo3ObSuScJt98RedPRYPiFOm2Q657tyqzZP0TZ2cIIT2E
6xX94zJ3wy84GHWqqkVyhAlWRjw/A911eu3+cEjQBqkTpe5q9M2W5Uqd/RrmFmIADH/zfuQo4MR6
2sJPE1dDpP1sFY3JGqyc8CkxQOUYto/2BBRCAGv7MPR6Udfn23obZ3T/2hY+C95dW3r09bSmIrqQ
+KjDb4UHzEjJZvjNYee+qLqY7zzP7YsOm2z1trR1LqP5UJ4kWue7g/4rC30aDTdVZb7n1XD+ySmw
qp+rsI/gRLm24XgiUhImzy7hwO5LNtkA5naijNRGU1sAQpDuUDe9o1Iy0UAzOXFcN07sgjoDXN5A
4g/fXAn1nxHqSXIsx2su0LAb1amk/LZiW2vhlhD3XACZtRI27jybmjZnP5/DKAdgbgeKTCPPUBtg
35MHfnB+RyMI2v6b3lWwYDvwdvGDjxvqJcDCyemAN0KjNURHYeX17wYFk20g2kTajFOMncZ04WOJ
69gH0KEVBUnRuiGaxfhHZab7KqOn7t7Bg9pfbybTocj8PLZORk9yiit1iypQ7Q9SL1/lmcoNmsbK
RhXikgfgh5LpNdLzYfzye4y+oB10iiI/Yt0VZ8PG48vPVnbu4PotGKZ2wDeoW9+cPgH8r92apkki
ZUG9F2rKb1KC+Ci0nsZ76LsMlZutCz+/Ahdie4HAmtoEYFdUDgzORdWbArQkX+I7/+idZm9poRBw
6ahKw31UuAw3pAtXt5zY8+EHlR7a4lmD5v9WV0DeXdgiNFw3P0k46CbbuZXWsGEz1U/U+NZRJ/fw
OuFBuoeXhXt2PsZ9F0o4iDa8Rq6rkyxqCAVDqLzps2Y8fPgxF9uGUp8WXpYgnWyG4SghJIc6NzZh
VBbFgXGHqM4zS08zMoHEB85MRJJr5nsaynu25BAvVjNzuMzQOgMNNmyKYfCNnZo4DvYp8gBja+cs
Llh1uHNU/XbZ89UGj2n6+P2DTS65+0Ht6sjjHHcBlEjA+o3Vw3I/Nzq+HFMi+iq8Bv36+H2pWGTM
tgHE0WrYDbi0ON6fBvXIwFzJOhFHvwu7gF+QTwHXWXfaooAr0C5JE1F8AFNi2OZswQtbG3E7ZgxZ
jsN/FiSlhLwLrjCNdP2I0Z5qlQqhmwzvuG8dbIVfnrZrNIYWDfNnwe0CKmEb2ycD5eh7pLz8W8g5
pC+J5RJZMZl9ULPkYxY67vls2YkkyVjuSjJQmytAVsNXbcWjDnCMobrKhZqdSO7LgXbYPoCFVRku
avs5tD8Act+39p84nt62LAzqmUL4RqxW+dgwV1h0jHn3SZweCy1QBV9O5H38nX4Z6Dxmv9hA07vN
2GxgDZRSQ76R57qrocA3GmcZVfZvKy2U8fvWvmJvtlmM5Fpa69J8/i6LSwUp2obKOO5NZf/23UMA
MjLMnWdnQoCo6CngO5bcOU0nXU++cZuU2HVu9WKlHEC0BigRu/BCyUJR0mmezVrM6+gZnFVFVtX7
7D0+7ErfwcnF28QPiKtS6FHKOjq1evlMQZGZ7W+j/EAW6SyTQKxM4z/XH2rgLMqjPr6FECrHSdd6
LQLu2SthNdtRho6uB9rK5e+U3eKdH2UwaMRyvX0FvkSuBTLNXTdnBBkUHivgY4SsRvgEpqhzPgJt
RX4pHCTQMPyXMl7Y/ynxWBgFMFQsSJPvX6O3J72zHRYwWPlHywJzQrXcZiCmKQihl29Hd6J/YTmE
IE+OtJWpFjprkNguWRN51SgcfZ1zBsHQpy9AyxsrhzxHN3mKxvKwFzPDpN3V8AhEPCssDho1otYx
rGciSBzLzpEd9qi32Scet3uGN3ECYz+aU+eJtivAd1UbzQ+8WOBfkkmRupCtP3jJURmYxZWZpBD+
RlPJ0fD3JhhMzm7GHNDS8BWSW8r8mGqonsSwDBNNwGSRDsb7kC1O9a+B7k8JhbCcuue3ZixGW60U
fgBfK7UTrv2D9dngVYWr9a7OmKRH3kgP9lon8v5uwJNgIo//RinLqAxcxsOykmwKFlg9h7O12rbg
fhC/xsee4s8UP+Bgkj5jnvfe7t9D5tEwz84Iql52PRHPnjY9cvRpYihoSiUsMqdbCdFAs/cpiMl2
x+7GrWZbbCUIomS85ZHmoOt8A5FMKPDDUPLi/5jDhdNy9G2CgSKqyx6xU3riqBtB4sfrDudk4wsq
nPpgc3yV+wsoetuwmhbxwCsVM48j+YynO1ZuiLG86HJVYC6sfr0YxPMJs2h6a0rzKj0Teum93NeJ
16C6qOT9qR/A+inNjcfWGKWIuDwEok6mwUR3f+AVxkvnLrcaXqSCLlyBsZo5QK98vMhTaauDFtJL
ZZzAcJvrojnptTDzGoc2tSVngHX9xX9s3gzmXNaqxqf1SOsBwvnlh3vxmY3n1Tg8M8s5hbNOOAd0
Co+vQQdv8pSErHK7h6Trt/GBp5XrRSXy4nWDFFJmhM+4IeA+SEYc2hm1g1D0IpyUvm0EMtsJNsdY
GmqM0XTTDbysmU33rcI4JYKe8CjgwXJVpnuyGSf1/I60Sw+fGZB9Ic8qNPvjLljcsgczAwiDHJxd
W2BF16rYzbpvt3+8mpM+hOX0YL1uUNtrAis1pTuJyfzZ4NnX6A7uo3suPRJ5MWcjzQPOedT1we5p
QGGmAdLQr5gEK12sD3J4ObQn/PVDeRGknf+aIx0fsslc11CITV0UljfLb1WGmgBCXf4fTXKRyNc7
72vFHIvLqwe5fYyBN3/OxrwnG5T+kXIAcgIQ/YLLV2tTP34R72BmlbaTKyZObeNrtgtCj0sN56aa
n4Hwa3IGnRWSv0E+T38tPvuvgEOrMTtkU2ns9jfdzWWat9/IfGWYbRwWKla/gnnegKQYlDLAwl5M
yPzSnAOSlKWloG3ktcwxaBfwZApiRVYiTTfeo7JzWEKf91HFqRR6FUqV1WowIoPszF0pzglp+bzq
tSMNYWRMdhYl1n9rmsZchjgHr4YPHqYaBqY3vpJj14cehWSVfGW8fH4ODaKzOzd5d+sI+YApV095
Q93sv5PTBeBTsHbGqzWP9zCBvwVGVnscFBPLcIZEmGEVPWEfidnSxg0EJ1DDtSPxbGT3MIqEZpt0
WzOS4jOMPywr3mkGD3VCf7oIoB+ucEzqJMtydySemkmCZRRW++5nNqgjcQcZ85+qRrPkj46q9Qtw
LDAPnXP17ckWQTovg8Ud5lT3qlKHNFm3OUgFwynZj0jEMcrXhBLvEwdUu97feymSC+uDhXwNJSRF
SR72e5qmaSLZj4ENGTsDcVesccxb6aGBe4FJ1kzomVYBrjaeUwVzFoY56Ayi3J8MJuXpQmt6ystE
PovSyF45tApOyu4465a7bZbPQkG1Bs4eDcNIjzZkUVpCbWUxmch/7VrY65VB0m0fiVzaM0m4TIn6
rd0e/0MUH9c81AKe+AdfhOZrsIAdF5Jmod2fOvlUnHQSP1rP1OtGikr0eDXaGYYvaYetUqoRY8ts
K0NtyqdS+zSlTwU9Ik9h2jGSpS6XLhBffMdgoPGoW/wdgDBdpBk3FfJIALhqLK+qmiXQECPHStcG
Q3R4UNlnZdcqowv1esX/hWEwTzKCHCr8LBUlXRgnMbB6AL00OB/Y1ESr/TAZ1M/ZEXdbZ+R0tSOi
EErdAEy0dhZ5ZXClFHkKNYMgQDWMF6Kk3ZPjdI2FKMWdMZ0VPT1q9ukv1mdOeFFbQ02N8MUd7m9D
q59YApE6FtDPWf6ODCLfpi2PjAG4rDoV12GhfRnCUYE2sKf/3UQW3OqTcMYYaeIwHqw6Bi5BVBVA
xq5romrBa9yjYv9X93oz2Z4CY9p5J/BcRGp6KFsJBkbt75b8KQvfuFG40bPNHe8IFO3iSpRRFxeb
VVgLj3ee0r0Dxgyb2OkfSMM1W9fmU2FPpDa/RZ6RicP6+1ySATJ/HmFk7CfKCokZxKqTx4pNXAJN
v9J/+dTTxkqWkyvB+8uGgC+JaoL5X41FNZfDXYn/nr1pvkxIHFJuRX673EwgCmY9tDBi7t2kIQ7u
bC0VF9buFyIpCC9Ukq6wI1TQ1yxzg2xL9DBkXDhPXUk/jX2nrpzQOo35vRJ+WyqBH4fhHZw8fkmC
SDm/GXyxqZJH6Uv9alQk2n/lmCinGNKrYUMjcf96MGVqqqZIOqREdGXyVrognjVaYqkGBpVINbWR
j0YRcQi2/jXTwrLW2oERCylG6pJji8pgt1iFleSXN47GM6N3c5OUBG3GdoFYwGLrziM0cLwwE+yk
C+GCqTbYD1g+prZMzWQYaYddLQnkuk8/cNKql9NS+eES8z7PhGjA2xUHbd7JXqj1e26lik25Vb4j
DRniYYQ3FBThTuW5J1W4nJVqeDox7ZIGE5kRG7oYGROkX3eCvdZ0Qj9WQHSTk1244lzQYkMKc1PB
T54viw/5tSp80+A0njP0J9wl08102mk+sVmAMaKinFxtVn5nhjNsPAk6OPnPhOClJq0cAZi/GO2n
/rIgJxgRZgB6npFMh+MKfbu03IV3YUURTDvrep08kUdMxNEuBlgnKYfyEYxPHpcqLsFCZd75m27Q
oVronguO2P1Ld444Nq8ZSzodUp2rnBXJ/9fU8RzvL7y89XenJXL/Mn0T7Vl5xZ+qwQzhOjRjbV0V
voYiOywjqy5rkYnkZAzTUL0Yv+sB1+tSsouW93Wb/bn1dauqbZZ6IJwl6BxXMOZJPkN9iy61HSrr
EX3ba0uOKJwx54nwji6FcCj0zgbi3JaT/wraQnSjABZj0aQPTK/SCpzwu+2AW0aHQTTWEP8eEFk7
KSLR3XSKW/hykMNKQy7/Q5GzlzZ19Vr2KnJCU7FK9K+mjxTpJK7duZbxfyU4k5XRAvLSzxm2WOwu
eXEvYmWKLUy4O+a0PG3ZxUvpmSXIJWcVtkMjCzgRk1Ctxw2F9twVQdsALvfHL5C1kPSr6WrIgOqG
VeZ3rZ0rmzwv1xTfyFm1E7/4SRL3rfNorQiTInocoqYWkXMbnqS3z2sTphcCKiYqcBMorJd1ZdZH
yqYg5lhkiw3lvqLS8lN1q1vQJzfRQmcdDTbmbFDROp0uH8PRMVtE0i4m5hlqMhM2BA2u5xLVIcef
M6fg0rPujtk9P1yhxwcrhLWpaxfyB5/ujcz9WJ17KYecOW4iUODTo1/wa9pQ6WXUhTMp4N2yvBTS
KAhY+HyunXOupmDAtXSftugtAmi01NFBOxY5AdKh2cZyaiFFEOXlsh2Yo427vD1Pdxlw+J7wG+z3
eBtnWSFLOa3W3KEUsW78Pbm5zosTHH3Rv9P9nVXUTiBtwZCwHFoUF4c1LfSPlWczMAWOlyyRqOUH
Fw+aD3Huispj6tiq0gjsKo0yRfnhCR9nOQuOTpEnQsb5x9Kpc/dSRAh1dPdyRiQn5i7BDH4mA1PB
2ysZNhRi+J1zn5Hb0BaE2LESlmGRQl1Zs/ujdZEVxlCoLnv4aHBj4XdA7VudRJxqQcM5ypfnvDaK
5BzHuPhjvubpjbr6gHmB8LWwcYXAtSdKZ2qPFzL/vt8YSQPJRdHq2YcapenvZktPXNriwO49nn9d
aQUIEALiEYWIF9IUxwC02tPIAXJYv/EI9T1cnBXvXS65vE6LQepBW+8XmrUkrCoprvciUI4HqPBn
wBVF/rum+jANwjq+gPxdj0r0o1/EXhBvH6kLXLm9xYNi+I+9cZjd6IWRzDhe5ZlK8G9Cwf4A7NnP
8sTI40/EO81OAxD7DRCoY0azHr51DrrsfQHDxTs3UrCq82pzce4V1Ez/Z5rQXxRUKB3PDhXd/DSe
flKAY1Jx2AWMNO85SNHLgP4efQJlhy6zh2xhv9lkBbyXnl7qyfpyO4NwHBJsy8+7dTnfZrYjFzM4
C8UVPm0t5WgYkuBcq4M/ER9fDHdzcKn+WiSPjzXz+QPbm+lin8f/6YLrD69VIUYxy3/Ndb0Fj73Y
GystKkK9Q8RUYVYVwRfab3exyoasnE2bkCBpp2vHTxIP3DgGLyB1TkFG9kvxF1fUf15rXhcIW39J
wDu+3Wv7jETpCk4VgnP3Fr2X37miJJ58eugxVg29GAxuqxy7HiTWmCoFPQe+GyiDRp/+rRvccrnB
WRvE+7gx46j/RAzYhPWoTd5YqT4Pv/gIvEykRwRqVuC7N8+Qi+RdmCCXHGCOSwAsbxVmN53NvpA3
HwhJYYwRu/DZooTuQjlLjqwNEgPQToGOaFt71/JwF/C2nM3mpI0DXkAgM8qFgSzQybGEjhYVl6dK
FNgmECqP/8PXqxVwHfr6EnHWQvTjN7fU9QPhmIF7V8XERlSoacEOJOF5VXzi9/KOQwbULAZr+yL5
Btb0ffuVBjlBX6/lFpQi28A/tUVARILsRwytZ5DDRwhZf8TAgRxH4mXG0wScSmjKzUm5/qhQ0MVy
Ip2k8rGmA/77tB647X1jP0h8g8ymFwELxvGIfi9AKFmOaA/1CT8XKbKVZYf/lE5NUvp1FuwAvrTj
IS8cOC7DKs1Bxtmi4+qdqjoUiLiu5oz6ShRZpcvoUgMyEiqaI9+I8+c6nKt1/j82S1OggzIYAmam
J984GWsql4AJJsvoPONIIWrAbUPrwsre4Wjosi6Irlqr/SMNPbPT3b+L3/Aui4xY0Gz4iSNfsLLG
518CNG/Y9iz1M+QZn+JCQPJzGZJ0RlltvyMVqosfttplO8Txji7tPjBSQrCmd3hbwZ/ZIHWtvcmd
eyixVHe9VTp9C3WLKZkQP39jA3ggmwIt69wbA9fhLUo8iK3KnC6Nfo3W9gHT4hHmtMTSa2ywiYGH
sRLbqqlA2eF+2z8KhOOgcZmSfBS68dfPYvUTqfJ47g+J3Y68h/mGcbI22Pk9sdQDXEXf40QpZqdr
oFAM3sLUTqLpx9WogxYt2X9nbNnbYrWdQp7QEInF8orqcwziPpFCtZ2nv8PHGcUjLx+NZT5UD7BR
EZKM+MLDKazAapJPdvbDxJ3at/km0x9mHjSjYev1rxYFRIdUKglfoOwaidNGvoYFQo+LhALAyWkf
iTIYeyqkP9wZWSH4EzRD30qHFO/IuAL/u8zp5UP8SEyT3DZa7N5AI5rwvuFa25saf1Iw0e0Jdndg
zxNaYctbrmtlO/qHymQyhbxiPu2RAYr/QcmpEi443Coj3lMwRB1VGg6tEhHDEDszzCDw3kF/7E5f
/j8IQugFRkLJgM6XMTkY49d2rgyC142AvMvfoS5zRe5iFeflmjeKmchR1rMZHLm0mPE57y2zQleR
S76jKEwl5jsjmIOAVM5t8yxYDYWJvdKqLOQ/ouAVcmgBAMTm8yioj6iddg+ZlQJWMOLCf6TZgg0m
olzfU9VVrzMen2QC4vL42d6mxMWZkaqZYe+2h14ExzI4YLPU1AZvQ83c3oRmGJaxdc9Iavujewcv
kpXWxL/WBYXzMjUbRycARXjYMiWUopEMR2QNV2Cq00bw7m3CrZktCmvsMOAw9RgzURPlKO/8Azsk
O/Rc2dce5KkuEFiEb5QmkSSAJGHYmrpkksGu4mOZym0iaIo3gNmJL/OwCBtH9ppqc1/7zVpEswd7
RLx6Cz4CBuWJ8ULv/gWoxHFh0v6h6c2/vK3/5zRVcASWu96fYsA6YgaDAplCYAOgAnzZDHCStMlU
ibHwh9XAWuclVQjJJZzl/uN0+aYQ6wCvB0LTgkl+PWa4F9/Q0emes6riSLXMvsHp/Z0ElAj3dIrG
DKANjMtUni1d/pkRzS9Jzy0cZIXZseIGonyZo/Qpw9/TFbxJM2r5BCZO7sbv6XIhSzltUmAyBC6x
FXEVzoCjcuJHoi18djpv8NvDVCTss4Hf5URSv8y8SEJgwE9RQvuGg2nZO1S34QEwLFUS24tMS0LO
j8d8ztfEA/6vinxHFnpMyz21PIvOT1iLIoLord40Q+O10LIoMKz9vn5HNl+BFURIa1efaNGE6Pz7
93euXLUGZypW4N1tqqsysxaaSaEQInMB9kYdIWrDr6b+6+4GfYCkLWEGgLyR86pJ6caf+CQ9Zaby
d7USQLSdaEuD/5wmCKMsB5js33W16AgOtAFvJtrvTbqytymq06HiGm55m2eFdH4jCRCR9OHDE2UZ
FlJh6xDgKxB0lvv+yh8NrWXYJ9I6lYaAmc31sYqX5N6ik5dVzAxBOAv+At6edQ5ez6XwT4i/ISv3
ksVetlF9SWjXZrVq7o6yPx1Ydt0i/Fa7Yqxm1z8LSaQO3+yi6lf8U8UjPLbJWDQpQ9yHs0/9RuUU
h7Grh6VXHVV0i7ILxKN5tR7tuTD1FlQHXADk5/1/jehvKkVNkUUFiXkRIn2CYkB171bmZ9jDwM+J
5xPlFYPDzeEvH0tQvaYWp3HX+1tAuidxqCAPBwpo7zqXrKFLwgg51G1nbR/NAl0E8wt1UPEcBkOv
qC2sGVxkjoZhi1orx9vkD8pYWXcLFzk3LYtxQibsQm6JaIqqQGAw4tPNQwOd/Qf5QCLoLRF0wHz3
ATLbA246x4tgBpves9cza/X1lp5Ax+S68mp7mdjy1MQNpyIrVuQHvDCM+ZPZY3nM4JrbwEf2ucWA
B/D0/7APFy0ZRFxrtfxNh6cv9dSP32FBO50gMX5E0O6JwBQ8K9mtVx2H1n1gNhjQHjBRdG0EHlvf
NXkpvrzBUMcbDDZLYZjT4gVbRy5DuCdtdTeVN4j0lDIpHceeW+V9HbwO/XrmIwmYYqylQFwE9kP9
vH+2xB1IA4+9p+6FKf58KJ72qi8PfkIsTmKTswEF433oRLt9QDn37ehunCupdzMdSVyiPmTRZZXs
D+pSew7RYLwW91TQGZQkNEIwTbgBiZW9hd6MRBBWZmqy2WMHHL/nzOSOShqJZJzd/SfD3LJn3gbG
uk/bdkOy32Zpy0Uy0jg6h1qRPs/vA5ixzWw6e6vzMrrR1MdwnpRpyNALVKC+/51depaDtny4n+Hp
6oA6kxWEoOwmSTZxnbjWfD5QSqJhMvaR2G9aJbJdl8K/r4Kcn436vfxrxIf/K1fgfo42IbW8icEa
4eb5J+Z+ZDiNo8nkgqeiIJj4S18RD8T+TOh4PrpH6YivZY2Tz5qh9MVBUpSnNLNFXWNLXMOYTvik
N8RxaHoJDsY7wtJP7J63Zr/RmswYr/C6sT4tSlN7nUgMUVOdbONrSlRDtAXCl57WmnzudZblZ1az
6cM+LXJQytuKluT/q4v3jq3k8/xMT1MlN8s+9pz7RG+K2PH2E008qahZ4YLK1EhhJuVG698sGHZo
J2GtMZf1V7xMqxWhCkpteEpkpaFfq2BPND9Gaz8qznEVLK/dRv7XdJ7Asc7KK9m70l2h3fvfOoN/
5+jSS19IWpZY0glpTQJLi6H1biPIHV0Sre5+vBu2/iL0eQ/Tmw8CbqyPBSBlPylM5KMxn1bHwwRd
wEBxIpAQWsqxKd/94D26gOp0K1tlMc9i40UvT3ied45lRzUt41JqmxHA3qeDxDJ0WknJ3mFyIMvg
boY+EyuYZ3Ip/4zQhqXkjEAWMuTcdugdEB/mVkL2/mDkQj/4WVOAA/Qkt4vl2YfQoXuP2fzI8eIx
28kDD0Yhtu59cr5c2GwV1nt2w0AHZcCo1wQZJ9qejf0YaOFHQzY0YL0eBd74Af0YNUBY6ihosOyq
X7DEReQWIJqy6u+eaGegiVr7RuLP+eHTx1dmtCd3UPQXK66zW3DzZKO8lmBOhtwYqKdcLmD0cskB
9iOBwL0z8COSHoISrArjWoUIJPhWQ72rTG2cmWeFc4B3ZvLIixxKSRt+X8Iu6BWbFnhgXmJqyy47
FhpuvK16lj90+ak3+XUQXyXrmwZkE+MjHbjzHAasUUELvQa5AHeKsNtx5MZ+RqhU3+b2qpQnNlkj
8QT2LGnrYKMYgG6bTHyjHGnxUMdvy8cusfSxEBsWUS2YlaF5+f+xFj8AJNGZpV5id8Wtyc4MCWaL
lAOy79O4SDUX2iy85UHPnrqY32c9WL2p/wF0VGCZXstZEgBYjR3KK7xBundUVStr1aHiM9ysPVIK
OVSdz3IYBN2w93hGOusypQPubJEZVkTCgrXbojniF/DxL+V5Nrbm/tzN1jf+NiDCLxL4WBTpJPwB
SdPtL1PF3pQBwdS1T7O69avuGnwAxOWGFucysLv8Fj3wFgq7VZRAu+yw+BuLj0Mh1ponNuoJLMa1
Li5hNhb1/6JemXaTFbS9i12/YmyzMYmD9974otxq46wmIy3TFsJ2pwK3wn/e4exqPphN2c/5FPnu
B1BQMX+dAwu5zR5ix13Xp4UaLa6W3sMw1PPQPodg9hxhQlBbITBEFWnqF+atAgcfUwtD1uJAZ56o
41+dwLwqF54U4tbFktihDAmeFS9XqeZVT2geXNlikFPQXua+I51D9lV/UClm7WLoCh4akHVqXQG6
v9yusyHL84o7MaF+85w7YWYUo+z4QLxomVV6SJnMGc3D5whqzEs4KsqIhJjryXuGjAvkhNtCdPr9
FxVs0rW4EnfaU7W45L9cMOCTy+oXj7U3f4Uc8qG2D33/2HhFX9HOm9NyM4LfVfj4wtEtdDNUwEJ6
9iTpRAFD5MKhaJBpv3WM1dr3Q4gSGLvdQO5ysNgJlFCLJRkKNSxqQiCv4fyUUnaR4+dN9cuawIZ8
gHpgsICdcgMMjQburvmYmdg+tSxcbGFohQ8zSfNR3ojeBTiEGGUJztpmkxdq0gdMJYWmg/luS4AF
ljIIS7WeRQXU920fx4drr0GEDaEdKb3n4MZpBlIVmDrAhToTUmzkskdbFo58NMEDvFyzEnhpn7es
RIVONCIA/7nVE5Nwy0Lk7BtyWJO2wvsx1S8XzW2Mghd1417CWeELnaAA+gP4pnOZ5x0uNQGqwgOw
9kllmw/JlZgnD3SEc51UvBKD47kfcAyfJt1MR3Lkn5gMVG5UHA3FkOOaIEw21gy9Py5od1YU+cSy
0ErkOImD/73D3Wcqbn3EERZAbUM7yijAkHBUHPTMrf6R4Xe41PC3Jahq4SIbCdDBAkKvS6CF+BB5
BdPRtp3Rq5sMt6toj2Aw/e7TkXL+1wGbzLJ8LmNVV5+vwDbz96rKEe8snCK2/P36YCOixIENzgQW
jySTkz6j2ZW8ThuIBrlU6Wyw2iL+ZjXm49hWRNrRQhtEZaLM1neoxg4P15b8+FOF5MweqsGMpzag
YG03mFzo4PK070eYEsNYEjMNtYk1/e0ji5B54C1z/O1xBRVHEksjEuuSCvx4aiWkY44LzLgjaRcV
Myg+jxXqkNQ7ibyFxUfJU4dbPRBOl/NWOhsxvXqz/5RAsF5x6OgxU0ZPsVwimOgEu03YLNEBImHq
WvbmuaRjO2OA2OcvqhkRMfhxHs+yTufT4N606Z19FgH+wSxGnchcS8JJV1CpbY02CRY/jruo3/Ym
ayWJGQBz9r4G1ExetnMcGpH6V/XE2Y/3QzSMXDhcK1mzOgWRG08hiGSlmAUGJs63ixG4QmN7qEbh
g1UEjQ9ajk3qlKfwxSLWsr53liEv7vbx+8gHaslwpONxwkFGER9zPfmpGNsWrrRa4fb3cfiExki/
in2VbwTleUtXu220Y0v8w2l9vIjlX5teoD7P3GzrjZYZ8ixN9Lb06o6SMBeeUmrSCI06HNmb3XR+
FNqHXNVi65LyAg1VpP6Pi0warTiyIlqJy6DTi4ss3R7H/w4G+J+V+x+NEOQr2SwoFeJ+preYPtGY
OZS6C+5hfhMiz2YFLeFoahOP9lAy/iY1BZsxkFu5erKo7lzZEk2zNyY1/h2OY2inXh0AlJUS9KZf
fP9vgCktIMGtqq5KDvBG/jq0lUztdUridGBPEgjSk8EyRsJ8vrzSALDtJCOmDidKzXq7j7CoevJk
t4hTQTZzL5ioCJoeVjY5eclEy0EG9YQSkv91d/fPipDKokQ6QTutwJeFO8WTN8+beCz0pDvWBUkk
OA/fJCmye/of/bWQA3gYTvsCwYGd5TYvYiZ6pjUkPjTNQWsB5K7RhPQh4JoTmK+I58AYA+Y8xETK
AcnjCR6bNivybikrUZIRhNnyLDQk+zz7s+CseJ+P2ja72zf+inqIgqYy9sAmHpA2dbG7izq+/O/3
+H5TUlq/dUv6oSRvXNghpI1nl+G5E4iZYDIAaEmvA1jAw1+8OeXjEaQSKNlBNxOVZ/D4V7KyZpux
N5UU4vvmZ3lDB9ixnOX5ZxQDPbuAsu0CNfW7uq7sK3vEY2UEmmseWVwOGzDF5Z584acyAr7h7A+C
mbrnNcjChF/pjndp6yhJSx7xH8cCL30883tR3tfW8kSl7IVt7QKlWNOsyRNsXZY3Z5I64Ynwb/QL
OCvl5WC1HkVTCWxxSVpQzJNPfu04Y9MVPOZZmVpSs4o6Wjw+79EfCb66PDwQfOzJuYvTamkiXtyn
LLpndMwqNiaaVmMltxIsxeNGAypiCNUkuk36VXg0ZcMQZhZPFUf3X3Lz46YmXqfX5wz13nb6W4p7
o18Y4rhxCIeFr03PE4PNSDoq0lc/aBBIUBShAyx9G1ggf3skW6qEvKUbFxD/fYM+QCk5wre0Zgsh
/LjsQ3Ry+rZgNL6fAGa8pKfqF6t6/3q4qjRLBv72rgReuyANNaKtvkYTXe5jh3ThLL9LLDK5yl0H
tgY48ORMIjtL5zWWy2kf7LFSaZnP0H0ytVt157i8pg7vwNW3UAxdd980Pu2hMtb8PR5YO7A8TD7d
gTQOZ06jnSC3QLaCaUGlXAYVoWFOIvpTKtHfFmFDfCCCrkyc4PRTmntjWvBKxsoaophi441a9hUq
+UjqoiOWqMwEmA89xgQtlQ3RujSZ3x5B432cFvNA6ZbgFkO2N0D+oq3PhKjPBgvbzm3eYK08rmbw
Mm1x+KE2cqDUPkqk0Gwzc4TWhkNotigfAb6LI7aUhGPE0CSgKcTWc9cB9463RA1VQXJdq5MsE5+z
vMJ8npg5itNyRhc/kiUfDPGrjUGcx9iX+/MKomZ+aGFDbuogRYiVgpQP7IzkXRCMoLhScS8WENbP
HjuVOPWZNdn8BJZs1y1TwEue0CTZwjcdjTv3laJ/0OEMt/ETs21ANfSrariUOH213TS+QZPCgtuY
0wLN2693XooF3weF4pY2xJH/Xf3syuKA09AV8oDI0/vQpx+fGhXT0Kb7LEuA3o4Mwthkjp8MrchN
rFNa3ugkNTQlOoNCl3N7mkDXsj2kCjXgTRj+vIlA6N9z96uUhl8agC8IkDOeZPb1sN49xzuih8Mc
gRD3IbJRHJnAMDSr968TQ5AUrDo+Ojcbg1yHOkAW5/30rRkWfaZRAGrkig1pBHbN8m0Qwgs9V20f
4oxImW0wWgfpOcWFVKHIYfXCSN2gmzEHImLVKqUG/ESxFSQXzIRE+eXeZVlCY7APrxaI7K6j0qCh
rL+j7ZmMuawk1Izqh/Plz0AYiBCtAjpyiZ4DoM0MLZ8nhHGApONmfAtVm7tE3vh8rPbqCgpT3dwQ
f/wJ72+qgNWWjxP0bfYnZdwCNB663PswaZp3IGGG83MmWHHMmFmkGIYrMkjn4PK/DNHoawNwP+br
Wr5abNPLVnrCfMnRB30luvk0YY1v1GWyg5KRKvYyNpBH6xzOefctaQNtzx+uZ1rITPAEqSVMRk5v
iPtf50+mYgL+xf4rAPy79xMOYfRH9lKR0wFLsuxBnvFSvFUWSvpCzEOZADOsZFwzq85AGMHEArk4
rRPaS6C9nvS50pX91hGalPtNM+VRNFlHRcY9eiAshynQDZ/N6cnlQmbcy3u2YwmNC+AXQi0wxNwT
kEBgHq5V74AdBK7pMJTaQoV2CrXwSA3o75eP4U19WtVHA6/hOvLuZ7w5YFkWcoghxZllBDb7J6MG
+wQh1hCQEX8FDdVwx5XBbaDEUgLHlAuxnWQHr2r/qU5dVmaukDc9mDX+thtSI4c9RMPzJIMhpR1H
he1Q65mLklX58oVUUmZV4X9Z8kY4czZdZldfth821CaiqGeA+2B8fTJA5AZtdh1QsukC36GXRz/6
GhXcdSv/fY/IZ9GcbYS0gIEEjTlL3F5rrs8thc8eSTKWs+BgTiEx4ayzjgu/zmJRLqOYQWQPBe6v
PtRl4yx7F4WLJjZUq/67vOxztKgYpebxMBGlrxY778m5/RdpCvd0YNXbA0+6iWb7JRRAPrUDjHC9
4t8EGHYi5LtWVkluellXtkvQMdyTr7TrhI2TJkQ64C9F8F/Lw+ZjZKjQfqbcSYhuqFhrlWdiIYzG
RMhhY9C63OdwcIcz+Mm6peZydM25/BHIrMdI/Sw0HEwIwf6pg1oJftx2kkiXPk7k0t6WK4xNYWgw
LtYUsxpkfRCFkHm4MbmMQuAfQh+l8OFzDdT+DM17ct7OWE/msHGDoOe4gQKSUf3itpyfS3Wgb7Ad
SiQIu6HwNP9js6J8tPvPrKunKsFZBsOBa4vOVgyAMcI+LvqO8st7sGOl61peRdSZ7y4BVU3WVVYg
04h6YO7GrETzNaUDkOe5l7H8HwTpUNGB43IqlI/xu308Hj/d70TU9vmEPzXxrQiAoz22sIdAVJ4i
5ZlIgd/wbC+gOf1RDXgUcoVERaTSBCn6MM2pXVs3MX4YaU/pdEJJs2KSiDiDBw5/c4GStInYkGXh
NsVRwLu+GU5m0245LAsqThlePbsyK5eiHH21S27KosrMFiJQQ2EkSn19tCX8gKIFrniUqm7G/5F8
galgr3evcCduM7+7mBMeevdBRIi52pVa5vxhEbttWol87Z5QS3ywAKpfjhO+uoTuhr8M16ti0Zxe
GfgB4v1TZXHU8P+2jff4r+PywsSjeEiu+rBbVnUZn4koQcApcT2cxK15Qz3+ljLfZDhrdYq4bhE2
U4Q7vZSDyO1EFI0u6+Gqi2dN7bFibg/GzBQNyN6ip9dIp8k8/zlZj1v2ln6sGTDTK5WgP/HftAQj
yjgGHBBdHs+OHtnNipG/24SB/1pv1/iccLoiw/6roz0z6Jho9Ql3vEQAsJyAz3u4diR/r4bezZY0
ThMMU2+cqt6e2wNVNk1OsMd7A2e80hQa7y4RjPVFgB9Ez1bLyVKnGY32HNZt0iu1h+JSCQSpJjsp
KMAPNZCPJdDRki1brgskFjjaQMtXed2jGRukegePoeUqtJQcwYQjK7DSFnBnvMDThoP0PmWL8HhN
G3VUrkoilc4uLIwmQC8gM+MlKM3KnKE2SBaS9OpODAftDoOC0Hp7tZRr8O0lEaxmBBOi8kcQvh7C
Ekgz/ZyGwbmYYGSNOqBGka1YelR/0ohw0uKNA/yZsNpgUxETVMV2lNTN76jRRbFMp41EvN5KgRNI
1lMESIE/jseYm7JfB/UpE5UK24lBKRlt7N4BRgFj/YW3Vy2qtALaSrUGQP9vqFr0M5oP//UU0Odl
pFw262d45/hyppVyuK8Bye8h2HiEO1ci69WcNR3SpgXJryqSsKEpda6LGF9wgzKWSZGyS8et9ek5
zvTdfkYAwTh/zj0u6dLDKD0IlK8fQY0y4oH216sxkqvu5snLeCePJfxIAaAH0RFakhKpOxqUhYV1
krCBPKBlwvYcM9r5eFzvDTGiHff/DcfB8iPDKFA2oeZ4TNijNan7iY4Qcff5b6+QLcdntuSqRaRK
Nh3MMvJvy0I/oXkpquOUOcBao/UIDWm2QJ6Ho1ubKGkv3Za9qoR+gl/KcaVcLwSypLUY1WMSuIxu
tVrNcxwRwbp8OaI6+PbyO1hiOx6Opg3AsvHAg6jpMiiAgNuTH4Z67YAavaYpAeAWonbl88BpwANe
v1+ChK6hikLH3MVF9b13EMCpy3tugiAP8iH2H8nrL9RX+elzjSfLcy5px6BsNPdbDMRqS/hH0w69
eQZLk4iDvTeIPgf86e3CyzIIGR7xmj5R+jb9c3udCoDBdfw2kzzqUtgrQfmw9B6Rniqgh2Fyo5Sn
q1fVyUiH5A2RZzl1gl+Rliw6YuA9mE5NBvl+xf9cgwOhjPAYUITRwXOH+KUfBtkTNQxnjvEYqoEt
qjr6wwv+RDY57XqT+fKPoXCBFKXV1nTy4d7bQgFfP0xuHu3Z/ivzkzwGBStLvmyo78UghyljyBWI
hV6XBNu+AFQG55EtRSoO86dQoGr2zss1SWUCgCco+8/jAztNImjhmi3RwnvkZlGsoOfHJQ0hQKIe
+OYQ/JXZi6sFCJTo2fhS5QCgzByTXOj0mQ39f1M6magD344u2vzUmDXHQzs+GcFAr90o4p8kA8yx
ys8g/unH+lXYBugtnUHXjJzIfYb0bpNx9Oy0i9YgDil2Rbg0B3tKGMXDMjmAc5yK5weMUXD9YKxl
ggnprAp5RxNKGxoW84Oky52WlY+yFfjzQwu5uELaIRH0VtZt7XBDmUzYIzimy9kDaPUvv8DBw/V7
ciGHi6RbdUpjffgiAVpTrorFypyQo/o5RSt0ZxDlLrCzTrssp8/0JBn0G4rWoi4wiJAfrQvfniRs
waseM8f6W3wYar4lmk49dofbcAjhdXZNgHw/JEWHf+BVlfWEApO5dcfBzIcjsnINe1I+CiyMUEZL
RM+bBSSQd7JHPQ4Q3hmuiczFvHz3ury1au60zfIamcEWl/nHC3PC+ljugKsBfk+HE1aoO4Lx5oxd
Eudyk+be2sstc9BMoZkxZ08gL1/AWwF+UHIPVQxKLKV/KYTimFq35dKTSIzzJAV1nRZ4mpt7Bdda
YdIkbJKQwXOLlp8uxtsWh9cyCbYCK7CQjx9yZf7MOUq0RfdOSujpLfdtLzBORsCbu+Qqz7WdVOxu
SHy8OXxjMebh6Y+s0Jgx+kgLleXqFXu8aVj798mPz0Z4xQDWvPaPaB8DPcCEsKXKRZ4xNMzucxFt
s6UEwhS/uz/gJHLyTSVyeACI4xvk8owRPVwXvRRBbU1vHw9Nwr0HNEbL4rmhCAEgLCB4Jxsw41bK
eN2Dv6UpWJP0L6Nw/bvMjEZ/3Ql75Cy73lt9ZFVu7qOrQAOuRwpe5luLR6T3+ba4tjYHByIPfVz6
RDHAYvju2ZEYVgxpJNcaC+Nvpb7XUoejrChXVHrNpqpLJ+/tYkzykAom9twpCek1SuMcnbpDA4PW
pbAtJnT1k9hEmD1IiL3yH3SWIBHBfgF9wRTNqyq2DJytdQMxhe8ZRNJ/4YV9TIceiaEW5qi3Kqss
UDADOEaWob2060gahNN84By4FJI4Vt7ldZHyUnoKcjSOCYlvcO6hnk+cH8IQr/zntfa4Tw5O2azw
p5JH/XftpBxI3crED3a6QGHowPLXwSFq74COTVfnbYeyJib4a1GO7wIoTdD9rCgmWEx09sO7j6qp
rOJ/Lv4FxFBfcXUbViP+NWss/W1aoh2OnOIvaEO8JuMZRolprlRXUnKNuqt6sIxBGwBXJ6Kll4Lb
oakdq+XSCFi39tkJK9aI6DrjEEUvZg3xGBW597wHBpWOZl2EMLB9AN1PRQfJVGjmmM/bbKASNida
UWRtVF2EQUDeTpHkrQ9wkp6cOemSP0ZWSOxgE2d0leJBupI2XQlm+WGdkodIEOVeu5mt+WiiNBKU
5slS1GKOP4Vdwsa7SIprHF+4FK3ihYyem/20IhhELUkD7Y4idQw4pfrtOGMvygJECYkskIWyyi4w
BMXez0nyzrc2g46jsnmuQHhugY6gocV1q+ZPNVt1PctFq7SPv2PnUzWMbDzkL9uvD36Lo4dVVh3h
1ihCyDJ+7jSw3S5+HjubkhxyAxu+B7d4UvhS7nh0hwA1jOThHL9kTnKAZHIrhyFJX4IWQKMIB1s/
yjkkydClQnt226dpgyjYViUB3/nsuzH25o0cijkE0avnm0eImrjR7MHo8oHkrn3pNT0fOaOih/SD
KTpxo70f0tYtKHxy5w5M12EVKzf+GL+yOSTW4DUEmfvbnr1MYsuW3D9bSEsfYD0hlSvqWDYVn/gd
txxJGxVGUppgisZdEWhKrnNvRiYGrWXjEvUZOd5nFtQket+kTuuuQiUQ5rfS5KLoJZtFcIn12g39
rQiZMADMfhnhPBTJmfi7JrkRaH9pCHkRj7w9DK+7I6+6wtHoU3SESckY2t3hdWSN0N5qqxFN56Gl
DiW+ipTSVeN40HafeIryUQyw6AauE0JV0ha0sC+2x7Iyu2FZRu2oH7FohVWNnSJqh1LI3pnmhzKA
939WFfOU1QJbPT1ywJR0MPmdDJLV+t9dFyIMspamY5kLB5+tuO5NjcrnuvC3sYuMvAdJtArU4AWf
Y91QA6nrlS3wG5vwuJRK2Q27Vmj37m0s/OHzCKgeP529754ysf2TLLMxPdQ2gP5OCCr9zJYvfAsK
K+Zf/7Le7zEjWP+gbkkyBxQ03JJQf+3eypT+kpVaRQsHZ5RlaW1Ucq6T7K50TqRArQ1eArnrxM2H
I6wkBBBkTsP2IY2bmcVeu6wNhcypHoXDzp1dkEeiquvmPj6CtaumhtqQlPx1laegb8I848QxHwXI
kp1cOFTsB2LogbhbMs8z0zAf7oRPNG8QiaeN+QWHZt5TBQGKHk47wy9X3Jj7NalUhTDzwZEH5KtD
xm+NAo9REkPoR3yH8W7VQet29kt+XpiDroI5IBc1K6zjLUcFYeIEI1yFX6iMUuMP2D6DEA7T45KE
+GZzIFc0COuEwBYxbvt5ZXdMa/8lwHS4hrL7fg3yEVMdInItdeW1E1SML/TWQfEvsul39l3aUgi2
6Vj0ZvLDLx2GzQ08wNpnutzP5AAgSpTrSfFNT1RtJ0dVZ52iqY9QxQIBVGUqIj+hBoeZN/BOuV4K
YwAJUOoaLSiH84diwpCsOCK32Z5yVfvJI3ARzM+y32O02UMndw9bN54/vl0CBdFCaYuOt4qtSgBQ
LWVmajVTl0vwI8F7iW0YtHlgWBSs7lgWExdraPNfaePr0tlRpFPBq9gH7JB6ua89OfsXLWY6R5jy
VTJkvnA5cJtECxquOCX136ZZpwdSrJFkmDfcl2RDoAhiSVT6kVylcKibEVJ/1VwmXFq2Y96gvTgE
YIkhiR2VrteiJfuNoxub2KaVqHiEJN3jr8iwUDNX7xO7gx2TT0hhi5g6CY8+gY3raDCQ0NqSJMZP
Ywlx0a2mm3ZUglcKbpCQOmzT5HMLAcqB7FqLhtRXnS23UAuSYimUIe53ufg0QEt2sj3ha7YQQVII
NS1pwtwvdIIfAc0yoxe2ZDVbc6TXaVJvneUWRsywO1F/LaUihKXMe2QCRXUMb/wdLwbMGB4hyTjt
gtg1KnwGKf6yJaUg/5uNGKjzrSMPIsaF7NRki8PzTN/qDjkOdHui4L3qAUIQmSFtuzzoFlIzVcjn
NzaMCvD+tZ7xbixg/3twey/zTofYGp+7aXE0CJXVbcIxNTkOqte3WcI56EWtNeKGwUKuzx6nFskC
nPg3yvz9F4nIhGvVlgvtwHcjMRGGLQcK7yoah+cCtpn0h0ExuvfrpxkAlsHKuioBvyk2o2TsM6j3
gIf9GEHeKB8K+Xw7DgfU9nTnCMgPYY6pHkRO4SmsgoH8dYCn0FSbvWLs2nHQwF+HwUCoPxP//J8+
laBHBhNcaeYEfFehoN0mb1+DsU7K6zUH+26EQU3LJqDQokYUohcXHKmg94wA6oq7xU28vm0IkZDT
4xbtjBaBepQpF8Q+Xec/VcJdOB8RqfotCB0dSTQqrwbO5Vt9Mq1ogvMVMHBfa7+qZdg1b5X5SYTf
tOBwqpDzLLIYgKcQCW3B8c0fLUKn/SCogTJlAQKfSofBm76UNyTmZjQOuF64E81RNmMfAPvqukZs
uXHbMZAkFEqbZDtwxOuKfh6L25iJn1CiAp2aHUa0rWbLW+1bvhCvANt8ZP8MwiZQhXIS/q6JCtHZ
JovGkN/WFhBYTcVMLOpeZ36OvlcMNLTTFDsG/3Gh7l5DO4m9Efkl42OyYKNDuQzarjAW0DcQGzqI
a2hZxgZ9QDxUmesaktK1g1KKs1CoxyJKBnTmkBCrflxVYP9xp4BVc/4lJMAgRUeLNVOyoF0j4FtK
Y7NE3/Gau65ux3H3L1Uo6iFQJeJgOGAoYkwyiRdEjmNqA3OSc+bMpDBEsHMr9tUmqSWGzxzWjyP6
Ih8D77oIK22I7hLXwjiqsbXeSomrQs1S0Dw3iHz+/9eACrO5Kmb+E0pQS9d52jzbpS6r0ghxlNef
UkKzzxXuCVXy3PmntzhdcgFgN+CbZ5j4YT+IwRoLnIwA/OJKR/gZriSIfEzxnOb7cvj7RqOnSSsK
fMAO40EkTsdMA3JOLFPogcCiW3/rpATcos7bfowZytFGJT6b3vImciOxo3dfxtQmSFJkynGOc8Xo
/EN/h1z8Q1UodqXpSC0Q529KDqsxhdjLn2E0/oasy/r4AeVUv7TbSMD85fcRDg49nINfXWMxu0Vi
Pgz3nFNkWVgTrMmMKSIglSk/ZPBKUYhoM0uWRVhzddbtAGvrR17vnOIMnWWFGFalWwGcd2vLPUeB
jHWgAfJ40ItSmhUQ6pY58Xz8+gtt4NESwcBn8f48xRO8pcig/3MR+9GfEB+pcYjHgAFHvS+un7ag
DSOmgKzgrGROgzOjIBuy994uX1moGk0JizEDQWJFDPU9FLMQk4f8p0T8AdgYFaX9CAwab+onj/Cj
0vBu6S7igpxI88eSaF1vW7pdgvzoVcNNR6e96S+I1lgBpBYkk94XwdN+KV693+oLSnG+iZhjqq98
HJmumEgBArOt813IDolUQtk9EvyBZb41AY8BUhQX9ABJ8LFo+gXqjsrnLL3y+GAZy4/No9/bwZEw
k7JO7SQJH3HqegBZNW4NOTot6m5Mg2JnFuX+XLEjtXkTHsUoKAcrI8SQZ9bGKeAu1Z3zC0xBMQyM
RGNGGdfqr2BCzoVLNF/zi8Wbh3++otPXPygcq9OGpT0pC7gJtTYKrzC0mfqQFcQZnI9X9vb7VxIX
8kVpX0oLy+7twy4rvaXnxPjy/8maeNfXJvd3aSVVtI0IfrK519qc+GbqRMwqF1Pj6IYMnOa7bnFe
b7S5oKFUs+RQv2UutCVzdE8V3RIPoWiBLMHMVwwQ6OCUYOv3jZijvZKYn42iCVEh4zOsqFeiKcGb
9qRQAjZ7rkqOOWRTcWptfXZxaNaNBQ22on6JTq9MihJ3L3m/XpWYWo94V9xtWGI5VyxyFgZw/2+X
PP1E0Wx5oX4eVshhph+U8DEgVY4+sIGS3BXZyWHVaAYQEhjvnAxzeT4aUn5+e9czRhrCjDz4F6HO
qUEjrABt2zGr+nZLfuCC2ZFjGOsyVYcXdqtxWUm971OLj/Q+Yrujok5xcYrSrfFgeErvB5N34dLd
lVrqYvYWKwJBCtwuXx6LfM8QtLKYCb//gQXbaTXpaK4DHVclPlRluW0Q7dG+nxZhE6nFfhM+ymdV
/KDKBSa87TmIS5LPslCywZrLAce+Be8sp2zcFUXaSorJdhc3B13M7sUXu+8fVwYH34KfxtY3q9TF
gffotKvdkkoNZ691ZLs+qWOwQFueN/xo3cQT/dQDyqIQ17I0MyjOD3A0n7V4msivtPXez+xWbKO0
P7L75b1icrLsGCi21JgSVfYnIsuMgFQCNkCPV2cQtBcdQKrHqfD1nEu+KVwu5AYcg7cy8hP1+mwW
fNwwXypZlL6McR03zQID0wGNOfhIqKVwTypgZzU1YCwpjAuue1pF9zwkhA14iQDtmKq4NJhshwgt
X9jZL5549phPI64PrTYnasbi3hhQvO3RzUjHZxPIjya+fezHzR6yPQgRVTDpuKDKFVh21s1mygh6
777qW13+CbO0EsWhS8y3NtXiFuzQ1U1PKd6STH0HemZTxnMvuuJrtcmlYMU+tRwYJQjcCgblrTJU
s/EqC2yWjf87mAjZM7X7+PpjJyKy7x/5UM3ZhrQFta1iY/LXwRnJKAKEXaiqcCxR4CjhmoVlKgLl
5evRqcMJ4ztGuxkfTx+4PbjtJ39YDVfyui6pF+DhOkNS7yHJ8KenqLTpJsbudHee9+CLAqUccYHU
kLAxIm8TGhU+CGayPo+YAeuNEcdFr7OHQO9mf8J3Mq+pvjYcbHN5TIWq3vyGTPaLdMEbCvPonhfs
+7wvbsr69yCWJtW/3Dnvpfa5L2uZ678vOKMnKGYcjPqvGXZV+6Cfy/QHlK6bX698Z71SMOvcXGkD
w0Z/co9TZPtM6zYurp+T4g1QdkMRJtZHAytb25cVnGkQFIrSe/8UefFJPVpoBEl1UTcVbVwK8qVo
VM8rmlFLkr5KUI3U76aNH/bZYeGH/fpWzer/aLeoEcLrwuQIdJYQCQziikZ3Ug4zKTuKaqYf3JHP
KZTKUHHIPa5dYSroDqTv8uUiT1K7+yJd3Wqo9ek72MQnGl3WZdCB3nK/Gcb/w/zFXCzdN/1usYFB
hJP/3v4WHiJHC/lhFeojTktMtI1nwri5S5qGDP6TXU6GvSXzPtU6ZsCqHij+CfGGnO2yyJDlXBwW
FWlhKrSVD0cMFaoFaSrIp/QbBO2CmeDuKVRDRtTyOTzXEKA3LaTK72DC+XAD4Z1YllkJASeHc1hx
OJ9H3VMeswMcCl+Tm9CbqwSwzRJ9hRLZjiif6P9dHVSEiTioyLVqWQNzufAJulCp7erQVnS43pdt
BzyI34jK/biosog9e/oSggoZIr6ldxPLqkGL2JZcd+an+a3Tx0NYFvcs74tN9rrLlHc59wm1k8ik
7vEDL9GiW1PuFhR0HlR8RY0afqVMcv7QvqcFpw+gkUwkkKCdReEk6Lh+gA4ff7OW7RQJulMwR4fU
fI9fC1e3rW47JndZDOvfGYXxgs2weiq9SHdl75v+YILIG0QfjWL95bEPBS+LK3hHdOi/wuBv1QR6
ZSoGTD99QGLyEh5sXJSQ2EcUBIH+9xI3heC5r0DDN0c0sy24w1G6mQIRc8NA1xlXvFS060IEXNau
NaOE4YLujvOEg4WSOismg0fygsywoZbCrgr08Zfuv93ZPnja8v9gWtauW6RAr5FKM7yAL05xtXb7
MM4yQl0id0tyhrt1LBGpxy8szLTBHKhZFT5dXWqlW9Ya26FjgC3etnz+KUdYCehmRiL/qO2OIsBD
yX3w7y2TqrWIgQekIbHF0SkM1FuzK1Zyv5c7F2VsvGt/Tci/wVJJqZNOaVa02Hkh+jyO0Bkltsmt
uApBNKqW3Ai9QOLtU+POB/4TPY8aHMrwhW3OzDLaVO/E3yfqu1mY/P0WlJvBD3I8AVM0YVmstIz7
f1nTdS8ggMfC2i+hMRsw8hjNGWUHshmNWvVEnET4t8f8Ax86Xx6jR5zOcOTHY2UzoAdnlccxJ+fY
hwQ2dwk539PqLCRgK+3GRAJW4ow243nSrbFIbMd7gu2C3OG9MFx4N4wKLhyTM81Rg3Mvy0tH4wgR
cMXbd3J+z+C7KmaTtJD5EOUdlXvX2H+HpLR340CHb22k/8vIMBGm0M1bSXgVrKYHIgP2ZxJgPkdA
KOpcHFaZe0OdTSe8a7WmKRdqmUQb6tu67tI1cTQgp+EZPhqxb74CjtxqGABMkAKNTFuULVYVZh8A
HneKT2oGYdIlV4jbtI+A9JRboFJ33rAdfKTvXmAtS/GP0SCMBUvF20PP9W/AF7AluuJ5h3BBZjAx
zQC/DfwxSiZH79jddejFB8omZMrjtFYUZWgEeEqaq5jkDT6DsYcgiNjMtMCgiL/X8MQv7DhgVFD/
ZEYfmW76WHmP67MJSrYATKhC3e+shV7SDcVoCdmFixIaO2swvdvAFKMUPatck/jbSAfV3Iburl4a
xLy6IckK2r1rnnx8PoUDNky4YApB0uaR9rUGP9oic4ZRWs4n90vGLVtiHnjhwl9efcD/lyMLR+qx
AqLXdnak8jAY8b68XMX6tbfpIwIRmXp0Uj1oGW95FnbOF1TUCbLJIyD0EDDszp1uYuIWwn9RqTT3
dHLD+puJEE29jMbtPCRc1lwuiNP2kg0FarYWCckAAXINywJyNLRfs+mN13/IgBOi8PUNpApvzQv+
ISjEfn0jTowbvwmJT65FZn+j11OiZQabbnJ8IVYRTg/9Sgsh9wblfRj1aWtJypVjOlKg/JAPEmSa
w3MknSLpV70fNpbPy5MjVA93F4zWJuHZDns+2I8uq9XZEydT9p67aqXusIWI4NiixcRoWliMYD0K
BBnwNg0rftTdAlbgdd4nnz3Yk9yjgIxKkiXvJK6OlPuOJ9W5eXeyJOyY6NfoTZZbb+0mtaKov8ZK
zrdVqipiHmo1g/JENB8JeCsu6Ag189mFT5TUUnDIQ/15+PU3EBhvc5IEEVnVtyGUFth1uiovheem
otuczXoataFsqNPJsdoWWDy8Po/sHWN59IZFmC9h17UGpLIgox4ikvVjSUwwXCRopWqGxJsir8n5
TY8qkUsWZiywjJsxLvraWnBw9vcvMW92iTBgMjfZnMJUFy5WQkX7ZNemv4HdNH16TI42IR0zlx+m
FyVsarsgmlb1wXR6yB82uqy3R9j3Oc0kYfu0wr6fH5yAlz00ZD24z8Bt3L+dKB41uDTQuuGMVPXB
8V3E1UFZ99PorChn6REvn631eRT4QSu/LYLUOtt/0wNpi1gx7J6B8J66Ie2Ol9os2AEFpwznAoiF
4tUzAMfuNN3Mh3Zk2otZBtc0Tg9RA3lPsieVUNCZYtl8512kh5zmqO4Wq3328YcVbfzItegWtdRo
D4+gmnIpeCUIusgtO0j0POP5FOCPqT7M3ZdbOT45FaE4S1VFEACPph/cxdRfQ1DB9hkIi1QzFyKK
aoQEmJAAl5JfkYiX9saqn+kTwi6PPN3vVtuJCoLMRxnh1sXJLL+RuxOIamt+YlMmOaSnhAyP/oSz
1YUDQSOVWbWM62QjvGOm54ky6ceDij2dLHctJHe/UBlPcILP+fwQhaq7RLX6t8xB8osk6U8lF9Fm
ADHBif7kiByEXkIN7ECW4yXx3xvZX0xO2gwdQ1L/q7pTRpBOPl8EvEgRqj1CmefBPZ41jb0efzb4
La3O3c4LH6Ir+05KhjHctKX8DZQzF+5g2IhAOp5psTYI9WzBRRaRtjlrZngsX+IAPr98iDokzaRZ
RBcXcDoZsPfeALZiA336M7GImjxE3z2krqrHU9sQ0U48j9KhB/vwjparZsWnVQdU7GxTcfMKbvqa
TBZZUkjr97AJ21R6zb60GqMGqUHv+u7xDCDcs90sRL/Pc21bSC84ijwZFabu/Y/hzkjVIxtCSsi7
dVjuv7HAKMQFWBBfm2y+U9igMxPGDLaAqoG9hZJHCve2RLnB9Jtv13KhQq3ipdpwuIXCglX83zs8
//QTmraUajnRS9nn7215PdLspiJWmsrwbl+A4kne4ekoAF5vCIvmEYSKWjCRt7HcDMXOgV24GOEB
oBr/sJbgOghnyqqVQmct1b8Yg/+5YxPv/Rc2kdsJfnZ9qKCC+QvmNT3rsCGMlGikRTz9CKDQCAfp
HzFisAhK2ZLER2LMWmmP3NKsGEO84UE/wEFbSEnzKTptTmWn4BWR9pBXBizHmNWLACuJUsoMIFCR
GMhhtunB3c5t7XVR79OPpOI0CFhbFdXaT/LkC+l4v5PRjNXZEgAbERN0bTXiIPsbwsEkPEDQoiJq
4XWzRAyuvPnxx8FZJNpAiFZ1fZYjr/YuQR3+0ybCbS5fCWONOH1HeBHmnjGkwVIE7B/DErnm4+/a
KXZGjiCjA5o879WSKBk1Ar+xrUJfCTgXkoxgaL1/LlIZh8tVvIr4jxhxhX7tMY4jdEp4Z6sbQBZW
5zMzXhwTnwA2StVBwea0Rzleg9BV/9kJDOgvaQhLiaAcNwQSw7k7L8zd4wxZy0JRzItEkWAyYbDe
RapuCmzFNINmOQTxdTCYoZyNPLmJjapkyhJ+xNvpF5ZVRwHhySb252lQ9ihzgNbf0AE53E7SE+fp
f7M6uGRh+uXcQccvf9Zf+5K56q0rbZnkXaoGZGuUhpCVwMWRC0GTaJ2HGBbWc3ubxTqZ9oFayiBl
l0UmcbnEnx5p3sVLYLbtzdwUVMfR7FZulPisLy1CTWoTN1HCj8QjJP+XOXz2aBJV6FEUY/+dBob5
+zZbdFeQRa4Me/vzKA2V5z3EWig5ua63VmbZIuNcDEbR1Mb2urD1tp+dJdxPHhPY94xgzjupYPyU
7HO00pPTG6Fhs5+zW5TCcNXW9J936jcZbSH1hHHQjUgTP8mbbGRRePT9sPocnAKoifb0/Xbt52RR
u+qFrrhsoIf91m3qnFsRy4P3XMt1TcJ6B0RysnF5etN5L27ClH53Rd3xFUz2Zo0mZdbM431qDZes
65umRJ1QcdHDlN5LbIDRdyvfZmekSr3sJf2zRMnShB0pwpIfI5CHbl01K2OOanN9RqBymrhUhoQt
++JyoEazSuLwU+huA2e8tcm9gAf96KlK8V9vlzUoshnxtjMFODsPnKo6ZBB/gBcWO4DU2TiF2KbH
kKKvjBrh+FMblNPOsyLcary15X2H8cE47uI8LyQ05gh7bNklEbSf3fsjuJO82/8KRWDT89W1tKyK
YZWMnBZsyVvn5Sje75UdhAWAIp4WjXQMIQ7+pkY27RcHREunUJpDbhh9cKDy69vvkAP00mdD0uXm
awP/Q/LOxFgznEEi3Y4jyQSaguioOCLewl6mUVH3sxqizZ+tkiA57yOoE8KJ8YR5RvV2iNvN1Lwf
DPA0Pm7UNCS9kiN2Cr9yldFOdNx8fID/zF7mJrgaiHW+WAbZaY8ze9bdSaiiuiVXzywBbjIcrwYt
5J7ZTRBXzjtpBmKyOYsCw911u3o4fsP6DuvHsmIjVJsGJThE/SCjaGjsf95b5Bxa+sshMR/z9K0J
bmpllvTCBYlYhT6V8SmVHqqwevRm2QCSBIMhcTyVv6v7HQyoflKMW9sRCJWqBip8snm3651++DH4
n+2Nsp4YCFNX72hXEd+O2u5Aj3LRSgYfN7n5k9SpyO2bxgeld/eHNPzyqA6jpEgJWxPNM206CJW9
b7Yx4tyBekUH1VtFENr4+8fEprsiaBwOI5ZH8VPq9qrdOY3sfEpxBi6TWGkWKL0U5JHSouxnwPJG
XBo0W3BlxZJWYB54AVzCCbzl/xYISHYk7HLQbCXQzUN96yygPjfz/Ba0PE+wmqLbsQCnYy6kKUBa
zOdVZECKI9DDQ697jQgBWUkq+oqJtb5g15BpcNTUAhNQH3Ip5TFxi4u4opag/kiEbSa3o7eNUXgF
j3OBTee3WPb3NloRZDWjKb9g/UeLSSMHej1/Ai+8ZW4GezswSs4BXEymb/XXRtLCLVyC7BJuka30
E4l3UG2fdXQk+jsyYOtmmvZ9BDaFHtDppcHUAImuMXyqkIwsO/e1ebBnjl0WZFzvfmhmJP7QfT6K
4OhQz3RgxuFu95Ins2eWlmpi+lH5kTBNH36uAQDhDs/gyWlqG4q61GKKK5CL3MqTMNvGkSTIpFlh
HyVBRzFLGu+zlcclYnTw7jmHDx7DMazqmSTUI6wzco9fEScsbGVEymEhF7rde5cHxhXssBXtV4X5
0IeSwMgi+XkHCPY6gksHiBq7Kzbysv4r3GkkwUzft4qq7x9MjCbwaJXCM+sTV+i1MTyq2oXGq04r
ZUlppoM2tsD8ScD0GUVAzK3bN0R7RYojVBR8D3UJC4WqbejppvobKiZDVf7p/o/N1LAYU6MpcNLb
4A/Kez7stjEKdLYE5VasIKxKm3Igh9G7evqauoOMsB+9V4Uv5u3bIUlqkaB0SipC1XW+kJKjY7m/
VkP0MZrbylYyN1PMp2lvJW6jDwgp3+rOZw1F7RNxv2n25S1tEPkUyhC+JgnRMIw4Nz0BtZuPTO3O
5N4KbjBupC3g4NYXhTfFkm2zLeGCQx/+TTkFCjnhwdO60Jw5RuRRMI18QbyIry4hz6PxqalSUlf2
Z9PAE1JWPoS8lkZgCU/ixdnuwKWga5wk9CgLo8aR565XD+mr9GgBtwnM9hGjVNKkYAWv9TXAa9Tc
E0ZFfqpa5CjdJd1xUGkubxnuiskZ5YC2o8uwO7MxE2dJWacBQiyfheFx0DhPsr3VoE56l8vhslJB
qkjlPNUjSSw1I96iwId0SE7YJBOxfz2APY95921bnKaH1MYBG1p+hxG2qPmaBbfxvbJcF29HjaPl
WItokSqEhW1szAQ2iEYohqO26PZ6Ql8X7ih3F90Om9V8Xsr2n3WT8Ll15h0WPnfR8/rK1ZjQMRuJ
FBKq9lPEcwB189w/6L7yFR8GF+BslTFKZYQZrt4DKZO+ZWyRcd5EiOLiz0rT/w4yxhGkAOb6wuU6
7JxDssZkckc/43Xa2GYauXI8aGQQAoi5DYGGagrgdWx7VBAiwmWo+63m/j5I7Fu+h0p1lWTlgS+U
n+j7vYJTSdhwhFturKrJMk4Xuvs9us+aexpjx8dIz5aPqWBBOtii5IQmYspQ/7pGIUVwi7j+HFWa
fO9iVI9g/WvwoS3VtAR5r4EUWpux5qT2pCnacktaRSf5S7Y+I1HDQbssM//ludrMHBJso3dDbxkw
5EV/rrXyvlid+nnnqqGBGzMX3JBT+cWt1m9jxDY6PcA97qZhDxiOyG3sB54/Z7D/atZRuJxvkTy/
QhqzM28x3phugqSR3q//aZuMETJqvRzCpFzm8KQXQgAMwESmdvxFUoFmaZM0FjiGiH1dyurtf7IQ
rvTvpHMIi/KEF2onhxU4cXvcEmH7KOyjm3jyACjSBGBkvyMePBGrpTxeiEUxb10+7iiqUWFVLIxj
sA3Hay0rkdYGHh5VOnsxLuPofwlf+sROntN92TeZpdiUqJMn/embyzOJNanRNRZJ4vbtXs4a7erV
o8GmUqZe9sDrUm3Rit023Bn0YhZWMU16cz9qgEgjkIAio5/C2rbrQ5mB5FFPPt6sE40GiUJ1zoKZ
HRqXYW88ofhzM2u8T1dpHPbM4beSLy2GpyHp2GphuGYCWOck20l7SP7TRjbIg4L0BwM+Qi2zYser
EIWQ8UppKyO3SNVaMcZMmFIH/zJ454Qyh/E/vthuNm+A1ZCjzLa48uplEWhyNs21d9xH6AcJgBP+
dJ8TVhLOiYQzIAiaHRq2FCGs6phyzvp/g9cbwObRNuPmmos6ne+kSi7NxGEy54D7kq1kFuYkUZCL
X6Tr9lEB929UttjiguNEHYd3oLq4fko/fY5Eme6NMsTEVvAvSsV17DaPKf4+bD/ykhTQNhzZ7MJB
8Mvs2qTxYwoigr/57PGTJKYhECXVjiV7vBYIrkKnmsTGCFvebvv28mQ0LFR1BfXlCCuEI1QdB/kr
cU1d4QR116w+W6VEuFjuQf2pTYZ9SZrZhvIcIsQcdOP5cYysjFhFsag8i1+mNyG/iNlmCgmjb6XD
J43jTFAwLXrPQ7my+JIYmLz7AW5hebdBXuvCu5TGMCcH4f5W037FAQxweNf4QTgaA6eXV9gO38z5
tUpbhh5uk7p2Dc/d0dipJi6NeCB+JdUzCBS0jkkKLVydbMk2bejoNctra0O/1I6duk+nMJ1QZBKy
qCvw5yp6tW380Yqw9M15MppiTlhqo82fLrVB9Cz0pa1NWm1B3caDTstJKZmIL0jQqbV6Pl00h61N
riUzaUW6/msQgeNKBgczIDTp/f4P+P5hiw3JhQQ3sxYGrOY6jfUa/5Wj9iJUkNZE3WaT/evfyZxz
v/vLLvbT6RuBwkt7XEtHOclY1zNdWvRKyPoAKdvVP8IjJ9JVGpq128L0+4R0b84hVZQxFpoNiUwa
/5XAMfqu/Ou5+VQmO2/r/y9jlyT/4+gN7XCtjizT+MiEmA6ZIxbMIyP/9a0dPs50Wa+hFxOhZkHl
daCJhQZru8XQa1vJWRGYK/t0T7y+CW6FTrJSQMQ7fc9V9Bx/6DsdfppjgmamvwVbD80izoRHIht4
LDOxm3pZEy1/GwoaxGL9HGdrF+hXQWAAzEKg0jfpkbHmK4isot7Y9ObKJY7MLEtBl1N86ws6oMQm
nLZuP7LMD2TzCsy4bhEcWaPPCsRsHTNa6Ij6wNT5H5pRJ6+q04hI3Ot7cgzy1mjGp1Oo/d7AY7Z3
PeycsUUIIPEjQ/5W4LxqRletW5adRjdvXPKGkRFoVpzZVzfc/VQk3wXuCbSXB/sHGMmHSydjK7lR
ry2H+oyyq34uWv/XhZNeg09xSxOuXk9AgTcrgU+1blY7SVPwidSlmvhJQ/9wxW1NyJVxxNzvG341
/jDVQo8SxG6cg3zHOPArbyXZQIeR1HSBsf01T0D/qUREXEbGjuHFIauf1xKIhWzU4dT/2BP6Ft0u
/qAYUr29F4nOIRS/XhbTp3wYcr/SReB1+S687//0nKl3BPC4Qub+RM8S2VxVyOBpsi2y9pi6aeCi
l6+JBX/cl+g/UJtnjPvHNDQw9RB5WTNYlOBXB6GXdhkeKqraCE7uDZOhTdSJsZHExVW/qiYIQ11L
iMC667qwhHPCcE3flygBs1gPhQwPiXcFfg8kmns25aEBqXW2x9o1477AIMJScTPb/EIu7fTCmC+T
cOpZYQpqr1vm3Mp4SiLWaVfZgZGrs1k3VTGolrsSHrRfJSCKFYKikkTdASQZSPicMWehcaMj//Tc
aQ8IkiEdGnIthV1huqHd115Obhg+1JKNTiTbvxSpKIQrvaRsDmhVCFdBCov7puEggn+VQiuAGIxB
/4YXCbVyljeF2Q4NYDwmtRtKppFJ9baKFfRB5Sc3DQ5yFaY7k/UNr9gHHe/b1RrTHmI8C3Yf1yq4
rHeECQ2YLWD/J+ezIXNBjobbU7AQmmgeze/RZGti92mO3bZ0KAZJWHqxYAdRBdS8vO23QkXxd6em
ogll0T2+LF2c7uX8xwrGUgX7l8yVkkt3g7tZdIWfvzrKd0a7B3sprgKI4ZbvfpxQqZkonFZEqCfd
X7ejEeP4c9RYKktJIQuTqUlfr/gvYZ28juq3cyP9GxgrLoYYEAW235e8Awo1cjDM889EuIGg9w1u
K9tcBPw43uJVvX0toJTTxu3auXCiLdqVvDuHyf1Rq1eEQeBAN6A7o37PMCkMP/495zI8wQ1/Dwha
WyVCOLIzIwS5Sc7jXjbtbQYBLjDo7gXIDkrmYn8atcWSO6asj2NqHxN0xC+0DSn6wJ5EuVSe94zL
1i01Q15HlUFkqw4BvxtrR14yRep3N7XxeX50BsRmC5PxvtpHN++H4xdiEZluvNf8AHt3LYj/UCTo
vdyEzqyIcsSmzWBUhVnvjzHudWwzYHj5vrxhLLvbbRxtFQVrPpCveGvpuK1TAwaJAN1yJNCNOQYY
jtVdNDKAPGKqZIqyPwmGiiQIEN6AkPhEBuDuftC8pR/+pw1vuLZGIf/veoBF9xJCX5GHrCgKRltV
EAhB9eqyclc/DaZt2XpwgNCV1NIN17lFKvJBxNAaJ2PA1KaN8cJKWvgNcp00mS+ReyqUKQDLG3Wy
dC96FdOQjZEWIU065RNmc7cPyBcRUgFpaqUT1MEX1Qerq/23wOvwME5qMwR1d1S1lysjT1CQHswE
aJ+zKcMW79drMvZnuCTLmWjREiziHcCdXRoHkIfi3QesKyj6un7zV9CUPUJ5R9dbFrAKXVDBXzc8
9nIFvfODXDI5rSuyNjDCj6DHabHClnpxkGhp+Uiij2flqqIIFBx+aU8BWE9cS+8da9TmvL5PuWTL
xdylmvOsuJ/Z1Mb+boc20erVKeSlJDOZUGhMtIo/VB+dL/dRxx+45rb+3t/B7HR8c4g8NRZwb72d
1Mn2jMffuDv891OeHuERFVSjG9A2t/lc4bfjql9ghh4AoL05cucAVzoaAaYFra4o/v8jceiSTXMH
jAvMF+S3PJKGYcNC3DRflKhS4SNqM6aaCt4AA6GorsUfqcB8I4z+zlxawEf3+6MfHM7ao+V8GcVq
jRFJTuo8wa0rYuUbydoJqxJTvqBg3EykXx57UH4XB3NVoZrLfpZ5T8IEFTvqIcpmyVJYQTNVvxvu
Jjw+IjdKKNmHKFtvStSZA+UfivRfXXtO3HppE2jzYJK/dPRyrrlUhk08i7x47jpYxBWT9c5s9y4E
4NuzQGaUZ5Ro/tv6Dy2+ykrQgklmkVVaywvC4QrBCEfLM/XuhB5LnvstJkvOcjuclkS2sC2HqEpQ
+FplR/neFly35G8RuLEBaK3qHVDP1XxL5YLvVndvdtB0VC9lvRssz7MqOmavlzdBNCgJcXTD0Ooy
WjZb9NP7MDUI2B4+6Fw17bl/plLU6W3U/BLnnV/xAy4oBh4wwebHCfbO3oGVtHDR6GNvn4+zhcuh
J74tvzcHzenMvsXLL1SF3ovfdGguCXCRAkkmrvay3ZEYh7pF2c2lW7ny04duC0dBrSujc1yuQla9
i0tos4KT1WYKF6nl+r5uO1FR0ECAiocXceqhS5CYsSTeOpz8Ldq/qGlGVhEfiy0pElAQngqTPBus
WWgwzjy6NsR8hPciInWXiqNSCPXdpZW4zeNLvDVG42wg2FeHZZD2qYKzsxHWwnjgtlnyGbjbI+RH
l0FRe7g11CK3ioaK7VrIyKr62Fn9VPbYyjhe9P7Qfyh+IJ63kjKKZL/kGZH3ombEYS385VYf6p25
ru7LI6oFhQBc97SK6dc79Q899kk+C7C+ntFm0W2PgutI6jU7UaLGGJ1bPhdBkcSJyBL8+l+RVzKb
SCH4MmTj37lj8Lt4+X0w8o0AaNR4VsPxg71oHJIEO9JLIhtBVpz4NZomvJCZGoT+65dR/t+xM7zn
dLrqw7bttXBeD4F2YcW2vGTyCPy8cY/EpleMQyJw/YkwgTaMFFx5EkBN18hVOO7k6wdd4NJf1uZM
pNbw0RJ20juGTdHUNa2c6kc7bpMHn29sSomEYcJVjw59YMLsw170Cxxqw1kKuIbQUb1PR0ZiKiGq
V4LTauS5HScQZrDKhKt9x0snuzDCyKPZnMBVu/szgBABq4UffUEVL6s/LQIAbs8WJQGZDI2GaAju
ONVmmFrbd2AE/9uvm7hrvfE0B/dHWAQn2o7v5WirPqxHQVZnkf2pLjo2vQdavszwkYzTk/qeii+U
KWLjpCpyKa2y+GTIBETbKRLy2E8XR4JJz7gODRzNdZjDC7J1/JyVAv1EN8e0mT9JNBYU6ckh5555
jJ1uFjNZnUm7KvSRmvLEXAHEFXNPio7lNUKVhmWCMm2T5AC493A8B+v0Tn6zjNsNzXTVi4ENMsUi
1ZEW+pFcyFHRKu4uXuSjirgaSgMSb83TlVCxFWtltY/Tsac1hOmzOUD630+oZ5furSaG3pyrB7yp
zcmmNET4g74fg6W5Cw5I5AbJe/Hz9qacQlkVtfJ31hRw42tk+rD1BVM8Sxq5aqXFoq9zqcxkeY9V
KqeUYtlI24IoSg684dWoas2/TXX3ER7VlSRIlUVhFwZ/rlgNwNa8m+PWxXZFBLip5PMXq9ngONAe
+esSCYJ2gajjFmTqxWzMLhQgQtxIidNWf3HTYwnGHUKpsTaxxjmGQJCXnFIgGW/5l+Su0IexYq6/
OVzDLTsONfcxcvFcM7ppWYpKaFIB8bZkiSvAqR7+YOAqwZnd5NcSkWtCwf9xv2pnzMAGFV3mhwzE
508hJ7HKIamI0U/tFe/1m/O2XW283otsOkmNAfL+EIul6EWDC0c/vcKqX/bnR0+uluNmkCTBlEAg
Nas5EwO0CwqB+wHW+j3ja/SkCkw4xXwqnIknKT893xEx76AwgVCdxl0d2B847/M7AFAXiaFw5w16
aHT7vyv5PjIPvY1y1WYp7DsVpD8RQAjO18vSjGfJVB/P3xePbaG4CVswZldiYZV4OsjSNnPR0C8E
iwTykVb1jotWHtIYWcoHexSt0l3aAaK3jP98EEmvswyLdASTNs3QubeXRfgagyGS9/OVPMmn0tfr
oEV+EbXy8GQAusV85WxQ+iM2vX+AEWQlxCcrqoojrPqxm2D3139HVHHtYLSxXvGWet4qg2H2aN6U
Iu3Sk3CpQkTsO0Imf0hjZM/8YFlB6LYF535WbZB2zXiVvrr4OoE6RCLy/Dci7tA94dl94yVJb0fd
HuIADSCjpxgdAA1bjA4GtDmRd86HtRejIMezrusJAciubvQ+Yov0R7fHmDq1Nvqa7wDt3oAYIh/p
JqRF9ab2rDzKO/wLqcLM2B5F6x6sY3Qe/Nz8fBSLQfPBlZevC49oyn8B00xKG4+P4DMgSHAHB0UK
3DDmUdfG1XKpAlrrzMUiTJ8+vjsSUuDRxtItTvTKzR9/cPd41CmYk0ISThWZFeBjhcgRggr0JpM3
sBeqdMd+nlYsQVOCewFNM+uH0oQayfe3+F/bgCx8BJ/JWomXAe7R9U/h9AuenozNr5fCOW9sY0Nb
WRQ7EsrdqbJMNzeFiqsPOco37sdh/zbhQD6t5xNyem3G7mUI7gwjPlRYhihxHl3+FDbZyKwZE1J7
SrtBqXm6TspRQUy1avwiYC6WXn2JypN14s/LJ34BdvsAk98GJ0mxquZfIQLhatvEB40VRqRcooBl
Cq+VNU/yQkr7brwadTW2I+twvw25UR7pZ0r6G6Mw6xo0wRCY7dRt3RwVL5fCzSgkCXTdgFzKvO36
kJCZxOssC5u8o6WvAQoMPC1aaEzRZm/H1YO+yhFda5PTfBKOw73XvSQdSMDt5zzen/iMTtPrsL1c
9TkmNX0LE+CS+eWho2oVFdXupb+tBWBNgNw5KhAtlvvnjyGDqtAYXSP632j3lBH6d0xE0jGIGKzG
K6dAGTujcX4kLYyCw8tC4acQzRf5McKaunnjCyn7ZU8q60xZB0RZ52Vg7xmzlunVypO5sHo2Q2dO
sVkF+bLNYMNXQTCtu5LUen25PE/9Oh0Ch5BILKLTwPZYpBE2mAqYYe/PsGVwd5/pdA1I/jtSKB1J
2uy6XE82XoZr6PiRhp3PCX5PtHY/WyLRhhc/EvmlHFbjcTWh0HrwosbcZ+jsQV2pBrrU0bNQpZKc
V8PYCYcDFToExqvBua5AFEa0NsDtAFayFeBFpcMg/SVoVRA44itb8EacnKCt3z7yX29YRRMeNocH
YbtW8FUiEAjeXCd+O+1w/22vnw1B6pcF0TuBzOF3sb8lVia4oURHx4hXUbyiVEZpoS2goqe34ixI
PRPfR0MWcjOTOtqQ4KR9fa93LUv7h0eiTx8rrfb8z51x3ysxfrSO0fWcC2C74d6Vi5suDpQv7XAp
wEtWR0Z/y4tpG90RANASmTUb1cocY5EaulUYynTZZ7eUojdSG6Wr++8MssuZ1HASJdDm6+eUxt4E
dcYws8RnTcRfE8ZlEMOMAbgSw8Z0wjMLkqr4RdTH53ZloxA+B5LQFbqVRwUevCi7CL0x1nFNyJh6
gyZptH/Q9NiCUFWrdAP7gtVASBIq7y14QIZL65elz6XNpFXvIjmor5CdxeoakpefjzjwTkz2Kb2R
eDHF7ciN7VDR3wrD2noCXtHteNTSqX+Mx8lDIkwTcXHJ51ebnsttxK+njdZqkbdJg5Xc1WFJC7sR
JB6BMVmEc3Hqh7CksrgfhVa4RPigQaaUkLQ8E0uZ/hjtYaQI8Y+TWUFSf9D5XSeXgVuh+TlBEDcq
08YkuFBnW5F2kzFmu1XWjOam3qUh5V6AnGVSc+kTpu9zZbMe/PZa9ltNU70uhturxEGryuZW9m/o
x7VXLFX8q2ffjuJQMnf9Xo2YJnFkmVWzC73UDq+Kl3a4D6GppU3CfIHQhHzs7nFkaiHuYu8ErtSp
E5rrEWQGGERz0Ncvc2PO1HYSbVFMbb63tcBkjv8mRWMvDbnJ6APJEFmCIq3QfpTO1AlW8InI+aJS
jWu02U51d1VVKx3u3yOiQQPTBNOg9BQ7jbafkVuvfBDAp6Vg4YMXk5nSOhv/B7KegReM0MdkKsyw
E47gCUNVoYICex8noK1Hh5qz/n53j/47zNJnqyBjkVYz77/vDnsVbKblRcpEETqIXTSSWkLDBPJN
+9QC7BGR3uHJNTDUwbimSZ/Vq4pvTpJGHRzQxZzBQaE5C4VYzLBG7AVejccE43I/SyMg2tBeHUNS
1WL+5foPrUCqbCi3yW7wdjPIt0LSHNye6NUOJVIQ6z4x7VsSMnzq7+XhVjDQ0B2XyRGGxJFd+D9H
oN6MvjkP1lAKVAFKXtimsegFnZ3bcOEe6+AB1OgFLLHI/CNbZXYANOo1hvZ3Cl8XkFYbYajvVUhe
C1EDln5hqu2hDZNeZKvMItKb31JIYpr6IDX0KweXISO5MhbVCldqrsRJUzTltuPBziPMSIUrfeiw
07oIjM/OxCdxG1lAgc8DFyMPscbnTy/RBB2hd+UWOdUz/chBZkgzkP5+7nVHkH2m7Z828U5pmlvd
nNHw4mm2YaTkKlfzJd2+hPSt1ZA3smJ9cfSATxMnMLp92cJaVHbcAkgaOeEXr2C2axs/8bIQ+IuJ
A607FA0h2+kwekU7Qp6swUUDquk6tzftxBGhQJlr6+LK2H78N2grOKP0rpm83kWudaa+JevcNNZH
jG3XNMfhS7oKUO94JAQcGfGqZ6hsSB0RBTltsqx4ILFZU3rvrhFoPDMBIqL3Hi94qDAGoucIKEPO
46gQDGl29fXU9VqNo/cmOc40LMkBTEds7+LzEjntOpnAWXN+wlBiyui/sY7DUyOEEPwuUJTqFDZ/
Ti365ZPEYgAUr3diLTaSASZmLcwWfJlmrhrYihdaaKd5ANOt879TTDBfAqL0Slj9mCJOO4aWKnXI
Kdj0PmbPztcuCIOYMDd+vc4/c78jmYuh73OhRvEVpFtRG48np04+L+y7/rTaSM7Nb8WndYL41NoK
LI/H/r2cmOajugh4LQMnxWehcVRQ1X/CkMnxjPo9nS1w3WEqWEZ6b8oWcx9B1aHigGUQk821hCBT
JjchEgfklxddlQk3R0ZOL4ypJbvUZhb4Cj0pufnvt8z+gxafx0LK6eCn5OtaxG6ic9vaaNDHW9yl
yVhHHOmNqgjMUFRwDaEw/2Pd2ZGNj5C80bo/TAWupk3DMO9ZVjPcKX8UF3F4qqZi+nw2w7Kb4vhQ
M9cg3GujLVYdzX65aI0dhRyWpGLvh+7+KEtADO2MbukRp23EcU0z4cvfIxeAuMNR9X4n7IwtSTwi
4gStHPWFod9ZUmqWK5sk3OEPx+ybiseuYrm/rYeyt0vyeupYjcDLVTmZNnt96rPFBhsBk4KWioA/
kFXgfx570Sa4s0tD6Nu+z2xJ6nrUv6/6NSsKhdDR9UAD5owrXNzQj33EyaTBh+RdcdYlKws1dAYj
aKK99ybydvQ04zyY7SjamtgycR2ikyOFhgUSpZ5QMfqfoKasDkjiojvQ6uvBDhY8shhASkLzRYm5
Rh1rvMWi3RxTfGjr+W3GW4w6hZznysVK5fIwEM73zD2Gm++2UWfbUvUURtzHkfPGxLetOp4HJyAs
evxJAw2b+9XV1Fo9WV0MUDPgz+Qd0moDrpiaYfZFXzLfIuU7NzYP1q7ZqGGMDcP7CL/jzC58l35M
IRfYr92ZM54J0+njVYcP2CwH/lXSyzk5Cwk3LAr9A4yeiYlS5QsdeVhg7bKKlU8S973NyZt5CagP
X2EgKC9cJnW+hxy2M+U87yg0Z3KnWnC/WRBKroq2Rm4Go7FYJKn9qzIA+CmosHHb4B7yhOQ4ugx2
xi6AFBTEqLmcTnBRUkfIKi6qRRy4paZN8r01IbZGPK2rwNoA0iDb0p+dUGNsKeKnLMsFNlH5XOkd
Y7VtQdLAuU7aEOyACX29LOkvt+Ya4ryLfc5gGTKU73Z4bH76dsmyeeDHfSER9TEUzexh8AJVe2tn
PVx8UGtYlW/1QkZ1Hzz0F5FGoDWRxcJdEWTzCgFAg0jU8Nj51N93UpRTJdLsRMjJDM/8umH9FumS
aQJUbHDiHXQeGYpFqRGQXx0bSoAkmllj87H8b5v6dz3HWfPVh9VHAIGfLgkIRIQh5KVdVXeFJk9e
ZkTsxdeDKgSxFgUy9+j1tXGHYoFZbYIOOvbYMiSK8X8Cj1PJ88iASMTQEwuUMcX8xkz+vTsKwGiC
gmfYHXtvxzPA1Ma7Q/5YM3rQORlHVmer/x1P6TZxIcj8B7ZavzWVb/M+XfmxyptqPkugs2zwS8s8
z7mHy+23xhNXv7p0OWVNrDsdeZL6bZFEPkdTbRBEnTG+6t4+cVZ7fV8sNI2uRIrasGuExpKqRHtt
dhg7W3mV7Hw2CVAX3iRJbJL+FfmgQhYnjerb7zrxKmRgL2o1SteQABzxDL7k3VgP+ypQGkYvRCGn
gmAPrNCwGSPa1poBRZJ4xpxWSkhOzyeJi0kWncpIjSITNU39IQzI/pjHbM2XECLiC0axFvD4IdTT
hYcB2aLzkJ8pQ7Zr6uN8kMGOnZ1/nZ+EOxLsZCydDVE78WvDE2gxBB/uIpph856FXX4HtRceRYxJ
mWfMrUboPgrceCnRJqbNW++9RPH/F2DHqpUmq7ijPG36BEhQ/cPaL+PNdmxKXmQwgNugY+n/NGvq
7gJblEYm0sSl1B/DHMdZUIwvDXnriC2/U4nvBK9N3hCurPQhBF49O3UmU6TNgeoTtt5D3m0qJUDJ
VNK5DOa79GA185XvazL7hKZ2Ux22NmPZQnqDmnbGpHOz97U7qlTI5UFBsvk6YSDlOfBfrCTaZfvv
tyhnpT+JFNr9cVgtOMyZnEKmlroTtvMNzUjy+/YppKbUd/UFKGDvXUHrrYLQVhMQldJgHmQvpAA+
TXn+ygY2E480qCLLNy0CNXe0c4VSL6x9ZeiTCTztsS94rpBT2WgM8BG7q+YxLGR6z8j5OU5i/8BO
Rk7+6EKy++b3V0Fm5RQ2UvPunBd8LRswsnO+rlE7UsXmmUc2UDEfdDzftBHp5/yy4RST5qsnIEbN
gczegpwikkqcGNrjore+zrhI44BXDp9OhJE62f0oBj0xg2OtzwFPUIafjuKQjRYVeQtlMOkjOPdK
8ktFRS8/bIWKdvvhMT6K5WPwko7DheD37hraraJiJ8hRIWDMOg/8uhgag04thJYHwlbTHhqfVYi7
Ugp8t9TWdkwUWzaLEbekNtFFIo+EpXGU6aS/8lKEMZR2/WAEx3NJ0r2gPPDToUO3qj9IV8VVzFkv
2qseAiesTW2gAU2XE+dPAsEcc2ZhV/kF6sCXA5O50cQBbroswVf/dbbD/jzsrA2gxgxWVJ/o6qDC
XrRg0UXu+lezP45QY9srT8rIXliy7bhVKd1NpqwcRjIca8McY/qiiMagd3OOZQXoiotjd6BzJtMk
YerVUBuIlpoNylgsTlbeFK+uGuHBe2Gwj124kHC/Ad4yZhPoFerBXCFsCpHxuCQf57B0Nf9/Oh3t
9kBuV/x98zoPkjuv1lp0qym+ak+4lijHMppi68kIXhY+6o0KkVL2Xv7NQMvKvF+Zui7kW9wQZoRR
VMlSgEcp8rnuD4ofk2ObbIVfhNOCwihyGAZeJPEjoScMmqUojWO2D5X2W01mHzKaln7Z7gdk79b0
/2IxxcSQwhJZm07rJkO0CTSTYwB2Xhb6Jta+xJBeg8HUCN80eZPUIp2cyaCGTSrIgiCJ2Rm6UE8v
ROL+g85b/x5MY44V4EZGawn4JZGAv4q6d8TvzfA94yMto/7V1uun0le89uM1mb+e/mnUNRLdoxt9
fU8EMdu9vo25A+c5ZPYVbD9nbzGkdS3SMc0cMA2gM6OuobArbw9sZBYaHLU6Z30rHTLo102wrbhX
jKw7ALCifny1Ir5RMp/7hVz8CZQT5ZpMBY/ItjjGNAiE2wySthOkZ0EscDLayGPPI2kZYsWb4GKG
LH2rUYM81ktKFurqm5SbumhP4ExsNORKyyGOWkpwfk7/fFHlnXxt/KQcOXHM+ePbXJEJRs+wa7gk
mQHPY5ZRWPEZJZOJGw3MM/fcQAwwflhcxuxYTiMtYnMt80/ypNAqq0v5upU5on2YV3QjDxX/z1P1
lA+P5y7jxf1tkGfWEe4+i98eUx6jpt1+BVhs9rDQGOCNcpzr/t5A5dUPfUVRyzpx7hRO548eU0iS
Ms5+q+rzUbs75I6L/mWHPDsc5uRT3G4TGJKddybjwfK6+WPbqJ3E57DaTJiWtHHK7bMAN6qh1R7A
Jq689f/9sYJ4SsAbCn/rkILxb9WmPr3ndDJimk8x+kk2qpMFpR1/ag3k+OjsKdssi9lP2sMZzjHU
Hp8TsRl1TIZAHtmZ7oTAb3P/5Va1mfl5jNiF7kUQ7Ogqgp3iEwkfdVTCViLCK8ICgAqZlJF0TFQE
IzbW4a8pF6rrStxt9vu+dA5aCKN/bjY/lvJhJ8nBU47UvVqkgvGYhkQX1E0SzUm2pZIww/9WBFIL
5gN1cbgjwi4fvzgl2muMFHCwjMvHl9ooGfQvYig8zbhpVWcqvvJuMjhFVy1X4dBFM6BJpEtc5X9u
oUp9AbFnric6xKaN09nfoixmbwJwOOM6qNSjgtn+w7aOsU2Mi03e+w1tVp93pUzPfy9RvhZRujzp
NFM4oofV+wFvuwV7i1Y3tLcirGsq5LpqQszWZu/AG5hx/17GNv2SFx6jkEt1I00AvVAzkPn36B1N
GraoxjjNPYBg+Sy51C3/HIGtyx0fx1hx0cLmuTjwt9epTnjlEXlmrClv2LCQFn32/LPKfSgWUkYi
cAJqFPDOC+YTKcIEtf+jwUPEAhSXJuFm1jk5yAu0FcUipzX5DPqVW4rVU3+v8R6Ht+oP4nT++ory
kzI0Kg0LA9uyAsUoduFr71xAtqIImGSFARIEuyVvqdXrjD7Wh5yaDJu81LWYt5S8wOHdfS92E9bz
ID9zhcE+oPSoAqNs082AEHO91fRIEka3bma3y4SNFXvKu//n+9u25OPLQAE8/MAJ0z2vbdBn3ugN
U4A5x8grW7Z3S/vTqHRG8ip6opX+iEqqz5NoaAZrP8aFHybC10IWxt95rNuczEFSmu/jLb++Pfko
uu3JYrkB5s3vvou53+uftVSns33Tr5TBz0NrAmnxJGYA2fk5Mj5u+2byeqH3Cm3VY5Lc1PNHJIqd
ZSKc+tktjLR7OIMkJydcpT3ExS58XGZdAhZqL9klDsnD2nToQ/F5KmZUiWqznY/O9HqKHnJiYxkd
n3XCy2XHMCA2Indiu1aqLSaRZi1P9jniHKreHLtZk4MLrocz89aLHNTDMT4DNZSYRhR/OmJn5o1C
mejolNeKmXZcLPjIdWYcR7AjxQwjDbWCsfhEh7x2VvFke2M3rQs/2K92gpGEeSVZJuDlXbpbx56J
rvf4bJdsROps0z4WkWyWvPkfSZgY8GbUJxZUl8hUgt7GMmrSVa6cfyhT0WA0pexfW2+6p4aLHGsl
vsBn84l4I7tHRODamUb/FLLOoc8yFyZiI3CTafaz+JLOBa3XPpeA4N2rXiBWjvZ2/5cQxF3J+o/b
WjAfxFatY9cx8Y5vXQE7H2B8cE1aimVp9w52NXQFD7KLq7Sml8tXtQfRT+SPVJKRG20VeVr2gChy
KP3oGFc0sIFNjzRngDKCwYrTM39Xpyj9jPQJyLfZEZeztZkok1YaHafLrE8RvEUKhoxdAg2f+T8/
J13J6mqMLwyVdCc81abtqlX6D3IwpP9XCJ4H3hpTO6h03x4TA2J+Kpy6PS/mvm5BkWNuTTbB1H7D
t0aO53n3cITJoUVfrIuStMyn2D6IQnMgBGkG6y88ooCmbJuBMkQ6twUr7j5iUEr/PoR473UA+f+0
8+u+C+XLEEpdvXULlw3XzRPnd5eniUjosQh4m4BkkIp7s8q5iYYnQkkTZErQsJ0cS7YL5TtELIk2
qePc3iXUDVIAAa/qXXYxkX127g0tCvBW6E9mglfoEbU5WWlXpn3ONlDXKxSuTDyCHes/wMGfiRe0
sqhrsR1o3qQSE2loGJz4icDxs6+BZvGx7FNGtBSkj2KeK/How9pCkvHzLXrWv6rSz2/1n8ifv6+T
p8sMj3L/hPJ5iW4kmChNszU0hjBG3MEBlGk6qrWgkcgbaBLQ4C+DRdJtHdl8pz+95JO1kk5Dfrh/
5rrDqKN0SmYBZ800XZRzo4MpLY/Ph6ymWs/rMzLkzZ0h05VkQZ+gvhODe/qcBgf2y+gvV2Cuy+y+
IL/L+NsqfR1vR241XcDQHAdxbgQidZOOuBKYlP2mMBXFVWGXAc5I9lzEvSpbMzRWLDLfw+/GeCI7
sYGWiYpiDf9wvQvGKl8xKJLg/Qv1aez6qy1vkXKhZyXNOTSaaoDjHtM48TyR96C3Lvg6Axegmx/C
sMeFh8pxtQLComSxiKsDt0k14HypMsjRgVgbIPwOkzaOfmo6dtxHza9+c91ojlWrfuIOp4mgr3fd
qrA95xREt1ffuxTv7nqf9euvHE4Df5zCGQz1DArkiwc/7JF4+2EBgxXK/60voUQk9AJqragH/W5/
UuOay4DFy1quld13CVHhQi9Cf6ZpxXQEj6n7X1HHdu8lInt0yh46e3TzH/ucdSlWDVs81aS3B5Qy
10aJi80+P4PkLtOLEYzIe9yECV1gL77qOavBmWls3yN7+2gcmqJ1lvydoFasPO6+YR82Pg33lWSU
bleA6ptBZV2bNsCjh+YrWKOPqb3MZIpBRdqimCqws/3k7jiShNDe0KRjebaZMvbLDzrQYjX/qLiL
cmCLg5OQe/WJhvvQSGpaHQOvJBDuZitNTqzwKF9Eg9Mz57B6tehRKKElPx/GFyQEl3xbvAZWrisl
XWsv+TuEh6DA0MNSvFs+pCKO2Aw3ZExIFvdYOe43XkQuh/E+xwG1FFGoXlLj47hy/elCeqEVy/dE
YuyJpIS2vSAdWZsfY20ZEHPOya5a0f/v8T6TtvbTO494WimejJaOLAOYOJ3IaMFGnPjWOZxYd3Ej
0sVf4ReaH0MZvf1az/NdG4gaYs1MxsNNUc2lCFDcny/ozXFop2rVQifztxv42xxja5ImCsaFa+T0
xO4/MLfCxgJKIGmYR/hjaZObKRe8p0x3JFLUlO6RgYjGmt0j2aeL52R9Kzk4DjAQ8THm8J/waqtZ
FH9aGFbLlzHbvRR5ueLCY3LYk1FIl2Jbqp9IpbDB1oC3driX9bk6xydGueetXcHsCND1jLSyE90b
iRkTaMH6va4pt8BNvfKnKEwIY4F8rs/BzF7KOx7snrOQI3qd0gHaTZeE61jeDSnMrxC6bW6leGrs
rjEUU1pDwQcVrejLAlZDuQonSrbUqk/xf+OK+2ibbEQUoeRzz5animmDdOU2SKBubWeuUY55vUUu
sPX/CYsvtRIWJxZi8borUtGV8QFGKB3S5JDSBPq24iZimiHOtkPFNzTyhhv5yUNGLgmvaDMASe6U
eT5W+p/qU9416X+7lr/U8fbR2gP49QjUOCbJhLvMSZWBDG6iEYUWYdKZn+InCex7BnoEn4dUrOaV
4EoLoAcFAd4DLgiaFZ/OvWYIzQUm3hMpAw9AgX+FVIxbT3zAE0HMzz9DouF/xCdDKU7Kr7Q9EK6u
p7uF+i75uYb8p8nvf5aUbKtFMgzCjB3ownhMq3TLwLmDtZm+ZC9xpsOFN2g85OFTn+IngVTNJd9j
zk8dkxzUpm/L+i9kVyS6KrhYDtBSK7Ak1cNSobaoxHrwIb7+g9M6fevROW2B2XRqHZalhmc53F3X
hYbtJwIE3Tjf3KK7/ABH13VkdCmdd/XoG2zwoEOjFB5yVBIA59YY4mFkGm4vxE2pkxPkN7SS5tox
wuQBHN3oPh5gcGPojRIwzUjNbT6igSQPIeNNmb++DaO3Y9iku8dQ2GALjAVYFyz7bB4LnNoJMaTz
Q4/8FB84YSSEM6+aHzAr/UeSr5kFPTuOKd1ecEZv4zbud1xF4nOlcNn3ncxo0YSlwzMs3fYd/IqH
GzZLq2L51GWeUL4k1hYKM5qrdoo+K3ZYwc94EoiiB750uuvTefI8eV2BvQOPONqvmt9VBlMbMlIA
Ak3zU+mCeawlCtHH8Dl2deDS3AH4LHZ2kGc+f31TpssLCewzg0dNpWMzB8z5kl7L8IoO5yeVqZMt
oh2OCJvd1MPxM0+v9n6WdL0NJ6wC8NAbS88uGLuvh6o1Jc1GflrDvZzaCUr3UIjN28RR3D9CBC+4
LwxEgH8WeuK01yiDJ4e8gULQwsozB8HhNMuNX5le9ZZ2Ha6AzFQZyL72Z9wtFzXA8qE4r3et1XdT
oektv/e0pzbTRUOLnDuUsydhirGCPSTx7uUKZw6x3L9C5NmmJJ1V9eHwmQF6rIm22vu7uGZYQHIx
lLZkwU85CzcTyFjZxWvYFMTw56lK0KT7/mS+9apeH+Xwoib2c7B92oVL/Jg9gyu3AhOF+ELbZZbq
YXQl5Bv0d0OXc0ELw/V1ASMocu343SlP1Ki+iAuZVnzeymcGYXv4IMjTSKLoqCTsFPEYjHwLYGIt
9HiyshaIoMBdEekBtAfOFaM4jJpyJLujshl0w+o+LlAyH27CtXQ/fIUNm3VjyZIF2qXoJAdd1JTz
7Nbw/YqJWGCY8PRMOgRo6m0i514B3oooIPLxZ6Gkf3lZDnOTTbmwHuVEvX2CIzmUOl+dtsJ/ANKx
zDmRqJ7qjinEOEq+kFP23G8NgKfZhYIvmQDJmgoLpzYLIksgYp80eB8lp4BcomQdY5FTDxz+aVI5
CNCHW31st9blrziob4XQxZGmE1JecoW0+AllhWW8yrPWvkZ/+rXFRRBTYndNZ/3hB+SOPwMKtIqU
58Jr0p7sVRzQMjXLSSqaPPA/EV/swcvjCyH5KP93T/paH9JV3gFHxZedBscnL31YhWRjWNK6MYVw
TE1gUB0dpbMWMln6AF6qE8Ke5n08TGl+M5lXhoH+bqS7TSbCfseMZTLL+22wjR/UXzMHkgaVi9p7
V2QNfuX74Q5QUoq0maX/LkgAyDh/RdqiJ3Jx+Cf6qy3YQCrgTyHyJ5g+7+9QjuqcQqfcY/NS3v1E
XEtKp3MTmGIh3jt9j6iPiTuAZraYk/rA78SZbPnqkoVxuiiX9zRofXoIXrfLWktp4eQ9eiH9mcjT
vvaVSeGk3F7O0SLRCp4ZgE1xrk0nH5NN10gTSWYaJACp7h/ktUmqp9E0CVl9ZsIN+w5AqvWSNnlz
GrZjVmspWREzBw94csyH4HQ/6PslikyyolZDPrhvzqlTtaIXPsHY7wm4RzGwACGXMEhnxlNLt06p
h7O7k8LhHaVmRZcWppKjVdJhbGivbm5P+qtpZeWpKfaMqRrldXTpDCiz+fSG0XjrfAs/E5KaKIK7
zuWqqDcw3aBbfZCxyV7Ioiekxc8kD4djzGqWXcwr3XObGOLUdPoJdJAWajJFnJZYCMww3PcxYYoT
cejv0ZqONeXPd3wm+Q77lySKDdApPApgYKGk5KOkduvzQMe9y/X0+oFNcRC6M5EK4LuyyxYiGeBB
cKRmRUq0N1hfqIuPh1C7Sb1adHhoRAD5fJIrfZd4oS6S/Rgq2yE0uqO1Qtppf9zsDRP+Da159NiP
klsX/x3lqbG3Gpof0TX344ZkOqjrnih71SN7Q9tY/0DbbeIbnvQ+zlfFrHjYoFNgmDCuSGvy8Dmt
k2V+TwqgxZEJRxGDjQHqFmhnsL22BLdnc/wT/EF4ywftG0GXoy35XZemlDjcttE7ADdIJLVEX6Hj
H+9smaPFRz8qkOuFBMwPCMXI/HO++zeCqwHn89DjRcP6hHU/IyFOUexGz1+xnv//QRqq5TiOwpt3
AUTUt+sBziVqGAFdxcKjwYoLep9RQ1CrXAlOgNQysrfka1kSGpUWKlCE94iUla8gUdQ9b2yj3IQD
xGKysSTA3eZb/V63mFWnmr1Y58jRZVSm0DJZegDu12RvOiZhZ3SJ2av1CXo1B4/6RBcvIAzKpAbO
saAEYVEYPFMcUkderAeEwEZ4ZFTf1N6tNh98+RtWs8qc//d1WMXxZFC0Gn4MRrsFvLmub8ywAIOz
r829mzNwZaKvMOpTEEn3mAxv4OUubjEaqFwSoJpHp0ODUHI4lUk2iGjQI8hUGVTepYa+0VnRhakh
y4/r66gpeqoPsVF7LAPT9mCVtSbjBeLW1fHtmKSyQxQd3wEI7ZN6wjISL6p6f1eVI+vEVQJWK2TY
eUL2PwhznZs9Mx0MEAecHF8GedbXsOv4HDjFZn9T9Jq+4CLdAYcLBR2BSp2kG47wtV0b+wuV37QS
qA2phwVb2YbFXaYnJ73RAdWRuuc0/vqObOrhz6s9tH0qETE6nmaJMGTtrbKWKveSc20f2ca2vvJG
3MXkV3aURZ/eFf9z5lJyePdpTzkDbwA3/0Jy7Ro+jUG9JjMs3UBfEx2AMLQBILPP4DTapwE0TBQO
IfMV1Sq1N3NEqoP0kJ3nBnXRBlsVeUQEDu1MuRZIKCIUJYijc2BTTJXTmWullOq28GX1ebDYH/Pc
WVNujiSs4CHFxV4F+SNJuAtIGhjdXH/ZwqpKqwcDSlQSYxkP99uDfcWZgHLmPGxMIVszTgySgbqO
VlGV57W8cQf7qlRG0bZxIILWczusCc9vVzjHHVWA3LVzqIzYMU54/9iswKR+077CpuBHu9qTDVFI
A4z0MH6KZ4VvphKI9cTnDMImSvo7Zf84LlhjPtOOXNpUiNX0NMAzUa1cMGLwDAHiKniTMlnhcZJ6
h+wPH8+nB6BfOmkxXgeTT8ZmR46Bpw++CZrgLgbND9GnmaGb7GgZDV+nKlWjT7EeDbkBUQuMni0m
T41zfLfdWz9e7EUh67GZTzA2HmDiHsyUTd2+ZTJkmWlX17clgFwfCgnJCU/OYt2SDRJy5j2NX6gI
TIn8s4auvxnguBJXdUyQQXkV9x3A2gw/UCSWiGDfpECYIrolQ+GZ31goovIuKrTFMp3babbAWqR6
YIfmQ+qsChNwORLvc14XLd5UqRoV3hBJZr69twpdcW2K6AXOZE1Uxy6yg5ZVHoitDHvtqHfiYpoC
us2I3MdMcLK19Fuk/14Q5kNxg/XAYu9zhL3GRaN9KQmo6XOs6eaxN3d+xhdzCG39KsYNnL9Ftayt
5sLy1UnYHDwoa6WY8ADmDc2X7DbjsSSHV8Yhe68+NqZegWsNooDyYOzGj00wrcOoUEbCHoogiTyN
nkdBWfqW/U6Dg+pTBmXZPEel//jc1lDH/xK3mDsOb9pAWkWL6NU/IR9Vf0QDXLpnRD+lAhmG+ABO
PdHBwgWco9v3ipXm0Tj0Pm1llfnTkpe1DZzoidLCSMEr415sMpclDm0zhPCUkjcEP/Ci9jVtXEO+
dl5QyEWekMewmTZGLJD712Onp7f6ONBXwhYvG9wH+RRltKbT7W41IXgd5oVi+cYTFCuVaoyw2ARG
/sap5Bi6bBEy6mCS8n97M0V/q2T6oMC3cXTUNoV0oCJZ99f2Np6U3dQ3hZbfKGrJkcfDMO3ZQ6L2
f+5T49T/EeefuOlclBQdEnqHR4N8v95HBP/RQkBLyC7fziP62H7qLHVmaUCMHSyMkZ4IgDu/O3ZZ
GFwCzprlxJdre6OtmVOgg5mmmYHPNvsRwvApijByUauVKfqkwh6j8PWLZ6suzvb890Wn13GJe5Yf
ZLLSCJ4CBLIEE7xJVlPE4dQq6tYfQDsp1iPgfl4W8Bv9QgRqfrgMkxLxWBuTpNIv564y89Rq87vq
QoVU+jxqvqwte6S2hqswQ7RvM6OkonaUIMl7q65iIGAuLNlJPs3uWy0RCh9SzEWdaGLK0Bg26ynY
KluwF6rAX1IACNWTdZHUe+yYq0DdoJaC9eu08xlq/wzkV5qOSpbsdVKr/nRkBRH6rpyQeGrp4qtK
2BYqZVpuaYJFbwFS6SlnRBJGUto/B++Qnj5WkqPO0YBVLDFoj2kp2KmdStX4yaTsWiDvmkCBwVvB
+pZqFzM68tM+V6ossYcIp9vaBJJWq0TqFRtFlmFuFCjrHqyPdLxTahbNc5LCj4sLaGykA6cJSA9P
N7vR9ObxSQGYzYmpHO3pgLPWptZGM9YE7kNnPCdoffzQw587CS/n9Q66jfjV8sVi9GZmYCJHutr1
BQJfGWLhn0fRH4snER8PafXnnwxaA1XUZmh+ucohNghaW2L7lIrE+NP/vVrBgjMd2V/GIeO9QtdZ
VYrqnhOjWy6Gb1jgdwOD89NKNQHoo/jIDHYhGJzqoXEuG9uNw7FEHzAuS/1vS+F/r0tKoM7E0Vgj
zbb2J0Pc3vY1xJ1vx4tWzg/UUJFVGV1/I3apMYTwlSAXIAnOkIAU1zyuQQ9oKqd2p7uMgR8cXfDy
P1mDm+ExUzhYQdLBa0RBS1Bp26qY2htOIAoant9t4oWotNF3qRHtixc3+XHqghiM9Y44Y9oM0+ev
uZ6Hl5jGv/QQTA24j0oSS+/Y0ceiJDvoIXBodBPN+BlU4RZYLK1IJNI6se34nSE4SUYw+qTUv7EA
RYfwu3O6qqcZLbJZpdC3/QmrHkiQQbB7YGiDaoxj13GFULUHH8f2HNq720Mp24ZyiGd1I0cmNPq8
slrSfiBndqepG34JbzHmN2/p+UJFrwHX/T0Aa1FpVtacHgLQJnUngFUPV0O+ymKial/VA/0fDP3N
dKuvL1qC5e65iA9tW2d/rNcIuGyyVykZOVASK/gCySezqkKVlrYGwg5/Do+9oyWgvzIGj8KmhL+B
j8GFiy+GHohQIFGyPwUSfbjg411P9BUpNhklVFiEWzqHlgLCUt5zwE3QUAWCqQaJEToiLRL+fVXe
7eHuNiUHuNhBXbMTVds8+zsT4QXXx19jNistAV1pu5xb5zBxhJ52aXYuFWByLgB58ylil385ECJW
YeElus/FDRo9MBGvHtR/XbONKj3d2w+bVPbv3TQ3rXBd6x6R5/PlO1m+zGb5MAaxg9v9UIHvQhuY
RFJVU2cWuS7lRCvlf5ncDDLL3dlT4a0hhPLPM7eA8nA+HxIGONjwNRZ6e+9wzg0f5IB1FaHwVH/G
kmwRRzqg7Y5b99IjDLaQIgqOj/2K7IYon+DpNTWW1CX7f3NQfHPwgSONpb40c0cTvu/GRUJiCwdh
GtIWl+cAx2fuVvhN9nrrFWy8v0TVPsE4U4KqNGrhLjtM9iXEHtBNXVTjdGGt9Ot9WVOGWpJObHHG
gkKHdf/u5mBs0TfkV/MYHOjZ8xaCeS07YC7tgDx5waXbFgWdsYn8+/sg3MHI4Ij5Z2Tqa18FoJhW
3SzK0Zg9Nb/TcbiMbV7fbCg8gcdDBYqf9S4EJGR0FaHpiHcbbRaQRCqvOgRestj6MYNr614OIZa7
kMLE4G80VuKL5V5a/TTVvEPuRtEi2oJEAaE6nqvfR1x5ZoIKMLUi2UOE2AZ+jyf8oX5cp/6yISUm
6uEtDMP+MXRqdNrwLyP6MJ6AmIMBHumt7bN616V54yH2/24uuNsi903MeeQHAD8jYHt2CrZ2BZGI
AtzILseBsDWJiVwEVy4/RsexndZHYeeqaUzVzZl1VNC0i/OwaVpCO7HeH8lV4mZpxhnDuVEqLINg
4SBtxGI8lp2i/4eJUwPBWX1X1BpX8Cs76O+iCaLKLPkZLVPGpjv+90t4F7KJfBRLsCcqAAdWIguI
I8ZCJEQv6J2ABidVXYiNTLdX69bEivbpu4Dbu5i/Zh8zssepJPfLTxdizrw/5DYVkVT0dsy7AN7V
fpv55P2MkRZamgv8GeRsxrXdlz8U72MWQR9UhrxlPnY6RebWeUaficrATeTn/S/RrtXfDi+LQf/4
tOqxUMDJN/P1ySZypYLSgFsbxHjhZnbAdIymxMt/uvNMSD+++xjKf1BB7PFgYyAtSonUWwq3kIZX
v7CGIwIOb9jsDeUg01zWPSIFdvhqzQVlKjpjXV8EFo3jyOhhr87MvIFgTBSGfzl456VO0KrBIGLF
RuhpixI3jn57k6bUPrqzc3A3Np15fBayR333qib6nvOeULh/PaUHDEyg5UAeewMrB3s440Eje0mq
MQ52zARj6pITZtDoHXrGpUAJGHo2AWouTSSU9yldKaLtp3N/CKds52zF0F+Z/ymzqBVNwAKb4rEf
V1oxHtQpgzJWYbw0DlGD7w8GY5X9uY5mivUYXTE9vCxQqcJ+MqbM2FnCGi5ubVTbX5fokjRMVLYA
DV/IZ3jit3Sdz0O0Pu0iA0RTW9D1bXvizS8BRbLSexzpvbdufQ9MslK2hlfB8B/DGSRdXk5xzj15
XAUYm0NBRdTSwBLyQpNG0m3oqZdLXArdZsFz+uZMZu2vYexvEDXj41ORPhWGQxjTpUvEOt/vw2T3
xAtiepzSO+o4bFozyWz8CTprDybRk2GOSnfVVXQFmhafL5Op7NSHFZKPXQC96N44lGfa44wKbREX
iaTea/fs7sBDkqPViNqi91QHXudj/Y4eJcxLLbQn/WRLv6vthxnDVyO1EflMTES6xCsFQYQXD1Xa
0N9jTgGs6iTwBG/ah6ZJA2la96myM5ellQqP7vh9/rWkd107xJoFNqfkl5w7g2fmyGgzX/HaSvFr
GxmlAxGpq9+LXRDwccRSkNMVcQwdzDasI4clqaNpEpiSQGk9mJ9YXc0MaE9jfzz6oFWFH8sIEMjE
4vDiYPC0Pvin0B+1WKtqMbGxg/mlmTfROm7KGbfC3RG1MiwvZFcNYc6ZjddlGvNJFZ9gtjhCVGjV
F55EF48yNCL8RwuyNhxqDgGQrbT66dwKnOIdNgEhhNU1xMVofyInT1rBAHq8oFnA+nI1xL4zKh+Z
oPZMB8LVIa1Y1VKzkbLM6fWvfvN86L7hGpOb6kROvKyhMnv7RQGEvq2P5DlR6h9fKZ0ZWtCIQAMY
cO1+0n5D3Q78WgVEetkbazGlKkYPY/18rkuYLvQSKLFht/8PW1sexlUUFsnsuiTUGZ64mkcdARQT
Nn4nX3QCZWAftJCOhAe/0MnJnDNwk08B4XgiaMPilQRmQp7p7QgIXC6adUYusm0UBhqe+dtTaHfE
yy9WmfH0yCyRG0n2g8H3aEpgc/9U832vRt/b3XVIVkujt2L32Q/LaNVAq1J18XFUCEHyUn0DuDe6
489VzSj7aVv4cB3JtWYOtCCT8ROWY7eZ5ttigw+GU1UxkcZEGwOI24rokNZsIb3M099C/bAix4kp
fHUiDBXGPSfFVhUOL4At3Wgy7TfU9P0kRot1rvYgDj+mydakMQFCO/4BOT2xQTd+89UX6Nhi6515
thhe6VQYr+9nrtNVu+KZ7UaYnYh1KQoYnKeHnx2iXNNoTLNTmn5nacaPnyMvYVuZtdq5EyjYo4dX
87ktXNkwOfNKQa/RB920FP+oj/Deu+wBoQBgf55h9zZLkB3QN/z/oUVX8JDbgQYQnCFhoz0RY6N7
dn/UZfi8j1/DDqHOqf/AmRBUM5CvH1sKX08n9LR2LUfHKAGPFxBFXKecAuRQhM/NPVaUXa90LL8G
eNcKZm6bHqyEPRhCfRZYUTjUdkIqHhUf5xXkNmD4J5rQgD6IzlYtfmFIhQcrRCKy8KFz8rCqVQGK
xuN9W2AlbkvR9Ebzghm/+T+93GhXDKahBLU2d0mbPB9aOuHMKTSQl5K0YsXEf8Z7mV/m1Sh1DK9j
bvtqM3uA4rffxWzSYxXUr0NBI00baG39NM56q6ckQBID0s8KUwhSGfvgNN9tNtpFyKCFwxYNKVYV
DcRREv5Bxx2TJXDhH9k/RpqP2aUHbMgILJ95BRnyYt8kqlPDfXN8IMpGppZa8OQPOk0+7YkrHvwT
NYEiDxuXgVZJnPjiYlncaZC0dTe9/tn5qVv489pSKyw+aafXUdHEEOkkiGSohtbuaV0VDR50Sb65
4fA1MMHXzkrFTrXnlaM5QgRjwoYNxC/PzO7h8bh7dhqwfwnwyzr3aIZwNFPZXaVRFGGfh4inrMgr
Yn3LE0BMlbIp3N38RgA5qZZIzgMAqzxTRrDjUlNTi9/RT8mFYjjyB0GvUBsBNVrvEVcPmoXbJBoA
VhncG3IKnPLvil63V+NdjMI3CRgfzRsDiTG/Ol0MBNoVqXlIEIBh3MiNGYsodT9ZqjliArTs+F0N
7t8uzbGKvPHGcJ8G09AYNzJtA1mCVhFbpETDE7e5Zvceh051ul0FFNBR0NPl8wfkK29Jnp4JpbvP
KYF595/HNFtPlxRevkOTKR6yGOMQpkKBxYGXAKkLIuM+QCWDxoPWFtncmnfko25UGRPGVtCnrmSR
8ChM0zj67UP3jPaa02K4rM4N93YjRyS4m/IPrEERuw/oEFA4BvPG4OqrdVGXD+2o7wxZOxRKnFge
XQkBQmlJp3QVfMr/0ATTwNptGXz0BM5Meazd04jTAd/B16fuKrTrMaYbKAATX0XJmnMKBDvXs+9o
Id0JZ19e0hilQW2nzCUTvq7W/cPhc1nRaPTTx6T86bhjWa9qayTyLLSbaofdEXZcLuwQ1GlPI9zK
4BwJyZvBnO2R2ZD1OF2JzAjMAk17RIfPwjVPT6LqVlbeQ5l1AxFScLpQM53Pjk0fZUId3YHpJUAK
1pcjGPrxQ/sfcalSkwtHyAdqW7pv8+x6LQ0FC7KT9WGEtN3EonO3LxdPJ3z6MN5ukRK8z/h3C8iw
WMjtanqwq+1qGOK7PR7/Nao2QjyKK6sjytVZJaeXp+EmEuodXCatbL96v9Bhzqr+4C0oLGZ2t6aY
pJynxQCzkqsJXe+bEyufBrNZrUlrUEClQT7QyIJKp0OwmsRPH7zobC4RhdSxzDIjIElbQl6Z6alA
hguFBE9PKczn5z9yzCyEnQS5ABIHmeXv9DWVbQcmS+sy3ef+wbBGHu+eYwFPPii77JVBnrhp7vG/
+kKRr5qYga4GJ2B3WlojyopF9QbfGByHgNDJQlHfeHGeW9+bIl6dDfuzSUTbtYHjGjWSQrMuQocg
3B8CGtz6Tq9LkzuBdvapWJVZqa5mHcBvcHs1O1ZyG4hTocvTVOoGP9bwvAgBRuIAYXj4S4CgvY+m
D0XrpDh5KA0l6MJt2Vq8Rp2PHLBd+0Ynm4UaIOs/DoUPm/OZ+iswVLn+pVjF3zdNQlPLQY0aS6tb
w4j138hzvrzgS2OF8S51riWXExd0NknEzGXrxG7yZP9vGHE+SxjBPEpE5D1gNivdKS0nTEzm9njM
M81YhlyaIfoAJXX19yX+1mqllqNMbs7/SWjMMXUcLdYEcznNAmoMHj/vzuJ+lRZGpzPaVLqad7bd
I8zSEVFfYZS58LO/mxO3b9hTAzuvMLc2ija6I0gIH0hvTAU+DAE8pHCraZz1h55w0ver4okm0TyH
quOZKo7eRgVFaWA9hVZQ6ScA5ByBAmxjPjosGAKMese6RCitjHcMHZIqMWSrWuJSX0/IhlfMAQuq
ho6rsTBgBJdbtaklxxILbKC68cIexhWrDGMsUempeUmnXuUZ96LO6VTdhUV4xHzc54vTAHVB28S3
4xQHKPtiuBRxigwu6dna8ebGhy65qVYnQI3W3KzNWtt2EpW8gl4H0oAQ+XudMMC/vCvLS30U3/kO
csE/8wzMN3exfDQRCUMkKopTzcn258+CthGJu62Uj+TVFFq9JD6BD+3nKQ9Nrdzca2Y/BrmqLVRI
KKYOi8XPOALjxT2nXaCvlVNLrSnfQZ4NMhEwycWnQ7EB3/KlQtEc1DEoWPp6Eqjhp+3JUBa4rJOC
N/K6ui8ATNAP846yzQwYBRSYxOfuYuGeDp7a0m3pf1o+wcc929sYLbkmgIZXmerFZA29LiquAKMc
f0QJf8ua9K9sQHn+pu+RY5z2pkEosdHTeCi84gmDDAQ/W0MyXnSDroty+qb2WZE3DzQg1oD62Hpp
buSBDGHnEhUZ+Jigqxh6i+nNwS5Bx/PeHsfkqAkOhxFgAy3tPJupLo11xdqxBwPTaB9bAbYZ8dOO
0vwKDAVxrOrZL3blJF4R1b1v3qK+lHL1JgfQxo6YB8fz/BYUifjDFof6PHeihQcbzl3labslv+SW
RKi/4jWLmSORIlPY0Y74PczELEvHvkuNY+6UyEc38B8mIHP8P1DipfsiUPWSEbBumIH8RdaAeFLN
zMV3DOk7YbmdkyBbAa4hKhwIEC5K6c87ANf2gInT04AInByuJWFxrsbJ1DkRWbVsyUqyhc9LsxDg
xc4B+JzpB+3N3Sb7lS9o6s8iQQy4Tw9aBxLzsmrqU1rztVVsBBZoZns0YdPEKbUfl4xJ+GMJuG24
bPeBg1QiJPrGTaU8flwXWZ7663bGoAqWOJItMCaYFZVTjKPNJn1W8yd++t9RGo+StzdH2oCgMBwZ
whtcUankdHYPGcDxgNohUHNGVYJr85y+p45/f3t10qV9eeYi5zMS219YqYVYLWz53KUvxqb6sx78
YIJop02wZmCqX1zGEdXx3KJJp0siC2Klm6X7klZkv7m63o/fiqeZij7Xdu9Cyyvt7+h62nkXlqH3
5iajxqYmbjGgRM85rdzBxwUjV/vYIfr+EZKrIoW13wL0yi2H2Ixy4wFjkRPtBLUxmvx2JLvtUDVY
8ZfEbFCoegXKNul9d02eolWlA/A6LcGbA294DZ+CEjiVIs1wkFmuGXQdALrW+lh1OW78/5PmZpju
/RLPHbXICGIleeslSBXSQ9aFMj8YTtjR3dsD0y9sMj3OJRnRjGXqKTK99hBf0O3Qepmb6M/ANUV5
brEvJWy0a8FFWIGqd8nFWCXbFPsPwFTCx6rriJvTntJkGrjq//PQupTKMC2/1H6wwWIXY+UBnXOX
vN+Q9Q0O79K/Wj70mMUWY3Qqpgt0IxRg6nbAIIRZTjh9+mB9Az+eIbzu2kbAKUgV9hgp5vnVbk9S
m7SqLLh/D1NfV6VByl4Uis0JrXt3SQVWcYGgbHwphSeblWg+wgEzJo8a9QTbnJ6t7iAneObt1ZgD
tmoZlAUWTUtH+FHZqR+Ji5y7ZmpZhVW7x82uV0lQkFQ6MaCDGyH8BwTai/fePilZBw64c2clOUEo
xwvqvrmuZbP62Py579zehnwSPX/+VFqUMzA4vd+rZDONXhOAUo/MSOXzfhCcAFYmkpgT6phyDP92
syTb9iGBgVdsQ3vnli5B1BApYlA6Fv4ZG+G5dtiqONJ8YyYI9xHnKqv0KbKBjO2qLi8GjdaFg0H8
iuL7DahsIvxD1MUF6Epho2uJDpFcV6fd2xM7KbhGMv/LVeZOJ4AMq3ncfmaEEadkizH5JRJqxcej
zd2J9TlEydXJ1mxeJIdlXNmKVoJWSYFNUf0WEuVMufU0uiex2uYULLuZl+GcMi4CHDIOfCD7nDMm
xHJ2sbH8DyJMXYlMdIk9dBOAFRtVfjIl7zDwPuR0A5m+LDB/RsQ03iQJPIMGBrpnXk2iq5vb3tN9
vZARS+3BcaXITDkwZEJsDv58P2KN+PNwID0PKZO6XtbBWaGlCvfwbLf4meh3E7o79wmpu6ros0xy
ZF+B7hLuVL9ZzbyrMoCY2BmmcOmb7mNmI2Zr2zbPREHUdU3+ek3OrOkM0gW9Dy5gElTTy6mj40vQ
vXSBi7tLsIKROtct8BFslMQzejg5+u4PTN9ofx86zdhgcbOVwc5yompr0pp2SLZvS3snQHI3NDfH
CATF7lF4PpR9VFlljMvJ6EUMpTCUNfovQb7VIXWRPhPY58c3qI/cwcxs9RIkWqKPJ52DjrgpTOKn
gXMZQqlw686PCmHhVnPjmN+3tnHyddfh1GqeLOgpB++KEy7Zjrtjz96bQEakyW27PlCdPCI2qdtK
O/D5/0EExgQ93CT3gFotZkCTTNoeMLYmo4dx8EQcJd068bz2Za+jX0YjVPdSwsqjfO0jyIYOpb+L
gFsTy9hfIzTVahQbChXCW4m/EgdBkgcfz4mzu0uY5bXZv7bVphR2Ry9XPhKzJcpbcr8am0obXlZ/
GA1EetpthwRLu11+N6Jt5XRwyA/c0OZIY68kR04f3LqTLeIlBc6zEbOTUiC6/W8RGmrNqj4+HWox
ohTKCoZs+IRRIxqJ3Lt0lMdgV82YtkL03TzrPKHJw3fnXkR52rYfSCi4l8CYF7QgFWmuy5TKAsQ2
hnR1gJC4CKkCtqrqtmE0Ys7v6lHanjF9p56fM4rW2zQig1tuLDL46upkAMR2L5ac0eYGTb99ppoH
IU1nx9s0fBHzoKbxsXh5qR8DN2HD4v3tLp+IQiO/uAJkjPywpHPR3I9EmmOCVYPvuAE91LqwW1eF
Xs4Jk3AIsmPmUND6K1aGIAs4nqJG9rMuBWGD3iVCGXVxbqJ1olcM7Jv1+3yvNbwp4pEXtqVH9Ucu
aCzP5PF5uiMW7JcfNe5NudunAiRUXzheuGrb5eUFbzbmKsNQiteC7WPEZE9QB39QEMmrrmnO40ro
MZGmH6X14e/ThWce76P3bC1OtVtUgpo+sOJA5t7VfOXZJD2tTb+/JzN8Q79OmprfegrYTfCPvnIV
LgFRZsS6STZa5gCkdHvB93gfjOZxJdAJ+2RjfPr0xbl+kLj8RCYwGzxxx1U5o1bFwkvH4foHyp6s
BBpvBal1IpmMRgn/WcoGhIXbJ3vI6iilkLycHgtW4b55/9uazxmj3vL20txaWyCKe9ee4/L4jrFd
IrPHoLUB9ZFw55/+W4NmLunsI/BNVY5slWRS276A6Z0RX177pvHq3YWCpA7VrBOXbSAsn2OXX7nU
q8Ry9kQOYxU0vw0xfXIVbx+399ofiOL44YvgHuug9RcMjifNgzz0ZyI7YOfsp1y+l8DgHsS9kCtk
w3ahLe6iojkR+XC4etD3GX0lzT5Gd/+bXXtAxKe/HH5iGtXgyTiOUMnXSwPwuHe1KIsPu4q4VgpO
l37tLJkSNKStmFuGKrBJ6T9bFkzipiJE4Cz7lJfy9MBkf56OlCNvxo3Us+fxcj/e5CT5moybkpu0
iWRDz4mZuyoTKbYR5Hag0/02RPFOYGTDZjP6qXVrJHo2lSCViFz/Wc546lxdlx8ba+Eo5AKlTgqu
P8+o2lmmXUeHKVSS+1oPs6TcubeXnVSFIt3jXkSICL1q42NEBvbgOW1xa16RQTwjsJ6xaVObwnTs
1nKVyk3TjC5UYniFlrbNf4dgaxfceZf52BHVVcqY0VAno0n4j/mL4kOFOXw0KYy4TRuJpPLpRXz4
WtMBROn0dYW5alVrNiTN+h0uRV2FYJ6TKUnrwdfz02XQ8CL8Hy+J0nS2QJqiYwgmO7odOI5DW5M8
bAQh/Du/W7lkDYeOeAbmXVxKmbp0E+g8X503teOa5u7/6UNKRoRIwMPTV3syF166hMjlxIFGNAAr
JQk2rh/s10cMW7x9ot3euuev3ZT7pZmKXx02Qn1PkfSWGBLdKdIuq+1vwE417+dCvzTPUp0tx/xT
SM6yvbM+DfXlx0Wb/Sg5TgfqE5NYmVH9IuQExDUgOrRGksoekaxjQLgwkgGRiwLOjFpm0GlMmqZQ
DD9a9+SUW9WVHsGy1zlI/gAe23bOs6r9O56fWFYBIyl9SOurs7HoS644AyD7O4DIQSLL6ulkE7RM
hw6qfmTV0wnMoMtH1kqeGibJqt65CeN6HAbUhbfY242o3semSP6/5yNDaRoUg657RrklDXZL8s+Z
oruGxcMXASQwYqAlsJkolz/pjCok5ZVW1EcRmKYYUN4rq2xwEUSjYnsT4nxRxRbWgxiDNEQ0yxmr
xExRaejejeGyeQqcL92c/MGFk1S0GZ6EIdWPdyED4YNxzzRTtTm0piQ04/v9cZvTZbwsbSJbEW7W
TlYqPEnZNRUkHBm5cc2EukUsm2OXai3taGcysNHsGHYwSxtRRtRGQZNmJ09LRVzfb4BO0rVncl2R
E6fp4z0hODqbnMvQOtKVllv4ZGTQelokKIN9ZnL8dkSgegBonxJN+gnL1Wrs4LDgms8Beule/Sa+
AKFLrvKYBn7t+GVQEWCQ6KZOwsJhh63tK+bX/ESAhIKU1eymSc9W+1s/l515CzoXtgGSxu7TUppX
jM68CSkRbEaToq6yCYXSZUD5VqobPmr3KwmupVAEUEzllzImC7KYVKxNak56ygV6r3tJXclV3onw
zPcxWCSRk9d1+/bXocfkV4YL9LfKbwJPfDSqpOypgVCinGGqfYfoE9xiYRDa5Nx/WsXgedcg6Icy
abqJg8pyAk100sQi/oe3ddbI1GoF6O5cR6nTn5YSh3jjz3szrh31vNMSoQIUeHsLNjyqDBsXTyy2
DyrCix0PEftog5z+UF/IRl/Buri+x0510VhPBFcD9PmfnumOehriHj0EHcYkn8t49z+32KV/3Fpb
GSrY7uMYk+rMKkLtIdHiwPo0cntLCLpa10SHB/rZNY7xnUC0R20XTansSRZ0VLmBurNck9AdNo0k
eCxySIxgvBCjRHbUcrWt1L7GU88FNy/Yj7fzltCEBRImUNcSI0vaN3JPoIXP5XLHI7Fn1dOL35Uh
tPqpWsVDIWl6roEXmZuMa1TSnKF3cCLF0mw+Ndk++JJ43EjnObfzglGlneLfu5D6D4KpfFTYYYC4
JSZy3cxgi3QNzZlkoEPgw46qb1d3kqRp/rMpjkRTZ75PTseKzPxpmoM2w47NuYKXxrr9QS5OORhS
FHPfnxI7VhNqYsLwMqTyiBSrJ3+Md04I7jyJb8X7XHu3cUNpvXJmD/JPqh4vUkYtchF8GVf2MNzA
5NUmoZjW6XgIiHH9ACAH9nsCq/zFSlYr6/3CtWhOXzmVe/aY9nJ+wh+m/kGaofIriiAHQ7C10NrD
c+bZnK/vssTDlVovRL5Zvq+B0GXl/9MbCI3IppsXtCufgcc4bSvQqY7vFHuKgqgw11nBVwf5P/Az
ULpEsbD/mOFrlpT80IxSqgrO7Fr9yLNX6USb9n/9lnlBbRxkGKLcjBRcCyhJjI4I25LAniODqVSN
o3yoeCU9ElUwPCh2ufVRGDIn8hDwj1fIDtvmnWAJN+4TefYWupzuDilK7AyzmSvgdNsoY9j+62bq
S5gUR66TiLg4ACLGSxAyYfIyR71kLKHqVmIKArEiOWClOpMYLsYqpQSsDWzN+B1vRqa60whj8QqH
xckC3wE8eq4aEtN4sK0nedebVuOISJQAGvSUX0Te2zxLmqB/hIAAyU0/FHA4TcPV+VCbnU/Gvpfd
lLmdyamEk0czZoMLVklNX9yF05zRC0cJbBrkIkka+Aorp4O/a7I0VL8xX9Def5ITQDoALUZWuU82
SQ4g1qMDepeqxdMqyvAnplkGOofhlzNJgRQUr7Lm3vYtLmNifNRk4UjYR1+5kW4FXSmmPFfupB1l
clANXg2ElBt6qR5QvGJFMvsLd7q5M0CqgR7sFx639Rz6q7T7xUtY23ucfgMrtuEJv5J2DYy9KuQq
gSkFbFDaBoJQo4riFY9PTK84pPIhlAgg+/daWLlFQo0fwNPdrnaTMyakSpde0MiQHCuc6xxTw/sK
9kuIMwCoCDcpshFf8AW7bdnDqqxhMzw48ZmYyPXzrYbbYB/WaITIZbhsd3EJaF5qA+vniqgmLysb
FbErE7rN58zM5U5J/cmoaSTtOYjYfdCiFjLMXYCTWYDYSfk26tZhe+FPzJhwMQoK98VD71ygEIhQ
EveqN9Vjwk9rFEVRqWayprlJOIP+tOPEWDtWvHujT93HRg6YSiswf2+UAZst1qvxviN8oPArpbIf
1gBLqsGXxxFlSUWMcq4X0DspuiLvXn2sHkDFuAEB2jNgE4Lk/ddJ0ZqZXzcwNzgVu6wLsvo7EUnv
ui7xEerJRQoHtQl9Z+JcHUTFRN9Xs1vAPxuu2/eHcKlMae/MOlyflGhKOHjkbYMTMX7oGffz8IZZ
bWcrzBQ8eG6pW7ez82ZXa3hOX9YAyYmme1Bu5OOmU12AFfpORo0OIe4wbI3eWV2N31OXPAU+tspw
kEFbFFSS5xzm77AjTt544vf/ZwWdn/erTjuOygIgD5T9SavwEiZteyCWOeCt9/exmtq8eu9y6djJ
EFpJiZwUMK+r3r1oKQrLre/NtAyOzxkmm3CouDl9F+UT8lwRjbHL4PlSYjqAJyYFy3yDobnLZEi7
acE40qPhKkRmTIZe0FhC6rzjGJhB/sGgDbORjx4NWVKb8PH728ABI8n4pvJGWuxo9kr7w0658wd9
cA5hQ9PGyAn8CnILKa+NIFoXgS4gsD2230eHrKUwQ7cwU24BR0SmdIz4C0COchFNYFDbu0CUgvPr
NRIHX5KUH5q6ahc0dg9way1rh+iyyQgnmYACm9UjAAUzgs+X48wBDgQM6gkg1SYC0DVCl65l58YA
o1fZdE7fpvICcdd9xqvbEeaBBpI5gofJ6nUdJUJzY1ZCzQH5RspNdNMqS7fg2uIQ1f170wq7Q9mg
rQ5Z7SCaC0ZEPiXPzUYv9NCj5UBCAl+abCmBBqCJEVPrOucGnan0v8UeBNB70UItKBi0HFoL12ZI
7Z3+YlP43P9UdEB01XGwfmThVo5me97poyCJsW8jeyx2QSTlLCTay5+GnsOS/ukqJvVfFu1WQIDt
bVJAYR+7zSRAaQhVvAGeXMhR01C44Wn+TjooQV5qJmOAFzyZKfQYTaZWt/L+4CPHHu1mlOlopECj
X4jfukyxovjvScryOFFBMh13ADGZ797I8EEQP3FjRi126opqqTTyCZe702Qa7zvDThsC2s/aHEKH
GxBdoh0pqfcIDpQzp6goGqc9oX388LdtY6YTb1qYnL4lRjG4dbZuGf9YQdhbkYCqYTxN7p+ZKe30
C7gHtFrbTUPsEWVjizENPVlgOCgvV/dIewT+mwRphhFeJN17BHZurZzCNwDBnt/avYszQYx2h25p
U52VaTSnbRXnvrFagm23EfFelKRr+AMnpzDhe5/UrGdffyfg561nezzpv2dmztnVMEd5m7kg7dcZ
5xI1f2oZE6+NQKr2YkmHnLqZI480vfclBxBpoGGaPHeq56rPAsGINNHof+tI37wTWg080kZFlzXC
0uCjk2WONJgMOMHCXTJXX4UYZ/npZy3QgvHRY5r0jydYiLENmDmEvgnaH2/ckloCap6Bz+0hZFb+
L+DlJvymeSejmNkfX902Chzgr5eRK4FgBtUJnIZFt90td1t8qEaeUR0QX5tYLvPIP/uSQ0XlKW03
czd7mqfne5+oP/jw0SxI4ENLblsUSIpU5D6db7viRzQPosDuKwPLyP+2TJ+J6hf7dMvgG4P9i5MM
SriDt+0eNEBcCZzq6MjVl92k+I1tjzar6z/1kSWGu3rIW/HX127wTlAkd6l63fhatwGbtbZlzsWX
elRTsZwg06wHTDSiwecP3tOyu7h54ki9EzzJ6e1oUgErMmg60ujiWghNUp1MwNQg6J37jGxcn6D9
41zz1tSysM6D/c3S6cNQNbNbCIUdKNlqaybwSVGCXnwg1BFGacl+tIEJL4D44Za6kqWbGo45BwsM
AIQnGA4lJGvniv0ziiOYhlf53uvWtmTHiWs1/zofZJLPJKWuknbauRYAh8pla8Fs+htfYJj3y1KW
YPQ5Q/b4MYI2J1fTePi3RrrKt648NLpoArKZdxb4CArR/0Qsgj4FCDUFS3n1fViTPPApsL1UyiIK
GHc6DTfM6joVzyH4AdOmf1QeBdoeIRGlW9wh1tKRuoEGVqeEEj1pSFoQjgHn6wMvKd0jFwoLmtKZ
3QmXgp1KEuGRa3+lsN5Axv3iHJoLPjH/W3vED3gWJ1cjorLyfLJOrq666G1W1CFXhmyd7y2hFxNs
LadvuMewI8yAbSbsTKBzR3XiSRfOQsyrIUwwrCAppmEvUadjN3lF/Bovs8BHWT+6s5zLlXRhaubY
LX4OLf3FVtneGqJT24mtuYVWyZ6Vr42Y0VKqDIGq0/4mUD1cEOnCoXj/J6s2f6/pNI3U2QTHhIre
77HmnpnZwxORztDlrbsShyPnlLmBAmEfVE0gv7dimcRrWABm4er4JpkwtwFzAG5RWTqmX0EMwsN6
s80wH244PFu6CCqI0xm2tXHeKbk4/OquGY4YkLjt47qszkFof2/kCfc6QiQVYe9gerM9fk0WIr5f
8/J1wViH7AjtMvDIkDzCVOueu8neFJtMDxiK1i/DQpVTraxsrzA9z+7kqHBHyYmEYJji6RfKpr+Z
90jC6AM2vsVG4pvTYP2X+M/wuSeSNnVN7zGtZy5J1MvdgGi3B1qih/GjB1wVD6Lp/5Vb5nHqIOtZ
SK1X6/vatxyKCHo3yUW5RSe0be8S0A2W4NTTja3uEtEKtWEuU5cJmlxL+p2faHWnJTsYDu2wNlBQ
rGwY6XOzE+9+scCiCD30ie+G1beED5iFLDUmHjZFyG0lm2BHuqTwFakm49VhfKQjTqrkRnMXjLBS
H/fG3xqXUBp2yTQA8VNQHOK8wYygsO60G8iyJ3sdtdUxvmv6p1a1mzBmd7g8MoWpe/0Sp1SVoJ4K
W+8kzK8wDuhjRxYpv8Bnve97u2kZlXK6XInJ8sgqtBGnQus/aL5PQsrKw88mstIq64SUhuTI/X/m
xwVuvk5Bn2SSoB+JAGFXQOIaPEOt1cDZvli3z0k0UN0oyoikMbADuAEsxu4zZ3W+OCCdC8YUMStN
Pls4flu6ls6OLJ4qccIUajKA2xyNxLp2AqxyfM9wZYAe9r+dT66Lv92WNodSaFAioDAeNZyyWtjr
hmqMJNq+x8GFkQ+43DGxgubIcR8jX0+ZrQoRFzUs5EsK/zHqBgls3RaAgjaSfFfJKGjZG+4uFgl3
FkW+0T3/vTafLQ+dGSIZJ9ONKktKidJUQmldV2Y5sVAzX37pGf0yVUU3ZQY3lWQbbaV2kOk1Q/YX
l/yZtPboSXrsAGjkpzhzQVp0pgV2QND+dRUK28cluytWp9ZRmQGiiaFai4s084FX8Cy8iS5/lTUj
oGXws6p7jJbamPirWNnR4YV0bXPOPtK+pb+pB2RVVo5+8qbi1jTHhxJn/2a/bs4LaKQTM39AZXm/
x3TZwyod72o40X9s19Cr8Oy6bN8MowVpOl4BNlNSx7bhlQLdKUJ9FDqdv+AVWvCpucGFKx60x0gX
v+HXCr0puXlgn5PYcXBKUXm53+bFx/MuBXP0nSi+F03cEn2igQ+w41EQrRJ13VJOy4Ss4ktVE9Yh
Tl7SDghM24TLKoOFr2+QPcprY8D8WJo4b1PYWEHgssULSkdOpr3p614R2Bc8rEvR1TgbeS805dGp
LNAoogskxdoXXdfoOayLo+kg2V0BgAoAmtj5p747zybedTK2pZxZ8p6TTR2P9ZA0ObxbnY3sXAoD
G8emAJi+/mm7o39/NITpw2T3kMSdNC73Ip9r2COsyOG1bFQrE8OYndwZNHPxe9qF3xvQ7AgmdW6f
FBPAnJsZpCUfOdOVG9QwHf8ZDIay5q8qL403Gp+VCFXeAyXaYEfW5Z74DvSjM8UGvXi/YpL32AxY
Ud3jYyp+4Pg8sx+G0jaC3sV2feLifD9P6AR4eKh0JhVIzbWADOO81GTYbUSJaVDA3Jezfr96ecZB
q4TrrWXsed7Ib1MJJGlc2/ft6JAWAj5gWYUZ0oKNcuUzS2xON2H0gp1+shuu5FnFqSuYwa79HqZO
r7kKt8JFMV5Slauo0DhwNtVfxTFbXi0BseZ4EYzBBIACrIhoEf6lJ1RN4O+Datkf9zkItS+9JLw5
ZP+3Q6faCgyHQnzMwK2gUqFThdtRrmPZfSJ3/Eilize8zjryfmYUgu3TqJXpnw6CUcITEoGk+yTs
OSrTpHhk6Oqz+Y8k5x8FEV9FUkdG8GYhLkG+FvKYS7Uof69C3zsQcvpWuXgftVprnxwNT+bbzeSW
iuILfesVev+P9i2bZC8gJd0KsrlXBRQnAktAbPWQhZkFC36q+hiw1Fy7hnBt8dD+jK3dHlsK657F
epM6xy6atGm+tAaxp2ElPXZl2jzpWWBj/drLVtOozOCj/KlX+X8unCgpgyaP3uD3qzuVlZqhFVFK
geclIDMmfdOjFxwwFbsVBA1XB9ileQbkMyAPHBEFllBE8ptzsFuthPco8XepAjoSfR+cOKqBIAWG
ylZPwhk4KQ0LbJZeUcgDTQwFUMj6V28V4rVtyBoDDOLKefaU+VabWth/ha8VzmwjdzXnCMWkO9R9
h9I6ClYjWwtgQSuIwAXgV9Uf80QyUHhqJQ4eRyoMydAS0gsFRHkn7sgha+eSZdN2OVcl0tzH0yyi
vH8gjZzMsJWTJ/KrsnubX8MGj3/YRfKsO90npq+h0dk4bz/0OVXqzSd1OhztMSTj95C3xqUlCWHQ
8pavQK0RlvoFbjwVOes0diOxNC6LOL0Q6YnKPZLb69RULjsCcqrazI+z+lLd6sZqQkE9kLeIfQFj
wwZJHKBvGJfJYgjl0hB6HvlRgjbiMW2MwZ1As+THcFgtQQVPFyHPfvTnto1RIeLwuE+FqTL3zda8
kC5PoRvbS6d65jn2WTwrQPpmsUOE8jcBEZIL2uJZEXIwOcwKAJWSDG0Bt/ZHciqhDlrwuL6opxJo
hmoQ5+ApLbLwhVePSWd0cj0k+niXLnRIHYCeryqRQkYVl75YTdaWF0GAJRiUbwCIaYQpe7wjp6By
lY1D3eaowxXtG0ghlu2ETKFw8b7KAjzjAdCdU1gTsYJa+5clt7gj8JixCb3qAG/NmPd2Xx4Cfelq
fxWN7sK4g/phuzD1LGARLYhx51N6uy9hqQ2eBFS9gbB1VlAD15DC20ctoMdNW9jvIRZIqV155Y/4
RFmwtgFsxnvVT9eek1D11ZXvq0jzVLowwfQFY+6LHn7CJPM+vsvIuyxCxxW13IEvRCcc4qmEl0Zq
e0kMZCnZCk/0xnE/uLSB1NDINmJyb+euYGUo03kinq5nMPHNvs/P5lNdzTTz6MA634JFxXDjoAps
1DIvC9qprjpknvcUZfxzsj9FkPnByq3nUJ1yH417lVAwwJHYYSX4Om989s+rpgDA2gXosf3BnW0D
WDnK5mydJwrhdBCQAs7RI7574NadNKl28fwWyaI2vkdWxh+y10CUpELYBv/wg1s1nwUNp9pHj9c5
mv3DYy47irBBfKHceTywf7ZMJdFzvzEnJ+m90JpDSkeKotxgUiPr1bpoXL+QKaToFIbQOqpd2Hwj
l9fdp7i/cufCDscS8cXtRYSXmcno5wtdSqfWPAUs9HfM1QERB7bEwEMX4sMsndlD551AYnFgdEBQ
ih1dYItD0LWAw6fnFm43ZnRHyIGHYECTJVFtNq5YzS3cty739mc/DnaZ48e0GW0H67/m0eQ0VPAH
nnKVnDRzDKfszgJ/20VVa4XE+2DsdNtlEQvM3kYy97iHbodYXMgjUhwL5VtAJO443L4w2WrBmjUq
M7pABLHoivVmQ66aFm6O6B9nOTEiXUNrSrd+HLnnQmbkaaDwNSKaBW4qr4vP/N/ZZboNrSkttjPX
J7RHmHhe+mJmBsAfJP+BIa2iijO9larDv+sfJl+GaKoFdEuhkgWWqX84XwQdQSFCldoxShujCcW5
hTZhpGOGkPR0pw5W53GWhwA95vpGLht59kYqU+m2bANUwAMdvn+Fm0VJjCRoLFPOKY53M/ex+/QY
+l00Lz6Fev61RIi7I0h29PqMFFSs8DZtikUtBL1TBRK+MxMnwJiUlPCWVzqVicnttw5Vga8/bV0C
0mEdE6ztec7wMXyUlh7caJQ2WWp8pGG2kncrNrfk7B2yEGw9POHRwVfRe38TZtAhBzU16g+A7FwR
g+InNErfKo0TWEVcyny13muffaXGj4b/uGonB3172e2850fViuUyVgH+ZdQun2NmdrxZwedY0G1b
BRjZlM2TiIKAlYuRnPSQ4Akpu1Amo/+bS5skzdXanN1dCVoklqCghRMvMoioIxjDymKG6BfmwFcO
JpuQ0rAPKa8Foz9NkIKW4pA1TVOxOaymaLaa5Uir6ErXa67XHa7nSCCxHS4gQsu5J+GG/353CtFv
5jaz7HgL4FEn3lgkitmO+GGOoYuG1ju+ftPUIizCmvT8lHi/t/ZFu+1PY87i/9xn963V+boGlCAd
iuJc6A0UldX8uzbh+CA8IeVEqWs/LVdFY6ZLIA/ujkGeM8jASkC/UF0ZbVNkwZ2Oz3sT2qckgprZ
fFR+rZxzCyyZigEHXDdiVdFmENBQ2D/KOJCCQedMuuLGTug/9wYlYLU5NiHuf9nriuW6aT/vixap
iUgs6FbZYxsyCHFE2ZvrmRpYEAhYmlpwgfD1/1DNQQJyQlDshWNCcHn28ZKRN5uHveF9szjI6jdF
80o/wIGw5fez5u39u9Si5MD3vGopp560tJpT3D+1Z9D5kduBaWR/9tdXOIXGtwj3c8sYYipTH9yx
FjUsfiLxImQB/2rQfbeHuhfh7Zz7cgkXBVss01Xjwtv5M9Xqjx1OvLc0RPkkxOt0Ljan85m9+XrD
W5xbUA7v/N2q1I/D1VnUg0tfxB/9tXL+O+ZaRWqq6K4t0JJgoU07TlFVM/wGdhYo19U8tnG7+xwm
g0ynZTYl2JqtrJgZjvuHa7aGsh4k9QWQO/IbV/zOpqUjLNk+TEuPsOX90+5OW+vSlWdypOZ/Xbpb
ucjRCliUQXytCJX/LNCHSCJt8t2tFTm+Y6gatRfxvRSvFBiAqsFAe0t8fqFLR2k4Hv/0iPIOFHcm
A9b7vTD8yIIjaAo9K28TYCEmJI+UT4PBEc0HIQbtb+sO18SsNDOtw1e1XTwfFVtTyp107rMCmVVL
wgzsTzXs++yRy8HhJ5jF9stba4shkOUCcOmyXjRCQ8/1dV8Ohwbj/PNELAqbBNS6y4Enw0VkKuu3
w/Q+93QvXEswJBUe779ohAfhYhCR4GNyYM62K+BmUCzhdrMiA2u9CrPfhO3Y7JUtOk3xd7HYpun0
ASdUkB/ukBtCwHNrs1Fb2BGpFeDnaeecvoGqTsm1m5vtwREf5xZQ0kTnZ+35Cx6hbN+0Aw7ZedS9
hencdKXbaQ1/HN6FGuv6jXqa1CudBn5Gnqw6h35F0Fui9BQhL7xTFA1ddTYBs3Lu9uBX2LjZU5FD
Sw2zS3Y/go/DSwilOan1WIVSK35y8Ts9dL8ZNdm2wlh2SXf8Br5fZslV6yRk5AD7EeYeu9ePyB9i
46BZja96H1wMPARKpAQ1NezmdcUZqiIo0D2KNHZp6sg0lYr1IQ2b6iO2XJdHciK1rUZkId5NZqnR
r8ayjvvtyNXkTQdTfz7R7azlxiHACdXCJ6gRQSFZF1YubwMBQPc2St3CW4Yg8cQQAVuWBHzarZGL
5quXOf+/DhqPHmBVm6QMYL1OGaCBf3/sLIblgJXAp0WkqdohNSnhzsRlottIKPMgDbiJ3lorwGkL
rt/wxetSFGkqNH5+dhOwVshfWXn38s6L7tUP/tUEl/ZL9z8c66EiMXFLvhjewYTHlhY/lxIPLq2k
jY3rFLwtpSH1p1mnL+bQAdaLNZ5+nHWmX/FFeyt1K/Pql02Y7ZQixqxh8n61c3fZXRjwQRtlqHrb
u/YoXDu2g8JizjmN1U/4pGwZxWGHVIIHRMySgYWM6POL9ZOIwuIddL39OsiW/x9FIDSx6tmDMqdw
C7+nJ6FPCVhul3B4XK9QQNJ+W83iXJfRFi7gUJDvmBY3MwkWTopV4MZcJbaC5oneddwyrl0e9kG8
n7U5nzOMoD0I0ozL4BTldRDtTHc0poM5S5jKUgg2DOLneqXrQ9IE4KKo14LgyuV41WsXNzjGjbmo
tLR9fcm0B/zdZFaX7/Di4CQ+W4nIml3Sj/ektlfewLFvxVWiK6jzAy/QAthn7MoTe00f8MWGospR
DZvRA+2pf7efsCoio3jD180KUodW5k/nerjZsfm7CyqTyPqZYg9agbCcT3o/YVAcO/FHXED3hq4O
xJXfFcTF5dkdjPT4x89xfvNg1tZCrHb886hEbeXAhdFBeHpxwcmi/Q4wNjuHCAfsAqV4xsagJa9o
hFcWHQuLbkyvNaL88emnGIM14oppaldGb7hqIR82IWK1QjDIkkiMN/8V4gqC1EOYCGw7Dj9b0E8C
tSPS/ZyNkHMbtjWQkTn14r1PMIaheWETRmbb7RPY8a2kK0+UOPqu5t84lPQEqK/8lPwKmlaZiSEt
FhJzVkHzC0oh90FPr/7FI8bdm9VQHJx4fusuKdla5SdVmBB5hf9Usx4tFseOMmN+jW8NKg0yIjBR
Q0tqKVDrA4Ekyy0eHLxFo45KRx1ZeOz7ceeDt1qVwvZ8eybJPV8A8jLX/62T1GDf134ZI3a6i3l9
xXpacuozL8UzM4dX+2O6UdvrObTlcIDa2NWlCuOQ8hcpHcWHsPhPbqO66cd7FkFoAVK10UzsMQs8
jn9uvt0srecatPxmhUSJjHIv11UEcItIhBi7M0O5csAg86dEqZAuRylixwgZmt0HC43jg4y+nUoi
02gXmugILepoaE5qpP9kXZV4LwL8EEROotomsWb8IiajzKYJFkkn3JRqRgdk5QhEm+xXPl8EL8v7
ib3rU+rnrz539GKcwdkU8fDaR2UcYZR6AhIQJT+Dp9o5prirLMCoaaF7nlVqmBZfw0dCXEY9xFvL
xlW3Vd12El6pNPN08idO6VTLM/sd5shwAt35mY6V/+ywLdTyFN2y3Ky7zbhXBHu4LQfKpqQxGJqI
lytjiQt9x1bGGDco0i6oFJ4sr9xmiUzgAGMyrHSXnewRXZD72Em8qNfFHkatkY3jq0vx2UPZOpy6
1Gj5C9p1XZt6q/SzhkjjHBYYYIn5kUPWNp+AGV3mFm03Z8cTQREpFBFENoUj1+Nb8f4aQvVmfpRw
n6H9u0Io2bCnmH+1kKh1Amrthknbww34gjcluX94LRGpAqQdc2tOO0+YoCJs8VMgApYxgMxIZrMY
vRqbISpoLYb76I70y344Mk3kWktdjBikItC2BBPEwdPnkLKp2CRb+Je746JUWSUiJUobQTn9sjB+
xXLoW3HZ+jHWNHFoa+wlZOKtW4j7CuOPlHjVc+bRD67F6irZnyfpC/iLRJzPdx0sTN36wQ/pXiP+
Q/m+jTD0hWlNiXvjrvv/h0fjzDx8R8eIQEc3dPC2puFuN4Pjdt5FZgzbmc21zXvE27D3yD3aHDYn
4Zo610/LCDmW9nIBdgSCwj1HVp5cnA8GQSETX9/Z4CcNyrz7+b8HQlUmU+uDO72MVlO3uYN6jIXD
UGskKSY12/etKv4eF0yHFSI6xOi4QWYtBJdi6p1roih9dz1vegT4mMh7jhkj6DBJaoMqifK4LYqa
BLgv9KTGBwRAUdJd05lwGdVOSa2mKlpHhuMNLQ095Z7k/EAqW+tKG8v0WjKtOjAi3XNh43p7kzoI
Q2okmCLES6+p4wNFQvunDLw3zjdunrYztSDPoS4NwmwL8CJVdxNLbtFoBw1KobglCzv3f0vVEnyI
7xJSUH1mylk3qciHGQ+O7XVygyZJbW2/hlHRMd2lwSQm20ZOPJJyDsvk/LsVIM/AuYxzdVF6Y5yD
ZuhfcjWyhVfzui2lBmY1Iyzf7j6yAbBWIwNZ+EDl594PZ5d8ER1NOz8K5vyhKVbYToQzrkRPWu+X
301oLYkkbbKzkHNZ5g3Uv96j9xiMV/DxkLjbaN2fErnjqGr8hiFekJVgrMxddPd0DqR/5jpNmpBw
KJZmEQZwJUGrDEG64+tnYkBBgHKlqmyJKrz0rx6/MLnMoHG4VnAIC/ej+CdrR1wNeQvTHDxzR7EC
SKi0uC2/C8y5NowwQy9aUNLGdbq6EkMWAMEf7+TtLBFAeRk8VOwWoEKanqUtS/L9lkdZYgx1Z1UA
YaDC7lNbUgzrCpFKa37zVIjVMXroHsWMbI5PfdaJ9QMYbj7b4L/FgBH1ZO0ITREKxuvMM25vryCh
r8jvBkwB88/kCE7B2N4HHwlpkA7IaWD7CtYvt5kFy8gxCRrMWNg7LP/NsIp+2G2sbxryoL6jRt09
YpWqVDL4pb+pbTmPCuacHDiq2QRTUxJrqWJx049pmtPrmHU0yULYk/uHiHI4PjIKWhwcZHiZ+fnS
mDlBqFQ6YVq51L8dOZ1h2+xhGhlSLVc2r6XiZn5xasyJoyRSlOkb3iD7OjLhTxbxeNzDgC8et6G5
Je7wvM0M+v3lRvpNSgiKUynCKX3BlYWzOrv1ZW0S+/U6/TUGWF09q84kdx844rMVssxgmpG6Fxfs
Ij0JwvFReL+3fShyrHJRamFN+w+JNE0DUIIi6RVia79YWPCTXo7bAzHPqp+nFMcHN2YshAEOr+5L
9DMrdKlbSC/Shi1pPWltPhU3F3nAHx2k08t9Nua9r/RLHwmSUiK1eohW2bkpYG1tk9pjKc/NvchF
+2GktwOl92Sl3eB+pZV/ubiolZMcVZ5fwNho+29K8e/feHD7RzBY/E46V7Nj+oHOwf/u4Nhn56V/
Uj4ng7Xiwn6oRQbu/OFppd91g8h52eYZbU9jsJ9qHmE0rA3s3kMKLKzJeWgwK8EZiqcr9Q3uCdSS
cYUItkKSGFr4m/wb2LnVyJn/0qwovxe1iS+/UU917QUwmE2tVto6+5TJi2E7E9bEbKUI879LVcmf
8/TNrp/Ty7hI7tFCnqPPkRDhfnb8uXr2V1Yy9ec4vxTBbExwedYBniUbT46hm7smwWQN3o2ZNDTm
STXXBRfwktkMwC3Mnu/y+UOSFN9u71tX3rBrFxcTJkz/4aK/j9kR9n21DDsKIA0ccUNA8i3N6fIb
CJPZB7GQw0QzEZ4uRB1NXPZH5D7i+j+hl/VzmXOC6SuWjkq1p1L2DQFamcGnA7nkvdOc8jQgsd+5
iO52iubrpT9P/82Je4V4XdR3IKpbcvvUn1FeS9T6SZYzJo46JB/2O/UopM9yniMOVXPirbi8OdSv
RUeTj3HSOlTrNwWkT3sPoxRxmlZFvSqMcl/x7BwbPxlSeb9neQVd4BERXrGk8IEN60ec+hWdC6rC
SUBtWP52cf9kYJ4ECYdwBbSkJGvQfmiipubGXLDImnPK30UKpuIxzy4v0WxJ94gA0lH2fth1IFxl
Q+0CCxB+b3+17jeYwT8BHnuHF4lSIaeNxhBHkPVvo5MywmSDSyqeuyjBPdYUW2aNU7eea8Oq54xc
JF7XvjhAgb801GIPjfwz65zDXtyZdNFzQXBXm0qKI0B69Sr7vYG38kJyzgc0lY2buA5+zwxS9Ebi
rGf7ZcjJV2viYbjETLMZFU0YA7bO3jEC3EktifJg9uoSyGQ9rKfpJ+ekuGXRVBjvdWbHMVhnYpdB
zi63f9OlqE3uXb6/52K9u3Ug5dT3DrHW67wtZyvvtPIgkW6pDexHxOI3xY/EJN9Oo9VpbrbAI/zs
OHfojGnMG9OmO5h6ey9jocdmlPTPUqRAvMCVYuVGrwlUFAWJSAghdHwagDLl/stn1A5Yjm+mMXSF
Pn8NdnvaeK3qiN1JsZ3iNsMhoqDHYyYlxQ4QerT8oWskvBiTgVb6aCSjMnDVcmZC/RLKpEpbLEhf
NOxDs4VxSD9Nm4f6WBNwu1s5QjWOa5I+DbhlR862vpcBINYPitFMU96UVcsECFa4CuHG5ayfK0pO
1Uk6ZX4F/CHR+5cPQSEHitLs8xIIrsZu/gFhOwy4iMjLfWkWrxY79jnKHy7XBk6gcxc+WrpbRcsp
f2c5dJu7hGnJ/IMpm5o7Rx+DRw4vc2tWKxyJGp8dv4jJrRACc9qUnLN0qd7trOlW/JTiPc74XeCl
CdHq6rolVXBFyN8N56q7srmnW7zLOYrVQIB7w8klQS+ANM7Zjttad4VUiRTKcctqyLxmpVAOqslV
8jyZHsJfe2BogE6nYfIjR85L4WtzOts8Lo5PHOu/1L5YiTUhZjEdsHyZho2Z52uXl00DWd04kBez
LR6gV7LP7FxEonxfX4svv1iK0Mb7OaXlSEhJVGtdXcf7tiial5w2jrPL2XsBulx7uyGITOIJhPBA
cwhjMV8ikN3K875qQ9RDFWlyS+ALhur9OLjYznqV7yhiBP2R4bTbvc+PkALbMnHf4rSaTEcFPslt
waRgC5GZxqZn3FOqAyqhLhYS9Xrr8KlVonGBQyIanlwpKO2VUlY3K3JwgEpv8zsRiz2NYIhVdpzN
AyrlVNopZ5uLT+VvhSjogYStVPsykGJ3sW+7d6wyS62uWfOBeO2+pwVRSOA2Xs/228KfVO3thsar
As3airwFke2OLeLT0KM55M0lpH8f/O868UYDMr/u3LsPKvC+hKEoJ8s+hLq0UGISipZrVg9hM1U0
1un5U31KWTgnrPkojX68BRIOlbXsEFWfFt1nX2gTK2sBSBthfvmq37s0KVjzjevg15CLQmuxDWb8
W3K+bNNvAg+Q+FMFoj9s5s1ZBjDcA+UubEInyfTSqMbNq+8q34Iyw9+f9v7yAeF52LYnV1DLjcHZ
ZnQ+KNBWacQQMyLB+qj8PO1wRpJkcDcxwRJAuNRs2vmgvJIKOsqbsWM9xEXcD5MyrmppOwyQZ/v4
1pNf48+idJD6vKAI97yUqs0vmv1EW8E3SV70E7AzRsg/J5absePlmb1K37M4FcYOs2aSDE4CVC1A
TkY3PmYyD7Y9U8qy5Kfr544W/FN+r4fxY3pSsch5S6BUrsCbYxrpQoJ0W0SZK7/UrwqE8KxDwp22
+8Q5R78XdLU3BgZHukX/zWBVxKisCSw6Lj3g9ZHS1Apc1JOOT1qpRRwNq8fdhuRpalX3W2NifaSo
fZrSWXJ2z0Nu9jLEGAnBoT/ZUJdZIXgGbi9gvR04EJAqkZ0MHm/DvUz7S9wc9qGhG7DPRLvbZwhV
mTFNZMTeZBURDQC2HzRi2xdWmQCX3sIEwVKlxjf3S66SaCnlEbYANC+mHJsd83hcmxry4E9chrzb
AH8QOAwHriDyjZhXgkh1l4++hOtCakGRg+QaSPKw8K3MXoA2UtYag2jpS16qUix/pJz310R2gyI9
U4tSl4A8FruwFTuDei7QLRQXjIMxMWr4Ga7OOqRW2eGy1t0MzFC1y0GXYBz2B3NdReM8P1VCvQpE
oeo2HHPZZW2otsmBwbVHJDqWGSdZOz6yqEjJyICKG+UsptErzrz8Xvh8xeO67t1PTdhraODEWyEB
APTK9NuVfeeVrQDuKPU7S6IBeBEAU9JvOegmnLmX69MoNl9AC8EkeHz/onXREa0Ara3ckWbe7gAW
Qavtc4FTYDmGyOzH/Km4uklnmETdF8ew6JU54/soz3WZFq6d0kdlY9/05mtmvd276DUHML/DAo3Y
VPpQCR/G9SjmlsFNsNzoRjM6MApPaRp99ODyRQTtfy4ygrDCEBJpi4kNLPnxNMJTSn6C29tIxI87
s5SK/xjoTWdVfM1R2g3QHTfBvdb0axa5nN9jtWlMlkLS5oK3KsB6UhYuXxxDclfJHbKgecxXtF9w
Ut+DziORBbnYLsAE0ZQFg85kmT+umC4M/0j1QFz5DAI6w1F5PxEXVmslVaKyhz9+VXiGk/J1Jh5I
H6w+LgpzqCwrebePrbuwz2OnLMDILs8UbzNGtJrrC4XFgik26cT3qw5XU9Uwp964QZqGKPN7rFdc
m9DGIx+d/7LKDLTGZQV0D9pgDT07hoSFifUknjzjEyaSqceZWMMe11VwT/yuNZR/WxHDUiNhL6Ly
e+qjEimbVfcWs2IdUd954PzUpC6yrf7dyjrJtBiEDc58/kEB60RUb6OJOGRcetdinxozTeFN6G5N
k3Ej/fSygAs12IDDvsmQx5hejr6y0paU0RMDKim2TkGGtVQ9x7gjZwarZ7u0EUqbbFNDL7ZhU/xA
egEYtWDwwD3vQHpCW/J2odqX8CkWe7siPK05iBNQwYCJI677hNI87x6jLcikRs9nQHdo4WP2hVJD
QudUCFMRap1Qq7Y2umzjaOIvxbi13KZSfSwxc1iZ6TeXGeKa1qy4O8OwOS/DoY6zBxH0dpWP5CO4
4/RyAnRmcVYxlrZwuc16QhlfYdOUk37tvMqiMmsF/W75vHH6l0DKe2K6eFDaJKkydrBJaCPud23X
o9hd0gd/jRBM/1IAojkfq6ZH1r2CLA+wRg7wgtX4V9qV9pFLdSIFifazXUa+NBsvwphI3hauqRVb
ul3LNbIA7v4A0YMFzbxLtQ4miKvhTFCn/7Syb1hsVY4Y4Zg6GKGBqF81k5ua313IwmIbs9aQEBnD
zqmnPjV0V/CQZWQyyHf8n1Vdtwj/3YFhyNkp74hKYxkieaKvOSvPqgWCnNQuy7bGgHgXe0CrySUv
YVb+ct71zukTCIhZsjUajfogkm5QocvXhCGF61zSZtNkYx5gddK+Yl6FmszVi5iLUX9enE6CijTE
vE7z5yvwZeuHGmHp64kn70Y2d7B7GZnb+6/hx268w6pWDkolP19fFD3H/s7yRXgYlMnxJE1SuYUf
8SU9S8HYsGfnyjOiv6hK8zI3VBIs8T9J68v5niqjnZKcrkpBBl+369lBVAiNBJmYt5YNrI/9xtc+
qeBteJhxpREc7N6IAW/UCy6v3qxFgedfukEcRBMimAIa+VfkM1nKPtOKKX8op9PSeZDIILBb+KxQ
wI5G8JcivbSh+R+6hmNcFEsiB17WKab32QXjmEhT+8M9u18TfvaRFh/0mrTUWr51GWibDOIGRvcL
Br5Iuu17h1jZnzqUxW9Hsl17XbLbMCsMDWjyewoomuoTEPu8C/+z64sYoApMjuyx/snrrckk1iQO
nESDi89En5cTdYTVqryxiFOQ9fUMYCBpVn15yhLJk3HWJopLLEWU0GiQwwLd1gTCsVFd/S3BZn0W
0wcc3vGcAzNfOYGS/R1DrGili6RP9aynhF/2Jbzr5K2gpUbib8cGgfotM/LSUVqW8UuyrlE28i7i
n/tSqRDPpLOj1xgqfFH8TuFr36KTxC2qeMZ4b3pqW0zrrNMGK8LRsaxAFA1RO51KeJOcqS1sKhz4
Jbei5BrdSjAm2FgbSdW8SzJmDrHhe7BE+UUjR2YgJAgt6xm1hk5+dnNtxrJ9HV+Y/XBgbWOzbcPS
P7cNHSIaAWpY9E2HwU7fa/9q0ogk5wG8SjXYONs83Qr80E7Nrj+hspGecv6KzO4a+hqVMv7gt87u
6u2xNjunotKkx0wKv0cRDEVqV9VHzTbFY4s6hpvRPeJNUSho+4iy6mC0wBbi3o2n9cfjbh9IkDKp
LTpBsRMkaYDtbgPE6EBhU24mFaqyuDsserdka0Qi44CfotyDmYdEJ9FXFokT0enCP/lKstgIb6I0
iB5kOQxXiv8Hzea4Lv+6YsVigeChcpIpsxLHI1I9sTcJ+T8ewFKOIRJvT8ltXCMb4zAUDyoVUWRu
J5S5wP4wGPE5YA28DXWPAHskLwKRYbz4+gdmabHMBVioTiWZCHU6roiIcBsi3t/XYyXkaDZL1hqa
e4nM2NivjBVfvdeyJEYIdbHMD/YXZ9MTSuQBQe4VK5gG5hIKZAEDFNyyrlnP8ZoHco2TKNSGEUIK
dyKuPTDEJOvyG+TiRDhaovg5l9Nuv+csbFlUqsZQ5lLT32oBAOuPJPXltFtz/ob7aFyc8wiWJHB1
CFW9h+rsH6/mIHR9goVsxF94d+u2l50hyG313nhrAlU1qOk/Mbze0th6J/Iue6/zmsoBCz6DSk4m
NaFPQSJh45nhCOUA6ue+pje98yPI/mbQAtSlE7YzIhlODSojq3gOVcYYLFH+q1ZOlSN9llunuH6x
xYP4gpgprUdvjyqpjq+beQsSxfXxFZO1mH/g0UW1rFfMDNuCU/2pnO5eyvFw/tVzl/e54Z5HEyoL
O57oUnW1gIc7OrBDCbLtGMay34IS/Fi1BrxGsP4ldHhWbqI1r+mbQL3rEEPVhcCos1o3n9qtaZfY
U9oIcaK8r31HY5D8nOHSfWD0cgy2XQnDEEhe92Sm4k+/hdF5OyoTejM0HmzwibubRmcQ0E0df/Ya
xniQNdImeVJ8aocSq6gMFEJ4eOCJsIb9aLckX1isSO04ct1izclac85TAIfOVwEJ/v9Nv8Ix1/k4
LzpOmtRtSS6raqFznC5YVD/o2zr88vvzhQy5ZfgNgWN4sbgd6mn6SkF/Vj8sc4fL1rTeSaoseU3o
TvpKAacaZfOptF7NRGhyzylbuxkCoYiEftokxQMvXDJGUX0FjPnAHE+7X3B40THYCFJFmHJGbm+U
uIIj4v73/Ww8Kk+tN9/Fmlmq0SHhVXFceeEF/pFOm6dQG56uOxn0E3cB4C5/jd88vKxqDVlHjeP5
/Bt5zQThF5r4p0PGr7Dlk5mu67UhPmHfmgkN5fVwDtSJMpKLGd/wB0MW9PktgJgNxg+SC+eNpd7j
STkOecEtJV/o1naNsYlatpS7N7l1Ro4OMX25lGGCWysUTLHVUPQMPewpsJOHOKD1dUb3aA94cglJ
GYRMdC48w3ATDG/SIuvNT2IjVGMb9zMyl7QTgc5mhF8VWp4ulOdeT9KyRlCCRUPtxBkse2Mvng8X
OVz1FCvXy6xh832SSO8IrEeimcKoxeJB66LJ34Hc7OLML7t5vdnQeJetDGJq1NFCF4FNT9aV9sCd
X6M/21rXcG/2ZxG49WcTBUGVUYI1mnaqRjTZCTzddM8tmNpq9wSahIRh2qRrAvyMDIAXrpXIsCO+
IeLbdXHY5oeEpBiVkaeasVaVG+BFE/UNnPvgfkbMOX8TM7SiLgKwCELeHw6oiB5bVBxmmoGP5iFf
7nFA8Sw7ZqgUbOmhgaRcgUdpPt99Oi0N79cOdvMiwtojEWwM7gxIcVp/a9iVmZ0keuugoZI5OIwu
V2UwrtNJZIclkXNt+en2AhlkVxRYuXuvdDNWxXwitSOm68yZYyn+CWpcLbbhIYz+dzaoTGyaSRRl
7WEng/L7fiFFQAGMhfhZDVKYKgKPBPvT+nen4z/60KOlHNUCfX3JLVfcWDDe5VBhBDaOSuXasN2Z
4X5BPFFnwcpXn5otEXCnidt50AEJM4D3So+JJ6kMNQYPDe1DVprLVN5qPuXrwErzGtmT++Gm3QU4
EN98G5GNtqhhe/MqthRBPYSR+dSlnAUFqB/L3HTsSjNMiTZ92JYViUEaa2aWcr+1wAB3q+l2LCzy
bNaEUhBNYmGk/Jf9nZ099co2IQQ3mnk8ghH2gVUfXM3IQrOakwHXFxY1wY6I+QutEyEL/n3w697x
kQ6peviZTMrDIeHuC/a18msKOFQdJxrUw3/XHQMvuBR4M8HJzaqE/hcEHRhYJpAbeRhstx/YyPor
dLpFUIbcFRQVY1GG8A3GCNIJq3uMc6LHlUrzt/ohBoUpntgbWa0hpQw6BcTOdWq0U2vlIbCbaIbj
R5ZMXsTpLGY3A/Puc6fMueW2COyZq5MaU20OKyGYKhjsOc/hsOIglZtCtieYzKkpMAdVh0DzuQ3Z
LuJ8HdXpQcrQFua+YbIAZiDpa6rZdq0PEV4VQUCXA+Y5wZJ1ZbSwE94vAvLhMWfXNJ4WKfjRRNwq
ll5cpMAV3SgCl6Rl/D+wZQPtbDEhE/qPJIueSTQnWP4fHzXSTDa8NisbmDsY9jFeplBsDhOuTV+V
tBoJcJZLWy/DyH4oDr8tqxJijxvOzvs8ypB+7SrnHpbijQ7t44DaaCrY6n43Z6NLVYHrfUCO1GqO
D++cZvA4a5G5Qd2Vm+aG8hsjxX892BLbUI41ki0Sc/Kj/1UT6om2Uhxhptez2wV3m04vHD235Xgb
nhHJ2+t5CELtOzXx/mwjZlzrpjBejGQkuUv0Lpynw9unscp+Hxj+Mba0zi85H429CWhQ7eG3j5Q5
tztchLe5SJ1WjR9pZ1PEM6IHfysfTZ0NQOjP7gpxYaEuFepKmaopIDqb+rPOaE2cN3moB0rrAGAE
D+FHMpkoY4konqPALx7c/TEU/s82gRMQh6BSFwZoe9eosWwdBW/xTeD2CCVS+A4YEZH/Ue1zx9yQ
pBi1C+/eyW/Q3abG3CGswhgz5YiQBhIdI32LvJFUR31x1ZaEGgzRlqed7Yl/ce/MS9sON4IQ1Plh
ie3Fcl7XRRWFIQMalLrjwZgHpQu9kqfL5sUhoBFnyOW+gk3C273Z2CyMc471XZbXo+MFa19giQzb
07vnA02nojboTp5rYAp0MjShJ8hCKmtKJps+ZJmpgm2D4Hoo9bNYoeaaRsRGb8+CyWN5JssSwAJT
oaNDHqklFC6cKBv6ZQt4romY3+dPaA2PtvKnZSVZY/v82vdEAv+TyiB3MqMUYpor6w4gXlboe92R
TXh3D09C3ZRHLXXOOzspI6Da2801qcifeC84wuBzm0OQ2U7Pc6shsq8qEYd8z+j8xrwT4UpZOP0g
RpseLcPf39H1q5ZjmIHBS8nI3AC4/JPXgHCIi571f3KTjzQfv5agChUcTdIJODwZcSZ/aid6xlda
trx7i2m1iRsHMpMz37Rx9X9jsad+RAGlj2aC39FxEVSzgxURsYWYvEtEE0uxkUCxa1JRVcGyJz9Y
KANGtCqWnDbcykMpr0M198Va0XHFK4EmXl95XPWULRqup62WxwRNr+WJIUmaeGniSFjSy37tPB3f
8eO/7S05s4QKhXteWJA34Blq5z9/i5f91Bef5PZtfe/IQrLU9YIZktoXmkNtskQ+TbLdXT7wGpez
+Hh6YvZwrZ4S+D1MDZumqU2Gt6Y9YLcy3dJqbPoMTyEbue8s5O0tvzGSJkVwlUmmIZEgtkFJqY/V
m2iYD2Hg75slMTaJM4LGMBY7OhFGU74HA4bK+o5KlkHhcvEmoAtjG4w6U6mwY7/yxWOGkaIjmAbO
3PRqluKUgqIQnQUwVAI1ayhLGae9FgOoaMPD57Bp66FZ1ufmQpkDpCfdBe0vPdajEHxHMQO1a8jN
Ih/+lAE/YDI2Fhg2ai07pB/Nk1Oxcx69EKZWhF+SmZguC/tjt6DrO5AoeuHZPX9yPWY2Qpv0IsGS
FENGSdxiBPJ8VCrcTJs7kPhPe5y8+bzgf7KIZKnRBLIL9kS/OHSpXsGPoTTQqL2JjWy1qtBvKWYN
zWoIYbB+Atbi6SMgU90WhkY5WxDoGGvu11n19sSl6TRCBj0ODqPrpR/JHi51J45s6xQ/M5z8t+nF
diIIA2qzMX2YPdGDWaXm+Yrkry5vSVJhEwg4wzSm63VSPMxlRmTmS9XtxP2MjRclSf5Ew/QkmKE5
NSp9KutQahnLDgzjOsnTN491rhMmVmRnn2elcTVA8S4U3aMYz82sxEN52zNQY3a28ypd8VVaSV9V
ExwxMSAwaFlG+T9deQ8Ns1X56A6vBTehxQ2LQVqfUbBHHVcOOSlYPrVlf9tFUQ15Wr8UK5IT5VJj
AMp5uV8Ux6NFl3rGbx9gtuIgk+KqGmzg0yXEjl59RjCvv3rGJcwTZlbdittOsEt0ICHgpBDhtHl3
9sSHnMfCxEGG1yapbssapAzXkwzhYMX7x9cMO/pNacnfLw335MJKomyftTD6QDJVPYiHO4mZ6dU6
tkNGs3H+WYRzU77oJX1HZiyC9F42w7ol3knblLfbkC08N/IBvsWthyeh5aPNa9avTAm6FfTO/QfN
3nJzsIH69r7+TqagZrA6FMfiFLcWEAo89kwmEuJP5p5Lq31i2FTRLQS1+MUNguSfjhrCJFbNNwu8
31RRCrHn6L+yyalttJCRx0kUs+t8W9G9LYATPmUEO9R097DjHnW5lv4PguMQePgU63Iios2Z2IMz
ediIRqgPomb0JtQMt9Sp25ffjlNxAmJEsj6RvG7epJkTgQzSvqOPMvGR7dMUkBMXCQeIHK3Z4cuV
zJxaA+mx8o63IIxbqWXaLG5QzKvO/HxC7/sXUJUh86HW8QcClv7vHHBeJgAjxldtuUeQJyvh90Ab
yNlAe2pHD2nEiS//K26wgPpA3sqTw7qyuesBrF1lbyowk76CNZfO5AXRx4tpnI0z+kn1zvQK3Q3Z
bMcmckIp8TDVfdmWLInDhf6RA+4mRXszrOHel9aEbnhuL8AGNnW8kUkPIKOpfzNMEpUAfE7IXRRh
lUiDBv0BlvnVCR50aJv+qvkZ1s909090lc3f2bZoWmLjR2Y9ufjDeFp3StlOhKg7b313rm5ofedB
3PZMeg7QxKCKl4edNJ+WjMsnLVR7Dc7ZrWFwc4qewwSDGGIYkam6K04TtfgJthQ85LuC84845CbM
zxhw7YKnIysKEsfwQRJAn9YhahYD4NPiabra/t2VHBkhhlDJZNSb95wrRfdKXLK7DBfuEo3+TMiV
OZG3kMb1DVaJivmZxMChyi3LhFvSQoJG1pcHG4sTmE/EEzJ7+x/dh0mhIaO/V3Xjv06H3m9XSCVa
ljuF/QtIz3Ayu9EOD/st7h91J1TzBXjDu3JPrKBW0qb/+Im4VJXeZtffEtVWVv8s3AIC3kdQhXsb
3A+Xa31EdBpFu5yqHesbzgQBpXR7XfDhoOS/1Kfqnidb5VGnVJRkDSl8MlIa6x3l+bVLvK9viUdT
q9dsDHXQKFjxoeANPwt7XOHcxBgL5anpItzCzDjRmhLa7DVEhcN2ly1JpcOpnE/yRHyzYyGH7td5
sK+4l8sF1uVSVyqSQv97fvZEWPM1ePRRxC0A4FYLad2wg8x1NwyC/x98OzYKnALRAhckcxxYtUh+
YU+6TGYy8b6QVEkOvS6Avz9ht44XJ04dRCdKYjV8VWYd5owgFFLdc4b9G4kZ4AKWXNuV82EwUGFa
WZXtXET+O2F5LWcRiCSjyigGi3UXMFpq/chEovGf+Omy0hpMfhcEKuD255Hkz/XwOrO/hU2OINeV
863aDmGFOcgu0w1h0xm2b2yk5P33PUG09Qvsoz2Bsld+SDKvlnZXcIbbOxkLqvzsAYxkL0jSnLNO
yRwgl+eypcAh3SZOXwycADkRHv/j9C5SOzVOVizz8la/ZAqI9CFiKKMtWpXw/WWJDnysa9X9QvnV
YHiBt/uZdf2l+VauSPr4+hoOT4Ti/rdhdoWQzoxNGQ4raBawf/eC+ZjIeshkFkS7YvpziiPzr9d8
fcN9IFd1AKPWq0femHm5XSvwxYgOoJoW5exFBLs4JnEg/e2m46ZxpZD/xUBw7KsONaaSh7Rpb1t0
udFXYch/9iBPtyDyE4nbV3eUpBhIoZ+QVWyZrYNlGfcHJOXuMcqJCRcdsX0Id+XZamba/BbTkVFf
S2X7cwUdPL6ie7bR5Oom8pLMnz2Wu/agZodS0IWzS7jolz8YHGNaZdRNzAmgqYZbtM2L39GmnrQr
C2bCF3/etSEZbOWikf0oomKF5S1Vxso9E4w38ia4pQIsnLpA+426l1D3soaRQ+mXwlNoZLo64pme
rgptrpDDXt7BcOTzIg4rrBfhzdEz3a4bS+dBo2HIbjO4PqMinVNPpjVghzXXkSSKa0K+odYnu/Tj
SxlqVyttY2g3q1NBmbRehp1Q4B06ooZcaiGSneJZgEkuWuFifqQ2BCTyCTcAA404o4fG/sitrzqe
DSEDqiqzPpFaQzKFBnu1VlQWgUog2ayLFF/oph3SGtiCRJ9Y6AZzLhVS7SspWR+P0pK3t2M0Uj/O
X1YAk+PZUySpU88sHvYoISHlXnWUOamUgYBMjU10GUdgAsUoeowZIkFCJjzotjDfVc0gzCQoxqGp
NfuWfrbwJgT1pcZtARknX+UMF5T6mZunaCfnNnFfrCtOv/smEHk+uds7WI+8/Kog9lqVbzTb1rSU
NEADKHrNJzCT6mmPRsitnrVsWW7h0++zOWgIbtDOnfcivHlNG9ogFNLOFyXz7FxJxoPkTVQ9HXSb
fI7DxgLXW9Y8RMRF28OqiNrnhphHwNvup7SjF9pxAwuuq4vIacSaSl5+/jg8igJmODDuF+YciiPF
8Dx9eHEskaNfICmaSQMgDNjlM/QYNJ5ZNJFEWfuyGes77AGc8z3ot7bWw8TOspwZYtqdP5uzKkJk
4OPBGbEbu1WFlSqsiUue4ZmUaKiyywxFCSZ161JDgYooFOyhaz6GX/rGJI56ESQpZxSY2uDULF8L
54xJdreuuexUk5iM13CkogvXGAEW0lJi7vtTzax7jGXchDEm5ImrGQIKwSj6wy9Sk4/1I3gf9GdV
f3kHKF1cnJXTXniDJtIMIFoiNLpK3rTX9ls8Nq4KJcVB8AacS/ft5FxpYRiBZy8UOsBLKTcNKhgN
5buA1rSHaP25jYtIpH+C79Jne8xgmUbdQK6kTRdiSKfUUHKOGA3jymFkRmrbMtR6EOcJUUAZysjG
YJJ3jK/hBzcILz2+8VWozhxGrbVq6t0nQKqW35Q8r0vs7mhnv6JZOAhjvs6yqmA1yf0RGCOWnaWc
ksneSTuPbtQvq0A9sGsBaqWbtFr7KBQFU3VUGxqMG2YutFgbyt9vnqdg9v28yCEllD2rN0bLMY+g
OzAx4E55oWnQLDiqd1wEqUx5qMTIOZah29Xc0xNtD27apEv3rZP9tCQIQphJ+WLpzzxUJeN6loe+
4heJeHkqdtH82Z0gvfOusd7qBRW6nUUjE2+g6YxdEV8435gAUqL/bI1QGD8jyfeoMzJMf6HVM6U9
jYfGK0QKJ5vUvfRQrl/Vc1/JbEvm6zYwdViP+bTV5aCyPK1fEoBHDsQ14nQlWQ9RGLvfu1mcAcPU
bY19M0fMKF+7zyBEMYQthlGDDx9ZRWfIPjt8PvgaTiBo5zw6d60LfjHuRJYlDNSbzK/yWaaWntYz
l/fGGXPfeepAswB3Uum5K8J7zHnUTSuzfZpt/ahiLflXS619xEXHKG+TPwZL58ikWvaFLakyJGQ0
3bdl4TYDC2shGJV1Rrbmgv6GyEsphwOBoyM1wAoGHo/yRPiQRxXwTz7xj7d5aS8XvJTJrf992dSy
jgtfl89JRAkseVqnuZ6HY+LpIrPDNEoowVJmObbfn7VqrERiP9tIufM6/3jreQTz/3Hcp1tWE1Wy
URnBpLLV0FmeYsKaXpOnD5TpAAgWSkyiGgv1zKlhn6jKWyqKx6hfMiwqoKM4uJiCD+xKYeYdKFsc
v+mZiAiU2+caAIQVj43a94COP8bvF91f4jZQiPCdGK9YslwtsmZPzbAZrA/qrX6mH34Oc4ULoRwL
+rZ1nKj4X98KFe//AsH+xwQ99GPpvgwf325sZHo2AaJMuODGKl1xhqwosO9DdArAf6Y1paHkSRF2
HUYK+6gTB6HW0GFswYQX1/3FEW53s20571Eu3Kf4nLhYqbPs7r4QY9i4H/zWAW85r7lNjcrxzWC/
61uVo/xNdvTiU2jSSemou+8HwRmeggxJZgjshNZTjkRgTwvliQxOqx465wkcxlyoOvhP1BPr8Te2
NXAG4Vuu2f25VHB3qSGUvxng/0kyqYgyd2+/iAyHOtP6O+1bMANo5E8NBlf4nphgchJw/cBtuaHz
xkuV8s1cH4yc1kXnCkjjmiSOjsVs6oDrS1Dor0tMHCLcwA5cTKosm9KFJy9151DjJes+kdZqLj35
kDPK6sQxeiTBsMp0Xdm73QnzMr9p7Q12ejuvRNtF5hlvaYLOj8cfwTxDHjpeAlkyS0y+eN8ujzty
nLjlUkyeqlvll8NPBpHb+sDjaeptHvgGg/r63jJp+6btTNlJy2H/Ae8EqPO9wiOrlW++Len7Qd0s
gv+35zda9Zg+TY0vMCHTOiXozcxe8eX/phe7uIHifzmamrF8Zg8RUriU5sERNDK503HoSzvzmR4b
qDFcSxD6oRFDb3VvieezI+MCPz0jGsnsp7rMA8wrUAM6apB8bHtWiEDKwoTvfOWqblcgHs3eZfLm
uhspa3AQRMlHEn9Lb97AmFV6QhZprwKXUT5hByDcDQVv1xmUOxUDjFURrebHRM2AsNV/oOLRzEJ9
1Jd7cCP6O6H82VEIKTfN9sT2BKUPKHaAofeqUQoNixP2tlTjaVKOG8ZQRbnFJaXyUO14NpfUe0fr
d6zZStA+3AYFb+nMDkYwy6L9pyANmt3qSwyUga5IAbCjUV95ynGow/u2AZpCmm7Mguvb2ufy+kY+
RGnDGJqOyAztKcYfc6NRTcrTIA4r2p5qXBHcL77EMzEZ/sMrbiTTNLQDwRNSbIQGlPRl7VNNhV74
DLgO6K6/Ojj3o5VOngiweqyFiVaaGlPJewJchlobsSbljoCZ99KBn5aVQ/ypzawmQYRVRMLzJbCM
uQH/W/j0w8A+X1sgNrCgue2b35LwpW216rl6PpV2NUvF12SvVwqlbfu2w1GGp5yIhaaO0jJ99cus
ooR3JoxObUb/bmaWVo39HJzH7UNS7jESrjCTw/zGKj3fDwHbDByuh+SfdHkz5qhmEWdM33Binzm5
DBKD8LlPRug/VjNe2sj9vW0Q39fknL4Fgo5c32dWIB2u55Ywt4JWgwBVmIy7pdDVpsvV1px72bSh
aJS/zUVejF+zbK9x9UUlFADbkNTu1+g/dSvpH7UzVZ/kpMeLgbu3zVJyfl/mJ8+oNqKgoUG8kQIp
hXB3jcV89k3hGUNiAKYVP9LqDGCDsH9yhcIpvCRy2LDlhh9bY2ut84251NnF4RLYhLyCHDKk0hbm
gphF2RuRa0Ot2tjEzeg2qEgMbpxEQiTbWP1BcD65Yd4Kws8NbvxlVyoQslUqTMuSrdXemd+Yyc8l
yf8dUns3DoBj3y5S3mtK+6hbRaTeop53+NJB+hPZcEV4XPcJsXtnumehvwiVuluplT9Mg4sQWI+k
rCqsEvsDWVgwufDeIJsEVD1VgIUtqrCgCK49eOPLSHVWH9HbWKVbw1dgZetDSKMw3POIkY8TUl/X
KafrgkaxZjSL2UFRyztKKRWbe6rKbiBFWC1GnIm77mdVlCwm28t5BiP6nh8syx6FjkFK+6jKJ7w6
BLe/s1kX4rixoREAaXyea9hVBG1+ZJRdMa4GnHxTHkNsQC+QdKkEWYXWtuX4T0V89fdyuXHDHtrA
hyqcOHKEJvsDbsyOLdNqB1sfSwkiEnjPMyYOsXZ3W8SEVruynPcv98XINwHqiaItkcBx55d48w/U
Z54FbtGKyfvb8zo17/fzWqKg4uewiwgiCW/NU1e3XMKpREmrEkQy3bklACZsL02g1XOrSEaTrZMn
3sXN+je58Nz5wu6WgN2aPY/1bFhpc1duQjGhuVwZRQmf0haCcS+I3h1CB/ppeXhrzoG4YZQZyp/B
e7lbtvqw/xgaZRIa1I9lGopuJAVY6lJugP6LKbAnmfVKb40bNXSz0GCWdRfTOATd58xp6ua2ZKCe
JswjR0cs0r+0/w23UWmm6BMfT2hnvoUARBCOP7EccN7L2TuasIhG7FR2oicI+N3aTZRG0P6BgQRh
ocuAbsJHxoeLxmCi1/5azb0690BgaxpRcBhmATi66XHp4lfxP66OB4yWWVu8gMzVQ8Lh1pdtqORz
ZeP/IkzKXj470cPp6qpBDB8Fx9F54p1cVL4aCWzzlWMtsM2U5/4+yG4KzDvqpK+Dms0WUmWhTNTe
l6iuI20GHiCKkU5/56ybWddJYLUd2jDf9ZaRB0xgIts2W/rv1MZJQxiBhKOZGrutt796g4fsuwkK
98nF46ZXZxPJ4ZCWzazpSd0tRNe3kBgvrfANdz3uSaoiyPh2iaPx/lXtigC5xXvQS+en1wr1PBvQ
dd1dd4F5l2/0nEC2uJKG9vfgt/x+x9Hfm8Sm9bUY/kZMO1+k4clkcfbTHb37WDfNtmN5YbIpYxnm
EymEQOcBA2v4hoenL16gGHYp5P6UWy7L+NLxex9cd0kQBXZk77kmuwS44bzKNBfUP65YNJpDPWXn
AyrYnA1m4M4DiK+HEygrSZ9Uodox+7WmDIirKzo3lpJbv0kjpMF1wkx5ev+uXJoITBcQepCrQ1B2
o08BJ1jfPKQySBOx9P12+Xe00IDxgJ0Nt5YnpgNRmQivgEZeu/q5ISJkI2bbBaQ9dnYf0f+PMAs9
WjnPKgHq3o1iqjCRxuPoxMiKxCEuKO18b4cosmheWQ+nxQeGO7iSduPvcCjO7ZWMg39aBoaGnsLL
AbV++XkRkjdot4BkLdfXk1BKOEXo7UmE/hG9qYZAtMa5wIy1iXt5fpsROruOC4c4O/6niuHn6twV
cWKti33CLtTaNdRrrFeHrflnmUdgMer13Xr7lumgug6z9nF+A1L8PbysizK+qBIiFDS8NGRQzq+Q
9xP2Z2oqiqirKR9BDSvApgElzmA+GivTgAtOhET/jQhQs9bM2CjZcJo4+Pl8YlGy8eXUXgq7bI3Y
ZdyLvtk6ctgR+eRRO+IgZRm0iXKa7PcUef/x0YOgODSrJR4h/FXvzuGjcAO2aXeTtHo6vcMgAgja
p/HtbXA49/7jmzIhO0y90PmanMn5sGpcwPb6IQa5n6SABxVEDmQ5lchwhev+K1vHhMK+KleUv0HP
qEFUW6cms10aolGUBANyYErXklgcjcVMPYBiKeh+qkpgAT+LEQY3yRbOXMeXk0jMXnCO7Oxuct5K
vdw7eq/WJCl4NV7X8geFRRaxx+h8JS5raFQTy2YzJDeu7eETW9SMypfr4yDLuM7G6GW7tDvppK5t
kuonvqMMCGgt1SlBoelJ67nj8uyuNkkypLcmaTJ9r9I1zZSGcCN1gxIFJOdyxOXXr1HVirVw6+Uo
EeYVwweez49zaWLUCCbhrGbPM+tPzoUj/q2KpMiylyBH3PLt+PA+b5kT+bakpdpF8n6oK7dA8uXV
oFUVNnjMNrCfkiLIJuQXWwh7gQzsobwVkNCfyRTY3FSgCm0p3eDGZ0sPk5Bd71DELc7PhRSxGN38
lrOePhVE8O1SEG8wgEb77XcsqAqriOtbLiKI/s+6AbLzV94znzf/P+sPSBv1w+wCahokHl37kJO2
OFz/ZIf+lJmqV3S26FMTqba94CnsJ3JLv3nU+y1xLxPWFiJ94d4G+9exz4iJq+gQI9HF9QlW1xGF
H1Bv8GeaU9RmspZNmpDRIJHJ4h1rLOHwVN1vUC4gXgP+0VN4LiXdkGjKYBxs1uaURszxhlkROrg3
yIHL7K+KfFX5qLlK6NALY2fgtb6KBMN0Wc1Xz3Wpx+SJOKn/QUlzG8r76O1hHa+aqhJRSjJDLz/D
RVEIx4ssGfFH9kaKRV4is6/Oa8ls3KTVHOTUtGacxEwxgYoX1ePkKrkIUqltN8mYmGVsQGg4i+oT
WuvUG3Okz0+NsadgkG95h1oQU7YysHVZEo8Y/+nbC/JJklNrvRUlYhizTGRYMssV9PO6FzCXtNc3
YhCIeHNIvt6HVC8WmjJgUhfzU/Q+LWMyUI5SdO4frIpX6dfsX/p/8Yx5clrORuTzmxhosY1urRdG
7ngAk4cSQPVwh0rLkAJWEr1AhrMVooJbPNHEap6uTAr4lDYRVhfSGLLgWg835RZnxWBpOW/Mw3ld
3bls/5oihA9Vm29ffNTe9bnDGvP5CqO9AuzB5tGDaD+V5KWsdy7ktJf8JMKBIPcOoBCrr1/QQTwK
eeWqJODvmHPPJwbvNStAdMQarTmT07K518oenllrxRnd7TBpTtUIfhksDwxHwOkXsqlhlOxNE66l
MVtlSFl/UpW2X+M4pnZonMxwqlmFrTcBO+QJRqsDABVMf/XeuIvCoUUJabF7+HoWChZxlDIdblmx
v9ol5k5yO3hC/gbksAvG27B9GQFx2716ViI0exa/nYgYao1wKYeutVqK7yOdeU5xAPuimu6AfOGU
BT2wlEVWoKx46G/bV8dbArHAQjjwIutjDCkO6mOggwWj3u1l5/D1QHUvNOsX5z/bnfVrcFsZjj1J
nkz5IYHJYckA+Mzq7N4g/vsKYCUP4am/NSsckkWC4FXWrcOIguigfzVp7X3aB9awMG7uYPeUNp4n
GcRjYrf5WP4/jxQCDAwC/HGkoH5UtvM3j1bMgXPcXwES0h8DQiGE6EpjTcRrkL3oBZw/VtpP1DdR
VDuPQ9cxt28Ng+7SCGhjKgT1UvRqbLNXiMl+B3pBoU5ve/LjCT+2Orcfh8S/LoI+PYTZL/VMYOc5
qbQZCP2PgFpv/BcPAwpMjIN4vH59xbrkNfH/dDL5nZ2jkVq2tNvZo4uTsvl3v5IXEl7VVVAoAbcm
XxEWZi+lHbjCCwAqDSIgBhLF+Hh8uRxonzAB8Z5yjOicQIn1WS8Hrrk0JJ+jOjA4gnaK4Q3E11xB
O6wlqK6WJjbQuoVDhn/2myVaQ1c8VVogQYBMeI0J4lGOh6DteyOBoX22RHPOD7aHsWV7Nczej+9S
fqgiXg2ks6ecUQtw+LDllphJI04U/lw9I3nOprEmG7DPW4kkxOoj3gHiBxpPfgH7Vm5561DNuQJX
vwOK2Ho772sX+MoCybeXIxM7bti/fGvrQUhqNGkvKmJpgRkiMZiuG+7LcuNc+0IB+PBse12XlEVe
XpMSB+DXEQsz/o1mcWcyLf97kg1IvZq8H5p0E86ywwq6SlksfYwXc5wO9NNqYREOSF8KordpMMap
uX1aJp+xM0HFtAEZowvwiK+nqBoA8L9LV4ZEivZVDmhsbobjY3TYVkZQCp0K5e3cJQkYW7hEx9AA
GxpD+FdZwzgkDNoZOMX7BK0KbfEcoqhCmifkuKCL6fHWMQCKE2RgGHJ30wVajjaiDNol7jnEdQuT
7XC3p50IQSspdP2CQLLILa0KpWtB3dW9TjPforRcVweyTXmQ6dKQ5ABueqZfgyg3gZmSPskRHo8p
Cxm3ZfUTZ9lcplhGbBzK2hQLeLFoFT4Mo+0luAn1czZISZSVKFNVr4nl80+1+1yzR+sxLC929gy2
eS0H/LmMsLN7wcCNl9gTfbTF4VeCeFMsw/s2UfYCBpHZmdzcZal3v1nCvOzXHSaEs0FW5/mGF7o3
IrhaxmmyRvSgaWyzrrE4DRdSM/OLZbq6dOEK+Ns3dm9nUnNdDgZbaR+hwr+7OCfucPvixHoq4kIW
MvQ2N0jIDuxDZchZGPqUP2BDNyoFychZtVK3cx3KomhSpp7wgexj4rV9L4fGmgfo/6sTyGpmO/cN
amgfa7BjsHVIK3f+lT9polFSdk1YtR3P6bQMUpqjQuwJkG7veyYjmaB8nvyrMWLmTOqrpsqPqQT9
rZuVMPmsY+eKOFl0L+gIos5+UDrpcpj+ERsw05LOpaWaAn9TBnZX3quqGSk9HKhK7wFUAxV610Iz
8jr1wrEy8rvJuyuvzkcQz0pvqCnTooI1vb3NAWjbq9yZMYnNaIN2+ScYYg5Vb3jL/u2Qnvrgf68o
OMXEC3IwvMVZxnv1Uq9qj3zHBVg/ASwHJipe7MRI3WD6/hUJhMSAbHSmGaE50Bwez+IGXvcdEqnR
gj3gbtV8tAGim7JKIHNmfZxP/UpYMVG/PZC73QRpcbMHPBZ8QFjdZefMKAFnSle7w8uZfn0PzBJ2
dAZtHevT0Hnxh2R5tJy74uLTb96jtp7aliIUb3wlVjECab54atZ79uTknXDgBDOFa0a191lqdY+v
hVpkGJfiOTXiogOhF1R0naoxoBSu+HaZ8b4eCdXxp+37uN6mG0Vq5UrGg2JCCdsTdkIjBsgdKgj6
NlQCKR7V7oOj8bpozIDhSwU1uFmV+kGeBjIepK3+R1URWWBANuTCqvIjZeEhRSsxdjKlJJ8w/r7s
hy7vMXKa3Fp+tIwSzI0wSj/lTE0ZfHqMxyt0jAg7RrRfvPB8IFg78z2CzCpRUguENELf5rzdshIr
p5eOaW1wLhAQH+EfGQp9wwyiyvg40VIbcWOfnRjYpuC+uJqpiUrFnFnFTxB2aGP0a76blnAC85cr
FKqCyAmcZz/bXzO57ARdWV+pUB2lMGBpT9gBJYJLo8vQ9bGKGr9n3rNb7Xw7/UtUGttuEsLghn8X
iLX0cksxkDAI5knfTZVySwFdqQJbTbQs7cwKrvcbUyR9UARdP3gT5Fipe+atts07KPqOw09hth5E
IqYrgyjHO7MkIjqOZqKJQZfE2KMjZEbl2i290KqCOMc6Fs0E2e7P1nmKD5dG30HBXV5/nZwCgYal
1W+0lM3I+XMuIm+T32qDK2nXjnH/zZNjyloIaZGiopadRvCNjpZOFiuzsW9Fy3NtnViTHM+keC7S
HxFdmVugGSwskkeZaHrHqjY29AthfjYF66R42jgFrRgcpgR0qJfgSQSvCvBEalr1w80GaoIfr7Xj
0qhzz43cs7LKVaS7ESd60EONZQL31pOSls2PTCWZfZyvz+p7X1aqfhnYRT5IXDspIDSe+nDChvzx
ACnb9GgDHzg0Ybo19+BMtziTIqbj96szWDBwQ02bJcd0YxIZNbFU/4mPJAekRjWDTEZZKhxjnebF
q0yzDixzBk8zznzEUb8fnEEPHVnC47CN19gjeJJP4QV2g8D/C4W+FohzkPZwL/KNm+GxpXp5qorD
e9FlvHMWMnT+VyAmtwLvWYYTACuKRKJT2iRxcz0kVRj6sLZt4wvw926tEn0Jm+G6GbTCYbVGZb7R
tU/hNF4TBlhi2Kfte9r4yavwIw/+elSnKp2yGvcpX2V/OAsvtRSItgOiCHbhSbgDe1DsmfN2wX8m
3JKEhku0gzv1QXKIBVDqGiEC6QEapDkRx9G/W8VM/HaFfNLp35w6KXFz1DBEg8y2U0grlhLJKPpl
hFkxFoIAkD0ygjxCpj/iy0ko1CcKDQrEQxWhaLCcg+LDmVSrVj7V9jLs9EM+kPsOJpC0Sa3a8dYf
CI9aNE/R0a4/YZJJ+Br9XoTm7dOEFqX+3UWHjObR971O+6z/bDjOE5m4Bhr4v8vpkQy3xMcTvTiS
I6nN8cTf59MNbYYX6ZV4RwuKp3hK+xkXt/tTLxd/h4c/UQ2fin3h9j6Dg9A79+u76UYWaa9mKi9B
qBwMBYg4jGuaKAzjL/iYIA4ZQJyArP5kGJEggSM1HmsNfZVWeqPCuQwha3isWn4OSL/bhbMNcqPP
iUJoOdfu4bYpPNbMYwnvHJiK2ydGySmC4EBdtzCiNknHmQ9oYErxQbXZ1T0PO7JGwMsrDcOPNNSv
6IWbO+xrzAmBH24K49bdPUVq3adQabyYF42SrsNIUAFtJX66E2w8YYTxp2nyecRXwvFJIAG0jl+Q
Yv4FvhyGsyrsMTP+FDA9jET6CpYrxZlilxBoR88aeiYyBpKXn2dnjHtlNLK+DP7A/GvMudWZvxj7
mcFnJBw3LL/kEiFu1g9YoPMi2F/SlV9kIRaNh95LIAKvb96sYN6JjvL6XSNfI4tRsq1XRHTuIjcK
jCZrXpb70t5JRl65/ndDW4aDCIYrfX5K9H4x0LowkJt59oBp+nIw4Kgvr5RnzLwLU66gKiKJQ38H
ja/b/qzk7CcbVUnp3oofECHvmCZe59xuotQJN4F1fcg//tykhxkBK3UKRrbq8ZoveUAT11cZsJBB
WOucTux06Mvj/FqL/4Trvh2jZpYw5+eM/SSNDS/OYxScLgF1MonqknYgnvnlTT5WoUXDkoCyPNMK
VFQ69kj7bBXXPNSQnkvT0kIaJwvNV/SMkAJf7qOVS2LEihyKwCq8t4N1NHmHpcNdb/+SFvHILqAR
ASvpxLwQy+g33ZKE3Ti7KCwWeqt/Zg0sr9bq+5Abl6QivUn2brZDc3coMYP4feokr6ZLTDgiV29G
zZvKAh+EGeLXx84e6M9p08N0K83Uy8W3HHIwhkXTSx0nXzgR1vb/0yjgtxQNr8mH30CuW6ctJna7
P+EpbUJsVq/r5BheKupmjh4wvxxz3DlNOscPyOAccdDvED3VBeMNRz4SKrRamI2rvKuwWr0wm5dX
hiNcSd8pakywkQB82wQ/C1pHg7ifXaSWUAjavx8JJlL4sC69BlOv3Cw+gmMQdNi+Ch2va/V3chC8
nWXcI1cAoY2IwhY2cT4zzIjckbrAONmj2he9Yletu3216VLoXNFDK1ri9LbnEcXvcqAC4LI6hi/k
aAoU0UVtkHvMUtfuh0nfbD7NMfGu9O6gG/r/PCIBRw/EBcFfS1IAZdm9qzYaWtdzEeLUwuJLe+sd
OF3QL66fDtG0IyWpYVEJi+pEP3D4KsQaB4SOVV90h7fXSgogmFW46Ts8tiAXiLep0kmiMjsWF+Ru
DLzjiSFGixJ1+IM6On70Mr0bhoXLBBHbvbQdRS1yEkYJdlehHxcawdMivt6M0czAgKXjbQhgPb/g
06tpr1evt63YkNJdfIzqlWUhX9FeDrW3/xkx0WVMxLhDE46RjTkbQ/CsVKVKRG+EntSTPDgXAQpp
WLF9Sf1g8RtMtaJY3/SFNVbj5w/kPfpvzgGVY98U4mpfTYiBaD9wtx39izOZS5OA/xddGONrBMj9
NA1OzOz46kkjKIeillHOFB2VyeTM7ooQlWK5m6GEDnz00J5olNIc63JtTh3xkyCdmSvjpuSqG7/V
xP+Jotj98RgDYMyWfGnby9fp8ZM+XCcfc6c/eCvYuxY68EF8I04NIbICvwiMy0MgXOBpe+mzS2Ic
cbuiOXkAgzX4KOUxQuKfv+GHIp/edchs6HzPAa1Ew7ulBizS5Qj4Zm81ebL0neHI1lhrgSJ7r+Cr
dO8DIYSCh75z3gcBIAZw8NMJkqpkhrEvW2vGV+KQHPsQFW0jIryE4rv/L/7xfFTmGIISvItWbgWt
V7yofv1bMLeA7/CGJL0wgMB/wcxRz3dOLftNij+luTJAvQ8gG6A3BLN8Lwj9G9GbRBQjof62Kf1V
CZ8TN7/5D5pIU4eVAfMqT74qgG7/HariPuNdX55YNNYB9b/TKOv1NOa24Pr3hsr+4yO4AVgk97y7
mQMlWstjpGcmr+zXFu7lrk/fQI2uuGU8LDLBoqqIftTmHoH7Dsnr6IpAlyssRxHdOEPrCi+rw6p9
72Wi/bEGPD2y8+nXRPu/+YuvyI2ypwP+L40KBG4Y2gqpiub1yEjay86hdTy/BWU7hrnBNPACHd7m
gbxp1dxEMMZjkvL4bgDs1JbtneOZwAmkIrAWlITHXCH6FWlTD3gLlhGrxco6ywzaCbL5JyYgPpYj
ibG742cWFCWkzyAZcV3TN2jtto+1i/DEbdNhn66gjOQWLch/nLr2371VKq2g8ix7BFJb3MVO5Q0Q
IiD5ckyigSZeWxnAwT0SAqGbQEGN0zWAzm2xTC7KpVWwFgZPmzD04CxIEyTU6S2+Pl5tptTCIkO0
ZGGxb4rinJzm8mlCxCGVPRged9NqTN9Zw50ZaM8OZfB6ARW5KhRbjmv520hZ35pmhWh0eUleX3Kv
gpnFRZmuu/ua3oiFUQyqo1fMg9aTdCoLEJfAmwFwwL2oVB/TEKOuhSS02RLqG54Mnoou6LoiwuNI
0lCwTZVvdklackRuJ7G9VLWOBi7AIEiUkbMignK4L1bjDz99rNTQbW2Y5VsRSV6R2fAee0bEKYKL
keD2pGLLS9XSWAS2Om6eyjru++bq1Bax0CeNm/F6C9Kn2fzm+EnmTZFm+VD5QiAejE5N6JJb7Axu
btWpKWeMBCV7fQ265hb6Wba1y1kZj9iu8qrUdokDC5lKHpqM1/UgNNjfgbMM1PAJkzg5NpJp2l2c
N5m1UWKe8DwrDyPnmG2cTK4Zg8FG0m75eM73p0g27BMUWof3/V5AwYutitqUp+uZcnOGShbyxz1b
LYqG9BaphbPzXe+NkDeV9mXHwLnteECvZkdYzxikgMIjqq3Fu8xX7N1zcLBTCrIehw6PsDDvxOHb
X44szKaiROVJ9C8Nv9f9rOrvHIE1OBkQSfbvl7ubd4Un3ZHBO0b2CqkZA41JdWuGFBwKX0WiGwld
HB0IXql7zCPUqcRwL/X+2CGXtrdOHFWn1+ros61F0DjvlbqrFGGtlOD9RMXEOCUGJB+bDd3eq36E
HmKMKFfx73V6s8iydcxCmtxmm6B4ZYP++Lq86I++Sg5Vom/5fEqcnNdFZB54+4hjN+AEBbBMkiXt
iNyRHDb7QYXsq497RSpGf9lNxxrYuByGF/ApWrsP2K33y7uFgr31Ubxcqa+c6W97i7J4dpaWrMKu
KTb+UH7a4bBeBIBRX+nK66tUCOGthlxHWYbIY2JsE9VZfL5ejR3gu4Xcmc6q3N9J3u/aFo84obeO
VIorribqLdWAkn1NkOzRO9fjIoMbHj8Z7QhHswFVYSftOsUD+vkTsjUARE/4Mve0YaCEHT+bMIJ1
tUBhz3AV5RRZr0wZbae8zXdtbBqyzf7Ix29r9f8VFn9bBuZX8jhAbe9jThXDJnamtJXo5e2TTjql
w6M5K0Hnf8JwtHCs8wtJ0rjUnJniAwUHzSOHB//6pC/5Pq7TXDfsURu2I2H8+LNr6QO7F3e1b0xf
nBU8Ks935a4HGhHVJDs571Fe8dmXNMu4vzxAuhKGv/clcMhGX7IrPtRgg+A4SWSCEaWmh3YDKNoZ
KPuYp1q3TUErN4PXVEOq9jgMDgqheot7APfoC3x7zGgpxG9gnoTfPmMPc8jpyGvuQsfVkccrm2SR
XLue2HEaeXVsW6QLuQqJrTyn7I/3i7SNZxos1aCsTSJi/je+XXFgwnet1Df6e6ZHVb/z0VLqL6/p
CkG6n3H7runzFhuRgQenQQbZgwH0hg8lFe82u1dOrFDTc/rqNkdmkhzBJTpbpgNHipqmrf/QyEkD
m5ebXKzUbJsUihm5pz0o9AQImuFGOiJIF7w0LC+cStJ8gH5vat75Hh4Wg5Ss92EQd1ZcnBHok48b
Ci5wFjcQYvw5zAQP534XX6PsRq9Umd+hwe0BPWEu3bY5sUF47LJSh2CWuw2koYwRuChoju8VUBdU
QgK5nS5/XmSgAkD/2maAiG0v6LqgCKzZs9WIF+3FjoQO+u4IE64cJM9Z4dzamBwKpbOzIVtkBoJE
vkUlK8S4as4D+I0/GOVmolgO8V5teA3fCwAD/FhJhrGjMhC5YZwEPMrnQKdfd7985muZO++P9nVB
h6mYDGan29UN1BeXdG+gI4Srm01dTnBegEaVcfYj4fWlB5BXf0WzYRJA2cFElBMyOkAxkON8PRmc
UI0Md/7p/UaGuD6sdkSfD8gJgpCim+YlxaAnbLtkgOlSi0flbTjkq++dPA8LbSpXjYvr0aljzlds
v7LD6zCanNlfScEOhF4gIEBihTcVNgV0XBjGz5AC/tFv9MZalEwk5lnbIj+9gfYCIvhHcr1n9W5e
MYjR0jgtLNtXa400CGIgyfy3Nyrt8/TkUxlchjXA8H1/7vD061ozSVV1JvORaCSczXN6dbhGSSo4
+ouLQ7jY9PSoITSkp42GilASPZGA0FAJ4gkY+R+psCkO0UO8lnTINrRcON374YuI24Dcz8UEO1fp
1biNUPDhdJsvN0NXPTsEoLpKTBkp8EAd4rdXLUfKHT72pj6lzTG4bYqhmSkb6c7XRYlLezvB8hWz
J42LvqAdQDRzu31XFV5fd+v/SpGmyIvNrWV1zMHWSJs3srTwhE/Fau44LqmnIgP0LQtHyiqKNCC0
WJmOf4kekh+ByUvkhYXwgf0aoVsn2k8HAFYWpNpdF/KgP1cUvBNL+kIzzDYqwom7wfwPf/eOU/LI
YBwdoQ5uurZBzvGplC8MzSXN8tXSdk2RCgdOYALz9dN/b4KSlrjxAmXpjluADMSJFzjp6yYIqZ5s
qF8R/hYKMs4IXoLeBBHbq9IvLFDrTdV3rUryF7xCNfc8gpIkY6iT243QhGmImB409mas4sYpCoJO
KYYf0JWhAikEeYcBbNK1P3J25ugajryxMpM4i9CiI9gpJTMDTkLAuGYVR53xqIUSIMGWWUPP4Ncn
uW5U6FiShsB234efHt5QcqifAWm5fXJbW+uuRd2zRydFWo5FKLbJ6iQw1HstwrqggGtYJ4SUuZoR
49wReGGnTHStSVhqeVhEz4IN5J4VkHqu5dDlyZiuZidWGLTUw+7wfnLWfdZMy9LOzxKxEVcEvI+5
aMh8EQ8cleSdMmv1fvXMspN65cEJqPq7+l6oDIZEyKcO+7aoAkpJZwp6z4MWy3piXkEK255BhR9K
DnpeDz32OQJY0m1lFBrXihoYcmpBqGMO8EcyewJTv4OUCjkTOIa6/iC08bpqWaiezieXIbBaKbYQ
82T8VKetiaxTBZ07AUr9YtanfILRn6r6A/bJ4T3WI1P4tH0tNUai/oO2S1n/orwx9FJjwnRVTJiM
p74c7MfV8GyiYiDmzUXB1V4jPAs9J3YwJyuI4PdfVwHRA5B6XyWZqhwmuxaNNTNNTxk6rAM4DXb5
sAwoEIWiSTb9SuF/Nb2XG+VL83UdyYfb6kiAG55VsaU+dapjjtpBywLz1Bpc8l4VkG1c1Xja87j9
mwk8Qq04w+sPxkZFymFhPXf9VXr+BJWbt+OGJIUDrWOfFF/UE9p3U7mO0w5iWqmDFqZ5VZ1icypY
PEWw+fddx4EA5j5RMcPMKXUOOsopOCjhLgGa1wEPFeBdhShJqJwWg3oyq6fJ6xOBrCoFnu4QwZsQ
pLQtTcxKSZmiUMygvECr8QdsMRbI9DfQeUiVvTWRwLIjvEYz4Qp3yfoUaDxos2Un0uDLBRgYHF5D
dU9zzWXMtsqdufC/T+//ltZJaBi0IIkiGwRGWLXWfMhI54Bl4UV5Dh75TID8XkikNS7CaYxwHfWT
L5qyI+l8Bmw/Zw1KV3SL1E7/g8TWuIgho6B/tYDcNnUE9hEAn6g63qCN2o669waNoTePQNhzLwNq
bE1v6t2CCWMMzEl/MQUUBHRtfAlZ6qRunGg9Iu9EVPg2RNYpjIhIaOzL7DlpqrA2ayaapghEdSLU
zUDSDDeqX8B3//0uUk9RZ94TfjyNsGohypb79xolUr4pSYQ+8n75BwgYmEN8VEbyMXXUoV/j6onT
2CLpGLFMWA1ATPb5rss2Uts0RQ9r20MI4dFBVrAAPz6cJ24ihbb/WN02VkFPzi8KvngtT40W0r2N
5Oq085AXybIpDhTAzoZBfg0E042vyxNT7OqexE+deZzPsfP+N5qiWfQhPrBA2fNLvWTgIq1asf0k
fUGuND0F7TxP5kfu02phVfwyGTJEaQ7jtecOv77Ywira8nPzh2keal42es1Q5Xz3prFj5IIXWhvz
b3RgjJDxNaKa7qNIvcVzxqKhItJaFdNhNqVpS8vZFW0ekP74Ek/ZXv5YxPgsJ1MQg+vez0+vekk6
quU/CYVwch5LNT5ewDNzWwV0uLhcl6IEFWtuEmavVsNC9G3DlTZC4/Af1hX90urHpmuIPvZhXvrT
jRZy5V+HIuLkyP+jxdmTO3BF52e4bQ0j1AgBFIsnS1mTSVvabNO0aIK1F6my4IAMKOxDusaGoDPM
fkt9/Uep+JMc4U/E41sLzMIy/NYEn5YzLlxnpX9kIls/2HNRc0SiOJYckxaPa9tv0pBtxIF4vsLc
uCeu6JuOWnfHQ39wT7rp1KDuDNneZ7G7ziqrUBTgaV52GuXsG0Nn4YsySnqa8oKSGDmz/9enQr+8
QcK8RB4tVtCflNGv2/5cKcJlaSGiWAvrC8TPaWGuRzyqsBXW2ULU96HSeo7hDUBrNQuY9Ex5c0Pv
THiYhfZNHWqgy5YqwtSK3p3YsoAIqABgrQVv5Swo8WVh4ob2JCPMKTPzEGeZCjAgKxtzUByFUsY4
qve239yeDv4mW1U/i/5w3Gkbk2D5lFX5oxqFNzF//2fq58X/I5jWdngwuOWGVzMjNAtlcjSRD6pR
5GMFk5KlfQZ5UtDZ1zS8CHm5H8GbCPNBq1+7XptXtNscyak+cGDMR83DFMuI8uQhVjb45lVr2Afj
Plg9WXbuLVJ4bnOUf7e+3SLs6VLWoQA7Y0MwOzpstYeUIXqV96ZkkZnWid9WMKlSCB0CfxjPW7xx
EZa8h1Zcdtq3rQIZyuk9FeoJeteQjgYof1mmDEF55RuBagEQWBcQoqQ70H9wb6ZDgAflTrZV8KH7
k/tPlNsEsmOf4BMEr5LGHAwGaTi9hpJg7eRr1pnrCVmO1tmPxVDjS7pQBKJaRqyxntry3qE0HnJm
DsObnPyktUS2GJuG6Z15JRJMaolyXrSRUZ3o5pR27SwEqVNI/HSYba4UH6bnokzfuSfJYxMMviTr
gxClBQPTlPFbHc3Uc0SBefB7RkdWgDXIWYI58p0GN2YdHXIfm8vLPVwLSIsMCWL19c25p9u8NWus
ZaVuoFNO8MtvzPwB64U5Mbym1rzswx568jeN3QyXWMEkksBC+GcdtA+S56Zn2VVRtzr3Y5D7IZcw
Icb8lXzT7LWwz5ZV4ucHhfj0n65deK364QUQZOH3nH5rWVwH+YxAcurhPHd4A1pWoS0RA8TLvgBK
7E5p/627y2RjrvlgFX4gEeQmwJ4zLuEWlprguft4N89F/Pdqjo/PacKx6ZgcZnOvXEvMprmAVpF9
DgaWGnz5bl5riMT/J7TljHMhFhBsTc+6aiKbkqzUQ1JIcmJ9NNlBk2YsZm744IeijWCQAGgxg3w3
9rV7YNpsltEhYNScumDlsAqWdJeBF2P7LqX1TbmVWerrOlNi+rZvI1xNT1KMmmm5mAXwDVqO5Fp8
D/4VaEdJRFDRzs0vgbkH0NS7reyiDBgVgsbN0SqICdZRzkRbg6Ru8srP8+nTdlvWtuVNMfN3D4oV
thXuItTbd8D5RvOA5z2oMc+A3YAsVmjvzdfKPjEynVPFfeumiFcJbqcP4BZ3cSXx1M5SzEi4xMOL
NDHERiG70M4689ax0wlo6lCD1MNOzVOBhk5ISVfu365rjyGW+m4SCh5Y2dY5bFmofORbusBUoJ2k
IsPSTQZ1Bdjpyj8BBWVU7c12iKalfC7AujqAfCIuSUlNIHVrf9o8Veot7ZvBe1z+XbIj67gLyAqY
21fzusbAGtOGMdr6YF7W0YqTb7JH7XZA6qpaLcDhF5xBsChlTIEikhSGL+bYVA9N1+hBy+pp4enQ
vwHbRJIZC//HHiOWiCBXk0B3+pYFduvFVsb2VowJlMhyJ18q/Xq0rLRvJZF/gmnJu51f7i8oyZyC
QoEY2bX+2uD/RUoVrFZuBnRrl8M7mYw/Cxf7FB/pKN01YlmQVCW+KRw86jo7ugC5tMzCBmJazQdY
st5uUnTQ4nveB4brE3z3pWqz3n9uCfobf/xLxiqcH4Yz3VNU8B4rnUMA6N9R7mE6sGpoCCFPm/+P
KmDXJrhKhu5GIX/cMNNnhWc2EuTIGMxgACJC88P3/mlAcsqASTlp3NW/VLbfCFCqTDKYQ1QPhWON
mG3JFvo/x0Ry8GwuknBJZVBJ9OQv3f+xnn+KWGBagwRPuiMRDoUDFloTl5WsODsy0XvjkGm4AK2W
hdo5THDWUFATNf9uAJ7SLHiJrvZuo5MNjQcAgZveBnPMi2uUCYofiyHkPkRJQO+fjux5vz9iLD1g
P6RhqpB2sGra9zHuw9V35T6APOwNsqubfvYWIojXNnDvkgKrkv+X34OwvbOvwf3W4JiEpwVlbF40
U0udoukoKz/Mr4dqvp5Wuc0g/Qyse0GO+p8iZMH1+v2XcGxUp3BI1R/a6jrg6HcIFvqbLAxYY1WO
f3K5atF0eHvQ4GyHZgfNLPceDNd0NrmBbeUaSt4QcFBFLw5n/BIsyeYZogUfFt1/qYIeceIGtF6k
ZfcYCSuFxaA/3r1Lf5vS1BVyOepB7elzeIMRr3h0OzHoJLL73cqj1pyH4sgZOv73ob2p6bfF7ezo
8jIAY+DpiQw783KpLIqpYFXou19jP3i+Evtctr9ERubhZaBQKHeFQnkFwNRxE7nkyFueW19IC4t+
BivqsaJJLfPr5JBt1Kvq67jDe3ujNPOdQ1yIHDMEWnR0n00iHktJ5bitK0K4OHKKH1XAcYhGhHo9
iIbdeRe4s/QXZa6E8jfTTiuNJ09urNZtR+A+7ntDLqLS0iANqKbwPg70nQNiA4jahJXRnHUMPj+H
EiEnXSGUP+raj/tnvlFbqiF+LCLmCNNMZeYM9Nv4vwFo0kkP6aIWvLr/fVN6Yn3aPNrhs4F45OJl
67Dih5XIBOafbceAXGTy/7I0ssuIYuBX478DeBf4kcpKvaLClhkiB/zg+/wy2BanMlwcthItLbKm
0+nnwPVmn91aiMlo5w0NaevoYyRG/HvCkAgfdDrgmIapwyL8VSqKnjCUPiE5pdxRUvI2zL52VpT6
W0oWcaHT5dW5MixUAVmkf0s5ZoG/uslfBYIl8sW2f95QYizusszz+WFzgntGvA5bWOkUU6+TX+Ea
Bo2OeUoJhotRZtFy8zvaz/zjIck4w6YGKbE0IKHyCvNoUg/64zwKnQDVgEXTC1Ly3w5itYuAAXYV
gxL5rbd38nm1MoRHGaZDCqE8VviQi1cwylR9ArrG+UDOA3ER/BjXhei09UMkneKN0I6sbT/kQDTw
BweijtuIaw5ZKbcQZdg+xe0Pc9EaN44M3tcOqPRMM+5jkahq+qWu5WFQxyfWduk6HRHPvvb03xSV
S8SF4awAtJjcakWQNegYE3q/CsHHE419QjxXdl87v1x6vPKRSzuuSHPkXIHntCERqi9p0hgB/b9Q
Cb1BoVfQOceA8M2QZh042kQxpEKDnXi6UqkDI2ef5IrhBZWf1O8kJim0gWK1eUSBHPyGtsoxnAuX
kJbNZKpnlHIDwsNQHohVDZIEZ3dhplJDfIdkuARHQM5QcW0QbNSMqNknwZzTfb0wadA0ct1d4OO1
4rEm6A0NkrWOUQM6BHZ3hnfxzP/K0oQVPRku3wSw4tW7bCfyOMCUZbARf42Dgvjw45lpU9NaEW3P
re7sevn+KrPABuBmgY99BJqDUhwV7MD8GdjsNe2uU/IHSa0ysEYUptFmcBO9eizjIvb7mBQ4ZzYd
O8Y9GXb2T8uG5dq6K/IVx3rQmVucJRiaHuumDb1pALoU0lv58C9NS4LczPk8nGckGWFlWyDUergj
NvJNIazfMsgHlMWZ67cpI4xCeCswb43eFdwvo1ApT61cJ2WfxPSHHz20msGTWRxQKjBTDuM4/rIL
zSN6euTrYFddhwbxZ7clb1/KkA1/YiaSDOh21eBwyM2KNaHO3yD3Yuj3If2knnhEzW2hYtuMK9LT
vpIiz2bbZF31XHpqOasXt93jKFMWLqLb/qeIKdygyGvP7cxdCUKmsYtkWQ7VkAIZZTCIJMFZXQdC
sedTTFqVL6Q7zsacTFdco6XCpGIRYga7W+QCr7uHt85KKzMcwaEAFp9cmtecCe/kEGpk0Vbvx6PY
jeswznCSe6rYi51nhMGqf5iS9OW4qKJYAdk0fX75zfJ5+RQ5o0WcCttfeBD490ZNOwvTeB+gh59P
yOXzRez7Viy8Y5J62xWer+mCMy9HMfxHoqiPIQRcKDL2PJ7LC4nUWXrdJTGJhQ1eeGxFXshzkFO8
yqy3MbR6cKjSjIJdnuRIxGyjPZLFqkJfUnxr72LYDYT1E7KLJTgIZ9hgFfzbasAcWQhV0eKM/AkK
ZyE7Kf37trZDaFLoJ6vR3vkIppmJ1ZuK1FFop0HMMEUk+iDBgF+aCwq75XNb9gTQkHtucX4J6gKT
TSnYLwIggAVsh3QMf7iJPrtpNrIoqvv5ipWuSA8q2GIw9+IXPB3lkeutPuJh5WtBwOKnS3ykoSit
B/hMgvAMB09/VH2OVnwSzH5FKN/sK6ZjwHxY6zL2xga/MbzSiDRM1b8kPIfLBmak/RYkA/htJ6ED
Ks6Ju0vJLWhUjkljGRTUWZp9zo+cWzoTf9oKhzkDHsTMKNBfuDff5UlFQny4sXf1g0ENt5lqvqvn
/YnS7s5wo3Rkc43gquHSDrwpgMqqzCEj3MtPhFacUvB8ee5AIOiLNsqTFgHpz6oxXSbcgnMINh4E
kdglh6JQp89W+Rv/NdSeu8yu6jBYuoAoro9L6xJ72srxJJ1ZZLFPKXmryhKqHBqHcUdy5VKt3ujB
WjCmVgcCc6Of0kE7jnwyHJjXuTI66S5SBAmkdRpWsZz/SHeOn0gPfYqWa4B94E+GY+sd/UBoRMy6
ocQjC6/NzBxJIMWKMvgLH+4Bo89JbHMSj57ykrmDMnIPiBP4gYl2HMyetuX6raUrUDOq3nL8judm
ghcDEEcgo+eWG5ftNdTfQuw9+mrtMX2bCeG2etqX5VKd++2myTezSWIyAQhqzBL2hLsvEDnScjLn
8DlKjXElqf3xA+iS3NpwbtHHvAHjQMKzI1acf3/jXjUKrAHxuMBLmQXYUYXtUWherN+wPD2FxuCy
JlojVnJK94ZLNBtXVo8O4OfRFQQox8f4bsMwoIVWujSMsQcOhxmCtT4SWm7aWFBpE6KsL8wRi2Ss
FFR0Ae676NzD5X5q1rQP6qOVP5bXPXIb7+ugmedgmmZW9Z6BBnFAJ8t9eGm9COgddM4vVVR406tU
MUSWz+TGA0Rf9yTejPMeNajOVG8DNMyDhk4Ih1yx2Sz7Dm/Bl1Rjw44aXVwGkvF3VIL1VjyjFIWH
MyAAnyUbveUvo4XvfiGUvXn/vjJtW7RBWxLqbDE+A5KXsuGpUe3bM0ElrNRWIAJEj3HCYzrl2jIT
Ccaz2FLK6lDRLveNvn0+5twMEujlKuV/cfYo80g+9nieNsKiQ7xvqamVPckgaL8aTijnYBgn0FMh
1ZDWli/0luRyr3iy2exSKbZGWtA05CqsyXEC6ynQyeGp5xRyDrbji5ebl9VkopmpMt4GShsXirjf
sI2KzBz90LTLcWhB6YjDET9BRCRfbCquPTBBVmX7LZFxPwZn/Eqe4y9JFW1W+42PdCaCxK02rkZL
uZi0R3mCIM1IcBhM4HdZrgYKlnI0FXf3RoFUNq8AlFPiRfrk1DzGZite7L/iwY5LlFHMeMFInhf6
ah2yLG8jMwycDN8PsdqV1fm4ciGrR25NI9V0xVU0kV3cYJbOQuWZgBQ1uwKvz3QbRO6WrHLIsa36
wn6HgMMDKZJMbQHkteDcOLs0De3Z1vJeE2b4fWDMUCw4/wu9B737A6KZxBO92BGJmkpyOHIkU+qC
4DUdzT3WUEN45/fTuYRJU9Ya6eJyXGdWl7A79qLn9VKszf78EbC7FOsyO+xlVbg6Uz/I3kc5YGJH
q+dDPvzFZAbisjt2pewepZhBCLDUCb4OIKpMMCjpcu/DAAsA2rhNVxhZiJnqAQAPBuHSF29GmJu6
lqjqSrvKoDEdqR9siMVBr/nFPw927KdC5J/rDc/ZlubC/Q1H1wqTowpbBTN/V/oPkcB7OiM6iIja
89WhHiYYhTUYtM4MyrG9PbY4Sipe7Sb4Fwi/DqNkwpu6zltroBTfY02XgQbLgnkMhR9EDhKQll3W
liDIyc14YynUY1XONROB53Najiiz2nIgpqzgR8xVR+Z7IjJhTd6ISqjvyRCciPHz3bp7fhzg/I1l
HJ+4ihW2C5stuT466LVzmtCWpbdvcyMH6QPnkSTFiVg475HGBbqJV+nVSFFNF7zsjdDmMrA8eNHX
Agz97FW6l3Pud2t9xibOdQATpUrdGjdtfengV0t2wHrFBfOhboCypfjNCak80UjyjvZJds8qujd8
w41sMSfACHYf+vUxgkiZbJONPdCs30ItttskkhM4i3BOIr3FykMTrN2tRnmasYfTBoaYXQMZ9Zxi
4Rfxu490E5iHIWhmpjmjAFA9ANDQB789wW82zrCzMCn6L/R4ZIa89jkzFtT87hsO5gW/1aRi9v8c
Z73QCZ/kBo8nIIBIjCMC9zgcJ8RF84tuchH0jVM+FxNeUjYwX8vs8dmpL8UHHj1aOv8OiQVb1BNe
oGb3LjYFz1l0v/NHOoRkusmwxMs3aDeA2ml5PWf99NQj73FXEQ3tz6Quq4u512d0pL22L7aZJnHZ
dJrQmuly1CpPB2V6BLSI/Ptk+XMPji0cnoaDU1FbxwtgPR0DM6ckh490OP4daCSqQTFUfa+q2tCT
MbswAQCJqjdOG0G5DLp95Mn0GeGUcDV1XL6TR8m4kKgfCaE/V4VxEaL5MdPLtOffpmIVV8S44C6J
yOs5d+puVAoHtPIHqYRuxwHkOjGq+ybwVG4nY8YmyfVEagiJNIBgPzt1g0LrJUs5E+P8yjVIvGk0
4ujJy1S03j3B+vsdJrCKrrwJ0xcP1DX+9MfqTEGQEw0Ys2KOigYptOvmX2qs4Ew9a/pRPW+qJ18X
y3PTGvcCj1I+BltcXsRsrr4WjGJvKQf/1NnTOK4qR2yAcrfPXmlx7+TPITN7w11nbMWLZqkGoXKV
oBlI2oIp5/5aEHD5B32W1N9BIzgtznCwyVhL8qWLcnbsfkC3lSAUdDjxzmHtWb8Rx8c82Pa1Ai7P
W0PMfiRU9h65bOE/GYvrh14wICB4BEFOs/nJX69jSK9pXvqibm64Ic117oS2NcSWml1iVJ+PO8+h
0kQ/SvriMG+70vx550TvODGKwrVKiWKT9Sqo7DrkWV0CekSC2OOKqEkEO/W1mWCYt6SXUMyAcE6h
Xl9zoKF6t4SRcWOL6yvq/8o6u2Us6aS8uj4yvhgYtHDCTtc2ITI/yHatHW3XZuBkYWVHZbMRiON3
EViNdRC57vj5DBKoGBju+I7O1tXnkvc/5wXZ81CLtN6ouN6CH2yNYkCeYNYFBE8fgVWJ11OD6tsn
QjuraTm9c5TJJN33ElFqeDsLkDlX21hMeIvlkq97MB6aekrlLSyT5IXO125R+iEZX68bFxXxWJ+A
kjnythbH6G7nD0Ki0Yzhi5tFVPEEZRC6LH71Vbg7IGTXutHcf2JVy4+zpeCSsKvTT2YUp6P/tVup
8aMkINAAqCPClVpJRPu2KVFqCWAnitQfUm6afpOQ0kjS5o36znjWP5PrtCT3QOs+gl4aAgO3lqJR
FGtpLc9xbYtULG5JM8kSLK4/9fhjCLew2lmkIFAOQZYnGHChU5QdbAwyi8QtWdMD0iitgC8w/pkC
byzXiu2l4pl72HKUkdUGpm8KVJBIBXWd4xJY33IB6JGMJNgutx0rh+Rw0lizPgDkniPqf2VEI+Z6
OCV8OOkKGomOEdZ2YqFkyofyJISO97wKbSiSqmFJTDQ9ZREVKBOXdY4jmLtMnOBnYNEZXOXh+yQD
2kuBIeVbT9pXtrq+g0UiyRt67BRpbm9kYthZm7Zk/8AAEZkppnu6PDW3GhT2aUIaod1HJ3M7WnNO
D0wXHguMM8Xu9tsFvdBTYdwwDD0y4bwhbLiPq01XXpRSstv4NIXTHVUMrhdwG89byTpAEvYXqpOG
PkTYQFPYmJ1+9xJCs/sZksjbtc9VUEUcsPuLdV25xy5t1gelk/z/JbWtIH2VYVyBFvxFJ5HT6et7
mJDmdc+ExY/hQW50D6rnizF4ZxCs++xRjrpWJmr5e+6lyhyK0eGOaH8k6JxzNVMM/DoxU0hqf9+K
DMYfz/Rk5yEAxtHUhaQWy0aOxH3abs11544hfOI0FVQpwznPpjtmeyrq7gxzUHhtzsc3vhAAuNXT
1bRyC3ASv1XT22DWZHoCBpxQ3CSEbm5rI9vspPRvEASAFv2B31ZrdxZcq9RvDlXer4hZUnuu6wDI
I7pNa/+qQntf0m0X70DX//QNzOZwcNdHRfKC6+xBnXeMm/TUxjD5ciT1HzXSwhX4NjamMRVJ4Hyu
oP0+/sixEsL2povPHXeTrypZsGSbaoB00J/H6nBecUArCshVa5ffhJCajHTrdoJ0fBukeaNawamw
ZDp0t2J+n80VlRaF1t5okeEJMejcVZs8ms+XtWENu/ZE3ltKDaOXsSKODn4jzsvZ7ZuwQSw3ZDiJ
LMIZQR8WlNEw1nlQJS+rQz/7aU+uwEOMqYAnJG0ECruVXA8dZZoLm3kT0x2zlVagMEcWWlCWnxRs
rfG0IN5xC19zo2aVCSa65nMMc/XMKkGIZXW0Yk4gt9y5/YJPTsu1GnQXdTe5grbCWhijaXYp10WH
YEyhbRaxLcv7Hgi5igPINOer5ow/PGL6x8Hu19z/VjppyLFe0YRRq/NRCWIawtd1wSCMJY13o5G4
SVekC1OD/pXjHG8UVT1UZJFkKVp8ErMRhHb5y2zh2Glcr6fDFBMh3CFaWqLcXABRTeZzJrsb764T
HABYkxliPyAp/sr8xupsgkZ13sDd7crB52NljDcU36kGRETlLHikSh4/CYWlfvslNO9NWY79D2QR
wGKTurprCA1kHYww9OGWjAz76DijJJ7GRnEgStSY3mkHS9rmD0XEGlOlXFyMZi1/e52rWv13qiEc
JlqpONBj0EplotdlhXTKpJYqB9guZMFY7fDGIempClxFEmRqvtjOWrepaNTFaAvyvaNs/3E3R43x
cgn6D1KFjYhvuMXqnMfEKCLd7DgU6r14KRID5FLaJmy75IIiPB/4u2tVEtW7eu2spgKeXFx60lHQ
5lJCYrkqREbieMHTy81Iqtjoyvby8xvTHoylHfm4NxZKBzUnLdSKClVor+l8r35DreBd3/bXHl20
s8iNxTEBz0i++e1HiUxYoYgY6Lyf3kHmZx0xplTmtJmEqh+0WkIRRTJFuGAN2n4rmj9wh1HLGdpY
ULpxztMjBBLv2ZWlCuwE3xFp7pdMfbQVz0bogx2g0rFmesy8Sxhe9/WglausxhoIN6iHHUXzW2Ix
vsgZYvH7URjRlCT3s6jDnV5VxCqLsL1hkei6g/mgx8eG9r5/7KkOlYB42yBcs+clx74AzDAFOH8q
MfI3qKnVoU0UDC1h6pCoOTKLOz8taLuJWziEqlAoVoHHOROaduvWLeygte3jHxV9JWXuaHCWgE5i
HWHUQwOCzQLDxtUeyq5ES/t0ZmV04C2iDn/e6+y9gZ1TClJEIGptN0sbCq9Zm4ust1pukwyMB4n0
QY//HbNaDY6LTk6m077fC6pD3o8TODUsIddhvZT+8bQwXqdjHphdEKcy63nMnBWYHu/WWyauHqi+
eM58VFFgDsM32XQx4uCA/Qn+Jf6n4bKTZo1AnPMGiamMscuMgWspnF2rsvOWrTEUK0MUqDrHjZy4
9K1NFz6JwTvUkKqjpuNGN+0BcZMDie+h8YZZjPsseTNvVdebFJDoGL5a9fqF56h7k5ESCGTl7I6Y
4XDQ99GYAmdFhCNxbVM4pxgNyWdiRbawVzABYfa1Qe0tEVijs5TJ0MW6TriWFHdseW+ZtRmFr4QE
6sPdAoNvB38b/neZGE0oMQj9t2vTxWt//n80NS7cswMD4uQVZgvZneFc9ERriSftc0i10/CCHAOd
5uocsHf5gSYhm/TyM4sLL8lc/jBLaYIclELeSBs49BFJFqyPwSmUKk64xwsQOKQ5ErYEAgdJE1Vm
MCgx7Wvu3HXO6qed802Thc8SjrB2q0Lb3Lcjq4IsMEgs9XQfJPPSNVM7PZYTjoSvUd9Jqb2AMLrT
T8H3U+N9p4QbHSvuXNg0UHG0XcxUnvf731htEFUT8y2V3nYjnKa1JEByHew165MAwAk6BLoY619z
vi9Ygm1XnUhjqky9T3jxd/jXofmPwCXNVEV2unBUezvobuyrv8b3bIRa5Ja1E4ElfPfTO5ufnXdX
khrKWOYFIlCVhH8tGpyqSTXXGO+9FaSyxfdG8Wgy3UrCog5h92UhbPJtM0h0cD1fiUtAx4EnCPSy
9VD4kIpGoVNePju6+8fwqgTfeVN3q5K5T8zus/dFI9k1VKZzRztOEuVhJehF1OqXX+iMgIINuP1l
bpa4M4ylbXvO8rYgqA8f6Rf3iJsOvIGTlR5hRRSwD20jeZXSDjYwXh/zWDeSRKtaxvCiFJzlrB9V
jW27OYQiPNl7ADA/9mKx1WZA49rdcGgOjMQcTaRIXLeihJuGPcqmz+/vvlxQsuk6QUBFzULu0LnU
2/4rblur94vZI88yyhAjhCSCzBx9N3Cbnf+jagqb/wU/4zxnhYjuNz4CP6/0mugC6vgP8atE2ehw
3qWwx5+qvFophgWEDYb9nE0kx+P30UXytApQZdq2dBEr10nDHbS1EVLPQaEN7rlJZpkzZJga6j7+
K98ii9VxSZkO7ug9oav0cAIS6t+8vluBPJ3MbLKshgAJI/q0gOMypTjlpsksUoiKSIhUcbFUjei7
PT9HItoE30KQ+y+LnPNd9WWPGv+pcy3THtlsSLJ7f5JXSsQA0owdUua/td772ISzEO5So6pT7IYy
CBmSBiJ8qbf293OPQu4L4h0wBSjSdxKykPVtUOczyn39jSOsZkIrHbaBYSreiT1zErVf8Z8ZpLmH
o29ucbjls20WxwQIg54iy5LQYR4xuZCZCq5PSDLSFkDqw0xOp/HEE98sR6Qx48OpduobkHMCJeU/
6HCcVM43DRckVtZlpEjJrUgy9BK8QmfBCKws3y7LyzpZWxPLWbcMc0IucDSOorGTVyWst4EpO3Ny
oj3Cdb7zvfdJ6y4gEbm3Smro1/DjNJzm1aFrpBvgMitvRg3OrRnZWy0mPJG2j9jqnlehiKskY70H
v3ZHHFUllPkW8wMhES5zRPWkwPGlWypPCCSmShu1sSeUxd64na0/fN30J8Y+qh+4qDL3Sn/80Sam
0/UG2W/kXIFGDX7TS5s5saUw2Xd+YjkN7mVhMCvMGIrVeTROaCb/XEarUqS424ZIzwE6on/v772N
RCXBo65Lf53XdID/lxd+h0s61OSXYR1r7W4llpEcwYldoC2AydedfYA5mkurUepGz+UWy7RaHNxU
JOAbbwepebcY5O/UvgWRHyH4pNJ+6KQEq4sGNJ5X0cMgfam3W1l5nGXmeB82UrNNyvxdTJD4Rzm7
DlLo808sKHV3mpTmFkFCPGFA9D4s4EONKq/n4DbfagQwuQHT12+t8VJxL6Wy0Onhsc5Clw+n+iSO
yWPt6P2nE2z/MOTjY7ca7ONyfA09shn/xXJ73DiVk9Ibs7dZwfgTWaZOxG9dDMlVRzKYWPsqHfMM
1pBp38jmQan8zPuFrTjM4dL0wAEqTonW5a/LUcBdVRcjyxEq8d1yeO69LRy+4ybSJ/LhbQPU1QoB
E9sc+gJPbLIQKI62+/9orc03DamK9N6ezcHdLwBKI72HUeGdlXtMGGtZ4Cpy/K2J9OaI+oecNAaX
5xfeOh3wr8E29NIrlamsUON5aIi9iJrCiQVQRqryAUYy4io8nq8qYwq3j8u1JgteVFCITbMvWv3+
/6Ydr48Yyjyf5SC/ZwKricX5xTgA6oTRxWA8ndAAZEdSCukGFjAePOTK+IaFNUkrZVng3cJ85hI7
2xPIHBBKkbpV8fYNULCMH/QGToZNMoJOCavw5VzQFH/9xrm4jXlKysrcQJ5aNsV7KAst7bwUyk7G
bLhY6/TpTUF+VR9J9lqBimtzNBP7Gh5fWpKr4r4ibn53WVOawsh/hTHIMu/2keO1C0i/ANz9SzEI
xdJ5iQy7/dFmNTOe4+SEumZsmde0Yh48EEzWR+sG2SjW0oLiSZed0ZDxbz+kJPIlqt4+EJ89lioN
UmVk+P5zGELY/kKAXbudmUrx3nLQ9QD3fqTjVMu/MWMeaC6S4QwAlEVKfTgFci44UG0fXFSSdrWc
O+g/YqyWnpACeTFqENuhsYrCRoisCkdmLXki0KW7gqOlehBFd4V4OMThgBIbbujehCSPEybynSBx
sVybSQ8rTo/IzL9Wj+UXU5C9O0NXC2AgqlbPXibYMmCXWfuVr9CZq+ZfVKHVtS5gX5+VjB2NBRkm
Tmkg0TDFsRVhxkVAIVAYsCWYhN7qdwxdFIAxCxqrn6Lk+fkr9FJu4AS2FJRbgOP2YfYVoEJXTkgh
l8XMZDHwIMSQHcM8Z02qFKjxhnyPNgEpwDkuSCHv+Xk6aKqztmhMYbR1ZcHDkXRlp3s7Mojt651d
rfMYiu331wpv1TF0sOmHnChm+gmUEjrwhu8ksKiHrlyP90jfXHivIptw4cyZdnTDJZEIN18BhtcZ
F1DCf5VvDPUK0lER1DSEa0gpwHmxo4wUPyozifLuz6/RwsK/vYGaM9HWvts93WYpiXfE6Ura7vjq
KLpMfclyiIqLYRVGJ3zOXfu95o8XQBEGt+jOofcRZU3YUOLkT8vhaV4/YVKo+61BU5DNMyH2pF0h
TDiuwTcRHKRb00TWupwgOHOWv1cBx5QagLlO5qAoSy9ECVnSeU9QlMW5YuDAPPS6B/JlqKWjRQsq
Ja3Fl7K7JVyDB/U4WMVuOG3ccbvn164BeMtee4pe6hhCmnhLCW2QqGIXDQ/1aZV9gaqADoCF8QYy
9xyrn2oA1sadwQ+laQXEKDs99Sq+MSXXLF0Slg85vKlnlJ30W0hNyLG7rchofkKsU4yxuSYHatQG
j4HBf8dc5PGfJanCCKIrhRrJPlhsr7mFwY+iMfbjVNeX0ZQnRWoiBesqUIcVZy3z62aBwOXXJgcZ
lHVk41nfYAsGSnSPReuveHIH67inAzUO8uH6dTs5vz3kQvcrs5yZB6SMc7sFUSXXKI+yzQjTW0Gl
RfMHgNQ164vdEIp/rqY677omQ4JcabPTqDHC2HewHKuWsoWUVriGI8ZUJuQ83dq55lPQH3AB7dgk
lMs45P3zOwd1hWVMzEaQkHjBqFBTI81P12UnFd+lY7LHApCtSlFFj6AjdEbT5na7LHQF00H2BptG
6gHDQSF2QdRhwNnE6Ahbc5+GumGxBHwYSx+I3cx8pnGIjAfJzX2U48fEt0oNdr+/mPt1MZi2s4Bi
IAHcZhgdT/xbIDHrv7ubZnxkjb6hOmTiZIDBKNQ69nkT8IQe+hI9ZJw8TPFyWcl0VrPIR6dOgChP
Jxc4DKA2RMpxDr9h4n0lI6g5hc0sCHq/RN8hTfKuJfX0JXroCtZSl+eWP8BOkkeJwS/liz6Nt3IJ
QeqlAb57AsjxlwJh0efzwioDDwhNkTa5711W9T+HcgEf5gIRbKZ2G/6Mq+6RVkISvlOA/f1fj/xq
klq2x2NoEWcN3LWlx0NqNCcK4jJj4quacYcMEjefu61IEXtNtkPWrWscPEgdSY5OAviaxAgDwzkn
aJfhh6gmEQoZ+ZESL/Hv2TghXa9t/WOIpdV1lrniN6PEsYOKJS2FlBtWTTDJpoMM1jWpr4HY0Y/+
JEzr6TqMdk6CDjY1qU3ZqnMdgq6wzdDVZacNiXDQIKBUTxei9wVZkbN6sr5m+uzNpCLfkhOXfnBz
4fzmIvZiUxdwI/4pydnwOMncbgzDrzNKk05plTWWo3iMIbBtQL4jpXBXvP70p6No1lGMWrm3Oi7u
L1W6fj4CkfJ8KGVdZuRFyrZu+yK+fXa+ysefCBItna/SnjQH9VehM1xrPXxDHkZUNaHOtL08O0uw
jqKuZ1DUymOry+D6il2pilKiTdKSiJWRR++Zqg7dr0KVOAUxcL+uZmb4LENuRNGA+1G/dIIbhdZC
lSvlI2xWdOLTUSS4wPPnd8KfS516WqfIYQhMLtZA4tIomkjh10rBs6OqvUkUhWMprVCz6dVOvKBu
8RxsRTqn29uZRNzTJHoCzHqQgbmDuEIX+1WhIeOdQOWDekBkEqREOUSNZp6G0hxQ1uml2dm6hgMd
Y2epNG4JUZ5BpQDqDhUgCNI4czZZaMLsqWVShQTToSHw+Z8KF+hF2bhMat9kyg58MZ56335sCT4f
2kvxWTXNVHU11JQ6JR54iYo45MVRlXg0VVOySfl96Mb+/dX3GC8BNiqZRXxlCojw6RESiowbdR15
JPswf7qDuohug0vHbnx3vsm0tP5B0qQLGvHAXF58RoflHFoUdS3Y/Fiy2JVP/pJSnlyYhVZSlLXE
N6UhXr1xWehq2AvRt89FI9uzaovGguvwsJBS0/0/jNLBY0FTAKGMZ+iM3befB/i9NffMeagtuzfe
z0eW3mwHBDkKELu1wJT9C79idIUknMKeYqIUa2cG4Qgj9w2kOzPm7nxdBCFFVVnvcbS2XQKh0kOE
C3iqLcLc91ZS7BFxZagwl5GnPQv2G4rCgy8VJC7ibpApe1GbWjkvtOjUXx8gAzvF2NULk1VNELgj
29xCIw+Zud7yBv58T7QbxJ+Xxo+aFmre0/8dsketVgT+e2IZTvJ9BlTVXVgqqHwIAmJ+qXaYcTaA
Z4NcslMwfQrKuMllX1WwfKBtrNgr7KKJ7AU4edSgAnHacEYHLaV8Y9ts78ecGkchd6DtqF4iQhq7
Uhud+Bg4qZGtuvwl8O3fWBZ6cd+ky3zMaMT8Qp3KAxX4Y0XjBPfmqFnPxOvqj9iayrJIwIqqals6
XT4bs8qCW36PJz3fF9g1sMMN4DtjOH47weTSQPtycvRX5lWd1HLx8fNxP4ZNEoMdB2FPiplsAbWF
Y/R2Kuf+rncn7XUedq/9lVCwF/WFBg9C+0ch5cxCV5w0ThdBkV3cUNOghnmLfMkEKakk3PaiOLZh
QKESirpHvabWj6AhQfKxSSz72MXrEAdRhmJN3mLovd4Gh/6px412U4v1qOj3GHpT2nVd4EM07dcc
toNe7qVXqWA6Dr0SBf8Co9DXcrWI3yOSvi9GEgcKH/5DgTZghA5IM87rYXNfru6Du7B+I6FLnMJh
FEh/4GdZWz8rxHQ+LaiG2iy3JMMnVTn9DqfGtk2WyXNloq5mM2NpPQWBTSm0IN2DQxMAUcpQmSEV
qEBb0vJxyh//uEOWtz0+J4qCKpQtGD01kwggwqym7gqGlaEuqHf7pkiYb6ZQ2mXgydzfizQt2HsY
2oZKXNsGKLb+JOTdIALbCnwrFHCb5tUHYiMutvfQtvGbo77ybfq7VRtH4AZ0tuANr0N2GYvDGQe8
nhu4tATbJaPPT8aXBu8+VMCNhF7hJvJu43vVyfiquQK5brS0HBZw2IJZ3OPwjphGueksPnqlKMv7
+OQfKjXGVfRERGMelWrOfaaVbfXmlgpun6WkpGWZLaeKiK/9Vrhb25LAbrjENXc7uGOCD15g5Cn9
mb49w7onEkfzQo1oLDGHUflxbpVHmi1ue7EVxnCRxrV7IMjsELks9y6d9vVpYkqOM2gIXqSTtiNJ
umgC5l04EPbWf0+UH3ETtVFLbxF+X7xG0GROTmSEibsfO/1N3FkjjcyD9byR2+FUdDt8k5n5FAef
8QogrolkI3V9HHw6VwO0UXq0z1oawhnV1Z0roAZ3aGIqnsnBs/njIod7tlpF9VKIPa0nFdrUYfov
ZOkRwUkS35LeE5nbvYWdKIhpeK6RInKBErRCNksZZQRIHqWhrF2Nwec0v/W8sq6bLvzxXayd8sKQ
FbGktyB/sSGeBvABJ8hMC38B9c6nLbiLoyX4rh2mxp63LMWIXCKXh6rC1AWaoaJFb6o4WTID2JS0
W6Dn+sDLCiozocpKYNyUiLuWDdqYDEkZaBVXjbTV/MJdCM2/oXzcx9ZfZWI8KRBbLT7W7P0rw+D6
ZRz8w+MjzfSnzcfeoRp9gFLtwUlC+QeK48EgS0B2T961Obrll9T/B1iODS4JHMywo05PBX30p8S5
xpd178YvYCdkItW5V13jdEoJ3WGD2spXBollCOJEz7QBLd/oGzL89abMNi88SVxmMDMjMGlRsBUt
zROCrE8oaj8PALUdCU/6UgsBeFxBexd89AouHOLHveO1XKHN65SO/TOKT9YEW/f2zZ0yo0e/AkiY
gGLmCMjeXCvhTijMjn9/3xBPUPiH37JtyylASB+qFasvCOgWFEwHQYiEbohn5C6U2NMFYuVCc+re
kXmljFd9Dy/xAM2tzNn4ROWJo7gTT3ySwC2FCfGGS4uqy4O+cmSf8ITOs6RPvIfoi01l7OYqgMB6
Nll/YhvQE7i22kXBnZhrBu8ZzfzEnIzntWmDPIwHbieeR8pCBFPncvV2o+BCYBoRKREW2GXXr3PS
0i92jAh+b4zK4bRHzcwXGWM5PTYi/CB7kRIrlxvpVYMVUg8+lXAan7wbGs6Pb7b2niH1d0LGBpLB
m4F/HvEFljFGI+xMEOj5QykaUB3bkrqjyMDNa9f+lQpI54Vgzje9yQoj9pWdYgUQsNlzhZdJpLCN
6ajcqhm/2go0murafD8csVCxk0Q/v7OXjgkqOZK0GeclAuhNfntkrwfUOPsNhQF8jRee63uwoomr
mZyUc40ciSHUODF+Ktz86Gyz6zipSBw1jrfsLzaUbbUgieHAxkin9n2haqzqcYONBs7SkaXFAvXz
YdMZDTyPV3kfhsyxaPBgvPF0c+mPBnWS2/apPNv2+anbwfujqngdxH1JCTpBCPbBA/dlPncQrRV/
jnPrKtZRdHY7gdnF+C6/tXExtVKIVe6A9vXdmZ7AOMu+IGcRTK/Xe0Gm7hv7dnF5FDtsH3nr+cx8
ulX3SavX+GPhrrpnVsQjbCGwdws5WTkLVwLOXdg3dXzXmqS5wbhO3xiG9Xa3PVxj8WqceAa0Af4y
3mQvc1hwX43kSAjk06N6UqMfT82+4qhIrkrR65Aikvm0vgyg5Q/i8PcnNntkx3zlDYz2AsWFvPCt
JefSHVzK/KiVZfnYcUtUzxTWEM3XdeW1qZ69f0LeAAVmYWjJvxb3CKIl6o220ccSTSuRiFQy3l4t
s12heWvM2vW9Iy1RRncOYtxSh0tbObbsjwJ/hj0MI9TmLe9WlUFqKBwPDSWoedf2tYlWQhCbcsr7
4+W0WeKq8X5uzI9gwyV+R+cwtr6NxUzrBHnGBC+O0aStAi3p5TnLZ5mr8zWYvj4lBkvQsiT3f0Px
FzcMeZOHj77whnemfaAEKP8/QZLxAFfYKyS3jzXBMUBDEE4Waf3v3CcoKgjpqtY2gQEH7I62UFbp
8CkGH0bZl420F2JDjMxdocdEypYgwdKoNRaza7esdZL8nLNDzGuMk7ilXYVdrnFQr9VliyEO5+IZ
zh3CC9Cq0W9XBq9A/CbQD+GagBDOn4/YEnkR9F1lF2uXrpYM2odMZejtTolNwf4YmzkoM7TmZbUM
chDLakRQZwaW9uTE64NUtijFzqXxgp3k7QmOkkkFsWMen8sTyE94SdAcS9urw/P87V6nuXdtseTe
tsIIUoXkUM7V8GJIK/b1EHXMqhTHMJ1GmKBYjciBiNTHwKqPUYnv5tEEWcsGvAukwOwAItwLMwp4
XlktBNtgjJLiE4Qq9TJ8mg+YxPG3/vJz8S/hfoiKS+skIt5VQGstX245GmG/G6pve1kSCB+QS2IY
VGrlBmQffk2IWDCWN2xOe1ewwScUjW4l4zC46hnaTmeT0jwEJ/oirMbKyxCuY5yus8kNT2j4ea3X
If3GH5JWwsFvTjB++w8Ge4V2sVf99R9Sy8TpdT5rCEz5EIjA/h6ll2uCI2mcQu0Pnpp4PcWt4L37
DxWxMOUIc0dFOGbYHiFH5HCZe8wy2h2Sl97HxlZosKWDliGPLIOQenKVMMxte3WGl7eMX5BaWTiO
r2KGgoeVQNNLtiKgPSm3+Mfe5K0ZIuZtdc/hrAJnRFMuWgl7L5+U0R8Y8uEkjOBmCEW5a229BVY2
YVuMTslp9g8TEBsOjCdyrs7f8qu5Xt+3pdmtMNX7fKbwTmQTXKNwyME60JymLobB43EDIR8oL5yz
YjeEKlCfH5jaTSBnFCDEwb33Ft7XreukW+i499cqpjzCKL6QBcByFWWHdQDIZW3LY4XZoo5cN0dn
iO/CfulkDp/9cfRObLZ4KAIi889IJjqrtVCmIqsg7gw2zG4mcYSOxa29VlXv948XM06dAyJnuEIe
ig0tBOlW9ZbYq9uZ++gJmgUvGyvPBdw9Lbthj+MWxXfPEgGmYynNZguwl9DekcpwjcL3txrsTMlF
tCjAUk8UWQNoNGwhzIZ5j0a1g86K+PrjWeehGl4BdK866mz+L9y58ceUS1eBcRZXMvoSUEVL4u06
O2Uc3gSlfqUpxx+C3/BiwhSfotQ6WE3oWOijNwuqfIgXlTDVY+kVtWLIjJpeaGS3zDqGHl3xEugt
9gaXB9YsQTsrkAyX0DRzztK6keo7KcgG6ZzBbSY2xtMOPsErCskcB8PKIqBBeCkIWPODIKcOER3u
4gukq5pvdBWpeyCztzzpNDyUaXL+SuK92A0xqrVfWmE8ryoLeq4EmNIEemF33sjHTS3un2Vj0rrC
upwx327AU6EdNU4Y9khh4u456w7dtqgfbMLDsj4I10FKXmqVvN6aKeoZNiVpZtwl1eJW+Zuxlsj0
0V5TuaXTWe2FjBeUftUhOR/3LL0tsu1TiFmn1fhVQ9WdVE7b3caU9uvTMYs1WNSj61xzRyPrAkdj
LOD+8m4vwpPVhhAUZWx3R5pnSCuDBuXlR98q0016//TieOPrxCUu6T8Ryv1WB3VNkhfhroQMNP1K
s6am/GwVlW6hjQ7NKgwwMVeCsfWodhbNCzYz4lta07i/Kb01FLXMS68/sgy3t6eJ+ORRslES9Q4e
DpKhLFNHK8u1qTWNarWR0GGCILTOfoS7qXBDysIkFHSQwxFGme9e4AWgQzw1YWzQBvD3KPjJeXgn
NuNfeerS7lM4RF4NcLB+zXNKxRoX9d8RAI4LGTWj4+dmhqcPVImEaMUj6ybTx3/jSdRUUX6DueJq
6LbHE/I8SWAJw7PiEBJ3U8Ty7vU0sZaPvx1jud8tj3LiJV78y0LesqwnJGClhe96S90CBYm3WO6w
ivXVaYLuUQdQKwFou0GWb4bBKadw9P9M9ylCbKEZ4MgS604cD6XjIKG/srIzoWhkNb1qgXkRFX8R
BzUcfmOfeuaNBMY9z+MdL0/8q1yrZO9VudC5QyZ+At31u5+K2rc96KzrpxoN8QG9nwSMPqDF4FVa
iT00SgAIkhcz0SZyijxBXB+KqresvN4ZPbjtgFiD0e/x6z55NNHhqmEccI8YS6U4jNB0R9NQ309n
V3iAOH9vw0etV6MPMG/0Qd5dxRM1Ty6ZCDWQGkGdYsq7slwwK/B8F+z4GmyYoghR/RmNyEuIRQik
faGrLzmJtWab2nc5a9hy4b0AGQn0yfJI+N0J/QxHfhAyvsO3onY0ZWMgh0Z+qIPWpukgqgdHU1o/
VKBHLwgP1lLlk2fizXMXDuKfp0HcGmTafYb3S0CjxHTgHw/uDvwXTzBiMronc7YGrp61ULCXVxVM
z1SWCZnSUXigA3zBEmfEdUbjV/w5uGGpyeu5Ev4vYWiTAygjs13TrPT30LkMZEggq+BpUfq1qGoC
hEvIf+VC0ZewQvcCHGwWeTuTkL7iAW3aWiUD+OBqkuTdUS+N3L3fItxmRxWqenTR/xvQiEr8HhEp
YVykub6Lv4wCdrtFOFlV/Nb/wx2pFzWv/vDilIktd9ZFTTj6EBCoGhatm6LqPsDbh4PtYdq/p4QT
q2GZPPjCF9SeA28lNOHT22Mpb17b4ddGy1UCHVH8uPtP/QmjaqvIE+Mi0+ItPfBolSOc1PPBDaX4
gFP6G2s7q43hrnEOmVrcJ8HW0lUcCV1vBAkpzgy1zjqxBmXj6ISLmCXYo/5bYnSs7tCewZSzLBt6
8QzIm32rEahfwtyPmOdghDfto4XlfQk34UPIK3xssGpGnqtio3L4P2ztv/MJJMI2JtdOLaAX/2K7
NfwwIIWpZHLuzgZFCN7CkQMMYUNsyQ6wBeS8LC7Y15dbZMqFzukbRZPPgkm9RrOuNkyiSwkWdSzr
vyz7Y1ije+wOkv2H5nB2aNCrW0trUbwK87LeYYeudIIPdK00b13Eo2ye4XYgU9GQaAyWWHedUYL5
UVhwTWezTf7gbFZJshCoWZ8yoheI5kTUA0zkAnph+JzBPEBtAAXQ9+E4fqGZzn7Hbyj6zL/n+X8G
Vx01GPxgKVB/eiOVoei1OX2iCicyuYmWxMZgmQFg76zfQ+uec5lyVWa09sxcafszlj+v06NRz76w
xM5nlBuPIgYuEjNH5tx/noPlsJlZCT+Y2JbayzhnZntaqm7HV0A6DF7x5yBoXL1O9NEu4YaQ0hB9
RNd3eqR+d64rmj81WS7sHt0KAGSQkHh/ci0JMS+Llr4Gi96srTaRxlZ+kg3Txgc1yme1hG7eoa1t
9ewmmURKvkEbBkpPRvVlx8X/+xiiUtdHIJ1f6cpd5LKcPfz3JlZHFOZR2rImeRHx4I6fuihPBTnC
3IMO/611yFkZVCxRy2PDBhdaKxmvae0Mavgaf7jadDa9kKqvPbKAJDUnvXc5Uk8bolpsX8e2lpSS
PSazQSPiSz7T0jpY5J46LymmoGxRG3mZgKkJ5Nnv7rMCs9/ojRn/NMsaQxTjoa6vlu7t64sbUw3i
fZGSD4GkpSad0ex22MWu4YevUABo0Ki7sacWC+zbuaI3gh0W8UYiKSsGey0pzCYMu+CFZ1Du8QC3
68snVcykMuI2809eI0gnAAnP8O+v8oCsp6QamfrgTlmE2J+yB9RUx6tP9BLbgtSdgRovwpygMeQj
nq3U28bFMwAsvzLalUiheEtb9lDEw71D/NG33Rim8LpqcB82pWFx08Q08WJfuqRMrwUp3dbLzzcF
K/6XHcyqp24h63h/97hupATYT8Bcg6+PELIy+w6aALBgT46aQEEH4S0rKRSyignI1vKVH6Y5/6CR
O4hMgHPEV3NueSilyr1ah57EO2U3yneuYlOl5a7cN1UukvDwns+4hILdDFUUcNJ1CuNI26IEMj+T
0q/kZU/wvQQzFPmhtY6nASckrxsdASThmIpBtTkiPObmzKZlv9+Zvb93zmpjmJCkG1BVcQHkvNmC
AQ3slVOx/RyqNkPDwTYRlJnwYMKrOQt091Vn3M3OQMmK6FyfA8fdqbbbjjN5UU7Ut6x+CYOOSdrL
teEJ/yiO6FZhE2GCxLdcjhFTZtsBjHnO8sCGxquaaJCyQjYzPHwoN8VLRSeLt1K0Fwpe1UxoFgkX
KDNU4+e+jaWqrTi71OwegqstMW26GTLOafJhZ8OPURpIs1j0GdqLECQjdIZhWhznJe0HvNHFw+Yg
O+ndtXP37dkO2HFzNfCfykE3y8VCBlVOGucux2Y7Z8XC3Pj5ETdYPXDZBkyvtZmwNAEybs3+rkFS
v/OJQmqy2/sm2ffOwTxS4cVYyeHtEoGrSFJmPZBHnUJAGev4+lsbqZfz0BdpjnbbHBQe038qjABo
XQZX95LkDaTlOdWRgUb8n8mvaICS6UTFluDjA443Ae+Tm5lSUbJM12q1eReObwxpFoom5zWX830j
iqQwnCY61IWsICrw7Ay4PxbcrWfn7/F7RqP624+TkI83BCH+DHRZ1z5A2YnEuFjowUeetprjN6A7
WAx0AUVae1uiKTinHQoFbEV2oYMRSGlmq03RW+nVCLN45uPM/zIiaRRt6HMT//BOOUhCR4v0W4YU
qymKG3RIxn1xctsFwnvxVZ5cZmP3U4GWP6ZlnkdOV76ZHHEmhjVW2+czrlQvCBX9pcU+TCPVJ+Kv
vhKld7N3zvun08+WfQ1EXQA3Wj3NXu4lwBUan49lRr4Gq3PncKQK37b1SRKm8u0s6MQftQSTmmqN
/WC2F2H02UgyQ4RytMwt1vlDZvn6VYbqDB5zQEvz+bSHfBGzoRxIT9OxeHhfWubwLkb0Q4LJSxGR
l5Tm7HDSAEzw6Vb2QeUO2s9D7ixakcUMW6Oe8Et8gQHqalpSx0TDzX8dALBeAAzwXzWqgMPv6ITE
VRoU4eSjgW9ETG08ISSZwIIbXQW/TFObcnF9ncZW3OQdHuqhDo++I7CXznYMYmxdsYo7veqlntUm
FCBNa4ml+DzNfHUX6GAJwQNUsZOVOmoyEh3jbLBtbL3hcc4xPF/q1YmhYRavcAfkEU1McZLjZigY
BKv+0cADOCp4+xpnT/B/VNHQc6SPkCPDTrl6Q/7E1pFnY5PUgcwpK0mDw7+cI4oWWFVr3Cxb4Gfy
Pdq1Eh0CNp3w2FknMysuf7uk6OZ39+q3dc6ytjz6p2XoF5PgAYzgBFpxMu+sbQMVhzs7e0DBC01X
ACfrhmp02OdQHHQPDNeUQgFH8MYH3f9RWSnejqmJW/t5GMUORmrkPwJvo/emUqBAyFW+g97B3wva
iIcOJQ+I7hRPSwini5TbhWkHqKpnyUxeFVXkddXClATRJeLLje+OKg9GMkcCAFT5GXKwwWMgAP/T
GcZ3krqc8z78k/qFmHqyiMXm2bYuvpqO6SGFi5awXqigm1AuvxDSn4GHvJzi0Sr5b10w9G4FjObv
0kHHlFwmnOtuzsw0CGR/UhsaYCiK7on7YO1IdJoqYdcqbtXIqlLb/8AMLHHi5uHtOZURuVf0luEZ
wgsgNm58dGv4PxT2dJP7cgS7kJ6Q8yHf0Dn1qMDQm5g2zwHP334DXDgp0xuPhY6DSG7GvfHGOmZX
2byp0EcST5tJqGpdsESVnAQeLU1vJKzxDK9+whcSFszFcEkcd5eX5FvwkYipjWMsr4Y2uQtZGauU
Q47aYjwF+0cix/h8BUxaCWfjR1pFl8zGHKGzvuTxeBm68hmzGO8V2W3W9UIM6RYpoKRy033gRTtL
cM7dcRNnEVJrxN7y4T3d/vgjqhHNNbupGyxCiVCT41iODxEgWka5mOkglQViFYOSVPJ2V9TJijxj
KJWPD+uXaT1qbxIaKpzxf7Qw9SEFdMu2Alq0h9Zh9981PNBhMdElKETBL/QVryeiFc7WC+h6ah65
NZEhdwvgPqS1a1YbJLVnkkDcuQ2vqVBl4YuzgzORWeh9QJIYnGA7iJhb42aZDBufYMuOlEg/bp2l
ZKQm+qFf/10H93xI/19mXdsE6tQcdnnSLb9MJjNVBeVofK/ydqcfBwh8dC65GVn+Xz17VzEXY5jc
uR8il5Up275Pc9zs5uy3aU1StTDqHctp9qSuyPacH8lwgUmUtMT+F4NwVYeU4feEBy/omJXDvNL9
oai+h1uhfUryTti7vC1bNKwYU0lKPM3rXivxCQyVYkDxNY/EwVnjr4Y5wUtHrkJ9vJRNxF6h9I2O
CncmUrWCN5Ib9Y3CknjSKNujg7F+50u0D+yCWkc7owJbuIBYNq+s97tIHQa3iLqOkneJdLVxyNmz
W9t+hHkKstUkSeCpqaybz/G5FrOuAjYmND5V9pTLdpyO/BWHXyTsboJyChE2obRg4MBvKAaobDHD
epNtYiC7c+CsZg7y/qor4FPkiXJwKchnMaY9+zTn1AG90Iz9pJ4Bk/Gr2HHtIvia65IQ8Elr+9od
zFFvyEOiFVemKHTt3DmffYwgpdj5PPtOMV3GeE7QoMMAcO1d6f/fx6ZL35py+jAmQZPdaj+DW+Rg
G45u/7OZ8V1Wuo7vHTHW37Qd/XBg9kWkpoqgLRqqeDtMYGfqAFNnyhDXgI1J3FzUmda3/huZisLq
bMk3qWcbWN2xKrutvjce/ECH7pJ2c+ikHJeYX3XB1kWPMmcTMgB8weppgV0GgDtJdiS2SMKdNcN1
bI+rL6Sr5a9mDauwfm/zYif1Q+ewQvnq/8Tnyrd44lq4/ivwZeu/7F4+KhqT3DzlTpru4/wxoMA7
KThdbua9TIl3F35TySDi+p1LHIT0npZbtU2/wx5JZXitlpirNnudEHZiq2pXXRXti0VvMQlyy2mf
aGJWMQqC24CuZMezCNFd9uWxxgr37mAymPXEg2AjYO4YJPArDZnRQU7paahSnQLUYZiphjA/A1oa
62m57cGiYjyjGdbnEh74TNaoBYfKAC00jZSOPFPMEVjKHf0qF0mF1QamrPyJ89W35Y9rqihmcJCh
IYTpjiEM5ChWDmmfAIlDtV3uQL4iFk2ENyAQKOOeVQeQsWUq879MV9WcVjJ5L3lBpXiE7/EOSvLq
o6gpWGbOpxfbXCn8yxswxmt0jf0u1Ukb1hNPONLTrBwwsXSI3VreVTjtyXOuqRF8GXINa6/OkBDz
0tp/pF9ijsXWEyMedxRCi9W9hogWAy2sJkDabLYUB7c7cfU8iEQRk/l43/Fg7wQHpdA1bTmQOOx7
aDiFobX6M570Us13z7J+uOqXBbqTATMeEj8As6RNwhsyVkQILG5GlVRPdF/s4hal7q3MU0Ee7+hq
n6poK+tWC7IRuFXOsJ4eyQGfu1A/zskIz4ZsP9/Vw+D8KCrwMqdSvzxSXmLnN3rgMmCLFh6l/xfB
qgoVPbAHFDPpzd+c/O9eRjWMGOqboqqVnRar93uHuAQB/BuoFkXJO5Eoi+kQznvuJYp6le/IPDC/
RLKIu6twj5B/n+PXPkODxZ2m+iBx/X9VPolQhaC1shs0ILYKKhKFYjvTGdeZwdzzLfg8Pknej3Cw
faFs5xzqo213aeTcOPu8Ou6573opO1oFlOF25wURTZdzaC5o9d1Jg+RaVN9hlwRASfVe1NtSTELZ
8UovLgauJwMRh4kof0OBgzjbzhzW+QlUdSMfhiQHEW8OzZ0cy+aX84HSyKozksL73e3u/+5J4JkQ
rTJcp7iNTGmDanCac0U3aS81E9ZwblcFLYDsEpm64oO+jOfHUE89DQSCjKd6/9BMz5yoEx6OO5gg
mLblhnarf8RHHFQgRmI2d+BUiSUw7h1hFxD8SrC3oi25ZbwEiqxEzMO40P60fB52rs11vvsO+ldF
xcg6hVDHNfhTBLvv7JxhokdREUtqaZ0S9v1U7ICNOcVUHlJsbY/Vh110aBNPQfDVUa05OaGbLAB/
f8P7OOAvvg5A5HQCpEJB5bJRwNXy/cNiwjWrLi3NfEEb5gCt0TmVgSz2JXPa0O8nBCdCOSurOmEK
eS7Mcj3XHGpBimzRjQfbBd3Tz5w+8883eCPTkolLrBEUSyyjf1nzW89UnWJuB4UAafux9lmsw+IM
eq5sTI7zpUbMuoC6XxAdNO3S2l6jueavJ2Y1pCeX3+rltcYawNru7PX/J1h9N4964aZRokQRuUbT
B1aJxZf7Ae9keeXerKA6/8ieZ9QCQsgY98ttKUhxjML86zp2aEH0XYgg3+hCb9jnTO7rUD6ldIIF
PVR2QqE1+PYynNAuqPhAQJaalSxgrSn1Bv7RlHxoTRQCd8II9ZY1rkYE80hShUKvthR7SA+eCc3r
hjj2ZAmaxV4KS4AfNX6mHsEhGLcBYW+IeA+4dPzagYpj1AcHThoby/tRq9wckbvXb4d+MO1aIEX8
+mJNVDvqGo1UiUjcMz2FNMBnZWsBZxpRhUvz3UslhNWj2q0IclG1+EiZMth+194LdnaMzBooeHdH
mCavMF6gHWafHrByzU8CEeKZeykrtweWf9iHWiuzTfqZRyYI0WCK7LayQOGv6kMQ71DDUpSBh6gz
Fa/IyXvVEzQFG1aru4dnOnaCmBu8ntaEIiN36Wzr3p1jlqwXQ+3AIwsiFTXsOWCk7qG8cL1WcDOR
G8axvhAaIkHI6GM28oLS4lrAT5jSdTZlAgtM3B0O7ZDB1pwhANX1Do9FcDubeCEeKCZvZjR/APiA
Bz0vAT7AasRBKbnOHcoBtcwKxJHtgkT31ddBFpMOLRIcHNLGFJk3UHB/sAAgUjV0k/fbF6+G79jQ
Z8CaWh279niWszujozeDOLWUNZFrkobdabMPl1ZyRWTMXpC0ng/seOFBr9bSdsVKYQTV/ldeOQFG
/x6AoW8Fs/n4CxK48m8IBJaSi80y93m2vboYgEn9mL0cgMeOsPBN7sFXRPdDGrIZ/soIspLIKhrT
D7Vc2cBVL8/68J/xVjQRAkI9G0urLNVXMw/6ysU2mArdKORBFUs7cq+956g3pfhNSVKb5NlSD3KF
1yYLt3jXkxqKNrURMRf5nbWPZyEjY6WBshxd2kTy4Lifk7xKXJA3tlyiwSwb8zUI5KX0PMIM/K5m
d+TOR3Nw4goteAL5rPYWTVhcXsNzEeGy9KnDmI7g9PLxTaJGglLF8LeLKm+XTFdDSuxyhZ9mMq54
kACNoVpvz2rnX6r6MWUnBzt6ga2LX7AaJW0rDsjhds4oSyupTmZ4v0wY4VHHuVDwsoYmd0a1Y/Pt
dIjkRYVgJC3hR5+NvR2iliPrz1xue5iQ9sdlDUSOqf/ZNsONE/Y8sHodLrLLkw47b7JvW+h0txO8
JZbUvoXmcvqa3thJcCVXrbBNGwjQBsIPy7arMCsyCwRXwaY4YJUC7duEOCNZII2jYuBwQsKFUYHQ
OIToNewHPO3dn1TC4KJiC/bmkDhOkwKaZVOh3XgDOwLYrAitNpZfUoiydVvAWV4btYZM10Kb/f09
B7eNc2w0gzJSd6ttQCk07GoPSaO4dxRjXaw4TcV1BLBdSKAffmwwKtOFXKKmc2qsbDEbrCe+yy9X
N+5LXy2p4ygeyRARAuudH476kbEvtArrmZPX90kKtvveoW8vKqH7FmSrRVv+PxdrpYwCIRg0VA2c
ESgKU1eef0BNSJztsDfqmJBqbkYtcDM6JhRCzlCUoG5tIfG4L0Gig0lZtf8+HUApDRkrGqiUnQQ6
eE86MBwpetiB+63LbPkurWd2OWvCb9kmEscmL/t9NRA/MX0+mQvM9aCnxkyIKFw4N3ILBJFfCsaT
wUvTP6ERuZ4AdYstSEePA2wUZi4H8Aa1lHVgtrtHiSqD7UCoZB6xACqUuG0NmOJQyGP1owb8IIsP
i7UWp56MOfB7aSJwRU9BtZ9gLeKnAwHEyTZEBvvxL3XEOnQus1PJQkA0yxkyaAHp6Y6aW5+FChJf
YFVUwFc1IZWhb8HtaiL8xXJ4nh4tJLnhE4Hkg5/lTr2ZuDDJMN7rlZrZqM98HgjyRBI7mqjvknk6
VWg7OkrZ830c3DmlDkhbSMKa/1mD5Y85qbjgjhWqITHijscd4m1MSVkTQefo6lL5K5KZPpnmX6gv
QA4xqBz3GDm3HmLIwLa/Exuzb5w/OaS8z/7WKFHmiDOXAt0fzine3mSAiAj/5gQGot0pGWsDMuaq
c/LtdbJa/aA5NTR5fHS75xGKQbyAdALcKXDAl/sF+lfZ/4Hc4ziNCM5l/MAWA97TwYrFiBL44S4K
oPgeVAW9kkfXx+9RtMu32mxl19LcoRm81stGPu7gAk1NdG/i5+Iir7vDPa8amNycYp4e00c31qXT
ripNWvg8LoYh6jlfCcjR1H5AcqKSiXFs8OpyimRkPls2MgngW+isVgz7YqE6Uio9L4nQPjcqGeuz
mbsJrMOG92kSgPJttuDvaJ8BXcshiHe2bEifiqmQpS4NDX7Y3BTpnC6ILtaDJ2FxawCSTzKdOIVr
kc+TxQ89kfJJr4c7oDGvOZ+pj62eh+TAtzVsYvQOGvapW6vTvEd7uKzCvA61bE6JvYqaCT5Zhsct
pDq+jvy0mYthia3Rq4Mdmc75tC/A4nCdDZknLxHdJxj+guTgasv7p6/l0n9aPG3qy9mkiMn960ZZ
j2wsGlA0Hk/jiEeckPc9JCQ47LRybVMA6fgAWUMymiT5dr6GaUDN/lJrzLYbK2DmzWQovRSLYCQC
A4DyihqAupQrifM+g+FYA7W69YQ7AJnjFrfjO8dyJkMDDtuHnDweMnv9TqgdrqjxPQXouXWrvotB
cbsoJ+hwoENx3vY3hsMLftvi6PG9C5YTWxgM6Y9vT0B1DANgwvkCGD01dg7NWqLIBJ9JCHe+RYuE
ZQ5PcQzx4hB6GZjw/dZXg6ULeyBYWJzLMQt7cp9wxbh+IMDpAJxkSDPE58oFFMkxhCsaj4JPZ75H
wRuK2jWTw1i8NqLOhuuzJGV+CEdcUQJqEZHT8Z/Nd5c//zuVNNc73cuaiy+8VF7N6oQaCmKljZ/e
3XqEZFu5nubRKB4FygETigs5uGyUuDqglOHxrDZE0bi9I+MrX+Ug35njHAXAAX0YBr5lmSsv4Q1j
cFnHllLCiXhES2tRVp5Bwnb0F+vlLCgTti0cTm5m4uhEPeTWALAdbUzp3ThbBZBjVetDgJDotZWq
ymnfcCwMJfPGtsejvubvSqD57L6I0h4dJQG3jIXUDjo1BTsHG6+jvfKFu4ck8Ee8Q/QVDderu6D8
Y0cI5mIEuBgD7KXr6WpML+bdahRZ/OqfSkhWk3WIQrNPxB+Uw3cr3TgXPuvhQLovSwxfO0uwOr9n
amRIgtKS6KvcZvadtWzGXJXYRJfd9klcfGLlT3/q9AXcFJ2z3vh9uz7oLRtlQrqWI6pG/qmSheSS
MkfcgzKYL3ZjU8IUfXqnsVbhE80+9QmLfCKZIhDmW8zruG//yTsrx6uWQ7UWyGtUxhP9UidR+4Rd
1BIwxoFSKwjJ7R1YRtWeHcwiD2siMqZfwEFiDZqWH/atK8faRWqfOC1NNtQE5ihfoQ8XfBqd3BPt
Nu2JCFYgV91tJp9dYbkmdJLkD3LkMpLb3jg5rPqPPSOA7yS7Bx2yUWL934fSSbKGB3udDXkGrMrS
ilh08leoZN8bPdosc9AjO2DBOMe6q7FUM9f0Zg5HdRXTOoqNqJW+yEO1WhPBCvpg8Ga/nbPjKVm6
m8ynUmYOUXZ3i8F0NLPSQX/jOZ+yUCzg0GhyjNGvazozStpzE5CLqBPOnfmPfprdVgAu3BwOHZzi
RZFL6w7/14Mh0Mg8luMXKeOu+0jb6rEpzNdlAXRInglNtMQE6M3tY0jODcIoJ8EY6WOyGwAtMmIA
jsnAaDNrcedKfRnl0sbUY/Ez1Jf4uCL38VXqmR5XcYVqlq5DPDpuaoO7a1qaQ7HKLMJeJp+RBZJP
X6dmJ7mPBp1dH9ILS6ZzGT/Tng+76/ksMNW9s2Bu2BZa8T5wiG3lsmES6iLKF9fHvrb9cGzIigIU
PU4MiNTO5xQHcYpmfRoEczGq2wkHI8vM1SVteCh9xcObkBYgCdFrdGy122EIGhiB1mdCWeFtaTNK
SaGFQjJNMuKrhQ8F5NN5YdEA2lb4sEXpEb5YVxuTdwXLOJ4Cx0QQnqpN/Jfbh2puTP8hntId0mH1
ywXnDzYJO8iKg9J7m54wyMo4mcCZ44vSpnuwvEhnyMjp8fVz+yf4fBV2FN27wltQzuBNW5D+GtlB
3u1fU4jqp2aRBlbsgEXMbDDf1mgVneIepjI1P/vnnCCRh0olXFxnUx+Wz+H8S2kSqcRsCy32zlni
1QlVPy/9Jf7r3FmWHgQEnE3TU8iGvKOU7NTaMA76Prh/CBqWKGcfwO85q94pheVFGnF4yHvFC5Wy
vOcuplqadhxjtHEGXE1U8u9GJMfeWDYyeKTUkShbhj1uCwOC5hrT3/15j5tL+ZM3PnFWNoqZ64go
K6wo+I6NSmD2BwHWWF5rTax1DH9Cv0FgTRjrcwCYNISFpiEouBTHY9ZLCffriQEWX/rYjyBNKKpV
QN1+Id4dxC008Bexk+Kdq3Wl+G/2LpmiimmyMUqJ7gvcv6A8x+887xarTgC5X4IalMMumM1G1SNU
7dc2UfAZZY6u422eV7cdd4F7Ed+vdcumVisZ6bmnvVGZyuEP74ECUvXuVWvU7TZTONiZlFqyyUXJ
jgS3f9rkwI6gyX0Ea/vhmgc2rMJDtocyqRST3SzZShOuDPkN6o2IgWn0TI+qahd9n9vu+USMv+KH
j/ZKAYlh2pcVeW3o6k6k30vT32ck/B/+AutM+4KSQTgZqN62HPqWLs+3Le+BapkdMrdmlGvDS4lP
DvQT5jkYsGSaJKcBW3B2aQi4bRh7WbmaTC/IxaQVRRZTGSQy/MBnC2JGXiZVGGNnm5H3WbStdCCu
KT8asQ/rjPzX2xsCJYpyWX/MAmvEdoJhNQdYoVlwJaP+tcvswqalc45Xz+TsGYDtXusI/ZVMBQcu
lf41gva1+O/LHa3pphKd3kCistXYm85Occe6RqTvxR34EaUXVD4GfjsaLU86N8IY+sw9hCZrlgZV
oiaD+VEJPt14NT/vhP/r8ea5CymLHoW2mowpKL+Bl+9wNXE4gxNOpFa+C0BV4Uy402KMjEX/uX/n
PXtWj2obd//3a/HaxVgIp3Yr88+jwXYM5eTpblmEpSuDW/jnj/kkg/l4cDQJlUTw5oije2TC58cN
3KxAjOrTy86mVPTFyeBiYZHY5zcrxmZwRsL+VDeHD+MnpPL/MiB6UtcVlNZpD2KH+59u0m+yGDFM
uKJc/zqXczRyhWLWQFReiwD7ZZuWIcJaNsPdkvJnn2zF6ApTLSTh9ZCJBUpcNFzPPDFxxgaMaf+K
G9/3QaowA+p+bpl5pMFegtOx9oX4t4J9toAvheuDlM5oO41bRF7XjOKY/zmpI2IgB/0Jlf1o+WU/
oVO1/hW+Llk/qjFVIiaVE8Is4VqVkSMJ6e4h1oRFvOvoaC13gpG/I454TasEyPfNNEtCWZ6LHv4V
BVaNOYtdWIgm44RHL2mgHCMJFMGV0Dhp1D3L6OKplD02gVAaeLoT5rWReuBtPDRVp7Ic1/YQ+XmN
m9Og9q5LESR5ZsrrbwjBJJkdNXlybzSkyoaf4rY84kXwqYa0XDMiwMVzeA7x7F1W6rVcCyYzToQI
bfZzvoDbYyefpco4l+64RmdiGDc7A+M5TWx/63eIHaX/ZaPm2/yFtxiRfFE+ejrZmlEzUMw3sHho
BiiJD0lBWSsGUgbEw/rAYUB4Q836DQ4AiqZ9NUMpx8lCGY8Csut+/Pa49KV20PZUyO4pz5z1Z/oS
A3HByUHcgoShrYW8VhXIlDuSs6yEwHgVar8S8UPqc4Wuqiwisovu3MccKkB9GcxCKWl0PMNbtYun
0AhmdyxfoesnT14cPij7wSBGT0kCRr75Je2K4OntIKNIxisihwSZQNEIk733sQfgrjveb2y0uDsV
TdEHyNl9e/WQboJmET4Y91wpBMd73GghgKJQmxx9Czssij7tx7DbHo/uQl6GpxtAY2mHUfhBnccG
Cc2UoW4bMq2KzGNpzaPqfffLqcFpK+1KesO3W0rj1ggF1VODWtI1r18RxM38EUh+4gs5M0VPRqdc
ybwpbqRqJNcMzja9esR4Fysr6A4m86gRHQj0/h7ACx9IiN4QTj1W8PQdasWkULUd4nNYw6rmVHb0
V1xQsmYzHIZ2zSOoLkXjunh4ESHllbp2b740pgiDjLvICqat+uu0i4UL45b9yYCSM/r7f+uHokAI
m8UbY634cx1HqgCB4G9fC1O0NSamhAo1rxIyQc+AmCb6P7oAe//ocWhoBr9zZHtbyxcAbssNd/by
s0M1Unxm55W+zszf7rf9cEAoU3o9jyFt4h+/G/tN5f9h4qsZgapjxO6k9OpztcObjBsXSYy8S7As
qPmfYhfbuYRmS3bZhh+yYp5xVZneJyZxJXFrFHrCZ+utRYulyDg/3EYd2vZxHoZT+fodhM2D21s4
ELLnVJ9Cakvf0Ozy0OVbdkH0s3NrdRZXjYYr9Ylg1sfqZEmrOgWFJ2ey3yxQ3RnKR3nWqe+6bjbw
oXWbiI3Gb26WpLPQ5zfdtuW3tfY5hlKDaN0B/rNUmee05fulB6hiEohfy/i6Ivdb7IUP5rX9aDOj
vyY95lUNuhA9CWPLmnkMe1sKnriVaea8IgYbbwkWGgYVGqDn49UL2iYOjmcYNpnn5gG57UqMGuRQ
IHpbHeX8+tO6gpejzrYCcYYmZX9pHaY1IpnHeuJogSOxb28V64mG5OTT3HHCwZn0vDg9ndPHn6sD
d15HmNd9nTtSFGbQMsl0Sk//XLGrz8jLRKuL4xtHJbESAzkESqOi/nk34Ol4QZkko4GqoxK4HG1M
bsMP8GmInhTJkeu4j+y4B4uTpyfB6UPX2jmc26dPgFqIOPU9dXRMj8//YtwEMePWdEdvYUFtlvUW
bvV6C7thtIPc5ML93qyl+SiPghyibIXrbEjizTzuuOpJul9w4zJjsWaLA0hcGrADqmFtr/1Yivfp
rkGwS9rYBwhPVgBeOcCwsXrmEdCB8/sgYet+DG0M1149finWS8VKKmfWXtDi2nqGoGjsDk1gsl5i
RoDIKXyXlN6mt+Z7vrXsa3T/ZxBpe4nzgFPdj5cHAknH3GEovzMIaeaA7TE4y5lAvUoD2q9Mm6u3
683a2ZUPMYxBm8FAFxJPJwfzHfi3ZLr1TjqjK7OGmGHkLRszM4Mdd1Jbvebk9iaz0VxdPlu7uBq5
W+dWCXUW0XRq/sGA50vf2F2xslCokVdX4kOqbisgfi1ijxXEesggCpK+mzTyv1Uin7iQIHIlm6SQ
VJDXyfx6YddYgaaxPglZrzATdBC3cay+rfW0AKvTwIc3N4fgIal6jkH5Cbp5pvmXpL72ZNZg9NYT
7Ioc7mm9qmmJXeX2d5vP6hCEUDv0/zeJeaOWt1pfzHReIc4YQgpqFROHBuRlSRXvjmN5IlxIkmaE
IyHHEfCKg3Y5Dcg0IcY2TnEss+rwRZ00RUb4fNl+Y4GTe+hPS91viyascgZ3nl+D6ZIpLZGrtY4F
99WE4ydFH4ND1RddxlXE63mFt3iZdWtMYo9cXc+jZ5BAPE9cihTfssrPdg1zxY4OTRx51TsK6bzQ
DXOqT7KrgP1xiJW10WC1qKOqNNJ0/ofNMAK3vcTWm9VPPx9wTvvaLTP4iQWPK0QZ67DWNMmVpuzX
0sM8EBiIJi5yIFZxIVo6MQ07bCq+gayTn+/f59dLzeCsCWP3xV/JKBu68HS4hNE1jR0bgPyF0Dv+
OO+Nd46OB/fC4h+GNEG7xOANYkN6w0/o9wqPND5GMht5LfkZVSXFUTDXL1JKsq0OjQ8KJpL8jXiY
xWSBmVWrb0miexOdcCEOIqHP7qlyk9ly4nHFB8tWfh+MLHxqmQV+hl7hkWTq/6hXas1k9lqc+eUg
WWnmLU751v1MlZFbtlwTG/00VvVE4Y9TMoT6cEI79Je0bRUj59SvnfZqFtEI8xdT2w48FVs3/GjW
lWBKXLcVjXKKcT/zH0lKK0HkRMRxa7+mGRreP8ZSwkkALdkP2czLFGeblmWFmZZ2YHkHpDIpNu9t
mn3AEnAzxGSOhxFFIJgRquIa2geuLXJcrItCit7C+irRXSVFAhpNOgKGkneu0cMCEEYO4O9m/UVa
b+HyALjJhITNsQWI1DQpPjvjqexe1A2vSfjnb0YeH5tzjtkd2PQ3r8327w/14/nNk2pgOwbSiFj2
3SQ82c28xRoa3Xx+lPDCOPjvfr4PVj1KYRdX8BEOOeKCYzHbY7yD4ACOhCaIC2OH4rh476aPT5v9
bj/UPIybfzkdAWfUbe6yNUAtclaht9a2yN4AkRo18YstHcZBel9wk9YuYez2+TMLJ64WPY8vpTP2
W+vRGv3tfAcPXGnY2v1CliCtxVK3IaNDTV13t9Pt6Znxgj3OL/zDC4FPvWKvRINq488HlC1HdSVv
uxNjrt0iDP9wEJRVeUWsAY+YZKRf53qjMAOOx1SEKgHKLgkZ2x9QdNk1vrvxe3apV/yRir+iytSF
hSxY/9MBKxDo/xCVjzzfvw6PYFKjnVp0F5SwnFsrVebDKHHkzvqtKTUsj7fsozs7Gh75hy2cGlEz
8q0FqWHnvollnC5YVlnYN6il0iyargRU7b3eb63axNUlSp/EROAO5V1sXGvAKf2KdWEU0cNF2kuz
UdUZmRIeNZS0a+WarRezcnJFYQoz9irpNekbzLl2FBKJRG2MOLINxE216EJDpDf2iU6KLapRKM3k
4JCb+P0n9rhNbbxxW8fq/+WD3Fsr8hXKP+bsZGsRpC5vDV/hhEvzfiLLIwIPULjDqhhJXGkh0XHM
2xnUaSfe6KAtG4KP5yjSXm19jdaWkIhUmiBiy8tClUbctiBfnzXw4ttWxhYyaRPMWjV2WKlYWuLJ
ZoQZejRNUk99tw1NvxLHbz0G8tB5yIa5TDiZAJ1sShXKO9+DkC4Y5hzFh9HHQb+173qaPUrDjVRx
4iP0IXqbYyNXIlJ9aF9eRyQUXCyNGyq2d+tnTiTWi+AiJ6R5q75EHCcJaYww7xTxm6f26NUwowkB
7i9jOGH3igCR0OQHpA6gkyKf2mQzUbHVAMVZxGc50+BBWXiwXBXxuu0tFtCIs3tJz/R3ENxYqWXu
EDLOMoTaZ/IXBX/U6V2u/37GxuGvjnhJXLk9eVFlKvrl7NIhrdpE2enDltqESmmZYhTthiZ/C9YS
tMvWe+W/I6gYRCOKW+T4lpvjHEQ7ekDfhHi/znz25O5NGxfuR1ncEiHLhcSabllpUuZO2UKbYfv/
giSOTYSl7koz0z7Lw3sdtf1kafTi54fEyd0dMh0S36igld4rh9wNk4qHwGTCsPAGoKuDZX2ERnoF
qHekZMLTRjcdId0W83neLErh1oYO+CmRKqIjMPb9HsTEeBVpu2ahRVvCVkTs7iO+0tFenU7GIlpW
Hwh4h/3bUwyXdZ7wfQVzDJJ+JnWnVUsBx52JyxAc7GdquXdA1tgSRlHMbWlWU1qhSbKSrfdzVWiB
FoOe/H02Yx99d3gGnQPyzd8UyN6YS8mKe9a/kXKbcgNE3WjbJ/OB9bY4GbbC9YuloI+9G3bB0ofZ
35n9kfCrebrXWOyhtJftjOAMwDWoSW0Mk6kHUZC5OEl0DctN3AgWoPC2RRboF5zcsDgkShEwfc4C
R9k6mK8zFWZdXqiqS4yiN+f1W2epUmoC31eXUIRhRZcao4R05/6HGzYnGKW4mlK4OFURJF9HwFn3
PiqWIz+LrfXJ9zG4S3pBw2ZPvK0Gqkq100aUBwShStGayf57AmLOVlKcTclaU890l661CWJ7BRtt
CJcV0rbr6vU/nFTQlATQhL6p66+jtqqJobgeVqmIqpgAsxJjrr2ctkEtmvlWJwJLhGSTcE8v/l2Y
GDEyh7YK/kdPKoBjlqIo11pfgRdmKFOI+dcEm95YNAM1gg4+lLUxMakHZieENSwhf4jjZG9jvU2u
L1V07NQAE22NqcoRW31zBO58tafYAaTe5r/1EgQFhOB7fPRNKURKJkeyeGHOzFQfuGArbhEA9Mom
KXdwc+sSgI+9CSP116+KkZRvsUd9hspPJ53j3hvZrMRE9h8az1sti+L9/sQ0FLeOLZZQc6PkAiRF
+9Y7mUCOYuIBbI1u3Pvonc2UA7HF57p70OcGAKo0rbAkxqK7Spacn5HSxKLWrsCyoDdsBxwrxFsD
BkUuCnUwjG54XiFqlByFEVVLksxX0+SCdpvyjL+hcAJaW2asMNQZpEoPt8JCAidED9PsDp2mgIzV
MzxLE4g7d4kL9NOhTZJsufaj8MBg8V6JwjY27LJgy+/DUDsQ8kOjKXpkE6iSDqZWgrVZrzOnDpTs
VgaZywtGHJnWgiur8Ws7FLhxLfxG5x7rLX9wgxFJajTRZ+trEUcZezRm0z9xwdO5gEElZ9agcZlD
NKhAz57h4dmLe+u+2HR1L5xDAUrOHXPGdK0JkUzX9mib7Mq6OfespMWT9cH9+8vJiNQ7quffHXgJ
UKsPoM6IyvSRnk1zRwfvpw9yUbS+k8FQQCCAmuetrc2qrOLxrG4BXNmSM37JDdLII2wa1Lbkt212
xpsarssugf0PH9GZsaEWyAvATaDTfR7PLU5jRBJeQvzQj5F5l9qIbHtjDxsnSMiztp6fq1/8HYFx
o0JQS0V6YK2UtMLGOL32tHfoEsQDdchk96wlE6zQw4Ffd0c1fang8bXLgLVYJSFLRaHxeOE5QLGi
W5BQ3qMfmc0k9nUJTS6H+f2sMuMjjkkRaGy2lD9JyR9ljH3lDpUy0dzIOlBXGpFkqUK8Z8I9s/rz
CQ+eO7pGrzCSu0sSMFvbyCzzHxJnuzu6ONTLnMX8ICYEehDJHXJZfzQYmwMzypFEufLc3QZQNew0
hSCFpGf8VEZ7F5u79cTtuseZutix3yfDVAP/GWZG2UkInA8hdTA/A4VC6drS/A2CGG9ql8uZqxQQ
z6AhpLjafeQZBZ93D2u35gfyGKn2ijsuY9nceO907eVVSLMgAmbsiZAlpxsnV5TEyEQalDBmtQaM
JKTpTTnln1BIsLMHoacmajZXPBZaTMEYOvwvhIdhpajUHZGhlePIKKwWWUKe4UHJZTHSJ+hKvhVH
e9HaDbZZjoF3v0w8Bj8P3K8URz0586MHHN+/5Z9eFehCImARsb0U+0FbIbb4uGPIKpKAYrwFJlBC
1DyJp4TkCnEnjEzJbIEcqI4R8N4KAYYHKuhah4SOO03VcW80vFHdE6itU6dBixUKcev7jb6X+G+8
uJMvwPubBQnY1qUsz1/RswGWpgcHQAut5W03keeY+ptXUeZojZ9Em9dq/9RsADaEnqz+CmF7hh7R
Tu/q2D/8JPDj/d55MZkTzabfGFqaJZRRUYkqG7vqWzvWWooCV7yKLR0Nj4Fp+hIYBhD01KfAqlix
dpN129BWg4AMHoXNibtKycP8VzPWK0JAl8PgHDJDqrtyHYSOusEA9N2QjTf5WAWtgaR9NHdhCspG
pqJMZf9LiRYstuBlrSJTGRJ4t46ktgY4u992R8Of8HYQVF3eik5CroLwfmxJBYuEOhx/U2Uq7Il/
77h2wEbvM/Ya65fMjCZykz2SSN3jUmpozKhUWTRbbaGYuAleyP9SB4QWDOuXhFyUrfOkbAJquH9O
VeyWwHHHxyh8UfXb1rjl5r3amFrOSXfp1CUMqpkA6yjjL1iPoaO0qaT+XYiM7sI9d9k4MfPc/Ain
jR6rBBhSi9CGyJV8V7z9yxc80ZK0znLyK84Ns8tPr40iwkPsueXsszGaplZpFW07ajXaafGlpuvb
qv6rvJnVgmljbV/stblfTlJc5s2AGVl3hbjUnhmxuojg0ytE6/XsXjz231UBqNnxXPbfGFpPPsPm
dOj7dEYKbK2hOokakppEnNyx5+uK2ZEr2Nlw5DCiLyKBkN1AsTiCmQeDobmpdKYnHUDp2OaXhm/E
PMI+p3nRMkh8HY4Y8Rk8jHKSaSItYbq8vdW5F1H2uoLcZRuRHK2LwpHWfNfgmQ4CtdtQk2//0aKo
oLNm5SoolE/DaxR6rqXixZLtsVqUspNwRfBK7DCtSn0zEXfCuMjh+awLFNjP4Qtou10U5eVLJPia
7s3FPFt1xF/cTgaN5jx3Mn5AO9qUleG5p8HRcidEHN9p4mKbfRubJnK6nHvEbm1rTeH0dWXIQgUV
Edhp+hsksEIU0sSHjYBugeldPTNkRUxZANOWBuRlYQrZzYyGG+aLWjhCp+8H1iQO4z/+6VB+Rqk8
PmAmet1Bwa87BkStbe+OsmOGJuKnLmaK81+dzApkSjvZG3KsOlmEFJZWB6C33WO5mY8R0EEUcMzv
gUUaxyR5ZVXZe94FK/2kereGOwB+o8XRnmAOnVZdXUbqFg9lchVDKx/AjKehXPxLDsmHNbnLb6Sl
0h5yHCQ7qkRLfOVLtSFnoyd49TQ5wdIYDyPDUceO047BYxjpcg5f4aOSfpejZggU+SOS3xKNYV8K
9ELsz5+YL9rFqcICecamS8bcWNFUL/r5N7N9RAyhXIJWTZcxoq2Nh80tVYHAHJa4kOjji8OfHQ5p
7tcmbC+zzN6HU2HbskOmKobl7Iw44zXDW5FoSSQsQwkwzyM21f0WN9GEZMm8bd6dzqpaa82lJlh1
uISv2BvkbLc7biOHLX/TAecyuFxcBrr2ibqRn+BcLTGiPG3vrzdOf5f3yyTyRIiJ3yuC5k6HA2LX
kpeKYn7ZeQKXO/hsAC/KE2CTBrTiVHQd9RTUZXGnaGF6TQd70537BEw6Ddz3sODdc6XS3IPV26L2
Aj2p9ML5kh7VjIJTYLUQnF9GjfVyR6O3aL1hSX6eh1Ruu6+CWcdcjdgdtAYX8ADMJXwVMvS7RMNf
N7u0tQbzFO9b3xxSnwAv+uQrCqbcShQvov9WlnIL1SNDsXF5xLmMlzk9EdBlvekmJXFXQj3eicRX
02NFTehbrDDbPVKmOzUtVx5Ot3Lv7gkmTSzVdR3tbAglZ2VeC44UVkF5zWH5UtYMkD0J3tLBMf9N
0wwPrKkNUaoBnTyyJqfvDif1OiHmRe+nErnPblgWxZIKJifkf1C2G5N3IdYXoI9vcRdiPTEyuAHH
ekhmivFN4KJrhF18lojRsh/FQ7JpZvWNm9hAVSc8fs4K69r4S9tN2h7NL6DK4YlP4b2RPjGziEOI
Mzf1/nTxO6qgSqzroR3FWdqwjakpEb8QxC9yxtemyf+QAY44GeDZM9fL8dpx+BlyWxSz4Q+wOBlB
7DZjWICDTxiOtGNGxKA45ceIivqXltpP69pU1ikmOa5KMFgICw8RxSFbNTs74wYb7E3QizuesGQk
YaF6Ag6yU30NXnRU1hEmho8cgnbcpzOOlXVRp91J/J1C1Vivzy4dNKinRp4lVZuXftvNlyOjy9h9
FXax9dEB7kf3PXjS0L0tDxv6XcQDcsfRHqm8OxG1fRiA2yMV98tuTuJeQUHy7d8oGV+SU8J8wFXB
S8rsAelyG7QI2KiTWQ8/7RKj8q0J8mET7g8SgT7fegWQLuLTO2CIMfCWzSVkpaf3zKilNGqtzM2y
K0CW1cuilEWCXVkHRdu7AZiGQiMYHidozzymeNpMTfuFa97AsN975VxixiQvraRKRQWx/ZwTtQJj
cWP5aOf8taYQKWiE3hLLTMBl9R+zxnr1WhT4yBlKjSxo7+Vi2+BO1Upw3Pi6XRmGpfR4/zCJthTB
7TxxENZMbRwrW+FldTDZbTOOK5SFA+1WzFQwdfMNdHeJeDVtMEAz57Sj7kbTkd/8BrJSBIKVo+9s
hJueAYWsr+KmyJa7MimXcp/kdGF9B5j/NK01671r5BXd0JnkoM4JNOAa3C5DUIk8cjDXVj0qRYg3
Hs9jeP9tr0zTyOikxAtEolhWzgCHlI3lU5UdenMXMEvb5AKueNxp3N/xe3C7GAH8xyefjesuR/Mf
wzeRZYbh71ZAGoYshtJFWOg1gwOO4LrACA+bcfIAmlM9KKULOeJMXQr1TrACHE4prxOo/5Wwdy+l
k7TTz9ay6Y8NLirSy2ubwBCrMicQQUNW2I8ok/q5LRpF3KJ8P2ARfW6zceD3D57/n6ZPPSplIVxz
VdNlxMHz5S/+zM8bypnKriIvSmTCXvdFFgtp9X27LP3uGzV0Qlep7AazIWHuD1FAAplLd/iFBZAJ
FUZiTf49vv4R8KeC9WWngjpxKXsYuLJ+IxYjwMZDVTNv/iAsx+3qnmvjTnSXVvRXrzfxWDE+rPYm
uckHbiIiGHgmxjHw49MzNa+vkMQfavU8Eb0E2PTIaFRoFllNav3K116yqQd/VUq3hiUJU5QqOuZo
xWQKdUtXhAK8QYjo7lCw+I9AuYWRe1XOiFUqSXupUEhnparrW4R3AxY4DrfuXdUQGWJg5ww02Cyn
l0LjO/SapXhRBiDhaKhU0HUS2vQVESfOEDevdqiCjT7h8aE5cu0W7tuo/43GIzr1gpAJa9JCBl9e
nFQXHU7x8qOxTZW4pksLNPnWi6QsCLbaLm/xElAZeMpQy7OOx236b9spNJD8NIuiO8jh5WBFNJIp
yflA6DPtA2mo3X+LmSMwvlAMmOKpxvVj5OQf1i89q4ajQA6bClypfWUNQJi3worqznN0CLO4Qw4k
cJF58NPGvTeaS7Pb3+p5FOZoTz2zHw28HPOglBzF8U8F75lnIWr5HYZtd09c8eA91Z61jdMg6Szo
fN4XWQVzRFFTXcGQ0Rxc6GRNEdkvQscznsPAwLGpVcD1uNBDZhT07qnXejLdSIF5+irWJ0uA/VpS
cjMqyzVwTWHWLhLDurDaZ0euuHcJ2d0cSYJsj9xBKgrWyGZgBpqMrQl0KOcf/LZmVFzDjvJ5irsm
17MtK7nrp61nkas1uBZtNjqjm+VVTByn0/JRn96pCUOqMVNXbHnY/APZuse0eqZI/X6x0U9qWchK
NAUxsRJakFax6l7WDSGMGThPZzgiiSBTfG0E/LbsWOvgKiqRP1RjFBjCyMqjDzkewmuZ2lmo54Z3
Yktzp2FYM2MoxRySz0wtFNEssfEl+hAcJLZdwt0E7igdStBt4/HdBBQ8bNpyZenDa27Ojf+qepSP
z3YUBm1u7Tjx8scMM/iQ2/uiO/Re5M0EPYBkk85BQQMXk/+YaLM9OV7xX2g7v3IsRg2Nb6uTasrj
dIHCb4ca0hmFqHkt0Qz4HnHkoOap0mmdznQnva42V1RmyW3ZTpO1W+LmzmT697Z0Soewk9RaBLZv
6Yms21qrI7Y7VKW35LNqrJlH1p6ZeXwyEA3/x3KP5+u8JogQwRIMtRlXfXtBmMlDkVOwqUYG0xFR
poaTN8WpGFmlgDjR1j5MVycZCa646UdBg0tfbdZgI1Wgc6yWj5YUwkrdC9dUIStK701QeROJkHPh
z1LI2t4KR+v+CCbK8lLXKsXfny4D7WFgNm14I2BvxS2lMShV9zRUw2K6lCbsOwZ1xXzTzFWIHGA4
ZMwBbll3v4bvbOaDGk7NBkraKTM/90yMKIpFJbxH6PYCXm8Xu5eXA5Ml1Ywsuq8PzBth77tkWXm2
BJNvnNw08hCRcBj0SuDcynwEYRP2QTjWF/Z+aryZo/g5Zyqck5I19VatT5rQV/U2Q0iccbSmfldD
fibje+o6rbVb34lCoalP1d+rPa841jQg2qKNotQtZhayQvT8aNNJa8sPrNa4iJJS/zWniJhV4r/l
4DTEhFnZ7fqreR2rn9tyPG0zbfOBqab70QaitxkoyVSzo24m6+tuas5OTXqVQmzOPs3wKhv8zWpR
GWLTO2hsiuzrrgx+USgobbX79eQxgJbgf5OnGvCrnMrlFftpQfJsy45LRUlbq6wIT14cJRyhoVX0
q5522xiaxHnA0/ymsEUM/BI+Jh8s+QMOGz0Wc/S6I7jccGu4eUyhbkfcNsHJsF0Mq2m5vLGfE0F1
ItM8cWL5eQX4LPxbqUkDOb1bc1XTmu8E2YSQSUJQLJ593v3kC4dcY9piSrj3Km6PekpB41eq67uT
WNvd/D1Xqyuuc5bfNgqFmz7z7pfdeeRxnu6MglFXF4XRxnOzse12KYQYAE3iu3igqwbK46zHtiPA
mtPMlaAGgZuUadoiOi3bpEFgE23FWlBfgCPaDJyZ61CLADx0NNcn8QegoyXbz7v21p5IeUGzPIy/
q6AHNt3+SxjcrW3HtAPIMlJxV4EDCL0DmNWCBsLveFYKYCqp3JepKktH42ZZTsudfB9vKDCHABJ5
Vm0a4MMhFfOs2VmoXmImn6l9KHQNhm3nrkK1DXz5jXblWKKwNZpT9wZuKb7EDtka9Ej93Y7r9kSf
OlQK5ZkDSdT40fdxI7MtEnnByi2S/l3NXYm3tBQLnidzJo50hBprokm4s6lWj1CfreumXCQuESlG
yoaXiZC8X3ObhmmdGoeNe9oJKbg9dxh5s4QXm1gi0k0ExcyVBq4hmKn/jp5wj8PZrNEsFMMhrpUF
rnu81/lQ0HNnhhtY6x6Z/x4k0CpyCfoOiLEY4p2YFRQBM0vptzrV4hNY2IZP1ma9+1vWmi3YAR3p
ypO2VQuy2J3x7WOE+M7FpLzuGMaKdI24UkkBWznUySdo6k8TqlbrjidQxsLLm4p80c4Kcy29Kmbx
t/OMWnaOVm6lLX2KwxjR8bS5raLDlyCC+ml0jnCumwxzgosXacVfia+ZVbTCjxWosR0dD1hj3ah+
5dWQa+S5bVahkL/noja1IrvSEI3+PycxV/4c3G/rOjq1CHdnNGMKmUMhJU9rvUn3RlGbCEySeYhp
v53m4bLWRyotfOeccGJp3EA+dFfZEiEx0Bl1Vab+brmnPxI3cQOlKMUgh/COsyiUOVe0RUCIRdxO
Vx5BoUnl78ZhKhusq0cfz4mU8V0c4p1Sj9pSArGyJ0VHIxPuz7eB/mJHf6T+dvpdc7cKNla8kLqS
JgwOmLuXMBrMLMSSIMqLvJnXlGOJRVwozYIEfvXQXY0+TS8fPIbu316SZP765xU2Vx+zxmjOngeF
NbtAZgW2gY9AKewiXurpgNbbTJCxwahV0Yw2ob3+9WDQ73tf+MAFo/tZTjVQo6uOCaO3NeWqZRJm
5lTvmf8tHHXYoBVdYOziVJGfoqYYxCfAz1SLCJ/Qdh3JT1Q5+Z2Ry5tuwKGtGND8lUwqFrbpe0ft
47nCiTyaiarTCkgIj2/oBq+oW6HxhffZM0l9p1CfdkMdLsJsSBF/z9EVOqXvt3AP546nCbb3nKUP
64vQFucU1uvGa5DrW18/hjhKD+finO0lo8rFF6vM7Jm566BtMF4hD/qc6u7Gd67mEsNj0evqr0bv
vdmro59VeP/iGl+tBTv5aeYHs6aQGCb+A788pnd6j5/1l7BkJm9sDE1JzRccHM2qE0BKQOsxq1rJ
f+Ux4Fd4UrqORUbWt05km+V7r2hJzasyirk+pHl3y8yU4x9ccC5LEiXlhrU91S7z8tSV7T2HfKUj
wYBw2OqGkhmH383/vJLk0pOfJiHU3p0zg8x/hAfXr9otUoE6fQ1yZzEjSq1k6cx7+xaXLDm+9st8
gk4GMts5BsUu0o9eED38VQ3RMGtoqVQTDxfEXfGf34CJs5TPqsZcRlaXHXnlsWGcqLhjwLaTAtLA
lgFZqQrUl6w5efikY/sNhKyZ1It9kwqbiq4EL9eEs6IrfkQF8hbDtzeeP8RBKVtuqZGFNHo4qEXw
F7AUidH6BxS9z4khhNxBxw+b/Kg439pcNpOZZ9K17XZUhDsrNZVM+3mcPB94/yOahTAkfAHfBX9+
KO2tL9FcQU3PBolygXu7qyV8PzH3DEBwg/4u+6qDWUh4CwLCBDztKuPpXnTJx9pDBNG349ZvkU5A
IHbYW87Etu4LOhim/Dp9sUoRhcLrPYfb6rj+3H4eEoT9H/xXqs2ohywZcJB4Y0jfnnMV/SW0tf0g
LuKC8j6UQQYdcFatJAlDa5wshPb6eHaqlDz/vdiD24JJX9m0DSTSaqzyXwl4o3eUjwIXQ1FDiGOO
WjarrCB7OVr8ySb1bDDBI9RLvOUBwsHHgu/9E4awgmA0fb4dZ1zDvmoHeUaTOo3TD3Ia+IVDr4Q+
x/Wj5g/QX/e0zpasnggupwfmjyXipujcUgFZ/8y6+RY+/IDJbLZtc/HKMHtTF730BY2bzbIqYnPB
YIUHT3QJPbF2KyWz6xodG/F7BBk7ebP+ivDp9IpRXkbGDe3WUja46wlXCXHBYiBivu8D/BmEpb1o
SpaiEOyJVyX/gdtUngIxC5s+s2MHAFo8XMKgz4IzUhBld5jVbW3Ljr2wxXousNm6iWNhc9EK3EWM
lh74bD+FvZSRf9e/WmFGBQpb42q2KdnAS2RaR0M3zw/9hunMP4ALuOjpVzDLrs2OOk2XwcwI9UQX
BcxuAr8yf86JEWKXeo0afbJO3NfIeg68tHE8l/QrbuTqkDWOxAcGF6ydlwm0tvh7ajtf0Q38jDVr
E2IqJJYaawDDMIzvUb8sZp/fafGKvOFzcayv2IicHDUXGa0SYWV87dm1TZ1VFzMsM4KMVldOMucI
7bOVzF973KAzNUODf9Qmvhsk/axZ2tpMLzIuRjgMxIFNuQvCkoHVDJRnxc58zths6KJBOynnv522
mF+c8Bdq6OZG4hoclw73cXBTeGb/kZmt0/LMmiOhV04MNx20ihsWZ69S8+QtHZX1rXk8121mKNSQ
RwxDB+sktiP0LJXB3Ef+bAge4yU80XMNJ4mLE0K+a95i7/YakCPxyeiqV6CmbQSBPrgT7YiB5lns
B0aNMMJAEJGJAWV+/blcsSEgO4aagMDDUR6pWXInjHIYNPNTBPVHN36rdgOzyIxMKCLurjvc5Ndz
9EMyNazYMpF+NcKooM8L14XYpQ9ew1qKOu4HD2jivG3Fl8i68PLxZtGeAYWe8uB8y5hnhukis/8B
khx1SXn4In42aGuPgEatEoUFy0YdZ7xUoOPoIDHLEfs/l+UlPH8oRTnrmFkJVIvFIUzMITkE6Pv3
bcXO65GoxptxrFWeDa1QlGpQ+qaA7K319Yk8ZTwy5GKbCORBd5GtwvvyVHX/3ImSDHWySxgfQJbV
V0HAm9bd7OktznLd6mFdJ8c3071IQzoUK3VNiTLe8qcdyqsMHMo2mhtfdr2LZvDxhW5CT2a+SeZy
5zjnvZjFuCdZdEsb9QdGK+m4EYeaOUGocKBtxiDfVX1/bTvSYlzaErw8Kswjcrgm1JxzzjMEQqBQ
9qCj+srfCryRKWTQHOJB9A1iMSbBwdr4TR7Tm9BbNXhcyLl+VMNmjsiVoFmnnMZVw0SOt1QW4BGg
GT7Om6uiCdtx5sn+RtMzPORq/r78ob7FPbV806EY1L0AwQHZ6Efwhf8PGyll1T6JcBH81BdTYutQ
OJ/tNzss9zwMi4/MQwrC8L6zGcZImk7kmUHtUhQ2DXcj4/QcK/gVYqNtFgRQMS2S3OslpEhC8xTl
ABjsWsmJYb+JTVM2dPjGgEz+1a17Jmf13cK3AkLVqENtzJEDF3by4yeT9vAz53MqDjA1ix4ABMW8
b526757XLNBgGmFIuTbT7/BSzBbpLQnz7x5a0Z94oacx7NxmvGZ3f7hpdypv/4T2wegHCfyrYMIm
rthPdLJhRJajg4+goFeQ/Q6wjvMjR06knut0XLqxCU0WGg3aLqqiMw9MpR9VncydpQOw2tOKZJO6
xc/SnEPPf2gDzcJYgEkpl7uLYjmdv4prUZIIYw5jKhE74v2YT8tLj1zv2DClq9Li1MJi+G+Xx1aj
U/S/Jgc+WzFHBnZVfgJKc35bj5ndk/kQCvFfGCRS0AKj7l56+2tLjsEGj+3p9iPGqEr4lRYsg1p2
qjH0EFxX9LaRAgok4akgZ4NLjWwZGTPuzY06u+cZMhMYorwR9AMrzG5jIEmtEpowhQmxE570F7UQ
5Cuxbbbj+UwC0EkiWLcLvfeyR8m1bgNkuaTiAm7lVk24WygOK1cRHhunYJzCr2lMOgmvUWgRcTFM
TCkQIBnDvPUNYcDzIb8SLd8RyKYLeaFE4iTTE17o4OIxwbIh3fMkYAE6yB7FRBixiMKC5k2S7Vxd
TlB6jyDOwUppPBwH3+A/6O8MA9wTFC7LSycopzyY45027ESULL08b8aC75S6El9PfWxJCXfYjDwj
5Zjez3/Qg24wFziL8gn8qgI0ZlIRCr67Lh5S24ZSFhh/nCzpn61HwgbU9S48Ck3rE0DVQsH5/3ls
OzprRtpTq89/PvBfJY8hyQWGjeL3ApqBVi2bRFWXvIJS8BQ6EdVN/Gn5p+55t23EQ6FrYDm7L3OD
6y/bDlKm6TRQP9Hr17pA/+KtQS3ANKIIztlOiqMsN1fXN4yV+ZYb1X7vrJJFqmgO6L00OPOsH/FS
tJBCUU6hjplnRqtOuosri9Wg3cJXlV/KEc4qKf23C2B82yxQST17Hjb6bCkYaStTE79ci4tNfbxu
Ics+pyNf4JBe3gVUeVPTnh71sB0iqKVQKslqCO4cWeLy7dZDB2UKShTT+Q6PxRJhWM9cVcvz01+O
GGqD/GFcLIhvl0RroDJhCE1AlvsAetW1780nu3HAXwLcBrGE7rxUR0GnNoxv8677pPjyGagIFBGf
4S8198dPuDFhL4Q45exRAXwwJkWZTLEYWW4ZFIkx5+Lgqnu7a///9GF/l2Sthl7pD45ZDf4e/oLK
mTS/62oklH6wb51gNwT9UxtISzTJ7qr3SwrS6CJhOySD2m3DbWAgF50X9G5rtD1W0GCqI22hkGNl
fUe3yct2FdKcn0zRsP4mc8eQAgyXRsl0KgAAQq9DbsSTmlQY1eaIrHFE7s8MoDY9GX2i5K0qGOoy
T/HdKCSyjF5qSsAF5XumCIPZCAY9zQI542nD2J0uMESEQMZNZMv91gNCHfJrnVI3yOO1r+cA3s22
4kDoUNWq7Jf5pt5Kiu1W1p5Wqd0OcA97CpoovNUiEQ5BT56D5hqJ9lKXhPwIcIWd4gwhiLMEcUOj
xfsUAx0xE772TbCdya8wq0ofRM7wMPPPYyhJmUXYLC/bKvbKJuKay3UWk2rPZVk1mA4kaTJVEmx2
EgcvMR4zKYRv8JSB1cM/2A9glx8Iwfi+g66FjqrO5kzZkh7I9t6DCZqkFy+OVl2eXVyYh7gvRus6
RitcJBIXVX/BFlpFJQBaRyyHqohD0jLtevs5X1HAHEWFQyYmkPm0LjkL3rpSGnIqW0SfD1VEF4C5
j7+1UBoBHK9cRvXfSg+jmPMF6pieQhHzHzbg1Brbf85I8jiovGtzuDNfLVqiZUODvHKzYSM8eUJz
Hcd1vwMnh+SWMg1ny6efuGLZUVHbgzkAFy3kKfEEMvM41OVPtz6TKtvufeDQ0JR3bFJEKH+6zOOi
xcOMJ9smcvk4nQHq1vRoVYcQ0zZapG2kReFtjksV+HUIqIrhEHEJx8fFzf46bhuRCWcfpSwCXbhe
Wx9qU4X9YXQLscYnahPmlQk4UZyrqKprMfI+N2QB5+DmHZgh/C6IY2AC6lvfhlHEZCJRvW3l1szo
TgWEZV7aHtR6M4LQBuDCOCrqLhF1gCDVC68l2JRUzvOyiqkH2+GUge9rpPp85DVFz+12ZoGxLN+9
bqTMr4wvj+XiqvZ4bbw6U8dslWsqOnA14nDcNaKllrEBTEVA22/lTRBiuo2kUxmx7wiJB8aOBl+O
CDXyFZNqigPDgMBRak1qruIUPI3RWAbNJ2f5s93I2fvdDsudqJx2ZGrZmKTXkh8GYeC2UmPguI+0
2cKapg3RmJAaAOvkIGmg9B4Uq3NRO3VR5bvkF/Ucg7MCL0MaUlIIjjp9GRMAZA4gQUDH67cXwLuY
UceS1vLoUs3dl/tnNZGSj2yaX+xqwTcpTbWRlU5uQtk2jRtQqsQZa1uYPtvj23109+p6YjP/93pV
M5ZjzYjv9J++pKT6x+s6ZxzhtMjba4JrsvFwW2Z5fXR9KPTJ4whltJpbi6g796dqOpplqhUqE4nh
iAezckUqU0RiIKK17pmUfzWaVQP2eoMrFGnU6xE23zaTtl3eWf9Smrlbx9myLbwsb+oPyEsxbFxu
cMTqgolWvUZclZhnppuiNXDLwSOcz4Ih7gGq0j+BNlDw6nYmE40WTtgjnoWJaLw01/R6V9x8HZwV
8FnfH+l5/nT9eSFSK13BTh4JAt5P6OyKqJIfwYSbWVQucIYHXuwCGDvQYOkkWWqrC+nNJ14P4+Hh
gzuPGnzuw3chxyT5R6nT8ErHy5A1WeUfAbZT2HQbAO4zr0YXBJ3oho4x5Uwxus+SebYQHagmUhch
f2ynH39xmtuEyGSy3suf6VdyNpeZQQ8RIInzRofZp4oaAZrDtQi80tc3s1p62tj+rJNmgmVkXwe4
xS9teq+ZJLEC1xQ/B23wjxxq+oyytd+J0vSC3c0a+dQ02SS6Mw83D4cx8GI63jf1IjwqsSSwJyAW
rqQkrRzZDRXqHmzKDY2qj9EwGTT9k7fzePF2SDypARaDmqft7jC6ThDwCyK8IoBr4eOXNOlrXB7/
PigFi4YZRv0TjQ4OULUhKG0BnU4oOjRHbxiN7AZ6FpSZp2o/N+6KQqG+iNA+rdFyOGuOoKro25Sw
AR7UvOw4/j5SRJhbtr+LPd2fun8kz3uDWZRGxvh5Mehlf0aw4zKDdZT74L1QjeNtjRDWVpFtvmRa
264SH+t8NBxETGrFAa7ECMNRDravhv5EKPPMsEGsrgT5n7cCL32Hxvrz3Ago60QVvwNMAbWiOvhe
GlNg3qGUqeTUp/6bOe8Zn6Wc54GZz57kkcSpIeQPcGjTnaaRjgbc5eenrmVayziEDebGPvrlyydQ
X/coFF7L7HxfNXepirY+Jv07RY853E7ZbPo8cnp49Yg3Xgm2aM7fQjAXbSltUyGSjjYHneEidcsE
cpjtAMHQhdsEsWzFV3RbCXduuEqH1x2QHPMbm9USeb7drHi6ist0vAGb0hdH7S0DFaPBF8+L78qQ
wU54FGAtNMylhkq34mYbrTglnjthglBS+/FkDRatfXFkMBtiV+4BN4JiLONcQhP2vr5OFZsWr47a
LC0gFJwrHIwiDtQ8BKTZUcDwOCeN8YO3bsXwmJ9S9xbV7MB9/HNAflLe0WU1UoSCdiFs3eS+JDlq
spPITozswiLxxQX5PlaTOWxRHQnOHK9yX5AoIAC6Xi0RhPiQhlr4onjfRMYVxnSsip8SXGMn3zIR
UoogfB+oP9Z3eyq8FgUOeE8f3jgDrKmv9fJrwDdSetTPBwovKSI9kkKT6koqkKsJkYyypWOroVFy
DvDIzagSqlVdBrQ4E/6Wa53ct840eDP91aVaakesPXmNUrv3Kca+tfFePD6hhZKuNwIqNody7d7n
Qy8TC04YVLj/KcafZH8xan7zG+Xld6vcEn/5qvnzB4+vD5NWa2H5Ps+TMWKlqovrysPywUPnLXG4
3l0661/f9F59FCeQoZTsdnwq2A1zWo5fhPLYxVlOqWeNBxtzkrMGeOF+wuZJk/Ur9YpHSU8TB9Br
wbe884ez+X/7RUN+A1/hdPemeRKm+HW7kVwmQKqwfao6cAM9ShF/qLcl4Qh+WYQs7BJeEsypnIxQ
VYOpy3oATQJ//Dd2lOofsV2HjNLXkgDZxrnZjpBU90Ss9lCq4PaxplS6wM6cWwx4hMfw8ygzREDa
KwNdvK3+i19L2UElxvEFDC9k4lzjZN5m24nPTXdbNlZwM5dn6Qb0AgASqcmCFd5tep0bAwWqx3jP
3Wq0qUrO7ymZvsAaljc/sm/58s68XF9D/NMaKwY2ND/9FfnOizGu+AbUgCs+pbxGOuXyelpO3CzI
AyudsPsMEGl1crZskA7uQMH6cuTp3F36Fk9w3Cs/J3VlWpZOTUs69hZ6yB7ylg+4FPvigFwwICBb
+ZlsSJrOY5fSp2TYYvKSlnHGNbQxkdWiRFn2vLB+q496R11SrnYgDjKiOs5hV9d0+z4434jn6WqR
y6LpRYWpRJBr844Gy1C1r5NxAzlyyHB3Lpkba80LGhXCCLhZOTqFJ2ZoP0EMoGINF5XGcysH1pC8
lLH8dQ6L0T+F4fL9LeHVynojMaH44xO6BQ+wcren5OtSE3cDmkxjRbEAW1ikalJF41E2Hu0wThe6
Qp+ZtBz3eIrnHsdQ8IOfls/DkwW/My0Jfjbrvy1Wd9uD8xO962pFC90rqpiiKWpaH5t29smzFD/9
skxJv8y/yGJ8IJ5Lfz493w56oCjtN4a2GQoKWsZ71VP1JxsMOGwfFuuApwM/hdAHaVfVq+xwVVuN
o07oywD4tKu88wt42BBRhzurz3bbXp103v+KOEQheFenz5ErXj/Yz7d6zkk8PS78K3Vrl4Mo8UTl
MWeYUYWBru/j7lMLW8kGAPqnFyMU627W8WJaYW7RnF1j0EbYvEUnDwyWEGBegUdHTzTrj9hGAyxe
Isi95DfUB/jggm3AQhyElorIqaSNUAL/EqFnVyCkIHp3ifzs513+O7Iscr9ajY1E1uvzaKOK+dbu
YrPGd6h3ebi6wQ/SexeVVdAkxMzhy334Rw7MlCxLBSZtEX6tXaVP4PYqoFZLV2pqXcCMnkJbbT64
576zMpB9Luvne1SN4m/o6KfBLVuvhRhkhVBDKdSlHDAfIRaVxhpw2L9Q5b0kx1mPF/Wt4Ikdxt9H
KO4CszLfd8ui41bC//xa53qZnM3E/h7Mh/08hiCUc35+oZfphsXIdBgH+KXVfQA3lFC7XdWrDoUm
lUde494NfntW+n4GjXWot8AoYR+nJ9nAmW755BWxiYOEyNG4thB4HlAxL0DK91pkK+bEzabRNLhk
BDtfYOuROICqA/6pZHAJ/LdUnMYEYA8csn0M4dzgCqZim2EmYcgZQUItKpNIkrdw0bnJrb5gX3xq
Db1JhS1Bekq8MIDSwKIjocF0X1SEG80pl1FiLfsQO9w1YhV6sUHKmSzlJRxTh/0Wb8ee0j6bbLtp
B6IwhXUFfh3O98kLuw/rypdlok4OrW4u611lhZuaxNU5YDMYuFN6VxVOayxEfPyEEh6VdjreVSu5
cS9WbBANEqs4hA9jd3HCmHzmQUnIJbln3Cor6BqeH8dBLFrdOZSD3r3lZxRQ2ZXoBdpwc2kPFNOt
1YR6iX4/zPRUYii3FlqJZ7TzdmkU5PcJtQAqQ7I6+tq0Ls8oGME617RJ6FoDC1dXCBEE+WkiTWlx
m0mfj9E7T2bIIw49OaPnPt52jb2+C3lT7p4I8CpmPXUBN7mjrCoMyVB45T/2CKXGGEG+sqahJVVA
aL8ZPIaeHzF2GhsbMKHa1fq+AUR1kHO6mtiSqE4TgWykcpIMZ5RjYCTjQ+QkAyJKb3RNR5twCXGF
QKN5at47X2JyDChexeSqiN8kOdQJGY4jcwIQnSqDhprS4mzw8Zzo4Rgmp849mHHHLEnL87kvZt+3
dvQ+6Jnc4KRpWaQ8AQPJ5Q+/LxXdlpy8mjSQCwrv3d5ljHAIJIMprRLcVwitox/yM9hPQZXUBoK1
d/EyBV8es3Yx1JrJvj1pdYPayVwgvvMHW3hyk111633SX98kYKS7NrPdDBDl7KRnmfgU2JTtixZr
j+BIlfIgukdclPLSth0GHyCEo9yNoo+2USAuUr6jYZhODgaIXJ6kAUsU50PiEnf4s4Ku9JNUmkwM
vU1OKR66o32IL9Vz5s/EebbWOjXzYyKi8kZZLaZsxv0xlrfacXmElgO8k8gWyXtytbDiyDSbKIzT
yv1FyKmVM/NQsYghFyZjOsPy5sYA2jAICFg2PtK70jRH+h1nXD9EQLFSSxHlOVL31gSlpXUZARdC
iDqAR8fdwyql82boSWQuZBBql5Fz1hBdsMOliK1irFf90Lpc5UXYPee1PbLVVu38oZEhWtSnsgN0
RjlGPWPa4eqpK1hnyh0JSlxXeVKCas+iUog8mXi3dI/0d04xew3Y1ujYVMLaxYtfKMa17SnkIBy4
o4d9BZh1epszSvFU1T6e4/vU0AHrpl1GHoff0uaY5O6nc2Hv0xOQDh98mGMRL7K7AmM1MOQ8sPvN
bd+K5KbIyVprElCGPYxM3sDF4l0nySS8rQfTYXqJ1xaf4YBgmNLFj6mIDsnJu1ajtwUpLKVqw/6Y
oPIesrIn3B5K+mEZIgXG+rGOYiIGRU8NDbIJHHSkt2Pymjahml9JJU6aEO6eNt2+aiFUDot3Bygj
vBVds4BK2sI7Ga+7OS55H3Q8Ef5IwNs5x2ztu05l83/HpU3CCQSYl3NKSr2wEjs6WTLdWuWivJ3y
ECvyz5fQmXcG2ufPY6cCyhaWhiClIN9Os+qiqj5IFn/yz9+EmpzHqPL77ZI7tc8uKuLdVZb0MPUA
qLFp2nMLYo/gKha/IjnsENpi59O5KteOQt9X92h7BKafT/w1Au2ASyNKjH8Z9D81XaOmlRm2GP9y
prLsxNjHNsCwwFkicfNTNzG0q0wI0cNHDfpWKwIUKADWK/KpiiOXaPltGW60h+ptLm53wIO73R4Y
p3SQuqNGL9u73uilVy/L5ee4f+aQ3NxUHqjGZhD1h80vAUFqiOmuH0PPCzDYxgD1gf+HhGkAM1Dx
EgjUYi2QYF5ncXNy3blk6m3PFjIaspiDFVJSknvHPw2Un0VdrfajAKRWcWhgJLGdZXhMPF/OeGPR
58d7aAad7LruOvTBCYE/1cYSiWzNwUsSKUgp8jQxgdvTRqi5rSLofdwHyGuqNCbWD0g+M6SRjFHS
4aD/s2Ciury0+Fj/5kVEMsIy3J7aZWJH5JIjZRP/7FxxQygFGEmWmLw8gg1h+FKkfslg1h7bCGYA
MEopg123iu+7Vv0W/VBQcNT6yd28D37oAmgZcvhqpJWx88LI7VL6x89TaAqX3GPW8Z95fxhHJBQa
9EkGu2Gudi7Kwvcf/qiGNFa3hG1uCtK5F/q3syr/eOJo2By9vzWNRy6XAc5vQxJ1OImH+CPUze8v
I8OkBx0/DqvYvsYNAp4IJrO77VdeNkWn8ItG6BcRID5PchE6lbsfT7Gg4PSIXBIUYCMuswfNsIJN
mm0Ph2DpQieSIKsDPQW/5LMIrmNKX0u2CB7sIOb1msxkPKPuTwMpWB0lUI1e6rb3hCNxgzVEbmsA
aD6AVN0WGO4rJO1ZGlliX4s6sbO6Bs0zQ7ywKJo+YFPKVwD+4YqQGl48f3czB60CrJVr7bVGymuq
eVpfxAkQCdHiOry2Vi90PTlWz26ZFXUCNnCcUjJLknrhZd+y9fxLWCnc85dpyhNN1hGQT3SfRV/A
CAuohtsUKDM1fLwWFFhrUwaS1AOzdcBooTzBvAB0PglCUnbEQOaoUJGXtYz1kI2br2+xplwzOWin
k8xu7JvwUOFPnyesnHMqFVIKcDahvFGYc+L8pip+TAgF7Ae7FoMeV35qCy24PTh+YBOPh4Xl01OB
JYTECNWbR0uTLc71zLNkuWdOF59EnGL2SulEibpJB2rafzdlDTywMBZDownorNlsSg8uz6nwk1lj
9Fowmm5xZ8MsiYIMRgJP0O5EUwzItAf0p0I/4O0g1Dn20NqSNaaxPxdbGCTry6FfBXJYT35y0FzD
2+vexaCxk+Z9wCnb2FIfc43qiNpLXBjhraBPWh9NkrbeZvM3flO4K6MPQ2dwnAMKg2jluzG6sFLx
TY3nPhc2MxzaU27eQOVdvCdjo2RpLBI6QyAyb/SOdI+IlW44SD2bJFcZOaV8+SzG6FgEkMfyXvAD
bXNOcTOVVEcT72b5tG7SPMbl32hi2lH+9cSGTV2ctEhdif0+FtvP30kfSube1qm9E2zGh29G6QE2
s53ScanP2iOH+0k0l5sKe/hDxPYhsdSGKIPXTFsR0/J5RDMCEa1TotWM/IxQ+RtKEyK7V/cxTuRe
IbjGrEaKWwIef3RAoTBWOZleoSKEnuIyYu6itlF6MfTnme9G8CUU23NamnoD2fUc9YueAzzeCvMi
4dvZ88HDjE7DRw8GSqCJmJcgfEEahApl9kEz3djm+a8ME5Yt1NRYSs09Xs2RcY1A+6JqYD7TQBxJ
e8fc81SfVxYgP9onNj0gsx2vjrx+l9R92zSMBMsU58BWHTxnuqqzHcg8oYL1vlqz2qSvy5SH7JfU
rGJrTXwTdIa8nDLq54JQceMXDoH3Rk7Cg7OLGZYrcJgdytFuhqPPIeGi1eB3DqXNO7ZPhHZNUtv9
H4QdOUTbnv/iT0yMrI+NjwucmKC7eHTo63eJAHknISsWLUonIPG4k2wbK+Y6YbVEn1rTvYlpjJ3H
gZNMhjo7ToE1gBUf1ckl81eCqhMgWeC2GDe6euT6X4LBwNjp/NpYI1wNbHSCQWgH1rwsdWCS85FQ
KnK2k2dHLdLzcPnmgyTTyQXobj4Si9cwiQxGWvbzmQTpIZbhJf8VrZKOzofcvF1r4wiSbUv3dFST
mqLDoxJQfMDS/NrLuztDHNyAp/aQPwIzVWLvLiVnH7prFDQZLGwFJN96R82hmu812ihsxexON3il
f7EvozRx95STZkIhVAcnAUa55kPgatRa7cqWCCzbxp4ecvjMlwOirpt4pfsmhYC3GCnSbbxR8/mX
yE55GBo7UHWj8hqHEpF+mfelH1kUl9tYpTcJ6D0/xHYf37AH2vOQ0UWjktR7FBZJgSPgrDK/kq21
Sbl/HsjjARrwjRVllGArK4iQwd/OBemYpiztE4JF55EOo0OZWqalV2amQKH8fJQiZx9Mca1qbHoE
hXRcQldpGUBYBMxePuixZwkZpBQCFQRZaMC8dZ24HHW/97rbf7LBC259ngXbqsz9HzN8q9oQTfwi
hUrcvzR3YKAvezovDj6uSNDKqHkxqKltVo59nU9ZkiLrpiUVuwgGnjs78EH2wmt1/zbRt66Pqojg
MRa/w97AsjIOOGC9A+xlGLZz4XZR5hB8B5CY+Auneqj5JRINxlLi41BSnsZvWAQcBOdLXEe03lm9
F5Nw5RaNJzkYveip9d2iIEDRt8UahFtgKkslRfCiIExRg3RJfy6ey2YNhPDJYRd0TqLKAmVgyfIb
58gBdv5q9Xj8F36ZBJge+//OLe4UFmfZe6qhI//Hk2qqQkcH1344g4QLseba8BMQS8ihK6WwTN/N
ozNHowNsSGERjcbCjm+++BuQeNMVa01RvnyidBPF1l/I5hTQ07EUieq84vs9zG81XNVSRiW1ErMe
yNWsQPFZYTcw9EELHcNHfZeZI/U8ElmJxefIxEB/14HithkAaMqQs7i/fNTPIPt9/mrGDT9lCfxb
598GpI2TWiLKvLVO8DDJ9OlgEHw2P8cK7yjG7pYJnfgSy1KXTmisttW/2e5ijM6DnrQ9DZkUwlh8
p06lEGLJolk9xJYBSnOGJS5MwU6C9mhH3lasyaD3DlD9CDRrOBx5goRPcZFyKz6eEKnmzdFzCPTs
4zRglaXCyDLmOxK3puBSrfzMZGxcZc5xWExo25TeP8EOflSqbC/mcLhGmA6NLVuQi7IwZUDWFElz
BiBMgNdDkYBFbGOkHLXBGLCXpyMubOc2Q6C6ZbexLJaiuqsjapLiNh7OxWYg/C9jhb5Y6Gnt5rjF
Phinbfp2nh4ee9i0MNKHVHPMT5vE1nEnnNDkK/Yrt+HjtpIyt8WZ38EyIO7eFuE6VVYGmvE3u+Yq
mEVEP0Ats2KuFC8cU1U8GDSAgYiEANoIKaNxcdbfDiCH+PAomuV5wBKalGThQUqCWl/iZahhjV8f
JVPc7CVd9eW+pY+uJZFMUMvKJvzfjxYOPItCnlV9tsL29NT0ctQNfgjp1zD4OUW6t2V2EOspN4JX
FpGzIEYdCK/qCXNpCDv/MKqlhUDJ09Mi9ESvDQynvj1MufUh0YMFrVzwINwEjb+Dud/1tiskQ1kt
NptLVzarnFZ5BiOd564AMT6CjdhM1VVnXRKI29u/wMYT7vMmXzeMc7snyCjUWFVn8k9Sv3d+Kkvm
gIP0u4mBnVIyjZZa6UTRMr4jE4NNgitWMmVBxdGQD/RyunWQbPV+pg7bBSB5zHPdcOoL/Bjnenzl
mxqHUKrnNDAaRVtuasfsGC0dhtRIyJee0CyeMSLmOaDw4TYQQ/uGOMaqm6dvCm1gESxLzvXEgFzB
TQ3e6vHfQxn286sv9zBQ0sa7WHKu8I6OHyb4sujKSTZhJOKh0u9K5te8MAeZaBIXxnacXontJW5N
niKrPK+UW3J1GXOmhmKFgiHGo69/8gWx2hMc49wdDjdlwVSoTNXNoEqLVn24DyF5tU6S9lrPougr
2u6C5c4oih11SRHE4zxfoNqyV/l0Khrvqsu4T6icbaWkH4OklacXlAfRjW6oclBma74K1+mEbjPp
3Qr3WVtsuy/eBjJGLaYbx3UZFDCkWDg4jCBrUzfq1tALHUypn9oHqtnZVrSZ77CqguU2LmtHM3yc
KuWPqHz02kyYVSXRBPC2LJm4Bd+jJEFXR7bKQSierMxz4EVKfkbFE3dQZStKQiOu2HuCTh8IZPl/
Ei13CsJ5vMKgaYJJawbZrKAKUNazZ9rMV3e+BaIT4xEIokOW0QYfcuLIOTlXSONXySKAQ8uei21N
UWIlv2ZQ90ZuXhiPoeeGtnahA/O/hx3TnL8s5MFwKOhUMCRPNc7Zt57mgoInRoZ0EM+Zn/Cf/q3W
7eaml2toc7vUJ+1c5FRsLuS8nzu4+lfxKPuqp7Y57ZjVyH3DQO9x6MQfxYzPntc24u0aUzYftjSG
qFnILaqnhvMzoF28uKUc6Op8nyhMHHunC2TZpq6HKyHQSGElRW6mkT9zcoHAGEXDx0pr7rqqsaAF
m7ArPdHQAQijHPx/+Bz+M0zwmFgDfdHUNmQsxRk6Gu2cX24+poD174KCnKgKxZzVBBOpGjGSPS5z
XrgTrKROOVU1XFAdPj9HEuHw5xVeM0w/OnrKL5xCwJ1uGDxJ0KjEGh2wM1HtS7eZPsmYFLIgI63B
pQS/zSp6v9VM7jfQ/UzmCKOLVjKPQUXupRSFzl1YhT4jCZpk6Tg9+iV2TgiMX8o6u459/qKg6twq
YznSxjSg1NPW62bBiESp9Gw2+WdhWOMOokN9oRn/gcQaEFa4rgdPtrnnU8aDwfZgqDkwjFmkXw2e
Qa3rd7QYHS5vc1F4Ca74G7RSMQ8EFdrFUavHjbQjEj+BKdpmDgP5PXQobKXadM0lGFHVGg/FlUos
KwZGiEm05/H9451LBjmzX90fbFdlNZfYHMguw2JgqPVlSibbpYyXTIlhRpRooAFTyOpAHfBwfEbe
JnaZDyjX1zqnpem0OtZIuH7iCPemlFLGbB9LFFQK5ni2H3qDLhczyG2xUT8r5J+d2TOwq2j/+r9b
Vbdb5dShBkQhuzuIOPg/Ag+enc+jU9PJnBOZswjs9F13TYzqfvas6oTC3w1d1nn/vl0O2dOGjE0J
/6ThwWxgELQV7zW+OQ+BtZOAR2KN95q8YWSjHKvt9EIU8dOPU0hb57qEhKs1WHWCHCsyBnvnQPYd
HLfXCinhxpaS6kgeYo/C6Pk8fN2xvTK//vYe5b4Wa3sGtWzzxO8riw81nX1ar6DFHCmpAo9XRqpR
3nHiqgxHmfE5Xa6jgFETyaPpAYodig4S986vKqWIB/J2fDs3DT/ldN6JChl0AxlaBXiA3GdMI6t7
Lyptg39/FewEm+27TOO0FrZIIChxaN5s7FAH0Jfh+mak/gWL2j6n4kILhSNU8r2xwVFpcT1xBBPE
EHnvxSE7W2XHDalTShnMjd5fSQKZwWn/Sy3oaoj6acPzU6EvtfzZrmn6iLsqObBp8ExzgP/8i8ON
ZM/OkA6uQRK+zZShnNBuc8IJL1sJHo8rjhKCBppIlGFR516r1NVhfJRoUd80cwlq1LjPWyyCiDw9
/O8k+7NITICI91aJ7k8tnvh9I0nqFm81nV13rfB9XFD/hYnSBM7u7o8W14DimSz8Cjf6mwx0h5dv
YMXGNneAPUvWhm3OAdO4lruNmnyfin7XiuqpZzim1T7coIFOrs6HAXN2nb13fbY9kuOW48V4DWlI
LypcJtNNvufTtkR22+0h/ZcNmwYZKrxxMz7RwMTGVPiKD12pWUqB8/YFdilejPKasLdWcGj9i8rS
lq/7Jqn5kvzrxe2n3HrTIA1XDlXBkJzVHXYFBJSKWDjHCRSPzLpiWk9UedFTu1pBP1vjBXxPkuhm
zWcBQ0HUgwMzbOcH8ejzorDKTQgZaJ9ypNNLTElfF9ScjriIlW/N4LFhWp1Iz7oEt7FdtBs1XrJv
gtMcMPzyx6GwwwuOPbFsmjDHXhGtpZmAjQtKZhuuZXdYh3GZnvTrt5fEA8mATJMY0+p/9GyGZS2o
l6Oe898wSr/2G+WeUfjcsPy3LJlqHDjSPDcLYK+CZE+SaGsNOidylb14HHwZJgCDC+9p351aW2Mb
1cMc11ty+67MGUygs5bKUROO5vEAVDNN1cGyaPXTTYe1jpuNL2v3QRo5uhTmnlyknv4ObPFkBJnu
P8T9exf4wb/SD0ZAWqV7212kS0e1QT/vSGX508XUITvgFt6e3W9Yad0Pom5xx1kwKfnHXrJ5pRix
w7tY5LR+V8fBvXB4UDPa1vayjOZLxCSEJcM0NILc46WmC2AuoalEi6uyjdsqHazOoZOqvSstIPFJ
1d60b1ow7K4DsFQwtDkydiTcCKc0L7EBNHOPI8BRu6r0Vq+CO5hVnv/geS8tmFfCtic2qUsoK0il
SwF3YS0bDLvIcjBPPQgu2FDOxppWRoG94N47fpIOkSJC9iz8Il4nwVBVhuF2ssbertxV2KqpXibo
gG6/NkkSUvIonoBmav517xLBXj8ArhR82EhYEW5OPlevYK8DUR29tRk2UbSStl14+nZpJu4YzzPM
bWQlcMC7N6XThROfcX0Xqa7j72UY2/OyQbZO25GB2VcWmnbFYQvBZ3TDMfy+mNQCxEs+fCmhSHX/
JJgtUN28zkdjcbG2zhK/P+oVB0jyfgrABAr+7oxBsWBJySQJvSPpxHLiebJZfvClBoyDm5Cqukb+
6Jqif9KYoOALVLo20NVRT2uJ3cMBf7Vtk5+uEvFyr1oOd9lpr/FvgWpynhFiqc8keL8f7iTApHpA
ObMHiSfMajsGV2JagSYlaf+A3UPUNdodF0oflfpK6TKfjwcu0r4vN60BqwRK5TZ0Vo+hahwu8h5a
MCaOjNlOIo/HF33gooAqlR3LulNVOa+Dw86FxnEQwDKyO3TRHlzLuUuiXPvkT9hYRvyzoaquGQ9U
rN5NQBPKTO4GPNkmmqy8IlzcrHF096bh0vRbeZGpIhlsSnC2Em9MseF8zxlL8BHuw1/FNRNg/+nL
b7YNiILc5i9bCrfzwjK3bFwflsLA/7OKLeUlpJVrs7ZwyjijSIRTzkdG6kts/uP4+YSXyGfINRGf
63bIXuXtinlbxCJmgGbIDHmWQTiEeWNKEgBEqSi0tTpsZ3YKeBRDaWqGv2+tw3QHsOpUI+s4+olQ
BV69fZtlZjRR/Lt8k5y51Hi/ZYL2mGjnOMdH8x6QwNCXNVL4HBET08RaYMpa8buF/4zM5YUV+hOe
+GMt2gBI4Dwzg+6D84EQDqsHuU0H+bz+UhLSXbPAHam6yjugeEua9uk/iq1mxXiR6vwDZlvhaueH
m8N/LJAdd66abvTfzs0JR2GpxLFWyVSarISIlY8/sherEn34YFk3whtesiDdfnVyC9OdgISbvvVi
PKLLgtG2xWSrRwMiOOKhbOSkDDQICWfYF+Ntsn1Kjv6Sz0t/YIWvvqADD8IYe00XJwWJkW6/6pi4
9XigFTLXZDb5NnYA4n+YZNHmhJOa5ezhEf/qPhSgXnbZqyOOCSf/OnFZYDqHB9YAkmZSDBGT9WfR
TYz20NdOyzAnG8LV1UBrmBKh/BaUblwiO4rRAJfARDf8rMZyfolLU+GH6mtSS8ScTk3wuwsVqZnI
nWaM6Mlzo5d8Hg80p3W/dtSNrPTNnqBm3be83c0TNxY862igujo48auTtpmN5FcHOtRHb+DZINBf
yTy66e/CkBwVeg46/4O5a929iSCSbZFXe1EC/tMdWPZyBJPcCFskfM7CkkDkU9aeh5/3BW60xTox
xxzZjL7L8XCqjnjCw1ggNBCCPgTgZcmPOm/AJ1sPZVfcE7gzDXrOT5SVMGT5E/5j7hG2/fsoPVoj
JFT6kk2eAwmvCy/bBW1tUtNPoYz46ZBpVrmc7oBuD52z9Lc4IGSS3HmImCVtL4CE3sA2Fs+EvYYb
riZ66+ln+eqGbzz91QdjhQ8YONXzqC+Rhs36J6W2ngtzPbKDmqJ8fmv9A0xwgMZwUUe7FL/1pt95
xV9XnZvWbqGBgfh9GfV8yUPfBxfpoQTeWuGsysmSNBO40FCwECf5ULuzZIPPkpkQmzC8KDzJBpnA
2s863nbQ8igVIycSP/WhCalFgb+CkSRkWburjxb0TN+VD7qO5sprwhtJ7hhY1gBtEeAsEgLFLW19
jo/GxIyh6VPjhKCJqdU5qTossc0Ry7EEr796/9uEuavEFn01Je78muAcTLzxA0NYp6wDd3dHCxeO
gDrTfXoN9z7ioM8WCjaOwYN6wJqUkQ4vsWUg2aTFX7qcuBkT3xYUKuLafPsFvlwLzVJgeSECQ202
kbDobGDz+7OIOWjd+ZEqUb0jKyvkHLezQrX2Dcqik75KU5pJswI8bNizNRaS4r5Ypg2QntUUkyS1
eDS3MvYs3OvMN0UkUNLloACw50eT/eAcFmALrpKjUD1fuKdHQeqq1XfLXQ+je/2URC8UPUoujOhY
XZgkVP7XhOdiLDyUAeyYkzvLwTNw46LJyhMFSZ1zRzzFF1iBnL0HGm3ma2xv3O3MXjSqwNhjV75Y
9gSZBMgdncwo/KnKAFd+xcypFrB850FYBgGsvV0J3qkls/4pBXI/p0/wqEE1ZJL6N5EYbeL1OYSc
ED3JFQVkVbHyuYEdq2x93IC/N1MvoJisfIxjfHFg7TBR+6axVGRL6zD7tZtAEoGBY4DDTKYrmyE5
p3mOuPx1oRBd2s3bRAtBP/bYbJdeA/0VbXsiWQJEvLMALH+rMjOvl4RYuwYIqYoVeI4gIsP8yXHr
Safnv8PyJATeR8ggIzl68Q05V667Yz6E6BMeKM20DNKqX8ttlPGYVQeYJL5Rpxc9Jb0ugia3bDOx
+gt9ErGfsyJUgUxW1XbA9zTioppn0opDfM+kSc7EBQmNRqEicrI5WWuW+hyvuE4ZvouYU7cs4Y9f
JBiNrapVwulFI95ailMBOHZeVTEDqdzsXAu6VkwtIkXbgHGar3qDexPbWJxEzRUKAiw8hV11x27v
+FBaivIr3tW8tWdxKndO+nHvCHmY08FYwnVKOu8L56vjdrSqWf7Ng4+Ah03+pT6BF8TFBAuADsfd
kqFhSZbw+HJ3OanHpXNrhbEdXUobjCrakU3tRRvon3g0lMgTnC3AMQcyzuHbDr6JiYrRqmIhWtR1
NGnQzeDUICIIWdyCuhgKkFTRONlazHwj6Phv1QEZb3OgGJ/p/uLhlR6RBrwIy/rdAE6dZA1GvtT7
VRJIBgQ9vplZij85vBDMmHPfzTzTgaS1ci/eHBzNUMgO10PdPj4/eRSUF+ZcgCYKinqtdg6smCqr
wtMIN0kvz9PLCGiI50WfzK8rWChnRIJbA8zBtQjqbukUelABjFfjIcANBFuONGIKCeeiVgubwBtk
o/2/0f/LhCC7MTvJxcEBVfRQC+bx7nRAqOV0/pUH5lcSRqxvASsa4P7FTPbFpzXJrfHVKe0PmOIS
rfIc/RgYUSha0qha3UsyOZyg0hrsc7Y+zjswRnJ14W5QDt7p62HgPprI+zgkHUotuWf/LKP8uDCu
pPsBVHMECvvYpTebvINKvr3OkmXGCpSK2GMNXQwnz5gZY65+ycUtNFpZgz0DCMhL78n98y/akAUK
FzssdnBrzMgYaWmabmDY2iE8gkTz3hwGldUlC++yXuxOEs0dRSqP2HHkqEaDlFi4eXJDyTuZKFDS
HmeI8mNkTpYtWzcHBQv0+emLxlFmx+UqbIKtlv7LgL77RWvrQqNZ2Bjk5woJz5+CAed4Exy7V86J
A+W4tGxQEIF+3cNVQCNYSvS3V+1RcpnqL+SGcTSYa3e3eH7pWsYqPWkJVk8J9jKRy8k1ZGap9YH/
im7lOD/9U93bNeyIjXMrZtfoHQB9wdsH71GfOSK28DAghlB5Ui4vQuanlZCwqTtbkiwRxtA0Zvw6
gaXSpW5fbs3otkftaeFozvd5kLmoij6U6sKNkYaAjUeniUDBipW21J6fKQhIaHUvTgDdJZxVZNf9
qzqAGdHxDK1Az5OyTlCxW0jKeqRYdTHiaCM/f8DAJ4IwJpnWHMOFetkibLmJooS7+YkhCKy9Vus1
ad+4E+7ftVRpxY69YN08JT5B17dKlfdTj37Sd4ukY5OMWWS9JnS/JlX3QJEuVCOCh85CEF2g1hPR
+zfBOP2GR+Vj4cPdtqsP/W5YE8had7t2r8FCqgqVmeDoZKWKjSh3Yh1f6PiXqjqsEQQQkuEGIXCN
LFJygFX7QnCpwLGXEPgF7DGaZEcQb1IMxkbR2VBQYgzybc99lKu6HX3sExlZ1VLXEzBMRdzYKoj/
pg3znyV+phRQAqRGiW/B3u50KnCFqpJVzL9YtBLoBUmZq3GnNNPP31uPWgv/417U/pMkTjFs4BNY
Hnq5/gpKeY3//JeYPEr9/qzBuq3V4JuYTrTqcjckSziL8NKvqvX39mW7VVW+KAQGO33RiWchL/ye
SpF4hbD3U65HtOVsvmRESzAiIAMWe6xspkhANlnbtDiMyMg0QMuZvXt5a0J0OnGoBe97uOIRgQTz
gmRT0Ft/xnkZhK+B++GhtX7UXrmGLyV52AIWrE3VlRgga3sw4um1Y1F3ZZmdae8vHO5VTECMTsUR
alh8RlW5zxFGeowSFrQX+Fh3Qgn/LqlpWbL0t8+rxMVpzHPl7X8VCC3Inj4YNBAp9bh+bA2nVq7H
pGfS1ZdHzT8e19R052QJ6u0PyLkHUpyBP2Jy+2vHD6pCyQ4C91K7IidGMI2pOpV4bj2QXplsFMIA
aCrJk8TLLmG54QL24Phb3e76AcT9M6l0UhNWCMvZRiSy9n0ENJnlcQyvXhkE5QEmaF+8UQGVfPxa
WdoskJetV7pqiLl8sWBUhjMSI79DpowyLa8tNdzONN54sllMoN4f68BmtQg9a31LhFLxlNRyXMpq
kmCIWqPe9ACYi14p96+yqCImWwYVSzxelEoKfayzTGvNon1rad1VnRTkiNp0nVhRWm54XwOgLcgE
1n5vUsMy4iyffUIAniLpSSVehPd4wElMG21Mu+82PZ7i114zXPbr1MHPZE6a4W0vrdk+v4qsDdr6
CNdh2swxUyvuwoYsGvaXIDEuw5S8qQI3W1wAYT3v42KEc8GBuZkPjbJtIUIgAeaU4EgMXogPeYNE
gLLdcbdrluL007D5jPgqHSH3KgUHQYwgF0W1BQuhN5c3rMGcInqnSNvCZ2CPUSSK2NwKpcDTyZfn
8PGyqddWl+ZJBukOqpWnKULliwNUB5hqINf9DKsJeBW10o8fsFghzgp8c+Eaa2aCjKfB7SkpcZeA
wiQxZAxJjZDnan7ploan/T8FuZ12/X/IzUDEqx+FlGSGefMDNneoCA9uVKNcyYCpZ6N86fNpLm6A
1OOJ3W7SgkliiyC9RMx+QkF5kFbfJLUevaSsArX/OIVkuCwzNTB5Qn8Sda/ksC+ddAoja3+4MCgX
/N3mi1m6g4UZbcZP76NWCeG2SbuSj5R0+5l8V9meNtCvbYoZpoBsDAPyTSNL5Oum60RMIk0L0dpe
8HOz4nCF8977/N31OJaJ7kUWJjDP5EhomV0QDH1yV9fUlylvHUS6i21XunKs6v+/J4/5FPsANRHt
F6li4Qk+Xza66fV8KK5C5NfO4zyG6juAcBKq86Zvt1ufQNAQLfp6AcgzZlMv2HOsWNWM1+JY4J0w
Q1+cX6VwhQLTEBLHjcR8B1ZdiFny+gn4EN+Vz+aVnSl+sYfAOSWqrcV2xKj3dvQWuRNbczc/3rDO
tyHiCDg0Qmyi0XI9Jlw9LbGjuZJNj/LsS667v/rGfpCFNFSYW9U38My1XPtldyht2eXZxxld3aWO
m2mNxDtxh8Yn76HcvuTa8v4T5LqrYwymIYPlwDTJYJ1ZIuBjL4Mm5h69LpelratkM8h1DGOpdmru
cbppT1RbTv/bk6HZ1dvLUYW7xJhvsZ/D4u+Tl5RmSoLLc0YIkPudfN3A5H8yXUYqR69DTlxgxbOw
1VJD6COtr3eAXbTyX0MJjqIXdnObSEyimQC6WNmInq0Yjj0xB5ISm/daw9v0u8T8ax8qqRCE+pK+
bNF2Ev0SPd0egW/O8ezOrM0SNNG/M8zMjRmJM08Bk0l5+vSjubL6S4LZFW21oOyeDVHRa2V8Q3LR
lCTG6A5F1HnFJSSfPes24wemtJKT3BIXO8Vtmmv/WEQHqWyy2rqTKCrPr/EcaiTvW85Utq1SgBSx
kD7OgeRiAzofqFYr8hxaeu3BHXt0mMsmmHUnbsSE8NMOdHHL+bd6itC45T/RHhLN2105Ir5l71So
C8tpuuLOsun6SPtbX9ULN85HbwDt+sQOU9pvsCFhwS9iF82935BodppgLACUtJczcP8CYTeNXhGt
vMiwEVTi7LUUZfHOjfrhu7HaENgEZRuy+SgxpRP098RX8nYps4GkA+pRiZI1/mgiJaMW2o0pGHWW
R3txdfbP6vqVrikIrwq0JVDm0q1bGJtb3zdIvFM+G3Nki3eIJ1olKSWBER1wAY1V9LUH0jJHWET/
98GmLnEKfDu2t8q+6z/WIjRxrZktWjJQSAtLyIP4aft69mKSGj/9PBj6Ri7Fhl+r9ZsSsloV+e+g
FFWtmjPel+D8yp9jiGkNyHVf7EN9JfB917VvQ1GV6NXSYSUcYp0mhG/PkPpWZ8VbjghfcvKi5t9M
D4jbA2KsvYsmfGh94PZi+qRCmOJs5kKYVxl5l71ENi5hqdoW63NnTbJXdlq4OgshwYW1wmfObcSJ
MWNrZ474vY12NL7LSfoPpwSa4WpVhLzYhZ706yHlMUR4+LUaCDn8sJSF5bgNc/XGubAl5ZqsyYuU
9MW+Ts4W6E5ij0WASZe+wqyk81A81qL+c/D+RIU0nnt+gV0ogNIWAO6fo3yBomCwqNzW3sZPgZQi
RLk/F/mdMqL3iTx8r1uIqVZzVETfEn4BKpg9Obvv1e1u3hqcht55oH4yopgzlVvLxokW1kWqF+vT
r8bByLkDhKd12ngb0eVXQpY/rxj5chK8R1Vvjv46M5MzICBsPFedQl6ufW5uM2L9noWVNsO9rLlr
yE7GA3UpgVUzEYkP4R+CYYhZPUrmX5ONeUQux8AJX5u3BWPp1ebbYNp9bPycAVvWctcYKb4q5Uyg
mvwhzlUp0jG456jU1kg5VUWupYoV3iQ6+cULxpOaOCDnxemY66jcX2FRSV0uHrvCb5hoalkV6FRg
tV4sqXa1Z2Vv4XYW9haMb7yYkDw14zDQvHyDjjp9jYOKqGZo8GQxkOBinK/BKAC5zDFDHxSbxXga
fnkDyL8vPeWSwQ4wxufBrrfMJC5xQVbBQrmqgu0vn5GRyuandIWIiPSrKO7ZPzVeEiD1RP/DiQzQ
ce/0n7CgMbtFW7HYQDBD1DPpRX3KVSwfaXH299RG6Mjd/KYw0vsOxuN4JKAwU5kboh11gTY4TfF+
4aR7aJXf0Tv2vLXyjEkMW0qqRBQ3cbPpQ6VZOMBPlEpVZH5qDV+Ho2vMF69+GHNhUiO/QRUQx6dD
xppMLtBjKml4FC01aqeJta7jBuIxY8y7Qi1nhKfzyU2BuqgJrx33lPDymkQDMjH5D/2gRke9ah1R
P2PTFhda8+o61F5mPR8KPKnMxyPLmoglLKd9OX9X9eDQcXtTB+IfGEWw4Ybnv8yLtFmjjku4eBOd
sUlmD7wZsyp7kB8CG1jboUQuaSjuGT7BWEbhB5VKUjgn1aMGomnIN9sB9e/IW1N4hHaJHakokzu+
eHn2ImNtHKt2L3QkLNBX2qhxQz0nX5BA+538LQXinGKvmEVYw1nTqbm1Bzi4mxFDQezVs14NSduV
sbkirkw1agU8fnxctber9qiWq23roZlngnBzFgnlB2p0NFGyKe9fH9EAg5RUlyzmfmfvAuIFjNXi
69nXk+jwlh76/2vt780+nvss1TF9YOaVLoNvcssBNcNsxNh3xzUZ1HcVULXxnKtUfVuGZU4O8S9e
WO3JxiYjG+kLlhfDo0c5cS+S7Xm2vjJ7ASKnzRrcwbZbavCKDO7bkLmpOMsjuuzgANuqGRygzzHj
rZ6HcxUiiIJF5ZXIllAfbQmDVLdBhIImps22zQzU4A+8C0hUZCG/0hbvrOaGIaxtIk5UclyJ4mFH
40iXXliNicFiqDseSuF0gVemcQPa+MJMGkZbqAH+VPOJ2NNleyiDCqr6ddY6cnp1uSUJ7adnXXb0
9XXmmisPK9T5Ego2+ob6yGXHRva6G6xH3xLlcYL9uvJmInqKwYGcK9NnqG8bOfybBPqZqpumEGwo
L1sxyx3kYIua8LDzJnwajSgPF9e0TyQJ9gTojj0vzpqzK7ClX/SmyXXERV/Rc9Ru9mRwR2yF+rpZ
krD4zp5ptzVBRdC7WFlgkY9sWhwGW6cFqK6O7cfg2tVVAtF3SZzfS8kjF6xDzlF7GqySgl8gudHZ
ObuKpAA1c8xfHIlfv4/EPai5DJIFbqtKa+BfngoG4OzGipvTvrZvcx4YSXhTn6ZIFYeA9cyWtn0D
4jd1OwvpjmvzFmjTzS6NbOiHVzTRnfZBAb7mdUVhX5AB+eiU1MLb9odbLRTcuWBzJaxwph/5tIv1
RW4NPtfrQXNzfSAGyzvIMWY/mOQTic+4qH4E/LSHSZLvLzAQOMpDaItFKVFty9txqQFVWc1+dKg3
t/TS1Q01WDBkv8HlGyhCfzfIRV+eey4vBcNCbfV4O+Xf+n06gl5anUtKvklvqTLO/0GKfnP6ImLR
t8uaHD/MWrO0gD4YHHZR5QFjUVCrT5KGdscNZ2iHfy6LZ9YKxUQtuJxLBYDagTdJafvzZqbo/ZyS
xqnWoay89GvG7D3MScMHoVB6wwnQLIo0FFckCzabJIR0f0v1gGtMfUOOqbh+8mTpnOX8mXEZ8Nfk
UJTdTwheq+AG0AebL9fDjZoUewAhUVb+zInCGihi2sS1Vyx1JBgl6lMMjWJtxtt6yLmrDOBr39dt
QqC1T4Hk0Pc15vZcVzaJTrJ34NNNzXJ08mjPKP0Y75zTJi0VshrsOgmUOQGe8m+SZg88BnUYwFVk
fZeZ+8C/9FgosrNl1MJ2jr5ARKQAjD3Z0LnscWYrL/bsLrDXOX6t1XSN0N9rlhwU2Dq+4h7cHgAr
VsvaI5Mt5kPMTxddMmAaX1xpNPELID5BURTHNGFk/POyExW37p1eVcAkKSiGADlXkJsJVBZlg4Mc
xUbrL/HA745B5dFBrrdhcbmLKYdpNVKPw8fMTmWi65JdZ0GUQ1EHgxSMTk/WybiQ8OSxigXP7YGm
fn+sP95Sm6zL/V+hinUbX11omQdCYISuYMEvWubkMLjEoRjIe+07J9kPxfotA61ETlSoAEArlNXh
AEJRV685+A24sjQqorrhte6nAcTUBouhxW1RA5G94DDK7eUlltznKYTCOGuofWglcLMD9YAVNlXj
bzecEwapdpXRAzQ3pMtgVMUEVzfx8wpf+0SGh5acu2coeO7U8BsrXpWJgsz8XdxShBbY6TsvYuUN
/aAmzse0kmTEFWCbbU/wLBTRYnN7DH0moGW4Jq4m+hUaQeZj80lFRKP4ACZ+zqy8o1BpSMlG7PPy
B0j7cCYcXXOzgeBwNi/9XklkvEajP5BvTp8oAZlJzkkiwhQKsPLaRaKGavazIf4A/UXW6r3zQxFt
5tMYMs2gEqYxVoOb17J3HH6+mbWgKbuNum5rVhzkJMIhsV+xzofgmXbvjIiTXGVBSXrA9wi1lFA/
FrauWzGyI0VS7BzoKJeLMMtuIbJRsMy6uNFujbB5HIA68oig5ocAUj1GEs8TbKtBXOtYge2JAlPG
XjVc3sUdWcDcygefCmK8g9bJn8pINxftxBCAr9BSR0Dfy/0hgv/zZRKODYeg8XtfgswZtpoSNlaO
goT6BOnmhO7tRPihwEnclSasz75vBMsYLZJKvnTUPUrYUfwDbcFISqrMAkgBEYUFaYRRiMZ2WHbs
aR5PRSSJGVt5DjNPLSWYggYwgDhtqkQJPA+uszoLwuC4Wb00hCXzRj9yFpkjkktXjF1rlysF0TD1
zE586KQngPmVnUw/7g/07AbiHyRZcN7Imn9oDtLFxDXC/IgasR0IYQUV+7WHHFujd+eiK8VYnNML
azQ7TbFe0S86k0z9IyARXGkQQ/C1VpN3rbBTEkHU9e+9WQzkTfQP6RkPUCBlsCL5HkNtkUwC15mL
1pONWpPhB+nQwSSopGJfcbk3IgpPSAOtmRw5/cPmvD/ivNyEu3A0HNLC9z8Sd40W7AXUC/muT6+I
1g74/wUIcoseSwxtZ4JGvZldBaG2OjWzDKI4DIEX2yWPuoCkveISvT/FZdQgGYdLsIagx23WDpnH
41pOrx4KpuvlbYd0vaNMykhrCBfpQ/He+3GNWkaeo7yTbvEm7Vxqft3FhMLqyQmpQYu6mm5jDShJ
LajsSVJuwy4QReLgvm6wS/PWL/Q6N9ROGqtZlQzmJ4bowckIqShCIDOdXkpDrChowqOe13jCHVrH
VPFgeFBdV7gq3jv6o0RtdPyHgrWNxBZbvRFAOUu02hUfxbuKpI3QmoERJSuLhNTqYEpIx3qBM04i
aNRlStMnsHaIcsD1yX+GTuZ7U+lwJhl5DD1yY8Kckjr2F2J82c5vyxa1RXV58WwT/ehEo4QjggJ9
7WhyylvINas14wCZIsNE55LnWQuD/XTh9pZT1VWYp1GpP03SrxQPNQffPpX3EZm3nzxssZ0EONRz
l76XVdsOp0k/H3krcUNN6AvlU++0U7GOnAYgo4w9KPk2aXB9E0kFb2ZNv8JmRuAGiat09hjgGhCp
hJtCT+wIPEEB7YJmFMvmG+Wo0RZc2xMw9IxtgJvJD8ZIkJkzj1sNz9xVigaMbVQbLKYGRpHjicmk
BzqLYWf9UGOdw0/ay2DFWnWTtNpocbDoBvKUjgi9N1wz7fradxFaZ3mm8UWzvUB4e9RSe8umed+z
wG1f/W38h8Sux5OkHxGAmtM69IIis91H89iIhhWd9izSPlc7MfhDkRamj1iWlDgwRdMZeZRZ9t5F
WzYWbpGqTHzATjgdX1Q17JKVVM2hk9aUP/rT2mavVKqdSF60Q7Jy1BatmfVmcouETYEcXoWKCn/l
R+0xquFkI06W24EPKq35pf3vEK6ZK0fVRzZm9/fuCgaHK4jpDSNVqLRVsIpVn3cjR0GH6/XjQSkp
oQT4WG1EAhnbxnDXn+0rgZb5s2w9tlHoZrZwAMJudmrEWsDECtyXZoZR6n/HPvXV6O1GSkWvImMs
f2G0nnzsydjm/OeWY/AtmYkoH3hxcK/O96GM2ncTyVAtC5kPN1FvSpZCQDq9YnCdjDBT8NLdgZrC
ui1HThu/gnXAgSO9JQUEaHHIpBMCKJfJHLaLLw5Yen1YoXXkSauv9MzfHVXgYPr5nuR3QFAyJV/K
XKjmJbM3B5JJOm2WqyUUCzDhO8K8ZlMXpBT8msoXSIiceQpFHFGPHof1x0Lx9JDcb96EhDQAA+mW
cQYz/oNJsNAPbaunvQlIv0WH4LPUvSbj605bl/a9YoTvGpuZtylKJ4Oc4vhi0FeIxGMYE/tdTOiP
Z9rdbLDMBRLktDw7oCwMptE7TZ3FkC3daahjmVLiE/h7si6bs8weKHfh8QpODDB8eXXksrQX8cB2
nmmq9xffIlBUMTKHUa6mFJvIsjwU8KwfRkAzXaBCAW0bNkYa83Hlg0sfCSzI1p399ii+GebWaHFu
pLEmsn+PHoj0l+kdPRwuLecWrH26E7Dn5zNfrWpwxJisowxro7dro5V35+lzbUhY8L35zGzOvadl
RjfFwlxnKIed0OJYAYEv/hla0eEgd0Z0oC14Y7CDQrbvNIxkT5mchvgu+vBS1G8t05+9KjyOyCh0
5o8gOQ5Zb7Y3M7/XhODnWlZ9Uq/3IYpR99AuBmbhdCDDNZuhBIkew//IAPHM4sD4/JtJBJQeLOei
ir5UuowjT/RTlxc4Nx5lljmukqYZCMfsR2LiNsCf9zhCtdRAOzkA5mapmASLcVTmF0ag0j/He4U6
kf2RAeNiHV0RT33KEJmHHKQ8ncSKkw4LFRsYHB43R1qWJvNff+yYqqB/HIuPzg8aivo3RRrsVsM/
6L37zHBaKHhOANAfqj128/O/QVFLg8l0ixb71/fp0nsFLLD+hZtA8VE+7MkIbrbv0Fp9yobqBxsW
f43XiMh4Xv9WQjKocCsmQUBi0tYomumjpHJxk6LXnYZH0aQoQdhAggz2AmgDImlPMPLFyD3vwae1
ltVLsb1uA7PV21Wbkws/8bWzssUSTWkJCeXqLyXhSnon9fojAlJNWkF2nOp5cHxH7EetVSbymFjO
l0N59bk/MyUVWG0QMnBPK7J5oNuotnTkdRlyAXxbDRXDJwDXsNWTf1R0mWfSiIBgtIpch9a3tRzy
tYICmGHLutxmD4OM62J/P2fsYIKJIux4HhlWLkkHP3H74WFbvbef+qfqMfWQwsecQTt2N25djPDe
3pMF17z4t29c2Gan5/zQ76z11LAKThvEsgT2wdBU0tJSMSDOuQeBPIn91E440wGPo9MjxnF9ZJgV
Xpmrm1fDwxzkYa6l0VouzR+xcax/5YfZCTi2fllPoBAMHirX01rpq4sOSyd7skoV4vZHRg1mZ2DL
PVolzLBUr8jVr+oTNbEKMdJIavfqRrSDbYI9SUS0+9Gvt0MLziYbAGau6FzcNLQv4akJaFm0jLkB
mpda0OHNZGBKS4+N1vPJM98yoZsldnQstTQ08bfOBqL9+EVqN3S/b9yVQOY7ktRjPcIQChgLeWJa
lyAmvUPkD/iM9k8SrwI/SZmlkTxBeU1o7KVDvYFesdDAxWguveXW2onlu5jb6Bo7g+LVLSXKO7Lf
FQLGATf+/lJTdbIYPyOhGj/VRmploK+tXn5MYnid8ZqmL5jAdTQYwO6exr10WCmerZo2DRtpckkP
EJONReGRmuGOEG66gr1Uzrm/8Ulbofs9EluUuaDXmn1R3+rF7r1Vii5vC3cdbZVz+f3Qd+RsX4sH
bHzxEvLoHRtCn18e2R0ieSwqeMzkG8bPBMRwTeHy5eBrg3f/hytozDgZ9Ip0taC3rXuAfn/BNnZ0
9MlE1osiT2u/Dng2m2h/9EuACXQ7z7npkvIGsCoq9zRlmg3JZyhPdpsTCqPrPn/Y0rA0O8VMtQKn
/2qvs0IYQT75ltaXws9oBrK/5fBeGyaXCVrZrcCrqcrSRzqtMzsg1NKDqE2cDY43f+wSViAfQrTR
rFgnVNRzxFUH67WUrBfbkYyZ3OtZiWh6NaAmxkCkAjbNUqK66yaNBKDhtY5KE+suFJxb2hpcP/i4
vM3bQokuXyKhyfy8w04rq7xDET2I6lsYQokRbbGntBO1/FpDVBmwnLynxXkkNO8jKIpxP/MgySD9
QSB8d5oqYZ6Q3sT+3JZvAhtS262YiC72TR+wKvU7MfxYhYaTE6/IK/HZ2G9Jd/6oJsXo2GNSqFOA
PmesqrxF3ldoEyHxFjc8Q8uXM+c3HUPPKf7eqmT7wwVYUjyLrAumGGjVY9oufp8sLEjZFczNO5y8
FsHkD4kSOwp9DN64q3VpMOGyoag0lDKw9ovhfGyhkBd7hMGDoUd2hXrHooaXh+2HiQXo28Gke2rr
aG4WXvxptr3LwgNu9gczNThV7l7mw8ZsnCJXGUT6d5W35ADFNj8ezfY4zju4pqQ4ILnenCazHjM5
ZOZQJzfRjnoY8Cvs1hju10eP+GNvkWppuBBrW4IHZkG4ES/3UMDzs9KzzWGzk7Li8Agz0A8pVBsq
K1Nzr8TvDU0tqLcBn3wErlkPYDzDBR97P/FfHi82YWEHrZvkDDwlgCxG5q4p4hpFQyS4BQEU2SrM
zmgHAHSJ011K8rNL0U/QHf9R0OuPZaxNimQPEcQi/P1UoW/TGZosyJQT/OOpdHuL3TpfkjfxjA/h
q80NS4vrzweb+2H+E6Gq616IB3juo1uoV+Lb/Dqk0fC1zELC2Xg3EM6tQ67UjSCWZUfNNdXH5sVe
b5Fm7AeJSm9dKBdWijR49gOuXWcryP3DoBf2y7j9CPanySR5uubRLrkLD/BnmlsHeBdQZbhzC7kF
eUZi1ElY4Orysa981LyoB79afwoKAC9qsyOSb2MgtFapARW2pRga4/nClLYAqhb3QiqCxGIGlLmQ
Ew60wnQW4BLrUqwZhsZLzyujPHCVl3O3Zfi95/KUu5yJWwPBXY7tQFd0mzqnjDMzuU9fX+gBaCyP
P8WNmhPKJ3snfEv2ejZPES6PqS987IgdaciRcH7QC7PoWqHp/Wt9UScu3qL4FHL0YeDZsSSJ4fAL
3jrtHz9JV/9cIbW/XksU9+wmgYhPEOithU73cnzPXx12+rAe6FFj/5bSufDR60+bidohJy2W8tMx
wyeOMxWVRFl1+k8v3bsSMbUr5yMJ0val0OP4e7jdhiovF/+5eRQCj2hw7NAf9mVR6kTP88NajTRO
3MDpGrYUmkmdmcLUnXoZEJbRwJK5+V77dFVVI9LhkqKMal1U6EqH3TQTb/o74u6QnkLFBxs/Gm5r
QeokUkC7JSVIJ6QWsnSibu6XcRxby3VjaT4fkbDTv5OQ2VZ7IBoznyxnY+ojSKDBEam9HJ2uIxJM
/3hfEwLcaGwII7tqkCv1zlr9wWO+N9WFqOkS0JLubF932KuOmkhbcLwRZmiXr4chnpWQP8uVuJMn
6KSaNpU0Z88qb7DhbSSAcunZB8GVt6pfYS+ylWpr8ED+HclKy+FTTP76wcZeIiS4jMepoVTw8S9q
u+xeYjID50gxiETblizfqb9u9Vo5/J8Q2UaOXuX07n13jJk1/1utDg03ipZlb1mUQwzSqjO176do
jM5TIrbeJmMrKJaO2RbJrevel8HyVy3baYWodfpoESUMenXfBs+thhZpmeFIFzdqw7a2U4LjTyx4
UXH7asCOltLXl/k3QoQNKt8tSjn3tGFqRNJsg2a1HGz9Lbz9r/8OvdjT1WqYzk2xpNklrLnlFEN7
ZgTxy7p91Mgv+xTVF2NowVw55leXFxT7Iv3YZdK19pgdNGm7UFGomLl7ZK7qig/kl8+ELNrHiiqZ
grgOk6n9MpW8DsumkSyA5gBCByBxUAsLU1jsze7FQO/xSSEj8FQPnBAoQseFwRs4JO0vUjbl8YrK
IpMzCOWJHBYkVElZirIIqoy0igZxQH1m9gQKqryahISBOSekEDVGgiEmwTbMAzkXFCVrAk+rC+nk
gTsnVpe/S2InDzdxKj/VF0pcTFJ07pH8caYFktsp+nShnkx6O6mqsolQrvhkNAZl8cFXvbYGpHyA
NLza1nEPZPczw6TfNiSmrq/U8ci3gBTDFa36Dr7yo3e0RWuzsVJ9ISO78izV0BvNv1dzU4Jb7j/K
NGdvPoD/CQbFiN+4ngz29pjbFqzQ/8RYCSIjesgdVFdb7OlRfsd1ECfcBLrI/sQJMsX8wtIEa6/e
7PvBeGOtNzwd29Q6E0Jgu66k5oNnYdwc62ZVIhmSaZJg/yz8x3FB+fZwqTeOJmDErz9VT8/yih8Q
CpahTIY1XsBXut2VCvYh445E1x3+xcYoqS5VT/EYPBOdRvk9MuURMaXFgvWp6qyYeNrWvLIY5Rdd
etdOCtxEyJsThgx35Qe4hGX7cypCbjBWbEOVr/xXrOAOqZXz7cfFwxVQgWSvaKfHVcGoVerOh+YY
+kFCcSM0qFwehkZ4xF1UfbV24vC5VV7oLQzlGxTUSqNUKV3XeEwDAYhjsmJVg07xJcvWR4gr8cvv
ady9MiHaO3Ye1gHjApIKAvB233NNtYVUx5F1MC/3nihgs7M1aAVOd7JwVhDu3M3EupAVZ6RNDbhm
GwRNcvSfNx2xTSFd4jRQlLVh/OdqoHlkO/wmdGrcERmzmI4aUmLugdjbGxJezbFc/IlDaY3lVmOe
3TcR2JI4sbGB1gjushAfXVWz8duxMURfs0PrRYHGJX221NotEGl3PD/FbOppFaQjI3gTeZvVUzIi
PaYVDNYP6fG8F7pUp3ps3cqOfIihq4nRPwLkhKsCz9LEbbxKQLrdvi+S81R3SsytzC5jWQ39/pV1
rraglBaFSpTQkeb1hH9HuqDHJ5hYUy8Vm2JXAEQ8Rli1yp00qgbiWvy4bSvzXWuN3FOM3LThha47
QaTLk6E4VRFfgRooFb+KfXEWi9f9/2gzJ6w5yWT5IvERJZvDt5liNnoxYsYNRHfstLj5PVkzgh3D
pu40hJRUksGVlRgPsApsQ23odoIjLH66xpdoan94v8xYByxXtPlUmbq1e+bgd/gOPOHHX6m4vEp0
PJFdWVudC4IhDb6P6g7JUeucI2UhMxIi/9ubp3M5TLl0LYKeGZcQ9lZxbZaddqc2M83kopUZViOr
1rsM5JLvHCyRU3AnwQ6DiU4RMvo0knPHgmDdp4pKhi0/2o7VhUydAuUSRFnNQqeZ8UhcAyR8BlLA
94Rg8bdEg6a0XSGNUIpdSTE5WBMgCa+d537UhnqQBX+fQrnHkkxbz3UVjSZu1fX/OiOwHdhZuIUl
SmvXC/H6KzeNixYLZef4T3BqVqi1ShIfniLeuhW1sK1R4wSY2kPEWf8AqrY9m8Q0UPU1+wDkcC1A
bGYFN/hF7akj4kMMf98xyDbr2uIQ5S+pv7Z6EceXU0HszWNN/7IesJ67KD72FCRABQUUYRNeWaXv
odX/BiQZV5rbHYhluoedsh2bhxDRd3EbYG9sVyNmysdr3Hfsys/ge/CcQNf5tmtAZxEsF1lQYGlR
/bTSIvjmCuXbYvn33RnAToP9j63SKC3/UOVuw5eVkHhjqTSpr+t2aEIkAsW+txIBUFnAC46DcCMP
v0hweeqfUzQ46YyedwI/9XKVzU9iKDkPDeTmTV8i+fOjXYFKgIAyN0myKYUbE6eKzHxwGc3iC9Mt
zADN0l4nbshldUr2s6i9YCwYM5WEKrsKkBA0+isct4REqQr0kRAHP+MTtFCAZfbzM/cU6eTNV+gE
qPdi/pO1NE/BZNb7tdbT9hl8E2SVQpxXCRD+gdNX66cUPu5OlxGqDwOu+UNddiwBKwX/2VscDxIP
R4ly2aa7FzOHL+xAoIcF8kek8UWhbBqvXvxxJILhvD5gZMtX4pP7TXeBlNAr9wMkuQBs6yO7Ew9b
FnyO6a2zFMEhWzMfsh1L30F5lxAqrzSk+bokUDky5jyWfz9fCSSkWbyEZz1rL2RHM1ViNdry06Za
KFV4uLVKwnnnzwXCUqekWcBVwv9/H/cOGm33wOkOvMA01zSus69N+DUBTGbhJFNk3UtXbzIwbdEZ
paLizm7yQ0WYwbzKYlJxd0sIL1DpVo2Zs8s3FyOSX9yyF1fvYpVG6cxJsnnK2T5So06Z/Fi/OQWJ
ojgTL3TTXzgXLPPHixwJCtHi2EIokvsCNTJHFxSqhZYlVOCn6SNzbLc8FMsDUr52wIpHiARmgepd
7svo34HQvxE9Cc65umebB3lWyK9VSvgJfp+Lv/Y0CTPIN6JTkt9DmvQp6rOz5Lq0HfrMbbL5b8Ub
8mM4QCj0CpciYcnmuyOY1jKu1uYrE/4LuLzsK9xFLCAATgEs1J4r/9kVAM3UbHpyYJeFR4Ik38Sv
Z2qjMDiR7m/yU4SY30vynO9GKwyz2eJr5vwNN68JI9f+XLHmLVFYxoJp2GmjB8wwDVd7sS4rXury
BXjSq2G/DXaSMA0/pt8VlWj3vGwYKOAC1mJzLYgvzKu9E6DkP/O8TxOtIcN443O4rSHcoYon6l0G
IZUmx/aQso1XJBqPDf1NAlUg1g6FLkyhFgmQ1uhIpuy75GxGHzyDfwbZmux4jOyB5b0JydT9sgKt
YjkJXY3mUN+EW/FXA5/85ot7oDG69io0DODhqKyn4le4ZBnZXXFsvj95wXc9FP/x4w9SxGHHBJge
Yj6T9zaAZF7+L5+kv5eq5dSS33xZWO8WjHG0dunhIdUt78/cHiASSxe4pm6y70Xtl54sO4+0TNXL
OmDROdg3dQDWGbjU9WteXJUiUHZyRoiqEOR9Pg47RlDOsg/65ptF70lsVrQNnc5BBFDuhCwCs75o
jlv7XvIO3Y51etzwUfahp2Hv3uuFukDMtbUt4ofktxPo7yLX/u6Ykx1tsXrwr/YiOitiABDTEC5H
e4S62PhrptYSqdz3sjI0AsvQUJAvK9HXq2M+2tyRelHjcMNa6EBporjBmbaz5KhG2lKgUFogQeYu
K3Wu0OzaRM4KBUK5IHoLqs+Y5ebVYKEFeM48iaPWVzr8dHY+kNFGpMtRC67E/hFcfuwdLdx92bWY
x+G7S1cui7FXiABeRrXavDecjtcZ/tKV3Y5ZKEc+cp+veJuQ0De3iTovKA4R7+hu912mNXdjAB7S
rGhkR7sfLIipuS5DSZc1NzAy2e+dAlLNMW19tJc8OW0YtgIxw0PKlZHjxXjtoHDg0kbP6AbYRRsx
ax9grb8vuBSslDsmIM9I5+heDKOheeTgruAUyZCpXOAT/0IqAU1m/tNcHdekhRDIIpAQsQee6UJ3
Ra2vw5uBWTwg3c8IKRcxbTSUo6MXgN7w2d0Ibh4/YJs8YbHjwsKO+T+LY1tiW9ja5wvVtVV2mvb/
U7w68sOVek9m29omAoNDFDwkD7BWwV72rwGdHGs/ROvN179IEasnRfj6vF68KRm91+XJEGixASI+
leFQfyiUB08SKj07eHkR2pLH3BqzeaDrjuIHOkj1B/9oAA1xE0jgJ4+iRuA6WK3rognE/xhU9ZPr
izRSnR6A4PGPSJ1rRNL/G51jVA0UXv25eh1DxWQl2GTGR8ZJrv3HWfGk0f5MxxANTegra2P8g2uC
qrWcmL+Qz6CrWcVEtSIr6d/39XrzZofJ2oDEFkCmeOw3J83Nyy+oXn5k70jJJM58oD97j9Xt+V7F
1E8Xm0CH8JVpk7gckZVcZGA+CcCmwSO5wQEHehuRPPv0nFYBMwSaRT/9Au2uG6zpnFIPNHFFMcL6
9lyM54ITuQjgNLKKKVhakuJat/iDkuv5k1STbEooy3R/Gxw+OMzDRHkiC6vD7r6bgCRQOY8TLX4d
0BxEPMiZdhRcaBWCzCN4/63yCdZW4RlheMqSKc92vEODmcAxn3r7y5scMzVQ75YTG7j2oZzKEJxg
LOTm8g/eNnl3tBVk+BzUZSQUQgHGFxstcckgzEt6I0U1nR4uLVZPzbNefcztlUbcfKDkwsjeCQva
5HazpHXAcx6r3nuqjx3/UyDi5xZZSvedvoIMqytuBcq3a2CS4mmasTgzjc33ph8Ala80hiuzdTKu
oEnNkSt2yTr8hbYVUemsbDez6jrf3aXQZs28OByWm4Dmpbcd5DvRrubLdczRrl/IzRX8jUOw8Uw2
ps1mZO2cX2l4X2lxnF+ZqJvBny2nbpLxoXAD1VIli+QTQetp7teGcBIihRJRdUDbPlOeN1xCxlL/
EGmQv5gmFqAwR7V4jkbiuQvrKPConR6Gk/wIm8dreNj6uCBrPXc/fESoa529OSd8RiQenrklmy5k
cWTCZmHo8koOIEE4XKKxLEldzEfiYDhP3CggmJqPmSQ9MBrPpkcwBFcvhaOSrn53UkgZqIe/wRbh
3mSsuqLNQf5vMh/tE6oPzzPn6RkZfqkt8YLz/B1bZf5gcv9cgbBTwnuRpOoVkEVXv2j4AdLjsMDg
mo4YuaJUgksiZn/dXrt99ukA06mmK8KQqfWxfEm8nEuArTaHZgR1t2sf4ZV87stU8M7EqkKx595f
zfUsfORn3CRkI72mTXt6cX3JazdEHBAdtsYZaVpNpR4AGvdGla7F7WkiIUTVockNVh99xtFJbVdA
6noayGS/Ma5qaHCBvUeT3WbOWaKjiEqGgveT+kZGSQKw4iO8HYxQqvhrOG1nFo/24/Gj6CLn90Ii
iJwAoRWqA5FwEoEDsVDMVeetjzPwHA4u7Ea2YtghdV4bjn1NRe1KSoBKZ7ZMFaT0wmcHzAwkhFqY
022Io6b/FImdjKbLevVNj9PMDMyn70gi8hyuEJrYBBV9h+ru8m2NBAhBl4XO1H0GfCVVbOY5GH1z
poKQ0JyzhTptYqZuzZdiTtl5C2EN8BYDjWdPICXYslb5FiTD0OnnmwO8xlij2/K6TN4kTFNj0iVR
o/0atT/oxEaKK7Uqa/nqdAWaVzFeKo3Mo36cZdC+ka1GYuj4jcJtYmmPzYFcgboOQGPsL8jVbmwY
NLrRDUUDV5ekEtYHOk7R413wa7G8/pZWJFaFRpCSJ3Rrv5g+QsSZxrzMjbuvsPTBCCrplsyaJ6IH
KtJ1cnjU0rT2IcAJcZzcmAOzK7vvFCdc6VKPMIAJiSkeW2m82Y36G6er3evn0M0ElQ3zr/tG3xDC
uIsVHPX9GyARpbOES1MMnQKLhEr3horhwzJLR+Sd42DPmKHXsTDbMLCv6P0qXqvaRv9UFni6pFpH
RJ6Jhpp3MKfYVLL7Lsa57IRcvqKvsmbfuD+Sfv+b+nhP1TuRFczjnmmzgI/n4+4tohWIxPc3dTCW
jZwFw0zq44T/Do6vTotJGGaqOyXyvAES1c+OP/BCrqcglH5TRLYi+ytLo9vTxH8S9TME56u59WF0
nqatGyqEm+W0oO+hJQTbdbJdaKLt1o1zxIewgzbPaOdSBR+4y5hKQZizgs1hC9jMjDMopV2I7i5I
mGTnKjllOuUCrPtAoIRTVLpWBaPvfOSk+nUv0IL+8wmYo30bYsJv/nSG2weUt58k6x/ErF9t5z1X
kYq9866HYe+1qpzJYxC9EUw82yUW8Dm5rFKhLVZpI0MBjIT1d2bp2ox3EESi7pEgrCL7wijoDA+7
rblwJ+gwqtCdTsqR9cp5WzzEgKpNKPNe++CcOEyy6d6Vs/M5atRlvkfZdiDpKD6ADfXP9C5KpWRP
2VzA1NtmUb5w7euAU3EHJD/367aKuLZKZ2cKZZpsDZh0ncFw8y3JHlDzQLCQG60T9tnwsXllDrJX
LonxjhYX62tsrQvQZbL7LzWFXUElhUt9Zd6xl+OYTgAoh9/lR6fCBAYfECm6YaNbL7eS9+txeXg2
kbhDeiqA39MPledr7y3lvBc5z8rUoXEdC+I08ez33EC9jOi1XodATLrqiQTBogetiayQ32zLr9/L
w9Ki6pkVbCuvhrK0nhpJIZ57KBY8qsppdRQrPCcRLRL5wN41i9Eauz0oCGB4jAO0tqjk+TU5IJM6
6LfShAfzvyLCOWQPKplIiVfvCCNipmSVjcRiF5Uoph/1dH5DVZIdtXNcr4bcAw7T2HyG66wsR3Oy
mHUhsyfEPaDOrGTaIMnITEkQ81IW7AnXH3rZ98Huraj8CbH1U0EZOTSR35zCQgv19NpVcw/gcxdY
1eDOdXAj26tMxIwQj9LXE6NiI7wAsryM5JPkJvsrPnQCaIhiprirkRvcEJPrQSnDJyKqzGiXUocu
DSVaGATTQcsd49Tfeu1CBSuue8IQbju9atIXwGHeUivensAsEwQYCT85FOuJq8EZWbePtnz0TOu1
Vez1GLOXFmWDTeZtpAM5GoRVuxu71+FKnFhgX1zva2RC9XkuAcQgl8AoPbh47EK3DMwNXL/Aspt7
kHZ8B25dks8Rqwt3ejy9ELo6Wc5plST7D5i8th0ft4BTTd6YGUtkpHMf+PRGo+/lT43Q2MZnknbD
r3zWgYZmXYFvnPPojmDMj31BA7hSE1jy+UbV1TlwGFGC9tC+E1NqtfN2dPb0RSXayzHs3Mfoc3/J
82ePZkZNO0xP/5vAdP4DeauDvEqogtCadtFqG1xBjBERzSKjTk5V77LJhLoUJIGFN2+mAbayYrA5
QA6ZvxVjCLT5gSY53zeRyko0larE6bdnw/U+lTNj80zhWOaCgVcYLFN+aS5PFEEBDKYZyKapEXeS
Z9aPQwylorvU8KYPsgTWr0eyNnMBSptT8e0CsLpgc4jAua1JIS93OZ4l+rMEznnQzh8vfXXo40Dv
cbmYVLL5IB8kBp+HJ5/fp2wMx8Ig59xhhPD/jjHLrPe5VSCtlnhBmS3bPXbFLeQ+ftv3YpfYtaLe
OvXp6bfSHwrT4wOr6/67JmKLZXOvmN7Wq6RDXFSf56WnpcXv3MuKFA3oSmilxmvulSUBjsWvy2mp
IBVbLOK/tUmJNvBo7dJ3gexmXjFg2ccpZOJ7MsZd5f1czM7Fo27+2Pdp5PuUsK4nQoGmvvj6JiIL
Iin3b9CUw2A1gA017TwfMqMOkNPhlu4rAqE8xfcF7R1IEgWQYldifD1qiXUQ87F02VKEI3zR7lFX
PaCQ0CykP2HaJm9EiMk+rzbIzrrQkaIwQLuZGXbrdXIjTdrIxXkLHp6DZ98W5tN9oZfoJXfLbx06
1FVUI/p0Yx5B5fXJgNVwSXcF+6YM6tgVtQKM6AyqFPFMYN67pWCuRBKuwzkqOAK9xZWJEUBNqH64
Ndki5zFuf8fssMcWP5Z+Cig31R8u/nUDQ1xpLzeb5Zc3xDVudvFFftA2Poi9UsiuYgfmaHQ9Nb5z
NYhMQ66fNov7b//oglG0A5LZJNdDTxfGnge8T6GpSGEz/ecmjcosWPogGfPGjsMcVHAMaSSSt6GR
Od3uBbv8ubh87JBCpv3PfignLYDzsEeVZL3EaSN6pxMtBe4S8QT16g6Z5Hep7PjWsKT8bAyyir/t
kBsPrBNphyQoNwATTOy7colB434DpLjLVP9enB3KqKbuRDccZEsJ+nNeUwl9866kZl0IYIDG53Ju
eN8pWpPJjejhXCd+WN1lOJ6Rct7uErUhlGq1Xo7/mYFtTXvK8ULpZU1GVWAXn9Sc3f1skJ0gZdlE
0j76yy+HwG4UyJ2+9dTd4vEGqDYhj35hz2HNzNX96rdtUCz+kJLJLC6/qo9elt1GsbMFZ3s/ZmtJ
6StBNP4Dst9eGxTuzTpCEH73BfZ8LZgP/MUmNHmP25XbIh9h2JJaOAjxvPVfZ8+lcVjGfUqgLs2i
plFYiDGIEtGjfHiVTyEnXAFgEi6a1gIqV0qDjOHI+OJmuB8SRigbt5XLcLotvmBjcqd3YCpnb14L
CEC5fHozl4TeKL4qD3EylPVhXhV6K6NIyJh0G08DkDl0TJs7Zi5knX7xDUj5BOoSmWW+ieixBXtI
Pke+6+G1nAfJw9CHT5LrlBZxtPFlvUT4rIXkz2MdRz6I7pqZT7m0rW0UWMuemxcWEJUoZQpb+ug2
rNez8Ah5Zd/FOf8To+D9F+EkS+hpFaFuHPH5gjAndG2HMZ+TiA9Rl9sVRN8zOTN5ufUCYcDqNvWY
gLI7z1SUzT7XUa1fulV56tGDUXJnvY1q0rBlYfxjBCQGV768cwRgq5gdV3BuIDaal6Dqwk093+hY
sA4tWm2b6hhcRmEjHKFwwwo2z/tg4t2guYEGdyXay6OkdBbodSzDVp+FPUzyYLOQOcobzb91D5XH
/mqfESOkcxHb6Q59FjE08HEETEVVdQ1mi6B3Epg5xEuFmhFv06nVSJ5JAueX1vagn0A/9kSB5YkT
UnhNMLIorcyliaaVGrUIK1o58nYllYjL7z+rHij1bONL5dz8pR3iKcLpOGpV5ZUbEOFKmFVg6yeJ
KgNmC05gxkxBMPZjbwcBtesK00iqgmxMLwghKDNijvfteZOKnx3y0NnA5Ygqnn0IMXpgl2G1gjaG
mQHllbr2x185t9PS4PjbIUkYiPiwOK1GEzSFv2m27+8QIRW7/Kd77E5LN4XAc0jqPeFeLYGye4L0
hNFQQvtGn6yuUwfePX1ipODH1q+qVsmwWHCpAlJ2SviX+LgxHo/FWh8x2A9pjpblZvENuX29O7M9
2UvkhInmYm7cB7b9xTf6kC0wIf3qzIeOdNXQHJDi9JveSJcWjDw1ILV4D4tB7Ul6CFyKa6CdbDoL
JsI4wkXXlEsl17Osyx9mYh3rCpz02EwCUJ6G8axcLGk++lepG54+sHLZSvboLLzlyEJ0gkN2ADKj
EY5QP3WPyZPcP4i2vglve2IIiMhnlRVFKNMXDPVDdR8J3rtMQQIn+e0EDnPwOUoY8c2BNtRn5ciV
Ix7aveIbhhTVQbWzZ5DGW5UzgLNkC807gs9SPg96tpaSYjJSy075u5nw3eHHt0QuPQ1u1yg0SmDi
9rgJHhNdwFAP47z/dWH6rLCWkTMpJ/UYPt35g0odnVaaT2p3Id5bLPHQ1yYZHYgNSei/M56ex2VL
oLtAFvLp8DBsX+e3wkDTE0Vg64GKuk08XzmbuMAzm8CZV8xoZlXCxT079+iFaIOrg5f1bto916S4
MpGFvC1pofQgx6pR+OhNAzIeWJh0V8tiriP+fI6dXU2wdXRngQS3Iqb8AHBRpznFKMC1zOg01LZ9
E4yeJCaQK8EtKTpUKEYKjGeI0QjOoGvs4DjY5yOSK1Mb54hkbv7zowUATqgMi9nRR/vmyUU8x//O
tEivorX+i9hIVsgKffl4c4bI2AKmLYmG4LApxZPya6tC0sSyxn3lGUkLuMETboXLTU/j4oVl57hR
JS14e08rKRJhsr9lpZ7ljuCHv/qfF/hau+33WhwfV/QbOntNjWz34Gjp9Ili2h2HTyb1ct8q+Zkp
LB4ro5eVe8XCn1QDgcjw9ew5A1oFjF5KuQDD24G7zaHkg5G6fGHwjtPvq8o+z5vAQrdsKfZP0D0O
OQyVXbkUHk1TyHemRRoJ96fT65rCLSzYhdiEHSb4ae2L9tn+nX+bPrPyyrCnV5vmuEM62d+HdHUH
jfj+8QiUDGMabFwWKT9Ov5UNparIt76PAK9ZE7WxuBoU1Wiqbzs8j8cvY9Rn7JAOQP6UU75dU4jI
0C5Qhr5nu7bIqsTjYoXziTrQgQgLZMarGD7hbkEMD7eFO5z59uW2/4+UYmstvDKA+r65aULM3Dr6
/MhztlMdvmR9cxd4dtLDbo/TjZFZtDRpEoJ2FoZxXYNiio1pJgQD1Q3D/5ENTfGtn7OpsIjuriHv
EimqptHJ+IhleUaQ76AnTAiYza3zKhlqXtfeKUZRtBGgQ8kAI/DU+SAcq6VPFm34CUVTiQJTHc62
Y1p20jJpNzjksq26RT8SzpbGK17yXv5zYvGmXW/4/VHbrn7of9sOuQfPpwJqpAValSPAfBgVDvIc
Te8dOPGmfBAQ/cxRSofQfMISbVjgpTy5u8iicQvJ3mxPRfSXmMjKWPkxxg/1NwXZPJ4TARFBEDka
mFxeHddOTCcvBYr5/MBmUKrD9uovqInRX7bHM2Ktqy/tjHgVMjczE0KWElc85dsZOYOLtqnY+u+R
E8sIrEKN2Gr60BCmFYFPP4rid4HaxVyWI6CjtKOTypkRnIcpUpHHlb9PXOlpbUcP42HOlq7asbz4
qwsYzhTxjg64EJ6LELLBPJHbMSPaaqINXR/vLMOUU3pYRRWAGtrikfL339LdLmy1o6edXviyi1wi
C8CCOU6t7mA5ZVFtgJL7Yjmemw705hzztJ/OmZ02+fBu8Lbn/OldEuc8nCX6qxdspKbYusk7u6FU
vfJTTF7U6L0XZsdCx+CKqjnYYSDHFkR6JkqsqVUcVGXWk40q52jrshlx6FOO4/8GVqVtLYNUXTph
gnM4cr/KHL0EZ3V6M80lpe1BTGwTxjlAxQ+Oqr4SXvAZcbPdc4JqNqwxn05horNeVRc2ojbh/9kE
Kz1PddGTirToBZR8wMdc7TX/sXuUt3hZZDM6DZgnnPzu9J2ntBgYf9jDTi8eyWPxhsKvAGbODgev
Fv2QrxlUXgkegJNmRup1T3ffLYpy9EuzQde97qknDIfnHUytgiGcd6W8/rSl4ccIVNKekLl+ejmA
l9p9cx0efbfwRvoAFYg4MpJGZxtDwUzUbhV70nTUrwmKoTjbldRGPowhHC5KnhoOqaoaf/I9FpX/
PjtGT/tRTyOviKadl7bOXBTxFO4FqQkirMxCznUaGapHPX6232jFP9AtCLX9tnmlB7ozl9qEwp9U
+DtBzvwYvss9BWNBCqpcXsy7OK6PrMUdfTJ4kqjUtZ+HBQG2XL19JcPqw4NClZyfNZEqthcfBwik
ycrU842NCEYanHOUp1kxZ/o0wkeRiHhNSYeAQRsHihtm8Y8C3wmOCuZZx7FGL6JrjizZC0OP5ZjD
fwQGB68jfADIE6TwuQsQm4XdcjrOH845YFk8n1wCZZMbwErD5h9J02ETpp/Hqw9ottkzhU/QN3W3
cbbkxy0gTDMuq42j9BEB+ibQZSIpUQ4KJ4KL286CH1mVM2VDd98+bnCkhi9vAuAbUGBCuTdYl0jp
HjnXZERg0wuDQEtcre13P4+WDMbFHrLyNlyTjet3fVwxjVr1SJrKEnBWBQlwPFjpjmMhsUsE0UtL
oIHohTd72fjvoKRFAnVSYgeZ6k6lKeIl6UUD4bZlaQLYrOAqM1Q9MmP2/Cmf6/Z/JU4ONuai7d59
uAHIqkZ0i7gd42ce9eStpYXZM1i9f/l0BhXxKt1v+amQvQDyHTC2cWdEZbpiIFT6McDCvqUCWHpl
zjX9q2+gpG5gjoqfAEI6HRM0ZxU1revEKjA1V6s8lyV+evwOdJuHEczE7b8FFm4E4ztDaKrB7xco
wnBKY/Rzn3et1ArhRh40wpw/FcZWcNRnnpzfSb/NaobCOinJxMrqJPmdnpIqXSQ8bToTBbBtYuDu
tY1GyEzDHEKFj8pWhcTunHq5eI8d89+f9o1yDXdM3n7SIQujUi4RIWh/87FT2MDnwrpTrjqu7KHg
r58ZdLNTkZBXVNjD9Jy3+3DoYxNyTTP4IqMfrhYIF11GnBcmsaOLjRkoBxxnzViTbyDO0d+xyVcm
TiVq7uwQ5pppMS4V79b8q0b8jeoOzyI/2LF+m67QqTYUFEXcu2ZjZNX8OBzIQtGzYQMk9E2ZbbHB
uR/Xc36zXJOkUkrpXqSFNlhcB+YYkuEV+0tdRp9zmYTfZ+6Eb0qIKH7bjOKvSDvwRlkxoLZsB8dj
KiXUPMF6QB9e6i0MyxIvX5hv1/Gthu0Ec9hn2I3xaDEXSMGwpalBHAdMXuUHeYQkbrxYSnLsZSJC
cTX0FYQ3Y+cHJ+fm3zVQepz6Y47VGtJUduBir8OmG9ohIyEBJxgmpT8tw7B2TufRsJTHW7Z8E4Za
1YeM8wMZZhGDCP5wvHVo7supdnfWUAqRR4gRENIJmVWIn/so7I/9LOdwskmiS5iq8tITCuC3GsHS
lgtcGkOYNl6K53P2xbyigy27KtnMCgGcFUTj/GFKpsgridKvP2J4phUfhroQoOc7mgdPaWW4gL6C
NTh/3H4WwXF1Xq0HQP294MeaaFp19AV5Xs3HzGvB6RgFbLUj0niVdxXNKj6tRK7KYqio3LaeFSwW
zD7PhRUanOX/EbbHJ62uz2EZW/pLv1VQsBy8fcugAMnUjJOfHCp4imV3KeC9/9fCrXh/2DMl7KcK
6H+PMRdgL+qf02EUpCOXActyIih0Cj2iBIcjeMfVG5eukfzMpPinhNdpSKYSUG9cNwV/iQUU2AsX
bklz2rFfwRyS6JKwPfBieXNcrcg7GUottt+m98zgNC0NepTeKPZ6g2YdNKKPkT4aTtUbrNJGwkJe
rOKR/nJXPsYkUlhXBkpSSB7tcUZOmRfYGDOhm/xaE898Nd8B76m/6XHlhuLtSG5kjo8mUtXcGMC8
Uz+/6jr263WUtUpS2yhGAeeUjdmm7TlrsKqZDhXzpGdt/5zrNWLMPGpNlr57dWgeb8yuRtghq7H3
N2ozLXMh6AWL041fYmPA5bx8t3OhEgKpJZ2c9qMnMSjzBuy0GnPHe2NPJE8AfVE3DtwJqJuI05oR
vZ91LWSF6CwjyKSaI1EzODLAqmXy/XhC/qYv4cs7mwnViuPBnuJ2JzVG5kx2UvXNON0JK2E8V7el
a49H14N01sfOj9vMfEq9/RfbP51tW26drsyRPGf2aIDh8H9moeo7GVVMNsANjlnW2Juj1YwkEwH8
2Rule3jTa/LsoOHuNhaGzQe+5unzlBuLiBiiPbOYDboz01C+35WkwRz/2emXy8GVWCEW5PjJtVH7
+1Y4nda8n8QpzdYSn831R4hIiwoOrU+VVAiow5/aC4oGw+Y2fInF/8L+IeHvLFhZ8ZiAsruhD9G9
UQLdty6xjWDqYoJUBdHT+ze7Q2nBeQ/Ck/mZukFjTOHZlx5Nz1GosZRPuQhwGi1UK7woWlyTp01j
sW8K+pKSOUK3xKtvkIKGSeI0GXONqUHmn6mXS8+fNCcdKSdNaA09T143jV0Aza7S93HGYWV430ot
s73alZ2dpk6gc2BhVPoFXLee6wHKXglhKx9FoUie/QWLamf3u+vB+RIJaIwAWsr2pVglTpmTrLAX
QrO5LSbm2EYyg2RjEu5Vs7/dfOMpf2xKlXnITiyTB5jkAvkeZGHfzgS7XSIbXXw9x2qzJHVqQibS
D2DeojlOc5mkbNQNB5+v+xN8yv3guX96fgL/JxQ1oRnat3avyqhiSXzpg1jr1uswV8YZsmMyOXR8
DQO3TQM/BvMDoevsOwNCNWpTEQ7qqW9cfNbjnXAXQgIg7bgimnNUX4tv0AT8IHOwx+rrR+CpXgsb
LLnF7q6RNCIUiZmoFCaTUQIL9UcbFMIAMsv2cDsBY54bkqT2c/4CtNVto4hNjERs1fTsX0030zPk
UFRE2Y9L8dGJecEus0GIDyj0HIZG/dQElDtzilo49SQMUAkzBwLdxnbQDkYzlMvt9HdS+vsd8BNW
GpMcYogdAuXPnQshKapX5fNYRQ5Aqvezixcd9ROl0rJwifeDUorn60AF7golNKt2hnG1QNhX/1MF
jSdBkrnMlFFC5KP8/sMRW8FolJmIVsLulYIZRxQNQofFS0eWo2qTr5qhj47Yz6rZJDSy1T0FVSnQ
byyX+atutFtgiXMbum8fQ41HpcF1lq9oabLf9+szAlbeuLYubu2Tzq0Vh/B/+PCozBGQVXhh2p5A
soO9U+58CCdPXQhHhIShCG85dOGTE6OykoUiTltU32uz0JRxxEYyInJr0twZodgl+bC9AWE7I5w7
KGQmTWS8aakAbktzcCqXXLpRgwFplyqhFfGKeQYRZLi568NwjRNW9dyd565DB8SU/C88o9oF5SYB
63G6hwCGSy0XGFQc3EjbnjMatB8e8KE6cyHn45oCgDq9PDPUnfFOMq9UeUaTDIfbbLxIW3keZzoL
MBoGtO/4xQ3rKw68dDrjDzVRBOjnj6RkWTwlpEqhLmbYMQSfh5dafCGPyxe84SIyFwH53SAYsq/B
Q95EpxCFtoSDmYNeygqw9Dia2fCOmQe9hpQEPanSj1bItqdkG4AgBBXl2tSKuKPYVUYj1zcyDzoc
wRvLA5gdHerFXDNzzXIGsjVRWD+NfEADV9n+iKzHvZZsW9RdNk1w0cmwGYHjM2TwQHh1NMUuM4QN
EEf7D54x4GOecVeI6fh0vIhtCMOX5OCi5g5FFYFBvAPfRePi86enjqu3sWufsJdl41Lo3IFDUd+b
R3kLpmiguoQdkvlagqGyJRsse4ZHHsfLjzTnlG6TGUh5SShPm0OMIzuANHG5BCg+Fs/Q/lSUiWpd
za/DQj4fytFYOtxTCAB8PNizqXEX8B0FkeW3Uwrbt6aaduDdEVfOrzP75N7/fAupiIUynMKk1nzB
O57R0Gb326HiJs5PzdpC6g30g+24FtgqXfWJBAmbZK9oeSoS7GGmm3Yfseo2sx84vkTDiIzXG3w1
g0X49cf6ftv9gL+4RCmK7b2X5nBYXWsSZ68KDTpg+7McNv8rAoJiSGmyY2NzKNxOsWts777vHytY
mxXLfXnhcy8hrGEv9xxkCTxD92R0ftVkYeRu30ZnWdYsg8bdvkvL4tkka2u8HgIUO9VxOl7V9ikS
KNTASZnjKEjPSUjPo2v94bCJWcgAcT2TaKaCl1D0jW2PtBPzIlrFPTfB86GqUuNiN56LEOgX/35I
2djC3oBuqe4xBhad3yO4XO83S78Y9HVwKsFu2+sVmUsUtBoAkjA7VznWbttayVIhsjGWcuB7krO7
dDUgcSkfJcawU5LbaGb4qZNsx7OeZ2eJDsp1xYwcjdN7eu0dIX3aU+qvxl/6p7+1Iwz20/bj7vZF
Hqo1cTOthb48FgqmwdOqxUKdiPKBjQGLH88p9Hg3wwUCq1K62f8CG/3wjsUsJfLpj1HB653dJrFJ
prWzgCU7BVrFQ/NObu3C/QcRNauM3Kd+AlFHZbrb6/f1QvjmdVpb8fvE51gVqK8WMIXiSjpQdq6W
2EGIqljPa2qREkYWsfKqTJITtJ3osa52NQ8vewQ1gGqXpR/V1WOqk+ieZw4Qsp1gP0c07pdbfPQe
6wzkoMZNCPuapHXfSkvY2NnHQ4Js20OwzJCQw5vj525acFRRuOWA+a5+jNxWk6QrQMkwZV+mOPIN
Fv3QqTNAylOdeb+/7wYWwcIRUKHbUsYdg2Mjx49qkV6XBtKlVAtlm8O6sTn5FREbMPPkW3wYagWQ
8soXoiltRWguejpexbihQDs0JZIQOTa8/0dx4O+ZRngrygQdzuiWObp+cIJTgx05irQKMV4JJoYU
DhwOg/qUq317XCiziAPdRFzlR/7D1tqi0FtT2pJQ77qsEY6EPtNJ44TlpSo1f7+KpVyIbftbBSzu
RDgufJaEZaOtshBpZ6wsiySUM60DfprOnB/glW7is1zSwQngGlUzR19I0dAT4QmcNZjbt/Xjyp8m
nblo2EIOoZnatbgddd4q6ACxPKlO/TzkRQqqCVVLGhC9aZ6w4Ggf6Z7sbW/b/OxzWAl0UzTmWT/G
XgY/1sevr1peXXJnA+qxE4dkB4GXmCj1jipdu7rfOG58g+asHg+YD45QUF3SgIcm4TE4WqqbfKtS
RQgw0vSMifiQb2rqSuRtmXF2lUEkKIx5ZQ5sdN9dX1BfxZOAsgOFMkC6Jc/5sHjXz9wJF8nYjaVR
VIuS3F1WLl1fNEzM0q5fbbN/z/o++S+oCi8YoQmaY3sJ0ujiywhsrdC4P+p0G7wN1BZDmgssegxp
nVc7lw8hnbqPd47Ovg1Jfv3WzQ7ib0ZymM9J0UWBBQiy85LZofdeMVxlkDvjmyJIBugkXONyZzSq
gSca++fzwA1YKqcRpXv2MLZ60IlmBLggDkCa4KpXVIFrCb6/tj8UOtYtRK8019Q6roXDMtJ9F0/3
3CxGci+uhbZW2d5afWuaDhTP2+grL1pMGEmb8lvkRdpln5z03LkadnIEQf2jCdR+2BzSK+XqavAJ
QIY/2URZYkUDZc2VSCuett5jk7Mc8TMuYwyCEEwpD+NT0CfdrMOMKJD20DgoxPGdkfFl7zxPk1en
+AyEVQTLPUhf0+j0iq6R/MqTzYUCHYoC1iHkmypY228iB+9A4Z9m/0oRiJ9ByMMCiSef9YZr8dr/
YJfrLELUrFqh8UU3EVBYBXDCZKNksiWzG5QKzVUJaW5bWL6NTI/DLibtbT/fXjyIgN/kU7mO9uiB
/lcXEU5fUTHP6DsN6t7enckWEzLKvkh3L+L7yZwP9xWSj8+pHu4bk6Fj35GPh2iiQaMoBMPQS4RM
06eqy4qUdE/dfteqn9iIjIIVneiOwlZ/bgeVsKyGKgQW3Bcm24iFEtmdIiYjtKwD+wi50aKAB61a
YznFYsmXrYwEFWaoNmKFavC9gCIHB+DpiOf3kO+ad8zGz4Lh2HqRsB5ZRkUL1uq4c/NNIXY9OAOQ
/DAYCfiaxho3XkKgzbbkovFvPY8/86qx3h/OmfbxpA6MPtMeO6dnSBhD5GCcaSdbPeMw2XKd/eCv
8w/Q2UzJ5DldxEmrjv7bTaqZpLiSCIhw+xDRzJWmcbYsPwVUlKw06tcgDm9lREQpMHUaV69Hs+kO
Qi2nwuQrbCqxJ3dYFuidVnMB+2q3cr6cDR6hipQw/TX6WQkwaN09+RY4s182xIhQC50YdWqbo3nz
5ArzjGkOHuZlpKENaCIm7/BqvBe+iqMhHcWi6QbI7c1OJ6Z9yL+40/4vTPg02LNToYdJpvh4kv6R
silOuDAAbAZMdVXGxcdojyj0aqtgEUM8F4S6k6d6XE4NGArxar9pLToFzswYXZUEj0uFOXsUm8aH
0uZCAw7eAjYr/RJNyvlRTc3ovzFS3C7YxRrib1THOi1BCyRe93aynjIaA8X4W54j4s0bfj5h/5HO
1OtwoFk/u9+3g+OnoN+51kc9m4XXki5E9e4jMd6TuRuDvlrIaOouPESToHLPXdqOHTP+5fMLTH+2
7ZjfrVAEO/JQ4T80eOQM8zh7/2DSW9O6S7nymllgKr0Pg3Nhbm6yRlPutJJMCzNf1r+e8ThHiYoe
YUOVIO0++skIsuq3qqGYaww05SP+62mFWpKXr0g+oM4A0rZPjloRvoci7VF8LPJlNs2y0I6DSkuZ
35Z9ExwceBZaFJnJtcBdRwqsnQQQKHBsgka8JtAaSAufGhE6hm9ee+pt1OPjh+MOyyV1CmUgpVCq
pWLZyQhvo5wOFk9Y7VGGjliSH0KqdtwXzrZjuRPDbb2YA3qat6GrXVfNUPjrndLMxFNbA/f8IMim
DbcFA171c4aCDztoLd+aaZdOZzWiWvlsfQ+7/CvGSkKajWxpCIciLANNJD9BKJwHziiQD99ECAdc
+nHLaoQnc6Z5+m5abDwNx12koQ30a7cbP5ZXBGIhaM0Z/8LylKw5euUv2Rliumu4rWS615LKY/A7
rbl795ik0FCeMkKK3MM4jodgjrT4xaWtgILkhWaYG4g9NNMX0sIwPgBTKpzkgGdvO4958gWsLePA
0X6WqzBr99nblR56oQASnuzkYlb+JdD30dx66LFRNKM01MHMRA6S51sIIuNguZB1293r2eoIJQf1
Pauw7JadGUlMTNzD3cHfzf5QFIeFE67hhLdFs8rLH1QtbCpkCXJCwV/OybrwP4IlHqbpS9ZPzm9I
TFQ2DnRVJ9iXn/6HGw39uZ1xeSNqDxx5hfsF/wzh7neLSVy1Tcjy5NHWod4GATnXxUMnxmOwiHiI
szDmRYqxII7S2neJxlLJ90/6LbUwpqtMnSwtDE2knvCePXqw4FGEMYOzHm1uktyGY31ejhmZqT0x
y0tIWTJwjLW/0hJCaZLVZl7TTaLhfFy0pTCt8BL/XriVGIzKEIGt1D96bTXYILecidP54PUgVnBm
gc3201Ki74UCnt7v6x2F1Yjmj230fSt3e98dJmqwyMVmdUg1s7JHD1Zj2cf/eycwI763CTSUPsSD
ucFuhEXoxiB98osH6H4nQmVcJRKX92+CbrVn/fM45PiPekOQ7utza6ISVS8s7xheRK+UqARr99/m
hRwIETvPZtuTakaqB6aVd32lp43q5E2kmNzxKXNyU8SBaaGXfu3SVgovJhZO/h0y8i1/C45lrVX7
33N2Al6bY28wobLD4VLdgoJJnBQ0++KGFHtJe51Qfytojp/s/s3ZTkeKeMPW9uYJwRtP+vWTLwIE
+bgTfolHs8n4eHmlLGiiceBLu3maEaOJuwQ+U6v/efzjHJrObpOEZ47NWqtV897GAyw2hMnCEyrf
QM6LtbQ8hy6Z0DIufntXh/KM+evYLZBYVwQ95qDseeE3DLK5GcIN7crJ22FqQpoll/yXNEE6l6LM
fs90ITCYh4YBu+hDVcPHqQwZEM8AOZ6DawyJa+jsGAzoRY8UJ1bKCsLjIjcmGdrCUKbmAJvJd5BL
/CQE52yCAPindszCErM8lqkamxXzCiWUV95M+IQB4njNvKHx4H8ZCbwLVC7l7QDYa99hWF04pntv
HBzmIbAxDLAs1oQaDCKy8DEs/NHjcjPQvdqacBdnXBwu7hW3RV0NAueNW6P2g7O6fOgTONSFtsfL
1ReLJI+WaRf3M2n5/h78tisx7lHlj/UdW5qqbHRrERcsgaeqim9TjuMg+i9wvVB8PvrvOSOu5zUK
hIs3Cq16TcOrIDJDKS/iqnbDcP4/QTkRrM2JQab+wq0t9dTzBjaPzdzsKPawZczqy3mh9uIqHASe
e3HSdT2E1DfVlzphuhRHgqEersDbG/3JFiux58izQ+lB6LvMqXZl+d6MRPG25rRyrk+bb9/yIbnP
J4/wHYtNklwymTI+eYWBe8tL6KBWEj8yFGbXrQUqcVlp/MzHsnYG4kwbao9knub6qI4GkSR12LpP
8dsG/iGSCsSI4DAcv/c/Wf04iyEuisBBhOURBMvaSi1Dmp3z89T6gYKloI1LY47UhrYE7TQvZbGP
yv8Gr+rz+f4GZbilov7a0H85k624KaOIUvoWJLRvMB2BUsK7Sv0gTr1kbJSmInZ7YENIeKfUmyS9
5QEPuzKqZfVlePQ8appvgoQrHynTPpHrC4Se2EyfLY0AZl5vufBGdvqm173unF9mhYUftCcyvKi/
kvSkESj5Ixm0icu4E/149XLCmCcmfRd/O3HL57ZIzwpAD63/tuuXHRJSAGuLQ19YROpfkm3BVdqY
1ahuUx/6WRdKa+gyaYbSynQOFMEmKS5GPH8REQVB2G1p/yAz8h0XAoLBwBMPWamBpq5SlFldZDsI
pb4G4wpWzFs8sJJv7MZOZfcLmqz6bmD+jT553VHq8OnTrRRg96ONLbqlk2cz+E0UmnHQX77OzV+k
1R6d/WmPvt1yz7OsNEOk1UCBOGxzp0rk8pX0e6MusiGszxTPhaxyymNiCNONOTXUKoIJ5MXr4A1Z
duRYRxbihZ5EYtjdwdxXEFZppwoa7tUkb6aqVFF8xMO3QUi5R/7AcCr/PaYWgV3Drm+oCOvCZqDU
q3VnDnC19uGM/HPGnL01/7iotmi59z1gYeCZMWh8tFRS48e11t1YzZ4+ZRExxiJ+9PcDOwT0O0tZ
3jPS8VBpaL5a2FNpMdRwNEX15MpSiHLW6KoEUdKs2D54+TIxPSHVQ3NkZ0IRQITDG7BLyhUhpwHy
hvkd2NGMFvuaGYVUkSuG/wIc5QC+D2W3By5m2K7upkO/QMtVQ9fx6fEZb935zDipjkab3PakmP4M
CJnMpwlU/pSQYSnffIQ01fO2XJ1UVQcxvENOu7oD6HlKjJpt46l9w2oG/GE83SRkN1hZBIn9SOYQ
Wp7kKvMzEydAG5r3dxuKi4pZjplyN4OImsmmIC5qi0Ih0Q66zzEUdGQjrrY2f2EjyJyfHXeOHwpX
6XB6A2yPjb6lx1kDl+Js0xDMnV9JQW7zDUXvwPIM6HYw/3961Xlkr6LBqVFHvwyc8G6sly7jSXC8
oHRDbafZEJrGo0aqq+H1Hx9AubzCONgfv6/HolMD1O9K+43ulAVnuYszgT12alv4MuWQytABPVQO
fvhnbtg//tPRvfZ3FBqE0atlAV4BogvqY2cD3p5HhesVJxGHUN9Ec3tnhbO8S+1Uw/VkTzVrLfD5
1nONK75HOYnMOpk72fAzpDRsNi47v50/IRwBnLH60QzgsVdjXBf2nYZnDQsNcgzHL7F2DPpiNber
ZkFO/GXy0dcyCunP5jUgCT1SgkD48AiqA3YxGXSQikMFNqvXmc7aJA94rWlPobYAuSLwxMHxC+8T
S/iFtFYPb3DVNdnwkxT8UE27dypWIblrjS10korFUP4MApYrr5tKq93oAs5tDL3O3KAjaRdw9x2V
dOa00qncHxEzhjSZCgu+1pmxI2c88QNtRq+rlIkfIcICxT/1tWR/mNfFLTzMFvPsRIPcRTLuLKZD
5xcjjABSCaZIK7jjpB+N93h1HDpjF85Jr0O47XvvlN+kO10PCu7WozxZMWIN54Kbc9zGN6VSzk72
tHNausCUGk/3amqE/gnrLDYIHLN+EcSv1g60ro87Kidj15jG/nbzsBWq2ZqhAe8diDhbhtlofNC1
E/emTzexvHARp6j1THdatDlgE+kHA7ZxVAymcyEXRz2lUZTPePPemjW9LvQaLjkUQ9+cMMJDMeeM
qUp172K6sxtfPfBloi6k9oXHTZg0Te6KZgJlKChu/DGPN/PvuqbSqg+klDf/Y1R3J1/XIgnut7eE
lWL8NLMdpawZgPgPnovdcs00BgLvJ6UhT5mLceR5EQoOnHXC/AUTByYgVeRIo4B6Xoz2dxX97vgw
4lLNaTMCZevDauGU41qu8gx1iuNWzw1UPiAaOVn4jLOxekn4MICQi9M0TmM6lwsnBRvr7kMmhq2P
Gs2fDD6hur5+UCySm3p8qFiIkVFSpS6PqtsCUrykQPw4hy5TDwdXpcZIY+s/sQJ4ScJS5OK4ibCt
vkI+TYepj9xokbxRmF8emm0bm+kMUs0h19sHViyQ5LncYur7+J4RMmhMKV9h5HB18tuF0d+V6q+K
3LRbDBayxn6buqu4+1eGgDTRoHA5pvemLBTb06GSIHFKsLmOVXbvgbYNqpx/ZXPwRXJpG7WImuHs
LimQAMZsKDySxNSLlxzd/2xYjeJTIiblx2bvy4LYEbGmLb5MBgXTdQBSQsLAD+h6feeGGitdqkvb
ylgDeU4RNdJrULhkWb8+TpXevROjeCe7uxniJ2sFr1iA2gBHzpRshJZdz0/eoLvvc7DMnB/A+wjO
1f9xrPN8F2Pm5bQCLm+mepFeJK23xUDHERWZgyDNFNld9XxUbu/HpljzVkXP0OcdgIkPf+fi3nF9
Cczf4ZtKXkdyzeAAi06fx1KXij6nXRI48InG4/YpmVF7wSIrlqVG4ij7ZohS2ZN+ZA4+Thf473Ox
/FAunMcoW0x5eP+XX1EWQl18wBa3VPs+Q/ZxWAAH7SJUqUBj7kzDUe/H2Za1y7++5x2KmHtlOOgn
CwlO4vlnznh0BLZvbox1RHv6U8tuYTCbhNbBLL1QeCmSf01krWWxXgvfmSTDsFO1scHrrq8f2YrA
UfbT+6lxvGo0GapywgsdlACjGgUKG+0Tpx9aTjIzw3SId30w8Ds6/LmT2ViwHCZbPHXrwGXMOsDS
iHi1ri3cMpqaIF7FaQeJuUXvbemLKVv72r6KnmczUE7D+u4r7qZHVB25Hvb3zj91ffssGrxUWkr8
2zHqTTOm+UjgbMkX8/8Go1lwwCyofsTTl7UnvkPDTroGQPykCeWgfe+1om6H3LLmsGMDB0nfdoXg
XmNbHAZ0bN4fhjFhTR0gBYxm3EcJ8I0H/gHr+tOsbjM2HIeXgPxGicda+MH9mY5+P3cxbtdYaDQz
vTPJYlbQTQOs+GkV6F0MpdkOHJN1x9UDj6X34qVAZwlbZwC25YkJZApsSTKUDI33pBy5JCxKG9qd
3YKlt0/DcbDqeBcDt8gnCLvz/aEm+/DThddcDu+lxl0TeH/Eq4T9XN4s0oXc6w3oZ2zeQba8Tu4i
Ps9HJR68nvh5S495qHHRjxFiAdVWbXpKa0kfSNN/mpkSyVRvF2BoArzJMskuE8PNREq7Bz6cTwMe
YQhGzdthEvn9Wk9gS0Gkw7Q4X+AeKpiEDa2bg+7AuG+icVFYy1WW7wj8No++iw/1aSIqwIK7jD7S
EiY8hxRSV76PbEOtHFsK3GeLCbXbbaNT6S8n8g+j1CBalNiJX9Gw4m8bY+CSOI74WuCWEud2+yQL
zwlzexJPVfwFLoC6bYta8pb/lz8WnMJ1SlAPQSGDrPHdwgVAXqpkrPmuoDJVnDMAYBU6T+hTUbT4
X/v/W7ZnU7rfqufTveme59l2bnO3+1zMS7CmYInv7+4/3F/ZsjPPJp/vvzypsM9/J3gRzlxc9uWS
shHO/cwVErvLRAvkVe6XpA7UAyZDGmutXK8aC1RwfDg2jm4GzyegUTTn1aPimIBF5qqsmT+2GjLZ
wR6BRaAE7NaGvpYbKflJzhnFSjU3USfrb8nl8Shr4vLeuWErqNbSX1izfXqyha6NI9UMsBaHR2C7
S6fxcp3Y6/l+fA+J+FIqEtnsDP+6newpUl6zKUNAo+Fg5WuOC0GUoQSzho0Gq6t9w5243y8emQwK
gXcj/GqKTjOny00z2MVBTN4dCHVK/kkAPBbRMYIYgoKESCjLvWY6+K4qUZiS/BpG9mBNvZZY96vc
eRX6n0ftnSfScsmjbCWv0V6h8lDjScBYQsm6teZF+47wt/WwlhYxlnYwJFWD1XwyAmT4ZOvXYonc
kJd/s9JstsQnnxPBEoeuqOPi6bIw/9Ge2LiEj8atNtv7/WArcTDE6EnrRGniZKkv0U6m/SoEZOAI
7F7bUNV4/4UNQPhR2rz2Ft4mrTJ8j90WJNgb3m0FnWenfimQFec3UEKXylH4ZYn+qP6YnvIMdy4K
3qMPkrh0Eyohpe+rkUZXgfcpkZNDXU+aDy8klSx4UkDeROUk4ObsylQom51g97SaqSUKgwLHj8oI
zha76OXwyXdv70UzGXqSCF+LxVQ7McSR3ZAuygDOyShlX8OObT4x5VZQJFLTFPqsDDkFeniR5Lab
c1Z1X0TdrPLXZmu0wOcNFd4w3QEu1LxVKl/92UpEQ8Zjm8p5B8TKAHIL6VOb9BhNqEiqFrgZuTdr
ZxtbnNi0viYHGePep7Yqjz+RE7npIVlnlW145vh8GgtPst+OIROirv06rYOsR7Zv+HXVBQnji1g4
Tx6XWB9/0hJD8goEN9Q6v3PyvtdOW+e47mtVEPyoQeBzywEGpvE6CUuT6IqJvbg3ghDo8gZnizH8
XUNTjXvKiYohauj2H8rpqpGA7Rzwj8eBAuPFMYmKj7JIU7POQJoTYklqmRGDZRJj8GDug4v8r9jB
4+pdEI7ALbMVCfnCKzmbSlTr6pfbSYUicgaLOo9/XeauaQ6/Up0XPiu2wWPYAMo4So1/Sd1RJMCV
YSVhhODihCfe6L6UCkfXaeGCMrBvziKPI6IpexGwRxHwUkdz6wjI2O99lS31AiAfNkuQvII7tnqD
hBmNLRpqv3wBB+4eASe1AYNWmnGRes3I0SA+zfhkC5KOEzDAzxDmmKPGRsgxP6S7EP4vlTx8QIMb
+7GuVkhVuwUZNqJjf6v62rqpddGTWOxTm39NxKm4QyLn9Nx8uXUL/T5Izcgg/tJsMAiNkIOY9glE
gG9n4YhZUT86iubcC+47CtbUJi0koeF9j3xMidI6Uf0VPoeA9b+P+fwtSTVOpKWvP1gUKMwxEg3n
dEkC3ocMZruMooRm75w9FlSZXzIbn8y+NjzXMdli3VE4FoTiaTH5j7LY+zTuudxCEbGhi3Wr2w7A
4FafXUCnsr22tDNxcgr8IjwTTuzJHcsGq+BBEzsFM6kk229/rQbUCHLN029IR96njBhuTbn2/0s6
9cUotBKXWzP0bAa+mdt6jgcRKG0FuJL94Jox5Z3L7jsAqiZLmLumGUrefL3UUFbacn9RJGlDmn16
j8isIQW1RLrtujpnfoTEYavAKJUW4YVhVii5ja+Q1LX/9FFKSLYXrtCQ/dOgquEhjzcJQMluDTIU
AYzf2om0+z9z2Z1lIVBL2gAbyOERMhWuk68aF/VaAKztvhvuiP3bIIlpBlnhsn5YeybdPZkwBRaZ
+hxMlFt5Ew08RwG+XhuJUFn+qe6n3/mdfy/nmSBU3Nq1Y5KbpumJ5V24ZLMuS6iv+d5H6PA3GBbb
zvBeT+NnMQTUyOeHX/1AnPwfGAb7wyL8xJYjlBicFLT3T2seERSS4m/GPVoF6igDGF96exb/jOti
ICAU8UHoJwnfCsb+PkbIx/+X4LeKfMypdlEXXVLVGGB5n/xY5TrhSOsU5Owgn/t+Kcqf51B5JfDO
VZt0wjI/ntJZlID7uqS7xAKuEKTdSmrd2Su3k5ckrbBX1QPXKEi0xl3H2G4ezD8kKMNHQM4bcRbt
+Z5+Sb5sDy8cOwC3oA3uEv6tFjXJXleacpiD+V8Mll1DJpMWaiK7G+ThR+J3i7wZcvzkXKb+dFij
COhE3HHdL4m+7YifN53h/YDrlDJOxm/xkmNPNJD+TWrtaSZBS6OCqMIrSZl4DucIwYF2UC02yc8H
6AyUOIyoSmDs3rjgRFf8ZkLY6olpPtUyALrMJgZYFPZTT5DMT7FtvPi2TVdf/+di+EM+o+lM7MaC
9Wmam1WXsr3yu7fGSdmQbTsMMLYusjhyRbzDfCyb0Eca/+tY4tX7xw7hY7Ayf/hbBGreJGqU48Ti
7/X5hXLb/Pull6/Rxxgko3+SdN1GchZUGMXH0jm9FDdmhXGvjfbvFfic1bJriGxkWe+xzAqIS8IJ
M3WFibM65Qzbj5xQ7mG5hiR5esam7xfT0UCQVgnB6OhhjQT6RxAaxW1dbx3GrYEoeO6dn63Dving
sIgpmwnb43Hn/0yLtTm2Oebu4E1BQmxeUus9Ed9oXChCC8hD7q/4OzTpjFZLBcWP4ph1EAZxVUl4
hria6qJ8yp2IQV/C6N6lhi7TwoxKQVYi+8tTl8T/JhCxkqQ13uTPmFb0ZQ4qh+/GzMTn3FcPZrEO
jGNhXsf4QSIjOjnf+JDJuHMllwuuSWd4c5xM8nIjbxsEsHwFjto8Msm3EMowt7jA1QhgvxOKxNgh
84SUL5pAzA1paNkFpIQXjAdM+/JPmEbMVz3PljbTUyXbdLv8kP506j3Eq3317LuZMfrlMHs5Pt4S
e+g0XjJ5PC37JIlhDvSJuRBvyn9pmi5HINY1qEt7JuBDUdTmRFR1SYVtmJLvzHGIOsZU/IZPr2jU
pKc5NIRdGvViT51f98r4khOMha6AFoKYBMkpr/WgxYvfmFbhPQJoBN4ip1zimFB9aNghwhI+n7ly
QZb9ZChqUkCqkB2vjhO32Z4EAbmAoJEUJYijPK1hxNnVLJBW9w38vLgNJdxtiqFVRQzyJVYW5PMp
6ubEMHbfZNJimywXKNfPrLkkDLlh6XHBkqLN7oiBhkgcwac7yHPDRfGsv7nayM5n+mU8BhNmx5V7
VNQrVtZ7ggKLj0iefqsAm6S/RIJrHpeyHhx8gQkD0l7tKpT8oz1VL5e+ZRCKh2Rw7t6AZ5TiPo+C
f5dcxLcWNpIhowZEQIY5lmdOWtrlUx+T83T1PmeHVtb1JALjxskJPKuH1VSPEoCnq2RzeIFzV5jt
qifDo2l4EcQHCvNG2SHT7TaQGxfJN7blVjIqh3OvDdUYj7GkL5lq+SjBswJzMpb3kcNW6xuuXEue
+CXm86Hh9Hg1StXwEM4tXDUIu/JBcgGdxP7YoIRuYExEpE7muPlScI3v19JuzcYJx8o+PORKEESD
YLiDL8s0bZBGMSs3mtbjVdn3jkO1SMOvMV0bsr+m3cy2zLg4Qo4yaPCOS06so+KqQmVpqIlIh8Dm
adNNG8lqDXg0w7vgUYyUPDuWZ0kKXyNpeFf0Gma6v+7jVyN2ofgC5SqEBE3bmRQu33QU9H0iDlJP
VgQViKqNGQ3Xz18rjywtxrpIIPWOQYyH5nMGhNyg11jaVI7D810fbKxuh0NHwJRoXPQjgPC2C91h
AXBs9XNJiH1tCEHc/8hq+7N09vUizH67HxKgSNUMggdPEVsnXcXOUq8lhEgSfB8p8Jts3ZF3rt5j
uZ+6br9lU+N5MmRtyiaOUP1TyHU6iPYcerOLXM7UVTGDTlVeCPjMLCBPi9Fufm7QmtjR1iv1mnXm
KyNpeqiI2KDen5OHRGObn/KXusLH3S4SX9HXZQkchejGO0QY14oR2dbh+ULrAVZM0AMRCAe/Dr2K
TYJcYJfUGfMxb1ggul0PLmjBgzAyp6i6QF2cWsbLiun16dXRE5hGix0GR+k7XRKnVfK9+SN7Tyr3
o0tOG/xlipkFLxidKtZQYDXAN50fdqoy/t4qQIUuJsj5W9GrhN1cuLYXgtH0CFEoX5CSupIB+9cC
zQLEGPQw6Bl5JcMBZK4C3fK5hfa8vxRYwGMKf+wqxt0f79VTOyCOMB3fQW6cBpOueGz/oShO/YX+
dYNaBKzns9uoBTmHR/YfMhAmtr/UjWvxqnKb0uBX486tOXsw4K9L7mr31eDRCkp+XZ4RM3LPQMgs
UMNoiKPrrfATcVx8nHh7bFtZUmlsnmQa2yzcMs0j4hMeby1tWTQ7yuYU9d+iBhl5KwRU2ieeCHlG
Hx4oVh0xzEpPDf+w9MFGCBpfbmKdtQ4R/BnxSeOv0QPMUILfFx2g7w1Pi+z6kAjIx4dqXuzFf8cc
NZvvNxEDqqx2MBbnPnWTTXXTESSeheGCKrWNHKoYjcFrKFHnbL4lpZHAx/z2EUhi4LsNOk6ONCRq
CYpY8tR6jtO+AiLjcNeFbT96gOxw1renmkiVAq+3f2Qtt/eeuEg3DAPUrHib5/LOHYdTfNMivAKS
tE3DbUd3EmW9ZfoJg14EOQPVE17fM9NPnd2GnLyfRef4hDPmkBLRHUpMWtaL+T/K4edCx8gm1xM7
8AkdHQfnUg5dVkefI0TORE5sBuuxF6SsDXf0oQ0xW+aqm5BIPZzdYWjJGtVmFyq+l6hevZGaojJD
nSTrY77XJ6dv25gOZTM5e9hCgurbEFm6snCLUpY3EpRGzY8m2gHOh5ZSoIGcu53bfxy2sTFERANq
BKxbH0RmJ+om+rvVfLvGflpWziRVvSTpCxoKD9ZtkF+DetuFS4wqz9oDlBZKstb9yjllM32deirU
7YSG0vwnjDP548jMajT+K+ZXWJoTP885es9b67TOMCPJIwtVJ/iVOh5zdHp/r7fIQ5odooGdqnsE
Hxp9z+fz7rWETB1R0cjbJcW8s9W+a2mu2w65UkICAjJSJQ576X3qBNWgcDx1dVA5Rvz/w/BQq29E
xJ9IpZ7Uwi5kbCJGCV5jPF8l01p+eUszIQE7h1F8Muc3HXOMTXeABA1ykylQ6OrQTmWJ6xXLFs90
AYYR4uo8RIuYE6RhD7bxMWMXlWbyzlxj34DuBnsx3ruUpH0QRAmXoLmqXz5cqiRi7QGUWR/z96Bi
GEjKstCRPkMDXTyeg+V5eQh7PI+S3FQth5g0D5/CLNBs1n7h/g4aCOErgUn3nLxm0i+5w4NffYNl
g8zuN08VmL1EbNAM65wecqiMQ1LC6pepQVOaxu2RdNC7gC3SnT8CqE6BD6UMcmOeHWNb7oD4nNtY
aE22PO2ejXRdpeZh6b5pcdEDItYhi62nin4Zp3zPvZf/GLs8Rs4Z32vM9SwiJmmchcks+C1F1771
K1XI8ONjsnUG0u7kkDsL5gM1QSXVw9OGRigBvw6SRdSGtM/T5NeHVvGE4k3sDuQWTWCkU0+rVnmu
IbLfVLtj+u9zXkjxM6QITj8tU4TlwpF5n8Xwm+QRXX4Jd5Yo3osNzSUTRQAuiM8CIYPwoU8zfRPM
M47aTq0Z8b3IF9enSMarOqBpcpaS5pU5kWJ3JLlpOIW9PrhC75/mxt8+rcTwzSMhBWyxQPy+fscp
XUsGzgOr+NVxBNfbmHSOsNbRkvAtkz37+m+4bm9kbAdZOJ+TrC0yklSrHR40XBLjHONyqwrul2VY
fFGgL7LByT0lbNE5qGI0MHzJA57EfHxxcnWhb1eNQodXycSsO1C3nvZzopuz18Ebxsp6r5Son4Iz
PHaO6FnwPi2ZYREKd7p+xTX/1fpxwA3DllZU0/meKvNOzenOpt6AOH4+HxVmUkbLyWZl0fYaS9DG
49c6ent6RlRgzoWwOmqkvrOrReE8GbpdDehMIeXe1O/0RCnmhC1USKuP1cfQV5nDB90Ed4H/xR3n
JgzzaClCCvYDnpqTAeRDjaoswgR32FXQduSB5pb1iAdEuYUN/NJXYTs7X7degSd1uGFdNXdVZ2Vb
cZuc7TUMrSYF2/ogfO7YimLuoiYFWKw7ywBIa3nC4O0lB6JZCwA4s7QfVnQz4IfqGzZu5Nzo5B3j
ZEjyuQ2ljT+hyW+ASfN82PJnuncLR7Z/gvtRQukegVUNd5WM++5KQaEw2VRe+sIFy7C4fIed0MuH
8jrvGKzby0IBJsqoMtshhMSsmo5WSev6Zz/frxvMolHhybWeXYUnmt9Y6FmDA0AhdZPWtORGQR5Y
vCJDVSl46PcwqZUb61zJpDKLxUfES3a2jN+1LUQ5rwhrsyGMiYh2+VQm6ScGp/rynImeh4cecV7u
5SCxv8pVFrdfagKVsS38OHnln35lICqipUMiLuYieX77TR4q0qgMAWXj6IPGsrFqcejDEbcqhoQt
pyRclUAMstCDGoGg2Qg/tEsS+yv5j8BDmiiMJD1s5w1rQaWxAsiofflG98OXUFm9odSlaGccw3cN
85aukWrpLcBcxP8dVqRn4zcuoF3O4TxJQLx+nfUcXhaFWkeIBYGEzH+pAb+Fu1+fdfwjnFyJaAo4
Zer32Hp55mwoPx+zJOZcvJYQfpj9qto/D/KKK1rW6wv8EShwtIbcD3lcq5C8+m08HpEpIAMM+XeV
IhNLGB5wYGcKKRvq+zvzBgmYCEUxo1SY2k47vN3UznJyEWVHQGCGLOibq6PdKgrRb+NNhorahXng
IY0ZxHouCCN/4aRr1VVrIJ9lus9Uk2hhBwzzFnevqvRskcyYO2AA2svnI8vnRTE1IkFU717Uv6ZD
2NuwF7d0wzY5ayTF2vqZf62SG4F9PUF7iKygwLY43c8j1jX1jT907vmyV0va+wLONQn57eVOqMqT
T/Rg9c6o4ZsjUMqnQL0Erw+ZfRVnp/RYWaETmGKtHh7TwNW1N1PqVnd3Tha4UJGvZ4YK7PAg3HoF
ZITRxh0N1lOc5e4oPDqsk8p1nMLwrxs4iZh75V3OQoRpxhcIrtIqoT3uE21paLV1ccilXsS9Buc9
MOK/1bhYNhY/5j49I3SziLvOUjVl/66D85IinmmiwLEr/OXWjOa+gtyHheLQJQEs0Mvp3/poh8Rw
p+uB/NVB3JsQwH4BnPcbn543IT2oRt9iqRiyUr+kverO48xspn3EGtVXbyi/QuEhB1kfHEfICKGo
8+OaXRWLy/CVg2UY3sstWYYw8131Ygdruyin42Dro6wtkJBPWwRllgkhojoK+rJsvbAet2mM6hTJ
yfP+ZZM2Ex1AjdRqXIGu5RtPVbR5K9X/0ezUgrOj5/fyG2jZYNPil1NsnRnD8TdD7vsgW2fcdMao
CnrQNbFvtddwPhYNP5GwG3yvCnLcwf+P2qSo1CWHXi4UuoG5IdZgN/d/PPALG6v+C81GkgD8QqMB
/7oAwTYJYsDcJ/TO3x4pCPYZw1IqfyR30wrnwak0o6kGJR7SEKaufv3hnU6NoE35D8ZANp30I7gM
0HHVR8RCNADg0mwxdJNVIv7rO4Fy38wS+tYSDQIci9skUFZtR1CvvXPq29Vx5wjsIIg5hJgjsCm7
mzh7JcTVfdL6VK1+Sh0+9sJa8CAWoFpTf49S0ePjbmtXRDvanSMv1QJwromfcf6KndgtXEwU+jnf
x0SPmY/X5pbKKchirikwECYVuGa6kTHlMxD/WoX+lc7u4BgAXehcudIvHz19wwIuzv7ISge4jAVG
SpciqokK5rgZ4ZYznZ/RDb8jgT3xqEpW9ZML0hVdFKmVpacuXHLR9Rq/uDbqJQwKB1eTGX2j/vnG
VhEN30oFOoG/PLv8Y52OsfUJUMNUQSrfaCyZ2IV9BP20868x/8yAXcjt5RuJFtiUNucg7fCH9TKb
JjSi2PMgr24BY81tjQgistIRdMa8sPSo7/0M8W6Bnuo/hvygTA4vUI2kC9Yty4eAAr0V66AAvl20
VzfMSnI9Anb6cIN0lLXUWPx56raA0cIzeXdPRripw5f9jOwwRFiu5pYgHWo+BQWF+bep7gbCPZst
mzAiKgczIGTFkM7P5yVHhkeUN+ZXoxvLaQPB0Wo6eEj4oftkZtM7/m3mNjhx1To9a4VAAKWqfLdi
wCFC5jKmzf8RVwsKy2prki2goPPb6tZa3/2h55j15Z+5ysXPQ3maCyyji4KWwGQDqbjbVVdFRvW3
9ud6Ez9KC5lHY/M2C4mRN3CbpU9rwHLlRWJ5HjqNTUdhHzMygP0zYqE6t6ugNC6MByTgr1vCYfdy
ia3idlw7QnbKv+ADZIB89Gbj0D8+7pU4DYA41AeI56xbQhe2OeuV1qtTXRJ4yRVdyvIggYrPjwdA
6H/qj8DUteyUs+ubn7fAdoW7AgB8exQqehNbN9Qk1Ta8oUGBDQGgj/B+vScQpNfdfYtXNZtkoVfa
IAarSIzsDMT/q5HGZZgBYc09/dpsSkYTXMiomM698fsWdTnyK6bQ2gJUc58N52uJYELLMdSV2mTH
839tYraJWTkdC+/7YdFknPQYftDqYX3UCJjafg5PWUZ0AP2t8XqLLO6jyG56Ssf/P726VqxIVXJU
KKd2dTKU+wxEh1kedW32NY14emDosY2XlxBrsrXbGSQStWwwpP8pBIUFZNx9CQw07FA+Lhs/MvAz
kj+Uqu4MAae57ZH7+/BDweC+nB/kIRQR+zAL7VO8GcSMRYak384j0jJszx2I6IRBbdDdMq58WgqY
kQXuqbW3cPecKUAg2Msrq9pWDwmZz4QvptWevRG2ZOOXToTq8MTfiUlb+DLD8Jr92dTqrVMmqW+9
wp3zZLG64PpiQyWD10zb+74NCf8AsPmaJQRb4x0ra3BXtRcXcdGzXmydtBF36sK/MD50sg+I7Egk
kemqT0BcKMFIrHm7UuRARIj4kYSXS3JpU+mY0y4ccji32PxzdmoTRBbd57SN0pE+vge8nSpJ2HP7
UpmEC1Nsrp4eYDYeE9n/f+ZuY6bKVhkh8RH/dToyXUJV7Z1IAyqwgi9meVaHH5slmwsMKDSAirn+
4iKsoXBAy9CHJZyXSKsp7mhUJ+wWi9eu6lold0+6wys/FB3cq19uEM77ng2ult8/VcucRDIsFqdn
RMAlyAAlRla0ruo2aivs0ExkaXFlwgKj+KeNtq9ZPUAhIPl1L7OLAIbttBe7cqR4O38PsnacElVz
ya8zFxQrtccZMrmUP9feGt2e6J5nEsGcM8qRGv8FYqMnC7dSqgU6DX+T2gumZAmCQtxtt6IiD6n0
6ty2aFb2AjtRdNf4akefy2wJ/OT5WO6SILW3uFH08HbVREf8AAI+Jkeq8Je3caZnBr6w+nCyIcUe
e8zmac2djSBK4AfVM+yjwTOi9AZ8CTMdeunBcxr6FOwYyOtnB1RaFDkNj3Q4/ESCdzWSEt3mq0sg
SBvLKBynFqBwxJgyxeIEcw4qtlxL5LRV1nr7xV8MGQIjfOcHQjh+OKuTNePQYh1o8UTk1VhGAChz
OMqahhtzCw8YY0hVZEsEVj+xskUcAsKsdumKcGMtWkqExNoLFVkjQ4B7+wD7gcsyxAVXQmNBpZip
NVvPDxbkMEVJJFcYChUg06tuWQU47LHoAzXHQ3ymxK7BXYXverpESSNZVK/VBM6njdE99jkUEg2q
+/GoIv5/npbIxTX1/fIlHiHE550H8hIQWWvBcSDMfxgr0HpSEVyH4ZxFb5v0nbJTBVFvPNHDAQ7O
k0ORC9mOg2N9f+a0TRDl2vEN+xTQuw6o7uGcAvJCWG1802+7bC80Nr9/4cGTDVdnMTYTyqGSUg5r
rfDbvKgXGLpb+8+Gu7pnahGj8rUhR4g4P22uilD1Vc2/VqN2weZhw4az1/xCzVYW8S6MExCMXC5R
TkOrl7pfyl0GmOKmgTvvDh3jx7KW1iA4+lExNLtDSF35zVtdg2soGWcjh/y7RhGMlxDykwCxEfSW
51FDfwzBX7WmdUccIl0B0NHBA1S1Rj2PYFd7yY9iqkCRJo1zicX/RC4I8wK7hc4OrtY7vgOfDsto
PEJen4jKcS0X9oqGFg7I6jng1jq0dxq3LtHL0GE2sFhEH0GsbK24upkbOvCk65wdWE6GgxH/qEFv
uMgMU3Zy6IDtJ90lTWf8EWY/3E2foe9Pw0RnrHH9msr/MXcZQRkpR+o9md44Zmw3s2+0W8y4ohXR
UG4ous17dqclqqT33x4Z1uL/yr5sLOrsbaU6xi/5LPPZ/BBnRop6F3HBKVV/akQii2Fqz34B4+mb
srj6MTqIrSGZJ0b1XQKxZ5q+3jdaawfQv7thmefoVvHJ6AZDKi7VNjMu93PvLrqcWV08DAC8Xsns
8ibxzNSsPcgWcFSO2xkcI0lPZAAuRuZhIQ0AC+LAM9WO11o42Sz1BZlu9PV9LiDnlhZwLwjTnw7R
+AJ55COoKIfS2CVBoPT9dYtaucIiMYClpMygJkNDId3CMUDd9rlFb6f9JsGD6UC3T423RWnVUd29
7+Gq3ECWphXte+rgAWopmNpvt8wtmbMKZ1gTkKjLIkq2tmQkcBboaO4JbutAV/aX2rrJIHx4FCvX
L0p+dR53wO9rbyp1yuv9kvsTWIGEGOr0hkcGxCtRmfprRpdPqd2i/w4TSXhIYqiuj7yLlvVzQas2
tnpiPAM544tVetE4wTp45blDbkziQSVyNDeniDfNB6Ud/PdkpHjPm1gjbaJX2Vqg2R21FHa8YzGp
X4KnkTRW763wmb3GwCC2fw88soK55BZhdK4QFX/prIlx3VKgTUWUONgyCphNc47LXp00nMbqaVtU
OzIwk6RE+OhwsBDWOdPVvRrGD7NNoWr1UVzchg2N2YHGCkR5ZhTyVXT6t1NxHDYh8FtYsuk5JhPq
V08iEXZzCnN9ZCF2ZsBZR9ELpw2/exO+WSzCRrDPnB88sWfw2XEvST9DVJr3SHGZI3GX8YOc7AFs
g2u56B4KMJFbKNCA90DEj3HGkamv1O+b+VpLFRvuUKgdG3matjFc8eJEApKtdUjPOX72pcMMpuS8
tiUHaefDPsCma9D0ubny27apJjAFxZ1LzKkWmqFRJG0ffwcjRo2nhPONcec2ueDY4S4LRCIc8aZJ
hl/KIUbnoaMAagZclO46m1OIUl/o4YWTxZT5k+NbbCcUVbuRS+KAHppE+JRRNQ0SnoBB2FBN00uz
eEeHvIdID5M7jaLcFSAN6XbZi7Iyaq+w+YqxWFBWnPq6r+9xPkybAOIqKjjWDpbg5jLlzd+4FrCI
ZXh06sE3jidOZCIhu26bHZwJ6yyAGqmxTtqfWZTl9fTJ2IZCcIUxT2ORT0vFxpsjtz0NsUxTJtmp
7GGeaZ8tYdktRfxTFZJcsgV+OEOa/rCJC4vN/WRtMBm++gS6BAMB9MVVEDhIBFNxA3M8kF7DxW1c
UZeR7xiz2jXGn8EOkwrtDPPq8PdgBykkgN+PWqqhX1xvWjKbWRy7lEh2EwmVlr5Alk5eVYnl82EZ
tSqeWaRpeBq8YXLS7EUZfO7poRul3pLM6eJ4YF2D2Lg2u1ULek6gdl1ehvuWhUS+MOQF8qBt0JtF
wd83VRt27CVZb5JKXonybLW/aU/FwHh87eQGqSn7JA7FHpf8xVXhSZwbkSyhj1OxzTAeE8x1BwQ4
IyHj2LQFDXm0oWJBwgbRDpMoGoztOB9ahCK5wsBafSY0JHp7iLW0Aq2Di0euAgsGeNzXKf+5FM5C
wOepR+xl0xkFlF4gaqZjcUL9hhigIsGN3ukrpd6LlIifXIiaz7PvEyQlR7vgjYc/po1MRyBH0t7q
XE2cN/hKi3x6R0gCgwvhB5qaQUaRAd0bTkcvX4hVJumMExc3mUKU2gyAsWQhImSAHVdrPiE1ZD7e
AqyzGNdF5gznkmn5HIu4zk8TAIOn0LTm5FOWg9Djh3yFdIRP4n/8E/TmJmDfwvXYu2qEfKvsuu65
ujzkMMPZ7lq0KxzIZmnp3p0c4HMofUBcMTp/IciFKMYN5cbehmhX8fOOWZP9vwJ6OqaqsVSyynQr
PfdpDT5vVvKLF+AzgscuOJhkk+WvB4Pd2eNDs6KAxtQe1/8SlBhi5hEN+8vrZ8Pczm91GCDzRP6W
SJFllN9/7Xxlphv8fP48XQ6uXTw5Jsw910mZMwfARlMFfgMhM2PkGU/g0QJ0KoesMYEFXaI3H+mt
FnDBfpnPyrcKP+blTOUVg2z3y3/hzyElvuA0c6SC0yjE8bQUDH6q5glBhK4pgrfSemgK2O/zgobx
dUq3I/XAsOXlgQo+ZaLze4bnsAT8mDemZgSeWJSYHJeDEXpu06XWqXg/VL60OE2eUhR9s5GJWz4h
dKyVlV0JKFoHz24rZtgfa7oT4rlsQN5q0NlpVuihDXRpTbxg8Pv1yDFx4u+7jAVIolTCPH13Ue/w
GI1MZiNW8wjlPH4qrld8Wg7mhVmVp+V8yknBp4KNwiRKrmv6ANaSVsKIgXbXjSLbAQwN/BMqTaDe
zQMBi52/PwkQIx8e8K/8T2FrPZeQKXbhMhyQbkzVnx1C4qb/FLjR3oG2YRy0raEokUzQKC+6bWWH
ae9hVn55w0yKkatqzROFZ7is6s13RODxLJsIdbp8W7pMfkUZIU6rGVnkTfJNtCBBBCFQVkDV/6pB
jtLL0o4kS/y6F3BkAWyrsF/BXaFM87qndVd3mo5tefUjsutGjdKbOhVzOAKeLpFa7N5UqkqgfqoO
zjEfnnLvk3Fwcfmq+cYLSOD/NfAqDGISF0PWpjRt3LX0+1u0txOztRqMMCH0udE6R9l+Bk0U5DQH
xYqZ0tgNgrMttWwod5iMLZEgUBH7X1pdQTtS3tEa4DCNVYna2M7bWuny3myjutH5GTD55IAWsR1b
dAykgqoeMSi6qVN9HSEeUAlV3NESaIcSQYWVuKff8AcdVx/az6Ouge0Cr8DbXKc6fbsrhUbtH092
ENjsfsAztQIlA4J7ZU4DLHU2LHF0w634GBJpSadWlijtGth2ZQneiGRN9K3bXM43yY5W4hVY6JpO
uAtsTg77OF5DN9LIvXeyX3aAuZ9gbCOQvIz7dclMUIBdBazBIh+fejZ3kJg28TVlIMPZ69G6GsN+
fdd5kz0beMkG4n5MPIkGvMOivkd5h9P4+m5TcYfCRP+XJ8IBfd69xKBer4+jl+PRSzOsFsh2+5bI
cpcWcWuWHEfHC0kSQY/xF1ioiBITPypouJkSSNLksgqFC0mfdC4XYmZeROLau3kkVzF3CVUU8xjC
BlgPO8+bCXclLRn5z6WcAcJZag8e9YdNhJX+qe1zIpl0+4oRM2jAFlmnK28I4RIqKG/Tpg/oJ1UD
KRJ4Zz5iyEGpQTdP/tgdHKgEZoyd5bP9iZ56xYYHwZfv5LhjH1MCOLLvJ82cUnkA4hiYrGsefgzc
MIQlP1C5ygt8cDAZFMFT3om58ibITk/f2he4p8Tm2GWUoRpsQT9aSdv2PCzrRdB5RIyJ8GWW5Rhq
q8rPvL4nGASH8Y0sA3jEx4jYhAt+Kabwv6QhPjDF+Ph4R5b4li+cHwrzrqezv7V8gfh5w6CF/FWU
Uv/eb/EJz7r2DumWcgYwUUExqFa/QSDV1+YiwHDtTpztpuwA+oucv2AogcQe3WrXrEYwNIqP61kH
oF2+TVrrH20RbcRzgLrk+X5MGKTrjJhA4+SaaoCrdqxpJ5RoW/2j57RTtlewA05s0HYR8IDq35MG
6sk45t+IWisBE1ZyQh3mzt32ALwQVOdbtLVdtz+eUsp92kqqx5rOfLVyzSZjSHPC8jwcVc4nYnRr
TFoqU/S7hw/KBdG+GuTdIDiqL+NyzUw/nkSoNdNP8p+3hkIb5X3GWdeJDEjJtQaEMmu0ikJtera1
llXskYDbzlumf0G0MjHEZ8IhHpPuqk/7HpLqBpwyZLy1AnHnJaUZjXDricvkaptzAc9jcimtBzBy
QkKaLYPsp/OvIdTjKyo8N+DL6RiKpztIGNOJPbSSP4cNY/2+i01WmOrTypGBSit1YpDu/JDuHAEl
JOguZ8gjfnibiAgMEkjMfVweOpbPXqA0Y2qisdqvmpdxSEctI1GjG15vMsNzklmrrCzJvzV35FO9
U/yQqqAOAxY6qfwJi0XmWL48GjY3dBRea0LQaC1xD7psIrlrKwbI2FlfOjrAJmDk2PpL6Zu9sz3X
4QPrF4F0Kf9AUBPkj8FLIR+H8bqg30+r3pNmw25RccqstfOg4xjc/gsntUCZjwNMZMtqjaj0proy
+4tAty2iYRyiF5vQu0HJ0YW1RZop0/Rzl4pq/NJ/8xrMx3iADKXkZnWhsv0pLdZvgwNPnY6r/LZ2
SpRv+lcjComkqahPq8d5y5P5F+CmvHd/1YHCWesjVB2Jt/rF1tMzg2HlLwjly8hlybb5hkHMmZWx
os+KgfJY+iZDOIChh0MM2BKr/pgZnykk/Gpc/5tVqae+jNDhwBGJyOtON9YfJ2ZEQ1lYkEITs+if
4XfLhkGC2+mhi5FlCQWtkH7PT/Yr4t9acU1B9TXnbZFpbDhsopmTiy7/XnkrXMpyVt7c7/VCzDI+
wGEIek0nW6fRTL/Y/ZJPZzv1GaVy2hLEhrx/PSVU4BD2eIYE2xK3TvKWaom4Dzusvjh9alTY8ZwZ
7fveFAQD6f1F43eZQsvNtlRReO2KKdiQIOOSXXZZxwZUc11u1nA0fSlPowzYQNN85IbbR8J5vPQf
pZf18I24XJqw5KpzkoFcUeShYlUhReVqi17sffeZfkT83irayEZq+jckK6zZjYQIdhRXEK3Kx3c7
kQKIkskkxZGFcEvyJ4K2SZsAJ9wXQgAGJ+v6N7UYV4HSiYEnOQfPLw61o5Oean95dlp65ZzcCmFz
ddPKbQK1+tw9XfgyPcrfjsCPhaR+vhIfsiGK51V8NcPhI10gp8lo2g7SiggHq7DzsrOxXbriSObe
U9AHID4IZfMiU87IRs3U7pEaYYwntGZRtYPuITwpcbJGf1u7j0ZAr2TmmI3Y6UkENBE1STH4ZThC
KBZZ26S4PfKc0yFM3TyNPMhG5NLGznSwcSagOih4hM8GA5pESy4P3kGCz7Es6J0Nu7yhBuMbO8SA
S39VD6bTfPhwrFgtcHtpCNLwZG6oNk8zmuJZ6QVBAdALEHM+zoHE6q4W21iltiEJIMhRo2KCozhT
UwFsykZL+8qA6JUKHDWwF2+eySqi4iVd9l7UrSJa8miUs/HlIVFz0hF07GKU++pOSvmjEXPJhOZs
JgzbcnCFkofkpvjFpvj3nHxLNH4dgwT7xoKr02voAIOftTM8xunoPMrsin5CzytkLUPfjE6JDtVX
yWxmXssu8XSxJFjbU9Qdd9rSe/wAFHElBfsyWjFSVSo+DUekZrM7GNkqHhkukK/XJxtxpVAhnVjY
+lSfkhBVbjECrpzLqsopVM/4CbOzVDSQyeHo+fC+0/7weoaDxIIqWWh9L1rI6kmThfM1Vz1ozFpB
+i7SAAbL1cgydtRwXmb0LcZNlDLIO08n/KrfNf0fTgX9BLU7iC2ZC2C3RCoqlf+44woEeIxzuB6q
9XoYCE3G5ZDMPm1oT+eo7VEp5dRSkbj7Gowkyb/yt6xMRk+CHsln/Je2ozxd8klu+K62kin6yC7f
oYpbIrUmxx509AR/VBUsMrXJ4jCPrhkCvz7O5nMv0GkIF/NQArfjVWI7wfuBmHYQQTPEQGD4cKX9
Z2bW6G2B/YqI6GfaujdxcoOU0tMZCtE1l4ExLIOcnuNw7oZykc5lZQ4vq9f7zVEz8ltPQz6BwUiR
7zSFVCaVzcotQ7Btqh8UBJfDVaDW+uTUPiQhOowWHS93lKPrWBqwz4y6m6i7ndzJWCHrfyXzZ+pR
IUo2LHvryn7kBa9whIZ5NaL5HJYDPwsar8BZPTkXGZAxrquiZNiHa+zsSm5t5EeLvtyzVngMLUi4
biHQl0Eq2vvifmgVb4tewi5w0hAoqzrmx2QNS5Bx1VTwM+3btvdak1YqCW90t/GrjSHGJWYWub6p
5AF6UewC4W+NlDa6wHG25GTUfTVacqFLyQBD/xI3oEws0gcKRH0IyRLHH9e+NSRc156WiSs6TJas
1/fCt+q9hJapo/97lR4+WnPZEGr+YQVDffVnWDGQdY8SqNuH5IPRNfvFKGX7PblIguuejjMl1z+D
PAM0U+sLC9EJZL35y979+3nyrquidmna4T5tqC/aOtSAgeY3/xPxK5rpSAVQLSB6J475tCS5cpBT
R6gqeh93ZU1X/H0QmBZLViRhR0aOKOzMfNm83pRfx/O8azvMKIiEBATtRHTnXHHz6FpDX/uqljVG
OZrNBAnPLCGGqNKbE/kmrkLDFm0BULF9XJtF9phyj9qyHuGTGna1PilW4xpUD6oYSiKK3YmfUdIo
+xmLmqQ6vj1IhEt2yb5Lwe5hbgUE8TRIrzeqlmHJkRqEkUDDOCfTloDzACAlGFfcuGwK5V2/1e/n
/WJdktEHsfup1sj4kvfzGMW+XufQEjmHrX9YqqEMBgqKLpnXGGORo2bnz3Ify+szijmiRzTKG3/V
ceZ1SMt3kKQlI4xZLkhN3l35BzM1XdYTO2mD+ZuKFAY9Ueiye/FZzHgllN6jbqHDAqnLJTTWkvPW
VlidV1MLbr3ELy9lOCARFhWAMB/lEdiicI/v6axGc8eMPhRMJmRAJsaJplEmf45ut772ftDeKCpR
OjIWB6cj2ryxRd1Bqr5kUAJaImT9XjbhOpqURrZ4gkH8aAB6w3s1oLMhWy6mW5jz1Do53MW463Cw
rzevAM20BPPaODLdRQeGFWbLoiEqQZyJ1B56xOWdR8cb/Iyphhqdh1eNrCVFo1weo/BXogUVoEKI
b0FMr1bQlozFiK8a5lGnH9GhW2RIrFeGjMK2+d5bUdiEwF9DMBcm3FLQe1k+AyiNH2okZnsxXTUr
FmjCWBUSvMgqUk9Ai1N/lzgqx/j6xe9+4zk3k1l1qolhvy4aJskxzFZu8QpDPnS0d9HK1OdAqWRq
Vj6v804zaWN/tXcOiEt69WmikyNfEv8Be/vIl/0MQYW1BFnVgUtjS272/CC5BlWb8u/Jt35EXtAq
T7SNbabQOKx0jJ57oVEizHK9LuzsKhbMETk9uLHCUcbAeb3uWU6axgMVC5ezXmANzm1tBedEE0FL
MEmH2XhIzYZP7FVWIrGBnS61hSXnIxwCvq6W0WBdYcfuhMmIcTQ6EELtZAMfAw8n1tvpnXFjFf5a
i+mPsxm2CgdcrF6KqtAy2aFgVf/4zhF4quzCGxmEW6eIxuMCBPMBuTdFWdvG5D0fIDu5bWs+QKYR
jhz8F6Qg5tmEkzvsGbqkMT8wAwRUi9t547HEDTWFirQZr8/JUj9+4qWxc0kMDhcLwM4A1IDmknXs
j7nYf18AR29FVVD2IBAFZSn2dI8oocopQ0Xx6UYj29Y7qbgltVq0O1UZxXYJlDAj2CGyd9NVx+iA
Zpp8wEweSL3uR8F5AOW9w/R+0iufdNcE4ldJLACp2QaDovu+Wh557wSA0YYJfQO1v46rJN8XZj1p
Somo0PqtY5w7cR3IrDQwR4huB0wCOZNo3aYbRifn8HyK656BN1hY9n2sGfla5ZG8iP8LFGMjB+lX
dTOJMEi8VEYangr73jFEIYOuCCuA5EYGT4xTwTDIz+4e6oWuVHLK0wsa7sBS+IbF1Dyk1NveP+RZ
flrxrIMmAp03GgWfoG0VRg+lZux2jHNg5qmcerVtdRBFGTF8mgNa3HRounoZIWC0TWLVKpz2iHNa
kb+RN+i2ZdyJ8fNJVi+poxswLcsWxhTXig9TlFglAlrwViZJpYqJeT4uG8SmvUea4HFl1YOJoIFh
jdxd/4afpZj9hdrRg5stfjyyvxfBfi6zwz3x61Ef30EdAa6vHwZ19QbyIlfIlGDlvHfmKZW+ZcqC
UZc3H+RsZmfrdmEff/49W1YLPNNnX7D2FjhV4PPqZdR67eKWRvXpk2lRSfEZheI0aWNd7Wf4pdrR
FiYS/5e2qhM/b0k/iS4HpxjgjFlQbhEaM09j3foZ5ZfkjAo3ucv2PC/dGvntkYCRv4OH3lHU4tnV
3O65gEupvk7VhAtuX2Z8He8DlFMjEDzvdP26ZDvNOBfU6a5vWw2Mul2aprj6oefxjCHn3VQoljCO
YeX03V6xkjzLuelpdkPdtUQWl+jTzgFfQcxH5au/mKZjoXd+s87ec0rCa6fqCxkiPOHWR76c3UxS
Zeb21/KpOcg8ya2NZyVqb5LLtoVUZQIypm1QPQ284+y+EI3yEkbJqe2X5AJU0uxkSUdssfgfrbC5
rokW1Se0Y/jremzALVNBhHr9vrBr6oak+ymeLNVNWdJMYE41IflTjUWvF5vGeRYKUWs9y5PmR9Ri
9ri0jfjQi/qPWyvbFgOViy2Oig+2+NTmghJzeAWzXrVHoXBb1HpVlf+1ruL+tbVqGCtrd9qGMwN/
Pk6cyWW8e/j/qmYO5l94K9g0FHDt/XDsyGF8B1sWJh9276ALQg7DnHI8BK5jcy84u5DRVSKB/qiz
CTATzfg5c/7entgZrcdJykAhlZhFfEd+kNe67hHr6cVe9bgxIFW8PHaRo+4Dl8yN7VL6BVtVuqDo
rv563AhWvEAUOm9OZ6WYS6fOkjsd2IkIy/U6Y0kP1ih0lFTUsRjdqqG+qOcA9YSs0AAhqE/VNDJF
2AUzR1GkhzIprHCo7sMCs2B/z/O2K9ce2CpeP7Lm6i2O1HqPvN9gxF6AgjWah/Z9FlqCSaBUO4Kw
0PhLT23W4ajL1H3KQfhPjS/JtYlvTuzYvmjikqPyAWafrTsoxjCBIPIjRuwRnbv4Pgzl74r+UXcu
NwQ+ntqjP3udFtVAJ1ZitYo1cELgsy1pnyk9xlvPdcmUNqzC3jDwzQIWz3ruftZ9RoooX4I6emTI
JVrz3rtQ81PDvBRdWad+lyoYPHG5xngpN6S3itOwCyt/zYqKneu1J06brV98vs2GCnQFQQ3MV9lj
ywma1bx4kzEWECo9cwBKyEq2Ein1u+hKPEH3igYb5RFe+w1R5LWWtWYyG14X93W/Ypf8de18c/YD
FZHP0KvaJMCITQHn0aZuyKO/PJS0IZ3Ne8W+aWsCWRzBcaNLu0m4vl84xYciGaLTt7BAEIBnCkQO
Pcnt4w10Wfxr865dMFMWe3mQ0vfJQxSVXLCHwIZbJlDbZ/1b4eU7taBVXuWox33v0imqgs+0vY1S
UVYbB26divNbMCFaI8zP8+yB46Ghxl++Ntxp3zCNHd+OcgM3E9AYf1wi3ytoav3Hk2tuvPQ36OZq
nvE736AJvGngVehYALp2LtvX+EBkvqfDVb5wYdTuXqdB7iFBoYYAAPGHyPUbvyyXYCMtRhZhJZVC
Mc1QGargazAQTh80m3E0Rk07dwvB6QTdnc33eiYsMs5XI8/yJav18i6Nn31mbwvIjNkExJGjIYXX
jTwwulPFDvceQEEMBrzuq7xIZT9xJn2CopSeivBCCu1JNQgiZ5aUR1HgcDw0HHnzkZmUimJrmZOd
SA0yDC230lqXE/MVClEv2tmyMBP3BaaQXaah6QdL83ymUXjePq7aMxF8OTtW6lSuKsNfOSAveXWm
lAFX+Ly44DF3vHFuvLm8VuplC5NrMskzISoKQp/Qn5U8dkJDEnnzWlELGiJ3SVtzy22GCPO7grct
1p6cEzkFHJB+56F1SZLkLatV7OLN29TDdqVj3KBVJzOzPRpLPvgHf9rt03XY5slcjtaOA07seG/M
4Axi/4VpSrI/EMucoI9XseyKZ4+kRLkknYxFvd5B2L1KfMVqCLh3xs3+ZXmetWMAdBw1C/2iikfX
6cNFBbMfPcXBk8yHsgtJ7mHCSisZEssri2rhpBUxiMMa7UIgUV75ZVn09WiyjqkuiVVlxrN0r8np
gaYvwG90W+d6fxUWBK/oVlj0dK7w330HkvzfwdU/LQsnb9etjacgHFYkYUQJ7UMRdrvQdHAGF89B
3wt1L+/vBsRXKU1+ERRIxBO0aWojOMwRU3akJqGU1W0sbDBa0QJJ/m3HXg42ar7UVmhrJctPsvnl
oopDJj2U6C+9k09KuguOABMjoNXcrUOszNwRTukvJU8g7gZjxlxlm3ex7SdLjUw+0cD83fgmVHg/
ilVmh+5J/fZBAqi7QTu6wzZSIemMNJp8xatVhqatfWm31/nan2f4tDiTWqrg/5s4jwxdKDFBfCnE
MBYjCBhNK9HPjdQPSCci5lh/AGkx25fijHl5+7r8gUuyW1KMLGbSc+m4b0PTfImU8dt1FglwEKAJ
6v2pDqrr0QLhL2LTPlOzm9m5guuOeM3tnFvqK7XSzaYgGa7cQ7WMVcA9l1met5PTBJG16pV3eUMc
pSD7whhH1fsdeLOVTuuPPq8d4CpXRWWIurQVz7v/TqmrR2tMlBt07iF7nYkHqMAh/jWXGEzsoWUT
tGBldH7wxwPEEB6uwsAECbeJERRXuFIFrmN02/NUO7nRS/h7HhthXEaund3CJAt+nUZ8YP+zZHEN
yjjQNeG3z1Ypbb8aPrifxiSCXqkdBxL3IhCBSjqeL0UmmHJHMYlwhpJMSrDs7vxH8S6mnE6yU58T
6OC7qWj2fECOoJ/OOIrZarxDl+Rrt4s2Jc/1VlmIyBsCT4Ee0KAr+K3D2xhusl8ah7JBLMLVNOHS
lBvNaWhgvLGkvpI7Z8C7XjrH13dd+zBH+pwWMcE29SzwdDt1lRMCsn64E1XsftPgRdWrqLCCdGXc
PTu64heLwgFcBuoXXyWdFFsWdbJ5DPPy5i1l3fE0FdEieaF+XN8RXYYKLi7C1Lo7x6SM0sOWersL
mXjqbxufWF6YQx4Q1Xfw5TZEK3DBDK0RoVgCv/jcIXCVgFWPz8uAbJql8uOTgwkD52BUXRPK+LDu
7Igw8p+ysKyZY3ev/yaqC/4tpjNht0YorbjY71LDO0lgoShTQULhCGOY6Y1EQHI/okd7wQeMZJwL
JRgqapGazI1UVQv2ZvwNbogW2TSaAtEQBwt3S6q2RTSJsJYGbfXw2NYDRGXK0CjUqWO7/ThIFjVP
d5ggZLZ8uophhlvwcbAK2iEuaWxsyc8XkYbjTojcNU/VKbK1cqR5VuMKv3RFS3BRDZwHr2jzAM3j
aJ1NmPwF1pgcMWHdqBmc63O7DSESaiEEc+Ru4TpnXHO0rWAr6X1WLs1ddoJCb90CdDCSGoHhJk8k
AWawajTpA6sYv5AQ0EIk9aWd1W17NruplPZvOxDCJOdISYrAz/9Pol5MH61RKsi5MocyjMuF0QFN
Fwi8PpKS5kBXbvC/fzy31G3SXnOy26FabM/PiUx/9guE+bJCpmplxdk8RWXOvY1XWIrY3GZQ0zAq
7RWHyiGcUK4gY7blYD+VxBnOyP/qahRFaX0vycclX3MyHW0ZvEMKf8GKKeUdRpChUuhVmmTpACPK
7kpP0N2JMdV50raUy9wRwlRxugDwGzmbyHWqKRJwBR7yHjkGffRmWY7JRdqLdEoqJ8sMuuk2ifDF
RERhFj2Kf4RbA+UcKkoEWzAiTcHJdzIFIXnvTSvSsKL6eIDdEmSN2iw/DjWu8P45UltyzDODqa3G
j7Vvmh7kDwBIjD1fIN9BUJT9GBHaG3VB0H3BeNzYpFeL0Dgla5tgl8Wq/PrU/lQcQjZZKLBoI0hY
0RBhPysyeN73WyFvT7CQFs0rhAASY25wQhF7OXPvLkWkjSEzFY/U/YePconsYBDUloPvSBNF0aNd
575QfRpAVLavqxk88YPeIRlHXON/eT0sOh+3/AyZJ8kksJ8izeoFY5QLGA9ikhrqLagcmnbV7k2q
UQeGqqax2iNv6nXNh2qPaD62qv+O8AkdgbAfS2n3dcM5GWYGEKEu+551Y25GWMF3JLGhAQ9JuwOJ
zD3JHDo3Y6hmJCCAn2KzB3C2MhWnhrXqGLVpzOcH/hCyo1jBoLbyloZrYDvvlLx9MskRzNPgavEw
XfxkxaBcbX55fKEQ25rMTgv9tFBnJbcGefZQyTICdFOmQUO9KZ939ePJePbf1ad8pGb9sjRrMdg8
/VkBc77BXeVZd9UrafNSiBsSNwCbxw3ySSU6Rw0+vU42WRNXponaG29Terd14B+tCTEI4G6Coovv
qhE/jtHW9MPByX7UwzDXz0lQaOPqmzIDkqB3YtOQB9f/iMtEL/1vGUIj5mbXso1/o6fDfLrFzW+C
+hkZvDwekxd+Yjrsq6pvip3X5A3xgMKH5yCCfYxiL6j1tUf54/yQdw73T8aBckkamwnT1+gKI9Lk
Uxtf46KRnBZU9pCXXoPjq8jbHOuZPdEnUfpZ2aMZzpl0NFxZTi+Y+cHioKCCFmfaAwvhqu50M2z8
+1/qN3kxElIS1wL5NUoiHTGRAc1Pnk9q283mxe1WvV905Yh90RfLnZFA8ZO1hK8ZOO6VZDMdpkqR
wpGcNXI0VDHlXoFBOQ8ON9ZkAgBONbFJjjqewarKV4pfnlZjT5G4LZNtsTXy8PN37j3bQwI4TVn8
F9Lkicoxc0SZF47uRuwbzRwYKgth8bPRVnvLrn2qT//Zr4PoH5PUBkgh1MVxTuVkRf6OOsY99bNL
CNt29sQIGuExmH79W5b/vJ5OE7C0BZmKERlZTsfYYhLnhGDrh65NshtSHAwd5cnuAN0TGRlf+5Nd
P+NXS6qOsWo1W9K8l6AzAvUyiKag0tC4D3QWwCamyHXU5csplecfIvCX+BPdnCy7T2d/hAKrCnes
Z39vCfKdu18NXn+iMJwW0UedHk1gn0gT82LqUdiN5tmuNk6EGNq+dHx/viCmiBC51wdk1t+aVs+s
RpH5bog8MQZXINslLfFEfTKnhYNrXoDdq59w9P2c4apj/wkrVDLgXOvUQUUpHGEwpGI0NcvOn9n7
XZ63oP62xREscBhF06AQKLyY6BbNfrBJaxTexY/Wl3dWWHFJRiiktk8QhesTQQWgALm4uA4qXaY2
unM/OpezLLWoXFVIiKHYw1Hl+EAdRnTOnuWL4DbItlyGoxeQsr4JjuDdjVksjeRQFipdA6P700Nf
zMFSqwaZIqOoIxMJIDlj9tHuvGunMGYdDiNMS0VgRfLcjKjNskKo3CgRlmMM4wBAslIoI70MaUHz
r/iD13YUCZyzOaxq7xLe3KuBFieg+7dAX5XVmxcDqCIDjR+NCFDeS1aQI9mamhbDHQY4v4JIFYJr
uvjP04N+Vv1wdW/G1KPsD8UC9LZUikbVII/ONyd+/IJ9BbDv6NgE6skXkd9mCq0QHFQp1wThMT68
cbrh1Q9zD2J0+0HW8mtRkzugTnJ30P+Yo4B20aUlG16izsf1R4D1n04wIDhYqk5CL+RY2dDsEYf2
pTZgLJF9i+xI2BVPRAIkmjT5X+eIcRd8RpPHCzpGj4nGEKOOePxNmE4SySLc9nBVq6sFzOwwiWKb
SCuQWiPiQLjUXI/4aiRcpwXJ2gONKz2a53nhf5rG/a9o1ynOnQaQnNqgI8jITPukt7XV63tQ5XNL
uMfGmAtACvpDbn3V6K4rEsn+eeKyTiAiXOgthzvjL66GZ4aqH5Sv4FdWrFiPuFjBpAv3vbesblGg
+tD0AZgeTF3LJJd1yq6/c4dz8aKH8PbZD3ujl+z4RBYMkCcOqnc7JfWDPDeq9ZfKlklJC3/CUHyn
41nfOHKK9334MpgvXoA7Wo0TaBl0kB8LR8PWGTkKeIj0kt/YH6z1cy7JOO5iuyZkVDGnN1riZLVE
Oqwms2LigiY7j1L0BHHDUYcy+zq+z2XRNUq7s2C+AS9a0SAeI/U8kdMSIpxQpAQCj3womZCct81a
PrBULrVOOzYE5166iHAWUH5njk25D6z1Ots6SjRJp6SpnPjaUuD1j2uEy00jV7GVYeaXVUqbYoHM
K5kEnX3UQkvPU783Xt7hE/djhXFnV/okrL7iRFxijzDsw/j+59QhuwkbLwPHPYuLObnlLsQ31HoE
D4Pw/p4ohzljBX9Yt7HaSmnVIbX0zYf0DQVNw3nOIT/G3pmmu5ccEh9llZ/EwTUzBi7fqW6ZuF7K
tQ3rxxzpWdq97Q3Rh1fxE2QrMx7YjlW29JP/E+aN+HzGYN1N++o9UylhweNzUmm0Mzf5HMvBtxNz
ryWXrFJb2w7XKpM1tE+/T55/gSckkjo3tBqW+eI6eFj9QUu3cY9vi8y0kS3qj3JdFo16UUt5ooVr
m7y809yAN51aJzb3zkO1dDLd6WcmvQyh9cP/M97zB5rzi10qfuh692M9bXVuKBrvHMCKpnHUJYmW
yJuRyjV/siNears2MsoiisBgWQopvuB/IVUrt1G5IIQoXwe38n8qvOLGSwprC1sSpjH8ofNYtCYT
x9Kp0R9RwhXqgHwOslZVK19BzeBnzdbabG9YRaX1fHIVyH/Bk2Xq4rgEEBB/MzAM5hO7Xy1qsQ/9
baPqzajeSVFiMF3YLHzeUFL0drn6S/AzO+U7eK/QyDnyrmZUEa/WU3/Vvv09tV/OJu/aiHbPiuy1
CMDIc6mxmZAX8JMgjaFRKhjtkBjjjIw0XMhdXrwtA2mJdk2tZH2scnnOTYV2ulab6t+ysjmScF7t
d9DxK2QjXhVmKHXqE2SkjTGBCUkUBpDDWQ3ADf4qC2ezvRhKo7po8X4lex5fhRdCvhJiI383kn36
GhUIuO4TKF16UQXv21iY5CHwVC6ydkk4ZnPxlnTE8u+Y586qjODZhbq5QOSZyRTeeUWmOZ7gjAX7
yCq3YTQp8SeFvs4e48u6yI7iXL0ZSL9DR2uHtiZvVNsnpbNun7wB5SQZ3U9jZYkQHANQDMEN1dyp
HHAfQO7HudXapq068u6EDazIeZJRa1bSYHMb6mEiEWCBEEaQW4ty5djy0zHWLYrZ+rLia/T/BrZl
6+QjqjqYELHlr84tecmtGx5uYu+Tn4VT9RPvrpdC1VJ8ecRVQ1lzefYPb24v8V//YL1ImTHTxFbt
g6ozA7MsxfiNBzR54CM53RfRj1M7EqEL7TLh5WlLwjkZ8Ef9OHfydKJ35Q99gJpb3wb1hBcHny1d
lSzFSqlOiMrKat1ZLqOxY1k9zEzWLb9NkIUYhqQoQLkrAji2ztKbNnmpt/JUG0uESR2905WBB7Rt
EKRJ5b6MUGYQhWNC7dLTfBd15cbQOHj5Uy0tEfWyI0EIH8ZiYgM0x0ABjF+QUuMWcy937zO7uxrb
6QsAgXF1tu4TTiKwGZyrQfcuCNInh70Qpauu4evMiX1XNGBuckqk7sNaFbejexmzUWbdk06VC2Q5
Ar0TJaB5h8kzIF2hWlx3cK72K9lE7cu4g+0Aa6bvgWGLmQFESUvYrKH+aU98tZThlDdYRjREoesv
dtnfpVHMDm2o7CtAts2tiZQB/7w71312FgthLYe8cMYf0h0o2o5si75TQFbwIbRp+hgcC1GcnpUH
fkqhdsGK5zShCndppwdIijUwtrAopfxSCShoo/i6GPJZprXlbmRcpJVXwlU/U5Mo3hGS8Dl4oL9i
yUIDLlFD1SZRRSuaQT/OFmwDKLjo4wGKq0katcCShSX77M6+iL55/MFUc0/yV+joqniBbY++U54c
nquQA1Rby3KZsli8l1nymZ71nAF+KGaZnlAAJKeQ9aj/GjAJtGSw/GLjoNMJbBUX4m0hm2cmrIvy
s1+tscZIl9kNpCsp3gh8vvTLMkMhHM+eEpoR7fiFtk7RPoh4ivbI7+zThusKfvuCMwKLecJja6ss
ijWV4B+E2qO0PlPblJ0l2/m3YsaeH3enpfuCpAcGolLKsyID112XxPfugXfeqwDoUq9BLefqJZ5x
0K+Cd2knFx/dNFDZarXz3n51TeA5tFv9C99K8jScBjCARkxSsYLtDexDJ2xBe7sXz+SP6q/8P1od
2iu84EsR4jFqPuDuaG3mBZTW2mou6RmHFR2Odat89tnaIPUpvlEuCgDQYEaAHW6eP6mBkU0OEvF2
VH4YF+xLfCgLt1KjTkzEtxmormIZ5yR8MB+AP/LCfuxcE1/PqhYNj6VIsqVDNOnM0XQaHZ5Vx5JO
06J+aFVCL2DWqRLedpFtvXbX5VlXR03ZCZwL7KVvtIPFianN2lgcOWNvrzD+RloQOpcaljzsnzJZ
JivfHE99oXZi5HRvDpfYSGicvmo3nS2hzLq9VpoLLqCAEcCLud5dXNXNTd+2uSHPik2MwNwsWRAo
lvK0PSI11/aTy1V1x0c5erqsMmjnXpRepYpn1cV+MHNz1b2gfxrzkfN3A4C9pVmFTcteEMZhTPnx
Ju3NIDtsiCghi2BkwzmQkUEi2QlM2f58nb2Ej9T3Gvl1aNpdBLqanmCrk1Q9cJz+NyruXew3qhE4
5OfkdatROTwnIVgeH1v+n5eqi9LgUH6Az5DgIv5IKWzmOE9hbVmn/8P7YTgJOrbzCTHGAOjQOhHa
JkWitOAA/d1N8FKmfDCAY9alByEgO4X+t7oXSXExRJAxWFrcljtPQHi1+w6RHe2CwVkO3dvAt37D
ld/FK63vtzUIxcFo8mmPA4tqMTFhMm2vQzPlv0iYY53TDzzxO7msrBomuNy67DLr1+qweaUmRPEn
utmEsx/wTJwT7XCIdILCS2ueUH60x/pIFQmqpySxIBoACTylBJWe23e/d/eD4zF16b0g0EF2dQLU
46cA3Ryioirr3Za82aDoFk9qmziIaVrXZMnp0bgzQk5mWGxLU3rBJIpwK3CfqJo/nyr2Fz0d57Z0
pHzS0HDt8WS0Cd1iRg+o+DCTFpriEyIGEfyKDwc+xmOtNI1FuO8XoAliQSBXShP5k4sRIiajbJ09
gNbgh2MgWv7CJPRnI9ognay8MzhK+/XgITEokyuyzSty/Zgy4ZSmn9fvRTY/VK4I42ab0Cxvp4In
A7aEwRVuF6Spnaxu4g3FYos9ci0WtbzuU1+gmMvOnnGTzbqQVnnloRUj80wUp7lROW94M5brN1kj
d6wcu6YdJC2MXT7CVyKaQW8mOuQIPMKixQE9VjCAWTNPPiFgubOhO6ksG+1P0KPvNu+b7s3Lj4PH
jeX9JnP8Elpt6oibWiAXUm/sTjYfFKeN8HBsaC3+8qNg6DOan+uj3+P1Ln3ySlAu7nwQg6avh/DZ
SToASFXODdMAJZVxTVEYHVoNFBL0LT+lJ+X7jZvoLSbmj37NeiqRiZN6cr/trsZAYK/9OW5C/ZaS
Dcoi6lnDY1W5WObmhMkfDgU5a+XwlxWWvoRihzqeQGGMi07UTl34JPUOF1wueta1mhx0vhXVXVSS
tFNN8NXRVSv7Gp01/GZebOItRHT+1esy5MNBp45Z//rz0pFPzWUjmJEPXUGAzDfTLEduj9nprFgb
JGxmSwLh8kEp3N7fCHd41jnUzfihjpVVdpNAGWRv+stWJsXEHq9Q73zCu0KQpJKQLhtyrfRwBXZy
G1T+pSk7eFFWUSkWzXfmvBjBO1FD76LShfpOZ+/gNoAevICi2adaddaZhY9Ta5N1t8sxniycFyqz
uz+PveRq5qglAAwWyJ6MKyTpqAqImf2H6HkNdHvzdO2mdhDCejhB8Os53ur3mnsQi0AuZfYmwvkL
oP5xY1kAphltTblUDoI/YVarfnJVGP90CvXHIslavCXAwV3susG16aahEEWAzRU7FZphNyxJxaj4
/LyAruyI/N97rGNDedt6DyhpFUTJfN2myNxSJpT84fLZAZtI/GK6fnASzsByNVkX2ATi5sMMCrIy
S48u1EYqU9ePpJz+sRhR3j2YCBSS8IkzaG/SHKcrSwtzGSoRtYW/8074ti+iDZThDmqgF4tFA9bN
skZR04omfi1ur53kRJDpF7lPbPDs4mDQMx/88mRCIwHFLyrsvrqYKVHV9rfN4vki+BI1IIpQx/os
WE86tOPfMLLoU//oxEIfwe8thVYrM7EShmhZOh2Aqzgn0tWrdBjunxD+K0TSrG8CsjRjzoVX/uBe
dTCaNgIhdd4njKzwijwcVcpdBQTkhvdpsjIGqzV5PxOGGi1zcG3kD1DGdDB9KsXO8McOLPsxp480
0H1Vp3V3Lf0QdMAwhimLK0pHsCogO1epnbDpt8DjFM96Vbn74Z7KPedMkBsLWG9w+L9UoO0KfCV1
7flQdcNIXIpGpva52r4D6AgH/1Iechm9AftaU9N7NsbLNWgJiWveVlckWnj7RCJDsuFSwnfijvXw
8OmcSFFV1YMnPFpWMZIcHlmvCEb+8RIpVUErdSMcEdQL3UDsAoYZn9COc6Sw6O9kWH62PjGNWG3U
Blam0Q8A2LxaLdnTwDOgI49TJAmJNCdzWOWoVNWb3g92PnDKRGrO+W3NMP02TnHCZegiIDPQsXZq
xB/8kB6i5JB+YkPfJK7S7rMq9pd0V3ruQ13ZQW/E5gGhCMnEzGpfjqdPj3J0a+Ci5zBhgDuU9cGj
2O+srC8yNAV8dvnxAEAhyQC7uVBxkMxfEa4caf6S1ghMroWglxhizSxBKx2jeJVQb6yh7/A3C58X
CrO93sKXVxstuB9W1Af3+pa7G8/0yTQDmGfxZkZWypqu3B8fgmoM8wBS2Fan3HQHUOqjDYvoVQOr
AIFV1MxuESB+Le4lSbt1UMf5Mf0JjXaGeMG9KPMr5PwwZXXnY//eo0Xh40JlM+EQTVQFFQAvnQMO
uBCU9GzO8r3n1enUpeOLUCOYfcsNix0xjapxFf9IzaxQVPK07/2CC5o3vSRQbKMtRq61Jo7OOIj6
T6rYrZzWFZTdMnQyzyphJhUJzHutRK62E4Ze0w5Xc/4RoNctmOdkCwR2+K7Z9opXkgZ1SlmCyeel
v9HIxuW0ohNJ17NKJeFnBJBos74E1dvXYdOSjFCG+cKxgbOEZDZ7tSLCMN+1h+15fVJQF2m6ZFLw
MEogGONzIb8x+MnnuLPY/+SyCGcYtmo4xs3YbdjHHkn4OipYbICm74MoenPAVNs61ENGGyWcTEss
rQmDw2gIK/gcSdtiXVNrYQNjiTo0vi1Pp9odP2svJl2cmxY4fGJ6fUKETYWcxxTv8mIjw+S3R6P+
mLz8wcoGoSyhSygiSuE+myNXNhjSb0ecm0WOfDw02lRr/4tgLlKyTByeilyaxTljRkBI61PxGKHD
ceiK15hrrhNSVsfLq3+/vr4vFTVS40hF/EteFTDGIat01KiShjqkL9u6nLiZKac3pvVyAnrRpqK3
H2ABznCka7KOeVQUxgOUTfovxlZ3XXlUN2DgVJvjNZCK0x9xIoVWaxD7YOr6wuEdrHjAbdvY3igF
pa5NsLNKWVfH4Xc6hwWxop87HvlK87HvtoYZ9mUhEYX5ucM01Bat3HUT9pl+0cYbcoLYDFblHBM0
YKYqwyi2A/lbxx8+ESWqEKq5/pYNxWCwD07dUKeb1A5qTKetjSEGBbC3GUAgvE2t62vG0bFMUlO7
x0X6x8Sso45N2DxL5bgnQ9pDhkio1pA5RMpqNheJnRRpfDUOEAHQDY0o5L8b9RkKekRHLe2G4FrC
7BEvq5WZglZCQMdwHVKviRQSEJUfjilgw28SjIqknAxQp5qVjxeIfCoO+u7Km+BLlCoszS66wkVP
I/s01ND3oTdqB89O24frWtCfgh7B9ThBiZ7YBX4haxjmlRmWNGXl3UV2HiabLNMisJ9zjDlqLpV5
5Wy2INi/JvsywjLJOwIGt7yZDUx4oRFMVaiJ3YK3Z91AoOkx9fNUWcjSKNzN4prBFZp9nN0j+Hku
EOnPIrCQ93wv1OgmkEzkdjq4Yk/JO5aIDsqRSGvtZCScC6qVY+F9BhWp7gh6jvLdwInvpL83s9mx
QubXXss80bnwbI/T3hqKrb1BHYXKgjOwelsnxsdw16FA5ZNBapDeNsRgoC1y7KkfRtjItuaowgxY
FDbyaZMyPecsuXrCHNj2noQ4Q2UfdxFoygIEuKsBRBs7Vur9r/a7q2/7F36ZX9TDkuzkqxUVqaUV
rCtSfVtdQNFcudf1FacN4yBP9SOcnIwSJJcOfLjO1SSwpsKQdB9tQftpBQveQnTU3tavKdWk2fkO
69Xj/OqJOhlMmvsmzAoK9yOfApKYhZpaepmAaHRWM4HEmKscgNNrci/xp65no4FSwOP+wgVhZur9
eAj1KRjgbYnKCGYoPlaq8GzjV0+hO19pM8tTkpAYwSe3Dj36EKNztRH1YH3/Y5lPpDvwZRVrsVFl
j98W1YimGHJDQM5+S8tU00dxMd+YuniXQw+4jKx/QD3nhoqa+SNBwAbLy8KCgs+zRQFfXzJ7nH4y
0hMVtp2ebUqpcEoY4y/rBBbiUUod8ABd0Zri3HsLDBOJlCIuBDsOtmwCRRZMpCiwXGL0iwu4Bc01
65zUFn3mn1K0FbqUKmMgEwCzcUm/Z3i5ZpbsOc3Wgm3ure9FMQDXdYaNDDkGqGwdmxv5+szyD5Ph
QXgT1lXvL1jBTkzrWmsLCn5cNswAg2OH2nVpsOIQHBQbalwgiWLs4pLAsnv1QCA7sg/jyi7/wFWi
hilCH73zMNPXxCFrIcFOvmk07TOwwTAGFOk753dTHXEljAECHcin7LLCi0nKFLck2Bz94dY/4wSK
2KEqTPhoJVSpE2aCOXV4VfJI4yvKFkomzaebhUnPuUkFOFGlHRSvHJfzrYlBtamh8UpfyayJSb+k
WPinrpM+Ay1PiZ3zwgkUirgkO+CUs8wwWfInsh75ue5zdRzusLOw1NyQbXUrZo8pA+ZsVEI415Ko
ahCH8Iw7KwYtdZlOvkc/A852jGGDsT3PJkEh3MUAZzxaWDD4N0PFGID9sUPqGO9oUTxqWVee7Mx+
pYSWDYB+o2mOZgcTYM2cKOhwxIhNLZIDbSnom1Bk2fYkpNzny9T+0Ci09RO8nVGvIOjSUkpgpBep
ionk92IuOhHVF67XkBil+NYf25nszBhsmtF4LkG7dD35ZzHWuWKl4BGH9WP+9dUlNDR9P47cIx5P
TdwZbbk2GsOuc8LJHpgODn6PQOioVMeZ9xHraFpgy/dy4Bnbhsls0vhqRhEtDPuG0ZtlwKbvV1Cq
xjdxtHqfybcno83zdUyUajves9uh3pxMIK5IsO8XHL5OFwOibOicCBLoJOIW/JuSm5ZcEBetE0oy
JNHLI5n15n+2aCTFcVMtF/Q12NH2jjz72jqn4FVQ2dlRxIcifmaqgQyh/fsd6AVb/Gx8TM51p88j
qbRi7ad3aptbgBxJZd49gprNtnRvzYCMIMUauUksckr6k4nx/kFfaD5EH3s0mUgdzkoQWXZKMWEl
aR33SxNHgwb4cS5Ok/7Ceu+IsrEGJioSH643D1v1Hbl6vuQYRt+WDFwHDxpSQdz1atRZyDndBagG
aTBQhJeNVJqBK140BGSPOCI5XraUkEHI54owbJ+60ndHbYtXiMDNvivXAGwSf9Pe/jbjEgBZLfSw
1wlehyCpR4XfDDvrbGdB403PqRCQTB1fpPg2xCqJOHDnRHv0vvWi8aVV0SKJyZQ7C+BFGYGTHgzs
07j7yjEkCRQtPeiCNpr4kBFO5QKUJ3k3xmIndt6rouWPhN3bY6zmaSa2t4AgNIT8rCTjErq0yOXC
JatIqmJJYlhTpH0E5HKnryIwNyR0PH9a9t8GlfRGSwLHdA7gvm8DjFVE0vOZvsUWIsLcu6df8PbW
HHinWHqUXXGPWqAPxgVObJxAxIZlSq1wrqYtFRmvB6zET+6vjUHJtciAWWL32GkwWJc/785U3ci7
mgih05z/gbZT9wMJLYFlNw4L1WGnz/ibAQ0iqZXscZkPVHv6BgXbUsreyczoi7HaQjgVocmtz2os
CKgwrsvVV3LKqp3RgmFvbn2BtrY56GM3o/xjZg2uYRa5ufDcEOEQEvNARc4JJCpN0IeNRV1wP6+i
ZHj13awYRIgeLDahfjp9slFwhWYH5gm/9UtYhPgYfSggQOMMmCF/i69I4eIIWCXarhjFGt/eKiYZ
SbozFYdSjRBeb0RC5iTJ1D8aiyAzwLhYYyIO8GWQQoX6oL6RKWvC6ZgmUnL1/VblsQ9njCLD8S7O
Ueo8N/f2DvfG9xcmZf3rDCaEHAYIhNVafjKJJHCfpSVj0RrpTvsFunXQaRoDn3CTdsKgRRiWk4Bg
D2PAXpP2cVTP5Imrlr7boH7asXQqnqLcV5m6v/pIbu6MYrZXJrT5BGYgj0lvR89U5Q9O2jcKftW4
a0Sf6mW0GqglEIrPR1TSWTdCygClqBk8zyIZ96GIZyr0lC1BALlhypZjsO3Q7QjB/YmrvThxAdHB
X3Dz2CiGMZcn7da7073VsU5eOp/r89CfAcgZPPr+8JFxQe8rQUD5kgjhYLBT/qBgETXSdZR6gSZd
2LeZgdxHszkmMN2/bha6l3+0EDiDe1mY1UKRjr3X9+LHVIhXvCYrcDEziAxVUAtXpEHbPvRV+5SG
jhUfHrP2WrzPkQLLBuXrbkakeneog+U8BmVAL1Ql40lZYuDQzLcyZcOD96ZdleWTHVQpcLxTl6qz
Mf6eTk+Rhyiaeoflx6Af/kNS4hft55M7JOHEHxJmtBdYk/lcwi5YxgOLN5dUfwLCp7qevEbyG+eU
1K5ohVsTqLd8xTcQXrHonPvBctCRU7WSiyQ9xfOqVTSY8C2eKMIYSR/7jquHU4xU2Xb6VYW/NVeM
rlUurofkEvczErU0oU7iWJRWqDrWQaMil+IQYyu4uAUD0rC2kuHfXaEfFxL6RLOn0/Vf4tNJuDSG
Ny4i/6s4gIUn3TZENl3GSUm0Lj+Mo9+mAvIdj6b7O+8O0S6VvaI5zg0P3CDQT8AmCzTCatr+OiV9
i9bdYZIjsVxo0JurbWqr3RH9z3bL+kz8KYv/e/W2YIZIxBeKj1mq2zYHhjQVFw0QamBIw5JnhaDd
zTI219xRD+qkRKMFLEsuph6RUp2Y3+8QwnIMyL3rhRCEMuvFxEpqXu/GDKHI+S1SShfYaDi3KvVV
BuUOyKZT0pE1hVO7bxf9UB1bD67Vxxn2Pc5LsyKBkjz37tJKIi5YsezNx5IlBz1sS3noAh2/K3OV
Qtx/qeSlX7MRYJaBpG02+iUaEbVbgBVLz35lWMXt/TTyJKBKXnCfCP5AgwVXgnIOxFT9VJVMAn8y
AjdiWD0RDC/C5HRo3Ao1ZtjTHQarzzN2rylf+Y/uQ0M54QkP7LMCU76QnJIQouKuyX3Uz+C6GedA
zJtSe0DAwYJTiRAy5bg4aZl4oPxczjvh7YRjQDfySHO6Li4IE4F1xye9UuVQkZNr6JtWiSsv/Qf7
1zSZUgSeUKCihpmxXekXoGl2eRNig2g6wrMn4rqU0J6ogECwNwvh5nEInjmTuOKDSc4bEAIEhJ8G
4uOtpcorrwn+UwNaX7hM2HwB6biywEW3sybDuYmUxaTyPOWFioFD8bZtnu6CdGzIrAGGHJyGYnxx
g4OJ9AbqYcepe96j4uCyKLrTcqiZTlHgy9paVAutSUpiEdIG98sz3EjDEll5Rlx8hgt4/2tw52x8
hQvQpLGqILpWXS+0yQnDUJAYV4m5OfKZwzXX2n6c9qv96pUOw41Bleo/SYhibaNH+Q2SB0kPBPZ/
/3RutOwDoAphh4AmocpNqlnQUYpp2pKuKAG3RAQWzU93Cw9XWD7RMFVUDIIS7omivKabrCN1S43R
S4ot0lCsvwTB4IxwQW19PVOet4koBsHUlTKPGbjvHrbV6DOjRUDXlg8L5eNJwxLhLKAp1G80KODe
v54LMWmKRnsi6InUud5NIFgRCR/4bpy6xqwlWxtN1Xl7kGToLGmT5Tl4BRoazNUDftig0Blv6s4+
yUEhMLnjz04jd7S4nKS8K1IzeiXdz0iSObVi9D1pu0w/m8mefc2lD6NsQoxA5B/oVBXfXGx1q1HJ
xjZ4Yam67T4rXnIrbtWx+Zr6ShCt1LG8FxJHHDL4eU55i7GTyVZgSOAizIgbfkcV+bkOoM4OrXAa
xcHKVsWgS7RnQKPj/HEJLigrc1Szv8XbY+XjySsoTsvPsrh1wgw1mlrmR2rRycFsLFcMdN99b9oR
s8rX/lzKYNw2bPXcp/XVZRYr2YYoid1xk6chunW9cSu5KvLUwjyES3N2HKmKEd6giepmaMpHN4Sa
nb3acwpDg3/FiI9wNf/qx6Eg4ge+Q0zydAd50dmHoDSZYAzSwfaX4yofNPAtKfO0b/9WO+7rVso1
EURqXaalIj6RKcuoqjdwQdFYq6G1V+8fZIWqRpbjg0MpHpoO3rUttx9Xak2PQxT4/7JaxBE79J4l
S/v7s1b+lktO7PIW0Bfp9nsH115mdehzT0VgFGQQcsrUex15jVyaV1OH7YXSLgsLMBVcw6QU8sA0
NSh3oTmvZ/JoMrBEzgwGk0yODJuWs++I19vnQH35mdegs/mOdE/9zMi5+ET0ej9zuS8yS4hutb7V
qw4uE5XnsosI01XqcMXqom3qrDB/9ro5dN68Fz9TdWsNBW3n/G5ZrmUE9/g24ZVAZDtD8ECNAPzr
EUYmGLxfELmLMLfVlzyepdcBXorjrR1TXiwEXANL+kYcA5/5lHCccoqZvntPbufgFCfnHbN5XD83
otarRUhmf2zkRuI1VY+Bp9uhV1VlGmOCIoMLDWVEyUOrQrZSMuBSRHTVtwEwfNdDafo7k8TuaK8H
qyG6jjtJw2Dd3C92/8Q7eQ05LF6Bd5wZBAfS5P2mejsXw+33AKsTZZbG+ucWwPkCUESvLvr9TBli
PRxma9kAV0EwsLEjnvghAau5OpWcTyE67M+XVJZOqfrhDbN7kFZzIwcCdqt9mSUMRoj1mkltz8ck
FsAPzVpvqKEd+Oc1un0C4K0ESu8ZLMs1w1G0L2hwi82dtonXaTSlbIcxQnRMYVhw6C3sN6zuqHk0
JLyE9ZP8OUATpgd2F1m7J9tVy07qmQvMYqS3LPHgLhi9pJ/UVonQIFUABa+Jt/c6S1NR9VhSflDn
6K2URxr2B3XehkCDPo/zXNQQD2t994N7H6JU9JFB/GdLf1R8j9i9mdms0HmKMVmq60zOXFKtMUAq
K4Ea5AzDt17Sw5XQ63xQaNW84INsvl42D7TPw3Al/709sPfV7PAJn5wKup3mOhH9Dd+tDFk2ksFP
gRlctqw04X3jM4fOqPxDUpp+kP5jVQ3YYZmSP0ZW187gKxih4i83JlHEbqFqj/ip5lvGB0KiMx6n
J/JVtyld7AFF+ISoyInXKllmj4Z4X5iYW/NJU2kExF47Q0c0kXequz3wMlQ6+AQMB9kmzC1NHgOi
K1pWvHy8G+vFL6lf2LS3+uoDTiVP3AyKtvhjnnMDSChydgMJ1DRIbATT1WnwnlBJu0TBERbvuxOq
vl1l+dfLTYx2xLusG1dE4XdTik8z/YZV5F1wlhGkSxp89bIdac/0Z9E4scAOE+9vCF3LufmiUNbc
16W5cwRlyh/wmSq7fLKSrUSeAGbYgGwuOWfoPn3whH4c3lmDwoCvSQeyC9lSl2rvHE8RsjAFcZGV
q2hl65MsSUIM3CG4XkyLv08TC73gMGautrea3fdSZAJOBMkm4/yOZg7pFa8d+bGq71cR1D0WsMyy
GWP/8yJeoqA45IBk3ini9q/IxLb09QW9tU2JtIToCmwr9TttVmhf419m/P+OjCdbwq3h28xXHDBk
EJWF21NVFNHp7R5lI1SATMm4HgNw5D9E1L9LvPCRCY0JM+X0+B3MddND1h2+YmX90PsTA20Zw4A/
Yt17kMZ0iife2WHHmD6XhxJ31bTLMgf0pxktcyzN+i/jnFbLNw3equniABEftYYhg9lAbUFM9hcx
McCIBKkK1ct3YXj88mxeB3rGPPQ2s2oFMjamaqou4YzbyksU792VepPmNzXPJ0+VHLZayezhAP1r
bqNaxSqoy1Lr6djmTJocLDAgm0OHMR06Q4O9hj0sWFqpSFsB1JhkVPYP/jpKz4/gTtU1/nkSdOOu
BVsLDN4Qnqi6zkbrLHfAizH1r2URq1citrUqts5sL+mjNpM4jaxFsYGbBNYGKLiGwtGVNz5eFG8e
u4shdIE4Q3AqCGGuza2TP/fpAMFGEF4SBcG3yQmK+JSaI5GD5+PSb9rEn0dYplAGNtJZtegzRM9G
TiO+D/862mzRnCIK1US67dH3MqChkobn8wfjUHc6p1yE1o58U45MkuSowNp9NbpMwDAf4C6C8SLU
aCwsufRtnjNu3JtbKO6Ei1wPik8cZwhsCdjFa/fV/5Ui17szUlatzjRKA6tNakhXhUGTgXj+z7ml
kEZ3XhCcwcjZ8a5RA/p87bUFWgPkENtcEAhATBKlQhAwB24cPIvpw/IN2uEc5KMDMhuTCblMPiRt
0g083TTfNEPswiHOiG7x/LXogoL+Ghiy9NKDrO4HXZ+MhLSoewfxlU5ovY/e7I73Vmej8E4/jtPX
TvQte4y3kNlAfd7yfyjpmXa2Q+zvJ8jJAT73pP66zy3BTuevgKV/wgDDMxAEFgLkindD4EXAYr0v
8ZMfYWLa6V7gqMs2JTXlltP40dgmLIsAXRJcQjEAahn26ok9rfAwDvNLUMWmndoPgSIJu5Jt/zgQ
lACVNqqmmTFHI0zVTm4LriyYPMQj/NZfy8wl5NEnpVN2sPi15GPVAWGyv/ybOgitiEt/bnCmkWTM
srWMbpELXGBt8yMlFzUw9Y7Ub9tPaceuQoZ+UG9pX6pJ6SX46bEPcmRQQrXE2r+scvUBkVTeTi+q
YJGlSOxyteiR6CztRSJzli43s1/x91AsncF/8nKo2IrYe9wX2IFS6m1jIMWwy6LTr02teiSFx0TT
i4DHNzHJBaNRUvUp9Vt115vnvv1Ke6SHZ/d+7HbsKgyQEPQYi+bApkapNyOdc+x+yeROQm1vGVCQ
nc3JY0h+tKPpjG3R7bXADSCcP7nKaegY0LFZOLJlYDTZdyWEsY6hdLdqNWpJ73U0PUvTd5zd6XC0
KmFq6fKGyGCwIDgSHvKrMc4PPTJMIQugOQJbXs6fbg2zdT4ZRh/BFTtwTrfrozNriQyhMvmhGgG2
CycsL0nY5pNqVv2+xEmWPEa69+iuYgteEcGnSvr2P1sVxpIo55Jvu+m1w8iNPaVnuvXFpQ26cNrj
ceqadyFz6h1/gBTNT9dKfTAsgyWZiiR0cOgvAza8evmm02kdjbhlCREx8WUJGtYtDa3dYTOV0yoH
Av/8LvHKzsrY5bfgS3oGnviPbkYly2x08wtCv2CI5iyGm8npU105S4N6SMkFwpbxCc+pZVlwgDtn
L9esq+HAx9vSuPUjAlET69fPmyQJQ0GPkItDj+ETTkFb7db7ImdsgKSjj1J6yxLT/4vLWXfbD8L4
J7HcPyK34Z6DGebskoVV9KzDLSD0hOWN10/1gL1Zdp/DvHAL/ZZQ9LRbWweot0Wh7Y0dmZPPA2yC
6ypNI7Dl5bZGGZJIV+cpQrKvpXrAetsk6fGtwr7ExkdsKHUgIc01hrvZGfcE/KH31SVrNeX0GWm+
JFMKoRVdSHI48KlR2DTNCPnSDia3ztcW6ce+aysh1FMA/Akt5cfZS8d39FLEO916RzbR4FLo6MBp
T5d6YQMsEIYz3ntqH5+X/iScI9Qd9yQy2lvPsptxaXEV7GDoKNx9bM9RoRqVqv+/CBMltbZhVlXT
Lza81Yw5k9R+ZWju5w7fW+E7QDn0H4gGWsZo0jfzSQMqv0QQhsR5OKCobEPu5OVxHC0/ibQafG17
J3q0XSV70b3OUKl157isKzQkLbL+iikcMGUzCTa2P+ZV6Wo4Blh8UJ/GdhYcmjhJCU3cxf72QbHz
d8KSzBP6Q/TXYAB7vw4xdbpkP1npZqHhcxts7MxH1FtWpEikJmKIFk5KajPvvgdgO0Y83YZL4+i/
egfn5Ncy9aU1rzrzeiQJ7OYWJHiJPMvO/tytKIfscKdXu6Mfq33OAF3SVDyw49u7nXjhwkV1khhs
3+Lamn2Y6AXC5iYlcjgP5Aecd2pXfSu4tCQ5mROlwGUGOjjMosKNBUonhOemO2Q7QO/sRJlVTjOS
pZdeGAYB7yZwfgfbVhbTmLuTcqYn8hXMOqb+lpMbvAUXbavN1tPU+bYjpso9Wh8qf1lGY4vjixUu
sCxaElUC0WMRVGft9pG9FPWnSxPv/yj6UXGnx6p/AJRuNgYZNBpF1Tl06Q5VWP2e6IeuS4tPrxAf
bI9/am30lI86bng38xZ/ChLNBzf6csLaDbk+2l5bMquXiiZjqA32LxI7ftIFkehpbK+Xz2IXY5ks
P3N4W+8Xy9Fht2QqP0TcVEdP9PjVjNVMAm5Iz81GYRx9vBg/jAgB1G4Y/3s6cy2CDY17vtGXuWoC
eW8ZrwRRInRcjukEOpAX+utvb4UgwmdH3FlxZG83hBtyQp3h1THtiBPMCUQPXMl4AdchYKYZ40Dk
AKkEDmu0Ju2JAjA6BGTj7Hh4/ChEdZxCbXEpMrUMM0prnPGK8JaWs/B997LeN5ByqpAz3OB5RHrG
pSeGKo5VHwKXurmpNlufEfBuVp9KXkwJIMOOBFYGG15LYbZDGV8rXbk9it8w2OfvwXslVp9wUxyU
CAOcljPllyswtMKeRyxugUuax/LAlXA4f6NGJmzJu6QSxd9GNX1yBscVbDFVUuF87S3yVFTwVI13
CrAR0xt20BzwI2H7VxwjB5i9hWHdOUNvL2Ucs09N0WSJ4/YmosruCl5wJgg+CKVSK+ijbSxzVJQ9
+0Z/OG2h88Qc711eQ3RPhwkscY7GQBP/MGGEXHGeK6dByuvc33Ji9uk20It8RsXqXIsS4xM2RaSh
MxAXYyLdoQjKumN0vYBPO4hsM9loN1vjR/GH0pNO6+cA9Agcigzm4X0+5M6KhAzgtlqxZsZcCLne
3r5v7W9CDWceeRK24f7tKjIahaq9KIcENlHpIArf9mXeI1YpF4v6CoPSISLYJN8RTcUKGIw4lAQX
nn5u0ZpUsTgxgwwz8qoSvRG6EtJPCLnkcss8r/OWQdM+c96090wRq0CUN4FR7cp68ZpS2hi73+tu
o1KbyycekSlZmI6AOgHj731L+bx8vnAdBDJT2CKP+n6WXjg+7wAukpvxj9BY5zqcRLkwOaBSOCON
c9Se9oLzxwKC1Bqm8apTh3IOQUv7A+DaayOyNxdAhEf/PoVskxPpcuRbwYZH0Hp9WRH95TUgUQDL
SAVR+qtefWzA062iT+MM31psC4ous0DKu/8r1gWdUfloNt+wvtIVlMf/7H7aD7z4ZZM6IVAtZ7C4
Tj8POEzCE+reKXok8YkFKx3f02HwxiTEtWFTdpZXjME4c15QrjKWkFRxSBCPWbMP+u/eA3X6/UMB
Fb+N/FH4Bvq1VtzcURxJcRTbQVpcFrzsBooyemDO70N6OY6jmxECj+IF96CYmbTxuIQJA8hlzizv
OP+TvFdbVJ7ZSDXidkKsMPJ8BvVuRpZg4fe1/YwBLes9goKeHU4DgTWcunJgwhq2yyJ0AXlNtWlB
HC4Hw8EfIHKMkyAJTqf/iAXKvEoCkC+X6p9Gcw4WF7YWBWyuIYS6C0D+TDA4Hb/oy4oxE3xpua49
Xzoc19cPlk8wpQRy4GK1oED2nirVCTAU4s9Z0kYgxzXQh26VHk+7qQaog+fJVsWfnNwM6xLlltvT
9aULVpSqnFMTsA4dpzPRXZtTrNK7mPIRFj+0liYopZlQVrkb2gMgQB95JoJIM3FywvpC1a6gKm+a
O9jmKkfEUFikUayp83+tDlnnpfW8zFfsYj0fCQ+QhGtj9Tq9g00hItKHSnQ+bg01Y+SIjPjItnMI
mHMHGE3M63lP3Mqcn6604eMqWqB3OreGI1dxg/Qy0W0V8N5lMOhWZLsc7VaDnIzHC7odycPA3RQC
MgZFYKpzJ5J5gLxTdtJOFNYhoQz1YecPjKK0XnZu3QyL+nOx1RdS3CdeyHtCXUhwyUr6F6u12q9j
t4Ouf9eTxod1GhuvIqBwZE/slkKNaV59N1uN94qr5ousdasoKgxxraimDp3oSJPiYtcWXknh25Sh
uw11ne5CwzjfSWBJ9eDDzrp+BZYLIVPdu9vUJT91P9CBKzw9V/qqsEQTOk89ExYhmX517GoZJfia
JrQsIy14mmceEHU4+pIbL6/u6a4RvUQr8MuHDV0Mcd+5WrtNGUPb0w24/okhmQFh9MzL47ITaQJI
0CFbe8rBjfZ1x0GDrI+lPu39Wf37Jd3VF3tJ6PKuYxjfGlFJalu1OBS+dj/WibtLdofv07bzNQpw
0yQiFSEXg5hnm/dpPBkV8TLJr7LwTrrkcVajkQKvGTsGdFSZ/mfAHRzdRf8268KIFdQhJYZ43Zus
uIpA2AxFw9zq31zk34hdt7An7sx291GmLnhJqou4Xxk3E4XBf31s2NphHiqfI25QEtCrGA+MLuha
HPWOGWzNiMdpAnvMmSSmqLB0GrpbO6On9t9jwOOqDMO1DSE6obZkQMQpUSGwPjhH1rVvR11SJXon
IlbbqdVPYAoB59fjCrbz2U5jWq6uaY9ptEDnkQNHiwnuWSiXFlhfyhHrmMVKVHu/sN1LClrxRqFT
cHb3k2okvWdOlA3VXWDz83NAkmpNFd523Od0TWT3JfhEgdSvpHspETR2infib0PFq2BBNOktqsNE
bjO8Mp9NNc/f3Xp1yXIjZEbLsuYU4wi5utE9vDWPF9LT0uiYic/fFOqr+HLxo92jO+bpqjUlxgub
0DMrlIU/JMDbU1ckmc/How8euaTHv7U9XRzB+g5MqK361sRJOrNN/ouPk65UmD8hJDaBz5uFMHje
lqo8Bhc6c95BRs0N/UrPtLGk7t7juDc5FeL/Xt6ldXqCiXq1ImRdOgcAOJAdbU9FCGDk9CS9z32U
lQ98t6kdRL9yanf6YOZgbOajEWcEFgH9d2ppdMWksS0PrvuEcp0Cl5mrZyvunTlJaMyY75DXXF3g
PLSJigQU4MdFx0XVDrZKVhfGtmw/u2AR9bjUNOfG0aLh8eHt6UW5o+LRQDi0YaNYFC83Kq3VG1fO
9nAhSr+LkSL3RpbDev4wLg1DjTOUIKyudB5RsUcnWQryA+N1nbD5x3iWA93kEcAb8xdc22AMNOco
aTk1aT5nOlEVzs/wJdn4znPTlEy4/9VX2FF9Y0AI++OlVkymr/SYlfxMFKXxQT712TuoWB5xVU56
rcEiOZj8R7/iE0KwEuBWMUHAuT3n4hEEJmK0jzUIQS7zt2V/483W5twX/SX7oDRrSpeXmvO3dvHt
g2yXmIGlPkJRX1PreIoz5BQCXGqZ2rt61f1K/TUF4/RMDsowhFMJuXny0It7rpLFxz3j7u5S4rvr
stkih2FCB5MJTJ1dDL4bO52+CqQCGHIVScfv11Due4Y5qBYBv5JAdPM4PKXUfLzKpKDVMIdelep/
++PbGPTbrokGHora777vnTgZ4z1bbwsIAVL9D+ly/JOX3dDdWhZ09LzavzpAhK4KR0gF0R1Y9uZS
2/AsEY78OF3+ItG/5IbJP2YafqcuZd84qTL+XIrzCjumG/mfkoFgrUPUkjM0aYOAG30/r16RNoUU
l+DCBR1K8TMWEU8/FeqT8J3QI2uLiMW3d0ie6zoc+Vjb72DFO/71a0UYhZLnV/VcpjAaTQVMGZM2
fYgLjnNI9MHjVPzIYVr/KtLM0F5wm2Nnh5HirOtaJfoIBRg1pNkM/1sno2QtI7OrY+s8MRzV3uKn
og8Ec5Rzvyadh0LUOyoHmEj10qSxGphJshEyLhDIgU1I/C5u8vwslDhYtRVCjseRdM/C9D7bHkMI
sILpTRl13mNAYqCaXG7sTn/BIPwDOaAXEePmbaswzfbN6tb8FFjbZLxs0HZNe+JAHkrT1vX6ox9q
1XbfrESfXbhCOOC81Wi5wHH3XlkH2QfGE1Em8fQX04emYN10XhSbb5UugzL28tt8RqBeIhn4HuWg
HNwYlzqqln1G/8mpGTZNkEk+YQr3WurNAz6Bb318ga3e0JhgyQvmGkthQwRYBvEIqftJ8xEvXBkL
vIXdLxbt7+3sLkEGTovsbFk29pHPiJuGSHNGMXsVHzcN/vJg2Q1YBJGnC39hR4yGF0M9hN9foZ2X
bSN1PF8ydTL9jWiwC4yGbxkSW2oWK7I6AgQW6OQBxrCOohCKgNCiNsTmCziS92By0MzNePkks7qK
vDiA1HjL9TrZXBFtC26F1jGJgoVSebVPUY3HNJI43QRUFjFz3WVsNqFberHdkuKPGZERnMhyVLtJ
QJFQuGarDoRO66yMHrES94UFbJsiSsxQ6KiVl7cZGtfl0E+hSbbwX2nzomRLV1gqk0vYuXDkgROg
CQSIVsSniLr59O8Cz/CXBgiq3Utx6sHnBiZmyl+Zsoe/UtVOsaTEpbQAArGwyFqnhOBFYK5wDWYw
v87MEKDpvUZ7wMOdU+WgQAjFSf+0SKvAiiQH/YB1wsutjcNIrvSj7bIdRdWaiGut+XCCx2UY3tXf
actiC164lXSEt/93sSumu2B8QDEqyP2O6IsMRIXuSbqQePoi6Qg/ZleX0lulPu2DIc7cfe8UWGJO
hmD/hf8zwcxnFjqZB5q7BfblTRSKVCtkUhlBbi8TkyKpHJkHc3SwwOKYnqmZxgMVYw4/mL2gnOLo
ieLRL6kC7wtvvh9jNjb+qf9XyAlmDstCZpaewMNDQh7HE7hKXciiuICAN9+CtBjm5DH4Xg39TUbt
O/vGVT114jlJQFA2hK9VjZpk1tEpW3ULs5YUlRIOOsKDCUxmLAzt2xgHJsyxIuwo1i7/qW460eQm
5CpX9WfXyutIYMAweH5kmPvzyivyxEsU/aQO3DBjuNucc2KeZ/Q6uX9u5zOvaUwKZel+728oXpDu
QdApSScHjaDu3L6/JkxKB7Bal34bUean4l+vk5yG3wX/WNYWvg924f5WVxx+SHKX/IAE8Alpoky4
di9wdw4XRG6P26UeZSEqLyvNwv5F4xOI4xxEzWjJelIO+f71b01aPJj+Dh7oRG2l6CJ5UZTt69le
IUyfCPoP6s1Buq1r/kQhEbxYuJf6wxsDNZOUL+uj2F4I8gAyWcPAV24w4WIwFRmXGcnVRX5oQ6HO
228sgAJwBcuO541Cf35GDCdauFDFzqXNQ70uByVnZPzYlkGgLbmKvGN6x295poi2ImoK7doh+49q
3ztkTttF1rCXa3Xmk7dYJ1PyDYm8zL7qnnjc5npABT/bVhTXOn9IuY17Yl3Ygg0N2C8qHVplRKY+
LfPwtqaXIEeGu3x1Qgmx1tsNcu3rs5+IRBgpbMVoZJJFB+g/kEii5MkwR8/R1ppV38+TYgWaTFB6
ZD5frt3LvLjAqLiGUeFxyiitxZVdYZmLqZh6ASzUmy0S01q/Kd8573JXWxxDapa5Y1ze13SbramZ
Bh2QqA9DUz7Gs4s1sXsiDaXTb8Rc6e/RwTYrrPR9EEsGZMdiTdme79fwtRSPwQUlhg69VNIickQE
nnQ/2+4tBr8Nfcg9UUF5MYqQNbgeevTTOJ5bsm/FqStWKGTYYciI5EhmAOLjnM2PZonqrwLiTIea
y1vLneR8zEpyLDDYO8NWuEr90+J0jE1ASW2XEnSAlj9a5xqpXgpfIM4uAebRkjLlob3NAV4HyjPk
+cluoS4U0U0ZPikvrS4iozZYnAcv9sRVf55hkMfeUxlRaWYa2VxgCdM17KCxhjZNB/cQ7bUVrvBF
4SD6ZlogJQo8d6b0bf6/GGxZw6GGkIgfEcLSfjW5whDHU141E+JZHKbmpebpWcxtwZ/YuAIle8Ci
wXDNotD01ecK6Exs2qd+46VgxHR2XRoHVdiJ3FcX6FnCbcSSUGQKgzH6rVHNDvyg2J/IM5F0KIxm
bRYkVJaY0GYj+kasbGWarImL1tvNQcNrsz1JR00AKtM9QL0cbKO29THzq2AD9v5uDS9apy0CXlWL
v1fZC0TiL2/ZiZyuBwCMQPGKSUPu38a5Q391rsMgnrHqMzJMM/FGGvhPIrLlEFXJ+5OKHnYIaOd3
mKWcAIOroo2mvVjL4h07ZAaA5xhfcyBIipXubv76tLgOsI3btdr6eCsyqinaOlFLaawcm+HC+U8s
W0Flp+OhDRMMFB29plj1De00FBDDpkUlcBYWQZi4r0n+5aTL94aTzcSrlysZbvvR7/ukW8bFh44u
LJarEoW1gWqEB3pRsWqf9bu49Pi6D/JF4nBEEdX4asp3D+hxTST3mHPsd51AOmaPXO4H4YjXSYrL
AtWlczPcPjBsKoX2p80q0qp5JXfITtMS+bZmEheF9+d1pjRK0IExkXiDrU3vVBVKIv3c35JZloiF
jIv8LYP5T2HhI4Coz9A5zxhBwQsdzSVM8MaJcoo6/AXyq3b0W6Thcf6NgHtbUgwpNEFMFMgDqhGI
77fYOnjUTqAe3l3J5gh863+zdB6FbQ5L9QtZDH7467BWjS8Bz3OBLKHqysZudOJ6jPxj8mHNBVnS
BNdg3TQmDOstF8FrNROhqaAe1NcO2/cz3se5JWPf/Z8fd7/WC7AR84d6pffWaqIkfhosPv1Ag+7g
OfXMTgG28lV7LO5rnqUiPg4D6LKoeNeDyMKaDcfSDD3tHBSgAxwAzWrTqj/dwcDqVQJN6dUa7htu
BTYA7fyoy73aAwmIotXgmc8OlXWq7clYZk1R5jQTs0m3wXA3fuaoMHZLSo7yDQ0Ai3OFqkFRbDv/
Cu3RgMyX4LMNB+Uz6axhL9YtSndgFQh4RAV8s4TI7PLOb9qqNfX1YTu8eO6Bhqx7EJnVIcGnEMbJ
nAiU+A0AFLTMditk79m2yHauOZHOjhcW0kQlV/xPOR9LoyQ9Qbck4aXCzOUejv+uJSF6NkxH0d33
15G/YeRUZ9Fzp5H6R+0RPETqvsyNdwLqXeRaSAATGJ1CYPCNc5b6ANaGWUfOC8I7Lx2ThaRX0WvG
33h2MnBr174pkIRdvBCJKt7qzWU9SHRELwrn6Urux8v/9dxVMDOB3M5v9gfUeXEP/Jk0Tr+x42Jc
OIqGNi300tZNwBsAuMeSkY04mvU0ku6cNZd1wkSBYhezJNRpIKdJmPeK9J7qRCTFRKY402Do/rAO
W00hvFcOva70wn27BiY1yK2pDViA/IJ7n/EriYvzHJFgw/waRNM/J3MwnJqofABBx3t6w2loroh8
fjuqgVFXUG+0Lrrde3wtGoQZitz2cT3WLuC+YYOd8vog8eRNE9ogA9MsAvpCkPwpHmAffbu0UZ6A
b61V3zWnhrW/OdCGQdwYsJ2btGZiNbbYgeQtQQtssY/QZ2Y7jQ/uDgzbI+rh/5fqlmtNWjzMzFs5
6G61bNEr78wE90XIwRIqzelOUY5RgdKT2lmQzdzpfJfswyepj18WYaux9KLOhKBvtwHzE22+Ml+8
L+kdilAAahCf7W028lYojQDWwmLRFlVydceeMdDygleQ906X89/dHy9C1qE9mPhLSsKBGd9LFYDr
XkmeiJ7WQLmEeGxaV+VgMn0YELj8sAEUqlF7mX7mVzX6WRKO6R53FVhpxh5Rj6BTtzAVMCQxkMmQ
j+ntzaYl2gSlVuv3ZrYm0c0L+V9fAVDo05DGBzuVTHmMzboo2g5fLFW+95zy/rRVS+xpsGghMbgk
ETOeuoz2dtH4Go5SKVqLUdmIOvUQgCgzZWH46PON20JdkS/cadek7LvoXWHSKGmDFojZvqyKH7D4
R08R3UJvXdD5TBZWy4T7LmaVxcWJsailZSVWIirhqyrE+b3TfbuJM/3IdRoKm5j2T8Op+SVw2nRX
N6fUFzOnej3027KiKIMs0OnrwBvtEBFny1cnGpeGA4s7vd4cPwDttUwKgRnaz7Ux+GIn9fspi05B
9Ezi/Mr/6nY9nV3OciPuYadm0fUPuHBa53OwnwFiY5BpPIOrm0hqk6eZJ/7Jtwm81kshw3W8woMG
bz/FE2FE1SSlHg1n1YSZVWMD49CWSsMYeB0jy2QnXdjNf/3abZkjihzvg2GxPdrLJDc6ypamu1ju
dj3bdZak4t0Bsav0OpMoZg+c/InuEtx2egObSyxMe+PgziKYz090KuRUCB1MjhlUlCwtqh67PONN
BHQn7so+69EJZv4Ts1+kL+mCRH7lpYrWCXlNLfYq+HWDgq2kRd+G3OorlzMO4wuEO7FJ/MC0WWtR
k7ewIno0BQmoM5lo9Tk6W9IyJZU0/HCoLBbYAUQ8MVZl4IXeJE/KODvuZ6aO03VPmCCDSar2wUPf
D+xNjSCkEABdyxjBd8SOKP7JjFZtc4WOpBES12SKwm9Fi1gZJ4kmpbNYR/19S+v8pRDefacN2rOW
/SUSU/be/HgTTgCmGoXs8BZKQIyYL/f0gleqV6BaNAMQoLOASF9z5J5S354O5kByZxPnv3T5vRn8
gcRWZV+n9zlfaIpykI1phdnHJ9weg5WVHYVVbLfAXakSIQ46mskWUhc1c1jzJaIb2Wt8FLjoqvP7
Op/QFGVeNWBs97lIf9hHTS9CFdTp/Exxrqo6UgvBOV0eW/6ob/wZZHS/sVGMETlE9PqapkSoCSbJ
QH4i7IW7FWaRLEHiLGh7rbLNpOzwBCaqGQ0yfWqqueNQfJ2KGxZo304/A9KVSlPOcYmgZNancelr
x+EKXsrqXv8n1ZHNWlcoqXg7MaDM2JrJ9Z9putWSyImKNb0gUDB+etavTIBlPGMcHDwX2S+riYys
n+rGo0rN0/Q2s91VrSgDBOSFd98nO1bUx4VmVQKf+i1YId1vIRk3K7Gr6IdnDSU6cecnX3BIo6oY
1rP8DSKFHuRtLUPP5GANXGaVrI3BYVhFFcqT2f65u4OQfi8E9+fsBQL7NveJgHPqqJtjrxlw9Hx3
1PwFn+K+Up5Y9z9YPVnXvg5xhCe5pT80JcXTNJxZUBBexgBvUougAtzXr5KB5XbKwRCb3vGpw/fA
1ko5SIu+z9D11qVOtsaostxuq3PDd4qOXoXPXpq81FBjTxnViBohTAxowbtUvz76u6x+OkL3iz1+
zAgIwfb6y5U8oXu/+H66TqIsJUwFDOsYj0vJqYFXl/1elgX/Oq8N7r+1hmhSfbDeZ+3Zi05ehFgs
9nI5WCnIEcItx+zr9fIG3ke0sfY+Gz8LWituHkQvKvr1wKh+d3T3xcnqvnHKYJSwnl74b26AuXEO
exWS6njHDCewOtdBJkehg5yctSS1vsdT574TiTZzFs5pM/NShMAPRBuS0GoizYzSvAmo0j5gzvgs
riioivHDbIFbdSUadWeDp5YkT0L0nWwqEAo2dNz3p5e3OhdE9zmr+fx+rBmrvx22rapHL5ake0CV
pABLHSdbSmMB+DoMKiHSKTjqBrj588tkUm7mZrekdrH57Ee/o1X8W/n7qlRaTQhBHS/SUM3Cqhrr
d2KO0fkGixgEz756hF+VoMCRvy4DIxJ3o0bQhvnYW9YNW9ExwvyxNfKtqCeDwTaNEutajT47KtUD
GhCtanKEPEgJZ/Liv8hlWzueoWn4JLxSvn/BvGAVONUvYfEAAW6VVLROjudZb6dq4MPqOmWRpJYT
YNppnCZSKlm9jY5NaJutg6YV8iM3FW1uCypNclQbywCqHP1GqSqLX4giBbCtUrMjPgK8I5wUI+Ox
yT5oYBudxwegHwpA/R6iE/xMM1eI08mSqNUygO3Ux6lPEUIo52ekUW9goF6jSNsKlESb8iAN8Cul
B+6X0pfVepzbS8d9Dm8PgzBBHomLMDqfi3+X16VNRO96GJLM/BRTUmZiMgIfl6YTSXEukVvNSliJ
xytiH+6wV+cjF8+3aiRF5SaP1xeP1+Wgnb04mteYny9B+Y2BVMUwOg+5+kuxHDgPlHVhq9YvUsGl
JVi4I9dYzjjfEAGtwURUsmPraXAV/3QJrWDT1Eh78E7OJU8aWEAbqU3x97DBA5eFZzEN+JP5pcd8
pYWW3HT2ulZANnX7zb5UuQ33GLoJmKtL0yIeAlWWSVk8OT8d5W4FjUhJp3c5OiLvRrm1gY/OYX6d
AVi4uw7byy/QG7SJBYjvhf7ZN1y5UEDs0M56f3w9c3hwT/7ce0hu68SFnB73ZIPrahsaMoaR0WJg
2+/J+ryILoONXAbXtRvSQduxpn5nRIboz4Rqj9lpMfC7PG0b+4yiDtYvI729Z7/F46a1AQFgZ9zR
ZpiA2sIwLGPRhf7fSOrcuUl0aqgXOLJw9GBPfaO8M7CRHTdnygrUNqTA6u0wZkVT29E+26nQmgWn
dPmvA2ZV3rsJ4vkK7TqNisqJNnS+yxYNAFKmQ3bihMXDTCQjRHhPhi14P+jJCS1JGtLAPfkP6wJc
dJ+1zTsPsV1PtNIRmERuk1MVcDI50dYf+n3zf3dHPUI2nxCQ2xUmO2e4ugtjEegdfCVd08Ky8gUV
74WrHbRQP7o9mxoyAe8oY5Sv/V6VxWgCmvefKkO94vozN5IKlqUranGh1kG92fx3aowZWcJQWXO2
2velLls+FAjdgKl3vQacvWSD0AaQVkPDCybIcYeAap/sAvFawunACnz208bloe9CfuVTQLA92Rsx
k2qHLxQGSq7jtejAUkU6JEcqT2GF4jmh99QxzzeyvGzjJZrsEcSvwuibvyfEioaqs0q3BU3pheAV
m78rRz3wYqUz0pZXbSenwQtTKspfhIPn06W8YiNi7SRRnuM0cwpzjmq8mmLl6jabjEpw+U4yqtQY
TMQumHR5AEt35BnS1lGAI+RcXNbwDVCSjoczo6nJw49qfMIY5uLYTTjQVMNO0e5TqTitPnGhkVx6
4r19LXkHa9j9KdpvhbD0JrQIkD0688zJ8y9ihpdr0JIzKFJGJrhhwsO0YARr4bGDQYqOArTOmN7r
uvReKmtBN294xI/p4JkBDlZNMvV83KEPGve6fQ/W/EfOz10Xy3clhxbOS7cEnzUzh1iS07eZG7M/
KqKHoeK9TKmpTBjzsWaGOurIF5OGI1LSx99Ubm05qZxZt3GriTeV+QcVerB0+81VOlZXGxlIWXmM
/62SJJP15jvqwjpZFoXRyVD5wa2SdJUbA+8XszUsSfKCO5GR0jlOqiiWWpXVjUjiJrknicdhc6WL
DZuossF9PKOKjAUt4QuW86B4Wc1Qun1Pi1nn4vt/XpOKCx7gqA/LhSXRjT0i6T5+hgu0dFb8E7Z6
yguyJkJDWlndZrJqRLzaTj5hDjbLmdFDHFFamBH6FwFmwjSuGC8WY9hVATxlwKaH2A1D6h0lzl6g
7ogg61n28ZqVMd4Z/Vn2hu3G+3y18VgagmFLK94YcIg001API+TifZDDKPVZppfsg+lYfRYN+bEO
D3PDoJaebn917Xbs8wYLx1CGRhUw/pv2S32ioeiw9axEgDmb/UuDUhwBUWZzUdSQV/ySY+Re616w
nPIqgzx9ruaWhoMX68/JOW0Zu1+sPxszrGhTqfDDkZAPYkovJQIYOmPA7IrbQ0ZpooUTIlfHBGOI
8OVrVrQXhNuyV5rL6hULAqoNLK4YTzXZ/QROPc3JEdqeCgLoArgBQC3UYOhWbOFxMBG+OC0L2213
fAYJvINCW3b++HjIn94avZ0tnXZ1UQvzMfvVkuL1cebjom3dhl4yUsvDpvx9p2uYufnGAuQJOpTy
lXCfWjmsoetOOLmwk7sHZLbH8fa5mT5aoX+0O9ck+Gl3EVBuTvwmlcgMIbKc8L/lmThgxmzc7raj
4FAsgqFOaf12RZFxKo3zm5j1n7q+p1PweP243zHsGLJt/0b5ub/n726gbyOEumqe4z/iUiMxIS1Z
rub5HQuB9usv96Ey3HaX5uU0B/PFkKwLCR/JaetCQr994BK4n5/80imGrZ+Ihh0Gs6+iHsBXYdm4
iO2NF7rWH0mmOHf+513nEBvpePR7ugO/mgHHZAt4ePdZOtz0Lh3E1eYIAxYW7gNTZGUXutPkx90s
Ft8uSbyFwhRHRuzV5dHTMhokkB3prRGsG91UYHw22KYLgln6P2/VAGdGYbnt1fpQ9pyB/5tSE2kK
1uCZYhkCf+rDlEnFWNABzpw9nEmSFSUcFuvYa55cdlPhA/zyMHB83uXQCzjV7yQ/1mzJGiHogJKm
aKHkrmDQc7kJeyTSn2hedz/f227VmipLlgp8a/8aIgTYNwvUUZWuOqn/Mu0IUtopYwo86dLAUyR/
S+2RsivPfo552xEOrq3RX8LznYas21DR3sZ4/GNnjxFreAndR4J/7AvDkdWF03xLt2mS8CblMFMU
24B0uFGF15mIMK5bqHmTPMFwtssKTi8+5p/HwiMVEIbUwP0BlXvsVrZHRhW0btWsGlH+SrU+UMX4
prOSXUwQPIIJyubj4Kw8uyjYUDEcWn3OC+yLfkcBi5l087qgQkO7qtjlItUqnoI/lxpLpr5bb+bA
Y92rNbVqh5CF4o1WqzOryrQx6LokX3Ka9o4O5IUfzMJ/7wfZ6HdfydddthNh5o8ku1bcmKApb3ki
xFJdiJ30UAwyJg3WBgh3Jpy9ksXWQWuVpmC9WY7MHbVPFjEON7Y5+GS1WH6eJ7QdDtLjuVn8V6k5
VJFqp0FUn8UKbR7046QwXrnBAVBWMdZduJt/7P2lnBcXp9782kNNQ8jIb9KB/Ays8u2B3moajq1G
8mK1g+z1vV10hF7I5RVljitHyERwtMtwp9Wy7UzC0mRSIbSEUK5E5xCRsq0Jo/RkOQl9HLRoMXL9
35cDgRXfSUI6THuFRSpRDo1HGKt2+R8jP85zCk34wcvsSXC02X9ht9yBKAUANW5dgK4E8gJ2TX6G
XzLwuSy7lqfeIS79wt9qy5Om7bGUoPOvJmn8ju5axIzhNPYh9cI7rzUSxVc254SyoZaTO1v/y6O7
LVoVzRiyiAtZnDcarQpRjeZHaJqdYZo5eLys7bJgSyO7sR36b7cPqNh4hLSXaEaLpb/dKEkPnomY
rshuR7Q10fc0IUWqDfno/vtYZC64ItygmJ5RpOdfFePKmbh9X8g+x06R6zhXUZS8K6o2RxEZroy7
ldZEulumPUpUtTWPSSCmVHNugqhvcrBkFjx0s7deccrlKP6pm6LQuv5ltao1xNIyNQlTZ+D8fyPN
kOeMHEy96/Kd41GFVYosogmxGIEdb5dpUPQluKTbhMeBU8LTcV+dUYtxEpK61t9uhThPSC0dQOEX
d2j7R+MxK2krFocTK78O6X52KBvv3VqfUoEzh406LXkd2NprcSy+LdDOgVQ64w3XmTgCdqWMZAJa
Q9ThKopgV3LFDhOZDJoNmf44YHDb6AWxQwISzy3rBnWA8+YCeDaiC8puuJpcNfp5GiplV+6pBn/K
c+zcihFuCaTsexzSYl0j34LyMjrpo9dE2W3S69wNoPdjw/AQ/4t5VxaoclxgsGO5hWysbmrpk/Jh
OhIdFUe2oTQ4SlpmZvB8Vlr632Fz3HFy2cspQtWR90vrQ76z1muoPoifDgZTUtlOI9mb0s/22idP
tsdhZBtdCEuNYehTuyWuBs/nclpLXXmQDMPO61XH/YRIQlw8NEDcYW9UuGlOkdUilYMpWZPEtsAr
jJcFVoJEvlJiOuv1+o8Yj4b4otjkaB2/aD7K7hAnUdq3gvkQkjQZVqdDO+MD5Dxrz1u0uqKEhPP7
g4K5iv57N6JG78XWTH6Nu60vC9J1n8Blu25N2mivfwaxNAh9TG3ps4k8QH3skkLLs5JoNNmuRmoo
HpihNOi2ZYmOFqD5Dyi2h67lwJbWce4njMWtSZhAJseGtRbaAqjBexfY+QHc8EOmCHS1coUpp1E6
lkokxuEi9WKWJa7KBmCsKGbSDWvgL6V9PGDFbx1YhRgxZwskSNcGyFU+FvmfMxwWC6cpYTj2r6ef
/zX5FMnXLPkF22hxpU76i6ptOC0EpMpipkCkfqYwrnxbruQT8bIOtsTKECC8UDGhnqoB9oOCvLlx
gv7WKJkJjZ5CMxVvoToseXo2BUSnjIp3U2H4sEND277Mh1xiW/nTXxZ+iwyrR1wDA5xZEgAMqR62
zKk7JSR0UBvEZFQBploZ23FACnJlDQVDn76dy8SPZgZpoV5Lshst8JsOQDFW93e3rb6NugCQ+rqx
ZkMOU7Qb+OosctHqhi0eu1+JD0236XKOV13UTADUUgrvTyyTQVl38E4J/846jsdx9Og7Dd3KJsbj
orp0eti0vN9wkWUHg9jORluaTCzXh4V5/Sh6SJIr/bw5EAwnoHmSr3Y8FOyNQmINvdVGiXtlhC5d
R+ltqRezMGP6Mv0tNefCLwmtl+dR8YuQ5NJFM56AjlUaWyEKLFAYI9xCVaS1WFxQPDPkvXTW3kn/
BaJAtBiNLgkAVxazMoO85geckD/TJl+WVJYkEgPgzLX0j2C0/pzjQRm3c4boY+pGeCLfcbcTpUKa
xMhxStPdnycKLVHC/82k4OgMgWTGX4KGvEK7kaPBqfiGI6wX4ksMTdcXSNajQDZgc4+YVrTCeQEP
YLIyxjcv1AdqEpFs+0xxUQgwb3+93Rsg7jdS77Z3RBTJ+NoKuYavt4SOM1OgPEYkQ2/2dmOeKqod
QarMMcS80yye3MHccFb3wFzMvF8eCe9TcabT/D1+GjN4emX7x7CjZsJ3ha5AtIoCyhR5MxcG4ElQ
x/fIv1xrDnmVmKkJN1fYZpMRxpzKXZTLe1khfb8KWSRrOSjNInpVshcnM1Pnrl9SDhdibggihDSV
1/SJD80ASr4IjCRr83rq2UGBWO7nTUd9jImwPSYJWowmssmm3cfZlXtkdCD+C6OQPZPKpVqe8kxd
x5+PA3lv8+Yfzk0v65UKMs6zh9QoS3cd10C+I3oF1hiZLOx3cRnsKD+nho4rjIGRisdknIJsp4Z2
7HDia57QwW/rIlIk7rzBlgGVjYsKkPzgvb8D7BzUw2+OSIxXqHz+ge2eCAarcbiNsulegMEMHAjo
SyHcgspM6o0j0KZ7phMYtT5uHqK/XtTQ2DH20N0Hr2YylvqXTsJmOp5PgGO10y6xB1CoW36sywKb
xL6RslHLWN+p1BOZMSQcdYbGQlBc/B25/vJWX3DWsQXzW94xYcTsf14awP5rb4ODElS4TiRWIimS
NT0L+xz2HwZkQwcMUUOKgCM0t3NGrVe+S2xKv/OvgG72H4qqvo/NnTrp8Q+6VU2ATBZk0ufl5V47
IfYWaBNw36156rEljYh1lQENOjuOTSU/QgkFu0A7NGa4Y4jHKUJFASrl0qnZvYSooQjEWOx/HUWe
zawBDR2gQbhj4kVI0277kzM3KFnIz+XBtuV/G5n7GsLPGc4BEx8UjCKoV3Pp1W1ltkMjTLEHD/m9
/2wg+bnwm4U+XSWPBK8yaHu/ekjrzFBERspa6zP140PvGD/nMsEd1d3V7TO1twv8OUOvRjKDGErH
YS7fjHCUvh9haOA/CnDidrfSH4I3MX9FINsbHx/sC6UmrsQlDSslB/xsME4OAs3QpEoKM5XVZLW/
w+fvN8t8XucvRkLDJoP+zsncTU5O/IvvnrgjaO54j0Vr0K/mdUOEnIQYu2sFFEKiLjwo0MtFdVET
mw+tE90zWJIZNm71g5FxJXuBL704/cwLX9/1dGBMl9TTWiSO6op/9hjwuSE6PogKbz3g0/Uj62Wk
Eur76D8t4s3CS/JNq3yNMRNZuI1WRZhunNho3bXWGnr1iO6QrYFppttzCjERgEqbFtagAEdfrIkK
rcP+4o+xd+FcswcqsTDW3l/53qYdyDJjLd38PkhIiQVbFwO2TCTzy5Ww6DlkR/BMY8VC2+9O3+P1
rooqGh4dHlKxKMM+6EoXsJlFHnietq8owjb3gmalOxfixLVkdJNW20mzWPlvZK0jAuS6NHvGliOK
ZB6lLSYwGFdzjDAErvvYyvXEJDYkPQUmkXa0B1GnrdR3Diz0W0VpnV6ATzAS5TIFtIOYQjO2onXM
thhIh1K2ZAVmqL/iNd+XlP4B8kvm4/tbHJhLkZetH81/IgCN8A3NGx+hkAOXb6dbnhOidtxZ9ja9
GE537R7mwIkkYQ7093R7KIcY2cNciS7pUhe3S/2n3ZPSM19bpZwzgtEkg4lokBa/+TivIAiI6Oym
Q+aKHZk+p4cG1u8nq8GzCbsHZ8g2VCH+lmnCC8PLSTnosaUVy9pyqZkf/PHXCkBtFdRsZQaRUjm4
9wj9R5VKsCuJDxLp5gwV312K90VbpcLXm4GkdLXwrEEG6A6YNGFGF7JyHL3HRyvddOjBQ2CElp4R
hnBClRpgzAdqxFVjDumFDpQCh7fTd3RlDRazUV7Z5hJgLA0HdIvg95+wlNvJniNd9H4xFrvaWC4Y
geCIaS9i4aT0I5Bj7YO9PK06A72sY1sRtcx0e812o8f8MeQmN74x2ijyVshDHLxp414bskBnMjSY
ooQw5aJVH0jxhtmlyrQJ1ADdN0rQVIjQWZIAy0cZyCGNiercV/W2eX76ftaeG/t8HwcCdDkbjFzr
dt9hYU+fGWJrnd3+/Owfdey2AfoyjRVNZfrorjX96wrBAZPellFNRaAkCJ68e6oAb2YF3cXY4vPM
GjRiauzwv65M9e0rl5cw940weBCPnmKctLXDQYaH4qZAzFsAGyZlLkWISvbCAv6/kRWDWcL6jRdJ
L206D/CC71pqTFf2nwj/5huHModCzXJDWPmb6HsHsMVRNeTVAHRpON381iT981Hwq+gdIWLjbgHZ
0Gc35AL/r6BK9mXLyzbJsJiE17xmb87saCErlecXCoCQufSC0fVoFL72YDMIF6O/FhhjLcRd1SZ4
bvNQHJWVKHFqNLB4eLCdPn5ZbyZxMpqO39fR/lacuIBg/l/eC9kWbfGiIQSWPS093jGK11llQ41k
vfAbLX1fyOD3871qqlKA5nvc7RpAdr2PyQR6VThuf4PeKcv77UQaM7wJpoqLqrlkgn2/dCpOvljQ
RHpgbdk3DwmUtSKb+1HXbj0nE+iRniqfufo7hMQ8HYcJ8POG9rKLbeYqXlGt3aijcj+Gvlpraq+4
zyA7cfe5gMswuSs+SW5U3PRUYDoE3q3KC3ms+mb3UrPrc5iaQrXtjALEP6r1OVWcHtOOLTJv7YIx
YDQF13M4l4oYVTKVbldlTF+hD2lVO6523n8z2AQGVMtaMjrmQaB/IlTGlk9BplU7wxNG+laRRTtz
Z4H948nSWeeqUUrW+9+4tHY2Jev5/IGp2HG3F80ROUZWyy7pdb52rEoGkbGjX/WpCLiyU06AK5+e
eMlw6llIf9VQlLwABNj6v8ctGusmrSAuFxwVGXW9LU7scvxW4iuiDzVD47OkxA5Ac3Tb0voV3J1l
5c/G8GpRkUFz7zQZx2hxU32aSmNSD47FFQpy7aZVEBa9zlwXVQ9Gr22ACxx4Zg86rwlM5OT7H+83
C4AvPyuHSI+hJ/x2DGoQruvywdc+DWfJ1ASWcCm1BhH+qzn7EfmPbIdIK6H4FgTH5HUMPxcu+kjM
vKkxY6zWvk1xkdgLeBpTMGyQXWv5JSKghxYydEBPTK2sX0z2b52uorKKZqXaOTz7eT53DEk6UuwY
ar83+AXaR3aAuGtQtWYk4BVPAo7S9m7xTpVjM6UaUc7QUuqyGmE9dcHe4FvC9cUwn5dC621LI5gq
aQXk9VG2xr0myugIuLUbkSxcxlDHIEyuFR3ZWsBzCe3Rg70Nt1Aoo6IhKtaIvXHxqCRvaxC30STS
IL2HdcA903Ot+Y/7y/b53y39MWkK4RuVkdBtXvPsPbq0t6DD8E4HP+6oqeMqk0BjXelxesPe6DOQ
cANrCnUz+8x1zE99TB91Vfa19MZSeUNGZx/L0DX3uSKxDPbovPiDYBFlyuDnzpirLgfYx+O/U8VY
+lUScF5kCWOBoGaOcaMn0bB7i7T4mvKNEhVA1BKVa/Mx7VGn/+4M6+5/LbmyUHwE56CynsDnTaQU
Zk55GCJtBx9nPdKg5rPTFOAojNL86EzD88NuZ++b/IGiLuZUV8shTxeVBmgN65ywY0nNvqgT9/9+
xXFv/XUehbuWbs10H5GHzNrBpuV9Nhg9RvXaQ3u6ngxMRW2Eq+zflKwtZkVpAKEmOFgY21WPlFGE
Xa7v2dt2AMDFPT2S++ymZtJlQx5sMrSJ6+zCJBw5Z1x7o5PAVtnRUjPiGMrLy+gk1oO2ov6lF0OL
1wwIprSrKH2MnZkNEkUY2tl8Nd7oWGkWtDvvtfO1cYpotGkYCgJyIe4Reu4OOqzQNfCk7XsEJrn4
cZM5GMut9yyrdQLjO3mtih+HhS6AsCnkhWMRLjGutYVhp/NhkfyPjgY2XHPZVdg3+nCRL12CXCS/
h0DxTQx6f5zPa10X9GHqi6mZawpDdCv3C81LX9dtJQRMqyOmrInY8TcQQeGvd0XtFS1MzIC4mT6v
px2kP/wLTTiCr3UM3VckitBQa0ll20vqZsFibqRjwacxWtRVxv5MmmHRNCXTSDngKUB3j90HKylG
QYPikA1HdFthX9vxfasJnjrsdghOL8W14HQDbtk/SssPXTMrk+LtBdg+MSTv9E3X/oKRZY3rboDt
wVEcVgdA4frEk0K+GufxKo2iOSt1u73mqHGbU1ADeXkMvEYo34VMvsFbfoklZ2lIlAssg6I5QLB0
2EuPB0z3CO76arN71BJimdEcO+slQZgrdK2BIjzkfmbHznZj/IyqnXrGa5gBP10umgErtoyMgAMX
UQv7usFnzsNBiAmsBS5HDO2YFDidAtlPqTwQQybtvxOblAyc46HL/9c5eYrnWyj80jqfw5u2SHg4
1NG0JjSGcxbBRlvogqG0LVCxgAfGSFGbBL0QxCaYpQylzZNVT+Boqyt2f6CSO8H6jZMJiJBpSdoE
22LthFWd/424YxrMCa16f+6Lnc6PJnONwxoREkjPngFgv5+ddztguDqIM9FGkF9OjcZKqkKZQcte
pUpIcWBZaGlr4tA2BnnhvWsVtAISPfp0pIwM0nxghaYrKlhSpLHIUU+iVV/g135Dks2uGxV0R+5V
RBnd9lHG5BZ8NlvOere5ucsK2K4JZhSU36PGubSYDqCB0bWqyG1JXyn0rNdTST3/4j2F+84IGHpj
QPJg1L6NuuMcxJsZSJVTU5bcawXgghT4rbjnl1cDN3ZBtV4lOCMjN2Sv+fIcM/s5aoUwexjkQqta
qjRzoXcsTqBz9rF5Zh2x0dd6ao83fsogGckD7i//LLVbVEAX6QRR9ovstRLOqGTGz0WvUj6yd0Ke
hbfsoLvOp50DCi9qeFBdjHapmuZq7XbP/8FrkvHQgj6DGVNXCSlwQ5hwgU3WRHKscAKntDOBjTDp
rcitUVUaiZIKBhvQpkPOv7Qk+hlG92mLkAxHs+Stn9GSPKyeUYKYJXmjERlQdQrW1t6eUf4ZPHQD
BMtBHwXBB7yU7ZdjYLfBCTVgbdQ6cMjhQgFb6+RYTVSqz26NhCAERmQx4Q9QTfq9injPqWoRIE9w
zt8ca/aarlZTnMgqZWxKhez/4g975kBgxHWIqqSmQPCPH5d5H5GmOlpCPG1msqPl9GKfn6kT3da6
IQVq3gDZ9AXA3f7vM8laQApgYdlsOztZBgB6xQVXBqke9iwLfHXo7fWmwwnl6bJJ7Q6qzJZC7+AZ
Lrfluq4sHuUYfl0daAa9mTcr0v6FYIxp4V+R6BUUnOE/Snn7UA3V+4ga/YJk7VEHzUoegucKdrOM
NNjBDIJ2fFjnceUhBqz1lgXOUwAHPM2pLfUsQKQ1yxNUcI50LrA77IlIEEeivpS5UMxcVG3cEIP3
Z5fMg1xcm2bBZRNW7Gs2AcEEfF1a2BCLLk/jQHGXQmDA6grBc41p+bTBwsKevV4lurRzjRMff6+n
gl+EVz3wYJI+pVsYvaQ0RUC41+52I7glQ16IUtP3GHamaDhl7iy9fp/GIflzIHo74W7BpTbuT2Jp
9tOLgAlIWNkZCrFkImlOU71ZKf2b+1PLgw/3kQ+Uu56TEKX596FvXjKQvqbOuwSZjj3QMem7Nmt8
qDC6w3KskB5KOYXKyri1wJvwzwzeOBX8rIiFVMM0m33FJz6+c7mIO189RZmOV6uCh+A4AxXc0Fep
GyAvf0ExdNMgkhIoASNo6KDAVUhrIwjySOKE58jGEvRKTjeo3JnMxrAbmSYNWWg/nXmG6vdKlokI
nucsfEP7qj3FKOE+3Inq0WdQsyY/rWeSxWvTkvK0xXqDqKHSaJVPKUiDlTioDHwzup0O1fA4HFat
pICN+Cq90Ob0EAtM4aq/Cb3Sr0X1vvgCF4z4k+O3USBOWtZt84FMqMqAv/e9Jte77QH9DJo+HhUq
NzFX8ilOz18Ph680hPi4LGPlpc6gwrq+2o+E0CoB24NuVid0Fpwg6iiBVmcGwr7MaJIxSuwdgpov
E+bQ07OH57wysZbdpRGa9J7uXfmZyNFw9ikxBncN6uzQOx3hKzfTASqJJ8/suntLpnUn18nS6t2o
1Fg0i33k+SzsNzDZDo6FzXcCLSmG0WzVOmAxzcuH6f8NGaNiTuXS6l+dxKhQTuOAbBphASd3Sn2a
fR85rlqq2mP0c+azcP7kSPbaJNFiRJE62A1lJ8G5n7ut1zvKY5it1AWaiGOYjkTIMyekFl5NDITs
9z4NCTR+zk80yGPD9LoAYgeMZvW2ac6jYdrMj7cXwJQH3W4fqQgnnxPCtU6ALRNDHVio6+Puq8Sm
sZLxWWPLn3XYyQHlJ/mI3dbvUf2bEzlMhJs2xXz6C/v6Xa72AcAbtGYlb5Lt6uxKlp/+pP+6YSEw
tVB+B9CR/Q+5FAbMyizkTpFEYJ8ECbjc5ICHQVmSetzn9WUpHPFw8STi8evQeGYuU+c8PQiKHT0H
0EHDazsQ4hqdXFEgt5hXgfDrsmYCrBGNeU1girwfIb4Mj8MGVssuXPOhG00hhwMp+gMj5ybxC4Bi
3iORau+bfzTNrSr8jPAPIUd7IQtyEl80cceWNcSyDUmNXJ/Bnnim3KOYYFkXRdUAqRvEApX+e8S6
j7QBGTRTrhoOSxy+hyT+jIxyEM5nZslMcZOGGPSIE61cG4aJk5EFS4Y085afsuYkZNXiTOaX3ju0
6FLpCXN4eije7Sp4Yf77FmHukixptKNI8APSucAkTQkqs5NrLlxKlEtQZs3H36ZePcBjtI4hq3jI
VTU5tB9Azb0+0v6x0xwntA87BJSPc5+udCI5mgdoZchmuXyZFEbMgrDeult/z1Uic+tyvD0VbY4S
yDaNbEo5c5W/r5IvsyQ2VAnBoUb+SSUqJo12SqHgm+/HfKGrLbeKggC+IzWOLtGeo7NGe697VVTc
TzJKZrz++xz5xOdiVGwbgde6tUxhiWZ/FGt5Fngq+yJH083ywAqzZExAokJgw1yG+3eww+Hesb0r
2sFc10fuQlvnMV8ZBLyAga8XRQef5fN4XY/rEeQmWAHXMVN47yEPqXJQjFFGcK87ZYUmkQMhM4D4
1VMt9fvFJhdi4z2rvwAhSUsaP6+J7/EaRSqiSnSXwUgX1meEAXMt9lx/h2Hp5kCjZkkuuvRvIabr
b+HIVqehrzLnOxBptVm38AIy/EGSKyQYJ3GXiPTavkD6dVCcU0AHHM8DJbh2gO/2LEK42hgFsthT
c3k2hNRhbt+q0359MF67qwu/ExT7OrxGelW+BtAjIeE5VdoQsFJzTAfvosOlttTcCPKC6y7J09SR
smlna0DyZyMX5wIqXdqyx1zXRonfF56Yyt+WPa0y1k/XiIAzg9aRfo8TzJtObazcyEVcgHavCw9/
NR66QhqWr/gK4E8gzW9aJxi+dfTIdmE26zb4Rbcx7zMw+blBKY2GfEmLLeoYG4A44Pfw4HLrbbbm
G1Q9IeQVYCPa1jn5wJl3shQKRPsd83pLTHbwX/SxfTWFkdVQmXVeb8sEIkFJFSeKgPBaz9rVuHgP
r+sNVDj/QkeS2GMep7QjAguIdnjfCnvtYxhMuAJ9x264Q8bIpHgQjWyfzhs0yLBM50xS+tNExN9/
+7RFr3K+yTjt2CDuOmX2uAoaxkCp/wIUew8+d8CDtBCyCN+2AqiFWY+NuDDRHKf7buOyINyhSNt7
Q2VOTc3Cq1dCyhgQ7ZPryL04AECWNCw+ignSNcNMVNgXv+Q1GwPgTig7cZx/j0GhU9BfmdYN4AdE
EWbMMMjhdWzAc7Y59EMfWNQLH5BbjH2WgF8sxzb6p9z3iJWEqLLI1z94a6cAQTQhz43Z4imVq51b
tmd2RPJJRtQWc9TqQ+wm7GOp3NAn8jXc70UesdqwiawLmqbHIhEq5fRnSOVe4GO6tt0bOLHPcUiR
oECD+hiCoAmW92/6jTBQz7NlqNAzXm/cX+U/wc0rf39IKMYcNYbUvA+0laGLJ1agSwGl3nVqNnS4
srZypIcTlYIpRjUCLVzTVymhY2pEdbNMU91X8FSd41nzS1JS7+xWMUTNF24jcKXrcLslC1OBX2a7
5h4p9nXdrq3bxSRvT7dn8lFMBX6B9wROMDgsBrbwW6qKktZHExsFgYbN8/vjgvSCUoO7jcezPtyh
89edL0lm3QkC7ktxurIw8xIkQl3HrEGAfvr553FWK0XdYz/9v2Ilxnkj8Wt3VsxOErfefrI0UWI0
V2msM3v9i0/GnUIiTAQi/jWrv6BW4zVbrrmXxqq3rqwLwDeNDeyKKq04DIwHjAh2zSiVzKw8uUWU
EXy+NWm/yNuBYEXa9Wa0GmuNVYU6/sca1QXtYc2irRXy2qnSsc0f+0ALVwvuQNXJn06q+hcI5bVV
Kwi5Gy4XVME170nIQGBALz4vZmp1DkH042j0ogpFIU3th2RSNEtHW0hGvK23fYLSTEEp2bu7zSWU
WewTy3qKORe0Xf7ofoAQvp63AYDq4WteThfWOb0GunndCUFgAhFGrourAKRJXEE/2Bv4iZP2XvKH
GBv0d7Unpn9DW77qDT5bEMPSEVJgU40G2jcF0bN+HcT3Z9EP1RU0bfCMXZfpC15JlprfbMSVRpYc
7Lc3TWKX6HQ56eht0ZjoMeDl7JKXPo47Ik+GBc6W6g9HbsCO2xbN7MX5kqC5XVusA2WEIJ/vezn8
h/yM/CjIhBbU4T4A+Et8ej9g6IMi6zTvd22JRtfVWN3bg+jWTZwDvg+3iSFiTfVhLfQNR28dxd4a
Ygg28OAa5KsGtKZD1ME7SIpENXZf5tpzuSQjPHpOIbck3JaW8ZfSALeGlO9uyTheaOLJgt0cydho
q4c5kldbz0tIUPrM88MGVxkFkX4+yWXXQUm8aSHp9k4VTrz9H/hJWay3QMwk+/JVeaRzdgyGao5v
qzmJn6fyScgDsrVTe6xfXHuu7Y1jrY8uUMeipOhINhDDySNUjOuroDiJhAfOgNYfG3PNY6k1yxSd
4RpExcC1ITSGLY0WsSdGKvTxzUy16oJKtbuH6gU7SS41G7e3buQOdFuEV4oDPB+v/JncJKCuKIp9
0e62y+XEWb1nL/WuKNGaydI6RXrn832eCN1oh0IgiU0GjPfGVhpiyAWkpgmS+biVFZyUQTSQVnyK
Tw9TCZtkIozM4FdrnpNVZgJNHuLy0kSC7A3tV+2G12d/SiqaDkTIuq6zOaGof5cJVfzL9+gJX4QP
qx7R30fkPftay2ZNS+ZOauNjlSG9dttOSqby8IKouCDRk8fZJXEcVeu5oHgVDv4l6yoLeHEKfL/K
x02XJYkiGIO2c1cuGwZ3ySZV/cArKLV/z5d2hU4gAu4qN2qz6kW5MiwkbdrZaadPgeHMIeDIC+8r
/bO5oWrQcoljSufHGOkq7mLQAmj/GVUHpvMl4Cg86JWRv02mswxw/UAMtbX3d6BMBdRQHu6N7Xf8
VYAaqTkLWmf4yMS4rRIDLLT4QMGy+oM38JUjx6CaN9cbuI09tX9/nxkOCrEPOz9DaeJvxJE7m1Nb
mb0Do90aLYHR53NQRp4/B8YrWci6/ey+btQpzPVUg9AzelHtN538kicfyUC9bstEv7vTCwdmxXSS
k4jL116i74PC/kDcY6sjW/Jx0LsTBN9Ii5FWCVJdh0USMsC8mCkvUVQCKt3hrLXQ3v/GZeDy8ETh
UIVFxzzZ6SymvJEweyP607NJNrDBTniQERa1vge8Pu4Oj/oXjnk98abQTMMcKZGRjii7WJbCL/FZ
Y2mWV5DISdWhZ99Pdfv0QNlH1TalHAeJ3HJsVs8SVxcxrHOgH1U6PHl2DYps/fE8AQuJZj9ZbpJq
lMTvOqtmYWmBpFhHBdckKs78GW6egtlZxmju8dFlxreqL+7z7eKQxrKpBfQClHna21zB5Ziu8luD
vxuGIrD4aK6/xf9d92qRs2vOOzjEczwOenabmtcBrEhemCJ0y3XFo47k4yOLoxFXW8dVM7XdyUn0
I9upd3OKyRdR+H7M1uwj/OB683aQXt1yahTMQt47j5N/3BmkjKWbdk8S12LOu9GAbuGP8k1GhILj
4WBP5UEtRucqCTKvt2AtpmopOZPxVrW1lsCkJAR1LJTKOv1UKg4wguUYBKlKvYdkKmtyZN8UIF9V
FP/rr5K6fYrBZpvvWcr2bvwywOp7fFopqrnBak2edGwKKfMgswMdNzEUjYHgQrBFDVEwdUoLv7j0
60EdCdsHMaMWrbYPQegsXjXwY0TghxtBGyg4R1UDmpAABLO3/mKKRpkMr0l54+PCFNS3wWwjM6QY
ozvOuQYGPylDj2W1ST1oan0hna+w5TQzWA0K6BjKOgkBsYMjPy2OnhllT2KAjooDmMv7bkvlbyfj
4upmmfAt5GF/exTKngF0rglIG56LdCWkVKWuOIRPE/E+E4W0eqhLqLOCLtD04REub//3bXWDxwtE
p+EV/TtY5yDXhScF1D2UgKNcMwp6ck4aLyBUUVPBBmbDC0yjyZNOkqRIYsqkNfmnBaoZSaYyLg/u
+RipAt3kv7BC+a79JRg87zbdl4kwlS1xZy0EyzzS3tvvv00wP5U7eW5vrL01Vl2IoWPKmfaF+Gi7
qm17K167ov2FjLqFoSlRomcBMDwa3lWUL1cvfmFfNDxI7U4ly8EB7w4Q8MUxImjiz5V09osWW+6h
vLN+i+tvc7eJ8gTQM/fSUjrv+tDPugvJzkNSdkwknrfW5zjQcaaUd4hqNXdrbN8H+6DWpzvYJ7UQ
+arJT7LIuNOs+utYaxGp4HzJMCR3ZFC3Zxh0Hp/ER5eDZXpbcCaigYUGe6BqpILy5KOOUdU6ujGR
+oFUoy/tMPUA1kQltCXnpY61m/zW9F5Ej0ySQL4baqCr6/7zYROwwfZRlRTxYeqClbP692qKPfAB
mKzz+1HE/z81j/Xy+3O9K0+LLVi5rQD/gKxfLl15wLRqMx7ZfhBKebCr4a7tSAtllh2JPmXkpmZV
Rfc2w2X/FINoUUg17jr2KMjwmpqnumHwKlfCnWVdo8auiypbTQuul38RxzP25f6zT1mDzFTE2iez
rCtS410hO6FvZhRy3Uv8H2FMJ3Frw4iYctfjIRd38ShaDdFxVAXHMNy2K7y2nvoPv7Jkf5yq8XzN
GhkeHQIGxMHw6OK5ZP9oDn8MkNs7Kuajw1nAl3CoyMD+piG72UBDuyKO63Epw1gMdh8253Y9HFl3
b7mzYVwdghbBIRunr+W95xokt673pFtnOchltr3kRRf+Kvb2fNnsZm9GTK/ZBmVQarHr1PSxTpHP
XyY6409FlEQEOAT6pVzS2KgKp116qmH4NxZqKy44XKWNaO6eq+LuwIO2grGsxve2+BjGByYGmgHf
XqLhGq8OPQTV55GEr9WyZ37htAWlTlObSb7xRmK0ZvK7QbpatCh4r/AeQff8k7AQgRUkMIaCjXET
VUDqWbyix1gg9I3k1/6PuptAQjxLoLgDMZFE/rS22+MIljaLO8JGRQIer6mPw5oSIPZNTMyGqmnl
Mq+58xqgnEb56kcVqOlKrGYFu1r6VptQ0qFWJLDCXTeoIz2Ny+cLVJWnBwstdx0Ym9Pq57xKpHqw
NVKV99gh5ho0cfvnyq6QYjE/jR6Ag4LGpeTAruMkrLoBTxNIdp4wPFMRbdMvJPoSld5WruK9Ndgj
0nRlEY5gRKg2uaUkb05XDjYFIUB7FNCvfJI8w2OGR6QeSg96Q29foCK6eai1wgYsEwd5n1et9jvf
vM260Hoto2xRXdgTx0sIifUYlpe39moJlQLWS4cBq69LO1lrx5fsrPcn7LuTbf4AA+c4loyq/K5Y
jOsRgim0HDn+aD5SjLAHK3+oCAL0eLNZQ2sNngEZ/WscxvuLu6nfWFacLw/gMDKAhDpQaaRitWV2
i9ZhbmDmDzY09c191aXD+tN9ww5khdRQJfcCgRHm+rWF5strf+ZebZmLL1USTgtXVsTlcWP83qa9
xvBkQTgtfp2rSTD9fKiBMIVYwf0ic+VNMkIm2GdaT436q3xw08mvSn1YTR9VggnkzxfKa9tdQkfs
01xnTZRAcKwtqLCbcem+ALoY9G3JHXiWwH+qOf9xDD6rEmgp2NoN9XSVPI0GMAf8ng8yvMWCvbdN
cGhGgkzkxkj7/psVCr6gmWDY6c54Qbs3YbTx0jCXPUeCrr72mPhStq21ojahb00pzi1d3OEOhW/X
ZUpQSkk/9P8nw/dv3r6OXig3wS7qn+XZQFkuJT9GUHBq8rnQxNVhqmaa1Qd0iJfbnk58W8lNFYvJ
mIojA99cjs4k8Tnx/iiglUWt1rpf4sV5nmG9GSF/VzNsNosWvL7f8QLrLMbUGmVLqdfXUMYqHwHt
E5xbhHzZ0GY+0fRCW74DwOEfkk/60LwvVQSEqJE8cibAWvvNyokP9VRi12YvTCTZuLkhFq5Q7gr0
dOiY84vIImjSudOBZEKeZZz+OA6GQSQ+6GBBUPiWPs+x8nowkYYe4vM7/5BmHc6qqTAbpGALySTQ
KnUlVGSDtrdHRjqo9GdrSBT5bJimyUwtH2FlbjM7uqp86GhDB4c2EcpKtw7Z9y4Q561wXvGsCXK4
72Aq/zbVvW7hFm37wyT7/kjqk9sT1ojJVOcJPGwWG9VLhxDXiz08/Us14RoHQtTKX1+GAyT/v6EO
WlwB1WWk4oSH+JhqutoR6i9YHFwoeyutMqbpXX0U/wqtKaKAUEfMg5QAGud9HBMOXWDWaNUvXlAM
hMlzGX2LyUZhJNvd2uNMISHqPQUws0pG3rIZ0VZ25bccb40Dkroep5AFPVCicqswDnfRiIbgV3rT
iY0/eCjLdKru++eF16dANGdKGPblS0QN0eK/RJq1kSaZsDb2EX45UFDuwzo2K3OxHrDjRwewwG0k
8LMS8gPIBn56v/EN/DpNh4IxCGZrNE5HpExFphnmYVTJHfRh9j4rj+KwjYtEV0/y7IXagcLir60K
taTHLxuywHwjGJ7Pn/VxTlR2Zh421KDQFpUOU7eAJSmAh3etoUQRZPkiyutnDL0wh3kBL7NIYH4q
WVAmk9JYsVstZdXlfwDkxx3K8Gaw1fohXtmUY8xrePFS15MjM2OlFmC1wvdeIkIF7Gf7pMQhfnoE
QXbfHUYWwzVELBf2sVoBS8c52N1icjlzK+leOQa4cAw9xamK4AO3+KjdJQfOp4HX3aYD9zmDSMXI
Zroy2eFO8aUGMwuGFsIO3Ztf4AYacf86al79OiR9gjEPzXRxHPAG4ypthgk3Q0UeIXc7/cfXYQU6
JKXux23jDQxgue0tjOj/N74NkHUgx92WF6OYq7O7Y7Aph1Z4Xqi+JPp216aI/XnYq73Y6/H34prI
/2hoFKTRgsWsVG2+pN9zYg1kK1pQ6+vWlcdcxKcq0RKW0p29zM7R6dzah7yhUqZ+yCbf1Eikiv9I
JxDlNgOcNKseLmzyk+7RsIxMvTF/kAvnMsWXqicqpOpd4Jc8MXQj5cCsDSAGp1sPEoL4NhQOZaMI
JWh4r1fvMJsJsC/oUjOOiWqQNMMDxj55j88svpwBxBXXc/o1DxPKvhRzJA9UGdZtKrG7UCw228Ss
cjrNLYyWvmN1Unv9145x0z/barWuCsBRhVpWNBLiurGj+0S0L9pHVo9Tr0rxp0/kqH7gRGWUKx9C
z00WUl5JSxsFcQeMSTPKSRyUc/aqbW7kDsQ7ST7LGfL5mqhLsYZzyKG7InrXZmQjDvIsXP6Kd1Rk
mMUZ/o65/bcySzsEOYo9G/U8l+yn6b/PBLDneIZ72RMprK0Z/nSE6nuGkIL9q7pkaWSTpAjdxrGX
LvCPUob8d5O5UVoIvCR3I1OFp82PiK3ZLUWsmvfnB3wEroOUa1ISU9TOVgvIISszv2GPCNpOxCQ8
d5YTohlky2Bb8CgeVIDK7/OaRWElBI/9YkgJ2r+dgR8EWXGkyFdhwWZWyVBuOgXgL0Rg7HOS+TbR
WEp51mTitOzLzwHIAZB4eJHEPpEX7bVav93gzLG54MfYoWOm7TOElgObaOZDPZyjtkPZrmpWDIfi
IvR9dPQRC4RnTZyn0uG37rvRHI5Qi6nGTGqa4jnMTcKcy27MSDcTj5BXt7Lk0JOKPStXt4fu1COR
LRcSwlEAGeWN2DmPgB8cdj+YLJZh6dQqOBDMzOnTH8lOdQ04dvUHynEvaXhxrdkBmraxkKIa6BNR
MdEq8KBUEB7I1tW2rkW6mIShsu+VDWF4fTkJ6bdUDmyoi3NesAoLWpWjId8om5JOHGKAbA08wDvY
ZfKLYkwcRfeQLnCohE8i40ys02f5kSInSCTSfU84TV6Ugr8pb9GAmT7W905OXm3TdmBu9rzval0N
hDoyoUBaQmyrmtl8WGy4PE56+8HsWM+jKNWhaVEhyI58bYCSvHvJPXUWI+OsbMSSLeLEkugIaIAR
zkip0oDRix1bZsFAuUIAqmOyYr7ZUDq7q+rQqDlJz57ZpFquO+1zajvut84pK/JB6XHM2GJnUz1g
me2wFDl+N/lIlBKE+02NP6x3JrCeRs6hSWZlo2m0IoERet5aFtffD14/GY2dzgl6Ez1s3POZX5B7
pjpvL0aPirC+OIRfAaumvjGcmCpigBLZ2DJ1g2YT63rDjFNWxD53AA5NPQhs6LCadqFc/XLbYq3l
mObJ/FEdcKgcj3WMz34hTiNjdgXzVFy2i5IGDsvc4qJ30wgxSnTEqSzWlVQyHs/Wn6VDFnjSDono
nIjqJ0jpbJ84XYuQwa7cpohj01sajcMN8lqdbEXyVbQwAzQ5YCtaJnvFVUCLMxhjmU4xZ/Ft2wp/
ASMzYc7HXN55Pc57k5zQ9TYbJUtAzZH7pCInEnNg0WLctmMT/LR4kKOuqDMqgUDueiyVtKA9pn5y
Dt4KHtGsUfg0nr99WQaUkl5JSGmmf2QixUc5ZW39jtzZZX2dE3Z1tRmUh/rd2KJRTGM/1p5AsM+R
O7Kn7/iKBcMupf/oBDJmpnKwHYV5Sql3dsb9PeOhllf6wA7WcpAaBOOLHfZ55MhScRjuZ/0dGtO4
UfokpTXp+OPRZzX8gllCtjW+m0M5njx9yzupy6Vf0R9o+dm9lQ/6YmwMgXRh/Cl8aqpTiymV6Uyw
EuL3dqyWZ+TigD6sJMy/m79Qv15qoQRueI4yldFiWs5+jCZG47LVZpYvFzeSxQhFzaq911dMH/sT
W7qjX3gRpxK92hLjjxvVEb9R76fpuTvWVI0iB+nDBKGoR3L7A3rpEw6po0Y+pgpMebuRvQalnqRp
GQFNX1th4SP21QIRlGtua4GW1U3KJzBP/YFitaAlrsuJ/wWERH4f6Urd1+LhBSk6527dXehgPOue
ER4GxXlavobbqy/rDO5gHB6oL6sarwb39+sV04HK/sh/5v5vRrPsb6r9tpuLbt+JMbl/5AOAPJKY
0LaLfQV4/vwEL08zKinwK8pULNWwSeTfOUfAWyRgvM0CZmxNooSE2HpEeAbFhGDNDhQGjKdARGMs
dsNbD8aHEpRlpg586Ljo9t0OV8nTjhEVVZ6Mwa/EOJv8bz7U5XIu0zs2jnWXNpe9R+zZjXNm7qX2
oySQdt/9dVM2O1KyAq89Vx7qhFNMa1SLiKRpCMtijK8KCnQxBU+/DVPD3p13SE0L5pvxX6BmPiet
mhCU7Fu03I3/CoIKErAvi81aK7j18BE2xruiUPTVWRu5zXKnNzFctvN4LB8nRIg6MJHsVoEo5POV
ooQ/qy+Q/Km29jss+wGqORyz2YEfQhvPl4Drkh2MdKaCqw7zzLnFdzR1WYUjrID43R3BQdFt+lCo
2hT9drfPna8G/g7AkCCbhPtAG4Ni/gyfjzRBOKBMMi8ic+0tA+guvkORsuRy27qWbwWtQMOem3u0
yg1WCHpYAh2ol/HBP2SJez4zxw+IQS4ESyDfdiXBfogSftgbnvJuoIZ4zFzkSUHutfh4ma8+vV3H
AteILsEpm91rhCeJsuIDguSwXep6pCAdVuSOp61Xdb8B3nIM1aH4SAizdfsmuYM5jqyPeJvUx3OH
sjT7VgNv5zpzU1KCOqrT6OSB9rJ5CMNZcp/NiihNGPQCMF8hqPmZKvfl+MPdmTQC32WO/oKGXjUc
8XTMLHrxV7upiVtQWdmcCWYOa6/nUuoSZjSUzH+JAaHo28qMe87aPPTRw4omPQAec4+Sra9jQ+Ot
ze16Q+7ziGZM7JzD5GSPyex/x4WsNB5qpOtuzUveFbyWoV8sMDiU5wo0BqB0T0gLpHenvv8oNrTI
/OvY9B6MBZkGoBg64GUShp2sCXQHxCCNbkf/xt54C60ivT5Z/Lp96JnQHwIW0+QeF2XmiqVxLcuU
a7m81Nq1Ex6m6PRxyTQGdFHy1gXJNaCrheWzh+S9XiIz1aauQYvqke5cdKlx9i/+6ydkIYJfH6CQ
sj4giDwO8gWhil244Om1aSExiynxpBfkZLgfeCM0Xs5Nkr+ZDQDLFUgzqjqhUBlKVQLNzMcGv/3Z
EfS/ZYFRxWYRLF33+PzUf6UMXe6a6tP2th+DRcqZyvrlROSxQfAxMCMTtj75QjjaC8g+yicxmGng
aL26y8kCtxk7n7eCz1fPsCELLkHbYSwPahxzPGJFttWTuh0wvOlXKrWh74YG8Bez+HLqlSn4rAYQ
z7bO/nUAx3i8KUM0+ChJwxeQydsDiPLtybS8hauJqi6AdBM+pS5TZH2rJGbZ+FyCz7gF8xt8+sdt
DAk7sQSuEfgLykG/dkHq/wM8UDdb5sR8JcjAE717ZP/u78O3D8PQdQwEfdCvJtKWz09d+9uTzeYN
kA4I0pWB8AVXJD28MeqwuiWn8AzqR9XJ0qt8inexod32HdbvIOowDMUGN5qoQSW1OJzkvLwEuHCP
oEwwowaeYGN/KUVADRaWtUFRdzcZbQiy9Clj9mMlu+RcHUXLl4oA00uIxLSMyKKORqp4BM9DwwQZ
C84MATSe8rla+g/XB0+Gc89YEJGaEdkKWQmF56FYHoy5JzopdeiHQkXmg9SP3teXsFu3ef0/7XhE
JZ7EDq7KarrCkSZAig3iNhKdeLxzOydR6MJnLlEFK143oqyY6FfS/U8zwpE+8wQSRc35/cNijrDR
tABKfgxw+4pGxoOIuUWqiYttfxhXfT2+OSVm6jLbio/Jl6AA8rXt4DJJyA723r+wa0nObjKs4zX2
XZDLvIsJUjwNJYrfvKQiVIpjJEyv9XQHElawtdSk0djAbf/uVh1+CPIhDLL4sgTjdz60lKCOjH5I
Wki1t3x6aOCcX+2B65S4IzGUGvA2L1w63zyXzaQ2qqpjoksu9I7iN08OW526E8BIEJs75vcdTCnw
ivHgD+rif8BR7+JkdB8Y5/oB5kbqfBrHW7wiYem1T3VvRByN8Ullh/6I9Ga4LHRxHie2Aipt+FWP
NuAZfSFIHSRrG47mu+N6QaWjD/eR5LtIzH8HKQM1UAh2HY+lO2Yp2W+RJSpAf6gEnkBxPjZcGN4E
IM1gTsUcK+toDk7P/usw8v/fjUZQBTD+SWfBpjT0GiTn+4KwaupY+3MNDEDZAf4YThZHZCiRHdpY
MnT88Q9MM0iQUPFRkNCzd0rwNKvCdWtdZQDyIR0zcyD0yfMohyg7QfzTXdQefgGDXUsJA8S0u9mZ
iXoqm/eyDl5IkGWhDZB1PRtIgWBXspQKjCtRIn3kBOYo7bXsOmXg61J43Ftm2PDuWFC8Anps2f8v
637/Xy5QAjevw0+NhNX2Rx3n871yhm7F6U0On1YPB0H6LFqjCLHlB8KM8zvo0ulp/mVlYujjia8O
74GyodNM6Hk3S56Q5qjxNzuxg9v+5IvMAv21ypo4G1hAnQdnQhlaH625p2e/5RP0Ken+7+TNPGZH
AFCgn0/aGhw6H+2/9T7qpCAOGYNfEFVCScARjiPjUYI5myyLN7INCNvk0I1A2/pLqzWoJltFpYYS
kjHBmfqNbJYVKrLVAX/Rm1soIDhHgeKPAOKYg7g5qdi2/t392gUWiRk/SZCNJOJLFhRVToze8kn0
BuIpuZSs2p7R75mDZUQopt7wwSYFYzPddGPtDhWTEYiWNni6XHnLY9rNIuBBlybII+b93WRUnwr9
yXrTO8UR7Oxh5KeAMfZ/E7pj/PkeiWIdYCu3Ei37gyBDMUCSAu1Tqi8IPg0e9RKeub4f36xSTtUf
shZokBaKCa2cY5qsf5UsSPSBXtjhs+NWQEAgmQjfSiZ5qJXYKvukXnBcSle38t1F09aWl3q6mSPK
7fig+O74tWzdtaS93HIweBr349R47FbmZDwJQAHw4CbxWICt0Vl2dPwmcIzCEYxonkpPBkkoHrz3
lQfzaxsoJUOQjEibFoOkFXnG5je0/dIHFe0VllZq8BEIfaFuZLKj+a2RIF9hAj/Mz2UiFQQBc1v2
3cA3l+0eFZAsZK4QygcFO3l8HPb5W4m0ooQ0qZUi0BCweowJ+fNsbxSMu3P15lkOHBwjPTB0QHF+
G+/TLEjPwd8o1sepwySRVGCAxDZpzp8AncZFSTHrxYHkf9iw3lzvk4AE0IbOHyVqIiXSyK8eVxtQ
d1tGTqKdIAnL4FkxfgHl4zHmo5+FZuJJhV3DeKjYzWntbxdwywBM+neoY9WjWBEAShpAqskOHXdC
kB/9iI4MXKx86o0WREnQBKCYjxQeT2wjYk2uuKdWs+VA9NMxVRA5xwymSUPDFS2eMICRDYCxyvh/
LSt2KUkoBpZSYsvsQlyD4Mm1jGCmxj0Q1Sd1ObEy6GJIGiJlexdjh10TXeZgpnvCJk9asrkNOy/6
d7J+dcMRkGWv4InsFa3lKyFiOUbM7FH2T2ruTHzM8nk8ennS8bl1lQPhtU24q5uzNsHA8WYIb6Ed
UO0JQQ9/xQN5aLNOE5Rcnj5xKb4q0EX8zsOcF1SWP3PESJLcewAhKYye1Fuzn12IBpcb8BGzURB2
kJRC15RFjmcFEx/LWzFlIsJ/LXt/P/qHM1g1ZYJRRUNCVljxC6zzGxGTwWP+xDKGoNIxTVMhChn3
zlhMFm7gJ7fQkeiz0rGXjOMdJSQ7dFIVssUzoHijk756YrCcroPHw+iyl+8qna+IAxq6mFrTxYDJ
TLViYcu5bI5G1bKEP7kaO44eeftkXPifZUhE7QSLjXEC/GXs8b8R45/AXopSkmMpSK0Ur8c/RqOg
sZWuMqltEWaWx5OMnXAaRM9W7X6Ko3VScnw975cj5QAiCu4+dyY03p+E0RTct1k4GsAlHh5VkIAK
6/PbP//lse6QkxFDSo88OQ2gK/UFSCrc1VnUy156tpt5jypjk+xI0SOsz+wg654pJZEUjciD/fp5
0PtPgZ4vxr3JH2bKDNKerjbsTZyqXb4WoUzFx4kk6CoWJMuU/wR+zhSxrQQjpwR/fuzWx3o3RrgP
bJB0yuZ8rZHK0oiG+cCjcQFOfbI1Co0HHO7veMgd56KbePrkDasleDeqiriJP9AKfmCmhFSoif7X
Yeo2KML3JPlkkl37zxkmd+0/wktu5tzqej67zbzpfuC6og4dBs5jHzTIur58xaaMPz3I8FfamWPQ
h8V9vUkW60aDKxCFsSiWLpquacD4C0vRxQwkh0RDXGinjZp+ZlToP23BZZ6F4Z2Iwfjb7lK0oqqJ
orCbGL8ReVw+vjKwCd0nRUp9CXo5M/lZpo2YAIzFio80wYF/4xuxwsuFvBYeh2h/lhb1b6PyorTv
USakz/m72brfRW97mdKg4pZzJdyUESi+QKlWtAyAuoS5YvJKpipoNdDgwVRFoWr2tQQKcVh6CXOh
vtAWwcpeKxgrLW0f34acq1J3bMtkqtqzTK7T8U4XNtGAz584hdznOwB++/XA2XZbaH+QlHzMzTc6
bri8Ve7wY63KGpROmaYJjT5ONp0rcwPfap3VYcC97Lh+0qDbRr0sl+mRPqQNiS6zhHYEDPHa4mDs
XP89op2KMQLzH6VFQIMpTv+OGkDICW6UQTHCz+Y/JKwkCoZO/y+1vE961FDQb1XwX2YDzV6DBxJI
QOOKUvrErCUZnWHeV5Y7UaqHxWlQqvZLcLMX8soxLaVn0DI6E6bv5eN0lPpmGMDGONGRA4SEFjHY
/Y8dyzu+3ody3zi0WRcmIHgAkosRBxA0H5BLcO/gmKop9hu1qQYqQMfHtROxnnDc4OGsVESP6LBO
U8aKKiY6mEgFR7p0egY8FLcORTfx6hjpvqUSblKc3ArTD+XwXA0f6F9z1tuESTCIRRn0QwFVikGC
TRl7l4KguJiJ3gsB8AMAIS0mb+H0ocieMOv9phLSzHLQ5azEgsRC+O3iLKVnXNSQfyNTJNBsZRRL
xnqcS0dcR29eUQoeC4flIoYMHJ0MTfu3ETbPAfeWtky2Bm2S9qVuhppwrsHBLoUAddPHUXt56oHN
0CzzW2BBpoudMH8aQqK3T2QvhCLVIcnRxIogtYkAV+kQlYMyxUIA6lLiPdV2a4/zvNJ6+vtt6H3Q
/jFokpi3aPcBLhBoq5Dy4kqGpwFJekiQ259xDI1ITmK43BOHf4wRCKCWtTh8JKHh/pJxw0BQUxrG
1jlnoDSKSblFmYsvj1mlJCkypp3CEvrnk/DslO9QKqP4Tgh3zAeIyWFw6hXDf4bkpl5LnPPrbYoK
GVVXaUWqhF8IkvFjugxaH91xFgOes899Oondp+AmiU62goiT+V5LqttBMwuo85p+xJ7magXi6H0H
lUfKq70hGXy9zr0CDMbHTQD5Dcc8t6HmzsKV2FSwP6vkDHuP0BOaQRmZf69qak0JqLLjZ7X338Kz
hds92oMOo5YLY34NbCHwboCeASAKvD2IDInxy8A9hpGoQdc50wdFs62AW1VYrEvp+QgENMrMFn+K
AheBIxqbBEfikDZ4feJA0+7toPeaHe/IEYnRWop4fXpDplooNL0/3x4A949qIMwIxjLk+NMfq7v3
jsZKlif4BeCS5t67SDPcyck2TEZIdBwwr6fMjSblKNNTw/uSaudLXpTc6SFCQcHrLtz6/Kc9mxx0
NdRtISUBLOveXZ2o1ol3UcDeh19uFEJ07AX/PQLHAYFXDQa831VvvT/BgQc4VZZ74rrZMWpC4gcF
LsMwtL4s5EoE7lEj3Esmofm2TvjJKBnhl4ltSBXUtGMiSBn7SgMcP6z3/tjGn7SBtYpfJSiq9ZJP
QchBksfx5cOXXyq5iFaxHNSAYY0OvaK3FiXUSwaN06QuLHhFiVEDj19aVaJ1HyVnJlkp/Uqc5bdB
OBs0HIaQbzE0NgyM9SZn8Z+wFFnUG2HJA9XER9qurajzGbb+lCGeVluAbPP3y0povKf3FkMVb7eu
dqNkHEll87vBUdvtI+pKueLm2AHMRVjd6S0H/zEEeOfJMGnwj8zGESc6EZ5pDqEoRQIvnjg7m33z
Pq/5xV4chwE7eZl+qhnd23WTeoKfj+ac9jrf1KnluLwEkilyGeJYAs0wYlmlhN8Sr+FAgYylFubn
U02DWHOYOaQ3BekStAja35Cx1Xy5MmUSbJ7GvqtOojCwBqfqyrfBpvMb5g2QCMv1vLW1IT4aZipx
xQYeD9QcF4VdAtFGl1jeG0chfK2P+rv+aeI0tTQABctcU8Lg9Qr0vSP+CPPy8Txa57hjpj9oV4vM
dG66YnwiTnwo/4tBmtwgG4HybExzn/U35TNA8bp5Mt5vly2uBber6D3TsJnWKW0M0nS3Jt8GkUJP
NKf6ALKKHmMb459pHl80xqLZ9841Jp4Sz/HeiaFDqLaS4260ssSVUcW+3ZAX8Q2iVrU7kXJAl6c8
Bhxw/CHT7ovMwR1cSJqEkqKORFfNL/qnay2skwKTBbwJhtiPU1jPWM3djgkn5FfnOrb1Rbj9LQl4
vvAY3RdimzrpBm3HqycQYXsw9mXM+xAzhREuBhsNUTGJewVbqfucHaNLbBFtumInb74o2S44qVa5
Ej12Nb6GMTu2dq69M6z+p8nLzx4Q3fCi14s9vJpFsuQ1E50Ml9WWO+XGoCByInSftP3/7ePzHM7i
uuuOeDXdi16Xp64n4bJphT6IWwpYBLOgFpVI1aixohKylNrDvIkaSyIrNEeo9nefQjiQzwz8wXat
/CaA76Oj1JVAUXDGbvRNSntBj0tLkfOncNEziLO6Ra/+uZGlFMwikGxQfFEb6PByiEGRlf7PksaA
IhdogUlCzscBOvj64hKLXbe7YexwCtvUBw2RPKaR9jt1FSzfTdBbUGlJ5UdV+Y9WIHrmlQ8JN4nQ
EdHei4Ql4DVa6YNgh/4b2IFLaGN5kp71z/ftFDk3v3oAmPbz7yaaRyYLOcseV4RRo2sFlX3GaUJh
VutKELFOqGEQS7HYZyww1UstWMUtz7fJCaAeyECGGYmw82aYqMJB/VoNiNnR9aDVvBQZP+XculDa
TiwDhoJithmARmthuzZpr0F+c41uUYJTRYInWU1r/n2xES0/Cp0lI+L0Gvq2vHDssXP8rwnHciUy
d/ul/1RjhqJmnvfWuaMk2LF/9yV1WYW7QSVZn/+FGVej8ypNRfNO7vxwoCUPXWZK37ruxK0RJrWC
HY6X+BAFZCZfyIyOmLW3TE9Vn58qdK998u2gZN/jD32ijLqCXE82Z+/0nKXgt4J27RJHjyIvYx3i
b2Cy49tgSJy3hgf0WGOP/c1km+gDNHE32ZVhsyKhayfngv/h9eQPCT8own8RkB312sWSPJ9R3khN
YQyCj3sGu14pRgyHyCd/BRKuzw2oA8qYWxbkbX1uP1aIKzPui5Xnw9N9RwkJEG2fXpdda04iu+9R
NtVWRQ8smdUhWWtU3mnDeeylmgN1EX2R5m4o8T/PdUjJwy5BXhn2WmIa0IPJFd14UlF4yVRPd1PO
EPDbH4yZsJ9EAgvw2bcyC2kzW8171yIIyWk8xt8m4U+NAaZJP3EaL2siX9vhvcLOpwApvuLCyIbK
Qi0btq/WEK5H9TLm3QGprLcUr4SdmjVmuJ/u7zzyYEv/lkWOb/fLzH1Mb8zUODukptmRkn0dYeg+
Gn2aVR2APodIrqsxATAllfXGX9PFoN5ko/P+zK55sSmMIHDJKAjgVXAWjFnfhf3vp9z7Mp0brAKt
ZHWDJcqlCS1GkOiCUnUa7G+oowZPc5DHxPDlu2OVi70gLSyfuWmPpSveFGwf4dCFZptvFJ8zefMH
3pX/K1+gdh5ReDbGpTf1RdZZwjQN54EXGeTqtbgzRsDYXHsDKK8lTOhnVXryWoyW8Xc7xeYb1ZCP
1cmfUN46mMoeYE7lHS4fTpqPoKWwjrUihcLbctBpgk2GobaB/vxCLXDwFiIZLYLBeRadlYETJdhx
0nxzNyGMTsJvai3TPCBA+iqqctbfX/efxfO9N162QAKjS538DcR7NGATBC+YLb/ClS3T4ciIaWRj
+pVgKXPPnZxu96zeNzjWASdmeLxJsqPhx/0MQ9GjSDsDxgPW/l6jG13+I0jpzxFgN40eFbHz7hPc
mBJ5igQhhY5H9diTckleFtTStF617Jrs4PHstPLTzQV1j91bkpDe13ElULGEFEZncjWbfIXL+Q6b
fDD7w+rveR0Z3SOvcfGt6tWXgcu80LRz2Qw9RMfsi0+NUh706Pj0mO87Xg/Y02sIhHHKn4cJC+3a
n6sFiC9yIPitYSGmtaiTpm0rhq7ulnFUuJjTeOPznuCyDYiuxQ5euQtfveGl422KOExhPmLg18F2
rhnaTOqSBotDGyQunDnll8f/adbVAIk8cNkEzCCH6P7j6WSRJ7omLJpqIHTHejmpesxAGxsc+Yui
K4pnt+9H7yWWli/bt0u8/0DnPmuAJO/i2bfUdoksGaP0b5HRCbBQzFfizK+6ioC1RjZW8+CAT6nH
4K1wEpXtn57VlvOuI4XFm0GyIXHgvxY/lIrB+gBipifREIXcb9jm5KlCC6nwbL+FAllg8IrRWIAg
s8Ozlxu7Ph0GuRG97aBqwMAd2v1XDJ0Q/AfnwCWwjoH3nWr2gxrOs5ZddAQBab6ioRBHSUt+xM78
8J1Cs0j7RhcFFCuc5J0Rtt5g/YFSesv1hWBn+EnjJaJiZra5GC1+nbLM40+58T7wyFeSH8KrS253
zSTL3ndf+sX6IHbZowep52FTa4JzTfaYzTeo6/tc9S/souOh3pnbpbWJqo3W8Y/ZHVxrQu7Gc+7d
kDGGE6VZucEPczsW/CFZmSA7jKhUaLGbNMjKZPNzaKzPlUZs/IeCxXRdODfBy2HinSwNYFtjSXPc
bsxRiVhGB3xdPnxdQ3SJ6Z9aHCBveCsTGU+BxeYsQ4vM+Mlt1x97QYLz2HgdYHN1T/huOzUCURI/
CwbivPRmqfXEIHyf3oCPqAx1iIirMv7aBJsoQrjEr67jVzsGSgFZe4zGL3yfH6A3tzGI42SyQTYn
ZVT8vptWuwHpUfC9SpnypYg646QUot/UQPpe+V5BMv6ysjF6+dJoYn/TsVJTz2XKbYopmKVybXAR
pwkANvnNx8PvqLmDSqdGN9UEU82w2HdISHYa2EGEJD90Vgj0YXjt3R2tJ+b7jMV0xg661NoVpNez
1K3xOf0A1pkQgLoeWlHYkMyH3JOCS4B50bfTjdAsuQd0mjV3svAyh36yJAB8pA3OrhIrX+IuIMKV
ZI5SvFt4HUgyWUb4A3m+4FXDhtqgKXNtDzpKUBXSEl4UPjT5aNYZLpN7cNPBDI7fD3lQPvSDoO51
i8hVYBZz5ITPtURJzjiCeyVhQ/Tipw1wEmrYUnnaZOhpba8y+iV9iw5ZwLq0fXjOwor95uTAFNR0
hnxkvNHPe9a6uEzox968fmHWIMYoDb2ik11SaJyzZdOdETjqOXkE8pEr1WpowMG6VHLC8/Jvzv68
icQG3YJPBAGNeyEFR4TXHlw+bInXh+NWRppu+RX+Hh/zT9BxrKHtq0o+EXvUBQkaxTUQCcojOfHM
YWy1dZ1CT4SpPoOjRZFev2mo0FD2aAZhE5w/2KZ0sX3lO9f22Ixq3vAENQOeFNzfvQehHUn8wNHu
s81URbQkm/EGIbyNW9/mmXPwynH+BzrogVAFTn8NO3Y+i0OvpqNotducpKCAysLu4q5akbUYvPnm
z8NVSvbAdOt5fpqtbLmXvTwSDTHaH6Xg5Y6LWhTh3pQXX6W6j6kmuSAccNb/nvwFJ1d0yofgJB5y
aQEI71BzKyKvlaVdXmWJ95alRrbZdv6u+590XtHBVKJ3+/y3aB2OSJCDpkkww7zA74nXx7VfmEYW
IOxSr8xq/v1p5TOmf53Y3WDUFI5JxNcniT4Nq0q95vOuw95tnez7DVVkh9v5E9u/abo4IifspMS0
0phovsQyNUX4emzLc3d0eKCHVjw65wm105HghuQdXkHRUIM5sxJr3kvfuKmD6i8mkwADuudTTtAe
/H03jPJxKiW4vWe2YRwK94NsNb5jEZsesnodnRTRvwN+pvWVggTDCnnub4lMpyedQfHBpUYjLJzH
K7IM5bALnkGOy4wI4Yc34N9LDQfN3D8g0G76g5DS5qmxVoxzDXTlsLRRreOBS23+03fTsPMPb++t
4Q+KkGhnN7sQqr4aay1vjEBzsZVqCoR+5MfN4IxAuc2bHYJm+twUwivIGpeP59rO3OUFplQVvDjk
knGfchGIhU4xewr9sIwcosIP+aPXD0JHSLYdSycnsgRp9F2ioiypr4yREFxtik0wmBD5vAxuXLku
GHLiuWpWttnjqcyPeM+wTwgzZ3hKYA8ptDXZaTQ5EnUIX2lsnvG3ZGw1eA97bbRq06ogwO9JRwjL
Wv3KKCVqQFf/f8jRYJP+EfKeDykNo6g01bvadGGdWLZOas5cbJ0m2e0VttdVHhyvTE/OujfOzjNp
C9PvLhXnyp4wXQES0vob6baNv3yvZlyC4ECS4kRtx78s+p1LOMKejMTFci0WWs2fDhnkdDJ2QFVV
j0NhY5jDB6SEvQ4jbhcDN9jcqU+lRNyFxh3LkML8kqX+oTqi9INKWu3/xYOftmVLcmWC2hU5wyRY
tVCmvzddwDhF56y0TlPTE/Y5zpRQTuVTucR+t9KX6TC5YiCdjq9T5kGB7YKvOot8WoGWk5jeSMTa
AD7h4G7JdGxQd3EKtmEJINMT//NbaWRRJnTo0lKdL5x4uVF8wVSJiXp2djdSuTVTuandZH0E6eCi
uQu3PeAbF0xQb5xE6XqJG67jCZhd/RGu0Vl3m+XSsam+dOZsbi4ULefty/2/EfgR+jh3/eM7KDww
ZIfRoAQeE750sSlcAxtyQbEGFWxOaltVAGhs/w5FsH9IFZPIArimYwuxl5wSdxk9dqzqiTognNSU
vcAsU3n1zNskp2BXyfmFmA51bBP6GBb6Hs7+UutzkBdLu3W6p78r5GbbwlJ47KPJL9+Uupxkfm8e
+jfkYZpoX/h/ckyx8MBoyJEMR4Q7qcUMNfyhhWKtCxTrzUB7uzfr3tETzN+N80sDxB2YTXNh3NGR
zl7fFk9XOW0m1efQweD65y9mYlNbVy7X3Agonh7mmRwKl2c8gPtS7e+Z1PhCrKdMPWDGle9BVQzk
z4FEwXlkXXuEEI1frCzYYdpEeex2MeP42Hgj/1zsPBFgxuDaBpcPIEOgSQQIlB40c6Ls7ZPChqyD
hkcIclZ1VKhKWRw0oMGtklGEvz64UDBukXyFKZndR37u97/R7isq6ptel6LRHP+XNIvjAEPN7V+2
Oxhy++ddNS4NqC4wjugNMqm9cMCAIS/LcxFJt3Rn2cD3U959v/FmMXez3JJtlpeVHm2S36NLXbVt
HXYgtNOM/6Y0guLU6ezOG33JdqPYoXArxd5PR/QKYqjJZkY4IskA5M6knxpm5b9MaTqU3iBKE0Yz
Ecz2deuO4+H8WRxG5Gxm21BRKTVjdfliZY9T8jPm4lwtltlqGS/9WWvqmGYVi6U3rmubK1DZGAOK
7WY4gVtkNRdss3TbMQ57do2z+vBHij0Co9DHkIrvOVfW5G/HcBrHkLGO/IbPQwhILS0oebiDspb2
3Shn+1wqRC39Dm8/dVeU9KQGO5VXXqTSBZvmTnnqx/Io1dl7e5CC25zjC+uV0ai2RYmafVX2BAmw
QqyihJ543U3D4vP3hBXZH6udk/wWA4w+nqVtXkHKttFDUSTTHfDZkgc6mDC1gc+lezNIC8XfEu6g
bdaM0jtP2YDBw/it/f/zh1lnFF0TFV2n44/g2LzND7mEaCCA9ukJAovHh7XsNGla8BLuRb/39HCV
lYLTOTHSgn4QSwMrqLps9xfW5OIXz0lMrbfr+xWMW5NU6TF8aBgKdO61ySPb123aNymLz2PSIOZz
ZzD/TgfSLnXKvUSEMssn2TMpO8lR3gpBbfWiCWCdRkwPkeZk4TA9gKCJRU+u6LY0LimEijbl29I3
WB01X7h7lDZPOIQSa+Se8sKIg8LJBA3c7XYlf/H954RFDf8b3zEJ/SeVIcx2ak4Jh4KgYvcUQ4cO
fVZAD+spWRJwPeyQgwxqLYdwGfRkSxRclTv3V/bBvq8/Pj88EHKWjE7O4WuqBXDLSGzZVdJ8uaRe
kEr/5FoX5fqGrTn+qDled6ezq6MtZlosUYl25xBKUPMqMIEtZ3/qHfQ99DGwaD41IWKr38LNHu0+
tLG65g6RXHdHrizQNMgprgYVg5iY3I61XWDyEYOrLM3yp03+f1HI02AAo4uRfIUrLz0yg0j5itaP
EzqIhHc48axupS/AXlFTTEcZmAWjSUIlg291D22g2ddiB4a6wWllJ4X0AhvqoD5CQvOc0bRn3aZf
L2UHqC4B1aPBQNUlFjPMz1tUDS2qc/RBcQT+zo3l37HgtHfBfINBs6mLUiD52BtWUtV4XA5wQxIy
cD7kcBibjgeK0yyTlZTpwpumZJUTuu8Uy2yWlS/AGp9TJswu4fsnYmZ01k/Ea3WH6qJ8Xw8g4QsY
GFxOoxVV8VzWKEV+Nm26QLw/2jRnCtM+U5jay9u/nr85DJsCTlQaIVtlGaZ++Eynoh/+T7THeI7l
to66bm7VFOk6KoK1imqGs/KJ/943+mtwDGKV6pzzIaY8BPgWgtDd0YZ8YykAbLM645u73jqvZ/wO
JTVv2331V1ahISE9tNjrLVWYbwStuCfFEAj0Wa+A0atkIgjtSppXj4PuTTQDjSFMFsSWRvImgB4L
SnnvMRDpVyi0zlmfHWfgHPTNn+RK3S6F8vLMqxDBkHfeDR+6VyXn5buRnxEikcfgq7dknPaCXOX7
JA6FZREDQtcWOH/4OUpXsHLyxtQ1RPpM4f7LvdxxUVYgr+GWRQ6L/WEeOhuFfHUDiqPRqRiU8jFA
ihxdE/xdy5cBXZc/Gx+zMhQ1r70Ug845HTp1uieY8xXw7sKbUhHlz/i7rL1PChSmTOjPttpSqWIa
2NKrcBOsnfPS5vIIMNIjSK9Pph6gXEngRaxb+oITYe5yxxez0CV18+Vpf/oxayzpgx4hwHFZKA/1
Nu81Vdyon677jejUdALS5ej11eIbCvgpS/RJUZvW4OWpJoR8yGWnl1CL9lXZxmV0jcK4cnpfrXCw
yoWQ3MCiShPDFTi2i7Sjcwkec2QPve3pKMtn5Ob0E4QzeY931LZgDwsLBAVIuFxk3C0/VRqoDd1u
me8thoW57bzxr5bQ0BjXzO2hbSyLmNVctv2wWu82rftnYJL/LFyG+rwAGDRu1nbJ6yw7qWmnG5ry
F5cvkLoC2OJKAZoJc+fvpRQ5KUV0kmuEUwDVTaxJWVkpLwgGYJm+pSJHPb2rFnUl6hkOCU6mGygD
jlWFyDZXvJydRn7snCBNNos29s6fskogIIkgJd4Gx57QDWu1j/PDgzmMIrZacz0pbzUDdo+bDzD9
Hgd0DwpI3BeADedChQJtOGI9+UcM3WJjenkfp3yZJTZ0328eNmmw4HePQw1McivyTKlWwhB6PGI/
cs4O1fdbR/TXqcc9p9NG1DA2iD85bVpuYE3XOf6aOB26bpA62eAY/cZrPGZXqINmAwORO4Nzvrfg
eHwnPtLuU5V6mqh/j357V4bbIw8zwVMRlDPGHLn97/GhnZC+npryaVW1jI/N+UAozkD3w1CVh7N3
BpM+ZqCZVM0tyEZveSqf3+NbvhAOrDCZIYkFFFAyhYIa76apKWGzF1IUcK9FYw4vr3Ekwph7kIj5
ke5w8xXyyhtuEby4U4mrR/3zKzk+/rOsy/h8x7bGY/NMToTmn0keOonmDwcdUH8auGbzBr+x5aNP
7X4aSxfUFRPc8j4qX95FcYcL2Z9x9jR3GvwFzsvXzgIytHEy5eu3OGEP+CufPXBI3aJu89DTLVkV
NjU+e9291ejMdXVpuUnjgMX9wjgQ9LQUsvF7UJl7w5Sqr84aJ+1rveQxGRrHNEdTkjNk59rd0XjF
zE00l3ZUQL7JPUZamexclx0FaQ2VtKYaywhseEcvUodX4KCHY6/msKzISRlHdN8dqESfnZU7wP6C
p8uysFjgFOLPLsURXG2/JRU2eUIYxiIiMcS2hc79tzuIr0uXpsTgmHDg58Ecjf/DRqdBnJdDBdpk
c6/bt/TuC7/mluY9lsjaqJuEbloS9VP9rLCMywFbKHGHOYOpdWNCLvRD0ty2B7T0B6p1g2EFi/zb
FycahKkeSMxY7uulLG50OgF5WwJ4X7w1jatWD/r+UmReWSB5vPmnBKPigC5uZEeZFAotrIJGQat7
pe2ibTLZnHYjZCSNPgKlpLuUDK3CKs4mxUcn2bTNwF8fGSOBpZUlWcYjthI8mZOYpywCxlz4WE7j
ueT+7AdC3KcNT2igrWZSSnTPXuj2AziaHqgNAHvjopj3C5xcmAPZNkRYNgxIV+hClqlP6/KrU5wQ
78lrt7iiiGvMjsz3wRDv9MDEPX3bguhqpZs/Sqa8ycU2R6p/zO3qIHxbLAjWrjzJey1ugJBn/E5O
6FEHev40AeuXJ4taiPH/1lumitILWwtk6aBFgb2Hm4BaO2X/E9JRMaq6eeLgHu9oa5/DIusGHsi7
NvSbLI4naL2nfxeTp5ohsaGFtaL9Pby2v1htas/PUp/ewV2LF1liNJeQyyJZAN8V0HCbgZTDwFJG
Ucz/KgbgtC9PgGgyj7NlDXp6GCn8JTgr3+jXGH+gXd+f2IAIK6EvDd6rC9w14LPlYvBPnX57qV0f
m6jx20qvYv+eq4Y1nrFyXUmtImlU0nWds3ZRDq+BbSNpRV3r6nERgBWognHmXz7ehMmjehJw8TPx
scjea8wpmyRCwnWmqEvwthMxVf/HrluLhOnIkit44V4n4sisLly5W31s1zuIBMPgt76FXFs0DcK4
3BroLI3ILQF99cOaPbbQ6r7FEecqdhoIRZMwY5HI0OGUJKLP+6k4YIdpXePDFjaLfUl96s9ItGwu
/s/pqWuNJUNV4oUbeLZU3LKc1iuDIBTwywElliHwQqL/Yd5o9IPaJgAl2+Wg4cjzNboq3/yCC4Z0
nKM236VH22W+Ej7dG/U1U9EDeXbC9/ge76eRAiFXoJaEJ84gQmVtBDEf4hP1OwjW/yxSMwfyZVRS
edfE4d3CPagUUVT8wfhe537b/XF79Vr+YZF90He0mACDcfAQgf5JUb8LEkHNmaKAHm9KVEgVocDD
Li+ZIc8TytER7hNpuW9j8hBd4JRlhI8PpxY9VNlLh0x8VN575oRUIOko/tAZhi4w2DwLfn7WsU4y
0prqe3i0wRFmDENXszDi+d4xXmlGxGT5uJeJISYk+5caZ2MjIZAn4lBqcee5QOrUmKIAmj7Pr2Dm
rdl7bERPkyAD5YqGiP3/lsY3CK4VAL5LHWqqZ/y5L/HePWVPJCJPjR8BRu0Z+HemdTTvCaQO39rw
E/NHThwvcXA6tfdeJgJF5R1bB1kurX7/X8sOQloZGEGqyaTM6CvK0AMI5paO1XUbV9LbpTjWJzOf
G64JHTEmgTu29ckhahZiqe6nam84ycifhA4M2w46XeghfzyU75FZMngVHlaLw+IXAfbL7d8KOVKP
kzJZxVDLb6gj0IoVAwI6PU7RM5mwycMxHJvkFGwoul2OiRP38m9ARR4c+3bK2jcze4aPkeOPycCU
xg6Gb4pF5gxpw3vTwWoW6vh7cY0AI8g/6Q5idQc1cHbHsyDGlF459ns99Zov2aPbG25VySjayYxH
0pZXXaGjM5fGqO3tg7dGhSokoPea1D0duceqlzomN8d1CnQy9Xwfh9CM85YguUWZqyaIqoDsgcOt
y9S+kDzEOEGaqkYESQuQbJBd7KIY26QVjm2jUNOWqyA34MgcuZU6DEFKgieEnoWh04wAmJUxIj9P
fkporYhTe6QlwLUpVAF3yv4dokRR63pe517/KV27L5h0Qhjypo/DLouYZGbX39L6mHqcUyUXdHE0
kV4hgUP+EAJOVIUChKJDO6fHBsbenahW+NAip9FLDZI4rwqZH5+uDcHs3r7Ac3CQT8uiJH8tDILU
X6DREs5XJXk/cTcXsClKM0JxQbaSLb+nxba9Axto32wbSUcWWKrIBAA7OjKm1ZB1jJiLDjt08VnY
AsTi/Blm/NkAZWrIlLuFhNn9rG6WwfL9vfdHjPDwMur9OToDDUFpgpe99cWs0BLCpxAfg3BGrgE8
9xcIQD3A9QSxSbaDAFo61dosYrpY6qEYKB6VX+rhxTcuYkZpcxvZfvsuEDymJoREKm39Bndwx7qs
6KlfwWG+Gag3bWzDq3pR+qVPZ0e3H96jlK34SPNiVyNE9bR2GDgbBYZJUVRaNN9qzEp7hhaFS/gw
YvdLG2QsS8yNYFq0EZohQFBz2mDPzG69p4aI2vckrjOtQO6k7lyRtFgXwxFKuH1IrUkNkh78Hutp
0BTG/YVw+C1/YN9kutYCy4D3bkGcVlWcx6GTRla1kXFk0GgK9EUy9aHn2/4wfRsCQemZf/weFc94
LeOA7dMDxwjiVHDr2j2GcaQ3AQGfXvcHEbFAwTzTWRDOBsfMLnKdY3y/gLlepD1LTTvnXXHCrWZA
i9618U0mtRi4ekMz3k+xJWDrQZd8wnzHoA2NCJYwzmdrbCxrZONUho4+4cOqGYFrzV/PMhOz2agt
dGXxdUn/EX4YVb4UH8Cr2HmnliWfB8NJY4G+6GVv0Qh0ZGSRvne2vKQb0xYoy4k6X/8+ZcB03/tz
bj3t2rHQxCKLSaCt1qDQu+Zp+pWHqwErpVVWX+HtGbzGNy2fJbR1dMM+fTkyDcC1AHg6QcHK9tBm
tjAgUZxXR4sBERuqkob7Xm/qXEPP+LdWotHPqIyqxa0K6pL2iKK1csvZh6EgRXrWgFNh/304ULhV
iyWdNzuQ4LiyJWfQyZotT0YHmFIzuq0NmbDB0Qi4V/L3/VIwBZ56sXXF19k2XToTQ/11b+/WMa0+
ELelhlMRT6L+yYfmjmXrxlEIupZu+vhmdjcAmu51Fo7Y4PpHmY5ouVPDEy4IfFdFDZrkofLCHntm
bXVeXY0wXfrIl9Pv+K/Ha4Pd9lVuVkoTGfarIOcJqsuehKg7cQnzGVhyS2tNhobZ6D7az7g5SkvZ
XmMtjfEp3jGN019oyEXP1IJ6dqBY7us+5KL6tuplTNaqYQwgMSQBnOQLGpkAJAFI+FUZQl3XfnCs
pMExa5wPFEIbpwpe5WXJXlI4cnTmhqj+j51doYYtHqt1OeKlJbiaO/3j9PUqOe+kVK5FNa6SiPea
IeSa6xhEEtXKsexp30dYQ3W0xwZtOJifD2lTkOp0PA6+9e9o8JG8UOaIomBzJLBIlNrhJfuAb56h
MUnFWW+3Llb6tVP0QzQYwSpeAdCETyA0s92a7tH7yp4fk1tF02L0AYz7eww6qZgQQ4rkqxvq6U1m
kbUA+rPOz83cl6yUkpvN5kzupjWjK43iqTl+r0r5dXGl6echaHS+s9oxg+W4FSn3qpmdKjpchg+h
idTy1fcDyaptaIpye/kyU35g7VY+X8bCjLiY08yEFTIhEsh0oS7XFHqNaAeT+THPoxoanutHLdUX
RWl5QZ6O0Vfg0AHeK2T2lMilM73ZeDyMgKG5eJY7RYHhJZD7Pkxmu7eqSjwq1eH8VdP0KKpqVcu1
GcQrYJiphPuUEDAkZTPhdoNXOMyMeE+xmMBLCKVYhrSP0SAJWG2e6LoOH2gM1WxmUdK0Rix9AyCL
fGP/9XpQp6lBnM/JhV+Z7PwlUeXOo9RS4sj9F01yH9kEAjUIZAqUFLqekePJq4N8lB6juwMILPoi
F6WicWrBw1eKFBDHy6cjjpykpV/t+ZkoLOLQ5aPW9Jvy329GyIowVVAUbi35F45p2tQyZckG2tex
hPDStkFoFJjnKt+HQA2fBJoIFQjdjS/xdUg/rRo2BO+6Kehbz/4vA3O5F2BnvFJ8hoCwlkGBYGO6
SP3pP/0hzTtLPGlMWmfmBgnPYV5GuwOyThXxupsrThe6nYltA/8QyNcyruq9hv+4iilaqqLJ/w4v
H4luUsHmdz6rOqxXSh5stWq3579OYnAbZNLGWBwswXxrlFzmZvFgG/ba/yMADmEQjSFWX3b/ZaS2
kjFrF0l4PWxJV172a0EiAULjdQwIy1w6q+D53Koudam0Ho5UEDDghdSgyX7YL8y0G7o4U51zux0g
WYGPorBWW1HX4eVemsVyE74eQyVSpP8vxmHOExKIj3hAQl25OaOyg9rjggH0smi/EQvgRcCv7kSO
Gf3w9SDROP3/BxyPf2vbX5hJwwdk+2raxTDWDO3kfceoOunOYZSCmZIrScdbq74+tktmibANjl3J
yWbHkoKFD07or0/bwc4nwDbVJRGOep+O88NzYAg/VzZTq0QlhS8278Cx57LO+PidNQOWbQPscxyT
GYXU9KoHxTPA2iDFoS52oYQyfU1kX2P/F/8/Vc3VnYOIKFrXxPR9tjnqXcAGYWjD4hVa2FxrnFBq
h5fGjjep0RAgxbY5V2Kspzhoc7sGJn/POilk/j9jP05udEio7NLvbIpJNK01Fr+WaShaIJfvxP85
h319qfAxZHP8gNDhTfOnsJ1O4x1xVoJYkmrTraZ7gXOdajlZqP06Zpwf/4O6cLwqxIzKSrPrkUJH
adUbBkE4L5+7yoRGQXnxzgzgscFZnMJxRz8eTskUQpbk0a7jAUr2lrpAqBznqQJNDX9rzScSezeg
DBeiejl96hgrewtylgLJwKlLnYbHx1hAWDeyVi5wsFUMnDb8FD+7IQI2irBIZhnyOuEwOOL1EROr
cH9PoLPrJycPNwEFgz6pV9kPU4ws0WJQeaWw5xOSRxmOpRbOfFbx+1RI0N+hICi9nt8k9degwaGf
8x+NptAZHLlMGfxf4+1ZxSaiIGN1pOy1/Whf1p/YHky3fQfiKO20ACYIO1xiuAEWMu8yVSmUWvlg
QRJptGp6A3VeJCNZAmt+NTz4UQWQ2GiF5Jt7DAzDUDCa4NE8N/lXbvkwLBtE13NVhMu7v8uKqVzv
IryyHo+A+3dPPdeR9LdBoaaXOUYe5BUeGE3FofUN4XnPvyu98iLThFO3UWzKHLVQrxRmGvtcl3xM
P+hl+tx6Ismu5Q7som2FOwe8UA80EluHnL7jDkCPzpdb6bMwnw/j6FDTzN1izMmPkhUeZDXeceX6
cuBu4XXnZphGEvamGrlaYkQYVOB0voCI4IJOCkYyU8eHpluiTsjI5M+twUTdrWsyQ9JYxzgbvSb/
ESpuf/H0rraevKZWWtC8dboPM8S5hZ+h9LFPr5Myw32F62TfDP4GJbiuG9B4XeLAICl8OfycfSrc
OqYGQt9BnsOSn0eEdrWDQDaNPP1+eR+Bu3GDoPbrg335gkWtZa5RRxGfnTrseau282Vrpe4xZrlZ
Oy4s4kO2ojO1OyZf6Hiqs7Xt+p7k/8/i/Eduj5VkqTvOxDdV8lO4XJVFPIMKkkci2TZq8uXyP3wk
BLr8LVA9N4LK3LE0WFImYzxvgOzcD0HYxDFngAXBQjMllTda6vMSm5S11VAvaQlaxyyGsxarEEYX
6W8j88RAQVwY8nvG3/ri9CYkYLoOG5BLoxlHJp0awHCrDswz07aGMxp0/LC0fH924ToMPgfrQ4bp
3IFLG2TzmvR60Vg6g/ogjnCv8oJm1sJz6tcyyU+y6i8oMgXiMqvCvII0lCWJeY7aMNv9MosfLqIU
zqDkX3ln6LpgZGmSQiOh4yIdtGCXWe9FdLEmJYp3RsAe5SP6EchrG/oz6knstBHpG0tQd/z0dWsy
71zjpgzLp1z7U3luf+sVMv4ypcU1+bdhf9fmdItP3QVQ9Lzhi89hukTBSVswxh/c7VpL9kk69yhY
rcdR0tuvC1WEJqSSU68StN24r4vk0m4ELjpEQ4RrPrNPZlNXz9XFRG+tpfLgr4u5ZXOBt1nB6t5o
SQUBtW0xeQjcW8OLagEHWLOr8aRZzrFSn717Eq5/X5iJg04R7zQiZyMHsjOrQ0vXGEkBjsF85nsp
l3xz/NpkFyHiOhMJVMXH30yVWVBFRK9khWPAo9hsVMrYHJsJm5ej8uC5OwjFy7lM9Fcu8hMyYS9J
siIHdW4LAGFXDgUpsEj+pqlfIxUMoR1iLjp62/wHvnFNKovJD0TEpwy7Vdy1HDkgdgKadI8nfwol
obVhw6xYAf8QJAMv1eROIe8U5SRMMqukMsipx1xy+eu9YdpZJTn6fTHkh7P5e0NF20pQ4qrpV97R
CeQDfgIM0Q8v9Uq+P6o22yT1vxdxPloAY6GI405jRNxfuA8Y3fhNM7gZz9RmgxbRzE/U2bJQwxtO
7VxVqPyzDAXcDhFQQtUStVpq0qtv9WRJkxNvvJtzIt7+wrTLr3dPpNoHQpCC238WE+czmuL8hiJY
Fcj1qzfp3flOTBPCXBwyk7KFXImhVJKxTxG404pb6wigS6O/w3YlmO7+ySZDWF+5gGtsM9c5CS8e
yYAX7BFt0QhKomhbb9PVEKlCoJ3OKGrN5XNu4Ki2a/88cxdwvz7G1T1Rm7tAekNdxdNZEqVSLpTw
e27z9RqIdj1oqSntrYChmg5o17mlXQDGGyKk92tTWNouR5HS44fQbYYiA+0WiaAVdy2D0nkgv8RY
DMyAQPOKQzTpyLOk1CM6POygWHI3bNbNRQpbpOpqO/jXphDTkWShIR+ACrM6mvznOOhWAt2jErWi
3zgQs+Mjpd8qTmBNoKtG7nxeD3gQCMThd64PG3ypHqt1I34cYWBVEFpDNp2YLP6ITwkS67keA3LO
d/dWQdEQuAAhadorj6m9RIDoyx95G0AttgLMYbRBFTvflhJ6Jl3fhiVPdu/zIulk12sXOnNeJe8v
UY5MJOB3el7JpT6X+j97IsU8r9K1SJmBDyhCIj7/zMk6tQ072sWR0IKd299XRM6vJk+ZmRnA9JDL
N5SHUD4WugETwLU/sJEMRbOXni9IoSlZUWfN6Re7DjUwTIFXV1Bve+JrwqB6/e5XQAz8wig92VDU
D9RKZGM99NomNY09nbSHkPfScMKY8DDNDrRUZEeEawQAIKYHt2us0ina6VQ8xDzHfQ8QwJuvR2yY
6lliH80nDNke+BleY3Au+Qodz/qDJ3pcJcCMWs22U/KdZOZiQFCsM/nXC8EK7/extq6vIuKuCe8a
wVoqfUCkf0RV5N2VlEUCL/Z41FyITvM5Y+B4/RA+xEWCecS6ODgPx+uQWDwb8Kf+jyHzldSILoKZ
H4aN99+27/Rr9SrTOCD3WA0JRsKED3sAL7725Dhb1WUVF8zw58qD7yCSt/0IgnCLujlIlBEyb9p9
/CdxAcdT6yaxr62Fl7WaNVmyGsM22pG4LjzxdrVPoIdIh9nQKPDRNb10Y3y69D5nXWzg5Ob7wOIA
raz95ydCEWKbIuEHTBCU4ViMYJT1Ks9UxZCWN9PBVyLuodZzSnsjE4466GED8xt/4s6B71BfKWtd
M2asmOeyEmmKYLHPFI+XRvijjT2Auk3gzN0ThojMpJuXAQ9AcS4VfasvCGe7InWxE7KlDzFwA9Rc
FnW8NwQmtEPlK9iyCLWIvvWfoQ7jBM5NSNnNCk6+F76YfsiC4TACxTrj1KQ/U4V+okz5huOrzWYM
EeLV3HRlS4yTO1/t7oXnhktvqGAGZg72mFtcBExHBHDx0HnmljdX+kaKO1qD1Xk5tQ5FJjRhSy5R
lbRs6uwMW2Hwojg2VEIp+90MjQZpNEr0uCmTwHJrJyZnP4i205cCtBmIi4nzwUiqVthVqFe4qSVv
LWB4qZcVO3e0/0zX3fpDe6jzkWMoWki3YEGZpyIO6t5rFP20LpP9NtMgmKRsxU1nDMHU6lfhhoD1
mN+RoR20D37mv+laqeTcThsNh+XkTPH1kEsLh3RX5quNyy2YeIzR7gyVYu31wvK9P44yA6xbvGnJ
tZV3gpuH9AZ6xiNBGCxHgxxtIPu3ajAUXKqF43mQed2H1kc58UMzF1u++KSz8GSVQDBluasucpYn
QRN/IfRImoJxLI7kh3sMZAp7/DSlQLpeEmc2qSPNVynrSrs0Bv3tM9T0Q8dMW9V+3m9HequaROX4
esCH5PTyiizioGQSut6nN074bmb7OGxGUkwzIYwl8KjgY/jlUDA8EjPK5knV1R2ySxL7/NlXlucb
TbBJlSNxQ9vz0sNUs28u+eWW27NC1zOiDHPqOSt5id7Em/tgmEP9/GtF+e5l5zo5aqh0j96u6F9F
jNq81eK4GMvGWs3iADSJf/XPSdgjQCEaQGWyGpRtw+Y6tBUNHqfQACCx6z1XPGMIe7hKfT0X5ppK
AzK9ztLogYBEAik19DXsfQud4WW8Flh4DT+mOMAkyLw1cbCnuNdqWCa/jW1o8EskNA1NR5azB+Gs
HcKlr43ZnwtCWbtBfGNgz+xQqxMif4o0THMmcaH2dE9a9IYyxhxhDpZa9K43DrivXyaXZBP698hY
D1OUNgkCWnx7c3OGuYq/LCTl8U7WV9mFLpANf+o3NNd6gckLQoB/Gxr4mUMqCIecXn7Ui3/pm0Kr
c4a6vw0wZ/TKNVyJhVXgwesIJ+BVZSIsvo0fnpK1PoIWZpIPn2wWMxXgrJAaKFgFMXy1bkZhGyzD
80amN9j/JHj+ZBNM4Y5CNWaPKe1AxaU2PmzgXMVrISRR/3uCfI+D2uxesar135o4vGJgYv/NjVNY
F0dxP5ueWHrcCEBHfA2v7HLww+RViBoT+Xlr3kqDDipptkh243tkXC3FPw6A8b8TkDQAcmSfdiDJ
X4jjFlhZezRQ4jRRbboWfhylyjJAwYVOrUdC595izanG9QWdsG/qaRiKwgiIUjhigJfomCFb/OzR
puJHqBG40uCxtzFkC3FMv8PSw1SkRQnm6fignk6SLw/dsDfZEuLA/HeMDRQWvKDarx87VI/T0nNl
vcrkKryck0yQQaNwUfebcJf1MI2ghGlOdUkCJyac0UWqRIK+40EOIqMdA9QbdmlbOsxRX9RGLxn2
iqrxZZEkZfKQ/JZpfxeIN05ZU1YNZZEKuDyw8MnJN2d/nwUUfRpdkzT27HAMX0F7maHTu1nVXK51
E7hgkw+o8t5BOtpk7XzraqeE7W87pdR7gkDVS5HtpjyFACfIsPJZOgEKtPkVO3fgVoikhoI8kWaK
HgvXfguc58L9kqi3jIqZ3qE4MCHaNh/LOojAjVPJhH5tIkSRe1JdYs5C9ZPk+MDYL8//bGKUTkg5
P9cvxorNzbUXbltSabn36mwvmmGGTwmFoZPJzfNAChQAXyZnmx9l4AlNGmso5n4CQY91ToyKcsb6
+fhTz/eTVpblUnnUVMfbAcSXaa+6AQac5OhIPZYNp8ylDtuPEJA2IBcJUoQBldNcC55IWQJghB2J
Yw8QWN7zs3lf7O30PA/iW5Y7ewaC0bEITNoGJ+8WLxqNaisLybX/EI5B9iLk0bAdTMVcRPFlrZz2
wFYjmfynGqPXI4tTDjFqHs5Dc3EhBZPH7nc/vAMC4JpGuHETi4fRL0GNDPwZAadWDnuj6LaERjR3
ajMQrp+QDvXB0OzmIHnVdxvjBk96Mv1RYmIn7XUsmy4glDGSr4tuaPcf7XDiYREvyQRqvddAXTW8
U45rHePALhNP0CsG6evUP0cJEbooNxKoKm9lg7a4EGtrbCEZJia3woA0g+AfLSvvOgkOoDf2LyZS
u6PZndiIufJmn2vZE9RAG1iRSsDA7rN/4+NSI+NO01WWV8ZZjTUItVapr8uUaC8N7zqscKEf63+O
RdTLPqKyPWe6XYjkyaL1rsrXjHq67NMTNEWrtLjNCnXX0Nwvpi16lbo988MblW+ngO6AQPsHgAUJ
GRezUSg3xFX2qMcp4Wg2NVASm0+9HxI1J9Q82VuqF+RaCYksmMGhWk2KM957SIveMZRDB15ApQLW
9QyRZ+fpnq3qdhIZpggfQBaQqnVy3dqCqEAM8JsYWJZ/mZU4J1fqU6ZDEPLG6kcA68+1Hjc/2mLZ
j+0myTRS62cKlWUlW4Rcs8E9YJL5OIhb8rOjOI6yL7TWsSqWgnPPfGZdyT0o87C9jpl1StFx4lMO
8n3XBT33tqBwznGPTLRtVlcIVZP7vBFstq2tOidU1sdKXPEEKLeDaC9cVly+hEMBIPBePGS3lkGP
FXvdb1PBevNkxylbuYKM82PTFUJY3Yqc4Mwp5r/77shzFnIGg9+8wDsQXPGEj4oaHhkDnakmL1tC
zXA22mVJCVC5JwkNTLZt+SAIFXcG0hGKgvcX4+JZZ6QoNCHFxyjZb34pdz/TEgpFCHxs0YBXeUGH
kPailUZmEuWhOUKtRceGSBxakATFTd8dkkmnai1N/FLuu3rsUXnHNJ1p+sePdXsLO7N4Ol8RtKbQ
HmPYvY1s15ZpJQulzG0w14VENhJdueGX+gwMUDrF1r8Ufjzznpcai1GzHIjrSrjQekPsOZzsat4m
OIsqs96P3gWAM5GzBosZOj79zFuWL8BN/zLpHKuK0b+XkxmA8ka9DH/pHVrROSyCpW+WMSc3Q8U4
TIYwJFHjrPd3f4ppmSIB9ks/Mj5SyCGkW3/wbc8pCLFAd5WdI51leCvhRCWI7aEtf6Gz+UpW5x4t
/VI5NU2/NV8QjLk36rvO7J2alCIKowvaNqIUT1nsHorLUFl2T3oPzw0FxxyGNtmTvWa1/ZGlLYK+
Gt44vC9UZwnw/ZUGMAC/ZGIdI8ic/NqDfvs0D2sM4RoFnfpER7MH57Z9Ryb3VUI/Qt0m2tletI12
EiytZGZzLqtm1bI7CV3s8Ds25AJdeMEW1aLIk6FeEre6IHGIPgq+4+7fQLEaOsGoB1hwL4FmWqm6
yvexfYHjpjTr4En71sgllr3dqmmrYvKIsuKBZWn4fZtxYVHB6USBUpchHSjd9PBXhJdYhmQSZdFv
P6wZlQZyNeKJHv7LKmSIVSFyFvXMHGN6RJcwQ2EMQ3tPb1fHdNrzEhsgnWVA5aKrav7ac131o7PC
ivLNHoBeGRosW/8Xa9URZiX+vc+EzZSJCcxkjY8itkI5co0VDLQMD11zIxOsusgoFM+ZCkMMCZUb
UnvJdeIl7V8g0z8iS/tU/WyJdxGxL4A38d03DRXW8T+ovTqSH7JiXejr7rnaGcSAQknJMwUv+xK7
n9BIU+wEgTZSN1Xs36s3j5qUZCfw7bCI9cYhRlQES1/JbhhSI4vmZHLPjzZE52oxe+83v/Ur1ShN
ZL0z+/jZprgGEp2hS2H8tL79ZS+WbQr2jGVfVuFP6aATdoeNtDIOj6rVLA6eRrxGItn98E5mY54u
ejgamyrDKkRCXyNuiLOmv8vMPxqFxGldlY5sXf34Ql9cPFecqHD1CmO0s8Tn+S+jlpX5fSOiBnKY
i5fo9J2k0d+1e4UK7Er4I7ZmdcW7a19kfiNd7lsLCzllVfATkNROAl6lfmRRunQbXnMIdQVLq4Oz
FjqJDczEtVkm6yYaODyDQmqGcv1OGXz4hGQLpRzhxMCjBtcRXEYsvhhBv79vqPGu3ruEh81Ii5m1
lGIGOCmEc7w2qu4vt22F5MCnNYS+4MEH6B5iKU2+2WF0M1YLe3HvQHOTc9bTB/2UMR9XUj9Dpbze
+/Bga6UUiW9MmQcbuVZykIvr/AoMTceY2bNy/J+U3tu+rB4SLq+6kpxJzTfUCyOdIG6Tv26t7mer
jf7MsspFzre4zXe4VHCfBarZcCDrE+/RWRWO+/BHg3hzD6NDnSiQEVghncrhQbsA2spqGsbQhnFS
woeDrpixKVfTIyfTX46/3/qOe1tvPBBSy0axmr+QlloxjZvlRy9PIVqHRx262JkSAawmN9P9w3ri
W/0JcOLWddvWkgJY8R/i4LDhJqvG8+zo4BLP247J/cTNND7aAPoPdNvok1Vy94J+KSwI3W5AzqCX
yVVjcjNwL9q3LZQC0etIFauto+Z+WhDy052zDZ/DCjZIrsi7zUZOOya0moZocNesfy28j9v3ybL+
+cHYJp0mQ4fbwcFbYJoJZLEmfoSBIQEthMC4D0sG1E8iWgJkLKIqkIYpdVCjDugB8b0x3YpU/Rq+
zru2IdHqQ2LtyJ/knsk04nfwOiHwGkm6zqJZPIFifEWZkoNuVR0LRnKN4F9xmToOCyL3/jatFUJI
dYzFlvDivKEgeBESpVsDzA0BSFgOkaDPOB7wpAl7zjEbJYrlhz3j6vdZPwR3i6/IPkgU8+zKr3IS
GDos/XNjLRE8LBdWfyloieEhp+sLy54b4H9Z4sBdtzNVovl7JG+v4VE468LQZxLCQCXBtrcpN+rH
Il9FzzZ3yppwmy3PRFAcwFeBaSV9WE+fYbCcPjomuQPVNuXjqnGZ3RfY0QOHIxd6wspbFhsJmmb9
ZEpF/mqIIwhJ5RdImgGmsVmDH/fHPrVkkuB68W3zRJPKj9sO6PpK4COyp2bicV9pFJ+ycVzgF1Z5
Pn+fVXO4LchCf3Ur9Wt4vf32GnGbhjbXBpCYIKLINL0Gz58Pg72hgomHaKLdzVh/0/iiM8cbWyKR
whugAVb8li3kgMOPqvPDzDUjWjWfu5I1ZogVT5RWAPFoAqvK0BCOQnNrsQG6sCGx/4pG2uCCJH3b
S+MIaI5b2akQrZsGY7kHB1nsgntuvzVprniuH1gfudhzd8v+oyqFHA5eTP9zOHR/Dp4I3AEx0XM4
8mHmUtLc0LiHSjweWnw+V2Bam89aCmSoArrE5BdXAdRfdSBWsxHM0DIkIr6UYpRIKhIN+d64Firt
I688z0PafQZtXRZWSRuIbWuFYdils/jWMTlfsu8w1C+WTG1njUJBaLNPNHI5KMvqhwFMmIdMXPEk
qyYK05ThaQp+ThhDoN5O7yshkMlVTQs31C3nMIXU+mXuoOeXIkhuXZIswLfGMaEpEW8Om4dh2Of6
bNIsf+wdOW6bRkXDSk7K62UodaJkgie8giLmauQPrBpF2llTSI4nxnhF8L8kQFao47BQwGsKnlCs
dzw64p46J9P02mJYBfxj7DSiL835AQG/WemBkHE3TVT8wmX0m68uQWH91OfNmEvHg55MhmVcPTLr
/L+Zf95QzaYzxZ+7CHDEyrXgCmlsVKKX8NLBxjXjf4hBXDwGLlAVCybE1Ul7HueaSZh9ZAEYPoDf
/eNKGWzVU23jQPRHOOt50iJb/0I71YWKzljLx+8qgV+Zrc8OArEC++VPx7ecssK3VTCGjMcninN8
58Cl82RKmELWQlWGDzksrIqzUKP7ytpRIZK8p9czqvNMYENfNukjHLnMi4GtwGWeOG8blaiHSOI2
B4XQsimt/Bff4prARsvT0C4v5zqsZmox7epg4zGciQM2h1RYO/hK7MiYaQ36+XDJx8jjEaRjCUt4
0iZFXZGDdsWaE2Wr5Ua2gQNNH8cz0zgaKxvNMR38gKzvuemd6NOwoxTcZ7JELxx93cYFxkYgePSx
CYkPxDqweUHzamMYZ1yzIlvnIAeO0uwu1jB4oWsi/72Sn2h9zkVcnH6A90R+je9Ptctl6BpMDIXy
vS07f4PLcbE/HvFsXYLgyM8J3YUHd149/V5+IFpmj6DpRYSEQEMEM82TTIhRmZtyfgbN1ubQIbCs
6gzpnmvvKt0/O3KAtyU91xs0o2LNMtpl5ZdwejGR9sDNmamWPV1Zu3f/pNR9AsOckIYhqprTvBT5
D2/wJIHWknZ4L1zFyKlcuwRVbHmoGLmXXgNuTY6fGimkAPpEIpWmR6RvuKvgMIhb/u2s3S67TeM6
RDVr0tzWuZzjGBcH8zIldQzIuAnjTWJBbRoWN7NtvlkMIAXdtgO1eggupomHs+GkZCU/IvpzRvQW
DAA1IOPMmXUZ7c95CA3Xqcf3K46iQVVvCg9HliwVENW9nR0L279J8ODa275BLSLTZSP9h5putizR
TScRuTnle+6apN8Ct+bj9z7CjplcDoR6tUJfZ6Pa1w1KPXRwpHEmQfHqHI4s9ojarb2pZZ2gw510
88VQRztNgHVGnwgODAveC5ozNXCrOyvCyBg+N7YOpgvNn+/H9uJ1W7IZVcfmAL0OHlZx/oWhJ/rX
0RRsZNOZUEuLsQzh2hU6F5qglFD9vZB/pLzs7ZmkiWzNQhfJ6+FDixBiksgbEPcHQ4lBgKneY3bj
8IX3mvKTk2D/wXh6wuX01BuzdWWSYP3OTk8HBurJEfuTJV1xdZHUASUjfw2yUEnbTGUtECArzCUQ
6zThcxeqsA6mrM7XbV6P+4+fs6gBaEtsQmMSTRVE1aBpmaeC4XpvOpJnbi1GvW9O6aUlYPEr/PYw
GGPZRrbMgSM6qd+DtD6NZ6wYCq11+DMr/wUK1nPOD27oz5j9a4Vybd7t9GXMshqSzUoCTGxcXHaa
rilA0/6T6Re604twAphzpguYauT/D/c9Kmi9MwJtErjmC9RSgl69pqH+vQLdQF1tWmqObzBbyGNg
H+bg7YOYUjzK+03xYLbcmXyfnoIn4UoaZfJLckcRMcXcu2nX/qJ1gnXzNZ9mL5c6Ye4aRTHaHmz4
R5zXI0b2z2Qa8uEk/WK6Rx3Kgocnb1OXgABajeYr/SzLSlmfC2QY+6+Bf+jLLNXQpN7TIwmK3xMI
dMATiEsH/IzzRRxp8yquNnlag98NaWXh21bu1lg9oz3+HZKzrULBwhQPMU6BdWFQ2i3zqdQvZiQH
eK/utjv8Smswc+74Q36DpG5RNDEL2YkA8N0d09ctd7FatYiLSdcoevSnQY1QOYteF2tkxJET8SkI
DIQYC/gpYCBR9sEUshfymGath+sdhdGW1Y+fjO5WKDqRF9wZuYiKc5NlA2dJL4ZF5ZA7jsPZNEwH
iZfneImgpjIqxgs86Ccltx2gmV+1BeCnHB8xrrSvkM0HcH2aCCMLDL2S4/Oe2rItG0N86bSLB7xd
H075JFYLUx2liv3BnLBIzROMS4qmADfuhOUD2wNWEtKyrEV0n4RPsvtCQAvGi95trsUhaUC8EN03
NWlivQnoCPt7RJK7UpGUAhNK9AgFhy/6yxiiBZgHhoJkWK/CNhSyxS6UERT9hr0TOVWLtQue9VKQ
qRR23EmLF8vZ6N50Q5o5kpxg40H9L8qIaAxKEQ/QT1qSTkir1hds4+vEKA+EgAzf2rkvU0RvZEuP
rs9LOHhVCcxk3VF5080dbvbpZppa3n4k+9z+xdt5QJE0tNDnqcGhJD+2eA6SjyE/YfQzkms57LIE
FM4SSrKfaS5E0biZ9oNKPPdu4W/4Kv6NqWoHW4bSFY8SWAaPDPeJ9eb4kwmDBsS6amRuuylH8PVW
jcUKtmr3A9RXNcyfXGM2D+C4wJ2AlD2ioVpL29P6cmEA1YsXxVo7AcGZFH26e3MFqZxxjek65NGW
CsubQAnoFta3hVy4tdoG1WKivlIx/GqFQDOfex26Up/MtuMKUNJHZK6YUqNgN4lv3GZYIELoaz6u
oKho6nLGbU+FcCXjZReYJHXS6Oh8fu50pavNrUo2VygkLMP8oBQZ/5E/3o1KhPnBeEjm+f3B8LKI
4FhTDHctGlNNHl2Fn0YKy9W9gYI0H+GW2YRSuUCT1PfbWmhQsEzNQF+LVm3XbLufmQbUvuvtrcZX
UjBtxz12/UpCulaptGQCdfh91qjaCTR45C4jXKccBxJmONzkc8JCPEmAO83L5DuzWPSowq2s/b/7
F7vVrqXDB40BoAz+VNsXLmAwsuJHTnbz1bkN5YtA+OHbwrh3VPk9Atce7WSJ/iGXrU6mWw2O5FnH
xLrIHbDY1u4Agh2YrEnRnpj/J9P3DbaQgFnPn/4o8sxQ9UOWS9LwFOKj0jLrXjZnfHsfvquISmjc
RyjcPtMA9p2IUmR7cXCRqzyCbuyAhzgMpXR86n1a3rMKJcifVraGIbC/Mji99FGozGVWqJN9NzBl
zKSO7Ny3QMpmPtpdwkD5jpjNg3ecvPZzcJi1me+czlptb9GhSKpLMKvWpaB+N0V8Ws/KXKfRkyKy
xZiJWf7hUIegaK8Qc6kxb1fQqoASZ/q1S7jn1Gu6m5tL+y0Iw3iFVGF99DmDfMvyDCXHTi2F1GuD
HCtzzojD9NUDLrLyx1/Ah/+vTUsaep0Grl560Y46egPmL8+OLjpex6rLK/lhGWfcl/PRwKmMax08
NCPe/J7q+eyyne2NX40dZg+GPCV2sKDpTd1akXZqTdmKYYnDTW1SMGF2mPiyXfvdtyYCacNaFDcx
87i3L5rtpv+f2HSpIVZiLqQauZIBdMA0kTnHrGpbhY5oO9xdzz0t1IYGkE9UXtWs++aC2yYkOHEw
MqklQtKCJdn6SpEzgyC87TwepLKC9eprS2UIINNsO95/8pbouJuuq3ISKh/0rs/4DbnwyG3BGpmM
7sfhQdb0El1SYHRSdL0wkw85KgYk/Md5zxwFVsjCszNpUzY3HwKuT9JqTWIi83JLJGbOGYrETRje
58RA0R+hAn4epAnD/aTmonIUUAApCA4gSXLNw9p3sHtM6P8w/SETSJiYLNYJGUmOZv8626o6ibJ9
E/O3BCJuqKIt2r39qVaLILenqqscg49N/qKzp2HV6jG1zslO0OOe2Ux/aAMH05Hjh00p2dw0MGbv
/sC9tVJD/S+uLdLDf2d+5s9C0FFGncERulNOGzrkrTLuP0BSF5MsE/zuZFd9qmAclaoI8umXO4Hw
gZWOo5G6Bx8DNENHl2aMTj5IWkz6CkPLkTUgnUAuop7i6BfGaE9KosktQMMOtGeT12Bzg7XfbbDB
mxjhVZB7vOcpXUpq3Q9BJu3AusgWCsOBVQL4648jq/fmbYrRDaITC9SkeGF+FHuj+rz2DwUltudj
UFy3XhXQOmrpfNBiZtE52ZHl8NYir0CHVTEMurlNP95g3oHvJEx0Q4ZE4hjG6oIYsgXIyQVpnxc2
wuKiCzMv3UAKrxI/YrELbYWkadFNeZxR1mCyqBsfSs8ZEdqSdJAYezug2XssaUfNu044+ezk6Sf8
eWGo2ceS8gYwLswPbqIQ1u2Vn4xm/gFVq7uxfesVEbJuFTlkUVpXUfavmuPf7AzLgs+cOvNLWtuz
lIPN5PtVWZEk1+YU0gU3+pMRzLD38l2gMnKH6WoTNVZA1iDjJ6Z5ZoHCsRxKF6gYoR6WRSdU61P0
c7ObiyS5QXBf9sKHuisODAvKTwIa3mb7VYac0+1LaY+8mSSYL8PyHQnmtJmPuNNRT34p8uf3uZNN
QCaqaQG4LpaB75GWJXAEGmaK4ymrrZRMDe6fTrnaO17a3vYGKjx9Wma1DxZcPO/GpeJVr5E5QnG8
CDM7BzO+ZHfqmJxYiIn6LW7NxK4aEX0icpnRrfIH2EA8RmS4Day+47N/aobyt/6h2KppPn6BRSR9
ugmd99eMklq7UpiclO3BG8aGBAcOmvJmW7/dKP7lHKCZX8TaINCO1h+66z7jcgsRmqERyZRTBjPc
U2KrgyJvTDf0tJpVzsGCDloL08z53zsCCbnCLkM4NCdgyZFBd27ogNclyuW950qCE4IxKbrY5486
IRh0XHLSdOXgCHBbOI1GKKOknLBLhppOEZvatPuSFVv6ShqN0uM3ewOAwrXCuKgkiKAn4/5lEepk
HTYvHjt9ME9QLlv5sT2tRDxvNfxOxsNM509qAUhYZPfhYEH96Sz836YHzIFyJ/FWpQTNXlaD5ULV
WrPK5Gv06RBfHr/uY7eBa/OSNEtKrxE0K+4b1S2glNZWEnnuR+6Bxu+NzvHtEc2jq0WAqtJoTk9M
VbvH46totbZQwAFtc3eTZa4E1Blj0E10Gd0cpx92nrAQZ+CLeuqxdSbqbuAdhGWIpbNW/mhLX3/6
ASmxIYuoiNiiFeoz9tYaFOyVMZpxgBC6+4KBfqEthl91RNOgK1XIGTLrqkj5me2UH7411Le6lScR
gZsUAMxHkCCVtKihM7lvaDTyyebvbde1Yai1WQ50GxXvtPgQmtxx2wKF+JJvrKC4kcTulTG0jevZ
5YoicQ6DJsKGyoUZbT7ZgB2G5pnSYOSFXwdUg3UFNTuMD1rWGIlC+EK/INhfhKlVPdPligEEiLfa
EUNGjmU6yVZDL+AzdHcsxIhDr/1bOhN9q8DI9lkdLcP3Aj2D/KTOhjePtxd3S3B+3oFPPlcH/D7E
unsuqtBy1rLImJGWdZJy8l8VgquSF4CKRQsTMqkiUrGOelsb0eV2MJBBXY5JXU9Za0iTfhXYEAlm
vsx00NayCmeRfSnTkrfH4NFoMamMphenoCMLl/BCJGtHvRTUImN8edf9q5R8LKkRk7YhJf2LuJz7
sNsn/aVFr9wrRBTtKaxpOdHqbKBhD802yrrXE/oB21p6dC+W7CO2N8FB3kTPRw4dk60+iIqxCMS0
SEIU2uSH4oFI9QiEa0CysaV92v5wQS0Y6tfeXP1/I1wu9smWK061gLS0CyEr/h5ZbftT/l/+GUnf
P9TA2JrPP+B2bwA3isoA4XQlhdYFuDjKpYR8JMGhcbZubPL4eP53Bpf7lhKq7grDxZPi4in6KA2S
7G16UaYwZoxn420MT26qCvlVogk0kQ1aEVVBSPihlyh03VSLDY1oMTvYAuzxa64LgWfjrnv7y/yt
GgcS/Jseb60Z1R06qy8Y/1KRA7Ojk6kbNRsJhw0c3Vt2VxBnq1pZaP1PlsDmrhMgW+v6d8uAgn4k
EH/a6GtVjadFR/TbbHzbl/S+1t2r9KNDScLeZXhFX1IknB+UnuproNs1TBekXvsX+8UFRV/QqfyF
ImpBYjNHd3QCQZ5lP6K6dfYvTrxGnForeq2s9+1je/uCHIHOFudw7eNu+DEbVDVf32xEiMg9QQaD
VWqm/1ucMEOU2NVD3ZVMPGGODlxQzQ40LGbFE/roqcWacsCEYQzFN3lYv96OhL17Jh86niYCdJ7w
1G8UK3s2nMj3uM3lquKyHvGI/+vVhwJD4MIL2gOanC+aktvm1rTPmsJe+Z8QLy8o06/8iY20Hu6/
AFtSCgf8gLJNrXHGZmxPuCYPKfqZAEY5BOLa6HxJH6OFAYQFJMWNJO61jgeXQ/BB4u4PGsl8CIYP
eErpXFuEvlDwZ1npmWJE0upH0wUV5EtKm/JKfdRvbHhoe3S7WPhfkMZQsfNxGxaljt4fHywENXRR
UOVAyG19A2ib8gARRyJW1dmNfr2WyMDBVvlDKOnmXbFWAf5/jSzAWJ0SYae6Uuj5OIh9dVxO37mr
ElF4Fe3eBzwg6+Sn+oKj9vRkVk8Urp1oOlN7HkY8hN191I80iwr/B3TsBTq4TuQGNcQdyaxE0zPc
GDieslVi1iqukgudFnKtD/Fa5FiEv68m3ZW1PGEtReTvQ/ZIsZ9PU47Wu8dBj8r6irHnXNCuysRf
WZO5QEqT5r2feD7O7+es8MR9SEkokCqohGn+Q9s2kUN0KmTUjowbmHshc8fEdRW//b3ijUxJGJbb
B8aUDd2LfmmJoT40bs1BybNX5CYKMFDviJgM5KchjFJlLJSJRbI3B0scuFbqQWRDyx0LHuU/YZRo
egDNHYR9o4laCsa6gLglrUPr5nHFkKgE0Feih2+gqG0XnUIlRC2lSIISmbySaR9ozpyrCilxd1v0
2E/Y6Fldq3gLTiFiyyEULARG3AzIA+4/c2owXAcU65g6fBwvksL8/LcrrfSpxywrj7b9sanyQTr4
SFAR1puJJp5Z2XKP4USrA0aGR7MHqR+EeaGLjXYfc0erNT+n13/t/hzV/kJA5XDx9I8Nz7HkHoIP
z13hKmiupuYsCtn5MjSIuP4UOrNIcxSotHwKwFzE1pM7xczlmF49/0dGEouYmNyJGqEl2cCS1NAx
0e9ZGp9tJknKJGZkwewNLyATmuIVVwSJnIjseV5h06Din5XBhfW0uufVPz5sEWhssg1vs7HWM6TG
/yDpGHbXHnZyGwNRHFItYIG5aJ2nBuHU7I3t1kOV0MOhhWP5QUt9DOXCLHI5hWw18kelugTW/R/M
jlQBC7hAIh8jeIy3eCtj50FchZtfWvKPjvLrrXbThdP+BbEVNUFmSsr4scGDALYXhLcNtj9FHjTP
FGCQ1a+KWlY7+DPFNk1oXfwT6LnKGyiYsGIMYzqgdn/y/LznV5DCoUborcNzlwSx3mI0rMTn4rF1
qWBeJ/y9fV6375ouubKnqu5VGRzebVvfoxZsdO8jODD0sIBRCxltPWpFPpm4KI2W7R38/gzcAysP
VNC4br6pKUSuZyWWwY46V4XBqXnej6be/LRQqgU+eTdJv/3g1veluC/oQ0+jnN6QoEVf5GR7YHYG
430wZ2CqksCXzFpA8xEwwiLsjyhPMtHj08Xih/yrE7eJYCFhRWVijxMNzQ1kN2A2B+DN7S17W4RS
miUrpM1XWfz4oCaumRbHt475xRqFDL43WYBUfqDcTms+94SIb4WBaHEfW5DXDvAFHLisqM1qPRUW
X65aWK0KSMBA3UaGs+qlnKY2NnjA204AywYsMyD2uCIZTeXw6sDLkWKAhPVyio3cECx4PAJsfZMv
ybZD3NDIjy56RNNBIpmS/N2SJE10UhMHGqTFGgvPpvXbPjMaEQ5Y7h1oqnXJYPz2HuDk7qFWhliJ
pfUCwDVs9c00IpQY7F1SLK3rpfnPBSZcef7BWPlgXqi/phI9UEx0n7BAECnB6H7CidNysWYsT0n+
+O4JZrnvcTDoXfWmtBWzrRkPNx79t2uXX9Akr81IzZYmPJdUcwSHZ+GzyI+XHFrj2lnAirCq0rXz
7ly+EFPNYYuiBOHR0cvtTI0e37wOHRygJFXYo6lj+UVk/5ElpnA+B+GiqNwq2GPhWjRZBy5yyzS2
A0eiORhcA78gexyzPA+777VHAXHxF1lnniied9ZcSBdwrs2t52RPv01vZ83crbRB9JtnPkQecose
APsosYe04Dga3P3Whrm1vMCIIJvW7d4PVCPfIuTStd9eMIKytKi16esYCe/P9smKUu+JAOI8p4Vp
w8N0YmDJEoPG1HUdeKrJ1IfzuTsHDHiUbetrCRPLzqf5toXUjGZn00sVIorl0Kwr7W4l57FF4ks/
9fI7GopD1GqaXsmgEc61C1tqlymcPQlFidsW9KCs2UXKImdrTbuTzhppjkh3+5Ry1RdR9EXfVyxh
t3chcBEv+NNlTn4yJOtcccwh+7NqIJVCAnx3GNSQNdF8ndSCEA3rfsi9h/Bqx4soElYame1H0ek7
O8LME35e/SLtkx0ScODY3q5CAtAf1tVqy6AXzuTPu/hOLucc0eeN0JDYfbAaN/NOsBwg4RCSIEvD
dQy1nzNW9UY2W0cDhztUZTVtt4iFsQQ+yIbfWkTkYLOvzdXBAOVb3mwO+eWxeCY++ZKj0ZfhObhK
MHAFsMtWYU+VijqoxSOeGd+4v5dXgpMNYZ7Wc/uqxwxdCzznxovEz1h5OIcqz9jWGOjx3JLVxKyc
C7ICFWzOV2cRNECUzHNH9oNCspWsfsH91icQKx3ovTA4zXQ1T1BSQejmoXOuqkKo8uqrBYho9PqT
+pSxKwmMZdZkRgyhdFCGFqT9PaH6g9S/7YYlKN4mD75FH6VgWmpZ6JeUrYR6KTRqMh8PjF6PtRNq
PRGlKM7pA1WofWKTvosRRWzHV2d+aaHBTnwtJVv6gs/7+2IJpl5K+LO0hMDfMtLSliDhfwEhyMrt
jnfU6n9nrYGHUp6mObkhofaO2src7zoUXePUO/clnfJrtoDeu21zzb8zO4RMeaLJSqTY9vsxVKsF
Eb9hA6n8F377M+P9hHbq4l/VNrsB+IgcXaTMwB9q9qbDCWLXkJWEEyxIXlQz6daSBQTbBxyCozBj
pZi9DcEHeDUijnbEPIGKjoRRRDRyXAoGHUWsH49A7dKk97TJhFNBMM22o7lJgYSxL03jKjuia4oK
TtRrtSiZrQoboElTJxSyU7urCcw61uQqCQcVTGuhc4MYboGB8aT8ITAZ76n5V1rdcVvVTA63gE5B
NMEBnyjt5eBOdDKvSBpPhgUWWyC/FBb2UUW5lAYgI2pN+VglOIwxFORD0kNIbfJsGpYfjlJc6nyR
P3DIrwvsAgVKUlCY99M23g/zVuLWciVbnnYjAE7BqWo8XjCte3SrpgWiwgp/7pB81el26pXOWO0A
29459kFduJ+kUl+GA9jWI9uSJAmT5ZLvWBD58d8pD+pyUasVp21KlLKrk7mmfYKNhdr6v58H4gfH
bxKhXyO+0IyNLobBFHFvbMHyVWOVG8VTUP6tdaAKV+3K3VzGoemrGpCG1o/jI3Bek6EBr4+XzcjJ
TwnYAWsp9qsUER9yHhkJ6miaa/6LocFIWAsJvOt2N/XhP3Dp1vpNnW5XqPlCzABgSZjtIevaTUlv
YVGRPgq+n/VpkQCdg8XIGG85PrflBWvaQtwU1qvPNyagFrB2EwYGHaEQj1ibuABWkkz0iFuT7ZjI
9bn7N5Ee3043BlmGzLpNUZYbKXQvFHgYpuXNtSOCRwr1OGy9qjZklwufnegXI5+OdqocuQaWaiJt
WqMu2ayMcbLyzOqOR1QCCooJv8Sbi5vK/sDDF/jSm7gIAUzeVjc2ticpEEtzPE80NoNvbgp8UWk7
BGwmrP4whk/zB7PJ5TW3XNV7hqOijCGgZWWRMtbzsYDWVj+JSRkqkSigd/rX+Fc6IFmpCZ2TGTXz
+Br/tL6QfIke35tMCD9ctds+QwJnmcNvDe8kIWxR5+w1KVLFSFcYk/818cMEuoSTWOeccaNswNIS
4aHQdyCQ0n9hKKXZln9lelo8Bj2jSXvyhKJq+sHy0PrHggrIfHpSpc4xkXzOQMURSPNUrYsS29MG
MDJSa3SAO8Me23eeF2qAwZ0BnT+0A2xrGU4yvv/mu8SI358tLuqSUTzKQnPd2dbMjDrOuvuAnBcK
J1OY7r9saQxVYEQXpOek4yB229fuBVtOCPFv1i8i8FQ6W8xoLVNyr/pketmNIvUd8s+Ud4Cm+6uQ
IeXmK0xbT7QyXPlmCDoMWwVQb2X1/XbPN2lP2P4/xhxTcnwXRfkvqVuST/1cY8xJLFNq4iqbxhDf
6y0AKvdxQVoXsU+cYLVEC9sZHzf1hlTlEYyzuPQNenzvMx8K9eZZt4Ohd5lIQAOKkWpO57zGoBv+
2C+bSWjIR7Sqc8pKhzuCRSQLtNBsAc3HPz6OsUiE7IG8z0yswnZeUzxSzhDUHAucwVcCgcK4p4SJ
tbo1Sszen82hTfbdnXgJOXZ+VR5d2hKLA0VnOg+186lO8D24So2Z4SHDZQgMlBYJTudlVKBVKH7y
P0Ac6xSsWC1hSuDoNfJ/SzAplR9l79V46Bv/bMCPPgVJP7KQMQ0ljQZEhRKkR2deOhcmPV/2cVjx
518W9BCo+dusbevP63BP+w0Av5JWD2rQyxg8Zq5XIM+IoEuhqmLZJF97uSti7ZcwxKOSR/1CkD+2
kgrwPtCFFG/eBxB59zpxmHB6JsXnCzT8NztRoPcrFUFSRuDgtLtPxkOnGZKe0SyJ0XshGkKc5fTN
3grEwhXAfhgfZIeHexDeASyiaH9v2mpjPtPsg5zxyHCjzt5fLDc0Up3BApTfTeBqmFV+ms7gtWtj
enRgSaxlXpIHz9f/rbze0R/5Ax6yaP4L6l7zH/Vw4HotOdHYBkOq9SofEL7jisg9+CYwRSEmuslb
ChxRlM+N4ZJUqIv739DNMT3Gl7BIroPAFu/mRpj+5f76UpqZdNxFTCSv9xDAaSyd/d/cFTzbIzgY
DxCGDQbNIV2q9yWHiZ7ZgK+yvJIeMIBdM5xxGyzHe9DKR81mKopqMaC+zl/XiuGPTaml7U/CXrJJ
jZtumQPAbc/aqtHPhb21MeLz1nuV/Zwv9TvOBtL9tGVVvq/OJ4ArhNl826SqUVcoEPLMqwFDwWid
Tf8fanH4cTCCc9b3uPIAzugkWXZqGlH0vGkqmr2E7OBT21c949kNWhPY6Xu0mm6fOrTyDQR2/lPv
3HZWnBIxAaBLIIDaOG4c42B99PixYuDFsO4AQ3A7N36J0Js0NeN2aD+zbXuTMz3+f53J58UZccMQ
qCRBcyOzrdTI9Mp+SzBISuaoyXJ7Jp1VnZx+a1uUAVscMqVdSZ86Fy3FU28jwO6Hl1q4L3j49wb6
cAOaYVdEAMSWA41wxXYmWLoj1bXJCXp292Rcd7gZQdX/2ZIBxMQrngwtcpSw788L0ekH5+RcXLca
0mtJBb1W4IABfsEdD5zSSTnEUappQQoitg+LZW/HUHlrF4nzGHp92YbT6VTKv3vfxnwP1LfPWvtC
ojlOPaB2PcMPvrgoDR7ORSxFK2GwsIR6gZMXVuLsZsbOWEAr/Xdi9Nm+nIZTiICFZzZawPO1IK4t
HrwHopiqz00pwvyEscu7Mixn6QvH0ujxTrI+vdAA+iDmC8bzcQ7HLZaMI/xwhayh8Mvf5bmB/tJk
PnU1FyZcpzdixmsoSDNF/iAFbkQm9D6LTSvXV+yfHb1QK+licA+oZB1DdTky4zaDvtoVq3pqgapx
gTVPMBTYImstt1z5b1AZpLoQiC5+iyjJe+3KcXGTWfu/DTuttsAgPaYCWvWk+hIImCtPx4HHXmxC
/QSItg7YW9LC42yuApvEt25xX0+wFOxSmJr7zYIYJ+YbCsNmF1nczuVfDCwL8UjcAGXM1U6yn8Oc
g5yMBxK3vPLd4iTnnQMbiNEvmPHYH5WQOzzyh5WR4uZR9ufqDtwn8rQRnMqeNSSO0YjugNM3+Dbf
JZu8jya35TOX5xoXD2r0PEtNX1IkozR9z4qgjMd4QjFADX2eYxFJXQBo+6eFFqrLoxa52pzil/MK
mdrnEyBDfXv7DwSypf3MNAy16TZWu0FqOCm+ClRiGpJRux/nsrPW2D3mIEnrQOHHaqomNKrFWIG1
rE1sjIwK9H0tUFL0Zxw9qPwzebn+480Qd7Vg98SKgdNYXMGBXsGOQLBGA7RvHMHNVfTzvJ0p6+5g
O2WMNiJkrDoZ2ls/wJR36U+MkztYb1VBszpi8wJ2bQHKWeH+SwtBJjCCHmY3SaGRL1wp8lfObn+w
U+9YeWhH/xZp/V2Od271N+jp/u73+e4X+v2JxFmUSb2a/cR//8YbGrPTCSEf3S7Of128EuekxDcS
rCEk1aCQF+OmE0kITVs26DTguN9KrpmS+Kqj3WGycDlFPB25N16Fysyw3IFwa4r8EQkOVCWnQPha
GzIkRKRuZ3NtAnDZJdrx2pnN5ojsn4bI9ibxmtkbw9W3KONVa5cym4XC9DtqS+Zhfir/alx3Ujww
WcayQxemFxF8/g6lqnUtsz7/ooB2h9cx1zBvZmjANNfnb95XEWUKb8N1yeCNcuiBjiIHQTRhlSJ4
HAJwos1GL1bGP1TdeKoHheIYTIl8UaoqZQxVUXYB6RbWnZ0OBdcEikLzW/3B7SVtyu0VSFnRd92g
5DICTlDG2VGTn98sEHOn9kEy3n7YwYZtXlICI1SBq72lK90zCyEtc5V+5BVCUTnsB0HHApQWc+Jn
D97zNo1fjiAJ0U0DxZmrvJuqXM8ED9H9U+WzxUseYV89oBGfUm4xsY5r5mJ64clkHsWQX7ue1P7D
Vdv55faNEp3Ei9WCaxpQhjBzxy0/9mbtaQ59QuCf2LkaP2K1X75mtBHIZYztO1wBTjH3eHRybbet
yXJZZ4fMjx5GjMwSWN4fHqNpvdlZGrTfTvOvLBPRzEURhZbxi3DBfxktrZCoOJqjiXoro9cbs+HZ
YkbSLXozOqiMSy0DJXF7gzoKd5PYES9lCFCgyqTLJkuv/S9maAu4utQg6O6qMWTn3KBzNLKGymgM
waOzLLpFt5hPRxohElUls1Y7FgLkKNObvNbTlPwndKtIbYnrrP2ivjc04Ywi26pVe/iQs1/0o4Uw
CHzgq1s2Do8XPt7zdppV+pXo4nl8CfWFZczKNMuPtcKV5sdf/dnhQY7dJL50AgA4qxWfS323X6ln
8SQu/aTK/r73sJBcTh03ejWBodhjeh4DIGnER6ylPVAaGfQ5D1uR7h2pjB/gslFk4AA3UpHh0KI1
8AzSbTi774x0TLDyQhrgU4vF1qD8j6i9xmhlp7MIix6VbWgSYx+nfWa5pnMw8modkELaAyFlaKg9
9ufKFjLYOYL95xnRVN75UQKT26+j8v75eQayPNMWEVyzuSY1cfG4DSKQJXQWDjc5WtM11MODGRym
lI3+empx37QH9dFD4q7x2GT6/qF/iZZrCGXn1JSvgawUNvHVL9+E9JqlKbNLu2L9FbhWLjtQJ3Np
YONMgF5uMNZnNmRXeNx/ejBXh4wRpUx/Olxv8G9GR+Y9sOa8itwZpBHJBnSUVVFFKxj4Meq/C2bD
vTeVO/aBuz41EUgTbIX5fwEKiUaZPo4cvDc/qMetXXiKg+UU/53/eHiVtf99N8zQ8b+ENrMK2r8l
8gX6hCwglS7eLMMXDCbbOyDSpdE+y2TxFlP91nVJ1jGb5IKBG2cuVNd2W598UN0e9o0ktQJN6er8
YrE8uE6eickjixgDPKcC0eXZaxK7jLki2VlAtjL1IlA6JsAtqIShFIN22S4SBTr2lew2TsGQOl4S
i8iRJMKT/6XSRDX2+G8UuaK+En076GR72LtwUQ3wdyFLM3VVhSZphUEHLiWRnuGx5XCEN/yj8Hzf
HogoISHpeHrFAFRUhdACLtIdm4YoxtRoRpUqX6jOaeQufR2ctAZdckJzDJDeTxD65ssjC0m6DtNc
7lxiE8joM/lZSlPifIOvtqE4qzmvM9/u4FESbpAK1jNtH8iPZIdtjtXSbAHI5tj/W0os2Q+qpvAG
O4DImu5wiQaFw951pRwvQXLGNmaAf2APilYxAMOR3PiPh7xiJns8yi0pii1nDNQXHNdcKBIWIly6
qI2T4Kok35BBzInUoNhF7yTi0xBq6ngvpdi0H1aAY1M6XC/wkcAbIRQLGVa6gzukP0Pz6/64aUij
Plm6doRoeHaVUYAIo2Bz9W30B6j7oYaXhBT5iALFxBslUBHUDB4KJX2VXuqMexudyjgikYBBv5an
V6G1BmgT2WD7FBAqMj5cErGxtYaPBOjGRJFdp7jhhWOWmlqitCUB8wHxobVx6fptmGjhwaFgIr9C
g69gAgUB9vt93+boYTGxdY/i7yVOORfWhkTsxFwxeTnBmVXrKQk3u2I/Y4rq8fW+niRX5vsJJb8f
+D/5Go8aRbSeMTvr1zRiLaxEGEYwMElk8GrulgTnuXkxOwMy84VbNgZn1InRXz0NkJeNljFAjU0o
q0I36ECtOI3CqQZBUQMpQCWOWDVQ1kT0CpZ3jzVX+kjLCp74TGDt5UQ5JWLKHB7CBfGafYkLajoD
kHlS0NjXmXZ5sQsdwoBDnDZOKZsc1N+pm+pFux/PprgdgjVN37jYCmC+NIuk5XIQBlt0g3cRmWjW
Zuteop29Ygu8eQowiOpyr5+znxbzC6rUS8FZF2Aq5W/auZqVmp7G1GM+XPiccXtIo8Vd89OlGZMD
swtuzkty4B5fwbQiAOOoVZH9uGl4fEQE9zHHS/cZYySvx14KtMeGs/bCMndgkDwNktUq4qSoxg8a
jpFC7S9QfCvABxW96jux10w5/xT6VXKD6ckap/EaBmv6mfbI2nBgQaeLh0DBRX6t4swImo62AkxZ
69wi2oYesMFqnfOt6hPn70xr1C3l+gi3ny2F2SeFvehf03zVSKseDfCMJkcUBYzt7moqOKHdcsnV
4HjlhYh/oFudXPiPKd0mhzqwH/5UyL/GvxVKUWW51NWBcN7L+5ZF9AqYXciWOPJGDSjpiECpuC6r
ceRVhY9RSah/vjue9G33pDggpl77QkEHMspJEnf2onGwQ8oGeRcq1EHcoiSmNOs64BumfV5QMbNC
EDfHu+62SfzZXPQEug9YpjQfXtrdMdGJsA+MhopLKQeXA1MwOm6NwNeUA74VeFy7xkgjtLKpHzP8
omG95tHKYvtI30FCauRCEQ/Uq1mXZMU1wEhZv97wrL5Mp8/M++00nXeN2o1NilztHdiuJOD/funR
F8bnu5pTkRdln+8KHBjMz8cTIWdip+rzgVSriHwBg7MNvhU2nnoLQavsM3AMSvSWyUgooygjzMfo
icng8X3mRijaHwr3mjfbpv2k53eSMGEkZoX8WCa1qrG4aJ9WJpLPQSrTapya2yi6WbBHrYG3TCfk
WxZ48kDNZfeK9IRe973158lZc6KRoGrfXFgJnoKZ7oVrIkJkJsYkwrgUaU+SjnahzRg/sRWDpA+T
EWOQgrW4NYLV+VHJyi7GPWffaLJ5LR08M1cdrsq0oS5koGypdCTn/hM/xW1uVdbzPX0FftpdzpFi
Ror5/qzNctYJ+JCgpL8rqH9FsIvVJ4ZQFJRGM2qlIA3j2FKMg24zsaZa+7IXxNX37JcKqHlA+Xrz
cDrjNeSYVlYdTjSH2rpO/OxSKGojOlOPVSDh0eeaOsBw9SdNo0PK4vP6WPb9DRHKb5TsSm/SJg86
kiDdVVCs3M5ASGzO3SU3ZLNOgY+dwjcI+JpgzhwdTZZt8ZZFKCn1EoQotL69FdZVBRyCalnkpipz
iRNKzrnNta5JVVJKRL9q/A08sqq1pQpZwvw222d6CjAJa1VkvFfiv3Amh+DWgChv+FRlPvTrs9ER
vBDc4SJZj6P9W9NSD+aE98Lfoj5EkITMIcSFICP+xwNBOgX7iqfN6AyxD2Rz7pImZGO36zmC9bO2
P7KeKXXp3DY7vmpZVKF4pikFQGP/zPSd+swXmchaq2JHnu53uFCpDD1WPS0LsI94nNjVWAXhfIZN
pYsjC3oZDEaV+hD2vs2Z2SwYcAhdkj38IrNykXH9OjvnaTbHC0tLj+T7F26cb9zdztuC6jcr6P3O
RXy/sstaMbDQoFkNg6WG3kBuOZccG17siPlUi3exurPynuRBABz/hpcAIaBTrl8iwQGD++YhS3xi
4TPhbH/Hh5hwCwYZQgKJSuvdc4QTw49hvTAtqLibNp+Y7flh82TvMPHk2liuULY25WQ+NntUFukk
eaD25B75q0IRZOoJ3GuOYW/ZJRFQ0PO2kPW9MOYjaCnSA7kH4KObuJazs04w0vbJdeAKG13u8vJ6
+TQ4L6MR3vPK6oVEW10CK+T/n+2tWzgSGEm8WJiKdmeS1Clp1LLdM+aX9Hwtf6nDbuniXK3g51Ba
Z4dM8599zHhBnfcFMiLJZkWpq1g/DXfzhPhLEhzs+H6xtSh2IOQgGSzgu8XJsT46fdBLcRSyG7Cl
a1KOtSEIS7qK4nS1I3mcTd8YtzTLJ2Z9THsdUhIdHd4O9XnoWaDUKPo0reLfS7w04Xg/R3I5llmE
zM++ZsGYZ+t0u+/6QhAa0sygWRJEjSWHGemUweh2x/LuOcbyJ0GMyhP3YeON+C1dYnB6A/Ks54e7
Qyyn41IKXfnil3Jorn7B9qdTw+jE0XICsxvwRZBj2YK5vlS3jD5h9LDXobyFT87V5oiGREx2tWpW
xjh/eyMoorKpUtH9TnQj5Ng9sSiklsE95xaFYB2/A7JEV9egnaipOxkQeBoCG2kqIvRXJcXSUUve
GLCTuN/Oykg+DjGh2urv4GBs+rSvH+T5CeOORw8Ja/marPWc7mzpHJ5r32ITbqaCHMH7450ilygI
fWjhIzgAhXrTJvjtNyXam+3iyiaR52IZrlBNysNfuuLbGwurqZf1KvpVQZyq8udsDv88sVF/2jOu
Fwg/dbuWyH61MSNyFr+6dGeoWas0wt6N+Y5S7P7NalNVh73QbD2ZU+zoyPS4HEH3kxB8uubu1pTK
9jy1VHwvTFlvlFQhPp12voinj6vwAd70+3JCL3jEz26wkQDgkSXtR5KAmnYfE60J3061Q9We6Uab
hhjFNxbKPaZ4t0w3VZNcsbUP6eCmU1y1BpfJ/z52+SRggdpnJxYjroyD7qI2S6YIME9c2ktYIJhP
rSHOvJ5c1OZGm96qmkVNAlUOSP133LoLF63lY3X7sx+EZugMhgJsShQsVMLiuTktWMnPrXBN2eno
lu3xu2pRRPOVajBeYJE5CDxXpOA17PxFugLdXD85Anym2tX4+Q7a8k0AcMYEVMf6+XSq0ylndvNs
0l9DtmZUPe6SEgnIjwWXK5VsaBwqsW6niUYJ2vAdMGewZUgFd7yFFAtGfrRyhZJ7hxacF/P8XzBn
0TEOnxoj+EAVpDvejH6Haboidn1wKaaGmh5WKCYZO73gJBeBaiVpU0XIPR+07jrxfzbR3ypANIpY
b7T25A6F7tpODec1hhvHhAbLjBxIuKhpdsHrFaiDHDijOwqTgVz54tPJ+PfDemmdfQ050M+5TQFr
JTtb+fWNsCLfktOb39qxYRx9JZc+k9i7D4+ojTwkaZUgVoUEg+Gj4L8WcUMAzkP6HOgxF4PznNQ5
v3JAelPnPWaZmEDJljF1xWWrS9zhbe6mn068DPmFbqNhiKsH/XMwUIOsJOn9HoXXUcfobYtLC9dK
8UP8bE44MDZXx23frlg43f4PdkN0TLdKCP7YJP9pJfnT0i3FK6DgbOEWP46dqYAviBeJWVPqCAy0
qB6zQG/amqDwACYs4g7RnWD/HnDuEdDmc84jnIPPy+8irxEkQCnbTfWDl672A4ML/YLa2sv5u/dT
0FAQTIX4p+loGsycYBum7bcZYr1pASrxNjbXETgoM0TxZZCnqdsf2EdPfur3jGTP2d2RsP6BHIHG
g7dsBTFLJEMLtA5TVL97KdaX0lg0+3KNzh8KNWBhPqsdJNCkGxkZBZhG+mrh5goU8abdcQk0TadT
ht2RjulVL7EWa2hLUuEu5Rvb3cftf6AK2pMY+c/dS9WgI2eyK5OIaPTrkHs0BL0gxlocVZzBx3+a
F+Lg1CfdFk8qJPH4LUCAubPvl2UcX4Jn2Ok4P2ii7fJAo/P43rN9eQxTwQH3XGO9EdxaxdCmJgwc
paIYUExwVVQTwRdoW2H9DsPKaolzMzS2mCsi3FDEclqdghE90DHBdmSqZ0TvqBy+jUCJceUrzZPN
3GB6np6dhj+MlOi+rQYgyiKeMJxB7KHVaWKj6qlke4DNfQhJdfFXawDR/Lsfwr5XbvIx45E8f83+
3oEsUWeua/7e/vaFe2RgVdTbaAXCQe1ryUVZSOj6J+FFMCiC3c9xmqgVgS/fgoyzvz+Eane1UO78
URU7yzJ6nDeZDuB2V7sFGh2ksuTohS+rwT1fnjwLmn2NCMmBcIr74ho7ie0i9gPb2yajJEGZIXhS
HkYFPAhXoStH8qaQTWOXi9coWeF5MG6yL4Lp9RLXUNhywHgrO7nSscrvWLCQaFn6Hs/NGHVT4VAs
7Qwy7RvwXbt6gzKvc0R7T+W/oUrs8R6a9sASJhYlzP8NbGRieiQ7GDWIIdxWniNDiKr0vrGZ4Cva
HPFfbkDgRFqfiycelSZKr+Q/DtXNFDX9pypHOaMv7Z37J1MKopng/JGFI3JKPJw4QSUOyHUHPj7e
GCfS1BjNrC8phhAlBHUslMtL6RaAW01HpEx/ZbaiQXAUmSq5ZBc2SkXRUMz9E2P8+Tgr707XMiar
izkrwBH8g/Z+44DPHu/FgQM4vHE8nU12Jeev9GcHGn6MrpQQiJ4huvalXXz/PlZoIrZHNM5L9Gic
S6ta9+APVRhyAbaWUW6ovr6yVqOD1cKhg1gygleQ2nL1LMCZMNIh6HXQPAJZBjg12Q0VpkVCT0lP
KnPSSb+z6tq2D+GtYhKx6NSj+Si1MJjtO84sGgURi56mZdfeNAo6f/v5kCW/h7uednVB8DMfy5eW
nezasa5qNn7C98/Ix9hbdR9ktJf6ypkzzOdYmxOFPeP0x/i6dm3wr8BGzdBAgq0LvvedMzLX70/8
E3E0ZOmgm21u67DIbXjSnqWU+uA2qRvK0Jsk7pDkNJevbwdD5AGXHnNAodbixzzJ9JwOOONqk0Ii
CmOI5HWMzLFM42gBvGkZm7OUH53245bYYks0Mq3J56S/ew0IYj4xevyJjFcwJY1bkEIeiX5xod7W
xoDKjkqXuwfcI/zJsrecSK+qoDWQFe4izhtMjklzfmjiOA3DSo87nP4K3FN7G9i61vFWj9qCWQpA
dc8mQP2U+CL34D1KAn/TsG7IGiLmUXpyAFCzYsxqLGCrjXAHfk2A1uwwHnOg0rADkeJd+JMeWy+M
9l0Pa3jZAnpvYfIsXHrJmplj6hvRIJYfPG0D27FFaIZBVJvcsVAdAzaHePrKpBY6rquAsD9BXzfi
UZKmfTyDfeRCC2R7+03szDdZebsBXxDPkHHqfNnWWoogV7010mjFRqC8iKiEyJCWtizMIK1sjj1x
wChhZQ97r9iS4QaY1kgZWKh1MvEPjZd2DL311ufO7D5velkATiW2rpx9kVwbibfzQcUltro8KCe+
1Db04q1j/hmJkLG3m3GnV0oUQCr1VUMF0XvJ+8G46EV5D3PEOKM2qfHo1L3H8nG6OC5eOu3b98+X
2WzeEEeSVwqUb1jyvELhTXVBnjuAUnYHrXkO19o6AnuyA7Ut9CkpnMVdEAYV043EdmfoBAQOGetU
BMpslMq6jL/8LOp+zbItWvfeYp40QPn5xTZ0AodTh0TRzr0t8Z9e3FCwflvhJvjQrVpB9sXrNIq6
ZCuEUDnVUGNAzxLmpwa7MZPgb+K1nIrFXjywRzw5PHDmefneBpm3EsvqjvkEAKTIJpWVlb/kC9ZR
ur+SEQsIriPTMFJhyBaJtrLvyS6aWGpTteUbA2RVGcU4TqresnaQugbS71qDRttO5xF+lPTSmd79
x5vFDXWnb/lhkPI35aKLWZUCImrQtUdZHfG+wBAMzRQ0BXNnTVuYgk8CxliIdj4LBT4b87G01nPc
sKMwWvLLL1DBs0kix/P+n42XDzt/2ShBi/BAyWEqOgqsDRDjiO6HBpCp2usFQXiy7Bh3+3AYPCXo
dRP4dnB37uZM6wcmSw0k6HMSy2m2DoJbujOwyZ+SxFOgsiuxjzVFrq829KOgoJcL/uLtyhLwMBqX
TnUDoboLUhhIz+6eK0NNVYNgdiCtIsEbJGGweWwiWTZqZGpv9NFgK9GQmJNkhnqh8BmR5CWgEBUU
0TKlASUPBEycWUSnySeQLQJ7Mn/p0i5DALZwawZ883GXIjUSr+I1m5awGuiYnKlKWd8iBCDYzHt4
l8d5muSUqmeBlRbv7T1If85+wsuQOhpvc9xBxv+OmO2GktZ4/Tdp+oS6SmA1zhsUaxNbmiWHPOjc
NVGWHy8ElMpdVZdjuqdm1CXN+azSLwVgEaJUIlqIkS7YEWxBF4+CXy9M1yj8C8YPlD+M08vrv4Mb
ZnObLn5T6hPSjgQiY4neBykcJsN/j4f34ZrwOKJRsB+Y71Dew9XaWeoVsdaPGET0/ridnicuxPUu
q/AuJwJ8cuozKghfuJaKgE+wYETwwzneTM1fBy1UWZLNmtJehB/BaB1yYLe93H/oT8lzbe0cr4gf
RsBy4E5xaIRdxJ61A1tOMPavXjBhU8dRg7cG6RY8VL6LmirMswtQu+9lamYhUgWumkdgYX7SDeyT
nv8A25HM8cmcKb+SUQF/f+ywaPLSUPNGh7GTX2kFbDBF/ANZqqIu32Vaw1VvXAmhCR5OyITsUQdo
GGW1sByhk8sECGn6VbQLz8C+Nu+HGR6kvZ3fod7AZPzinasulWLyGkGu0takfbS7+vYrUE4whuAV
S2FTzMWlpQ0j4k9D6zmzts7sP3KF8BvKMTWNYaIx82EueqHSi09yYSqZvouVmGdvwCHDm0EvbYbg
JApPkQomcL9+czIN+s/3jx+nRkBMBYMiXgQ986asehmN9y5N/mnSOipnJ8m/UwQPrJmB025JlB1/
m3RHISTRGE9rq1FKpQaJQmBS9J3idCmXKAQ9OLx0/eC8DQbUZEqDNUNmRGkvOdYHot7nHXI95iya
IHo+khe27b1ho5tXbsEC3RJK4ea6MWiBvpgnLc0p4kb9np0SgciCGgIAiiRl2ImYG1/Au+xuwbO6
lbUN51m+Vwhpwst4jJw+gHKfTI/XPNZsK7GLfUdU+ECDcYFQFoZLGCW5Cln1Qoua+OlF0K7IhqQJ
dKf4QtUKkj8cSuVQ3kG2Ep43JqV/BpSuNlDTP0CGjCjxXfLx01HJk9+ORJIlYens97c332WNCOR3
9VlbvXQJlKhTDImd9Adxf8qEzOFPIfTD0mysW8nfq+/QZv8kSH/c5voNXxhLdN5GZlNZWN5G+3Kn
2g0WOV23QpT/6af7XC0MOAGT/elF7sfilPJzCxLizsu2s+TPcMLKLDmG2GgKIx+rEKn4/EtUZIK4
xBEmNRv6PjJjS1etS9maUruK3I3MMSnyARqCOjQuGunq66y73J99aOsM6F8cSGA56KJ+d5mGU/kI
6Qck5/FyiwhIRgeUkcodY1gq6F4bd1M32yk+Fg4YXHXvm0eXIz+GyokyCbeRDo0OGv3eWTzlYOR5
3xsSqk6HFeUgp8cn14jiSpANUVAoFEN2vqhRP8yhhZvh0zfb6Pp6Bg4mSGnwJhjEa6UAme+x3Icr
a91IEDLNcNWQd43dnoisMPI4rxyc3kjp/skHvjFO4XxD2OSSAR55gAIklSzdNmrHrj8u9fAaO16+
U05QjsvRrZI9UKBSA8E4/WgqOMSwOgwuuCwC5yAVALm11E77+x5VXRvc0PfTMWNl7xar18RFZnq4
XxpkAW9XlGL/75XDv4ezhPmjRfi2lxieHfdT9Tq+9Iqa/DpwTdxhwFyt+7bRTeKriwhHM5LWz0xS
o2yA6i/42VsHMlEkuNfDfnDpMgErOU3uQas86lsBg4EImDkoUfIWckoJzGcikcMSQ1aghVEYMg6j
efvvEYGHIYvbzhLddUB/ADr6vHZ5HjrcimUD0EjJff+KFkMnBDZp5ghM075NtSIKjn/LOdGocz3b
a6eGg0MZP6lHb9GmjCg7De+07bFtQr+EadHn9wGSrIPTiQ/WDaVkBq2Zjp17UlLvWxxb9BJGL3aS
ENrC5FuhCyAYjYkcmZW+b2NRt/vSDKkv1Lfctzu1GNGvChDK64k35ZPbrng9Ka3mEYoBNt0GNL5P
Xh/CJzorXsDWHjW3+ItBbb1a0udm21QyOtKoiG4AvsTdbJ4FyUo+K/v44bBz0JegB6MbtggxlJH9
tJYApymVo13n84O8Luek4mFaLpMHGhokWLWCl6fTrmQbaM+SCawx7kN6pdjH9S+dbuNIdwqUh+eo
kDmQluNojKq+dMPKdpaStZsEQ21QAlqy74z3FciYj+eC3OU5XCjw0gchMhSAfTlY5rwE4h0O0m6E
U+SJUi6SjCMLVjZC6vIkqIdhLpn5p6O/VxGGg6qfJ6h8Idg6Z+qmwRkCn3IjYdRtXP/H2B6016e3
iavVjYegxCjpiOWaf6P8rSPUnXhD2YtUXsjnz6JTdoGCNAesHsp+Ta9zNmGl063TP2ztmTfUjhDM
BTJ2XvdmF3nDAc5aerTntdZiixCmu96NbpT6XXboyMT61h5s9tS9s60RKxM1YsIQ0n+C9SaBfT8a
WmCwWoMzRnGGFlrSqg16FAatBHUuIlFn/kmfr/WvyYGfF7U276Iw9feyp8jEXtU+tcsRJ+1Ar9Gg
kVkhH/YZejuVMayo9/bEZbQoxwmZz3lBHv2zHPqTA9Mz5liyOjZZULpYh8QuNnG4Q0l+f4MvNka1
xlQBIb4jMAXdguMcnhEPzLGGFWAc67/DluQWoaoNmR+KJeuVLjJeSORcnyWuk7CZjx3USp+GUP4L
7SB31vXXDeJBNY6978cyQnoE7yWcE8Vp3DdxuCn3WvUlFU8Ks4xuOrB0Q9ebKk5G0eA6eKz9TY5F
8sAPCy2mxqXHIHSvL1xdEXmAyrqAILmgZNNCgy2jmnufRrDSwhJlYtwl0Epoawknxak9HJmoSu5u
Cs/AZW5K7kqzZL61dHKpLgBe5RaEeeNn/a/6Tok6FFH8iZlg29dFO+HgiKV0W0xxwFQpQL1mwSxy
GkLEjnxmfRMm1bi2ExiT6f10RIXnYJdbH3ZfJZHPNDYV4gR6H697AeR6aJK+5etI0byO8Wca4LI4
ePW//9XZ7mbLMFK2IIHtihGwaw5ZajbxizVwxx/hLQmCcM0Ct7LgVxHJfkn3MxII0lYxmEXoC1rX
HXTYssTBwsaLJGVBcSgI+OgSnEHV/zIJpqc5CWDusS2KMVohmuyXAB4P99TllvTmVux14GNDItF1
7DwEdzoXS73BB25ViYBv+HV9PqlHyo+IhtdRiObqsfE4hAo2WNMg5axgOGj3p7PgtpmAMdQeP7XS
NeNn/XLDAWLWrWx40p5E+6j7zWmS97T0Dt8Msg9YX9VQPUXnWHahArwYgYv6wMeVveaNYNydAQgy
3A9v9juHsul2DDoaHgUcdMtMpP/IbtUp955QMhfw1Yh0fwjEYpeh8HRFCC69anSD95ndEOJZdXAy
MlsW1yGjRU6kb2NgZMgSQs5keoNKeijZtr3JV1qU6yDZNUBZDPb96B5R3KpV50Gi4mnjDUmZnP97
0PqEjHX9pgR67yoHDLXYYiRDbEQJBPRioEABk78kT4E278Fju7aPCc0XtqS7iXfWk8rwszISanu2
T9j0A4/namBBkADisvJ1NkmZLnzEBhftLo1KE8ejaZrVN5B1O6eEeEmL705M9/CTpaOxsMe5KQyi
3+qOlvEwsq4G+SIln2XkztfOYvGnXBQTHwO/jrNucs2j2CB8z3ZvlYblfKZc4/zuTpYa841RJovx
Ymwv+uBGVAZElJZ7dPxyLxgDkl0wIBLvK3XqUanHyoa7vGZdcSIg9I7Wy9ec464jXqWQLF190Qc/
CWeve8AnqQSImSefk8/VOUCSgoxPPi3Ajq4V7omx30pe8+JMbWW8mAJjv9EkYYclS5VNxVTQDtDC
t2Dsr6UZ6ROXkg2f1C4x4s5IQuEl96Bv+zvGMx/qepJTLjSfX/3/F1/tpZ+FaqzdIriw1Q4ZR8Jx
luERVAzs4Hfu9VsStFwOGJqIAGmamjcwS4e7MVIYJ+oa9aLg/GLvoP2KfmhI0YBxvvAoFJb5XGUh
1pgnBe1SU3X/ZHk9raTSonUI7DTzsLDK+HasCVO/r0FIscIcqWhrkRQ3FPYkLtWgUEWCTUObmK65
ErD4syFgpLAd05kG3QZqnZP/ZaRoh2ce7wr9Ui8BntodYVZqphTxCTXH5S37yCu3XMEXsWwpX5DP
xo1qhJ7vJI8D7GfT4SZSy0VBc6buFHB/n/28pXuQ6xm785+t2/ckxQzyyaffQ6vCa2+L6RhujCK8
AP6yMVLmFtTr6+lEJFNd0woQVR8gckFQ85mnlpgEvUhm45MvEgJV8C2/SlCC6DcxYZJvxElJWm+e
psdVbzNeoi550CQmkd5II4ylNVOEwILWUlcHNspscwXMK6ojQBxpA1Wl/JJXbHJGaZ/nLdvG8GUk
Ovdyt4IpySawN1JbfWUWB7FkL4bd1mmvaWnmrqIe4UAQdNnhwiib9wTw3ZjxytO4X76kY+21PQfK
+tdT7g7uhmW8Yn7RRU259XTblCW5nYza3vQcqpIl3eZC0yz1KXkX0sHcKNNxfCHcfRPok6oWrOcp
8aUf5Y7jJLKJu7msRx61lm1qmAQOVfC9Y0mEgnaZfoggic1RiI1CBIRjeWiqliUH7LSYp+ug0jrY
VSOCJNt+YC/2nAPlAPa27ZAk21v4DQW1oumkzBdhyIAu+ftzBGzviqdtbn+MxBBIzvInf2XEgtXu
3fvMtXe48/fb75dAVandhR3fkEAmQ9XKBuACrLHf2mcs0/GlsLsF8WGMgIGJhaMd6y4XBfhh0QfN
rwkPDu/Kf4I3kV5lBTsim8MoBUFg4sifHXFXGb3sRwnL5l5jJTRu9zRJc08CXypdiplP3mmDtqIs
ykhjxgzpfRfKmfs1cnJCyU2w2JAp6QFazxauLy803yYs3hzj9KJHOih3ENhMT4i2FMIsQGJ//GY9
i4xANnVRccwHHqs8DBo7SLT7KzKjdpgbP8/ZEGoy7Cgnus9Zh7y5MoYB/qTlne1koj5M4TbgwpWj
d84D1umr8SOPJfZEnmNi3LceKQ9W0of1CxNri5A+MG2+BqSWGzIEXP8vcEA/DGQhu6IBYHDBWxd1
676t1W4B5EkwBvujLT/zg6YVZXPr4QmxIzRErHp5EQ+Eg2HzrAVsUO35b9sWUVoYSYK+LJ0XC5Xy
ihP9k1M4noRtwDE7gM4gqdmOixOEfJgBzJB5u7ozWnhhi48YUJFYy5j9vEBDzXJ4nMu62U0gpGDV
s4fT7HNMsVp9A9gTduUOzFGD9uFzc/Vf0TvhHO3otp0gbE9OdJbmBdth8+M8xQoiJPE5B92v+FX/
Vf1+h9HZ03NlwQqBs9bR+b4JUiRgl8DsxUQsqwUuPynSQD+BybD2deKoreCO/yZdU5SDUdb4gktM
Myc9RjvcTFMBhgxqg7Ia1iT4HjCh/jT8a/nrcg1gNXr0ljKjVT+nxBQNObKsvLVXIcWptM6nlJGJ
ZLs+OBikRA1Kr+zJE95Ty8zM2nAj0PPkjnOyvIKD3Z+yegG2oSOWCX/UXJWIkBqCG4uFwGI8bsVq
2yZMugryoACBpCk7KIw7szHhqD/ZX4MGC1PNoLkrB35vpSAXRvu9ogmlTYeY7LgSy0oZvkJMPl85
BUmxx/GA3xEE2q4kFkkyqvRtZ6l2hnnN8gy5aS7ZT3V4DCzDjmYK73lx/ut22Hp0aZYEyMw6ktKE
BHV/5CBKDYLU43DKAYYalzWwcliYox9tS7mLZIA1RYQqpHWC4F0uF9ff7SmO5Qvgh6mJvCMQPSwg
nZBFRuRIhmZu2z6to4NlJbdL0e6iz3iv7Ecilg3lbC3D01hiZSrs4xMIdELgktFMef/0G3VbVN7g
l1fVTK19VJZ3DgCEiMYTXB9hLC3hJj2d0Tm1+cCN2r9bKTmh2ydea62VExDyX9g35kiGSYG7pIOe
M+uOGS7YCEPlolw05Pk3ZwtMzU47afisP/JmkcyEITzVyOGspn7R5yW00k7KpcwSGIVfpESnZrKb
9zwUaJSvKC8sbRFwDrzW+aBxzr69gb2Gshd9BRd38rs8fw92TCw8JDzQ1ZC9Y9tH3tsab+gmoXSF
Acj7Ew0r0MQ9nzq10k6DodSEYKmrd2kzzKst0ScsR1sWUWuetgoBFu2n84GjHll+JAN0GR7E8vbw
xjOiOR2gJ6CGD1PaCg7CYK2det+Bpm+BVIghJwSvFelTOMrnfylW8GNdiMRSW306r7h3ndGsnqow
RtVgO6mZMu8KAR3kZEqDrgvMcjD6snZ9xfJcxtmVGtyxxPTsqrA3KvpkLyajmhiELYhUnsRTNo/c
edNvApB49B3/5kOFueXb4/FIK1WotpMKXw6vBRTwrNgbsheJhPIJKJaH+IIZyjxBS9vW+b7M3B6V
ZpP1ozACPdH50w9bMOPFEr92r0qXNVMnVcP8mmUipAtGI1XD49D61Q9ZQdstg/0hTqpk1LjqhdMO
Fj9h7KfAeIeK9tLbsnMvuwrIkD2EdE0ok9+lkUIprVunH03q0ISgF58mD44CTxUCCCBSm9SI0aau
LjVQ6JNTq4uDP0a5+XNYZtp56doF1htEYjSbNbwHiPC/E9AtD44I5/DyhnCh6xOS3q9SEeG0D9cM
bmI9lcRQvJbkiUFLg2wSnO/OcnA34MpErrTGR/lvjIDNqwE6bo+oal7fURgUxHZcyn55S5V9FDpP
tEVQteShoYpqtPxvEldGhKUXCx0oV7+kmt2hzM9DknEOabi3mbVCDpx70gDw3WZWgKjVfyfirxnH
s5gf+Eb57L4vpr8EA7k1BIsxddLHgtO+iTLkNmjcdB085vHN7ORthv/HQYt8biyq37gMRdbD03g+
zCxZ9AbqcSRpU2tHRGvZkCOFmU3RzrhETlG9rbTJZB4lFg0Wbh8wE/HOwC8PB+V1rNbC2JenCLwC
0DImbpG6QelXNbllAu/KziA6GoiPPp/gJwsYg0NTpmsD0TqL7qCAF2NaK4CzTX6brw6jE6HiNKrr
CnI3glvLVQe4kISAon3RLkSFQW6zpNSxe2SObyq5efKkkX4oQ2TxYkf4UMzIM99y92F+EC05hYRA
Rp1dINx/vuVJoO4EX1iUq+804LtA83SQ66aN4NMKpvrj9xhDyTsTYoTbuiFlvP3KyvFlHLWPJsWR
InEvNcaWV8FoY1/CwqDeTBHQBP+k4UM3Gm57bq18xvCJ31pO2tLQ8omuFvleBiKZcSRSaUxQqeEg
4OIQq23kVXsIoQtkWMZpf4jmg/5/w85U8C1I2U8a9hcUzOFm/dZftnH3KahRMVapVqu4L+mkbjkY
8n9bZE9Ip8+haGtvVRcqq5dhSXNmZiHjHQqH7IAisFcQIlOlUkIlqFkAesJSM0gBg+gJClpnZOrO
5ZEM/RxPRw9a2TBkyAwaClUNnuei/fbXmBmSA93xEoL6G8oY0yxi+FArCwrqKIYy0jBQYWs9rADe
qoBL5QwkC/P56v1yT94jtNi0hixsIvaPiFcv7bRrQ0SThYPfHECHDDver4RQ8aKj6+mWtfSnwFhh
Xem6Sn9Oj+xmYgZnH6/48K/9aCU6+ZD0ilftmLi1vzb1GBGoN/qNAiXDFnfY7ev4ygLIoEE2AS+K
p0igy9cNjpSNjfwtz+IldrW73idHNdSovsI8HmJklvf+rLJ9h3QW7Teqwlzizx5Ab+AmISh5NAki
cNT1+z+e5suEYaBJQIKoNjkfY1h6FkrYdrdZ29IeWljzvHCTQkJpbBmGvSCSVGqL6CALd2cMKvjS
U3oPsw2rZzwU3QYXroCCRROx8FrUTrOEoy58N677CSoPEEpGluoUasFX6q8vyIgTMcKqG04qdY5P
Oiln/tP8lRnrM2h7XSyIydX2PP2G8Oipod7a6uIkxgDckSRmkhYflLWeGV6uOTEV19H+cKdvWUsM
/8QRAhYDet7zO2sf//hQaY4hnBTJp7klZuNf5nmeIjUtzqjyedy9Umr3xtzp1sf2Uc9L0FLQF5WD
r7JH66mTLXJ81vz6jSwBZlFqSKDu35nRnChygGvICS2mpQ7YF8ilx561ivqmXS1Yeg2ZtvX0emIc
X3Nwgp7bxS1NbCq385Z03RvFzvDqENZyVc7jctivZqKf5Pp0Ild9JZDnsADkA3YRAvzq6BFNfqpC
NTEkh+bd1eyNBQ7exA1xZcYKFanXHTBjpK/VcVFA4gEfoesl45EriT2XXz9StUPqo8C/qlKvi0Q7
VxqlHpWYcyl0D9sAx83P0M+jP7hZwh8Pgd57cRzdnF1ijrB/ycB3IUt5G+mIeH55vAwCowRkMTwf
1aT5OfCGlnXPv0fla4yMGZHFckUEIxJyCySui4mMaCfZBouiZ5HQ4/3pa5FPBhERjBDbFSYlKygg
FLj77lY/tuYbG1k+AFUrHi49jnblMw2CerQAT4anfQ3zXhvVh8SaUAbBqrwlBGfm6P9i8ZqrBg38
LqVhznRDpA8LqcantWjKmwYIlfUQn3ngmTa8jXtDvGFBIHNBGipnaDFD483huTHkdUvWYnJskd66
8baXLlOiifEDzqrTP3ogDcX+4P9IylwG7+gRdqZoPVm/SdDWmDy2xNOtscXM8yDaCm+NjKapexzD
Te9DMuUf83SPtXoTJZckekocMlgujSWDx1Ua00saO/XD9+o6QFipCc15x+R1uLNDxF1lJtKOzXAR
/wGhdkzsKARjEdKaUIDg+EVoURAhRzo5MruqaxqC2KfOs9DCYnC7dKqTNpKg68XHYrzcF/SWJEPj
WEQkbnJ5OIWi2KS4GWgc97Pd2eBqXdESQ6tAcNIH1pBUt2oX2tfEa6aHPb9elr769mVmmKotwC2Y
+QlUqloDKik+sjRxowC8adR4tIqbMLnmbi0sTmzQ09Wr4wHPae6ntLKn+qhxka6IwEBwkvfG7air
FxwdL+xFNyb9hmaztotU2CeAshTWZ2V789fLoFCLvFSkmo5mTnojMkgqYs5xcAXuN6vltzz/Otkh
j6URc0FXWHUYFE2tjgr1fOLBFf6GVgaNl6iABgAW0yUFwHwqsglKuEihLEYr5NM4gay7J5HyjACI
keIN5P28uemyDzFXN67UiL3/hCP+mAWz1n36peKtVRYCPfWOSyR4gY0vR+2QuQwpybg3/XIh37rc
YO+tcwBfzlgvNVPmrlWDkSxpq8H1y3sNLanbUbwfJeWZ297y3j5+EtBP5YMhKwBouikiffrljFzl
yyRWO0hCkr2VVhXAGDhG35ILckFAMFVYqnzQeoW10cN173IC8pjm5QZaU1Aa18HlIZmypdS0APqL
6NS1nuIs8nr+HTQuQ6Y7nbXsyFn10p/AvuPt0IKA7K4dY+RSOriVk2itg0r2lIVvbFOKLjdT00Ur
cv5cvlxBRCVfwsCVG7B26IiPrmL3F+e7XfIFCe8BUvfesuDdAf9dWWrzyPhYApB98GnXmDCSifn2
DGEBpZaalav75tlUr+2YLJEO5RLxZH68sjKZM13KhVkrQCm4JKlp1atKvKpAIL8BJEs6GcCWgGdO
vSCPtxe1RutmxNW0EvYTpB4UlC+w+KTZpOlbRXjvsuYOlIA5ZJXS70mNRaTmQpqQsyF5E2G0U3Wp
IJC6KJoakD0qw8q+UnT/LN9X08rHUeB+Crtx7XJGhr7yz50wR9yblQWDYcp+4ou4rzstAGJ4cCbR
oysx6nCOy1hQd3/CHSFR+0PJY66a3FJtvbQ+uqeAy7JTNojr2VIO7VpLu6oxnlvPesrWpouVRiEd
we4wAmUnR9R8FS5LVhZL5zlHVyw2vRO6mpNYRiCvld4GEgCumo+M8GbZnasDRjPIc6O/fGvnE8L+
rITC806HZXgMBYnmygy+bTTRtsTB/pv60snPQQ/VETne5lHTs9XVdoB1KSldP9IZiDcVr4cYxbFU
Ab+mxY2YTGtctyCGGC8mlEIG+qS2YhZQR7vApcNVVIH6T8P4DvD5+FocCwHvZzgCn2mj4iihO66j
FdipeAKSSq+bYnydmBqIE1pj8+ZVqGEfiK9yXqyTh6v3LZ6FUhfQ7ajcf8R82C068dTEPxjbnMKg
TmFG1X7bdVWadorq3RYXeGFbUbv4Fvft76S2OTvlXkWcRCA3Ylp6DzwDWfFWg+hySy7g00mcQaX6
xojT6KbEMivic33kc1FnP9/dbWzbNlOUR/fLgJ1tdUiRNQjtz8iq23tgaSHMafQMJWI+MsJpJ4gn
zVu0FrW5Jlg+rHO1FRBxYoEZ2eugfbIaCCNpTaUGaUXXaUCxAjpwf5a2Mp+U9GBX/ZQv9EJjVxCp
2SBl+AmlMP+Xt3VylmoJdFZx8KpArd7nN0yUzACrDi6IXdPq1bf94Dn4BPmYVBkEEdWiy9rOQAbc
GI7Pjgvn0xj+yT0q4QllQKNx+9Ap0FvWUf+ys/FOGmHIwo43kcVPlZa5aav2ZyRAWGQ76ukKqQvF
OrBeo1bPc33mRsEVQa4YZ34QCKlmGuIT/PpTuPotcJ+LuocvTQxUf6bx4eY6u9YjWQNEDxRg/m+Y
PH1cPYQD9cRMullQpmtCZJRQyJRPzRxvbHyrTLH1gHdpzmWFoWuwfKlZlxuKvEjzizME30bGCBJ+
0kz1ytu0xv1Pi/jbtmEAPrWtm86sEiDqO4BrBbcRc9hsyBOijLLZuRSa8z8JQRCLxIz7m0q3dQFh
GG5xrvQODuaXktgZhJ946srgp1hbW/UFRVpXRuh3XjHZR0g2QUJt4SxijwJ5KHyTRU2ETReU3/sy
4OKzWscFdO1vYens53cZK29oTD7LsPaH9nbbHjrgCb6PP9UxYuEYktk5jPIvYMypQ1dMUb1XrzYC
luQaS4OyVcR8HxWL1KVuokFv5uQifwbRHaApTCTAIm693lpDKoreaO9xze6LhBas3VLxCF4Dadge
6RteOBj00xLOhvciSTtpDiZGXAGzHhJdrT5gfAAZlLtirPIVZaQel+gAfEMKTVQdiavGT9jhP74d
sk3PLbozQ8dEXxPnIY9KNwju7o5wX2AAKauqnB7K6YwyvoFuU1UrLqlrbziNiVtqqfcoV+hc0iBR
mtn51bWgM0DJTENY3x2BAi2BzZbPEBDwxJ/mZ6QGxwrhn9E6RSOy67mPM+haCMCMy/Gqfa3FNQKU
Q8ie45MIWeLY87qFF01PDKRGCxPMLUIVrOvxB2J8Hr8g26tr+yTap4rcT1FRU4slTiqEDCMyZfTz
Y8cpKCrkPQqDmsYUwad1swkuI6DRBNue0Z6yjo9T9eUsi8m0pscmcd0ArK32H5vZUPWwB80D8We7
8UUo5enGron8OloilPWEm03ADkjYhegUHOYC++NjVBxykr00AF81gz8VBuSbTIbKhwRqHMw/ydyi
tGTvTSIT0c48+Hpo/1ATxEmpEj7fwB9FyToty5RE+jScj6tYmbBJgwihVEfzvh/bGa9E96NIMXJF
wRJ7Yf1Hstie6y+t5M5+nI5A0LWZ6aCAQM0WBpfFzRshgIDs0MspGrtwZg5s2WX7CxsrDgxxgiZ2
sBmV1Pv7yN3Wkv5pIDl07cjT24apjQCg3JatPxGRYuf4CnQcQCDUHqiv1dxNWULV2zLppIxytnCJ
m/YDrOlKvEuEj7l/mE7CcKUCF7hVBLCMHEG5caQRSfgC4jBS4KXHlcALY4dvmxPoUmvO+j0IoxuG
9JGeAK/BgTy2mui3BykSkBQlcgpYPdB2sSTErb/gkvzJkoZ/zJAY56hIvj9/aQKACXUejVrwqXHD
dOnrq4P2Ohp0+iRx18SX/bBLxE3Fy+6yfZHSYISx36sAAYKUTr5Mgxg7/slr8es42UtyppdTPFn6
2wgrvGa1a+FgTilhQpp7/cK30Lbll+fXhym92oSDVe14q4lgif9VE1Az0mt7Fbl67PYdyxfJaayw
MH08ilbAPnjU8v8OiJCWcZ5sBXKvirnuSn2uCNJAcfgZGHg8Hq6owLRBuEaNQYB5F+qAWzdGcIIm
is/SJfFvSQfBUZ8k7kISbRNeuIWRfA+Tz78DvzA/euhyvA+sQ4ecMjQz1FlrE+reF3IDCp08GQzz
muBktD5EZf0W62AW6vkP9ft33qPIXcsJh7g2GW4CQGrTflN1kHriRAH5fOKaailwXkJDCSc95s/a
46II6aEiY/gA/TXwX71xYtzhOZqwBiXMEN6UO81jGTXb9xQo1wSGq2quYbftikyn/VJiVHcKf9FT
HLSVA0oDK5tV+0mxQg5ir0uKwW/Nxzcl+tS9GOm9tLzeHa/sJNCMna279bP+qJ2IGXYxl/qRrBTH
d/vUDoeMQQZimRpOqzfQQSxAeeN3c9PemQCt2X04FP4K0dAF1AVCXaoULUSHyNz95fBaHCJ1DJ04
lct76MSpjsQWMyGE2vSJvJzxzj9oLPeGZIC4PXsNYdnjIvjidl6aiUKYlUmScCHLpDxggPBEA+LH
8CNb9BG7qtkBKMfQukU+30H+Y8reuBJRm4ea1/t9rzjAJFjtU5iTmkivAxdW4L4yo8jG05nJT9DY
sViwOLzxyzSO7kTYikjrTe7bFvlQuFqKR2YP5KEuPiYw360pp5ozuDZQSlR66JYP2es05AJv0tqS
s2aBMkleWW/wN5p6a9g4YGE88nbAQ+016aJmOPigmoaT6T42zEsDCOOW7t2KPpVqegLOfgT0Wb0G
JfSsPQdRtEGb1wYPexzbk7S8lY6WhXE278P/KeM7Kjfb1fIyqe4hmSpIEtigrh9OkmroF0qdk6wk
xNsdvMUB9fWVYCUojd2UnrmOTa/MFdCWXEzbvcnjCDZJK0FF/eghkc9Yh9f5MVdJsDkLlou1Ql62
L4DQcwa4IzDd3htbIaP/PQhrTtxX4Xm+wPIxhbGIU+qpKJus+2wu3nkZsWxHOdgYZuIHud0kxHeL
SV0ZkqesB0FDDuqbBhlKpTZ9PVSJZ8rKHPiHFG6fELJga5n60CMKuOH32h2brBiaA+z9d3Dh5k+Q
0E1DdZHfwcjSePAkFC28Gv8uxgpG6M6YBuFIIj2TG4KzzQiX+P1dkuwfVghFY9tc/8vZx/Daqd0w
4NyhtarRCMBz1W96x/Tsu7tqbfuoZZTXPYN68nwLlrag9Of5C8KV9naK3c/97FwWjq9Kh1LCsp8j
slyXpGeOvPeuPi7blq90jSKNgcnXwYum0YMbUBrm606/huandajr0OiXAv2dVM+tPYdhfExa0q2A
oF2QZ5eZEOdD6S+Jt+GoKTm5X8MWYmFDYDRJ2a0YC9K8ABq/QFf0pY+jjg0CAN3qFhnPfJYf1X/X
uPwngSOnGT49X9wYXl56t7bgtDBtrJuUvLXmPjmH+ekXoqdEV7ECjTfhxPLxrmHQPj+rkAEBG9eM
/gobFoKe7Peuf6W4BlM4bskEq1NBOPtMXFske77VxkuMGamoj0RO1IVSK2pXOOzVV3wJ5gntgZuU
2CxRXbm785vLr7qeZlTYK/ZZF4hb6oC87PRIOe7NaGl1LsHc+3uCFAFvNoaCtjwYu0NLi3L+FUIR
PgYUyNK2EMi8ZPsFaPY9n4jnOXnj+L9UGAgCifH6UZ4hSSRYlqjGX1Q7PLdp6MEGUah5zdJOLBAc
lKMxPhcjjKVFPui1anWXnZ2k3OPJ/GPkB+QI2cXP2bWat1w2REdda7m9MvK8RUv2IY34O0qG2NGd
L1mCM8+aAQF3uOiy6J+5IhkjWxn9VrtN2Z70LiiPBBiiIVifMjsfNmtFqL4FxtQJzISBMGy+dXM3
+XWKJraIJ1zfCH9SZS3LSSxUrb2H3z/j8aoUDXqcfPLYcv9Ets8Ln1Afyr8jHRsNoagF4f0uYL5B
xka/oz8/tDUY2yL/et0BARstgsfxgbK3bkCUX3wbP6zX5iH+pEKnI3ub5bv4OBaLpKld8WLYgWAh
HvpxKTLTfJ45BxzOOYQjt4p5ZxMFpwLPO11MXdN8qJm4yL64pR07ra2s5KgvrP3HDROvgKgtTwV9
8hm+Yl9H/UsGFhOBvV8t5cMYD0JpdnuFdh+fwinQxuRBKTHJZeRlTXVuEkNQKPkjFsRCqfrXpmur
1RcNzCd0eWL6CUtfm3dCaK3QiWTrMcvH756OeQotBH4/SiMU3CfTBoteOS7t07jKv59HT9NErFKW
ApfP3L2tsC7qJY2mXxQs3uOitSQpJkKo5yMrWT7xN/BWdU7oMGL7zu/JOM+f7JRaCJl5UC7UfsP3
KPnEXvfsjSg9mBYA84Xlcogim5gFoZnO1+FO2y5OoBGo7aOYdKwsDIDg+nWQeNcftRKApooliZNa
gwA4+chkJkItXSnv0EiylWEs67gGLIFECpNvL651EohqgEBP28/xdiC3BnYwRb+LjlvJ69wfYUyV
774fXTp3ROTWs9nlhYnLz8gLdf2Xj9QlmSH07hWnRdDp381OAbGKjtDhDc4zRjkZZfrst/C8C8oo
mlhXfzA90pQcdA9VJgBHhmDQnrtC8spb646PvbT5k1LcosfMZ3MT0GMIhzSA3jzIEVXtYBPsSse/
0ozaaQ0QKMG/o+6SF5VGNszYJq86n8vN/aq5IJc+7YBV8ceW5b5o+hZ09Ip8C0JTsZ3TlTvO0rkH
mEmuqA4Ro3w3RVV1V70n6wD5SuwSXq+ybInfOHBoCO686S6eA3Wzz8AHWAgZeVzy29vEgWMCnkzO
hhcv/QtyjIvO7gpU4T7jVMSvMzIB0ljyAPE9UZeuazz6wLrFV92Ij2ImvdqezRkYXe03b8qeK5jn
GK7R2XSS+Zj3z2b//jMnROtrXNVYL8um0qDpqCg3F7bXGJnc8z2s9gEoxVvnpunDGsgFyjcly5Uw
MzU6ADnDgrIkGRKiDnh/ui7RUdKzhmlADTwMafA/X2zFzQoL1TI3ZFNelAwqcehTrJqe2rkREz/J
jezRdgWeTlO/fEEAPY6/MsU/qDH8KFiee17cJ53cnCGgl+cbgExEAcaASFzSO0A/Knn3r+6VoZHs
YmkKEuhC/533JfJHKaNJ8mzIw8LXkhjzVTSGaxGfxkmlOzGkszvhaTWwmAGqGNRJOAGh8iZ4YdEd
Qk0PHIcynU4cF08uBrke0nTn0kkAcEeFETcZ54DfexqUzpCsptw0/aIvHBWl8dRpvJv/148wV0Y5
Vtc/kKQxsHOvKZ2bstYDfBP5TTviW73bxTqP0hCrjgRMSj6e5f2Xw3oklBXOe9tJtJRBfcJOQS+R
uD7R16NBL/jjCOZQYG+yWlpehMVQMW9zGZGfNqAjBGtfm6ABQmj3rV2pPgCDto/SySVQQtW+MAO9
WerMCLeKZZd7d/8c4kZdSvo4DToUdGoE8GUa0BhNBRy5o51lGg3CoB0GoYwvp28xSIdXNb28vRDf
rKy7kgBtI4fNdpZIbKOjTurQjtEAFdO1/82CC56MoG6cFRFcFu/8BzNCbVhbOJ/PlOy1+L8siT/i
g8xaTvcalDEmrcao5tMKvpRgjZx88dWDfRK55jgipzIvp7XbTRW7O9u0nS789bjXNCCoF8HoIx2y
qidthoqWsSn+BidEidLmywT9CNHryy8puL3BSAK7Sy00o9BBwJxo3lvHwPO6J+EJ/TV2HF5VrD6D
qUNAGW4lkHmZiOoVRJR0CwQV1mPEzvWksuyMu5iEUiDr4YQwpx0FyXogdJZR17azCChcVrgdF3Hx
wkrpnbDw16csFG2vKSaHLwO8d+dzM4J0Eq2HCfwRikMC/irvGMfLAPPK6wxgHeqH8kw6Ge4pH2uT
kq/R2kznjXWlZXaNxwgmt8w7lhksXUkSAJvNWcIYOcS2jxlrx4luQyqU+y4XDXDO+9itJ0OgYtOB
d/2CZosT8x5K79VPCF1uiZWRBuMsto3mQ1bOFOqCb2yQXIAxiTNlCaABo6HxaJJu5IxGEAgc4o3O
WFB36QeI/Zyhtzw2VcRknPzYHu51bmqw85noFPLDb9l7HdDZGDGwqLDV4j4p8yZU9y+CVW5gUpKB
lDsKWBxg6FhIneDHgmHCsiQpo0BMqBwGlhSP6nHFCFLd75C2MMEKHYTEGc6amJUpuscqn8iXLd6i
wO+cKaQqANQHkq2KYNWuCqWKcFEsJ+M97vata0ZeAdmc1lI6aXTDfmEpzus8sfv+uWo9/PR+pom3
kW9yft7lkv/eePrRYUy0bHEXcmAhWZ346p9lbWPd9c/0jaWq6uAG+XolmbsH8GJ+VyGfNYXAuub/
iY/Nb1JDC3TH5GXmTTje+e0CdDE3w++8OXTrACgnUJUgnBQgzVMt6KVl4pCTSCx+u4w3mfim/0NV
hZurqcg4FBishlECZdfgtjOcBEvxgTsIxfrpznkGFEPkGcC9Lb5+t/oM4iu3vAjoSg2MzzizdPCo
lFfq29mMpib87pP0YqFljcSSHTwq4yKwQ2R41ZOtVlmwEny+d0tU7SvFsxSqYjhguS1HTaMRMGXt
rN9BwCBYyUmwxvQbStmEw1HV+B1jc1QaDD81Q2GSiuVwFwOmQRCm0Lx1NSw9sa8x9n2blP+1OZ5h
HJsi9/2W3n4uxCeUh90MslLZNRvrGmAV7TGMkqZDcC780GcC9Q1W9rQNM8ytoiEdZ+7Cig2vqrGv
vLnOaA80q5yts1G9J2U3J1m3/lERSzKY8SKcjBMO8pz1IzcEj3k8dzoLZDctjUXdKWr8E9dhwMSN
0btmz1PHpneZ8UqCdu9BdnSV26CjLOPbRTnrWaTX4VHMhsc2B7iuJXEqQ/TzkSkKCxQZ1RCpd1OV
okv9MFhkPtDO46ljqKSe/mIA4l8GUpWuAjJtVCVfs/+NJnGJe0DwVxTdvIgN5/Lf27Xp+osKfwpB
qhmV4XeC8WrAxzu2Xs6ibQMqnhoEAYeru1/kVSnfLkcn3k+1sFL4iwNifcpmkMQ68R+cSNHZuRCT
rfBwJQkmLG67tADcU5VudbsOhNx5oeV0RyqY7IUvMtgavcT/y6DoKZeRpL36aniSVhCf5XJBbK8G
AKtNFwRHufRet7vcR0SVtz1zTkQZv4v3QfPyi/teMN1hIEUe7b5jKG9lt21opiRU27VFdrgkoX5J
fkjgoFHFPQIGaVqHn5xnyZAHeMCF8c+QKyJ2mh9cVPvgsAqHZ4o5DyAr5Y8UD2Y7SUjvZTQX4gSz
jWnSZnlyJ1IqZ1hTb8dYy2OXtMsoZycyN0X7QkaOpy5meI8/0pOcqgh+h8qtTVj5Nmh1xOO9ljiK
ohNd25erFq376mkuSbzj0lFcf8zg3Ch0jKGAyjjgPRa0G2G56a8ipyUUCRR4pN9ooCSlN5LPQ0uj
E9N6PwhpxcmQ84WXkPYXTuwTkS8sSHMMbY9x01xoR51JiiA5pR82TcI7kENrGZYa8VlagsRc07Ag
LSlczEVqIWkKIYlTRBAEJpjT6CqudFXvrqA/5WG3/QL6i+iFxYhpIY7X+MtdQLgJBWVScoqlatSQ
Fo0cmlHs1PmdokEgJ6CP2fSQNj1Ff2AV593leaQVep3C15hc8WflG+LhAqou3C9UeKaxF9xf3tYo
B17HQaj1ckmt3G8kLX8fsGwuICh0nT/PgdUiRGJ2NO/+fAYg1T3pc21hPlIW8Ml7gVrzNc1Wy8Kh
WMh3GOayNAAMKPEFEnNJMFNckaEkvUTuexryFyJpNCJMGNytL8v/H1a4NTjyPVmFVHverfzWPNPw
H/GbTLIQ0z45IwGYQhMhq6K1/MkUgam5RCEEyoZu8jATmWuT4g1BGQVkosM2qEF8QETJTMAQHCr6
qUPzPxbBfkA8fQmjJZRmOjfkrLol8i+N7PxMNsDxRjm6HNPvSsrJli1ZoJHeCRIXV0+9PrARF7Sf
zvtt2suEeVniRhINQ4TKURUJDmYQH3RUILCAXCJdyY4S7RoFR3LAhCAt2OAa28zSGFnEbsvQNH4/
3oPLY4AeiKnyLqPuiy7RED98lnL88FkM0IycCFBvGxwfyeAzNIycYvk+Fk+r5d+flIrX0g2PVKPJ
jRF0JGjI4xUlWNmSiqy5GhQgVYa4RT5OlVLfaHjt/oge33wJRHUUl8NrIkqRYDVgnqxSzC6oSKRt
81wiH5rg7LB9IkAq81HO+RjkuIWDCEPcDSnRhG3zIel1YgB4vu8pCdYZVhBvWCOCqBDJYmoYNhcK
23kfIwKtW/dm4NKmvVtERnhwJQcZOTExHfHRfmn8ymngLSxgKaTgRJwTAIWlGX9dKT3qZXjkKqss
vIO88jwmhzMwvsuE/nTu1NOTJpFJC87/AxZHl0ls9uDVUB/HQWD7p1kLnEe9SbCGD+/QFxKYd77I
G4YEAfOPuKppZsVweQleCpyE1heJIF/Zyew4p0V/oK7hwz2EwvOFvcLGmPd0kI1RtWDjhkptPKd5
kiByE7OIjCRQQsU9oZlpKDd5PYTjDKYMlJWxQOg3IKiHoGwaCvJ2eNfH/RGSgtVvMh+PcRBSSyQP
JoxyQx3++hgF1ziTxrE9/JRdIIx9zjNbEYm9ZWQy1P/6XWJ0qgCOvSTG40Z1jTueca5gloeCl9z2
dt+wF8+Pzzw+uLo7lHSZbkUmYEfeFmrO+TfupKz3B28ekaXSv9gAwPPWczMPwfbjoYOKZo/tMxOj
bqJPEKbT5DRyRww84Pa6MTp8AvF1dzbs6idP43jVWXsX2e//aVVusLv0X9FPxFhQ9CdI8k+1ezT/
kIFWZKRbiNos5TqgzAsSMt28D/iqU6hqRy989DSk3/mYQoxnPCjrz9hg793WE+6OZBVEWbjzVKl0
8DDS34/38+iS6D6/aL7A9v+DdZAhvcWJknGaPo7MFxuhiYnJS8vDNsRsz3NaHoeXKIz9vLQG43MV
a67jkAGBQgl5/7ZoShR7jgK83mKiUIq4RmJCtifE7rg8nxnUlJ1SSUT3y059SgxN1HQfJqLHwtY5
A+lE6fRVkSlV2eWBwmLC8RCi94nXRwlH3wIOj7gDx4mJWkD2dNSoMXxm3iCdhC7gB1mygrmn9xBe
Z1hKAqUS29RjVvk2L9NzX+G6jw5Jf4pAXDGnC6N/szi2HjlCBtO+FapcLKio5TjXLyItU/b13kvb
W12UyscYyundUAr3HrZHQ3XLXNfbgxeoIUlDMaRImvaN/MH3ukC5TmXgLAz90oUdBtSi3KKKXUKt
W4XqwkxH3LvL6npZE2t/5hSLcDD8B6xvZPv3e1qnLiD9i6xXBX4xoaj8oLDAMAPZFg9ybZI72Y3K
/kKecL3X5j4RCqrfMCEG+t2uk3bkvltUrkGaCoL9AWy8lW3CVFj9bBIEQFs8wG2C2pph58xCaArO
XcrmidLTzbsLFuy7YdaA2PcZ9ZCEZ71VFWF9hcP1OEjTvo/ILaRIE5iboIC1t8JDekp5JhW4XMYU
vUP+Rt2AZBLmkwTZCA7iP0LnJsskmpe4U8tIGn52zaAC5SQ744VhfQNOOzIpC+RCQMjjAVWbjPTB
TPYwaGuvDGM7nO3k+WKa8K86vMHQchpCteraHthUKmxA5LMY0IdJcEPwwwpC+fH7+M4UMVXwOwPb
x7v7TXjlc+mz1j5EkripMyzDhZM1YKF9bukSoU0P48CLK1T0yqzjrsD2so1MR05LvK9M7N//+ZLd
kYvBb7DRgDaPryG5svtnnY9xRcFX3jAE4tK5+RNoR2/zxx0qcJuGzcySKo3Xa/i5gs3k4C+AViV8
gcXzv0MnIBafy6mZsX7ukecYY/9lCDRZFP3kKYiAfnaE4eP9nQipWFsufRH9G425IE8VH3hkjuLR
4VX6uMD6fvDEooIJYx7EhKsE/SHnoDc3wqLxAlai6rPofTJzfgLtcVmG9EhqD1RrpL7r0gZ5BMxT
f3/CXymctFASDeopSuNBFuo8F7SLlAOKcv9fWlPlqE4IeHBUgWMjDpPc4TcvX1gdC6WNEfseoJ0i
pqGBDCDZursbn+2ULpmG+gIvPg90zZc93tQ3KoF6Y/sgc783wnwSU+774pPY58JpxAjGQOE/MFHL
TzdQILUVE+YfSS5nSBtf9ZTjB4F1u/NpVDHg6OOxXsxOMktpH7oM2z3iXcjYIfcS4MXclXsTkYij
gJJgX13+g98ZJm0I2Ewm1Uos3eckyfise/zx+KUDVkx6cDgEXGNdmZCvLk4PHMF5ZdfxSBrwYvF0
Qz2hhYMmucPdwuGI6BlfDTbrVNHMXOpL2Qpa51E7OaW8LRVjQTx/3O24NJLdi8KEqGUu/nWHP1Xp
iLm/Diz6GUL/SYFW3qzC4amiAH7cv77YaUy/UmHw3EMZJvS1tBNctsPUjTsvmlg/ENQw7lvirReh
3+HfQvVkraq/hq/0KsmOg/e26OrA4eGAgyOZom+A5gFFKnq9uldXid4AMGwBw+RuOFKwsWsO+HGO
jAMGYMLwmwdy6cOWKMEPziR3Cm7VgS1xJw3isC64IAPJ8lisVF0cPNtvrx1iOZcqlXUkJoccYu8y
fU5vL09TI9ELS9+qQFIJX0O72R+XUkEViZcfJE7LcYp4gU/X91Kh6o8LErHLZBIjguoKz82oEZ46
JuYF6S/Fh8n6N63e9EDNk9CwlliLOgv65XEL9vif33kW4QvyB7HvycPRqcrj0v/XGXD7JYTUCSaH
SZ7APY2pO5+/asF3Qht+3eB0yFJKEYHIkKtzeZCgYs1YdzrsQAqlsSta+/8tfa3hGWK55PRI6epu
xoH4Amc04PXZDMt/Kub9qndm6W0Ye1LDQnGTXNMwjbQMWMU67pxQ+eDM2M99sFnXm8mRPW1d3sSi
+9hghZXXXSCUjT+INMrJ7cfKMoAAYber5iZSzOMo1SPnPJY/L6VN8Ne2PpZ4k8OokQudZikIt0J+
g6ho/JWkPBOuBdVToi5cfUgOvYzBLuU1jjsne3nx9b5wKR6UYm1GyR7rFOx553F3MgYJNvkg1qS1
pPTV1b7XTtrd7FfDZ6oE14NIacLmQ9q6g2DnyjHAXcoO0F9AaqsP3s6hEUbxNganSOvToikx5UD5
GagGzk8JEkt90w7KTgcIYd4x4knhNCAtutEt7SD1xGJnXpSZOCketzI8HfN25OdQrpF7babGwHF1
21YS/DE2/1gI7vc1GIlYOUt+3ajoUxCL25/gfBdh2qIQDer7gWKkT29toDWGKoN1Rh9H+70va30C
/aIcMim9ijsiuuGAXFSn8+y4GfjiRQFJLwjRQ1jzOIFwBkRZmtd3g9tI/fbW5ybo0XeRZjvatFZo
B5ATo6dmrslewhvJe0hI08Br1wHnf+lZGVqrmY2rn5AqeSFmfF3Nl4veLu+8ARjPVE2G3/mTx4gZ
MGRN8Cd6Fy9ZG/wor0hNCz8XKFePGhCqRMSVidSxP0yIN/yzacYMGv9Zaqr7RDAh5J3xT0OKOgQ6
KpdGRy8r1G0eig5qBUPdbss1RDNEsr75IGCJ64KkeVERf1ygPJlSStDp7PdUOdk0y+yfaUt3MBh2
pKHSTOopiyLAd3yQ/ADrI958b+xcoM9TGSWObr+XVKWoeiZggmwRnSLY3iqb1SYmuAUw8BTfywK7
jv0p1HzlgNqKgU8nxgaNJ8wPy0SXnRn66Vxi9eE57sN3RWeuQluBLpyWZr9hKVuQ6p4MwwCHS+Ae
FKb46CgH5v84HSH6f334XwmE15UNA5kEkFaLUMlz0hANOjzMQjBuL4WjvBq4NC6PW6NIQFX6g7lQ
sec4Df/MlBRMkwmTDy0/cQGvecPEcwReMK5s+7dqCIiVilzFYXh2H0KFRe+VZKxymjg9Nv1+n7Ca
2xaM+dsLCuGMgcmXdmflcTLzR+tp5MI5xLyiP6wOCh9QTVYj5748+Bye0JCtm0+IMCW9HPJezUYs
okgPe+611lmTff0MzNN7lK9EI3k2dePj4GHIalOrmj3Wf+kpj8rnX9V7xqYp8Ub/8IAoCFnoNzgG
gZ+S5hFavII3umjLhb3WZKRLFGAsXZB8RvTWep+r8EP61ezEuFTI0Yp5wk/H0N4jgR6jS/9sSDmm
KeLmWaFTnuGBcCFVhZYaHoG+SZGQFYKwmtE9F+Z5CFv86p5EUzIJmHF59PEhR87KKC0qF7zu3aB/
Q1xvfv7ddF0rLrJcMrz0tsa63zq6F4JjKF1y751yapsvrbqvVcMbMPiV6OEthf8m3e+a8bDUb3I/
bc9LDAaS2rGGOzTKgFbhdT3MIKg9YX/Z6eZhMJr6NIH6D3OAv+9EJ8nkAQ4dKaiLTiCiUi8/AWTu
3Rn9ZAfrtLNVj8cx9YdD5DNH1cjZZ2vae4m8BCZj+JxepncQ6XWLTvT/F9R9J02URk4YtY+UmiIJ
pyBzXgyEBdqqSgTsNhO8DLFi3p3m3K+jlejJeskDOvw25CYBHG0x+9Jnzfpk00Fz0lV9+LT77YP9
RalL1P7rdbpjKBqoSO+IwJgGrfcHDALlAnsDkmKH2PlZLCdl1F7Zdcd4JYJURX1D7YLpFPtUUL6Z
AXpXNBtEPqKAvN6nK4dQIq4lZt/cqryQf0OTAZ5JBeyhwcuD0yArTxWQNjCOqFyIVYVP0sfyx3nO
YQLq+LmKrtFqFBE0WeCmgPtPSGbc547Luf2FZWQ1jAF1zP7EnObyRrRprQh/uZo44hrV7S3X+Zbx
N/xLpedjrxpI/LhAnm6RouSCDyfpeS50LSwPU6WQgyQy07J1L9lGw8WBEXz4qQrfy7Id4H0amaIF
AiVy6ncBnZUkUY7Nqzny6wHYj0KWXCFU9u6d6G9zyWWPAfEdmy/XXpg1B99NJUdMQfW+MCzaqUum
b4UveqZIErSL/fNVpuWOSA9le2XrtmV9SgCpjyflt9rqU/PQiSjS6qJK2Kj6CWE39rVJt7I86N8s
bW05DSbY11x//yW2a7kkPhsHAZLhB3LnPHtX8wk4LcsIIdo3iO05fQ4jqEwvPSnzp8uleG3MIHgW
qq8FBEL9nf57BgyvHqdRRhhfz7CttZ5axyKA708C2Qs15sZ8kIFfU8ISY90D0+MnVojAQqoCO0yx
WROYm5fauTe9EUv90hMYvuOYZgGRDJp6mpFkFMdJVY96mJqmW0QNIcHVH1xHlE61RLvWUNfT/Qwb
3qLNqGwf+glm4IZygoj5nTx5jEqjJod7RnQNCg3runBO5MUz7s3a1FE7fOhaLo29Kd8+IRX62ehl
b88AhgX1R+uMNDIqD2Vas+GzwmTy4pbZRK3guqG4+28VOEnxOqVDqGHtZkdsHT7dLMqMlfXMWrJb
ZW2NfcM/yo6kK0yb8ayW+wvotFgSGc8Wm9DJR9GMrV4A7DYLn/dfW69Hd6Wjp6ppwh4JtHE74CgH
2RiYQtJwdjY712sDQoK4iNy7YabcNEu6JMGNoo6CfFdMY/VQ4dCJ+HrWKoE36wk8ivPueeKHHVyk
aMamu3zrD/2Vrpr1f9m5JK1H4svDmGJ+y01n3qie0lwcap4wYdyDYxmNMTEPWvfmmIUX/M6sir/+
tDORHs/f8TGdJzPD7i+5ESIGl3pkFRqRxiDzo/vzPyopHYf7UX82iQVa3cMcb5pwxMj56xrXVeDO
SusmmacOejA5NGq1g3+bV4VEq9WaHGa9yLkxNg/wtnZ9fF8w23IDnsXGGHgIVpHKKdbLZ5eyI0jA
oBht+C92EskDibOiJrANsq3xDKp0c9KjI+Fk+n9J4SHOXJBhR3s12UMgBSNAsq0r5bGV3EB+BTns
7J74wzMDI0yFNAMlxWiqkQl6J1WTmnX8YRtqtHYIuLMiviiZq8MyXDzRtbpAx2kD9MdA2t6TulKk
Yvn196wwfZDIFcyGg9d7LhJNyY5eoVtxn0rFmBk/Icl2vh26/qRStxBgBywqNcyyGaT87hTIkPuG
JCF8/c/+s9F1SyfzvT9dfkVHlJamIPtZjM4vf+nt7YZsiQgzdYvtMvYm+ICpcAuAZXlDJ8i2zCos
qmrJAuOIcq++6amOE1KHXbtUN++BXMZ8zYnq+fatjSjfNU+yWUZW5WHEer4idpMJX3SB4xyAUjhr
3YXvZ2JZrJZ2rYaqt+s2AImSgHB11aWrGxPzGJYbLVI9pOqIIDPLGY99SwCYousjSy8nQSJ8UlO6
9GcxJe6HFXn8RPywDMDMdcZbszDnl13ONV8C4dwR2tgBUpAL5IKEoa6P0hwNgIFvkvr21s15KbzR
C/oJ85JRxI1w7BI3DLEmTpInRzj8kOrLai2LooOCmo2W7SpfKqHea5Kmvt4v5jo6Ch9FoydBEwLb
HpFd4vfwdaRmE5TSsl54EEQ0uLcWWH9nPz8DEckPRjeiNIUZgTOJ+SorsPYAn4VEFX3xOhjM9KtH
cjNrXDSxRPrVMR6epHK8L5BSX4Y9Jjx/amuZDl4whV6259o52Eb6dL9b1LltaCQye3MMAPNOqzT6
rH4pSfR5v+wK34TQacwHPUauLYrbwXHGx7gI4Ahj2wcnGOuIU52IjwZ9pFsZcwOf9TlCaMaakmzw
DPyPBzmTDxkkxchvZCKdJtUjxR3Kss5iMFSdBYlJk/B3LEm74crrqBshBpe/CCa53HHmCS1Hssqk
xW5CvfvEF6oA02v4rZc/Sf0km40THCj32D9sdFk6NTcdO3m1SbdbYisxPjvhQ28yPc+J+S1FsyWa
51wlHjCjDAuor1DCXkw5j7rRfAdSXXqdoIN2TZVmQZdXNKv3ihLivtW8NrUUG0RYV7pfXlkuZFal
aRLCdpnUvZzm151RlSkeUyvwkQsUL26yVht0PEK0Jo38hTOG7xY0t/9/KPrrwHewzPMGL8uP+exn
E37FFIx5iGO4gMmbeIS6ih7zCLIs+B2/YUmtf1pQsUwmIa6+wmvXblKAH0k3sLvI7DQ0g4h1fwBm
pqViPOeW/HTI17p2doLRcuFvyPUDRkUspGl/nKwCNZkcoId7nZtJR9FNgnfupwkxZUyuryVZaTJd
EgtiGobrN+yn1OfMpOpogXeMu7EM4RCyMnO+WEIbIdCBuEyucyRf89o4jvVSkHDhZjZwLOhrUKAF
FnP8YjLAvZ6Vn7oE0a/vaZ/OixCpby+K7sQTwa+v/3L8MLnnYWP2lN9RqjboLlHxf8ofOf0pEmos
J2zHa1lJE+ZzswHfEK1VPbfv0tNEeJvI5D2EMeUUSn6FZA4MsnhC1IS9oeAkz0yXSYxwdbzUKr5t
CgIliIJNJFuY2m34QpJkaFE3wZH98emFXxRsWFeuzy/0JlWPRUDKDblKk2pabzWaIi32eBEY1xgl
tpeAUOL4SfFE+ATYsVxBsdG6MCB65I59l6WVxZNJxBZRDXRwxJPuQVyzpMXCZ46fl1Ll2vtDOJ26
3PqRIONKvl95ptvQP9Oam2I9v8lWyohyKg4zU606bsIcslGAmnkI0aveHDyRzRXDs27Ct7tagphm
mny6f+rN2WHv16oq77KdM5T3F2r4qbgK0tHs7N8PtBawnXBb2CC+fOaIP2AM0/ZXL+atHt/1CYTJ
6Ue1Ww9qo1uIYQyQkqUTzL6WXafQCJCfIxe50E+KDfbqPlmjnAwXGPLTV6NLAhPTdi331H6PL0MM
gpSPjb5erMrLKvbsS0uSuk7TKD3LAF3dLRpngRhh89W7kb5q9wR/DW36yi5r3rhvmtz+BZ4LPNqh
MoyYuXgF4Eh5Xe5a0clIgh1wRIc72JxvNCUxMatuNLsFwP5Pg8AnYlrQeG1BOKKG4NC5qAeIgOT6
FCH49AoCC0Dm29zoy4qOGI8AQg43z8CTyAlSreXDx5pfC2gaXOm8xqh2CimGzj0/Up0huJEyY+HW
l+/MF2qIIcgNUYG3jQDsXvvkoz1w77FxkxINlqyEHJl1i0q42aPxwtwTTPl7hwzfEQKU4F3tZo35
YngpUCmcoQyA6QjHEdZPY8nzRra394a7OyRCzIAfQWa6Ko0TugIcHESRzFb+p5i7HJPbUMeeCCq5
TdE8kbB7d3rm6rtFh2yO037sk5rNazOb1e8LE+FY8Y535M5vDK//wOEX/NdpT0DJ/pkj38aBUMEq
PLItqKzQjd4RgR/9ZBP0MVysM4Ap83vGVOFr9niDqosktkTpuICMvxbVNipDViU2PooXsI6LCl+s
YRTJO/09WC8jBo1/9AflagzlOdNxswj+3rX7nrnNobPYvmfPGL67ByfXIgAYtpWIUskh7LzcxdhD
Bq007RN+KFafKRpm9GGKptYvpgVmZWe6yvnKfCSMfg1HxvyEAQxlH8jVVYLNvZ046mo7SMjzeHmJ
iW0aWcqg76q8HWnFFjcZ1t5i9mW8JHmnHmgqVtO7rlimh1Awu7KkszR9dF04vNMVsDimkME16no4
SwRgdWORmYSxKEptQ80zRIExnKmhEQzF02TpNkWVi20sEE0bWNs2xlVpFEVnTbjRPOFQioT0Ju5M
hgtlzQt59z13DueV+9DGIkFpQKzTFnjNN+lkK76iNkOiR+nso1q2pwzEsMINm25hHEoMw79npVKY
TwWFIXWQEIMKyKUrtyngGzN2gGC/IDlZkbOUOkaKp6s+gSzDsd33shSfZefuwVBpz6B9Ea1oSBgH
lq8u94BV995ngpfasqt0sq0SSkInw1+WQOhXtyutXpyhLrQbOOTo7HYtWi6yqq+2TeuGqRLmOeEV
ZuSQd1Wr3ZTKR4/eoyhjOfgMz0G85I9S9yGkue2r8GDK+U2JeiZ6yUiMaUnsSvGLdhVw8codz801
lpuka4Ss25tgvlVv4N6tWRFYbIMfqIYPbncaxjkVAzfdqdwueh9nZkVAjGhh3pJJzsymSj6mTCRb
EMO8cj9UM2jzHssbee4WosNjWc7ejaWbyoyl3oARZYHrwi2I4duggeefObyUKipLhHYBLwss33/I
+9p2Y8J/YKhwxri/F/R6/aH+6skluOcdBXZcWMSX0cJms1WcUkHETjwywGPnMh4ybZec0w3OvgUd
sQLJZQlv5pJluDUTArz4y09XbUdQ/fzlq2VHt/BwG1/Mc0bx+gizS2Vps9vnHyl/pOQz6ZkBE3gj
BAD2CD5ZzfMMkZ269J3C3AsngwmdhzciMVuSoiDjqp5H7IHgPc6os70R7eNw+fci7dyvfXLSVOeO
WKfIepWV0r1Rjx7n6qa9WKPIaZTbcO9x0VMKONZ/NVtjpK3vb7wEAI4AzHFcGUxTWkKCD763muqW
apTLzvImUD7wmZlT64igEOyvo/mNHAkCzZIJ4ggUVxpdM0YvEI77Ibo6W8nME6bZUImXlvenkfvj
318G05XteHokHsmPq5O+2D1vN4SnH2bRmLok26zJBi+rZLdtGxjkXePjKIwi1AbXP5tuNDlLIHAx
kpVq60RvLiy9UUbhYAvHPpQntpL4H2SZ6m+SoGkDvpUEnpPVTRu6c8BuuCXK1TW1N8KLxAXLWcPr
nTzXNe3hDtR1CoQ3RMDQ8hm+PXT2gBkt1uSu+/wAMMOVWY9k8U5QQX3rJqvYN32MQlUswftsEBJe
7X+Nk6GRmgn4H+J0zQ9SbXD9C+fJG0pO+59CH+/bIof32IaiBjkDJz5ZL1G7iO7+UNlc10w4WaWt
Y+QKIiZnmnySYCnKczHR/R0FYlWemohkVas9J53aQG0eWVmf+d9O5MrM9ZrSrcUOGmwvRxQAbj0l
JyquddciRmGyWPo2Xu0ZYKhH1N52yXIlkOpF3iSv8iNzSkXOY4uqaHYbsJ+Q5Orv84V5ghG2oDbg
iDFaHlOmweVKw1jAj95kV4bo37Qhgv037RTaDqO1ZYU7ozZ2fjA8fsc2bKDKfuXhhDRtjMc/KsmZ
aNEmK0cInU3uuuFCpQAmcTQ0/g/rRmYZqy2wN7osj3+tVfgPG6vJBIgpkwrJXz74+/OwkSh3X+nl
aPnUZtHA6gmMTwZuyI6JRQ/ufmGVx41iTLpqGb90NVTczh1penx4qSLtHEGO1xLID8LPCczOzbmc
4On5XbkHzDjDjLDbjoxdbIZX0lTKDFod09NUthsSLeDF5tYHJPkzRvE+1rwvfD2yN/90L8ppm68j
BtkhojYLLt6QcNocKfRMvUNpfxJo17SeCPuEhozqU+OGyaSAWgmoJXznvS5TJSyVEugFQKvPfi/p
P0bgWVd0NMAnN+B//xrF7EpaE29rCmtMQpSxzMDpCFQxVaY4nkFSUV3SyfBIuY93X+ShTGWjtNk/
0SCLdgNf/3h1M6UeS8AgbDW8iFQ0e1vnAVgsyiUTDCSfyMJpVlqqJCCeTq//A3be2droz9+ogkBO
sElWB1djyS00EaXk+GeX+GZrvTTRWw2S7tN1iZCWd2AdNmBQ0WVwyjydQ7I2mniHHnCXpK2FTU+F
JlXBKms6eeJsLUQpFOMXXUDZXkEWsaBHz2JW1ukcQxMbIWJZc2PRnFZX/8aHgZC23/2ZbIUNBRF8
eeLXxhdabIA/NspLMUPXCuiNFT5Jrzxfli7FmQzAJTlFnqH61Gj8KkAi8ov6abK/LNHmYCESLe5g
3i6yp0ZSpJ+5gY4bGoMUtJ/jkktDzKD4WtAXN+oaDflZobkASuYn3nYUSwx/DpIVYs6/s+sx0kqv
2gr8y1A69aKmgj7Hyccelur9M/1knauuhfn7ZPiu+mNAW5+GqKANulIImzxsLGljNK1XrKGZXZB/
f9wgb8O5gTUUpk2isjybnBx5dxJGOAllJt0Qx5e5B5+XPE8gZ0EbZ0saOgwAiOzWbUc784d2MRF0
z32j7+co0bNgzRPA66IcvTAyWlBiqlF5lYGDcM9dziePrqIZ+2ebNTnvB0gOw3rR70cVGQRIwB4y
Q8DZAQxlSlRywBw06AU6RPcvQylfqY604jNIUIAboWlb4uFts9tdQs6365Y5CvW4oyR58899QAtu
ifNHNpQbfuiGlHk7LI1Gs+t28DHfgjo43jXKA2bWfq2sXCYAEyE/ZVuRBHqH/xHF94lHwDq3ppqf
j175vuil7RU8kGEC3Q+NyNPs81xyV6qquO9QyaIFjOW9bx0A5Ern41m5UmPi3zccajpcQKVP6uQX
GVmOQlnYZ3ZbcjMxkJ7XkaFSOCmGCmalmgeHJ8S0sEpkAACFkg8ArqxGC+e1I8oCSUjQQSZ0t9z0
vg3iB0SBDccUfS0z0dCCyKOJ2UU3f/rYQDODD6onaxCgWR+1NwDvzdf91t+yjE5+mlmmvibPZc73
b01KjuKJ9y3bg5v2tXgLza16/6wGc18HS8J/uxyTZl7Wk1Hu2icv/ql/RJfC6jDycpKcsPig+oxf
UawRAX2hib864Qa6XcUJQICIK/UzaMMOdTLfKgPonq2MA8GRDE9a5OekemcbKQNymgEcXq9J58du
pZph1wqYNVbUk+SNhUXcF1vr1BeNwDYHKznjIDRD2LOf7H/dRp5osB0JZkXWGCr331Wg4en9qNiP
RHEs5I8LghApcu017VfVmIF4tWBMvdNXFLqOZ0KTjDpurrqwBcXLlXCLuKsql3QGVP+blz43ZCV4
uDVT4lEeR2FMRYUJPsdt2lCyoz7x5Y+XjoLjd1IY+EpzAHuDoqTOAdj33vLh6Mm4duaWlMR4pbHY
yJQr8vPhJpRXl7CDYfclvPV7ODL2JkXcjDX/E54l1uj9M5j6pC6X7cGlThjPlPdA5ktICmkGThDi
pvmPQPKG9q3VTRQLUO3TNQNrM04gUrdsfQHuC2I6PQVIVuTUrpz1nIMiFs6YNJpuGRWKSUN7LGdZ
5xtookesxDZe6YZbxeyIZgdDCbHNLn9pYli9hz+xqLOUmCZv0D2uma3Zpb/uZ6ozNPvyFjgf0lao
HXyj2qBiocH3Nq11Jgh5kVJylpktKmh3p/Md/BKqSDQB4R4n8v6uS/zopL4yn/Ap6YSowqfQyghn
UxweRp4EMB+OpDXdRN+54S/kEYwjntdeaF8hZtZVmLuNeyo56nuVWIe/vbCKTuCT0Mo/jnaC3Fg0
WUCzypqH/WTEldAPfKaT6y9hzfX8zF1JLMYMwPXaGJEdt4p6RaIMZb13A+ynw9iB9HfaO5oHt9Qz
iDyqkYla3ksvg0BVYNFAuawY3ZwpHOKNoDuL5fahjKVz5qscQF558YsrYQ0Od+TeIKjhOFYDGQ+O
KkxazxaYMDMgTRQpG5vjs4vsYRkII17jUyd310VvAwd+8JKNTzoKVWm+qiNlYL1NDnamKCEewfFy
bZn5q0qMKm9iqe37eu37zuWk6epSvHsodUHYWurotfQLYZMzakB89wnzM8WHUVCskrt0o5C+X4Lm
oSeya8eNN4Qb/B8eVr90IVM/VszTVNheVaVe1ZLRYvOE6+IwILHzVR3tlwSaG6L+YpTI8Idaldqk
9qdzpBsALWoFvHmZ6w+4zEbKzcpCh6WqEnxbsdiop8sVqHs3CLBu65T1YVzOsIucTxvAHKpbIkLO
GFZyuD2FiJuKZAhJz38LVCHo0owr5PereP0Hj4cWdEUmIn8YppZXChTfqlyVjw0Pgv26KrTTnT2x
ntRVL0xjhdQVswCnMfhdGj9FZjbrf7eqApufQkKKBsoiy4WozCD6Teo+vhoVjMR9vrzCs3JzcUbf
Yqb+uvylTaQ7EWKd7BhJbTsGWRg5VmIY8Khu6OTUDVvk5sEaAFlBJppEJ+LCxSXZadm6xfSGfTt9
r6P7361J4YxNk4FK+RDOnrn4InVO8rSc1hUBFq8tDG96qwOI5m1Dq/dOVUa8Ro6Mmh3Zr58VkUWp
tylYgskvCrw7NYHSZBISdR4vysyuKweW2MuhqF2Ji5GfeIQYeqQ0Mk1UrAFROmCaGMCA8aDPtFu8
XUjJVgj1Gf9K/EVg8MP08A6npbu32lkJV+AeBO9Y+G7fAz9pHZ/cnAohX/8XIQPdL/GSyOYkBHJH
h76Sv3KdIvEwv4YBqXsIcx+W/c/Zo+/uvXXgMWg47cG61c6vIWNW0qOa+XeX32+CHnx9+6ai2f17
4YBIAXrNBVE4P+PvuzP4JKNZTvw9CsBuojpzzV4HVbaf84CWS7Cv1EAuItFlURpD/YcZq2uqsOB3
j4gmIulatzX8eRnRvxQJb91iyOGPUpvm0W1flcKBh73g7Xn0rhEn+8AgGRkIWaVqeOhQ4PIXiPB0
FIacqFe/8To/T5zvwTLWWfwmW27xj4FLx0awroEdDkn+j4d+OY+/TyGsp8dwr4VZG/q1iOSfFxfH
gib2zf4NdQeKufFShTULYEZ61ayZERjAO7ujayqLdQ8t4moJQc89AIhSoOundtJF1XXn4x85iitb
7FrXVOukkWNezipVcL85eHb+I5xYbV3NU3xJ2HVt+wkA1o7iXtkN9OzQLQ1TKT7/a/CYsU4ATPc2
GboBVgI5IaTetDeq0j/ONmPmTASOImsVpLxUiNLwo9JqnV77owrJ1x2auESWDY3z1WsqlcHocsYq
Nun/cwIdKoNWAzZBgun5NBk+fH0/Z5BLtDnYh2csnNg8f9vOlTHydLxDfV5NCFrVYm5ModgAIj8k
UWo+1XB73wPUFauua+12ZEtQXHxkLZeZQFVd4HrmM8uDdJ8r4lkWGd+PETOYFF0w6gsODceQWRzU
IuMakxn6TMdzZGB4t5xMyZoavwGwg+HKnQb5iDd6qHntOuApIudmzMeQNTNzqZBG50KEQlHoBv6o
670h3v8oh1CmMoCB/r4xaJvYf+UupZtadTymU/QQR5Y/eXiJcW3mnRvWJPxLqgSVyG5453zsr9fL
+reecYWsblNOLYnYEm3wcl1/Q+CeFMhx02wUmqOBW7PhXByqQFSGH7I4yZk+j9TFQi2n+ZSo1qGc
lBGCWfqTNGBeoIhap9e98HBrceKKwpCcewzslCCIPSqpZat34HRuwahXZJ0fiO5LQK5mKoO3fz+I
oVlCxtr25lokOpC5H8KmO6UbzufsxC7orRBjEM0ahNFrWcfeCefQ0Za9+2WYcq2f0yd47WqlRus1
1lElohsA5kUc/oRydmWqlQV/uh/04K1fwu4aAjIhax0+1fdFyllPKbtPfPZXZMQFn40c9hFbavdd
7qGFVnKiHC5tsjAnY9NABSVcaFcNZeHcp+5NHwSIHinCTEU4hbQqIWXqx84Z5bD4pHSzmqVB6sRC
Ce3T/GhYBeu8YWwdewPMao26kjtBOkjvbZjTHmHtG4CaGcBHwSeP4XFJ4QHZ1S6LwSFa/k58c8id
3qbipDC+QPjXfeWBLW7LsN0MClqMQGBBFj/ygc+Y1Wcuf2SR6elP80vCUc37+XILJiKPegl9hPMH
zQxLO6aEhqFCqekxRp2foJOiKFvZAWdgVCcIQktaRK3DQQ/nk7eye55pyRXu7mLw6daifGAnAWn3
SUJfisKGyvn/85oftMA78bERb+0YydX/T3ukJvdEG3dxTMungIm4C9Rb/TY6hAwMOL76BjFUmeND
V5loiDhMG/3QuWczq/sQGBssCP5RmluzCJHP6JIDunt+tz5/0vKOncb0EWBF76NLcl6x2vNnCxqE
Y1sW5AvJpKWCVdN/03/sfQWZWud3CK4shoW4O81m8DyTO1hpCn3ol8bdl7xgnuyIQrNPmmJgd+tI
0QmtvkpF7s+ze8qBEzCQ8T1PViN/Ug3jLXEYioMqB8bGZlCQn/TzG8Y8tt0CdUCi6Y9wSd3ddSjS
UTGC7YwtK+b6qyPr2D9Z6RyNl1Ns66lQWcfhClp+X4P+iAoaPN+9WOmK6CtSJJQvx5jbnOWkE24K
DkZOK6eMswRUQBeUzmgE4NYa8WoHBODH5LwVY73HTFeOZa5Je14t7Of2BNW2Ty/utrr/X5uUI22X
L4V/2wepWJPcIQUA2NAPuvsaovAJ9TpjdKpQ9vpWNnOCPIcguZanxdwsjQhEtLw3/9VZRyNkrw49
e4JBgAu8LD6e5DPULQ2c/YvOCUio665zfVsmlZ2IleqGU3vK9EMQIm3vgAqJ/vLHSp0O0gWQLAYO
edeTrP+8N2h6ge7o6sv3rx74Ut4Z2ONqYq0jj9rep49Bv5s+C8rYiA9sJ+/wbv1F9wCccDMDazpI
WIuDdbn6Lv+caQYiQmhIR+dyzwcN1xm0cY7KtTvNqbIdapJcGgIEEa/vLfDJB4Y6e7fNGrFE7+I8
jW9iZFzgqldAajCUfZQVC6lUkAPN3s1UcGdhk+2xb5vLtpzX+C7cbMU1KwtccE49HzfXsEcrn30a
FUEJoYkxKEwoF1dcqlhvhQLAenqOvfpN2jjvf5aUJO8YlBqinP859MtcZp5jTy1jNcf/pBTDdIYP
21VWTwalZoH1T7HDBA4uQ1ggDoGMxECac8k2A9ZxBPGqTRMxKbhi4B1WCyFnSvifhmsjxAc7W1+j
+SUjfzSWGfZWxgQybFt4evoP85mQVnm7N7mmi+cIzLQBOLMxLER7laeKf+sv7ATKreb5wn3yVv6Q
7zsqeVZBB7p1zC3xSyCennxoL6Wa4ZuJFhrAdFsL/uM0pD2gRRChqoIpd9AG3AJCtBHg7tAtStL5
24pG2DV2p46fIgac8ZuoBzpxQothJYnKA0o8feZirvAxoq+ZNErDypvGxTWwdRk0BpWh9/xgn9R9
ApGaz3eXKD1Yb5oJ6kg1qLiWlIG7/Gw/JZ5Rm/pqeigmcsSd42mvEcylc3aUdQuhqCyzsOADPes/
H7Muqo4NyJw9+FfBEPPpBIvjOiMqOVFuXsbaMxycHcXXjq9EikDnFMtGfSrk1g8cV3bAPD25jFi/
pTj5cS+6Yo7+9pUF51cNxqM2nKQMsw+2Smy8bopKxrjNwipfyMi2F+8qIMHobpg6YsbPxrzyOlgT
CjADNkv5cc4Um4qj7VNIJVfRVwwpW7ZvE4/e61q/M7YgY6gsrmt2FeNe3x53gaBRBqFCkeO0/JkG
2JxF5t9hKQXEwRNRSU5kK0faQSk5CAEXVrmZO6IamVIGPMaYIyJG99Ms6DDQ0nq7+iZ9uTG3lbEg
gy9eTP9Qe2hZrKQcFF9uHXnLMYJlJ6HqYmLbXmMNZ+S10EqJO0SBNXjiWKZWwMUP3GjyOzHWHb9q
gMszXSbb5KQRQL1Zvc+eK6biBIT133K+0MBZJEnzZ2khe1/XkBCAmNATlYtGAimYermaCywc0BtL
qb37HQlhkQxsZMzgNZEGNQnJsriBLwVtNAZuaxpzp4aN7KtI37R/mBwlb+F7/fRE42MvrnFjzTdO
E9Gs5guUCoxqgbegwd+JvQWmEUIevtIhUnL5jHSgD0rxxJH85XcgloIsnVOPos9WsFdRSaSMZZN6
BNWNdP9assGie/HrLbcI+BdGwkZuxtb2gl/RTgo1hsTE4B25fi6KBQp/Z09jko2GN3Jg0M8K8f8p
MWN3l7GSaTO3lMo9XArjqd+Lf/ZPQUdW0l5LTsh5zILH1bQoZ3osSbIVCPKK+Ex6aPze286/SHaL
wsd8Oscdjq1PbG6oScXcQR0mraLjNJPr1Omu2ptIg+kCFJc+NGq1vDKLifzlPuRjyG2Csq+q2wNA
vpc5gjXCMOK6kWaGgw5Oe/9BwBjPbZZ3JSD9u6dYOdykUHTF4vyJcSowOh1MEpO6oul8TlnlrXRG
flS3Z6vZWu9XbstPQebcJiJNoyV9uRSAalKawviltDCgGki5XtxCOU01xsrroUfv5RZ/Th6dFJVp
1Ms2/ysxvO7HvIH8VVBD3ILQaN7pCpgbZcT52QHIqt9qzndElH29/Y3DPHvgGn5+krUkdUaqBM+D
+VRvTCmeNeFCdVATKcTBrJZ9QZ2dhikuFYnIJ/rI017ohBIEurW+7pbhPGo7xVAh3BsLYfElkwA3
x2PuoHMEVGR0705O5+eaY+LkN1/W0IIj4crUjabioGKdd18ETVPQAQltFJPXWo+eKK/rapIw4g7g
k3jDz+4nBMmY+oMOi5rLwEDlWvYDwSxmLuLx6LLdKTiGP7nTTibvUW2e0MFF4bdddFt6TLfeavLH
LNVVnt5tkaH0r7ATHWuHdhirWDu0IuQrqSX5NAHEMOkFaZYDC5IG8uasjNRoy89iBLyhYpMGDdre
8/80carISJ0nSlthZTZPoc24x8Q6vzt69bQgPYQtWKRzIrqRyqK5iWp2xWplKgNwtJBLpmECfu+h
5iUV3aWOcx2aXUXN5PAQCORVglsooAYTZES2SiPUyQtCQRC4BFS1MEhEKgU73CMC6vrZryCrRVoI
9ko8GZSu0o7iv5P1U1JVR5xongbxOHjsNaXNWLbX0kS0Zm5r5CsoiVNbIFD54gq1ob2Chiqu3seb
r8ZuhdGgUkbt9uYXMfzUEv3zoiWQmjkM8ZgD6WEZbgBou3C4aNkUAoeTRZLzU1aLSWzu5U76fLnG
GW66PjCLg06FxAyXy8VRzDkfG6K25LZ/v9oSqK1O8uTcCJOEr71Q+uxqfkYAXDmuc9cMBUr83hyu
GCxgEG9XcGfttADTIrH+CNeRbqHAmH1sdFCtaqO9hKYxbGdK5fuhT9nYY947grSCUcYgm1VNEruB
MwGKTgwKYCyMDqxm7GZ/ouw7Di4o1ZCUUAczTb0jNBg6Brm0emiI+/j1YvwpS90t2RH5Y/w1gp/D
IL5+pdgsHJBRd8hP8IP70KpS0wsneZfuLgqM0nMh0TJZXdcpFo3IRbZe95kqUaPFLEeQu+s4LP9O
ydx22wgO4P8+ASUxhp2+uS79ZwxCbfUDRXQy2QHelFXwkUJlqQYXPlcsG8oXjY+14zf9VUAX1tVl
SMGdwWkmxlf8xY/Kvp02XgbfhRu+AnetlJ4f05UDWcR+3Ay+lJuayaduH7NPl09ag/1x4bqSdqul
rN0EJAO8gK3zh76puv5ee/948mVZt62XINkGT3wsPFzHJMLCtmniCAdKmDCOLUBzxnUxDJ+Lkp5D
I+T9o32wDyLWXYw3ysUpT7vNrYUs48yv7UguIJ8lsUTEibBalrx7u8wpzgz6jvn8KgeLo8AzZUUy
DbFooFHLlQvh/AO9qwTu7+ugQYJPEmnYDOiI2HJjXLm8YmEOV9Z9KEUrbUZeV7u2RIFx2LY9feuz
wNDvesPBgm0ZOs0r+TcUsiPJxiewTZIheWRLXcRBG5eWjqgBzJ/omGMfWKgLT6Z8844fnrkJ19as
wJh9fqvT/NUULinbUeRmE2DGu3ieM0r6bQxMZycBIO3c/j7URP3ArGSzmKsJDwc0piLUdWlafNX9
iHJtXnJcLODVDjeM+qy+lnyWQO++ZHvDwWSxlhTo0U2LLIps5X40hDUL28CznFDYTsP+ncnAd0C6
yc7jjoRsbEmS5YUtu7hjJa8+ehIov/TRoab12L6KaCPMFoEHchlDs00UBjor3n9VDy0jd1QdXKb1
4UhHqgxGa2G/rGLkXFoAbhwe8ff5D3VtaPqE7Z/rEKf/xtCQFAuF/o8sBtxZjKBRZXrpxodgyb8O
b2+cHHGR+MaZHpnPBKra5mS7ALr7Ywc27s/OGi3gqITbNDnkcBKoZcHz11tvJOW5Fk0E9e+voBQS
4ihJftSy9wUQ4f+TIKnerC9uz/sA9wk/xpkh1UlSftLodYd9SGhj0QMUhBAOw8ExqgbJMHGcoSce
HZiE8ShwlJJCwcLWT0u5pyvzdgHEa6TAPVf2yYIrx96o5hu0wsZl1HoCXkDlB6sc/OgY/CoOjrSQ
+KeR+RkWccXiSZq7bsrru7xSBn/HFLDSKE2jICf1fejfQEw/jOip3TJqTrQ0xtGt3uMsDnGBOP/h
UF+u5Q+P8SR0cGPZDiEHd8yBcQg9143GgSKuq4bkzmDYXnqKUzQE3ZrsMIWKAWZJQNKpa4TB3mPt
mJFH6raFS24VC4MmwaCCVwkyNyOZ7iYIGk9t3Bw1rrobOvhJaF2Ug01nvGdCOFrNLBkOBQSpIhDt
xsmCR7f/ZSn1Gm9I7M/nr5avfi5FAfpYeMSybQM2ryAAAJHlcFB219dXUbRK6a8ipNRGcRGPMyfX
43daXck8VnNjVnDePbH35Ib5mVe92NZWHeIbnrnU+matOeEgxcuvcSknM0qyNuiXDkVP55qNd8dq
YbaUWz7mQv3+PhhdJkLi227n6ycvIoGvMVxT04jX0pphzumzVz6K/tClMGIbPZBdo2B4Edu1POzw
iOfr0H4kc7QT5nz83NpOGvdzx1Uj4t5IABdHeXdl6FNJs8CdsgJ4ZjPMJcH3GwhvN8BjJVBGwx5a
BKERu21DaojuiBofKVWHyQLYT3sfxEn6AZPlMzBjL2nSYuWJNqi8Wxel9jFNHUDN50bTWKN0l9wn
NzGfyhIptm1l68qAYViprEB6AUpHDIePmfbsXKbRDCoz5Sp+7KOzR2CXHyF9C46bZ7Eta6hrR/zH
asdqFUZ4Ce7+uL7gaQPRkUq9pjghy2cE7AfzevitVkWX9SWO9hTi06MMxuqJRqUJMfVSJgDHhvM0
My/1Ytu/hosNhUpy3cujbNyg24qLW/Ttfs1v9IYxvmiskCpRBjItxvDi11dTJBSXybzlSvwwsmc8
4op60a4o8BrVnsZcJv8HKtrQ1NN04whVMaZ790QrKklSJmHqI9x6bzuIE52xCUnSHotPa6+YrvNR
XGVDTISJ61GdN1PiUTAqD1ebO3QlUz87Tl5JhnapeMhAFVsJrzcna05RjIojsKJQCZ9P+/Me4suI
3/7E+h5bjneqJDsfgSue4bOc0X6Dd7/SLzYMZDJECq8LP+BABfE29sjzecL/yiPeuZOxl1sJZEok
8bmJhEx9kXlFe5fkxC7fchFxJYDa+jRgmu9QE5ta24ymog07J64i5tp4rUkppbeIabkrXJD1slUS
OghHRFOP+NZZK6nAR8kEikqczLYXzAXiE5P2nZCm2t2FXFniBVXZQ7PQ9AI7BQyWCPZb8W/GujsI
jIMW11xZrzXPsWdIpb5Nt7dtmxZmpHFruAjk9iQ2rpiwoj0R1weKFyD7tktVMsgroPeqOGqB+lvL
HhetWb8crdeg8BgT/f+xnAOm9fKnDTbcUG8qiqCQsqdB7ZarsQIwrOnQEI/uL8fBRxCb3hblH1Ys
oQgk7Ye1ZJxhTGcpHCkjAFkQX2rvdl9QYxjxie40TskcuuEEpAfs/5p8oIuHArjAHJ4rkRtnZAzu
V1EoWZpG58QYHn5C7kJ+smybldoq+wK22T+6jB+3jFohUpkQhN33wiOMsLUP6O/SOtepsr4pxDB7
gQO0sgrXokZ0Q6mM9M+/s6KNTFsBbM7i1V9jlTg274EL1WdTjERlhEq5ia81KxgbW3eZKsUvB+me
vMAv5/Sto4Kw9HUW48t21w84xWOtHhS2lF83hKKM+Z7C8sScSDzE5fkA0RG9M77RIsEKpBdvgjLH
W17Z6Kwu+h0Vl+TCxTxW34PKZRDghamyIgr1kYX4Yv/aktxXsd4FRpBUPoF2l9IdMoV0yMbxWhhh
xdq56j1NBQLaD9uYkUEo5WjMboR6rxCCxZIQe7jzFH9iaasgyENxECwtTx1/r1cvF1EApQFOj1He
ZUzU44mZmzWZWEo78R4cvZn19vBIoDrzxw8Ybn9dD33vnTvI7FVl+YxuaaKEGKzeFjS78r6C4rm2
Jqn0DMT+hA7i4l87Ooye6xmIkBeDL7ZtPRjN51lzZ8IUJOb50DjJdCgjiTErHCEXTPCxliwZlhuG
a3y8Vt2bB/jkPq4xGoNznFfh2NGhl5PggPLoq11WccY8YUxgUgDOEH6MFZ1VBHry02dyE/x8VfZJ
/LPWPGIPHCYF6aodmyFBjKl+RATQw4Zhzth3Q70PJ41F3jLohCh4FmwPdTOc/HpzGKhJwcF352NB
2Fh34Za6LhChTF5vhIYZcnkJJ13Uw4w8OdFvXhFmnjfY7XU+Os5d592PGQXlwuQgNy9VKg3sHFn6
CETyuKm9C7nbX4yIjbtMVrUjq73kf44ul4ssIwvcz+SnAOSG8xN3qQobmc+7yoBXyUFRKUuOgWp8
f2UnuSF8zZEzMt2Xmnv+qblFRxeVnEuXPPAvUMRqHktFYzzlE6GSOb1hSDZ+KHJG+mMKF3j/aQ3x
KSb2XmDYFhW7EQBIm37lNWN0iSWkl07QsMthI2I6wHQcuBOwIoeF7NGriTtqchVqgoAJ/Ey9PTNB
S6QPDsi/VWjo7ZulmQzzhtqAQqAA7M4tUHqeOy/1aXFOFJWx7Deau5u02UK60o88RG9HAv0w1dbC
Qi5ck0ljk6ifQFzmjgLfwwhrZcrQCf9lnW90vaTBGVEAeN/Wz616Ldzrc+8v8Xi4630gKbf20JE6
uLme5Q70BvVar0QeaPMqSRmfNgksxzW1uQ/XisqAuEWhDVq6ABStGnh41L+YE7Ls/YHI2SHLqYO3
WTwQGg6MEEmwNf1HmBlbzy+RYT+3iQLnpjB6W+4XneBlnwaY8kv9pUHlQkMsJvNYcuTaOCMm+ykP
ReXOtayV0RmN7AzgDAhsVPNVZC7oPS2MuwQbcvmprJkgqmRfVmRfdsv1RgHQFfAhvwwH8xMtbgPe
rzPG/dSy9grBEX52wmxb9pWL7XuYE5pBab2dLEtjaoNIU4n/V09XxO9ZltYlhrDaJYikZx8KIyHJ
XF+iXAFAdj6HsuVcqGe9d8VQW5vDTO2zny3iiyI2EXS0nizaIHgYNtd0xScH/jYCfglr2XCtguNK
a8MYI0Pw0n4vtKhY4FnwctCTV9figv3AlRTH19jl/NJt7kYOgj7ajSQ03XyCyE5E9rPvB5cBi8qu
hcsZFZp3wETh8VVMigv84VY4GvdEc/YLMMy3KzJ6HwIPfAWSZz8OtZa+H+KeeluoLKAiGn0jNTXY
Y/eBNtVIFR4rlZEHvolDX8afRhu3ZsH5LZEu5fvleqhhrUPgR6HrR5mWUW/7oXIRVmHho8Y99q4D
cqnoT2Ztm+J27sh6eaILc/x7DKr9aS5rT3YsvE2NBbLeZagdxCvWzI0oL1LSEgyXMDrqwW36hMLB
gwJytw+SEzFcGDY7Mf+LAKc0dMZW8cYzLxc4JqER0igYDhE8Xes+SDTAAoUT15BHIB5IJhhqoSly
+BSDkavIMQlS09IqEQ1+osbzKJnaQNQMvXIl2Ny+LyAJxpjymJdo1bwBYf7Bsbtlib2pa1jkBgER
yRkwDtuu/5Q5DR7mVJ2Owwr4n+GmXNlb4KrHQZMa57dsrF0YnDyEkl5OjOR9GD/xijGEiXRj23TI
D/9jcjrl5hEOEv1Dre8KIRZBHFLky2jz+Pgwk9X6Bvp0PRtDeItrvr04bw5cNmfwBTG11yXKL/gJ
qrp6eRNjK09U5CBf8nbEpTF3astj0QEcf9QDxRKvX75vU5s/5lpGz5u7mcYHfSipKJ6CvOk+CmmS
R37o2ubizh86fIIj6tnKfbkUHclxF7GgHmVWEIZAj3tbpAbl79tGCUP1ZBCt47Q+31mgYnKJukLc
UBH6p5DlVQ1BreJIjK7PQPXioQCsDBoNG1z6t4E52iielt0plWSMB9+v0ODyBtxQEDRxNch5KFZZ
+z1NF64VvJVKhYJdLkuUO15gKzi5jlt997OG7uG3+TvYn8vjc2URRm1IcViuHVTY+AlpWUmBV/HS
Q8akOoupfVu5rNJDCm9ZZll8jQPUWrlN4zVUFV2M7vraqd3xaNUwnM/0DNfNWxAK/qg04K/7uBE0
aMqtnqv9YknheHNHtWSBsLbzcj14ZkMxziHwB8Qb1PzMg4WOTCTBycVHDgnB/TDBGqHDpYAkqEFq
Yocjxv9lCY5DdG6KRcROTU8kPS6C1e6R9Tpfqw4P/f9mPvzFroRGJVlcF7g3G4gcGxpeyuYygazI
K/hoXroLRR8Bv8OT036sVta1TvjWsxSV1utaO1Ki4ijSfmvbAkO63Wb6x3U66oXGNHGqYoO9MWNP
OxvUZTQp6sg22mGReRC63c7iUXIJ2ZeDoJ33mRhRpD9oTThfATtraRlzqJYXL+nHipmeV+c+Jw7D
Q8O3Qa1FWAjneSY2zr7pjcxfSVS9LxTfUFTB4ZsbJEedQG8xoLj03GIkXi3C8OiApeT591dEsTxb
GIg070kLb597iPPvb1LinbnXxXtSEAHVjFCjO0e0hk9QKfdko80PeMRlnLO7+OtOBUaXZC+xNYzU
9OX8fdJN33ZmZQImLOWtrzXEhQ0vrTkEfbZOYtvJswxHEWkgOnc5bi/pSO62XaJO/S18gllEptfq
Ow1FjP9zlfHTb/mYsFFs8iceu61TKvmK6PFcKgwl7ReXtlUBQNTmDeL1B5fM/wf0kwdRg/Af73Vh
paxApwuGnIC73Jxz2b3B/OsTVvwn6L+Zk4jMy767F0T4ZP+whA6lpC/hl7t7W1iSeudFNBU4D6h7
UptlZ/ckcyYewsKemEkYYnKvcSc0cymKJnbh3F2qIGD7GvygB/pee1U30HryvS4Rn1wbchSo6S4r
ABcfPXQz52QxYTNbFJSqNWs1jPO4ayHt3k8cX9uyED/+qynN4+18/ZwYeGWh1pABzZx8pf/J1HX9
I0Jq7VOXiQGjLjMtwGBg2yE2A6loNssutH/89wzwdIPEjQZcbQsVwZyG64JffUR5FOPP32fy/bj0
5SLDScVkuvdsoyKR6jO8ylgl/IHp8YG4I/tXxyZztnzxf4CKBiJz6dkyAT95zZu+DKNVYZAd84lD
iwPHzuVb39LEA45Nt9pf+rbDNhHWpdVrZ5lTI4qDlfdCLmGfIgTpEdiPrziNiCRok8/a0Q/RxSKe
FnfU3Gliou6Azx5sAIuKgdBxRE7NQAMXfCKFaPEBkViGozoPeunnHAabDGUJ9+PsLeyjpJ3d0pk6
EZEYS1eaG6p2oglsBdxPFzp4btPIm+AlyPhiY3LNEQf8I9ErBA2+ON27YKFJkUoWWBNdc0DmHQ5Z
qf4kaSps+sCYPqmiilwqHIknkiBKWzVSM8uDAHI7bo6bW1kkp5Lxd+BzfkK0xJH8Tsk6pV9c1Fq9
dkYx1JCPAuJ8Gn4f+rMPaZogHoU8Un8Ld5Rmj21qcpAtIBZjfv4h/dbYpOJw4R/qDj891iUpZLLZ
444XnWkxNY52iWVdBBIIVe5lt1IJnAbnJHEifNNao9XfOq8z6X+0o5bDhEnK4DTqB62w6Z2SXZTV
EmlyVxP3RC4+rEwuin49u1YZVSX7dhUWX0LNGm2tfyczWSGFRD3fMuqro3wMHJi6AnlWjIa+sHSa
F6Pf7pFSMtADHYi7tprhOAzxtZAfAh2nyoKdwzplipHl8mscVKBzjCf0bXLlWsdSXcjOwhoRr5Dm
FmfOLDpVIDfaA5IEvt9BpOUv5eDLnmpZj+afOwzMfy2PqxUiIf3NUIg7S5/nKcIxmedbK0zfWIRN
4yO8ckLlIzej9hJuxC2BgmG6JIQXT/7+Pg5r5FoW5Jzm3JzRwMtd4Shj7KiEL1V42h2YArtqO1vF
7alRXsJtKl2Rs08JyB3xbweLwsOqVR2jmuNwVLuoSmPx65pWpwj/5+xg4BHX/Rclcqps+Y280qYU
GamAcb5wgPk5jquQJ/ln94vBNdGXp9gQ5ugSNNMPdqExNWASGC/8NDPubJGGsYQWoPaRu6jOl8gu
8q2uenipXX2RcrhRLIgjAVkKz+CYGR1RZO1GA2XBjbcmQD3W80PKhhOYbUlPqgGTEWYeMBVyJ0be
HkGsc2CKAQ7wjpc4C5WrqwmvcTkpvITF19/0PX1FwE5c2ceTD/9QpkQ4/POVCCRNZy/MA7AP+Ber
BRKHDuHtG3WzsBHGUgLsUxfpr/j/1YWnmxJngvHniXKmbO7GjKJUpgAfFe4LoCy3/1EGd0CDe8PY
oo9SCgknMLuVV6BSzaro/2jRET11/VK8otw3p3rjvn8b9sBojsmMD0UvvM0B2OuQEtAxOUongHhv
tT2X18+b/uFnY56V9/sUNj4yoiwZITcoOQDt9BdraR76zXVwXgn452zR61Nsph+MlNYKJ3W0QXNS
/ehkcqlWToD596+SxPvNE9XVeLk/4PhJvHBh2payCluNxAKlRpx/c4eh1dyAkX4uvdpBwlpqkU6r
DzjY/MTwiEQeD8j7j4oEDgsEEK6LaLWIp9+HBq02KIyL3CM5fxkBXUAVTnijck9dA5uTgc9v2lNm
sZ/1kUV+vaCcoeEmEmjLrNwc+s4t/wECUkr+48CUi41wB2v8E5t3zTgeB0mbcJAszLN9C+fUgj0L
yCR3PsxzUD1OHZnWyphfKLCit9M6Mrw6xLjS2u1cJEpLH/yKJqX93YCpfX/zRdZzJdB11MA4vMGu
TC2CprqGg3Kj4l03YVFiNdWSEOX9FpFvwqpr5sGsQm3UFG1f4473VslqW0zZAF8FN1mex5vRL9AB
KGysRFHhHmz0DgpfHQmv0ZFxFqKS9CUZYA/bU4u94Fm3LqcsT+NT8EDQJuKcdyqeh9MCycCZJCiJ
Da8qlzpZuo+Stiue7Oi+TnU5102Nt0bQqA/gEH9QUboJNi9B/XbkknXEOqesDiLBxqmzysrCrU94
Wj/TMBo9klClbFk5fJgwzIm9XJ+7pZ/BPL+bwh7HcEm4o6N2WwzDn/cEuQeIES6diteaOwWheeCJ
INoJ0cts60DXaaZAl8pM0aGFLXifnrCcUxnQQ16dxgqXIVGMBQ+UJCECeFpvf7+Vv8G9q7YhSaAS
wFFPcE/ys7CJScguRt7Utw7e6/vdDbEcxhqTrWgWxvmpoVx1aZlsO/16sd30j1A7jCEv918ozmDT
FOEHFmkp+gTBm6t+AB2kD4O1NCp28Xqcgd5+FtXDRHC/VW0UaNtTRkMbF6WiBbtl5ASDrOlyucWr
RkeFMxAE/WfmMxLlIWRXuP14kXERfBXLScB//7YOswGal5++P/aLne8SycQp1qEhivhHdW287eVM
j23hZ13hyZq3R7tptGEIlhp95e07NLGe9PWvcmcrpGvGIbOGRkgnvIwEwlcbiQfKJzrGywNq9fiz
Kdjht8vIXHtbHEIhGDn7PcsmGITU9S14gb51G3LcoFnSHYF0kZenm9k5ShlkUgb6WOJG9f79s1ts
Jkt1GxKQqDteg8ahzSW0AixLRonppZuwKcJjf8MS5OkD4URiKSSM3AKVhAL+EHldjPiQMQZLIRT2
2F6CTSIiuir8FTLsiC9TlthHV50uuHjNvfeOiLsd1XGoGtVMDh2d4IfEqWWxHtuFhRE9KE6pIslY
quPqUjatisz3V3/P8fbx6TjdADAWYUJKGEKusmEzjAdHhvzL/GJgmBGAfvlEj3/BzJclXOwt+f/f
+xZFe29enh9FB0/tPRNvBvTHfNRDEnUp3ZoPF0uJod6h0A2B/yJJ6+UzfNIMVHG+4Crp/kncatij
JILNxTc0OBGrsjhW3sRlm2nDXEVa/q+KY7uUP+WudgCJVfdou3GIPO6MEvuwRDCoSIHOWhT6z27v
kcjopzuJXLbf0CeIbPL5LQ0OOLcSz4T8lrcWrLhz9yxzYvrgiI28CywWwCtnmZ+KGy306/BWbC5J
UfCHOv9JdrIuYFRTXkB23KDo+wkZUEcFTMNmmPtMnelC7o+WldK/fF6saluxy8bWs3NlT6Fj+IlC
DUo/wCPwghfTscbhtVaLfhixPTMYU2c/aV7H1pOa7n974jh8VskkZPwGkAecb3NwVvc9yBdv+SU9
A/cpB7Ve5ReaqMvDOlDzdzZxMh1ZsP0kVW7rXLN3L/V+67y0Wkmrme9e1mdXYDMozirmwXErXPNq
7pJ2sTWXZFYgpqjsjd78/+xJoMMIoXTxq1gehosdMLtFFnQsjrUQxQ8Oax4ftknVbABYC3musUmg
FE4e/SviZ6Kcqgmy1Qr54P3N31lolqcogyZ0jJeLyROe5ZTPkhS9xANKT+O5CV2iFOHvz2NvMQT2
Nh75xIYsDpqID+aZnaoxfhYcPTVuatpy55g95K08cxgwRprHkU4qUTTdcduaaPZV6br3Wj+P5FwC
tJdZipEHl2ah108rz91fw+FJMhobPM3JEmImo0p3a9rgnIg2g4koF6ZA3H3Tbywy727FK7MMuCnx
gpF6E1ukN/ezeEj3g7deShmEyMOgxPanVlqa++0I9q6ek75vw1Re4A65FF2jeKv7fYrDx1ka4xlP
hpD5B1czAgaC1VPwMMlfdZk9Fkd1p3Ep2WHQbMscff5+RQDfN5ckQN0UydyQGSvsekz+J3yEtczd
QRcHjg5aqtmYmdPbUvbiOlI5qk8umbn7RpWCok+E0i9frR27cUmEBpGt+JUB9rDTILf7cDO4fm15
ixNserZ27xmbZN4kimkmVOltxBYIqYvktI8x7UJ6aKeAUcVyYGZi+It5o8Xw+cNEEHFjmhFc/VO/
FEFNkXR8Ynit3iIKFOc+Pm+sJqmqIUgJa4b668bLqNY0p/GFXS7n9KzsaubBF/3x0gee7aFFiEkI
N1/6SvwKebU/vt0dhid6LJgiRrHtsEaAlFa2WRj7D8dyiGLLofczaNkXoLwugyOeFdjMQYD8iyw4
JOmwbGNjfb/cuxdp4IbHZtdkyKiEFiS4aUWUg9JjNxmYbK/66l7cFxNAI6wmJUQRvKRst9W+L8ls
ZozH6PNXuF8Zh1TdoAvsBWlXKX01QzS2O3rrrG8V2MGFgm+fQCpmUSWuk4SF9KRKTzLuGSfqnX3Q
WXPN7Kw69qx5qttEeH2xXDH1hf7w0lXXQbeSLiNR8ybLnlKOJOaUgvc6dWznBuCtJw4F2p43JErg
IvCF7VzI2r0ZC/2F691F/Fh2hXX2wgw+4Gu3AK5lMfEIKRKzJakO3BV1xGWOPRhTv8tqVt7RSG3u
ByIdybo/7BLAkQZA2BKmxvW8HwVMAk2rOqxS4t9Hq1Uc+iRWoAPoeLYXRClyuGSOfZBkaaD0KmLO
263HWe7Zk+/aR/3ezYXTHLxT1WM5ORHnkiCVK42OhU4gou+uba5bl83IFGRJS6+HzZY7D09D2N6a
YfqhWsu9qjzAXGHXq+CRSHky0MGpfANPB1QIoC9ZJ4aDvZ9lDt/SHWa9+BAoDCf9vcHOjkqH32EL
7b+RVHENcofSw3Y4EbRqz3rjyEYFSJvuQCBI43Hry3hvwbjJMq34BYEs4nt9WTDspWpgwxqAR8ly
qP4MZgVpsvIYjNIo7rUsogHjb94m8DAqQQdd7vFZRiLSfXG4ycRT4Y9wxednkm5qZCU/NyCJWNaQ
vjIZeT469X96rVFjptaPxWGNX3dc9LrFx5ccc/SJoBjxefjrn8Vj3FcJ+3EsFpjV5rPINMJBem+q
Uy8Qhjl5ZrLv98uMpN/Sl1Hw9Fqj/42f5KviOAbimLKCH94f2eSpIHU4ePZuue+TWE+oCrNs114W
TEmkvB3hw5JRy1j0VPsalWtfEiohc6fc2NxcjtpxxziEwp1dZPnmmbqtgYA40+yyokZrSgkiSXg+
ZAFKl88Qr80oNRMzlgM296oh3gm8UqqJXop3S1zKjvaZrqMcr5DNUqTaKATYwYQ+8za6aT87BsHb
iw6JGei6Rv1rzIOK6dni7nHNyuW8PAkgRR1m0zKokcjhGjANg8U00qEEmBj/3ay5Z4aNzWrnsh2X
/0u6dANOJZy6ui6cCS/69JGG/Qo1aVuF/+Fzs3eCOVRxpcel85F6XpIz6VZtmxGN5MwnRTDjtb7H
qwe+bSSLlV7/146i0jiIkfK+8M+Nbj7sqVGaeLuMiPKKk4uEKSkNYeV+TZBwscupY+30/ao49kTy
/LKz2Y33rktR+9ZDQTEidZxOxs+GR7TmFgMwafL5I0oYgf6lphWsqQSp5KJgyR5KQxnP+Xg/iK4R
UWNMT2fuE/YN7gotoOImGD85O8xw115lTJxlFA/5aNPHSU8m/9W0uFV5yXOZTg4KOxRdbMbkwoDn
WXFIIQnLrt+zG9Ps40MQ50Sh+idHYtceJrbq8pljcf2aVqeOB1qMfIVqgAdDfCvl9c8HU0CvAkEk
OADQiyuGdSdQooQqraBEyzOSQMC+MiyJzb9PowFJsne7iQkuxMhVdxFiGdyqAYgz4a1OqDQU6rTv
66KQW165le1+NJkRFebm7Ij0LDKq868DUm2SDlYqAmH28e6soLHscg8DO9eQ7DEfZHqDpeP74FCV
lbuT22gYoHfO63x37Mg07wqpiCliBb1xeuijOEkhEjM1exu+oxXb9DPFoOYCmtEqPWiXVcpa+Yk2
UanIcT7tuy6p9p882SOtCrDG1+quBGJcHYTgpEPdmUdkdMR2ZA7mgp8w5BsGQKeSb1aKJOlUOSR6
j4asaHYxrUHRF59R5U9q99Tt51zy1tNgRa5l6yCxkrVfyN+yoaNBs4L2kvdcKnPZV5iG6nxyEPFQ
eGtoBXzUJ2269c3v1LFdTainWc2lw31Ta4eLHUbDuJDkvbnm5xiRa95nvvsea5aongU+NJh51McW
xqb5/Pp3fS+N4qL4hvIDwUTh8njVj669YYnJUaINvWxteDmEgiMtgmPxjZ0zmkYKq3AAOJj3ukdX
MjKm9RP5xtzsbdSJ5sP2LYTZXOiekl0polVjhhouJHM9RKh8vj6dthaDXC1yApHNLlUroNL8NGWc
1Fpu2Ay4HYRyxmMXDOuIPcwkz/fPX4hCYntk1JBcWQCoTSTbcYQutmFhx2OSOqUKUlKpwC5HyFHf
I4LqASiLockCiNiVBu8fnFw0spTjejq/QzWYMFqrzuVJxZ0PD2JdnuU84u4OLcLSdMaA791XT4bd
Jr4oijxbVWVCnrHUyM+S9WA//NUiJxTdTikkpxauKneaLCV+roCQLWG5eSb0niiRF2cNxYEqL1Lg
zGv+lVIshvD9vCPYy8aG+w2kQJaX03DP5E0uvm9I7B55Tp68s6SvHhzqkb8o5cE32XqVmfpQ4Jlc
qBYRa4nPQtN6KpALoiPpiktMdCTFceh9RSYsviJfqS3hESCoqY6JvREd29ufeoE9x0PqwH+R9wKl
LARCHNpBKiTWC3vEKW+ZKZONZ0g72ljXikKajDEfFZTL6BnT6d7YXrtVHNi5vA1nCnYV7/xFt6iv
OnvekOL8fihHXuzABSfmwaj7gQnEX4s0kXN7zjak97xu8JKtKk/Js3+bDTP+DCO989RvDQOmc/Fd
46Zu2yZ3Z5xgjUFGPxKz/cwPE5r/dkt0tz3FGWXQ2niu08tmxI9E2xVOOX74hbh9jwR60boPjgU6
E6G02NcCA+e/zt3At0m6DkJEvEQ67v4xvAzPEDHLyKq+X57PTid+cbqHwlh9Z/m/HQTTNGZOIbaF
lgKy7RDh95PJGdcT/X4fKvgn0kjHOx0pdkfuIqEDjh7pEUSu1aU14QEPzR8CyundBgaqUXl0zrHh
FDGh/ZyMXL5Y4CKsA/0TvoPL7vrSRkApv2GS8dh3jb3uAME4fGPFW9Q/yaNKXPaCAk9lgZcWs+AO
fSsTHGU0pe9haSJOC9plorNs+FyNZKDvHAbwRUw7rfivMaZsOnWzTzNZ0O7BLJfjGkLHXDfEYVzy
Meq1rLeGvGb9FD52GLJIlHFm1KigYGveQUuHpcbf/+WiAGfdQPnpqbdQS8MoYQL2MNlkshL/h6ls
q/qWenXrcb/ITzuFm83VaOVPy7rumbkz5b59p4I2slgP/HpE2y3LQnZ6Lzo0ljXjTWvqrn2n4pAt
XsxWZ4YdF81Xfndpw7sO7qDrNWYg+OCqkUVUwS6t07Qj52vSnuz4xSL8wn1UxxsbtIwIopfMoH6b
fqfEBPDdTacCEfdyZEcXgfvvLE3ZSHMGrBpNdfaLdhliWT8SLZ8PA4+oL7FEV5qYqYDhvkGGGX1u
xvwv5/GnjEcOFqv9IBP1fpGgVR7anBGutTGzQJVsHB80EV4FPXYyRsuBhNMGqfBV7+mtiNHeK2Yg
dR0xSBew6rDwM/4Bc4z5JhvD3qzKng3LALdUbesx+/c8JWuK8XE4SvSwh+k1AlYNRBf+5hfM7LIU
IqEAGBJIX4WdWI2lM2+1nX8gVlA+r4PKySjXTZlsT/J0x2mKGhrk3BPmU7L06jQAd+dDixMnDC5b
3EtmDkgqR86RicYhDw+qVG/IVmFo5aMmDYA0DpGUMe3LGVPEPb33eeEcjJCWRzxVLpk0KfzpWtFt
qcRnq33s1es/ezJwPtHk8HGYpAWlplS3lG+F3dO/pvtGhYIzk51BA47YDHHfO6iJnLd6GYaeMZKF
mIuXZ019Jr9APvwdNZfauEBYqpfl9ubPncsAZXjtA2QOpqHnLH8gEfGovGG8qqXLtY+4x7aBzSw0
uaBE2+G+7LN2at85lab/4uFmhFezSdOSdR1FE9Cz7pmmeoMZmOGt2KmI8v1wGj39yzi9UZHB0hxG
yiKYVECjmsGSiHiLVzk7d7pavFyEdzb7GamJTdwQPcq1IuoMd6EYaVaPyZB88L6BssYyi4by0qas
wzjuKeg1Qpg7gldDbKLJyUYQyzRHK9t9DarwwJBPdk+F9YM0d3CAq3Jr2LpcxTslU8NT7KAv+zqM
l1GxXDlLDVyneAfTV1Yezm012wxiC7mPWk2JbVX+bJg0B7491lZlfbODCrkZaS1Siy4Wi1bTZo9F
cQ9arboV5NKJAF2vAdtsr5arMjriNGLJTgY3iKebHafgHN+hhxKs9kTiSN5Yc4TQ+jz54cU7FBFq
h+gat5v67XygiO/BakT4ZqIDIi9U7WiBoUzSJ+9+RLvneFuEu2R2V4TZ89+dManE0az/8fmh4MCC
qSs4iGOy3d6B1OpU3Y6+mEDarDvf6+4tKYEiJXjFDR9tCxg6Li0NyYjG8yCopkNVSV1J39QFcu9y
2LTc1ippF7JNiCD6GnWpSr+y9LDAkC5HQdZJIGJhNigSblaEVZXM28X8LkWURqpZRfgCIQ3apuAn
8g2YKlkNZG1zdqCqSQxrjChw7IBqdmJcofvx+cmFQ97XG/pFh7WxegpElXEbk1W0qzf2wCP76B+m
8C3MSDEpx35GhzcEckV0Xn5sngxt53M5kQ3OFeA03Q1DE3STsb22XmGo8CQRkqW+8X59Pw8xXzat
fJKD5sHOm0+TnDlRHhW+ntlMl9Y38N7MbSaBUkbzxdaW8sTlTH3Kn7kCa6RyLZzEw7LWkOyadKYo
8h59QuqLtTGp+Yfnr9RIfLYpOSmYy8jk1TCDz9ROGyyUZQabi1eeO+6qSpAzKKuw3ugBz4NfadjG
y++OLxgwi10FypXaS+ScsOTEmch22KOTrybe8TeqmQPfkcmlWEFTTWR5EfQVrTJH9hVQP+vyROgp
ZX/+yIHnlV00R9IFLahxCZxXR8tgTYw/eQMck44leMFb6K56K5Ogqa2e8xAvQVLaz8Rhd9HW1ESL
+5kt8gm7NCkDkYGARLe1Yqmo9yk2S1Iw3hMCWI9pJToJi4FUTy3f6pA57penocA9HAhfZJNPmi1A
rWckJg4ei+AbLT+2NQg/CWrxYB8eR+c/uqZWHpjDwFrlxMHpqTS7gW79gWly72FOMz1CxOrFuFAw
9zUOqWJxfJE9CeiHDG531xlIAZ2JkYtutwruAw3oTLtZN02MBSg1Xzx+vtalncCFitLG94DHgSSn
PEgplrDkL/kkNy6JP/yFd85Weq7k3NJo9q9nbfVNii+e2c+d3h4MfXxHJs5XIpwcvJ+EOun9/gUj
Ew+S3nj91M2sQWwdKr7l4/3dVxkkETsPDMIaMzCwq1SIXkfVxrDLm6GftVfsargyo4R3wmjpxdg3
BXDkdYRBx/pkQ2kXlJg2yLXfomZ+b7R3zwLS6phG1ENK1zIwM5oZYM0TDde8cYsEmFTpPXmN0hZI
YuRBmRrsZgkRH2cN++bMNOp0LDqVMFswBj9+3WxI8y67ncgioppADjXFn5yj2AlZOkG1tBpYtd5u
pfgnydszcSoNQBKKNGgM94oEpFuh02fgz6+UUMaiGletOMefwCvSyNjjMwOSTDCQjDONYqPb8Bz2
srl0Wp1rU971+rqESOKjnShwrSiGayl5pcOWZSMjRta1cWxd75Pd6LFGyOy4K8UdBmx3C9G8zR12
4nofw9cWvil7RHJ/X30u+F3OYtBsF2R/Q3WUx8cZ1GAbM4pwhy9rfxMB8elX2CRFHl2FQRlPC4fh
zwvSt5C1TNtUVjC6q6l2xh9mkVeCF8j2dJNwqf0xhTx7yAPia2UNhZvomgAMfl89fUv1DpUfP5uq
WfOfkL8/linsyjBeVRIi0isSxedVV+hCa4xZuktMZLJAKdDm8dmBFyRbMmNp8MyDchBsghUYALY5
Ew7c8GbuHp73Roooq5JFlMCtawuLH0EgwJf0bpR4BTRH9T5EoR6SfALrmmAdwXwJIQm3JpRbBJMc
dB0M+l+oc5xPmP7m3rr7qMQQZSSdn7buQWrFnb4hbMuDathppI7TXveJijA9E8xF9WXRNPIXYkiU
yMtB+h2SzKwyWxPXuGopOBNFRBEYinQnwWz+Ptn20oUMzB8HJNFlvSUvdbQ80cVBgobQ+iCgbmzS
pXme21Fd05a9op061FUh9B3ZsvG7GDLndfOqaAm2lwBYATPJwQRVp5nAqgjZ2bLx5HKryylHpufH
DC0M7PHFindS7XG55810tWaV2RN8Yq/swcKtdQfJ9sgXHtK1XEUHjcEj9Cjz4+BI3P/TsEvGxVFh
n1KM+7Z9ghRp42pWfTvHhA3dfUC8t9C6Qm8v44I4wQcEQ6hyY6GdYsp7P03SUGC3dBDz7/VXfKyw
U+TBweSZf7ebJ8N0k2jSO2lnDeU8ex6vhWpFlrWDgHy3pC+Py/4avpczLR/6lVQX7F1d8/VlFCo9
PgrXgy8ZH/4WlWpkotMBdtKwuopB9DzKfe2SbbIH+xCAf09E84PmB6E/VhrfrpDJP+PMLOAsrfkO
ID0joTQEMaHLzho1GqwX+t51uOJOPq2jLOmQR4v8DUp7mBvbu0Vt+xXCyFlE4IcL2LC9NtyC8JkK
DgVGypnIe6oMA2zLyMB8eE6X3Lz+GUs14x1G9r30004vQjDG7I6nerB72T/9xsjZ7AzKWHfTt3qG
1AeNvSPueaW63jNXZCN3PAtQ+fEYYX4bFisT+8J/ogG4JeeG/yO3Zd+2W6U054RYCU/kVTh7ukTB
79TAMCteritEriE2dtGrNQuhHkKsW+Hkk+yr/IUH8DTtaXC5Q1Mb5J1WkS7jkV4roZxqJ+NkZiCR
RQv/2zRq24saOfa57TouFYm7a8+CfPxEZZjNcchDqv5AGZqg1+THltIqxy/3WVBRKOxHzqO6RtMq
RAzs1/M74tR5rpQfl6nNXmw74JhN14kn6Qt68JD1CFffQFPyTI9OERQO40xWNrfiUpu2smVlNJQz
1o16Z2BoBlUkuqGBRoKYOh0JZ1VzGrvAbdV8S4ZNYaRjdRXA38So4w398DJoGTYS6ufaizCZ9joh
GCGgfFOiS7eY9gwK/9+CRVft1C/rX5cR3znU0VDSP8njPchYbl1LrYIpkTWb9pr1WUdQLC8pB95e
2bLxgXAZj5JIsvGRI9bC/ey6LU6bVTrxtwfY0XGR+B+XcNLe/6J91XdGkGuswLcMQcuu88rXUDf2
ReE7iv5HGMRrlC24UUqRWaXFXlh+11DSGKJibrTYYD/vMIrnAXI9vgPWVkvWaey3uWEM6j0xwv9J
xKWLVFzuk7G8FpH9UFLabYfpK3czeGThDK0vsfg2hHv5QqrRVumxWhUbAjtRTH44KTgIzbtBdlhn
4JYbHDKzL7kzWitysnXTQSxe+o9zw0In9qdj/SfHYunra8g5n3faeBIWu9d9pfnNmJ1g9uzNS01P
yJWVKDKdCk6OgIuMMneTw8tExquCuZMpaT1onnTiNfzPq5rH+4S/RIVmXBE/Qy1cjf7o1Ll7HCt+
m7g0m8YGhdPkPTEWRfKV6gAaQQ3wRSagosiBwVMaXXFQDmHzmFdQXSfQb4AxarOBhsAPMu7J6FaU
Wp1NXb/ehO1I42nR6URdq1mbfNk7BBfLl2FoqzGvs6vKsS+v1GMrxWh3aNO65n2K9ECaCZrmP88C
98zNf0d8sKRcsOznZHVBlXbTtnuLWAN3yJdO8/i1QNVI/PsQ7Io/9VigsjiYHnJ4AcElDBNc75jd
D1REaoD/goQO0kXWnfT7DjB6LBRfSa0WBR7vboTirwKpLLuEyEz1nIeqd1DXuFhhMblRbVx+m94o
3dHa4t1VvPKv/fWVlYzj3GlV7ZpNJO/CwbL/zlBtHZvl2gBvDUePsje4u0OPMaj62IcgNLR4FtKW
mTm91u1e4EeFPL6tfpSnkcwNyiIrsnTCeRiHFxgw10fO/53uOS3tfZxiafWL79IvWYJszNpcY2Qz
bsoxX9FA67JwgDjtogCTzGs3I8kIrSlESaUvCbtwLD8P08rfiHeS9XUZzeRSILVRZOSTt+cPap+T
db/MdNAwSX9eswntSMxlUXqtiDvH3NK3SXxJX3kB8EliNPRvj52QAiAl+W4HgypkSsS57Vrt4ako
szIg49vNtnQn9MPLPWpGIM4G1zc+JAnHqlo2cmT1Dl9iGo73BT4Ddh0nHccr9k2p8JmCXRQ0dD5D
nwV8uQdE8fIXujBxyZ3w6f0RWSu0BZxK4yI3ZCVbqDNvYVOrw0IPbVn5idPOdnd6GfG8PCvGr9/5
ZeaIVnewnMdBw44swTcFOvoxcGX76CmXkk1QEcspRchMWRrhu5s9KDbzHl9pgIuj6xacn0KilgjY
fgIoCuldYGQ050V8ndKja/GLd7NcNvWA353KcATKJQrd4sm41WDfPreSI0CTRBvBXUumgbJObLAB
7jAtjNoMwTHwyC5aeOCdv+hW9Ei4IaSo+BCqSpteY3PMnTEFL8R27i8nKqmQsFnlgWzhPyZjbMYZ
fPT8fK/9UlqG17wiRbm5sE1FCoErHx2e8Z5VvEDM5CadHQF27ydsRuwUo3OidZEa0dU8pJoQm6Rz
iBkVPXWvPlksWbaBbwpT6nM2iaUEHfDOLktLpRNZuP6xosMK2K+BqaWElg+cLSstAqYKQISIYhgT
Qj4jk2HRwC5fCspbt5+GrO5Rhh4iq3odrXf+I6gRfeaGB2FB8u2yrHxC+pFpVfispRfERBP/E5l8
Pi7LVZo6vVKotdYEfKolZbAgYe3QeRAM0xdsa6AUkXI81prrns+RIOaPYRlt5DcksxJl2TbtInB8
UN30ucX+ZoBiWo6jXi7LemSceZc6OBEe+WL9NHdQ54ImSRufYflUSfwceAAsMXEl9E5wkW9MDt8j
+ZHrBT9LiwxcpZqE5z3e5WPSCmkXX6E5Vrj/2yCtJgoB5OfoJsnSCTQKDzUryYEp8odY3gC+Srdo
dT67w6kRihzHCf90/7MTWfS2iAczHHfrpuWHx2ET0YVopO2hCmEkCEXV9xYE7iHl+7iTu0PteYyY
VL15JvK5/0TXfn10OjEi6MOoPm27ExWKaWeZPw3HsTTnCfAMia1JbXzUGHRiGrY9HznW0N359lLY
bCkhJOVZ7G6qJqHlezFJYaMZ3OE6WXOzSyqxam6jh6yTLxGrZf+kGmrIWmMMi79Knq9h+wb41t9p
2lgjYrR8KTDs5IMz8HsebygbQXG48ba+bRAJkWRQWQGH8w0ZYCmaIFzzw3nZSk0oJV8NwkSMLgir
pn0cPS9S5I6Kwl9csG5L+kvxAkCHC2w+k30QmjSbsyBOyqn/dCxgoC/K4nuxWvRCF1uNcdG3uRsl
Qd5cyAYV3d8kBVuNpC+mrGcenegXfByyFSHlK84djTCZoazs3s/kpI0ngxBZsXRjKeYaH1jULuIv
TI4FWJhQXvgaJ9lBIdeT4b4zfLVfkstWCU2GqbgtCDX5fEFJws9MU7cNDY6Cx3SupREM05DJNbvG
wRjhl8Yltwif4uvm9AczPFjLVuVJ5YqiwVcL1a5rgI250lCD/xtDfm3keGb0uLmF6nnhWsuMOFTl
EfgoHgFZUjXihiDLJJ1LhR2ZqjKuP2mWjUWD/GH8I9BDH6Et2c483gb6RVcKegrqSfNMLZtwxY6T
8rkd2hA/WASS4Gb2bE4xX0vfcTOMNwv04KhVW9NmoBMJJ/BD2ayCZMW8hIMNfeCFrwfxrM3dRLd5
A8Ti4yWY1iHasH0D3cJOX/76H3j9aQ64/h876/JUtId6QDMKh6YtePL3HiCbvsX5S/rCTZT/4MQw
jOklCG0x2kCJO/Zi7iYXaneM2uKgRVarezxcwhOtkCU0FEt1K5lo6/LuSx03ZEBJ9NnxIy1HzJmK
Tu3iGFTXK+MjLvTSSNowpU/PmuJYpVJ/RZw3wIesCfP77VaMrCyyB5aGymWesCOB27buvIA2qKox
pts1ITboo1dLWxE7gjQr10YrGDMvYO0QOIQA4glfGt9nKhbi6d3kMMIv5ae/hurGb8Qr4l7nrymv
jI0lavTnMJ+o8ShW7TOMTgriCX5OXnMBIJtvrVqlpKqLjXBz7G6r8HlfFs2SiJZmMIL5N6xG6l5l
2eaDI0IXUB1Exi2E3TaC6PTBWejRLSiyTeLYHZXIAUDq7Y1WUR9oGwudyshu3Y1k4sASzvtjIgcu
paAtu8nuxPqtrsL3eArEFmU9NV+lJnIrlRPd7Lk5rCwk6htDX8HWD+6rwIcUEN4HwQ9jA3Wp/db5
R8UF/4Oo+7nbbLNtziFXxGRItJtTPcYfmGuXGPZ6oxaRrcF+5i9ZWtGikVgw97U0PHO1VHUgNU/H
iMg9OO8Rt3+CIKoED87CgspMttQGKWaMyvpvM5AcW+JRDiFKrBqcINU7RKAB3qMsH/58eN309ivh
066FA5waAy16aWcGlxiQ2SwIpMvHhEyufdFlc617KnixHglo0fxXcip9DlylRD4mQPsfL9oX2hGz
BdbMRX9ctnhvGf0qI4gD/UiCJbBcY4ePobitLcYXj+OCOryCBLWkAyq2XaBaSHwUNLIQqNyox1af
bEerDOwU7Y94Jpvh0yBPz+RlkgvDSckYDE4jYgDoMtexL9Y0/8Jj2FtVALE0fcFZbCFJJ89rnf0+
UytvbgVwmAA/jTJVgXibq+7O5Vfqh158YXGa46tdWleE7D8M9aA/RCGVAq41ueoa/gdp/rA5aY5+
FluROEoo3tSBkV3BnffVIWOA88IInTUv+LbOZfmjbjdjhPjNRRsvYcZ0h2Mr2CuVf7mM71F0Gt8i
VeVciyQKMVG+iptOQ/0jvDmgyZiXDhGeYz8eqfkgTCEBfc1EECYxbP+P6+qXl1tumTU81EaguVZW
l38hcOQ0/0PwfnTpk1KI4BleSGeJ1J3xMWRh2kz7ondaq8hoCo7iQAeYaBc+AWaLpFmjtHA9b6dC
6hzEKZPO/hw8JgwQ4OlAOcaSA1worrKXUB4gkyAW/tPBIC4Ww69GdscwbAwoulEVMjjmPw4My0Ca
icZD7GEH6n7JWplBpYUiXVPHqQBSjdmhvM3ISH6FTdb7gHcYNEAIYkxT1eZUMItl9rXMxGzEhdfr
qy5/xfAWIqyGvq9teqC251GjTRzfmHCPR/KOQuurfjZLo0Zf9hOKF0hvjhZ6s0Ynpbi347FbHgur
ACArEYGalnSPrBRXjDvkD6xVCCyXJIxwYPPL16gt0h2Nmci2ehsPJDHU6xPkUVbu9h7Fyy83S1ME
94P0NYo4fT/lX3an96AKzqT/qLUX+W7OT/idgJiY0Z0Be2Vytcx7xE+6VxaNNI1QiMcashKCekzZ
NTFGg5A+fVQ9Lt/OooVo5r3KuDHYQRfbKdhbW25SM7/Il3xVdKZJJnZt7u0Lw7D5TT5a0DQZRjue
VjVd8cHFPEcsB5QsecHAoagexv1Pdxp8XsReeeCY3KepFyH2rQseN4tf83e7Imy/K/ZTVe/c103L
O9lgP0xoOnajwvD92PVbPuPA9bfqJ2/YEi0+KJocMTY5EdwLIBG4LQYsfpXL1qClkCNlqocrAuoR
2qdzckWmb5GNqW7rOqJ/TKSLHyNByOe+ThuO7UM6JPO00tyStvrIG/eiDhzaeED8Kdd8QyD4cfk9
0Ttl9qS/+6j07j+yXpb4sw9R/Y68pXAAZMj+tApQyiCgX4MjMhrPYV5NpVql3OhnjW9d4JwUZpK1
TF1wWgVJsChT/2zx9NVIGaSUEw62hLEEoo/QxKvKblAPLTjychGlrRA8+NgsmbfZKzJSG9YKB363
3m0MIbAlSVK1xAL5Ra5GQ8JBcEfN5tUKglTPWyhs9/nh38StaUfZ18smB74vd4sFPQ7/a++bCNjj
koIgp6yzolWbkJ0tJBq5qsTy/zztuiTrI7+wG6zXsGGUmF8wv4jjAPjrbYd0Wqqc0NiPmsIOVGg4
LeTXRpo/n9E4FFkbufE1Tmh8e3JerY86RSlTqSR9dAuJGq+KWshJNkfRntI0OJMhHHqbllkMx1wv
8Tlbf8LGNtwEkCpdokT4uzHnLW2xh2YetR6MTY072+TiLUcSh/H7jjWXIMu7feEmYl1xMzFwxSQW
0URjKMsGSrTi+XR3jFpeGqfwK8rgZ2zl7gWUnmqVRjyjSP7+8B1EF2cP2c4p42hCaZns/oF2o17L
eufMJiiyLjHqD/nJEmT8D4l8m1mF45XHCMJjZR9mBZm5x1Akt0v+LZ0q4S++wQkSLHTwwNBS945u
7HlKcgXpi4rrTf2YXMaCjk9tf4tZHzRYtZKsnfGaMw991rNI1EmhQFUivJeWSi+0ggaZdw3dyF+z
JPscddz6ahMelgT0bUzB+mYjwcL3AjeqdSVwu8UHTMNz+NCDywe/c3BcbR053OGSEEITMTDoPQQI
PdNe8colHi+pH+mTR5ODRJwikgPRO0K2G2q4sIxZzwWLoNMpjzFdM2u63IRJnAAHvChrH81zEcyM
IZMqNgQvGnfqXsGy5A5x66ccyl2Z7TnsMhUYlgfOJ6JVq2BB9+YC3Hu+5JysnkLXj3d8z8ePECmu
TUcRRDoHpuPP4Hxzofm1I4yh5KoqNk0WAcsWoeLvPGSyyXHtjbAuEpHPX6cCl/4HGK/chiw0hkrj
EdEEgmBi4vZJJ8OcmwrhrghVKGy3x0cECybSMxvQzUWEqMix4sxXWUk5DWfFc79nTtONHaeEagCH
1h7DPJj2vE076FbqNfxnVvJge6NcWvbH7rcrN2zhAzkAvBL3dOe0i2biH9eJp5TQsWtVpgYZcyLl
m7Z4VDHMxqem2SPJhrqIceE9Pv7ycbRly5iN6yfw+qf4IknNMdyfULgLZkoTvvyBD9euWC0FVswb
BxNiitD6NjjY1gkodzvvwETuc8dltE3vJ2APpVt/Cdx1ccQTShT56yn7fT4jCXhsbhjXcNCzMCye
6xyWIlTlX9BTblT/1gi9qoGdxGbQvfxGve/iLUKTsM4I7ObmJAkiPiJV9hlCJ1fDa03XTcPNVUKX
7cyqkIvIaFZ/CqC2iScXIQn6MZtKXlKNnZBLsNUN5Gu28O9KEWFn+E5zlzL5/dbdTt89dxsLX/kO
HYP5qA5aIry2nnj1dvlWMBdWUPLKXNGPoGBZI76K/lFZq2fkVUD0+zsVVqk0SUY+m1t/rhtNzhtn
RN2Qzi2c81NPE65BzcKIsDfIdB8ZKwVPO6AIO7cbf+k2Gg+U3r6KzgOhMiQcBTFjys0ktqhhxFYk
2mKo6OJ6jVjb3QoFfytzd/mteXNCYBIM0HZRzdNagASviXoyrCIpGX5hFx6hDabJq4u1jbAQHHBD
tNaeSxlV5fCeXeN9YBiCfFQirHlw2fDerSv/FQxjgynnW99oCsxQgb/m3/AuB79M0ymZMbpGjd9Y
uUX3qYDStYcA20npwvF8OXm5WxQJZgGZVwQheLlRJe46KqjSsPqoWilQ8mNB+rNrfBTgPoXgR5La
dzuzIhdFCvND4+EkVpZN+aFHcYRUt59MDPx+lbCCnGIrf6V1F03WXW9j01SW03Yr1HSUEFCDx6jv
8cW8waC4+BxC4BwCD3q7RsunjFBKcCE5kn7iRs894EQ81wIGn20xuEYJfFRHudMDnnhAMEpab3Yy
rp4Pe8dKI8zcZBQfdAU1hizPp6CNA6kNCf+mloQ7dpl/IycjoAVLQ6G37cNrfy8htK7O2nBLCfOx
GauEnJFeQxiyeQWiZZw5UWGIY/IVsR8hmkbSAfFRmNRThBlLY+xZfPN0sYucscUkYUS2phZmKpIl
ZkyRKRwbtYMSITOv9XEbK9EgtirZXOrmbniXe+5OBhn4yYSCS+JU3NdkFyxJwgfhcvg8tSfA6pE6
9VnDnrMU5JvFshBGrtdXrsWVkKXYmr2bw+LkvovWT3OgBL1m46RXKgBLThEeTpTn/aIQVfVE+72K
jEBolScbfEXRX2sMmnDRVonTWM58zXHaCBmZV6MpILcoJ/cspEPRk377pGGTEZn6p25L8Rrsdk7i
vJMmwuwRov2WTTwufbTcL9nfggHJsD1rOtVhMPutx+DgsIXWoydCOt0ras2BFvuI4HqfRPix9n49
DanLIFu5F1zol2ydc3Wvi4N+G2dL57F3qE/6oe1Mf0z655IbUvRiJDBY0yXYcxt7JYwy1Rw/wZOw
WbyS9GdPcO8PbZNGhRT4EEKs+ZNBXAmzTwV5wSFnUuaGLkCabI3GRwF7m+xglgRNMNYrEyHYN91K
WL8ruWUASJGwWFgfhKkWAbs+TPlL6ItHPA2yk1DeNWlXVVRarG3++bmWK51trZXgjy6hiSCJYGzt
g8xqfr1xv2lRbZJO7bG3FUbIJCc7aDR8e1DJhRl/UBk48pqEpsgkumjf0yZt5gTaA18pkfaDM4zA
pHQ7Ym7PeBPjOKMBgRroQAXNvwvUYGK4RHaTzVIeXVkUpSWDmJ6OxYNWPBuCqjaol6xdh/o8Mr3+
FnDIZ+nyjfslA222yl7FIo95gc6f33EeE3/VN0AHvxuLMjDaMRzOTpsaKig6j1EQGMOTjME1UmrI
7jReufCqHryLaFIXMtuZMVIm6yatF5ig2NtxLZ6yycGLuw4yUESF3yBUtltQlIGyXKQzuzfjy2le
IWmdO/C0BJKYcgidP2H3CPRa0GZ6GQluigWaktm02Gxo0WroT+Cbzl3u4y91R1fFLcXmYBhDHFaT
043RnIbfsB1k8TT4d+nWEH+1p2OnOkBl0VkDOyeojvl2uAI7Ag14kCMTz1Nh8aoIwINJcv2xU/vZ
ov9xTQKTQxzGnhDqnIdydJkzGUW6Hno3ZtnUtEZRFpB/S4dzizhoScncwojBZ9fsCNFXHheyIVKo
0b1duvVKDHa9KIRbjuFC4yV1Rzz/ADOfa0GTiZTL+1Pe1sXTCFhq5xQaXQ3UVFC/BXvyYDIaXFqc
l+Ro/+Ef2g9umQSvwnhblZXYuRDm+VIcqTk0B16qOJ6k/YtWsxLgywqjPqmZ9uftEbvRr21sVaRp
HA40B5Ka2Wne6R+TmfrcRDn1+mit8PVFAHtJXocm749PGFOVmzpC86OwM06UbgIZ0MoYveTFf8+t
tNf+HJCFluvGDHLEXihb1j8I8ixk1DWs53FBswJHF/hJgak3wV4prdAN50Z8AaSWagUP5sGz7j85
B+QBy+JoHMREhaEPgo/25MzS+JwzQIyH7zG/aYsH1ZN7gUGcDDBCz4B1o20OzROW5cJNUU6NMZ7r
WFGYxwLI8G06/MWoSTMJdH9G5LYao/S2fcq83slGsLBm2UwMYl7jk2z3sOUpurDurAGTDHrhFB+K
M4rTXxlLJcbyKXkE7sOskctObhjt/pAP+KNurd8T0ecjKIxYJxh1xnqoSoR6B7UfT1xNRYoqj80g
qFQ5lPTOXkQgIGJkUSNOQ3tRj6ee7yJtOVefdPf+IGKy5gCJ2UMkpMF8fBvEO3Rh6wtBfSsJ+E/W
LC3Eok0V+5Qa8fuT933HczVeXYc47pvANZvXpQ1sOOW+CBRdS+BLnLFk74lljzajgjDupJ7iaWb3
/UCggyrxhM6qMiaqzBN+JNmGbfS3mXrEALknaITJKc9TmQECpw8D4/JRt8emb9S4ooAn8uM4kxEn
+N2pQ+7na7NjxhMSXOOLy2QFX2X/qBqyN6AiQjSKt3Hosdtw/WlLuCIR96PdQqn7v1SlqSl2uGdd
JzrQEw8jZT2T0hOBffri3VGthjd5ulkpJTRRd2DB7tUQuJS+9cxUQ++Vas4nQ5CU58Yor7h5u+F0
YOAM/GaeHIvGDTvS8YkBe3Z1pdIMbto5eSJN7CR8fpZmYy0uaVSKYRB4AU49AidV/mJqQhVA7Vfr
irbaghPbkSXK/w+2dRPBb/RZI3ZS4wDiQ2mXfk+39JoLWzZhUr6Tgqkkl6RsqaGxBErWeiQsHain
BxoYKUmn6S438wlbmyUql29+MBXe0EDUyXxn4npN2ip5ah/idd0T0ysDsentuRFJqd+7w8Je65g2
e6TA4KMYaWDPSe/5fTKmiwUqi9GMXkjA8wMgWZtOd2RLpJSZULbilKBQc6zZ6yRDmOWdXXntHErW
EIJ094QrAMEO7MziRpeH1KotuzpFERiT25MSCsaohCBjRy+oZJ9F0S53Ydt3o0OjlpYOYD8tqqJB
mTOYemwWecmxh4cO5mY0+qxB3INw1LJ9hNrh2PtnWAMalBZme/p2kg4L3bGfvDEUxea21e2z0/Hz
8oYvkUm6VGBf5p4GU4O8neiTjfVjTYDgTuYkK/cgTAqsyQYzoHh+nqiA16hT1hZLsh7ELPTjs/mS
nW8mkQER3OXyZ22MCoZ9r6QLQfEIqxXRVcrECw5bw4y9D1FJbAoz9kDuAthpckL4HKqDp6dj8S93
TLNby/bF63PxQb98vJSG8MkX4OrBnpprUc2klEgpskWOaJeYYaA7U2WjlxftOi10G7mFrGGJLImX
1wrgA3vNyBhYIkOApTagbed6KRCPyxjI1dwih6S6VCqm6mGclJwj3K5KrFim9QcyTuBtrjd5AuC4
ioMRwLNec1Zd4X6Oi83eU5ZCT3DTOagUA/4ki2uVbSa+Thnbqs9ac0rbSEi2JEDAkU4Ml45R6TUU
n73EKDwefXqNjpKbWFWyWdBHXuxN+Pu2q4WsQLFhB6lsWuwe0OpMLoXmczoon8wzKaNmKDBfUaTQ
AaDCRf1hOkfDV168kV642vhE4iAc/skAg0TGlsckY/B6GI66zLS5b5fPdFa2z9oLYWCIOcP6Qbcb
kNHS0ZzCoog/yZDsCdkygr82QR13uAscfOvJ5bI19PFjaIy09Ma+1ADKZdnMBlNIFyd2CBwqGOtP
DhnQAXyPrynWRfnMhIIMUrwqZKgIfR+cI7pXrdJtVxf7ojiEPeEQrEAhB6Tr9AKrqyW1ESVDK/Gb
ZYGva1VT6a/X4c97mTVcBNNEJfSh0cYmbPMIbp7Cfw1Wmq9oUoPLA0DHUZyLi4RLeUtjKb+tNGrB
LhsrhNdpZSONUZSgfHj0UyU/ZjgFm2eJmsjP0C1ox67gzFYGeL42AgM0Bjv1giiv0syMPh1EQcCE
FP74Zfa/bSOkYRIXbKdBftQZH5PAU+LiPcU5TBQI8EFbg/UOQvPWlXusrDYjGS4oM3t82+0ahR1P
0ALTk75a2hb3B5Jj/otiR73klFMIf9KbQDNXJzMh7vlOxYplQ1mgY1Wx3t4EqWg+jNeG1X7QHofW
CaMlsWmJWTyaXgyhvxFRiS+DY+IHGoT6hfYX8G9Jc05+sMFWHyQZL489uOX59eGNajA4iw7a1Vpf
IPr1WchIpO78zUviPObM2du5T4+9+2a5Ql61SjKTijya6u2j7HIPCJv7y0Zm5Hw4SfnIT/eg56jJ
RR+fVF4HmGBirDs0Ak16xURYMvwj6EYnj9CFDC9Vr+jG+9zAYAXFsQT43ffvPa5KkplbEDOOAx4o
De2m1+lKjgRWDePc3Jb2CudJpuc5cXilC/f+1VXzCX4U06cwcJtnNYNXwn+kvPpKVR8dtKlGbu0E
rsbf+hwCgrOrblB0tJvhM5IzdWZvWLURAGCXhLHdGtw6ju9qWcLtLB3OI+KGsb8B/m/1NFOinK/6
tGxP5JB7QLaIR1V3BZHpKIjlI2jKyiTuZbOPaVkLVJ3p3Cn1I5GCIlDB0lkjZK1eOm0V3lt9f8DR
qysfxvS49YiwQXywJSOQLNHHvwYhRv8r50CR/6dGz3QGd2Zq4gYE89r0jaWT6+CesDbhsjWIqQAx
u+fegVl5+l/wTNb7gzV8plD+t6hmzm1iF3rdPh20vLRgetx3R3OHXTRxszUEFjkVGhU2lb7ZOsSL
gKKSfkl4q16dgApC4vg5Ev1+wd/R1Qz06CBJS3JxBvBx0q+f0v65XHal7vguc5WGHruHhldw1PMN
Y5+RwVR0sw5b/ktH/h6Mibn67Kzyc+4V3t+R7Vuu1fqg6ST4UqQYG8UP6mbFPqgVSwQGpTNHRSJE
VPtq9b6obHadjsuSSNqMzwTtnvJO30NDjvAdUpnF5EStg9CCCiO0kUjH33Im/HUtH03nbsIAeBVS
mABuORwm3/xbBy/AziGI3ayPXD+YPcYIFdS5CyYl42q9nubyzsfaLwSCukLgcKv7HBpx2t96PXbR
XtrD5l4TGVp9ZS82PwvUC1aM61/8ae0FbPVF2exF9gkEylpi9+0NO7apwezUC521FbP7qZndFtwZ
vI32BMY7u1xKJVbx+BNSj1cMN2YN4QTPOQcjjpzX7DJKpPKY+Op1/BhyvHXlVg4Jk64jDD9uoBFz
EH/gFgS7VkYtidemWVdegub/f3rs7CRJnRhUcfvIaMMQSbKXr3VAExkTuuVDb0qzf9yjmna0n5cZ
MniKPQ3XhPlkVoV91x+qgKFdXPYzxi2O0a+JacxQZPoP/lDmo15Vs/z4E3zEga5fA8s7WUKyflIY
9tY58s+sGRYDKDJ5sPX97c1HXK3sClCwPGNAkd/coS0rYvrHubICg+o9FnWQ1q733VGBQvkzuKx6
G6pJ3oqwG+0UHWKUVwB1oEt/yIKs4aP9Gni5+Z4sTX9BlbAufc0wCQCyeF/xsu0PNUsVeozgMQtl
uH30PYGexQ1R8PMDk1abmWRC+SLF+SoizGDRUpk6PPwZQlz3MNiPWrATU/IMKHsnZpVuZ8HK5mKZ
R4zZXjTJO5NCe/OA7ziHOApmamADv3xkz4bw6w/dJOhUg6GP1BQXTrEF3SjtfSG7AHLm1B9Nv+t+
WbhKydNeG3DIjC9QYtluiOhqZrN5TjSZHcpf3RbTd1BjnZzi/F2jpBNpJstHwL362EqPw5NEYRgK
aMBpLlVzwle9iR8kRqi8R0ti+u9eJAtjwYllJos8CgvlJ70WfOjZOTnZjQb3vW/yDVzCiPfEtuxl
HoEpa+0PV/BvAaMzRh29juwww5a46blAIbbGVhkVRLVzPX+t4Z17F4e03Ud1MP7uMdbl+yND9x9P
JXO2n1LHG0f/Shew+NbhUoEFMhbCtggq0UdANnILp684Fd8hCA3AnitZSrpsLR77o+Jak/HHcW5U
YXaWAR9EVbGa8g/h6q9ZABrFYendsFngvGtc7lnjHCjBuM8yAaUkj3v6A1f0UFvvQnEuvMSXB0Uu
MZmlIElvswcEAnN+VTNmn1mtiQhA7VoS/Aa368g/hlc2EQjdSgqoJ23Rh+GxXKuSSIWmwhs8SOSU
XVK6nCKS66OkSF5G7TgZaMrfOvgUZ8caN8vSupjvdsgEIUaFLpbM35xsdJwLFPBfhVa05jZKZop2
4enr8+3N1lFYqrsMuSr7IKg25+6hBCEV7+TbPr1MfHt8FYmZuj99Ht3iPMpl/qUxqZzGxn5nydcW
Ty4Y6oiWxRkZuSpvg+stQBU3v5rqyb/ABQEHZwULSo5/sc4295HcapTpAaW5Z8407FUYyiEXpVox
RDa01znQPTWk0Xf1SVWp9kJlukkFijz+Bm3f9BWiKVF4pkx/IpJ3hOXqczdErwn1TEK5igRpbEgg
R5Dcm0tY9gqOsjr3+Y5Xtr704RhT1M5mcFewcOECro0T2o9rImIjOzD+ZfD3N+hcOzux3wrCPZhk
fmyiYoiaZ0fJyz02OfypE79EqyoY74hLOHsBZp/RFVMFs1grJtmVlP/0acBaq0GkmbPHN5K/i+lr
DfYwWauVbuk245YNY8bgpGFHT+fPcQsD1468ifENUF4QFwViNTZ/koSswSgHx8NS71jNWQ5Wa+IU
ZpV14DS6Ig4yhJeYid4SryvAeSMxi0X8uP6xOoawTt/Zq6FnR5W6W9KCC37UAfbBeyXVohroipBD
oJ2NrF6sr67gphUHTV9aZo9aB804noKLNr8UjwRDuY0QOjIwZ5GpFMmfclzVmENlBqy3VyprcMKZ
6OSjmBQsIH0sVHNn18SeqrMnRB75fC8m30MtprpSoryiLCUpmgPVHuVOOt/wTkZBFjeVVqmPwo0O
lRY52d+fSW4RV2zb1k7ytXvw5aEXAUNsW5CQYHWhVyxNmWHcixj/huWo7qv1rAI5E7FKHw4LCzIg
vNdgHtVgmsvgR0l0RGEhps2furBMpjo6u4mW3KOsAE7d6EKdqtSgxgneFgdrjg/QRdJYF3h5MxZN
Vw+yGtOEbaA3xJ5Ci2rXOLIw+/fi6CFZ9Axa1kf45g4pNGIjSkXhYsXX4kiCZG11+K7NlrQn+4dp
1LnEwY2eIEjikNdWQx0kM0+gw70A+mVFoRVXS0WKoUoW/tZRGt8EW96VSMAI4WOedOciAwsNApPS
2aasC33IU5nzFbynLpRxq3mxA6XEZGep8Zy4tcpUZCNUKLuMJMZ4DAIYFU+ZsVdZinVbBlZ4Qcxk
UkklLUR0PBdkol9dkoGbFn7JDONsD74zAWe2XCgXWMu5cGQ9rnipdVH4mOQig4fPtWrmXcQrmsAL
qV3cHCLD0RCAOJ3G9tW9bwaSnvm+3xaXp/dyqrZSVmtKWJlu2A4WG1POCnN3r7V/ieaTLR8nb/rZ
jeIqnTmEiLCzec0fd85VP+cfEWf0zI1uSG1Gbl9HL1zcfS14JEg3PX37oBIKBqtL+dmD4leOHpyc
IGZEE1gGtitOmb7o+OYBBpD2h3vWfYRXg+A5IhX1X/WekpZG1tmPItL6Pk/p56pl/nUMHDqZyi0Z
1pTRhpexenW6K+qd4MGLSsc0HsU29v563WIDqftwAoCHwsQt4osBIvEoOQaQtP+10meJ1BvMYEPT
UywN+Ny5ZPABt7AgDynFGWxGDlcQYm7g1FvANhl53nBJYXBeY+BKboVjUnDltUidPbeZXFu+i4Kl
YhcpKf3n7gGTUONnINBnSW8BZKGBw6OwlLsxCH7FBZEiBXMfzyT8AhgP4o55wqp65JFRQdUKUIpe
iDYGc2hSuyhkgeRR8TsCaReAxeu4foMCTWKjdA2GoSb69BwXr8YVIdwqZ37YKo+bXe+1BjlNeywl
W2M5ZEPqSvZEJVzoH1ENdGiXTZ6xch8EmOkc1gKutDfCcyXrRF69bC97NnZsmHNpRrdZzGyAnjTu
nGDjyLn/JCkLJD3ZKWR1x/npVM7xNHEBaR3ZXpWGfMud2EsRGakcpWsLH2eqzDPVn9mYeFqE1jWy
dD4zfMZkJXyRlKWOJkk85/tzILgP4WKt/1mwTV/kO9XIT3xk1bXjRrh/t88KVwsB2YwpBWMwIVV+
OG6RpV16A8iSg7520fo9sj4mtE+/+4gT0O0PSa8If3VYMBu/96C2uVrHgn01hKLdkpkbq36DgWcN
3dPAfPzuNekvTy8ZPZt/pXRtkp8zWeim5Vv7xaAJH347D75mvsE3M+g+x/xiLOnR60dbyZqIfO5M
8THDODx990TAOEC2SpX+vdjDI62MAdsINMRNd/Cwnue+lpZq0gYshkcnm/rP5dVt2k8MOhTJYh+D
yAPml3cUQK1fTy9SqVUuhv+BpiTmY48UATthtEEH/a1SLKpMLH3pA9LzX/gNug/a0Vko4Dsn0mky
8LavnjIHU4NBB95FcIz9Zwm6p+C0aJf/F2doc4xpC27/rrnilaBAm7ALJHmbYOKmViORYfQy2maM
6eEOjr+o2CZz99a2gNotS/wSRM7NnM/aLmrnxIdD9tzIIHHIIwACltVbXX2Y+WMLBpfKiwh73Rzy
xBTDNDPh9n/CfSO5Y8Hwo4QDj1x/U4p1GrO/3ZVebrcrqmZP8+haXO7tJTWE8pzImRzqz7Uvjss6
AiboJYNhR4xCD9O0c8Xpx8NmSdXKf0VMn1Od0N3ntuCgXGJ//S757om8g0XqGb3XBeUapIdNpJl9
2sO419zivhBwtwVo5ht7edYtHAXZHUydGfweRRV/4i+6QlpnD3s9JH3zpoYtNzzYthf46D9EMj5O
ysQmo9nfKMKZ3fFkmtABYSZ/CVASIudkiMBTGhBdsNqX6TznnSu2IQAXqbvXYtWJ0jKV6RYt74kW
R2Q2OEaGFiOmG/pPBbnW3eWKDH4x2Ny6HDzEa5Ck36n2wrCEBy28zScnR5hxGE0NvFpldq25X73k
1ZNnaZA1mlJ5lZE7EG33LobQHRmsYmWXL3i8vdvMmAFzQJrcTUi49Bk/pjK4jpmWKoqU7e07K+xD
Ny/q47ErF0bGF2BVX/973QsQaSSeF+6VBgXJo1509VlxhZvqz0RHskCr+LoB4qjk3z7q2LnXc3jV
XEs2zO6NL0fcQxQlRMj8ZoqcAQx1l6UJC9LmK3qPs1ymvqEd+sLPwAJ9aEW/gi2DzWuDJkg7JUpr
np5TiRk/M7Wwh4WRuvlQ0E3jX49QlZNCTXU5w6CC5Cv2nz0n6poNPmSox49ZloNP4mKK7KsF3IvG
Qt2A0yHV974scoAzq252rzfw13ITpcSQFsJmWHHPT9ONzCu6IC1EbBA5aWGGE/K6pNmoj/mN8Owe
A6+CGCBU0cs1bRLNYtX/xZ8c+RCwXv9CUGpDYYdyBqkdhLWwx8E7VIxccg1qX0j/lNP1oTbQIdCn
y37ILKLD2kdQ5Ca49ci0EwKTqkoV5vvFA77ZvPxf/tgaDvLOw6jIsjkT0juxb6LmuNACCyJ0W196
/xQh4YzZySxQaMWI75Qd9YD/UsEVJ0GMKd8YayXh6twDkigaHChXN74FM4EtVjiqT2dzSqT2Z30S
5CE4RpYz+gSSmCAa6VtFn2mWIyli92MfbUKp64MI7rs+hzx0oI1N85QBxM1Hlc8YNon55D6x4RUe
yPbjEfi5A0iYQ06WjPj0rDWjimY+D8d6rxggzxPe3SYRhGLs1GREzgou5zMw6ZWOhAnqB0ikfVT2
F/avlP7VmoB0LCoIwNX3MjV4mbqcwfylgHvljoSwV+VpJZMVCs9KJwEh/7RNrAnis3U9GNSKnTVd
WR+qV3+3Ay7tcZLyrOCbwAj82ja0JdR4yaDGQkWhzeGpA+2k83woR9hOg4DlDgQrQWBf2YKvqu1O
iNl+EOtZ2BZv52MlIvq45WYBmQR/35S9cZBAnmxHjZjs3tJ7y5Ab3Yx2YAJzv5vUtUxX7pxsIXB/
gMTj2lyOOKenjiCxreBphjR/Djizxc5iFw9FuFpY6VcUi+Mx1ULeVJKBytFvjPm/Qzn/JIxV8Mey
0OOZjdn6rTeAARm8ZZR6OEcbc0+pnOepy42V0aX5kJTO7zdhGCemLdEb9BsWUY3TGoJEsDDCASch
zJbM2JQTgHVVRCNsKwO9WBhr9babheMEhLTrkfPUxiYelk4Y8z7kSDtVYO2dDNPSFiyBOQGywDVZ
z8k01lSbsHVwItaivP0N8EpU+zGY+q+tQ42kCP4O1a1/Vsdizr3QY2Gdde105gymVGkgF7KJS9ak
QJLjj0g0UGmPAFlginq48ox4GKk9L8O6F3curIVySG+vo8vDF4L5CLIvf3CBdtTQVRRT+dBMktBl
pD0AimM8ILdY5dcyzcMlz/R7LKouwODF9KT2Z+TRrUc8Y/1lUXSQgCARy0KoPxDQf5sMncKcP+yH
eDb9fVoMhtrBf7JR6etJ87iJCD/LsUaK6L7AxgyDs/QkNdRa93pejp7sFUvZZezvA2mAlTd1/pqi
K6Fmgn6RZhP8wTeUGhx78xxG6rdO3PiDTTjW8slhFAgBGp/UzUvIXqHI9tPPPs8Z69DX8wv6erhq
fQ/3AzB0cN+pVwCFiwF8ne98bvEr+104dsHIVy37bms7HrTJLWKiG63S5xhnMwNMkKpbM6Xyfzem
XktMnmYPHoXKoyH9GA9UWEJ/mDmd8MfDpChOt8kHDJE6Y0AjQU110/UTB7636i9Jn+aQHZfcaALX
CuhtvRq26hktuEpYAsHCO7R/prxzt3lQb1SzP0FoM3Sj/iajvbFOHoijgxVGA8mI0SsLb9s41JNQ
alanWSz+ynTxDgXJQfmwvijOByk1nxvY6Nb8f/UXAvNTygic+6D+Ls86Urd5fA6iUxxvPKVICUl3
Ct46KPdWx84sO+w/AS8P6O/8/E+XF/9gCDFbyLrbwYS6Wiy+F4eyb/607PiEa+8yx+1u9Tomq/Gi
b0fJPvmcwMx4aGuZuTW/I93dTR1nVk9jjbEYoVxaT3BNMdrkZjYKS1XZ5SjKPoVpjLOoDcK3CYZE
91wNRpJtDEhWIpGabVP/31+ex96J3R9z2hSa/oyfp+FHSzwfpk1wng92JlDV3p5y94PclTqPsuDC
AZX7G4MqLgeuUcSmCNki3V3uuRpujaU7sbRCe68fr27c8OKHXFlyzFDKIPAMRTKU3HmWhxLokLKB
jYOYE5eIQcjbwTuhDjKetef9OmMdUiL+RVJTnndCvyzZG2jVYpCfVUd/CL3GSSqL4ebI6s+0mG7P
BRz0ek3MsJRHxqHUKt0q4EBrMeLXO8B7bzMc8+flIwhfo/WxH7h9BBZ3k8fvh7Jb9v6jQM39pzu+
DdN+KPE1HS078vtwn+JJWtWzIzcKjOdiAq6Qd5tyF4CapUHZyZkdHp5Ly6oRc8oHcu55bIy//P7y
n91zM3O9AdmDd5cdaThTngnnS2qNLYYTpbSV3p9oisGwzQ2z46xumnRi0abLpymbwWiqVvj5iQ+3
aDr/bmQMsEAdq44s8Oh7THAMldlM1SeFrpanBfA4S8hSGZC3kHtCXXWsVWM2eIHcIZoA8X2oOQuW
EMXkkGel1cdaO+IECL/+1y71itLMNm7Ukn2pet7oApOY7TltwRt5IVEOvA8/2hEe5pKDhop74M3J
LPeHZNKfrQbaMNBoIO7zPO853rX/b+CkAkNi5jsQY9jJBfvRYTDj/MJnf4sBpeJFDm8XexHCo7sY
4VYS82D2UO0bNWKER5ydLF/PUyZVRnBRmtUNI0hodgaIJ1WFtQMSKuRZpCY/XuWOQ4Pc9Iap6xHQ
mJnfiDv/Mzmcp5CvQCIlalzx1va0DEtdGE8mTzSnW7l3zJFwFYT+mj6iLx25R4F7vTyEeSmf/Osw
msRAzuriuRPtwAWZBtwPVQIG0g8Fee6V//JCMS7pUNECbxkas6BoMPmaFmx6zUV61Ok5jIjXFE3N
e0QZCnMp4CHh1VgGO3ukcQvdUff693vElgeTXjJjagX5Lsb2LI3Z0KBFjkGa/MtHtI9yajMl6toq
qirFY7jMzzKvZVWJdwxVNI5zGsObdygEyulIl/r63aPZd+M6LVOZU44i4tkOlDoPl1hhQqQXC1YM
oTKworx2ehVsTWeoRzG3TP7vZTga63yDGuXI5E6eQYiFh8VeY9oe9v8HOn26swUNqGNdp36xLX13
Hko4valkh1UVqqqoPS93Jsbdau+3+JOMdi2B17Dz/812+5yIeVbaRVmC6xP0dbgtesL54khosUMv
+D22DpQya+nBV/kdRoO5+v1aZ401luDhnvfwbKfogBMrH5zuqJdQXEDuCdU6q6Tnc2i/LY5W2s5K
R+w7Ns3/svZEj3acj9Jhz15rmFKxGye1gzJHDIiwgz90BviaITWNuX55cukO4ObkDCFJEEynQk5W
i99WBPPsihnV0oAueLtEFcCBhWesgtgmEjAGbdbhhQ/hMU6OoMCfkMi9oDaJz1R/3O/DjeQ+Q4tq
v9rfhmYWIOZFA/XmV6Bc5phtSX9JH2SQoj9rrylbokoElDzvhL6o0bBzUDiIvE6adCIN8bxTR1mt
GCe2rY85DYCRSE/CA4EemCVGodMKloHAgW9HTuFh7aQTbKoWo8qUtzMxvdIbPc6L6LCCDRumrj06
T0d7KqOhgkAnla0J5HJDUlTcn9FygUnQgKAsRFq449qkf33yBhHUoTT//0z4yXVRkeu6bYe3aOqF
MJUxGyQUOjG3vh5gVNtHGORoLMvAaU/WcigQB8qtiom+OuyZ8XxiTSCoG+axFXrxETq5dUvCAq+x
6IWJ0sDwP4gmf1hfAbAVeU8bsQkwh3jh+uMLPvzWhNTNc5q4LvMkqDKh9e5YQSAXvWAFpCIdq8jY
q51LTI984OK6kYAgRyPH48PVbdP5yXddHt43D/pxnmejQWCTncS/qJjXjvcSk7vLZewBn1LB6Qwb
VtLxmJNqei53Lng2fVHO2saj1brbXYJ930/MRd48HFqAyC2kVr3bx23YiPNwLOkWD7G7cQM1lux7
M2sH7r4BCa1SkbqE+wqJPX02W9u9/fE/Qb7jWRu5njbUHgllfgKDK+nW3CEukUj1w23teeNt+0pv
cmsRDMaZO1A53hnOsxXxuC99tFVH5cHWya5wWvgrPGprITPaYPr5p7XfbmKU+8Q4cR2LE4T+rpzY
8mhyh+2w2vt3TAVdq3IYbr0nw6N8wtGg1zZx3HxG6uFSo8RNF4ALTkzA+ezKV5Flf0xsvmNTh4bJ
Rdd6MPgKBofx36rCabEvAWQ1Pd/i8v9KPsp+ZjChUkQBjnS4kzUAUrMaBQc6KzTrJZNUM0suDGu4
uo3FFrYr+PK6j6b1iedU/3CeECmBPLP+7c7HDmymcDjJBJcLY9iP+Kdbjy/ETEPkmRTjMkDQcRHH
9YCFShm44ap2tneo84q5I8kQ8R+JIcbbs00nC9dcaOzRFrlvWOT/K4IjMO45FFu6czcbNbhe0rWu
9Bn3dswoHN5zIwzs+S9+IIBsb2X1EG0aCp12RfWyqB4HdSmm9ZhzPYHc/DmnHV+oCAMKp6vgcRA6
IyIyHDpVicdB/poZgk599ae83T17UVMMj0hnL3eXwdebURoQq5BTxV3JOZlD0O4oyE4Kix2EN9Qz
57gLTFMmWyB3yIcT33fsg4BQVRdYBkPKP8TKv9aYn6jaZbkZYzS21+mAlYEIjQcfTVIqHl/b/X2D
UOh21aY6OJEAsNFFBGrRMYqXzM7uuVLj+U/xYEYBb/bYZZNf+Jg8P1NZJgPo1MyzgKmPrMmIgU3E
B5JuHuQsTAFe/DtKuJlg9I+tgHMkWRUxIQsj4u7/7m/Yz/r6DAWMPxjMcUZ6K0Wz2zgTETj2KIE3
BlOCfXQj+1in675o851XszsWOzZvkMu9numw0ZhB3pHysis7scH3g0be5nyz402/ILauEWQkMRUD
T14h34mFoqu7AZd3x29PG2tryKNC9xIegDK9QkhsTqV5vukdUANAYCbFg6dzzCoCRgbC2wDGch9y
Kgnbifdlz9T4vaOMVFAkLOLJXGEWDsVJNnmN9rnA0Jx1+h4acuqZ+ES5bWu1QHWdVOfl4uj+d+Ma
WhH4KvNc7tj92D2O9NryFjjsCJ6v+gmcg8YzSNtGY0M1WBuDCRb+SKrpYFOTcExlH4qWY5+6HcjO
NXLXDaT0FuOzfw1XKgNXAIw3P9Eatu4FjgPyttAEgvE2j10Ea/xEsJN6Gt0me4VwebbYeWfEHMq2
IxzMSqoTbAzOb/xgNxefd4BLWb96S234UpJPthqW6fkTr/yi4HNnUCIR5H+It4xmgNBeuDBbp7ev
o1chYLyMv6acIi5b00f4ApDbj9CPzpVRWlwq8F2s6OLo+lHCnpBGwI/jz+oocoAW+dgOupAt1ZYA
mB7akbI/pO+CyokgG1JoEF7uM6IvQS3fX/5kF8art+oqZtvIEanS4hwRd2tq+KWEcWBezYFy/GDH
czAa79a/hvBzCQcfwmjD4+2PomZWQR1N/hG6KuPZulmBg773Q79Gb12RJOpitu2s6uOBaetEX33p
/+7UiF2Lx3Qu8KveM35s0+fJTaH7GPX/+Jb5aeG+Vbz51+Nf93xzJbdNMCw9i0xYEGajURbqYD4l
1poafPgU7tDhzl5B+gD4q3NS6YaWC5nLmJo2V+RtEwmA8U3tEkmkROhzfeSzcyAJwIMNyrLWVZM7
RtsYSbEcX5psacZEL9mLJFuBgtQTTSw1KRX7abocoX0eJ2vvtxE4inkiHpXrVwLtDn5SH1MM1FAs
8wT0ajOUgC4ss0nC14mcpyCsbOs99uMkpY/Rn4R/dSV404Xs3SZOMWwe2T9LZ4N3f7nVbG+dAdR0
3QkA/bw4rBV9samFpFWmbbJYUPtqCwaeNqTfRlTCmzz+4uOEI5FVeNbiLOIilGP7GXao9qTA0vI4
o1zmOaJPobYxglNJeUyjVWT4n0/0n6d0rLgHOT5Usky3XDrfXGMOYiAn1ijXTnwNzEFVbvnAZ0MO
LIXrZe4Pz/nPPBG3QY9B0rOCvWui73fOaITZcIOw3u45n02eiDTSktRJqE0W7CzibQT8fBkSJOXH
d0154hNcUgF7sXi5VDoXKZXZIP4oaimktmukCLQ6fy0ar/LQqjogo/l7MQdDt/KJP6ts2GTnq5uX
+mITtfTc74TWZwlhna9GWOHRObAW8TOsTxBmSlr/GOhv5nVtE+1RZGBtHC8fp6BKwJFniB1Yzs7x
nCKXDJewhO/EfJtAQOdf0fqP1GFqVIU1GVWLo069DbELqydkVcuUCL9EhiZF7j3ahVy3SyCpEO4Z
+KfY34z3ZyeUwRxxJWNzlU2VW9sVyVTuzUN7hiZ1iJTd4skkFWl0mGa3tB80RY1dntREl37VbCpd
q5a9/KFIDypTjBhTHDxHpGi1HYQZkliwx0LTLwyoE4rgz1U+kXjTwsu2WcstzsMMY69O/yfpC703
+skqttDzCV3KfgU8yfs5ceJ/31hCOQMzPbzSKmZUMSLUlQTvYMYZG2zbS97LN72RDJ5Ha5Om+Z08
bqFlzkWCD6XcgwadRKAV/bmpNTvfdWi3EZn2FgrXNtOdMQ4TcWnSLSpqSWRcDYir+TMTYUbsg0jh
OQt8TjLJuR+hAk4niZskTiVC2ZeX9KjyIRUPvOPQZHBMSx22AagNa79vnXvGqEf6PP6zwZO1j70y
awoAED5LKeCf18QiG1NfrsYKxhnVDA9/la956f5v0ZS7XIkl8fxlDxzhm58a9qSIgu5S/HsVPIow
TMlUZWwM86gUmk1p9zo1ClHGN1QxByn2E2+OJV+4jf2HQbwo0XEeOA1Tb15G7Z6wWdb0/6CJvdMW
Eh0tZMHRsxjshwi45/V6CVNiMTIJlnM5isHRm02Td/JjRQLQxAdSDmnKX1UY35bgcVdLu9VaDpRq
gybfxNW4vJvt8loHsjCEkfiNUxlZZ2DmU5cHkO0ohQiQFRBglw+wM4OTB7DWgiVh+527EcDRrxD0
BKAiIPMO5GU2h8F902Z5OmGniTjSGUys8p516JwHYP1bzsh8MfWXdfD+uUZsQ/u9VNpN7/EFyP10
onpBOvdPSpPc2m/CnOCSTtAjilsvm6SW+0a5ItcIM452jKqbgsOe2jfkrnCu9xzpNMXdWKcn2AU7
da7eTIHo1wjkUm+LNGvmQP62pW0ovUtv3FVTqvgazxUNqCyICdb74Gj0X3UkqLYwh4mw71jLRlEg
UV07iATKbI9xQodY06255avwdu0oiDZa0ny4ISA3WHsa9EbwmvJx5EnSJbCXCqX82UTh3zXJJl2i
qCU0PqKpftiRnCmn+FubxBY4LWGkSBkAgpqQPuLJB20oNlOKn2y7uw7DMeDYsSnUbTq22ri/+Ixe
XKtwEICOKNma+d02perrG7klHunn+nACZkxGcuIJL8wGm6l1QwtNBzsI0zZs4tykGq6jBEg3gvAI
PMLiOIHExOJX2x1AUQHFtaIXwx6aRqUDda1MI9uLcfgBYvA4ud776zd9oDDFT4vvg39y+deys512
OY2BOG/SB7uDOA6u5IkVHT/DFfBDamPGzYeKXn/YpX5H40o0z3xZfyf2f87BVtXSxG0upbWLlcAg
ioG7wlpFUi/AHVmU0T/Auyg4vrnprhQE3Prkl8ONzhJOJj+TAUTL7vgohwWfpwxy2a6ahNu7+VZf
kRw9t/rruqY6kLhxPNxO3ggXQfwN/ZfX01kgGITMz6suAm2zdebOELEOv+dPH88N2SZf8e+XokDo
JDVWOwCTCyl2wgxbB8PegPXxAY1n9CbdaPUXn0ytwgwdPnRotm1IAEIO1DHPRjycCv/8O/+/tMgX
D5+8Z/nCut9l7T74jd5eOpVbDW2Dg+fIOTf4BUhSU0lN6/v8UQfvCOIKf9IKNM2Spum0v974r6WF
HUcDBHGe+JjdbO2ctW5zp9HaTZu+0KqifekDXROYszCb/gcWt8FKCEiaaHt+Wa6NrkQWVDHDnPdu
V8ubZMc/o2qebhP8b2o8begCW/BgDGeN61X6o8njRhGTyod+63JcmAiBcTmn9FQkH+iNvEDnL+ap
BDPxUWGadx3FzmQRWdIfQSACt+NI0ArnS+y+wELG4bwidTYsQV8bLeZNLlKwUoDBRJs5QrVi9pMc
Gj+WMUdTFITtpWGT0hNZ2j1UK/ox0qnOpFWGQsAShQvlF0Xx9Plc8CfRIrQPaxkPF0HyuV9/+8wJ
XK5tElgAagkGIWp7b6DOk7GtRcyhWkLjheBMmmHwvM6wKPTiTrxxwy2wgED/Ljg3XeaX58yPVx5O
Pk0dWakcwl2uqb1J4xLD8YXIyhvF/QCVhLgR834/xpF63hd2dE6s4LMIDC56ctlbr1RezB4TIxJr
bzMcAGHOmHN7Q1fpLQzZnXiKc0fwj33aKvxw/6pkckuFYfSVWD0fSoOIzfNDwZue14psWhKMttI2
yGNskIvHyF7HwLh3ANFodSqZa4VfhXOGmPKXCzrr8wvqD3kz+5VsZYMBt3Pw1oODKozDpRaBDbft
cD6II0dMvf/Vfm5kP/R6DcKV3VxI6Tfh5sPJInNrWbq++sh9NzWb+VEQkYQxwHEWPry+eFoa4Xug
MkBwlRrsRDs7eaFOD5WoSZaln+VGC8VmuUjGi9jM4LjCx2jldizlN8RHBBScK91dZNYdWRMQpzBm
j+acB9BYDrDOtnOT4zoWVbMO+ZS33RdIMQNMMvV7ZyoSTtF9yxVmbm9A0kVOj9qbgFz1bSN2GNOR
/5EIZpHJz4GjCpiorbRjAoxAwHAAhWG3jbKeX6W+VaM+UhDj92SCaIvJ2HxYyQJTRhzC6CV3llG/
9+NKF2ydud/uqBTFrRMXOu1IAB53Jx5h3/NuWqq5xxb3tM+nFwPG9co6VQA6L5eQd/ijdYn+Pf1O
NWWZ87pUS9SrbR9DwHNJYksDbnGHn716RrT/itkGlpM0jNgSxzT4XWg5SpSYTOP7x0e0ok/vLxcI
rzeM01GXAtxxoPY0d9CMI18ccvF3D1YPvHYg/Zb2vvJ8vBb8eJ1f4mMVrZtV9zvsTNL7Y+R1F0D2
dSCSpjUKqrQ2xjnwxXAfE7qkOc7fGZ92b7irVvGqY6nsxSPrv6+6+0GdGkdKJ/155uJBrtBWV8mw
Z63drqH7/oN+pH5mVImPpn9c6/8u098E2pEejXLaaJhrqWgVgEXjsUB0kPz9BVFp/vrW0SNjUlMs
i65gNfbS1+bsnY/3DtN/pk7DrmViDNAoc8S9ipudpnVVFj6JgFRotQxpKReQrM+d7InmwqETpoN1
0md/acugaUHwjfidM8AQDpLOnus5dSaHoHi4qrwv3mFHlmHrBkoMmVdTcYwYSdfuW5YTsZUaerMd
pjD644mlsfrMk5mF6SzM/cF7HgavbPGApjRTNPWxdIARMIa5qzn2kHESeCOAPZl4buM8hXyqnMiK
qaON5/773f+utN9iiwbtPLLfmAp0+siUQcjBQwHijxgza70quKcdjqCuAgxg85C2OunbByo+WGs/
JPe/HOtKbk9UDIExUsS4vUdK4gGCZfphbwuLNRqWIFZb+Ruh8TO7gWvDO/wgJiKCszHBvPsInkAv
S/J7YAI4D0gpXYLS4eYpLW0u98GCLseAAwWptnN1Nm0mMozIAeCiEzuG/WBDtbw/kWX+1psrLEzk
t8L+OhwmI+uOB77DF3EbgBG/dA0jIlZ0cn1Z2Zn8Mx54Jc70uAL2OhLwYkgpdaYIRdEi8HtCyo/7
wGi87C5ZCJmCwM/LypwUr7idYLoWb9Rr2eqIGKw+du04qMD98kKpxObPIKCr8xkfwaxao5HyYyT/
IZYi4BGHSF6MihvZE0svx7NbUCQLrJbJMJsXJ0b8jCr+zRSpiCwY191b6t2OkiY0utUZBqZchqAT
UsBiAtd9jdd8FF02XX79K01NsT10cvnUDI4euuRjD6T/wPOYuGfBYF8ch8e5jcZPzDtKTuFPjnGN
QwPW+b+q5ruLtkyxCFFDhPkK4nlvdxza6oe0TwMSIAX+za9HJiGfMLsStiJokhxhlHPbeU791pzD
Sxm2aZHSy2FyKBkaNBVGilehdaMgROV+T8h3hpU90TaDZi3vDxHYvhHDT3D/2K6xEinfOwPSPocN
kOH77E10jdAq932zG16XJaf9Aem4eSQgmUz+vTeBb8bdHrQ3c27i/+tS+qe1WbjDttCxt5uwhtGz
MlFVDL0r5mt5Kf1niVt5OKLoBHniV+UV7REuQh1C1m0+C7m9O72kasNGX2nzL9gwiyoZGBDCjWIP
2zmZi+gegLQ6r2Lh3RDKIH/HwNhv56t8kOLOqCeswxfczT0D5InwLY5GRr/2bScABSnb2eHqeUd+
dKakJqESvLEUqqizBulvGJX7mtV+Vr7VP1fuc6KuBuw41zfKfgfPHq7saqCLNMwLOLwXR7OrKCor
0+yJGrbkAogWp3QYTxoykWk0nuR54wceKNosZpUT2tnPMlrNOJ71fXFA9YxUmA8dmSeoh6T5+48V
GNLP+cwgWSqu+D1lL4wNh5j2ewKl3CAS0C49DVuCEoo0NV3Oqt24gebcCp0Zj/9xgugHYZJeSpZg
jBZ3cuMVEM3fdAti5IcOStPGRCFOTkMvjqyKREfghMGD0KhUPPaxwYQB9IY7eYr6ZNNCRAGaqtv2
7Zm5Y1PeZ6+XOxye88ZJwmCk4Zp2lkNsla1DKFTm0sH3QVEnZHV/2fxqipIdUxgqWFF1mBd2vMff
kpzl7fEG3mb22CazYsV7xwFFDjuAvl37CMvxKCuho7f1znaXhh71ytQfmeBlLFRBpFwKDnBei3bM
i3lTf2lGmPNhzq892/eghsWYGyiADghvtJ0ch6XTEGedRCAm5lUOm7DhlrTSIxIPAfInx8zPGe9o
dp5QmqbKNu+H0M9QcitJJVWSN7i8y9v4C5HzLlzW7QNfVJoXCvc5S/3LDi0zfvSFOOi3tdngEr3U
LgC72YZqL3NwrTxLiMe/1ZpeASIhNIrT0SpP2PiqcjiQ0WSvca2mlUP8J2xGewCBO9uy67rUQGWp
Q/qvcP0uuSRRCTXAHKnw9RxVGzRP2xKRYQE6lPD9bodHYEnug3rhWZZaORRAX8+Sb7Y7vq45xaR/
MwnbKSy677/EGLYrhH2214Lgpl1n0xbtu7FVe5X0O+AcyLXJxq99ePOfzyjBkXaIdsOuzfnQUP2A
BBy1QXqIgJkB5PA+BLSeECzmAZHhZhBmNVysturkmpmK4yZqbpgCaabpJj89C9gfbwNTQzLk7xSj
QpngWtjF2768bA6nq5xS97DzL7VIAaPgOsGUs8I55YaDzEM4rs7SQYii6lpxdAKNHvZC9TXrw/cL
wABkh4QId0GSwlrPXctMewTbYFZThhXAgcIk0h0WKkP2mlgtTp/n1AuRV4qvi7e3bt/ovo4lauVS
BFxo4s1OYhw3aMcEQMZKU6O+8yo+LnQoumJ07u+c0uBY4Ycom5q/KDMWLpqqE5rzkMZcX8occaI+
dRNjA+4xrd7wXMpo94oSGAvEeJarS9jI4w0ol6tLTazZDpzE2fCvHy59CVGbZPwDlQlFgJ3maIKe
nCKGNC4cgfF+EvmLW6U5vWHqh1tFI3E6IuUA2NVQoTtHlxszI3QSEK4K4XFLHhr08WJEVcr7/HR4
iAlaNab/2q1dOhEQrK7A7W7a338CsRLP9jPk5rzTPFHpHDDXzuWShnBPQkxurosQz+wq3K1HYEu3
hloh0eCB4+zGx2sALxivORzCV+Ol9VUR4JNesuMLTz0tzr0kg7XKD8TL1oojkC75mqfHNc1m18sl
DMS1CDqhDlxkGKe2/MOA0xXvThFuZsn4CHiSqkVHHEeUSDgTypSOuUnPiKu+wHpybKZv6wt49Htu
xBt08tTX+u6q60f/JcV4Y5/oa6cuGfhDKmSaWz4IiZe30Gp1DepeTpO83wMPAtZ7sEqVo5jwQXOh
Tu83LudZfVlumsYVvXmhfbjAK84gJVQQlQvx3XXoi+4ZBQbiU54j/qa+974aOR/pn78eD9DWZlQE
m5+qGi0qlHvobxx7nbmyChuq7zlGRafb8MpjazlFkU4EmbLbXQ2RZ3SjvI1eQfImuODT4P6EtTGG
zDN7vaPe5/nr9Skx1egFoWvH3NphsHtZa56lc0lj7bGKzaLGjnJpE+DYjb/Tg+G8q083X7wtC1Bo
rjanD0AyoArTW5FcfHMCWNW72iVrFpgoHknK4jqc93xe2MD8+aZDMMG0U29Zw1Kh7GUOH8EGWb6e
XILFhJq/lmqqvN8AtkZ4+euafZV8r38gvFEV/9cuufbPbnM3MUqUQIgjSbXX9mjyIvK9CON/284F
qzO5JHAqLCM+lX19u9XUn84ZkvoJEMfH6O/i4Lmi/RC3HUjI2yGTOE5nKyVkAxbISM6aYZY9Ow0c
eko3cNf4/3HKoU791nkj4X3CcoaI6bvt8Q9uUbYMv5E3NKzO8J7K4tHoEZIqpQmd3xj1GgFcDWwp
lt+kk1GZEdNz6miuJA3Q/uYNtE0gageYHjlRarlA0U3pkS89Hel607T13HVWmaldKfWys9WDx3Hm
Yv/7TgXT/2jT9OW0prnd1NZQcveAF6YCvGYWkumt9ocTTdNhhzlv+y7uHb3//nsATWOCM3ONjPoR
zw2btsUmAOCjqigR8fw8AEttgpK2+FYfK9+KwM/xUtj0se+CfgKOyVNRKNrkydzRGMOPU84G3/o3
O6ybNwgQNLeAMBHLViS0nDo3x5+8Xlj2b47VSEl5WcZnTHA1t9HRKqF8AqQP60mEIWaP01sbvqLw
HjuuU7QHQW7CCbrlYuMs+lmO1eyAmy7JR1KPNKZjrqR+YDMxpdfDt2ZjjUMaXs9YWe0P1pexUZRt
HZXupMLy0AUzcUoHMyg/cHLeVjg2KscVuXYVnZrSUaIXjEJ4yawnSp12mySSqPkyzA9534YoFU9M
vMUNj+VK9iJjaSwCuuWQfFkiKvlqC2vPq3ybwt6YN451W/5S/rF7d+VTpF6yhbiHfpWN37S7doMw
WsJXVNu5eH30H5TkFwh6siBOyZ/InFbFi5/RU6rcueWGm6/lia8D57faUkNdon6ezitM2oRFV5Ui
WhE+jTdwtyrb+k4nxRiGGCamjYG0IyJ3a3nU0YIH6a+y0LePWOy1qS9WlnKEn/ReFN5BEQSdATZh
XVkMHZoH4p3BilUMUuxQEKNWuwhNTZ1jKTzeonMKTgfyjINmOXK+XWZpo64IyDwTT6o0QU1QHj9q
X0rXQxw5Kc5cVfuybBz+cSdKEbdTAyrFltzu9CyKBj9zzlQuXdvWMqCuMAZzChvCMpoT0kGjTnQf
zG91tP653/ayYIryFsnzPw2YhYj+ogw+4+BH+2luj59YGPFGwTuvG6Xpe0pccQ8fdGSk1cDhe/UX
CZK2JZgqq7Ad3ZX2lJBm+hFktDQtr+cmsouZ1KiWMlUC8e727RtNf7xK8JX1V8cdI/x13zf7Wo6E
A+sWHr5VRTut5IpkcV+kd1hGGfA9u+iPVyGvtE9JKZ5fPSqiH0ix3jjMymvWV4zqYDnu2ZnnMh1D
O8+6uN5AZ34wzMXgC1ctbhUmpm2GGNCHmwzdpXwMjHAc6Yx3OZ0HuKbpCUF1xi52lYIPjwgoo8hw
OgJfpUF5pwuKklqtuRWo1996FmVG3BrwdzxBUoMOksC81vG21Yh/6L45iMwFFIPjxhLvnpt8KcoA
EwQKLIZhCmgPzAnZswr998lLCIyMM9LgrwAGFK3OylQiM7nOaDEd6sR9H+0Imw2lv9eB6mJQh75Y
orgr6FbHgM/KLXrUYhEZ6thiEqVkibBoubdpWKKDAKzVUWhyp0Z22/d3wAkkCQAYZsVzgrEyULpy
wWoBGlFtQAbySHjXyaLqD5k9z6S5gQVkVNfI+ryQrMO8hcrg9NnR+O9COzy/ZsydE5fmc7+WNXt+
oKWmBMXaf0l0AEpt8fiq4Lsyg2ZQ5t5sdDPfgrJvZEbUfpOjn8RBYbvUYVioaajjGOSAA3iSbpPL
YphjEi7lc5m5cWfUY37GzI1uHfIbbmXANl8faQo2WKFS2GvCnnSJ+8PCXYt5Dss6RpxfO42peL8I
GrTjwCDwqr80Jcv1TDhQNy3ZJuH2/KP6jbzdTPT5Aj19e9gwKyfLJ61lDGmuIBCE8S9OHwsJ6yt+
+WBWnlCtbHWDFnjvGhj5fAzdhUlSO/HDmSgsZWC4vHTcIK5iRzIFDXzAZFvIcYKRbRge4fm1iE+f
PlcvKPRKmrazOnBkbMY7g5ReZZMG8iB91ET12uf8StlYI5/GQAlt30f7iVgdOwpjEoAOcI4YwAVg
rKB0xfdo1MIOUWuxapmgcmmiwNmE52fBU4vFbrPmAbZ54L8NX8JbcgTbanEqEK+2CkL1q5bC+ql/
0b4UY1R/SotPaRWtgUvcO57gW7f00DKaInd8Mlydf206azKE8SX6K73R24Xky8F04eZciwM7hZvW
kxTa5duWQDPfYD6FmA1Hk9EfPIhLXp2lbtKXykpAp0y0r44Kfg93PObvhONvJiTAUbrMhGe6je9l
erSMdfzq7kbSeu7KLLXWxhN9esyyHqFPs4K1zgHVxpsX/IHFunNTphRiPxnQoN1Magt6Ce+ioCcU
+zd+WNBEBVaPHPRs+zFcaP9qW/lhw4cIoIRiqKriTuqqvHkVsE4D59rnpwoekekfZlFG7O5YAsf4
e/YHck0OQlfWOLoV9yq0g6f9ta1JkHE6DfrKoOEMlDtMGDS+v0k9LKhkHN02+EQAwS7Rp9Eb7eGw
WMC7WtCIRCEZm+aUZpYegVXP48EMsmF9syjuExp9u9+GR980N9qrgbdzWI/r80gHLYrNq87GrWq9
N1dDJME2ESQSTxtTOfRjCme7OplXqYcEltxjHGXF+kDOwRd2bTmg/oi0xhfpu4B1NkpxQE/FuRrS
z4gv0azuJLeb1qMyw1clFbyNer2XCAmr50nOs+C2lnnneGfQloep4Vlv9emy+/yrP33LxPfILuyz
BrzD1n6Ctl9CaalosoyojndphL/3xQcVDNytxMACDS+y+Uhh1Zq7t8HaPZXjoju2cvJ+SUoLYTEO
5L7UXMxBjD18r3GDvpVMQd4JOruAat7JpCoigYJEpSgZqmHPIRMHCrsSVUPRZF9dlTKNgsv7WcYU
IHsxdH5OQRa20zqAqWX3PC0lGHZUV9UmlQQmtmeS9XQZvw1PwgsxGTMt19zrM3fYiov4AGDi2rkO
zX/RNnw+R3+ndohX3Lf/9MsJ9JsxpuvwyP+QFfom3Ns5mqPMUHXCCSvRVU1bDEfaRIQnl/4AztBf
zk10JEfgQONh6jF2wH3VwHCekQ/KN6BjMMOZfzqW7Jz0rnCVzu9GMcuRyvKA7WJfmkzQF1Ked6lb
K8s6W34+nSh9foK29uOjA1a2EYBbtdmfY20a6lZQjfkhiHNxrq8+4NGiuUgyFsFG4GmZZ3rfRUsp
DaPRIA81K0XULWpgyki9j7mTf8mfnVc9PABD+7VFgvLqgcRcosPJ89mBJqYnOK901Y3QAjg3MA5r
ZwrVzIea0KJVKZUXRlYCQi5xcGfKEy2YYPtBhEH1jyCEk8zUaA/Us9K0dINiRKt7jxCJhvt3GLD3
LDon3rJuXHQwIkXJr12/iSAIJHwou3ukmlnrL+U/l7ynxDvSQAgl1sYlZoYyBkIKvJkpRkgsOhGQ
L09SDfQiDAbwhR0a42N+my37e3gnzsPGu1hRho4AWdLPAdrmJ+SHCdN2fCjuduTqSJLvJVbjli5K
OICIn9tXm5OpSiA1l/+af3H90VDAs7Do8nKTiQ41nJwo36rZOux538quIWvbk0+InlVZlBmTWQpf
AOWFsnqukaTCqFQuJQ0UGbKxX1OGgaT2lju0asH3pUd4ArRFrNg6/gCJLz2BQMj7TPQvuqi+o9Cj
hq1tK+bXGOv9zNZaWAxac524duHVjnsvFiiX1BMavaPY2ppJoERY8SIsqb/7TeXr9Wz28K5ogiZR
XC4POdKM8YdWftYMS/Ymqw82qVJvPyjCfT1CFGXeKg6FLjZfszCtvGzeU7KE5dGrNwT6OiuouM8L
0zagfKcsimU38TMlahX9Qkl0ly1dMlQbMVpDiDaTdz+waKvnu+Eu7n5KgBbXUKtKJ5K+7hOdy+ac
XN4tx4wzmeGrI3wRRmiGdGeZV9ffH8f/RBg6dHP/otoRtAVM1DpdChMcczTYAHIYfnHhwAoGuc3F
cGsaZmq+g9JBCsqCyxG0nPEyYste2Tj81ktwVwA2yOS6bKthgTX29NkmAVzVggIqF6qZ8bdSjOqG
dydx+jec7shNNwBMzFGSKoUg4Uw7bNzgHGrbp4y1FiZC6cmgU+hXTsteFwUB0szDIRLq7NTV/8wj
gO/OyLYe3UcZJf7zvY8ARw7AM2RadrUp34cWkxBuTmAC2YQXWYqWPVCTPij9b9j9HHzBbTezztUG
4muV1zpHq607vcjbVkM8gGr3FFbCGIUbugGqLAV3VEpLIxlLFLhliKTpHncldEsN+6SawxE4I1+j
4gfMyUDF+AnVVIWIf5OpiCtV2D10LI6SMThvJAGhKsvsrIwMiA0L5WLE969/C8VUI5WE+D0Eht30
/JN+8Zn56e2uQXV4qo7D+bBNXNT8puTq1PL6fc/2yCeEZBsjqXt4bF/wddrGNQFnfNQRiGupDZbL
gGiYz1PpQjt0Wfyg5iFHsFfJe1O5PrExu85Ean3Hg5inHr9yV2bg7YbiRTKGuXrlVfA3YBLAmgfQ
nsHS0ZhN4Fv1h+yNe1QQDyvXIHMHOryanurdd7gD5JwgJud9QZom6+m6Jtzswj4IYwuf8M9AIYLs
4HvXJkjiUuG8nIbJPdsKFOvnBw1WNCzII16BjHevT2db0Qn0nb+mLOWfQsCZlX7RiQXS+PmCqw61
dVCxsJWWmSj5EKrHzJUtel8MvCnpHNFd8V49hTShFf/QbWVAHsUsUmk+FGzj7ZY+LTQLxUbemi6X
64/mmrHxv+m/PriQ4R+xVcDIaT1DkyBIPNOK3SrUmCpBziKZBbEBleCKKDEUEaFhx0jd984SI92y
hGSmbviWq+VxTFTggqR5BB/9xu+aV779A4QLfg022shPFTeoAA/omjffMK2Y1sG3lLKWQ93QWf0L
Hx9Z9r3T6AeHp1ckH80zJ23909hgN72Fdh8r8GSYYZkRURF1Q8/wkxwgyp8Sm6wRZT9sLGkowT5Z
vQ2z+AwFyyFJopoFTuCaaNPAFc0IZO8q/n2RTCBimNA1q7ZdAYTymGnb0lne/KxzDtuVUji9fYpg
QixeVTpXTeRGNVg3llAIt7I4uTjsSg5E1YImrhrDaycfGBKealVIyRvFdsc1fJ5TYcnKd/8Uzq8S
FbTguGv9sVAKB8t5s37M9WAhLRI8vMQGO1VM8QxA9Dt84iEwuXOfhejySFIXyolwHbR1CY0qFESP
jlvpJBl9qe+TPsqt9Njp+gDJ1tKlynzXbPeWt0KwtrtlSaKhwIlHGfLgGgJ55ixLRUNfaUo3oFpC
t5N6ZRbMCIdj9rzYa3exT5uzu/O+s3YxyNPp7TfRZD3b+vOzpNFU/MM8uKD+e8Rcz7xfv5htjC/7
gvHQSIuAGUXfRUppae+9TvmZDKV4vfGW6thLaFodxB8EbQ4mn08WwGikuT1zOtip+Urzn9KKbFFn
PVwZaMqDSGfwYKQoInhyBF57a/1+bFF77p4nqscOOA9vvSUdi89Nju1jKIzo4+2u6lkz27C6ljff
HlsJyB/SC8lBZK0fZ4mlAymw+WWZhQprdODamVKA4M0mFh12t6xDYAA7IsdhD1XMcpDV91GMS1Sy
W+t169T1ukDvPVEKo+USJk+De4Fv2zEqRmSivn2o9KKI9xYzlqDia6LqbmmbkUUbJjjXnSvMQ99O
QQnwTltOQZ1HsJF75bg+WsJLNq9G3b9vJtvdyKdT17+61OqVjJ42UQatVT8i1P2MFdousVqHakq6
CUUSCSSNHXfJXa3qIGrWOcsOY8/GxFpsgoIOXKRapoyQ2dTjWBO0dX4PMguOs4aPVR0henlqo96d
lgkJZ5k7csGgByptML08ci2dkvH7OgUBdQpc3uD56on+zAZLXnVLqOuZc85YpThsQZVtNjP1UyFl
lLAQwatfVLKqJZuMepQb5xulLtiMhyLkzx6JIBwLkPL60qO1PFdx9KhXNF5cQM7N3RiDHzHSmHXn
y+4wjxYqnIlQFMkKhCvf5LseeawVyFPln3iFUrFnUvp1fUazlvdw3CtmvXbCtrw2qVZzO+Ner8ru
cWX0eNuihLWavBFRK1hreTykY+ns5/Nf3kxx3lsXwHNJOPRbk9eG4sQX9aWjR/X6DvstXpu10X1T
SMweV/LiZwpQEr5v5IpKhL1G6zIfUB4YygdBeNdBWSI+LdNtyz74w+CG47pFh6/9Yd4oENEMk3gw
eW9OBOiiNuUE4bmP9vJ9UvWgisZwJKcUpZIGswBkdNgec2OrYlDoi/oAfQblZpRy2fKf9SXmfd8e
ZoWjdV1D9N9pxUY9T+o85MH6mOoYG/O09p9+8mkMVkiOdhBi5eVW0d4mfmnQlq028hau/hGNH133
zCmX7Yvo5u5ckITrj/MxN9/S/VHwSx7ZzoSpF1WYh6AL40flY+yqJ7fvCxJDjLUPcLhYJhVosQuF
jhkwJWwE07m5xcFudLrX9tR7Omggqaeus/5JrkvTgXWxMZA57t2FhYc/ZfWbZ87kR1CCy/PRkZDP
Q0MbSGI5/GXTX8wNVU8KBKGn3GKCPMkE5xNWDqjAAsJmxq4qO7Q7sAkjgkRY4T9jWRdOQ3ydwnff
jlZ5kGn4zTy8ugpPiEhnsIGtBKrEViQ4DigU1KfzC2VS0hiUNiY2pPRyOFtw9ZsoAVLY4UuOozUl
vR0pFb7f9uFMeMub1MCGllrl5JU43txP0OVuebWJtrIcFmvKHL+uth0+yJcp//W1DwuVrm5y/6R0
XoznVqmShU8UFx4wAG0IS5KFBrF3xRI9QXb9iV0SxnYMJ9zdJaOgAhflSzn3jNrEVhrBJ2c3LGht
ZAxyFQPpXw5i2QNG9jd9MnV3T5myNDQFiLabkg86Q8nDVrZpXSWXQZvNseib66OJe8YCP2sK9apK
wIRxZm8RjtV4FXlR6qN3h3IHdqKDPeKHA8VyGMdm9t4gDXd4NVx/8t1GfRWzrZErFyla5eUYdF7y
AGaKnLdzEOzVTY3xC1jVzsbr/9rJ1S0jS/bPMPaZrdiKg+NN85VrXTEUY5S5gfrL9ieaHS9Zykx0
JF0C1Rku1nixdAd1XJTDcEOukEew2HZNAycZ2Vqi/8W/vIwAJjRY0x6SxKmb4wexHu9Z7qjutCYG
BsISFgen5LrNM9n1d/0xbKMTFLfXGIBWjS+E1STbXMy57fYygR8RNhtpUbHyy7MM4uMxILJLWOzB
LA9eqHUw8r4z41Y+4KMz11JosYvttzbv4OXiNSuupCCM0FuC/C+wZbDvBL/e0EMtQM0plZiTD/1E
XwZyedWtzCPEN2kUrf5WLL8zHQKzxM9EV67a4QTsY/2RPQIuzwLbhUM7EoYzj8hC80Cwfp5LWXdd
4k1lOQVoxGEAALhy2UDcA7L/A98Lq/h+vSk+UQgqgcpoBdjAYLWsTNDHI97vnhco15KBb4LNvsG9
sLuXo2E1gQfVdHdykHSyOCp9m8cfekWJlSo4btFzT5Su6wbeHBuS+t24Gfe/EAnRSbAyob1NZwua
C2g2Y9OrYGjtibbEGK+PO5CDWqehWF/Pk1hKH/8JG6hBEGZUrMIfZKimS28KhJSsRU2xMj4PCjWT
sBHgDJR42dkQLRB4sccgp802wXyAyyfeIPwdu7b/w8SgWnFiro3zeWaQbGE8D1KqHUWQUP07FpQV
1n8XwkYlmVbELIL6UJPm07wVUcUCPw0TI9q/qytem3Gk2gR4Fyndsf9cUoDUE+oXcItsqOD+f9zm
48S8KhiGyLLuFACJuFeBNIy7t2cTo4mLg0WgGykkIVB/85A30RF7cmOn4T+EE8U0tXGYKChjWw6e
STLj6dnloQO7SpdzWPG1NIkCCQqDwKUKcBMFdqxDJu5KBO1rN2xfXOyPow/BvVtrb5HoaJscn7c2
CzGTB2F8Cau+eT+oe7dVJXYRsr6XjWygO/mMXur8G9lEqqIcmdTqmuXKvixdzWqgpkWyoA7hhlOd
5oT7o+oWyPYFHNoghnYtU3JcPXvdoB2FC3oEi/gegbmAeTndAfavNEmk7G+S7Qgd/to4r+8TmvST
m3Z313EXkW7u8haGppk2hdsmbg4h2qOfYPzfZi88JFtjDPCCn7otXG0NyJ//3bti3NMaiOWXrf23
lIQbknuQGFA1Vp/ezHax1hnAuvTyKHYqRklo3dEJqsiAdH/GY8Y8Ti2qFop3FO6C9MQ1iqC73jlJ
mf2b1d1470Jiww+pOljuvbSVJUwo6BuruswCRCHt6uUGTZ0WpqsDVzbSJyq0NLNm9gxHCvQzIXmo
g52apfl9B0hfHF092tKWm0R119mxuIP1/2JXJpWT8ZwQhlWGkiFb5mmomd6N1JbCncJ5ddZLWwlc
MtbkFqNp3OTspHoWtz8r1hYzmoVqUBckbkOhCzI5DI64OO5wH4vB5AnVlR+EL3WbIEApKKGfTiyZ
vsVzRGFV2N8r1KOTW/tOSa0dEGvsQ7w5dUCocSLHWCyepeF1Fx25WdziwsqO0hRF4iI42L1S8kL5
es/LwJGcUydrftj6ItbfFNdQBcD76nqo4UD8h0bkWs3SIPuBtqMz/3kEIyzyK8AY2zIQURzrgezC
PjN5Cpgfcr9JV+dLobzhwx0tB1qUU+2bhxuxVmZ3MNOve50q5WBEGon1jGDlIGYTFINibMPy9ZK4
+8SfujdUIhWD+/Zy/tbdwpD9cNC9ckP+rLEmyvMu1oTgqtXGg0+MFrp3vKKNJ7oxYFMDJwNOJTSy
KTKI7SO3mrPGUr+xHH/gFkbYNTCQ8VWxlFadxhqeWxgwUPh2m6kwYhIxU5af6VHTttkU7uDJnIWV
BYy1Wor/gOwivDOP/Eu6YMAeI057+zcpP4tELMUt2RYdniN9+783P6uckktOFgrD5S9yd+WLnGeG
YDv/z2WLYJZCI6emtxVSp8le3o2Oq8WlFO50abfZ/1CkU0zRsCFhtDrwjILt2H57iBSEygY4OTL5
AQXwjiP6NwEwDKrqsqz616aId/rfYOIms1GgHw3uUj/TWRMLk4msicPGIy5DQF1FXZM5dtuBBTGX
PeftaiD2yk++gNLnYNEHhFauhdCLNnaFsQp8BLezYlMZT3+qAPfQMqqhqFKmux1NtPKz5y6J5N4Z
NRySo4RtBqRZcBVVyRo95/mq9LbtHhmiPGRj4Eh/EGRcvIqfYSzzDlTYIDo1k+YuvE2yFbYKZ8Sy
bkm2PGCMo8IkOu4E1JJp+ZOzRzeQXTDHA1uVP/u5MQdLs+pfyNFjCFTp/1LudTkYzkz20QBZ9lM+
Lv05092g+ZBXtwkTXwCMF/x7EAP5R6/decoAcC++Y78iZE7dVgkj6yw7GqPzpZM0TQjaQZwXBUXe
Revp5OHAveGdYTv8wykQDPyQW3H8XqKRqF0E55FJ1mhDwhxPhCjcP47lCi3xISD6x4qpf4vHcUWV
6QmQfFoL7QL8bpmqcdS4BYJWNEfnB5FVrBILa0we6+WTfuU07idXYcaHVRRkf5GVbie58VTM54Bv
v8OD8xU6AqwWFWFtnsya7LaH8msHmj+9JCVdq2j0VE+Hf6vZWLck1T8OaB1gcVyc9hqmP0Shsbzg
PEosdO8Mlm2DgN2s0kpxlIp3OndtzhWn8zMT1+VzOBvHCB6/5E2JPyClu7m/u5IEGSF16oolm0Qp
Q2b8m4fU5aXel6DjIVSXloL1JM6ogQ8/i9XNaqOgpphwbNlP91f0m+75/znwUcdHUYleHgpj13nT
mInk90Hnw4S3ptOkrtm5UVwS2b4BPARuelTBO9zmalgIxXf2ncYbJ6dO9iZ1gspPi7uaxsjPXxaY
eXLJwaxLa5fXR3GsahY9bpKqHMixoYGcLgq6lxMc9DOOsgG54o/+nt6mhmsBHzpGfZ6GvXJ+15pv
kVcwInMqhgLCJFYVWuMkyvqxv/qrnAIZpIO32CzhRvf+C6LORcOexq5GAiH+fLiQH3sLTPuOU/6z
uxFX6/YcxPPeYPPA51ldedJgTxi59fZ3NYGYaxmaP4kt09WMOjx+o07sDqLrxGR3mNVjs59WRhh1
wb8EpV9zfyq5UuQjeHs28sI6kZbFt0EfbgiRUmUkg1qLQ/9uSJZhJFQaueYE6wAGfVLx1vULWF0N
rxy5O44ilxFmBxFQsP70w/Q2so2cmVtRljpBxXvq4yIJYdNqreIkh/nUEWh6ebZGgi8eJ8Z0n+y8
LGNDDkkOWQ4xgQWtcf6jgQPZspT/zxg9UE31/dkRLtJTJ97jU6KhfcOp9+uwUnUbKJli57xOthAJ
KdZtJRz/fGKa96FVhmwJxmSKnyIdPM9f3zWpydIFw36+N5b3rtGxSHQvFVJnRn2QvHKc+qMz7X3A
wyJgZ9Wg5s8BTggXh778RBBN90vi+SD0Z83NiQVhvt0RDO8FM/lRjznFzxEi6JsGtp9CDL+rbBZ2
C/R6NfYifyJHLI2MfRQUBewjXlA01qWRtzOGWtsXBdFc0ZoeuSwnmLry16gQ8h3vnSa7O2ETE9Fh
m9HkK1J1ia4vkvoQup+AcGa5ghWkSkSoBSLx6Chz+fM6BRS/os8X1OPbEIGiCKqZOxstLjwL8p4z
MktJIy9Ie8Mk8JTmHxACcUtTTrtQpjA7x7f4QspOWheVB3AUOANOC5p1182pqiFDHSofZwBIlMIW
55jfZNumBsW3/Hsj+kydLLYzQWCDmIwD0j+3dGbR9Bo2BpuE3/JMWaJ4Ry3McXDVE3JE05ZD9KtM
lOF5PVEUNdTOrbp1QbebIvVfj5kTcrGqq+rgRNcu9ipWII1hnzyxTKQvlpitVTg3Q6UOhQ4xPtry
VBOcfBd9vf2Br3fEtOdQrLjO1vW8/+VQYwXPZ84rOLnB7aAoDOeSkFCTgLrj/n9h7v0gbM54HsSH
Shca8avXKEiAbhmvPiTJOsMHb6sNbjaRKx9um1BWY/fW9PQAS57qHrr21dAMJhZru1kWQRZjTYpg
3c7slHPTKCZFWPUBNk/1ekZdR1ikw9k+ysakuqYAL/DMRMXrR9c4lqEzu4JVdBqA5u/sd2G/LZ9W
wRUlRYY3aknBXEIlODLtzJZwsqmKmARFBwnB08eL0xgcc9dvZOeyfl67CBD0Rz91+icEZkD4eM21
IdquOsoj97w0RvRKQXOYlOR//7sIXsB3SNaEOnTtdsmUnuuo16znuCk+grsxRDTz0mL9QEtI0ZMf
HV1oWdUXTpWFBn9JGdmNXlzmbC1t0VNfx5xn/aSxAdLNkWijZizjXa/r5gP2WCfqSXc9NfOVkGQ/
BVpgQvRqlhhoout9JX+ulTUDAslJWTAoFhSdds4nxjOT+202obYZQYUKfM5CL9Ht5ygIOTHYYsrY
rgvYd2crvht0R7+OZICgCFpxpulfCketiHeHY7EfKdSgyUTb9f3TdqR+oyCHqLBioUHoErZdzGwL
ux8/eVqGm+VGr4lIVxXQ3UD9+Kl0panHcNDRCguz9WoB3kpEw0KqybM9ap7P+MRk9/OweeWm+0NU
b/m2bVaA5N5i696sOvwRLUJZAl4Tluf4qJdk8IfTVWHQ4QxsagPjq7iKEtFfKu7IRXus+tfUQt7q
t/+fJ7C7Qj1ilEfyssW/GUNGYJPzWFcjn5gzmPkGhVrxHcKP4DncWeJi0P0U1mqHVVA7axZFRsw+
WYXIqLwZ74t2MZqN3P8FPKD1ksXhE2exGYnLRzNA8Byll5z7lMxK6YQPOIC8uRCqa+9ZYWxR/1+7
R72BDW7qZn5it07q8uuY54u+9FycyAGyKWyT4aJ3iSKsGT2BT5my30beboB3cL0zSsKSYUB8XNo9
XWGT6qHH+mThZKDwS7AyV7t6ji7nBUZlyjmx+VfTXRdikf5dFAzvJcDLE9b5KtwZHkpSgHVos6Kg
HsvSofv1Aum+wQzOk/2cxgmxF70QFBijr6s0Qpf0iyUmuqpswPUboIbqJ+AjvQnvIDSplR0QXdR4
pUAg0clbA1SFWLEGpx6q7B4yESmjAxpzf3HZ+XbqfrVEdcOlw4tdkV+WJeu4kXP5L4p/Cl4FKWDN
iKglkwKMi67DB91VJ7/SCZg4aGHrG2Ah/nQz1lm2n68WHoeqKRjF+hpOiFEy4g/eHO/1LJtjKt24
tJbjuChVhlA55XTV0zSgLRfCzYdmIvIXHSdHfTwNkegSNrDGIkDuzV/FxA5dKwFOO+tHiPvZyXnh
PODmQWM/YZmQtyO+64+MHhiyJFRNMtPvEISnQBhDXlzlYQIAkK9ejHs4++QzFdpCHY8tDLP5ONNM
cnclq/seIIwj6VeDlxZdyCQaU5Obiju3vtEW7KjgOovnJME/YIEdzMPtMLKhzESbGP9sAfco82K5
yPPikkfjg0J8Oza3pL9JgHPxVN2vmbzhCN37XyghB8C3sY3eOYhvI5UboiUjGN4XmRQM+bbLQa6Y
KTieAVJygPny1IkekINVid/WlbhuUaJYVjAiqhfQDU1I7+7eSCToIK2+pWu03TNIxSgofEeYabnx
3zeGjmqYbMXKS5tgFmyuTXzkH7ECmgMxQSdo0EWemsKKgRsFp9jDm5zuvxiYgXU0QgqJAqG4Hdil
+HRQMhVVA6fCNGFQ4DXSiWhb7XjZuBit4Te6K1In6Gzgmg2bllaTQ0hYbrIT4uromZRK+MHz7i2j
GDfZK1G+4owfo0u682QhBRxS8CAIUyx8Azr2zGWBqYYBa53bmZcb4bi06OZO0K0la/tR+N5GaIWL
jSPkNwhpk5xNa6lMwjhcZajocfr++mz8YPZDCXQRIzSruBMED8SqQIUhUEkRXb7FwMw9YGmONjwR
6uuz9FLeDy4dhVFPETD9d/CAizW0wGRMmT33My0Rg7G3HJED3YtKFZtDVL+Xp8D1dl7IAdfbW/eh
hrOhEQq//E4kd6LMUQshIMkvHDKVnWTaPK6klA/+1aJ4Ccfja5czim41aFaJAxyzbdT1gnCnasOm
blC657su7kYZWGTiPZX3rANxXZKhX8GsYe/2Tcgnf/pKDjc+We7gcpv0hZ5tyW95O1hDR98Yth3Z
PKYc8PIG/6EnNTVzLY64lyfoXepakUzUuQAuWGc4c0sTRH8XzIfYaXmg3ARykgj5ur1dlk3Xr45D
I/B4p3RUu9mgUinn3og63v7+TyT1bPWdJCySifByMteNWX46T1VStj2E2VYzbs+RUcknZVlvQMMt
u81xQZn93Zq5zeTHilgfQ9eJaZqzoXmaILvmNpsHZ/FcxGrha699rlm82PljBA0+gIe4mOZNZDSt
MnTcIhI7HLc6OmpLPqENEUzGmVm6HLUNUSx86x3Gl7MEwXhhsxFCaa3pLfrIlLWeQQVRN/zEsHnX
oAWuFebrgAKkmpPxxsRfNimgU4CK57HQq3w2d0fr4ErdXxnLAZITByJiidAkrFECxrZGrZZ7xJLn
XbreHqW3GSNqZzAtfQtnivnbLGZhoSKbVM6laid2q7SLUQIbs80rPk+lBjQXWjeiqlarT7R/PLHM
rbLaEcY+Tjb2UYp8ERRD6A+rUwNGQVczRbun00aK25jeSEttSmuQI9mZoI7z1XxnsnN+NKKDq2T4
lR5RvJfLadGxNVY9uhDgMhYcpXEWiClWtRPcnWlwaNIKbGHLNnF+S0qLeHnuM7IdYw/cyfC4DSoQ
1z4hrpEhT/dVxFzT/vvY53VF4mDUSLaGDY1n8PmsCArQDx5vuyD0OLA7ACGyIZ0GWrrkIa3006/H
eKN17ZRo3XyDewp6xeOCuV6eEmQSCC/4m4CswKBC7/1oBZ83FOB1R3/df1ALPfFiTImOD/CZXQYV
ofYRn212G1I27W+sYBqkLk4KOof6bMQJdkCamEAMKrhBd1TO4ieC71HTdH+aJNlY1lf6bvTTxe1T
HGf8dGf40qDwX3vcLjDEeh9qYS3NV5VBBsabZg3jdF124N4U55LBVqM6pqks5MC6DTOO93MWemlz
w6r1WzKjJabIM3H7Gk9F/krHDVFRBvPx42zAFZraENuKet40qJ2q60RZRd1mP+zioRAdyEVSPJpc
EYbNnx3TJSzlf2dVog6H7iFcYi9ISiBnaqBBojeqHtOiuOKEdHQDYwAZGXO6Tmn9hbCHKZGlojyc
+cM33FsLPuCk8qPkQVVdijAzq5gQbfyB+Chcp3M7cHZXai5mySthz3zTnNPdrhNCe9UQGpSWXxoP
FQgKl7Mk4n52QA7v+DrNbtxO4NkDU2ip6ImdDssluAHi7Wyd1Jn0OWnr4TtH7z2D29G2oWieYOOe
egEv6gcr4iSzEJ+jZ1pZmfAPbUEqjlYu/N2EYyMXDTgWWy5AXIIFc0l4hfyIWVxG+7fgsmx4Olf7
EES73ydSwQ2JA4EMMMBGCJQw/Ie5v6FVwpGrJPK7EWBmKaNlf3iV4KXsykUVkZNl8PTHRa7hei0D
8ritcOm0KmQlN9XLPLrVSZ/JVAoGArdATyW+JwhIaHPMKKU/TBl+jGX+7DmbGMImEPp2siiNSS9K
u1g3toP+rcP5EEhm48RsGTT80laIHAhi0WS1A57JLyfvVdSGDUQt9SB/WUImvsoHu3Rsdq5qo6FL
uKHIlD8v88omBZq9foTsRb+Y796yTilDeBIZoMhN5GtBoX8SWG7yidIYZwmGP8YAGx4b1xhphlOd
olZlf+ahGHX9OxSWUP1JZdnBRzD3JhlVgPFDMdMptTMZTUgnHsMcbZm5+RHI7EiDYIxt3JxAbVkB
B4a6pb850HG5QBwcvAX9kCnOf8U1IdRhDzlVx19aVkRxz/eLmubE4bSlcYFRIqBeL63GmzbZUXw3
ewKlCrUPCENmk44VcLmm8668m4aiqKtCHz6K3JkRPYPvjhPQAfzYslQaYpRci1uvGYDc4zeDH4k1
JCFUyPoW6FlS5G6M2rf3feobf11rYusT+CrtYDSD7jw/sMVRigutbfdlZ51FbYW5kgFZey2iUu8/
KHPCC/kWL8wRugc4mhZHP8VxakcaeHwgY4HrVu2afSsmfx6Kln0ZJYGGvEMRFDQwCUPpAuzfGpYC
t20FRjmFfDY4DsJ4FsvgkMiTAUD/zzzGIEtB+wMd49BrCp3QxeDs763UWRMkGELNosLHva+VxKG2
udUZKblQoLxmh3vfI+f20OAaG/VocQCep2GfVSrs0Qhmtpe+19sEMWfraKoAscuJvY2YRBwcNwN5
MmlRMYLoOQwp99zqoZMSCJPTXV8FpyB62wlX7BDu2fBeAQnIlwhMEomBa01HcCcGivO1i+d8utvA
VN5f/F7/Be3aMVBakVEqeE0dmlilk5tzqsoh66q8xPDRLX1k0ZV9FAaRhYjlf+ei+2mWrJSCgWs6
NAf7ykgGHlgaIC8Ukmyw/ou/4KaF5R+ncsH33xSPCaHYJEe4zKIShH2H5jvb/js7WQCAL/HKYZgL
665x/qnSDjJWDpF1vpEk0zVSTObCOPVhzXyzPT8kwJwT2r+dTXpSzEzZFDYNgktPXuUaub/WXRfn
TrSDjypS247suC5e0CQr9UyTJv+sK7IXKEqwM5EulSH1aMA2Z1d4EMTJAak9tZXHRBXfPxY9MgNQ
KaHcEu5Tvw2uTPKtGaGlU+MOclqSjZZZOFGlDSMJetmEyPTuTa2HIV3CQOUR7LMREJPnbEn5UHui
HbqxDLhy3tXap6CTOtFBM/e7BFh1r5bcLsHgi4FHwlj9X0cdBsl2lzp2uVlqX/6UM3caeNPbZzem
RE/3z9U6ofU3jqSclVPLcSEAHlaDrEwDEz6nGfTplk07lk6y5obs4XdH52lR7W5GfVg1WWV2g12G
P86Vwt3Hy0ITVVOc58BH7c8UAC/sfr7o0svp2HhWW2J8XP+8o991kb1OQjQtPgdUldBlqNgVg0An
/B26ntbFbYATs8b13s7dV8GxveyE4q7c/z93mKAakiXBQiPX3GEgiodAvO2a1v9ER3D1MkHrvHOf
rQIXE09mVNOG9/f0jvDK8m4/Gek8wi6POgj8LOYLjP/8uGX56ob91tPfS+cHWP6NgCnWWZhM8svk
Bt+BLjdGBcEnr/REhL5VIarphwfEhiteF6KwdgIsomoAtUP0vMRVYdCgNsDDPDjEoY7+8FGr+J7c
qN5I30ibA3KogoELZG8xN2y0y24ImS4bv6xFQNRX7MJXchBpUmIT+wsAoVUbrp1nOGno4qRGgnEM
lj9tla9CqIY6Q9iK6naa5SWPLzpgoKGj7VbbfKLUEnODytbZomy9ZJIlB5g/Mm57/who14RRw4KY
eNtDm+0bay1N2K7kjdsmy6PoZ/tEXvUfGYQHtWQosQTPynNSW0EaD0f8gxRWJHLCpWZIvkS30Xte
DQsA4vEcJEBBfNYjXz7h80dw/8tS/20olmIxVKDvY0bobEPQgO09zyvq8nNFCMSym0GG9H9obwcY
5Q+tOPeEBFE/5/Bx3E7rn9u61uNxEWAcSy0DbOWfQ0q2uZThrLQB4sfCpNkOTPRzRbt4jKmBpKSC
OcE2k3wdJ+gjHhYGQHrIjzcTssv3E0SFUzHFLfss3AebFesAZTdpA71O3hCKH0pnp5VnakxrCLwO
t2LUEa68M/xA6VfFgqc40S1uHhD3kCv1YtmLv8oQwKzCe2Ycj0vVCmv2EAbAM6PA/U2QuOROEJQa
hq2xOXE1DWC4/COFyUuLy3K8FOztKizg3VHaAxWWdLR+sktKWSGypRcILY3KD5biev++2ECC+5F5
ajFI40n1DcB79oC1OkNTyFATflzGElE310Mlz5jn2wg1sy4kMUo977iRhOK2DzBfexFJm4pf6Y88
dUD1/AmvclZ66P/uMGMlY8SC1LJc5WH56jHnFOKM2ru9S1fxZVIuLM/D68mRJ4dUWj3hLmuEEolP
rVmpd+a6TTn4dJpE6kEoqk8BqZQW+873PO8R8No+kDwpZ3rxLkA1XN0l77bTZmV90hkWxLLZ1PHr
+7bbQF92WKMC0uDHN0Y2IS7zEgrB+bNFAVxBucdlHBPKJ9Fj/iNEukXc9MqHT3cr1h5ja4GAfQVj
FQdTursOeHlVseAdupPyb94hrPEgpu8fM75p8W00cQDZ5p4H9JJLUPXsdXjBaNK1ZyqVHSBSPHvg
Y8DcojcURtDCYX0lYyb3RH8bQrX4CY2sW1LmG7kGPaQwR9NaG6WGvJYQkOttpuLN//fTE/LdWp1N
idjYKc7JHTmfylHqgYZFlW47nwWxsggw3YYJ6jUUUaw0NXRyx+idWwYY0NG0KBAVgk1+7VCMVLUD
ElrthGozpq2Bvh3Ky14U8VdxwJOVJXxZffBqSWAWRfqPJZaZRfRz3Rgu2dcKnduUs28BNLRLfXWe
+lTNJf0gGnhNe523ti7X755C5aCbhzET/vtFltsEahe7hMxFgrkkSja9sxcg9xz3oadRGC5JFQ8A
CYLCZIZ6RJYb8RUZmnzX9t0ihDFEjFAQTXoxnKysDng5o2yuFnN0H96Bjt7k9IIC0luyYlAlYRx0
aV/G6WwkMaGXM2Dv3BVrUGTI6+fviCw0kRPMeCM85ZtvdUkx+OMMXC849BnhQJodKVdtLSs9Dv0p
DT83yV/zmsXHb7YImTgU+NvHJoLxWK6gWByi4XiVAGHAgUr/v3wysAhzxOsn+Qs5KBsw7AD75yCn
bQ7th4LXifZ7YQOUukxn+rDMU2ipp9aOHfW90zPkXILzh0IIJXc7gQCbq/eBuvN3du8+taHHb9Yx
lt5HzmJkX73LunV0kkNwlTYD0QHsDsiDvJLZz7HDPujxzbJxskKUkjSiehnxjhYXkKXToavbbGgf
4FOnroSaFyjzcrAUb4IOv2DtPu7uFo6ezHaI2huu+12WsEDoS3rF4IzuNWFh0zk1N9fP0Ndu0rVo
TszOx7mdysf4iCJnM8hpnQoe7yOrpu86LL0UbGc/qGMW+5wYLypNWzHcp+BCuUHlZzCtJL+iEtOU
9JSJTVy3qRrL1Kc8EZ6EdgOpnDg/G7+VH9AyyLGLILtWMRIK5xt9aBSAJQpr6F0n1ASTWyB8/Ciq
kFJ/yUPQybsC2tM+DNzmpW3dVMUNewT5P3cNJ97Qf6eYYaqhGJyi/LxaN+uvjvfrIs0VXxJ0yznX
olSzwEkvEvFi1/hWrclZhCdoW51AWvzkmgWdg0a1s1J6zntN9oWTTFaGC1bGrUoVv7YNvclsrEXb
2YgSMEILUhIhZHhZrZrKfgEuelHUSO4fIj7j+CAOQbzT32YrsIuLyDhFohMxTIzmHbXAAnBbovcD
IBTYffbOGG+3YMwKkWOjVRPRWOjJFB5jeAQq9UUJrKfY324vApx+k4KCO9UYtszKi8UHfg+B53P7
z8sGTCG3xBvcr00mtoK0nKMbgaS9iXkzFDPbfxSUeSXF8KmEQeGXv1AFXxWi/D6JV4ZqH9uwSCXZ
MX6uXHB7kV9HM15dHRTqr68dn46n0shEE/QKawt3u9gK36pBOU/Qxn7nFJDpMcDWzrgmI9THHlpL
9WeZ1OYKQA4oivn70QwCWBfjJIUtGAMdg+OPh+8D6TcJB7quyQu7pF0jgl54C2btpeTtOYvjRQ3Y
a4Gobu7Dcy3QDgACsfhMcX/Vq5m7vrUeh+MB9xocK1wU+K50X91U7ncBZj4H8FR/37ASZ4UlaDIh
OznV+Hyry1kwoibiNvCMItISzXzYM0MyxOYhF0o/Fke9nOjk4aIavShouajIKP3dkhkCHjIeZM5a
hWeI/fmk+KKDEd/xTm5y8esaojWBJdP9q4m4SZF6r4Vjvt6ekDPxNsLMCUfnvvgcxxQPvmzJaB/q
Q1+joj4yYcinAJpFSXtd3BuGzp5TqMTTs7kIEiNEr3lAOyN52IteDb0RLDzZRW1ThuyN3J0l4Iwr
v03cFSxMTQSKn2mBmEwMExnFp4NVVk+0i89AWEY1IoQPe19Rkbt563NkMV2ikWWy/r+z13C+d8TO
vI3QM0v/ugavS9uZnXC530k+4fgPNiABZkOd1quM2+sgT5SkfULL8Cyk7dHuXPEXs0o0sJXBzU4h
1Uk9Q/i98nChs2lFGZy2WerOJgqTBPh/XMNPo4xtYOKyPIum/ChgCir+zBQQteHC5j07uTye/sjb
GnYZ+ulJ5PVse2tgXoTXEOT3p0PHyfeLfkLie7bXNcwbIb+j9ghnlaGfTAhzLuc+ZXCUH1z1VX7Q
98PMrL6xU9uksHu7zVHlDoBgQlDxUag5i0KIwfti0Fn4MQfFT2M2IkpUskgLsL1AKjKXgO2uHAmF
SU3Xj3PsW/2CPpsRcavImjkKxU81SLFHpPSKf2E/HfmCyctvX9uGfkM3+zixcmf6r4SczHTp9dyn
JLlk4lIoAcLa19kf6jG87cQhGN0tw4/FDEqyoNt+GuXy+TEcSwDa2rk/iScFVMpeD8Vq0LJCyqNe
H1G3PnaiOxI6qO6cMV2Nl1am+vZWtdtnbzsPjnPFDqV7cIN10NY6Z80ZaEq3VznngDW7JY4jnsgK
j87x2vLS9srk0o4RDdOc6uXazmekRSxsSQTh44KVrRe6mIG49kD01p8YPcKV2/Pue6fP9Lw2AzdY
Txzbh4QiQ59mGiWDSkb3U2QlQHXVfaXHjbEbGDFfReokXsI9qoYFJo6paKp467ulKNyd0aF1L5Vj
O4bgL+zFiyG01aw8y8tmjwcrOCpO9+hJNEVkOuYOQ+9a26A7s8goK/5VF5oAgTcoOq0oQ2AJ8Mv6
gE12mKltP6Ef21Bnyay6SJclnReBLLpzwRacCfXdh5JyP6MxvJHC+/J440SPmfxJhwcZmNVjw6mO
fLNRTwXrCLQlNWteBZ2/L6jNTJhfQzCOw9u+LedQnJKyTRDTXEeYWZ4yFFQUYmtcd5uulHorEzUo
lZc5uNl0XT/GuGp+aKL/rSEdWU574HEXePH0ZxUTxAiyD1WDLBWwFuMNCh4HUPLal4MxnsUgO/Xj
yrBoD/AyEXUhrSEAVHn4JDUcqxpFFJwPZMj3o1RCMq6IWJjRtltvAYeCCCCm7gIzjI4gvKByfhi1
x1RvOOBaNATNhfb6pY2TPPyNxHFN02lFGxd8LVzPqTKsJbmY6KOZrBB/PRqiqdzpHnrZMOWRRpOP
GitHLWXs4sGmZco2vbE16YzpYlDLV1Lc+0gKe/mHk1KIIOIVa6oeqq8uAXhvfqqlTlRyoWVU23An
tScgYFXbD8WC3OfM1x6WKptXfKKSfwHTJWzc/rSXzcljNDxfEUv/NExCaudrWEqzfj6qTm8SiLtp
soN8Eh2Sa/ywZX1b3B1rv7eUFkkbXyazi6Xkf+efoEiwDmlxkp0mOaq6mKan6cx7hFnsd9fxNYwu
DlZtm7An95wpaGGP2VkuyOBhdNVSTbEMNZI8baBW9D+OBZGrcowQbu3wmvA9cOwyK7NVe9v5OC/d
bVBdh9NjcrzHQD5WzQyZIjlQlUDOVP2igyEEcCbgDrX32ibvg2J4oQA+P+L2v2WA0p7sXbF6+g4j
mBma1RIDRMayJnj5LwZxN9a0dSvs8WQZL1TpCreD80qxKwMAHxVVKBa1osWICTAKJVGMsDJRRFws
F7yULo40Ms3zjI5DXBbk3K3A3+onC1Me2eX9N6/jzFj2faUOnXOq5+/gNVtN1kEb+ycZBYKAshWi
FdZKmft8aEJgd8Oo2tB7dyXF4zSiJzXtY+oTtTjBYtvNNSJNJcQOJ+u8igFP/9ULoXIMIagEPGbw
UgAVlFZZ7T1Gh7z04ilOiupL1eI9WeMcqwac+ZWFaSCNMdL18trNGhc8Ngn4xGtn4fgDLBnyY+9j
GBG9tE50vNwWDi3fplBwwtAPkm33gkM0nbdyx1cqHrprUupxvYEHZ6mnBdbWxyhVHEl9BkT/WSob
U/m+izy3EiaNCJJYOSXeVi/kdgxdrgV/n9/mAQkJZXn5e1WSdV9jjNw8hWsvD1Tp0OHlk5t0C9oI
XTLYfzP0VdeTYDe75EyND0VhtxHFNYphiK0jfwmFwCnxp0oWg4HsuqUGVcc0/81vzqkWcgdLit9y
ITXoc7ZZJuG1cLbkUZux9ysu5FtoNA2AwA7pzTJAzckHcpggz8Pe2/bc5KlnyMtdcCy81Av71qUf
1121jabcczSF1aoWaz63k/P8UAW3MuEGvUQNQ42XSg61GZ2fIZ4bbl8+8gjZJUbj06cQ6+wJtR1H
wYFOoy1BAHQlmRQdrOe0/VFCX7RxSd0vzFdtUv7K3WdSYkNAcBZelCiPv/8UOw7fzBjEz9jt5M1o
SSJO7oalc++azkMR8d1yRvVH6eStIIYjQkLohvFmEGhqv+78mdVsdDbqsKw130VbB8MAQXL0INbp
CdF0D/C0JP+xOogY36sKYp/dSAizMWRsoEBuSSQUoVKIEEjSGoe1fO9A9/iQljyf4iciQFJ1nZMI
zmiWDXv4+ppHLYWAIxJIQO4o0I90sbo+aVALor2YcLDVnUyOSVDkXO0YpIBpgtvsENSpMtyYMF/k
0vlrJ6gjKRoM6UocXhb1vWItNUVFVLDNK2RdQC6FD3VLXS83MYCXLCxCQ4f5m5IKTAtrsVpzW0P0
QIlppdnxipaA8b76/drIVf88BJwOFe6n/jNzEptVmPVYkyyLGAkMNUkUf+vVPs6CIrKz/Ad9u46U
XpH0EwBuciMz98nQ+rh7elx1UJyL5VwMFs0TEwRp8DdhGbfi5naS+Fiyry+X6vPUNoPNPf9yEn8y
2UQ0/jAjXP7z4jaRJVh0V7zjjJXuxw+47RIkFU0GejNGD/fY088un/C/Ls7e54zG1Ur4jo8W+PRe
Fd9UEK8O3eFawWKpzMLHkOE73KEm1VGbICEStmwWcNZ9x3P1OMeSuU9U3YKo12y71QkOFehCx6fl
gbuxB/KQg34o3rmJnUkah4ghpPn7nDSFq4gNWHTw8yOAb+c52u+5+5wFwFTDPFTsRtxNw9jR2knm
u7ps+dlm+sUFcd7z0lpB5gnvnWzHztEbfSYWmFjUpf72Yf6bw2ANrwsinHHztUif2a5fuP0ALe/H
mCR3207T46xK3hVghw+hE2+J5RNqQXmQiHYHK3xrHpT3a/19pgmPErvAwXaCxHwnZ32TUsJjjbj8
NdVqTXeFt8S9c2a/LeedRFd9BxTvQ8dDUTyWXdw1cbevgzHJRUgKHy3hpdjbYl0QYA6wwuzK+7oF
BQHpmu6uejWTJOV+e5eQK2XlDS/gi1RS4MrS1D8FkP4gYZI68ZwnF/KcrL4c77o8qpckxoNIQqiS
Jq0t9Oo6BrkWp4p0Cf9TyCgrC5nAtDSM7++JR5RCP39i/2mgQUc+IektNSnNQQhP33tJFJOqJOP5
M5JwW/03fXOX2mdaJyvEt9TzGszTeeM25mzyj/3LC/kFXw2GEQKOXH5OK2/oVHa5yBnQV6AK4Aqv
upCPACTvZvGUY6hb9G6FfPB09o31UT5WKm0KDZ5vONkFepDKiGnyhpw7Mu2jswu70DqL1j6uJeoG
QhpSxklFelhLZbPFQC0X9+zCn4fAtjZ2o86fdXo5E3kn/ZFYUbGRzSNpkCJUZXC2sBwBqbjuO5q+
68URrtvPJJr+FAjrb2RuHNHT8UCZItmd5rX3yCn8cS1OvWmTBSyzL4pMGTyJsP/QM2jBuyDCglMQ
7rjw2CrMhgx03BvLRJyIg37unxJPnc6IL3WyfsYMuNBPgHIleL9B57HC5mQkyaV0hsp6JNDvSrxU
659l8zAH+SfJmhBH0QSD67trL9moV5V9TOJ/PWoi5hwii3v1Qqk4NVYJTsfiFHKX1rsg1hMdyElR
GBUEaWDTzxQxFxZYRBd7Ec7B0fdakX8TMmMONuN7p1PneqFZfU4lRGGqDSk92xN4YmicX9YekjYL
J57h0U2O1BxWjyllYLY57bdJLwIL4RqeDGKjw3gB1ZbCJ6Tf87v85MtCPpc6/Olm1YuaOpUu7K/u
Y6w0BR/BiscpTs8FIPZ/HE10RDix1nPfvCF6Un73mlAT0ZH25rFzyGb4rHptmgkDjyIGs6knZnHI
di9XObFtMTMyK76JwBGz2jQOtDqQZB/LnicQK4EIcMkTIyas84urdo10DRkpGF4r6/CJUf+V70DN
feqHY9wf1gps8Ajt0+tAGKjYu7w1R+NCrSMaLSZ/QPt9LQRz2QZyYgWGnlV3FAM7VBMxJI/xXbob
PwM946KSGCJnv+LxQUUTWNf1Qk3MLGC4UVR3NVzdFhqPnsDVItfY2KoH+noQl0VHru+R01kYcGvc
dWKWbQYe64uG9E2sU5dJN5wQezmx3DNUdf8pN1Xh+4lG7WRdTA0VJNrbCW/NDXY2JDVOKNrdXyZB
IqkzFNp5+ZIxfx4HWtMrsSlPtIjxQCPSE5BH55s6r1KVEh4rsXAqZixqMsTWMNjP/R7RSqGyExyu
NHqt2D3lZRTyqVLxI89XrkncaY/bgg9ZfOujcLfCdn7Er6oavAqaRlN5Pv//1v1Fvu7yU3hMQ/vr
05HkIWBrjqsMNtRQbmWADE6amzuxB9Riln8HWO4ZFhytK3bAMWPuoqbF2BeICN6aOFBV8gWnfS19
V3pgN8NmbJbNocuxDY8WMjyJkcs5ox7eZRh3M0OSB4vEJcyFkwkCQB9L8hkLLaY/RPHKhGZWRUZc
6LLoKSjFIJLUOoVQwW5umRWJq0kX+UJQljDpZO53Z3PV8vmiiYk0ZkjjrSpqPgrkyV/2pSmNwNcU
GX1sHmF9AG9do5jh5mEcmx74DgX3xfLGkV59jO8+qVMDechN0pP7zkvX2Ab/B8r3klid6yqF1ri9
UXOrauXdqAQ2NUwqEu8YRpz/rLFWYy/S1kcQFMMeFw216FgNQFWxc8O7Q4+730MhmWWaymQZ8auP
e6/J/C88oTTv75uFH+yu3FylYoeK/DIZjFVesY7n6KRz0qzpDtljwTqcy81vuB9zLCKwGAW7x7L9
O6yBb+yzUo0M+YlGBTsrAwHJ7zzl0agJlNYsrEd59XOrDZsLU7ydeWuqW6PXX9630iJf4rKLqkD2
SBW45VEFuNM17ptgp+ruDWBp8sylld6TDbK0ce0ZK7y5l3uNFOyylcYmoauzus+fpXX7gl4x29bB
NQNqUWYlKQ/dSEV5aeg1dgxwDIdQTuBQsAGpMDIXMlYsQbvjDAzxEW3FNe/DpRpTyYfMSugTAZ9p
KvuG4gb09SoLnEbDLTqkYGUfweJISyvsCviFKwy7Ax2WE8SjsMEjlQRVWOz6/6g+FA/oe7lO5CEf
XJNxW935m874K/nZ/gEH+ShAC1zTi7qf7Q3HbZ8XSQAXVd+oW9LeCEZRp9l4vYdf91IwTfPFUnxa
0Q19AKN6oXtzTb1/A3Q9kq/Ck7LNRMg5K42I5EUNi6Dm7X3FWYe51y1c0a4EUbQ9xBDngzq+QjMA
ATV827pyBXwVm12BnnxjVv9j8q12ei6t/RffIUTGhU8GeSPgPDHI9UHTdFihoCpeQf9u6tzA9npW
5e1S5UK4yRtWaKIBN8xYWY1iXgNMMvtaw87VutFVCVRsSVTSDvWeqVU5Y/30+v2W7S9+ouyS5MbU
RFXuxomyTtFhnyD4umB1oK9NcIdpYFoth3wqvOUKVjEgu5i9VZwJ8E9unCjiwhAxROzcPvxnil1B
kI9QCGydivaug+i9OpmutWH2jJhJEfA5dB6YipNcss4XZI755UaMoBXCg6oNP7J/Le1l4UM7FUCF
pbmNCM0kl2jsYSZI/PVq+PsVA9AGWeJqaXfwrTIEGzbg7qjUvtFoUJCYskE5wfjCr6OUenJbq6YS
iXAybupVbfUvbCn+k0bw7qf7GhWSn09QEwMRNALx7VJNxF+9ArCkXYkV3Dy7rfyDFNF+rVc+ktyS
hQQIChYijrb+EbG7a0eOLWFQ6i2JYSfvSDboercXdJsyHHDqee4u9KaKPNV0wIXkEmMJe3sbsytd
wFBAZuSIsrRLjBv/eUtUtpezhe6EOO9GaPCQ+yNZHs65cB6YK18ozp7BaX8NXuzMPvre5r1pxgOD
70P5g/04tKxyscOJ7CtcNY4iicpyJj7ogk+Y0qljqPVL2RgLpHgjYmAHNxsYdk7lEytm6VhQr92Y
dG5A1/IRCXiFe8TB16lcdDLRGd4tYT3H26aH03AmBX3ik9hpRc4QMUIrzQsj/+t3N/Tpj4y8FSqd
nCE83/NJECVzCNHKkfmlJ6FreCAYvzeTfrecJUbgOkVpXA8Sogqo3jeL9jiPvJl3aTmO6wsrQomk
PD33Nouy/UQPwmg+nt+iYJC42DSHYFMUrWD6Hpd2v9RIXP1grN0Bh++Uds4uB3hMK58k15bBW0O2
lg0c884cn38ph2L8eewOnX1Oc5RQ0t5oqa/3uDMDVGfEzkHyY2JcVhRV+vvQySLjqziLOb3mIfWk
GysRxoFzJ37GXOUz/0udruAgY130jvNXUDA+cmzvngelRaskByL7e6jwXXluteVNdp8W4nKX1N8m
Cwi9kG5SDvO1q5kQFcq1txcPSTYw7nzNGPGDux2CZhuAfqpsNmP+exsjh7fmfra/ijRjkbzmKyPj
j/PxIfO4WlLyUUmwkaukG3DyI7ZRvkfGBMeBeL+gUkHF5XRuyPjJFK/h/Z7qAJuwHdTvpe8P+fRL
s73zm0K/nY7jY1E4q8uNXVkyNbvSzzG1XHrDied1n/Om8p9P1KdDgviPy/StDxAurzHGYPh4WlGW
5w3sCmJNaKJ1msoSNyawBvL7fMOCDYLVb1n87H8ageGQO2pmEa3lSDlsG1z6nf5OW4q7wxYwRUOg
JQVq1DHBqgel0zDfUV7MuRqhwq2qs6Vjv9WG7vPX0fsO0DdAY2Q7VzZs29KCfCxLrAqLGLtzMZ7w
zTMEmuBuSNYH7TeNE7YTa53sd1Fc0w2x8fC86H57tfIfe6dNnWhb8zqB1gswkGqV6KgZibx8DUSv
4lNGuzEghVFEfrr34PHg3xbNZEr8FqgjgzCwF7pESb875zaDMlR872pLI8QC2QSz1G+775Cgxr6P
xDbqZUpmFD2cT2L9D9StX1W5p3BLbaxh9cOxS2cplW2HuBNa+irTGvnvxXNDO88FHoueHboxAPGq
BJidLHQMKZCqyAmrH/bU9dyrnFQ9e8C1SVT+e2qM0btfHqcL8VmamI6kJXytpH8GC0/DSuXHmscM
RZqnVgjqHYrXImvy3isDKP0NfZfqXByMTQJ8numpXQmVoBKh21Fe2N/Px15QNeyJFZArKS9eg6d/
QzeViFM1cgz+9/TOm9nl7YGfbidRY0OkeLvAFTuaCxdsafUxmwdOfLc8afe8utG/2pDCNgeSIGot
auZbu5KleRomyAOHhDejEGOYKq8TUvgL6ZREzgxHwgHQnRAP0Pp9F2UhdBXGA9O61DBf4ZZPuNYV
E1iBIpHTPc6AfOn5iSlma3F7I4/GzbL97mFqe4fCqP+vYD9YrOR77OU8TQnhnMU9Fu+yhKiRxCkF
p7LzKeqeNU/kGY2/vHyyLsHiNXHCRLzIU/3oWyt+uSOUSaGXz9eUzQslU3qRbiN62dTtMb3CNP9f
GJSVONZfbdPjYIXrT8Zl4SveFbD8ol0syny02TZh1Tmap7SBgVMIdBmb/Dd3epMbxK54tRXLXlH5
L2I8jTqBes0gn/pwpyXm0a9hPYc8mEmfZMbXgpwHbsUy1JVhOsjmbOHZNLFiscuyLtz72nVyfRMW
tiff3ysnz3+FgQ9RphcAw/Bs/6qcfOjVDpqXtOtZ0ST6dv1k+ednl/ZC68lNIVifhsuj8aAQiWbA
cXhkeao7kifMeekXzULQCMPoZ6uG9t0UWgA9hV6xpMHIvZgc1RrVpNkUO338eKTBO7bQAFZLzEGx
y9RiGvYsOcdQt08WXQU9pSItxABgyPox7LbgvXvsQBP0amHfmKjuomADR1bfcbCBNkHLFNUu7dmE
MX6zKXR69ROJa+usYyw9F3l6Zrk3B8ER8590aG+mm2Qw8KRP2DFg6claXZcHmxUhM8q+/Pd83XV/
31scHwTlWX1fsaio82xVsc9NIVyY3jC3b19k8mlNzHNjRbdcxnZvDLwpqZ3cfYjxJvcEN4bshUAF
NXQQN+Tnv+t60z/9DcIg5BqdTne4ej9LJRecmjLHQq3ooRngIhclJa1n+KNSU97lZHMJVIhCiH4j
MRr96ygqY5QCIkbEySgWP8Gj9lQbJbOLPbw7+fYoO1+QAWcaPGtRldt+MyLBUqr2Cwg2oHRlLdhB
g9csoo9ZAUty0ogZNSY1IXRIroiAU5ePAynRHho4FAkFsEdelM/FfoxFQbnGCLOOiTxUsfyEvqfA
iOuMPp/dhaUUKhujcjsOley4N+KP0IiJ7Zn6a0l5G1np7RunuV8DRt1XWr/obOD876oP5U5BPOzX
8d5KryFdPBHHQ9Hd7mEHXasw9sDilxDHfyHd18ThEv6LwYOS/8cGTbeJfDhtm/WuY2QS1gQSqUO+
EEu0hy8gHq66SvuL9qU+d2+Ln0E2lQ8k4vE1ieha7glmSUv9w2QWhr2ejTuSxlTEeOCSi/5+Zvei
CD4YJSORVXhZ70bMG65SRDikgFDqnm//Uxddt/F+iAExoFvdB9PBSF9pv4TCGro28Y85Id9Ggzm/
tIZ/ZgpvpTLiutlhBvFSJy6Ye3wT0gakMbULS7CjwxgJqrME6xRPvoQP/xwvBRIRVHuYeBPeWa6V
KiTrGS4OdyXjwfduXFExYU8VBLixxQ9NBxI+e99xqr5AQvLoF5cs6o98YRNI7g3OTnhopOArLgwY
Zksi2mo0WDdtbrDWOnKHkfx2esj3nCSEUA7AN5BRophNNWVUmAJPb7PFnCwfgdlE9E5RM2f0Ifix
cxCPISr4571ki4aBz1rZVhKhD1JCFzYdE/A2WgixqHDhkdCGZE+TFSzaUGoghzDDp9cI4FI8iA6h
sK3FhgonOuidyKDW1MsjzPm6rTqYIHV0SX1P+GVf9q39QPTI0TNhiq4kqEYupc4WqdOIN96UiC69
JX0P2VuSafs0vAIbwilW8muBfJSsOcGuJRjWs/6cRSTnxYMmvcTaNpzERP/u+U9s3tbsYVdYnQYX
oDNSe4Wof4QT3wlk4f1eb/nnDLDKr81FI4KjcUHRGEQ7W1ucSlGMDvS0b3s4pCJVZNg7C4aw8tGA
nWtQBEZv+FWEpDOA4vxQk8DvVDpaUs7R1u2I9vuzwDR5QP4w4HOQdfpE/1SqmdDKcr/QzIzAwRa/
SRkbhunufPeMIGArcpDJlXooVRetvLFAolZKC1BcsH/kzCE8IIuN2Rj7uyqnGoeykoCNz65PLMhk
7NsRdnbfww4xp9tHkKrBajr3ckGpfRmG4fRMIO7+SeHooeatZqy1qAZD9d6J6qnIis/53VJ+JMf2
znOUpSI1iwsyEBvgDecF8y5tbgOZi501KAwM3hvSon9UI452IBN/B9Ma+OiOHHZVRhCaRHKdtpzR
ekmJapTBTKnnSICuTCUX5o4/4olJuIVoV77lYiU4X8cHbr7WC9rl9SkW+UOTN8ssChIqGHX4uEUp
g5IcYHY6CqhP86ZRnAqDsk2ifL6lDEDdr0mbOdSae9tjV7DrgODJ2RM9+BWiQfZ/g42ePs/IWMBf
o5loPua0DRs7DMwVhyMdCAgkKRHRZvioA+SmBN41tBvT9p5aO1AJFIuwicxm/afVwBZHINX5+6rj
5MyHdRSPm+zzBowPXkJkrFyn/uZiOyHiMhSjMh1pbgKZko7GJNZdvRzosDkVw428fRLrJZxvod6z
FxsGajQ/sacffgB0AL6KHSUHheeiheVMlLum416tO/TnlXANIjcnRDTZOIjNf+gLt4pc2fBOnWoh
zZ8uUKXsT7oOiljAq5JDpLj1NGCwpD0/bGMWoFD57RSmYmUKttg74SUk/hmJ36FhLjJ+l6nlAimX
0m+Sm5H0Kt9PUqKTDHiSJOPje6Whll5saIdVeNvAroJ/WPF+hdqbmq22VglI9JfMnMJcMOcs7iFv
An8BivbdiytV+YAyRIERo2xdhs7Y9OZ4O8zffHxu+vQ+MOJBLrFrIjl6+EecRurAwiPlMOIf8bPv
OApDlCSwuuQhTobaIDS4OOXgn6ehDbuB9nA17R0Mox7LMYB2j30pkJE9R9ZVcsfUMBbvmzqiLz/G
q+btPIQJvNWryZVU+OLTOnz10neTdH4OZRSTMyZPya1bPsIqfcFfne9huGAEBe2ElqafXzjtGXq4
Jh5x+EvaPYDhPnSOciegeCJYZwTAgmz/DMB31saiXwp9o9TglPk+ThUb7Q7gKqKDlcE5928u4Yxp
smQEW2PpocEQArkfVlEeDBWGZ/1u7Oi5SYUjPSoq0hZKwU/EwQ3iZTfotMujhSylSsJh0PxCxEY+
EnzbtTri7whvVhtMAvrMt5+UiMzeSw6oAwYMgajTQU65NFqtUtZCrkxzdTADWRpTKOrVcvspDXVs
UZOuf8BGWV4MYYdqvVHuJ0xAIr+TcvyIGpNXcGANs1YSVt9Q/PuEokEaDquE7k6IMAAlWcUbhF/T
G9D1Sj4ZbC2oRfyiUFlyGbPkg2iXjTs+UkSnTjdvmcJBCC8MlmAtY2X7PcH4zd4p76xlHfyFrIDZ
zmPcOX55SmOhxthkpT+cUgysIiyhhcEWJ/9in4QchLv5lVgvFPk3mZmJkAkiXf2sL0Bd/dwLhpwG
vwkVjZcw5vf5sRBvjp9Thyemla7ah4xuIO5xxd/ZXh7IUAggfw4bH1EXwm+i8PGlQB9RuhAAeJrv
uqtHMuaXFpzgGoRjHKvHQYXpJQHJP9cyw3VjrfqAZGn9VB7B8GS3fKMKwokJL6k/TmkbFN6CfpV7
iYkEIzhZDtFoqOd9lcZN8aPZgdgBpApuzn+EQxIB3GJSrQd8moG4ndCBWGm0lsASoiNkykYcqnuA
+3K9pLJjj3SAZShnhSbItD4aOIUElVvXtScVZ2yCNj7Vmd+jHvr0d2kDENQi3RIESyVucbqRo5La
KcqhWKAbSmdFQkA4my210IOLgz7sbuOFGc0Atl5zKnHI5mSsbo/Te6m7XoFu4mN5BgVLZDBS1URb
6G7BMMu2ULxWdpb0FuRjhj15LkmY7FT/i6c7AvuDcaEXA0lxOvZUVV7hrzquSOQ8vi2atWNqQFUo
50IVimnNDcvwhaHRpTF8OPm+iyOv7blWf1QB+qaUstUY4YT3FlP3g1qgsb2oK0bukJu5Ht3kb65w
t3IucwJDp6wl+40JZ7Y5tgm0VKaYX4uY2x3uGCsI5r2Npq6AQv3uMYMMZVuNs8y8z38AvB4qpkGh
V+H0gwkIJv5OHfEJVLH0QB8F+1e3ckgu1r/MqYrihQai0yQxOikR3cppnEauxk9Cyo5v8fuuh9tK
8n3Msj5e2X76Hcf2xmgS52mmeiC234RYjegSoMS4czKyIKLMyxzyDx/bpz2ZoP9UsP1Fzu6TFwf6
4w8QOdSEpiJquh6GPKGfyWfrbLT5cpXHln2GYdopLaFW2Aoby8dnV+PD5Vx7R5m+8z5jM7FWWpjN
0FF9amTkZYcD2MR1/F7R+pbT3sL8Y9PyeZgvGa3Fl1/SxtMvpu3Ejdz5Opjj7ywgXWa50wsB7XrK
1KSUALrsl6f8gHdp3pzjNzk39MuucHXx71OcPN4rIf19somZSU2sp9QsHcAdeg7UhSqN9c6hIKUU
gFeJ7GJWgp+d0REsLFOmi7stGNtfOW1YbLuhiFsPJbyzyHfHu9lNmtLKpj4HGKw7OBAsR/1Styza
bC5i2vC97T9UiZAKKLvxacKjTEH00G+DARTi+Jvwk+iEQa/2naHcV0GR4WxUo15hoxM5aK9W898N
aAqLW9CQt3V/uwGvjCk3die8/Z2SXpbl+8iyibsMza8i9N1VjhVJYnLqNFUpJLak7WuUhCCd+3aj
3+4dmngIdTv6c35F6MQngwEK9/5pqi1PEx429hwgPrtk0c0Fl6Qk1CEGU2taWE7eZwyc1EHde3aX
V2BqwIXQjCMI9W+v7jaDvj625w2a4TA/iHGvRuU7s4T4GXtWi71M1hCM+0Dof167hsjEWAKatWh2
gdgSxQsTNSkTxYQ41w4pvxHUV5tAppRrak0n/0dzTyYm6rm3RBK9gzQYgQcqm3csJ2pOPAeGhCJg
hsbmhBkRlQZNeEXADQL0gDD/HBgi0EiKv9d2i+yKnvc2IxSk2u7Mzz3Osow+NSltSdHWN0rDREBU
XeouPqi2SUTzboe3B2jBLDhrN8yFUcSbjfd3xYaProRyv/KODaOEd1J9sueOwYM2vxL7Ad6ygD/O
37b7jKO32dyNpsjGNW00vFtK/g+XHaoWZ3n+QjPbTyFc3db4tZ/qg840YJ1Gy1OdG0ZID7pFu48n
z14EAuxuBfBmw8t34c6lWREqm2pHt/MhljZEKGRV/uUFu53VJOzDFpHNeRv0HVyPs5CC0CQm+LZL
Ri4oh/5SOJrsjkPBK/HuCdZZuqCV3dvwch4Yp/CL5+ZW/X5xHJ0P6p9YTa/4RA73XAmE2VRhjfjW
acr8J+4d5uUsMRT0+0UxVoQcc9mXYmNmN+NqM1YZRRznJJ7MMawTNo28j1lDdw2P4URuPIdABda/
ScpkASdpOCgJyDl2m8CLCJnYjSpHrCcAyDNWmpL4BI/a7ePKB6tOT6PtKOY4bJkxf53GoqEBvDfs
sAyhMAAC4OH4GiTmY8YjXw0W5KyKxy+eggHNAHXiDRvNmWkxUwzXfOP8JhGM7OZTihnZIyBmKCfR
L07TXe4FigslldR722E2CD5dC32kNbMofAiobLc8PjAoFJIFN9yoWVnYIRdZO7mYxPy7idCxR95c
Q394mOOlchlbVY6kBmII34jFdHe4g9/RHtAAzefkWMmx3uzzsIQ+d6jLc5kJmFQbn6qkYmbjl71c
HAZaKBKl5wotPRfklosgpmrVRQ8Vj+oC2RmRsbHFSJZOceUnB2vS2H6vcdokFSNxtslmoCzXJyxr
roSblG2rqa89A/epCv4rUwGV5zLrP8vMVg14eGpIbUy/5ea0k3tWggaakxRedpJBgcRsn2pGwfGe
OQXHi7nnmFgnqKZKc9KzklWVK83LLUME5RRnRKmryv3gA8BmsQ/d4D+Ljibfx2j0BLHFm83pnf42
NuQNNMcGtpcsQXbYATCo8Js+A/cWFg/cqd6YYxRAc4uFYltigUb9oDUrdwmvLyT68fDu43Y2TxMy
Fvv5r8B8Oty8SiZ6wNTVn1iLuXGbQ7B6AD3dAxVCb4UuR7z+L/xpmwZye2S8u9v3SHDt+r/qOEvZ
C/YjVE/QTUa9i6eEtZWFJltu85rqjBqU4cP1e6iErRuxDYi6tx7aQD5xROsJ5zNrPFwPBuUJ4wfX
EzF8hS7N0bN3FRA9kVRAonpe/qqT2/d+ufXizDuatAF7X1zxAXWzHwXE5q2A2gWmVtN9KKzTi2L9
99VrfwEt0ebsatb6sKJaROlSqYkNH6PqJGeRYs6R9Y3soYJqbTj+0pNaW5DDOVlkEfdakQ6CBiEv
XxE6A5IXWUXrjYv72W7fZmLCEQRFBYV1a6bI68X6nCHNYlu06nu50vmZ2wMImDHESPntmHK+QI/o
MR29P3XFotxPACt6x8zPHmaNYiU1AkdRswXodUrfy+z2WOqtfgL3GN7rsThrcR+6jyW38f2SdnH/
GS3M7EamK0BwKZRODidAiThw5CUHfX48N980zkTnBuGQp0/4f/vtonMggP/GJIo1gOeWqrkcDi9G
jx9yJom1M+nYXGVw+YloK9nMrcMJuieGhmH2Nis7KkpQT20wztyGiiLO6/0NIe0LZ5878mshGLER
U6QvLVFHIksfsS9v94PPA1S82zIUES6SEY8cww22ufhfg3kj3Wz5bsZigO3ev5GbISqGCxbBSL6n
owbj1/YNegS4YIi966maEYUsyJ0f569LRvhyOPEbP4KiY7DyEN1ksxNdk2APPp7uW+QGV5n+kEfY
MB2jp+BVenQfgWWgF2UyedmfvAoZ/1XFwP2qNi6NB4v0gjNOAXEKcnCYdG3VMXQjoC/Kcnx9gqkV
PerGEGyMgL00qluEgp6mGAMvF4nXSNy3GB2xvbUy6INfnqoVS+89y1zWrSzPZXupP6mAV8XcNyj6
JSl/lxZ+t6E+yhKul9cn+9RY7jcRdnzEWTaaoyg8Q+GyKHgKn4wSc0ZB7Y3FHpiX7AyiOQaLeVcx
3xY01mJ9fuLyi+1scaCWThMs66QWlDSGtWV/FpHA5ahthuPOMXUHntXT9mKOiNeUQ5f7rlHrPQTW
yz0lCl0L+AYY2oGNYS3w6HJ9D6M69fgND+Au6infqJT3ZtiNNADqgw2brMi/t8wwGkr2C+u9ZRQ1
wriKcLWA92UiWMs5kbUqNd3HVQub7cDXBpCohPwO8qW5O3V+I2PAkKSknus6MvBaDmTGJrzhaKNK
SidWO3asVkiGWenYJujEfj/rNR499zpE7ognR15N8Nxrf5z59dWhpOa+7nlmGJyqzHj2uuBYm+fe
RpsYkkiDRbbRrgtigM1/LQcBskKcfMRw5/CHmcauzdoK5E6sr6cOCVfZwJIvxQRpKNfRZM7SS2ym
j90d47BR/kMycKZkRgzq2thZUhsev5ByKL3xk6EUgrKSWQZpTPHT3s0Rk/RLj8vzuyaJGiZDvHU+
6yMuCdnp8NkDme5g3ekm9tuD25Qkoc09DGmJFQMLsy7wzg8bxc2yC5Zn2c4F18D4NYT5J0RHvnTJ
/U3/JPwW/HNMbo97zQcx8x+AW6qxn0F0DrQFdLK5ptEgOwdaQGMGO2+1h88if3AvhbptHYDM5Xsf
miNt1O9YGpPeBaLpVIokRFq73qd0I2iSsgU28TNj3mE4KmdIUR8GkFh7LXS+Z495NNYnN1O0jWfe
v/PpL36m1cq6bz3s79yR62Wh2CSOBsrmlz6aFY6zoqjsuBsPyTwPAOypqG7zLbZvLkMtdaS1ixOm
f2mWp6Bdi3gmFJb7kUFnTwu14C4RigBgmYIRPy3UkPQgO/gv8/DMrYcI+w/+gLCszwoqf+4OvaRx
agpavhTL1KHrOZNZhHLuSY86I5efC2+JFhoE/TWV6saSiahw7iEaKoyOyadE80Nr1+l/IFjmb/SJ
XNr/Q8qx1Ppauk4KyVqnogcVOAmxzPT8Of2bdmmdfQzncxO64r9RahbAMIRznUlLHeBtNx2of0VC
Jj80LYa7joRKTJc0KMAixMhec6Z9zdyWBpO0NzKF9NdSFxHlw5BmBA8EpXRM7HzKf5M/pEOO/7pR
5/AdL4anmve8Fl9rXhgq/MbD0OSKbLt2rA+WCpxsax84dYNf7Bo+ufmi4zJ4M3lR+q7VfxBtnCHF
eCsAovJ+f27Wci+PsR1iq20H9riEiJ0n9zGDM2qwEZuopAp8SrjrfXCg8o773WYyWR79AzX+EdqK
uTY+W+sJPC3duoUuhUpsWCIeJ8EKb8MHNtN8S+ySf6ZoxYG+9HzE9PTAy3iNu/ZjHX73OO3V3qZz
oN707Vk6bROtTCE/0StF1HK0nyGeKz4aGDaOld/yJgX7SHhPmPHOMMId8XWGTyh5e0AdNeEL9650
rIVQS8Uxyge1voM88tRKjAkNrhoD9BK9SxJK8qLodQcDELnVyXj5poyeFd15eGcY2YY2XqGpZjRl
/1j4xM3qHXAYd77gqWynPUli3Kin0q+vvOO7kYPmzAsm/c8IJXIBFYxZzXMWSwSETxdzri90tyg0
AKinIQsn4bC3eh0T6GDedT2heby4Zp2/4W3ddCQ3g/Hndg/nQ3uRt3YPVZ5gykgjk3M4OehXejcx
wnIfXRYpjHmjI85jLhhRrAJoOQkpEPB7paEKwewlLiw+1Mb+TU9IW353OOBxSyyBmlh1Fj1qabjW
xKtSD8fT377UXgxUxOqOVv8c028ptlc8eqXwz8prQrBmEPzXqr36208sp8raF66cTx/rMIBnT1bc
d3ZGm/TUU3IhV3JKQ0HppqKcZTJAr+xEUDhif89YkuPtO3gKkW37CylrgUKgXi/xlcN25GR3ZJJ/
KaMlLFuBh+ugC1Qjmsc2bG/qtnrbFtZahJo4/KSYQG3JEJ7nM630lMblcaq4Vo2HW3blRFJHQGPr
ZX4DpdmA5xO8VhDN7OltIg8Ro6Md9uGi6OBMyoIcY0XaBEvyPdjpnUGklQRZjU9uIZcoGzvM2ZRQ
jtbLRDVryM9BPfr8epbL1PfP/PzoZdmGrXzK8qcwtg++5QKVfnpVxip7MOxaOPxxaPlkHoJr/x8A
zZcd4W9r9nk3u3de7BtU6dwfk8+8TAykxNk7belDufcTRS45A0b/vBLGsc6ziQRt+MovhtGJzDwl
wAoyHmk6UXy1lvWS7J49Z1F5GHWXcK2B/YtU8oNoGzKDGJvgIdf+LGs1JClvOoR+Kqxfr+84+d5b
Drjcd+bj6Au+qnFItwuglr83PtojySvZ2W3Kyng+dtmkYhLaRZkW/m1wZ628azi2ZB92h0qlXTFp
y/mEOZmjI3BP7xPIsRKzlCVT3CrudKPEDImNfiB4BIN4whTPU0+9WY4I1EnAfZqkYat5KSAT8OzF
NU9geNztejkr+CHF4AQDJ58Lvv2HsQ/HQCuTQE3iblqFGJ5PpmIeN9WPIiMOXgw6vCr2/3m0uQLo
cJJYk6Sce61of5/KT0p3t3F1pMgr8II/6+D2Shsv/dNbuf+nPWjEW1Rr9E4OTItOH5N/3vJjYr6i
hQED4YvRY/8z9OtlKX+0BMOZofPWDhNI1obMaHOgYAnWD5RBF2ZrOUFUDpxbuqYVIJMsd43oIusN
SpPks/kKTAfv1zWFWo5bnHezRyqzilzHMBgRkNWLl3xe2Vma8ZrGgzqJn+Su4Fl/3+WETOdSB2wE
k+j1BQGooUGctyMV4ArW4NlXQgspcE+JVUj4opmDmGidDXxtUATNutXd8bLDE4G9W77HgpR2q5Cp
nd1OSCvYDDMIeisW8PuCGGleI7LoBuO5Pz7QaR2DTew3kkxBC/McxwyF6BL6o5aHyKHHvGr7JtYM
uhcVVUnROYZ6RQieeziFHaGKaeHesSKpSIP6oaz+fw77hmizmWx+fnvBRJ+/FGj7tjPewb35IXmt
9PZjDc1qUTRAU96WXdduqkuF9dLVjPjkIVqrFGfAly+2AAD3nCy8esgHvG6zxUndk5TBMKM5MGDU
+gy7LifYKiHv2ks0hWS8SlkGdt5k9jyd0IGyu/FhGEv0gXqu/jzrDPyeUjV53cxjFSxfNqtiSByL
bJAGpMoJl+rvJefvv8/vuysxLpIRvmGloVkSq2kFZ9Oqegxz2crccJGhksjbfJMuRrBZ77JTPLIs
BtjoXJBHy/GXnH+GY5gONzp+LKmpgGqmYOQTwlQX6br6cS9h0DuydqZlgj7RGsYu4wkXmlZbwq+0
rdetdBgvBXVz3m3tZ8hZ+SMzTL4NyNbjqwAmPgjAgsdXpUD47JJV2YDCdJeOEB+1atOVFo763XxH
IqCeuzhVkzkloIbOZ9NqDuUsEY0xH9bBuU62WcloCCEXXOXNgc6LS50wnqUF4m7GhR2RPq7eME60
PyLZR2z3SC+K7ZR+2uBBhyVrOz9PUGLjfVsxDlS51tnuDA93vKwSoJsG6ZfvkZToGBZhbXqPGITl
gsspDOEX6XF15DVFpzunXGMtrtV8bNCT3SbTf9vFIdF3IG7Uof6NDt1S+w811ySpyHZcbBieY4l9
5+tK6LelZUYoDh+XEtPcwJF/SgIm4tvKOPD+GVkmHP+/bFA+HuF+PRfMzlYPuMidGtLgsHdrVS1n
5f85ACsXxI5ajLPhIAeDmCsqjiv795IC2GkkjA0Aps7EFJssTkfs3hT7v1arvA5O2d3v87vxuxw6
ppgYRgekNKtjbp/vqJW9bdJLVHSaqtq8WVXPQNnfAXcGDzS11QYZ23/Imh+nWSfe9pdAOYcIHIHD
ZD3idtDBA6RgvLY8IzfIvvwNr3VCljSXvB8Mo2sbc9WUAUSLL0gPY2fxYcaxncPcGATvIehMU6Fv
9F7dZI6UpfY0v0nkkzWQDLHaByidLIynmrV/PFoqRsUo50O8nc0ryxlZqHHotnabVM+6TxmCokxz
Bwl5Wzl4GM158ypb3Gp390Ggol88BYr2llPMFEhj99MnxfpWkwRFjnKncCo/k+RaiJKoVPEfA/Ct
1uUAP4vIPXgxRD1xjVj2X+SWkwupVKTu3n2X6dHln5YbuESHXufSCZShcO/f7HWoOzXuHZIAU8zY
mbxhWcovP/c9eEl841KW71S3PRY4ZQl3XB19wxneL9nCugM/o4skQZxF0Prhwc//+TgvxNvMduab
om+Da88XFdEBd0SEVCQkGr3JcJ29KNZO/MwGbxKQwgNhzmpghSTK6gThG2ythPwYC8r6hLeSW6LQ
Afs9TqKox0AhvJkETuo3kjRFDZ7HS8PsTMMpbMprib4Ly26RiohGyKsWKCPbY18qz2eteKIcbHsF
bbLkaJtgTA/Cx/9YWMTwNLhr+PURqotb+q5SA21fOPBDpY/vfMblho6NCUNnOCqyN6azVBz/rubG
L6dvkiuCU6qeFqME2IQGEuolyMEs/Y6HGe1xjjNDVMClETU9lBT12L0XVyIsLLIn5nNRxbB2MHk2
tA20VCgmIlVLTyHP0LaD53R5bLzXNF+GWCiocanTChuy+9wetw1mQluubDCJDN7nNh66UPC16LyL
WUQVxuCJU4nz+5GEuVbrl8Q9CERb5N/M0XS1BuUS0nVNyquDNlnmTfEmirWg6cT42T2im/gNwS2O
xgw65BbWobq1pZx+3RWR95HjwR/6M47Ghf/E2qGckXJgIYU4o8mXhon0kQxw2FEFL4vpAsNChoHP
8XDidq0Yw+EV/EkBYovkHKgFAIOqh7FiXa7gXtMHItxTBeOQXJZNWUvbhnqw5YMQfOeMACFIVeXk
hflRDohy1BROV5+NNiR58+ZGHCsnaNY82U4005fOhaP0dVwYtJf2goNbTH0VsSn03YBLXBKQgvvR
HY4R0k5I8iDPMV9NoJAsODeYprgDqiNfCtV3U7pD5JX9weJTAlIhcvHyp7NrW8s4ci1xka2NV7gt
gyX4OcD/InqamemNJLtlc6PlJhmTGBA6biGqnIjlJ1U8CdrqLQ41PiQhijCB4SsvQSNUa1CSJa2s
o9mNihZkPPO9cffcxSBIdYLMHbXYalHpHzKyWpgVdNn6pofsOXu0JT0FJaF5ZQBUFale+c4MoxcH
PzDWGWg//Tvs5YNS6QzHCUILx/TAKe2tVhU5ZBDIu6HQxYipHu8d1TxBSAQhCUBTN0qXUS5LYdSV
bGbpPOyKrSrADB/oYTOCdjn4geg9NgbGnpqtyKsRSozBScewrCa+B4UIHo8fOamMEJpGu1BDZJ61
RU45HcmyeJXIMQaG4xkNVeAfxnQmvz9nBeW85jJlkMnnFrw/M0jmgJmZqIFM2itAWVOsuOYzSzGX
ghzDPIEIKbomZK+9TAnic3FkgnB6QUZRoPMHiGXh2wkBNpOWOHADrtvJwhKuvcc5zFUuv4oQ+mG5
fBZgvcxO6ZS+FkMPCOt9wOqUUiSvxWUEjOcJm+ITnObmB+fTDSZsSug1Phk4WmSSwvolgFYdG8Bz
ZsPKPYDv88lWinx3j0V3Mm1h3kq+WXiwEd9/YKWhcktImKbt/hOT098sZShZTxuyfjBwt5DbFHOD
UO0CNhkqYUsPmLS0V2C4PPZjXDvXgaUYpY0r6ZRJhUOZNR3Mo1+8U5gasFkkWDeroivLqqgE1v4O
pAo1OzdbQDxmzwNzxdpb/BzRPQNVegXOUEqxHRIPjl/P/Qu99GqVaWNB6q3g4rPpvOJvFN/BqwWm
gQ8cqVBBTiPcezyjq+kauTXZGmLImXLREJE2e25Mw4mgHa/ldyfwdO8ez/IMzB1EPzZOJwrQvuI2
vIDsEVQz15LEo8yrfT3ujR/2iSCmYJwTYSd61mx4CHkK6cW/1SYFRoza4vMQcdazAjwBl0eusM0M
jpH+ZmKTekZFU25EpdAAzaI5Y19V3BKUz7RBludvbw/DObnH1NKMVMFT8KtZbME1MP0IFMUFPx3B
w/wO/T7ysqVgBsgGuWp/fUmB9vNKLafgtE2qir8+eK543q1coEibkvltEtwmsKXqn5vOy36bNQDk
qb12/eeTLrF24jbTjycStK3yntsO9/QyFt5TEVoiuXyN/iCRvbzMzmN/52d79o1nvsouRYMhSZOJ
GRxqsnUiXBYLoFUeBuPHeDNIGTijpOmY1y+KsVlgMxB2rZ6CcDF6hfuZGX5s+XNhFtausBJWsnlh
5mowMzJHlAx5CZECOr/09Tc9ti2fvezIwu3Acw9ZQrM2m0a39mvC6SFOZJaNftgkmtVA62rx+hwM
pod4C6j2uuxhkEDjJ0Q9iFIN8Q7+JWBk+qduPwzVvfqgXFWhZE6mj/7BL1vUFOT0HenJP9OHkFWj
/7PyVgmXN5MihTHpAK1j6pCMwVdCOS8SSLZMcpmRyY0d4//SVjARhARNyb4WOyeGvIhJxUB1DA+3
fOOeAE90O32LQE0SEEdtSLVUU0XYHRmgmBRCYkD4ry8QDSkcikyrGhkecwfvXUrYOae1YHz8FKQz
YI4RE4iYrgBDQqdXv2o96iVM/YL9oxRboYA+fKxZskVjm9JJAG+k+esCzd/V+SKGAiVkXI/tA1HK
c8kgDSkjS67D413Nhs8V2/sQvswZBsn4O3ts5xZpvdsJMI7R78EQqZzRoJU9M94/TnPeVRKc/MhJ
Uj4YjOKIlXozrRvoYXQ0OnixYWqa3Aga0bBj6MTIwMaTuHt9zso791u2/nBUmUulM+FuNqQ5pXin
ic0/MaA6gZ2aJvhXV0sRfKGFehdYozrFnXZXU17fKohiTpvGn9Vo9vd1KwBgH4MkuKPO5h5m8KMC
oI7EUq7wJQGVQ6vxQq3CQaoA3CqiZbgAQZpusalIvwJ2gmEjvvM671pYoJrIPBBkm7oOhGDED2JQ
kEu5WFkeSu6sY6Vd9u+A8WAu+8MjBLWCzwfl3/1vHr/EZLO1UmXSItfHSrMjh2AixhMMn88ajAXN
iJMx2yPqeI8M8myUDCdv3oxP9Y2CjpBiPNX1lKprdWwbGqqJ4JUzjelC+Ed16BZYmmvsh/lRbXrt
UfVbWqIpjc+o6/GanQJzchTCjLj5drhguKjGX+T1FOrvP8XyfoH9g8jgxTW1lFQr6inZi+VRPbT3
LoVyQPsr7x0dLeMuGZWqD1M5/gKQtRfJbIuQNRP/WtsjkG7wlB+sbv5ZTPDA23vqHQXzGOieg+bS
q6Z4M+yiltkoUzJ/DeknLM13bEQDh+zIJ48//Jurn3DlaDu/gSw6lUmOkj+2wbfCefRRTm8wAS5s
sTNyoV+PFy2yeMsdSwFfnJ9PVKiuDyKIahn/twoR2w3SDFOGXOK1Tarkp2EIIJnr+UlLRkzju0dN
klOzLrAHP9CS37r434uSweOyKgsUpycZM769FCDFAf+3u46S3y62rgGe+Oyix27BgihLb3MMxx5j
V32wnK6PsEcUE3HRdKVTGVmtvQOoRvKDjYQNtpJ93Ti/C2Lk5IK1WCHFLTELTdbLGJzHvo34y4H9
kE7Uy0pNJrQSpsOFyMahwtJyVBoaRfHAoNRyYhjYE1VbAX6ryskqqkh0n3WckUtSmLcbGzNZIDNh
bcTronyt63NPUN/vF8EJC82Q7jZyQzqPxyCyqiKgr8IoZ9xrWvbjFpqoA97qvrMZB9jlM7699COC
rYwBtecYinB4IP0iAylkzGmh0b0vo8yBgv+EVzWwcwIzVjT69HRnLwFLxR41VoCvZ/jofgDSP+02
3+/cpqilnRRDsB0fhHU2tF1mpD7hylJyKiyZOJyGRaEZnfwuLKtK2wsgcvBcaHtBc0C4BJqHwhx5
9H9Gan0IvhRJgZncYu9OVcTFKsGf3NRLHCKeCPKSX0pkX+2/Lqyfkrzp1opmlWuYhN1CAWg8DPh4
TJ9jQfJMCyve+fpRMTpU4RLaQp4HYqkCSRJ6TO1TujuTRmxMtIwrjzX1ODKyYxPLgOpVbynl04qV
2bvIChm7nWyoEn9QWXI+KNxuuUeUPnHXuRhWams+VoCOykGsA1Gc6NMaUpERzPx9qGs0o54WaUvU
yEMj25mowwrqXvj0ApGe7Keuk7OzCDpXfbpoSqolVgQ10ExeUeBctbBYlNgkMbXpYa0xtxhkLEwn
GkYeQC2ufRZwjOxWxNlCz27sIuxxSJ41ElqzIMnJ9wYmFclXLd2CH+Kx1LTyx1R0vJ/qHXFL4EoR
TP4Dj7RWlYqYmQoDag2FjxcGLO5AYxrHO8r0dpzQbaJlX3QabXIKLoMb1hV0SxG924ge8XfxqZqw
4dKIGPuze4TTKFPxYpCkuj8sDgH7dLAVufANtX8FNjd7SYKaiFbHsqTvN4UsPs+Dv3aWWrn+z9W0
Zio2T3Ez/CQuBmXZK/6PP2eY3zdlg09cyJXC3nNvfBK/m49J49mD7eapZubrptvh7XUDuBQgt3AM
NYZni55thbFMYTCDIxOT0vxVoNKYRtYK7BU8LvEY/bhVK5TUy8h9vbJFFW887RCbgLmk4fdgqnzS
f2HaOUEmCwjjevMbZnydLVRgfd5H3gSjLhCzQvzaaPypdXCWvvIVpZeHHZ/prhoOVLBB7E56Ebnl
S/pZCR8EYumbznOOXfu2ZQfGNuJz94av/bIJiIYBsPIfFlOVAKJQuqN0D3t4S6srMUmLGhisxwi0
xkj1DHGrJyucwP4az6kjHyMGWFuAbcCaNvnR+QQzNNEvLrDQd+yICJaoJVL1LswblWEwc1EhamvQ
7WrMmGMi+HcIvAkjT3R0Rb4cfNW91yEpj4pS/Fy/qTojYEfJkNvH+9qZwkEXYubmmmOErWP+lpJx
aho1/Q/JmT3nWtMjljTOBQ7NOs+XaYyzGl/T7EOtfZCTZ7LlWOLQba0eSAaYurKy/o3n131qC4Hb
xWf3qzsAg5HmxtQQXTOo5EDzdSZY/MRrTq0K6+vbl4vAcde/IjyoMTEdiTLnbXWtWxYilVeXO/JV
PrL0pXCwWWM/UVH9sCT62tWhA0bj0HisqSWi9ogmiWgcdnGlC4qmHbXPEaXeFuJDNxKoO2uUkb4N
+vE3qfNpHu41ncAvDl3qT7366yq8jo5CFWu/bcZ+mF0/qgKX4U+svNUrImaA5Gne6UYLwnKDCYdp
DM54iZkdt/fbBeNRNnQqe2mFMcpAVZXW91zXH8ICgDnEzcUVRPV5AME/gj4BcOI4bkGP6OPDjkyF
Awl1xN/4t0Xl262mwQIEPGD69kqSTS7UN20sZ7OT59Xk25lR2x3RgZs8G1XP5jrNL51KEslmnLLg
jcGbEvcd4AAC5cVlMfZjM27L9LwrVO8HsYNHhpsajCm+TP50il9GzGtMvIqK0e++rwyt8aywpr8E
bn/jscd9BLYUL6ufDJDTHPCHSDyVHmBAd1h2tLPU5hkI9y76B5WZixTJF8ZPSO8VqNa/iXOBrRS3
XGO51388ntOSzwRqnHLt78efIraD5xWRLDpWdqW3S48uJNoLA6IUa2JBFbTxonxA+zeJoupzDOoS
AzZcKlpKtLh/oyQQHYOGuBLoVE3bzF8ZE8lfxIzDlMb9tEwuiYyXxsPBASpcmdOYmOovQdMjrgk6
IyP/Lx2vdgzzTxwUHuDMn+AefCypLHIMRw4hvfzfpqOw2N/imlr1gOjIKYEO3ofY+S2YioanENZG
mENAFdoEjLG3FnESO7j9EEcULw/OGNb6WuvjI2L4nWVjwE6DoFQ+Vr5joAXThgj4qKCcCVYSipP8
m9YVJWY5E0/QXa/bmXR8325NHkKjOkrWWwtP/rJgREUnS7PrSwvZ1Q7BMoh5221sn5vb+eZcBlc1
LTLiQ1RaKlFIwYF1vNBUgXNzSPK2kjfYMHfQmm8khyUSeWJNKiYYqed3PSEtf8hWNxp3R646JlSa
9AaY+VeF5giXacHzn4otOf6SsqMLdaeLdCSLYXaxvg5W7nAkCPTPzkg2OgX+WmcbiyGH8UkuF6vg
hNHiQrNRqEB8xGUuHr21sWR6EGa9yhtmxifUD/ZdZ8VN1IPzLY7b1/lwEGrt2O02PsJZcmpHhWvQ
T20au3xKmNMI7mRu5rkrni8PmYmftipgXRQFsdBZjFILm+fhUD3D69WgzzX/XaP3ibh2OT+MkxJX
jdsV5//cBZCZZg6+0tMKD1wKnTXl1RrkSzZvmnCEEL8/6RGtJcjyPRG80pqO0/vCFAnQQFtHnHfB
tridFwgnDn575TNO36BRf44QhWaxb73nQwSiKciJ+S4fhM7ZKor2U6nHfRiLC1bkKiPGHQgKbFkK
hRYTw4tk0AJs3R9nTRgQDjQisiGNkV6fydjAunK29RYIbAaKIBX5EeT+YT9HU3/myZf48ps8XIST
ciRSX7mfno1/iBcxua3EWiYbAgH5ZEV4o0N88ExKjQVdD2WI1YJ/UfJ07eBDN3Z9ywhxZy6pJz1V
91ZK03uEZtyBROQLY/GCRpINCbUZKUSuyd4QatJwTOotYAftUonw5QpbapShfbOzCVhFVi0O3HqN
CI6qe+4q7EeO2RxDrEQfi91wQ9xckhYtHv4NwstMxmTFp5IvhFsDdAeDir1puEOzIWKE+FEO7mPM
pYV7/9Q2kwAye5/gOKP/azxGJwOTfiShxtFF3BrN1kEa56QnpJft5pazlJ4DuQmHC2l/81C7z9KY
2O0JPz8CzE/L8MaI5QwN20duDGMKjq/XK/j7Tmh85G3uRM0Sa2YsGtNR2kz0nyhK2jtFi2I/RNVH
YX/DI9Jo+ClijMkgjRKGnxLEkxAOgNWDv6cgySgGdDHIq2GOkqHVxnLmGMQYZ3HxM6Tzllrs7iN8
5uZ45yASEgWu4cF5abJ+celofoU5PP6bqdg78jflEkag4qhNcQTrPevMVN4+CxInpc0LQRG4ZwtT
bff4KZrQy5PwtJmeJHkYPl1gBPNGmfpWSX4LArztCPwutCCxDIwwHsrSm6AJ4tlaA8uylOrASiTM
54E1ZpfTI91kWsRNFbTSGmYeMQl2Pg9yA2QPRZP4vcnZ8TXdp9EUzlmIQ0ZSAs2F7n0mMPT8B5Mb
9BNPquLNDlxO61/R58BNXigRhr79/UqA5S1mXbxqgdKPKC0oucYy85J/4ip1QhW08DNx9ptu5XFc
rvd7vrev4Crwwe3IFkilCC/7YLu+mywLg3+wcFZpChUi7uIxONBBq1czufc6XYzMzT7zWU3oYEzt
//4nPJx020+VCj6EFF3XHdn4eEWVSgCwisIylRN2GGhC10R0L6Q4sSX6OiPFcMeHrA3Z9545D134
iJ8kahf7DyY5TDMTWGUxvNn+1cKtuEHJUNF9lyhlLSbUU+ol//j046aPhujF8CD+xkDDSaKE7ezM
sWui3ZWxO9SXZ3j7WHwX21VICtRzLN/x6Mp5XmmCKA6rvtuY+NQQN6B1Vy0lfXHP3EF71KSrrDK/
mkf1bdtWn11Wd0QkLydL1uV00R/u20WMGvZxz/vb1T2srHx7GTd6Chj+/L0m8MOqn7gWF6X7E3wG
BFvPER8e978qIHV45qo81hAr4kHuAE9snhg3ikCYDcvh+61I2INlochr2iaOes3CSYoYZsoBtGDZ
ZnH7oNOhBTDCZkC3ywSi13enYlvbdEmgQ+/MzG/oigXwXyD2LCNvV8JOxZL/NwDU8eQj9x1aZGj0
2osuUtPhv2wkiCE+sH+NkwT2LZm30i1uh7Sl7bW0jhT8/03SH3qJrvyQGsTKAOHCKVBoLTykrEn2
z7/LO9MApfjymUdAyHgRPjK5wnBS/3h87VdjMBKCCEW7lcilYqTfUt3IiKgN/CUE2Tljyb3OgNYX
h8tKmVh1uUN6sfRmvrDFUh6NxMTplRJ49c9uolHVTCxKbj2kF5rWe0fyDnVtvSZs065JYUa2ZlJX
AplBKczjv+i6VndCvFktyD8PfxKkk1AB2iFOJ7iljvtLwd5HeO6J2VKdCi9qy9jV9Q7388SP11nC
TwKs5PmmsrkRDy0c/FZYG9Ppcd/azsWLDMY4wg0r72Og0Xnhdet707gm/VyO8mIT8Z78QbIMwsUv
K8uhsqHHHWeXBEcXIB5JJQ7NkBk3PkJpsjo6u/O2J0w9kOG7sbRYx2Hqy1KCI+rmp4h5iv8z09Of
y/nVqDHO95buZeXQKIwb9mpG16pVPyFq7gZVNyIO80/mhgeIAvI1rXFJv58MjzlEWG8d28oOMHCu
riGTlhoX8pwXXKUm5TYpp0+/dD5jToT2CJbY37P6vsF6a+7iFayoLy/zw6XIkiXVLF4PM69Ec21W
v1pcsARg9kA9FhdI8QXj+zfvX+pz9xLykutFj/HJP5uYrQK/qd/POfUsQWi7TSvARduKQvWLRJOs
ljIoBElguifC/jlwAtYf6S1Bwj0d9FkmZfc6sWCGQ2I6N3znVCars+ngYnrT8XajM9hXhkTaI27j
8pXsFrZk9JZ94qU6UWKyHZ9ktb0P1OskjpVailCKLJGnDQ4bqSw80/P0Dbma3QEYgQwq7JQ+rU4S
VAzXojxdQa6RusUHsPIJwd+OJZkUaa3jpW+85XnwWQ1yIhJPzg0wcxNFfbK0Q/IHfZNuqSJmkr4m
auyY5NKMvw5hbd65Ru3jjbReqODUErm5QfEz4DgYIYOrPBgM1Dqs8FYDq4rB4GWk1KDW8FhKugu0
CG8KdLpbjecE9M1FQUZBhz7Yvgd2AH/qDf0eh0Hi0o/1jVGp58uAVjYhGrdSUrKyeTj0SGcwqWG/
fKC0Nmtrug+pBfQnIU3x/qslXAgQbL2fxNYyFRDjJPpLOt3Is4057pckEMQm9l8EyZeRe5lw0m/u
0d+p40SQtWhYtJg95IcVVv3QIk9cxJFFCLvx3ZC3vJPUGYfkwFktqE3x/DftU/nRo4/KnehqDQxJ
f9sVoX4z0NtC5A1Fvd82Ln59GO+ufQagEuPo5kNXTGfG8GEn/2Hd5oqcGnAbbTQ3OaZ25y3NLMsS
VSVQu3Hh4pZtg0h+h2krS8tUCzp/QFC8ZhhzkrCOw1vK81cKN+xFve/cppcku5qMkgPot1+sB8IY
14S/rtKJFJzOSD1EC/tcGjRL2QoG0P3ZqzR1hM9L+96I0rprqVrPORHTmqfWs9UjviqMaTDV8mtV
w5kgd6yh4khVVa6j/A88fPQpTyf/blPAp0m5/OIKszWL5Y6HF7BBvfy/IyCLSd3eyPuOEOjD1TL1
DC32VTPdY8dBo0NcwTK9qSGuJzEt4VhnPHu2mZtnIVe9326T4pWDULhbJvzBLoAr16jYr3TkMypp
Pe9xDlDujqoaM2EpuuSvkGFwvmcaqhcN+Ky8s2Kw9sHDKUP6lazP57XP0zl5csr567wJwJKB9iUS
APT2cBhQpboseoiNVcHdP2h9mG5+od0SSMjX7z6fM+pB5Z7yvrEEaHzhHUhixtwjtArK3WbFZBqu
bzhucPQNpsQoE2JT6KnEGwHC5xdQwPey56muBRSJvZ3gtTKdNQgE6KCtkc7LRbhcMbHpAPJf55v9
WXlfCm/JfB7oYCl49HtIXTMTEh6smX3gEvuLkO2V/R91JqBiT05nFNUQU3rN+sLjDgBio2n8Tq4h
yDS5DFHVt+7eeEgFIaVbSeVHSwyuWtrmZb3VB4L1T0tesSzCOP8tyy5cl68L5pN8maO7afU9y92t
rNJBZ36NqrTxDJ9Z4bEla/SwYUQlbhUX3YA3gTD0oTWf0K5SOt36FULz6NXUxbK14/fteRMbFX2n
+UcWhj55j/FSE3v/N9JQ4rEMa4m1UzpUxeHkVfjcYoHUAE3Gut3tqNNq9a6CNQ15PlkZdmn8T1Sq
zuEeD2KTY48EKWVrgwYZj51I1hlQ4GEdIBw2dVrDwgctIQwUpe1yPVFiW+9EgvevfqvzOkwl7eiD
ADjIUDUZplTwr0JDkZi0pxK8aV89rfCHV/D9CubsBQ8DtkxTyYzyz+votgB9S5kjnqEtd5mt9JmZ
kfKPPrS/YMyp0YaQF9YpxRkDKvAYPjeseaOSTbtsdS2HRbNf4dSjJE1KEYiLe5NdLGyZwAbc+GUh
BAVvMQ9gbokdPJzUMNKe1/54e6RTLAjsWiqv3245hdUe2JQl68m1+l1YEakkkx9osQAdzRIUhaCx
UqAMA/D/yqun0JhMhWWveFQk4fQ+9gBYP9bg0ls+/NcKNvXNTArrGM0oYeiebPORlzGp8TOERskx
cd16LA+eOgPXlttFOen3+TVaimIhYXx7stAGJX3u1tyq1GKJLIMqftUx8vt6dtgmq1/470sQ2h6m
AxlfGpgt3krP1G9h5fDxFQIAaSpbU8y2JMLapQB7teOX/00ndHhj+meGB/msRqqs3/W148GVVXGj
prxTE0Mlp7jmOOxHcJIaADoUfq0LM7s/EjAqn6v9cu52B5CaNTue64vugoBv7wBtDjGgodq3yK1U
VWdtk37jMZq0x5+kVw5CeCqNZV+8hu+/slBw8rS/gehbt0bQXOp5HxEcjtAqHSrEJjm/fAr01aLR
mvvvpj6RqOuzm9102jRJDF184U5c5ARnltF9IAeHptyxKfYarDuO5Hz5x6Emd8cJdSgA+Q/H2SFt
aV5RatgbJ9HY98rws70VpjnwWdi7G6Q08/M4+TITd2XBXrW5DaPLPJumAaUgIOXm69eTAht0IzF8
6u97lJzHtSBUMO88Z06zvDd0duqQWHO8D6gPoGbecNi/gIRmAGnyGY1cUYrDV4v2N4B6ZhZUMrqk
KA7OmAnKuFM+7wCIirzrF2v7TN/TZES3E7UYsNxnGgsCBqW2QPAiSfuPRvSFgcI/NGuUojiQLMVf
vmE9PU/pAcPiyfAOesvqh1rQkSLP8d880Suk85WsO5kA89WaWUUValFlCAe6if0aqCGYbSHDevSy
Vw9ZSE/SsaNlwU19Z+DsxVhBRYklPNIjkbLHbKPYyjZGDnjgN/guFBqzICxarSfp6fIsONTL3tQR
G8n3mcOtqT9+0VxttcL8H7VudQq8g3e9goG7Q/i1M0x64MrqJmwxl1Og3E/UwLeZzfyWwlln85xl
cvRZ1U4EDeQet7UEPccyesgBttFaKRLcd8RvOI4nVpoPcVO+VoozeWp4SMiY7Adw2a7sAN+sUUSE
X0b9c2Pj1n8Vy5lL9XIebUnfflXaUF+ccg7YFUwahnX0nfLW8Rapp37mGrkOSkvQ1FcvaW3mhBrA
dTStUZs6tR5LkEdZeui6C8JKeECpO0Rw5TBxmY9LFw3PfgIFRC1fFA9F7OBfGd/89aSmJ6Sg5K9H
kksPW2+2NOt7svVaxXsfYOZAt9AMEbHlMoVZdOBbFCA9ZnOONaAyHHyIxBzxTjaZEWtC3b0uewKB
kZzyhknRDGXQU6B8hip4SNHoXeLKFXc5nSW9pEZuALpnUZlXiSxTdua3RqXpqQlYDOOwEI5uSMRJ
E/XrJiQmtB9ZOh7egHMuXeCXN5C8mtUn/G/9zVZK1P77l7KMk5HEfrLrbHWWwODlIr5UdYL7LdQ+
AYjquqaJrTNFCzVvaCidIjmWLckkPOmPB3tDj9fNf22fI+3WkKVxNdRNQ2SafRQJS8vShBB90ZjU
GeWPiGLnqweJwzQORTpRpdpkJfM5T8NcmibVJLnRNplabcYw6zFZQW9NjYbZNCTSmb7FTW+KcyJh
Hgm1mPcKeg7nUzP7hwWnyoB0icbHTRZuzd6tf0/RWbiCTl7q7yN5UHIIcKn0UbKbwNG3HbvznBS6
bDyVW3fCY/n1yoBrzPuf3IldB+q9dGEoh04NIjzaZihvzResa8tuNvTGd+Ozz/SaIKF/EiwNLJay
58fhyVzEzEzghZqT8TDr5ic4f5agC66RFX5fw2149RsphtUIULICUOtNM/Lqfkqs9zeZ9TobR5Tn
M6FPfXSNa2U4YIvYYmwA9hPu0Ue9f2bbaLHF62pEmyDNyrfJ4xwmASyq+PErlclCOYBC/ycKpM0H
WBLn6iEOEeVfNFIlVC1DRoFMDjq380fK6b6AP0Sl7eEiNSfSDZb1fC6eKqY8zXwzF695hXF325pi
xboouPdyc++8wm+cQHAtMRVYTR9c5ZiGhQXJ3NDN+d0udMIWK9Qs/j1gm7mQoxVCaMZYE6MqYZcp
50Pmueud155ywbzpQqXbbTxP4b0j8g1Zwj2Td3R49p7/m+QrVxoHyx6pyzMmrSOimObyfRgfJKI3
L2OOkd6mEQmHuW3Sx3PfEXCrK4k3IQSiK4SkLNhomIo+I4r+U9cf2mNSCNxhoVBKdtx55cV2wnaP
3oqfPGuGEubn2FbR5Uqa4sfRm2AJ5KciyX8a6JIVZqCPVCcqoiV3mbg3yGHN44jfBKUU2eoNiJX9
a0GVMQ+C26JTZLDlZ4ayC7okraAazIaH0ajc2nAl5btJP+6lDohlESjxo0V+4NN7oh1uVypR0t1s
DjhcjxsA30ZrZ8mesj5PHpSR4/ZEB1/hHbBw8DifQ1F8h5cfigz5ru3hkjpw/ZJWecJsUkGQXKpU
34VtlxhUfsbUFv3rPvENd3WmbQyHqLoOoAf09pnu2lA3QeVO741Y5Y8jIzJ416PQezLxZ4Yd+Ewd
SzwqjPCgecHkfGsRVccXApCGcCC4ioasuswxcu+6edM8kvuZLGwGMVyrQ15kpojdHWcjTJYsZHM9
MR3NIdYfMLxxdJ1Yme5nUcnobGuaWssGiM94DAcPzE7HIQsjdxFg8t+5LQl8q3WLKqmxTSpZFvyR
Z9JtZma+UtjEyBr0ydun4GcDRa/YgSLL7y2t/7nwZHhH4sDHKZd/O+x0h2hLCSSrza4h+6QOk5PK
QsEIb3BG/ScAaokRAtF9m9RoLl9HM3r9en35PMosb9jHV9GjM7hYbykLoC0LRZfsY2iIDEv4ZHja
ClV3OH/WrWav3TSyv3WQx0Zx5ItGsN4651VjP+KWkNqZBwReGYv/FOoGK+i1B6DdPP3fQO/aXRXv
e86z0+RwdOgW9Kd3/RJ1YaOq/6rmQhIa4gZ5Fw8elK5jUGaB6BaXYQ3PnLmd1a/wwNNREdamvWaU
r/E6VmUSofX6/a6kbgd2ch2w/XhEkUnhZLS69O8cHYNcDYPO+cj8POl0Q037LesqlSocpC/8lMmS
quFt2HQbunxL7iCcBmv8P3ZKY7WistHuNxCzOW9G0ic07HCYw8jm2W+79lfjqezt5evCZ97hvpM7
mXr7rp17YOAWxnodmOwRhJM6Svcu1857tYEUbBuBDgo6nj2LT9PqEruJw2uPvsoWgOXMRMpsW9ny
Qn22RC9Y/AL0Rf387PPehFzDWLhMx1d67TWaC7MFyjePFIRy8HfNSoxLsV73sYSOGolRd1Yo44M6
wP4ygI0QdS6L4ndDtxR4ep9XPdzJSplX0FzSbAlLxbhzwRx1HciP6d4w1gfALMmxvbdsho/pzMRH
0WpsSs2Y4RweFl2rFs7snHy/LeECfynhxPdLxqUmXbBSs5Z6aisXRGp93jwWgtv4O1KeXMB4McFW
oxR650AZcN/xr7K5mPVectDJzhewTR73M3U/v92KOEkgusFeyOg/DBMTA15wBuh5LeuBmn1a0kQs
HCFCVQGIfPvNkX/DhzUNUdMfSo5tYEYORhxbOXetsdiyaafZNHE0OfuKeNf22qLW6XDRy8AGQZi+
70CqcD3Hy1SqDPqOw+8SRGzSRiIDT9Bh+uWf4YtppI4A2xsBRDUfKvy/HqyjJ5uKt9zHMG+mawy8
no+LoPj45vc/LkhVbiKEYPIaBkgylDDGXPP5u0QFFWS8e/0jZfIq73s8e9ww3nEg4FZa83MoCgA+
8STPAa+yFgsGQHlwTG+wnsISlwDzqzVuQ9iENXGUhZXHS8uGdUmPxaydx+AOdqgCwRwtJx4t6ydR
Sgg7Q316m8V45N4V4ddg3S3JpZzGWJGUX//Qqd7lC985IIrRXMVVMhoMlijdOVo8iuzzJwVEnZnH
qNDAANreDzhCbeZGBdxXaRyrINIrfUzF5VUQ80t8N4UkyzIznX5EDl+P5UtEdQHYpUG89ovir6Kv
lrbN/cPNsUK7wbhgdVGT+ppaouYeOLQnqxquUdzVKMyK+WUl0DB7io0t3GmYd+I4AYJBx3Hn6T1Y
E7VUL40bCnLmbd48caaq8v8QcmECG4xYrWw13jnipMGXipHhi0dX/AeQG2f+N0aFQ/WEkW1Lori0
sD/E25xhl4AHO3k1vcetO6Fd3akFYActOmJSa89U6iC7qShIbzHUUaAnN842PdhVA4tOEmbkNvCZ
PevhcbwOqc8sULsLSoM6S25LkkvBf/2B+KfVId6ghEeivjsF1Q/S9GDBlB26VAGW3049ThOYDv4p
pM09cqJ+MGb2xIND+iVbcvKeQTVJ3WjcWEF/Qro2KWF8eAZ1WuNnwVPO3q3kpjU/pmAyTDDsXZRZ
Ly8PkVDlvxPCYY5oGGsxmCPMPj18ldHXHYd/B/Nev/bHfvu4DS6basyGSuEaQmsN2m9R+hOyu+j5
Q60ErLw+GOlnFfLoMHIwxmn/Pa7aG2iHPNF07zpZMjeLVS+plfIYnPPGEEDbsrF1EdX4BjV4jSH0
7uDqyUXVRGm4jO4tmb0WHWLVEjLQJ8xo7Nrcl0vWNTaE4VQi4r9fieI0MTlM0JjC1iU4eFDPzYRX
OV8ispPtoHBcYjWIkkfHWWSGJl70I0HwxB7F6CuHll6jjTugcMm2itM1YB+MUBzEkR/Z1rIixoQi
sIsisoPWa1JXKTUrGBaPwuN7CYDEnfZn0B9nNrdPaLKcbOd6DFRYT9K/CDrlQSwG9JK7qKg37+Et
CjjqoYlBgAovL0bwpvMBbO7mR33UsmDjNfbmk1oK2fqDW5xXiVIWKcXZHND3AT5HCeSiIpbXkmT2
Rtf+OlBOGy5eaHDrmndbw33lLzvhaItLdG0mZdTFKSoe/Mjd5AauHKjv3edlPiXYaRvZsLNoKH3R
7K4/zftfGKwbGuIn5PvA+maFESuMtcUbUIPABy1yomJ/o2BqnRaHsT1vWYqwPTNahQ+9OZcIPprC
HUuyu6AZYTQSGPsrSQ69p+Fhb33O+kFgy50x9O2+OnDBd025UhzAHiyKWgaz6PTICizPVOe4fw6q
wtISOolMq8JwRdUcdVfl69IQbw+XgAHVAUeW7fD6vpAdjQXtidw/oAmeqtglSMhrdzVNoNb6iG56
UT3EL1jKCTrnmH7Yw5AZ6LdZ7S7xJ70jU0KBIPr8CrSNxxHBmi6PzYn7cM/cyUzVSpQYJTa+lHex
sp9GXEG7lIFzQneWsc70eogdRkQf+xq67J5AZAklgOe4rLSUeXqH6+JjtBE/QpWAu8tDlGxBMEHy
mYzk8qaFvsIE6GWggPI9v/RqvRtmrjfHbeRcxoy0+cx2zvlQ0cqkN/QeHJjn0oFCgHQweQCMPL07
SA7WTh8yssMSTwxJ2AD91Nuc6Slb73lFiG1Wlm6Wv5lBErZWvU+9mRQY5ptoSU7tsxLk0ZHYAEjI
zLi83kR7+hHswz/FRzhK3ZvMGI9KgbxE7RvaGbTToYN4tLJtN8UKHhSMvmWe3cNsZ6x6ThL5Y6cP
0Gx1MP605xDDvIHaVqfU+xKEY1Ycvrd803GqxL0xs/1XXTuKKUtQoImDDWX66QEiF4m2Ls78GoBd
yPQr9a8X5xV2bAlteTs1RPMn+wDhYcGBr2WpRIb9fbdlt0hqhSU6YSN2zU7MzuC2itiktX+vL7Ya
KhGbPhRGyWyn/N9lcZVYavJp8qxP5k53G4Cch4DADTWIMsxf869PaiwAo3pD/DJjsdwfOR65BFkD
1wmW5DV1jFn1eg3hxtfZqSmNC/7LmSR8yLKRksW4XQkgE9de+xUUix+xkxODh/I8elMb9aI1wVUu
SV9hDC6vdMzNDwMMTOOiweehBD9yLvX9Ff7RnbndcOHGAxj8Hctgi9sR4VmacMAfeY+7ouejcHNW
3DiyMDLdPCa0Dgz4z/ZTtcNJqlTomO/4hhjdArZ+KuT3B23+A3PDXNAafT7NXKEcGzg6yZjTkqWW
jyMQ0XAouXbqrvJ37OJtc3YFXJEn2sKJs1WA+zcb11POBFdppvcG0YE5DOIbQxsioFiQ4INCgx2Q
4PJdskCD+TSbQN/pOzTtyrtBgbCvzpHcIxvO68MY2oONX5ZAld0b5FRhDV+8BIrJsasscwf31vfj
CmlPLpb5R4cHTZZ5U6PXOiAeBwvgmF28yVFaYWPhtv6gjKj5/Vhvn9T6YXcFa6jIWXZvd4RD+Y4X
G9sDAHqbrCVjCtrHCU/rgrNJpRH5Vx2a7Qj3vEOYIldnY1g/TkjDU3yXCxAgbqPIFHbI63yfpLCX
bgBgDkzN21gwS1fLYBIEB0x5JMtMeBIBDe9k1tTPewrZRKA13i3biXIpPDRBGOhJp9vf2ChI3FOo
1+5AQKzzRrZ/1IpJrve3eEb/LbvUvbvfJh0AGDWPy/TqJhOsxHABgqBBSwJK8S/fOpjg+BuGzoIh
BatdwT/g8DKLWMXZkVcGyK2guT+nB4ZlOZIeK7Z6HHECmNGXLy++v0jVqSVmkKhlSLYXfDlRQtqY
DJqeFbkD2RuOKgNNfKa/3BpmGHu34bvgyCi6CHXYC9pfRYpk+BVAONzya3nTRvZHNEPQivgGi1GY
SACFCYGhY7y2CaienV+G4Wa2UBy82FHdgwA+YH9aR+B+gUtutZA3puoGPb/gxlfYLKPQC1kv/13c
GSKiJ1j2W/A/HF2EBCKWrxpCbcL71328ltJjSQfKSXdoN66qnzNoMyCt5al29adUWHtI7xJTjYeV
Vj+uGwsArQrUL2gZwo71V6Z+Eb9vVLjqGmpv9/vWCQjU0jweMrej7Z7dUyrRcuIM/5SYJYpXg9m/
OE5sfbz5R5Ulreq80taqgAcK6DgPSdy54xyuiCFhi9YIm3mDcoop7gZrGMWPXN7ER+W6zU8Gax85
YS1CfgLX985Irhhiol1EdfUbVHSPoyG8F/z33R5gOZhqXGuj6DOpy4/sDy+hbyFJBJnFo+fzO067
K5f7er9ecBvP+4rr5d4MA1AmGJo/wLTijK6cKzYC1OsbXJ/H3MNwZqkPD4QNYelzdGeFL5oszfDA
yibL44AmRnt248h0O1/KgrjaO9p8dGADU6YKrUEdTE7YtpBkfN4Yo14l1qmJ49EK+u5+oucyGEvv
Mzv3q1i/5wifdWPsQSoiImLw6+B2Mv+SFYwjXmBmpNHtCi2k9oGbjSf2V99hVRN2gZLU/8PeozoE
oAhtbWW4JrOauDK7pa/LHWvSTjeNxdQXvLumYQKen9NGggmqAR+bWtYXyADdfRw2U8XPSChJIx/z
BvCgb2TdUZVJCAUhRK116LtHcgKJhc7sh4Rudvq/EolWaqq1AxeO3l2VAvPV85lPLxlQ4vNorn5t
0u/OZ0VIXXbSmx8jX4jZFscLVLJCZEoSD7qstOL+u+aYIlf/vqw6dyK1bRqZ9oLCc9SjfvsAiKBk
UNCj5WXrzNqWMOjky4rgAoz2MYP9G7sJl0eUTVEptqfNQxf/L9GxtRoP1bZlKh75iSweq0zJ2qJJ
lfJrL7ZpxSollyUMYMTyskKtkDhFWtJkfbOJZ7YllKo2vprWSoMjz+a7G3VI1bPlC3N1AFiRjggr
QIsq9w6dLPPe8NFiZ0x+as4gDk5UXxpcG98j10FloGoOnc0LL7TQP/a3jq4iyE0M0L+LWoI25t4H
W9sxiIepTvhd+CwL8rgQtZJ0MfRRX6tde2Jaq4qLgHc3EIc5S1DAw4rpGDDl/2fXCruAANnVhkPK
i3sPx7Tt54hmIYIcdsorPjHAtZlE1Zr0At4WDosu3CCayf2qRiaCZilLMLNinCGiYNBXvZ5HGJiC
bnbd2+L3Jt3LwUxSEyRE7UqgshPj/PaQGU11TUDgooWbRXyeVnOk4Cl9O0BrOG694qv3GQCsNOR6
AVHG/ip18jKcpYcbiH5Gi6t5mAgpuReivDQUjd9JgtLcr3ByDFmWQyR/Jri9nj1DFKrefOiQ59KX
6jMj0/Wo8APiE/9Bhru5r5k3W5wNIi20kiTqPCgEAF7cJ81dTU8k84i75s9QruidT6m0nx/psgZh
cxC/VRvdeUHX048kaxSfQYeUQUsl39m5epIW8KFDBSIRBcJRryomMoXE2D961XXkhvFJKM9uO+3w
JHgUwl/AScrIdHswYb+Blwx83T17frzUMAuqolDGOM6rlrXb6qg7CGxB7QUV0Z0VyRT9UwdbeKFx
qIWccumyoEdHbgGFRClkRCBFirL6cKbYTziZF/sVVXLHVhQ4SRRGxY9QsN6C2+xVwUysVvOKmETj
L9R9cM9g34OX/5TCCJo2UfeKcwTPdsWx5g5vWcX3/TdtYHzqic0rkatLxi9L+m1tVCE2XEfnUpix
QRlpDdfYtb0uutVy/Wpq59hVOHHvEpH0WaFPJAOJP/7kjXQOrjmUqOmy0xK2YE3oIopVIOpbTYsO
XafYlys0rTtnZzITvdDkDbClFG0onBFGRIE3K7fix3IS5IKeJgF3FDgVke3tD2aMPEnQcN2hTDQb
QXb5SKoC5nWYW2E6flpxCp81gX75g6EOBgZ55sFEy7mIns9b6Syj5n5nBBgdRf7UD07ZZWwTUorq
jBt6eejjXXQGGlkL08GybwktwEvUIQGCpk+vnzK6jYAYcTE/+r7xSpMQDYkcHipaMUAxUQFT35ei
jSaXiA5Ok+LbJZMoxpkQ1pUGDn5ormiaMLbid0dLDTJjfNTLejK/x3vu9QfuCQgAZKMioyDALIh3
bRTQtwJzB4QQoYPIdc/GHIqufKmhxVYvsw3KP7q2P/jH+JFHKJIxRdEhDnC5VXRd0SA6ang948hs
zdMRzbNw4+UDaEuOwIcL5nA/Tv1HNVQEGszbGlZjMP7+OS6dLux6MxXTTLVSnqVu/RLofn5lplnn
Zo7E7ZvHhs2VMb1bb1ezFfpBo0wqX6StAuKFLDddx6QYSBiCIHQutaQC0EOB8XOMDWJzuFUUrbQc
CCC74gGmcWKAblIADKww/8FF78GNz4BIJETMEhaBN/7TtB2OMk/P8BD5vCY/xnb/rk0vIDpOLcgR
ckKV3z7XSR81tKHIieFZOpnwy4JPmIaWyThWzxXWAr8ILqISBHDald+tyViGHnW5maWPSQ2p2Avx
wn09hrykP8t9eK/spJkPIc+IEgKFOSiI+rvjP7+K9tmsGdStdGtCutv4cHU6BRiK0K4aaHljRNTK
jiF6p3ZAl8kWhQCtxsnTX1tfeGqkpjlnti8jnFZb7zIUmSVmuIP6GK7yIctG+k0Qr/ooCo2l2Myj
3GqjR9dn84QHkmmJE0NGtW3a9S7rm7os82Q3ly2x0OYQprKwo8oNq3rMz4ZqmxsUswIBQ/alHPWS
UVvD1xYLMqo7aiQoI3PFYUCv2p6JQtPqZLNn4Z6DJT+2ePWi5qPIYIa+/fE4J5WqmG0nime2Ih/f
7Xjt3HNKS71bSn1rvKXB81cavua7SrgSBi5HFspCCm2R1+GQXxxQ/jmu69S4WSfI+Cc7fmEvS9c2
H0m7O1qd0f3DIRmbqvd7tmpeSwgxw4WRBEIbs1DXiW/3/gQKTP8fyWNbHoCkE6JR15QIY0Kt3LIQ
6bSgmf9LYY3RRQKz9nvOFW2WxdiyhmVK4DbWMqpxLoiOLVe5Ee8N2lMJPVvPkGrslx/NQglLNLtp
3UVyGAm8It3Yys7JYW5cLUGnUEkcHe1h3YwkFuP0v2ti6XL6SJcJBnEi6V9TUEicMjnBPpIH8UFC
TYb6DAoWA5eb2bwy6YQm9b+EqLEgOJvKqORbgfcX16vfdiWHxTZHOQhCW9obWadaxrKZJNc9bq81
P/eK1lfKPLp4SetkrrXPEMQF6nBoilI2wNE11fIfwPA6NT5gF9JbgnSpbgjpEjNET5RiefF9TJmC
A99brkUyMUJvU2HS3z9Sub3cfMmOyP7i5B3IcUPbQM9MEep6fq7EOC/5Rf0f1XF7l+WCr0OqUAcd
sT0cJX0k9p4u9CzU8/xWPAZF0flQmtDPxPaC9imRe6sFEa1qQkRRE+RG0QWMzCxaLwkn7OKMc3px
PZDWrLeZY64iCnwWM6x0rCCsEGT3actPUSTnEC0/b1yuFx3IbMSqDD9U8ImzTI7Uh+2UOjtHcq9E
tAN4Mi/AZ7T7P+kKBIwMyqo6ot+LrYRNHCiVdwI4z3rPsXtx09lwfsI+dntEeFV6BFFl2tHoXNv6
aYUyJix4japN11is0TWQzzvtya06KCfmm77lgMOWMUyoPZf9HGTptTUesZ9dtdqonKZCcWY+eOpK
Z2+z248+QyBEymTyoOnvJgmIteS4FWqcmNtQTniFXD6BZ89jhd2p93hQ80JjtW/N1ID8/k8lnzB7
z9ohmmsJkRXrrleVLZUIpqYcJarad2XPTEUG4x0F+dmM84bdlzjq8lgjqNfDI4e4ffLOdk5fV3wO
sl54R9cgbgbHa7i7UJqre6QOpSu3L/beEQ8erFnft4xtIe6VDqeYhxY+4atnz8y9V1jUyq8PwT9Y
NGUSacu6yuWnu++RxqthkppVL7xeKN/MS94VGnwGyliNzbFDnmt26rM0y9Q4/fqOrjwY6dlGGKbB
9gc9m7AkNeE2x8y8BHZKVSXY3rqKe5nUECdrbGel0CKC8mVdVUaRjLrHkEzzkBzqbYLeu8KVgN8t
R2Nj0G+cCF/KbbA5rgHQdFKg97HyWaEWp7MJJSJYbyVbP/AAjdbBMRjQYdvajXZzm1SR84hk8S98
11LpsvtZukMp+ICLKrD13LZMCZLkfiBoeRjvokedfDVrbV7HC31GV/UUWUbCaYl/n4LPnA2qVAe8
8U4Df3ptYO9MkpogkK9iLkcTo9ijPj3UISDBfXsbEDebVDMxSGmXTh3BvbBF4RFFPWW7zi3pzuZO
4CpeRTgDh7c706o7enDQfeUf3q85arVdXpLy+ei9DiIogFaZf0/btTWA7OMsGegWCdJ90CSEDeBt
jQpTerFi9A+XzNqH2YiPU0Yikv/qKCXP34fJPii+r174AtKsxhGrJC6fbWn0Ufc+HsbczGNMLyyH
M8eqSNqwiOI12tBUK0DNJQ/gxz4B6Zb3+cbkTjPylXbNsv7XFh9gf1+2LVWkQY3+aV7rJNC8A9Nr
SDqxPB2ZILaX3f3JO3IZFJ4T3hxrz3WwP096JXESpqheesp8UsU44NeFVBuKqIgd/Jre4ZV7hUJI
mgyApSvs13WUvn7WMS3KUqPfmKRJ4ho9zJ/Oy1gccbozLV2VG3MkNWSC7PKOzojZLJHVlAWlgfPe
wBQsSeJ09M2T02LXkZgqWhSNeSrYS5ZmFiCUgYYGSpr5KLDUvRm1Q/wpJYb6x5TBj4r66qRtLWvv
iw1x6dwfBxMTdiT6FQGP0e20mXaqbpiM2orKUq/Kc0bqSyBMVqT44z2vTi8y4nVnj46tgeld2EMt
2b131xlopGGSbh4NFz8vFwNgexIctcapKA3jZIKYFeHA0mOoItz4u1wcH5WQo0DVb9lEpeAAljNE
VzIbU5HnRbbB/RxCuhw/HxQHjDlInM2wbIXlYqtSty3yHImaz7ROYs7PodAsgDuADQU/Jw9FUPi/
YJbFyqrLoxTUiNsF0w7lYrUbhqoO++XB3Aqs+vZpJ+5P3W6uKowiqp3pqdSGzAhIo1qqkcu7D455
GEQaxqR8/xSn3KySYxY6yWTG5e87vZ4YQuXp4juDCKfbp4ElLA38klEaQ1MZh/17gGX8zquudzpR
/iGvya/owd7d2U00hNFX8wbKAF5g3mOjBQ2CbGndAtDY0FaJcC48s5Cd8BYuXDZt0YozbQ9PoALU
h3s4Y5emWR/6WIkCwb1yN0XgXo3lxzDNAXQsrMHoRNo+hBO5yMw1YgUCwdxP2VSj2f0Ibuh/w0La
HY1sleQTu1ivl8FwVEPmT4XNIZ3yAFKR0B6fAEiFqNVDRKsnb/DSwVj7gUZjD1GwyiQnLV28OTIh
37xRiMRbd/T+G9WbuL9q/DE3a2k0lRUNoBhdVHg34Hba4Ca0hzrq9scVTEqH0f41wjgr7GCHEpPq
4cNZTjWFtx9jxyy1rk+7Ckn2GWXsR7ZPnwvyaPZh0V/yrAEYUeOXhCY4xCpw42nG9eMSFcjDUYYX
ggnGdZOXukLCp4vwWISJHXDwNLMPwGwbQFt3EBiKhCbgTx/47wPLv1vBrkSDZOQcxRI9yyXuBIuC
BAETJRqBkqF+7cn6FMUh//Zl1jQHf1ICRpeD+ZjLR9we8om8rmEp6eNhoT1vmCeYjyG5pB5pExnl
WOLb2fL7P4fjxO1TEJUg97Ou026v7EU47p6djVaguYQZchKssgH7wrTdhiH4RCuasS23eDudDrBm
p3qb/lzVwOLzQTTrf9JXg0USvHr9gMFQodiCsNEtSnzVNUL66hlNBjSKqK5ZPkqUPnRo7GgZ2dnf
vqGLrBL/uxe2264DSo4nI1ANeFfOLtjvJV+PlOTCOZNECxGM9ptNpUGOPOjVbUg3aXLlfF18B9Np
QGXVBTjLzZXFIAVUadHsTqsJFmMAxr8NJUbwK01kHjepG6WeSDeFdAlpyPXWr7f0iFqgwilBOuxH
pJ9Ob7Kil2zGlY237TEorQZG5C9oyyJATivdsnD5ivgTU6K3waDO8WY4nq54+oPGlAJVZLOYTq4R
b2I8hv/Vu1ZAtAHttulbf+TnrevVbg//lYiQaiFk0SI3GgQogTAZvQRvuZgp2x7bW69EdObQ4ZiE
+va1LZVpFqkiSqkqQ5U2rzED5tVCMq+HtlIu8PywsW4bbhzhMd1PAGVSaG0Qrv5nOXgvufaDEXyK
1EIeTXyKjV4TXm9ZMm/JH7NVh7TUSpEHcKYBoI903w1tIK6svxfz0LXY9RC1u0MMMC8Y3RM9K8nL
ArYocL/mHKLFzXfeZG2zA/oNGypZz4glPND1LgpX2ge/pFYhMVPLs91uGESCmOHxzsbZG2CIZ0jE
+psvfPCC55idqvQLfk2bWW+1fjvAhFwcmyq6KTwrqgBDE9mh4j8pfXvmetzkeTaGXThceNk+gW7X
0a3o0M5TJHJu3NqTBkq5KP9Obp2wYLXbeFeCgxVpXd5ZPY4X+g1XZqtMNf3iG9KvQHWiMYb1Av4I
CUbDfzgAfDqlKTdvoRRW8rK8D0PFWL4Bj2xHIC9lPlX5mjrzENkwZyOydocWCk3kWfqrMk4+F3ay
M59/Hd/xoK9BS+WKQpRdXFStjvgbs66xRY+1p6SDpiN6f+NF9Gy0Gi/iOdqZ+fzSUr+EnDlheYS9
sN1JN/pCzQ35jv1+uPWKRTSYPhsCBUCldbKzxu7h2vmjuAxS+XAMVWMkX4yCFnjJ6rkrWErTHIp0
emSqPcThQFalV0VWyHtnVmQOBRulZGhTQ/1RyVBVUAiAZOmm5j3KCMC/vlrcw1objcXkG53BonOF
LvOl6WnNSHhx1cqAKhcOGRaWkFG65ttKg34BzBqd/29s6PiQKSMGUOzSxYPYJomhFja4ZLMH6ix/
AgK6sNSvNLr8XtTC1mnrRn47KWhAPQqLV+0zCV86UV5j6JFRd7oJOjcIh2RgIv6goqhqzulrdYPU
3YQCGuc4iC6U3f9TNqTqnC2K1DOeBJmXAF74quut+db26bB+O2htK4mZO9z2keYJc7o6cGKnZid8
qfl7EbGKFLeL5NKVUNgdYflTzyCjpNh6owLzAi24/hSFS2R5FHYP2EBPnYbfy52BLC2EuBAvsuUs
IwzsQWo1jOvEpxuBDrNpgoSlOUuf/9WGChT/vF2eoc57u/lMrVBcRnzIkw2ZSA74/85Lk/R6svVA
WXQHgiR5dZzaC15t+v5CtpKjKjAqHnP7jX83vAHFID2Vo+O7vKGEO37mlIbGWMCSDtwXDezi6CO3
JfLqZ05e08JyQ5tpFA7AhCi+H1Uz8IM0jp11gBGwoepbXkYDnN0UHxig0HffvY3wLPfRCMIiyKgl
S2xEOxuYk3qRIp7W2RvlQTtog45AUDPz17LIoBlE/cs+zUvLFNYedub0ohOMMc8JMHyUGXxndN8E
aLUP7A1IVXUVhoE7sXH8ylTz3nRAGrK5oce/2T5QMgxIU7kOqlPLV+Mh1bDwmwObX/nca3TF2mgm
EUkLxaRDcgNiIszFjfvVnZzb3JIRsjCTVyRd8ag+iJfKCg0IlPgmwGzNZY6RO8G+iwBo03XRQRwr
2rKG9CsyyXkxf5wRMLfTUWn9ONG7vmoGqtbBj+vgukhg9MBj15h5214wwU4Q2w7Bhbh28XB5PebA
vJ+hrJIySDbkuT8gb2QjWXdLmW81ZlPofH++mSyKvC/dZExkYRI8JmfuRr8i9CxS5KYfauyIxYLH
iGF6W+MTNnYrY3tmWJmS0SipVjkOSlX9U5ZBPLHCRHuw/1pQvJe3lC6VyczIbdTLEwAxcx23GqNH
ze9Mw1HjDBNnw+5REznDqVym0yeyifQJ5KawDlSSlKGvucOU5QEMvKUz+tfV7WvQpPHxS+r6zNR5
8jaqTCWj21EaLqJvAjo7DatGNHmK+rERZ49oevGUS4fBsSVBrtR81p+IsINeYoKmtSB2Ceh5DYBz
O7D7UAm5ZC/8gW4hXZc18Ly6xqvWX6HFw1Pg9xC+6PfC6ak2fA3hQOO1tFUgoQv6kYBS0R6/aUC7
VVDg2xgyRg2dmJ5r6Gm+dCkqx0AjgUaL6A0WJmBbm8lWJRB/FJIUJTBY5rgZCZvGO5SksYzuvL/X
oRfiBMen9fjF4EF1AvgtlUjfTpfnKFzPHzj6dRkhcdAP/yMS6JSeKH33nG7Y92O0uLwV82F9gQ5a
xLZ1j+ZluoDatcTFXfU7JRsYwq7C2EsCyxsYnV1v4g5nK2mL+egLrvQC7QLwKXV+OcCr6nkPgKf3
XNjHj+bTtrPSwvphTR8BHiOryZhxvcH5VFO5vEMEfHDY2sHf9IQONo7IGr9IiWdJra+8qjVwjNZH
uitbAHkPxv53yfYNEqJhX5jHH0g9DBPLdOV7HRTadNFPdPok9MH6bMgUZWTZbgrXuehacFAcTnq0
QnsVj7BFgVHcS7PY5RD5V5Aw8+tYXibUn1nXUHJKI9hk4mSRbsV2TwIs2glnoAKWotUrUWWD9baG
xuv96oNh2ZXYvzCiLTbeGMCIvf+N0fJuBKmBPnLGX5TTPbzwHSjtx8geZ9yg10jU3XdiHSjbjo+p
q3vXXkQonBxo1xAXcQ9BxKSl/C2ziOYv1ycp1sis5hbBA1PpSHJAzPWkJrUfCilpfqiC477ttT3C
4KniXBCof3CVDJO3qdUxvtK8CqmZPyndoMqKaUPFJW8MH0aHLvNDAqr+7KlZq/1wac31kcxwCyRu
skZGtfqM14XUMDTOmLqL2jKdCZQI8qzU9AqcnWQDvwqub+YHt6HsMPHoF0+7xOL6UQZgxK0YEZjt
Yj89afaarZZWb+yYIY1/kPfZARpj8/IxIbUpckNOLLsls9eTUZll0Lb/YIxWP4yV7GQ9Mh0LkKS0
cH4qT1cmQwwhZAK20Lo7zcKpB3pmePvOGzmL3px+GTUHne5w1q57SipJjDAKgPKjoFQFzMCsE0OC
a99+X6UwqXeZsjO8pE3i5JI5wSNRv8igaAjWkWHE5DeSOo0DRy2DqD74l/g3Np67TWQj8NsYEK2f
nEnHilgx2PbfQcUGLIyhod+M61xW9PTGILrjwu6tiGNFlUThOfJqgEjakQSk3iB2wnwEuApS54nK
MltAitcHwhRbIWRWA0DbFMjot+ZrNCzPkukNngsuMpYmsBSeDal2kd6Z7U6wvTcvBIBYGwWzDcC8
fWCXKDaCZB7tg3t+bJITeiyWxh5EnLhIUYyq4V+9VRIpbdExgXIgf0FhKYXbkAAx+nt3wIajFi0N
EmzSxPk6tYfNrEbbU4ZFxKYV+xVKKVWS/a0oF0b24H7EJGEOTJT/+UFF/QR6wEcXtEJEQOxYR1Ai
n8cZm9FUnPCCsNqR3OWYTVN+hP2JsGsE5/S7tWYcNV2qPOIjLKBFrkiifj5S9fgqGGvEtygADZZo
TGRpnt6XKg2PAfeUSt+mxplM95lShTIxr64pHUwhx6i5vrucQ/gtG95J6e50z76BeWF4g7kXtYAc
lkFgcwEJ3SaztYMzBMuN4ok4nDNb2NoGWHNi2c6jtSy5dP7uTWzWVMdckv1a/VIosBWj3iOPWe34
IjUP0lClGHS9Gipe1hCO6K5k35iuxMYhJc6p6xUvCa+E1qFq/gviz9NNdI5Pzq7yJfCXwMme7SUw
l91oqXy6tGxlW2NPKicezAIAu+mubufCv+geatOKZZQ/YnRKNJycAZnXlCKJzCgk761DrX8OBxRH
4G2UBEqEwjXi+Wvtp2EnmuMi+ayHVmSbyfUMK1J3hOPB4kaJjun23UAK9zLjJcTyUjS6SAEkfXSq
18vz9k2aLfpMn82ILoABTjdFGL0b3YzjLBX0hLBPoog316DwXwtLf6eeJDpftDbTpS5UXsyigJAo
KohQ2x+UnUJX8sZ645K49nC6jj1jA135UexnEIRoyRGJ4bNJSNte+xT4+mn9do+vVs44DJ/u/v20
V/mjH8JFvgXBvsfuLghCVQpMyQjzYR0aKfBwMWpyhqw3w7Fw9LyghOmXCjdUJYkifq6v0VRatCtF
6BxPK7OcC886vTKriEYZWEnXIR/fRhAJq4t7MdawWsZq1W5lEi/0Zre3gxkqaIzntCKFGIN210On
euG8A1ZkRn09/IIwlPSYR12O0zHUizGS8ZiXUEnM6qwEWSlITqyWxZpINXg9umLaQ7+C12AhZ3pD
+nCCG/VrB3Rjd7i+sSV14oq19lW6AYo1u40rHGIJ3myfAJLqFDauASCtkQxUM0HhUz+TSjEDjCt0
LWbNzMCUixcJ4fS/IoaIgs0P2OGn+Pw88+4JDurWbGxNApCqIMCmHVeSqUTOgICk/rGMSMO4WZJc
Q9H6TBfWlt55lJ8wuyykQS1SSJ+E7nHoE1hd/gW5nPX6FGDODqGU6dO1EVx7aS/OlgGqk/h8rZPq
h3IKOSkOiBZ9oRLZx9eQ/IA16j/aUB1rS0HFMxUO9CKfSPU4BJbszFccPhf3gG3Lt82I+ZBR0mZt
mXPhofxjawOGIuJ3TTWdJzJI2A3pVh6iclbwpLaWiCKS4S1iImNR9JGK4s55uJjyu8fJXomPTRnw
QZ8yhMODBlrGZgOKY/+YMKY8IeecU3EXiuiYtIybt0aCQrXUtLu+gLvCZ67fjKWGtnwC4yV3vbX9
8zv58o/wpyEpA/v5nRsU/3sXzj0RjvoIbIyDTZqPJOcRC37uDYw4r0S5xrXy1Mdh3cnbFCLGYljR
PBeGDGr6KqIcNZdntxYUUG1L+Ybcu9tppUNGKyt+rNGLXZ4wU0LoxGAAQTAq4x9og9B/RFv8Msjt
hH6fntc3psLE+2djqDB8a3NNXCqnuB+jODyP9S81OsQyCaa81Ef6vrmzBFLDB3PociRUlof0cdVX
17T0qBUJHyZP5/BXUW4BzSNRoZ2KRBA/cjq7doehbrhyUocZyKEipcLUDyDGUgMjc0Jj8FEPcEmd
fYa15sR4ib/YWBtHbfVaOXUOSmS7bzDyOZ0okaOOM5WgmoITI9486VGhOhOlx57vaRLJmgimqbdU
VTWvBjU2W3xGbLb9ulBjIC07E/329cFNsBTwHnU8ztZ8GIne9X/s+Y/ISTeHiXIc9Rbg/s+tNwqA
rPyAlmSWqIHqfseJZhgCvK497CRLwaYAKE+e2dB60TimK8X7V3NIKeFmEY7zIJe2BM1S+EDQWhlb
0KwnY+PE/YQo7dgtyWDiL4dkeLKx0Kz2ooXira5lrOLC728Ju20+5z641E1Ofd4n0uuv7K7CNH93
Pjg+I9VNwanXE/Rg4DCbWkP8XrIJEoY2/VqX0gJTAy6r1DRkaSQhp35nEOU25xKB1qEE1jWMqWn6
ox0Edr1lhX21gRpBSeoUVmCqw+F2pgkVSzNiElUD4TPuIf4Q+l6elikjOAEgvbPsvcCh9xLD5EF3
Mkm22P0twhcPStf//VoNjRWRm3PZIBdETfOPrsQAiR3Jfh4yYjwV9uRjtnafTteqdElAczQArrSP
dlgM5uN71ionqn7e3JB8X3O/miLEg7kncVo/o1LKsLQ3HeQD9be8tCGUEvj6/4DSF1r2jz9JEMfk
J6f1NcA8uGCIQn3iIGTX1yS8zI+Y2XPeWzGpytYI5v2r9JskAYPM9z828Ej41WmWeCe4Q7D0Hgwa
/XcJ5AKiZgYOaTtvkT0aOSwX2+iwmA0ivYzhXkSIDXiPKKXDUCdTykkXhbA0YKx1so1d6yBsHHFT
xnUDy+wN41yPuATgdkERumQ8djRv7c1Qh0GsMyLbQR6kZPCGuN5IxWvIGiWZvNYecuMgTfqzm94h
QFvlZY6eL9421qEolK9kC2p0ZffpZS+rE18iikBoAyNuiTyax2zPZsETDbyz9Xl6641v1BLmRKby
qinPQzWMhYdnGnHeXDWb4Q+d9Tm69Tqat6/XwSWbzv+f0XhvOp/lPHGabM3r9ctHErlXGngTxuOL
/3gK2N/ia1RDZQEBTxKhGyffdDlbDaTtAxNLHeI9sgzZ6/V9fFMntoARvfYOr7yCLkvo5iWRt7P6
/B838OiLDv1Pzs3bCr+U/RflIVKyjFb/11PZUkydFJmMxH+TyOuKQhejLvSQzeyPXa4yxwdClo0H
YEWz1BqUEIsepu6s5MuK3IHoHT98AL8NQNax8RaE0qUm72sml9Aoq5b4QkNDUJSIamdoZ0Nlw+dS
3EU9sgG9iVoqol/XvDVIzbC9TKyjfFIu1RzWko+FOylruosuXexy7a3Xlcz+ki9YSfnfJh08zrom
jm1QJhTqQnEfMWPbSTNJNevgEse1aftovPh9uqRClrnnH3xf/FEJ9kNp5Omz4SR62YKxLnnHnO96
Rv+Kuit0Rh4rPojvSsKBYh9EoDfY3eMVx0TTO6mHaE34VTUcSKq4L0jk4DPocqkaTAWkIkWr6k41
2rTBUpBGI1uTVnoYlVsRaCRGzVuWjmEadk71HOUpS1uMGwa92KmIfCVDqVx69kLdlnRMFs3qTgkr
+MOOPacXh1ZKiEMOnG8K7YM0tytl3mdLEsGNS+nB1jOC6+Nb5t8x7VsUvhuS+FCgXOYNYCeoZG2w
mpErktipt/0E4SPlyolvAhvw0yqILu+cubraQIXuzTxLLZtoZs0R4xgTXABiQrPJybZsa6u25KZn
MUhTWBuFjb6feWT7ewmCDVGMAJHEcyYLOCZNsxTaS5HE4k8MZOaXT81RcXD92LznthLwVsfRWXvw
0Fvls0JJg+AiZDdxc3o1mKoWcX/KZw5B5qUPvBnKe0E5fDLsaupt+rw/b+r+w+8D2vhh7aUYRd7X
mYsOA26BB+PCfg4EwF/36gxCnY2bHDcK7q16dL5JgHwbgd3NPCuCK7gjlvXhGertNShF9knilSWP
Vjk5z5vQoWCWyzKNLycAmRbcC/bBPaYoMtPyxf+jMjp5+p7g/Aqfq2fIsXw6ScH2X279dj+xkypZ
bqDk59ROiulkvRfAWVPHwhAYkUpXK5sPuv0sjFbzIKKbsqxUB4G4bCrUhDKM4QdrmcubYrdkOXjT
K03efuPQjhzpWC8CsPWXtfysgWqoULCYoq6pEUW9oDZ1ZGabIZ0dl2FkNsy33UYzLTR16bY586IZ
jFjQ7akUAjHODXLgEI7rL4b7Cy5tE6nZ2+nmi0f18utyKXe6Va/iXvvoJs+wbY+XAR/FbFiH9APj
h5X93SjD/ckRxJVW/bBEbdUL47nEZ0JBKdLJEvegwOV3VZNoDlm5OQQ2SDOZ65koPLaTmNWtVLbJ
NZd0bYrOjq+b2pAR6Rgshc0jJbvsp6w4ZmIPSfxAtud/i1juLqf9kxrtiDk795LSqIZQsgT9XuqL
pBdQ3B9BIKfp8As5I+S95vCmO98Il68CeiFKOFt73cRqSqqVDeiQFG95+NLoBd+O+jl52GOF7iTf
fO9aI3QiZoiCBtLVpf1/3xP1NKzKWaXaGlouv0GKv+3ujqbEBVKOyYgTS6wt9ezMT6+kGLvkQE/y
kMfHknnVdu03bbw9MeBa15IyuvEQgzwIVqrTHRBl6vFN6Og9P/4qXVt5ievfWiO/dmo5Lta/ENec
knPgPXX9K6R5vHxkcCWlgf4v94pAWklhR4gJEYq7oyCsXHQZHZBWb5C59SWx6sCy3dsCr+2pvTFW
CEsVY+TslvXtPJFPlFW3A9RY/KDyPd98l87A60rB3EPawzKZ3AxJeByC40tHh3CqieVKod82qKhJ
L+PZQLwGXVT7fonHq94pEfAUH8SQiQV4M2zguRly5RxOAcCWoTmI6g/Xwi9iHOxxsw1qLIHQEy8X
Vbf5jFpHwCAzSk82irlUFlTKKTjlZGrSmw/hx4hb5aRav4OYvpXnWI4GYIZMJCSDidm+GNrRSFg+
wFYhpEZj9rQ6bp+MR034HOR1Qfz7U2AWQd1udY56OGbDVWbyaJTyvGIFgyOIAuImr7NsxnXafnts
/fqyWm3ZI3IJu/bwVtgKBVxlchZaofwDVVGxgmxiXKXrCuVlbdJ9IJbnwKEYGxPEgTXpyZj3MB0q
MbxWzVU9vwIt1j57zOn9adBeA6t5yTokNERgrLrYDEK1d7nA6iFBKMo9m2Hzn2IuiAGuiAz80+8X
gAx6liOzGpafeJvhU0cvdXGWHmCfPgacOOVCT634SZsq02IJpXjnfz/hkv1r66+fly6PruSWoE5a
af/QMR+QrCXPJvV0m9BbuvqFy0nhJcV2PwTsurhqJlgWRypNDeCUceQdfjv7mJMvSYvpMS51q3wn
tiE51qFLGrzcEt/BvaEEB1VvzI33RHe5BkJgXYCIWGDyQhTYGwuHfIY6yxdARiIWGunU0hxnkm1Z
LQpTMWzxdfUIkR7JVE1S0WlTy6Y42Zo+2q/OBrbteu07239g8NVQp04XahbOwkeAvpqKP1gj6RXk
fv9In3AcB1eksyQGis4j5FdAjWiZE3CO03IGRsjHtP1TRDtcL300j4o0Aj7Mrqzy0T4Y4es8HkWn
yZXNjVgY4A/pCuURBW1V7AniLCnAV9jozxWKaifPzyqQSvPpD/LufhNqTeMTkDQKMeW0O+Ol8Igm
qkqlFUdJju0RkB1JPNWSSiauf/+/ohO+VrkL0UHmD1u6xDnsW36jqJmTeWHoSABz7txH5i1dacFW
kmvVY6CPS6hnxhqSsQLaE8fRABvMETahRsyhg2xuCG5qaAkhrbYkdZ1i2Y5mDzdkUeWamBh/eqP1
iK3BUmH1NjiNt3iP7lkLs8GuQHML93A37/q7Xzx11lCRj2M7AzvLFnO3rzr+6yqcwPskuauEn7Hm
u51nI+2dUUI6G88qW7CP/dQYa1le+wAD5fl3kzrDsdNlrk8ejtFLYMk0LbPXrYLdEko4A6QiY697
L1U+XcqkK7AQL9qfLDJJL0v28PZjwBrs/zAj8grdfK12+MwoFuJ9xaSEX250X+GL+Vj6blzX9qz9
aE4p9N959UBKP2+vgM8DCEvnVxxShsAbjWAImEDXujwgoC1dlJ/y7+T1lXrF9SLntSD6E2fW5mgW
c+C1sYxHt2RAU1F3hRp6Pq3LX1BMeKnkWkNepkRjepXfoURVXtN4CnytXBKrKNMQOmmZAeuAdTWp
i2UhL/qWkSCRbufpwQTEFDozodLvMldWA4LlFS00QxrlD8k3nPFFpsoV7XZu82/n1BgHnVxF1eA1
dprHL7dDRNC/qA5trvFgukP+LAP5uzkCd/aZt6r/fuJD6O6c8YGi0r6B0eLmEapROXHekcogILol
oE3R5FA+jnv7GSdtunkpekoLnIhvNfJIOTrFFcRTZn6WuE1lYB+GBdzQd4Di3SqSgZjFdHUQWnpS
FP5JdCeYZy/VEPqpnrDzBJzSfoYC4Vi34RiYwMU7mzutLAyeT62MqtD+mC0c/kGV9i0Y0mG2MkZ4
zNhXtZFCfbxHUKQPlYAhwlhXPeAbKlCqUpaz427HXrI5gJXj2IKecm3HMP4bSCq/rqgULRlstONW
xnAfRrq/b1w/BIF622kfwyHcuh+LU7RLdCpMQa9v4GnJk6xTJu/Os1TwWtPLoUpmw2Jj0taVVY3x
N4J44rtJ0nKLU0T+pqcBCgRFpu0KyU2QPmuGlEF4B1ub9DsDaZOBcpytg0J9UKeZvUUQFkcJiJyQ
wbamjoqNBI74LOPcB+KVxSbj1/JkJ1t+EUPVjVC7zSHVRerylVWpafs2Z0SqKO3xWytx3Hz1W7Vh
giG/ZAScZPizourKzzt73J6PIN3pTu59JfunzNjUI2We9EvL29fxcVeag3DBKKGU1Gtu/fbXQaLW
iJHp/B3wBiRPXGfHEq+fAeysceiHAzDMqv6Q4oHWFN0t+CXiWTlY41adaM6BTc8PJBCXuTtBnzti
AsvYQ6VF4yH1fHlcTpDik/9zqYGe88JloVOcN9vGmwfW/SLEAFCUgx1l9LM94SPGBLY5pXfKGKP8
P9kjdFV70pSaOsNx38bh/YhA4tuDlcrFuv7kdPibT+hh0wjx+e9LMrBAXWGUeUBo6FF4Z4GuvoCh
++/1cTdsMUQh8eRnajlPh+3jNSf4FjX8APXFecGGWSURLv13v0Q9zclUSrH3AnNx7zIpRl1xfeAi
kfQkAnUswNm3PoO9XkNSik28plFb88RNT8BuOAD6ngBWfn07yiOVn6fGejKMbVB7GgngblyzFUW/
fzxM6jiCqdKg22oQTARB9iE1POir2i5AXD+jXJ3cVwlTc/R1Q8aGnq5f3ACUzU1doU6tAKKMPq8Z
uiipqeSm7ubmVPW0nM0KvuzkDPWVFiBJyEz53dvRo4I5r1Tw7N4Y9zA5gO3XMyRj+BCuPdvxoayN
MzNFmgZF2/l1Bn4Du2+Cox2cPCRUC+zRPFeQIH5FX5SBSwb5r5DU8IdXg7ni4GVcZ0hmGb2tiPab
ZlNQS7xnaPBoZ8bJQfQkRvtkOlln+w/zvi1wkALQPJTF3q+cVC9n/PuWrtIzLdZ2rtlc5eOssNrF
VRLoPG0+0KGk2hxQ37VIAou9v51MRstJdJawMVkHW4JXwWb0WGgtXR4/4pqdLRSRnlsv54vot8go
pvMcVUFRg/UEmNOg0eEV9nVCl/1hZqkluDn097SHntBD9QDIagpXBq6CH7zYhr1h5RTqvUGSWxVT
Ht+tKJNTDg59U3cCgeOM+vDK6A/aFFz8F6lxB2OKHay9rWc+emEAci/u3Ta2dwoa7UN4uWT0n8gI
lyRGv04J7pHJYn9TRzvBdPhSsraMEC0tLzmreTis4whgvS44AtBpGFhNxzbmkDivfwkTMB/h9iCy
EWrb7ZS/3uOsxC9pGphyazo4daFr5rqZpltt9ufryd9mgUbsBpkAW5B4wEuMmmFwsAKN1WFuAJxl
hofbVdVorDTM/pc7KDpKZ3LIE9ZF+ScWqfpV3JdBdQQ1eb3yOCocJ7k5HhR46JJYn0CHFhn2HcFk
bp1lancDN+4e2uSh6sx7iLXAtnFyfH69nnB0sJ0TFWxI5V5h1fVmp4pIVpTWWdCpYUwBevBxfvhS
LRiImKtqA3odkpE9pZWz3ZReHLW5e/Gw2ph9YmJUBPOqShMr4KV/w2xFnG9UD5hQmGKTKrfVoLg4
H5wEvJoNs2fjajWu6gXzf4tiUL8Ox5JYv3W8E+5KcZiwpnd3LrdBzlWXN8YhVGd1nQazdp8yCkI9
wsF13Lt9t1VoiKXm5RWC10Ky8RLhv/lBsJ91AWR8bmgzOtttdMNUqBi2YYPxsJfDjtyqcFEehTqE
sYWsANK+aT4crkuYYi4WahSZq65iA4T1lc49aAiUgQZ4PqgilB7NYMd6wUG+hutor2lOh8JIPrlk
1xEb1LZkvVhoKFY4tF65mOVymBfFBFRpfAYHho8b6raVXpQ8sw+DW5dWbisLxIq+qzTrCFMxxN4d
Jew6VhZyvuA5zzsgP3QRzMHuaCT58ZpWn9U7CksGZSQ2qFeyTCRGMJZVmgeBPt+Bvj5aPeVqhaBy
zflBZALXBJ4AzX8bhG+uvAcDcZTxu2cLBFTT/3mlfVi/FNq7fuJnthIa8QVEXNT+C/49d6sZS0qW
xBoRlBUroWLQWJ4S2iXuXOQ+6IQ7ZvWqTEgUqmMNEivA770pv3Ug5/PLgoG6/NyNcOVUetOzUDUM
FEQHZ8TxfN6pV/k4cSMXK12+J7PnwNGD5tbyPYTSONlDsXMYmF0+TKdTgQ/vQ6db1Gzh7G6FnrNl
6IIdrK40OcsD7RxOzJWV3a3Vj43Mu4NtNxC3KhwpbO3yfh7XrtLdre2bgoOsA0jw6eIXNQTh90eI
5U7jVsZ6Ah96vxXpRi5Jr1tMSISMKSInhcusaLR+6g+L3E0yT7tE1eTkk2a22WIppJIAL/Hdvlbo
+VWmBJ9fFuDq5BVHApsarQlfL0Org3OW6sKvqxsjV7hlxUBPc6YmHZzMeOTSJYCCjlCUenIh6Wj4
snOA9EERsTK1boWK251NaWYX3+wegF2P1J+yXJa3OhsIydp/NHP4Cu1p1HKDVR1ph0MIQ39pZr4K
2LIpC7K9HhV8gnGJKvcHSnUPH+PqKN7CiRiefagb2I6vRM8p+6mh+l/NQwTnpfNPZI6iKGcYgiuv
J/TJfMGFt/kxZ13DVvSFuly7JYEjnNwx6Vzp8SNl82UR193FSkSphj3k+j3N9kuYfE1vDMCMOZPo
7ZY96oi6c1bsjr1QHdwEoxK22TCUpHNNAELkkCcB7MWW7HVEyaM0DkYIm3SPmoqRjMFYLTgMnBO8
fTvVnG5K1Gl4pc6K8GyIVByVemo+pAivcjZVOML/UZ+GMOaVC2UCSypzTyUDbciumTMElYubw7/4
t0v8xe9l0M5LBAHSTNuHfC8XRy7HgqWnJhM3TLEHA9t+xxegTfVWC9kGn17mtHbQEkh70cTsDXN1
kqKdb0AI2bqTMBVV06ZKqHd0pjrzYwHw2Alkh+0CXwFSOgOpwn3mdk8Ur+cEy+QEvdviWZ2r+kpF
dUNzFiDB/ovb5IL3IAm3GxhzutfRyeCmJmpy7arQfusCdT/x7u+kAby4N696ocR7T9xPO4GhbKTP
OJjTBajQl4O8rq89uj0T3TTioTmiAofUbfZGSBCZzcM9gFStyCbu7kuREFzhRTf22uW8akdWCTx1
xqSfTOosJ+Tlf2My7jba+Z2pb1o7juxq1g2H/ndijn2Mz6dJihAGX8uBwuG4hHPZ3U2A6OiMKCwU
bI6c19eAKdom4OrDRytSvC5vWzrrif54yNuUpooTTvBszqEf3+jXR7RnhHkph4sln70lijWmPPf/
NmPyLIobTFkxdEjrcZgdPV2ZDeBGI/lCIyqQxWQkEK8CNXFEiwed2zO3xd0rU+b5ZbyoMEdeSuf0
kkTb0MQRHFKF6H8OpU+xkyfVYfrDywbFGfwVj32p67p7VUB98VAi1W5HAdqKt1xDupolLVwbnoS2
6rSQpZLufZB5Z7R0INoAVdAmkqdH1xdety+S+WI2YDUHHFGA4vGkEFZgdU4lUIgE8d9zch35qJrI
ZwNHLSb1QgNN7u0TZz72qFHOUUzvV05cZYFtVmTZvDUdBWKMAyAFB3wcUDaP9c7XZzAnzPZeL381
Mk2gLsZOdzCp3JrM1eKLNenPIob0ClFO1qNuLJpdELI1aAQ6jvHYjha5cV5NteqCnRMV+6KnTW4X
tJTJcUEsRT+kssaj7gDAl1xsmjux2B1J8hdNU70xi40PYq+OACacJ2yZw/QApzKgCt79lHnWniOY
nUAssCBLUW9jvpoR5gpb7Lgjbyn/wnFCioNzgrcWMenEwzAO89L/SVo1AJiNadNe4ZlNlZpwhcbh
6qx3nkBRp3ruGuItjPaJ5ImbpfACSD042sN864c2SHtZzlXqXVgBh7FNyd62D6FMZr7Rteulwgpj
0lkxxGjPrh3T5dutzLyYVwObkaV1QJdC/BQ2e3R1nCfhQayGlcz9LNxAFEkWW0X6JHYx2iC8rVrq
8QoMy6BybQYCsmoxY96aHUSiT66gfo1HURDTykArZkzmKR6gPn+2Ni4LpiFCLRUEL4KoZcqFdHQL
ato5u0Y63LLPjCH0Ye9i50F+5LXOX6none/Df4ajq/sRQwZt2cINIShYUMR2i5c1hKBD9lPi67xD
yunv5Eh4UlstFT6EZHM3INkZ+1zC4mOHfLWB0Q+SRNeOMby78Jrhmij6hpbxYIbu2n64aox+gRVT
WtHavUZxBhg8x8WnbghKOa1LvPW8GKosH+RSK8wvmWDnivAti7mZPSyrhLW/QdXfd4P5zlb0M+Qz
4aE7QBL2/A7FG1NbUrUGbLmDBQw5v0e3fbXCtyHhaMP2pZgQRfXjJ7z9QLV4lHpk6mwtEDGlRkfJ
fhTqW/i/RNpQyBHEaQ0jIpwg9bo9LcNzXK95RgfxLLSduVc3e7LlERxMtLMzneWaIMowRStuxN/R
RZNVpL8o7K9YzxNYWMj/BIZbNHFrq0KxoAJacjkeizfVF/2zhLWRMxIaFHgP2ayp3kuw6J2DjyxL
C9kLhd9uWVrNNJfTqdyb4xBF+gfPRpATAiWb241t1deBccdVvep1nRxEpny1QK2BKDL9VCu2ZNCv
yzZB1kWesqwu6RLot4ZSXuNLbNUdJxzrFzAfEsJdeg5qz87KETeNJBbaXHf3B0wod9mUbX61//5W
qdbc8t+l2i0njG3gCGuCNT+aQW9229zJIJkCxTNO6cbOGH37n01xX9FGtDVq9rrb97RXa5BR0k+5
qanX1fGXhwPiqJspKe2/2JLWoem1qirUJbQu/H8LP8J98j7g5QSrmr1hzdKHPfjCvsqkqfiaxjLM
r+fShE32JRn55K7VPJ1ExFBwRzZTkJyQS+LXzGQKagY48BX23jAesINd73J7liHPNcCafZKpDwEW
hUz4cLC8SLzo9Gdlh6n5H/lGSj7LwdcI07KX7u7QG8caHKeZmmGnB1FQmEen/vwngVpgDzdU9hN3
DS5OKegaGJovBE7nYpF2yIB3enUUv2JslpR6QCRGt6JIw7XvYxsS9yPrjbDsGg++iyf9r4xXHNG/
fw82HkOy4LYsJGH6S0biFUR//zrMyLdZ4lyJAK+f03bQCy8jzSIxa2lfGPY1qisjL1PCKLh2wp1c
EbwKC/JNoNZCGGHOPyPhkdjOM1VFypTgrGEu4e2RtwpF0IDbSTjiDAnhZI6NnVqPjDZPbnYyLWnq
zy3YXN+HKO0/qY/5Fx6XBXnMzXe9AU356szNkrpzeVzseq7GQTrpTLvQIfGfkFY7ZadV7i/dpt6a
UQVBGXtqjs1uCuYWaBcQHMjRg5NDBIVsOhp4H4KbwA3xqHQOjxR3mIvmLIK1i1e7kVE1cocQwAb6
QmdizA7qzpfiyLghXo7UoCZ1bs0if5ggbK4YyDh2Fqua11KrY/4SmoUbqY6SpOl6KqG4oY+Ck624
MiRHZtW+TGL8GuWF4MZORA2LomG9gDrKmUtXTZjJMO0tgUiBGFJg6o40zCtign/BsPIoqNuv1fvv
rO2NhY6S4NmCO3e9sULT7eBaCPKeJCTWiPRCr9G2JRhMDq3dGoH24OpTNzVtHO+PaO1wnBIChIub
NYPentwgYNRhUuWJD6l5Ral10Lxq87fN3TqHNw8i5gE8U/rfGpB5hdNmRn/IPkZQsa5yPDaeYV0T
hzLvKuzul1RPsbZfR3zDehKxy9Pc90Ec1OuuB4jcRNZk+2uN0BIKqXnq/bknEDt7oIXtmdMjEH0V
FvWLMN4sKITFEeCHq3spujt0CC8Z6qa8jN5nvaeE9tOQtsKLohw7T+SYjl6MC2NalI8o5uln8YIX
8ZwW47DxDPXpEW7oXJ5i6IjxD+atKu97COsJNiH6X25MNLTeH6P55zPqLWaCLATfzWoy5zO9KYDu
ljs44gOEZq4/vvL0KZDkS6jr9HCEBGJLjYP3rehX1HlQDNcqa+euErI5+EhZSXmLLo1TEIfER5FO
GFYlnBN6DjC0FcydXHg1aLYjJGNIMU2+t5zwpLVwmC1dg33Js6M4VJVUVaUy8ULmtqmC0GeOAGEk
6EgTXTRw/WsjYyyKo3md3Z8mbUcIjh/KWjP2sm1313tzaKbF/WWaUPPL3VJeCtrRUecCPUi/0q9j
prvsn4HJypjbnjKZu7cW8brptuUjFKkmpjwSdNdqzCDkQwh53PtgdxIceuLg7/QZONP8h6WMbE8u
S8oyMPASQPagCYFZg14SE3UkFF5A3yp86TicqYIgw1BjKfSDtjyit1J49FeJyAuBjIvN+M4zG745
LGWZEc1qDeCzdgCeVi1h76R/FZrweSbdUFztDl5SSgBngiliLWmwP3h7/Slp7r4DCA/B2U1EhxRK
Qrej63BfnWbIFGf8w0L2wH6tQucEzJI1vsL+21jqf0QRuX6eAonyt8nK2p/53jFsOF2OXjJTuR6q
L944E/EUdhAtUFKNLbt2TV0GxDq9UUr+3GHHmEdCQvBVr0yz4P3bgqEC/0OFjEsdSqTzE3xOOk6/
tyLChuA5E7T52WdJKoLluQValN52aoH/YnNONf3q2lkmsDrOMlo8bWzGoUmXg61n0167k6GBgfzU
HSDCm/R8xdbm4TLvvEoTSk7pXAIXvYCxmY7GFrJtVBqEKzwBjWvq7kv2LN2dksY2rMi1dKoxZVNk
gUEBZgMo+/Cx7k+PWCeQqwJbVU2ci0zcAtcB8T6cvudcbJUE6Rh1gBpmFdlJs315c+O5UBbqifGQ
pCmceho/CQ/4hHFDdmgSBxURitVSA30pkth09mFNeUXMyF/Y3JYIyz46XGAqqTUYwMYquXhImSSW
nNUa76k16eQc3tMjPW84H8pHD+2yfrsJICLlXAZK5jF5MOELT02OGOvpNimZiiSWp3Ky3OE7TQ8N
2pG1d9RW5sJMMrWbPobrDSNln9eZzWl+2lE31KdafkWuFgX77G3bdnHGE5FlQzcUqWQTvwwOPVvj
XThEFEtBgdArXDRA4drKA0Oq/gkhKbOp2n3f4eLQ+0ghRa1gcvt1eXBBA2FqBryVj3iAWLy2fxwM
eP8y7EleFHKoa5+S02iFeZl7IU503XsGX0N0u0SnbdYhMle3eimvAQUNscGmEyH9I7dExSk7cUnC
GuKderW3fCRO8QEgadJXH2aEtEwM2VjgvO0oNFeV+5w6teAvlIjcmAfO3oWAyGZDAJTw8TDaa/XF
VBRYozuU58+sjQ5KWsb+1V+Fb3RNAJsEc/83Db2powz37SUTW+7mGiY+mRPhCWxV8Bq9uSSKfMDe
iDDcW9K4dsvEJY6o6I9dRXiVjMz6DUtGbQH97F9eSuw5sDFv35pIG9bxJKTnymO1Uz4denofdgSq
VthzFiriuv31Dl9ikpm/dvCHFeiSvhO3/Yd0wr0J1CwQFbVjbT4agN927Gx2zIeo807gKsyJ/EIg
Vtddsc5efdzUi6ToUl/EYM0CZRhFULJnu4K8Yva6BR7px0JWvzP2MPy1dzmOID/x3Mgsh9Joijo+
CFANm7cIqBkzlPB/NrMMW4kcQNr4oaKIfyOYczUOBfI3ua7dgQ6xZqBUeXUeDblcNipqwT6IvhFj
qpxjbHAXbjO46JU8557CLy5DlVo5cXbpgaxTylTNZzKAIhvp7GAAnWU8v9/6GooqEX9ElgmY8sjD
VSBu4D9HzSROmqH0CL9KDn5C7T2NYVbJtM9BAnUUxxGGXKdvg6l2Gimt/reHxLvphuSFssxCnrJn
ef54EtoeLGFYyv6litQOy9VhEWErcHF2Q2NMYNFoAGMZQ9UaNYyuOBIEmL4eWRK51tXeZhrPmMZg
KW/6SnP/pFsgASsxoZ0jKWNn5jZ4MbE9RyB0TAb4GXJWf3ON2Jgo8T3SVIUB/l/QKgFeFZgRttUP
khioTRl7RYCgnUG1GKVhWDgCcdOKZDzxGICSpJDY8qMDeryjC4Ufs4OsBl4dkTxefuRPD/X0bHwl
TZLhDfKc8RzBLF/Ta0W7NqXDFslyqW/UeG0XKCqDAunrLUsRpp43fwd23cyWFNnx11xD4pJHPvzA
km5yzZ92WvomYI0PGUGXM+24CmXjXf4RnJ0AFuL2nbvxv0lENp+aPw0B+wW6e6N/PebhHcOS4TV9
bkCiGonD77ZC9OFvhVJnx50t/F9puIwThepr21KiTK0oOX/wcOZ1BrLOo56sUnIwW5KxwnfnC/15
gFKVTs3SYjI8CUZ4iHzCaAOMt/dgSH4WA5EX0ubSwfQf5e3O0HbNhOHrhcwNouBWvUomR1ci0u+f
X0kHHgOySXOqZq74DlM6vvSRju5GaIGWLLPWd8pMy++zlst6m06knczT0/d7z4FX+WVM0TlrOnuJ
kvJ6Rl0s8H0fLX32ihv3ybBM97vPVqM6U/E/Ypw2mAzi9PPHMFNT8p65zJcGkvFxpAmIcV1NS6B4
rWSM7/7ExXhWowqHgzp5RJmEhP1cUNGvAkRxPshb2ebIjmAtW6cNdSyglaPXFSJKYtGW5gyXGx+z
IVOpOlU2os8rSXAFnwDWqRyFC9WZ66oA1fvJ4f608F4qLQzuK0GDKXHvnLqaPxkWygqFEG3SwmGk
CUmBGtwCTFvgnU2CBJzxjNZ95v0YFtWeDpZ5dyS8/8RgzRh44ixjRLV9JqNjVzVXSHNCyH7LSXxn
NLwK1OR6BeP58HDkw2uasocac8tHNGMYp/IoJa+6nklrM3b8rsHcAlVyCZRbDCW81NK8II94bTdE
x8Uv8PiFiMbdRl5oT1fG2bTmmNWdGtLxY0pvQlzsEderTNi/b+BKFfvrwsEEeXhHEETAwWHvNH5J
jA0+LJJdrIOYvbg18qsLCFbdnQMv9mfixJtIc+r8fsjDA4Q8zMvl66EAmPA8JY2rZChPRO+Pp8nO
/FH2XZ983oe4HXFNod0rNiyGjhffH743wTk5NPloFY/ybJjhjR5wE3R6E7zSGQFr8302iTxs4i92
wPKTLvTXlxAojiKRTRdPF8T4kphnsHMlurJOwpogF6LpGKCL84Avy3HWVkSl3r+z4/Fu7PAmCPjp
UCTpKX2TKrdKBSH4xS9GHE2dhwlCrWTEw6ZgFJtJTooH+3D0fswYTsa4sMtfDurMlJnvlVqQc/ZG
LC3LNT11pOmhxV7C/oBeRdrnPSm0NN6koGNf7mCEodoijZT4nJzAxFia3Wgo3V6XnboD+WL6t/S8
rYF8pCFLB3FhZ470aVz6OT2VlobCeNp4BQcwJ4iNSqr6KHhNwggusYHq1sneeW3WOnUrBB6V5H7j
/uH8fodpP+6mVyaA3tSfyjW4rDiHz0mLF6MyH0w8FaNHqH4PW4UwYQ9SC15HvBDa+9Ejvpmy5OoB
rd99afQHLexxatGF61sikldNnQaKVwXfJ5r92uJknyvtm1arrX5tnfs45cR0j5O8hmWaRATq2VFX
EbUKdpY0+gf6LmPIzdMPzhskKVfAnHqsPPvikf0Gw/Kn6nNODVKCf2HN7c4XvpvjRkpclo/sMHSS
jMiOzsFYIV7epsvcVW2+Iq93plFJ5PSWLLcqrMux+LTrN7MpJCu0VKuoxevSi8WM295zQH5Ls2wn
1KRqTSh1RhWm5Z/fDRmwlCOd5BvFbu+Yg/5wcoWes2ufAkaPvYdsVmWdmfH8w4wFQRUzpLdW+ug7
MVuIdMjPq4nvxTmT7gwKmWDX4vvdhOZqAApf1YJkq4dtVfnSs71h+04FTqWb/ZK8XZRIk/EMvgxr
sfaLNyiiHDPX/AXmcHrFG+B1vKaRJAtfsLus7iNQl0FDKPZXf9Gqjo1aqFovM01hHf2sn1ojkFn/
k2D58E0iI0LpHt8Vt4xlK4YnxZ5olnIToqcCaAflj3b4GQdpiCWaGYjt5Ch4QeNHv8d79VpkmAk7
3dwbFEehc/e5FmE8z+Hp0iuldVbslhxTzJjIqW4F+zp9y2Al5hhudmTANXnoednFKa7eHZgWfxLJ
gc1tccOHASDvz0x1WRSWIZiqBpIh3r5EQLJLJ+W9IrOdn4YEkEhu/8mQkxro0fRV3RnToeZwOqWY
VfRIdT++NgH3pZBysWDS9xtDPo7KsAlg84h/ymXHNh2avQKALgQHBznZH/a/Dk7vzmDvYlrdVpJP
dkmIhf77iusV2hWk90+ZFeaAvWUnZ5vMasKzuGIk0Zagou1tGE7In+A2yWCFv/4ckdIubbdNv92o
Dd+sgH/aBvdjjYrEpTkyrU3p/fX0Ukc/oaF38Pn0A1/jcxDssCvTlHk1eET3zkg5zNRtVbfTkW0E
OzrW9VvGAV+0PHYsaenX2NJXhS4js7NFgf/YO/C4N0SpMK865A4/UVllBDYjXbcJMbPQZZ5Y+Cd1
qRghqHS8KMCqrHpbv79zbjTgzQluTOsyg46m6/VAzjr6L41mVGeuJO9loQTvO9VkgJrsiPyxLY6O
nQIjIDoaEYl4yws9xfaldsfACWS8CZNfuzR7meW+r1KyQM7O6QxMY32sv38VGhfvbWxSbbE4BJRS
b48uznZ1bgD8xkGRcLUI062kLPRibkPm2yqFt3jW21kI5tC9fOdXKb8Ziy96o2Wx9zfLMcjzR+BL
BdFuzYlgkVcRy5jdXdnQGZCZ8WgdE3H0PJlTyRvEa41sew3AM1PrdHxkiRF2G8qFylht9xjvR4JE
jHfIuU+E8AYpMf1kHrZ/TPn6PemJ3uDe3Hw7NJsfkThK3YwZsHG+1X1vu8NtcMgGMA3lZjTCYQsH
oBYomQWWNMQzRLgxyDr/E91lzT/KzLZr5UgPK9pSbIJikC/qmcYHxS4Tx7Ok4NHnWDMY9LQN3yqC
1NvzoskZ3ZRl9xDLvjhAYQGj2aeryO3ZRP1wH78b9goi2x0Fv/O18n+aLxh40cOcNmRzAEEsC9B3
sNxRJRWWCvpEN6hkwb+NsF8HI1yHAy2dGWA30QaYA62iVfcz/mkFM++CRVoBr1CP5RQ9wDsvYVHB
AlEEAe3JYsMVZOrKBDrBgJW6Vbp798xg9nY6K6av6J4iwKg9TzB9HEmRGXoY4e2n14o73zcE523m
Iv7LJAAM8iUt+a8hV48NitWFaJTi3xUpYEXgjLfi6hAN2JrfUMn0BoneK7bTw9FxcPHb9vNczNAp
IMuByYrIz19prYE2not0DipY/wrR+YBWhBOCmrNf58MKRpgJYa0EYRXykLeFqtpg5NH2aSXebcoB
L1Y16w7QPrcueFvCGXi3v7BPnrdI7uf2S+BPQSfPVFqPJ1hLWNYLGh9gaeVs4IiFObjQlEDSPVQZ
odXT+XwuKhg5oA4y4jPj+OXADoL+GkDeCA29bJYrKRy9zzN7UnAEaBIzYif/mWMckss77TLgFZ9O
EysMsCV5EJXLMVMRNoKcng07/Pk1CJb/wHD/s9BHvqVY9tf8O/JxTw1GkKbuWzHRDSWeQKDPYXk3
y8LnU37R0PdUGhZ++B9xE0bhPSxojWUC80PTN3xB1EAGxYLzhqmAfBuZKEOezVUJrALlyptc6lAm
Om4yuTax8p8aLq72o9h82GXO9wzrBW7OUviFZLwHnX3IHdd0Fo/9krGOoFVLi96vpM3buLfL2eci
SZCKpw06DtTHaPXIhuxiRcpJ+1XNeu2WTCLp1NEmBDv+rWWL1uO2FPJAMRBaciiHb3jEQPlAKpZ3
K9/fuy6wBfXKTSUCsfQNEN3y2pfr1eVBwl6cdEdaWb/ZfAzmPqT5B0hRuE2XTl4DI6FD6DWny/vi
BI/LaucXgJHXbln0T6sXdtobfsN44OYBI+aLWvHuuGhKdYChA57F8wT5FhbJgzLu7pLqgOpTBz1d
kn/NiccontOZzwgLvUuE/gCXGPYZEPC0NwqEUIc3taFCi/ZtMHatQ2Ql9tZiXsxB8I27mI8aApAt
usfjHYa2TAGEdAlLgf4N214ZVXsDEolZKxW3+YDxjdbjLMuPIlVwf86siQ7OamUqy/C9V2VHNxN+
c+EivTEvPuZuXhJ9BA2OaU1F0KgsMIUgtA1vnhgPuQAXpSVhdFspepFnB6Lvh0FSwkR8BZKZNISk
f9grCgI5q/melIk+n4gM8JGyX7S4PkkiKqRx2uPQhmJ5XYea34kP1T2sREoEhyTa/8TyPwsLceDV
rdnnVva/dyPd1EgVoVrj/hsyGTwGfhQUk18RknGrqLy0E0NBY1AevGacC/c/rxQCRkPyIXE+ETVy
mt/bMnEnmZLjvl0di6LvI65sIKLgRnZkrs5g/3yKCaciQFIt4Mi2cp/v00OP7I2q37xOwhoFEMtV
U+5adqGOyb2Bbs0NMiEZFmj09Vjb6tOaVoFYpTaO4IQgbFbHW1fwAJ33OSwXAKj2knZ61aUU3zUH
Y08sBmnjxJGOI/H7BMUwkl5GNmwB9fCQL1Y5tvcG0IIOZoUNCXcwnfocKzWfBy90SHW+CA/ob+t1
3yzh6IxzluMMMB6TCNwUTn6ARCx2giKbOGM4/G5Z9eTuV5+ufApbaFeiN4bzorD/y+Q9EDbsgmVj
qYihUA5b8fIcY4qixYppeON2rctdXZQ16CVJLqRqoRb1c+fhM6o9BLqEVQfIyC+Gtub66n6tM9uA
3K1JZwg49uqbfbFp120hlvp+JNUmoxoHLW0s++A5OkmxOSVAYvqLEiAxiB8ilwyzlCw7NdH0fsir
5dyQnk4MINn+GIoNfPzcHcnRxUo36LWSSyzI69vEMDAU/RslPeiG3D2OBeq4FSvILyoGtjfBkQY/
nK09UuRaBaeEsTcknOHP9gxGgmoMTgMdLSDPFWlFINlfVt4J4BhA+wxsrZ6xEGGHPB8rFY7yGe6X
zRVkvIEoi5Qvg9JlSiqdYb+AlmHwZLzI6r8GZvFbHInFs6BENs6twETNpNNQ2tB3wUs+sqNN3NO5
x5hCK77ABFCFAjYHKYOKLRCphoGxdJl5nzB4gzA6fKrLu7OpxuT9uZG00wh7Ts9M/hEOO317Asy3
0wDxPvsoRwpecjT8REeAl+ccKJAUpJVeGuE2UvYFNA+aUzoBkAd0WJ6lzOsiiOyWX2kpffqyfAd8
gQaeaKlZB9nRLbiAQ24nEOLzI4YXEZq+JbqAHqaUF1qpGTOwxTr5hlDa1pl2tvCRqKAUbCmXKWt6
0PV10rkPATJPYZvoCgfp/Kn3sciL96NtsKoZbUk3V/d+Ttcx2pDiz5vUSfjAsrrTBkeCR1bsDl7c
0PSSvB6cCw0bdsgxuDCCIezAblt0HXEWras5ytw1nLSzGNH7yPes8LqKytVDiAQsn42AePICkbRv
GfqJsn+Nl52JBQyF9ac/8GJGbf5BJjzjr+Y+X57btqBvXJNnF5TPC7tkhhM8sPFTFDRBTPbj3g1B
bKiejou0Er+Ne1B3b5NiTKuAobqeaVQRykkVs3pY1w+aNLa2qOyl1mwgZpLWkz4k7yd4JKS20bBq
thIrIQQJyB5EMX//2khbtHeoLxwsHmxMEpozjANnPG5floqMP9+8jI+wsSXNEVVY83zdayWs9duI
sP8o7cAjNeK05/n8r6J4zOfniRo22vrZnyWHeqxxSkXJA3meo3bKX9J3vo63MQv07osJbzPfDsD+
zbbU5ZeLwemyw7yIaor1YiMzfZG6c+/Nwn96mTCTYVnzzBEbXHc63vascZzNywDXkBlC5VsfJU3w
F+7ROKAs+M7h13bzloVAAp+qPLTwGV8EQWt1dkCH8LIuzO4AABf4cisIQxFwsQdE230RIg67MMa7
MtqcZZuQW6CuHvDOubTeraU1IaiEWZhFuLxQn/vNNL9UGHz36O9JCFZ34K0EPWFIVN7nngOqAODg
hHZ/uhVF0tl0dFl3Bh8wPrm6xRu/rmiZCf1yQ6z9tCxrbXDF6b9b1gGLr3hGN3/pchiTgwwXvO0e
EbI6R7/4jJnDKOO1nf48U+D66sY19yj14e0Uo6dabZoy76AOeApn0yDFbvmbOoffytw1rVCsl7qJ
GNLQ4pblI68bv1FVv0wlcagWbflPGUlwZNE5vHiBuKU0TkR6Pu+uKCb3I4SDOBWiGgi7X+EL6pZy
5s+H1t0Bgdy/GvEO4W7UThJA/YtRYd4eWnSe4H1tC/d9KxXmviEdCpytnRh+4tyIez+AQzdW5odZ
0XkdwP65koC03Nknll2N8N8TYp0EFvQvZkqSjv8O3liXxLgZM/5z6ql0ds+b40VPA6YCfEjwsw8F
omRR8ZA1nSgKBM86mzyBRHf9B4ChMhOf3wD9i+tHReftZPj0Meva5BTH0tlYNfx05k3h36FMQW90
fdAZKNj9X95hre3HmE3AH9at2EsEDvPsuvVTBgzRXx5Iw3VCfEfhmulxztz/AVP02LqWT0EyO9lb
hZsRmA8jpbpWb7ZExIYvTs6XF5kTmTpFYGPA0S1FUQnltUJFpvRkhmFOB6CJQVccdwXQA2JoaiOM
SIJBhlqD6aZsQf+XnsNu+TGrYaD5AOxJ7jzG9h20Df/1j67wOr8N03MBFt0YmYYvLk3Lf71W2klv
2ZgWZfrfOtpc9JeaNhBG4WdEVZX1aMvlQz7/STa0b/89C1FxZR5b9arDjuiU7FZytt8F7X4Vf11b
PXDUxxjbuDRR0BuGcMVAJesWFIGLnt0wuFh/dP9gUSzyz3kRmBXANHMvLNXPrsLWwr2+0GQBX9Wu
pBtk/Y7kchqfdoR9YRzyN5m6p0GgI51K2pZqNfZ+hbsPWhQHV8XHX4EH/S6AsMseHhl5h2S7USiH
LO19/loa7u+IYT4RIL7glO06gu0F2TznbSIA3YoQQivt3rZvtHc9eN3tvj34MRE+MGBk5I+orRbW
ZD3uJ8u9dbo2Yb85vUEVI65cu05Y+7FcHXeVQ/lYIEBUnGVDdOPujPACye60Z75erh0S7Wy0z2TO
zmNME7mg2GEgQntNVLzkSx6qUxtxigfLhlQY4jedhziJPWesUooJpgs5Z0i48vzXl7Fab7k+XdHV
JQjIBZmfA4U95ZBXehYMzzhZMataQMG9NSqLGs/hEwwVZcrz4u2QqcKs5AFq7TIibO3o7M3qhTnV
yh8Tb2NyWionyrqhDNzVZyWcGugbpMqqML5/GXCWmY64G4SIau1CxRdc6WrWC06QCayDbvi/7Ta0
OB7S57hoX9dozdYh40zo8smoAG13Qd6qDNyecSkCmgQJInXdl1Qdd9AsIWBtCySaZeK6FZFi9zA9
ql9ojm5dw6dM07aVmKMH5PE44Fimes6cp7yZmhMDo2fgu8b32N236jGU0oQxknyjd88XMTcLjLfU
xJE9BuwWQ8fpnMaHr3HAef5xlSKD683AX7qlMLo8roetHps395BNnV5FdGTPiN5qXrdgbHGuoJw+
7ljYWYxUENGhPtNpuIAreJBPl2RGNGl9m//OPJ73YEXq5ov4Q1Yx925rywbcUW0bq6GZEykV8bHF
xwvAn2yjOGkRH4mPWOAuydNQBpGPmVwQ668pltSkArernofEcm7NYVkke8nIiIY2e0WT86/CEkZT
FIMbdKPLsWcXAllJBuuubi+Fim9xeAqblWv1kB30NnMH1Vdjr5ZLpb+3JGrobP/pxhTXKNa0SsIt
qbpYtTi7TFmvJpcfujY0ZeDo9ObqsBEDRci3CAYJREXvbIdk7MMOOLSbmDGoIq50+BcLgvTUBA4g
pHeyRfLV6GKh0fNrNE0BVxHVY7QNrlfvXIYiWEnIQdJl2sa1/FsUzM9wnrSMUe9nRrM6v419o8MP
0lDsSM3zSPeOMO80UUeGV3VQG7v/OUkcPl0KRGvtwTaI9Jyq4WhQ5+F4pIgJwFhQyj3Lfy4xJaUd
SWJFwD0VT0eH3lo/0BuaiNTXdw/Drl/FhwtP30qV+GBHwXbF3tOaNfxBXMH0NkFhOFPARIeX9q5m
Nj9dBLBf9UA3eLDkn4UDBQY2/nZOdRLsPbH6FSB9AgTt6GjzaeSHwGlhdIi3l71ulohDzav5bI7k
c3rTJmem9zcfhN8tEJMPhJ5e5QJrmzzjWPcvOIxbjRXvLOeur4+KgwUr4u3f6BzYdGv2hMLKtnYi
ycbusmglnx07ItWlEoh387u83xrik65jTLeajdok0YfQoT4diQ2CGrjvYnk87Lk5e2KUXnpd5hiZ
kpGPcmOZePMzq7dpZ/j5ApZO0qdVvyx/pms5FdHy7NpySibVfNZZQHCGmlB771L42zPGFt8/HQIv
Lr+vX7VeOwTvuvMsttHRNw1s0lFdsrWd9llCc0DnOp/oVh17dEk22xYiLdmuQ1CikqWrIPSM02Bm
ZzQZln6S6bpZnWvkKhZiiqy2mqCyJHKbosKoiuGnX6qYf/gfR+rj0Vzw6MjnJaigiY+e62zRTd4o
KITCMgA1inOPTuRvG+E4IXvFpGXuANpHVMO1trSZOvqMV7O+l+2MjJYwQdiB75WXt0hoOijOuoTC
6cU9khgWgOvFoSP0Npd9S7XRZe/HRmgEiuVZW5AXl2wu7CTtXRa23l9sBGt/XiEK6fwhPsWmr0Ei
aSuGWfpUzdwuOUwFzlT3hlwAjdLoMGzkViZc+3nLniGSHwR0x1/BmU+PtfYbLUBbRr+AQY35CmOD
+3GlpgpwysHCA5MT5+7o2XdbgoYJq0N6yZZHsIhsa8HbM9hH6+GD7URR0t8JQh/DpEnY/sJ3Qo/8
Z1hqOahlWQyBt4pA63np6E22KJ5moDyM10+3wpn+qvL73kyfwiJ9q0BOeC61vBUfTuPUDE3f5uUi
8rBhCJUijBhLW+aGzUVPYnW5Dz0SMQ+zcJv/pZzaQOKiN4jbvVs7nyFmWXZ8hRJJ6r5yx1Z2qD7G
qPEhz/mltKXqlKMW4EPMOVIsQS1enmBqMnVRBLrTjj0GcH8H/3jiZMlrEWRVGGGH8S/SW5HohNfF
TzIREkO5xeod3ChC8AMQ6Q222cjEGCh4+wFTMn6lPSevpb4s3owsICnRiqQ+cM3Uyk/Eo6O+OOdY
6h25CK3j5syhUEXVBa3+WtxBKdtYjIld5bhqfnkHti7h7BXEgICK9Q9ITf1Y77QemnnlTANk0atW
83LNYErZyQo7Mb4hPmOKwBG4wXpjhj2ODwLz/4KubE+wH+jt4oXn1XVq7WNtRnqtKMWde9QH2/9M
33jZOQ0SrPX6MFwVWoQUc1NEhs2IMQxs52d42KEz7MYy1CDX50s9LoyTMdLCJX+Kl1SsgZ5y9Iom
vDN5VmRbzysLtc7Ndlib14g4GOAHLuXEkv3782f7saluJAXacdj9fzYJX2FZGRpahJ+6z0qCHXc/
LiXwEsVjicLbZgIPPkopJxzK4krgo8Im4u+lhnEFZudpQ7TpsX8FGp2JkjZ7U5duLTkxLWoTNzoh
Tkckieu3qpzqZYfV98iZcMCUQhIiL/PzzThWMqRhnmp4kddwh+qHSvVuhv9Qur/edrtvkrI6i3kP
lDiRauVDypTFn7+q9miKOIaB6MWBOi/EUMhaZef24irL984izdldRsek2Kbv6WbMR2JNBsHoa+yW
iT3y6DymCxLXKyxKQVpF9K8wNY30DTVEBkS3cE7OWBTjFkZRMOUbj0SnpeVyZnsPLsxkL6K4J3KE
RdH+sIdnvCRkHDQTQGpB9dFmAgJqmDtNTFtIVtdERergzg+C7OErjCnZMF5kbQK6iHXnjqA3Vk4Q
qy/S+v8S1srKXVwzYp9HHJRxQ1B4zfIFE4se8GzSt6safgYOyxT4KMTV4QlFyF5hNgj1UKH+eoF8
d0Pi+qNkw0DhhhO2i81/l2FK216MYjIbsrdmP/8BFqjeXb8SfKYa/IL+JrPG3wCqCqDkuOf8l92i
vaE8JtvEtlA2wYVZnk5btVMQ8KoS23cTEFhTRgcCJEHYfDYq8Wz47Jcid4J98HgPbEOCi7no/1I/
FYZYcBjWrTW4hL6T795iNyA+LquC8QrLNCCXtIQz5EyqhSki5qPowb/Kx3aCE3pyCJb/bxqLlkdv
jhMVyUgerYXOWbr/vhf/I9ZGOpbGC+mUveKQQ5TDYZIQdWEgXcoSxcsyF1UUbXp2+HYLT6lHV8bf
jhsV19WdNKsdNO+Dtb1TbqIOnsjiFlHdtYiz/jkL5lF8C/MwLg7V5KBwYI4sP4K0QDUD81Ncx1Si
3CPwPi1Kez7ar37Kbwws70Q8q/B4zfAKuF7xjwNc6q4uIU9w7mn2KWVFsfU7KUgnIyhz+63a2KEM
toa1tIDMMaC0cLDqvLhKlVVwB+3vXz+KSpPHYaX5ccxl8mZVHzO6568CMPe4JBNG5Lmc+N9rUWB4
8N2aBlJDOSFIwAstWOEOrGZhyz//6bYHv7ytAkuuaNyCcvbfgjJ+03TRKCZbijx3FSdcf411gC2M
He8bjCQ/sGzfYzMlevEIxBJpNJg3CztPkNJHqEJofdlcjqB7ELcTurD0PI0ZKcWk7GoiPMbw+eCu
d5/2NvJRtHAPDK0PgdWfh3FxAZm8s4f9gQ2YF0wacGrnnXVDA/UBXR4n8Fwx/Ts2RZ2MHmJ6+wxw
6J3kLyMxohQ4a7ZkGXXzz/syvYUr1JFJXlkeCjf2D3wxB3mFie3UH8m5hFs4GQso3CD9wc7xrJyt
TtrFw8q+bG5ULB5Jd1/4ZVUI7JIXlnUkm78vNSS5Z07oLCK/J904pyshpzj6tFloLkfaqd3CNE/z
7kDrOY6LNkHkGQlxganom1IGF5u2BVPMCxx3veXPR5Xc5XJIS6f3/isQ7mqz0gEq5pgZJyRcQHTt
5OKe3ukecR6Slp/jK0mx5C45ZPs2O3y7hAF1SUEgDC2nTrVm461uLuIbn3dNmCLCoeJrx6zhSRfg
Qtw4zTp417Mm+4SlC0YFiJsjxyBoAFfD9NmkPVWXxSaJ2kk7aDjYn8MDMjM7+B4a8kDH0avM/lV3
A9d5UtCobI+yKCgQFd3tXTRPWJm4IwFgyuwY4dhpkxb+JUBv39IcXpqQQZYg10NItFJbQ4gMVtFR
WldaPRqQatC3YYzhvyYIn3MTS8kKKSEwjF1oclfTfyQj5ifsTE6Ixr90m77ugTY4UWDunXI0DE/R
0+lx3Nmg/sk/jcbTBAEhrnUkSZf6fF2gXwqqlqw4F76IxGgGYKejj6Ij5HVZl6Ck0GprjZlDDNn6
aHG55qcLtZOoFKW1/r9AoqYwyejp52gGGRvgCKzoL1+v3jAjE8aGoIAj4BA215Jo1WA89hDz7goG
AkKOiJcNuICQxZrSxwLzX+FylThl2DC1hTsRAyV5hSYGuGvsL6ZM96B+zG6KPLYp9LNk8M4WBbUE
KeXyc8GMgbo4WlZwj2vuoW5bvbZGtw49ygNv2gDEAKbHGKMBBocAjhtuN64Py7xjNvJH+hC1QBxe
9N+UIFpXiivhqE87833Ey8M0I4o9utl9RjFQsOX3MIv6Fowl0kYc1+aKUi/GwjlvVpnroS1MJOJk
DLypImpv6d+x3Nilk7pN27TR+AK5LuzpcchdjzMytut3T9E+5A6mGeNIUKd8+8V5nT+kHYVMp8bE
LSUdGqVBZLuGZqvp5T6xudblHGRu7FGsejeIvqhNK0UZyllq/d5p+36QDY0NawZnew8QwL/AurjP
S3nq5v/bok8VEJuEZ/Otqc74wcoRXAggy5zk9DcxGG+B+5fqHP1OSFeBJmIB/VqyzEEXZWDoFtVv
TLWszQQ+JrjloOGC48FbohLrXlEHWItPwrsp4rcTYa2njd8D28G667jb2zNPrNqe5AJV9UZvXvtA
4pPdGJra5jROARMlNtN8HPj9J41mPnuBPp+A29Pg38kGsEOAzGcVcj+MyZioknYvuigna7I534LU
nOcH1rI0qDvwvXjK9YPtyg1rPfAiLDui0GGiHp2qWsy4jU8kl7R6S6TOcsonm7LU9Cdh0j2Du9DT
rAAtIb56ahFmEnHqEYEN87XtNZb7r6kaIr5egGvXc6qVwYbioq8355/2TpGWIb2dG6N8SgNHw9NH
pnLwJBd/Q2LjdKBm6fKjfMdKGZnnahO4QQaD+HCjv54di7/KMhiU8rGsyv4lHTWgVxXmdSYj+WZr
w4C31Ohu2gnMpIwA+aifNbUZVc5fMDNU92p1rTfhkDZBEVCR0GJq4ftygs5KRljZ45Md2qle3jpx
MszH5Loz8E4BuMatmaJ2azPqd90jzma61sy6nufVsN3WY7UmVWg95tV0PZFzKJZkb+01WZLdsAPI
L8drTpAbTlSa/0hU+vgSLs1PC/u1KDXe39HpFbX6YEma8Nalx6ytDyg5XYqyz6nnveY5hJfSji2u
FOPUylThrckRroKrKHB+t6GTD8Lon9Xm6DoAYHjjS0vPuuv5ddQOiRLvujosOD0UBwWwTVKambA2
cWjPa1fxoFERrKvZ4g2U1KgSRal8HTw1OEw2kxFZZFcI62ljxJPJJf86zWyAAdnx0opzsepgbm5E
gSeqOhH2NvMEeZu38Zruf/wCfaoOruW6DzAmdo+b4cf01eaFMPM2mhWOs/CR+tL+vgISUMDMojtm
Bd8537GIR9uXrowTcTarRwK/oyZK69Gb2Al3REPx0RGohePleXkOY6dygDawrO7GKKbI4T+FRFda
FJgwyLxyx90BXQhvFKNcLoRM/TmNqWCFXS/slcV2j3kcoBzQdVEMMlXssvlB706ixVU1pgkFafkg
nsSE9azUBjxFuHXmjA0EQhTRFIghFO+Vzvh4fxQEU3xA2f9MqCMsN0vwKxEt2H5tta+GI/9G/9gR
YjvVwoqgStle2IgY8Cwwj/W+4RmT55Y9Z86zEeZmoB9sPtLviUd/F/m2518UGj6+nXtQABd4IwXq
D2ML/uZW5s6umZqJ51DnT3kaOyRrFpGQEen3BP2XMZ5WkGu7RkIBlNFPZdYpvJitYyQq96WkIVIH
pFbU42UaMFUJ8uQ6NrkX1l3KlDXvvhzto8SnLeODtq0e2M11WP4vXNGrf2IAOBHYJLIMwo/PNxO4
xWAb3WqzJCjhxc0XewZracVdOL0JU829Spk4DAZ2nzzALXb9xTs4M1VoS5b/YaVP62LnCLuy/WRl
gumstkl/B4JILVmFw6gcKYQOjSBwjZVPNPJQTrnxQXFsGIYoh4FG5F+iBXWZxnKjUlrSXwmlZqpm
xvjRqPqHizF6ouyx7CCIllJpVmDX7HpuOACtKhyNvUyXJoKEge/7ObrLtJb8ROqcNhAUBwnwHcuK
ylaRjkK3FSNmht06G0Og4M8lG9a9OQ5haJ+gLMcMHvUNyvDG2lpW19CgopLYQR/vAxbGDeghmPy/
vSo72u8EGHBjda+1IS9Jjlc9iz4oHjbahhjt3TUuqaf6/H1NJlBsIDDCfzy8RSB58PTyiuWPm0xv
7qZHvb3Nsc+vZylkv6xghCYdn6vBmD0AC6gJWnGicIgxUBAGczxLCYYa+j7d9w5qgH+qGH16suJo
VF8sfGVbMP7+vS2Z4yRMC6KuM7HGsKuEmZuWdkiarb3BkfmtbeArx7cHXnFCHcWTJ+DOBzeHKjJd
zbqMu+pOhVyVVhUoLw4vMDhajnSvsX9GhhgRpzKFv56WvSJQ8j6eoPKKnVr5JdMPgqFs1rzP0a1e
b8mKQlp2loU/yMp9CNWy/P0vO0pTL2Z+Am5F9XK8vqyO8d8mCTnuy4f+nSHc+UcLRtSO+HLQ5WGj
ZwFBXai1kqOgr4d1mZkqVaYbAml7ToL2zd82JJD4cw/GEF1oufHfFJOXyyw+nc3ho+kOcicHYMee
QKITPOWCWHFSTdvBbXOev1G3uZ56/JeSFNImmOlvI6kZ+kicosaozCpHw+q0jOqnb9i41RQmauXB
T2Y0A+SSwOfYLMKpkw0AEUiMEyY84eVZG0C/e4xXX7hiGJIrMhUoOLU9Ce9Qyg1Cq/KUN70W1Frg
vc4Kij4VyNgFG8OkMPuk/n6Nwfy/T3J9+bjssjL6/JWnZO0exY9UzILmJVO1JY4WDsMiCZixYghc
WCdVYT+dUXQCs/gfbvx2C1kkys9TkSyUhlEtSCCuMNn9YrqWzf5VjAOuPWIh01KBPx+vFHulxB7g
3twm+l4vXjGnWnNlC+sDa4BPqCKKRXLu7hYcM6r2oz6dq+PpJYYux5KKqWKXeyeZQEg/zLAVkbXS
8SOgSzr42hNyekk1OYQT1drbgsUqlynWiRItp/mdt0N7eH8OD2LlqbY/XSwub/LO0/+iRG+IAjOR
n4PtAwIhBkDmfrAaMtXYP7hSpzBTSBFNhO8+WglbbjJJ2gOYiAaqeVtq0Zpyg2MBV07X2Y5NZBkv
t1Upka5hPvZsZzLsfFcrHYlyfcNDj79hayFHa9Nb+erq36+zLIydwaG/GUh1ycQD2j8DVC+iqc6m
OtEX+DXkW7FP9CVEQtY3ekjNwvQJZ4XJJ8vabyRrStAVVaRVsxSrR8/rnJJoxHrCBMgBZDQzyDhF
QNgN4OagfSMLad4yjT7202SmiLLDvtD/mPUKTtw/fj9X6P+PXtQY41KY7oSuzXmpAM7FPt0GTZuG
ArWDI+t+Ow37HXSSe6Q4TJw2NGHe+Ef4OWbJ956uNxkJZqCojOAqaXf5DiBn3fJyEypMQWAcBsa2
18xEM7r+mCm3QaDHaR0/iKPL3n3DEu866ILlKn1LOSzDsyf8I0Nzm6wkw1v8op7gwQd3J2Sosyuu
w00yp2vPzdmVSSsdCDyi4aEOGXeiDZkw8IwsgGfp3rfyUvo/rpcAy+EUGubSeMsqjfuakD839c8f
WOR4hgwiwQMiSh8zuVz/H7nkQRSeZ9197tiE8CA0v9IN0zXuXabM1fdXoiIoEkQ3CqLhGXv5u/Jr
B8cKqHG7mMcSPvz+F32l/ZzZBf2XufgkGPx56xndBRl8/wXF85Ab/O5Avi3MBqyB+q61rxBGlDi1
doP+zw+4G71K7CM+8DVYmp/+Op9a+lD1EHVZeFKGQOA9gZn9kYEKmVvMfEcOk17HEmXX3Tl3VK/M
VSHXj+aJInrg2qV2g09Inb1IK1BgF9QvwBJGQzReSEBzcXDyNTRrZ9wqeNhRcFPEnVKDGWHdDvLT
u73gWPp35N3orlZ+PbKjAyN/4TsT+nG7Pbfb0XlkP3iMNz7bHz0QN3RhKhO4LouuVsa5+ON2/XWy
hbfCH6Zp3kFVCV4XhWKETT+4qVp8Rl1HGBMVuS+DKVYsSxKjXfdRknGXilCOyNeiFQYGlMG+5gsQ
KIaUV/JLZQWsYjwqSW0zO5eoBYylej1F4HcC4GXe2IVrqGPQ3vRewfqYwW5QcStIXPMf/mrIWRsq
Zcb1HvfHtiu70GXGZd5Ednw2DNLlo0xhL13RuwxquM8S5hLsHn79tF4tyHNkYasUD+hR8PfZfhXk
PitjdfPU9W/Tben1NURDjOMmNn/ZwjytdVF4aAHMUmAYxK4Be9UaN4+m3HU1S38oK17UH78J++lt
H/Wz0ICrp+YO2RuGkItf8LuTEKmbRs0lkZvv6JPDliIh9/NeXxF3Rt/ZrHqonlcFu4WtFqC2YRZ4
ir/vn+x8XMhaXErO7AFfXWlhTqqAoGHFKgErrVb66RdepJFu0OeieN+BnmqRgaWgR93MSIdonpCd
1pp2bLK1SwcaGifB8iAX3fPvaBLqSNN1DvFy8UO26rSIDMfPcHRwEow35XDAZsd4oBhW/7A8802x
41+bvXMAM7ndRh5s2pEjL62eDD5GPGxW87RFricpNBt1phJLd5Rx4kmkzQkoR4LJI40zQjcjXnvM
rTqRoTy2KqMwgF0pw+eHGZAiS2S3XoFYrKJwEdewH6zGuMDgAuZSd20v2GH5zYQwHtbgExM2QNkp
iYGG78tpG0abOA2tHlmo+skATWEWecSFYeexdWjTKLp7WmEOLAz1ECxfIQL/K3OJq4RGGMHckX6R
cDIiIhfDI73mS1OsXnWOPoXqpBV8ZMhp4gppr7fIeppAPYuLlkoezAej/HlGhWKbmXo4+jkUUX4F
X94WyENI4UGu/NbroghThNwlhscvmH27TN3u1z0CpEWOmySTu2lyHhO5KjFOaBq0jyWhoHU3LqJZ
P1nQNTxGKjxwkAdWu982YydPjLDQHD94a+Xx1LaGBQybZIoObrgCOBADHs9hpMDbc9ejl6YzASKD
Y29+13Kb5CurEco3Yu60rwKVCEK26X0wZornd6P140f9D0l/qyPLgKpJSrSA0WLOMxMBfA0P9kBM
s/CwUVWq5JA1Fi1mWitUXG4FNl4/uDLd5FS/d/IijLvRfvzQ22D52kiyfNDWemBtNaS2XnEaZq39
cISWHn4KHvu01PScoS7YPCx8XAB4XdiZJo3K1ulvDO2hd8+aMWTbmEaxR5zCnynhAwBNnt9JWCPA
tNpUtA6fjBBt6h7WFpYng+Om0pqK0vMh4rswIbrDnWcHMdsfbJBLbSE/+wd9O7cUitH0lO1aWLff
WNe/oLIiSqKYjIMF6MQ+wQvvRy8W+WVcFIuURfAPidoGD9ZqvVOExT0Hy8MDWRkfDs6MOWtKC8or
1dR4yRdjHuM2yoJL5RwvAKheLDM1sVumNtmVaRRZT4VGQwbo7Y3zKkDciRs9Z7hECSWWCEwtD3By
FD37uPeCq9ICrJEsYR8FjloX5grfj+5ZXNhSpkfoog0HBOw9VcF63GLPtXDlAWSCEcqKVAy6wadN
BmUWXKy7SZMTtLjTfU8TdSioaHJMFareCE1vmZDxDQtOyLSh/apmN0396XdZCEjVUtUEhjdX/Zx5
hrs5eSOIqtHCA19ShjJJPQsfDe79oZBBOIJe/j2NMUJ+EOPweh5SjBtKW8Zz790wY0A7yWxFKjIE
J+EeKJ8tR38Ny5c5+U2QwNvZoO+VRJ4vXJ600BRMUURZ4YC0ye/yyedPzKXnPNQ1Kduf5vD7wpks
DnT+ifVIiDkWwD4aLUY+QNWs0zpTixLxyfsUlkaV3aXU3PXcmNuCA424tCYuhCnwBLKTgqNWq6iv
vMlINs6QeLX86J067sVx7FA3FynRjiiWyjoV+VBBpEV6liZFaHLVmEdCuzXUfy66WaZREB2iRy7x
qqDLez+cyEk/QPUmrsZqlihVMb1xtNNhP8GrVqOe8N/cFbLTzIx5RMzJ2m5DI6pHAMTUBJIXdS27
ntoff6YRTgtQgIHGpjneDYvKF5DYgsUJUyqUrcWvKJSUztQu9MIuqrPxzSMiupm7Fnrv1p4pOIHL
z/gaJ/L62ElNjzIES6Swf6pk0p7s0A1Zl5QdEib8K4Rg5rEfMH3eQ2Gs6RykoaIKwH0Rrsdu3fXm
sx5YADXiAj4NqWTm+oO9Ng7uexHxYQY9VzxIh+tLgF0BgAWzP2T5h3lipc2rTJzF+ZlK/vjmlNXU
gY6rkSV0duPvG06h5IQX0XmY3DT585NyAsGPITIHSGCh0ykVPgyHMyrfJEoyBgBMOqgW3LA+bG0D
185snRPRwZ9Js8QrLEs1dXjX9QSydKV3BztqtqsgiCIp2zeZM+0uV07X9cdgId8m2g0NotPTTHrC
KBx/GEIkOFmB8fu7xe6XjcoZYedZ8NnjDQy3uAfWBlZyG9Y8oRfOLNES7oF9WX3Auislic3ZIRGp
PbhWpF3KKFMljK6H9HE6hbMDpk6ifv1Gko1vyHv1uv2s6e9I220KVa8vZCkBwC7nUBr4XhrpsFwE
bMFqqzJiALin6nW5CGQ0h2FBM3863B5CL5fZbWi+FfZtrsCehXT8GLAj9TGnIZQAf03q0jFYYG9T
heUizIl4Swpf8P8yLsSXW3w3yhgc8gEZZV1mhmYyiP5fWdegxrN5aRkyULZql56yqsaSQM7ZSocc
DHEHH0YNdKdpkWPkeC1UmKKOeHe0IRtZ+/YplbCNJkp5WigKfpeJWYg499I8Vt46KNePuos6u/HZ
ktBI5emUBQzIRHfkDP1kObMMNaXFNWm2T99STfVXF9k+sV3JGHZ7X4HfFyJSqys3078eWQfHrcbX
gaVgcy08RbX65OwRZGW/0+3lhhCcJeoTQgGZz4WTiy2scDBFiJby9x5OvQMX/Zgf95pboIUNHPaN
aiJjixFY2pYRq945iYiD4ZtEZ4sS1SUfoCEVxfj33pNkKNaLXEa1hh7RhtHLM+9Zwv7g1ea/nVsH
txvD8zmSCS5TVakW5nM+92GV4FvovCtm4qo0QSUA8eNvbm/pHeIeoCJtkG/AFlf6pRBSrjdIsqyM
p/g8BA09NCYS1a936FXXgzHw5UH/FZjl/6v5H93WVd5Lz8U9aaGk/TTFDXb3iIFcb7nY5EIHa4N9
85c3/DtSalde+rKPK6qyMOsZLgHg9u0KwO8XaFd7U4S4gDfIeXWyYwv7Esf6I4Pb6nJtoL4RVxu2
99D4r9m1314hMZWXBcKhwX2cFzxuTgn0cTRU/37aK5DRzKDcdMSrahnEi6kcvgDCX8cAEjdyJdHH
UkrHWM8atgjYHKjFofTZhGpiHwnp7HKREkpwNTGiiHnaqopH8pzX7vITW/rDlct27w78vIQkz3Y9
RGjhXNLK2kr1hulOqtIG3fKBFfSWcq5Q89x7FMZVOeihWEfi1PGR6TPUIv8Y8fq58LSYTBkMe+V3
P1mBfI3mfNqyZD3Wy5hxppO92GI8pyurBjVMZOPOaOxQirKHyIAqFpmdGdqNHQfc6Ay7PfgMAGCH
+EQxiYFRSEBjDA/JRO1IyB02LrMHvEnxPkQDvMSisNQgC6HLHiWIIxjUgtGSDNb+R0pYxAlnnizI
ib165XMXDeqWBkgLJuuffqhuK3vmNVW3Vme1VgkM4yIoY8E7f6jgMKiXY0WZrpeAIf4Smo9Fb6WF
JC2UIBimUyvt/Nl+Zh0VyM6AmLwZ2y4OaZtlRemnY3XS3tu+BVKXcYAlmk7S9lZYS0KAcnUw0KMp
mkoRF/Yi0P3gikYGnvmSeWt/jPkx5LnMuQNEIt3IvrbjgExRkn/+I5MoNUHAveSc9GNLNO457xYr
egGX1v43cFcOCf/BTKRpklFdziKoeAgcawntpEb/TSaXP45TEAQDElWw8tWRh/xyWuaUSqHCe48x
oKvJwFpWCaUJ6Uqir3prF+kOyVPT8/CaEw5kzH+6LNgsyZn/k3E33gV8NDg85Hm5GyXIZpWDH8W3
6WV2AU3HC3QlgMtdAWMeLM262ZhfrfpO3Cyds9wNcgJl40/lvEEGzNR/VUZZG59YfYmQfoLtPllI
OUErDGSA9II2EmSFqF1UwuxTtzUnu6Yvm1ktViaHyO3yiZFP/oVhcmPNI6Y2di8XY3BN0dW3HWmK
DiD8miGs3I4yXMNG0JKjAFQwmMpW1Pa9x+km3rEDkaxh64zGpSUQkoV2u/oebx7/79eDZxLJ4gUZ
PvA5D8z7S4/8NpM8dd04BxffFZI8Km4EpbEPa47Dj2jAPTdqsl82wvWkBv/CfZJY6uUgPKOnnthB
n6ckYVSPWvqIT0BEHl8+RwGblclXvRxBPLfSooB7rpiOavBEnEleKL6BpdRiWEYOj55f91ZzvYSe
oH1JEmEOpWDdEBiQ21vXhPYmLYqUmzia5vhHcbIXEMZ/5w1vd8J7LoV4wSl9k29f1DDaoBgyQmf8
bWwFYLAbzF241veREKJ5wWmczU9kpXE7uVVhFEYWBIi06LfZkktsm+YcEthrJ2k7+1dZR4BC+9dk
3cWZW1xW4gpZUiNcBD2aVH65oF8laF6AQFhltEAPS7ddwNvZPxy/qLfRFxxssw7ZwJ9dtGUEpRU0
d7aVKUobGbvk2HdOcq0MqwcXCcebjUiEK3u7+hg5RSyAMJufcJx9AhTuSCpYW/Sns4eZeix1NHFs
+lGpMtQih0diuWpjG3OFoVJCFCRfac1zsrEN6l/mzJeVjP16GOdS37KkE5UN3j9+3RFrtWJOXYZp
1BCtAx0q3mufYJDpJtfmWfCfMQGRvAmoOykBLqZB5NikcDGDw3PHIYG1d+YcKrVFzNLHkFJT1hr0
N929XcWGGwMZpEBCL4IzBzjCH/AmBBMKKqxdFNd2EGIslw7PrsHbqOX/O3zv7daxT96AAWsbKmQ4
pN4P01whAtzissf6c09Rhm6VhLQ0yuUw4IazAtNon06AdWWsHTv207uoR+P8fonLQljkwDXIyS1k
+VH0Oy7Dj5vgxIpO/SizSefb6UhVNEoGl9Hz/GEI3urm1A4qm23hIj6WXEEx5YBHhxQ3yzf/SQel
hCz8HMiPKMte/6BovaPIdS75HKFNWr5Cj/8Q1qOt3QVdibii8upliUR5c21j++b7QUj9MiOArqd8
bz5BPFtasZPkCeLG0PERqJXwRW3Vd1bOzaRBQWYjZYX4Gec55au0dmeKxuWB/klWuiOJRJ3i7EqS
XV1AW+MIzeIW/mXEvzoQnZe5USlPgpDBam2gpAk+pt16B0vQoDaGWfUp2VVX0QOeiskKPEiVDwtq
Jh1fG3DbxN/Iam8cd1sVUYmosWeFhgL4U5HaCg9uKOfu+SUalGuxXXyhAW0llSPz4bz1fdX7tnnN
xfatH9CW+GefmdjqlQs2i863j38P4zbZAnG/n/92nbRj7E5zduNGxpR702uTMmCMlyXbjT4F1Vzt
I4Q2PqAmqlFdws6fmvAxzAOHJDqAwEy9V/1kszHo/ENNpY7O+NbbJ3O2oSN8aNrW1NK8JkLtQJhc
AxQuKrggri7GtOJaQAxvF5s6RGB5d6K4CaPZ2oLNvSmf84X2M3MeVVHF0Dskvq914GFuZzPct+/i
jCOIzWbec8gtXRbxpxc2a6f1AhX+OTBWtnkuUQCIfdeMDefJzpXoR8SoNh8S9eqXZXW1KVPQgU0S
s9Prw5RqaIra4Tn9ydAUqyaSnlMtAxg21plg8kI20MwczRlzznVX5ebQXwMjjvpfTW8+LUe6N5o0
u9Q55G0uAdbR9lf/4Ry16da9qB4w/VodNPbESq6oHKeK4hy0dvjTJJTi4NNk96BjMD2W6UffKTNO
sm0bdois+nP80/ORxvbkLTrMVmvdayi9/b1n4EVMsTS1MNkVtOo1NBW9yweMc8Rom+7nxkF3vEzK
3dKu43e1gFgJNjvna7Vwl/yvCa94w5scT4pt3Y/Vg9kSIWy2ukdg8sQrzh7o23fRtENvB0YvKkxp
H0SCoScf/NG9Y3kYJ6zoPZ4iASPC07R3ccwh1OK+i5iyx9Es2hxPBcqtqiypVNz96RRPfYkKuZaL
F5D/ckoK5cO9exQoEj+rDCnSr8b6qPzEW8LdiQg85uddjKyoJrsqSyjTDfFoKXW3yfuQ2zJ2Vw5K
NGZ8mA7Z/tkHb/EYbCZBWNM2sXurjRE98wGpV5Nqjhk1P3cY87vcb8EsIuDX7VnPve07YWe7VBgz
hhf2Q+Fo85+EgtAik2H+hiBNw7JwcCcXUbZMvZzmfUGgF//6NUENCmNU3VvUZkxIQKhN6Oql/Xd2
gCm3cSQ8vV7QTu+UKBDEoFrVTu1lXg9cT4Ppv3sHTNFpEp1KNCcO+Gz31vHnI81ht3bjUZDlxywH
OYxpbx3KPys4iYfgI7H+FWJY3lXHsVFrl2G01/OxA257YmL5CM44nJW5UfuI6uma7BUj098hoQCN
hyi8mml4O7VkvE8yyYUabexZVMAuoppDqLKuxmNQRcDiZu6QAzLWW/8fJQghYJUW6iVoCzU+SSIH
WJj2kvprBx4TyQ0gCP9Z02GlH1Em/QITo/anv2uXGXz9xY+1ae1UgiZUkWN4HfqqPmpBrC9Veke9
ooyYWHmPxh1tpTz2YJe1K2ZXsEpIYrxGYmNzIDlnY75HuSGm44Vz5xOTiP1x1/eNAFPFhIxMyGrf
Xnr1a5BIUdUHEB3lZ/eoKhCSa9CBOjv4sTFPbR+eVJ0JXkeMb71OJKwifwOvyf9zhcNN2tw8kwDD
neQ0E2kcxEdtLjJhcNr6isHEY6wPuRuVLuflWhgRfXYzAn6g2qcvVPoNUq4+7F8ypVAn/3Nj0mG0
ZPAeVe59dp09VfTfNW19qTTsyGGu1xS54ed/skYmBKFH6eEe91UWgLLZKEJJoiZ2DIeF+1i8vKee
N4z2X5LIhRv6EEdcXrfscxKJAGe/bAKNem8Ix1AvioGhC/hvNgJ0KUV6jU5lOJTLB205TrosSABn
iU/wn1WhNq4LLTHozUhCfs4cLp2iUK8dnKAknOMkcS316khp6Xrv20ZWo5bwWI/IXOiXASWxOy2r
Ax7MRFdUEf4TM3vfCEuJhrRcDKOpkbmUbM7hP7V1PJsCU/k5ULyYgvtTYvOQdnET99cpmj9CALKh
rhxCX0NLTJerJ+KkqKI7yVUujkyUg+Lim6XIuYZuJOM9W/9+T06YYLIxf1eggQwjW76CaFKzs/H5
5DDenCkujwgEJAWMxNWP1qg2rvoc3jcPolWTqTcMeqTYOUk8Zxzqsjj4/hVPVE+2+ayCMXso9y+q
ao3Jce9hMJpVHCMKyPf/kaNzDIG4JC6wz0VPdZMS95yP7e0NqMCWSoN/Rj3rd9+ltnasrBy7B8/q
dq9gaigZZlebv231Rmbfx3+kQfIpRiDWrpz6ime5sS8smyjRV0PfyKoM/v3F8HT0s60rxvf1did8
ys0nBuea+GhBwf29/gi1+DrFDje39BKsx9uv2pAmqloa03ZAjjEh7OhacIYw+EU/aK4DDHbX/7qI
3XDnVe2hbmYmgmYnN1KPpkWct1T3E0y+6MXBonTRIIBWcDJdKHMPszu+BoDWr4ilFmmilNrbajGP
OzN4QLB8mbFxUU9uAIRGbmAlVSRaSPz0QqLKhpXcDgdejErEh5xbyzdb8VJ2+pSWn8PewMNW0Zs1
hASqLtlm5cyA36hILqi/Rw8O99Uo4IRmUAPi5P1AGUi2K5UIkC0IyWuQqN4/K2dUMUkPnwcXJZHh
ydXowPAeszfuqpfpGdLKcDwcJJUqHsF+v3bK7gMEoyVAx6aOI6zSOy+gic/GVWYtOuBis6KvXlan
u77FOXcjYnqHfMiUkki5VpJu6yAi2bfH5+28N5WmYkbI1/XEkm+mcuYOhOf3eZD0nhmAOGMyS2kz
sGq/FAEA7sbKv+Nc9wfX+EeSB8C6aTUPwIOs/rVeSK+LPcq8aOd5dCb8ZCuN7xDVXHetHPLj/BgV
JM4RPJBkSrQahI2KuICgacu516QmPCPCKThOkigpXz5aeFYy6tzxYBYw6QBLGAwb9EoosPhaEteL
u5XFl7q+EdmKHreRnYgR6PBobiJYmSdDRn6iaAKAWlGH+IbgvncYG3EpDujGIeMYlEmOIZfiQna2
3xp8QvfdJKc+JruI18VxRLR/7ipEWvcKKLNlT1UtDAoxyygSKGauN2owXMmDTjNQyM+QpSps6/tr
wV/ejsAaMUc+MWn/hBvkSNn1EDu/zM5rfpNFLyx1zCERByNbp9546h7hxV9eOcQ+KHMbLsE9YNaJ
Xv+Sy3kyrtpnbOINNOnsooQqFWEx/qEdWhZvvzHYPuTQDRroOYVeWxMnKB6aQzYUAJ1YSNLLHBAA
+rvjbnW9FBYyS6MlIi8lAeX2ShxlYshYyi61wAIlK9xsVNxJjKhhC6PTQ8Zh/IVT46CrX2roBOPv
mQ/hwG/R0yelREZX3j1gbOPRZ4k4ti6EAz7BdXgrCHfrxHwm6IBWY70mjc676rNz5IwnI1aRqmmZ
XvzmkKtjKwujgPlZ4U3X93VGeXJwmHv3GeZX63X0R8G4kgwShqYSiinfYLLXAhfSqcCiyLp+WHKb
m25nCmufN9xfJtq9FYD40cZC5nPU6hOEwk7pI3t21eE7hVmctREiMVLSBmv5Uce8Ri3xLTPua+2Q
o30V1S7xDYprKNkhFbAsRvb7OIuMKKyxdtWLq81jxCHiFq+Lc15Tw91PrVwXxNWn9odA/dnijEG9
Pj9aZ9+kD8Z51NPf8XQ8F/5R6Fmc8mfghv8G4z/+e/SAsrFgXo+a2EA3kot1AoecTNg2RVEVr3BQ
x1HCgkJ+QsewEw6CnTRHo3rV8LAxPju/kq9xZ/xfM4PdiU0Fg9zOEXdLN71Q/sl5spNb7ROt8c/P
dQ1l00szwz1Q+DPJW+iRsJTYKaJ14B7fP/alUWI07GsWx49aVnFZYU2FOa8uwj9+kTde7mwwnBxa
Et30XFW289N+dQdsmioJqk0xzp3iEb6J42oMPV150TRv4CQgxxmYi7cUR/zPP1Wu8+xpOeVHoalD
rjWg+5QzC1lhZrBIXILIR7SrR3Oz0q6vA0L1T4U3TJ3WnEEZDuAZIue8TltWrVYcL6ktujUiTvq7
QLYOTcWPAJ2bOVHhh9kGW9o68ua7cpPqSKBmPQ3KbBYyMc4oPoZo+HZewOIJSKTvtQnvU81MIL1p
5A+mGMiz7KmILTnyoEh27YOF2wuHApP48382GKQCssj9ZxldONXn5+fQQ0sXmr5H9ZrhGZf/MAkW
qM352k+Y9dri5YO8UMJfsZ1F+LjT1xoZrZfDQQmUtO39Lt0xjDAsTReLzFRo9sBhjl/RSQ6gy3K/
/Hmdfr+he1WAsSP0SwOfoiLrtFpjJy4B2ahqeyRPlz8m9iWz9+UtHU1wWRSWP82iWHaPoHH3U7AL
IjrC7Retlj1g4BZefFkNo8ABbz1r7SysrPEMyBMe+2ufHjXScnYndQh7mgSTkZvX5JpR3CJ5CrNa
3CGTPdXZ1cixChIRsBbhobqD/a8+ACe/VRbugGTcOwfXdPhf8bv9xYtVQKVZzoKL/Qdk4/+mEiGF
OlY9mSyTkyHhwgcFQf7ky1cy2md8/+QJngkyyGdOzfB8yYciI3aso+XSdLrP4jDDxLb+v1z9U56L
RrmWpWzGDC7ATJPJgH/TO4ygeWKTT29PXwbXIhmPoxwSTLuawsDdnxO1FSTztNKmN31wmqNM147k
pOgPgUM+INIbPT37ha27tF8c09ISVuVTC8EVWGdj7PMCJtsWf30ivJeNShqZndlCXOHZfmlzru86
YCH+vHM4oxwQNDZk7FtMowu7rwiIzV3pz3n6/wJ4P+viVRZBYRlObAN+zBT3tznmfm5hzFEI9xi0
b30d549U6+61vw/W56CG2cpP+SZj4MwnF4yji4kgPHzUhK756KchuNtcw2yls+q3gyd6TlfMRKy2
7JKgQGXrP0ju+SHL49ek0L7srR0z8iBHZcuGJhm8j7fz/+AAOoIyBt26w7Adt3Oo/9E0it9BNRqU
RYq2JYtOtsu61NIzC2g7F653FqZfkJfzLV9xE79yaRp2M6swRP2X3SwDpJPhNvskCb/EuMs05CQE
YLidSvt0veIQZXcHUA95zKKZ9k9zuXa47B5Q/TAqp/3g+bt7c+JC86uuTFmu5EClsZRANb5rBY+Z
Zt0SGi9sBE17bySURsTetqJ0daL1aCXgUO6w2F/HTpl9LGTumKTTOK2lYrfQoN7ceLZ8yqjFPnq4
T4X7BpvAq5UPCV4a1RFuKU5RHzROP5r3Pc3deoHroWTsV9Mxjz8dJ6Fo58qosu1iqV7thvp2iF6/
GJdqHPnj0MlugbIHgXFMhPxfNHPQ+W2IjDY3LsJq2kC+64YigUg8syGskYgyK9cwX9coMzWs7XtB
mMKe/DxPZeNRJfsT+yvIRkqbgHXU8pWzoqJzONvU09whSgcwLlWZZibAdYBAaQ6HhtQjNh0yqyjD
KAzXA6eKaIOlXSBFNNE/90vhqOfihwLeLRZPcGNRHLHMPjbQTZGiYm19plZu3zHjoe55I5G+l1uS
UU8gegVsQDXDGEstKBVSOtYJyJ0xid90ey1+L/TC43AaFielCXwVzQMlnZm8WaHNz2DKz/IW/pgk
Kqh7gPx9cH4YbQgZKzGmLaUImWyBHaZSFLmg3VKda4btuZlu6bkuMPEt3xTKKnSZvQ9fhJuhVRvo
+kmLDN9JErK5LVSg+gkZTgTvK+JWqWdqfK3l6gJpPR/ptf5QdHUNn4qXuqBltxnCYvUsZj57cVPf
yP77nBf/Ro9M+YTIqPZi77rr+ccEQ83DalVavOASgc5G6RSFBn6syhTIdJXScVOgxBreOwIHPv1r
UDpABL8DWDuHknwe1zkhKg4i+o5wevWk9J0VRCU72rJcU7flgpffHCqdPy9KLRiUwzREXqu/OkYy
oJgfCgo5lLAnDrbsdNeLbLI2RkWfV6nqTwi+0hZpVEuXNu3Qc7DI0HHm44yMAbgsUsV3mSv8RwyO
qPzm6d6S6wSjPkqWUUv22G/FU/hcPB/vJRu5LrIDeweZXQ7qLtqthXkALG7KDktBrnVkwnXgoeP1
4s8VLelwP45LIVZh3OHkFr+N7TksS+SgDZNo2/qoP9mGckIL/sA1+lt6iK1qmfLxllYvpBerQHd6
J9oMrQ7AFFpqoMO3X5gfjcBP6h7Z3u5yl60dznKAWP8BRbob87vXueS5kRTEheXTwXEXiH1P3W7q
2A6FrWrQNn6w94/kWRFiOrv2tAcnAhw7wD1L7Qpghua14bJAXAWMvC8rVY/LN/qwa2ysN2VPJg+f
KSPo1uolLNROnsMulXLFkrFOFlPpag6Bdfyyqd22CmtqnSblrNYdSo+9c179LvupwutSNjd+tvhH
9y8AKdZbZ203BtSdpvlPtrJVGqBj9DtJrsywyy/Hn6WwNbkxdElsXbBdRA1fJ6j+Lkdv/Pto95mk
DJmCrnnfWy7S/KPbqvtuLQ1zEw9Xf/chIGtR8Mk5Xh87PNQh3bXuNhjvgj0cJ74rj2cnOe5BZ9Ab
nr+b3m8iSIn/Lod9QyJN5C+u/xqX29XuCSMPb3kX4JfqnsD1p2je7yYi2nU7JamUZ36CdeQARb6Y
vDkQ4bS1Nhn/QUWYORGoA7W1q9xG2T2XGl8WrCcWavatkwER/Pp+nGuxc6v0xmR6du6TJ5uYX9+v
zZCbCJuvYszSQg8mlDXUO64hT85SGEgX7dDUuQ7qIYRTaKUhLjcG7+fd5UUsoNlRRdsl0WjfB01Q
UUy4Puq8j/bIqvTbpjwV88OC/3u24FavllXvhEhJEPwO6sQRZ/jr6DDobb6Xtp5IDu7wMmYzmOfT
agrZPWJiKQ26Fwc8IXDbrJ8RnJ3xDG4P5Vza/lWD/dUKwlLgz1Oy4mtLARiJ/0hWqQI20LHxikK/
dM6ObJbm+jTHMrpNkwubYJu2wBGzEsT02+YZcyimdvoyi48dRPp53pCidg1Hskanwx9Acj38G74Z
1968vS4pXM6IqN9dH+nY+0PQdiNdrnsnBmYVQ+36YDkZZVxP0RlL547UIPLf3f+0xuZzQZfY19Qt
hQUz5mY35fqWI8yCMNhXDgpbf7LbvYluu02UHQffKqDmr8/zl05hR/S/SsiPFgOwot3o8rv1Au7c
oTX63qiO8lMr0dXDaIXTPDNQrquJ5fizgJOy4UPb0Z8UIM2iiUqDp4vR8bAt8USVzULJ9mH6+OaR
jU/A/AXfKcxYj78JuSXjpaE3ytu2+ncq0uN7kXfps4lsTevrX9jxa1qQtALzAaL8U77XnLx9xSab
HChKsII5yv08yi+9GBIWx7PiQYzEdsZihfu0qcCi4t5RrAjlqcKiO9Ab+6vhE8TYAXnu8Fl0CyHV
ef1FB0MDQtFYpTy/dnRfL0rzsSSqleRA/ZIyvWcMTtJ+0fauzyiI/V8dfdxpDpM81Ckv0sk5fKn8
pbh/XNhczm5ql07Sbn6e1yaV3pq1lE6hFzqUA+vhE25Q7zU0f3mH+fbYpbl5xk7Sj9ntcumdQC2k
FdWYaz1DeEOsgBY1hmEg6k5v6ZXWm9C8VnhrtaetrctjACD1/MAg853hjhLS+GADsxZql4klZRcu
NRi3JSQQmKqZXGtiwwU3Je7FVHIAbHovBbRv4Pr/1b5UPOWEqzv1ldAhPmrAEtnkCXUnWExQVcFa
5S7xxjysr0zIII7uCgNwI3I5+mo/oVDqjKWLHFCGdBdQTgsfYaDtLCVx7QMFx/re5g8c0g1hq22U
cSPy9a6+XNX/O/jkYo9HmHdgOAoaTcQGB/3MMnvXED+eAwAHSMdhkELZfgZObfOWSBbEKeA8ZeEN
CN/ik1yMovHfXqrq6aS2p/VtjbInhCi4UUkZpEmeEhxeuIKWmoyYn4lHwaL7R0bf6VDxS22FZHcD
1jIPtPtz/S9H+xO6XWBgyuZthSFOy7wj0NcWtV0hU6eTJxScgUPPgdtcGS1KCl8Ak6bmzDSA+qlm
Ap8gltC0O6PlsbSXpu+WaRzq4jhfgnk4vDXpV+4EWMAcMlhcO207njHf97Jy1lBNLAgOlUwEvO5d
x2Sk/07vc0oRM858zJPbzF1mrVocV3VVv3uIQ2dsOkApAgv4m1PQodajk+FqhkYuDKcAntLR2qk3
r+IQERY5fOKEdXYxcURYCSAcstRtW/QDMjPUDI3DgyIvj7ksUsWs549qxe5fLSwUP9t8Rw6l3RII
SQKdPjb2uJ29um8Q6tZcD183nP/1sZruo9NUcmc991/MEE2Yju7c/UvI0Dz+pJ8BqNY3I83ClLPL
dZ1ca9s/CcVwrKNV2I4oFnRcb0Am3uW7sDPEflSC+n7/PJ2vWYhFfhLjThhbdVlL2DP2r4L3C/UH
9sTMoJigLwiY6E8bykPeqWsuRXqAjXS0XeBCii7DcuzD1oE+f1t/SN+3IART+Rm/OjyMV7jTuLkL
l2qLfCoUvUP+yhg4FX7n+eLKP9bAEnyIskNRi/DwskCZ9cyVguhmD+YZW4WlZwR3F9cN3K938Gn2
9Ss78U7nVREzHwf32GavJNayRIvBe7HNjTpx37O6PzIMW4z58xmRuPenJ43+DajEICsPvDH7D6TE
Vrrp4SdMwE1d2KVdggAWaZZjcBCnQ3EN//WEOl2tdmzZ+9fyrtQOUvVFEG3nlelWQyY3+pThx9/P
xkDp117/JVmTY2sADsY2z3e4er2/ReOpp93hTPeQ/u5Py8NtVOCzoKqhm4KbFRbnDVhkBw7lz2Mq
AqKSgbWoyTzS5nxV9V9EPUXK8nRbkYqLdFOEe/PofAKzXNazRWCELKifMK1J3WEYOxu1XEDmGADA
xTfqt/4Wd/FH/s31xvg9HQxrsfjxCec6wYm+TYFPUsSOGVFxFIpWKIynQlZogWSM5TEaI/Y2u3vo
FlRSNvR4O5DzS9aWxC71Hm48cgACJQaW8cCXBGZc89QDjaiKLAaka0SJ7FUEtWRe5tVszfe29znD
jne3MhcZL4iy1jyAWkXEKAtpZ8kvZZdwAFFzSafuPlbwcScLNwFcgyML/6umD/pwdCXniTCmQ8wB
dpBCMVixZ2GKa11VOPiBIq06ZXc7+IqD7/fRuRh2qOIqyYC3qwZ7NAKynzJX0GfLcZakbXdvZzJC
IMlNzsw4FH1ji7qQeWuIYa9daqNLdZJyhpXHyvLlqGd+7SSxAtH3Gu4rmnVSjhw2qzP0fqIbkToU
DyFkn6ckjrFPdsbcFX5Wk+/29IwCOweJI6/qApEYI/YMalc8LENfE7WV432npLkGrK1FDOF5g7jp
3ze0QXEcNBcsxEnNGKM6Z5eK09SNxHv1UbbN6XKtP89CD3KUyRAANucyUHNPFTvVcwlfE3bJVWRq
HHEen2ZK6MuFZcJvAHdWKOkRduXettpXRn/BnGZZ1qTtxmfGl+CTZu5m6gc0YbflzaBMbCesKyDF
9u7lDN15bbTsUqNNVcJYPAtpg6liO53s8mUCZvBz3f7seKrCuaw1iUVwvDb3Tk0dGx41dkt7VsQj
kTjexDs5DM6xqSCCx6u4Mth3pxiozvqnazq84bO2KXa2b4kNOJbaQj68XXr5Grdn1T0+CspQwzda
dlVoFkuQsWMA5ELwXB/VAGtz4PnRopZJDcZMuWMJuC2ZKEBs/cupRCDkuFvtmusGZ0fGNjn0FRir
AJt2+NbF/VgIoMIHwH+eRm1PYistum5w+E5YpItAaDlSTgKsxiO9owyiGJOTGZq1GvS1w738e2jx
h1S/kPyub7OJTkPcxj+8oVEZjK+/NE5Me1ZLqEATgZf4E9qPN/Hqc3n36TcMy8JCgwzxDnx/HiNP
PdUwr7spEqweoFzF4mnrnhueBnJKogeC7W8X1uGY2N8sd2fNHhK+fRoVa2G4wOLOUgmS05aUtoH0
biyXCJwKa4nKx2AIeJWwy985oUR6ruzp3QpHwybG8VeuVSL2zFISZWPD4e0UPiJIlR+IJKxdxL03
pawiPxZa/prco+xfCz/NOgeTS80tMzzbuTvZ+nlVmeYb7312UMCsBv7FSkKx5HWYsi8pImppOCHP
5syQZBKFEubLf0meSapk0pGKN7UTw6sx3/SA7bEmZCvltucs4pdGn5gnDqdLYDpJy6L0wy5c3tIf
uGpjKR5Ojhd9ZVxoejK+mcZCrQHwRdIYbqBukFoQ3BAaRiwoDt4kwpudtHG3eXUsdZHfO3wMixl+
t6BtXnJLAyqUMISl4uuTkI/oz+yrX3IYvohLsNjm0GLawn4bimMDCaT4wAyLDiSKgU9sELvHKg51
VIj/P7n0rspJs2BZ6akG7gxnpNCFQEgmZdcxjM6lT+PkjkDC+bpQUyLJg+/pahiKl/6EwraztYlF
CaI/oQPMWqTm3uq/9AwHvlg2B+X0qTQuu3z0ZBRdSOttB2PpM+6/XTFD4w/Oph4EWEHoF3hxTTvh
VUnN3TWiUQ/yqKO6NSuWRRtDtILUejW9oSs0PEZXkeLRtBWtlNEzSszvbtCB62n9uGmN2KvFlPIq
J2ZJ/iHk+Jq9UT1muMadcrB/vclQpS0spjcHcjo+6Lf3LGcLw4nVo2NhN7CYImRld609ZakDJyNd
lmJyCGoA+MOw+kZew5p3zRCe/HEUe9sLSLpGRM4/OsUCfn+BNEjK5rVsTeWs1PvvPcwxOP/8xgcv
w3XRNUXKpVd2cF1TbDXhbUGw/be0NaeOjM8Ee6Vrrricd3UPinGHsJNz35K2gTBpZTNKF3OPO7We
46lhHvJcozUi4wJnv5p5f0a1syO1tY54FRESj7vDYNf9rrqK2zdWDAP0HytUh2AlzkkuHOjuLckq
TNcCDSkXVzCvogEneAu8DTxuKa+yanpSOjABGTcTpAgEmhQv9mmyfc3GIHQkiKaAuWEsPOjRb0fI
cWcy5SRdlISBH6El+HVOPw0F/weBTp4LhCPnoQSzROvFIMykqMgMDRVXXYrmzyUxzyK/wddKbkN3
7snYn8vUauISZCrgOH8fqhtCw8eU2GPOcAp4eNx56bS+W8zxDmX08jdZvsxDBSNeSTplIqJk03q6
jd4e5o04cXLeMMLHjt1w8UqPmcSBMLYQkEqUe1aZtB1dz2xXm1/X8+5vR0lRIMKiF9YhQ7XfFwjh
n4t/J1W64OekgM4TxreiFXpruMKIQjUG0KZhEg+q81wIDzXsC85PgPbeflYov4neTX7/ph5xLos9
8yZJqINJJLDe+/HAKChkgFBvo9g+PYISlx/e4t6t6wqUxCJsx35BB5rwGtRWlVr1rKMF0/Ha1SEx
utIHP7P68s1GUKmEmxgY1+0J1kk4Zfbbrulws0Fk/wTQ2eV7K94JP3XDCr4vchKGMVQhKRd3Q21I
W4Q9GAKCgIr5n/OJ/PWpHt1vPl6P0puL/CZqp070rS7U1+2Q7/zOeyaqNXZCTS+sgPsYTOsC/6J4
vr/mER96Fg7mjT4peJG4lz8KzCkhDHN8fW2MBVcJQTlPtPzhiZp/VOhMb6eVjx9zX2T6eHwnvCPN
V7IaDDWXSsFdwef25iCHLIJbngmrm67fIQeAuVolObL1pdGuvG2riq+gJCAx26nWYnKJj0jQb6ws
ExrujAnv7KLduQbFKcWlSIh9+6NR+YYLOz+n9l2cnjWnKmSE4TA+r6vnr2srb+S7Ve5N8JMdVOYr
Oxt0bC5KFggUP0ZAO/T7inws3nBfQb+NNJxK7FteNbrSwqBMvjhJN+UDtiAbBDebvRFlL7sKMnOZ
ZVTyysdmp2z/yvTZwtuEW+kCE9LY+EgxL0Adc7o+BnSAoOEiUHqUN48XaZ7FT31UYfSlcgPGfH+T
rKfpqXZfxRligvIbcEmbgElnPB9X6F+kl7DcN17vuJm0srihB8R4y8q4rVyTHJ4x9KL636fOuUHY
M7wjOZujISyHthPgjmUAqi+vArWHstLfBn5CgGhl/GJmbTFt5eX9Cw4FrZgWk2+fqzANjOcTkFIG
ecptgJMLfOcgIB60KR0I5fR7jMlWx0380I1q3U9268IWVMCs4voZEpKct9ZNY+cbSd/+PPrrvEl7
E8Z6wk1Ol0z1VZ/rxxVl9XJ4gJdYrKC+387t5m51E+CU40HbzzIdmwu955aaAh/xcETurkSYWoUN
nYHkbPGn6SmzSs7riwzwjOVoUbob/qW/mSKsiyArWSA02fW/BKaTmREz/SIfLM+cjlJVFzw0CmY0
h2QpfQ8YP0nIDhcDSwbrYOXYidvLV0svtqQIgI7+uFMg3fEjOCZAgsCWSjafotkJPzdesvQnaR5q
ENo1TKjc3u1dJNQ/PonwGlBEWbqLG94XwkeVvRUplUZlqkeLy8BtJiq1/3umS1/gku2VAaCXxnQy
SNJOAypOfTCGtU2FY7Q4BKCRXwOBlUrkHlBbYuYTJvZZg31vpBjPg/lmiyob6L8POqodP7w4e5nW
9kg90q122Fraeq7JqXHWuQv7tWnbGS5tuM/jM4IrJ0nJXstLn1A0LXB4XQN7PXPx5IAJX+zVRjJ8
2fsfQfghS3NsGQNa+LYDw9mSS3JYTfCUWKGGVg+txb0ihcrkQnRT3n8KFUbXzjJYQ3YXWX+DheDu
e0u1UNdiIMR0Ffpgd7Gdr6etgaBIhwmxnbFMRP3K2ZdwlaalNFgAmcNk6rvcMlO+5ramRTUOPuHY
duGgNKQW0KrNzb4241qIxvbAyLXI6i2K4FOuNjkyvR44MrU+KgeBlBALjAJP3FA5O/j3CFnoAtrV
saaG+Q53Sa371XM7gayORJyMfu/ATaJq2kBqNz5hMuVYoqKpmcv8BF4utpW2bgYqn5IbhBNF86pu
UgY8DzXqVmNJd77MrObXWQ1NJxutn8zDOuqN+I0Rs6RYt2hjbVnd3dVDUW4G8hTpxSzvFaql5Hjv
tFVI4wX80HaRkVNoIQ7DNbYQ2XOIQkuQXdDGG6Mqdr0wMInsM+5fRczTX/sG5HylMs3EPZt6kONh
C37VKt4Xe5iyTJlUHdUPBzJzaxjkpalQSxDy6kP1B6ownHg2HzO+GxiSCkHebtsS/tbiLWDjKvYu
5x+sw1mD91+U7kkcjpZwkHibDE6kVoH/PeJJs8cSWedV4dHmCowR7TRDA8VSWyLVoI7R1T7Uv0Gq
XyB2EcP9l7Ekw2Sh8Aa3knWmc03PRFNsO+IgLpj6f/DL6t/F3TXznefOfkwyOzCMi+NceilLCMfI
qDCUnbC6mpHT6a25zXGDZQkJnmWXxgZaVIuTLWzx928MuQ3nk2migW0QNEG6xV+o82YmlJhaZbbb
Af2EA8JCjPrtlBjdK7B7yHbfnlwF5DqdtWy8gwpCyEzHv9I/atzkhA5EnGwOFxDLOSF7J/zV2xlj
Kma1S2/JbP7qPMBarP/u8oymb5BDhmpR6xVlk3deJDkmV+S9/ZUfXzWOErtOKNUEtPFOaqOgORtN
NYpRDMyuMCVKpo7tiYxwX06FV7lkAKPcpRdItoZWi6WVotqZ/1wmKcw+RAzTRIJpGhPekidcdamm
NPZ6emBD2clMuXA/KZ/QxsBSWmVD06emeh+I0C276Zn+6XVJqJdGiFYLMjgYvHFk23xPfHwO2kwY
mJUxzo9NNsJIWcQIHyDfCF+GIH29oiQTNcHdD7WJcsc+STzdP6wBdwPXcQKceyejieEvGyj1z3bK
6rUsKMDTSoScUIXAR/UpKcj71Y9eCKoI9K1Uh4Di2gMqCX3Dzxh1twtm2VQp8G8JhrTStzs6pWus
c6bufGQJUVkHNs8XossR1zgaHp/Dv2wBgN6OicWTrWu6IHIUk6goHyEyKY7w+o8inwubdy8utRzp
pmCo7PWv/YxRpSXwDIhjUygo38ZznIOppdGMPD9kFitxMaM0i8XaWvpsv97B39lOj/JiuDtqrTle
P/gVuZYodeYis4l/qNmOjyMu3A4T3mb7cEu2Z6eUt0HGWUlNlM9O5fSVedkFbJDPFn6QS6vF6uzA
4FP6V/38/FkH+v+z7+qcP1etw8oEoavwAQloinxkgERZlLmNglgaE1KpSKS+zavA3hSH1QtpHvEL
5UVFJCQFnXDcxtO8jMxRfYdA1f4K1FYrxAlK8w4NlSnWuUcNt58KI64bM6zyojr6abHtbMa67da3
JPF1TbYHCjkOm/DfKx8SAZTWk/lD45ggMf8CpRaU/85/dgBxPLzvEld/ZUmed3GFMw50FARJ9vao
9uW+/6h07frWPEyAX7r4SuMMo1jJt8BFzMujbJaJ5AxUcfMnVLbJvDwK0HdILCLfVbZxuoRNzeTq
GwY2uOsEfu31+49VKzY6FRsxmakNvl0yhZ1M4RNIy7+FrmMqwMcl8YiBmhnbrkTMW0yy5Fgukq8o
fieFGXsHRwBobP6mrhs0zvqWSasjRhnUUgfTBUSCuCgXLBhheSstXC2vxXBOmlHZ+kPDd+FX9KHp
6L6KXOCLC52f7skP8wCN7zrRkbyDmbj1bS+5xk/rU1Snl12gFxCQq/jCn0OjI2KKQXnuGn6+Ty9l
L5RVOoefAuPUr0DRdp0PiRb6iOrKFehKInmft9rJ+pzyjC9ayu3/d0yyvlOUwp8+0cZZz2IZeGQa
cymOvEA8YrW+1HaSdMnPiXzUh8QHyY2ZIwC9tJW65eqw03YVya10PQwMEK9QXK7ZrEajnxKiHDwc
tAqkE3xaXj8T4HIXQ67Ijbk6aPnSLlr2n2ihrKNa+AAdQskAOs8TlSMOs40J0zvLIyUmB77HvYwl
f0Tp1kWNyOmpAcYzwFGjjquoWFtmH0PqsmrmFLBUJsEYcS8TcaZyUsiwudGx61GFCJ15f/FfStyw
BqxXRrKdatb2A0SttDhriGaSpD+2DGPeSaJyEQ/CLZsuysg+uphAUxLFlrvFB8iVZrYKyoArjZs1
DeMsUJ2fqi27gk52Sl/nvtUa/fcIEbdtEUzE80QhWc3Nk4BFv1mnOrCEvfWfOtNJLRsdib5fu7vm
2SrHo9o4RXt37RVAOLIy5p3eCYQwXaI1SGH+jMkGu33YulyZ5LzpKpdazHoCe6XIMBeN2VxVDLDP
eqXFOj90Vri7ok07NNEJPichw5+J+1m2yKXomVZge9hfB29ybIxSQQ7pIj13UDIJWJrW5KNpM3Ni
aAyN1JjEx+0gOulf813hnCYItoEUysbhpTYJf76PlzUnxwFK8D5qpHcLJguJGw72zjMCMthoz1oU
uA3VIgBp6nffXNND16uJT3ZU1P+MPgqXIxMsALde+8jgjUk+uQ7Vva5mF4zk8zcJr7L2fheQY5tS
1/1wY4sv6gOwZwXSw010R5LUA4EB/VZOI/+eqMJngT3z0wgff2JcWuO1fTBdw7soWJ8GmrMjGUGh
gmEIURXGCOMo3CyHxF7Cdd+9gXn7AqE12golNnuoLwNkp2i9JLsqHdLqPjRdh8oDHKFiULcEcK/s
XqchJ/wdCrQYHnxMeBLip0O+7uRfYg7olhAw9vmQfpyKvxLi4RXABR1Lky6RlIz6gn+gSnaxiwPR
OZBk0mDQ2hNkLU3TQrf+kSaWu/w06szVFYSO761p0R2F4awalsMzcwKHmBFrhBgaRXpYvaNfH/Qx
Nx+lnpcAMYH/hx9z2g/doMGc3X9UQwNZmt2fb9rmiR1tqVnaqyLPWHC1zOFtq8djLMweM0/aJ11a
pltYuqLDxxIzuJmQuO4AgwwtYbIc1MFMS/s+3tAb1EEaaAEWXBPmzmsTk0YcoEnYGmoUH2STEf0/
6wvMgqIqpE3PHOHREkmP1g0X3I7XyI4szoOhqgKNiMsoGTBONKeGnsmpK1JWVmxrgLUM3gNwb3vU
5YR244OWapj5uScFWAZh45Kz5VHqgW1CzHP5UP6G4rMiaZIecl9vmPZoMuZE0MqZooI3C/u6dS6w
62pOv18khdh034IjdwyHLiFqUdQG0qiM3X/0LG3xFepXzRq8tXk26JTzww9Ncogy8yvvp0v61A0A
oBKbOdkIQYrrQ3fzlRrGLr9qCm+XOaVi7u+vKBmEgVPprNTTk4lWQntGGXtEnQszrL7wwGJnHQro
DuFPoVC1zl7yT9Upmt9y0qqUktovH/Rd+xYHfJIpTA6j8KS/Mzk/mKTzV0WTvOTpgGKKEaiBakMG
wCAhLLpkQS0GFDb/A5fCEOICBcfAam9ciGUnJdR1I9RnEEvQ1zqlhWRaCIZOT3iA7bFIgh38y6B+
ZzVxOXCpsZgx6gZbthGW+TCSPh750GvY9fl7rFI8N17ZiBfapvZjQD4JXOtiF6rKMtTabTy2Adfu
GimK1ku/zHWQ3t4y70Mv6TafL99coeQWh+F5/xNk5Ucgdg0Xp3g8u2CLFQxlts8OcRTrBComHj5k
RV/7B/vT8aMy50SaAfyqsxjnORDt1l+2fq3aY1azE26dEhi3ZIe0TB9AXLWzKAhQL524b0PZmcEw
OvWBNCkeWGnERJN84SpBO7efzJhdYQd4lnVu9//dV4YGkhkLbT3/tUUF64o56akVv+oSOAx12lXy
JtUPp4oR1REz0F7qWqPuONJ4uMReFR55UdroBvETAqPHKDK04ui/LqH5Y6/e2zAY/TtSuGIK3UkY
kqRqHiAfDmsccuRlDgLQF6ME/f16Y79yH4a7dNW8OvmffUjhg5S0Mxa6Queo7ncpUkTUeSJmNpBQ
dq9vrU3td2KwGl7QNpjPaHNK3cO7wD2yfBVqRWxvuI4hf3EEGVVyjBurOoRIcak9M/7uGk9bB2je
CfasQSa6uFLiWLpZysmFmCh9mggRXs/RnEW7qZwZOdYTZxow97I2CAJK9AA/VIHahNPezp49ZG86
/zE7Ry1p8pD3DjSubX+3qaIbTg2qi5yhH9Q3aD/ryr8/xnMDQfvtg0a1xNt0Vgtnln/zdxNoWSVw
roEiBRLYjXw106T/DnIm8WSAWtrd6tKXzEX939zLEWFAbqDpXzMtiH/dg3hNQ3vmuyeRheFCG0dV
L+rOQI/IYMgA6vG27/Bm/lA6UwpCHednH4AJjqFutW55c1e6LqCxjDmdUFVG0sbL+7pN2nYW4fov
wSgSdkK/FmXRynNB5el3wHz1nd6jP8UQ7gTfwbXC+DlnWX2QInkl6CRjd9ust2BtkAwamocMZh/j
caxx2uTiJDE/eeqmDZIINpTntaZXq3VL2ekq1Cl9maH3ZovKtOKYmR19A3xVJozK5/FBh+biuc1Y
SZxeEkd8eopQkuFNeIdTDZ9Id76F+DzIDNBymU+QcHN0OwGs2ZUgC2V1JkcP+8ht7dEXSPhij8iq
5yWLy3CtFG114kK/blqqJrVgK5PYN9XDQ9OlykzzCGuYyv8OgywDofv4zQ799eBKuiUrPpF4lnVT
zQ6L8sc0ioYvOc9z6V3FSjGb+tz3wEv+XIhxjfUsi0crWilQyux7RWqabbqkAg59SzV8xt4HJ1/g
FuKXTRmNBNz3t1y5MAHteXP2eg1uyZkUEHUBap+bKkYfFszYiuEsuxsQ5QlNotiTINsX2N6cZROH
C4myYN1RH7qasBHa61qs74nocEXGw2ME182pV7OMP6M8eS5TfrSj8zNr6PnAK56cUQjtCYUUIlZ+
9YEs7sp5dPDzBIt9NbLaUKN/5v4tgPxBo3wdrGhbSzy5uFRscXlrsoz2jcZ9zcn56YXvqPK1+Xh6
ngVvJ6ijWV2S26elBtMzd1ohZeE0Az7DTeITVsku+MoroQkhefIoErM1rPFrGichMnBdfe420hDR
vXmS3WgsBKTIqpQCwtYcTSyaT8UnOea8n4h88a18vDTmH1gpSl+mkiVHpIlzhWhCVnyOudSWoe0s
d9AP4esGpKfCYygdHc/eVxSVEwPpZCTybMbIIqfRikyqA3TbrSUVeb8lxrN82BLTUfhn3nxnRvpC
VS5NaqqZromnVWvDq1rz2yvlz45RXvKxj8qlKlWSnG6Gkct40eS7uEjNhgHmYLl/vE8akG1ZKFMm
ox66qZq+Id4g+RLbdhDQXll9qr5wwyM7OtQidnXSXE48GhNadrvJzmGfCafvNuc+zcx8FMaqCGpg
b4Ru4g6AfEboWYboJAmpK9J+yu/GmE/yuBbG64geX2FTCxosRoITIBurGmMBlfgt26U+GJnjEFF6
ilFGgmwGrIxuRpsYdpMVp4JKAJ1/hzaWd86oIKvl6VPF5IuOi9NAZdNVFLTNkPzGfxdKLcES5iIE
mIzLjfBtIOpEWoKY2rq4AeMNHUYL1ulbC9jDc/hX0aTi4zYX2lLE9U2VfcdOZ/FlMTWy3D7EIRX8
QHwdCrBMgLq652PzacTcPy3BisWmIW5UJQK7ZPkHQ8FxjGnXzYzSD+dJmmdrcxBanjogs3nPkE+O
sDJz0YONeZbmSQ4GvaYN581A35TODITnwH41D/pG9nyqbSvHBoRlhbCdkldA+qijKYWYqb74qZEt
v7AaW9ohVVDP1sf4mp5hktl99cp9oKCcu8BLVhMJ4x9Vn2ytBTZrLgS92/VE1yRad8I0CemuRzmC
Wd7AWfP8KKwgaUB4nCTr3rAxSLjRMk3IvPD7/5q+eKNHRg3pP1S0uOMdWgPTnZHZb/3JWgZekY7r
86pjsjgwnRoKXkHxVQj1jDV0gb/zxEiy85hM/y8rpYp4bSXQ6MaZbDH5yvuZQMsaILrpvk6ZGrLM
psUVIWebi/LKUJA/vgECLQWrxxEECf40SmFLR9P1mQb8QKyVPRK9CcBr1Za1WVSVuuI2wq2YgtLU
ZcNNpIxYivtWNs3gv2NTP22VDM4NUR12aj+7apwOj0nEYUGTSI8WbwA/0WF0kpUCdU5cWWbZDKoM
xqWM6LW3HlHVj51SaGKL1Cn/5MMoh3KoO0u32XKEcBpKD4ivV5cvTnr9sj8/ESObrsRxWIXj7SJP
6DeTvVxe5cHX5Gqt/OHahw+BrbyJKTr7ouwGhmoQ9EFOI7UXD8Ww6tdtaJHZb21MZ7cZuDrqv8K6
eZp9RuAgIivFdHbD2/LkDd8NU6Hs8pudTmKkYIbWLIgsLAtdISwnGZAed7cy4Mb7qSmcE/CYricz
Isa/6uh0lgvlGbLH43JkOkZCIWRixIcdBkou04ZhcbONAvJ0vvDJNuZCu4Evycy200OKYHOnXBZe
auHcpfNGAfOTw6NDxq0VntVf4eWFICNxzkCO+/22vYEYwslnk24ZMQj1JQD3uvzdQ3sULO5eNAOu
eRgx0iKiZWXXrPVIpntRULIKkmpcitAuuL7VqDvXGqaix5xrWD9zlwRF6bwbmzN1HQgaEturspW1
V0QfvV03dHPe96dtHZl69aWlZ8P+DkFz788r+32gE4SVJigjX5acdCCD8KhiaOPg9NoV1VvHYEvy
dEnb8mXOulEQ45F+uYMSXZKNwTX0CxWxDsugQc7s0NugJX8GtJFm1nikw4+gUePS/i7H2eCpxJ1g
iEbWngfyyLZmz0lgCiIgm4vlmTloSAR0YnFplLSoRxCfsZU+y4ef4e1BzQsyhqJKBwnVd7Ofq8u8
YcaYY8q9GkY1h2mZnZDvlOvr2zbWP1CBm2nWm/lWmwcEPs5aM8tRs//2vQG/FdCw4eypA7zyy2xB
JmbUVu4zE8J+LQgddzWt3istVErWNAhnslXMzEtRuekm+kkvMJCtmrNOu0X5lomQaizwsUcKfbvB
IEEmZ2RfTuoPOglxNfUv/aa0YyniwCUIZrXxrtxMrFz9H3b3keP9UsAODg/7rL4gGd+omVoN9Py+
AY+jB0zfP3Tse0b0sCW+gy8B4ZctIyYot3E9X2r24YJV+mpATtlfDDYHMnAfz5oXz6lB6Px1rLfK
FeYfrFLj4mQekVCETurkA6VNGW9glvlCJJGjGSO9+X/EzUiGf0FUetC+EkAAjlGuXDT+jo57M5aW
cRqYC38NYxBV8z6rQ3PLgBiucKpZJ34Q+8AIvDS2X2BkfXNuGzirxcBiU48SnsbJHa9+gsLdZu8P
TLakZDmBF4SCADCa3QWM4kaGgFxDJaVEITNig14mG00HA/ttwwfyXNCteJBU2046hkO6gdfFXYEv
9a2giZ8IZK8cwzHeT12oQR9exXyJPvy3AuJKzO1QF5+H8dWe7w9rm/AtmcC0o14fcCFp6QagVlds
Fya6Fr2haA2lE+z1fUrvGUpyQLEzRrcStGxmOyzW+GwipzBrOQ238NuR91Myg2AOBdtZBkRYRxpm
BUmkZRhHwJ0IDQt9Qds7obUH73vX5fES4WqPyrBNy0qpLaSDe0D88Pt9PisnJZvMzOZvkmlS7Jve
dU3okE2pICvpFqxpRspRUH/7XiK1t6FsYl1nH5knzmrIkemS0zD6W8JiuBzumrmGdCFdhzLPemJh
8r4KTvRv09pDHLLRAAOkewAjR0wha85NE1NrgQYO6HMsZqy27Zp5mSyhUsAeLHmoJSKBdykcDz+l
uikL/9D8QyBeQw4seb8Gtai7Ua12QRQ7fhchoZ6eGmuZt1mHd6s9MJjW1Wl2PTgEN6l/SwXzwakb
SmGLgeRV7vBa+FPEZNg8D7fVjeNbtdNsKPrVphF5MqkTIyGtcpvDO+M5r+eYTNxp0UXUP1NPTqR3
WJL8/1mTPzlTLni4L40ffe6sNa54B2CEqG0IvGSaW/acA1Bh759JSnCIgYpFNDS3ZqdvHDj54ZOe
3X/c3T8JIKd3rDfcS5eetl2f/gJyMhLSjEG5N+X11E+zOJemxGtkqx0sIPsGOUOZW4r0v7GP9NHv
t8AAnMTnVOyAG2CwG0aY03qECTME5Qu8CgGW8zrErsFSICUg/X3V/0fgiWXewI3Tm052zwMQ1yKd
TNITRAaA4/LEPsNKHGrItO/cjYBpskCkkQnGd1ke4VHAdEbE8V00U7KFjLsd7n8pzC3xtOGyEfDU
uWSh0yeBlyI+i8JElMpt8FcPDAwxYR19nyJObaaRUr8tJdR1OIR4sWcG0+Vt3cTVFyPYWfIjSdbE
AskEmcpZVKrMq+HddZyKZhnUfCo2xuDWmYI5SIViahvd3pcnfw78JxxN85OqJghl82V+ScpuahvN
1FbCDOlWk5DDHDa0rpQUMy0zTz/5XCtGZCzqfzysNCdFHYAnt9HmOjsSm9ds1MF/BPuJFqI1/YVG
MzhTbwWDt+LQx603C9bP8gdWyrRi6Bw85TacJyJbydJuHS6xyl8SYjpHpI7mEmeZJakYEQ0Dspwg
VADpVP3oMQVH50wsosMCXxsAktrO300HvLGdDOEKC5v4NuIRJqNXcPsuPdTU8E+6Y6G/yDVMCWIo
5Hq2RrHRgdKjazr+4U2c6Uv8k/6OVUuwb2dbCDYHmzWO70fUD13/b8g4emQwc5fspj2LrXbDQPii
4uFt0HySDqZcpvXebSeaqlKarZyYrKQXrjnU4Guj3bAy1FVZyZcZhRh9L2P4YywA7h+ZftnaYpMn
U/+34CGjccmHtYh4+9Skihg0fqH7g/KRt7Ad0HBMrwbIwfKe5ERT2whpZe3cK36UtR5ClSci9MCe
M97ENEJQJqReAJ2uA+68p1TVWvHQKVwUwnBMtbbNF1G7opWhibDCttzv9HqHWWfStu7Nm5ku2LF8
BaxC/BY3VrNVQP9eDMbsGPCSTytSZd58LG2trksCTk1dJ6xBZc7q4Ikit2HLli3qbYq+dOfNyW4W
uOPMB13Z295smIvanGGsUoQ6nj1aH66KiJFwUI4DVFlBfMm8u1ZmW5rsOxKnGrP24KJ6pbMYyTln
ZbQsre3hRyNBV5WFH33rktYQsfz+bFumI1weJTDF+4UbLzl0fFKNDA05vjSLiauhEucWxdw/ZX6L
G1Zm1yIh5gTKAx+IHi9BZtB8SSu+/no2qvJc8bZYK2vExKae4D+gUDtr6bUF/i/jO2BFDmxU1yND
AH5aGMUln9C7l6O6seubfaKcWtS28zbp+PZJOe9nyLuOYCCZXhZ0BCH2sxdowgorT59w1xt4uO5K
MdE3qoZPIUgIyJaRotZvmXrvhB7iDkYpcxkvwwM1idMw18V9sKJWyz89tUw1LeIlqtKiWwgrCmLD
cX5/eB/VModdYmc38u5CzMuugm5q2GYREtDw4jwIFPzUlNS2+GMhj05wCUHtXrrYBi03YeobTs5u
+m25E+v9RP5lYZ51XgwmonsGBv1gi3Rvw8t5MBFP8Dhk5ggyQv0/2godIvPpMm5PK/po8yiTVwbu
EhsJpYjVgfi43zKTQBGT4aSJdYgB2e0E7eeoNZO84mbbcJl0DYvF0RdM1O5rFJ2H7mn1ymV7aElu
o9p5+CgX201y1jfEnId++cL86TtZErVxX4iadQl7ME92mdsvyuzRwG50UttaztLikA1BmuYjtuIo
BwugjCOjH2cY2KD1MQBEkHIl3ZLpZmXA6tzNFAwak1tePfSwIlg4n60qI875IndFIi6AWnh2bowp
NG06PPbhp2Z0tDAm5MhMIfkRLHKYoJ5ph+dMs7AYd9XbUdJDSeeBSBganiKV2A/ICzwpeatOQn4V
fhwKhHc20ObU1HAp29F7SranywLmrZIOORAhXOH8BbeISiHoSnBuJoi0/8HB7eBY09rc2wtHM7U+
HokuyUkx78KatdO13i1O08unpu3oUeJooNp+AHzOIR6Hv7SSNHgdSkyPAprzxq8zDsJOaUKuLBA9
s9ZvQ84kDMqo1ZKJ8q5zZI2E9FII+VyRsQI80pmiQ8ezX8aDiFJswHCtx/83/sa7Hux3//52YGuB
bamIp4IlZmWVbV0umXOdldPxAzQbzzDF1JxmIbyx8RcCjhH58EaDZbXMLiOALqEgvMNDrw5euum1
QKPC4fud8528R4vP2UWEle0mv0+fvb70ktDpNIy1j/btvDelVDyxL4Y5yFAo4cnaTi4Onpvexa+F
mubkTq6mkQ5yEr2FAVX7LhnCkm6xX9jrc7Zpg+3v26M3e3Pi6gLTIhW+ZpNqxHpd2kca6nr53M+f
zGf4qN6nQc8dp5Q+83K+/IIkWMCFQ4mnsc7LNmibTgqhZRurfF06/R/+cISQPL9G4j9xEBYEmDS5
Mci3UCE2zZXT1fFQQWIoqOAMzxPu14uA6EQYrC+FRnWO0/xxVZ9txQt56q0cTva6cnlwZ+Y5Tfia
Ii5Kx5eShgRPrAhsAcxAemMDCUSEgvWCPiz038Z1+RZq7Sv23FoXnquLTdy41FwLfP7Q0Ble5k+h
vk9iJZ5E8kEVE0sJWmakj0qa82B9PZW6/1BNd9DST27ciPTCVWstHhARQN05Z1ylN27DBw084lay
DBiVEIoLeq8Ri+V5Y+h6tEPAkCNLyPbzGpelN8McroqMYXwz8sn+/vxjDt54+5K5rlrc74IV7I0Y
EFTH5UvsliPrW3wFRD2wjdvQXJ7aBJ888mAP0XBoW/C0m5dQ5ziztmVpucatn8WW8fxE9RnFuTOu
yLcUo6mwCjO1ShdVhTbUInrvXMm0FCZ5dePc6+5WpT5yTbNMOUrOjv7uZ3NClTJHs1+9KWklhrxy
pZ6e6bsKpXpb9Cc074VyvAvBwr/2eujZN3gWJINDmivNfujzK1wrqzUwtrcvtMOrt+EIZ/BUzgKq
qTa+1nfIoKc5pY4h4Cxcy4jqEDTv94GcECFaoJji39m9BJaLS8l1IUmy0rBCYYEoeGyfZNqrUtgE
BE2OlxdZoFGek48aW6ehZR1cnCl5S1yMAf8pAPUfJzvHmMBu1In5QhAp7IEL44L5G4JGguzy0XWL
LJypatll0suIHYrSxTYfQfvA61n5yXd5TH1oiYQg7cW3MwjG2zcDYIFkSOTfDyYrZHHgL31dPDM7
3VfxbszSGYzPBYdQNNfUw4zPE+YWSEeGYHHktIxsh6Q82lhOvNhOVMbdcO7KOmoeAXuC9VJhckZh
kEYPL660bJc5kJLciUluZxuYZP7gNxX0oi99M2dKRx7d8lRSkJxEKHxLA0PBZYonGZttlmIoEbt5
W/UHUmmZBsw4ub8EnAgPUcXmEku8g3VVLxzrrqRkb98nJU4eccpW/WvIzCJl2c2envf7AUqBAj3v
vGI5bJcdLdMt54yS52UEiJJTQZiC1p+QsW+eGRrAvJZbQxtvVAQ0tg5i+3M2q4kQESpuCrngxiJC
leUdtgSbUZSf5SN6Zzk/PLkY3RPGpTaFpMV5CXh1wszsnykshEcw0hMk5ZxXK+Uq36YGWBwMq7PP
TXkUw2HQkS0/jWV8+0nWqy+Ix6O3Hs2GPOgrvYAJja24TcT43jREp64mcpJqMmS4ysXwyYUPmO7V
pFgclWauhZd6jSacVgCnTLAQtFZ3eqIsH9vu1envDKrGeEgGBpKizri9DMstv10maIWm/uq5o3nL
zy2ulVlZvLCsNpglt31rzXrRvO9ne0eX4OhyOKrmIUl5ZY3geKGtoTI4vEA9GS6RlFHeh9//bIoi
0tjdtdjAu0Y3LlwmsDvR8oGrhlhV3vF4Dj2U1wuRo8lzbiyJ4iY+3gI+7Wzlipm5jf6hfj4gANKW
g1cHwu4cQApmqc9doDndDirjwZCccIpwKi+wYGgQjyr2yQYy9Upj+vU/NFGiOkkzVJlcNeZWFt6u
EUU5hOurO/iOcc+CkzoRx3iKczF44+yqg2CUM4AzJJuxZHBZIDDXOZNo+TF1OIaqvmo7EfhniCRY
O6Yo5fN5vpxi1L+33b2hUlQpJKzIiY1ccjQbMbUWXFGf9Y4EgBGJknOaf+xuyGgJ2UkIim18D/Bp
jJutqV7lFAJfMjpFIzgm6RYY7d3sF4gctpGlXhPy3cRpIm6xrvUeOjMYNSCwW998vDcdEfvH3/4L
bV3FhXQ2wkN8x+GNCfV+mu0AS7TUea26PUkNH3ib7w12S+UuN6PUkfWca4I5jwI76DXLENFESGTL
9eTVTwfXT2v7Pm6/k/gLhXYQfUtfUZJ8JukmWLIG27yJtZM63qaGshOcEMS+qGyBAu0awTsTuWIq
T/0qyR9dg5EnlXtx3aETVthrImKi28clYZig4npOAtLQ3c/RDfeCpGT3laloNoWlKpfORYKoGMY4
oNAnT7kAVzM+h7KlzZ1FFAlnqzoViW5sJvjOymm7irnkmDVEMOaoGBdIrcmxlM9ZH5eKhNaajuzl
BWr47oSrUqxZC/Q/Qm09fGiywbd6s/ImZilG5FQhDPcnPwQxVd7V6xs05LRHFPYuuMsLxLmeIjJD
xweMqmVcD6sqCl+MzHCYzYsdfeEHwGlfSrS6bZ1/OYfYHVRN9QXDuTzket9hTaQ+MEI8cdkwnNfN
+gv/6kdwgcPnA+UCQXGhy7gnS5RU8vkrPOG48+ALRt9bt1LM/ZYqkQDtfeJuWcWJrQvzCj6xPeE1
Ggh2gYpK+SAc3j97Y+tG4jNKwnc/gNItPrzYvAA29lvYvDRSCHpvd4d82nvnqMOPpxXy5bXuE5ce
ynPFNDb21W8j8L+Nf5iH8TRPgZ5TsYOnG9jjEvQ0xnPo3LUJdwliUTkB41xzFHv5uOok+2H+n8pg
BD7sKL2perWPAxRXIcEjGMRo757D088KDv6AYKD7q58QWbsCpri+Np9dXt+5t0e1AjvlHGjv85Qs
fV4V3Tfo1amDodRxU1Rnr5cfdAJOrllsb9bawR4cGtXp86oVBS/JXDTWwh6pLuJldlHfhHJF0v9Z
7+mVWKVSiRUu6hVmG/4SV4QOHt0rtIMDN1dHr3q/M5ADfp8WSmLeXrxZFfwwaGmpDQj3+SNGExAY
fgOH4XVnWi1DUDQYLjYNNkaZsRfJPQx3QfLNFNlBBpQG7u4mj31mm8ZmOV4QJD4jSonS8B8hdQX9
K263zMo53iKzisoF4isKfDASosufkG9jS4XY5BNEh8OJV4VByr5/eVYCfHibvHTArtELIL2N0eIq
i/onpXxoIZfWbPa8CX/VTs4aI0nHSZLZ7mCLzi8e4xvJteF8JbTHXaJDvJ7rSBZ+E1Hn3aH6BbAY
Xit73iv7Tu5eaQiGwwfv9G4570FJPgQp/XYay2vjP7c70B0JflhWdd8B9h1vveMa6SBJ8pB0PXnM
ve3k7Y5wVDyPKLoeEDfrH/UQkO/6PC5gjFkB4RX6dk6+cSriQOLHqzzu5uifu8RBKycJmEkwNywu
rCesq9lpKA25wCl/b11WDftsFSzeMWBGlO0atQjFopw5osZNUGfjcdAXDabjzSGfquZiFblaWU9S
2mzygo87/6HGVddnoKfv7FAvBUS1GQKooTucYtdqek8o17jI0cFRkXN0zpZRoNc5OSOnxPH1G+MX
J3FMinkQfjrQAkv5791gAA/ud7VtU4eg+SJ+1/FkhCOFYg7PghQtT7zTPKE7g4wr9Uh//BFLVYqK
o0ychJlDa8rFM62GOpfv1RWADeNxMhNKWg7PNvkxHB1ur/S+68VXNyak9/ws57aZmB+Fzpdim8z8
XvvoqkDuivz8OOpcIUAZ3UkuNb5vhc4nahZM5OoDR3RM3H0c9RkL9swBtSlRYlAjfiT92nnmLJyX
cSD8YxnDUBa2ougnvRDVLAHlf0j/kUdoz/aKKB3jlHOSFZG5F0/vzRvAMXduNEfy0Ail/oziqaCY
AzrXUhzoDZ7pLs597gQuSzPqXynKeIpZfmhE9HEDr3Xk3vfmM8r3AQvaP4VcZ8Pp1YjANlcZGVx+
p2c5MBJ2dc5nmzWMkOChRexPU7eFYqV60hrIPuVlqbSxCzc+v3l9W9swxiqrubQsYNU49w+bXrc5
zzvag4WF73aEMOZ5muPZXBLKs1qsA9O831Qia2ubufTOrLRdmVhz9q2VvdapvvCWm01OV8+l6sdQ
FfrQdG2Mop4nxeSbk+YFWhtwmNHUSz5dnOIkXzb4wUr7t3nZ+3spy3Qo0RfDwEAM6Xo3EBKwhkgP
CsydKq/obU7YicfDbdX4rXZhfkE7PjO9TgTgkHo4o/An2vlS2zMxs4ES6bKCQvkWWe+CtcwLuHK3
RPD1Noa657nRiRp5TwYnU0Kc3GEajvpLQHmcsacsfZRNZxgRylMXsRfpWGpxPmyG3O2EMNnKy6j/
UK7beFvO7dll0O6dwGhdmNXa2izppDWBrR9KS3CD7DA0Ratdg6vTShqhVhC5230XMBKWm7K33cut
4My5NQWjIuocDoY/fHHFXIDPMQWqwfCjjc9miA0MKepmO9YNYK9NXUCDug5aupephn7zVvgtFYlE
XMLMx4GSR+argwof0Fzb0gZtWLlB5DEAcAlujeL1sq5LveefDQiL9n00Is3E6SPBrZOZr9JNPBET
ffOFWOp9EVCQEs9gv5a/Q3aA6+dS1q0p4L9AsAP5HUq/VHSjT2lq+NsUCQwMwBmcq8YMx02GxShK
jnlDUp+onTurcWCB1u24/iOIXYGtf6SyA0pqMG6Ye7Sye4ViMjAkdKaRP6lB++SUrPlcZqAHa3rH
2dmByhTefX4gFQlVaFNpFPi5j9AhFDAGGtApv8TbZJ5hO0SAh+nEPuZImYUf83sCK1VfGwFevqa4
ZirbKche9v6x8+ct7/J2zMwBEzsYDmoK/y+ApBN8e6Wh/MdEseaI991/RIhXoYbc2QO7fVZuLbqk
Lq20rOu7GPmmmfjYYwEpwVpWzpXGnyNEgTkj0HjnS0NWmVl81/GWC4dvxZtu5swABYuFa/3296Xy
DnboamXKjuY0si7m1kg0eYzEos3ggNC8j7F/MxPdXc2di9vYKxwJai4wi1Exuw+rLC6sCoUaKkaV
y7EeuYG3lohPW8pkX+JUVWKRiqELujg9QM0ududipkNhKkJTHENM3sK7llrzgpyZNlu8g/+Cpci6
fx+q6lLdTLLW6RgMCDg86Mv9L2LwZiCY8SZIFpPg7YXw9m255A7l2UNH1Sh21RzuQAhMqUsS6k7O
AdgY4tUW8t/sV4E+vRxTcEScm3p4Qfm8wehd2rYHCzs24HmJoTdHzWyVHBG9/9j8UcgZJGvWMBMg
XSzdb3tuR1xpbec29BCUG1SJLDfIYi0G6bvT7rMpP8Dn/3ZShyva1OO0d3Lhi1Heb/y0Pw4tHfLq
en1gp+bU57egm1NF1u5V1TfDMjghbCrNpIn/FlJHAcxqlKJ+Uukz+9q793rVqp8uyc2tIS94bAyC
GnbBLE/dzAPeO9GDg22tnTfhQFX3/HplCXewLnO/opxFPxU5oDHpgCz+tU5YjlFdPPyWz8zHH445
oA9v03siDQxWAA3m4agf+WmpBzbtCG3JdDcmGDxePhE+SQc2ODdHnH5J0HTBnyxG6jWmCCljlBPY
HWeKn33FyCXMxxoePqVp/iZjYH8LNDiOWCrDtrCBa+vFs5X7Kch2Ou8WTpZY/feFY9eTdIBZe05O
KG64vCj6MNY1buRfXK7kypcaOzT4AIZKp5XEXA36mOL5H31O1JE5DTRxxO8/EUobTFmjKvmRu+4u
jMrk5F4i9o0tE2zxh7Pleh8eWH6Qwk8A+/mwQ/Id7musPvMMK43GXXLJTAJHThrIGuip2S6Yrs0z
c5m3HHEwYNLmV93VSQ+fRiY/3PLIpokfFLJr+iuYwH98ff4GqHxNyjxI9+5NHtLu3eDSSEe4q4Dd
48El0qZ0ho/k2vf0NxdbkcU7sfhHE2u6kvoyl2a+3d2aydr9qMQRWkp7/Dy9nbJUSQBHHN3nYV3v
3FcD9sWxjdhtdr3Q+R5SmSqMFICPIF51BdMTic65gkfLPOZBzqy3A8lyGjA5ssNWMP21subR6eI7
vlIZU5TTeuTqe20gR8WLEIvswbQwZkw2rsD4jOrT1/ddShHW3nuiMg51AGnKEO2chEmAuzTgEHOX
IXhed72mTerXe+cZwn3T236AOh29w3RhfLt20JATKcIZBM4iKxLOSlHzrfIxBkeqreGxnDnGKQAt
RlhIzKYy3tAaK0UPAwiApwt692HmHWSj6L4I/M4gpxIFdAsDfFk92ux6WKXBFaNqTB0DNP1M4s1e
6c9u1lMaSAlSaV4ZrG+AfGr9YvPvxEcwkpneki49a3bj3mGycpHiuxS0yFTELd1nhiwg9YIhVrop
Yyu5wvQXGsEth8GWk9WJXa9yeqyX/5ODs1agL8qM9aMpakvacsRbFp1kNpGPgaGxXBDevw/vFOHu
1UMg8ZOIjLA8zLLI2I3PbgLHjc9S2S+X7/lUKOmBwkl9vsM5dGTwFRL/nU/QQStwAf+Tfgoalbn6
X+yW22r/17Yl+n0NTEYUqEA1D4CVkO2Os13H0/jkGyd1ptSLsofxFgfsmaBKMkO3Cb3lP9E40dmX
SxTE2dnPIvhvzwYC66olEfXPsy6YpjGKrSknZo2xDQS7fK/e1pxM+hxBy9VfQI2Scbc9AlVIuWxH
PS/Pju8Qp2wuzLfjuAHU5oyB6eIaY1IGTPonPQg9R6csSxs+K257lGNFbRdD7etyO9tRmGhXTZDa
ofkd7h5bTdhUa9uGMWOtjEZeH8tziCdz5KbiLC8/xFCKxXn2texnVpiuxt7dydp7D+fHoJ92Jt5g
CJ8gmVs6+r5y58N7bwhVnF+FSdz6vSyQn1uMzhfprL7ZeztU1Ohs4Cs/z1Yn6pbhqXrIhwKlBwaF
ulWOwTVeP6at6j8PGTA1g6WX14bL8vh9qGvLrSZfgHS6fdFIXKImzkMbnMnwsDLVKPVIeZDtSg6r
lDKsQTEe60UTdd2Coh5XT9otPFuxwQkz3TZ9KF29ILhziWOLrDIuU91nZN/acLIXrI3krXYUzL/y
pBj0vvrBIAFzdu0R7Zp+pHvQsOMlr93aEMJX9uipuRObgSXqMMGzOwf83v+iPTW/pqG72kN4M0Zw
ppNpwMslv6bxqOg4EaulKF83Ab0/8U3eZaAvJnhEZ5+G19V5CI51pxO77BLlARQdQpMN6pR+9IjI
j40WuIQJ8Ef04oId9WM2aesSbsZ9P+PeW6WsS0WG/dL7lD9R+iOXUdx+koVauu+ZOxVF0+bZo5bU
lTIkCB51zqOyToSRfgAfS06niQ4A+QXbArNmDpU2yVvlqKdEZ5NrRQTHKypeBCrLkPD4NvvfhJg/
QDkNe/MNHrFRm+0aGkm/BjZthjguKAVjwsJCUVmgk0ZQWdBibZUvjg4uub5oDfwpXv1pQ9ctUyfY
kKs4iqjwcIQrUKo0k7vu0kn9ei8Ify2j6A0kTK1HHSCwEsDgkSaQg8ZesZjP3cy6xByMDmmSZThb
/m7n0uw6E5JZYraerUOe9L+WdvmIgCJ9Qq1bFL4iJrkmPFM5jevHk7C4p9lydg70sGStq985map9
0fW2zHDcDc3xgJ0rFO66eHMf0sAl4pO/deF1xnL3q5eNiIu1XOG2VbnwfpSE9x14009Mpcf5OlGj
iggRzPqpkHb0A4xmrxGhMPoDuOASUicHS1a2XI288i0OfBvLhV+0zcgGY6AAPkunOu95CIvSL+Ub
0v0RXIsUN6dT7e5sRdHZBB5WKCKQU9djk537+QCG5BF0ZQLFRV3ZWqJL67OnSJ7i9u4s9U7rM99x
8vCx4i1pZxY3+NmfgRDt8/s/Y3lo0oIacDgmyOtdVafoFngkhVnyoQUPifDdCbUOOM2ex9K22SSh
+TNJXMkF600HwfqdU3XeWqJhdu7PT0avEsS4E1pMoy9Jq/VyGA25E4JB3WbyGR91r8tzqnJHWAy7
oArLMjnilY8eOVxK8/QMlxprCoizk9vO5xGOFcBU2fok4YJoplPZakrkIPpnRoMHI5P56GddnFal
kpAX9W58WlXqgonB09+H7neg88xJX8weeMMzUYzKH+a9jwzmOByRZ8g15lJ9ULdiJxj2iYxiM8iA
7hie0mYZrc1FPGkKYa/SD8jvpD9lCNj9rysLfOz7KO3/TwWbKYe18G2rPHFzkaMtjLM96Qg8N5cU
CnIoWg0caGw3xuZxE7GY08rocdq0vKjBopUdtBKqeSeaN7odBzB9LkAkL0lviNKVPZEDvBQtGxJ0
3r0LKQKJdeS3T6iFdynMh24bZrDtqQ602IFH+OSdIU0mH3NyrqRQXlN6Gp6qRR4kB++NgtpDEIVY
KCoZAxTbi0+cdFrsCLYiVnaxNZQE2TY3NFT78sHMQPeEYedpIUojuMtOpTbRUJwDbeMkEayGWvHb
fsyUY9Qwcpzpnv95YjN2wOA5m2dc3RZu8huWnvtHlcSUvJspfAPP2h06FaDPLyxnP7zo7R9N3L+W
fQVj8k1ryuhgZvbX4w0KTceR1jb308NaQfqVVsde/BS63V3lHCUJ2DEUKcBUDQN0+441/SFsTFbH
5XyfIfnm0qxjc9kkXLkqxoOeatL9SEDpArHMM6xVU23dyv5RT8eNF+rdrkHD0cs0pWTVUH0Rzio2
3w8JUXr0kGlOyMIlaGtPeb/3TL19R6xZCjbgoyrMO0ZsN2SBYZEjZow10+X3HEnILmWTZsEWS3oB
vDSz2/daDNiq9KJri4F0RQriuScA0Ft6jgcvZ6PaQCyGS2xEXsrvLoiwbDJg3w/xGtQqTPBOopLG
pvkWrvVzEj2Xc6/xenWbT9z+K31dCXq3OgfZ0n9LdA3mNoqUCT//xnwPKQA3aD9ig4eW8akicJxT
J5GPvWj3AjWAnoko7DqeX2PIXymwPNJ9xArM/SFE2fUvdc+C8AxDbcjcF6HiPao6mqrlHtCfqLqz
9e4xJgnWVX684Ac2zZROg5GhHrxVTmmNPNulHw2lh9sJ8vMHw0z9UBAQDxNWIakXpN9r2m937WFl
W8Z/b9C//y5LC6ZbMZx4ekmM76dM5HtdCtWj1ea1tKkkW8ib0UxU07RjLKU4J/aA5fqHMJXyhmfW
4vmz/FEScfGznbO+kwQblTKvA0c053w9yEGW9ce00NZs6shwLv4QRxJZCB2vQRkhRwhi8E2oCXC0
e4madV2onEWU7npv4g6oa6YoiiqA9Mil/BleSt6UPbpH5LwRHsTGpi3Txfgo3Qt6xDKeWyYoWaNm
soxOQAMW/hLM7kJG447wf0tShrgPVPtUYADBt+bZ8U9R5xPC7opZnE+5yCVop7YYFwMLoZruonhe
l7lvjTEC0UScC2nG9Diju3YguUboMrQQR6wsUt/WlNjklBgl0jHifT7V2af+gQJbBKwCDL4Oi4sl
8z3KZkekIDF0cc24u/iMTzN6qXXGtqx6PUVmCSHk6qgrxS9wPKRBussAy5C4EsiiiuHkdzySYoV/
LrRiEmAGEnhX956uR7U+CJt+U/+50q+r2bzDFE70ARmg8sHUnHOUc1sGzGUUs2e53+d+DprSDFFD
S7ll0yEt0dBTzNrPHyJ3nwimmA75Zns5ZMqDiMmyU8HiwohiEcBLTJ0JKqyK36pLfKdsQRtk9yQ8
5hOmKoOrya4YaUoaUde/rJSDfsT3h67g9CNWvra/VWw+VjRxFMOYRe/zcf7UPJb7Ftlrjsrt1d8+
uaeXKcWCdsbtcQQ0+vl0d6K4GKEBMzaGOpidwjzEd/syACIeF2d8K5P5jUBYrScenq286qmotzFJ
ks1BLndONKkcl2mPrxAUAUws6YGZkX3FmD32dOcy+BuULLPndO6Hmkv/34VFy96V92v/iv4Xwg9r
vpIo3EnRfP8yyaIML7KWf1Zt0FLhOrwV4wheck27Q4Lg2OFm/dua0TlNQQnbM/euXMY2j11suwft
KCOqcdzWDIzvff7AbmmyT6/VU3UM3x160rHml33WsdnSHQUH2z0bvxiWxZBcGJNt7SCDNTfP+Awe
yxUiHtdXsUJyCizkEaLJSoARxt09vX1CSNR1sveYc3yOWqK9FgnThEu5qf8BUr6fpPyw3ffkg9gD
eoxzmHuzhqFy6NcfknHp8Qp0IejHj2AIDxrxQZXj5GH4AEc0cRolLdN7U93c4BXHrgPoU84irAX0
nNNRnfX3ygvOLVUzkN0bzyeQqchANnrTdn74BqiMn1gHV2nQZ1s7DvI8dSFz3bl1GrL0+acvHfdm
mbBIlS5hf0Z+0rcRjt/+XnyZ6s6vz5Kbu/n6TDOfxC9CfquLcnwhSta+x3NXIMFGshFUutL50kfX
fyGQuTve0v7OI3A3lP00oURD4yUG8hseT+bTI7sdE0cVX8GjV91y2SQ/jNWWQ8hsMD6+URn6N2VU
LbdtT2vzpyDIdICGVIofNQV0iF6UMtIIYGmCTTpfjr5mdS7Z7d2mdmesI0m6glmVxBNfCGg+3wn+
4W2zEQPX7C2EFWLhJo7bXfAHRo+UVWdSc5fIEMVh3BSnD2gTi4iitlvOU53OLuDGwiLRkDxruDRA
JeJuRSlFwtuIh3qWmycw3/boD++MctRLOSVwt3VXhE+BqOjRqKVt6oe2SI/lSG4+DfXi7iYc4DsZ
OPsfEGfDq+N8VXJT4MILb7XAg9eahoCKywv2vyj/wlUC4KizGqZKYSX0DAygLxM6EhIE4xthKdo6
wlFW3qLpgjRTQIJc6F9Ahi1dxQBim45MxZSOnRUOjZUMds6Uj92iJOIOzyg95Gd95dJ32CONG+l/
YY9x0M9NE9fsctDSMR3xmNWlM57b9G24cqDjuI2GEhh4YGNlIttOTi+cKHmQXE1y1/z1BOtzyEt6
OBcBMzKJ7rAG3bfwwEpLCUNRqxYGmkbEEqdyvvg6hsG+Pmmi6YtGxt5YyijYclXz9XczRJTbigqN
Mr4XmoBFxr/WKDg75KxcXD3L5OucwR758FclqIWMfQYTszgtM/DckUr4+XDHiPfK616JINruxWw3
l1HsfCbnVxsRA+s14BxUN3ILPnQdd8BpYyxRsQzWu6XTJeD4ROxkbP+/eeyx3uXkjW5sTxHbTG3Y
2ySxukvPdg1OXwlakTR6mwz+5iJd+hQaEVV/X4LR+arwIVHJLLaPqFmSOM+8J8ZbAQSSiu8J6scd
HjKRyBU8ZyIE9KmO3yALiUrxdOUiXtHP82hJN+wOZLJ0OBWIh2YDphgi1SglKvIKB+qociFDpaCM
9o2IPzBg3uZE6Sluu0Qhrj6SYA7DVPeDGy2l/2UoOwW1VuqOz2eK/mC/tu5Xc16l5WQpgIWD+l5+
CjD3P/qbiVuWb/6jbHoa5ukLUuHvLUYAL1qjX2BY9/JuffXjIrEQw9cMoihgA3WU88owBcNjNcrv
aNQAIy1Q/kmZxiCJ8bkGqvcLPcouerSh94DEkEHvuWFhDvMoieWlFcn9OWRG9+f99Le1I8ZtBWvx
TXHXcaSr+g5VLucxrpcrpHOHUincmIDILHEtWTlzjm6XABgoI0TIIqmwE+5ajwPc7arY7wUjfOUp
tgypInSvsU3EMbxdsOURcIWGFsEl28KmWgybmho8r0kXq6mugDjfv59BSlonsRTGcWollRl0leFm
shCn4Nn94VUFnk0ulyg22KtfPbsjks5ynQSJwtfvI1fLasYWxycj4nw5KShcoc3euNLo/bkDeUtr
E+krG/QDhthM8g0Tjhvheo1RYmNhl0ljUoCeU3xCSd3QqIGHWhygvGbzTbJicZKV1IaiiuBg7vx/
Wmg4Po9x2RtqRIx6LhtB2u23Ve3Mb65GPvbZfPr2yIqz0kIIaZDWA5/d/LPQMITQt7piJInAyLUs
HhwfExoFhuDLvah7RWiWjwtXr/eVma2N52WQHIyA+mXt0GADA1o/AZ0xpKZ833DsKE1CZz53Yk7d
K/3BLujKoFZKQeYeM075+yPxi7hAmFT5A6j3jGB6Gby7nAFvnBj7ysF3t56NPfI7cLDptU6hJikK
wlF8FfGc8nM+73eRZHAyXNGyn7G5Y+IYitBoUEe5CZ3e8MTfu/4U9NpEWtoCQk9U9Ks4cM/fhM7D
ivomUJripm/ytF9oBl2Rg/thFsZFQN4/Um08Dxwnk+x6OaKxPRRX88O0GQ+wQ2+CGpPDFBtdS3Vk
5MMiswUfBio+aQjX/gfDIK6qmVE91OtotklyzbiPzVcjmxVqA5WDMNRneM8RnIoyAQFX9k6xU9kD
6m/AFBLWbDX4nrQhwrWLclIS9uKUyz+3yR0KbPF0dmfMJlV2XQuds+xZoPoVIsP+/vF/+hfWe+OR
lUZ7iWFrp1o+7fNORmPc1SWch9wPkpHGpg/cOyQidx+Oxz2L1Qj+sWWpNuQ2E1g3mKiY2afDu4Ai
2V6VNJST8N9yF4VGFoELocp5+R0SUeXKuv32cujc6irAIFtvHlVwveuwWz5+Xd2utQQwwmbPbWvp
Ko5ZNeqjJsmhB36nawOrYHQALfRqMyLMrTemLHOCXKiwITs1pv5GtE/W3tAnoQ0RfWjWgZNGmNpx
wR3d0pM87YPEm3R78BENXP6DTydFKTcKAhbB11DF+aNZnD8C8ndI3UNxLAqN3GM38RrLp6Cs1s9o
7RM5PlG7IrL7VbkwNbUUrIUl2z8+UgNdYPNSJv+nuzpcLpZWRJW3JVw5nBl7sBbqM+lTQK9h65cd
5wgeqVhObrPMpBRoo/4PR3105pVDD5kEBYywwazeQww/DN61k8PbYTh3sK2x2OOOmbJfVHbyaOG7
t/Vf6zrShhn8/UCsTdEKRugxqNCmCzZGeB1F7++AC4Bn0yGiywIbXhIzKdKpDtONe5YQxIzYRMCx
8Y1aShcNzKy0AhiE/lPYQ18BvNCsWC6OX1I64Bo/Mp/QLxrLukRmKYwws+VI7K33UYEGdu/prLtx
BehnvNSSa+WKzykpnLxrNfZdKkr6v/xpHqc/zhoFpG4/x3CI9zUTapb886Kz404GKvN5WWMBh43I
XJdPsmgJ+t+VVGy+0rsd1e8mTxda3Q0UZxnu5i2RKPMgLqIrfHjlsgb0evtA6ooSegX8gf1h27Ge
KjSlB2Mo1EElaBoRpz7bM/5alllDCwSq9hmyqLmRWAgv+Kl9bey0yAsIsb3JBcX6xGu+VShVHLNl
Ho6vkYgixnrypcRimoh/8+qu6khnseNTUImlsrhd/q0yCt49EXrFNWqJL+qYtcPUhSHOKWHmCTwx
/DIsjMOjBJfyep7t4/raPZeGtwqxGs4o1ysnpPF1pS+C57DNRHM/6LHKNIH9yh4l9yYWTnNxQFpf
dn23mteCRmak+rorKQmFm4BRck8E6BFoncnmnHAT1suNHLWbmkaCX63BucKf9gyT1dMKVfS/2Z8X
M37evH3kBGjAU3R67w8aBc3U44GXgBdnG5kPBY3gPiMj12ufmEEutmtrfgjNX8KMoVrXNOuk8Sr4
W+4wyrfEQxXHjPM5y6NnsWUIOj/FEWr7km198QZ0nCFdDzHANMoLGtdf67SnvaToGvD+I1xDxkxE
kIUyFQewuM5p3fKfChhPfiG53mnkLZs6CVIFlOsTFrPeAzQ9xe/g/tBmD4XqQP+7V1gd0y7nSWhC
/ELfCqhfXbp6cM9QhOCRY68DSIgjayCejodDrE+Xh7fBTqruTkxUmLW//7r11I9apFNLz72mr4z4
QA3fhCy9F8CdLJT8MYazg+HuYNiX0yPQelovbSnGhH09c/9VBD/zFou7R5LD+Xh+ZXuPVgmtEen0
pWIWDce6CL15ofm8tuMxcJGgDiSBsRiDcOegy/Pbaji2iT3WpWb8trnnBgxg/Hj1ric1E57nYY9Q
8hZO+KVToSW4wnCoecE+PWChhDnQSPPcLg1boVvf6n6NBvxQmhwGY9T8ei2BKHNtz2Br9fjtghKU
8leG1AVvv8I/m/LzIU0o4OUUDJOXEYeYmVdKx1qOltCZl0dssz+8q74V/gO4EfL/IeKt4P00/zHC
5TJwGFgvvbbC2owp6lmv7GWZRaufaJnzkPDYdaNlKk8sTJyCXp5K93D7Au0byu05TT2uNXUiQfJq
LkPb0riyYKai/ziQskBE2lXoymlytQoSL83ymk1qsf11pDl9C94tjOyc/wBOlBDGQKkwbzQtkJh1
4K4R3sRYEFNRSNbQzinfakp9KzG/qBQcYU0sifjNbm9gb3gH5oPuVBPI1NQKWPofmRPDvFqP87M8
cg7WyBps+U0wNCTcCQ7tpDqg+Gcllam7NDCCmWNkUGz3Vac6G3hvEHFX4JCsShc9yAvx90Y9dJa1
V5oAUXxRTbWb1E4/pUp5yvMkLxMhzjwaReEF+VKK7Zxamy0dHwkX1xaiAylJnir1f7VEjB0TWREA
ysq7me7ibJGTb3+aiLnaZtuaUqFDg1z4on7BxPEwncgbNpxrQSpyizUAIvT+S8BzvwNDfYjVOBKR
doTLFRS6+DzMsKSar7eoRKm3FHKYAKjviX2LEsr8JuavRMZOsXVDWDEYrmSneTbJm/PWMM0JtMD4
GLfGVJIPT0uVsOMUmGbIH+2Z9YC1///uN0DjO+CaNL+O3SlQ2Y+ne0VPxxd1qy8Nc+piwUWh7f41
tb7wPYrsDz9teRjiGqPHaYEgerrLg9Uk2mCrXdTkxCKbgGVo5ojTP8QyWPlLSIocJppwx0FzhFLK
1KxhL1FzigsHDPw3YMuI+OYQE1cwFJJbLW+mQqeiHtlh+52RrDEbc+EEc4KR/EfwhKYeWzmhIx9A
4W1cC+9p68NLdWHEG1L0SgWrHyq3JetigOyLxwhhSmwi9w794VMCyX8l8EIuZxScH6ay1dKQoYSN
e+o3oKsnw8/Nu4PMTiqYkkrQ8puLgpSb7Dd33PJpfd3L9aJThoAFICZlitknxBjUJnJxyohOJ71R
P2vKG4YgTTT7QfgB3WkfTmaSs4umRUKdEwiBF8hVSBs4Z7owEXVZxuBRDe3T/3P8crB0ReCtoLMD
HjpuD0h7ZwH6jIPaEl3RnVjk3Cpr7RDe6GAS3DNKKtGWOWMTxBGPGE7/xrnTK2NxlW3A4hEUyo20
KUx50+qZ6koauRqpuUWb9sECQVHnsz9zy2Gc4+V1iTtYaCHiC6bkqPVE0rrpVvqHOoDN108CAGmD
HQoPnD4x0achEQKON1B0YToS1yYQsh5VssobAj1LJm79mYomFh1lJNdRy3HLyNIyNR1IYE0aKGFp
J9BVM+aDCywWFp+ZHjchLOo8iZfWguOxfxTRhjU9Hrk+W4RCd1QMgMU2Y8WEiwBET2fM503k0kqR
h94rIqwndPKlBh2whgIVicuntRbFI5iUVSEhlfDmjmzZWEE/BaW8NI1h2JAAuw0o188xFY3osRsg
ogiO7SDL/PHhCiINLrC0buiycjyZ8DCvS97Fd/vhLMLDGFTajcmS4QKKwhLrO5WQbNS/bEj9PWBo
Ud33h2EY45E2T6Z9BPu2wC7+fB0aoSyQycw7KCTHU//pYo+/61gGlBLiXlgnxXNE15ef080ubNqW
VY6pGS+Q8n5T9fs0xRsTTBx1nmDerWvv4InOQLbvpAmGyWRme9zdC0wkkenyPIzkkyq67A7XHfNK
sJ9OeI495A/ZyZ5hoWqBunWrwnG/CvWUCxyFH8SkXTQsfoPrU6GHa/FlYkR60+jOZjUy6ZxPXLCF
8DZbqblfYsLEQXPsW5IsBDAMfOWpjk6Yn/tCvxVzOhH6gC9kbrQsUD4W0TgO5yGAPmpmwkOUq9tf
DrHZ9i/V1guOIkJp1zs3CC6r4ouTmSn9o+L754cKBfAs3sBVT7l6L9DrJMFGoDHUfa6zvt2M6yFZ
pya0QOapvfBiqLTLvw25wjx6cCR0zbMd5nA4I1bhoq/cq9yCfkZjh8MH/xnXoKVSbZBd89Saa2HT
erbiLbA7AbvmvRaCKRzgr+qZE1Dv3t654SZQZoDmV4/x5GsmlWqNT1g9DJFeBEYq+b1vEh/kstRo
JgA+ntSpgbkgnrn/CbNFsaAggJpTLyIrD+joyw/FgHlj2ScGBSehRbdWa2RBPecvuwhCc5VCCmYi
dStlctmv+xXelzY+jxWAdfgo8xOblLdxgIR1nzNfQG9ky8eS1jrmnBV+9AYfjuAVilVyjr2yE1ce
W6RhFw8edoupSfuTbyxeQZmE8fuibuLkkEOm+YvGLfwH+gHMAHdS63MNjITo6LqqOwy1Xvgpy85q
WaL086tuV7AmPlnaXvlG1pYHY9GH/rSlRxOYGMZoAe7QYq5WbHppWVlH7ULxpLqFOzejuEATZ9AI
a2jjT5X/2+lMwX7mMPo+792Zwd5IsgV4562p3+f1THpaq1epa/QSw2rYtsNNz8t5wTfMPxrzn2RT
HuAfHQI6wAECoI6fGz8vFURy+P7j44EucMPLeO1GTB1/biUnfusVh4UUVxshK2KzhOVAKSjYQubd
a4cntvKTLc3PfAnsNZqCjGnPMyIrOp0R648gzQpAIg+Iy0ghuaRyLI5U+rjzrI0KDZgwn6PsSkj5
+qUj4GjSCDxm0GXepHgOxk0wc1xHkvElwnU6VUdkl1w9GN34XAh910+oDjCgFVjqg22jN0IjDuQM
AOo/2pO255xeFdKwLgjCm55XDcQvwevCEv/1PdHnz5PEK39qf3xIBEyuK6+wtDBU9Gs+cPSogkEp
00lrX82BUZ1Fx9eoCAimKGPC+Nuin8vzYyotMYip9fEiZsO2sMp13zNUVnvdRlMzlZhhvz+MX6CV
HiXV9St09GZnywDk1jJqtg9ojbM6gKcKu0KTA1FKKQsOsRkASVkRHaLYIu3uOfzfNfkiH4NrzTdb
Mh+yuLyxPP2yO0GjLAooeS9LCqWx6ox9JkLsZMpn2skZTSVTpuLP446hPN/OclIBKtRFFcNc8UXu
7E63iIgURd+pFlIqfQNn0lEeHhiVX6u0/0tWoO0vtGtSiR2rhDMPIb4Jv31Ojpc249E8j74ZPiNx
RFrtnxo2E313BlBuAa0pbbf5JV01+18YhjMgefxm2gAkCGhywsg+MfdVEYrk7i9LiCpogDRwOEp6
Ix2KzKvIpUQf579DPjHWPEY18wKvqMwMi8kdh39NrDV0zNldAxHDVdNAYoV5HShhE8k6OzqaiqcD
YHPWgLMl0IR6WY2ukOiRBqArfU7DhgkXHKbzB3pMJlyeB82IEJEXc3cLCiFEP6eGFOuRIU2GSDxQ
DGY0AjGw1O6r1BojQ7v9PWVbHF2xmVQi8N/uBT+X8FQFJcEsVpIxvzII8OureYpnDEUYufkYnES9
0Qw4crwjdgf9bWDVsto2odpYjmRKqcMG24LinGcTRVM10Pba1pqvNZpsF7clTXcSeAkE1qDmzxAT
3V48yMiqQ83CRpcTgiNeGI9T2z8pon42E2zK6Fdya2p5i/AtCls+CUYWPgfXV13iJcwC0P8/8A4Q
PVA1ij9OHsw091OLBG67KWauRa7FXImttPIMvJSJpAFN9vCtQtTxlquVBDyqa96gmX8+KgJgA+8A
+aMUxBkh8tF+ixsJC0MIPxKUwQ24MoDAred3fqAFy7MsV7tsd9lOBjm4vZrpU2urXE79x3CjD2ux
6wkgx+y34qydCXelUIiNRfPiBGH5LOn2YHR9psLaonU9DwMbVRasUXlBzjn30iZxbwnTuvqAiOWo
D8Ua1S7GT3rCtDgJKtlF+8YNSuH/IiArI+RT8mY9FYK4j7KqdMM2BiNM5RXhrfXW/k+MjtDdcHX+
73RnBTCVluboXvKmk3CuLssQeVf9aL+knnT8WVuxqVbSPHfVS04uPy4OXxyOXw37rPgDiuqTFw+e
g9a+B91VyW6ewv5B83x9DXqyklwGmDW61bBtnK+VneRT5RuHB1p0tBUXxxvuEIsVbDnT5QOE0ge3
6WBJlIGdN1YHwaslf3C0Cxd7uHl0c5TplG7JXJ9yMKTfKwVB9CUjo86hxZj0jRALjng/zpysy+pJ
NubqW3CDa6Ss5kCyfcBc3nlE68oa2uGQihuF0v5sWvHzAFrx0pZeN5qgFEWbyFZnsyyznNJ73zrR
EiYwxg0sHrFbMQSz+9K6TOZnoI9n+z7gsuuvud90VHi2JwibpqCfNMDJIOZ1HleW25E2nGICvEn9
uQUJ4gykQrwuZ01z7Cj63aPnFaz3g38a61DLGOQwvYXOoowOVdvz5DcsvJzksw4GJQK9B5nK5avo
kKfrpT3/0pTWPPRWKCXCkDhQnB9zwz3jiS995w+xwm+YDPm69AYZuEP3B+pX8aTKRgZIchJf0wuD
dLk+Sy1NgLW9jjdZINLow5fslRPE5aSk2sAzZzRF7fwlDzYyAHpR53UC8Vm+Oe8E+4tX7GolsGYT
tdyQaTV2U4rRUeFOndzUjDaHCf3uQn0vPx76AkiYWghi140ryMqrgsjrOr6eRh0Ln7MSoCjMm4ZL
NhZdYKYLzJcUqH43gontZvfiA5SNcsstrGX4B49spsKwuXiqc8LJo+3rOkymtpGa5cMQ0oCngfy/
TRlVC5L/8xcPXpdo9PcdAJUT7NjjIfl5pSz6GbFfigl6fjpTEJph0PhSDmOtjo46egHyhp282f/3
8h6+oW33FjmZAbzn4yD+9HIKiXugIqs6DclV/FzhQGj+kxuBUqU1tDOS1/u/8ZXAyay1+GCMpQDI
QfIGm94wUa2WbKJL/rR6vllrmnSWG9a8Azy1A2KzF/OZL1Gl0VXqxMXcldhTei8xAZXY1OLE0IP6
VQQHjqo00IMfC5BYo3kWjOc9MdOJ98xU0IFGODWANQFZt2J1rJeMMA9DPhIcHFkz+WCkUaipI/tV
38Nm1omiCi9mRCLtZI8tgQs3lCLtzn4BWJpoUh4Oiax3K+VuJtnGX8iF0RTm9dtJKvzO/YEoHuSv
yPKPS2upFT133U06AwlC//ux+ZzJiGCddsgW39X7sqfz3mGzK4Kown2qPpU67qyToGVh949t1VCX
wA5oCkn7016nyhCkxAIE9RddMAnj480Wqt/tJcmtF3G88f6CDx0Jmsnq2euIFBbxXFRod63r62Pe
Qgb01FJovffED9nLhvVJmj1o/ejm6upW8kMqSr7GMzm4rXg21KvXGkiviFdUKZBLmRPxVwq3EN0c
aH5ofAbV+99yMTe05qlE/DLR1QOOcUEIUAlQKUrlCr1WsN11BafsSj4NfYT4aMbPl6VZjryRnpQl
rVQOv5YZojC9R33BUC725Fn4GsrfxMWfggdypu12h4peB9H3THVoZrpqh9bxd6Kyd2Zm5UmjuSCg
4JfAm2MBcW/3paigWq0xl9UVTTv6q2uQGPKtfT3fhy+70F6xafPzWrZLU2ky2Ex5Uvq/p2ZpCz5T
A/bSfwUBoOewDbqmUEu1VmtH2LQ0Jpz3W55rsSCMFnYQ43k/GSKx/TMxkiToaaYATwLD4YNfji/T
efthWiX54yQmeOmdWUKBNd32bqGV56xnJyMXt5yG7SkGAmhYLYTKS1CfZE0QBCS+sFpBaRAaLBVp
nxXXeGSCB5zEb6cmqh0lOHM1+RMVjt48rr++JdBt3sFvPP4ehK2S7tovmyU9iSgAOe1TC05x94zH
/spg12TToB8nHUi5gHI6/fFgP3gXfugiC6Bxtsrx/lemxUA8l8hHzX69Y+mf5qJJUQ5N1j9I2Yik
2uyLEzDFrE5Rg3X0MH89G4ma+6BP3fJAHqVnIQh1DxVjrhLZqZ/LlG4ftW/LXvV0d0YV5yqpTl8i
bIVCW9A+8FDKu5sbac63tla9Qn39s1gWNdmz3zOiSjcOB/kzPoYfSKFEiMklzoy1zyPMJhh0wJbi
aGn08bmgGtG+ti3LmK1cWE1HBQKc9nd30BqBPgWS/4IFUYq54Qi9RprbT3peoaureWvIAdXbmAcJ
br/CsNSNlbydwnV1u+/tH6O89E1Kql62QBNVArU9mDFN1Fgpfx2HHjnVpoGzB+YqMjoOdp5761Gy
vo4mQOUK/ovbWyQG7+gu17ozrAbf3zYsGpSXXn0Qx5qky5KjuoO491lBWyV9UOzMUgPqcJE5ooM6
VKBGUH8fTbfxS5qhMo9+sm33MF3HkXWJblk0PNgSpSHw278rI0o9Qb8zjnC57Oag4os7Lab7k/gW
byclplMrweWoXMBPNFN7FcfpEoUbhMUvHFcxo5q/8GJ4jf6iu8DvlI+yQl+T20PvHKMShIV20Ahi
/uCdkOPG+VJ/dsqLP+efE9ThWKEc5xE+GjyUbD1GY13GEk+61dU8Gv+rRqVp6nRS70s8/mc4oloh
FH1v5V8kw39xCWsHrsGu9OJ0UeO2GHvHE3z4FRJIbyAcdp8Dl09YVTMS79I6jMSaPSPZudIi3ad0
uiAOqW3f6mlkyUv6k0GjyLqSlPHU+k273yZmHwHXSfEHavOnkLibJaItERbLONJsLqa0NMqcq/p9
cGFrN1zZYDUhXJGhoMt7ibwVRE3udW22EN71xVOtgUdJPBlNJ4nI4QN9vP487oqQqLVPmduWoKNl
aUBk6MpVcl4k1it+P9uf20rw9UVefl30Qq9xhG/h86rj/YJtOM5gos1Pnh1WDwlUFy8dfIeLw1ra
ay3IjTmom/rhc6h6uujcY7VYZLMzJa+r0O4GrD4Rc3pPdbAirnNzKlWwfPbb22yGu2AW42cghkUM
BOOBwuzz+tfcc+qtUhFQldar8JcdW7TcXJCy0ygaI2nv1KnubwUUeRtQTHGUiYfJlXOf+QCliNi3
jRFPjMsBCfE0nnf3hO+KHq42HLEqoqMcA/v3vc7a7DxgJ2tInu56sZRT1tH1xoA6w3LIeyM9cP9v
xzR1kL8DQCbV/6A7AMfXdSQvOKXogdF56pPTJRsGnL7eR+zsRnq+zhgetcB67SF4wrIro8upn0UW
QyurbOJp33HGoYqwkmaLmf4g6opFjpLJjYelXvAg3td/37aBytN8FZXRjGDXqYh/9uV9Fk3miCyn
qOas8m+gq//LGX21FqZT6WYBgdAC/jHFRnSyYSSVPMbz5id6kQlk9AQAmcSRjgzpDz8pavFnX501
Pa5OOq1olFMHZIBiNemGjLuR/csas6EPyWYp0hs66MdSWARxHe7MBRqSWBDlf6w0F8PpFMDA+/Pr
93oRFkHakf6uIkR/uRvJe4U58TQP1YXLxNwQyCk+RZ+hx81L14X+/qTVoILDA7rezGNrx/UW4ens
f/9UiHDcAlC5hHNi0S7hAe7HsX7+bZusYjzE9CuCvK2bbc8Avb8uEwAYnv4RzdxEMbsSkAK3P58U
15O1Lwr7nlj+A5Tm+HLtA1uspHck8IEMHsqYbQs/wLeoNBLtftRrz4jmDMI+BDIv5/v3TvpBcfS0
kQVeodRD0yNcV5AHipE0tlcmSxBlQSd4xbve6giV9OKOgD9wZbFeAAwfXgs66qjORuX+Tu8SfyKF
QdOUsYTed+tSgKyvmTjjz6Gwv1K7JXoyn8I2ksP3/TBOPR7ot5pWS3Lw6Kh9bPxyh8PINcyPAsD4
Gfyje+WLjrsXR/l00qSqSxxKpLReo00EITQLTttoh5Fw8jh+rreuPs4gQlbPKtHK4ajTCHsuY+xw
isnGtymfi2npMskgFA19bKpqnxL79w8aTOKNWPk71mm6rq3RjgdbWmCkXq7CwNiXkFUP+5mcqGwi
nzDlp+RsmxdFCiTfErir8Vv77NUNcn0BbMbasA9wCBW9WzpXIXm05aH45K83Tz07kO1fmtdIhOzE
8E/QYWs3d5VIDq86td6V1vSrFZTRtXwiOYN+cU4yxnHz29MWXxbPa742oTtO0PDSGsa2eRgTsOKL
kav8YzvTHf8G4Dh1nk5Kd9BeNUNSM2mTtle7uhfCc/ZXavI9leYO42BlUfzEXF9CMp+5EA2H3F1C
xo/0Dpk92GjgDzeu+n0LT635ixyxWszV9Y8+sKKdfdP8nDIyyAdN53a3i4RBCfKY+Gx95oRBP32N
6x2v3zulh25xDQjOyBBa7DV9sO0uUewrFTRnHpgleHfdeH0QwLT/4t7Uz9VXr6eUWLkNwcVD9HBd
7OR1WFFHNkbTciykVHNR1hcz6N6UxZ/mVvSeWOtNxBypvxWy6BvoNhM6PqYu2gjLjMiQC/+bviYT
jxD+VdxFJ/yHHVyAZL5wz4nILbsWlm3gARrFQSMf/N6C1OWuvuLFi9xzHkUJ+9D4rhfUMAQD+7Cl
JMQvjEiYT/axzTFHLLke/cNZ6YhVSNtdsMqWhkxgMNCthaDUPB3yWxUhdLE/hWrjMQOaLc3Q8lmC
94OLdgtgsoov6XtQ+gi48J9qwW8jgfgvcgKqdFRFfBdegp4Q+YK51B/70WJeoVkmFnnMN5u6AGKX
Q19J521OfKC/mGNfaTMD8V9TIBtS6LnQtbUdz0F/gv8j4XW2TnfSYpPfTZ63QstWvkhjAgUf7UUg
GPGEAppx17+r9i2bpcdyS9j57tUVKYe1vrFTWkJuKaG6wF1Dhxq0iqY6r/ZWvSTxMcUIwgLA+bBf
ddYLWcK1jZL4em40RroYO+ljtsfbZXciEiKGHiaH92WDhEB33CLr00aJtTYP6ulOZWyEuGzfQCzS
DOsZSEP3lxioaUgN60BkddMZ7mdpKTKOICHE0ZDOaZbfmkSRtaE+30J6CoBh6+9ZT0gq1dGD89IS
gVeJ/n6NSbTk25iQjg4+HSsWVplWbz4f2cELRZNhS3zYPFdltFCotuAV4n781wFP8zl8NoWsF9eA
5zX0bGBmb/LfmcJ0rR9NIvSKZpOuuyEvHtT+qUtIaJ+ukT0w5WUetO6/ixyygLgvdPOu+2F8HWkD
586WkLog31+3o6RIElT5333lyNuB5QXZSgqXK/upJHhRl5eghSfb46l6j1lIiTE6fIbwlVIYxE/H
tcj0jRjF9VfIbBzf6Iikh79CkMWaZuQwpwjGF+pCLtCiZZxygZM5cfw7qpC5rRpBXH5xHLk9edjj
8FqgZHvG8rO0wqz1KrEZJvy6weG2mBAGGUqwmwsPCFXDSOOCK0cXtO7+pvszR0622qU/XqSZNwIn
zyYiQv89PMA6zOnmKAbTj86GuzRlEiYkl2cnwu4nn2T2oV/Uc/zXmVEoWDlmOyRUUjZvwail2+zt
9h9M9HjymRmDP1SQMY5Li42DqZxGW/inK6HdYuvBs60h5nTZliaxcMXxxENxegi9NZcA96HZfYiL
qu6WzD/Iv3MGw6i9xMCcmVawPxbHH2CP5HkBzlN28pfdLG2UfZqeGNdTHTL1SM1Xszia3X4SL5yq
HnWyfE6x8rHAmiPpsYoDdnDNe5ObRbLTVR2OnVUjQJ7XmF+rU6gTOeEhnvsfUXDsmyVjfYiEp/Vu
dqaHP8jT1AN31KMRi8LbT2HQpoyqBEfGu4hGnwy5P5XLXWs54a0HI1q5p5/+KGNlIH52oY2Qklxr
CnBjHLuLo/Ue4v/npazdFORPPu9uSlfdkGEs4DxYaWgbqMbtxXP9n0a1DISykKvnVGzHqOZZ9oFl
cXdfdP2Huv2mgIF4hPxbmbDOokWuSR5XS8nQBJ4zcmdr/NtLUFbEq3O67WzHl1Mi6xgCr67j84g0
I8vmXDjKHiVN6fBzu3wnh+ZfUt735qm62Uu06fUYC6KVXzk4lmWV3rQZCt9PPdUWPHl7MlkSPAys
gcVCb+94JhFb0w8EH6BBGZRfihZnxlJUtHlHDH7H2TOmr76T4DjB+EgZ1Y0Wbe0bx57oPBAkVzoj
1NvszQMkHizzEWSuZdfmidik80ygz6h3h0JsO6aw4UDwrWKl81GC1TcGbVjd8/DZ0iyWG20xROOY
ESrVRq9L/sPreoJPUvR4g6DOWUMArn81L+BG6RaCe4ffEJGguRLSOo/X5Ul80thXtn/Ftg+5ItKT
7jlM/XpHDwNPYssjr227THUnVjtYpui7RTmHibmjnO4OoQOyqjgM0krD+thttY5iM2MBuFRlpD2i
FxvoUoeAOEUv1f7JuW7vXqGuEy0uymL4jqQbFmC1GOaKjYIYd1ebASWMnQK69ogrVtZVCxpH1Uq2
7co6/YaSxQogqQxzxizsCy/Kkw86LzUDHImG6KldDiJWy+0RNy2nZzahf43DhVBMFICgHUcUnnzI
w8xa0Hm2R+GZ5hC3Rb7bnf9s53yEUpMCXOitzTslrMpSLx4veIYHJpAumcEeh0lvc2qJIRwNuk5u
ZGB9mMdP+muq5ZDSDnR5YnGwlRXx7CUdN1Ns66yFkZBdys3H3e2WYpIn8m443XefpmrVNZMsTEkY
/pODqXQ4l0ATIOjKpH8iIHji1uCHY6hn+NaDsh2F7vXQFVgz5+B4W9X7abXtpzq3W/zvmj9xk5ZM
WfN3uRKh2PxxEutctf/obIj0ToUizMpwd4Tu0iv0m01nPVVY5/MI3IKMeUNnt85YPI/N7GIdLW67
M0OqWE5KyuM9WzVDF3ueYz5YyzaPwhI5ok8z4e8FOlCSKaMQkTdNkBuK4bYBWkl1thk948URWWNL
jjANlFV7lzSrzI0rXKwKgZMOq0TQKShRhyKPjTouet6o9l+rePuN5Wt+BPwVfXMOjMSjy9ERziRA
xMA+XKV5PFOzmijKr7+jjNmadqnaL3cRlcOAzUHeH2lalasHHPEwGBpgfYt6OflTBEonw1m1yO6a
JlKM/F/p/Vrz3ry6kz2UbH5j2+VW6WNWVo85OqowwVSKk5LuzI8sul6kQOp7PRldh/VJMEPrj+Gm
BS0W1QaRAX4lZ0aj8wEaalof3YGbgjY4q6WqLwT8gVzca5R8+K/vEFcENUga/AMDUe2bBp0SnzVB
rRVQs3Km/olpZQgUlsGDpjWyYJMjgM02rkqmr2shyKzrRSQ+I4UIpVX4vWGIMPe3Qxx93HiX/xX+
REn0yJmkSNtorRqcnFANNiJ1B685GNxlyvj9QnQJy10B3laqvmQZW8j460e2Yn0HQAvOalWL6gI0
PQZBq/tpVOBlQdqcjEm8sXvnRfIfEG9TgLjpZaaNaNKSF1qCTLmoqnYnwrzxCOKS2p2UtV+VaTRA
A8KLNZR6xrYvJnS2GAKA2KlitDES2T0995r2+sWoIpESp4MasSIWHYcvA+WTYiaaZ6xuaRxIkuMl
tawBETJQT6od5jcx4IuBOeEBZmU314rebygNHElqa76JCFyUJdGzI1iC0dJfDyKElo654W4Dc1Zr
/Nx3R+qMpz2UeA/ZOVIKPMle6WZUHt8lHSrp3/2W+VF1Pw1XMQwVRD/6hL1EZzKHjEZRdOHsImBb
IWg+rkRx9XLW0oK2Rz5xMdD9synMJbolNeO6dVotJXsF/ZlYWvFdGIO/kY/ctJB6kBKdVnVTitYI
X6OCXkfPfnH7fW8AMhVvgbDdoJsH+DBKW2Q1AoMfYOoavDBVumMcImhy55jpu0dLYZKypAfbi/Vo
XbOY7RjfzGoeVX/1h2jm+NPBmPfNvCdNmkqghm1ZalzAabPEPwl630NxWGqua95ny0kAl0Czqrpx
lP+o0F51gK7Zy/5R2F70L6s36+VOYylJVwe3Kwlx5uDXbfnzmdnhmMwCH4UeXU5+YKfYz1u1mP0u
bXZ5eVvGr0r73VCBrMRFMdi0dcF1K5hIncO3IVdF1ujDXfpzr8D0d1lNN2ZIqEpfSkorMql8tz7Y
fH7bscANyvWCF5jbWYcJwXQZ3cGShEgs7F/shai2+SdraaCS9RkL28GbmANgV6Eoju6pXd8ufCut
pioCnOQlIJ4o9CccMi9msLWbKK8yZIiEiFk0Tv1e7PMTv0OjB4H2dlLJKuVT4w95Vg0NKMjnC5ZL
yeIk1KO32qKgXrmp7+uAXhjExoFzVuHFImuIcV8An5qI61GwM8ID/3wbadF7mErydsKUNJwLohq7
dcDFPODvd2Pd5ClPQQpJDnehrHALdmwkmHh3xyv5jq2Tnl/GB4gDLpLKK/XAZ/TefiJnIVcC1uPt
ByfuB+YYcexsWWQ9FUcnPlcAOh7r/Mwyf9qSbbDwuDUuhNoojpkaV3zZvG3+iNreFrMIXARxai53
PoTm6FnaE2CBI40JICOQtdrY7bP5LpIUPAZQHCS3iSw67dzFPPFZBT0sFKE/hAo0DSc8L3HXFLld
bcSNQ5Cfh69Oei1O2SFelMut7W9cMRbohk3X9vFevYlatQOa+ylu7H4JqP1zkIQZxqlHRqv1prmY
L1Gla5GdMXBmBp2jZPj6RNcUViprSz9/I9Jwx2DGPkMzba2AK0FNPpY37ahoHkNB67qfsxsFVF8g
MoJWdToZaKAbYCv3Yovl6Y7Y2sk7Eeb0z5zluPG3cEpqnI1sy36V2pTkd2eMgv6M++KptRAbZyja
9gH5ZChGW32kTU+sj4/jEW8zUyysb5J072XTY02AQXfp4Vl75i21xiK6u6b26IKvIG2NI1rroCfm
STmjEIn18OoskliFplnF3rF0I3wSZEuSqyQ0KtYtFGI42zIVJ+LtdPKcGr/ue0h7h0CIigUDYiR3
J6zimKWoPcaWMZ4SKOqpYrrMmqFOrsbPfIW6wPKOqMSPqelkHlCT+rem8VL5rSAPZ4sZLcbtKZUp
KW7DtwAFMvDluoOC4fRPS0i5FrEC0UFoahoCXyQJh2uvWpYsYR8mp0pNWa50jdY6xQgx3QoFuuMP
AqTR1jnerdEYchUT1IsoNPLER1H8g3NWmy25skt93S1c7NoFikBjggRRehXMzZhKDvq743Pv5QYI
Ew8SNCy/lmHiLae6muXASPR0Wno2/Phyi0d04QmHD5d/w2to8nTcFvucm6NQohyL0z8EeF/qu13+
t1Ki4UNamCrOAg3otYljs2FgdINpv5M/vDKLaZ4Mr+WmUtapeI+KzXACndCdpiuKPnRDIISe8KBv
+EgaoBOH5lLPxvzEKuyghnjelFSQW6PYmnd23tsvbaWBuHP7hPTp31pmAK1mv0rragFDo90hU1R9
VmsWCek8PBPXX8UbJ3/W61yZ7zF7reI+O3faW7Ob+1OU8uKVKBVr6133MU5MPhLAl0wkI4DF+oFL
wO0njcJShkhiwTwwHJPBvJVydrglDHv6hjbHEdfUixHcjeF4tE1whbQ6iQIxdSYql+d0RtAw5SwM
tfoxxdTHo+cdaGTp5BYb6Wke43ZICD1uyl/eTYpfX/WX5HXSZCwomcL4jEKX/dTm93a8PZZWTphD
VQ7Uzx89xrN1Y3QXoqL7/wRUBcLogIzjPF60x0Zr9d4S1UFwIwzPjrts0Z6uPkQaSG7n9mjRaexY
Hi22zn6PSZm+at1QdyitqM4Ql+cLQ6wt8eHiFIC/a+xxQoLguvY/Ud/Og3AYkXp6CDJahV8oeSnl
LWH2+NJC1cZ7OxKRDPoYVISxh1Op8ik7kDPNVHsONv7UxIhhQhEpAH9h3lUjYuG+aOz/kmG2DtLl
2asl4/Zt4vHrMwlYx+EB0CVBarehfFSB9AqwnU3hwUnfzIktZcBr/HmjNXTz3Ku3qoJUiIU5czGH
o7F+7Q7bUdfNkfwJduyz47jurNkoTcF/t3hhkWalP8KBnOg5gmLfIp5HsdLOWGUcNuADhqPR7RH/
LFiV6W4Ny6hUl2iBvfaz/g1HjTAAO8/FbOjgbYcPB4pRhGkzsbfz3AaTnWD6K9Y7uWEogEpAeO9l
LnNNG3wcnOUEzT/v+sOYY6ReP44H8tQgpJbBrvK4ABkhJcOfKGWLgo8GjcT4c33mbEY//QUll4gx
fRBytuag7dB7kRlWfyeo0JxU2CaQjcXSI/YCVeT+1HISDCdytDoYx0VwciVuFe+S+2JlUGeWxR5+
By3L2v6bCEUy4bXCZho1plLyZrCQXPmTdl+8/4xhmmaWMZy//lP54zxHo8jzevaYzKFqiPISf2vj
34Ilup9pylD6XXtvY/NQMzMsu6LOWDVBZM4Ium5YEceX1vcA/EYqguzFNfYnW7+1L4nDCpdE0CFl
KpL5LXG1CZ/hGS+BiFzfAVBaFUorJw3ey5ean06oAerUF5ENwvYPAQwxwugKqhT/3YFRVZyDWxBu
Jhv//XFV+bp73LCXDUTt99CYPIraIZ/cQIbT0AikeY39vNoyQym2mB9x8ZIW9tCLCA4Bs6jEa+bh
sflQkkjQiVWDfHAVGXhjJBzrU/44fqdAtKi6sgOrjPasMIxg+x7Yhkut4Ft7A2XW30oCciRP+8Wy
N8zpe43WNExVsUyYkgGPSuMOs5d05QXiC42ouKDJMtcqHlqZt2JXmj3/1YhD4IiH7Twx143dtcoL
a9eL6E855vTse+srJTxx5SkEcYtVbIXSdcEo4WuCROoYXkVjOolBpe5r5cZk4BKA0OjFqU9qKGD0
v6N3qCS7Ee4ZrtM8hEcjAEtAFy9Rf0OwHbKz4yAIk/+tyz/NocZpar4rxyXVEiKPN8SOpL2bIkh2
IMq1U4KfSDPxcvQCL7a4+GY0EUPBLFmJqE6T7G6c+kGn65doDgatxXzM/XxIuW6FihFOxQ9HVM1I
4yUAMj/zF9EeiZTbNL/nc+Pskr+ekIz4Vj8ErjzX9APhQ4ImUuYItcZudhdY0A3cQn9cTBNPXiPP
5ZCi2r3KIIxrh5CmKACoAOcLOIXhRLU4176DsM8SHyprCypj+3uBpTUj+S1A/+ahclO5qSyup3Ra
sUV+GyXiW43u7a5OeqF3uMmsBxQhtEYuQ2v48BTwfBnXcy3ZRDIyjPztIOvqEX77v/fmpEm6dHEY
rQIxihrnxyGjIUu+J6/VLhQXYspiWG/eHRnYbUIBmqCso6ukpy0DT7fFn5jAd6XME3tSOQmZm/qQ
sorHncEZElq6L3T5+DOCE9TThPhAhXO+0qz7vChoZnsKe7c9DR0okN+ewHOp1TXyUQw7Ncnqb1G0
o4wQ3kGldNsBhg10StNZ00Ih5di1uWblxs/manQ6c+o/lGkn8nVb4jsWIRuN5gEw8Ey4ZaBDUFLp
Xwr2cOePmsdyEyz88U1OEF+4PBeB3JUDJ7VeS/WXmGSZUhvn1TqkXutFYvyGlpUdJ1QbBgLO6bNb
yqF1WsXC7Ef9KNx3ZWIuHl9EUnJIkIMEfEUStzSA7QUU3+X3hkc1FV7wFdeORS2ewDDcDN7iU/uV
CaVc5aHmEQaofrUgHq9WLXkaqUwyEe0Ok+4brLwS8cq3pqIdQWbWfDlpMn0iMJLlxp6ixNCN5FyA
E514nt/wlEV7UWyumAtOHQVim7VRxVIpUMOqVqAmtk4r4LKuem9XuQGC3++3AW4NJpHbJXh2mOce
TnUpGZOS1tHmx9gyd7gWy2m8VEL2rxZVCTM476MsGONXH1k7b5LjzwbFLO6N9Sc5Zhy7PCFsVH9q
1MJlmI4SK1CjOz3qpBTDLDe+vx/2VpRq9VMLP3QQd9u6jZJ/5P6YhX1NQbLryyZXulWBM0OMR8Hc
SiRYlWs3/USWQScFkqA66JDGot/ulE4TZIzbroBRvTzAvf1wfQG+6HaIe+704gt4/8cPPuxgaUUm
ARbbnW3MoAv9aeZvFrXqyGy3oqN/b5g5ZYPzVEWm+wGB9fo/MBLAZSCfii6I04bugoMtzR2ZpvL/
xCeL1vp6U9E912V7s3W4y4Ezlup2HlmqANO78NuOb+sio02IKfStJKv0o8jNMWVuwy86ufkTiAUQ
Gx6wJ0jTjMVzEPegl9gTV/2tQkitVy486EWKtTJtbj8co6OqXS7CFLpqniauYMgVZdl4V/q24pvg
cnr20ok97KFoVTnX/TGzsdeFuJsJ8OI/DqEJv/cdgfol4EM/ORatxRc2up5fRWlXF6698is4eUZt
1f+wDSP1oRySeJLu3VHR8kynoNjy87xsHGci/PLs+vO9UBq0wCK5SxiZgjfvFY8JGjw5jNz84dib
Du5m6UQgxv1qMkeX8hcZHOyeCrTQkXdlHhaylaYQL3aLsS+C8UBJBcDIKX7ME+lZrpckhdcG4Xvr
eKRj8mD9ia+wnheR8Cekp5J75TJxVorFWlFli7hBE1JyGdi9tG92kCtRMor6srFWDrdO7bedDUt/
RRtG7X390AsBCs/bTP5mzQucfUkApRe+WvGD8S3wECFC7ovUZL8MtFXsmLK2izw7u7+enijY3xgA
KrAHgCWAxr+Nh9opH6ICXFtyWnXxMJB5Nf6VIhy1uHorI/CLntqnllOn8/NUi1ClcYbNvNiHk2Kj
1czL1jeILbhUvNejOGnwG6IQOG6ta4qiyVim91alNngSH9lo1pBYwteFYXVZPxxlQeUcZQCTsF2X
RrkOf9wECcPYlKO0TZn9Bab/YmS4purso7Q/g72MlebisNQK/yhsuRlRZ+ZfyPonvsjzwMYrhAms
yRAjA7C33e0GyDtqN9x6OhCPmfjA1rMclQA9jqWFsGWW+QI5/bQdah8dYpsginjmTuQDSCYAKa9y
UFcWvBsLVB8lx5AuvS1n/vZFhGKnWatNfaYthlkMuYRbO32MM85s0lIf6Lm35MT1A8ye/cvi5xfX
uDrglUkmEw62sNoQ0V+u29Tvw3X+L5bYt2b6RryJUa48rgfMnU6SIwbAH0Nd7avXhyS3AveVxth3
hy67ROQcveU+C0xjJ520i95YoznzDIN0cnTS+66dukjj1WerYz086iXgysx7RiwxSXRqcV1SGUK0
7nikWlfrtopB4oXb2ivXljyxG/kYxwqjzDEUzPRTJss46B+IiT7/5y2SS0YTUreHu21609CG4fkz
PUFVzhhbe/9plgyiFx5e6sXso9/jUqWgeAUzCVVRpwFvSNqWghxXdiaXNvBkKzNouwcarYsofkU/
LYc5qRoufdJ/FBV6SY/56RymMO3tP9C1Ukv3dhOVPiPHBt0o+OR2B42NtEL/OOI8xiLEucRNjSPQ
BDw9aMqubn51pKy90XewnE+D5yHwHsgnoBSJ0K8lKjSfZKD8ZhIeHGIuupV2GSzEwStxU2Bf+lia
y15ytOeeWwIVIomXWTZ9+QuaKUI24Acehhrj7rB93aHmzKHKKNeDJUS1TbvCuPUBYmBhosJg/mu3
IZCknwN4HE2aWPaXuBjJ2+JYXCz/s2xE56YXMJCSgIvFgEpP8tOkN5zNROKIy75fCqJ+fhJT7TK9
4woDfV5zFO+07Hd4b2xQGzvE4/HzIoR+Tgpmo31HXRkA8Bk3LRIvC5Vn2sz3wqCjIsrvJaxZmCDf
RJOdTSrv0B1f4ivjT1Oq0rzw9trM+up62RG8ukd/NoOQPm4rGbEmKa+QsURvB6uFBi8OLyajEuem
d+pvectw898eOgnvbPUn6yI7mQQyZZm7YIQocY0amXau4SbuxsO+jz9l1nCRDYNPXuXQswM7SzCu
kZAT3Ly5DEMTnqOkQU86BjwzADbFGd1bFMDkyhCgE44aDctjlQlBO1Ki+DmWiYXWSpdOvIo/EHB/
dTgyh/IpAnp7q6Hyv0MR8urVoXxv4N4rfWsJyEWK+Az1aUG5O15BC8FQcDGDiLqi7w+JYaM9DgRu
rOanPuUOXMddtTF8BTtZQLJ9TYPpj3TCP/RgRmDERXnqGFuRyEbPXO3i+3BttZAGeMaPxYXKGQoc
WbqE9lPtJTDoQkWll2mqQ9d6sKjkne6exPOUYZLfOJx4ZqIKyf5bllreiJXiU17KJ1jFNBOfE3DF
EyTvdWN9OgR6krVoUDRij70pRWsKV+cLmcnUx+G9ijpp539V5qWz800pbd81Lj5D0tfXhA6/dpFj
+c1scwqUHdWUcDXwbQ4EUiGTi+Rrr5QfyPNRXu70XfjUUD+w834gMwDTSCb4OshlwuriQOrqd8sg
9V7dd8pM9Sb5yRnp6S/GdAsn5BCkiTmi8a+ZjHkbx3cwNK2qDaeZMcjF9bamgL+b6UjKlpW/uPbI
ZgQrgOySyjc8ByJ4+7XOxq4vDT1m7B4mOsyFXoruPK7DyfrakMz/SvR0OsFGDtp985SolTrCpZ4P
Xb4tDdVnL24Hho4Gp+6VGMeljvb4jJ4F8+XmRYJtoRSDAcfjGd+7rv4pTBlLJ54ja4qgtlIFQUC1
SlHC+Upd1gwe9VDgARCVPyGSz5x51On7nUJ3oF99MDhVQ/645D/XPq8icQRFZ/u8FKcI94QYZpfR
y5LC3cV9CY90Yi9EM8hZRlkAdRwggDyxBokoilUhaCu+THRaH9ehLSXwzHcHnrl1owzfWO4gkSnx
Ve0KWQ7EXhFb4vKwDLSpUPYl5eFpADRMWXGJRhlzfyR77cLwCJ3PfKIzruvZKRXfpq85DkTlHNEx
wVM/Bcq1AZBbxwj96uQi5nGvN/GddsuNydMTAK9WZJLM4rq+4AnP1l8FXM8vjo5pCNvxcATCGdJI
c88O/T3IwoSg0iayWUKsAAUZ5Q/klsqTcln7pSmwSRGxvPZkAv5n7U32mC/Hsvb2Z2x1I6qyMz3L
wC0Y0EAmAlqzP52opGDos1+0Gw8SkTOfY7ph3pK8itM3sVfeePM2rq0fG1X5yswapXzwYgyl1ym4
CHzBPouG074QELdC9ZPpZya3AfAWHIg9h3P1V7bRDDxEaKZupFBSjmwFAgm3dNDtRS33WPNR2+EH
50zFY+3jyyU3SIahmRy5WqHd60aWL7Q/N1xXWflVtgSx08IlwIs7qnT6DtNjXX2NtAVQIlBUyRUL
ucjYDGpUCGx0hWQa6cnW0fv6ZNpiyyOUrrUynRWg8u5Kqc+awTQREYMpYUDaAQmWO/Z2JbUiEbCO
QjG8QNyJzzuX3xqu11jMFmggXfI81Che8mmvZLF5f2tCsuAzWE7RL1D4JJO/YAv8xrDt8EShaX/H
tOlSu9MpI5joKIgneJPuk2MqxCPo//DlZHOIIIjcsD+3hP3DKz9N4i9Duo6kS59NYfoOS8FVH3Bv
I/Uuq+uA2EmwKuVynFqewlh0hAyTlkyblmAhaby28F53ZKnR8g3Oiws2cBJDDjifAS86gwBpcgzm
ySSetbLiAqjkkvWoRXbOBnBG3xNryK6C3vUB93ZoUTW5JkseQMxo0sF9QlVWBmebQ88Hl/CK+/cS
iePnA0craipfax3CHN+TxNrAiroFtkNofuG7sj9GYvNh76hab0keyk8nVgG9CKYBdlfsRQXIkBMm
agYRqv8y25ghvNrolbYnq5FcYfjpczyjCevzZTBQq5YU4+pRGLhfaaFryTgYppLLcAMI08kzk54K
xKeXt8rFfv+dvVyVNnYrEKRPQObT9eucHfM4uwp/birwqwbNsOFh6iLIshZXcrlcrZlDTeJZJDmk
yki4avD21X9mdD9QY6yv2dgJ8REv2RCWCnza8Fmeclt2ufpDwh7F8g8AeHXkn/AGLpaJGW0JOkZO
pKXtG4gEmx3ktXAxD+4RqomDE1U5R9M/Cnmekea/fmJCXlopZPB5+i0t7o/8qnSEvN62YgtC0Iuo
N4OTp4bTiYktd1GGeirAds1QFjCzLjyxZy9LbevYdGKB8Px/HyP8PSjDQC9loh+4m23T0mv3WF0P
D0Qs1BJ3krz3BJq/XHg8N0iyanoDoaIVDCymANT0vFmic/YZrpJPwDneIOCjQISmhHl/Kmmf0FI+
XdvSGM/3kYpy5JxHCvlRmuz154VL006MeVaLkKt+SFL6b/Xv7gczH7XSgXrlFRSkTrStUnbajcCo
B2cmaPlIIVaw7ofpUc8sgF0drvsHyVypgbsHSF+6aBB0rDiDiF9rIpIHkuBAGVDh77gq+Zjm2DHU
+C5eG3yj+8bnr1eLN5vleCAbCvyHK8Z4wNLSMTfBFmHCDtJNYblAAj5ulwQ9F8JcjQMeO8JZXNr8
vEW9J0/cXnHY/iO36sabV9aRSSvDPXPBO1i4fOUA4I3ei8L9LUG56EhlOx1gUW66WIWXWS0wUX7X
Ty6mGPiW1p+CteQXxC8FlWd9LpH+ZpOjO+zyfyflwM84B6zKbB1wDHpOT/QF3rXK7jvFRaTn8Qef
6F5wYgvPLG24r+HUHjzyv6aCu2p/8nyeXcBGTQ0cANa5BT+vqBD/ObY3l6KssSgUMWt2KEwnQvXU
Baco6naubL8GYlS5jd3q1z/5GjcygoJH5M1cftA4IRpjs3HNQd/Ow4AIx01G3yYyM6mATsWZlc0E
3I9G1+gVEwiZrVZikemE1F/zKlIbZYFrM94YLlBq7OBtci23jhbeIHL3G7TTtxxUMLdP1SVnGrtc
vaE3E8iQbLVKCfi/izofI0olttFb8hCd+VLQ6Z0sqeiq16dQM3udzy411NL2lOSdh9ywdemhgiaK
p3DId0eLxc2LWHMnsyEZhSimPlu86H+K0rTYCXQ/6dE0zgXxfcVZHnFBWS7vmtwhuLUIz91LTo+Y
UVtMZxY9KYbozEnbNrBANWLSmPHUK0cz0A5frPFljhtpCV1oZ6X9nOVCmNzVnJh+/ENdTvIVbHV0
4MZuez7uuyt/WYA55QBUlVPupuTSywzsl2atLUaQB/usNaAaRzc2E2XLkuxOR8OSltzIkpRNX+dE
ts0EscpJwMxrnYEhB4RUPDQlTYET5+CQ8Y4+k4fIoatX98l39RAh6FuDfQ42X07oV9Yv1/b6psOZ
ZZFdF1fpgx1yKx+7nBSDlfwCc6QLMj1oD9+Nug53W5WD0O+yCh/jY1ztpeLAHpEzduzVNgh2+Wlp
PuMNvvOCjGTFEtQkqIFI3njLZfacDzUzmE/m6Yb9RNXdISNxmcd4J6wPVAyA6mf1NUVPoBtyaluT
z4jYLdrdpg0hEhO3PCyYGcInlFlGEb0+8uUUFqzGvx9nBO+92ogrTAHZHSCQoXpbiIUslAcbq1SW
Vr0eyPT893RGrzX/6wjuUE6yAWIwjV4po33CkQCZiCBVf00RofxG0EYHptB0pu/NTIv7M5atx3Mo
1c7G7SwPJDmeCN5MMb/Sew0PIqemiqmY/rWx30Y88KLjiueZFuorE5c+IRsoKSDV4twgAI0AX/eX
OzGDoq+rdt2X+zg41dMUtJ6Lfc6wxQZ0SLaMplnSvPth2QV8r7ZZf3G7va+U+Nwnrizb+ZAGnDX3
UsdpAG34pPTengAdNzpqhBGvRjwJgRFBr9wZEldfSwIL1AHbQZ/XN/U+NoP3Vq+mKkBaU5GEWCR3
VkGhJDaZrtb6Fl+7c6cO/eS4uM0ahSamJoV+PsBovSC9Z3Go1JvmjktIkPuc/Ocl+k98W5fCqwHB
r88jdXNoX0mXtDIAAiPXdyQ9eLwIidH2IreLvvX7gjJb6p/eJIhglgP5fDiU00s0iXtCTD3KiEcT
Hm7f+bm+TlrF7r5L3iBevRgcxSDwl+UShOVcoH4PexdWP5Ph3xI/5drEtDYivrehudSkj7SS6cDk
U4lZzxOPRcIfcx0A4DoZeLTrm01NRdAgBwSTqOTsYPmhPNOwDJv0v5dWA8lmFe7evKaPS35FYTt7
dJ7vQ9UJFshChr3YqrhWKCZhQn8Mfmt+Yz+wP+kzOOdZMVNUEwNFggJFDdTd1Wqq9sQpIGp1karM
O+87lfMHh/8oBIh1yelJA8HnRtgf8eGv24NCWkIwXeJJVVNyGQYVjKlYEXm1XllH29u+E7rwFDWy
n4V10pYgNUu9jG77wN3whgNRff8wPU5NMvT6XZGbiKvwl5MQFJhwDf4bKJ+jwx30Hx9HYxd1YSem
y0b/DQH4zxZQ7/jxb14pdpsU2uZHbM6kY+nEmWYt7vBu3Tc2Jn8YT0Rcappm8q9NYIiizO6Z5i55
Y4MBECYAlqd+QwKn7yBF1PmRM7N7oDIOwcAp24AL001Xh3YoWMXXwWvEMS182oqnKGr/G5sqQtfm
MHNaKTb80UEqY/tRjM+tP5Gq94sRwxlyGJYBiwkOS+vTwFj/uRhDDrM5/oD3GfjJunX1UZ4oPxts
zIq0XMumMqZHLRiuBKX+bNJ4L5RrFMyUGae+069zVVO9DN8gnhWA+wFF2Vc3PdimkZsFQPWAm8rO
E6tXuQejwL1QgE8btbgJJ41m5Nu0Rd/aJ+6v3m8KT3ajPWGP9TkcEx/QvoJb/HkHfNRXBsQsJfx3
8ELLMAImmTBgJoLXQQ2J/cNqcmWs3v5QEXjabfWU2Dw9DoOSSpdNzNWH5fdc6ZOZH69vrFFeC5PR
YqMMYTTnDwG8xT5p4J20kr+5CShG4SFmLH/xosIKvWW6/+W5g02g2++0dPiMrxF56EIBokp90434
rjW5m14T62DjwP2FQfcnnvsaog928B6GgIrbSS8CQVhmRIwvj3WnlV4Rbjs9vOI1w6HjCGQR7Wc4
zs/CpyV9IfWdf/kvB1Pk1iuaIrGQJEjn+hwWpuosBsh6lcsYUCLAMPaDbrqRasb1gO9qqd4Y2Wqw
sAUzXPRX7QDwCmFTnO148kGuL+/z/x8NHphMSjo7PI3swvog6X3inMo+9DEnbDnCBDZbqIvnpjNo
u5bTb0BG7yve/RCCfS1FVO13kFWsmQCg/DOfmLsnOI6+GGdGW/HKB+LU4Y3B/0Bz47CYbdnKyG+i
i/7dRbVElBI/4WGfNjnMLtKg+6NyQIavCuWhRGBKULYN7x0eApyF8VxC6KzjFV3aoAaXDhp7xS9W
tmc6MGXnlVr9nNuV8ZGwwBsPImI6ltKBkFMyFfhPp+Qd/LTGiY044Qxm1nw8lSmEREpTr7ISGzoo
QZEASq3YPc5wS8vKQbCdu6Jh5RenPnbrzU/k1KNVCP2nzOXgJqNt5rqg+LnCK+WxKc46n0RNEsej
JwfzabalckeZ9lWqEntRfwFxjEldpU3TS3HNsoO+Wms2JllpBKyrDzfPpbBYIxLHzZjjeOIyt4bQ
JP4XO85hkrCUtkFlQap2er9Piu3ySIhAEn4qywYHVbRsJkBawIGhDIXBLhErN0tScPQMNDQ2TK73
auQBC8OkTbGiK+lyarY1SkKGeYskXlTr9tCFOR2rwLBXpupNuhivPra1LvxLpN8tLCRSU8+BKpNA
jFLDtRpje3+0GN4N1VHUT7q4X72MKcpiPK36GsQ2TkeOhhGgpuNr4xDPYtzEPOYeCigET2cVS1lQ
S8g2LRDTqe8BgokZYuggzgpyRYbTZUJ4qoxM7NsX+NwznEhysxsfV4t2TQK9/R0DEn+cgxZ0I/TO
n+IgZhRnYmajWZUf2wtWGEdEBPSATexfKnS70Z5Bc47XpRPwXoF9wYqbPJ+NJNx0hB0JmDwzldib
KjpLpzZt2nzsUYAmSRhrAPuIVheQShOQGoriSNNaIikHfMsog+bexAgzhD4T0seTX2xWO2FHeATD
GjkghGvjvaAXBOqXbnqh/cDNQGl4gYD736eN554YGn2Km8AYJKWa0E5micNvVFqagJ2HUCNMK/8v
MiKFALRVluWxRPB5m4Udoco6bQiXeQMhz4az0XmXSdWKwkC0LcJSjFEnzvudFGSnGH08RuwZ3QWc
G+/NPl74WjGiaI0iBPSnO0YlyN62CALfQrpsOfYORWo4o5+CNscrICOmDaRy+S+lLhMeAsbDIMSh
BUkRKvF064lYqP4lwP0BIeROEF+XoNtrhpB9WNBMGYd2CB+Z2Fk68mecEgCvbza2m8TtMTrxCtAw
mjJ14uArta/f9kvhsGlMf5/VP+ZybJTULu/ohMsIji4PvcW8/afNiVcFiohz7zVq/ErHabwDf2wz
p+9aMnvXhmKX+5x8KinMZ88GlftG4B5zDorxA88mxFHL/DJ6aTCDaMinrbd3SGw/jznqUbYI14xG
DLhN8OYVvD3Jnd7iLGCBsiPWygAoAQ2GNTx9JgQlkAMf/Dwmt6xS/MTdOoOim72Med+MCNcsfy6I
morYUygbUfTLK1BgR5z3bjEPjCZaRCpQh8es8lBzp75m7lV/jVsonTUa7cvla0XCx5GNOhLjn4uE
3x3AYLjvPwqC4jEG61g4oZQb8gyfAD4G5mPyZj+oe/8F7gMIY6FToEyEzXsPdlnMP2puStaFYJVu
cnN/bmsGPEhZ0dYefQP9+oe4i3KlIGOvjTgMk24hUEeUNVYX8zEp9DAjv1yIEVq3RZpuRbay5ABz
0J0BYIxqFtplJiXc4HUp5lNdiZi1iww/mqgUzlYnqpcTbK21brGpQOMw4Ab7oQuvmrUzF+W6zPNP
k4Ho9TBzHTeOrHWPLjlS0pPMBRbkXvSjlPM05mPVJ5Mo9p1yghEjMAlRfmC6AyiFFU9T1OavZpt/
RDB8V8CwkIlQxzNfp7YlKoKBGyco2S4nGMIp2LQdasu9k+uDmyfVYJt5B2hGzxfJrH0tG1mTNeEO
6b50UpbklKlFxhbzwC+BADWjImmqv8w7OMoyjAFth1iKeW7Y1BfEiV7bf3MQyjti01mKz8zB1/jD
NC1ShR/o3Dx1FG88mvfhciU2fllMBaGdvUQzySIFg7nSodyOF4EKXsTCMD8RRrE3i7jTcM1yNNkA
OFrW8UQTG+RTymOkMP5tlZDbi+x6xan+ypz8T97rsQYhs03hFFF7kjWdW27iafMzQsAeiiwrbTKl
Dt7hP7ZxHigkhxbyVKIfoAYlLHtOBey8N4DC8bk7E8PTj0M8g4knbW7NoW4nQmMAwgUIa1xfu1Vk
PH8nwCWxfeEOm53mwhg/maXdgLmEwcQ78NTAGm1o/OJuiL16/1ENApkRID0cDxMSkLcbXq73NiRc
DhrCEMJyWCVrRr7S4B1mpLpAgRubapapDrhaKV80JBWDbJ+tmeR8iUGTrHZyhVnmPrCu7r5TZPtl
yQZUMJSlAw2GKCuQNE8OBEK2W0LR7xxGB58DgBWxbR6R84JXORPWyifN3PE8tpxcR4U2HnggJIrg
W80u1z1jHxu1py0GS0Y7yljR/FDU2a5cz/dBimLJNlqBD3EJu0zefWm4DMAnFa1XP0votS130Inf
Og5tV2X6WKoxpf+sbkHmkwxvTk/y8GWGD5nZf47ZGqXaRjiRAKDJBArWnBNE0I80oqBYLR7fIM77
0mIQFEgINPxaHBco+LYkHkSVA7F1EgBPyEd3/JfxVhlGV3FdPz5QtQV366/vHWW6lRRljDYvQfBw
s6mZo01qUBqPGZSsT1Aou8M8q8a7YYSN0pcbuhSeWdOhAAPOKhsd+szHKLRakVPVR8E+w8Pq5BQh
tcrwgtM4+jnEjpC1SJMs0TTy6hv+YAbo4fBVxWeybMGj+XW0o395cmgV8uGmseUJAlP76wAO9CNw
VZlMSlz5GabOnPYd0yYKu4ojtAtKwSayLwVd0T1gR+/MnNMGq57QTm4Nuehb+HBSI455pcTVQnGU
B41qoo2OhLf9hfdzeSeTtnVyotLtZ9YXujBVQM5iFTTN5uMqUPw6wvgV6D0OnEegcyOwMGBwCChl
6Do4KOu4QSkKNYtdECA7ZfOkohnTEYDDVLNlIyQOrXlDCyXtxOPMfEcpZeQO50rq+a+Yh9vWNdTE
RuibPa3e8gNjrXWrtmowDZNij/7W/DMaeKSd7+Iu+DKb70xlbimw9BU3x8uMPknf2OrSpIdmwqac
2ar0V+eAfBQzJE14i41BCMlFQQc8e/CSWfAgQ/S/OLAtNb2QnC92X/gVLLGa1pN07YVTVqXQ1QQq
DFvMFPqA6ykQsOX0PtSarkIGOWm4WDU8lF+9xpRhRsbNYUsYWw/U3S3m/TWo4rFdZySfcmjCj21m
Mih6RmoQvHjaHPCb5sBs2da7FK9mOam1uz+XmvjvijYn6/KUR5PTjxPKWt5h2CTqfxOtqBi8Dwmv
qZoW4/k2j7sZrlkJbmUj2H7SwF65Bq49zyNV+q1kh+5OKJ0CUQpnZa0iuVNLWMMyB0LU23/nOKQR
azj3fILJOGOJrwxiutyRx5kF7T2rn9YERWRngJrAL/d71XI1eTTwTF3RDmhnWMJnzk7GFezqul8i
hnfff3i0ckvB6DNZETpzm066c1dGASySnuPFgphF1BW7fRTNQZGcLsZZqqRevNCYXWAlJ7lNw3Mg
39l34aqwbJ7RvDaDn1mjLQGQmJh3tSfuWIqS5UUmJ0uyjGt8Nt65J3R2lFaf2svg3uL7bFiCDF0t
DLlMRoVCH/sMZyfPIgrK8MLrx5cqah8fTLUo7ygUjrxrmBEmKOmrALPv3rccCyfjGJ2TCnHxBmlb
+wlcxTkMLpw+pjKp3ItZPwl4OZXY2P+NjAGdR7NOtfpX1Ds1Ix/Jzg3sopbk7+RgTDrtuccgs7+9
qC5O06fMfuO0LRnTEUv3jiTmTfOpf1+kES3OzDv1oIyQ3tQ8Pa1ZubVjOXERnHg+htGSWeNH2Sd/
hfvHOndwOrLGj0DOUKb9TRsqqhuSG6IvGchRJOeGSJvAum8Jb+Vsy5d9Qw5kawpz34/7d3ZYrxAC
ff9A3zCnU5hzuAh0bED5fVWKecaS9vHkBk4DW3APPyXdQogAWG9HtEoQbp/XziW3JF4V3MjHibd5
rVWJzVnUlQlepBnXHzhzBLTYygIq37r7uNN28i2DJHrom0/Xgcm0F2pHD+SA9CdmaQ4IFLB1u/fG
KQuiG5f+A0NRPDsCahX7oOHjSWJJSSLxH3+PCbO9utgUqOYrAzc7hWYINaqEB1I21eskFppwtIGN
86BsZPPRYs04HA77vksyV+vq8jBZqO1TfwgnJ7Elw0+JGwIKYHlsVybjfC5OtDMCdG4WlM7hvCVN
qc+mZGyYpuYWleb3alTiT/Znbh62K3U6syRRbQYj3aaMrYjZiurl85JYLyqdWyl8YTUBK/ZzS9a+
plJkki34ghUqWRqJYyjVwrfDROclGqbfK7MYltSNI3AW80sR01yH8aH3bTEdwx8JNWjW1NxfbZn+
o70OLmoJzT4iK1HS3g8XEKNF9K+BGvcSzfpZuXS79yUjeWaHl9Oya9EO8VperlGnvfWRIHEoj1Sx
AeTjjoDlRK71OYHtYXiNA2KGq1PgRy4mvlzpK+Ax1bhDuflO7YFdUqDFEbLwdXP4kPG3uB4v2MHg
msjSX3N/VFzC3S7/K+70Dz18aFGS5lH7tq+V6zwhKyMkTcQpt/WWv5l0AM/yup/xr4Yo9lGe6HK0
AoQ4YamH0GTehVce3dSQBPjkIBBHSKLuym0wiR97Dw/a4O5tC0V7s6c5eNyx1LxP/b5pLpubpQwS
f4UT6B3l86JhVxXpgq+5c99waaeSRuv6DXroD1WFxNglvUyBsLb386Yg60nGVq+zbOEEBygxsEZ0
n60C41RJKFXrJmQzLOTBP/neUptMccULE3VTNeaVmHVFQYs7kRnclYvnl6ULF2ByUVSe094SS+ER
w/+Z1vE/LBjppSVK5j3i1lEV8uuZFY2L3qqFgjx9j65hCpskask7WE/3ZRDIS+6vDe5OQ3eaD55k
B/k0DJVRcJaGoba1yjfnqKrKI2iQk0OVE7dWE3WHI4zQAq++rezsg93KBJtBBjR+I7QZu600GnK8
4liTW9g7KZAk5av5caCXHbN8f30DESvOvUknzLyAgdehSs67Y1XmhgAYyeSPcTf27Ps05c5zjLS2
PrCVtYSWrA2nTm0khlX0U0IbTxAXBpzYvQ710BWQvdiNJBmaB7dA5gwLilhvnY4Iyzss+OAj0+b3
STe1+2y4wEav4j71I4XOjIL5Ocpb757x55aTOrFI3rLwOnRPSjwT/SlRzw9hI/eameoOw/IuKOyN
hyXRtkGsi/OXllHJxpS9Uf2Z3SVMI3sP+HEQyMHlOb1mCKGB5A1jqzXGvMb1oDstbe+RXXZ+SgqV
xntZ71/zV0b1JPr1WYkROjokUttvWl+ItCdc0kjBTmymn+crqvar1cUwzx7rpObgeY+QeGiaoxGU
P6wO3PBh+6Ks1+PLnbH0xepdT26e+PsxEiki/gdF281iifZb1uO4AB6jbTy4VnrjIAX6wsDICinq
pQQJWHzVGvO6EcdqApSjWTtO45CrwzPTyZrx/0YTxxVyUZG3kzZ9yRo1RAQIfneURwGHdKBy/SoX
bOF0FnM80v4EQklsF2odqsqj9ihXNzmqjkGCVijjAv1CDZIALI75o/RCDyHJK9XpWTysBZYFgE6Y
zNgk4ailxPnLoEZUb3jQc1yJSuuQ/FVfmaFMU5EapafYqHeMrkHpo90r6bnjnzYQg28JMo/tu1uR
4+j1qBOaS+xp3r7lXaMUTQCYNGbgSxFBS9di757bE9SM+8oA+rcddD4MqmlK7VqGHJY3efs2aGtX
ZiZbQA9VbUZSV2yfVBOJxKRxPGmH8F/lehT2SjVhpQc/lGiE/8DLD1oVQuXbTOHVrND4hFRweriG
HdMddl47xq/xsFip50q7pl66rmVUJGH05cyhfH5CXQn0TuG83PvcIc8PPYAgHVdHmy+RX4IlrzfY
Hqc+wJvtvSP7ZCA95AU1LOr8Q2ymcTsOyS6xF8jFQ4GMn1ZcZLNxTvvmX38z9MGn2Lx4/yCh8Wzs
WQRA1tIIH5rrc52Dg3tMznu4P60WDXkyoNdBJHIok2vubot5V3+DQNYC+u3pZ2EtHVzy7IvC+1To
1ci6OTp1A7BPj2a4S6wLWCdS/6Kcwu0lj9Dz2aAog/4ane/g6+lvQhikiW2w5HtFYRhAvMR58cDu
X2/SI61+UHDWgczwLTlba/f6ecLl2oMuMXwQ81iwFvcvFRiMz/5DKdX8AblMNmiaPiCdngkmRJjT
9dwFxaCtjlShGamiN9HWxUDsA3FvFpbAueZMeSGFO8wrANB/fKn5MkXHmZ+0THvCZrfuqriieJWO
s4JBSGlbSqxYFg/qd5UVSn32CHvoIbjKSGXQzD7lpnAv6P8UAshhOnoSGMM9rFueE9Am2WbQXmQJ
M2+JAz2vpZG2AsMkQvtvmD3dXh8VGFyUTle2WEq+IVTZMoqgEjYtzrZB62Jy4sytOT6AKz04iPFO
0cFrZ07mNtGBh4Vnv46GalXM4fsCG8zkQj92w37f4JU8gqKm7+Vds4jYhXFumrBOhLuzEBMLEpeH
FiNieGS3WgpQ0wZ/o1aqOeEoLPJb7939wEvDUuM0G9rL3dGr/dBhn1QyC/phTdpMYA4dep3WJmns
toGWb1SFilrTkJK/mGlVBMKUmZc0doGGggtCumunVL2PF9kp8qb1434XhycPOGQfT4vBpYMVY84+
HDgM0+Q9GSl1c8umlAmIoprvCwGnRMYAgdGYGzMMlXNVmsggOwzs4TxsexWqzONM3cv5ECH15zo7
hj4qlqcr6N2MfI3Hfqz3lch2bRTshIBeaUWMKZWWi2lAxnK5C/V1WZOc0RuzoLvLZ+V57vbebbY3
eDZ1wSvqL8dVOYCyzQ7Id8riR5im2vxJ2uUF62VWkViVTfs6EgllhZRjsXMgfRuF/Ellf1+UQAor
6becUHIJ7CYaQup8z8ubI/Q8ZKx6RgesiHdeYp1KU/P71iChZ6M5CZYD4tucUxnjj8V079N0Is30
CmjQfb5Zyt/ij5y8UOWnw2GATfi1W7c//70MexWhKNmwHCchO3qU/Wll905o3wUHRhn0Fw/oS+4y
5NZHEhRJ+jdI2ZG/BGHKuuKrW3jDIl3zs7fclweUgPdhnkuPDeReS78SMkswW0S/LO/V8K5796bJ
BplOkUMwFKT3EUKDHLzFnDWiEYZ75M5fI2uBoZ3IPDh3+6AvF5uKS1gwXh5omYNCZZwsUeJZPN9G
JXSAXamA64djqpp0ayBLsXgSB3HEYTuMRupZJNaJAUDjuhm8SXlOq/iw55UocuQTDS2cpGFI99SN
o4ggeAq1G7ZJzfQAj/FiJdaGnM5mGiWvxNt0klPgEiaomIC0VWLyRtKCyE6P4vrEE4jtx8ugTfnC
twOBNvDOJdiWSE2SfioksA1kzz/DthyBfDl0reVkpKYrwYrSBmS/6qvEYywrpPkI47bZt2YdfL/E
EBE6dc7fydIIuRKmm4RGhldRDHSecNkaXGV4Lj4QUKZWECDxY64gSCCUfxPV0v6u/g2OcZh//oyZ
45dAIZdeH5FPhHRJw6v3jDYYFqtmMU0kkmNbFA8MHonb5NLCm2JB4QHeP1N75XAc8VbWyS55ojQ9
7RYhHeVxELqI3sSWiY9jFKuew87r1gUXLHlc40fJk3AEHCcL3dMHuO/Gr0UAcwFaOdqZ+JuTDmMT
1XzxXT/TxdGMaGrjqCfEw/WQP9R6hbdyVvGIQcSlOQUgGSIeXV/Qyyw9XGcayYaiMH8j1OlmOf9D
cDfTJzOfq8/emMitrgkz5U8KAIu8iVYWNL2cAsq4O/4de9tUN0MfrEViwRqD/rodTkxLaxBU1O0M
dsvhv3IMBM0X1fRR+qv1CBL+iYcceYKPHP+Y7WTpJpMnYvrmEHzHUGx7r//0j3vSIC/krmUYZo+8
FD84KQAotDP6jURKu3eOwveejA0OVfkmfNIXCkbvSEN4fxVaIcw8vNoiFkNFS6PaKRTnzujG7DgB
/zOlhfPNNeHaaP8ptgpmbRGk03bGCB1AM2X6WkX6GRP8qqMGnHT+rb9N8hL+x5D8KhsoFYRKB6Eu
MUjMvaBJ6gEsK9euccJnWBbB+0qmNmPy+dePQHymxuo6fQAPS3GymHd5DJJpJHz4puuRpk8ab5Gl
95Z3P9ihFwEhaTaYEGIB3ederImWSJRjmk9ms2L0mnXfDW8hXpT0QORA5OEoLTayzuVI+3Qg17Pf
d0Dv4ONU6SitCGKRhyt6l0/UEY4IMhOSCaqFb7bhMH1SR7HMCP533PEab3UJWTHJujN45Tr6aEoy
+exIjddLWKdDSfrx/hF4P/J8k2mp7VzLOAWAKexVFZfsXyBYcsBzrqo7IuYpRRKSeezH3vKUevOY
d+rTITNznRofiFu/kHcBkb9uSDb8i0INsM0bCUPbhXF0NGKLc1CixKv0M1f0eyR2dESO8TsIJOIE
iinyCAaD1wn8HUIcrCXu8xHsu5yHGEKjcbfJD7QQ6baUni0m/RY3qrQMY/bzhGF5XwK7p8X8MUkw
+xU7QU6EHsRt5mLcm3z2A+zSNpWkXJRGlhFp8ZLpeg7gLpUdIMIxKA4xZuQL/7/sAFjotPMFDicX
ngnsqy1e2T+s2FWODshKmXynymOUjuVR9y1wAQVHbAr4C749BQ9RgnLuHBcYiloTW7iL+WV1Kcpb
zoODmE+Kb6p3+PgZozCpiQs3wZLan2Nl0eQDbIgyrYw0iSdRtyvYB/3F2Ui1IBOci5XeFXXwVRL5
POM7N73W5cgdEdDDY4hJ2l3Pf8+bSRe+FDBga6VeTkpGpD5afyq4EU/R/5dy+0X2Eu8ljluPNoE9
V7i3RR6ztcEYV9j4juIQ74XMgtWGNG6251qCsapZeJPVkWSLWfvMvbk8bdTbaoAZ/sGZUTTHZzTb
Xd9pUon/XaeIUiWMJ6+79KYHpTGlvc6P3e+hNdKCGueXXGXicc7Wfpw4pBB4vm92a66iL6iud3XI
ehX5gVyf60Eejwmb7Yw6JEuYT3fw7rsD/nO9ScMJV0mgvHOuz1dZsdF6dZlwFjbJl6uK6HGu2zMw
S9UDkx2uuR6gnXoBb5fBRfsk9HZQX8x9vPZUBidxNl/axLQfBjK30+6Lv7MiKvKu8qQBprfqsNeL
9EbfG1p2S7b8aNpTUDA2QLHM+WG0R+V6cUBGCpYP8tBdJzfQL7VaL3AjsejNT/p9VyOP5s8axRBh
NdliOLXwuqExsRUbYBdwupFhTvS/0/LR1ScmJIC1OwKWGG1ISJwhzxle5PPBTuwuCTgL5oB4Ftmc
EwYttG3dzmmOAMMZopwrKFkLatYeWVgeepCmaMtdcY/IfoWTLdNlyOFfIfa2ZF7aYIaI5165zBSM
uKwQxXb+snFCoBbWJ5QCNWUfYxWMbLtjrY9NLt4f+sSkrqkJvBErz02OBGtJ7jkxRdXVyfIDeGLh
oIB4fwVmk/bQObMBvJpLb29mkt3EYY8sdII+U9zhJ2EyqsjUV3Hq2nCv1CU+Mg7z6Y6P+PLwr0YM
QepP10cxtV0hwb+VfWTnuBlRe8abVZO3pPPNFE9PXAp6gqokL0A/5LitZQM2qPY6i8e3gP7wr86p
RPDn/4kRT4i/+5mCUC97wK7cuxg6MsZ0rLIp6+N4wPGNI0vz42Mv8+lN+AF9aiBAeCmS/ZMY8rYC
Rf6f86RpGRh09T/9jsQWbI2YLxg1cAGjiJQ/Q9TJVaW9PxS4aEXnqwJcGwNBj729V56/ak+BN/PJ
kFwXXA1QstRwLteLNokwL9FJBPZqFFzHLz1awQuuhXyCBy1AdkSkMfd7F/4xoXDKywmzlbHUDPe0
/iTezy9fdPjgUHCwg0pSWINjFW5O7yPtTSwXlXm4oMOyxjWuCPIhViAp/NnTsTbeYb3JRqZHqzYK
Asadd0mtsrkswxhNSeJFS/UvsdY/k3QsVdzfKhI2BomIvZwPjyMJq4v80n01EvQaoRAu85BIssno
EGPwjT1TvRgWx4dXabxj5Jdxff04q0ntNhprPx3/64CR4Zi3XosFVUESvT31JXc6upCnNmwNwcqZ
U7j28kF9y4eIb8qJHwBjy3ZOAxaisJFSxeixZ3+Bqrd9qQe6kDiiKvdkOoquaN0siWdmIPWZYFIj
WDTkrYMLreUNxu2xiTdRF9kGj4fzhrNfA0BhTcNbYDV8gzyOhQIMtR59CqekT4Pifbqk457sM17P
d5IeR5YKR35O4PccSr+ceoxNyWaOJSNTxo5DtpazdmzYRSzGDiwEkQECkiMSrkJy7J8iefS4o0sD
r9ruT+HBg+9gjQW99MJgrwCdZtXMBMiaE6lPDic9aVvcmrPo651QMmLjKbbVR/WUFBzR5tU7s7JR
WlFjim+1WshgnjoTUP8GTPmgUodNdngyjex47srTUYgV11nKiiVlWT3cSyf03m4yosKQetbdFqCJ
3thblI8GlJu97wl3zt0ZXkMFI+udLAW2vtjk0PJsooqL/7ET5oViqOrIAHD5YXBRz4C6ZpUmTQEK
08Ece10CFXgpiwNfJqGky9tj57W8aSQh1h31cpLXtlkBF0eOgrqOV6fAM10n+NqVe118zjvl7sDd
wXGFVqjy/zgULoIhPsyZqNS3sASS7XbylGo233l2ODRz8JVd7+JjbqLveTLdeK+VmdqhjsTRhYRA
agp95bQ3XdKMLfq4+NtsuwRBdP4vB6ylzdZ78LJ/Eiy4Ddjsv9AsHVOvGHFId6KClYPMaktnoDG9
Ba9cCN4Gwcr823n+n54hJI4/O3OnlSYF4ULc035S+4DgDo1ujfCDUZuZBKC/MHDuGcSnS15uQlAB
BNqHeP09N9FJmgtP8LM64zPR4g2ajjjkg76r/hAEM1XrgvGWYR0qPzyxqYpx3WOwjqocjDiA6Koe
CjHC6KD1K4Ums650/8syCwrb2sW1xoVfbulLJxW3kQ0jxw+wefhtltwKlmWVxB1G1UQEzvthYfE7
Op8KvhvjCRktIOfnSjS1CGYfakX/x2s6/Rt9tlq1YwH+2hpU0fXxfgmF4mnWWfOe3wNAocrn9dCh
j+QmJMK9QEy3JhCOgYI5y6N18MwC9afHXVyUC7YqQAoxAWXyjbRyO7EXFuTVO4ZsDmNA5b4qbgCD
EJur0v5QeLqNpo3ctkTcG6dLeAwbTNsxoHVgNi7zTXeNqfblsoQ4+dX4fDxa5nBb/Z089KNnozq/
97vnScjh/QhQnRjsS2XFe0eXLCj2cwStoj4PdPapJO8uGxbRqO89OX2Pv7DoImx++K0LWn7Ld1bK
fxHrJw2E4oG9Hh8JlFS72XofGx06CuWGUYOKKJJEcAzOvthkQlYrjQbXpR+iUYMlQo9LlY+MxCRj
2ik5KltDtSk1moM16A0Tmz6uiMt4oZyjdSGsyVERf4cjklpsh1RCvCaxBVOy3lV/zhZUEGyAPgrp
Yk/WVq97dbzY+/d8KkZOR6TbMCfMyQGAQFaATvJ9dZX266YuYD8uJU3oj5Qtx1P8bkjzo6s8ZZ51
tB0qJf0MAYCgk5blae22UuYoN7jeO5nEdfDuTnXHHkT+DkxzYj0nyVMycIJbZjtHtDcBsIYX0EHh
NLdsvXgby4c2fu4uQyaLKT4zhRjLrpb+pu8V+wGSPS1fTHHW+5J+HuHuyp3rWK1bbqzNeCqAXM9V
uXP6poPDabQcn6xY2qXfJGgTvaYWUdrZXmM0XJlXy8Na1LWYRcJv63QCx3kAD1qJNftL7MFba30p
CeCSfLWNpAwxb8+6mUsNmBxVxH0DjQmuu6q+TIZzcKMNg/DY73xdVIyNUyZetZCetkl26DPTFa24
grcSN9aKPhipYb4D67c3aGiKQoCFQkxcVA9TAmrMTfcBsKyEttX+Y9nnk3P9d/t1kze8H9c+l2P7
vln8J5UuBjVEPijVA3yr+NueIyLbTLnzwL1lek05agp6sltTq8zMXugSBQBMx9E+BRzzJ43JPgq4
b/Q1bRDpnWdonO44CEwUxiM/snDYC19paQ2rq/m2mTW7Qk/r77Ihez61hgzDn8HvWZ5RJ79+DoyC
7+bZEH3uTc+1I2adnVFAHUlKKJZ5EJwl81hLJrEKHhLtIo1YuATY00m5BWUpESC0VwYiMaqBAxgj
ni5Mpd9n/pbi2vjIjOELDvY4MOfcniK0DjCSZlHjr0qCeDt1ZmC6fv+OnjRAzqAF8OzL6uDjMvVW
RCPETNGC5RYl5KBU3NquIN14elrZUCiGz6maRIbAc5yF1z/9LzzLTiWKcbCEzjJaE8fcy/GNOa1H
C5oktpWdSl1VwIaDEsLPY8eQWj025JzMC4nn/PdoxyNHobnsNKXY2X0uKaFFvPs1xGHHpgqcdqzS
DjMvZyhWbg5yCyCCRXrmW8c91Hu5GeDRwVjwb1Exru1EBBAG2w349JEbFQc0zZH4k38SM/qQ2x8G
5a/e6fAhsbhzwq4FEFMr4cEmO5JPecn+T8BHfK+VUMoTfR1GSwL8NxdXOgfc791D/QtieLZAnuRm
fIKIp82AnUFSsK5sqPu/vCaPkr4RaFU7ZmBpjb+L8TmF9Ijeym1jmqFnAx4t740io4KyFRYL7dbU
XCptRoJlIc/2yL7dSC+WQt02UEO7ZJ8zPjmDFNM5vWFxLxbMhREXdt8TsMXOEKjrBcgZn7vsnDKp
wID6M/PHg3eT2KoCfMZxbXw1Ld/LKLnEwE01vdgz2MmlMiomzZF00knvQuGwDrybxeoH2e6JuD3D
h+y//dg0F2T95KYOQ9cSXV3o7hMbZAUBIM1s/yZwmIYDMJ+gvT2+Z4ZDRr3ZsKkmpnqWf8vl5Cj8
qPAt1hA/NSu/h6XzSzBTM73L6CB7enqP5ORMej1DsxYO16Cxjq8VPmqzgDCTiOgkTZyIHFwiXPQ4
1qpIejCQkKylW6iDNZNeUcAl/6qv1PoBEULNo4hJQXF8d/IXswS7nW7Q5MuQV3AOgniZtVqrax05
ikIN18whH0MlesxD83gvbQB9FhF+cl3uORvRjgyMImSzoYH+LxBAlCTMC1meFpCC4AE74vRSV9FU
A8uiVAhO886/FaaFEesNzduAGPudHXwq0F5q4fbkKJnWTUc8bB9yg8wZYuuwA0BcdVBAEd5dovfp
PJExUbf0MNV7PJcAlSusczqS1NTlYYoEsIcfVpI4HG/49CtugkWd9Zb2eOmY9aR98ia9Ymhu9B/F
vTMZOrSWD2Pl8uvbb+evHKdh61hFrcF+Lld+77Mfa87iB3Yr/m/3He5DWtftauHcc3EWz2hictgL
azZfUmeBPDFVKfttjZuD6vkdXDhb0CCkOwdnEKmNh96wHPb9lSosSvSLEBgUh1f/0jm5+u6W8xdE
7KrHncmGnQ7xDRTxtlTfAt6LbMytjTXeBxgP5JDCJIiDhmlBQV1J/e50t6J27FZxxtdTAW8Zghr6
yyaqGAI6nQvlUd4vSi4GyGgyPvrSB8ZgCAn51NNPLD7vRhMlyR2Ley42++RZp1IRWaEjR0h8/Pfr
jaiTnZcdliKQXqrR7VFTvhSrKWcKKURsj0EhwlRf91RbBnpPniILRazAARHwNsccidWhV8d8LK+g
fhHz9+tGueUnMk8/xrDPJe7cuf4PrdVD/uZbpAnuTzimQr3ob0qpiuZsBOxOW9yaewmlCUuXtFlO
45944108otWQdgPF4hOKWIterV7fBDT8N5cvbMC9coXw/dRjuP9+NOqcicDhpTZJHLYQIvhZzetF
6FX2aVDH6EiXXAUNNbpx21qjipPayL+wG21ruYD/spULTRSzucKE/zl6D2KI2/xgX08EuuC2ZWBS
9qxD+U3PMSVsuOKkagI2HZTonlcEXFIUGWO6/Kg6E8Gp+DgljcbZplKkusroPvUPWqhZ9Orq/g6z
uU3kJyAUe44F8aCAz6MjiiCy679WNX4mlf9FFKmjbGDu+fstbwWYP63GTZ+9VjK1ghERHLl/ruVd
pTRjSDXS2BdcjODiezaU/0lKDJ22+qg9jdvTrYXogq+Zx9yTREZkaBYFluUcYW84x9Sl0MBQSSB0
Nz9mpopvCI5xGfYUQUga///id30Fi82lqKR1L2+0Ug2f5jnTywl9g6wZRgvyyTZqwEAE0baXJhnr
j79HF0BI1I56Gp6hHX/vHR3c9aN8mez5IyoWfXr9CmqB1CWjCFPnU/cPi8mcRE4ZXAb9MgScw07X
V7srISvND1WRZz86iUV4iFY63VlWMOKI/3tHZxcyPob7KZ/b0eBMo196Fa/U9aAJIE4TVEDw2Nfr
MTMS1dwm+kJnzVqE+iq2pXoY0b91zelLTdb9G2JaGfww+Ha/T9SitEixoYr1cEU8Pe40GzOB0AP7
i/Lk+xcphoITVR5V3VF07WekBDOXZy/XosMPZtVl05tgE/QOG/HOMo9+JewzcZvC9tjQ7ec00i8e
gFVl7drXkWr5K+qv/5xCxQQEKOwGEnmZy1+8ow/cREKzuSWuW7AUxl1lXKlsUO6zSKKdioUDiQd6
aWfMfLJl+VL455MiqODFTdFFXS+ds/jMrGMzhX5bfaYUvmUUb+JzL2U2RLEKQbnGsdY8cuNt4ULB
WCTvDG2T5FJ+6tfRQBKilTgkhQh2vD0wmbscxG2ZjhLKFuhyqTYfJHfOeN2zGNx8ZiH+MAqxjoK7
SgxpVXkEQgvptq9jUcALsIGcQd3GEaFNJ85Gq+lJWim+bfn4sVnHL05kSKn0dVGA9v27+1GoYpcg
Aif9SvNrdMCQ2PAGLopZksKbN5vb0OTnhHgSfUseKm6LPicxWL9TKiHJiYwF7dZe2s3cC5OxvmL+
esFvvhv+sY0/44DqRBpZXpLmqo5zTWhKysD777AJlr1xJFDS4a8+ZAizF4FkNOeJRMVj2f7Bh2t8
p6ERBwgMe54AtAHKDaGD1AGSs/xlpt1FkgwZIXuvIUdrAUs5XlWPDi8SqtVWBbTmmD8EX2Zr1HXR
jqWYKz+JOO4Q3iwelvSxL0qoIyNlrfZK2HgVpmhSa/uOGuAaCMjImI+sAq460MAqbAKnkl4dKE2M
/GwpG86/GluBcGZGZcrGcTjBgZb95j4OnM6AqUH0mEZT+idJ7WAarcLR0Yrbzbbp17h1AaMsWzrU
jhsUlsk1/71UvqwURLi4EkRrKpUB75DndZ/mqcId2Qy98lxBP18JwxoOxlUWmXe/yFI8zRta0VFd
KMFN+5nVGpQt46TnJYcuOnJ0pmoyEMbXVHGYfFwC1vgICQmNlLCtXd0zHrC74lxCcLozy51Zq20O
2EKzxzveD1z96tVeiTieFkLyZTLG9V3o2klKz859DTP8OVqY7bjFQPIa5RRA5bh7YUgzlkSq8a6q
UJBCElZnsIm52KMVX9E9oTuf4XpHK76xpf1oqMnoYvv2lvNiBhpFm7K4NSYLL8rC1eIXO2P8vlFD
PmeQd7AFsFbNxsp0aKcu3cGJpi2eweYZhDxiug3izT8920e3GBi8zUXndeo2awiBeeSzAWBmQS32
fIPsQomPtdnAMSNPIraHdbftUiV2l0wRVBTlerVAfPBhsT4UnGrRsCcMrDv12J3v8xtjGHvYkjuz
LQDD3TPB12yXA8LPzfaK+URvpSDaRinCxe77sBiPr+527otYrmUr2TRLWndUAlyREKVnibUIJXmp
BzS7653ydi3EqafM7B/Dlo0tH0Ke/I2QHOR38cwSOxCj9Rl8D74JuoB3XP08SZsysYHKL6uWQa0k
YOwtyUFszrt5rI1TY9fGp8glpDC/z6BEYfq7TSY+gSfJRKgbb/8D6b5pu3LXSyummk/fSLICk0fu
T2iggrBkNQIphubIdtWnYm0gbUV49/BC0v3Eus8OWFIZRYAaIxNguMLNYHFatTHBFgmuZsN1O/5a
pKAGBXEzmAPj4/bRHujjtbwAuyMwrIfQVPD6mU6VLjWHYKv4GZOuRHc7Ygtriu0TCmz+Ye8K2tQx
0iCtbCa5jrRi5jU7cQGAIhLDs9RbRTN23AsTa2gUn3wIf7mp4PuabdkiVANzKYpEu8EsSlTsEbOS
4GKOoWdNF3Hm+ViWWIt7OlJcpZbh+6DjP7cTd7C05LMYSjWh3uCoFBYPxshy5GtFQEY64GyV0e61
L1lDei5vJ5HDfHc2xjt9BGZnuo9DNfabrL2acA3Eimx3WYAUrbjCAFjZo3WyK6mVpJCk9hyPRrVR
eYSPetUW3X5Pucl+LHK4ur2TdMa+kwr4grunyWVJKukrjFXiLOQ5hlO/jnpiZHVhOvoDVtoquSZP
z79stIuGDNasv4lr8oa6r91aMSpyRENgL8MIgTyl4pPi14moUwCcMQmPj60EiXjjRVAuuQUZP5GH
cQVhVYvSckbEfHBkBC82jFw4kB6MrnLzLp2QNYy+I6e2T1DIp9UwYZ3nR4RvPShS99xo2cJZ6+nx
B3c1GnxkC5yDc20h+KcWxI9/2z1UMRhxXkTjGHXyESsoPzs7ICosKNUZ0w8THAx71pvplSoEUte9
8ZM4BgnbrEcuXB019xwiVUE+xF1Dx7+10gmFxEBhIPy/TFRAIT8aLRz+4OOnJatPLwjBZ8zMENqW
HXOndSh3Cg4KM7EHftQtnQY5iYN3m70q3FTPTJBuU+/us5LL6az1y2ZsOPsNPCNBY24XYltuhcz7
Za6cUFoNhiJPNzPHpkxtsBrJfSK8EYpgKJVBIGnvFmcE1T7fJK9VGy/WTfzz7XEcc5WjrLsRRu1K
GLdsKwRRz2cf2unQYTimHLpZn6zKkM+RXzoHJWzccCseS5/R6ix6FICnKkAGBh4MaoahisFgPcUA
6cAYb7uxu9/VSfsnzQPC+bw/tAiGqyqKAMzmcyfxevcpzm2ixMg2354jSHIXbPwGReD76tUfAj+z
IUK+twf0KPmetnTaqdjwKnPd21RVoIQFxh8cr0V6uriJo6sFqXvUSyJVZ+XCUWiEQgLTQfaFgU/h
//0U4vbfK5onrzIYYuXJW/oVy0xpEX0N3SKbiZQQIlUUbI1Qzi7uQp3qSEptVME9wKIAAdvYQ34C
jtwIo0iaAw0tLe7r0hg/8Wl3HaM0d13Nk4bvWb5wwZPpfn2Ag0Qt9k37fIeH34fXNyiNPMasDDD/
BjGm0aE8TiANE3BWkArZGEcYy2BAjfURNfgmaNWLK2BBp1GC04AepHCqPKCEDNrZ67qRkkx2K31a
Wg1bphMDXtl4PhoaOdzhzl7mS3F1EQE8KaKUOgGLmDgDxHPTYycK+wrDf3EV+Rxrz10HOXasHZjP
hQKQ0EOicDMNmNpyTRA7aH89io22+Q/AswtpkObkGHXIQlZ9K3nZPLd5S3xi31Zyo2tyRPIoz2ll
iBQteGIiGFmvfpLC2HLEXvZHOkLRLRRgG+CSdoRh07JAbJbDhdmI2xKRk6ivl8gDdgRItFHVHqXH
9LVDLwf17/MLYBQPnvyldLoTvkJo8vaWPyE8krT/3vXA74r/kADOsdGEd5ngrx97c1ai0FATObOy
l++A1i0Y5bVoCCjWdg1DkzzNu/iKI4SLZpevUzjZ2bdUOivxxr3QVg46nKXhPq7nWWx6Ebx7va4u
848Z6/LzISvShOIEqebozksXnuy82qywVKI+WrUrV3hocXPAK0eGOV3mugL5JSJyGjloP/ZtucjU
0513G05K1aEN0PtPhCCTqEcfkuekYOUYyt1WJ+8LGfa45pjNtq4hkNPNaeBofnCF5Mc+hb0u4UsM
td2+AIZVz/vdMF3KpHSJ47Szk44Sg7sjj+rbG72CLgKxQuzE28++HyaRc1WZglYVT8O+BkxeYy3u
tXlNXQ+7GDtMMK+5yNZUJA2mmMb+n4ncDgJC7olGij/9FmF7g89suZI85r4F0c/Wq7WLShbMKrb1
8qqin975sxR/1OSHgwLtb3s9XTnGGLNG2PD7JAVmmyGHPZwC0F/XmUqY5uS0cTFcEiQZFpgOwdRw
mE8NpYaR/zvHZNwJzBEgo6V0muma9mPf9Kr6VckTXao5Qqgu6fWLrkGV3w5U+UiXE8iFMuJ/DfiA
mXVJy4Xpy/DTElTydo6Bw4FwF7VaFOtTAYu6v/GLe7Qw2FCU7WOwmNVhDudM0A2spOTwU324qiI/
HGae+q74a8s1JNIar9GnQLYaqMRDcDw/12RIWVrGDG8+ydEm6Di/AcWAk9zakfk8dubQAO7F11O1
kUSLqZm6dXtwGaLyqKgt/hfQkAdCIwn2RxvoxOXeW0mY1s8TH17x/I259M7oHDD68229B1O/BApI
uSY7fbPASFWvJbha1bJC32h44leZ8xQluiT4qnUwGiKJPdYdmTcoPF6x+BvkT/H7wYO1cZD0i2AH
Up52w1Z/idW34z6gXnL34YgubIPJrY1TWaggy0YYGYjKeaarElt6yO7K6w5EF7zxxBCu0cse+eSO
CjzAGif2MeemZiWcihCnuXq93Nb7WvNZCKfWowsZaLZHrUKmtzknnc52UnRvgHkqgaEwd2GXNN9G
MAAxRhEUGXfcVGLdi2wi4ryYtDrpX6Y0gzSYIbSLy+Uis3cB9aAPF4xzA/YFv2NAvf9i4nAj76Z/
U0tSnSKQL+SV2mDNiSfqCL+QTCXetfhefkpRkVTwuOwQQFW19uz75DiAF3NBqx8dLoWHGwOUSmL9
fD5adg6ckqWmCfHihDM29rrF3pwA7edpK6rFXBSXKWmxDxE6yS3O96wjz2nvw3LpNIXjeOdsD2Yp
HQRedlb6oNn05C4OupqRmc4v1ouwpBe97QrPni1QWIYsyxVDns+W8cA8NgZFMbtnXNnOLystzJFu
tBLwItF3vQawIXor33peu75GMsl4CxaBlHec/LL6Ej0BpO064SMJugVLOVBzfVSIb95Uojril7wO
S0h69ZDuYcKACcm8vbRdP1nti9VNmRczOpDed5UK4sVUBYK2nmGno5l++qe1Ekc1OCa7OPSwxchO
jwcVFJqtPJvS72koMAsH0iaVvMNu61W9KJ6hOGXKDXAR9Veh9sTUmjAeTXmOaHhsQyOwBFVF1rdd
C09YGkVy7KszY180pqHXyLBhwAsEKV0OIft99rc7zApr5S1Ja+9U8bFsBA3oiA67tChVhCwzDIi6
B7UaDiWneSNc6jc/stjjQbOqa5cIOUVjBk5koOAkw822W3q1QbHiu7gNtR7PsNh9C6sy3s1lDzDo
lllWL57U912aJ3WtXgkD/pEf9Oc87iqdwTRQOT01nKGb3YqUBkKqObS9LLOK+SgBlxoo+2P+x3/m
8FdSNBZmvFx6m3eLXubUechBrldrzNhBNbvYdYcHiQx4gVVZyfch80OerWJFwDJnJE1zAP/5PgFj
pTjWmBFCWfd3gxsUwc9PcUFNM63R70sAsuKpmkRKhnmaoWKJQbm7cXhWGuOGVQcuen31OpHFhRkH
74EzFhGg4ivieqygJvuEvPz4/h3CPrFnXMz1cDBv+ma8SxU4j/Jr8bYrwH8Y3oD96zTBFQN2lVtp
HaZ5ZDZWO1NlIDScZ3DhLwrLr871UOz+tleduWowUHu7onxuv8j+lsmbZ+M0Dms2uRlnBdn0yT36
bqUnDGoJ+UJF2/i0X10RIlr6wZl3bprMEOizek47ZKtGoZ1EztGN+MxUJ6GDz+YsxL/68mqsBNNJ
xjEaekZFIXQtDmSDFVw/oNNEFL/Y0kRPQGnhcfUPubOw0w0LDQ8jIuSvjHRoIFCRkofI2p2YmTEB
I7jTtNTWWGeV1avHAdJ2L/exAzSLRVGOQ/xZqtQw1Y+03uXbfnyq2yiY2aruZGvuSKdzoZ3lMEyH
Mbos9844Xbz8yFCrVNaC2pDt3kbVZxfnEil1HWYAkgeADRCTBCQflqODosjuPzngFake99x6u1im
UYhjg12c8eo+YPcjx0L5xmCpoSSshQQRKxhL681tMD7iA77Dmyo9ukJGDEj1h8awwMy0DyyqMyu0
ndsoyVlEfMfREoS3l+Im8OnSPtO814xRq0Vx9lF1np0NF0sz3uYVtZ6CLnfKcwck2PIhS5QTj7b3
GJlxQxrcztE57VIDUevnN9hgUVf/iVxYHrEy5r98EHJ9zNNJUuu4AgqZFi0hN7YJqL3lQZBS6h74
0xwdui4UaBOwoDL8J1Opq6BUZ9HKLG5SJS643hZZeruDH4ziMzCqZG3tlGYR7mgj0e7SP5Qnw4f7
tQo14/1gA6gbyqKDk+NRnJ1KWOthajuDgwwFBddOKY94v7NBWzljOaXfOy9D0VacTChn9R9K7JAF
Cpk3+woRg0WzKfeVw2wfOiwR70YGIXtRyrd3fYtxexthsWmD2LTBVQVAriuVzHtR0MR26SldPzzm
3FaPGgQlyDfoqjVdALBQu2TVcOzfockCo4hCGpLOH2C2IDaV0+uzlB9lp6FP0GOAz0L0f0N5fyWs
yY4DnTrvYz7HdbTgOk+U+oE2uG7EXxtz5dNiX3O3drySHD22UP6kspaD0+jL0tHlhRmtqh0nXZAS
j/aaMVau/cb2yghHH3VHS55UnS7a3EDivCjoHRHpaKubF6OfDMILs7kLXEVl463PI2idfXj2Dr7T
1nQhhYV1zoKS9OCl3/H7dFnQ68jNm1xYjhBBmtgVMKR6cblncy2JqCRK9L2KzHkjrEQ6BD3znZl5
im19DwFHcWDAi2zdrsb8SuLbSKEmstNRzADslWRp33ggpLp8qw9DmSJMidCPagZ/xud6Hm+tuhur
rASac1rdqBHmg+11pO5nuWkKLvLYROZLLEAuTZYV7bTrdSegb3WYeslqAqRasRLQKAXeeL6Dn9UF
J7+C2DbsaT8n0OVpB0D1wZF6k+GfClEr1V0Tz5k49+LN1D7UszGm6hDhOqaeldXh4n3lnWWNjP0S
/wVjl+LofvZ1r4YFXrEVvHTZaDs0o5HV8GtpbiAuV2K+alprPht7pQYDajtDe83KYGFCCAlp690E
yxGyoHRZWh6ybWC9FMkM0Qd2ahh1+uYdZrPxYsfkeSd5FUuq0fyFQkm7i91Y/1DP4htVbBWuT1ec
epzbvvI4CQk2eS+tZQgi0k1zvfxAKvHUadCf49/+BrUEQIISvensWPpMrbpJazaSuNrMnlVA/wNM
14mBmoo2W7BpSyEQKxBrszlGu9IrsGV6o9DZdd2i2LWKVEeXmIFHywTk6tF4xLIn+7PEDJF/h4KN
CzjC858QKsC1d1+rcp4nXpIiUC5rdgeYWGPxnSuN+eQZZkNkSyr4ZHG5R1UqHG5W+Gzj6YXVGYhP
WCIufv/JRFuNO6UFfCL4f7z77M55Q+IYYsGBLO+ZxVOfdn3Fu7r6yvnT66Ecz+FTDtiHFzA5avv6
8nw0w08BmJh15Va+t+VipwGL9A65xgk5r6ymuc+vQprfCRif9MUp8G65kcfIN5DGZFCmSwKGo+2G
51ojOXenhVC+taohHOurm3+tytiCeotMiHs0UNb/6TB+ktHQTFQxoz+IqB+z3pvHAd83BiqL+x+w
8taLgULHYvvhM8uYBca8mKUFVK1m54yCxP6YB/pRvgf6R2a2AX+z6CmYFZrRYP3l5wMdZgkK9/2Y
xyiYenoSCcLQ6YQaJNSvwWtSnjPx4RD2swZbl0L6Wtpc5eTw6AlRYKVDOo7RqvzIcPXNPRIlpdeD
ZnGtJlwbdYkzqWm+kslLTD1cJaZ3quMphCSwpxzpDh7P+ReNOYhhBtGYEJpt51ilzQ7UYpVAs1eu
92qdjFiLMx7BMnf2lkLE8HTCLE3T9Fa41YeoMGFWGva09TZAnpMeCEp6L7YOuQbQsE30FOMXrk20
eadYXWnPmV2ZYOcgFguPqd0IXF02ReFajw02JZWh7wbil6DD+/KcAUF2ukIbBMp1pbUaLAc7fzUI
R+WdukEZbIhsn+lI7V1+PNKFJaAkjiTmNBzMjCfvBnfn9BF6DJgsj/4MFx0kugTZSD6a7x+/Vhrh
2cxpIYZbTUYu2T7EywX26Jct4ksJ+OGUY/TzULo7gTttaYCsryjKrnibRY32XMepveHmVEsP6EAi
bwtsNm+MIW2H4kz5LQwqi525pxDquESpkx+s7A1bmuxpEU+DuN+7Q/D+JQ3ulH81o3t3pclSAK6h
0U9ledBv6mKmMmq0WMgDkiRqASfiERnqqBuKXHbvcnVw7Lv2LKp7kO/6or0TYwJ9A4jpp6AW3QDn
2Y+l3Sx7diANbkL2wZd7hzEaQPrLHbpph15zJJu/fXI/z7/VaUopqN2F/RIU9hYOldPAEA/tOfJ7
UcnV4wkdSg2XOfsIxrPOm0QpoBLuWtSt/7fGwInkzFuD7cV8DAf62eG3LD8kQcBJrY5+dPJZ72RH
cAgyWDIGRONRQ+eHEp1J+Q9ZHvdR4fgtMKT9/yuQSjrxjj8qB5cPsyu5RLHr0b/BS8itBDLNnCPJ
IUbEsMGObG8OSdTaN2bqZ/DsQfMNFMIIv73knPp8mrfg5g23L6WtXXd/sFK1cjGKQ/9c2FS+wq1Z
I7AMu0H31Hfi7sShYqIT76h4wKhMPwKzZ1iH/wEC26+2KlokQoTIqqmS6M3toYfNkfowDeV0+7ur
HK18qNMfs8ncPOSgcuLxExAeTWe0cQAVZGrkvSK6BHRdCsFOSFYHnM09CqhjyOLQY0LQsBkGQbPD
n4GI/XABcpcd1r7FQHc6TmsCGjtc2/Oc3SWaY/qfrXwGJhgPTT74AGoQliTA5PQD/o7kb8VuMhax
Y1tv7x3L1R8jg09SzttMBY8GXQtBOXY826w/jOfGQgGy1oZF9WtUGtNGX3owJisx0fJt/YwnyWVr
luLb7qC9dndCZefS2cUENcURVQuir5cVwd/G88xMtouTpGhzGMOA92v8XFJiuWcjRUMnAxJkCwy8
YOGtWNKuqOtxBHOal3TsFU6rQR8ZCSqyoYEFYpiqaDfRDu1e2mjM4VClyJitSE7eeCFa3OGtDTq+
nigndoL3zQDlDM86+zWSGkgYTKmdcSuYLwNQK/gJW5HCcuJ/aBgQU3n0qJ55tEl7RiwYEzJE85Ox
t75LbrAHLtQ9qX/gRksS/apdBQGwgJuiCb5+MRl7YK2QQ0w5l1bJVDkYYWlwnvb1dI9tj0HC2cik
cDZdIQOW54SrLmSGrMVGUFfbSRTbZUCCJJJxhkYouN1LwJ/yWaCQQcH+fbrpE3/TdmXcDkBRnQdq
y8sln9xkGn8bufHuqGN8AKEZSA7whFRuetF7993xMNsNqlpqnx6KRtccAUakUw7iLU44MNzkN4m+
UowQ8YkTCv7fMDWSHFgp99zy33uk/nlTvf+Sbg5HNLLfambW2jth47z6t6OhVBqyd2FNb1k+cJT4
gc99FViT6xvbg4M4/jpAaa0BgdVVecuQtsObJ75tc3dgcVg1P4+aN1boI5JiiVhTnO75Qutezzt8
V1GvMm+fAeYhyJtyksRaNKQCPsgBV35u7E9WhhjmVYp/hYsXqEh5EogxNIyt1zhKo/Y+Jfb8WFKT
SJrjELFGm0tDKy/2Oce5iujMB3BSFZV21uqxcemSzZn6HKYgoS84kzbvDxsuUavbvbDG0hyBrFNq
Ow5tEAzsOvZeIqMRaHG9fXmDAku7rsmsd8DtxId0gFZ1iKaADRIGQx2cI00b7H1YTrYd9XwxbC+c
SoOcpnuWRy1f5yv34GFj4mBKl1K42sjpD/p1zXjzVUL2VKV9S0LAhLh2rQoF0XxKOuKbUwX/meR4
updbbmzrw44WcgjHQbs3f++XllasruDnXeCexCGiGufEEngR3blwUL1WuCpVjGGbZdij/Ye56y/9
dxBj6awXwCrB+OQeJiPrXccxkNOix7jTqOO96ZAPGk6hFxNXqKlIMjIL8BOII8Tk5MGU5pxKZ8sD
p42L9wYYzWKi+h0q89Dy+0itN9Pl3XAi1kCo8T2zHJ4Sb8TlVXChRdRyBh/gWqhLMYWSIp3AV64D
HwRiYqa8Rl54t388HLWjNiRR57MYmrKMAJcyqo4JTo72FjyhhRdxoVSkoD6l+sc0PN/08Ufv8PoU
uAe2HwfkccnWmdofCLAYBJvBmJtkkPb/yTbpuX03NR5Ws+BRw0K0+CxJxrgVd3/8yoBZCo3rFefu
fgY0qFxEqZzxsrZo9N3Wl0xjrzfvilHcqNLLE22ukoZfHyRpELfATsmI4cZ+M9ts9/Wh8zZQc38Z
OXWY+qXZ9EeuP/mTX9tVha1XhjWdfssVAaH0pRv7P4299YN5EhvJ3theDIvw+w34aay5n6IuYjcT
51/ygNAWIyTu/8wwSQxMjK2fiE5HVj782dVrqMK1sd68Z0gUnV3f/VGHirNwJ/yRphBwAgFSSfbp
iN9sahTy1Vq/kzxcCDoFyuiT11SFkr2vPtm4aTVMmHmS/DKgYqE/1boTShZoyMGrSrQChVvaderM
CdWxl741DqruOwXJVluo2+jhtBw2GlBRo1EufxA4KwqPcn0PtFucKMowWKGolHaabEAGXDab5xPs
DBl+l8SyIiySI6+6+rIaCpRKjtHo8g6/WjXyF6US6yHlhSxy8nRGTNUxBAEt60VpjVJrhPcq+Pqi
W2FsQxwxZjeuMetKZlPCRKFQ5y2EU4Oktk+QFB54QZZY2lerkTX9lxg6pUYs+OyJNB5mMp6yaPnF
OsDQQzySpPqlODTGzutuItjrZor+QvMDKzqkdD/tamZUJRG/hM/ynKTgeGFC/Nt0NjQwPSL4eVZU
lvJ7U+jzX6oQQwGLypEiHRrTUxiNJDcIg/ebXrS9bhpDdoZzQFMmVay2iODoSg2xlb8pFdFhLJ18
Bncjw0KFpoJo+5AfzJZhQRurAkohAlxiZp94254OPLDB81P1l8TGbgjcxwD/TKRfFGsxrQERO7lO
9ojZrbU2QbevXHk7HefUo4m8OfZlDsDWUTxQL50XdcK3h/xuVjuBqPTBgE1J9x440h85tJKRcx2f
Bp2KZcf6BchNzuls1w83ib4N3cs0h/i5B9dRC4gCeomut8p3peJgsvC9KeIp2lagjrhVJPMKWnxL
Iq/mDE7Vd5hVEX0b/eCzNrBO+y5FNaZwBo42pteh8mnerlyhniy2AmLt/TjV+E8rzBxbVfYO0ApY
Zg6J0zbXv0JRWQ0XJtDESQOystSRRPrKjsr8fB4+xpqKjQLX7ICBY+Cajepi0eVzhiVBqrx9kMjI
TwKmAVFDkGFSobO0lfZhEuVi5x3w2gEzZWnlh1HAgI++ZoQNs8TWHhlNHJiMx7Yg4VsbFTtWoc90
kuXFtGPLZ0l45IMjyZrSxAEAsNbRFs9sVjB8ZOeU0SxmTfJ3FnZBMysB31QLE6yDU4QM7k9CNIZ8
qZRkEoD85PZ3bMCdY9PudI13LFkkX/3vfDtiaqIeH6OC7LLhYJ9tu82gGSCZPseEPtyO2VJfeDda
dhrRM6vJyhi2Ji6aKqZIbh1GFSupdeouwXjgqpHkPQInQ91L8kLO2S8E4rGyWnOTPYtwraPt10zP
CM6kquLIMyXmDFKeFb3XuTWQ1nNp6SvJd+pt/CGTx27TLHEWBS/Q/wJR/gUCYBpoBFx3MDSHtZYw
jLLUZegGfan4LJh1p6n9W0P1N/ARvGsyqfEBkrEbIP34ZFBJTA+OmluxipA9jaUAwJll+Uegnav6
44pTntSvQKvNaL7KTgCJEu50nn6GRKsCA1Rqdg0Mml7CGv1ygbx120AykPXTvMQ/t0ujfv0PgN2q
j/BYt+5Nl2Bp9VYhe2vjMFxrhAd1QecTrXX90xif0KOFNHBGeh6ZhvUEH0+hgZ5+4jmkR05hDoeN
srptArNnaXBGyv8csbkBVqTJIzIe953G2wdaWOm6ptMxetCj0pxrtWaCmp1BXXJYYgXsqVLIkpwb
uOMZp/LsGouyJrAElZefBMnHGwWXKa0fm+dH/7IOmoXDXSRjEER62FhqEjiXrrQOaRe60Cy9zFR8
JuYKAbMytK/0jquQCVx5CBYWiqHcx1mfIsygvgXSXADbzGVu11ZwG+hIC8M+UyB9967Zmo74KYHl
tFqwWVSx8UYUnGkqTw8ipB+jg7w+VI3n4/Xk8IbBkt0SUm5o+v65sBYHPKCAtcmhcnLNjmvs9IJc
0DTwlNNcZMnuFzZwdjFf0yEnOyjtPOJvna1ERkRhoUIcYHZDP7+t64LEnCx8E0zfLIJyub2ZTApd
u2+hfnagULzABsanH9pCAqOATWnQmAigvvnu0ddq5ubScQ7vAWmF9sIsOnlI0ev/rm2VscAezHrZ
t1nEsf2sp0kuugm8bpp0u1CGVgUtpCQdfPdnGJM4xC05/kIhMo2xI3F52wbv70gVbpi5lYKWzlmY
hD1kdmPyWQTj24Xc5BvYUcES/FpXaFNq0LfLpBXPzDYI21b7teDxL6In4FCiNXKwlsTpA04qSNdz
jROp66IeJRBrIMnJbnSCfF2YY1vyYvZIrRb/qc04tGo8MNFSYO+vf95+4fSY285qbgZ3hxNy1b3l
72vOocNtoOL+Hoqe1bcvUlwb2x4nEil1sgjwkjMqqEbYg4KXypGg3UZWU2Ub+RMNbNaziAQ13m/n
Q4+Gw/fh+cK5miGTigonFji/fAK1BrBqWdQz+VtI59D7+V3biS5t+dWGGn3F7dRrAtPIJQtmySB1
PRHfbU0sMznc2hVliuPfgepc251etT+Tr6zyU672CNFlxDowV32rG3QESMDTa8hwUkbIuO7jh81G
Kz+3I2C4eitGm98h75e9TunIWNNAz4QxipqiI7VOIhZ/VgNkXlmOTenWJ39fvK+awzvm77L1Ncxk
5bkxPKXahOwSafMNqD7OO4hbkKBMSEPwUXaiFMEiZthQS7F52yqTUpQYq4hYtCTbRpTltFgCHb2f
A/fW2ycL5hPx9amcBP++Ezl1417KoBBjUAqzfkWhIl0G0ZIN20QEYeIc17mH0OQALEBdo+iMQR5+
iEUauPKwphhkU1cOwZOOB37ilPjuwb3oJkJDxXM8rpsSp6/7C8J/eJhhRuNLdgs4JaqoBYqbd/Ov
9eTLQw8mEnmfX+ggV87efgUWIDrXdnHf+H+PRjee351fI4CazChfioWmOROnSTDXb04Wk8KjLTpy
54tkbz8rf11J5+pXGVgHF2hFwyyNpQwEKM+E/xARbS4ks87p2nDYjs1evTIqLwrv1YFcqGGYoSnf
cTbNPAgL99/CND6buvAYmKL/OlR/60SUFIly/+TRBAf78jctb9BSHgfvs4LyQHsL7zF67xKFl69z
KjIhZkc0mTGhz7KmhGsvkYGyP0GKJ3LhUchTrzS0dJJUWTJxG3tYuLCZ34gA9VjUG5PVPPw2fZuv
qzLjxyaAMVVQTGfzXKna55O5W4Zw70WsQ55iChjCR07IlX5R7k10i1KLzl3rYKLeQwTX3rJCl7eN
ABoFOVhaGvs109XF2UQaCQZkZR0qmXYwYQQLRftpxCRNssmWmxhpoO5f71DIIi/mgM0FKvnB6C//
CvhDn1HFXaNzQbJfL3T9GrptaiAHAfuaHrgXSiKB2OVtfl3No+NwYjWtODdIiyoPLjn+wEPEy8hq
43ftZw9fXgzBPIf2vn/KDEd7owb0McPuMubh4lZTCfLHclSbK5/jG89Dsvxja7tUqMStw51IM6QA
Los3WtDZ7kJg9GdsHoxrsW8sBJjIwznMfRvgYGdi0usASvtVY8lnX0QSpZFQyXc37xeqLusC6H6D
tz1venwhkYrzbLJpPPofqOz45jQtkvQnZGXOQ0I6UWExwcA3lZ5fd5CqLQWTwOlgobcwBgeNCQdU
iP144/LRqe/hYkQkfyd2tzpLSXOQMCtWg69pe49VCRXFNZPnyK9r2q73wXSyWBCJyFXdhV9L4BSN
MGFZMMghzneXHoPhUKFTw12OGDNjB4kaiD4Rt9M8uOedQ99KaYXcv+tAis4hfxhpFlAiBUFdBV4m
YpbqRTiMxCLXfhJ9SMEMzFUzPKErFICqxADzEpekaMmk5b7WYipV3Gu+86mk2It/Vj7QN0tgZcAg
4l+6FvwoxFvuwwMpPbe7KEIi5qiqoTTLwSraBbSs3Oau+BOVxcFoTcJaRLSp+5DpfAbsXAeHxPO9
lTSbpDKQtAxrfsMijocOQth3bShdV1mLRVuFVwkuhHoKTn64vlLVat60ys3ngVAOPkVh+UVJEjHN
bAtfeS1NDwOrLV46GNx9PUy/nIpj+JFpb5VSz6ugOy22N+4gFjU1jivoBQovqUS7WCOrL0So8Xr6
mu/ZrIOjg+mJ8XUd0+qQCRrICc2GDdR6S16Su9yb1JTd4VgZp69zViGZkomDCYHTh6BMMdoSQwmy
/jNatukp9B19WleKj4WqKCjW1nHkxYKYH5x9ifazXQ6zWcsB2odJDx61RAwMpLbzJLfib/dKXp2f
ASSnHM1KRHjBzelbmx0NO04ePENwi90EYAm/VHCC1w8sCPjGK4QHW3+csS75TTBUFd28KDq+DylM
6cjBQgCvBXQMrbfV6Mw3K3UjKVPQIGn54EIx6WGU9zmcwpaS+tl2OscUt6l1J/LWAq/2QUqOZlpT
SXNDoLJ1oN1fhHqCLgkROJob+zGSmV8eFryCwOWkBpC40ESRgoi83AH3W+VJa1CeTsOUMc84S7gr
j/H0ynT96Yjk5XBEn9IfE6ze6clPtLB2z+2o7ndudoL7TQuriiYASZQC8X6OzKBT3TGUlQLZHjMk
J+V40z6vCU4jNWS644PC5aF4ze6tUq0t71WqikphpY9KpMZxDxod+lh2bCUFzVBx8IE+bXx5W/D6
5z+15DfF2rLYfb5f1+LjC17lO3DU2AaIfAIQvO5TpRUF/FTjhPqgrkz2qmqs8qhnKjSRZMNse8//
l1vjB5MDmUayKP2xvJ1p9Nz8OkJ6YfU5DsfTzO3YE9vY2Ylb++c+yQu9+1R0LQUlnn+Vy4elx87k
s5q4obREKOWv3A1i8rjY/oeET1zin7FBou7+nl22gOkJ9mMNHPt6PswR7gKwiHgFRcu35dVFF+O+
t1zBjOXWESrEehaSudcoR8CNg/GNwGP/M3tDqFJPgrfXopPblbiym3+a49DJRGRXCDIa19JQdAKW
V6L0EcQy79zXuhAcB+XG745lgB6Gvkp9pN0xTLYM+ENPnAhOPsyOdSx2VpYWxfktK2jc48CfUfSq
0p3rVoXENSD0gCYfPSwVdcEYCH+cqOs/iNkoyLxcm9GK8ovN1IramxdvVnTs2xf0upvnjd3aJqzb
hYwt6+N7rrmI+EKE2lmdzZty6n3bFixgxD/lfebFrWzkjHOjg3ScEnet5ERl91KaPAMWBe3HESRh
eLmJ1dErXcr2sRe4qEPd0o2hP8K7vkEgQfNb3ByhD1joV/O7Xh9lmugZbqFjnloqRohNj9iiWem8
+YuBhoNiKFUn+ORQB70xt3nPxlzXFbGeZYoTvc/zt3QtBMSFdFO6uHqy9r2d4bxIn/JXXdVRCVd2
IEiE0MkJ/9Mxm6PqN+T9UykAVNCR0QrH1IEicOEY7I0fAi0XkTzSEwdV/WCYWVC4wgfaO3PPClvX
Rh4WAUsB76dip1mZKlqII3xv7bvM8ReBb8n/NUo/OLMpRrGaycveC4gScSaiWYi11L9Yr3UztW+H
yZDDRJb8NIbj2Kjsf7q2XR+jHagWlhsG1pJZiEUpcZ4f+Bkeet1rGXOsE+c3BuHBDFaoIUOFKLWE
Iw5DSS4rPmaETeOAUEd509vvz+Mnj+22xmN/7CURH5S1pYu8CwihD2fL/rYTf3R9mTf6sBI55nhw
MuDqyC1FJGDdNXXCgd66bxVZYReboCOUEc+3Ut85Jot7ZBX223MqjHdyFvZj5QszJWnEd0HFdYap
VL9r6xoqY82Yu7b9udCQsh9ApbC+midokKjNIGqyPm/q9kJNtCnm+owzuP0wJ9y7FMz7eSk05Rkw
/5GpLWlyUVdL5fE5Rwb3rqQKrE067ih3yrrV1umiv2ZK12yMC3rEJ414h99Xc9LanzuetkxpEW94
3MzDSUzwbNDn3rHBgjxy+Eu/Pv/hMFrlr8b537U/uP+2Z1AwAVcjfudA9iwgB801cK6kNMaSC1pb
CTueodGS6fh4W9mQ5IF/RuLBlZ+4bKfX0gOyiYDt+rO/L0H2Org21D8CDeh+i5vjXBoRMR6GjzGR
2g6V4EwQZoW++Oi5tkFCx75D96bxVsamCg/omFuXH1oSl95mB8U2GaKWBUPNCqjAUfXJ0GmOUMKS
C9Z1kg6xP+Yew6jIf9p0YvMeuMYKnB+goeoHkPeSsxUXvMWyR/7di2Ki54Anut/LFKksI73LY6BC
dJ1OkAQeJWJu8ExdmgkUllG/qRWmKGuiIYAVFHBnExKWG3xmUcILDtQcj1zZNI2tZhdnpFtnnmFr
dhyBBYZzwRjVs08ylNllHPqp1dwhWXRGYf4gLfmqgrC105jDF+z0klTAtAuA+R8F0pB+Q4vmapQq
CpBZ8y9u8ytoOcj7uVYzdnWOaOp3izB5K6p89Gp3aXOcfJ15sza/NIbUWJjT/5zXzJm2/g3QKTSV
tHk83oBS5P0hwErJpx0RI2US8CNZTBZ/El/kTbeGXNvb6IT7/c3AQxvk00Fd65MZ88BOleIIR+9i
L0UBLalxvAsuFozZ9Ef9kz4vHHGBVOLmHRaEaw92mMtdOI1RCoo44Cafs/1ISHXgHzAWDth7TjvU
J21S3qJkfHOPPUDzPlzHAEfY0HMkehgYWoQR+2gYJpvxnKIJ1aGS1ovmhJAEqRd3eMd7v/6rH+Vb
wd8rkTCubklClmJCOhhNhIqpSxxW6q287mYQimohLcbH23I0I/FpTgvyyw9sm4RGqlM7hB1t+Ly3
G0lthTVvzYos6++1pc/UR+TujjeT3A8wx4WEs/N3QQP5+WtXi2QuYLf0ByOC2Ca6G8sgmgR6PFFJ
Kxy26KmpYjkbs66CG8c+3np5ZGHUefZg+vMMAhfOjMpyp0IEOGNt1hZAc0NP8MPvrK3EDKw1GHQ7
NU0fOhf4kTiBgnSo3K2IzX8cKb1sMjf+IuUzJDn81GwpYqAh/bGW2i8VquTmW64Iqjr6aoEaO2mh
6zuY8RXr6KiD9Cy8DTXbF+DWWNgzZ2A4wktUY9r7wIzfscUeA/iY6bkuZ2OETUCeLao2ZWokSYth
EGNM7EJu+T8BB5JAKnBEuPaPh2rkAvgo4/DQ6URbYLb9IINPIdj3w+oxRe/GVVoDcE98Bbcsi1jC
jQsbsN11JfFzar8QsfIklnsNS2QFQRgawDBMGu6NyNhQZSAek5+eDEuc/2anUfAvNwu/firWsqd3
nwxbmF+jKyKw5iz5QrL196LdO9wQMqdBQZGEU9eAUAL3Y3vTsU+uQRVpFMyALPWi6hDW/4O+3wfc
ofZxtC/tBjA+GmNhO8eQzv0PvGKIdUn3UslQytC6zd4gg0etJaaBJIY0SLVvKWSeaEiIXs7Ez2EH
iO4Qc4LDpzEktfZLhevHEoAiewHdebkN9Q1jQjhVVm5P2CeUYdEUbYsdCfDvI55fZIbdLaktB70u
5iWRQkJvsMphnijpE8dZedCOCyo1OI63UudeW43Rwyg5FtcrUXsYzjzoyqdUkesV1pCfsHE3j95b
PvXbc+9rvvcUmv3cLXZCJi4tQAjJdCwIEZeOXrQMp5O1og+K/QY9PwZGSCcAIXl7ypFxx+DFQGKH
ECRqhvaCKcZ7t8jyWAhb1wFHev0stVky/jDMLYk4c/axHvcxL3Iv3XgfzmXLD0H6QlfCZAVivA5s
RV+nBM+UYkb4bxSw96BF4i3kp2Ql56tOQyKpZWPiQmhOptUI+zzVEd+WSiyncQF8cAZwkzHX7tgs
CVX0v6qizRaqR3I3pe2UY+My/e8VdQoD3q3hRCZlDb60nRaGa3VPc3T5KVDsr2/wzIMWhYA/jVUW
yfeNZtHQCCbxykz38QOvVeDf0e4jGFI7+6mnHMB9ILYDWTpdFtuyouwdH+7WHv+3D32Hm+rGNX5h
Bg5yKHtKBWTMryneA2dOqRDPMiEJxxyFECthEVAeEJOA3QfoGybN+NGSOCSS419DWwPnX6VfXNdC
ol+/fiLuRcmQW9utKjKBz/u94+bCENoa+X8Y5uzJzaVakYMykER5R0HyA3t3j3uhdlJdrUEyOS8e
/yuJk2E5d2475PO7tXi/KdSsRSGDkarewVJEBnbumAcaiGM+K9GJVIfaVtVT2+9c6Zd8MFI3pqd7
Io8Kun8vqfBPt5aA95xbKkgTAsc2HbrM8706sBqAJHaHvvLYZbkJ9bxrUWh453BB08syIE7/PDVX
yvsqBzAo1SyjFS3dC98NiXDko1qmFoTJtK6U+pyA7SVhMMC6//PtFjEfpkTgY8nR2a26bI5Yj4Gb
4BBiDkJbctRgKYimRf4XvBf6B07MrG5HgAzu6Z1PA6hK3wplLUIr0LR8CdQretwLkOABcjY4hU0x
2W2kB1gFVv7XQx9O6DfdZCY2str/RI04My/ZPIUZ2ouAIbvsiXauJc/rVmIKhQdJ5HjRfR/Ctl/Y
xme/C5WN0KwqQCcEbRpCcjKkoYVE0bdNTojwGjO/5V0dndPbKBjehZ7K2nCbv0dfd7s5rZtPqnb/
rlxopyJSuCB64OlhorzzzZNjeVk1gvN2o5cxvzVI4cpMP8Uh5I3Ztg0W3nCAUUNacRwpKJj7qP42
Xs+p+2oPd5/RftJgwEziVyMeI611qyERYMyW/w1ttxwHGjPZqT/W3ljBDhBrEZ/ZoQdFzoVi1E/r
V7lC4dvhtNG5k2Y42qyezyE//0CmucM8PNNuQq+W7StmY/2Vww0BHB+LoMvi5jwnpuFpIvSzZjPL
47NTJKBSKSWqNsdZYr7+UJ+phTQ9CjMWodVDvubD/VjXrNMlJJht1Ukt5Og2oUPSbnqFmRIQMSGq
af4UhHIYpfwo/7vWridDANdtoYll9Qnk3DX/nYHaAp9BluoxMoIQh6pCmvnUnz/3MSOOj3xc4Qbl
HnjTBNtG3ZIWk1vtoFOiB3iuBkUylll4/f3EgQkRXXrPEQzoR6keLKJo5fBl/GtZqA7ys8X0ZDUi
eN3GROe14K0kQqqPhn7IwP2xn9o6eMqStgGxrtJ2xR+cFPPP5aaxThpFeg1DwG+70VblpVlhiFEY
LoRBAXy8vPabdB+n5CwTF686fEshYxhF9wGed6J2jv6XI7YhihLWSfTOuFgbf0/T0rfR0GSZoEd5
p6EWmwxdHkAJ2taV7myNVo5f3hG/+P2xbV1fE3yws9e5hwEanViKzbHyS6OyO+3/X3Y84zBXNAmr
TfvKqMG4hVKVWqcB+lNrbCYwdfnERSYZZgZsNznRngknT5UUzFXtNo0SycDhnWN/cGCDTyKrciBu
Q4rzahD90gV2zjZIOPJ3UPWMGQW6/qFgaeM9fZAlewPFdL7fscBe66ruc73TdnGDgseGO01qq7eM
Bwvzg+b8t7pm3RGoBWDOH8baB7jOyg7qm9T7Gej1jT4GXoJNl+0mIbGw3JFAK8ozqT/p7c+Wagjl
8hsqVG2l5dsbxvm/2WxjcgYox89glzj1GRvwoT/ZC24c4GuPoJTy6Zb5jWHNB1qxpbG60NK7R/bN
W7JQM7whnax5xOsD+xKMTlD/oJgXz0OVOfERDcb5Kr0yH9ZnICYURS2jMXAaKknoOjG4Fa30PWbT
eKQsfm62giLGrwmXz087I0+Yi+lcJ23sdtaTtpxAUXPy/l9M/AsS9bDUYLn0pjMmGEG8zAl9md/I
1zQCfLCxKYr/piFDd7UxeD/9U08h03kxR5+6TUeBAhk4wlBWdKkCwbxOpn905rOon+CnvW7RafE4
FR+MCWzlgCAlXzNjKFhyO6vUS6EkPuB1y7gl534qWGTyeWL/hSMi1nedBb9nw4cBObR3/6zfroNo
JDpHWFm/5Z53wAf7yKNjltLNtGsPCY68tauisTSngq0aXtX+F7vCPpQt2yITrcw5cndbaawe9XnA
zfmkkpEGxyU3i94hyaIXXWRtVVQpfnZQVnSIoEURzM7gKWUUignlimhcSVg3BgY4T+SpvF48THML
6zQ+KCmOCgC8sG/KOuE9sBEB/YPWAo4KxqscXOTOI/ttHwu4lG4SaKUhtlV9P7jr9iivXammy76K
DCheRtDVvYjdg+BsRl6dWmkoEL2/0m/GTeMYiCc9+hGRMJritblov+qiPCMh6ecb53FLtICttAM4
9OKffxtUjkp/P/U40HDVC1XUNfUNv3uvMFt7KLCCdUYLbQkiCihz/JC6NNUZXjVeuTjvC7fD/JIj
Is/F3PEMvgDSYBYN2npHkNLA+PsbgAXWeDLAJMO3eZ99eA4ZiDtGQR2R2oCknuMTGBQA+NzOmmgE
aaQMhY1vwyr7TxgC0E+zEhRZbxJisx9JWUelOOxQ7WxoQjdSig4KJzsj73/qU3QhE81sYo54ly9Y
hX/AiUf3jpDcjMenLOW1J+5PiOEL8GKy7B2Q3C2wbmGs+gJyJBhGv3RYyiStl7+wwQFGy7A71dmj
mdKSN5mmBCQUfMi5VjKySVp4vQPutER5yFM2/Rmq3rqeBBzUiPdfY5WUlFe9n6GojUqTbENAT5VX
u7XJ3XXZW9QAZhvbLwyD7nOqR7xKgOISsAeqofDHyBEfbDYe2BeHqCGrKYCyplaF5akM8M8hI+ah
Mn/8bdn7Jybr5p5CgVF/DkcYA+xvc6slbY2G76IFysxTVJYx2Oo99BLyReX/25oZIfXo3GjEa9Y0
nL1ycprPtDapM/JNspNkX+NxBDfUEcFhr4xZPsIPbfZubrDMnzNAJhatvZ8dPmVLuFvnoSHzsL0F
cgWInEEfh9KYTdSzrg6f6rltoe2ydlxacYzXVtNt1morMwp0/aFcx46L3+gkxy19HWeoftEzCNhZ
aiLimZuLGV4MHwi5ndM4LeYKiuB/wh7TVrXTkUn4/8PqBPIxS7OgIeVM/RVFpSCxiKvl06lcj8u9
VLmqjvn0cpsUVdvUggXCTtHJDMGKuHUibC1HNPt+OO7yIfdaQkP26o2x0r2ezFQ9+mvMzxE15Rip
IJYzzAQMgoIO5ahRSGsWArfoq5KA3UmF4KUM/qiFHr6zaRa9F85JyhE1GgyVTGpScILFuO1r2EOz
IqqKBhVONy/LbRS1Pko4FS+1tJNagNxlbLdcdmQaE4m/Y92HXWzy39j4sITIQ7N5Sjnfgk3gbwm2
XhGCtmu+H2Xo4DC495jTLOqydaLoPDeP4C0L8Xq4qxAQuJH6dmUGJfB6udoRy29YZdhEKFz/+faH
DLuXd4IzdMIsCOvFmjReiCKSyaJp1pgrrkTmmni3tzsdzo2O3k3Tvidx5WeiG1eyO2OwBic6XNdg
dapeOCbkRvWqGvNBGehYdkuzv+KgpMok/S82SbJaryxnhQJwmWi/j23F3r3FJdsCXRP8YvUuqEUU
kxGaSzhDf6u/U+rIpWD7SyFck5wrQLQ7UJZMmMBXM+v5iuw6VoNYkdJaR/uYUrPqLJxZRfZP/IeK
c64y+bMxzZYuQt/5nOWqXjIgjlI5K+tKgo2/sn9H44cefyFYmhWkdmXNiWgKhC/dwMGjVPRFK2BT
l7GmYTd413TDs3V9szy0xjufnQVjJCehegtKpTY+Vm/LhZeSaVqSfnycwAQiQcCQp+lh+FuDxwIw
d0/gvodD4h6Tc9aZw2T9XUK0+taaFY+W0TseyusuHOwu704PaxZJ/vNKHKldMQCC1jXhmLeMythq
dNsYd/W7pgxXtlZpge9iy5JQbgwh9D6IDdHQmpazC/mDBBzQ0rIhSseL73ZklQ7YvP+7WjBOCJLx
Se+6o4ByuorfhrW1UtAkNbSJNiq4ZlGvN0Q4ktCWgWbOwswFSSdMHp7CxFSPMDlx2iknIHNtMzhP
04d2v5oZfAsGX/lvYptmBsNigcAh/pDnHFs0MRpdkNjeZGQ6AHlGzrhBOIRrKGR5NRIXhXKz0jiW
+jNm4LPm2KRDUT0RwcO9NquUlJICfcSt5Nz1tXFNiH6+AgpPXZx1ITANVvUrzaQ6MWGZ/we+hhB9
M7oH8p7kSaQRob//yQ3P6CoOB4SwJJxS76YKtIfvg052EN2gDmIvhBevzPtXqhbiP0M0i81gBvQs
9BYkEPa3klpzTNoSSBYK55XCei0YKoubisyxsrHkDYRdApZjRUs9+owI2qM3gBuUn1ssMEa0Tmti
Ji0CRt/4LRKYjEEzXoHJ7fq+kwpC2B1ITOJ/7hjbxYnd0sRUaOCmScnSguzDQsZviEjHueuVl1Yn
mNeci7vpw/N0OE6Lw7sj09T57ctHClUZO7qLHXnhM3qkJFliMu81nNNpUHkj0pD+gRKep9hFrmCL
rtZk5ptbrsUaSVObsC6oreowGSFdzAQUxbetcvJtqTD2akW2z63cHZwv6pul8yPZQS5m4Q5tTfZh
6deavUIWc57Sjb+SHCn9hgbLCdql6yxBxImijllQqsjm5uEsVqJX9Otf0ZvMMOHKk+fEFKRP7gmG
1NgNHmTw3BrgqSaI91TGuhkeS/Ixea460fOlV/2xpb7/22vxEVl8UiVhMV5tNaOI+tcz8khLykBR
nLHOTdzflmrDalCcF2eD9bzcwNwZqOebYy4ppCTCsz5oB7A4HJWGiyFx/MaEciFX0EiI3d34Jocl
ISYIjZoRQA5a/0L1xsTFLPvtgtefhStuCDkISknQ/EoXOMYihu4Wf/CIKOBwwr7/kVlPROrdA1Yo
SGmap/ebUPgV446PNHpwYuHzcINZvCzGklVDyFuJFkrJCsfxeEUg1RG9pOiEOlmNh18X2HZygV6O
4k/JmpjLcu2wcTCHJ6OJMYbZ0pnto4xWTcXgiabTHgTgzF1mXUE+a6z4JoRk1UZA8HXvYBYXu+lm
JWy8qATqMCWsZjErldIHBcahsS2uYaAGTrLD+yvwFqwQpDRR+zYzbPN/0A5UeusLJ+CviK5gMCbO
I6uPCFv4JG8gnBpdhNN7ij9671mnbyf9/8JTUK/p5fV6YfsPy5ciPtR1RmVD6zy3Fpdpa+wP0pIH
d7o4jL/Qkir227G1T49AE+CAeGrBe4dulVqIPeba5FzW0aGJB5DGWUn0kMELW6S+dmEbF0N40CoE
QSO5+g3NY+UBfeAXqviozxpowkhizYWdF1aj6Ar8TDuK2G2GGKxnpRtl9AM+adBWiNigLjn7HFSE
QQ6RQqYh8QtPXZLgnKgWNahWntUazrXN1zZeg2KUm4PVeQBc3/b1qAudPrYCtIedxH39qT8l5nTs
7oXZ26Xfjx+D+iQfjq8DyEYUVD6qN2jsz+XVNtEYrpOcz/xGgBeQpfkKQxKZBGEd2Z08CvgvURan
z2bySuYiMahHNKCbBKicwuBJ0Hd6IvNQ1gl4QobMzIuJL4SeSDsHtViuvBzY+3TaRwQ5Qe2ado8g
HKjbEWHhMcCXfhJmgHmsq8VniQ8EyjdxBD0TSZSWTzFA3O/C8G9YiY8AaVuttjsZheih9jTZXenL
SfV1IP5pdqwzvrUs3paGFc3mxmzQq1D6qlbL+vd+YFS1WGdnRvs58vUDRriBTRvXKO3kxZm4U6Tj
je92MGfHN5mxtwY3oLAOWVt+NomimyayRwXKlfDnT3MsdP+3i6cYOO5aw9yG6W4fEkUzq4Xdkgdj
3SuSUBJYngchHziNBB+2PUNy7zjWWaC2W7daqon1J9CzJBFFbYbZbvfRgMeLIv8A4/47oCjyj095
PzyUTBlZr5mvbyMfZ19arvcZS5SiTYA/O6G+hovC62QlZN5ij7//C/36FgsBIcuvu052nPZ31YC+
v7ds/2/fwQq36gjGuONOT/g+7DNvw0qg+1S8Kv9m2yJdSR2ngGf4sBXByZkx5VWVFPUzv/WIvEhm
OY0MR62ch4xXDXd2IBFQq4Eg9ged9M02MP0vBkXhTuxZvlJfz17e7ESpK3KxRSKO9Ai9NPKj5b6B
QVXvQr1/GxKTRSz4LZU8K6UTjs75zix6CmvzUgqlx8dv+jwxWezxgtogGFsabe0jDILINTCNjoTu
/2CfLLof52BNuprBFABJaidW6CUhihO/AxRmZ7YR7jD2EIxVa/Ln3lKnWcngva7zm4wkOHfykfEa
7LaaO73YDPL982MICj6Utnc+ECjtnb2a0S8/JW1zNMg68kexRZBFapVn3pEp70c1oL8FC6bwqWGm
a4va/nTaqvF1tOC9YqkQYIAJl94sM1mAJ71p9PH5KNxSzR+NBhEvlpPDcJwT1Jp+0R9jAXcPjU/z
C2ARvT839XZuqzRXUAmhaBahBQiQNax16Mvb7W2Qih8WkNsx7q7gAQbJIfyz7Fw7+PQ866y6V5T7
4QYpWV6DSbUMiGwS1yVTvtUM1BT8rymj6j576II15H3u5Virl6x4UJs8r9EY0Ok6xg53w6Ll1c5b
Rxon6nVp+/nlqWB2iDQR7gmP4UrZkVcLI6uhg/Mgew5EsRfLI4p37/5mQfHg/6uTpSKrABAT62W7
TwOhsVh+3+dEZus/fCDwh0kFj/oECs7SgnbtZUAMeK1wXXXHraig17syyr2hnkmDP6XIMharWM+i
4pH3XNB5yBlp3cDRumVpljHsssPDV4Pc32zJP3j9FZ2mpEVyD6JZB9bTOoXB5Q3MxbZYKeVMETQY
K7L+MOgMdRKN1nDXwgVsBWR+yF7jslf1pp4cSGm7P+YUdO4Q0QLCMLYSxsJBJQFSB4ONs5v/wyjP
U9J7mug1QoT9FQ+NNlUzen9JXFn5CaFElLzHovE4whcQ+ELvhNyntERSq8MOdB5PyrLzAjZA7qLX
KXSzAZmvpmRtMMWFKyvHk2nSWFf/96xdPj+h19peZ+IPftjob7O5kRoQH/xFtNdeFT/x64XuYUkL
nJCxBpMigO8UJ4RtcyYz+lRWfMkRlzn16CrZ2iaLOrtImSL6mDDMkJJlnp0lg0LpvyDDxtzYVo3K
wB7a06kKXGzRpPeKQNOeNZFnMGf1NeI37PZhSplg+fHw7zKaYIEvZjeZ48ZAOAOz9Sz9mbv34spk
MCUycpAyNWqaRsATo3eXuRLQRUsZ1FV4rUH5eCnj4BOTHs8Dw+hosiAjdyKi6i9WYBLcVhNMdWhY
jj5Y3Er/OQZt7lPnXxMEUWkySxsMQlvDUh+GSPNNOJ71EdS5PICDqg8XkOYn8S78ltMY7IUkkVG2
hjSv8ZJUdPyTTu3rSh6OkB+SX1nA36G9njLurGZ0JZtFhC2oIYRkvRnQlIzgOfjpYxuTDCm0i4O5
d3KzYAvrj6amxljNPcbFVSL1k7zxENC8pTOSlm0eUtn6L3rXPpu9y0KGYZlM6HUC3vCfXL2ED/IY
tgNwlQC594LO0/IwrnQV4dTjy2i1VuWhWvYUwtoJczIxFPc4jNtixxQa6j711NWdfrBJ5RSLENFY
nOxd0MjSglDb3nyj0gHwlxUFQWWohHaRrGd68kwQ3eU836fuq4AiGq1Ly3ul4r1b5VzqEdzrmqca
J5PyPyKMcygtTZByw9NeBYcRrJP9kJjWbOybQFoZ0oz6D5hlAoaiPXFPPv4w1clggY7SOey4/FXF
l6sJDrjWNGXgxV3PTM9OMX0g60E9Ftdx86GY5O+Y1ZZeWt82sUbnEe2n4i8PapAUA7ALO3atSNpE
5v8+BPyzgYTShYZiUQMDI5jQ0flOREkKVxkfiK3rWs34LZoxqEFsozLuvd0CHABnl4Y9SYEv/SWA
wrt0gY+SPpbRdC3g9t6vbj2dAHB+LM5BhUMKsEHOVxURuxSknSYY9jy+k/vvTlEkktTowcRuML48
5Afzi/uYdyXiqKu4iiPlAmpTbJNSHcG9PgvMQ8abv/FGXpwJ3f5yybUeVNOp2CwhHp2J1NjfFEo7
hdv6Q0TdITMmskqxFLfwsBYegswtMrFJILGYyEBwHLHOE5p/DMAF6eZo4Avi6aaIypmqqn2x4SZu
UQylpW6tBmLuihXUprYq3hMq+4KzRmh7Z5dPzKZD+m+/ua83A+ZCfRB+Z1A0Qjj4/GSRtmRWdiV5
NMXxonSU29O8WsOCWVgESmyrS3x+nF/Q/Jas+jTAEBG4IZsZlKHJl0pkt+fOrUwYWPeSPo545Xb8
UiXz+vCz//nvxgqka1wr6CcQwLIJBU1Q8C0bbXlikyqVFkR+AvolKbUQG778lvpARdNa2xaOM1S3
kws+9l0tbS1j+Q0/Mu0NQHTJR+80oacx6iGC2DEToCQvzpwkOcGtftqCKs/qkZPYjEJ1nT0Lfdja
5UxWHcH4xtz8EVhZIdx/32lv4M5VUGgxlixXlbXysGPATLjSyeHO7w15fN+us7LHkytsCZzW89wc
4I53bc45st47Xf3V90d4DvaulFNEhgZF7aXKvbR9uPqv5EVZgYFdADny45bSRK2ZhdHf+gNq7f3Q
bB5A031X7Q9tPaAzIZQwsTsAC8aRPTBVOHA0fZWiaFrzU9JM3s+jL8I+bFmA8BEUoZItRa3C0CWQ
2QmwbAz0lTwrJt+ygH/17fnEqgXAsIDTlkiLIsPqriPIocFqyTWdqgEWkiEGAonG1HN0sZwH7afT
LrH1HEiOMudSCycoaiXSwcH0ApklC8HBGdXziPIYtqd7qlUvj50raKfYhqYmaloN37nVHi95+KXg
2QutiRRTiwY2SYWEoG8CoNclkIWO8IHO/B/MtIZoig2Y8VflOGhDbSwqZLEnMhp8HJxt1TXzmAJD
69QyXVEXFyVxHxH0jlAPOJfc8lv4gs2+CdtSYc1zfzdNYjcxD36hWDARwwP7XB+bFLgvUIVW5peC
0aDT7mfxTjuCqZom3bzIwjAsD98oSOnlQT3ooQal+sa3DN8pKdG5Sio+H21p1wSjSq68linAyGaf
RqiME+KgX3/8mxSpwm9GgDQnlawKm53MOUXRjyVsdFVTJegS7JKzfFpfzbi/B+mwOYP/PF9QuJok
Ci8rWs7oyOpP2UVHhW2IxtOwDgnKwTBeZ14cYbmY2dYbrPiil7okOhtMKf+IHjGY2ZzwIwVdhruG
EEPsBgHpl6r3bhOt1UH+XZ4m/Yw+Sbp9VIN2xPKhNqXmHwzhKAKUwxf0k0XSowqU7K+DfbAPW0eJ
LJos9bxIUAcStn0NwKLei53NtbeEtauuZ6w2SaoihyA967Z6YCyoZ1isDkqZzbtQGoynBJv6loGC
lZs6KJSzLpYVtuWknZeFl2GT+7L5xkT5w9jMc94ACHj/ZBGL72HKd6U0Om7SHwUjTbyGfRdBa04w
QWKyNybNxNelxPjXOMpxZ+VjZG4RdqT8zxjVTqpvtYKxcBEC0Uc5svGxD9WvRfvqsJTHVRBomudk
GFqSQDL35rAtC5jnTNn3+jGAYYV5kmE7S4/+BZKVYStVfi7bYYkFxavX+7qDSIDbD8V9QdSTGSiS
dLjvKk2bd2jf7KwFLFmxS+97nsB4RSiipN6H9967R+aGblg3hKb/IktANbo7e1bNQ4h5r6oNzdMO
5y4cpTjvCt6qe9/NGca3k5IROD2DBBph6FChFyw738sZxadB7ov/U9dLZDdqlWJYPBG4Ftpfd+qp
azMQn5GnssRd4bfa667mOsYao/FCrhRRolXatMnqH6uxcyLkNvh7oWEr4aqA3Y2cE/aN9irnFw7y
tvw/EzdKFOxh1leyFe5e6OYCOZXOfvCG7+H0RKRzKmGLSJ8XnPsilLoy0M2RvQMfeZNcTwbeLeT4
QW6khR6hxPH8r9p0bqtZOAq4dqcv75h/Wf2usIXXQhTXqWc1DPc41m+2G7Wo/xNnVM7KmaBqHaX1
9IKtxBCSojuz0tvISLS/mprWne8t/j7ExfcCA+8AFfuz1SVz0KAKvTCwgShqu6fs67BGBhvasj9G
8TylwB059vkOTEdPLybfMOk3P1WwKuYGoXaDp/6+wbhyH1N0W3FCd8JPJYRA5ulQ68Hh4vYxcZeH
FceXWKbxbrDGE+ugTv7vSIra064su3JB/V2mstgZg9IB37i27TVSBhLwuhXclsgWNb6vUF5/GsYH
u885+aiaucBkW4Ds3RhsdrZYdih5v0YoSFaDBHaCuv/RSwxWz9RIBO6D7dZsyXznh+6TG7cCz0E/
S0Gon/5trZYyVe8bgjSPuWSVPJP7qiT7h3MAcNteLXPLMnNY0F9Os8QmFFWVUVoRxMrp+M4vdFAC
Xdlr0HND8ODsQlrI/0Rx/rP0Z+HWclkjJgqvaqGv7Jdp63Ab2i3q6srrPYa6vHwRua4dGxdLdUOy
b0ZPmPQZ5ZB396/pO7sgxpWFc3TpKsiJy+wQB2Erdizj2F8v5M6dsY0ioP+88eWFfDKHOlVhE5Ps
RG9qv7gf8HIdGd1UeV0s7dTnginvfYeJQU1e4Qg0ylghSaG2tbnpyEUxm8QZPBYSR0aKhXqlyWdC
RSydG4aBxnOcp2gOrZsNW42ZVETbYfF59HfKHekNBQ2NvYxCeCjSHwP/700rWFjKKjH6c+qwAJPz
cVXPmeQfnnlBt/kgRo/kfhJ4Uh/XPBlPaGEkzawIH4FZuIqNjAP4kLVeONhOi6qYtSJp/wCa6SGw
QT6fn+DEQ7nX7sta28Qjf4eM1ZSaoUBhDfZZF2G7TKMORXkqFd6h4253gNQGT/MRNOL6l5Q0CV60
i0J9sWErPYlY2F6hGGFuHegfmrsWL1d3JjunjYr3RIOTc2k29HWySLuQGWJprpwfPx9gjFbLjuiv
zx9WY76sVR9etO+RIrda8h0Bp9B7BUO2is+bfvgH5KksQflWU6QZIc/sc77AEXtDLShLLacMrAXq
HToJRolr6WFjjUPzfwW/wnK/VRrobGXP5vAXpyarlsvl8VfJgGUCadPc0fsEsaS7gBJwBs+t5zoZ
1PSOaq+eTAAiVTZeVbE2eh/bTWjmlkEa91XoHLVfjGQmdHDtwxfUHruvdtTJTG11SYm4QOrCvI4I
kU0vUtdO62AFn80AnR/2tsnxYrmP8SZHXDBKZmxxqMV5c/AonJU6if/TNzhOfIe8JMDFXva9w5SB
5bIu1lxaLiVgRDPFLZqgSPdAGupNW/ZSfZjO8FfVwFq+e9QdtGRA4gi3AaQIl2jAd19T7c0yzGUS
WQkjERVqTSRk+MPATIIrjdUhE4C2c9oRnf8UDIigyTttSMSx82nDmO/USL+F2jYzMghzxPx9ZyFV
dn3NZvLHmIdK86PBbh/BsxNHg+LbXXfcE0ZnoqxIsUZA9YcXbzVpttfOsxFsUArppnwcKl6hWpzA
VDjD2iSykjddMVgWt0Xp7uxQ5Vq2V3aEG0RffnVTsBjwXkEQc0F51Fs9DEcmBCbewVZXoBdCNfJ8
lTXZfJ9UuBOHFk5mGfS+c7OEvdEft5LLFbcmRNqENTyl/BVinmR0Cb+hDwPWbbaANrngNq3JN2d5
l5RM81eREu/UGmdJ9HeVeGk9xH2Z6NgGFuHsdOEwAs6i/R3I3ztpJUA3c7HxhrM4o2HxXp5o1axI
ozLr/1jTDtHaW+oIbxSAE61MMHolFZdliPpUJrE+8DmiPaOhlxEjMwz8HJ2ghCj5MxFqI+UurP8M
KdEiOnXwnmd1KTrMXlOERpr4XOiDq5sOb+Jt61MsUrco3Xbl1fFpYt7CFQHawr0Gaz4247Zl2Oq0
ndxm5DAD45UtUyfcwvDciFViIW9HAdrOb4lJNFrp1vuktGkqFP51nXjtPr4bMb1DK8Wh5qUnyRDT
PdzG6P2Po91PhKKKXK4JKhRXUtEw6jQHN25yJesMi1qYEKc2AlpWP772vhwc+CAWNuFgYYHDMXll
rYE30txP/hotkYz3VHhHe0xlOTgMvHMiGFqA+1fJLuDNckFaxbMcg+/wVkF7zqj87m44bAD+1myO
kADLVJx6ajgysi7wDDVM7fnjkNlWYQyDl13q7bTQgN1mNMdwrBJrfdszv00gopdcincgIa0gWKXB
UcBxahnrXPVxfN/F2BTonaK2boMoOkgeUBUGOrB3YzQaseawqKuiDyaHSgPFy9zfv5eeH8wmHXUn
znAdT0P1lcgx0G+DANfZi612Ug/6eV7WyJB8bghddFATbDzwwQLAFXzp3YSjOzJbaif1ZUzO0jAv
50EqIjd7563rixngOFkJ/kz7xyVp6szLhbgxcq4N0sT5wYiqbdRRwz0GKJl8qgLFjqQZcOl51f4O
3joMwV9AUdk2ahn2QlfmjgrZ6tW96ElVJGYrJY8jcMo1EsFkOCj85+ah/RPQqeMUSKLW2V71sHkB
6G0Y67tW8BR+o/N9MMJCgxMqcuPiD1BDjxJem8AcTChmoKWPxKCrCsr/47O8nuk442H+E1dSuh/J
EVrZd+MUE6yaKvGZjw24lBeuwK3LEUcAYcpj3Afo8d7sQwlRzO4NN0muXe+C9cevkdVGSNvG00HH
kRLJrB/Y3pkYU18dw5zhO0Tp8dR/WHxWAWFN9epm3056yfwZFrtq/rU6EJXqYgmRklGTwsdVlS3n
83speSelmAaNUGMYBBZ+l1boisMVujM0xl3Mojy+IRmwonAxwwWB/JzMcYeAUXB9AP5uwyia76/m
aGQoORB/83VptREy8UfOE7WNhzA9RxJLzzi+quhbCeNpkff28t75jQWORp40sCMQXz+YmBTJvu9p
r96kCPMM7LvpkGMlLizFPrNo1Ab165FAtKDzG6o/K8q+dBXeIZrOlKksGFGym8tlLL7pUT/DqVcp
xVylx3V7vU2sDnOnNeTNjzb4SQoh/OjhfF5kA0hoFREJBx/isPEAvuN06R8cYykKJVAci7Gc0T/J
GTjz6SIkAACn/Skos3HZCHZitVdemLWncaGX2zxTRyBU5xy8R5oepsc+0opD97+oI6bPgD/nw2zt
mS3NGx9hew+Mm1LnKHNx6zTdT2eMGKHtNawOsJAbnAA2k2JK/lk+ai2ALo0hVSa2oeZ5W/9fXzZq
KfyoQigcOsHvWefUJq8kLdbboj3xESCK9SrE6/WOPHwXLnQ166H8xyzTmKzULLvwUiztISTF56qW
YiV0eiWMmvUwQJ0PQe6n58Ntb5TcPcMHjy0Sk06jM/s87JNdycdR5TKbI0VBNqfjcSRMh7iATkNy
0t300NGspOjzxyy4Jao8WUguK9RGGbe9ntlIuYU/vZUf7ITBCHqlJn6MEJs0AEtebOrVRsf/EOsh
43rrNRdFqgJYqvkTvy7Gw1iUxG0XMXxZhftLXGXDARUTRMhGDfWTiyeU+BepxZzwshsd2adFhPuQ
HlUS0pRXWAVCjLxqA7wIJNLI87rJGMi9E0NcSBykpqODLv0g/nYLLc8b46toA/GV0a2U/QWi1F40
W3zhmnxhI8LH4EAZvyvXA0xyiySQL3jKiJLAjfv9p36KhBCbU5NFIRU3rDLy8LgKbP9sgMA+fEub
7jcdEWtWZ/16o+VqqPuVAZrl9XEwcLn41AxaFKnZG5S04W4XQjynk5BymVuG/5jnZ/rjhmWMUCrs
kflwFTQskjcRbEXrwOmHXPEicMcIjxH4nD1024N4TKmmhhbtkGANpRHufp5ITGkXqTeyhNrc79RX
GIIuZSp9hjX9LNQoTL35ZbmM5I8FfxBfTfbF8APYoKJdNaB9YwCE1QJjWuS1OkbGOj9C+/81i31v
3+HPpRsbS3KGb/6psJgbyXDzYLFl/T0V8SMAJtaDfqpChCwl2WKOxWZygw6q/NfRXz7LYKpMJOz1
hiJY7YHUiFmF6C4EGLLxi/AToHNS4VYcVAJMekUuOdV72z0EwBlZK3BDYK+V+S4Z8Zys0F9k/E7z
KnROAOxYpDtji1gm2E8KytsawEN1k3/W9m9MyiajiKVKtJkd3h7lSWVVUciR8k3YgpvU3Gwzah+F
8kI6djEb3NwGVf9jMbsGYEXvwROaQlGyDsyHF0qdKl3hBY9clFxbmmGf9La911BMWfN6vt060iz5
5kdsYnjGrb2nmCzWuVGn56LdBgWSVKlaPs5Ik0ZbfYIXK6WXbNycykEl6Xmb2ublmb43KCTRCulJ
E2GrUaXsIfmik/WKdd0bE1TXFtqw1H5G4evBKUV8AJsyLrIlJXGR/+o9q434mPNHlpe1yL3N3R3P
kEaYt6BJ9gU2Ztveoa9ooes+jApG35V9d3RwF/2pzwXCKKfq3Pte+tX0u5M1kPdYA7Z/41E+7owa
XSB2R/iZd5m+dXUV1sBq4qZtNkaAbKfjBoIGl1oWYdS5ftXw7i9PbXWcSBqXSFpEd9vkhpRxUHua
Q9SZhFsA4CCZSIwSP3GWhlXNvNEjpdci9YFWzR6UJC+C824f8RP2eZh/3ZEsIFVhsFoGgoWClLvC
QdfSr2Fhg7duEMVkRclXPwwNvpGjq7jHCpfcCLEj9F4TmhHpx9P4ttz1HpLa3+XvEotbNqMTUt40
5n3dECbToa6XZ5ikfdc8jiam53p3yaWH+sWxH300G3LbPIG/ZnSV/3X/u4txnbro7R0RHrrr76dU
pDhSMCEGIlhUTv1+5WOh2uwChkPI3l+E/bhUv199kjfHNj1G/LRzUuIM3VoF5gKCRttwjpfWv4az
QBsarUaAtZ1v9J9YyrmkZ7raw8hGh9N5qbPNbOZVDfzzfVSkFDa3Gv2rsvO0AdE+Fssgk/ZUolXx
SJZRzomsFVkRxOgczi6Gu8rDDrgcdWkeWguoOaKdxv7Zf6a1izQYdJlWniiR4HBiyAvhnDzchU+0
nvKfvRJ2AyuutD0tsl8ylJ2W+avIv1Oerof+rVD1AeqZj07JhIXuK2OCUoU+LJ0RUfSuEg2EIzdN
GPRmqWyngHCSOgCOw66i/jcOHnwRiJumOhiYAmsnB/ClYZzz3gVfo01at9OqPiKTQTIFRkNTA2ZE
8agNyWy66JA0nwY/liUw6KAa3TA7fJ1luVElOZSYPhcEM6sy5nlCEMUgDoAasbARgjHaWthIczIB
Ai0edd4SeoSVEs2Y99tthmh4oSmYpCSq2jK2sPGXW0cNAeMNY9bBIz6Xhe4nU4I/xBWJAvBBm63L
pESWR9ILzOgnhg7p+yuO8dUu63kEYGSST36BVhLYOAtHIbi83JSH0/E69ESlbLHhOIYHgCGqQq7K
XqBOSH9H4CycJOl+PIu80DLrMechxHYw6/Eerg+VRYwNtRchZ6GyLPsX1VxXOMaVw5lYGKGJsbCT
uyJqJa/guXUIme2MgakJSOcYNY8YETUi5n02G3DbrKMWo9EOUWITSzTz3YjEAuiQJ7/+zP34Kj3v
eVJUhwGwnzOTJCQm55z5x03aISpZdBV9v8buVZxkt/UqCaMREgHiucxk57sWVRCPOafftkZdmQ59
cOa87eOVyRQJk3Q3qt5FKz7ocH/sN0akb0Xu++2KOFmJhLI1qTbcZxFVjI7wv5o/L2zMOxTLBo1S
8/nfOy8hfxV1N4fzksLqJS3JYA555kT8g4/IoPsZD50dMDiuNQTAGVZg/XJB44lrqst8mtHJ8kIU
+qIq2An2oy7SitGe3veUeltKC86X8oJXTOF19ZzznIfc2wF9Cl+ZyRCGXqdpNWmG5N3l/cyVyAhl
tngw+iwZ3aDLNMspQBIc5wRL0xtXUTbllXEE2oI9DtUzYAjXumjiw0sb/WOusN0Qke1KYO824GbL
7Z0QnD//UdHfyxS1C77xp3MMhJa2X+iC5nwPV1JEpisj8pZzonjxdcgY+qhYjWhpbjMMK6cuhh1W
Cp6Z+4C+o2VbePIIWFgjQvyH4LLhcTQVISwzPgwpx9ss08kjwf10qNbPRh3l12XMZf1n0piS/qRr
rNZLFf79RE2hYGDQMe23GP/ZRAPrYB5CkmEsyHT0UckX05DHZYvdbKCVgUGByNxiGHYyTqzcwBcO
NVrEOjJA/SslnhElkC8SHd96nbkzatiymb+CpakkMJ75sL3Bq0PJ/cdkyIA90ByOo+Fm9T/hePAg
zhfrJ9PkvQmYD044b7FH60/GDuoMDvK7Ku1Sednxwq8cEgo+VBQ4AdcpA7aSHTwTnFn3S8Ydvi1D
7LXr390D61Jl9MJeFouT6VwonMfs8reQFehEN9qAjmLMe6Cy2iskuqIJ6Z+4+VoNZonXixo1zZ/t
nm4Lxw+JYj/NTWCQfOUHVEBQl5hKvY/q3rmMNBP9H9RJI8exr4DCXXTX0P8/OhQZcQQeyUtGn3zC
4KXqXHpG4OS+MnIpaGBmt3bgLD5AhaXYFuVQ7dUY9jkDJoKOLTCK4SiTrAktzA8mFl9n1X9ncA1/
SnUSu7RYXc0zoBMZ4TlwdTk1HP1pA18vZ4ZINg3z47um+Dvo9Q8ZGqww5Om65i5q21xLGhDr0LGZ
fTgX+bYJUXjr08ludt2g3E03BUHO8G4/RST8W8gL+2+qY011nSPvjcOH6MJfr6wzcUuxCOBiuPhW
CJtlNits+HEf4XbOjbz4P7Rcwq2hAmKA31Y5BG4ogA0nuOvaXMDt0uK4O82LDpXmYYedo7DGG9rX
kDJbBqsG0IMD8tgHdFZFQYys3ma6O+ZxgCpUA63iEjRWUyZ2OEIfSVGjbrBawftHU5xSauKNC7NE
0IS6N6Y1cwdMuwudb46Dfnib+9crleidpIpfhBNF3X8fxqrg5sgRExxZBvXVDzYLIWqvYZIyQmxr
GFx+BvubFr6mOE7iJADlJFrSrqPB4pbTEQjY4Dyodcz2yv2T+IFAS+lJ2+TNDfjE5mIw4DMp89dP
/bGI4EgAGr7qRZD1a7eZVAIqCEyJKofoKkwpXB+lRqUukNWkyFm4TFzJ4iHfiNJctLueInrsMITC
pcGosZeCS2ULE7G0LNyek9z5QhOqf6CpWGdhHVJeJLDSTGDXy9X77AlXX4i6Nn8ZfKtgfa3m9BPv
5FnYHR73ObP+Mki5OEv33temmWrbt74OUQAUlnx/RfO+ItdOtVsSS5iRWNV2mK2nuJI2nDMbbm3U
9TVghy3QtHkjB2sLVrwZPMiP/gZlS0FhMRrCWCS3/j3DfdI2vMIReasuucFpW3deo+wUhnuDRKQk
jcwm65uGPmlZzIJ/UUPNo+h+OzJvZeB5eDJY0sF5+bVDrilLl1bnQoUJqdDuVDsakRb0W5tgX9Gn
50Or4oLOSlXnhwUseswmK07ZyP/iLjw4Tr8UsEbQc/3OyVPqNVddWlwhWzdYtiTV68FoghiWPM/B
k8LYB07sNS1UX5bSDoP6qd6J+Co7k2ix6Dw017VzPKKZ4gNUjpp3ctL6uj6+1JwR04gZCFqIDUd7
xUHO5PayQlNrdK6UOzhqjZTWKH6Ct/Io7j+GrBDBaOBn2R7YnmisE79sDiwtp19laj+avTLAvwAJ
WBLUkVyIcThhKrDZouiEiqTknWkXsDH/0uL6znjhX8zkifxBmfpthg3zl7tm7CAmMnm96UCmC34m
LSLnP5enomDisqVNQnSZZWR5Jm7Xj1mNp3omUgv7ucQTkG+hyvZlzjBzgN8UZvmIYsQtVcsKsG/W
ANiMVuqVQ9I1odzkjzUVBGFJVkUgtCWKWJQvsJKGBneKCgIkr88AtfYhfTbJLC2tS8hsUz/sHHWB
ZjizXxBGWVdBhT0NSLZH8rjH54u+DW2Ori3BcsIdGeRiAzwjx5bBzORqs4R+zkVCMjXUdPEji8+M
2nIWpZb3sOkKBkckDbqozmnYcanpXYBhGCEBVdo6ieI5jgg4hF5sQhRuhLlP26NZthup3ZWRLYVh
9uIYSmvYiKc9CihJR7FZm3TmyL5teVngkx84DpwmVAGhPzfswIpAdfTTiEC26cYs5QGbffwOlKOn
UagSIl+OJjexPtiJhgmo7nHS+s+VswusUxnrGlsm+SWVsp0Xjy4e5MVFG6LYz9ZWU2f7TT914Als
oRfjFQhG3RHFFK1znNcpbqkuu1XEIkHs2DVpT2FSo1GbXNdfkuTcIJeNV0FjGB1wSMcmIPlMXOAD
OngRLapbCk2Yd2Fhwiv2I1cSYUVoTGFG6oFqtq/7rNmjREeEh0v8ZyzA7oAWf5DN/33jas18R0v4
KH/cfprfzvopZyf0y8gVe1J9zVOTk+Wp/xBOKa3CenZkf4egaeEf2jA3W/DIOKaGTJHakkgC6AX8
hRxNbql0MF4dUAZC5VzsQNsMIvhqd+iQCYbyGrYI0rtPXf7fNONKaWCloYvBp797ihOs2wUYku5W
Dl8iyAmS8QDeivLXOqEk5/ujXvJNXeUl2aGUjqSBpNMnzFmHgOiaiXkRIt3t2FO0H2X1sexsTjCB
tnod0oV5eQzPem4LRefhil9f5ybM7yjrb2vM31+UVAjK/bsZ3C6org1x/TVGdXv3XwpRxqe7/aun
pi4FgGLFX2AGyRNCXzG+1Szv0/7weXqzyjDWBou/ijY/fvLFgdvubYFrgkaZxGVrc6PSQ8ya1bV4
9SDBRK8wDPAuzlRRMay+FKdLXuNaaVyT43ll7P7vJckASBwiXHkZpUJA/QhVMx6j7eezk5zopgCL
q3jSxIYSkNvAdHkXAopOQQFJo5mdMNGR/koDDfNrdg0tTm8TGfhtv6OAcQ8HSbhjSmQvcco1LNWE
URIMFMPVhsqS0QqNoyFrVsSJgncwlt5WeoEmUVJsjmG8O99yYvXBBi5oohUfC7sHuGg1US1Ezth3
BjHKPeVKlba0LHqes5+78WLGVkJLcHjIdlehCC9AygEpVzMVVAG0nsrvGjJz7Ao6RWwpfLi3pJ7W
ihb3cY1ptw+rH1wLYpwhAHYR1+8s5C1d8W50Cfm4TGutUGg1kXRByHa3HDRys5U8s1Szi6XXyWOf
tGzx2ldxTL7CT1FopGNVXyDD7MxU2SOjTAlXBVwC7dZwHktF0jidder4eSe08ktmCw8HpS9i6qfp
9M6ZUfKlYWrKHJA1aQQfkioIB9m39n48+Dt+VuF4Rk2lVTwpTs1teG6ZC78Eso1z6D32Ay4y0NLf
ISV0eNsZtjiqg+jhvyw33bCHmX/WBs9idkEpH7WWwrpFPa/1w4kUEF+mai8/RpeHPGn2nWTSyf3e
i+cWD/yCsgg4a2avDAaoaPjkK14US3j/gspr7UrnuiRl2KCpIXK9S1ag7xcUPZvhK371gW3iXeSO
+tWEL0veGPngRGnkHLGjCk87QBAoVoHr5h0OzwSiNKQ6dxe/yqaWnBVwmoIjqglMIQci6GtuxxYZ
6UI30iFr5+0GDVJf3CTGRE2M4K6WZQYCH373RxSIboyFQujbqLCFJsXetciJMsG95//JFTYYpMQk
P1crcuDLBSlKhpO5yScjcPl9EwPSNr0ITO1eDpQDVf9+heW0wPLthDSGxE7tEvMaHOgjt5HCVMOp
WN2GLZ8IoGslS8CkLE8I0uy9IEe5gQ3bm4rZMllCamr8yCys/Ye2N5bLt4lPws4kUSXG6/JcaFFO
+X8oB3B6VHRjekdfTkah7w+UC6tjeJj+3IIFEP1stylSNmm+8/1bcUx7peAT8lHP3QB8oMH8Wdc7
YGyH36UYmfUieauw3ugLIl1BvqMl/j+L4YWqM8ag2tLXp2x56GvMQw5LRIAOX8HlxOqFUATnbMYV
ROtj918LULDtXeER8flEofI++/n5HESgezJ/tf6e2mKgSjs551Be+NED54ihZ+NjD3vX5wj3E1Mj
p5P53gGtijwAmD3cPDf2De8JFzUd4YdHuNbHFMNYqeZk8ixdbgxZ71kbH0VJUbyhATj5sOxmEZXA
Oun6MHd0nLuzse97TTATRydYf/BNkrGws2fmjRHH4bqb4R/cHAfDS+Fy/aqsVQytzR8liP071i2e
4Sn8v5wyCm1J6fNE97oyRNwZgV+sTLsfXJtnaEp8f1O0SyBRgRRc26uaE2kcegg8oj0hS5tdtMYb
m4b6EaMZLNOWHQVKLnY7s/3WQydo97p1CH8jGMSzjejZgx/B8mhK2UtCiR3UBLOcGYAtsa9NNfUs
XW/NZhpc8mqEije2FULzPWljNV3v785T5Rt5VcgFzU3fML8Lm1jXWHoZq7yBI2NExaxXMr3ECwKU
pFfqqjW3NjoLZ8AcLshesDk2qIUPbJRhK+E9YNYEcfXGIpHSbIa47i22duXx1cFhm3m6icWk9HTk
Wg0di0/miLw8NmJRJpxMKxB4KrJKu3K+/xUVgVkZFg/vSANB6ZrX3oz4gOkk5W7wIz2NSf4a5lyb
LYZBfN/hqfn0Q+p/boHsKC2PnC85qOduVKHKOpwBJL8vGkITD8bBZ/K9tw68JY8kgNZqCi+yl4UY
G5ZVaAfN9ma16qbmgKur3Tglnv/GadQ6WKEw6dZKHkO1OXOQEWXs6PaaxdSSj1C4+uARd2NLzgcN
Z4saEpHL/1GQ6UWcOv9/hpP86/WawZ+X6BjPMh4z7k66DyejpivRiAtRmaOgssQacCs6IvXb1dFB
Z9lJuoMEQQNP2zihrpT/aMGWiBF21g6Dc/At933mfvnRUrUwWaY7SfSx2Llx5BNDM2JAGKsTtzDn
kvUqvuQwqc+0jNjbjJPNX1VGFsdBpn+61CDLLPKjuc8DzOrG3G3M81bOMZpw3MJPrqfv5gC1ePwE
aXHNi6KdZroBZGZ/4Km/16/TzQTeQkYPAtjo/eBU0BXe7XJDErTLUcB969zWuAm1ni15M5GRv4yc
qbRzoFEcmUYLzaM+SrqjQqRMTkKbmBrm4JOPTfqGSJeM5XlJi+KNJ6/op9zTEmHALm6a/4XNoL6w
vs5TF1DtVk6Xc3GcF0oP/SK2r6tS+F3FWqjb08bYchSrUqyUHHCb1MaAJswtel/8zLz5VFD+Y7ML
kYrH19LAYcrW95EXewJDjOh0/mFdf5d1vGh5CnSWRc5v4VtfEh2L5a15ri/fea558psIAAihrFFq
EXgvCv76GbS61UFxSJTzNiASDFtsLFunuoqmoBS1fqYakO2j9P9EWecFKoxSHMhhbE4BMdEMTc8f
fXByHSaXiCcVXFTqWT/6cOlCIm4pTGZJSMx87qQns+HsAQzEfyXxlF5RVIc4wgAsrTVUEbDDvTlb
wZlcNr0g9fmUEwuDsNfpsarXppqZprLzFs4E7FsGH2m6qESq22nlYLRbkunT+t9uP3gCzIfK+bTT
mQt6ebI85p2JwdK7y8btrVbFfpCP9oC4n31fAsYUq7010fqRXyAR/DJC45mOeHJRLf8x3asBG7CD
bqGvTRFPCdfZjOneDtiIHsFFv2lyuZlFmy2eSTKdud0Nn0Pqgzd/vHWI0HP7tb6ADPp5e9IB0SJ8
O1Wn1VlDFN2H4W/WYSGMK8kgJkq6J3DKjyZupLT1XQrjAsjaBXoGSygAPrMijBXTqF83NfuI9/TN
qGZE6tI3TdLCpfVWUoylgr1SwK5eve+/+pwF3nek5kKy1jH1tuEY7t6gXPJr3JfgSMXvfkP6/6Uc
lVcTOcc2qT8bVr8nUpIP+uicfajP1kEqGoO/AY05cim32y894mYtnAkYt6R0wjtxwE56MmtgqO0J
3mirACBJ22DVJzTXk0K+iuo+9F2lhBiI0mOiHd6Mqk1O8AYtk1RsqbrfoD2m99uWPgtR6x6DI6Ak
5Q6LHoUyZTw3P8BNQe01rn76BLxAVNBpMspUeXN75XUO9kird5ai2S3M0EEkr2lLDb7OSKuyndZs
43v352uJsx5ZxorV4STWvjjkoQiuyJq/5jljMVpPxBz3ssLrJxuR6imjtQ43mZs8tJXwBJfibCi7
fPZ2dQQaAgVREw8E6eMADlBpDiJD2LNDX+SBjB1KX0ty9l6ptqllXK53e6hG9+R8MUUE6+znTiyZ
Nh0YT5GaS3Lo0Vo4Q0bj7jDDPUUJG7rUGZQRe53NGmKg4Ju7Gyry241Fyej2TDD+ZjM3GHIN2AIB
su1j+YdI0fhqg0SpUxmIYJW5bhJ39cBpOHPpC7IzMi260eZAjvfk1/CJtNEZH+l8IJB0iZMZIv/g
DmOT1aSobzJzHo807uVDV4NwxQ+8IVXNOpW439ZX30F0IYrJH+nwJQ93Zj0MMNbb5tS4/x0JhCKY
qQhL6x8vGCr4gOc0uZq9AFm5FYtF5bWL8xT+SFcrlB4EcfRtVp0RsTBpP7KzoclnKEVHuLD9STtQ
ilrTDnc6gdMtew/zUnz0ibBKKu29aIb5lT3+eFQ0JPsd/1C9IA1XeRMmvMRfnLSOOFRiotYrAD2N
ufvGGVlrVWhi3m1mb4yuw4VfWD5lB+hHlBl+roXw0T32irNBekk5aIHuvZmJqX0z6NHxuLaFIKdh
XeZdLra+3ey7zK8CUaKyaV3tc5aNY9jQzMCoULRfMpKDcOkzVtkJaYJl7x4bJPa7FPu2rKD11EIi
gF5dA9mULNKeoizuUTT9df5f4xAnpD93t/qTEk2ts+lpcNq8JVYx+6VNDNZ3RMzfTg4qzKL1eYam
/I2fnVQWFzemUEURPD0XycjUW8ik/lqAjOKoIrDAD5eClibsQGRF04xYTGClxb0MuvMmsHgtPXav
D3SOMkrRn+g51qofZVv8u9VqI/GAyPEhEu8h8bsAu6I+v9GI3V3GVlfTHTJE7eI4rcpo4K8UdWU0
72eO4gNt9dInmejXwAJwgfIEwtizUC3uWmLNm4Pm5KPq9nPllmxbAXxVEg/H/N5DftYxc/USB7PR
8CCeNATu/uc4s9uZe9NJtUqHt4oIMnfiA7FyV2xDYWtI/d2/4fmTjjgHe9tUDDiCLa6upPt7Z803
7vJh3wf89QOTMbIH5mkIEykauc7FXhAJRVTLA0FgvDIXlWOt70mUazCERYT+zjn3hnKcV4br7NC+
sCHFHC/HrpVjFcMFvxrA+NSjH9mLUsAYBegKBsAomHweSx88Vg8mWfPYHwtl3DO+6QxAQ9hQQuF0
6kNFfIdRG6+eF4L0CsbBZb2piYpV7TGNefOz5sWXRE8G9iskysjG4SRiGVtTqjJ5TYg+KI9gQ+Uw
5xlHiliNv0iJYxZFMJ7CEvIjffuZLfKg88jztKwW+NkDFTg/cF8exurJpjhB0ubWu0iw2p8T40ZP
Fs5q9h49BaciQbTR9swyRRT53XtRd+qr38HAmNKEHMlpXRx2nTQpXNZvSUArDrTErDsJ7s0sId7W
8ibMXQkMHL9CguKO1wIL3+a2LD9RjbrmTt3TIYzoTq+d3qnViXO+JxieUC2xR0y2fDt0MTjUE7C3
wOIQzWIIr1phPFZypvyyNnWOZyoc1T0dgbzdixo+gkFeJ+8PVdjIWjJwl9FgzZaW9YvO0pIpXYSn
pbqwH0M+rLveGNm5x8nsgbNDMQa93/YVazCie0f/k0CTYFVII/HdSiZg1ZmvrxovGuLDFlhpNAXJ
5vj+FWEyl69A1tzI3OCVzrTl3Poj8h/Y/YYxvgo7Y7ak9Cd/AJ/s4wpFjBR79fQkxHnK1R1gKcEL
UqOYEIONcVmDn4R4yjNSe8KsHGVjIUgCfamQ4e0mJLBP0+bjzsUmo04lrF7Gv2LVHt4BkqMwX1Pj
Swp5xgTSW+o4vbRk92iGUXBkcCLtD6bXXQfpwie8R5SwShGc2q/D2mbmbzL22f7jLMPkY7/HaMvT
qnm3omWhCKS7zQl2zckuyBlYyZHV7ETY2oucxaPnigKEPoXgB3/xq/KD+BGXd5Y9meSqtQX+31Ap
wdqY+rLqd6+9y8QIr9Y+uNojcGD5Saj7+akV5x5GWlhmP81bS4NOmtOKAeMV1JDmJ+A+IfrDC4Zz
zL9utuNHPnK8A0wE+5qQS/HsdA9r2siXONwTG9XlTF5LhcVx3Rdc2hvnUKSgyWvbIxwlQPkvE1KH
uqWuDivS5g5gAkK4P3Wsx7aG+OWew48bscC5GiN6i9MsZa/b1mUiCB0FHpzGqshpB0AjFOa4BsW3
DWpNJD3fCOEH4o7oqUgcBOx9dTlfA/r0HNxkuHCL8hC6xTngTTHDu/pNc8mE4H0YgdT5ru52Zbcb
1pNyFLfS/6IQW2aKUZrHQTW+D10dyzV7O3Zd2BN7LbGy8QwnZaW1HiXrP18OrL/UzZbVM21GBIst
s8aXITj8If20ar8Uqsn8GtbO+fuzNXKh49Mv4wEpNg2OdTgT2BYa6Pt1F0xeBQriqB60cTgoh8XS
dUPDqAfAen4LEHdT6YzPYkAAMai+RBqVBieWAC3xv51bUmf8+2jvz+T9uOxlzWwJgjJTvvKTPMWc
vClfAB2PoTTi/Bt51a8VGF7qG/Bglzw8VVyCJpA3ebP9Gkf3GffVBafa0o3DIr7PocXEfxjGujny
8tSGVgHnueRGjhy1hbpGegQuHXFncIDVl7X/SzTYjtw/KYQJKuhOhwch+I1qPr3wwXIEp5jeyqki
EiZGHGMpsSyctX91rYspKMBzYoucJ8/oqnUS1INfq4RfI2tr0oBrTrmAt5Y7SZDPJT/UuvI+YyX1
+IMaE+h9uZ0JDV969PDG7gttcf6bgDQU4Od3UDef3FpJ7Li495yoc2dLyaX1PSqdaSoRWAMo2jlp
HBuBxywABqmwi9/TSGQxRXtDfx74Mu8WwYSFfFdi/xzPU+naeOBISksCm0Vi5aNLBJEaRrgXM3ES
+3z1zwsiPgW7lNREW4k2066UL1CzchaC+A8ezrWLFxMUNFdbz0Ep7QdE6IYFyMuZ62VkGDgzDdTB
4jK3l4ppmeeNKQrNjnB6qKKlp9zGoiGbxCkZfX0m0I/MS59BfIKYgUdYFRmZg3ERB+S4u2uMafOb
iwX8UWaWe/IJ/wre3MtjpRebEeGdGBgw+QsiGemKf9s3z0aqKViUs0meN6/lJNnrGSCOSklJ+ofl
SVh0Nl5mQdat0TJeLBYTurdAkMk9FbqVtLaQxdV4ivFkovmezx6k7N6jgCyu4J3zEonjuIHfGzF3
yWpBfm1gR3JYSgQ2722TFtBq4iZVNerfpSXDnM2V7rUsbpAVNUqAdrg/jICbYg0Hlz8mtdfl+yH6
0UNWGtySFxS0SHvrYfT16H0DIEVIdz4khsT+aYTHCXnaQJmwurxXjagIsFOBG1KFhkHpGdDvczWF
8zyAeK4JSi9P/2xC81BDmIv0Agys2SLbjiAH3bLNdBRkGs7ZyM/qXTvnXyNvaB4y4rdBSCZA7ufh
WrcxHkmewY1qM32VFhda/ABNMT4G101FOwssO0zewEauBzexi+44P2x+A6558wkSNfxaatZWBU+7
0W5vHRcIT21tJgDIJSIIM8uYotYN/q5mwrzZspspmfbzH4w/Mv3SWYv3YafeXHb2BYOAOgv9J3Wy
6UuGWf/haZUZWS5t5BDmVaL1whD0ik8cC6+8/eR4f4o+3MFySQ6lRD9dUi5rqloesUXfTS1tIkJV
mxvgkP9O8R1Wn8kAj6gRjjkBZck9IBi4IqcPER77OAw9Cle7Jx1oY1gILQ8Rb/XHtkcTtOJpI8Sz
GDXObWRh4fjiS9W8Fs91lRPYk5W8MVBzxmA8/ffgZ1XtA25/iH7qpJPe75viBMZYdEKAaUjtVrz3
XNGqinFFYm3n/KJdFQJctZR1INmcflnseORxclEIw5HaTN5buCddx0rJZXkBTnAgF9CIqnFZ9FW/
Uoawr5HNPA8ON4NDTsRtODzhKV0e6JT8L2eCWE+Ia3zZZrTWGeFIjwoijpONEfd1dtRyQPmSLJzX
AyXiejjy25NGFiW3gIa0+k+qePxj7kTmkfTRoZSmq3Xi9hs/L1se99bzJFHEIuU6WeKH7KyrCvqf
5hp1aSAq6Uut3i9sSfhppdI0SJzeFFG/zz5sEpYQyVD4XkwgyhE/j8dGgcedqpPk0VMONEKZPJnf
E76N17WB2ZefNvS6vvpIobA6wooy6ljb9NptVj17Ml6fbrMm2ca/20DWb8qBlzBDR8+mcTOyQYQQ
1X5f/Eu4WLYwESg6cVAR1O75BITIUHiDa4lvjx1A+fmTQvCMO7Lcw+ibz5L3WDoCWNG78WghJkN/
XL0lpnUUZfG9IlQlS8eH89iLW+6xavG/m2Ts65MG64uki119AEylNfvirwawoRUG+HOKJj6hTPSx
8symRMFCoM27Q0ejR5MLkrnm1wipcRD+eBjMYRTVHNG5CQwHK+ekNosgxNYy4xQKX1iigFVndB4z
kgF3kuMX4S01dP+n/doMzA3cHXHO6MAAKey7DFd/zgAk2gFJSI6d2EwI20exLhMYacEy4wLtEvIA
W/qsdYE35xXwLMhdY2mIIDFm6Iqc9heADeYjPunaOG/3M2mzzIgkAlH1tjGqQ+QhN9eko0NZ/ZQD
vyOqNCm5lMEJzAPhGWjmkudGspadIcdIXcpa1cmMW5n99AocPT1455Fu35h9C9zd+WTk42JRxiB0
GF0Jr7oiSj9hKkGlu9iMojWSvoSLNsLQxk4k33e5Cng7CIj2Iqr9bndYKuasPS7FTR/e73dV5H5B
LTK9PD368TR+aHT4mP/T3E2OtX3PaxdmmlmgEkGINTfESiWe/ehHR9JSRlbiClYX8IJKq/IUtiEm
tBNts6D3N1zhyX+0NElkhuXU/m6xpC6VV1YzsGdsrehBmu4kJ0/uZgdXXQbG7CV5xqWIbPex+EKl
hfQ0WNzBCAujMoQ/rcVgdg40EyTN/ShEjTmWIHse1azLVSiWf6DcDU5MHznmI1pxoSDmX81UK1p7
sj/Ud2seI1B258TbnsgB6/bpDCUeacO1wZ5Jaw5MEs6VqK8Dq0b1K7GuFAQusQ+LTZYjTe/7jpFI
S+mtXATr/FUHVvuw1Taezk4QMx19NHVIRfy+dXBaoCiOfs5rmk7BpO+452CuT/6dmeUKxb9VwM1Q
t4nQw0XA4LbL0YGrFRkXcxwBC8pZG5VeeKkdgmjgeB0Wfy0p7T7CndxaZ5GDIM2A4pvVaT9pyqLl
JQ5UWngZKKn23vH5sm//+CFADP4urM4sPRotJhZWU3dMbICnroiN8ZZNqGrSmvVgU2s2zPzvGMpv
VD0QrRVi9vPeQA9X7DK1VKniLOWtBJKuu/bTsRn0jLaLDbFyVFNQ3JWqrNuFhdBQQ+cCKCWp6Gyz
9L2y7TgAH7FKZqQtSurlwv/BkvWaE7+HZhO95knZOaAA/O/sd/I5xuu1/YHAC2DYw7rT6c0AvNRN
E84BqwgKGES3jOxbQWnFHG4Fq68qAwigDG1VcSUgNoH3X2zfJEmkhOnHO6+VS0lZ2XdzLt3BlgHv
LXh9662IrN/a5phCJx/u1cnjQZIYUiOOBPTCABeVQXQrmrcV0cY9LPYI/IBYDlHcNe+omh83tqmJ
u+i3PuhEup4rfFbOvfyNmTvcIgjGEO/pY3suOcLVjf+YApOB/gqR8stXiPFbUV0+6+Y40kACSHY3
NFTKlrzZ+YylXAuq5aftrMtebBR4/4BPWwud3rcknDkm+xSkCxKXs+epXyhP7NzQZyoQUw/JiY59
hOg+udh5lBKVQTqXTGqe9NJjz+VC/DDw2xeKjRgnYqoVL/FS3B6lGeTUJt4tkXWDBy8Z6lz5Odjw
+K7IfX9iqpKz8/tCfxfb35ODh5h6lQAW++86iy5As3Rz0GpFmAdwxYT0NuwkPI+0eN/PZ/0MCCQs
V/4x4KO1pn98ECYLA6avd9+Q3vJw6J84EmWaFunqpR2zhdlH8l523IhaLkL+Lmr/quB7BRDgL3Wo
u/gViIFJxTPLe4ou4pDKjwpQWnFid3PGcP4mr6no424PM8u6YqO6bwQD2lGkym5LU+b8h8Y6Y4F9
rQwO/3DJfnvvyZ7EK3JgM1Jsetv7/9KlDhyKCzjDg9tEDklSwV3QzPR7NSgD7YpEwe6RanGL1FoG
mwmLc1RFUmRFx/mRzfkxyN0m5uxd//a4rAQKIcu1BnqwGGzQrJBpEkn6Uuru1MeBNtLtdKbHQqWi
9n18PmC5Wqd83WrphqFsprFobO/VbWB9ircvCxMEkD0wSjDL7DWKtqByHkYbiX0Ca5Y4s/tnR9/W
PXV5pwjJ0dFKjIwUAzrLUKcgIq5/U87Gcfpni+8xb9H+rFoys8vMXliZV+qTwrsFobwaRnzuBoFt
+wrSu4/snU2x+gX7Ue2rrqpmxO/saNEp18+6X8bKTmSu4WlXHyYptsOKussqmg606StogSXX01uG
V8CCohkm8uIPDtLlybGyILg86ng+jZEuzUn+jC7BNe+4vOpR2oNp1hChdZBwcZaqxGY6TS4wJe6S
RnKrXliZXkvUZk7rxOzewQDlZTaXGBAbfvE1okSyv6bVmISE5h4VbxOUBtTDmGFx05KyAmW+aEb8
fBXddB+KncGNASb3vZm3WbKbqV45u82BcHMHzRI8WjslVFX/d/YmaK6m0uoIWWg84lKtcYHcK9R9
elTXLLDhl0MlA9hhDEZZzy7U8ytOzNbt+wUiwIDKMHFfxus9dTSvxYjd2l4hKqecN2BYb8W8m/XL
86FlLBp1j7ioMjiz7kAjwMnMHGYajG62g72eV4Uxu3YylwMSuDgoctXlldeQZ4MR2HEieSQZgIWi
cPbYncUVU+6GndgSMIttOdu0vwMzKoKoQkjKCyFBUnL8tHBnMNzMZPJynHqu2FziaksbKsp+RKDm
LRoVbGNcOCISdl6kXPbKBZyut1e5jT4yZqn/pmJ5fgdLxN3yfpEemZnICpVQYH3YcBTxEbOrvAs6
AQkd1N7agigZeS5ZQK5ppKGqDJXlmimpb80dMMzNI5A+sSwKmwT7KPZfWO9li793D0V2hfyta4Nk
FUaSPlWrT+nqPwlgF2B35ZfGRYyF8FJH/hIwIuw8EOgub8YWiLRCZsE9GHUgQhmOo6zEq7ttW4l5
XGct2Fa6pKlZ+3bQWrUL1/8O5CaJYuA2DPfAg37DuYu2n+EVLtADmldc2plGYDShEc06RnviB/2l
q3x4+WwAb+XUPdrSDai5RGr0DgJ2DEYvoS5tw+Rh42YDvaU0+znxDvSdxppoGpU2X9QsdAZ5Xuml
r8Z+nLqi5/M4pWxuHQXdBC0UvR8tKJNUZ0RP6efBf3Von4o3+oqd5Cc1T0kOzEv4NCLuTSo+lwXj
lCD008tKxP2YcVBTCH+vup3AQUy/LukAEeDPafuLzEAqe9N+rIVQM6299QRZVpzXQxqSLF9pbuZd
8DGsBbaZ5W2mrYrP7UHMMskBEKMJfxOjEkgbPjj96dHIJ7uQ3YKsDJcX6+pHbr1/zwKYJVQAKM7k
N8V9A+s+Lc8+Lr8cW/D5GKBhecVaKlsRLiWtx7KXQMxA+vwx0fVHmIthKgXrkrhYXzcpHRFX14Wq
pFZS4uuiMFpdors1N+BQlp/BUlXfwWW0DWoq4J1xKhgcink6TNVRAGcrmmWCLRxSAWYp6cAXbgrp
8o6CpnENvrFfjY4LveMYT1VSvcHNiE1O0d8tC/3Cy4hn064p08D3MhezojlV1ScnIYJVLyiUE/cc
V6Wf/Su0LFGNgjzMO1QhQfj6Cgtbt90jCjvEdA2uwN3oxI5zD6jbAsF0k0Jet9fwNI2iWxJRltEc
vaYw+NNtIpduBcqp+sLJ3a1vV++DAU0HwIaYh2qUk48KADUQm2A7ox6w57b1pvAJcwloDKT8t/g6
sMMR0sK3sk84Bd2buQ8BEFF4HAwkAAcRyUD9B20drlqg6DIQ+31kEmlGfKW/JHjvOQiaH28S5Ogx
A0Zp7T7RpAKuGixESmAhX8bhITOuGx6NnGfY/N1vWjFM3Lqe3becDLHrGQdLMhYjm5WCgTmZgB5H
JlDXUptBVZh+0pYsW+a79FIpiamFjrb7xd9bJqJrpqaBDYH60ZEO08QYyqX7+IBg4pTy3xs3EkrK
A9YIWrhWNFdF1RVrc6yF8zEKnYAqkdKePJeZG28GsGJrR+obTHML4GAjuFnE9Qr/obXd21SuuRYK
ciPsVPG5+yxUNeCjNUIuUZjTMavCD5q1U8G3X5fMKtY28CyxRrDtg0HhqRAc8L2X/ydcyc7XMGqM
ZiiTN5H0pj9GBvD9cM5exVlU0TPzkXZuZVFZ43xY+A7j6OA+A2eCQKvNQm443bsmslbtaRF+a1Bx
YOu4q+TWkijgf1WdjpSut4enSVvWO/8UtsWtoJ6Qm88spfXp52O16Ohe4DYSkXNsO8DtsUjV6TUz
AVtRXsjyRCqtOag39YUUJRbjJKWLdde778IIBVQmcWivKeXwhKthekKMqTduQvh983b1DCE95MIi
8g6w5SDGuAe2FvfRqNSJ3uwRzJektVJSOX3pcL3JqItXD9c4HT6MI+Mq33p4fzy6OkE6FfktQ63a
Xs17fZ/3aubVfvecP5jUf4/6MyuPkBZlq8WoFnZevlSHmdwAY2ONNb3HRc6hOMK7dBeSDJ9wrerE
PCCsvbHo5KotV1jfCivL9PduKoMVaSRkumiytjGt4w6jXiP6GKi9TM+Z9zDvSzbebwIbcgYRpZox
mUsiIZrW/jGOSbNXEPFex/2h9z2REDSkZqvZthWAZNrmtUFN4XfahcnOy98qEGdVEQbFyBAhtkg+
BZNpCRvQalYPwGoo85cM4nqQbwfEluy011ATnu390WcNAoMdax7poE1GVIsqdpcVt+/l89Rq5B58
A5/EU2QN9tL0yW/8MWqdRZbx80vAPq9ara8M/Pk/x8LFMYZMEn1jt6XeN+israQ8SKmOSLskBY70
MI7UHdHlMhnwFgz6t/wW1cNGagwPTbfT7xdY3wFkK6ubQuzhjHG3D/05WuZXkoIjgMCCVGYF7b8z
AWkguuRXE5eCs3FWza52siW6THzwraEvDy8tKvm5NB8Q/Nc62OpnyprclOW11qrjWXO9YkfqYHDl
mmXPcEtvdIUAos+oc7Qc3xaRyUJH16F1EEUkaMNRTh+N5miWbQOHaypzWKOHRIxUG0awExpVWxFK
z0G39vyviBRSrHkcKxNIF64mqLFnUfMlLYbiguduB9Ki8EV5y5oPF85KRwXSJIiFaL51WZa5dFTU
4pD74yq702rAa07exEnWAHA32l9s9hqZUpyHl2a2kJhLfJ0cUgP6tbOwTsO4A7MrwWaNJYFu9P+I
LhSqOyOk2E/GCsbLmj3ak4XYrfkwrb+1keaN8eEv+sPx9jnTN4Nto8NqTHWQRejdpW4Eh8Tb3PDv
t0V2OXZ5NsoVxBf3jQsks+I+6YqDYpGEVf3k+5BE8HJvKxkchzUiA6bn8MjGRHFLHagO+lye8mMS
RCvb8arbLLDICXFCw7HoQeE61bALHY1lupQ7qtKyet4TDlwXIw7bFpCCuXrMI1OJc4nkVsnxBNwY
28RbgubiZAP5H0DO6TBhHvrge1XJkjU1t9B8PhMIlbea5QO4G32E25kqiN1HxmB6wfAMFXrk0HZO
o/cnwPYTbz5PsqNzS9c8EFQ6Kr4YTP6yzt3Nl1A/y1pgxvN3LP6cH4CBZ56jProTeC+rCnG2qWhu
Cc78VXBgidMjI6fY/920QJdVNNq3PlVnHrmXDRQZbRK4T+JcZbsA3/dqZ3KcphqzVWKt89u85Inp
07AM3p6Kw9DFUm7eQ3gYmDPNMap8ktYUhFE50snVhYDIz4upTtekGfQdEEzWJt8p6+9k/HSV4D9A
Ddv6ls0JTbINzNFUr0Ua3NwHsF4COll04Z7qG0tqTy9gog6B+kG4wY9DQjfrvPJVWLT0rqgZVQ0j
KD06xgx9BF0k5KGm20lSX8F0rNFJvUYCXSiGJ8rbF5FaZWmi30AAM38U1y0Dxnr4Wh1SDaql3RWq
zOlvXNB8yCQIBOHtMDKtvDW0XeWO9Hdc/I8NvGyEDFJWtbpqN5Fs615PehLBAeQwe1xs6M5KtVtx
Ind/lfdvqs5BM6lBpkX2zMrqrgSE+skwOHmgVZrMLUg1VV8uXJZeG7k24z/SFoxpugKiLwd8qbN+
RHGadcI9Eq7Ndl1Uc3kS1J0pgjiI0gzZzIMhyXtK7gQcUtJodM/NNqWNnDzfFxBmtlICOCpmPnsX
3zQEHkE6AiOrWB0g7tGStCSfJdP4LHK2tb4UQp2rqDFLNePOMnYv3ocrj/+R5RjZYMw/0/mp9tpl
PYuoaUGuB8EsCznOk/gg0hbnD9HIBNowSwqXR0yip6wDEBo6YRUbbf5no1aeA3/kLFjb5TqYiacX
6MpFO0jXyGWn6UsS4GtbKEMsmWxTe3muu2eOstszu6sddODAnWWexICvXcNS2Q/7nmpVscdTlNZv
FfQL2+RrSU50Kam0iRO9ihjRL12i2MxNl0za49gHJS7WnbKtqOv1OAY9AqvqnnC1KklH1pKxQKMh
Nls2pbvLDRNlEVEiKq56yEBsiSzcMWb+JT9coiVRjQpp3P0Efyf28ISqkCSi/LnuxDlpnNGW4wA0
4NT79HEYB29z8Nai47FOUSWg5ILObwRhnDTKHtsr2B56j9Lc2/qVOwofEuShBja1ElKaa/BWfLzY
187FHdOyvUXjtpylv+KCSmvZOXbnRtmyVOFwDKBx52XoLRf0h8MShtFhcsmPRbBOQcKO3id9nEgO
sT4A/oAdVXWasex88T6XHtyZ4TSIUnOOItbHLUND0A5ya+kUzUsz5ERejZSGef9D2uNhNXn8otgN
SMg8u9ZOybehqyPx0KhS6pPtT7+eG47juS/ObtSnhSF4PUeBt2Rbo2DFOOBghOQv8PU71vHreGq7
cyx/j7JVFtFJjLYdGkNmy0UzJ/P86Y/xFgzWGNTOJou0cHOosF10RhDeP+VAsbh844frPX7eLjZ0
+mDz/JNk8Y0J6+TVpjmV6BnTCYDDo8ucYqFGXTGvQTAWV8sCGbWb+Xh6CsdxmSNCZAuKf9EV7HoC
GFcWmaLa6eJ4lBk70qPicmwPVJ7ECmy10iYSnTs3tauJp6eLRpl/vlDFhci3ivJ9xNAppnIYHKLp
dNeDqh59VYlHkqhAK6XvDS5CR0RgeimmgPpJz65vlEVFJEd8lVvybCoiW4T5W6ig2KOgl+6GocRi
7HeF22jSE8Iurw79F+MFZkwz55ThkIZkHYnYryP5lv78Z+QL3d1HD+A4OkLaS9MARCs0yl3lQHu+
TbOEbxN+jSB1qHk3f+0sYU5tjVhqHlQM1ilOYzE96hxcb2Q+O8uReoaYQu0lwNJPVW75jGlN5u6M
v63Zk9MJOdzVQteRsMgdY7HTE+ScYPdcv35A3UZZvvR0AGJawnPPh9Xy+GhJZ+oR4HGUMAVnpeay
2llFJE1Msaq9GCxyEZd57jFAP50QJD1JQ53mZj+EH4ucnhXV4TJ6MMK71R1p23z2oShuZhBvQ6Ih
fup+xo61AWwvepCMXGnADAaNJkWZQf+7drnXeGS0/N7+S0NsB9CuFMZ9vICb23Akw57TOndT/i88
WFU+y7jCl7x879ld7aidyv3e2q4Fjdc9GrHFz1bN5d7Msdc7s6J3HMOeZnuoIoGUwwae6cCG7/OK
IEf5TFs8z/R552w59hqg9Uya4M2T3siYeGpru5nTGzFKyREj+XXMu4GKiVE7XVxwoWZ2ywbL30Px
BYsOXG54cPphyDKOd6TaVAYSserwvCwlqfCQZxDBMFAjQPdQh+BfmkLEMx1qDCT6KOUQdDQWX0Va
YhWK3sxp67NZurX77XK8Z9Q7g9414Dqiqds8SoPiX+VOf4SRsH+OuF0aIsZGPn165C0fgiryMnaW
FZBLMpHICnSqcidOdL9do+b2nG3r0uRGHFLbxbmaK7DdEBzO6crPHMHuRPmGYVwW9NEAmfaRdvbf
ImiS2aFNxEHFvH5qLAx6cCmKLPlSH1dQ1WGpTLq6PSJoxi5onPVdrxtORe6n8iBXQ5fJ7814GTKI
2CPNbxy0L5za7462RAo3OqEduuoW64mPoH0cz9cGX7rcDjRMf18cOp99b2PmuL30EigUBP+xBzKC
rHPEuIRMHQ/sadjxBoHCjz9+5goW9+oQVJCJewcpAKYHdRbt29o+lqOg3xXngG8k3PzGlFBI2RdV
mNHZKNCylcQxVol24ERYB3rMDfi6cNcj64fsCla2A05DE9oGv9eXTe/eKpZ7N8lifkJa3xGIdrca
Izm1J2j/LjKhYkvNO9i0Co5whBxBqbMT+jtGTU7KBdqJKhRvEpIHKYrXnN7kY0KBx9LyxLwoYWn8
18ChdiqwcYgImI7S1ecdZH40BJT3D/CMGRUVXAD/kGiYe6xW5YsQb3yL0LLrBUWLUVvnsUoWxfZO
9+4GqnMHH8ZnXuNcYUeS+1SvDKm1E9uQehTaifa5J4DU2VgsrBScjjbqYwY0Ox3Bw8xOFj+gFure
47icGX1/uSa7azrK4qv7Ve3VzP1ueVLvS4UjfihQSHSveQ9hMPyKVTXpLD3R0OZkxZtQTm5me7u+
s25k2Ft0FigKNRXG74K4p+8PsYE1Bu/2+jx+QjsDaM5iee7LIj0hQaKv3W383xhiV7ljI7qm1k4F
BqDhkHsr1G238oxLEOaAUEQ98CquV4FnYCLKOMpaDi7+PQAvXhrnbNQHhu8CGLJD/RvEXtbu8FHU
0HKuFe6cVicgdYZkHF8msEEZW1h76O37bUSXq0V87s7KUoTlgo8G0ajuMt9Vjayq+TE3DLJoms62
syOSj2mvOh7p7O1cIHIcKC1acztzmzfvqRIiIN0ydOkWWpFZRq+sEMBbKlYMAJmYHFRsj4ewG4cp
pmNz6vPOng/1BXPWQoIL2L7LqrAd8yeoWAE5HPfx1q/uegwmDtadhjKMhHiRaPc3Bbvnwj4rgHsv
52j1fb6AX4qY49b2N0Nxt6DsyY+z581f1HofAUhTeA8192/eWcAA5E5vFDYHMJCf+RD68BgN1i0L
bMDOjenuuo0tB7wXx/4RM2pDMllxHHWhHCAac9glOXITcvGjd684ioTVwnWzOWhBExypxjbA0orz
ePUcCE6FDQRfP12Yi5vZS0IxdWiuHoNEUIVpA8in4DBAsvcDfXdLzyD2emyxkeETpawnCcti91YS
BuW3gGjjehi39b9Ut84kB0TY9XT50oFrsY6cExgUjHyQ9QnyuBqpQ3Z5+SZjgU4eNbzSZpcF+ynZ
Z6fuZam1XZ6XITeWV0B+xbAojmF/9cd6a1u7y4XW27Vs6xv4EWIpGQ69vVilKicQDURtEQY8Itkj
CrHT+YP1akAs1gjDtep6l7zNHVJNReyV10r/JsvB9vMgU7tQryiBAZoXG29RmBCqGnzlEWyCRBee
54axWM0jHQzd4C3ZROrXE1283Jj65veQe9tRsv+DzyAlghue/vrNSr9dTA34h5+H922zeF2No6AA
QFnknQ7o37J3BthzxTcQDJaW6N/qMEDv6u/T0iPf4wjn13iDCWO9/maOOQuAjfeDX64FKeA5/VS8
uIbeg0XOwP3VOyTzQ/gC+yJ28sYm+NKSCtlZ3M3ew4FwW5bbU+Md6ZLJZRL7LJ5o1wN4OTjBjU0h
M3ssUdjw5lvYJjztkYR/N/O3t4o6ulfGlZMp6Y6ZY5ogDFQaE0RzjoRjRP/MSUJrH5Bb8ySKjvUx
DKzBWS2hFgTkYvW7WIhNQoZHIIMIvqIXld0AST4PtQWtnWS88Ej4ECl2YrwpBs3yH6YOgO06efnm
wuGjBjl3R95k9v1R1eSwf7NZypTTOa76Mq71XZs9FDdnsqRSWwx5toL/ukUd8ZaetS+khgaWocPg
Oe6YHyFrZbaFaGgxHemEhrkP4mYIHTHabU+Wld5996g6cT2NstXQuSvs+9P7CdbvazABgUzZFYhQ
NI1O8mGWdPFTjAq7IDlAaPSlG9tFRLuV55v6XDRohiT8hd73ejSEXZGKVeihegVAT08d1EXR9Xom
XIvN3vmdB8dNWAqxi/DlhsRuy4LESsMwp/JEoFASgcOhgauu1NdIyNbVEOgEAXAm2l2gb8bi7FqZ
psO624xuRebvpnxs9DBdzyCd9V/T2GmdX+5KqUy5V3kL95C2KuZoDFUcJtMZC4Yb0w+rRNyTGkaP
wt3OulgeDPtrGMizTN3KqzxcRXNPFCVB46y5uXwYr/71WIwZVFAJYcnUadGOLhYPkBE4YnYm7dS9
2fAMtyg03iKOu9TCOQhoLd4s4lAA7iyf2AW1t3zTW9B1rYmC0pHQGD5LAaQ0Tyo2dqE0V4c4gdh2
34pff1xEpyUCEQeqp/YzNed49Vl6/e/E5tTL6ilNYC8d9Sq2REVMVPeh9E/36/cn13+Flp3/OZM2
PNyqi5II625mJwTFgKg8K9rn6R4k8CKTXyuu/ZqK82J60pdU0jSn+UrDx6Dx+mdci+gyJuFjB4EE
tXz+kf9gyOOTOcFz7mHTG4vFYbSsUYGhgNKiCnUXCvmqGnCIhnmuGpGTgTbbmZGdx7CsFaviVyX+
C+eXgbDMfYGD37IAu2IaTyb4Rn3AGK4kZimnz0owhFo6xm19lfZNMlqieLSsFejApuYgHgJ2wo0O
gYk7Iduk5dkiwq0skDY9Qg9p/wdy/9+MomyltBUF/CrKSduXH2doV72R0NblQmJ3KxHV9pUfs2HI
URp9neGVP+S/UklAP4YwE/R8ug8tl2ZYQt8cq572o8NbCYqOXcZ3Ii9Jf7F7Gck3tSnBYZaHv6xA
iC2Wt+Jj9K+YKG9rluHvS+ewCqh0Xvon/MPV0sejcuKIDrLkedz0aG836HWxOwXOPe+vNo6qW2YK
mQSvKxwL9UFzbjCNn1uDI4Mst+JWpU6mjKxICYHuE/S/E6krvgTkUosnEbbnDq+ZgiaFhV+ApQvF
oGgM/vARQ/T1ilHCJLFzHIz5dAVTf5ybHoRg4U7EbHyHQHCjO+uymfZzZbUep7To6X7Iwi/OtVdW
8UmO94FOfsokXJ61vK623qBlEAz0SE31Q3drhqG0OuOYH2yKRf2sPLILsrmO2bFHfXN43kWFJgP7
L4coZMKxHUgJRN0LorhJTP4AsDqoSRmz8P/hG9lzMkq2qhu8zJv+hWMo+AKMV+K4aailmbN7oklL
iOY8XRsVK9hblEX4KphLCq94gz2TjJZzlLfHrPhSF6G2WteB1cpB0Xs9iQP88QdN7W923RwQmKgO
QmW2HitkINX9xFxv1QJKEBkwAUdSz1kHLIkmOflem+257E2flLowhUm0XlC99A9lelmChWkBznyC
Of9P6ldgaA6u3aHQ3yrW1/J409Raay7h5atjNFL4mgcTC72ncTbkHbw0OhugC+YpDxANAEhFGU6r
eKsJ3YUnzCO+A01uJl5m20/G1bueqiyvuULN0g3vU8z1Z43JzrD8DbIw92KZ+Ww1RHHi2CsouyVx
WjFuWr44ba5VfdNoJW54wh8BLGufmMrLgxfx/11tWWLC93HoWGroIHN58lNrYafCslIAi91AuJwl
WO7iEjfq6aFKtSZE1zpQ/T8YzbCRz2l3PXU0rFCQiAhTBilO+zdnxhzdna9Wc0nNT//F9+mA/jPz
bGWIvRru09MpaUhhImZUgoN5+0UVMPZDqIAHEu3pO4gt00LQf0lkvSU3UnL8eJMQhk9Y6vR4EgAq
yovsqKtKrXIaCmf9POQdgx2Sek4bHOzZ6ts5veWEA1DTH2uVUhY1jERqlAxC8Cam5rli8yU/jCtT
x0J9sLF1lb/1DEA1rk4JzNobv2wcyKdiM4iFydU/4auzejCkk7Xc+x6XTBIO6kGTzjotcWKBSyke
J9Sv94bTi1X2wJGEw0WaTwFPMmlBlnLwp8MwjgRgSbGGQxvtV+TkoQ5ycW7Mpvmm+UswaNwsBFWl
J3OqhuVg10y+rpJo0LCABsFh0UL5mn3GqR6RQiL1ovx2B3MPcK1Eh8dJE0voqlT16qfikcrBivGA
A3xSGf3WSo3iKddJlo926OfriQ35vekVqKyvEifCmQScgHV+EdesnGqTJ+tq09nEDLgAQZ6fLyP7
tIf4a0GcQjyCmyRt1GzxQtzD+zeV5E8uShJKQYLXeF2mcqkUMlihjvVIU12IUx+yYEFxcjCchGec
bW85j+nqM+HxqUsLxSOz+l/tKMfN71FeS3T7b5ZsCiOKa1n4J4Lo6tI+f4+k5/mc+EQoXtLvPOxF
WuQWijyJsL/26NOR/KwIQuhSgUzPWAdT+MQYL3XL1JG1027RXGqMJx8pJBn5U8mb2A7G+Em8dK6s
0du+yjakkgSWDDisRLGvun0FK52mMAT7dTOrcrATUA3QewmOwn5jHlKgTxAKJNpx6bs7PUPrARZ3
2UYncsjuVExRXNgPnfOsIC/wb7L91yhlERVKEYxvumsdMNKoIjXNUeU7mZNA76bWnGbnMXX+9oRb
VxWj1sZgpxd077a5lbm8VAa7rUQOannQCJMAasX+0cExSMSlyT46Jfm706t5FhVHCnLzb+x2Y1C0
INV4g5BXIbC9+155L8AyR2hsvOK5dxvaEpYfsR7iik+jZ91Y+TSAnL9dPquz/VZMQO7iZt5pMll7
cq04eK3g7KEKLDBTlywA1dd4Y532l+eZSbGnLkEEeCIFKT/DVlsC52qXZQ/2X8OONQqQ8+SZ76il
nJ6KBXrJpdKPweV6nR2VF4nMNpR+mTxQw4RtDHtRZY7Kl7N3bQneJGwTotzSfR7x3WQfwa7B7iKM
NS/fHUuKTGMwN8kv9LwxeGaEZdEF/WWMnUtxFwdnYtcMkpjURlpeQP6Hy2nTM4O2lKAZjliiOs/D
i/DVG0jR4cdCRVSvzXkRGVUNsqSvto6+pu70QiHa35XfsU/cihh7RfGxvpt5duDBVObEEguJeHoU
wssOCtfz3dlai9mYsxtTetqqOMYopt6xPQeOar5bJCXN7B9zQFTiq91sWNn7H2qksuqv6B/U6q9F
7m/3uVlzuVVgfabLup31HXfRkIvoiqix+x5b9k22RvLlS+Yd2kLXp1fz+DheaitDMK1uLhG7ohNX
qDxVp8FrGDKxk8tqsXh/LAltdYh6sWl34WMtlfqgUj1r5ALayhktv8K4GgjrHPOL/jrOC/hvS5Cw
tHRw8okPUI9z7Y6EYak3XkrNw9stT782oSbPbaxxtoiI6FaZvj/hLH8wAWWOUomM6Hiz1t8X31wn
GTtFVU6k11St6FXuqFnjoYsfE0ukUaYHWPExvmFje+AkwXsBR2MrA723DoAJVC2HOQQ3B8GV5h+5
XIqVAYqW7cUWiFeIrGFPLg7xzQs743dWEOcwqiUWST1ltD+SphMT+SGcwQpdtz/SUbp4uS624lpr
YaeatXBPnS+De/uK79MgAJhRnllOlT/wnnVrQMxx6JRFgZJUkUzVUnhXj9qupxbSmIDV1O9tOojX
trB1rLHbwMU1lzpbascCdNcT5OP7ZjkPdFc4LGWVhLaHSi4AqI3GEW/afwtTG8ZQDp+ZrvXYTdOy
KQ+1jg8AaUOdGIHCR0UM50QHJkF5l9fcVYkDkcV1QfslQt9rvrw4ky9oyeSf2C3HNdGPC0ETx7Jv
mER18kAHGEn35V/aYRyFZK0nQgGTjXvw2tNQ0Caj7mmPCCWAraH56Y8gPR+hLSl0JcnyeOG1UIS7
HNR4qKpynExV/pBb1FQZIwp6PB1Ty3sfrYDLosmXvzyw03zQBLEOb0j4Jy8BlUByacql37MRHMXK
P6Gfkf1KAXHtZNdX7KUH+RG6SI+/Vb/4RUhLpXkke4VSfry4DM39+h6k/FdmU/NPOeAsB/ZQTSRL
01ebv2NZDDHgYvfRwnyttlZJP5tpLaireGmC7W91FQ2QJvnKeGpNN7kSyelZpijw9ApKWH/l7vlL
4g+5chlmApfCM3ayWKI171WjZzAz+gwhK1Tqzx2dMS3uSEPYzZAlCruR97q02Ue+1jkxPdrR3iTy
gUqyJQ+GKncDWpKOoDEKNSpuTAoDHeGoOkAypdseiu2foJCkrPV6pvIG5QIiOKyYQ8O5+fZSzuZF
72rFj7cjSeSkx2LPB6hEOS/I2BZbcQutdY0lNmUmEOlMAo1+4Gt4iUkEK4u+Zc8v+nXWbKrE0+0g
9dJIuRvODcpgT9VQTkpncsTj9KtnQmihdS46ZiU/j+c5gIfkHPwac1C7rDhK/JiNEDz9/2kSa6Iq
144UBXijaJSFbV6HvUEoa4HcbohVs9/rkY9pWkFCyl5O95TWASqeYSI4JCfskR3gpgukzo+aFBk9
sYqfNl30JAJvVapMKmE4OtTIH8pDdKbKLefjmnkPRMxsPc/N1F7EHEcbDpUjCu4uq5nPjOz04ffl
w5s5U2DbavWulef/AvPIsbaJ8d1kVoJxR6xuQJAZlS9XgecNqy/rQwpYRo9AQsDY6VnWMVKXAFgZ
eZtXMsKbCBIel6v6Qqt3+QQ/4Sgd4Nk82UJL1jymP5vYx1a2E+IMvMVBO3DK5M9RsCiw6n7gWk2p
1K0f7GTjKGeexK/T/13PxPIrbYrdC+FwNKzOWfcLOy1AbZqEDw82ejcjVdMO/W5XZfxag2UiNI5E
C3zELBIPnUHS/C/lzaHuECQ50D8Q9uw5p7MHbNjfsRcyIxwZU/dbwdGlvsLzA6/PILfo/lbJ2SyE
7ep/wH1C+SnbV428ES9LoV0AG4juemzgI3Epwsqe42fs9gZZElaRLMU85jLpm9d5mMOlGo6bj63e
dS3ab9QUhGbfHM4EpCeEWWKShiovgLFt1ZWMqvepoFV6iKFYXkXdutdq3nfgAP7j7iQxFsp9alOd
R3OHbJ6OMrC+rsp//fCQJNySEENGsZU7nY51K0lSm+2aM179ANaOhFMRGeapMo1pRN/R26I54ex/
ATixLDsf6EhhlwOJh2aJEOAGREfBWsTebf14c4LT/DOpxrQJ47L4DI2R/buv3u+CohSWUR4ridgA
h3/6S9onjvdK3jYCav6sR3zjr0lHLRVygC+1z0gKB8luh6LD7bS8tcM/fG2yCb05Kkd6KbrOyowa
yRpupR0VyFPs3KQz/9KD7pc1xvy81AIfmr71WlWuCDEBv3vK+MnrgbzBSqA9FxAlLiiHk5IBWMQ8
i2S9HOKB3gEcL3cOXE9U4Z3tmxP0vVk+QtxA9JFwkNDnQAg8A2sJsDwjZvqJBBseM0HJ/hopE6jU
IENDPvO9tFhiJBVqLSXATjNfNA3IuzpOwzRlJhR6vZ2AHnwq9KvUHmHRLoqhmKKfan7wPUhvDm9l
aZVr0K8DhYcbflmHRsOEWGfuKRJ0Tyh7mHv6+a31yg4ymGZKkEFfRWjjt9pKd0GmBp6vVe39Taby
SQhXTl/JTWHSP7cpbqNTls5h2IoxuTqflIs8qVrEmdqeuIRyZx16LAndbAfo9F6w4DB6kFxXn5C/
lE0CGidfQyOOwnpG3BZ5jKwNrthYurFwi4kTsnJb9qGIWRdwp+DhTj1SU6ih1+HviXThk45XjJEo
qDtwEX4CMlJt3qa1MhNXPW5xRjehfDcZz8FmTBeAJWdsKOBSKqjUZCni9Eq/9gVYWvvORXakrEvV
Iia9UJa7VtjRUbCsfpt/GTxpc/TQoOR0dAd42zMEVX/MPLnOOmcr0dJfNP1Kr17UXfpE34bZcKuk
bw2tR9PNLZ48NldIxKNNi82V5mmrbDBRCH5h+7O5dD//8ULBYezjd2oj/fAt0JL5qKrOdslRaZTk
9Mcm3WuqcSWGbRuIolPDcqWxF+AyrSWHbFX7DTQgWzf4sKJXfrnwkUqI/1BWvvGCK9W2ME8Z0YCR
5D7INijkb1HyRUPkVRNpn9sy1aip6XdHtejXBb4KQ/WiQnY0nxMueEJz1A/d611foqyJ39TQUUXp
k3vpsw0YXoVubjFABlHc+XATEjyalsi+GTjZBVc73vQu5Tam7hgHWE8+P1onHcGVD2hlCdtx9AUf
t7JiXvZcnGawKXVXzZ1HpM4RbL/8Nn3nowSfROdOFVfyj0wOzl4XfYuWhnO/iVo+Iluc82R8Emh/
KYzMyVvI68VeKOd13cKoF6qRdHGBFWu+vD5qxTyIwd0BSm20+LnXIUmO8UlziFiyggXV1oHiS6HW
AKjXxmNRtACovLwjqZoR5fKGkrKCzQy449a71UmfEamPCjfHAvc91AqSpkolllhSXqYjchSQmBvA
CPN9Cy/CfuTq6jliL+V3qcehySiz7gpJQH2WFeDSWB9xtdjxCxx6sLqFRktdn1xupiSz6atsV/ZU
Isv51btAWt5fylm1PaO5AMxyRKoPvnE7YCnjYWT9gazR7VymX5WgTDCe8UALMe3V4OpEKtL8W2OT
GGWcDbRvNUVKJg/2ahujCd8nZCGiWvCBEt4WHBfJrulv/0U1hzba3njCaXrwcjwrQVJhVpTPYskP
MlT1EM8np8NhhAOa07hivHNVV8SGUdd7cVtRW/GghXwputSqbrpfHm3Jv7dM6VHCYRZ/IaJcsZp5
ESMQ1RI5d822OIc3AhW66DFqWHq+V7mkfcfIXErOdlpDnxZ3NAta+0+pOG2OCwWnGThp0Zwymltj
T5OdHsZvk/CPONwsrYFmiEK3E/US1rad2d/Rwehh6wROUmvENsdRWM6wtzy3OC1OH5049mb0AyOf
2MBcuCcbre9AZCdxiebp27Msj2RuQOkXBFGRHMIqUEnantsMNhbzN87ePCGMrrbQWze7Xstf9fd1
UW2r1vnsKzRksCVvD0ev1k4lV8vd+WsGuK8rIPfyi1f+7MrEUcn1aDac4dd9JX7LdridAiHcj4xR
YzzXg6BdMwcnrQRd1RYLM9QDqK793qFrdnhEluv4Bc7/po0+nhdR6zwe1J9Q2bbm5QNDWiXqkwhx
+xSo8NiM1Vbhlm8MCyJ8Vzuvgk8dsA7X0BOtrshIm3gIoYiExc1oYF7tlyswDHOEw522n3pxcE3i
fIggGiPTZtDMLIJkCXo8ThfIpkgUFJ/RQgqYKZgZ4JV7bDFMwHpQrVDEkMkr681BxKXnhJM8QTdK
4p3qKfYPh3p5K5Dp/oV06zJFkufXS9uHLOFsn2/R90l1E6IgocPuGm5YRo577gGmFAuxp/sgchNN
0G4mC5eAZD0LnJEieVuhX6FBcv8YlN3s32guSrjFs5aGSNM/zwYMsL7l1w/KW9Q1eZt5HYv2+qgI
6ntOhUz/qGQ1DS9DS0GpD0J+NV3hly8IYQKIqccVrnsmBLtjcql8wkwdQSR9G9IwPW87HKYeZ/HU
d0WB7/gl7LrqmrH9cyAUrTDx9ACwXoZdwHqFcibGwGfcT8HJPJ38JeIE5rqo+WKBO79pXfS7J3By
9cK4IKhlZ2eQIbVzQonjZQc3FGplj/h9Mk/3cqilVQIYzTrgCl18S6yNfDaASXHdYrOG4pWvN+W0
3kTh/M3wAWkq6/wgMCH/dNJx5MR+Aaha/6wYS3Mz5BqFZkp/SeRT4vHb1nlNUg3f60U2YrYd81Fg
MABvNUsWjuQ7UyQTpTf4A3ZTN6wrADylmtSm01YxS8NEKrNG2F+jCofvzuxLjDUIA6UhTDg3zdjz
1IBoHCFIIcTlPPDQWrkAquMxriXwnMMaWKtKOWeqH8CGlvAp0rYX/P3Wg73OZtrhLBjX+t8WUvn+
1Vc8hafrjKTee6AAWsgey/JDgCe3jlL6ZphorfquSvmoADSiyffY5TxrqohjROrcR8MOPupKbf+H
OGTewgVdXGb8VYDyJE0mkD3T3Wv6w3fYB9yUZW9f8G4pt7tIsurfeibgGfeJ4n3HHPR9vX+VkzJ4
TqRZMGQIhPU5gPl7Tp3yyJ2v0XgoGVD5SvJ1LTos1VIha6GdD2lDTQWGxL7UWbRNsqCtCJToM/Dn
jVzx7+VxMqQVt865ztWhiwvRbCoQSerAqICJQyv/LGcBpFVc2Cxz0y10+iVcIf1DeVRlJjM1gc7Q
QT8FJqSiQn6vLuY2JLHgYBsF+AF8LwBLsxfXaQASeN/np/C+bD8evQpG45HULynjb4rlz6UpLUFb
ftfMSSM5ViUrFCncQKm5Twg3RMcrdfVfyK4UZiZTV2zaOISHKrHb+LymYwyUG1Zcrg+Dbmv9RmZ7
otyyMS41GLJLYAvtELi1ad+rj2EqDv/WRFLUpsgUkf6aYzcLrWxweL+HtQQO23QTfSQaVqxmXRvL
2adfs8xjU53YHOJk7pf6+MaB9KGjAwYLVo4d+nnSh05ucfIQmZ2IsEhpG9guEcnvpuLn5BeSTzWx
NSjNrn6qAMQy/rntnIdB/ikFNULKnrtFabSQrEX+1/k1u3Z+c1eTyXwEufCCKJAumHOs1so7IS5J
fVU8K9iHrFnS9epk/3LD5k0GIBF2qWm9+7CLA/3vOKaGUSOangsEWxXer+u48PnQan96DzIvVh29
xqhs33pJWJn8bwvqX9aCYp/jRkuNtfiGRNnJHuVLaL+lUvV6PYwTQx+vAo0+RIuNA8zNv0YFzvkG
misTmfP0U8pPwvKGHfZmbuTcrSqlEj7yWvX85qFl3XzV/mX7rqpeapL9OMi30gI2dRmhAUJHY+Cz
hwqLsglavoEA0fSqbFFu/DFP0jiiy9E2XWBeiTLyWKyWRV6fG5lIPwdhAEWpsjbRarG5SHO0w5ya
x48s2PG100aTMlE1SMzHsJ52PyUKFIIGj22wRruKX5G9fRr5Mb0hqHDOCjo3hQpNcebSQ3+BKb+l
5DMv7aV4WeipK80XsnJExdC/OdSbDgiml/Wp5Y73eXZNYB9lzUu7FfzQiGFOndEtN1InyARXUVC8
chY2gGpTCrhdpUFy9zK29an8Vvke3h0+h3DSBhrQ3PwSbU+yULp6I5FIPYqxkw2tvA9XcflOKFPg
3sqGcpwRdi9mLxVFzWOlmZPzqMoiy8OsaZ3C9xaXfZLxUSoPS9iH6qMlNuLQOBFeWlM1dgpXENYe
YfbS09ZtWcs2BKdubApcu5Qa8qzWSqjbR10ElhQwTey7dGhMiYNak/oidb6qu+Sm7yulRgTmg4wE
jyLxhJa/0sKe8DmstkLB9/W+rLHPpRm5CxtXgzAfrhHQY2NsfpeCYdULY0dUrqpRlUuXSwJ+04Cb
7qrx3IVHff82lTnvRHl+vFbKnDXa+LvZb5atnXnu3M2vHrI+RjYO/6ga+rQvgG2BLLTnfYzJNOOy
vI+q9DMfeQrk5FjYQ/nWGvv+XeAA2gRObMIQwkWgSNBJLkCdCMQjGL/WychaIkBXIhPOdsAVtJW9
LHaWY8VlwnX3EAzNIXPVUG8zKy150/pnBoKMhmxZFUxizRBT/M269C36ulY8fhuLOZAfgQ3CyAnJ
xSlucPGG9arkmIhWA+56a6fL1LtIMqjY5WwrAbDX6EI+MggR+OBO74bD7VkwgD5Jv92osKYVtYOt
xmYNXoZlBAHJ5ariWSwMOjeD8KL6EmmYWYglOEJL1z+BtB7aLDdZ4pSj+xJ6RYHJiALxAqe6CXxe
Qbf1981JZhHsgvFlB+xHgrObdENZCS6qSkrY8zStKPlXlo5ZrY8e2o0XiiCAfxFNZKxTG+ijwqqv
7F4tc4UXPtu2SzlkAPYJoXev3ICOYZHN+3CPraYj3wN0pKh3OoX+1ss5Ve29cXZ0vC1xrlxDKve3
z3R5vfoRseWfcRP8J1G5SN4K6XrD8A/AaDNdTPW9ozVwCdigTunsvLb/lGXNHvIoGiyabWH4Jb8v
idUET5euFwcF2+NSw3jaeJkDdHrz9Bme6qB7+5k33sG9J62M0/S1GQU+XHLYWV/ixILyKTapKm+m
DnbbAQM5Ql65RfUYlh4nKgEFKlYaiR7GqqhzDakk3FA/OrL7Nm912JGtjbIIccwTY+K+fAjmWKSa
xLRaPBrw/phH8U0VcpbYory/twAP37XvWOq10OqX0hELiqRMlQakY2q1xBe3MsKM3ETonllVRd86
+DYWHv5FTZwjno/yooo7Z/13y1gTYkp//2cukTYyuPLBxFnPTL5oruHeiU3CCC7xWVpq+koOKHVg
AgNU+CibIAkzlX6yZU/i79EgYa1P5TLS7QbOL9owlzlkLMLyNz3vEJUrfD9iXJ/MwssXMvKGjzOR
P/R4ToAEanrvbrhay5HcVB1iIJhzHEg77e8vePkwRaWj924aXTWhSeIjBdsixy/2r1WdNPuTaGxJ
U7kbi2rxBg+gcjvQu8vdMt/VEq3jnHQkyWbyc8ldelI8jZ/YwBISWFK0cUUe9ui4jybj6AFFRf/5
X8qRitpATc4QXY2hNjreiJgSHuurWhjx2thTRl8DL7vk5prOjARO5s5JYJ2D4zC0tWmobPMc9GCI
alheHaa/3gLKZJm1zPZVcSddTC+OlIK82KXpD6V+O3Uk3hvX1GRg0b7dd6YV0eg938F+w3LanZZb
OUtNIAUK3fLLJmtQ+llmzmQeWLCsIXArvEDr1rb6GDsOsSimsLmT7BDPnu1nL8gKWn1aZG66ic8d
eb6LBD0/6Xl+39aET7kTqw8XdgiqM+ljtRWGRV2b1WDIvSHrDxvrZZYZVPWt6yk4CMXo6rpCwQW8
iA8FX4YubpTrpzcPnY6BB2JT1x8LjdWwAre+R0/WB7qapeCK3nFZ20WdeHXFa+SDadBtmacOqPBg
Vb3I728y3rMKuemauY1E95BOLDDmICsRKT9lLLXHjbkt6VZi8yACgbU27RyXDf43F7I7zRQ4LiEi
Q/rPZ1JklWkVoXLicVp5chDCQIpQu8VAv4SW4CLpaj/InUjfMOGd580tTSCTWGo8J+a6A6sKxvJJ
cBoJG1IMaw+/fXzQnsam2eau2RtNEOGIWj5q1W+983r3IqrgkinxwZV7WRHjQjWzKlWxNPq/wdhR
KLIJda3KAYIrLBuhKs9q/FRlI1fZk0oTS/J7dBnFU9DXkPKKcyofXIkeBMcGQuAVliqFiK214cdN
D/gu0ebJ8hq7YQFZsFyoFm3DYp53bPFAwU3FadUGAnZnO/jv/gs0xUURVFbc/aq0MvyixesBcneM
BZYra9nojuoB/IYd5n9TFHZbFBuCeatKtKJxGMBYfFdCzVcuW1Uiix9aEeGLIKbrYpG7j1WuacJB
uKKIhEF9ho/G8dODAHQMS19YmzuablZ4CsG5hOGap2Rxf5Jusp7+XYqe9V+6XkYlapwXaUIsMIjw
o1llCbMwTyZCc+JeXwFtRStCYQYySf913NSKtjl4u4pYBdTB5d0msZCDL6ho29S7W+N6iOMimHu5
tqHnppuYcxTsvpuUuGRQO5rCUFJXL4tGpUe3khARIcKs9Q90J+55ZAdiLlsOuO1j9L5hEdVvHBQp
0GIhlJpz1V07iBV4zwRXQ5KPwb3PS1kcZM+EPFcQxwh6/e5LGpfD59LekvdIX5fjZG5+AwH38ysm
QqzRZ/k/1iFbBMtyleC9QCgIvk8+6vPIrTPuFI64s9Rv26e4+XTS8f92JcWmd1g/0oqYC1hzTwE3
P9cJ+5ZcVnaS6DNK0tPCjWPa5kpYlHdSal4po3UfhDgVzfgiDhklII9dbnsUuW3X4UhU7a6DIRxa
gGWMe6nEMWN3MpF1aIRd/37lfGq9xANZdHMlOCT+F0p9QjjD2zu2kEXXnlXxjKmtniB0YO+wlUFw
/MB/z3zUonni4dkn9m454hLX0EcE8MVq1rMeiyDVB1l1YAw/FBPMi+n3veMmDKcqgRa8vcEW3JoI
vj8Fq2w8jRzGMr9HTILQa2h4VXTHta+GRyjHVC1qQ43YfG+/g2taeW1Td+K5JymAPeNERUVgFP+e
ay5NdRHIcQrm/C+5IXEXQHeiyIXxqnsT4gKzqfX0FhcmlktlOcJeM/2uU8xiFsQrImNeKo8r4BX4
i6cHg53cwgeVxdF+hI9gHfJAsfkLeK/OeMvEVRENPyGYLR6c6tjRqevfcslOxtFKsHIEacE3g4HK
35bYLVszF+G/OGXe9S8bPnPqTzwbxxP+6Fkg/ALWaLPdQ797oDRzOa37FBSFfnFWXHoqK2BSbM0C
WZEbSbQ6IRqiNYhyp47y6SYrP4on/PNNxy+t4pq7mdXF2liyEUmOmrc4wm8r5KnqVXO1iBOZcITf
4UgPHFwEqu0w16WgMfRkGodLoyYs/vhBEji/Imz9SetFP14Q2afFx2V9bFxh+tQJSghjJ9rEujeh
hz76mH9CSIbzl9nNqL3tE8sowS2FXMf+q3dgiS0yiTMhqbhOCxlKrg2/V2guH/qnFUemhPhwvGp/
5eZtuttD8R6WoSRiAqq/ybDr3UnTFN0QZX/KeZKpqvFLHcvrrsLGcaKuvQFQUqKr2bhAQ8u23wAh
0JifbnvXQ5zGorO6bPQzgggIjsdF8z+JtDHZGWSheWK02tnKn6EpXmjuVbE/ceMtrpI+ZxnnJwA7
cgFeeS0mqRWkWMmAe8TaoCRBdmK5eZK1sIyIOYjuPKmv0rvCVL5ak+Pupy7UGW1HhivJJZnFCiwK
2IhAchtXosuqYNx00OmAQO3eP0SU/G7E6gCNMIeQc42OikkdXQbKd+AUI1XAhHydpi+EY1BxjvHX
QlXPS1T7Z+4zVGPdAbfmb2MySAabc0UyibY7j6VbwhV3h1Q4f+m9+EZ1vn8561SfemOUT2aDwh6i
k2nJPkLLMsHWMp3PB17IDooBSn0MgixLjxs4iNwgHIx/Gl0Vy7Od8HrdD4zvefoPF269ZuvDujtA
qbBkhZxtS4CLPx1pmIMpotymT0yKza32gpj546/H5WcNMJA14VSUonpX6SnI8aPaICcH18298Dbq
ITdDmZnWOtvzvH+wMDmzbD91y5zKNDQBTH1WaeUDZmzxeMraY9gQ0gQKCrCXLTM4fg+yy35y76fC
PshmlqLImw5dEoiVq31qELi7fimWBfXoAA0sVXUtp+N7XboLWN1doG9CMfHCbnnYJKZuzdeZlKV2
nZemsZ9Nsc5JICOI1JuYvo11Wf2I5VbRV5JmJhsrAzq/Xx0hdOdxyrOsgbK8rfK7JMqTCkxwPCxn
p6AH5ezPa4IzMdVuSUtfqvOR/yIRhMa/zeiNyOtzY8lnpYswxSDs7roTxWbyVoliVfvxPjfcna94
1L/AZv3+41siYr6zJiugruC9CmhpeLwEBfwejdemcdk1mx7rKPXR76uZEbExVv3XTa28txFvHF7R
Lr1Gp96o7peAwiyNoCPCxPAuIYlL2rrOzHtomNn8pcOX1D1QidqsgPFk/vRx+N9MX5Q9OHb0iemV
kcjxACbgHPsoacYQrovPhzUEWZ3qcFYeZPV6jqknKvZSgr+UjHWMneKcB0T/23dgj0y3J9FfURRM
wP3FRGPNRt7GwX9q2JfchByD9cCa1clGcxg4Ddf7gA7LS796Mex9DFLhP5ldB2pKMMy5wlVHeJA9
ZBoQh1aBD9BvTjkye+LBw3+CIjKtKNlTyyFB/e8ScngonR2nJ/UQYT8UcLMxRAgbJoillk43UJ9F
gX5hFsJpvCTLG34h+2qfdt7ImFe+gQlNuDZ2Uh9WN9maP2sHn/dnCsG02Jn7jWbCVM2bwh+XTepz
3UAcfGl5dUdtF/C5Owc4fzW0UCIf1Qpb3xWVFkB38JMHs2hM8z0tCUC/ocN61qHneg1MuCV/KgVb
4150EE7RHAt+OmNIdTB2ERWeMwZo4H7xekly6ZtP8dfhkCPICwdK9TZsZZARDRX3t+XBnA6Xf1io
dIEBHd6hWXsJKT3vzIAj3xMLFxt9JOV9HxHa8/pwdDvaEHssb/B/ZKwA/KzzJeMF7YBezc82SOs7
Ud1AzsJDw7UjRIklKeW6tImstqM4J18jNzaY80QdNqvNJuatinkXs9eOH4CH3HuroAPXUrZWv23b
c0fl8qxFnMmTIvuK4dWngVQdzjqkP9jzl1CHB7Jb/DoqeCoVyvZB71WxzVNE2B9NRi6KRMgxwR42
Vt/C0g5c78Pa+qoItlpgsjIHpLH8HalufAEitfQ7QPG7lchg8SixQLdnMZPef8NMzta5/QA/2rS8
OQWKKa3q4+AMb4AHZNJx7XZTul3rY4gMr497rgfgmFrK9ULA1k1PR2KN+DmFgeJqNhmL34Zfn0jU
YxR1+Q73s2foV0toR1AGhY48RtX/tz7adXrTRnfJJy+5rwUG+EPR8zHJJ2ODW1TikbzHL5PbUksI
/aBfzl6pY3mQjU4afL6hKQUlON8WMgjty30d4YwYrZEZFGunp646e103XRYIhyEP3Rzhv5vcDjhx
tGeQFHcLMkDWjkKT8+3njP4AMDsB6SzfFk/fymFS8WBBTyH6clnoAx2G7plV24JuyM9HY4DHLBKg
yBC2hglK1cFpd2CUQymYkVvzIqja7Ztxlqe5SdguTgd0k9t4Lnv87nYy3qnnSn6jSJoMUfiyE8+t
9jjG+9OdxSeoRoMeqzHAzyWxpq3or3BzKpD7Ca/bS90QfKiJTvdrjCJdQb/6hWayu7PHGrpVIcn2
EW2qgJ78GXcJrMZCd7dpU5fQKwa4Fa4SXYjJjGd/fAHxP+5Cn2TTX1QzCrTxCB8/KCckG4+Q8zHX
bnWzyqEeJvQIA2kmrjqPwZBMLeLrpKs7Jt9RgzjbkrIPORSonZLq4M1hXK27RNQZuCOX2tsbm4Ty
UiXBTwOjp3NYbuBOCnIIybz5hU8ZGGUx5U0IGrYbN04Aafh2cFDHOdgaQd1a2MvBkQZhGHjC757g
ZCmUW8SE8qmNhPjtPqHX1+7er5dWdWo8Oo/5NZyo9ErrzYxkKOPsB7tMGFiuhDLZHubsFq0gwqGT
66CIYB5vKF+Qcn8RHYfk8E2FREOGUwF6cLMJX5CsXYPshLzUNMabBUWBRQip0BE6n2STubIQe6Pm
+BG+KUFNZ2r1ym2d4IZKfsZ74cqLq7Cl+Irna00G0OhaAi/hgSe5y65b4dGAnXU77JrzruT4U+RY
RywtGsZ3JutmO8bGpONfk3TQyyhIB9Udx7yqJCKhmDqfckiS7dWAWZNCC2DGURNZVzNd1MrzzVxW
1uEnOSfFnzEoGXzWjk0N797MLMrqYzSSd9tM/4wwRcrh/2EyxEwsbfklLRzGEcXgTT38RAvCwQ/Z
ytUwgF2OAkEq0G8O50H/m7Z7htEuJ26UcOCK/P4lOGO9YHzTzXPvYpYfRatwGzngQfLDQo7DTpCL
8Zo4b1VmE7Z2R11532xNbBSTtshM5E0DIdVu+odUkswD/hKN/4nM/n/KPzdLTe3nSe92jRHWsIJy
vpE6Lb+8/W4UZAS4ROK9iztvXRcc8XYJUXoFo6FIacugF4eKi9+2vczhbxFaGjiTdSg5wZIiI34h
+jZ2PePlbupT67dlg1D0voq8YweH+n5gsmG3oVHWe0XnyJwTCPqF/5jc+taZSqsTmJ/vQhkzhTm5
x3iAbEDeDF8/E2rr+6WkqZnYhUKundorgdTa1GGQxteATF+qfW1XCmIAnsRRKlkIaBEo2jPbb9D6
M6K4cilr1JrZCorbGuFf7DpwFCPuRzVqqIN9HY9R4zOKoN+EBthyI5Qvu727ctrzQc/2mRedsYet
C3hRcyv7G30SiZax+C+k+byvycxZCTyGbhqZUApgP0W6LkPqMMd1NxkS42lQyLQ06aAtExFZ8FLW
NNbh5D5s0Cay3qbD3BJyR3oyX3+Vo4AOCUI4mWa8fQbJaKGx4QX14PsZhei7B/iwbDBwDvhDP6hg
7JvzUs4HRrGlezJk3lT2x4sVRZYkYmAtazTvzhZ4RrZkdblq4MqXgSWhApBt6iWF3a6mQwRB4U9W
etdq94a6+dwiHHqcfqciodQM2v3E6uPK5SWhVzIw8lX/Qd0bcs9ZsDnICoarce8rg6JfwYZObuV3
F28sDAeMWi1uzU2GCJBddjAGnAwVdPRKkL7BbnuPuIy4LhmZCr9agmAHCXYrxEXlm4L6/JxyKS+3
DMUcg38MMBGRRGQ7aM/pomcV1213vMm1PcJPWyLN/IQYfj9ry5+9jIjIjrATvZ8BZ9+nxNfYbPWk
3u3ZtcF+0hD7Uu1v4Hn/a6jKCbjVimeAyonI1stwEVCkL66IzTjUpyd9/ifAzPalVeien9ZLLRVR
yPhzGU0y/mHi86hML+kL9gfLl/HBPrTHxUponpjfTLrHpCQ+gSseLBHSVSm88PZjBk3uJXvzahjZ
CR8Gi0N/C3rE2I6HmFftAiqKm16nrY71sIleF5CPP65fCJJo4ox72YrJg6YxFxUdkjH862pg+fUO
Dmrn1FuejuPmtLyi1LRX4ow+ryrpjXD41X40MCOKhD91FBUsoCk4O+GMenXEFtED+Zg7ZIFOUgPR
2YQW6q/BNOFJeZc0y3TEu4AavvD+K6PpYN9d2I9yzfuYj9VLAkWWd0KzLy2miR7SO2Boi736Gp+s
ORDrzlkPohEU3gPzhZR5lF13uu6KRhjq6eVpe9vX3GcttK4RcdRXOTVRVyH+avC0rbYop6ezz8Hy
1XLBIo6fzaR820pcG4oUyKEktVwTggx+1FgZDywhFV4MvzcJFysFSEFUGQ4f/2o1YSXa99YzqiTf
G2YfjNiRMNQQWfBkM4lUELjBv38iA1HKuSeurvf+YKiNVKrMmOTBGDs0bzQMngU/m5OM5cpTVG9+
6zqXLClWseS6RAzCqwvES3FMn75h9jz9AP/HpfqkTiUp2xtxZ2nk/V3D+tkCbSF/dM7hYOkhN2Qg
GDcL2GZ9cFfYaK/8PKYbbBma1Cnt00f1zIvRdujiq0p+hllVJaRraSlF0Qy59LoNmC3Hdz9SdqAl
Q8vDNTqM0COIgPSMNqqvYpvJPnLm3009T+c3uQNiP0TQYp0/SSAjFWfH1oGYhhGmFY6yfRfVglYH
yebiYCi8PkA4JfF3qFVjHvga7MY2m/bvxxkryvHvb1E+wz/Iw5A7XvgX0NZbHYf2psQDSkEJ225+
ZPubUo91oqbFrPNiV0LypuldeZ/+iRFZedd+rOQ+NjM8K477AcTVVDh75KmH5jrTxz66LGRE+d4Z
76K22/7xQvas4Ziy64mblftoD3QjwTCZJvnkAJIUaRLJHklXvKO0OPVUkxZGC6HoBYKI3/n0rwEq
HCzs47ciyhRWkMVXBbfkVpYlgvf+BpzNhMTxybQSyG3IYGsFyFbsYOjo3hwc04eznwk5bfbzaWk2
bjFdJqhH/59Xylv5Km8cfQPKItS1APvcaTeKaZ19117C/5TtIUSFF7x7ABVNr2F8hhqR2oixOCha
lOuL355N3Yf7xmOhCBFr2mXGn7dE4rDfcd9p7pfSUWDBepmxPjfl3r9XRIOCAxq1tVgtZKjSRq3k
imLTQVA1XxS8iTJeGUe3/lm//5xEZi61zXuWT6xO1RFWqEDU8itbLVe6o4EAKrGRgFp4go3hqm0y
gaKkWgG/2wecQdL9Wu9z598ft7wpxMWL6kqVkCGt1rBxUBekzfU4UeF8+VGML++WwMLNRBYtrNYJ
nax88XeNpjOxrpOt5AkRrmipV6J9knliySOh0a6M5dQgj7Ut6ejqYoPuhcxZANbhCkg8KyT2UC1y
VuWlZ1c8rJ5SWHObFbE8qsIaqNlVGpJhccChE6yHCLYnwmzzhkACdxPyAJJAWYniOw8W/csWY3AH
jPUfgaBW1rukJa3VAVLOm0H4KsEuwiC+mRmmOydQX3dIF6H5lbKQ77SWVuWv87fLw4h1djTLiJQT
O2pwdjjyOicD8ruwF8pIIyt/7UN+ZbCo7HCuho53eNmereZKODz3tLMl8AnBn4WkIlpCISq1XSPu
ob72XFMchRTTKkzBz0WKowgZmTK9jBedEH1/jpm8Amx6FOG8NfQ1bquvXll3WDwmbaG9HsjhKz4i
7J9TH4L2uSFnpNkDQTzjXLaSGeU3zR+hyFfxVm42EwllLTer3iG0+cDVuxwFasU+BArR2k3FBl1a
YIkDimLCpx/1P/bUZyDKPLtJ3a5HzjBx0CkF2xrOJMVgJVnNrbq/srwcbgb7IujsJx1PvcxOEfKk
P0flFJxYyRq0dZYjLvxtU/YMii/1ynx5AVBc5aDB6u11XJq7nQybikpje9D8Pk95ImS7XZUPbKGs
rpalinXaeoepi/nSXJJWIoEQSYD5BXW7aCNASqIgy+vsdubu8ej0fz0Tozh9USkoX3ZOmB01eFOw
FSg+QFWkzGtMeGF/OCfP8OhHDlAgEZUhkr3FAgifQabb73WMr1RaKPDijZbX6ln//aM0Ei4ub8QN
7vxxo98gYL2hRGzzjWL6jKHPCtp4RBamskS7rpl55k3XzF48jvcktTAcZcq9WHSRMP9L6e6MMn5Z
4cMK0jdL8EjR4R6Z1BtH1/zBuGTEUydBfY3HL9xus6t5QOoMuReXKfOerfu/j+4olPPLEokn3aZ7
g+VB3aJqPZZKQspV1sjB1qiPdJNLsgqdta/at6WnHPo96v3DNOzdEImXt6gNjpnqyiTH8FcYvppX
SIK9bU3Xx6RR+YmlG2z5+vKNsocvRLYJMGQ/osJ5U8wiV4TmFgfWYvDd4nY0i4Gh/YJKB+UyRD2s
FFtwcPgM22Mh5c7JRUBUdo8e57e95sTa/E96CaMSiO270AEL8N9x+jtH4M31ogjnhX+kj5zUrkzw
4qOlrsavpLHFTQopL3F7I3kxn8lIzWSjEVYc6+aOzv61TM3mBXWzpV0MbGDQJypJNKkZ+v+RqjZT
IjWVecqeTykLAF8f1GOjnxYUBqZ3I22DXMFG1g3Pgx8y4kLXKHjYbiBvE8XGv+iAOUVTfHqDkoRe
EEVZCSEXC3Wd9kmtpbT0LZd7xOzQ3aI/bjIyOwDN7KXsXZXq1RAXjAoWXot8uKDA3wG5jvnH9kFv
Vki6sFVC7NrlqzJgJSWyDamYraCdoyXXSlKvFwhBM4sCgLxi0hQ44oJPbSHHKdau4FZCKUZQMcWk
Yz3Hh5K0+cfU3UhbfGs/evG+RxUuGLUzWFyBGb6j/RqlZzxMOF5JB7AU6PLEntfv8WLMTXn39ux/
1tULs5c/bYw9LvIcipP1QAkTD1Vx8h9HBdkuUSWFqR3eMKLDRfljywtw02pxg6OYXpKDuc8oc73N
XZ6ojQvTxDT5feIldqT2TTNoJcCSzdKhYw2A/9z5s551mHkYNwRChm8XqbKLIKpPkxEMiFs106kO
JCUuIZeasGCk60MtuZHUbg1lOLA8tOVh03bp07SyTutCLwS6sP+GAvl0ykBiCI9sp5wKBF2R2Fez
fkGodcwzdDcSfbO5IfqjEELrLcJTAQlmn9pL+roiGqFOkEhFhfOSVS99DYYc/W2R1AimAGFOTL4P
c20JNK4PN1VkWPbHXwkj59rDb9ZqGQGt3HoPMh2xnmi7fg+7WW611ufCzlDX4LBRjp1VMKtvvqWs
I+ipxOHids4rOfXZ5n80WHqn/hJT3/ujd4j2518+8hX3vQzYx0wXeFzrC9j9ZldwGOLarJue8FT1
HcnINdVfqZsM4yrYL6U/xcbVWaW53pl2EJkqW4p2mK0LbV4IIPkKNHuVJBrS76YNg0O4vUG1kAoD
M8JyaeUBOEw005DOjOwFFaGhVF4fIg0EgTgCwxt/FR9ErQ6B7VDEMHilo8bJT1t5neJMwfyMaCJd
R0oB1p+WBy7ee+nEshXnA4IBOLnI4Fzq+fxy9Fmk+b+AMicTXaPihe0ZvKvtOMZvMhp+ZWLm60e8
Gt8iPg+HVepi7frgkmIJ/PzAhbfDLPt/fLLcRN+llo/egorkIDCg1Bym+EcVYSDM6VrE+lXvTtdm
Z9ieWu5ajIrnxbqemkgYnGQuyFdU61+nr/W5lWzOemxyQMYquaBCseceVbhtbJbdkK4CLiQtaHsA
eRO3RC33asagyJesv7qbScFO4vLcKSq+4NhMIeoBhR7WsWBmdChtCtfLlBESiN/BxC5G1zG7vUhJ
7WeuydcgiDQ4BuUOuPDjR5ciPtCpL957Dcewyav6X0R24Kn8Yro5ZjnClVroIv1wAwtAm5BzLmXv
vEhMgF6d/lMBk1V8E7UiUEQFZMw6SNcuGNkQGMRBqvyhKMW8WxZ0V0v3Kx1Fv8QDsWTNC+k3sOw8
Y8784y5d9g9i2fegwWwmrEva4x+Q4+d1AiaeOfId0CleJVzzY78agQA9ETcmsmYFxo8VZq5oRMCn
+48F46TeQK9ufAqMAEiVobnva8Q6T300KisMfhS3Yy1NJBScqfupsmh61swT4VlIaTZie6xMPh14
inetaHK2SeCarDBgR424quSscrscwUA6X9Ai7tP7Uopbkp+CjAPEtPQrzInYQdOikRZDc69oAIAv
6xvhMD58tBmy77PnMhZIiFDOegUxDtPDsbmVRD3Yxd4A09UqZUNYXcVKvwl6sIm/DsQzQqDgwq1M
8MKFsHS8UtyMX9Srm19GG7cz9RRQx9Q+cwuHyxqYQPSO7GJCbfNbobTHMr3z76mQNMPPtlvBTNuF
MCx05BhDF+Obe9iDoaHo59hiH+82e50fRQFnAEWPYp2FpImZS+buk9iOVyI9kSPZJNWEkzXVcTdA
ssbPSK6CDPgpIRSpxImfgq3BoinV5meZw1izdrvT+PU6EvEp4xq497I1tT9sQybfTsM/UbDgjvOm
c0tEpdael29Xor0O25dNIPWMZGSc9PmQ8PTxmNgA2a28gUaiAiVbvIat7JM+SzMT/pAu20Xnners
eCD/BTZAbYLJjs+jVPfCArN9kqtX6X42YTlQsVMf8F7YofnXv5yIMVVWHeX2gEmoi7tUSfOtdf1O
/JpwwYkS6vmc9Lv1VMPkr+QKiJKZIv/3ti06pS/otsoWOF0sQ4aZSp0RYiMWwfk4sr7Rl2rnFncP
BIrsFTw4+2il2yI5NNbe65qlAdMJO1lTg18bfC2+j0OT6jtttTxxa5I9kbRF4Q8Pbb6Kh7PVnV+e
ZnIF2wyNB0LS7inxyt0TYimMQ548CvbkLW4Rg/0LG2SoQqWIrvzpxlKnr96YTh6efmB618Zvp4C2
xInABqHfaQWISY0YNLhvpLhyRzlV51nPNFkZfWsbF8jkjQPvJFHTIdQdQX2TX/lKpYzSzPeGP7WB
gRuRi3kmDjbJOLTSDrGRpEuz/CK7v7P+k5ktbKzW0xF6wC0bVZ5WfJ1AVGKOX8BHfFe3y0WZE0Ro
yBMaOqk18LV55WsOy163nwofMzm23tq01Q3RHKfBryR0nE8JKPxRPbERKitY12S8db+oDo/lADHs
bHekrDEgJRMz7dyp11qHhd4DV+9crCY9HNTnWOtsdjY/4D313upqzRAI704aBXiV9v8oJVE1u5LP
yp8cCdX1ZfPLGtz83QSiabx5jsu5b72w6Z6MpinxCRhrJ7arhh8XPyfqMLvsIXlNrhx3UPO5NYvK
r39KFahVQ6Eqv4r262GhzBee+krKEnvV2/sELOt+xkkxXwy7CAiOBP6zwKeE6dCJYbFU2LQN4/QY
Yv7hA30n2RlEufTG81FF69nV90xQSmWXCh0zSKCXZd0V5KY+UKE7OQYdr5JtN9+NgbpEl6IEki/C
2zIWBzDpIAodoW/EIP0p8NHfwH8vZWWd+h1BgrQRxege5qqyDzlV4OMeEBf5XY7TvocKx0L3TPK2
zfxBa571XLHX3+Mz9fy/v+Rak+ZJyuZnhyT1apT27Wo4Q5dofqhUVGa/0u0o0iJcq7eEkpJ5U+5N
QPHAnDqplziEZ770Mp5tR7N8Fz3z85MvAUh+k6aYb9EBAa0//vbxEQ1EsEpS6zA42RNK8/Y/LzmI
rVr8JtQy6MadeD9s6GgnT3ZtVKptoi9heCRdKtKsToYdYANsro0pGDxf9tN9MEvO42FT8qTcOxxI
og6sbE5F0+mg1ZX2ul3PqlqqWu+VneFeCjsQOyNdYXoe2ON28gXAfyNrTahURgrg0OcCl8i+lqtI
2xAwTOa8XPYpRclRmhoFHmw0I7i48nTi7K1L68vN8TmD1x/XswzGTz7qIuwu7EJJeOtK2NdknwYb
2Kx+YgW2jJE1LasG19X3J3iUEj8GUCiGAZXIFcbG+tEWBb3XZcusuiwHul/0/0ZUeB3hv7cBs+Ge
WMHkb/QkQi0hJKdRJ5j8zx8itNx1BiC1OIMz9GStB7I+RnuwGNIm96h+D5mGBCv0VN6IG8Y7YvXT
28wW14h5KtdfBKWOklusF3TbSXOyAovWoNayDS+qJUNh+terNt8tCemqQY0+gLyQduRxe/yO6dId
OIC27q+ib3pqCN/mqvX65GCQQkDw7Eh4yEriyN3j7m7CxBI4X36yR2jSZfjmEdp2N3lNHk00iU9r
PlYX8gDP7hnyyyhJ3QeztpfilkKH9J9bs+M+5NEZF2s8lE0HoV18Z3UxpkybPcARPiwAEY/OQ1KX
sptReli8f7SccmqkVCBhLEb1jTY5bZI4q/foFxTBlkzbLd9TRm19PCLRjmXFjE4MO0vtc+g/YStj
pNUu8Uo9V8kQ5Rr18VwJxu7ZeK7YfK4DoQYTL4Brrpe8zTOYpga6lmKV33BH1F2p1Ff6LveH8Vxe
rCo4GFAdg8mggz1vjb5YoKElRI0IA9BReJsElOLEujVKuCD6Nk/lDqEPS4jwCPPO2Oh5JI61OvnA
y2GtHCKygf2p7JAoZmSULNPem7lw62wBVodDVI8HSZhVI9PU8kk8g2IKwNB/tJBvMk5LXZAIp6HA
kFswH4zUJqk1lEZroGuUNaG0RJNyFB88Acp/L5RIZESvzh3JIB1vRhCSAUxRFByhlU15HgXYnbrJ
869BX+AeUdhGCosN7+EMmqLOHlwScXfvK+owLSekhSRUyykkDCfJyohid8iNmKJfxsTCoDfhAgXf
qDx7PHPAU92ih3hQCqDmIDgzokC1MBjdUKcTkydQ2Q+mfP4ez3BlYEeCVI/fFBAGND0IYZ2Pk59P
Ekig3e5fhHooIAycbm6IGzuyvzZwEOXdyaO2IiJQCNdZNTpH6yaA2TJXRHlexZmPi/0A2BRjk5DW
Vv0hkxCVT2i9fbnZlUwJ8MzXWRPMA3A2L4gf0aGWqLqJzz9ZF8dH5PSSpulfa/WtoPQ5l2CR8p+Z
np3K4mCFmlnEyD5rZe3Yv4g3mZS4QueZB6E5RbT+R+5m68QmrV0E4CbABmZ//lqNqBSp08qN0+zh
vnHP/5br8OSMGnmBpaRQRe75kH3NspsvzIW2JBHkeKIzxRTo7m+Hv6bMOWqxppALzqjpbku6/Pry
ONXp7+yZDOS3q6/RfTpVPTYvvMzztiCwgmR6VFHvZLcReFXTFbRX36x/pvX4xq6WBbBj1Wb8YL3a
3gTB3ozEfOOaKiA/xsmPwluIk+0Q1We612nQdLttvdf6hinSieaaS80Bmc0DcTnJMonwd2W+0XEN
+W8+IrzXQMADPYjsTg30W+fddKxe0hRiygYmLkDiVyff7bBqXOC5hh3crEv8dvSUMERvymXzl58A
R0CcrTTXy+wKhSMnTSMDxNfBAXvnW3Cjw5GeLHwaoELn8C5UFA06K9Kx/lF/8bDrjJiPOSpkY+mq
3IqhoDoDGbeJ42WnglemHUzEp7h/RAdRGnwJFviaAMBA+iVZJ5wg/hO5nEICX1bYuCBZvJNouDv3
rOdP80JhFUBkQGQiH4V2Cn3fc3+ECtg9fcN9qM+gYbbVk53Jouu8fRYB3SAcu/g5mwpzOljLPY8T
m1HIISrx0qzMUnHEI59+CHTuag+zD8v8s+WR7fgLv9HXw22V8CHnhPUeF1vZPOJvyb+6pzIbkxrh
82Uk6sl00jof7x+pXX3k5XlvbUzkz7mBUhUtGGoBTBsCNIhApx4cTp3nzBbQqXoRP+xpaOm8GBJZ
l6Y21rNA2+DFS+Z0L/x2kL1s++HrCli8vHYJguMcRg0AXyZMAMz1nLGKJZpixDIxCIyLFcktk0+8
PsAxyYyZsVBBU256N80KM76OPFTCFBe0wh3kO0QK/EZ5pjMoxAVDQYM9IfsD8dhjsa1VYTC7EqU8
a9UUjv10CbO4UMTjuWwqa3MwQ1kvyR4nfpanjbVjbx+8TQcovA8gr6NRsEEyLv5yNdkTRqRSbw59
7XsXRk7L/8EmBAMMi9HFzGhN+f0g1k6a0D9nDeKqeZGQ9k9MZf2fZNu1SSAwrKlZ8zSCp88WtHCB
2c2yP5tbLhFrCVPxOvyN+VeM/oTu2k0Tc1CowUNV385Gp0jwDxL3Z+LIjmCkygKFFFUAPL1+YCoI
BG97edEjabwgfpn7cCBqnfUzkCpmKPSseJNHnbd6tFIbepOB+vxPQrIjdSqUInE53j1ID3UqFGhK
kK4UD7Dc7mLluy/dkt8JH/3gwAQDVUYlf0b8W8+OrNll+vw4DuhFxnEpg0OHCBMMhgFsEtTyzCkh
L+n2zuvtOeP6HUt6wA8VMFbyj9WyoEk5KdWzyDWAF/+SjmqN/bSGOC+V8nb7SrrChZQg4/A24Hzx
cI4bAjSia1R/9fU0MmkBwKbf5yllY3oOSEAdKlDW4XezbvLSnkiOhUWfcSRBrsmt0SNjHHmIvSA7
71sr4B6jkqHYZ6pPnQehoJAEx/xK1ZWXOIhAafm5sQ0cEZRE/CwGPagROilSbDdgb2WY5jsGhqPm
YiXkfmx+cma2JAtTvgGx27Cr3yaQsKwu/bXrSc0Mv3NRRRM/eQ/hhJVrz1TydgBGO3EbqocMbmF0
F0/KDk0KsUIMMj/eQvOIY5bK4gspU2I0TDeV8jZvwLQsqoRACKwhTVVJ0CxJrou0qYTCXrFYFBgy
47eeSRqfXiw0olIiCKWtLHmVLlkljBaz1b0IhYNhjEiRmT/OMY7c4nvajjX71l/2CJExUU648bsf
YWiuPcuyR3D8fngQExqzHPwpsQWMspJD9LV9vc50PlYA31ci54OQB4+RcO/ig8v3PLdDtYjgAGqC
D20LoONnEF1rw6QnSmWSQruG/SAmYc8aGZa+Xexk0DAU4kIJeqodBBbTYT9ASj8nMkJ35kl30zkV
2RisBGJmDUijbCNOZswafwdt7JVvhfXRf53MJFThjRdqQKsrk+N6ERcljGl1ibxcSyyUXeFOQS1+
vAjZxcDQpzFhxP5G6yeaD0IFODdj66RKPdYnO3WOH4YCY/V8IgNZOLi78BtDuHUCvfgzvNBQHptZ
jbxwuRjqGoopv7s5QGowl/2sPrgPefgd1rltZez5oO/NZxxjp+C6jO9OzpbBSRAi13PKOLlNyfzR
BvLGFdH2b65HAEN129CgApD7zs3amz/tiCY+sqfAc0sCveWTGn/tPT8yhANm0xu8R1VxBJFlNloj
ecNg0KA/bWx8PLYn57Loi6ov9n0bfeUKTireF2+nwEWGLN1hIyO6dgVnhT68O0vPLO0iTRU/e9uZ
j0f/MCCZdfe5B8EiDhA5qz7P8u2wBGfmpPTAMkoRzks+PQpH4FTzisdkgeACmd1UKj39GFKHCDTM
C9d9ArEgeQGERdy8anSrBAeSSI6pr0085vBT/qwlNmCV4RLDg2JOG00q3yo1PbuBGELMgvJAykqu
gDJtf8/m8Drj8SyqtFGgHhQKTb0bA+i2kafckijKmfwiYJAUpgkZDE7iB9XiBpT3Rcbc+VTIWEDu
+ZPTPu/tHYCl8pGdKs3ITyKhVwASIlEbSSMytz0HyHgczaqxWe8Tno2OhQB4NavqIjhjvSB4KpmC
q0Dk6FOhCg6tpWMtzTDYSFhDCLBaLe+c6ouT2SxxbuXIq1+9hBceWHfI8Gy/j9yExiNtHfmll9fT
6xrb1a7+DoRMqQBICQgqF70nrOD43hFtCm7afWVL5oxV++qlOoYjhKtbXaxl/J2GUqrf4Vnvdh4a
B7ReMgi3pgqhrtzWfOBdsL01Am4+5RRVkBos/p8Srf6NgbaVIAKr2GHdRDAp6MQ0M5Gj32uEJ3r2
diJ6w97NhLUf8V4j5ZH3FnnCwKRRB3ewn56hMCCXCLl5GX5RWY+01ud0Vey7nzKoRThbFbjrjomU
GcNBFrYAHD+uisy8HZRB0mH+xwvqwxEzb20D8SPQPZ5s7cXpc36lC/cEtSXA0fEGrErfHFnUdWE/
lVKwUu0SeomeHvjmHmaGdUvFWG0mWVRmXuTccwGlmdnVOP/kk4aw+KkCpZAVdKB+hclkxNtPeEM+
2Ym8VfOo/cdg5RFYilJJvNtamS2wfrzZz1KTsxvleH8arL5uu8hvpr9nemOwkHS89hHmPk++1KmP
qXiKvEoVbAD5ZNsqHnSqi2u4T4jK9QpqlzdH3A13kewoJlsc7AQ98A11vt+LkPtbzehLgBm1keUO
2qiDlqXISR8R65i6GXq0AyCigSgjqWQs14ngyupTiIhI+TXG3R7yoiCObgDNMf1nwlhi5LSmy4NQ
MkjDTZP3cAK88N5kN2z65sud8b1UdgwPVD8w15jDxPlwGWNhUkDlKMqpYdGUDPWklaMzyIzbH3hq
60xj3WE8dXkEBceQzXrIC7U7HyjrgBwSP9Kb81ROdwUmD2bTcA4aolU7LgY3wsRXsS3YJeA8ur1i
hwd+CMVwfo2CdRDbJpaiESbq1jIRQ/AnMcxP20Tfmy9wiF4ull7HEUEvQl+QfjVBWaJ5/J4/GdmC
CcqpuP+Es9FdLC/TGyyxwVa+PQFveBpHX6r4ugJvjJUsOhoBylxdJrJPlbhh1bA9MLxnYs9gtWKg
eMoHcL1LnleTsyd0mUORx806IKjQdcxz2MHkDVereo3AUd4GhlA3TlfKWLxTfGPja+z3kIFDt/eY
yrNaoSBS6AlljnYtz8PXnlaaCptHM2VpXRbSk1Xu3A/WM2HjKDyOQBSVHy8Al84frY1KEfoK90Rp
xOeGU1DjYzDcf0hKwS8EIFZwMewmfzKUc8M+ESEm2Phzlx9jFmf9U6/xl1P04JZH9MzIhB/huoCl
f6uhZLAJkzFiyJIcD4xKmcsRthccnVcNI9qk06L+HKBtjI1iM2hOKor0Y6Ua/uQViTYFrKsmxgTb
XhEdO53N1+XCyGQDcYURSFyE1SuF8R72tLzghcfdnWt9Yw1krrD6nvdntL6/U9r6zeQmdRcsJnPy
YwtxMZx2Re44pTUeum6rA/9XQe9EtZ8qAQXGth4Vbco+gTsyRqq+rP9jvOVZS4xLnNhcIkWeISEB
qM3+70NyaFTQ2lJUagSXQiwWmg2OXaSWBMpyI+zZs3YXAZVkvUoBCK/U7FCjTHDnQ6pj6lkfzirt
ihY7QJG+N56Ga5GXP3uXJV5MgmDYOUPkDcKtFbkAw6lMn5tijdhoteV+mZtWhbtJwlmxA5UeSxZ7
QzbuPGjHAawtHsTK3uba9dQjRZqnLbojRhvB1gDzaBVXKaw2l2/PieJKVm3ZyNazN4+b07SVBDnK
ykuoTylM/WfD0v/NAsWxSsBIEgMUmSq+vo26dVfQ+W/DBXJQawJ7lt6fM8Nm5VbZ0pgyS1h/pRxI
Yz5UxadEjyV9V2rPETwILFUDZG9ckKdS8ITXTXfdYXzt60+1XKyCJXDDhafalmpOln5FWyJ1WIEC
EPxHla3WdclKpY1XUCvqLa0LGHSYBQSAGzaquSsNt2b/IcbwJG4N1Dr5/vdKKVlYmC1nNy42JK2G
GjYCf3bOyVGA0ee1f94ugoICt/VMfKDq9OdDS9+1zZJ2Da+Cf1AYHqZlDyJm/5r+nUZd6WTaUP8+
suPqkrI/9ZVItjKWyXz5YfrBd+rB8dWSXkIWlKuclq909AyFooqFAt2PhCkUWX4TKFIUXMsnLfdr
e5Nd1y+sLys+CR6xy9slbZ537lQCQjUPTYyPfRRxeBU1S3afAp5QEu98SSHZvwhiT7gXinCMtnVA
TKizu68BSzLOh7LT/2PcjOQrybiSRxwL2kKDO+WNwwgV6D7cDtIalIMA8gY2gdU7TezFQX1X7pn9
YpUKi5DZP1NCmJUKi6NbJeH2jg0rseS8K+tklt8rXXfHsbtuD+YyjKgs/RRZbuAluyvq3QHgj44S
FyubPuy5SCUjX9rPos97SzF25mBR/GDBYKlfIqp6RtF4iV0ENuAsb5csc/KLNNU/ZNkwYWUu8yPW
AU63iD4xPTP2/H2vonW3wyrvybs5VDOjuRqkIjf2fM4KNACamkQUJ8el8AeYMBQBFX5+MOurJpl3
AyKLLLy1OjtrGTPg5Xl5IypzcPa2tOPBmTptbzLVxrJtZSIYLYK5KWdQMa5n2tEA5t5QjY8acduM
q5dm3f7NZQ+ULC4WfdxENcJetjxjryd/nZ11KmlPygsuxRe2KZjS+9QFwEw5l4GbbYx8e8m07rZH
bgaeW2ouX8PuOp/0NOxRIVbBGw6ZYNWiPuR0kiVXMhxzZiZle9vNcePq1rzMwD+3LXoXtvF8zEx7
6jsosji84o0Q75naJN8M8ErtfeJf15xci3LJmeWUDWZCGUf8WBBOeHUEWuIDZrsK7WPWaLo1dZJP
sI2j5N2YfgbJ0sx020NqPJkqg6v6wJhWYTmpwVvs7MQt+8/OZ08TJAu2zwJVNWwDqfo9xl57oWRT
6ZTQDXcdfKfBMhTw9UVUGQ8vCDrZ+vxvrL1em9WX2wZYrAoOtPHQz+F1ocZEJsiOgp9oMpxb8fZT
Efx4MvJhXBVG6qwARb52VwJVsuGgm46ExQ5UmFKtibUj9MjF0L0GKV6Hg13wvaQegF7EfgGLm5HN
QaGQ/oiVfozNvLIdZd9jLzKUozqAghP298z1V0lAcZQIEqEI+c7L2pipH4j8Gynr7drTGF7b4rHR
AxDq+lDmeQNxc7y66zadIrp5Ky3I8scf9fD91vxmfvy6vb70dfc6RB0VkLfaZNW9jtajd4fF+j4Q
pfh6gXJsFiQebVAYH94R+/DQ1XJfp16iK8BImk3dAahY/HILyg6KkGkvVUHbHbwWCkjczg9mANlc
/z51yKSRSW67dIq8vGJzCSgyNkULeaJeNnxwCfvBX7vPIx3OFGVOwCWRG5dB5lVEDboFOX6vqGrs
EKMyxTLEIHYqle8TsenyodEDoLybfoamQNc61talhfrmtDC+t0IixGmYamY0H8Jt0E4cbPZpgJjy
p6Z5IxRIAOGVerKynKxVpRGyeMPVDiWjyIiiL3FhtS1rXEFscc12FxNLuiD27HAhP1KJrjpXy3km
fj9/J/L8J5cjD+0jt1IvzQF7zv7E9M8zC5ChLG/+iR7Kf6sKdemAD1Tn2UcVyufKhS7GsKtm63GX
aByi6O1JEAK437axgIZPsE/qhKAqPhpYth0xIdCK/nn7m8x6nUS/K8ST0xxdr+NDS9JArEqg7wnR
Y1ilze6/qmDDeF+/cd72e+UeY22y9gEiusQf58nn05q2A3gOHb5phd7p1RaLqiWg97PL8inGSE81
UBOmOdJFGybkxMNF5qWuu+RD1wHsm2TSkGsG4xyDobVfbCsvPpiAcxCG7d/FdO4iaaVE2zNhvcSt
mt7QzzTTp8QIvQIV649a87DRf/XMf6MDw8HXOtRFEMeIPwAr8rp5bmhPf8OPMa9wBB9FwoTix/0J
BGsHwgTn1CzKf4EHsiEQwgxb3IPK7K6fwGKtiIpBI3ugkdSsv7MCzuxUxdBidLMSEtAE+pk+laM5
CpyTwCTjXcjyPpyYZ7I2/BeJsgboov4hNszEs91O9lOvIctiUVC4k0QkEnlOg6AOag2tP1PAqBdy
JR0rfRQRKNoeu/unLywNd6AuW+21/vyr0gJz7MyzMHv87Z0LXzYs2D9h15gQSNUtuu05A+ffmv8P
+WTSUPjLwCE2kAbGExNEgjLVNiGIaPlDebiz4CO5YBXXP9yiuWNxyTGw+Wo2LQ4uZoNPeFneVk/c
swkEElAXz6yRjAtXgmu5PKJqRA+vtTWbJNEytRPdBskQcVsuHoRTkgQvwrkyQcNWRPoed84uqTVy
cnw9NHcinXU1pYqXXTLFiV95ptwjd4K9eKQZ2uwhoDsdAHGdhuH+RX+f4NmCu3kvDWCC/h+0JsBF
+QXGx/O8JZ1H289/1koqA3iUHBPCe9/QSoJGsB5Dz1NNvMSAiMRnCVXQsdVyEPdWe2SMOdIIZnUy
LFSW+omNsIXo82UJuUUKBUSdQvAFIatpUEf+11yh3HqZfotGgR5qHRhqdSuSJzjO4QLmNzh4fWVo
b9klIf6nvIkSl+QT5smvTLtvleZOztaM45BsnLjO5+E98kxXKOKLXwVUju0YJ9Eh7u68068VCuzy
awpt/hmyDH/wJtZeYP/Kgdo2XcMTydLd67YzWeeff1SzABUNHA+bnjnZC/4xacQ7lPb4NvArO4e1
VNFrZDJWASnOLXyaukq35yJCxmylEmob53uFQbg3S5rh0yNmNB5BJaKmPw7PyWtGQvosXLD4/Aib
fGWh0VvEuANLsfJ6G74Q1b1BV4gIW4211DkZQRiYxbRvD7Va5eTwUIapUvX1un6qtZx6xzmqAAi4
6YogaM+gTARdkTnQKPk88vgLfTgfupIuX7vpT/fe4ip5HZMC2OaT9GSsITGVHjVL1Q2y8d95OsMQ
7wH//TTY3CD2tWvrRXmIoJa+ZlncyFYY8CBB8/9WR/Mef/6Ix28R/cGZDRoOw2DG16AQZaneufTg
A17SQf2OoEMBiRqb6iRlRzBtVyqjX0cUJAS0jIUEXzu1jTpOWcTqmUTVVqS/ybEFxRFuW8GDQUFB
rMbwIQqzkbSgADaYNClQLCP1AlbUuEkMWHwLJlrKC/cy70JMi7KjRNsPEnexGsTb7huIBipDm+/q
utQzpqS1YlG3ha8d41/15rah5uvwneaAS6XKMaP+nKTy1DXHqB48/VzndskfAxzWq6YZjJ3WbNwm
cUVrWo60nmr9NT/Da6EaKjPL/EIIbOy1lIw2G9SoY1gP3WLvqaDlA/RfMWqQOlGj23+WQbGJ11ZW
mXbA1Kt3xwxOshZ9a+xLKcV90hFUL1cdr8ZlGUlGeyJWkLOvsJHN9Cp2YGS8/qKGaCGHlhisjtDZ
9pEFCaKhVlfJtJQiWyFUw4ElRUkto+a3hc89OWaaBMCzVrO1qo0JxD2T/140b2bYRhYHgVLv141H
DhCcNP8y95a03c/sWy/uZCAyCXXikq4+Pze6eAWPALp7Giu8NuThSN/RQsoCnuxPAxweIZJAV+/z
JAyF1jKhcjTDQrqEMQvBIQyyJf2ktdDjaVKOB0u+Lyw470D1OEMmO55H4XSewQSEw3DjOPBXvUOH
ZEboP1iY+eOg3zOA6ursGm1PIvlzVMYCVFMqDR5j5+VgHlpdRaVJJzDTOVTxaIzTzk9eCee68mV5
6sFoJxbL6qL7xgnzDFD24N9Bu4VfEKMtOvimefrFL8OWnzYHD/OThosvvPRvhZhjLdTbJSut2MyE
1eRYbsKEw3An7XWbTflAJH91EDoEyDVAoNBbFhA73i8yD47lKi+Bd9EWYJEv2eayb+2Lt+0/vjM2
DdDsGd+rnBZRDfRrbNFzKdXsHoMCwrxF7/ai3KFhD38yg/g8dn8C4sR9SuOkcR2AZvXa1/RVJj7Z
pQdPiL70TBKBlaI9UdGDvMnLZTB13n2SMEExRHeegTyAeEs9LhxOcUK3luCVpzsOumvZP40BOgEB
wvvWAPp1eD3AyS6rSSZ4UnWPd+V229n0chD4R4AIVFXOSR0vKKZ9esdV6oygTHF5cgVykM+R6lOh
oEFnmtWD1yRLTPo/Ul9dFLcW54Toa9FfyH++O+AQgCI37lGcR4Exj3N0Elq2N7nho3bQCE4tX4b5
q5VjRtunv1fXLc4zgH9FVJ/ZlfVNXt3QFsokeQQkXEKYgYyUMQsVNIVDSglQK/SujK5pxZhkS2ul
x7sZqxU8sYBLbEiNXTRLt6OvdlN/5u0DOBuyS2OjAbBIcfSg8/Ypw5LMQKpS80bPBcH3v39k01Rj
I7yfbLAQHMwFCJgKthxecI655HaoJllNiEVgIkz42e1d0T8DoD0FpFeLwO1idQKw/dSdfUHuB1W9
UtWUNnUisyg6/T/9VBSM3WoIHmXToL5QIGfOez9ei5G5nKyrdf+StpxJ3ZZbrC1qKrbcjtpTL52y
reSq5el0MrqbC7LnRZrL1I0j2lgCLKKK/r+4aLssUBwmqPy+3YpIYVOTEc/KbGyLmttlgeP54LFT
K8hrjPIW5ZCBI/Dbupqzsy9W7GdjWsxxoum3JMkMltmlZ4qEGV1UXZ0zx/umvR4OGExYwykMSA9T
niGXSfo6IzFBJCNUJbFtrHLAbU26MNHt9eOC3ZXoyCKgFDJHuMaTyTTBnJolEw8zyKTQrP8iEXH+
ydnTVgBPGaPfJc2FR5AuxK5SvCVC2l824uCeUpoGz9Md2npX2tPynf8xuwtoJWJp0gvILw2RT36O
kgLlCgzkrRQV7DkOPXOI9hjukfuzhduA0JrYRwQw/QkR+flvu2F0LlQGjBYaeuaHj7brf9pUAfmU
pNfMPqH6aTG/3UywPNNCWTuaELVVztJcJiJyc3o24lUMgG7RJ9URfEsg1EuTPF6MXhx+ErzmXguj
zA7chYAKtfXzsQJjuON0cI2OQR3HJsMn/tayltj+ZJrqKqSmXPrB/T8U3lkXf0mRYp9TQAyk9Qgq
8dYLa36ema23nnnqnd6UvE/51rsHdXjOhu1RN1dAoRhTh2qbN/J+BuElx75cykpOWka8ALA0hqo+
hvz3PI0wAYAIcUYqTRtLPFAXO462G/1VmmrC/vqtTsOBBwnxIONLZyx+I0Q+cbLWv2xcWoj8IENv
ptlyrv0KcfAiyi4/pXaSKKPBqefWKBLJJks6eqR4+TxYvhXaYHWxlUaHWQ1Fvq7mUnh0+PVzLv8x
ubPdYSxx47Tj7iVgO9Ywh2zRAc3lzTdKR1zhbYuKNtXbuWm2C8NF1thP+znIbNzb5u/kBDbCW6FC
cPkoCK41oB5JqeB5zhBSfD4KuAGLgfGEcJ21ju6n273d8M6ItSgBaz3B6K/uLgXpAaj4ZhqvvBBm
uzx15QRUEv0zr9BlE0tOPwhk1kL3mu0nJhPgy8WLnxA1ebQsy1k7xJ2J+E9J9ZTLfgmmBn7L6pje
TzUu3Q6hNCOwfLLyV0IFIkmYHugd/fveYJjXtBk1lL+knXFmsnMookUZJZvTLBPC4sw/Fgp021MT
c8nF8r/cCpzcw2I40gIDp71i4KNMAZGGg2Q1jEBB7BQzi1RnaU5bs2YbhZ0OUyw+yQE16EBNaMEe
GQe794Pl/wbAyaR5kqfjiQHebfP9yfwOA0jx5SY0ZVYv6qg8W1fOtrWITtusspKnwQzWHagONcyb
ZX8N4M2t4z2YUJpSx9T9hMn+T3Ocb1kiObOiyQ8C0N5H/TYk82n2FovFfr07NE8ocKuwvPwEaA5w
ezeOkP2yWWQLtxGT/eBc0y906a5x7dNdybMjyCXlVq81rd79WzWLQnyFKF0wf5FpaGFAItAOZ16a
r5TOtMMGeXSzc5VijM43vzBvVhTjjfyFGC1iGdV+OwX4o88eFoLhgaqWoWkS1gp0qJc2dV9TQTqP
vxGob3/ilPs7o5/9Frg70ZikkYosO1dleWStBUw21V6QCBP2waGUJ0sja+5VQDj81vOFoYgpRCB7
mO1HLvdoJpqY+xkjIIuewU9pHJp/XK3rgaf9zG1YVgtmADTtJ8cU4ZXnRv22eHPGf6auOd6rWIKq
p3qtTmsI9A9BogehcFHwtQRTWqHvIJJ4Fv9JQRTGFeduiUyqB1WKnhuH63owiepd3BYRUGnGCEk5
R8oCEpYCI7/W2Ux9bAKDdNRviCOyJ+kvw9CHXK0PuRsR0jKSAJP3kqJXZfSosNSYjxAVCXTeGqVc
lqDjZz1V9+gPrf3x3iN4XbmDRYMqDh3oFRrEaPecxX1B6uDfir7NtRFovJP9mNEmXTx5BGDwP+Kh
UvasyqylP2JTZw6U5xcZsIrpgijRwK/NBcv4KWNyKaSLN4ZSdTccy0a807gyvlGljxFfMWdxdtoK
h9TLdcNAJth5B0iGE9cTfafkJlLSi+m8F1yABhRBbfnkjw1BpcmMHm3Tz0bwARN+E4qJr+DMfvgV
2cQYhne9gHZa3Zi9nuX210dHwXFgviXQBJxTkybUZe8hpY7bY3xYgi2KZ+eTLoOXidFIQWaM9ktX
tF490i1kxI/3rgdfyH79ENBlAqJKl+AAcrvZyl9eIr9rNNqKTiovmzN/QrI338S5Du8MVfYp+otG
zwp08Z8zCw9mHUMFUtramGv+fo4+Ek268WErYcDi/THAL6DFUvZAOjsU2PeZDZKVQlKsBG2WW91q
2wkZ2+AzbwnjSOALKIUpsyKWfJ/njNqXpsiQMOaO+S1H9cH1rCKEC7pz/jTZHiXVTy+XkrGMhIs+
FRvHo/gvzj9cPqlJcQlDZS1DD8ovAAj+4spKdKaJEunCXOfZ5A3FZUalaGwo97Cb4BnSnLWZGz1h
4kj0PZFMcgKkc07Vn9euPXUYr1mP7oxQiFYpt0STa+JtoICyCutlBrX089mUiyOss1FEUpWxWe9s
hj0r1tVc1CZ92FCAQUOwhymg4omeiFFnl+7N9EEETTnpfSjyHE4Ux02xwHkQ22xdcpBpVMvliwWR
eDXyYemtW+jE9fVS2hm/tBDvaoPhpfdRFB81YCQM1GwedVZaFpcZnGynoMZU+Kkbuh/hMQgiYDXC
h3ApMHIBOxkQIG/sm45jyxa10WhWX2JLOFL1YdYQS82CnnWCWs6SyAruVuaabEMdSJygCBxZDACK
EYnWvmtR2yRQ97B9m6H/ORHCwd5OmIUK3Tq1HCpkWXtzeGfv6oy8vxyvGeRSRNSm9iBD3HtOX1FZ
OtoIxvnz+dsrgzi4fcWy1Fi6dAprfUani9e+aVA4W+AMxbuS5kv8/Wzia1T6KeaNP0FJ5U4IJjga
8vpjpX+rXWq0NaZj5tG6aWigRYrpZhJxnYs/o6Cep/KOEMamAAyssZpMZn3/6U4EBO9goyCqBT6W
DP6PLB1O6yrdAQG/HzSoJvIU5Ej73w4DPIrs1eNQh91gtbhXUKtSylR1g2nuxQK5ywABHaTqMJc0
37xz9H1f3DkjBDdDhYwGkqd+Cjs3b7VNUXR8GYrgxaRNZ9PUv7Pl/V7WVT5Md8dzpLP159vMuKRn
pcC30MeoJgjSJlTtqLqSs6bMQeSR8fvEFemmiWnqhLmZZM/U+FAR1T+BEi2yflVbZbQpRO1YPWsz
OLr/FKpfXPHa3+FuvE3byDFTOcOi5hcasGX6rYbaabHaQj7OUbLxEJBF1VnSm8LiIKXSuyEKn31s
PA9yZjof5024yUvKzp9xuGOECFn1drruo5CUnsCQJ4BS/a2OGMft0oUgvo32j1o/S+Hn2AjWF92s
QBY6lv1jMNOO/6omuQaZkASHfYFbgZ0dJ5ikAsWRNmLs9QAnrSA/lqFGbbwJPimticW3ZpvwRyTr
qaUFC9VK1t4Tf5QWpfKqxL7tHA2sW6BOfW2RehS7T9herHJdEg6I15JIkWdA0t2if9DmsDgtl1Ls
rXJX55rkm/MTH10hNDLfsZjLvt3mum5Coy7/+OKmFPGA3YhD/+uQOwBlU4byR3yF1IH0AwuAjc3V
NpXlc6kLPfqpi+7LEjHpCfcnXCmaTGYSFK3prUE/ngFb5OARx47XkJn6WD2EV55g/rOka8WyZeEz
Nd7y6riDwjceVO+BV0NAGXq/5Kcw+eh6HS4Bq7AC4ViBft/lmUQK2BuDHKf2FF5H5oq11BqeIB0V
kHFH+ATSMOjfVL5wnK2OwVX/drLzvrk3JDdLQI9+K++5L0qabnnnZfu7zOv5UUe32mWQBSNjEDiG
jRJph9cdfD2IalTwbuk4ka3sFZBdVfsr6BKtAGE4YE5IjQsbEjd6K5I9p72C+Ug/mZiJTDDStcQN
TsUOef71tI0FqINgaMRRlmcKcJNqN35cR2EqjjssaXE/wXJjsEFxA9oOgDSzOVQofEWmXuTE5zCI
Qj9Pj/0owwLChegxPB6zBn+QpV/IpcCTIOg1umKkXknGgGah4p/vUdKstLN+4guuT63p3nI1iF+2
rYzghgZ6swBQvMJXemYeUqNvHNT4jXbn05A3Cc2ewiP8bQbwFNgnHda98tq0SoGb6uR9vLSI30Fv
ha+JQi5KUR9CEz24bydEV8csLhRGz+eMAIW5zHi1aZObEjmhy95WjKqlQ4MWWZM2FH+iTR/Nz2Ca
0obUzfnqwPJdDtz86gC0GkxQFE8h1h0U0zT8vhlAuyzWGdN+a9vukrw85ZrE4fZNI7nlCPHN0/no
963mYJ+3kuEm14xiLM8GC9njGlAT3lQWMybBSs2Gj85V094xxKo5o9zRuapX9SfDsmJs6NObCUYM
/l1ErcyzXM2yg/cJSAHJe81Zp78fPwgYDLftw/kfz7anvfM/C+ynFv2N6SHyl2D83mDLjjoTJOlb
NY8Q89upuF89UFsQQNPqCuBbs8JRDfC8HDwy2nHBjk9Kjf0eiJGHNVkGwLkwIsATkWlsD2SJ3xdM
narl+5pFQtrURjB5Ld9JHulxvmpXpFBYjzYkwqJ7x+LhrVIo1q8/RAqs6stJjRbm2txOV/U0g9n9
CHfUmdPUpIrdM18UirQcN87Yj7Up4Z08g8baUhsovFsvH0F3K6lHINBf5kRd0x/prMssFwmjw7p3
5C811/0jzAxjCWR8o5DbHCRnzU72whtG5cdWNId0FiBQSKCsBCiHQoN8J4lCRgmi60gRTZy3zUnB
u6/nsVs8qjnKNS3QeFtnWQiWT/U/pXrG5M0vBMl/SF5OAjUdverdvgEw1fVZLLSRenup5vBv+m9r
w50ILQitmJFdWOiij1do/TTslPLga485E9R7IKNPtvQR96RLJI3Eun8QNLQj1MEOh9DKDUaUqLQ6
LXq79ZyaKSqwOdKwZQf4DSK25U7E1Dow4lI3TKe9dH0JkI4Uae/z7lU65Q0/ElKEj0Fpk6tz35r+
4DGn9v1r7UehcwuHYi5LWrp/2jSOMfZxfS4WzwNWcgCIyrD9f0aqaPf45dSw6wDrUY1Y0L4tjVRC
lkK5enb95ysJqicXMKK1u7NuMbRJTc37cKTOy/PliTRfsC7CWs15UbIVUkYQwpGGEE811IWSqvkM
LQTdodlD6y485CjfhSQWajOCrmYyuw4XSfrD70fN6JUI9DlQIhKcmarCZuw+tM+JfjAXEo5rBL2n
HjQlOuqz5bfRZxXx7Wlrz3M0vZ3hnp4UQbNZXGiGY9foTJsFdLlpPud/SC6+WKeXTDmzmPC95RQZ
d8FyoLbKxMMmO73Qg1C5uwa9OLH4d/WCiLU5GxYtvwwRrq9b6lTgdaDahYvwOzreHYhlV8+IUsW4
0AzqjhhlBLL8bU51EXhfjnPhRpqNONwx7E0YFs/LfMZjGkVM1KfvzK1xhWc8P/DtHCV+ble9/PQw
JYoL+xbjQr2l8Rn6A9pFrocqFCHK71jdApRlzlXZTpVtvDyIYLaqISkol5CZb0BoAoYX5MwNl6/D
41aiSVGN2T4VVrTrdcLNqoLmRvd9+54d4wvON2ZINJEwm3uLQ2Khs0XKQq4nauPorNw3DYnSp28r
hOAENdLro7U5f6ROQN1ICBhVTBgoFgBCZomUfhfcqEHQ2XIO6DYGsSW0D1Pt6BmaGGdIm+BbFVap
WWt3TXrEzPErr1bZgaTJCh6nLk1979ACj5zqdYEV4M546lgYKcmYDThvshd12wly9qu2tlFpICsM
Lsq8GTnoccwfBg5iXR6ggj9SG33lwNqHZSas6gYyN88Iwxr+sPwsttUU4ywcOHGDj70I/fu/ILq9
vcPTzTFWcnfVm7aDYSWS9FY9Ui6QdmUeNSuaOqKBFJRTGoXkmEBfp6Dm5HNzTEUQvAIGmlh3cvdE
S6T16mzQKVxdmplP/6GLJPtY43SqrV0oCwz9lZOycqsavJVjhVqdQMCSf2i7PrWCmC0YRiIFTLA5
Um515RqY4PcEFjN0yP/OyqOi6tOXIOVFkrg9TUSYwn+bYzHwmsELVwGWNdX9+KNLisVpZ1AE38HJ
N8aqPAvF+Xn9di0XNtZVjrzxkD7MZP4brL1E9zdA/MOq5lacsRYOBKCLYPHfY/Qyu/irkei1slee
TIzLllDQxUeYCP+INjY3ZQX3U84myy0mcJR4bDu7MN8kpc2bKa8eg4CFmnD7lo/hQYZf8QtVv+QT
LhHTPZKu9Z+I/rNCHor2Oc44bw4wWGRTvj61Zq22GFBgBSw1hVHC6+maaDfg05a2yLZGJLC8b6V5
JlJfR/wx4zNix1WyTU+e4vqRYoj//KSX/M+xGebRageU6dhTYeqEZ0hcdWomGKn11BCyTvDPxIMH
8aCBpjAOyFjOGixdD/bonvnv3Hsp1Z7rwLFsgLnnq3UOesDtq7dHt7jORIwNfkIargpWhSiRliyH
mhCTdtJMbml4447XgUaI/FVH/7LxTcRa+bi1b5+mC/Tgmbb0JKjLcqCdmnC3uN8UjwFvWvfPyKVm
D7As5bXU/qcmTWAu9InxPGV6FpoEZ7wuH+p9XooWRtbH7OVm+aQugTG1EnJ9WkUHlKV2noZmM4dC
aTfBAks0EF9DE087JTWuWnwcGzi0utHXc5cW+0Wau+oJD03Mfw0ftS90A5VdKmkSnUIm1jFHwajh
7eQ7vLU0Ql63H+ORSnxy95rF9ZpuBd9Q9T8bSLXdf+ncG99cFwa0rVigyB4qVyiSiekBkCPj+XcW
MNKpcueNaVlBruEwZZL3b/ydje8Twg6ozcIynXMZZVcu38c5gYaMMMr8wKHBNYIHpkYAOo0hlitV
PTtV/AAHYq5KabzGfxQOchMRTxO1I7kNX3HwvKoq4Av3QYB4GESF7+Vs7/Tc3RFF/6fuvg/qEFuV
8I1xZ7en0/vFhFnkimvRx1LqPCCCTy8vgdrC4Ypwac+RXnC5W1+Ez3ia7I53mwmLkBke6auiyRQf
PKOW/uVSq+9S9r/2MSfEadfu0oJTt+vp7hL5OnRW7k4QtRNoIyaUnRwaxgkO0oUt0s/J4VrwKJnY
pL9plxx4fyKlr1p/zXFhaYI8lYEaCTxWdBOn/yOv6rbV6giK7cG986HuIYXSaoZ6afDzWFUpa6HT
IKJ5mVs2zshYbb+FibkFHMn5RbBAFx9X1ri4QFJ3YoogHPWMKZN9vChAxxBqSMEdiZ/j5HM/HrQY
fGShgpHtN02LqE2GGHaMac7QdKiWXAnDb6t+n7otBUpcbNxIQbDznBfQORJ3h5NxFkDTQFm1zhXg
mAut2fz3CZffZIP3XVTmvkl1mU9Nf1Hm7NaDQXDU8X/rOGktE+Lp+R3HznoBdDJUIVOr4dm22sTw
M62gQjl2wqfLWB5/GUrSg8U/zXDi/D6ztEXDvrcEHgAUdWVQ+FZYtFm2p2k2ko/OpbqtGqp037md
FFCL9EmmXAbwonUcjlpLcCSuQmkV5oqW4hQK704XKkRC8nSSugB4yzEMlujU0G9nkOAGQjtDwIQ9
gSv3K6pJfIjkIK3m5GihfR38aEX236Rji/MSs8UZF+7hISYLud9wwM5FzLkku2bF0s4JemKjDidL
Zdb+lkt3UBRi6+kRmD+TUp4/7oOI2BHQy1Wfc0BNe9pruIK5Vt84Bsm3md1OxbH99TM1XWMnLwcD
c5OxaDb/+8P3BMcPahlJ4chFK3IaHzIyhSUozkBSJqvvzzMGG5wc8UlisAEg7YDmYqkwSEG2CQb8
IHMiB639fwp5KVklyDY/zlLpgPBL1K/gx1qaRVhh6vjgE8rsuFiEFzjCbNb5UnMa5yJH6hhCcbP/
5ZSaKCd8CEpiakgSwhr4trvp9lqgq0LrNeY3iOoQOCvB25CEkYGftby2u68/2NXYZ1rfGDNV2lS5
GeJUGKdtC3zps2p+9cek3lNaKh3TPJPqELWzQiXgruKtY6SHfv+6PiTMwCQma2Gp2O2HQ/e2vsUz
3oJsyZscPwZePHE95rXVGb7elZqNihhTyE/QrLUdC7gawDU0ojISutaiNNEs7j8l9/9/cy6cR7He
fTCDcAPefB+fFwsYp8Hyc8hCrq5UA7aElbnrPhb6h0RvpSieKGb7FzuOAGJMvNhqndxCB1Jz6uob
dXL2u55ioIAEP6AEeQ28hlm7oI3iYXviVGN5GUGtDa25/5Z00D8E9Ip/UezNq9wgcU/6DVEkvNth
iYv5lEsarqJaa/wcErMvQVPHX4gRSU9+/nl3UJInexjI5afCjYE+0U9VqX7q+wHwFP8PUnWgNd0N
Q9w25Vt0261o/JfzLv2i+CdD2EQiLZW0ThKvGip8KjIwGPYrjlfGhidzeUoEwhGRtGzjef36HAFc
YOQumzwZoRwEt5dOgZQjQKw2O4X9vS/fZr850ma19pndIMjPmZgIt6woZkuBhOHs0TxCCu2iKJPZ
4WyEp7c0SNJtfKrUD7RIkWg8B0iiY+S5pEmptqHUiM9HrcP44f9vMbm/Kakd9TexZHE6lpwCJoWm
Ss8Pbl+LDQ0t+u6s2eBQ2HRTmZvq9JVc/mhTlmWr7Pd1C3HOMBEfDJ4R5WDnKA+QrGSVqF5VWRi2
tyDRVITaAp7Kf5zaGNe8k9EN8X9E+WVR6o/9piRlZoW8ZYTkPZR8COT5u4H9W0qzKM0/b6T+MTlX
vHtPQmv5UbYzj9EOX+OhFbHl8lM6dzXNWPece7z2b2YPE4ADgDrj80ZcTmiQyMfioYgAVpj4OC+4
niynuf1z/s2ziy2HwfcYr81I0YnbgRjkpfcJ1KAJjhX3cAyadBldNJ2CMRgHsSwbmKAIUGjWviiy
QYpKS6SBswDJ/pLBkZYORHouoCnzrGrSdJav3tamRe23y/9xiNykldErdr6yllidDB6Ad9bRCGAR
V7ICRffS2DBKZrs3yh5JQuM5xvYvRb4V26GbrOe/BePb+IgB8oOEA9TvydIlxX/u/KiXA2aLQlB7
oJFJ8imdSeNqKyydTSv0uyy7wcBO5QXq9vOdntPdyhqbwr+3Tf/i19bIJWRb3jjdC273eIhhmJf/
G00cbF080sit3ZHFmBE9dNcsmfBy6l8M0jjgzUOCgfU3+D60wUZTCnydsI7QIcqPwFSAyueEGD/H
36VTbG9qDaTFFbRdWFALkwUy3umGZwTyTtLLBGCtswdXkdh1UKK0KxkwFhxlb8Suytx79kQ5cfgp
go2VC97VacYHEWmVEd0ZS3jXP7NZheMKNbXjcqaxrls/r3RCmU8H3NTqltaX7w5/5bxk+uMGG+0f
tcR4WyxE4deyWdK7pbAfKl+ejEmNLGdQ/MkLQw8XXUXaH7SHkq6M68OmwfoNGHM7EVG+txG7M9cb
s8UFBb4bdSCt//MNRPoA+jzQOOGFelC0uR+ScIp9AyGddE8Z5T4LYaAY2jmsYWZ+QzMAyFiGYfqF
cKqm7JfukMmbx9UNu9moSUX5KQvQiZOApudNWbV6KZqijhJjNQqAh/CQGiluGC3/Htpi/RAwoMkG
c+1JTOBOSrDALKRA3dAK6ERFmELvpdBQ5gVX5GQFnIjQNWHdVkZvwNZJsdiYvyACj6nMrFiuIRe6
epl8wfy2ufZ0N8uuYRQgvA6UCsCeTGdEYPfHPmrNxDS4x0z6m1duHPp6qO3H7J66XZ/sZhZPBrMZ
3Z1BQCkxvhJ1MouL93SCmjakUYEh4C10Blg9WFxWlgPxqQB0xjDwG+oroAbBB8/ZxQvHZbRMT7y7
QjQkS4ccCK0ig0mZOBeOQxgslkHnhH03cZ4d6i9ACzWlUMPeUBAGLcvtx1r+KTdMr/i5A639x9qz
U0jjugSIwXwzMBSMRnQjQskSRZ6YIZAQgtDXLslxOeY7zAWrMMqYkkd5UbPBx1+R9ge7n/BlS30G
yni9oeU4FBzdI9X56YI1QsIG+SQjeL5tjQQ6mIygVaef8BbiKPSgf+Uo3qw0fS8E6WcAwiHRHkp0
dAv/3jAdLpN5tgkuw3GHhaxw1eceA4TxMaWQ8bggnjREGBgZDY2/AhLYAf3GaF2IJTBn3aQJ7x1v
pp8QtaVsP9g2w1fDuBbegdmFvscDue7Hja+TvDr15FGEtZ3NtEZz+GgkizdZhf96pfm0/QOrEOTn
jbLw/rQ1x+/oM/Uqhx89LAYWctOhW6d1CtwaU5aU8WRY1qbgfHW+xMbvfl1AFwsS/ZD/eHDHcBw1
N/q6tLsfLW1+aC/W5PeiSCeIWtVGdPeNIgTxGObsG951POfaeQhs246R7Ht/utkEAzon53bfD3vg
l79asSkxsXqVZYVjlLs9EsOcJ2IZ1s7ES2S9BCTHaEgOyvFdzXw2gn9YwWX+xdspK3R26sUzEDT2
2mRhmaiTiLEiq4tYUvSKCuRIQlgo2xM9AsDWmjDujdjE/sf/kiCQMLCi8fJpW3TK3+1yfwCPfbsU
a1VQQzNWDz6W+XGl+hlJdA2JazItxrShTQ/TYIF/UEIlnFvrOCKRLFgqcOIBqQtVjo4QK5KHllaQ
2IdrkAvllpX3LwhWK8D5paBi3YGsci0LUC83hrwG71fUHJlc8FiT6SEBq0fUPKN00N93bGB9ebhY
Xu1+DHDgWJEtF7pWcRMYRuWIa+Zn3ELF4AItUIOqiLKiExOoNE44bis51nVzEks9kEr0yRBX8ssm
V33S3RXHyJSwVzKeWONkTjM8QOpC9UHlChn5F8815WSc6TbYk6Wz+4mkFf3BC29DKOQ3fr+XWXoU
kv9MVHWt+A9OfBcXahXNtY80Cj9gxTuSIrlo/Fe3ow0Xb3j+/1aEEkMoC4J0UKto2u9f3RvfHjmD
XGqDX7SyXqZycKJjscqMESc9dx7WcHmYY+VAAEY0XJ7MiTD8NlfygRFqYwkE47MXFy+MF+VBMO4B
dX50UCFbsIChBy0PvEp5FRR9KGogWsSnOLJTK1DmJC3aZ82NVGxzCabrE5xj//mVlDq/U20ohIri
xZ82sK3xK23MDdLvUlJCcJPPjdWEqwPpvKaQ6TlcGi7jcNm/fdVwuSYKqeEipxrDDqbXO0FNIBDW
2lgxHODhvYPM6zepeDUhQ/xWz4JYXbMPRU2ESITGX3NE916CojjzDxZch4FcMLYMjriIgih3pS4f
ImU54gPiXoAcD7JgjRMqWNYap13qnheQFSa1IZXPSkCcxJQTGQWW2hr/RmyXbd/3TKkU/Ny3r2GN
ArIfSZ/fI3C6lyXk4vh2gYk/7TFyIadR6KCTeL1UvYXddFoT6j8Pb5R/Of/uK1eQBf1CbFOZTIwY
wOekCwMufZFEvEEh5L8Xu02qX/cqOrUqlyCLZXzedo3ZOz7hZA6RtrASffltGqE5W50i6jduZIwZ
x3atXk9CkzxyhL4nO+KNgbYYq92p/rMsu+I8gboNqFakuX5a+7KryhGWwfC98LvmTBDsjxppH18z
togYlkBS7NoTAC5sAXr3TEJwRtjnK9E39bBCQ1yWOoZ5BvR4WRje9QRAjg9a4EsIm/8D9N3KWMAb
IW8px1MIjeveVYovfR3EB89wI5r6tdyOG+yWlL/XeYBuu/TblEPMTAMaAfQYVZK9klCOYZX1umnm
aJldG7osOei4+CF7bQy4TTmpR4VZ35pkp5dbOz+Rljt5Gz51jPkEiuO79P6qr6VmbiXKmSPokkG3
KTpLAzGmUUfVFOsEyD5xI+MeyLONfvlKY2gbrrC75ba+m8qVfKJwXnXVQDKinTjcMTvq19flxqyS
YlJDQy33zwuWopx7RpgCqj+mjkdO0G6nfkVA/6LEccWSIVzR7xbSHft8cURsT+BSwuYfs2WMAw4N
Ami0A/G7+8Wj7mLVP1KsaFdUu+ahoW02vT3peGEu0UfM8252WDvVw4yh83RUuGUT/75OKr3g4q7P
Ia229UGz7TVQAxqkagKy9NIer6a2F05VBnJG5qsj2lWFkLT0ZkkfFisSv+2iViXdwSOVy0Vp/PeJ
CpiD2zrYoE9W468PcksonvmcOhn7TqIKjy7D3LJLxJy3FAw0aU9IMANU+Ze09hRwliyTH/EvHPPM
pawWRkYrCibDHmcQlV1tL2lrZDvPJwyulBdBKZcIWhXqeLun94JqfHWAFXGp0LznBnPws1D+eqSv
MUvQBVIZu8S7LesxInM5HJi5MhjN01O/krQraTOVAW4mm1UIh+Zft3VpEhix/2qZ9Dxda8hKKtWw
W1MsvFM2XDMaDJEUBZFFV0EM+RJpVJnk8LwtT3Nd54IJoMstwj+VcGVr3ltO4IJELOKAmNuUb+sJ
D4IlkePYEy1JjKaP9hLp89uv20uXNmhei/ll1WC2an2BeY1ARZKaw9F3xULei8vNXqRJsm0/b/Pp
n54pFrgQDvcglyaaQ+XRgYyBmo9fIIHBZTGiD+YPA30OagxjjLAlZ/0+WF0fSYHhOnpRzvgPcWey
DYj5r7yAXWonJcrwgl7smuQNJtymrpdBLT1a8k+PiORwcschuoydQAsWogqSO3UGjNR5RR1+VOtY
yxU0TOwKD96R7QTkglVmjCppd3LoaK4p5IGU55ePLFQN8c/fQVfBP1pxl6ePN6bCWRcuN+8sYT7P
z0tEel4knY0gp15cjWtoAg4pj7jRRc02USxzhdYqlKhBHcnzhClMZWaA3YCtNqeXGntI/jrRtGfo
naxn+/60aeNUZ+DyzQXUHX6KJnHrAjKL+Cj4Y1Qlrip+MHpSpV/HzjgZaMCIscy7w74htWIWJDN7
Q28N+TnHlWJDGbiKK+B7wZ7uMZ/iJTLjQmim5+0eaeL3J4Fz+mo61yzYbwbIL0Ij7S91UqxXeJP/
TFz+grmHRfZz0afkkRZoLsZyoWi8Yt5o6SDm633Q+CoPMWE9W8es2aO6NelX8kZUcLCL2kyOrHVE
jqtv5T4ohGUnCFHp5FMdEGtyvP0k4v/9T0sdyu9XEJNhEYS0MbrI2JrL+ffip9JrgNRqq/jtz7dZ
Y43d8LibvkmBHuQPEN0dBuKxX0OvfIMS04iic8OLsFUX9r0M5Px22Ermy+R1vgf47v/UEmxb571r
3S1vb0rNo2mt4iK1X6ojcqQEUJc7udqoreUNTZWzQzCdRoq3MmUZSEBS23QGFT3XFW/xbCo+GuD/
UzVOPNArZ43EuaaHVOCIymCmbJDsH2Qk3bKCAkr1hc9qQbj2EiQsK1bgpgyhDQ/vsCZFoDjLKK7n
ZJsGE1rpy1hWIWQrb6Zvq9QsAQyBM9sWN0MzqbgRC3gllW/y1z6v3amGxdpAxvCiCAMeClWsXRl9
IHr0mbtl8kweaQW3BVh42SixPC98LUI3NaqTgwY9iK2oWucuPvPbT7WcTNpeV1KPD2347xHMjpHq
bY0BOI53mD3C326KJsLubxYLEZVOSfvPLAUM4Ce0F6fCUVKf4X35EtfM+RNPJqa+9sEaPYlcFuOt
wUOgpK5w/wE6et6WfGrXcRJZ8lawNqwqF8CwqelfRNbKvL8zMnQJpkX9Dhy8rUJaDvrJ8dVGaqUm
Q8FmN06YH+QCU+EkuB7T2LxOgZaYSGrIsx5JqY0nWpc2aV19U/sborxu3UpxTnkIalM3p3u2HYsL
gadRRwsesb1yNRdZvPBrq/MIKBe3TbVon2o1pkhN6pKb1BrYJErKZFai7nAy1IRzAt3BOUgV0jKY
S66TWYotHMqYoU1NprtutfJK48+Czrut4+b/dq6EyE69bEHffA9d9ZqcaAswfKrxdl+Cj7GKKAyH
bGp9ab/b6C9WAoZgZ9ND+UQLd2+xGqWpYha31z0K+dY5XFHZGO1Ym3JREOKoOx0utfcOkdvF8KO/
wVFqMsGk4gKNWmOWkgYMr90twaRCus0KxkLHCNBMw5dfLQynm51EhvgN6A6r4pD++BLYdedOcMyN
5wdADVP6vTJNCwURlu8goMoUMvddOSKJ/U8lXkzH3Lf/OJPy9WB+0Xc8pN4lVGTgzr3vgGEeNElN
zo02EUBxZbEOmFaUwsxmPvBWBZDePxfPWtFDafteqBvQbU19RlApsKK3h9K1P/OY+iqLohG/Fn77
Sfp0kTuta3saKZa83mu3c0ray5rUVICrZOevC9nn9DeIlcocL80mm00a7pvHewzZMqZ0lwfsh7Pr
VJNlLSRV/aHqNh/fDhl3BsEy/gIq0jL+gofNxwqXrvTag40cNREI/PTFdAKbgxOodc3AymxfS4av
BKHMeSVQyKvut9YQIJCGMUZZy2hKJiYdhx4UE9gP8D7bhvgowIxaGLQaG1fe2Hc5PdQRahZR6nym
1T8QlpV6MRtmyo9gJhAubcbPKqP8Qz/GzF2es9qGcHyLwqOw2rusz5MjAxCZnamCnW0LRsNGkDej
9ld5+QZd6e0Fga9b3XEPrXMoJBxXN6IiaaHpL56HNHTd/PPAKmtvnUB2rFFaOWVUit7H2UrfAor5
k0QM/4CipLlKROe8dWtBKJTALp6VQmuutrTzY2PreaYB7AlorF1eJYHNeKLVciY6FM93l0CA2ed6
1wshL9h5++BVxKHMFzzwkuuZ6Rp8X+0n/QQincXQ/tqB858eqktX4f441boh5iL/HekG8tjlCF7A
5Etbsy53ip2hbPHBpD5co4XmIxY1St8gLrTRFJ+3tU8KKFOJRS8SLqHyGtNyRPGq1QlExnMnbBeS
j4NBJdkd3VKCjv5XMUklYfgH6O22nIuTaV081BwWaw8JbbXFPmHOZ2d8DDMncTxJ67U8tZe3Pyqq
pPyypXBTviID8eWo3w0Bzash+8HfZiym5rt/C9Z+Ty3DBa1wS+UVQYOVBqQzOiQV7sXcK04GfseF
vZKk2krxH1SoQTp7AJKlRukaCiwxcWZKqr4kIQ8ggdZusEgZowB3kMDjsAIF4d7rRP43Tazqw2Lx
gkKRkomu1/2gN1zHwR3PwON09W14SN+0gaDoyCZnkkoUIyJ1IUPR/ZI2LIAj+0n3Wr91d6oTEEJO
C8xb4SSpFKNQRPBzeG68iNO4nZt4a31FXCOoi6J7dri7Djnz34gkNttX60PWhNTLtaNB+S+3F6An
8fJx210vR+LYv/OnoFhYS4YmSjQxbzGIleZcISU+pzSXAjW2xqVqPnaTqcjFh4Sx8t4D78/eSPHW
coTaE1XJK8nRhji6eojK0tT+qxjCvrd4PIhEEfpmbr6xZ+52JDVV/ed/kY5j63cCphGZb/HegGJq
9U1einIAVyEbk7tdbsmbIYzNSA3fqoznm/FGm7032Dnbavf+4NfIJskbKWQn4ItcO1DYRkxF+1jZ
R6N+O36bBdwy1o140RmZmIKT/qZbcvupFAtxlDer+6wTx3wVESXk/mxh5X4IXEUW5RTyxbzxzm66
cjYMkQFOVZsreyffJBHAibK3SgOM99fOoZ1nw2F/5UXJO6wRnEdHFLSZhEovZvTNpgFq7XS5kK/T
3WZVfsRgGhrUH+QkJa3aDiyYgsKjboHQ6llzSq0dTK3/ChDsxCgB9lVCaNF4B5PzHnU6YlZhGCO5
wFbHYVbrAIuzOGBptU0ipV1R2Mk10djXFpaL3nvVzl7EcfBIgp92a/2xmQaUdqdMLfZjh7dGHmRO
R95Ab7Xv4c6uomZxooKZ9OJVk2pm9+65S/7tzxEwZqIJQh2ZUcdPZdACbbo0GSwTrFlIzGjMCgMO
7+mTX8S8on86I2l4sI51GYD4GImn1gMg35DcxxiSHbUzZdSh4CltzY3TNZcVaocKsEbJjx4oqrfB
0pZueGBY20YYZh4VAe7P9SUD1L2PDmQa1+T9XCvlS1V6+rN1eTuHTYvL7JMiYky8itFCBydjR+Gw
7xfg7UkICQom+JhxPovjoGzdIUdqnkfv4LCR17yzEJHh1G99O4t6DibK/woqbVZpElA7jJJhABMg
J85r2ts2pI/I8sriZDNcCKxxM/vxIxE59sAz+0jiEJl+WGfC79jEXVVNcK3eWyhV0jlBKWcdzwDe
mtv2XXa1Bm5PmJNv4LSAM+v5k+X2fvvcIuPyQqfTHPSigdNwOdHVzqerZm9WqoS3XOIsgNPmvPl0
5J3cEty8M05rrNU4MlXuie+7ewdNfkD1Vv8VnaFOYadKylfyMArdp53+8Hk+xDe8JzBDO4Muf44i
J+FLF3JFZAzI+P4VlOEr3TNFivqCn4s3CgzK/IW7AuJ3zpCK8ygNXtRCKqafMEaqV+Xpz6AY2tLc
zB1SHPJbYiwjw/Of/CAuMDDm4yBx3vFigoa5bj10Q6wKMz9OLm+SK+qAWLeIejXP0yUAaZKjvo3P
2xdi6tbRRxwdR2xyztrtHYqkwTNlJu77BAdw2nG98KZ14/z1XmxsUuNfxWLFG6E49IrChn21ABzg
k/PUv8wcrTGIFqRg0MKjeh8Js/U5H6MHU29ZIMn5UjNSM3/RFWgrBG9J8jTmE1LOiSXtadVuiTom
kDII75iYsup/QsoBb846q2eI24djgR9FmSU5JaGCbsMqUc8QyXQ++1aAtq095ggpmLs6+kNywEn0
rS+fJK5DvyAbrzkYDARDgPc6dgyeBineFMI5788dkvFfzUFWMFdnyewtz2c3zzh3RigH2tnzs28R
NKtJfoAAVNpD6aMvlrHZCHeeUzR2lV3zu4ApmL6JpP0D8u6jWXcT7vuz4IB6zDDaYtyajJOrSCjy
M3rV7sigjAyqKPRDBMDegcdoGwNv5qIl2Vpb+4wIVgE0c0Xyhk94QhQCvoYtXV1TeK/WQrgbd5oq
iEhRlTQCn/klWZEW5/bhXLST8Q+TS/qkAbzF191eIoRxxOoJRo08sEB2R3jC891HaJy5nRx24/72
8w9XXtXHXm9e/0/13G4uE3FhF9FDWmAw2txqGPaFgVXnOr/LM+I1z9PjFSX+XAQSoHLbxY1aml8b
3BKz6Gx/O4rvpWk+oi7nvLknbwx/nBqMl1VClppyLVBk3C5lbWGFkBl5+oKjHrtJOfSH0h/Vzgyq
O41MPNBbaZzQUoU8/bJfX/TNo4XK0rjjGHQXdxOQXJH2vMuMFBRh8rAJ41qzHhp+Kz5phsqQF0Tw
KRk/KYHQilQ6+/QtlGrKoSMl9gheMvkkOSHxrfoTJ7OJ6XTQEfYF9p2z1BvfsoD/GJUmAyf+GM4k
yiTwHzwtlP6R+9ASrQ+vr7n8P7HI3yynoroHwPG42gJI1iKA4oPiaTpAG8YuZatgrX1wqPakTfnH
beJ4qdXytrlIbyGYpdfWGhVFkX0lSoSz3fGIdYQ/VTZV/orUIYqlhuBI0EN+YV/XGSLiPZNIyaEw
X52ojA+fw3Y7vnS3y5lcOvLWspV7SfiuCqDo99y9vGskACd6ZDabuRRh+8NUNvRTUZdl7RBnWMhK
DNMSYfip0oH7qdtgo01z78/ia9+ELQPg6axvfQdRcz42x65xqgEurh0+TrOVpsS5N0zHv/kSYjrX
q5ddC4xdOrhwEVxVur7jgFslAk+YLrUk55RCFJn6wy4rSHQts57897tphXOh3o72eedlWLBPlp5c
7UnW7mEXXE1JJGz5AJAJWqxk9NFDDxymZXg6AfSFmcDwgs17g1fuDCYJonJohg4EAfImgUMkk+PG
lvyOleB2f/WYY8H4kY9/HeJdkjAE0I328BZnp2NfOSGpI2BBTrzGMdR91mkQY+3ewsxb6NeXlu4O
wSlTTQgd+R9t5y19VHWRjuqrkPVLW0kYA5FwdC2l23OfsVK40s3e2TEGtkLXWqLM1n6OHQHjrNMs
N6EmaP5zRie9DtmPT7yKOtvGzvoTWCpJQCgIZSnwTZaxLiiuX90vB5e6Uf8AfiQjNcDsnoo8AjOe
+CGEbFK5sH/QYExS4V8GagCt3fljNVp2mzwCH4h1ZLRPlW3XbqRSad1/Uc4zzVfbXZtBwaF74/iO
R9gHWzUB9o8sxILJHOgFwu0omUbFHxf4zsGI3C+JBESWsKrv7npG6CHKnGgS3N8VxiHsDCSx0aJk
xlOaHoxmm1zlN/TdGy71t70rSP7TxI5S2TzidMqtNfwoZtvxyMuXSUuiqYtuqmtBe7y+Umbxlz0z
BvRlSAyf2V9MFUNf2fNWNEERDYNKuxsQpPa2u//SG1gjfy6rq8/8HZo7Ckxh6lWTxxcRc7d2GGrz
QizVK8+EXOe+sOKp4doIi0y1/uTDtSvtVl1qj7aEcyn7u8hmt0Pyb6bdhg3pNdyKqVbkz58jghfV
zOi8Lds8+yHfdfBB3CTe6Mqibp0Xwaynth1ryX7MxbhUEiahoo+g105nONcsx8LTYqvI+8jabLgU
qDpiTFuTviceogJYK50CyZWgFvXiOkXZOPkKIFiKbY2zQs/0i2CKhs1WElKQr7MbgjuzGtsf8qhe
H+8SDmuLe6m/+lrhqn5zcAhbQNjGwBOHVICevXYXEjrLRvUEfFDT2hbmSxKdwDZ0ElMEd8VEaU1R
IVXo7jGhvIeXuVxjpfbTZAk93Aem6ykbl4Sn56hUvUBICDKjRuAgtBrloUsjjUessCu+sdr3pCLH
2T4cRzCD2WKHmBYMep6p7JZK4j4Iz4IkRIOEE7eHUj1hI76NFsw5zfNCtajG5fBwpukWue6j3MPZ
BBPIQ8Xv+bEpxlifu+QvminEkVl7mHIcV0/JZG1Xu2GK3xa9vQ/cSpUzft9bZMYmAxvmG+r7KH1t
JqISeKBLno8/cmSiuoTGADE20FSlVHuejradED3qEcImfKVGil+4JI4ohc0A0jbGeuWkRBzvgoh0
8BV8aQQiFO/vmuCQ4ZMsWuVGZY8NRg5eUTKMR09/8nkLmFaMBuMXVYGLC04seQ0NAv9pXwRg+cKf
fPKQq9cgKstDk5UToZTu21hi0TaHFvKx7xAyk+z5+bezTuHyfaRTnWuV5ZV0xMaqQ0baDeNBeq16
IgzDTzyaehgNk0lzU9WqZcwMBl6GhHsDYk8GPQoclmUMHMnm+PUIDj/So7/MguhKrs69GojmaPCW
bEpV3fq8A2V/KkoBJUbhfLm1AVSn+8o7RpSPk1TmJnV4c2byut5bX7eNXl4ZDoIk8WemPEnmWpzX
psROD54gLVrPsckBxIyWhv2A9oQQnntEq0GUVGcNmBBjuUnGe7bZOGiSfkC1gjdCBjsBu8/I1V6L
IzfOxQBL/DqorX4dVZ2tJdTv1k0BLth8Y7qmq/XPFrCsTWcLpMstOTHPHCjR91rdRosE4ulvUZYp
9k52MvH1h5geOhH5NYxxa8VPAK8qirD+NtU3feyeXvLRP2Af7ZCRDYwRrcE2w3LUx/9zSSw6gVpb
l+U5mGPh0kZonSGTUD1oddK2Vsc1PGO6genbV0jHZpN72CwMbc4s5/7ddibln9AVteJkuju2IThP
Nbv8NUCia1kzNB+JOYkc9d7bHOaGwh4SDPG48FoI0lzOBEu50ViPeqsTMet5fabeyUrkfGG1lZab
HkZtogiCBECf3+I/9nUtV8t60GB5ib1VcaDj2RrmSUSTMIc1NbB3dl15Jc6KBOv+QuQfLCzH1REw
mD0FNIpL4fqMvUZRKSIeW14MJh3/ZYLwlYFu7X7HQnUhrmmwEFoucyWGnjH2ZxQGnO/rKmAQPyhL
g/zScM+JhPG2+/FsaH2x4IvwUa6HmlOXZo1mAhX5sikem3Zp9Gd8oa7QFIqyiS5w62vKP418Bzge
4NH2p4iNpeh8+hP37AydeuEHtImrASOVjefY6GurgFzl+LbTUKWWGgxvFe1mJVIsMHCPBep//Yck
Cv/jQm+8ruEiso4FsR3FKu90kFCq1F7pAo8TupAxpEY7DNAZ3L730tAOylnxugP5QGUpmBDsjo/n
hAtfhZZVpLwdNTosmhGVc/2K0yxG2LuyfX8W3NJ71mR89eyw3Yev9cC+Gct/R4AW1drsBSVVjiXn
6VVCxj/7dq7Br3CoiAD6V/xdzKJnrRn+oavw6Loi7oRb5TXq+gv6rfCqEM5qtPqLnAShJBl32z7N
z5QcTA2vys1V/D5wVk+FS+LKqLsLCek+aYVajMIkwqTbbQikWV9wqcGs9Mivzk9rW5G3BxiaXcRV
6wPw16oqtGPJc4TeirmfS2TX4U62ZJ8Oux6Cj7E1oCY9UOLpz8Xq0Jktj7YXEjsZ9yxZtWrM9N4j
lR7aQtAIyorQGHNyifUmsXNe2y+gCrxCc4oJ1+mrNivQPxoIIGOHSz1UQKtSUa7R8Z8Nogmzf3xG
/1NgOLyvSu9d5lxyi/V8XAsvHOFMfPtRFiP2AaNomgwmtoVitYv6rSc7xpj9APZeGV18Gok5+yuV
WOwAFL/l0m/q+j6WLZvrcFCS1C2pcIZtMbdY+ST/ucZRUiegj5k4PRs6+JvoG1kYZBfWGcrxcTX+
kJG01di3tC0YuvVYQaqskZqpaPH/LTdmj9PvzkA7Yf9xGDel9wWRj60RdpexAUUR++Udq6UxuJ32
QY4Stg8Vdba6gb6IZhmW0CPpv0nQIKYZF91Xv2lNZHqd+zgsUM7RA1D9NUer40jEoiEbb6I4Oe17
UAaLRzKVIKDrhi956dipeaCpI3NQjtnkbsojtNBLUBFjNMMOvw7MBfyV24dSK1jLIK4LIS9acTKl
tHqx4rUMn5cMK8rnZa/ByiP9onu9HRZSE276sK7AZp1KozhyrhFiNu5KGeX6O8duH4e9qXqtbrCP
Q0l9BklA1DjTnVEHQizKNSPvJRG4h7wm3P92QMYcBo8nB0gG3T1uTlBu2BTh/zRPL+NrRYZN9ULG
ZK5SLwdRW4gn0LBeTpp7Tqbyp/FhyNFnw4Q6joWo+1p7VPgoyt2afrRf/ZF2L0feynIC2VZKrD2m
nWDoKQZFRKsZq5MbnPw344/M8PZrYBUvxQ2CFKuweJG5zNv3N6yJOLGzqlrXtXnYDHgzvtK16ttd
QpZJTYB6qFR8r8ec5yLe4l+prl70GSQFUHyu7ZqxYo5IIBfrCyYFZBeTubMNBPlwFkKYS2I9+N1E
myTVvj2wWR6/fEY8fZkvUEgtMcZUyQRpEM/j+qUs71t9YqVP9VJ/fOzpBeYF3h/8ysXPM58StxOX
E1IL1gfsVMOXa4efXOrgqILk7H12G42AMfdV6XNhcgrNizohnB010XXpaXz7mlhCkugzbRCRYxUn
+p1yDXvsUa+dzZPpFwMbYsyqVmYaVSddO9JNxKGAhDSxgLOjvP5yt4Jb93BjqJlyEkbWTykTlpGU
ZiJ9YQYHFtQ2s4+XDDpgoxGGhR+WAyR32lGsDBENhmNQ4lhucTnrzKpzV9I9tkLSz0sjXG1ffejG
toiR7R2XYiJCl/j/kmdq2leuRrRcuVQDoyPp6YZWeXsu+Mi9cHv7NrllumH2E6AYVhWL0FvShXRK
2nC8psm4rqTX32PeHe0oB1Sx8jhKZioO+Qq5pZcsVTudP/dqBcy2FbQiy4doSpDkU+vYYMswZqif
DJhK6G21wNPYSUCsBE4IKIhLpyT88vlwHSa/cR5FX7SzBV3XBEpd3trHcDatShWTE2V51q7zcC9c
R7Rbj7Tkx/qtXOae7gSCIqj2OyIlCRdOvC/vrl47nUgtwzZAfEpVGESjuzHQwGhm8C89CvNsHSlf
cX8EWPd2j2cgdkJfQ19eKQ5rFbm27YhtC82W7EKECdq8MHQ1Rgy9650vA6+db1TM6MnK8M7xwQ8w
N2/PWK6SJz9j97TIpwxXdi5LxH7CxKThJiNOKMBPfALFxnr2bJgWpb82N93/5eCPiqbFirl27VCF
0X/2rGyb/qwu6sjP7Zi74SDtDlRQALXtefPoMD3Cy+onl8KgvRuv2FR6P/mo/GWnhdf4CsTyM6Q1
IeAPDRtEv8yGb2XdO3+mX7VmmVTS6Kp6LFcyb2pkhHkH7vk5z8Z4NfmIdJZRDdlHz5SoCGR1PQS7
NstNzfvjsVgU15eZRZ+rGcl5In85Ugw+Sh0lkzGw5XlhITCyfPn8w4SRZ+rT3rPehlhwtJlaM3Nr
zAlEhuAaUyF6MohmQ7533hf8Uu//DcDMg4vOC4KceugCsP2hI8A/Tm5/A/vuXzkcSez+Nn7Jpgiw
gwhUZp+GidUpD+2buttFkYyOqLt7qmtG/Fyb6/eolEkPBiyE15cQz7p+SLjILBp4bfLlyKbjAkcz
NrsRye4Z04W+4bMwgtDFDQz1EGfc3ZEj1sGIJTZKt+3Omi8lV0f0ZkYRwa2noHILqBDuhCNexneX
a336SmMpaIB709FWVYjODHwMeIdm4xjz9/ENDtZMHommPe8aegTeuCYhaxB/pFeALj8y7MXJqE9V
6HvpWtXzptIcXnbTeXR3n5XgAKvSydeYNhSbmfte4EcjkSagAkQXxanpac28lQwyCIwPEd33iFoq
wpdliS7OF3Xn3Tjq5rejgQ7/+ks61/nlZYSKVOjFtDGx0EJmg4YlOtDSd0sTM3dRorKBZ+Ub7a5B
npBR+8nvkCP2TTllZuq/2XBGGBMEGxFDh75XeVQQlO2MlPdCVh7JkCBAbBmfuLpV56fkxR7EG/x9
IknC0N9lrgsQHr3dCek9Y84xuuYiHhXnhktES9wp6ii0nT0ss7edZ/d0ePqkakagDptQBF7GeT60
a7GQfy8XC6gbkEwK1kQdKMDyyh/dnPO147R2LyNRoDdx0LRHfBpopQNv6vnb1V9uJzqdESAybWTB
RU7HnvGu40CkJv64nwutYKXRueMWCQLmaKDzohfkx7GFzbgMQ1uW/ww2sbbXP9y05GMsgsBJ8+Dh
WYeOEzTxYvaHuCG2Z3x8vikgv8B14DzZtpASA09Pg5TjjgpwUE9FaLbWIcCwZrVaKg4J29CGJZCo
noXlKL946RcjJ01gWFAqZkLn0kVfv+N4DtFvNYIJ0+/mztUuWbtzJbyP1WN98rXCgW+LDQFX64xa
fu/vlGTg1FK9eH3a/2hc3iX2XppgB0PcTT2CC5t6gwvZdGKI1kFMX7+2fssfDIIX52opFcA/keUn
CldVOEfoZDAmbZ7YL13uVNftoCChqYMIQAzZNtrNSSLXflGnB+wGMnujg/qijGyWcG5ZpQ8scK0i
pGdqi5Ibn3CxrX+jTyXJiqWI8xRVZZ2Y1tL+FfORbvolqGgjhHkSCfa1umZjzCbQ7v0wCPnlekYk
9vQAsg6XxoEVYllrhTQ85WdW0qXZYfMofZBN5/sjMLsqDclxVWB33hXxUaSWqw4pGgpCh2ZQEql7
0td1ZOcWATGPzEf3K+gwfFIHHd1/F0kO8CTGoK7HoQmtZ+aM19PDMrleBmBZfcZAEENGCLpX2R2Y
+Bpt948sZ0/jjvgtk40tuSPRbwQ0B+MOwsDFqG7vGpGvgfe+jPo3qgOyppL4a1IgE6WICtUJ+JZN
XRrNsDFMLZH8vjln7E6BoNo5JsGO4WW9C/EhyxY5/fTUkBQJ/Av/1zPebEtseMvYL3p/8RpW0Uwy
hMdM4gAFnmPPuMlw82orehOJif53a89Gk4pUZddWYEsoMjfhHvqrd/URVFeoVfZofF06oJTiWREC
psw/vvXF5JY6vbsPnjh8/oBPNw2ZNaRgckalXinvnCv2TWCgYsxgdlvr6v0g3LoX95UBVJwNImeZ
URj8Paz+OhpfFKZYSv3DmylfsRjDu9YKnaiDIHQKDI/P9jpfZbm9wfmYKHK0QR2jUUkTA3AsadN5
BhKuLhF8c7c8A+yvYdbPkQcHASt7LKa9x0HfS/48mCcnPssJ3t/75KPZc+bTv7H1HVZAj0gnXUDd
tglcW/OB7HgjVB3tMB/Sve4dT2Dgk2km5v/BVGRkv/fjeXQwpTtlvQoan5lQmNH6cog0VJMcyFob
Jc49dxDDtgssgo8xZx20wQwI9C1mZwXTw2Gz1P4B8S1WLzoE+cyhD7EuXiZbUMqxU0fMYszPLxT1
ly8/Nom3umqrbVRiqJlt00BgxFpTSyZizjmpw/aVOrOvf3PTg55/zYahgccCF4kORvZ3TqEr8OL1
78akKz6jl3Xfdg3J+SWvnmlCayEiFRvg0M4IJ8xJjsTGYaVUgoM1LQs4HA4FH8f/0pxyIEmSH9Fp
vcyd+1pRfrp63yUUBrUDfr11HrGqSCYCMw5Hcxxmy1L4zdrrqmaD489fa9BI4Z7vokD1H+0JiR9X
nQ9efUpDOSM5YEOLN5ccrBSgCY3k7xSyk/0tlcsrKYBzA4Bo73bRZyZIqqM0fnF0IAnrZ5ZxNgwV
8w/trXgxsAB94mToSn9BT6iKm7AavflRz/ekn3ruE/I4mi/hEHp6IfrKWerOqTsQuQ5AwecghBKr
a3npKembFhCjsCE56VNyPLXTLvqMY3/vijsiiRHcUv4NPbz6ZvpmCQACUXl5SnM1hUk1H2sw9GBW
VVhnjj0fuv7uIgo401zFYNWTvNIJ6lgBMvyju1YFhqMdhExDWcrKiud31OQTRdHn7vZDEEYMatik
6InNWor+6tq4WX4IEOid3VivtXPOoeSvP5NvNGBU2043kccT1kQGXF0KGSdfOTeea21p7l1zc12K
mzSQAa0ypqrlhswmHf995mXXI/cYACrvDKhOtvYGPkCC7etHe/OeDKsTmt6fh3ALW8aWl6kP9erf
kj23DYO7uUFQPfjpAmH5muwxptg7wb3eGb3bS7sjaGKhsJ2/pywiLGxpAWxRLWHYy1ptVmhaVeOA
CGBR7MCpnvPw5DG5LVicT95oHLXkQ+S2Af+YtzUJQVAasddvF+5VwkFIcNEau7oklKQIVPuJsotd
4wYOkV6x9FzDWxJNXpE05EyDFVvTSl9+PT2XtFCE+tQrH3VR+gyYB+b66TSK4DEHSHCosihLH8CO
N8vBL6plpq7Fv+PkrUcQksBcbm8etvzLRKQjha1c8EsocF58MnqRJASCuZlAoQSZ8Zdujft3UrpF
7rRxbQBqORA0OBFOIKr6aYpSr2M9gFOtTQfzUgByTKzf78xaGdK769N0nX56FmGuZ/6aWmRq5Fud
SUVY/YpToO3cxMl2Gu8fmu5nVOHP3yxUvK4/O/lsx5mstIus3SsmE8ctJkvHFljy+81d2gQOSQ0L
NfqG5uoO/1XtbnbLuTCM4pNk+zD9fFUs7XSeVOeO3sRytY44TiUjKV4rsaysViEOFVONb0aWkbrc
pKM84umPNTpxGXKDXCwDHMsFiYXdsWlclKSWyzlvxuxAHL8t0jCoJ312sXBzWRxO343K3NetawMr
sswDVjPoFb/rExmLIHlB4e5VEciLcAfPVPMkF4hF/yjGdYNA0qY8V2zCwNTK8518Vp1pf4rvmhq2
4fbwAyRmX13/JqrEzrd3/QTnHjt/d8+Q4NyPZgEc7jho8iDNVtzFZ2FvT+eSNsk6EttWGvFqAqVL
Iw/s1WmM+WCtc0KpxiTOyEJQWgy76UfT6nMAcNgLq5PcShhUXSJStKVm9tbCHaibwbf02nfh/60z
4Y6rN/bd0dmpIN2kBrSAUZQTsi97LLL8ko1X62pEJRaYCW3cx/Z7U8qHZ1TH7Gbls0t/oBdU0inG
IZrJmuqxzjxLEp5/vuFs2skhw3zuiEiYs/4P9gRlcn/NAg8ItbJI/j5IchfJOjqbNpajYMPCiyJ0
rZmzoS7Od75RqblnwewYvbIGIh2HfdP7hNR5lA1XLukOhLW4R4ZjsQT9sk4NjWAXBZyAGAKkqnd8
DaCgFCNNI6AkMLsGQl+SFKF/IjIUWTWV64XKIu/0prbi0LRS48wK84GDPJr1ywJneaiNNcjaHtgy
BxTHnkqSRhtcOvfmljNmM6CGGeVB/8i/IFi1JnIhUt8sG/6klLfmiIi6vj0/xrX6E/uzmaQWtIzM
TVshpJW2eG7WcMbRO40XuCFMRQcomcR7NSlSIOBahb3zcyoBhGaMXKsmROG842xZLQsLLaN3wQLQ
9UjuSQanJz8u9w6iQZl8FFubX49ffEH+1F5FXx+5au9tjw2FVFcns1uFES/XiqPXrLUw1nP0OXZ5
xnla4ImFXh0CbRvwSqi+atmp+QfQW3qdMnBiUotg6lxzqtQ9ElK95/JTP8OwGzRTCtu/sV+0RL9/
k8s0f441tIiALM8RZpDk1a7Mxi8dWiuW8tZl/xGQ+phb8lyg/CsURXoAulDegCmqzw2aXHu2YsZQ
JtAw+HZ9YYQAxouPajUiQpphlABNsed+jdvGs/ieD6HRiDIRrPDPJ+7IL7gKBJrY5c+WiK2ziKa7
pjpykE1KdeWbSGKVnB/VZnZlzzzyR/OLkuajoEwuRbiU6d98mhOAe1lEKgS944RbpMTv/SlektnP
IAeCuc0k9c/FP5JkgFF6GjRR1kgh7W2PNT7tc32FNLBq072crTZ6lApJfw2vlG3AUUhUhIyd+v9I
TZmYk9A0ROvJKLeD6Q/fqYH1XsfCKmymqfQe1q/anvhzBInDIAuZJLPM93qcPJGSEwjnWfzXnr6R
AMjvgAsPgdu+JEY+V0nVDa0D0ywtGIaSoKqdNmAnnTYTUM+ftqgqeUueK5dV6R5d3I6nUIC4Al4H
Db2Ih9YE5LpLxWMVn1QdWEhG7EoWjEqiFsBODOSD4puvpvq+nlCOtbqF95/oueQAfz/aRlCVDQDd
lf2xJfpm0tZe/rJmXRHZSDKkFYaE9D3HRrPX7gzSlsutsvJk/V08uAv9+wTi9sJRgsHFp+eqKk/V
XJ1+aeUIKA1zEW3EozLxPQaHxKUedfW+Amk0QkRaTGhYfHDnfCI0IA2TyArFBCYuz9vuuNKuf8Od
C4o/2QfgcO4Qw9C1q4VMd53SoB8HSw3dGCK/rpIhMGjDVVlXsLGzqG70tQkuaIQBsRS5IRoJSknD
ZhTv/KYDC1M0qcncvbo0QYolNyUvcrvs3IV7QaR5FaCeRIrDjMlu5DfXZOaE5JpXuR2g8gP4OsvT
db4aaK51iNg3Vicpt6UqFTP7M+6wZ8mr2EoHJ/XIUxNOTp/rRyO4V6wml5bZte3M3Heey4qMD6BD
F8rbRwEsHFfkAJQukI/StJe/SHs1L9OrT7er3m5oK7ZXQ/j5pm4TXLszQaDkF6tiFK238DECuXLq
l8GmxjR4X9swz9FDUfwaopd0rEiSkvw2KfpPNnkoH/yJ0o3CammAT1e0ycChpojGJJipBqq3uUqp
3f6adTP7/nyFJ8G9BL0huZukJBEaVwcPklp6remW9l1G3ne9yYTCxOMzolvnlTxCHaJaP0g4BGxT
yHKwlQl5fSGrjGaTtlDSDhkHcd4o+31GD+2xMzHEuaqfa9/CP6hZRREP5X05PX1yVLWbv0pCkLkv
RXjza5207LAQ4QGbkpIo4+qXe6JZ13H0jLprFVF5yHk8RqQgOYGg9tBjRHICYqQy5U3mhKzYhP9o
r3OP5flYkV27+u6r+yjr9L0We8wRhj83T/bLMnEZVQflM7g8L+wnlIqbIgnuZ121T5DiLKuA3WpU
Ys2OjFe3FHH/SNkEYRqXZfVgpilyV/KXc9aPhK2ICAzcoWccN+z8EkgD2F/p1gqFv2oFl9XmoCnB
3B+gZV4hHLoJhGs29q9xeWZ3E3ZrNGs2QJijUJCVdqdSmxQtAGSbqZwHeK6I0OQmmT3X2XskXEP6
RaXXZbkcCyJl3pfAyGKthoutAe9Urv6Dt0whXSI9rEEei5ZcXlsbCpSsT1ANfHZWskXp5gK/txOY
FT30DeBRDsiy6VhToWqHsB6Z3WwQ79RDUq35Ca4XC94BObHQT+A8UCwwFbP9NL240hfANjkfkUt4
eUKKwbFlUADCfOwMNKwVkI3TA+w1Z+yF5FgXdXySavvl2NxLcXJDhVHFZdiMmQJZ5TPMI10t8toI
FzKgp/EaMiWEZtECRT89pVUounhLQDRs99EKrqdOaknlGYJHu1T0sKASi2XSI4bfcqwcr7IUockn
uBD5qRh1wfHJeDdRutpsPv5KQnhS5szaQMi5cfojb0sU3dwl9fQz8qQlU+k1gKH8dtOZID+H80Do
FAKYZOJY7d9KBPy8zRKkY4FrplOE4arEHK505UpS/WYLpzwWZWMOHYEYZ6/BzvzWdJwBh9ijxEpd
FMYJ9wN8XtcUuB7coW/u2cGsq26ZRN2QLPZpSg56qXbBhTV8Pj3t2qMuITSYpwlIfWTVbhLvH10a
zEZW4sLqAu4gLYLAyH1k9/w15MDFpsCaRhghFPHvrko+Y26lb29kIgRhjwQkrZs5Z8GbWgWQOg4e
UuJOUGK/yY3zYzxtGuBwWo38dBaWudgEuCetfRtaIFoEjjARjnH6kX7umbQXol4qzo5BWoj8ibv9
lkeLYprbq1WylwntBwxWpfqCM6VhJDxeobwe02o5s3M4o0ndClB0ws10IGMV4ZVFyEsjOQpgORIZ
ag8zcDhPXU9GKvYyD1arQIPj+vnx0WWlDpJ4mfDSAUF1sbmsOCBjAu017tn7OBrZK3ou7XNKSAAd
Ux9ccqUraZiWOutCmqLGvj4l14+2umt64ZBagwLUV3rH1wC2jc6MgM2z+AG0AgXO2lsAeKsJRJoZ
D/3wFumf5RLUwocs1iU3247vfBeyekmqVOw0psCp8RHP0S/VYAEWXbxvuxvegHxTfULb9rSp7E3q
wDFZyYlfFu1t9HEvn/2plmSbhlRG/bClGTeBRnRqeM5ETypQpUhqtJulArpsFcW5ydF87uNV4wPO
hBSxVpt54EoHlSrxpAsh2zHBbyUjoH6NZpSWlyELiZkwvq8BsuNLsvAGuf2IQ37a/tfXcWP5mm9V
pcwrW88sLVM+GavLpEZ+bJKI45UKkfuPYcZExSJvUlbJIAhHtp32C9kVyiQx8pYdSpQMR1z3PXXy
648ntUPwSoUZl0ObL5nMgvry7H2GONJwzxZBi1UX2zchXkbG29jZXkWMUZYsEOi5aQP9NuZSdYdf
jzIoK1aVyMAyouzsvK/N8ewsPoEu8N+z8XjXSMlFBs9K1wGBBvtyVJVTxga7sUQjdierhpSiY0D7
JML1MWMURKY7YuCOr9ENtrIan8uTmKcMA8mq31kavAVYp7vsxFzK4I0OWcEuTv/H8Y8DeXiCgPs1
I2Xe2/JvPSup58UUVLAue814aP7bMzgGrgv47dn/mOHpBwXxsas5lYaNsWHtimpA+1KMRXKhB5iB
qTgSqWs8QzksafiYIuV1gV4s+mUBjIQtncojIF68SU0+bmCqdey0JOpZ6LMzOEGatKzCYkvETxe2
SQ2sUfY3lCiJxpVlMet2Zz8utOraSteG8YpzlTVRYpQO/HQsyC7qQAQfApZePOOvepAb3fzXaRf4
kR468fNTyoSxp8GXm3tennaT9Ikf7StUe7+zaMLAykU3i/4tzeAXMMM+nSIgBsn1N+uHL+ylepKB
ZO1bFkdzvDdJELZbrHLwFcxPh5J5xz0ikmcGrgU2Zd9Vn2WohcxpLZMQgCYZ1423gV7+8ru8tm2+
rwqAeJIhoJBrQYsgQeyuJpTGiuMEOMi8dGWUIVd5OSFl9VDBx9gocjPlA+VxCm6XEjcNASf5xj6v
Vs4CFEJUcWxWfFpk70UEX28EsDdzZiCmpGEUVWmZTGdKqFdOhiZaM5mhvM0zY+1b3dzM/T0ViWCk
sODu0yoWeCm85vh1foRkyq3SGgMjuVt0IHnIYrXiJU0zV4h2H83b1CNB7IdYNO8O9JSh/UfPf0NF
NNCfSgK4CFj+sSxHP36AzA8IPJSsbxrJk0zWZxr9bpHR3cJiUC2hbvImF54Fi+gdyh/Z9ue8jUD2
F9h0+rvtaznyUeuCIxSf0DyxlrlrL6+lnRaWlKNLhGYtubZktVSAjk/3dP4RpoF4Fthiw9t97j9j
Y4/JE23Vfut/wk/wnA/kRv5oxpS21FsHaC+ky2YqlCCYmXhc2zH5eRQMMUqUNryZo8BdvvbbUzIP
pGmF9fQ4lJVGVbLmAHIIoQYQOnzIqkAWxwSgQYrYwbzFN64nqlVCK4wR+G6Zukxk8Me385SlJ2WK
uCOO4N3UcgDPbtVGWO3CtQERbO5ARJzsjVwmUqic0csU+8SNIgvg5UUFs5ryiKWRa0t/710C8b8K
ZHlQo56MetWaRPQb6rrA5+ES4QiCkz+u/HUZ+AAtdEZCXa8V9Qs3E5bv0EBz1s90RAHX6DeBbcY3
S4TrIRnTcaiPMNNfhWw1HDTFFxLw+f2ihjuE3WZTjBcZQlCiRiXqGGXbR8DDV1NO1KeHTM6cPWbD
/eRpQz9TVcOto4oUotmujmDOnhkkHI/xgM8LIq0cWmNwHu2CMZRXH8744jrCl1YXK91F/9QIIE/s
fHzWaBUSIL6YifJN3RpZ5bKkRjgJVKtiB7OpY/ol6eeHo4Buv6uSg9Pli7ZBEHIep5vlCQQvRvsk
x72CcOnb6LIduVcEDznjxlXlNAUGT6x0Ms3xj18C5BJZ5/Q9GZIbJVYSP9cJOnmJpcCIeACT1e7L
8RFZFs+ie85VcuIaFvqonrp5qTmoyT7KYQSS1hPk0z/jqWzEB7czyTi8tazl9gMIOTHw8pvgURFc
yWmuj7K8kQ8N0s1Ukz/BMKwlyCpA4kBUeFNX1uguafE7as+T8Oj8JswkN30X5GU4Bw7wFPy2bTgV
gPGmgoo1g05jnMec/9KgV5Hy+LcN8mujZt0onMkCVce2tj12dStSm8U4BmLeUdxtKY/okaSxTRdp
sWFXM+0Ay82m3xf/x/TKPJ1ABwoleT5NRoAbzRS3IFvaTLQ4wNLDH/dnzkOEYhSo3jppPAJjHkFo
SwmI4EQYA8QshDFsyk/OQ6yK+Xk1kQoJp868cNT4gp1Ie8IKAjIPw4AlwI5MdxxjJIRyQIK/uVtP
DXtZR0XGvv4hhE9HBmpkurq8zITfjcG7SyYtqWB2f0fySJtr37YtFp5O4ZLnKrDv7OZB2vhErYjd
EoLawOWmexbuCiXsVAp9In2WXQKEDEauxiJDa3hQmIvDunlw6JSAjaGJa94KB/dr+uJWRQmgaOOc
lOY6uTEJcY/Uo/441XYub7eUH8qFwo0LFPxKlKqThc0YGCp+H4URw7xzmfA8biLWqvp+G5ass5nP
DhT6opKYqsI2CODR2eZOfM+jZiw+pP17EAUEI2Sa0hWsZNc2giblPv/fjyVgciEJDU+HCGKGinaR
nrIYLg7Wc/cnzRxJ7Jv7DaeicctnqL3SmlHXGHs8LSKEGPAKekiau03Tp9t1vIYQZ1MZRD3mdM4C
GMRkWDz+XyYzNAKfIx9mt19L+uJL3UcE/zbQEQ9k1UU9X3PkD/TNqjWiy1L5OlQ/UYZbqZl4y3Af
64FslyUGckPQCrD7Cr0vCAZi/hcAtXRYKogVn/kSEBy1G3pF4TSK++bZZ+sozhu3O41A4Fl3Dxmt
I4nu97rn15bGoST7G1DHrMgQVEpmaIISfvSZGQ+7nZQWHFDXrt4X5R+1iM7I9nodpff4iDYdylaT
UeHPC7fEYhIDi9HMi9F3Lq1xb79PZMTD0an5a7/cSkVaZi9RyAMJ8BzvXHxXInLz92dWUg49FEqB
nam8EUzyJvOhWb+y3tugRXy25RjaEgPPBrYeBgwMmqkDq/jpdHKv+BXYfYH/73Ad+yva+QWlmelW
EpKrj/+x5BNWZ+WUUXNChYjHhjABqY9M/gTdESnAVqKXzlsxcXqFvCpFR89XfG2qc+0vvRsnzzfA
z/ix/0k4CWtWlOpiMY8nKXbMaL9b7uepDvppJSs+WtAbMwUkKoN7mL4+lTQwH5WWZEzodCvNt02s
Z0hWBfCY2uoc1b5d491KDUL+DJyPn/rOGv/tpqZSHpJOru4LVWLy+2HTwO/aW728/WgeVqwWTo6N
qtIgAKYhLuPfn2jm5kIkWQAaxi768GnSARUCLD+3Ox0Qy0pj8MLx4Z7ph/C11Sbo3X3E7pabI4dv
MN5zOvI5ea5v9XWWnV/SJEd8omGy4zn9l8I3qpYN4osh90cDglOWcNy4Hwc7fvLpXcH5eOLsP2Qd
ufcNCw7qcrHtUdpSkhhWOOq2IjT4uouSdyAMbAwg+RvMIg87SDp2ShzKrReTZ0T8iAlIPAkuIoEf
979OGE/Nqam0qHnFRsQ/P3qIROrJdFZpJ2ANS17+BhgU5bRBkVTCCx3Wxo3CxORX6xhnQQP7tLTP
JgxV1J26vKi+A/IFcBqNU5NPHxJsF1Yz+JyxT4SRJpb7tP6dE+SBAA6K1eHV72UwB1Ow6L7A7YaS
RLtK92otST7K2E9x3zsnmaMRl2TodfW5t6UBsZ4D9XN1PXGKVwLgqFmhtl9N4yuUxOnSYd0v4ZOb
xJotkrXn3ZuwWJiZ6PhJ3LiWIIlDF4anfKaJ97Zr3PXWyn3/ar9xjyt4bxCQy8Ti4mCzS6xbIpgq
d00QAryjs2d2TrXg5A/bCmlv5OvJc5EY5tNz2huGF07EVgVBouJDNhIOLB7QE2RGD8CED+F+T7Wj
hBfAB2NDtngWGOnxDcJp+fBpAJpa1K1nSrvYQmHNGO7RPfXV3T1gA7c37t3Gdr/aJ/koGZlPX5t2
OPySya88oQ+coLV7FAM9l16NQ0hba2ysJCiHeq8qeblRXKTDUc3JIT9cYPns3Y6re01Ub72kShZs
995oUxw+7ftu46CHWulJgFBH158RbF3DMTSYHbHQ9U4HeURRJfunCR88uCe2GDLIbgVQNyyx0sbD
UDcCu20ss2NL6n2ImktLN8PrS02E+cMKb9X/xIpUJ6WcdHmfNH9/M+wgT5lxWqxMS48VVjwdneO2
eqbK21+igYkxj8NSuzMqtc6+p3daQQ0ru+J9K6HV0fFm10nyZaLck325pCjGjjwT85pA7gXVDfsa
TEXBKP/mSZw2iMOR9s3cgM1LkKdU6Voxqql2AuwZ6/iIS24k1aSj3oWUn9N4cDMMuCcoFcnGKooa
gvJKteiUCrzPmMBoiHUS4NZpncr2/00pXWWBFa/Ia7l78zoAgu1LX3HWDiNuwEZJ0AJDZwSXLtlh
Y3zop8IUTw3MbJPN75OcvSoLIvX8j3/hJz7OqS0J2pItsRxD79ztGX7Jt46SVIyTYEXULwwRMYmz
xAjqdpg2Hw0xJNYe5tk4IsRfQk5Zf8ABhZlaFzTWHXadKaE948jFLAjQNGVe/qecYAnst4NlxblA
+vuQkTHQ7TEPizEOKrpKdiGeyGO3En6+XJPaqy01d/hSBJwA/0mNUlPKPBkYphpSRcz3RikURLPp
RwiKuQodBLm2UTuYSQj9Ag9SNJgasXnwUMpipfrfoQDwvH4R1mbOWIiwX/vVmG0xkUSid/qiLqRW
fb6RZRb5k6N0+kkePS0Yr/Y9LwOJ1RqiLCwsPTCrc5jd5Kz+Zx+Op4uHytARXARxjtEcBxPLtGZq
pHtkz78AqT7Ie3ZjgDqlaX8AogC83LHWHpPkNAnmVvxJFtUoQt3YHCpJv8wyESDp5+CzJhQ0Rxna
temzkI60L3+r/Y0fRexFh4ogAIqXn1cZTbahmffsPM2NE5hCibP3vQmKh7EWtbDIF7OCJIJS/5pA
QE9kNvjz0ZcaqXTUfhnLMYfY65BdCxgn67q86eb15f0uMU1JYkWTuPmwk/8nf6zIWblU5Fzm2zcw
jOA8Rl8j6mlOixlAn4RzdShNqsP1fckFGHrdeFg5WsS275t34XjY3D8NDOF2uDYaTTgJJaoXOCX3
2JjzykKOtrAXvULjnsxrlllF0YaWH5W8Js7n7YMmG6pX7YqgJnB59icgnMhZuYgpzx+zhcmYoFCj
pJ+gUlcqGmCEszstdD8KFkK/RVS5J9AGx9lNvl2RzpKzoCIVHIeHJc1M9ZbqEoASRr6nChAxaJD4
52IcwmdTM0Lw8W4bx3lSgpNMOVcIGVpR1DXhJekjygmTAFy7vkPZ/8XecUHZKnhe3p6XP4HHkQHF
3+uP/a5e73Dh2dm0FkqbcaQjauDXHQynyKBRH+2MtKds53lD9HFv8ZXA9Ls878YGeqRwx4GEoMKh
vxvjgUrFrTB+hqOOGeNkQMztUad1VHqdQ97ZaiRASC9xVW+RtHpvQf1T23XzzL4nKxMDXmywg29P
Bib+AqVlAp0U3eZkABUa2mV+SUPALgx5qQ+k1pQoWaZfjCQ57vx/ELo5oeSePQCStgdH2WBtuVQ0
txyoeLNcQYVBDup8YFvqdTJSn/w3v+DZ+nSDpai0nvWZsV4Dby4vZzz4YK1iLe2McRQZWl8tkdkz
1/7UTofiKRJsfYQNDTmUcCSPuNgTNXHPrSKGUcY6P7ni+u4YFz0u0C9s9E3iAl+AlZnNU0MfFgsi
gaYQOS/9v46vvz4mMN58S32dDBH9+d5BoCDzlEcZakaG+9VcwU9RZ1QD79p82mcODJNtfyHWrF4z
ljBSm6eZrijhtO/bZM9T3v42Lia56N/n7WEl9yBA0NjZiYBnY29qv/XShK9SNf0rXmMEgWFSzl6c
cd8HDQcKM4Rjeza5OWKTfZ2FzpT2yFa7fdchcNoWlfqrdjfyXnRgFEWUnms/t75VsR5CvWSD4Z0T
jmnPraBxCO9LMnueRDBjV9FMx86Bvm4v9RDts1v+ufIhDw2EC1wGTsSPaY7dxBJ/AHSb2akB1VZ7
/jSbJbkaG3Am1BnFyyx0SDsU735bLhiLxFLpOmbsPV0/GyCX64tD2l53OZhHi0Bm9tetPMi8WYCD
AU+cp0cMn0RKGotzb+vEtRvnfry/5/W94RsKQLwbHe3JMknGA7BEGs3nHkVty3VYRXYowwmCY4FU
l2SeT7lqTWKZeOKD0sYhI3Tfrk3DDnjwWNN65wghP4Kri9JTlbt2GIvadn/rO5UkV2XKiP1sxkrl
BcfXI3eNJ/xCI6GRqdvrk0BnQ1NrJxG6iv3PTa1OsDUeqc3rX3JkEZ+68GvFtfO5ERhjDiyyN6uC
n7DhMGBg38D3d7z/H/aftRFGdhmZOekaAYO2RGs/jrdQbqtKMJJPbxZ6dK/sUm59E/q5HfM4lxns
B+cCYPUaoBxYRThil4q469GdtB1eIk0sHH9JzvYCCnsY3P3tI7NodJw/qjzD942UJ3XpM1Aeq6B4
SZZk+w44edYiGj4fuP4gAqT1h831c6A3l1Gny32Me9pjH9quCyL3OOA0BpPPI93enhvDJMpzLxoz
D4WI34tvvO3VdWQuLDNthxQ/D8gEENI6ejrsXg8ssRVf9LWd5JXoWdlIwRcAtRra2DVD+dcTrrlP
iltEoAGH4mG65dvu3hKRj8BSUDclwxmrixAKbAj9Z2G3ZTnmUybQTAn09O35CpN7QdRwsxfMLSMr
DiFenG3o/NeIVW/Hb0bdsHyQzkk+M9GGhyoTKCyPUkkVxo2fecQ+LY/d2CIT2UUl6TKvuppT4EC3
+VKz0XQURrl9mpSI0g7AtJ17nu/eJNmScggwj82LzN5L4H/IhASf49GniDxACUVrjCl/FSwm4SWL
LwFS1aXo56lEAMbpRZ2HVFYEX9cgxxMi8dfoWdrtMhvDWCcxylyCvM6Yh7XGmALJVut1x0UYFgYc
m00r0Szg+s7Ywe+fX5BwyaMB6p8HHjlPdyy0b0Rkt5V7vG95PxSb/RqJc+Jbam1aKLvtEyU4w0t3
XjP0MnmueJRFSx7AIKeewzwpYvu3OO4zswpihu+ETstH3yBpmrOHs5Ic4O5K9SQ0xKsClclxj3rx
cLfbbMWPFWxZMk9ydi+9G3OMFSz24CnQwqzyklYc63IiROKSGyD3qmFCNsVWCUPGSm4vO+IsFqV0
M3rJElj/eGvtwiW71TOpo+QM2TvOzY3RXl2X1dg1R1oVvhFWi7y5zP28F4G6kujDFEkeFhsaD7rw
u9kvFBNy6Ve2MDVKDv7r05Hb2fJgjwx3XGyo1/4BtWRmA8Zrx1BBtIxDESvfVDumma1oc2csm8I9
RXMnQTJR/ModkfPq7hMq2RPhrafQy+RYGezNKeoL97oXyIeRTFeiYZZcRS90xHjK6T+pT47+XWHJ
lAhjh62z3QLyo6Q2L4Ib4fNgNA2Xx/IKUeZ85qYzojXAxkb2RDjYQ+DfdZSCpD6wu8vc43irSsn0
8SXYLamhGgdjXHhSE6dutGE2TNEmGLwSTn0yUKz/WtCJDDp00mLbz6cVhvFlTbjb5yAFauri2N58
q0xcirWkUi1B/0VULR9DkqIyhEHqURcXLMebtyZVQA+9asOX/6gCDDH9JDb2yA6jB1+q/oDfyL+b
K9xILYk7iB639V7hi1OPbsZeleqklNh9U9mhFvkyVOLCagzEsUU1AS/Uh4jWlX6/XIWef/HUUYcc
sJnX+tpbHo7F4eTa2bevVuTKhsvnfHOE25BywxabmGDws7soibE9ouI+aTbJiNf+q5GMrRCEj0i8
Vpg8/WnVE3kBkOqyIdksR9Qxw+wM0Fr//Wa1VjaHoeFBGMbm29Ij/2RYoB8efUupbg6onM6+gHBI
Y5MAsL6/HH0gwT8PtFt2AP8JH1v8mecB5hdLvHAN6VYMDNkFa1cjU4KOmC0Rm34dusHbJvHStpfy
8+hj1uy0Xkj8gmSMwQFmCjXqDT4EnUXtZkCC1IA8ajg1BzHxf76ZVMQIcQ3A/UQodt0K/rOlapoO
Temv/5kd9Sk4Un2akG1+jYtNukrYWKJic6GcU5G0+KxD2xctCxgvmoXVFLweHugGnDjccxpJgUqW
uEiBJQ9bLUE+vXLhrP2fqyGc6ws7RuqLI3RtjFYIudFe6nepdBCTLEeuZQcW8a3CsdxV5qpy4rjH
uEMwsnPqu8Q8cHlT15GRtes8aesWffgW56AoisM+5fLEf0vEBwWuhvCwpIN9EP3E/+EtDD/5RvIK
HI7wJweZVfboCOcxJZDFA5FRYgZK2z7k0EHvhNameaI6qhi+mUWokunbSBYbzqLCZX1DnXXsQwm0
yDD9HAmMZEAYSoVW1u3C2SjSvfFEsS/xwKGO/9wPwWsyJBMWr3CafJdu51Xkbiq1RjKrmos+f14k
4gysLARDLxDD5vQ31U02Bf4G4VDA37boldn3fV0wWePgj60P/kWOlf/r7QOmaXFBTjJ8v1oOzCP9
pXY3hZC/K8mb2J0IRBWTYleGyICOG4jY5AUBCKZeB7yWQqkm8/7KR+ReGrUeHz3r1+Ogh0wCkzdc
ZADwOZ5T877axax8AAX7f/MRzEr2m/TBnOmsbUpB8hac7LpP4ueStfJEmxYK1I6MwVf0TaaoDRas
en0Cg+4xrYjZI3dfNY8gwGf7AqJLyazZ5HL7lPA0qI2gfTlQdsdU7oHsYHD09yVpgWPN9bg1ZN6g
4x3wMwV2BVK3uvpmZytC+RFgDzRV6x3gX067GGN4kfxn1vBaqoJKNhzzaVMR3vcuFQdRj4EP76u9
pR2sZVO7NnHRSbVIvBrtb2S+hixaWW6iscLORuW5fcYp04ZRn3SPU3EFNlehwhxtlgzrUKzOjwMD
JsSCwx+MLizVa66oWP5caWYH8BwTYaqOH/gVZ5BZ+r+jvt18A72VQyg00ZDWSmwFJdEt9ySuKPP0
kkQpnvqC2xfT7994+gHHsWJZwXs8bmWPn1RbN5TrXUqpA/wIOGH3F/xj4997r14cvsy8SPdDn6pL
mJGzhd+xqF53zuBofy0wYDnafYZPg+rRl6VyU4lNRf40OMx6ZAaCg0HHcFE4GthHdIi6tVp+XLcQ
rsiOfrNjMIweoIO7Grw58VPnMnIPKoSZkc41PxkXZnMm+SKzZTPODDd/KJHiltFBBXQ7UwxTGx9A
yry5wZ8akAD/OFyh0y3sKFOk1PtY5IGdnRL5Dj6rDSo5aDA8d/fW5YnBlVG5iTLMqUrgVS4XK6VW
1Mf6QGBj8W6knEy5rOtj/+Jr3OOAlldCI6LaEDjTcXc7LebJ3szjK2bChLY1uTm7ohM08wzAjAl+
k4Qxqq6zB9XbVydk6zpfoS5G/htTE1oW+EQIduYxJVZFralRkfB27pb/HjSyiKT/8FA1EuHccu+/
iIJT2BFrJ/GP2EW3PnGyCUaUxpekrzwhpjs5o1YLtJ+m1mBZxcdgO063xT5pTEojnOCV0cNw7TyK
PkEYXEXs6N7IFQ7hcy8Pu2tCaRawF4TaVGqOtwWFL4PAhQFpZ3i2OhIMcGWnYjQmBypxpKRcnlfC
kuV15aYcCefLpfK1qTNUQwSEA3ozkvFy7piOeF066D4s34Vr5mopF5lcvJ/Zn6s/J7zEMWS/oPo2
Y2dY8PzCYsJrA4sRhwAxTyvHWcbl9viZ3wiZslgMpUzS2N+hPRpZjOE4vS+Nr7J2JCUehtkO5ftz
F6x8p6/mxEW7CCKK6PKgXhuiakE/ye+JbmIm2RMV4com6LXOnOGnEqRoBXj0Q8D/h0GiiwheX5Ql
nXmsYN/RCq/JJoikPuCmarKEGqDr7mhC/naJSF7FVZZ+eOKfmIsZ5n5e3h/BpEkQ+QZAWZ9jGX/g
EuZ6zanWasgDOSxY6fq2Un+m5iaMLh/JZq/6kFxG+LZv+vmjNqHF7kvC0suOZATOyF4t88WoFHJy
jp2qCLQmWOG8M7GMy3iXAnYtFalbfPGAcjzhlkxMO9PQLVFn/nMA/cKjBw8kCxV2J4HQJGw4pdEj
v32SV045XuosmlOs7uK5HDUfyIn54vOZq2/cfaCBlmgNVK0DTIcoW9ECzH1cjEv0hNVCMcrmK6j2
aah58CteuC/TVyNnfbMQ18Q36l5PN2ojFZSye/GVf2oc+auJ8ickxzGXYwufSsNwlFDlN3529xeY
FxuVFOR/7KzTW7bimvVOIZghZbAav2sXgYoiPFcqcI3pgZzMQ4pDcvLuEfMOjCwKJnNiip8zbitI
dZCvqHY2gKNt78VWBaGWC03/xlPOReejfr80KD1FcFpAk3Xk6zcZT2n95tiKmWMp5P1w5JTAgf2V
ZBDTaISOrYxTy7o5LSyWBT9DU+F9ELhiEwCx4PoHk7xa8SMB+MvRWunorJVI3jbQhpbEJVosUCqm
u1u6WrdNUiee26gnjdSUa+YshAIkN8UK8jDnn5EF/zNo0pjdsXdjD5W/mOWhbjo8atM5yW3SY6Pf
U9TOP7F/dbAMOgluWD1/FrCzTE0tM5D/3V3DvxmTxxLB+AodvGdnUoMQyGuaDUPrg6EGveXGg/OT
Y44q0YbW9XWfIliP9IYeBSQ6KmVhmpQgeID18vJFGkC9qQKWsBmg+5ws7e0ZfEbF/8bVIpZzXId/
iQgUJjFLUia1QARimOJyeFrHgC/EwrHO0IKR04n6XP4ZGbZqLdQ3B4Rdi3WrG20xVwylyrZQvobv
iCM+YEcRP5VkuO6O6lPmbaPoIjqOI1Z3zUcv0YpepIXde8kZQltTp1EC3Gj6umgESs1fq9GvQzLK
FBDCA4n97wIgZ57FsJjbZMskyyB+1Ni7xbASrZgaRBSZ0I0scIbbh6NsTshtmvxFyujShnRK1S4o
no7Bt7XeZddiSKz/BkzTXpvHZVLVpdq5NeAqlLDG96XQADZN1bc/O0E/j7H5atfQ0DiDL6wdzWsd
wK5/evDU4soqEuug98y0O5+/lbF/tq10BGHPtCbxbYfY2fogww1BykH2HUKevET7YEluxIOcJyI+
Qx9DgCU3Vbu3/IBGnMBjT9sMhYbAndEw1scaiAICKTjngo/uSZQ1qEnWUUGJ/AIJKTVMWi36wqNE
J15Gxt2aLfmzZK3V72GDbTmvHEOoQLh3Yh6W1lMnKqLJyPu7CRguz672fXpR/7xRFI9v6+lZ4t+m
gN4jIhwpnHNpi/CzV7crRyhVVFBWYFC6vb+hd27d0dWOQ54TGF4PJPz9G3MrKNHhqYfuV700qlNt
X/qY+68YZWIxg4x617y/60hfq1BWU6MEpcTFPV+ztvOdCSIliy1dt45ONeRrGG419fHyv6K/G/Ir
c6x5IKaQL+Ai3+kVuBe1zMEb/RPorIm1jWcckPlFxZ1wExEXZI9BhkEBoAJhhYEa2N2FGSkWKaUp
EVGGLS0L6E4Apy2WF/wyf1yZEDtTfS5L902CZbyRyEkHQrJhRBh2+ti8EdaWtAGTXBoo/FTt10nG
UQrKZZIdiLeqKno1h0cBCr6RqvR8T8El/qPP9kCeAOc3n+g5tcD4G1PVcNVs7rJNGeo6n6Kp420K
r+huu/QeQl5zuCViPAidQXK9i0UYtbz1ptjUwb0kQILsaJe/zV3nf0RlChdHzuRwLyqGRfL6ouz3
CUjsGvtvFTf7MTnLCqiKkDycsPSq/82h0yzzxb683F4OO9vHkOLvf913EJ0a23E+VMSSQUR82Mm+
vIo9yof+5JsxknqQaUTQMcpEO5/QcbcxFXmsZzY9vzngsPuE21xsr5qkJ1zJMezP/anvQIHmD45f
2+KoY+XU3bv3n67kDDhbbtK7FGepCSvmbHlVxksxFwyF0MZ67REHl496EGbyzvMGOvCssRTIlkyN
BcWqW77bsQEZ2C1dUuqqE21I+3xlGgRB4SuZNh4Q5+Ezh9vbPF0dXwSvGg8Ia5LAhwOhf63ls+mP
zUlKgJv8PXGcjlYYIHNEsRu07jVD9zvKto0XoXdyKaKOFjq/vtg728pU+8cQBBsRj54NXSKjO//0
njp0JPVu012ZfFfwuN31LwDpg6PSBVtL9+6MHWCpC6GoEyJH03nujjpyD/2E/t/I+lJrJTeXVc4g
P6YbDJZLQycMV++ogPE7DE5q3RhiXkmZDQ9pTavk+flTwyrYr+GpcrItstwSSGzoicEmHwbx+FUe
/6+KSddJD39Jy2udG5oV1Zj9DypSI4LQHDz3CPmLM794/m1tTQfd1LY5ruRn0p02QRDr2UhR80SB
17bS6xxRRdK6b0Ow/fyHVuEx1Ay597MKxw7bM0meXxgxXTZp1SZBU1BGk95SKaC2dbM8JCJOlWdx
UpGO7Mry2bQEweWblqjBgqVZTA8XpvbwkDAbGLC/bN5F2v1OV/K3c9WhN/Zu10BM+FI8xfj1dNNO
zBx6QMIagXX4/ZXmVXITgaQQZu88WSjDkfoaWvb2MFwx2FUknCtLJ/NClebBq49hZXjrUbuD44CC
gRQPgxCO7CYhOOp/qn0x/3cbRNm3by37mmeKYmqwjplkoCOERSsk3h1GjbcsdKnQOC8JPHLOPFtb
ddZs9Ldk0Du4Wg5r+cmlO0/UrAatSO83669ALDNCVFEZkf1yqW6NkCXk4c5G7rDqG6tLX9mySJMe
43hQ8Kiz8Qp3OaegueA1VL55D7cOVqkB4ayIgHQGNpmwk63sxAKzWMuqvCgcecCH3NMeARAh6NHe
f/0ZfCPVah85yGqo238JzPQ/OgZW/shi6X6Ux1uQ5xyMtZiUsguO/kdslfwxlPzMpTk8KetXUm14
78mohnDQaUs46SV3xofG4l6mBD3VyjA3a1pXyVY8siW3HygmolwV+fw4lPjYvWhE8o+X2ZP9mRdT
BOiNqzMpO3qUxI7IdwZ07oT8sXAzCNdhFsZ4mDIpPXsYiM3ZgRove0KB2GhvL+oD7ueNo1dT9ihy
51ck22g+liWeGVtg1HckfuwyovH4UqQUz1WLjYMKhqyBFb17VST1cprrY5py1J8MQPtmsv3vAxPh
bbpANzhQB6tznxWO0bo0FfZVBVnPhpVi4jgNaG51g8QD1e9mDUoibDGPG1Wyg9ulmtiuVJsBWzl9
+q4L2hMvwDUiO77m8xNUn/P4llMrx6x8Oz5klil4o8EkBzjpofI4/nnFHGSOr22Z8cGDgt37jz4Y
wsyWq9mG9NwAVWFVXxEyBiFprsk1rZ+A0aA4XjMZCbDhUZhlu9yjDOLNXiscxssV8aMwN24q+iaW
sP3NFgpmuyVYhjt+0y9jjU1auE/TDESbNeVfy38WKwPLb4s5y5aUPOWNGMI/JfXs1mXKCTYiEVo/
gPcyaKXPQ2quF1Sno5jryonxd3lPwe2FHFH2wFn9QsFs8qQzrUGthS80F3CpgL/fstcBQBTXTplW
lfIksE09dQFrCP6O6+n8mC6cIoMg/Hd7u/o0dVD3ZcScf8m+24hePuCCn/5OxbxQfXYLRZD6lgyp
ImMg8agUv/orsDVOLQbRMEXNjuXYCRf/iKM83G9zteOo40UI9tsPmZfg4j9Rs5NU2w6Nj55R46Yr
nnqqadaRXK5OMP5uc5TIep/EWPV0ynH0aNxC22W08mmg21QsLWU5JHLtSzZ1mJhtgrwZ9fg+1Mgb
G6SbG1fvuyXIexQWgsm6D9ibdiRiUgyOIT4u4uiBxqxlu1xMYWaei5LtPjWLFQABeu/gIHABl0zw
DQs36F6kRpStgLsl9jy/7PquoG5Cf3mkMy7z+1A8jC9zCVt1NLoiTTFpeFu68vnPb6UGCAs1zi6S
aQhUCJhTyOT90ZExosnSd/qewCi0oSAaHkol+5nVzaAI6E6Fc1RAbaXXAUCYmzv8PdBqJFQvJON6
0dxbix+CZmYpkks/ULNEc0vG87t+TonE91zxsFezYUMAZdMJWWH3eCvL+DFzUQB4PRTBLhRt7vAq
mS+pzwNXwDY7EokRkTh2j20vmdeLcQusK5GnSxHU6glt+IZVZHGsbLhZJ92OoyaWaBG5zbdYkldL
dyV7FEa3J7g1Rc3j3h50DhChEj8DIiwogeFtX0hw958E2mauc0Uk9RiHVQtMa1UmnP1fHK7mfsC8
Bbfg6nfqCr50gY6JXhKrlQyzyAdD2gaSoXyJoD/u6r5F3WZh1SyVdYogL2A6Ru78LfMU0kRL/w/L
iioSFfXXMazVJo8XZgfplQCYSQfMXgpUqV/KWFs6lzVl816hjW96dVwKkaBf/cGUOwPHXZhgPk4c
oXFLop+7zaCWLTrBQQnjCjIvQk3/kJKXSeATjbkjm0/NDfSLf8ytn66jxvWJ0hFeA02mBEmKYBJn
cnCyGb3D6j9NoJi7uQzdg6mGz4xm+4i22+poAEXUWUJs0U7ZQRqQzvwNGX8A9gwzKs64gLORHn1m
QinAOFcnN3gqAHcV9L0KDzXfX9w093mHx90sHjlM7WSTM2m62rJPgLSUqnEDozxuBF5GlE29eg6R
kwqdFciVTNn9EtteAUS0UNleBhB0KdTw9vrtrCiOw26mZv8tnRG6vY5vBJh0nl/ePB+A9fhZpJhH
jjbTB+NQelOO14eFTG5SA00hmQqnyPH/bLvhM+oAQU7WUVXKsALJHqcOs+i9dYaeMKYNXbzGuvTz
qHkvrAM7n8Pzon5gAQ4TMdMZZ6jPm2p0pk159WKrGksLhjQ5YNDpo4+HZz59YRJPrYs1yIkmNKp2
vjOXRgaCMSc1w5b9yY+ONI9EigdP6S0f97n6hcFBRSXm2UHP+d/RVI48oC1tNaqE5zXcoXA93+D/
kQikL75COgvfwREON+YPWOceK/pvJ67mOsnlF691o0wPlW03/Xhx7LlEnoR7xgvaBwqjbiBizfvU
KCTE1ccnsKMxP6rE3zwAkOMRiLj8RW8Eh+lTbt9dUovpIhs++wMklk5qRlHl/cqQMExDumFToZHg
A9GIqm2/BdjLjMbpf9RjwafKPABJiX9S5AZEq57gcOFC964PR12/TwGD485YyvkhlhzHqrPP29C2
ZZU9Bp7Af7ipoE/Qi+fyfk8jW3d9aDxTeTdWXu14YYvXa1wYb/H15L87ah77r+1cobPg1uDq963K
GGwL20C+0Ynv27+zQq9o4pAlIeeVgTP+JV/P5IoFvyFvR+zo0W+j7iWnkKNafaADpxF0lpyppS7Q
kqYzT8lbveTtR7jXqyxlbhG5mNbsx3OaXnvhqVll5pWSlb5mEalXSMtGhvvJ8VYoUyeFX4EuZ2Wo
mrou+C0b2avoawNClTySvAws0t9XixW4XZ4uiSFlsSnauraA50zCrTbltqnzTJaS4SAu6mJSGq7b
CMtWSOzBlumSNcovmcGXWx2+kFdhBgdSORQmyZ2O9AHFEPyWYtTiMJYyGtqOddDt86KH010AdmCZ
vozYlt0+pSW2Ea1lfzztKF7yjDk9lprTmnnZ1XRjevvO4VMah+lx/v6Pnfw8VPDdUGYCbummHy3C
7oZGopIse6WxBUb8fFYho/XoA00WbbHxitKSA44XMAIpBzP4+K0CUhYllXECnmwMhc/i905iyDn5
lbodIHuUGRIwFJ/1JN0D25E4UCVsojlHbbyBf93VcJGP2dnkpFOlqxWARMmAjONhl/3ZTrw4lVJw
DIelShK8V4hKgHPtGjP1QcV3sAlAdaF8i9VJGyvNBjQSmg4mYfrwwsiPFSGwKd9bzj49jl2fU9Gx
owISK6RocvsHW6KNL/V6PJi3155+v6VbGTVf24221o+D+xhTr5sKgZ0VA73aoFXzxuJFbxIOEeGF
qo+/aW5lRdVMF1O+f7M7Q/lADz4a6r5DcBGwYnY3WSJNSC+1Kat265Ui1guoeENmMA7jj4uxABr/
2EeQosBWiKMIJ9snWzTuMwUGjNPp/YO6r9eZRXWJiPw8bidQpN+EXeTU1Hk+sWIyCXc44RI5kTnz
bJ2bHsvWuRaXnFD0XpClF1VZgc0Zz29iRguslTRCyD3tGMlPSktAo17I3TiRkRWLp/nuNJ9mZeTO
jfVd5+S/xyDPJ0Fo9rOeGDSwUVuxhEYpzVR/FAw2g3FqZUI0ryytiE8WbpBGRJMHsnlrOX1dkHc1
Vim6iir6fOPzaz1kxkP7/Lkb6lxoRgYhJgGM8/qQq3vryA6tOMbJE/fiSpYnEQ8lR8CGdt791fRA
ojzRxJ2jBssvGytLpS6HWBEUbwKZO3nk9RviJdR9YiJ+5F4IJ6ka6iM9YQRf5mnBM9Muo2CHbGrb
OnApCGH5gx/gkke2rebw29rPfU5jE8xmE0QkBzExnhiJsX8M8b8WUKi8PeINMG2U1obcXl+eF4JK
P6VGN6mV8iEgh8htajtYD+mhnGLhfy4HvnU24Av152TKcDoLHYhTF1D9fDYGd9/cs9gUEGJV9NGd
cy1cEurgqbMZUMewUW7D/tQ5/WJMQp2k+JMB7vYGei6A6ylgPtvTHtM5jt7972NL4VPWnlVQfjP/
PA65d8yn2XOHp6M1BQHcRlmZQlvuZ9zTIWIE3D6pgNfvMwB/FyXMhyIiF+X4FvG1GIGvt0cOLxS0
6VMKdnQ9iElOM+o/ptw3S43oG84tSYFumND841e9+Vp+OjYFQas58DoH2GAInH1WnAE1djlJ6nDK
qa2ABgk2pxY8G4jioFVSYjtKLjWJr9OdlDT+EmBUE1KHPZiNGjcKPfpSa4Kcf8GnsEw9efX+RwbT
RfNrYDrVvfEE1n1XZHPf9DE3LJZvNlLVn4RxSmpOtRjDVYjvRqw3uPAGil9F0wuDCNqR0jmpLJ59
S7D9S+B5bvp7eh9SPP86xP1czY9yjFU615wxkFJqX+9wwpO8Q9vGipdCMs0es8HIQ5/aQhmqeHmo
uqZmde1fR/R4brQxwdh7aHQLD80ENCvVxwsj4HIfDYLTkknbbIILrW5vtMrZ4LruKdCWAOvdC39Z
o9nynV6VHnCvUbR5OcwOtFDRhau7FnXf894+htJwIU81p+bATS2LYi2WpJfHJmrrVgNI5vGSXX0p
AkvjU4mycdrlDaUv6ec+znkInsMDTgc8nVj6rSStUS04IYt6kXJ5IHZR2/3HwoV1QJWnSwbtzY0q
cNwXKPYtHFHYWKErUb1D1tkqWMWDURQX60e4xizpXEi9NNQekrPQrfsDgHibMW0Up0i9NK7/vjGI
MmzNfI1IpQtPjJGKHoGhSm4CmCnEwtZPNM+n55hYdimxpezwf2zOxqeY7e/G2IWjB7PPnBcWoN5j
uSjbIttJIQMdvqFB5HricXh0APmnlmgVuxTbLnoika2N9eyi4/WX62vyW8wrxwtGmhsh7lgbcOqM
ZfSDePmnMFmnvOXY64cXi2q27iLmtMoJ7I3u/0A3XT2GyQemcyvh6WukRgbQ828XXci79FaJBm91
YHnZLPRHEgDXXboNLNLzo2H7uUwiXJxlgEFwwbbI4tf1jZC/ot3xRL/R8UkbGJx5wPLLOdlEjb/M
ae3WxytuqJe3Ll/Ry4riAZJ03CWxHOQ/HDRnftlwaMMiJB2MZzMfzo1RWXCZNR8rT/Itgv/q9CAw
qaoxS+6tYf8zfOcdPR3mQAkRWN8IA8gDBjZZ2yxJisX8ZKz+r3h1nvC6p1q8Wj2OcrWXUKQcya4D
aZ6vpKG55DttEi96Cg/mzMeF3+s98NRoiKLWO0RbRtTAtsynb05rl+YKK+2FSxzv0LfXma3PwSbl
o80kM9tWGVSSN5n0h2K8zntWH0bfiyRO74hcN5SMC2Oqkv0ClyqxKbkdhzR7mF49FuvN7/h46lnv
9ZLkhDjVYLSmRI2hifZjU7CgyqxwFxwQCUfodMDBOCgqlRrI9jogSrwiWkRAHxUN9QKP7OoXsqBG
77LM8nIwfpYNa/9p/8Ru5+CBOWrwt4dAuVaqzHg0Ph28cte/u4Ae87laBRw1RRwgSwcSeuuecgcY
jxzOc6M8TH0bbxKUOsa0lWQQ7D0EUC486XoFqRzpWAq2T35+XHP9Q7+Oibo7y5LigIIzarGlFoo3
9Lf6bYvxrYdfKPraXvBSSWdYQJ4NKpNePmeMWJCoPHRMdWLLEy2DXsWPJOdOiIRRXvxqfAwHJbj+
fEvtbAVJI1S33ELYEqlew664htqMtLhQMf2LK/AfMDWOmIVBlCRYctoiv2bc0LKdoImZG07C/I5s
JsBfZW8iuIEoakH5Ix/7anskBNurnENTLNuL92Doj3x2p/WEx5AIRmzXTUCacUuS7lQBvQVScTUj
dPbPfJIbaiV2aTWI1oHQRQBLZiWg1EkXo+uvjPJXGHHDBtQIx97Z1kclxnuCkou9Hzkfh5LFYN6G
8HffTRSqq/FqmgUji0tgFg3ONb0kulhZDo1xxOLjMqkGdJWsNoSCrHRbiEvB+UqaOJA23YxYBobj
2Xf+hsNF4YmYjJWkOa9bHQXUHJP7cT1xE26VbYyTKK++sNM0WPLcErM1y9ewQ33YsIDK8l4A8ItP
dVhKGF1QPWlMACMr21CEJiOFstCwhMoqaldd03vxdVrJqs0P/dHLnhqOtZ9GMGuZ2yjDJ4ooHE9Y
P+r+keejyuvu2A5TPLIIjV9uJQbiDlafzt9fdC6hQ6szYczvZM+wyCHJhAWJLmeUcYxaKUNqNI09
H5yyzhPaU0geVyQK3UPGYZCkx+u2t8WGOfD8ucIKNleAdJmmazhs1wl1g39LMmyND/GdILV8yEV5
Vt3j8kd9J1WEztyz7QlCWVulspa9I4oRFPPqC7ow1Z5TGtye4LU7+c7k/Xuz6TpR4r4rhcyEMAjm
HLR6BFN5guWRHc3EjpoTLgXkXK1xc01RtrSo21smwFrN46mkoEuuHQ7MzoK38QoKsZgVTMHFGevE
ej9GuNDggHlU8M5q2Zx9My0lEhhAIL0Hu2jJzLLnw7ugOJcoZESrNdHvr+obsACbb7Fpi8hrlm9t
mzNXmweTAnH6eef42dJOCH9Nat1A/98Rj9UfoqIfy972lcdpPv1ppA7fX/rVopD4nTVh+Zo1/Vk9
UHSD2Wf9o0lIJ0wWQOL+5GEOdRgn6lVbYa+sdWsKbks0uCHxejtieyrfoDuhNqKlcxSemO7a2Kxd
SYHesLD3DgglCHWQPpM8F9/BZ7439GkRZtR6h21IXjh+ytqZ+SxyQ+/cKBB7w2XmCUfHCrKAnPOq
5dNU/7IqL2XoFwvleVrUas7KdWR/kyTOgyoQYvoVDFOxA+f+jnFzacB5oHfKm9305UFtvJ9tlkAw
wpz0URYsyB8qY9FlTx4AzZds8EhR9YNVWwN1nzRD7IfDdlsbNZZNQfOZLum7Kv0tosrZsoP0MPH3
7Z6h1F1PmGioDxQjiZ3R/dqK0kUpDNpNh6tjmik8MCzUbok5x2DptWG32xkCVIULm7MwzOKC+GQJ
RPxXHUw9Ok2ne+aP2GZFzV6zg0r3a1uSzSQTJYuLWYXX1sAfDM2tXJBdDbAJSs/TXAMLujgM/Y7Y
5KH9rLkybcFjb1GggKW5Z6kITX0uACYkOz9yvS/eqZo+C6mazy6cwJUVcFQZ/rGwM8DOQ0KLsh4r
vMr3LBLX5Lc5VTzC1nr0jGFliowGstP7mz/45K5PcCzW0ccdV1aB+skhTAirzmDmIDm66cRAA5o+
HUZz16P3X6vm92sO5AkVgZzflBA1ny2AwDoNcuiR03vkT5kAPgxGC+4FyBkyEYuMQtj7Fe6mcOhs
lDraXbOWRX3E7C4jimzjDVnRYixEtwa6qT3IB2PGm5NZbkeNKMmjfx+2OOv6ngxpilFrO3lHSzUG
aaWY+qc2LIasXv+iBAb2mHU593cGXBtTH50Vfg9TsRzfwEie3B0+PrccPUJzfMdYmTYGhPMEamAM
aAIRvFnoQo4BWdLnOINibiVsPDs9AZ0OqOZpPhBILXuOE96eZz/HHBEeFvZ/mybv70Fhyy2gB2II
ZwdMqPM/RaU1mNWv+Nhr0JJ4434EhohiR18dtbI544yBstWyMU/XMlH54akrZbeyHOAmLkNzMZY9
466eNen+sgAP9n/zOXWjIICdj3oCOh3ShppFquKD7/aBi8AlnpdrR1N62QA834UOyjt7K43pf19d
aBnQP6ryuqi6z0hwLFkhR3DFva+P9BHRH4CCvctmm+SqrOKYeZY/+V8Yi3sgIBiTCwBdqEogco/5
dOT+QQuxuh30+vG2+Aj0SKTFA9nobOQH01SsN8MKpbqGwDDPTXpAPfbXSnHOZ3SIoFB8ka1JENlT
XmNfxAmaOsVL0JSiEpw6BV9HtPgqT02fllLKLgA2geZJbkXpFhngLI4K6TH1EzC1xpeh3EXx06hW
SVjtLD/tU9kHSl0eoOYKUcnT+QbNU9IeftG02LaUHkbjMEMQ9Xul3Fe96lcFmm9o74nifDSxd6p0
z8nyhXmk0LpNrjuK8aJFR5eVdazAEOlyb+FAnsm7WdfEKDAZngAgqPyhkM8XU3Yc5sBstcGusnYD
5VcffVqnNBi7EJqBRRdUzh/zWVpeSMLIXKIfZisygzD0FxIXEB1x9koghtZ3rBAzvhrX0Y759v+F
+Cbd+oqs+pm8Fl31C4GYmzWkf7H2tfSLH9UccqzH2SfY5J8mJxcXsDjmXx9DE5LpJXRRO3z8/k28
TdNosLSV07UfOxNt386vmnS+Zhn8WygVqXJMT04RXAUfa/tRvqpcPlO0MmqLMaEsPMqepfv/JwLP
ZL+6bplk/38jyKEaIKELgaJM+1l6K97YD6ocZK2xkDYklfkOKVkgcsWZv3p4F4H0sjRH2FuZKcUc
48ObUKP2cIsM+jHfVFbSOC2lTrBKgX25AUV504JqBQNWZheKnB5yl8nGVgWWNLcp0gsxkA1Rd79a
T6+URucLzg5vuijJHJqaZzhedCbG3scDiBNebt4MyyOW+Uud1qfaEn3e7/mcJPe6kewByLU7yH50
mEpfACHO1pR9Qq7B4+PzR2y/56IA0ZW61xSxXGkDag/VDDYECffRRvncc4POtu54tfVmM8E8Y5vE
OvKubIZLFodOQi5+p4TK3LBXL9t3eAWqJoploqxKsMpcXvohh7x/0QhLjy6wrhyqkUOoN4VxWoWz
RcpBkCR4UaEs/hreT4UKQXiA5wL1+F9KM2dL2ZkZppFERgjQW2s49chL2kd9uUdnPQ+ZvCjgtpA0
hq2Jg0+etmVWTjLVzNVdWoklBCDreDcjZibteawlZ6rrki++0NpVmIFBKq6jWDEoK7HEVB/MNmdN
IjsB4xT/BP0spkU5y2NHAT7rMbE+hD6NsKHHWhHfX/g1Q+wx9CtjQoQgl7Xi2VrQXz3vONv3H6AV
6SCRvO25as0PlDQ3N/G9FvYTKFMiOLYMq1deepK6PyFgbV705gjD/7iUz7D3RGc3i3FHRmvu8uKn
s/8X5ql5dc9goCf6yzQUbH7u0Rdnz7WlnFEzrqBkvWlxQfmVQPEeQ+7MWwMBg5HxeRnupvqbUD6c
sKiypW1dqjfr7qpU5Grh4tkV9TJZhgkUtzZRaVUsoDHPBztVTDbsydlkQU5DaNopNwcTKlMQ/L/b
esX7djnjhXnNeo4SEdlYYNVi/R6jvVL3xxOQ8jOkhWDYySoh3H3wSRBHqPRe3gTkbypli8v52P1Y
8fVr48M2lCGMK3jp6wrcoIhIvZLcZ6FbgJI1ubZk1GIe4E8SBAewd0askaWEiDs3mSIn1nHlXyjw
cxv+UuRS8mgwK7AtE3rbIU/V1cUthWigz3CKhnBlgrx7+JDGpxHuYPxsdgyjinvQsdJ7/FPjEcv2
ILEsIfOmCToIw/uqz4s0/ZRpsFPLIzO/NsFRahfuSARmx+UzgUAKiOYkgpHUpgysCXqYjwp2KLRB
w1P3MJedg1FVtUjihsxzBiVBpX3nljt6ujF/J/P4LqZ6K7pELUReRImkN6EKOH2Z004CVCtPZMqT
PLKDWM/qaVaWA0IK8rLJ/iBVGMwTFRkayFZaE5HO2Fz00lliyzbGl/xW0SBXkutDEXnFCSsprrVR
wAu9R94HrlVOXtHF9GOxe/m7zZIydi1xTjJq0YspTNAAPBaQhjSCm1h8+hcXmJBIr1QF5XFqRaV7
F5joNy+UxT3Tsf3rqEPfVlalXVSx82tCAA5ddp9uVCqkvyhA3L54dBqr9N9aKtXzOrt+TOAXio1P
ysl0Cs5AyWu7oqV11Ur0ZhZMmPlocikBk8BjOKT+uNkMYgTqaO45PjEc7QbpBkX42rrVrf7B9NFN
M8g+qLJD/g+KvV+KnlhOH043zYAoziSNvNFm/ERJ41V37OQ5j2siYJJqpsIBAkvTiTnCfGx3bkPy
MVthKn5mVN+hThJLFxlEOgxHsh4cwLjOOigxmI69fMpoz97pKPLWO7oztQ6luUJAWklay9UdgJt8
vhenZv/uvRhiPR7/Lh4EM9VSVjX0MkKYlMZv+cPvJBi401irRPmcUhAqKHjdR1+y5PrB3iJcjgWc
wM7JVCSFpfD9CiUWuFM7lFoHBcvudE7GZCW7gcGTEKNzyDjL6VYPqqKeZoa4gIIghqaaYPoAmkXZ
MmyGxY/f0kDpyvoLeaxS0R9nN0rvBiOUyg5tjw9vs3WkT3TKe30pt09Nb67ML3zeuLlXNFFv6z5I
UoqwrKEblGth0jHQTr80CkAz/TUnMuQuvxpdjcw7JzCmy4BHUpVwsK82sBlY7sWDfTkll0sgJDaW
t9oosU5LoF7cHO5E3J9foPJtnHvq8p8d8PY1urmZrk2BTO5Lefhx0QV0Joy2D+eANcNoFrbiyvO0
kCRiSbjhqoHi0tAuu2EYsvV0HVR6R+Soa0OAAq9bIMvzS1eWz21vm8qCOIA8V/lJN+xl4mHqSJL2
ynr/A4qosQbjKSdrgqXuvFXvVw1G33d4bkUPiPhRciK7+NMptNn8Xr2FmRFJ3FH9sCRXJArWgyv3
2MO0FhsY99halEe9GMa1mpsAxWt8Z7A2ZJNGX6MpxuImRgds7kM6bBXMd16BV0zZ8aaFIu7fBrr9
6bwCnIahhjRqrgBq+RX+Ug3SQfItCaDBRNFgexh4wJHO+kvceishYCr3KSUE5YALkhy6pDsNcIkd
TBXc1JXwSlW166rQ8DkgBahe0dajjPJNOG3XDTe0SARrUSgAGz6Ips4sw/309pCxadPe0f1hpdYu
vdXb3GwKF6H+NSN/66AB4ekXWIUJUpkBKwj8pRV4j7Kp5rV/lKmSNB1U7Y0yuUz27yQHe694JGp/
dKC6adz/WjZbFnyYN8NKGg9NyxMSEgUjebA9HIzmey51q3nJuvcw3860cC5BTMDOpsOgSAo5lNR0
uRv0p0Du15Df6EOZcsD0WHNOmzHsiNs8X8enXPHQYub6H5IYB3s4MUYyunvxnlVr1Ql87G2jddW+
liB7b3G/vcYwxCNwMsRSDTsXVYOd3GKfjl46FuZ5X4aUJdJPbVQYkvyIcVhbrDS38gQ8bBNeTk1m
j2qW59a+rDzQlKcX72B+5oAFBKLVcdKO5jiuZuj4b6k5ztG23u9uPonTvoQQEioe3+ygFZyBh1Yp
N+maQlHIA7WHoI+2s1W/RJCs2XeY5FKLgGXIeg8D4puSg/st0TRNcS/kWQognlg7hO4wpMMN+bOo
hqXdC/V3MW8VbzgDujeHOCvhz5EtcmqP4OMiFbHaAN7EY/FZdh7oOyi0F2jVVa8c8Tm4Fn7BhJln
oQCQm7oiQD4TMbEe6Yl/nOnlCSjIVUhGWnyOh5bPq2XZb4DaKr01YeDcXmHoWAPuXAsJPPE1aU5z
7XoBQpejy1PosFGY7btcyRz5+Z2oqxhvlZThXXYpVho1qSv9HFcMjHy32dMpx20reRmHMvhMD4D4
O7QsTMOK0NizD/eQPtxibz5NY2rTFlO3+y//os0OoT5hAVK+n2ywrZL+/h+EijmFck2hYaiO1eQQ
xNqgHzYaCgfaPR0sAxoAn8dqwRXUU7B/b4U1rldLLBpEAg26KmnUOXcl7IEKDV/fKokXEcwLjtMW
m7BkeHQyF8gsx+UrvD8zzJ6+2pLBjY+iRuCKLQLO9Wq2EtRO8lVt2Qn1+G0+zbseOiwZXu+IuN7J
KZnmqfpMr5m4qgpPLMWXbSjpk9/k0eLNGjkMztX5QN8WbGEztU/gAmWj537sXZTb5kS4cU4vM3mT
7TLwkeGMzE7msGEHf5jTi/f9JRoIxkjx41lobhgAcskcWODDhG4Ws5K67hqAhTxF4VnN17Ln3dJF
zMt/XqvP1WKYQhmJ51JP25wzTLL/T8jeyU0sTYaA34flI5wyGKArHd3Wr9en7tihrXFgZuyev4gM
2QyWO5g30MFvZS+y4kBpJylcdhlQdPh5fUH3JF+6OBC1PwDLC3JQ2vB45RFCT4cBPtzaVHsLrjML
ZPi8prEsnoD7dxj4WTuLgFMX/vvJapQMqX43Nfw1ZWKNYlbx27SR9p1iYXguXe+45wI5FV7z/D4z
admTQGeZrMjsFZboe2pICqrTOLRDrRNicS38Oza/6Bj7ROEHlnT9nhu1ExOM6AzMnY6EQPh9bcg4
+KfRbg/6CAUb8rKDyXdHzpZj/BEOdjRTVFLEPemOf/w2KlXo13JkErhp5PLbRYr0cWXVZaweMZpO
GQ0eSOoLFvDRD3z0H2gLDiuU/TlJxXWRru0yk4jXEO0s+edsV5EmWmlyxy93YaOuVRNQFt66QEn1
ckChC4ZMOLK6DYgi+2Os+f5f/7q8aYoUQw9IyKCAN6a01jFuQs6fPLzvl1jaKjcgWG7rhDoosY1L
pcKquenWMuoGm7aUDoPvAWFouf6HRe8Lc2U0EXfIXVJgt7gUshviL8pOm8fHipVj9UXwz0HlU5mT
zjTls/boYIW5hqSGkWeZ14NtulC2kH+dUQrbwBWKfn2mzeHale3Vo2iZHg9oYpu/9RhwBZBBB8Q8
2XlarVFZvLHZ/UMri1SrBE9X4vCA6pOLD1H/L1zvpPJt7buV1pw+TJjgOCvEwO2qmtEwrk/UHlUb
Y9GWJZPXeaMLIxTnfmJN39qiRZZAD71d2s77j9zFDXqqOEU6wDV98MTHlbJ7PGZonPpDFILCC7jy
kfxX7aNYEdCcWHEPYCzl6oPTxtjiws/7ks+ahRMqeRfg0qcAdy6MGGhaETzXQ4ueEJc7HrT7H04W
006mW6YddwdwrudLMd8Lfvt6yJK0V0Ft/TDvez3hmJtV/H7OF9QfwvHZzXJDCvfD/HFpq1nhK6JC
N31CgAWs6n0GNWKTgTtZ+1XkJeKxaB/2JEAcl1+anuho9BZrlygii7YugJ4Lrp4x24a41ARq6ri1
AwTLqpzgFU70ZXGsYZ+lXdNQtswgSfuQx4CBn47gIozskjcXuu0ku/kldgjViF9fzhZf1sBd5ZVY
quSlZkvws/wFm2v9u99fDv/U9qQ2c57efaeLOZqP/RN7qOfIkmFbLuBxPZ9Slegf2MNnLOXT2a8n
vEJLLk5gnFzBGFGtZB2cR5KAqEchB3k2m1Y0WjqOyg8XFzsJ09f1GaLehiwoZ2sfETRdTwH5uTOE
2lfkhNDP501xvkMK8aqQTdsvGCgQ0n4NMQeaWgop68+BmVctn1lWOlwR4yUqFryFMz7ggRLR13Jc
ezV5fNVL1mJwrIP/eSLM92q9auqVvdt9U+PdiVOgnBlZDLH7vWBMLwi5fIerVpH2JScoRKiX12kh
yVoWE71Iqm1L5mzEUGD1U63lGpmtlcgsUeVJl21L0MvtlXlO4t1ZuqCIWFCHqeLwD9QhLvD+Hkr1
KHlAIS+9x6Z+7Qp+kSptY05mAeJEWilkU/rOsZPC4JaM9SkzUIE6/v8CkmPZ39aG/RUsX7+azojn
FtdzVmVy+50hgv6OaXJ0x8Q9iYj+YtTDhxpO4M0BsNviNv5wJiwQtRwtlqcg9DoOihdNYrKhk+AX
wyNKgH245CjQJQonLzSMEyNZNmiN+HoQaKDswDSa6gDbLDXCbUzGEXi2lz39JlDwRzkZR54WaiVN
PlctHgJ2rCE5H/HKZyyLM9fffK12aVGUsOkQLiKf8QOB/0gfDpGrFR5Z/Imn9I3vRyYT+Udp6wtz
dSYcWtdL+1nn7HfiHM9xpazK8twHdNzJzpmtn7V68LWaAcVTV+UaGYFvRr7/Ycm2VH/hc0QIOnw8
XPva1KBkFIJcTpKrXCebZO2a0SCrTZISO3d47OL1RC4sddfW4cAbnoIlHF7RyRWnmO2lpRw06hm/
iV72d1KCOwXoC9NDlFs9WQbze/4Kkce7G9Ra+fvv7wj7XdXva5tskZpJXM5N36QyHqRR802hmWxG
fgzfVxTAMdJtZgtJT1/2VKtnhZdSMnEvZVpqbXxSISXYmaW6/6CHtgYD73HtG+RLtpU1BJNsCdfw
KUmAymB+eZX/vu4mfo96oxLiJErcyUSiIigC+8Vgfw9YtSnQ/HvsrsyRH/OU7pBR/LompRN7+ra3
SrLbULtpmxBiO8x5rmvq+4eYzaQHer2AFSEnaExhpn9qLQz/u2E3FfQtZwOYy77FNpCwgRWmGU+v
54+Kv/7yT1RyPkPc9Ip4IkTiW4xfXpKps3YZFUcC6XVgdYc03vJz8puscW1vq1GVkrovJAG4BreR
6TfuwOdse9DQXb6gbtSVvvowfhihyoS3B6AtTI7Grl2cFVL/n0TEK3V6qC/U3QvtmwyKOLbV8Jba
W/PyY2++7aCg+g2MtEM19r/kjhHeD7Ln3QjgVX+vwPraf1DKUbBrap4SoTngB/FeSUMtqPw3V6iu
3CPwU7E/CCCaFrI2n7h4xPJrScYIoyddo3Ono4kgwuHWAx74+8vRS5jMKNY8dtLBXoEegeY19nKB
peq7EJgbdpK2mN8Im8mLD0pxy/tKIKz8vNOMjGARqIuD1AeXDiMdY8ezSK/G8C/1WpGAsiO89VAx
FvwUB2+1yIsFNIWGBY9D/dAfAjImZOv3Qx8DaxzyfGuKKRsE2FKMHub/4dF2wlmsmGH1YCOEccFQ
Oz7aWE2QKp8UbOeR4nFiD7XsTdTGJWNvghdMSlHcuGSsJcn8QL6RNL6e+Cyz+Rx63c1gr6v8sn2G
bmBJs5H8y+rsiRGySjAdGEItcvXWIlLvM/7sWFYFoa2J+HAyefFfcCga9oLazSLZpbvq36/zC4CG
jbsP3A3rQ/dnYfyCBcKPvB+pptEUSkY2YFAeLdlTRlI6FCc25dd2JEWVmu4LXyuUGkssims/2rOR
OYfJ6Db4YV4bL+pu7SbLOi3JGtYe2AGVu+uc+Gzxeh4ifT5ox3hMQiVTwQacjEuA/YXiy9wHnHKq
AKBUL+dzx8GZGpmmmJmIqpI+iNqfsIbtGEsX0FDOg2P0trCuxZ1sv4HACXGGkLP2SIhFAYUqbI7z
tk8zwGVh/WQksVRRvZa9RRivtUadvXyNnWfoHT0IsOJKUHk4HQwbvO654aAjlZWPYJONcUrHU072
nbnnPRthsQKJBveKyrMIVlbk6YQZRdtOGn5xC8IMangWSu7p59oeaay1obneS6A0ttUlQD+mD3yk
sVi4RJngcm4ScP0O35R05U3rky5mwlhMR2z/w9VO1xin3OPDA0gtDVzY69uRHAv2DLeXf93jsEtH
dA+LbwLALBilzPI2WcZ4xi5hNzptqBxsT7yekTyV8P9xbW8Q7n26JF+m/lqLIbtmO4Mo3h5XLr1M
E6mSszpEq+WzNGVD/gLFmB0y0Yw+lT2t8pDBbc1dZR7Zr1lkvSkg1LioDWa/6DIis/XQ8xoACjUN
jVcC4whND11rFhKhAWIUJRfumNsER4/bIwUOyL07R/zOlNi69KKULBMLtsuv+efu2XD7fveApIN8
M/EJTK3owr7WKasnKoKew1uSIX5SyxtoQojA5DSWuQHvpqpuBgHlLNwXUMXWfyxDa1MKrACT9Kbg
WPMuCKs7mHFvYyW+YC9usSDNejAGcLUlf5kp2Par8YFAgMvIjTbN8bdMcPgaCtAZX8Bj5N9CqQO/
b0ntIhdquSkt2kwqnoJaF1kPeNc0jVtvR8g0j6VtXWqiKcAQy7bmfDw5bXc+UwUcrdcCwE1aiWi3
8tu8RaKnwowPneaQl0H9+q6we3OasdEhtHdfbBiqvDpFQw/Jyc8IYqsTTUsrTn9v8TOD4hBXMIDY
oJNe0bkPJUMHWfMEjiAd1hDvep/JrZgWzwyq1zJS9Aj4J5RTGlH848AUWT7TbLZGowmbAq1KmeCA
89XpfR+A8XORgI0sFf5PRYXHJQewIR13AfLFhNu7MV2czZKM6DQYsNz395ii5lNgHKa7twEpR1jt
E2UfDSutAdCzYarkedchAM8/epq6FrxAdDyp6Q8GEczVzta1zeaNSkRa/yUdTl65bgjSny8kKQOo
eEhTYBrq/Q2FKsS+xn1IV6ko3pHI2MTSTxfWslWvQmWXZJmMfQu6DwJ/PS1Wex8NMOsJj2x4p7zU
3J4bEw6X0/f00RRzSUnJcjizD7eD7Vq7Lm/FQoxFSavw8tm/eDWqZLnC4aR2AKQdrGAYUkeZrCrV
BbmIuZ0TS5nditObg3UnA0BUHHfr+Lc+ChKKcpRGNhKUp8K4+rYkhUJcwdIxxqfnkPirYy0AT8HY
O652ixHKb0NCsDR9vO7pc8DMZI5M+5MIlWGoZAP+rTMQ+NPghQ9TVhwUPmUJ0ewW6P/S7wzf5Dql
vGhW2PrUQjNFccKFKIN2KvT09Pquj4yHbgmA4w370MKwjeERSE4BLbvILhzHhes5xdroomE4QgvI
KimE5bGFv1UvyIjUeXrOmI8f5sqwOvJjvDFZZY1l2hjEKd+R7Jbjklc7cfORI5C6AZ71/S6KYBMR
eFSQeJKHFK80yQHiQ2JtiiKNAWJt5MuqkIBG1rziNCY7OFZHpFA5LneGwaLDVysvybrOkPgKUe9k
O15N7ZwyKb4nCfum0TCPV86l9psI5T/jpZhqjpDkILQ3Yn9kwigMDAstcyFwJAniNTvrpYsXIfUv
3CMo4/rnfeCjtzxMOVy5w6jKeQexHpzJEiNMuO48gqHth56IsS4D1JKPLnA8HhTIfRvBnFoicOJG
bmyzg7jlqIfGwSEvGTF0HCuyfBmyQrviWFZGaeNqbxrZEX/qYzZJLrPNZXRtpZNo0U5IDtECxj99
qjrPad5ZPmBolvVeSsVU2/QaVMHsP8nt5jrxnSFaHUKsAhdT5lzk+188WIuQv41fdT5njz6G7pcJ
hV4tsYR+gKf8kr8ML8y5MRXUHwY7NPQqdof/ljKfuTjUIMthVn/sHjM08rTN1DGgQDtMgr7Anvx5
j70YO0gjta/vZPovHDZpI0DCUcZpzPMqnR/88+tbut1c3j0bmO2C7wT2PVZZNHbiqhc2DWw4r9GB
E29OjO7hVqe6b83jo4iGnKBVe9zgxGmRHpAyd6OYdSd0Ot/H9vG+ZWTqQvh3rS3J7Rp8Gl/Unx8W
8Ue7tCYNX6mafLgzwNmUsOjpvjq8B3cXxChLDqC7GczMtDySPidUfKcOxFcMmebRdkkYx79jUEmb
53vf0LREyzYIVmPA6y1krUJ6Ey+JDwnqVlMuS9W3twlM64j+e8SuvCqTchjh0vIV56m1fiEQaVUE
CevCxff7s63a6M/XoNtUfIFYMjVMweBwCD84mZbLkQOA+xgwxrDa9lB6kA8Uuq+FAbtD9pyjvv32
N9ccFxaDOxZbW1vftR/oOm2UQ0hXmiXyQbsqGDdMTMLp+tPiRqrQaIV2o/5xe4JyPxWDMYrljTxa
xg6mee6SHpLcV6LAFgwMiHtfEcypLmW6zA6foQAHnLbx+NlCJh1/JNjE5jJLrZWV27Sj1hpkK5+i
NYxdGjojg/FKI6rvLQNzvGO+vTwdEOzMfwqwqHoGr/FH+pXNeylDi/cW82yY6QnVY0H59eq+eKId
bB4KQyccwEl8nInc6DFFRxR63vVqrr0z5ySC474utk+OLPf1x16wIZkNIZcRMz7E34W+CcJd0MXp
SXusCl0ZH20wINULyJcBzt61Q/T29zKW+4fSoCiFct3cSBeGILdbie2OOOJTW8lvRVQr+WJKoHkn
5k42f4jPKDObDUcI6sewfodnmIS7crkgvghZ4P1JUgQjmqOZWfSquai8MeRgMY0bn/8FkJTJXdf2
EbmVEccPu1SXI66am6yoXxTGqJYRqFD0dZkqGIdSNQHekDk5DNjpu9ROydyaH2WAWcnvoE/Dkz9I
OaecmYg+JsZ5oq6P5m8sxFz7ALBmEe6nQM8YTb9WTRPSL5NS5b2ikRxYbuF5hXJHyN53hRUWk/23
FJXEBcoCyEuXJA2/YxvyeYnHMtOlIxY85mXST+DtnvUtHwOGd7ycYPJdPcewMags5r+Tdg4nFJb5
JXbk+RyDUVR70EjPGtB7js3gIRNlYsSVhMQByNQtTeS6W6UuoOs4RjDKoqDuj3e5Unp0EHmoPWsi
y0ofVL5FNhWc4yONUt5Q8kkl3QG+RhKhLfOAEwHexsQyA0vVvWn3FoPCfTaGQNj2WWdR30VyVVjO
p3pS1Oc6PGb8EufgrFe7cmChS+pJTnR5N0dhzR/nKS0DCmTlRvqy13dSW/Abk1S2IZkfza+U8WiL
v5MXxfUetm61y7hiq45V7IlxCOjhGpzjCiz08a6UIE72ic5NWPh/YvwX4DV1SEO1vkEd3aQbj9QI
MlT3+Ccfc4dy4P/1/A39snLYjBOwvXAk9dBJZPAlm7Nqnu72ziLtpcmRXcQVjJTlfTwCeXV/STWA
SAK9K3bYVOGFGs5JaL9FyZYbnmOA4evcHqIEturig3ACVcJ6KpiqRp/lv7n06TQ/gaQamvOS2BlI
A+Cw+puH8Nb7gJFEP5WfrrXqrZKWo5vxPJXL1f0+Y8Y22rULsh79UGNqcPyKMNzUxoE07Lq3Sogn
6eP8nWKBZOykzdHjm1mwZp8Ivlow5RN60k09zIDgl/qKW0Ak+i/xNopDn6RgIqfN2BTP1hOOqH+b
j3f/jBT0XCcT87a19oQD0YlPUwtXwSSw37KXs7gbbQwN+Rfg+8I/FjaN1mzS+hHa4B9nvTwt9LGB
JPwtrp4oIzVoup8RIvpbv7lTArydT3VktVSd2J9GUdOjkovsGt39Cxp9Q5mB8wTg0FFFTEsSy+RX
fRW1Aeio7n1GxSV06vThgWeSmSwcLjPqELr1z4JHx68ZTUVzzodvsxRJmVcEokHnr4PreI6ClqTM
SN7mZg08/HjKhIgHlqyEUGJVhOHaoEZXZfAn4IQgOSBGDj5bAeP1QVWrA93Zuk8/0Oo1CDRuqckC
DbEOVf6tcgO3a9fdcXTHMNyTNDe3nGKacJD+PBmIxnrdQwPiYGH8M55IwZpM4ejbS/Q65pZBtOAy
h++V40NWpalFlc61omDut0cVSREunmHu2vpWJm18G7AZivEfM+lackNbUcgAdPdaPPuqMdBXVFBS
6mkb4kkPyzc/dcVJHU2vAh+N0DTZ/LwSkrGy4TLF66gDCI/LJ3bzHtX4ZA/LOyL6h53eEb39NQsp
WkkCvaLo35XBnDNWVy32i1NEeXuNBWKwSn6OYzjEip0Q1QN6NB9Nqyng4Rt9alOGGhPFQ5s7gwFg
X4jza4b6WEOmgmG5bqQfjj40eX7QzUo3i1WZRFlYV34yDM3YeLtV+cj+oTi8R2mZRb8l4oaWCkH1
G7AghUxpYgm3Asx2Qdbql1+6HQN+UpKZXnMQcNd1N1PSrFVF/i0t93TQc7UwBgrR7/ErUzWNDSkJ
hr8xE7YuvTidfUn4uuodzqG7pEEslLhtr02/ysTSWXacc58B8G5IaUke+Lng9XC+6F/vc46OQcYd
87taPM7u7dhu9gvmSdWescgSc/0BHw4x2M+ulkWeYjHq3DFysBwOvfX1hr79WuZtqhCQ2NNek+pT
dBnu3pHYzp6Ssa7QII5FUuFhItF4ZtqDmAMTdzsYX5qxamU92M0AfENMLve2IihSjOuGjhbJIjfh
9aVesQGowscTobudrkHArA1bIcu+Ns8seRr6W7WcNl6nif5rQZet7u++DTqNDs+yKuh6a7fRVAqM
kKrJXG8c2HXuni6Q2L4Q8yo6ZjoR2iK4KzC/rVTqJGGAtexTKc/zJd0PRe5UKqfnqSflPr4ECzMo
NYPejGQwLW2Z6EbbGavIhkicE14RuWWSdRumP9PaibHXJh7U4pG6+c/M3msutvjnMDnJp5KmKtO3
QMBy++ZtVRc6yzWRg8E6wzNOFgkjSDVpU0w3wX9BKS0D2kBk0DBhj2R9lVNsanVzOAewJg4XDepJ
Pe48XKq2vnuUQtqQuwZULJIWsxhIJzktrAYO+rTBQjPrEO2nMfvxLpRP5JzYyk6R/3t2wfVLioK+
dU3MOH+8bBloVFFQuIqeT8cYFf5emU69WPhJH4szeR4gtIAdQ4CAzUh3PdgwWPo05OMrX49hrnsg
hSWKa7aINvZumXQLNn/URqmSySRSNIYuwAyJbhmOAIZ/aIcKthFXu1zRGE73GSS4TiBbBDVF1XAO
Mw31pRB9LtAeY4xLGjV/yLy1/B8BARZ1xs047/6PqKAOCNwlQrWubKaHWSyLziTxDZTIGwKj5Fgq
clO4dGaIVXqk6RTXHo/FddFrRHMyB9okhl5psTTDMC1E2My4MI/5Sk2oRQmK1BlHBQSGhSgFUk7U
Thy9V+DC830S6QlbiYPQ+4+Ik8JjZtAYpgDw7vM0ByMWRoaLFFm/cxys4PCFdXj3ZP+A6cIN5fVk
2t/5L5XkhhjCBMJcbz3+S6tkrTYUzyj5tHMe5+A5yElgVwBxfDMQYGSah8G21FJrR1xrTxOOaSYN
ksG8DOqjr0Xd7d81N+2uCP8n2pAsqfyynoyL1rkcmNFXeXmP/10Xjq19J1hWaHpohDwvMh7qtp5N
Pa/nr3WcYSVT7FNuLPRNwqDk+Jah1of6W5aWOGyA471lkwdS4v4BeCpc/np5kINGVGm9GSZs8YOP
P/7OB4nhH+Ogfa9rycnKVb5G7kaTDMkwGEjtvSp8yog9acPY7wQfOUign0ugL1W+Ys4o2h0H24nN
RyuE0qlYOmmanXEDbtpKX/wHs3NLteC8zerV7tzCm8uB6p+duDwe1AUXfJ72An2eshxyN4sBpCTH
Pye/4QPr28NjbWXYvaibx2Mnv/mxkzWCxh76dVpAiH3uYr9JZVSyVbS5jjjUSyRtepApLU9HNClX
mm1CeyOr6b4xlLP61MX7JSjWj9UjelCEZTL4sHS+XIYkrTBrJpfn5M/HqHF+33a9Zji+Ki4zIhD+
/w+c4jLDmrJCHOAejmoRjLFUjxP01JjnX0aka5l39u0wiF8b+pyb2HXJBIUu6M7PaokPVPl/ql83
bLV+NVWFarKeM+XZ+2nMV1Ee/1K/lRHWyMH+u8BJavHTG09cFDvrUuu8iZ7ZqaCRg6JiMRMKcYCB
kJG4wUqJaCn5Q+0cqLajtNHq0uywG/33Hr0VM8HgrYKIVg6kFY7MvEl7eEK1F8sHagV4MV6JDPxz
fw7fwEtxQtXHOz1YVpegAQFb0SJqo4GCOE2YMfnuMJkMK7oI+NZavfRbCT0x62moIsz16qFmjFMa
EjDapsO2yqE5b7X2un+v/eK3SgwnsoxRCyZoE0CMZiE+afvP0bWCZyd8Rm4o1axt1nzvarTTg0jb
eywckqSz/JEnk1DWt6EvN47SXN3fYC/MSwElTKCx9eqJyB1R+lUC+yepyweWn3X/tv8nuOKZF8i0
vXkYupWnTXcxJiMbEwEn43BIcoiu98JlDGrwQSVArHLhdremJTSMf4/PWI19llCbHiojwynPzPMI
7bNRR3BnI2oxP7dJnMi3KtJFuVSCX0zDK5FXYkBqCAzwEvXS8Onfzj7yAvnwi1Lilchicfp+RpQf
IZG0qz12Tjn4fyQcdhKcbZyek5xQm/yXfEs9S6wTYj8e9JTS5cEa2mGSJorST3O2Dydhz71lsJRx
zHBPPYN9gP5duimfCdi7WZz7kCTnJONlKjz4TSW1a6RqbhT7sRub0E8Twc45L36iIja/GXl03RuY
9UPS4k0QFZVrHJDWugTmUrdc8gxNRYQO2PJVUiTOp5LqvC8OE6uswS4Bgayzbu3BXeaRQm2oy2OW
7GfE9e4Ow0VmaUAvFML/iSK+ISNodA4L5r1oKNv7hRvndDnN1Z2YIuU2eaSiJayAE5WmZo4YeP3F
R9WNPeUFFunM4dIG7/ZGhLJFCe9ZuLIvBs/kJmAuU6wum9Y+cE7Py3EEomQBHWpcpl399HSGXpfx
6v5IA10GEcrHT6ilUALJgwnbVHhIol2B4kM0hx4xI+7sFMg4SOcSZ9Wk5KQKaR443WUObbAvo/lL
BXT82uy9VXTUIHJa//6vPrQNOMm29VcfT2EiMfpGqqZAoV4F1U8m3KnWKdhnJSzwMya4z8QhPuRK
k/Kh2g0xhvwwu5SNi6iixChHGLpPXgadQuSOd5lQAjFxT+grJ87MrolshQnuHgQ42sx+nA+jPl4m
SUFL1TrMsZKom2377phFLKKxIeIccwT16fB3fgJgCrp8Wtcu2lpC0BTR6z7z0RmpyTG6dIsrpGRi
VVnQBhXd09FiOBdYx0HLn4eaQLH4dw0+waUUif1yUvd/Zd9Js2qw9LfH3y4lysK0fFuwFfLJ60d8
GqBMSuTliUUMSBcY156wetvsngj4AD/BisTB+1W6Ck3Da6COXGZaRrymwPE+S13oDeTd+sic0vTo
Dgg/MaUMCfmwG1790NJS0sCi7eoBDr287PGpvD94Xe3MfcN4u9a8iCIf5c60dvYvvMUs8LtqLPp5
ba+RPzYbnRrUEBHDJt1QkU41Ae8+L1foMQvs1o6K10Oyk4uGqln8PtddiQfDojSY8zLf1giFpfIx
eK1wJlAuRIgYvE73J36Xgio3r1aNiSga63m3HSiBZ1/GRGwyewNgBjf+HCludNQj9FPCkVY/77Rw
+AbqylSBAr9VMdcCeE4K/TM+uDp+eGA6o+he+fDs9AYTaGEJvzpHLjduk+UdH4K+Gpn6IGVR8DoZ
PIErm/rhFSXyXvF0aOKmg/mPAMFGhSLdAqvBqnxecCtpSbtWsphJ++Nqn/l26XxlIu1qy67xLgMY
sBybzOkFroopgZusF9RU4BXZbE1avFUcazyS9feFil7rVFCGwwNFMRYl0OOElOV9QP29xLnkdATo
9tdTzAzx1IqES1SRWcbz6G0MZxjLMRKLbf9Ai/LeBgA/0mDnwRxHLNrs0P9wZuiJTHZnYIZwG0Ty
+TusEsIKAv049NEqlG0ZfCDFhi+zNuUTghGuzNm3QhNd1CD2P62u1okm9pTkHqrifxim+uvboZNl
ImufobSMWS0X5mQTnAtBUvNMl1L6sjoMv9ukHVNXplAvCS3NJY3qioz+ThClmUUua12gGbC0eVHO
9+nCi3fDRG6ySb55Qt6hWvbImCpbBc80XiTC8m+hqFYPrPDuowiN0LuWJMrSPQN1syaiNjAZHgbK
20BbI6ZQXdgbsYdTirloYG5rR7qsbRBshKOclNXlkKUqB9++dWqT7o58/fx7XQu4eEFaXrUEEH29
agznaX29/mL862VwYpH9eJg4ylxyLWiBO6JGxrZQkNAH3eUZ0D48YpCeqpJ5h3fk9AXSHM3tdE7r
azShxorzLXv4z1EsK5MM+3vSuZJJoxkc7OK3smUWUKdASp7Jkp/JXNgIw4JXtyVPuKCePSsAJREs
3RvL+evAFS2vaL4+4eQkuoA37rtyCv3Ziwu+qR93+8IfIAoGmiSAQpV1MhuE16Lhbis0J1EVbvOk
L8wioMwWlI+75FJhhUBW2idVp/KHRSdBAd2hIQ+CVEttF0iSPxcsheSKGLCJ6KvNQ7CNLVKuLAVY
tX0e1YXbeU950jY+BZYVWlhMZ5+YeSG/lE7yiwztLJjPkRzeEd0hiUfk2KLEhcqzinK8IvXyW8uH
zE80ygE1LN20b0Ls9F4LoRPQgKZkauxAi5wQbzLkYiMfBLFPHtrhX1pQ7MN5ChDSRF9FV3Zk7cA2
NGE5iw7ybPec7Bsmi8GwjCJiwAWKBJV7UZtwAU3YKXaDojOycpeFEQk2AEHi0g2K/hvkxdCrH2GR
QYTH86sWKMOLHSyW4gbyeydwAlzCXRIxeSgR2gTkZww4MjHqFfKLMH8j0PQ2oI4iLp9kB3kdST/b
aDWFsPwE6CpgimrOltOKLR9Gn/mTqQIAM6D/GM7Yaf8k3tFlNd4rrKNHMZFSuLkxKKsOUQRncpx+
oolVo6i8w377b4t/uc5M6rfaA9ODgNWGG96mQoZgOSOE3UhoAjTH6vNVkov7oEQ+3uJRw4cd1X4u
zn14xYRwHVOnBoxH8w0T3SpX8YvgjrRU/hqLesMDl65MLUML4Tx1s04bPgjkU9eiCg47XqanFPqj
75e55vR1J+SJNadoS6YrUD1E2Z+8Wmw7G9Sw/p41T3D4zIFUPww1dnY5q+CRjiFY7B4s+t1WFD//
iMv3kNkXfSbEXCGwO0iblxjrQEL1oea1ky+KTB9hE9/+3806RWZr04es7D6Qmo7wZ8seHYKpMQUG
BDDjuliZpfArLvE3FgL9LuUoXt09L7UKDp+J+DlTjJWnuPqfbKRAbFVCTIiGcrI+JpIubxB1IdGZ
0K8vsLtrWE7QL9Fi+HAmlQcMnYWs4Vwg1hJQ/w2zlfy2pAFyFjkoS7nRZ4/jzepGSPn7u0ByUOCD
jzm/7Yox0nvzf3RXqm5nRvduj/lMa3w1dyLgFq8QWXEgMBiUozmX02CN8Z0/c7PPVQxlMqxX/OWr
bO2C9NancAi6j7y0VJmU1Gb+V65QNFWGptaA4wfZmCawp2/n/qbEV3rY3/DF1oKpNbSr6+wzh636
vtCV+ZODY79vLBugFvYpS6f53b0cLeDGitvuS7JkktdsQhGN4Nkc3ym3/Ug0hy2tC875SicRilmC
ul/r6/ISUvi2IsJ0qt1keiwUS6hr4uIEBlgLCs9R15EmDlkX7oF8IFvwZ2Y7AlPo32mM9vKrqoca
hksJ679fqj3jClJphqY/brduFPAmowzsHKnaxP+EsLFk/ivUs7bI9/LfEvd3LomV0Un5OQhSRbNC
zaiYt1CIrlPEJHyPOWnxm4kgSCNuGXqxV0MHAXDNINZK0vIFr6HEqqP5ArzwrOUVeR/q7Zut/9nl
YYjTZd7Xb0bEVVAMoRVFzr7Rj/4SYi/z9DkeY0qiR6arIBC/D6+9gzvcAYAH5eerI9ArUroodd2p
gpoYW/zTNhBXAU6Nl7RaCHSz8NIZXhpHcIOlTiWDnv775uj2t/qmtyuEMJe5Gm8IH7nc8mLWyXtU
nDgDIs12t6OUm4r+bZKh/lVvzFJty6rSX78zQAD5f1yqPTBuGbS1bmB3F9oZiahaCRUroieCoCim
ed11BjnLODGQY9J64r71mNk6SZnbBuYRG8hMM/tRHFy82hRqRc2HLcrzatFV9S7lGLL7Zfxz+D/g
KTXxMFcjieNNpKugKOqfgN8823Rk3Jws7pkRYD9mSt6sy5Ux7oGMd1LTfsg7c4nVIBpkXqgps+gv
qWmTcvSkDhFepo/qGrgjm6DcREgnROXu2bJTwwXU0Eqddqmo/HPyFbVP70proKJZjqj9ogTc0wPS
dYX3gkt8z+VeDBP129CDMwdO2aBv683HqlN8lozOYMvJo3ZucIxbnsPKojfK4uDDGCD3f8usiY9n
juJIOJqFjqSkpg6t+8iNvURgo5x8Wdm24WaiAvsmFx9Cd8RPh8UNkN4xxoRZGhquDL9W+v/QCcVR
fB6odssaoxRK8KseYEHrNKD2c+GVICrny/Y6K25bItBATL0gACc547vepSRoWXDYsludUqWzDr3x
WHduQxGk8lsj1ZrmpcyWOUsMIztLYRNDts7TDUoy0Xz2yeNpHruiELgsD/TtHK9kvrrJqzdI5ErS
fs0/H/Fv0Ziy4cPJtFoFiDsKPp8oqrBX+GoUbLGgXuZci58Mj9Pbvl+ncnhRKEr02fX03J/snXR8
9sD8lEZD3tY8MglS1A8Hw5zK9o3XpWfeg8Anrf1AMieytlyh+A4fYCXiJ21iBSSzZjZfpzXyduJO
jvCoRYDc1Lgw6BeLCYRXXvN88y7v3X4/BH6mEb9iSKvkq2wmiXotQncWabfb3tMUf/zC6Y67g1MW
bqhMrppxAo3aOmnXpJymI2pYn4E02eKSlSiZpdiznBZ9goPR/HRyFGO7fvlp88LhNJjKoVFf/jqN
JLSrHaEtn1k2kJt8mvnmVZVbNgSmEWtBqxRsICCTG0vt4EZp1v08q80V5NftwsEW4pso0u47iyHU
FxmSMMicurvazcEN9lqYdAvvoQ0Xj/G4KyAC/+78j8t0AWBJGL1o39G+ad8mas5O+VCRPVZhk6zL
BTC0BjLfhNcw/qBxsM+XYSLgT0CBYsPY5IWR6L+/qOvw8H3vV7XvMcpYsbTwkUHULlzdULXwXByX
rvWHqvKDKYIGdSjiG7QsQHfptjA27QRMxlEAIsJ8jS7MQOPkkmigUAzLNu1uWigC9Qtq40oHMPQb
T0PsvCVLIQ1CIzkINuqdSAfz9F4QJikTQ1koH8qlqg3IQhNpPXbtrsrpyYUiHMmaD5vZ/7D8vAqy
6XzXLr+239KdtrUdnIjHQ9IlppxMI+jlYE87RxBiQIr/aZQC9O1zg++cao6As6poRHweLc5uC2or
zWBjNITvXSwAf+1ydGwTrUGiXnLgowjf0r1NCg2p4haNK4FLgh0ye4Lc7l61VN2w7IQxylWjvecE
Pm1L66mbX7IG5etHlXknfIFWPL6rQXjXdSUzom8iwtAcl9uR/cTV2NvO1pEJIySoVjOctXzqqD0N
SbzRM4yLM6NuRq6wiBLxsUUT6U/VCP4hUE8nop58F34f29G3lUIJ9IOAn8dN0D5u3bfGVVX0PBz2
jvhTu9Q9DXwFGQbbQr/Z7QVDc1CwAWEoQcjLJDFWEjZ5QwddK8B0B0eyztPgdZRTBTlbHKiENxf2
R/rfiiCDE104xyLrwNTKf4epuBbVUfgRs3037ld7K6b4CjeYpl3ae8+NRi3oCHrMk0FKlVA9qclQ
7eUT9OOwFq8s/y0z5vrynXImcBCmgd9AHPWn275rT2YkohLiL+C87ETDZEI+/CbgR5apeGutmfl7
HSgL4JaITzZW/nCiOmlDeiHG+G1PMfdluJD0OV1sxA8ooNZo7IkD51E6Ww5633yJUl+gGNqJnjt5
IHB+iTH/A/xpdbvS9DYKJiQQ5kN22DK/FQmUUHaT9zEKogeR6VZhEzqqc1LMYqYEqMSFMS+HGpKz
6wDeb3p0ehaHZGRtSsGbbvrkEGxsMIWW92ZEdS8zIXFaDZJqKH+l48QnCfwQzfkkuSpuinq+IjvT
5Uo2abmDt/T9M6rOQVQ79hqkABKKkgExnJyiA0puhE9vw9qBCUy1rAVBYbROixq8fRc+GKB0a9R+
G2qWiK7so7lsm87N/YtLLMVs2Odbq1XSKUlDKtM7lNc53f1jy90so3tO4OcU35xvMWOsKi0Ig0aO
Vl8FV97abzxsjkjwy668/iPcK/YJLxvdr/u5HFtIFTEcwu4L7cS3hHp/69ZNqYdvrvxjtGVgp81o
6zk8Qkieto6M9bRZkia6T5TjTwR4Gy5VIqu4CIbe+6lFvSEJl90NzAXg4lJHZCRQJIX5VBPfrdhE
BR8bLilo2Dl8WmaG72S9lATquYf045f8QALOiEeo75q8Q2UqaIzIr+LQIPuF61pRA/EM88d5m7Ft
CKsAec1s/iB3l+USYd6HaLQRbkxDqB3TPOi2urmPws5UdasUUeL31YQcumQY3d6h47BEtT7KnYkH
q3H+msJeUWebO5EKRmL+785gJvXrt0ekpz9f/9kavU0pBvLgok+eB7VaOltnYuM2AdRZC3sSUsyt
QMUzRr0FZph81Pf2XqnLuuy1A6YrJR0k10OdR/65zcv0tF6BkvjSxvfngImOC59a9AL/v8YudGgX
PixXAaDWCYjYkcap7Tkqo0+jpYHfYy9qrYyiZNqEH/TCj8JTFB3LyiXvodkZfnq+bJoSiIJDsDBe
dM+jfEXGbtS40R/SXwZ/CFWaiP8br9/n3KgoPs5sRzkAiiHUiLJYC2gPM5AE/GwNzodY8XxI7riv
LUnQ3KY6oGZ963LdKAgZjWJ1GHaPcU/wx5QFPWeeqV1esimKJNEsCIl+n4+xl/N6+oCaTfk1QMbH
G390zpl4m7nlRl/2VOGZL7XXMhD5Qd6sDJZPtsUNl0/0gMfUbCCv8MOeqmutoIvrvoQE/a+dgntQ
42fjtpNa+dbNKFp0XmyQ0VWtqKTmtM/pIMOJBCSdzVcIHn4f+1H6YnVg1lJK9djyPvgsE8tjR84q
TAeEPFMYQAzT5E33hJaZZK87Tu5c9ES0ZmYfgfSQCB8F02RpQs2O50W43hKTbV+Pls9g1p689DPB
thBjdH1kDCuvqxpDcBnv0jS1Uuz2WAQBal7YCmkWBZkogXkytE8H51obRf4tFu77t+NRDy9jnDdC
uLmW59/iCaoBXOZ/r+70X9NQxJm9cQuVVgIgPac4dMt9Kx4Wyf+uSGd0yKppPLpYzTkhlko2I/IL
9fVV19YtPMVH1v4qimLsUK06vn/crFEu/JeypZPerrXIFcwFxIaX+krl24oBKQXveAvSh70kufIf
k/Qu2j8IGlNOvvkD1IbsBYWI6NV1R1c+oZEYwj6tlyYLhBoD4P/9vemTPP+3aMVVIhUgzMrrB8hI
vGvRa1z1yFj40xDDOSCyIHdUHsqGbwZlyD2UPKjFIwxBPEQHQnWw3KBMkJt6ZESwC7kIpiTE/Gu8
GNt2t5CHd/R63hD9joZUiyFXHAnxnbpSi4SxTY6/WNg2ZXf429C23ddjDzzumwOnFHEAmfxhdAlO
oT730IdWVJXZVGK4TGnUuFVRE+JXN6JmMiuTqskZAyJYB3BdUxkR7sAnj+vI16cW2uQIlr6s9Tv9
mqdzdg1aAyxxKHnTQvLcPU63Eyo9m9Wvz1PBHDoRZzc6SA/UcyEHzsSKEaqjbFqT6OXvQmPjBsEq
1OupION9ORHK5aXuTui8Z0HYU3FpmxrQk/dD8+e7t1FqyYGUgwaMQyPKeYbf69et6lQ0Qy6NEfLg
2NkYUM7Bw43+e8LxeWFuXSpTkVSXfFNK5B295Vaeau7mfA16VAqRyNsfdlOjVHM03925XfgV52+j
waSJC9EEJy/YlYT381ePeS+oSk4dMo5JTxauLew7eaO4Lw5eJgH7IQDwZjvC4Szj6chz0VfiKtyZ
6QphJD4/7mjEjS0AsWTpXMny/WaYA6Xo1/Hxe4jeK6TqZclRHhywlv3VVB0D9xOTQ8OM4Pj0uYgK
1cjd+TLpE2JlYbArxES5RAm7x10TEaxNqZkMku9uIMSe5exVEqM1eORW3e1b9+q301JyVQVHOeyp
0CKGqmzIrfPA94nsKEcWenymnuNkSSGeHtPSb2pv/WokTTfL7/jQdPGlTBUBGnYes6Z2alDcgQaZ
kLPb6E4eLcz4nI7cQChGDSzXoO8YmgFT1eotG+gDV/uR/xKl/vKchQd0jLc7tDBPbYTCGp6JHkWC
IoXiWw/Xk2uKfZzKlniUuF+wGYgs5cDjDaccW3pf/IxVy8q8r1RwLEWj/rWfaKMk4sJw3hIQWU6e
LmOSiqiyd4WqLfwgOrBCgjXBJgPV9V5sDDi9iJ80+qNJl8oCUdNj0AStjsS3dHBHntuy/f8V4CoX
zwKC7Q7HjHEhI4krwedTEXvsTZekOy7wBcVDFb/e/jKkYwO4RdO13njTlPldetnWLNvESQs84MM4
MSNRv8jc7c0HJB3Fv6AWAdBDu5HU1yBP43CURja/gBpzvR/BYhaBO6nVk0GGs+Hhd+sEsWs7QnlL
mcvK7qnOfi+4F+OIdXLitxP0LVpkTVFJNysyBTnRDhomNdPh6bLS7ABmcg0UCTDY0Ziv1s6xLdPF
rUG+M72cqRPSivR9kMxDPvrPyuu9WwSOrR12TnZrXcRMpDaIcxheup+t52oGWe2Dj6I//fPc2lkQ
YtwY63N8WRnr2yBdM6yqhDSiFUkiEVU1rEHchOcrtnFkxuKVw0wrKHa7Mr2itZ6fD+MCti6Zv5Ne
Fq0NvYRT2TPEDp3m54MvMoxTJblUguTcoP5MwceyEPNFX9n+8a1WVflNBl1vH9ojbIrWmMLvxioc
WBViTKDWkKMdeNEj3S4DFye1xX1i+RhfEdo50lwupWHCbJ9gaqfpoaNQcJ68JJCOK8mI10HQpZhG
TXhR5RBrhamDWOED+MSplP1MErJ6HUKC3QlSRU59cAk88WJ+2WXeS7gGLhJWwsUyAIRQ7d9eGCrj
2W4QgnwY932kDJ60BI2/UDnFG7FffE6MoFdvW3l5MKJafKOh2NoBfck4X5m2WmkETcwufsJ50NfM
kyID5IuC3FNmxha9hmHcnOsjwsLX9CBvcky/yzX2A6bQaq+XC2c2b1YsBvrdxmIBXtfF6hAhQFxS
Y2eURfjAhOdlllcRZ+ZKv+7c1v/0DbaS5edQM9shdcYPr2GvqInUV1XUy57/bll1Wey+7aT3sAkY
ctIDvdf+Ekk7yYXgdmJYZmSjJ04FtcflouiPj+Wv9YUzUVgKIvuDjEm3AsfT7z8AjHe2Oy9Rk3hw
OIbYntBoh1Ojwk0TJaSgTkVgERaCuguZYOxSQot9JdEI5eEk0+Q4TQ1fkiG/Lf2YqX1DLkCHAq3N
3ykAfRo8kS46OqXlfsSSl+QfJC5dldi0eB5NQz6eK2LqwSBH0k5NwE1wxT1nX2GD5BUk0mGZE4kX
+s2wkmmmaFtYIandBB2d7RlJ7x0QnnR/6D9PiBni93jUR/cqSzMg9G7IxB76xrHD89kdu9hTGXJ+
AP3cQnIbTK1FHMSoOajOhRNV6Y6JOZGKlJHmARBpz/HcXGq/JnByU2OoRmGkb9AYa/39FrlEdqj0
oMfeNOf76LZF/Cx4Jp5pUvR3FLysBKPgBfqP0/ZYLfg3E+IdPW3CHW72wwaHzgynmgIVEuha7lUi
5y9pObLR0Z/RYhp39J/ROkBWmH8+IrWIiIcl1Xkal4LXs6/h1Y2b6WjJY7fZ6JLtw7fQ6cNERW0N
NVj7X6FtMnQTpMrUnrGJ53r7K2Q0BbiytUEkR+DV3hmfk+b33MHPWCbFsZCxeaK+TYU83q2+la5r
hHjz+qXK9o7uUH5B8JFbLoBx60Cc/3vjHozvBoeMZvzf9MR9CKl0Wa25af8RELnn/OSbb5/XYWep
gGK/bFEMwmaQisWiFJUkZjeJRuLwd6azJfQ4i1AldFPCT9BOzFFO781ayROkWcguDE8J0g+zd5AP
qIaQaWMNoYSGDkDGbJsrTaKn1GpqHKKyEJY7bQe9Ox84VN67NPnmKh1WxgLH2G1QboK1Jgz44+MJ
juQBjsrY02SF95V2RPmYiEbKIo4WBbA03vjSAYBqGzDAP+j42nc7k1/TQ0ceNOL/3QtKdGfAr6jW
jQiXsCTnyKtAyJPB4f0MfOQSXxi/PcfY2uhmmHdI6hEtUxaoWqxI1CEPZG+gLpiIr8ebFnuiyDih
yt39FfAJ0sRsRQ4F4RgDK+NSkKf56bD2dt/JHObxgReXEG+vKzVogPXJKOAwR0GQHJySQRnz4XNM
Q6VgBnndDBdk2BMskwg9WIycDdb5huumXGqrpvnqxI38FhTPUO0bADRnmEeb+H6BrQGMN93BzA1c
ydhlI5HOSs/UELe1kJRJFWyvi//+oeZc0p0zDKgs+PLYzhfMWlfzqYD5xwG8zMnK9g+QbTJiigFf
MOFkSOtPXYLbw/mPsFsdpsxlxpacVOcPfVN+wf4UV3IdRgsBq4M3DIL5wf/mc/3xN8ljslqU7bcz
VIat7pHKU9pTCa6S6G6IRxF8rZqM9P6UOzBti2JxFfrf3UJXvH9snzqhzeq9vy5CSbvNasOtqY6U
G0JVv5Yt79kw52yj0ldNRYSRQAD3j/OsV8P9LVx0jqAGl6V5PYKoOEizoL9oRgXzg2STSGhSccr6
dMiWEvS/9di2M3xCjfpD47ElNQwNKtsXI0vtzVnv5N4+tofuvufi36787qFO6KWsqgRJq8Dwu+IJ
bc90zUEA5SIvJcjWwrLcmantt5ZRg/Z0NXnjDwoKZlv+n0wN7pns3gV2r8qQBmlSL88ZyBNo1DIv
Yn/3lMlUKKlvBywIbcH1OYugGeUzWRbf1zJj4x/ER1T1gZz8XAHEJ1REtx9MXxAvSo3D75gj/qto
ekfBMcaK2sX5nJdkvmDTyYzdtspjGoc8IWgPi2KyJ4SNyQWTrmrzP1Bg6rpkFdiQQ1/5/5zFxCxo
PrKvzVzpQ6fg7HOMEM8rEeNW8FY9ZDonNkyOIvGvZx0YJMYM7E5Us3sRP7ahH7tNGViC2azhDHcE
IjLqV0jZ9XVbqqcVpmSPiQy/7g8wwUPl/OLfLD2xoRUc36EMkuKxXwWNLJrbCyiS8NMi09Yb/nA0
ldrb0ng8O8UyXOo0vqW4MyNpFhwZxee99doo4/OtCytYc01IortpvMDz9p8TrvM7T3Ohz5e413bn
mEnC/JOUT803OBgF9d7IQgE5DRN3X9JmtMBiNCCPjDHFmZQSVwypbfcJHgG09Sasd+gjANUhqZEN
OulokDb3RSXrhQ0C2DJtpgjBn1rxavy2BLqqsIhLYDTRD7ShAcvBiOcH4LMed4RNp9Qn2SUlW6Ql
wCLF3cnNgpnJ395xxbpfqcF/Y/OlzGfj2R3BbrRKEPiki/VqS22xt43pm2wlDhOmHHzG6dSHjUzM
sMuKbsH6dkxaXrBevdw0MdDRmt51HGbkzO3kTt7nn6puZEEm3FozjcM2qqUcZqsPOn/Ra0No7Kgy
8C/63ZnxTaj1G6m18H/bhXIDptVCH2rQSOhxFNoOIeMkjzP9pNDqIJpcu2xAEzhP7tOZCDRnr1Mu
awB9/N0JpH5X6ZX1/wvyXOJNcTzX75QsqWmAXVXaFRDc2R3l3ulM+3htsNXRHyQSCXIIvMrjA8H3
wrPP7K0ESF8IVWv5/ocWNGCzssbu4GiRdjDLqQ8INLGYihL9Kpvp8ktNcdwSBC9RxnC8j3BzQzhX
mPCBiwpeAZ2pMViBSCePilJlePPxhjH6sBQcKpCsK60e91ZPC83X4Ftth8LzVtwep8QXnO4Nn1vw
I9iR0Mg8BziSsqYRy548v8V+LsV1LAG829GhIqppFXt8DvMBtbbPEw5KJCOEhUuLDVodX7Il2+AA
gPHJp3PV+KyM8KbWILLsrL9Rbwu4pnxcrpFb33eKwBj4g+trDXI8MFyMwOiVThdONcQqFO5B9Pav
UvudY85R6YZz4omqp+F9uBa+yeROt8Xl0UauXAPmw4E+oBwlauk+oaRVWSoRgqM0MsNUcQ/WrPqp
Rmo83rx9P2xIuk3zQBPE/EVLto4OFx3q6KuhLLuSCMPpMc+Ng59/JzkFpVvf4nN12YYCj/l679GX
C4ABi5xClQXVxBgvYM/0jWxua6h3dnvMPXsEgfeAXQQRhVNlFPlA5vvMAHVDjz+9VIJ2jQMLfivV
ob4DRlpESssJKonE/whqe57EV80eFJK0AyrD3L3fyu88E5uEwOT0bCh6JcklGfsWa98VMk4XmwVe
xxr3KRnDOG4gfBNhCB373Sn8Ckdf3HBNHIwR5Wd98+7e7d2V8KW8pWp4yphD4aUG4UFjabYsA7do
Hscq+mQep2ERufXX9HD6vRtq3yu63nPeyLdPVtuX9+Hha9KkGCwWOp7sqJcpogFqwbgKSSy4wGV9
ky2xdOK94GMoHpjHfEpXHEHvCUtKy26ayf+EWFGAKzRxViRgBDwALPpQimVAwAaC76AGbFjIiCJf
7Mqqm35lRA+QnS2K0ru0mpYgbg1T1hG/nxM82dY24lR5TsT8BX2vbujfStIvUYIHKC47G/HeSF+L
uJwzN+vqEiBZ2HKdHvQd1fQIyv54orLGAV7rziFgHZ8p+Gmqz0au5HnCH1PbU0VXhXwwm7Uia2JH
2NChqfQeOSMz3cZIBSeP+TppYUlF4Kq78EqEcVCJ+A/GYXcMbyj+LkMV1z3ilbsAeNHJWafPAmle
oZF4zgQvjyRrzDGltxj4E9wMK+KSe/TVCX5z0q0By1IGRD/cn+Uuhe4RAeiQ+AXhefpEUvvXcW9p
yNLamei7uP711NE5NsvQfnqyomUhzvHsXvr2KukHSl6FLPrE5IgByCPe7rIYkt/KeH97FUvp2EUM
Fz69W/TnTrFnuvAwZqzpcg1nU9ej2TNG1aLSiH41l2S3+/GlyAv6nok1y3IiYzTJJnc0VS0jySuE
EBTRV39mq2+WTIeZS0npkuFZyJ6Z5TlFpFdOYI+I+8X4jQ658MtpIsqXY2iNTeZjjKDj5Zhr1hmo
ZLVN65oT5n7fBvc9OUud+fqIcrOq5fHLYneqYfXeAro5n9aNjaLHJve6TV3P7yc8VM2nWM96PrAu
pcHSLjGKSfmvzM2HqS3HtakQ+0ZBAkxJUxg93v+VdA6EzMq94HiSmNf6wkJRcarqhH46GQQTDO+4
ycCA0WdWPYsC+bORZYEeNbGHbIB+/YcXICAWdSI0AYHmIGmbebCqr3dpysDPzIbQbCrjMA9TAN8k
ZFHdympbElbUZlQafYR3MJiUpSu2gwZI67wiUx6cFckdUQNwAhH2MjHS3oDa1mEKRW4pvQJhgttK
Zu43Ceic7c8SsLL6HmgtaGpQpSinwueTzYpkbUpDzhWS19PS7nSquGNQuCuHc/YTJNXDP6PorSx4
C+3Lv29uiTpungIMulnqYLsjTWccVmo6ECzzXzJCA0RChz3oH50cTPX21dxHFsyWmART/1/vbmMx
lXbqbajgc1TuyriE+gOzsXUm7VWkRMqvaSgwJT+uZQev6Dkz2PKopSme9rv1qkE0UKkJgIAacdbZ
s/6Iehnltk/MxzgjG/kmAiI6Xpg7aaH/u+74nm7OOenIW71kePtcCB6cLsY9ULdtnSKxw1PmnZeL
4zfK3TzmVbGGJi8r063TlW85ZWBBbL5aJEczHRAoAo0+kbOh3kxrw+t2OV2TTbXFiqKl17j9KxFq
JihWKO0z/vRpJKJzikrw0oCxZl8orScxg4YJ07bOVwo3KbeEAjPwFnOFqWWPJVHF1duFcm//AFcA
W8DMryWzp/2VhZcAoPJimf8TSJk5kX5nzmN21EEHjyqDavZxeBpSGj8/aqA4JVIXoI+Xccy33+jl
tqO05maf2eseZdcZdE8I+DaCY9jkCZv5f/Vog4LhHDwipPpmgsbKICNU2SZVEQA59nfGNhlzwSSa
cLsyH01Q47qnmCRJWumUY/HdPv9auZlIVXYNKRvJ7hYDOjSiYwoUz+C/hTAoVil+PQvd7L8gHJER
hw2Ecxu+arrHJO+qU6LiszOOa5HzMy2ZOe1nragXodPXAsnaGq4XREEMAOKxr97U3EXpMqJv5qr0
PTZyAR8lGg74amBAKts0jlqbJTYFYMenb9zshb+8Se6rI8xh8kDCSe23WRyv7nPFDx/WS7J2rxiS
haO3SfG/DvtmbsLUxTbPx+x0OELmcSHXuZVe5IxVBDlinu8cx9miBcdjwoipTVKqQ3aIfk2We7X9
uDz8u+Dm9eHDafZS2zm5+E+rZoYced3sZwpxMwLO24nnj2ZSiEOyqxQD6mEc5DUnyhwbuVTdbIXL
97TmdFFVsRyuvXvTPQ/Qvahk91ZWZbCmZixUtBaE+3buz5jdTDwf4CHZBtxB+MBafP/TJx8Na+JW
JrR64NJQSrbpvrXJXBeW72HpcfpRcXu1gAsgxSJ0wK9NWTqgHY5Pz1NKkb6DcAgdMUK5By6MjKtk
rO1bhoZv882DOLZwcTfK4xGV5FT6TF88GupfF8JQkANos9btduhOI/UcVpLLud6d86+wvjiP8q2k
NIXZkaHjtCxKcUrm6K2pvxZp08JSlTpf2VOtiLsCSlJMR2pq7wYXc0PCpUq40sDpIQwIRHxSSfNh
2e2aqZ7xqICSChJOFZFk9f81t4PPeYH6G2E7ajzG+LVZa3LR3m3lojUDX97QrfSXixixaLTNKlnG
d4qAdtsv8MyPxtAvSTitgBctDTnec1nXVB/7xxJSOZDu45Jqw2I1L2mvIPVBWYUpQO0uoBvPCVWm
KL76aPr1DjBzujOKwaqGLhmiObmua3n4AlJ7grO4v0MxnPBFQPTqTFLTAL2/bg57bnW3am1rXz6p
+lPsZ/msa1dSDDiqF2ogWxrBAN2L2LdlCn/ozqVM19PYyQvQnijMFG15W6qlo9D9JUp22Qj7s5Nw
P/0Gk3k7KuFtuGivu11T2oVje70o7TEmO8yF9ozoLJ0RfwIoiC7h1Xo4keAyjDA42Xv7WDM2csf9
L0TtkpMM5+K3AZ8+FdWEEmWQvrLrVhibUcGXGocE0lDnhcnk5/WQvPhhg7sRakQGNNeX6yFeZ5ix
0GlonYqXxRSAI5Af1+atRPvKvfSjXlgXBvwwTz+GhC8ksJXDOi+HmUiXjlXWwt736I16alh0+cau
SAcfhuYMGfc7IPUxhFx4t/U+OOQLPcr7ou2kuhAfNMm5uTd83s/SrZdbSw6b6U4N0ABflyBUeqH2
9bLX8rdKhW2QllqZyLfvGF7VFruVukEcUQIcsl3MCgXCeRpCNjM/C9SFoJzYRO0SuXXXaJxDjh3H
H9vsjGVpXoHgElmDsv9YQop93zM3BbMGDwrZf+E13i+pHUNQkvSyLeZxCVG/iE2TvvqT4X5t9psH
7P/cF+QRVNYj32fYODx7Qdjdn/Wql4G6v/84W4FZJ51tW2TntjIAwKqlgBUDHcPXOnCdA77RcvrQ
vBbkD/Y6HcdebnnIPBxhxrEzhOSoMi8lCTy61WStLw4KGnQU8OJ++JWEMjFVDJIP3vTKKB4mQLXN
PbWM1LePP5IFzrKRDIPVPGXTkYmPvKtgAgHYAy4nVZ++5KoL0NppYXOKs35wikKacWbEWIiluQ93
mzXPFh9gJsijW4R1zk1Oq/0YVjC8uXEfW47dvbOElIRIbVAHrdTPyhlHGqmf9XpPu1KGKNVTar1E
hULJ8JIbZK5OsQYHBiYiAnsB4DosHBxcFmMLv5n2WcHJda1Hmo2ztPk87ZXbl0TSZZbDuRtpaxId
1a7XdCtrdAV1GIGFoDCumbolfRcpBsN2PiYF+YBGRs3HkYs2hPBzNeoen3Nt6iNAZD4EqoEYjPCS
HliHf3GegIEbDYyqk55iyG1ROyyfQ2eMFgnbQJE+F+k76MgEE+/4XLwyUFABw1N6tUZNcvpICVwe
iVxWC1+XlhWzkcvhSSMpN3iJ6LnyynMTd7Q368OPcC8WKVzVcHy+Yv/oy/EqmLqrh2IuViq4Quz4
04U+pCsSt0S2zLC5nqj575nwgBnmaiEK6q1pc7RMPjOwcbxCjTBUfquoJF84cSpLN9+LdOUKH31n
rAIK5fUp4SYpCIUGjpmSDgW1M4enSppSyrKqHZbn25PlNJRDytMIULppAPkZcq5dvFv2e5YiycvA
xk7Wq78pGyi76ssrJ95E9OoIieHyuwPNRnr6z3OCw1n4Ag2dSU0Y9bq2YDt78KOOd8Lg9S7oprni
mJH34UP4U7wdfSZPRj32PkiMlDj3/95tdN3LjxOi1qdUZyNBToAeTLkv/KsNs0Z5aKpdnKIrloHk
t4n7eN/SAuCMF5LgnrZdIQvzIomOznQscmCv7r/jwlD/Bl2/ErDxyZpwADPgJF5DHYmyfmP58xyN
3liKPOkGWKc+D7t8r+CNzCX3pPWz95iLi4BxXYW/MuLD1QqmemcXNg7ld2+liyyKZ9wCK5pjIDvf
pOwyw1ittRgO7Nw6etCBNY53+NvkYI2kR9Oky1SVWZhp9mBCKOY8GaO8PdMao3QgQCgoAvAsieaI
EP2AiwF79VLiOKdWe6GSzFgcewLFJTG+0klmYzDaoqC33i9vNvztcWLcUc/dPMW3w892W8of6hlW
tHLx0eQ5gReV+vJDRc58LGjh4S6GI01lhgWUPs/OBZAvr5pLgLHuNWMYIUhvTyEJoMbhZhX8S49f
ISzGGyiJT7LLi5LIGtuUHuCch/cDK5Uyi/OIMSqSd/vVz4ChBqBG0JVC0jWLSNym4EF0fHRY065P
x/PLRT6xzxwZSWxy9AoyGaOARaeea7918tc4MLW+t9rT6SgmLnxgpMjYG3aAVxxC8jHBNkmtE/n6
iNisbhAsTXhOvH3vzvGYAJ3eZL6TubFSROCZvufIxEP3ggRUZZYdHzcUO7hErdGIHrwqlK3mrX53
gIZ2Zo5cCEsCKxArfmz/tuheSElvyOMSAwekXZOiRoNCJmktdyMtT/UboXfXJkq/RdUUuLfgQLFv
g+CyShlg4CeLemoRCHNQu4qBlloR6zo4AbHSDF5jAi7jsoowIluKU+hOvH0jVeXRLpLde6+9ms4c
+s7hs0mi8VDZcYcMRXxD2DnfH7AeUFspmr4WxwwNJWPk8xnFVxd2UVrY4OAA7cjJmfiBpQJeJGGa
BN7J5ouSU+KhAGH3v5zdxVjkpetDcLzkk8KIVz+rsXuT2beBWy6Q6Vbjuy+O0rv6Ns+44IOsyqqk
QW1jEFzCbcyYBxYbbBR2FYra5nZKjLhn+SRgMGZniluQLT1z7TQRYy8y3+v90xhreRPEL8/WOSF3
JfzehqRoo0BiJq1MdfZm9zAswvwx6Sg4PxkB5woxuAF7Xy871JlImdofe+U5W/hBFllVbxg4Ortx
n1O0UO7w3ckdZl/4mVL8+fNJTEV4G11J6XCj6c1AqUWkqn7bd1Eddx4xC63ryVYGd9pBHOg3BTFW
RpaEt2gGR3aG0gBR5AukMa12+0TY5TikVAivn362INhxjRsyn5uNPjjmrc34IGBgubXgebnjsJfp
WVL8M9Ln3ozcXFqg725WUXTwOEG6/hYy1gAABaDEefw1YOUrvIbwig6b7vKF3z8fSXg0DHGVQui7
WLBRthlRHX/WGLz/41n3L5bZqFXhqDoIkCpxZ0q/RFnyt2ZaFiEufKEcex0Ouob5vpd6A3NlfZ/r
aXcJULvkadrD2Mq4udrnu1jghWp5jBwrSCi1SqWAFYLZqACImx/1AkAIOm0ImV4ai9hJX70RfN/c
YnDjtg9P1dQkDv/jzorc6Q0QZCs0Sp8Q4QJxwob2MzqL8qAtFCSN3pMeZ0hoFGMREVkJR07saXJS
CgqHn2f6Vfg+9/nC+V/Yv9IHIK+/8YMvqTZjQpAPboPeSg/7HCfORVKlShITjsMvQy6Zvgj8FBYT
GNSPdumQPLjbRisr3tN9p9eWRTmlBx2GBKtqcQanVux51vSx6DkSVAGYnTfgBFLHM1WmMilXz+w3
iqzbLxkyGUHSaheMwiC22igd/vB0EK2W4OhLWfYym2O6BJ3sqsEFSvs1SM0acLHrNRACjWVXaaqr
WUN0iYUVdOuIS9v/8pX+UvhvmCpT/CRNiguYvGHSg/tv+3ztjV+YP1Gl2yVIDVIVgtfVdU8bLqPw
VHMY4JTenXSaBlofithrZlMK0HtNd6FxJil+xsbgHktyiBnwiSITjEWEWWM3xYBRLMDwWG8FW+3G
oVryA5fa2uTMh4H51GIIiwe1ifLXBlrYYbLZnscjgJG2M6aODyLnV1vF2AmXT1+Krc1b2m4YyqZb
WHPDlD0Fam6T+S/IhfQ59bEqZVyc1d8hOdlFAwpzka+agF56meqtzdVd6YGllL3EYxvgOq7H3Z9+
QIApD21Eaf75qn+WZ1uth1dtYGe/+sJ1RaYhiAY0r3gdXRnOtThkfaLX1w750B1JhcrEH3NE0rrc
qGfWf059EUrIz68yRzedtiekjTqzjXgecu5KDczXDqUlvoIA7zFoXvb6GEa0KwFhAEvVam/QtonV
+ELInotUK+/vQB5HRrLz0Yd4xokcnLsW40LS5qNlwRZG1+d7g09S7UmTqsF16vMQRTWkighZxgf7
MrLOXmxwYUCxDaSReDWpLtrjLlBdPaOQyyYuTscnArpeMBTZI8DOT35e5990h5l6kPCuD2dUNIKB
H3VAMHRkg39FpRhYxzEKk7ttThAxvX63TeNEB1eIlcgU30DlBv4I9YKGtELKRbLseBKqm3OcK2NW
S0HldUeWFwwnLztxIyNDg70qkkFOTmZDYtkFXjVQvtixYUmdAqDGigeEvIjrM/mGZZtJ3f5dnOyZ
EuVZVqyMEzrwxr4lOpUHfx+fKoxf/AHExZJQkKUmJBKk/3c4988bGGgG3cnsgTeaRI3P4byZg7B+
w5xwbtRC9aabCauWog2wJd1XKZxARksM1EI5CD8FOE8/xZLCrZN1RX58AlK9GQL7XobeDDicAnv4
Tfk/ar0mvp3EaMsQQDtokfYwZgDQ1bG2BlyVe1jYXCRQwuHCXWlMYHaRtuKQMx6P+JcI3BjlmpCw
P8V9jzTWnGCuMtvuLOW3GPqKvfwQ3CNOV0nHS/E58ZKE6UdVDAPLE/k/VMWGU2LFkmwRYl/1y6+U
ssggmxUqET9HPYdHgEzeG34nclhORqdIcJpooxEC0exSp6gFyMP83Vvi1btAsYLEXqTxSagWC8JU
srToHf5Z9CPXds89wb4DjQOB7l2pgoSltlp1MacZtjpv0zZ4Pvyyoy6QD6WtkMVWHi0QHU8EQsXZ
bez694GdAdH6oQLD6oqhCsCxsXoQIAyEUEzZGkyqKJwlKs7vvws20YchFwiERHDNMwqNr5lrpjY7
KD4anFoQ7gHcfrZHs5ImaLvnvpaaVKnxhbeCIEgmIHqNEGGSEkjrRSyGyGznjE9yXblkfkVUSVpg
j3e3uW8WOpslTCHsP59cUQZ6bQzlAadS5KYprgY++r4Tu5rzb2v8TfNDGVspNI6A8hVl/7yX7CI2
ljXUSMFW8eU9oXuZHQEllH2IH6ryAt6R61cCMT27I15g+WcATsK1Wu6cuEF4w6cmkViePLA1+nEe
1KCQC/b/XJYgg550Bk5mIaZ9ov3cj9jo8P/y4sdqX50xV5UbdHcjvuZKyWD+Ca41DsatDiPdqI6o
iDLMJVEklQ/NL0FGI0mYGn31MhV0Pb8dY0NsEucjwWihbaDuincIv3Ldf90lJ5Gep5p6/6HliDvj
NXhZqQSpGoCM5DftDC/8RSDaFhcy6SdYldSDL1Q3TCtuYC3qd5hHF8VsoX32feHC/9uI+cd7up5J
qgk7fgBqwLOYTlCsDNVju1/62kth/3kaKzM3Ezshf4wGO3xAY68KOryBAV4a1T+7QDKZPX4SUTC7
XKdRScJDNbnb4FMgN6ogZUyAkN6dIqk0F1Rp+oRHoi80G925O1RxpEccQ3pnNEfLMOJBkh/kwEam
b1/+h2BAGn7BFM40KAzV96uzkRcSsNr1BRvAnnStYk9fbcO6NptpqGlm54Gs90Sa5k3N6zrHPZaq
lNz8ATj3FFkqZs6zI9H2p0tk1/Pa41Nn3BwvQw6fYyqA7mPSuu8TSGCVg/Ums8GB2Sw+G+BYWEXP
ER1M1tOvnDizvRT8FBwgp1pQz90SbFsPvUAkTL4bt/kFG8pLWcTKQFLrLBQnPHq9xJjYPETfHjEB
yymY3HmvHd+ROHhQDUbeJUHB8Xu2QF1NIicWJj7r+QVQz+llC6Zkr3dsD67U8XyovTXI+37e3C4l
JCM4/RKhYqg+dDf5lIc0YUjTnOB7fQN16Wah1BRfKGD3us4JZtB7CJ3Lb3lIyUYxtOipWDUZyown
F8fYAH9Cj5nF9gX3zZZZ90tylyr+MvQmsbKYjXuy0YXox3ISD5paIrfWgborgASns+nC5nag3rlh
8FXoHAI/cWgs9wPBpRA+BYZLMQDznHWLjiQnCSUZEF9LMNxWXKyLuzj6LOvU/eVl8q6HG412BfOv
J05/8CdW7VRbmLXayZF7BaH38v6kmO1pEzlQiyxW0sBVTyNNwt1LSdpJVfBdZ+Ju6B6DHzd9I1Ol
w6vL4vGDI6OvJPk/iUbBq/gbduQjTrFgnrI0dKZ/fKjsY/SDhSI+iD5xShZz2NTQriko8/3i8Z6s
vYtnsYsh61m5VIhGsIf9oTod1B8yt2aJK2mOStE8YT1CvPZI9RpDPXME1h4oFkC+I11GxAo3ojpM
Ri2IB7cW6Pl32wDOR7bAB5ixmP75tleqL21P8cu1RTlgszqiuQvBTf9znQizkVztfIzhKQ3KvcOX
O1Rrux8+6KnN7JkZc2YJ7S7X5flPInKJDNco7Vn185QTLRCg0lDnFWYA+8mdmM8YGGawI/RG0fcH
LwSHdzlYI/pAl+ZxOrpT2hd/drARvK+A34rQITVwgYxBqdB2Nojwrh+7CKKzO7dxzgAyoFjUEbB1
orfTt5Lcscg3E/B/dmtA1AzUNcAi7Yw0TDYEVH7lFDihUhxiYPCo1MjcbRiQiANqS+Aj5jeIzqO/
3zvau/9/bRrtzqWLwwcfWEjuR4zZZ9Q4J37jt2vBGf0PTNvTafZx7y7ziJ8m4MnEpEuClvE1v8+j
YIekyR6C+6w/ipBc8DBYT0MNgWih6X6AalZeE4096dXmxbievJRioAnPu0YYyCAuZzrH/7cIVDMT
OTnEmFIPm2fFurbYmA+AWpzYGkFgKScX4jEGxoNq2fJ7DA4v6TuTIMcFR2w6Z//qLjY5WtStgMff
f7KZmk4Slq3aeDeE5TOy7wVBEAzPoVNFmn/qBntn1kuMnKjsVznf+1Hy98vSkqXuNaA42f0M8imu
JYJQHNc3lANJtqgNN8SZAWPyS79HVkZKBKNEyTxR7r7/+m7FyUnYP2GXQ435fhLelhW74I3L/xT6
QP7x1KpuHOFKEb6yz1AODeYm58Y0aQp+O1FYNkrHPiAS/sOVlU7NfwdsCXE19uT8bNxeAY6aQC87
QPBK6/VC8AeXmUrOI5GTrNcZ3JgBpYTit6P3z2afCzLuH1r3+EYXEzSwwlkILDWkC6a1yU24CV/E
lvDv/38/L2rp2Qz+qfE4zKtwre5kOCVIdp3r8cvQUEoLVrXNx9zzSfCuwJMHSdsEHo8y7S+qdzXb
cC2X2aExiUG1c/YSAxp8j7cjYNhsjf0LwhpeenWpn/yftbX3IgZchBjFLGx5Q1AT5KdaivrQoyX9
yhmFdkCVZ1M8UwO6DZIxvkDVL3VlBfon/Uiv4IM3D2RqKjsHpTI9Uh1pLKI6KNL6n0r6+yOlKZ3Q
GJXGfo0QlYgYILRaFx3O6HECb6l5wfZnOw/syr2IkBoAJLcklPSSov1YLuLg6Y2PJxHPF3Chwq5X
BPbgMkBHL+MlV/67uk9O80/ffExYK/YKFQq3frA92/0ns5iyArtY7DA6IwNmpHfUPryOT+C+b9Bf
XfGQZv0FDAEmM0KKuhh6FgeVbFdRbSzT7b189PQdARfMOd1R/NJ1w88GiEOKvg3LoHcdDs9UrFzW
LrnM8cy1QrgXJt3Gc++FhvI+QFprWNzKPR3PlLCKNDr3283/VIwkH2IbKCvYd1OlUdB4zRYgJpd5
kA+dEzSraOX1H21TOIVXMQV/wDeng2C2nSaYqzIwGfKtQnZYLEFXA8CvR7maSNZWkFrBD37z/cAi
cIaW9mefvYI1NngVuiZRNjUWPdDjWZ3mG7q/OUgL4H22pLYEqMXFm+y3hCzmdrC5WE4uLQ3LJUGA
hFIBpEDZXN4ICWRHy8blwK8qdPwymfAFURIb4eM0a1l/dQ2q+sXhzP00a04lJUmc2jdz9W37QyGQ
HgXBVVMd0VLlik/nSNNSt/npRJOCirb0Y6giW4ew82DGb+GQ9ujZhoom+ucCAlOM459UHmvf9nr5
UC4TUjy7jmCk0x1S5caa5k03VkVuN9q0x6Z5XC54iM91HXJlHQV57dkrfirULWKTaLCz5SlKqRg/
ui7aLVrW00LHhiyFT7hR/pKWJi8k086b3wehmG8Zs+ldbasrbnU1a7EICkQt/FcFX2adaTzmXfLh
yfDjwGFpqSFVNgxwiHXmHdHuu9cGdESIZzq2YBfhgDa3Ok+AGcnftJLXjNHlOU2DyyEDvxISOmcr
Xxfai0eCKBadSzV/D/K8gb2vjJQ/m7kl6U2jXTEkrZ/zMG3etclHBDFPtpTOR3CPJrQvCNhnDVTI
eATlDJH7kzGartwlo9SmBEPn9lVTEBMsoR99QJTCDYlXvhOJi8o4GK7e4DZ/dfjI/5V+C7P5kSsU
o8iT5/UFsFlWVqxoJpGZ3p7qVIVa2K3RdadyaZmmUd05KnvG/jLZVIX5y/iG6M5uMR5cEMr63YLQ
Q1yzqdHumrvvwDDXJCq1Goun8SjwYlPmihboVUbJ92dEcSksEjYd0P49UAir28YNs8ch55rEUhz8
9jTgIQcKvL3L5nSMrdwjQl+1pwUdfxywde8nvtdN19OiyX2RcV2ACEXUW/iSFPTWeXrDxqMwb0LY
ET2mC9VcUvWuJY9DS8cD90ShgJZq8nE9T8fc4rUmWQMy1yYGhTlu/KZIGuDQPr12IZ06FyJqqddN
ofLOfC1aaQ0zRt9wcUn8v1hKcUGCSbbzai6jPusbrl0dHKztn+P2f8xKy+jE/L78W1s8+/cfibb4
6Ta+0g94xj6BuIAKdY5zpF8H8cbxtYPElnDPSsLkNV0vOys7GyJT8CNa7bczRitHlkJ0RW0PlLiv
SFV/rcQ3CWT7sWbjR2rHuSy9xOXyKkrY5+XK5myt5lCCaSlKdnlVM3f1x90UfM9qU3vmThSw/m5X
p1oCxrJmogEZ1t6W3UpJLuDNTF4yjzm00ALcUmTy7/l7VxY26fGwxRdoNf51rkxRqOLVMImyMEoV
uH1xd2qR0/3rvFiqi4JZIqySWxuyRQJLsPPnfznhXxHORqJOnGLHUZ+EpgsVmlUpVyfADj2WFBgK
gB7x8H0lPu7orlVgPx4OvnGEd99FQ8ATCfSqaVtF/P6SKXBKELN8kfDcucJdfjwmPlr+k/15Vshk
yZQX+0r6P8ekMFhZpLiaYgTYocgBAvDYu0JNVR6ECajUNIB9b75Rdlv09O+QGrivYse4JoUjgCRN
qtEKoo/PfONhC2zN0rdMRwd7Y2fccnaMd/fed4Q7mtuhPwWYE3pUJdNgBQG38q8bQwaXLiJ44COU
sQwnL92UOOjT5JlK+P+OL0HdLrcbtHaLz7VFUdCImm1C0r7co7HbprnIcO41JyXrjMwmFbYSTwDA
Fm9RncPgJwmaS7Y5IMDExkplJCdmztLOMgY4G3gpg1HA52l+hFmx0NK4zAtkCIrVKN2htF/h6Mtw
lDxUXU7IYyp4gRUOGUKmyeWn/we1Vns+7p7dyulIedLwptk3mDbx8tcEU40eRemALsEEnRZajRiO
8Dnzcv/FbN8L2VGqzBhLbQC4lGhCCeW6IW1+IqA78xfcEveZv4YUu0yncaBy/XLBOgoLGUUbWWwu
oMerXCpS0lKGQjXcnr00d5sABEzDCKR+GzzLNHti8LlO/brMJs77l1RIS7gbLM+p9zUmXSNBVz/h
sW/W8BMw91VbD5fwFfzRwQ19YqnieHIRgdEJrOHud01oCFpkE6+4mv/YNEuZsXdp2kuXtIa8w6sO
UKESkgfDZFZy3WgmVPZsW10uCHSPSzt4I07pRf7St9YSuMcjjXvnd2aulZ4Arhqh9hB7EZ0DfFc0
DJahZTsQ2GCG2/S8OkkaV55jCvrO9kgEsWcRW1zRQ6UExMEGQWpwy6ovf37A+U0vDPjAvCtkOIIv
urzn08mOHptgO1AiQisZ8lYlnaH7YOY43adgqMNX5fEE7v1ALiAIKwQ6VXEHaaRXWMy614W+bcQR
5P9dwdNlm4z/mzGlY6mrXff4Ba7KstDwpMFSxDSLVmWjvvOR9zvM71N7kPdphQfV/AFLsUhqTiN2
y8NpvZvAA4lzD+3g2RSaJNr88WJjHVWxSt8W2iVagyfHvytnD8Q54PJ3vIrAL0/uqumggE1eRCtJ
cmAEPBckxVSjW0Osewud9uoLGYZKcturDneftIstt3qg5X65Gblh75OPnCHFlpkwADL+45RoboL5
Ree4Z2TbNsy45TJnP/omPe+V55NKBtvPYgClQu9ZiQg95RwqOvvTzIApWg2Ae2LPLUMHas9Q5N7u
z5YgDa5nGLQQC4ZyDCrGHIdV59dMX8aq6lRHEVp7y7DtFOh2SibUzuz5y5AaK8IFWpfE1V7wPR0X
GkXl6tuvueAmbi3CGoqN5BXttvCr26aC+++WD5PNEF+waekpbO40OP637CEgRyTP0gLcb1h4oi8s
nFYJvQ5L6NotzAGxXzt+iwxkyoltKuxyFxx0XRc/Yoan8aaY8Hb6sykDPm1bZMCIl5jWWA30rPtO
3PAyVvGoLiUXwQQ3+NCc2qFfFn+g4CckASlfkj8ObPOhH6bXCtLawInXAtiPf0dDEciASXhRZgIP
X1TYpkmtwxzJTqCul5zndYyNQTpiMt+wjou9I4tU5yqJ8qQWgS06ca7I3wcrKwfFDkqEQJcDIvEH
2r2DuJy9eik+cg+geUupVTXG3jWU0cAS13UnBZiOBUUXr9BonvOss2aFggz0rbPkBv07aldOUMPV
EQDonNjXzXOZvSRAwpAyRp+4Celo++tBZ9Q7vDTzagZmQQSzDGUhH7ga7cbbsKz7uW2wAj16CU9w
QVt1KIG+z6wUueQr/s3CIFqUUa+tsbYVBePxtrDDuuxzljBvoamq05tNj1UJay2Yd1xZ8rD5RNuw
L61F6ipnbnVydWhGKSbFLedJp7edjHC6wrgqEZJzGzBkOQ8Aynk67yYVorHA11hS1JcttVhaShXB
Lk+PYjSTicosSNooU1Fkoexry8X7kVvlSXN2etHofnoPSNCrOBaJU7UOKjzf0oOyhiY1mPTJ/L02
JQAtdEI3rshqT/zkKJJYNC8oCzyPbWtjwCznPq42325NTqG2LaiU9hHxahSSpP2WVh8JMUu+fILh
7f5hXSaQtR2cvbxUadjoB/qAvNv3NWLyMFLA/LC1fZbQDDCi+ycnog2qMfHOjEeUbjjsGDdF82e9
BgXycusKvG1gyGla2MtKtdQqBaF4AMkXIAFmCBxDS2SDrcXPqoje81gajmW/G8jFY8ZtPBMl7XGV
KBdn0D8ow+V9Dc33Lc+U2yQBrIyab4/KmslcQEhJAG8pf5CoivUuTwx1vcHYgTnkw7lZXpBs+K+Q
tP3m7pJUeGB6BvGU4Hn5/MmXPuKRNPQrLl8nwkpnUlw7WrgpCiqoJPvRCACw1P6t17vO5NLB1iK/
gXXxy3FmFINTG767u5pmjS+239VGwoiBlhA+bHnKEqdSPOMBzWPS9ZTfo3PptTCaUWHWc0kG/9X6
yqPE5qjHZJ46vTESQeg5gnqy1C2YF2mJuyJzpvrL6INcw3qDYFCTZCAoVNvNZsB8drQIPHaqNVot
S4tODlHK5sS9GfRLELNOzHcW0e1Tudt7UMAd98nmaBjq+UUNsUsu37mN6ajIGzm/X+UDw5SF8qnh
7ux2i2wo2WZvdxqpjVcehkqRMqtFiBZn5lTv1krtY1W3R/NHH1ULorMt+8wj0r8PxB412Jwq7wYS
LDmT1RCYeObkKuElil6wmLwIubADq3Ek4b88kCewB3Jxe0Tat/LJOAt5Q3p5cDbBF6mfoXHA1Vh9
xE/lsEMT/vjBAh5yqdUNfneOf1cRPJB1GBNd5gF8SPu/OxerljkFWru44CVZFE69VZG6OVvK+wEs
p56i4Sy6j5vtQ2okwVmCvh597jvyXQprBctUphCVAk4zruAihn2LlBeG3gYD1pQvZkxWb/8DC1vg
/aEgwdrgh7duzAUgJe5bGF05qSp5n10ELDyYpxj2lu0LTRH/Onw5ZER+4+nmBPo9UX2SLTwGfSB1
++VhHrZDhyFpE154njlqvjLGBsNeJwjgfRTLtqdmijw8dqWp4Io49AnqQpbE5ZDDbh1ug7hmeCgb
OQEPgOg4bFKE/0cQAPhEslBT7aZH2pe2o9DB7WkWsOKOOTTC2S6ScUK7+jxLFmFlyh5KJhosrunw
j2DY70svb79edi/nJ1svHnoftW02hO6pqS6U/Wk06lwJ+MbkASn+nqtg6UmP1Pw70ahXo4Cpr+gn
NxP77kHoKBSxYqrJAD6bRXc50f8WCoozMr8W2yQOanh+1HNL2e+Qh+Cv8phc2oMfloLAWyW/bmRQ
IIOq8bSUel1kObchbRZrO+G+mSNXvUTNSd3qMR2xyfppkJtoG++Iv0sq3YC9rNGOIvFOi2yMbIfv
Q3zomi6LQPGCYLtN8/LUF51sjssHrTZLsJptAQ7k4MqfaUUn4if99BAURERvopROcCMCYC0K87io
AbtL9NiIMYroM9Wq9N6E/fXjn3CnEgsFrwGBld6wjDRUpI72RM+uMjZswndAO69FfoDEdMsycrIY
W0bso1bUZL4Tf5TBYY8tH8bKXy8J51g8E8cVY4mn59TZ2n0m/WDWubut1R4UPVzSsXpj5yCJ8zpH
jx1dqFlABit2MlHofn3hCEjv6PhJ2TxkX/1OyXwI6OP6xRxYu9w228Vzqct2dOpGLvWKS6MT20Ou
WThVQuHMv+6LTyENW9GY3ERiG1IMnjej/+bxkJsmzp7+ekH3I6XmzaBV6aSFtFmrgo5q2x+1z5Pf
nK70ExqItRrAhDfpFDjoHrdAW5N030uAI3e6x/i3dorNv2WxT7dvPeD0T8APiNycA+O7KkKnkl/y
adR15ULgBnnawKos82ooY1s+6u3L9cHx+2wMNaq91lALHb03JyskTnrP+6wwU1A457szEInpKNP2
jUGEoh9Q650SgAhf1gFAS4mcIyQfeIizxAZ8WJAerzHzYNoOKvhAYNho9dpKXeTp+okwVQARxI2z
9nzQsXFHdCuS/dvb8KCKihoEaxe6nuq0StBp+g0fWTfpwctU0JuEL3IcTZGthsUJe5zp6+1hmid9
BjD/8PNFNLFd6jWUZvsG91u2TZnXY8ujbisoAZ9Cs13FCkHOrE5wheKC9ZINCDM3CE++q/rxxkyn
ei0gOsrixFcMis7Ja+G8IJC1bm9sm53owujJn57QSh5TOMGYBEQ6Qj9P9Qdjd/hscY6cfvF1Ej6o
XS2bXgeud1kgYyg8lhu+S+alLgC9tJs8k5sZ7mZxFtWXtcuz7NAVkp1Qe7SshwRE2q8mJYamXLYv
+x66Xl0rX2JOpV4AxkJYU/p0mcXBbiWYTMGC8VnXK5FJSgaWsdEHKI7UI+lcfmPaz7dMsUKs+qRZ
ODLZZKRjWq0E0u5H6GH/DmsKYqSt1dfKUu+9SptJRLZIGjIGG55Taj+97Jbvsx8SDe7wqlQheUjK
20CGf3GUrZDor8I9e02Qptlb52WeLUqSBw37E9O74BqTkagACsnqNkwtrL5hAUbUh3Q79kEuL3hv
R9WC383gvu5DioZoJ4XVoTnMS+RB7TVXbIQAN3MCZg4o0XvwNjZiIduSVntrdyOGrfl+3eWqWTm+
PgPJBGUdsQYRV/1ZoYiuD5VA1Jel6hTMSJCjQhnyazEQ8Z6Efttqe24gp1EXHbcC2X299s1bRutr
w0z9f2W3dIzB3PKrNGd4W3tKxMHSgub2tsjhFaHZhrqLOIjIJ9Q0bb8XzuJXSvbFxZHpT+YUdoMO
9DTaLfcB2vluu+B1kDs019caMslTJmxMSLtFeVLETVSMMA3fannZaoFbNzjEWDB4BcZqc7UIHGj9
8DlTTHfVMmXDow5oA9V8KOjH+0nDUFH8foFRVzZDVLlX95zGw2/600bQQzpLtbglrV761PkDlV+B
Lxvp0FCvf3O1rwmKNPgyLN4/d2AlDiTvI/g2QH5KsTEEBQf/xRoo7XjZlYKO+tizMzZQxTk4dhhx
MBxt5DyuXBLajvb9ZUZs6Dbh8uf72x8xF5UYvmmfQhZuJGqho/bUSElFqb32mIIMakiTMfVTNHfE
DlrurV9FXjaJmMbi21PDKtGZqAFSGMw/E0FO7580+0L65y3QehTHSOEYVMVRg3vxF5+Mya+bPOe9
VNwSwcy7R/yhPdawHAPxVI8x+6W2uTc8b0bWCqAanYFTsQ4i+LmiDgajTzXzmxFuKvj60BL94adb
aSFB6dgLC+RaI2uzdF/Np281bS5aBe5DPkAattAzW1IXsZfykwVuWN1592N3ml3NFVn/5bTl/6J+
p4i+mZk0CZkmP7XoRXsP6hIBR0M9+i/WpbqG4QwoOWcl0GJVX4QNKDd2SXWutnQcyD0sKzVf+phx
3IlxvKsFS4uxZESio0HWlPndZeprlDKdg6U4PYJ3LspDnPFk+rE3mT2qHf2JuH/AyWbf2k2yK6eo
26R5P6HjtA3wORoEPfKk6InCsqvjW7HAp1taIdTnpPw3G5j0pMbTqw3UJok5ZKx58hwsY2oCLlD2
AnpiqYYC3CgFhM2l3ia1PeQJSIriI1788dGcqQSFKlH4u6uKsdttZKS3qzDg+7iHs73yEqS/wmUd
wdZh1ISXD5aMIrtGCY+xxJ4Nr9lv/2leIBN0hVca2oeAV5Y2JyTyUfigLXtzyJkP0B0f5ZcyBj8r
amHReN8wq0yGWJrXHBU/LWzJH2zuc34BZg35XSSDBdVmf8Oo5BwaaR9qM9Cp5z67UKVCwI8Vu3zg
MO7c7+TVLz0yrArvObAhHRUBs1o2+Mb+/2EJFACUY39bXrZpTts1E9JCRDA6NqaIuubvclelK0Kc
DVo/cLT7QTJaQGxZKPV3yJKxI3voOaAmAoY41EDc3ooBUaIqYu5QZWJa+lcBS6kSnAj6zJkQW8D+
2GUvA458ZOo7XzSWpnWsMOX+xo/jpRHluMgY01aXWdEOOPJjEmncEAP+wfboZArxYRnUHTxeeSlJ
1+Mwugfo/gI+xcyepJ4E0AJq9VaKakQyoeu1CWhx3Cjqev/XfwMBzagrZXopHGYBgdTmeBHf5KRo
HDVWPoYr0Njdy30yAAsDz3uIcbMtegVA3ERy7O9SGR+nPSb5rykNyg3JXO0t19k0HlvPMZ6iBq3W
AyoZ3cRsABjR0QVTScbp0miGhKZIhp2rLsGYrNKWdbHxz4/RUKks6j8mcazTqyaykK7OU/8PnToa
MoAw77LgCwelD59yujon8Rci21TEkAKAsy2J8brIEk5tba7JWGA42vpID9BS759JvV0j3HIPmrka
ilBtzxpX69O8k/OkpyyqTCwSlyoQUcms0E0JntiscbJB2fkaaYA4QuqICWLd6fwb4/fTWz7zEJSq
uP2qnR7+YmraHxphxubk91cpFwQbjM/jxe3SW2ok6zf2I88ohr6g4EOBw4QgR0OfnNQSifh8f3HN
gOcK0/Bi17yA7RWOWx2raCyVU5GW14ue44KKYkZxxyIEh9US6DwfC76Quwdz5x0oTTMvZYqTxtB+
uQZo57T+CtW5CcYyL/8hIUUzXiK7QPgLlfLXmn5gKp/84bmBLyeAxFtBLOFjzxTWUtzsQxEsXbG4
Y4/vE9UvG9Aoq+gnKXaTEYz462ltd/zYynnQ7iRRCRcTzHw7glNSQ4tPB+4HDR7DHGkV7t6ZijGS
c+R5TVxbmnDmasGDKd63xwy8bR5ZeDNiH2tvc7UK3GPo6V7Ge/Ci8TUb6o1R6dWdDYIrPze3nJev
bFFIGAewrA1b4hmaYW9DA2Dm+seZhZkiGmaBhZ5+wIBR3EJ0zW3tgZps91chOJQnf8yvrMjZqXSt
K7plWHIKRuvDzIkzwwUPe4vyZ03QmQXiTSzF7wQCMQhwfrODetYt8jcXk7tSYWX5Wx1W4UuzakGH
8Yi8ANuOwPVir7Uj4I9a++v8ogjB5cUgvj3NkAGdTFg+QkAGVEVkXnkuKBtwblJKz+sa5U6A0uHG
Dmrr0TFObAfHJyfgS/THFTo96tZgtETqCYf2p88IBgHXZMOpGn8wTI1NxlVGdlEZOaKTQvLYCfJk
f9hLCd7CbixY7eM9TwS09IqMkQpIcU8oz1UZMrYHxaw+QHCAfdUh+iZtMdL4bvzjMYY3Gwqly3xo
zY0jJNFHjsLIXvlFgo7kEgBUPvQyZyWmUkHExN9wEaDSRUfdd3RQ8ceEW5TjTkwzEdPeKVnLHrOL
Em9ktDvWUiItiTtKfrOZqW5SkcE+MbfSTp3fqssBQHNVaKdzVlu90iYWmnQ6MxIYv15m5TioZ1mE
XKbJT4BEQNwUKFM9LLgYRAeoR2tvuCWm+TY/dQuqNy61vjDyVwflnuuspdIky8rPlUWHFOUXO6Vv
I4ua1mGcINKVc01v4ydQBcLzsbxT6c/D1xYJb1u46WejdcTqDqlUfe+6HvghXoxX9vPb8p5zVm2g
srojzzW/KonOCdjypdlIyLwDgHf4KN5iUBryENFdYMtzZJ7apFeacX/zBTL2yK9VzDItY0FDc9d5
EQSE2w4QfKix4BaRq/lWV3gXpoTOhEq3s2MLjsifrly180Fvvx4z7XAg4NBEZyqRGcMM8+NUTXS5
J2Qm1yymV78b7CrZHCqTdDAoX2kJKUTVRHOY47xm0HdI9VzNcaDPVvY+0zL/hDHBfE+9nGZNjTeM
5OlYaxlqphonYZcgSHR/t+lQANdj+DHQNxAqeyLPwe30i53u8vI32Qh/uX9Q2jil8pRQi2MCDPrF
Ck52Z2CgUMx0raOg/HeHqqv/f55mFxb9tzHZ6el34vczi12aPVHc2tWwQeT9tnuVbcabV3tQ0m7h
/hbtVTm3kwUQwHKE67pW5QpVYcnaLFR/MFYNkyo3iCcqbH4Qs0TVqaubimjx6nFUzPRtQh7I7sQ2
M2sgC7rQoeeDiJvgIBPU5UhziRLWfns+8zcRm+uY4j1M828fu6uIGM6Y96JtrGdi4ajbw1RrRBVN
Darl6R9sv2INexsDTUwZRp3l46KmFsLD7l8lo/geGoaX6rEFs3G38ZsoZViDZZVi92WVGJdC5mNL
tDG/30XGT5ibUvp7+eVuJ3yAwuOAftKz/7X5qk3wNM4a5WjB0rrMOgoSlBmpe602eWAdHZXRLURK
fFAYjj627GuTX1BP5rAx+B9WV/M2jnODpJBTgnpNTecUUKD0fh4xs/xkjrWJ3Tzg9cNgSqfDavkG
K/fPWY3aJ9+NmO2iErx27XGOQvbSt3HkCh/SORoyy3wOMy5PIKenJdkRXAs4DHdgOK6NzfrfC2E2
Iu2gF37EGTFWSBH62dnktqXZ30xzzNQZnEsJumZoiP5pFRK3lVKUkvj6FOnAIVRyqSedg8uGbGcW
yuBgO509FIWlcIjMKMVuxj3F7S3/e3RqHnIXmbfGf5J5E1CCsGzi0VBOSI3wtwYfC3NmOIlgnMRe
SIfM3vShNWbJRfWFN/gQOzUDUYX4HkviNT5WcWhMoJwQBCr02C+TcxqRTCyICnQiMINZvivdqDF/
hB0lnIhb51XQOxzJRlFBCtezeJD4MsAVGVJr06c2iLS/frNBW+7gUfsg6zDY2MVo9UchZ3H8C+GO
c/1N8Vw1AUrei2J6r8Zpg8dLbxwJE7cTZK36xyxckPrO7r/+VU6zTY4wnl0gOzGS0PV+/h+SisKU
HwUZiLttEvEDWqsARdY1/gYAm1/sWbENBeBHnbtgg2FktmKoa4fo+fRHKrHqoPjkVErYpUa5fHRi
c6gaGq4wlDimJKLtpk7qeKYyZX1+Kss5JPQcz7PefkMkeCJjo5mq8ZDOI4Eet6Oj9NwIRix1FERg
GdgEt+k5ZXIBhGO4Nhf9kXd0ZQ2dH4Nraqvipv7lfByNzAwcD2dQB19fihnXY82ZpgsWGdltmiA4
xaTCz3dEaDSJchsNMFIRir+sG9KQpim17BxomlQD+cRHWmCZVxoHD7BWJKwvEd/mbaaRHO0NCH8R
KQcXv73ajDf/kCbNF2ezdkWck+IkpxgUk68etIoirM4WnbhfQcACBYirc2zKZyzkHVVYN+6KqUXQ
sTJtwa106UXfD4WRl1NUuTOeaJRD1bF7/S2cIWfUu6E+ZDdY10+egBLPNPW9tTul55R9tzI9DgL4
kLCjNNPbKEhmixb58ZVRX8YlRmV2gxVc5LYYlxFBADgpEmFaZE+4vZteP5ZJT8wCEr15jjBZNU9Y
jgPixj6LloEn0e4mNPTCrYq92PhSo/90S83KOH/AjC2lc6bkLx+y6hoSAW+vRIERjUNXt0pBxBwm
vx04kN+EiIfabvL+sHcxDAjJl1ixwaRBXkpKGW6xlU3L5Mgp4MwVhiImjSBfFZVUakRj2yDuWxEe
R68RpsyrhoYFhrCzPQAsvDRVl/5Vd/LWVrNiEePEKf7cpK6kfWMumdkkjQHtgr69ykiTxgDbi/0J
Omm3r/PFQJrElzfSZ71wbsykNf2nV3xmSl6Uh9C69ONsPYIr8sYH4JGRNZSHbN8kLqXkrLJuUhtz
pt334kAF9+tbjzQKs3Hs/C9GDNugPYbtaXJjgYJxpPg+V8YRgrMyhsbkmoa+Qe/CqP56uRbkIEUi
GG3F6PoP5lAmkP4LJNMs+okAdwG1EOlumZKRByUOYbjTiR9IPPvQidG/fS03lEdmdcVHUMCj2YNB
D/3v6dc7cZqv3U2OjIxYDw16N6fdpmBoslCN95XufBWjdaRRcyg3/npeiQQPIOdYPx3Vs0rb52DQ
0aibGIF5iAnVA74xaw5p0O7KfPLB6oZuLu4FwE+KfjOfO6T+6sXzKZadcrkaRnhO0kJ3DYfqwTqQ
7JWgwZobdhZPwR0bX1kcIEdVr/CpadEoJOAHrifg1//8o3J1vMvrEyRs3ob6sDoP3SK+COcGnEiG
qRROpkHfEAWkGG05usH02wCZESvsCN5NCMnLeaPKc8Qs2NZcPh9zexFMleRTAUbIWtuhECTaU/ZA
kNOwILlh9ENcTALOHiX695Qy0VISwRXqVd4BLSYqCnYUWIIsXahMBYO7SdwxdGC3azVP+04mb2ci
/mJk7QusRpyz4VVFVUPhs7PtyZvlyKJPXNOjlzceKzZnVx3RHNTO7GGxYq5+LqWCkWDzwJPiQ7gA
9iIxcfmrzy+CMgkldXRMxv6vMPyLeAP4jGbKcBUoMou4J5kUNL4SJDVAE3DXt0+y05o2pl+iq6fG
rOkJf0xrC4f25oNdTkAStl9oqrjCEw01Ur3Lk21rxit7LPCbTibAnFWhMwFIr2tX1u7XWoxWukQV
U0rV0QQv/Tm9IoFiN66Hs+iKNR9Ey2k+LTcjBz8Vi2hWbYK5LpBcK74uXrfo+7r0urtzujYyGHQ2
Fds+H5ql++AkuHlVRhpUQSM2sqmcJ4Ig3aOW8ZF5FjhdnsJVn6UvVBk5FFtvt4YgTLr3vQK1Nn4g
qNfJ8zcirLgyR50rbzd9gDQFeUFs2k8AqVn/9nFsYz6H007dJotz6Ez+BPWjjkpzRth2VasmIRy/
7jlkpm/RjJi4CGAI7dJuHrztH0fHZa2B6vIUArICdT/dpOpG8qg3AnKf9d8l29hE3YNxZ8c0+jFP
M6EQunmb4HJFHuEfp/HfE3VuEgBElXE44VaizLhj/L4D2RVSzECxg7uP01jDVqI8itIQ/eM8mWIw
rqYbVPmk3cg6cIqO21RXgOAMOTyaS9hqcXTIMV74xCIFe9AANSoSCSJ3fNQJghkaez1NxEuBKBk4
YEecusyILajBUJOicFGfzRNOWlsZPvwt3oVmp6nHh/CNARJ3JGqbLGO6LH9B6P+Yuza7Y4/hLmN4
WDZAeZ0Rcq3MDzeTKHInamix1sbRaUfVnH9Zd7Qr7lCIJUxbu71NsI1F3eyWHd6+tzH+/K/hroFT
bnaC/1VBwoluH6mS9Z33f5zw0UcbMN93srJKHaxrAh8OQKjHzCjCeDaRGRlvWJfgiINiYgXZoeEx
K34Tn+41Y3mcNX1a0o5n+keddU9KQE9l/R6s3IYZy+bCI28C6JUVAWL+Iv3HlaY3noSASkFbU/Iz
jNADtv9CP58cZ7KLt0XOmC1IwGOniYfSZkgujYNvsvh8hLEaHnKaFnySjugtlBwepPJfMsL+5u5m
Sh1bgD9JEHxcvPxWgJdkf0pMfjae79x3uTrXHaEqf6WKha5q7XvOHjzxxBJ4MeNQT/x8yioEYQw1
nDW0aj4BnXxBM6KmfNcnE9W1h60yhdBBC4tCy3t8RfepkNkTCuzpHC6ZzVYhE64cUo1V/BY2nev0
W/MeKPVAKAvvpo5rzh18nPk++XPG9qhbk/1egzH3PBadnTv4qIZqCmTY6NhLDzBPSMYslYNnrYAm
loZ+/ZhYnEGABO7YlaREig+DMTEZ5hjTt1675nkHIbNyoaCdnnebTADg2yTHKZrWsRsl51nRFXoI
QARTRleNJdpSubIEwfCbR+mdpOnNJ5dmev7fIcvM/d0DRNGsVGSkVJ8cT7S8HTnTZsZMukQWlNqT
IHvRF3gkdJYfzn9Kw/b/4HKpxnRWFvnY8HtqftwWEbVIyC9PLMCIFE0gQxk/hqyZ+twfEeh8wcgw
5DUymL6oLrF74s+6WRcoOO0A+1iFtMyPUDkwUf4k9W33lZUyM8j2rgH8Wi0p7PXZjpVUuNywDBT+
8i147XtY5zLybqIbTMWcRrzDMyjw5H/qo76MqZjhb89wZhysmSdujcuPogcnIJw2xALbZ0F32eED
VFvTihZWWYlPxAxm3r1uYLLZcUS9ZWGV57pZXPPu/D54qJ0VjtZcy4HTzfhDZ+S5gzGuGxA1e/ro
TXr95YIRXuvv+nl7iRfVkp1ErEQGz28+u+vacC+8RGZ2rCekQUUcdKahxLEqan7yrKgVD4Wbza+M
IQ2tGEEY4+sYTXZLwzwdIhfwZxtxUUbmyHwA0fuZWH7rDjA6ThTsk+qGz6rmne3Sl0rxtFsUzoRd
dVEDRGzHHjEdq+G7Dh0WhImkSKllrEA15cwww9HPNZ/upXXonhI/F9420R36EtbWjoeq2+7jWaps
lzaf5mYEuTF83YEB2sq8Abkokz7O/YpKN9B9YiO/iKoY7MdLbwcWRYl7WhLmjNdUdFGe9YzEmN2+
LCrzqauvO89W2bgEaqIC0buHaIpTRoyMJ4OiyCCa4iFUROeSS6aQ6qfoCw/P6e+XJqbsIttnKGp5
gjauJQAJNDJOVqgE34BrlGsfvWWQAd87k8t4fTOfgWXXKMFL0hPDMfz7TOAEdtCnw/JNGPArbjhM
+QRTQnNACptH+Qn4qq7D3Bo6hBtEF3j88DKybbEIC3EWdaAFL3oBietyd1LShjLK7mwaZEojx2lO
kFN50BoMBNuFNMr2JyAb5E7eIb3S0IYKS9ZoJUSml/ckmOYHmQSrOACAWbccor4mv2mUID7CmJRu
cRP5m5FwDVxB9KlbmRMVga+0qVl6n1+Rf6L7OLL9wG+e90cCNmFjQHiJtwpeIsDUEqzdGAeDhZ3T
85kFhkwMZeZZsKREEKKB1e3s6w7siDJXdIDDpFY2C8ZYJ5+GNOONzrKLH8OlSrLkJ/OlzcQpdTvB
onmXI+oYt6vtz2aHJemhVSa5Vv9pv48j4snqiYwBnIepZxfX9sLwkin79aoTLS6onMYXIeJSyaxv
dSi8OtOg5cJhldvCpPCrwFKDAPEXWdhFRDXeQencs7d0YC9TZ21n4xdOgKaJWatdTvcqi9Zci7wY
OUhKhHezRZCHPpuJg13chj070OrRRxeFIOSD5s7mCbOatGWJ9ah+4Awt4Fn20gwmpd21llqGhNjp
A6iIyHdsu4yXUAWMcFyu+JSKNKCp5ylE23OfWLE9KGc6fZosg0AdOMgOf/E9b0mqRXxaqTj4shZL
fgTdi8vWgZfbcnJvDsV5ooIZVjhmWB1mIQr/nb60aQHXHFYzytI6CoCG1ZSyIGk5kjtJAn7FAF/A
Nc1TKL1PfayIFIIQVRaAAdEzfpxo0u6FW18/5KJvuo5204kd4IRfoYKLZH/97GuJFZDozJw9ZJbY
lrrFLcc8qht7uvOPLpoze0wNAepbLPF61eROsI5HVT4c+QtLHUF9alz+UT4z/LDt1iJUKaEj1fUV
P5DQqUaM6Oe/iNk4CT7s6QsqH4weqpbruX0ZWrrdghdTQSR3JBQwzFh633fCYDcxhL3yTghbYGtv
MvDOgcZ+p5qEXxSFp6pVdjA/j4c/Rl2U1JpVCw1vhneLVPp4rvz6kaAMPQknyqZAjJ2MNAxj2z20
nSmafLNvO38lGhxMgGJNYiA2azKLvyiMo6AkUlwraJiy8LRLUmu8lr4LOMSgS++nM/kU72cqNG2W
UdjCfyjg2P0jDmj6WWNCjHs/pn3oimqhKgFSiW92x6sVc6GUJxWGzHQ/KoRvg9w2gQS5jSeSCA+e
RXFbqPFhA2d8/Nr82PbLyux8RdgijJgYLPSMN3mGCNp+qD9kBZkZussFepNN0H5fQGRRAyksvrby
hBfzkFB2XgOTZsDP8Id4/R/5IWuq/ZMjppZYBBEqWPlyLlD/YNG4/u1S1z+0arCgkcP7OKYsW1yT
WfW7/7aVkup51ztmPXEkERATsNrezQJYzyA2zloBTnZLth9cMEysdwt1HVPx/kxC9F3UPyLbYPRz
D6apPQv80/akqNLcYCqYn6Tmq9NYlOGagFGC3ceDvhC6LnfIXS1pjKRfRZbirx3Maw6ijV5UjwED
exnWbyndfhHxDQsKxCFcuu+tDeROsRAzOXX3L/jDr2kfuDIhJ3cvUPoeylQpGXlrIVPIfHWand4F
Vp2nAPatDaCBNq86HLlqrb74UQQvrwPgee0oVUWHLTXrUfjNMWC+1dMOQoZGXmu3YVxlR2QtMFAw
4LGp3lOVVKk9cOUos8Kyw0jOV0+CmY7QRdpYZqUnApxohogw9u2mUDKOK09oQNoz+B3M2H2/JNXQ
AYmwBwUTpmxS77TB+0AG5rrljWl8Tb7H42KoMZ5FBvmcn0qeWQoNKDmkHAZe7UqhBFsoccHTzRon
ciQ6mWz1XZOsjFKGmay3PKSo8BlJBUYc+2j45xIJX3ep0UgnixWzkpI7WEZNxcSW0mC3yLxfjvZs
7rF3+BR11OW4rNKkhspncGLG/dEdjfusJvZAGB3V/PAOj05E9+W9AZhwL8vp8FP9IXg5vsz4RWNP
BVASFhLVqBwiM7gkUzQC1NCq3kNqI/iV8/BRUpFm2ozoszVtUtd7vE1QiznAKrcdLw6qnMvqYh+i
ghcXV0d6O2+jZoQ4/LmlFH5X3zVDonRhG6Ika3AF+qVE2fK3FSIO7edyvD8MBJHdMlV1XR6OY5fx
/wi0eZznaPXPTP4xMrDhwNu3n8qXzub6bNBEVHbZcE/xTTgqwSog+UI2YjLwU6GUNqBHWD7ilwNn
VtJMSK8xhISnlOXcsIJwy7CBAVC6jFDytt4AmnM9WDSzalWJd/uJY8IiaJFz7pB7cyfumlAkcU+6
Bat9CUA6PlSPHScwjccbAttzCuMpxldE00Li4aKUE0YaHcTOTTJDJFzTtk9OXKIQIy1gvDYT0nL3
S0rMd3sSnX9Cc7wDLnL2+ipEMSsQMleqtJwLMrnEfNBhi+wI48SnlWCW4lm4yzrUhiU3+dFwREI4
BINprLQkiWOV2xraDYss0DM+53q22MXA/BnzulJVcIowej/ShLtWTJeLTtsADvLfol1LRiZNGmc3
NDYEOWr5HkXinm3Po7jKK/x0KoZ3c6cTmdJmV/PUTZKgnnAqMmWQJeddDGKBVPSlA/O5UtSQOEpQ
dFX+XI3e4/VnusOqEsChRBKQt338N+lHKYFIPig1HwQsizhml7kOgG6xU4TNod6K3CwmLRW0roD0
UQHLqYZOx/jFFuNuV9bQH8+UyWVbRnKHQgh7zSZP9lwUjCMFyTLbZrzKnJEFjIeJst7AX2hP898I
cbIgCBp10oeaIReDxmPcWFtdAuEP0WS+IsCEgk9iUdcXebZs+oZXbGQyJNaWoZgFbQxXcKX7vtAr
nM6H7Szz2vXc4TfStqBmp38BeL8HLOvk3o/g/k4WAU6thi0PRFiO+9lnlI3v7pIXfZpFgF2UwzXb
pPi2wC8Ib5CFENqhUS31yc7TXRFBjlNxToM/D9FOtX4aJAAetk17Rd3RBn0JZBT1CXPWc81dtkEa
tmnSdTtB3nvRqwifYCm5/D+kI6eagvRtyVRqen+yD9k8bEUdcPQvbwStaGTSue9kCHxDNmmNWvg+
un55dL9B29Hl0vzTRfqPmV6LmBNWPtBIFLhTfNJClLzCU1GlMh5sH6nCoBdPyjyIMjoxRXbtetoj
rrrDNPgX/yAUcMDN3ybXcd+QZ/DVY5eBH4zdoT9j2nIe66j+8iT9bUq3lIXVkfOAEypoKxVZ3gEp
XIlW+1SIZ7EMnrTvgDE4aWS4hnGzSlxz7qbLWlAAEN+Ul0wK9UiH5K/T3/YsaqEcbZEFJ4glH08I
3gLWCtPpdy5ORVZPtI8dfeumGnUQK0S5x4OoCP4DrQ0uG5lGpCjsV6B3dhB8VFdL+5fhPoI7aIk1
fMKfjDaMa14iLgkbOqHrD+jw/eDsKwBwJ7PI5eMaK4reOWu2ft36RfyOyhcTn9c1ftVh8BU/ytPB
8vbQ5S9E+FvFctprPXmiLp+9jupVNO5G2m/DY6hFjNCIcGAU9hNbw4sQnutNRmsVoTZowIxQRRi1
KGgRJUn+mVylYw6gMdilQm9YTBi8Wr7agiMS1pjd/W6ZZLys7gVpkkLVfT6ERByuuWoM/jf9uucZ
Rx979htTVyg710sA6heXMDFzS8D6XT77x6+D0I/C47seinyZrf20H6JVkQnsV5TWoCLVNn8kQIYL
Na8QC0xx2+PStu3jm53HGFyKHIQdSMETYrdkPK6nO6OwswJuUL28oz+K2R+0v76T06q5jk/DeNlW
aPe7jpAirx/kR2QYsYBhpKV/YK08q5Xm87mptrcu0yec4Bk2lqZfaClexPedgPkZd5RovmbhKVeS
4ZmL4luvJmQ8TotI3P92S7uo74amgMz14p6jp+AsnixgRppEOuTI9W+zSj3Av3mCGFIrnEmuf/B2
uU5NxdiFKBgVfwPEmx1Lm08HG+QnUpQ4EUY2Eb4BS0LVjzgHfQGuDYzMAs7L1Fxv+vwyjV681+bo
xZHHoluU3bjGM2Cp5z1FRxfVzpFIUQc49TZe2UWYxoeK1yL7CWZI81eKzDKqfbCvpvB1qsaCPl1Y
VahyXvbLL4u/iofc/oH1ThTdeRcHIh1vs07KJ61uwD6Dfng0AjdFwqlDOAfE/Zi9ARmSUhAIyeYo
crc8eQbwg7VYQpi9qMV57IzhstOuiRnzu4Ijob76+N5L9mDyPTY3lDCuq8gkPtNEYKAJDaxl2tXU
XV7dVOwXPlFs2qhbbgwQEnmn5t0RXNX3vL7Rihf3Tn2Yvn01nsMorTvv+ZqKyHpJGCoffpspJ0ga
zwvDDfUSqXoxXPt+cWh1eKPJAEo7J3g1fAriiYBj1gvY3XCwE/vd/3LHVSDAjZn3YJrHMFFjvY92
tFp1aka2iZvoqSG8i24BVMys5cWfrbgb8aPPoONQIJLxmf9MSlev29jTpW9fcdHeAkotdELl8nFx
4+sfoNOtbgmaaCAHpKtcXifrksUCwSJxZS+ohc9EZ9yilWV2U+mYg2R9/iX9QwgbcnDU2LNUy+z9
cWn60/8LnCrFYVsnPYR+ragtHTo7ErfCnAcZHgVHosQvR2O7VnDx9VRSqfgv7OPg4agExmXQBjVx
CfG64Clwh2wOid2gEdXQHaozr5vgs6NYV/DWKWy1p9r5dm+bT9eTnJUXT/lrRbchrZJr2NDtocbY
LF+apTB/kgOcc1GfrTkytjtWNjCswnVNeQuyMycNLkSpM5vHhVj2AAkKysl77JxCSbx84eDx+1ca
0C/uBLTzVxx+e1jToTC+286m8uWl6n3MFBYI0w7Op36BUjuPeWzpTEmvQZquIQ4RlFXytQ+vV24I
oY5H/4rGmhsvbTSoK/FWf8iH3wULT+aMY3Ps5BK9NOzMuHFnAq+ZO3+ZIAgIm11xhOlLybxBz4dn
liVsGTK2OFlcttzg5WyLVsTtkMp3Y2aRfKfbtOLejc4rTJH+SNq148NPvJKAGKM48RQMw4062F1P
YNM4Yzq41mpZVmoc2TJdujlmo4ZbYTvV9zp0jHraj2Xrn6IfYd2A2ota//csri8t05bfRJEB3ull
ZCXdI1U3Qx1CQIShwtDf+h6wzIKWTXKPPOOOJM1p5spZw60laxd075hc+M4BDvLholTpMr2sWCcv
KLcrIpcPGG9LzY72Rhvr4xDtZJZSkHnlRPTQ2a3na7WdaQDxMm0w/tkGj+SR4IrCl8K2OUbLUAj7
qUmKV4NkmU+31fMPlaafH5bTlicEdcIwxTZQD9ay/AtiJ/G99axUX1VsVELVBMH0KUownO/m7J3z
F8tOiiVeMsB1IsaWkihkGPie56eYnvqGtD/W9CNUUA7CZIbVRhWCEb4yHOJ89gvwYsEXb/b9f0dY
dbj/0GYO5a+NmcFAryzu8hdSnIK8KgMu8SDE9F49aMg5gscOscNHgn4M0s1VS3afLi2NykWmiRBN
uyXhcUBYIrNpgNcaA02ELwMPzFnuabsnWkZd8r+PiqrcIBD1ztMrntl7qXlMY8HJQx2ypfAU6dHj
adsGI8W/VhMrkZDqO18pMq/MJQ2hbsl30Ja/GzRNKhyQgzalCpk1Wx64qDgCF2Cr0NC3Nq4JsOXB
8brCEjJ4AxVEinme0FjH6C0Gu6AQGCthmu6z98+CF/5dMdldMK+4iQzXAYK9DDcz6AmhGD5hJrmp
GoO6hRfFYXAb9kEq9oUupqx4arE2W3Gw5MTz1MmaNI+PSdVcT1eNDYNx2+CFS1E4Qpk+8t3+3fnX
Ju8HpQ+EegW9iV/dZzYeEXgAJenYkEBvtaMKgNupuFzGg7+XvViHIPyY0eQFfbDfFbgpArN8GEiu
bwfy58cx1I7JCn4biqXoWlvH2XmABCGM0FYIs56OW4PjEjEamO6VhA2iMDemnerIebC2lbi8+j2A
vRL27DbAFDJRLJDRLrX5y4h0jtll0IWCVZt3zJZGlrOeAEbaSZ/devkbrQ8ch3EZ5VBC372b0ds/
5lurbXIqng8wgRrFlDBJfg0k3pL9SrWOYLJslW83o9jzrnRdWYevcuJb2CJvZ5LDIox5oVZtMNUo
8jTV97LHto1x3o20QBRrX+WsSLcfLdDoLSuwfKgg1UHj+tmmsun2UFalesiVgXsDy1g7NZqILh7V
RwMCFpdDGNniqhNPUihN9aRNEa/fVe9qlyDss/fS2ejjFDh7AviAPzZDrOcyjNhQx20zgvEJ09al
CXY0Eviba/BBUIWAKeWmJqdbQ6MnJQX59MivRe8XIzImWa783vzh0fUTMPUVvRLEAuJqy4ozEtrI
v0L0SKDanRg6z3PI4WSbEAAFRWV37pAqiWOHgDs11YzNHFuZrRWpnzZ2lhLbpb0n43e3iP3o3ur3
wEgghWDqm1IALm9Ltvgf6Gb3V2/wf1q1lEBCPTlMka+ZeJf+g2jjqabtYFhLWCdRiAcan+Sjl45L
DW2amWpIb9T8J/g2cZZJqFUIBEgmNOyvhZdZDhNnnNQVEhYTcJ7QWlfrUsczFoLiz16RfwgIBLxH
FLua6LKOSBS5WU7vglCe9fNOTO0FVz+RubOChfj9M1Ydd5kjdPbExTY3812Gp/yfA3t5iooYVZ1l
puhMa2bcIjbpzBSnjOH1KpXLhcnqMbcSF+CDgtWmIKxtJlbqBrF/4A6/pGR3dVLn+4LmwfMTshpG
OopAL5/4QHeKNzDRG8DwYWIi/y5VCfQ8Lnv8BXwqzlRJDQqZLTynWvWAb7El5qgwDo8uybY5gko2
jPNx89gSJbIywrKip5I9wiPFiT7QvJ0rowD12B14qIY8qdBJk6o/cBxfCIr7bwapyYFSGqJurw15
gNjR4MSulkRtlr1LBbdTT1plQkD3BjfLvrtFVx2chSXtHq12FyMWLGil0SZsIKmPlIr7J6ek+fv4
A4XV7sqY+YinvYbSJqcA/crUviwHgsEwtvemlY6ag3HEtD8W0KIzHTKm6rdKE5NTd4+b4HYUjfc5
d+pyiqp6HFsbtrBjzfIEWWRQBXbF0yuYrsG+AvvYAGE6jO/xjtjHodomJ1StjpRdnCJktmyB3Yn8
QugaXoDhmwnJFQCIrtWL+wr22hXjYfPiKpxOc4wm+InflmR2nAVC3bmffA6HbjTMOO+JdkiVINi0
SHSQhQLC29mbFtfQrCGWQ29XhspjYVBATBHoCT16pXntzLQWhkyF7nLfw9VY/5s/E/aZ78lijN/a
gqRNyzZZqHb1s/aO9CC5sMqP1lOEs+jPUyGp/+B/BuiGQKDNmW4MHD2Pciel+DBXJXPMwxArq9f1
Y7ednivRCE32iE1kyGqSki9PUf7bQKUa6iiTUU5I2ISOMJEen4YfW7dmfKAoTBf3OQcOQe0zh6wg
9TTmIJtO98wbaiQf2SYY/RWygem6HUbhXRk6u12i7yHSoht+elYQiI7InVUkzoPyzDfxF+SYGSxC
B0+u8But8b5QLXkJsZ35Rk8hpKE5CbrzT1KhzumL147xjY+1ia0p9mulF/7JTxgJ4vyAq5qp+HuS
AX2kZYjkKb3h9iPWSXLy2M9ABhhM4vI6rf5VDIdMe6pGFPHX9djlv3n08kcu2XDN590qB/MGLEaf
N/c4lvxO3eAtGY6Cy/a+EcWyb0MmDbp2x143cTvkc5Y2Wq0qV6c3V6lKhbFIatcJl4TQMXBdsQiA
2CvVfK4BgKaoTa3x6hY7ic5E3gOgErjZI4g1vEm1x9o+xewHQVR1DyrPSh0PVuQ8jzoLJGfWauwL
4/cZSeTBralWI77Q8YndO09F+BAlk4QaCM9juU6ZFNMRGZr7jqYyzxKfhW8TfsK6BHZq5PkiRFrJ
6BHA4E+zn/os1CBe4QaN+8YM0fN6++xDAtc+w+txUWb+nufp3w06FaWyd2P9iavrMgbrLdL6VjQA
ktYdCsw1o7O48cp2o29u7v92c+05vT0w2RayQZKiHPaeA+QCbajApi6D8WOs6pdGNrEc1dkb2yNi
tAQ9kXYMpAjYBjhZKZi7UN2eYOhUjcjVXIobr0rIy4xfcgghteoT4yHGAbLuD/dS66PMLTjouN6Q
Jf7Hcd5m/EmXcajpwnon5WRFJYosWk6SJhxWu1yqzCqeyKXBk/GDSddwSYWProIuvi9mD8QZpaeW
JWNVlgIlfj03aDAn+9jbmex6oOZj4NeBeKep3ueuMuaJP+ItdKOkO3D7m8Jnzpmmu/gRDqFIN6J5
L8X6mpV66TG5N79sfrSK85nJLfoWp4TJ6eJhRWXpFp47/H4S39bCt2Y23AtTgqddSizen06TFmLg
cmcq7HxH6sJ2nRRc3JSnsdCMGPLmlfYAxvKr+EybBmsB/IubSu72sCHI4Z+x2oKXYsw2qiH+hGKB
t6phjLDplyxAJfqZF8ASuVLSpji46SFENsHWKRV0UPGW8+bqTmmhbBxWSKk4KI58+Z4PYLq5Bxzo
pK4jY3C9Fdw0P2a7kWS9VDOFcZZ53nSgilMs6aLfrrO5MamZUxTugkyXqKntNwYskZ+cMbwQXX+T
LDIihFLhtPA4Wv21zKTJh0DQSdoGUGdRVRkD4NIIInyGKgF5LfpQNqU3Bq0wtrsZ4W7GcVob5BW7
i+OjzVdhWrd9bzjxhE60Xk5nBl2s+oPyknPieeaLTMd+u/Jq+d3F9msRYtKsluw5KLfWUun7uBRM
Yy/eb2uzdMNEQmlE//ds2oiVI26JbmH/WrxaiogFA/VwfxqhYodlTT/zxX3KL6oJq8r2IEYkXYi0
dfqu5f7r7b13QcN3dV66V+luWDlNekEkHkEi0HyCv8EayMqrhcMSPNOZiUc1dLQTuq7Wj+QHOM5o
znDMC5wNRmAaLlFPupeCjjZrfSyS89kILCCxhuDO653aH8bjx0E0EgJcHzkOESYqRopuzgWYKfpD
q3dBc/sIIQuuQnc1Ngen8Zfjxkez58nEp+9l1H8gEHga59kH757vYDN2XBQtbkHoQrQTvdxjj2Mp
1lHxz+n/7tm19+Yl+1oOs3cRIg9YnST2bofeOrnrl2o6Ai/wfBFVydIbicWxoXoIsaoV4pBKzgvb
FKZ26GSCtz3AWl4gKFHl7J2w8uOa4XB8A840vX6T9yCN/CEbYmfOT6Y/vay883NWDymLish2L8I4
HTnCBs2UtKFgDHQTYPcnXM6gZtu9FxvboTlM4Ew0Ya8huy2CyVqgGHJvgvKudtQlrdtUKo6QT5Yo
hpk6hhcT/Vunwl3kSp2gK9gaKnFFnw7tssmif2q9tL+7ihrRQfSQFR31q3hRYCYrMGDPwu4DN8u6
ok/kNJXs8uu2gJ6AgUiIe5jFEUv4YIMIed3SFm/69K6kflXSra0YVb3wuwsnrT8k+m22rjpt/kYf
pnWYIo+B49vs3y3Z/WFXP4nZ4xTz+/7MgD4VvB/N4xUIzgSy2BFaHJMVADQOyEMFp9gpxa4ELeBm
+B9dYxm65kH/zvbDEvfd7WWz1s+UTtQopK5D3N1z8/2aAc1gcr4QTs/27gfAdF7c9lR0ekvTXFeV
ljbVepw0wdPBTgTai99sEO0uK5lP4hNVOwvpxvMUXZEXQQQ3/AM0iYxg6RTfcLvoR7Ty/VWClq2Y
NrQTVwp9GYkdiAUYAsE7bLiSwSvlx7JaPmIO11g+78fyoVT5mRYlH/SkqoI0Vq+gKBpac/XTgm0Z
aYKS+eVC0Vp/WlBljCTr/nbre6wbabcWEAhQ3HD7AZNuTyVIKb478+3wXm9TGNfHRhiTmkJUSZqO
SKRBAmjv17iI79eerQHfM5CzEpqaFOygH/tAA1MRpIjvGQLE9T0vtapgyafP5JdX3m3b4hPyIgME
8zJ1SICYbFE9J9ycfhG7nsT07tr5smQ370Tz1Q2c7You/98kAry1THUJsvFbh1pOLTkglZ2d0+2c
Ni2gS5ndbA/ytB0+b6o4THCABowgDcBa33jfyTWeJfk141LoJpHw2UCVVJVuiKMsuxuxFTojAXwL
Scx60qL6n9skYrlxbbF4wxnf6SIS7jf4jnUpwK7xHf1t/K6EjU5XAEJa2jv6Wo1ZfQSpHPVX8M3N
yIPbiFnOhPUxU+X2v7/SLNSe8z0f5VPIi9sAWHQEFihHjRjQrNh0gazWM8+fZQT0KVtPFxfVR8d+
oPFEsjakF28kFqZ3JFpU4FPSHTmaY8BI9vcK+y7SaW3koJzFcIeQyelvC7CKvkkEvnVSugpBO/2O
BBpVh8COR74vi8KaPpP+6CBr2JHdkwqfDluBuptpc/WenmJpytHX4AtMR4Yzu+mXI1wjIrLT6edy
Quo/xeUb5qemXFH0cTNe/8gUgGwPmctZTfCs2UfjgffI+rAUu9nMpc/9t/AR0qEeNtxTTEUHIp9T
4PgV4vL+bp1deSyKaVMQIJ5FctBmWX6Yh8WdxQQFjFvnmEW7f2jOuCkY17pkUAF3YMYnnx+3K6vz
4q/ez8SbJbR4d5BR03YIWcvq8JmNVLgDJ0I3VBAO89xSLIYaN7m96224ei6qBOSeXzn9191T3MTf
0UxX9ezTmjEoF9wm7+d8HpQIC/FO1UlGI5VJJiI21bRL5kLYC8qtILrPhW7i8HWy3tA7IMIBKEqT
KXJa+/CD3p6VtMsCh5hlSEH1MNmZXH+15ZXGhnzwfB/gbc9x96fICa5C28N58cEp8ssHNXpemPFE
y+ogbEzlP85vOB8Gc7JLH/vWBN5sXpPnZKSq8/OeSjNgjA4BqPPuP1Z2Y4kYL1VALtaZ51bFeQoI
S7QkpJtDabsNOgsvs5iMaOCwLvHK0cKoz3vbX3/FtNdAvrhB20EzxJTpFf1reRPEDnjNCqASF9kO
18tql/kGuRE2khA2Mqv5CuH+KIXcoU9eA0E+EJ9+GQMzngmgRatyPse46DA6slOCIL7uSdY87WDU
XifkLKnLbwCF2UOpOL/9W4cgVqOICoByEFWQ5JeKdilPuKI54fCd4O5A7REvHvBQQ9xdd2YWv4Li
AmGreCKeOD1wWwp4bXBEM/hgPmfCFbOdIRLkpJINEEAYl35YKmUD7S4rp1C+96rcnaNHQO+mjI9x
yYQRZfErAA+3hSkwLTtRG/OUUA1SNQOI2vsv5drsJf2cABJ7OQMf6sOC9AV/sZhF6ni1/11vQFR6
O1a+LhCQuc3FOiYFNn8ewgK2nfqdpt7CBRhCuRZ4bb2IE1zeGGnMF3c63IwxoeAcbLH3lIhfjd1k
rx0h0be2sk5ZgQuvJVE1LNdjELY69SPVFMp/HI6DL2gzzHUighHciZfwWi4P2rWKAeIFws6S2dht
MYk0lb92hNdCvs0cJ4NaOSP2no3Jg0lsmYb+ZBHqj90HXs0dpe0H6MnVlA9KLv/RPK9juSbonAsC
Jumg4FJ4Kiz9JCMHJcV+8RlUg6yK8Jx7yFoCBhR5/UGr2Pk5xp2s7kPUNZh8l1TY8TzgwePD4vUa
VsQR2tlKsrpAgACR7ZKASPCb2f5bKXyJxXUYYlVQyJy2UZy14id0418XDgL0EdyXdKZlz9ahdL7g
9G9CSn68NHGJzP+aPFy3GL6UVpCodH3VY4SA0Sm/tULx3UV2eY5SXeqxWH5HH4n9+R0icn962mC/
I1xZSBu9f18PE4gO8Kj3rGPlsUA7p9bO/pLtcHqsWDebFkwrSIhVV30LIWqktHpzB8IEjrZ2RTQp
2aapqevFXDxSZNTv1zmIfwVX9jMrVEhzbCWfcX/ReogVuV+U2N102A1XiozaJOEwFV4mPBh7Oe5H
9I61W2D9/SsN395hKj0IjOHX0sxnSAVrvmqHu6Mejjo6xHLVZlDfQAMKiF8iy1MomWPBDCn5KQiG
srHL7uPIKNKxExgRXrHDxG+g7kTWoMhO0Zjjfsq5AFjch5+paXYgAxmyTjz+iGd67r2Fip/Awlua
uL6nvncGE3FU28Wn4C2NpUiIPxRSsiUD4C6A7TDOIQUU0lZPuYfratEfQOuLSj//I4NTZWDPGfCw
sLYNBCv/LyiSl05/mHpLdQDmP9VVoje0eHUb5jum55EyJbCFS5OFHRefyJEoyUCjJ5LuC4qY5Yjw
fXuRW8ZYz5WcKZR5UWDBoxqpAWNj3mapcYJAjFCDdl/PzbY6V7Gb17dgk2+s7jTcvThKqsM1fiS/
jSbZinOPFNCIn1UGIsfYKqsxmlO4JeR4ChwFEsmB/E4nb8lEK0C4Y+ZmwP2ZvwtQ44vvAN+ugmOD
aEIhfedEzauJie929f4aqt34yMczqj/hKtnDnl0x3Qxmcdp/Xs+TzyKBmOrp6BCfdBDJ4zHMzpNf
Iv8w2leJFkOUsIdPkuyPzyJ58QpeLtobLsKl63YtiVilI6zsyCRlgzeVky/FKrJ9vXOVRu7u5Xql
Skf+dLjxbZfZ6qAkNR4Vvm75T0xj+As0+Qku8uYlLRPnrTxTE7OEc6IchFVPJutUHQeCQcdXb1Ml
t32uE0epXyOQtQmuX26/zW0/pIIhEbudvs6OlsCyInU2cqD0o97DrPv+UfEA7et5PH2MLgZMQx+D
2Z+5ugXZGUo7bnpIoF0jpHfKnLmeDKC/JC8Ip4dWpjvSduGQlWV8YiqrvixZygNgRimO+WgwJ2QJ
lTtJuGzt1wl14Rpe+xrWyswBG7DsMOYP1TitL8NS5Sfi6h2QoQXKLLkJqcVHq56Yu7MWMf7dTsTL
uNJXaYqu8EiygxG2R4mTVbnzN9xkTuQ+GwJzN8kaWijLSfSmaGqoIpye5Ym+sbshSoTgAkei8JUc
G91EWnS2aQNYHmCKQ/rypNxwhXEIQPfh/vfulB8XTqvnXLrs3kcbNR6gulWc5+2DbXT21+qj5aNt
Rh5qmjlDqUpQ+ctxS2QI3STya3ZaqXDgm8nn+87P6y5/W6ci2f1mycj8o5dz1trej9mUpfQUirLu
YD3Q0ht0QYbxFYR14MiNYECvz5wSatpXl5CiZstOBGveL4w4nC2QUobHs296snlYC02z/2OX6DNe
zrGaGag2bvQq3rqTZMm2NosemYv7NTbi8B2eY32DXZdtbpA1VRcrALnZNSrHn4Lt3j/aeda2R6ho
MEMRS00UACUzAGtPfdEjkqgyvzIVoiODqU2UXJXFcg9ToM1PiAMUtkWDpYKseZShA2OM/IYa0nHA
AXXfn2xWTDG8AHpUmNTq4tLGyUpWMAI3rh0vIVEchJVOfq1k4y+pSee5/ulUYZvoZdifJsPEvAj3
PfbIsBwHCZB47HO0jX+iSiRExToTaUqoxjIdIVYht3AzQ9XgYTWwPQj/qJe9plQoV5L72cAKsH49
Ld3KGvvR3GFAIyWhP1tpdXFUf3nO94JS5h+03958sIWYZewff+Owtg8fdz+zEkLzkoVO4DjmJ/4R
muP4bLEREHicav3xuzxb0upBOHGd+WmP6UAhtczOsjeQO7dVN6uyO9eBXVnD0JxE2v4esAAIezob
QbtfZcJeVy4DcL/N3RR8/v4KZ4ldSjWJSIrjfY46QAtkCmPp+ZxZADEpTOKl4ZRCQWtQpi2/0rBH
UoTzl556G9qNXr9i+xIjVgedFQl62X3lIwfSQ1Xx1my6LXKrJ6AfX4KUdC0yCxtl5ucXpCWa663g
rzWexbHGwiqegpm3JaWAKyGNqASzubuyo1JxQTEnJFj6Eu+IgUASW0xguHpHKWmOGvzUH4gUhnfv
qGdwN8qzkW32YTGukBr/I4MFmCn8rjROW32DVW6ELvsigL1RgoeG2g7O22y5QKvZEZdNUl4hDznL
tFOF0AIwz9E/g5D8DUuyujMQ8Tkj5GsRIL2LgxcPEDNpHXHuN9N8+r8N4LoMp8r54NLHC22iF/Df
9x21tXQPcj5YZBq1XHaa2LirIFmnoc0MES8Oq4Js1AHNQoLApEb/qOD0F7fHSdxpUvuMKr4uGsSW
lblVu0uorlRQ1HiUQSAPSZhNhGWLOBJlj69J2gfmRraqS5FbgtnaBKsVR07ds/Dp6vwbLVA3jHaM
SnfbdTHzwrFynW2cqi75NzUcIuUeN2Aq7+4/mNwL/Enh5ZnwF0Y+LeI1q4xB0ClkcsPgjRaa9mlD
VOBp5dclgVLSzheRUCDfhlRNyOQOOhAepY4mjnk5WZEEUURILCykmHMgsNBKMlow/8LAelbpUPPK
aLcNS45Yp1piMTuhx7RnnhmC+melR+x6DN88s9q8dtPA3lyZe8Szji8IaCCD3Xe30HDcLO/KXNZh
4xTA2ds6j9HGyI6Qg1LuTRs28sicC1xTVvkKMhzjZUM+07dKWn4BeZp5HsICLee6TUdICD/KmK1A
p3zM0jC4dYn9UJ4wgKcKbxY2SieQg35wvAGJS66d5sdJE8801cmuRL22iROCpRkVQPv69WtAi/gu
NLzxX7Sr+WcSRcox2YVkVRRbZPe2mE3IJC8VqN2We9Xz9leadXYrOdbqcaX5u4F7APQM2CPp1QVV
SVZtgJGsWwY/H+ZlNwnHriFRUHbyHxpk73fp2/F6Bjwys7YgrmMrDAlY6CXc+AY/L2n8WtvNFDn2
JMaOTB0mR781fhQvlq+P6e3NoJWk1wYYDeabAafOAHriIit7GgBlHu9iqcpgMYVSYDWNDD481kY0
rpH8r9dQu7pBHn6A8o3EShyPDOYQQYVO8V56VhO3toayIc0g1BhGhQnVhEEo7rX5U2bVF5zPzpaE
q7xOd1zedRnFAJY52y1uQixO8gUqi73I0M9PnsjG8bLXhDamXjt3onfkaM2h1wiMrHwK+pj27dhH
+ZrF9/vkB14F1HCir/S2/xjA+StKaAN2GXfxxt1n65WyPIqCa9gWfJZqDlIGGEXALRyz418JIW5F
oYEbXKEYSBQK4rIb32MRsnf2sARoW9rT0BEd6C7y1LCDnCZNHd/sgETBkmhziK7KOl6x0/8rqyWE
ZdChmVHxLZnocSzNwhTR8oYgE4kysYueA2ej5ymMFPO0M5UUDHDPLElDMLzittuUUYYF0hBR18Iy
BLHuWHsaP8pQheKPf8HzzfPXdjN6ByyQOa9i6YJO7VZHuMJPN3mIh1qLugfD/w7v6CqFnMFlmEHA
TXM8wJ2uyCxtVt5ha6Yzj7unfzbFZ91EsBUfbOBSWQic8MT3UYwAXQ25aHW0tQik3CSZX92salXS
o7h7wFaVh94/FwwK55sH15U/gMDIVXBaAEGU5NJrNljv/K2Z7CfhYhvNwc1wQZEwoxA6rFANuqDs
FXP8yvWmwflFwtQVVY2Neq+urtE8Zjpo/UPUqGFB2BjIOlIspEiGKQwFqeOJm9C1NMT0t2tDMC3a
z1mg6DXk1F5HnkDO06WVcfoS5rYcTTW0yTaqjXhJJCXgOZvcrREeZKxE4YC2Qmf5wWH9Obtg9BkL
+zZWwna1xMbesvOcYOMK4nE55CJPBWAfYUpyAuOVVsNAXGtEcjHkJRPJcD/l155iAr1dXSvaHc1N
jFOvMlOGwe4Ho1U/HIjXELAID3jZQBRqVbT8Z8PVQmzZRxlsFuBXbQN13dNkLXfFRe3DAXzQdpJE
hajyh1TNxIDg6jnibX0/TZ1lXQuw9V4oyWnH9x+O4PMrYdJ9kugfs2Yi4SKa/IehSF8VOkJTxuJU
hKsww6oNsa5/qVBTIr4wt1enELJ0Pv8ia5DoXCAoU1husLyyayxdo2p63TWz0pBh8Ga7KdinxRA6
gN90boWrnVz71683wrnuHRhjDuNlLkv85/Iy1sAl5R3Y2xGeZRjQjEQZnuI6O1+AwgAEc3ihAUVP
qe4Au0mu2VpqMPLiXQDxTJe0Fsiv+CSrzcEL9Wj3BcsVsy0BhowYRlIVZjR6JN7gl5VBv3xMk1ej
1h6sG021gBJnm3+2K0TLE+faPc6r5s+A8BMDRvbzFU5NhrOAO+AUD0fP3Iy+sCYBPEOehlt/gCIg
2d0oVjf+UghT0tSpHQeC0kY8zApaDL99k22r3CboMPAew0Tls0FT1GjX56k/vxxNJEZu428p0zAs
TgfdxM5fqRmRC1e2Q4E4IRwSClZG3JVt5sEKjTk1RXuts/e+2gnMHDdK3kyURHaZBiEjO9lqQ4R9
zDCWkC9qsoXDxG0K6sHnH8ktRXdepli+kBwxtNLXVeBZnez7WkK4XVe+icKYepM3vM3xQpnA6yJV
dW3VmtmJaqGMZdyl0QoUGp3y3V66kuWz6IhMrksHeBM0ewx+A6iztmmV5zmyvSfsbScmk8+c597F
Uy/ePE0kDZuIFlUlvXj87dHSHK8P9gGpHLvsOzuPsm7etcIad/mgXY+MhWFP20MzZAPqZwAOYvpZ
n1fR0gK4pGLJzkOIQUA+w7ZzQ0RpEJnFjgRHQqQBGTJR+PbFjZ7562cGt/sVxCgWeY5X6aryno4J
Ll7XelDrN6NSjNXJaNbbrkge+KJomg2oPA8sob9n2J4l5hnzusyaAFQRkUqv5WsZh1/wBBsp3WJ8
INjZIMDYL6l5CgFdR4/grEX4XTFRWeWHacBIC4jgwt6STP2mxfFB9etl0APJPE7J0GzBRqzlgbv7
GQzzRt/mlYfK0fc6abf0HFurlwkJgZdPjVGJR5H+SM0Wig3ouWnxvgX9lycs5lh8SoU99GhcRTEx
lCBBFQPMqVf8R9py5NNck1+kI5ekefhA/2wevVzn8GjyLis6WA1oMw+gIRldzJ1jOyN2rg8gcBsu
OrI765k2kuKShRZofg8xdI1a9gfyXw4F/LnmEAs3Vk0QNwZ5Zhvd6A53mz1ZKv3uuhMWa9JerRYm
c9yBzURaYzUICa1A3iLnpGcST00Yr0cPl4dfjB2l1OHkrIGF1RGG85G3kOoOL75pRVwX2Z8qfNBP
GdonMiqlT48t4FKshxC273FKwupkQRubMve4Bvm6mobc8gpdUtiotRJBi+uXaxvID8APNBD3cmiJ
SVtIjRMi7iV67dlf7B5PRbZaubF+b5Ly6SrMg/y1W8K1M02GQkkrC5I9knnDmyj8o1VvgQF92Jtw
u/fq9tFOUurmlTV1TldRW0T3uuNDfLM5T13U58lTl3OP0KCAOVA6Gre+GHY6xsgSTLV5E1ZqMj5y
hXKc7Lm5oPCLdBv8pPH2C73FVM/biPln8Hf08RpCWddVeQ2c++vWDpYD2sY6RrQ8MeeshYEBMIle
CeaKjErgMzD0T7G1TMIC0ts5uKaIDCPgXO6lsgXljwfd3HcpSiLmmJ5j0nsX+KNj6cpgJSaGAjFW
qQN85NO15iRoyoBu/GSbWI+vsiyhZ3H72Q5bohmRdrjlZPT7x2fHl0UvdVp6pE3Sn+IefxEkrC+u
d87IpMmXW5PJvWQ851a3h2aJjiZFhBASraXO+0PUYTzN5oblH5qmDEjzPc0nflAc5d/zw2XYrdCq
lQ991QgDMyhFpAcRY88vJ0K7AdMeAVEqsFdH5Cv+1gXKN1lWfjQ4oujuosjKqQQTXC7HgBXYmvos
6xOKs/vAyRn1/M1D+jy4+sH4DjWgdlo3FwHi3wdVQfCk3Sjj9oii3SgUCeB8kbKir1ihgZUX2c2S
ekKp5WHmH6RpK8gGiX8WH0FHtVxl0X+x+dprvhLTvvNtrn565puo0YXwTZx+aQnlQTacgdEetSdK
cpW5wUh9jtGIN0Hc1//8wVY5lYFbjN2myTk2pqgaHwhtltW6FMxOx+Me3p77F1oM0hvNuPmYPvUj
wwvRA+cUoeVk7GFev5cyzzru8eVmAIKh63thBoupcI8LtGuaLsH4y/FqKoxcDxUCRF0nyp5PipXB
g8uomqZ2hw4H//JwtrhtH8TLg1FtG3eLyv0v7H2hJb00IOvFsai6d87CHTgZAyKmQvWIzQdqq88C
lsLbgqGSW/OHnt/EDpxdV5MQ3uQ8FdrTWqW+f2k/iEXybiRw6ZNn5XDT1df+HlU3hoV5KIfss552
LWWYlGVyQyQqvJwSx7iKW1PgcixXDSDVBNu+Qa6RcbCZ6rBhGtVVhHKcTvkRdBACKylul7MY1O1R
xrNr1098LBzxvTTubVg7bh6iVJvpG06O7BvJKG32yH8Eif3cD2WioIPdSg00KCKBGaJ74d16qnce
2PxXe5xSNJ6J7cYqNZvpn5RBWQ8ddjslNLFlu9sOukvjotzrVppkjnxM8l6r1iyiRSTAQEhwNnjz
OSLstgeDvJsDvL3eO2DYkfuSzQMOkWbgJrYsVNiCbfmVhsakAQxI7SYpo7tURKM74V+ueQARekEq
R+gVOSxlrFKQBZO15MqDneoqcYN5lNaEuLFRY16/+p3qnTX4jbtkjItKCi27aVBBD1tqsplTo3Bd
yEh95UzA40deBR7GfsUlBuc41qQdm8NGLR3qEvIM6tOhzNMJI7uNhioUNZ+frkX/kprSuObSj/0C
6Px9y9gF8GsfEmdGFGEM97CN+gZ9UX+Jv0RQVe1UkRqsQsrHnXV1A49yTozAzfYBwBROc4NdIOH7
eJdZeXOqj1WxYzUTiSIO0KcZRjgn4d39ZYvYgJIdVlFKHgsb63rlPBTtc24DFBJ4RUY2bpiWZmca
hbX3Jz7si7OJTLrpB/TVQLJDeoTORk3yqmSHB7jIpPrprHvHh843RUem8yKBtidcUfDFLkZnvXuw
GQaAHc4WeXZW+w3pxJppYqP17YEDfwHbVGK7Dn/hMNgNUpUEio4q8jRGmPTs0cacMSTloSWE6sKQ
HD6rUb7/5uRSflhQDIUNQMTZHcTeJN7p0fWfLLGQA37WwN+z1HkxqEGp3eIXZj7hNcCk1YhMSxu5
1Y1ZmZEpyG8CdSoMhGOnjiob0d9p1t1IA0kFp8zzDRBM98otfTXN346fxNiW7aJQOWIV7poupo7+
UeUVMMrErMyboLnSRNzqxpXb0gxtcME+v0r20wsBK9tkeWgsFiXuyzTwof+syhzbYGi1+BpknDtE
gn1XtwrNUuhasUaL5M1YeaUH41ousVoz7uNLB2peiCX2ZIVoc2XSdrSKXAMDR5QvIIqfLRJ8giSN
IslQYgaa/pR9TxhteSvdy4eq4RcgayIPHo+HH/iUbAsQFYz4arVE1ff1j9Sabx2eMJ0Oe0sQ9TkE
PVJAr0ctd+ObW4/R8CJNSV+jOCRiyqFjxWQYwNcYqhQMEwM3NnT6Y/Iwjdwtmk6sTWSEvvUlnHsX
URmUR4K+LOdLJWhuN22QTAysujXzkXYYkjttQl0hISbcr33D2iODkqBHHYcqQvuJtYk+MPrl11Zj
ZimxWgQ6kJ+yRbBH5d++fhXdU9u210d/w6NVlcJ06G9kM9ZHc+rsI2DDEOPQLmSlxbGfubQOo/pe
sv/TJ0JdwDr/I5V4uwUO3dVk0Yo4Epm+/so1Z9lFIzPwRhQhIZnHRPWpdQlcSfYXb2ELeuP67fdq
8ED5g0I7CFnPEtICPU0wSaKmoEQzM3Gl6F764m2SomY7QGceRJDSQNSwomq3PWM9UGQC2dhVKCZG
yq7U9mS6bX+i24SYgSvsXkW4B62wGDFPm4+kNCa9gOJG8IygvFPNvz5zQYV2vbOcxMto36hPUOkS
iVlQXff0WuZXvr0kTVT95aPfpijcUPPIMBodOoReLpnpi/m8CIgMX3rUqreF/4wjlzjcX/XBhWQp
oCra2n0rE/dm6nnGt3oW+5RXu26/CYyCHbVnBwgNYijHPqejccl8rSzQYh+NO7z2Yr7LVe6x0det
T+r/80S1Ekc064VFCor8fKL6KIQEqzHlHL3BM+YOWu0aNIkp49gUZxISuht4ZG2G25YjX6M2xmx5
pdg5vEhHTtwlHFTkYKrdii/oczel86c7SLCTEwRD8wZzbw+gdQo0I//hQPyiYVxbbhq+YXCWSYD0
7szdgmN7JppGrnc8vwikgnSQaEi9yiIvY0RSBDEUNCsgTXNYhOJSiSHa7btO8/iwzLjlLQsD4bG+
ZcR9OxCaUZD8olWjWjq4WV96CQRgS2CRqfcoyPWvKuDKgj84nYeWqHF6xAjHB33tiaa8PVNrQv6L
5QrMU06gmBQ7XIL1J3Id5kS1zwSWs8gqgzBvM5JvN5pzmo/fIlLh1GjpVEGE2seRaTrkPBO8b/Rl
Ep3FKlDEVQDC1TfsValjXAyNhiGiUh7g+KyQAIe5a0QNDii7V4Wmku34NWgof5cm7Vn18hQPmAAP
aqRT1mUaom94DR4IUbl4CeMdZ8wrJRTAxOieOCsQKXk/I/3wngXgswup/mkUvp3nhtKe5n/CwN1d
hDrRwFBCOleLm3PbG0ARqSScrOBBGLdWHaUBo3gBzAtjlAFqi4LWUl9RCXjUkeEWEcSOZPg0rnQn
De8joP/scCsqy16gV5KgZwQ33p0nZPqK78Gkyexs9V/q85qVtF5hUGbEqxjCUF73KZvy4qu0g5pu
fycwcwY5FLw8oS9FzGsF5VQeBPKqqu65U5sVhft2Rj0UIle3x6g5ZY83UVG0avMSLrYAutBGe4v/
l8R6FYiZ6/l1T87DrX0RsbxwhAk5ZxeLL/nFzVNYJenG/bSXnqjPDd0XfPYPNleyqepZIoqXfNt/
bF9aAV8Enslk6vN5m0/gmEcqOtAkKwXrePUGfR8tLEsWM5TMJcfFw0E5ud+QVw3y4p2QgceHjK6V
grpTBJgxj9JziZv9oSBHuq+RFOO1CV2M8UuT8tjvV5X5/0shPnygmMMnQl7+crXK+4DREbJ0zSj5
83I6rKdJzvFPJeBx9WwPCr1ki5hkentdrau72fsUVWRdZeAq0LOlj7fgXh4gQnjD5cZGfvZhvlyp
Motxb2UHdXKd2YvAkOkdoSoykGEgLqi2pdbdaN8UyKrE1ngnNB9ACrJQr7z5+TTsABL5sK2DE0hh
fVe5Sb1TBDdgA7BzGdjsjD1PKz1vjRlWZhAbOvYZeKBMJdlzBynB6aR5ECSd6xhNWdwPrx6ZVfgt
2Dz2+5W1YqwzEUWFzhNZurMn9LOGJG2kgSQHe7xVlXk6lYIBaG8swIJHZrT5cdtFjy5Gc6It+kor
RSLWPNjW6m/shUjoL3uHBbdvSsXnErPUN8Da4RFJM1E5KxRbYOcCDasZbzc0K/UNH56EpTFLWjly
x0VA05LyVmNHeIFRUZe5LHr2Z2Hx3/PD6Ee4RAXg+18nvHPBML48FNNVeglVZsYikNfivCfn+pNF
vQknXgtYVqOj34d3nkqPRQ6bPE0254BFhusTUGCiFQSWvaPdr5lLv2AywLEeKZXVDDw5f0NZO9ZA
DexuUgEyRsqC6D6r20sWZANUvctLrk+q6+5daP5dwOlWfFVOYH5hJL3FVABZ/DI7bVuLnAWXmp4K
Ep/SFhZ49CH6hoMeYkncn3DzqAac1wJ0wiNpU7Zvr/WHY84N73pJRcXEh4vRRHBVOdfa1P7d2E5r
Ixu/wDoxcDYAXz8Vea8A7Dq/nOeihJ7thxbhtg0/CUvoUKYLrtRE71oT9t6ed+KjQJnsZJbzCsOG
es1WHrBtpPO5XQE1OPJLxV64P7FgGZd6MfPXN+y02T92ZPR95wd8ldU8M5smsxQ1hfN4iAS31STq
uuvXhMQ+wNIr7r4R2xWkKxFR0uGRJCWpkXFn0a50BCcW6jID2C4E+GkpVdq2qyhY9jXtArFe2COc
RVHkY2e0nmvBeVDksFCckFTTtdELzo09eH3lg4SFV4ILHqHyN027lFZ54UpLunICwUbUOx8z8GYQ
FEiCJEn0jF4ucmbjDV7TEZmkwdIWUZYV/wNKto3TSvKbJbtRGurnmDPEXzn1R6lCOhw1rd+E3Tru
WLVC4rEc8FR6ZeDgHwnydVSv7S4bcMBE0iwM18Ep9f0mbIvBvfkP8K9e30SYLGupWy+04GXdRBJ/
Y/SUG9ssaWc66JMgORSTPT6a3JIKgssFOyfw2Zyh4Ohh+YRe3oD/5kOnJ8P+/ODo22KRKjnGghfK
9rlAZLVg4I/PlsWYZoty85K1OaabQch9IsuSMbSk4ji76tzyyVySZWKwBj+mvfTGDqrJlCP+lC7H
x5J8SwZKSCssrzvNjnTCXeSaVWjgUrqrrSPqSSNz2LFggFQf3B76rqylsTti3NKTY/VXsRxyj2pv
Oi1XV+UuipGqfc1CZ9EthcP4agwSN8OKFvCyeRoVWx1j+sDEp/d/hxGYN01KO99+kk5FPdLU2LfS
VqozliAPDE+gqwQwxhMWjAhg03dQNSJIc6N1fxQFP/4xjFl9ACHsHAs89toCheVzChZGyx6DFBHV
O5caVBebyjDTMTgN387++k0Z0Yu8mW3muqe+XSaEUkFq/AGUKlZTzvhSYYYiiJPd8fkoK9LN1EG6
tN9dVXb204u4i9Sl2e/vpDGQtOzM5sHTqBqTAXhj9ZuoNuUMYv1mp85rA3GV+dluIN71iT0N0wxm
j6teMjvu+3imJyldu/Bm/sqYklkHHbpx9I/1vOr5rSa3oa3qdUR1vLx9oCX1lgDuLRC/W+I4Bd0u
v6TH5mcccLVRMJZq+uikWCGtPXGdQroaFvHoewkVOM2HFoGgeZW9C20SfN9RSbsGcT6YggCMKmVv
5aEwbQr2iqMXV+hU6HBU6CKIwQGOD+QZMrojKFu335AMRRh2XGLuGi3JQfjZ17ziGqPTgtB6nHnh
ZDynn+QCq309I7O/HNdpDg7OjGBjMNaGWuET995tbcdjE2i3rtsYr4V1jWIeSG2nDktDx2ONIhsa
QDLcqUt8ezCq0wA9dDQxBkejASZ/gbdW6lJ01MmIGnyLxtuPab+PfnV2dJKtA2O0nGlOU6UFtWzo
F+DGIofxj2HkqVPnz+fjHdYnKzmMTht2c/guocMX0vAb+FDEZtbvkwxCtzQh1C6WVYRvEQOIFC92
2LV3EY4cpoO6Uy/R5kLgSfTr7fa7Rz0V+vWGrLS7xdhDlKQ6lyb5UQm2tV/jBBNJ3SiiFqkfOae0
IY8ZnVHmAgDzmbaf7CpqmAkS1pUKSdXdRMWdvFlMEI+cVsLcdGfz1ouljauzkqGIqSBOljv9n3/q
ATdAxMAG7H5plr2g/XrtspsBQmWLGSQKRfF959+Ke6kXHfzzEbzwqLkFwkoqZPku6K64MH07+UZP
iuLj1oD1u7XJshmrZRnKeT6fogMc8R27Lpy3ELJFCtgTJzHnV6N2g+uFbThrOo/PnxuNgkXEYcaI
tUE9Bsg3Sauc0+L8DjosztJJZWDWjR0SnZ6iaCTJT4HiluZQGeuc7FHKvHRuA1YxslukC9RwSh1e
FWWJPH9wtzv85NdGhULUvE18alfdoXR9DXv0T2QP3yEbZcPg/7UhzFN6X99xaCGUy6T5TgtDCdss
YuL4O4SMRnLAUA+r+kAl0OKX2rr2NSYYI/0wwP2db8EwUN6uUFi8gsm+PRB18gWAWUmS4IapN17c
wzIi8qLoqjXxgZA5+1gROjSwQN3I25PEiTGVyWaGSPcI6sIIBns36Hvm94A/HK025zbnE6gl/+dt
JrGoW8118773s5MibXpDiqqx9PN2eYEaEFKvgY7JVLw2z3C2ZffwSFStOkYDticq8Ot8mDECXMyl
/yDRVS73vx/SvvkYUUeVdcaNr6tdxpAt4kMZxkvF3PU+hODoaLv65ulYfubEM/D5IGU+GIaIqesz
NgPTV9qwM9mOHru7b1lXqz7pYOkfoWmfsippus4MR8DAEm1+zJYAYdeBLJpzaDLQrhz2Z9c1ag7Q
NLcd6P2lSD+R7eevGchEVXW2+28USzE/tgzipOyjoqVfZpDU02+R8zbvLA9+TlfRVvGjzo7z4r6R
SQXPLbMC1PTN6x705hTVE406UB7ratun+roqJVZdcbP3u1VhhdvdZ6Vnxm2jypNCF4yUO/2imfdG
S+4fmTNbMUNRM1mHw49ETCTBnIXMWz6erwQ1p4rtAx6OIPvrre+6oXoBE+2D9x3Ov7szM8iP9I4K
yKq93SnSCuA6pjW2bmiZ9kHOJz7kj18P46qFpqWcTsiyYBR6zP1yx5dnVhokmzHSLM4iCN7RLe9t
7x4q8eEuV9ebQF2zphaH8gFFKV/o5t7qpHz+1At/RAkSN/YE55BupIMTKB+1qe2kA4sl40HmeaMa
htk/aeQA7nDPA0gp/e3TPLC39SWs9UKDRT94clp1VlveIKtFyZFhSqtWFmUE118I1Po8Dtmlx/9y
4jFQJ7ZcQaPUChN8j7h1GwRotvFT/KPRQ8/clei39jB789cEGVjmsJc1bDi3u9J5hGxuoRBrOXkd
CdoFsNVrfPIy8Nw1Jjv0BO5MlBl/uJoC8mo+ut3pEoC53Rh5hUu14qKddf7ovwvg0nK+9DMU/hDu
EFrfgBFH4LQmSwym9DiAP0/s3WJgFVk9kZgdDhr4D38Y69Z1eXdfm4bJw8JEnqrUPiLyJYezHT0r
2IM7BMexJIdzEYp5PRnkKMlGXC3DUJ6bGgY/TvbFto4kNyLRWsPRVx3oEOzOS8amJqjWZR5zivoC
ZOOV4zBHemv/mFy1IIc7/GiLMbjox4sEtRKeMlwQ/lqwKNflPxdRXdGBcm2Dez0qQo0lejYRJqS2
opD3tuoqQOS1eT7DYIH3JfAE8ymh9KcpoJ5ZqCQq0LZsaK1/XkWHNh8OqyckU5LzUihoemDGOPlt
SEJMRpoWcdMZuFYA/AA5wCOdlIusgZ3l7Z9AdV2MeXqaRt0l6ZuyggCqTanSaFdcd4FVk9qPAaPB
qLVWdSCnDNiXgW6PwTs/EL69+WScsv8+41Yx2gu+4TsDY1g2vXcFP2oW+qm51YvX5NBjqfYLJ4rw
P1HUyTOogSXES7dYhWMvoWq4It3KygonmJWc502Ccr3ZqaWglwM4bj7r++J0Rrln7ydQyh2ii9pQ
k4mOWYyNcnMmgLQhu7OZU2ZvB0/r1rs2CLlk0TvwTPzKcATB2QarET5B9Gq+3VPEI+TxJp1vbaer
VY+/c6cxn8TrXmnJpW6vAxyEHVu3vYnXb8xCzTD1bJqoajb+FNySaLLozFBlSvIVS1YTIfb3w3fM
ogAgSi8nGZWzM33LJnm0KkpVeOgInsztgN7hUZcuB2WGyBfbnfhNfYcyQvLBoHcRzxf32zOnIoRi
QS1ZI0z5kbYbCJKEV1pMemcQyksPa/LQ9Gi2HoCYRgMHK6GQ8MmafqoetG1Lugagb6HDh4KKufOr
hChJLMJC5eU1iQbXIzOtaBkc60LS3Hic26nmws47oIooJPHSgj5MA/a0aYqSSCOFj5llLXbBW5Ex
aNfLfTyl1R9hFT5t5Jd1cpM3e/gojdFb5PNdC2Z4n4XpI3985zMmjvH4vxPjp6I9ljxbXm2/fxD7
KCAxcwrcJEpx5INhXrqkJJQoLYkO7jROK3OIGSEaS9UEwrK1WKuQVJigK6qbinzBKpTSGka4JMqH
BlnjsUXk/KPmPz3krR2uXDEv/kmqpTr1Rpdq+POXoqfG8Ja/GCv2m/dxSaXBR5Lya/r6w4ZXwXwD
XfoG+0SwgZrwZVj8sPwt/NHru7LjoFh0OW99RXl25dWeaBKM6rAIHSF893pNErJiengHZqGU7Lac
dglcyxv3+WEJP8seQebWdVI0eonWIH2rTL4dcAZ5r+vPV45iyRBR/OYRsBadLnxddbQAVy404fI/
tlmp3wlaK38ejI4KgavOQwIHxKMUzPmfMPr6YdgpU1fvLXQMPsRtf41IDTJ2TThQE5ggGUn+wzpy
e+AVBMI1Gl3cTC1xkHvxZd4OitxfLcwW6v7+Z48uu9ZZUYN+IPQrjjD22Sm7NnztiOmjDL5e3KFd
hAU1abI2RPF05qoQt+rb2S6VfD0vHjLDy/ynr2z3W6A3RuSJd6u26/b4SJWYXEHQe93qXF1GVgB+
3QsOiyAznAKxuX8aiZx6+THRlbqYMv9sAnCEYztNqmpsTXjsFai8HOv2NW6pLzLfTAkgKQZ1/oQL
M2R5PhfL6dRRkB3O7l+M8v6BSphevoXbwHOajG7BJjSP+aYRDDGGHrt54tUAd4OyqYm6gBSAOFG4
ELTPyAg7zo4goA5wo+mAT92exiV80y8jWtc3he4hVRWrsd8wPDPOi1XKKkA9CHKyEgQh40MFcXyN
RWewpjSMo7hFVe6meK6eQqf8XtKiswecQgg55xTWn5fRukiTFKkRJewSyC43xXPC87D+matM7Xa2
nd+nwN/0dIgVAlusIaSDqPfazxpKsXXnt+Yj1yV61GEMWG8CR+WA3EV40pnru0zADzq6BRwSTt5K
enCIoK5tsldvCLwvVhDH/iRqaAh0e4epGXE1BbyPSNgKS7m8lQM8iWlNE7DdqwFyl9GOs5PWSRcX
Ol/cTw0CzX7UachgEpm6WqOsdbQ6t3SZGd/AyN3Fa7G4RfpTWN95Tt6B0HvvTw9W8Njgq7baulGh
0FULZPGxLCjmp83dy7K2LWat57wUG/roBPBOg/VxZotpXi+g/vhosWASiTs2G5I3UqK1wyNBLfgj
1sftGcYaUwIAxny9DX8Q8dCNx8eQlMqu21372XDEd7F8hAnsTBVvoecg69GrUhwBrIe3zLVBjwgN
YEsoeQ7rbPxxRMzuW31sVDEJzRxbMghxpVJsA3rad4U5GqqQtDM7S+Z3Gn4BGNsw49fEUu/Q6uo0
H4BYDyCrzYwfRi3kfbQsETel5rC3K34BC3IuuBxuPrY00Nu4mqUJdOEERqOGYZuKrBROeLIp3yE0
vArgECWjghKQ55OgV5cwga+2WLFOxOzcEZNpdFsrlpaDY7pVOTXhzPbdEi0llgwcBhMId1y0Xb72
XgD5hotBMXTVpsdPdsMTKBgPCsg22YtC5gfm02hCkQ0EjdNWKbe8fXnG4xuTpldZqdbUcRKzRujs
GhEWQN0PtY2LmcPyB5+lUcG55hljVn3bzaESwEQLedtQKmUKnQ1aE1K89K3hFcnTm113YRNIz78q
B/F7b69g4ZZ88jrEjJQDntXdV7D8DNzJgUVuy73cc7H9KTPbAPAucxQtu+ckLd80uZlbUMHROTXU
8hRuthX3NdVcNK2ndBTYSh8KqCz/mnCyUa1r5nyjLyfF1ZQolXBNH7mc520z7CtAKzQaW+2O8QxD
XdTdXM+nEhUgPcz3zDt3UmDd8W5hqmuJokiO0ZuwPvl0VN9XCbpGiTcYBaWKn1OR4Wjlqq2+MDvS
KFtGOv/tKJ6rw6GCQWfQkMsWqJ/HXqYLY/lRSG9hi+LLGlh2anzoim7Jz+MLEC+bqPf30YdPiGPu
TvRJ2tVPRgPzHUSgM3sDZ+yX7TIC74qsGBWBV/DUUXLsY2CrU2nAKkJsyJ7vWvACxzXmYbPtBes6
Ylp5o9T7nIkAbQgX6AcVyo8XiInMB09IaL2JU6+kviuzR1dODbl2aIVD3mKKIfew5LJgS1xGXCUp
wVU3ibDeXVjfXAPCs3rnAZs54OJyw694Fs1BvFUj2yVlgRJPcQOG5q2rGxOKVEsmomt2RCXD4xZz
8QW7ZVbEdYywKhNsJQE8a3SXdgIoL/qpjgvF4DouN+GrC1xFCTRDgJIjHUFp4QGsaimlmFX5M1vI
hXeED16ZcrHUUcTIroOQRmtsgCWx9Sv2T/wO0RPG/K2KCdDlyxG8oa3leKeoGG2s9d6RKcBra1bR
6vbhp5X0RV9sDR60VbWKbNSlpbr76YX2jA4fyDjZ1tUqshpIKUHEkqDxteKF6jrFMDNT5d4rlWFl
dgsv9Hchnijqo90D2cIeOwYP80goZqRpTmHgTn749ARbz1+u/T+hlkdJrHXHXr92A5C3b+2yAPIn
2ONMeWW0f9zYMIlSbbjPNBdHXStA5AnRoBp3yuvM7caKyA9ZQwJr68nq+3/shlRhVJUF1HzYrnF6
jeMHsE8xSrKvEdrYOWAh/7B4Ee4eIORAjwghXS7d/3uMfMkXDaiRGiqWf3InJbt0ujgt0fFT10vr
y6bLdO0S105G8iAsDAmsxyic/VB8REhhC1LVyDMSF67j9GXynhMrNQtC11q7a1egKQP11vMTAk04
uxnanLsKruX21RmaqoNBnvEBiF0hXE/4X7E9v3tuft+7JmLnUTgWp+IxuM7NhrXqEZcoAiEnZ/nx
lQY7rLkNiGc+0B0YGxwA0jCqSo7z6HHBW4lL/WnV3n8GF6c7g52brO7y4bx2jO9rK7RzCmr+1d3O
IIF5eyGGWSp9PU0eShtzfwNvqw9P9IGaDZY7fXaap2FJo7QDAGkPO/atPnJMEf4rroJ537ap/4oI
MbJUQAPltrpFaJZ2AHfNsTCeV7cf4uqFEE3qSoDbsjbGqavcxCqkhErHLjld/S6kqu/H7qj4e/IT
FcCR9fAWMhOnUZqwYp7ufFo98YSdvEFhckMcsTRqBsu38o5gI/BNua+BnS+xudZuASRUPPT59yX1
Qy66P2AUQyxsN+53uPkd9ghoKU1s1/5DxY9KSBjMIUmNepTlS+7xusaF5F2miNLL7Q54kfYBuLv9
TygFE4oTIRcJ5W6vtKN0G6tVh3VZe/UUFRnqPurlYNMQ1pLhVXsfZ76koS6VoroS1O6IB+tfxLw0
vjkQMq5DaeUgncBWFg1z0PFwyFkAL59Xl5v61l+5crrCbU9abH3Zw2HMDTr4vPjnibyeDZtVd+Wr
tvvBSDrVlexkPnLqtFGtQGswM2Yb5r/XgEs0PceRonZ518+IvFAZckhVK2WIKvEFIXwprla0dMfG
0tkkOFq6WE+u+G+mldvl29o8SAhcjfRuE7svUl43o8Cuf1KkEARtCN87YevCXiN8pk5BC8G7B5cI
gGUk3MkH5+WYHrBAwvZ1bWz0X5V/+r17wLNYv5rGeffJUQ5F3I5qQl3g+Zj6PcJK8EMFVdJc7+X3
DOPSV7qCiBe4rPiwoniVKCrfSsAPrbRn8/IS8BuQGDbVjRyM7hO+eYkjHgLbPYyhIuiAXf122vOC
n1rnQc7U4ja+Y+D4jjqo3nwBJSmpwHBNDzxmNr6StOai9gK/z3qK2HiiSnLb/i4/tWg3BJ4PfM3J
mdkkOoGGTaKR0pM9gfz7jmF9TVBVdRYica33BSVNyKBTdJGD7ZrJXJGtOaOxbaS2eNXv14V63/0y
DJ1zaoL7TZu86hTh7E0NbXNnirN0BgrIdqjMGflMGb/28sFW9Qhym5Nqa4ptClYR/o4rHWF00eEA
zDno6ylLBK+TCWMaKXxLxdmsokzIv4Ak3RWDhs0ehh3AwzyfkNyPwBFBGW8KF0gkNNvl5ZLANwEC
RkjuUMnDyg/WzBfUbe20VqJhPbUVHjUmpUzVUcaq7i2oLv/5vsHdO2gxlNo4uXLLSqtAQtUGAKKW
pXiFbx6/XYtDwB2Urnz9NTY8VdYkimu+wIDPFpmjv5EZ5OXYOAITv0vUHjCnAGMCIz5ujczmOy5f
GzK8ChvKNwdYG/H06eMxNqr6yz7R24I1K68eESXJdlq9pwnJctIyn9AfD2787k8GsKkhjZTa7vol
NNtS6FVLpC2dX7mo412vL/ebABaPpFXsEZibEZYtTtz5nNAExW6pnhG8SGzt0bkGlqy6lg1q5XoY
LGD/62GLb9w3V2EnmeGJTc2TOeFf1Gsd4Gpm8iwv3NaomdHflrDw6XrpqejmZHWtDHD7Nkg5TMVZ
YZqQUmh2CoKPzASScYLpBNKQjXifLqNSMoX5+7OlKOd+RwdPtGW867qc1AziLn2dt4O90KuJEIxG
X4vWBrsPtHZXlqo7wjJ7I53oCmJmTcg78n1UlVyKlRYSyFISm9WL6OWX1Utq8OLzkGNuedNGc8TZ
gIuXwTf7A43uPQ+HBAUn4pLDXmWzjO83qsczi4/F0g0du0dP0MO7YUgxV3/xO4EZC4qVLhT4gq4+
5Ob98oB7IMTovNSm0+GrIEsVdbCiGZTw3/8zjPmW4F9o2/qZNqiAegFy3oXRY1ungY/dwnlKPYgb
GPpxssbq3YtlYCS3hhivowWbVTHtybl08corjAmJZxDPFVyE+CGXTbJGsUkMamk9yobC+LzGyhu0
y5CQTzLtKHei+yohEMxoyoDnqLx3YWkyXfgjd/6XBubHxyJ4oS1i8p1r8ANPyUPyYQFjhqf5orPd
gjIqGhgICEN0dK1L2Ligxbhen/dMrjxV5ghs0FOZ9ekvANttZj612j+L1KTJ/1RP6JpjnCojQG+x
K6FUompsHNpkS/GcXg/MVFBgDYIgSiTqTQVAPhbbQmQ7WCDe9jkb8wJaWtlo6q247Ebmmbns9jfm
dG+dH5Ji2Nrld1Wvtk7Z/rxjC8u18Fe+1eOENYJ1PS3FLTRpTN7DKUECc5a2o4BDcwaWEmN7zw41
JBHdLxgYoavmIpE1vsv3jWSnL45XhP7M8XFIyPFWS0MbYl4LsZcXgjuWk1N5kAQdeo5RWCOqblcV
sbWaLJy9KQAEQxTGbyW8ELFWOailEi2HrulczShKDMq2nqGMyidQTmzyOwO+pLKnUjg77TFk3hbW
mhpizQsHtnXH8xlqNM5rCtl+ymvDmpybPNUVQiDJ+F+gira4cDtM4bYtuyHab4/NCsKYNjU2h6Rd
W59EwXsdWHDyNbHnVCRuPmn60X+Ytzu+1LS3MJnMnQNuB2pkUdNpFPQhGF568Omb6LBuj2VxEdxC
gFm85EA9PWBUSWtnML2cEOpiBDIZT2Ucoa7zaIbOBJdYy14kSKs409+75Cf37BRD1+fLhhamnRfT
9cFKmLmgO4YL/wFN2Y8U9Hy42DS2S2d5SgnOdvP8QXIuHOg7RTJC4wGwV3giOoDQV68w6htFyLtH
5RvIj9zEJ6rKciwatpFzM74Bn2mqk2/ukr76ZdtjowTAfLoT8TQpF/yfHp+oPuCAz9XS4UonYAP9
Kds+RKTa67de3LmYqKuQUPhNf5VM7OBcoRDif/YQ5KO0FJjKJJKNqHI1FZojnJ80BbT5p06SNlLv
LkPTWB+nDefyrb1650+NiiPRHbV2ao2X/PPyCpgZLSaMKAafEC1xhTSZ7lvtLV9Crjy08rJ3o+St
jKE4+ImWK+ZeTudwNS/8rDbQUsctrF13LA5btGeFSYrjSRY8Ey6BMYpllzt6pFPb4kLPNQxakFmy
q4ThSLkBOuFE6MpkhgcqbBysx2TW7zMTaDhA8ERQgChjomuhf65hZtPkRt4fPx1LT172Oni61N9L
Qguy8StRPmjBRWNNcvggbZNaRZLTewWpyZuzqf3p1wU14PahB/fk/Rvn+3F1yQv52cjyEC3gL+zu
U4eY/bdqeJJ/DUaH08qm1EsTN4Lu1xnNzJxEaFkGQVfoB+YpO8msHpi3Y+joH2bjgeQi1Mghg7tE
urjnkHQUGOESFu8s+SPd4D6cyyxqHclzeJ8YF05Zz2/+qg3BwAVs8MUnhgl7pbFQVemavvzDbMgS
yykVJuPbz97jxyLVHgK5ZdeMT8joNU9EtdTCWMGzdKPlfUgZ+C/BSADAMGiz6AppG/DYum/wDfB9
rlWNijcV8MU6kYZGLa0bBzEjRDH1cWH14w3EB3PmSsQ4a2ZFyDlZdUDr5ftaPCz84UvHUwKAk9Kt
goobTMf3/IHmhKY9nIUcTVjsM5j1nn7BQf7MKIJWXDf9W39qBks8viYFUw/kPALproGV7mmtPPjw
yPyX/lL2BUO8l3oY0VjBzxvLXEVr9Rm6XGf1NgMiX+FKMtkbOjCg0SecMWjDAHsBLqx5olqMDlAC
K/tJXCtucewde1dfZVa2G4BmyROsrs2uunz5Von1Cj1u8WL3WsrhAnW3pnF4Fid3w4+T+zHXTY4Z
b78F/ecTRNd5U0aj4FbItDVbO6wl0MI/CNscfO0yCTSUGHLt/HR6NH8PhRBd8eboic6hd9YqNQn9
g3eBEjrN3+eDHAXn+4mYmTNLQmP40HAfWb9mHipyR4eF29AeCxpJt8epJCYsyt7Cu7uQ0/Hbu8SA
dxI5Kq0X7DMMRSwGyBrqawZhNON9eiZnjci5mVy4g6o5YGBrDzqGYuKI3OlTyNMuBehJlPIla+Eu
OFp7jQKiFU2IYuVwb2mFwXuyOkJtH8/4LuS7gvk4MTVOOBWNz7cSSbibtBKfdYoHOnrW7z1GqKNB
NCS9tqdfJGnb9Edf9M+mUiAwODcjiJt9YOzZgOkWaihdKfoHzpMz0lfURBx0/WzRuXNlq5CrQ1oB
2h3cEQ7vp3zPsT4s3e+MNSwBboFbKwytWEwdWPYhTcKKN2pOkBUGM0wsDSrsR8e0rtAEK2mp9uSZ
YxQnYM4L9uOFaK3YsERQ9jkjR6hixczWV6/62DtCeqOSKgSloZSCieKHnfzMwSdg9zuekvFO8gZg
+AzjUQl2rRLoQYYPErNBlC/oAT61vpP+WN3iZZjkJwvF/3swb+CczDZNm/hcnwPWSxH+NEpvoJna
vXekJOSaLrd4hkKVAY2GEk3yUVsufPHsBTlGAlb04x5lb/8Hiy7S1ygifu6ErbL+AW/aGbp9+FOw
MD8bXh3RNhXQpUrapExkKF0/OD83c/wuczERHpTly0vZIrBUggh5/MkL7wN/uyttjtHSdi5v1HMM
k0QhLcVC8Cl/Fyq2/oOZpIg71GS2nWrgXEIK6PL4+FV8Qp6l+PCDDqCERqw2OdbBQR1dMHqXAve6
J8kZljwsn+ek+8THeB+eRFmrr96wvt/JqfzPb8yzgfV3dChFSwvX7va1SCyLDOo1tHlWAPFzMd1p
D0gxf3BV2F19IB8gJDKO/aBs6DmQMVoC94J9d/TBDzIo951+blyvnYA+tRaZAzgr9Vk4cFJhajhp
cGcFlT/quGZRIvv/PaI7tjFcdY28eYhd19l+FEb+E5oe6qrf98EbXeXwzJz7Gui9dXy6tInbP4Q7
pisXG4h5YIXzLb9i5gv48S6++6VUmEu+5ogAEpUr19G9EkB7qo5bC4/ndi22AIDBkeYXF9ygD1kN
SOAjlAheU3V6yVULM9P80RbZ0RrntDzxWa4FW0rwhU6fRxUe/6aP2nnTsG6Xko4ZtPUOEYocwbIP
jgM8fXZJA86QYtrm7StUxuYshYeSJ0B8DzPd4FJr26S2PyEZKelgf52zl3FbjMqdHMvjm/Ltsms0
ISEgwS20JdutcffbD+z/DZ+URDe5AgOaR9K4k95IhClKtRvYV/60pg/LaF5FAp0HNzyJ6hHOHoWJ
Jdn7res2QaEHKG/wR3dSSO9Xc2fxxkqY4bTvC9SMCs6Z0RU+RtRvMSeC5j48sgf/ARqWdNvdq0Zg
xkmWbUBDk+mnMNjLfVyeDGFuxOeURaYhhHRpLFi6d/Mlx3+I50RvtQZ2WdJY6nxL5mIMPXC+Ryni
clAJ3rcDVAVaeNWe2QfWHIBbKJaPgQWx1PnjvtdkTCpfmMnfOrT/8z6A5rjTv+piaoRwiCTa91IC
vrloz+SW545BpnJdpgSAt0TSblidX7M0lvtyNl7hzUq6UcpMUAt/Q0zYmKFUo42mjRPdc0bZTSAQ
f0CCSe4uHbNDwr28nrWArMgdAYW07GNXm708yyovYe5ozl9Oza5HNFfGwXq6Jm0aQ86sbPAdeWkn
clP3BdCNi4+fZZiJWcTVOnK/o/Ovo5tyLeYjuAODkZvaPfVsur61lKg+h11rz0U9hHqVFGmGDZ+D
lUkHe/KPNxwAsopVS8RfrlJsnMNUfwPHe2tCZ2CNkkngdNl1xzBwOfIWLq6ySACOaOG9D+O61yBC
1zhvlq2hawsisdQeEI87MYQOMSvkFIZz9GQvrt0fFB1c849/WKOkv3DpLQn0lzbSTPri8Lq4JOqR
57x8yYE9OT1Dqo6JrKJK2m+bnQH7Ze6N1EEKQlCSA+81RiaaBa9aBvjRW2HeaAAFIBKbOSRTnJhL
XKTLnCExivu2jr7nuDK/nhnA1ChA0tlSGsYmUV6urm2qivy68gaFfTiX264jt2EHlv7voEiNgMUN
boMC81Fvssc/mtKNEnC6IByaUGKyA18abb+yrYZd/f9oa2Ma4CoOi4SIKGdB2IOMJLC0LJDrPnQu
gfzFmd3lJVcHKZmWhbZJ5q8ZBvLUaVBRzZPWu7rGOmwbydluXJ2Xl8PwFBU6m2F7kLffwK9Oeun/
ozVxpTgOOw3CpzuQAyexBBmhmsjMlAA92a8m5C+99QQqMOjU/QGxSXKdH5/gXmwGr17cGmXy8PNP
fNoRx3PYFMucmPDSOiX1UV5dak8ivj9g6UA5qJ+vNJ5tBCftyd2pvxhQpIyGthD6IY0kn/LM0vqX
apm2xphr2+DPEofiYTP2tN2smU5XNzMt8ct8O4S8gEI+BytjxOclKxuTenYzYC8mdYz8kcYoqhaZ
0b9YTV8u8N3suVJt/5B3bSLy2mX9b2e01O9ojSIyc3MK7dr78Go9dizIeDIXbmf7Vj1Ja1GRhL59
HFf4OUQ4cmj664rCXZpLZNrsKT4jybwbses8PXuiykUG3W4T0PU+xmVKLu3eQMbsl/DHd4mA+YzI
8Apdf7P8DyWl2y4tfrIsNlP1yKE0ezQr9kqGp1o7E+GlOHGLqCaIzSfMiSazKu1ZS53jmu+jmwAK
TFInCEzR/qUvU/ZTO+ZPAEy//MKYMzQPzuLZcHIcUE7adCjV8if92rysvTmd2GyIlkH8CkTV0S3C
FHF1qyMeno7FGHAawNfb/GscGy36HJBnopMGnnwg4RuYRgxhNEyIimwX7rGKstGnCZ+pjNwL7tgY
wkS0ANdCAFtTeSEfKnvrVC3qWyZs1xkl/FTceXWA8CF6dZFUHyJKeV6FYABHvmoLM3REilSbh7ea
KrTGDjKJ6A+ezsrvyLEHbbmwvUGRb+T67Xp4osl045amjzQzhOBcqCWZYvYLu6qmZyf0cxED5t5l
RJrLhAPUctkaOm5n0Jb2j67mr17n1j93/SWL/vyTIFoet1kVN9E7q1tqSSWjVrAl7ngF3UsbT9ev
tgUmo4dyMRvrhUoqSbUHJQNh3lqsVlD8O0MFottAjQtVdyaLwixQX7RgH5RdNDectH6V0aiX9/YA
y6b7FQU1h8lDF2w6lTTT5ie4KIzYKcG/O1Dybw1Rblsr0nY0hb+00enV0Uurw7StLBzojdp6zcrY
bF4JsEtP9qlNrBiN5r+pIKm6tJsxVRfzzSRVM8vt4UaoQFS+Anpcg3XKBx6M2L4/nch0/a077fZN
OS3Q0UFrA7Mfdmho03chfd2PhxyHSc4ndNhe3AYsfY2ZDxMcFuaJq5l37+utuHxDhwfVJOFBpaZO
/j5tLydqDUpiA6T3NWVX+n9Q7Gp8TX8OI/ua+Cn/HoKIqpMVh5W6baRHv7n/CqZogqboAPodsHPt
Af2AqFStwkCHaFJX3Vy8lHWHXKZYB9Y9ilw+vLRZO9Qjf2xv+y0fp4SfPjoVEzNLjIoKcft42b18
gpFuneDLPgiEbQIIF4JSDEnt1qCmv3NjByYQS2uBrV7EnzLjHjhwNo/Ye/7PydgKIpk9FHyCPXlN
TeNysCVwYn7pVZYx//VxLwP/11EO7Ur2hZd7l3nMRbUbFCjhJO2Ck5xbnZIwi7gWpiGQhPBJPaKU
VlY69SLcfSCCCAUVnGjywOAAf+i8uNQGvx2FUV1e4zWzFlFkZHCvi8sWEjIBlOVzXBFg//ZbnV0E
x3EeAaKhEe9ptw8QzCRRbYDED5kRy5qpW/B+N8n5XBwNrmK/Bb41yepAYfznyF3Kyx8q63C2GJmM
JsGhUucWrkMDeXacQaC+ikWgWePCDcWSaEVJDAWQKk6SvhKD+TciYBosAfWBrOqS66Gl9ZGaAuBO
nf8Ws52doe40rDeRoHqyM4cNF3RJwX2CQM+ggabAkOmQxwZlWCw2eTrConpCxcULIYI/k7+/q2e7
l4b6lHkKBTITWuli5pT3yIVcVKCmEbFoIM6vu0b3E5O/5+GWdrj5tlkHQGCGvJQWOkRtj6sEO2wS
rrmeGjMMWXub3r+051gEj+Hg24KiFFF9K+c+ZUcDou6NxDzctvUd7gTUfxKGisMbsmFbMZh23yDu
H0oVscwq2RNDptoTLmB2ufavZwm3Jhf/CtV+aaLkgiKLbcsv1xxRpQt6G8jGRiJUIzo5vvRlVXlQ
IFLv+MowuL0uT9HHbohw9ep8YAfd0zdL4xQ84BV/MnN+PlVRGefT7dkiRSepTjRFh9yVXYiedXLH
W43Fz0h/0LumHsxJzr8EiOen50taCOvFm5tuLkOo1qmnEH03RfC8zLTPQ/3YHgarDz3wxw1UMgyL
HOAdDbheblWkV+sFmb6MXaUoriYgIs85eUPQ4+qcEIaHfhIa+070WZfvWTrkQLNwtOd7He6/VK/s
1hK7QTHjk79lhrjiap9xCWwr8sQYzdT+0SWkSuX3RsFikslD+Y4Wy8hZquykOf7Ns+wxXBNBQz6v
00aur3MPnExhzieKpv6F1+j+j8Bvl2RsFBKWRvQHoDIbR0fQj3b/tIBYZNYybkHME8KGFkXtJ6rM
mwnBNzIR06YIF78+k8LSF8TKbxPt82NMnvXOBLejNMk4nMvbLhVQMbaP0KIaKbNi2REBkdKFYpZe
GNi7RsEL+/hqPmB6T5046fV3pT7ydr5XqOJxeIL/ThrW1hVDUQVSqRqvmQu7hXR39ezooTGBvfpX
XKzVmPY1EZRoKFTUwh5uXvrl2iYDSJshnMDnJMt4RehEerLgj3/HIcXY5lg9OvJ9MVtzPFFFFgaD
EUT4OgcKhSOfnzw9JbgV+ZN8NZAuVa4SvKdylOWh5WTjSWiedGyZpcDimwL8Pn6Vk8iS84l+sg3H
W/zr6r1NVj9gH4aZX9tfDt82nUQKHNELpvOXEDv2hPvGuxu4VGavjW70YuYNOUXA0T7jBfEmgIvK
qurBT4wzgOSICAgF9uNKSD7Z63UbTdmlDrtQeXHO8eDYVjnDwzKUw63bgGzrIqxubde9tTXQg96m
fz/LAUtAysGXUWbENJj+E1Yk8gsnx4oGQlbFL+WdXMU6w4QI38FDamgodegPXjTyRkABcBiIBtIN
mQGOTmDoHOgFotuBU+djMdwcyulG2h815T21qIKJuhTcKTrW3gSSYtVoxsCGABhheeQ1vnXM0Fal
kHCWnkZjOzjTvmuIbct+gk4+sVJXFBCK9ja1NMlxGMhbTeqk+Z5pPaUn+lTnZZRgXiV4MTcBEjI6
WEEd45uVepvx4+k29MPJmzVQJYBo85lURsUvcByvymWET0+LXL6B4oZQRpA/x6Mry/yr9ZwwPD4r
6HiuoEAKdeGtF15CTlKBWYNy6XY7ymZZ1EWLLHXaFTQQ1TidRZq2HQGMMyi2/n/E5Uq4UwLK2Gyz
rcAXTKdvzAWf30jz9cITms0Wn2fvQ84uRkxzOCjjZLqLGMVMG5BXug5LrEcOB9M5qzRt6WvQQ9XD
JKlpi8Mjm/Y32xkSP/4q5d5iKoraWlzZ3xKnTaJBcxsbTgpPr2IaAzCOVf/ZBVGzNcPb9COxOFLa
Lx91eCmDnZACEbDvYQkUSvVX+iQIyQNkvEkRvR+xc6TUVOKr82x94LXW591OfngCu1lY+8DwFsRa
pHFOHiXypkZdjSigJ0jOGFO44wi2udgKT8qGtbTCKyyH/Qt/QsR21BS0glebx5au9UwsQHrUUq40
PAniEpLmUchkFBqSz1N6y35NOlbfrAc7CdeV49As10Lg9b0LvcCW94ipOiqzAx8yHFKZCedfkVPO
xLxSSuE1YY8u2dp63yxAJMHEmczibsBusgWUvinQ9fAQ24Lrnjc81VBjiSRDP395TBo7qPtxnnql
wRtPCbS5/o02+OP1ypoBmuSg2dx9NDLEOX6P7rlpourl3FeCjREzf9kaUzSE8MAP7W3SzkkXviIr
v5dBGBv/w/VhwaJrVlSMn9OTQ69lcxRZzuOPoErx8ZZtlj7z6UEjOAYYDHQBgt2y7eAIcfuYBPKN
9V9Cw+E06/MPQ4wLkyOUesDUGQzqjtcb081QUFE1finNdoCcASX6JWc9EKDzRf42OPPyHILgh7Al
m1qLk8DgljaBy+qtK/Z7aBT/MuUp/ccnfW1xm6Qc43El22mgIXKmP04lng+Yaf3+iUATbGVCXQex
KdJ2nl/kj/gee1JCFwu/fetk460gb3lXtgizdY25Wj+d2szny0YTbYXrlQKsww2UZ8nUGSlPkSGR
25eblqqFfwWqNFLvFlAhbNOR+xHGVuZKeatGaubcI26E+0/GOG0bI6A+QsFVWQvQIfUocUzbB0th
9BIr/QQbRbKODIc9uJUqwmtMFhgi+tjf9LnZfRLUxa9MDJcdAUCcB7gJzgddVxcx1rdbbJrxg8Pf
GNAc0h0OeI7sgV8wkBHCutCagrNM/6Cxy4VCLfBRXdxjxf61GpRT9YVmorEjiySxd3BGxbx4WQuz
Y128Yf242weXe49SWbEd2AvpQfZaK/96KyRd6lzB+90kfWFiZFCNWbZ+EF4OBz45eFktb+zdt6P5
mBqjiLxyT6TCOykKj18W1Ji+FDCM20A+90JkSXzmBkAm47TMJtzF/QnWaJPM8n8p4aYKUBbhhZdt
7HvF15/uorlIFHCc9Ll3j+xC/E0sECoBtO7+E7EcVV+GvXXG5kwQB7jmdLfYOC+v+Yv7S3Src1ww
iMOKDBRYl8/gsP+K4LkQ4Hy/pLPpD2+UagVJqpyxaRIsL3fKSVdj6PgUCCur9k2A6aCSgrmxwFxw
Jfd33b0MdKp0R/sTbeBn7ImoOaWaG4cahR5rWvoAW4TWLwac1COOkmIM7Zg4O+y++2cQ/ClgoTvS
XZWxji5ebN9Qa/ODE/DI+P2gbpeh45AKlOdFkzxn/kqN8ltF+fjHoO5K0ARFZzW5dPVUZGcKGS7T
Gkz7GMOWzWsLvqiBEz2S36uEV0udz2NPqgWQjWnC5O7Wl+8Y/kInd2z6LnB0UbLsns/xJ5S82OGD
7Jm1SzINseesxxY4pmkQPADp8eBlLyf6cXq1qMOAGV67rkQ7gtlK3+SBvSkIogdcK6CkHwqh1bki
tWU1HLPZkoYk8ezij2neU8cH0BHxCR9OFxxY8Rkvny1SL2a7Ny34INZKaXSmK4sVfzW0sgqxXMA4
4MGqYYdiVeIXPNjgPgypGcvchSx2wMdEsUCZXKvVBRx25D/ToIEH27ovwLE58GlzLgx3n8mlZ7V7
L+jtEUuXUWDSa3ogSAvqYGzi7BNCTe2oztgOTqCCfknw9kQqakfBzljRilo29cj9jw65MquT02Lj
u5f+EM0DhF2I+8Nv83c5nioZ6sR9E7Wn4ZoX+Obpgz6u5d7ZhPOqWV4rE/aeDBmC0yVJ7ky8d8WS
zgm/HS+Vy1m4FlKPdL4woUKDDjhiKfGyqEIlBwQLy2S3/w3fxKiySlPp1jsLtYAb+mDHUK3N+XEb
K8nP7xy1N7GIUVZr47vgylY2Jl2+KBQ46ZLU7RtiS9psWIxtdAVw8EA9fO8USLM6NuQQfO1HQSVa
KGyzAF2R6xq0aJLiyTSZ8L/iNpCBz4fdkypdMZl+WTJmU6/EPJoAw1tqa6ukt96LILYcXSPAEopt
3olMcPqTura5Bt8xoC0g83xTs9yWAJUoMu1r/eliQWkMomGdRIdRk5JKUKl3DZ7Lv1pLYVzgJA6r
8z83Z5x4rE/28+mDTHrw3H+T++iPxYmmFGe6L/+2ELjFRBuC4Jca0oJPHiCH/x8SYFLHLLL9eW3l
bzVEjMfJ64rcROcjcVIoRZEEUyzo44oFTT3Owgv/g4PrBRrHvgqbRld8MpYTrIWRcqPr+qJ5STGR
PFfwx1t0nnf0giUBrWIF7oUE16Pr7iwQ9cekKnwoXRXi/ERla36G+Ak5lsT818WLTWujEX5t2Yig
DIrKJpuaGKyn1M22cOB1WxIfKkK+zHG40+Q9QtdUcSfp0sGbpJc2sXJBCr6QfLQV+ZCZ+x0f1sQJ
8KKB2oyD8/qadksgo8HqoIWsdRyhmc1Ppv475DX5uFHqANypc83enN9dg7pUHFWs/BfmAJneNINE
hme+avXppgrBENwRo7lN5Hox/xD+3aV0i+SLWdshJbNyBO07eDLcmH/EvRsfgiFPhDgrcu4WUMsF
i0ToTdgxMS36BlvxBlnUfLevErCxyODSxmRsRfV3Lwq18GnfkJsTniiJZXjVhLVu0zxIcFAwZB6c
CbNrM2LTDWQsa+r+zlo3P8sUMd/t95yYSO/p0D3CAion4oPHTnsf9VlwkV9j46jGCRVqQk4BotgB
ysU/DwNXu52AtIV3pOxwvnvBZ3o9/aVU6h/fsi8oxkB8LH9d5CRqBGVI7msViiDVg9i0VAo8ydev
0GmK2eUCzmylcWKE7dDQF18fvAIVRFmCpDlUuaeXBODdOMDmwZr8gyxwyIUXLIzfIyZYiWbmxoH/
vdmWzPi/QBNNNEwPEIcrnR30UnKg6u6QtFoScUHsZXYQDq4FgZx4xk8b2MuzAIz5FuRxdMF0XHyv
QPdeZtFBBWMzTknDgUqWikDBPYsE9QhKDczWoUDUrBLWk/ZUkiOGQndPF5qF2DfFmBPA6gMl8+Av
Hip8WV6eYxMCpZtMLV5b5tEbX/Kaw8MQYxZHpGZx1QhFKsd2a/KFG+OaOZQesc/o0mJrS3LGKoKR
LlOEFuioVb0DI/nTTv6LVmE3iilm1FuljLKgHo0EG5nhhA3OazIuogIn+/Y07jWBISTaKNQ6d3eQ
+8G3tnxuk9MXxkafFRn3VbjI0UfLp4gjydt467t5KKRH1fqc11CQYSDK9+K3OHsVkEiek41lVWhq
ubxT/AtlOTJn+roNKlf8kS+5eBsYXaswtRuTYwxOV23RGqunYe9M6geyrJUIHpoFpF4eNgClq+yo
JJw5Wle8O8jErCnXwIa37ZNF07v1xUBr8k0a1A+8EB9Y/erb91WTWBgQRztQzDRnZw/GGZJAiOzV
K4KJTf7zrtzeNwimvoZTRcsxJfetQMetJ42cruHX0ZWkC7xlaoeebvqbT/pE3N0N9lhCZl+mtTRG
0fo0MjmHVfZXR3kKoNzZS+JCGdWDdN6rYU69l/ZyIfaEnd6mwhIQhPoTz4liPMH1NusaoM2g4jwq
g8bhgJXb+oTHDuPjLPQp0RuG7LQ+8ieLFMg5ogLE55g1wuQmEu+dPij7l4/4oeiTbsoCFu14t1p7
f9h7qRIagKGSYhv441IHCqPylxYVEvhnMQViff007AnxZc4HB2wOeCJ53i4/zU56+VjlN+N2C0pw
1/ABjK+asDhusvc/Pd7GRdSdCUxrdOFERvugGETur7KVvPFS4JYb6hq4kQuM8SfWOPmb6wb3DIL7
G38DsOldj95vX/6SgX7xMGrZkVjDuvuS+ZTQ+J7ZTCXQq+hnHA/wZI3vygfZWna+DF8k5u96S12W
o+JR/Y5IHzHggO2rrjIJtAVo43Ue19/Wjw5gvsKPW8xTj2Zn2e2rruUo0iEuBfw4rSgqoZdBK6PI
D9nxD9PFZ0YgZi04mFu3gf9pBlw6ICkwXU/CXU1TInJis0dJHhz8+SeTk4ycbMFcnCuN0u/p5KVl
7Vx7uQwgR+lBx+07BqXW2bdOBl2z7/eWj9jjCY1obkgQ2jMYtMw//BMlt85l0VZnyF27CI+wxRNX
aEx6Xo8x/XvlqSBVS8tMZ5+FGnOVV1iiKZL6TEI62fSfWBD08ajeCl2TF4uMkxKVYGfWzfdFCqu2
cLPwuujNBIIlzmdzxGH0XYyXTepJM+5UkwT6PU0ybLABRUP9GpFaJX6raP+VwIMuJlqHuYTtdb6k
WdKTWz9UYfPKjNDP+suk8wcipJ6LLHvs6+wVAWIc82boBB2aHfPT2jzhNe2sZb+MIBzyyJ0i4giB
7mkfF+cmUqB/0LlmQQEqavpyqp+V6u+2FO1hIQhZ+P4mFwmJFQqSzGCwKTFaND/MJJmN3oN0ttha
siPVNHWZY9kF/XL3du+vL1dTlUfK93TJdc7CVdiJYcETLrLOVTu1qd731kAClxAnnk6AObFblveJ
/8ADv0vFzxEExPomI/B1Pgh+Vc9ea4dDt4Lul044dUlIRIFd8vprOWYt2OXv3fleGKE4xHNYODUo
MFlJX81auV4KS8U/vUQY94gkDAhGv4P4Hj0IwA7tJyOi1q+mvgUg5EtM1AIwehrPAtCUrXEqM6MD
+lav8IFot3rKyHeQfCenKZK7NklhQeemg4X6+FxRmn9+/1QOB3OHL+jhnKzf1os94PxCwoki/gqd
bgj/HUKP7R8xOP921B8JmldHl6lNn2Rxordr1OfJHcAm+clXSYPdYp08MLsadIpq9bB6Z7SORtb9
5zJtmUa4V2BuabaRFlyK1xM4+McN738tkENjqF+Vv9y9e25mgiBXxi65su3MK4jg3envSUd+sGGE
Kk36s2uOK17i4Z/tC7WQaOTFXAHRZ6wD/SB9WdP54X+9Jv3coV6QI/jcAFHYmR4w2HlZM3uBvoGD
7xuEjjuINxxmPXKDnc8OP4dJfwLuCiHoGFJUfxhMijb3nKSZokuTS0wyM9I7ellY/28FtFlCzDD8
8IK+fzkVz2dO9+5HLLWrPzitVAP/V0Oe9UppTCD/9xVgBis3wVqLHyhXO1naQo4y4ROn11PCI4V2
3O0CXhMc3fXN5cJGL5BFfLfVCgKBWoFGRNq5aZg4iX5L2XuyqSZD3E5dBU6HXcVOQGaOalu7RoNG
gFab0SVqPnmjbj2HJOAOq7bF/pQ9/yONobdVRUzKJMU2qIIFxJxElQllk15N+dCSqiOxxTlCIM3r
p1IXXGxV+EUXPHPCs3BOxcr/DSjRFrRLjUVDs+TueMIavRLolukfPck2uVBXuF7XMXJgAsYtyLR/
rWbOl7PG3tMQLb0Ol6cTHlNFbDrCUULKxP8eiF64ew/wN4iUEqvG8CQPvWukmp2AeftTDN0Mhn9o
NWKDi6VE1rLAHmpOzjIlaO/3rSFSLSOVz4GxJsqD9HOr5hzje8BwFqSWz4Fi3IQftjcfDoW3JrSR
5tylyCXZixn5zu8mHKxEmD4H32G5MN8IBq4R335PqHDo9fiuJeO8dql+sRrBj77/wh3xpvhN5y1v
ak06qp68AoonrIuZ5vEDokLCo/dFcUx4ECBNeD96yqHExU1BDmzKCnTyuN/G8nK8N4l0jGaFnxDq
NVTPPsN8ye0rSgYZiSqWi76Y33ko1iZWjEuylpDk2xUTZTpHFHTdxol/1a6vnzXzFyuUUqmAHw95
mzd4/N4HYJaIKo07bosp9saXCEmbE+Ah3YK1ghy/NDQshkqrHqPbMSZDSBHeMNtXWTxvPmJtVwHn
O5oOLixqX8/29Pxme62abp/79QEAkE8YRLPJ0jKXtBn71itCVzYDDSbgWwBi9WWVB5Ul+6BxzkIz
wDuMvMToRaKG6R6jIJr9e6dh+i9RBafkaFeUp14f7EdtY1k7gyxgegaGTLqtF7/r/OCXgAebbLO5
J39RvsT/SjSZhowM658KjKXt9ZRg7+WKjzduxlB56gTsRv3j7VwRlL6Iwk7znKg/tY6XAWYvXnWW
HXd8A+ETQXz6/pv9WYYiqNVHAtp3G0UxL1aB/khJQI2wAZHUGiIjpORER/YCe5Gcs9yttuJWHzpS
MV31EbBHY+NrmK8j9ZCeHEmgUdYl+xkn2BQiaxI1X9JU6guhqPuLepqnNAtxOewXjb1S0ZZw7WHI
v8q3dS0hw486LsoQSVyxjCVLertEoyDqczsKuVqLPGjLh/znQE5fnHr/PZX2SRj/3jPNlCVOwb0Y
Wt44oSDgq8tIDh99rgnnU80xj9h5UTAu8+t8cgQ2D0d6b6syr0jQWPNv21bSQtLSJgO/LyyqFOiK
2H205sWDS4LtuXoPaTqucjOubob4jzFukjKL9Cc2zIrGxsErB0weJXvViMT9GCSUb9T9yzaRZghD
lCmk6Nt9xBq/5NGM7C7Lu+A3TXgDRWdob5CM/pBiqwpFONK+cRCg5ChcJg0iau2AuIz3b5udHr3h
tvCE2zby2k7jKoojWeBAO0rLzn5wy2eJCVyd/aaKhZSeXjXL/JYGg75hrrQ2M1MSzy/xtViPno+Q
Z13Xeo9ByLPYbMMucJW7Xa/3ZLzi/10W9RTPTPiAMdmy+j6qQnX7ue4PLKqW/fnuUXM8A+PjE+nM
og4ag3jQaDgucMeGJ+2aKUzeB8buYDXUG8GZoiSz0bL3n+neopd3/AqhBUF4l45Ch995Cz40EZV8
oyZgdkWmEQ72kT5VSm60CdreoaUyQcvJBk7oZuJMi71ha9N0HMoswNCaFESkpX9+bD3xONhHdw5N
Pcj/e2vmuXeeleYYxtVrHpfX4vxAtPsYIYZlmLUlIFerOHc+XrGz9Fkq121/l6j7a2sKjBhR5mWD
MLiMwkhGWE0aKYWmDbj9vhHgDXLOOR2xJh0uVSMh6a61uFzFIFlZvsZXeWhVHNTkyfw4blULm1q5
kk1wDt1KrTK2R6g/QZxiecAK03FEU6yg5lPTWKGZoOqEb43RJSmcIHOFGK9gmcjB+jM8tPnT8ssL
mnxlv9hNdL68FYuE3xDTSiHL++1pVAx9wVIaRwHi4MEL3whPYEImtHRzZSG+Lax/po8csIWQcDCs
vMhSqqZcf8cdithxKbetviJpxCa6PGPbqsU6Alsja3zbNTd0CKb3ObHOXnkyup1zvbS3/XHsSND2
LuMqDBO2g5U+Fs8ZJ0TE8FTdydUUoSDhQg0BbtYdS3KlHWkHLi790gaXVAqcpvW15yTbYj29dR68
OlLmMiX+pPQ5nxOoJ2e9JrDLsyeVpsH7Cc03iY1Mbet4Kltx7pGZi88PpihwtZB1bYxTWFWmFKO7
UufDH3FCzhG6bVFBZdgH6pxywkGiwhiE3Pcm1Hm/tjIRnXvNO5dVxWdX/edLPHi+cK5l56mQSTm1
0a2UvA4u6CGpHICTehkzc1PjBoBS6URP+8xQkCbpDnVrQLisuNTcDHT3O1TTI4AsOWgyC+G5Sogo
g3KV0iaIIsMR3cJR/goTYDH31XHSNpiP6Ex6lidzqD4bh7LzZbwbLsToD8kTTyxrwvLJwAeHPLF/
8XpPGhvnNiV08zxPhPamAygJIgYuDIaWDj/9VOK7xdVyWAZeF3EcHlWhGoPU3UmXVIuig2V0PHVm
r+cllLWQCj0zH75vxLW2MW0jrT3+rGtLuxWbJiZXYQsAJ3hbg7TE3PYZejmp+mYIsOpcUa0e2C2w
7X4hzQsYxbf+jHbTJhzD8DLHMsHLGnkMGx7RWHFnHJDx9x+JXozNt/tySNX30O0EFqF54CwdQDb4
0MWQfm9SHRkTm6Xn27O54SawS8BAWxxBUjpqQqjV3Uqq93G/B3YAmVJHaoxic4Wb323BNWMWCVYv
XVVxZesqH6CNZ2ByzH1USSyi3DTO1g3D2tPKFEfZbcIW9ikDk6CqRt0H+RSlQBwDNq6wqol9jmv8
IKSVc/3v7ZyXne5qu0WT+viNCh+e4CXLs42aFhlkOLMCu7AaWNxA85mZmI27ylI8f8Tq/s0Duky0
S/XLuz6VlNm/NITWntiDkFzdwsg0I70n+uF4dvlCn3F4molKoppozbFODyU+u3DBkqKJhCUEdlEI
may2LUEI24W3S0yWjFy8W0wraY370R4W1c2fkf4quIgriiJ9q8YY+eZQp94jjjs/S6Ur7J+4VGZ6
xq1zQ/BeF2yl14Oj+d6WlIOtcLbPe9xQJRJ4JeRPTNiLAkydB41JT69P4HqfCH+2hHbotEP2H5Zn
iGlqJdkAmoxQDPaEpmhLvqxZlZskx5JPg8Hv1ZIF5giz7UMgpCuFBzFZNZfxPd3iAOxUD8dvihrD
Xjx2a0ft2C6ebKmom5SkmEiRd1g4bG9epCtjIL88Nl+IIxjqEBqAiueMO0JAy8pOc2NBPGIIr6MP
IpTP2qhB8zNAsHzQLpSvh/ZitWn3mVcvRvX29FY6PvjSCzGQwwedRj4h6wwmnjVBkMpRXYJLPBSk
JRNi8rbt6cIooXx5hbt0/idYido0ye0KiSlgPZHbs6dkHUnPP34mhAP2ncbMu3uxM8B45NKmYc8G
vgkQ/wpXFwPQgocy2NECZ3zqCfs0g3/4lnRUqYW0T66p3AXxgJEFYjgSONHwhiztVw0C6gyMN14G
fkwCT52l3lwHaVGspVZW+8eB4zpQSmZl4kGHmFvkCriTnqO6kiong2BpdBT/3NtPtRlxiQkWerD/
7Rx/WhYYQmHka7grc137fLaLTzIAMG2DxSazbxTyQTnsS7VaU0BmqYy/I3a8qkHsQPMIXc/nKdy5
IqcoHw5QcybEW6YiEviaQW9DdSaQN7Zc7HY6iTQ93EJ6bor8ekrOBUTKnUZGF3KzM17dmXtqzyKT
x+cta/cJMclS7XGEy/ECmz002JdvnBXk2kKMZOzP//WVYbLO2g0OkgiOyj/1NByh+xArNKpLlTc4
1UUFijPR/KOEoN4BLM4Ooc5F0buwgfzK/cjjiZEuVi0N4/LOJMyBmarRGYyZCqTxCASi3awl+bVd
tQb4bRND09706pF/b/Q+8s5QNbNMQuWZgoYF3hGQ10Y0cKXFH38DGnY242RtVrlWl7mkBymzeDx2
63Qc2POXTgNWVo+Eg/S+1KYKPTCoNpaUaowienX6VZanlFMzUqU4Wem+JNKJw8sI/BHxAKWo5jTo
O+LmanAOnWjwJVgp0Me6csnZKn3UNSOUuiSFr/mtskuB4Ddwgxr0euWihak1o3XLDeE8nhGdUlM2
yGc75Re2Ad1J+UZXFkHxU7W6YqRn3O8ndNLMPqSq4h9Fkmqweg/G2Na3U1gBquWZQtHip45bC/xX
jcYJrjLBzCu+qbV9+06uL+revNZx0ajSwyvAaArjIC4IH6a67nAwU8TznM6dwqwISHPrqBNyKnCu
nrKJfk9w7iH/Y4aymdMyI1OPh0lqmI3zMUYur4QQPD5J0FzAunmgRJburfTeRv28uD7sLZ+ijWsQ
3aZvZJhOp1Hw7uu6a1R08WlP5IeaZT51nqSrCCS45PaPg6bMQxHwYOl03npojTKBkaA+3+dQFPYN
3S2W6oqrs8o8Mm7G029ycWXVbi888ALayuVB7bRo9HUSkqDJQ7+lI8UArSt9WFxsoqOkT5PsU2PB
rlWskW3AZC3UySapA0fMESQR2e2Dk6RzlP/k0J5ip3l5fqyuD1PLdxS3JkZov14c4iWF1Kvn/NuF
+fC6CcCiteHxRLqC7QIrl7PotxbV+21oJvkytqb1aW+U1Pb6wCJc6bZQz2+Cz08KmHg5Z7McOiFc
5fxIPfyTHQCm+sdF0+EPCctAepHPie4DOIr2dZD2nz6Pl1zby+MMo2REn//5qKcqZc2EysfqDjx2
NBKjqctb3yxLv0iVRYxxwifWZY2BL4Qa3rO/sVJueR0X7EMPpcjZuojzQ3aTUB9AImUbdP1DOila
mwl+acadWBLJnefVTys3AjNjxsUSyPpvFF/ET9r5Fw/PndcOivZvSi24AF5thR53bMkpvKcHHSuR
r3sc4KnFqHduSex2cPLAmZITx5rAR5ns9ZNZaLg1W3P4sdqrtlK+wdBO0zEpTSQknU0mJLmc69MU
VTYGur/QZLbOJAvCXE0zy3npIap4ESTkM/GwexeBa7u+HaEkHYD+sJoDeg9T3Vt7gFrVclcnmokq
hfg+0UzyCp8nF+yspq5bHxL30gN7OacNF8zXazCqClbEmJIi59XJYm19AY417EBbCys8kGClCCM2
vfZ7HRIb5wa/iSYjdZXOct6ltDzhU9qJjxTlKlgSG/mZnExgdJhps0x/qMzIJrJ7TslEr2pfE7nZ
9mnAI4WTL9C2fssKy984OvGUq6HHWB+xtI/oQmf9fO2dHtGD5303Z18hPd9t3eTZK0PtdvfobdBr
XThctVeS040qZfceHb0n81+YqVXY4DW+puOvqhq8ezf8XvEKW5oC28vtUrb8N0Tl+JcV4/SwgAdk
hSRMaeat7Rlt41JFMQq5Ee0t20+oOR88GCa11p2JbtIRuz9AhsYPgefwFYOE1zOMf937Qg/qEHoL
O5uKQTnrEBtjUM6DGAlbZ+ob4A7NHY3Pzz/etJS2AtSf6XjocrWOWyi9a8saOeSGbYT0EiIy/zam
c0K4nILquHk9VJXX4nWftb9bv0oj+Di1+i7F02Lr1wFZemRn3Iul35RkBfpN/4C7wbbnoRysG438
BNhyw1PfmdIjP3i/rpJzX9F46Lk1TFNY2O7fvgSm6QWOYcwBHcO9hEhQbDSF3h02AfnOq80LaNZ/
1DiR9xRlgPryccMxv7XBbH+2nI05WcK3K31GOKtmVKEpoSFDcKcqLuIUEwnxvrOVIxB4MwDGzWrN
B4+iLTpxRPycAmutC5W9m4krP8BtdSKKd7MxRTgjHKeVgh3bx+nksExJ/4GJQcIfyUHhkpDcxH4A
wPB9lGiNRuWxtyrnimI1uMutViFa90QQ5QkKFWpNO6acpCV2TfEo2/x2jN2+LEwBxsZAdl1d5dOl
sP6qyqoJ1jCVIyGhwsklE5aarnwkPvyRrX45KGEwUE0Y5gIYKskmpJEtd6Z4ECOlEI0h2SRYqD0t
oWaFxj6VxM0LcYxEKSD1DC7/1nblxl8jGyKUMs9Ed8tPaot7zVtFodG/hrJc3ipy4nNboxaXvnY0
QXPHfalF55lLYLWah2+RRT35XbtYzWpYhU68wj/cshQ3PJDsFbz/J2wJQSTM8z9lJwXvpzPKh6vr
uPJ1mxPCqGYN58QpJ3VHITqaCklcXb3f0Br2oam9zvuqNZNTHRYsi6Tkov26Gzsj8Voj3wAAHPma
l+apWLLxU2AsEPQS885UIXwUWnLFUauJ2cgdegHKwAbaSICdlKG2GET397JMrOrwXZZHbXBfVtpz
mfSwpZmvsYKPtlVkSO0+UdsCu+KmBdRDekN25yhE2WiT7LdJVs8Ar9hcg/LQvX6dO+OEaF/Eeuct
JVBe6gkkpzaZg9K9DxTw729hUUiGFDeSfk6guPnPrQ0WXGczSz9Wj8bXMNNEFnbxcsNylbYiKjF7
ddaFHNnwqDi2Az9gpwUB9q0PCXKm0CRXXwtjDZIxeOHBYbNHDtq7RRfJT9/4ODeDLSmMqJqNEY4p
RiLGP7kGQ/kb8pqzbt7mBOSTRpYXH7NYk5iE+z6ZunMYRWM8GGSnSBkrBsC9bYl07gmJi45dW5jG
1dDvJY5tnCUZCaj3Yi4P6eyMkILNSgYl0BfQ0yO+hHBMEKco8zBxUiBkcTfPD7ZcE5/4aFNyHj02
QoGwF8lBJPGk3lHVlCttKTWA9LQ2A6QAgTxL4ixhh+w+0Oem+seS9s+sF+8uHUaZ39ny989AxgWI
RSdloMq2jP1B+n6D/iO67pA9aKT2Qtz1Nnmlo3okYct8LCtmtDrlI+4cdH/7rL8ri0a1ogOojBl9
bm5DGEuQZPXqkaOAJkbBLaMXJoLgQiJUbBDS+/S4w0wzYSGTZ9QVYnameCMNyrFvESHUqFyFoGa1
hn+NrRhbmBtuSxOhrpZaN4YQuFju3v9NyPO7yylJKSylwf41VqaA4uV6yaZ0L1vcKpNVAZHRXnom
j5ROy7i+QPMDUuVCvDqgUcAUbJf93AtoYg/Z53d3tBIvAuQDjKRpVIeW/TiK6772KWLRf4td3vU+
/UEbdCdB5gaoR3vvrX8FM6xXd2uXjTIS75LE/V+Fu+G/G4z+uC9PZNdxS7htEOvzu3PQM6G5eue2
/TNWlActn1DEqSUy4e7qiB708mSHwk4G6D1eSD8exl16TvutRrrxLCpLeG+ouoxfWpQNx9PWf6xC
gjxPUhhYtdmVFPcVcBNnah5iSezQYq9oKtBrWnOsRFwYjl4p3Q4D+LVXLiOkTtTkP6BKpRrnc2GO
IRdAhN3bHNNw9nzOgwi5wtbWT2CEDspSVAHGpysbblYHJa9jMDdDmX3SFuiLQLByBw9DNgqThLan
goUlVhyUdBKxnuhoBDXZvqq8DWx8uGaqTpP3GydVSn96WB4+atQDWC+WdrY+4ielWOgP2qoDQr/U
ivPJ2iYl20QDOKFYbZMOmCaQ8rHLjCIjWvIx8SSkeCnoOwgW1zsBLyS4vSB6LR4a5DF4DYabwECv
uT56cQcH+tbQ+tUpK2hW6ynpagZjGULyQqB4koFznq5lpnPy/hKqUDwtteco3BWdHlyaB4qKw2bY
aGJbnMxEWvCxTyb4JrbGtLm3olZ8dx5ajnFIcfVv9gXE41gavW4pmDkae7Cwor5ms0x5GJFWQIos
vWqVP6zpOB7pLa8mH9u6WcKbAhw/2tumTy1sZ/CSmNzgHF44prBS37p/75H4+4gmNaMhNToXmQXw
NqsPLgqgRZAqzt+F8jvjvHiuZJ/yT5ThSQX0H/P78kOJyrk2LZ83UzX0OzYy8rtWgmsj3jmtuM5/
YWvx3llIS8/ciS97ykZlLwR1maBbjZkux0C7+Omt306W5NPC7q8PNYQkM3rvYO/Xgna3SuD5PkP3
TQn5W6slwBIqQoEOhe2ox3KsgmX1vn0/EPzbGwzcUMtIdEY3B8/lG/hvHJwjLKZeIFk2CUydyL4I
8scCFyioUtdxr4/RtID6u5Ao4TU5AJBMTdglbOlTVZrxRUWeO8LN8LJoopfNCHvIOvTdVXjxW4Cz
E1qxWBeXkWcMdQ4mYQ354wUMHevWfNV6iZkwbeyYlnsxip7WjH87B22A4qcqEsxfFiRVm3FDZOmI
z8+CALcFQ5MQbgebymlb8k1iiOcPcwswixJG1qnAXYxB2+f6X9AnzD920N00peEKfJAqzcNWvPdT
Wp7loszx1BhAFC9HGeCGAcb76HTZXeR0Jsnv2SVvz/JwgQq4tkXk64u361BF0bBFarX4AyHWWExh
3XdStz4T8seyAL7BTWcgGWaMrVWY44WckhPr5tZaU9ys0pf+5jYhw0t+p+DWIGWE3B6P+nTE63gA
PLTz82fTxzJyHMfvcR60msJOX8i6UgwMi/TcF+rd+GrlHvA3h0nsi+aiQvgiM9kE/w9/6qQyKXIU
cs5708SXu0urTMj8JA2NS3yktxHinhdaieNUnyNZD6qIkpW/piREF5SbFLaZ9NJeDAkWmPWyVzmH
IMIaNCstd8lNLi0ZKWEqjKOet4aNrkxkEazyT/DCGcFR/zWWaEgPgrCPyvrZBzclry/B5Sb/WDNV
82fYXTetdck+FwD62aVuxPUDd8fFSFOGRhq8omX240oDKRR5br5oZLAKZW+LlsCiKZV3awOaJFsU
eliyTMm2myHv0nNt+XPcY9t0aCdi2WpSQr83k5ke8JMAMn5snIpsGjbN2C4g/qHG9KtbE9nDqc3P
K4WhgROZ5cloXo7tGxnv8ewqjBkal/I/g1G0SB/HOwYHyUnXNOfLybS2AtoGrhSXSrMhYzc1g1ne
FGs+LwrpMDDQYecQc8wji6g5H9lRuhBm0OtRcwYxTerkQiHEmXDU7awotZ4NNNNgs9U0BR2/07YA
5uW3hG/JN92secDcMc3+Kxr5G0h0BDqTbQYv2OwHBEXuhkNd18ggHRXFmB4aq6WqGhcCe9n3+dZM
DA5uL6MHYnUL6DvfqoLCt4pzqU4oGRlL+fyWYQj438IBgXbcxL92/slVWe5TWlINKhYfsY/dQ+io
czwNwbXmBAK4W4C4HURs4kXnR+fizGIIZzRWnNXVd3pffp9p1AiG6XIYJoo4HTCnA3wbSbqPO/Yf
Zvngli80HsLvWRVgGY3km7+bGkTEM6AzlPnhKcsyKLorXyRmy40wqwOB17Y9jWCnEA7h7QqWIltB
tPhaJIRd6y+0igivgC8ioa/eklVGAb9aGYZCgsBR/7GV0g7acld8icbY51VfmGX+JEKxUhJW1H7u
fVDtRZAjKUjgADiyPk8b2eMEar8YfaPfss6pujxcb7ooNhIuTBaRkz5R7iwY0cxNp8sufSmkuI9B
cp+btAoMRCWPXoxnWgMhKTw3CXrPlMCTNylkY8f4beUE0joF1IZSXO6mX5lC42RVlhmZv1totJFb
quQiiAVKS7aQaPY8jLE7PUpLy0mnDrEqciew44L32w6wG423WWLJiEI3UaAbN+VTsTyH4yO+2oFM
oIwv4xbVgP5+LXhF3CUw6fMabUVUHT3nZpq0Hw2O1PqMGR/o1ULnhdaOf/kukqAzatXXwiRh7qeE
plv0mjbX2RbsmOJxWCPtcOhtDmKIvVBAoChnSdy71dDMwOYTdZCUVqxOkfsCMF0nm9Rxb8FWT9Pw
UQKS7d8JHXZJUlXREo85pX9mJAP1YYD+jr5GmCG4WV/BJ+UYCIjrZBtunf2h95rgamVuOLTTXBLJ
Gi7R0kFh2egsuTWOXvNoJCF56TL5J0jmJzwG5aZ8zqR16nL19LwcUN3xDLD7S7E+vj5niD+Kt40Y
SLgrEUqEUju5WOcpglxY3zJ+2qhbOT/sgbhmfRmJsliQ6b7OT9rZcBlgFs7dl6aep0LWDvktoNTb
K3Z6RgJShQp6RoszjSYzvjWPyHxyY0SpHtxw5OCXrSKelIRxgj6loORoBN0uoBzq+j8M57gz9DA+
m9RKL1UDC3V+RUekVuc43xk3oySQyht1h+6DCmVlH/+6ajzZn2IqRAUya3fHwJO/sRCZveqRlobp
6nZ/T7hDbBE+KzLLZisMtzgWyaTQSb70tTiAEkJHQ7mVphgEOoQaMAV1Mx6aL/mknXBhbXSh3P4D
ySUmJxotpaBQ+wzhw9kkLridRFsxfJu8aWmW4P+F7w4h5knH2cAcIs44pbkAisC666jpqr36rJsi
7JWVK/v45jNWrswyvPny+4A+zN/pKbR8gmRFmv1yW5e0O5MxyfrHeuy2OvrKBp+PZ2EZrupwl7vX
ff/ZREZKPTpgJie+CqU60GKbqk4br2xABhWFVUPGfxhWB+tBAtLx2pgzDTVRiRuzo8EWNkHlv/9F
Px2HaZdFkwVmQVt+6pNkgEp9hFllVx1oLbj2Wa+B4jlZDH57rZQ1zYQ6araUXTR/SjIbtn/yLnSQ
24sJ//SOxW78Kvy4NxWGI40Er+b0h4cKu6V2GxsV7nn2vhlyueJpaOV/fMcGB/iYObh4Ay5afSNd
hGYok35rr6T2fKT0NgKNPp5ykr+Z5anwDtI4TusA+BSyojoMPtwQVf0jiSbBXPV4FRIPnJTlOFjC
2vE1EorBwRIveWnSbLp9qZc2PSCbSFiXw97Ax+HWfpybQDpd6AqTBEa6pZVaS+qGwBn/YqYHg85/
r++AcZY3Haxb+AqaMP4RSeOAzzkQtvSgfwyWGHixyYk8sIF6Y0X6h8hARWNG6vvz9Dw3DAdJxTIG
yV3QJJ9WwCFojDUy1VkwVKecVJSdecYy/+z0ewDuLLnX5kb7s/hSznHZG1C+CniGw9VhOCAoSV5x
YeJ8XIqhwZBsK199IOx+evhNcq+TvsVj8edJXl60w5jV/S2n53XGYMcBE/YBt/GDflqO364nowPm
oFczGgxQfTtG/okBkRoNBuSgaxp6L5E2+o6+1VSBukH2iCeKWvBBlRbWWkdqasBc/KgaTT5hGe4u
uHbr/U0qhqeNR71kqyY5TAn+cEyXr9JLEJpp4O/M8rmw97Y81Mp/eNkYufP1F6y2qF4ToUEGI4Qh
7ST63eTDjyK0Ne/JcfwjLjjXFYiIs4lgABSCrNA9BRpgTTqQ54QM0IYeNgE8tEoFW0ui31/wWxq3
mfABIxPozo6Sp5+lp7d9rrFU9K61tYueQe5Vo1AJNp002Bgn8rOmJR6wkf3pkgLzSD6XMmEJI3ne
ZiREN8cXm2gP1dNqPeKkZ0wuq47zMnIXmXJOvlAFe3gAO2CUrJZ52kE0Vj2MGfkfGYbJfKiIgZjJ
jJXqq7kkcHSc9iMZ4iQuWEyOqfvkzUr7mKxtMpcu724sgSKyzM8ytIq4e419zP4WaP2fRXXIGdBK
rARIDGTfTihMe42S5s/QMjrVA91cKDxuTZvYWx9Sj3Is/jzJ2h07M21ZCpcZ+tqiU2VrPoKhRoBh
qQVGSepYLzj2xzzfbgxiP8QjfjxKYIFj0O2o8Ljh3bC6PGizdViapOrsgtUFWCig4x+G3HUhmfgA
2iPxs/+pn61VW/E/TbO/RFrUpn6UbaP98Us7Q5hMy4UstvyRbtbdr35fF+F4V4f9lzAJ2Aah3a/v
ynOZr2At+CqLP5xO6BzEVuuSucsk+QgsPGTaRouypv/bgGtqggKWeUftepJ/EkGsFKT9RbtEtPWF
45tnPCECaLsNiJYiQeP4a2098jX64FyJQteqNNbQ59fQNHlCnJbvaE0W42dNx3HWHUG/iXqZD+lH
BdMLwpo9zAfx72+zR/Kpf309qTt8r/UFIpbBzx5sMjWjjTe52J4TCUwMp5M0LCj7ZH/qCaGYjsuc
k2ITEuCrTr7qwbmV3aawb3oAtx6/oRZq0Yqsm2aMBViql534Qf+hODJgDUPOxCv6dDUDKac7JwgZ
+so2YPH1sySVjqeFvBqeMJ+RQ32hYOc1gZ3BMHiHQ80gBZWVx1VTAYZR/MH6O2R7QjLoMCw/rwtX
RAQXJYtWCHv8NwX8I9w/35HrjZb8QmZ2xMf0ROR9SmWqH1dnYw+Gl0V6wm37bSQ/MLlwxV21W7WF
S1WJSPDr+Zw8ugxT8e9gB6yHmgw3l/LJOq8HaNpB4A4IyS1jLiV4o0dhjNk1azgmc1JSJHc3G/HP
3Oep+8BXALiaffm5BjExrCEtTWW40fYGcW6pZDIF5n6/Hsa7se+My1yI4kGKZC4A+Uk6X2lZjDqd
1dRSnnQ37r9+PiftLmjsgB+bSmCmpbpvYLBQtQiZJYfj+kfqdOmwG/0M6uSUYfsilPlNDNLchE8O
Fx+OpiRHJ8TigbSkI7IyUS3H4HWK/TyepLzF+xrMQATJe8JZbw0duTwDnVU2exX4r0qFvCSaj2RK
oiyZNu1yuC85AviE3lF1MadauEC1NdPWczb+UPrw9JCFaiS9a5SXXAKZBTRkKxRif1OdVSlLTeX/
yD6ESD3yTwUkf73F6zmuoGG4SNpzd2wIkeMe2Cmp81FQUslF3SujMYB9ut7NKzmFa5vHWkFl994w
L9J69xo/Uvqkv5tLtOC/Z77HEhDW5XeVgYQIdlumOC+hzVnR7imFn1nFqH7vJQX3vFsPW4TE5XQg
whaMxE4HID9m6ioDRNMq9NbN65MTon7EvRzzu7HknBAIbBkq/6ozQYfgeosX4wT2KUPm5EfWl2VV
qsz4lPPpYFSM0a/EQJfROniq8hZgqGBwPc5VOfWZOawFhaSHeVfm3k14/2h6pmxLXD9cF100KQPu
NSaGOwadz81ZmnLRLFQBE0maUgHipKjhOynZaLD1YA+VWqV+iicRzGzt1dNQoQKj9/lddrXYbYMu
OK3vEl1FPuDghR4BXfgQrUsva0UrrXsqsEvFvNzDz9vin39AUeQUkSAxG4PqxyoxsLfFppZdkfJA
nHQuUVCJITBa4hVYPGHwvjnwFiT5/E+UqIMLlt9PwAx12bAB7y+nyoTvtU4bnjVPqsyN+JcUfwF5
eThlTjMeCac7+90Yrb+eRKjw0wGyJr53eQJ9qYmBKSLi+QdCmKZjryjB+BrzVQ3IU9aCwU5cyTc0
dvC9ZbBxLsHF4sc4ObV5dat+u6Gq1zDf1dIe6Sy5Us55YKweXlo3YlpBzJy7yERZGO+Qt6LY+aFE
Zj3bbajtZjqFu71Q/xxJwYCdZQp8tIb888KtgsbYAMd35uX/JCWuMprbCrUdfO5ROI6LbHOwpYNM
lH4GF1nJKOLY0GtRf0UG/piVA8K2qfkGKJDbB0hLGyZtuPPJu58RzvkdaxflKRsppb8vPZ8iDul6
nSBAFrb8uREe17hd6uv8+l1M8TAN9tBeK+jIFSuJQ6ANIIw1wJdoWx3IfZdmapYxhghyYUjhoLWR
z5ASUC6zpNAywUMNywu9P4FzelyDldvCgcX3NhamZzuvEcbG1pcLBdZ8Bsd7BPwEkKCh+uaXSXpF
1VDbt7fpR8iGCm3nnt7sXa/J3BwtKQWZ9JVvxQMEx+yRzYhhN+smICOkTnGeLehr9kBNgi3E8EfX
+75XNMpM98+GcGS9cUI306e759ohY3DIeBBdA45f9s7+zfJ8BkPS8rWPNBIVfYsUQkI7LgCeFFND
NTpmt7KbiTAUXqF+LjmXM2+5sJaUzHJbPIy9QPeXwjksWkvdCV7dmpzWnab6Xms+x54pIY8lf/7u
DlFHD87BuhISp6qytSrXN1xgoDxWKOJtWZnpQQX9P4Qk0kXj7MV3Ar4tk4fTy+rToTinYvE5yUY0
uNbfgDABKAMGb1ebnPIB2elioSE/4RMOdkScMeXQWdu4bQSll1CJTq5JfeuGLiKJ9ltJ8Ih6X0EA
J6m14kIvRItEKr0LgKtsNbfVsGijQbwbD3oM6JPTMAjctUELcN/MAEZ0haKbCDrMDKResbDQ1Rgv
o+6NoAsXVGkJJGCPYudPhn4RBMG7Dv17FeU5F3lnbXBcqqpoa53rnFX1cTUCQaByVdsmsisFjmuX
zsLleez1gfyanCk/PR6y0HDqDYbkgWVryURoDjkyRRkUC3Wg6wEQmGg6lPw0mPPF4st9b3NsLV8p
/3jG2NQxF9zMX5/ogAVImIvMjc1EHjgGt6LE0qhvWUxwxCwS3JykcbtMwVGLtKWCsj83aPryUO3s
Ze4DpjiRblZlfbMCVe8RMUEAoY8fzjn3KogSMSSB3/DJCrfye+HoMFtIUiXQQ5wDocKZEhAXqHoA
KRqexLmMQxGDV+p9JuCx6Sl7VdKlANiUY9ZbTonaluP9OnAJjIyLNq1gE0zJcBKigiYMHN68Ouhj
9OO3RrV98/Zwuh+FAROZ58AlTeE5Mw+aTCEmtUUnJJWehDmMer7F0LanhhtK1QwlhY+YiEKnVfpD
eZ10xzbHOtdrBN2d1NcriBZoC4yBiLkJyU8UoEfrs7XWOoyyZYSfYteBlyWGX4vmVYbUVhj02flS
ND7QjIMcoZpaoWeMGC+R2kA5eBFreaqCGYaeLqpHFHdFTAm3pk8jlIZjgf0N7U2r1I462E5O62Yv
oh9V/TSevM7yVyquAxTlHgTxFdr22ZpI+nNQzAhcFqJZ69aglk4p2Xa6BXzatfurwEaEztNO5L+A
/rojuZ6qtZL9ZzTD0llnwR0pgTMOFTCZugfOWyOn/KESVpDC6FRraoYcNkAOWbRsFlcn7wrKgxrk
AL8i/bpiOVmzMogMiccx/gDprcfuW1/BuILo+AtZ/iq9l0WFetli0OeHcSdmEVgHbHRJ9VJ0BMAb
2CQ3nLxPDHQQajiRRyvDEPQghZREl8soM0hVCowab6Kg4YM+rV1jWsWwoezjqCfZVCgyTqz96jX0
li86U+27m1hRrJk1ktCyTRIdfZX2YE5Lt1OXNO3Q2zvxKImADzQOqjOgZ2CVBPzmUT/aoGdvKWKt
ofaMWxMmZt/k7O7DgTcL9OM86ubFd8eishTg3mX6MsYny+CRS9B/fRePMmY5hFALfhdwP27dSa2y
FkCewtN+75nPiwXhZ5WpkDFyywajAR2qPctQwRUouUmSHpRt6cYjRBfhJA4uke3TvLFRNBSDGEjz
SZv7IdgZTErr1UnG83KoTEfJxDZQ+wH6zY5ZG1w2YmsT3UvU0Tov5IFux1wiO93V0LVQ42O1QDkW
a/wYrUoJV9TTNTKelo7fxZLRL+nYCE8R0/xCgG4EPzK1vsxSJXgevyX/8wr7J5mebFQKzolWuF0v
zCsrK//4GeS66i7UWpt+x3+pHhQk8zPI9/S113CPq9L6ElQfNfSPzDRP5VFTypBwP+VPavk+dFMf
Finsdwwy1qLTLF+z9CKlCVNKyqlOtbVJx//80qhDN4E+43Ynsm68vJhHDtdccXiUTqRtMIMkZv32
vK5VqvW58rKCJ/RjXy+sC9BHpGgdJc8Aro+hEaUhPOf4TZExy6GBvMIqqljZLKB5niwCwYIxrab5
69iu3ejB6bH/hNGxiZd9tUKOzMu6uNJox+9vi8Frp+cvmgDcSdCQCAdy5kd0dUuRifF1wQM4xTEP
IAgzVhaKdA/plrkKz3hNA777nqmGvaO7aDjn4DKliDIvBM67uAuGBzn/G3oYpuDA0QWKeUpHrqI2
0/50gwGSrX7AbOjbe6N58RGWhaNpZ5dJHHPLUYZJIoWjgZAxcnCSe/wRqeD/2+7/oSj5/dwr1dYK
tAvjatinVGvVawhmuh7FmjwaWqlUPi4kTjQy0kPlofqQnaPwwtglIQNUZ82UuBD9FVuD/equIcns
HecH+8XS/RGyxPduX3WtSpWS1f44TP2prP1Pb0y06QOze1ELsYdiHvgOTanGhFWxi9zau/9Q9i3V
FcpShk9K0ZRqNmQ+LN558vXMe6Sar6ZasxFE5f1om4GLdNTzInhNRx7jFN8fv42U5N5b7zzVCyKS
VLQiRipjy8ttbnQkFNY/a7bpIUkycqzu5RwfWOii9CWauaDrDs+bUBZIp74TnXq6s4ZvGxrDs1A/
zE4+odMPQobIl6twEdMzc6mrwM4k9P6SPZAzt4nOUgnU32Lp0vWqKK/COm2quAL5Co2G5o0uhIXD
MkKOsCrUObtbJg9I4ckThQDPF+HZPhF+UVD5qPiMWaT7l/f8xD7aXFv4bOASZhi/7qriY6/Ev8/l
Mq6Db3DUHQkUr+VL6aoLshmLk5MHZCQaCLQQ0+ucDNkG6P9mEkIQORpgB8/37lIh4KUaZZ3kqsod
yUgIrNH0vEs6MfLPwESUN4skinn5EneC6UrSkF2t1iVzM7gYaClM7NEBVlwJl88NX+MVqtBceE9V
KseMTpQMTYF8F1Pt3UHHleVTsDrZpqEi1zpAPkmmc23RCn4HEnbjc+Euj2cBjv9GtOkwAph1dG/q
GS18eo3mwxd0Nz9cmGV2zndMslr6u1tl0BFKMAlNuMe+IkNCZl2ZPYD3pdQ4lX7MDElK5cKyuAZf
JA6KGY71feBBsCB8W5Fdi9wOOpHyu/c6DfUyBGrrncRWFl0MXr01YP11LHpY2yKRofPKKPm2UBK3
NlcfqR5pMb7Gun5+jFi+4Bwly+JyVGABtMGnG/aLzJfj4A3kb6Rwsmt4peXvIBwFDHj/BmSgS35F
82NkAuWjo70QZGSeuaqhiXafG88LCZUTvFjne+7Nmzwdl0OlvpREpBcwdc6yTHwUFQ4+8VNHPF4H
Zg31c6AN3Y0I5fRDuD2N/SqFs3/hH7TawWsDVFI0Cx+LpHyrjRguZUOYDmKWuVIvRsQDhgTDi2za
vm/6ZhwFHfsLA3+bYGtAj9mX0e+Sh3f6tgSzNOmOWZ5l/FjGFu7jraG4MglltcmhhCjAfBlz7LT7
EgevtNXw+NpQXOsSlEYwnxT4H2D0Lhfpwbl/TGFIWvGYJllS/sjmieLTmR+thf9TFLYF76yHB5/B
Rv7JAhsQ4U/W6+Vr7l/hMQO9+2vlwYkTH+7xX4sIwUNGt9I6GvjJwtxSzDO8Xd7iKQrSpxJyQkW5
qOYmeAZM5xERr0RHsrqUaS0Z1G2MrfJQ1jb4nYYbJn1S94qfsXUDV/OnVyJ9FwtHQz49f42WxJKW
JZj4qo9EFyNeNhTxS566USAqd2VXQRN9azxJ2GitJfXrv2omxJtHGgL+F0F74n6+Xf8NHLaH10ty
UkAxK2JfRtI3SesGUIjrUFP0UCuoH4V30v9IdyqfalM8gp0pa+j3GG8ZGTbFXswSbI3yWIvPzHKL
QBviLCsFpFZrXaZXxjzgOoRzgt6HNEIJkkMACMKcJcaXJvttxtEgn2KjozHVouZZsIWGSmgJL5/E
XnRfptbnOj1rUK4WRY0jOpaA6ZREHzphwjUc0Dk+YvCnkRvXWsnURlH2i/VHllCSaKovF+0IPKYY
oi6zgs1IV/XGGvLDkI7lxhy+Wf5U9VO9pH/mriIoMq9eBMEaogQDDJI7yV0dfkKw2JIffU2dPiI5
ku1jIc0fQGMSDEfw6WW7O6vCUP/cwF1Npp9AUW5URDaPbLv2xwGogn2DqkRLLelSdKJAQKKshQbJ
B2pmmtA5FRpbKWr00XcvFB2d72i7OEEL4p8HjJtLRLB0SNzBSURdd8TmV2QTo7f1G1stcZn0EiPN
2QEjx+EeJS/HmA+TG9SfXqEPab6SKtgE46EDRBxkzIAyFsbpYMHvHvRXZg9ouygYuMF3W3IMpRaX
kj4k9MwBNVcsHK1qkazjziZ8ZUZAxtNvCvwwdc2b8nylf6jspkyuRwxWGzDKG6jbXf/q94MVp+Fa
xA7FTeV0/hx4G65ZbP/SKFPLBzUZ84HBB+lxRu5QuQU4zZQ1HQooQyN0M8WV6PnsHM3dVNzeRLwx
oeroO6WTSnjIk/xxvXTn2HCV/OWRe+ejJqFCiDyTcw3HQo3fwRth3S3PkQX48pBomRXqeopeptxc
TXl5HtWpIHpB6qLIg2rdOcHXvzyOm2QMY2wm247fSMWpGhIn7DvAqlvr2XBNyxB1mHaAiXfDF8s6
zz+MjCntF3rEUkFqFVUnFjovg3Mhecm7GRBe7y0P9rN5s2+9oqU9WHjPWXMN9n3v7c9Hpwrf9K5a
kdHsKjshnTMKcaPHYQreAOj2AT22W1XysTjvB2ie4R8IZe09fQnr/lh78xu4JAjcw/3Nk4ZEP5p4
4E5OEuHE7HpLfEKmHA1MEKoKHkCgZE7IyM5BL+6Gc+PYf/R4VTMKsqukT4QsE+CY8GRv6bxZ7bvz
PCm2b/MZHts1Bla61GUu9AESqJhuQgHwzpBMk6rgGID/70lv2VrvIWE9ewkGytuB1VQuhJC1q2lx
MqlCGv9mr0yInO0GTVUp1uQb3rgnvqkbOqdpBcu3VrC8oyUzXWjNQzaH03VFk/BHF+VNfquR00vx
4zpMQwZQAiHwk3w8jdtvRNiQ4IRDiRLj0R95xBg7Inj7v6qdIc+oqMmpywkEeUFDHI+Wwiw9sYmF
H25HI1iuwnnWfUdSujg+MJ0gJnJ8PlUDqI9jAwjW349n+x8fJNBa2+4ePefJb6nuNjUt5kVJ8eoN
T3imL3r97xBC/2/4EEE2D2l0T6I4I9Rh6uzqUCE09G9JgeXmdMs8puNNscSH32IyU8sEqH8acrj2
i7qpWCpnUcenbC6KpjTd0fgSWA7DILy7PIdonE+YFxWy198yQDnAeIwRwyXCepFQdCJmKMsH7Mq3
8DXoJ1Pbfl3jxPX4kPd8Dzqj1VtRxhsEBLaJmfwtywB6437+XETD9taY81k0D5iT8zsSbDVIxUq6
6aw9ISLIk5xjHHvk2ZeI5OPDl2fVhqveiRVMGPaO6s5NdXdvgyLyyLsj1i1CQx18Q3yiKvKBfVFz
D6XwB0M60yuEpIuybhFbK97GSx/06Zfxju77Rh5VatqeDXD4ZiBrWc/dM3rXK7UjsyRYwFHIZUur
Plpe9ngTK62L9AlqgUIvcWa3WtaLckqAAN0g32laHIOYB7cglAMvpczzpaygso9fVMdmjcmE+Xf5
Fhci3kFdETFkYYoVQXZgobt1dFipy9+wKgvKzSeS3HZzMDxB2xlZDb4Ua7fAm3CYytcPq0wrzS+I
4ce6y/Qbl3pNrVYT4Nb05XR0Z3ZlSzEWsv5JNAW+FfyPUWNJLgDCZfyhWceNjrzuua8WwzdSc0Wu
zMXAj9W9ljkkWrnB56gQKauT6r8+lQ8Mf1LURUItf5uCJt7iDNf9pIlav465kyeG8YQ6yrknfLsu
XdbxehBTboHHb8L+Utc0XJNwoHfriB0p/G87EJhY3GzogHXetofo4GNOXiqryzwieWrqyqAtV2sJ
7SuznfjVCaNJ99jIlysJWyQmL6cnaPGhy7oXYga52k2PB02QhGGWhzlmX7mVRSG3W1rFcBDLvT2E
lXVaBMcnIJwJif+G1FqcSVFqlW2hJkL6bVRUhqB2u8cTNEt3faR7euQx+K+bnmbx+cQU7cvz34HV
0fJv/rAt7Jg9d/MR18QirzVtAVkTH8/LGubz7j1DADNJq1sCrgxZmCIL5Z9c190n2DFW5NMqQAXn
zpOyWINI7/pktiqh2twgAYPLDC7S1F6VlGV9eXVYKuTAyJLtRxswhrEVdtSZ91/2/yrGKBjL1rYH
SoKJvwEvWbk4/VteI1ljKLqD4FSABpo29muNy9USK5l/6e3TPurKDJCNGzV2L7GzM0FIyusvLaKt
ya1xumS2EjI6XpTifif4/cMGE25TdEUeBz7FV31q4nAZNYbdaiY0UBdVzf7n7Xu/5z2WH5sVpD+6
ofpe/XSGrXAcr1dUtq7W6OY0tPYvaZBdNB/UFHc7XXOFJZi9cHK6q/1350TmbsAArHZRrbdkuq/7
ABY6TOO7ylP9DoaPDoP1DIqMxxfOaR1ifJVl2z27hom4EjmQFjIheDXSAhjotFJs8KmnfWG/CEpH
gcDQHEPrq63kfENVeGCeV/X2t7eLNKadcPdw07t2Q24GFWaxRmD8iAAiZ+jEf3etVm6HSjnr8IoE
U4Fj6B5Z4bYICew9xddKitkuSHkYrwOh2vJlstq0gp6BwafcRjCx7JwVpzERXr/m8StwPs2DOH8x
fVRPYDuqGybxvq3AbZbWT2FD2+29mHPDV+QQlFQo2yYZHwHpg4BvYdNyp7ZqsB5Xpn+qD1NmDAFj
fZe3IcvygDUlPx9AwS3aDG3M44q2Q6ZBRZtZaYYthjDWPe2YMXxDKenMj3vT+5zS5O7tCrg81zkp
TUAOomTUCNmtM8ozxwgxkyQE3zJdzoiQWbXCYpyzyhuamfA2jyIdpU+F6u6a50aeywGmYJNlVw6l
AVB29fDSHVlE/MdPm+SvgbWobmrxCpdRKw5MmBE3s9flsemvhfZj1/7m+BI61lrsobWB/IXwvTlG
LITMwB2aCNOggcgHajad1pYTmxjDP3QvXk5gUuUM7qYXacjgAJVUB9Y/0a7DngYx0OpHCrNE+I5/
wXGb3LfvtWYsUMyMjoEuQuXRH3zxsraIrVLbVWAVAYQbDW7LAaudhzdCnq9HNzlcudKO5nEf9/tL
1Xkt3kilrwH1vjUkdwn3LSiyhSx7fLL9Qi2dXVw6rV8nwJt7/tYa1bARYn+tJT7gzk725HBtHMC9
rzPEslIZ3wo5nsTLpA2lry0oUro9ZorMR5qPYItjDWSDJ8af5OU1o3BGh/C6v9oIFiMIomBuIlMm
MPb0+rb+imR51xEnGtA9gVZ16s5LsK2+CxqQJUh+1g7WJmUs7aTTrhMXG0+tMvX9bOgFWGrKLF1o
pID3jJq6E97k7AECDxrtpnfxAhT/AbHh6+0ARRcy9HtDwcZiIXtt2kS5/mVp2M99wRVpqCtg7OiY
Te9Q2y8BaGPOjCbyUE17fRiVLXZlVNJMtENWPbYkN3KPoCQEBsxaze9Enu4/422Ca03vTVqBxhhc
wX0Kwb5uctPbHDMh+SxrZl13qlrw0Gj113u1MmTPSuTwxjgYX7Dmr4ZEb3Wn2FN9H21tCN0mB/u7
q/TH1fhWLGWNpSeaC9cCZmcdhDVTw5VaZgwzQ/Iuu0tQpSsPjy5Ena0tPt4tzUReiQt92YuZEGwp
wlxqmCxEtbukYeFjGRy+Z50GPHmyqm800xpGmMvIZ5jQEBrc9/8Ai9TzUjsJ6aLCldG8RNY2H30n
5T7r/WpPiuUg/qNeNeDX0koRIc2UU+XcDxD99ZcX9mNii1P1UKDh20msPjlOO7ytodsZAC4NBajC
vxIhJpRJcbyJKh3qjTmOSyQ4ShVONfocELSipWirz7FkLdMfDsqYPDNW8B1k2SDEFaSKPLziFEFh
Np/nKahw4LWPUXP4O+HLdx9Y4kPjRXsNkBX2KxPd1v+XZgGfYq0YNZDyxe0l55dhtjbC051DixVa
jH96AiATNlAlv9H6AtNRagch70xVEjTUBuM97Kz+bT5K76Qi5h6NS3Zd8Q9/m1VZ08Q27WkdnWJ0
vr7AFvDt8N9cNuCeIhn5KF8isuBMP9PkAojzAF6OlvgaZ+y/XujzdgafEfJmUDh+vl3qOB9TQtKD
+ujjqLNzOzpfx9QHfetg98wgSCTc0oPd9MszREWuPvH3J4TwvD0SjzlZAtdMUySgm+mNOfG6SXz5
GvtsuemfMZrJObGKskd95j74avtzdKmhOGcVXjp2ul6Vi9FVk7SN0OLeNsP3JeWisCjbBpCV2l1M
5377wwsxoMxi65ews34qngMoYd3zzA3/w0hhczrq8UrtRhLFs8MTJNqzfwZPGjLiT0RPFx01xm4E
qJH0SvSwMrkhZRd6VWZSa19nSR4ZyBe1U7REBt65Vu+x038Fq7LQuwjozURlL5BPBDDH9wX8Ynyp
T9o8Z/TGgJCBQVjUDwj5Z3x6LZ3qBM4CKijc0G+bE3LhNb5sFm87gry3IHhnwqvQqtpbD24CP6Rc
DB+xLJj46XPRoFTgFwboW+s6DL1bDaVRuft0hEUbc42rCD2bFgzYIe+rwT2mFZzEXi5Ugd8YkEZA
hlr+UsOF4QtDG7Uzkuh/uic0UBnLuIl22cCcYpNVffury5kDB2CZklgcD02ABUHSDaug9JY2/sxu
R5ITBQrw/RXwo0FF9Z6YHknEJUw4suvhEDvDZ9JBZGDke0TSqAcGnTRmP3afEQaXVJuC+vvm1ye+
mU34Va/vvCrsNe9UY8DuApEMPOmw83tCffmBxCLl4iB6zlbCLks7rn0u3EUGjyWJ/qq2oKB2p59Y
T1bg7xnnWz/0zwq5joLpGb3y1U0Tu5pGINxAtciKRa0opnJ6FT+CTXv1YRKZJPocZ42JbTN7KXkC
LM2BgEftX/6UkJZoTDGDhp0eV3kVECAMfQBj/e+OnyvOv2658oEKHsS8mpEeFglwuNCJXKMnigSf
itmQ7DhDcuH5BB4vUzRp4KScv1uiQ94YjEvlDfwGzhAKfyqJc87tYGSzT5gnoa1ocHpQgHW/jov/
i+D8DW0C/dw6yE7/ECvWWHRQSrKYEFvAQZZMwUnBNPRSgAkJNvVbhfEj4zoD9NwOhj+rNTLW/CQg
Nm3UsQ6iriBqZEgUoFlHMdN6HD0dd+VW0ptdv9aCz3qFF5hzufquqModzszo91EcpQxeER7vfCjc
5PysTdljVob6iCYfIAZ9zgG6f6ocmyTbu9pBMHyeWuLjK2wapU50LsnUvIQUp6ezr+Qiu8cQ/nKf
HQey0oiYvxOYUEOubiQoRDcX677iQfUlYVuhxSA94K+kBwG0kLbXKNLnARwo6rn0G6n24zt3zzxD
DKU13RP+wGvj/FBp2w2FI2E1K90IBId273A98lgsOt/X0tqZqVy/Rt8c/ODfhCjRjCum/EEtty4m
vGLKaBdEOQyZcyZcA0+ANsLq6ft74jvT4clbAtJBnjsEhoeugqdXxZe7xk9HbKp514E80frtbUWs
Fmd+81gLYiEwSlM99QhrFWErdnMgowq5K5WD+PZEWcMR99QwSOXmuE/NLO3CGmHNkllwnPK3b2rx
ZBcQ67i4LZ9TIabUwkUnovtPUVdKJXr5uO+MtG8O5T/UViNhaRI4+uRG6XkSV0vENjJ8AYSVhC13
bmqsIc4LSt9itwEQhESlMhG5K0ognkivu40oPg5uesYklY8a2pkBKBjFSW5rYeQz+FyZQTHBrHSQ
V2f8Kg+coOloaHMleukfSr3/m82VCWkmh26111ga/mQvF5NwKx0cXED7eIy3dqxuQpI318q9SxFT
hfEX30bmnMj0v/2UbbmpEMD1Q5ecmGx9maSJ28IywvNeTsRwUredJG+EWVP5ReSRA2jWMo1+WdtO
JCLtjPh43ZkBtsd4bh29T1pbKaslbxrz/rX44nzLzkgG9Flk5IYajI4YlfdC70clM6N1o1tNeJfY
h0cQQeNGjUq1cc1SLSzFPqZvnvo4vtVfJTFl/GFLGBTfZvUxXoWJgeXA1UhkPBxBePc7S46Zp5QS
WDrDPVra2XrSbVMh8f5UBSRvAGFGu5+mIL9fGIwDXHr6POERqLDeyVLxK77/wHNBMxXdDMHkYA0G
YOGuDHqftXMKDgVQ6I1wc0tsDc8Ybn5jpICKnBDhkASOqyJvD5D1lOkjlpXqMXGDhngZZXxUJXuM
cmj9G3kHkECEGljuFcjVYqnLyuiC1FunqJKwhuijo1c/wnhiYPgVHf0Yw7+A//KmPjSHch3v4ZWj
pKVeZiQIsWjBOeL1ZZ2vboLVLOXS+psfjSKg+EBdfRSoLMinRq+Xx6dVYLW0S0FgsGAeibIw4H9O
ytbHtF4Ol+f5dMNTPYW0QnEO7KRcppVmcDP/MG0hBKQD+WhMXt4ndK7TKDT1CDEgjbXH9Js26i4s
/Q5V7Z59L3Jg0+jMkJctZ7KknpMplho7lIu3hg1X6uNXMe38bXgTP/h1DCklJnrLD7H867yIVd5/
270tm4yL52/RY4775AgumwPSz5g0EveJaIf9SDVs76EKS+GmzZ+dGUub2FEM4XcB1ZWt0Fy2vsH5
xhpQJXQ+u8gJqSKcN4CscpRFdxJEgIAMoiLeCzkkpSQDPjS1hZglQ3gA5tenN25JmQGVk6d2j6y2
jTRFd6yaR69bAruA+gQ0SzMSIojCvrOHv/Admay7vLiH3b3xt/nIHtxL+7zes/OmPYVbRy2FHfK4
+xJdO2tFm8vUveklqO3gVWQ2nk2K8jFVcD8upvyR8eMOH/FGN4VXKthwbWKu2eM0MRPExWdtz5VO
QtU6LvuYhx3tkgewpYvDRFZGYUcHlVmX2R7SERl4QR+1WDqfIthlNgbYRZMbjHj4N/Jzyjy6uA15
6wzTYWW55FOeY8ACSYmRmmbJP+4AEnYAdhmALhDWC/f2B0CNr3+K+95BT84EF2XGxAQQJSWI8i3U
qL26/F0c/7ex5MpJQHkeDqJIsc9/S1h9wjAe1alyzyQJbbaI9QfzL/BlUFpN8H8U9KNcwW5CGGUA
q0WHLIe3fiKR7niEZpnWinAj2YKZZz9D0nFcrdFWZIz00VJOJ2T63UHaEZ/NCBuYMdL3aS/KA5bO
hjgythCuV6qGYBvA0eCt8dcNaj2FqeWCxgSJWK0Pir2Q2X9QGAyxTULHlBaQIcjDRfifW1mMqhRH
EOyS6z4Fen3O9gokX87OWy3FAlseNewnUiiEKS6CqCCk0uoUkWlyWmgaZSQP/U4MJZaSQgnZRL/b
XIHil1jHZrXQaBmWheWIl6YC4lEFm0HG72oUevYDzl39IapvdEykzx25cGDmbVev0pe8QrcQVO9s
cQkZiSienvYa+V64zCo3fZxaKP8ixOuVrXnqsd9QleBrZGEQlGPkb7f3TR8MleJWzwZHDwVzOUCV
MhtXsXg0Va1hnH7rgKn2TaVVJ5UlP9topsFHnEhsEF8sYH3Qra9qIS++wG2kmPppLBgckaTOzkQz
MFwo+1xyTgAoF0aOxqrEyIovSB8hm6TkuGEn6kR4/vNkeqjPOiE0bJ2OJbnwEhy+bZYgpbwc1lfG
2YK/9QA88YSaUIFGU607AGrwJG6OpSy10eH4YcWWaVcgXIDvrHxa4q2jQHjcSFAWjSdWgN99p9ei
ZcsqNG/7xOjBws2uUpJK+/ZeWbJfnpbgbka8u3PYLO70rrZ23D6b6RdtznOPZivT6EQ6qReosCLW
lot91mjqUCRZTD3yXgRc5+nEQYCf9FUcPt2aNW+dfy5b6y+CeJyd58zD1abLqUOlFfhub/Ddvn5V
RZmSDOOLbV2dXm/CSULB7mBSrIE7zhgJ9G4DKhdPbBc1ygx4t2cB9xLZglyAqC94j5OOySxK52h0
aaewUAq0Tpk5uyZdRPl4ItkXNqp0TpwQA21M/PR6rcqK9W0ILurcZ5bxyPUCXsXEmOVBNlZfMjBc
RBn6TXdwTXTuD6d0QDbXzIXZkEu0pFCSh8d8kJnmwbxyTzZvTZHb4MwTX+XZvC5xoSv7IscZbcI4
YeeeFzXL9wpCHKtAZ3VycLgYx3phxvHOVg09Ua4k2jg2GpN5iXEcjFo1So6ilQ3+jaIB72KtLNNH
Kkb5KJSKMl1zoSas+HM1R487J+Vf0rMYCFXLi8TNaelOVAzSCLd0fbp1FamyiNSDvCnh1FTtcRDG
kNpnsuomlTDRbo4G7Z2V2Xr8E8iv2jDN05UvdQBJhQIxKiMmbtcBTTLb0EO148KTXKZ/6LnTJ77f
Emdcf2oTs/Wr/XiukQ4g0034OZi2iZkLq4DkD8fcxze9zzXWnVi5QrzJxxV2wrQ/VPjzTssa5WlI
GaeSM2s/3GYa9EiFwcBXAtNmOjMRRkCpma9+RFWhMgcHyXnQQaFX45hCmAvwKyFQWjb2iaG++n7/
9/kj04PJKEVZd5XN+Of5SN+lpqQU4ot4jG51n5N1i6qqKQergmIKNnliIOVbjDx2FfIudw/6GRWj
Xg5Znw1Gdw5ADRxt8oVU8s1N0bha7oFupHnmprlWY+E1PrYhpnIczagNscEGTw3B2jtKrJbW0JVb
KpAFxO7GTMr3eCYhMhzCmZtV8hK4smedF6g3NbIGYv8J7K1xkgbytwuWcPxJn4fNsSpKk3btOTZ3
fEKNXVdFKyCs2IX7IeCXVMwVRCqSlg0viEN8mho0zmGHrzWaluwoQ8NUpSiqW+g9veZ5Hd1rblFx
zklddHtvnt5aJOkXcpmptihjZzlMYbxJhXhAReczwmCVwiHjTv/J1AeXzDqHb1CU7smlSuw36HB2
OGdm39qCuBRXtRQwVljwRAV9A85RUAFO/lHdYkDOlg4me6BzneCD4x+/n4Stmq5PL5GRo5uFMjm2
TCydmCynP7ZyRJwE6Sne4YcoZ5ICPh6iv+RXzCmTSIbHTcuhqplhLpA0V2C8ERU6lstlO5AoPiyA
XzaA9J2nyLqXBowhUENM+Y1RhBLt/Jx2Ee2s0YFLUTYccPQt3C4VsjvfUe6nqRGEO51mqvJsdv8l
Zw8pbykYJljcMoovqCiuJE3ZRLYjYuzNjGhdXNArq1paGLYYmit9p9AWoWczvzOc/IrHqfHbY/g0
19dvnUOIOkf0W/iPsGr+RxkNooxLGQE9xWuAwv/bIRWCRI8UuNNU67E1E3HBsOaxXANn4QKskVFO
G7RAVuQWGiBqm1AdU59WyYw465uZK3jjr30ma5OCNQ3w+rfP6+xkGKDz5LUczX6QbVBcPw01ts8V
Xm5NrAmJg+6Bzlh6ZypLo91AVzwXg7dHyD8XLbujZ7+mNAy/FVeeEnfXasWstkeVVoHujfqlkZD3
4307Fv9HakNYCZNgQIvG8hoM3OkOo7dd69sbVDfzHKeHGmL7tdFHloHjJ4Prwo8l6j05qpYTssKv
uojKM8Iukj5uyY6XNDU7jEFNrEP6sPa/lMtvw4DRHt6dHlLyhFu/2klbFlNx+wqfCUpoi+bcvlOK
IzvgZpoHTF6itirtmXjAEYwyV4wbHW9po58HA/VCm0ngWgCbDBuqc089LOjKkgd4/X1iJqId92CU
mMYGbavHE4QqVV/cjJix3GAXv3eJ7fxRPJExhw8WSCSl2GqfOpy30TysAwm61DgFTXePaJakWFbs
wC/bofE3Dx9I/ljvdEaOn4PnII3F8NC0jU/7Rh5U75bGE/Eo4qt+zcZZLqBK8JIv4BHiIOR6J0aF
pCS3MkzzEEvkJeTdgAOvJ9aHSb54PFxmppUzZvCiBxWl6Z97yCimJa8yMEUT000IhgNsuNw+pOUF
mA8D2mClfxIy18VMqsxs3EekqQC6EN2gXaPvc62y4bkK5J7lXsNyfXgz+b177fETPNqoB5eTfiXR
y8rMwooMtoMkG22vomxhe5A3VRV/v4mhvnSi0ZA1GVHfMzA3Mgqpedw4SwI+hElIOjuMeAHIbq4W
czhbGiiWEyxj6IpIJqqmxJKBe/iR/yal51bBPxGIztQZj6Oe2lYkKd2QUSeE80Hw/QYgqbPah4nZ
Jkn93LVaEQEUyhqfO5RKAXFNllGdAKGSqMEzbyGkFhAdiu5w0dd2swATL+mI3fZpFmbbmnXxuGeV
VSklDHxXqaFXLqeiJQiLLYPbGbp9GFWzRqI6ECAKTky4pMLNLclXKuqaYocW8rHuwjPq37RV8wFa
vZI3mlq32wYUiQ6KBhG/iILGRjjBj709U5p4HXFmMVXS/XMu/884gBuMOBdsRuA+mJaA8/3qgNIr
WDCcXJ47Dql7Ys/8/D9U7elIFisyfqX5rMTsQVlgGWqwUs44gm50yVl1Xz6CypFns0cqfyFVxWT3
540wMROqXmG3MdUJ/zDSolng+T6/14K6b2nMNpXeWaS3PjlGXjZ23M0zrx+DzvXr8QVWA5zDirDd
1c16dHhxljC9XsNtkrL5SR9jkTYtvKcxso0em2aFKm6sAQWbvatHIk6R+XJoU5fPJYCHZ+qTkp/g
2DiSg7+HKlGIpSm71c7EW7I7f3J2BhPQlHXs1Gvxj3HGPj6X4tq2IwC/qCw9CwfqEPpJjLPwTfPC
pL++gEqZE3w5tDrjjWGVV1g14/2q1SB7Cmv59gpAGZpa2kVmTtyZMHf0tPDW6UUDaL67xiNkKZAM
vHlcZk9gP9nKlOADVibhsQsuNj75Sb9/jgKjSrbi3XW16x4xr5vDLvgBbAaWiMPmED9xB5S0iTtW
2iarFTNyXjHhldTxQNOGKIF5zFMevZnrSIEgDfjpBnHixjhTFWoUmPiIvYzT/lv5QNSeNyn4f0qq
7qEO8f9a66WYMvcg9UHcJTqcIR9bdxEd25X9d4yi9NFFMTAB9y1woxhiGh3D8Ol5arLVo4rjSBts
ELzt5JAHplL5R6bsFUeLbz3quk2hLDSLmhn7iLbYmPrW7gJcujktKXzLEx8ZsCwIbSrmcZb5M9Mg
0i3mrVmxXNrhAEViADVsx9YgTKfzd2jpHzFRkYWl9ft78Fm8ItEK/eMAn04tQ6sPerWsN+9vwlEm
c1+YoFbN4ruQXLvr4BxXjxgAR+lm1S9mqCfO0wcEGT71eZz3nheK39df4v0Sk/8cqnYxn2a4A3/E
5HuQeaRfoPncUe/CFysdIljvXp6fXqla+3PoOZD/icubVh2t9x6Qm9uSVia23THm+hh6ruB6J4yP
A0I15XBgy8w3nl++Isl6oFrOENgStXYZQXV2UlkNd38NwcS74g06m6PPlxmHD0lLfn3CGiqh3zDi
i7guxZXDwZxSE1rvmildWvB0gvnSy7IAIQ1EMd9bQal56EEJOzu0jUAEPYA90S1ncuEpx8HFLsGc
lAleuXn72PEMOQzktlPopTOKUWu+0+5ARMdZvlL5LHG1jxts8kSsGVEJ8Ah+dSyWyuQrCT8OXw9m
2uq7gB9mJbo4wJdGkMBSyughiUquLnU0nBADHIKo7EtckErm2rawHRQ3Ta9UKGJp/LJcpC9xw+lU
rrT1PV1NZ8e4nA6o/yCqJBtWFwqbn4a1cSlwLJlVk7viEF6+nCoydrhGSXKxzR944m2ygzzcUsgM
jLXhwLQW6X8pkoQROsnmtlXuCl/ASDN2ZaLlVHIUZL8pxE9BeUxjfPPB+qKiuEmb9RN5wWnU445m
V0d2wXJ+8JpEh0c9cmM7enqBHRK38qdIKq+1Yge2X3w6oTLlsXGDzy+GesT1QDNEyodRa/jmbg4K
ALfUuABWfvS0I8The33qgatd3kLtUh+aWqZ9GeRBmm99xt+Ny3SjgLmmhcuQg0i94rCvyar5O7pw
xNxRLEW0wuRtjMdZbejjCBpRtZpHzp1moRxkqKStBOIJUfmltsB6c0VAJE/QMQ+IOrzaKnA6+8+J
r1iqX1YzBdUh0MxAW9zdP4Meji67wf5CTRBhpTIAJQoddhKTbqQAaCqnGFzsNBWgWWPZ1urP7thm
3xVLX2geggsSY3ynOTl5/aydpAbivdxufq7y7QkqYcKLJTLpT9KgoQLpB4z5XeyzbVrUlqLLjb32
+8luRvXiKuM+JfoEckUBSQNRB6Slf4A3ndXz3cIT5I/JtaN6kr3XGjCt+gsXIbMXEUBZYuvQEqAe
ppfi2ndbo2Xn34NbH3L/3Cp91WkfddhOjkbxIaPciAhY2y6LGMA1IZHd3gW6D3aziXWPcqo9nMUw
PZQC59nTTC/XUosmYU42l/XRADLK1V/QdfJVAgJTROE3ddl9a7LISsbjwy+mX0804KSgr7joLxFT
PTabxZ1oHh0Hrb1NwcbMcwW9nmL1G35w8Fnq5vKebHkR7eaDWOnNTnULcGJQQRMmmjsjkYleJbcY
PgFut7rJbRQn3e59xsVYhE7UC1NN0+Yo0WYt2EcTr34OYJEu+VPJBfg6QjNUCbWhba8ix5nAyT/l
1fKgBCMMC8WOJQbsGY/qUwZWIAmZZ6gVjTjNAnERzBq6XiUeHhDtnMWQOedp2A/i0PGJ+JjYBovj
w6RSJdFRWI5Gzdgg2t9/AhHzgL4mcxMiKGRqk/ThwMt55Na1wjupoa5bbmKla6xQs+6PzczfkCjR
1fR94SJYJYwrPWq3ZhR573EbOaZSyQi7uRB2GMxGDeEw+CDkYJ7AdXylQpT6/BqWCljV9SYoxKZN
TGscqxxZPxR0Z2uci71fGSlbU0PtsFF2KkyEemjjbQNkoKPSdnGiP/si626ZBDjOs1x5m0eWVgPl
1Rm0meUn6vJdHFUjBA7nRNhNvodQw63V+mONKMguffU9WUTPhkhxgMV9XVieVa+5aO2AVmaCpkH4
iKTQWPrylsBH5fE3C7dQ2W98wxRbTNa723UamrWbdas8U/xf8zy2FpZKOa544k5Hz6f040Ib1vBG
YRxt+UjT95K8xkkImnIm0bfFiqRhQ6AEwEosY09lUfX9JQAPLZC8uiLCo1WGdv4ZE9uLfw3atmNC
QtNoDT7y4fYx9PYU9EKjLQ5D6jr2QOh+GrnZ1B/N/DwyeAPDp46qBdUFok+gk0m+jl+/hhsLeJU3
ZbSU/wl0PaZgbkamd04WguivE4Cltk0Wzs1bnQ6ExNob8K4YXXiqT2TwQ3Hxn4y9nhWCuIPzNnZM
/OTAUmaT+TbS7u/GrCyIrYN7P6fAZnHmXXWLaE9Oi08OqATn15WHbJDGPY6b2pXzSs0EDKYJoBjj
yA516WD8j1eq1mu+bdG5V1VFt/nedZ/fBmG2dURCRCtysUmKbRkBRqJmoqisywDd3mJNtBM25dj7
OKqM8+EWvysDLQHdXL3OIxBfMLJdDGKuSIFcBJsJVxZgtf9P563N+Nmcziu3ZG87u9Si97ONG/8+
KnIyJHvXMZ1iJYUrlyPvVp7wXDf7Z8sRBYA+TaniREpmfOJTw7zyFNPHXjEIx0AcjjYQJZ4zfbvJ
ITZqoL8R31JjnjM/CYa5/ZZAArqZdI+IgDEhEonSVyTsQKLyxHi4/+oLqAPFClJvi4KfOtdwcsJY
wdHUYYsVdn/sYZQzuFbu6+GYXNMxVkzWDDGYRUfeC9bCpLC8m82LQRxV18XT3iqdpX2txRZbfM5N
v1KUQbcL1umGPCg8a8uk1c9Cfn4D2xV4QP/N068rD2Ay7Hs9MtLtRuepDvPFGbSSTVrAMH7ryWH+
Y/or6EP2KuCn+fs7XP27CdxczT4awFWAkHmxY/RoUyiOWKJeOIkkwuMS7m1g1MA6uxBUqzm9Z5+i
VLU5jcldxA+EX530cncJMOzbK6qWXdh3apoltIQKOkntLyqlHu6/17O1LTczBXY3PZLQSlgANjfR
q5Wg/xBMWdi/gwn//COFHvJekAaOS2GZ31+o79WusjQvxd6OG1KEd5rwU2da7sJ0f33ky9AfWEja
r55/+nVjIS9axp2lSX+YwTqn6UsIlT/N8N37f6ELbgNg9JIqbuZYmrk8edxCW6kQvszsvq3gJEqR
cOO8KnQAJ39osfUtlGP2D5ff5fOcTkH6PMFW8v2etHpm5zPivJGc1KnT2t/ep0o0AHFtkGul6Eez
IVeKPNWIg1lAT3jeZ4Wb4hhHkBBOQX8LCeLg06eqWsUO6frsef3+vhaw+4GSOTsOX75L6C84PR0S
kR0toxex/9L5sM3pTE3NwJcMxJwnI0cz+NnGIEWUHkOnqWfXh2wa+5PdUzQWto95xqkQ83pXWwIj
sXi4WbVcEhS7wNkldM/lVOtXDwLeSlUGvvjT6FQlEoifYV2WywDTFR7uQ0vbbdpCORgiSy2K34gX
4YBNvWogBXhm7Khjq1DAkJUzeZ4PJ/NMpYjWwP3RbDpLlc8r9yK8PrL9JWcIo8MX+3QnAUzCnAws
pge5zJbWvDpZrp5+bttr4MMynOhiBtYYE3J88GFS/YCZrUUbPmdgR2kUzIeZAjQ+V4V4AyZMqpXd
8k61SXjspka4Aml6r5/HhFbFMBB9SLvGyDfz5fShChN8XnPDTdBhMmW0G23PclPhhSjqQdsIb3Ml
f2VWuyHi/7h+MVUG1pG34SugkGh6yGLT2nQmrnRW5A/Ws1gWKpUuxGIAd143HeImcfA/xsT4JySM
YppOQId1Mk5zycXTIyNyzDLTN4/CnuHTXeVFC9ZZ7SoBO78dHC+6A30LOF/JhlzmzuuHupHMmQJG
ssDC/4k46s5HJRDpi8yaXJfzjCjVsC+Saj/PRJdZlKnpP5/+3z6GEHQESIzJQD1U1myK4zT7n4QN
HQOBY31nr05I6SqIdBF1/GpfwLi2gL0HzqeGRdk07kuwMj47rNG8Dmf/a080KvYTVhLUOWWlHT+1
+M02ezSg9EQnxb+Q8JHi4oD+3vrMPlQMxQC9CQB3T5WTv9eQd5M8nwbJ9gujpXhG62EozjvJgqRs
I5GouSpzO7OCEfXiOE9HuLy5elpTpf+vVahWkRqZ0wSGEVH+4DwNkOQ6b9n2OrdHPyKs8zlNyWVY
U6XoJ6g4nk7CaIKKufgrK3NbM4GxubiAj/xR7dl28Jb1V30+Wk5jWYq2/+d7gQkwjA4S3wIhDbL3
F10mAs0n6UDtXn6YbZnD2CzJlLqMNuRPedXGzuXOXeVCfAPcjOsJ/gYuNkX6y9k6sOsaOWX821dC
iRAfPL+9RYEtYZkNkgiOf1O2juJ/Zsn6Czu58eZ4qAks4UhJMtSuvx3pkykl1E6UoDEbEtP7ZHCL
qGzk4HD9J2wrmtpR7vBN+6cXGdMfyBee2OLkm5OUn0l5pD8oiUpUrhCOIBs/3hqFSMQgA8ZqDQeL
Ax7DgGUBEF7PZfTMqFOzI8p4/9UdIDNephWN4WjI8nJBoLcqxFivXOv9NacUpqbdbRqPSxu9CcTi
iFVWnNBXGQTFYpXwojSIsX9DOl8QyXe4PIig0hZC9PWD1IZTWGA+soKiik3HVs7g8fu74ugudF/Y
zJXUHprb9KOlUcPW1JEWxAWly6D+jS/MhGqxEpy0d1vY//XrFVSI9zMvQ00FWJ4C+by8mIGBODeG
y7rAGP29z8Iau0G64PqBBjQsymB620gYcloJMdsRp5fj5ssSoWaT6ncBgva78A6+fV+7Ic1/JKH5
LPMkYHWb8BXVCtRKUS4P1Z1ut9Q6Zcv9hr5WCtp/g2vDdiG4+ens5/FmH2ixtQkJHJUE2eXvmzAc
M9VKNqGv8/Py7tsvMEn+SMluJwgB/KTbn5Rsk2jrIZRWpBIlQqwgrhV1yqwRVHh9h8otkCwg6kh4
pIuOTRUvVhm8OgqQIL43g4mHyGzfAIosdO0ffYj/zYIa5WcJ/Jgt0uxK7s8+h3Ei6lYSSM9ctis7
/qIjTsploffDHY3o2pNGh1Ue0lRLD/2oxfASfWtzwGy5o7JsfDDOuapRV4tCAdsll54+0BZxlQdd
KIDWfWH3bMg7qsHF/TnSdp+tGzbVpKwPwrX8LYY6fbfnn9HpaTtmGih0YQ6xMgZvs/JkXzsTQ/EU
GIfGZfcrVD/pAAtBOF6JJ+H1TfX4ndb3J1ixPbwqXsrfYazXAmyYwmCU028v04UiMwIuHzUfYT6i
FIvSKA0jlyX6b41ZBltW5DMCAT500qnh6sU9tOUkkbsJsKRNreKafN1BNQF5VcAJ6D/X1SO4fP0a
5C4+4cJyuikhmMB4NVGswLD2e9DoqTC5bzmAE1gV3q+i223Fvu1bZbAAw4jmV3gdOC+n9xFbP21T
wO9MH9rOv/YjtfbDxlx1H4w0zyukTDKWGKq0aJhkCJTcmiG7gG7N8rAvql/itutpMoA8V07zFz+E
TI+y7vvid6uWiY8uDLLDjcqFuBm7YIWJHdbMlvgPUFgpXLusPMTpUcjut4d3UMD7cQgh1zvo6OB/
51EXH98GirdG/tTRx66W0yT85il6ZkB/wd+zE7yBEO+S9/FD8EeK5Dsk/qGKqGj0W1ICnryt5LJm
CEM/GwwKgTvEiDMOxFVMficYYNE3hefgIjWrksw6J8BM6B5k5BbFlnODB0OlwCtekKCppJaseB+J
wxxgp3k7FXm4V1W8lPXnyeCS6JuXn/jUoAJog1RF6vDSptZSTu0jlxQ7/zUO2aRWySV8o9hpzNXL
OlReLnPs+uAsyg4PIUY7rE9kf+AiKrDHxZzr54xdoLaHFry+L8/mXcyYYbOYwRNhig922fRL45Sh
LMm2qxETaq2hRj9nbpW2ZRoxLaPV/kpwrQP+a6MdglvIF17YVNbNMW+X00amZwFcGzy6a9YcA6rj
ysebCcxKCSgRBMnoTQU9BlEV/dr6q2QBmAp4be8PabYhGIE4AyBo2zVxC9vipUYyGUYGuo/Rgwur
tCKsArm2LicCye4dvkHSb3utGr/SQ24fbrNuv283p/GFC04wovSPo3sCgWg9ImAre9cY6xz0xhV2
tLyDK/0aH+KNozjVr4Go02NalNjZKEjtNzCpEQWNaNtosIqqgG+NNNUh13pTrS6YwDwE2SIY+pzC
NAViuGKKHmVMDNtaHyIkhzyY6Iyu7m834H4GUfSv/FXVEAm/adgpD4L7GwRC5AHOSoH2iXVh+Q7W
4yc/JjW8WmchmVbaHdONDNeRKXlZDg0fE1kmFsh6PfCWx/K1vFj4Y2mhEgg+VuIPBGz2+ktFQKNK
FPDfm0WfhXgMURKbv60RO+XHreeGGujv0Fpj1VEke8VgWCzXWuZ68toLnZgX6RUCzr5anVh8cYBT
BM4+kDjd9O4o2Ugl03E/9YdIguFbys7sPYdgJdTB7iFpvXLEU9kbPuEwjg1g/L7VZ/LYDNhRLn5O
Jpp4TvhE/TFYHiLINj703rPrI6a2hpewdgp6MuhgmzQ01fmvL7Nq/Gi8drqc6kIMcBHWfxw1dxGd
J7cRuLQbR43t8cC3LnD7bgoU9m0P0dohHM4qLH4zSVz8Mafcf4tOLzzH3pPZg15KbW+ao/Xr7icQ
lW89I5ht8d2OXw0lW17ZYitHu7PsbPCzBo/7S3DwMtFahMKd0AFrvY0hzRpF/isuqbfRqy/VZufr
/xwC8Z1Jbwg4O1Q39r9g0pKWUOmXY0+7OQc7FLAW6+nPi+8teluKM6teDcEHXuR3oZZHtwvmfozP
TgiUoBA8ltPaIOV7ofR7JKQ6VHCJVwHucuvL0FpE1gSU8ssKKq84bP4UwOkg+Qd6GVuDKIYFr2va
0+TW8128/PxQ9W4ctEDquE/boCYgBdXt+qpXEkkqZ1Scmzn238iI/5OSzwJZGAqIc1U+UaF2IUyM
kwpAfDDw/8/vauVq6lK5AZNaMLSpZP4kYZbYXepL+QKmLrt5ZY8fHZameA8xqxfX6Wr7sdnR2nb3
Fted4GwkQJ59ULqy6M4a0Sir72HkR20ikShvNblApKb6xL7PNSU1dBiD9M2rGdiPPMx+g/ajj1y3
7iKeDEaxyxWbx6Y93zQHiZrwZ7ns9qiGyBH+V/vN+I63EBXGDYsc3gYw4Gofd/ngXAusyFDHJQHd
L3oS/9Izs5vfSW9zl7WWOGThSCfKFLi6xmI7dhAgezfAHKuxxg3hNfyXX8cZf1GpE3A0GXEhM7WF
0x9DS9auoiRabXsnqAO63ivisppL6np27swZlNI7W3BD0kyQ9MvxBPIbpssnIATt7fwm5+CeqWDG
jtt9lzZ57Ps1XAZ3S/lDte6Vq6K5H202Jn2K/DGxslK9vypZzWrKm0d9VKO19LwoZS+TLEYe0AJU
PHnlJ+OkdIKtSW+8qTPEtmAVW/4iYZpsVSLzVxzonw6Otlw5Dm1ENM+mCHoZytsgpipo5SyKvcIK
kFCVKfMVJU8ps9iRusaId6YODbD3B5YHhsk+iSKiowe8pF3D6UtQp3d4I+mJwYSpNcCrIZceGA47
XWCy24DU+EVSc9nZQWXMttpCFQguz/Ulc/sdZOCmaBEbexY96oZYqe+wQI+pd1XreiU+eG3rbrqi
SrKDwvRS0ezrylmiuLQOlPkF0IsnBYYzeKUKz+MUusAgXxM7CpOhgvoJHbjLuXnJBU9w/mQwxx+d
kdWyuG1OxOzb2JObVzn60dMGvQvVgh4cKANg0JOElz5aQKsmWMSmNm99CkopxJwE+ynDHmW6uW/k
TKPg1CR46HVyoA8T/gMWBcqh6OuxU6cs0kqKYU8GrNfMxUokQ794lCOGz0RrvSDpHcZ4/UwD+Shg
681CmTWzX4iJWazFOJHaUnNl+5KbR93ZKc6GBLD12uZpfCejZDA/sTHcdptc8khVlp7KbNMgytTk
avmhQC3qqtnED9a//4dAcWQfHCDC+fAPAYUnqUJING3yvdnZXXUawqH6ZvWbXPbRhytHt//fEdvf
Zzwz6HRHKQUJ2voIaPVt2fvS327DcDuE1J2Y0+jr++aZJHkd8nrKAI4nOMfgu2txWB5Um/S9Cx8L
SwL+LtiqnwUh87PDvC2f7SFqHrrT3Dpm57B4UbUlPI6UxGPZrbXAO9cWtaPG+6xmKXZl8tYRGzwn
WtxVKZmnoS9T1qFRuMHUMANCDNZ8Ho7teJXVoVRT8lI71ny29RSXG0XET6CHiomG0YdejgVT2XbO
+woQwafo4pey1UncfW+K1MGAbZvAEvON71rMIaYC0geWsdWzviKwn0bxakiCO9Uergvj9U71mRxh
7nQDDNP7qWXV+1JRdFfkRzvHkzlcw1zkOxegCLlVAjA1l98B+K9RF1vSXOhw2syGJAY59uJHv410
TDR7SaShFuzIS00MOGs4y+XvawHp6vKolui2C6CrFzQdqIAfEml0xq5xpv2N/dDS4KSaZKwYOA9K
rMPwEga2WNqEhV0vALECHrCtN7x9kxIDn4kjsgYWXnWfOqjRowZGrDzzdhWGTc0ISl4aFspLtVW7
rpRmTNmN1YaG9Mf3yL4ETCRJf/7VJgcQu9uRng2oGXX6NtGKUiQliaQR+P+Y9xfvjtNDhkcmBTQN
uS+Xagwl9jiADNIYWnkzi4Pk7Zjv+v8u45nVk2TPjnnbxRp4dkncQGhtkRJy0GYEdYv8Bi+8IswU
j9UMaGGseEpTkNKerVjQ66Jp7+apxJ/wmnJHGTOHL7nOlfyyn9p4K9DOWx0vWsq5FG1euLY+PiwI
qR2+lugywk/TWnJ9snSCAjwiAXgtm3Ilt8fRHgwWdpeJlUi80znD6x0XBVQIxEFk4McR+uN1QxBu
5r9VIFlR/1fVqfeP4R3oO/nOHcAaNKlJZuPzGQaAXt+X8DvpOqAg3oGSbz870HC7aHXgktcbajJr
v7AJCVz2pdqr5Qe7sCjBxlwrP+HdwDAyqUbj/CNBA6wsfiJHhuUTTbk7/U3zwcWVgyrm6gtParOl
tG74b3zaf4DUwQmew53847gs3GPfjXubB0jUEH/v5I11hoB9rYobboapKrVoe/wgz4obwXnHQNd/
paPAvSMqrmAon01sjsw0mjFYnWtnYw83xKZPFJE/PIU9NYrcixJFToRAt7IdVXbhBL3Byst18Cq3
hV9cKQIaRzvgJ0Yv4AnWCqUIeO2wB+5PLQJty3zT09rfHD7cY0rBp0XMx3osvqepWItGvMImgyBM
kRWiL+TU2PreltWsK/JpYDe4W3HqeZs8SMMyXrLmySpwr4BJk+Zrdg9A/CIKWvSoz/ThDr/aGnVq
VjjwKmFc/+qG+94P+fey48UFEaa+y6L00gKAOvC9IZ0Xo/b8av54GCANHCk45te+u8G7h0DM6uwS
qnUQdV9Zo7HoZFfd5iupJKCUbA9YHLI/rPZU3KF10Q+CXLRWVOZ1ZCse3l5me4ZFYs7TJAoV/uM5
CsCAz/jTUMItFAibjZZ0LFUawMgxxkA3nVYClXc74vEl/mVy3opd2Tr/MsnGnHqkTlNctg0TA3nZ
7ETEW8LZuhww33oCbQ8zEPdVi3Uu5c9zJ0tPlzlu5dYDGxI/r9065Mw9qpkZQWTbxlbBqMETSWSa
vTN7Z1DFZeAAwho7szb2qwiFSm0jiyM7jZsuAsXSNk/nqxIEgUIbEr/+5hAgbf3Bg4iySe2TlEj2
mC3NH5dZAyohoRvYQ1uS0wr/vdpYAQUA2m05g9O2r3JbRFS1BqbfaoXGx9m14ifeJPYJrDuwno/A
AIZrn50MZWMNSjObT3KDr1PybLr5X9EhcdBuMdrb3o6k2rWbfq8gNRHdivjtib9MZUYHc3AjCTIF
C7zSUFNvslMk+O4daViu28/zD92GamUBeTW4jfduOPCV7GBGzl6h/VpoCIOyZzferaRhf1RiaW9F
KFUoA4FnM3H29COnpc+l94Do1+7ndBT56xtPIEgBKWpYe6wPfRoyoZnqSPmuTBSIuKH/1zo72D3C
afSmLFUngi0QVt7cLO97/nWwwzK8DTzRuaVqbYncFO0KGoY47Fj8k+30ZlCykIDp6SNzspDusJ7A
lwPATkbeshxbJxsiYmSuZFZcB9vVanoESpE2iw1+EE6INY7oIcT4By5tmaL7sEuZkd79Itv96rdK
6ntmPYha40hgtXfr23zCBfKyYIhKOdmm2Ot+ujtp6VJEWXptBpfGLDBMhwvp7I0NRJfwqGJ5BkGW
YiPWoGbWT8m11nnHLjpkWRkI4u1drBFGkndREPIwFYpuQXUvdeDWn/0b9B+cstDBmO7GMkZ9l9ez
Ew/nHjPfAEX7JVR128G8e3pSfpEqsZ25ZXQ6lkMIaLf7yx5166z45stf3BdxxB3UMI5W4muS9ykO
78LcBfuXaz3yhb7vLXun6Uw58CZP7uhPkh/3bcQGj3mSmjR1VmX75nYNuSFKfPwXrPfKG9fE9OBz
fkJEuAL0EJACjZ6maK2pBt3Yuv3H6RasXVRXyEmSMWy2k3vAsBBBtLFLhXLjJ2geUf98EI6/4duL
ASZLLdkNtCBi3uAss8StHVeYpPp0BC5fJ7zw8sBhaSzTbP+xPjKcG0lpi5IuBg/zmtNVnYPFI1qj
xdRxuA9MGF5ZqkG5L3VLH2lnbYUy4VP5Q3O3GgR3b78BOdACSU6vqwX4VK4duzAFg8wGMThapJnm
BBWgQ9Mv+DaZomRFvPP9YqOHk2iRtJ69W8Quu7j0huIxQwmnKv8CqDOF7A+NfHJ4xfOBvfLWxmLh
cGGuTt91o2iUJ94n5qEYOS3umaauGIETMSuUZI2OG1NL1oT0nd4E8h1cQipsABag9EbYgFkOcgPQ
MsFpqT6eTwJGLzgu8LiIgGVH1AB1/HCSRqRRPuokAFLLRgX+cYwLqK4Qadks/M3j9Ajoak9HUjeA
5R+zM8atIUkrsGztmgRuOBrf9pluds2cANsVFTmZPx8HUU239PZgRTCwcbV03rQ/B9BpVZN/nr9m
be8dPXgMI8jlJZfLPYHOTDMFfaYbSpsBD9aniyYdNDchjL0qc6SidJVVPTvGDq5cGxcWLwqq9JEr
MEK5zHQ0xeCfOQmNazpCxh+vw7UMIsoKfhvycHY7daYmWT83qMNqHQwdD0wzwu8A4DRTiOaapz64
s3qDmgJBSznAnlY3inBMrNor+m2nrVbRHQjcJLi7/9K8HQ3Fx3SpUt2b94/6nPiVYQnhROTP3q1G
UFnGdhx/+PwcH+O+43Nduu1LtMYfJJ4ucMgJE0SrMGCLHFKpL9R5EDgX7w+x2ntMtSEyaS14Smid
eIC/AaRtXHS3MMzwVljbzljTMcpieBwjM/IUZkUIqxEN5GqyjfA028Dt8LJMgvnBE9/zTXIdfajP
h+SkHpkNOVSMku3k3q527VucPevbRUUGjYcSipgXCR2reirWQA+1m22erZY0nIxrPeN/eszsMabl
IlXGh5IRF6YjAjGHQq03RQfEMk/giqdTHR9+eHcJgV+AOXg8sUku6yhE3Jv10mJ6BJViFcgs/jKg
g6H3i79Tsjr4TZsv4MeYYx6r6ghDecM7I8rUPDzytzd2XmyvLMF1AaWNoMPM5f3EaWMPEPWgQSsY
g7+xsJtnhTu9SSYNg/KMzCYp+RrlA8aC2hmoHVcugd43LFjbppHTfEB89WWFqLAPsaRlsjufTjA5
yoo7btLpmhlIADB6j4+/IzUSddvlX13kCoee+6Ct3PwwQLuimnSsueMAUJLvm/bODtlT93maYzLs
jU2/AfxdVZbG33f7lEYAkam8pDkTDSdt4unLrWCJrTFomhAanE080sB76GtoX2hE8vevm9xZCpR0
m6AE93fR1DhbjXgQzDCnRId7zwR+HD7vp7iuy8QakDNeOCp3INsKaDDaeJ1ThkHy/XjOTdOnAAc3
xMcCGj0VEWTDq0+lI51NC8iIs8dTsEx9RNgr66oToL31SdEpgiO4KesLl3lJEhzwlT/q17WZ13wn
si3FbV73pbZPtcSj7rQnVbZn3w6lu14Q2/ttruPNBtzIasDgbgjkgsZEJJbIwscVnhHaYKjKMlkk
dJW99ZdZRj/RUxM/ebDVmp1WGwbs3sZACWLbgCG2rx+IxUnz+n0KO2tUagxGvOsCd6BtQo1EOlSt
qPwJZvn/crBYeKEtSeWw1qm/z7rocxdd4Rh5dsGZm7CNzLqw20oGNuUkK2I+Mmrqom989YbapcRy
vET+0+/IrtrlygV8O0F1Oum2zGvxNbUNCvwDfBXI2pK8mZuP9iEkyWfjW4DtPvpun8eoFkeD3pBb
mJyqfZq5l196TTnh6OFcKY+rO+kgZj+hWsXPyHN7RMwSv9duWU5VLiKkzB1rZ8EwgrORhyI6fW2n
5h24wQI/bDcpihR1/dnYXK9S8v5v8eOhMYMA0kQhkaI3xjEPppkgsoYbHOh64P88OVJd0aNV6ZkZ
aPbeRQJCQbJU858aFIMBU7g29p6bAncISEWnzsdz5amWZ7+ZI8PWgqY11nYcJasgeWVZR632Pv2r
ok/Qr1X6C06hWM8zAGXxpF2LZqSvmWXx1a8Zx0zuKrsmfWEATli2gRYD+sQU3QKen6BA36PtmDMV
qHUcGkqT1cFLwfp3qrNYt6zOnIZegXc8gd6404T4mCUpYo8OF5BoGqm1DA3KfdRhLvn/DpcPuItJ
T1toMEvmOcXTO9pbzf/rsYnYZVey1GjX2eojedFDO2u0NDfXUP4O+xvtCtc7uOzyc5QgahlY9AZ9
F7nw5yaRDIxMZhFWlJ6HO/0F6h/hIwwWfisc3yPc86nUgHnsiOU3yRME7eZjSM28XH8nl0x+WNi5
cT9xXEP/0iqcBdKfa7NpvuS2bF+H+GATOPme3bd5Ik1X4JO/28fJgyVJ6v/qrB8G6hpZOmAzOul2
Qb8fN8g6Pr6cU/w65uMO8vCkcMAe9HIMp/Rssj7dRtleqAHN0tNxnPek5n3KenTy2fLRqfuUwFRy
uRz4cwJSTPWsA/JTCjMwdwKvRdjhB5GF5+cpUodd868tp6ssZyFO69jS6iYx02UabltcrGKNoece
bFSbPjH61bhtcIVN14WiJx08y53pdWt/QbXaRlzYCuf9BYpa/O1NjlhE2xNUmrujBukOu6DhJ00v
BtsFLJH8OO7GYPJBzZd2yGCWD94OljEfbbk3rnG7QSuDHNnJwT7zB021RVdb39yAvOAAs5czTTid
upzFuiBFgWgIJsjM59upno7cUaBFw6xeooV/TVR7WnV7hgIOFr6kAgGgBrMbF8Ls4SqtHzmNCdi3
bbiQ50Icr4NQTb2nNQ82FPqYPVCcOC7Zfn/y+SkM50YOMEzAxsNQ35KMMxYEhH7tEuRL408I3iDP
D5Kp7hrxsxIeA5a/SykV4wBh1yjVht6QIM+i0GbxmbMfr/vYFtcuHZ2I680I5/iHtbZLHmUOszJp
EMLzOkvIqFdbnwE3Ylj1uErimS8CX/u3ea/FXNdEGCdZ0HrJ+IENs68O+hhGKgiQZULR3JVwuapJ
qunvYwwdldWGLIbUqP//WcyFpeMYSHehhXhUB7iOIAwX4IameK6vmpnzsmimEzSiFDDKgbvZuj6G
Ut/38ptj5XnSInK7F0I/oMp1o3pyJ9laKBSoU/llGp73wB2NMLP6jZx6Y9VkgGk8McwRWtVHiwja
wNrcn+S9cyQY0EghE+jvZP3FOdDI4lW2iQsCpWTcvQ7bnzb1gtKUHUY1XBE9lTppKJrEPIByfwzj
M0XhMaCvcLPqHHkmQtNwokZtRmi/nfMX3ErkW9eTg6uWLda9Q6aCRBaOc7bBT5RCjNEJDwDPBD/q
bjhkHI/M5CqOF4Pr6A1pY8EHdbWr5Uux4yv4ltrJ8rwY2mT687yb2f/EHYli5M2j7DBXmajz/EU1
YKZsvGukDpXzNH3tvk7y8kRp3YS2OCqsbR5efgSz1/VeVcNnRVCx8PFdimgDOxSU3uYzjR4jJR9c
MfHF03oAHw6/dHWf5YdRNWEa33VXGoN8NEXKUrff+tzeYECnUPdseqovsYI+6pB7xaE7SwiFpKyE
Cnj5CQ8SUH84OOPaHMZA6FNBXIuji7DyvbCJZngDpqS23liqQtX7CwEVVNSz4gfjBAy9nyyvu457
fDLYhbza/KZ1VKyfAhcixx0qAy56bQjsnK/g30oztuUreVjpmA9M1bAc+9RLXP8AXA2Cj6FHW8uR
QkToVi67pXdFOSJxHhStScFn/QPdIDphc6WcRQpuEkksyyaNCnZn7LV6eOKbDeuO+1JBJuXsYTOF
j3RqeVCiDqlhKv7I1ygm8d8d2hXuscFaJyz9O3UAR6x8qCoTlS8nJ96J+W2UHgEyXSmYxzdWGOg7
2vaCGGPB0DJkoJ/mNhdv10qAETOCxd74xVqQRVxAIzl+0PYne5ZunYhTAOBDR43RnBIae9ED4NB2
1NOE9IdThWJeNkgu+/hxj/k4eRSBSRROCtSOv1lWmFCPCBfpIJM4wG6DVQfNbiboWXJyWTVi6mhi
kiaYiVorFEm8wZt92yG7aFOn9NRlijjh3RoYJmq62i3J/BjlQD6Il4yHfWYO98+vxmIz5AW4MdvW
AtlaUSWtBDnWYEFhfAMZ6KLoCANIrIOQpmF+MYncIivCGzA/dYrQR+g/71PBRHTClpAAJA+c5GM/
ytd1OZMH6rRvf7AV1xLUOcTagRwiZKNJ1okSq/5jQq/74tTwaqaEpQ2PC/KGkSoX4aT36+CViQgg
tM33ZodLU4269jZRR4Hl/14My0g7o41mjsTn22qO1DzJ40ECf7eVQjcaLc4j9LjkhE3m77FDuORS
k9ebf54OqAutQyS/8uhaZFkQbLJxnjFqIJANOMs9dFwAH5g/tXNs9nk8Z54KrnCwuF5904dKEfPq
HJldKw9eqXsFe/m4NCUTciPCS8AAeqk1r3g15HtVvkiHg5gR/hfsvE8pR8ELkPrfqAczBxf+8Rtw
EE8EOLPFzBTwJVpO4urMhxnHQgBL0b3UVZEdXVaBbb1KuLCyrhkd5oWkjdoFx/jULIIOn+KQOqbq
TMqZcbct5gd9uK3Gy80OME0tU3e1pUdUorxsQgK0vKlVhvHhwlJYh8AXQ8xe3rdO+oXu89uL9MSB
05NIKFe5CWeuG3MWpz+f6CJMyucBD73kBPpU0c3r3dKgyzsE5iR7i+RlBktrAEU6zGiY8z/FzLZo
bRMwEA4IM504d+7zXFawHMsGnDc1tzPHNETPpBIRllA9PWI1Xeh3cD13J1J+ON2J4czfbRFEzd8t
P8+pQE80VYKehFourHBbND4Tb1iqlWHZrgleunipaqy+w8QCmFKKFwkAUalw5OU+yrCndY348bUD
0gphJTxY0VOlohJ3Il7cz/4dCvRzBalywxyeoOLar5HSarZgeOosa6bql63c4kp+GpCA0ZAQkfaD
51ezSa5lsNySJT2bxUdktOb/Zhk3szBH2JRSxIjIPBeHdkRBRVqjJwX6g5Bawqp2anGCeDWi977d
BJWsvLVDY+q4SfpeiPRPDIv5N+cMStKSVlkhXBOC3Sbt3xzhayx+0y9yQT2FfSAzv+1UXE43b0H2
f9+waZNlWVykMzE+50Jg2kSis/s6xdqeULE6MoHZXZbTZuk54aju/Rg3qWyYvcjBj60e205o5nIl
F6o411NitCyUOwN2PN7xhxExaKbGXHr5H7qErGJVhhOSdRUV4i6DUrqW35mxirB4Bf90T0SXL1Q+
bTYRsZOM2i3VF7Z8cNYXUUW7l+4VfrUy5BRoaSw15zDIfj+QSJXLvJLaVIlYwEmzrlf5RQjbiLtW
vA3mLNsW4EZINsmYFAgmR7kJmBiK3tJgT/NTHtyT6pLGt44kvWTAaxJi5xl1jxTPn3EVR2veBf1p
tOm+OftdnwSue9gZIyYu3FyCXnMewzDFprmCmidShiAM3cb0Isf41I63WNb8mAQAKIShCivNDAAe
dB8QceH42+k5f84fNIrfKaEKIaRbA/2yi7VnAV/UMvZ5uY0zs4aWFSl1yYDGbTv7PvuTfAuzvFQH
sVWv6WTxA/A9P/iN5ZUJHv1L9QjzUqGAszZOZNo3HnfDZoCGlBcdpCMRXubPpRZ6n4okB3RQFbl8
Uo6SeflsZ+n4C0V1b2VWGPJV3hPeGJtXJIv/qob6je6jyOjQBNPAl8KKqjOHhVb7SlPSKB+g3kLA
LMfKoh2ficUxHvXdzGfB1HI5w56oquAsND3hyrcItmhEFVEnTROdvRyP0J5CIQM/y48XDajpUDH9
j1KpLtXe1p9o4+RbCKLfpagNrdQ7JdI9tTe1+Rv+2Z2AXtH4ejJgizLfrg9n37BagpOYhibCLDzC
o0nEu2hm30dt9a6J3zyYrQkLNmt7ee5g9wvcnZjezz9kL3Lp36c4I/e8nkPohwW8oE1848ijrQ2v
jZgPIXa0t25vOaHH6HRPrwEQoZ0cD13ebkP+A43V+gNt9RhlByM/5A/K1Eyc9IqHLefZfBVWrFri
4TaMkhBv3mRzRerZo0Sk3DaT8rEsxo9dh3rOxIpttfL5Lkv2OniKGNVjjltIVqhL9Z0AoXvxsvAM
urukUF9o7Bl7iVY3+haRHzF3+zTBNAlndrj65SgM6+x5DCSmEQfSg1shgfBdZJZo9XwyF899gptq
y7780ZAGf5ObPjyp50jUzQELcH1YkuE2QJ6fNvdyagNi/tJ7GZl3Q/4q+VTrhZWSTN25FdY709la
qdqh36p9EnYGf6ZhP43ZvIjAazbN/lURljttLi1jNn7uUS5jA+CXIgo8iSc8QzqVsQqhuJPnzako
plM6xnJbiFv+2rM50Feve8TkP4tWjRBMf0mWso7GIjsL5INL3nHxiQ6MoxwChqUA8/pesbzf1KTQ
QzbsV5fEIkbf4h7zn10IbRS2oGumFCqjkWjWoxq6DAYOP7uXEiLKQ6+DdrQYNRyJRUG9UBfXHwdw
teq2gfeq8CeYGRFp8ocDGgSa3t+9rDzXZ9U2aGWwGWYuKaBGr2faROfXEYva8uhaFzFzW65Extd9
ZmQIRSIpHEmhelgMmZ5vtLG8WX168pWdBcEQqw2v/npxGwMNHUov3YgF0AadJJI0nHOBbsl7Uwo8
HgJ3GpJYbXk/BRPHA1F1+X+jnpVIludnJAuBFpduzytd0XbVeWt3MYW1KdOiIoMH9lBOlTM/tejl
VnbN6nueUBN5SXBY0iZUxtDuet376Y0AH2vCgv6qGGG0mUNDZ7K1X2j3d9ceyGJ5Ezq+M+O0CA9L
BhRM0W/euZfg80q65ap2xKbLSsTbuL0J8eov6IOWrqZmm0R8i2Q7WOLT8f2iGol12VwHOj0ZtXBQ
BouD+dZIree3bV+CKEp0pJ873Q93g02qNsJeKfrP/4jrenQY/VLAdU+jhkFq6axhcANli+z4KwTw
6FNMtTFtddiA+ayiE7s8M59zCSoKrbOYdpZqUg6OE/LsGMm142jY6Je3L4kS14JGfeAig6RbXrGS
vI+2SyVZ8o5PmNpPJGnG8yVycVKgaPsre9cGg1mBzBJzfQ9G+oYZ9aZmkqQXn3ZfGC4IFaj6iksL
e539DFyu0+wK46hKEVtOq+V5KH7iAGuPjxdUf6UHIoppZbuI5bvBoJKqJM6cMWqditmYcon6ndyF
/HF/pZZijF3CWkIQmsB13t21KAWW4EXt2gILNdZ/gO9ooxXFd4ompZqx/fT861g9PagJEsP3toHc
xSWaKoAga1OM82uUCcMqpMrYEQSthyryiOPVyZPJcGEEeh/a05YWrL6EmlmOC6lB4VGrgZRqiXUL
5rpaprkv5l7xJmN/2h4DAl/w6Q4IxNZLKOff6Jqwx2mQsHq0ax9UrVTn4p+yVStn3HLs3Iyqfu7Z
rQ3ifjwmNUvsgu5UhxRCTnH7KcH11FStri57zS807M5GplLjKvniocf1/0OBv5v4bNPc0X9UJ++G
7Ty2rMOPmx3y7aPi7psNlIJpplHh1YsB2jOYeytBGHthXluXSnMtsckxvheM6xS48I9/FpbkuxMK
jEw7ztKWs/CJtBAyozy0ueb06Is8L4978HQojs0fQgNQ8ppTH2gkTQaQZfi+2xpj9mM/N663uexw
PQEkSlaysBDadmTFKPTS3qf0WW+9RkZz3yI9ITLDTv4HianJLDeLHox/Q3DDMrR2SfmfWOj3xfna
DP0r0cnKHlCg40vI+FbbmOBpdYKWNvUfmOROx///zbUmjcEwQ+CAqx+ZytoV6McLV4IRKewvXqiB
8YDtqAVulGJ1PlLEaPolitgVtAG71PT7SooATpjHFxCpujnj2R7R5YdXFz6PeLsIDCpni7dfIDqY
mBSubSzRTQvx/wgZMUQs0yS2fe0uW1atJem+DMQAFR8FKANbr8YvzKUBIEmSI55Ope+FjzxZcb7H
oTXtVXNQr+bkbYbqcQE0NKUMYxCkFAJiSc+hneilzTDx0XgbOihFjBHMWsmgxQubsQ5MRynAG8cC
oJb3i1SFykLaOzO0Oee1HMFCx07Ze4asv2UTI1YCq0j/qNc98hw5aamU90L1MLzLWQ1N1PauXsRX
NA46rT5sW7h/p2u4E/KMyBmjC7nZjpjwDeEGk8hdShcv8FnSw7Jblz+o48c0OyZLR5grm8HMYN0F
bh8xw10bmV/08jzeLuPIVzSjgBp3RWp33xqLK4oQFPtKN/dzjCs8GC0e4Yr/5P9l8CR5pYW7g9Xh
V5wYdfddT5jMZZ2wmjyCZf0SXq4d7s0NPjQZXNa7ju/2CabvEsi4Oa5WEOGR6k1qoNzDX7x/HJbn
wjX1HPuLH3vqkStzxzTdj3JMxuydhOURwAl0Tnu2z/vwalf1TJdBQoca2fso+XYiq8agcYikKHFT
xQjgwklWqHETkpJN6jmVBkd6L5UG/U64edGQz/WnywHQakwQwPt4I14/+JToUbiUSK6WELH8RBJN
+QJnPtGO5c3WnJipE0m0q6LLDXMcSYXJXREeMt1tZGJoEzVp6K3ollTeRUKbMDZ0H6ALjghscdWc
0C9K+SZ64z63wNEYKeSRejBbXlVbrZUtaL0kMLWfWAL+3sQAsHUkgtaPWMdZCqsWWfyFtPM1Tk0C
/k6YtZP9EFIBCGy4YLLOrJwE0T/QyKjQz0rrpfBfg8BDTdFxngSl0JYt/7YdjkzaIYqTnH7eLxWh
LueR+OspoCxxnRKDFiQWT3lsYO7h2v+3XTu8YRKfpTVpZvkBb8U5+Yij7F7eknQZiLGNCNYafqqq
iLWTG77T/8WQnm0qcQvmKkL2kWd4kawgmUqk6hX645hvAu4jZ1xiFlRhLVr72mGtN9WkfsppnN27
Dojn2yfRcHOxjtNKdgMqj7cyW0xL/lSTWdKbMSDTlbcPIH9QcPmlfnsMJbTwGoaaSZMCos6onGmD
ZBW857IolMq6MHkbKbAn/iDkzLxiz2kzLxGUFhiTpktFdApbEP5Ful2y5snwLxV5tpnU2A6b4O/q
NqotiWqyfs/R8DLKz0l5TEaFAauI5Ss7sfaeEN38elD4zhkkwjGRwLgH39MvmJDG0p7OtuNUcM2A
RFnIMO9GpVvcykuRQvdNMeY7XJNNxpcck51iNRZjFmztge/0XnHIy/vJTlPBYKSoeWJh40RosKc6
Gyq/A86A6ioN8m1ZEQUTTPj0cE1E5SY1dSRkp44nuXGY73QYmF/DARs2wFQRYSRgHggp2mX5xMhs
JQ1vVm53SPhswV0OPhU7MrmQxicanp2DjBR8Iu9zH+R4Pk+pFn4ym+dl1G8nWkLdL/CkK8f/3IMl
ZhCdhzltIEaSzD6fShuUjqI+Q5WO/mr7aF9PU4yivCHfg6ZFj1frb8OITCu8+0yeUSW/xJyy0+ga
FGkPDavw+Mbc6ApoTQFKLz5L+IXpDCTKMnlc3lIFR5XLGFnAQJYS94rKqIyze574on5SOs+mjmdN
EsiGJIBBAFIAsAr76O7VpDswcqTGwzREUAFUdaq9KK84M8lrA6+b5M47xDl6Bp2QgSKyKa3Z8WAp
xs5dzYxyGjBnHgHj8FlKcP0VpTgQ/PRPzZy0fwREmP8cag2IH/aaiq0UBlse5MivBVfPfFfgV4gP
Pxb2hQSqLKnSl1r37dTxifz7VWg/yI7Z/xiC92tXwxS0mG1GHpzzrh76xNDqzVU4t6sOFjxbb5fF
GdgKoM/AUEOIsHJeDGKZF2T0BjQtLDyVOczP52J4DJvya9WqCijwMNUaOKdWgD9FyiLa5i//Yzos
nwhuRWL3dXruSXghE8szDxjyFlsMqEfm8rLp+KZ+Mq5MaAG21nKKch4mWRHSrlJT59oTlvpm9z4D
oeKTZGglMTldHdaFcGwx+wxaI7IqFzdAtCuvgWlg7S9DgA7Mrp5wlpdPB00sBMoFh2JGq1JkCwJY
+qAXG3UQNw886UdoMDiZwqWmL7gFyEcNTkprBu7CfJU9PALG7MSsIAl8Abt9mjBhYMseY8I27dqj
424WT/hS3+fCqD5du66NmKsiwkwdo9D+Kb+K80O0hjv+bcvsalHCWiTgJFXWqgS0jaDxC6ehlfIg
rKqSXbuczfb3N6LBkfKz/dPtP0RABLK9gWlAj4FR6xXXaVm+ovBQKUT7Eyik98yQsXv0BYeJI6Tq
CtxnRNSsyTlVPtTQkVhciwO2xZZLbQQhZ4HjcknN8bOJ/3zXzFASiwiyUlogUZKrJbmt6vtxY2b3
WvCtGfmqJFKBxOUJ0s4ImQ1Ouc5sT2G6hOErHBkSzKD8JPVHzUkeaLxWKOChXWKtpytNrL2/At8M
8cqBLjxIbhR28ehExx8G7zu/1XV/JfC2IFuTW76j1obfxZX8PyAiF1GoBJ5ciPhaC3T8NG3S9pcH
qEc6TSrY8868jIlGvve4UFx2kfMCZLxk6K34CNki1NlSm0jP5Esw+oj/o2WdOnol5/bNSO5Ilflt
wKPrBIJu2jYcLwaaIsntwaR8oJ2EjjSOl/w59jXi/Db62Nlt3eokkxMgJV6StRxG2HhpN2yZJMf0
nPXNfhVLVeMn8SHkwUfuo+1l0nXuKDmARdZHxrsz9wISADevmI/GcdM0IJUry6LX2xtlwoiiQzke
jdz64S+wiIG0czzzSu/O4FjTRLZshhyy6zjsx7xbrleK1HnMruV83b1YsaFL95cXbWgXxwcOBkgB
a/VlGNBdIgsw5oXG3JLcwDgqS7/WoB2XJwyp6As4yvnSVXdi0xISw6TbVHorjeFd60GNZD+Eeo0u
LpGEzZljFy75Mrt/C+RBmmvs27QeZwSKceHejJjJ+eW9pV+ESzFbGArWyqSfq8BQs3H8ySVtiily
jVsUNH7xzQsg9/8iw0GMi+h7TXFETVRl4JaSpnJQWBDavVRV+ysmPEwzzRuw8rP53a7qIbyTBWwP
TG9wAL+rp99Taiiqq9qNcdI7xmz+tiWxYX0CdSfoApzoJPt/+p8/yYblQ0BjfU8dZRPlG+GKW4M7
G5ir/6XeKByvVTgrZllekZg9VSkVjSL8RZifGNVyXbFXb4XZu0VFSkRCeERV6qKST89Xfg3JurKT
fqkPtJngoaWKiQBDjDXGSAw6qrxSpoxnTugcilfOO8K2445xf5E15KFLwc3pB3Q1bt3mPA3Ks97K
76N8kE9JgUo8GRrXoDgJ2BKXFzSRWDpwH92qRw1V7xBKg8nkfYpVJvOzz6Hmo8YuKHa09deLAGqr
rpV0Xcn+I3TyTTnHyiKqW5EnIuzgH5w3xy43II2GpRV6s9T9p+P7zZapW7ujlKAEsvtqw/m0BlG4
64/aPbfedC1IgefSA5CHkgJoaNHTYPqZd7FXgGmCSaCwN0XT/yGytPlDuzy26PPtrPCT2dEq2SJG
Wwieadpf5kvulTZLtU5w0TS7PJmOSthUgq+8/FrB7WcO4ldd4w65a29hKlV0/4S6K3kaRBCoImW1
NieulbUE44vOfJMx7n3lLIaKAqj/FqUuAeeN4QAcUHdneCZCuegdhRiWZ1BvQos/JY13zlQgiGDM
ztFmNEgqIiH7SxZYsRuvW4JQP7sg/0WKtvR4LveHKXO0zg3SvG2vaAXM5PmAUNGAOnpYpyYGx6oq
ovczfKgr/fC8zHVqKOdyDPaFQduNKuVcyEspjy7CHQXmar6q936A+t769CXFYdaTmJSx/QfaMuRO
3f/MO0VdHMU43tOV1bhKPXRQ/uIRBcVo1m7q/Vp6cXkXjhjL1rH6zCRGirB3tvzAJd3u95xW5Ftb
6oM3WDVI26rR70H4LIbvRVC8xFJC5o0PYRZrQ2LpWKQ6VmxFjIcNAXjQODks6a3LttYw2r1VWZHR
ERl5sZMMmum73RrtdwvgouLWg5825j5jdf9ZdatH3VklDCBw3V0P06GC0dK1HByEvkfYvFA5rmob
VGhI35Ne0SFtp0TWABJ2FU6DslkVQdCyIE+kYTFMaqtJcWr5Sq2OlYl2eyUh0W+ahKQaZSa7qPOx
fwws8irKr0wh1o+Q4SU1rPrWykYupPU7UbUaef9IDoWBvKb9NezbCTZWedfFAmHrtQzImRWiBsOy
MNkeGGWxVuDv+0ifPUEfbKMkSxLxVU9LDNSv8KFcd7lQ2GIWNzjVnriprqmi4M/VRacQJDurlSw3
/PMgqAnzSUrica3KuC6qdWRhkObi55uFX8r7aCSn3Bf36vUrs1Cwkf7/0Dhxo42uZv3mtG4DvRmL
7hQcdh/J9b1+/aghJypbokPjBIcGRSd5coe3Kj8vxsggt8c/x4DAv9e3/vQFNxwUR82S2x6UiKnB
g0MFyBBeal7ltigeBNdvarnQmKJVm1kLjcX9+6NHhtfvpk6Nxs4Bb/Lb8uLVMBTVUyIko4hTubSe
W4wWAJqdO6562avykjNUkLEEj3VFygc/17NctPehp/JztIzBJRk91C0UD8hx45I5JgD97TvaIBqb
/gWIQ8LHFMtE4rJ7x8TY5iS0+qS1S2Vh3Ded24KCUl+dBQOGJCvzkNGjj021nrj3/AxcnI5dR1ni
yhaZsHMs+I8P3mXiOBTShDAMIgnCKw8cOpo7eenTkZ5X2ioNeJR64Psp8Ua6kp9Lzg/CP4o9ivgg
1MivhQDF46tOMINPZJdwDrmuy7+CLYQv5d71TCdeuaJ3vcL0ZQY5MlRusAqIu+lbDcYMa52YMH2u
mX456+QVV+a3qkNfR9TtiSfLMSd6w2OpXhzlIX6Yt9/fsF/fKDaAzB2vG8oMTubd2bCNK7Z6ftpI
qd0K076YEWdUhzCtPoao654PqJCOGLDnJZhir6ytqcb3zOgz9Oh+AG16a4aX2yYzEIWnsO5FYMI/
1fwPPG2yKPu0+pB/nwtIj7+eg57UG+UPP8AIG+J7bFOPHsbt3ys9OQ141GQcon8cjpNWmCgyKrNF
CmZ6vMja0BgpBrYIs1gABcGjobosgrp5QRNB3kBJyYeBrD/4tjJVm85MVa8Ty2856fM99suOWDZB
VC61eYiHV3fPWOzQl9Dgp2Q6MnpZQnMbElzyfPMnrlAbR9zML3qzLNPyg555yddqnZ928b2Vuo3J
rb8ONFiHijpDIUbKStbUHtZIPG+zOj15AQwcCJJlwYGET6/tUDB1rl+WbdUagfI8LtTq4oDouX9F
727Yq3qwhQCpIVjKFQPkyt2vKpJC2yidY3aecKi79lNmQYdQDDdZMMqVY55466AoPmsRC0P6RO+w
1XsYziDtzU82BocDWijWgktg2XeRTeosXA/qrVwgNDUJEWWeL3XmSzmQ8oXi6N9kZW924BXX3hRx
wVbH1S93s7KSZWT7V4jW9UaBzpJgigpHTLrQ/kmXLhkEzeIqGZ0WUL8Wm7+HVtepmTPzLT0XlFd6
UDDCV/z8GcjtrH6Zi4SBh5CcbEPozUeXGNl8FVbj82hzlgoPsN+orTwlog6xHx3gZuYmfk8DkawK
I/IOiInACf06w3as44UIQhU3F9/FZoxxOkB2cLTDpLOxiktcXc5o1dJzO38gpZImZ9XP333FZG5/
7Klq7RwW1Q2cR0GblimDv7hl/d5cjqgpb4Mf5lBD4D4Budk6mA5cWjsUWAouqoxw5DpTQRIyoKPy
rtVE415HWYsiLCrP1giyT8X1n+QMrOGlJh3/tkILhuYozjpTAX7LaaRkV3zBMWWdKFl8NeeJOmsq
RKicD/VZOKz1RPpUf//37fdStCtWySwVcR7MmM+4PydjrlE1cQtqMXmmDW+um3UGCL/EpYea3uc2
WbeDzT84WpYxJ59nHQrkd7FLlPIZdSw/mNkFyMw98vWQ9Q32/o+wtEcfJjRhNY/B3ljIHBTZRPQ9
OjD2fZt30IPseSuFFvHOwBcZpFPvgbqM7RQ9+DqZ8KOZmN0n3bpizp2C6k0JECO6vPG85SDEGg5t
aSKS43H/zRXk74AclAyrYEVo+3RQOVMRuPLc6tM96k/WpxIXDiZx+EIGMiiTKQUwLIbaFs5WiirW
aVa4bPrpGdz0FS2cZX4HCcQ3GxHggKJM2ZLcbTwVeDaJqEeuUgq1U2JsCEt4MNNAGYCik58GMw+H
+Bh1zTsjzP0VGAczWv4Q+6QI3sepDkoxuk/hXW5pAH/8WMRwJOLyHle2mk/I51Ck51IZQmidentb
HnRPSVeWXKWmPiqlINjIv8RqHaIIxlOhrsWE0YAXfQJF8m1buKF0Wli6AZC5d3UTr81iUw6m8qWp
J4mFKC3dW4q1W9BbGzczyeWy2ROzczH+jwP6YRGgALWNPvXDq2DQJihUCDQve30ho2InF7CoNgBj
T6IdoCCLxCEUyO00+5ZoQFBZIuEcLbyNOdQ1J3KfGFKSGkJB/GRY9Wo/IHwPTTC/Dj/nfCR1CFPr
Lna1uFTDCPlv74aTGtTn6nKWyYzdHK4u35YTEAajQvqIERcDGCLsAzMt3ZkeQicfimsXUI+rOmvf
JZZKZz7qFzgbJKGiHLT/R0B0LgIW0yM8e8XE4i18Geeq6p4NPlCGa+iZdXLHNIDzz51Hp0ysmW+Z
pPV2Te3kR7lzmd6lwIavHBOENAZ60ohPlJK1eqydavXIFk6ZUQhou6KcwQ6nSlKWYXnhJ/MWxqd4
H9Vc8QwCK/HRPB+NCfXoQlRCvX/oTdTfiASba55vj3rLaLZBgj3s3gaboFamFdGhyv5eXeF8Lx/T
IrNspS1xM6/of8u0pnvW5qUwmO+LCJHwulz+bE/VOXddhC9yzM3bMQzmuv7foC85NGGNtH+TSZT6
3KdWSokxZtzhwHPgT19f3k+nVtTuwUljfoUMJ+PjfCF1PEu+O56r1C8MJZpDlHPZtw4rQ94GarCK
EAfJxLaxZuHXq7y1U2itpm8bos8kCqV0I6fDEFHxGlvrXGEQugzd4giiPMF/dhovWZmw8VI9RCuo
O4oyKfW7D6pEWUa5LkmybkiBjffy/Hov1Qk59eInpSvOa5mbBLdFo5rIveVKc8p3nM/efFwOcv+i
1cg7CXUJHGaLFJUvUYIoUJUs0GYYMVr94rya5UC66pu0G1384lu7/G1HnO63Q22y6ZfqQi3iMGFt
Y+m2tNwjq2fInXf+nHOnIsxhmxUga388O7zqNLgyS5WVhLy7bw0HtzVdCUXkMvmmnbASy9xbFzdw
lhgJPrvbFgwmLZSNMLJvRUqj/m00j4JaU+kOPshFJl5f9N/BwLUT9c85QQx3/KD9oO7UeMbYLLDg
2y1qNdMtaH07sWtm/r0S4jEmmiBIF9hqWxwerTatrNPm0jnb43Eukr+HqbmWjkih4qFd0xh/m0Qu
EvM1Ye7wQcOU4yIgk1NbyobY6VXmjqg2W8CSDoRf0hWstNjgefwpTqeDPe0IM1I4j14EJi82me8i
Qq21oP2RVV1d5mxOJxgxy/tQ7qxA09D4KoEvh4F0lgfDIip7ClB48SseIRJKYwbsq6EQJxiMR9/n
DuNXLs66tGvGsWwPe1FdaHPbIXzYlDK3h41FyTD2u6z4SgrXMioTUDSZvo3UCa62tGABT90akYJb
x2YcIXQfuECnYaIyj/1UUQP5PwtNGHRtSJoSlO/pupz27ouepfxI8GZH2pJNudd2mOCsTNDiUJHh
ihG1pzYiR/AbC4NmPpyNbkV6JOit1ixWqEzh9/oC2JonZxzbeR6dB6BWqh/ka6J70B3teKQi22BQ
Os9ZvTpIcHiXe7ABsQJi/EjgQOncnBmGVg8Z2KUFG0MKf0uHGcTpX8ltCtnS6/Y3UhOP4K0yAJKQ
CfOiz6KfOFG5I0soWUkmw+4a4xb7iXHSCCeSMf6/mryVimTO1ucCSZcET6wDYZCOz8+gvKYgLPDl
9HVLSw1jAI7bUYfNptlI8fUwOKf6l3Xn4MtkLbFW1GWRGyaCL1uYCQ+C6qgAfEdcvqXVkrXhshYP
zp47dKRYRHKetwSIyhKNJybocxa6hu+4Cr9t7EKzXwxdWvWtrgFQ49+WB3CvnJ/TbJS/o1iPsq1e
FI46NxGy8Gb8ciBk9OtjftRenMlz9vbMsL4Huoejs3/3M0PkRi3vnJ9jOWID95wY2c8kbIUH52kE
CzcY5E3fHEy2DVl+ocTe7G4E11ZzD17zlpDPhQB/FnSNddzUrZlqPdEol4bJZbLpM0hxhwqDiynC
ObpSxiK46PZgVo6aTxw6X/s3MT1VJMmAatOCzU8/QfGLTO/2y1L/NCwNAo5+PYpa8cpAd2Ovt2E1
WhvWWabbmoSG0440hJ2uja8dffiiqRC2WZMJU1RXnc7p9sIagn1f44ra0MJs2e8t0bx1JxHbde0i
LsOgt9zqgL7XqKIC5Tv/3ORfYTBJR9furUUP+4gXmbxuea2VY1dnHymI845Tk4SX2CT2N7ZK9I4i
sJTcNE/C/43bYtTZ+GvpmCRBwHxYdRGl9WGbKfEd4AIKzVKQhLqZ9BtaviaPjTIcNk/cv1s4NhZF
tevo7qgUavx1qp/BsHGsss1rhweOMFXayxVsVRA1WZ/hVufLbYDpi7JOm2uZ+7TbZEH7euyguYSZ
BKZ73mzAcZj5ccv3MMwi4TBKp5qohlL0dWxDdC4A2iuMcDSX+EQvYy/5pAJVQomXSQv2m0/W2Y7U
r3MWwF0+rXtHRlSfGC7hnGn5ZDU8VIy20Qgvkf+MgXMF0OgLD+kFFgiq7+8yHxsGkg7HD5hJoq20
u2SE+CvY0TIID4Fa7IT4rpFbPuTTkd48TRO74+WTf9BKGVI+HNpt0gQX4SCUAycJd4gVwWIvrS/X
ZJpX6kP0qxkzSJ7kalyrluFt9QTEg2l9UM7jNl95WtZ/5JOxTiwTJfgQlYY/UFSEKhJd0n6NSWOB
yMKiJSca3BY+4GIgs8l26w0hcCkbeJAVPg+Yu84Y4XnsLGO9P7eY/Vzn+istJvi+rlUkcME8o3E5
VslsW/KKbczGfHTTwy+KuULbMBdGqi1OCwR70/BMwmgxtwzTTz6xcVDzFE4LFs9UIqV6WOAO5x6a
pAV63IezcFO5AClY8gyAdqo4O4tm9gVKt6anm50kqOq6kDohODxU1/YNsXo1Sm0eJrlPoJNRj8Ck
JfUIwCRYDmg00tbgFYLSriYF0QAypWEeLknTUTSvtoSFs2GiBokuAniMYOIY+O0byj2yFNI16PZL
EM24pFYHYbuqXC8bxcrQnPp0qkdAuRlQeqQEFBDSJZbfISHvdLGtOIWJlE7aH9B1YfUPShjQ4sbg
6NXsSzXa42ZzJ05JhM31514iARLtndOsF0NMGyP/cX7Q3Pg9dgmo0iEL1EfkZDMCZODFzfW3I5LQ
5Js5gFWkNMQc3G4rHgiFx1jz+G3JpXoNE+nCUpXxLqpM/Emz5wdPuzs3SpVL8Nn1z7wBOHy3pdSo
8tMs4UuPtSIsAQyrhQMxpeFDGByNRI/gfHB8KGX4bETjvwfQvc99GVWzCsHnJpiE2fBRIAIiVR2c
FGA92B9N5tOrlCejKnAuL8kcbuvgd5HmXyHWiJa/xpbY3Yb4cmB5nPbgpgtGwrEXQpePRT2Eh4vE
EnozcIz7cUmDQAQsr3mYLbZMdSm3Wyy5/j5azcXTLfKG26Keo2yGszxT4/938SD7YtlTcibNkj+q
QU0A+YDmBLVTbCTZCIc1rJEIGj3pnHGdld9oeCFf2AlvANEAleBfPDxiEdghuXJCvxVb8BT6r2LI
+eeIaXix6g/59VAk07cdmK9khk8A6V+Frzg6dpF0BB0MdV6Mk3OLq0OrPKYPUHT4gNorYpsdwWlV
xPIRo0OXIghOMUAt84Arvh02ogms3ApTIN4RltIC5ytV3CE2w7iUDA+EmwlTQKqxRTt4Jg6U2SV0
vVL3ATdl0Fq0mLUKk7sufcRXQ12vpVbjxmarCK51z8YngeH1y68jHIrW8ELzk8POjZgpdJw7URnn
rabxoc1M8IM1dqD/L9SVtGYgroPcc+HthIO9O9NXswMuurHEJoB80SG8MVpIt1pchn9x9fEUu7ny
N1l+k+LMb5IiljZvckls8JQc+d8IXlgQ04xiVVtgI7Ypq0ZDGEa6jFSHHa/p7CB0rvhWhI4GVfsI
NZEIGw9x+RMScRIppG3eIoDW+sSXBKaFbEeIK/zjJxSFNCANsxzG5q19d1Hxho+D0+sFkZN1eha3
o9d+jStirrVt/ov6F44cligVFIMN0p7wbaJz1MbI+KexEBTzDAZHjdZJ2TkBWQU+qbMHQEvip1tm
1a4Qh/8JiPKviQnY3jcCdmkVDLZHnq6DuwQl85Dj+WUkmzi+cNDHMoz7H3KLv+wVw9D02vQHnYGX
UdDMka70gXaEfph3czx/ip5A7ay3/+rFY7rHKD+B4RjdTriME7T0QlPBKRWvuCtuZach7SZHtgOw
j7cdoTymeyFLluGtHbBbGaxBt6GMwRC/SXy9FxJENkcCT38hgNFH/ll21pIbSm4rc+HArH18WrzF
cZ8rpkxzaT1cgJ6qCNXsqUXmQ8m1SzoCBJPALS0piBL9upvNztQ+uFHpGgXnobtbYr7jutSbWprt
yubv2qZpeaE5Y8mKRHwjGQDgu36BM8MIGt5I6WRB8COzrJNLqAj8njn9qzPeWfQ4ZsJjfEqyxe/q
jF6DR6c9IZhG1UN1NkwJ0Ebf3lJm3SBppCV1Z9b0/GBhomENh3Mp8M9bk21XtMpVVqz/YKrFT9rM
cPy9/b07snQh1AUSAEsmVV/Fej6Or9tvPtjPJLBJyjYPTNY/hSvCsvPx4LOv+G4/HUIWSpmN4J8n
unELxaH2+Ya8FzobVFMlTYYL4JwJai8AngayZsWZ3riuesRgenZErH29PzpZwh8oviBzSjBrjl/j
98Ktlhd8srBJSHd6T7LijmPZgsnvbOZxGhCzKqMK4x6yUBir48T+io0gKswl9gy32i5J4MP0UQQJ
Z5L7s3zUly4v/9cYAHLXgdhrjhGnmeuQTpN1GBQl6kcRuHw1Ln2R82oECSvPBl2MlO4X5eB9f/j2
RvOjPi0GGEngN+nWbiWNo5vF8OzTbJW6msSL+7TbZacX60YqEvhnagI3LPruyS2kJqifWc+ulUqn
+1ofH9ffj191z6Sf6wBv5+IB1geAstw4IFRKOSewCIHDNKkJ9PRI+jzUC5RDbGg+dLshZmqc033R
uZzalrNN/OCErw9fXpAie8ZIrvPTWOWEz6pfufzN2e2sQIMoPZz4bdJe2ihcyg8PHPekT+kDCgiA
WxTqvjYPhHbn2gHswOhla6U4OBNKaUVpRsa5gzhP2sLSBkfVGBvF4//50yyzJLkcW9qyVgU8D76b
Op9zGm7X345l62tiQaV70B3IajSbrwGZzV4xYX5W8SeJYGSto2MQn/dJnBMrIrqlv8o/lJchzxme
kpc+duZLSwY7gLAp+cpuVmhmOlqbzwEEE7mB11TjgK+LC8+/Qle3IaDJfl4w17cJlhuVJ8tJwcxR
w8gqbWikOelytbQoIXwhykUoGUtYVVjvT+vdFzH2BrDkaszE5FJbitdbSTQqIYORzSHt4T3IymhE
EQMyKBpEIjd8N5Xgmic2g4CBuBcAoZCiSm6i67xH6x4AtOx+0PCuyh7B6qy6L16qOwirGIpO2nmf
uEMYNBD8DFyd61n3+Iyq/9Z7Wf3JGKVCo8x1FF3xQF7klyhQGIoSmU0Jr1N0K35NKlL+voC9le0j
o0tVl3iIv+6UZpeiuq33aplGK2ZmT76XE5tJSeIhIT2th1P0FWE8QqGS8V6zEfuDlLsXry37DZCs
yDrRByeUog7bEce7hjh0cVYt9Tfz+CKthhckBwEP5jD8bx4u+DS6g7yFwdtsO+BA7SvV80NWwStH
rfW+pANlaoP6yrEWNWDTw++4NUT3vvHWYsHD/3iTYN2TZI7L/yh1Z5Lan+hFQoMyRavG7efrZV4Z
0IjN3WqEfK+dghBKzh+LPlnBDoC0ryaZ/vCu3taWA+p+SzPRNTEwFfV1OQTcKkeXxje/3owOehLr
M+QXMRZ+mPxUQm40+ZD3QPZy3ntnf96iHtr0wXN6pjtfVKYDqjHrFX2nmeQBCGqBZmUBkgon865p
QT/oQ8ydM5PmesTzE4PDI3toBdvW49XrxyPUcm7X5OsZQJUTNYMHObrWkY3q+mgZ3A2N6Z4bvHYe
kcT0IjcG8Kec7quXo5cwmNatQLwVD73QE2Rr8sRId3Zbh3w29CgZ71zEg0yvkPwE0+OA7VsuoMSt
ldv97BgMMdwsnA4VqBhqMd+afjmi88xcZ4hdvJFsgbMzA23ctBzxHfP6DtIMJoTuzcjyayT/iVV1
VjLj/nMBTZumlbkoCAduCLn1j5SEIRHZprm3+n/8025HDIJgjFdncjJY00J8AN1bVH6aE2rYy+lK
Rp5Gstwb65tx+yssuzUNkCz6gO53In2B7gh92mKu0xiqJ1xDWPO1PdulspEuZyPokHj6cgfOIYEe
cM3tJOocnDY51SNKVDVVVGy16xqI8ZZb75r0FVnpngitIjBq0D2Y3Py0aXvmzlwzToCazlR+ggPU
jD8A0PDxGgNq+FCLzOpTSnr6B8GCKQqd5xnsD/0TyoQ2wkPoDdErKngaKEUcy3m1XoUcpYfiElXa
F0+cdgbqSijBHTo3IzVfYwC0NA6TmX+QoN1Srg2vPwQoy1CVqYWTDOc1q4ZjrsdRS1gpxy8IIi9u
7cJqEjZIXDDojYlCWycHE16+jAlkOvpmro+60ouv3XtAr0BcrODEuxxSAOxjvrd8LHFk9l1pfza0
rAkbJYcTAFIWdQcbjEXqYJv4Q/yGCkbMLZXCvLzytyHXmhJJUqE4Sa4Azrn/wXPrlQP8THeaXrYk
MGV8/mOfAXaOxs3omsWm2uO4WbPHPXNZRHyO5Pyg4C9VAtxCzI/548EjIiZaJC24EvVSdO8ioSjK
Gq0jHaVRrhMYGLKFPVG8DwzjSxcTPtZP7/8941VMtN5x7iZGG82R90DoPUnGVJlmSvs50iDU3wW4
68zvnNODoxNwXndXKMJKbQchkOcB5mwTUWvrENQYvY3PKLQRBy4u7CNiLKG2cOUZEzscRrkeomaV
UxdwT0lT2EUdmlfEJiNspTntzxoEAetH75jOM/OKF9cLey+MVQr/f/7C4nTRj43WUT2jmQCRQXWo
LQqlUvt05J3wzcnfRO+7iCm+uVtSpv40QfQi49Dcbexb+re4xo+x2WIgjoNm6tg3ouh43caIB2Ir
6/WBkJ0g+69jATUPW9igaOX9GqT4jzjY2wJ1gVttl0CfdtwJ3v1Cf2fahPYmNHo0gSRRRSOGHR1O
sV5zhBNyISM+kPygbgliDd9tGSut6DEFadYnEEnESpsFElNOGIY5418abYRsaI8xNMeJrK+zmEPr
BU4DfpJpWMe+cRGbQmgOzn4kw5qexz4GWx7k7oRRhJDOeQvtVoPOlsF3RiPFSYRkkXr3OaW0ABgI
lbbkW2XBtv43rxDV2rJ9cKvbxZBogqw2lVeP0ENEZxl1AJTI7TdN1LQrJ9RMT8z4X33wEjIwR3BP
dG8zDOKLrView6ok5nat59+HbWwY3WkhE4770C8M5/Q2rA6P7C/Dbj07JP7vuVw0mo7BhRXqHOAj
eqcXvXbN+SL1N2fPBXLzN7mZCE5cJf3vvzpZmOaIHkX0ESV+/JoSXc/fP4fK6GwpOjVeDgSE2WB6
yza8caYgMaIUVIRqu9qsOe0wOiAsZdhvgp4848VR+MXZCAnOL7dNS2zSkC4h0f40Y+jw5MEfcToW
OgHAe7h95h/ZjS3Xr5Vv6gA9r7K70zL2OHsJKGxTIJvmXsuG0AB/MRJloEiaNbKH8P188kJsVhJ0
bOA6xVmKEnAnaG7HbEzFfpTS4w+SStVLMlUDTrQuqZXSV8Xi6J+FQjvBzKU3+uNtH2Xf+MOqkaLS
8FIqf9Chj9jp57pkxVWcdyXoiUUG69rAGP33LwdFkswWrCwkwl7Ve/sEGH9mekEiJJgdsoF1hpX1
PNXMiej/y2V6uKC7r89DinBqRQWs6WI76juj1T5Hrmm+eZLkWxdkVlJHVET0HiEzJpLoLiwEIp3A
lkjW3FtKtlOtzUScqDvUkNVg2wkN9muit8oE1tgL8tVinwnUWSLhl9ctSf1P6mHegtS6encOllMD
1cHpkmefvFpuSxi+js2pFjJrmpxf7DbRngSmBf4wk8M+h94vFou9icj8JvX6lACX5uICXkwlb2KG
H2NK7mHkJ/Ru3XsFeWlcYGfUD0Zfcqmcvi9gdSi4ChLBSK1ygrGZi1V2eUbAFcGWD9BhCoa4gZ/I
TvV1N9tD0rzwkk2fYfqOJUaFX0UREWl4sL5CbK7WrK1d02SYMKSm0Vcx+zT8EZFtmEd6Oj3+Wsz3
v5yt+A/VRlEYwY+lWSoqEeiiupHqvxlVO2eFl+ocyFWm3TIpW3tDI1Q2zFFaxW/gc37ZGAkyEx/A
fxkJ8vMQUbvr22F3R19YPo1DReAoWvPvsFuEBTNklu7fUSAVT27En5AWHALpC5xJ8G/QMfGSyd+L
6L5YcPrHvEhhbIq15mmo9FyGvdEZeP4IzewJSDTjLh+gDON8xm/q0vfnAyeLe91BgNLal2WbdHyE
PSF0mTxVGJ0SJmi3y0eShmtAN6c/rMUiU/Ku7NCLJWJlCy2N6pGThOdJsOcObyI2q3WB71wLC/bQ
mkzyoezZsHvtjcwtFwAy3fiC3zabdhZUMJegOEjjREIGFVH4Vtxc8azwHiLHxC9WclUlOy2lVYql
VpPu2b3qY3NrwL/Z+kRvGBrdj/KjWFTKpje7XX9wOzIxHlbvMuiPMP50M3/gzaa+E8O4m5mdGPC7
eubAWR3J7uMLp2+yvAfQUKol7N2tJjb8Jar4bKYaa2IFHZPxQU94f24bV8U+Gdc2riQpXj2AfFhB
7A9ONNjTqpH/toLxvQZs0xoId7rOmDWr0xy5gDpaMuQS9JwBgmE3delS26rrfJX6VyzCEUpQG7CW
z9E5N8bIur3ax/dPPHqcShtX7sxcAetVrvK/J9+Jxy1X4VdZlWosgcVQi3e39QlmGKKyJqaG3Y1m
MH76QkV8AxBOUdw6cKcGYcs3hF36ZWdhCFE257ckgdGSxIbKTyi5ZRUAmUqpQ/WaMiS6wStJmtI8
YGdj922V90DxcsKkDn+KL9+UJErUpzMmlsQq79aJ25Mf7eGXxrnQoS6lXgUTK4vuOiWz5U1czCtq
tCmOrSaJP2oQ6n+18mmF6Zw2znWXVUQSf1VTa95Dx2E/98PBBc3exNucbrblYA3+aZbW9SUSFXeN
Pamy0SWnsofB9HCX+cpwbYkAcDTCAUmMkKYmShQKYasAsJQLmOvrfTHfyGr1Ham6HQfb63LwkCEs
LLn0nSZl13pVT6+uq6La2dzE/tCJF3zTTWkaAkqsDED7Mpvxc/ukLcimqdjp0nOetHuZegDnVx3j
d2kxvbjkRI/5OdqN1zEZSvWWiD9LfNR0G82KSRGN04hu9vEOf47L64NweypiAnA7LWp3yv1SB1Ft
18gms6O/SEfUR1G1zs1RrbhNh8YF/NcrqyS/frYZoOX/EafvZvj50jJ4I01L8FgTaW890Ce48pAn
qmGY6I4Kr1+wlT/Ig3tlMHzi71x/wzYfKu8wErIwRutX7Gyxdu68pb6n3uopRcJPk8JwA/z9QnnC
L6Os59YpGC6doUpVNogoKvne+GBwmgnmwXJZL9Xu4mhi6XIwtjuYu0MiKPlQGriCX53M6FRD/ZQu
lVqTj0L50iPqhYtgzeaJL4jhqIgJiNC478UUqcsHtHJ85ZpRee+VBZHemAaT5+scKdn3e6gRxQgc
+Mbf4ynJ32T4WzNQRR3STG5zpTkAG4SMPDE3ZWoWtiWiAeULBEF6zRpPshw9U3K0Q26l321zMGma
cRUbOYK+/mXbf4ra5Dpb4RtvBXpFDp6nKSasbjqFMZkx6ycnS2ON6Tv1yoF4EoTrCDC4aehVXi5b
enKodngGrN1R9PZ1TuFYSjeIY8Ua0a+EyO9sFGVYiwWMVbNuR6+Ycg4+LsddDlziBUpjMdFhQaEA
hlrIhUptNDoM7lv68SXFYwrldAqcGH2zWq5s8/cE6fLwGhAo9Z6y+d/5M2GIr1gRlGT3CUoowYz8
Sea7o/q112KgN3hfxCs1xBu7Klr9pE6ojw5VaxZk5gaXDttaE18LvxKPLxPDkc0UuRu/lg8Mk82q
qBVVyiiC0kHvB4me9E6Z8L31rscIhopfivsmuV2od7L2oXk4gWnRr3scYFvgW2QRqWyRMCig9vhW
whx+fs8losHIqG7cRJtrBiHfvODzzPUXQ6e5zS3luOYBBijsI+V0WLV8pLVwvafBaKxx9s8pKrGk
71qPDfukF41NaGMqE2jSsRRZaehCwfEW/0fJqCFSqB5sKcrfXCIKG1hWwVoMupFSZ80kCesh2pIh
yEYiBABwDYehiJEJp0iGmlO2RPAfXS/ykTNh5cek+1+9MG2SA9pg7edi4pKhWJ3nWPmCxrjmMnOt
9q5F1AE7jAEFLuXysDOTR3b5H4jKT+COOekWHQcE2qG79xV3xDeWb0VKlvTogCu/gN7hY9w1okT6
PTw9PY3rGFUrvkj0bFr2r82WT+T3WKGwlzaKxkcr4nLP6FvMP6ErrLp8L9PoIe3Jfom6QQ2CuDcc
th9IVkwPwV7AwUhqtIUFdKfGr0IfJ+dc3hFKf47LukLJqATLkPB8ZTnRJe1DLoASqnLNntqw+if2
RNOXEktZSviUXr+CE60mIMjVCWWud90fad4GXqo3ZyjHPnQ86o6Chmi8wlKvJtE3h7UkUD5dO5CK
mI6fiBcSU61nh4gciyAsDQeL7oI7D9dKeXMhphAfKLK5RwIFh3PZratBhD8f3Cf64UKgjrK49/uE
Tag083YGObwyF1hV+7VB4dGqlUnl2DjF/AnLb6M8R5xAZhw1C2DbEsRN6f8O0okEhBN2Y8tjy9BG
wFGmb1uZzRSWwRmzohirpjWHWtgnCP3IatlvOqiWzxemtF4gaaBTNueoZJobaJoVDXuXcEZy13Dq
ehoPcYbDMtSg3KucLhDixfT3/knveVZmftW2JPGvw1/d/05nktTiCwDwWtU9X29/7P6MEfCNPLch
XUsuenmusE44RlnW2v0C2UMJan6oxiFfMf0Kdsw71oL2JGG6OP2oUxScDUW4nSsCPQrT/E+S2AtD
zXqq7XRJ1tYpk5DIvo8Dz0V6335EKUHS/cf4Il1Mj81EaC84OMdhJt7fF5qQSFtthW6KFY6X343P
ae07pQw0VhOBBn+2mcqSNjVW8cdAiDoO5puJzvb2F2lbn/KWr1qbva1hcoeqf8BzpEAS1BlcyjeW
QuMGjjmksmtITHnvrhkwqO6dobXgxh6SledVSOJS7m3KhZ16AQGhRvqBu4F/BjzmWUYXojPRsYo+
4n9cbYEkjtFcY50fuTTyNcbLuy41RmYaZUMrXrs2PS4XxnKIG9Yt4+Iv+p03oD5JRcPcGEcCqjj0
BriL/B8iCNWELdxCotd2L7Lz65KNFVkuN5/BgoH7u5tPY/+SdYzMxMyqGG/Frs1ZYelpDnzp6/1/
W5eBeBplMu29a+DovDh8BOzBJu7Y9qG7vGH8Y0unoDcCAT7iM3simidSBbtG4KUZAMd3HcYo8DlV
16KzeLVA2rGzlRnfqPTeawmPUOfXQI6X/tnNX40GNKZMxosYPMF3IMk7NfX1wyBOD3GjiHAGTt1E
nU1cLqRRtW1yRlc+eHrrURMY8c5PVNk/ZsEpVuPd3gjRLecA8XxDXM+BhP5C+ktwBonVaQ7AltgD
gXbfPZurgnuHAlZXCj5vRvbravWcxgdorazbCrbMZFR9W1WfhgalmR1PN0uBZZ6pkrAqKk/o0UN5
HmgiOB/34c+9qXdFl4Xtgpil01sS6VZ45TZt72z0JHpNsRHBxgAwavUb6pxQHl7ajCqrg+Nqspil
JIgvIGITB0NW7I4pbmCw+jMNmxupgsa3nKnepmMOinkZsRlL/D90zdqC8l576NVvhhU29kXwThcx
g4leKiL1FGP7BXbHpsMoxpURw0cYh1bdkfYwwTf9TwYwC6FBop4ShLjEL+F4XguyqfIIcOHrYZ8N
vFKNsHIyTGOUcnGdQN6GhE7Qd5cMh/gKS4snUGlugibmVCVXP0KJNv6iFV6Aw/7zy2JSx70wkitN
jkImImcwC5wzrx3vV3pd9ZZl/xoT5IRzpM4qaXJkD3DpwsC0lUYMx8COhKtJkyA1IucjWfRzCwGj
82+bebf1+nmOibDWnnRHDTaEp9AMucGw/KItEO4wxs83PWEt+KTqWHjUywgz7jx0oRCmB7k9HRJn
B1Z9WFYn3+82mq0sk5xqfj62KnQVaC9JdWSpZXTPZUR70v5a1ja3YO/KKZBwRZWEp2vybRiHibe5
RSZGS6UJzO+/rjnb37clABxd9wkx1Jb8qvguNXJvKFmcDLP6bLQSfky7KVQ/1K+WAH710UvDn6K6
8vR8fm6eAOWHlPC5bNbHDicqTu9D6K0EZ5gxo8fyNwuYYicvsq9gVcVnKiDwG7ZQmuQUO35SXHCT
da12w9gzP5mvxcJOI+I/gJWJ1h3JJKx+SecEJwayFEWacQS5Dntwp1ocVBxgdLV7Go8DF4iVhCHa
XY/XD92PbwShF7KSQwolGuLEdCJ1YUzhSkHz3m5tHjWCdjmErMHTrUDd6b/wnqV6H5e0cHrqXEXy
bE94K5IL9V4+VmIS5wNlBSf/jzSDktsVUg45hYLmo6pnpscPYFyjz+Zbea7lVRZujUSrgdex1ZFb
NtD2f8bJAFbsglkmhIVAnYmMzT0zsN2Ty2lJRraGDccbEmMwbw60mdjttRz4461j/Vm9IvBmuzvY
VwiRym2DJiDMf15k2wnZtx/3xh+ViUGQK90eIldypHlaIO1mfg3F2rprGxSgl2t1qwTYsOShG26S
O1BoSWd2cVum7p87Ep5hbXqXt1soMvEAmAKFe18wXoF3sbmux3JqXjKfgILLdc16iU4+/HfvkUiB
dAUtjyb1gG4yFlXtKwsWZQyoSX/DJ7RyMeK9I5LYSpP5nsTiaIifpMvHVuTyEuV0CrrAflNiSbod
rUtyl1XC1j28bdiL4N7z7VC+qTXOTr2qSOLNvyI4im8Bf2RgSZFZ+R1W6u30tUtSUkqH2B1oCxYK
jug3JNbofZOxY864ZTRrwJCuMqG2yE0lTNbBS6k6sfNxfB9nNcNHcFwsC7Jwyt6udapuwUg4VKMl
khpNZYS0p5ilztAgrRgE3AIew/Wg6jUacY2Z8fPw71Qe5wzGHdDvHgv2AVCUYtNnjAl9bEhQt0ZC
0e64th445VNJnYWFyhmQn0RaP1Ucs337vQaDBISgkrGDyCtHon2YomnCSc72Jn4Yn+kPidfVWut7
E0QWD8qXMto5edhXU/+prEtsmciLz7wispAwIvW3TgUarNBlosr2T0cvadkkAf+VOGmlZb52vESK
7oLEt7p61js6kNp6zfDgiIGIFpt+oba+jUmqobps3wnUeYZJkmygS0yI7vnjkDUsOhEgXIKVOkbD
rzsvNzP5Wvd11lRqMTpKdzr3HBmxPJ/dQWzGV0xm6UzP3wQ2uz8zYEeQHwxRaXFyfaW+V9yfypiv
qSjrMxh4hM8xAA6vDnZOtYTDFuhEkizq+RAYOOc2Sw/zweGOZdxa5PHaRfHDaAjy2wgOR02DZTR6
q0Zklja8sMNgxBN84ENXJ2F1qhdriccOvdSHjb6a7lngoiA3VHohtOuIeddl0g6xkvcrHyj62J3i
Nfp9ugJQqdUloJE7HxpnJqcHvawbuP4d8VIn7ZexkCG+UOW4wTVWVEQt9gOVckl4P3Ftq8RL5KXz
lvcKjTD7kZNz76phye/xevECD2B8zut0SDrQzwasIFGOAjkyXYwTaXje8Az4YX2zigb2nsyuZLUA
8ZqF+YJSYfWqeEJdn0WBolPfqffpk6sKUspNTL2tq7BN9WJjHWjEyYInVxKc4vwyY1xOguHJOMUm
BsXNUyLO4uTSZJzHQZcZGMyJ8SPP7qWMnYzaZ3de0EDYQMM7TCEsbUoRDkCJymjAp+Yv9NLA6ySQ
A7WNBWH/PHkJKCwwYYxT//XQccOWtNCtj/e1xpsG+Zm4pXn+8JkqMpBr7hrJBI5T7+mFuGaqm5FA
il3NzV/y0m/PWcm6XXenbczZtotgl8ra0dTxHa7+bssxBlgMcSVkiHAOn3jQiwMyN2CM3ubzQ5Js
1mwLgPHFZCtFMqCR8jMPbrIENwKwj9MRYPMzc0ARFiraF/Jcf5OdoBI2ByLjIfydJPoKm1tFCZEx
+jM6tfutfJhrvobcsD4gflLAzKjwIO3kVD1/Up3hwyTKcIMnX7PkQBGUJkCDTPCUx3Vq8QDVz52l
XIe32uvob9a44spKBLRffVZwdcCMViJsutPvTx6cm5DSAEUmg1iUSfgdTjHgkudEhuPi6TqG8GDc
01q8/sw1rpSyVgHhyLh0pzNKmoAoJx6COIXgFX1FtoHKwAwO8B/8x68VfUXpnlAOyZapKBQEKavw
AGj3FlxgeBmGpahLcUReNpVg2hrk45LCp7WVVRS8UmCFRGMAU74bDnCoZKljJ+FgJbqoV8ZZg2GN
zPBwplojtjhA3c3cU5T2VG5rjZ2tJMOA5Z8f3m1J3qKMcfnPzgCFtxxD4OaVF88svxHLTOAaRG2M
/E4q/IWxKNzlaOXZgS39Zc5DYIa8pQrnE+bOlNLrHZSDxIRktdBybUQQfbDfsrjkr3HsyebNnKb/
gAZ+vzqnkCb4xd006Ovayqe93VutUbiYOMxDPp+c04bNApyOeHnJTEW58irGvZSO7f7sBr0lu27i
PzyUyECyI/P/TFeDybIACmJroSwnTvHiUjtRtobyXCTyU/6UjLZL7qb0TKa+tulCa2jkv6SkGsxm
jhV9nupZl0/O24s90CmP4e+dIqMVSLVJXocM9SacrobBJ1zQTxAOKkEcGzsGVoQ6Vx+gDXUO8J2o
R8PT3Eyzdhsl6iyXV5CZ5NvFD+tYyXppw766vEhK3j/VUJT+AmnEe+p3G7rXVB+fAfU2C+GFfkAR
R9z25SZlXSvDcDlrnFlzw50aQtCbbaYo502dYrqEDZTwaKXaQ4ZFWeXTlNhbzeQTO2ZJryU5Rs8C
u2NWe4wRjCkdTYAJf31fCmBcr2zAw5bodvb1n0Zp1vs5FcYeHKE1eDfPcCMPpzdtNeRGnLrvZYzQ
yHeEfiOJTcOzceeKLP5+beOF7J04KLVhys8VNLIEBDk5Eep+UzDwGb4uU4B5hfF28MyjvNRoNfkD
qfEquXPixw3bGmSeLCuUz2vKlVHmMoulups8nJZ++EjsfwgVGTgV1mJoMN8wKADx/YWmgC5mkZqw
zhsBH7X47d6SjJeo13PRIa73yE3I8j+Zt2UZ/QXZll4Na9amz18ZXitZFhYMq1oYu0/RyKia17uN
GhRU49+uUzHMTiagwrzB8llieAiBl6WGc/FsBXvhgvAnX+X2UMLmCmh6y3QdPCwDQA1q7wwZYBKq
dZs4n+Op6CNTVCNgSGVWwgh8Equ0E6ETqENMSiJ2UZ7LKsyKuFB4IoD1kSoSwY88/48LNfDSkyoy
S/B3dOb/8aPc1n7A7gokOu/Le7a3ECeVtZueSEIBXuAfolyGQ13887E+Cm5Wiq2j61XDKTID59DS
Gx1eMWtm35Mbiwtq/49GnZEEG/aR3uiZxNvyBDDQGcvKaH+eR8aFsowMkEg8NZ1aBoL/nze0U9ei
Ur536aCxb+YXzqC7QC4QmBoDzRO18jrV627DQ2qAHxzd8ydJ6BDDVtKxJ6osFA+H5o/W2cN36qPx
S89BGBmErB1vFDwXU3eBR5mpDoiHCn8VgZIgEPO2peBzPaIOMlEEH5N53vRf1fS26O3M7h8w+NN/
ngRAGMi/V6RD36tjuY37DTVktKORRX6Y8pZlm+Xkc8JIOteZlb6LF6T3u2hGGqkfPQhxMTG5L2pL
pZD4Pykjv9NhFsllb9xgT8wWI2tp8jb2ifhPap/3lqqdShLVQIS7/3DyzMdK47XEXIZYdF2scKFo
c6xDWLWpKw2DWHxB9QtG2aEm029PVel+kaDmTg06ZFBBzaEVALpX5AnTuTWi4SVDbTNgzOcg37RZ
LNZK3rgq+rpeHyD6uGY7nNy75bMwccm5tgd76/o9Pep+rV7tHwdFiosU8Ngrce6HYR2F1MU+rGAS
6A+qMANAUSM66+rOYM7tYc3PFikTR7vb4n2UQFvp1h9jW2M/pwOJqaGGXI+qje6hZB3J1DQZ8HmK
xn6JWbUZYgh8Ff+oHCFabWPiSZQZDbnIYiQ3GsTbXC6TN9BsOYbguK7sKVta6LjrI8VhIWWlVIY+
paTdqrj6aurMVNRNQ2cc6UGWn5fChZcqf6V/ibmm+QZFHjqPMWhOzoiRW1HZuXk6WlVka6ssYlpY
vzn91MwxjPDLJ095YVWxff70yWqrw0n50jLZYiWapDyni8lLT1ryBm/aRKkBQK0Gkq1Yz6KsyW2A
eXTjNipVtLTX8ekVelWtIKIF+S/1oOdHHrTNuiGL6j9fW5cVIQHK6h+qH+XOtdHvzxeLmZSmRewm
+2J4OmE0c9jXkjjPPr/WjfX+Ia/5FjRkJjlH4PiyDPoGctg8ABQQ3rKCAWRUzQqcOEP5iinKWxWG
cpRbLSPIr1eGIk31QYz85j52gRQQSk1q0eClv/ab/6pCGoy+LzZ0EKdvbJL+6AFssRu96CD4pJhH
rbXl3+qPHZdwF6vU6XQ3FFyAqWZHUvT2rpnfwYtwSdT0imFKo0c8Vi7VCqKny5drEdHcZg3cGlgQ
nkYJI/IFoypmkqgHVicHhFtHmzu0pbH5b+1vNb+X+vlwHHFFYZlyme8lBou+2+qBCKyoe4LwjOEw
MA0BFc3FFBqJ/fTjd/W3CHRcymfWHpk47y12um5ber20vjtz1uf8rJX41uUR4JtQvv36DDdceok6
ZwElibFnIWwunEdXGpNUUVk2klDXTlVY75R13URFbHINSp2pYxiTRxSS/NIZeRC+s9B2eEYgZcwb
PKxA/7iOMu3HxsWOJqAjVesymllPhZdpdzfnxGUMJygAvfmtNE11lhs19wLa3Xeyv+Fur25aY8Gp
cGYhjCLnQoX6Oar9DF7LTTkHscA8/j2DEnMEHjhj9YdAZ+3NOaXgOqgfexk9USJLEEGx4m6htuTV
3wN0B96ds4Ut0FeL32pgSRLui0QLJ7R+UbDuhaGbLdzC7n+bW9sXi1XPvxeHDYM4J+k2HZDRu0sE
ydLXoYRuxAcEUak07BwbkW/RnChn1MyWkmSwwBTn4RsFbGLq01NPizzK95mBJgLXWC5StNgu2+zz
KVxe1ad8IZwQhdo+IwGwpFIQBT4A7rgXkIkSIcS+cYDcL7ETPLa0EQD3m+XM8Q2u216g6CLgC2oz
5Oa8zKI8CQPqSD6ynZwTcTct5A8mgwjtAzbCFRksFaFxtrkuJOFr5JV/hGGZQAEyNimQ7Bl6Y6eh
KNgwn2zeXJimZWB+1gBYoCI3NBVwNsoIM8eIITzlVkyztubsN9ozqlWG5tDd8y26+IWRfjmkyXDg
sX0Yik0cdIKQIuiWdrSsoKPZNJYv2WIIOMXNNa9QrmdsHX+a9OiolIypTLBknZxRSpBMJVO+4W2u
LNJ3V2IVpW2nklSXxbQxgnnptml7mf0YhfaCJsrrNFshDo+poMAa3lDWseC7QkDN267yrqhJhnTN
WApbYCejSrVY7UEU68vybMobZDEJW6dN4+1wzrAz7qt9oJD0keT+/GpHzBH3VXJMFQbykK8QZ6E+
RZuu86g/MD1lSZXycVNpZstjhyJF1vB0VaLwIuFDt4FmQPks8LU3McfdlHkgxM9BmWY3F5eQDnBF
yq1XZ4kGicIgN3tzj7rqwrofTtLsU7HIk+6mOgNyk4WN5zOO4DT0yGQfLCEjwy5hdUvrCdsxErvv
3KmyX9tjrmbApaYGozFWAlFFafw/2UDDFI0yIKfvSH5dpmq6hCpZ4l7UFzkj3iSr7ms3nqOkliMH
fuxRX6OaieAPnOPiasCehbQnaZBOTZntpeVCsB8WqANL0NNuRlCZNgLNlpP7tKdaJZDnQZe+KN/Y
Re4iKRr0VZeRYQh/KwLbuH0UZuWHa+CP+tE6Z7D36DVNpbKXYbQUYMOVuWqAVM/xuO9tam9oi0kW
RHeERIUoiny3P3rRebd4SAsoJ07Y5X0Vw0i/b7ZkSneC/LesSDjlUH2TX1gdosgRxlhY0stzlyCM
zG1UwW+60/ABNda2RTvYXn+UzIbK4HWk8yd8EOCgSrXlXdWMAIK8b7pLJxtpp+dMtvan2zmGAIhr
ipPnAWnMuAnBduuf4FKRr+jsl1HA2cG0sM3Tv6TVcCiMOqdPf3M6Ycpovy7HeJN8QR/KRFk9mWUM
vQIz1rYnFFQDe67b+2BB1+qukD2CWbwKHubuyU9yMJankSqlVLDEMmf0LicIzXXp9FsgTPJC8EWD
8+jhusWCO1FaKE0/kkM61SvLFtqONjADwhVzabG5SzkcYjhNByVpFtEzJ/FeVP1szcC0ypUDN/Bv
YuPekBfxcDiaHk553F2ku1jYu5oz01xclTWswaJyCufxB3qg3zA5PbXXBOWFXSJuH3pcBVpYMfon
qdQbWvsYpbrgsJgKEprvVQY25dtuTZ60y0dKvSb+hrOSuPb7dyppKSk2HUru31ZMRZi9WE7d7UGX
gBURf/i5PX5yZmQDlTqfLV+dWLgn/jpzrvxaKymVdfOmG5Gi4fZHPOWBgo6zk2NoLXwQJAJWcAge
1SBZwOo1MVIspmCFPhXaR1B0yivaD4FJ+fPuSanJWESZPQxetQeGOh3BUePRPGprTy3sGCMk56b8
8NENfZ8mzexPtsucchLhK4OpS4yRC6xEbuFWyyjO6QYD/tJzD9/e/UG28xsrMwHQx9TR2KQOHLce
KaPwd3YqE6wu2zBl0S5b29/eZTETXrnAzidXQm9+fXnfWtpHvKkPneuqVc+VAPG2Z1u70GKmYkvM
v8zhPLOT2v9/9aNbDfF6jn/WhbzNLM6Ck28KRyN2hRK8HafDmgeePFy5Pii+nfYwNH8b3AYSIH3c
EPB6fihZmiWLHoUMO3s4c3fzBJwOaUuOrQfu2zRW3MPe78rSgKgK5tfpuBFJ7ZoHBQkzQ2LYCiHK
XlfVQkC87vEL86Y0I++ybS2tn7KyIguG5VPbPCWz55IT/0sEQcqvMHcAunTMdAxV4jMZlyaM5r5j
t61XHb8ZHK9ppUMxtgwm4E7iWgArqph5EkEGpjhmwdHuweiI8/ojTOrKFvVCF2VJrtj9zHVVRtYg
Kq705qv/ri50wY8VAc+LelzoVQ26F9zjg2Nfksq4lh/Sw4P+jde8a5iyUGSHh+nUhaaotYyGRntf
zvb97dnkhOa4/KfagAQuZPiZbgoFOBaNJXabJE74EH8w2z08o1vwUmGvY7Ugm0ShltWJYRCnayy3
eudPf/Ho1fF8URZ0fc/pP+XzK8NvnhfsEJ7zr6n4mVWQQ7+kbSqyGkgHQnEedL9C/1xuVf/A5RkW
kzJZAx9HkSE/JS/KF8M1HlLdx4HwIU0KorkKkMezztrjZZknc6vYJXxHelzEhadt6qzZJ94zbheB
nzdSVU8ZyGE2FWkBhvT+Qvia7qdf/caONDdI+bEopxX0QUGrqfYET/zEBxyahfm3208e6Tjiow9y
w9Et+08YnBt5rnptcmdNsKLIlPdGLoNnQf6Z15ezo61FKKLMIYEyC+2RdwMUcHbkVGbcrECOG50y
rKh22epRpBkg3qc/ShNJoGIkw4xEbS0LRfO4JH0GbRCw6A0Z2EmK2/J+N88rR+k2/Q9vbWgJzhZy
uAVeo6+G3apKpTZMJQklh9lxU+Ykxtp0uCvMdfBivCNAdWoElGsHzxgWNPFr1hWypHxAYdOcXnkX
XWbfUR8RajM+ZXhvBhsbsi6dc8MvufaBz69iWgQUVZ87RE0S3wOhUMIbT7By1vc5AWMy0EZZk0Ik
zOMpn0dMqhfq8IRTCEBKok8fw/U5y4oztp5cCbRt56rqNlT03JNzdN0gvaIgDdVCDpgC54a3cNTC
lYlxoxRVh2eMns7KHW1Qe4huvbcrAIblpVUC3AsFTFyoc62pxYGOrERDTaE6SosXxEvdlQVPYU6s
Z71yCVcDjfh6tLgqeU5G67aHLz3BO9QEKlrb+BOb+N4ycgcEm2fem87IvuVNtVbPoF2/XCLkSUQF
tIQEQUJ+IMOLdrPYMWKx/ofc95j62WUy4zq3qKiNu418iuNOrg74IEGrxS+J2hN0iOkQO05bj76g
ZFRrFiUejSVYStiltsv/G+HyWQz8mDs1R9wmmFm7dbJ0LYbNcGKvHG1j7QLv4hHy/nXiZEe/OePi
7worsM6GixbQIl9M/R1F7QPeJIcqgZWe4qWrEPEA8HTuE3GZP/KLEhNFrhH6jSctKPtijMz6iI5E
AVhR32hBUNgTWJvzFi4xWxKs5RxpquYUI8iv8FTcUuie7vbeSWVbJ6Qj+Fz9CxzwIGv1UG4BkFp5
jsux/ponfhojNpBE/uxlkncArlAoxL/7WL5Y3W/i5/r//CpYNPIbyTLuUJ3pwf/4nNjal/i3kols
WjXqHbLMBNOpNDeiGBXDC1eAxc74W3mzZrLZJCjXFTDItuR289f6iHERAOIaXCKOCePtEl/TZLoF
c77o5lZoypoJ0X7P6aLbuDwN667m7ijOFMJ70YWvtQZL8CoCUXCeIswxEAryBhIRXWY+9CRkcDjp
GejO2z3nw3yzXgc7yg7AQ32OABGsa7vrtvY3hPe62f6nwF2R8kjrdA5tChyTRiV/08y3rlT72HQW
4z1CuhKY0BNvRkr6A2aw9m70CRcM7KmGC9dQ9bzSu/IT9i6m2PbRMQ96ZIFk3qeFcSAYMBTftYok
bqQiH8ovznhac+eAq+PLLy+LlVwFEhvZ6w+lHH7rgTxWrIY2nLAJk6LZhmKlAQCMAh4mEFpIHUBv
YibN4wKzYzDtXilUt0kOci8drBWWv04nuvqHyW+9LbuxlFiWSXmvL1v8EGI+IEMnjoQmVT9SHlt5
0nAmxijyj8kveXhsgqhEI0T5zZsvR7VtkPjpcljlAFx9XtYA0k6Pn04MbOY5Z+00o8WEOHFYLZ4P
F4Ma9WFeE+gaEcTfBNWuOL3kQkQ0RsTjX7HRm0uoChw2wl/QL7LfRn5yEdVRnVOnY9HOHb6kUX98
DQICO6LxJX+FF4dm5NExSJGK6HwNQP4hUpad0vq5kUgfTxYZ1kPqxk/sboC+Jigmr35XkHw6XAj5
wO4Q6cpL/7e/bISLN8DFcqqKZb+d+N+JpUpl5oUeqJODoNgVEreUjw5yGhXia08k8bmXxkoxKQO1
y6lSijC/+lWRO4rwvxqRTKP0OMTkYUmBuareK+m88Il135sTJnFT2pFyWSXe2fUtCmmBUmy1yAfV
cP2F7zQpD68rirEfgns/5V3CbbkjKYP9J7gKrXiy+ogjTs3fT2kXIqkZ9P4sp6FvUYK1W4tGuQbe
erVlLt0k8x/xOuD3obKPWFxqVfvPcRo2H2aclakqSJhEkTtw4n/tGp6xD3Z2SV690VSCHjcdSxIV
SU3Tx+DFkd3bWHpjj1ZJevS0SRedGnCDWqqoLACtII8UQbBkqN1cpRZDRMbo63vMWoC9VVnfyF1f
SdIvVJ5ZUjSPWHRSlBxjuNwr0gJ70jGVYT5/IXrlKpg1diqh/WxH+cD+/tKpfull4i5z65Oz+t8o
+I23S+dvhsSknYCWUpjPZ4uyOS0KV6uCIhWDV+zaqI/ewFunWkfS5/1W44wYginMP1Gn2Bi5Sh9/
Xairzhx8nLiXh0smMuBHxpWv0djxZvPNyq7b+KLA2T3niF5EfzhWKTe1FbiLXVa3jsQgb2VHsGCB
A8zpyu3uWRASZALNvWd5fsb0Xen/OMWQ9yWqRKBmPdNokawx65CV7uKU6dHRLLUqh1QOdlehqAGy
wax4j/6ciA7cUdf0lcRSFubfvRv5rXJPxrGDkyL4t8Sn1x4On+rEEhRoq1aNav2IzaXdiX9QwIjD
H/gxCc5N5dhcPYFxmroHrHhhU5X01k0YpzP1uctDiK6z7sRamCTk7yAPucVLspJxNZTtKYipGw0B
IhnhxUcHcPt56CBWa0Q5HFjQFvlMqAu5LySTWmTA4ocTMlv7dc1FcVUc2l2mBX1QfxmVlaTMj0MW
FSXhxN70xZaPi8LgdEdMcyCoZclP0DI9E1Z3sBPty6zYXPB87EblKfTrPSjzW8eMAY1HIRIJBsoJ
kVLfWYcPFsFlcQOtE2RfheAwtwlQ65xzged6fWdHWkt7CmQpI29Asqy2RoWhc3tmxa3lHsKm3MY8
bvVyFJ+DMEU9Nq4CHIoQVEypxv+FWHtzk+/LohrupjE7Rp8mzs7CNIlsfeCdqt67K4p87cp8C+X6
UEOqw7YQsHsYp0mgwttQIrnXj9hu6Zws9qYmH38OCaWAFvj2/v4tOo5PTuRSek2iH22Nm+QMYMKM
LRHfePiy8yjalii+q+O6rXRyO5DlHlB4FuNRSRnauJq0pH23LW8vslAnEHPUbx+4q1yRwwjBwu1f
TP1eqmQZc6YxLYvYRwehWKwslA7mukJUSSdEy6HucYQYKSpOEU8gI6gIHxQM/bkVWILzNFb8MUGj
M3I0xHzDFct3qlvIbtPPu+winjvEnaqNSl9iDPQqiPvUuX/0DAMErRCFvaWkcK8R1e5aN/RMg3eS
yH948TbtTQuThxnQ13GY6cHTNLdbMtL6sfB24QxLjIFk69n9efXytPsooKafZjrOd0+XXPssHwjb
7cr080cbuRYrXyIYN4YfIxA6SNPMV1muflhVs0LYtXeztxCiRXBD7ifWfymiK2VvEvkFZhiFXDzX
ruWwF3ZZsEcngwYwgzNUuDSzKFjwtJe3w7uFC2V3BABQH+0cU36Xnnbzjv4Zksf3LZXu7XtjwnEY
xW/1U/ATY0H1IfN2bhZZ0kg/cNBO/0LhxqawFoNA2wQR85vt3tsqJkRxlZP36UWEEKeAH312nk/5
hAEUtml+euFV5+eLPg4nu4XlKZ7PjhegfXvPheG+wDl5i1kZjXGFkT/gLDW2Pk9rEfJjCuZAvaC/
rpZBuL6kvutL5kdC6gfAQSo6Tff3yzBfklQ0kC5GocGB9h6oKroy3Frf0PUeIIR3Y1WH2EobTtcH
nVfSEyzfzZNutUxt+QoBMfnMN/KJO2dlLET/wAUIZ0KgbkWzzH0e+/YWRUXS9ldNgcjEG8Qj+cXx
NbdjrdP7M79CELUXMuyLhXbkxSv9hVHxM8JF9QJGxRpKM9KrXNKuJANzjND3mH8Ej7BivyL6UCGu
m6TCycbXkWH1HYNS0e8GUpHoz44y6/zZ8WdG15b/8XXa7eoOvVLyBKTGrsKJR+vUYBtohnMSNvUW
O6DM5Ghjm1E6h69V2hUts2O4L3WGQ033bXmu1JWeAGZDJbRvS9JQge5ldNHy/f8rUD7hoBKAnGKU
Q3aFF1bpuFuNyB65hDXz/lZJ2PfHjYwqkePnDs2pthiboc1nYICKGncD/6R98KaS7phlJe4fV8yL
l7eZewektnVCu/pOf7k6CBnrWkP8cXXHwahSLWeeHghO22g8RUwkfZWYouK2n0FlvF6Z/ZqGciA9
kNcdX1bzZJVwVNIJsjdH9DnfvgGT1QtO40XsL19rCjDrY00+zuhq0t85JpeTk7MqTtAuViYnp/a/
voCuPlA6sWy/kNlmjycEfpBlEZkQbp66obgRfQ4gqFZZax9IgHqjycgzaioO9Q6T/ACgU1kJ5e3i
a/0/+81+9WB2BIID6VoMPFwOKVS6JrBdAPu6cmLEu2e05g2eHnGYtNeGYnJJRiKS78QpdHQOJ/q9
WRHc2+CMerj9WMQCq3SQGxzCpcVei3skYLjaHOsrk3JHDuASdyYBCIXItbgHpnQM7KktyNVS8FeE
KLbWb7i3HC/YY2yh6gDl9ld/8FQyHLartl8wevWm1W88XYBItxwFWNlOT0n/bItK39FLgbVT/XQC
tRQpwHUw/2zGPfgoO3YKYzqP8frUTjVwJ7qvcfdtapA7LBCP5nk/a/bEGqG71dO9T9rUB6N7BsK5
Nuih76k1iNLQUpXl8NV/ckNYfcdC3sCEljKxAC0Bty+OQ0H++lHJM+tagojq4IWBZfC707B74wrx
fjhDX0LQJCfRhXJUJ53ZKh1WWlOhI+MtkDtohvjJUpTmFAXKHWmzRgcVbE6SV5SrfVKHoiQ9LA4J
Fy96zTEc/nQ4jzS0HJMVWm6qk+gwdr/YX1YA0fn9s2y3c5XwIyrRdDC6CejAkJY1GpPcce2PdjOg
urg6PPj8D94d71seC3gf35H+sPwePMT5DwBksa4dob/atTVnag1GJNkd50b6wdeYBeogacLPvbjd
s4hA0/jPY7S+qJ2dK0Sp9g1mSbKGRPQLKm7sg6PSWCyr4wWvfaPXiTb5HnRe5E24Uvz6csRGMn2F
gJSG8MnRfdbvJXvdIJC6hfPsN4r697JgFP7icLLsFKLT22W8CCJhwvpCGqDFHNcqx19B1Cnpn0dA
u5rC9h1muCCKO3VJjfm/6ST/nuAsTYlic4+9552gbhIZ3CYJn0UDrkIrLm4Mkjzz2jrhSb/cfOOm
mi7oWZBVrCR01jz9a/VZK45oa+sWJiD7sE9FJbtrg/lNg6Kz/hel45veJPMj9uZ5gJYmt1Qnyj7F
mr4Iykcz1WOV9j98L67AmYhJHJLuT0x4mYnDEi+8eLjOwOzHXT5103YOHsJ9Xc+8/dDjp9JPSR4I
ZRjHqv7HwSjyHj0f+JZt6Sehp1sbIOSxeR5QMzt+Oy0dBXnKpXKl2rEGR594+36sZcYSP7oT0gVu
0ElHiAceHiYxm3FslkW6C6INzqf/lSX97oG0lU23CV4gAB2Z1D9zgi4UiN1gH64mnBAWtZgdx4S4
povXwGpg2JGm2Rb0CTnqJGqQDagBWE4gAGe+iOCWij3n1e71bljZrvrvnaSvvVR+SAj+9OuKChq4
ClNDzC3Rz/hBrVceSpfHZ6E837dX7RYbyPOn20fV6nI5S1bSFgSlp33BnQLBrNIQHiXp6vu5pKUw
KCytq9ultuvIQmobJ2Jr8Iw8Gkao+hnpvpDNOsuxmWw9tugKUAdE1/nxMV50V9q4C8G1hl6x0GSW
3heKoRfJ1Ns5old3cqLX2N7y3+A3mp1vu6ewLZz8fUzUSsGSWjQ2t12RNaA8WpL8RehhxQN+PJkF
vV+rbae81BTqEW+NPHu25aFOIzFKnHHWx9jPx1LE2sbQbsDfi1zIMKt5hK02MwysjGv4UZJYzTaH
aVeLwRr4Q/5879tYLVcp1x1/eYX0KTiAbDtT8YyOrYU7FS8Grz5pXeonO7s0+/z4bVWiIGsx5y0Y
plHqynXs7r26kRaY1Wo6bTRtdGHjM2LopLuG5s178rXACjGe8DOwjXsE8spwHGWmXR1HxokJBLPE
0bGUUvK1LJvaA5cRiWuCvaicd/DYnpYc/vzzG+sYP2Wk841F7JHOysP3/pskbzDMm4gN1LUKVtyt
lxuBEVAvyZTFoiq8/7nP303qZRF5bLCTEMfp9nqsMzoRpDvngQK+fT3Ljwo8/l2D0mpH2KxcMIgJ
f6rHUM4ytVMgPWBCKDPEmwOtwTUBgq3uzVdZ9M9HYeXryF2xubgBSuT6jk2outklX2hwOwyBwul6
qicMNS5qH7VBRnkvIrHwrxxl3Ji6MYRFQrDuDSY3lcXvtpTkA18/fICCOdNUOz85QzYgYJovMSIJ
ptN3wxoVz0v+tTkavIwlVZ4nZtzW5cf9VsqoA8uaFN6e2/qhq25IIHda6CTpjKLJRmL9CC75p6VC
0+IM+cCZ4U8KP/KMWnh3M79DJ4SWemHq8T2V1V48KCU9vARokrsJaBghgkksL3daHSrSZo/MQcxu
aAeSPjLmxMgDaix8eSCihm6yvDnhSqIO/QQv5Ltg15hYKtDzNt9rRICedAf/X/dBC8wtfA4mTPIe
icwg7rZoB84Z0JeCdn0bFhEzCBbaBuiW2evgtOJaZH5/69wOkVmgqLURIDQkI2txkUr4FAzjYrZb
iBGrNBIAyQBKmNeTsf4dsdMtUuipLha/UiSrlt0LsDwVnl5QGFPb3rDhmHR1ISh2Ygs6QXr32cgJ
ZMz7/9gs4yhJIvma8eC5biNjpXEnow/mbiLcfM03kVtrzf1FMjn1dmgZU5QHN5xGX56uLYtbsYP8
zb84sWxJZCkezKwiHk3IqFM9PkQmeyYXvmNtgXWA7ftv70D3fJUkQDE1Jut47L1tudtePsOT+T+X
vfkeVrTSlknwql+HovXTyL+freYQMhWI3/TeWVU+ZxPiYQ5u7pQpGJypUt1egaXJ4Z70I5pXVPtu
OPERsOniYKuWzAQ5/RNoDo9ZJNA+RijYL3cgz7URefpSSGuNLV7f+ZgUbHEF9+RO6nBLjsJlRE/w
id177yhYq9zTIlywhFw+0aG3cswg+IjDxAA1LenMcZKpCu4dnEOKF5j0JmX9QJdcNw0rcYX1GZhy
0BxhECJ1UPB7XiDt/FarcAzOef2klIHKmOx6ryJDg+V7/0C0ppFsUZFmeEY3m9MR2idkzDEpy6m0
hb+7drx11Z8HQicCYkPie+5Wj1GnaYTfrp3DauguXF2dNz/fHn+DqlwM0IQjdh3gswDvO+HaVXfM
40p9DYDhXc6y0ZVZtYBLdmZ57H7+LkybpEmHcpwsdUEWK453nwmOjjQFk3n9bzcqF4rbWJkRHlzf
Kho7nF8/xbYWfiUBEqLYviAv5+lUHJpyB02nvLr8JasqIdKD8ZlNEqcB67fKn4FCsyS+ia9fHxZp
o6Mm+30o9F+1Ncb0zeESX3rorshjYePTFwCJ2Z50jgiXRjnYEnxrfw04G7DPpXu3LPRKHZjLGOig
jTqR4DAsL0BktmWNnL/62fTTgpXm9f9q5gn+z6OGBxgJ0u2uvrXLK0FjgQzv5vP8aYpSaAWvZHsj
UY3SEtsE3Idscr5IVNSmi3jPoCexexwD6Xhp5nP+qVyh4yeerZjPYxM3BnvCdx5UKjcJdf5q6ioX
2Vck8rVB6noJqQgoPw+X8Ee7fPGiHP3h+FJJuAyp6cwIkFnvPorOeLLIJVqk9sre+Pef7uoMgIOV
her6FLAiahX1h+j0lE7x/+KTL0Tgaf0aoPlI4OBuy2Ax1J3JLzjtNxsvfKt8HjJqaOxCjR2MMjAw
oP+qXfBIm+jFCqW0jy2ERRWfOgvfC8HeLx7F48aNdWc5JqT0eO5gQxWEdO86OQswp/gL6Juav9fs
0EllXhJWFMPnhGOqpFYxX6fOLZUUtNYLEG/StWWDq5nuEY7GSkT9P4ZlIJd9iu1QglkGIiCmFyYg
51U6p7yaz40IoHhzRFWsAFb3ceYnLdWlxVkt5+A/95BQ7mT3U2inEb8cLLZkRembhkBmPiX7Q18h
mAV2dkLl0czzH7y+zDeEE1vz2pqrT0d5IreH0eCx821xhrYKiZ5GyIWHh4wWSXiEEuD1XPvTcbMx
D4j4pVQhiRHMeyD+8YcGGPk+N7aP09L4dQMqML43Jc3JOfyP2LOHEbkyrhmt7Cnl9Zi9FAI1WMnI
4qvzPHEr2oF8UevzDPTAHTrK3a+PBopw9YALf8PUC9ZmToLqUhWL/dUOYghGEATPYMFFg+TLeh74
nmnSrFbLVxJ9Z8HgDfoerXbvmI9SiG1Wy0nV0C3ADiY58NvBs4higI7IQhvzqdZnlLZb7Z1IViz4
isbkBB3sNyCbUo2Z8kQJzdMEzKMPCxeIkrSghX5dh1vIGNRWcCDsXx4D0xbQLjSr0KuA/NRzx1VQ
6l1323JnUFEu12Eu/nDQJx/dohpxVQdk6WFQeDV0mVvQuEQHMivTSNezZmrIBnkwz5QO9LyAqJre
inwi+fJ0T5iolXaoEkj2oJak9KqVkuKZ4fpn6UiPU3uYRdKV/oSc11Z2Db70LpX9yruWHMfNBuGZ
8t85CW79ZJxwDdHnTxaSFgFhh04UwOt0/bXv66ECfVD6dzkzOTo1ThqxuTBaTBXAWjp+g29Ga+5d
oHoaRn0NtkBxfU88Mbh+aXqpe9sGFpvc1UKs8wBHIHGxomowbeHgFytGg11jW7o1U3JZGPyP78Rz
ePl4Sr1Im4gnW+IDfkkhJQsBZ5e1dOJZCfPiGMA/Kpm5uMdxhJK7Sy7rpXptPgC5CE2rRnDlxfdE
yLnJayXHsKWpKTLLLok6eXOdJlisG5upxQ5X/qnCSWwoN2rL3VULbqvYc/w8ju2/wm3/+K3lEs0W
zezGp6pfW6+2dCKAo51PuEiYUhXQbSnjdlZWHDnJXzCKqvx68KmJHP2euLKVtNw2ykBGtJcQlwVl
AWLG/zfv9setr7r6accsixxlVgMJkB/mKvIFWr43kWmyVZKncQ9pwioZeziOfepv/s5uPxDe9MB+
eylugopi9EmX6/gN/XK76nNgFDVVDNxA3Vf4k2N/OrktxM0cs/5i5LHX/9uIy7O5whouFSYu49Kx
kJZJU1rG6n3jxU0i5zLKjDF2sWYAygJ7IAjp5clsLTw8/GQjRSwW0+9+/2rjaqOhy7bUsm1J+xtA
ZcYoa5le6ge8+OAJQsvVtXOhttTJFM+TNByhU5Xyarw2nS+TOma3Sm3La6RxddsCmYOEVaMOYOWq
t6pTvUHiRKaTsk0+QX/oSr5IYko7EFWkjnBEnvmtvD3j+qZkgYfAyXx7lQhopdd9Px6j4MOBrizt
c1QqWGI8wki4tfycyJevx8B6Dk7L5umWGRgSPiw2s7LtPmh65EBJ6m8ENDY7fSvlqivv3A+lpv18
llf9RH+SrAef+leG1ZnbE0APZBaPuANAK+HrsmfifqrpR1t6GhnjK68Pb+jSyE2fkWbHcjwIQgH8
YkhXpTBgDPV2ScYCe1eYPcylyf4QKTkYB/q5h0anYEnZtXyUHcHTjdPhXWbPWjWB7fYR/w1Kwa1k
ylfNWodTpopd9M8V4+kbPsuedMBiPR2Yd7FpBJ7I4CqPNoFjKPbKDIopreNOBBK8y2CQQeBc0c3E
uT3FttuKdbEx51ozFRVveg9VgdPfmEIQHUR8D0Xzw3hAJQlAIyGFWsuHY19mSTX0AhpG27G/w9I3
z+P5X9VNZuGLzNHEJ69AUYp6oqxhtch0lqT2FfmGA+WSl4wuLJOD7Ra24eZk8awLeGL7M3yZWz6a
VMQX+6UgUerkvXX+m9yQZwoqKNQxlmb9OBYE4yR0sMeJBbSsLzj0g6K0RAslSYnDLsauZoGcp0Rg
bE5+7JK9zKcW546xwRNQ2EwdiDdxJLZOj1AFoPxqDw+LVLIjbYI2GobDvAZ7K5HYXYCvxkzeAQnh
3BhgJx1n06NuqtubLDW7J3rhWPU6AUuvJDpL8Vi15Fhjk44MWo2FK2oU7nDVjZ/CP2Snmj30nERV
9d9hRzgZcHx6b44zF87J5e0IuQNgz4qXDXU34C1EWCkBMsXdr478OyOlxnciR4J49gv0l3C1r7xm
R/1spstO1PtbPATpLBn4QvK4wMKYLgsJJTecVROqYEHopDmN2gJMgdeLQftW1yJEpB6CPy2czA3Z
6NAmQcUH3ELjnYOt5vtpqkD3cWYqqlhkGl1+3K3iQtgi+WdDKP9i+/qF7+qI2ic1b5kqB7KcBQP2
cuw/P/KtSq9mQekGL65KdSGIynBwQWe6yHcdXTyKLvYaA7lHg3sq2LbyfCZi9MOsHIzD6iAuNNsh
HJvzNXm4of+JOOcQaqRX/+xcFfMiYn9E6Wk6vuU8LiYdMcfwqPKFuX/sL2GrogvJms6F/U2K3v3C
xF66d4oVK2bpV7vG9/EgtVaY6XbOzxDynQ9GMEm5cdsMjhkwlrqlAvRZtUuzGvcSZoP10RG7q2tr
Y0ZrcnmmGsM5Gu3MMvygO+POjNfk1eXIKs2AGkKKglbsN7FyhJvXnLc0enxOTfuvTgQTEuEOSvyz
HDiICU80KE1KyyOu8QCyrd2+Xf+AhHEK4sRenVXrHefc8TE4jgyFHYF8LP4uDwKyd1zhZfjwqlIg
fZqaH5khD99bot4r/QgvFxf32YnishtVOfeLb+MzcPYPExQ/Qo0xsQ2rdYKfOFhBr10gpnzCBPI9
VDarIsp780iAMzuEJPZH/lAmQJ1CIsAEX9QILXgRyJJzpwmxo1cm0j15/qfrwOIK9YLwYms9n0X6
Fj/4XdPFFIVQXRtTdQt/jf09J2lURPotbUDzYJ3olnMCY1waIdC6qWSenM4B/4NMyPFkVv0tzJFG
f7pQLU42zIUdnaC+pqwIkLvw0hPPl4iMMQBdxkr8VpBdd3LOW17YNblf2NCvpYsJYVqKU5lbrdDj
G7ZxcDXyA0CMYBSVZgtG+VGV76WUkAA/Lys7zyWc9oI/zw3H0qpCI6siKCQRMhx1pLMQULMS93Xm
jD4X49cZKATPY44QKtyRihEQsNVNdvuJOKDPXio6hyBNWzVOfKmVukO2x1ZJcEwZWYZijibzX1ju
jqBySPeTq6qVVV4t4kv9ievm5tS2sM7uq5XGhSd5bZu65kU3pV3PdB86FdvIo/5NJXC0TDG5/rWv
MBNp+K+P2GMLB+SgDeWhwpCiiFa7q5zYn5vz43V0GPIDrMAAQyM74PysJACIYWyBvEQRslzdxitq
QE5LlmR5yBOyvmvr1SgswBeJdHM9YIXCadhmN/1tCcdlbBiAxpeMLsGTs+dPgnHkT1o09hNILVLu
0cFI6ueiUmfH4isVKoLbDnTyvramqGdoUEVMaiHmGAjLo6DdWguAhqixaSEVshnJ7R13giueNNNZ
bTNAlqgnWBasOO6Zn1v3fFKL9YnFnmrGmfzSPhQElW2VDqaNbPtRNhJv2Yjr4XuRojohwXGZaTGG
sl+gbyjdMToeTmS3Ck+d2mCupotGp+THjRINLqwdbpMuEWerw+k4LbRQf1dnlrCsHreKyYFGujBJ
wwL5UKl9LvlAmWbjIKdd5G5Bj+FfOMNm95SNBAOGSXONf9A9SnOiBgjM3mURkYSa4Rh8Xeu+jQ5b
vyoFedbl1oyDBdr0ahD8ny1T73xPvNg4qeEnXPk3dKhYSV8PGWdnOJp7aPGUywsR4N5Y5uOs6Thx
pbpqRTzty1u7+mPAerkX4O/xZX4QXAbKV61ps7lk9Fi/L1ZCtf+h+LhzJQOXgq2vwzk7ynYeKhMc
B9fYJ5g1B/TLhAH17wSZt/8a8mHnGFfUqwlA8jg+rAyxns2fDbnyEdV0xCxScsgYeqdzqGrv/cH1
mv8Qqeb8PZNQsah+PnUm3cmS7ZTmB4KQCR4+NDk8jed1AR6bV5fBqEo5WQYqWHm5gxCYYGTWWn4t
45j/k3W3/CwcuUEtdQ1n7UCJs4zWhOJF8EsAnqSM3WGWpBG8bQL4P5Wy1u+oUBBpI4DLwQTq+MNO
AU0EhPB9QQi7Xyq+CbMa/E9ff4zT07Xdq9ucLEIxi7iFC2Cpu6e4WuR8M28qsRNHuLrH7i35ELEB
M1kKIJhIvtS5ac+Ta8FxPHQGhU7kDVapdxTEebkd1e1RcsMx2M60HoFQhNSAMHGwiiFRP0CDjVdM
9l9t0XfKpR4d6h4lF1C3rZUOKo7GKMFKDGIzIwZBuo6j/sitDXPca4W0Y0ldWyCBuoeQv7FrMJix
JncYZPMMxHu13R5sRf6hAeCUmN1ummgXdSdGpsGK2rpoDtKwKywZCKm3pi2IywlwvZ0z2DydSeb+
uYOf03HQ/ZTbYtgskSWG+GfbDgrUezbf42R5XPQXnltMdBGs3ZIlKVAs5m5vb+Lh9wx4/fjIrxf6
aMgSbO5NAAJK1NuStXE2Pr9ATipcxnENXR5jFvs982TMwhjDgstjnVAzb2uPvSDfpgRl3wEvoo7q
mck+eG9VMHFTBG+o0KDgfOGGm/1z8ZAYrekbLa5xYsGkERx8MQ9lAQ8r15+qqIDdCdf9qwS5BDnR
ZHvPS/WHCNrwmuOB6wb2AZyyVk8zh+3r1XmlCn0bq+6tgdz53IdgX2YtGWoNNSSrmZIs4/vMEGlz
u1mjeqbcba/e5uqgi1BgHnNpUzqsBdvL+wAYm1SdqjfpDDA3OzXAc2WQKel1pmGKMYYxGjK6Jah3
GgAKwd7brXwqWmpU0IBmuaY7eMXTcDzg8BlosQdzWZOFmdbmxgKI4cu1tu27hnpL+JAIQ4TnJ39x
SPl38JW9fjI/Zlq7snNGUdcaVuWqDHfwwEGmFC6Czx5LZxAhgV9OqNQ+XFxkODsJ9PprMf9W3AGA
fOmOnHvCjvozcX6hY6Ej2xh5p/y0vfjBVbxMw6EtO8qQUK4eJsp/wDgvL5s7J2WOvz6TByejkifR
mpi6Nv0Jgd8RHn8XmYMlIaaRu9ROrTWiORKdjHNpzioTFnkWwbWvQv1dpoBJNFNz9ggOmuU+gtrn
57Ij/afW99JV+5uWh8hToW2RiWj8Yqde/tDmPxH5dMxcSK4vo35FG14cOjCWbf819m+m8tw2n321
lUbgwH7kYFmW9RDeRiaVGijdMX/LDdPp4ixNZ7BWNMZyDaoNYPgh0t+a4vp6Y19InV/bZjmRsi3F
TDwjsd1PJl9nxFJun4AdYD7X07iakDgZ3wW1WzLtySvKn+HulGzdoIxb92RPASuIH2T/WpZeY4bs
XCjRpe/AQTwiyZBn6R1ClLJuw+7gwdNXhM8nXVo4gIvkaad+gN3ezmFfIIL86unLknzZvIlBvKor
ERYaiH9zUPbEIrUqBV4sP+IJSwW6Ym9QBWDFSOiFU5zxlouRxwhK8xAfYRoh4+ZQgqSsYjv5cZE1
od7g0M7WpJrwSBnY+A6xtzGDkan2a/vt4qKs6gzw1B32yWORcjsTovu25+i/vjYB0rrq4b/KCycq
XI8ufdrW800gPsoK1O/EebZyzXJ2JXxzv2JDMNzzCllo1rAd0QDue6VVX6usZCq0Am6XosmEB34k
B0WMWqEB7QYRrEzEuvMm1up/Z1j7Mh7aalwGoRcCYBlVPsvmpqjb1SMWKqrsp0gMddrlx5ue9/zY
3/iQjIPtXPEDzfmRKPImooeOuJ1oW5bNNj0K2XZNgkH3Cb7sEqM7UORaIqNkjCZC4Fj/luDPlb9X
aiy7dj7ZXavPqg3lQhWedle0kRKDUHKCx47SzCNZfpAfjiwYNEhs0wuRjUIFZVq8wfXAJ9N8nxVS
UfLqNSh9TySLnhVSrbHc/H1LyZPvGZVdlx3S5u4i6bAdt2D0Hr8GPWi95N1tNISOvV3w7uhJ4brb
od9uv8zxdrEuyF/CLx1Mdg8jor0U/wPm4sfVWovOryG7sd8K665WpN/rh19+dkZaqJ2JjmVqjQPI
PNOo9IuZo5H5ylA4pt3SDRTO1uq6GMlIKWhxPi8tNupy6poFJa2zHfy5Mz6uPGeOyqzmI4KGByoT
hqB0tKNy2ef8H1bzupcZHa8Jm5kp/3l8sKRkHrTV87n4PoiTu3ymMh+CUYNv7OSCLDF8MmHmZdV/
ehv/bP2ljgkCaPhfetiowZdZHVDZQK0ZCkvlSFhBVAYY2OcMgHEiTJJGRARUop6H9QTIOAYPvgKt
laqNctjzhBs8FbA1i8W1KivmyKmWFZbZNDS0twJeJKAQUkKuGTfd4LCcB21rD+OFq2Rsu92x0Yao
F8XFQgFwEGuGBTgYiipGfJnN4nwWt8qrFyBZA9sQUs+wJiXAqqja5ojUB9V+l0ObBJkW2+kMx+5S
07l6+aj9EtPodS0VdgWwMYsMsJtlArKBEGhJiKcdPlmrK+cI0PTOQt3XUB+cZRFm16fPMoVzwkCq
gGxx2U5gHWb+7Igy9G3J6p6FyE4mU/8yeoIhvdVbh7Gu3ECHIX0jZKIPYUDZi9Y8bqOXnLzqyxNT
gvQJSfvoVVHcp+fcOcbiWcqphSEwooeRpRXExi349crdPm4v0pfxJZDvPACmUJ15+guHCY9GnqES
jOD3R9RJePm9Qs0TOLzfKF1YiGXbWA8SVY4leoE8X6WWM5PDurXoCFDwXsI5sW5MnVMhFfiL0vu2
gQPNY6DwdLzEkR5/Pg6OwrZlkpaftP7hBfAjxYa1+0EceR0qK5upg5TzEM1mQoKLxDKLN39U8jyB
div40Nh/CEZgbz03T/P3NHBAcBh9Rx3JiTCgPqfchalZ6aYS/kogN+YOCOipoQU5U0FPAdnF5GOA
vJn6euL4wbPDytjZEi7PcZG+LfikjugwQM+90nHD88NfCQniXQHz+Rw6Fj4GhxRr7cpoR4Yt+wwz
xh9CI54akkWt8bpLjG2GuqVYBVMyuRguhNHmxR+pH0IiysoPLTgXtLLF340ev8UJa7CpzZD7a/dq
zNq7EZcD89vxr1MV3/clXY33xaUFlOCS2bMpbM/Ezgx7WWcIv7NRaVtI2YUyZux+vWds2xCCUwwV
NZH3xcCJoLXK9yYTh96f4lZDbo1evGt1Eh4g5kjn4Z2hwxdNCnpQVjhjFY1YlYcULhT9pY6BT522
0zde1bf7VIw0xT/b7mcj0B23jSAUncvuS8sywEAVr14a/BfynkmZTcTbjTmOdWH3B/hFGLlOs6wt
FXcchJ8IKaQ5rVR8qZVSKvpMcmbhvOU/WzhbV5xrfLb2rCNMPWwWsEEQln25VxR5GlzPWzSmRbKX
sTvlPjbmE51x9KwsKOngIKVhKP1PJu2xoztW7bwa/XA+YNWHtrCLgB54px56wCNJgDROngt4KYeX
7YGtO6CnY//RdSoLmXJUEvFYTG7wsEoEcZWRPm/l3Ru01gzQ3iJK900NsOSBk7DQuGJWCXsdMmGi
li8WDM3nsJTVwYs64x1a2rcHc4vNgK003nJHHmBSGi8vTHJP0OGP8hgGUnX05Rtj7WkNergGPpVN
iUlOhOmzZPsx9CtGkG6EzzodNXHEaeX7F9rmZKFJ/r9kmOTcdLzNSyQmgy2xzHLG5wMCsoHeOHHb
jTokXOcOPu24gi8jB8c7NMgDta5ktSy3GhD1+4lWZ44uPevi9qdVs5I8tadncxOKO7TgLobrIiSs
kKpBKEQsnGbQcNdDyWD65jWu1Nc+gpSIK3MV/yeLPf9a3SMrIV/M66x5hilAhiraKfcs2uhY5FDN
MiSpPNM0YswwH4nBjU7xm7MdRgdp7WVI00OECzjgr5McnHZHUJT+gN3B+r781Lijvm78B3ekSd96
OpWvDw7ZdSUwLYEKa5IW5Avd4L2i785SYhP8sw3rKbtT74DkILIY+j6vA1zO1rBmi6QwpV9MvF1V
WRxYuRd2WAHP6PFeDcMayUlEfx5UGt2pjFuBmxO7lm1+yCX7ocPpsR08DmLBWlQlDcu3asjyQZhj
KwpJfvdx42VtlzjOcWtDlqanZ3fBCx2crwytGr6Ebt7+zqIifo4njDlFlwiQebR34XpoUPCmzjiz
8yrdEddzMZA57lbkxKLylETX7pw+Tw2cchN5anICYmE+bKAAfVONOkkL5dyzIipZ8dDTNhkluprd
bvaNM+9/jrUsgzG8ry7KRvWSyKTO5z5Pxi/oDzd/TlC5fA7JcFfRmfC/8P/jhE0UakC5eDWSJem1
rgcj8Zll4Xpa93OrOeryB1wOE3N6WQhLTW0J6DXXqcAQ84ZsbvKmhTvlltUatzoP3hfAaZmpqsSl
cbyOnldJYiQnepPeWnS6Y9T/ISOsK/A/2o547z9hgXHspaG/zQpy3axDfItfj0YxtPoswmx0mKR9
co41pH5MzR9bjhx9MW/GUTKASFy0dpKc2+ypinONTRrd64pKW6WMQpobmXhl8J6LGB+MGqnHYH5M
LUs8/6YZrnmWsUT9hDXSsA7SmYx0LQNLX6cTfqd3dTI6aEI/Xqx3x82WzcNrpG1RoVPagqBuBYDJ
he43euS4J0NHJD0rrpUdFXvMqDcPEjId6u0SSu6BACTHi0EgokpeMMwFsLmF4KYePkZu8MB0YIOJ
7sIJMS95dKM5wpOl0TyMlf0KcK7FmNtpxgNxGOLVig8nwevKzKT+er83LDaaHfVinRGG4VnmPNTZ
haD1cRgt5VsNML+1HWG1uuAWubOEWL9ILH/V/rvnrkv6qG7T3j8xPghljhLgL4OnEF/WM2BalpEg
m+M2zFFpgj3W1AFUtQp39Qzr0Jjx+V95IiXQHmEve+OjvYQiAZtO5+moReODHKZyr8tvszNHaMbK
BeUGUtA0f4p8VaonkEJYvNgxZdCBS50kpRK8rL6kxJ3IwMH25JAYK5I4muvVD5rWrGJ795lVqu9D
GahpQ1gqyF7GkJ3yXaaLTTKQBLDPd9Ecf+3fbglIrOdgtl7JNDylScY3j6WwHFMfoCBk38LvqIlp
vlhu5Gd9ai/yJyuaSZiAmkOJX75tuUH+37eqj2v4/5XgpUi8a2qvZTVwnTg4e9WGyDgn4XpZyz9E
6FlrtUotu9q5UakvdNbZTkLhfH6WN7x94XkAKTo9SLaKnH57cC+4qaV0WYC6V/LcZm10DBH0x17O
n5eOwiy+1+ZCHsYkmU5gFHWSaVoxErF27J0w0Zq55OKj1mHjY/HoycoIiBzhqE8YykA2wW4JWxMw
XeG6oDWm/lYWAXiUMR3Z+Bz0gsp3aaT03AJaUUcSMCfP83lreOZt7CddEu88hnXcMoUiVuC07AEg
Mqjkp3G4x9PndrZoNJQEKAd8HIw5RBD6z0mOE7K0BQ/EuZkpZScuFHoPDyoDsZW0X2aslbvoo4IF
49qSsKV1thMr4C25BsKN2i0Bgp3wx4X6l06GO22dl/e6AI2DjVYWGFt39ZmE2gRC/Q+UArVx0QFX
0YpoAchCDkB5NWVXV4/e9d3eWiEwkwUnKPvWOFzDwkOrY/jNr42X+7UnmmCOgrTIBmoWnzD+ZTnj
oepZcGYQtgHrGwxZHXggugv+6cYuQ5KMQ7iGOvaj84TgG06vhJ5Vqro3e647bkeNcvtGlOGhxeWw
Hxagn0cjOh3NMhIt2nP8iuhTxUQEOzPIt/4v7SAJ3jsw6oHr7gVUiY8C8LtRFC8gJd1V4QJuleZ7
JmpapyJDet/xvMnAisBpTSRg+QPg9vEk6J3DOhtn2oCntNVifPwJldV6C8gp1BBWpazTc8oNdmPk
2onKCQWtpzKDX/v0AsSRwbwwefESxZjL8udyRpsLtu4FXZLCWq+vJnKCUtvHerq5JWAytVcIDVvY
LEsLbmrzSTEoJe7LN3Cf4C/nwjOWi7rN5X/bmE0h025t8B9/0xYM9cKQwwC/fUwnG42Xfndoqr+B
a+4mJflSJKwonMU03bZzXmDZ2cOsFh80SxldCfciiG+h0dsBjyH19gIf7Fj3UQ/W2QNQPwPtmrTo
YKZEyOLsEtW7A4TOvD/Ahdfp4C+KE0zISRTxOMtOdS6sx6/P3dVXvG//tgQO5rJDGENvU2qlkQxm
0a0wvd66e5KWo6eJgnhyTWukPOC0g0eqVovP+8xJCEFq+c48xvDoSJi/F5FXl8SPm2ZOjm/XvgvK
acceTyR2DGhvuPDJ3/O1/TkUVv0g8eCvQO6RyHux8rIVN/kRjlbuC0FMdnFeNsGsjaxwas/TCnyY
ZAA4ViSr3J2z9/Ldi6Z+kyFeAwsMI2QzIcinXIvaEJ7NJNKnEwhCaoq2S3p8SggoTiNn7hI23RCj
KJDvhrL/qN/YtCBfmV00bnLpT9bAsa8YJUO1XBFpnLmasNzzgUbnnTG4IqIumuH7zMgqCDQzu/af
WKofCS8QzYxvoXyujLIPR6rAk6mk/bpR4KsLnS7It907SigcBzTLbObCmErA6Lh+A6TBZdyKbtCj
kNP/KYC7h5WlW5MT+m6jjGpR66b2xfeDU4WncRu0yMtexSd2tCNHt10jvoE//kcR2CYCuZDBeM0E
StpzbMWpWVeXjXApXJRCKNlhdT6o3E66ZHoBLDxe/oFZZa+T9CfA8Z5VbDs1I6egptC+swNy8pgK
4FOzxFdMMxTTOvstim/8WTcHQ1l6tJ/LJhwkO2b2LwYn7GZeT7o+/Wxqput9sLIj+8+ElRm/lVOL
bPIbfkgSNtjWD+/xeGjDBBCoWM0ZhrGVcmX4b6uyeorihTRFH5wCfbqrtohJN8C2X4cnBF4db1eU
7Ny7601diVELiG0VRi+DUC0XKhPWdYHd63LeWDhs/e7ioOIN14PUKarAw4EE8aGjrK5uY1SOFrcJ
2pMXRRg6o/E/ntLU5PgUxrUlygNnYF1dQkO1JnQOE+Ctkrb+Mmh46NKwsPR6rmzgXtBxE/Afpz1Q
3sewu8sTqfX+eHrF5AtcuWi2ssTRRZ7JeP+otTApUvuCVmCPMIsHyfSItQsWZNXG0Q2lQSu+HzMR
cD21fMtjDoWRkDzxfI53I9vff4neQ/kOxb/OsxywLZ+YoOuLY/IMCR2q9aPv3NoCpO2KYOj9qZ4l
QgV0GVHsN62OsGJA6aSshpZyMpLPRBqYC0V9RkNAwJaDcW8GqpT4JlSXXfuJaxodQtl+dlCo/tLY
V/6TeuxJm3iruiublrOJp2eQ9VphOpj/RRoifZBKOd9naElM9rJSe5x4qWp6oQdgsHGRBTsilOje
VcFq55MTI25WxGMavUe3tCNTYebTf4YpDPW6L2ZhDygOEfnUPvBnDrubRYk5gqUERvpt/9frMzm2
ntAXgF9iOn9ZAcFiKV4FAOeFVIXJVkVZ4V6r+Uw8qN9TA9YGyQAHnYF7f4+OrOOYPQwZiWwS2oz4
JDzWmrr8ZLOwCS9Lw/ivGjfHe2wTaPJuPz1FhXCdRyce+77K+qTPweenK2fkJOw0fvLPqwXI6c+K
YumwMEWbzObcd+UQtd0wJ37f3MgjifF5OvShbeAsyn5KteSCKrZ57lFm4JJk1hII5pprhmOA4wbn
JAF1XXNV9Cqq6uEsHoXruqLnjoWvRG0ug5eKB+h+AQz08pK7awiie//n0lP7/Pjepj1+J+rVUHyf
lkJZGxMZsNN9hRucvnhNgEf9xYKGTYWRU1e1Xy6j2eopH7aEQwJwS3m4eAeqlLVEALPA1PsNQ6N4
ssVYldLCw0OilLxEkiCCakd9y+QHyrQASqYqs2jcUWGLGfG9aMNSmOhcMchPu1klTl5sNhbz+utP
oK5Lpa+MvhMgVRkCO5r4mj0DUgyXEQoKKh/eKLuVOgYgP0ZW2KpcHb4R85eXThHV2h1ljK2B9DX6
yeC2Hcxlzr/cgwAIoUcyx/yJqAlcRZzi+/eBJx4ABX75qsuksvVDMPDbyMgNz/fyuiRji/FqfzpY
U9TjyOJ0gOWMO40oeyItsLEK9VbuChxhum2iGkaEq6MR3reE0nGstxm7HKVlyGe/YFe8HSr5HA+e
ZnPosmP33Dw8WNoUXmTpMHWVe7jO6Z20QI0Ir+wAf9O/yidT0g8PRni0Tc3LHdU/dY1DCqs5qzce
GIvkjn5RT0spGg5bf4ylyWyIi94GA58nr7tpBEIvVB8YqAlFglAv+1QiosJUcesTWW/pPzVq+WFV
HIC/pNrk0d8NMQ1PZWuMEKHEUihsbfOWY6v2jVhKGNpy9TDcxm2QgZcfEk+1+5H03yROzMg9w6Cq
v2IEbjsHv3aBp9wIfOAp0zo+tX5HAPnB9p8clVQWXXM5V3HUJCDO3r/JzjNjII+yGiYWmrCH95Zb
R1xY3f7SmLlP8wVbCfNaAfDCGSGGNrjFwjifgVHVOq2rXgDSBY1cEiDmH+euVg/GF/lBYbmGGdRA
BM6WmDTzGeHnY79kT7K0GP5XCgIa16a5vOxmZkeAC+JQ3gQsFhpZX9eDvWJfM80umZEKOlFnFEKW
QFlAGqD8sXW2TZ8Y6CFhqbkobtp29xuycMeU2Ba8z5vRNe5t0YtpL0p8zzYuTd9Pwea1Oua3EtC2
VdV8veFlDzX/t/H6QxF+JHh70qaemvDsoiR7ThyG/oIKjW7+n0/KrQuU2Mnn4h0xLh0q3/4Z1NeI
3U/5YLHAk7GO0QpOMs4rPVvNcSpYXaT8uzQHqS6YRQu19i21fSdUvB7jMkw9YxES7eWwOEhqXlDt
g1cXcdKKo0KiwsnsFISHZ7sAJES/lNzLeW/GDToNS/wVCgFfTjrxvBRSRqgTtg/yxYooMPcxwIrD
eK4PSv6n26RPShLLG+pLFPVHkfNofIBNECsjFcuBRb1vysDbbUyh95JTK4RsdcXf4Hr0P7KXGyCn
pyg02KAUlUX73A51MXMJG55EMtvb7sw3zTqOnS0UTaTcVCKrubZJDTSpgmwlfuA7Mwvvt7exazh5
cdkT0KDxEucbjfqASzy4hgjyNtyZLtuWyPbQIiGziOmX9BOInnDgolZ/lvbLHxwwvgUyZj2Vn2fv
E+NYjSFLvkoGouBMiNiWSrIsg5JjUiiIvcQh1RSXph5BFhNmCEJFfHy/q2eC/6qgqLo5YGeuQgxo
nV4Kl/aFF/HWvO+NnsjzSp8cHGGTs1sjLC13T0Q/WmtezRMHaC6iT4ZXQ/6kx+q9MyPYjqszJZm2
pmG+mNxkaViv/N3cKgNI62lLKmhduXnd7K/jDsfQGe+CGTRAOmmoR7vy0Vbi2Wdv8QG4F8FnRqV2
UeMAhjsdrnQnJeWesh4q1/yBKLHD03ruHTvBwbwuRmGR1Cs8CkW0lAFDE23UEna017NeqehI5CFg
46A6IvJ7pAe72dzDap0kz6sVtJz+cKV8L3vPp0syVPVm/GOWvNOwewid1RmS3PRugpLpuqHbk3GZ
GJ4AMWqr53kbR79g9RcZ4oIMHSUpvZCar1EXEp1Pp0BNzVeVjjNSZddYDySHQu1a7g7xsObFOw1R
pUweIdZx3+xH2ZYfF3XxChqOAXVnIC/+ZEQW262zHwJ9qdS8MZuGy5r25DS5S4on3M64zkHsqk5F
G0913FPicBQ0GZM2Vi5FiQGNZS/1TouEi4TuCmt25EvHfAtnO7UcfneBTrbKpGtBY4zW8Db1KhR7
NWmsEJOb13jWMw4FWPD0JFvjilu8bCoPoXuXq/Xd663torKOpapbR1WKEaeJKutzxZNK/XVwE77T
IlCJQVrygRixwIhUq8EVaXqWQ9mpumyQjIr8b63/0eyr2RxFUfjbiOVsnHYW4Mi8eW/t+G6+lkcH
X/DHVq6M+AdEjLYp/lmJPQYq7g9vC8lZ1Ct3sKe8SHvPyISGjunpjjCd/ZejsCjfxM0V18Jggm6I
jHYqMvS4vWeWccQbSYYnd0EI/EGaug6tpSlwI88GNbhlIwEJwDWureekBU+kZgBLb0v3NzgT6nwm
u8xTXOiNCmz4EwlhPG1rzdxfjxScbkGCUjKoLaa6Ths1QPheBAH8rnkI5NMRNHxeA67SjvaTAUvQ
C8ES1pfDR9B5r1nPW61Kdf5XV7gWIwI4V9gYtTfuh+ipyAxiroZJDaeFY9TVzGNZcRiNv1txuPNP
28HSmawhmzertXA7vPrn9n5r0UpT91RHjKtyEUuXBf1cr3P0QQlSJoXwB65kKsAUMvsRqNDMjyIt
YC5ddqVnG9BPXsBf3YjLc7r8rwn+mhyF/5SoHavWdhXTyY9UD1ziDwgKnC8XSBn19OPoPvIGf63S
LnAv+WHRzPQlmZ47Qh6IDPABuhGh7+My5GwxSQo9sCjaLQDvVrXTVba4EcepIiHzzp8QaiINYmQR
IAvb29q0g0qsbb8mTuuFl7KNIgJArCMvJb1FBWubmsL0AEB0oahKcORacpFCoCgHLo///wQiF7uY
KaU20ir8weIkNUITuDFLSY+NPKrBiE3HsWN/2PjxhAgoBGn+PVCnhaxODbdsVvn4YI7yI3o2sxfG
qVHUDYeexM4C5Fp7fZV6y7zvMAerszyOxwNb63M+9ZfJMG08XuKXhwckPc4ZRMslz/IpCxzKV+uU
1IaHr58hCa9J2oC9WCH7uTfTYVP2OX45l69ob7cBTAe9mdZzJofibInXumv3xw/aZQO6WTXxnC/c
iMFCVITRhT0vS9tez6NAgOERmxYNPI/muLINdw93/nrxAU+/jtM7fx7tdHsJ4ctn58SLmubNiGMR
rjqtUFT6NKw1mWTEPG7oC22ZbaRZpK2NPd9K2NH7/vWg5SxhJgL04uQEEibrICjv8Q09vMD0N+sY
JIpzTR8XsqeCI3jqyUsasXkGXzj7dI3Vbd0MI6G2ewrcErSbmOBFW1BfodkSr5xtZf6pfE17lQr0
Xyb00JZF6OdNS7G7HYo3HVa5F3nEwQZmSqiFh30PLUvVHIRipeUggMdDJWvxZVUr8OJWLLu2QWRs
1G6GONmjC2iH85wKZakuYT80tdU7paVR8u0p548x8xGnFymDBmCUEIaD870Ngkh3g/yEIb5KSmRl
DMVV1vQUuiyxn4KjumBCq7G0BSB0VOx8Cn4BZbmCR1jZcEhfLf+druT7unRO7uY2jPvsbrTB/VUQ
I4txpFh4RA4fjKtL6dQj1o2CRT1oe0qfT/4q19wUUOoD1DTf6mII9bzJwIyi7w+/NInRMILnHWHg
HQNY/ekEXqQexu2VRCcudTQ33YpmdpoywC3Y2ddLYc4utrCM+u1k9Okvv6chrx5dFKYcXbS2wcel
4vSAwCQKkPicrOAeUPVqnbRdjmbGaz2+QmJu9xsUy2X5O0ABxeNyhJKSTTogbDTfFocTWJ8EzlaY
ZKKvvAgni2jgpilZv8pJrXtiFcDSP/6FeRJiaHZ2vpt7Hxm3zZ/+GA1J00MiTW2LyRY9vB982PXz
tFc0zObAaYANANas3ftVbozqLrYkAUi1Xs6ChDLshKY0A9lE/620nMC93cDvQU2d3rAv3aVfTWsc
Q4D5FhqW1Qb7MTaq6Jm0wlI0IFB8xX8sfT8BEU+P9G964qLtKlF/772ZFyXWTrFQtJwHCurXN4+n
HioWZU1EbWDoEMbzW/8FjaK+sSqH2Os+VZnF7EkcnjUzvASZM2SgVig2l6k+2nDkwfRINF+5dqLu
r0FnSTX3qIf/Z7yma5PK/KebDjWMGzIiKkLSjFtfCAlfh0CJAwnvHXoLrfJbFxQGaUh6FyThBntL
l6RBv1aOpmhZOYrlEqL02TNnvfNmzYo4twy5RDp7ohb1Zn41puYr4Uh1q9NlsHZCHftYLBix/D0y
DMCXr19HylGti/NvKqISjMYh3EQseMsb0k0LGUzw29ZokewEKBG47XPvzSqtyoyDSl918ftazQ10
fYydYP/0eCCgSHE9lCSEfJxT5t2gB3OcJvBX0PsDJXIUKZhbLGY2hePTEyOyzXW2L9KzkHVomzpc
HYSD/P5kE8TafO8lmP7wNK4zhtrKaIYrbmrssWcMKyCgzR8rbsu5taDujXJxixcAhHs5zY1SFco6
GXwlVfAcBvLlC4vj32N0rSCFdkrvkVYuyCaKi6NfWTIWRo6YNQPuoRb6fAEOpP/CA/SL5THfRvfo
cElMUrAwupU3krKAXVmYp6dtLRgSlu8CWI+jLsa7y/1MwWkeKhfcaVwkEdGw2eVemUIZoTH6aO3/
396mY3EvvnxwQE7qlKUZ8jqAPkK/xZ8ApCwHMUqUAfn1GYSHn1L3hJzIlp06LOt2myfyavuSK8Ou
L79283ok8FfpUDSMMR6IVFOEiSgZFSdxHUumCO1PaLUYfzF2InYQNBLqww4xxlqxM7tbv+IseffK
FAK5YRZlu5N3dXpUEi+7oqm2jaQ0HZm6Kvc1aARIM+3duUbV5RosCvua3Vr8rZJKDKrGxMzUaHmF
9mAoE2RKyBgZU1RdKLRb+xA0oDRPbrzDc8s2ozThlowRvex2V2+FaaMuNuNiGStXCCw8bItOTGtz
siNJplNPHrjCnTrkZrTVU8w0Syz7n3SN8U8np1pdCctKcKob70sgnruKgO11FpuLI0hpoiBRao9k
cMIynAxic0UItkApKjUA4o4mI9I3a5TCT8/CxZHYclMDGkfxkVgXoibgACZML9dW0dye0z+2rN2Y
5ci7YQ98gRcLvmBn0pOtAfc8ssJfkhYHCcVpLuzPzrxCNt4cK800ah5QkGUtwf4o6/xu+Zf8xGed
ov7KB4Ngp/c+MXhRCJOkIBpHNKeoLIHIfJUpjANAyk1V5U5U2KWGUhZoyt5nEwQuISRF4MTgfgJ1
V6hWv0n0KFIuaTzXWpru5H+XoEvySoHHG9j3G/0gMVjLW8Ii74D1wLwArL7/ejO72k0LRUgzkO1s
IZFpbUf492+0aoY/z6EQxKDRW6ZA2SCOtyjaOi6jtMdEqYcBlU7RH5O409lWtUolHhaGwO5SlGr5
K4TlVZVnT2R6rfFTJyNeAs3y13FM6vv1qhL8wzV3wBWR0I9KsbtZgSnQ+N9kgO29ljboMIaTAWk/
S2pXm30Vlty+7NjGAsJT4JhJg2F8Jyi2dR9WfBsY5ZilUl3tnjnHTTmFibaz01s9ffag/can6mc0
xbdROgf//jJoD1S4qDmQSQ2Igfs+IUOE9LtPU4kIzODu2OtSsTHicUxutntVaJ3kkWuzz718/Z6P
iq12MxabDPc4m6CI7xmzI1ThnUo4wqwdNeFAGtTQ7i7xwxHq6oc6QhzfxlLUO71nLLIVqC6UfK7A
2JYzYhbmrQt6kevl4OKfcDIf6b7mJHOsr4KqvJoQXVENeY0p9GckLLFdsgm9p3/mt1icapDVRMwj
7jidNtDXln/ataQUg4KdapTq2xrQlU+W6i8bXXVIcGAwMDoi9BWgUpnKNU+U9ulwhsZtozfczDQP
Wnaywwj9lPXtsy7+//lg2m8azQpE056zStQmskQyZERNj0GtKy+L1sIW5nq/4Fdrah5OVUmCB/Mn
MURpEOF1mJqxrvY6ZybA7PfYxzn6T3T1HiAu0AatU/Sjs7Kp+PpK1eIgexylmYcPpitAq7XkFbC4
gfY6bGqbDYdZVdbeAykgQ5sqEOIEB/64V7kx/5Kd+4srX3vNeXHG12us+58xLRz3HSdZ2kF/3qAa
DOfRhwHjuP46w42e+0o3/c3ZyZL8Dqm4uGjQDZQ8M6KIREAfLa02uwj+LLifmLX2FRI9OoSFeKrm
7OTfEfhcrqwgtx1LaRs/x/Jg3x23t7Mn517E6ucRMIgtv7/+KZHHxGG+r5WvSb0LkTKNMTs8IFSG
DUwS+NUvYjRquNyT8jVSP0ZsMjZwjDbHrWzypAmHV6eaz2OctYtOGfJsl9ZSSYLgdVSI+utFaRqp
pVacR1t3KSmd+njX41HhhV19YMLMomnYnTEUfvRTz8OADNQ0WkwaRw9zYicFTvO0uY739JOExu2C
cGvuKT1Fe7TdiaBMxUDhKFFcCoi9kukzFRxfxyZZyBDJuSENlK9h04HDcdbxcU7gglP+m1pF1WXe
Ec5Pru34UWC1zi36VtJe7Sun9etOcbDlS63WWAvsSV0zO7B1Nkl0BAZ/o+G5vJ7y0K1iXy/nRQ/0
2HR26ddqrMeD+RLgK1O2iNvOa18mTTSS8vMLFA6WhswGYvzdBJf953WouWiJka4CQ+hyZCNRmqCE
P0+eqGxMTKWXNt6J1trwjSMu/gCpMM0INtZLBq09ws+lMMN8GmXuyzBaKNBoUhd8UwgTH2cL/w3A
UqdTfwLms/S52FmtW1/SemQ5xycydGPwhasEJZHAxJeS8JvqTlzn43JwDL6L31YSjk27iqFZj669
WgKn8by4QWlJDb10b023OOBbuqpjuJJdA355Tj0ruMrRhoTG9Fvc6pn+mLu73pVovKKR0aqks18p
YYT2CRStYwUPMHgRs39AwI0kyWxgjDqTcuEh3V98TQ+0bLZN06T1ZAXMldGW6GYg+cXvAc6PVxJV
AN6V8Bt5VU8MKJaRzF92Q3biJV6SdojM1TOHn/MeWLJmqw3g0l6S0cfi2hNJHCaCSAwdw0UKR8DS
GFJnLpfBzJViRPXRJx5OyKdd5X+Hjq6twTlm2sBlc/WgZ5v8Ih+d2q6MnlS6fHrw/r0lrbY3fFJA
gqOFXBI2HgPsFkwOQMNJjhAfdeQf8vW7S1sv525p3275POJGNOzERgIRvCW0kvniTMhIU0spC8QM
kkLu/Ox4PeD0vp708rjuNTIiHxioimU5ZitxCm+OLN1eqmprzaABCb+AVEQczf5zl5mwClXoRJti
F4LcNgNK6Cbv0DC8/FrJwiaw1BQd4P1b8gXfYLn9Pwy6GLM0hMapK788Prjcjck7paXM60tOXjHU
jQCK6gX1qCKlqeaD2hgWi5onBryCIfRM3Saigc/ECPPk7ckExTOMLJ52LqJNjZhyM2eQ8Zbtn2SK
jwKoG6JM5ONmlnR7T8XnwJH4Vk6+YW3pQJs36K/sTkL3hzJ/sCxCE6W2QfRW/lo3eVGQwz2+YH80
5+4h/IuS4lr/KrvJTiu2yCgHuv0reAvBW9SR6HZutXpQrVuXfwAkB/HDaCdb1fwBPJppx0j5u5m1
ENCGfLPs70KaeGYsX8ak+670ugpP/mTUtpnQpq0c/k6vYGXfLd4wW8C2Begb8dC5tRAU64ADBJTA
ekNgiH3eVtQpPtLvv1qtb3DcBpXQbWZ9ICvWrfxGsFfwHU1svAxdnycKtGrICaE96glTsoCTGiiu
dQCQeSDrJ7v25jDrw4+1zDkA1nN2O/7gaC3yBGC+Rpv+yZfLgXVkFuyeSKbxr4Fs/t/YtF+9+ZuP
2DkOZmw3al4DyuGVdDvlQ7+zR62ixXL0s3IyFRG0s3d67hRWM6NorTj915Tb6b054DrckJRKrD3u
/yfJxrKZt3X3RDQEwM1g3utw4cf6tkhKyVf4XIxGfYSC+uWd260keDh/GG9qHfa2HquTNk9Nr+aZ
aYEpGJUEO7p4OtQyUl6+HVT+SxsXQpe3dcO7hDNC1S49VW7w4xnknzZv7lFBrxp/JjCpx2tGyWht
KrRveVV/JRorYSZ9qVYyYcMzN0gQsfXe4UjidIpaNUsg1dalLNBvcKFDgFNZcuODUnPSUCErvU7H
GJFt0XD7kwS21GVPLJOPDn0fsnkkqhluf8CMnjp2swk72IeWDX6nkLCOA/Mqe/ENXNBcpFtr72ei
CyPvqEuJK74NZRI0TeX7BnF3BwqXHdZTy7O7dEXCO4Xu2kfJnrO1nIOlToChTVIB2/BiNDs9LJXl
UXNQOewOoMa1XnfFMwyB5hlrf0ArFta2lQ3oS+/TBzNOvyvzcc4ZkXlDXCcbrAauM3k/MJCya2WJ
mZ/VD4NIQGN8o3UGmoj936tO5gRUyt3+FQHZgAlksoUWtPQLcqeHbIpyLCtX98y+5w7/vSeY2cTC
y3W8612sfejrCNugrrBF5oq1McJX8KjOBymL9aqRBr1aYxeo3BjOGdq2RiIhQsGrQs+k8cju6lS6
G29ElQgcFlMVO6NuWfzVy/XfvPDwhQOJeL8IoUxmjOHs2IR6bsL+dGsFAh99HM/hLNz/Mu8naZt7
rHAXEnP+yapqW6EKeGdAeNQ8ZEVMPHqgZP9lQ30A+1/1mxyvSQoFJB0W1elWWrcrsCQVgvtbHjuR
sdwQrPK9bb918J1So8NRKiec428IwEvhTPUos/K/IMY0OBKCzcVT0rqNNCarcTu+LUUtX7w64Hpp
jVG7DeVKH5iiH/jnEfrBbvFFnBRbUZqiK+jConwcf1EGEpMTJNNbykw3ol8bfTZCc4ptMf7r8laN
+rhyh+LGz5liAq9gtua1Id2GzyOIEENPY8nYVtHm3jPB5VWnpQWx/qneMSjXzQb0I869pEFWv/qN
EnUb2NFILpfhjPQtkNG05Rn1C5v5DZVnwv3DtfvoB93IQpSH4l43PnmtKDTmB7vC5xSirjp2wDqH
9xeMKRaLHaNt+x6mdSq2WKCbwCulV+80gc0oTXxIMmBXCea52P/KeNhfy3r9G5Kzs2p6+Uxr6xvf
FJnIcqQyUHXvN6xNfY2skqYZmLKP4R7kGTbp5BYAH7e+SSUXo5zt9j0TY3pPExFLPdEVW0HywRfs
iaNvpln9iSWFpCSOpq3lpJo5KxbgTfFFuqddGeJvJg3NYhRtnJqVvqb+4SlFfPf0fLx6JwxYFNDd
h8VHZA0JNALRmrWsZlwYMMMprOApEWMc5rf9OXI0RNkpSZUAfgEA5m3sZG6M0pu75WrKPNR6xBY7
4X/XLtSU4EMQyDYwPWL6fn8/lMyte6fIPluewC4ybFt5SfCtfburB5TJzoM3ZJj5Z6li3v84Dgxm
U1O3Y7ok6QP+AJAXZLGsaEHL7VrcjMlYIHyp0PARSVFgHfSlzueBZFCnphmxdH3v+S0ZZMSAmMkX
4W/K7CVFeFZ6/noZHhoTllkuuexm+CzSgItONcCBxSKOeBf0rEEgqgVgTOXYM+oC/ZqYNEZZq/UZ
sFcuv26FkM4Fz/1zdxoAINb481TvjEjdaRSe8jxkuxLiEAIxCL4xbwjV0B0YyJLeXDH0/AdWuzmg
mANjClqqqVU/FZCh0JaaZJwGIY7eN49d8VnJFaLnLgvGFr/NcaXf/D3OWeqqktUGRBs3I1wbFS7u
Jx7yzepaqtUl8LBkms8q+lIMqKt2eT5rJUaN2MVzIYCUT42pdeOQRlGxW3qqWhlYu5YMV7iyQWst
ChN3QS1fGHdgzit0w2vOnDM8MaK60w8uGYGLSzjOCLLv7f7nb6QqhAoqTE3bfIH7LxwibaVXHJoF
EK4lRwEmdLIaVj9ocIPnKKi7QHQsXR6Xe8toglTwppfQW8Bi5Hp7F8VbUcv0Ay1zmeYTrE4+4Mta
oycjDzvwWiIhdauXZBREsBRWmAce1JbRUmhQsIw/9shFx0mrke8UUbkmZU+C85pdCDKzGbLWJoNN
nCDQlCgUWe+FQQzfkVHl+N8SEkvlN+QnRhRkFPhQWTmAJw6HSJ+QiD65+Bpgda/4MbLK2g+1l1Ll
deyiKItAI88ni071y+42Z2lNV+b9zmL5O26G2WD/6XiNqLBjtITXAuIpI6wHxuSCfnEnBX+hOmN5
GRcVSatNv+bVaxF3TH1qrU4+Nx3JXb7i4LqZwy3v6M4WSxutJb+7PWhdj0oDm8XGP4caBRBgctpq
n0fDhhHbPEbX/z5I4gW8Kn9V0M5OypkqRSlPLT3ARTfh/D7BZN1Xb6CY462/ie99vvqDdc07VKb1
d2MPLB+OuFd6ArvaweEM463cXcwajZsVbU08LJN22GDGo6I5YyDygOyQSm59jIa/Zkaf2VHGXyjW
ZouLJGSeMQ7gPCqnYsjlMuZx/vWyPALIpsQT7gJLaagwETPK7/07OQa4VgLbeufebxO1KQmDZ/6/
t85/NWtP7V64gGDXxtV/L385/TccNeImDY7EWMI+wt6ZcJRF+wCK1EIRo+DRvw2e8pZvo0b+JeOx
hSp6KbL2ESS78e/vkWAKLfYdyv1a4nzwvK+7pCY7e/YnaA/DW2HCOgdRDefm5/CVsP/H81P5J5ii
YcYEwpwvPV6FZDUmPpKQMGTU3bsogbc7Y/KfKxfSLxCdpifmtJ80Zj3CRDb3hzLEgzi4W933yH7y
+KOiZFUMb+OgMjf1E919RdBg3UMDQZ/Yu+YREvdoXwBxDc2LZlRXjEIBmmnIxknmeKbfYoInYYLm
1Bt3VYmZhhCjZUYZpoRJuQ6pugOl2q6zK2aQo+Jzc6KMxO/SwcKCjggGDIJmtkhgn104swXauY/B
fmYd/4CFJlMOUcNfHMF7mBaa73bbHDH3CgJlEbWkV1CUqD0KUcXKuXH3YGKUpLTz3HFhSYuTAWAa
Nv0ZmJzfk4SaUMaQSQ2GwnO9lx0S6i91o/nspLMV9yhvTxvMBO4Vz1uurzIadHhS0g/x3YUsGUmQ
w1ff4Qf174wbOst+2SnWQFcN1j5Y1hwn5dNT11/rnegTQDZNxRXuwax4DqbjScwm11EVmC8B4AuL
jxcbXEhEcf4frn5rbRx35RGvaVUSEdWxtEhgVDvBTQQ5zzxldpdPm2uKuhTAzlg/6OxHN12/g6Mx
Wp83QL9QmfRqFdc/YtYXJxxrqJ9Ahnu4EW1ZOuhbWLKPnuP63GT34WQxSVwk8gtTCJoxx+uIPVxI
ktZ1EcaDyHrEpVlMd8cJ2YJg3+j+4cgWxb29Wu1scAxTHxj7ZFnCGET55+cUMLHpAhifegjwk0an
xngsdGr+rmpDqXXX8b9HGHWLmdAVecRsCxhiwf3rn8eNC2qfL0ubf+Dt2ETApfcuxwTwr5SXlP+S
0fSQY11Lm0ko6j7ERg/IaunvHbCAk5inktyLW3FLqm2oQZqa2NlUzKfNtBgRwouUk3va7YC2oBlV
RNY2/2WkIiPDL3QahUQKhVjQPwob3XnfjRYiqLNjCasBcE41APaGUDVKgylht9MFNkOuvSdtH/YV
efGKGTILDTTltJkm8TBzadKCN+Bx0EsS80jJuHqjfnBAZQm+Nfw5un9HwRJk4evc99gqQ8sEvB3R
BdlKoi0CinBKfWNoKWotzhzSJTkgEtPd2HTN0HCR48ceS4xQW/K0zthqFF4VzOFoGKoPHwO7okXX
mS/ZKvr4Nq6Kr4cJUkzvwMuf8+Y/10nV/KKDdwOXjaVOUp+D5dLWb9MV5K9pxwebliVcmkWdJl+s
ChlEaEQU+QCjOWygXi62o9EaMtAC1RqRdAeNS3lhcaeDt33hxgT9nth8LVNGgB/AqmLWTibfSJHO
Bq192p0W5srcQVl/z119IzGqDJpIQJwK3jh0KhOtr+/Nye92/06p+rIksV08vCWRF03q7IpkeNDs
1zdtrcVzDsky2o0Q8a9PHPSFiIFZJkChKJKq4q4xH+ITryxRzyC4lA6XiUjH5C4eHGyE+4eqJwh4
2+4F4icFOqQJ4fXehD7q0Qzxott5ASmu4qwBCtJaTTnNqEdp0+fX0lWouotQBC3rtxuD5GZKxAiV
yztm4V0+0qpxXbjvlS/dKn5c6rQHqZfb7zHsuSwY0+egCoBXCEKSSW1SSFn6MaF4+7OmarNciSFA
r9f8/87YdMftf0+SsC5mPO07Jjy5qgqUu6LtEPmFd+jg2aYiDWXweI7PCcm9oVrOCRwaxq+14yYP
JzSHr89TUNUBial8M+BaroCv6yggS4ag1RmV8axAeBdQ27wa5xIUBRsMeVniyzuFNANgP1Lpa2nD
NJ6eKpXHsWTq6h50+HxlyEZ0woi95NP/s0e2rQXcnM8qHr0z0kuspyb868iWvZcMdVyC0cMQq2FD
KeE+2eZQa5wdtjHbAJozKGToSClQKs2Fq689+VAVW02tQWOkz+wHCqjJ1fe+A2AuKRV1N+rO9KWS
vrfeqSj3EUN5/E4uoYEMNbmWYbxpQ8lQ+pJ/7NwPwmhKWDGmNFKohisOjs/MVufoyuLmSi5VikiD
DeaFnS8JKXRRdr+Sc9pPO3nT2HBY3chLnu1+tI4YIwfxqswFF/d49DpE48YRoQRisGS72+WqAzZH
ugK3HSJ7Ign9l5WZn54QYuF3w7AvWaCAUSF/wpccIqGbYF9XZR91Nx0Tp5627YYgcmGEK6TET0BV
RjOCFCTKVg1UlFfd1xqHLeYH3s0miaa+m+wKfRATkA9dO3lrWfYroLz6yjjsIv+MApAEhU9mlK28
+/pvdKSa/ekRbmFxb5c0GHWBYUe12AYFHXhMHAscJWJuPJPnd9BZw/iBJb+XdEKJQ/kf1t7rE49A
NfyYvkwPl+GfLWjkspKyFxqsf4WbQj3MV5yujwCjlDK6du0HrmU+5VdHX3ssmB0wBUlSjbo+cjFW
h4j+KEFj2o9/31A5zXUmE6XkQ7nI7nZtO384ke4Fi/9t89WCJpkoeyStqEAsOHMFwpC1IhsxdQCW
BHG4VuHutml8iGTmbQTt72q4GUsWzYHg75uCcdFLOxkAwzK6ON9lneTq2WZFmxyhWBW/eQFgypw1
1rVL77t9/tpQJTf71pImgQICwtmlnQ8dlwipImEwatSP2Yso7YoKS4n9tTqa8jkURfgdDqJKK2j5
Wyje9hAsseuXF/I5HtkNZNnx+fMmcVaxVDKexDFnHdo6tUxVsgQdSyyEQbJdngfwTpTzlqjOAJhy
iqnWaundMNGu46uzwV6RgfIIVlR+8r88sLPo24+7KWM6Fn7jl5ri0kZOsB6+OlLuk7MckbsKJOma
ZLZMSawW0RAUqD2cmrFHTwdpR0XWubFlgf3z79fmAC6lvAQLzbZ8wQREp0oBVAwITsDmbmpDutDU
HKiAlURt8QY4JmXvoiKsAlgvtwhegr+7E9gyNIfgXitr6popEAalCgNRJeJgCmzkFARRfl+ywe4v
4EXtv62ZQeSATpXyt7Z85TYK4IWyoSVrxAbcqhbPJFmjZ3FK0hMzlz4HfO+NEKYH7lU4q4utVcSQ
OerqE14D+ASEbnqoJF+/SORCVvux1VcDsDTERneaVa2m4KtIz/D18KG5pMmSEqgB5c7kSAVsYLYf
jB9RTatL82BnKAB7ODiKIiAUpZQH5eAt0N4R8tKWWSl4cyp0hs2DlscnzNNTNYwAPQHmok8zJ15i
1Q9CCPCpcX9d8wNK5rC4eHEAqiI8tYU7dXnSQoa+YIltvBrDIgEIjxfY2v+QVmeDRtXuJfU3FysL
81OCRdAYP937txF9ip/NJkQVyWhTDROWjNSIDgNxvfg+jO1+LoT8BTOops7bCtQFZCjRb9/xUyaJ
AMhkfvfXQ2u9wLrzvzayTnj2WpLiKusoOgMflVyVGsKP5+FNCt/JpXRR58th+et9hFoYr6sHdKJb
AeomLoxk7TTKzZsN3fq3/v3crcgaQYVLIf2DC1xAtzoLgfxyDyQtB8yMlzcp9T46SKwGHSWhUp2o
AizpwT/ibnFXb/v6AojB/WfYOR4uLafvOwMyNHuE1s3+l31ajO2RV6H09KTdz89b9LMJDV4VdhEU
+nZgpfma5Ulaan4YoSFTG2JPth2wxzIMNWTItx3iF6h8ceByNjaMEN48pdBdAzYTlKbdlyiR/s48
Sps6dFu5PDbqT8m673pSkZhN+vorK2TniGac+l1rx1ZYZrP/WDFxfvVfmC1gCOHDEjm2HsGqZgrK
NYmEdf1VHUWvi7tc4LANNIN7zWNGqs5uThyJOEt9v/gobU7fCsplaWm6zImz2KfpSr7cYNY7exo2
8JJ44H+SeWll5BSPtiaiBiwDBhT1EugNYWbIn0OPDB1SSvgeAsDnqfW804LKQ++S+hchnsrYVd9a
hofj/dqfEvByYrjCb/DcHPH8f0NRTgIWtCy0CYHtCAJnmxcCrOWaVVlDJEgupT+eR/1l5ZmJ0Jak
5xXH0+pN5elBOddqnjfGhGH1GzLwNlqBk5oYm00mS5+7pILN9+pnFVVpvtaPbztLkt0m/cq6Gqwl
vdqmAjecBGAn4wPO6qP5QNp14bxb1tYVNRNTFey7ehrgiX2r9nXzhEPEB3B7NZTnSXzk5kKPWAfZ
kLAuHtnRiFy+zvvawtnHXl3x07TUKe/THe69dTewg+2Q+FOvk4RBjHY3//9EynsiVO1sjHstlJaE
b+bODOFdgtQeQJEYplkkUx+xxO91QL4ZDCNg9u0bpDhcMIwHcK9zr5VWG328GUoRAkDRQkM5+ZE8
2gaf/TmUug3kiBKBxSYijrFoxNLJ93TF9q35CQmWRwqwQJMdV1a6kstNVo6+k81C7+24oN2ijlnr
0xlezVmftiMnYyRt5wJdG0VMhuiHZPL7CfImPwZijtucSjRutBXPlIwZKMezPUGXGULY9jm1p05H
CAx2dYo0IWWFae0le7GVFdYgy8MBoPArnAlBjWpCGOFg6Sqf8JtInfDuWCYFa6UvWuQPJRMrGvsW
hWZ55axdswdYfQhp5I6CRivjxW0LJF9buTbB+RYU/cZ/k/ZmkLSDZ8lAijqfoAXMNilD7o8khWpJ
nUp5rrLYuUqNqcmLnNOdmKefQy24mSkhBi2HBK5FMpg0H3BWcKCwu4l/l7QWYqikluxozFkWP6Ax
UMVqD1yEOU2t0DyO8HngKhKTII2YB5af1byxPTTV2a7bpdfnSdXxbAAFfH7RJ4CDXPzRTAf87tvO
L2Y8KnEVdPse1sizUI1n6zPQVdOMjWFQC+kjOaOwhXG6tnUnUPorsYTP3lOvLvrDX2u2iadp5ffQ
sJPxVkkTrEQnji4EQlVSh6Wp1LZp6n88gL48g1HIKVRcoBywDPnrpDkwfw0PiWi9LO7WKI5y73WP
rHKN0MLUbHjEBdW0tnuO6+4Jdh2S8H7HoAnqhUquZ21W4K1/+Sfs9Qyb+KjzeJDU0TyfsEmuJaGn
WlvNNJR3pXTIWJ9p1cwPrYgoDSKALE0XJpxX4Sx72CapsEbQCwdOvFOBoX6EfcuGewUpP2Z87xze
NBsDKGjT0BOzL0QS6H9GnCzg0n8X/Zs3w6EHcJK8KvivGeYPor6h9NgD1TX4AqamDgs89C01eNe0
eL+ArMKqJrYyUUH+XMOhQEinayFhI8LHIpdZfvS3d4TvwRUSsrhmxLs7VGNtIVrYMvtqXZAAZM4z
xg+saQNlh8Ec6A+jhWAW5v2r6MpxU8fnDGdZ9IwFwrkjKpoPkuij/ONmV7nae2fgzsaEXwXXWayU
oCqCkHmo6WLq6ocDFvqMTfqjetRANyx5kQ87VCN8+pSvOKuiSf4z0qMFeunzCM6zY0A399THfycL
raE07iAKF6bTai+MSbkj1SsQEqT2tf++3LP0THeG5w3TiIvBWQtpDIkUYyWkfDye6KFdigkYSSHO
LOhiHUTJQIZ5ORG/fDVjTBcmWH+hcmLwsedDKyqnUAYYTWV5HcstLkFYq/H92NqyQx7wX1vkpdHv
VOTD69oZhezgyUxi2GPPinOmzs0IbEkVtno767M9QxdDRlFsXdk2qBtXu6GT2kFCKYNMVD0LJi5A
g2egTX5CCyhINWJpNtWEjnOrG0WzrxSWhckAIcBTtmQNds2TtYNdnpGNajoZo+QeISABIwaONHGC
3GbbFxVmRtIGSxV5FnGPOHFyzy8q+1AUvBXc1Dhh7PjPdcAZzmOTJJj41RVOw2GkiF5hFnDgSaJ0
IJo50aVR+nQjw06kHx/QPA1axqAjKKcpIdcUf4FhijO+zfbn0h+/nWhgaKvqebQl+5mSLlqfyxQk
kMYTKY4/4EPJ9oeqgSc4tsO2wW6diFIPDG3QI2nGRwdd8NW26cQHxmeaqluzaLognDKlhdtShlXR
OSHLUxKIQ8g4LgvZIZKa0gcAt90oqWV4/tMcB2zpaayG3K0BXn1xcS1mt65rlJGFeeS8YaDJvgsz
pYO5bDjXd9VXlVV40Wk0f8CPDPpS+44KML60Vu5sXC6CrLaW2BEYJ6xqNjL6kGz1S0dWe9wplABl
GCoRoFxaP/n9/QS9mdD47N+PK0VWhjI73c6cbMiD+3x8xHjceXQI3rQN3BkKQQonviq3l04SUGzR
GrhrEeh8G+aikSdIQaNYI1pf4kySjE4t1LGpWNZI/L4kgSHXzM1frpd/kUPn+wQGBWGmAgwNo7b+
ii1mwlbNgOneVmariHqdoiPVwq/VmSvZ6CCeaHzkKJwU9hO6/zOZQDuqHGmFFUiHONKkFo4/O/FW
rZMciPqBpQFOiB/dRwxDp9v5Thy1wPc+1TxfnT02tbnRygG+MmCb8sBYVYqaiSxqWOuytcCljB9T
QR/M0gVRwBFtiO+Ndoexmf++gTEHfWKCHzpdyCY7K5e9+VvJmeOnPVxvmM5T75CcGXQIvKqLemF0
tsoFZ/5M+xncUy655MY5iSJu5ngThNj4eNWVHx5OC/5lIq+gb9ivV0kE/F58EIDLHXFS/yb1mvF+
/CDSSJmWCC4y3Y9MIzHhJCvATr+70+HkN20hYNdYEf3OYUBGyI/lA+AWtKYc/wBAgm4H07XE7Zh8
TX0+vRSmFAbqpVylhapVdNlVUpzMDnisNpfudthPCbCeIFCRkhWPEiEnXpR69pCzKNcLYJ5XFiMh
Vgwszjzh/s7xOGqJWso3MEnQrbFHJ2k7CoX32UMdJeu+GFPOyFWCAvlnloufRLCrNdA3GfxUUNlY
e261Wr04n1ayie65CXiVKMUIUOl/YJvUgx8loV9WwhmYnDujHcD002bbyQPvEOWjMizrHsyWB3EN
FVMUHbhNuX5Pc5dmNGOp918ZxO/Xb6PzgGZJ0ZL6s8Uith6IOz154/IpjmKarSDkfu6uW5I/Xs1v
kepk3XnClp68tjqHp+YVdJJSjWbNDoNKJlQ2bBVDSU6T20rI3VnnDb37Gzxp6wCNBEOcDZTEAAIM
2177EmeNW1f9wvaLmJNiJcPt3V8sUfTDSiW6ZUOoPRPZKkrAK5m5xbbonJ15oxafda/D8+ckNzT/
Hlszcr3AKz48ShQc0s3itQkehstKbO5oW5v2Ht7gEHCYU5KUVrA4nQAr85+bBK3uHObIXKqE0hPf
NgkosAEO8CEWslGFOC6vXkPmr6wa+6UVTNWP21x6rxq5iLj9vIJZOIm/L+Axqgcf2e4M/s8U/efy
XWrnQLH3IB2da0hmHPuGfqISnvDXfLfSxDjrfcoL3hCU+spm3trkYjMP8glMOcPh/cx34LGPjWxK
88cGdhQJJbH9sSbVSh5tGXquT4Tj4/DRvwBfNsgdiLx75KZoeEjL40kYIAoRklrn4CuOo7grbJqT
1oPujAeIvSCjvuARcMd2/P3GkB8mjRYmJ25cIv24CzB0UQ3+3S1w0dWO0Z4oZHqOD6goxH0c1LD5
Mjg0FTacJa/+M7Vv9YLrOhE/vOfMkTblOumArrSdER/XdSfGieFceduD/BDVQ6DGKCwk/EbbA9em
HEbWKfl8nAo5q2cy5nj7ZzmSa9yi68S8DI+5L4l1TQ+hN+gsHxDYfEh+iQHdxcDNlmxxdGjngqXf
SlngHetCa8XWFRQsbFQQy+2KqT8/yr5bhGfs6fSotDCp6rhi0d6o8rHZEw7fh1SPY+UU1p9QSQH2
gYDB17XX+AgXMLFOwfVVdpRzvzOkXtBJAZp8RyF5OYJ2KxBe5HRISaqyrMOf24iUeTMoMVuff3S2
ngEu/Qfb5OgRinkDl8fth369hj3IOe8j+et3/8b6S39x0RdfKC4y0qAQz4UasV0Wvhmmgo47O6/t
69VCqCvnpTArC749GCkoBgYj9hYxb1IsRe9FuZlH5pmHbYi6ZBjS9EOXnU37/Ax5EfjT5IV4DPYY
AMXDIjtayPpZQRwprB8nbIUghDD6EtlYIvB8DiJODgGsatcNfGc/DRAD2/cXgjLxIB8iBm0pre1O
n3H8aZUvuB/3HZXRa0UzkyHawrY6WjOzFQ2920Ko/PON3hmNzUHGAviAjbRZAMbWjSq02fL8/I0s
2ZQtbiJ/WB0PbKm2rNlalbgM1FVPJGSVVOMzQlORV7XOaUaEXAA5NMKaAY7V/Vh9FOqb5vY2XDe6
G4e30CJv1vUFoicj6Tbmv1SfTlyMIScUC+WSMKKoj4kjem9WQdGNGrznOpOkZ2C4vp/vnDsEQnNi
a6497cd4QMQresC+gI+v+SNjrO2G78dlN69iH/54uODKRYoOE6JM1ssJgpm79kLzkHPwEUvICw9o
pzTbjfsPwyDFxhZSL1Lm9a5wLBHOB/eUY4DKL8/QOiM9fsVs10QpLLgePvuE3T1VOErkH/+dtyYl
UfHN+cO6Rj50C/sBIHcV7GzEg1veR6wT5wKL22goi3GpQN1SHSw3ZXShNAlVJtcsxK6cAnSAPGIv
k0wCmB7dgQ/H2D468McaRFZEQ0J20JyxqbYxKo0rHxrM1IonaPBuhgW8iRxQx1Lyz20H0sfvrZnN
H03cyaj2oaiyTVsB8MF7C8u+FGrwsadTOmBiYRKiHRX+URu9KVAwAScFRMr9zQxYRt2kxfPpvEHt
1i8gBnUNJYqirOtXylWLStxDdxzlEYWKpt9aZaJn2WvChvX01oFWT0Vkm1PWaIdMjQjkLunRKKZ3
nSHpkpGXfUt6KnUGoNIxpnd9AmS+oCr0MkP/fYLu5bAVNn4uwoXEOrnUtONkfcWn8BZp2cXuwWwk
VkPlF4u+DUD4sRcVpzW/ugrifQ9twXGVD64rt5ExhaFtDqPtwbiUtKI0laQ0gz++Y8dr5wLNt9q6
jVmXKntUTFiRQJK2YV0WL7Ni+JwJ8F7MPBTf8GGjntHLxsVcx+T4vIJBaQYHrM3y6JS8FE5iNL32
VwwhvVnQKBUxwOTLnMcKR3DHDmeu02SpcVqDhUICQgu2lmxKKxtndaY+JnhwNL3tGGSXz9S9yRZs
fRv8ZoMjEQYuzcbvZaRrCQS1/i/GXEb8Mo7dMuyhLT1Y/xa2SYTraEagNVPVRQ4iVqS9cQ5j1409
LzkODAeJEoR7E3cBOakNvAKKyFtovLWnlC7iUg3clfyYgpF66u+T2ApMnf2rffumGC72beo18Epp
JWd1zCjIfZqVTn8V1ZkFsNF1X+JASvCAR4gq1nCOdJQSEdKVxYUo4o04F3+ndqbzRsyp83raVYjj
m3e3PZtBWHoATyf3K7jNKi453Llb6t2jHuNOm4tF07SX9TnyeMYhd3Pc9pki0zOL4ZIhZ03mspmD
geXqxaRcqvnvBE4THRJd9N/94EntaDyYY2morDTEnRIQZ1RF/A1s46YUDzaQ3KnPTBicrUv+vgDf
QQQ6kvIWOOK8yNrvJnPebd2Wx47Vsch2xM/+H0ets3LMPmzDe9tgV9wBEPZ1MIPMQma6UhPkMc3O
PZA4UmwxnO7Ysw9pLNSm1OJfjVyYQsbWEs0+mCsYuYDT36uOiLSuyZlrgwoKHVj32/ZtXHVpuF32
ALAlW6lpEsMqsezoYM7espVl9l8SzHVAPfmOmXGk1xxRKNr7dPDIbpB+74JD4yTwKZtRNMmOCqcn
VO4fa2JBBYXe8UI0NrCCOowxzA2xgcI3glJnV/HeIPqK9RWLQsRcVOT+Y3bf0oEtfu3dFWDk357H
OQZNCGiep1LEaVwYBnqnay9J+d1xEDJksiQ9E+fFd797N0MKIA1bk7WF1lEnUbPtmnPkmO9Yl0Ni
s3dK5Gkzls+9wXx/KA5pjI7b3VLuLoARbPYWWQBA2cpwYthRW3KGaMn07R4oYzezZrh6PnvPZWcq
5XrHQBx2q7e4SWKZAEw2tx/Mp6qmutqkLUm4+iZJA+sdJkUbHJFPn7xb2ckqHpfzHeYU4r5QcPps
yM8QWphD4IZUcF9dNg0041XBhe71SJhlxMtd2v+VG7t6YguNyt0J0NsNDt8K+mQXqSazInSeeub5
b2LiK3Dgq6Z9IcvNNClWxuuj3Xc7XySeaO1ipwmIYzOYD6hMuPI5eIMYTvn8UWSmD7l8k99rCY+K
5jKFw1ak/H/tOzNfE0PBBnEel0FV/Xm90exqjhzNDaXTHToaurhdX83n4rDfrlT7joWmqEHPPj7P
0jV0eIo/P2sJUoUAhrUgtbnKEL2/+Ynyp9SVWgLZvq/Kq7QSo+odZpduOVPWxczDtzx5sJVUWV3c
6glet7a1YQXz4PwebVeUtrokmqDLDDYTI9R5tNuOFtXZs55SJHLJQIgNncG7/NNj/3MRuV2GUAq4
h/voGvpBclnMuELTufzzsmvJ7z3YCXfjCrhSt/17pVewVucqu+4uJwo6BH5bIHgbGjyVE7HDa/Nj
i7tN8iGHJR+yJOKtkdewqX3qDeSurBoKANIe2xZ5j8MhKG7Rz42gNP2AuNc6GvBhevcxlSQm0sYY
ZSaHzeDqiZP4kNWb6jGKDPYmQAQWbKDsdjO+DL0GOEeGHuSJSgwoK1Q3cLd4Ro5YhdJmuS+DAJF/
JWe71iFfga5SUAJ+yXyco8uLK8lWoErfv6Ua/YAXTES2czOQlCI/9xatunbddcX+V39BcHQROV81
fzWsinadNbYsrYcLru/MaXqTLwYEwIX+eAfrKZ1m/SSuWUV/p1VXPN27vu3LOvmvLAj7aGjksYlL
XiW/BPNVppaNPrato9RGWPKs9TxJU0ZCklGyaKF35HDKkyxPR2ypIa4Zr4kTWEwXqQglowl6d2iC
WuNaaZju2DiaN4NArVe9gSJY9HFfTh3jSzIeqHlg0bhbqQErsFcEdRU03JFuW2eOosdKVqSGOuFz
JwLRGPXmzfjsHyLsAuPeczEw/RV8mpDDFzgQFAh0VQLcWfeggtlk03PwVvJiOI68wDqo2bRSduqC
vFm8z+pZZMDcaXZyYbkfWGOVDPA6tFTB7u6mTQ3JWMITB7fyR+vBnLHAgSh5usOYtfKagsVWn7OP
orY58J9PHAcKA3fJ7H0ju1bQWAOGXkXiMbpZQ3YiXTLMcQ9yWlA1aHzq/erFIKN7Q+aqxFbaoTUt
vfTHbBQbvWzr4qaKkyUO/YiDV1F1uQmdx7Gaw69Ld86fdlAgvjxbME09ExGSl7+AYau/0XjA0t0w
RxEJIcF/vSkhNRVZLvtc1dabgC/UqwfypWn6AkQOeqjo5UlCoPf08qNAnlHbAO3zddlsrSwnRukT
qfsPm0kpQzjVda/GBMzsoJLVl/vfpMQdcCrpRElsI7AfW0Mo1aH9CKAZ+X136M15jeblIoQxk8Xp
RHaLNKvyIuWjJzMaRoofZaQJrErHzo/Y6V9vsL6R+Srhrg2v30InE9TM3hQ2IQWC5cBvpXYHMKQN
Nxxar265yP57+JvP6HyP06+7ZodQpLlEv8zTCZghHS0jqOi3805dcICykjLNp01zP9d4OmFqSANr
fJIMHJgvDBn0LTas4QpivRcIfwMBI2Sc/fxmAnlzwLSltw0yFrJXJDExRGY+fUQh9bo2DmntNRW/
t/wypID8OxEZyy3gdPkZvc0NVPpz5Uaf4o0i/ZM1FRQ4uPA+Xf9c50hYq6ofreK5mio8+e+pcBtF
4K4UjYofqam5Ygq3hsnLCPIAdKvKYQXp2OtBNQwWSYeEdGEv6r5Va6QjhVi/hH1yAncobNYFNKs3
8JTpeX3Y4xX08keeFiQC5W2hUmylbbcib3kZo6LmTjhVBRNOOjE5pD0dfj44Y/+x2TnDjD9no7GR
wIXNJhHhGilvKBS+Kc2tQ4pvHZfVefRRqMDHgSGAkDLoBpgfIQ9nJnNVleITRSckxgoRSSDqO5ny
lm/Oz2RQd92IFYe9DbVHbWBuI/9sbsInqE1axvf9h6xeqT964viLf1jfCSk7sWu9IaZXqaV+iXM8
BP2M3x8ieQ9tHNod9pfJlaBCM3qRZz9KdJGoOemwGaKp+UE2j5ob7iqDaznVdOyeoc9YXV8RX8Zp
ro9S3F2EwI7oltER7n2tjObb+vvsiZWY5/zqoJ71bEw5TGuu4BVsn/F7PWQI93SCNohbK5twk9n1
r3+KDXq06JMRViVhjcM0Nk6A/eREl5cVtp3RBqd4esU68Ua+J7aT1r3jKXuSMzvoNIZ0yi+mKlhW
9t/UFXfUmA3DJIXjvDXtCL0e6Oh5L/+kGCYWm8ccw8jNUNljCLsUsRBhZInGdH7hhsMNeYeGWvr7
2C1IcnCq0t9NvEXtmoB2kgtq2XPCRX15GEARIh4JUNIXn4mjBx7ARkdRMNgxctJgYzCRAm2AiSwF
I4H8SzlMZwy0rS1eAqzdE3DMxmX74owWDbQ9KyjEsRnnX5WAn2t4XYgyj3e68IsS/6JcwpSuM57C
HxRVySr1YcSrehHAPMnDBB8fLSd5uW44jAucdchhw1odNKtHpBWHLBOCgDmaUOvZL74bupCWCOAR
ZvjCgpDMsMFOGB8hd5nf1fAUW9v5P7lGtxsNjQ1VYDE033aWb57dw1IhsPlNQWif0/jFSOneIlDh
awBKlVSEcOeK3bsaLR+zg6s1HUX1QRAH0F3F8vXwli+Fdi+97+8TkHzffW/Pg2XiC727XKqVK0fZ
u6MilXiSq9c7WKy/riUzqmB43Z3wDgLsNlRkdz/gxqxKjpGJwaKsmTWHQJEKpX3EqinkeQHJ4Gv1
pM/BUEurAnJKwmwzz3buyoZ5SZJku3WnPaAaXxJqAOmMnXEPp5uTcpudoa7WhMRBtqRIdaj1eQeK
A6ju7hpyWli9oyX4NDPScnf2xlVxtKtkjd7FO6m9JjmW9+vCWGjiWshunNCPgWfNFiiPj9olxfIj
/QSCwp+UsY4vw7ZTkZuI/uq6F5646I1pDeHsBjBCSgWpQEjJdvv+ZaRju/goH7w/aW1IZ8KdQ93E
gGAX8gyu3BM8aAOd0DeaiFi7BBk7DIaBq/tpHauhmmpU2MPK4KL2suD9dPv3/eh/iGLnanH4IiA0
3PxnmahM9i4/26qEoKIulQlIDC+1t8Agzt082iJxBXit7RiCooTvWCivow7FKM0CtSt940DbxN4W
rY6jBkfM+Wgb8ikLoVbH2BdkPTREZq2pDZTh1qyC+Fb4nIu9FH7MEjcE6BHvkk6k5VxrY/CTrNjI
rD/ktgNMw12vir0xzDbNKv4E34waV9eEobIh+FK/lENkwUQsoVBAUDKebfkCgRlYtkN024vECS0Y
nR1QNZDCZSyMKYiIaUR+tobI1zGeSi/ehLgsz8UJ/LfKE3gUVYIsTcHgLEx2R8vJp90huekAq6EO
Rw7Zy+zQohOI4M/bJZCXPVex57XA7rSLjKlCqIUjPAyD8TSqJfVvGpcVynIGg1bWlTOGR1CDL52C
dWoH8dsrhcbXNrLTgg+RJ5ygyx9MIa78Vw1e9DIIsi639mok72Og/vQmIZB++mbcKHQiI2k5GyzX
ekzaSjXz4Mc/xHmd5zpUtBZcaL2vAZldiYaASk79HCAPpErU/0MBhXTqV4G0W2WNzEKSjkZrLdqr
9aL3OpjBTI0VYIYPbWQALeraaBNM60RI8/hvsN0b+DfuOy7IxGp2FB/w/4ok6lwZAWgFUg52T5Ei
4Xptq2FzRUoPVsBTPE48pl17/mtDXNtWozH8sjMG16C70YeRm1PxFe3zsUA8d29kSSdnSNpUg3A3
h5e9UdDg/9IFDqzXPiwRPVmwvzkkYXX0EkYILeHwGXFLTgKV1N+v5bFmrBWgxy85QbN2HCaG41Yw
G5kRAqEsnaQOTPekBPwVPG+gVCw/HZgbfQ+pRL++CVMpdX+IxW0b22CleVSUHn27UZ7tSl8CysfX
79jtd1Ovs2sT3gmBty2aWggARnyWUZn0YP0cfBhks+7ll/PRYBq3gOJqYTNWK3t5TkE0HKJvATsr
XUsGh/+YbcmDCjASGlTCOSYl07Bt95CB/Px3HM8lMCQUaepQLcJD8c7cRY2htCaFe+5dqDmye3hJ
aIFOCYduxDc+QZXGa+UxCgDwGO10SVOXng0GHbIxWOsgMisj/24ZPEs7V97aJ0Yh4byNvYftk7ma
pW6VOrVyvrFKiHuAjnkf+f9hwAmjemXxgUb8wyrHMTH16MDrtG81ugww04EQPXxa9N8EvhZXm/VR
u9DFCrB8SoZTKkaja2qEeTKDoJNgGKcitxX1shAKGfKEt29SP3SSuInKIDKTxhyzWwXNFIz4uw6Y
kiUkLIo0dCNrYJCBNZARy3oYBxfseBDVCInr1yxmw7H3c9ZeCUJH54mQdzoAlNP41RUB6Xq0O3dg
GieZttWVTwXdB5gc3yhsRT9PqprC+s4j7pr5LF49s7FVaHPcvfYooCHHrI596kuNrWxZ02QAHrfh
tpHU9Tvvxl4j+azA529Z2UYC0tm5rt8ReRkWnKNDD2op2AMeekf/+ds6UYqfbe4LFKVAyssDNjPP
vraOhdQFSdRH9CnwQLNyLID0ipeG1S3pWk4X1mhyrxC0ipJFPFQB+Tf4PSlazOJRwPUdgCQVz556
wKH2GPWMUTakBQGM1ZjPSViRAA9Jh3p+PBRlSlTkweGIKT4pSyyW5bevT39uQ6v05QH/RqvZ6R+K
L0UPbGTmg49uC+6mrR8PSSIFhqz6fPoYHLmznOkP6m022TzJzVl/TGDSfocRM6UVXw4b0kMJhRBx
eaR/HRiRPkUey4xckSUePYOdQ8VisqHvtQRpdky+jVpayFFCkmCK7ivzVRQuyDxPwC7biCkF7qEA
IYxpc/Yv/xR3OMup4Q+oC07VdSplCrBT0bx5Zd2fOZULXdEVubudGZWjk6iA7oQ+xH5Fkveuk9ER
Vd4YD6pRUNaoI+AbYVQAqRAZ7P02pvH7J1u6y/5beTeun4iZiiuEY+FcHbcqhzM5ziq0fEkGRx/V
kuzQFnoOndQ78tR6q2jSc2KM5Kllw2BTOLaSvXaT9M6wDD3DxfKadFgH33L+QrgPvbHPpiDNxU99
Y7/e/17uuagZG0OuOUc9Ptp7WEpqB7uxpLP56QicjxCUhm5yFNDEcHn79UjjcGhyHHZAz3uqaycC
fDGK5CH4gE+42zt91UE7Okr68327LdqU2Y+U17By0pPHXD5N6nGZv19osjwGteiBmEkQogIiJYEY
usymEF+pvRoBS4q7T82E+RkChxiieW5JbeWX2mSQOXcq1fjkZ84Uhr/l5YAsZkDCFUu2ch2gaoi6
cl6d0C7Lr+7834rPYiOCg+q2AeABXrGroaCdhEzCT0PN+kKibVGTMY6x7UmW5EGdsNVvj564UECS
i1haqHiWtL2pQYhcIFON8/cGVg6YalzaxQZf6qKs4q08r080Rra5ve5Zkx1aUgLbUKUMdtBjk8pA
hbqduHG+6Jr8mNiMumTOZ8gntu3fQt7zZMPnvXO9uJQeTGamXyQY+Az9bDYeAueJ5ywpQqyKCIGB
d8RcM5LkG3oMhNv0cJFvlGwNPrLAdRvqJnytoY7p8AvGXMs1Y+GeHjb/l0IgUERKlD13C8flZaq0
oSx/ZA/FE0FR9R1VspBckBrSnkVe/VzAoofST2FHnfmK7fKxtZjAFhQTZtOI8CUtmKk3eIBO9NVm
16II2tUDDginqzsSB9tcK0Amr8LON/B/MePtBCt7CuJO8bwPalBAyUVni3lkdFyojS5MAD33gs92
vFbC/Zt2UBhJmGXNBVk/ZpA6HXlFXS7OkySDSLkm3oWaaD5uW/Oi5CwFSKCg48CtUkxCs6dzpx05
moTl/KnFSHOtgqi9kqpmjnkBz7O49pWDlOx4eBmzgpXiWBRbhue4FwVjS06o51v+Q0EQ/pH2Ul7Z
KD/wUUyDT0v2GRFJOqGSwwCeJzY20aN6V9xg1PMtO4I+EiTJhBWRj2Hv0N57I3MF4dCkYU+Pl7oF
NUbsxa9XxjTr68fpxD7WGgdA0s2wqGbS7D62+jCjyzqTpIgZBUORiDZT70kCNXOPBHYRRi5VrNAW
Ghn3t8CJzAarhEWwQxvA1+7gbRIVSJ/Jc84gMDXRorbcWoHiUAa8Ct4I02kK3uXH8yM44wXuLyve
ols4LpwW56Zq6sNNdmfxmkT0M3DtiHAkSQ+930YkEaAqHhX3trMWgMv7GryOFj+dQ7Yc2ipWqrK6
K9fUwhCK603CI7E7cGXL0RCdgbqrgynCQXfpAKwjs84ztej3fLKIY9t+ZTRZ+m94dVbXok2yD6sv
OAPUxvaVH/Ych/wk8buYW8A4OLz3ja15ZLY0OtpUYGUP1iav56t23g0sIjKpwVyombhrEH8WM827
l9iIh5aSdHKJCchL9ceRwrWwnuyD/EFZ3EQj95F/LE9fxvQVZ6xl5vsEKkVGQJaULJskGf+Fsi5f
jThv4j+oh0jGlVQA4hUNZ2bcB4hz28i5MQM0K7X5oBwrnjsQVyPAhEwyMzxMqeZ6BhvJv2rqL1uJ
4mrObx6Qfyrm0ZQW+KoGcO2s9BPOZeGt72NVtwCUXgOXYFo223WN2kYaxMlQcgtXHm71y16MN0+N
rnsWm4beDMTfOEc2m1eIUGQH2tXGmqoB74uWBKz3Y5T1pXrqlNXzyU/AzxgNklXtAiI9htjaPl9x
cDIZlW2OzCjKDR9m/HtMR/LE81oOX93harg85FMbtuopQHNikkarcWBz5YmkBePGr9hLDrz7vMJY
cv/fWrfcoZnPvAsh1AFDTHlToB6xeBw3IMglJbZV9qedClFVPY0o+TPEZkUVWIJ8FCV8cB3tdJ/Z
9g1fVwvk9Q1+H/wd0GawXmzLMiXqnGOYshM/J9/kEZ0pKlL9gCw4axDhXu6NJB8sxtLn8GI8/o6u
l9YYjHp0brmifN8VbGXeqPUnU7BMQTlhss5fsfVGGLMiMal+k0YPu9ZxCfzWtV6vYAkHpX4QQ9UG
9G+M4Dq+MjXx9Dk9oHr9HaqQyxF1Q1XPeNkEF3le3g0xlqai8C97R4AGxXiq/u7Go1EfqjSEyaca
4IGUz6wpPeGFAXyVgTdth2vQb4K1ZnWKZd6EgxGhI0W5TcEoEJV8RkmVC5tm8VtpNMOHxPhLw/LZ
bYy1gZSiwWBgxBdUvKVYNKjBpqzRmmNZvJwgH4GztUXZdyVq8p5ryHDA9gWFTvlZDC37pWCSmIpy
P1VuvKpHNIqvQUYX5tfbrfYMpifEUYY0sf0hjFpYCLb4qdkS60QX8Z/HXNB1o2CXTf+PMFvMfLD7
VZeX6lXSWUiOTykhh/YJevFEb3Fm0wCoBQI+MI9+9FfGSnpcyOvZDP8UrmgJDWLC4tcz22JHim2E
VtxZ6ZKPN1yEm54XIqbDRyBBgiYk/aHon9r8uWKkr53ppxX2BSlj+7FVq2lGWlZMtkiJtIDT2rwd
fSYw9CQtTldws6TiBRAAYe8JSI/LLul1f+VvwsbBHGHoLGd0MQderiTyGeBBZ/Q7CHpdTEnXs0YQ
NI0RL8CoUrna9RZtq2wnNmDIUzlNbzJmWan6h1TW42J1l1sF3SQENFKu95KUfkN6TnzTgkKo7dDn
ZLLyDZ81MAPw3lJ0s+aD+MGjN/FPCCybLuEwqqhmfyOnWOBJZX0ZEhjqBMDIF/SZyrnK1h8dnxZB
CeC1KTtpWSi0c8SqRWY+EJL0yq+lUJq895jn5FsHSxN7NRUXDwIzB5YUb4kC5dvQ9LR7qnEGmVLJ
b/aYeXidrcP5WqxPU8dGRZpxT5bngZoYm9ZjA4vfW5TvX7n2ECLRZsuDdz0GJmXYwhC4ScdnjbF+
s6zlZ1hfzIdKwI713fdhrcF/IlDR05u7dSQ+WTckN0SdMHD7BV6hic93jVUuAtwsEJF8Mrf4AXNf
K7Ey7vNn2XmPWGpZtvtyXhQmMJxslMk8aNAeGXom8f81HTVrSWoJRVrLfGNx2r8uz1+5r+j9lgst
lct5OwMAIwFLakcSxn5CXx8HJWw0Cr3ZYHndWGhnvKmSDpXriF9AkQA5n9esNjkXI1OUjZjkm8VG
t/lwT7AAgb+ePOCTyKJsFt8UwLBS+zkw+TzlugHNB4XmPp5/rdHLYUXEEdzNlzxVJlYlQI58NwM2
7mKlg3rsn4cicKjMmrxixboyhHmoNhHLLioPTqML7QkGZ7cBYh6fmdtIJ8/s0dX5DplGUO2EfOB4
LsfgSDkFsEgVhze+NYvVyYqDD35lBlf1dU3K1FXNuok5TnFjcTZt54Msf/xM/fQ2VogDH0ng45BE
DR5XFcEsNd9OjgqgIb1zn0PuAQchvacUzZpvFt6s7FY/sGt+Iry5+ywgsM+kz+t9PVq7FnSqtwft
u/9RIRS7ffgFI+aJksdiS4pYwfP540b1sNxzpnSvFgU//JCavo/eAegB0uR4XM3c6aF4SyYMwzWD
aXTJt5OKATZjMpuU1Y3vgi4FhVxG2sq+HgCzmfOdsJ3GSO6oIxgZz8/IjpZEMJrc1XVQYRZkKeLW
HfDt3/l13csbefjAOHpYxA5EkaYsLJxc0ztPTmUrydqv9hfVoS7Kj9ZfQrS+1is6fRNgOFmdg1NB
zyX7+ltOGFLPpxfSgAGFTmMhGYqzzI+q+SWrgAIny8geqYmLQ0HxVZDBA6paSU9P2Y/wrZNfzVuN
2TpdscD+1clbOlSRUrTb4fh436ijMPu1qq7VPoKKgtNjGZwgPoxmZQbVdUB4NmSoDicuNmYNFR0Z
xreX7sEZ8RAqsPf4wMgYMMF7uR2Yl9QcWkdUyD+USEL/q+QzmuUKyM0vKf5Dd9ezHPRTY5o+Rw59
qTTOyeMOLttxeUdFRMv3T/A4VuY85gTMitVp4YkM7K3QbvA/G2OiSZgC7W7t4qUnJMNqu+ZX3JfW
bXkPWRSBZqmPz3CGncuI4rmtLryplrTZBHde8e4oZuw5Goa8P/s3rCbCnJ0YslFTcFB3pPM4cUID
aIxSI8niZYBHi3pqMXn4p35/v/h+uQgHZYZMTTVXOCNE4hp9IIMv7niT67OSk2mj3um1Sj6/hJHo
ZJsJ+AJxfTT3/gMZud110Jd7JTp69TNZWzLV/PNarAaasbVuYkCUS8gTjCZJzyd3N2bQRRmoRdXa
0a3WFzi+edefvUtkapS5bZvCj7uuLou4beyRB7qeKo5jwwegJfgaRuJNaRLbvz8xYgHwn4FeAP9g
vY9YU/rbN5Gz9HtcMNdbwoRxK0LFFIyonQFgvir5qTVH75BWj103ZR5bl3WYzMEIDydHPJiqnAdh
7grn/Pa4TdIJKQtaBM191Xki3PG9qY8fe8M/kvSQzBPsj3ZgXK4IRaiyhMhj313ziJtnC6i/biTX
XpITFZABjiEfj6RsvdaDuk3g8eQoOFospRbnL4jOKK6M7V4mTETOgpHZ4rX9nDl7wNrJ62Iwc0qP
pG8NAWHAw9SFfKk31HWGRFTIZOkxuMaTqpWbWu1ukt7MY4qF7n7PyKxUnauGnoPj3d9RlgzEBtoJ
PFwwvR/HPRy737yKiYuf6fRLFDinIdoc/4TzuQCl8xoQf/Ge5WZW76aXuo9r+tVamX0/iX5tnybN
KpqjEIx/6UydnNDey9G9ukTUsTrBHhNX+DEH8HV3Ti4uIHGN8svi6S7ndr7ejdlK+a/RoUzXhziD
zWE5HYs+RvSE9G7JfMCN9MPCVHhGgyiz/77ooDaPo2mDGS2bpUhtPbwWLDzWJffCMGxGRB7hJ78l
sKcajGn/zwqbiOvxjoXOQ8IzqxfOEI1PoO+49NDXw0I8iz9O+FlHPJUDTGcbhEM0fYHZVoyCxpbL
Ps16EmGZ9kqDHrcB/nNxiUqNVfH1U8w1GtY1yTcFTVFgSY4CHxIktwJjsUc81hpCPD/eKRue7+RT
Up9XVe9hszRlTPJQc2kahPcUxkbVP2tUPu5g3qFaYXNfTlTHA+x1ELzECVM9Xz8IJzszWnve6BP/
n9K26s3uCOOmo6GiTODPddahrbO/GNVhlNYG/wkmXCwV6Y71T4YmiwOp3kAdIxFhNWyDj3AI/OHR
BFJUfslLe8MlQiszh0UZ9Brd3YYoq/yvLM47lvpSzaRn/qbkVcxQiBjlTOz+In55QkZvLB4wf6TO
cHYl/ocI/K0tzSe7ew4wzINt7JOpt+5VvrC4tmvef61xWZckoylXLJ57YDTlXGcem2jv8SfOfo07
LYdGyVw+BO2ulpl7EW+hFEK/y5pGR9HRI0z7XYEG1SAGB8R2d46HhNp9zgY017GPUoTojIzo4K9X
bv4KMozhw1CUR5BWg7DcvBJ0y1jAa8WhkUIgv2FIpGrqLmDRDa8D4YZZRJfjy+czD8Rey65HAIT7
aJexcgWrOfMHGML63qtSHJ7yaL4aOuPy8SCUM6gmhWVmMp5S19B1uqWtt9ShKRVXDCbAYSTGm+9N
0lz1XmMVOMFCz+P6HErzQbVz0JJUz+rYB48zCSySUy6cr4SGUQYxMQdF8IyQjnwviPD6+C3N8F+0
dugb7D9girk8lgbAoacH148BgfLFlIFevfg5jgkMLf8s8HX1hEkkf/18r51IelX/W26u7ND8p7Q7
a7DL+X5gmpALBNynUn3f9gmIKHK0BqLlcJsIIGsMl4OPUAXe0jg+KenYOJuzuKqKIe22WUdO7K54
JVpk4hck2BscFDHzJ5zNMnIaraAgVIDqpIn5eF2MUqTb7hzqIu5lbRC/oohUWXGlbJRIKejS9QaP
Uis2mMb/p+CBbSojWZhJxWXWJK2fgysUZkKnu1usSwzLL659zFFoH2dw7Oja5bisAdUyqgtdxdZR
7WvSwWjvLyrjG8/aGQjpzinozc8wFsUAF80Hphv8ugt+PfNvL1dr3YBDAw/JloF6dC965LEcRU6Y
8qazeJtOqAnEiQC7jySkPfu02OeDlWCQBNK8qABWqcbNKz9eh8UwRkK+b9YaY7lOWQPCjjqRI8nv
aKruchq5d+LsUu0UCRScw0Cnc8QkC1TJbBtn0eoZzE/r6WFJKBV64a6dLNr62dZ8rXlUBxmtimxg
V2/YjtOQsw5LEg5YeOyGHB4XgzmpdeZZRra7FPg8iULCqxDU1CHFairjxlJoMcpWNnu3J4ZWFYpW
6k684e+DZmLHx9sKCtn5TAzSP8Cerm5Q1QrE0Rx52ZmCUjAvZ0KTwJ8w/J1qfx87EWQdhv9deWIk
hHtt2djJRItrrbQC5+agPmTGWUGo6J8ZwXS2U/1CGn5dhC8Ah8xQ9mIUDh2rtjvXy1i0NfLw+hhc
dNmx+ItO3gW2aJPqVY2g0FvbBguWFh57c8ypV4sA8eKxTxQCa/gaCAggqJWh4AHuJFs05mRnnzGV
JwUqzb9dtSR/p3cU+OB7f4OzsiFBhC9SyjfYvTNG3ARBuD9XwnJsHQGcWLTfR4yAdaigSdAgcatP
t9tas6FDGQlbLEYxR9gcwLWloDyK72heEp7PMojP1Bfae6/hJjS0RLDrmSKGcP+3IRtHEAbPJlhl
dl9s3wMi9G2NCQEqV3ZMi5fmMa7iWol9rYucjXTJIv78hZX7pMwy0AOh4rHM+HTKEo1vp3SDVjzq
i5W97LJ30GgU6o2pXADxBnGBIoAQxoFnpfp+xBsSa0tj7DShhr4gaceyWoepd13HHcNqDv+O5/ID
19CiGIIAHFEeTDHrYcnkMdEmMajh/PCj7Na+fivbEpghnzojHuMlsrC0oMyMzVXQjwTA57lA6m/X
2lsE/NImnWV6T7wcXwNnBobyBw7GhdgKwn9g1RxojqpikgvFemK23ZClcujCR105RPmgl6jnVDP3
iKYsrIRDtv3TmGTTkpbgdEHNF4Z/VFeVOuyLf2TEC+y3BEUNzD3pq1OH9u/p07C4MmK6bdTf9jAm
Vf4tVP/r6xDlq0Hr+6ms0/VR27T3XnKTABpl2M32H9ufRDMRnIfEeor3nWx3/dtAlVPhu1+cChiv
c1+TBcfdhq+pgVu0xfSGPdhr8g76Cb+xxMpl9fU+qMSw/iMvXCezwG6YHqQw00Fhprza463IsIka
DjaiONfrSocADsNbMB4eCT0l2I5M96DbgDsxxP9rXNrsSTWGDOTDrTh94ne6LlZTsnVLfq/xklVa
Yaw7UbTpZSyQHxz8B2J0kqo4KjqiGN+kiH707/Z0Iwvt0M8zkheijFrISuJuhs/YMT2G7y8GrFxc
PNIA+EIAIp5diQNJ9J4a7y2oegSoD7gyMb7pCChplb+KLl80TqsI8HvEGf+zyKlsdYB4MnWc/SIy
aWUYAf4s17Q7SfvnPxt2Eqn33whDBacmOYloiW/hYIEPAl4bKzPpIHUQI+dGVwrpoeSbT2JuLsvI
LdeeCzcDwoyAqBlXf9JZf//nfTvDEyMqtlNyTcrs7gLVfbA2z64Wqg0fzrhCWr0W51/QbkDYSrR3
Zfd+RQbgCieXYRHs7Hiv0ktUH1nMNIaA5LxU9J1yqVIlTpqpRED+h2HLDaOabxV47oPYxMcxqB9S
SlR+HH6ZfB94SAW4ZrxJEpBV50RB/79BTwQ+TdX1PFPsuieBI11rkoKhZx5GiWha7wjM9SoPokra
Y2kRqHNwS5Ieh3cHBLsbvK9l8tcL/Bpm9HERvprlalmv56JxdNJwPtnllx/t+BD9FjwmnghMB7iD
WvUN8EOlW0ddS0Gojb1JnL4t9DfBUcj40i2xITFp3DplubGigpy4OWq1XdYDz3ODnBSB8eCCWUyv
BIyeXsaZ564uPKBoXB77+1AJ8hWfmL2BvA/HhKpdkgQFOVSRxW5iNsP8PzVVwhxrL3QLQNjaM0jE
0wV8YfvUsYt7ZAd6yNA0r5Gp0A+eDL6y3Thzp8v+tToCYjTstnTPgQEatCFENHSdV9HRSnjt1RC7
o8czDYvAmlcq+pXLKO/G1Kxxnj0IzqnF6Xat1X2S9XAtddxPBLjHdipYHt3wTsnNMEMNLPHC+5Bn
3gxxuBm1GWfobc0d+EDWEn63pxlM+yXRquLlvMuzhIVhxUt3xR8OAh2H7h8BYzYxgdb1/5lUHl2X
QghFfZ6/xVsI4ogPnVTT+NM7g4jdP+NQMnIqU8A7tUuOezqgjCyb0o0/VnV8S9xU48HB4X/AFjAm
hmg/nd1mz7SxscMI56CDwbxd2/FyOMVdlLhZ89ccYRnEfvhpx6/+CytuX9pHexetC5+w1gkgGUWN
tCq8rEFsA8VWfnRoMGOvneKKbmvrnbaRU81eK6NcYUmo8W9KIxaJSc3/r2ODtOYDev30FTAEbH+E
glKYaneQlqgjMhV/hBIZ5A5jr0AV/GEoTssaE45c5+r9Xm8/bYizPxzaKxl98xZjDUPTQXrOgPj+
3w6ONWvIKJ6wx4V4CdQLYxU8/syJQyF78JHXhcvPAfgW5fwamY40FxgN28/8z02ZsjOJ4w2FNkMH
WCtlFbpC6xV96V45bx5C+WyJ+ZERxlMhFLetFjQwY6FrjZtyvdUeWv6zWihyim8D8691GZl7PHys
H5hJonhqUJgwt6XBJ1/np8UVA8ZL1NHgi/gQHHh6eYrfpH7ywYZPgbTAPIQbHLPuiTcklkxUgjrs
DWhTYHNLVwwcRByeuWYDCCwrhEYshltQi0b8v0qTeDj0JFKBP8CuWFd3//Re4GLENG/dbuB2etdI
4HGlCYHcV2XyIB2RWZxr8qz160LOYSFvkueGZUUoj+mNoxz4ZyLZ1vnSh3Su3CzQHzI26PWlvbTt
hL+O0w3DnB6g55zhwobPTK7p4VAeqBUb4U8bAlGo6JtxLHOdZgX+NObyD5mEL23nJ4sEGbq57F5K
uC4l/+0a3wGCg9vReT4QYfH74qaWIiEgUHv7CzkcQh5cl+g4ZncxsJv5QiCaJD6MW+BwzXK4xNO2
JQTldIvX+UsYGT/MaIKppjRkEDSIBhXPrPZGRljgJBvSg9ywWa0zrsUnx7OpoYouymgUdIcRwKyf
7jKd3ZKOAuVlTcOcLum0CHuaQZdudM5N6LxifrU1aUFozVPb05nGgSNsf92OiJLLTsrllKB/lUGr
kNYPt13tYRzL758DwfzZqql8/ijlotxO2mQgWn2EBgZ2pZdTm/hjwnLXV8SyeHCA8JlEbP374Lv9
CH/EkM2EM5NZcxhjeFEQwQZXfCvbtgfKwivSqspLZwRymrUoIXtg5Tre5/ovNtb1sDdaIB3mab/j
IrxzG9ZHQ98UECkl+ofkzSueBulteYGhVrdviDCC+cQ5FWpSjbJG7x8vhcTZwzrStbbkMqQ8K2Ns
9sChDKPKIvHWggBioF7a8BT7v0WIVuyjgpZ7hPnbrGwudwt+rXcsBCzqDyxeOh5zKTMt5DlpcmZ8
ZH3lAW9wHo9c9aB0I1XJmndYvL6ccrRo7OqHi6iC92JQCatS37EP4SSx/xcFf0xWYK2rT95Vr8vH
LBQkuDv0/qnAMKgeHWC1yQJrQCkc8QiAWqkfaBIvup7YoZMenFT8gx4gzrhvIjpx1K9mwi3k2YCS
+lziJ15USOWi+A2NjzUAuZKJ0l3OfobWlSHt69t+/PIVGgrhLFoGLyY183dburi1Wk19HRQuvHr8
MUvv3oQPwRL28E4Y1MARh8ky2NSTFM2azOhuSPc+kEz3JRgT4WJ4YjH9LCQWSGk7YyTD13Ue/nej
bxxC1zi3st7cpoNJfdE6u8gPi12SieayjqSSkiFEvxwwMy3HkWKGDKn0/sUO1ay9k8dOjG+utBk3
aFDo0mvm4twXLK9q1NyQquwtDzYkVP2nZNvP2Qfp1BxrMo2uzPAaNG9Px5SQgCRIBxE5m+phL03p
ruTx0y4nn1soMISDNetrsdQpmJTf7bdRPbcpIcfmnnjfeEZvqMayJzUDuRpR7I3qVJKfaPgo7ocG
tRDeHbg0ebtOUrQsL481r+mYCihalwIgu8Duwh6fCA0JxWxyRXAOMTDdDGgEpj2Z6n5UT0UOwntw
uPyTgF6Q6ySryABW1UK0MdFz7/P9N/Sxu0fMt7GN/dcEJ61OLc9ltWMrLJn0np8/oHMJVnabZfo+
KK026ygynl7SusPLMg1ulLX1ALlBhVfkYuZIHnBlIz0gsO4yynoIW/LeQryd6R3r6vyKfsO/x8Wd
SfSov/eBBO2Mx4VwS4d9Kt8whwIhHtjX9AT7syIxr3+mgs08vRGPbS6klyxtBV+RGXXYGHNtfUtD
/a1wXbgcsRmI133vuEkw0qUQ2SOBr1wYm5I1DhEfYbh6I96wM0tiuzKhH2ZexNOZ3Nu67F+dHKat
SOVLRBRzrvxDr19HGj3kSa3eBZKnjIlbQw3Ul2hAF14je5EpQroVF0Mr3LHM412mtxwAVsotDQp0
EZFrlVtTT7L5zMHZyTMzy8bm12eubMNYKvhnAAZTYzn5RLwVFKOKvnsk/de+CnOM1Bvo7vnnwXri
/d/+kLlfw33QQm5GUpubSK6CxHvOjzht60Zl3SHmFlCPc4ESB9yfoPdwjjPCkyW5jNlGEhgYrGU4
gd0Hgczym32xJBTpd4sNedI5+3GLwrOutCTVNZYLnp3PEOxZ/yEk6u9nzFtOitRMR5PNW508Ngo0
nY8Xoq7mGo9O4Uir3BRkTr55aIloX/G+0my7kgXiycPGzWq1GsIx0CfEtN1fDU0JjyYeZJpUWLNv
1q4qo/smEICBCIvgbMRg/eRky46xpP+nJIm5joEUXgZclrrlT/vLjz+rUuz1i6JS/JuLyiMX+G4d
O9gc6lAThaLHztfNEmJPek/8j1sOf7UoG+EQzR68eOMEdNLh+vM2g5UGx0IvNcb+7fX8iLr9gFzI
xcOhzHAMgDhb8bsJCrNDy3gVAI91eTx6wum1/zA323gPlPCTx98DBCrnik7DJGZysMZ2r6AWR3Hf
2h1+Bv6RTv6gpjMkXfmfhM1xgYEA/JCGg9q5Oyqcci8IHTvR3PblK87HdFZ+hiOQLzt9to1gCcoZ
nrXzi3eGRISG48iAkZuHXRX+26ph5km0PtU5njKXnlAYGD9h/ESe1KXlhQZvTtB5sGKAuam1feMJ
8DlLdNY1n9L/x3iAn0VedTgReUMqES9LPo/6QDNWgZfcppbXiwUYS3P06Z7umEbbVJJ4a74CpNu4
Wmosmlbs8oJ95GBF60icfH0/4YUjMEfJMBLCQw6OCQzoyH3oR1WjFj22H1yxLL940793ONv8XIW2
XedmLnCWNEVB53ql/HZLVyDYqsTj0uW36YHckYlR527QNHT2Os3rVeK3VLR+JrhVh8Ch4hE6wwrB
6We17Bpm+6BkI7K9hoblsCnjCQsdPXPzrmayCG12cnxGO6jtaaVEdqcTg28flSVSJPI5fIp08+zQ
JxgKfBDSdqf2u8nbEN/1QCZCWra2RYUlMGqGCspp+UI/NcwUMuVzfpYk6yWyY3HGZFnB4bgWe4gs
Ac/zjD8vUpytJK0TaFSqklbNPJFbWKYAv5iEtfDhnjBmbG3cJzfB40NFGRFOg8vRreVB18pYpTDI
TWyntVFIqXhI2DJNc/hzEJjtaIEcnyuQayBK82iF0Tm/fA/0pEzLMKkGBxD9l0tC1D7HHo8G7qon
CyOijIMAIYWe+GC49UX9UXLEi/Hxr7K1Op6vQz2bRclZu4aJ4x8MXDPAoK9r8ptdmw7NRMEmWxg/
hjtDt/9Fl9/aYNHK1E36AF5VoNIpdbh9vpnk44TqHKuEbyht6woadr4b7s3Tw/+9cgi3jLj4FGXm
B7g2b0VffD0lC3teO4Csn6p39Z/CGkopNDrRlFmBegX0nfXyDKAjrTrlE48DJL87YHbnVAsFbm1M
WELVoSEsdEWvnlW3mE904yrQFIm3V/NiWjNiIumQmrMySFq82xUk24eSF3Bnh+8BWLACu1zv7XvE
Z0QMBRtO4xEROSkFGSrTU5uGMCHno/qKYsEjTWccqIvhoZ/vIGZjqkIaKG6iIKmztY/NYdV8Tfqq
1FPgyqWViAzz+NeIaJFY4fmlrNeJeZxzcKbRvVVwo4JTq6ONJYnFen2Ag7iJ7ROuzxlFKvbNASkx
OLBDblJQMC/Ql/ZVNbAcKVQY4u0a/rMaebCkRzVHzlV4aInBPo+nsWiWhYiWgY2zz8XQteTTSDG+
5ocZhLK4m+M9Z80bkFLXm/5iH3KJTWyS9ehKgEQO69gWfyar5xVV/gXfMTTAR+oHqCDAWnI3yR+I
IXkCcbbgNNRG3llTriHkIecmmQ7ACjRaXwApqz+nVdnhe3l/uLtqvbs4Rt/ivTRSCKySDCrUXU2i
8FXsjZZy0uP2+Add89aX7z4JmSb7OtjxuJ6UkPLQmIbr5jpLjRfD+3xAKOeGSgHkJ/dWj6zD8kqn
PPQsWjdndbtYNk48WQywqTkmBWwjl0x2Haxc86vZt4vIOucgs54dYwm6ZTaUFp7Wi3znLQZiDEZX
grMy5/8dQ2lBOYtGA9gE+04IcNtjFgl54KZ/DGDQF5DrQM5c3UUuaTFlmCDHQLb+XaEIcXNjer9/
vOJiDRL3C/v6pFBAlavNu52xHVVZCq/WgNi8STvyZzXozoDG4mLo7FK0+PYaWA8nBifKhWQFC8/T
fuk7r5HA6C4F0LiI5YgasOFBnPG1p5S7a66OdQCLgqmQY7F1ePux8/2hjZqT9o53EO9mD2caDyEB
MHGd/9yxbxbANAJF1b/peWkw6B5bQOpT/HDMHSYrvmMLk2G+jtp/UJQg5H57V1WHI6z+OKpqVvgD
U02UIsVi7laYBO+OUSMmpY5aaBHrucmSpbFfIWQkptrxH661Dad4W9/AaaCqsB2pVJUFSnkJyQM9
WUzQsiI1h9m6dthno6YHtdCK5WSko48RDjK3wqprpEDrzJBP3Oies2n42P265Ovlw9aPKI1Cq4s0
83ow8YDFIKDpAqnrh8bWzHQ5JQhpiWLkMIFioY3aLNLYjEPXLKyAeRDN1cmg2hIf5uwncW+U3Nzf
1eHCtmbD1VEZeN1WlZeDNIyIEUCI8H4SqI4DNe/gbmCHiG2pDMsjRJcQfoZ2+natwcl2q2Q/wSwA
GpGPj+3chvLWQnAnO2eaowgK2/JDSL6AOfj7ob5F7cbrA5BRD0MQvq46KTmTnvjQToZy21H47gPF
9+TU0LVqvsnKhW5TidF++n/UdCVNSIoBIDGhBY39Z17+nrFidy+TKT0AtoQUF2AgMmGhIvsHg2bA
ZvyW2txDyiv3qtk4XFvmfZQCG9VXRA7L7J+9L0mlxDnNR4a+EPJM+r3E66CZFqVD6TXvJJN/rFJE
k1AIYABNRsYo8+xkEYjzz9P/0LKstUjycCPjVkGZoShjpywFqo2J5MPB2iLHb1+Ttcfp5gjgw+9h
S0vgHlv3TlOdGUyMzMPGPzZt64I0I+y+0QH4goAVKgiCfHVMXChaXGxl2YIgPDoc19Q1mlC2VA+2
MwCXDxM7bKHjz3crJVAiYrn3GHg9C1XC/3o/Mf75EqVFVZtx3Z9dEDmvKS+Ixo800dGZtQi8hwWF
Y9HzkeqJF09vlJ8CCbjbbZrVu8LdmQP59qVBAIRH5crAZ3ownvWyAcesqxd39nAZg+VI86lQQwWm
dAGAmZKiL//VDQ9ntpcLMwpdLYVIDtA4P/vDLKTWg+PCHrjnyDR8jxbY0qgn05o9GddRfUtzIXQM
l37a8blSaGt3JHHhwOcu1nJnCOTVQ4aYefo+Hk4eNa6oWDeQSMwOrxU3XnjBOwEn8Glkxd4qK4SQ
ysLCYvMkCWv2MeYXoFUk1JbDbr3sgoV1VCpOcY/cwObPhncG+t4B+SNV76VehYap8OhWH3u+pYM1
HgqZgqfr7kk3xJebM8XHw8ydgYnnKUNFTV8GX/UrrvvktyR90My8jEWaarfwp0gdnoXGE0vDlFUy
EB7RcL0D+PEezi3ak21ykdlp5UqKEFD8p5A/kHTlIjTG2aldp2zB3UhYBgcTjwJaZCi8I/7FP5yt
uS0Ko99LkhjWwstP3AsHtdEpUGhWyTJwjvicvAf4rLVAcEGenr1EJxvnb02Nm66IlKIFzkDHD3ge
UWwafy0XtdCYv6y07XDEVY6Fb6LHK70dLA2eLyuBKx61yR5d1nXL+4R7AhgI+J5XivYTbQ2bmaBT
DiijvZRFqqmISAXUUupTar9Qk86rWtLSlIvWCYv5hJjIAJ6SsTqMRcrG80hP6s7DEjla7LtUcx5E
PnnjNLXOqinKclY0WIF4YuGp8ACD9PQUEcw4f+0d1qfmTM/A61VVhMawsC3iY80CvCGecF4e7xAA
W2V0/9+spnscGZGlbP1/Dp8/Qo5TCL56ihq+kDJeUqVxnWJvIalDOfMyJhwFDamKi9vyUzJHjrpN
v7P02Gl956CPckDdqMYMc4KYoh0SE7DAHgSkBl/Vtxn879FuPGTNIQClTOy9kmZjmGskfp5wqy5p
G5GdtilqA22ptm7QooPWYjDmfMDWNigqplhPko2WqzMapF1mDnaScqFaUhe2Z5FxPJS5yZUb1nT5
VPpPHWrQLsLXWzcGalLmSTL6/9OaEV5L3LLk7Kb07jVkMc5yx1G6TzMCk+vpy3zKmbxFgwaLVmYu
SVpxFOMYsuHEqS6D82e2huOJsG3V6IEE0D+QG4WnSGsQOcL1Q7LD4NuE077Ji7Fs6+HetzyxlDUR
C/XsejP9HpT3r9armyo04VURaozEtlni3fQlXN0UgtcBJz04R93VMqqvVKnt8u7IBjUxW/O644Zs
qWyl2d2RDn1JAkeW5hol6mX1HKtU3mbkavDF+F1VEI5JZOmaFK9fcuU6fZABdNgL+pN8enRAce/0
b+cX0KhGN8XuE0F0WHo/nCnzWsrwsJfgvOPQ/Yyh2QPa3EMt3EjmMgjz7Rwh/ngMcBpAfdHcdU4H
RqEwcDwLKVcp1b9d2eFTwhP1Jafv1KJZsGKQd2GapvhgdFIUIOdHDp37Q2/o9qOhQxIXeoCivnsI
eu3r0HzOqo2F+WIQRs6JTBJA1icE8Oj9lU8TEafjn/ApGYDggtoK+kicH/a9FjqUCuJO4FEyFR7V
QhV6h8YtPZ5ZoOOBRIPkc2Q7VIfPmKe4ERCMot/rEfOw4un7TGV5JkIkaT84nGyQf/iWNG+XkGQ/
AKhWYJINKtEG5UcpR39KOMPSqVPHklnQ82Cyx+IqfbhdftYv3jSL1ohLa2LB/bgQkjfMqZJhcZmU
ULfzRJel3Zn841D5mlO67kinKdVOfhWNzBU9VnLdRyILQLsYIU5hwSWLGdrj2F/cpxG1PuImT/AL
ld50eUEdRwInDpOC6eC9luuaEO+Ff9OsyXrDGbSWt5H0sfdwzlfSL/nlEEW8GCv/xuDy6BRRyhSs
TFmUp2WdPVz09O1I8p/goVYayVwWbATWqyX2s2wM6oOaBsY4FGRAJYt5DAvpjIngCLkeVUY5Hx2w
UasgQqABNyhXQJaxv35jrpQiBlYM/RS6pbhzXJgNlBU/NbTz0n7AORH5tRBFvzITQdfJ6ydA/ZCn
hP8DhuTHZvIBTvMkVLSi+sM8TeRkpcgzF/Er2ZxwFYnTSWjGvVxR064kHUO9T0lbb3M6oCAdfLGh
koD/NmvueBaGa3nU0gByWZpSgzuWfTDupF16fzBGcdjEU59n/pVMW+W30JRSTcBODNgU8RirAbtW
DHyeJRBA4tYtDJK5VPdizsos0adARuZq7/dicJJWNzicc0sAQH/bymZw5CVex6oyVzNVTv67dYwp
hM2PR6l6yPAIsyXAYeKOY+kkSUZD4OIqr0zfH3azAGLkNad7WFhw30FvyB2bXw5SdHYYSw8RdIsu
056MNbcHrD9Cos40hkysJ+J1pAe1Iqt+0ANMbT2HiUo/x/eJkcrPcEsG4fBsinNnYcCmPIb6WRZ8
Y85DrL2050pY+n12uHZ+5i7MzJvXh/3/h6rZt+XSi3rCHUbjHJ/Q6M1H6sSjZ400wribQGZBo+n0
Gg29ZfK9+KoLvSLw7HN8ZoLaxI9VGByOpyCUIYs5SueKHofYXUF7WZNgOACVyEZ7k3T2gD7+Fcl0
q+Gb1vFRUoDdxP4XR0LqxJpRelN1s4nxnU9e0gndxdJVVZqvBwT9X8mLH8X/0Womn/mKPskO3syO
zE2zhuMRwWwmq1WNpJiP5PXLtBt4WN5U7gNlX+MkXdxCvCwQsOPRTxZOHGjAlsKVW4SDmc6kX3jB
XxYQT86GAc9pHN9nWaX0aKvx1gqW/5uiTGihooEy4VwLpe+X6uwAJZRQR0TYVI/i2bi8ibF/5Aps
daCG6ode9VW57clw0eXVfPTr7alHMqk7f4GJyv811iAxsjqB65Bk2T5N52p8XKeiChoiySz+zW8k
RREdLW8SCPi9LgIUXLC6R5Rq9PWQxt27lIUFccymb9z8EZcSo+zUSGTFJ3DMapdplJxJIg+2oqpM
cvY+dqjMXx+M13PMWcHgOd42U9XlyM1XeBrm/mlRHPF/9QXrv+qOuTkkHlpO6KLullS/wXPMGV+q
S0dNdckJmSIan+5pde0AZmGdWJy3Lrd3mtaRJfdxDW1zKFgR3f9sm1WJ06HxU8jn6bnfNwybQLjn
r3TxkviLGQyptxAFNV1M7IjXnV3JGj6IhYO4d9RZOpY8y2k4zzBT1mqhxyGKvmFPdUS0DY+IYgTV
46n1nIz4Q8CrMIjB1/6SUfScrWfTN0wk0jgXtDxUfqOiCDd5mhTc5SZM02y6kRtIjfWvboHdMOWH
54rq4bK/wDdJ5fpb21Lvl2xk29OohEhusYJGee1eMCjC7mOF1rdUd/AKm5LU1r4Uxbk536V9KGLf
EvQea4ThMGT5LfhtHUv/rDgJk4+khmuZN9yZ9MknqowEqORlp+bEjRVBvNNsQQuXscUd04YYYO5i
8PMI1Qk7IdoP+RWJCJNj/KX5CcNTRnfrhpngGRajaC/jCf1CJnVg90Y7tjP34EpC/ROmpNFLAAwX
xuRNX0THXom6tuoqmEW4zB7EFk8sz6mWGUs+6BmFkYmOT8h7BMbMQXZJk9YL7vBuLuABGojXaV8v
h9ZYypKtwgyQdZXYFSh5R2hG88I0BdSBtIYZlQpGlc1YR2SFpYGeQuCAjD3MMXy5AhTvcGgp2mYF
t0bbaIQxGvtewnH1TBUUJY3RVEqBNCoA5YSGtKedyxHDR42yn06g4PAnE0v2bXNkQqztHEj0WB2e
vOTJGUtyjZrgdYAeBQWiFvsArxjSQU8nz6ACT5bA2ZMVdu47Npag/sEUhuR40BqIz+a0nvdUJnMR
lPMZVbT1llCD5rOA9QU/X5ARhPDka9FtUumxiZeMGh5glLfqULrGUK32sbUqK+JcDVjVqYvxyBDq
GwJN4fBIlH66BTR4H/p61YGLskSrpeVlJngM8OJIAeQua+Xkb+DYSGgpe8J9X/LT4VJ+JdZb5v9i
nOLXAvup+zszIDq7Qo5oLbEdkDjP0tZVN4vBwNC0dqkG1mbfOo/RVGF2WLUPT1o3nm0L2KnRdlg8
UxxMAjZHq0SFI/0Lj4E5grfCEzE3jfBzziiZJVb0QUIwtb570rbHhz/13jg/VAoVBiLtSkBEHLHF
uUNnK9xG+Qvf/8bwRCtp+ShDhE4iWyZKjGF69I3kUGl2M6ktpXQzLT17QI86YyXdEFDQvNYzQxUy
Qm3HkIhmozHSMH5LBiGprkh7BrxGlDwZ0otN7HaAa2UVdd3u6vnUNEpY85t6hZrMuo5wEJr+WVbp
0CzqDorHyWTYLhRJLlE6BDwI6SuOUvK5nL1pRcWF7LziPHOoCIXsOqLI45T61m6qxShfe/rokj8/
r1JopZ9x3CbEvJ5T8xVKRqECyKxBptEw8nnMIGs1jYDNHPvoPmKRVELnBBs8NPqp67e6YvS5WBzQ
Jspi0QfZT8paRi5iRyjnNjw0DgDhSJBiGd9clwZyU99Mk09tuBazgojWQkES6vBmlpua72D/DEKh
o96aBA+9bDu8zn1yC3807ONLkrSEtoq0Qk51juK+yk481vjdRxIwDW9wbwDiT8vsOydPUCaGTovs
Qd0V82ySwRnizqwR7N0NYDMTVdgxv9GGgKHml4AeebIAvqn6mztguIShjuZEr8TL0IFqCvfBHDqz
9WcnffPOs2klbYljdkTS7LNxn9ixq1rqVA+fE0LH3P/U2mgoTuDEOB3T0iuPoO7vfYnnKqB9e8tZ
bKibU2jbGUN6U4uH5SvkbwBqyPgDDJkwAmD0Uqcf+anO3p/RwgMD6TeRBIVl1d2YfQaEUDQ/6HQ8
KsLjBH+j4nJ1XIcVbIDc4sw3Mf8QSHJiW4LCJBdXH39n+EYtAQJVFXiPxgC/gNXC9L9h2aMxEezZ
tUZ/HKs+gngpoLgG/YBjK/8IX5qk6ER5VeEr8alktH2WMTBhWRyC4kiuXiHvHHBoiz/wS8G4E1ds
eqvRvSgnVvKJSU80BguIEqoST105wZuT02wd158beew5Y+XR6r1mjxFeIT9eH99oddP4M5bybJ1g
qCvbPY12qdXCZmuHvMKCrHz/lqMQuRQOtr/GZ+97sYE+WKIeV/aenP8yqQ/P0um9zTFzX7k+X7+R
qBR5m2sv1tHdgudWuROmap/ATM6BXjqCP3LeCRN2baapyrgdcxTgPqG/DSKXS8K/uKTRBZ86qrCz
CQJ7Az+FqK0vbLkqZuFjZ7TI6x8TcRU2jVZ2BLPOfyZ5K2HQKTh5vwv6cfgW3hYaREYItC6aqAlj
Xrg8HtsOqxNVNZ1bfk9cNbCXYbLxr7cRpsQ0O+XKi5YbYwLuy1UrYMzTe7XWNXF9fUH5mbHWHCuB
lwp1DvXI8NCun/fsinXgp+xoxEcV43FpDMIjQS6YKJ3N349Kflk+wHxHTtItRQ5aJvrj4w7cMlfN
0sZLA4IU+jdanNAHARq7lz9PKJF4FADHVxzKm/ppRfyMmGQiPVEADz9tL1s9B8jA72ooMb23d2Lk
SfHPRCtDzhu5IZbt5TZBCJcajpvG3us7llkFxUxRbrXacqWhY77WixPwTbhkd2Zj8u4Jh/IWSb9u
+7Z7DkdVApB6J9l/V7jfETP5EQkJ6gwcOB5PbDbR31lVXZNsyogMy5G1aEdE3laD/BIGMxqOzd1l
X+ESKApcpTWeNvsauiSfIfNmzWttU6ubiOOIwAgqjOQ3srrObhalP29MvTRy2GV/GQJT9kCHHpin
cERacUiUOyC5+U6Xa0BfTzaKA2dzzFv1QguF/mNswJmq9GhDDIiYZmrMP4PqkpqWAJyE6OQiOud5
M3HSQPrvjYZVrzrQ+LAFmxPnxIF+IPeJyNHRLxKf5mXMzYGQhGTWtscjiOdaFqpV7ASininDvShA
b144DqM/BR8T5kwqYpTW9YYCGoy7C7IBYxcdYmlOGucYORUP5B7jMKXzAI2/loItEVqZLl15DQG3
Ql8qAqewjbwGe5KRR70JMEkeNH/Bum1biwpVL8E8JyKZMEsANhN2s5CK2Nw8QJLD0zDkQKg1bAGz
s6ATEDDokP5uDBg73uXF3EeLAMM0r5Z+JZuLL39jpvQ+tffEjHQ2/vWtfjbQ0QXGjEEw4urHx/br
KLpH6AxNA6F2R51Yn9dAPbIdGqqoFD3Hf+X0XczbqIYLIqAq6sJquV4hjco88cUrAVW8di1G7WSo
QbBA56y2lJEnZfYOPhVCPfyQJYwlue8bFganpsRfQq+aNi1awwO+BuvsuEVi1Y9Vp4tFSs42bvcb
IWH3PQSkwriF6n+KxYBP4Ko90U+WIKbZRz+Bx4QDnBKY3MR8CQO6kMhiskHK0K/d+tiqFzxBcrHe
8sjS+mNLHfzQAa2+wDMKlC7GfLgMXk/SlS7wNAK4340eRRkCjmPQBGtTWZ3pcD1Kunwzv0/uoWiS
FvfnHAZQYz/C707Uu2pQhhdeTiVBKsjhBuFTcT3hUBiTZl8gKOxIn6Yn2olAzUmu6ZwQoKYSn9QB
67L8WGwig8kVJeKeWo4/NF3bVfE9jWo3NVJZMbPmZabZKv3OoSB/dDnzgq2ldu1qXGTCru2MlKO4
toWRIbUjEVQRu2/KhcTkbmHGQoUabSvRKUFm6cZJt1r22ORDbHP2hhpPoQXvMl3f8S1qn3AQpqfV
U4/D/As4atJwgr/JPLbHCJBjPstudzGiQ6V5OyJoGFIVpfrNqsqtkvbm7oXi429q6sHqL3LZxUvK
EUayuA+JLxyWp6T3SNrlRVQ3zpQ4GJgfpW+v/kOPfFi5g5jzswqkqzLXpysve5Qcrbj7JHQycPxH
VZSrl0QTQJBrTuQTM1cLUC/n5xMy1xopbBWWPe8cs235MCovbv9yluJojRaLolTGRhWziGTvvYRi
DEAC94iv2XOaw8o71mZatC/SWPPN9IpW3B6skk0Hiw+byOv1iMV7dGd2ow2t3VhQhLkmMxRez7EI
AP4C0y1+m/uO1hHVu9by35s9TIruGjAJGfhSKxs/p0aQ13SrAhRW9ezvGJspSdl0UGhUX7XLa33K
p4E/kA2BAZK1z0CAfWaJRhJ7IxX2OnBpCKrI9WPg3UKdc1MoHRyGPsQqoI9TQxOahm9A2WFemIE5
LKU2CPrHCcgqbwKVW0ZZwfpxeyJU1uHEzu435YrfFZpir3PYuhBjZ7/nUhX/+vVLk/OJ4D/RRh6Y
a3mY31LlkjrvNCBuuC0K6E7Q8PqU1ZEH46I+RDDiuSDPstxLR1dGiJtV+tPGouh1Kg7dO6Jz/6eD
fNWDRWTKquBLe6WIezRY/RiWaR2ylu9swiJ08wBFAOSZPN5/c4tvcYWDEz7mpJ/WA8z8I8Y9aaH1
1g9K5/FZ2EKFn0iFf9ad3QgSFeZsYlgAatvFglfM5HS+RrFI3Lk+J3wQt9UAap/hkBBhiyXX4PxW
J8ZyiGz8NwaEOb7KVpywHQnv8ROryUWwAd5WQ9uJXkpwMiCJHh5eEuNmxpKQ9MM7gf6jhBSxRND/
CZPBM3qWpGql8Mdw4cVB6gCLuQBn9LnMd093oSERH+1Zf1JqdIQFvedmUIdPBbqncCDZkNRiq7Fb
2vZBhE5+ntuWF40hTsu+OtCozTYhvbsXL5tHG0A7m4/v+SUyPCPtjLRCXHmcl1o8p28YZvAPg/ch
AKmbfWnC9ey4KZLnWE9LxgI9Cqk9iMO7vfe6DdnH4JxIgWAjOVKGxGOPvxGwF+ENwL/lkpO7aQrn
f1x2zoq/PLBOpFlIAFLVKNV1y7eR3eecVpTQCFalWfzvHXYKVA9Dnf0bisBwZ+cDZHaQoAfgnZ10
XLLeGkzi1iDsLV/JwiFlSeiIMY7XSvJ7icwPH5eu6WrHTsqhoGo2Uvpuad+m25MIe8a/OuYqbosv
IwiNw+QShoPMMWcnUsY9ZDUcVDwS5SnyxLYT0kM8GKqo13rNTkT+YwAlzgfBSRKBd61vBbiuNQ/4
pwvRipAagP0ajc/GF+LrJ36fDLZhJ2wUMdYvWL6BPyW2kpEIeyspW0tXELSC5SkUImVw1yr3li5N
o6vwqxEpiO8nbddbPfB++FSiJMNhqMA2YDP6Amz3Sectzdpp/tAO/fCYvJ82qOpMayxKCgBHnnxL
Rk6ep3ggXDwug53BeeT2v2Oy/uZTf9Vauoogq9GzOmBGoW12NBZ8KlMgDN3n9ABY7sddtebQE9AS
05rWRLWlciifnbBd2ygnURM+t4t1xmaDSq+D/vc26iTQAsfuUC9Bdo7yWzK+bWQykLfOWSM7x/gJ
72i45b2kexLTP0TRKkMKCiQ+kW3HsSupZ3xZ+XfclNYoo0M99tnoL6MtjENGhinRYrZqAYYu61Nw
72ZYUUcxnXmmXpphXc9qs3pU26uZ9XJM0NW/GQHstuXDtJIxpSjsm+pYNMY0wLJzT7VzqetA3PV/
AEnpvyZro3zo3m32bEuTzQpmDeQ/Zo0x14EFKjEnGK69Ek39iK/hLScxw85BUYF5oXOMt2zRVodq
8oFRJdWVKMl5uVvhaB3nU2X75xu5XUVlyU84X+V1OraOzaewHk8o5LKjQkyO3qHYB+w82k4U1FKC
WNkmxA8323BpS7BqdUxJsuW7QvwVtPp7sFMdVZGVv9y+paWQfJ5pLPMQjnPuBAsEC2bT9Q/2zXUP
wvFvXXiaAQ7AjDbT713+Qghn35tGbiBvdgqXxl+a2Dq2559NN3JFuwLCIna/D7U8xssiJg0YgFOX
jpei/lv5m1zNHd33lr2leTSf74cGh0g+IQ3FsZcB1bjXHrfq48cIGGlpdWDlo1CPWmbvcHrlIDTj
cu0acUBI42HcpWErO1oqbcXu0TLGPn5vY2g/0TT6s/f9X+mwTMZLuIAHF6iSRuj8zBcGtDxu2G5F
j88Bg1o/+nowskkfI5AWmYLDY808W0I0SdhYhne1nx5Z1fsUaCGSOrfyjtcm32pd/yj0XLgIaSfC
/pQrAuw/AGH+71ADxO/WQJZpdfyCSZ2N71GGrHNMKvHgEFyS59C1U9QgnSD8owekWgNcQuMtrMIW
+gZXa6HxvAlM9QDPN7QjUSEexNgrU8WN49Ca2Xa8zBoeb022P5wNWpB5k+h7usfSC6+Lix4NT8pd
RryeeM2Anam6cQqGvDV8xuVH/R19BVFZRAWdmTW2LIjagGkCtL9+rXeccdLr6F3MbP40SiTQgUKm
xEObUsP8y4o017rdRgOXruK8hTBw3TdxcGYHkrTELMHX1yt9r6UL27+/LYJ1fzXF1Kf86XIzuLBb
O/XCAcFeBQ1akYO3NavqOs7d7eCe/wHojKFg507X4ZdyTiGN+acGnqjlyimK+0Q9+Nf+dwQkcBgB
wSjxmXh70TNuYe2ChkaCPCZii+0OFGyLgHl67h8hmHMZ/F+S5LwWr1DZv2+mGEMKTGqMJQRCbwg6
0Mx48QekCxsAlO9apatQ3fcf1/LidvKbBh9+vh5h8tITnIAtaKocflfOkcUfW/u61kd9fV74ZEPS
kY6HcNkZGmSOms/IAOlzf9nmIW+iYo8Ximwgb466R35k9NcARDWMCGvAYa90WxyMs6C931lB7U1a
WvWTbTDRCcg6VMhHBVGKY0At2VI8z4c/DbWfGVDKkxuF5E0NVxSlF+cBkA1oQIpItyjz+18yyETK
jX9o0U0BJEyxtfZFMa4gW98vaODElWU1pG1gsFH/aaLn/P9Mcy5T/Y4q5OIxSbuMGV0LiQvXXSAZ
oBc7eAgysTcWKFZPdThxxqx7eH88XLy7oUjAWmEK9JuDRer0FA4pd90dA9i9ogx53oosiOxQ34Rj
ou/uH7kkZ8xtaQYSsRY69sF6uxOowjogcFqHnWuxmqu2lXMHuEnZiyR9L3UDYGg8LNZHhUMvvaRY
QSWIC4jlQFW2VXsA1KsUFEeLnywyGrguRcoxi+x00yeOjwcSNPD9WShUMzUolYa33wkLGDodMKUr
PRu22RUUehlJ9CTdT7pAG8BmynCnpHT9lBcyO13VuldbTrByylCclPAGfCh7rhkfDGsp8ahF/kXP
HDHaSfNntAZg/75vge7OJPlxeIJLX9t9ofGLvyTo7AWBGRIBZXV6M5Hq/SWUfcJaaGQcVtLbQRPE
R2p/cU6aKk1d1Uq3iF2nZX1GeponamQIq1Pzd9epYvtcMNQt/ubLU30Bonfa41OwjNXGgQLVdv8D
i1ypJR2/M9rOzvryz+a4KFqOZxQcDRyag6tBT3tT2yv0oqkEFAd1tE0mp8drHFYwZc+Lk8GMt6Fg
/79xtlV+D/RL9Q8Ck+nWu1KZ0BWhTuFVCR3uPRJrE8jS5g+zcwB/GnE+LggBCfr5oK/kKKcFjW4q
1rZyru8iuuOa8JBkjKNqFl2hrS8cMCqqXoy+yVqvdn6tb8jr5YunuKIFVcK027wcumBvptu4Yl77
ygxL9KnOGNTgjUfoYN5Nv4ekY/DZlGNMUwyoXL4ksIr9qXsFwCR1Xn5IoG1xVOCqo/qaT6MOtfv+
HDkStRlrWj0opoBFb+g4EdBLYkK0uoDjDlHhZAVfJqriZ+LBS8dwa4ncqd1OJGZw8XYCdAaAg/JH
efH44NeVVXakVGpfUHwLf4NTghvLez86V0jEo8ZyFXvZwiVVx2vfLlGlKBYIKtRgWupqn/eo3d8A
xmyQKSBObeKv1QDuPCoCjedE3ix8U9jFy6Rj66+YW0ClWiJDQa2kNJ3u557lHKmoOLUz4vh8uKGi
tjNwRZKs7eaz1Fnn9S5gxC3fPzM+UjVjXUAX2QuKKGLBT4NR9ZRmkBhWpPhdAYufGDin4pqbedtN
AsKsvRX8af05ySWVibYTaxq8tz9ZmVhvCiIgs1GbA5RebLS0Nk9Chm772rLBbaG0jT7YdHGrGTdI
kro6LKlvLK5ZFU2cArx+H0DXdmNWgy8fmCcDD8sEjOrYQYyfL5rqwbxT+GKJGahZbFEb5g5QR6tG
QEtAxxuOyzX0rftr7kYFQPZ6eKej/67KxSZd+A4BnwyISLEOs4hIykjk7PjvAmAipPcDxsRo9s72
2TWBjH7IKDDDugjeVG2gMYef7cz3IFcAs6+Vjk74cRQcO+aFHvLQ5FefUgs1ypMXLnfYeDkN5EaH
ThntwqnnrKRnsp70NHdjVEgI99EkH07j2rEQngMDhQrmZNsXycfsC3v9nOQKtV/ODW2uJG1Q8p56
258O6xm0wxQ5BEdSXSGHA7bhVjHGkXMV8L+9Brz488YxqeqNb8IZZHeLgbR0M6GEJm0/w9mykqXH
q/MjyAQFa1I0KhOSVpiW64c6TghTZrJlKXV8wFHzg4cS7TFgjvCYzmfgIblgueMliWN1v3hU1ia0
kVdxurZLf1szJvyWU/2uib5wr5swqKvReo7ktQDYEA3VlRZJSkewZHtiKHUSm14QwGTvbydBGGJM
Vic0UwBrx4i0XfYjj/i8QVQn18u55MOfdgZpOUe1JcUYXfXfAd+HadrnGQTRifUjOtDi7aEy3ljx
Zd7s2zw4sAh3uBhBeSSmyEwUyu5OVgEUItmotYNWX+uFogFUvnoPxEr35/O/5YMCemBokEJ/HFqd
Oor+dmZuaathh8WwucMpfrn9mL2AAugDjpSXNsqHEInY0OzpaqXzeSivRoW5LNF9v0Fq21yqgFWe
rxRNq8KYsjlpfzzlxTLVPQEhS7i1Tm+ESsb8LxhWTD+m+ZjZ6Z2yUd5ABtImj4cZ7t4rsr5rV6fr
mHh/QTr7Kpt99VOhSJrrCjr8PQcI6s6ZX6nnW/0t7wpZjMdyOpFIlx4B+VSA17R/mlDNg7/deRqz
iTSDeQYj+7SGCc4xAnL0ETF502HDn3+aEKqKriJtoj+CrDj2Ie7emwHq25s3L4MOo8ultU+cKi7L
17JXMwl+/boVW2cyvpbLD3MWtAjYDC+I28JeXzDuDjoqyV0GZ3PAzccIJHn4EVp4HEfLaZEX3d4H
HgbVOG0b/feBPhPekWAG8jKJstsyL9cQH36VEDtMS7QoDoRgXmGybHQYi8SbeKfiFX/8jovzbJTd
bFudzqdK5cc0oF+xKgyP+M+n5vd0z3A9p+kWdPBolJiw+K6PZPSpWIiDNH24cTcpGeLSDVfYKv01
hbfGS+9IEfPeMMmCE9VGknO5RkKq1N5KdYzhkM1n7MDQfvmAB8OBGG+gOn5hR76LOYY/1OVYZgmg
EtwU9uZ0SK3Wg4e5Tv5A97GwqLiAuu/lHw2jJ0FJBUHjjjFo3EEzFxDHlUBb+rE7tahS9P5xK5HY
KmWPpBUC4w0es+OJt4SAyADeJnvywdp894faNQ/HnDY+YuD6vbTjlmUVQ9CF0W4k6iQIad9aGitx
VetWs4G0am5kmMIAXnNQqiZ8SVgHFrvgUwJeiOE6DThwM5nYXBsqn2VKNe8+IX5SSaIUPdU8l68I
PhCXwvVp70XV6X1nfcQSwJg6rT9Eo74IHqlF0mtJzENNXGCLZ/VM5xx/ViBXHWIyHVorkriLuEsw
4R3s/6z50tWIsnEBSClNG+G+HqbggG6C8ghiTpRH23fr5u4O+wWwnZJq39+076fQOGBAYgiEF3Ty
97DogXnzVDpHmf/57Tdqyaf+r9o+Ain8pEi6qH6ieGuPWToKLA63TL+dbtLENiyVBc1vs0RGkuJ2
TinHa+WXkyE/TCr0nzl91ftPi0QRwyRXg74d8Yq9JNbcMNaiJYR3gKMKq8DHmgPBUYY9B+KQac3c
G6mZqglPhICAMibXaPGBziyDgjR5Djrt9G3Je9k4Z/3lw2/NHWD2WgKVx0rSkX0SJVcfnqgbQ2Dq
WZ+UedMqo41hnDyPGK/CDo+aEsl0j/+3gbdRN0fXt6o6/EgZ/LqmwfncUAOqAiXjlqriVlMcYJeg
bnl1YFvNQRmiPETvxV4F7dSXVxAK6vssuQZEKbUBF3RC5acBCiu0hI/PLM1uOuU6QXcz06VOn+Nu
7ax4UqrojrZ2jTrqym4nxbzIsy+P2wF963Gq2C1zztFSWYiu2iZfDdqXu4Ho76S0hGqeq+ehXZ51
M2+dESTGG0OlD8fRM62uRX7at01HieZcCwJZuXJ91j2OjopmV2lNWNTVsnMfjlr67ue1z56nLQDI
sF9qsA6rC/gVKs6wcYJHb/kNIEg6zUdRPYgICWjTb7PELgpIyP2LLoawzSrCWUNGzS5P9V1hR47z
GxKM2rORi+90o1Nw0TwYFNruN6bB80in5p8Q4+lM9mSHwvCDR6HxWigC01ste+ZMZ0bwI/xMILLn
HfdALb+5SxQIXcrUL5hqW3gvP+8hUvWWlYnnAY1B3b+Xk7MRQlbp9ZV72oqmgTLNwMSfEmVvhavN
KBoK09iRtb8x23uSW4EU1mLU5UszeZvoj0/pJjHERDnqDTXAUJk6ESNtLAcQ9NjScYR8ZuCun+Jn
pWn1wqoxywGog3+gzzkHfpm8T7NWjK8MQ18a2vRLj9agu/07ABJN4ZSeAinRS8gVIczuGvrDSWc8
sEAhBSuaMke7qFgL+Vi9zwetkE5kck6XCRGflaVQJwvy6/N9f1ogi1d/dIcPWLDf8Y9z/jht9twp
0V5XotIVRZlGUYUznAnRkEtDLPzZ9dW0DKBxoFbeKZUK1mOZT8ZJ+eXqeZoy9ucgLFq0qZzebKwL
vB78Xg29L6jv4+cJx3Vxas1JM76EhPZBvhL9DOR+b9ROfB0lpVejNzhMJOAtC8kesWB/SknEm2Oa
iT3r/zMpPfcn4tmpf6jIEOzn3+w/z72ZY6ePDwpyAKcmUFPKJ2jL1wJvSaZo5rBVY/NXB6RDDa+v
FPjeyJn/GPvc76e7yCr56m/H6ndDc6dmAynfLNGRCcKXxirth+PwP7GJ2Gq9hcXY9RhuTsleb4Bg
e88PE2PL5EvG5k1pSeEO0AJP6/k70a02s/tRIOdgTjCNo5IOh2vVtbk84Dm7P2E46QBkk5l7Yv/q
mfExFizpb5qrTixdwCujVXMJfZlvweNPt7iZOUCPvZaE6D3nJVLnflMj6jHvFwGXOnutAwNsX17t
tB6j5QtsNNTtqxNENIwpRlqmKHYCp9TcmVEJylejtX1v390L389J0wF8cfeo5ncFIHinqEbZCml7
lvpXv9HiYF06s2aHLyQ6u4B4uqBaEufspqvG0v85a747h4JbAo5+T0T9Vrg9rfpOPv0yPA1WdwpG
VGRJzdnuoGGt5V882Y5OXm5FcgL4S98vJUmvka+2b9/gA60uHg3swbkAq/0VCtQVysgf4MvqaY+e
GOa5gYSP4lOxiqqSEemc5O1gEKs5ViTMxuClRkYR7CKok2vjW37O9xuiggpAZj18AJumD/IYS0kU
RHGisDVBZkdCeJGq1yNC/niAYQyHS2zbq3SQOLlqVkVzgsaaXTV86QNyDmSkfHTCsdE2g1xGgXSR
fSE5e4tasEPY51/sVOUit4XX6r+YmEuZjDnw9FqR4kxDcYeersV+rna0fPCtNCJEhGR+ZWlRpe9c
SYn+Unq/5W3UqDcwjRj32ZHTpkuoMI6873MkXbgEjXFAytfTJcf21Z7WXytKaCPAP4NRwGy8ce65
XKQ+Z8oFF4lh9oPPEzFClrOgRoibYdDS8GC5xkD9TzUbQ26rglXfsebacYcojDBxIV32unP+CHhE
fR9gcpkMKepPHQXA/Y7li6l3u2SObaShMi0d3PO5M2f/6oQtJbncvLzyKfkM9lArxGDZ9FCjzJBL
c65CF6gyBsIfGYaxxTOjqs0Qv18j633kRMn0hMzStoEpkUYw1w7YhrIht9pgJwiAtzWhT6Dbe1v6
UiB69eUmrmp1Fz9ctUbs9c9PhqV2MmN8pULulguCecNtg657bQWlG/ZhKRApa1DqCDQqlFN/AIjM
P9nru8Gm/8V4KhNKsIDywc3ube1Ape9XKP/PDpN+K3sX0ZFawsYkVhNP5/eR7S6dgQc6NSFxE6sB
ZDUF7QsHMf2d+viqM6xEEdNAfy0JezwOsYY/6CuwVUsTysRTG/4Ai5n6wihWhEuATT6SAS0FX8W3
resitR7/JkuqREeU8Tbz4EBt7ThbG2GLN64iiOcj1GW/INwFJbac4kynZuUcywRZc346rl7YO859
M5XeqYK7qQNuVxSYyFNqD5LsfThLWVqy8UUqmyNGi9f8Ux4/ze1nSHDlVXFRON/PttzufJgXwY4l
c66hz56y2lSUksatngJB7ooGdPC82e+cb/n3ozVHiwKHfBcVsaZ3MJkd078NpNNppvfLET1eo8hQ
usL92wlfZgyNZkvHNJCCfscYRuZPdx1TwQa7qOW5aDsCZkCrs5+SJAfxf3bRnoqO0biHj++4r0ke
/qnkklzfo+NnEuFu3L8o2QDy/3GR8oyep1RPBRJ1F3LsE7CSW+qmCC4HHWZ9eYLD90x038Yc8DCj
0lCor17seAhmgLikwwwspDPbIERaRCYiGLQJFqjwGzX86Ojb4SY7LWdXc20LfjpXc8Cbi3xDZH9Y
iFhYnB3jQPZ7WZ/KO8YnjYQUJNHgV/DeL2Azz7BzejsO+tdZHiQbGyqsuTYbAacBAUrZJlP3pwg4
KRkDI/g47gkpchwqRnZf4A9pYlCFbYcNbRKE400cTX4QZ+lABzb+IcmLMbZCe/GzEELSkwYCpfAC
ELUc9WeLbEIPrcBRYZ1Qt1O8ujs69I8YrcvmBr/4jD98d86a7cOpIhQioQGxeLjH+H1fbPuzBE0w
YW6cMqNgQCfSwSuu1wpHv+gB6iDv3Hvxv+rLByo3VHGN52vJWuAJxmvNu1dEAoBql+YzK6Fn+dCo
3cVmt9DQXIZUdjlRFdpdGA4CPFMzo7+KxlumTuXtrL7odeql29IT5/JBf06dZ6mRajceCVBab8p5
p7wiL8V9mcOC5xxEI3+F+BO3nwdRqigyLy2ZKZNc9fwcCvimzX4LSNagoODT3DxkaO5khe7/QH+x
pWAKADZtpx2ooVi6YOvo1TnFE5nr96T55Uo4MIYC/11uW85NRC9sW5BjgYer8FhAMpSGCiElxUPw
aGbQ8Wkf0z6/5Z9dUh5/3gStSxW4Tzq+dBbc1j9aPsY8Da+4Wlt+qgZGwW9dfsMTUpSDn2vGYV94
XnLfjzaRy7vokB26AiCasVMlWsnoI0CPiRfQ7boVschqOrqfaC7KEm2maHLm2ndek4EfsXuy8Trg
RWJa15ydVkTu3JhWfD3UiyFvmBEiXkcPrsBuUwRdXX2XmXrMlRUZrZjFT8VfRqKx0Fy876oPDSlJ
bN5Ic0c0RVEzdLfhgnmxnosE4hcP6xLa5Ti9sj4Jxp4sw/69doEZxjAbraXd9grkC7LlplzSjaCh
rDJEly8JNZVpLjx26saPwGX6dAAvlD1PGu7xuMIBHreF8AHnCZsqiJpj18WccjenGnCAV359OB13
LN8iZRwq0YX3RTKGtKrcrJLApcGVBTTaiZRulcjrFsfX7o6NnrReA/RjKP4CIogHipvAv0dANXWQ
1xWs7frMFEYJQ+/5QrpPmegJCin/wD+UGpYYv8N8pZBmA3kZX4lISNgqFv+1+ay40xcId2X1tzXw
B/o5kFyaq7CMQ+zwohDauNRdpy5XEfBpqMDYy+jWNXZ1A9JMoVG0WkrB//wgk4uxW+wmRaFHyJJW
WVm+35NE8Q2qvK216KA21EGeUCfTw2ir3k2517skL1Y5QR3VbQ5+CmRemgvYRsXxoNLvO/03WnXi
ATH3C16/HLzRcloGqCEmMi+FFOJmimBZ/1l6yZKkfjeS5kdjfBCIGvJfQVYIweb7eUI8+S/Z0sJq
DLLnkcPnHo5eKfBfypKHEAbGAfPGbCYA/wJobuzpmsCrireOGm2TChb6mbi7a1zT/68hH8CndzSV
LsdSKkttSkNCFN2j0B4vKDAis+GZYUyOYI8g5m4NmGXjdqdUyLkVFWxCBTjx9F7h+TeDMWV5I3Oc
D4Jd8tyvTdx7vBTPAkZTmtG5usGnNhQLmfifFBRzs6e/H3Soi6I8JonYQx6BnSw3WxCiLQLiCZT0
CY2jSoTPfvWYXNzhpUo95xfEtWNO//z0rKijvTxFUe4zSMhDsPlsVPlOxvChCw5oJKceXOd9VzG7
Ubu8yaPSb35SHXBCHmxOZG+/UtCh+r5t8n475qQ6mfYSFKmk3k7RAC/eG000BEvvWOjfdlDDNWIt
7mbUCRL4oZa+f7OmkNevfBtysiApIY9SmRmVsP1emvWMUS8967ObqHo32rvfieN3765mgx86yB7Y
5kr2GPdI01uWReyaci1LqexUaZODr/qTRRylZ02bTb0tDogwvnNiHJGQdKoVXyAqwLEsQilaCcKe
vsCYEOYpA2sNrVTomjHVlKm0jBqt19thrFR1cznWe03be5gvBpNIvFaRDoyB5jB6SGuerg0TuqQY
usWS84hnbOdVfgMIScMmOk5huuXfac7bM5U5qzEXLw2NYUdEbva+Axhuc4vX5xZbDaOCT5p4mQHi
I6gIBFvucU8hnJWuIguxFjxtSuStz3/WkGycbAgEWo6GddqIdjlLepSU6OOBdCtpIN8tWmEEUU35
tNdLdHdTwk2DVCfCAdquepLAOdBEopWd5mT3zGhOXNL9+/ATU2Pn2wxQZggvijImuvAH6JDVX08O
XeTvypPsPrxozTeEycE17sHNn9jBxaTbjzgpRcD7nJ9ESY73y3OcExlZm0pCLDU4GYABJiH0tRZA
87CYp4Y2DA/eEx3YH71K7fvnUcLAYgOpK+73Mq9Nvg83VIvua6vrGsUKqXcUe3Gyg9Qa0A6zWlyw
I2EKPMCG+8dlqz4cW6YYy9HXrs1GusUiNnpJy9X0/mejqfQ7H+HwL3dGlcaORaqLIFld4i1SgDMT
BBkB4zRwN1JXCEiVzrggzxe8jdI93SWjHFyAhRkicB0eC3YsqcLYtdoIEa1zUuhC8BZ/fIGURPnU
DKDPC7fbntf72RMcjhonbbBoUkBNuGfdVIyZeUEu66vqP0Ef5FDMouC44nio5htyfnRiWxtYcQjU
4L6MbsgzYRpUQ1FhjnNH/5Mov4QvhY6eCCyYg4YydduTF0NLXtf6TGtdiC58oXRLMBdnI+Ufvs1u
mFafge5v4mlCXYiI42B8nk4EX3Ft9ytGKiElOQ+7kZFDfwH4ONBl0P7PulY3sKyreC4XO9J8vN81
LGqstwChT5AoxguPYWZi+8DAQjK9z+yYU7lTy+DA+xmreSEXhUgQvqR2Ud/RmpOq4O/sfJrrYDs6
8V8hUvMRpLd3AnQ6RXonbvyWY3yL71pN5IdY0YrXXWXAt3GdHy9waOHA0NL0wezsNvQQYKW89cl6
J8Hh7RllQvLXOC3jMJSe/Xx5GdTcFBAEATHuobWxTVEv1Ht7pxcckgz6wB2CTSc18RSRZs5Jnzw1
NRz/7YzHdeUM2fmqbQqKZ0X1O1aHVJjeZksI2tZi6kp9s0ZnHesOt8k0ZMQiLPBi7RuIdqGNrxVZ
e2F6gREyRb8g3WCDcRpGabSxcNiSPyJnmw33I9FSZj5zaBP36ZUSh5Nunr+Nzxi2Z6TAhb14R4gI
jIcM+pkuEcsaS/EwY8PTZw3/kIeq/0MuI4ED4MoWsiDwcEX8S5GDXEwEjmVd2edDEYoeia7Wa28H
2fqrVIZ6qKK+9nPYssVrviikXTP6D0OGFSsQDJihaya6RGcjiHedLICvgDzBzeFv80umPyaMwylz
jqEe66n2Yg9zOOTJDNLdusxEUJ0G4mN/FRuM9QWDvUmuyf6P84dOUQZbEVbYji1m9W3vOrR4h2v7
uoc8vj67XhDYS5fDoJSNllarWbPW9tae/P2qW5SBA5dL2XQU/O3l0Iruwbc0WhSF3cmachALAuVZ
Tw6MIhjzLeD8v9D/NZn0muBFeLMmeDJM/j2t9jU76WZcTwzcOL6bTRFMO+sjt6B2hJtagjGk9iIS
t8vl2haNsCgO9skAR1TNbvbosMaRaJ9y5dbUgvzl+3pia5PTr2vWFj72FDnIRv3hSksQRF735txh
bMlFplLSl0mVOVbk19Hfn8chGJpkJSAeQ7M0Fz73+hPa0bJoEDohuQqUZLgP6PCgCBgi/WbCOYgN
gWaJF7cGOr6cw8PmGxG1O+4CY9FIMRSJ/LtphT/LbJiwtdQCq1xVJilq2zsfmhvTwcQ2P4itaADq
9A5THnUkKbYlIQ6qU2h0DubYlHbw/9vXcOBpNKp70nY51XRdFkdpUYkpafq49WCwhy9+bLB5sRvw
t76bnCSp8wwwStUg25LlRrSRZSswiOUKPUylt6MyKiqHccDOCgJvO8i0kOmfcucdglhg4yFVSWyF
0HAvRty1/G0vFvn1+tf9NW46c1bDFzyKF03mDSBpGB6P7Ut2yuCdR3ZwBr58sf+ujgMQB0fTtsGR
/5w8mr1KF2msDaHIe3/4uHtXiXN2Jd8tzU/k2WAAfkVjPvRDpaADPyZwfA6CtUyMBrDuJRM/eWx8
tNGN3/huS7zaApAc88htJ1yd72s1xOt93styR6sLKixVnQm7aiS12pUGTywt1APFUVz4u65qyLH3
8Eh+pUpllFwFoqr+EJpTXt7mGKTrdpz0qXCBWuVQWb2VAD4FRWzEzJxhRv7qit1K07qk98wuChL8
ElDCqyF3YVL2I2BwpXC/PH+dy/xkJUu5Ld8Xx/46gAQ5B9shQHzoprSNGyrgEltIb9qZbP1jAd22
jzq9LkkOIEbsfVMyqVassVHdJ+p7AkAZLl6ttlRSJFbrJogWlLNiZ+jDrJBD5dWi74iCyZgZ/t8U
/GBmYReQvABW0JKHFlbr6zkzTwzJk16mCbQDpa1H9P3n9TKGxbhIwsF1UMIMJ3BhwUdcraCEMdbp
eSD0IA4thpTm3hqqRmK+YsxEoGyxMFmqsG49tjsWN/id+WWxvNht8/INBSIEC3bPhZ7BL/q/UK6k
gcFt0OVfYGkpIL0rh21pT5Pv3xBrAVFCP3DT5UvUQgh88m1Q8G6FlOK7cnUFDMURLWePct17qVrH
+J1DzasknCkJEjR3t7iTjTyfQQNaGfTJ4cWyg+0s1CermRX7YC6bpiKR09HO07dubf9I2aTU15Nx
D63YfE/CHi+eR/Vu0HFpyZ2p0SvnqPGzYudm65wtz//FMzy0LwIdZu8Lfzb6VoJug/9MfiHtV6zM
APYkLcu2B3WEnjUghrhBJn/kdWjx88yguhXM4quyDyaYJzSxspIYEfBBFbaFb825fN9DotjxSOzz
ReqSvN0QtnidrkeRQRGFitAUVW6qeXKTov6uiJ86Eg1QRiw11uXwZqNq5Hvm3O7NnxgYC1MtlWZf
0G9gVL0rMDaUJt/MPICuB9MGSwDZSM8xkNJyInWTxvfpfXBIju6lamV7J7DaXG6a+RItVlME2sLS
Lk+hAKLbWLP5GZr2yNCEU8stS8bHmVL+ZksfNZhzEiQfXa/baPewPOFetQbKYU6PBHHXF/O2zrnG
YgjMKgOb8PDbBl0u/Pmi3fJAEgI+7z/zlJG/RZ8wJyZvMVeuaf6CTtWneQCuEelWU9QrSL0XMaQY
nlVoLQH9hQLo5tsOe1StfuGBZKnMpp8NsF89nxX5zF55JwbsiQJKgWDgQ7ZUaGHscFYfPqVJjsl4
94xB9/jK2RP4glHDfHYYLQV4XW2ifIHxEH7yVVBgydY9mV4bG0LX0uCqqYqZRr+5jpQ/Qb899M3P
6lYYc1853xWqL1AyFwIqBYcWRHUZswJsrCh7huaI+MYT8DVqqcUf4tb6JZuiTmXGHYVIATa53VNi
NDsiYF6ELGhdqk2IFXHH8O2RXGNkoZFJqsFrpIWwHU81iiQHwXCy/lheKPLxZfycQO4RUcOsn5qe
/QNAbvW2fW+d180fgvlHrCd0kUyjg3OgmtsrRSAKiaDbK0ZiKG6A4Ecov0vrbLdNwpw9ztNJnXhf
b/b39buZt62x2avr5JF1n8/3m4VtHTphtWvvcVYi4Ip6tSlz9GRwQDJRfMbWehrL19EqeVaWz0Mj
DlsSArDcds+jI3IskP9sFktolTE7X2tU8sDnrblv1Y2hNXEJHYT7kN4bUIOcozIfolAPtnUFsbDu
J2SLhFnchBf8yKfENaijxrV/NykuQ1JE6k5clI6MP8SGE6bSLk0X8aRz5xUgT/qdMJBVMTSjz0nK
6WYChiej/lstWFPF9nmdf6xgGheHqrVi2CHLcP/uhAYhm1WcPgkTbrfYwN0dgzL6UkfgSqKrn4D1
zyLGvigl8NLxp+n0hpe6CGkv0AgxRkiOTd9lhvxcWUSivLF7d3JDP51vCgh3kow2nOG3ga+GB2bb
QCbl2LKGLb3lMiNogX88EBzbL6LEFSAXm/tKA0ck7BI192se11PBWF7z6ZspVPgtbe4YMbGJn+i8
cyFj9cqLMegnvXCtwQB1EBLURU5J7ftwW+mxLDfI2XWBNx8tD31kaa2BQWN/IgoJQRFAi6mIDVcw
H4Ufsn7TZlCROjfGmsknFDDJZlyAAmnr7kH91Y0rwyMNMuXATqw2MNVjLENITOa1Rv5sSnf/X2Hr
+xncJ3fIQtiYbYvCahPD0Q8fklvZR9UQaAs5aJvRMIVAkj3zNEWjJjJx8zWiBSo0U2etekVzxV08
0PM6V8/I6KhIlou1otfUKU5CTu6/f95wOtSG4HBaJgG7lmICPIsFEKl53y/51g6m4XkJA29CFRRB
hvGtZ+HxLmAxVS2OdR8bqtQgGxRGWPq1GmFGS5SIOFfdFz8zzZnLuhBz1IFMcVqxVWqGYs/tuh1V
319bJ8l4BZ1LF7BoM33O4+TmuoJBh1Mu8jcC0d53U0XjyuW9EPok9USfF9JFlhwfUxYy2nXJ3H1I
rgElEpMDSKvv8vMzVJONc9uXSEYnshKYLUB34IHqmtQ/7O327eTvOYjhapOZlt9A6Iz+8A6ZkQkA
nkomPYobCNAA0V497GjYCQPiY7K+H3MBc2kHsHVFFzlJ1jUIyk+Rl0DGUhCXYZ0XBeydP+DZysP2
tr/gv+m/7gzMC5lbotFSfe6igVSjTGoIk9eqcFaKs5bTNY4ciYqEII+H68giP1Gyx60DJOvW3GHB
pRiDLzXSDJRhPHwn+xv68Eo9QZwaSW0yKBgzMzOucptYIApXs8smTSsKTdLMlHBvOFK/USm7eK4D
KCLCKOt8U5cwC9stSVaUq7E7F4D6JRe+hviE/aqBmoK/FczEYHiuAF6tFAIkzJc4SFhTRI6M/nPQ
kNppJtrsJy2sZwWNZeUkT4eEk3Q4K+XrjIE6f5+Rp5+Epb4pDV0bI6i+sQYA56DSMgniB+b4/+Ux
c90JBwyBKJJ1xgxt8Zc83BH8gHUdrbeFcNj183WzODeoym01MKSoM3uk4plDu9yzLS1AmofFvY/N
5r/fQnMaNCferZGS8wRUIU3hZ4xM6lzlMHUz6a2bYVTrWlgybZ11NUHcd1bAAQcm7qVBxGpl2o5y
QJDHyN5CE3ofK2cj87Bhcx/Fm5np5M+pcGpGFSp+eZ8urOYeOoiKoOCe+tV8u0dtZZTdr49KldKR
3q97RCdhil1vxyhJoLKWei/1jF3hFxADbfWUaFmokiUzI5lyIWjodI6rBtxhtut4KxhhchOdIW/D
rNyyBwROuG4Fa+e7mms5JvcQvDiSqWeFDdVFyxCTPusxrkLcxBweF8ud79l+MRBjwRKJqo+7wFyj
0HkxycIUTHHBcMd0MlnryzPBlx8N+7NKIre3ZV5Lgw2mGpAqhl7nIcA3f/lHiqWqmKw+j6AaH2mv
1WVCCaD9LD9bDUQX9jLLZJVjjSv0gX1O4MkjQ+szX9PW/Es8rvbS8YGznhn62gPupV8xL/FL3WVB
/iAhFJ2UXhjXntNXmxF5blVjXi6fGuUnlog87wWrRs5DYpQbRXwKATMpvPrqB99IQEqmo9X6JW9U
g0dsaDZ5DKAxslw1dAv1Z6F6XZXrm+AqoERiMVn9AQ6p/W1CkUgLeyCdluOUZzWFQ55h2RiQbinM
pYIWAQX5IpbAIe0Y20ZulhxIxeEVws9gNSWt7pLEr5vBO7tMCiLb0YgyBtA5o9N5H7WTDZDD+qXm
dNt69tF/5HnyM6PkF+Ir0yuE97sBpIa3Uay8oUFFw9CRapvSIPHvsUuoKt9cQl/qVxk3ZQ9kz3vd
A8plZMCjVgu/MK7yVIDFHWOVOwn/50BeHleDXyCVj26BMY3TW1e6sss7Sc929i+30/AIb+2SEjxS
N/rnTK94f7Bfignz2XJRx47nIQR2QUChT+O4UbQRLg8vPmvvz4Ejte5awB42XF/+OOtt4fwqIP1z
0zsxLLDviUOHSCbx+1EAdue1c5/FDCDkR2tkQf6m53fqUm1ycOL/0+PnBHQJxqrUY4H5u6uavTQz
BK3vSGpcWwYJQ7FjaicGoFoBfq5uW2SMcxB1L09l7XVwdh2dLcmBWrAWABOaDZUwSvNZQjyGzjei
TTvT3r2bpceE+pkLc5MuPbGunX7al4BaCfmVARpg+KkJNa2YYP+3dfZeBhHCk1mKLO/IeSiL8Az0
X3S3f0jiAwX/Jax6vsVrx1iXpP6wAPHJjp8JZ5zjZCu/NVsj+UEX+t20EKnm3kP5fIHYWMCJhuZd
KVFhl39QetLVflnqDJmYuw/r1/KWN6uN7grYB7C4ZKsH7eD2/Iu+dvizd7J2dryhTLNrsmNoXCDH
L5x6ouHlFUuyrm4ngTS9WPMMebGo6oJezG5J79st8S7DHTqTDO+Q2mxMnJdIOyKD1jbg5JxpRBNA
fqRNtpuqHPRXsrgx+6hHxa14ToDApbkNwew0ZupX/jnyKzFcYQ9dz5A0S58qxzJ1NHfR1v74oeWL
HjjM/QZ/+TPb8O4EDDAi9+K0cQGv7e6RQeI6Yj6gJU6wOaDGg8+t9sFmeqj43hn5Udl+lc7p6Drb
1cdxwenVa8oIqDPCORZRGDqiwlgEkSMRZVcjbudx/tCR9XhRzD1+uuJKHWHgPnSz3HPMkvEoFpzK
mRmgc96CW/dWVwIK/GWUJVAp2PaGpmSkestDU/hCASpz6UV9a1xJ53BANhWmcUknEXTvCeNqXi/W
MtZF3iZk2FU7zJ8mUFUtxNqqtKl6eZONxXWrIJcWERajqeo3dci2ZZsYTWSlhJfXvy7hFL4BA85n
Pb6r/DIiPUiODuQ2yQqGiReRgiX6dsdTCPVDLzruePEF3Gg3sIzpiYuj3BkQO2pg2N5R2JCOixzm
HxhFNgs1MwSuyhME56CDwe04HVlvky28PPdkNFyvDZMFyIqDZz9tFv1bkVaIAvlWh6JlyEE65LRa
KQXtCOkTHGtHMge71u2RgeD3Vi9Nfc/RR8ebtAUiPjTezAWthxoE866wHYK1yYlYQ2EnVtazUaSW
mueLbXBVV0WnpeHRLluw3wx1vZNCe0itJCrBHt0OHRtm0ncRV8mxxyXqZdftVNEGOxOHCTxhZApd
ENdFn2orC3Oroityt1yMzom8p4XSXWZxE7qsJi5KpUFqtNueqKInDsPTaCJngR69A3BadNygBJb2
b2DOqyZtLDVf79i6ZBR2EItPLBqfV5waxqNn/VZymj8AIDsfVLMNZ9dDPHbgr+1/yQOLgiSeH4CS
MxzaDk7zdMmwa4Vucnu0S99UTxvnj5eS/kfRsC48HfQN/ghIfxEKsyXVfKnBoSbbPBQqlAHhNBJv
JHi+gX37q/1E1Gszj3BiSPawXrqZ2Y9P6hOe9c/w8Nz1Uhg3aprzvNDk2t0B114oOhZZEpm2c2CD
DQ8qPTQvpi5Hry07tpqD0yT6kKDNK4SUHSCm7G/COMgMs4qsFKOjfPN/rolQB9P7rGtEEz9i9bb7
nRsjYWcwovFqa6eqoJ0EIgxhloLVMoBTRq+awWF/ZiDjueA9WFl9qKORU9/b6uwKd/zZkq7dfiJk
V/Ao05333X3dGcljNYbGGilFvHmtNFYeheOIcGIoc6sBexvEzq67iShoVkaNZ004H1DOMy31toV2
aloN1MwCsbOEO961GIuvcqv+z80WjrKTlaKCHuurYvQKYGPjN+6atwex54mnsdUtmwFmPMCMno9v
nLThgRivwftXLZLUxzoJ+A0VgONwTDBrQhLddxXfdSy5Wgw1sU33sh5k9kSVa9H8dm2ljlnQPcFM
orG5COi6lb2NwAhsQcrx+AGiPMzj+ubLN1lQlmO2eGSzwR6SuvhLFzJQjyAhNQd+YFw87dbFEk/A
u5A1whXipxerzYik/ofQPSCfADl+FZCc5Ml371H2nuPFLMN/dQecsor7HqLSmHsdAcLFcHq2PEh0
Xf8uRpjaYzIylibzRtkyZjtcxyMIRnK8DKC27V4y+gDouVp6qwu85gPO7wmEcKo+YMyPeYCif4xl
JgaMSQuJeD1Me43bEEdkPXUCO42U0BdtN+PA+VNqVXJDGpMDGjsQxjaXSbPKWnxVLVlN/heNGORg
pcJGCil7g1fcpA6nMp90osNrBL7F7gPgY48N4tRMfkAz5kpmLvw/IKYBurdqh3Y5zq8GkEKkE5QB
xVFD79TFJRWomwu1JmAZV2BQjh2IZ4l7cO9gTSnPCwuc9owhej74gI0nDbnsyeAgPRKuMmucQok7
T156Kb7JkcKM0rCgTdAyElSmLcLiIzTpHBV2t2NR3NiRnL956dWJTekvmdvIjnq4G1RcUmiRSQQ5
XkIVdIuYAeh5F0dal3FY7IaiCueSUsAmZW9UhHzrvt6WEIJnRD78cq9f0of15l76mCmruI7tCX5+
nB+pzcvHp+o3ui0zHgHor/jvgYcbCrbjhkCgSnzWA+qqGSgMedMj4EVTM58C89hMmXVRON95DYv2
kuQW/Irw6CaqBnfENqKRIheP0n4PRDuq6xsO79jxV3Hfz3aKPqS6/3CbMYAVefdxlPO65NXVwdcw
plHcn6hca399gjbJ4cm4ZgnZJiptuz5qcVH4RjpbvNNpkPvwsSEOUW25ZLUr0WqNvQ+oOKnLNW03
6Z0ZbkA7BwiabfNoqTa7nz4k4VO1OTcQ6XET1pZ2zLXMdmSm99u3bVGSApK3R1iWfK9+gGYjD+DF
91NM+sQvDQ9Sjjhqgj4ymHe2bYxHwdVbEDz3/B5oyx8RMxWxHCZpae0x9vgxLEbpg6ccp3cgmk4k
8Gh+wgWB4Igb7C+tBmxmVZaYOw/iYxwgvLGNP7gBpx5h29kFD7gL8n2tyhLTd9DR5zt6igOzto51
FypXTUeQpeZwtr/+5YL/JXLC2v9FaSowa0YsfNfA6cJCVpV6QaXrSScd2/b94tfVl4BLQEtcxiUT
wYzr1NHnF9OlCwx43tW9PVEcRZrrtcuxeuHwliO1S91Soh+gaV13y/OgMMi7a281cUfGEm/WdpvN
hMyoOV/8RYKRjzBIaxSIgbcIV59fCwf5xGJfmE8bp1NxNWsHhNjjSkA6by4m8To0pZyxCuNMEwM1
9O6nwGTz1XOcwrnJVNVkhik6YGoVaYC+2EZh9gw/ytWxthBTws8LEhNFhlwuGomyR6G27zzfDszg
Wgu5lWozebnqI+YCWVktIZQ5m1cTO1AGYKdhLbd7wsYFt+tYfj7QNq1BTPJhzUXySmkphac4kC+N
WmFvPsxudyySHMTaV1SXNnxlq0Zc+qAezMxHs2JxDGUmGe08ELm6o8F38//R6JM60iJmpr4HjSTg
/4Mw6ql20JWmEkVTTR7EqIfo1XCiAkGO/vMPQYmwYbZ60Pmo9Gw9IMhkPrSoeQH/ELD4GuFQSGXe
0ibWMeD4dgCmnat6OKYf0UXPUJ3xSwUnAnHyFr7eo24MOAXm63Kbg30OP++Qw2vzhhc+JXoIvOPF
ZKbLNCr4XDxL5ykM4KOJoz8msfeGLvsnoFmmNnza6c2W4o9BXlJ/cd3H/kugsnU5bh+s9EQLhl/U
JXIlqsKjNIl19jb80eENQt5tQ+FVEh30t/3YD1naLyzcjAHhdtAVzECfqQmIITHoVBXwqaQ79uWb
b/3dvduS6xZ32eKex38MyzOczQYvpqDdmtu7Ih70O/Ll/iXdEm5NGW5PIIk5F21Bo2TS0VfuxjP9
kYoFTXJki8U0dS/toIo73kAphlPHhCNRhR7IxkeotXOvCrLYdXP0HRXPAlNtEhg5qsTeF+YQF8OG
PprCE9CsZRZXHLP+kcmq0EdE4F/pBZqeu7SGIo9HfRELai6GBF4OZ8HLFPLhGZ/GikosINvAuHGU
hzHiYMeR2gRhjl3DkkMMKPUETuVdD3oL+0zIQkmY0xhuWTE0nDh8NVxVPTJ/nQiSy6jUiPkaS0Oo
DCF+3CcowEiqOois6YV8yOYHrBf67BcQjzV/uPa3lLm9swQ2HUHzK6qdbH/ssU9mlPgV+PGnn9+p
yx8CIwtlTiyF0VJWg06axtCAH/aEPu0UzMttBcJHqJN5mNYL5jRmd3on9DOwLncuMpbsFfHVzTPp
UFihwRW94XtkGZXKXU4Ggf71i5k2YztsFBoUdv6XdbkzczxLo6EJrKogkA7KwjWnfaYzJRR3DOv3
fviTAAjDiJLY+r6smkzog7vrm/pB2UXH2B0P8MUnCtHhbKqGK5MNHwvF42I5runrba5cYypssNjh
/NXZCi+SwF+TzqWKjwun21F7ly+Vf+H9D/nXA9B7KxC1JQ8jigtYN5H+3U3unaAJ7JXOUaSADC+3
/YAL22htTvu0n9NbRhQi/XolWVHS8VIzypmuYU2eR7I6naH6GGT5AeLCwb9sJ33NHuwUHaZD/Eju
NhJByXdGlUzJWSuT23pw53GT+QTsuZ+g20Pp2lEW3Onlo55x5+WqUgFU1eqf30eBuKPE426+iNxR
Zq0MIOKvvMcWQWNKlR4OHAHPO0C2OQPQhZXrF8xDu1//aIkHVYmmN/XjmoEWks2z2dfc020W1CJB
zMA57UPS+w0DkC87q9JEmsq2JPLbELI5KrmeQHj2iDSL1WHtzgnNGXfqiav7d8HTxAYARXb+a3fg
iDSfBFGXfPe5rAspu7EikT/oTA/0kO7wo5i7vwXqFEfkCMN53x7tABVKDIj0uKK0ZdHZ1X3jYcqa
BcOluZOZiizxp4zqfn6H3YcE2AkoICB4mO9HlwQHbLBa5lAQqEx5Y+ysiyPtc0c8vxZPqyh19SKb
FwMsq7oPJZOYVZz72heFcUoZVCQJjA4raADyiSPaLPRnfiybBX7ZvwtQz9x0Ou9OXvRRKtqn8JCP
Ja6fV1UCKJUjdyk4lI8H3hQ+nA9DxhK4H6zVh0nKPtW5Z6L+m40BVlq5TDPJFMRm+zMpaDEMBQF/
ic+fLiyvsrt3PBYbUQc+W0Ad3dDHuzWcAdMYBzZAHIwO2CI1j+cwpCRn1/nHsJeBmJeSHIb37IyC
GToDrXpRuDi7bQIvr8fex2zWdX3PbygfxZA/e8pQ6X11/yx10V2GRo2y8s4Xgz+PZdlMFPZFFQSQ
cu9z7aUkJcLiVtYM8XDQ5TyrdrZCMS3TfT41UguhE+lyDROh0F3jLCp3CTmz9ZN3blid/nttDG91
ARfLRLlVH3LqdrGGgGfe4qK8V2LZpnWQhKfmTc1NLjVUYUjtndgPeGEuCldqLbWOSeKm66qmT+/o
Bqelk3tHJdC9/B5VLTCEbeoNzA2x43zW41p0Ai0LHIoVEhgjCilx4pK0BDkm7QEXmZpPi04DCsvA
kkASSftmfTmntYZUfr3mdqSp2EY8cB54KhzhxqssR2UdwAFwLc+p9fPEzei/JW4+mC0yafV3i27M
HT93koW5awu2IfAZ7csw60HC/2WrA3rLqpP/C/44yaDYVtVovr0X7m/F5URT1EF3BZW+0qwuwN9m
DXPUri1jGBn46euKkb/irYe7y+Z5Lv40V2QBz5N+p3THGgsGFZ+hR/0j3sbFmbnmpCQcx/XXqaJT
OA8iW/nYsBt5Y9Ryi6W5PwfTzgrQuR7dPRA7Gmp0Mj5sp9cFW/+goTARaa0lQcw7zKts2vFQkTnS
wC/oFvigxbufzKWuOgVmMt6yRAz1ElJkIdmUWw0AwkVs/IOuBLt70TxF5BE/z+FljCB0bSeTvXO3
ThJJv8OnD411Wco0DEc7n59xqsG1fZlHbdq/cPOIDmV+jH5nTD8tMWZDTjmjX8GM+N5goR4KVQss
dApT/dOK/8Ayb5gqsm/qbR3i0Nfz9tyXZGByeu5VclKSJgbatxCWLSZb6n+ojgE4TlXHAmKvsOP+
+c2NxjKBQdJVSPRZ4XyD2PCj1cd7GjxWlzm33VDIVYVf8NHkbSvhwOCKSJTEy/zt4c0B2NC8XY8Q
J5i0ErvqhZ5RYJhcwmc1bwinyHbuNHdvVuOPlYcbU13dWUx2FYeMbigZTnQGmnVeJxirtLIR6eqG
+dEhA+wFNvj7kkpTOraNb5yPkATA1dH5H+UUSL3ty4ATYyOTX4XffvfCxwE92asVhyjXBIZaUn8u
cqr7Dzaq8q03nxQsuCh7V4U3r1ZoIUiJXOcOFRpSB8AKlu2hRS3BhPtTG5D53d2S/jpLiuODx8PO
IinTPIHtt1pfWrc9dNgOggFgpS0/8IM84+4TEbkON29amNfUmxp8jMy06u3L9DW+Eh6iAqEhEMvO
7p3TJxJ0Dt/EoxNa1um60+V80uUrUNmx95f4V+yjS9k87/fi//u4fHBjJkOOvl/OSY1HyvN7yRPa
NuDOCy9YzxdPdIDKh3qfcbFDN7UDlLakrLdLkSJM0sjQchq5b+4oWZ0xC5wWHHnQqGUJmVsa7UT8
Y4jkvftmstC+yTbWtmvDoLcOw7Af2tBpFGcwYCQ4DJWOUEzTjJCrQLwxUutTecu2QuPPHwKXlQ0z
jayEYgEEsahIu2Km8UkJx3h5MWzsTEctfrx7FiLz6B+81NEia+WIo3jFjIG++pr4I6hjLvUaAJPs
RhW+P9jMpJFtTV/HxbSvfHQwnwIk6Fh8ecBaHwo2ls4r0N6F/YxRrcE8WsVKqEHLdNBIO44mce0S
VSUMKxWrYZ5RtybYy/3SVgp3qUTGKJ/494hi9bsscIRPoBurphfkCqMyDZo6FgxoL/V8AdLjyLYD
ebcqHKaY7ZwxTjczIQsiEuVBZf601mvnEdNUpIikEI/vdb0zHQtIr1h7GbcTqtGo7qnjWbX9zlg2
V9Lko9r9Ey+n1Yvaj1ATNipojsrqRtc6SiDFxQG322vx7TZ4iEW5qP4EB/flLRXNHZ9Vy70OERJD
BVTkqU7D25ZgE6HZCpAGYuqeoBJFIgmh/T5qbaorEC8HOgX599pLN9tzx1CKirPL/vv3HhMsGfxQ
CM6i7VuPprpDEL/N/9Kx0jr2EhC9C/91WqO5KDl+UMxpwSLQ6iQZJ+c3ZmuI98ZBNWer7aYiHJlS
avOMIjbBbCJG9abShcMQRUB3NNmqqLm4wIiOlViLvetZ+3tgp5jbiDoKRDZ98Cg5BfHyqD5nTYlN
A8W0DpOAlSdvjVys6Yn5kVvLEZvEEXp7Hqm8PTv8MFUJl1Td+KPK0iycEltJB/aMb/h9Zg7RbA/E
UQ2rMJ8Vie4umimQLpItfabtMVcgLdKdZOsKM6srRmUB4wDNU1LjTZC6dzZEh1WteFpqfXIKbXx8
1IH4Zm9p3WkdoaaZPASoofOrHg6MoqAgspY9JGvT7Mk0T/MUTQ5F0FwrTRsRfweNvKnjcVkccNYQ
5yHIXKz0t+yOTxku9rQD1RCK2oLPfoi+dQwBj/bCeleYi9L/gZCsrDiEJZdlMHHHoYYPr7iCQCEG
An8gjUnNeFcVQ9aKXSf3Q+yJiQ54eUG1MQrAX8h5FKagvtC3NVaVer3VWYQwDXcuKQazxty5xUU9
N7dbkoNuJ7a0+Ld7fFhsS4caGRTaMsTO4fvAJ2jk4CIvyrf4ybRtHwVmRz1NIpkcQDUrT98sGyxZ
jJ6k684AWWvlCePq8iphuCf7CtMNAsMwg1eiHLnSA4x2VxgHhWpcJwIxWZThpXLlXIFJ0hEXSnuP
BTMFh50ei+x7oGE4lNSsuKWZJG7u89wgXNiyPOvNfeLdQri2lpmmV0Ed5QQfZioFMe+5fQNXaWRo
ULzqtclC8QawTMovcr+vqP8p9hssVkvzcfman6HKpPKR5FX0rb6NwlZPiz0wZzRQJc2HfMQMrQli
TDICDvkqB6xdK56EeUYWw5iaceTZtV9hbG8L64UozCRNrmqKRxd/GSOxYk0r0g62Ih8yQUSSjWZz
8VDjFOGNFh1iPulnKD18pne0HKhAVLpa4x1GNDwSkMSGHId7Ip+G0LEQ1DdruQOUq8scCoa3MLCb
5BrEErNOIsBNghroxOFd6dCassfSb9QXtQmxhsOW+3oJmBYpIlRSpUg+/Kx3ql/GQhXBvVQSVBQL
y+/D/FqOS5zLszanNWdFqRkPz0s+JmyS7KObvs5Cc3CuTDZ5x7LIWslGC/NaQ9VrJJxlEKr2uiOG
sGxn20TR+un28RXrLNTTVY9uIbvF9XBhzPyqNg7FBgxe9cDd2TGKSKR/AGht5+sxhvWimYVth07O
jzeiW6ANUER4JCLarPot8fem+v8yU459HHqxzxAOSJNheqthQwAxSdNqKo8QFDeodrlL1fb/kvrn
OsXxHilB3zdM/6yuozR0ir9rCgI1Qt8fkTbTwABHdQEcGnMkd6j2A2T42C5N/odRjJ99i7VOfbNA
sRLs4onoEJNsJGIqCTP6AS5r/d8m5YJ6L6xzPt91ugXU5CIH8JItNde3+gFDdxDAaVtXmFpXM3A2
aMcbOKJ7GhRaXU+7b0QbszWhT2vfxdbvFNYUO00ZqwUJWN8rjmRuV32SBiC4vS6lnUZ+NFvJb/oc
KtLYwF9o2VF+dMSZFSniBmbt+F0HJClT4RmywrF721ubeQ1Tf3M4DiACyzeSzQeIrofuvYHP5AgC
ba+598RdRUm0T8T7ZyAY8Mx+7KfhhRt0Lme+dd0Oq4v6Gk6K5jbHS83VqfOcPiIeKIuooZUBIANB
KkoODSN2Ck6AfQt9hKsGUvEJOnM7eAwzln3TXqPd1DPTVuv6f4uO/PGQnbZfD35k4uEzEsI89PAw
lJCI55OvKWehtMVY+UwyBrxUVhNcppBPHd2okCUj8RpxymvjHmYgbb7Byqgy/5+esBRDFX5C5BYS
+FvjM/Faax8qP54QQqQT43wH7hxXDQJWu5P1K1FUEJWcqPZ5e6kepxpTzvu2xkHVjEa0d0PViOUi
Mlhm90eQttbY+k3IyYY6u1P5hs1/lpocOpprU4p0wjLHQprX9Qi1v+khFEIqQe1DdrmgUjsTaHnn
KzrFg4xSLOgX3hjlnHhXmUul4gJrWWHNpv7lLiE2hbxG78KsyJPIOMpbkWs1lHuo4JD+wizFM4Wj
kSaqkALyf3u6vaf5ooVyxsOB1S7N+pyWKz68EmUgkZafHkRT8IpAN8LCZiwR9yZet7MZy173J46r
Xs2QcLVTY6WpY9HqoWRdGMSAp9TSp6Ww6MBHo2APSo+iw6HgFkYhg+DbnQ0FePtjr1laXo/Noa6p
bqLQ8FJrvVKw8lIVDsYGa/KtHQEzs6+Gq2gFAPFvxLIbpWuugkq9f+Flavm+Hml2KdXvZStCiD4z
ozE91HkMVcFuhGoWIRYprJ6NQ1axYi5N/76yhZgVV5FgRc91WHRffvwOXuYNm1B+FZXN26ud6p1U
OAPwT2vRHzBML9YIwsa1gMHmZQKiY8VzWPZp8V9hqAfsfOJaRtXKQMgV3kQaxRJSimy2Ku4oW+cH
aA6HCn0Vr7brv1+MPLrLWhkPl681pn+tkRs8YBVvjZO2YQTlzuh2QA7VuTGf1fclNnisgAMOfHNn
ibYeaZDqC9I5sQA77aRTo7yiuG+iA3Eae5VNreWf79/Y2glSZs8sauEAMIHQt6VPuY+AatPb/k4k
xT51gDN4Hh7FF65OVxG7KN3sEdOsCBqq8EUdoz2qAWu5FByT+Fgn2eGNnN8QxV1Yu2Evq34SE2OF
A6iDXjxNgbMpf5FK8bhxyBZGkZgNZ25NeRoXXTyU/5hEmEGBxsxgRwNJUqRNhdTKQVBc+fPFq1xK
d8Mwqe/clO6k4aCcxBsFuXdiF80hjA20nDLspSuFY5kg7WzrrPIwxunvUJ73P86BWzSR+L48Dw5t
b4T5W51++LzE8R6DH6WG90YOc/SXtn90Gb7hvbz9PVCDIj2CAHpbkzNooUYPfVcwv/2FvgxJjEDm
VErg0/3ezN56c6zHwzI+nm0t0ZSqZ5Mitdzo/ZBcXJNfxgTvzBbVyCLlkYZxL+pbaon8SNQaOz5a
FpHxy7+THGTo68l4qq3yMbfPx+jk48yqD17Q++W78p4b2xTabaL4Dz3vRMRfGEbm/a+n9ZW/gS6N
kODjSZLPNiGxB+QYydqb0ySAgRl3x+1dO9+uLnqVPoNgH3/AHkeI6bmfRBMkjyenitMJn3SRHqmV
UZeDEsERTMGc4Z+/mvEUQ8yoZN/2B9UUBsRd8JDtTNvETvBqp2kzfXIfp+AMqIC+PsSPNld//wXx
sOzjM240V+T/u84ce83dA4K22QHVWYwEUPfuc3L2VFpn1cTBvVkT8Byv4/cRmYNxllzU4+hfwWtK
1V0jIDfBcXo6yLCs4RDUuO7a9XB1x0SqwrrwYXvW/69w/tvqqWY3lwgCohAqSTDwwigkkXZqeapp
5Fhys3qS2hRn8smxzkrxU1hN1vqWiIe1ePdqaEJkfCLIe4I//kTQOvEunjmxIArTBrgATu9CIx6W
ABvJPVnfJhlHrAWCW7Z7NGPVaHV4GcakndMy2eQOtn4qYKNyzyARzm9zSs3gLmwc9eJVzKmKofJZ
3c9vHJosbumVkVimkjGS4CSBlimVWqUK4vB0fItDlPBR6Je7Sh3EEskW9MFs5HktE4RmQky6WUqA
AMdBtbxuPBytYcDYEMWME1Ms61LRVFO5D30Mm1Wn2YvcF7pzPuoNVQttPsISqu+lUco7RQD/jl6J
ssZhBV7GBGZNDFFFkmKzflhZ5O8VpW89tIfFCj6+xaxflT+TCKEozGuE++yPSczyZNa4Dph+q0+6
Y5/P3NKfJn3ei6MosxohGDEz1qF2s7IAPZv/shQPif7TbhjqG/dfrInK1JCECTGsac/5RkOxqHrD
qvl0kNE63pXZRJ7yjj2HgvQJLmnDvz5hLM54l8J+uakVjdyeaWmug56mpgf92yVwnvH0ChRkAG/f
YyEZpy3o9mVfKXRTyQzgG9orLU9FqdxgvaL7B3ntqNTqN+KebmS+uIeNyc+lse3KVD6LZ5afNNP5
t7Dmlh3ZOscKI4pEqZjzxUY4XebX+/1ahgGEDMtrYFEr8yu14hhN/xjUgpRiNiaWIS8ax9sMxHUi
oK/gDRu2dF0/1EvncAmU8JIKNkfvegPf11zQ1Ryd0yJuBe4QivhNG/hzq0VepP9hviY2gURklD73
8mhgWflPldb2snQHUUTd75LOZ2YyLoheNvTl60ILinMBWgUjeFFzj2x94FK2Mv6uMnvJS11OnafQ
Mc2mrCyTOQEkGfPYdVvvl5Z9RBervAbsnSQVimekI1FMujajSHKOO5rCaRo1O6L7Rat58Btx8eQ1
bcuKVpP1bWp92nQX1O65Zb7k9CnybXHXDgyyP3aZyknTtqle/5NxpSChPzltjzJiHXUenlz7BGPK
25VCsXKxjkVH1Vvk9x24HP4+1fwqmupHF7TvD5YzgAFf5RkGu6D+x+zY+FX7Kt5sxIa0typuKS2e
9d0czCeVqwEt7t+fPr9aezHMVehNOXH/UEckdJ1RVqHs8amYt2ZDbb6sfutrZSYHCAPJ/H5BqZ+i
SAfHRVlu5hhTrJWlJBzpQHQSU2g8fc9T+eJp8FIzzMTa5wBbcFckrWMAHfeqxIUi15YerH2kbJ3/
lWSOC75h7RGR8lFOByBX5O3wILUvFZgnjwFagAdVcJ0av1kmUg9Fh/cET8+siZGR5yEDZ8A9+Dqx
joGR8CLsnOel+txqOsVpsLUz0dIEmdSB88UaKE/h/jWFO7pfFnniOxRT2NJVzQpfrjp2x7YEl4vH
BD0m0zkY/ZrOjsHTtyFONhQo6vOUVE7uc+ub1pxLya9WEz26LfYCdJkfxOocRD4v/5T/PmKwmfOU
ejA/QUaf7XfpVJMiFhTZx5zXV/Cv8DglzuR2O37UbGy38DA6YPrELB8hvGdmQ9S0pVp9+7NWIACO
QQjOAbeztntsSqSjr1DnOAbmqHZiGujrMNq9TqHIZl/DDI1IRxbYWyboALhlKuExRrXZsUwMRfPj
zVTklWJKoAaQgheHbF4pjdvvSPAfLYHcfvnRvOVzoyPalU0Gcn36cJez/3WQl5y2yKjuo22Wus3g
TjaPBcxH2Ai5oEbMGAQHAhcHVAlsqkcDlxC5XXNouAPAzjMDOLlmHJ7S4XFM9tyyndyIYB4wKbwp
qws+p+AFhyO5uYAsT4n+KD5qwDclEoerrDzx6xs/hiGM3/qFNAseh9vflQ2A40SbIBy02GJI7wvp
Vq6X56XJA5mQke9OE3cG8+C14w9OkF5mzjcw75isZ2GB2/Sg04b3SQWOA1/rCQEPMKh/Mm5VjWB8
xathYhHK7J+kmGATy60RYYS9Sd8prMe/dsIPzGyI9CwJLNjULlnXiuHaDA52w2Vqhspa5ltsat2P
ORC4jrZNEaOBmKnqAQinQAYS2lCidpQxDG1VL34AnSzS6Qe/77onfG4pIIVyffKCxEW5/sa5RfZv
pK/b6/RsmO1OgfPFO9mGMSCY9oFri8S6nVBaZDwLop91Bb3tFyKQDnws+8+LvxBM60LhhUX8YVz0
7/EpfC4kgFehLulPfPBJhDFW+WyYRw4rFa5j3DQmvuaZRkruTkkNYj/hQVtCGxjhc/BzrJXFEky4
BIlECRLf/sKvs1NCiGwXpRhJGoJEwdj8zNCNM15gt82A14jDgrPh5dLY5C7UI75fUcNlE8ZfB7Sf
YNhqTHfkULkRlizaf4KC39xN2JMZ1sGogeSGj0bm/O5YnAi2X40m25ZjDrI5FFS5oWd/t9KdXfXB
PB8Jz4YK3brOQ/6Fewp0edMIxN0lJaonMWM2z+gKJLf3tJum0UWSEG+WQZcoQZzwvq85Ob5gRKvg
2XAGDSudjq+gUqoRydAg60R3U8Sk33aul0zIke4iL34uiyk/xvtUc00WcBJmJo8ipRk4dYvJZhih
Vip5LBnePTeHwSGmPF6WPCIfBMVwp20Ii83qCPsbXXk8ZBpxRgLTxAiaZxi7YFupnrOuFaFMmxDr
UYBdGFgn1yMC4og8OWfasYRKuFQgVYeDTOO1tGVgc5jfSr29cWEz+ytVF1k38k0ztunop7dfxl94
fULPW4wbGR/+yYDwIybGHvUDV188RqueKVRqm8xm53kQZBC8okFCMVKgLZopdH/d7Uy5o8/t8YES
j1M/zPAHzok/wqJpFH9SEXcgsnF9xAxVNavmx1xb8B7fnd2qh2f84PHpZMSglZmWlQW+HjpUtjWc
TmHBAovUA9+hWFmWd07/6xzk2ekY8m4cclqKoatZc2ohg2R13t1BQtXn5ouNtNBWEuB4rO2aRTwb
Impfb3ioNclgWkg3s/YFYf1AN5MiFgiFeNJFx3hEIwbx1UE2wy0JEvtcJOZoYGa+rYX5EAbo/s6v
bM6Y1cUDZGGSaKoaw/YTE7mZL94LbCsUAfa8kuC3XkfArMhXVxmV7LHqEU63E4Yuu33hWIpMM/bx
z78m6zQxGJX65dIt0O4fjrg0JAYvmw6o1rXo8gSuLIlZPjpuIs+LGDT+X8gDvgE/ZB5BFm7dROZc
7BCIVFp7ceKt3gk52wwqZQ3wMDlJWFACtl98rrMVizj66ibSsGTT1lKvEI0xAV9ErrqbecKKAwRV
YWc8WYGntYKGxbMRsFvpUhov9R4lFPiqMkaOdexj0zZ4B8FSrfe3bdIgpuqxdGuXXz836I7UH+bX
oH7TUpx5ojqUaMmNb2nIfxcUUaJJTK5runQ5LVmTWkZRDclhM5GaT7r4BIG8tqNSbBnqKU7FFvsW
rX5vXIfv9ZB+7sV/NCwQiIpVdQb1TeOiXH6PsrRmlhRjYvEDrHiD0uvm0IeLESG8Pz/ZPorS26kd
JgYtKK+BeAWaPu3yJSjP7yiaG1HBnN7U68r85LfdFwgHbO/QRLoc9s5/7VoiYMAD0on6ZgSmAFV7
Ct2rBIhIZR0XgH1LO7xigmOaP8FWfz8wa4SMDKUtEeuSFx0ZIiJAVjMVWdKbV/QIsg/6WV63et/u
G9f5TCw07x52GQFPG4WI+brRWmCNZz6fm7OsV8ZsFxTuzoThdd9lw+M31VtGAM5kgT4z/ccQbiWu
enVUjAV5j7fgZs4vI/dnkU+MZxmzaYfxxiNn4sdwjte2r8/lGLwqIrVBHm5E07i4D6wlIAoLBusa
zzr49UBZ05TicGzCbgIW+OPjtZp5Cfw8v0hd6C+CkULmym3tDysx75/K2vtl1Mv6giPDNBy60rvB
bchnMNANGQqZUxU7fJO86/PPkQnDw8hz9fPN/2V1BLIJ+yn5eXONOkKaabyQj3PLByTY0C21UBvj
kQIMCYOkIvkngBCY/m6JDvhR1nEP61nva3GpfIAqwLhAR5aJw39rrurnKwNPAB+FpQtEiS6cEd/F
or6EKiI7ncEBveSTQgdSjxIBQ8LXuPW2GAZ6Jxw45jVWtoCFRLopzAjChTGKF7GvCx3yTBlSZKaK
QDcQE034fqNvAAMrrp1Y8uFF8TtG1BrrWn8joZjZTf/L7iVvcZ4Lq52peXC32uPdr666S6ctphMN
y9q2w/xyuFc9kb2r460J84Dc54+usz77+hJo+nu+VhwcYnn5I0V7f/e0QqKTtBDQWBphsLU0D4MM
hIG3I55Pfza9hvrxZqRahmBiQtPVh2WNwb521D9RJrEMXtnz4krn9ZW9MYJ5jQi65vbHv40rx4n3
28mRyoPiVYpMQu1BUQCB40KpiIxu9KWKvT07VJ0j3TeRV5HhxE/lZgcHry3I32ZijlJGs27bB7rm
dQXyFStYnGlpb/soC8dOD9JqWpHpxA0r2Pu2ASWGsBreaap7wC0VZ4G0+mYD4/g4/K54CaKfVm6i
aFMMXQmuP58mJtD8aXccuD+b/IUISC0n1mwF9a9PUK5EQKhPg3T2NXAzvo4XM0iFC6yqB1eJDzyR
xNrqjgQTXow6B9gKuvJO5w06T/LH+b1RaaQRwvOv8FTniJpWn+mwTAi4ZrQ/BOQdd3rvixDNVB6Z
+4zvLvNYSkqQjEVABcaKVNP9oX++IBsd3Qy6GP+ApmGst62A3dNwlKulH9eGR9cLATKgtbQcO1T3
mJTG8D8MPE5QzWRknq5Sc1y1rfSO4zFo6n1P9M95ekYpaJuecFjQt1QbfEN2KPFvpMWbPrDFZ8cX
e3wKpA62Lavq9S//Jqwhlgt5OxvhKwtjXlrO44Yk27qATHuNlIEry9TWPqh+UFJynZZwJgavF+Mh
/B+MBRFAWd3YVHfnt6uGQ/DCGIPEvdO4xxLEcKPPl+9TWFzANR448mgzHMXALGbMm5t+8x4IUlWB
bVj0l3HR5R6RP6OVOSoQ+nAphH3QgXzja6Y7EAAQzxDLvarSg2NeJC0R1sS44RYJVVUp7WX5qRO9
H1+HTVfWYKiY5vD4vN03E+jPHTrEI8HZSLmBHCGoqU2T0SE7TVdrmLjfZH4VOHZBEv3vmu6tdZr/
XafoLxzgwXmqnaWxiyw+hRn/DEhxrSZQOmwVfWY5yQawAWTQUqgMjLleltXmqWl/h0U7VGDZ07iT
bpT3loR+ai4YZM2jCEakVS63TApS8NKgKIoGuw53/N3zlKZHF9tx1EDMcbSlHd8Sjdf3Si6SsJXd
Cxq8aq37Imq3ZKipLs78hspxGeNLgBQmmRfPYMUytHOZ0h3VpkgYfq3TRKEB9wW5jzJenDNkusOj
WqI0sQ9fCcQ+vfGPQkbMTmQ/UFSv/w6rjAJ4+gi+vNgm4mDU7ugMFvhdzeErGYcmGzzE0sSmmPzw
R7FNXcf0IoJZn5kuWk59jNH4yKEP8dWZtKCYvYMtdqZSohP6S1KwLkwZzN6UbVzoRNlW/deX/aRQ
qM9MhbmRA3UTYwy16OyKsYEQLyzY9Y+eLkr4XpsYItbAgFszt7nUbz/Wq/bO6OSlwgCrJ3Eg2POd
F88WfqTLJdc/XCp7ZYyw/wV4l/bkEo2C5NTFOH8xDeBRtviK35u0m5MAx9bWHcZPe6QMYdT2XvYI
WbIRmsZy2V4cagXPh7POSDUxlluxQ1+PVOG7vKc6Aos63hJ+D4pdA4IGAwZktejb2PHhN9588Yaj
cWc46gq5/1MWKCBaCXKUvVQL2Q2pjb6QlJKyFq8AR+CuhP8soyCx0WAhsbe8dUJ3HoeDxb8yHXX3
AnQ79A2pg+wJ69QcEPEdJ+nSWDKij1Db/Q5XGz+brLn/izfquGLzslGRW03HLB1Xcy5PJS1+APet
r9R7rS6uWtSoe4p2D93g266sxgqvqQFDvXrdYhUOdLPDRj9NJWc9kAVNea+P42YGxH6+NFO156Q0
n+cmiUdneN8Lare5Q9KjVmaWFSqfKUhdLoSf3HMrGPkNWbZrJTyboKyb3xjUsUmNMtzZ8QpHDcQW
GZ3tJwXEl35PQq2HFwoXh3G3u2R5Sh+FBkGYsmdBeb7kVGQjiISniFZ6Y4udvHopOvMYGBeeTVLJ
5tEMfKbbDYFTruChEuvDu4G19WQMWTml1AxMn0xj/87DOnpLuWe4gV6gHvAVRycw8a1mtJaiiY7F
J+TC/vwZnPsvpW9esUC2urPFjrNUe1ALjF0pkGPIou2Pvb9DPuPwZ6AyN8o0lOKLkRufCvFLxQyL
CdnRs0x0ksmrqycTmP/gSyC1F4m1hgPQt113f90FT4I4cODR6JEYEi2LXNrYdOCkokSOb3isHhLR
8Q80Vl2Y3tpbKR6JYSBrH7S9LqH0Kq8gsO0aNklFy169unuQHL787ihm5BO7DDqkJb8onnoSW3Nh
8XMSpPUMPiEhMPiqzaH/9YxcFDmQ7ulUO7Xv+gCN1/zoa1JcNwoA0iZwjTaSQJhFoxAH00VJ1+B/
SVlOfxNXMXDzqem8yWbDoKOY9/KscqTThqIvCfpEA6zLsZ9PjldFkEt34Y4h4T3rGphseT26jUDx
xWTesuCUQILvlcokZCmO9sEf2V9rTRQQtyE+h9HAfyad6qTVSTYZgyzTF0S6SA2Ov1uijeKColxK
nkKrTiY5uKgVSvvvzYhrlMAsZTMt64UH4C5P9tFCP08mhmvzCx1cttwAB6E1YBK+M6Vjf6jYEHnG
VYtSnJwPw0Jwtt0ZtQM6+3Oq7FlZht+XGXPrY+RIZxzsjorh+JnSGO5H+hK1RxzZy28US4wewmk3
7JlVWU5rjxPE77jQES3EJON+91injcqWEdLQ9H6xatvKfd1mw4cbSZwsCVR4XqhZ40UNYwpB1274
dJVVCNcRoe3RcReE6I/aURmbCaakUXov7plMPWs+43svGs6LBMc+rFefuLFlkhaOPfn7MdbFFOZ7
7rFxC8X31FvGqIcgqly/eKPbTfULUsI1R86mbvhYAxA6LQkE23X3xsWL65YoC7dsBIZGyVCO+MU6
csv77UX/JjVw3+Ix/n9K8HWYYNJOFL1U6uNEhb/Ebm3KG8vRP7G9UeEkIey/sggdI556/8EQPxMI
i2LZrQ+6thKic6+mUaSHAAVVuv02OkZphyAQ2ViAQ/RGxXSrdRcB/IlwN3mCvg31g7QWDViXU+GR
s+7dIfwA3ktRehTXbNH02QmXcV/RDOJhaVll98PLpaH9kU/DOj9sHzBtV9njb8++xcVShrlMbl9X
bty89uJ+HywSCh/52mGYey8ThJVZDhk4iNBFbYjVaI0neM1Z08kJOzNelwzzMd979V2xud9KbMEN
pNAGNRJBemSdaAfh5PcQsbS7NTV1I9d7AnPhCJVFQizrVd8jsl+gXx5zcBbOhJl6VcQtoyz9kNLE
Lh7GpAfIQDb+92EhyQIItTMNko7u/YqHt6qaM2jblniNN9zsRhQDErgaR0k6+Kvd9aT2jrg2DHdi
/DRfJWdalRW3hLLxSqkRpYr3PFqUtSdj0DY2In6xG+y3kZoUacl8h004YQ7KnIxagrYYqtRtVoKx
HSGbJIx+aI2mwLd3Tk4w558Rligw7J0csTcz1Lu8JYv+Kjv8m+GWcCl4hd0BwzC2AmpPKvjfJbgY
XDoJdvFc0f1XrWNzU3rUIueAJf1PvGcd9acpbIDROdEXePnDaoDWxftKfYS9fMRrevILNyWNy6qV
mDtBnxuKKabjv//GtXMEbke22yWlN1zfnsiBzJIzXAPFqvf/FqxOUZ614ofqQDZNbLe9LQnSH4fH
pJdt68/TeAVXfeww7YPDYQsKL3ep0aQPpNmXPfiq+w6B7XTdLqHltv4HI6FBZMJsynf1QPBq7m/8
6ZS7MXBrnxtoWoktrhRTR5x5gj/yiunJFQAPmx0bv3uZXHmtcuPc1vfK9gJf6rh+MsxGDRhMGC5S
4PVtzHu4mlFQ/Ar5Q8AdI4p1g6k6JVk1TpVmi/nM1hRVl75i7thQv0Zaax2P+pE6cNqOb4w6us2G
L0mMHwUBRfrKn+3QzXjnICALScCZe6dw/vp5wPvSEsTYywqe2fDrj/ihZi1rH3r68YcMA8VQAeo7
CfPPy/0heK8E5cle4PuyQuS+t95ITXXzoufkvlVKqA2U8aS680lEY7x58K1ztCnQ0INcvoWfzQBy
7kQRrfC/BFODLGZOamOxRlV2YBllklCHvZgiVzcTwJXqBVjhL+W0HfawmVhkGBV0NOnRHGZFyNTW
yI/8jXT8O8TVZzQIZnQmDyRhvaNf1zNmbKoUgO4BviASOyTOoRIoLAnIjt1ATu+Evs9jRVU9NJ9J
Lo3hGqbmf0XNxOT3gul+uVoryASIDKRosFVztBA3A5rFiOS44oUGT0YQpeO8lqmAAWLaHGSxjIlD
KyejdHUWfyXGZb16nPHs7RGgEda+SSrYTG7zKgjWBn5PvSzB2UdV5BG7StOU6WOLXgv3O+LMSlgH
W/p/iNePlB8MqGdhvKXNsoV23lhSa1qwOcCsnIfc9USkJhfm2OR9/jzmRjY7sNOSwId/EZyBpE3U
UhcW4ZyEAR+LF87R9CEi0BUkY0e3kIycLWxaw5q+cm4OjezJ1fjbYjnz71g5SINrPtl+p61wNrDd
+MTZCraaLOaOfaQyUj3xgXIxrenP5CAh+kho7+1cZAOwxSPiw/fKARGXhAvSJj8ax0GmVAlG75rG
vZtE+gQdQWTVh+WIJvZcgO6Fnlc/AIx+Tm02b34L3cjvZVtr3ZwwBVezivv6tlRbeRN/OdrkD0J+
5YhcRlhhdq6AxQEkf2bEwv86CyNLQaPCZ0oJIi0Y2FR7bjRmSDHivhIRTpsOLA3AsCk0O6QRSCjQ
/f3OnCU2dnz1On+QEHFWW3IfFmwY84W+Lx1nuIAKGLuN0PngZMaQ9y5KvZVRdd3/89cRMEGDkvLX
G0glROnmjIINERu2yeryHBJOUUZTPhvlCBCmMCgVkFPWzdFhyWYiq/eQp27mxAmV5SwVaHStU+vZ
l7/7VQR7/0ncFQpXsOCuONOB2h7ETwmGsB/2mxTGjjBvE9kQz3dFPpVynMHazBYoG2WFQDiNQGrs
fFsMb9yxNo5TiZFUU7y6HBBka3ldgob03fuitLlfMCjYudGLYd8Td4UwjGmrsZWB6yCPDUgHY296
47V1xylF8HZMRXOgbdxhwgUQGVKoJOiqLo74jQc4RkE5s5l9eGVKbuPxU8L5RVU2NqqVD8nMVNSC
UvcksHw35HDLifC1PP1IXhIkQ3R7JAhzOVsQkidGBunk8ss6dJMIs+etT6OrAWt00QvbFxEpXJAP
BUOF8LerDEE1q0z1cqwoJ+j/G2dmfIMQoBcsqimOd+lzYflxhM9QgG9UU3GeXX+a9xCgzpj3R5dL
YMcaGMvenJqLmcYpmVJwI10aHIKYfUFYZ9zyKzz+bdIsxGASp3Pz2x1trGJHUu/3BBWBuGk0ZUx/
p8n+VLtQRhEwCK+4DLDwx4OEk9ZGBrH9librqrQZqUYiACrEhSsOA3l0bEIFaNY1wkFZcEEe3VcM
uyKgQvDcOR2p0tnQjvNk6OKOrapfdA4IKfFT/lhHxideQMpo6mkQICp66zmZY97vZcl38dVwXQRP
Jf3rhRjxlPuy/0PbsVmu3xjGNhVOQYNt1wOMvvTuEW/ZOFg58hjllGGGmuQzHegLDZAqLxghKDCN
VO9ViWwKDrUuWYaa6wgjtfraoEm0V/7p1LEbIsHjkwNzu15qsAs4x++wuU7obVuqFkYv39d+tDfq
7rl6hHOP0SW1PhpfoJPk5SnVazAjhSuhwkX5LUVTrqaczXsZyTZphB8pZfbPD646rFI4bdX/PFuq
EebWFC5P9XfEcjQH4e21nTfFq4cDABXiBvFkwc0VyxrRPGteTCrZsKghPoq4n75RApvNrzGcdsOa
OC6C1ouGUsFakaJpWo7z+T+Al5G2oXdLCZMA+ioidzbmSWDOI7Op6p1aP3xEbDuaAqmy0ushvFao
eTNGQWydyun3Nn9cydlvJXUHotZ64D9Yne7GUJbdsejjoLmFLd+rekSmV+VZ6UvlGZRhvK4tUmpx
XVRhO3uhEIKwi1CB3SxYRjun0p3kUV+Rlyv94vIHMy8re+avHQtKEBLnzJxopfv1Oc0HvyJgSWHZ
2qJEI27LHJVXgA5F8GSvSWEEyoHMondBoFm5LvpbxacUTiUrQRxjxPIDnooZwfk4OjWmVe15FqED
Q732ISC/VVgYprcW8KFPShLQuAA1j3GPJHkOLDsiem/X9xJSm/HFZSSbPwWe/8UwOrlMvS1rNg6R
zTGhpz4uZy9m1dg4zABiCTGWo8Q1F4TMMUdAeJseoG0ZiEaa4goC7kKitDclGhhxSB51RkH0lMhi
cJ/Q/N6P0esDiupdjAPo+cpHxVlWiR6wW3HeaoUp3PKT5AgRiN+GrbTQGPVdb+rYUyk43HIy60k+
7Tw44VzAX2DeBueLlJWfYi0hh/y4SKkV6BHifbuzUTvpq8SCHpe6r2RPurxsakUor+dHkRgofft6
i7XV9P5LNDhF9Yna4YlpMPuI94SAxwvDYYgi+6A41AJO4cgqdVNgoIZ6AuFFi95u4cLtk7Snq7j3
7bxcUpB3e90YgKlZLd3dtcpZQRaCyTYi80NI7HTRS6FA5MmavMKSsEEuirtsp+QMg3aUEf8ULYbw
bV1lxCukWI+GxWARLdP5FI1FAM2gvPS6iyoj3/8h8ZDJ3UeCYMFFZl7yqYTD8nCuXhViKfsl+Ao/
Zx0LPPhOfTF2z0skk6wIni48GcHsLzZVAvu/AvnUDGg43pfiLKKi53C0CCfUVu6RqKT2NxMNmNDZ
X1/jsTKukxC0NpEK8katjUFKNannQv7feRp7KxHYuAKJHx0S0rz07LaAiKz9ifgzod7u3YLxYWsp
cauzAMdj52Bd/p2D3ti/7uZslJ1Z4Uo36tma22HpK6Aa0ADfMI9nzySUmJtkIwKdDrfSecGooGDN
w027RDLmgDVE6YSxaurtOI7ltrcRIptEi24z2B5Yb6HV83kCm7GJjjo0Sxxc7+cQalpB+4MDua0L
8otbcr28wtfJzWD3Mk/IbHRFild13PASrrXhKHGvr1pQoQr+SZSWjvso+i0quaCMD5TAVADCDGo6
0OyFCaz5ssbgrjpZ/ForxGBMAROjrA2xnR/ufFutg90R10I/4W9QdZMatPfMzRlE+lesL4M4QN5A
4Ie9JPYqF8hsI6Qf5E36gXvIeC03bZf8PkPZqjC2WfVYlLJgkU1+20r7rwq5aUpjY9fhlqn3a0/7
rIJsLSWEWW1oCUva3ikGjDnTGyFBPv4J8zMvh9GL2iOazSTarCuTXO+TWOUteQ2eUbz9h1xBNE9P
Wkr2nVxf4jvm4G29EBk6G+3J9oW9FU4mqKNn2l5v2+yE3kr5lVDFwNLyTeTaHegjixKbJwdFf+Je
VISNzE9jogHiAWA8tB7W2nhJjFh1tZAiHbEjWnP1JS3sokVVXFyOpUnGi8KiovS44F5dMrj7dO3t
d96xVZ7+yzvnlAgw5+nxub+MdaiaTa0o3NvBH8erRTWtd2u325xp6JPYdVTt+RAqYg5kklV5nZn9
AxM12ocPoqrEnz0LjGwcxl0vSw9UISOn46P5Qj28czG0eQyGxEnwwxJDWJMDt2TXbACq74DLVHz0
cogeCKmJ310YHgFU4o0R7sqNJn96Yb8mh6yhYQ0EIZw7GhZr4lcTqN5Qk2DWIq8SZwLcO/XQfSdw
C1HbZZYVOEdPqKUCyDKdJvtl2HwPX97QL5fDbO44WTQIYV9E3+j+1ZM6sWjLTesIrgRFu2QbG6zU
CQ4Mt1BAZfVQ6QIVj6tgqxPhW1nn97dMyvAxiL/RlYCc0vPAu9G6oaYI5NG9PT9xJndPbpUVIhI4
UoDSC+/W+tufhPODun6dD3KppMCcZTxD03YOpOflx7vx3prT3R4/yiB3GaQA3dP3/xt8BiMpc5HQ
fDgWdSIDit4JUuRU/lPk+w8dkbGXLCbv8BD5MQgG74oYvixojChmGT/rnMULqkNxzUBb7+PNurup
w6iAobkm1lhVOUPs1fk479VHxYPsvp1F2x9tlQg2YO0pZI5vCm6UjOHcH8HKdWA6+urDGYbg95Sm
Z2JKavNVWNDWgv3jW2F7QAosmH1mqeQ07OguLgpIrUorAfhXF2ic5/5G0L+4+2nTAS9uOgzmjN4d
8q8MHvG0j1Pz3COryQZ9e9LtOJ8MmrCklbLvzeDNmxR/w0afsHcJYkAvCqDUuZiMpFodyfuMmXy3
Xs/AXKbZNe3Ozgec/8I/eUfr9xBRS+e8+7GjbZ4EBAva9U76yHRKjIcdBPUWZlv3CwxySY8H+Y+F
BvZRsfFNts++yWFzcdecItUWkFwMRxaJJ1AdjSUBoAjqc9k4Vy1RP9fPwF1gJlzi/ruGEsu9eDyr
a5pTSC+/v76LdAcKhZeGhiXrK4DEB7oghjzHUJ2KqZ1/W3Czfai0fBnmVkiiNwKxl3meSTO4UrmE
/vUutEDxPsWI2Kk8swFlTacJ7T8gEYGKyZQe477d3EXUWzltTKraZstQz0/DgQmXcc+sKxGy+yqT
+IbyOcPper0CwnVYQn7SAjXatZbSkFzp55mfL4LsYUNHrkIHbev/9jy5xqaMyJ3fMkdR5RU2HrGH
9+gINHJ6IwNqBLElQQReyiUtNIfEjdPVPxiWzhWEogwpDbmSU3IwMm8HD/zHhyLtclBBRpTKJHjO
Ct5sbfaVun1T/WSYepOQ5lxbwOa11cf7SpBNBHk+W/BbenTKNjgGZClMzW+EdIV5kAmJh90vQ0fy
VJk/tY32gNpWiqdc4t5evHyAnptAS+LGghFDlTIQoXIdgwV7tSB/i4ywMJgGNVweQ+TDpWAEZ32Y
26PAge8ikA0GaJN7ft2hlBNfBV3Cv3Mb2h1zzxfqbJk2DKMlxg/fJQF22EfLpLABAmMG38bvJZof
YMIJTy42PItcopjxaNWJ0pb6BuuSZXdai18a3goTWQ1IJtrL19qKfJwS7fU/Ach7w4PBl4l7MUKH
Qh6jMBQxp7TQ1TUYpPLj0N6xzDbe4xxTh7MNoqDFDX7Avkj8qHZyDHdXU6xFOHvMNjblCBCt1+OO
rnlxpQwVeXeKylAmqi0HjCWXTpgadhN73atbNotX/XbCN1uSVJYvsYuvZYXVekCM/bE+7KZ3gXPu
oUgB87aesiWa8oXGn70zR6PoEt4dYzwtl/pbySAOJPqIJemIyqX4bhkEGy3lDmNmYgkl9FkBEnTr
7/wYaBzx1RfKZYUU+z26xmx0nG0XMlv4G5+BkiKhd4UfupdY+fnr3SsFSBTxkcKw9wfwhaqnfW9H
+AU+yzuZ0Vdk1GX7LJ5by9KHNB7SGwDevuP/J7wcnPepMpvaaiRbOAE10PgFh51EsHSh70mgdewW
X8YKHe/+RAAmn5+FhVxmTZ0iCxdrsZJC+vZr3bGW197vTLBy1grXZaYS6QQI72d4S+2nTPJFak2j
H9wbor2Qn5LDOdr1CwLSs00UqtcRD2/4IPZeRNj7gQb42qfAOk7S6p9nApfL1LDfwmTUZchoxvF2
7r5DZG1j3qesRzHIOhfyhngl7UBPc31n8dGqG9S+V347PpSqX4LdP73vj4eDNa+rpz6y+uUWvQBu
OXSJzOoM8sF2sL5iSyb1FmEJf974kIysL4AnYuTsm62jfza2tm8wmgoJrurr9xA7T+fqus/F8PYP
pUjhkTlNEUaMp8vC1TXiTVbsozTMhXJ8Nfa3uwqH4MgljueS/JaxRulDAZaITg2hyGX/ilrESMe+
VBdDzSB5WCS2i+vdvt8LP0edEcl+TQfHb9v28f5NecBWc6xDa1/AMYxv0pDeAuIgEzL2jZhXnpgM
w30rF+gVKKkNGtpyPYiILYUxTOvPnIbszRhmp9+0VMMgeRgWTG34o/QFeMplvu4fAymh7BLYs5kO
mMuN3WAZvtc6K6nYEnF9BdqVs28bGhXVt9JZVpQdEiFYuFdom5DWPafiJYghS9DrHbgQ3o9lTIcP
jtubmxUDTxkQ7jTwrEOITAw2v997+8gx4Kphdp7GdHbtpOce8LUTMsxbERveBHbkd6oTNAeaURms
1OsKtq6joWYMvcDxC42l0krOHKQQuOzjGFSl5CMNVeJ5RUBEUfwXEosLM87BFvIVH5afP6tH0G0k
HQfeqslIZGUnvrWAeamhPJxdt+RDtaMPYCwOuTvgRaaGvFdClj7XZHMcf0aEfOgdKkclj6lTnAbv
iawsUxkpfTQjzRX9QdRVwma4d/jNSSwKGAKU1MtqsbsZS7cGYOBHzzetQqhD9gaK4scyxLQ02C5U
vPm9T/XAlAy6xUko7EMyeBUOGM9Gzklzq4qWdFoqrIn6Wj63aGuIzEH0U4DgCdWEffkojKgLeoEt
aBp0wy7vOLPDFGXRVFujK/NZJL0UwvtdWi5P7S1fTmLtLVn09RfBKoO2fDeeGZTPFAYJMs6yB5RC
WfpsxXNhINPwZ8+WfeyHJdbltTdC6Fjh0OqKKWPBd+6suZowUZF7pq4kYbGRd3c1jZDCXBcen+qt
D6grLgcpuP0pOuoyooB9JAZuuWs4EkKcg9C3Q87RVZUjnayFa4OTC6NpTPo1vi9lYJjx7C8Tim4m
fgYaQuAdCEVzHwmbtD77d8U57xuG7nWg4+I/H29FckQzwLoSV/fknx+ddpMXwynqdMg6aVOy2N0C
Q2WUlTOzEMIRWUGSQxufWs+knXuqZN2NcVmP9xd4viI3Y+I9wfGxXf41gl41zwTBZHn4BG8jlSXb
/OtjCuFfF6SC9fXfk3qGrVeF4HZ/23Kue+ekpkPqLQBzDiMIHLmcwh2dJ/+x0pjL6vzONNfh9z2w
g4Mi8rUQlbbOFtjLp68AiGwyySV8FCJT9QxU9RuIARgWC+eaR2P9JdgFUFuA1Ph5la934SIEjHdn
4LT6FkhqbASb3m6jXyAgLPjDbEU8nbZM9b7GG60QuLps1waz/4Ih7B7PpTjCce92PE4Ja9zXsHpi
uKhA6yJM/UGEuHIvhAZ01IYgSDPUKdO7x7vHVYvVEUdnJNPWQ7LkT+9Jc7y5MiSGby2REiOwful5
65NLTy836E+YlTXj4+wd81IBiaM5ZReE102A/WZg8Frem0bEJ939N++z952NECtslJ3UNRf8FeaC
f1wMT6URYuCH9AUqbz26lxzBI8qYY4yAMWoFpcduglbV1Cf9+Mkph+T28qjTO6oEb6yqQR3rFwTE
+kKCpnTc35ffPbE8P5kkgH6d+GBHJljCk2V4vNd5AQZK0QmqFG0BbbDpzjn1JG+Bn5eyZIWBkXSJ
KoZnY5CMBrTztyPH2+leyCMlJZ7UHMd+G8IPynPvtr8o2wlZ0pDoGA/iazaAOZ7/erA5QmFJseZC
EKeXc85KYhREDS7C9Fj6tjSkNH3H8/iQ9uugiaULukjvgdC9tpyE8NJTE6XyQwT62Yot4+740CO7
eVtWj0GkjUHwNHxx84q3exLaiMlRKHKZPtBFgrPSz8E2TibdMX3d8gr8OJbMCGhmyKDmGawulWsI
aK0O0wUK3NTMS9piwuOsptJmRP1Xr3VIYWT74ARLvmEQ0m1GWQ+CJ9qZ7GT+W6nArM7BBfvZh3oi
n3utxf9BeAUBSQMZGIy/JcFmbTDvMzzWHGt239lWy9VRDX8LTcFAHK2PELWO65rktH1Bmyp80Lmu
XoNZH009nJ9g2ssZ/K2GagFTVII/JueKqilvdueEtl8MBh0osKiSqs3v4JBUHLHHd6Rtx7L6koU+
LEKBoA7xv+H/zSCxCnCaKCeKiRG68QJTh52aApgn8Zzr6HDfVXVu5t1QFC2A7KyR82ANuZUQLVHp
yfzsDu4a9zH7aThjk+Npb8itDnf8QmeYG6ujWsa27eug/qKO7ev7a2sn9/Ha0adZ1oy1faf37oNI
xYWG+QE3FKT3K5HUGePzKPyPMlnsCkQz7F7QbX9AerrPfhEiNTuvgWqT7YHchDR6AuDlS5ziEBXl
WIBaGDLtmH46UQoksSEOJFXHRZ3TCO/kz7uxNFk0hbwzFr+Q0DcfSwY4xusC4ZZ+yHq+1Aae0p3Z
oCx+AKGxHOIhM+VwwJAq0s6CE2uf5FbyWTj8L/UKdH0QKJfuskRuJT7XuzBIIvwcYBAUMdMRYI8L
Kd5d70XFH9ffPlWdxKoevDMqxiDT+n+OJsAE7sh8XRvG1+j02vTkJtjT5ZySu0f3ZHEktYpUcxFi
pom0Fi3wsX9l6iazrV4XvzbC56xzBa+BOIO94JAC1d8hUJamfroSTulhJjHVRr2vKbR8M9Uks8G2
YIAoGiqr3mqV/uuRKkPLUi+V/YM94MP7rWhVQaM/0DL3bDXd1tO7BJkLfsOxvnjXiV/OvlGvn+lP
0Ig0Iu+6Ihs6NJKbWqKlkE8serGF6fa0nwu/j1H4l8FTUIcvKyZNZEjYPN1b1jFo+QevBCzbC5sJ
T2StdFPU/DyU2iGmBUPthue1lV9G+mZyGvk4NdyL/3a5wx3Ju4O9Ro+ZAsHSEpN0P6hk8+xpLJJC
OnnRVYi+H2QJzt9rCPrm7K1LylOOqYtwM+t1d6RvAm89DaHGY9UL76MRPM1T8+BdZy4LVAk+x7s7
YsKUuHp9Ag9cPqAmJ/cxJHnYc3d15CJlMV8wDzBMY6Keb+fdtuXuOV4lqwl5cA6eHU2g3LLBXVZ8
SdbfaRMQxNQbTKq3d6bK8CX7mHvaTpOzDVJgZ+Ihd8UJzHtPkiHpAp/IBHgZJg29V0T5V/J1zEcc
Z89itbR0RBWP+2/Pal6brIyYY2tYnnMjUXdSiLZYNVsPxRSwvMnBXcFQ+ua0OcvGkTEL7eKPZ+8Q
+Q8uhCF2sm81BAns02/rAp4/WTszOTCDdFVyteanEy5Y5R/z5KxCk7ytin6cNm3s6pPWmIUxR5eo
ysmb2scc0NZ/AaJEKfIUr6RbjY4HY5wQE0fL1uP+0nGVxtBczQBz4I6j/ZcRUF7DRSJewzL404Eu
OpqoMBNHmCH/Qw1vyTe41gDGFCPVw8VIqR+NvSwu6XHtkPqTARUsotEgVnqa8eWi2kPRrxV99Fao
hz71U4YLrEc/2LNLjVWbiD3X8F2IBwj6FJL88aSZ/Vkepf1mLM7Jeax/qQGcr8pCaKRu7LaSU53k
1xQuTzYN5XjqeJs5T3D97Bb1tnAUebXhvjZIhCXSeFT1npNtbWbNc2K3cgWVwHYIX2tyXHIVemJH
GBEau5+GTkTlfdpK2Syw+8u91QiOYfp6C8msIe058QgPrdMCU81DFiRn8ZjqofOoZAKA4+8oZ1CU
Szk0x9qr+AyH36cfaVWLN8g01DCHeQLb7uHcfTlweqgkBX8mtURicZHAee+Ajhf6lsIckE2Nfz8z
ZVV8rVBUvTD550eQj9g9lOUN3Lz4YseB319qDx9qrEb7HtRDalR2IXrlcYdabZw3vUvOTy3Y8oMN
CghltQK/aggEHwzIADv87q09K/KVyIJbFM8MPH7lf3pLeynneLpf1qliPZYjJ4oEDOKOuNBcas+J
79bV5brHhOUKqjkl2Rn+O3vzouaKRHmjCXqeGbZDR+mPx5xiQVfyP7DYXRfxpqjcv30bk0gLPUrE
k4BZvNTdsMjLVXBfMame0JSL+nObEEJ7XzJ9uNcnY6PhwGigo7DF06YWg7rM0Fy/rBGMQYZRnLzP
49AHYsbtPKZw3XxOrYDd9dK6jj1ojSjMHx9CDeky/zJjPJwKkj5w4b+gQfwhLBLF+wnsnh9E64rU
GDuBKDhvGpzbmPls+jVhf/hW2A6e94xALduS2agW6j9TnmddZefYv1eOXFgi00OHwT20JHm+P/eD
wvHrehb8ib/+6vNWwDwWqoW6Q8Qwe7++m/lp6gn3I03B43ZSpsUtAbtaTxNJME6JwNuHm+MtCAL/
mEhqNpCa5m9Aya2Vwpf+7YEtDy2GfBcMp8Rp+ePhpReKXSNVzlWC+9R7HmXIck+IA+cHrKxkDoyF
ZaGrFm4yG7dsvLOMpucIUs3J5cWQh1KHVs+/SIqMXiX8N/+5tUfF/GN8VoKS4Z+/rHosSNu+QDOf
SfG5UAezbdv0b4F4JxiHpixQwWRSJV4apmWgryWZ7mtn6DSrRYA3yN6JpOdhn6cligBDKquV2Vyv
B5b35KvtszReQaGDKSuslrxvV50bW24nu0NekiRCBrsTFeXi5GGRrwejhpJSEuNqgNKrMXIeibz6
g3EOZaZ3ipKZ+ln+UVq+jQlDKlVhv1LFNowYVraEHOL41tgYD448HmEApbDPYquhm7g/i5JU/8h0
MJDS02unCAUTL9R5FjehI51DGnd0ArVElfJ3CDevFDhlqJHpWmZoKXL/qzPtRQI1vxJZMt315DPK
2sJiqjhOFTRlLJq3i7MumgPzFJgA7OM8REoaoop6T8DxjtZAeSy45BDtH3BfGIJ3Ct4ecYa5dVQO
MphPGHD2+udAOSwvYSWPP9IrVAPDkkD+AalaO7eRBana8u/AxHyyLgNASquqLpiYt96a6SSc0s3T
MQfxccHhWPqCkCv5kwqrFSlfQNptedjDlsPVN7LkUtbRmRzjwu/Ky+UVK7ZARJf/E/buAIwcVt3g
IuXDWCo6lZwZI6DmbQNW5v+Cyw7b/+osRs04NFwbIFFU3mTawFolnupEEtWodD/pcs3bQqvVVHLA
0gTj41nINOmAAV2E7aSj8Fj+RLPrBFdnShjpn8lF4ZWLconvqidlIyeTv8RX8lWl7ez0QYNA49IN
CpYLZNXCWeZqmy1iC50vFtV0Q8YHltAYWcQ8QY1Jz+iSPiHNQIeyLVMVoinRbE7je+a6NalzPWCb
lQztP14vKRNzXluhtYbmj4TidcTaEIFuQ1rYdoEdxuKI8s/25tXQfdlWiEdhCDnnSK2Rc/gddcTN
nWRZjJ2bUYHJzDCzkRcTTc3SW49gRPRdCuNUuAeoYA8QCCoCMbunFqRzIr6LJg+k6nMGe6fTae57
hdZWVcvNdYpbg6INq2mNtpj3gIcmSoVghRXuoaYRTxyaBSLjngvTtMh8brhZnPQIhjtEWya9vczs
sPGw6l//RiYb3h1lxyzGKB3ElxB42Enb3T0hnFBXX+W1QKrHhyD9N44aTVHT4xZCZT1M56WtFDdP
ZJ4brlr9Q9jNS5TyuXYUwvu1drUZR1t4xiysYufPsqIu4+oiQ2aKGrwGuswqjt4s9fohpqKRmvUL
0NuqSV8ES3WUrryYVENY+slZS73Y+zpySJOQ2cEZuRKC+gKp+ZwwrNEQvt1IVRuCGPJrIvArVZ6l
c6wW9OLyN+yZ7MGl9Uvnu3bK1p/eou55hD3wh0xSI47QLV6DkbXVbmYgTmCjuGrtpNcKVHEwKlmG
P/FCAesz1hnM7SkBOgaejFzsWgY3KWtcLA2dEp9oERcGvRicZej6Vp12HtRnfwC+1wZo/J8pwrdN
ikNwjipC+TGXJN+69YmaqhdI44PFfHGiZoMnRwZhK1YY7D+xDx0SDXOkv+vv0SnVHgUNoLoWYt1+
XQwgOzoUE63aJxvmPkvBc7/Q5vnp6c7u/Gxb6C1AyDKxzfAf72Oq7/wG9kdZFnjHTR8rejZQtP7v
KZF3JKkCirnIwl3YJuAH61RTs8tslWapwK5OoLiriulmwbJdJ0JXJtTMXQA54LjIbcXIZnyE20AK
Vy4r56sI92dJr7qmQ11Kd010S/qVXFT28Wbv1PONoXUB3UfMyFf9F/z0COxMKVn1GuQUlNqatczW
dUcYyZ8YQtfCgBphXkHnFc2dUJGhDXnlBtImEjvAtgSfvh7RyAQsKTyuVdNnRtNtxC4ycUdVbZVE
6ttTdVt5AgV8oiFOUW8lc1hqpBepTH+B/Fi4JY2Y4mCYE9ph5CR5zzmT5YjNPofEfv3hjAtkLsBA
TCivClTRWE9fyt3mjICeOiYklv+UAvu9/Qg4DHqNlWJewlZfAVSZtMKoP10Aov7BdkzicviK7Y1E
F7qxoHfTuGEWvRwPjhhSsMTk/rQQK8FczaZTeryzFjnd5QYckeHVyL/nRgx6MdSckLoofiYMchpJ
HQzlW8sOXgBgpbCUKhxpds6TkUa2h8+i6stAtx+nASX1QpZhU7j41FLjyhU/ZZYe0NH9990M4LOp
30MJ2k7Mf7bgt2qSkb8uuqZtWVQ3xNSLpUlAoM0JfiPaf8GTJVRgCQB8PGSSzY9rEx9jAPuxexCB
L8k6OgDOJIHW/WHZZY6ZZgqicqNlLMP8htM0Ls7ZTGXgWI4LN347BmbpVDtSOy9LQRKz/3Ijq78B
d8xtCeCexb2MzqCNaZLcz0WtEcqpMFFoXi9YMgBCJNIEbmufGXqj8vW6DVntIbGu02aWODbJhhfN
oFIKcDDBIAgm2/JiUhwP5h67girYAP6So2o+rp8NxQJvCpaIfEHcQnoUAkJ3Q33d8+jadAaYLa63
F+a6AJ4mJT0N+QpoVrdoeK8Q6xe+qtEYb/LBNWb3dL0ccf2sluwiNKD6qZl+sl6WSi+WNTaueGcE
OLye/GiDHWXe3zo69ZoYxwYizNNN0h/nM3OVrHsoOJS4mMKl434IjNBs2jiW66TQAW+Gzmye4Lya
rGFVgt3ttP5skaVLGkkSGABdthf/J/XcPbRrlBzYmvB+t7ogkO13NcqOxnXdy9ra39JEbiUwOw6M
iewVUABXOvMNYa6+/f6Nm5446GnsQ9rLUellGLU0s6PfJbacjGY9ZSqK7yvPuV3jdaFUALdwLBgn
HcJg4TBDxh8bytwEkc54d5HkcO7zRlcsvHzkwSIcR85VgDCEVn0km4YfF9A5sZWSJYx05DGwn9WH
fosS/m9hslrkkwtgyPPYaNpM7E/ZwHnQBh+DG2yDp1VaJI0WCL8R88n/aheLeoqRXxV771NXPlj4
W3BClanjnAJnrZ0F8InI+C+o8UYnGlvzGb6WgPqCzbLG1BVbE/8O0ORiMcGdF0fMSZat4oPvTqih
T3TSx0+SDD1YXS2zSMl4XshuEdE2f51CEyrDh9yFvlDruFuLnh5iBUaxEJCG7igtItorqkiwerM4
fhB7uE+CwwmtTQ3atX+xXtJNG9TffGkbkLjtcsxbG2fQGtK94Qfl+CBraHehh184h4HgVN1PFZPy
RA9OO3pFdj5Wtdyczqi6GFS+gcUnX/khoLd6ep9ilMs7Uj9haER29MtA9oYTP7DmAvcNlIC1B834
8IwXc7aTbAFB2vMt1NLKDy8CZGlbSWUYuJfUY7B9F+0sw+bqG7dwBSg8QyQueqmccWTpyE+pQuaA
dw+g7nSb72qt8e+40H3lW0IbHfZzXQ4KFTrX4dkioJJj+XK/D/OOIa8FpEyaSBcL/sYH8IZQy6Jw
2BbEkmEDg69QVvMKAJXc0jotXyMr0ruMg4gsUKr4Oc9dNvWo/kG1bD1AVdndS+IWw+o3gNfpzG+9
jvOBCJ8G86hX1mscv7G6gx8AAKvwwuLj/5EVl95UwBDxS3RriqSXta+6UsYc+7xr6MjPyj3+/FNj
tvhhu5JZ6/w1ELH03JN7WP7i7asd/BB05sTj1OKrWKcqMrc454gIQfQN+vKf31JnwbwKG6n2MWVo
P+aiUGezvzZvbMoyRguaaj57kMy8IaY6iLAh2YD6nqsFrIyH3Cm9Og6l6ZNUTuX5HSxW9TMzpRCe
bHBZm8OdUP9y6t07gMbrb19o/5uo5S2o+uaObRQEfwniOz5Y601R1MgIa0upOnParapQVCQea1dR
HP48d1wI80zfMz5pzO54tuscPBnPGtO1Vg79gaNx1N57oj6Fc74Q6RNXwlHQLDx+EmqYoH/mC158
sW0psqELY6q9iSo31pHzWDZwhm7fCLq1S/1vtPTYTpaEIYJ/1GM1d+SRePr4O0/E/YPNhVL9v3fA
nZvubx1EPp5lE8GnBHvZxu42lHyEBCqlX3UmPO0Iylq5hzNS2FFdxb059bQ2fQH+p9QiqJwL1HH9
9ew4Y4o95aOYSlcRVLrANt528VvIJ8IyQ5wr7ErGT9gP4SIHQRwdHZjkUJcs9wJei+7Kkeu7Olu7
+IoHfI7MJQ9yDjPa8iUs+rDzYzqKf2sNJkrNLNvfou1DWYzmnj9jR7schDP0ZG9eqaz7rBcP1MSa
9sKphy/xgsqmFBvvAmdtMoKNQ1/8qwLlCBzZCxkp87p/R5TlxVW6Msy37a2GefdMlYYciQjMDmfT
STwbiDzAht/qkrUkO12lu7l8fZvbWaVYXQ1H39BOD/xJYZcOFP/YGGtz9uZkNrBlCDjfAoWzrKFp
tbrwzLlg6kXU2wgqEEpzU/9irZ7oqv0nChBUXXk10+qQ8NGu32A08ox623t2H+3LLqctTAhrE6lL
h+Dny5doSL8mDZGpP5TuXG7NyX7kFUhQcJTZB3p9AqVfdl9t9Z4pRW3ZSJVi52GEzkDtAkWN9k6N
rc0tVBmqXwoGxyWYxCCfD6cdfx+Z/QS8c3w6ravnfPUH1twrOa7UlJS74Uo4shb7O5KYOzLDFsZx
7H1jleTlNXwOJZQc3ld95Aj/ynkflq8IEkLMXGfBAg6XRBJ6y9Vwbtnof7g4vsJRk9n53u8PyAiS
deRnyicWD2kNsUrfoDXU5fvesWkYkbfgm+TunsY0xVxyD7fTZ0gkUqhuZAUcG70jB0SJHCOo1tU8
Qxt0fL2CAsLDKavbfthZvZ4AmyyPMLzqTZbrSpBT5A3+SaGZYAj/IEPWQ57VToUINY5sL2LUvsBu
3F7pj7i8mB6cJMl5M+M4drchUEMCea85fWoRXUajl20NAo1QQwYTjvABk2a4mwjXc5RIzqiXOq6Z
yCIUZRsOfRjjUkdlp9J2mOWoJJdhe3djy/P8PL04lK2Z3t7Nnvo9oonVe/vifPivmVUCFVbeF0Bw
0ARsNTHQXBF/7/yiGSHrZdy8gl2lU7umIMUUhAbVs0PWElr0Kaqn2MhPyOMrRWiEy07V3cQak7SI
Y1h2vILJx9B70Io70Mea9IfQ3GZ78hBadgGAAvDol8/yy63IZgAYv7QQsYv66FoTF/i/fBkTOyJL
UnVxwFVbT0ttB08U4D5xF3OKoB/9UJw+MRhf70ei5DBpD+7l3YMCpHA1jazqkjOin5rExvDVTxv0
pDSp+Jtc8oGNGL1lDkIN0UFajeRE1P0wUoD05XTaUdCC9cerM6g3A1WvwpHJxz8QY2Kcda53QW1J
ha24LWQZ8oJO6t9FV/vWaWM3nU6ocz/Ms7aE2isu6RxuknUFfu91qSb0v5ZesoQQomvIUjgcmKGl
t5PFTx32T1BAot4js6PPuJf2J3w7xYt7APgs6rbR7hcVpat2CC05vt2f42P0RZfJgiCgXsaMzPU1
/3IHqDnOvIra8kkKQ2MrPDSVrAyopq/Hv2LasJcsP1a5GEljEzyuyLkMMxNBxRezVmPIe5rDnI1J
zfcA8oaEKa0pXM8dRyn2sTsXNldrxuOlLYZl8SIsHBzS/HAXHUrvdb8RkXZ5mSMnUVPe4HaDftXn
uCVkC8i2qCsf0N5TFnQhKNnKzEyJvSny1q2Pm2rFkzfxZmUYX0qlVMYlXMop1mV69OV/LaGO44gr
frzZPyRMJ3ohlXY3kOcGj687ISiHcmuz9SNYOHWSW3DgOenbPz1TIs9wxs5XKk3hUZGs20gN4Tpb
GOkSusbxBkreG30U1/ZYIWspca/6thwut/dDAUvJS3+HF0akki83IGt7LOzWd6pvU0wsoZjQMO6k
snOqvEbr4gIA+O29Lm0NjS3p4+6P5lFy0BTEV66z0VslHg1SYpekLjWmyjRGUgBZXoT3gqhBJDAr
11SxR4GEhq2D+nTzde105SS+eAd/xJtrIgh0UP2QsXTV1sZcB+agfCk3Pn+iqBZ+f93xVMvYTSez
01I0reqjDgjcFQ/3SEoVPz7xHSZgJAepyuIdAChNz0WMqkyXLZFA5n9Q5Cx1QKOjAqiASIs5ZDmE
q8pYfIkSpZ2GV2aSwaXqPZ9QMF0J4QtEYG8U+W6w9t9Cu6PU3slIBueCjMM5EgGORD5+/9y5/oQG
pPSbhkJ9oABQ/RD8524RHnTM2Aukr+vR39y1uJaJcsUjwI7/eUnxOl2L4Z1ENFOw41rd1dLl4Sde
dyHIsP8YBy8k3ZhJ/HPuC/XqmBpgO4o9NcFiYDMBQTfvgJaLYz9WJoq2nbdVTYIeRdxl09N3iSQ9
juB7GGQt+c+xFpah/rg/ZvCI11hpbss/EFgiXKwn4ZqdM3tbNE0HnhEFJfUAj3R8lsxRKEjaUGzA
6Oe/SoiDxscKiOwZtSP3vuXJMwjpHyuSHb1TKMgA89UL+IStblGAt3CsWu9dmpcgknBy/4FirhgC
ARi7zpfEa8R4025PjUeh0oZEvfR4ufBrmfOXCeL0TYKP6flCzelRjQmPTS1urjCtXJr3P9b+Xilz
AfDphiNFoCWXmI0VUrE1N+/FvRJW1QzPumcM7vDmf+iYJeyRb2QbwEqHGuBOjkPkNLJ5K40JDbgF
BwvN7WRp/x2X/uYl3BOrC2pVQuuJobqxZaJOKdOerSOxHlrzimwEJ8G3vjrbvd4lQ5l7+ayj9qDS
tUGxwLyDkeYyJh03uVIO8afq/YMex/izxeWOmNZJJVrtZj+eB/ZEP7uAGhCcBYK3YEQmnDzW7aRH
Xx3k8KgMgjA5KDvfYXPtQmjuZwO6D9K/QMxUJiV7DktHiARzyq5mg5KXN3zlNTKQdfyxtK4mOWLR
l0h2kGbGx1lQqX/ijOQIwOmRSnzP8J/dcToMvqkUIuW2pNddUXrFfZrussUMoq3cjU1lc0BdHRkH
Kp+RI9sjN4yUL6fbkLlM0qHDTJcfu//T/i8QPJ6MXTIFzg1VFXtA8we4VHrSLAIKs2Ewb6cHxKZm
z7nU51vVS5quRnmJX54vAA6dYCVmgkmYFoXxlXu4Yk9RyLl+an0mpjTgwb7x0sOL/2YmPf1Fwkhx
Sk7n/w8Tlp842UanjgoJSWxi6SmfN64CbBYJyCtal6B7YiU2xUe6QuIiYy/FIWZYTC3fx4IObT5Q
BLPae+UechtYhs/2qPM3b59iYFc+ODjPrm17J3Iv+yS3mNijAYtiw3y+/WULc8YC23m+5h+1pfXn
sKmSzL+Hts8+0DEh8rXcTQ8SojdMsJRseseOPpAtBUp7K+Gc4pmiKOrO4m5WI4xgPJhb/dgNZ9ry
VtKk8zbi9bk2HqQx2P3zEnw9ccTq62XTXq2rktiqb67APO1I1huruz1Y75lQ8y3XuGE9bjwyv8GZ
wCSFsfAftD5rNPozRk0O9+nrZ5vsqFa2SY+OdA0fuv02TFT+QJEiOchiDEch2nSjiZMzZa3dpIc4
n4qEYKFEkgfzdLUcwgYlG/1lxsHUmpCpmfyHZ6VZzmiGxWIxvk68cHmmUUw7poxKk50e0AnSBZG0
IWRHzdVDXhzgGv5fGNTZl7avb8wmL2aZtD62NHPo90/pxK7rHziFMBrc7lEiczP9WsGccYNQ8uBy
DEppIr4gOrAHXGxxG+IJhkHwjghCzqe8/yUoAzJMOUoUs79jokPDj/3Gt+dkGqO0ynvQ/KlH3648
QJdqDOVV5uL04YEaisU4G6+xAmI/4qZ8MQr17jhjhtJea8EcsgJUEsZhAf6TRF7sKGVVfpcUGzU6
8ruJROH5exSwcuZ3EKXRbV9OAGI1GcxzTV/he7v6We14ooUH4dxveJlzuIW2qFBZhrP5TcDoxC5U
1y+zpEGxC/CvPGdR5IaW5SheG6w6TjgPcdvBS8A344peRNSeNH7MBceuIhdN/azeLm+NXaUBIpcr
VKPi4qpNuO2c/LFXQpeyFC/5j/Af4ScGeUqkvUZnzCCRbIOjtDcntepC80wLgiaCJoR//84Fz8ZP
kwfvrD0rDYhlHQsSCXBH5oxPCFFz/qAwsiflob5VSuN3Ly3Wk3fNafn+nRP6jQhA5cFom66Yf89t
J5PbK56HZJWDx5ptnJCfozBW835t7zyZn2WuanqwNjcPb3t0Z/2w+pNrbMgDR1X3+P9lagQDKlAz
UmfzV5rV7+lYza5DBbr0KOvKFMM1HdC81RdaUTw/G4fazjk1DQWJEon5Zr56yBcjBvkdOspovmMp
80TUSd1HGFG7y513YXNl74feYEPlh7c4i6NUtY6JfA2PDfU1to3+lsFeNUpHh2mXjPvSZZ775wnp
y4bI72KWfOUq746tZs4Gs2K9cJ898CfQwXniEYs/TFy6yFEckCKfwQXrdiThlk8HFTYZca2/BZxf
ELmLpY7eNupl+G1Fn19YOrkahdqGAdN8DQXbhNysNikDCbGMZV/YR7ByPkcqkXecDwOq/cu7dZKS
sBSdeAb579KzEiZLrHMmz294T7rD+UlhjAEDDnIIC9LdsKhXcuQO3DrWnhpCaDCOxd227/b0yhLb
9m5lg0QNmW/478eo1z4qDTWPTGmxzdxqZZxSKnKAgy8iybiCETDI/n0+mFkzaCKDIwn8Kf2d2+sv
JesZD5Xae/5L81rIB6XQ15cO5YtWoaU2kqxiMIXxstHxMq0INEqqkchyVso8IQ4TU9OE4+94rQNP
uj2xfNkL5alCtjPUVzxjMY5rulOTbLdMVMOc0rGSuXvRV2qIPBdq/fiYiS8PJ2lT3FxUMAwsuduC
Rr3DY119ADOooaAWOiPXi8CA5Qf/ZfcRPx+E1JWkZGjcGHnzzIVW99HVaEOg4yxgaozYgabkZtR9
e+MsgrsSxvX2OkHq7m6tXe2IZLtbHfntT6rwMuP1j8ZARkqfDO+IqwfDK6CN7FSxKpp/0cFGe7/I
NNjjSSSY9CoIbFg9y6AVb6Ks1quxT7JbcJTzJwvM4bR1Qi5wsknbSTXO+Sh9vFte0UPS4UVOLUTK
ybhmNO4GMeNqQUGMGBcQCHkPTBhWfJP33SaKxIPT2hRoYo/U4n1pPmJc5gNx4hvhpOPjao9JKUUo
32MmZDRzEvpdIwbCK9wy+I2bSClsFXEGvR0b1XZBBhcs9nGNYpQVGZLNIsR+y0Simmf9rOoOSo2b
1vbkmK5oURsBGcugeM3ljOavFITFNsFq81OJUZWLaCY+l3xAuAUJzsZhYE/+3n9uuP9flrKfQB5p
rB8homoJ80woMyHRO9zX8H7PVTzzAiZlpvWtbzRt2+nMIR8C0mKsutg9Jl9pPwkaHFzQx9Styxcy
xWjMI4w5nyd7b/3OHYWaCfoZ2URkfPJPpeoU19+D6ECbYeD9SZRP9vSPWSJfuecOYY0za/LZUoxM
HNmxw5u/s2fkyd8jMuIK6yUmBLqE1QzzxC78HhzNvSn4hLUpKfshJ0OkETiqYr8gVNVK+M7Ipw0u
As/Tq9PE79hBIcrJ9DxrSv2+uY83to21Gd3UYHMMKQ0ifhxcPi0XvPLOmJIGEM6AVUO2wuBLAXj+
OmqYckpNOSscv/jvl3YLlvJ4OpixvnUO6wIR2VTGmxFGIXfmTte7/TG3khL6L3qM33gxMJK6e/ha
s/nnUU4vnhNKNkDkZOP4nS73Gy5MiTu0iRLTc3ufWxM7xJnr1dp0zFYDQRQaHWG93Fju3DfD7Jln
Pa59wHZ7/wCX/3e6HIlC6JzHiSmOBr9bX1Bnvf5ODrmmxsmyDiAIADKECcn5uNthSqDVBTiDFkrk
PAK5yt3F6XIddmJ0u2cbH/ATHKpGFeYs7YCUogj5JywbubwqrpCoUb4AHQQd/iJXPUMyk+TZbQu+
8b6UEyipR5U4sMW35kKMCcw/s7S3ngi+V/Vk6BHBXSa/bTX3UJ2whjtqAIojOzOZlEBrS7DwFp3k
75nzuRr0mTxXfMNe2GOr4WZDT/TL/rRkKIbQ3Qom4u82Zvflud1wGlNZ9m8g5opFRO/vJznOcJa3
qREPJsZN/Bgwg07J5jV95XbNm431jjONevOJXSVuhYcI8Xvr7G1H2RDDacvkLctoebPCH5U9h1ZY
IMiKZz+7o23z5rA8GWWrkLq3QVW8ttBFxUT3DZcBi0m0lsnjnE148JOZgqwcGzfJMJLEIC04ucaQ
RHwn6kz82sb4zWSzo/ekbrRShtxhuGpH9CiYKRDrSFGD3hp7JHBfuqe8L/OKsIUMGFr0Bz53bkC+
zctNeyZX6uaLu77Jo+h3lOTVePqY+tvBL4taEzLYJyE8xybAf7ZBcK8HZQwHndg6kAbHC32UOWm1
NDHldqY+YAFAL/khztCe1mopA8r3Z5XCUe3aIiGFrsg2RZshC4JIf/76LLgmWozynmUUdi+FmmQJ
izASib+/el4alWAjqSGhvzT+rYJme25avSAuQVrvKQkq1q+cp4tLFUWNALMDuHSKxLN4QGf+TMXF
pGoggXULw/msv0cYu8oyWbq4ZG+Z4zEScckNOtwCQQiVjiTToIZdzMgX41tVDH9c0XwVQiygYJHy
tuDeg8M+mY3YeNUNBuRumEGO2Mw+VEgP0sTjcgTT/wE9q3cVn8VLwBWS/kztbj9ZM1bshkmXT0f2
VrvsxvWIZNsGRtzLkWzNCf6RMTTTN07Cf8lNiQBsT7ESQIiksZEYEX9oDkS9GUM3FGA4tUvPZlpL
nVjfIpkZ82ZSWGr9ivAJcjp1+PdhOw8if1r48Nu8ZBM1GXqTp0N1wVUlUJCY0YPDj+cxX1B7xK0g
L4ITz4N7FRNGrFHm6NtmqPxP0vU5ht6a9WnVCX3Y1DBiqX5F/5OYHtQxQr3SD+jzmCmZN5F93qTC
oW3dZS8sKrk+pac0DUAW+0p2Yd9/GfQmuRZElkBQizRBvQeUqo/22Jaq9fvOa7y+0Kefudev7621
dEqWwkW/pY5H9jJ16rzhlhCCJY9oIKR0rAhpUQjrShrh2gKsSfb2qZGH1SE00Oj0nYNGgKVx+9EB
30JKLMJpyaryjACBBPwZtoYTpqD9ctkj7FUpShwrWNBWkVu7pyhnYVw0ZjWR5eoj5+0FnApFV7Mx
qOWEwWei+FaA/BTEZYl70KRbZNQ2XzKkHcItVXml96qojlfFjSg0vOi2RxOSxKVKC6tuMQIjHMnp
jPTZ3N2bVcN1beElytOOEV3RzO74Ouo7qclizDXrxuhM8q6pHKCP/jZ4gfdgDiW6KDtTfyQ0stDB
cBi+wKewRGfF/7VqrAy3ZNpPa8xuSwD0s2pLThkJ6N4ArS0hlRMKkTKwT4c06S1+0/fpnLyAPBbb
pDQS1tqrZrKWEe8mS9A++ucQg6lBdzKYy9lTqO/sPNEBHssZNLKkD0q0YiRsGLIKUf2cgWccCo8I
Gv17XvXcNA7jhW4ELqvkiZGbp23Bp4IMkvqNRcAcUjjf8Vc+aPy7NSEzS4BxU9Cfye2gZj7XkW7o
p2QnoCvGq/ktN2NNon+MY1RuHo/+p45RxjoDQB2voSmWj7JleH9s2AKhgOpfTqMHKXjBt0sWqOx6
2+KKUVO8ismvPVDx4UYkcjOriMH8fb033zCTUDFwALAz2xOFhHTY33SQHSWWjq7G3LWmm+MpSzFx
KD+2+5IpNYNA52T3rrz58d4yQHPFcxkIqKVUxxVpEPbePehm0uveOxNe+zuzBG3YrY52/lUfY0gD
jO8sv8nhLzUQHzEWj0aqWJrkZ6b92NCeO2oaJxlFMmWeyMm0Pgf9mJHecdg+cRs6RSgCC0NujXR6
7CJyX1VND2uOAqi7yQuWhhC70ELl4oCWKlsczhZULG4tOytZRsTRzxihoHWaGgvBcPI6ixNGuHcX
mW9fXZ6bphAGPr4oSk2smvdGAekyeuqkGqdZBPMLAdf5cbs/8JltMZL2XOWPaXeal9SDjTecJBky
tYgtt8zczGM71ZDVMr5lutO1EbTfr+zqBA1PDGgWvjm8uBIfvZVRoT+0O2oCGRsm1tt+HNXPRnBx
frGi0AuyxP+gsk7KajD7Nhgv+L/W+CR7UagWUZZSPUwthTWMp2o9vBzenJHanjGi3F4yEZm9C3oT
z+p87D16aRfMK49Fq7od20XP9YM9yGY26q7lfBtaRA82lAOo00opAJcSnvwLkUtQLY1XNY+u9Ber
fRWbP04SgqmWnPz372hwkKkFFGnulNd5dCmCJyl49VEXKEmt1FTuPSWsEG6w14mASDF1D9aVhSSp
8VUTkb9kaxb0vUKLdBESfVCXYpZSK2wFkwD15PedCzJsCzVHywlhBo+U/y0HTwX1tkg1XboNaUSZ
lNr3dzJUUIqOUBw36NGi6St/0ioQZKBHRqgaUEVH2J5joJam5fO8OkQK5luZUw/eziUb+tKgNF2U
jYJS5ZVKOyLOvo6bD3JV95wuzweQ9XITaqWV/65V6wbZQ6+6l+HmD9dAenFSDZDOuIBKUTknpOaq
HVRo2GXHIFlRm2MIskvRvgEMFwb6/yysiA8EpiIBs1j9l3KOsELQUlBjtCHQ9BwRaboRYhdepeIf
lnaraPT6LYX94kL30XMm4biAwcwhhS/O8F1YmGbZAjQUQqJoScrBhvQ6kGvl5k36+ugZHjJlOGHz
oVtpudodq5w3eBAvXB3LDcq4Jzoftx+s5Oh78RldVAE+jGT7OBIj5mSJ9wQQi/GJSnSRiz739QpK
mzZGi8yKycuVS42iGUrk/pNrXr6PWMwH1ISFxQ7mBq4TnpL68ttq+DMRn2S3bV3Evqdup3ult0Jj
GSbl5T8ybWVUnuCYMjMUMF6+8nQHm3GqqRGcuWqbPp4EljfoSPB7Nkk6AKAnuYlY44Q/sA3ai6YX
ajj3ex+LZIE5VkNA98bmdRd6GzZtyubNLATeXN8ppSiz+kuAVCtLFlauxBS+1o6woc98jihqqs56
QAf2PbPBNsQI/qJ8kkaEIrutHDos6jV/gF224Am/VNLh4m4XfQsRLfiGZkLfCFzx5odnmgmzKTDL
v1PubaywFKeLizHqvSgmZg7Bz7q2OF/TDgm7vLshQVMvPZ7uIW5JO/bE6cYsRltXiQ1C08NsL6Gc
nCMCYpAwDdOJcEcmShONkzXXTWaoLikGsJ0OU+suvdDxYWDBDkYDFIPwSXHBu+IbVzOcqzPuUcet
hfKrk0GPip3mq1ukXniZ2ZRyCXoc0KCXW4nDEtcBWcjiJc718AfStMWk9UYgC+3JWq/6t5cG7C+B
lTTHtKqr6N14acCj9WpngZyQYZw5HIufH7ckJZj/gueqf4AC/xnXnq4W3DlZPiR+Mjt51cevihVo
S26jH8waYyUZfJjBknuodZtZ7VRZVJquEDheHN5ctYU/g++zYvuaqnuYqL+bfK0xMLlA79zz2Bdb
rMmM4Xa+UgrOI4Qr4kfWAooK8trPuqVVu63JNm8BPr7SspQfQE2EH0PIKXgExUxKTujgpJBHDa1a
w8xS2N7u2QvmVw59NYnMKVbYzbLaLc29Dy0+7vSZEYh5sNVrOxEvANe0tAyaWaq+wS31+8TOXj2Q
+49SXEonMA3X3hgEJZh83YCgqhj0bwqBzxEJ2L/vCatfdLoYWAfgIG8hauq6jhqvM4ugVcEZdAU1
FB8ITGnZGk5h7eQul5xvSzL/42IUZ0NM3RrUzVYCYaEHQP4Uo8uZYI8XgQlTvzeIggCvPOzp1GPd
Hsef8LiulRqsqaLpabZzXV4qI8+f7uRu2v0zyaXzc658jOsqD1XTWS4CEu9/dRh1m06gFtIzPQqW
lCLd8MLcS9vcLVH9ViuZc+KuNw+tJ0AwebmHjI4e0kqC/gHA124XDk5T1p4vZrg7BMiYNpbHNvmb
C+FzcV1m+maLuaZsBq0vGUYy0zu/yo3QJqtTcaFIkhoUrNAmZqSY3TRJcSRS7wx3bs+DRb+ON4e8
B73Jean2D6bS6LLKWZ/T5BhLqmTU/NSLR3qPjIMRv2+mI0axJCCKAY+RLMPiJBBjp+d7d7SeUHKT
tgpJA5uPPZN3QizXpK85rvqM7PCZQVPyNqorYjK6zdrlP3R5hsP+j0kq1qwfYQWuAPNaXMRkgMe9
Lo0129TaIVbN5Diy3VU21ffhH5EQN0MYab75mGMc9J8WOztYxLt5SpFuJ+nx6Pb56SYh/SX/lPHO
cFFmaOzLDq4z5okt9+e5Jpz/cBP+VD0nosz37GZxQNMIPWTxuDJotwZlZlHSBlAgK8yVNffO1rJN
I71j4L9X7V2NhoHuKlUICMDm53keiPXC+U4u1Uvor9xTYlSwPNQozsq7/YdH5SF1MBr2acvkSXgb
aSor0SuWVDkMvYA6n4eOqPiSJylkEi0mQDgvrw8HweF5nWludcq5++fs9qIpQkK1aCv5EukdAQa/
j8v/7bfUW2mmW4HUNpdlHdxVq+77gVvgZwBRj1xt29RaLLustiZ6HHSvCcL3fl3Mqmpk5GR+/7tH
tukpNa6+1RVRc0QB3nb7vYJNBMhBvrxh2ThSylvd+N+EctrJ3Yebp465PtfMiQyljjnZcCc8Z6hD
BRDG0x8q87Qh2EZmwPPmZb2NPd9dNH6OoGECLK+VWcnI4/UYjrF9U/gxDkUIzEuD1nJni/j/9Hgs
bPDT9H9xHpeOkxTSH76TraKtuoXi1CyXT7ka75aTxPQlv35hmDsbpJl/Wh+moEkEPveb+9sIYBKa
O164/CupPzEBgJ3pQibf7lN60glQ33wp29+wnhTEFvLA5bYcexb7pxGF4HAdK5+6iILMtp1WK1kb
w651h8k8b5+AvIIQZHrF1KQpUy3DT61K8v9EOKlNUfMPnO1Ueaa8VIgqv1Z46BbnJyICURwpactp
laOwNQaqCwSSx/7qLR80iILN0kqeFnBE1YfJqavTlk3ivp/f8AU0ddKdHNnlM1fiVClg6HTY7Bpt
VUN0jnG8Z6f5T5tL2PkQT7VFOxbHxXFHSQ6V/tqMoTwrJpqED0RuUs5VgTUmiAU9VGP107/AtRp7
DM75VJyQgtCEmkOx0a5iRd9qz/fFAwi0PC30QBLrQ186dKJpT8MWZGV/SXn+xieKXuBfVhpJjvjG
ffCcEXA2pMJXFs2I0ewH2MlKfq4+2LqwS9lEP6dmU1O7wf/kFdaGg+DYOkKWpvSXO4wiIANE97G/
Jdfa71Dvw/KHsry9JB0ja6DUKyLsw0H24GbcGumGKrZUl1szk+Y7O/WxqMwWQkpd15NxqaDsZLps
9OAS3glfg7TbfouqR+DMqBV0fTHiCSx9IZTPgMLEYpV9PBJeFWIUn+lmNZzTcw/Q7hlGja1WYlxq
mLxvIqQ+jzxYLehoTd2BvcJDcd4cJy4Bm/AokMuxTp8xmBslqxdxZqJDTlKtdregc1Nc0MqAIB75
n88wChJRUB2f4rgPuZRB0Qluu+bzsb/stG4UlFWoZ92r/5Ql75SmEoSAt+CryaimDJwfesDnmnRY
wAJLLiheULPMiVb0u72AGpRFmBUyRbPWrXjZelkOdhsPrpj+UXIl9tA/91OiXwY6m31doOMKIOWH
dDljDA5imX6Opl7JQtzb/tYnEI9a7uGPyLZZgklNqA/N7VQo5SVz2BhPEkqXHs3Mn0h535x2S/iv
qpNH+FOMRXBoYrPHPH1BSGscIzV6OpJCc2qsENDZ+HcrSGZUYzrZ6lMk54DPfJAwOUoa6KXEyiQg
sbqRhPccm70/UUmt4sLCk7bdLFQjI5kGTghEoZifruXf9n5JnXuq2WiW/NvvGzBNEMlaTg1Izlh0
3Wyn4bmrCsqi6gihA93ZWirOg78CRyMBIhhzfFWaudNJhG5INI025NVW1+KbkvuRyvAJXMycQyjs
DsoVdmjNmZZczZaQxk8OR4C6GvalsZOZm78Vwv8iZqScK+Zmr8nHLRYskCDMBPkISBbvGqxUpABa
84ZKLKF+z6I4h2H2yJfl5EEkCbdaXxJqTLbdq5rjcAiORvlxLN4aMrk6WW8LQmx15k1fR0U9vpTH
W3BflVQVg0Gief+sIYVTBNbcspf7QHMI0S+bqfR0YxSuzJ8dLDcCJrWt/mwZC6LD1NW1ubR3O1Xo
Sgs3zQdC/40wYGMABA7XQHG6ra/aj7HOQ9se+PtSrSfhmetI4ikj5kp2cg8qBeOpJA2xVcHZYz8s
zaBLB0nBf/nP65TTd6jMcuIvaxisP5nFeFKfwMeMSRSzcuRxf/3EPnmdFSDNbH+dq+bz4xY98qao
nsKzXsVzDeV9p40GowWmhhGZXBfSU/nw3pD6o3bhXdgcXpowynw7dJSrPTPrORclzBXfMvyG0WF1
kl11TNmc3etKLBZpdJNdKmC6MhCuSZm7Ebd6K73o/nglQL98lasPg1FDkIC7m7XbuMsJBtnOuImg
7Y91RH2Zdgc8T+jLXNtH43lxrL0Q02lMFX9FIZvqoj48Cgw/Dun2y5QaRWGf9/u4CutQBRMscDGY
ZwV3v7Jj/n8a9PUoYApphkL5iKzCmfr4zY2QG4BzIGESg/S33EAylGDQNEq0b3do8/jQ9IDfSk9P
vbM31BFTBsTMG17OPixNvqDTdhcAezfYxBkQ3h4+LwEC27gB6TgTallVANUfgxO8GX/2EN2AFnqm
IMkLO4KABFzxreGKIfjUM6jYWs6UZkTkBTxyoo0aZVMDncuNkqysZJN2BKESSep9HCj81n/7gHJc
LADFK4l8YhKBhdLPrGLX2HmtVG2aLWYbp+7qfLgPmYhK2s49neQmYWAWIlvsVGR17XutFDJ/8fhH
hiCjJUSSaFzToWh27356UzWe0EQtxmsLCPAfS/BBf3QCP50xLjhUCotX+XHmuI/HUiRaa9/uN/m8
lmLdNfkzIFV5fxi/593oLP1APNYDiGSVAGM+YE5LEyfdLIuCSFvEvrurOPLZC2ClUe0tIIjezR2c
pCH1fasjsnKW/W4AJyIx6nUZqvKDPll2eXjOe5CK/Kw3Z7UAtiLbOo7Q28P0bn3WlecEP1WKY8rI
xm5m+WIR6cIopiXQj0pdcvlzad3/pnfQvpgtQTYhLHBNyrGFGN32visBdvnvABJ0uDbaxMG3RbTU
PXVH31OLieCUhz6IoWZOGAHzopoZTEiTgUjYgoI59IjzaZH8U9hO+KlH3jeKwRG6gjOt52dtE6ML
PCyfLF9iJjMF2GCFyxX5RrHhhBViMeBsKOUou/umdFworMAIt6eoRM0QOxc7VVLHL+llHG95eFHc
YWRNHPJPfZEzqvwgyTMKU671HC0WKB1SQRdwk2ej8vNo1cNvYI4N75p00FtvZqz3g4tIy/ptQD1r
NTbskvBC2c7zJ0KQQJ3csIEzilXeNkq39O5+3vDPU+Qe3f8/X4ixA3c7Z/mcRsPIWuaOEtbnm8M8
EljnofuYnuN3KEAH+eMki2wWUXGOgy9AENzkNwE+JnQ/dFdK+/cry2OXjncQO2/6UJEzBVby0WuM
Wtw/qBNh9OiVm/Zw28Ne0ksJRrHRQg9Jc4FMPUJ7Se1cq56ljtK9pvxiE2JjlYqwCAwExf+O+dbi
zX37KZB1G9Oap4YseAeh2oa2ocnsM+Kiz3g5faFkA22kP4bBpy8Q1/XBJ/jAlsy5VN3i5GNArydq
qGo5RVRyqelTq4VGQNWbedIpBHmYSlEiL/Cec0CtJGT6Mspvt4iXnjOwjF2UQTrFgVGjy/tPWjxd
ACzltV6FTpxiQ3X5nmlcYkYao0WqAQyYbqiNvbdwjBIKARpziBgpajd6pDyjSsijgimgKMAbX8lI
VxvU/l5ni1Lv2PDkmTYqf8Ue+Fo5NtToWmxiwX+Qzmrv2SSh6o9oTsnGn5EZXrdEBaMoFmrBpB4B
Ocd4oc2MiQvje30vlrhCTCr7k+b0m5cYUtDaQ+G8NKX7+CoQmnnvCRiB33yvjspn0VoT3UAkc0YZ
ONdNbmEqRsZOGSQcGwARXEk3X6BXIS/O7DVNXnw9uWU1gFx7DdTnIRGgc9fro4tU8m8uLEHgmoRl
yn9cF2SHm+BoNH5tWJeEsaz2VqwYwJBeOMopSC9aHdYn5GbgwlaqcSPKZYz1UR/Dpw4BlerWwRkY
hJhP8QAGuvsDKaj/LxepJbP1jVUx1cUew7sWM0BKeBxvPOd8zWu6OHO5KhHTZ1NfXNAURLxbGdu6
Wn4juJEaxUwkn/BvYvcslt3X5aCLqv5doCpnfh9jjGlFL2LU+RELZnl1avqkhzJzkaElXyzxcWkQ
ieC+E9HtwXnikVXqukDPxx2DX84c5NSB8S9g+2zQ+NRYTTlnDtnCyJ5HSpU3iKOAaA+Wcl6l2Fk7
GCYkpDP7+f5iHeaZfE70U7p0QSSk3CF6Trc5QllwX4wLUyRHbWE9SkNDOAa9QyL4yUFXZW3BneNU
FF8Brz9OKRGNcSe2tZ8JZFTOxlvk5Th3cGlES2PxGzzaOJ4tnDxVrQUvImKNHNdN2l9eXHTySK05
r8GWsiphGxy5mqcJnVNj1wL+b0B3oTtiHkTVLrmosR24zEOuVDu2ROGSHoWxsLVbVYaMOd6y8kBA
8q5Lb3mj8hbq5lmPghuLTE4hVXcBoYVrIyhhxafeTm/E7723lw3FIe8D/w9ObcxlvUlbEa75Cc4S
+k8XXYUeCsivFqQZrEqHln2haGlWY2W26tXoVlDFzmDsE+TcTiblfIPoSnmUKTBKgqpUCD1DyGlX
+m+W8iqCuKIG+3tueW3Jl5RnlOb5uRpyOqSlRRq1GrEq2JIOLiGO2UMPNN8/qyPMQX1p8oq+hHc7
56TykZWVlp5DIuBsucBoim+KLQK3/2qJNBQM70rAXFLfMruNbH0fVTexLV/x85Hk3mjWhi3A1iwx
epkrB9Of+XVmW94DL/Odz99s+OUsGXt8qjV6ojmSdd9v9YvUX2Q8z5n4QS7CEv4gPns+GXzspVe8
5Ez/Sg7YOlFV2Wf5loWeSaQih7hZTyTmoIiyji3OU74z9D48eOoN/nn1srLXm531rsOIlNB3VZzu
/o1mN3SjoSESOkFmbvQBA7XesEWDRp+ObPKkuGdG3S+tkOiY9rYiDaFjlY1eCCOM9VTdWqTWlh4V
DIPaV2I0R/c/QHuKcWzs3BQoVBTuLcIBvtNvnbySIYoE/licE2eXUIsX6KZZjc3IVNHvlU9o0WWr
u62W5/nhBnEtRHACG82pvu1mTynHK34MQ4EI+8hXqTq7SWhKIm9g2Ah99bq9n/wVPYGVKkw52J3q
nUI0lxVrVVPyC2pcvO5RuB0/xX+fNeHCRHsRHdp5UrNZZ4GzL3yh0GO17RMt1NGCKUaisog4/w4N
0GNH8Scp4QQuxR29Rc6Tu22GVMX87eqo2OuZ6kuDKluRBAqNBJundhTenE3aYX4413drgtMRCDjR
jZAyER75cwvmVhGL7t2ekn+xaWLPzjPxpOvfbujmWkxq7eVH8BHMtQBoGE/EEwcngJ5diszHedPo
QmKmAS6B5Zj9Vg+NcgF9F7VF7coCQi2qROq3eVpm194gs5dfGi0aLav6XisJIGM6FbNRDOh7k1u4
1H0xTghhyAG2wVoUgPNf9g/KTsVf/krca9PRjhQyb+E60EuXpRtOH+nqL+mfZn7hOOH+8NhnGWpN
735R03P+Wze6qnRWy72ct3b/+V7Z6vKbcZIbe4GpyRxRhKhJ5zyGXd2gMmFNr92PbqXynPOiFVGu
7hhq/NgHLRDGK4vXd6+sh8dKHf4Tn9ykEZY7DwSjpyfXHYxw1F84RAZBKaho1BTp53Jxr0Tigo8l
qj0KCAyrUjv2jD77J1oDIwBBY8vh/sNBffH+fljDzZjwLM/FpmJVeTIxR+hVXVyWOXPb5Ec8WuKE
bwSAdZlGmAHbjQErpTtCdZQTkX0OipN4Vl8AesVTAKU5FpjakOXgMkm+E5b0anIaPrE/yiWPthFb
M1G3U76iAfEC2v/H99wbPmxtvF9gbYBDX+WEaxYBYWq3e1WhHG5xFFq/WMSn8wIoQAwahcAEGBRV
haOEtOB/6q4cQOfvF4UGLEPUeGQNjnsRFmMgNg7EiAq611KqjaaGuQ0Eqr9mQpCfHzZtOfbGXoWv
2TKSZlkVjtkBiZTit2gIym7QiaXWwYxlZK7o02kQzbyOTqp+A7x/gUBNkZPCYiQIRWRfkA/J6nhI
whaHXL6m48lOMbzm/YXrVNjNqre7QWJW4HpAnjUQ9oRU6Ry+dMCLJwNx3hiBenpsI30bVpupyHnX
U+hqD2PLydk9qfdo+15ocdtb4+st9umqHmkA6WkqlTGHEKuYVhxiKBbLPcqlH9BJl3QMKF7UTNT8
aS8S1SR5XLHK93nNu0CSW0mR2yzBEy1BuFm24B+fOx1aQeRNjBDaFac897TyJKoRNIcOMc41eCEF
o53P4k1GKQG7MwzoEccsYn/LdrMGylDKqflqtWTFsAXmj0Y5IZUb4qQnUojAioJ4Qnwewp7OXXsF
31s4HpLQ9iRooWmCNI9dbYhEsWx7D7UPyADcQ3QoVDfAHG0QbWY+orZASCfeDx9M7phqiAAWaJy+
w1L4cD/cXZW05nvGl/toxBPt6mtipCTFqRYKKt4UMj/wywZNsD6gHbgE/TuVhJQSX7SCjtToUeTk
+prBOTfTpTwXK+w1EXrS/pfzH0dVtTneHd4Uz0nmqNQlG3ZQk+Ri9iD3SQ04JYWcrhi1GNUAKCrH
SqJ0S4I2lfI8Ls63sX4T8lrOQDZg79TBWbP+NVrS8yDyr3ku/SdLKf0KcCjjXcA1jlE7KOYkIT83
tp+lWjobkvQBr6yDylMdHql9pFgEqZtNGbUSdMYa3w2k8c+YUG9Y581vaN/HzjMdoHTrFwy8m1CS
mdQLWw93LVw7bDcHz1AXW/w3F9mihgYnM/0qEcBIsPh7Bk9PyaW+occvtGnJXULYGNphNY35K2pq
/8wI2JWsXH1V9R18niHZrAzXC2IjPuvMvt52PMTNMoV+jAiJJYyqjz56aHgfTZ7qG5xANF09nQSN
IG4mEX+Rgzuk3jkotoBgr96yHcpkd2Ph/pz6R/anj86jXx3SX/KVj+kvGdB/7nkf/MBboWre8c/i
Q6uT2Ol/jkPhiTPgYcM4uYqjHIoYGQHjTzxIKgVEjymKu8Te/zY773hB1lIMjUd1dqWwwFvfh7WN
m1IbKmld7DwHTgfsfl97hmZgwez2YDzEFw+4r8B2WbsZRpECBt9FhrDjBUscuPEQxL57+bC1cP7L
2HbVAKCrODyDT/FGFaUfNpAfdZHMxTDZFsKaN5J1QNQE9deJJWAnDjOsa8z+YHmMAuV8y9tdQ+7R
pigsS/ecmSZsI3G2M1MhpcsV1hDkEqzhJyDVB8CYiiHt/mjX5IonFWQgbxUHdm0U3818iV1cshox
iJZZkmJc/hVwuKrDgclGJ1+p6J15CWEJvzjo9/5oh6ARyAeDKxXRf1PuGhOKgzneizZqSUI9Hx0n
tAJAiLmYjm3O9iHKipua+x9CgFaSPQSs+wyMeniFEQ8carpYHokzGETQy7gVlCd5FGQ/Hj6QHztv
HXxSlwMjDRMrL1Y5B6hgWicFnbnzZtBwC/vWLSGP2wIfVN+goVYJc5ZTfspCGy/hfzVEmHzEHcnO
QlcSpebylDUipQkbkTYgkqCeaaFC/Ug0KIZQRCoh9+JLAcB9syuegq+YZ1phaHqrYmBDwA/rNf7Y
rDjqEAljOTWN1aPsDdfsUnjYb9c+F9ypCrrOj5Ui8nw3ODQj0noNgS1qRb4oQIQaAnsjXD6TOCCP
Tdg7G6ZdhOfTfJCeajlmst2TjRb7gZdp34H9rKExIsVENa6GgJAl3q7mQeLJPUGVgokbF5yqAB/I
SepDs68+Aah5Bp1SI4ly+O93n0f1Ikcmh6IN5GLONAn/SGV9OpgqDE6m9vvSns0qLCpKJTb0lp49
1TN4nKqbhyC3HtCzxoQjFIdouHvWwUnQBmc32L5e2f6ndAL9fm5B3/hmQAxd8yh3Rixux3kkVkzG
MgS6JQ5KG89bYd5V2Fn4V+QbXV37x2P7ggt/5FwRIFfhFUimimSEhfFdywxGp8yc0+pkZLKcUqtV
wFOj17GTkXeiJ6dFAzxJgKlq9JBB8eGGpIjY7+/i0kn0cAMPsTB/CzgLZ+l7hTw/I/4Wz8yKAccM
bCrRnPff0+WVTs0jFDVipiz0PU/ZpLUNtpFU6UF5ttaySy9rP94tiOOvNxWaBQ36a1TkvVMsRbxh
enRKNWSnHPN3zxuuFCbR+gf9zyoKE2EhQSGwzZJrQ4vwyEQuK0X7qkdUXycAHhqPh8bADrttW20Q
NGAIdVxmMZjPBuHQPnUsINUyoJeSdHojvXNphDqiEcpNyLs0c3j9WEZHOMP/X4liNkQhNYJt7mzr
D0NcjN7mxfqsYeR3sakTOPjNqmvwB/OGuW1U/IwllVLYwlRYV41KGtFZy4Vnjg6wv62je2Tyn6H8
hgxAV0XUA9vDGR5zVf/eOQ8IEAbsjLxL8Ak/jEQTIZ9f+QXUiBmnbYntBrLf6vZBeNNyWyGUj1Ex
EM6K7i+z2R8etwe6WQ27PqF3bQ6+6ZjX5xdBsRJDqiFh0jWGgRX/Eswz3xl49+XOUitZXUnvZhnV
/ZqLD4Mh8yIcavFlGz/fjDxJ9/awLnEJsnY0YkGx2paWJqtPzeJixzglXn/TPx7t+W6wjNoF0xrQ
4oWqBOQxoEJ8tplqGeUK5HrO5wPKRgD0WaZeklH6FrFN378XgU08x8MoBY29wXJj3LuuPAM7/TcK
9d+3QVHmHKbxgvfHnQI9nnxbEe4vX8gNRH2+55UQRJX+O1WB6a5neerQC6Ui5nzdRtgozqDAfOjR
0QwXrE7loBUxjn3BbGovkAaiSf7ivFlsqcojzSxavrO3bH69YFnUYKsVbb7uMO9aU9GNKa18qBNH
WQlcwrdKWYILmIQ2y5GcZbMCoyuzA026eDHaONf2LueBPj9Fw8YWg4IlQDckdlF+x13Q5hDjrKC8
g//iVUkd8g2hzVcfIk3rsjccSn5+i0Y/IYubvIARHxC/GMNZEvjAFUF/tM3F3Tz0azASYMX1C5fX
JIrOy4LiijWzwC62Pg82dSCw+YN60tc6z1pr7UdpMrsfoKu7ZqyBYK7OgAwhkTtLJv3xI/06yLYy
xvRl7zZEF8w2YS3qpXRCFxvw1iRgU2ci3oZ94zeICDnzGOlJhiQhy3UvDovzqYwRirZoNp8v5ctg
oXai2YuEcaUGoEZrwJJsECouN9CnE2EvaouaPKmYZysrJpJu4WR4xNuq5UvTaFxX+L7LAKEag2xj
OnawyBFRjnUk9GMu8R/x3rdDy6Yh3qN/nB59kDJS4XALwIxR/6+h/etH95FVM3yMyIy8L8PjsNnJ
JwBAOt5h+S2pZuT8QKpgE6Ti8dnyig6WVLD47vOyXKo8HfTh5VVl6qd6O+hMv3sndsv+PXBWg6zy
jxYQ7JrF0AAgixZDevtQ/GAP0CS9QYf/uZCVFUOcIAwnRtBjFxXl/GFXdR10g5CPSdW+rI+2vbZM
RnZFRISHBXKUxSSqeNwah1DTCQ1hKAdSTMgK1L94CvWw4eVL9la1zn26RaSsWsX3ouMy2x+uaRSf
JOV0uoc+Dq6JFwG+vwMFCr6Ee3Sbj2M1dbJo0bEkSoHzY98aELZZGcPgut6QjcypuOfyuhvFm0pI
P6eKzUIHhtJNg2kPLNC9YQXpiyLfbWjsFWAR+ojFjp6byXHo933WLhh9+OUlDFgfyZpOAMHQeaM5
qGaZ7DWn6v2Tb+a3fX6Y4BJeRenUvIzBtmKHYQcTR87X9EqCk9Qq7Kcf4IM9dZKMywuv+UCVG2x9
zSMnQti7kLGnbisGcu9yytKQOyIw7USN6VT7uOCODxFdLjXO+Mrojhmucfo2N3oEim1vEFMIiJ4W
m3uDU+Xxp8lAOHZNQmMopQ7+4FDMNvnkigWOBxjysrSOcMJTIrubnrMXi2W4I2HAw7aE/pEfR5II
t+GN0ZEEam1kar4Emac4Pbr6zYcg0q7nkxMDqjlJPFtZXKgxneG9rpQRPM0GOhXDGQDXAaWrZUAV
44OpQ0n0whHYKBFGd/uCRdJLh30Mb31PO/gmcBa7h/RZnQPBtlv/FC8zdQ483bQ0YpivG8U/Mon8
C15roerpCP8P9TXulnRkzuDTQFv+uJuH9P2akq1tFcEXkvcV2BpFO0ZMpwavut7ySU5MqVXhTfK6
KRs+1wxzIVi99qWhmQrIiqQ8mxItGBDGYkNJdoNWfvRL21RmiglPvSV8FEKYb1QCDdiiHkrDEi7/
eyFYpG8GsDTI1SuPGEWdNNFObDyet+A6gArElbPGW6P5T4scOO3v49pDv8heoWsigljWKurO4RTP
EOFTwx5wEZlT2H2HlHRtfk/25iJVBEV/aQ7svEEJJ2/TZ/lbTO755egZQuyH1dxnrYclgljyfJyS
nhjbrsERpN/FD9YAFfoNUDf3gCQjbzzLYt/+0UNF3vDIHFe4vjLjLeAJLXGY131OUCVdOP/zHDQJ
cYz0Mz/gXDEGsgHzWNLb4Sk54Sh9ccaZ5h6PFw1nrw9ZfrmwdQUuPPSgF1QWcvGumHyJ7Na9yNbo
K1QzeTm3e6HSdE0YhxvEmHCrn0Ey8lII9qcJmzVhOzqJSnfIt/z4b/0RkBMGd+Cg1bsmdGKPL9NS
+II4vu3qV+IWlEaCi596Ov/bJnV7ZVuUGEDgv1+eDoQZaaVy1aBTYmt2Zmw7mrcIDJpRZXwvyOLT
2ogo1f6soEw+GEMI9aIUi7n9RENAvFcK3hcTosUmL8mg/ub7lyhJEXAncEsp7+5qWcNSBDAqC0WD
cPXrfj4t3Bu6z3SmDL5IGJSyl6v/nFY199DeY7UJDnoVfgYMNCfZ2aBxzWF1+zZroz+81cmg4V6J
fsTLx001S2BJxdLSxsW02QAc5/lgfuKVcRlHii6gmP4rfPUZyesR653c2yG20Xner5W0JmecQc0q
iCLL3QCIgmSd667nUusnWuYgzs+puXbeBTPT1tB4CJZu/UdkAKK7FgbmrYiAdAbFSbX/ZgMswwfc
eicsMQag0dkn1bpwbkS0jgw1UKRfau+VB+uvagdKFf1cISa/SiOSXFO0q96U3AhpUSU8x1D2gLKz
j1brMZuOjQhbFBqUo1uiDEC7V4A2ud6/W+nS+Cf31KYI5hlvaIklZMJsCoOiUWYx4MfomkbKvmtB
ahY0lUKS9KOQyD6jbzkIObGE8odSFRS7hLOhbOQlZ6X9BBIOk+k4yoqAZCwf9vkhxCFtL3kAP6On
IpOb6wByY2XVITL8Jb3WfiveySu+/ssikocs2D1H+RXn/ka8HM1gSwIaNOlmuG4qsLtCxvtju5Cn
gE0H8jGzh/JDunGmLXiRfoiPgfB9g+Nrf+dykiZxgwbXV8KoKHdVxfcZ++3f+b1Ej1hrbqw312hF
K8LbxKHy6fc/jvYxyhm7u4ArVBBWag41WP2XQauZCIOCs+VzZI0vUdyaKTYxqezAQiDGjXhQLF4P
upW4oPzkGbF4eFO49aWHY6mbHFmiQirhOLt9eGFXMebNbgoFYbjHB+SeNMFc1ddYdrXm2Q+BaeV+
tUVuCrU3mFjpZlSTcb6SO+GB6aG5TY/Ch0weREfLbdiYd1AATjNpa4yGdp69Clu0bOHjhnNiL+fT
BDFwF9QDaKO0kB2xKIK9a3VGeHYqze6wounFlul6AB3xcSkrozkBzgIvwoVZprPMsT2kqcPXQtx7
er+pTohOmyOfpIpRQm7SnTBHbuGcXGbMt7pyTErjtHbYuHw+82A9jF98E5zAF6Dr4w+JiupvQI1c
VdDJ1EInRdjmMO/q/DE5jTUF9o4LWyta5tuNRszn/DVywHrps/5yWGeQ1VfFnR2+weWABT7yKvFi
1CjxouMDI9UnwifwVd8V7hY9hRGODAzwypDWHB4XQeu04AYQHRX9OSBofmEgxIn6SW/VqEZk4iyC
426ISxbhIdUViIDlaPSFfinl0NHzGKbZzVH8dQzLRAJUuK0PafxDgAiIRGbMf1Qz6gL78VaDZN66
kExO0/wkcOaQkPcZLWnVxFsFsxkGY+Tz5L9JV1lGCUnvSQtmCQRzHe6Yfm4ucG6I4NS8HnNVWF0o
naczDLV9G7WCdUYW//i3QtgX3hMSAk6srQbNfiuDTw/X4VWvTJBvY7wF6IaYWZpJ/b4PMj34uWYg
gTCma8wtR/LHCxjKwrZXjgyuCYOUznEFgTVGeBGMHvZTyoOC5LyBsHTfw3r1E/MZY4FHbULJ/1/p
Xcojd9FDJ7/Np8xd5aLnmTrZoZ927r5G6OZpbDy39aMuv3juO+CNv/LNXSkCz5fNQv0d6EzNCzT+
3zDUEi2oFKcZpOvbENTulYjL+mwDnMBValee/dqI1VXqI+QOEGV0VfrXcvRtBYnsZr88pLa0NfUq
m6WGF8kcn91ZaPg+tm6yl9Muc3ODSn4YBACDLAN+uYdsHh59SA8Bl+HTqEF5G2gY3QWS42kaYVbN
oHOPrGggeB3aSz60TTcHIlX6DMukGBFQaDyhT8Jf3Z5be8pyXKm+u4jSSdWocBLJnS9zRP80i2oC
DKkOUuVfFmzonUiCJqstJrmz3neWjt3liYKE1mvuaj1rETVt4GmUFdymw065j1XtmpZ4f/1SkruX
CYK5/6JTLvqtssoKR9IQAn+7/wjGSRtJoMn1U0MlbAnOYFndsi93GlFXuO5EF7w7W4TWpGTbC5uv
W+cgEYMPEJsl0nUGxxHwhu8AlwhKUWZUeSECNdf3utyCaeKPB9dVpxjFI0b1WJpf5Ah1GZjr/kk3
ECn6l9FXgbiJOxw9ZTDYSlALiuaYtm3DNqYlfCDeLWcxmq9RSEkKga0KAT5R2xN+IvjCv+y10UeW
jyCrFc3j9f7i7iYPIC09hhtwrX3c8odGufUhjOw8h3kgwDKuGjxjxAAcwHNCcZeF4e7TiUqhG+bb
OStwgAD7oNuYaZygHPMlC/m9TNf7OUduO4He8hESqoJwpmKZcFtSJklOhKepvIWY/eNwKpNAeIkN
duzEdG47Id3mYHqFAlEcbP3M4wllvlrkhwwehJfKae5FUgVDCVPTVYJ/3+eJuYQF4YUCWZlW7wQV
LvdNleK+XcAFBTox9JXdZbqeLYg6s7RFBBC/yvGv+oqTEbF4buvnBlQgQMfZH21bFR9GMoTAsIGj
W6MPwtVIVb01N6de9kQTuu6Iecmehnk6irQZHw4/G5S99mDmwytCQV8g7/xEs+dw2/sTRAFE1Ozk
U4W1OSciVWnMX+WgsDNYknQbDboUs51Z6TGBgIvZPdOM0Xuxs2NI/goXBgvcUwbKHn0rTFBBtT27
ywX/Vi00KvN3qfrpHWQzYNS+uzTdlrv9oVs6nfCOU0WFDtfnTediH+hBsGzI3bzJ0bOmTmj1mXkY
bqdIKM0MUvxd5yOj/RCTc/CsBJ+yNP5k3gjwwarpKR8M1AwaFgtj209i7OgwA4JuDlenkI2aqlP9
yWVime2AIgA9QGWnII+eeAkb8+s5kdvc/3PZjmDdriBv9uknwuT7xAnKUwlvfYBTJ0Z2VJs7la78
FTTvgQyyoNX7Lcbz5Mr6X5Vx6WBFip/l1i0rqRWTS5lSPBqwgbdAFijYu5VSr89i+adpchJ5nPY1
EX1aJF/vZQBzdyJhx5XqnF3tGNeCW5hCHC7jh59T4TqoFojppL56js/xf5dYGhMeLHhUBuuvYIc+
RNYKhsVTmrBTf6FeCUjnXZZAElikSgnw1v8B0HkC4fX/MltDMxOAvcri+spDqGEozBQ/9uh23VGq
PbYFqeqKlTYavtQzsuJDsyDyetTn6hVit4/5mjRqOlv+Nj+ktJGQgQh2llZ6sBV9peKQiFz3dgDI
tLCHUTTvi7MM+cBzckjPI1mVpQLYggf+8mM+aYTdns4bmA9sJzItwHO8zLQpp80E0WWdjkpBZN9W
2dfHwiPVHNWNa8biNRxffgdHyy97J8+ldO2uPdILIs6imarXdYPBUmvFlbzmtr91Nn72HIMcr6Pw
p9rmmf7poAX5V1EA7u1Ba7/dG/R8VFcGn5T4z/BeE+AsE0JCFjRvVFgC3DOczCDKw5r31LzJGBIF
m7mWCjZBwEbbE0+A5xGw5nKYuNwWw88GQEI5jrR8kUw6QUXGfbuCo6eTLinUlzCFZaGPwjMwoRE6
2tgprUpafhMoE5ZNforMnXwPBYKJzvfSDR3ozuHq7K5/9vhxWkMeGE9z7VvxINNSrhaySzd8EIhk
NSGXh9yb1yG0gLMbT2NsrttsKWPeYrDteXVvqVk6058ehZOQ7IPW1Vk80s5hxwr0hq8+4xkd0l28
pA4Wbcizy9kbkbF+9+UP+2XVG5skeJ0xiwJKGcrrzsyY4VUy842OfaFMPN1fd8DzJ61cIIeKhR7E
bdcp/E9EsrBgGHa2dJ2XOIku2p+Au4+jwR8zJd2fnet0H1Zzv2FynyVR3+P62iYHMMI4a6GNpL9s
OYlWy+n4nGJIa+5+TNXMPbbb4ouS0ob0Xp9UADsn3OOq5nbfGLywW/cR8neUXMaK4pHTEx6KMJDE
SNQNh/BP8w+PvNTVRLvGKi3nI7/UllISEH+Kux/s1x98AWbvRtFUTtQ1splUazps66KTQXbwCJZS
6grE7pf8HIFB23K40UrQPwWYQYFLDQ5HRfozYUk6FhWoYJTMxUMWAvB4RANPNYYwP0GrAQivXyqg
xXAWM7VrgepIaYRUom5qx2aaYOqRZl0YMsQwADBHNcK1C6FhqQdiOaSAymvHo3J45bMRSKj0S57q
/11v1BT5MbgmKbVqIVgzFtLcO3wC6KAFw+JwCm815fOWiPkbzUU7rnXdHPxtcHGxIreeQlgzWEyU
GKF6Ez8SCbtSCg8bbdu7udpYJiDXslWi+/nXEQIXppvTnpE2SudAxKhsN+Zgo981h5cuD8TaEMQT
mFgvlMEw9rOLPUnW5/zRC+IoHbStroqz81bxH7KPMWpcM7aGN7LJA8K2OIfPdfU4f4+r22cU9DmV
GaKX2F2bVnxxvT2HIjUqC9gVVDl2DDnhomlm7OLJPJrLuJR3UzgbPei6qcE//fby+z2bqNDU01fH
P1IpdHmBNa1EdWN3MrYa9Kc2tMu3Y6l2IxdTvyK7q8CTR/ixyzwPo7/eIyTKLRk9DHjdbfvFaVhw
oKlUBmYL7enmvCKycxZWAsqNwu/rYWH/t5S6oGyXllEtTZn+khnYPT7vx2ezSzCFksTUlrnMdl5L
vyEuF48oL6waI1AIoxZ22VaogDbWfhLzDeIZgkaZJkErzUSFeCw2c3+IyqFXh4KIUF6iPRogUlwX
X5o1pdKh8RsCXpl0njpDJBj/e2Lu359PhEWhokJx81hlXlwf4CdolTeQQEBo6fUG/sGs60OsqYQa
yZMbvLh3FHX9U6Gy7p7fRal8oD+v8+O6XfnCUXu9G+fSnujMC2LodUEHIl4crRJSqIumHb7snBol
iPOTjuqZzvdPgvNKlHWbegImLaJi2E8jLfTyY5UfbswlljPwgXiyy1lw+EWMQ/i055K7si8EXfyc
k9I1Nb0/Hqddg7j3Y6/0ocpLe/DjIXp/MLRb6w19OJc/RSCMCionQq537Pxnw1Gr3eBNodtL3H9g
dn0BYOCDYaZErzapm2oQGmwYs/k3nnwMM8xxjcCTKUx6KMPOH4Y714pYDODTKIT+Yf9BPhkKNP8i
jw13UwZqgHTeKiMIYFOByLqJ/Uge5r15Udkyh6PLrilECsyeyb/zEEDWyiokDjdU9qaXyaN/8CEw
ZQsEPsOe8C+tnKGdnbfqolmOk7SKSB+LPt6+i/V0urA3yLcEPZNBaIAptb0P3Th2Az/grLK9PPjT
ew2dLppm28rWSHBvFMGCaIArhsCajcNx0aN2YG4ArI3kLCZWivVPhkzB5bbu5jdRHDm5A4K6sOV0
+EnGKxa529/eEzcTjMnBNqds45iNWb0y5e43oiX4iu4Onqh3CG060wsCg6zgNxUwTbJtjyFVQNY1
m6kHXBBUglJ8DUMSG+VjMYwke0PYjRebpnoZaA0e9ZaHKRErtEjaohF7GVNikCZVRrr5f65/gzdE
9W6E1VUeKvaolFGvz7sYJivlnLcWZTjYu7zjgnSar9Wnx2LMcFpvS+GcRQyff4x0xeBGbpa/LbfP
9jgysuKGWV96X/B5PxfgqbdRnZeQaBL7Xszen2OrOvPYt3aAvAehsRnKz7U+Pqf+u6TghbFQCRUd
91VFHNaa8mC/ki+rjd/UKCpAENm8xzAObl/y5SRyChfU5SUH3aq78ynK5zSnk13XdGEK4AI9PyGf
y2OZWJa9U8bypEBbWcCxdpD9fWHu9/eTd4lbU39WtgMpbEFScHoEjiBDmsnAGWakIsRfVPWShZly
iiwP/L5528DgUG3ez98nPQJTNOINFQOJfVQeVcy2QugVH5qR/yv6V+OmwY9CIEA4eI1e9tjmmOOg
BC9JUIT+OyKPtYIAKDsGl2fNyQjdkgHOZ/uiteSw2hvrkAo0A4sxJARTnJSygy5RiT5FdAbrZI3U
i8kmngEmd0yi/9SQXB4Z4VKcvAHuYlAEd6GrBewSqCUiKY/4nv45QvXZVCgw7UJyYOrpRG7ZbsKa
l05bSv6FoU7vCADU5LqY4DVsQftY2jWEz2dvuZahZGFn6OxtwFmTeJa72Npsd33fbDp6jyX+IJsJ
kkgLdQV4mjSQohBQhDp75OfnpmWzms/bj/ToMeRwCPfTpzKSIeWs2FyJot2b5Xlr8tAd4uJf6/XB
LaMvldof8n7MFrMJ3FAG+6xeNXPcaUyVu5pRRd3IasDp1SlmANqyjf0B0fBlE5fCYptuxEoIcbJc
hVhEkKMpZWZDgdtuJjYqeHpjfC9wkgdikRwTqLG7olYe4wBAxilZchIFgzMCDFr1H5BgazxzAaXF
k1ctfqbfRC/6IAHyDGd0K5llTOItbZTIIgjM+57+sM7MYs1mpiGhBlfWu5KexcG53zAP2Fv5AFxy
mdN49kjNwe1wlocUFxW3l5Ev2e06bAJZnRyvQWbKrrGETDLPpTuxwRLtX8unO7hpvmD3hnJKxepn
gf4j2K0f6UrzCNSkfY6ZDpaSE+A+JE1KVwDF6MMYMe2TXn9rGb+IM4k3OSqwjxz4oKSJPkavaMXq
VqdnOezhVdxJy9FX/SHAgR3GxsFzzMUKFN9O/fmwtAEmKz+8pWMZNLDWYOKxdusO03jJaWQFrWfU
TsS1XJ+YKvbhfruK0zwMyHt2j6oIsqGxWsqEVr8C8luZroje3oOB4h05NPYDczfmGRZwz+116K/3
lyZf3xmGCZYJ7oJhQbgcmzTVmTjAI5LQw55vmPgru53COuYVbfhdaJrWMJpvNrNq5Os9N/PjJTgs
Lf19O9DMqcHRIuyS71a/THNBJAStCqhkDHIWXA2+0gacwveUaLm2XS6fai0AS5yuGaN0kq4UDuDC
WHtvLIEYDFznYnIMxE+gfbqWdHUD/VQtvmDK0oDQuN400PjrkoJ6SPPzP+cv3zBndjODmzeio16A
sSD1lny6/nvefDhycwtu9j5RqT7v2qIVXPW70crAYdcxP1qqJnFUvNgjlTrXi2L+tf12lFIZfRDf
BzkprfnAOi4lhFcVw1Adg3YHAUzmnS3Yh3iqD/awLfmD1ZrQjgW8+FPWmnMBNprxS6lP4M19D2pn
rcXVR5qBgR86pUa5jGIxtks3O15LvShaf2K6V4bCBpjrp4M+U8yx17ecw2EsQXLAR3MssBpGh6AU
2x8xq3/hj7IdXfTnCSeeFD7NDvia3uQ7p4sZKxBMYHmbSKtGLJ6h+dEssUuhLBgkRXVpOz1hltIY
EIk2i1nYN/Z2t1P7BWjmvih2Fplzk5oGQaQXO6dBCIsgJjqkzYKUlRL2xgVZASsOHf0YXZnK0IKu
6eTyI5VEYHyPYIBjVGmeFSvCfXecPpR6Bx4XU2aCWXvxUctBAmL3WxU4OwwsT8FzaQ2dlb3NUxQs
zVUCK5OdTp2TLffueVfr5Vd3TWmQDwCuBTk7uyx5rIl5VKuXHC5DO+lzEWRACeUf7jM1xjfqPMBz
0m2tJdGmTYHFvl4jjon10Tt6A1uLuXxRN009OEPH4DG/f6wFWWl+VAk1u76xU6yfdZhxSnR+jkbz
tt/+mJcnPxNCRfYBuOOlKHpKV7K8DDbg27x+lqPjatS3keOHGN1LKUdgSmdxTU6U0SHkX+5HrWHc
jSM/l8Hk36VcxO7L7yb6Qx6WsxYu0ve8xOemPRLZlPozlgobkqrl6vIdJW+eIDOU6QIBT/LAAvto
trn0sVmQo2e/QaNK6i7gPY5O7FeIeB9/kwuFg2ij2j9aQacFlnMuIPgHYtczh6C1Te0Aa50gROUn
T7Abot1igRsPGYHcjNEZ/yWvKCDl8y9d6KjeoEYrIbJfqlPiDs8enYPjUbUAT8c0DyxVizD53a2x
iWtVCvXD127369D3eJefEdki/NYrW8G8oHvd+zrcfcNtdRjyLlQDuttVao41paHc85EPnJ5ExzhR
8Nhc5PGNwByorMAh7489VuY4opgsVkcU4SJ2rA+9TZrjoTzkWiTXsPkPB9Lje6YACseECbAn2/Q0
oup9i/qXTWw+yLVxvTFYQxUevIWIxvByOLSw+UG5dYyYKg/11dlmTaTkmsnKMc5guORKquw+z0Rt
JmMSmNR0eNFRDi/ip4v6KbLhJk8X0Ate76sSjCmNzcmZeeDdlQUNe5DjzDUjIT0iCem/kRHN3HTm
5h0pVLSa6EUSN+grlITmuWmwmcWi3b3vZZ74UYkgqxeEewMgZPNjO14fJfufGEWLH2Kxq57DzgIy
HK8AFRtknec5Mk4dAFY4QWi07WsGLUHI28rwyjhzPMsrGGDXkSozZdvV6VDtE4ep21NPKCWNLMVW
UzSRYf6/TFAm0SisAbaJFhEKIr7geDjuG4d3FBPC9AODfxcriizRr6kmRXBg6s2cvo+mUTjgykME
aoTzwkSeHe3uxP+UQqWypOWV+0Kr6kl6+c4IY7rWIAuyokeQGrgARmeVE8ngvA8kAvBSMlj4d67s
bOY/jzgPx734ws7vTh4E0i3SZsprCng+1JOkeXhcFRT6LydlDxYVh4sJnIPQGy6khBIEhYOXZw9e
R6bx08kaTFikq0xJjngg2HJbT1KuzeRhtjNqYiLtIXfP15PdRvNNq5OMCZU7Ec3ZJLvQOj3+tYJy
3jvtMfvJjLFDRGo3In525eYrhzmQ3hrPNp/DJgC/LoC5MFBDgasN2r2KgjS7dzYNCdp8Qtr8ZYZ1
zZS6yzsv9ruu49mpvX5IQ+IetLPXapsfe83ljwNuDtQDbgXqVrYWNm0yOhDeKovBbIaqyQ9APl+/
l63dgfgnDX9DdBRFd87hmWmImsV/xb/CuTXr3cXIYyo5m0PmoSKLw7Zp1bs0pBQ3LsX2DkNTnXxf
Hx6SGeYcpJY8k1l7+YvvbP18mGsa/jYuCPRQucpVrPpDy4Ltv74tYP331YPq4OLMlDX8wiVrUegL
F/TA2doEiZcZxqrOaFtFSELium5PkuUyQ+f6BaNpyoncyxwROmxCakZtXZu2EBcqqzAIfdR6XbkG
t5bgouJ8NOjUE/dcPYYksSfAzrz0E8Gk0XSma2q8RwOMsrxVAwTSr13MLOKlEXESaDeu5QX1UlN7
VblvIKkRIuZIuvMAAHx5kyBo+x8p0r4PU/09m49sunN8zNLRQ6Y7tYAjONl+z+LcD5N9C87jykk2
pZ7Eft2BWFGTl+jLsb6EwnsAPJbTO1kdah/JD60myuWfZCXDLV5ijUKl++kOqLhsVecYjU+2DQpy
wvYfsRCtTN0zhCMddj9kehrAHN3W8JUb0+A2Boh8v5tKusV2d/zexzRR61L7z/5npvng7uG1rhSS
vpy1bYSAEkmEIUlf7v5VUZMA9qBaLaWFhA7tcFL7d8afzaohQQU4gZuSYQ+NShIPOZqPVqKvAT/Z
3lFNwFw4bwa2OHhNnK1v3zX9HOb61k2HG1L8VM82vOHT5zE5hSLqGreBHFs8z8r9sVcMAa53RXb1
JMbxXmpEjyKCp1u9VCFY+YuVE+lz0H3mXTRW3yCHKj5e5dQjFsQMsRZFpCfQFzGCNRxEXSg6b4pC
fYn92C34dTSgjZwhxGe+TeK9dY7Z9MlVIGSd9R1DyNyw8k353fHHEin3g3yEehiza2JGGtnucl9L
ZqzDiiB/mVEWIGGmUqdYRemBhjrfpgnPLfV3gsZkbkgXWuQUoU66lHygNhM0TsXEESqxEgiNUdBq
n49U1IDTVe3S9fFemhar4092GxFsQd0NlBUU488c7O7j8Z1t/Lv1ZGkJEXXus7HPS03wfUlG7vzS
jR+Bp8632jZMoPhHOuVp/0KJ0fvVyYdpEOEvnMFkSWnSA4UtdB6YwFLKad5MWEigMaux62tksGpR
GZOQ2aKscipEWuAlJIPg3bvlDjuNEFjZqONpK6EV3VezVSNnA4xG7nujcBKtbG9LN5jOYmChrDrG
OXzQyssWlb2puD9cyyk3E1nbn8VGgHmIn3Sxy8fBNGspC3DF4ZN7Tve16v95xq7s/6lNYXOu44fv
n3qUX1S/AfJwwf3GXtKOZFYuvQNSVT/RP1XOrLV+e5J6xjFMf3K+vjvFRHnnqBUeNtUABJIwDnW9
wa6CIfq0hLzI01uDAiM2ECessqbKQ1ST7bjAMlo2n8fNdPmO7yr3D84Q8tbx7k5lbnZj9r3Hisjk
kgRwlckjnhED5hNiNjkc6YwOhmjhF/gJuKUqP04+bcwbmD5yXcOIBRUQLsIvPwAZ0wLraM1lU2RT
YoflA42WqKd38RHrPw/5ti3Yl/FWeT9WPJ31Fj7yvHo3Yqb5IFEamnBHpDo3I8wmnIXzWb4ii1rO
8DUkHkZMbZDEf7g802KMm4tPTBi9XpQJ6N/fVah+TQIoESmut71IA4p8GyYg9m0QoQ4M9DAJj0VH
6DNQotqpwcNS/Na0hfY7hPKj4OGru+gAXkZq1LqutbWCfNynccTlByXaeOl2UiLCmhahaC1eXVt3
ZT8tjTgIi+S6bSmaQN/wZg0yrOSsKqp0ACPteXNxVXdtOn+8XyvoTJ2+SFuJNKBh2GLEe6hJHQPS
0fUX4o0CZOKT22AslVnBaqL2VCTuOF39YxnneISrfU4JhxM6gRL9RQkO0BMzzS+lGmuDz4a9Jn2D
NNhbSGPpw2/kmVV9axm78IdaXcdTuxUZxH89SLgnYmvkuCS8NckCb6WJrP0cYRs9L1VAkkCuC9w3
N952svhVPxc1YmmBrgERWKGOFzJKhnxAPYHSMrD1THK6CiKVlg232tEXDUFgEkRmtZ7QWoHhHy1p
Jmaxz050bM7Pvkb4hW5yIsYOd0Za2QnDlSKgGEVtQ/i4aVN7KxERHrQ9sT5Q0aq1vQJC65sYxMt0
R4R6+zFRJhgAwpSm1zCLixGwt8rAfJt0gePi7EADnapWcCl783iZhhxC4RvWgc84GmsC6wT9e8Ln
y6SD+ZFlQ2HuzS3vWWaeph2dIcbwQFITKnX+nLg3ZjwHrB6v78tzuDW4R4DD2IrfVPZFwK4JbKHx
k6Fmv4OICGc1sixDYV/WrcvYhH1CxAzt/791QpdCIZkTVXypHJUkGcoS2wV1LdGmF0f3GuHgNEOS
bL6L1OPDSoGxio8i05vfzyxDOuIBwLKN3R9WxX8t70ZI6E7OH8XgYyIhk92fma72vEk45uRKUveM
wgg7esowHk8g8TZwMw+ciDI/qbLIvpMXJQmVWVfLci4zFj1hm46UH/v22761ldNgri7J76AGJ7ru
sFK+FE93ZNIOp6WeUmS8JKHNBQCC4PCcQAqzTDC/5ZIPtdS+kuY3kAoJhMf2HhH8Hs2V1/Wl5313
SREktiXGGBC16g+D3gvgn/e9X71kovmieJcvebJLtMr7zcw1YqOYW+1VEi52ibgTQ+jMYbFRRy+p
7DRwNosCNTCDHiDcqk1AqsSXAJAuBgeFANYpp5Ml8JvCuIaJu+5eTjLclcCaI8M+0WLlwRpGSbSx
2ix+fsR2JGW2uTqBpvZb72UH+38UmaB2tmipBVdWF0jb4iOTdpKPPTY1o9q55BYyBNjtWPHGwICQ
W9+iG1kIVMfWjLzn0g3RTwNpjOd1edGXXYKYnvGahNN5c3UFz9lLW+XjCNIhTc5wHykZlvU1yRYd
F4NDg1RJh322AXYDe8qjvGbFZDM7najSiCnB4ZGzgbeC7LLe15IX0liQ9/Kr/Kl0+2IHu19rVonW
TSeVId9NSg5Iv7es8ORE7HdUVL2ecCqRsCudfcJbqdv3jYpVqo8cnwSgkmzx55KIG0YMUUeL7ZtO
dmGGZJzVk/VrN+8N7gi4lRv5rvao5IgzD28JyR7YnKLFSUTIcqaChttFFaL7ewUmih0hor9tbBii
sMmKXMVnHNtmcIkR+h9DaxyJnJpZIV9CgSc064m3tF56UQBxQEGrolzf7Eh8/wwQC36Ik7Ey/Rgy
LNaFidhWm+d+Zu14UtkhhzES4dExnFe2kjdBCyLkcOXPAB8E/3ZPaPdTSsewg1ekVc1kdD86UB8m
yfe0t6aVj3pZz4OQ4vpfK/5VJr9ze1RYNguOalb0KEryIqOSO2kGlRTiHz7vovtD2Ag2ehKtGPj5
PrajqqtjVjdAwcFlWeoc5y9h0fF5ffMg7y37M1o0R5Ub0okMwZQzN12d3nSHlB54/8/AHPvmlvcP
iyZnk17XhA9M3HL414tbr8EL9idECaEfnaKeaxBeDNzUdCkqKtD0ivUszuQOK2kiitLW7xTGHMmk
koFvI6rv7RFN7nLQlWA3YpF/dVn9pX55fEEdZptwrBTmgEpvOouF0oK/vKH8MKVhnUT+KYmUpr4F
/NpDE2ZT265KzNH4UVZA8KCuNKBSZrQkH/eup2WXkDHm6ArgyriZrTiPXepKoWSN/J5LsNNYa0SU
zjXLA8ymsG6MbGGZIxQtpQLXy8M3svA9ta3mZi9K2AKmx1bu90SXICRJyuJxKPXsaauWb/jfJa0v
lZyDNlhXnt5POUOmS5NSTRCvBkNXi7E/RlJufozO3CImzUIECI0JCjaNCSBkeRe5QtJfCFiitPu2
kX9GJVZr4WHQZ2B2uNKxJBQe74aMLASVmuyYLMeBajSCXIXwDnQEtYxasvsi4+81Ig8JCIQHkENN
gy3j8KfbayRUDK6sD0ZBv3wX3Yu9Fmc67R7AYan1L3mMlJtkcFjA1HYi/rcSD2zQa7dRqDItUjrw
QnL1j8y9rE2i/U1qfQGuF3VAjNk1zlmD06UfCGg8U02QS4VpfnuWUMDuEYF79RylO8HV/cBz2g6w
sf3hfKyf2qFRpdqCNgtomFw2LgFohMulV2lXHHnrsALIx/uofS7ayZrNXg9mFe2r40/BEmG/XrhO
AIoGfhMcWSKDIlc5MhCz0BlWsuFFExX5OlYtR1P0qU8psDgUgjfG3il3YsJAQYnwPB8XSFMH8nwr
5Cq7bgOIavo/BTa3EOb7wIgS8L/WfAPLk6CZet2YN6dHIWRV01hoOEakiNeBvjj/vICe5+TwLFve
y5WjgqnhmdB5RzZ9NYrCDHYuZTaY96BKQmpmbwkT/BpSJeK6Edq/d+B6fyQDJja/vVXgyIn3P52c
JT+FbZvAfnj6Ni5LTBqPSr2lBaDviSV/VdTABx2vTjau0NUH2DBFEf25eSXfZK4+LVXS7hppo1Dh
ODTX3VGc+uJHZzFtdFgiDl31+I8nge5pwcbc7gxDcR8Xp1NYzVXY5n99mRPObJW3wfA7xj82g1iz
wzfBUqUsfaC/IcQWt39DZaUymJK7HUzXiLXT5NjL79B1qYw7Hgel0q7A4nw7M+hRKxOMsT66laOZ
fr0R36Q00L+oqmcdZtpH1yz5WcXy+4tBDMSp8r9AxYl2X488HqQ19BWYgHvejFQDhlG+yGO6n6nl
6AFcRiOsCR388uJ8trsCoyIJMur0NOCvmm4JwJu3Wh3q5JhbB6nmB4I6r6gxiEKxd0pRU/raARlk
lCiXzigsPa7jFYyd5ovyDdVBlpt5qUgfEZeQ1EwU2BIuARGw1sftWlNkJNJMZ0BWuBWWSuGkiOzZ
O7jitHi3SWamIG64NFJB/N2SY3f9kzQi10Rnk13A9CbOsJl8WQlUF4sBjnQIpu2dTEctI5cOfF5x
IRP0myhUIR2Gm+XTNYR0ZpwEEhv29YHUzQg4amBypCnNqDWWOD6eRKusU4blhlQ5NXuJYjEM4UXI
UAOYAHbQkZ0mmpv9EgBtJpISNSwbqU31fneUOWP10Bh2TbSRcOlHdfoABDcOH74Briq1hjUSowhM
DtWtNk2BLGqWbz4Fra9Xc5CIsBTYUN4KULen3cttELlp529RRWt3CyXXfpQgYhLCPxv/RxHTGJVN
MUS53gYLuAlC9Gz76yTmR42EcRrWRHcMWPV7G5eyEzA9QDa+u/x0zH04IxfvnvP3zUyOBF+MpED3
WfMpUMJgPdie7O2iCc0ujRz8cBjhJqGBcQyLI+EsTWK4SZeu1+ibMyRUnpzSFNC1uFToeWi295+t
z1ydUrtyUlErT3TuVv8ubmpPNo0swlMn1u3QlEvhsdwRCQe35d2bgHy/sfMaQpCSkyj6dlExoczT
4/CrAuPm5S6c6TJOkjrFeRkpJn4AvCe0Gc1Wic/75g3OrzCD9CcRp9ng3D26XB5uOqaflo0z59GF
Lc1HqhTYKvOtL09YzT/fsuccaeEfc8IROIZ7r2Muwr0oaEZDMYWO4GpBmlnWdo3kFVb0QjB6sKYX
usu23JmKDBEnrI+5+LMqxRwMzc/0ha2RZX7NY7YizP4lS4jYGc/llDpxSuW2SuWU0O9+R1PhMn3m
nSLmBaYcgGxvo6FEbBcPqefO+67LqKv/iXWlflYid0Bg/M5bkwcQLNzwXrANA8QiyNjMkPDAxaCQ
ZZigZIIzPStLNKSs49T4IFoWgbRi1770n+X3F8zk9GmyJapualCpGkHx0UMv4tTsZFbAvjGNrW6V
6GMfu2RVgB+8yPPUPdqc/Mppv4nkLnOP4KEtl9DE8pa+Y85+u2R2kg7qQuEkeuzhfc0NE3ODGoGa
GoTDgmbbEYAq+BxR1c7RW4i4jVxt+cl6Dlb4yI0UiCoUrEGN3sfi6S6Mwuke2tB4wBGQH508MffL
kvKps+rXqpbx94WiRtCPGv9bX5Gy1/KUpuT9I3U21P7LBmifvAd6ywrAtrEm5lS2zzA917y8gM3t
92cFlnHJdKJEZkgyyKg4dWY0rL8r7SW5QIfqL1EzGU2JuXmBAOvBAHE4sK8bxihH57TsBWT0mVpV
qsUZKrRko8LDyfDLOZ/zTMXqr55JjcTbHf8zKtUFET2+LTKDdc7W5dUYm8TcPpO8BX0cvbUH1sPy
h37QiEu0Xzp8lxWX0SVXAcZ2dIUhgJAeHzlS94pI/rbWGH7GBsfBW4eR+drW4GyrYbbyzmkIPHbr
jAWqov7cVPHsdcO30KRhzuRmpuKBoCZZ0AORQ7nDgmBXQ9KK39yfCxGJd39q7LGq+a2Dk66KtdtY
eTSQzFoIuAwhivXZ5zqQZhIMEBzmekE+p0eXHbO+3tjfpjoAk1bTgzPWB+ugV4yHa/JWRB58zJ00
6ne/tc6dYGBVlRAChS/QXUiq6EtIDF8A7q03MBvfsdYwcj2rSo51Fp9/cyc1+FHWX7abh/Iq22Dm
aN9HmHifG/XPoqlLzX2vzXa1pCET04RBSJUMPvee38UVBP8A0K2hWytSQJQXjPQB/W9UVyGkSyG/
L3UIKc7Y0hoEsG/ZaolWqkL0k1BkvXdfwsDqUTwRg6n11wG1qcgW4vFkm7T1TwRWIkRoVfq8pE1D
YGtngvMVtx1V0pe2zvOBzxphzTNdNE5uV2sOIq7PXx92u19FAes1HvkJXFTbZcyBCylAYb6Lt3ZJ
w8OICyp4vCqscIvzTEwaRy5prntXOVIPzfAN1w3N4k0Wady8eiMUbgL4i4PNhQJFRXL6qd1q4CKg
mf7bkXiwODiA9+yr9KEI5klqSEQSoZX5urBozmi/qqnd2jsOHVBt22JKp1HQ86n+DvDszB5WODVC
TaNIQ4Tqe/y6yxb7lLK/W9+5qG6tcY8BBI8KJQQ8fs7cAYK3lUMlEdyx3ml/rFJ3xKfuQ38NTGLr
f8eM0j57wD3coWpUZYSgmkhFWaKiKJvFVOhvUKM4crfMkzcXVe06LVTkWd5BTWl+GwVDBDE1l/BQ
tfFWkDWkHIenlsVzxz7IcKJOsA/k+DgG+6Vy80JBJ8BCK/DNc5LW/WAeNY8GAwMfikoOl8X+HosD
l8t9RBO2UmMwBNaruehQ30RdpR4YLBiPQfK26v+b9lfzhp/r3NR1mwDkNyaJmvtP7IvJz6Sspfw8
64rmrD+kNAigIhpsmS/JCblpnoXF/KBsBuT7YdZQeQEF2/py+uM+Z11KbTMTCLZSt67kOsHJ8429
OrfKuVA6PMkSbzrDFVTwbkNFKM+QCPcwW9n1K6ZgI4Dg171RSmKVOGSQcqNKPbrj8ZMVlNCVPo7H
CjJGSXIcTQE/Tydjvg2jySdZYzxKFTF/G0DpMuBK1MrO+rS3M6YfixLeAoZ/dIBez6bjAZfI2ELH
uT/H9YUu6DixZWTe9R4jt3H/ztwYOhokHGUD0bTLLGlw1tNuQVwXeKt30l/1pCvymkbVrs2SGdeM
SXsjxLpP4sTQ0sTYAG3gmVwx7H5xn71N51GwicFs8cSaxW+8KBlynBJEEWsCyiLDM/d25X0Z4fKu
UuM2uIDhmpZU1nfCmwEwE4LOpO3MV3bkjP6r1QLIFfE6IwWsLluDc6LpBxN8S62xE5zsQNiXMv/3
GS+3QgIbrXi0tV6NXW6NlHDCjUUbbSX/Ysqy0va12e0k48Ylz8Ss68mkuq7aSTVw+UZa4h1q++NR
yb66/dVX4qof9y8fRpTf268EZx4i6k9nDa9ttkTcb43qPeoJ3kI7vncvwH9lqZqqSZw33QT/mY+l
y+4yBhbD1f61yQzGe2pgzcviuvK1AA3dyUXKjrR55WmgsyTbmqQ+UcXdc+IMjy/bn/mm2VTqzH0T
C5elLRm67Bz5M2day8VERy/ctiXPhHJV8L222c7miWE4y3VkjT0ub9aIXoqpo6LmW+R9LM5jgAA/
TxD5bfJe85Q9p6HRExY10jdwqJTDyqiuYEKwP5YOrit9OlQngWKFRYx1jnA7NtZC+AGRuYoHtOy9
ZkzHXWuphUYgIBRkRihHuEg7dQSjc9+Ck0GlaOj4SO+G2hcYpKiUaeMCgDvbzHJcmLUC5PPpg74V
LUopRMl1XgCVMrnlYpf/JwE9w4Sm3jWB2w6+kFUGY157A/vHh+ErKwrToJLMBYmddFyAxvBoOqKx
1pxvtUr16jZZejK5TV6qTEKm2sD4HU4ZklleqS20dgFtfbMjfp05oUghum9j2znp/WfC9H39Trqh
TCTowVDdQYmlakzJISbPf8vfcDUR56XGHMu0LF4GnNBReCzWfq3Z88FBO7uguKeLqavj/xyFUdSk
i8LQYl5/79FFVvMqpq6JxnowGpqyc+HaVxhhc6hoVuVJXriRcd0dOOcsFVacCD/LStQf5NxkCzCT
at/QyNg2qAoipVFndEuySoGCw33Z4KvpnsNOZR4SOoCXeN/DTIY/qJgP5zetb/UroQFRzTRN0I32
HFQ+CvlzWwh96aBY53Vzktm3ZGjhmjd0TGo3IxNOecxbaI+OyZgR9650OxpW4GT+kOT21DQk17vc
WcJ+rDw4VzzONPxFs4nn/SrjibfP5kMa0W95jUc1tW+5tZz05lJTJjlVnoHGqUGR4kV8bmRJx2PA
FyU1DZlSVwYEP65t7weXPhOcPPtXp90W/SDgaY+IxnKhEGUiOTnwIonvwYEYIqqD2xFh5RnxTpPa
8NL7sfZWfjdVjO1/1EbfK6U2MHsd9YYDKeBUNrFd8su7Yl2iK4IAjEHZ0AfKtNPrESHcCxoW2MCh
AppJ91NQ5HYLK/XufW6/T+v6uKd8JZxXZ1BRSKasaDXlKSY8TX+O2f6Mq7M3WglhEgIY5LkmHxIW
r86jNaTacTHzA9a52sPEhLNGMQuxaNAFyhTH+BZY02ht9/pPplHxoYMi/fKzHlg8xgGzyhPKNVix
0vAfQJ+HRs6R9mVxUXh2ALTYdO/3Ral9WHUq6hx0TjLpL9cCSQdMAT7k1tFRP7VaSpaxrvh6JYMT
vcur/YbbnxLc5Bg65GYLuM+EA/3zOM4VqsK+VIk82O5lOQXrag5mSVW/A383Srp498blrXb3DkIV
8hnskbu2WCiTnmim1jJagX4b3ThVt5CKR3hEr27qWhgcTZW27P3etsLDM224tkzEeFwUFtvkXKzA
3g4l3SAdNbQi/mdI/ZgckVK3QzE9kIDTBo9LNlSUL/3ihVLUyhnGGmER0tAbG7f0gFs3ZmsSYB14
s8HwgIFVdgrzpIoTzTFIfkBFfDZQISmwaY3I0FJccT2Max78zQ04HswtiKF+S4ATOJzrxtF26EFo
zSGrPqAMSalIPJ9CbxdAIqkPmP/5FOQZxb9xFICuiiXbtx6+VLpcRlRq2QZ+hnYxBbhLqho6Zv6A
dqfvd0oP7qn9zDWLFVyUkJhtz5U7u7ikSsukCgHlW+19VnHV0mAdPJNJPeockjOwKKTcD33blZhB
+mIVn9IpuqNvHJspre2teLpwBL+ORjdGgVVZMNkGflRwl+sK8urQwPZd/Z6YePekHfLym0J8XcSY
YAJuHVZIBXn7Np5rJbrpxohy7HAWdF+eFUDIcGqkXVt7FBXTHKje/O17HKYeH6eeFkdyHTOectq7
z84oa50AjgRESe+S9k1ewzb1w+FoMow59K5s+APqzfj2YfGplkqBEe8mt4C+f/t2+aHZNapmJc9Z
eiqUN/UywrCm1PQqwHl7JVivslDv4yu8oYppK51Rf+gLTHMwQRMI/OKOwMJlUXU6a0PS58C/aYKw
NUHzJwtppiiPGaqtFMWz5wJgPYpdy8wuH81FzBKav2waKfOmw6QvGM0E0guP07+8WBNFiHp0ZW0r
A141K1IutHirv3P+sFfrjIusdrlB0OD4dIstOlwBE3yhHrJUHdGjXHS3LcVG/yD1AjifilcQADsB
p9hTyMiUrNwqhNBbSYV58xaQR6K/iS2IVpMB5ol/lyyFo7bwQFalmbXdnER9SJziJ0XASkogaKww
QU5BAuVgIS2gDvnqJMWR/BYfmvPMEnmZaOgjl7ijdzEjyD2Iu4xLJp7PXfjUTGZaTQkRHDaqBEpH
VUeNZIkVr6qv1MmpQ1sIip32Qw0dtFNBfPbj3kiz5c/Rh+ibMj903PlALSIhyXuzlg8DS8G+q6CQ
wsSyP9OTGV/ylUOmT45P21kYr7QdmzxBdQiIYTs5gSmbWZLEGz63H9ERq4l3TuUWeisaNUKJqFtI
bh1tZ8myUEubDaNv8pZD8z78VVRYBJZ3MhdGIGrbXslvFKQ6Ub7qGKAqjMKhfc+ECdwX2ggQiIbX
TQMuz5gJvdELtaBcDen9B83w3FGbqIcs/09dKIYd5QiWIwmLoSc0NOk3hexNgph4QmOJyeyYz9us
bcmbbZVgv7iH7v7NgC9dPrspcDd6GK3r/Om2TX9JQtRZjEfpG3/vD1GWCg2l9Kf4u2dUSnKW9ZjJ
F2lxj7RwCK0Jzf1ussfgq+9Bn/SkceD1xOSm6N/Zv4dhxilTKqgCDATcI6Hob7fEXt66+itacRNY
YL2izqoxcdrT5RDfKJ+wFCjeDEi8/25Ph2ZgfLt9RHY85UVI0BQr8ZKVebDmmMUoDIXwyu0tIdMf
oKomA3sd5OHdR9FvR7ncJ9gZ7j1FMBRrBScoMTnXXYUfgqrLSyJ5Ah4R7r5pst/j7fA4Y3omIRxa
ZzCy8GHu517zDw2HxGqp8DBrpEuvrDWGv0eqKW29WZQuTAR5PNrMkH4m0uwPAtfTA9dRO0TjT59V
HTU9HMK/A6hL1TkhRCvndLJl7BVKl8yNsON3ScfyG6kitlbGIBes2YwqEA6ILlTMf7bmPb1ND5JD
LVOaP32KltsMVeBU5BpFBj7NZ0J911cx4EwmCDNae7vkZjmjROF6YK2ExZW/cuuRXV0kwuocKWH7
z++GotBs95MHpIVMRMdCQsoo50ofFX+J8nMa3IgPS2zRtLM6t5/H73MgyBHK2wKbKyq2cQ5oPFgT
uGKfPYQ8Dmh0xRI1qHfIDI3Nydf1Ykx4trrN7U6uuOHRXoWzJGsJQTgVe0dc1XgHJct4gv5e+FIr
u4FpYXVP+THpdmvekWRC81Jz0my97XE+g6M3tG+sa6QTC4gAPXKpgXpYNiBzDYLpJyUzdXhO2MEB
3dyTnM4eM/EeHBQ5AQYMu6AjKBynDpiCge/htedGsE+cIbCDpW+38Cuxe6ZrE03MPKAdZnYBfrgs
jDfvRbN1BRUIz08zojo5eia2aFMYjZ/RB3jqD/XOp0d8uAXVUXK0c/33nL0EzJ/UN1JaP2KyO1pQ
w/lW2xTupS/D6G/l5DufXR1a+Avlhq8eI+/vh4xv5E5vBVcGnqcc2iYa6M5aPrIRY3zlO+LnY1KQ
Qy69eigtuAg5En7qK0HNeHNGUu6YPPC6j7sUgNwzRxuz9148Jqx6Nta4aWN5YeY2FLh7778QGuSi
ZIVpp3ckrUZsqRHMcl0GE17ZShH4majL4IQEfRadnjeUUm6lLzp17nhskac2hJu7AwjqzQSbcfCE
3L+C/WuIS2qNl+E0OSz47a/uoCuKkhCUqI9QX1qVpId9r3oL9Up/4sJniTIE+hva/Z6iQWV6wLsU
lyrd76JjjCehn9Nzy5X+osS7TaQfO/USQP+zp0Iv5WCk8eoOzf5f01A804Lwr9B5JlTqeLCtKVyo
NmXNSI9SIYGhfa5pREp2HQvIeLcVowedmHw3Qp9rCntjOW1427S2wuZ+NlKqXKynATXKukVnDoRC
gdpaEQrwxuierc0pXaYwTIMBru78Ipqar4H55/AmAyxM4Uo/+4vSleHqaoiZr534bxV+NrralUWR
m8zxT3iNbht6xgpkvw9ME7OfhsvtINrrhYuRIASLf6qZ85SX2Bd4pqOcpeGJFtd19Bf8Tzb36wzt
4jfKn4BNWUG1uW59aJetcc6S+a+MiLt2e++S2GbkRm4DpGkoQyVweHrBbwwSAQkMhKTmXkTdyBWW
EcfIDnpHIG42uwar+qp6Z6ccvNze8tKuyCuA+bR8R099lSTMFwY9pwHWri7+zJ5EMxuIOWlDk49y
RoyJgpmPoJnXtYfQJFv4suItV5oF7xKQ7jCZjSNVKgDFPfGdOreIgSQN4E3ChyNDy6c7Nea68rhX
kJoZxZMY0mzoGsZ8LBS2bwpnZOrUUHHiK8H+gH5Lbvub0J8OW1FVX1ESwX7hXZdLUg3TweX9Mu2V
goBDAp35Ewc3q92tOSWfB7nE+aHN/Tm4FLJwFboyEeFBduyBJbMtPwkh1azcKTI3zECi/cu81ubM
nuYBRKY1oCy+aIJggmj75cL8cyKJ/cRrO5zQ/ouOLByebRhchFEEj4H6xi7879cCtWvXRz98jDjC
8zkeE2knGoaOKKU/xBKI/UhQVyihDx27Ir3dNUHBvRPhAJdMnFJzmhcmDuj6dRAzjALxis4UIUci
4kfP3NBQNzMm+dN5rtuqxIYHb/vBETmq1j9+Kz9ID+6k+7ayt/ys2tNANVg+k88P5XFbt+IiPOP3
Cgkc33qQZW7UtXnmN4y1aJVsevAB2xw8pPaBaee0fSdXHNhnriMj28HlLm7j3D3AI4TYCeqKm+IT
QQnpl1hY2bFl9TJBZqa+uTAgmkWMuogM1C83ttTfQ/UMHwLyvVG836bWwCW9VOrNprie04aJGBi5
wo94+BX8dNS3lOjllS3WInmtN2wTeWhW22JRqNj5EPx4iYHIJKaVDg3aH/1wHMiI9ng3lH3unreR
oQY2VI21+NAsaeMGTXEz/nOZw4fATiKLm5rei6oKv3NVsWQofzFE+MF+YeHUA8/TjExwOKF0A+rS
dBPmz5sOXx4BOfYTlhMkLXz1S2DddasPongA7j+cg3zoNGADEelxjqUy2nzEje/hSrdEeUrKaq9U
eHoi6NLj1BEcJGrINO+yfERc3stVVtDz+ctu38GuNxczmTMFi9vhgwov22PlO97q1EbaJ1KlqOj6
fOFqmNs5opoT26C6HiP9zhc3OeZUgOH/wTnNJLMqwtfYY4pbLVjXLyLIVIXRFJe6Diahi24PG4f7
rd4qzY0emCZ6fe/uy4dLjgBZzw6Cy80osyxk+4qcgfsGWrUVWIwjDHhN/7zM3PYi51t97473MMa4
kdu7XpoZ/c8YrZOaaYnBQLNpfn71p4RvvjSWVp6lSt0Znr5aYzk8WTBcE8fImfS51SE3HKJBBanE
gIDEjWnkFRVibAs5zC898tawd9tGluZtGF+osznwoObgTQyWOJm9gBIfpk40KioSdlWv9EOP7FOc
6EHNezVHZWbyXh836v3CbcMa7IOF/gnr3Ji6N/w+8KPsPHoF05wVb8nF92QVSXZTsbk+p/tNFXoU
QaHqsGBlrAmO8wh6po2Vyhai3jwbMhEzht1wshYFwZ19o8mJhHeu3L55ZveiGa0iB9O9AeYxayF8
xTVSHxPtbXBZjJ6GVeEvi2FoGmGRFvtnVU6FAzWoMatxsgnTUsyKPtpPBWDphQ93bvdRcoOXLQgk
MRqs00mc16MyuOlURZ+UDqV6FcZXBf9SDJDb+W/aeWw7EI1JjUVxMomdGtzJwBFCTVlmg21sTkv4
zcdzmgT2IQuG8vuHBD58XhI65KtwSdKa6YqdcmjbZ4XrxWHwfIvoQA2syjRpj0+R0Kr9b5tzZdRG
fppRb4YkXNt3Izes+/1V63mCmD40NASkrjJN/mcgkLydhkguy3YSfAcN1t0FJs8LKXw0bwohXPbz
gzRdThfWoF3WrWkIWn0jY84v3JQJKoRvsByM7JSBuAeo21Z1l/xgJhY/b6chS0bXCudVd/qOScnQ
1HhNf5CTIGrXHfnTEnAeaaaUsPcZ3UxhJnx0YZ3sT2mgsKu8h7VyTRb/lNg9nD71zvKLm2VGTzl1
zLMsfRFlmmogaHuU9NgyosGFxI4nlUFDwinyjLIo4smA2EEwU9bL9s3Qi+lEDF+qnpchNtbTK8oU
I0SPwOyYMUAV3S5g+pAoeW0C/KGTySC61r+Atz7FOMx/4OILtoDQ8qOJlXTftZGeqjqljUyAGIbr
cMSqT+1B9jE7tLbDRqYsibW2PzddEzzuSVbxGn0JCNXggDKcPwQikKAfEyQWNR8ZEwAdonoynB/U
nPM5l3HSdKtx3947ExPBtJt0a7Ac4cX+Wuk+Lpa5KtCpBW7h8pPT1RLP0CIKOZGteGpgF9DFLPAQ
b3txC0SsEizONXle6GKx+u5XWog3DwS97Yn19Vfe57jdgQBAe5bcMsoJhlvBA1lpeNI+/CLpvbx9
a/xAgctbcQtS7YoYTzdn3cEqhDv1igbxsH+TptZ/yv3vTNF79NXlv8VMPSKCB6YX9nLS1ksWlcKm
Ins2lht/7BBp2G47D4y3qGCW3xliVNWsZD1OP51M+Y8AygbJj8BHPTqJ2RBIPOg1ti+v826f+Mm0
uV8+ov1i+4UUxMJyqxP304d8mo+jRScN3g47DE/6OxfQBAgbcv8pE4ZxhSuFhDy118SKFRd3qTuw
zWszsWYkexGV6Uuz5iWa0Usgd4SALL8sr4erEbjDQnZ9iaUyMsDbViF7uSXqzTwLhmHvsB+nZMgr
+i1lyvFNtKZ4puVpyvSPE5M63jtul3dpKGIhAmIji0yD02d1fwnCZBLv0XG1XelRjz74i26K8PSt
VsJzuo8GMGpEhLCXnEkMLB/r0imVugLTDZVsV/M+hbdqQurU5uhiNlOM2FbwU70qx34V/11/N5ax
8zmuJgdDaaPqV9ocwy/NGdU862caLayGzc6M3VpqvgHjI9UXqwA/mn0w7hg120FE+D8K9wnj7ZFg
LyM1qn/0nfMLW5dBNCF5wLK8uGri55401BtRSoVKuIeqizZDf+WrNkWONHRsazsi+yB0CbXiO/vM
uvdU9TSCLLNXnjEUVCXxySZBGv1ZE52W54yu+9GsgOSYX/KkZyrHZhIKwcjxRdPy/FwMLFqzdUBG
LxKff8DJ8kef6Sr3x5yewVt5PD16gzQDprwRk7A3oR0Lx4uJbqgOwP8BK7Vs1BTfNdMj6bMvqkzu
rQ6Qpb+CTS6y+LK5Ze2SgWYwz/cA3o+sw51IuNbfoypM7C95hHpt9z9lUXqdHkyTNvTgToPg9bIc
XCPh58jJQzePj0ZRjdsy2iY20Lx29XbFEHzKuB7hImqj5WJDKKfluAoM/npcOAcYRa3ghpdxMh7J
pSKvLkZE7hJR38XQZ/eZ8J8ZfoubPOFnEwkimQi9MOMM4aTeCfx0oJuK3Rgmy/JWEz0Lx5NDJmnP
BsVmyFPsgBcnvwIxbB33+WVYCe4MzLJ/eiUj4VEqARioUPgi8y4Gpeei8Gzp87PhsWBCw7hhILWz
9RYI9wUt4rhm4Obk0/xryFNw2fU8Btozx01bzrPPKFwsnx8pJUXVaa/SosblyOMR3FSrsp/lxGcZ
u0Grrl78QOulX+qb4Hsgyh3Gf6AA7xcOmsjSR4q/KHAONvFTpKaePPBAOZLa9/Lt9j1cCpv5qfMf
yzW/lnWMSmi/FfpN5+qbIBG0JA72Ja+Y+WC5vA9foTKGIuqHf6m2phv0PC8Gfzmz5bZuA34VxAXB
gV5XDPvVRkId2uZ8PDmrOYRKIi43NKQW0x9RaSs4oRa89s5RJnAx6tdF7WwtUbmvurmtHD3CUsxl
dkyAlakuvzOtPtjpBQO2q02KujZu0Clhrgs/hIJKDcPR3FLfrrzzZ7BN31dNvdexRLplnLphm8QC
RVh+q6A32tQmPlLbt0U6TiY5VGjFeStmgz72C6qs7hosN8bFSCXrl45KTUG8/x2nN0kXlR8/hZum
daUUvOYQCbg8JnNePjJKt59Ctk/c9o3UM8MAZNkknNrxBa/dIA9PZmM5uEPU1LY1veiZuTXJjfcY
jenP5OgtH3dHc+3QZHDPQBeOmkElgTAA6fKnNmfpFqLACNlSbZHYd/PTbExStI6y/6D6xHPrB3NM
vkZQtIPD+YJJX3Lt0b4hYcL0RIwKUWDhCA5am78OoaTAUuJATdB9srdf4gJOLXy5w5LjvMxhxf6N
3wpWBkypoja7ef2DU39N1dsWdB74zcRFu8ETkQjTbfZX6BZ1Pa0YYbs0kpMGIhR5FNuqiKh5ERxR
pBDCV28sn/juY2XS3H4KxzYMDU/0OGv5xYNh2lc1NHVMM4IXz2ayoaqZeUwWQOkLJiZ2+eqeXtgQ
2DsCuubEC5zGxQDmVS81KNcaIqcC4X1dTYSz0ubFH5r7FIsy+fs4UbHxwrgMzgVdAZk7qHLHELu7
yUsa1bnwcj4eGFKPaBnTuBG8zsdHGUc1H9bCz311BYgRVQNiWvcn3ewrGElr5hP8zeoPPMfMT/j2
FPHgn7rl31IM3X9ZqZ7OanAFsF5foSVub6Tj0xzpxxSC0tWW+LGLelBIBT0BruBbc/tGPxQfOQop
vciBwkEWE51aV3ZTTicSgb6Oz2yqOfy6LS+4x+cUk2iHQYElP8DONthtGKveBwrKZPY9GIHjznst
z6aV8PCdLsKTo2KgO1EX1qMzg8X//z9CaUYoZKtqsX9+pEH/DRpDUPCr8NrvNWSMNsbMkJdhQnSs
lgfGcQCL+uQy4DvO9g3YtLJqc+EaIJ5NJwJCXgQ1amoy3kOi9vZAIFKTL0fpRIMnsQjx36JXzUnm
lbspsP2uD+QMpkFAfOC5DdEcFrcNe7itsA1P/aQb0xh/4ksjnpX5vJLK2hSRdMQvex4o/K4/MOAE
YgKZ6T68TWcpReCvrU42EdLM+50PDuii6EBmUycoVFJCICCrtuN5rPWYWBfadujrdmp+ca60diEX
yjTY3svOftFwqZFWUq0rJ4pNqdWB5KErAEFYtvjI/czYQ0EynOYKxMbl+HIlomNXaHzm8bmGPZVS
yyo0bL8NTN0St8IaudTce5PGS9ASIDklEZf7CSVh4dejjeMpLhqH0SCsBwno/oJ/xzpoePiTVkA8
pu88guCLPm7bP2mk3MyevSv076pS2bzVNiidqgPcLpmI4R7xDmXSdrXhFgJ9IsIj1qSa0Z/CvkgQ
yTXrB7AhwoADMqnU9g9CVDkTWEVnprbG7DoonAsm5Qf1pZGeRHEKp+wCAHEWvOfcOzLIE8IGswp2
r0x2KuEYY4BhnfI5N9Rkm2tvJJjqtzFwSm8P2+HwQXmI6tJWuHAPRqeUHQ+W/XoxcpXobpiSmZxj
s/p63DCjXOPu2x2l7fDEtzSU0k2+Jysn2Nx/FUSn8Sdj+pAVFDHUk16hvWH941geUjW603uxxuxh
9hEEf17X3eUWLnFsENmOM7Tm1iuMQZ/yqhqJBvFm2JyYyq0jO7nMottP/x8QIrR4a/4Oqkd/tWz+
V8JniQKujs9yKur/oiGTitxmBV5rebjQjF7ZhIkpFpnX8KvNc0pitdzQoFNQfVAI68JbLe5sAo0h
uowRGYGRE1jeesTEi2ssHjIiNESIObZhLKSHBx9G9G1BVysGYoPrwkPYqGXZI435wJHPNfHEXfzf
UzPeahynT0gmDM+YAzLQvBDDIz5dqex4dikcgGOvJC2dr2Hukxl613RFTvDyQqpfoDX34MBAnwXf
vZzivHgclUv8XB6od6rYjfLBVGVqm9jcGRnKXJt1cGtqcDjcrV1Gl2UohYQXUiMpl38vWjdLCt5z
orvFJE9688jPsgXK2FTbIUcINhF86Nc4aK/wyul9VTVe8nkx461by1raM7YTEJm+j3zeHkXzxDWa
4h5KfI7LU52nvXJpHwPxNUtsFfHXGhgReVymgiJENlu8e4shZDloIwQNwFxZwim4P+C0YaJEDfGj
IO1upR9mehzUSGRSWJBiWfP4CwGaPcZsRZ+XemuMuoKuh1uQGEgYBE34kVOa5gjB91KmC7kkL0UF
da6uSrTsqD4x22OVXexY7MdTYXpvEc2uGxi5misBn1r/BYbveWVGQ5Pl8x7uaxG/O4GGvWzp3cwp
StbW5kNX/OvM2FOA9xb6P9zrkZ/QMi1M8uAVrxJcrR3TIWx0fXe7mmfgN3RBD3NLACuh7g6sod/D
rHeRBxN55n3Gr9WCoTNnZ9RsvEBLw40QaZBcAm9Mtk68+fQQIDyi+akm0qtkqV6T/g4DD38/Reus
q/6vLH3LRdHCE+Rx4hFN7sA/a0p61fXf5knCFwDNKMXEgEHLBa9y7/ghHET/qzERfJ3Dk0qvV5mZ
PLS7ugHZVvQz+6QZhqcXFecvRvToIpHsr7/3+6iCyKGNBXL4hhOimS4ZTCHWKe/m4CPy4Iu2BnJw
shhFMEGPxPVJIuU3H1bzGTjIlEPZMC3q1aSYMftmHJ2GNl4BbQvsrk4plIZtoZ7f+rGxSqnENfyf
o4+d0IgA0JZfQ4EvnFzACTJosQLfZgnr9PtONRNKufsGBP5KinsRuV2OKfvMyfhlbvgWIaFlVf+Y
iiSns1W9h8169wAIYoMpiIpo5iQEGtinNxcekSeFxkV/4hkRpLsXvV0Ez4C/4NuKfetTQBkcLpJq
uQARv4i5DT4bBCfyvX184vxixgsTm0YQIOMyfD44sg1uszc2PnB0/Y8l7p/iHu0OYN0dOdsllfu7
xYEqsCha3aELRQTRe1+EP10atX4bQmxlJH0vjiUFyxgfcN/vFZaUHXMngoF6Xv2sHCRWSymEsCLJ
1E5AM/kBoO0/Et83ccK9A02gCrzGvRKauP4UQQPZm8wiqd0NeDmuYjPGfkrB4wdxCPV+jbBGq+bn
hPKqRCwrVh6sbmq8A+Gjt97eQAntRC9lDIxCPar3zSK8baZbsSWMz+8aq4zfvlLEMLZ3Fo0h6LhZ
idP62y4wPaoQ9NYrPPgmk9yyJXKXPEBu13UmUoXKe3a7hprNsNbXNAd3MCYJmdxZSXGcxVtczd3Z
rf7rJK2u3vzfhnFNiDPHE3SCAV4MoQy/96cU0ttDbJwUxmTtDKvYmgGSTZTtzmtWnSc08y2mp9Q4
OA+mYoXY2LxkROa47PtaPusZaQ38F7PWp4HO6LKfiS4m8BquRZWPghFKW0/eo+8PtVe3OayKYXDr
/t+8w7qApj+p+FjsC8By8V0lq6zr0GyH1TDoZf2cSlDKOOVwYIRi8sJ9HDIJmH9Zhvc9ZipJX8RE
9VFUXGiivQnWY5c4arOduQGnrHdNFUKJdSpvWHwr2kbvX1wX5YEIFcN8H/6aV710aZ53OgjLRO0g
oY60lBjWgOLLORXmcnPAwWet/gic4T/saUoKVkMlij/ID+rxnOgQCQaCaZU/oqoO+ev9KJnIijFA
6BDBIoYJTdT5uwbA89J5cqX2zNLfzsZiN2xMLtolTNEj5Ov63SAiteJGJTpFH74dsijkVAw04I81
MpJ0AW6PQKD+62Djp/184h6Xh34ak4rjlK+FNDrqUGYsXuBAEOMU95+jEy83UF0Ntgztm+W6tV4F
oz+3JhpC8QSDb3Nro1NJNrX5MCFTBhElDGif38C+YXxY9whPdZFY043psLoRWeOtwJt+jinuojou
n67IB2kdV/Cj4MhWvjqws3MuOmkm6snkEw3uyK2GdvhN6qtesf3Oqnca3sXJdV+uh4PqaHFLNVu4
RVd72bwJyeLx4IG8y0YKlfYTfMAtY2OaVqwNOTccbWeymXEXVhpdFT+ulQvJp+N5tQzfjO14OTRF
tyLC9xpoLx331Z+UNBTxPu5kwqiUOqWbBpUgXPinsKhZeN8afrpLC0sFIPYQLbhN2I8/MsU1H/my
kN51fj7Ge5HkogCzecKr+97R4vu1bT/HGfdHur0jyzt9TEY5GjtsQCfP8VT9LihcPH6U8w8wQmt8
amjyJI+3jyjgsgoyQijEeDMjXlY+0+smF7zsQxTW2+JHVXiJ2EDv/AdoPwEbn0doGcqGa7w52W71
k0HTB6/zVu2qC8TNBcS9IwL30MXaIZLICXY4jvo+7j97zRxEdBht+CYjLafwOTDu95tmvg4uo/MS
4DgAGnrBBvqK3uaVqpHOZNIT+VO+Nv+SgdLcCVJx+FxhZxJH4NbJUFCZjCP5hSiZObLaLuaMYizL
C+NGtQ5s760hBDyVczRlAejAJIoFuJx7PkcR25oECW1XCIx6CwdZrdoz0RUAw0klvmta0Fz36Ig0
NJjC1qa9KMnHLNbm3pYOy26Y8ZMrItww+gfcKqLzdcVwFbKSCEddMVoElyBtFo82cPxd27/K76fP
p3aVwDhQD0GU2323a8w9ykAvuy9rR2nM9IjY91iAUT/nSANv1dgZmm5kdR97F9RQz57FEtlFhjcT
lnlhCd8eYb2PstTiyTzRu6HRtX+LE0w1rjnOZ8LkNlapowFtXoNaVRtJRkZAENZUKI/GmWr33wNK
A+auAq8Bql0FD4OZ0eIxr2BW6+i6+vrG4qX/2CEOaXn0JXcFH4Ds308J8i5b5hywfKNrNGRyJ0uJ
SNtEJN+k66OHW/YO9UIM3HV+zMVe83OZxc3e0vtKC0wNfICsjn8d70mk6JNMM0uICYfZrvet/Q3C
y0usSB2wcxOBp75F+/oMR7BAN2lMTq2Yd1RKC5XC6+KfYxRTqWKRSra1ZSYdpt2RZo8WR09ScGZ6
56rK3H4Q3W6bHL4JfpK0NueaPZlOkIDE6DpWxamkxyLq5My05Z3RNQuBY/EpAls5/eU42MwG7z4z
1v6Lp7dqjoRqms+RFyG4p18PZDIehYFhjhN00Q5jMsd8uUcSfpt1SGe5QUtebY5OS5kZ6wadF5u/
5s0c2xbUnT2eCWu1zVjbLpWWfbndyT91Vi/5WXKDhXTxANmd/w5gYkxrNkiP2I2NprYs7AtdfOPo
hlk7aqbkHWsQH/mZnqzpit0P7G37jz1UEbOlMNRKIGYZiSVBLXz3bPj007zKDeml59AsMKrlj8f6
JszcM2enA9q7Jc7SVI+hZrgypzgrmmO+P4Q8SdUPbkUfaPPjQjyJMxnzqqsYazoUpU909k0/AveO
7ofD9nLZ7001+b+nQsiVu8LFHrpTQc8RlJpcbSFI2158a3clVjRJ+UdRQqz+5Zt2SWbBatTHCKEv
15rSz7hQ+nybr1X/R4PYYa8AFYuDQa0ymoid43qYa5oANBfZwkS6MNDGtoiz+cO0J+jGGtFTyyWe
WhXbZZGD4k7URhvVVHbDS1toVAR0YV30aNRk7jw3mmYaArQIU25mZpfYDnZJ1ZnTi7wseTHDOZpJ
I0VCodXxu6OjpzlkvKQRyqvbM/bPOdxfu/fPvYZPw7vzryw+FSzC5meypG+ofBk9rkIOnwnPNjaU
xp7u2x+Z5cfNdF7O/oMup3ZHWjyCcO1wt2w7iJGfmku9CQbOF7Gd1h7cmgJBNCfFmWnr1rw1LZrX
Ny/je++OOF2qMYkoxDLjzkU8VDaptmF7/mHOVJ0pmywGy77ED6esZ36wPimrRE3HYFo7k6A7RCZQ
yeuwRZQAFlhdoCR5tAmN1zx6gzuEzlOWo0hObg0o2fpM70y93ub9xmO9eQaey0G/2VmwiZwnlS1B
AVyn3TffJilTrmezQzjgmJNaJqGGLUiapKHOhcaEpACHNGdA3DM3eRBdpTOEvFdUW0FiPo5LaVIW
GbbTlbYnT6qWLLGYAezCpKSHn4h+KJ2CQA1eG9d/ZRaiQfQKbiNmWMM7ERBGHRPAVjHyOiuJRjPA
fzG1eyfsTUDI4FWUAPxK2C3Kq2H/OOrEXdud1yWJaIQ6Si1kVvRTpClEvswEQO4prLlCIZt84HaD
HbQpnSNFu9JlkSCzJC1o9Q7e/zI6DYuqtA7kuKMwbq2R4qmDsky73uPoErUxQZGA9hOAlQC16VXt
BjOCHB6CwoYyL7zdYKSqre+bS/TDCyZdSgFb0wvTMlnRTq6ZxuiZnYVX2KLB4aITD3JY19rQu/qh
ahDp9813j6UEML4kn1J2kza/TjJP1dgVrQWVsPM6QPRFkb7C7kyIonsKyA7EeZ2GhdkvB0GnpOiF
lBkG3IYjfRjvv6FgvjOjk100jAeH86GogOvaV2vUeoMFtWmmMdEaqsxcOYmo2Q5a+ZXl5EdvAy+p
TXK22Z2y5bXr+YG+/qzrQigjyiOALRJGPkU0nr0T+lKC2JVXKe1MCcFxhqg1isNDMQAl+eSypdwJ
gci+a55K4hzcF3toRC4RHBY8A/xzx9zwfxA4sWY8wtq6y9JvcySR3GrtZkeDgLiRyfhAjBVac3Ub
uHyybCGXdlRD9k3oPFetbnAQzIq0uhVbtvgQuVbjhsVEaYT1HHUw6B+gWtGuFV1dvHxfxH8SNt/e
Woaj04VulVhX4kyafW3qyvE9zD878sfO8huAHY3tmAgIEAJWh9ZWKs5nhfTOirDQeuWempgr2ryD
mA5qjfDXxXhAOUKe3wxvHPZISlrrAOfFuCxRIHbRepVrR+43hVmfsjd4wO2lO0YWyKgiOzSGX2hQ
S7ikQsq2rgBJpr+CZ1mq0FfdUPgEw1e5H77WRRVNkfzacUUMYBE1LBVct7fkwPxjlEFAlUzA6JQW
GwGUBAGnI2jOGCLfFPbrMO636SnsNOPzP91y1GbKV/qcDXBxdIqDTDPVfq9hUACtScR7eOHqAR/X
T3p0hSelC0KP5+j+fCYCMD5XnmGuAemHinJlGy4g1PlfishnBC1IEmnIdJUZgsZlOo6F9gGlt1a6
IT9jcHdOKtHrZ4hKdyBosg15+lHvJr/Ftci0G1OnHvyAbb0GGpgTJr2Or+BxByUyulxNktGx0Xa9
P3BSYApkCrJmKn7MvVsS1bnRbFKTOQeP+HZSZ2WozDRtfMHxPqCTyeUXJbW91WK7+T2vA7chQF1U
SGcO6ab71qv/Fw28xdbbepdSm6lko5A4XUHgqlwoiwZr8ZJ2QN9aiE3S7jg8y73Hg0bG51auRNaK
4HJw6taXxotPud1wYHEXnL5sKTRse1WFFrMOt7IO4NcbOx0CyNQ2Mfpor0XWL4a/tznwlfz5KSd+
S0/LZIAetzUwQUEGJbJ5LiXrQEgbPiTKmr5yK2F08EoSkcQykzI3RvTBiIHxQAKHHf7mf4tyC+xa
Vl4V83J6eu2Bg01q40yw2nIdcRaIRQ0yxydh6p/A2oABl+5xFqZ3y6ZD3l3AL4mToy2ONheV2uIQ
EaoRNGLISXQ256e7PiRm6+Dm7kYS1Jd3MMOh/IgZespFVC9eOZsVdaFIe3iiLXyAh1SrftrEv06n
dihezVKIw/VVr6plEL4A4EAi8I04DIqdHA12LNYivoTSSwKDdpjzvvEPfgFG6FvLnID+gD2Awzn+
bJbB+lF1a4XPWBlKEBQl8XKo9wsAwE4kLBQeRn9nbKGKDeZvGiNdA4bbvsWKOzIv7wjoiIvidNBH
qSsJO5TaLHUscXl82sepuPpc9mcgnz7WYrFAtuRRCNMJGE/OQhi4QiM/WneW6AHb+KkPy6h5yQK3
XZZ0i3RqtQBl4MJD8JLJv9hIrC6osfS9+PjEoPWZhGTJckUjeXeEm2dR4MIpcGEJ2tTkMPu7PUMJ
51/oTQEEboNlAQe+OzVDg3N2vno0hxTfSdspVyHebioY97WSp40verZ4h4MC3XEpdDvJgQDhFyJt
AhrfDVNUdQxcLsXfuRW3o0brVvDdwTpKtRLvuEYMV96lWJJw7BFzRl9F4pzB5tNFYcB29HkG2pgy
dm5uzklejNJGukvQNyVsTZlIppyzIPMXwpVrU+hhlSSxbn/KgEHOA6jd6roRMT2A3Z5H1VfGLz1D
WAZqGzryucCKNgKsG2cTL2yfE3g4Fr1a9+2fGNw1cEsqJM84f6ZgaTT5p0iS12zBw7R+5gsMvAIE
rqQHObRG/Wj6RIPFZZBFLeuIIh2qFqstgjj4HrkKh2UA6vcsc+aQUsv20ndcnu6gfkO9wjZwm6Qz
EzUxYLtSs17SLGCL2/RSZ5b++a4XdNVy78dNWhlV+0HKiuedMGT0c1evvmZH8eNjI+S3JyOTG4Td
wIYVY8Xnvq80VIxBaNgnMySSUpFPh34ECnglO1O/AhU4/wsRzYCOIaXQ4SFF/gp/0O7Ev61q7jnk
VeEB1xd9PxkVF0n8x2NaW67zQiyLjJB3nRNwgLBgJu/yUk/EaeEZbrgA9J9Cw+WhEGUrtZDksaSY
1WWMLQsMHrF8R3JIFhYEgoJxKLxg+9kF737+tFyBYxay86OlNY0/sDEfMxr3QEI7H7tkw9vzPICL
97BV/NBjxW/inOkoaTUTaX5B+PRqrpjeQe2NLcpwppERqUAreho9qQWRRPFYvkTaKYbA87VWwyj7
6UYjCUvnkfpM9/ybFPMkPNETeOX9dsKktXZaBwWYTbm3mWJbFQlhu5NfnTlrwzzrdOIpxjrSDyUF
umHBES7n1UDDsrZ4RJY5fZujHD/m4j9o1Nvkqwx4aK/sQmh6PqZ3V20kzZhAIXXIdUyoBH68COCo
ej6h2Vk5xEMQnTAoWKd3H4c0QagmDmYjWWcohbIuhbarBPgIyIu53oivUVfCxKROJ/bkUH7EUgMi
aRU8TiARX4Bzw4FcYeOFgfwqKduG0W+ajdDwdjIbI/msGtp3rGJ2RkCg2BQcmHc5TDOznzJGmgOu
ZDxyFqX/cxew+LQo2+cGkZ8QOu3WTqWTtbrEfvpB5B9C5LnxkcBnsFMvJIp8rzPm1qbXhjYkHBlH
RRMdGlBFd+hr1G+Qz0gojDw76ZS/EcvGBr4gaQuBK24BWDDjlsZGnx15H42eCJ4FWoxCP6P58Lnp
YwoLhGJTK+gl8f5xyzUbk58/IoStGbMJYl//DyIRgv0dU0wgfCraDwGHvUxu6ykDptaCvljJAgV5
Xm0ibJ0j7fG4XeHDBU6zco574sjfEAFL+w6sw7tEJoCdkMQ+FfI+FduuH+ctSkPlZ5psIvDJPIcY
yvo0sGkUzvrxz6hYHFtTJIvtnwzMQgqumaj9NJzfutol3YckknupT0p/SVB4uvHc0RvccrJfoM9N
2soDe8wnZoxCV8qJewNeZtC4rzJsAMO9aADVm/oDh3ZEoaf3omYan8LXac80RXO0Xj0e+zjx5apo
8uydx5HdX6zKHAHFE8my2PnoZAqsxIoXgrEgp9zSp8uAddGclAo+XOUfpWAK2bZhdpc3kNLHRnwd
Yi+1DY4XgnpnrvhFXn/gxt93jzJclaINnukMdfLfg3gxQxky802lFrutzJTlhZ2Ueeal30fP5Pu1
t6mlkKxZkuZrQgt4eZNxmIk7hTOstbkP7gChbhhteuxVietem4euznqu6aaUAgnaeXYkZkohwxyz
T3Nox8TYrxFoB0SUCIflYXzE0Bmicg0lf0Z9jUtjzccVbrx3YiDxmtgIxlJ6lNrMNIwMjQKQHZGl
/j0htqyEzSsFxxA8BHH+w/fOUL1nyct3GMmXR02iXyZ8ojlUA2CC9aW6FgB9R+564ydGQZzzows3
hY2O/IdWdhdHGZ0rFe4sQhIO/NEPCJxlx2o3OVQSnBrqNfh5XYE1GfOOqNEDMfjT5Twq1c+TpZOu
n8AW+QkOxEun3phjb5ipyuLMrvI8inon2siMJccRBmUiSfxOghW3LjH286YV0kqh4fs7HdoCo0dk
pi23NKL993jNMXc1FlLA0lKd91vme2kRUy3I7ONfxxQ+Tn+ofyjt/yiP1GQygrLjLtKDpe6dIJYt
oODf20eNtNxR/ln1P5idsDEV6xika9QIdxFYOpL4qsrfYc1Tw4qY2QidZJt7hW3ZWZz614NJuw+w
AVV3nSeZRFS7utNH0gUIo2nqv8HJJR3jN6klSTMhvL3g+CAHr91kPy/W/aguYd3USLFmN3JQDxcV
Y57poLoibMYsf9IrAx3bw5+O1dXiDfhwLn0JsqMNwrtLKPJirc6wnc5m/DjsKM/ebjo5rZt0mmKZ
J/Bz0MfE1U1XzTmhX2QKZtpFK7EPsWK1jMATHy7g+G04o9lKLtYYbRs/+CciMlYfpWrJRGRqHMaw
bAFAmDBE/q2onX7owZaVUyHimCb6tmyeEdlxo/4m/t32Ph8GEfYkOjTBrGYOZA+AMU1DXHE8D6t/
EsEpV7MYEsRH3w2anFNqvAcLoOV8Jw/L8/wAYi4WEfv8J/SrZO+HBzyxXVBkZ+yCzG1zKLr9e+Z3
M5buuRyMepxhSHyTzyZ11eCbEvVHfvKVgQw5yHfOCaegkKcIF2F2Sg0rthKFdLPxkRbScp+CkXBf
H74xX23DEbNZG+EYpIKrRoUzQDG5ew8KSiNdGmVzjrxAcXMEGOclt4lzNxZz6prZvmsaCiO/olOp
lhq1ubuJJYP0WMji5i7OD+m8f8OsYWWEjIG+jg9uH/CfKBnis//FqAmvm10nUOaJAHa8AvNN+eSy
wWkfz/c6yYfDxWvwxJjaFI028x3cNkHnhkCayjiBim3xFPJdM7I9KvxPzme5yvucCGli3vBcKlDN
Fk4twLQUyztd5il7w8ugCswmvG5Z3y6zeZDbtAz4Thj0OqKC5DBwNedcdqM6yZ9xW3sbU2F/cwy2
pEFq5FHZaZXFd6v3wYTXb9fl9G0SSrPLExQ7JfR7mZkpddk7mcaDdT0yR3dsPRX4tb2c9eZVh7W+
d1YvC8jjGksf+yM8vJt6BEBo8PBkiQlfajMfJkRecWhF6rEccbnF143fsnRdrfOe3hIjJzWI+d3z
B6JH8yaQ37LPMuAnnH46651LKtwfNwZX6jcDCPKDFYsPPVW/M0Zamlo2U07vbpZ1rzKfWxgadGGv
/skrL0iEvtRBG+DIqoTaVbOvekKaSIqlDlHOllz7O35BuFqxid/tsvM8Yv1sf3UXMeap59YUZgwy
+97HH4F/egcPIg5sGD+VeNDZExUdOQbJwjQtr2rsZfYk2M4AD6LvrUT/tR8cRoG4wyYyABglNOc9
ndF50IxJmyHQHgbWC4hjAr6rk04GiEUoDAFryAKkWB1oVl0ma4zNjSAQsP80A3VwI/Rs/YskgBfk
tvDEvDdaH1SogqkHZkZUrikUuMVC/1IC+JczoU0uYwU7TfACbA0P1TsdrueTV8SqfxLEwnaBqLaC
V/AeRMjPhwuxEP8CtygMLGUJ7ZPG5El8EzMHGFIC/84gfRk4Nkl3PAGX8T8/2uHLngNn4g0Z+AuE
ptxLL1i8DDdasBk9s/QKiglNT0bToSv1mrcPQ9rkTSi7613N62hAwrT5XEt9jmKyohkngWKUfUr3
L0+kmF2tgLtRhzsZVoZZ9fHzk4EROVJHl8tdqNzgVbmMkDuSZgLWNy5z28a9VsHOyyNUOhomCPMu
/s8Rypg5lB2NWtpc7BNPmhsTroGZE6FQpkKc7t5hmD3eKGjCha3JL7ArFMti+w2Ma9q1q1/sZofq
f5ILbxpBNZQGbP+mwkVf4Vldljs+0vONRY7nn8f+hhhY3rrq65+KCAmGtauGI7vW9QkOkObY3k5k
NqbCW0nBGSFnXa7wwhMzLFUXgk9oEd8D9awvykUS7a+UW98ghrUh7dV7mgfYMXt3T757meIyu6Pe
rcndcdHn+sjUDUJEMx1EvNp7LjWShiRkZujS2BO9b3sCgFQOnGNVn8jx00QKKWL/xLSP1FQ8oms3
pp0v/RGIeDeuM0ZJhvhC8dwHJM1DVMBpGLNsInNPYywwONN3UDR+Rb1NCdguwXVgTWuGJ4OjQsmn
Zm1NeIdM3eZAxV9iD5AAK+/szHiRp7nQpSP5r15aWqQkXKGEvZBVecnH/q7FS4BNYUyc14prjdfi
gL8RSNYUiMZyHVZ+fbsMwqMHb8+uiu6kd5IxWDzVODvV+QUFjN5nsGGN2cQ+0cW85mG9vKy7tK59
HqFt6+dHBK1vj7oV7Zo7jswkNuV6D884qkCr12gsQkfTxM6IenLHmsYcEIeRH3IfJME1dcEa+29V
F48AgmiyFDR1lFE/LmNlcS5JjDpgevsq5s+M9Y4NmjVNMfzov1b2HOfoSpx167xUf/UXFSJAgZr9
J5SrQHlAGlHggdU0i2CRvho6q5N3WSBgq6Pvn9bWnUljqijVLGJmnuKaT1d1uE7mgJWGk+s5GdZs
q74PnCmYB4GGt+5vsSTP+FVvxair2uwmEdB1eL93EiAltaqcLuIIZFRmvz3yOwMICQGnBsRo57l9
7YXlE3VAUjroNU+x3X/O6EerIE867ClrozpMa5NmsNeSDEaWYe/DfGzKZULOJJpgs5/dKkdbD18i
8Ip8XyteZUIGcVOZoBK+kZ/fW+HVuh6bnsQr4gQv+empqkFuQRoBU1ZRDKj9Gy+CgzJXrK8xpRnN
KxYIewoyzIN7QkFYCvB71NQaM2fkdW0gdagZb8m3Ll39n3KiN17gYCpfjwLJK9UHYXPOFQM4OxAX
GNkpUJlrniEmKY+MTHQgb9aTEVvrCGGJyiPWEXsFSMPRhIFSOGVydU7k+9X1k6L629jz/PKA50NT
vBD019RvA/IgRTQoeqDVOL2n3JxF1JycPWGdiL9Dz3Wt/a2PIvQh/hmQj3Yk7neeOI7izkp4FYoh
XQdSQSHaiPyELqlXzWkTnIkovMzSn0Xu3zZYC/Un4tzKiQLbZWMXYTiCVJUt5pPyjJasa/IC2zVK
ytfKOis1ucWxwARPHLqJ4URPX4h5qksamv7msXcwNWe46hRrfwo19yEwqzJfm15fqfa1oA6wWmP+
fZMHLzYPZhNTFHDspULLwDkwkV9zBqtH+nLh/ED2bXb2fZZKTDtZCfujjJKS2hocCuVB3WuopNoj
+Y1fR6n2IzBTfZ6cvff1Oirogi6SZ0qoll+7iidR1eJ1DHq7uDI1EQs6sVkuL161oG5YJS3jtYW3
07dGOQGfRJi9XEjfr0eIbKYzj52N0LQMzcJ2+goeQU02nY4BbWsFGa05PrIBgbnnjWmbG1AiaHCy
kaKYgLMx1WuomQoVvBei93FgOkMK56ihQgDposdKnv6oyESK/v7aHr9TdL4CZC5WKDvzBS4w4njN
KYN339kjehhi31EYyNvP7dYzkfO3V4CGB6BukJKmueTUjEElt6DousTqWHwMpd+CKqAZSvazULLq
Un5euZStk3GBo51xkgEXJXGq+COhncIPCexKkG2wuEVfX/sW3fuhrkAM1J3Uj0j7b+P5nb0ZWsEB
DbKIKR+f62s+lPgZZv9JIMDga76azqjPcz3dAXMTFfpo2VR/Kqtezi94e5wkmZLBde72tk0PtE2l
elXJ5h43hDxzUd5Datj77fRtjhwPYI8FTZXqerCpJFoNocGILmggIPJazkmujqJI1DH7m+q+/zfW
QoXlFUZorDPTGx+Wr1OPVbNk2AOqndGbFPRUykyEBudHto1Z4B+b9gC/fc/fcKPuRsU/7fUbKa17
Ef1QFdIuD/eL0qxNdoeQo0B7b4jGKMc+rQBgxrWmwRGOu92nxu4F4KsFGNPGXievpni3inP3ykN0
M8Tlf+4GqmV8MREMTry1t/LxqKC+eUvc1d4643YWcXAZuZyl7TPlrnrRiia0lc/lMxY8pkgS6po6
gM9e46v3bv9dXCq8U0cvVSorPjbK7Tve76WnNss5bHHUHzMCdhKzGdPGMnv5EZRIJ2gCFrfz3awI
c1uAGosnBc7aw0i1ghgES+l0dg8Z12czMmQF/mHgsEDjno93QiUQ0+aZlPw8o4t6YlKuA0JFs4V7
g5fFhoHtA4U/B0TuF7K0OAbZOt3S0UvqL6Z9z0MS4d276v4NCJc25chZpbLvXXrnxYOnAksFz89w
yDO+bWQo0Z04KzmRnsUsoROBGP4Z1ipeyo8jqI3eV453ea4zX9GfL2eyV4PagpIbJjCGQOtQ4gGD
Hqe2JwATY6TAZetkzd4QVRHUozvE3B6r9BZBCp6Byl7yzLT4aCEOUFuDU3CwWAPBs4V4hVL6zG4W
U70PMJcru3098lbfQlC2pIsHTdQNpVsjk4T1/XuyVeijNy6qjv43YWIJxOJB48dD5uc6/ZsjUHbo
c21ArcXOlnEk+t0L+UTNfsifrivfS+jcAivkfbZVW27YPBpXw+jWuvOTO18R9uRCH5KVmDlF3Eb2
PIziEo+nrRTvRwocFih2/0R6hK3q6cwgPGLYsHOSvs1kENyuzF1sLCIHZASSalMHDZE3e3DWsz0r
YszihdP9UERSLb0w/x5DnNvlmMC+jCG884AqY/QPT1q4aYkS60XHKuRQ6C8D9rX+XXyzcjlqn7Vd
oCazCVM/ujWNvDEtsXSfCy+9gYmD5kSvpLjrnFtInmNJokXnkFTM601ec8Rl4txOO3/qTaU3y9M+
+b0FFQiCE2Jb7rBBRrn8P7Er1ZL7/L93L175bU5ieo8fwBj+YaMQC0aGSf2RoEikgW/6C09mrMjA
vBlKu64APWSOHtFzZlPb6vPJFbXYRgJp11inY0SuvMpzcgqeHe2q7EvElofJnDrhJGGML5EvXUum
9+KWpJwY89DYsR8ffxccbDYUPDx9IXkXiIZf+sQhL4BR/08BRy+ha1RUtMpQyUpU4ag9YebkU2wZ
q7cdmo1TgMfHOlIs4BvfJNDdfUMXJSwwqJPER0OjxbhcMwNpLP7+feZPhe5sACGwfVRGZPLeNRtZ
MjWlDnz2R+0KgxC1FzWI+1rGmrBJjTWXErkzJ7knhLzH1bH8p+R7I4GBzmAWU3/zGjwJ4c3JiHPY
XtRVJJbdwPHP7Qaax0ZBhkEbWKhPV7T0FETGrQoZdFWb+lIIFs8WImTS/TGodZSNzfnmwUlJ/FHA
9O/qrKQLHI3howfLmzwgvSfdP39v3d61cSwhUpxi6jk6QWhiDBrFY7ydxWXIDlnVdK8ct38kC5vD
SlA8kXYXX2pkzWrgaypZRXCD3GvrwCIKTS2xsvx/wo+kalGB9h834djB3O3q2yUBia0mcbk2TgMS
CVJrH7l6GDaj/cNuO7gcLAZ/zy2Av+sVfalD/FGZpgO7iplRAmQBxOzCR731sIRkyPiPb2VG58tW
Hwa9zFCpzC7E/YI42jhCZsd4LhSKlmiskWdPi/cci0qjkaN1bdyb+bBKy3m71SfzARbpAMiANIGv
+S13DP4T7n6zOUWA3pPrcsjvcRU5Is68xbCkRf9ju7fSRbYeQA+Hwl9qdEavxcN4LfUSeEw5OsVN
p7mSQVzP+8d1mGQRT78TvHZt2MZn6fFq7cmBsnWiT3FssyueBuENm6Ya1XaSUTcShd10eaIwugsF
8VyXigLlVC1M/+jnQ0GIhGSe0rKVBUs6kb6oFkQZSutx+R7O3wiSz4tIxrwPizeYNlmKZRDs6APj
PlLICgIGUql+HbpyeJ5AL2oYLgKvugSpt6suIa5twRfgTxhfeE3wERxZ42eWeeuQ0IzC3bdK6ZIh
YoV6cQza0+QlziflH8Yc+NN9Qw4+Zew7MNPLKRGqs2BTL9wh2J8rU9v1iBOYKIXxN/L15huZIAPm
3m5vmM35/fELZGGNCBmbDR7Q+gJYN42O//HjNueHdZe/em0XYbSHcK3NMwa2OjbXeeC1+0lmFgTV
0d84EFdzOt+jIPiyD7Lf3EuD6QYPMf/WEcZ2J0iqiQQ8IKAI8KhQ37Hj2Jr8pCz6n4xvYMwWfTN0
l0CXnWQRXk7vLM5e6pfdsEcyuyn2/uomutJHhrcBa6aJhW5ir8b+mRydigQPbfAKCRW0raHkKXjC
Jlpt5OwBOo+Nw+JYKU6fAIZJ9wchb2m16Vk0wKf9rZcAdUSyl4n18H9eT9Yn6nfV+qLCvQuJ9QcX
KqUhUNyQR/4SgtBSxs+iLka+3kG9OE5gIh4tyPmhyXRe+SDkyhvonMVFiaZyafg/qdQfN/hBLs8N
/1hdmCjRJHj3h6GGTn6/7X21szCGYm0/G27e9Mn3+98h9WDiYXSxaciFmy/tJF8ddb1hDIHNy2bg
7NiDkx3E1RG+dU+ysqAX0UsAy5OTMevcAYY8IaWfZQJaAsETHw1cOTunhbXGAQ4vCQUj2yyqKRaP
4UuBNQ6i3QYgGJMx66kJXlCGpLX59W6QqJXrXKJj1gJ9PE6AewSs8JUASLe4WSTCOPWO+AAk1V8y
BM8S8KsCEFvYADhCicziLK+UzuLnL13pUQzJ3jilaVVqc8dj3ZE4xupJYMNyM56jBzYHarSygMXN
T0Uaceky2Pw5Spo8vDh44xjLbEWbdF053JRlh6Y0nktseMrfoNo6xxFLUss6rs4GmqYLFZgdPimK
asNReqFeueY/5M/sQ+j59jdmJkQqRiUgpYIpkH50cvI2AMLzkWV7+TWNktC5CFsXGA74Hk+yXYaC
5EBW2ZGPBniW1aJaA0xumWnZF8uKIM2SN5Jw9w2GJdCQz3pRqP6vzvCRL2dU5OTRwDZZzy9dbvSF
VGNM1um/VCwKB0oMlFMJ8PeKaQZZbAEwK63aesdAbq0WMo5rI/I0nExGQU9Ce0u7tTOuNaimN5Hh
fPVeaA8upylU3+BswqO8Du+kMP/e/91X0DG7yKypWtfraee8C7feUlIkde/sYGKUFveT24QI+/us
4cJwp8nlaI5zNwVzt6vh30X1t56GZggk92RJssBIOn/vdiNPOVA2B6dV6MtoxkVW7e2hcQsSI5Kh
UWnz+ZOkQUB7P/Sy6ybFsHH8rwUK86D4qlb0Fl1qgtey1Kawn6/bbzo3wzcU/oCCVft4IVk0hRwf
uiaNbTCa39V+8i5pyoe1gXlp3TRX97HGdZ4LMceVxwBYDsOUgJ93CL4y1be6xoAyjSaSX0BKSYD/
gp/uUIEMIsrsnIEqzDI9SIhPVYgbTtw/bm/k2wPbs8c0mVINaodlb+RDXKOKkIIIf9fQC6o/oDqe
sSZcC5mmNeR8G28+ef4K0eNOGmbLGF1Tmm4Ug0DrNhE0qlWVsSLnIhaWVJ1g593wCUpzl9uAwfh/
K5eno9CGpcNKjOz9dW9bceUcfQDtwawcoKkPlfok/jypT0Ci2hdGC7LdE4olZgOnBXu7/QikstJU
tHoB7oEcZNrzTq3pyHgmcZy45fj87vr/Qj3mL0hJCKJqdUI2kiW9x2bh6vSB5cjNmIH+cMtPDjth
+jG76/gBaLxeDNh5m8zXfT9RQ1GpL2J1yBoe5rUHJLgpIRM+GZO+o2iFraXYEtOi3K1Sg3Ze/5H0
gTd5DF8gEjKYfkLIhmbv3dAKrxoW+9gXxBqvPCjd8JPe2r+bs4sDh3szDYZimwzNwvHVEvYbq51T
jYPJExhCe1BEUHmWhSqfGGGPEkjpHnURK8eunuG0jZnjyZ1evZvhPJOPhaSQ5m5lENyYxzI9Engx
EkAAzmcE+7d4Krl6kE4Jb2adKWv5lnBUqxmHTQGQBzg3Dg9Q46y6dDfYMSXBLzdvqMN1OeTj7ZXw
W1m6Ue8pkV2l2XEgF4UGuREsstx/Rxxnsqzr9nSi7sxVvG+mZt8e9dSvBWRbspCgyfM8Y3jsupTR
n3KMnlQDk9uyCAFQgmFTOMjU6TJUoNRidBlNvZ3PDOd9Hxo6ieutqz4RHS6MNQu16pRFZtqAhWtN
5z0cf1+YWtJ0Kuk1+tXq7rCJoD6mkhQrtnoxym/8HxEluYrR7h9nfxcdGR4cv+/FwsQzoklw4U3p
npBq3R5cEeQzggTPLKpI1Ei4EZyORy2yLq/R2bVkBgADew63YEEF9xSdB3geefnxVcFDZNrs1+H0
iAIf3x6Fjj6whJ30yoQ5fWEHRDwJINkR0WWG1VEt2SfbpOQZVCS/4Gri9qjMGglWBAxsab13ubJ/
8O1RT9OR6ypsq7vHKv6DIggiZ6k/Nd1DeNnjV9TWPIL+kArfyLrfepjDYSX4FAJCTbW/h/nt84VB
4qo0dHmuAJeimVO8OpJ7vNqgBiGm3MNPOfOZtBdZQdtx93U3CaKp2OiDLqdkRoCOsmtUbPhe7pmP
gLdRf126AavXCQ+W8AnASu/WLFrx8j4uUvzL5ibMiqNXYMbHn3NXgYcSA0DS05z9Pw0OSvu2DULF
hgjjTpLljebCI0miJdC5MhbM8lcxF2S7oeeQ+KcGedmEbCUifXIck6elWiPIpIdH184ktzpLAN/A
jC1A0siBhtBEWBt4xY1xgcCTdrgORIhonZeMXIfhcIkvXLTXv0fjhEN1iwJ1iGr+3SX9uaulNzfw
0PluIMQ0LRy4XMDljcbKA4aeXRP1/r3X+MyKPP3WvAvzZC/JUAbI2QfCBWoemo1vULvdSonUAB/B
xf6cEPynigPsLOA8eDOx+5kDysIWujRPx4sf5LJd+bSx+G0YcyUj/C24l1T5LpS75mUZcV66fZOK
pzM48bxcgmnfwEgBEuGHdzau7t8v66dNMDMRW06p+U7mYWJC5FbuY2bszHZ0aC56vYUWa87dh5VR
2zJSAR5nU+YW0z2eUzHhHO+/aiuMgZikpxf03eAOYqs/iX2liDfSdVAeTVOOKNdptqo9TmvDIj7+
nvY53my61KFnZ6xP7E3lOpFOKubmNhiZS9otnUfLbPTszgXKLpDPuMUVf//3AnUn0YVEEZn9yYSb
U6O9ZS3dM+3OGG/upgubBAKfoymopkzA/IHObUj8sc3L+pkSP1wTrv32E37d41lDfBcppSltOVWM
5LMq8D3BYlB0X9PvSlQvi6pA/s1R8Ft9MltqUPF4ho7OoOhgnG67xFvuqoTj15NJMo0s3vFT5cDN
EckeQe9AsY5NKBV/upaEhmX7c5gEKzTgZC9Vvp7UPmNbkRf/2TJ8vrXEvl75FzTtLO2g8W4eTgVu
RER6HRCA3s962kC75z9LjoYPd/3sItR+K8YghCiVEIYUPY3SB2kIuK8r0ZP2b7SgSAFDiqQcC9M9
QqDh8+IVfqsb/5ttx5WrwEVJCNPXmveSHhjNuXhx43apiWj6nHXUx2253Sjt/cU4QdfMse8f6P7l
Fq2O2cayKxtwvjIJ85cOD4BSdwq/0rpXDGktOxQky1R1PRJBrDCKOiFuDVf9az8kBzk2avWEMyeE
KUJpGLTKGC+RPv+QY+efpB46brLa2SoN0XN/nhay3cLM902eFSTdpjt8pDHs2A6j/rWEjS/0uNDY
OLnIBr/KRd70CQ8AsW3aGItVlyRMUbWT9sesIsjFiha1J0JTSc9/kwsP3nFFmdGJMEHwb2UHoOjX
5hjk6iYw6i2Rxvksi9cNJqLKb0utl62XhFVZ3hKABOPIWV6uFsLo/w/960zcGuQAv89xn5fgkmEh
QY2swls+a3fYvAH82L3SQ/3r4vDhu4iKPMeD3xPoN/b0u230hCQizS6VSow8cphLLwHRwm9cvDdU
9zLIISGH+0i+GKrSWdKX4iVeFvz3fUwHzX41aO0c0pIe17zd9af0ofliXsQ06+Yn7WFubj57zwpo
fN++0g+XXd6c1UqeAiBC3KEG8EJkwLupt9T8XWg2W8k3OvheDYvNzBM55x9hxaHt0MclAzU8rl3m
cSh3ij/lbyVq9xA5WUby8i8SwUwukoEYoPv7w1t0TagC/hIMHhzTuGLhJtPkZsYgwknc/yRUN5B+
wYy4qQ3ME+nwFUiDH/EFzgv7V1imFIu3YZ1EG+gpolzqJ6xUD8smRv+g386nVyVAIuLgAm5Z+tP2
nJuYju+lg+B6KhVWdGrTf5MCh3Yaf8RLTeiigfvLvAVlacjBQt7vxL+5/Z0JVUuZ3fSNFvlQ5JHm
0OYdEdw4fORsZQLwQejAzzWibbz8KY0EZpCvYoZcOGus13RFDPECUudmNyDDA4ZtVXhSdL0BbQsL
BA7D+VzuZYUztRTTjepGmh5wg5gKrTiCgYKaQxELlZYfUl/ceMWeaQ6B97Fl96JDhZu3awmZiwAu
II/WZA+hoTGrGqtYFKWy33sMRbeM51GWhIp3nDt2aN3AlAjrYC7JWRbJPgBK/FXYzYra4P3HxrgW
7oqrjCLzjv7buGRlTU6+n+F5tRfhIPWgRu64T2Tlspo5XJ1mhitlDzRCdt33dlE2jlK1zndyFS2t
Y7JxdHS5aEQf5ZC/CQ/T2kEgM6hQ0oETtCWUZ0NTZFk1MvyO5wpukDAVaPoOTAyKGkSb//yvGX+J
ZJ0LqqZ7WSqrhLNM9rEfzlSUo/cyTSf3SRymqS+fS1Hg3/yib8XrINk0M2MmYrb/Nn5skkfsWSN1
y42gtx6TZ85Qchd4G3nCiDhWoihuuoMatbXDPjSLs56ZSNI9mcyhZnFnSYoXvEpU3F/DodvGCWJn
oyLdEK+ZAP0RW7WC9yesQP41TWK+gP3z3N47NAYzZIF9yWXLEwQCK8U9H0qel+Na/lh11rSrrEsm
xOb1A1VXiMSR8DUMtZZjD8lXqFVgmDD+vkTdXDZKg9riAHfbnY8+OMKxXLfD3fcapfVHPl/QjM4Z
4Q/5funutPqR1b/asbqMzt8TF4IqE1McFFtynR6EAiiwtzHm5M4Ru7olXJt4VRhJm7n8xXO8xvnR
/kbrn5gJ2SIzFv7ZGlC1LkGLIMq41WyYYOiU5QUzCASjwZkPxVYQrRduEADghx5P7hkfSW3nX2Y2
KVk3078gVwUlglRM9q/fGXIHxRjuxHLvwZ12lD4+6tsGRBchmeMwJddO+ecMtJYpH89yJPBzkg/1
eqyKL9gBSIfl4syjGx2eBxWbBVbRyOGktAJ5Wn7rK78gtwVHIYHNjDu/xiS1utrqc3UBvJS2S7JN
OPI3Vj1suuRfgtsqTxvaiOt6tj2QUkzrqrZqf/8MBJ3TXgvn6N3CIuKInaiRhYVx5QSFsJxYyIJH
Gb+YWp1783LF7dSn8XkuJHfaAYQz4XfyjtMZi9nJvjQEi/vB0+BU7O5mLuagmG6TMayMbncaJNH0
4YyXHvsBvyI0DgmB0WseXmnzCwhPhOx3npaJCsrL1weKF5GBTI6mCKcsO6cSDaQBTFYFH3qFJVM8
16fcfrOw0rlK+YuOJZWxrDEQevX5OVsaDJ77JEH4LJZiNlsclB26a/e/ZEaN1A7QRPEcZGfbon2i
2/bmh2D7KCFX4tVrjSWx058UhFKKhAJI9mZLjjheaVUqYNFA1RlWXamQUNaGVk/RalxdcBMAyPGG
SmBVgYo+2gvfNtFtdT/wYThMT2LyILyc8ilvLOIlxJq5Z+yIuMoHrXC4nhhnHpzHGzECRUNEzeR/
l0t0vT+GDyQwroITxjy5/vWRuZKfAp97x85jF1hdieFWBd3GJzi5GfL4Z0BIv1Xa0QYZF53Aqttj
fptv0FW68Fatp1z63oaY0bjILtaVZ0MbTbwCuOvw4QtDS7POWgnFza+I6MJfI/2sdwwX05K8IkrA
92bPvGQpIRDAWsDer6TtiPQXcBKWlfvaXy+BR6PYviy5X3mL1MDZtfQ52GS+/2eeoZPKhLAeNyX6
SeAMp3fzMNGcf1ylmwkNgIdUSyS2+J/ng5dY1xQf8cmLgiNKmh7rjAWqdXoG5io2ZrijkZQVNrSk
BWRjvAXripyYI54+ScjfgdBPAgZ5J4sh+j9w1dzvvgw+0koGA5c6Ug0oyP5AKpN9EK1Z4S3qi9hM
RcRcnQk61+UehUbhAQ7hzkeEJCQvI29qb3Cy2LGKbKuE2uZH+PSrJpJbgRrl3hUOVVWI4FXlGdhd
j9vR71mNMxRbgJZtMt7xF5AX89NZRNv7D96WLwQIUljFugP61fnEyUtCHLyBoftB42mG1TWHIoWZ
ddHZS8faDk9yO1KvwdJyHKRHCxZxK2JiZOCt24V8l9d8Zg2PgSDhunr45ata/jqjV4DnUCBNknMi
hRrm5rfPIWzI4D7fK4Ak+HlKx/9/Y93fk/gKjTT39GrDWrtT3xfgk8R46eQLqFfyIn3WWvF2eJkp
PeNAvCp9Ml1noFgRD0koIslhinn0XlB4Q/QEiQseN25574sIaCO3ipu3MWS174Zyzl4GWLzzuvmn
iAFW7yttYuO5wWdmY6n0Q4t7TRMfsOkYQvwIJbph/3Npx7d21yV5AePnLB7vUnFRmC4wHxlymzye
rnFWlda3AgbAgiEW3JwpVRjbJ/J/LH2y+mgoySuHzrzYJNBWnIZan5MLUljHd/v5tH1HedkoEXR3
TvMYZgOGA0F+Rih0osgPMS32orT83MdLnVciPvcrPYOzz3IC8K192FynO0KtVezRbDg5WfGnCIZx
qJ6+n/6+X2t9ysxYDhOJV7aJtE/AaAYbf2uBpZYBUz1Y3TlrLQ7Jt9mD7ewKoJqZO7sBXA/w40aJ
e42hFFNwEullcevLAlmH5dtjyBfQizILgZu6fCY3cRJnuvkrcCjwhMEATrFL3uJgjZHolyX/IxYV
cNo/IhmSAEBI58MFKbw8yJ+towg+On2F0L3PaHacMaYfX7Mszp5C6EKFmXjBNkf4ybd6BHBNiIYT
WJQtMhCBkRo6LZrEiBCvMyV7IfFBZOJNqtuVq22HaPfqlA9RLv+DkCLFbpbrC2DQ5VprpD9fOHYh
WdaKGSIizjqpaX0su6G0Ulh/7Mz4T5syldShldwgi1HEYF9Ax1v3cBbGVMK5DpXXkiRJCzVPMbnb
b1+qE/pUQjwjexxhgKthskusoItJ6YlG5D9kt/zkTyfAlfGR6iksHmzKgl4Kdr7O0gYDDmKVd6gu
z3XZhCwoew4JCBKkZPdWAMBsSYP1VXCsw3JkdmZJRjl2wwRFhSILvaqw/J2ALMjc+lp55LnUCFZ5
zJI5AZ2dLMUtSWeMoGw0zus41Fe9nmipulwqD0KQ8Wv4UDsOJcbqIoL1MWiNVCtBuLUjHMCsYq14
tyBgEaeGCOFmJV41UPIqfyQgDn7nD7qrYaHZDhIxiOXHZJd8YA4aCU+cHuiubUF65ChfwG1BdnbD
qWvJv6CkBNOrtiMdENSVsH5twIipX62vDrX5dAvqLSKomEmnBJNwm/x91GYvoAX3KxerSrKU7fuH
N7KAplB+urTmQOQCT9UwRYl7mqRQnmwwOeYY2MbcqaxvrBLhDrlTGyu+BKiuGguCn2QljZ/AAHBR
AO7GD1AuAtF9JUS9E8Y2QVPMjqVQq/SijLr8piAatQxV8Ls2X8mZMFrwzNBUfPduYu4AGbC8oD4k
jG3nnZsP4oWDZ07kg9yfzix03YCIjmO7HmIV7iocFpNUKMIk/oPqvjN6wp2Mfx8DGolL8uPXh58Y
Aos4UVDy5/jPHoyT/Y8tKUEFDq3fyx3PYMLKGyu3UspKgxg+e5u28cS+S0YjKO01Bn5bj6NC0BSW
8a0FYDb2hAkUwp7KYVAfyo/0ksMpoS76uLUeVDxKgqarkc1RE4olS68sXHk70F2e5tGERSwKM8zq
8zFD1N/v/ntG2W3INvaP20l7qJitaQRpo9+nnIabmiSoh/ZFdc7NBXam5hOymz87bCTUnIT+XVu4
7Re3dsdAg/IhWWSyRGsGSdJ4WerspkfzMs3tzhIK3CRnlw864/HcZuGQzD6WY1DoYoBBZvdpSoXo
+aQIYHnN6vHWQChJbmW96S3YsV3zEwCnAQOyI82EmEE7WisWr96pAQ7sYXjPtBjyFqO5fN6DUFNm
310xgAsxBs48mVAijmrGTth0z8ZdK7Iz7Law7Nf1EMWBKJP6lDnSia2GOxu89OJ7mERPaJBg1EpQ
btzxTR5LvDqH2rmEi03w0uXQQsTxKFmJgu5tBdLnG6Z+6fPGL4pB3nDqoWitiq7sS/+icTrN5hy8
qYJeoKAzr2dR4LmztN4t6jVlI4HzbW81dvEK7WdllLSCQacQK+vZn2SRj9DpoauQY2GMQ5aVLweB
DDDDXIA7c0eo61wPsbBsoJjqh4/UOXZ55kSfhR2k9Dpq1POj/flqRaJomRzle2yLCBoEi6yguIPk
hrfxlh4UBNXFP95a9DAFv9Wgp4rqz65dhZLsGv0DdkW3b2yqQYKnLDPrUCz1njw7ihPjKItzB1eG
E5Xp3EhC59LVpBGnFWyYWatXGA8V2voofs4GxaV7Go2Ybt2r1SD2uqHA199CbEkv6AExlnbbC23Q
XfJCTPy6zUEMuuW8VyOlVvEJetcWaBpSRiUJl96coVUrjV95YtdaJKjeaUbFuPzxmxi4lJs9/kpN
eEjIwMmaHkJuF9JA3NZarOAoBNXo9yD5w7N2eXCP9wUyaMi+PlTCgZuq7Ukl7ZL/zLjqQ7ZKm3zu
2qDJjmYztBu8JMtkXAdUJGbTnoQXby0Zb2aEnwfti0lY9CKjcLUgiFdDFGGEwTQpsMqmMc7/lSKA
zpwqUNgmFPaEz8DCtNyoAx8LdeOS0hR0Ak4d+KyfYyYg20n43JUCy4lv7HbNog6gRVg8DSxWDHax
syLKwYSNRaInhwasISbtJhaezHK6CNummy0Pb5P0lJB81Sea9dc3dFPDjTKUpPAwdpxCTd0eb6X0
wZudcy74+/ofrEyukUVZe09vekkboPGidjmqtVMM/7XVOBJhcKpFquRQsVOm/U05ioflUyrw1VSb
YL+IGktYVjnjwxO2uiuMPcmcGuqK1TJE+0xrYzp+9Icutf8U4h3GszU+3I7EVgJ5aGvkyUFkuCUl
8wkdpchs9Pe4Vw+gSbrQpCBg+RZkX2xvhwTcQPd1BLdpL3WgWYb3E0ACt4p5KXaNjZ94q/FLvZKN
710bsMvHXY+w0S7ajCMwPNzeeMsBbBfbp1coFSeB2u8T7zOV9CwK+3guzR6vjC5kAS+vIHU5jlUb
nOG1MofRYnIq9qOKSkROxx32Ts4+XLTXLLeIXIX9v0CHPM8c/2/UVuXaN1ylQRwsemMtB+KQMImR
bk3jcYvUWVTLsqd2uis9G7uQAIOSNMNlUc9BheevRCDbT3k78XrZC0CKo4WckRMTp6RvLKU5uz5v
wACQn0DSveCm4sMnpLLsU67Jo62vmbmJeQTJt0ov1zCVRvWdZ8OjYyhO83Y3LR+EjZBNNp1JFf91
P5JGZMzIS7YImqqLoJuJ6BVWktE3BGYHgv+pnVsBx+hATDntAvMnVHFyWzjqaoKX/4srCGb0sIe1
2Sb18X5O535RKWtxZnjCChrlObNP9RAUxHfBam4l9OSFghSZvppAzFSgwozxJx+fAEwLJwy3gh9j
gv8DUJM6gAw9UTm1YI6HQI0tNxeOFfS6iA7C6rM7FcxD4ezheGZKmPK3FBxVzilPPTuP1g8sntPo
sRsi5idMpEXfJ/Sk+YDX79v0BGEIbwY+osJCDNfpWkEwoEUtQrvxtaRh2M9F8rH7IYV56uIlKg7w
TOuzdqftN80VPxriWd2TTbeGCzeZLnGSO+TjkMxZH2aw+djnguz47Fm0S0U3jfV9XvNI8V/TZp6C
oRyTe18NbVMsyDoaxqCxMtT9+eDkv970Xuithk0fwFddo59BWijTFgFiSo0lnW8ngR04ZgPJtkJW
jFKCqGMgJRxo5j7WvWXWTGeRrjFmx0TgYpoBZb9E+WvUg1uw79W9kP+/w5plP0lCjPxD58G6TP+v
3x0KiaC5iyXYVCHXftNlbvRU4goniHhuHAGse/2knBWzgCWBfszNhTxDbmGFTiKQw68PmiMo7B9t
Y9aqgxH3UqYnuJG5tpdsX70ghI1Pf1Njkyce9MQH2waN4IcJQeB/Vy5VAevbNB+8bTDJFGYOeAUt
di4h3hs4PIcpoXeMdef7bdz3i1zT7jOyUlhC33/JWd4rq22f8KLjCXruJUblkQ5Zs8dhHnA62kGt
kJTojX/0a66Fem2LX4+tvARnpxdDA4AmWFRoqS5KoV9gkAZVrshfhNzKSnoKae+U/gApN/OvQ0EB
zNhNJhMZTk94d/w0dS2hQB4+votiH9+re41w1Sbz/iYeUH+3npOA13Qltda4KjHEC5+2GwnMX5fp
kkOMM9lpZKM8SRUo1+3pZVSfKWAj+cJodf9xUQ5+xb2g4rgAdT/tJd9VPGhLQJ/NPMeKj1z0guKx
MoY2WSRl57r8+bcUR17xtYidoX2LC6kii+qPupEJ7sYSKPlbz+18vc87S8J1LPYlHQ05tRX72h2t
rHlXLT9Y1feVDm5QJpcdcbjGN9k851wx+zv5jKP1H+m8lsh8yM9+pynYnWos3s4ngVm2fq6z3A+Y
XmdBBAQPcUrLFJ95/V3ov9Qh7Y+MrCKw2NKfj+jxE5/vCbBc+n8FKznN1+fsA9jxN61KTiYjhAtl
h03PA7y6AYAh2t9YNSXj6NjOCd1kX68vIfjMbBXIXA43sLwlO7HFwb8hTSDpvfVz4lk+k+dkpZW/
dmgqwwC+IPJL8uehgVsnEeDReEEU1WVo7CelgQFzuHM8b0M0mejKMyhK36c8Fzim65zFhhKSGptN
BiXBzToSI+cpJneT68OA3D9yoqRSMMFIIR14Pds5l6mpXYbDck6x90WNxZYcVbA4Ft8PPMfWw6Bv
PVMtsVcCX01qlDJBy+PFmHEhfWOo7SJub9hgsfg7TkCfrxPewwImzuTp4dsLpn/qvyf+tUTCWdUm
muzEFvfKFemhBxRaqdh1pNjvz8/HvzVEwrbcYcZuiAqxZlaWMW4GrvE/HQqiXJSsUHMwPB6fLm/U
ipFjHKmPZAzQ/njMjk/Ci+eoOj5qrKhLw/gVgTjE+GIwCm9bz59kP2VKRFuBVWr3OmsU68LZYaQ3
3qLqbUoxx7ZP4CiZmO+24a6mY02z3r7/kviLY3NM34K+2JBcdB8ZOeMZ8elWwQp86XhKFiyVbq7P
og2Eq5roKSOosE0mTS6dDRDS91ZOyFUSHEbU1+1nMaJETwX4owNCGTSKWONkMGuRNXQeVualBdAh
FC58SOYOsoizHtDpMVq9YxJAmdrNWG4LROrYBn1pDcU3oOojoxk+6J/vb/68weBIUwrWMnfO3wYc
yO9sXMey/tzbvp33+nZCV4Qhb+OHn44Aj5EhGCwEw+46N7xRrwhbOAsdxP/YmTZWt2YXRTerGsEM
aPk3rqpS7FDJQjs+vVnlPdz7AZC9/En6WDmArx8oOepD0o4Yx6ikkc4TohT6zpN5ISOTrINyiLNP
5YkfgC+Q4c1EQo1jyZ3V2BLbJe4ZNPubYykaDjyYGnHpBkWJ9acgIOAkiXaLflvLyykVSFmRW8IM
74bTIMwKG+bN+llXbMw6Mr0Pi+GH/B9PIWOZRKOxUJ0zTvc/dxq5gJ7CWev4Jn8mFlo3te3ngb8p
KLCI5P+DXkLmdSKyF2PwIV/8kKMvt0HH2gLTXU552byvhW72shojA7SvnYAiFEQuZGkAhQNblF5n
rQM/C7fwAv6a+WStvCnLD52mIavh9zH/7uxetE6fKh+OslS6cy2D5xaevm6qf3D9VpfPyOCxplRO
kpXX63y3ozF0lcno0yyqUiuQQSa2n+e0vnuD8KdWhanL6agCZ8/jHFzWTxRFBpdpiLLD4w0kVBWt
q49OFVh7jm+11XNvjFs8qlhq4DkSwhZDjgNeJJVu955qjTSE/W4LzLthXXPTiq5R+0ZfifF/AsGX
pdFf6Dt2oBRczvpFNGg/UK7RqOPyQl14MJ9o5xXragZE6L1wMfx6fc0KlUCE4IuVdBDmDnYdlHip
WqPOLNZmXK5GCgGn/DP3gf28GUQ+O/NPPQ9Er7YiH7Vfw7z4HHeSWW7MlOsEgM+3Qo6R4lpV79hv
qwfecPYbIIY0wZFiC3k6GLs/NjY5/5Bjmu8D+UwU7/xszrlt6MoUyWHOK2E6qqaG2qTuN9/jN61U
zy6Pb5Bo5nZryP6RVeHB2GHAmQHmA6ltr8y1mGy/gFP30g5k9IQhy7b1eDvY6X1p9lKPiZsnhls0
W+PdKt2qCO0C9MnDOwGgfuW9OJ5O8Ibq2eqpJZogwZ0sd69kYaNU876kGCd2mQpZkuCzpbeUNs6h
X+Wft9PgxMz+pPgJlEw/Tw3ewbbyPPnUmv77uHK26FbNSBQmBHFIJOskfAlrhqzzQIbhQCBeKkJq
hSsrmWM5RNZJdfAKkqzxsGDLdcro4LtDksz4Z1BJuFZ9t76+EAyKOPrWaQ9f8ZW+xI7BBsqq5jPf
MYTsIvlBnNPvkKj17uU5yaYBpr76VVvme48ccB+nmOjxy+eVRezaSJ8O7yMlI74XkvP2DcnhFDQv
b/PGUAaeDus62tXj0GWV/plq6IGuOcB0sUK2tl45WHRfsWXDe6vkx97u6+xdx5tZS7elHsL2zo8M
+mx1vL6SZCv9CHPRHedkGYP/GtrnbVewFEabtbxwD29dzyU74ta9/Cz6sdeVKWklazjZhtYBdghV
PqDuUigwrDe6aoNM2RHBBy5lt6M2uTLdpaSib4ANw7YcEvGEwgJko8vbBm5/c6jCWQ8zB0ecKY5L
KVAMUuHDV9M7bIsN5yvsySG+XmfGgxpU1/1UwfnEZwUxFNqvjejKXh/HLLR4elruVCa/6fIiuixm
92oP8GOwQprvA/EgY6EkXbVX3/7iMNvWxpjDYjHUd63w7Iy/raT9S9NmTwOWxfyTx4N9wboD8anw
vw7g+bgbgG6S1u4UjYeItTkoxlofGKkHxCET0jbgY17VoWSdlZgBBjs3unsOPtmUypbslTAzTHOA
tMMw6wrvzlLK2KJ7acLEYdEvytAjlvZ0c3BpP//AkwC1cG4ikpGkcd3ycxZnilgJ8nOXi55a0ZGF
36YdVRB3k+nqq6ufbNNOIfG3WcaF9UBUGFZyrzrfSKztZR19vV0TBLbtKFglPv/pTeOhKOdRagSW
/bo1BOakfq6UeXcQFLC9z5TV0acrTt7QKl7ktlTjrAgJTPgw3b/75Uh0UXbFrpWOUWngCFoij71z
BxuvSFKdsva56AXzQlfOxKH+whTNRr5hP0yyfFsQOSCYb/ZodBsAx8lOAlAdzAgkinnmMvip+t1e
DGgVjhBab68k4/xigboyCXiiTXVX/nrY1k1ubd5Hh0KgTXmKC/vXQQyWklHkwhR5/HIStpQwU/FN
WZTDaQ2DyecHuseMiD9RCTj0pvl7hQtbvMRhq638IococsUzD+8IQZ4815RxlVbOa8Qtibg03EXN
2oXrT/7hwQsNlTtWnHaLt6frZG6qcoXsJmfsZDlKXOcH1b9OSQ3t875ON2aPsyyKNybzZwUufoJc
HM8esQk01YU83Xz4/G64+1mk1KRctmjSlrwQT/NYMDQWn5tRNGdTiyOSwlTOdyBdw02WpFuR2aiX
Uyp37KLD/ibBLmmtYsAvHyZFoF1rsCqPmu0cYkh7Kgy945iwSKKQHYjAADUrIcJ5XROQq3zN4M9M
kYx6h0ssV6h+sv8QZuQZtT5L8rVtbt2SeJnNLE5B3oGQRXmK32l+rbnGq8W7rAKgoZYn0uy93X2R
xfp/Rlilw16unfUrJi/JsrmySpdO4Xq0UXz9dn9thOOW8GaMagbvjQR/TlCBJcYisZT/ei8VwY71
KPlB61/jVnFS/Hy4RTe1wFz6rkiBelupfXJAq71uBjnz926svBSCbsria76F6p9QZ6mb6oglboMj
mhYKF/e5JT9VrN1Q3/+1bdoG+VAG9q6UlsS6QVYKkIbDxtk2YZ19uq6VcSqFIDBP9o/9gJCmPD5B
N9r06f0k3MzjoW5VVx3kBOWrLO+RJZ/Q3gBbpZ0qNfmItWHCSHtRZbFX63EF8Tw/UZRShz+p5YNR
lk8geLhMfhAPXpF+P5/I3LKqzls27WVHuu6GJ5mMkTg2JJ+TsriZg2wQx8qaObCPXtCWq4TbcwLw
IiPv3vkduWjMM2isc3rhRRMqREOMIaSAdt8Txsb4JvjjoAliW+UCg0G16bWJZvJAAnXpi06EHO4+
ILcM6iqvDS5S8ogl2OFKIFteOguLb9vhWz8RSHvi1FbTc9rrOb+epvr42vGqvwfM1+Km2chp7kJZ
bOlxXcVV5LyZLiVq4nyQ4criqvYq7/SYzi3/avKM+uD4yY4hVHIdYZKgPRsuRFGjrIvABFVH8n4b
7a2/cT2vP9lSXT8uuyI5NMad4ACtKAzRxKoxw4hKnlIF3bzmR/uBY/CVCDqOae+4VkZbNS8WWtZn
l1nqCc0D3QN+G3sUjKP3q7JMVonSynsXV4QrKQHshJU0vJQju1uWo6RQfHbfDjbn9+daLC40jrBP
Zgsf82eJ2Mmal3mKGdwegn+Zb0QZTRtQbGhc7kTIoPwTJQWk4VwuKvISunfSCOz7AMju5wSrxsrW
HhalofsSm+gICCR81uqB6y/Bs0MdY+1ePuRd6VYcAPDuG8QWHdmcpRSz8U1haJa1Hlvlp1QApu5o
BS59Vcwh6ahUZMcKpEnUyRJ4QFU1Ykw9QSDLaIhImhEPZiTa54DbZo32UENpp6sWSAGziGbdL3pR
NEC1KW+4hjcAy7+ccV8uJmvU1EM45tj7+DZhlBERvV5Nnf8MejTJMHwxg+nwTYIcJ4sMth6FaKQW
bO4E7rp1AKEa8CfdNtlvztBYQ0pAfNneYYRqWq0Nviq2lfdbcSo+m/kBpD1LkXPI8dm0cEB3NpS6
KWKEC47C5V/xHdCe9tPqpgj1Zs0hecDeq1bDClBW4+KxSvXEFZKdKcAdOejckr5hDztWPlDXuunC
bvGfy99fMBC2Ks2VSQU8bP9SxUX1qI9Xtird4DatRPEHdV8M2xuBMRuYU4ezvJZqTaJ4MI9W3zAI
UcczvQvdsbKRjBUCKSjTi8uhsZLFG4gK36rWna3oNb5zM6Sl3+o1JSacJiZ6HlTdMlehRzoDZ/7G
7l5N6L83koyxv3LsX130SkzlI9O1tsHiJETwGU6aVdLN9bGyWExALgMjOz9Q/4961J8x26gkXUvP
fOW4SGIjYfrsTdtMZAl2l0m6XIY23J7tm8pGwvBU5eucVRWp65YsMdiWQyR01dMxS+qLFiOfbTFy
yyovVOPCQSMPW0CgaS6lBUC4Lka0o3IjhCeKy7yv3kUc8rDuoBYR6EGEIks6tJS2bkJi4n8s7dVY
Lh9tKoDEjx90KNNghTFt14QG+YEowxVZcSGvrqkn1ESKd1RsSa/9rMR+0C3GLDy62fcH3SriEzmv
bGweZnYgq78NZmAuk+HKPtHIj2JKpgkufVZF1rrOm6yh17JNbQmxW/ILZ8RMn70AMeiItzzeQ5hN
rPtQN2PH+ssnjcn5QZLXUD55g9yACVrcRHvqMdb43MXD9lq2Opk5gex0bv3xhbffIbOG4TqkxXpe
vSWgc+LJYan/GCBjsiiGIe2hFFsgDqdpXUx7TPdlSORkl6jn3/w42wnAA5rodJqq9xoQXR6P7npM
ScecBVEOHIbBWkBGI3WPg+0YSc0IrPEzD8uUimRHxtAjTTRhJxeC8IJptruRZRrTWVXt4+TqBfMA
VLiP8VALajh0WUCxeiQc267/do4p+twXC4E3shIvfoO9R6gaanWLtEIT24PvjQ98UPTLaurJfGyC
YaAty/hSns7TkUITGWQN/4NvzCNwfB8Fp/9vOXGxIkw6y9LY0VM8xyS7sAfmklAr0Vm6fdc6ydaH
paetilEOLATEr9iSfsLpbNue49DNJ3zdo75+pFw7qS4J0hL02/RYasstG30QK6tj7XF/+31FNPmh
qVHyXmVGTAHoWEvPfYZ/BXesMgGCe5M1hZvTVXwtn2GmWOjz43PIFq3tH5PgLvj7w/dl52IgWCiT
g3ro/99iIPcTXQqL49RqjNZEicUm1hgVZmP9yLvLlGbGkn1V9BmdLZbQNLD8u1c0WruqktuI1mEM
LS7GWsXaw41CUhlPXrGlBVnvkZlEu1jz5jNrJAEQTq/DK56ebY6wms7wavX9HjA0qDwDxer3TK14
8i+1MT9UKVUfc7QYivBaLemWlGGl0N+jU91CMBR5PWsfTYr2SrI92H+UtY1Lq1eGI6/twMdmlfPh
+RIpz7cerQnIQTIIJT/FkH7esjD7jrJ7sGCeCiMkJFaac23/SIpuaXMG+fOd9YW9cPqL6LeWwQ4u
uSpGhMKD4EA7OVDrsu4AsaY1MNd3L8R2eio6iogAZqMpwgx8/XARwRzjR7FvI8/EpvUEvqNR2MjC
S9nqHshNfaQjPEEJz+bBUBlgxzzGPoVHIYbVoTTEUxxlfmTV4hv6peqn5mXCnf6gtkJnfq1b5Ky4
6Mzk7P3E7irFgCaf21KGUuYp/Fhu/FnvNJb9dFocgN6aCtsdSKFGJkhd6MZVQCGe+D+Jjvt1CNF4
e9DY0RP7KV43piW4XBkxrgeM0FHFTKkuWsfsCd/3KjMfAUZ3dnbSL+tc5QRbSfMPRd568H7URpH3
0vxRwSdPyodl4OCR8HWLzMOuWhzKSre/2l+pNtAAU5D2qzRwktIxN+zZYgjtWLFpi1baLcHnECwk
DZUyQdY31PB5F7AZOLc13LL+0wKakkOy97kr5JKcqCLleTefTpPVuQatqesKixHsQhjedgXw4CWs
5KLkIUhHRpDtadMrg3hZm+MxFlkMlbybIrSHn5OO/tPybSlLKU3F/SazWQzNe0UY7KbF3SP2RMrh
WEg93JiZ4Q9lV7iu/+He2IpUns7x2WYANRz+TQGuIJHGmaQ4gHDlX7MFv3nE+JhWTXFn6uzFggqA
I01phXW+450mdmP+Usv6qJzxVXWd+1y73DOAOCQJzyKi/2evhP7nvobjQKOzKCA2lUds3ec1DoNT
612QFBsugkfY8H+RMRU3sh+Hch1QM1xDZrkYHLhC7Gx7OTH7BbLDx88VHzkFF1mp9x7CrTWn8SP+
7Kx3TQ7H0Q74m9eFTNAzuV9W96wa0iekI4yhFM+/bPM5oPFxpMcmY2pPeJGprN5ifYjx6ssxPRLW
s1ZgV2UICHjp6T80jPTLE78ngaYqQSpyGj9NunE+P9c1Fl7Aq1wD8wVJggETbSkYpGGxNfbiWN1z
u1qM+VrB3vSfMCfYo0C6Yc7K7/1S6wQp/77oCR9ayVx70VjAf4jfOGR0tjV7pFE7ZnPLlmpQrifK
a9Yk/4CgxJQ7bA91ZO//dmVz4b+w2RxlquaIDA15feloSnBzo3LHCzBzHk0OzV5vUE3x8gdbOA8H
RQaTmaXdmvWyW3faDwFTHs5waHFsHXQMzbCIENap8+e9hJp+1u20Mbr0B04hRWZZPyAc6ws1q56p
zaKJ1mAWVh24s4oGpNPovzCgsAohVnB1FvK/ewbZE169++12t8imHdvx7Hxp86Y5bcBUD4wWndqa
E+BV/Lbo3fL+7CtXyemRWhSSFZeV75H8ZN4mVLf65smXZs/SzDwfPmKzI3jA7Kk9gn63lYTVHqag
sTg5G+TsWnPEFdgjrA2CWqLcSFmnXfe3bDoPIU4osoF9c4Edwu/7JzJJDGU+GC/S+Y0it1VQu/99
ihwrBkkebNIAS/HPItV0Zb5PjlfyAlKUt9hV0cNjFzvzWB9V/2MbdT7o6YG9EOWYb2TNGvaPCUeS
0irlr7PlKyIxwIhdryxscC9jKLKPYyf1k5J/hSPkwU89s4gDFXmaoJ60vkrX2m7W7IvXuGcLoESF
VTQhAe/gpCBlwTj5BLqjrob/cibehl41zmo2SUouFMrZYRNs7AGxrd/Fl8BriyjZCo9HaODsSyzh
To13Q00z+1QEO3Y5Q+LfEBUMRNl4uJIPu+EiR5hm4O2hlyWgRTzU+d0o8F/2qfP9wgEgZt4lBAzr
vbnt1I0Q6uK8Y12PM8nTFLa+eZ4p0tBlJSaoQZOr+cm86/7zfvUACAivtsEYlzTh5JCahHAZq9ya
F8N2gluJEkmop9IwEXkkjrUaCZ2/T9JyMxhMUuHRIXrNj+aF+0R9HQ3YTLDB3eHhZM0q1YQEHMl+
iXL7Mj5piVl6t8qLdC0YCP4njzCMYhyeC30GcwLrikubQRCTYk9Iu/jz1ooU9UZO1K9U9qDdFWQS
scK7jT6LaCy2eMOXHXwXoZ1AxBbPPepiGcKWyqmzAfahESEn8x/WTfBKWIGWBP6CRc8in9J/zyvJ
1RvcYwhqy5EqTroaBu5fON9EhETBL1n+OvPaZQhy6mYvD77xCjjYc9WMYu1ilcCWCSDsptcR3dvw
bMNb2JJoeY8lYq04aEpSh4Gy/1iwsYqmvrlZzxWrDDwqmxWVIyzXL84BpBcvxNlAOj7Titrtcqmi
6/DI1KkX2IMg+jKzcLGHJKoYzwO8zpoBuZosLOjvTMLC0Ad/o79BRSFcWjujbcRMbUt7zRtD4MTh
BcWVAcxgBuNyxHAReJW2f9XYcBSLqpiei2y4K7VLVmBPC9f3dDe19PzbsnefWoE/M71yCuypH5k5
Wq8wLragOO27WxkqxQFlt3wzUHnmgVlj+7bUCNJnmftetHnUCnMXwbDOh4RsOGfh5jNi8g+bkJM3
V7xDAGSzucgpYlwZPbDn/aQzGJgVIPAvE+dJZqTSdgmMdg0dFOHnzTySAPK/6lF6YwRZBzctCL1B
9Z2NwA43M3xIQTasCNBMmKsOhf7gFZuShna8h3GZuCam1aztU5HldTWi4IrXMRFYleVBPAOV7o6l
gaQ339YMQE6HTiVgOmba4pKx4eiXN8ZhzXrcJSDCfIvSJlIe9JK6qhopUQfAnMaF83mTng5SVf1Q
MAmXw/msoUEIq+zdtNolrKcpFHaesf1St6ls3XpMOskodJmr4SQNp2/unLo9iZoTqby5zeKuquEv
or02lnKXAWhHV6EpfQEeHZCyZ832Zk/h1xR9t6yG5VQO+ZO7znB/+bLwg2E50liVJgBk7l2C7mKW
zFe+biclt8SMlPWJn01GZJQOfbeVHx04xU9K+8Mv02IPuZy/OlTiejcqF1zlM51glWMGYz3F9m06
MZfh5Hgt4s/l4Zt+eixdBsBCFwEGy/XHTiR1LA0+TPEtXKc9uQ7iqo3bqkp/ic5nrjlSx9ROUTzN
EWzl+G+dv8apzlQApCtfd9nTy1y7NU1Nwq9ws89SI11idYH6Gp55cnrSTQQdZ6Wj81q3tfrBqRTl
gaz04RkQflwQBfysaxO8yAdT0Xo6nhC54E4oFUNjoWO/48VLI0BCkCzaz78uyChVzLTo5T38Cmkp
zb8CxTF1/JS9KqLLdS4XB+4vaQ1TM7fan35Wm9WqB/fRAwbghyjIF0MPhBl11DWMxHmGldp9RQpo
gOXArdpglqR8Mc71qwVyu0gzdUKM/4U1pDwOnwd0FKenRpAZOjDCVo4uIwgnV6nELrQvLjsMaUrg
5j3pdjPkPbbb8/SFwP86wERG0vniOeNrdTgX+EaHpO6N9MzLJO2wWvLPRHmJzlfOyYD0khNFe6C+
iWGoarp8NUoBhNkRlDXRoigiL0Scikb5c7qFxp/HBlBycB654doili8pzYL9gh7rzrd+Zdl3eiMa
X0RlVe/6Y8Jemm94wmpxJguq0PKQ2tJazH1vJV1XIBzk7oGz0qAxwb//qNlWn5syLumeEyv2gZyQ
LpgkV34OGoPKZdKR7HD88UH2xYzHFVOeonLqQW0R0V2s8bWu2A3ZTQ74f+tXVdcamJ3J6/SDmJ40
mPHtEj1hMhqz55rmCvEF0S8rGKTN6SwAnyQX0RIbRgjJmMXwV85ns7uvT8vfFgSol3lqYK1CerWc
PpoOsP6NB535O8nnfjAZqT6Cpp12p9vHmoGEKFrMbK3rY0jtXkIIitGAOGLCV17hy3q4FGuJEqDZ
B804ltsaH8WFoE5+vcF3y1fYSQpRUU7q2NOT15EAu++isUbQRhh0kYFcmZdCRyGbcZIbL+OIAAhA
mPoEahhU+jAB2tbg+IcX7FE5nJpMWF7047dX23dmOsUPvAUBe9WINFWnnwezsQBYtHOGXgyHxui5
nwmsUMb1fp0jSJujYJ4KaswWKjKBQvX/E47rC+JvHwkt8WTmt8iYF531mJ1sbtAA7yDrbhFqujuj
Q2dDgPhaZB7sJHnDNGE43gU5IqqBDUH8GDKOCn8aFKXUYRBpZYZJZxFLZXo7iZYWF8X2De3jk3Im
Mj2W8DmJPk08gYnG9dAu71CybgX8jY1pGf6JfOFZN83FCf07EGv97DcybE36dIfwNxoUc35FqGtI
7IdREifyczSvlOO5XMnRsdIuQVFOLKMqDlP4TjyJNYUa6IAVlv31TkVCcoIHtHc6+ncbZyCzwoNi
CA7JzTvh9aAror8KNoFxMmHuhRXExvx4ggdVC4MWGjQ7JHx92t2LmwZT8SsrfTgK3I8Q9y37F5wn
KWx4l3aTpXEVKujiXONQPySTaa4/GCDXLM6U479gkd5wF7Php/k9lck/yTx2HgrPWEKfBzS6YMVm
JpLy/WHqr4s0F+RqPBxL/vaLnfvLFMqk9Ys7p8UDLiExeI13ko3jwdvlCz8yPv0zTz982jvSGTcM
2/V3ZOFB2YbTSKlUIXdfR/Ev5I05AuxEOl9R4JBUk40ZUe2lwgHBMM/SIb3qVJrEXWMJUW9186vo
F0HPs1kRDpNvbyQM/K4WGBehAh/7Rm7adF67o/oc5Fs21B8i7ncYcSdX85/v88axhWMMiPHVCFS1
T47KiEkQhdpyVho3H2iOJ5XCYJc568P0d6Z0Z4yDy3lXkhu57Ynfmw9mIX4qBjCcKQgVHiDz5Vl8
FN/IUx2YspOhfNonhmjxxmBeN9v6wuTnGDR5l3yfamv6LOdx4BuCBTB/ns6dUuijUgTdwoNzV351
vdUGXB8on1TzvWZ7rIgPUiWYAWVvqr+cNqyK/yjjeoDC2C9Km9EX6izqboEW7hsMZpE7nfGNoNJx
YCcanOyWXcqv1EWjNqO5/AHlIspULe3kM5X/4sB/UtneBpmCRe9ZnlsCpNBDLJuB74RcsCTv1lco
xfkHyUX/GR9OyaFesgiuC2/zpdQ0wePPjrzvDH10B8LMkWPawH0HO4LhqgVagCbCAZZ0ok5R6ryW
4sxoJEv52pE7K+Gw9D7oNaWmq3bxLCVe+qpsq5uNSEGKvpK6veffZEUs6b1tAQaPBojBuHJZhfpJ
6m3eyKkZ1x4tKk0VZKN6Ko2VD+cHggU/cfcbN3g1wrHHLn1w65NwUl+b59oFfsh3J1iNcbsX+ohh
F1+quQVpKlEyiWssNGB75060PGY5drjLMu5gzdFYnmfCU9jiYN/wwQl1wlV0R31sy8IOXpDmXQAB
k+ix6U8yn+rE/bhlPlUoAM6/0WYO1d6NBxPJYC5Wzi2gFtnQXrCfmRhzEAQMST0J6gkQVW+mjZZU
BPU3/IL02ho/MRxSD1RaQ3xYROWo9ULFoSaUEcwOzlIQUvIRHuZiDGqlHtb/6V4g2vzboPM2C1FY
BD8Zwz5wrq8ScrqVPxh5otmc4RWKWPKpKoVqMWXvcAUp6X22nefuWDpJjO8Xn4PuGoQ5v/B4pVkp
3fPefw3NxB3CjiTWBjTqqpdSUlJzQQ8wTlw47+xTlUeXhPOzPsRRNbZpVZnIPuTUsKg/788TZrvu
NYxdlFp22JZpGADOAZSI7TJq9HvcwXF+QZM5xHLGu+RxT731tn+pWoHPgw5PTWnG63zeZsPXUMhh
a/KheaPLboWa50PUeuZTEekiMSx75G9VATmZWwpYwQcaZuNgttkzG/aYxmJ+cxms82s2Owib14GY
Fh0fmj+LqgZd8rlYVftT8y1PeRXnW3aa+w90uA7JDK+4e/rzvm1dbDddM/OaZkmZdjxOicGbxvBM
6yQkv9eBAVML9VSOeeJERROVxmJ4Rl31frlptEzhtpRw5f0zd+iRWNtaM+n+C29JeA6pP7ypGQ/D
iq8tfReNRgRRDa0Tz0GolYESqB//JNv50lD++s+Fjxk13NxYhGWhAuORjN+m0Y+AuWZQQJWdiXCz
j9uacVLlXYtAI+hBetHqSAOaTHaH1yI0nVl6IXDiJTcICj59OWZD6SNTvb4gYCfnEry2MR10LpMD
A8XIMJAMv/U/5oJVx5ur5x+n7N9g3AB0NtfA6uPNBS8ojt1c8gW2/vY9vU8Eb/ZLKoji8zafEUUu
mK07RNT3qIV4VbDPjPTrJUf/hdSNlpAXsKg8Oj2fNkCgD2E70xb6iWfBReL2LuoMHi6LrUmF/qPc
qYqsV81f1uraVtsbixbnwOoDB+ixLQtEwE9ZrBEp0YFxF+l8E0hKXC66kmf8ypdTfZaWVX5XScw9
u1QO2njz2TXKAlcMpU8oZB1SUJbsO/yt4+jILqXeykS54LXu7tgikzp2WI/FNn2utIwhCQdt29uR
5wMKXp3InBl6AUM6fXB7ZPmN8RhoKjHjdmUZ7SU8wB6tLgpiZ3dsRSw106usbH4Nbipt8Y6a7Y3Z
vzWNmVAdtuSbp13DlZ1T+wMwZeL/euXbfFLrlxYMjsq7xxPVNgCJQbUrNl/ycEZIGakHP5l4oMMl
pH1k9n/goTGMOawbvqFszsJHmk/I2rA4YIJ+kQe5tHdpotmmTwc+C+Jhfduu0F4sBNwyfN3krmo2
bzjz+i0bX2p1FUJIPgycAbYIU6rk1oK38yaLXLXQnmnXxU5FSmEgvy+EilTJ9aExcd23Cot2MGRI
Or3rhBkmrg8EJ3vlqkLfQGryoQO+unYbASh4SlwMHVdoQbj7U9+YWXML5KSFsluLj9vQRztB2P6F
w+TxzmFEK9h6p7vYikrAh+c/+3R/AeNzNDqn3D6XSr1R7ReIwSXmmrIDXNlg8srQrl5oXkQz0T0V
U6HM/BBHXkm2bfJRfsbumAiuXZ7Y4h1Vqswpa2WhCrSlX8DFp4GE5gRrygBzwwJ976HXxgdv5a/T
LYAWcgC7PlvTTReh2lwbc8dgsFywXwdP/0CC5psS56qUZJe2DbmxOXP/24acMnA3In4sDfn62ITa
Db0unbAmb037a5SN9OLEvoOsHjjHxyHG2bnHEY8ILcw4WJRW5OsAdoEgpMUudVPiNOKHaolJwuDY
V0mQDpEH/hqboWPOyaBFLWGpYFI18mR2v7WlN/vhMoelHlFL0rnXqNp6NUfTpBSYVCIio0f6Qn9Q
NDfome6TrVC7YDx087n6ARmpO+rEWZXfZ4mW76u+xCO8eLO5uJ/DW/p2SmCPiB6uLW+p1FrSdwD+
1BOewEPvNt82CaqDdk7pqrg/wCih6C9gTmZKB2n9XUNH/r7ADBzpc71gb9DPqKSOCElY5zL6ZG4R
OIDSgYNWX6/fCsb/7HGofLIO/MIvBY4wTg4l66KGMbLxUdohNld4ACOUlUlY3mH25gtCczTByRZ6
yO3DTVS05L95ZZsk7JXvC0YmOhVhO1FyEuejvom8hivP95v27Ks3arviOFYFs2DSOG4yPHu10bRR
2/hxkTk1b714g+Re71viM1T8Y6jD/TKMk1Z2x9q3BpfCKGOoPthzGB6OofpWGysFuo1wsjmTECNm
e09u+yF8G1N05RulqvRN6AGRXPBwRsfJit3uLd0LZaG1MIaVE8w01cgrooqup6jb370ek4ox0dgR
IunbIFUrkJD3Ibwbd2TzW/4WhsvauCdVW4ttXLP8SCiql3K0Bq4wXUT0r89f5dxZkTwG+y36qYLR
mkECvWSV1k8NzjYNCUP/BUDY2KUn4osgENvVG02qCmDi5zUxo6vnNjtpmmrMqBZonPgjZO9g7CW/
S0XZS5CbJkfGzyBHfUxFQbooxirLLaLMX/blBEjlUNedcbDbT/4e8euUmljLjAU2xWNRMZSowqW1
tnjuXlitcXCAWUCVLF8hZyBnalyFAxw2upDE1IZC1ySLCn09zqSHOmJJk0aX9B9TiZtwKJdhMKv8
hskU3STV7tMM70jDZVV3wa9272fWt1ZcTYl5+7fj7FwJ28NcLbiFmBiTudR8RQq1HleJISNIFDVF
l3+HniJ4iYK2B+D34FRAMhY2efzMyKfxzXWL8IoEM0+JlAu80YbwXybv0q642SZT4HctnTtZIGRi
jmH+H4c/pJcyv964ANVc6bil2p1n+I3eGE7mPWWb8ETyKbeSPCWSorVDAYAQwVfmdcJTr8Nu5q6E
SK9LdSpJzckMv/G3aA0aIgsrffgq0+D6+vFgaIPkqf2zafNk+j6Bf/OVxKYCgS9dJFQue3+pO0PV
Qrksj3boQopnc2QPaFgwFCo/QExnT23hN/EZCW4oMx+bdPxdpGkJWJ3ZPE+eco53kvEkcliAT9Ad
ZIv+iA7hHwpSteg/Mxkqpl3G0nk3gDFGLi1Hl2iVfpvpBQGvbsaOp2CX5dx2OAMrQad9UeXepe8K
VgEaX1mwmSFX1e39IXquZuOChsujqiipmrPlWM4CbLZlVOJUxhWNtmOO8tvZmwgB2TCixyp/Bob1
WNSciPfGKjwpoW6BiNkVQ4w9sRPMPtpaXTIwCnEIQRvqFOIWDdag6dCKFzcbYvI2gtGlqTk1iLIu
sRVEBgF79vqHN0oStjqX5A41k4fTEP8K5qT8ZwJNLuMP3C69FfUrPbF8VpfyznsYEuxAjmSmvRTL
rBbplb4cjGQOzT9eTQmOwkzR8clycziwXWDNK2jvDCezr+mPACYD+l5cCIpB2Tzqi7eg/0csZsSF
OVIWcffSfR6Qb8oom+mP4m9xjmP1tWDbySR6Kb1JLv/TB3G0dtr/W1lHIwETuZUzOTCml3HV4Pc6
a/nnsdo2VlzZ0r0a1MYmKIwSAFK4tyBkXnTrAfhgL6FQoLBFnnHj4pOFZFl0lvI4htA/1RQdSL3x
GEtN3CHU1sE+K1uFibZQ/JSwRjsNueGFEfEgM+PjEc13qEokpgKtvTUd6fFrLh48h2vvKPiczTvx
wI+vGRqSJUQH3J6wIqZ5R57+i4nFYuNsy6simnil8aiDS/yEfP/2lqKI2rH9Nqt8sVKek16FyugZ
6WDVA4T/dQNbdpjE1xYxghjoeuUV+G8pM6iYE0J0yTZq6Z7+grRXUq9zXpXyM8966pDu2ZXJWp56
AwC9jpLD/weDorIbTf3N7vOUEBuMvDrp2Q6JEjyTBPJy7r07h15i7w1jwGzfCQhX5pLdruOFyuH6
kWen+e/n7tnYp94jLbf56U+U8THWP/8ejGtCVP3VAUfX1Ho1ENHH1rARe61mrf2icoHoec0hB1Xf
T93nlI+0IuaMIWOrORUiyeykjvpBXt9XKjS6RUjCZe/7gKpolvQApG06rnSGJA6ELrVOFQZImYRY
/rugI3iX9zDcU49hILlaVLok/mkb8C+W5JcNRscJdPRv9nASImliJBzmDNcOnAP5oUuthDfwH3Ve
bfIvLTKXCO3y++u9gvFKRIyWaTgtEMpmpEvbnY0JGxitJHIzIcECX/4O5/0Pr0rP+0wLxu/AMZhN
ong/1YCHGgCfJuKd+V+PUMahbnSTQozrq3/3YX0CjBbc4XNH7HWjDShR5LTUSAVTqz5hou+pr+YH
4ELTgPLSkq6BrDuc2FeHXEJWzPguwBY5WzXWWfHX9/Mq/imJepzHwA+9sgKNcLstePKj3Q9bqxq4
slYj/qf8bJ4zEIrGPcaQHeMUqM/ldvbZ5sw/ZIbXRL6CyJcWjY3CA2XXyE6wEvUfkRouFL41hxZ5
xp0oBMsGVMRVeEwAO5v1Xvw3USEXny15B7gv6cUCgaL+emPwcqKkC6qbcKxWgijzQVWfE2t8/oNC
BKLmrWCeAKzwg3nCPcpYWbqdlg+DT45z4xKNuZNDQ90lbCUqWPygjNAEe0mTIIfkvZhrsFyFU0oM
yFgTpqIwoQHAFrc1WWxUCwH91OOfS2kwQRMYW94YmcRoXMYExAqaIRRVtqcjjm3LG85nRutJ+lan
tGAifi8PFaJEAlK/VtU0Uck5ghnY+st7OKOjnFTIGEvuynKmDppDg2wMk0D0U9q8bD0bVBgO7d47
vW7ZL9jY8VzHklcaDRh57Qs0FxLIy6a7zEtYkJnBKAk874mBBu8EoUf4wa8NCVatLnqNN3ByOvYv
u/tFQXHfbzYL4yZ7V5F+5lxdh9ORnPhBnodIWh98Kh9OnaheyXO+88wIFPWUI15EeMZdTffrdw/J
pQHgM/5ARYCh6PZGdN4zVYiUsGrscPAHUyM9j/6tcx8VuLeaI+0P6Tq4TUJLpyOZPEoDsa/Lt8dk
NA0v1DuwdF/Dx6yZIFoB2RSAEuqeBFDTpapn5DVCxvj6PfbzM1/LUw60typF8xaNUgYFyrkgcIOU
VoBHl9kp132oJMLMMUtFlRlrbNnkswHiFmtOZYwxV6zmEGRD0RvYN9/t56fewNLo8+cKnLp1T2ql
2y2NuW135a7pneGPWSggP4BcJfiFBHpcEONFkg0P+p/HwVx2PsJhFPW7nVmp7nL5HDs/P6Ssjzq4
iqXHm5eHRfYys2Tc0B/TCvNGcBGIN+LbUARUhb0Ey5MFWca8wfocz5fVjjkL7vRzTS2wny0X+bh/
TeOJBadiJePr6nqDr1DOuZGOlguxu0nE/NX4MFcmNU/zExtaa0XfBWX0D2GTwkoJYq1wzcxfWcFK
6NTg3jS0UH8KDg3Y29fq/vBmQgEqm0B8mLxxEa4PGSxCIEGqLoeq05UzLPSabfN6JvymCQK25cgX
0Yqd3qbgg3XZBBXwigGVpoPfj0bz86eQSbugCQm0Xi85phB/WLuNSHGatG1/pjmLdnQHafe5JFbB
Rx/7Vw5hsk+96DSMzBmpC99A9y8MB/IhwaRGYu6WjhojxRdXGnLc4Ttwl1iU5gDGZDlejh1c3J2l
UKQ1jx3tczMm1SNK2HOwtMw2mMw6vTK7P0ULgvepUbpfUJFFnLUh2sfTwZjAxRRiDtZ3XUbCdMf0
Oh/K3T2Uca6BV/NmbckGFNPb6gOn4iIr0BoZsc7rwzeG9qMvzdGCHbbeZbf4mPJ/87x+0RDIElZe
4f19FIZuOxMZH8zumBiYw9JRG5KrjxXAbycorvYXII017rtFm2NBshAxcq5ea+jfkp5gEVR9EhU8
xJofu7eJURr1OH5IPiuLxM+CYduB3EwM7LMD1zRFovDA3zxc5t+W3RX4KAZq5Z2eYzoRCafN6zAF
GQAlUzVH7RCbDWEQiTrJrEldD9Gs90cUyP8xbwfli3AgK5hwXHtA9QyrXYg8nhyhhQzRLcQUMNDj
OT8OYfZOVWF5trl3xQ4vEJYmvNzp0PjpYajXxCMamEF30FP8LJA0R3/pN3XqSFYpy86xwWDIpBF5
wEz2/k3Ldr/8E80bjhkQFxkTMn9ROoR/6mXSwKchmg21O2ReoYDPaJwW3aTZrNnLdw18tvYZZYjB
oDfC4akZOoyrUnf4MJiEMvgksPBYFwpSIlset+LkpvQ0dqvdd3fzUzSllOcoI4kjv6YzI3jmJC9o
/LKI6qzXiGgpdehjOO/rzDXLHF5SEevALd4s9EhhSqJaJ3kJXITVkl6SkL/hOs4xmkojR6Ri/1iG
EtjUvny+s6/JnNloWQ+aenn12uduoqE53U6zMOo0gtO1QhggJogUDIeFSsWNVvWjfOZkkVTgsjRo
Rdcjz4Aa9WFDKSaToJk6yaDadaHFIz6mSdRM2TLzrESusM5uatvPCW0vAZbOSQyeCL8UNKo6OMyA
XuQ6Hzc/BT5hBc+ihpxq/Q0zTmaism0qkd2gAzC/K7QHoklnuzcoGg3pDy8Zw1+ZCLcMklk5aG2z
0GRNNhJ7N058v18GxFgzf6F3rAaQU4ug7s7mRKYXiauYHrm6eT+bLcN6ZjLHGlhhEZ3UscqdGuQH
+9WMEuwohG1noCLjRAOa033J5w5hWR7wzOCueuutgQz8zITQomngSDftnMM9eVlsq/J/++cs8w3U
u0u1pj7LzHJqaO6+uIh6UqAMKdHYiyzIGUTIbLuyHC1Vdpwlc5LkpvkN5aa78e59yZLSnX9vb25e
zlxSUV865BsFYKc7QbIQ5OZcJjJg7aMlz2K8Zu8jdGIZsGuW67qDw6crxbg6TxqhwZFJhpSCFjzY
L0ujnUMCtZoTkZiOXp8Fbv/PO0HMHKteoInYAhdHqjuwZYtGrwgPSrVWTnlWc0xCQ+4AkuNMLReJ
Ns3ox9bX03qGGEGVbq3Y3anmIK4++G8ztRfVlDcm/v1UdXQdmw5PRW9dhxGbGVRfArILSLBXf/GS
Vmv6+7dN8Z40ePfWdlhMAdhveMcDnTEmRhDFJoOmehHam5WAjUHkTdzSsFq4Sbdk2vst7GC+h3FM
gEZJt+lev6VU47vfeldkOAZlDEcUSUIo76EOhXCW3MocEa7xQXa4rq0RzAV/k1p/T1lQhVC+cAED
VIUkdi2fw7qQF012kP8fW88a7v0gvDQDtv1dBclGZSTQ57HbkUkuGOiQrV0SK/yme1G+qIUUFmOO
l3FXDMAWBM2MeC012B+8PjyufshyoHTD+VUIj5jZbwQHg45locNg4YI+DsmB4BG2FcHVssbdGiDI
jUT3EGinfnyw9o/ugn/+VAwrbN+VLJFZ0z2xE6F2WFRzhva4AHGcOFP1HMKsAfuJlJ+MegBwKNH7
KuTSh/aVr8vQCA8LW+0PQutz2P2B+E+f2IzqXW9PtoWaj6kMw4ZOSljSJ/0iH9LdOdJJuqx/4u3Y
xJW+wuGQGgJra/l4sv6m1cc6pAvEI678pN+OLc95yHCCmjNO+S5gvSq4AwPDvSsFJhl4YiZpaVlG
k/wolT3ZPaQKTvmwj3xFfm0ChMPKEEGbsu/ECooNjiiwfN0WLqS2LWHQKw1h2o4U+MMHuV3nnaFs
j7H4g6RoIzVAAiArFNQUkeHZBBSehUhQLSyPfIWmANPdbHWzCsFFE8vr3I6b03yj/52fwmB/5EOL
rsweZ7PEsVtBQ3Z7cu+iOSsPjlbaxiFQxpv2dxIwKIt4BzaM2FsgC7j2m1IjwwbqexkgeHpDcX+B
xscOqssqK5DaqQyWZQB5/mxrG/m433Q3eKjB5SLHuI4giA+almmpTrnOlEIMvcJ6Zvn4L2HXLb5o
RMzTHU74y2mpw6rHN8Jc41bt/5IfIWNrxTVpEyW32sXToNbFjXbK4+c1ZgnKVhefEiYM+ddjhNCw
skkAzw/87Ar0DU9JQqAYXK+HTZmF/LLa89o3g9jBbt8XY5a2c1FBo7Ja2XOlvg8TB7uEraqz+NWA
tspluOXelS+IAJ/yZVSQ54FmU/kuiaHAGGyMUSQBgdEWAoYT+UfyhjJX248ZmSqaFUez41FP20r0
zaLAA2uRl6dvnKhchez0/g9/z01KAczdQhXdlyCajZD1GuO733bODhipn69UdBywrskPsaOKHbyo
+IAMDX4HxNGHHlImJQ/BnWaXHBqYXI06K6owrIWP7/qH3Rbxb6m271/zUhH6EXwUGJLZCazVrklU
E0QBRnXldMWCwCwjGUyygdFszbdrFqxXGDIJP0RVKbjZFLITzPxYkV0uXu8UZPM7e7KKjs0xBVmE
7dJ+TIM/rlnmBjHYBo1s4Mi+jlOkziKYctTcX+Uxhu1s8octirJm1iwpLTpLzjyVrQCkF8XAa9SE
Xiu6Y0grszaYgUH9GE0+YvBKgNAhuepEG4dfI0sYtn202uMIR8DMLjnJRS3/ckjVJE1P/awJMjVo
8csiYlaBNG80mBYPDuvuJj11zwNpShtwiB7bpdDesHtKN0OrYsFmKHEBwK53iJhnAH8IrnZktt07
UwPMYcwMHkHPrOkaZiR17K4ecK2fQh2kLiMkqwgWlMUJeqY+eml0ALr+rHpvBprItHhApyQw6bwf
FuD9TADKADXgHNaKlRQhjhJodg3cB8egxWRx6cvdSzZzZ+8g9GW0HBp3oUBXT7PzXcD52JlkZgar
bnZgHid1konkO5dcfeuyj4xfVjhpx0jGj04AL/aGdZLLkxQE7MO4HxfbYJ4Rh/2PHOqktV8m2IoC
2RN/Fb9rMSmDBCcFOwPraJhHMWc3LAZ6NgCx4VT2KeCXrw+wbyRrQdzMbk7vaadgD8VKyW6PrIBE
tiGvhLMYFtEN3lB/k12CIE/Rq7YvXAkm+eu3CsMztQxcz48tbl8+Bm1o4d0oSlmYfhSxG5W0Hdo/
SBa4fmvVSUONmSR6b9zfeRCP8UQlUgImMeU8Tv+fpFgeMYrh3jg9/CRDuJcpBNR8EQBpWkURlSvg
4nJuUtZ+yKvMTBADL7q7C6IbyJ3UGYHcbhKze9ghB3alSvy1nTL7KCVS6yy/wr71rAc1oAG8tw5t
xdo2pgkhe9irDCTQxO4kcIUVx1wMRgsrrs7Uxz1wAOMP56MSqfh1Cpi28iU6G/HFofEkoIMSZK/9
+iacEcWtjptJ2FlAFIIZ78OmGxucMk0r6O3BYBy49JPHjCzm9i8oHwGUvyPEnDCHROAAlytgWTEh
dLMUHD//JYF7SWVPp4FdNo9ADdA2Fmje96NNI0L8mY5k6dVoevv955a+amdnryk61EWKDiKVnAT8
AzgLhEd5xkUPqKIftvHPGAYyidm5qz+BR31eKcXrUDu6pm3tfzPjYbodp4BRyeDI9D/jv992yyRj
JO7GNLEhQ+5pdEZJl8zQ56BSOGC6TmlLIx3PSE5QQ7Caw5U98acBPx2l9noiTWgBR7/++xHM2AOZ
A6SALtVTRwuhMwkaaf1ebiIiJDlRtTw1pKtRqT6rgld1oSjBzztBWlch8R+sveTlbOJqz6oUzc7l
SzOAAzIgnNcDvFt5ZkNbIY2yuFtwhH+fxBPj9XWGUE2/zhSiD16pVrqyP7a9NnL9BbZ22DW08Qw+
7JSebBphWUh+2NT5mEGX2vwxS91oqUrIVjhEBM5TcxnrpzIpAgrry6EgCUgQm3qiGcXyDazWj4qh
FAy08JtB1ztjwwm5Fu9Ze10lLhVibbBwwEc2BKfeqoOPmGnVOE2/0q/SPdApoeBA6OXIQ2foWYIh
RY4ejZ0gImqc2Nk0B9Ec2+y2pUDKSj3qdPNnwAw4gwQs/vkCC7R7qjRJ2iHkoJBS0D4p/o66uNue
sjaHBnSapFL0oSRnt4f6kHclXFZTZLLS8PlKOlQk0+Kp9OIa+VT8IYyIulYrhr8uy5AASOzCe/XG
C5bb4a5NJQwXHODqByhtoBDwlWiJhuIYhdwesTva9g7wRjoFPsv+e4ThWVTDcpN3/s14peIZPPcq
BRRwN5TJN6fDH+Vcjv1z3EPvxxwprJu3Kg/6s+HCQi7UHwshaLjHogfeKvNpsHxLBj+qxx5C5Pv6
vtWgOgwkWXm+NIP5Zoaz5/HnQ3jf/0R41XKXwErqcr8SmKmKR5JN5/pWFIaenFVoHntis1rGhRm+
hEcSEgoTG580wda4jOA3WvGreM0yqHmZ8uvRvrC0uV0PRiJsUrz5xvXO6CqrNMmSvjaOCe6OgUat
iHOm3tsBlzf8bFFMqGYUHJ4/NbrGHSVatpM/6yw09OErl/IJNzCmDbWarGQBme/vAV6Y/epzaLmJ
+aPZvsLRHxXTa6B8N3+m2Rv+S1CTJgKme8GsDHt0dm2JBekfCHJfcWOszzZ4W/SGFxoYSd945oEo
DUnvj3w4IkajGFNJ/PwMw2v1am8U4YSU4kaWNnjzjd0UqJQyx5nfGesGh1VGmXbCmrPw0nthN/nt
B0XBq9Tn70318ctraieksE+TpSyPZgLz267HsbqFAL6xHm/mRkz5czYnzrVoRr1nvadLJEGr6aGM
9iJ5NBE0bhv0ws9CmvJlzvLEaDFTIo5GUU0F9LSFFQH8sXRUZdbHkLTA115O4Y3wQCKEfifZSw88
2I/zX3B9aGgl1N/e/gwc4v2WDUMZtYZ1nias3eTA26O9rEhL454CKFbFGDojSdbyjqbT3fwa4Ne6
ZYS8dcPaxJ5Opoi3a1YGK4rosgQubksObR2EYeIIe1OPKRe22wV2X15ahG71dJn9IY2ESzaBlYki
CUHysGbheWDgZw4zuihIz9j6KZj8M8diJSii6kJo9BZ8oam2Nu4teiJwkvW3H8YQARb98FmLqc0i
dKKYYWQkkQYNdLpLT4msoHSvh7zgtIprT0nxgwq60Ai/0tB0aIIpqnA6QVLj+P0m6xwmYDCiGiyI
AubJgf+XaeKzeAZCRqwNhUflLbm+4lOgWk9mBAXVZoM/xpyz13+OmoWVqb/AQmtlJgeqgNoA9/sI
61H9lKgsxSpGdjFGMEEJb7vxCkqLFD54DfPDpMThN5qXsep9rSM98FL/SAEVDEnPfVvBIy5dEAo+
Rsuoqex+YTf6EInxAxjFQmBA5bGMZ0v4KDFWkUCJKzK5yuZ+fiuPVSYZTAjMDD00/JZeRu5q/gvP
vWt4DG3lRji0+bPhVlhWAbRXc8ZX0Nfxfs6H4BBDImc0iL0r1tOCRbYyJus75W/bFk2pRmbPuNd9
CXRNHH8CHZC6G93OHMsyApbEwYWF9QvNbEbL72B/dMkPAzl2ugL9iMNA+jC2rSnRDEsEiwS8sum2
mIXr1IL1CD3mD4bCNbze11mIq/26xsZrxLjvCtsLTGlXgZdZvUBWtiTnp9aTZ4K6MIbm+9o6/2mp
4Kq+617mV5iZjjHzuLMXI8sscUD2oFhEsmBLMaelZCswPxHK2ikjSIHcfsVEeyBi2XFTtsNBZue0
7ItL57h5Zhk6VQimCT1DPpx3r8TwmpecbY6kdjXQSpwhIsYgG06H30vr3G6Y9bHk8m3IV8F/gTA7
UCqEe7N52r4oF4/K+o/piZf+M2lbQuye5JtWHtrPUcDqENxPReG5Rdze/ejFJydBLX5YWsJNXAAp
/lp0BbiGR8cGZ0/9TWU905sBPJnxK2PLBLiuMoQvGxxjCBzKa6lW268USNxErla6CxyAwGvI8vA7
ylHcs3A5ydZ2/qoOOxG47dm1lJ9MSxr6D4H/SBIvn4toNUh00xYVNoIXYkxONAuUq+9RCOxZU3V0
KwSJ+YZsSUC+HnCHKlnI33GrHmcipBxF5Hr67woQmQVxbMBdClWifrnUB2X2C/CjsiIGWjBp4RgR
HnBBgMTARuGtuFgFtGqmTAZhofE8E20GR9D+i57BMT0g1uKx1M7RzGZeynR29Ove42vyOT5eCJtj
l+SSYsvh3AGqkOhTR/pNBTL6MFM37H4g6UdOlzJCZqypJLEmlNsRF+5fUimHWU+iGVcPUVzHRnPN
3CXVMnQLZi6AVAVjN1tIiJ3iKZN1m2ox9VNznkyv/sZRt+X31q0+ahNVCA5gJURKiQ6J5uYFCsHP
wkMJ5F2zTJrjWlBzrpZcbxxSP0AjXCDK6N9cS6fgd71LMzw6RyYtnz6D3R405rXgNc50yv7uyUf4
Yfd/4r+Ky5pvN14gIB02YGqsfa1fz8f+9h71Gy7AIL9Axhqu/o5zQZHUoWOEq2PxFsfDUroC+uPT
0AiMuRaE7wBTCiaggeEBBeOAGA/HhPgK7m8+ZjMTddovkoKwmJ86kuQPEDcp6k4ucrlHwqP7h3qF
94cpMiwIbixjiX5B+T9er+75h9xk4OU1YtDe1XHsP7vkS+HM9U+SUFEYjJ/Vw8wPkaCyFi4OYNGT
U7WjdD8tLrY6tdK/dxMx/haL4z2dmTay8jSB1agTHFv3bRS6HKK7XCvyDH/6fcIrIS7KiuZ8KBJ2
SFrBZV3RN2mgEyN8Jd5clfMKMh7b92+7Ry1uPVUkUgVmHE0FJ58QD9KCEClNT0nQESeQvZl3pG3n
xtMpahJ1iwvz3EskzzvebBJpsEQoB9LtaGgfiASG2nbvIjX+KlAhIBk4QK0VQ/LRnIKebhz0Qovy
DPZdKXl0birlxharr2KyUhegRVrSQJrYK9qTLxHEWjoRVgxuh1dn69/zjntY+qiBjOsLBnelInfa
hqX/S5J8V2sScIBmIQisvaFuUCiqQNUa+3myAQ9nhpk4J8dgMq1buEaKHrnoOOfU+Ivmg3pxEN3M
/eSlQOO80jJJtYVHHz/WA52MTN6kCIzwPxzk/Eij59dMPV2KhtQKhdE6C8KPL59U6kTpI8NXdwMX
iu0nHtKayiqj8zAfWXRjPXJq6moyZJsKsLnIVvFvXLyDS6gk/EyWz7J1AZgJBBSmCZ9zX/QKTSmU
mnkRnJKQlc2hOdBB1FLxuTtSzauj3uWdDCIPKzmXmOPqSS1HLStXJR+snUmGBs+4bsM6mpw6HIBD
JJxz6WGQOZZenU/j/q3OJoKnUGNsXCJRyOV86UuUZOttyjVYLorKu9u6bn3n8rNpEXJqB0fe8TfB
IQ+4Us05pX52ZuVhwnU34l3ROyJbx1j0xnc6SOzRatgTZrA/7ZP93kXF6+Egzhq2aUELtGbszxi6
XVmekO/7UWpOaKMyQZq9EYObFwmVimLUewfBfZZZ7hT22OoZCnqyBkJUSVSDDWYEDxvkyqVohk/M
cO6B8ZUdq45qunFkfYja6Gox9MVFoFf25yZkqeWBy/ZwiAYfBDAmy9OJij59F40EK4PP/dSSkOK1
dgYjXbcuQxd8b2lEltfjUHjIAYr48NXtc8M1BP78D1I1qdk1jGMpCXyPxW0MhACpyVYxUfWxm74Q
TZeMH/ZG5YcqG+J35ZoUk9kL9R1/8E7ExKHBC8kn29eOL7ovqdX2VkYtCXSPY743c2pb0YLM2Hba
E6aosvWXXOkj1xrRU3xCdg40akOR9UVz7PgvOmwWuZ1i0+hRL/AaZ8HhM+BR5L+rvoaLK2mVAIuy
frisv5a5LRopLCPCapGBROsjD9DyDc9CTYSGX64I7wz173vUG3y0U2TDTY9k74L8fiPoFAYdSmkl
1+Hxd4eh9i6fldOTA5kPPBwBC5cHVPHLeSepfnaLrMRvrS7bmZXXQ+OCTKzMkZhW4x+psSwUhLe8
sOpNPagjEpeImvD1q/rvGEfnlNC58coyeneqcu3JXkkgfqP8TstpfZqt8htLb6fIFZt8tQ+3p21O
8RMcSH3K+ac3F+PXUKaI1OknQIccVxBXF5+ljuXfUqKybN/QIFxyp1q6Zq6wZN7qRDd5XFtmd1ud
s5yO89rhT2i4K/TsV1K4j0JkWGgWWGwLGPRR2bC3UdQHtdbvxE6ibgDIgZ4xP6lrDht6ZA7F3t35
/NZksW/4h8WQ2/Fu0SnCr3kiyYbfCAYkgZnK8fwCxjB2KkuKg5GGG5kEMOcje/0oldfBECO2YB5M
RKwTrafZVDuuNVTK7qORKjRN0y+dOryVz082AybYN8FJK+57x69/FfZxqSVsHht3Dlz3ikBPuoVV
N2+rxbC+QX8KLhr9BHzEGm7aIL05y0uqTiZ7DqNu0DHtNK8eIi9pT3cLKT+JV7Ml99xAWaS0e5+6
ZRBUwyp4yip8ZYiGdSYdIT1NkWphrgmbzgJyajxBpyj2A1uoK4sTgFc7cjK9ku3wr75aOllOAk0P
ILKVNaowRyajZ5ABDoMDBvr/Yqh0kR7/QY9TbD8h8PhZfmQxOJh+UZXJhndc3fkAHw+w87q2hjSa
nrgtnSGr443IpCjrNrwSsJ35E6rrA1nHSpWXH+qZuDXisLPNnjO4hblzhkMuN53QraGLXAcf4IDS
hZSQGQrgCIYpwHkNMajFJUwBgnNk/UarfwEwvrVeelLKDOq0vt2Ogu7YCJWAa+MLagGL4mMc6OrA
NctKqNjSiTBBytP64p3uvifOTvcFrjCyyAAUPoK/A+KiIvisO13l8WZyYdbenOEAcxzQo3dy/cAm
yv7PsmApCFOO1UWCYRM2tPDnjgqmuOU9vEmBwqR0XlLhbXaa/vzbJVgq/Zwpw7535wUm8thz2+vX
wvfQkD1NVoaxUC5ljXJhsGcXuq6fcVfwVrymuJMGsTgc4T9JxxV19vJeGTj/SQVp82Gl17ODPxbS
CIfMltGVqMER9qvRmHNqxApZLqwej1m8OC2N4G92OrT5z8l4dIiuNQwkg7jgFUd0uqPlQuVQ9VCE
pMhypKT1/Sguqz0UZNJoTcbhcVpSqdEtlY910XRFDf+dUW0j4TQf1dzsSd06b2ySETbxo8TPhn6F
D2PXWw126OV/nZOaWe+PGd6iiPyJvP+87i8THBwJBTP6iJd36KajUBu8Ipzg8o717tntpnU7tDXh
FEIY7EJx7E225sskRfHZ13mttdbOcbKyGOPNVNJ6VCLcOZjVuNSJ2JSNENICylalvkgqD5Ij+b8p
KM+uG+YVa9e5QAgYTv53jvXLewvVpVL+H4tTLCY/ENUtqu7oBKwQAaul/fl79s1r2ivk0uKOb5pF
rdXezqiG1+w03zk9BMMpWWzcJYX273GH1dnFyTWkPEH/8ExUe6sbTFgbAH1uL9+yZVBak+23AAOA
GhzUjWKahAcj50vTmRTw23IjH+BRs0b2FouHr68A0Gm3SAe6rgkk0pCXNvqXjC2vQTQHvLeGFvkz
hP9xPTxtYkOTbkqaaxvM4mA1IkJC0CtMdsr1JDOo84Z58J24KQljBW2wRLWmH0QXjnV/pB7amvHX
9U7V6KQgl+vCTnzzTscRyMTbC4oCvr9ueHRF25ZDXbXEbBRpgy1eSu8+fuBdsuVDAC/+SKYf8Jop
piEnGaEzW7/TSGa9cajcVDD+bycu58InGYRgx8A0wBch7XI9Uj96nW4N81LomLVyQ8MGHwQB39lv
0VrM9CbONsb015cZvC3kaxVlErWemfqQ4P74Fc13AI6cbTJCkygjpBbbsCWxbLKuk2NiGrnadqBP
ijKELQwdWOnb9SWc4901HqTsVGrpjKLBGKtVfUIc2739kDGgJemL3nJlNojiLF6ITuVzofnU2aPM
vhkH+9Q2e9+Fowq1ltCcaVcUq1Vudlsf/uVkiRbG/rE9npw+UYEZolUDzDBucEnAE6mtNr1Gha5o
2nucw8VznIfoc637K31USnrcB6Gnh7hkqnfavTD/U2ftNkjqgKjzJkcU4xw6EuEA7X7J4vj5nXTs
5dnib7OV3RA3S6C5b2hkB3BA5xQi4WOH/c6/YksMbYCu8YwBE+hXKsu+KBxYWYaiEd+OO3WFzx1g
/XxyueoGO7yUy8mPUI3iV00+DsVDQ1PmDaL14SwtjgvPiS7N/9U8LiI3ekCyf2VARNZsGD3LzeFG
fpasC9y5mRZdgLGlaL1rQrmPTRyEzCGFiTa6J0xq9+2JXznD3Ol/xmcwvNqkunDfojxlX22Ae+Ii
6eaesLIT77ac1ywGbMlTvFAwNoTvUELhS5tzQlg8iqXaidXGWZUQMgdhEe4MGU812blO5IvuMKD/
FBlEH5Wr0+uazs9vk59D06zvI6UlnQpQ5fDAXEUDlx8RLL5NW1MBc/EGLJHfBkD5JFIUx+poQvCn
E3O0wpZLBUqauQDdBuGN/zpLQePSsAIAXgQ8VeYxfI5KQrOE/efDvElkRSyc8+Qr2BM1yQlTFef9
S+dBBJwDkktNkDBJ65Cq/fRcCMfKfV85v86MCXshWc8TB/WlMLTk+zTCGP2ya4cCKAHzRx53BY1a
sP5r/AfM9yZ+QneyVhynZraS55+jIObHcRQzr9HzXUvSHDQk6sMsauTeCYzY8lHgQNYb5GNp6zln
uTbrQ2HxWv6Lffu5vbQ5BEfK1i38PGGeHO6Vcw/f2ow3XBEDlpcH3eJaRRDv4n8LLKxQdeurVtbB
tIuM5wuytm1OAL/9o5LufSRpJ8J7ZURkv5jiQEh1rQrY7p9q8/vKbGlRdqr9fKqA3RuefgtrTMp8
bNSfqFaga6p4hYHvpA4gN2BoBmDIAvPppic+I5d75k2xPd7rHbhw+SzWVe2qpMGluLabFs9rNtoQ
k/d77JW+eOajarcs/AotVttf5zTHeq8vnbLTtp9l2MpoGtlXoUbChQ/5e1h7Kqhvx4vl2u8kJOCx
8KHYClzxVwdRVRlEJpTOyM+vyzxMZdb96UYwtx/U8IpEFrsZMzv9qQTSsOZ8LcjvczENaeNiDQ1N
wgRSiMo31rFdv/5kATd/ANQhskexxYruU7LiTeiwhjuSQ964iwQM6IyOh3DYwM4x3cOJel3t4NUC
1aILE24BxkGv8wggRAaAIwIN98yW9LMqNEQNOvsv8Crdg8s6rFIcDMeN8Rlchy8H8OviHqAT3W86
SJgpk9DWFIGFB9nQbr5c5N3F5lGUgPbJHjFJmhUc2uNZ/IJFr14TuKcGXfeAHLSEJUKtvcI8ags+
uJUXzPRQI13rhs/uj58hOxx5STXKNQa8B/srvvUe2QJKm1qc94N2jRfNDW8TPUQjOtJyK3VlwC15
UfF9wLPL0yzROMrhsh0Cg0RjV7Kb9PofcrHWGEj7ABWFB2a4vuzKuOnPDisRnughz8LHexE6T5kZ
bAZO0IrR8TFZNnfLGipe2CPwX8Gw5THAFQe0GIml71fyv3PV7Ux3v+baC07mX2Lp7fJTUZbH9qa1
pubfGoZzvlr2NIL9IpZZS138v/EljavieKeq0B74zcLpJyDoQGxznp44mF4AW2Vu3lyjjvQTg1y4
Tvu3dtVwUmPIccxGoskjgqrOkg14SjAml3ug0HFMWge3TpYNqKJri/+FRBqc4sBdwKp6r1jqdb9b
KAICjeeE6PMeD5FjeNGAPM7xMlnhXodD70jQLQl8j4dyqL1PRdwmnBc6bgBKxbOUmoxcny79i2MZ
m+cEADYGwr+WIil6G6yJgbuXo38jXzoQveLbX+bQOZJBB48qfoLmph3wcRYUKKLZs7w8prXL1rDn
GmTLCXbuy+QzrKkFH3G2CGeoXjy4702rtKDQYRYop5B9igX0GZIhQ/t/GwwwuUviYr3VbwUAU74L
FllezRqhjX9/Ivj/Xftt+twYHT/IRQhq4G4KuXrIITomJwomdgXx5Yl8fx94mTD4T+E4UhxpfKU4
Xi3IB7ugmEVeBQD5nHT17chClKVTGlfeSebCZ3dQtBpATqq5wyY5PLs5C1qokzGQ33z+m6MjXmx6
1zT0TlnAwkxf/b3VHtfcPZgn/N9Sy5Jxy8/IS951LQ7xCc+OidJ7niLdr4J2TS9agf+dlIcsOC3Z
XBSVkUzvrBq4wPhQNGkgAZXQMi/IeHk+K2ywagQoMTzuGM0uS3xgmP7D9scy02cYE8p1tVfGZw+m
6hTP/vyXpS2paP2Xta+Lplgn3xaAxiA2FSTJjHSSrM8Gyf7D7AeTUhvj89LuGieA1dtxTVh8Fo4g
aVhjuCDrX372aPRX+xzWGgg3KoHnMwTSLGfJC8gqAbsgyGUECWy1kyswVdpzniwDRlmpYUKZK7iR
ub6uRIdn2wJaL2ht/SRSmFQdlImui5vUdlevO8yTlfHfsNHg/uugSFEYaCtarT+0HRYFirV76jPM
L0CvReSUcrCCNIZeCPRoFKa39Dd8Cg+dsPYiPqDyutczbg1T4hlyw0fQFzx8aUxPzdP8TvpyHzkC
q+IqB04b0ZyYelurYdCXAuwsv4EIGsIz5U7dNEY11kNJWf/nUOcZxNc7xoKD6g4fbyGIx/UduPN4
N/mny1gB4F/ycZXrWowMD854ztr9mA+/wr9+1OdblTfzHIDXUZJZiFtOgcrMVgIeGfpjWbZaO/wW
eTUnjuozMLO13ZShbtYbkQxRjoFjD9GRsuOOlvBjfHX1o4rpLC+vGLz9DoUsiEcuM+p8KzmK/i7H
imRUwLdDqVp7mM19ZXImcz6L9L1k2TFm2gtKccvES/0nHQqnrr7N1HOjoX+/A+tIJ2JZZ+gDkPKZ
N2Dx4MdyUxWNenl+HJi6jK68bgAaF0JG7jmSnBM5ZEhOz2lUqz/bZG+a/zaaSwtGrqwCDLY2+vOs
26Ex3+dhvgUv7ga+zMH61sOyru9SpLQzGXuXkYU1vQw2oFNdgTcvokNRnpBZopezYxKnCLOZMSHY
yjHLmYQJLYe+MyGJLvFVeH4SDdH3Ywr0Nj9T4K5ZajsafyHylLO9jEeTozLUeGJ6z68SyLqL9q+D
m+uZLgpvCsxoY6tdp+XB0SHfwYF5l25Nsmh46TjU/iaDLn6Ef4en0uNguVfswru2/Ftm5+jkZzu4
IGM5LUYQwIb5B3kJq2Pu3WQ7qSeMDjjkiv81GC6wCpN3PxmuVBGCAG5Gdcgjfa3TsLjioDLP8Igb
fePll476fCb6q5nVCgeoEtefuUaEBkQdcdCH4ReOuzzi4Jj7LHxpwTp14ULed+m183xMYClvS90v
DSWA9evJaM04Ma5Pl6jc0gGjFSfR3YD4dIX1QmOHJHtcD8bBBwvGjZi/uW7DlwVGrT/TA1Wl9Xx2
fDCkiIW9i1bLHufXsuutMuujYAbhDKwCfvSaqwqWSWpMgiE1zak4HUrE5t7gFmrC556a7l08OJcw
ej//J9Q+G738Wiwq7zA8Jg071CyT/vSPOBXCWkAnjFiVhrSmbSR43dRj/VI21BrHpA9ntb6FzI0S
ymspTBEYlA2lao/9XxDrGM9+P7rq8+aqAIsO5RgNjwl7CvMF2z4eWu1kSK10U6mvMHs3reju5Eow
hkrakmkO0VC6hV0GCXkvDgYBY/OejyXQEKjQOWiFN/ELyBgvKV1QeEWqRSasgJZrVP9fofkd+efo
esDptDu+YvZRRvi/X+VnqwnK8oW5DHTCSyP/cvEofb2Tr7wSlgaFnhSDQ0shF9ZpZvHYjG+5y3hi
arjQhVSEwxEeXwiDCf29w4CdROo54Z4/ymvNvQ/z6jQDdNJzzX5zyJ9JyyFFRXmUAwf4XG+jd/RE
ChHXPdI9hRSrl+nAj/bbmUYoJ8/RkSRfM/43YXMwtplhA63lW4we8yix2ffrxDmbK1m6G4hgVGKW
Rjc8rOb2MNcaGBObqynVOP3Rq2ljZJ7Fw4ZLJyE7oBeOdtfDUVGsPH2kWD7wj6pyQtPpSaqqYjo0
++h5hAgSUVzejGgrPU92Dn7PMpg111g4IXo/iWihLFS/k+YBGhP45uzG0wuowd4FTGRPZlkhmhg+
BrUHtJtRIwcQuHKi68TNrmn5jhEOxlhty0hPOPYhe/kNFi3Trp3VvozFGBCamtLSuoC3vbzoGNrP
Znm/mMIchNMBOIts4kAnIu4hd2hGIPodpxsiff4MTW+4YIZXe7g3L9j2ZG83D0UGBgP3F4s/nZve
TuBnB+B7+SU02kBnYPSeA9rLApjpY9JHSjRI/WRa2m1ELOS9hhd634fMkErvPBhCf4Jvh7wVL6Bj
ZQ2jEXz3wNVxR4jYn5e8FV046PCASlvwIu09kuNWG7VXfm/g58PW4QAUgRYiZI1UUzdRSfrOYLEv
xWHSItJ9L/qcjJpaMAacHJge5gC11HUMF6Fxfv4UF8EJxzC+717aRxIDZ3gaguun681zAUhmIEnl
tQRbwseHoHhXu8ENuCWhg8r1JDBRfWWZuFLTYjgZdWCI7g2ETLYEojwY7LIXAgcMvKqr7E44aV3j
kjrZudOXplMlYdJbl0gQEjGCznMkbxPbtzqaDCokBGai4zR+atNp+xZPg8jVYlvO23Rm4b81FVog
I7a0wiwJOdRn19ZeiAfWbmF0xkS7QO6znwc2Gu0c7w7fCSL2l6DR3Kq2H77PDTu5SRqCG5gaKKBp
bfQWWf1wDdPZqrjUJMrrx4LkfE5fSIdBq3l/Qam8TqnDEVRjX3hK1LjfI44i09qfyebQYdf4KpPd
nGX+5UBab0nFj99DkFNfEeWQ0ProGas8UppXDLZoVUsOZBdWVgDxGrXCwlnVJQuhY9AsAUv6Z9iG
Jf/rQ3gYzzdKd2oNZa/8sCjRZQWMMFQGbto2B7aGpwJK3UiwZ2dQrCtcEM5ZEVutzD+IwdluiiKx
d2Jkmytrqe7sp87XxdcHIFs67gb1Vey9Ck7BwAETUDaE9AjW6tZRLlO9RGPTcBJMPjfErFpxv0cZ
gzyGglEhSa8zpS6dNCotKKznzBIoIUvfCXx3QDcpb6CvxP1oRgGvVpoCgYNogJ+Wd0GkO1dGeysg
DP0LXHXqUtNaMCz6fjaSX+VuRCGi8JiPTZbM2R9Fx5jL1h2HZYPOVpmFbgMgGjbiBMZI6sVyFzEt
StQu2c8eBPpKPNZcyHMOQW/Z+ps4ovq5eDuniEMvMtSWaXCuZxe2q69m9KVDsUURzojM0Ko8iyg7
KtUcJWKamjxbCodjLLJm7tYKn3NQ6V9LHpy65WsA/4P+imrgzpDcmXRALR6o1Ugs2y7shMKphsg9
PSED33WIWG+O14RqitUl5aRrzl5CR4k+QS2ro6JnNRdFhIA6sgYy7xpK19/BbzD7VQlB2h0QHjiv
QSlRZMWQ8bLJVdcXYIfqxkBvrhpOOzJhtPSo+nm7GerNJiwLQ/3EbmWDtFZ9fG622Ox1aYrelAJ4
gPEGEWCMWlsEd1oJGpnMUV73ZnTinGj5WpwmO9vNtr9wBehVtfeBbJrPgNV/eJXsWhAdf3ZZXLaz
YBDMUP36FqLwmfJCWodRr0JofLjtzAFRBbULAV6M6i33oYFMZNCa+MV4msB9iqnYH6pouGt+b6DJ
XLRk2qatUiy1rkjc/lmTU2j+Z0gEQrDoJwZ0/n1QelmhSZoOp2VTfmA+iaJttAx4kT/0R2AaiOEm
WNDjvOFyVJhh3YL5ChwQLx+V7iEXePQN7hPjqa2YgqG1YxFriE2Y7XoMwbHn1g7QULMTONYaEmcT
+X697oJS1tXOALzesNB0ljY0qhXfi5hOTTWaLuiVkYZPfYlWRXzvtcRAN9XoY2Tzh8s9O4/kY07T
zwaq6XfdB0ip4H2DMwOoCpSbagUMeSfRNMuBXPogdZou1ohyeE7+6uH7CWGFwPS+o+H6+WZ/LnDB
JT3VfcgYYoaYSJdwdyiRS+lnu3ReIZDSXBnyTSRqVNO3BR8436fykZL4U6iBsawM3h21scg8hs6g
YRKvqKBGi9zdKx87+dXv3pXVIc+woUFhmKcbkgAA5G37vmVwOhuN89jpPyRzaHHwsDmHQt87MfZ8
oY7ioVPvvyqG5oxkxmbMDeHRk6FMydDlQ5yBZVFBwMGvp+qtyDGAzqXSDVd4Gwah/itpUJOKb24a
9/n8k2s7spJJsym7kwHyMCgddQkQ6NjnUwuIsLCcawUpQ/YZdxNB6q9x5jHSIX/0C7jlMuwW7vHa
2hszQw6wQwAGIhINn1EWAPZaV4aKDlWQlUp0rqyk09+0wFKRm6Yzamv1+l20qG/NFMxLNvBgmT9A
ZZQ4OSAYDsV18osLFTwVg4Ixw3zj8sxl5+z+xKfa7sVpLdjZjXvDf3fxkLBAzR3ZwQKikLKmOY2z
Zu3Nil3y8f3gJ0Nji6r6t8fNo9AJmFBAi++1VDHekyjNF7TCd4qfFhJLJprMiQjZU/Ti3h5HOeEd
gg0Y9xCBfhPgwtMLzSbbKdD8ekIWZ2QEFRG/MY/QMaIIwgc63FvaVRkvbzjTxocyxz9q74V7qamc
PkDHXJy8zRaCQIC2+7+hvD08W+E1aAP8xDAtvnbvXdnz5G/Cjs0S0aY5sGIhepCDR4sOu1BCtSFt
AGwodUnlOiTJVssbwhrt0CHyUjfqxBIY6HfVgt/Ze3npqz3kddM9GzA/lmAlgdrbHVGgNbmhhqrW
KHuq1qUWoe6zGkar9kwMs2YNYzWbBM/6W6oAp1iEna06CINILvo1DEY3RiwZpWfE3woyFodJ4NF5
DP2HFobxGnFFP9VQpSUMPh/8lC9aWCbCnlJW8R/XzIQEFYVlbxYakcuOfeS+tAVR0c8t3eudJ3fi
x4MsuwexPx7qoPE+Nm6YKrYJsRmDSb5cpyy+3NnNn4EeQ8ezb2MpzaXpmvgrVxYUfxqInKWmt5rh
ZQ3/GnBjEeoUmlf5ng6XvbNzfBbLSu/MIYl79Cd4OsUmr2CBp5O6T2DrbJ7zMZNyuJ9L81zwyHxH
dD3bgOyqg/m84W1vS9o+UOgO1mxK4M6eCvmilqSMqC0ql4njcRNkQsl/YqXiJPOYgBG46uGMxSpr
S3fWd0TVJSuFLJhuRpQYwooK0L8yAVWNlm9Uqc+jzOZ2PyMxflSkgsrz4LkmuvQNXi5WzOVaT+C3
QtqlG76EZK8/kz8tjp7Rr6HcPihMQPUkCJ1lR+UJHv3r/im8OZQz5tb+hIJfSGrT/yi569Xhu+QI
nreuaWLy2N+1D9VcLlwlXXptbmFB9A3XO+v9h/OEMiRIxEujHUPAg68TGWwKiJumJusd6MiTOkyO
tAr8/MgRdvucUtf7l+uWr6erXGrukyrIU5Pv/q0mMpFFddSTkzU+2XRzJ+29dosaziXdtDFD3a3V
mV14SyVyqyTNvszH82xwy2FL2jAEJiQFoN9DaY5HRiZC6icSEjyZP+Vwt/+dVTL3I0jzfve2NUir
J69sXs7kmGVhYFlPl6ODoQzSmfjE1teJ9AhTsTNQ3k2kPmINwe4t3LF+/W+yLzESOdmNnZNtgBEO
F66aMay3NxFOabYoxLxrYe9erjYx9JkJzutGETkZsF16At5HBp+gefmjdX46T1kp0Zvxi0eMCPXr
1vEz//IB+fzCeiBftcglJUWhg+EcYqdZeTk5FRWn5kpt9vNMmZF92E0XlbxnuXsAsu5aWJBz4cCm
mNYyqf3ATttJGdzxqTrIipDKcAmywQ+LfrXkDR4PUubCIuQLdbqztSoz17PGSQ2ZahHnhg9d78yD
kpa9sq0yrru6gcMjXPdLmTA5mf0tHccDrK8tR2Uj0y0G07dZEmAJpcQPdOZe6xqzWWMnlaGKbjPr
kQfhllRkzEyAPY6iTIUyhhceKg1G4ziyEReB7Au9t+y1JQPFB/1PFbyMv0edpBTH9V5WRgsKnJLL
5/o8pUFzt2TybhYYA8tcp3knpeUj115iBEcYSxrq8104PR33D54F16Zu+MMZx7x7JlUIdVnhlPjk
LK7SURt9wFke67MfoOXg1W68nXH6s85gDq7U3La99AyaueWikHYM4HXy8BStQA4UTw9ielWs8n92
IXnL+ftOPGiOUnT2p2VaRAECfYBR8zzkXq1FE9+wZzQxqmQ+i3XzkADHK9e9E8hSxV79x4OjQUXN
BiLf3AgCCLEFRJo6lzQRWxffB8bMsDxT/Sy5CTpk7hSGX24bnJZoVsiNOwfc2+DlmVpGdbk90qf3
gFn6k+Gue28q0lRL/C/sxdigNGrtdAVc7oWbPMGmXG4Po28cS8NAMo1fgMq2hHNLmq4tlMZJqgvn
kpkmQNGpRvj2yPz+/A1yRkNOAiqytsl9CBhK7IeUNBul8Zxm17eDFvJR7DFjjr72FBBk9swuXvFM
AHDH6/ANGMuxnKxpJdHvopQhllUkcjPIUWsHccbT9KO+hwx03DAUwMxiQYssh1VySh9XoUwBZWQE
8Qq4qEMbbqEvX6SQfdVZQmkqKfpbpSWDKZ3YNdFUDwLw6+dQr+FAUolyp7KnXqdntGBkSwuNX3Y1
Wu4omDxa2zzXLGApBMB4J6eKp9WfMt76R1+HzRYFvQeClmx02lAqJ+p4MqkEJ+fRtjXxPRSzoRzD
ZbpQJeWiU0yU/OBRT3fINNh2aepIwj3T1W8PHomZcCwtZFXI8dTdcJEqSC1KNZrLGEHMYA4utGSe
n6sZNW/NCfYwmjQBwljcvGqw90TqdHOFzoEPrYZ3yBGOu310KyYTzHVS16XmZHCpoaSZkLf/xUYm
JpT7LEwlAOleN+ehPnyZzMTST14c54PI4F/jj9Iu9yx14ZDwBrc+yBqMMfsS5fR261gKJa21g1gW
TMg+PrWGJpEBt58yoBFVk16s4D84Hb7nP44MqE4IKZetAVqKIoOfSNRKg68bc5aSRkPSUvsiz67Z
6zLEtsYhYrj4yPIPWcaRhgq1XdCPfVM1tnVk8p8A39ZqtxMRH9Ril2/CWz/GIAQCD3rKbXhDc+cT
f94nKjyopOu11xjL6gagTFOdta2CLmoAZBOJXpy4A7nnVB4TSTRZ/VHp4uMu2c8WDvo77PAKb9/P
wkC1G1ZVdcbJ9XwMldTMba25RtKZ12CCW9X5Qz4/AdjM+uKHvWsaTJXVu1xALTy8JXaD9RRqxFK9
OgvXKQzYdzOeocfyh3eYLJck8FyCjNpRsCZr50ZljmQXhqZnc781PuFPpzBcVvjaBdgidPaYbKGe
NMaX7WliMYetyfTfltcS1vxvnxQR3I1AWW5Vl5pZ7ayVZP5X17JTVfdod8dA5SViajBnyuNHkDDw
P3yAtrQfFL9sLrr1wJcGiT8caFJVdJ9MKiE6N07tnMyHN+Oz4GlO8FtwnQcDpwkMSAhMO98XOQJC
G8oRW5cXsvJfmX9lSOSXYZVeRIJh9BmI4L+1k8b7Rw8HGGVupdyp09+rH0cUaTWJ0QoePakuGMz0
9WZPdyWUswjPJBF7oWfykU2rE6uZ7nc3cWRZ80SsoOTXboCacU96NzqPMYoic9S1qzeTUvbF6vVQ
+klfwoVXzvz6GnVgDL/7Z2XJu6lTObJX964Ve2h9Q3uyoaKiafgnb8lnXwJzpgBxZKTx+F6trMcD
pOw0F5o5LQpXR8rLlngdbTzbSz5WpZaRW9IdL5tUl9fTG2R4YNTCZu/4U+Let8pzOsXrXfnlRxne
8K66vz1plP+TzAnvXM9U1chbQphqP5Zs22KJNP5Dhis8H1WsTgHHgRwPzBM9LVN/QBz3y0fol9IU
SjL0fqjSx3lxya2LS0iuHvTBM0qhtCPJYiE9WQ9YpILZRwPpl14MHfo/99rUHTaLizbbgh1b2CFR
bEpope/nngVLXCamoWh4fg2RH0OT7X518/JkzAmcCorHu+LRiCOuGSmzvdg9H11T0W2m/vX0BFnK
Xu3zw1dsw4XeEjsXwUpwhDQ72avNG0JNvSOgu8lygB9gSxCcR28pYHFRfD2FbMHvxkVTgRoVuaBK
zN8ExZjJ3RTPS+FRsA4sLObaRNgE1Bqlbf6h1Sxho0gDWaxojg3FdhWztZOyU7zQBM+008lFNoV/
h8NmYUOFvJcL5Nc5/fcYgwkxqfvuX1yeIvQk2hHiYT4y85E9HBko+CgdZNqJr5d16+OGLTLOqrUd
0/pux6SySeujUgg7EHcaWBo457sIlTzw90iiHk4nQKygUvGySo/uAxy82UKbZtas/uj+3IaHCG98
/VDZIwhtCW6bKIXT7kHw4xWVYxs4kPNrNM73XfSfja16ldysjV/XjSMKMqJpDnhJYStPRs/ne7JL
E8suWpozm97Jr7EXmW9euVOET2c8x8jDnC0Qjy4Ka716u5QpVGfIc5XCiCuSdSzsgoD4QIE/ezEI
umUob/PQqJHKL1oiK8YfWMpyvSWA+CvctuIkp5OawUoBb6doMoxdrATTqQqIpJi6c1je8qUm9gV7
RdHcITbNWawpl4mLFXj18woNNtdITo7M3u3V342UGTfzBE6GZ4CLaV2xnqQanmG3yCPM5AT0okF5
3odjBDwitnvUwxJpWVsnceX0nWv5fetb3pV6oIiI91rOkMdrfzaeoYZ5K9CXUm+X2zdeskSm4H7g
X+RfJ6Z1wMYVGQKAsQ7ES8TmLnubmuHhS2w/loGYEWWtaKP+OG6xRyeh3L3e57EDLBzAYNVZsKck
dxzSJHfMt58Bb+cmFer2vsZbaVnsobP1U3YoZLE3hW4FlPBGHoRHykILaf8aoHCCd19VtHv/DJO8
NeskSBwT/9ujVmflry3BAa2FcWcaIfcZ/UNCfxjHI8TZpO5m9SfVaee8g6O73QAvpKV5vfUCoUTq
Kl9p1d+LGqmtRqaU84uOAuJMokhFYpk2mPpSx1lP+xQYHycC0BkyUsdkjGtvDoJizo8oX6o8h8T3
oAu5oWUg38Fe/GI0xH0EE93tgxRYjXlaTvS1XlaEI++BgbzP8vKA/QFHbtwK54wkjlkuZQAp0N7Z
zVHKtROYlhJ0R70ywzWEDDjsjSbz4dKyo6X4u/kQVq1JDBw+TD/L16zpA3oW0+PqONBs73jliZN5
i0q+zbEqfIsVlw/npYDjSFO1qHpaTw88UVc2/2slu9Ii8r76Iw389noDetRHKtwdJcUPh6xjrBBz
tqD5JgGRgVwHA1VQvcBcaloRuKXNkB8ee5HRqhYoW3lco/xPSI8H/hAwblaHvAslnBb4obMUvmHU
3vDytubdZx19MYW2rNFZXX/jSa+8WinuNoq/Kxj7Bgj2mYcPZsrnkEWhgKDk02XznogTArxM252e
GxKdO1vmC9Y7jN7VRJKUZIFNQDoQZCNMpHnzoKk6to+Dk8oFr+kvHH3SEx1muX4fO84KwWcVbDEZ
sHshZQP2066vtP+2GZ1Ziw/1icY1zWjBLfFl83huS35QEgTe0z4+MPEToQ6Bhl3M6SxFoKTOKqO1
bwndKI4tZAYLfjdznDpqvlFqT0Uuc2P2HzeHdWsiHwZhFeODWhqbP/gfZCcBwoXLjgBIyPXNn1Bm
ERJf2bebKxYbjWVvSrjo6bX6gHNNoAUcFSgJcJUYq1TyAa68H2eNGFcZt5KbEPLwcco8lsj/z0iW
hPkJ5jVuFIti0DifM0TJQMl2Lv4raJyauAqoJKwD0Xk/ahy05VpNlJtbIRZNg9MnkW9ZNc1A9mse
NvRHQlxX/inbUPZC04Q1AmLdjRUyneOBj/xAFwRMkRhXx91D+z0d1RSWhxnrg+dCARRr34544LiR
Kl78YXIKcEr289aSHHfWztZK+JWfv2u9xiAfGYdglM2p4WCfiraXa09DjmstukzcaFG3vgUelONl
i41KMeJxXt50aGnHtQN8vZ3VS8+7SwCiwz4wLBXZcjeHmCUe+0h8CHhq8ENDtZ7stp+xoh9kRT7x
TwmmoZPm+LgBglHizfdsrwqZP2E7emfWUxywhnKz+KJO20zSxY/AOEKWpftpNGzVNmu58U4Sia+a
5LN3TPjzVuk4vNdATaN51pwYsVu/zczBadellMKEpVt+knSk4nkvo53EiRemFwxgJb+Mil1M9J2Z
aRSUndTkaRBMecs6QMAeP8BmGN+4KZIYMj0aJ6zbGDZLbpgE6CvuODzqXGqWBXnqCigU1hivh5rS
6BJW0aSXxu6LjkYCDl2VXmteJI/YON41hy2xUvNFHfIf6hF4DCguchtwUVWPqkvGK6EAcF68m/kV
orC6Inc3LPUtfZuTaBrJRzlush6+BjBwbCimlzSJLRaveJtcn4faMZ8sdQCgo2CsvKg6N3iBLv9x
oEfLDvXWp8cSMWaBoAQZGLsDN+ylD5FahT55VBewDqBh7T1i/LBl7U7pjhlM7ZXO+EFlhIWpswff
r2I+wGhGUdmn+t84C0Z4YwXVUSqhWBy04/ZN4+bY9Ua2Z2XW6aE9m0S8KZifO+o12RsGTsjU3q1u
gJR4QNWOPxQpn8B/pe4rwOdDdFgTioWK7yLdfRF92bkKgDkO4dntpEQOh5PCEC8PpIG4Re2Y8n3q
bjL1bve9q1I/gqelBhvmRBb/BG2W7yKqbwKpESD+99viAKv4G4dZstjR394HSODBjJQbrb1rEaQA
iWsPzKLg1Yn9NUrYoze3wyR1LqPtnmHdiynpi3rlK95HgMDZ8ZU/MjBHapUs4xYT+LRW3Ko5qnwR
3Bhr4FF1KSb1XcuLmz7mZytduLdZBhjqTAibRQNsg63tXk7Vm6qezqn6OgoZNugvEM1/ha/OQv5B
FxoiX3BbbW3C4anDxdkmLqG5Swx87bBHJmErqISm1e8vrmuJB/aJDvrOnw3Ko4QNfZ/xskHNfA6+
M7kvmch6nFb+oCvxRuyW4dAnWHj1/8x2G5LjqrQhIWoRhkLSMFUncYP2Bq2YMH0RYl63B04sNAAs
IESKoZUb3guKIpTZDE1RGvWzcfJG33PM9reEqIOpCJ9iVoOB8/TxSYRl6YgA4QSerRs37qLQx0SB
7ozl8EeiHwNGCA7uAMLCb6P/CUIVDSeyxsJQbsGwCLwLBi/CzjUfuBpxQdUX780pDWvaEapWygOf
fgko8zvvOvOX9m7v2WFcnlreBesofkRgK33IkCWB9hqke6+pcUdp23KX3jjWhaL7Y/vS+UyqB6cM
PTRMaPQtVtoH7TFXQ8b/4kUZAeci1bnCTcW0aDmJRF2POUgcxL58jMKxhnGo7Xkc0XUrkYlzZKgj
I4Yez0CtGBUNV4aBZkkTSq0TCcgkuAs/+EVd474aAKREc0hFdiyZM2VBBCDyIwWRU4AHOJf0GQmU
HiUKIwqN6TlYiL+CN2/4Jnk72N0JEFpQhsmswzYgb53uyJAqopaz1Yp/wjK6KY/hgg3j4WKohWD/
xHMjd7VmxJjBdSlEZwsYIgxMvPYZ4Syh9UcdJNnEBmtHiW9OSg0YxioTvUciZNMwhvRGJTh3jSHI
yMD/TfohW4HJFhvcHms6YVJkxP6+pRwEbpRpW55oc0kw0VAGZIZ7BP1XYzOQ8SN+qe0dyKIom6XT
QArjXe8hyC6ASwUI4G9OLK9/HqTWwSnudnSzI9nHNbaurTILbZ+vf2m+GZuCsfAvmc3bNfichufQ
wiUb7FvpsaL+OH7Z+BqKh6RrKVG697fZfN6YpofZIwjZi7wDMt+6pS948jXtlTY6uOb2MmxocIC1
Vs7ypDoOk7KvIOrlTZOupBn8WWkaIKae5L3n3TH3+URFu+lV6THjgQzHZo7KzZ8RHla7/qn1JHcP
8eL1ZdpVzbDG8O/QMXSlZU9K3CBsQsDy8kTlQrXW+xn4weEeihBUDd6oe6bgLhhXKDi9VNV7vxoQ
xbgoEGibzu63ic9naISpTjege324+Tt/rxu/qseQqqrJQRC/tEliJlPaAJEeCwqVBLDZA8j/TbUu
mPRc5CMugjVFYce0+GiJ+13nosn6zSzA5dWerpG4sYYKu3TRBYt2caQNPFgS78eazQP67Ng2Gful
2qR8quTxZYKHDrgEra1SRQciRs5fxPi6PHhKEkW4IgKp/znzlLcfZX3YlxVLOTYwTZ8JHddK+mr6
mQAy3o2PQJm0oPVEBxXojaPbqr4PtqIgjP53dHu2QgtN/p1vhgD4fv245dK/ISseJRou9AyhI75F
Y4zCsg4PpoZxxdZGmqaDFP6tzbz+z5YfYJ8QEqBLB3pqvVmoSsp0SpulNAXK13EmXdduDaEkdany
TOz1KzzZRumCGtzRxVYLNNcuPX9PQvjC8DChWPZqL0TtPoG9kjZcKzYSQP8KtwByw8nRmkvt/COv
HrHfD5OVXRnUauXZpTsRAyieCEY3JmI8vXGDIj77lUIEtQ8Ykji3knnh1qqvBss7HUZfBJxlILna
mRoDu453e2b/LbQrdIl1uMO9HH2hffDfDxG5xMg5GI0xMiKhwj2FxQhtyfQ2LutyQdwiOdgbO9Px
6dRt4BtUQM5KIV1jFRX3vEfwvKrTdnX2YF8Qg+eJrFSm0MvzFW9UfLg6bFdO/AlelO0TG9otWJgQ
mOovyM21RPPbrQeUYEbRQ6xFsdmP/TNEUItlc2ZQAlVgmWLdk0UxIN31FEtOg5JGT8TWAVXsGmfu
SX0BoOxBK0LXB0EyrPQHKn6Y9LG/0kDGceEJSgmm4/OvMrMLhIRLKVRZ5IJvDwOn4GRMjUKaK7R5
j4I+WN4Iqe/iplsI+62cAE5ufP2f7IhcEh3oC10zjZD01rnAVYvjgIMBXTSJLdhjH6mrgex3sKso
7PBambQaGiK3hbUohBR0x8xoq90J+pwD+rXItVKdKV4khBvjOn9IiZ3Ye09FFXGOfyHO10v7o898
cWKzFxUaG5Jd/xnzTFXbGuqhWecq1JQYCd4AtETtlCxQ01ig86ssejtHIZtSHO4aTnF97oeubrzb
f+tF872pvlqBhcxecPzFpHtynyE+H39kVTmJZG4wzWouFfz7raJjoomkL9+UejzQtAeTM3NiIG43
q7+nkMQ1qeEyacgJSUn3/3KoFn/e0X26XmxTccU4aPPEGnFbU2+NpyrdTfYy4/c07vJrE1m4W8kf
+VSAt4O31k49d1yUC+u7j2YwzhMPlXwIIM+buS8dVHS64INIBgIoP9z8/mG1DVjxd0UolYuVBIsM
9OG+oPeJ9o9USAAAmWOv0Z4fNk120YPKzMpyVR0sjRECnfdMu9sS4kdnmujiANEXpdR+Xgm3h8vd
Q5I3+u3ocOaePMTk//PBRrZKhRwqt4YAjpxraDhFat5Gf8l2tWX/61Qt3YRSFEIpQbMR4CmOvamP
iufJT0Ea04y8Mqc9tnXKLrRQo311pWgJlWYGDcJnRK7VCNyzRPt7vFp/0gyynpJ/P3sPbkNulyb4
7BmP76RWCcxnlNI6apXtxUbuV7aFNLHSrp79YuHh8imPKvqBviCwjirtXTS4Ww02m0GSfMKNQ095
6eVw4dQI7JtfTJd7QSpw5R9LJCVYcjwZelM4pU96CQHPMyaxeEIELszbNj2Z9sqrpsAYrp5oETeD
QkoMOgosvfpfF1GlWZPgcvdHYkWUdwvkNKlq/V2a8bk8uI9n+Wd8rONoP37QMHMjJBe+boLIdnqf
AyEedMxNphuSPA+w+2TYCAp8ar8xrjXh0i0cbWRmdCVfRfJ7Q2YjXf9bjOqk9oTR8XZqxiuH1eNB
VSuit4nA353t6dihnk2CsdVSteuf9NCYdQW3m4vxQQeRWeefgKIqbAZ6kM3iwetFvEAnMnpml6ch
Cf+N2stsR5lGoP+fIt//UVpiunoJ9O1EJmKz9B4CmHcCxdB/8vW9lHxX8cU0q6JEU7D5yEZrO4zD
kZqFlhP2u5MsXJJ8QC8ZPjU7v+NccfGAeQitNYD193B/9oDc/+cNYoqVFUIiffomKb3thOHBL9VX
xCf4TN+aeyCDBlnqNym6m22ZKsAeOc7nTbmrHcfRh3ggVL8Dn5e5Tx5T3/V4q9VFtBFr/8p6Mo6y
Ls6DqnQ+PMCDd/GDKoJOXb/goKbPd5Te7pCxY0l2nxVuZqNKEhiodQ+WMa+Xy3Y8qPslsfOudNVH
HJAHrBdLfaEmVQi7H2OX/nYZOcpczcZZ8Ze/z1Vl4kR/mp0qc34LBQOsFSYYmkysSH46gihNuW5E
H1p9BKZyDsEm6p8IRfq0b9z0e0M5rl0Myv+XLNsTtm+G6TWg9lgEkD7OedSNC5a/yzu9xUenTmxk
1AczRgP8jNT3sxgEcx+Ig+pksaxWms1whaYhqLqMbPl6LbpsN7pJXVFVe/ILpsGMyQJ6rClJsCYu
k4YKwuATFW4hdUyBUF5SBkU9Rj5QzJzvDicNmilxSOwC+48Q8+0dIpsOpLSfuO2gDz0/y9M9DwdK
j+f4mgLo3nxapkw/VkkQ9khpDzJ/S4QA7VnGPLClN2jDHyRisxeKnaTWSuXjoR6r89EG+kyIWzWr
JD74wjDdjcvJqoiDZ9Ael2Iwlb+L7aUOH8shFISYa3PXZHra+naRIqC6mVaK4NbWRB9QlCdTnRSF
99AmLE7N4QJ3Xzfl0+01G8hu4/zBUM1iw3KCnuEUd51HOt72ijGRpWoQ7xEfPpIbwXq/56hyPDYP
p1G7po7H68kB8MTtIfBtPi/KoCHfwK/x1malyg55MDiOe2UhyuJoY0we94tsIYSOGnmG9GqPcFPX
wO7ITNwlvUAfzdNvQZeKCiqu4qX8w1RDlY7Ev2aCch7W6OkSM0YZXK+V84h9ZMpjsYXeUWY44/zu
yef8mKrQUkTVvZl6nUjDuaHsUeuYB2Vu9HHffE7VD5D6jP7yovENIVd5rS7leTVwZZVYh0pdzBYh
SGeuwPql6LVrzc6+Cj45GlwWCcFMa5Mp80kG44HOZ252ia3fJp1FIi1+9Fut0N2t8JQpVc4tUEky
TdSL/C+aS3ANlUMPYGsQ4VrQRuuWPwnIW5R37Jco6aMoAdxNnuvAsdljUDFhDvBdvDOO9jJMUV+S
I/HHT8ZVTQ0UDf5CZDZu5byzShglc17JW0A89dzH0NG7qiJwLTYVk2fgqDzANnkF+L2u7n0M0uQ2
b/ucrbvaMLsP2H/P8/lYckzfUARe/+AAmpBA2EvUWcTQdd1DGiLZPaF8j2rYhS1piuvY4m1LxF+q
Hq5y+DhCYlPPQb2189b5CoSAvsMbiR0mrgOdqdmSxaJf8O6HbutTdIwmNw25PxxDDLkUPJNgIcwF
Uw9aAuUfaHwGEBXNDFmC/WbLTbz3yJ1vd7l8zGTdLhTGdHXa+gtQqmUd0XZT9EaddkZKjBUZ77Jg
E4PyF8jZwxdZjXgOutzB7xSEUEZlPyA9K0TfYRkb8RwRYFN4Ky28DKH2fpvKK1cdr2F/XcB6UZVy
Zz5IHDfCbBkNGelQtJwrDHJKkCKQ/4VsRY5KlPWmj/AzNDSiUu19hIE0LGo915F7U1X/w/i+XfZo
8ALY38Hw+Jw52r5xX47RJ7U4o+UsdrmSj7S1Ftu66BaCYHSi334bI4Jg/feRVxviNdrhpWn+OV4v
Ng8cOb4pSQhJRAk1cvvlidcVIIeAaZJL9T1uGV6d7b4C2DkmgwX3ksPIXg0RTngn43Wg/oFSgqHY
UmS6FgZN8u3RGTovRhH+D81DoEWMg0tkO7Z/5H9ZUshSLPM9/Eyv2XKrPqDqFZ06RMrLY0K9dZUv
dkZHcdRRiCYmGQCNLSxx/SK8MGBfPdxgMiUjf96KM4LR/Ibl3gN70dpS7e7NXsWxquR1Byzfnmy5
EBU4FvCypom1uMVRlwMmhcCSw5B/5cFc2hR1ICLUJ435cJl/RZkqYj+oN6Nmv5TrB0OmwbJwv71p
ig22xPxABkZTGcCUyl2MGKLkvr3fj80/Fdgm9nx5A2nA4k2mdT1I+nQ+QQByl83f0SwQIh4+6qMy
hgy77AzSdZg3so4QsfkxI4HLcau922Zra6dqEvBl0GN+D73fnMDBGxRM96ZapqbsodSf6bnQFV9j
KrcbKNcCcjimmt7uoGKyjaa0luzMd1REZQv1U2A10zh3FpxCy5/j5xXnwGVP6k+8UBhBptjfEa33
87tWm7LEXeJJUnW/46zBqFUy+P+kCabO56Sn07g0ZjHyy/GMJoyeYfqY0U3exT5BNG/N3InGoyY1
m6G8jHO7jTsZqPurg3m/cwji7bgwlDfNyN3eopvqcJsbcKTT0iw8vIntuNT2aYcGO983AjBvlCaY
wXghcNIEYT3alSWOWa+zSkYWoAuDxFRlHp0r/2o4P1ihDPpYx0PcZXu7IxtmcnBTV9CGxNbwFs/0
CNkpsSUe6hvB8tqYOMeg7zyxQOSN/hOrEH8IsI5ydhx3ME54YlZmd0Ikk0cInkwbCFqDzwyQrKmy
Yqvjbuul1qYyR4CRFwQ161u8K948GFpX2//2D/lI41W2XhjL1ZtYQ9L8HsP3oyUyt6xoJ8VXuhcE
hqDVGBHDUBogbFstLz6d//70oHu2uuAW6Ad+tVWteKRjWuseDHyZUhMHUsby15JEONobFOSHyOYr
tZqIwLqUST+65DNzrKG1E5PO+Ci0ZR13roo++Q0pZX9o0Evepmzxsw3tyaDoOau1b0Gc4d53pKH5
qocR/iNbR6G0/J7qZktXXJpN0phn18c/L9890jcpqQQ64sJCoGCoR5hOc+jblnJ1JI84WqM92ZLa
xl3wQ096hS3edpe6oxxxhaFwT6uyRbzX1spmuv67FxMEZsfhbAOaA6eHigp2MmfVZ2V1ItcaJe0Z
sKlj7jwavqh77D5+TFaPYNa1J224Lde6/n5/lQr0mzq0OVVXtSxb9R9jtXCBl7kFVnhrTMTNZiWQ
pTM1dBe9W7t8mSV2YCU3f5eK72ObszPjWwLJyQqqEtbiO3CEaHm6bDJKAHU73WW8tsVbUJBrawWF
A2YduWEfBzjXh1x3zONGhAq4Z9aZ7cmQiclno0GZzC7VIYFyGXuHTaJ2U23zByep2TCatZDWBYux
91BbiDh+nm89rPb9VfepPiT9dmc1CqXII7QSndKhquSiqLR4v48G5EKZgCrZ9ra1BqnXOnJB4ENT
STFqKZrdtI0DOgqY5LZLuwoeyDjh9XDwPeDRaZqyHwXjpG9LUq9TrkIPyAJFVz3agK7QbgOsP9/i
sBgkZ1pdxWtikbkuL2xFaYBr7SdRczZOa5Zrqhl5rhLYIWq6rU/QqfGq3Nhd9SpWBKrqQVLedCzT
HD37HSrWIVnmqW0X9VmknBVaRsutJi9YW+4RG5Z02PusgMmn9wmltJJM/phXVXJt9GGG+KwfFReT
wRw0NZGaJuI/CyNuXBdy1M8blYydmg6E74Xf5QcUhwBWP7bk5eyy9mAuUnyOB5vTGqTInBmKdjTy
l4RJ0MUmM7J+z7I5/R7AIAbOgDBjxQjfQBdwgkvlFsLckQ7KX6DEw+gHi7wbkuEfrQHo6gxFllUP
eTs0OnJ38ABreDH0oiconQbhN0YoF8v84EOJ+IZa4iIJT109WB/fP7OZlc2SCWMWXKHlWpVXHhDO
4qgjjJsBHt/rhgms8bF8cQb4iMn+PEo5qZyat21CAri9NcDAkHtZNmS2xnYf/e43nC8+ATc5FBlh
Ztc0+YKNGsX3JxMT5Uv2eCu3b4f5TsN/K64tIcwLC8EDpj9Zt95fjbpp0HdE9AF4Y3x5lRHLk0Dt
Qwtr3MH9BVWn9I3a0uCQ6XFzoqg1QNdPa5xmxEb5lzfFfwwo2mjUby88p2bQje5zWstBMbEYVZv5
M/INFjxdBFAxSSvNofjdKq6pz2ZWYCL3CpD/YQXzTAoxmqYp5JIfAvVH6Z8knggaOu6P+TQnuIH3
0kNrEJMFi0W9SQSRQqVqAhsBW+lwIE6i0D3RgVg5V4OiPPpggwfEAPB1V83m4LbqAViwbKr6kLNy
l0rxY1Dg9ChEu5FEhdrs6jdehmTK6ABOdKZuFONGYKUwQb/gL+sI+4+cY3JZVQx0ns/3BQim7yhw
sworqaXlP2SlgCVpO5sTutbnamQz6tGyYq4AOmJheVkAASYEZRX12F+9fL3Rz0msXEyX+ZDpN1hY
c++HIu95gozo9SyyWyBl02C7XD0jm1bXnIGcz0Dt74igDEWUBSFZZ/M0wlMXdWp/lzkZr7O5SgDv
V4q4lj3wdBLqkG4jAL4BWsUlTpw5GhoHyX25VB6Y5ykxTXaizt0EqNmahS1Ur28/NDFNg9TNUoxO
JZu3ggxKT9EjJPSQPA3FP2L+kYZshtYERlZ0wd5yma/ClvMQJRQUD4M6zRNQYNUqe66WhP5kxfOO
Oe90QA2ochlqgDLiNVTyP1gyqK0ONilPRt2oHVXH297LSKSAMNRdhiDIIfCd/pQP93qjuro/VOtE
dw+L/Wt0y3+vxdnpg/UQtASCM3FtqP7yBJZdrA6yjT1DJKhWDlBGkKZOf7r9A9v1qqDlfzfJsTy+
p9hikP2OkxKovEjoFwtoe4sTaCo+5bMobj5NNroHV42dxsS7lEHCmusB/eCIO7fI5TpP4Xx5rsUY
iiF5cdtUh8G7/dsSwg8VPKLccFJzN0XQmG6xsw20Ct3qYpFwTdraLVB7tCjt6AjuZtU8N+r85Sro
+eOTQFbe9UKynSK1RyPYFZGURlKCZnlsr1rEuZ3HmXWxYa5MSXPmnzsciY+ZXfCh3TAGssWf/3Ht
9ETS3WJE1Cikp0P2B46jjvnxgbUyp/Fdap1C5BSZ/XDpDCE6KqSKqNDbrmChTAVWfRZjmdwLN93Y
sOCDBSk24GRNOioroxi6V8bLExGNKN+SWdI+EXNMOoueozZn6vqjtQ5dQ5JDOrYGS9nd4T3e4GZj
+cDIn+rxo1eRi7/306g0qgxHCdIFu/EI7kAHTK8SzLQxwjwKeWylq3v/rzQpO4IC7f3BfvP6S1/e
n3ubP7/3b/0ZM/TzSYNU/aQEC6VLGwTaaguOWI2WKyGEPhMtHeBiCGU+oiTuTheTB1tdfs388ijq
EAIcjDaSwt45dLdKtr1T5TdJY3Flx2tpSysisfvl+TUYUcGI69debcQeACbl6ygVaF0ESqQXLESB
0cezZ+wFL2yslE/brRRYZEHhWfHMO2PkHT3N4QZajuREaoEFvzRuHfm5pKpOPBzgY7aJe8FkCREP
cYH0US+3C+yi0hbit1uj6hWg2vx/8ZcXA70+5kiNpvsSHatwys1aktW4VWpMhLJNIYaEauAMXSde
DciRkSKZn3hY8AKOtbSX9+w0Vimwk1/9k//+jvCAjlCgalfzuynNreFOB1h5aCPEeZus0f/Uv1S+
pcj9wA+xUaKcjZl+8r+Zbq8ph88C2TKbIViDNIqxKe9Yc+wK+k6dG+ofPdAqZxMvG1QrQf3w9LR1
CJBI66seTyiBlvzT2krX6VvUjEABrXPSzD9xE4UTa1OkM9gNxA7MlTx0VbWwqaKfLjMYfXQS9CiZ
5J7tRC/cuFKkjW9xkN7ZFMWhfcrh9zph2JL45xYBW7m5WMk/xuQWpo4T53B/Ozy9nG7LggkSJObu
hDK4KwzdjmJR5HM/4z12up/V1LI0p7e8W0DmzNKt8JzbANlQAxLBvtk8g8mVsKAsM7r4Tas931Fi
4qmHXAeyanPiNoPQnryAr7rk0gE3L3jAU4uxcN6vPYpA4MR+mWjUKn0Wck2TXAEuDvus/ZCUwBbU
p6l7oST4J3eUuEmRT2Dw/XUauQEP4M61Hzm2Wa0jm2Enhz32k3oNr66o5zTKp/W79ieUo9J+IpDX
3neHXAbesH/O26C25MhIKpswA4c4RARKhj0S6kkwVw+MNxJXXK5gUGJxeELHB1LHcby/w7uv9Tr4
BhTsa96tn1VnRcFtWU7cHVuiJyk8OUUSeGj4y2li0vxLLSkoaQLM9rLrtV0rARj2jij6tajhTnDa
kKIPSxIMP/Cf2RGDE2mf/UNPEX1+rWe1C/xGqhQk+lMwFuRxMkjrSd9oscH1PZziK6Wf4e75zlHO
psg/1OkTTDZsNTIWovfePW0VKubH2s6WpScimsYJMdD59a/tMkxHq0V8MUq/Ny89USnRm5NQRLa9
xseOMwLbs6NbddfVw5lK1AlHEfgaVM9G/lIhffgRHk4WV8NRNxSx7okz6t/QAtRmjBoqN8cd6QoW
URZblInPt0Wri3nUZh0p9OsAyvgt0OT7ig7Bn+LjulpjXyhtmNq5WJ/x+c9/T0g6hKeQa3/FQ09H
CrXATgEwRK627/rBFrJ7SuUV2F9Kk5z4t4TWqCGbSCmuA1Dt5lFqyEDXSPmFDS9hGZNqzL+td5f1
jOA0grpQg5UBvG1a2PzOkwo3FNK4BnolF75uz7rgAgFvQypTHfYF/qDlV8E/eh6+xh6Sr2rh4qSU
IAxmkg5LKA53+Xh191OqOl52/AvwnXGVhmIKRBWfAxXj6IA3RdAOaqFKHpq0nUWHWJBxLm/lYXGT
gCTCAJhAvyFkiM0uNWTTgo0BA2FTU4QxL4nkMFL8oTgd+M5xS9HYSTkDREdX0B4sfiRdO7fN6csK
WxuZi7V5nHw4t7yJ5X3zPkworuwtSrQH6mSaBigQ236W+qp1ADYYlkpf3e/8z3701FzQnMXPDZ3b
u2Jwar/ZuxQY+ZDYYyVHMpz6H3JjQalqRbHXGFgRaT4KwMgoWhbCMN8SeQNNQa0ZibiY9Nfk5NNR
AiW7uNlvg8eXlA6PjV558HIbfL3SZmDPeX/s2CaJzcsvos50qpYFXMNWtMD2uL4FmZ+MPd/i7DTe
s2VnnqgLlADEZ0YUyml4k3f2wHa/be2a/Cq5aKVFktZHtUx49jyIy4+kKyYRfIV6bcdCNj8OneMK
1PlWdkAl0yEMRzrDDM4r41oAFG/Sd+QesjDqksL56Yfg70zE/9DhvbGkOWsanAm9r+qZzPClyVZm
XXvs8Sq/N7LUIjQY631wzQFx0m9F6MsDjQ/iH7ceqbnsvzneHdw3VbXIUec+F7JDFtQek5I0T+bV
QmTB/6zsnHChZOGRbFkYPW+yFQy/Qtnm3eEplzAN23FHwvPbC/TVhL9XNQWq3VOhTlXJKxkYk3PH
rrRk6f6Q2v0GK+vSWkeRFacGoTsT0pkvQRNkWUhtsF1TA5CVxmkHw9HCohmSJXbx/4b5XG+CcyDW
IZUKtUV0o3GqnyWCnNfHf97ht0GxVZzuXMoYVPwZFomMaiktabjo34v3tfs1sOL3f5OqweN9pn5C
gFeKFLa2MU0tjA2YdUHMEIpjdS3rDgRdK6fMf2fqyMVyt5XYJVq8c+TFuRKud0GQ8PsUwBs+4Grw
mQ7HOwm9z/Zx6HZRyxScsdiyokRhYQFyCnAxzOjVwcyJ38LJHKi+HQqHfPLtfFLOaXxza1Ai9dSl
/WoBVp6KKLbLWenoZvqj97c5knJepPWPLOJGrDO46w+XvJYI+p/ShsXxOalcnyhwko37EOsx2duz
eEY9e1EE77CVNPQYVZdFD2aYo3F7byjb6worGcO/Zwgxj71G8rlgJOcrVHq9j89PJU0q34ZYLFlK
BH0Ie6r+I0rqVwJY8szAZ4Ups6+nTgd6dBKriwbfjDwyiKdkvx7vQeXvM2UkW+tE8uPq3n8M5pzL
l09ddaq8i6HYIwFhYYDp/J5MpA8zovx1iTuey3olSWD/pN5Sg67H7LmfEinLJ7+0YwRpnzp2bAX4
F8V6Lj3QFdIJEd8ajNmvTqx8W1fFmUzUYQBv3k5hE5RsY3a+51zaRfEOJ2PHk8ALDFfIy6y/TBnR
OA2Ett91lyBiLbBUoPUDaAEFWR7YVZpdTymmbjZG3UOYp0Vt09R76lPLz146VSEUDUm7nhzElEcQ
7BljRd0hi4q3jGjTnqSXzT0nPw1SQr2pfDce5xxHQaXRShgVvYzHlFHbBqx4EbsZkzEnSou2XluJ
x61AMOOkkgJPqiJgn1idPDu87m1eVybExNQunQb9V8hRJPs7sBfltd3wYLsIzOQVTKKa+i0aGrkk
by9pjNKpmI6JOlzcU8INLJACQNhHaCjmzKlshap0I1oEsrMwwlXW9cU6v+ete4GxJvl3zfQvdN2G
8KbcYiXRKFWbExsqKDirkK/+sJiR01HjjKofkQFqfxl1u977hhXx6vOeKuMnpN+NBPk7WKRl2cuw
ycXWv2IVxlW3rtjuCadeWNw/4give7b8itJj6wThtVq23Z8N3mQbSGQpm2KJRx4dwnI+outMvAYt
++HXgCbdETBOoVFmi9h9IPi/tVQekvuJl1T6BO5nl1zm+sipMc3mn/V3hIhKpKa0CgE7g0LnaEe5
QkQUhyg6IX0qmQ/FIYFF2bW0CK8kw/UCp6EWXw1o6ARiGDm7l8URdknPMi/LXAyPdVIC3hvDq6HC
e3wXvelQq6T03pm6lPHdX3sOKnrXdhn2Zj2s/p4MgTDqu6lQymspPbQx+FFB+WG0PgRHjdCrEfUt
SG/04E5Tre+skYdPxDi9pFV2TCg70M2kq2lT4Fh7X6+hbIbFVsElG9eJZOxv8tLmPBzmIIARBjIz
Dz6TQPkWAOnErHtG+tN/AcHmbe0vZxxpxgXAnsmbDk9+Rj5yPvxRzwRIdVT6Xo1ssdjwUh6ZKepO
xjnIuJZhfd+sATKCTiug05K0eisEJmRi7XO4lZOt+DoqmOlfU8PY55G09A3ZZxZrUy/GvojL0OTd
evR6t/riMq40J/tPsiSnRTxilO/Yb7eMM7h46M1wz9l5XjI0PMpb3KCT9YHaG/PXei8yncNIFQXI
Z9sR6OfpPBq6YEdqu38MhYiUAy6yjXYCVOSv8uQ1NX+KGwbrjUf8YoBODdQty5C4lSgWj7KclESQ
qaVkEAIxyagblkhBxEaaBLBUR+uXl1RE/QY01VH4XyxO27u5kStHw0Dtcf8avuj4ZC4WxOcAZAhN
N3eTqbKrPDPq1spMQX9FxbndPaBto7Yk7yxwqJ9oB1taPs66ni7DgThuvnEEUyRm40O9X4/0MY/Z
vfya4o8gIIPKX0LdWFwGi2JC4SGrfbK7J3Q3SIv0xPDLKgy+E8Mn4k6SgY7LyJJyCOO9ynvwi42t
kjmR44ypMppJ+im1AIIrrYDdVgEHuBDpW7LHd835l6+2KKFf4JToMjVGdb77nfsqplwdMb6f6cOh
UI/IE4Q60APBGz0eN1MO5SMKaVr6lfut/gzBNwC1K0gNuVn/mxoimxNvNJp5vOFV3DBNSbey2FGP
k73OmWJkiQ2ALLKm3OTvrujoumNaE7eIeN8EdQ4oSDKvu19y9OuxxgMHgpLGJ4j3p3Pj/e2RFQgV
QAk2Wr7f29CCTpbnUxiPACXXOEc9Im/GpSMwWVD+B4Std+cOirPCA7yQTvspz/bkin9y9KPWRpLX
nrEUovf5N1bGVXmFsxAVc7GOOrAqwiyp2i8YEz1I4Prt1yoW0QCOkf+6gwy9PKHmem3m2lSlJOJ5
sXTaK7NfFZDN8+iIVWQBr33rnb10aiSb2t1l8fFbd+2MObn6T+tKYmwxAp7IET1Aq3O3TAwxhWd1
lebI/AchokisXRiLbJdr3OgFnNM+wqK1oN+NxhcJgfl1DiT6bMn6/0CwwKkXZJfQ6gdsdsiYTUmG
sbEr6NDlki4Z1Va4UCxIac89TNLx8R+5qGrplGUeRj8t65AZX0mpZU9TCKXHMk3+sXRwsIt2YWmO
BB0obS5o4UloCyUmRbxEe11hv2I6QzvoeQap6KkVkgJH45cAOfCvraUTAOIhduXVNKkJ1tW1DpFN
jt/ssCH5tNvfqcWh0ipFGOpNbxngzKFRsUx9QQUkv2E+1fXUMO5Ui5IZRPt3LNzAiwfl2wXIUBVr
KJnuzFqp1WkSauZq2uHTFYFVWzXr3P9q8Apd03pbUxGC4PUrmwaIBah4PVCavLYPf4FaJiUrYaR/
bk9ozN5q5JcxAuH6o3xV+0YLeUOrFG/8FGIWzIiktFy5pNRYphNYN+Jxj3u9S+fOadRZmJ7PMItu
anS/aR8UANscc+4OztU9pj9uwICRnl9jLjBZVz0IzJM1pezuPeRNjmVEUKJZAyQcohznbJZw9E++
+sYhZrAVFKKMK6kiagv9mUlzkpbH0JMrxPkjQS6o2pnn2DnJF3nGw9rh5mhfIS7Iw1TsAYqj7wM/
ZuXu1M9+4HGRi2Q9QbKsf1EhSA+lshLBBqYtMVLVOo1m5e0YUYmTQq67Mb8HeMKairj3PXLEMUS+
z8TFH9CmaX79bSQrPuRW2//JET1AHIbVdyL5K8YLci9pM+S7VLHbNjQjNsqgKhmxgF5HCoT13Jzs
ROod9qGFRP+I24ta2+ASIwUfYW4L6ku59/B3dyeYaBzh41nLjdJ4Rf5xqxfPVZqtkFZoVUu0dRUh
wbDzYBof0g0WhY3aBrQfUpzbNiUQXM/vcqZ8787SHeTLSyZY2nSMCyylhQiPALgkrJf8G/pR3Fnd
BDTPWgUA4g/IUlBNwWTCDLt+Vaeaw/e0khpF5iKIEp98ksA5aoeNil7z2NqpWuah6T5WfcVWcDN+
qB0esZEZTWLspDOltUY47RiCym0WrIMaL8pe070ehb90lSDpPNpL/cRdjP+of4F1wvoXMomHmErW
6tq8CeTXeJpAx+ZKdOlCSu9cEro4cIfdqUIP70m3johIKq8TNiqv/RqqK7T5AKG0YtdYxT79OVKx
WLu3wkiA/MQmowzybmSU5zl6eNF/x2/7R3Re9ei4363Dxukpr+0MSjQ8sCU9E3G7vy+SaDavquEA
PMOLklKYOsAsoNFWKmJaW+iJGzk8fO67iC3ZR+IIwUgpWxagILBpHyJOU4kt/IC2IcACtDwPT6uc
SWyBCGMmwopQfiSrALnz1UmuZlhauEZkBsbn4RLkoVzxzZRrDrJKs4xUklYTv1Y5pjdi4PgfcVL0
83cSNJ8/LKmtglIcbnlnFgQpAGawsB0T1iRUowyxQWlLIC/RXNYFPk9fJvx7bnf/dqfhkLoNfr+u
QNdXrb7lsoWuinK7EbwmGJ1Ect+0OjHFMDNDzF/MEefnQQ2oZdgLAc/4BJAhwQlkJXZITEyztmFk
S2yn85kem1UG0syr9r2eTv4eNbr3arM27f1imH8AIBnOFQRxnRtqNRNX+ZdX/PyNx078rlmoVC4i
/UlvI3HyVFQDjrCIBp4o/R+N8UsZ0f0INBVABmXEPpMyreIBQGL9fcqVX0Sblv2DzAcVCYqeg2UP
9j9LyrBR54uTWBPUTXdBtxoEefr84zLzN2fHCM3Zp+AWgxxP0b6MG+8sA09GIYJgT1Z89SnzN1Nv
yehWXJhedqw2IIuuZqqWYwI4jFM5JzX6GHkzLUtWq5ElSX8P0jAIj7ZmbZbUSYX4jHa5ZtX6Vffl
LbUWsIVbVHFBXmpGNqqBeOjjHk7OsKKENdDmDUzL6Xe6qk9Vk6eVvSQGSkOLl8762nhqXbTMIT8m
FmxmPfAtp4EylT70pc8WIJMrIQw4LsOHfwN7le4+hZ3FfuE9ej+MwuvKxV2Q8L/gXOpiQy44JOm0
/gmtq9ue1IdTfBBhD1DDyec1V5KmgHmGkUXVq5I3Sw9T4P1vh+klIu1DWBowgNHcc212PXXrPHRH
2rV9/gvMK7LKvw60J5GwIQN8y2EXR7C43FNA0i7Kx5oW6vVd3bUI0qun9MOeeTqIe2e+2RjRxDQg
SZUVl9F2cOy4w/AIiDYOsJWPLURlbnk8J3F3BjAVue67lli/Fukx89wtT9nxnPaW4QuJicOeMWFH
lx8g9kVeakskWrV00O+cGsi4dFMYIzmWqCeqd8ZNj/XUxnO63u6ec+QNAMOe2FE9wKGyfDIgGWxT
kL8cjUjyyKlUzLK2L7BTcsvaD9744IlZCUMaw49mzIl6ID9PyBCICzufCpdNFDeDllybQrHYcR5g
XsbWx4Bd0dChOiYz8MYdhqDaBFkS1U7z8S2AMzmhXAjrwDr52U7Nddo9ChJlaA6c45ROqnE8djXS
7fPGyJDO+3SHOju8u24EuKIJQsZSPNBkLmzU6XelAgtO6BZUFjUnZHfXtPawmCr/3AwHquGyCzKP
i0kYv/q2jB3TNpzyYnRNvBrthMjtFLlKmoQU/t2qeZlPJnygk8IX95tdBBxvL7i7BC6HBY0/AAvo
xvkzUFjvPTAQokgWm/C4ZDwGFcnt8MjLsmY8c4eqjxixIV2eQAAXw+8tRM78xnMeQVE82iSeaySR
jyydoCPMWLiJe1qt4skvy8ypfgCtU2gqmBPxg1JnT0vaBTHzlIsvITcznWsba5vS251CiVUEWzoL
chUxjS3od2Kx5JIBoZ47DBDxBVWBAAIIzI/5TPwiTSNOmRzlePQmNUkVWwtiF7S59ffO9DBaZ0Ib
doz0HZDLOTL9n3uuJ/DYQNELJE0RrUGgUkFEQVPbLMLBcevLeNY8HfUOnqMd7kmjov3zxhGXWLyS
rcJPRSyBjKzXnRj+BGwkSr6MvpJs82FR2VX8bhJGPmD69f6QoJt7RqlIwUUGIW5LdQOXESf1jS7V
uvthWkeVxvSMFKvqZ3vTt3DaXEtmwhaOkgqgDPHfcJi7UwojL483WOXKtRz/Q4zl7tarSMp/9R5n
vS2D7yyPkWjMC2opcbO97e4VfZ3llnFKfmUjxsPEtJQw/GNFmBzd/diOrRCGoORE2BndWtIc9QmZ
3mJliD4BO/MXdyt6VX47JE+BHp8p3SMjTW95zskQd+p8l6PBsoP0H/hfUwAgybtn1I10sNY33AQN
q/I7XL7rSQcLhNteF5Ui3H20la0B23BtnxcIJ6HohnaX7RQZPjDJbG5sFJhZP04EFog1aAOdzh39
FbZQxxe5PIOVjpeyb6S9Fd7Bf5zicsnhZhYJLhUcyrLI2x4ZEyPdw3KX2DeNNIiBVL4/jFqL8TQQ
VRu56HVA7w9HWXZkiE8lk5Rl0/UDIg1T9JJ6k9N1oEzAca0v2/Ysm2V4W5mTUHQKaokRKy7vVmWp
8xK77yVE2wORRortAFvCs0s2jvcovgb3BnoTtHNBMUiwlgLL4VWIV6/yCc8uSaLTy4+iB4gaXh6K
pMioPYRlNrHrYdBwM66wG17UbVk8hJynTI3eEYkpMSJl0d9QsNbTHcrPqShRPjJoqEmHp1D64SfA
5TXrHOQDKdoh6pOiucjoF0lYzQYqaaqBdalgaNFzs45OqhmDydqkjQSVwnElmtKR1rTm/NWG9CY7
hTRbxdRHedMYNqfiRYLjwpyJnz56nbPQNOPKniT17P007/7x91Qcn44aQG/ZuM86fLeUB6OA0CUp
ZM7PgE5lRjlqHzc9B6+gioT3Dza6bEhiWtjlAXxrQVXEJYnS9mUYEdLJsx49gBjXaRa+jx52f0i8
4ZDTycsrc3EZU3YS5u1CWAqtYsWDnYGbxJw1nXJunp1zi0S0S1wg5MbmqWWMSSiWBaEsIglwLuGK
zi+GC/8I0HG5ekGH23JEXWvnwYRoPIJCI0RkTeUSxbwQR8gwBsFvAOEdEtrd8d3tjWi7CESBhdaz
XZy+Uffrf/34e7If/Xl/dlXldQsVX/b7ygjyP8Q1eR/Zl/379pmXkpvQuyebz8IuzA1x9RvWNvVN
amsUMOsfaR8wAFsuKCLYYR8IKJ4UnbKED4h2vXVIeDVQ2DDwMRf7nJCX6GHaWp7tLetXojARjOCr
L1yubgXqFxmsurbZGWuXEzeNAqiuNNq0rY9dU9mh1BZKIx+2pnhyuHhvTN1A+xR/n3Bv3LTP1UAS
AuhUHZ/G1Oe/4VJk93NtCyy+q8G/2TzTy30InjFz04Ld69NAzcVjvA1FoNIc5Dm67SFQDeDUWA62
dPbTnt/Oqt4v6dbIUVJQIjXdvqH10nvQPVSWozeadb/pliWiUxxFfNoy5mFAT3VCSWN+vy20RcsP
dlHnOIgRQzIEawB6jiCB00B3IyO2AXOd3SeeLOaTUMRKpm22mC8MDVOhgEe/plH2B9lsogjETkYD
P4dJjcZ1mWBlPp4DFsBpI5alZRFGX/Zr/JZrWPZiyg1K1iaOkF9sIYYdESUQrUdZVbm7LnOZAtAE
1oj5ZOjAX2yYpWefoMm7ntVS61yEURRB8UlOyabHdLonamU7j8hgiBpBiNrTGbs/CrZQ+eL2vFPs
qnZ+L2zm/+Z8y8ekw+RRDZ+7WJN3t4E+xVCaQTSkBTkT5zmL7K0FLnDnDO3AiOio6TJAlWFosfEM
Nt0mGwjIR31tA/XWDJ9Hejra16S07+QDdudUe5bxUnIrcNycsqpzt6gtn9KX9kB3Dq91fHYQ7xim
RFsYK66fS+lj1QLP7hAv7C1pO68i3G7O7/pBYHR2iELU38aumP5lh7xJVgT6PSAWX9dN9p98vYke
l4kuTg/G1epJyt5Xhekcu+IyzscUPCheYmSn5JoeVG8ZY6wGfvEVt7ZBX9uffTiu8CDZbrnLiWWZ
S+yot/t1Ia+oZYFw1D1ad+YynJrLH7DUFZpMNdizIhCWI+CjKXCX9gjVEcxBhPsJAlsDFYSqqtYZ
0QWlkDITVmwKQ9OTLJMLkvMnInP6c9gVd0EAy83aCObKCXqs3l2dxt/xi8UnDcELKZQ0ZCXOJOFS
+aLgrnZ3ns/SmNnZY39FaE0Sl7dwbySjl9aCdOtLfmK65qwGk66wCMvqc3C9lxGDsrUtTVC8HU8k
evbwZ0VN3Nwg/vvsJpQkmUyTco6QwSqAqWNuZpaaVsVXywfCXjkXH/z8DlbDYFQcRg+6zTu4cSTu
yg4gXbHzB1Dz181nWNKZaKr/PTJK+zwiYz1qXYI3xB79CbN7v+dj0476O0Lv0ZGE5kHoy1Xa0EYP
vsRt8L2WmcD6azcKDuAHc89BiT+rDyuGyf59xFAepGhKk3cMZQkzkDPSBMKIalBIm9bT4pHvtn5q
v9Zf7PoMG9m31/UfEIpbsaY9rRLm8WS1P3ajEFg3Fg2OoWOx4KQEFJY8tvOjVnC8RM4ayCE/2mrU
sIHZmwXjAXXD5w+VY3T4QtDifmDi9BRpP6YBwf/OvCARHZYRZhZbHwhhokqxFrPxDZIvw1gXWjGp
skGTQGMcYkPUoSIIlGjnwSzWlUHzPlJRfCuFys+fSmQfm/7iNmCBKlra4MLtfk/AOedsepipfOns
Y3D389d5zn2fAVWSmybkqrASRr6sdJgInI0kYJcASiYypySiLJ9LOaxYh1503QLtEy1vbdZzF1VE
4q9tBHR1svOf1fU4FzB/7LhFK69mLpuEB46SveC4zV43OaC6W9BIb57qxUYqoHzvRlwxsMHwDRzP
GmFHJhEL+1GDe4bsQ6nYfJr59m3vXfWjoV49v4EaVhBfYDFp9r+eFFXfiMuzXSXeWpZVnk99evf0
Mj1CxLrilEUjCQZJRCJI3+gO6xjwERFR0jjNtAoAynnd5XJ17zbr4fhBnwvX81g4TIlT3vHNvex4
GCtsyD9SPziiaVdYliGHThcfelr668wlteLKIislMvCOjSgtktwTSiffSP9j410Xn9JIHjmyUJqA
LE+oKdjyd8f9Xt4qeaZ2+LiXDG8ph/ceNc+9KGtOjeLJax3SVp5GldbRZ4LYe1yPDFium83l3GR6
RHBWk2U0e2MqY/asldKvSk01cv8sxqMcdzLGkiihU/DXeGDysYmZTfZiCO3t36emXsKzl2lDN302
dXPQz/wK7+hdXZ1PQqOd6WmBH7bTYJ05fOiCAfnnPNUE4UmK7N3XB3vpPd3MWYupdmBsea/UtfuV
iedg8JFf6l6aAq0H5GKrkF7i4ZUUnGVS0vsCeEv/D42566+toOMbb9dDWgXnapDgxHCS8dywN/gp
Sdd8Vhetj2OK+RBstkjkNzMgUK5SIJ+rvt3ATjRs2+xHnQscM1e4tev6gHL/pNia5EdtRA9gP7oo
VRGfNBqGFz3ow34hvJqUHOB9ivg2vpk/4jwNzJeDwaGfYl4QCLRTY/tpDyOMws/c6q78CGfp3W1Y
9zNqgoR3R8rPngf0FDJpyZDglUuBZiLTgw+OWaMDEl7OS5DbbOVuloHbPb4HBuQp+CCNmR01YIRm
jqONapYoRjxBL1H8iV0PKzXLoluWwsO/D8gTqoki/fH8TAE8rekWWeatSYwMlscKcoOJ63X88l3o
EsjB7mEoW6eZqWNHvOPyDr5uGs3DwByzkhrkwiU73jAM3xbLsPNtkYXl21zaHfRyzNvGhc4GF3BM
BhiZlNqOyYZ8noIWhK1AHALSzDpBrr5osZHPvwaaPR3yobIFa3/yBABWLGyUr+ZGiPC8h7U16c4T
KJS9Bs95Jv57LtLNo9k7FusNCZc0eGpfVUKjsn/GG64yuKFNxMgRFdh7Hpq8MfVT8b3l0ShH96/R
3LsTj1HumvIKKAmS+8nzEFBsfrPbk3q4n3H+jWKR7737LcfyZMzV0vLFCKFGHEjBUo62iu0MwFnq
CbMNyqgvamiTuMZQyF73+nImvEELtanuz7BNaB6iXoZefGUoQrg0jp7YwqGcX1PiqMViiP/5E6bQ
W7uNWsQvWdlPxOfE2gOqpb0nVb7RRvgZ1BZjbzpHinqoTJou31g6x38cH8X53uDIcR9yR2uq3oHX
ZVxLC16R3VWCzwOk2QXZE114zsq9WujmMmPbgHx7N617DWFovf/AKDIqD42pPkBviEWBUrPnh1ww
jb5kMlFhHYCNKNLEoGtM39X4JmfEwkZU1GW7nkvlfVH9GaEhsPa52WNN2sv47Nr+0msUjtPakSiD
fIkUe23h8r4iPGumJdFB9kBQlCjWk6+Vlj4EqEpS3ScWERYRrv+89OjCkbx4DxP3TEuZoWoatLmO
EdXUCK5rPy1fp5eGdC0AI7HUAXvG1LQIWqU93P+8+W3kvM/W/TC6RtiEULVsdCnUTt1cscZZyLE2
XXzL3Nobp3lAoLC8wYYyZfwVOr/fgsfHy6F6Q5Cyu7d7/GIk+sGPmbEiLWKCNrRnTAdnub5yzT7r
E7oVd/MKNBMvxrzfpOIU/qqPns7XLnLC/VEzrcnrpOz/wymtWWI9QYTb07n8CzKBANJtJ0Vuw35d
kAXCWw1X2aYOYvlZ6QSHYrf+Moa2JM2gg+potWabgxdaeFVddXffg+eMNaTX4PMwBpowWzkhe0c/
vql3v/8XCF4rhFGhB4LFeX78pc2j2FN+QdlF2l9El9RLCbEIE0YCFwsjJ2c+m6R/NNikmiZ/waoB
d9Nb38thGQdDUHzAkRVVXsOPQqPGJVy8CpQ5WK3Akc9SilURYouMzBBkNaw2VhjNZZrhpF41b3Yo
T49cx41cy8dVgm7pLAxaa9PzPYvO1bMIAtZSHd2YeLfTnYDeoB1vGBz4Me8k9OJUGPNpRC4WifQp
PdIKWUt9aO4wf8Pzi0JNMV0Kh4xuC2BycA2XPOEaS7sU4EN2Eq/KeYHjeid6CpuKHyLGqika8qw3
W/5bknjC5c/QZ7/zWVjAoel/MQFf+sAwIUXcTTKPsUm5TsFwn1qtObSAzXkf+2rbmt/nRlDIgWJC
asq2n1EppSA1hVTVwCnIW2Soro4gVLS9wMf/01zMlX+80FmBJPigUO80zVtkxsznKF+U1PMNTU62
8eKvBNf++iLzagpw6E7hoYX0Q1DPfC+//6re0EPp9pUh6patVTn2yZVGo2ahbkYMTwgmVcV0sxtK
BFl79FM5rSYLcXeHELz22C/NOKwQ5zgqljOfk06hhcYXycps7THBhkjexG4oiWv2xH92Z7hHKKez
YKir1x9BBfZ19NTOIm2BzxJclZy7Dmo1m37sge3NDixYzO3UBiOWlN1r0LP9BnipAmBxkLpC+01Z
XLldrpouKNxA4yAbqBtntNSNgSmBh+FWRAoo91sbQHrjtPSCnhzpOX+EcrXoOHoX53Tr0KdlWH4N
e2JKzQuGCui09WUgLEmHkiOx319rc/iXL893E3GkwNDwDZVJFhWTz3ghBQoMjpkS1D+PWU1kKm7C
chOS86/b5NChYIEkKGEmtXumrv05R6wU+QPF4quCKgqHIvbtvDEDpSoflwQSTvSnW0kCd1J9xhtC
0LtkVTQoUZ73MeeNQhlYLSE64pVDyOUKyMfEx1YirjcXCMe4CfjJLou4qiIL8VrF67KwbsNtYBzx
SSisUpur3OtCcdjsdfTuaRi8Otc9BHrsNwz4wXhz0NmDfEyHleautPFIexNTGiuOJ8V1TGM+Oduj
py8htTChfhmJX81nVI2YrhoxXgVer47BK3He6lTSxM76h6pO5/ac35Xabg0ZE6TVirBokFyI3OSL
bz3JyFpy9T+7JlEVnJS3qx1rQlOH8Fk5rFWcDVU6ZmyNXKKtR9w2yJ8eLn+YgoyVodN1pPenEkTR
Qz47nR+S8AwaoQ3oW08hO19ihmq9wEiILI727AzXrdiQ0GIGoIRNtuUoQWgb8NS3xWBRq/j37XCm
jXDLyHJwQDSEEK88571CsPR4mW27mDckqO480RF3qUosQGeYaL9VPjurLAbIORKVxpBKBumGSeqZ
0vGSUwI2mOqs0AIU4jL+sZQSxB5PPwv2IUTtK51ppTypM0+lKJwLI2J2ERwv94HURJHftGFocY+s
SYKad+UUiqS1Cx9rz5XGkrst5kQL5shpHSTcxq5Pvnau++QwXKW2ueaiBaJq99Uby95b0Sq7iSzq
84TwXxfiVFwuxYYZ+bBaqSWVhUzDbl9r6lYN0rqCaH3eaJYoUgL95Vu85272QrgStsAnBpfuIAsh
KcZy8qFtFbpXKZXusQ1uR6zPXQoJj3m2GIM294POp/Vi9LWHreWO6wVJO8CJczP4drtHhlgxP+ab
J2Ec/f0h2XbmkzvLDtP1jtYv47Fo54+CV1+LMkVPzNLhxje3RmudRi7AqXjW66uXNoDKL6Wn3tPm
g6K5+rBfb2Zxw5hZ95S7eyUEaESJBIsDCAUZ/rH+Ik8zJkwXIJn+YO6KyQ5tKjucKXvJzQdZOVSw
O8X5YQaImrnBCUTEyfdYMWHsHfqKCAV+6ltbaJjK/WHaHa65ek5vtAgrWEquYU3tmmmZsy1kAKtb
uOJptWdaQJMB+LDgvVyX79vpkyTz01XwW0kU0eZaZY/t9DtVZ79ptobbWBy/Hr7F1g3IPFxim2yf
r8n53Ul1TOz+QSGkUPanaqJvy/UYOadttye6/0sTmxf5Lm5dqqh8+V/WQfEL3Fq/Bt+T76PlcYef
1OB0KTXd4do9Cki1uzlEA/k3VBFMC3n4Orje1tj4kJAtcQtDqPtaIrcKlGilYxgI3qKBUZUVQajQ
ICaVhHLcdTMu2JIFZlwB0zzTMi7N/iJZnn/KjyXHi/6GRhIp0J2HTB1gAd9fDH+c/im8l9vD1rSy
AvivX1eBVxd2pRPcE1eIha3JBjqEVorRfEiKlLOwQWm6ISPflK0lsEDebYWAliysZbbg32VrvWV/
ywUl1T7mM9fOtPyJk2Stu4uUhxxctJb8oCotwZGgWjBkG+NHnFcIZWLRhn/dI4R+6BdHkKHGqgiH
ohrVhMn+j9NAEV9Q17Of7LSLX6ZGymtAryhyYs4jvNyEjixRx1zCxAqayn284YEC42vpNjOJXwYA
MkWx1BiAFaTo5dD5hsAwnz8oJ+ze7gfmYN2FlFrMeD5+QQInkpUoS88bU20CA6AvbO7k18vPFD1o
OtD07I8V/RMKeb875ZzCpw0hfmoSbmKai6u20SLf2l8sqKo7jpSNzuCz61ShrgF5miGNcGDlABHn
US0sc/y3yglC3HbvpmHXbUImA8042aZ5Aa7f8GsEsLpuvnbv8FGgK//AqX4vXIV7XER1G7YtBVa7
E2QWJzZbFK9a5d0OE3yPQrrr/kXdxcqZh+h3Bz/ME96S0RhbRJy0Iz1rtdqatRh0u8PDa4O2lC8K
6xAcUWecAE6xiCF7d6vN9/HFSZTF5a8dGePkGZN4n1dCPspP3udPKxg9IzW2+fxmVWXY7m79CDcd
DWWRDc0Mv4NtchYA/8VEfHqK850BWp6OTyslO9RIvhiqcu5E6ii4wlBjuf9K09BEZ6GmkrDSJllm
w0CplkBl5PiIKVrUByiT+44SkWTWUx1T3UE3G0n7lXx9OK3WFmP8ufDvF0vNi6nDKhGB56DrRwxB
4thOHbTNmwY8nJVHxwjwkw04f+zfsn/9WP6ww/I54LG/FgdkKxb4y1SRRqgGsHRPsWnryo8TXNPL
5gsLPvcYMi1SSSV6NUmaILPKZzuoShMXVKYj1B0cG+fp089tL7wr+Wc3qDcsjO8iWEVnVx0ryjAS
DSqBq6XKVdGqlnM4VxZCtJ9pxoXCOdK5kA0XYUzinLA7YjEJSmsXqooeWbiT05RDMVkkKvq/cMGH
D1OZJgxJwGkX7ll1adCD7hBbMkMUYul3G0+1Zt8ke/NPwScuwO5uf+WqxEgiciwPmGCcdsbpw3Gn
0wZ5IW+dkrfi7oQUa4z74KGtYr5mYT9lsG4Ca1ylwiQXV6lY9AGR8FY6suwBiY+Bh9Z3WZFRK3zy
8WWWoTPbmJWXyLct/MOIn4ZomFR3N4/7xJZUhlS1EJkFAOtXgS31aFeWO8uBl0tjOCL6hjh1IEz2
UrQmXeweqloZmlMhSktH08snr9hMTYteDWyeEYtpVn3BxBbropFXdcy88DIzCzuCZ0VULOARSrJx
GDxDQ6+sUOwYGTwc233Q1Aq6Y+bzrDtG6YWdgxwi3eKx4Hd8AFwtAdtMLRihIrjqJ/dZj2V4nz7/
5HuwB0aMIkExlp5E68TdhqeFMSvCenx9xr0pSla9bbDD1RE3Gm2w+hTma279wJWJWTzyBLvbU/UY
57pobU8UdHFxvOA9K+3ZO1nJnEXYLZdieDCYtVRYTbs/4OoyFpJPF02S5hVts5iNZjJfqDwgVLDq
JqBckd4SBJ+aGfOPed1p5EGKXArH+OslR5z2za1HgoxtFX3CXWcBrMCiLfFkZlIL57VpvxSarFQ0
Rb/K2BtDS/7waAM45lOaoZa3wrsV1FQjPFt69H4fqPgll2sKA7qBoEhFK8VifdTNWj83s0uKXChz
mW0+nizSdIuucJEjs6vcfOWdGzxlFT7RhfklyZDIbpJEiCOMvTbhcuOn/F4oKzmbGQrxFDaAE5fi
vhjq2tzXa2I6V3tpngs6WSUYgBTJinMxjwbL4hRCXKPXHm1G4JWgr9F/lLtAmGRnJBgLbTRDtkTj
ww/oKTwUXANbqzpsAJGSym2+8YQtYbwB1x7k5Y+q/IlXPgbU7z8tIT1P2atdkopDhqSaVgIGdkf6
vWBFxQlNonPkLWzVNtNlqubdvQKxGnzqXu3nm+DwTZCEL6C1HWUUOXlnuxagQktROCjIKrjf2GdW
bg3pke3RXFEsTgy5hOiH8J7Ac6fYArKC4oJN94+FJW04MpD1k9pmsCo5p7dM8ksdL87jYBCyBtq/
MpxjsxmxiM2D9fBXgzTnvwxHQ+cWr8Fon8QMIe6G05GtfgwEJdJR3yrp3dXCH1VMMxIdXVAp8JRx
d9Rr+G3aAqBC7qb0p/je5kCkoiFlcOQQhZMj/KU1l1IPS5ArCpJRNYF3uPRfQp8/QUUTktpCF0RG
KAy72N8Vfzt2eWmrrwRjVdiEwDFmSYJYOgH2TZRO2o/f+zvlaclECj5rF6NO3+ukvcivRHOah/DK
v4QYPMi+QcZcCm+4ushBBNu+sPFeH1ENUkDocbgsEzWfUQX7j/ok1O0epqSvuH1m6N+B3bYcooJA
P8cPVju6Q1QAvyX3bUW++9lC1X/ljTOKusxh+oBM6d33NEovQv0+JgvLqGVTuIJJxRIqnfUDLHb4
tIJdY4z9rLQiwYXCyNum3RSllpvm0JnmS18WtBZufFqc58/3IJ1XZNPxwNA3nHXuF6psMAFwn2lw
Kvsk019bX2WpDww5PvhQBx58hjjD9hJ7iaTVvcyQ7JKxDyi6xdrl6QCUwTDFrtL4ML5PzBcjIe50
9h3lssz36chWJueeTaVgRzco8XBP3pqHlZxtJIqzErswluBeEXlbLHHEsFCYx2eQQ//qSV3pFjhM
sqt7HvYljP2cKsyWgcIBwZJW8AIw31SjTn7gnSnTnelWIHqvOoYlQB0zRPVqewJX45PqVnKyLar+
bKE1p3gKXhMgq74Vxb6eqxHKR5Iasbye7loUMzaX5vyT/T7USRgscBDM9gReOx6keTFgdamRN9fS
mw2zUk44BqKzcyJZSEJovxKmh0yxseRO63M92oqWHFwajXgatzGpdCo9NE3SsjcGkcUGGl8WIzan
c65V7AiOsCgt1Vepj7IyZjcm9MPnw6vv5yXh5nKXJodtjwYMhNPae0EbH2Vvi6vnOPI/JiaTaQzn
Kzz1UoBLUWkHcOd8k+p51W2uBVVblyP0bllmgeFuB/V3H5l0r4WNsN95okI+r3lda+fRod71Tg9G
rKd70R7fboUwPZK7pJqg951AaIcWLaT0JxoqOcXLgNjjpYxb56fpnPFHd2E58NfzcDojw+yzZ3Nc
83SjK9SDeNLrRRk95tVYxCfYFEPvrp5avJPihYG7JItcZ2zDF+9+9KX/lfClgPY+mQYv4YMewAzI
5givvR0/PXlNvBiOSTNB+X65xKZnZEiCCS0/QhUu859lbR/e9QbnQVr9Bf8SPup4IMy87MJP0LrU
tEhcRHJgHgbSWmD+TYjhymh+LwKsN+Vphezf0WT7NWu57j7VR6YSCMOT7BlHSeS9HYnjQMhgbSw0
ZN5+8P4GmsdRKh3vkaZezmk9Ly//6tcPwd0I7g9n61dNDSwqFDSDFGhdh4UO0Modi0Ojgt1i2T2s
wD6L5DRLF+PeaMuuGX+vDmySHWykOixmKjWOBkkCsJXaa+SxdwuExl8joZpRa2pNoUZh4cqh3Kgn
GPqytWAF10jrUhhfUXDw/U62/Rl02YNNtM2H7tYJD6F8+n3KuqHfmyijFcmOLo4AhDbQNpYSK3nl
tkBlGlcwY2xWY9sXo7/FCWPB5drmaSczJ4PKMbIg4GaxQh5t6u5Dn/YkQq6WXB5SFiD/NOgl5Luk
0YAR5c5fJkfaJZHGE32K+DOBZj0BAupGtq/JVt7gou4y6j5iY0l0RWU3VNjlQ7kygMFbgRa69+6F
IUXxIb1vxlbu2TfU87JNsKcucMpcoCkJLNKQXKENlA1bQW9cXxZ4YgbJ72BzVGw3o3QrWS6m1ikA
Ao+tp13L1wFYKKsbWn32ABhwv4jfDlObP3THvbCp8O6rVtf7lNFfyaVsedcsPKzlwetVNtVZLn73
fatg8FMLa3KvhHuadKXqczjNLI6PT1705oRog5FPTsi9rsPB6pYQ7/1xXBOKJIusT3Btm8ZcxB/s
cVuG2iAn1rnLjvOWd3Fr2dXGba454tqB8q8tjVWK8vIISwZr25VcWPpq3iALLQrxyUpw6YcyrsOp
QhoqCz/qYdIZ9L3FB4HHUbldAIxFM25Bdc6OuDkg5+aQq7Y2AwiPYgn/+L9oVVeDsBScalEoKSnW
lN3fsfboF9VZ8e4BlZ0B4o1ux8kFTTGMwLng/Q56qeqxKyZiRoOZf1L+HObf0Il4rDg8jl0TQZGs
aHyxNHhMzx7faIwsXkUENayHvgJb/EkvQ4GSsK7tkwitUHe4GQzWHSXeIARa5rsWZAKbVs2B+myC
gRJ2FU2FLS9ysXVJypwUnXNni0pxTi4xjOKuXDd7UWMgc219TMMK0CkHAqP4c9MhTTHkYbWi3jP3
fe3Ssm802Cty3pitGf3zXlpwENdgAZTs7A59HvKs9hkCVqrANFhDUCbPGs0WPDEBhEPOAStnylIt
reMur/3yIMNWTnAZA6dNn+3vM7l4uTJxM8DB2e7kHwKIGBTBrTFuAY3crR5UAQKQiXA7XniasaQY
pFeLv3yNurGFSBqfpcnPpnmvyZGOdh7oDnnZX1APZsj4A35uJoUtb9w/aiv8x7HPFcRuZCENehWE
PDfh14TkuAabAHk3511lMVctq06cnmT5BEzomJJW3kCwIdlFh8WLgg9tMtLP12jm5UlXfygLcJLL
SFIArNDftrbYLKOTkAZtcOOxp4IPx+UHJ+gU+pIvdwAgkKLrEvH2j2J06A9f/qs/1QMSXwZh2k9y
MSt6Lv9ktgXsz7LXMZcmyNKjeXAzQacjlfHtgQUI/mDIfZhbZPm0cSxL4fSIkYR4J9EYtaTzXjen
fFji5g/bGRtDwyLz0XC66ePgjtNLLvLWPL4Og+/HLyqLLZfA1i3YpDvJ4ywxrneBouRC3SUqi1Im
j85SVBuTAU8yHilHxL97HPxCLv/V5Leo5m1YGnXjRdvs4vKQ7i+TxlH+Blr5rZKHg5NbNnMTA77Z
zGJNf6zycaQ+JcOJ4CNmH5i9/FKcmNuY8n5r0P51vXB30wENQ9ukCRR8XyLBftCxJD8iqoTBQQaQ
YZH2tt6P9eJta9d44u1oKQ+0800KXGWi6tq8F02vngAQvdSilAVq520Ce9qlJtyor7gT6mx1v3NF
hdQvHymPpy3fXyoyk/xCWpD886sBHCVjxIFLn3VWqh5lxX3PGsSLF1OL0ROviZY96bdl3eeR7biS
Yz4OBo8bNsR7/HnlhCHahOKer31DH08tpwJ55/mTLWuIxXg4a2Ykf/32JrWUFL2NKOgGIMMBXtNQ
Fu0KAKqraCZDLK1fr5MAJQ6kZwF8r9QhAH4UPz9vCNQ4AXEhLl9qQP+Cm+nwQVKZ4V5Ibx7Q9ALc
zDuvraqHF1RJgChMOYkuJQvtqq+Cx22VG1WfokunbLoy4Do7w6ieLjzBrteupMb9dV4B4N42IAM+
HVkjlTWKp7dOl4nUEEZNSLzDj/SaouRFlubbTfhWT5Vz1Y7Bbg1p1LwmQIR8XPo0QHXq7r81vGah
g40NQWXSkwvskVe8yFf+1d5KkqZqhYnZu6i27VMgoi3WvE2Gh+DYbg3shJAfj0VPXzsIV5GhFH0S
YlA1FBHdgm0Ub4NDKyJx0b3nPzp0j1XzNlE8oZmv1SbVXWgNbawM6b22VmURGDyS56DmfG50MhIX
gZgGg8+A/3h+0UDpHuxoHkJZdt8jXXbp+AZD0HO1uuaUDXGxoZv7vpGvdO+EckgtlHtTpylLr+7h
9U+2lWGyEw/5kAHK/9UJaFroYHiMzKpyUBWiVA2ZjWwh+B/f8khk+JcWinJ8KAI0nJzAuktFb5ts
YJBF3GhQllrmHP2JYe74029haYf5UTAQdQJ3FX+iSmnoaRZQNxEbmTfO5fcTp0mjm8ZHbVZxKe93
i3ZzNUl2qMujMufv4/FMIsz4KyYRIq6lfgmXdp/Xe1DFVkkG2wEMzhEySojI8w2g6659OSnsSYti
a6uiAjN6lzne+/1kS33BHKvTU1YzZ4uWp+VcPpMk0nKO/GXqc1jC+KA2KIe4XDKJo0IXSVzCUhrF
LjPBLuiGJkxTHkxeRU3WrmOVgfYQ3pPdxq4rcQw/3snDQNySh9FYNiA3yTDJU8DZJAqCx69QY5kk
3BWCeJJ3BNF+wmZI8AqLzCb14ClsmKvLQOTn7UD7j1X6Uxj/LHfpPJQm1BKFF8RDJrz7kbEeFeMF
yI7Nt4eRr0DBNOguOLPonqZXMaEvQUwt5HE1U4qJeOFkSvPLoTwaIFgmGFtLadh1APbdI8QNiw8A
JoakFpXxWoyZqt4YqVcgRhY/xd1PTiN1oZKfTP+QoJrsHUF9rqTXD1VrsXRXwS25RVegp4MdPdSu
rl/3opYttNhgtgV3+pTRGPEoLvpG8aAU/OtXnGTn7+zdHCjeqnz6X9WRTXV+0eSasKgWsCBQsa7c
Jf/JbPQnYU3aTlT0gsxdpsuQxOH158CpglbNKNVNT4Pl3R0kR/omdopVlmy7g6Uxc2oJXcWnl+gN
E2UBKLnuZzJ3dveaG4DakZOIfv1xjeuCocki9YeNGW/osyOMURFJBjMX9W7RVwgEC+LET4SSLCIo
r/umT8yIoH5NgVCyKlWt1i2ea3XzmgImOix0SGYL3bwQR9vtLaGPR7kqrx4KMfXOooux/ivUc0hO
joHys4NlTBJc/YCzOFRUYaBcxwqkhS4b/l/I8pC0j7FqUu6+XJQIwC2/TZBesCQmeA3oqrWWzSgj
OKR/S8huQ7TGIQ27EuzUDWnlThHJj+1chRIU2cxOgs9KhKwT+gWsuoIeDCsRq/9rwlOpEUa93E3Y
OtwQiPCpJHoDPJtqN77QbQQZtWKHFir2s76rEBirhpXWaC5Sr8qBM8+pjgxduY3I0Kz+OUqG0811
hQKQX7TeHfcat4lnN/Rx84cK6nPiLxTHKZTtuY6WWgmfvYsVn3UKVr/smoE5MRHUbE4e5xQGD/D8
5dwfZqG6KrsKeHpCsu24UiRytD5PDyJH3d+VkbnqOx7tu9DZHpgSvzPFon3dgmIJe/Vvr50OdCVe
fNP1XUpFNzdnt0aMkzekffPS6IkIqA1xQ8pNi+xOzvx7mWNkQBy1fiM00RNRstWokEAlq/5YD1E5
Lrr+10dqZN3AbI9+01R18FopuyS94LhxN6GBXQ+6aPNI2uL5yAyqSswz8m6tCe7tRxXFwFN4e6Kg
beDbwwjBJD78nzK/RJ3lzfHnlTXQH0DIkCKu1CnNUGQMus7arVg4uUAftaRDRfwt1lATh6LpQvcJ
QMZ/VuCbogeSS3kX7val/f6vgmf+ogPdAe/kQLwqCjAv7lApJH2ZYdnmzwk3nJqaR+uDMeXjTuoO
RgvBzPCrbcmDxNUaQ6GrDREh4xVP9moEBe5GUCYf65c9spQsGv7r8w78zscuyi0mdKHjVCgw4zej
CgilIX3nuto12iRhESJshkf3bR4AXxLrtVPDlee2R3b/ICxRUTHtPUWPadgSNEeKh5vzgO99PI2l
1L8eAi7ycQHBW5YP8p+hor2NC+RLWf5pWRmsB2Wyw+tCucxbT1q8xxXAZQ4IsvDYiuLbfJcZlnp/
Uyde8N0G3mfAlCZ9dEc6MO5vZyIkS+LalQ1a+kiXxPXtqPtESE8WYHfLltJtbVGgKQQhg24BOoCL
I0xTw50JxgqAM5u5EDTnOOEgLujIg+GcBbRZRkYzu1D6uDz6bEL+o+UoOZEgCTMd8m6c6APLd4gG
jtALC8oUgtLKPCPhJJRxPyTeUSCh2FSfJDAM92PkEqGjJXS4AhKw9hrBnyM79VaCPrPofdEANmDu
c3tZO5EjU7wLA/Pdv7/4j0iCg9Aaht9OhluI4+LVo17CSgQFqwurNKO2THmnZzuEu11iRpeg1jsi
n8p3fIMUEnrIeTaB5mAjFbo8olW/piNfbsAs+CgP8WG7u9fBtZbWxdNtnTZES8/wSphouZlFqKGR
EoE2B1wuOHAdIh2l9hII/t/NZSL1fT9m/9/pGC940VN5FiH1uq7pD7ne3ELkmjGhbn1MzGWdVSsd
6YN4B5tf2DmvfqPUKl43fzodSDZxLbv4UGcgX4lmEbOd/OxPgGyXW6+lRTw2EHLTxhPTtyk6SvXH
ETBkjbIBlglW2Xze++XEM3IxHJ8xQX5G46ZHceZagq874ffeyj/J4x0MTvD9QwAliJLgg4Iqsx5h
yEaxdlOUveuz+ZSCntQDjAw7/dsarge/YWH/xfc+p/xztJrG1t9U/peS7/W+fAe3/YBvtiNA3xjp
MFFLcCo/wZ4GSz/6GUR3n/R7oC+rY4dkyO9TnVKEOmvPn0UMTLUx1/ZxCIhWO3qfaIh5s2RdCdx4
Km/soS5nrsZIef0fO6Ts0qV/a7S7xkCGuNNwFNjoyr7Aj7Vre/1sfJo3nWE3yPIKN+txIxbmPk2z
P/6hlAh9kD0mAWqU3UYmECNrXviEdW3n7LG5KpyUTHfJxOPEABC5DZva7q/sGlZxsSBl5T2Nt6z4
ssx804KNaKgeQyAkbJig0b1bMDs3h6Bh4DOggn55mv2AV+Ne04BwByA9/gnWl/uTih7faI66alsM
9nBaLZfczzOhHNPE4WZuDg6+bNH0A1zyEqhN9JY3Ij82QDPn7p9BnWNGa9Hqe2Czn9ldUsHgsFY+
WSsvkzGMqqPdDZFgFkeGaKWNzJwDysmsJ3wooemXjeNQIjgBPDXPm7dovNilU7uCgUpH1s2W+d0j
YcAZQL3YN6gkSHmtxHo1T1fg27jb1WC512lIvTbnt53+3ubTM1RR8Jb8vxFWU2ZMM1I9H9Obl5SL
5IqOVcHeWib3TqBc9KYxNZHRCG3Bdl/xWHpr2RDAXQPCPx+UyfGFf3A6ytF/+sbkh8imyaGw1A0H
4A2PgKdqR4hJp57Ge+jqlefxJRshCbBttpWE1ZoYo+Y6SB/4X2Y1jn138ACEqk5tHbM0SDVUxDbb
9OXvd8QKZaA5fR+u/H9xp1WndFDaJgmEUb21OcZ7qUnX+QhVkZkf+Q0sadexy7u+1TBHnr2KnP07
sTjHFcxUccGasmJ6AbChzBwIuyfxa5NGFmZHZFIAJTQbdb252+N4U7LY+wFmmWj2JGLPbYcTjofO
JFSHOL7WiZd+vefbVDQHGNPZK1lvdNFMDcElmhEtvBKbsPwK/d1TdtS6DZSZEtvB0cZL0X5V+buM
rVCHDDPr7dYJelpUqctCfNUmyAXw5R1ER2ipFsQBPc9EKQ9WOlhdoRePCA28RqH/jcWTG/cF8bIQ
HfPiQerNEOdU0wwSZlWCDa1j+tnS7OlV8tB2UWzionuMHtghUsdw7VosmHx+L55GlpALJIfIw7Vu
O52iO39FTcjllM4e+Wqdxr6mYAxSDL3sX1Zqln1X07DnHReYxbIATVZDLiwuBKTSKNKbr2dViQhD
CUughEEKNHd6xbUDOzNxWk5ZmkD8+liiyen+/OuKhp7FKMAEz4l7urkKC+Epll1NVxHrRcRjykRm
H7ZyjExfG9PjhOXymDyW53bAaOB+80P6ErRrn0DJKKJS1m5Oi/7fmKf7xE/EUcn1zKFQTTIe7odo
7tpFv2p5vRy34WoeCDdGOvyxZiXfrTehaFGTX+nt4DYsh1nevMzS/V3Uttb3Xiln0ylQIOBaZyd5
c2wDNWRMYbkIxOAXvS4VsYZNgOV87R6+H7YmjA7CtiwnyG+rg16TTOCMhQO3TIknORZBNdFuN4Ko
1Rfbz0TNm7bzKGH/hD/kvTCvuUDYZ8W8q209aMgFmVQcdPM7+b1fmRCiz3nPEK9ji1BopMs2TwNt
BLpZOG5LH9Ta3W5uFLKYHScIzlgqoxiGBeZVvyOHxuUPvrVYWup5JokyEaPOTfYsDAc1+ujycJZ2
EE3Jvhz1fERHMz0ZPFgJRuwHjBk8LWwhAeIwPQhXxnUb9DWj90h5y6SEZMiaySbSJQxO19REia3W
iphjOAyNNvsTqA/uqVSZe10apyWTn0mLD9wv0H89NxJ5W7CXFuSD51GGTbjpzfT1Oz3y6QNS1s6L
E0BsVP/5hoBhiHoGyFMmmDPlZ/kOEnIied2cXmIMI+7JkZhvrHIrUw7AlWwaB3kZqurb80Gu3vQ5
pgapRom1yD8rewqT9TeZ0/unqOmy9xXn+pPxq7NwzcWWC6wBfDSPnj+6zgamVnUmv7/ezYd7/KSI
Ul11HHs/ZqMaUnYo7/fQvdgt20eA2gDRs6rVRAeDbyMJZ0i9s/LFngjFkZIPFWh6Bil8UBLc06dB
ssPm1FWQ65Btx3lY5MfwKKmb/7yvH6EhJLWBqD+ueQA+uj7XHbYtt0og1WbHutiX6B6lGeB50Iig
/sLCWp+scldnvAznqB4mfDP3IuyyCTkekoKeo+R4kx2yNGsVf3GNcAf/q5aObzETl8m78VyJINYU
CiSellnb1RmXe0caUwj0zxFP5ymrwe4KU35Sbw+po+AaR8JL9zoVXoKtRJcycTT5VJ1G3BipVdwb
MQ/uTJKv3/PLh1w2JmXNmrduhQz/UNLU4pccEmsGivDYtdj/VynrDRXyZFop3iV/6qHiHQ3Zrm8V
+OlBO1RAXrjiUxjzMZ+6sUH0N5R3qyJ/+tKmEatuBDMd1P5C9rNk36m/8NQZS+ilIh6pL+pEECKe
UDV7urfM2Gh0cRm9GovZDczr5MJjbrZGyxWbeoI45ERMFW5QbK3HL4FGYGFbUnRghaDYopvyqBH8
sCGthfVRQ1A70EKEpiG3hd4Z7XQ+k5BNjASQOek1re9jTZ5LVPY+SXHbqJ9fb5nQS8Gtpd7RWvH4
3hEcCUQnG4siVrel8ZTYxPvgzOwBzSg9RJTkp29XjJo270QdlJuPGDgOpuDgCb7yGRWPygflW2/U
Qrr8k+LrWxCOcUszTQTS+c3twzMTbt6gE0puNL/s+if3q17aYAyCF8HDq4/jpvWwoUilBknMzdh8
pDxYHUbsSbQjqtHWSUfjBv6Y0vsqlsxGMz+s/cm4/NwOyeqWURHqICFlczNaZ3yR77Sjo/5/a9FD
2YVNUzmH+lnZikXIkBxQ5Lh2+6m5vKsgRUbHXcLCLfxwQ2Tf4GGgECtZ+aPNu/n9T9rzn1wATdrp
iMoBFxSeGj47nMklPqk2/ktJKRG1rTch9R4vf/9+bf6M1EVbM+aWHv7OTXXRWnKpoccGyFx6yn/p
hVzWC9RgMAAJTSjV1u9AnpqLW3/dCGxCmyg8jPlbbpL+2VoGcK7N2YrGtO6vyOhFSatAKaWdcqKT
JvL7c1JLqpOukvbz+I8SlrH/lDMMwbJgX2wen7fFBdu321cxWcx9QxpgER3h6FqowqwdmcovT6BA
aOzqiB2ZpbGFiXRaJwfNye0GOUISXWjLG+I4Vq8/LsI0enGjN7tiom1KVbhL2Zx2VcdmYiEL/x6e
3t54CGHV3EM5IFWr7RDTAdUyg5XRLHg6Pb9n60RBbmH1cvOuNN9xy7AYuXa8RgJsoX82TBmAzJxl
ShqCG6v2EXIoB4ylqtx28umtAudygiragRjB7flqf/KUvP6UAE6TxuNVTbDou7iyXKt+r9Bym7uG
DUcMM8hNj1mNlg7M0BN9Q5Zo9E+Ij09j+AoPuRSZpL7nEq7R14J2Zp5jxM2RibpX19kklzS0yQz9
c/0E1/tnwgDnwVj/wK24FY7IGKobXYT+STx1Q05TijcaDp2JhYmxmPf9XLX39pcSKZunkQlh7lMB
bB+1qJh6qR7ySA4xu77TTybWF9NSAuyPXuDThg9CHpfTa2FRjmJ7W2QuBAJu0CTo43CP7IVZeonE
8qtMQ0g3pSLmsPDWbmUTAAVWOIDxAfiQqj6nV17Ebmbo2yyDGGRacskIcDq8sgXh3jtAIyoyyp+R
/mHYCHh3vnHDIh7q9Pqf9SnAzxioBrlAin9bovxOnjtmYrbhFWRZAieQ1YBd/frFQ/ioj25ZNlx9
iV1HSZbtv4fhHCCsjQUPk4QYppNN8zHraKwW8BbFFk3R4z18ctRZYQy5w5m+e2hVo0RaluC3kG9e
AyCpyRcgDA3IVVO+pmt6i/fMv9K6g/MHl2ZVzT7bMnq1PeL7Jd2NMA0eEAiPSRyr1KTzXSJRG7oA
hzyXmnPW2QJfJQHIBsb575NYrBs+7QcHXVfoDlK2YuQGeEidnL0Vf5T9dqLeh8AXjcB2J61lJ1vC
TdUQ/srTdaw7dqycn2YUkHdPhStD9ILFubv23+fwL070qTg3CXpv3P7bnkRZPyaQvyDsC55udGHY
Tfs9lRKJwlupMV8axvbhJjtHCSkzuKzXJ6ImlQhy1sW30e/KwsWaIeak2WoUtQp6UI+CwYObsJPi
QKXNeiQAHy9Q+ShyhAgktBAZMf/TZrBLOlmwG8MTySavjQBiIdLHSOCnb6c03jX2aqDRAyvbSskM
NJm0yTXt6o6u8zA3mH2KoF/nl0o2K8N5JGqqvjzOXWEj5hR2MnUfLHHFxOZrA2CB+mFPYtO5cfk6
DZDBOr2CRdtLNSzGE3VapaJKuNvqxZGTqFRo91w7KB0UGgVjzUmNC678aYj1dVbDYjB522Qfv4BL
xJ6F2zwqvNFkSY92py1Dy0GiYzTk+unfWL5MUFwZB1It8QHaOsD3T6ontdaJCCE5bqRrG1UIO4fd
0xJ9q2Qxd5NFpfB8MHfKK9ftC3KyKFeZSmfG5h+3ZkYUqwo5GnKlzu5KpBbvXhBi/+/tz7lYAgJ6
XbibuCR7i+MDci44K2t/cVnov7JKivGnlsqeqvQAaWjfHIyt9ybLvaD70dtbcc5i5gub0yYyEZFe
JFfnnJ0nn+NRpta+or9meDlmoA5U7an4GDI7z81pBaLZZnEKjk0fb/SMAQtr3TUK4ylvaOw9gXyy
xN/AtIVoo8XN5mJ1L9DZFNwtx7DfcgxMTFP+genwuLvBGT9ICR+2ZSZkVTSiFcCUJPm9Psu3XRk+
36ei5X8gTTcC/ZeZKW7p4az8VpbxJsttbSs59+BoptZRkUVYH1uvuYK3QA2j0Olus9WDTBnWq7pA
tVfiD9Yk87BZcrVuSVPCnVAq4Fm7QXjyEpe45v/lPreqJ/QWbpzZS3KA3ohXpoi6rGkj1VTCd+D0
2ZjykrzQIvT+d1+30rUeHd1ivGb9B5blzpjkeecxwRbOHRqvAEPwfTYOy51fZV3l4O/jEnC5TqYw
EJ4EMDaXV8BT0Tl0A9ib0RkhInfWNHegoRX/EnroqCvUq76SpkWUwYJoXwb/tJz1xwjQ5Et4iLkQ
04a2aCGZIaya3QJJYWH6BYugopWB6uGk2WgEjYvAHmR7yZAZAP9cDnQsyGt8wNahR+9ExdsxEA4j
2GYPBARQg9eRdJVlTKsF1hRo4Ye3Hgo5b59kE1n6EIBnU6CskoEZN3vfGpXrGfv3CKwfp7W3e04S
F87EUXSDPg8SlyukHoXCvngBL8V4fuVJkbRz+ELAR50V/pEujDl8I5jFwF69iv07d8d3mloS5QYU
TZ++TF6ABr+gqz/xenWZ3IcUMwLu1mKrSN/O3HL+JgWYm0y3Ucvr2AR59IeUM157i2EkWA6DNDXm
4o733xk3dPJAxDqVyePgmsr4XwPX7ZdJgM7gr/0o3AXtLD3zPR7bar0f5om+wElxnSACCEIiP4hQ
mRs30SUrmf2aSwEL6mz16OxhSSttZaGMgA/Y+5kFW5ehp4LFrZXSL8EfV67LcpuvQ4HVt8DoDj5A
i79LgmH4IXqH1H+1ko58FAjmPWhzkO3+t0TK++FznAxRXFB2NqbdcLkzYLPn77W5ONzntY9II+bN
WlJT6CFjEvnk+fAqVyX27cC6H+xTbT9P2FTnPlCND5a/FXh8CnquS8eRl5wP0sm9dTQKSnG6JdAN
LY0JDvUB2kRoumbv7MYLryiWorbSZwKySJMtQBwIiLU4kIsawXCSk6/o6XeyEPFGqWyq5/bcazzE
VeCGhDkUAb1xmOU6YL8UMx9p3tna4wU6hHtvF7oHtQ41S7PMUMj8t0+Tyw3Pp04lTiAH5bpON4kM
xqhc36yTIq1uHCY6ZPzNlRipyQ9AfHaI40zzmDsZoTOFvCLZxT7JGmF2RRITAcx5z+7ySb7+lzja
QSeaDT3BrvNd+lEVuEAixv+wUkA3gzXWNjkCQZqc9DmARxfd8jsmOAu8Wc0QjVkPtqtP1J8NQGMt
FAx2GG1fkjrQY+Z0UTG099ho/291u3PaxLwBtFfy7InTnRUYLSkIMe3rWHGEyiCv1+4Pv4a58O4z
/d+Z7g4/TrX/6xaW7zdVPbWUVNz0q0rCxsulpq0HSch1j3JmCAnws8XoAsuuDCYTKSP5gUWYIPE2
+rryetvlSaafqxVNHy2Ze7/LQ6IIHxOFBKmRR3sO16Z/do4YjfNB00OnB4ja0Nkk/h5Db1g2Y+8r
5pDlJGXCu5yBbQOlnfqtLCF1+BzpI7gkfrrYWUdl4ZuyHEOIlQj9MOb4VXlAL0u3TRiXwc6qBGLF
wy7lKtxfJZlvzH6TtnEZ+69nONjE1qQy+ByrnucwwAUIvijz8avKN5taV3pbg+KnWjNSr0NRIJLk
/iOvi9d0ZpLnN+oG87rxWnzzcdnZkGxCZ41Z3UmsphnRfhNiJ5P9b8ixW7+vEe5m4v1l4nDKvTuJ
BJkYdzYho2auFHYLvQYjq/SckfuqJkYH0i/K6IBFamPvYkuHx/q1oSzrsCUW51Sb2LCerFdfV35C
dvtKVDS5Ho/2j06MSYb7go+FyU1Kub7TJgV/x5e+e5Nc4SgstMjzM2ZtPXLUrWPXmD8n/P2EdwHP
iKzTOXGEdKX9gNQc1Y8Z9oc2Y3TyyheR4m7nVrMDpPMptBcND406tQbkIythSmwKK7D0T+mnqNbE
gMOcHJIVURnl0moINxYa/kayRozBAx/wkajD6zTH/8vo1QlVthAN3WP1+zkUzCtVEINJOs9Glvkt
TqlsFverSXRcEqad0TiufW6wPRidedWGVwR2kXeZDJ1Oi0wuJhhP8CY+oERV5iYRxQddLe+9spYk
Kp9Td1u+vzCi2y4qUbOJyCPUAdilZ2ZiFy0/ldEenQdqsSvJKcXHwU++PG0ZnZPLW+UXzboqB6Lr
r8QthfRxhhzbdOXkxcDvPtoBeIzOG7IyJwtVqAGHbS/M13tq2YUB+mP1g+CJrMxwyNjnAsS6vRvu
5uHUPPGIkR7aaN4OOzVNQ1N5WpPMsia8V/65JyTccfEBXyCb7laJTf4iPH4qtGld8ECTCtsYxygS
k8e4G3laYgn5Mad3YrdxkbWDyAWvbi8hdRDiaS+JZrRrW7uAt5AmARsYiAg+I4nN+qvlYF7n6stz
7g8fJ2M2aKhnWaiYpGe7LicOG89lpo8UvvobAylya8xZP6ZsUOJLUKEX69kndLVyywG5nVIi+5r8
tsJYmGA0TAwKC6tuIPnH+gOlbhujulnlIvNS2M22KE6VycMv2eOQ0eQeOxv1HzB+Lmz0AtATtqkK
aeyO0bpqcCvT6wIqyoCH2isXyZzG+o6HpyvjeRNem33XFbba5scDQKrdpV9zHvjqDpnifjTU/AE0
jskag9jIvLBMAPHPFaJARoIDum6NYNml7a7norLu50tLhMii+/htYeQeh+gRs3TEqUQu8KcHKvUz
S0/AW9AVT3z0Q4Gporbt8MKyC4GprfIF6hgU2Pf7uyt7fMJcsL0ULWMXfFUDQCjdkxGujGQ43PmW
S8HNYGuT3OTVS6gTkeLSn4gmm0Ix+PsmfH1YAwXDPg8BF6jjdxes0BEs6MN9VrnTtPuIz5FCoguo
xxTm6j9+l/g2kPU7/+g85TbtT52qvMRMhJsMPT63OzPXcfpcFz3Z1IErqOIkqoNyZC3luSGrWOnJ
QDH3RSP/5LnQDtSCtoNh9METoexboHQ/033MvJnk+y5CDkxrMbtPiHWUWSKaFWVw+cpcW9Om+SRE
BNeSxbq19UEhwQOrLHQD00zRG4OVAmx6Yz885E4IFJqyIy6Iz4yjAnqVTAFrMSOGbxuauf7KT5GN
QAm2DM9RG1/DMBknNjXLr4yQNMDbmSsiHNbLZjfyyHxCQxJui04i4s7H92Id8jrhCd3Z0RCrHesN
237Bi49iDn07D1ax4hGsTDXeFWhCeRBvskOudnSMsFyzzvgaNsuHCs4sbxtxrQI0iszqMBE9cjCI
uc/ZSD5h1vo7Ms7IpJM9O+c4e7CXtH0uE9I1wc39ZOsh2SZ/aJvQA1za+IZqwVKddVjihzi/BDhQ
K9IodbXxqKsthLL6rZnI14yA0ZcFP06lOOFi/myY9/13kZpbkBx34NdWrxGb119V9rIOuYz2GRjo
VgVbSR++QaUN5aT8V0k2HH3HZhPk9vgJbdaoB+EuJn8T8JhXzrH21GVS4zxGup22TM1N8GsJhzVi
kO4XU+6LEj3XpLJyPg3Vv5XeSJTfyahU1RcqgpfJdtgp63wq/e1MxgD3blakv21THJI9JfKk1k/k
SpvYdJduuzxpg2mEWqsKh5ffrrOLcviZaXCs4b03o82VLYVK49v3JojLVbsz3BWcAgak2kaRK2pr
Kpm1t52V9wY7Us/zFJA6jnWbfmpj5RALHHnxbxPuWFiYHrtxbsdrlbU6wvExZpFSqCJGN6PJOlw0
G/0qq2t70xjqu/x7WOFyhilIjIQ7MaEkLUGjhA1rSJROgshnFtO/x/wafiadOpIQyQ40QE0SELGW
2Dd87BlucejNmtzQ/K2tpUtzottYr+wz3FHQ5n6PMN8bVbXet5C7u7+m/beSw5eqRH8Tj6zIQkpi
TQTt47SxoaE5rqbesd4uVwfcLFlIvQh/sP7vcwNSXq9m4/mrWb8otvgbVLQlvJJFpfGRiTSmFBnU
tNm5pV55VIFmcWSzwt+DAbY2ZYex/rauJkYMvv7bxJnVtoot1llVDLkuo4o4UCMC2sb7GnJ96M9w
pLZY9Kxzy+e3GaJ2ro/w7VTR0UT7SPYVapk5c+3YgZBSrUxOJ7asB3Cvyp0pYn7Po7oZ07UCZZc8
qt2q7/6iYdrpQaK/2JwjN4fdzaHl/ow66yhXJQe0FT8+WyVyHF2Y0AbshSNLSAXV1INKHb4wsEOg
B/Vt9TEf1uAxHCi9MqbX8O3I7QF/PG7oEgn1KcDeqbEBZUHuHTx0fogB49jYIVbPgh8Jpx7549Ii
ouiSkQRKsm7TaIWJnbrZK5a7Ip72sGURibwh6BQoBHLtazlLMphRay5/JbyC/NOnHh/iYGFsJD3Y
GqpUcqxQAhEof7ZaSKlvgE6F5dEZZC40E6wWAG7GgdnrE8UG25EhkxkVjVlPNAG+J6SdPRYYwxKa
99AKezI9b+F1IaDAlzdP55ONbuGNXaAUYyhnEFndmx9hS/DJcBmBpSF1EjFtIQPwQylkrzKfDKTV
SQZcMhcATEiQB4IjO/8pcGy5fRpip+3VeSRdA8UFFCryGIp1Ky0zKDUxZyogEd2shlY4iZWvxOWN
3A2+9gV86q/DcsO8P2OnOwo0ySDoRzixXVIOGdR4y6o8y5JQJ9/zxTMAFcfUWph+ShL7MUTKJ5J0
eaOctF2UZExVshllcAYyue3aD7Z/Kueay7qWD27haZU+3nGlGaW4qoDX2ng1rIHwxaXm2sQgZpdo
iEjx9Zi1vMyZJ1B1Od2Yb19q8dsMoaZJAv23I5awY8FRxCK4Y94LKj7ucUcO+paQVruHEehkEW0P
cVmBuPj5SJIzDMvI5KQ/7g7T8iwkYSeQqLq50t1WTINiiSUFgDk7aEjGdKtnM0oltI/ogLGh8mKQ
goXhE4s4EdyO6676R9/82b0LcdpyTO+RYZQtjw8N4joQeuEkKmN8Dpl/PM+qaTRHRXr1Sa9C4uK+
TbN6ma/OcvSP5hJFavqWUfaGUECnOkf/VfneDmrt3ci1ceoExcUQm1Q20sO2TDd9wn5uzPXmVQ77
KqrMIJbk4GZINx0O0Q98LJOjxeogrmVNViHWiAHfyiczoEI3TfzkbQoxvS9ksbRGfj34lBzUidYd
VfD1eCGv6K6fk60WdIawgshBGoGB0M0G+D52d6MM5vTadTqhG+W9/M5leSlDt8S8lpCYuGACYbBm
e+uvCcY6k3j+fMOe1lcMBD6bQp/A55qRdYCWjmCWhpYFODA+YlXX7NfWDNC3Jelpkb971671BQ1r
reBo3ZaDpl1/Wv9vKFVTNZhUvbdwGXJNFcr8kda1KPGYrzrdgfmp3uEWHn4Ti5XCVDHv4CZsahll
AXKkouWjeD53/Myd6JkJIzgaGPkIpJVSWjWrOpIaJgawBAndmN24mfYKFPbhaTJzrER3s8DvHaDn
k2hP7rVpqH/nOHPBy+4MLrKu06u9L0Hw51LO7ssBnhg0USIPN7kqbVmUYQDzKaYapL8N7lUMIs5X
SEIhcwUjA4Xh0wFm+AifIMYbibI5K5YA6PtO5uoZbUt2t1XQb6zRo+LV3cdepptR+cykEebqh6dO
8OwDaumK/jNuRD/QCKdheQmekF9i7HMPsaamHGN8avWZxNBn3e/4EIJVizHoINVLLBeg5Qwm/lY0
suwQO6THbEaVuwRlPfScOyE41ydhhG0mYUz5kntdSZ9pWEOXv2wFstTUiHUV28+K5/WkFTOEFruL
++5L9nY5kcqrPYRjP8TMU46/yHNz+Ti33gOvE2I2YXHdYeUR8ENBwEc8eE35qMFaxROUlTvf/db5
7yit/waFCr6KsHSX6da01lAlKatyi/5GdRoXYk4RkFtFGDvKxvozHjUL3Hj6WYf/n/kEQi+6rd3+
j6MCVKAMJ1RztCC8lcjWUHV1XcJ9wtaTGlTGKi23NFPvhsyPiUhp4j15EPcguhbBdcMxZd3Qb1P0
NAGblhrWA7q3fmUShvJCsofNF0B4/Uf0bEdZ+vzd7jMsIYeeUM+Mc2uoQXT14zjmRIDoG3VPCWs0
1GOLJNLozH5ZYCbACWewhks46hRJjL4dA+sNBQTUhoRBL8oD/mEtOvF9e6QlDt41S9RfA3s9F6hf
k3IVbyaEzs59SxNixr2/ora0jshcfLNldti2uMHkTXpkDmx09LVDkRXhkOXjh0Oq4y/8FJDWumYO
HLGf+xnMFhlqUNDOVbh+LavLfFk/FvM9ONjfaQ210r9MnBQsVaCmBwTYS1mgp3Dv97zA2Hn8gkae
+7GKypEKGdJOjSI2es2ytSbb0u2F/Z6bn95nS/mKIV9cg4QMAVu4XqfjS1EB8xSO+WdaeXGhHc9L
0ceSzlzMRWFprqEkaEVC72YEgFy42TMkc9c4VZKdAN5Qp+ezVlI+jmfkFbknyrmkIY/hLeDAxulz
TkG2ShHrmSeU2kReMIoUEzRW11H41lJkQPcgdmuu0nY14ZYP2NRW+EGy9hKaUxyymFyfOKSTIuf9
LMBP4unIaU7bcIwQ2/7GBUAlPDgrZcp19WGP2LDV8elTjZbFlDXcPzFAev7gjSONxd6uxbwswjqD
PJ61rdH0ueVaVCRoeRU3M2eJXuUteSlpmW3HwV9lg1Vyzh8MHaPgQ6h8hA45Pp4ZGh7SAOnNBDx3
9/d03nekOF56Hx/iG0mHWkhMmteJUlQ/CV/2TFid6tJiFE96kX5N53eqMikXDKReBdUg+cnmT9xx
H4ku2p2QBSaIdGTh94mOog7RkJElHncRvnN/dMnlYQUxcKIOTsQTcRqCe23Da9ETldul+K1ijZwc
Pa6YKCZD1tef4PISw63REikR75bkishYDWe+A8RNtE0qPdyZQODojJ/F/euDxVQyRRh5HRnSG9hr
Il++w1Z/Y4mkXNO6GdeNTi8YlpxjSqHpGY7EckJJU5iwP+xp/lMrDKNYXWXTj/LCFcqfaV4yZ+jm
hkApYHG3f1Sq7Ef6Am0e2Jk1XqpG33IwJRlGO955YVgaA0RVBxhjuKaIJ0WtayiKj5gV6Cvvla4u
OkdfW43O65cwusN3X4Gk4CEfkC+XQDSbSiQK1QeW+8cJAKKmMIDUM1kwq6f+AcTrv7n/LLZ1prIn
essuulOHYOtEIXV59wgR0ye80T4uWVEjJsS8mikddv+rSHZNXTB8Ni1aYn2D9wM0Ic3ebkXjQD3d
uOgYfVi54FNuYU/kaJSpcL4BrK9/Vc3wer+fv5ch/1fCpr53jwJH3NbT0cgAlR2Bm/LA+WY/Bsoh
+Z4H/pWmtFUys9A/eYLDw3bHlP87gNEft1lGo+ZYHHXl4jExGD6kfDz/tU4F/rLQ7hZExTkfD91u
V3+i0nl92w47oapmlY5hpeh6kj82iTDAo4dl3jjbrPo3D3cX+9jfTnnZi3qrokqNT8+4lHibAaUl
EjjTLAvZrtTrFfGPAvzLVsknvh8QlhTrzorpnxkC1/FnXlpKBj77un2vwUUWrQlXdusEPMQy5hA+
xI1DkzropeWiV6iMhRZXokRdGcV8mUE5O2r/6EeCiDIMjBjw4Po0WhOq926GJhQaT0I2Y0n4gfTN
GFsqUVrmaFottQf6AzzdB9Poh0Mp8WeKp6Db7EbRU1IO+Gx6xTH7h+xj7LwEyKKGxp5zkK8ARIc8
Om5IYR4QfSJ4RR+CeLjcrktZsu/NNCOoeNwFqCXnNtPBQ/J0fS6HdJckVlEgKFX0UqXMvuAhALQt
kulM1+852iShJRuUrpFGvHjKnxiDc2HT6HOzgHaxlS5Rm7dQPLTrBUFs2ro2wzoVDLueCSXBhVh6
NYhtgItdzPHHeoew3S2rnE8xdJTR/K44KGy+SF+dGf5dIkGPHUfAgFZoXqBF+53jfRju5v+l9An7
Mk2cgsROvmFaV22B0raWaCIqrMLBBLEX0zafEkZ24aBwD2pH6ogJTZqQZ+ZEQXjtWF4m5ET96ksE
3VWnL6QhLg7gRU3ISTH6DV676u1nU8fXZ0EKr36vKURqMJxeFFsaFyeoKuyn7TAEgEHFoPo/kv6D
BuofCu/Udia8+Kr7aFDdg4pxQRajz2Fj0+V//91k7HlpSBebDzPHj8U47pQf8IY45jPak3nUKqVO
ycKtbYtp9a04Boq4ya/Rk5arLKg8OPd2dsXvqXxCKvHh9yC/gvVqkklnEV56X/H0uiOg5hVDrgtY
mscVv5UEO93VMGRKWAOjFSwc++DZ9nVBrwxoQ7WN0H2H4BxmJLmRb1bUv/ECzRCbBCVhJgO09yDS
nmLKv3pMxbP0QTdTA1vVSU2/8TT5xYFN72Uhgq23Oa1yWQQzJK71pIszBAc0veuoyqKnbT1WA7i+
nuY1JR8atLhqUyc2xPll3aSF7p9WxFNVJftkXLdGru/P4ARENCWmyv+VufEH2sNsA9Lo4r5TIytg
ZWoWUWwJP104aSZWCGFYAZ0JnZzViMlKe+iPg2Y9BW3so9OSydyy5REhCiGa/LaSPbMe8JWUp71B
q3Z90VOHTaHbJWMkGTSmqF0wN97TbpiGBA+nkagxTBfrdpm4yk5vqmrg01vAmeFXyFDDGPY6N0LC
2hdnVz4fnb0bc5Y2sex9xK7CFSjh+FCm211vv/M/hkL8iY8WOVbRvDCzYefDhVO3ZAa95ZBX0uK+
wLOBHv3+yd2MJyfII9Popz56mfD6Kd3P5RiBUI+mfJG2p6gUiHnJGwM23GNVV35LtvUjWu6unpSM
kQFRIiV9ZhEBsePdjWOGjq/EocYHHdAp94U/6hVfQTAOTqDfLO+wBNRnh/wQfQCGFaRC5emrk/HG
k0WDasI9cZ0+2+Lk8GfXgUzzHr1z7nZH6lKOC2kLJGrzhhH/NyHsCf3M1aTwTX+jFT02kn5kdQ63
wmilpzPqvytbOt0SEV5lN/8r8Rti1heaQ1m0dDhKpemHqVRRoi9+UVW6ru+f79Kmhh5rR7WZfsPv
HejIS+PL0Kz7OuUBChZYB9NHwVYqbW2iijUCqcDWMbsnhS/SBR1EqLhB2LoXnbQ2CLJhaFH1UGZX
m/JD6aVDND+ObFzgG9VXfFb9TAn1/TWMSx7Um5M/mhDIy+OLViwSDou5G8nzc8+owB65ztl6pvmK
LRzFq4HRBNFO5jvKkWe4HNZ/JcR8IPKA6pYqJkMvxkZ9peILal6fTBwQHhno8hbMZyxsiARpcVWO
tKewjD7wGU/PEFzFyLXfUtK93Xe6vMI2QGYVx4i7e2hwONwXu/NEYMXHXq0fyx1PymexkPAEE7/R
QuVTtgfXGDOgFAV3qcbpM2DNQZmIiNmMB7j/CFLWiUsCziWze3kVVJvIGoUxU2VNQZ5vVXXypXGG
l3QhxEqW0wKX1xH7Fl9ccNQzLFf/NuDdJ81WfAoUUCa535a4j9JahRwt4hrKsgACSi6Ma+UM2K8k
NRQHEcW3flaXfQHXq9jv6pM0QOkk+Q/N20uetw5AdF2EIm/h7WhWB3q+MSrMDGAtQV/6f2dGQDKN
/vAxp1W5NQeN4HaqZj6QPmxmioJEIcoBg2UcP0BENKZaP+IoqY4yUuV7eyGzXh3GH47cgELRI2Um
V4EsEUX1q4vbUhUzGNqkWhtwLV4yidceQVufXlVfNZP/TTZ/IYbfw8yPgEAD2NieFmhBKlCYI0tq
EEtLN7vKlw5Hi3oOkZfiK4ziQ8z4YpsfAL+5w6MZ2+9Ahgv0v968V3UKk4Q5jYeFu8lr25eDzdI7
WwhOJwbf9DVgzJ+oYjnh8TTln5f/p6Mcy6juHlQxG62fnLiX9SEldPI3b01SMJLzO/Aw9O8Mnlkj
t79dAzUtukne3hu/tKyGNBBYGIBnkv0ODcK1nNOj81VYVxou7EuUNLMLLKAckL6T01lzrJXF+Ggp
cB3I/htMRI9UenK20cTYRWvL423QYGCfQpQYBehbXQ1/PK1wvWqXS6+bS/W87Nv+T5nOO/Dwos9e
2wuSe9+wEiidWsydU941VybD3nNklLZdbDZRLkL85mlmftMk3ppZgg9cTHneRprwIBpZJen/pc+U
hqDWo3X7TKm0JUiW+bOZXhv+n+2Wfwn7bKD/E1EXmyfIlliMMHFGAUQiElyrJPjcPaS2SVUM97pm
iUsL9rxN7MEsx3PGd2bf2nx7u/uiiYKw68OFrvsO7hsRv5KP2RGit3VJ/lKWOvr5Oap1LG5ZSH/Z
1+l2uVosX5z0n8A2eJi8Jnueb9TAN9LSA1YtjVQlRw8P74qfOpcCdFWynBYthygfwOPxWXmfilqQ
h2PQypJLXFvRbGgnR6/gapekbmFg4YHEPKDlML7OwDObMeSv6LsqnwDR0ZyvRQ6bdS7T2plxronc
yJIOlBVGg0y3SxFgLHZV4miZXO3uzsBh0DRV2fdd7R6Bs/rRSj/xoRwdekPjRWzp38v4GxZBzp6J
+HHvt16TuGicOHmJ/dfGH97qkCIZ84MNAboXqwCuKYaOa9BdfgUPzjdq41ASZh3cF/Cx4TMrtm5O
8IZ2JFBKLapIDpqiaDZK2UHtrmQMtJd6g3pbmBYjsQLenOXa9RGG/A13mA/0GekWemJ4Tr3mwDdC
6D2Ite8wH9Pok/+p/fZ1IjaQzhs/xdbwz3UFMlhZu8HkM0HkQpyoh3rxDdfsaSXToMwdi4aoePrl
jv6hhMv8NSTPFgitJ6iESCv3MbMIDbGkqgsqImYdmo/U8CjBJxk3d5/uRBqyBRM1Wfs5PZFmkbem
25IOD4vY1Cc2VAkC7rKhAk0nUdszX3OESbxz/XyMY4t/qQGH5rh8G45h41860Jz17mQlucS4Mgui
eXmC2jHmNkuHi/WGgv7YvkBE6N2qwEsgCgkVGiKmYDJF+MqPjmxT13dyBEw8XuEeHbzQTzjjHnsf
sqhRcg2Ep9Y3iFhyZwvQ4ePt9MCVeo7QnjLx2B2e2hc0RTAk4ChLlGBqfFERryIWmi/sjSMwSiRJ
IxWdK7AerdZoFEI+r60QWMW4rSyKBaAHWWX1bpQ4BGVfvusNjveD8WEwdXVASDNF6H9E2k+14/0X
vYpu4D6d+2vWeA0EVdpFrOfAmCEj0wBaD+46sAb/K2a4rob916IPf/4aUmnEyhYs2X8afkni/fAh
5fMcFeSg/8dsYULhms4Pn+w4F+OMEn4myxGClJjxtAkxMwfR+MqB+ZG62io1PIX437MYcvxJ7g6A
OnAC4ZEJ88pQwPCRixFudD3YDi76jS8ekxwzQ5+LSXZ/6Kbbdw4u86oBNwELR+mSVddxlHPMc+dU
Y+a2eSEeAgFko0k92zfahYoTGnFPPu+BxGgIJ7torqqz8d6W+gVQ2uWuU8d1cIWjuWXnsHezXfjB
KRjG50bSc5UacITFGM8FEuqM2h4qdXIfKjpgwADkERe6W1iOm81Y8Dw6YFw3Pro6HazJb3/KqXI9
QtfnTQeZpuFVCqm3/yzLR0mSSOeFYFbKztV/fN1Y91Rr1t6ACfKkEcPJrdekUDw0iEJfIEGa1rC/
6t2EmZDvfV7tvHE8R9KEZ8L1xoWHXSpJ20qPQzh1qKyFUbZzcdWIv9zyjvCD7v9ZWFJygqOtQms3
unIKjwA96yysaYfWv63TonlUKoWdeN/mBkehIdNT4oRR3Yj7S6w2VHYW7HCvQWNm/rwxxunBoL2e
muZJTm0Q5y4c7a4Tz1PjkB6KhDbQJUGrtLmRUgweTVkS3eFiStvc8l2F3EGmMAX/L8E4ufPYoXw7
Bf6gqFNaVL3v9+gVLtbAFcHMGNablzcrepFhHanVfDU8Pb/JpHFpUg0YxJceV7rtJxCrBhhPPCA+
JmrFKtgwR6XvnGY2xj65zuGCkjg694NTDQjzK6DW3ZcruiCD2cXpiDmR/4NAn9zNcvvrfGSNrPLg
PiXHQAZCo7ZEvWDrV/WFyQHpR9/cTC/nBeKNGutGIhyHfZwDjWFp3ux0vw42hMICZFSWULeeMQCr
dNLzn+t37wqJl/bJDyeH+pohDlWHN/G5dhlc6nffomCtCmI6DkFK0TBH8ppyYdLWsU9Zw9BSNrJT
P7Q5oCzK/Sq4j9U5D+4lUNp79V+nDFVNyfcwpl9QcHRglCOWsUUxhWYr55OZESZ7dhxhyA374Vh6
BQdCuB9v2RBvms0seQqayokFGVKvPT1DEpO2b1zs87SemzOgPrVCemi68P6YYHFR8MR9NSM4E2QX
rWkfPnah2aCeMouEcHANIGBHpQWTQmvSuu5Tr5gtv5LVsS6xFy8bM2/OCy2bJGM8biNOm2ZSKN3k
MsTu1YhmYcuHenHCkTfwf6RdGVl00aZxopRbU72J54wS1TmyZvKZ0rxpwoXoSwFwEWGsihbiXnBS
z0UiScPQb6ZLeSZZ9Wk7Izy784l8dE3uEIntBvmlgFUEHJw2DM0NwYpy8mIEB6AFi94qCKT47cgE
O0MZwYPelFKpoQLV+7sDqezsacpTXkzrutcQsO9xhE0UxWhVKOFRpnkho1d+ifoDYWaHXEpIuxRd
7BURP4XgfbN/YVvTyLvoCUrll9nXC7TA1ppDLhfm0/irFcDhrdbn3I9MGki++f//NKgd62EUJkKd
zaHy22xsDgBPY5m9SRQjUDKLmp8RbaDe+TFtUetxIeTmEycdymfRiX5zJ1WJHXk7+S7/+9caAQYQ
ReVIwGnJlQBl0r9K/z4zoRIuk52HBmXw6ecyOYZwZUQB9j94/CiBQNfqGNlbOxmlDBBdbD2cC8sD
gt+agLdqauN7RH2jDuyMRbqirsrvKlyI83NA8OWGHlYPduPW7aNaA94d6SjHOOE1SlHJxZ67xhg/
Ca9QSSGCkE5I6U3HSfwrz0OYlkXEPoWv2C/mhJQKle1XGIby96bSEVy8hG7Du/SLjR9GxoNSScMJ
7RENAJ6ce3tnuY4eMtAcrEnEKVm6bGLgDK/VpV8TEJGwlpgvvD4xCMh4AwbDNKNjEgXyhbFlOqCA
SZ9U3OGzUnSCU5HwxMmsvSVjKxA/45dUlnewnHtJtlhJvt7/NfgvIJSX7FcSt5ajc84AXQqpEJ5J
NMQeIswXA5iGaqKeINmsmnhIYuzs1KpdU+PUFNosBlLpzKHzi9pAFrX8ZX+E3x5K6kDD7/tx0hHZ
lbaqqvO23XI4RS7Fuk4p98w+jqQR+1u5slIC19CZUq7Xr5x5uw1TXNWA9qOs9RIhDLsBkgkWlMqC
M5J2DyyqpthEuJjQu7WYs23296fSZsVGcx5jr0VnuzOUciYR2yQsk82CxaC4tQZwU+LujXL4D5sg
xCo96y6Lo1O97WViMqSgtl5li6uWYysKnmcIguynZnZZKTBxna4bbfXfRq94xq5QSnZH8ATZIjol
TQuqj1Gcr0MD1vPV5iScZ0SMWeXS3NrH85i8K1DGY4KC7R5I0erQVQbjG6adI9lARt2C6OWKDnFI
u6RbXDGGe2IcVyuxKvjVSSbM4Dmu4beVufS5G2pOlsdxBAY1D+ni5bL+1VymIBEQMd3ywEKY4WhR
owf/QuS2FUY4FXu97n120gpidTVMJ+V6l2S3vnFkbT5IjMz6t/Es06TnY1CbXyeeBbfHF2gBTLNl
6y4axaDnb3yYaDnxnE0yylpy9SqSBC3Y5d7csG4acQ0WNY18wOfT1V526gw+bm8TSozI32liDObV
Mpr5z1fngTudaH+/7/7Qhms+8agyowaLaVpgAUJdRZ7pYrVqXgzHG8m4Q/HZHbS9f7/xLEr6YZDt
E1pUjG3ELB7NYcUf894TczPBVB3ABvB2VvXKjjmsPCwmZVFwogXvBfK65SjIz6jvbSkRLDH3QDeA
PWd0RwBwHo30pS2dFJb49TTXbN1x6qyaqTU38/+zgVKeFCR/KmZqmR1ALB7IgMmnm9kTrNw7dU4H
CchEOzzr6kCLxXw8oognMnAMpHmisyiA1X7q+G8sHFJIIrkZTjhVWScJtAE+qi3FdBZA5kJ4092z
MJn6rkBpMmYN5n4W1yNXazZ3IxTizEF28hekSprU8/DKeUEv8mF1B1ULHd/NhFQi+7FmsJxK3btZ
tsvfYqkCClAtFvupYdX05+PTVipunpH0hciFF1LRWm/kJB64RZ+wmAKWFIv0SlPMmYGbywqttLP2
yUlPhbUa2j1GBV3Aqs+PNqgdZ60g3BmxVZ+71Oalkpp2y4AndZoFt/Gr+cnIY1lz3hs+bFqO674W
kP5YT5/8qFpcd27t2gg7S2DAMA7j6Uv35JPKZEA91RC66RvC3tb7VxRMYuSF/hIUiVHl+FM8erlP
ZyGgTknx73ejGlrcb3sOldbvWSBA1udhKTtgeGuxsMr4TiOhn5VOpmdLxa+4Z5mKbAiX7MJrtrde
4vCm1r0wqIzYQAy4XB8+u9ZKBZsb2ZRDZ3noTSnQsy54wjze7GHg9GX/33k2IEzbA7KwOyb2sBbm
+EMzjGAHFz7IHNGCYDi09GIRBbDXOR0RJ1wb9An7aYpoYpg+5KP0bOfCvUHMsv8iTEHK/UeuTWOQ
9VTGvsqYDixBPwINZPAWhUBXnTfLzc6UjcMomJABzWfpdctXFWshM/ai9Dv6eMusJJnJErw2i1Ge
sxcz3v+xMWegMCdY9DUHAGm2SaNsw2edB0j/qABsW0G32qxgiG3kasisFdpQGy0XhHPdhPq1ZNg1
YxdtBJj8r1A3or0/GbueAphWfWgwcdRmc4iueO9sa2kfcl/uxNQNWG88m08dFWFLCMGRX5T9RXOR
PILx3O1MeoNNr4L23YaHw6nskUK8cKMzFn0w8bb+AzhU6cCS6VZ2CL1OYO4JS270audck9mbdh7l
t2DbogfS6ka79bLRkVo5Ni9Qc2y4XvO306PMioEWDiokpiDD04FMtE3RZAHu+dVf45hwPZQ7AniX
/U8g6K7EJJRcWj/3zWXNGwlBbmq8KZDyJXYcl4zupruPijnn7RowDL1MqVtFKHauZl3q+cT/cMnq
xZqc0nrrDU8rKkP2srmUL6TkSrh8VTsAMmPcf46PU1d2C7e92p4+Qljio1RZ950G4ir3/rsHdtr/
ea1QaPcW+jGcmxSdnt53t3MufeD5RriEnbbdb3zP+J6qBUkDbMTP1tOQ+2u2dTJLJGZWQJf8ZRG5
Clgv8rL/dSsA+IFyNvU5RyYJNsc7hmXEirJg/zM364xaOxKEsdNxaar81fqsgis59Q+p91kFUsm2
YKK/aTufA3hWDO0rP9RDRY3MGBLxvaCockL5CTa4NQrVlXQfRXr22jl/w06wsPlvlSa3FdWjr+iG
NnviDUsGSnqg8wTIrGZe/nk+bbljw/qEXrgKjAtpIQKtIeEbFge0tf5x1UbJvKFJhmT9shUcapwf
32Drbmgw9+iGBSm6tHG2Pj9EiCJYcqDdCWkbPBRDiStGTOP5Mv4ivMxnVPJ78kC5voxNc/eYV3WS
i6wXvZcG1UrI3DSwnhYOSpKF6b17csvZ/GDjj/kYVaCXEEE4CM+5CaNz+MjU4difim1eMfnEB2Ql
D7XDwkVKRSceIy5/DrkSLS2Jzwo3WxuGmVH6rit+R8Ghvdpdg1LD4F5E25YwsJ9wmbn+imh5Ov2k
qdCfl0BpZam2zS/Mcj2lZaAM5XNzBfKTD60YqMnC0MPWVz5KOLgUQZRvE64XEEUdrW4AbJDd3ZZi
X03wRYiznJZsg+oSWxjyrBAJvFfqC74MPdVQ7i6BtTt6B8yDw/niTMyXuriXIIJnNiNcySUl7QDT
MbSCjVkcHQDVGhgHZcrBbAtXfbl3yH5wQZ6OkQKGitAAQuH/qB8KXAfDmrXdKhHtvpJX2MS2mwOP
PHrr/duQpsyW/TNFfWqZVOCLit9XcGBJQ+MrQEJlicNk8mzVs0dbCTVEF/XvCn9Ar+wyQc1lZPwc
a8bLSeRZ+0UB5bcy7LfkG9sfRTwW0Z+6JgTR6oqvbKsBdhgYPfvj9SfAM0xHvTtc4zNQyo3PU/j6
QmycEeYt5YRSW4/iNe7K3VQ19KGcX1cKK+rgYPrnad8c5B+PwZ3E/PXIK9rrWTQzNBcprn+ed0iI
WRADTtM4QewHMZzFGP8hDmENYotM+yo2fOYe39q7MaodxRMAh5XN7D4EZX5PtCRJkefigUFgeYmN
GkXgPwIO22pdNrHLaN4bM5zTrJXg4QBIUJ5ioCIE2Sl8XNMW/HLIOsGrAdMqGy5XfAZEwWJhR2xT
klyQ63pTA1ddHwOmJI9YF+b16zi/HAm/ML/FJAINvpDVI8TdbX1uysCGN0qdNucEpRr2BURnimX1
w+CXgy/6wFHo/pH9sOhMa5FndEhnX90td+eT4dPx5e7RfDehLMavuUD9L/Q5Ip1nvtTDMQOmIRcT
QbikmXMyBt2KJw5nt6NwasBe7FdzaE9SKVKbrf3OlQTBVOS3a76YTtA6YUVitnADPqNZL68ypdJG
7xaGmUkxH5N1/QMeRygz/Z8x7s98XCy61sX9DTZR/p5LqaU3qfKUt0DsFYo+81btISJ54izo9Ock
8SqDNgG0WPr+vhJ6yM70sLnv6oG7kfOLUmKKLXZFSvKbP5K82xXtSEhQXuM67PNAKXnFuKLRYLgX
2hBzQ1Rr6sgL3fsnh5ULJFSmfZQvA5VF7Q/osrUxxOT2KulG25qwbDIIFR/feJ5VKXDeW5eB729U
fwYlMw9EkaYxFoY3WxFfpz/H/kspBG19hHJHz6sxb3k7JFrQdfkgyOfB4RvduLMne1rx6KVb5f+e
YGgVnmq4zPFMgfXOPQP8DhLDd3aS/06vNz9HzwcQ1WLcBKx71VnhxZQ7g9/PT/dKSlGvMVaDNxMe
6PNPy43oX/0YusfPbHxWWR92SOW3hHY0h05VTT0VtIY4uW9Vw5PwkYpfoZnfnucXwT2GeXDH5xTo
qAUaSG+QZeKfAL8QaDS9IBEhBZ9Ib8ES2qOjVSXBHbgzZW8x5CAVYS6tXQvUfgB2o+bWyfTOv7UU
XiS9/Xm58DRVRt7q4JRFvxF0Miq07z0HQkGd1ifwdMPvbqlsjZNqp5Q68LC1+/js2R5gOncaGlDu
4IXXErlZDOUARGhanbbRLSxZxmOLitPA3l10SlQOwS209S9xJgNp2AASlBnV9cGUB1w1i85TulyX
COgHhpYW7jXDab4ycIR65g/KjPHmKFm0sk7LD2vZjnKQ/1IYV+4/GodsFg/AyhbjFw3lfm9K7uqO
jXrnPTWSjQdLhii68aCZd8x57nv+oPid71+SXVzDLVQDcWOr/AC7kq7jHj7id5D6BthsctQStk1d
CzflMsoOTElap3jN5VXjIaq/Yk4ALZBa+jyWRwL5RtJXp69ozjrPGC07UXL0pNls/6VNMNTQsncE
WzVd+hAwapnGqlmDQq1MZ/ZyZ7KZ0Ba3DMFqUcyHvBXVhr3QEgbSzl/+T2KpjwzBM6C/GAtrB86N
hkZ9C6bBBWgpTFiDuHv5X41Svu8oloWnHpGGxSb7xMwkKD+nbyK4JziFF6WQLlJYvBGObCU9Hc6M
KIkHeIPC/anq4Ql4a3wVKZqzJJK4+32aLfJPK43Q67hft52pfNzFVRdD91dOcoYx4ET1+2o8mstA
tCuvgi86gAuIIQ+fpys1htL2F7rUD7vjW1oLK9Q6aopbTeIgPDqMdlw2RPqiW5nvzLbbjlCBb52x
3BBQLrGAo6kjIXEC7BT+R8B9tRuMlyYK/EQsTsFvAwtBcqL9hQtlzjVfWnlDo4YHbVB9mFXcN7Bs
h0OsWldSS/ZX7fX8QewOASj4y6GkK+RsWvpT+4PcLONHA2m/0FSI+HPsHt15QD3B50IkiQJHsLps
173WKuwQlYaeKsQZsnQlKXWstnqTV4a+NextJRSFmOO3Yw03XaENC3uSXWBjZuNFyCNAc1gNja+2
nlyrP8z5Mdqd22CPxRKnE5WSwPr8M5ubXQOtvKRNB5vaMY9ZCMdsgg9Wykl6a9efBYi8oUgJ/XEb
iNXqhnRt9ODxF4s1kHxgM6qAEtY1iVh9oNKRHoytHp+iwC1imjdRYvk2SWGy7U5EYJ9haUrp/JcF
yrJXDgBU2fnq7l+EZXVA7cuSipkvcd/OJwdPu4lpNNA6jPecAsuM+Gag+5f6NDI09gUWdgoDDghY
TyuD3IRes2RgQ5IKxOOqJGgF57Lgj/p/5TZBAF3HIgVuiut3MWva3kP3+NutQPy0TMyM2uzJvpCg
ACN5jzZPwzIO+OyqArabtL02W4vBfx/IAq+GXOO66JYMU21ua9HahLu1IHbRxNN6R6Wy7vZtVFpY
Jps2h/Ah0ySz7cLVjGmLOway8Sz3AAm+sVw0nZWccirMrqwlYpYauKrEOjIAuZVbcdCxk84itkzb
eg+PnoQzvrK7T1GUcMlRgjg8VNh4HwkcJCOPltCH0q3QkzgBYPv9ZoIIdgSD22MqGz1ffo10nGK3
BI1vPMX1mTKEhGzFJzqfsj8iQ9UrFn32fPt2YlkkGey6YxtjYN+a3hF3ErQZEk3mQkXu5AwKJuVt
2y+uz4i/nN4npMuZDqm/i2P4fDDSYDfH3glhrb9GKS7ytIDiZoCICocFPIqEkRF7pOmOOsc7DmzI
ypmpeyUTeBtJ+RwH8TLtzZb7kONN3eATicS/ngzi+QxV7Pcl61BPkndT1lho3Tsg9pt3zSUmsm5N
8e8I8u+/6cezn/mbblwoEghnZUYLH39781AymGvobvJ1HdVksv1PSo43onxGhYVDerh4txoIcwWk
0WKScyqHIDL7ormhyYOggwLRlDWPDGqbQbIvQkZyF+F5Umz4SRDwLYpFDgDmDBlVRGsKVfOtCUWv
Ls7NOHnM8+qUmw0n1435jkCsPDIOepMqKn7r0K9+ssHBU5CsB99u+IoYrHrIeahPS53/ruuNphv6
RDD/Fbccr+bAk3Ouh892i6AUOi9XNQmMJB4Jr8KBGL0T6aCXaMwkkMAXgdUsqq9Pg9EapDew+oLa
qAMEn32+atbyxdmuKhWQNJ102nzidoYWs8+IJzxxaLTB/8fFWC7ADRvWYcJGTJaBf/uvdRpsahW4
pzcpI1uoB1zy11ucg31Hflr2ufQTbGGTJeerZjCejVSkAtTJ7GazrnZWLkjuKnQ7RVAT/JqPCaWu
QXuHaIT0MHd/SGd+40O096gRlc5Bs1NKxomW8WNNwpl+h4ZSZduS6T453RVsExGELKPb/0hZDw1h
+nGTWtS/yUPxDkftBteUMGFlDjxIAp6zfKCqV9m3NN1Ybpfdpz2Q1b5wTzcjlFjGG3aJstUCmFWr
nF6yv5XevK5ayezbawzB+0FVxD3lIgRzhVzUySHEEqWP3Jr95RcJamy/yB79ADwgWKZTTUi03OrL
hbS5S4CWSKZPUItdli5Cd2Crg2/bIxAonE8rN7XaIzqpxaXgDskZZcpI0Msn/Kk+XxjoMmPxu5dI
fOHdLskKwZkAYSfjTDQs6dpAuZhAxfqfmktA6BLw1TmckIfDcqHJ/nrekPEwhwQ8uAS+wq8IzTQL
07Qy5EihH4LESb0ttUC3twuNE+eag+7yQqtmdJrG3OWJBT095HFRf0s11qv41lv41pTvZ9uQLh6y
7JYS5f8Kpxn3mzYf76dsrwxQi54UbQcn2QCl1O13SjWA2rcQkanlnC0QPf7cJKvevygC+hWlN1wf
6glX1ihZLqOqFuOhTg4w0C/0qB9q+rPxXjsNIEuau9zLLxv0HEFAnp/uSq5yJGWty63K95T9Xbp2
pQMkH5YZtqSwbs42TlerVxLoZtzG/lIGGZj0pWA34U8qsadoh8bSiFRssm1OwuV5gnHoLm8F8hoV
I5vmVgFpqt1otc1jrskJX1oYPyyTuNaUCW5oVo3YydQksN6lBcs5etWp3ugn4VC5us/OSYvs3zOS
0kVbZ/8QJJyoB6H02m1aLWuN1TlQa/RqZ7PwEDmMDg8TQAKBkoivdJ/feLtrRkR6RINaqn3y91aK
pjWBFcteSBEZY3D6mRkcL4D/UIEnBX5rWq5BE1BCTntrwIAiv/9uF4h/ei0gOpCv79s4mI5GXO/4
km4ZcOEQaxNnBQUS9tG0CnQi2BXckZpjzmuIWO9BD+nJ6K8lZgYMyCzivtj2AJa8h1Dox4fiYkZz
StFQdfNmLEQMu4T2l8yM0CdtXH8EtK4dZzVmfhBdlMxA5QgzGn0iQJh8552oK2jJONp0B5eUxlua
SFsPQJog5CQq2IcRBLxH8Y0BCTDEZRt1LplHMY/1oerNOj8RXXobIyL+n9DHuIbwvBn1UrWMtJiI
3em4eQ35M5rpRafhEeA4xSXItjPeBsXVQ/vJY920XUqfa8dYdg7qWSfGzjCKHc5aguMOtSZrqhun
+XMPjgRFOb6BGOXdmRCtF7VaECtXJzXX428ly7yVl+YUHXPDOj0U+Yy31b9JiTJPhr6mjfaNn2tc
IRhkHib5TwXadeRthAhjSWwxAEF8K2egN972xnb/CpVo9GgmYkPSkeiEB1vezsd/vZTDdl5dA9tC
9XdC/XicZBpLwnAVE98Gzgazc04Ge+YX82bumkeVgCWqmhpZNEIlYX6/PtGSPd9LVBVqeICm8fH4
yGc9+BEvCoXQr+HgFBbRfkZkFH78QiyywDhYsEC/hsRFhJ4vHrwiHaXESrbiH5UR4S0365QDK8Q5
llZ0I8peu5VliQQZ7Wgc1swQUlr+Ii4VNLAjg4z+Al7Ds211xMCWLdGPW9zkMCJinoCSnZtgKS3O
WQ8JNgbE7Dikfi9tyudKMDZZhEtKKBU4HHHL+BmdUf8H0bAVQymuSW0i38lO8HQa9bj6X634LtXW
shDEhG6CjHCNcUGCYpHG+99xc9fwtiJKNmpYh3iHABqCNogtBJevOshdHydpnHR9gq652mdrF7tM
7uzOxtZ6luyQJbqkRlPAJPsBa87ct+Dj123PSDJGvX9Hkkz5OJ+bNRoM/piBqTTqZSZ2sp3vSebm
2gbEFOl8r1DdVDB593EygNaT2l7QW9YoQwN3BRxai+jYh/qQ86Nh62bc6n+YvJIzytP6NcbYN/4C
sx8s5/NnoF84Q09O1KTVM9JowLj5fYP7eWUKYVuDCKtTfxwYXthvTwpOPt03vC8xGUmdM9usWWJG
8PN+kCFX+mf8zxm/BD3A+fbJELiEQuXuumkT3u2eUAcc7hDTl8l94ijie2d4T+asFHoxbu6c/S0s
bRN76f51tBNDzJJHDUY/wcpjRXc/CCwUa48g4XAEov00xbQjxjqUvw1HCgXrKCKuwenJPyUcCMCu
qqsidjGAWHYZGym+L2aO/Xvp/EMVU71eDDErsob14xmUoHSO5Mmp6IrdG61rE++7zPB0x8vaeRAW
NkGEdsSRUFHZJnX8VF7qoP9HZiRDu3PID2UhZrlg3WiB2zucF/zxt/1zmOMpzZrF12dJEFLQvNcn
IKdqk1WBkVHoqdmSOJFW2xdKaveVQOeahwo+FyehEm9K4hzaTOMpkLNxMovhccsby4PshkExiwIt
OF/fBWpxS3EJ2lzdbSqbDrN0IYVE2VYlAnck2pjyGUam2JxeEzFTUKOpdd6lK+uqD1u9DPB8Yu8p
9v70lg0JwjaVpTiEKp+ETFYPH30ZegGS0lDyAoL1JyaiIqlJnPSyO2J8jAugr8dihHgePCnIZUcC
7bMaIv2oq3Q8vvF4S9oldgH5Kk0sjGK2Pk5hi4kfVTXxJ7GdWZ3w3o57+/xBGcOBA6pYHTVQLtXr
VGcDZg28+qO1ikeHAbt+BdEYfuuKm7XtSbf6HtX1nLEjZoNH4Uj5tTt8OWTkXbIfoN/EQcW+9mHf
SmcmG45CXbOIPni65WT7yqm1rC3Ydr/i7BI1WtDeE17lSW50EzrHRfkTPa0hZHtUGJS+IVhPzEfX
z919lpsAT8nZAQQF7ywhp9SHsDQZPJoOdVkIzDhEDciN6JzgCz5E5DKElwrLNOKzk5rpkYrKcMNA
KNkSPvbDx5zli135bilB49nio+VBWqkUQlhCwkqw4MpOSiApIo3eRQ2kB8Y6aTSaJadEigiDXzut
gJqxIBAxPpwlnXP7O4MNuCto6rtHnrWo1iJqsewMZRjsbEB/CD8S7GpOjsXqu3dnSRQZ2PS1vplh
MOHoamq6V4gPyFZcpwT55S+RghA0IjnEvzS1CtQFmBBzZzr9QDqlbL0oqma2pYbMBwIUri4c99ux
GZEwlDpWwvEothOLkCJbbrWirIDlzOst++63bKy6YSVVh7oy8dymC9I5VZuDKB7+aR1lg3GE5WO/
x0viJcZY6y0iLcj8i2ry3yDPXpLmGu8gP4ZhljsHzTcm1k23MZvDXIWFaizlytY38nVDHGI6aPsh
Q5dKZV0cg3Wyj+5gyn3QcZwSnI5oswmLyT7oAPc1m/sGaINvfU7BKQ0m3HO+w5r8zH3I6XznWqts
aGkjGA3VYTyZapOQcY2G0Wq06nR2wpSDj8W8sl/YEmZGXTZsmWLAl0ykCob5/lHfS66MmtCY/Vuw
aBpgJ5uKVK0o93S6VByuhcLlpJ0Geq+KqP9GuqK3zpAJGm9i2JtYXZWV0Xx4APOXcdUDlX3vwbd+
LkLCDA3CC7yUmPtzn1PNUMcoQ+r0exIS6fIK4MVzI5JOASUaSjqdmeJ4mEEmAQMG+5l1h6wthXn+
6ZTc/NWtNjdMBCe5utUlm8AbVM94pvniFO7SfbxSvX7TW8jOu6McvQyspYnMi+fMaID5ziXZ99OE
J08qQK9fT+kYtP/JEHNTUdww+gzvGsTSdFuqsU7IEAz+zGxZNGYARxmMduw0V76avkbygMOdOsU/
eVTfRDuvD+ERq11LfDU2cv2o6l26EM92VChLGhFWbgModt3DBtmTCUWjCGnPGFhaR1jRMQouFKf3
0RAdHLBeYYRvGdL1qiwOV9ermdEWjJY0FdDVlxLOTtqRLMw9l/L8SxVjoz/7IVsZLpv8Cd9/ZSjd
qYPJF5LlK7qxaX1yTximAfOoduRursdQCp5b9dQvQ+BrIRblUn+263FLApIll9kZbCuS/UDJDqCQ
x62k4kdDT1hy0w0clBiSrdbrzZPXdLpWDuyySKh5vbmZpL/nwtzAIvQbcrbT6B5/mzsdzTaKckQ3
bl4FO4WMzGUJ7JC+aVbYaLjVTLuE/Cr1WVcRB0qsu633cQbyetGESrsUYujfW+HZG210Cd++McxH
75SqR3mnIxaT3sA69terzp2n+OSpiKUHKrj7z35fkXlusZhyuSKAIr7mnQ8myxipgITrkLePrQ3b
JPHPU2QfT4WD058niPy/XPRtu7pOu2I8H38nz8Ef1Sa0g4HzuBt4SnMF5XFDoIPNPtEhPz3jPUix
aiETzBnueLB2rdThl1K5RtBOdvKT2/1AZjS/IuqU4bRr5/JmvrMkPTKcvLC/TRP3YHZo2hG4DkWN
I8c5hgQ5FEiccFDT6vnoMF/jocep9J0St+6nXlCIFC7fUA2kUuKfwfQR9nQeK91XbGNqQgsQpJWm
uFv+HH0+Oap1XT5a10z9kLvGV2POn015HA89LOVlG2j8+xidLTraDCQiZbFmgxQcMY6dd0yvBaD5
P8frngFRnzEExAsd40F77WY9knG8nVoP026eHZpl6TkSBKZgk1YKNtXJyZmf4bTsCY5ZCAw+vymv
zGP2wQ3NtdjWnqCMnNlvEGQ1UX3za+t2NnAM8Bmwg16O2ptj9utotEr0NZsiY9O6RvaVJCUCM/h8
+ehLC7wRoZDrdgncOXAtbA4xDTMvkd9St+A1AdxdH2YGEy28i1ECLhqH8IlJ6GmUPrptpX4d57Rt
V7RSeisC7QD56UwoEZi9u+C10MZlM9TDw2rlYanAWNCpE8pxavi7H4bWoQoVTPsC+C4cDHQNUeMJ
0NVkV8vDNP7yj+tLVcFHm9iZxBDlS1+LB16hVfnGv4ujjjAd9HOIKky5tWBWTXqcUUGHg0T4xIKT
KsCyOKVRP9xlPoSdthKTsD9lXjf1gQKGgJu1r6ydB+/ZePJwB4crgK73/lm7jPisGdrWUyJ6+0pA
nneOwieqP7M42HeOTELBr6bEx2433BdY3QgtBxMPlzBKFu+poww5RvJsZ6F8UhyaUrBquKAmp4AB
98tNi0B+T9bpXZu+6TAXhNGPy1jf0bXBvIJ4L9PdBDpans3AV9LXQGwDB2P7f0Qc5SEHh+QKU9Aq
YGICm4PsLrmAiZY0f8NqcNoSAfuCa98WLKSQvVtXP3lCFnr4X/InD9HjwAMOojJKbWsc6kfCYXy1
3n6oe3xyrTJucxQ6yjGeFlWpcUTJTolNV/buRzX8zeVzbImjKd4el/4zQI/gKeH6CAtwMxoYxP9b
33ADt0SnJQ5CIMbz7j/UmFhLZCgeK5Q83CyEy6QhqKsjnWIY7oXv6mT3nOvT3UAf+ERGtrfEDpzP
E5qgzeVqZcUEQle+wqQwnnB8bjVRpO2EAHrqaClwv91NW8l04sWzeYJqhDnEOSivQ6O675aGLJiQ
NzXoVtEDshsjI4V0Zcmf4vbhRE7PmUcy3OimNs1Z4DCsMhCAsuTVLtXVkc5jlUhfeNgQtyu1ZSoQ
rZ98dvneQCBVG84qkUVcdm6C1AAc7HTVVC33ayakqKn+d46KnuBBCjYfnk0Pls93nJq8aJNipfuS
Klm8n9B5k7TGsPU9iWIhj2deNRXpLf5Vma4hOFeHToXKkFbihpwtp8AWwLzQ5z5QxRXgFc4OZ+ju
j1RJAfG2xYsovir/CBezM6zKIG0HWh50WwFAa8do0x1m5hSDBug9SdxmmsMEdbjEkKsSMFb6JGLj
/Azh4PeH+HK8P4faGkIcKPhB4qJ+n2i1n8CMlkOfI7LBB03TLvD/OE0O89uZ6GBnQ0eizDAXziGD
kxsDu+wrxKowFpYCcZLkqX33yYxO+1iJh7nWVIYLDLOKOPmEuNKuBhxfIoqlhb2Poi6zlAr7CakR
56HIQMIf5k7kQeuG8O2S8Q6NRpTLB9JFdQo5jrNz+ZzRgvjAHZGE1ujlqhvekfMpbh67dDLVb7iv
u02RF2YUs7tR12tpQu3+R5fS/aaLfM5VqQYsdmYl4Z3PsPeth1SfLKGwHTOvMX2n77dOtL7aw6Wr
mv03pOhL9ORmnMaTbAXBwYk86T0m/m+LcbmTABO9FPKOmYxerCJBL4u2Z4denRAhvyZG+UxTt6MM
DqPvCvm3ijE7LYoC/u00E4jePdOeqep8dSIIeA/UsDSGo0+wygZKgkBYMylZYTRtIa/zTuofXY5c
M4K7isSiTqw5UbEk3CmPbEfVE8i4wKNgSMB3OnxogoZeD4RIKItjq8FplG/z32N703r5dGPg6tks
cO+sA+tJGRIwil6A4sIgDSbJgGnqqEQH9uWkWI43fX1djf+USXD8Oxdb8PBjD3G1B+ngV91PWEee
/ahNv5Jlx295B3E5GDHWRphFGzJff9NFHeQmueRyVtSuE6mTryELvtE9S1As8rtCD5d+OOQtBdZd
/RPMul0HpIPgaNNqpbDjSELxXuYHof5J6GAouJVSgOz0BNriQ7Wnz4KO2exrmh168KfQVAaTFgZ7
u3wXEI9+Iwj+dusqBGbN2okARcwTQE96T2rwaiu10pg1oklllSLl8x4+ZcIHrFwdzDlnB3Z/3wKB
a6xp2GQDXc+BM8hWGkG0XfobAg3GJmkiQzoQ8nFNPYzf0wswYwqu4G0yYQU/jewR3dfl2bGKTPY5
CED1kD0uWQVVVnlgjF5V9zOjsJvFEc/Bomr3H0vur7Yoyz/CW1JPuNK7OJmeyYNWRCRvdrofg1kl
zPbrdsm4RfoM0di+smfr/y20S6NRCNeRtnQ/gY4MMEf8nYK6N0mn9talbUeNDJZXKVlkOu1uLoyd
oPGCo3lMqCRwiNrEIi13bt3bxoYzmMOxDDz/8siWeC0vBb6hMgF7RCSKrob0Kgad1SPiYqlmH9Bl
GTgwHTekA+yMrrFAL5OfzXtzhfqEgiDrxeUBuQHEP01JkgbebdI1vkp66Mj4HjLdN6RuVUffP+k2
vZbWbcUG+icbzxQfpgMdlIo7fjXGgxxeZz2qG9dBr5VlLeVwtoGjpouZuTVzc3cJ0qskR1dTP8PF
aHTpj9anQgNK+I37hWBXnG/G3R+jXN6lOniNSgfnDlS6i7qLCpwWvoupE19X3Km8Ks1z4G2t3cp7
AdKaLsjnPFv3bOJV2GvKTzbgMOdbFoWIC1sCOQmCq3pRFOHmu68SdSDaA4Ts1faF3nNzt7O5fcT6
j7smj31gat2up2cvss9AiruaFwC75mW6QIGhcYJKI6yU83ijvTbEVZfx74+5RXpel/5aMc94SqXq
vYC88USnb+dkDULFGQ9Tpw1YNjufJT5QWlRWrLB/0e9e8FD/RxXK2Wx3p3bEnmbe8wdk4LU2Nd0E
4Rfq1k+g3rWjueXHTWV83yOiK4wI2NP9bgMIJ4SQRRHG6cT5GXVOAGAP3HQqu2Lczwi2vYymrLDE
fSuGUMeMxwxQteFV2Zqdvrnf91bbXHAjxhOJxwg6jUtcOamgdEdYrmmE7iNOJMgBqS7R+MLuaUcS
S/lWRcl/AHMLk1htbRmjigWG8NZVytXsZQZHdIHltpcab4RGDvvdlxpGZlGO2cd6u+/BqUSL7nnj
jz3E5OPpGg615Tz89ScFWxn2tZ9fmgL2wXCPgaCxDiyJQIDMdPCNg7P5jhwdXMvCL5GhjbT8aUge
n5FTZq+DPAvvWy1x7XW5KsdM2N2gC4EPQhE1kbzCoS0BeK3TNiGryg771V3BIv74MtUj0alpxsxN
IjQ56AxQFeH+W8XoCV2ODD6ZwZKZpZ9+XSXDb82QfTi01qXAZ6weoR4ykr57DqGGwLYHVHLOpZA9
GlE0YDxhYfLCd2yrvVscuVBp85pPB5Pn0UNTHTkSOaZPB7tBMVNH7PSY+7jRenLTMPNvzEEyHPH3
EpgWUSsKBopPBUW74T1APDCI7PlicGdyBX51fi673rlGuMfFEA+y+rjHfBbEZdZHuJYdXHSBmUuY
9klTave9rRosmKWYHl9cgxJkWKHYiTnxXR0M7W7/1JkqgCHn11CH6/V8RyFAMvWtdJ8jJMrQxTzP
ETuL+j6Vxejns1S5qd+jcFM5thuRkbV+zXHMExfb4NDMUPHeOPWyvZJaojZBjKEX7SP77I2NPnRW
AmBsvurYgUYHtE8zAYCb7Wp+aj15uWxHMeCZiFGsQ5wH6RFUjjIE9w5VETVbam5cT+lEntkPx8S7
wmzwmWsy2j0UjxQ2plL7kYLvD9e5U5DWQ0TDyyZHhRQ8YyYmgfBziOgSyeq2EPfF6OhmPiXLfdQU
laUVTY8LYgf357yRznGqUBjDJqHNMJ2vHHW71WD682kIDaTlJwRQiMzuEO02mkco6TSm7LMIeyUk
rfthhgjXUW0MCoD8XeNyub/AWMKWtKXFRCQmEBJwqcsQfO4OWlfZPhNGt+DO9947TdUF9q+nqePO
Al6zJmjxMx62DOzOYQj1LgwwayG26NntFgk7lDTiLL+ZkoGaMEwCaAg/MDfGsCyYOZaf9pPIPAPs
me9z77DvXqTo+fWiIgseb09VjkTbIJGge1+PfWL1k/REofgneAjFXh97Jcfa0iT0FKoyRiOOjVIs
FzQhFLE4inHVB2HLVuvtD7pEhiNIyLeEF/nVJSxtuWZC9SBL32wnbXg2bQfDWIFDmalVs9RGPXnT
1YD5d189/b91AFbG0uwMxqLsh/pfX4xuGuvDqernSjM12zT3RwahEHAlxN1mgjSJijGKwSSPtqe2
OE1pQN5LDAUXFQ1gisInF2zV/sAZVaBnMMgrORRc/Lxfhml4oASgQjvXUR0XwpQvIpPXyYwUD+g+
zsZjJ2NtxkyAPHlTx5YhLs4YY8UnLH5buyWT+dR6ytlMwC5irpnLDQYFZ64psVtWswkVGZmbuRaa
PEy5Z/xO5ynpc6R9xthaeFjbvYJ1dAiE1AzjOiP2kprB+ppZ6jLpdYD++BFzpT7ik1eGnwPLWP8M
NOy8ikAMoJNPCsMjvmSa0WImAqQQhuMRhRKIo8sWFZBYjHrs8uLq1UsCdch/NHJ+G7w2vEMaltfE
2DHE4SRKNao/wvC4C5UypPBN3HsIv8+1mz5IZYl5X3wFgqWO4zdqIDcwT9jp3uHpkg/3EZEcpB+p
A4oJmdi506F1FTNqn87SQGDkGQNMZ3Pd+j6dBwDBmYj7XYuGWwLGtySbKQ2j1lkxIRf0eJSj/UF2
ukMx8Ro369ufGkVnXfu3sHYizvQjoAxyjx98+/8inwsKAgxzM6b/Y2rf4a4wJktskxy0hyg2PsFb
1GUhDHQtPFw7H3sCKpS+Z4RXCwbxNvwtUkE9+XqKayPIrb7b0KA3K0+auqLeuXoARKP0huTpKJfu
o3ZRYeUYogCg8j1gUtuY015ha7v/qfJjCkt+9eNlRlalYNPniJ7SDt4DwTC5CrUE/S/2WwZE8yTY
wMLHdAAYVwgCyH0uu0VTor65tXawuCTLlshFq5wuAhlGu7FTIAVzkMYmopz8Yinz4hg0FnMp9ck0
kN+K6exRxV/XRIB6jHxtJK1w4cQ99ZaOJ7NF7zBaClmcYzKMm/pcHD4Dkht86c72ZNxfJJEDLpg7
n+15nFOiaWlcCFtWwGISwNySR+fVEj6y2Exl5nUtkm6D7NQW88WPtei19rKXh8mrmL200Y1BcMAU
Rs4MxTlAzCBhhFgfHRRUM8pG90b+KpUu8rdwRmDjbH5Xd0y4q1eSn/tPnkT/kJHyB/9n7r/hasrM
5q5TNYVjoHSbKgu1wBsUCOpAVgZZiN5MOg72I+Zdch/FXS9a55yF7JzqX+8hBulZjKdptpD9DrMm
kpZrYfeZsHEiM9pTOQGQ6Pu7eWfPszPPXfqM1eAYnT8f54eBOIzvp5WHps9eKj3+lWmqyMioI26h
ZZa1P95F89UugmtLCcMmgvFAF711SeMRTo5royrkQJsE9XlOcha8KURqP4iOnJUi6O4Ub+pZq7XE
HNGeL7UiiqwAcTrRlSKAj0W6UTzoYsNzxVVedpQL+SMMUPeWOwJO9I1J0XDNq9AvCTrX7N0gsoSA
aBoyPO3wjLCIgDfAcixdBNZ13aLNqLM5XQNcaB4IJR8LTCavoRyW6NjEykVnMWKSCFjZ2m3VwiVZ
bNYFXzaHmhFdU0fn/vBVBuuo52GE0pcv9q7P1xOjCjSIkKXZrisftrQoH+7D6AvZxHEV+0Gjj+r2
UfaOd78NIDyTFck1nKHBt8f78R97Mkm88WWu/QepaieWYO0tnX5BVY164FleAYkMLIbIFeL8MsEe
hoGT/XgwKqTZj0Lt1znWcQ7BNqJeJ+Oh4KiGFFlBYSEGHOCQOGB98K0+czVhP10M0VWFVUSKJCYF
vOJ7E4raVnt5pAr7z+KqkxXbk6ARLn7UCopCNJhWfuYN0HgdSPwrFNFl/8skP6h9CYm0frFRDnm7
ThPFPMR275cCU5jJUk27V7hfdVNbGoCs+Q/tA3d7otoYpFNO1ugIdjvgDMt8AG00nm7t5N52NiwM
ihKC5ixNOXq7iUGi1tWQ3w2oXOBDYpssuQvX9tUh3tO7YRNVg87/c6SaPmbO/musy2RnqTbALam9
3l/aKd09B3PnbksXDJQQyL34BqxAFtFeh3fibMg1oONfz+pU993MGz34fWvdRg7aCDXH72oDRYUL
nd+mVdVmduWSZKjCdPX0D11GG4cwx8uFWChGkIgRfyDGNbK59pxcisi+Nfnu/LSx3PKa0n5GB797
EEZjIF8J0xoG+P2Ip/FXEv/z/+fNAEcTIsAg9WlBhHMh98mZbHVIA78u7m/ZKWHIQnElQXqCfKKJ
v1y9ulazH8r/GoDgL0Y7Ov/Q+o1gqfzXtzNjnMzMv/xcAPheaD1NBwGFIODHL5LTKPYUKm2pLfxP
lXbeJGyv4sk23myauHvLA18AFqukI/axRAkNInCJJLF0RZozdfkFzM8FGPnoywptTgYWOvTUu/Gs
9Ul+3hvcLhIW5jUhMyZJ334jS8Sfj7dQ4GK6jQLOxBDV8oZRP3kL9aGGYE1axpQR4+o741R/7/rY
qZqB7qxG+m+TY/mfNuMymiIP1VN02GZxFz6vp3D+RLgHxHOh0HSO9MyNC6Pca/VPtfZlvoxPdHhd
f5SUCgLXKKbFzDMX3aclbuHyfTjJ530JHtq3290l2UzqAxfgwsESpFMYsjnih1ZKdM9WHqwgYBpH
L8ZCY9FfHMjutd8TWTz3EUGs3rKe2MELDGON5NJtfnJxUT7VowKcBrOt9WF9W2+j64fUCW25vKUh
LqlzvBqzD9PODkceQpmVnZQZ2yM40zakHk0XBv4o1VlGv9fjChIm/Nvv7HTsX0UzXaK4A0nX5x/J
TrpJKf2tmvoNEsONT2dmPX72A4JwVcvWocLktjXMh5qOzrD4T8Z+HQ39x9BjHdeJPtpFwVhCxZdF
ROo1nsL4Y7vZk4K36ZgTg0d7qsxS+uYosdSV9Bs9kebQcRIoooLnM/EtvcD4D21ONapyinAu7W1L
ig/qS069oGzwlymm5RhEi8r8hmXx0OpqwU03NvMBkUVoVH5ZJ0lsWzJRkyTY43lupN9MBYLamEF2
YxS7ojI1ybhDLXvNq9kKegv2fKQfuedzE7FN8xeUvNhR72FQx+k6UlNhQFg5yNmgemkPvTsSLkf3
EyKDybOAH3aHvMNa8G8CiRzw5s8oZQff6+bdSgPKWMdEtNNUx/Mnzd4NvY7F0lV9NHqxps/Ibxal
fZTwDEsojpmw0Cbj/vFc/kVEDSIhOrFAp9U9KkOxERCiE11OYWMD0Xqu2HNq5FUiZx97xZ0ISmHc
zl5GfPx/QUIHzIBeZDr3sPXBIaIJaC4c0A4XL+chVksarI71M7A/q16xurls+0tXQVmIHy0q2HSa
Ui8aaUbAd4BfpgWdYObpaAf4/oCXWv0MZ4y/YjjDJpZURgdKtsePPscdzISQLgGX/NwOR66bmOJr
lVR3wY9rGPtLaHrj7hYXm/sDXJma/rd5BhGkJ1n7pbgzXhBZW/UElXAXw5VFqL7bgXvvVt1Ws/sO
za1zxYOlG+QkZlIKSZv8upw3XT6KIXVX9F/3Ag7EMFgJHhx3qxZZxaECwmAAO+8Uo24hCthNquHB
czW8txTawHCSgtxwRhlK7Yu3JKZAz4F/+qkhhKTQCdQ9YET0tb79Y24CdAnlGQMQaSYk7HINvxCX
qvK1X/3m5Rt2ZKyW1Quj22H6ka+BV0HleHr+LensVNOdVCYyI52+kZMnI8MVPEVkVV2tr5Vq2Nl1
dyweJRwYXWAFRn414cPtauC4sjy2Lf8XT0gQMxt4IX4vW5MNYQVWu7gA7xihoPLULNfuxib088Fp
9HffUmVh7ari7R91d30kK1H3qhaaKaMxXWVrdf/emFiBz4l7d5GIfEbQ1b1bR7HPciN+cguQG504
7a6RORzAsUUB6Y7rNh12x3KuZ4cqaWdC1BKJnamvtb4rFWdZItuSBk5NnFRkYNnZ13AaUSFH4Cye
2V4h0DRrQzyW2A9a9IFzJQqcN0qsRFyFJXjFv4UIg24uelcBBs52rFhi3kR1XS6j++fY7Hh1b2/9
vdUn1cRhBZjgiuuLig17O9u9gckMwXOYf1tIY0HiGqNfz0pFb3aDctxmJhCiY2CPTcqMFBKZ51aB
Ho+dXgc3BEVIFeR62OrWn3SCGcGwlLerPJ4UgrhxxrcaOs0xYwQnn4+o8nKd89zknuiSfl7UGqrV
0VdgPlMaRRfnNHp1jUwe71G4JLUSzyMCSAoKGqWx8FjRRC0SqwQGJ09PRxV5Gng9HCltbUgUwzBf
Ds2+/gvQ1ifBLOB6uahBBW1N+3bMHzX3Zf7Cvf0it3FlrlTvlayujmpI9aCG1vM/KfU+v3pVj5Nh
zaJwQTk+qrjrb/9bwFW5CH3jzalP2wXLOvFj1Nc91YUBX58y1uYgk3OijR2lpSqI4pz8lpI6dR7W
9Iuhpg4f1tKR49Lbnqr/sbdFbG+3wlhURm1n4mxCuqlhbwhB/BA9CaYrltxhnhuvcnLla0YbJHrq
a3j1mt3FW0cSKVB/HgAA1nBN8baBNn5DdC7ewQdXb0ZoOl2jb/9tfosqfPHmIwRjSRqd7RvaAfjd
wZAdUkc/LG6sLIWNpZTOuiPPTM0DNlmk2/UYSZKPd4MJLBZfRbo3ErHyPQLcAedb7LSeK1+qffyd
8V+BQ5t4bQK5xnGVbsMQ38FOjLjdAVM55w6q6cPxW94D1fwyf6dyBuTIDR/475t3eSzoafZq6gfB
S6vLdw0T+jLe/i2LDa0Kg0Ik2JTftal5T+hx9SnUq0PondDZS1Ht4PfSMxXlsqgh5fW0OvLjhuCj
jCUAYD5PtqtycDxl/19khZ+EIhaPh0rYVL8OEOD+9h0Bx3AYan2TrcTX0iHu8W73KtkJsdHEAnuf
6MC7tDl/nMgbMk/63KRKRe6EfmLu/AM9Je4HDGopvd+JFh/M147HaNoxOYpfOLNBEtAh0sm+HvFO
hquQhKIn4mj5bRCZEglBcY4BiAYOAkmGlL0GTNeL6y2/B3BqIL/BF0bvci750czL2T1KBYIdb2AG
82lHeU+VU6kv+Llr26C5yAZ1riTVRoaFFUHWK8RqRAtfXijDMooF5VjDHhLLEvTMBbXYf//DZsvs
cfQOv71VWWBuynxiABmW77oaD7l2RtTOTJBPH/fYqU2BuEbPWexdmhRa29H89FMeSldmHjiQuA2u
LqTpq29uxoKgxTNDRopTruWpzCnFQ2usMOc2trDrFM7wdzcRk8LVLljkNsP7dha37DkinfP08yzZ
5m8nAXuhEpYynZDXDD1uj1EuOc8ayYipZPnha2HphFfU+k+1quV13DPpaeGH6yD2T8jgFNa+7S60
2AgoBaSUEwun1xzm1QxiBHfub8ldro6t3wVJ3IkJImtWvZifcBc48N5H5Aj7udoEt/EHQbXN2JFw
wFkAosAkrKFGJsLGgvGce1vxGOYTn/CxETVSEDCFWI/2JoryUw80sToK8ckgJRrH6ORhC0qHSE2f
Smdqdw06HLAijIPR4Ig6Kt6F1pwr0CUmKxGYWdNxMspA5AfWFME07m0yQyT1ENsOi9IwhVxdEslp
MqkBjUn1GatelRmElaOC5xH8zNTC+cdH5vWZOLZw+GQXJ6t7SIt8ef5orRJtlpQ9HK6z5/1B3UPC
rEo04mjRa18HyjkhSZUMDzyN0VubXg49w89v/ejhihI2sRIyt/UU49qZbvm8EtSSFEyq4JYevLXu
SVPbvjeovLlV3Hj3lSuWUfd/GzxKG8QgLkqFXBm55aWIm3TTJvjXkO6vo/XYqkxNaN41iSy4YFjJ
rT6+7FdcUuFRILa3Jb+R0iv6rW1y0GjY3kxlOkpSvUtvHdP7cfilsKVQz0f0Kt0v4aQnM9HZdsc8
PfumU0Dyqcshha5C/dZcojVF7qzVZROPD4T2M4egwEuuKYB5zWW8k0iqyEwgvvF6aF2Wpz4/4mkJ
+tU6QMBc3lG0QxPBjDRaTJ8x5wVASHDW8D7yzeBTwoTA7zv681887j5Q0v0DXH2ITGxlHSStjYgS
9HZpNmMdgci2p8loFRkYXiUfrz8N5feLJuceJQiBlVx8ipv7z1tntGOAeCA5ax55a8sORX+286RR
9cPAkxzUt++BhTAdIe3kyYevju3vx9JNFy6djSP09hSuMstWN6R2qfEmhv5NRc6Jdd6cqdB8AIvC
L9t2NRjcMeKN6+m6K0X7P3N605RQzkGFBmD03Knj/YLqSsfSarPyuVOnIeJnMP5se95MnIM6n9qB
c88jEWDXj9aF5Vz8+iw0pAGoQxqvrkc/q2VK995khJ3jzTyTyXwQgRLXdjYOyzvRqFWr4zsDFrpL
qitsLxd4VS+IovI8YG3X7lfqRdrVFsp9QA0Ufa3i0Rjj4wtIcwORpvNq+UKyb6fR/a7SWNS1WFj/
qUqfmrpLZBif4juXdJpAJMUBukzQlqdGpH9sWve1frNNWXYgoL04Cl9A638Sb+ytJpWrtd3czcdY
QjrIghyOEqp0Iz62KM5mq4wraUvMGfXpHWh2hYKU9YmagqlIA3y4WlTN9kCAWqXr6NTYUCJ1mK3e
d/1+gK8G2MdZP9KN70RzLgK37Dsm2Xiz79da/lmj4b01Kdb3JU2m7Re4AcNd5ZHH0Qij13/MIUph
kg1IkUelDNKqHufwgRgMQ3yPGjtrruXvJI3SANSxINc5Y2kV+HKA16tZDH3VtN7GU1Q9rvNXx7A1
1L1LNv70rni1IQWL3GarnNuxVMEesBfrAqO1s12Oqmor8KdQCtyvRimoKMcOy5o/tDZBoDOW0iDY
RQ+cRuJJiSUjJv3EOT5VI7WNt89xDQO4p8K3Zx2ALWbq4UdtixZot9EQLQQ5x+pXfqYlC6naJahF
BkC7zPCC3bGfN6WNaLFUQP5gOjgAFGws+nFl9JNNB1TTNqDOLPRL1BnyD8h9/0Y+Kx2iQOLUHFjD
HLa6IvgLsvawc9XswhKn8LFXyb7Udrsk/w1hRpUXjLSgJhPBIgOz97pcjbO0LIyvgGO+/4t6rDip
QZVh9hfBgF8Jw2VHMIaxVgUnDXiTwyLPhiN3Jfj3X5nIlHeq0z8hpTe/dOHlLGhAoZ4/S6HzB4vi
onlDq8UlsE/4yGd37msocBupXNVZrcWXiRlfbwKgImdRJoUTy41i+PB2MZAAw67LeOkmgiSxmpa0
x3gQQJEU2WiVUtFZj44Bu5lB5fVw1piRlBKM9ALuhRbwWLIN99Lm5Bb4mo+19boliFQ59xqF0CLM
Nx7nlXXt4TP01XHAA7Q6ZpZkRA8zbLP/YB79/mIMU7xGyB/5PljTn+pbMGv3LNSvHno7tU5Ojr5E
c0EtwgMTpZApANL4Pl/1CF4dr0O+hSiiQWMZ3Z0m8vX2TzZu3rV3XmKrGryjVddjsyAzmRbz8OpN
/Hy3TCCGkXTssl/q74aJWZHJEIwTtvT7UjgMWfPkXmx3t8sXXReLiXzdT8NLxWgRwL4xWmP8Dx16
YaV3dlDSrgPdM0/UMXl9/Ug21eT4NpEOhAubb1YD6MQRvsO+mg1mPMDY/guGD6BZdeg2oUG/d7D3
wrO2w0CXQu3BBXFyVjpuR4iXev+K3dgb6GfEjmxsH04tzLHVfGLPU0USWDTab02ylpXV1Gj1hu3t
fYqkT1Jr6gVAzX3yBEYMWwGUncUqkPzCWOvvsiUUlWjfU5QUbKNxiUpx0pbzqEf4dclrHWrj6itd
teGBQucLbAbkd5nCEk5XIu3NXNWygB/4SUlVOz+kZ0VZ1NZKJygQSyFGM/347hptfPpps66L6oTf
MecDI0VuNuUr3twjrSns76cnixceHLK4CcI+sO+sTUs36aQxYN1bfcpLxwCgGGTq7G3YvAwPRtnl
8DVKIVAElD+rQKCJGEAEVm47r9nBU8GhKgMV1dNO8nzz0ajvNlP2+mJMV0SpZd/biQ82vucIwyPz
NV5UBtHZZlfUbfsHrtx5w5Rn3CflGyZ8AQOjsEc8UP8qADLTQ3VBhOXrs23sIGRmNDpqaJePCa5U
TevVscvfIRJrk9Y6bQhHaL+dvATW1x38hY17cPefbwTom2p9V5FRwgOYuqO8niPve+DzM9kEgVig
mbLr5vipCAiJwrAlGFJih43Vea7mJotOBRiMsRzFHJkkghstUjtqjyuXErKV0GlR0UFZrBaLF+5K
hJ8gVML/ME9iMJN4lQG0fIz5KrlGZe5sKFmzDKg421gKCUjBrPB3bt8PZTSgbwAMBQz4dOK5Mmyq
abUIHvbaEJThb5zRCvAaRNNzrEyB4VSY92w3iLuhb380zxzMN51FVNrMRlhom2TItNA7FzdpAsaJ
t9ZDkfo4ZJU2vX8jhbY3mcT8GYBE2UfbK2+n/gYfpZAZSeEhzm9rkeVvN5l5iqIlz6s20eNqNC60
Z0l7/OHxZjFKt1CDXaOXbqPccpIabY4K3a1aVGwzOhhp4a5nRaiSK67FfSsDZrGWzKrVxtIJRRlZ
+Kgkwgwfk854/Qp7HCHytxkXLpjBiNS9rVjNZmxzODuAYzEGC4GjfcE35853lTQc+d5ZdZYVuWQN
kMkgDTyzo7m0q/oXld7Aw8uqgSMeavJTob6j14WxfOFc6VO8MjcLF9Vv/ECnZ6oEjq9vLZbp9i3U
VLSZWT3amla2nU/8JT9aGpUztqvw8XqrLrDZO8vffQJrqMNc9H0QufsqdgAc+PefqD63kosRqIWx
Exq9jsZ26aIxZuu6gM9lbliXnxJwA1FPNJPVY9PywfVmkbfRNl57m6ulKJfwpUKZ8hRL+u0NdvWq
WWuHYoeQlyCv2LV/wLfzxx5aKRmYRgrpwtdsD58aOwqUqV+oIqDTqAe3Au3uA6K22135JGzL80N+
1uV4Jjy5Y6bQsa07jzkgF6a+JgmUe4zN5n53wdwPF7I8JY/JA18k7c1mmL0M3v3FVewapou7Ubfe
n85z5gSp7OkowBrS7ownUECR1BZfPp77Fq00HSdgNttEJOXGoD8Zi8eAb7JCTAYikvDGaPkLGLDN
9ax1jm1UMBd9Bpj1Da8Gk3tJxI5aMZFDvtE9igcXMtQ8VQ5OZ9mzpYYiaF4oVreG6Nd23KWDUuDa
Gbzj/zzKz7nZrE6QfskeG7KnOZUcuXkhvoKaZwI3gOpjm3/pHFyWl57uSs64t5CVPjje0RmwKK3u
Ojfwz3BVK3o7VwKaeLntAyd2EOg8M3i2CrMqaJQ1dny0p6tl5eG3JTA6KoGgn4d35dhl9zLSbaPD
PjOxiG7ni33hlFEqbRGLD8F1Hy8dZvkpk0rqMftXIMhKgSwg6m6lCb6eFmPy47mm2RnobLSsUKhV
k/eE9kNlydEr0OtdMvwuxdUuo0QxqS6o8uqUPukIKwwaRvV8UeWMy+zytfAkRbsqH/l54ZTXPdWJ
nmW9rSaUCcerQFqc9hDHhsPLLffpeE3Vu6CKuCGwZJb/dna1AL/k+8euogd5ZFN5tAz4oQV6Mo2d
cnfwlranAP8UK+FnIQ0ZIYs74VrwpkIVXw4e31xJjOYFNf/dWyN+LXXWj35IynZtsUl0Ybcy/4xU
si2hotgycOBfMbBBqNhTChjAtc/PL5mI3j3Um9ybY89WsaF9gPlEwI9X1z2VVQw7u8yvJW2HgauG
+tbZ9Zr5l3aQtFBLAMsJB4DtmHo6YPporUBjqf7Plt3t904UDvNZKA2It7Rdkw9CoLof51gzsS6r
3LnrFxFs7GUTObrBnqODZm+BbNbYMiHbW2nTXF3LEq1In4bswg9yqpvFSrhl7NoZvbuDmPWRTl3h
davFXGfWH+dtOIurU0IhhZXkacV/OtHxvtTwdV92qX8j88YzJJyef9O0+OKtbWf7hwuF/DncqhHK
eeCMBtsiap1/WrDiecD2QBg6AIb8oavTlAndApueuNdJ+CMHf4Tfr1+5bGCcIZMPE6MF+kOi6ql4
Uzh0+AuIFJUsXk079IO2I7KsGyjJq6AigLPEeX56D2SBnrHrRQNzYD/xarucoh+rhb7u9kCHghRd
ZWuEqWu/uAbUDezI1H7mHGKA/ZisPR0qQzHjkFj1fzEFSaGxoGpHrbjMd7sCskLZa36MDNBagvtm
/1y7rLrcZX2GWWNPW7PsfE2N3FOvGQuVGi5qI+3KWtVLqsxDEp7A5v0mmbmQ9/KlnOya701md71Z
WEvZMIKyVIQHOhlr+Q/fF5yUCtAu4gZZHo0R4Lsxm/R5zAFFwGyd3k4q7BTrlrq/dOXIyvr5T015
c4WFVynPrW3HinhwrwHMimFx7LpBUEDoDvxRcPhEKsP2vGK1Dpcw8xmArHtuggpTeItJxgicHbaM
JDJiL0yc4e8Lwmm8WbN/JJMUz038ENPzAbgxU3Wulo7jJ26bGPhBtVqfZNMiS8vhnghHuAu969jT
+axiPGvHTliqlLf9ANmuv0xy0667AccY7NXfrYQA+sb/94FqN1rsCu8SvG1AYjqKukZRPy91eHZO
u86flNY0fw2SxHUpqZNSSMOG+ZGpcizJU2RUxoZURRWZNLVXBkJMjDJWmPrV4mfBfb60jUs9kB9a
AEvc3DtvIrlZHxE/m1AO5Uo03b0QybH8avzntPwtxUYi+IWy7NI72Du71A3Emb3276WMyi5v4ZPW
4l7oG2bwHTJlCqNlMeDdm9Ir5bXRvrVQtOIUNNjmqlfwHWzeBP3Z6XxSBkOZMvfbOADQQPY8NFZi
R/oOMKXujocWtEzeuOmtBVcdew/fsSM/QaoTcV2xYzQZdv6l5YehWKITeNy7PzaZAwURTGKdHJOL
SWrUox5EY6WCWFmHg3KtMfx7IPkBYxk9yNjM/YJc5AYPLInGWhxZzeGsWH6KdK4UoBGKjyW2ZZsn
ux/xC25nV4I8ZHlgeS5XYNJi4ZD7K/KzIxlwAtF5bjN6dhuLpOo4KU5/OpgRaZWfAeoglQ60wGWr
NeDzy/yM68XNZUReScsS4W/6MBvXeQ8XZ5eXt4jAlHtes9gR7NRStRs5vGFWXkj9SZmoJpPAurfs
QWCXs/TghXC5Fxy8dFkOdKQaeL9llmTXGWpa76E2BAG38VQPRAy4W5EbvU89mX4bQuszjvrfko8S
dbaEBDJw4XU/Ej1C30MnNhQok5OS5nVJjfXqA0HeYsv1FlRi/Glrmw/n/IY+lr8d5bH+P2Gg8LHt
vSgo1B9ey4pD9K20t8+H6Gb1MsYahAHKAN1o13dkvrlXLQssZMCVYdbD2p7A1XwE/U0E5pTb7UYg
LjeMBBqGXjTP8G7ELxrhmFRYeYEfwWZaePcZQo2fNOMLKfndH4Y7NC1iC5wTIayULX9JMIXm8p0v
pdogsQJuR+W/L5av0K5jAWg0XGQD24hAzqv9IqM9RfQXTPyMUwuxEr48NFjcK+qCGMcVUHm/dC3I
mQNfGR2G3CUccTK4WZiu/9Dv6gTihNuPBEoEsPQ2N/6xYGh496ZNWfDP5Rm3wF5ssWrNAIfFwMxp
6BdEsmzaDCD70KB9gyQCK/R8tx+2CgczhvR2bxHzPPUgQHm0rM5E4IdTtcNoKxcyMHusWzpUI9QA
o5Q/joyGD+kZ74KjxEJcKDvJUrd+KT6oz1t22eLxLQJYIdcDUZLIF+FDMQ8JGaVRwKVdt2PUZ6l7
Qd2MNrKHHsxis00Oe3nbrrjo45xa+RJPPP57suAST+dXEfX4ZwXiCd+I9EqxICJLJ8jS2sj/v3ML
iuxes6udtH85ZsMDEJhEzo+Z8lSuK2mEOFDRIOSr8MVpKXRI39xTnjKfnT1xOuAycj9PPDQU6rBE
Hra3b5exUpK0wxOe2zC5PyTYQI1/IER56s+refAJuSlPJYj9jUSMrMjeO4CXWGk1TdH5So242zAG
w7jzvB8NkMKimT0LuUrCiNFKoNfbRC4iUCkmYMPHWnqZVJM4+FxagaAmVyray4b9+wRQrXBDRe3E
AhgtOST7ed85dkmgERHz2eCRZZARA7KLRxLhmYMmhS7AHUBQxZnQqE+zdjONCDdcTBm+oEAldfxX
9nTDmvwz3+qoUp7dstcpFj4+92QjnKub7sBoMwAoy1Sy6LHMWPpaoDErz6H5X1mU0YrqFyAipSmW
l1YZGmRSK1aEBRFi91gBOmiEm1yQe3Ed1iIipDkXbaWavBFOUjVvEr+x0E7UL+Bp1qmW0D1WTE0H
puqC78pHq3BxVBNF83o+4sJBu8rOPPRjRs2Nvk0LghFrZttIJZzUpSc3lyxFX43a2azubsgCw+87
3yDFKdDgRNs4WXq9n1dG2ykmqSb5ZR2yMlwiiGXKQNVlRx5bruagtKi5R5vXy9BwKxU98RpEtekt
eyFnxH3BE8jofNsGm6awtrEgZJr3fllDJWhVXe4Ov3TuCVkiwuiZBjyZ/WMg26KZPZrEL3Ig/bFQ
LcN2BgpR/pHCpyULpVABLrATWEGIrl6HumyNabycAlPzzXaISfUw0sA5eBf2Ot8se/qI3YndxMdo
kPuXf28/iRcLXDMatferqd2vUkrSj4f8eBm/bVAw3aOTXUNCNp8Pl6ocbQFWeFAwCWsNKmWQHyzI
EwRXpEseus/s/DuzZUj6UoOjEk+H3/5QJgGOA005qUmerNRlJGSOq8N6qMml2zh9ujRxSy8kxq+k
AfMx+zoo75gty28hcih/VCYyyLGWYb0qtZEq/Mizx1YJrjsjhthqJvQbrqqmPtwL+8csIdX/gAWv
vXBE11hM2PyAc14MhcU7kHo0ch6+w/48PlI+b3nTSDySxHM5kzNEZTyL5FCwpbbsPN/O7GnXSfOu
nI3VSizu1WpJKBZJxk2a5uU5UfmYaVHZHe0NkI+u4O7QfVatpmWpZjfvdCfkSghUIbMExQgXe5AP
YFUZ7fC7uMe7ePvFndLlf0JXoYfWGX/KM4fxVGq3diZKg778otJBjBX6H1CCWWpUSnEKbg92totJ
4fEw7gG9LW+ZI+xW6KYC9mq2K4s7sLrv3WnTCQ31SRqgkgftrOO5lH9TbpmJvCkKsHEI7SDNlE+l
BAP0x5EIH2b3RcaUu9Ti6mOxuKAFrWwQ12MzXjSv5DSCIyK1bl9lsqzcF+KGcPPXnBxL1QD252JP
GCbPAySnX9HLh7N8wzjrOQMDXQ1Gu8MS/KInuC1k3QMhMIsvD2vpbKJXcMIOflSv+5GKnw58G0UM
BfKad/FKUi5Ql6AJWvHL8vnt+H5IMPZmaUekuYVbiF85D54FdKpSTGX8YU6fiZ7JcrBlBkC2ttED
vrsgHtn1gsw6SN8UOJsZhoKiHYzuQL9A/pdSHFQQszXOlKEQsj/Wu3Sm4EzYUHZrZHmR4VKIXM3p
ADCqvlELaxAqckdY5oJ/CCEvM8Jl3qyciPh2AFGquer3XrEsWT9llEhhIcHwZ4DGklHOvmBbEJ/9
7OL54xIHlAxg4JcaebUJnqtPS/W28AeNCd721u2uGyCBdBvN0uUFNEe7G15Qy8KGtgbW86S91zoP
rVKilrljYZbYLtV4c2DaHg9BVj/ymUQSKmi3Z6l6fyqEn5xYteS6vLSTmdAC/dtd5IJYjrWCuKqz
9IPgzr2e8Jmxr6XLKTtjArJ4iY0PvyAyM5TPK6zjZXv2Oh54qLHcJL5JJpkDifEDlikiWcji98ie
UmIrFdo6J3cx+2/KyMT13zF1YR1TZ3U+GECbZLV7j6o+DQ+gg/8ffdHRXMWMTMZ1vCRdd2jKUz0I
p2cmkHxpNgJU0KtnYTk4B1o758UuEw9bCxy3Ua4BbSSJT5oY+WQ+r2Z+lfB6/Mwb+D/Lno5iMfrG
Ii8KPvfaqAXIOJeB0ErLgQdc7kWhbDWhrCslmKO30CT6Oe0Us9DNQ2QhPVoUg+iZQKOMAEQoBEun
3j4hL2R5aV0Bhvsfm05qoTUFTntfd7Vd4aChW/06G35q7uuZGabcZXxBkuXwYgX3ZCpbaZuCdTNx
+skdhxqCrs/CVw7Bv4gz3FpeIZh6vCvccNQIcOpodhHkRMJFbfp14vMG/sCYGjYLzhV+Dlw9GmnD
DIZ8AK1ftzXKYshktEoBUZg/SAxJqJp39dgBzVLczLJCkBQmkgObTixvV+jBjk1FlwUOiTEVH3FX
ruTKjWNWZSnVWB3VkBBuqw29y5Qq5NENOBK7Nvp8TJaOq4/Y5Adzu86FHwUIcmEy4J3qRgKP0QXZ
X9MRtPDWMH9JDtDJchGAvt5Zfhf7issF3JcGiBtQq6UA28EJP8R6M1/ws6lygWf0xHKrKunw2ufM
aO8+fh3Xk1upkzA3/AfUOaR9yzoB5D6IgFdEivyvXzOopet3dHiATul4uKPyZkXClDI2m7E69NGv
rn18b51jXnmio5CMNctWNrlkNl++QbcPGqw2HCyF3ZkySEPc4/VC7cuKH5nynxQdduVit2f6Xg6n
2s5s+Wf1vS1rt+c/lrTlDXVrv9nBqqy9m6HIFDEkCXky+G/Dq2UQAIhEwW1iKTfepGrqDfjm3BiX
nFjSsSCH0xwTnOK66SPpEHo7FDontVV2EHXZBJtz2QFOwoQ27OU8ue2hr/W9Nsy4E9D5r+lf/I6K
CDS9l7jEUQ+xcRfiixUVJTs/3glg9/uQ/sweAKBlLAMSxQg+ehEfPDSzxv4puXcBKSyz9tEV7BOA
IOakn4CjX4NWw2njrPKy/jL8heCqDfFIyspQxL6dxv05/DR6Mv4RWVz2j9AESnB6asdEGb+KZUCv
X47rbODqxfJ1G61pXhWFLJACEbUNmSMzrd4eScEd8PGXEjUZzrFm/P0x2wdAYMDkTWBlUKmSd6xb
rpjaLF0cJlyU4Km5eQ8avcFXZi+C6k/F3kCpcz7tUyv9otzFQbCFAcaKIl2JHGG70l+ofYcQtne7
5wPOvwpzj37Zupaz94uZHTeJw9uK6HCe82qxFybhanQU7k9WdeR4x3VaKvPVjoj6LvDbuxb5kMNP
mn4BU65KkrK9M/h6Xe1VxvZqK0fJPI0h7aSzDmx3l3D3yQZDHD0NwkwZ8pfn9EDZ20QgjgNLxInJ
HoJ4lBnu8aQ55B3MrocVZkjRfDFDzxKUOm11GOGaaKgpVA1CVZrlp3f/zq14phQKpebyEHDNcZ9x
hBwvj/QA1O0v03VywfE7JKo2Dhj9BGhGqWL4zQPVIIz6gF5Aa8KsQPOrWANXmvgAIQRlPfn+jkT0
IeqOE8Df5KCcdiUhMpqSaP6wb5sX3bZlnLuIDNVpjrz7Ia3oQPbSE14b8vSJeFyxfAaKJ365TARW
c5IiGCZ8b2YE7elqOvMTxb1TzJy7ZNOMu3QxR0962Z9rEmX5qZmH/qhF51kcrP2oOcIfhLGq1wCT
O4O3zxS5cpiYmj4YxaG0wzZWyUTi+2OCsfF3Su4r0sh+ARcb7NQSccPzwH8dq/KMX8SLtUWl9TkL
ayWchrXUgMxbg5GLD4w9UkPGThOL02qBhn7PtXRfSl3+tg34+VVjxenyBZkrJEqhLHDeCkZYpGdj
KFASplntnsnJpJ1h2Kos/eQV/hvpRzToOM+3Voq6HJiaq6izv7dp/rqB9wlk2sMcsDY6lQOtWBpb
nWRTolL306g/kEox5+NbND9+TW2ktZC1lL9SOEJd9CH0hPEa9oGUKSCj12lQKj7bS7sX8HLv4zE9
X6TyDjYWsXD6T/sU/IkDpQwcwFR6tBd9cSWHoRcwrUeZhMQSf+AvCaPj6FCiawE6q6MY2Rkf+gZB
6gEihv+xtUXIWzyPpWE+vxk3uvFp7vkXhmaaG0irDDZBVMB/fg2Qa7F6YQzNhpQL7dereEeXxJki
hX7SM/f88yVeJotPz65L3/lIJGT+YLBeF2JJqU9SBelbGUbJNcuMY3Iy70BRWOUFjQUdJUrUVvmE
TEIy3Zcgv3N8n6inKhN7uHV4xRIaaU5XE2eZBnYP0vmgDIHqfB/d3aQle73ogfvWM0SmTY4+5RA5
yKq/prMtWBDUWyUiu15niVkd/+twzeLXKwZ931k7vS0jRRbJoP5NXyrHYgOrspIEt5nqTSJPxvSp
/mtxXxS7b73yhJfWsOSFzKEX2PlGlMMz7hJrS1QGIrouB6DorQc1pA/Zp8eVXmkGWtbVj8cyhgL4
KunSuQfRqQN9CzNEGq1F11B9o6d05tzrNdqvsspzqFOYHe8ueSvaL/JwM1NS9NGer8mCFcrjVd5C
kdVEHeITwtWqXHrEFj4MUA1Qw3nd8FBFnlg1X0q3D1pr1HYIJpicAXT2ZHzLhvn31k4Rz9+3JC/B
ld3v+cSG0vCYYNsolaj51e8qsctyf8tAWBroeyIDzSTbKwUUBDbSo2I5eaOuthBnHEByYrbcSFwc
88bDmKNZk/fgbb3GRq6+M6McFGWbAhK6wqNPd+o5Y5JgmTX3VdhS+XLAMD6/RpEmDJUq4+7S9qnD
XOauSIlvHZ0CFruZeNO90BE6pKcFL9K2l5E5bSzHyM9SGvIvYLT54OSv0wuJiOE14Ol7zZGyrS6+
6Jzo4F6i0djv7Tdc2eF1BjpoK9SVYHLDwp0R+Yu6LFHuPzuXnbdXRPA77xBFq1Corxk2Hg83twSz
g6ai6+r3prG3JI410JxcqE1oPbJgcyL5Z8YmCFZo8X0fMmdndIUj7VnWC/ruTAJdzrsW8v4FeW2n
f+7VToAA1JON+ogwEoe2dFAbcbbwzoMs5HJsttJur48iAugVEB9/TJ60ZJdNQXQDmlUc0u2zet5H
huWl+BLEkFhVFlZF5DhQdXyRKyQJlqgN5QQ31OFIHURb4DhZ8zxkAFRK/LGIKVb4+ZVOCqCBvhtC
ZSqohdPTibzoxfoZC41MuMQW4FPlKE3M7H1J1Lc6LLvPi/xrsN43brafgiZFZA0jamcFB5xesfGa
zVYiEkEyOq1YyCPBQWN1l1T94+uNQLUMWdgDOB4sPBsihTRJOa6RcYaSryKhCtKJvNozU7KG/qWt
aWvD5076JdFlAm1jnvQJk+oUu2pdBEIdxP31v6AsWZtap1DRMLAEFdo9ktqwpIuU6vwJkIjSVQ9j
7qy9dPPZsNrO4fEW2cUfFqWj4OdK8RZO6FQqI/h3IUJVaKBwxAtgA7KIOgnr3o3rKwyx8XEEaJ2/
E3IZy5leKWKTidLBnztGj37jKz5ltJ4FRBweuGEWgdxGLCkDkzNr3T64MQORAxGWxw+nuEfTkwW5
OeHB9E56GV/gkG8QFP3uaHvyRyl4dOyVghuqFLj9S5a1UmT15T0awjvCzkx6t6kjs27zvbJ9lwLD
scWDpjAijp6vU7B2FG0Za9we8wvh30Knt0mixmh9h9dFJDw96ZG9dOCijOaRNbj6VhH+EZe3xdlg
oMVctXR3o+oxnehbJpf0isWeUxcKQo17rrkcmHjA2C5iaqEK8SZG0dt3J0XgLW8jRrV9eB2I22KP
RDE2jHnC4tWtq4rEe4r9TkUDvaN7mKpFRW+FeqzIl8Aor6fH5DSsqO4sXEWKhl1e5VMNIBRYUJWz
I2coQZ93X+91Nyf+3kSoLq8Eo3QOq5Q1LWqrk8MqbEtQi8kBj53hs+IRIbGYFX5gWNtQCz78db1W
eW2EZoZT4iBxYle9k3FuFA7sesS3Qn+P2EmtyEd2UJvgRVCpbvQnq/0zNmnFt6wkme3bVRz8xMR/
tdX1SCpBUAIq9O94WLpOO4+rI3+QywYHl0/gELVJfEU9G4QhORLNvqRHVF+RAGfA3ZdIJomZ+S26
zuJkMARTRB4DDkWyFDOJQDGLixd7NvZFyfEklNuYVF/yDDy9++wq+CTU+giRIGre6hebhrGtNQtk
2caN7+VHT8o819qy7tdit5yjLiZ8OCL6N+k5YuoP5IumOOtmbk79Z+ubpp8C4C+1ABsD7ZPMS5dV
MXPmQcBGz4lGDFadYEXcRXBcUuAleDXJxDLfVY9DQxjkBxvwyuC8opPHWK6073WDsInCpNIZ3mS+
rAKmNZS4553WMcWDRaLsNhjk9yVSXFSGLWianEph+xr6cTmoVAuZQj7SNldl4jhMn0t1Hl52aS0D
TqNRUcAce0AoFOUXbK0wSj2Snymcf8oCx1TCa98hj4lVs1UnhvEYsl6auOf3j+SkLAbHTRq6paaD
z6v+FAMcYuM6aS/ECC6SSBXKJlPMao5e6eIn7cHHnlt8XNFxr0y+SjUaAVy9SDz5/wyBFUSqbwFz
/GJn5YdbX2Ad0zP7PlPSieQs6eZNDOB3G0WFRpSX/C6b20HfTSBrAs+efoifB0kbxyHFD2ykJW2U
wz5v+gMwPPZIJ61stm6oAGDyFDer+Ghun0iCan0N5Zv7irdizeuXG3mxdQUily3yYtgVg5q1N6Ft
vo743aJM1yJ+/IIGOYA7yPIFJU1NYJf8xKY16ZGB0Sl0wI1Ju+JffNrw+vXeed5W/hXvsqpaopb4
mVW9tTqC0x+unRG0eAmjXhtGPKDZcbSY6CYuCfa33ePUZib3G1fGNR0G6t0aukUt5rNWEHH3xkxY
UoruCIw6oJNF5S3okzYf8gajHKSFkxeYcZyvqZ6DetWauhMIU0WYMZBYOek3ZXoXK5tVFGL0kE8q
5JYw8xuXB0GkK+7nhaEaghNrw/2ZWRYS1lMxKe7FJ/FjwKPgaPvWze9apKSFubxC7e6AYymcMIiG
GpvT5/+t1AVQOnKdPq4ExhcoGhD71H7fA7oyJMw7U8BI/gmj6ufJBEJ0OYEaH0naE+bGYM3q81mK
rQai4/f129y/djoXdBzIAMq6i0GniGNa2YkXWp2pn+4OJ4CE8vfrwHQ9HeI/yiLzrX9zPBmarMCR
uIzUqT1czXbq/WzGnM7k+v5sQpZCmwgYhK50cVh6f+Hzii77Cz8IdGQt7p8/RVA3mxruFVJd7eqW
KD2Bcgd+YoF9iWsbFYXo31L1gXDTM1fIbk03ccX7YjIJIcLzy2Llkxe9Vt8FJEju36WMlyHNCDgf
ox7Vep3GfghdRg9HqEZmVCmm/eImhyPKalkDdWFFbNGiqZv5g/fIPxZ+3DTms8mwoFNMdm5mAop8
J/eU4B48S6j1C4q4RzSxNFU3iL1BfPfhSI88oXmY3jBEVFF8XXyBJ/as3w8WlEV/xNgS4oCkber/
Ktg6X/U0NlM5UBMA5LA23wLcsJwOvv6j22HwW6FShInd0oGay2kFqYro3DAnRyEno4rXJrsUWvbS
Omgh5SfXF+ItCL/gnGgc3x68xD928GyD0jyYPWAP2pmC2Zb4nZgW5sUmsei4CKoRwHZ5Pw4mwqJ6
BLM1R3w79+T/h9IZvWg+MR1xke4/kMDnMZQYWvUxps50cPdvnliJW55ZtIqPwWpckMhCGjxYSma8
igKF9Rn7SJvYeHnyIZ5Mr05MJM2UFKPcyF5/+IqhQOzhkpFr64A5duWDZrGqGw93sGj2yuE6aeoB
Gr4j4efi5qlo7BPlPWphwwG5rRrWRaNQWlyfwQhPpQBrjKr1dnlggrVoLK7hkC/I5yDwSQQ26HHW
Lu1xIx50kzgtFDXgiGjOPRJ7l8zsKu2d/ELC6UdV/z/9K8Y2pGjVvTl560ajhc01PhY56xzB7cGe
tFmNGOUvxOtilMVx4agTkMnCk7UEnHYxh+etWILs1lc4a2TwP22NSdjWErYdc3p6AuwAuKpwQw71
4ij+1qr+FiabzAjA0aWd5chDYOWW/iM0jzix5VaC2zCWJV6hZIG3yBWmMxUdu0BfA6qerwb9s9MZ
g0RbuQj1v9xCLXPFh6CoziuTDAazFmG8wD85QGJc8q4M/Ct11I89FcZT4Ma4iOAqHPpdqHaR2sLS
mqMR9H2joTnFmrv/UIp110nnYstJ2utG3kV6neJbYCiUgDhGWOfS0LZkLu65x0Aga91zHaqXAaPv
UsjCwjpCfY10kQkZqnW6wJybEfo3EIosvsbOxzIVZdZw77LpyAmDi7kas5okVg1NE2ldSL4GbWsE
FhnsOsFHMoLFhfwY7g7XYvMkudtH68+HZF6UEx/PaY8z3q8q3rjPosjqf3gB3iVXWP6nS4/RR3KL
+wgrPLO90aJZfunNbWMr13Iil63qKlQx0R1keNxb1QsfJP8MCGnYJbE5i6yjmSL9+WAS6/hiRJTX
HG8N0kvo46/XPVOud1C1QtfSJNdmaVelVnL7fiP9Rx1E3zeAB8+LaKe99aHVsOWo4MsROnONNCBj
n98jZ+GJjb+XOtuIY2nT7zOOY/0wiC1Ksod0zY8LV89YYtvG55Qe2WIewrefJQFhEBejfPYBJdqI
9tAn9DdrysiXw/3Dbg0mjb8O2K/PQOffFq+NiZa6m2MGgPHAYeONagqQPa0GQsJ2U43mKritPDiK
FUkhIMBLyscb0m/CqBfKS+QFRQPrDtmDGJ/xsG+qeaE5cBg3//BhfuJ+s1VipcWVvSMx7XVaiEZp
Zi++aOaIFIxDXueo5bmjGB2uR3Y/HCsMOvdjw6nBCkh6G2xtw2IRYjZxR+nrnYXN61Mjp9MMefox
3dqGzCJwljZ2ZdlpCfhKSTheeKucJ2Fu8yIlGNQP4WHe6P3KnYTIu0gqzkCeAt4UA+vFgUK4raq2
Pt/ZYXpwIVfw55+Jn9RP3tiDccFPAhUEz9C8jx2tToIhjr0NOvYa07j2edHi9KkwKJCgWG8MuxtW
1WFQ77pbSG4zTgYx4kmE30IsFD6/qUp717IsdORYOQwGkqOzSAeHGzq7kcGiJNABuzW1jpFQdtPS
vUEEjzJkPO2hrXoezENrgQlowetFeb2NY2UDiIh3ZS8kD3P/mdCWnyl+jp+DlPSBwu+kvPdDYUYf
W5mc2pOa8yd45IcxPni8301LAaouoHmsJgfau/ez2AUM9mLJ0oTX5BX2BrqYOx1R1m0eg2Vq+ee2
kBs1YvHRpwVJfsDBl0NnSTDGFVkS0ReUFT9/9nW5GF0RKzcShMh7ciss84ge50QufZQ5+vjVn+Rr
gn+jk8xhmMjgTSwXonA9mHtOGUcRMyEIgrfC85eNrqwAA9mKzLPMkrndOJkwsFZtDDf/Jez2USS/
yMWiE14b5yThWu7v6zO4e+02gvbnj3xzc8gslvvjmG6UqdzbypoPMTikvx9NNKWqwnAy9P/FGn23
Brub5oQs/NCSn2ZNRtHZTJijPewYXaHo0P73O1kdE0hI+GCEEFG7Yf0sJdPg1PXWaeLCre93/uLf
zs7MeCYRcK3DUzzSHIoqj4XDYj4EkauU2n9HiVgIEifkfDiEqwjikgFV+6laS9wSn+rU50lUNGQi
CYso/lv3rgfKPVXzvvFCjFt4XYRaqVwxQY/x1fYUoHS6BTI7XXvr9r/r5amL4tXm7vfZc7b1bO2m
ptmFj+yAvDwV5K1yKqH2GULLbi6zofrGy6EbvtC/NIPfyH7u3jQYdMvIODgYYwUFkjmLqXaXRpKS
Qg4pg0PRaZjgReBtrML5e4+NAFcLhMC374T/RwdRqV7jkbzk2IMhgGG4Hi5wEP/dfdKG0mwgQSlC
grNdGdTo7JkwT8D0IWUaueG/RakVvKEyMnajFWkyAhK0KJqaVT9sjCGRkUJT/c0ARV/UKAcK8N5T
Xj+VRYlhXoG1gcaaSQpS11h4OOo5t5oP3H9WFkGWAndgZe3aHL0tfDn4Zg7DB9SqHLItJXUgM0+j
FDaCEE4XBHb/uTuNPilHZzhLmTG2VH5nhAhhddNR5j2JnybOuut5RrYGpBZMHzdLQ+XnzRq6ckk/
INGv8XaL5JKbM3R+z2KFKK+DUHbVgwPu8cb8okf4IAdScwrm02QvNGM0wnvQNzfxfF7qzU0tnDbT
bf4tkBfJgqCHKY/tWCuDefwJfz8n+YMuUTnCi2jW0Rhkpc7VNl/RuF967vtSqIkQrrUsOtrs32H7
i0fjuIccvE59A3yNPdbsp955+Tfk1Qpq13lIIzUYewnLPzs5GyF9fxrhuqasOh65EY7qXSo/0rNO
XV2NSQiZcA0TbTs/LiE1XXFUAxbbG0gY1UTrNGLMffNgZl3DtOCktf3mG/80T3Q8s6/5JNp15XYF
LOBVZddrIjDxxtk9ZU2lyvnij+37yiUmrNjAxjP7qSXV8RjzoNpSwQPJKUbysvkTZ173Q2IdNZL2
8Q3v4guoZvFKCVkqgdPPuvNUqgVqqB+9gUVe/Ye7t6800JCSvPL1brkmhNQsyUIA8+VkjQZrqVmK
ZtIBbRHhDIQPG++SvJvQ4csyaWCMTw/WSfG0BtlIBjOCC9iAXGpfi11j/HfRq5u76gHQVz9Vu80v
mgItZsMWDk58RjGwPqWnReXckdQBHBDUjzisfcqVHf1WSJlp+aQGdW89c5Mhvz6ytOZ9k1IitKK1
imhId5mAAOYeYaoqUqnobhqy4r729VOtPzlSCfGeBLiQ26YrMua92I4LSBuf+fkRebPuR4ZhUD/n
yC4SxrwlLSWu6xZJDFIH8BC8rNatLzMvtudpdKf1S73RCUIfd25DAZgbZkCpAhCLnUFS5CMZhJuI
9T7Dxu2vqRSZtnipUZSrk9wb5aGkk1iw53f+PBt5RwAJlOVLUQI6MDzdYXmWc4Hm/3S3ssjZFVRW
rD4LmfNtG7FANEppuhR1Mb/2oS7bBfQpmnt6fn3Na6fs66bzyPWV1JZImqvgrYpyiyS7z9tN/jcR
UaZHZ4quaD52NUTP9mmY6TU2HnPVL6xiC9BrKsQBMyoADPIfy1My+l+QXO/DH9wJ9vXwSSM3f7Fo
LXKcaIjGH88RDmcDnyyf+ZQxpjBmlPM5PCB+MNHstde7yeWHHWda2j0QkupJi0xQbTHz2lhGVkQZ
1RxOSsfMdSfLbB2WxVkZ4v+TUOUdO8APFvUWszUc/lbiJPgnL7IqUM/1CVfQ8eiAQ010OSSTR7OY
uLWR8SwwMT7mpcI4OHtZsfGQyHGDNoQYaDyf8gQpCHM4O9D1V7vfoBeCJX8QUvZI5cFtTJpbVkYp
4Y1xuMcy2iufmycC85zSQO5pzev0IWJqublPH+ttGdrY0Zod3EIli41sMtyi9JeAv/E5yWnZI6gf
yFhcCRwPt3xFTfMtPvrpJiwJ/DFXJNSkJOUsWhvL9lSvdoO9C7NIXd5G+cU0W+Edu/4DxoxFhJ2S
VGfOExpFuUfKBm7uESV4nFhCOU/vwc8E5Xhbgajrgjp9fc2iSDWPaj3lVJ1j6Zy/OBsCm6+/+VWn
/Iu7UoRMPLmOogD+6g+q/XbIaUxkrLIKAOuQOv/TDxtULj64g0xEoZy140mspcjXMTFE2owmORik
pjfKozVH/YYp82aSbR9UzAIu+AhLC20uvbO6aX5QT387/tht4iFJGEkbRbj2IQ/m0SP2syOEdfil
tL1pPnJXQVmEvNpvymwiIksPHLp8ngq3vMvTe3k1dUV+s33oX3tpR/DkTaGSuiZb8/4mFA9/HW6n
2138Do0aCT5VaOXJ0I822cgiccdUKJAOfGrUM6qzKUT0uKeEBMcN3SlfU/NIchY94qYNwx7hFjwG
GKHKjjVH0MM3KaejlQk/p7dC6/dx7EF8H7qXY3jBm5G9SjAxG8vRJLhSOl/rvih7FmVCUmW/X5Ol
ZmA++E8KEaaefId3d4WVfNpw0tKxav52RL4aQuzUPs1X6kwFKHMZDBlxznZ+rmjj/siNV5gVEvO6
NNbKOXGlODvDyDqwXQkRGsPK71qD0VLKun7mzBnuQlh1AhqXg66QV/2MUnTiEXx6XPCp9q7WgJbW
sE/HFdsgT9lGygmeJs/RAP8IbqLjqciWnGdrpiqslF8pFgjFm2fFWs99FajHFCz/4qY6Na2UQc6t
BJuBKmwdcBsHnFOHkpE49p6TGqPJn2UaAbB6uCmUDhYVmqU12DYnK/Ld9UeuLqzu+s7gsEY8hlQT
p9uA0x7qwdlC8WS3xr84HDYM9++ohDZTg4QGI5Y/q/ROJzaLaIjhIFZVdd2bm/3KpHszoOq4HGB7
nGL4iAC8nrFb/ppf2H3aIYIwY87i5OGRYPVyUCW4QMVHWc7zVS8JfQ/h5MHdjIPHoW1LTkvgKg25
qgXk4FSUJyanKbqlMNytBpskHE/awQhkfGagzznv9VtpBuH4TLgW8z2uyLmpd3j+mRLX9LGqEW9R
fLkAu7GMVcsTCNrsgRxAqAltE9bkWfNRiapXxraHHw5BLXH4eQKe/Of8EB6F44msohXT9vXVsCdB
VTZXGa+HKwTQ40XHHT/QxjMUb12dfWff9qNtWab+ptcD12p71bEjaVESdrqnIUUpLSXvyTW/ksep
Mr8qbjwsCNhWmGQAFdbZjuHJn34lnapB8kfBsYZg/j8qKuDKWmgqri1pXbFjSc+DbQdiB+RC2AG2
Ko+c74FYp2aZobwBmrbTK6332WRO8KLMN1VWsNqrkkFRNkDGJZ4RVU4+chlcbO5tYDXD0dOH5leF
SYdyFVEJT2BKNzy6nMZgLsAePpdUlZvn2HsHihiLFB3+8YF1NswJr8J3gbw+qHQsqviI2DyMKAhb
btTMTf0/2OEax5k56uzWkrMe7H3yFFUqslhSXGURgP6VXKf8qhgYSf4i+0L2jAQJnPhX0paz9kvy
i0LbPfQlBKLcsuehwvSjUZzDQeJTwrB8ahzfHYb+p/ui2fV7LodbZ1cf86bQV8y/PR2fJI4I6izY
u77xkDp/+RMwSP/tLwPOBm8vzzHCNR8qXsPHGAlgHeqsEe1G/j2b0SiBpMoRNVoFODLM2n00nOTq
b0KqQVAV52PWnf24YcfGGAqhMg3yPhMc6BC3Hs/Nwf0DtKgFULt1s4rk4sFUFlJfQOR4dq27Rlvp
jJRjfh8Lm3Z8KoSKcMvsqwmR9mLfdeDbG2TuSgOnMmmW17f0nlzUTWJCpC/Y6WxvkJ58GPSZR2jm
1/unzC2CfWzLrdWbrXvtWSsDgA3apKQ7v13fkSherjbxCrORrx01oKLoXwC+4gu/ja0hcfzdSVMt
NaOGjRN6JZrUVThDUdZJcPBQsEvuJwChQlBQxVkOxhnaSzB0NVvlkrKqHybHArzfK063kOmOSOVr
wrtKPtB6O+xgb1f+SU/dq+bHFYx33hXkXX7OZxkv+y28SQpvFt3NAIhU4KK39KXvy7WU6R5SOE4b
cpFKBw7ZnjDSst20Dvvx7puKA83wKoOJmLGfPRJRMmQHBdySHqc7SB/i3DMXiA4VQgzr/szKgBJ0
Dv0urSt7R2kziyl07QIVOM5C9nXPGF1VVscdicJOoehsSER2xR7U4DcIswDmk+ksWZHwpO1jnGYS
lYTAfV1IoTNANtj4biquL9M0covZeOkZzXG/a5+Fob8gkx8EWssKIR9o90EUWbodEsbOVE5FUhbU
uG2MW3Nn066D/j9PfO6Gf16vU/6KYP+TpfSxodVDSD6k5gyXfSyBMvtrsYfyJP/3uiVSwYNR1oGs
u9g2obPHwqfh0fVsKGu6mWNVwQl9dXWIpp5GMj3HWerdlFzudRYQDK8NM7UgKfwJGag66q1ybFA1
41gf3hJwSoDedjrVos1xoNsqsb12OaI/VYOLvJVEjNDZvrwLsG+GFSaTky64Ln3ST1YdfRg1ovEu
WO0ZHjbqDZNbXLJfrBCVWpkAhejT4NoZWLvUO7dZd8e+WhPbLY8imC0UKuToCS74gNlsnV3afY+A
OXg1MC55pMKTXjlS+bIDClgh3+GJf9rXv4J3ZiDoZ0FxNEkT5/Ybs8kFzyzm0x5N3UShoIpu9xGx
RGknwYScJ9ebBxKBM8Ep4EUgXaHuP2bnAYsoweQY1S5sO46s7LPFQguoRIPtXLIe40DGcs7T5npZ
khVX7+z1pIIYgv5HoKhkAmeCW0Ps9tDlTyCbmK5+XouWOwcB4+/Gk035Aeax4978Jf+/3QU17uy9
JGMoDOwMBc//spWDDvIuo0B6QTrzayR9MMesVUYnuGNJtWuzR2gQjD894XvsENwasActr8jbEz0U
zmPtHQ92CBKF0QZaLqvvuOw4qvN11cfLbQFWnEw+JV5oNS23VnqKkhZLuoDWIGPCktFJijbOSBrn
3PAkJxutpxgSzn7V/iCt19mdmgE911vrOZwxE8XZ9eSuTwLgv8R9hGkRQtV/9c9PHzB1Nsa08HtW
oMd3qkJC8iAcCCHxb3oIU2vXEVmHeMECCL4ZCmN+14rg0SX++esHHLiHAuG/laOR3fZIGtcMe2xy
Z/XLaIIYgwk6V20vEc/pElssPg4YcpM+D5cAR+uhj9F5FmpgHpv/vSgkb2JjMfj2lMC5BFM0lpzQ
cz/av2ZRWIqu6GM5KO6H+nCkiVboZxI4JU0QeGmyzvTWlUBC9KignXirasgkBqubVvBWpwCFhs1C
gbGDL41wjwtztBu0fUkd7amcySQ7R9oOL87usTV40cw6IrSjzxAK73Sr9ZsFh9Pd13VOnhDtJ3k8
xdtzFObcVLAwauAPOc6k1ugKffqdUuHX07LPr2KvuKoHn6CoaXunFFmi7mZspsSmo9Bb1/ZYedW3
S6R/Kma7169KIKzXYl9T5maQR4kBHHHfPb1hVZaTvlvWk9vb0sexy+wmxkoJgKHj+eB8RfdNLxgw
hags3ABgl3BI+h+FInhG2zkEy1PJPDpc2zzkIzc2LHM5b95Ib4Nxlb+6HioFmvzVa7H53N3bRMbA
Qtm66zVJzfPnEeoyI7Z9jOGF9jm9A6EmI8d/Oib0WEmdOfIjGFk3xpG9hLlw6CTMzdXi1vgglWI/
CY5m+BQdq3tI2pzLnoSsXPurIMaBA5wOKe9utpbCrpQP0WSdy8ijd1VboWZfmtUH064iwGipTbgb
Xk2Aj6zzGAsWfQAUrYFa2oRDg6FlEbYmTmrwTxozSqlAUZEXbXutcX6GMgpVNIth6AaWY4ilMOUO
pxSa4TbiWyMeSHKCvlQrrdc6l+0Dwav7G0P1SHIM/gXRzL+x43d/PMBGufy72d74T+M1nvcREmRV
81tShjqAjowWNqkVZRx1lQkJie/FdryucSTBLtZjJ1y2wKTQZMXVn1b27GXJutU0q2qmS3oo4mBC
Obdy3fFw7G5N5jHrfPLHdnLIt11hsCLACgCMOPyaLjc+OCk7EHD+aY30QgPiYU7jAjAVEKQR9GLy
kkqzCk97K/Xt0ealXQzcudjLh5xz2jSFa00kpsdmonl0xv1IC93MjUojWJ9Vjz43/nfzuPNcDAbU
5E4Q0b2nZ1T+w+y/TavP2z5ZBrxoSZOYlTIl4k5Zvx1IRD6Odk8aATEKq2RCHhXdhLgkK+u0d0rV
8AyaaGUEKpJC8gxFA4jc4lhyiVyHSzEw5bxiExSa3lMb4q9XTYjIThhLY8k2LhvHHqL+yFjFcFZh
g4NgunZlFv3pXaQTdidiq5O1GqEQXNvmFdrnXrrXsxWE3M9xx/3iJW2YtcQaKBOnXtuKpsRd96w0
UWNnWnERxltKkReF5XkBZmJc7knf85kb4WcWsTV5J1see7L+/GDndDymoewNJ8QzcwhUf1PlaPeX
mpAriUOfznFc1GavF0PLGlzWzWCCkPdCa/e52o7HBy/HpJ4mVXLiFJ3ZWvvRPJMVhALEhkvzQYo/
WBamcGwpTzJU76qlX0eyQ4/3dtK8TFXEbrjub9CbdEHCbyoylJXgrezSRyv4lsTX/YJq223vuKut
3ucQR2OK5mbwyzA5q9Vchx8REzNG5zXTq1NL9jy1BhxMkpFSuYtpx/hYsldZNsavsFabb1ZP1Byz
Kjq9PrcRt1oEPWts29Mf3pVfcXzVrogh1NT/9xoeeqE5dE8KFsF33E0X2z9W1Is7nHptq0Oax30y
5JGJ5TiTPDeIDYVgraAvuUArSdOa1i59kH/kSM+q8aJ2/TG7tQzFdF3l9Itn9oGYBZMUv5koSJ7a
pJLRNKRe1xO7bI1DJZzkBTb7M2Uaq2ZOyftF8h+A4++KNE3tO1tF+2u/xnRsqS6zngyQIkr0tW+J
AcMQbkqBJj1u9q97QY7+kdOgaPX4rtsgtQKlfnP6vQDPw56FEnYHvt+p1DGU3U6G2lphXWay26Ac
yn8VnBrqixYmzZG2WrCwm/qpLC8e9q7X5tZMvltUdH4K9EVezM5v8BRU4kRY6PpTEcUi6C9sTWLH
7JGarH1WryJkBXAiIj81buhH16AVubK1IBKUJKeUxVIE0xW3uqQUh7LEG4Yy90/vDC/Vf/pZwmr3
UWtYDyDt3EIV7LZRLj+qCQM0XSRQLZ8NdwANRUXZ56Jqi2X1/W+TOlppo/1n857ikhQFzD2iThCa
9RmjAOs+1swJvxRhewWbDlugW5AbJQkHCCT/Jk89ZCt+HH6H0gMyG1LcJGipwbNOjv7udB+/uo01
MZgFmNP8wnaCR7PqmDOGqVR4OQHEc0AzdBLw8Rh9O6w37zhfaJxTs44DULxDBu/C8/sRzswaSBsu
G+lv5bLHeK3ZoYabE3XBpx7Za+omjwoVFemBULdPZ2EWlAM12i4uV9YkKVxRBM5fqKqFNOAVpI5z
DQmAiZDshg+6Ef29lLcEpaHWvHAETkscwbSCCmi520A2La35iQrhK31j+nSy28bchyTSlYVu5BCJ
47jaj0OX5t93m+CjApavkbQ4Qe4nXcGxUV2wUjCiXCoWsyVz9u+HTtybnzKGEbx+V0EHGFg8+drl
Td1IW41dthMJG8xmnSughEedl2ovemmggnQaakvsFjUWelfEfYVxmb515AdRhKCL+bXj7utR9StW
mfbTGd3niy0/WeIKCAdW1yxY06GZKjet0oR/OezbQnrCvCvUqDdMLYSfhp2JgPjFERLYEGQM8dgE
DMnSlxL5U1dMA8WIQDKQgybu/R6Zrl1uJJ995fP+fdq+11TjRELOxERDJovj3tY47BnttJDU4wJh
QSXx1H7ycrTthjrb+LSZzxwxwJKVfLaFM6TVTcKXmpibMVrYZxhaNAkvCrKsSHUWIAUV6GjtflRW
CHZKZsjKC+gBS86hHemDI5XOz9/KMv4+Gg1S7n/uhngBeRrGJgVl/1oA5X1+idPKzN33lsN501Xj
Q1wwRXLzKY2y4Rk9cMP7YAHRYV/XAssvCXePwjjiaCV1/TJzgQM1x8kyUBddmRv13JDtQSocVwa1
Ir5x/5Mr8oTqnOnjpXIMrVUY653+ojUsgPPwpT89Ma/fqTq7W9rXosI4t8cswO46yYqadq7ta88Q
WrGrR7rXiIL4PwVSBIeL2hxeVJH4W1gAgxBPYpLb+tyRzjEGvNLHIwdwSiU/NDuEyTzg+ppbqgvm
Uw1tIlhTPzBq2IKtontsJwd7CvojIk62fYjhMF9pxv91e8lVNWw/4enK6FYgwpYgEYJtvmyzf3E1
Rf2uD8cF+B/m4AwFLKpNM7Vcy623TNSpkEExdGBKAeZyNACAUWhwOtmnXgw9rq1xWg0UR1pQythC
IS7ugb6ejFHr1Q/mtBjJCZYIkTXQD0wwskMjITrk2cb1o2tk/CrokrG/FBqneG7fmVaoa/VT/Bk9
Egjve6yVu+xOWcwaRyBC1O28eQ5bXaV41Dwla2Fr+oFmq9Df9ke4TJgk91Vt0Z8GkW3tuuvHy1Y7
5ZkgpE69MwXREPqpe0oltW6eULfaRSpYuEZf4/ryLvwAnwUc79zhdnghB8Ma6rp3XtXtkozOXlRx
EN5AogS8lBsDr+zTWVDaGLyRNilkyFNWiA/p7KQiBEZuY5mMu2FjaquWODr4+pwes77CCRxIQVH5
Gfo7KvIIMYBKzF4Q5YRZ7X4Ex3ObfQpUlh8hT8KnpDk3LF1r99JrxXijzbBQro1Y/brOQBzZ0J36
zaWbel0DAxo0UXZX7vz6ziPJRTtTW/o0gLKBSf5tej0NpXkYHvpn78jJL0u2a8/PmJyeWrl1ipv9
tsjSYP2/2NLHrpu0YIh9cs+Z4h0Rv7MseCzpIFuWEl1RTihq5uGIH1SHreX4RXhehlSTp7L6aiu0
2wNno0aOKleauuW4ATXvhG2cGyaeXnitqlA7y0GTpJW0Pz67Wq9HJcWKiyUj6SDvykDAN0Fhwy4v
CyQg/dlBEv8TbY4iWLC8pJvMOwm6MhMylv3aRw64sMVQCF6Zo6DhjEVDCBcTTHgXtFwsRQQu2Dda
UhsQ/uxTUEcU3klYPLnPKmUUjGwYH9gMMTAXaBMh/HBskOcCyOlNa0TDu2w9RL13pvwKIzSIC0Cf
XzzI9zQwTb1dJ8V+jJcTg3LGB7xUcIR+bmvso4tg0sIrosTcuexHNC14D1mCv6i8ZU7DnKxbL1CO
zKDQGpT15xBn8cla7EukKI897o2mCiZGS8ON/8TlAL0nh/Q0QmB/Wu8DrHeysF24hS4j2otk3Ex3
yz9lkmUMj5L4vgHGggM1kZKkaTqexg0IM9+SJksDMppwQeeXMDjqyctUY5JZEUX4FrLRslW/Zdw7
6hvqpRbnldUuh+74nEjmNWBgOGiaaCFHED6mnQAABrhsGbNWK1vdvw5KbwgfL21YYBSyc10JdOGB
8wodE+nRduU6ofByivp9FVNS74gBoRHzp6v9qAS7hK+DKYFDniNqPLzIgU4xRjAE2Sq+YWJhE+5n
YPvXf9sjfBen/hsRaiP1v7gy6uKtO4hK/ZDmJuWJUIhmCbEjAfc+HOeBxFCbt0vkD9ZMQb3AxnY8
H8RMdBYO2eObJeLti3RD4X+U8cajh/dMtPMiy5Z3kLyqL5XHVOGMlVlnUhACoc/zUhbycciNK4ek
+ambIodX7AndiIFyioRB1PM1NTAUGrSjwJDiCaCgTiU0aYWQYXDYNBOF9bcDM3eERM9I7elpbLD7
eZZjLbGlVx6CIT10uT+eN7spq8xUz3ry1SXFChr0Nl3Ab4SDmuIToukR4VYDXBM1/Pb04G3izIqn
UQUOH73ar5tz1f6ASP0zBmmOxPqDrATjhl/pUQZdiMqjnW6Ya1JdHrqqQRwDYAe6fXkgOv/gVnNg
a0uiEKxWzfj1GchyXjIpdb4VSHdEYO3PCeYcSvjfxkIvQ1hTFEwXdBKF0dR3PcDIqiKskT4CkzMb
ugBj1X/+IcVNEt2GIApVW6kx9IghbhjGi0j5QJCq7jXad9JK/nIh/99u6lrf6DJK0V6tqDd5dE6Z
BJQsYRt8vGOajfQe7EPd6RbIeAvYa4A5YFoAn5k1HnaRw/dK7CrmfrUFTJTO/jGFKyZtvwxYvGB0
HoIzVoIxLzDvQr+b1Rj2cPy3TAWhysSxaCqpqR3j78yYnd4mdcDNgE7ioAx7PUb8Pdt2TytKlO+M
nDMR85r8dgUsCIBe+xpZjVn9GRSu8yQVZs7TKauiUG0glJF+TY74U4QvAmdhmWcrZQ7EfEw58YZi
a5jRcJbRW4F32Gp+4H8pJm4WYuMh7fw6PLzX1XUV98n2tWB75fjpRtDQD+F1OaEZc4dk4eGCOR8b
Rmfx1scUzAcmWjorUZzdaVur6yZMXS+VBuaMlOgn+ltel4gz9BRd7B+Cy7SgOQQVs21OXJCimHjl
tYQMs6THbXun3E8AQHzhtZqdMzvARsX+V6/OVNaItEUXXcvnRw0AOr395rc6MCbcy3eGSWUEerm4
QHID4RySXTDOEwWGCsfoptmTpC4d4bCH+USxG7s5UWN420rKENyEoNDZyxZO+aSiK9P3q5tD7z/I
FHcAY6a6i+1oDE7Se9ANI76hrEpLIrXCFgnrQFd8BYi7zvsjbRldpnhDo7H9UvLuiDwZFUNO+pMu
HKsn2eDujPFMt9IxsAtWX3PffDEhbr9lXavLL1oj9wJbP8JehAhwXSjwjy9PZX7bMop/k3sVEJkv
5AfzUwCIfh3QtXrAaTWEPRoxerogco2ppTAtVRSTmewDXIZ5OVcIlmtznJdeaoxYX6r9v4cuRlW6
EaUzGShJR8GgmrRaeidOKnZsGS1TogVcPdlJSIBKF9w8ak7BPsq8Tg1FUCwTDmPytN2VCwVnOTJW
ovo4jl8VL8uK4Q+vPRPcEUsIaCPF6CKHGoI6yDErEou/FxoiYYOi3VhV2xDkoLDF24wPR1kWj4bi
m5RQQylXVscKkMKckCSYBsKpmUnYChxmzeSBcsoPiUt4WSoTmEh9y8RyRvSzIsDKMBAXQSEhRDbS
H5FKeL8qzTKnj7PGCPBJmbITkCJAYwsjLhVKpgbJb4LWcdUXoYh2e8SCGBRVOV/3r+WvRBT7Xa9g
So9sud3Z4RSwVtVF6/cbsSQTQNjtYOsMAgCWXb8wkUnDbHZlpuNjIDNPb9aH5eiwth7zgjmZHVPc
1ZJH3AaHpFl/trFB5keJgFjOPkjMAoUFbbPyvtbW4cW64ql+b81j+1iLWiJ347vB2XKWgWukzR9f
25GWUFe68lHNxO5Iz+Jn5f8ABtbWSyD8tDQgjNoeCs7IgjN2sGoCXsP++GAZnzGKZ89lQBgl7rsh
PwAuT5qT2Esyovtq7WXKk/InCuZ637j8tvwgSwBf5+OsEjFK08vd3bNq7etGKBT/+Lk45ha/IWm7
z5juW+Sj7y1HxLE5U5DuirEUygx1riIiz67CBgIruve5oXGI9DcPl88CLU6eQQrP4WSziIXRGJhj
KvO0Z3cwMUG1X9xx/9fMMsd4421wLhHsJm0Qbwzfem0tAtK0+JSUx7sQyOnzaa7X5uiut1VraApl
osOl+h0R0Ra8TPoH27hNwS+pUm5lpk8q5UGx4HFDfmfu7jQ0ClFzhoJ2CB0IaKbT1amhPlm6pX3I
qrAKulpn4EQ3xtXc+aH/D8Hmf75WZ3/YMpLTQH9gJbNJXA/9LfVqzS7CshnEUEQ1e9B4xFQUZUCS
tx+Nj8VGDawFZTxtA5I0/++kLGNhsFHTfAptmOM7V/XV74GDSoLMgmTx7jPjTKdM2KM8plPhxiUO
wBsduWWWh+M56VQZ3aZl55hGxMCNDafr1v+n9dq7x9hdsu7+z8c6J81+plGr2tku/kfmX+tEpA9b
bhBG+ZNH+4j3p8I3EwvatoFls/qWoa4gH8twd2niQBBceLiVyoUmj67FRF42jiZoHkefkotDZTnF
dvhD21LM7U7V2CrlIt0/0j4ulopPE2U5LQnCc0n5pNMwIz8IX8YpKMBQJiUctvVlyvap2PJt3u6k
VFKIXZrXil9VJA09FAVz7VD6C+EcKd1ztt0vHi3bteENKaqqZGuyHmYfJVUiVZFDWH8UR3TwAyWz
GqJwKBnVcuM4SqOyd2nGbVaAWRiRERcY3DYSCLHrgWyZrtpcrvyc5/NyxbNLLwx8KsOoFaX83tfG
mUpUmOxM89odQt0zroo9n/UqvEahArYBj31PmNmrMCN7YU6rSD1y2cYXycrq8nS3WiyG5sbC4+OQ
CcCsczDL23M1dosEYbaoBE64bfX9JdFObfHrz9KnLBeP17RwQsDdXCump91mVn0dZKz8f+fIPjIV
5aZO1DX0PEajk2YrJXP6XFio6CfcVZidcLKGMP6Y6dhZkEv9bOOcZ5DxvNOx/wVnea0T2QVIr/lZ
nTFtzBb3QEZExJFe2/8Cw9BtNEJMaLmk61aSiZG2jSm0yiOIpr/1VeulTXuFIG6kbvu+I0PqNKch
U74l0y1W30KyHVvx100L886z+z5vWWqdFGsOWGl0oYwh3tXNqH7E40vAI9thvNugxuxC+Wzwb3OH
Ab811Zu0CT+/rmexwnItqxrf+I9geG9HXpgV0wiH7h2qxXbu8+ukyhAdf1DvxZQhp+uT7vgoohwb
cWPouA6SlTy+f/WqU4A7rtu/QQukynCbrX+2q2fMp0mIJRKILlqt0Ppr8tSsC67hh6TynDmni16U
fkooTXO2NeMBjS0/kuN1aN3HaD8cS6srM6y5fxm4VENwUURdykZXs6qL4eGfrfE63ZcyiSOQlxUe
DZGOfr9MejRwlHVe/8SaTHu5bvKafGxJ0pE2oJMx0Spb8LIl17MrzxOTYgYcPsZ+yvh1QWXYL8OL
qdDt+DenisPT5u63YAjs1/TSnHeOz9EEYLLJcmZO0GK5VoxD1DKG4yZeDah05OSTRfWycwHlZdG8
0/hAH4vNh2vSFHCAIzVjnTuvqHARIk35jMAGs77+l5BtM/54vBp4KtauU+jTg85DpPWeMr4TFCex
Jo/WU1kyB2jgqGWD1rLpH+6Eesn/yZnr3wgE85eWq1t77VciD+Io8VpeaV+Z7tWUFCee5SghNhC6
m/09uPoVUZMUONgOzPnfUxjvvH9yi57uW2Fguiq7aPJlw3w1bKaTBnwGWMZRFEkEn5yLpxoTwrmA
q1LYxx+pHN1TBspvpkjKDd/ctbj69qeEIlc2ZOHaNXnyMGroazlsTCynTEBEv9EIf8XabMfPExPG
1uhcpFmXlmvjJkS6CBuDw76tGF+FP9l1M7YfArC3pvdzaTGigzm/Dsi0L0exs5ZWqYbIAKWrYNjm
5ls+XxR2ieHmBYILtWQG1p0v9lrM82vqjczK+HPlWRGKOh+n8J5NdHPnezVLuuFwXQcYj0jTOuVv
TNNYKCApBQdmXa4sc4qoEKsXtI6tCWeuh3kt6X5wVOEt4jzuKU94YsEB5+/OBOOFK8wfkcHxAoIj
/73m4fIKv3EGnADurT6M+WZ2e5r0CTesk8mR1XEEalqSqotl/EvegusYOFbrkbOp6xZkDnGU7ktS
owSTTQ8cd3M+h+y5pn95JPMUk3JJoONK/rns8NoFOrxuDRgVi4G/ZbJIs1W/5m5faydndXe/WteO
zv5kco79MQ59tAd1poK6IJ4aG+GUD+UjO1UDpw/VV25imwr6/tENLlPOrObdkyP/u7Y5an7izKwx
pTrNLNMJsmkqLcG/z6c+gwkk7cdsgOWuOoRS9HjZxRqcFQMD4q1+i35sBpSpVzT0w0HtDRnZ+XHw
35bxQCT7+E4vwQeD+S0bcohx3BOGfgXq4dLluBH6bFvqc3QBTIS9j/X6/iKOz+IQND5qngQiZTuU
FgbuzRV2/ErW+4KkyLAheQbuDB56/kamPYqtkrsaIJCW221deHdF8/r3861aU51xfTGj+6cEG2W2
sKxgsPSEEqqie0efHfOK15h+4X9Tut5s6jHoj5SU3JUdJ+QkNLtiv/jx6Ibi8BWuUE4Cgk1vu9Es
CL4bYaywGdS8ksbCzbdG15nm1H8HpHzxHN+kAaPC9xUJnhZ2WMwSu2uREr4Spxec44cnfVq+nl+f
jdo0zbnjOyDCct2FExHj9dOX6txZJ1QSJJgvcsbN1U+uPZPPOfr3PWZukmo9z5zgp3I8cF6POvK/
ZmQLJ/x6OkJZWlWm7ldPwdQBs0KbN+iqJcW6VcdoTqdr/AEby7WIFE5q/MxZP7k2aWwIiBMv4uMs
CeS7iIWqNnlLeNKiPp2wWpGAzhzioAnZUVVlBV4XoLTRk1diHOtY3uMSo6G2dZwoD+NE+HbYSjO1
T1Cj2rSSUjMydyjESOSJmoli/d9do9aJnclmZCk2BL6qc9jelCnVWjl/z98K9BNoZKvSLGancX77
dGd05ZbiAOoZTPB4KLs45d/Zcv/qy5BJHM/U2bHKhTZJbmsk1Kt/lOSKgMuKY3CNni3QX1dyjcUc
f62aHQHMeUC0zXCg8nTHNEt9smCqpbO1qtzC8EU/7NBvgNO5qmkf/dLotNX7NwTNkf9pXcTBoFQd
Q8lJNyOGQVdtdVoPrIeoVkJuq4M1LzXFidPXI0ZJGszuminADnmOgCfYXCwHlPM4PCFbVCvwXTe2
s1Ku7T7ZuA4Q8u3BDa8vpKRVL7hoAz78HqrdvwLxnQQISEm1nkoCof+pedbEwIiYaVDqRVOQyQ+H
LiVyA+cu3lW5Nj4xVC5hj8thHq7IeRyD3oeuAMAF/8noJ+ighfCB4MlVB+w8L7O+t+aFPH1UliMw
8BDxMdkAppaNSBXbR9i74+Lkb9jtlKg5FZ0zIQvTUjtjU5hl+lk8WQ3iQr2yrRAZ8yBdxssSJy1f
jzwwQ1MRlFy6DmLfDxkgK/P3hMaBaneDpsR1JOtqIuccKBaE/h42jhXmUnbpnEN1FpcjjrYeCLZp
ap+rd6sAtuWWa6653NzqUVnuMEVv9pjHy1zcna+Wcp1a9oHewYLO2TxqvrROQgmhU/YfQgeiIQir
gApXyZ/sjxjyWMHpZys3B2B6UoX3wIkGTDvv//cv6MJ07Y/oL8FW0Oy/HCB2likxqyyGRv9hrTX/
0viB3m6hthNmP21HcmamGZ56eA+tXfb05RLye3ZLuOcxsU6YsEHO+2VEX0BXV8P07wdmZnFNjXUO
eATjjEWpxY7HpIkgA/+/H7jUoQInXeHYJNFMX0MBm2Roz1Zz8fKR2GK2ZuM4w2bTr8cXobyJIp54
FuDqsi6wxOYJVxc3eRs+yqx0FSAMq4nx9TXyAMN+52qoQraAI5LUfRVdm0qL96mnnhno6iN+Le25
JK+qY6EoTJfKRORqyldVVvIP/QYIqLXTXeYufM0RDGSOtH9M5PAQgTiBA+mV8nZleJqypefOq43E
3AnBX29dLZUdbtjlFl8wr2L2LDA7xyGzDbT9ZVSYvmGq0fta123X1mgJzd6j9TE7SZCGL8H7jnwN
WJsW9yzuK+XQOu6cski2Ne7NpY2B0EMziVELeIOrlhPK+kWRGrkRC8/iINUgqsXJ+Bj/LCUBt/hi
nGN2CVBCMzTGpSVj8O8g5DkVf7+NUS1YbPmVXb+KsCexZqGUsz/gAhYxdCzjoQ638G5pysJAiHrm
e2h1NJoZtenvFI8E7DEmu0WA9siIYgxL5UpTWe2i7qopjfp/f7nmvVM0IDi4rd+QQHVaB4md0ulg
iqC1cVvIpfBxCa/tR0i9syHQd4VhKTWFBHE6xZZ8dmwGCswH+jx1Z59mhIHmhuZOsBku74h/4TLT
tVUcGIBaY39EwiF4e6jtWRS1yFAjnxQgeQtbTL/03fN/LRYJwX1WCC22rQAjdN9mxyDeKbbRC0RE
TeS7/eB4zI4qfMg1AwEVZb5WHlXpMjviWTBBsa7gWaPsXmUHHbpWnHe63AZW+2ekJRtjl8NuE6Gt
gMEifZkOAXqFd+lLMXkVnF/m8VrpK4BFPKD7GnXYeEbwAqPHAV/uSUr1IaadTlyix9aVqj1Wpp9D
R1en6xzfzcAA5FafKNMqzGkZHgCpD2DvB4iWGqvF+kCODdVA846ePq0JZ0XLCMuYdxYMHcwXW+bu
EvITA09ISx6vLp4S0tXe1G4Q5DLKjfJ1j0LDRhd8/UbjTsn7PLlU2TyChuBPEWs+9l7eA/cV3GJm
OR+SBvfrcHdv/o8guuiP0BP99XQVIy+Er11U7YVmnMjrtJol5ys8t8WYxnihe8jMA93PEfk99mV7
1vTUMuHMYu1s2BzW5CXaq1tQ2lhtvXX+rRbwSCt8TgHGrsnIh6PllYUWQG03vKtDRPkKBLErO3NF
VYTfdShqnHLjDTynbdS0PNaANRdCH2YO6DFAb8xiam5jj3PJmt6ZaKc2Hz7f1Q34xZ7PG7Yiymc+
HsVq8e/R1YKCqcPDJz7xnEeJ0OZWp96wbMZRZZwICvivz6Fy6x7mOYE7QNJrBjIK8cEFngtQpL9T
cANOiTcjGdA2W1biGhEhwA6mTorEvgOkeya4fNX/kzFjbFn4OaKWhPLW+a0YK5EIxPhpf4tzmtrW
g+CiG9z+tUiS+f32b6UyrceZ/AbLL6FRTtGNMiYpJlStOFgdVSYrmsnlI3t5XrBSwyXFNCovOPu2
at6z8QO1lGq9MaR2uZY8ff0eeP4IPXrCfgI4+RL978IDpu6q/LQ8A1vFpug9N9zBHcSQhUzdvKvT
NJNI5dDWh9sXorrMa6BdYgXfktNZ8v6l8yl3EqQ3hh0lFzlmvGGnVtZijdWYIqcvX5IiWJye59NH
nEDTI/rKrbiZWLhfHgm41WAvaxuh7K3bLBbMtCt+3iobmYF/zG6vMO/ujqQpKFL/IiDKJ920JNsE
UB7vPKYA8t07gqN6CbffgNfRro8mbOGYMDyGK8dRTpD8WXmRgQXQRNuzOm/GXhsKhlnzX863OFG0
U9kFHhQQ4jkuJvH5dpFsKoy4KjX0oSE17pBaLrZ1bcTFWeqajpYZGv4quNu3cwUMIzWmGQFFj3lx
lF6zxt+8E5f8mQO3k9xy/syZ66oCUyji2SYtDDc8wUSviqrQDiIH1JisAjhXYYjuRrDcrxmqrtHk
UjS0+3JtE1aw3ItY595Ad3E6Dl/itfgYsoiCX22Ew03wgpyl4+FFR9aKuo6yIUVNFsswQ0sth1ZP
gbpeoJvU+rhCmss1SLfQqff5IvsIbEExujKVXMZsVj2Bd2hU+M7L2ZUxG7S0WcnMcv8TDJekYsoO
xiivmT/XGRiBXzO2SmYosamEjW26k5rYttjauX4TjlChdiqwiKoaNGW5TmuF8+Og+f+b3enoz81S
pRtoBMHnjp/PkMF+NnAeyNQXli6DEACofw/eZbv+1s8tIsdPnchkmGrZAPdUGLvhWTBFf+EL8TmU
C0GyfjQV0lGiX5eSmPkFsUiJuyg0uVtH9sA6Xpt9bXfiKsgti8435+YOV9bG83YY871GlztFgoSo
YirjDGz1Ukboue6kkCx5ZGGRAYdoX1jwuKxq4WyUMhrC+qX7LXMCfQZ27LQFU7eIEv4A9a6EFxKr
15O2XBRMxOc1mF/boijwZLQ0WzYoimYQCNaXYL1O8uJOE38OrvyZd/WUsJsLmOIuHl8HIrgwMIpX
FwpfL7dQymXaCNGFd4vTbkfPO3ALZnciNSUCuCRYa+tyNuZaT360FphVimByMctC1qbjNmmy2SaC
w1+SzWhg6/+JG+6NRFnPc1oluhQ8tUeog3GhADuY3UjMER2DEbDHwLDHl/Z/OlmMYmmr+apHPiCj
zD2tlPD9MxYnS8C6+zQO1srzw+NuQjkml5QgUGiiugMlpcn19af27wguVyuQzYG/8T+xJiDroTkB
HV9Uvb9M7nHgBwBkvfxG3Fwu3+NAl2UXZTVx4/MdHTDRWljaIi0u+/S1M4J+++0FwLtP8OwkewO9
FLipvjkMFJm8KNVBjj/aiUreLd9t4Yzu3G9JsjRUtExcPLLTbsji/ADeuIOQFKu3Gb38GcGick+/
Psw2wRuclbWvVyIOQC3q7FLUM+iRp2rDM1jy6YjxB/vYmKaeIQlu/Y2HoSGCLd+ZSAXfFcA5Lod0
llGN8oBrVr7tNMjotFS84CyAdwsjwNRsDDxKxnpsr1KL7ldXXjdxpzW4BZtS/zx5n2wfzlInY1h9
a4NChwRzg5u7Y39VoS2ysmer9e/OMSy8kxBujFvU7QZGty2pFbZ2WMcRja4clc+loUOHKdddseOb
DgxnmpaimgNK7GYEkcg9WAkzaEeZPnIH2LJESQnLnOdUhDXzUu3E/MiUGsZNj/a8SF+v32OjoKGN
XrDpX1V9EQeZ32jHVADEaoJhIV4ddWn+5S7SY5meUi1fEqJKwFuuegMJuBlm1F4yH8YuDdOGAbN9
jfjjNQNcPo/59/vGxNGtJCQpPrO+x43yi3JkIFHRaSJl8jvNTk5TF2soI5TyK86ip2vy4ckOkbCj
eos5bYWd/Xv+pJq68ix22FEuke4yxW+fnhHE4axdvwvMAwi5cEyynlyoSKEbPF/9gn3JPnFsKlPp
bvlzMfv7z4p4Rb/WPIf2w9LgspYXC4KCmfQkuhE0bBZ7C4N6VDezf22WRPd0IoZKM6hM1lB8fAte
PGY57dipCqEUcs5jWc0MFsMbHhhl7dul2CRyKf3p4zUYEojL9HmYboRUKjvMAQmPstltOAj7PGw9
vbPwMLJKqlLwXPoyVQFHE2nAjVLAOD8xfs7S5t+OVww1B1cmrnRHnxpKUEGkR3WzGl7aXca34eEU
RscO0ilqQ5jDfWtut48FHkpvXK+G2qJmUPK+1wByiE+1PP6QUn4xo12azmRGb3kCH2F4Cjax2OzM
GiwV6JlLN8AbEFAIfkilDJJdHq1MatFcNLvy0s7/DqTnV1zA+6S/I/H9fIegYK5FSsPSrnJ9RorP
ppJniVUGurUTAmNWe5tvvQ0HbNmP2CuVSDh4Dc9DS378wNl2OLcDnaSZHaY8mobw9FWlG3gvMsrY
gnEUlepU2RNKgy2pBOnzWk6BY0hjNStt2/SbO8n5mr0Rc/q1qGiMJs+xU1OOl6dZr8uvOt5wQ/Dc
4KClAKVbVDyjtq65jW9CWDY9lWxlunkfL5eqi0aZCs6yCaneK4s62XjU2mpveUV88QYYsK1Qpb+Y
M1wKkYYpdXXLg39AkTQp33Ol+xxDSo7//IrWVs1MfxcRsRdbi5N9Mi1kzf1EDaOoMATDxAXrC2+J
Bw7SWr9elMBToqzXQ5gRU5gGyG78v2qFr5I0GoIE63cWqhIR7H/ybo9vnzLp54SCNGvXRr55Rv7a
2FjZ1Gdrfc+pqg0jf/PGCh/qMJFkgGpp3VTgLdfyWdPYb7q+jiwXPJgULqDpntj25kdKSmPiddLn
UsXQCv/9F8w4R4Cb/nAGaZFo7XZ5NvdzlFPViPDisOS9qoNPpg6Q5xyH0kE4jKXXfjJKnR3H69Rv
8e2J4WcqOmuA+hsiNibKGCdIURlcBvDpsqvkCnfNWb+G0DZTkJDZ5Fcb/t4NADFO3aVsx9UVhvOl
4rvROuJKhivt4GELIdv/MgUdMHdS8n1MuSl5iPb+F0laxMTUt37jle1vxX9uoPGuVEsYBUBSS5Wl
8XId1aYPHCEG0btcWblqudEXbmvV980AWidkg/tvtSri1a5TV09ObSlLTbf8ygdSFWuZ/Dhj3g8G
guqG+cVUHS7zUwrKEyjiaeeEvGbZ6TRfloC60VbsiTwYhIGg7O5LpZGOle0Ro1XaNZ2j8mvaqz5t
smS0trKTcjIF6qKFz8o+DqCM34TnEq7MIvQD872HceGbyetXgrh+yAJwgZzBoG2NJD2Ha0LXSQ8H
GrXyDKeNk/iY/Oxfz5EJ2ZouMQfaCPEth67RFOy74JGW77fzLq4V6TSpYECtS9cx7Rda4Ak7tdtZ
RFw0i/PBC3kY42osOEdaqH8xtnnVC+VuKIhnO+cJA+AmYuH1izBxw2VjkZVEjxUgv65HmFpneczA
9KN6/D7cLodKP6Ao0M3m4qFFDYk6GXY/7LvWjFa3aFfOYO5R54GPm02rj/F5H9pbFWmcyyCw2bBO
/h0usMl6BACrx2Bu3ACtCNn3Z2TMguKlgbwpXyddXBw1IkLc6jOI+169hXNz4wAfQFZ9BfB76SR/
MzNzJk5RFPU3gszncQrWQjbxP3xsXxzCz+ocA6K1544wysOcozANIgYHEyLygB4jEWs1yaT/RVF+
eDkQ9xLJRR/C0LaRy+pKBsJjJhz5X5PkQpSq2QVcwNUvz000Zqs+w5sUj5P517OTA6GGcIuSVe66
LV5SBTjLOWJZik+pF86B0XpBwlHZbkgqJ5zqtO9hRMORPeD3fu94S5iulWLu/qv62ZEbgrKwKhFs
aa1EUMyehfRr4gNRzkVInhFWweeUh2/Yg/K0p1H5cQp0uYxIqQOOYoLRnvDkNCtsUxmMeUH1GCS5
MBa09jA0/ASefQlLlMGqwjN7Oq4eBRLhFtlqPlzwd1a3I/6OxXKf8or+KrrolX1xjAXhCXLxtkFa
dPaji5GW5dbFht1tO/lSJUwmKVcNIA6DAL7KkorJIoCsqy6msKHbmyWxy6Gc7ht3iR1lBDJ2IyHG
YAJBNIE3EOUp1KiQ7zJTtMk2KDelh6O/ctS6Lk8ZuKd0nycM0EvoUYdjSLx+rgSrqzE8XEPYBb3H
NGI0p8A7hC8dsdR1AVdYub+tDoi64jN9m27CIZbgcmTmEc3dN3lzeS228S0KowSG1/N8ApjbkDMc
UAML97aw26TnWGbWZeACqXhfBn2v7lJzNdEvwDDokdx/lo3MJbMm0Hwj6Xcn2dGFHEM/4fbU+ENY
TSXFHlwNPcgTMEe4O4PRuz7oTPYHpSBWia1hSvvx/aZ6a11IQ89MKSGxREk2nQb3B5IxZlJa7A6E
yOCLUldIP8l+IlBGYIZJgLpkyj507uT5uq6IEGPeJJxKZn0mKCLZ31upgCmr2cngp+7kNKfXyDUx
7pCvP2p/naUfymcHis1LUWq1HnIWOpKOqW7JIqlexV5ULYn6e+OaI5L/+Adv9XRs4IJoa/0NFsnQ
yrkx2huPP4rrmLc9tfn9QeBluNJxB7/SAjGmXxkv5LUkKkYtQwnvGndV16dtk/9af3blj/rVvz03
LQkpY1fLTA5ZLbm8D4C2+gaJC4xr3MC/DDtQlN5HpWz5FRqTME0f26R/6CpY8cq8k8NWGFMmaztk
npjenASuJUNPrWBNYu2m5aBwyTjKE/ZUBneIL2iDUmnu1z92Bg09B8SWYjAN6uk0DxCql/vxCR2H
YKiMlTc1xmt1wYPhgNsDzNHvlP0GPWv3+uZYoQl2YADod03DyBfa66qX72bxeEjeNpNqVU3IdPNz
YnUyZwAzDiHjAcf0rHC8HgBm0FLypUWkTyQeyjfsluG8nPFaf60NBxzThFRiECqdK0az6Iget+AD
TeQ41DCVUnERF0Cy7fwRzizSB7ksIDGw9XOELVdltNh5kDpyjLqMTiFQ8fB+ZeUU9sHbmlTierpQ
0rfzakUygf+cOE2St4HYFnd2ZsmVeQ2ZIwtX4EEReXakctMVpOGfHI/sID/dk0sZp8xbyGpoyIG9
Bq1n3yy4X86NmsMuEG6qUB3cIXGlvhczjSJYyM45rkpTt0HTN88sa3Q5oiDBkKmwGB3WWN8Y8ABs
Ge6aieDl9q+0L6aNMtEyy1zlv1/XN2FybmAgNQ4j/vk/nYjPfUD4vP1NJ4AQhcxfFyFU5SCwXQHR
1kI2C+daUcd3aZtE41W7wVnqTA7wErKq61ExmSHbDZvyh8XqHGD8MjDM6Ionl44TvE44hr0PmoIh
pci7fSnF9u4/E7+hb0BjU+4MV9l5gpDDGpLmIcQJ8V9PX5owBNVQWyhsNq32SHyG2jXZ4ew9uOwC
wck6yV15I6azXfqhKOGQ4DghBckW2vp2oZ++mTFERNzW6/RbuXVbsub44PHeHUxD2KLP+Adq2vew
+HWmS6/umAZojyJAsSduvdli/W64daMsGKxPnFnyIryhz1yXmh5F5N5WFBAUFSEBTMnGWaezGXt8
3kV9FzHi/sB0lJb+43srGMeRR92yOuEftvHEBwRVd4erHVR+1n1C3xvywDzATbK0rfyrT6P3z9+2
LoPeW1kuktY753ltdyhBeC4owfKmofPGT+0u4ffei6zPP9R0VhvBPnyeBpZreRXZaC4NYjVlL3ah
KisLi09GKapvUIAI09hT4ifoesp71W4RNBk0etGIlDqCfr6SUjLCiXwHeuqmQ0eJk9Ry6n2Qff7y
K+ilKo7B/YEf8c8zxcQqrU1tcQKpqzGzDaZM7ahDCsP2+yOj/7xEy8G0LbVNKrxX8rVQfz9Nkzd1
H3ShZHyzQkCqKuLTFM5taxrnOkMfax+PZJlCw8JCjz2waM0fbbMKv1iyADUAwXz7jrgRqzh/l8Pa
DzdisR4JrbEXlgPohB+hhdnTIS6fHlxDBHczUzh8o05tOYuNqEtgMr79YAxNupEE/ySGx/MT+oG3
oAaE2oW464B+mJgvTct8YQdv5BGiNmekyb/gf1M9EWzjHaOGu/Fdgml9JG2yblQZHEikxIDqlmE3
Gf1nsaeQKZg8yfSCpnkkm6fi2GUtQ7y/3tqR7DZB6YP4L0FNvvuA4AP6ZdBR2jHm0N5sm0y9KbSO
raZg0BHv2SCeQedbPLm8jbG6+7YGX8aoZ8km+fXGkKf+EmeWaNd+XQ0b2uZTUBi+YGSJYPicAcsK
6mDImJ2lMbJskwy9DWUUnjecx+IbCkkLgnyGMYaM6fOjw6NyYSITgK3T09f8Nuc7kdsA6Z/z5Sz6
YO3yHBilasZFphyLKsmrWNQ250PIWK658hO2fgOVd1NGAAANX2ouaXo1l6FEH9NPM94KM0DD7LQ9
QVy4XDjP9eEWNr0b1JbBCSIy+L6/IwnUH+CEi8aBfgirx+nndg6+NCMHWF1pBARH2y4M0tWBBtuj
AQCgsHMF3TkVt6GC+qZKrEA96Sc5LHiADFcwGzSB37G/NzHQFNORDgelIXr7db8THudQWlYMSR6h
eUWIdr+eJAmkKc6CZK8qW0Cl15sHCu1jzUelAE9bIMl3guKN7FORPBHfvFYIxV+goQi97F7a1KGc
ZSFW2RIL/XKwW8JkH/8fD/NpL4ucTxaSmwWWEHt6ilZRYz/5e79AaIGkSZYPG1Ve4/8CMmpD/YNc
/AVYSrT+iDw2mIDQ0qvCpUL/OpFEjjSQUdbevwwrQCuV1e2OxyAPdUQhwm6ZEC54v5fG8Bcw/JxV
pp1inIHlNBKpWUKjOt9j8HXQdkiSePRJ9YIuoUW+I3XESMSzTOhyha2rhPySS85eIA31n+qXYsEm
BTbpQhEcQDsWf2QwnT+Z6hcJAITRcsEu5UwX+Eo60bROOXxTUHRx1L8AKuH0ZkhFZMcxtVMms61X
Cq3qD23bpusSqnFR5KTykU4pV0I4can8+ZE7EsOfdDIa5bKMTWc3k75X+n9wjgg403u68rIQbT4k
QQimvUVulz9ynjc9YOnJwZHuU6yAH2tEgAPBo+uaRBxc5hwrgsYVrVjQuTq+pSc8XjR2W8krvD/M
nPwQ3YXqwAw6yrZN8KP1ofp1C5xr5FDXy+MnziZZA+cD4WdveZUADSPs/lIJ641BbQqCYIWkcEJR
kyhaICYZZQSROpj8QsLq4myfaCy/vJBoD1aJKRuLwHsXLoWK4f0rsrLYRojvj3TCavAFl+tH0DcT
OnSae70xUOUrgAhKNF9dnipZoecan88u2azNnw0/k4xcyJLs0pyfktKOJuJ09qsy9RoSyQpK1hhD
h2C5bLp5W2jXnzqR+W5Zl253uCvGXZF6tSOBeg/lidaMWTz8mlHgfvA95dcvpD/YzdWXxWfBNU9F
3Vq9e1f6T7YMGYdPa+HM5/WSAkHk930JuGOroUCIOW7TFihrr9ZL/0k4k5Bk0QwfQxyp0lH3eqxS
MoozEIBgiuWpFfGLnn2pENzKyqfoZnyfp9C0V4BFE5E0EWn9Dntn4Gjf9ngfv0VFO7Nm/HYUmpn8
OEbIPjspLmLwUDB8dwB6Zdymq3oVqMX1YdkkcA4b+lza0srGFtWh3imkvFujBwAZZxlI0MKglQM3
XQhrYjNTdfW/ndMsMPUx9TUNWxbbacKdj4F3tOZ6wIEeLV8JZkkHgf9mN/KpvqSaCyQTt+EQt5bl
DraE9RqUjNEgqzRPkGL73vwCSAgej3Qn9y/vsfTELa6XgaIis2gX580IuXxRUC/ojPdbO6rwycYr
rz0oQmt3rN9nkqOy9rPE17uHTOgBGRSZOlGndXCD1hdKOG+2QlxK7IqgpFtDlHIKugp4Zo3vJyYo
NkG/NUV/RAjkqMGiPMEZCKtEffbEq1YAne+UZwqTufYXdRJmk2WDvbA+gmmFuilQpt2kTRIjg/6C
Hvk1TLeanvoY0buDgpDjwUUJVsWFrexoDwlaQiPb2abN5S5vdTfOrc156HL/7CZrBl4R1EQhyY9C
4SUeRCd38rbQQ+jJNO04ZeRaBaJxjRwZadOW7vwrnuIvQJhBCrNeVZOjaAnPqAtRJ2e9VTLhlgYP
lT33Xe9qUSlpAvuSBRydZ0KM0/xA3sau/2ai4xrlXhVyv7KBd57L6eHjflLRmFWCMggZR5XeTzrj
Yo3rUWUI+LdPs3g8q8/2SYu+4odtPqSokfxJwIIUUYBsI6GhHzkXtPn2DFwnkEAIiz2rI6Ievv5t
mgj1i0NLjk7QW70CaH2rqBGWxBeLA3Ijdd0x7w10/KSgrv07Rm4ghfCC17anBmPvgh11VJ8lKaDs
FtQprGNLXgJ6JiDLXlRsj6mHK1ByJ367K60y1KvtNV0QnvWse/85m0vVLkKNZ+Xdl/C6XQS87+Md
DJz+GgW0XovsTxYQusMcaOHld3FjZsAheKveR1qNfFrXJmaw4acQOhVd4ZCRPOZRBpYhx8sTbK/W
+2XQvT4rNE0RgVSaTIlp3iOuYQTG+W7Nlii9aBXt+yWlcp8EPddcnhBaR2c0rXQck/1tZNxjQlGZ
ihgC8fmsD6WiBu0XkjuYy3r2uUfJHc95jy7utWXfnXfEW/mK+WzoQbgoxRt9OGcAg9a0EfKWA5nR
KFsWVp+lslwxuAW5sUWbkuUpdVpcShjHPBFlxKrM20nJa5J9lT27U/8q4pet+vqu8TuAR7f0UgEx
VK8+9f7WKHfjqFZ9dUmm34+bBsYhTgdfk+DXMkEunxHIvsjn4Et33cVkQb3apQx1MhXo+AvsKL9N
Xc39LhUqNgwYKhyAQQ+3fGg4eujnswL8pi9BH4IBKgK2NTF0h/69sty/XlkTz7Kugf/DwRIdZooZ
Z0WNRGwcTAtqZsI5y3hROwrmVazse3YnnK7slzAhndWkanqqQQNLisAo9x9OOZYxR9DVc/rlruLD
0ZiQX1LJQKVbSGehe/TaPV5X3HjcVx64QTWQQ5gCOM9BUme19sjfPHEqdTNstjoHD9/Y55hPIj9b
g9k1DUp4f+eAgbrIrNezhr5eN5USV7qrlb9KyoeezluNWEQ21RZ5Pl5eW2tLifr23B6n980zom3y
QIwxFYhu2GY+e8BX2u1Chw2z3LU7Hgh9q4by1uwQdR0TL41IImdQ5wop/nSfsEXiQbTfi4p9/i45
xT1toDOyY/1K9nR410f5eg/wEU9EaatWyg8BVALL9X1AdftF0hvfn2CSo6BWIr3bC13cd8fCt0rG
n7br6Y0bRdAc/jcYrrod5henm/ElCWUQadCMP2vuO5TXpeIq9IBP6jPfLI972KYJ/N1+2BVg22Lc
cNAcxQwjlTvrR75V07Yk7aNWYYrFT5Ugf66gwCC46RYyht9c7IHi/bbBKNv8BFsd9PQkB7ENjhQZ
XvyBCYFkgNdcdSS0E5kdCMRtSN79Bdp8AmZgVk1dF6istMPB21fBlFRzDnRKCjdysTHo5pzGXFRP
JC1ZK62ypHSpKmXWf5ihjALrgaLR2CCEklVCtHpyf3yFqLXLBRqTn5MKn01PSIu15iIQxsXOccSl
RV4RKUejAWYx0Ues3IY6sHBCtDmEcIH05eMO9iKFcy+IIBVMXMNwx6YJIzNgxtA3uWhv4g6Ld9GV
H92BZsqyRGVZoN8+4a8SVDbCdaAPM7TTz3nhPZM7b4GKDxEKHbplizj8Y5PIBqmcp8PWlEE2NIk2
GBi/75qg5Wku28fcRIT25n5Jbgf9EFvKmU2+NzGvxe7Ly3KN9xodYfdDgvXITGLllQEprUTkM598
c0Son2NxDghArL2p0v1rumMBqWxBKwb/9HsH+nK3jqGYnstgkmoFO4mX1hF8Xulk/hhl1DcUvScs
n03Eiu7Sun3Ay6/0ox1fSjnRfPgJDgi1pCSAhiKxJASNsN5zDucl6imFG/qqOQtbUtseGVGunx8l
un71KnJ2qwBRkCcBgYfM5VRq+T29ml6jm8fbxpOpuZjlWYF+muACx1C/qeKnfXFdlS8sAgU8TKCk
web5i3bg50oUcEVJh205QIoa5Uk/dvaSrfwgW8VFXPsFcTBbBBOm2+5iSYAomkE2fgzmVRZDxlaU
jpnEmWa6Ya+vHmq+24ujncyd5SW4T5Fe1Pv5sTNofDiSIfy6Wx/FfViW9Zox+2PYQzt/gEiZLP35
52bkv26uvCY/Izfazwx93BtHImu7a/qV5PNIMMeHjmII4nrSt0+SytNYZyFktPNRUpu75TCkX2rg
AJe5g5ST8Dz6KayWC0P9U3tTUsIURtzDqWiLySC7lY5mQ59jR3T+XSwIRE8KMhUbCGVUteG9rm5v
+z4THd+poEYkfCclnwoKNB3K52Z9PBImcsHmpq2fn87yyapgA2qsQf0uRv0fDB+5CoJZG2/GPJeK
zH0Kf7RUhgCWO/67qDLwtaCSVP516q4wHDgv7HwL9cf4Urly9aUYWRxVuWwmf0WLOApDPj0I2jcW
lzmOidqqkFj5BCfXG3akd5tyi465c9s6eH2U6Y9etZwhR+iDnb1rNdb9dsZ3MV6iu4L/TNosDABe
5eNzRFkcTQuzQJ1aMYgWeuq+Tpz0jV37WAEKCt+PUTtNRCcapBbKFDhewdiE7H3o6R6o5MwtWYIy
XuIzX9jHoCwnbGFW9yUiMVxUPF5R757G6IwyUP+gwW86L2fUZp6MpPcx+d7iVZo9kH/54yfatCUc
7jtV7xT4qs2uHRN1BmLjphyVsKzu8khJYvj4b309E06lp6khPv5WQYScu1eKh2eX5c+4H8W8wrYu
NQxbZ76GwExkxrkWcTOoDbsdAmODzjal3C6p3vOgPE72RLp4WfENxXl/nEvs7Oa0PngwQhI/o5hn
2wA7fav4AGWReJvc6BIxhwhyLsJP1PZxAbswYJqsnTBOojhpyWfq7tfACEHCCLghxBrvxXjmmjv9
tJ8uIV3VsHEC2R8nAex8maaMKRpMxmeNNa8OCv355as9pkC4wcZ+mRN1fW735rbrzGfUyh+1HACx
0kpM5B16pMUyggboymYVRvxROLYft4xeL0ItOtmS3Uw+Cb9EM+JDLumSGguQI5pe/9+286IbOxFO
Mr/izoO6Ft8h+nhOoxtgpHGpFwAn6MB2G0AfN3+jRgbAKNy6OfZNoBazFyuNmtM5nLXLtiBPJa4B
wn6vzcxp+KOgH3ZiUf39YtHKXia+fQhmdcDYUUTHiGXwHYSCSE0t93PHQWUbx9UcIkcGOESn/aUl
Fn8UxJDVJ3Zjg5NMmkA8gk3z+MXqc1/jg1O+aCmvgWQV9WC1vcR7ZFQVoWNcKAwNTmImGC/mzjbW
VQ52zLe2fX84nqt3BjMntiHccQC1/LfObhSa/PW1/cGlHdDYUrqDtzHbmG/omfOldZRJ4mMDFTsw
FENlM1e7z57BBW6LHmjQ7/bIfpggaZVoH1+A6IYr3kRLzzMgndD8PJ0lD4Qiud+/wNoy0aHxbWTm
HNHFi98ENYhtcr2ij77W+PynMfYevi9YSgPs3d98tUH51sP/6EBFkcSesLE0lkN/S3EHPWS8ruy/
WP2ayAtudzIi/7b3D9Sq9SNCQVC01SaEctExjP7Y2mRAwiCiXCMNE9MWnGI6hFIIZH7E1+SJoKYM
wMs+t50QDwlX0Sn/2NaUuHqmZU5RBxk+j6knLKNtOxLK2Na/wkPnDjEiGJodJtvxyPeoqWa4YJNq
ha50R9wILGIUbM4q3siXhSjmV9LQkRjkKaWeQ8SiYao2Ay8FXvVZ4zkQzhYHcuRZH95f8BnBfTc4
NrJqzj5aNUWFN9jhdmld5CZYzNR9nE0m3IhpOMsshAhlmHN/i1i9feB8eHyOoP6zkovW4Zc3zIkK
5lNEPcNQjoqjnnjMcDI7p4E9neqbbFA5V082kUjoQHfSi14wkQEJORVWQ+ZU/ipAnNFTOk2UB56b
GWDWvlfrgiPvbM2+wdrRHhwFUJDF8DNGMT8ShTScl67UFimXuu1nGtmR9oo5FEoH4rx0Njirha7c
1KPULtkrCz9q+/ntUyGksR95+mWXNypOGA4PBn6c7pW6U6gj+N39acHqDMx2numQQPMgWuNrZk7F
A9fljK8cMcgK8Hx6wVU2t2LGjvNboe6+4FerWIRL7YQq0cA6z74PmXF1zub7LQLB6uaDl2J6izkQ
fDwYTyP3bLJt8P9A0HOMGehyq+iqeaxPRD5BTKEl7wkvEqJWkEe9DJiqzopQdD5TbQ9di0Q6XzAX
KdykjBpBrbcff7aUvWN9BgJKg5Ko+ucfe0bLdlGvqKcpEGPHdrlEGTvYeDoG1PsrnriD66mCBIWD
MyEXK2y9ytcb+th94VN9Vfbl4paA3MTi7HJLMj7pB+tI+VSnkl5Wavu4tFenoWhwvVXfU4TbikKC
idv55MwxI9pgUzWEgarKifpxNK736+VazDwnAJ4JDoy9j/Bx0GpiTuuyAZs5U7UkdvtDIiDFSYnw
OBKgCweN+7nPFD4K53WPO3SglVq833iEK0nUiuZ4v0b3ivG/hWmVFFmDDpn6Xr5qQ6t/zmFxeCKn
jSWwGUEJ9S5aStdYJB6dU3DGsArkrMDGSNTUfCR7lEZ7EegZBf2f80ULXFmclVHXM6d5+iOoq534
3awxYgV055LV12FoNQOlLKm8yeB+pAHGlQ8i6+LJgnuTWJg0TdiZmfi9cDJ5OmW9WCAyf64KF+rY
2xUrb7tpAl+Fd+UO1aZOY4/ZFjQE+ZEq9533AkGUHtl1WW1VfTUFun+67/ASXJEVYSJ1eWFEuwQW
OGYmokY9vDBK5Pqb7DNfSXUAhfd11U05P0gKh3oDB6e6PuGR3GWvHHQmH+EF2WCvCpgqrnKTY5bk
UmA5aIvmycaIhQCI7yJgaSFburp6Ec7nRNy9UMHzJQ9aVxFj+TsIsE8bxsFluW+SPk2HmH0TDfNY
a/uJlKXyfDrMVkaNU5ajd9RTjYgpd0WzJrrlPtkOYrkk8GbZyTD9uXIqgPaMB9jucjjB7romazFD
TqwzsGpbV3KPlRz4OR08IATQmA4dgYyF9bOZbzvbuQohr3EMoK97bXVWlIwKUBM6fVqtvlVJ1oJ1
ViQ7s8J/C2n87l24VLBAYTW3UIdNJjAr0dDHrPbi7bXcN6GsytsVjTC2ch16EbQSsszcwSK1Uy4/
Oc6MA9LwdyGXppJ+sbkjaYcmuUMgeJJxFA33xmhJqYafImtN8kM8/Dtv3rTDnaIUkTBtaWcLiOmu
Gxqqv69cMwjCuAQoCJp6CkKrl8VEDBHFjTUU/U5V7dqc26X6jeFfWkgbtdJpSoRcTEN0bqOGgR4O
Z7mL7D4qCioIuLA7GsR3MlMjgAztP8Jo5M7ClChZnuj/Q/PDTZ1hmEF4FKAjcBcKH3LbFobSDc5x
XZdc722YODbfEuiuWppABmSNGCbBCbniK6ndxRGPZRL6y98u+pELlg5sXoX3lnvirw/u6UMykYU0
URCGUmFr2B4eZBOML2zLKuGbKOvDrEqHV4RHKycwPPg7ogP8m2CU9GcYfLoxpZqCHI8WojeZ/h3D
qsWFoHdBBWwvnIeusz98wVJDHYMCUviohaXm8n6d9pjY5DsADTyBxxIk60oUqyxGL6Q9y5COcUZn
KHYpZ3bRNRDYhIHDXnZrlBwACiJxXPnkFOCOrI56KZlaf3p0lqkSXqPEVoiLUxRNxt4zdfElns+Y
asPYAXZ3g7VLyG32wOpFdQYv9ZTQ6zmXjwQfikKHx2nTzjFGtSVHAOWG6mp5krHO5dWbITl61D+m
TGHz8oNKTwDtH18rVX0qkaBW5Hx6Gm+7dn75vXoUTiaGiQsTQrptLK76uNFqHITcHT5nUsVMCgj0
VfLkwj7Yr/TAXdFMhnZXdn4pLEPAGvwihtx5KUK7Yojkx0KHH56wxALYSAoMe4CkvYL7A0DDW/hI
LJRFRf5t7o/NOxB8pBj+sljN9Z3wSkzNoMQnKrwSMwHCACBxrqW8Lk7u7aG/vE8tWJhKuhZETnOq
TKjojzbNcLGWd3HAVoHzzbecjYV/wwBAjScxOZi/kZlyeLWfPwlsYOJdKL0xYHgUnMKqRtPjH5EW
g6k7W4NqlTzLP5tHTQemOlzBZhSLscdcSEnKi1+a8S52YvU1eXbP+8V7t6O5vvLZ2J7Hfqnj6ony
82/wuPADsMnc4UoDxnfSeEu+BxBHvcMsY05uwAfVYpHfk6aiCy/fRHhxoSmFfZDQQpsgnfC86UAP
akcJ9BbV0TXyhjgtVKlnGFbih62aZD42Y6up2DzvspwbjMqCpBeMDjPvpcdU1GfyPcq0s6dSDpIl
ZORFJTYyTUq3/X0t3pZ5jpa1UrjLqELwu/0WDM03XJ8DkMjqVyljWk+fIUib/pRxB9qAEJcw4A2A
TFNJDNE+Hv2uUwt6QObFeA/TFpMkprTA3kFcyDnfL1JiODZHITHuISvJJiMGcSmPZo9wkT0uI6tz
Wy9HKyVI92dQi/oQarVDncvN48E9/JcztScz9b/bdBj9nh0uyrCQRzsTiM6z/8qytOZNPpzxOmf7
I7fEAj57W1XIQSquaCqp+PIpMisBMylxpcRSokcNnjFZYb370Z2/83IRgbbMRdZxd79iYE4ykGeF
W5dqw0mjAEpVxhpd1+plT8VUJdimIdtkiwvcncZJXNlhFGsfmMjlYLvVjR5yrhq5dayQPevQKIRi
cYC4IHl0saS+eDjjccbxh1XIy6ZFgMgcHfHF815QNSwa3POUyhvknALkwQMyIW5kAMcy1gOP+NJF
jqxA2IxKIFYgRMSdEvpNdes2BTK2eRJgnb5muWlv1T8U/sPLzMsPx7WiisSStwBqdyPu9XE2MU8t
CvRIe3/AVp35EdKuEJnffVXXudRDNNpO0qdNQD5vvrPXpWqOD9RMur9upFjU/xTMpePkVTV3PjZ5
GRU84l68S2+celbNJEoFcg3bQaD48ee32T/oVo/aS6FcHDjSBTgHEjU8oHNXSgQ/00IopmYNss3u
9abnntdlLvHklxHiZvKaAXIObuYzTZH0Kp7TtohHsRRH2s/29df6DQoOxfl9TMa77Ia6IAVDGXyB
ZZ4isW3c8z1mP/WnpfTU5OKEH+PN8Ha2PG5TA4EkzeUcGabpbWZUMwo0jNASwaV2neU4Ln9ORnpg
+8PKk0mSqNsVm8nZHiQJfs0dP1qYZv2GaBbgFxFIvlFDtBRNz/lR1WmwtkijBoDtLZL8B1yvsFBP
iy22pp1Uj6q14Xsvu0irUFNrw/i44RmH9tpn706Zhs31fHM3pT6YMQyDdjqZWqhE9pgHPRnTK8S7
imEqzUuEgXvKxCoMk5PaK9dOrYC4kIvlWsmlqSerwOnVyS4rfeaVSMYfF1rEQgkY/G5zqy9HViOD
iRzniinMChYntOhDYgJXsNgicdgC8tDkuFQu0HFnnnw2jOLbw6ml2uC5lJnDB02kwhW5XXAtUn/s
qxojUe2fqYiCHfDJvlPn6GoGTRB1A6s+Pn6fjxps1UywTGXHyEZopwWRhLUshowxqmOCEMeqtbxm
jhLbqVg+PXQLjHnq7TYiiyLKaX4uNQEtiDbQTibskvn287bQC3q0PgrByVw30pCN6403BJRO4izi
+PyvLF/zHQgrGMoMo0AkfE2PiVdmztTmNVA/KmTYtQ0uveZfDI5VHeTAr31mcX4y1LpX+xWqzhpZ
fNqeNPWirL9dvC6F5gF/tpeFkK8ysNDTkq8HW6/PrgpYNaerdFgivItjNMRPFyPsqlCoU7F4Njgm
XeZ8+P5D+S1UpAG2+oZDGsh3ixNP5+SuvZMOY4X5AEp26eVf2h+WNdumhIWEw9YikD5p+oxvk8vf
Ql34JYNC1LC3iUmeJB3mZ/Qt0wchuXNzdnULD8fCybfLOes9r1O6/4K1F3Yhzqi4tEr3B6KDjIyH
i3p9s4TgfsI7WlNmwYp/pdGSWlj5ym9OtqrwB4WcKC0fhlA/VhIDTYs+EkS/mUSu3R0L9sXw+W+z
8+9jzMftBLvPpRp6Fnnensl5BbwgAu/v6Sk8/rWWJB/LycBcXKygiVsZzHYHqu/B6xzfOXCRxQsp
KlxQ+1x6JPIrUZKmoEVkD2iB70zhJbtWyv3xKGUDF6hdHChtIPlve8Xj7WBUXrz6lba7GnlABCRk
YhpIWI23oTY89WcEu2ZNnXrfjtANYTgUURXNWg7f2QCJsdkD7vStGmmXaPBFV2CeM2PqOUM4kbab
+zEoFyR6Nf0Q4D0r1WCWkKdXf4Eylc0qrRm7kFuuCRF6lOAXfdr+64oE8btNQy30PqglMek4FOXr
/eorP15Dq8IA7xYwX/IwW3VPzEcrIxhHzwDp4EZ6xp/RwQKKT4PzPiYEK45+QX3OnqE+pmBbrwpo
pBRPLWEN32HCVv1F3h49QnfFmbagGye6dQneJjSaINLUYEhl/QbRXdqvsjoZGR84mGnJM7S4P5/n
Nm7bbvOwMlJe1+vP9zDCTBPu5cMLPubwJ7OpUwdqLA/z+dZx8WvGXvi0KCoEfK3OxjY6/BRdPBXM
307zB5/9lMbVAv/bRHZ6uv8VmeGtw1Sky+vEZyxUG8CJHHDcHgOoA0pKXszXmQSTpzEZAmv2vyoR
EJ2ed2Smi4gzPhopax0dC1lBjPkZizGCikLDZRfedUWIxt7OpP1bU4xqSR/7UlSRSyzhADLmx/PT
9uxiQzqj0Qf41TVADmKFXTVxHWKOI7fF6Twx2cCJbage28nDZ/QgMkbe2UPa5jouTaB9ZbLs9Yh3
KSUd51vRZGPpl9jcML+BVQxL4t7P5zpe8YD9rlKlq74QuVcW/cu/v7GzlNG9qWa7N+8JjAZm+meX
puVqS6vyhAXsNvjwFSGsnE2aXpdIYBrXYn//orwsSjnsLB2Zj3GUlSpQagjHjVILad1FEemxjyDc
8KLYI7myg1YUahlzM3oQCRZDHQYxs3ECOIIXk9FDX+rfnMYzzSrHNHO/HV5wDDDM7w3kl1VX98xR
blE+reZE/Ao71+eefsxU93nNSCPXjWlk7Zz6u56EfdNvbNdZ8+7kpO1pZyN8ur5whBQWu/O50VBI
bGJMl1UK1oa0hki0c+N7TVncz3n9DVznInY7Ok/2DjYuJHWCZ9TSbW9aLbWRVvFWZCluQBbiX4xc
6GCQEJj0kP0X25hBL95wQkE2hyD1kes1RyaKlqR64J3G/2F7xL9H9VjGz4O9uHYAH2IEb1+kV9A0
zE0z5vhAPnDvOb8PefrORXUVXD/zTVR3+vCamlLBf7GTovwmbsKMhplXdl1fUMqW7jXTBInRxHU+
wvCvtIrtjoBPnKd8+KzVlbrhx89CV6fknh8teNUwxJu53OJQEii8ahlclIytj9Q+Ef01sKAYX0PU
0B9f51sHT+mo+9sCHcWO2N9kRT5X6mqasFXnGE4AtJlvB/oIoWmWPr7/PMoM4cSjtS7JpwwbOFD1
rnumHd8D++cyANFA/xNaZ1HCzyG3zJaZwAODVgF1SouEqnevUkwMu7Yq83WTRXgt9u5ISdpRiErT
YFsEb0gmpKbkIgECD0D7NAiBt1fAC12SMC3oZtmxCwXMGa6LCnP8me4EtSORLBqMOhV1z15lHlyg
ACcc6KGdI0wX07KNNBqeMUygs49/SAiaL52M87WrPl+s7rYLqLxGrrM5nnyyfgxwX6uD4u6tRHca
L944LAwZp6nB2ETLMgx9rv/M5ZKlYLhYDUHMaQ61pZK6JOBXKWaqL50sHsxDNkIQ4NnRUOd3utqV
t6ELJVn61b713x/TpIzumsYy3BNR+tX/dZIyBvzbeUMLSAVGizsLiUzXT0rk5SzBSl0FwxvdpMob
9hUN6kW2d+sbq7ChVL9c9ttZ0LU9eNI+ajn0S08RJ6jhJsfdbTWtLtWb43IOXDw7NK284C1Iqb44
pScs4aMo1mmW7QVyT6S+9J7Dkpf0KN+Q3YQ0iWjHzZ8HIugDYltTemof+w5HqsK4dgcSZ/B5I0Kp
o1MTrTT0MqqFr1q94vw5VMCdpogQhKqKz0jnlawQCpYzUBpoH4QKUa0FkWLGdskoOrrmLu4PbVq0
oBdBaVdtLlW68Uepyxv8Wj4T1MvC1/6HZSWYF+8XFWKMrtQO2Hj+n7fcd0+7+l2PJGpwu0JJHvGk
iAI0hyxe543AVw84G6fkvTQjVgEzMjqPboZvl05ExqMWZu9ruM2mVehlif4jPDhEpjPiTGOcXEks
JqDMYJ3LEaTg+B1EDc509N5YZt9qzbDDm5HisA1NIQ4Cnj5RcfPtt6WjQjZOhefH2ZEgAPlKEJNh
Fl7Y1X4vcmXiqBoWFyVFlTdIif5jAY2IQ0pOn/gdxF+O3enHoxwWyexSMiEyCk0hoiwiaJ9lPfZY
ltNi8SeLRUS70KzKZ/ihDsZYraiQdcEO/mQ3Gpia7khYX8YytE4AgtuE8zxQzt9i7pRShoqeLUj8
5ii2ryEPeFhJuNQx8vGM1XHEOSxbAf1J9Ix0hxfKds7Sjv5rDwO3iwrFRIcHkq+sIRGPStuWpU2F
sG9v9fCn9m4byNKftqMl17cqZSj/qE4znt8Dghm7y3sNP+fh2YUm2P9Mdqchu7oc1dvNSIuEpQYY
gFWJvgGISVRWP85q7/fk7q7TUxRRVTz6v2W21cMMWbCSSsBs7Xghv7YzOpoypOGrqTSy53FT1DwI
ibdupKrGo4B8ndTcYNwBekxJUCjHP860LLkrbBcnlAJSlP+vwqWICUweLLvqAhE3SduZGpTG+cGo
gyrtz/4Drx6mgbUp/Ld0AYkOyDfWe/vAwC4m04OpHE7+OHewIVu/zgEN/wWINRUrSn6hZDDSFaL8
3/4i8bq+b9nX9surakmsQ/XlfftgenwzzUL8maCfPCvo6vqt0tGag+VdS89bjb/dKzZt23FBp/tR
CJVuo+aRjzsa1XFI1AbTk0qL5+i8j/q29GKmZnvT4jKtLgn8X/vXxDLq6Gr4ztOykn8QcnTACzb0
83ZKYH1LNOnlZW47gRPSKS2Go5ss4kABMd/xaieTx8T8NZg2ByWDvyZBebwWF4fFFMiujSW7lzOU
epK/Yr1/UdrADI5FOHmwG96ZW7j3UWKf1PqhNeX/O5JMZtXVir/4NHpZL3569R24oiRlp3C8MC00
Eb9hOusIhvCGyJaNI20ckFNG4R9DMmIViaCqlRkkoi6NMciZhhJgdcmJCbdSHxEqQp2o0zrfwmku
e5DZAFTbCFdSHjYHFt9i7PIoHPpGxPZCOPW3ayQCo66txQtgNza6KWdJFsVAxBIpWYGjLBh0GLAM
K7vvsA/Nbb2LvJFr8ED1Jk8bE/PLPazFJrANyFCQkcdgFsKyyiWGl1o8LUxjMbzobQYNTa/3FIM/
uIhSM/uoB2rfooOO1xqPQZmt+RS+QCkYHOz6H3XksQMT92fPyTG+iLVTMSUFKq4hfxChuvdiDjaR
vWeh1BGq5Z77JXgowKH/lJSyntaAUBfXFrqr9fBKN4H+vOyeSvdjMjLABm3Gzz+BGPlMrwMnDq/H
R6W7B5fPxAhe5FyXDB1jVIF1/7y2aO7qDh9aKw5IOFCe1vvt+Pw9szmy8I3XHhluNZ973MpZC3vT
SJYscIxLx6c2UFBPA4+7WcXQ4nKHNkvjtqmWZ4Yfm82NqR0w8SQn7PB6x9TQ5gVTu377AEpaeHXW
nHt9mkTc/EQpAgmyQG41LwogfcNr68rvdgW1+5Te9pUs6Yd5+mBAPt9PBMFyenptdvXD5bB8yKWK
Nz4f7yEqM5N1ZmrZDhgDM8IOjpVdVb5Ld5x1eohr+wW4RoV0b8fixKfaolw8ambFDQ8QOpBoR29O
ihrfyHcDFn6VQ3B1tSLpm16kqwVkYdsx48s0L0Sb/YlkgDM+OCWPf1aw8wMvqSxerem6A1o5qFr4
o7qGgBiGRrryJqX0ZqS1k34c3doHseR0AnSJ4/abK7g4karZJgbRMHcajKyA5Qn9T3ZUBmlYBffn
jTHjXM3IF5af+c0vxaQGGi6GGSIxnVRta6rTDqf0QTCJA1zHciwkGC8SeGPOUzHEB6Qo5crQA7Dv
jcnA+U/VeZx7PznOfCTE6VTz8MXnd6Vjy+zpq5p69Z9b0u87/rFdB2pZLOW+1a/grVDXVLMcvlHB
OWyUZtIOYDpyHGihmPGS7NQA5qfR7BGT7s506VgxoyjDxInrkwA3Dn6H8EFZE9+0ot3aQvVZza8t
sPsE276o1IqDxPuia/7DNQ9Sz5pQJGkeIfAgh+jXTvvOA4aeahAfgfKz/4/9NzNMJVWMa8xupJ5v
KKMLtGTUnWzgbj8tVUpMjaT+B9dm5jvrxCI+tT9n0lMNTDLRfTRUmnzRmz5S2csgQz34W8+WiqN7
SsYPh9nfXR2lrhaURozBqTKk1VZiaJULjtmHHWBD0b1QDY7qiJ6S9PDQ/8BYRE6TqmfvfeyilkSW
eREYea0GDIYAdwVjNCkq/rDgOd6XWNCpSLOa7jOgFqERUkDIcoYCjFLkXsM0dnQkQfQyHgwHK0cf
swE7GH9twG2Id98goOi6evT+3Z02vyvPhacVDGcOMrd4A2s7pLyT280X4i5Zv8SXyxR+fkFRsqkQ
yGy2dojD8JMC8nO4T5uAnM9lz7hqZWbNRp/lCQ3cxZ9Mq2Dblzn3uov1WX/DKQsDYI3mApqIJLcH
yKhvxVue5kWNafjrUsmp4xZ3MRjSNCgSgWvwoRSyeXD/xvFAE4TbY9gNMnK97s3jfCcNBRu2YERr
WDsxVFI+B5WyUTy3lJadxTMBD4M11wSIU1SxXOKC/dkVM8ISK1P5xj/+ueOMQlEIm0aw1Y2iJbvp
QhqGnNJ3FR7v/Llerc4C6ueihlnX7HFC6R+8/tEBqQJLnnuFfRXKhuhVgLNQH34oFno0sHTPzq34
hDBBPwl1EzRDWCCcvVdYMfWThA9oTYmqrRbRaCdF1hkQiV4N/qr+gMvAVvUfKulD/jvfmCWGW2Jd
FYYeGnfhoJffsYOVFuLUDl8OPki7+njOM307VK0Yh4QOC314mopPyW+l852lVltFG17QmXZi6oxI
BDVvop5QhWliXLIisj0P/ooYUvlugxmsD34HfJecESsc2oguEUufwvk+F+wm3Dj/kypLBa+vyKga
2pNOhSJtczIofvl9Xh3DZrGIFucoLCJ7uSc/HfIKNxi625ypX+DX0+shxxi04R81HIgFhHhsBae5
Qs7smmTuB9dzamngpf9k4UcmpFMlKy04viAliJVZSPCaHMUSLH7TFDswyHHTZXCdp7R0oV+9q4ym
whFwkFb84RTxJBgiBdTjPJZv/j/I02Ojv30gNIheMybZKyedYhLDVnQegs8E5oUYQSpwd++kFfju
s/56vX/JZgeMF+sI9vZZois2jo5gjlLw1X8h+tHFg/Zy8m0vMZikdg7EGwpisyHwCefuZiUbyjHH
YVNX3Xt2BSQ8nWGomr049OK4FwCrMlsRUhX68G0IWd6OU4JHUn3nw5qRQknf1kBB5Acgq4jF34jr
pl7x7BkkOesoSR9f/5tkRWHdmnpvnWqsqpAbFfJ/7mClCsuDO/bIVDRPHCIVCFpcYgOUTOiRAI6w
JsZpjGfDqVccGz5ihKOzQxDZ3oa3xDSIuRPxfz0pCaOANXPQOks9OjBNWnhh17jBq3JJhUKC1eP/
heK8dhLmvNLbVpL+9+S0TvMGO6d6itMjI1pOBCIaUoNRpQyB9PmUvZHmxdVQymmtu0RqIIOUO0cn
TlizaAz5AS9GcAacdMxM3VLX1Wf4H7Bk0GI8Ed0NF28Jt5+t/5vCIoHjKDVVW20uqGtLcx0LyB3X
wcj4HYDWetxLILINm9zwr4VPAb29nrqNTdLAlpNF0O0Hhjx2KznzX8TbVQ6nqMNvXy0HCfsMDbFJ
GwEx/vPX4Vu3+PXWoi3K5wTDu8uRWHtko2j/5ddk3aAp8c8HnJsOrp6jwayWpHUs/E84LjiVLxZ6
l8xusaWTfucc7DrVutJhCR82XGug6NEqpS6KOypgmmZMORCGyETHCwCdJoEfH9KckK8X0mRNPqiy
8T/Ortw9W8822+nj6UzrzO4ndahf7wRWfJCksUeATv3EmBtQAVSQVEc+OiLeUluL7ruTsJKb10yQ
cum29saBLz7xZpqXKtPoSuXEb4GFcKh7ZQRuJB3A1Mwesaxs7JTTevGvAvVhlCDa2Rb3fBIBCZJF
dRdL0VPRiYiPAK8GG1J0s6Z8GCDl1MUzJgHUKEAy+AiWWS+nJGNhFZnJx6F1z+nU2q0rukKc2u00
amPGVnAj1ErVS7SuGne3GgNcw0QO//BBxa2BxtF5nr/fF6erBfkU7GREbyh+0oJCRkC5asZt0fA4
0TcNnGUgDdeUwwyx6xtByh+VOX0n6s2RkDmyUgA+UExC5fiWB387AOQfQvEMi4Tc3l9iJZZCOEz5
0G2wsVbErF+kApqM8XkPPmOg8zu+V5arOIISVb2VyrbLBdH5awr02LVY2nm9HaeMsny7U2osaWE1
gwHUeIFfBoqR5dzRCHZdrOiNS2sxaJr71mLZs4Gbi0zNJDtkqzAQnLcN/KQECC/vJVK67RXEZLCS
PiYid6Iavw==
`pragma protect end_protected

// 
