`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15440)
`pragma protect data_block
giGA109OWTgnmloyaK8oODsiRC9RZVQFcgf9mR/obyjke8kkfwHUD0rFD2w6Qg5sKJtvAY8b/b0q
V+Sa+ZX24LFU4BuS1vxLWFGohu1WaQVSB9HQcsOWHML849yQr1UuXHS1H7VUn17v0E61+/PqUzk1
X19/pJmyYW1BM5ZHOhJulHdCd99vhdUA5znwgIeL+qkiU0sf11eCHljau90FYmDoD5m6woWzKvoP
6gHK4sfqQrITuaqk25AtWPgKwR1csWbXynMZjHngIasrLf7+jwQp9U7hvKe3TkF5y1hwawHe+qXI
mHMa1yWWpzfy5p5ieVb29m9XmYhrRxDyTlNv4ymQLieSHlFh4bpHz2cCPnZBGMhJ36Gsg1sx7rAD
IPLxwR70F1L3FPukc6qZVsL1+vSLvYcQkrjUBuN2hLvb4bJfdV4RkHev9LiOl7Z3dL9/ccfJmHPJ
oIeOItxDDVeonISQwlFt+bQ5ajDhE9yjmuAFvBLF+0HT3zG+SUav+xt2udkrBDevJO8lQDulHoCf
pMgN0AglRkl1o6Re1ta0PBnOxk/rErpTXrvgGFq+J2EYlQQRVcmSCvaHXeas8H9B+ZMOsx//OECw
8ZfQKprBUvE46tZbjxgKUMb72oOw4Gd496U87F3oxxIzLqviCOfT4OWvUes9N/PZ47WC5iZm6Feg
iZNnSNiqWdQ9qeaFXUn1QG3CiBq+6r+j1agJR/UNO2xb9PcFj/0nDVrYobjh0DzvxgLC4RN11lpF
5gLzIARh146tM+JNfzGjYOR4oD6QNU+73/C2+43vdA/8KEDa0HL+19Ht3xQEMR6Z7uMpqrStQafd
RhyF7G+4A85I3DnM8rlZ4Cl7lVC4DKvFeczgHaaCK/DMICJ4XLkuRTS32KrPec+cDy7E5tPigZ1b
Ss8fxKAxVpQhcNQWwzjdZQh/uOupsyjOBUhj6Hq+e2q3i9qIdMNqf9Cme2tWbT0GicHXy69EReOx
so5O9f/ppxgTvfyr9FEDdAszkFFVJXoLB8nc+/tsIBa/6fxYWlmfhBnuykzWW6LfBrc5nrenPdpA
3uHHaH6TWbhxup4N8qmlMXz536Wlqre0kNpAVkeWRuJaojWuAFkMIjUfrgWZMmFdYXMR0y5cFjp3
BcyLUAzkZY19YFG3LwyNzPIr8/lmQ/MIOqqf+pylJYd8ILWPnh9KlJRYu4Z5FFBEkekKOHKFQTxn
mZCR3J/efLLOyUzyCJko/lnsZPf+PrFt9E3k+2tR/MkF5mnjm5v5zzUNbvyKKw0Ecyl79RahAVu1
X77C9ewl4PVyHl9j0BACZ6sSKkVKPta7cyr+mcAjPlC0YMr5QOLV0ry0GO+2qq8PmcuQ+wqtfOW2
x5XZfIpZMJLUaDCtiDTTq43KDqs3zkRTYW8xRPMrK5mK0T1EmDnHLWoh2HLaZWS6RQdDBe144cp5
sRZqV8HF2oFBj1PvSbJkMnmdL18S0DQE9xLobC10+b+y7+yUt8gUfdOUUvkVGVKww5wV4kmq4pM/
xBXWziqtoOmIt0lKP44bEO44+J0tAiIN1UMJgUbNrSgoPYsjrvkuhFKNDmBSx7lI1MKJpEdP/2Ks
AN6jGvMgeO5HvJiPRqWlKBhjV8bKkBMCwZR4vkhibqytnqMy60xJaki7HdGfWzVgwdxaaxEGpby/
YmWxzt1v3AN3zcGPG2NpI5Yji3/IqWOeXOHnwl4qcBZSo8IbN6IBeQuLMqdIHg9+YjljIFW4ta2e
EUYorP1fAcYiYD56vHmdESfgv2jOBj9MpxKpPl5sYg7ZSkJ1aBgZe8HsDp1mFvGMX2mRL+cgWCWK
e6ZSZnq+XfO08siSO+rwgSxmaCBRaEIK6TZshL/iNFpvPMCHX7bqzDfpZrTbW7w3mZ6GKonl6QeB
s0ZxrdD5ow5b+ExZBLezePrQTv7O6+6+tQSOp4Clt9bjSdxoh/Gksp9lKTvPybi2EoQFVPgYg+k6
FZqI7JN2NENMW4VaWJ4gfY+DsUHiq43fBIiuMu6K7D5fNLoOtwzczPj4zP6WEF1fodxjhQnfHaVJ
uT+JxgPw93R/CnnoWkyyUZrk5AR0cOSu57GlMQ03k/Ls6w2cGU1G8IAI7C8BiX8lBYlvfyjT8uvh
cne0VlEs+OHpSWrFPsGGbQ+BmCpvRIvpn6fXZeZrZy6/DE+VJbUe8vSK5a7myMfEzWiEIitQdI72
PemLHUmyvTdE4u1eowS1oay0BtQiOAIiU7oYaFwme1E3JVtJBBUWqqo12T2QidIFwV91rjAKIt1o
ot3oNuw/hvM7eKv4UcvKfTMSGbuMlUAyMKLUG+dW+GlyPjjoIesCUCoGUEyBKBlRo3/o6u77e1m7
fravFgf9srRCn9kEPnC8Tqh/Fp/6mXFPydHHeTk5QToIyNDVrOz2FckF1wSZfrd+XaQ07Lu5jNhG
j2KWOrRPV9gvz//BWoWIakxcxw4mxHjE9GRtOCKdfYArFvsfrQWTw2H2aXSRfysb3Pr1z7SFCUNH
1oxXuMOdsf3N//jLpxzalhsjHOj/U1HXIjKqyBPf5UWGEbyCoQ/Xlgr51+3ljr+nbXgjaNz0PAk9
iJsIW6oX+zJfoYuVbpuSoVrrb6wD8m4G/jZvqi1ToYvQDQfls4fx2AIRMPkKFxqjJzhZQtupSlut
ltEuScOnqTKc4CI7M7Vn3BjM5WBPvA0l1wIakARPFRgRtws19O9ddVIezh7yBghDjG7t+Zzsk4R9
TYS51iyoPiyDdEIl4wIpj7e+GLtoU2zeXI3wqDG7QH1SCQc7HcJlAhJXEfjw/sSjWK5q5gZF23lr
OOytZxIOxLUrCwGIdG/2aF7v9Yxm/5TLj/F4Ira5ItxIzl09JkuJvLhPFNaxJoOiDGJLPB+bEpDQ
IxxSxADxskv1htA7YXkLjKccoNFMeoiTYoKxifpxDpDChYvvoWaZFLegPh6OAVWe3msY/EIWok8A
RtFHAfklk5dXlLfY6Z/xGCu2TMbT0WT05mMTw2QQu+Qsynw76AIqZU8vYwlxlbHRjeeWhUvYt46h
OgCTXRq6OEdmKueiojkA4nYjcHyjcBk3BjTbmj8uFKCvOx2fdny/ftejv/mK3dZQ/O0IKNDx5O1E
FrYH3VrrY08BmDc5+HXRCL+mIifOQGGBc33V1usCw1D0Alo3oRqpvZEirBNW/FtcbqaSHCYDcGSn
CYbexdGTuQcz0nmkX8Jigam66s4PlC3HffF9q8uV08k6fxf+M59M14jLrh+M6O5s0s4Sna3LpI9K
G3+3MtooKJ9rHxQx4lV2N0ceA0evP2oJgITdhhXR9J8KoI80IsyaDF35NqVHdba4UwwPD8vVo8bj
B8MIXHnwXYMQvRWr0cKMg+RQWJa3g+nsSQNvDsqFuMwiV7AVoqEdgoW5/ht3o20zt3mp+so3dcFT
Qk+xe9ANtn+fC+8WwcbmDIg0u0SvhbtuLbBeYy5c5+oP2U+gvukownwg3p93KmOKAYbmiwkHbRox
mxOhyzAsXcxpqDL0KUkCuiuzRzKxGYrRKe66lhzWlt6kXqNOoMwSlLYbvYCC5xNmGGRTh/pc2tkT
XgAnJXtSQJZ3yZ0vfiVfW0hWWf56pkjvgFgvNalLZH1Nq9kxWVB7bbuNbLGjZHSKDYbl9vxFLqu4
OkrSnSlUUY011/YpP6Usfp6bXIuKqGJtNkUlh6Ltwp68tcxIai+3QnzUGRa+2NBavocgqLCnNt1I
HYv5LLhacmtxYZ6xmzPsO/ov2BaLGNUgY9sqkCBe+5C9uPphLOeTMhui9zt6jWf71g8R/oibYU1T
iuoVF1gze72ne444x0/uvR7/n2Vx9aRsmaJcBpfDoWe9RHJbpvBFhL61pJOiGBS4q271BdyCTOsj
3D9AzrdSdan0Wz1IPK7dgigUrjcjwa3C1rCo2mDV7xLHCoL6rv+DdsNYsAcZiXwjTeJMJnXXpe71
zEBYDtNM20CjFTphHn4xb63tNLI1Jli+zgXRxHfUtx574dlK9NscwI6d6VO0bxyLhSTu+Y5NqgB4
8B06zY2c2E430I4vKZqemCnNlqLFKv8e6KvoO0JfZhmtgqchROE/zvxefOg85YOkb4Jk8JcoPSyY
uqjcy7pL1ARwFYbt1vMzrvx+x6GjTylebkVYdsOSTfSn8K51xAwh8jqr/oPTMdwYcx2KAWJSXW4z
7olpd2f/vBnw4n3R6FS/SNTVdtxAkY0JL7p5/mxWxNFLK1yzOlvQUJnr0u6j1fqO5QyIWtV81Whc
xpkn5eN8M5P/rx7kCb+pg9DtpiXt1S0OWC2w+Xf8bf6RLU+5JABMtR5ULASbDR7oTug1Arc9cHj/
mtt3EQdQ6BslTHxjtvp1A6JzOaS2ZH1KGupEB4Zla8beUIW6d+nBrNbszttBcAaLUkfg6LEg/2Ao
s8nxiBTAf62k+aqQBR9vALZeRqNKAhRq9bwGjaCJP1uYy1EyhzlraSzCl76jI4q5ShH5WQk+xliZ
+R0EIYhMxRin/mnQQRrw60+nGuW+0QmIBlgtU2QzynKKYcb1gAL0J0dNfDwtDhSbdY4HANSAizl+
pDmpktv1oz8d4TiVBvV2/ZH6B6ECQniijWbz/tKuDjHyvEHgxZTKR41khv/kJzkTYM0z+h5VR6Tm
UZBSAS5jGCab9Z2Xm+Ty0mSGiANKO27zo8tqigmAoyh1LCDBN3OyXMryIM+kiKSifXeajLNOFXmF
L6TkrHnxdzLmMliLKw4cY7Q/a4EUusuB+FpkpPKYkpTR+m473DRVNBDfnwKkUmGFX8w3Blz5Jtoz
ONn6oN34i2OUeqRFN8P06ig2abset67BQaxGnaXVchU9ZG5UWvnq0Tl4HbO6TzbmDgTeIsEAuueP
qbhw40FzUh84Ai/gY/9lzgmEe7LPKoVN49RFRo3EW7ocVeKPuk+cvUKKrc8GVCyTA3OaD2T4+qzQ
ulDig3GsdpV2dJNc9WIucpufpBYnHdgHR6wGsLnvz+3UbTPR3bNT2pyfur6li+cDu/Pq2cXLXw0w
OcAS2Qfyk0TBnry/FBmASxD1CO3tmJcVD1a9nL5KmXM1GfGNsx/UW8LCmC1L8UjyUpp0XPQjO2Sv
So0voBgHKLxVQ9N51xryDBbhdf/3EMVtwCZZq0ruF9ZLBt1WOarOyIg64Ec7km4A2/tNjjgV4y8N
1qpqbDE6TGIFmw2vRiX5WKIMYQ2CD/RvRq27prrBRuvd/n6GcZwL3wXWajdR8rOX7v2+XXGbWYGi
+cOYECUs+aZJJSO4JJAPZcOFwbA8xcmoYUtJ2WRgWCwirpk6X0349Z+R8aLcaY4nQdv1yi1w0MC7
2sj4ITjyazFLZphoPJpvjFllN8HcJMELiwXjfIp/0/UB9f2e0OQ0nodlvmZwQMnUfcmqIjbv2dak
oK+eDpHY6/lDtGHVk2LJLOD7qUjZdQ7KO4x0eISvXRTvabP2XuiEAEGv36IB7vqiOsKwYgXI5AU8
mqHFV5+sO21bE6oMOztrqpDoRxpRfyhLd+JUCnYK6iwi/GERevfQGisI/eNFoTFlJ0B5bHj+3mBC
Yf5+5rBVMiL9QBsJ4kMo2BjjQusIsLaPBWlIfLHm8x+1dGqxCuVG0KtHp3SZtWdnsoXPimqcE0/b
BRIjj11zXX9/BkWbmEWkU/lqsos5RKaCUIaT4LglHRmv7zYULqB1uiAGhQXEJeZ+/uAeP+LWNbDj
3DdXQoYbq7P0AUw5+4QyA0NQtI8hYwX9SnclK8FCd3GMsPmDWzkc6V7TzhUB9jKviCZGQpqYTVau
18o+WjQYXojIMKyrRqM+MIQmEjzQkKCFJrOoWwqZtaCezrjqTeIZvw94llC2eT/U8YgPKRGDYZIV
fUDsHm/xWbYOgDyZTEqecFp0v+5+Gl1UZiUMQwn6nP9Tcq9Y1a42yTqp5ENh0RWdWLi9eyvAMlNE
p1GhVMitz8KwJ5eRtxWs2BL6U9NljVWWRqaT1ugYkHbElSr8uqOoFYF31TDGWYIM13D2LVu7vvgP
1eHdelX6ceuywfXqcVxucpE9U3kNqICs4kcykOMvKZtnU1wcy1/yYRN7DodYaErv/OURxnU01nVd
LPh6Ob6+0vqJO3Ohv9oaXZD9FWvGuUOYcVjSJy5VaZA7v1ohnr6yqGO1o6mrtOLdrgT5uO9TeQOV
RUSkL1e3HqH99Z6/edWPUpPM/7Quy4K6E6fXwhPnDckVAJobpuT6pN0gNgO2qmdVLdud3H6PeEkx
uDOQ5ylHfQ/0a5S5MJcSyqmU6yqL7IlCFeWaRZWRvoFs6ygD9dxupCKq88PHmX2XUqT3eSp7fTjx
/szixjQgsDi7UgcPFM5X4aIU4/SmKlLWXdghJ1yvj/wm4qlt/2havrlP9D9NRQdVUOfpIV8b0pe9
V2T2LbSBeukzWek9Ee7IB0zzmQ2FYVfS7jMoPanRtTMzTDuFhbMvgFMdSp2OdQnnpFi7SXtH2BDl
oOxbuo9wepIDA24DTMdnEJGZaUByqVqKJGDYFiR09vV4mh/LSVqLVgKGq6Jdbczl5qaaXEqjwmUy
BXv625KWsRk4uTojLwa+4mKG63687GINi817DJlFW83zy7OOUUynFet1b9COV0sKOHgIZ6dwTSEs
+9CGYgJxpwcGmAiQc4JSZKiM798p33hrEjlGhPQeGppI/pzWxp+UTefDeJLbhzwh++oI+m4JQs28
JKLnTL/jCd947Wi40210Z+iq3ZCe5XNttPTrN74TtvMxtsf1j0J5Zdh0yLR+qks9YSLbqPnDpmrM
iJIKzwqUokL/Eys50D2Pgi1Vawpm5rYzCboy9n8+NW8pmqBfO1/3fqgJ2Ptj6lnGbcYg1VbOZfmP
XtKpozwlv6QFVfWAEHJDwwhIRYjEtVYGoOE883wg3wdom7PkyuBjVJrDO4GiA8T/15KmB+rebQFS
xglI51lF/OdgDhWcBjXgZLp1/AMrW3MVN5LXXb/cICEWJrFLgWN/gbcly51lJYUcREb2usP7SJ7u
1Et0mD4TtuBzjUQKJ5xZQdptQuiflMkIUS/E2+4iVHxBE7tNTlEuMWpp9B0XBhQADNWlUz8pZ4OS
K0vU5LdTr+Kq3ortXP2P+NIsNijqAYg63nUkbAHCwRGMtFBcjcg1g2TRlh3KbVB0qPYTbJR4GJ0w
5MECGWB1fMwUV+mg6fTqPlJb7tfm50P/OY22eq812rjseCmt++N6pRsc+Gujf2aOVshf+HcVBWA9
iT5+RcP7WJNgetfSyDMAuDWDTiR3QbPMcGtL9z9nX3kQ2NILIcjPhAJmJpi7VVVSnpTpF4hCtNMr
gQgO0XpHXRIlwCpXwIu8Mi4a3aTbPENa+JeppJWT6obOE0Wea8JdGzjlzRHJqc9tr6G9emQ+OPEv
0+PSGSZYv8V2TL6Xq27Y9VvafZUmSMpEWAkOd0/BjLdQi0FiMK9jOb7g60BhF/BHm+KFNBs/6F+y
4sR86Oi861sTfRoJ+zD0lXUMe/VAPpIoBl8xkuv1eMXqLy7WPow28ZosCeeVWMKhs/mNXGWhnqwI
B2bDU2h3XyQkZTzNxEYUlSUuMg1R+eNkA/SZHWEm9EUTW0amwBQanXZBxZ01Z8X0b2Wsp/xYpjMR
/vdbpe1qjv4d1bgPVhNWFMXWEgdl9QnZ2ErRrt9VsZMbgxHK1JVUi/MeHIfqYKvdwq4bGXkOlT5v
Jn05A4Rf7Keh9TkKApy0H3nFlXdzoWIVkNC9FhrhW0pKM45RtP+hMF18DToTT/mxGl1oixgfLmj0
z7qdMyPF0Ut2pMN6j3JhZtKOCcgvJwkZsz90Te7bF0CFwXsPerWzAjzOBVAY8uhzrVfwYounA8j5
2It5KJbqUUaD3oXl4TlvIe75bF0hfeBihA1zvYtv+6yVGrJZX85l6i10EU3TvTsDa/nld05gQH20
e2yanXG4SK71ZignTT9E9FpSV3VGVzpZt/n2iDj6C0L0gcuQgHfLhKHYA/7Ms5rTRe2CczhrnmEr
X/wCd9mVLQOmEUkZlzmGO9JulIVEMzXcNlgJ3JIpyAQGgsxhUO3IYDbYUHJWqSra7dVxm14SP8Wv
rf013O3Spais/qccUp7JuYb7E6pOVsdQ5JdztEbqdPyDq5VyMEfYD1tlP3ST6N+5iJc0ZNjvqhIL
TgNA/TNet2sI1aHIy8rqrq0HDnQ32cLVkI4GY4g3EaPy8usvWOVNI/cpIzKyhsLi5sthlSBPg0Lw
GXMTbfb1iyJSNQO/bsTd+DvKU4yow3jjXsBAGppIYsxUzeQeMJBPXsUlwaOgei+OMYO/yDqhQs7J
uazxe3ZLMFYVlGUtoKMGGQLPQkYlakWXlDJMtb4KUU8g7PWrEVbYl42Y6DRGDyZlsnwkEGjpI8VX
XOZwrxWwByL6G2KnRbuKjXKLHoeoAN7TKEiLdEdoyUMC5ROTwuugf2p21Xl+oToX8bRu8zDu4TK7
dI1ST35aOpnJC/o0uxDZ9JAE2hBVlvKTPYhTIuUbCF0b0aQ8EomNmKq88H88KnyjhTbsT8Pcd+k0
zZG+i4mZCTxOSFYtm7m4mUxanf2DGpJca9kCtykgYX9yobh1L2WIJbchD7rKyAnShRckUnqfKAwy
H9np8njIpZrDgybGZQhiYA3XH/szQLIKx//ScjuVn1KhyolFk4CeVCRvSE6XrxdZ36WUEmNZ58Qh
wjOiEhPrJifbnNsNPaMBoED+hFXXuLHZP6whlkojJ1l+Yu3Bb6J2BeASDkQB80x6zewRHHzkcOqO
M3wmOGdlBq1bqZyBwk5VBymSpF7HHlyZEINiX82dCR0WaoBbAqUTMzGro/acWe6SCzkfcfH7wW4r
ObTUJ6hL5T51ACwO04+fTFbc/QGiqan3UtDW705zYJ2cCTGPQfkNUI9+0QHPUT85yG89V93o77Ut
1Nqpi/3u2EozTcTAgTn1q6djEBY1fWdH7x9RlMONVuCEXXLXtYeiYTGD92vx6YNs+C2FbuNUXqNZ
3ug2D/htg5P5strLWPrTi1bsrGrzDR/BwFU+cWVq7/2XPU5Jip/drSTorfUPr7pNixknf4DVDejs
BYA+cXm5rSOJ46PZsbkiJlPSkREerL4IXCVgxyLO1Gccvp/6AQ0GbHbCgQHuiFzwQKSbqCdjZyLg
sNnbXw2y8zk374NJEuV6Y7VcTGwZA1bQ1343S8gfkledpmdBVRkZtyMIJgWhxKkau53F8uuAj+xY
vWFYiO1v79cszYFw6LbQPrac8g/SDHVUH2ggO6ujnS+6aQ+VtLcHcDBMopJvicmY5BhHsTgn5F+j
pNSj4WvmTPBQEnX+fgfTFBE6756+dE7ypHt2E76cQWQ4XpFzu8B57oWUrcplQxgeV/5OuXpj65Z6
BQF61k0O2E3InxYhJ6RvzrtUzo+ThjkUFD0/LsDRDJ7n0f8U+fWljFXxHOCbUHA1vvj6ssEFYPb5
uPMUkpkFesxQQBLLO1otniIRGN7Z/Lcn9m50NQORB+mcZ4mxSumjOwUf2OTc4eU0U+r46WTB2MBo
BlqBWrXe9OMOuvFJreUMad5f9+XQBvZbN7tr91OSSSXx3czf61dyYl+mCkSQJUZMDeL4PoI6wuDC
57bxf3ztuF0YFfnkSZDVtWw7dUoidwP/unmRxMTBuORLZPPaqCtujoF7oXeNftbUcwIns+KvO9FA
CaUHaPF56Lx3/8q5aFdg09cPl4ERLeO4WcSYV5On7isqJfJFFP/aKTgfzQ3UcvdquocUXzi+MEW/
ChxVgfp0n9DC6NQ1sp12Plb5k+toFCHWMaY7VRUNvE64F+yHzaW6H4oxE5LJNCcDrMfHd7XHMDva
m5r+p0grrPUP3Aan7+2XidwqOZuiBJNQwB0WmIj1d6OyVfFBwBos2p92v+uh941ajbYG8bOWANFy
VljeoMvUvNsgzi6Z5C9D6rfFrafD8OYKo7SyCHjTZIVxSpOChyQ12B3S+hzkJdiPltHwcj4zJpJP
wXDbgY0zK1LSOP+4R4iWWL7M7Sx1fe+tdz13+U+FjfQXzoaLlKBMNLIFThn/bB4Jee18PN9Lwo6U
GVPUY2MZ1wLsgVrgZK5HqARPbJeguwTr2aBkgihBzkBdboBWnfk3WS5+4KUKuzPJGQb+jBKJhLXj
WzOazIW9orGz6E2bSnkUWPOwNjQsaqCshlE4gzRDbAyuMfxT06vCRf+YazTUs4gE2t0Ovr9hvjW7
3Y6OQmmhshtsu5bUJ7j1T8ODPF8JjaVNX5wxXdRMpoudPlGn2wL+fY4Y+mZpZGlgzHPxd4cLkxmE
lHZ0M+W1rtcfkIL5oxdnMqQg8yRE82EbfmYfLIBZsZW8MoeMUXsX0vTbQvFGj1szSebQXmfQcRD9
35JT7uZEkWSz5PnfQ0w1SJ4qwVJZFVVXUQXg3snDtubFfCXu9ACsBXf8O/JPUwLvOBeTykOX50Qd
kS+H4l6jRBYXToPJGJWcrDv66l1VQDe6hxAbAkEceK5IuEdcQ/m20PLI0Zq/uhnRIPeTSm4WYVMv
tiiCNeWG4dH3P/Eg/vo7h0dVRJ+dpjkhg9cOLI2dHQTqVlsndLoFYKmaI/g7nm3APQDMga8D9UFe
3SXXg2XQoDzqr+XUHR+nToK6dU3ZDooUuDo3poDhTxovFiJaDBa1CQ2U8teFFXhOUZisgOQp5BsQ
KQrPXxlMuqrl9nSzCkDTdpztqukBUi6Lyw4z6b+AYlwkjuFcYQVTRH5n2y/rH48YFDMFuDJVOoy4
fGatAGFyVP/v6IjrPLwamPT0QDnZLubgHRczav77JEKcdQ0q0AbpoRDfNsCKnWbdfEm5b+USH8TT
SiWuKb7JjiT73dIy0JZyyq0oCoiRAyxmfjot/VTiQO3ixwcP6H9nUAGtBkcqEHgsJ/af7oT8CD8m
VWlBaV26BfFRdkZQbWexVaDUl9L4kIHSEUeJJdhkBr26CZFgXXFrS81lfpN5cMmLN+nAWXlykdA1
oVitfppu6NJJMinB8RCA6BqbrUEXHab9XOANaiMk+XQ8g+S5yIsTv+L4hXo2kJC6cntn/HdMqQe0
5gG4/OKm9eY1sLePwOvKKXaNWQxIldvCpnmojXxPze6ySjQ5yU8KASMnY+MqMBEnUBZ06Wlk6w15
XD5L598CtQlFhyhJ6L58N5NKxyEThNVt4p/jnVnatu47tlJBsoZK/s4aeAaHHwup3UxDoAlDxlwW
jRzNiuT4HVytZvcvnrbwUY4dBDT57CVXSuUTCDh1YqSuR8UOOFy/IAePUYNzPizRuX4mqzExqZPR
MO80oZ5cM1e6SOD6z8nqOr1KQUoRDp+7lXxbMtjDZ3AfsukI/zfhldtrCeIeS7IorkJMbpKSTdxM
WVJ/K6YZ8uET2HVHw2PyZYoSAsGSXJHGRF92CMtMHsrE4wDnBFzryoLUhtu3TCQiNlJSoR+yj7PY
0PgPJwOTgmCpy3tZvan8/4suzb6XBIMcHdqVdmBwwhKrZDqsz6i+MndClGj5CV9/rz5rU4011Dlk
IefaqAGc6n9rE70iqsZb2sJXsKpUhRSRD8TuQEGR9huC5iVkytzMsARTUKatuTAjHJ1cykIg9i2Y
RDsfcJ3Qr+0RaAKDhPeMeRAklh6wY1Zb+rrSKZEawNszrnbtvu4q0iPZ3lIaj1hJ076C9+3q9bG7
UiGwE/YhyVkw8JecbBo74X7ZBMtk3hhKeTgXcMvI7lhchtk0pTszDusJXmA5kbzn5GNB0TiEWXkA
+nswoyM/1UUMegSmdjjgfSjYntfbHuAFGKhEYplsManm5G5LmlWmxJw25osCZoyfwSNcesNPjsbb
8y+Pvy2sX/b/75COmbzMpTlHBF1KhBe3qeuMO+HCrcjfS+FgbUptYcubODB2VX7KDPXjJL5m9EJD
/C7RxZx0/eEg5pUj1EpIxnx8o+JuOq8ps6DYqPi4zzB8Jvd/gF+cbHDBY3J2NJwGacZJPE4f5woe
/Iq372AejrCWM4aBA7oCT6n4Q8pXH9DhHuHMv2AcuJwrtvU4NXMIJrxpmLa7TFEajrTVJq+NLEgD
wzPlcW9EddYZURsa3gMVdbBL969u03+92+BpOY6fZBkwtLWAVuXby9m/NUn68Se6OFBycLEEQaWU
4V6E/qwomMmG9D24rOYM5EpJ5i8esi+NEBZfdypltzpytEimno8a5eYWFTEiS5HDeaCt1+fIJsZ6
b6DbrLPNIeTsr85uPExTUeSWcthPdVc9RSO7GqyF6NpAFMiMAy08RrnkUccq3IfFyGo8ZurtDjCA
tazlDAF1cE7mQlxqivkaRSuMmEuzztu0J7hC/r3+8/o6WfASeyGOWYD1c/FJkK375ujPHNoQ6+n/
NdMc10/J35qvTBFMOrfCeo7Nvbj3BCPSNyCP0Tra7BdvBWboPx1XiW/PZ0ycn2kLc7FHOeMrm8I1
JrtFV25GdciLkUA2IWh4dfxGLakurWZvOu+lRmCnH+uCDsJCxZ8PO9MtqkDLXDdVD3cU1Nj4lAST
yVNb3nPPB3hr6sGMV5J36AH6UKBGVnHEFdLQ/1QBPLJLM+SAJGJZXIPkwXKlNaAe0llKSJYM9Lxc
gQGX2ARidxt/tyTqGstO3CNOdxSikCWrS+1HD1X2+WH6dCsb2UfAroYaOHo+iYOypPJE68Nj7zaP
JZ4BYyD5LKLV6kSGzVPlpECqJt0Sqmy6yub6wNw5nbUlPpRYk9uiLy0D2/b1uNaJ4gPRoYH9PVw6
akXdybLi7x09y7AK1JiDGCyXDjTmCUv/9VbZYZnhafMyeblZ47pU9J5NlSOct/B4rHRBMvIMcS7X
jE8hKM/ZSEV87aJOUFSEQm0lod4I/ZkhpqpichJ+0Dxc3Owplho17dmxWv8lR0pVKnB3g1CdzRgf
SYBoSi/OEL9QtSkfX7kwsxj73L5+qJaPLRaKQE3qL1l7r4/uI2Gh+m8TfszBIu/w7itmca953j0z
PqbTzijXARUglo3UW64QPwqzHqRuc/DaoYwmfu/l7kxe/g0dWqE3w+Ue6zo0F3ylC85GcSLoVnVd
QMP133tJvqs6lz2HILzdOv+etCyiLDluPxxpDSAY66zOkp2V3dfwRnJI4uwXgbFRW0b2TpC204Wm
5cyAT/TeTHhCEVsw+E9JvrE55htVe+vrtNmhZ/H5Y5nMWYWv+37YugnW8yM5Gy6AmI60zSffEDf3
DEX6xJR4ruJAKtQi8bc+diqgmXLTdLu1qTMVYLJbXyQacQCAHG+8KkFMksl9hWWx9FyB6fUy6YaN
Jf4iyeVOIKWqmJA7gylUknn3pwa5GW/nr9q2ksG+fCWyopzoKbA3FGLZ4GKbtOgA73x6tQkctBrB
XL21OrmjAleNyWdq7+7483HtCudr8NDI+g+UgOO7ULDFeMZwpGEhk9dyMfUPmsWS1cfLvvR+3/fF
g/Hfeut9buQC83FPSkzwUMMmucACrlTBxFtqUkAvnfe/Mg565KYEB0niWN08Z2lHYFUNRqmINQqY
bvDm/R8uEMRnrwzPIOkhiVg8f+BHKBOMYiWVioA45GzO2BNQzYW2ATBYPfA1dILxzHDBYui6RKUb
eFfDQ4lRX1emkTOrtA59xQNDiKtIQPMBS63C9H57JWh9ao0PfrTDhMLYLw4g1ILRo7vuKJ3m4+p0
MtSJDKVmnVlZyuXE6zrnjSIWl21i971mKT1VGIVqZ0q8AtjET3RuXke9zmH7b7Yn7MHZWtUPmGzr
VxhF5lO2IA/jtyKJy1+QBo08FxuvOuahLtZcSGRAlc3Ex9xNi4k8uElT7ye7uIFrgYFVzQ+wfpEr
elexkmOY8mtSlv2IQBXh05tCeqO4Ja15KPEYaGdSB4P33CK+OV08lpKopuwlY7ao7sKDpgxQ7Lu6
X4SAcnbbsRS55UgTkG5Le8cv38bnqcle5imVRmeAbKMsjerXGR4fkMzPzc6AHQX2QJYxKUe+Jgw+
0Yk21gLixvUsMuyWZ+ukut3huQ9m52ycQmPwQsxNHWy7ib7XvSLwUbS6j9dnpwuB+zKZ9gPbBd2V
SP8ySVTURLLdKWQ/21/2Z5il4whLPCD/Jz3wFisfiZmagpM39FP6USonEOmxRa4M7COd3SB3UHG9
ugNGlWXlW4rUScywRTrc1PDKOR9MQSC83VeFYAkf5Un4jANgkM6ism7kPMolgDcUmJ0BvslnVA86
7/rqoFr/iD0cD10z555IppIFSIdrNqiF2h9HtY+hHA1b/gyAcED/2cqFdLgY0OAtIOTkCGo6qH6W
dSccqTCyPcX/coJ758X1PjXgFWla3VkI7U+UdZSUVWVkIBaEIBS3UBUz4gCCvYmpe2yCDbsAtMjk
AgNRcElg0z5gq0+WYeDQpZI+ZjzZkHtIgPXIdN1YiHzaijs32zdEhgdhgIT6+c2t6PRQDp36zjJQ
zVre4SmIKD5pAmsEfjrclQRo+nJ6ucx9jSRNvHhBlqWkDhqx3mogyClev9caLOyvAkork5ldvB8k
8kHWHXAYPlCfxCT3/sQNBaEE/OmvTTbi0aGmRwGjl7sWoExPVo/aZCl3F/97mSL6XJZrj1dYy82o
Up2c8um0jcR9Mk1CFBkLVFkCS0JhUjdNh9ZOc4m1EQqwwVTua1xeIAiKlHbBGWRhiVs9PNsqxdud
rdq58ZG5OusYojj9xMBSrUVNhsVnzDdnbtswwyCXVLVk2q59edpYtGmMumqA6J981JKGxCuf8MJn
5Sqw9S3ToZGf0MPqPuLigR5HWWp0clg+7S3QM2AMCuvSncI5X6klSggooSpqT51Sa2W6shkll1DN
KJFcA7vUd0AxeQtOKFhtjGXvozWPK0Iish4KFG+42l89tVDuE5KOaHhiHjUkQ1eLw4lBzckpCjO4
uGmh9/73KzQWMFSqhYHVnGjub/UA21IfNYGZ/Y/tug32h7Ur6Y/G5JxMTzXOJRSmHNatKJypw5NX
tdiemTcAAJzSY6txWBhKWSY0qIt7GCCpEYaLTLEHdmVQaKFA4H+AJQ3wwk2sLmjkL8bnldeD/iCb
jhkMt1bJusyoz8hOl1fRpvYrumTrYOu9wy/wchjhj27Y7k7RApUy2DCJ+nwvE5RimuCN69pKFGrM
xJPliCyP0SIuwIOqZl9XawSIP/SqK5X4NifTTLUi+/CmBxpkmx6vHQU9EtsAwSJQL2EePAFEZTrw
FZ6QaHnv8xCqNh2FkC155flUvhnge4jBGx6w0mSBzbV25UqGUXlzI3i2C+dB7NGC2us2IxV1Hb4c
DXGkcH9S229+Mgp8iSgxQhU8WcUVN/D1RkHQ6MPzac5l+/YxSG09rQaswp8uaBuIqts7N1klIymd
+XwyRSzMeOdsjx1ooy8gwpFllbvnyeU28p6cBg1fCTOE3x7ZTs+/2ptmQRcAGz4MWAmeIyTEj4pe
XAhOs6j8haEuQ9kOE/CUenf2tJhc7wp4XLQQhlEeTZ6tYd1sAtcTRyqFe6d4Jt9TLiNp4MmPBocA
Kk8XwY2hmi0Tcb8yq5uwMh9EQrC50z6iJh52k13al5MSxx1Jn9I+mGPpcYq3UGz9TcXmGn+VlmrO
RhNt2oc3tzQG6MDj6Ih/7tSinqtf2GVXYQQkSoMpcUs4S/rwBdvLZP7hSrChYxQ5ODczne9KZv86
trZYY3Gij8KYyuqqKqzhPHaD7Ad3djSNuGykJNJr9uKXqNnAinGeTOf+35EKJzzBkG1BDLjN0L35
c8D2JEwMyL18cIRP/h5owxc3sPfIbBNEj6z3ofpbyVR+D0MLc05ccEtE2w9C21LQOjQRD8dPpvSJ
JzyeYRbxX18hXev/eSS/68xVlM5XINs/rrWNTCW83h3+HYQRwc416xfCIu9OQ9IK/W20nM6sdvnJ
DzcUngAi9JSF8a7vxDLKyrhuarf6qCLtTj5m3Y4DNcI6CIty2mSb+MEt9ilRw72xyZDEXvLHWpSi
ltgxw8OnNcO+3CcNmjakwSgt5Y9YrrAdrcNk7Cjk3BHYGI/pLh+1rLhnBdEU23AwznXlHrPHbrkm
hu1k+fOa4qrOh6rTA8s+y1Vo3VxAjTdH/bxoNl1ax/SUMMJ8b34HRmC3sDcptz3JQvt8/25osmJ9
MQeJZH0rNux6Fd08tj3lvBGxxs1Rum9keCNN/87mFFnCRu9DFr0kIbCaca0z+51j7peG/boBD66W
6BZZowHHMS8AsEh0F+b5x0ZOZHhlGxOhtuhe653lLNLZXUKtkMx5jO4m0ilrBLU8I5lW2/Rj+z2o
GL5yWPsNbXecl/dIpa2VyViIyjmqg6stblJboKqRiwEhKEARFMnM6ZBxjziOQqgoZyKUnl4iaD6y
q5hLdgLeTzM6M8UQ5zonkB9jv1EekgfBlyj5AEIphkuKzPBpOiJO/X9xodjyk+HHzRXPvYQBfaPP
Rj9cVaAglor7o/QJdrdpwW3b4NQqtwBvkrC9IMBVbdKihgfYJKv1+Z8ZxI0kmpsei/Yamu6kVZU0
1HvdzU44XgkAOt5P2/4TuAJsPkxVto+oZKihZ5ZC4/NoHxZwVrnmuNMAdLm0bqliQYvoYYO3V6HU
xuPICi2VpLPxFjSsU9jfeANPIT/KLIoxkSn6ijQlZRAS8inIlMW0F6oboENW6sQYnvT0N/rsYjF1
2xCr5BFgydqYTqgpZEz81PvY9FsIhTyVskXuPDKbK9QP/pZ/Ogo3M+GDTqPbcZM8Mq6/4zFrc6xM
q4AURKUaoUlInGq3I3q8AHq37MP3q7zVB/HOY2d9SN3fbD1vd2aD8U/aiWYr5SW9r/HN0jENa1K4
n+ClYB4g5+Qi2H+W3ioXkgLav+pRXCYb3QQ0tqLiuEtAP58tjuRNa66VhletCJHK1Jhw8CrzgDoP
dMnfvt1IkLKhAC3wMki5jNCX3w+uDC11N0AqbjH+Onr8Td3YlfEBUBRHvjYZF1lnlfuEpu64UR4Y
WLS+HZiKxGd5v/W/ZIeGaVGD+0MeDYIU9fFrCL+wbNd8svIFIvov2wJKaE5n4YAcJ/sE+R4QIEM7
c83mkJhKmWiJxMvS8NEUrGddKfdKeh1dvl3k2buk08CrG2BQ2FpbhbTGB55/LKIhvdF0GSxINwz/
6pC3imPtp4NAir9opvKr4HQY4KBswpHvIkV09YZ+Z/I9owKe+EkMFCaaX2E6Mf0pM4/1M7DK4g+6
IOCst94ohOzpXJSHeDSVz1BPzu9Lv4EyKvAdMrPtSoqKGb8QH3M0f5HtDTaU6Po245YYXaBJ590p
Qb52jCFyeP32XSbl68fEyTw0d1pCASi+T8awrZXc6UWqZcl34SumfNNHyu7w3jl3wKpygzsgf/FX
tiBKckTdbBql0GE7qttl4p7zuBbNyO1yp39wjpbDKsMVpYhL9asO6V/RfayfkMRnvJzyeweiD484
+RieTsFGwOUAK1Unnn+Ge/7mE1QGdkjbdhDJ5ScvwRYNN9seDfNh/+4cmX/Qc7vnkeYkg90os8qS
cWIkQMiWhL1N/AqV3Mr6SZWfXBti6oG0nHZjxvCVipsKra98WrwB2YbeJbkysCgdI90M5ZQqiuvL
eZlDph1wobg9iPtSPg3QeDW1+BP3FRfuNhvBGGUrVR80vf/QdKNShRiJ0YEZBd0Yef+wHcY2dD2P
9xSNzDmEDwx/mJHqskeC2vJm8/Y8ih8jN/mtaXiKF8hRx/KwNPpgTPkWtfoYeOk06DYkywWnrfFF
vyC9yuC/EF1w2l1Xhwgg1EFPpk3Cic9VUA5GUI5tLylstUKFcpaxzP8T6S4vBgA8jUOWt9VszeEk
xGxAGK2j4pV66rstTDqxXkM9SVu/vItC1A9nTFcaGkESZG95LqrBS/96Tc/p2p17qkfxuxbFmlpK
e97VcBT3PoVKy/bgPRAF3yR62IraTcinZQTS05H1y0KSjkskFPrNUowlbdi+Dg1gfU1GJTBsXoRY
R1d8+3B/jbRmF48WhhZW12LjXcCrrp1I88GyOOGc75tOQLu5u9qOGCYulBjTXkfurKAFsDobOYLt
iQLz2RAN3VaFSk7NlPOupoGhxIhaLUBREQD0rUTg4Dk6yqKUI2c7qumRgH3yuMHg17GbLGhotMJX
qmtLBknilCzLIkvJg0QPxI6tqZqVSB6RsD2HYMaA9mbIszSOLVAbGB0N6c4ETRiUlBtC4izl6VMl
MoFjaDcddgm4RcIRgwmKwlC6gANGDCKcSEIEybhGNvt7HHzUAfg2AJFSNmafVKtLZeFp9LrAwW7w
3qynQfELamG/VqPrkm72hP6AMT/0gNHlCljxw5CKgGPXDbuXzjNKcfnTUA/hs1W+7RYoQZOafe5M
D6nFZ1ZLRXf4fg9TSAldOn6wtBEcekHiMDZx2LqWfab1yFFHq+L7CdRHLaoCsf8GsvxjWBFr7OJJ
IENRX58c4952dpK4XymQaJnPjI4y7D5SUdLnykAEjUh9a6OBhu7CHQTslkfw5WI8mdghOfzGTfSB
h8G41dDPAoHg1zQurTfxFAvgoHmRxKTVwQj5cytbiyQpZYwiALmsdytwgP9FNs/s/tj3c8Yxj/Fa
HcQGVXF3ELbMUnVRZCDaBwFAtG8qqSvdP19KWVeFn1Ebm2UIBs6XR63gRozRXVwEcFlU+Yn0sLrK
ZHSbjcZOomSrFa5OdLYOIXjbKTwvOTR3Gcl852oI4dpN7J9lQjvSUUlk6Ym4SXdVAjLJwuxDuRym
uSf09AD+By2WWd/tcOw5+nhS/rZX97WYe2SKkWE/N3VhAV5UTZzArtZ+rPnC8jujGnKb7j8WzbtH
E8fdVgNj6hMzmmCsxltPfphqcGxGcKQ4ZeQfzF2VcKvNvAiWp3YokYB+Y2wpMhF9abi2IFJQYnM6
w9K/S+4WXN3o7nN1/ffqls2Vus8KJiilMmEHW6/ndDJDHPnYlZ1mdzRMk/ODn4BNtACmAC7E6Shb
+bKmyxZYPUJ4/auYBGCw5PaIRKZI9Hqww5TuhXlSpMUcCZXjfWauq00mVsd2j8g/d5AAmSmPzA34
YQyLcsN9UhiP7P4zjZggczQ6H0yZ8c2mettVGGfraAi0bSRlk8IVi93zeGAWelPjRtuGaUhrkyAR
xNj9IdYYsJiL/VCENAVSjOCAi0Z9dv3CAySF3I7OqDj9HrA0fMQGo/83UzuCWlCwR8n0xjp02VpB
fBggvUC/hS5I654UQOp/w+EqNmOBcFW7U4Vmnj0zvd0J0HLJ0lb7S5g7FrkvAyRClo2jSt88f8Gv
0jh/yz3IC1+HlWSW5A50druo+GmeG3ZwPGKFzzSn8TxNsV92iDDDah5ov8fWTiJqnTiuw7sW439x
9ADu6vKW1WtLHZ0LT7Cf150Dm9X7H6PePwNdoGVkadtFejs2hJiS5fHUNaxDaVRQGf5xRTPr9ycz
5LfgWqXIL7UyZwIb3S8CNcu/NiuPTLwHmlD65ODHUjKQe1zJ0KmZAotg1IXXF43xpKoZgGk0ij6t
JiDy1N0dHsyS6JKfS6kMHP8ygVPxqCrVr2NgvwsOEKvGUqCYc7fRtgCJb23i5z5kik1nRO23vX5B
uOTmjGiwipq17w4E6sNCY/rQBY7pxN+ub5W/oO2Pm1V33L9geGP9o0f6gakPXl7oi18pRbdNefia
n3UEAe49BC4k8R+c3wyRYRuiscZqCwQTyHEWYEuJ7Xfs+Lnkk0fcHXHKOlQCSuYSkOLD4TCq5uL1
bT+gslQF799CzEriew1uQ+BJ3LLe4ovV3fESzvWnrCxi1hBJFNUcvcrbT4To8dGzspxm3joNl1qT
j5On7aFFBduuwAXimLciIXV/4zWKLu6fnNCRYZK/KL2o3dWLFojJarn/Uvj3lXlDn8bSIcYsRxp9
xXb+DMVr6JhzP9YKUfW7Xk2xeoE05rhJ0Og26lAjkD+nsRWovN+bJ378zwYa9eaZbES2VSNezE4L
CcMGQ0jsD+H1I3VhTVr0AlKrybwsvhawwdPV/ir0jPff8s0qz77aKrYuRapoqUtT4N8Xmz15Nzrf
fRm8khTzdzBFR3oWwT/oHnpmtnSUw0YnNO0caJIboqiEiGUrVVI5Zl3nFV6dCme51fyF/4zHmO3O
jiDGcStYsmHdoI1azTA7w0iB+gMJa/nE/qYUyTr7Ue7kKMoKySyMTwwGt29foY23lV9ckJ3Q8yzO
cqhGjNjUASw8T31NWLkUr9DURRegpol1DfE4HlCwyZLkWM73gDmLScPItPelvp/IF9yTXe9VUlhJ
bOBEPkBZj4lU4MbPPCkTOcKfe12Cpd0rttZjqOAINnAfsbtJuD6u8VlszqJxUQcgdqiNjIQ9Ia6s
z4xtA2O60iQ8gVhJqI5KRQxmQ0NU9g89Q+Uov8ElcQccCwoTRwvIS0YSXuu8gt77GNjxpLMpAZHN
iHlOUgN2FYOuwPFOJfx4ujrqnKNAfBouk2AoE3Bd7ixoShJm5IquUA8fZp0ixZjMnC0i2kDWqLR4
2fr/NgUIcx3lmnj4nCzwhzONHi7MsMDwAjOqnbkqUnPCDD5HoJeK0wqut45W5/CI0vjngZNt34CD
s5tBuyonOI8XpLb+wpDGl3leYhFXce3m9UL3lQe5A5i3AsM/3Fw9Eh66TJ84xVPm4gMrdfDQC9lS
mDqeSDcC+OP0gxr/+DDypDiUyuXxTCwXbtc0/ikEdxaW1h4Cc4KNVZdztSCL3XKZPXM=
`pragma protect end_protected
