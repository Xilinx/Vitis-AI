`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vMl/F3Jn+bbJeZ6oONZAAPbmUyI8nO8pr+MpG6WMo4k8R34R6Ht3+nsl7K6UiWLjHiebbv6o6faP
VQSztkQsK3vfiz0mgF/c23PD8JWj7ETGP0YG7/BLFgTUnU0R5WStJbAfmyrJhPmvdd04Mn9jKgBW
zCiKn5dL/r82xVP0N3o5klZK/09H83hQFuU8KdEGdErKKJ5cwaFBicXxaQ+7qVLR9xqZt7WMrEMW
iBX/ZB8YJWcFZVHDielKlp3r1agEYaQ67LllAdiQBVI25+YX7YvopU6k3gtuHSZ6C65gIjDGiurO
TD57ihw0CDtYs1WbGFVXBvOMB1YDT/8fLpxv+g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H6JCs5wBp0QM993fMUtscOIxGEygcaiMQd6LzQYXmdRksszDiTXRFjkGdbzmkkYxrO09AXJIxJmv
OHYpPb+SCGDumIiT0ikq+4EwqFo5wpo7ZKS6iZW8uYULSyV+llzOEGjDiml8a1NyNGqtpXe8jicc
5hQvCsrJWdjqyD1Z4fG6LEr7l3cCowu65JYSdTLqGrOzQO0MBd8oZ3E54fgDZ4bDuRGb9AJFuNp1
G4+VeqpQNWxsrYseXTtdNdbVmc1PDnPFt3ghvfdXTUaZXaBfGuGAp9B42u8/ZnLh0JvYpU/0U3VG
73M89IkwSVikAv128djRBwrqNg3qmkZOQBBALA==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TlpXcKQUZk8r/Frltm1DjMB/QV34UgKJSVDkIWGmf4WGGchWGcrXI3uGxgffn4k2Hlk0dxVVmKZT
gBx8b+BtVjKvtakrclKcKceHvmtCTXr6fYowtGMegkF+DjmEjKTCBoc307lnXWu2l8ngz9ezOz73
wEYpyR68qSsMZfDvwV/x9I/bL8fxwTxFuL7fGoG0doxRn3jwmYM1W97BqrXwDLYe9FXk3u2sSqMj
qseCIHy6sXtgFbMwg0vMEDN+1XVBcncCHvtJQwmgfnlxiYpE9/nZCRWFZQq/CnlWiQgrW6XXH6rl
BzMx+eCNMz9Rk93sbAO7Z82H8PvpP6dvygmXsQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1498112)
`pragma protect data_block
BclYlr2aGa66uztbYnsMeVtqxujeLoQEdtorHfcM3az/IxkDZxrTvH9aJxWKKIRcN2UEEOka67m9
xLfBYCHcdoLj5i16iUOK6C57rd5wgIXSyZxe6StkuW8m+8za83wAd+QygTg0j8Uh/F2NYCgj5XRP
4jWrK13RUV1N+eJ8ye0JIsdeABe16ilUP31lAGZNkkC338uQOJwJHy5/nahu2wbiDIP8jCY8gyqN
FQiqbChajNOif2f8GhbsxqMb/qyGBmeaMOXXgfG7Gw2eEy59C3sTaggOU4/jYV01pzHAAGXPpgAl
X744KljSzxM/hyNGP4c4/7I8AGSYKuitl9rFRXmNCOQwhy1gxwrMV52e+G4HwrWjPzeJ6N8C13FF
fs+/GjD2PI8FtQS+iVF8wfYq3vVHuGvee1o9DRu0sUJFWq+437lWJW6JwarLRhuSiJ1Gon4zAaDe
XyPbHm4Y3T36vGnjO6nYS7FPp16O9BW0MkTT8JlIbhyrENn3r0ICmm65pgn8Ul8/6lq0osHgJsLp
4Du2Szrti55Cnz8cHoLcx+oQEffAr5oWrhaEBIEIGkDOaZn+fRW+bv31r9NPWSV8VB2McA66GFSS
+a8vTSpP5P5ep8jQAUkrgSPnsjdBXyq9e+oty/LIjkCDSimsWoSuRC48GFzyseFZSA8EkH2E959a
+Iz87kTe2GXGvPrOX2XyaClbtdzCrJ7WH0bdqh1Et/ZsLIDfFUVbnBheCze7oyxKmNPLMyRW4gbc
FI/odl1grVcPCZN56DfNVWFJlDDuVqnS5vRFVihcEaYISU2SSsA2e2JvaTAguVyBnuI/l1Y1jkBp
H2wuUertjcvpSM3TULX8wrdzzXjwetKfZP2yyHcVDnDIdCt8uWrLGWRpeILK15bxpONEJ7djDuM/
r3EAUTlaakRrpVBp92vRMip+0E83RBYyH1yCUMOWgKUbp5roxS2cpIp24n7u6W2mO7L/dXe/Qbww
J4IUOSUddThD0aJHA/AVjOIWldwY4drtJ7VcSvMIxeok31v+cTFGJ7ALqKPUD/XhQG7GR5myQOzy
aYR0ew4snfzJZFg19rrXBVgf/nQMbTMuO70oKy03lSjugHXxh6+Nd5Lu7iKAN2HfOjPqoKiGXx24
9WgIymw2Rq8U5h9SuLH6+ibCDzAH5Sqnd7iixMd1lPT0qldzaMC4p5SB3SgaOMe/v0rs1rksY1AK
CW594aMwWviSxlcsqL0T2+bPSQTimTzd7L/0rj614pICFg+MD24YG+ApKcQ9j/XBfsY2C0rBLVS1
OJxqBMZfhseu4n2lIRaAajurJi2YbcZElcmvN1hFPr+yhk6lcjZ3Zv42X/cROapw3Md9KFY7cw4+
2q0SYOEKHI7UpVQCcid0w376hvPnjSAkQoQz1Bjtticyh6XeYEQd75elQ/wOnQxUiMPtphtrWC3T
rB920IrNWhfM09NNNze4dVgNMDn6nH0o0ilCwpTP5ASZ5c8yaQKEx8MwFrYuf0ntXlEVDRSsNnxJ
0QhpCdVOqAQra7MXFm/aefdhMayZkLDbV88wUVC8ru6COYUyoT/8xgHbnuodON+rZPae2JdLFX5y
OH0zvAvXUVPOTCYvvnTVaX+CGjW1qinGoDOESpFo6cyvOFblk0izAIwfE3VybleUJVEWGief0um1
+3PD5jFR9iMx2GVGgD0SdzR0ZWjr0Z21NyWhqPRvGSZqJMZxsvitZHlKzINZAO9yqwvGcW5Ih0MV
O9v2DIHTelHI5VQX5v7mrJE2T5Q6dIOc2ODb4vwF91rc/L3+Wahn25tkaNBHy3Z9IxnXnVaHNmW0
hZWHnx8RSSof5BoINqCTxT3nMTNW1rG+bH3D70yTdhBb3CFrbsaGpd9zDOXvSgVzEo/ieNP9Eoa8
jfwOEMfVOotEejBIoOOFMSwLTYvU5Nfm0K4/aiUmSYrfYtdL7tYzVYJiyVL8P+43lI3cQKd2OD7M
HZWwhD9E44AnPsZaY/A4r1BtiIg2dxNQTgKE9UBcOJ6Q1/A5phRo9XbApTNHY0GDMmsmoQ0spy62
EoX7CXpPpqtkCuiop/0D8SUN98PDYZ8Llmp3E6k8xRUGlFhrtYHz3UZO4S9PWQBUgTxSw0t67Y9k
cJGJzYzRKJliesNDtoZPdBdcO3jEesJN8EVVkP8adNqzV+oHAJ662vSpn++GDJEXtgb6fxfkZYrf
fi2jfqaToRsmH+JuOaarOomLIU0AVKbbQuVUAveAsZkQYFZjxfWQ54SbjCWhQu0GN3nhGR8Fko64
GoXrrb1kr0CgldrVvJB3aJBvRvfm+b4f23X4KLUM/Gdb8dj2z4lNapR9bvKmjJy4ES7WlK/pPTJv
YuNu3E1Jxnc/HAWRimqKtgcFtTi3TapLcHQ9XM/+DnNSRCLD2a9jOYpybplcJGR/fz7+6snMg7un
VQSAbTpG2LLcqrUP28gJqTnZRYC7Wu5IWeJwi7ogUYseDe91ZPEPTC72q/qTX/6cAOhSmw2TGn9v
Fd86aiV3jQcLzRZO7WKzrdmShegCrkEON1JYciR0Hl6FoSTujvd5Lm6WqZaaUvAVWOnkb5bXxsTH
s2OELy2j6MRoRk47bJu9WEoJTZrLqH6xE91IlPbSLsHKeYWNjjmqAQfQo6PhP2YExe5XNCvBWQuI
SqYK3AkYBABLFIro8o9IU+R5vf/qHb1GXKJY61FLBIKu0lWUR5FDk+OsZvRBaakNIpCyw6CFEPfr
wwghunPpyxNTOLGf/TFjvSqY9fsbe0oxX3RI8r5EETDU32PZMOdSyF4GYQ0lXWsVV+c0RYJ65o24
wOHWh/CYjHNDFQyfW8m91nEKUJqfpbw5TCGH9Z7GDey8c4C60TopCjdVfjqVQ3lo94LpCUp6J1eC
cwawrL4gRRlEdJT6mh23BBQpAAkQxY2aw92tbOeT1Hu2JHWmUclAtKgoUcC2JWNm4wpsKRJRe6+k
Xyht5AQiA6CCUqJt/hszrPl+a4vz355bwlC5CheRyZkosnPYdwhAnYUEFtn/WFOFGjQAvdUeS6PM
bEX2LeYaEL4q72GuRyfOAWI1ysHYPuZtI02T32OwZesJ41L/qYazjRw9/knZbDlVpPgZSp8coWxK
uAJP6DmjWhUtTIEX9x0U6l0/x9PE+Tc2FoLe0eWevpGfKMk+0PVO1ierej94YxON/1Yo8K85LfSj
eZ4YRpDERnNQBXRlEFl+651XhUf/n+RTqKI0kcHkREYvA2Tw4nMSxsBSBizZIQC30drUNQOieNMM
2GVKlAYFgrqG6ffDHBNMcxwMJzJ2fycWcJ/3R0W2ngnZdBTHNW4W0eDWk5+QBF0VvYGZMAVXnjFo
xMWyv0JtwYeaTtdW37EcgKvnADTeR78Gn5tjeLkk3klTeaX/h2qEWSLo/o8VkriHB1/4zZEEAn81
V96nNDq0+hGlscJE1TpF+3/CXoBi1HIn2pPCPx+xlMz8fhxPvn715UAa6LgHvv2DblqbzgxVDZrM
lalVe9ScfZ4sXMhjUibd6pWSB7lPxKL6or5iWO53Y3V+pHEwIcOSx0DTcplF06Ut+POFeAO7rSwQ
2ptZUOF9bQgBaXVR7z/1lyepQvLGwo9Nh6iVbumChD6wVjhNEhArVYjKPIRktkKkPLbGgR9n/fFO
lH/mTpPEHPtWQMpfbJppx0JY2dvs0q7CJ6IAVcatdBRVlGFEnQAVj0+4ZE6tT1pWvN/rE/YJ53uV
zNrOP7RvHzF+S0i7Bij1/HCdqeqvb0xdILWRbIsiXrWuoA8Y0Gvq/5ddluLpJx6u1tp+udQp2TRg
20fYrLZqvZlPYTisS6Wo583fEz3dZo9OxuDJ4wwaCE5r7fkVj3om/7l0GlYV1+s3RZnzD5wf1m0Q
bvvV63LBEDF+rrL189VjI3IAOGJlQb9BKsctcaGboa4sNGXf6qSE8cGiTQxwb47/3fGWv2OpZd0D
xcvuKO2QKb33IRYfw3vKygF69lYBdpzh0mrukZ6jVnLkgG7D1SXgNCFQHzoEwM0v5NZmWF90+o+2
5hrMrXzVpWQinqB1eCo1RMnn+NDpPr99AJqzzxzLgWN3heB5wjUMosFalcMkB8h5tUJ9JX7kdB2p
yyWnKA0GO52hKGW3hwx1cenxglj8NgmZFbQIXkEygftV1RVC4sDBjtqBqRGrVF8/aubLtOITHRcX
49KuFaWuRo08zFvlAmQC31ivy3dReyNqPKILpR7iXOzY+PS8587Wzwshpb31p3r6QR3Hs/IU29sp
w2CTE8RYhOh5mn9NX9xr06HHUlE5c1DB9qaUXzaT8ki8aBOt4/Gd7Fe8CDj7wrsI9khG2gk2Y6u4
sJUMl6VIfkLZ0p8MbnJYxP2RB3SfYhsvldbF1UCgj0H09naG1vsbHcU5LElqfVgxBGHtTYuDl6E4
hHe6e6eU6fUwY4+AVPcb4AtjB1rJc+9VXp9YU5bDAZJ73/fXsVKlC465uam6qKyxWsNKMFC9rWPt
I6M/wdnsVnX1CASrFoPYws/fPjrQQR/PO9MnNfaKMZ2kkBo4BGvhqzQ7oGhMSa8lWuMLWWnMZmFK
iSxIU2s4mtuM2N3WLJ1r7OaVlsBqYCdsz7NbYJEwHhgQ7g3r5bwFqaapDfEwVR3gJKVoFBLNiAEc
DweZG8vcCwGEXBVzmBLxpf5HG26DzVMsi+fJtjwSfsSCevlC4Zc1AC3Og1ql7yjJ+AYtrfyj8DHj
NostNRauqh9lXSrM5Unjp/VM/SNGVl21G/kfx3IM4Ux0nIaPRVqsJWAoJf0mUiH3DOAyKgcYN5km
OatLiVOtprnohs13gReFeB6Dyp2gwiVC6nBhulxveCjBDpyaousKSixPvrty7uOBvocqAY09rYJR
Qb5RLOIeMmMjia3aHIgYFQorTJrB3nN6HsJn3abTVrh350l85RDEUsxLzOHvJY5FSjFlBjiwXc95
7QxZV2nh1whRg4MCOh+liAtQpr2j9s0gUsmKgYO5D7E5frhuX5K29DvI5FTl7CUcIOfkGNukwkUM
ISo1YGub58s6Symdaha0TEQbvUFkEFRVxQekgbdj+Ze7LflfPoLd1wPJmFK9rdkjEnyerj3f5NUn
wvjyppmdqSpGuxEZoFdtpfpPs3RDLlz7ro8rVMdC+KDOvwV3A3StCXyQd/bCdCZz3QffXhA0bZC5
zaqxVbnsVgRrBNoIwE5pR2XsdCbpimErDdQrAJXJ+gzm37fb92KtTKvaE5NpEkv6zDqdLtl/608F
/YMHIPqnnx4STirscL4e59frd9cTMNsVfyxZaEhPsHZ7BB4BnQLRxnr7bITTGHP74Eg5Iqg/wZM3
K7ryBrEbahkpipWHie8D49XB5adL/GT2oRmdz7MeZf3dVhgKoMHtch9zwP5NKadKbYNefqH02VNI
xIMV6cALXyRoEx/x0fxndCm98Be6XhRcibdqaVI7WKK3IIXnLHcUnsFrjw/+ABmxrBupjWe8kNmd
qg99fS+4eyLy39V3koqfa48uMygQfLg++dNrG+LlIXBrIwa4fmwrxqxFTYB3BOwP+vY3r/TU9NlL
JH01bmNVJZOUhP+ldttjckeFSwHnwEVXKl/6UYIn3QyuV0h8xBsmsxZiw/ymeq6Y/vHK3Cw3UAtq
zwQZLY0l2jKRYU6kwkv5mZdZZmwWuYHrS0G/PvpaMfGkKtboXT4mvD/fRETzUC2RpVjuPwMcyah0
HNwa2WpBe3rlLwBsX/pD5wbg9VcuPCdWFCGlJxeT7+OLnGBQnaQq0xh620Lq+xrCXZ7MbCiof/ix
r3Z/2brJ/r4nQ+5jwKhqRupD21OR0QKc/NEgCNngHfqrxe+6zjpCdARe4GAY0wqs+KtuqKBx+mwj
xvYAb1w0JpcmKuBQJbZUUrIuyBwoclrSkl3NYnIBBF2X5S+nYaEY53jwn8Iab+4YdQN+ABB2iylW
TrTbzyBDgCZrsyYmrD/AD8sVxW4WrG/EFiZMy6jjn00d/nF3k7u5iQLecVru8sLWCIfnxzUVi/fu
MAg5Htt0+Yn2fBa9dq0LwvNHP8E7R2GcvHEsJJobYCBv9TgO6rHuprzE/chnfdewd8rMuNgHmOQJ
1b5uCIA9S6Zm2hu/wL5xQxXD9F8D1vO8lOgAnXkJ+TOp8l6VCIjiiR6w6QZe+/sbZKnQp7hyeN0H
LYEoJlwgWLzqJATYl8BJYAxr3XtMua1Xh1GoRQ1vbqlc4A1Hh8IZ1MYVzpVl3AztCmJSsFm0VO/b
0CHuQHrdcOkEyAyKzzM5g4cTFf/pS/Da7CfL/sAtGKZ52WEUYv3bdBUCbf4CoEKgZqhuO9x8Pc/9
BsLbD0bPncs3h4IMc1Q4EyAQyNpTOX0oCFF5u9KqAKO/A5Lox3E8q2q8bTurISJ5A56e54xOQtZo
WxLS5a+8A15tEfLGebZEMCHAQv3yAnNPWqNKBQ/8wu6+a+609Wq63pOiPVekwsrDA3B5DzUvrTBm
Ip3JP6cQumV2y9VAaSLqEn06yoPythWAH09UORC1t69+v4s7EWKwURkBSkMV/4UZrYNDLWRqPtDS
uNoopizPGkVY6iyd66EjZ3st1258C5QKgv1G1WGtU/D4h4y67pt20nbSe/6IYvJmFgblZGuYWh3R
9CX1eItof4SJQdXzrP5rFwJhaOWTfYXef4+ZM8n0tTE8atxYL05pKBFNN8GbHISFPE9aLIejox7U
4EmEa6DrwIog/xc/urLda/7We86u4xs9yduKiyZ0jYb5UdxKQg2uGryT7WTppH+kORe0B4nvA7YA
svG7x4Iv+D/L2za4+bJrMovU9yW4Czvp0PIMkJ4ajXzo0zod4Zu0j21SpFFh/8J0kmwBj0oFbCsl
JHaM69+q9u327mutI4qj/Oy9vWX9w38Y5ktrn79iFY9SazJufcWmRL4UOI0iotRYhkb7yPUMtkDs
/9MyHgEXDtyN2CJx/byFym9qNzuoGgjUeic3wH127O6++mPL/82/8ngpvMHHB30T/Hyx6EWqL/Xw
s7SWOE89RanLV4da115LEMDSH8bPdFUSSv1jdRpRFcdD/yok8Xl6CgbXes8oKpkAjB4yIkSpYOLF
VyU+gI/r0tPeCRJsD4OgV70XRkwch55lB0YNAFCcxo1icNwMAPfkLTi2954+f2hbI8oGa2Vb30NH
CUwHcwazjQiLrwdFQZL5tBePkgcrQctFlKG1U2P+BrTdkRlqIv82Np+6T2TpqvQjht7mwAVju8cN
xzwiwFd8I6eImoew87Kj9zp/BYtWLcNqOWYT9EgahDykXpERjpU+XGTvhy9Z03Idobq36TvPyc6F
50/dwUcH9+ZGDNQvb5mt9x3HR1kEK0KPgLAOAoH+6jL8DyTriupl9x7Mn7WTL+jXqcqu25p8ac2c
zyYr298F5lkaJDDG1mt4bxs9tI3qgvCdv+EruHWGlNSlbV0N0N2x1ksqy8o86uVBD4hMSkCq5UYJ
Vuo99ofOPqqY/f2YvjOR9qkjmSYFVeVq1gxznW01cxFCr2V+qMb2EwaFuWUfWh6gt68UVT6kBrNj
PBNwLsTV/emIxv4CupZ6i+Mx/qMHWmNoNm6A/SnN9PmzYhSPU16gbFhwV0Mnw4DLLvQnG46OCX21
wkEKCqbbtHB1/ssaaUee3flT2pVG2bVB7Ig6FB/nNLzUUUfcBdueGIX8WfQoehHDyMTCcRf0WVjR
e4qI8SoxCVWnXLEoY05jbsIgWj9FafIj3S1QBp+gEb0ee/hRHhF3qN2z8ef3JHqK7DiNrf90Tk5e
nb8YeGxQBA62veb7+tCYx+RYblODDlBGJMtGxSFRjpLNwdi/S/IEpPSa7lkE2pslU9Ys7VYsyZe4
rLKfC+ZclCOZzvLaxWAb0MKxgN+y69KsFqo2PfPV15MFLPLkR1bj3BrXiMMKobeO7pMVSFLE3LtO
lrOA1NmI0Pr6GCcpLpw+qcv6f5AefMEbkcBViFUYP4On4P83lKvAhdLTnwUqU6Xo6sKx+13WSMSv
sNnT3hJAx0dtwonN5i9vq9Z/BSAKAj6bEycLCB2aoS+NcvKkx51TKxcqbLjpOp7pAMcYDl4J3ZP/
o9GNnW8ofr+a3WFnnQDhsQoZyiLwPOROQ8t2pepfT6JlbooMMGBDBH+tbO+KMuuywvrzom/HIUk6
m0HBw1tBkOVdBNEUM2dgm1M8PbVphps0wL6MeLqlVjOD95OY/jxM8PZXISA8GxfWUDUqhBm7LSl1
ad9jvnrgoBQ8A7yRb3UJo3q1IQrzrBAFwFoAFN4fp3bF1Zh2far40/x/H+wXjzGXZbzmMrLxdez4
NucJJB4hx+DSSkLbfM93IJju8iyeSEQCNeFmywHouR4Vtxe42Nlni5qAxp8PiCKpm4Uad6WgV0R9
FpLEcDVbqyL1ZPuM769/AH9lU9TF5oUoRCkRm2jv7GUCzNarpekqP0ApeHm1jbFruzfWVZXFK8jw
MyZF7OwVjszN1BmQGQ1s1CyQ67PjbpnyWC2UKpTt5JRsxSFmC/cXV0uwkFCbNrY96QIU8mQ6r+7Q
H1AilS+Pc4GHbace7U7R9ShKF8UE0G7VLw53v8n4cxZkjwb12gfMTlnr1q+SgsBtYqSSD7M5/fCu
uAzyOf6c/O2wqv5YHdDu/eSxAzwFQWYYzs/2ED8lm3Bf11rTShCt0TSh31qkCxeV7pLV3doguas4
VNT7AMy5W2k70oq1shGL7BL3puCa+QJmyRSld8JU3pDf8ykXywOQz9R8snqY6YwyExNYYiqkVVnd
5x6XebLQAJlKUFrGuio9iUs3if3Q3gNlXdRY8Tp963P1nBemov8AbLdJoNiawK/Ii9a8AvfQChIZ
9BBdIMTcNy0C0fM73fFbNgc8gC2Zl+tzmNRdg0E1rdq4nC+QJeC91njOA4PysbXFTOiCJ3tLFvb3
KoMjGqGzpw1IWlZAZC+8KH11Icohnvi8XyuqRYxEdis2isjpp5cml165xLEny+9AwYnOStNqzARB
b9MPiN0GAUMcINrbVOzjVpn+bPjJKSBQuUlUHmpCwp6sNzaR1LSEip+zyBpS6gRayrT2TJLNIo7x
nsTJmIAEHrYgleetkN3zu35nCux6IaCYTQ0dLkV9jrSA1lFV2YacwnDx/ghkyc9YMQ4TR4u2hOKh
TJcLkk3Hg2BYOIwjgg8o0xXdAeweooP/TzPcCocihMxoYJZckW/M3KtENLOxde6nK6N49xNYEeyN
wGHXybz5grjRgdfKAueecBLZDGjxDzIRuiE9AhQyAP+SiCN0EOtjj6d+3+RHMhMJ3zx8L73vQYYd
KCcaYE8cCceIgR9bX9jH38tKyXYsI3B3LCMbQtIpb6iCkNIOiCe67IvLuZ9ZlXIX3vR+K0MdrKbl
K14maklNyJJZpzphYh1bosrOFsrFzXd/u/sU7XVjeBOIp6WXONtPUivzb/ZCyNZBX+TtXTERpF25
HHS+lLTPMJzTx4qbhS9cVhJyTmTEA7MyzUdNPrvhXsx4WjNV9RlrX6riJq3lDId65m2ZiLbp5yPt
COqmonvURhElagm3Ve+Scnsnk4htmHSjSQLBXlyCHt1nUD2ffunKxMtKyLezBzuWdyVlafCdbOn5
dUVUOvi89/RqmtYZp8eBhD66NeCC/DiwRauXfqi/u6Ewv5brfHMp2OojvszmwpG07RtgZ9SM4Ecw
kv+CrheZMgM4+l6EortD36NOBw6QNNnmoFuBkYs6ZmshkinQzCTNOOM+pU2a4Pd3gAGUmvyEEVMf
kAkMJuZLoe/CS1EvPDLtiF13hxu3+wgbX56XoctqWKhiuR9HI9mwdBEr9fhyDm9pBYz/KIeMwVks
TlJN5Ly2YZ9OJBo4bupaFyu6AKmGtKNQJwm6S/L5SRMSLOXUmxYzr5CKs02ty+fZllEG1XWN2uIQ
7gKkULJSIcS93y81Y1yJHamXGyy9lHVYRBTboBblOJe0ay9oPnnndSsfsoMv1welkOzBQEzYmChA
GbL5GNwEzVrU3ewttNtich9QbCHWu3JgsKsfahcVVm/1wpXLnPMPDWwrLhgRNaXKy40c92K95KqQ
D9CzaX1Rn/wx9u3DE+tWl0iAEo4LvTpG7XFyepmsVdXn09VBhHLkyvLYEt/iBX02Z4j+ylIdyI2B
xhjZI+Rs6u1R+bQbDSjTC7U2N827UkISOTHOigK+MvvavTCUyseHpxOzaQHNDxiZbTb4vB/bJ6A3
leue4vMSK7c5dI2lBXnW3DUTOKg8CAG8BwtUvzakSRtiMbFs5Nl42YMG4bTRULEkqzUeytEkwNXr
uy0Ra2/K0GEGu0dMUjRZp0QjQatpEqaluArCVK8SYt0Zc8Vxwqw0zx1PSkqjTDL1tRSsAgfTXd7x
NwonDywWagT4bpqEwYd5SngpeT5KGX9ICJl4xet36Y+bzCGEHWmdOGX+Drz5T2fXlJZnKMvZyKfW
03zNQSdkCCR78i8z+jV49nnujrf+BYbKNM4asbF9yIx3UZd26RKpvo54xG3N/L/nHKOtWgdfN6nN
0ffz+QuHIw0szN22em4KsKA5koXm6CgU6lWj2rPErac9tG9iIO7xXQaipfi5EjuxfQB8aY09uEf3
/oAlCLHbx646ttlFR5ee1yrfwa3qsN2jhUFJepKysRwJac0xOu9XvCzl5fsHaIZH6/z8IuZ36LSe
/N/VmqsKC+7PlKaD1pmHrQW/o0QHkHn4qV4FBVjbGRYeo6gF3ylDlfX+LkItch1v7HHVJXBhHYnb
w2nr9rycs1KVMEl8RXfCZpbykldJRN4W1uM+eHgtGaZnDA8ve8ghC7uChQMdwm3PYfHe2DpX4Uw+
LcCoy1ff3352Ac7M+nGcmZFTQpyUiLMrOCnhl9vJRztIv1Eh1jdN5HTUduSGd4b72/DhJdzBlmnc
3QsuFPG31hCO+dDrqbZJux1BmVtjk+rfpONByTS/yzx2Hx9L5BQfs3ZA+kPBORIb0EB5GbLtGfv7
BN03Rq2+XujPbhCCJswpEtQ61md+IYMRbJy6eI9SSpb+wKgOQP929KC38NduPXZeYyikJ3KqtWvQ
i/5ts4HqDHFpzkLmeVsZHkDl+WRKJGcn97vUOYOHRs97WeP8gyhHFdwFeR9P53IlGbJ99eSMgZqF
p/CZmX/fOD6wPrhZuxV6ofozQgNQ1KI2SOV+WvJDvp2PfkxMssA11HDfsJidB/WfjraZqQErdFsV
HaxHT1177fZgJmf6gC7UPAR9Iv9m5TqaoMMfiMFs5ziGKRPQePWTaANe6CWU8kByiqySx/lr4TjH
zrvn/VRpmbd5XB68d2sDoZTkPG6d5m0XPlUq/3J9nhXfmSpRJ9N3a6p62qGuRlmQMBC8oPUkGSkw
KvNtodzVOdQkZxHsbwyFtIx0Zjw0h1fxh0J9EoRIR9oGhsiKthpX17mb/CGx7JwmgsJmr2G5NMlX
T8v7s1RwaVmUlRLui3Xusa5UfcNI7DZZS36Mg+NVbEhGJPkMELsLn+qRn0uKUlrhewFuYA9/pv/B
GpypUvUkl6Imk5uc5QE8Xs/Ux0tMq77npn/eVnAKVoywS2QATpk8N6v9lnERHYmJhpPemnObV6tJ
DRz/4qjA57MXzR8J1C8/sJBmUSu40XwErN1gkRgfv0ySNoBYkAM+g4hVEtb9DQkM6D3jyVlhGtvL
YOM32L22h7/4XwRy5HAErXlno0aKw8hBM56vLwlHPKqc643RjV+pVOy84xj1UogCutnqpYqxxg3G
c7a6SimY+Fx++wTUh5nbGo0Rli/EBrM1EK1wyBRr/5Pb2J5sj1bFIth9yc0ZtkRbyqv+sUvTlUQ9
h1IKpPllFVCWKEbYZLikMMN2ALYNweFCcogoFCjte+I8J+cdf8gWpm7VBkYLYTK4aVPwYhHo/xjP
MvlDUG6vvTt5OvEXmWxlXrBfUbJ640NummyfHlZm+obtUv8EGYJSzpK5l/c+Rk/kaPFSVgIsIfiF
3SLcoOqCu6xGjmjSB90tj9stFak/N8KBfSIFTiQmhL/Ve3nbH0qe55Wl1xoWQ2m9oejhkQFMMgTe
uTVpSwVBSBnqbH61/r5XV9AZ/eafnMAOoBaDvpBXbdrFnFoGdCuWxpIbg9Avnb23BwyUk0d+SYxn
ni9I29wbE9epkylsevptdslI3wK+S3RwQTcpmWkxrHbHkGUyGkW3pnZhhjQ/mKfBJub4QSVG7bO8
X0To6vPPn9pbN70wXTD2TBeeeEYWH0a22irYvbc9wLVf6/o8LN2phQ8gZ54yoX7WVqc2CS1pOJEh
TDYtLdp1K9P28KKLYM60LKQMgqDCqY75XwqKF2Zwl4JLrBaWjjPnxKwn5cq1xJxgEyJvUVhiCCsu
S2VyKT2jNJGqkTmKPMEI42btTqImIBdlOeXTxeI8atqNHF6dnMWDpYcrVFCSmERDtZiZuGZvndHI
ZFmboUD1NaESol6meBe/tI5/E3R5RfF8+t/wb1sBq5865nuDdnveuLPV7mVX73nERoxZ5Ls1oaw3
yW8T54h+oZaCwlq83pXovEAmL21c40xnJSY45Jgm9cDt8Iv/Lal9flxPjXPbUQAzBrfeG6nUxJ/x
zxLKADXh1qRrL9zRdg1sufbGzizgB86gU7ToY5N1xBCfEonAMC/2L1Xp/lBrJt3uL+PEtMjvbmPo
UbKioLiz5FBvYow2Zv9YcnNr3dGGgG1iFGmLHtZt9rFx/q2iuj0uYULDjwJ1fhNeu/H8fbVk+VQr
TvUU8HVHTl/UES5hXszk5zN+0sWuJWKm3oESElcIPamqi+22+JnOk8ykJuzEc7Xn9Tl7QwFPmEoC
k9ppOTnWYjBhHof0P0S/BFzKv8muRj2D5LmX0mSxPfG1eMLxiRLzatlRqtbIBdGoh3n1zKZmMPfj
N/HEWz4Q4Ad18Nsel+G2ErK1c52VorGyXtNAjDQQoixZNbDMS6mZ3CNMJ1B183is2P5QPtnXcrin
R29CFPv430HU/4ymwJBvVveT7/4TKm2cILTWDpyB3GLdAzT4z03xhyDiTSrgkTFRX54Zi3MCIXy9
bHN+5JaPnfH0qccLmIL6NZldGaFIFWRUBg6k5/JdKawhP13NYXnCKxo+Ze2/7BhYd/gwmjkAGvPj
jQ3ZXhmFT/RZh2B9pmm44VCalRTT7vF6A9LCJgHNyyQfmA7TXrxLtlBIGYyxQUq/el8VbuPq3xuW
oMEckmXlfmgR6V9KPSihs7eqAt3qFO+QeXAbr+H29qgYuAW4egdEAcS4mebMmlBXLl7eDYgYb0NG
z4kN0URQuidnbC/SxQ4/RuAZVEJO4XtJNGa+2aJNpMn8lEOKunUfgvfb8YUYUUYduiBQWtg8RhOv
yWBlHZAFJ+dhefuFIVNzg8yZRM4Aj+mN3ma276980nOALwyytSEjSRODFvgHmAHcAeZ6XKOZJhbE
b9f+w158paie3xHnURkLXHzF5mUEhexmlDx8jDTWppV8jRmUSm23huXfmrftG/IB64bpdIC3c04c
PHkVN5jTXljQIj5yY6WoL64QjWUUFZ4bU1f3VUfDjqVpJCnAhzbG1UC5z1sX7aTAFLlwrUmPiI6x
05lmDwmNErns8rb1stKJ3ZAPlaxrQy7Yx6oOnlQxVrbpXorv4W73zoZTunfJ7SOL5+AJH7Whvw1O
42xZrgzu52J7embf3Nz3p8a1rIer/Q4DWpJroiQ/uhnvq7FxBAPJhHvscc3n5QFHQBoFgOeI5qTa
/FkU5u+QomhLP1JK1FGo57Smipjyh4oRrLmNscpBtBWaNmWu04hmTdL3MkWv/8dKIoTIQzCCmNgI
X/q2xc4UKeqilZqySbbvKQHeH+QR2mW4stHH9mwB1c/QM+Pmfqyf1pUG6p6WJOeustKcVU/p+vGt
WpEqLk1JrnlY92PdYpe4ML+j4aP15ud/OopKv97mDCf4u54zC0cI/nPSSkLR22Kj9chRGCkneD0n
dLJXxYYZV3LbuuuueN/WMmT94eWPefRX7y7/OhL1Y6EnyH1FhxYsJdvCt7/s02CTS7z0qfIpa2Gt
SpzRssniTheAOV/EknTRSVz+E/XoxV7vToo3AtQGWDLunsVXNNmFyR42KocVkru+0evAw4HtjtKd
aRKEXSKNsp5RYMwgLRSutgOVnwxLpuOXB/VB+a2UBoejfqERTRIu2KjUqd/1nbjoYDdgRCkm34li
C9WhzsFOkWYWL4vc3PA4n4EDT+murtG2Y4q/LU/aRY3lY90HIYti3SEf4ZH5tmVuBLoANL5bJ0D0
vSQ++V0M/BT/iaI8t1JToLxwH9MfkPVztOYz06Vkj8+Atd2rZyiu9TVGC/WLa9CGFcTVNWjJ2PkX
SrX0h62tGfFIMHD3DiiWjDmfopkneeUS8Lut8/c+5rMLD7ss3/QOfYmAOLAMpQQ6KUXwvYrNr6gn
lJ60aL4a4Dd10TCXLCv3dhqoArjZywadPtfodB7ujDka4w9rU/L3PSVVDXYOpbax5US960Ci+IE/
hSMeLUOimfd0pho4xAUJyTnhQqk3jPyCLr9+/evwafhVDemvnWvxZOWjOwf/pDr3n/iDPGatjokf
rgN3IazgChQB0jL311k19++JDlgUlPUvbd5a1LY0yGXXYQM5Ivbd9Mlu5wkqRnfmikGnS46G2uTC
K5v2nAS5702QFZaE2zCv0X4cYsboiOKfoJjcW1QEl2O/m/dSm++r4PX+P7xyWRQpBMeW2pLvOhwP
C36zETeNjdVMRXEgp3uEdC2gQatdJaTHdREvxHxSILxgaCl3qC0jJhJRgUL7EmsaaLr0mboxOahW
hTCavEMIj02deswOgIBQAN/mtLue1io2lptr09XRNylqNzBuPZsh1eZJ7/C8s4+Rq0fx1er6+L4t
Iqsbv0h7o4K29QrfmRtc5xObWuMw0tGYnUWTiYJBdznSrBAIh2FI0zPfSZ+xr32/MBDUZsckfa1X
qlBwGp24YXK+Rl34TYpmKEEAQ/bos5cfwzSXZlzUgTTeKsfnbA7cmC34loD2/HkheBprZr9hqPGO
M5UMvYuiXOtFfNZYtfySKVzv1LIUzYYp93vs6mKPN6OQotER+qXmKZguCiBt1D+2Hii6v7zXkB5n
ohWAPn8Ed/5OtD4HchI4Yt2FJI0hEiLekf9KVE2HUcAgOD/2l0yyUbJT5chR6UM1Fuwyd9aSmZt6
4KK/g6a/qxwU4CX31LZXeVzM0Y5g71ref5Dxd7TfvXDl1acuJ72VkFpMcvI42tl5lKEa0GSPOGxs
PdjQ7Qtpjj0NUfVfAyY72Y+lgSSqNSsdR0RL3Av7CZlbQr53tDGfcZlUoUP5kjpANUALk9BSNLsg
h24mHFbHVWwpw1xqzrtpaOLhlODs/jBgb5L4OmacvhAVCp+5pOrmRoBuJQ2m2Sh7M0oMa1y3+Joo
MTrTvI3fOIAiEdWTTJ33jptlH4efflQE+4CbVNNqHeXFnp0CegpvUZthKbs4qh9hZVTGFuspwSin
z2MDvNi2wfpZ7U/l/4p95PWsXtS+wkjr7HWegmISFojzyOGhvO+R75Ufdg8D24xJzRep9KWX/Bti
dhxs63KbkMMqyTDJUPKYtLeFdHVrVc+Aax82kCh91+uSp7+SFfLcDebBgWscS1foPp0oG60wSsAM
ZdAdHaVgswGbn0nvbttpMEVrqYtbHqB6JNMb2NoQOnsgS24UGaO0FJLawKPuBacaBx3sOp6HTHxh
raGzz/e28Ql61iznU5A4JdIuUQ9GpVwH/Ervw98a4Eya1lxhVVGw9cHSaTZCvZ/otNkcs8sPTP7v
5ogEkfwFeu+gDKpNaxwXMzyz3eDxocFXcAk879Ln2wSHwUDK0yYgzrgUnA4O/REDl8fvVxWrujR4
K3m3BlojNAtMBT70uc+zOd//O/Kb2casf0isumlFBh5lyFJQ3jZlZPwYVnGUOs0e8rggtVIUUqO1
tHCUv17KSsbr+bIlrnh55jWt2LrglxHEUXO+WyZC3LBW02Y0OJu5I3C4VXtbl+b6M0PsyUdTwCuQ
nDDaMzRgg+xf+8r8AQz0+ASFh1NZgOSYF/y7bpZFBbMMzVQBZROtpVd7LHx8nnqTr9d9Tnouh62X
bpJdltCbsvg18Ts5yq+dIvrg2hFK9F1ZoxgGc+3tWmcOLRPUTu8NWF9sIWJu1mABGIkZkYfFkpHO
usVqs6qhJXSxKUUHC9h+3gxspASO+KDOg+wRD+E7U261xwOhvRnWmQUKMC1ndRgQ04X++L4PrV1y
muxd2r/gbxP7wxmWlPpcBy3zH4O2j/muAOqqX3CHDjlckBPs910Nsb0LZOxFnYFBeazOnKpS6/xU
f7ORZI5TZZCvhyarD4w/xUtEu56hwmiy+KezmE41Db3iAs1mxeXK2lFOTRHpgcppIY/bnUSp71CL
M7uFiijUWaFdI1CQ/X7ERSQMoQoIrdTr3I82Dzo7jG56frpEZ4/mYIG7pvjeuXyvb8IcYofGQ3fw
wpp9AnRcas+sc+x1L6sy6nJK1pyCG3iH3ufqgNwpme+YQpRrBgVSjJua2HMeYBv5foQgs53P6064
E3rWElyNFn2QNFyuH5uLsh4NJ/LIPZdhfCCSIO5iG8EU/kvp4SUntuDN16midyZtVgKNM0F8MwSa
cUgvAQnT+2FfnoobTEOzAjd1o8MN+acGGzt6uzGYnzQDj5KMMx6DtDLcwwmz51Yrz7lACTWvW8SO
91YFzxFyS8XE82xPUcfVKdgkfnmL92n7GdrrC7Z1AjB1fu7H1oBl1gbhKOC1J87nlTjuwJ5w7CAQ
bCsWeGBIqzPKS3EY477IL0AV4KoPtl1yYTS0QjwK64wqEwaLZcZ150YCcCakxK28oGZMAbe4URoA
zKa2MKIg/ZYh88QfdL1k8tJY7OuTOcro+W+8tLlIyi2CmX4BdfaydEIEwFFdWtBI6b7BgbMn7j8j
Xlfj89RoloKrmBtnnKPD4zMwOk6KAXHuVz8xk3717GWwHtVUUshBGhXsH92tb12OAFPINLukdBLQ
ouhI8TfdErE+4xWf+5fYSA7WxvPHm0m/zFgWMWaQIaZOYkeSsJT/XzaEZt1/8ehJR4c/sF8ODvDU
p4CiqXtQFVzzdKWbCW5d9lKpB36H+oak7rzxDY3rqvCMBI0M2LX0HFS2uIYYX3yJYU77m0LCROS3
0PHAh4O5EQDnvy3GlPuc5JR1zA65arw96I9njtLW3qltJpf0WUWBwDLv+gEoD2iU0EN4z/hm6Il/
sgK1TBkwV+65Fzc6dCneC9cd0bEJ2gDTtsmyTWBmnwcLlbZku7E5bGLXFcpr0ADvnF+At/b3k8UE
ChFgxF0WIyI8+7wZfhzGXKWVj5bOwa6h0VaT47gcHxxJhMx14sNT4VS4uMZ+zLPj+lvkoNnf3e76
4L+IRys+0Kua0jqq1yn/ch38GhHZarauxJ3AIFuB/Q+TtRJXZRSLOARfapme1fS6QTYgqtR0Vm0I
Ocw2sqJuIBcmjJ8mezD+CN9cUTiJ/64EvDbQ0jbSPI3god96X9J/fCTlnL8QOwDcdCuaeiK1chyE
X7+j8Khg0K+wBrKJ1aUMwbAtUCxCPQ1rF2Z8LWG0wMwUgiJDB3nUg0xAKDHpD9Jp4bhJogbO8koK
LUaD1CXtGjDaHaVdUQ0Pu6k2e2UNRyV9jYCrqPM943BrW/m7DyczEaYFupnGv9Zjr5HD/aYlDjNu
qt7MPTkrz6lzUapye8W6KXW936cfLHX/fpF3W7RgpDhXNe2oIKuABNI9+725tpOh1vFk0eyY9LhQ
/SsTKQTdYgmdLRXJ5Qcq6MJ+0y6/vakT+IOn/ak1EY/eW/M4nTlkCHht8dbLkBa4sEatV5ucyYvT
3lNn6l5LGEEXl6o7kST29rRg7Lk/ThFE+K70wiBGZltTJkqAmHPu4zZZ5YelBp9+FBuIB6at2AJ3
5c+zBlU8Tea1I8vu6ewOZ2vvYWyV8kPID+TOH8Rnt/9WkdOcuxpE2adUlO2G2t3uBSFlLe8jYeIg
9tYPKWnHBCBwnEZGhHJIwoMBmhJBCXOB9pPTEApEVTtlx3emAiLTeZTFCI+z4X4D0LeOS0IhZ0cC
kw3Jk0Ou8DkMUZaQVkXDr+tmkxaH/ferj7981JbVqSAMT6GWS63evv5lJubiMMt+d+ycpF9T34/n
1wFgIuPDHnb2t2ueQUpbHUYWdgmjwLI7qMGtLXiKQKPZ9frU8vR5Fq2k5ZbTjHEsMtndmGJeAj2l
w1erGNpdVQa/f2P/AeVfPMUAXvf+0yhYGO+5YAN0V5soJWrwwsdWZsZo4OKVyE3tbQWIDZ07Q05I
jKaUZSqW6nG72+Q92GidCZDxNHIG/ZlwCQSXDguh7cLtC8KDSIByn2IiQWt270qhtVW8PdWg+YHd
mKAwrTgZ8+HHJZeY0Di21yKDjZLqozws+hfP3REYgsZgXaGKuOf6M84bBghfhrkV1OMehpYGntlR
xYe4U6XLI5LOPlpyeBNBpJdK8sdiIrM1hJJmaJet9MYtSLktsiYApsPAG5SfAb6DBQqn0UPuNkV7
YztENo0lEqnS6ff0jh29zrgj4xl6U6i6qmpr9ld2NZYYwEfrijljHuKI8kfXXsiseBt6bgr5FSKZ
kUQhMy9RZ5S/0yKfooCf9lMRWnMs28K9M6xDgUmUuvjcj2xo/sdNv9ifO7M03m9nozMfOyCPKJFY
NgC3uHgebFj4nCHdjrH2lDzSMTP3Pz3KI13Tpq3qZFTPJjMX9AsOFqedMmInqImFf9RrKsmg8HLd
vKWn/zzTjc/eExCHx1mYrK/6LkYQ435PcttgR0B5atFI7CNw5hKQff5S6Aw+r5AuXTd729W8cohP
bbP2nhwgPvBBms69QU43xUIVmCz2cLkiXH1d3kT11SatwfRtjOc2AHvc2Z8oesLJcLt+bP8Zn0Oc
4CE94LlYf8jEhboubNGtgHX4YLzZ47ecbckkxSTMssXSZFWRVp+sF9D4sH7dkTtn+0MozV0dQ48q
OWKKY+kORfbowOr0DM4feHpjBYoSwwicHjouwEUascJvJH1sKBHbo6LQtaeDol5Xose4O/5NcUQD
NBde+DO5CwfnlEudinmOkHBQS6/mn1GuADJn6FIbEbBOXR0kSHnKVoTHacdQM9g6w0YPVtKcEhCQ
+R0OQULOxkXUvjiyjx9XUkYuwAMHHGssBD4ddSZ6zKyd3kwgvLloH4dxMK1Y4MkDLRwe14sGxTEU
EhE56LuInOTyeWcwrV7jDPreseRN1rf5mPhqhdL8ax51mSMbav95PGv1r1LTGahddk8qIwbI+B71
iPLqcFhQk6pl01HM/8K8bE8nMLMUWI5WpyKu4037Z29jromRCiRMtpLpBdGc+c6niGbB47b6P5Fg
gR62QwThTZmLLCo04k7lp0b9NXhxyqDhAmH1PNVkaHEN7hONfJw9+L7htwUj2UZBMZCUWlqOzoeE
Z/giUqNtdS/JN1hPSNwuS3MrXPsVBkfqjitT7GAiwawXM5eAHdqfZDZOdEhUmPtnR/tcZ0Dc2M2v
HxJAEg0fs9vgix4kM75TyhLMl5vudB916w9ZfZNomRVEVJUIzT4BVoJQWAy4+3t1KZZLes9xdoIs
Fjr1LVfrcotAmX8x6LOz31wP9H2ZFwZdnokMJt2EqkBcl84MtLTRwEu+CGiM4uhbOzqv+nsZ/A8E
WRHNXL/vEtkRTbhvBjOb4zXnEY/vB9mKi6Sv7+dFDQU9KHBw5+D+UjaZRA1kkBbwQhExxM/KK1Vg
1TGJl/ggWbyo/9mAbd1WmA1IRVmvxwPPlVRScXdkCxHxlIbM8gclRBzSLHkPKJBR8kLPDzGxnuvq
r2TGHpoT1DuMRBhcZ0ksMeZsceSBFFa/ZH68NSeNuSHCx78w9t9/p12i9K3nQLHxeM4PmYqln5Zi
gldvwWSewah02t3TxFi4HE9qQ/jCUpx9mWKDlTH9FRYK0OfeQW1UDlazNfASXqW19EvDrBP1Ksd0
DOuutaxO0GVt84Qb1SgGfWq/gNPnr83/u381p8h/u59Re0FU/f9sX6YGhSob6Dq+fpihFtFnw6sm
2wHpnG51kafJWMEKdTnCbiUcoVNM2N9NJv0T04eydhCsMzrO+4rSYyfKYN5SeQ8JRuTGnIsLmVK0
N+bqw0QK1FkZ4b8q+86SRB+7QkPDpARuJ8SM8X6hO006vBryQ8PFDLjFZ2aIR+XDNSlKC5iDXeYq
0QD99IChbGZsHDHore9Jg+Z0EqtdIqVMht7l3BFomu4Y5CGpdX6ogJeiWaeGKtaGW6joxADKKTNj
QltNqe3bd77dat78OnpPs7mjQKtdNnPcS3n7h3d5buAM38ZmaBd9wKhs/XzhkVJB5IUoqExbCfbX
n3bZ960wAB2DGBnFgh6qGnutqL7+U40HmBi/oJJvFXM2y1tfuImtWLxiTUgDDqVncE5Lzi7/R+Ba
bao36cj8irGKBbeFTMWfq0oPM0gmHZqidNyWrj21KhB3L8gjpqZczCXsbewzyqlAH8mSz7mmpxHA
Spz2CSBAQM1bGiYrwS2X+mmDBHOFe/HXbZEP9LMlNB1VSLsrMZaqj5WvLt3NxvE0gNRFgWHmx7YQ
vrkm1VolGrrOG/m5YGUymlScyH3RDOVaRqDB8Z/KyU8tf4U+BJLbO5Uk4DWEWj2gRW6KzXfIQlVR
YBymPBmy2as4IjinCL+Lb9xLFHEbWDUbWfAJA8lfWUO1bPSmp9Gz3WUWuKfSWlsSvKGYgsH83/86
IVYCh1gG6Udt8oMZNsmSa75Lu/B4Q2ycP7vPjJ4A5BZlW2snElCb4cgpcIJ4Yf8zoXgFzQa2VYR8
CMzaU7i1PCk70m6WTHxHT41SpHnPtYii0AlbBHzR3C3hJgLXiGijqPmBFKrb+OXIY/tcURVcJXeJ
FH6heXaL5pqFg0EV0Vmy3lBPiPtKWGWLfHNuHntgBnIZcef08Cd1V2MlMehSi7DbYWsayNWbkaIW
yFkDrApq8J7DC9SMMZjcsi/QtFiuRde1EBEQ41EnsUjEZountKbUvPFjildd+Bfm9aWQKswHMeTf
tb65wlPiTK5tAcrkCO2riG7ZyDPX2ZB2lUsn7/xSIca7IlKrBObqjnbelzyrSzSiwWsVxANkfSeA
j91TXeeFCLlCLzaZe375uHP42J8qQSzc7uuOoD5+9jcz5+1eYhhL/Az/YF3MWa2z8ACa24jFxK4l
3L9z0msS0EsAQt7SuCtQW2V/+Q3diuOaNsrvSWrzcJRaaCFQ7CSgWiYXvahQzqD1I/BTf22pVm/V
B4gqcagmzeMtsqlt9iwcOzmLcVKSc/GzbVtfXyrWHYjrzWC4v8vuoLhtFxJvmEqkIMTrRDq5dTrk
DWMwLVd3DnH93lIKinbWLZK1nmtkRpgTvIj77RLFLyrk5407E6DSECF/E74+/Zd2+lyNBlbDVsQB
2Gv3VIihlGt+Go5z0VvaAO32ku/x1JClGBAEiQq9vVmzcKbUtSG2N1USA6k4MfD2bfyBxnuJGgVA
/b9eGsOhocjRpTWmCctvrCierYog9vPMaunHh5UHVOl6Hb4rLaywosjB8besbon1tZ1mzK5dyDLe
vqDqb2dMqtleCbwWIK4oCKPH0WY4NuFl1D/cUlp3SvmiWp6WZXGuSUtHsYBTb2386WQLdb3G0Mjj
0MOaNYU+I/SD2sVPSIHQPVyZJwkG/k0MXKsFlSRAjT2oBeHNiGsDpsVi80jq/mIoJ/85Hj8D39QI
2PUDcfjakvi+e49avZBjdPsr0bUNMA5Y4Vf8buPZtNX59ESXnIp1449r3PjYPJrbsRAKPG7Oemwj
IOtbuEK7+HF7LosEM5MiuuIE87HBzogi2RaPUdB35Vcsj5rf6UAwCez2jlHAXZj0mktdPCdYkRgZ
NvwPcyIdqfFCLEaMKUUD8rI/bpuHnzsA1OelA5+HzbdZTI74xRRg8mORvxj4s+vJvv0qUDdRqkkJ
wXagx5fzu6Mew/TZi7p8EhW6fwQ9pRo8YvK/wxpTNBayXr1BugTpZIzObAHLdCcEJ0Q4aCvQyUkB
B/8pbrUXjAKdR2FZ1wK8lT3s1HykYCrEcoGJdmryM8bmtOt/7lmqHA6COPpqq0FygiCYbdVoXBqP
ESHu/DE69Xgna+A9XC/RWdfmg20T0fyc0bUPNogof71h5mXGmLZ/uoZMOesH0HRQLOFT1p61OrhY
TIB2r7Z7BOHHLbOrhzMbZX4V+3InQHEsqAMdnCloyRTXniQpZ1uxrn3cCZLS6NRsINiEYC70+1y9
xZnmxF1WldWcol/mpVksdxkaA6F1W+xDRMEyj//A0VgYgM9m2zDRrM0vYrPIFx04SIGw0rlO/IOY
7l1EmVSX9Ys6XBSQfS4XbkJGbkirEkFggTT312neOmt9C2bNMNDhOmclFVm3QtNIeM7sIui+npIe
ywVZM9CDoGEhEmllbJjelCa5tug9wm2RNvYXoIH+gpam57cyAuqFQ6S+fahUCYQ92aUIr2Y0HVEw
uKP6pUa/H161i7LK75PoEXq3ipC5T7YzScJWh2Xok/uACbyTgNydQlKijTlnyVE7NppfotDsr+18
mVhwbagE0konb7jIOPpQY5TPtZuVMc6cEWJ5xDmIk4EStKRwciHDVD/+IEFp7Qy+KMjvzhgyFNFT
hhjyE/gvTFCrfaxaGykE8xGtlyH8e1m8vYEjYwrTx/3+rjuXKahNVXPkL5nS0FpTIfojxAcRp22m
0WMp/63lhFQMGXAvqEfqR2DaA+kdCgEfZ7cmN/kBPObTBWsaaBr6DVWd4T2XvMjYxhCns8UaDhOF
XfinyHFYwVhCWniDNPYkSlYl3whItXYj3TGysJtmDJFLBg1oaz7dv0VWDbz/S7o95bauUYu8TGzg
W05NKLFKOjrmJNk73ZAivMUyjxdY30Z3PTWM6245HNyuD6YFfUN8WFh1+4Uk5xyIrTKwP+S0QRaB
S4rIwTQBPPVWUAkeolvuywWb55nDREZB4teIo8pE63fKJu8lhDfXzdA0lIwDv790MWPMA056jMyM
eNcpQYtM2L2CCoWHhJZRNmUwni18Ffdd0ihVSaC7xAZdbRfScNUP60a7EKmp9KOwdjQ2BBC2pc0b
9OZEoQHEGYKubHqqRfcnP1f19DydT5gDyoIAUz4RbjgEXTtSMxvjFvX4T9AV1vNZhB6s8cIiMkbe
eXc2/0l+MSttxaDMGz54ivT778QC4BDoYMtcRlPiJQ8FS8CCPnMV/kw6Bgpiqtu42oTg/nio0GRG
6EMnIAdM81L51kuB4Oh79VRAd5WPR7oV2E3bWEE03U4PaV6lM0ExO2nCB0pn4++l1wXzs95+5sft
mmKFJikAm/CT9sqk7F2cIW0ex6dxeZNukC5XfBqg7D7YXw+d/9ZLRykQ6cgCDV/d3PbQ9Nulv1S8
htDL0TsjNhb7N/yJG3e6ddHp9gAdvXRnljLgYRdpqEdu3vmdcfJPrx8aTZreGBaUc1YoFK2Zsg/M
mpBNrv+kghF7+DgzR+rcFnKywGtvTu9SPTbo8vygb0ryB5ykO1shqsK+GPsDv55fJvJXixDbth+N
HzdtwjPAV07fdKAt9cZa5NEGWuB8Qc0OSV0iETI7i2QxZ86V7JtGZeQF9DZNEgl/Q4YV7bUYp9K/
OvIfVYHHfSDOXdw3uHNhAee7GgFoCXEOjLOTD2GQj3cdFctXgVTy5t8awhRl5TtL7BmUCSSHmEHK
MKIsnAxhoIpHPDHfbh4zDHyf3WkTh2S/m0InLE9NEv+aX7fqHpoHU5YFzsPcNx+GpgZRXXW11dId
kFA9LHPmp9P+eS0XJqkGhjnuHx4xPBRqOXk/h+FU1BM1j2+ge8ldR5jl88fBYVBVV/Kj7vwSInvP
rf/d6Dljbhi9uZBECkTXWmBUYvGmkRcf/JA/V8cNs2NDcHI/VtJXAk2kKp2H66nmKA0VTkh2ged0
VRsiIrVCyV2wxHL0AwXwmHAU2cSEd564+YFmpHfMJ/QAIJhjQW1mRDyPfKdE3p2kpgIViX4LS+aq
wrkRy7jbXRDFzDgr5ZredtR2ihG5LE0qBCDpx51OItQUT4hkYVcKCjv5OXnIm3WfWMKLhDiv+kcD
5ZqMMbiIpO8AL5sUxQLRkL+20AHywqDGYqMc0jW5DmHZbq6bn8TyFCIgxhPWSHGQUU5VSMjL/LnW
2xe4wtNZbtbkrar62BAQEfDwl3989mleRNJNgx0RA5akC8ZmLozdXxMW32q78IN3pLhUIfz+fmpP
nqx26UF88ZgSeSX2cgdrWZhAJCBTVG6nJzKOsOulS0R9FhqZqfVqgv+G66sRf0yC1jwEPfE1AbCq
s8jmYHN0VfSpkm/lcBw8YkUrN6Tc1iShiWleuPME3PAblLovfZW49I/zoX6iph23Xf4tOnXD9GKg
JXa1apRc2ggc/t+KMbnuAanRSZViFYkdibDgbZCv2kB7LvXtci3evaZ76x8GUzuLpRh/3f95bkWz
cMFQgHSDFVF0FfmMF9gYM48WzOI0C/MQ9JE14g93oRvTyiiBgn+A/w0lvj3zpoI9ZRLD7phdpIny
h2MkG55fNv0dwYXVgprCEGIrjNYXo/ZkNgDEerj/+wGJ2KRD2C3ununN/8Mf7E65Nt0xThD+ov11
5C1iGsvF7wBW4F9SGtYlW7MLPDIthe08/0kHSF0Y8CxYSUByOVGtkPiJX9equ8/kSg86vPD7+ju7
cISKXCUudAkDmyLw30wtAZolqGChZPv8ha2EY9zX0VkBXzAvtavpzVoIeyUbs5Co9v5CSuyVNlCD
CN65DO7NZxeGHC1hkDGuy/7MO5fJymzqrX69i6d3DpfMg69CCbHlCpQK2sdU2Q2fAQ57AiqMbmRH
oBt9pNRSQ7gM77HiJNHPKpF0pR+WrfFU+QPt8ngrD570uO7GTYWBRjaf8yM5tto0Xf41Fr9i+zBt
UxxUWobuMp8oy1aa/wcFl3Z27YuPq9MEBD/yjlQBRYAWgxMETloK+d6W6e4d7Nsaz5ZQi6wCJlQM
nSimg/is/2Wcy+5C/NyMVRGG3eKnYVWmx5f7pzHNYhSwnmhk49VoUKAjmuE+WB5K3fDMy7gqj4US
jelr7HyYhFd8FzoSi465eCuqzWUMuZjBzp5yvv3LczBxxv1910QSfG3vBFKlLZotSeMVIpasXpVe
tm9LD3NUzF6q2JMUlaKCXG1C1oLpVWGjn5Gj/h72NshvaLd/3/B9F8yikTnUhKdKU279KdwcYbB/
L4pu2Kc0afj07liUkR3zko8lLpVcyvpvVW4P42I2VnMrC4k+hgZKgs2/Lm3qUWIloEK+7GvByzaF
NNkiiZ52g9CHMSQNhk683fjHsehmsK2obUt1C841GdGEasgEV54KiMKyOqDRmq1ueM4Q828Y+6DS
VfjLNVLdvsIcbTxZDy8Bh4YLwkAlvph7EnhBP0mL3iY6RowmUibhKxstVHmqAv+KhdJJ86y2ATeN
XTudVAKPi/NHZ6Nujaedpixd2YQuz7MBfxgaSZjKQV7npdfN5gSyrVHzzt2QZqXDnhjsJcVnDWHA
SD8yBMxrEn+7gMMQryE1THjuD0+6c1aK+Lc8c+b43bERh/m5M96SaCrnmgjKd5s6Avmmgun9FgMH
3g5eESzDVtcRglqfxTXqybWcuR6DKqWWF61NGm8iphuX5SciCgsKriefj3ujfI51fwIlBp1eLBpq
OUa17F+utK8I8yAMEjlaqYSRCci5/pT+JG7mlXMr/7mOMV9bk2ehdhQdGMo7W8m5cer5ouneL6EX
AuQqCGx31OiT9uNyZ51tzuwt4qebWHFrM4LhKX9YWd+2RxDHOwjiSCo/CkTu/PATitEZDrC5h3Zj
Ygstw5Byo2nLv1mY7qCL9/rjH+EJInyIzV749lthDD1I4DQaB0+gelUIAO2xaEk0usQy/WXPQBUh
V8wMq3q3YVn7cQ1KjKHsLr8CpgT3Dk4Fwf1xAeEMF6PqGpl0wjeD4pwhtKxAsNmxqIj+O3jHE1zU
Qa0KbAmjhhAwGK9qGXoshRRcdXCX0eaB3PvtwbGbZTMjBWrFDOTAqx5X8jV0+YAvaEZyni+7DKZi
cuGj5jc1o7sHNQi7c+ppc+4OaNnd83o2l1leWm1dTFrebE7SvJjDzu7AZlhwKapVAxDl3NZvCWm1
GjHOlJpufXRGpsQBWRF3jT6JLsyupEKps42YmD7gq0bKrnqY5FRgxmM+jXP36nPp4w4xT3aAOvrG
AhMxgoA8oKtYRsTcaqp66Wg6oVcBx86HXbToZxC0bOKkjbf96s3eXSVSmTxP597i7geUFgGsMbHI
oPWjV4vkt2hsEIr0kGTHnxLU0G6ia15de+t6RMeXXk+idnN3oC7kWmy46ZZCJMtSwVfr2Eu0r8KD
HBL5wF//R5S9tQ2bRz0g3NBPPzHJIvE+qcqXaCk6ANpxqBmpGHtVEXGxW8neX4r981DiKl1tMFzC
L3LNKdlCs8MvXZ/QvmRQD++GL8uAb2cTfG13c3I7Ki4SZPmYq+DcNYcElLcUwDXWCNPQOBkNIpYt
1U3PoG6d35QoAK6GKfCHiayZUPx3gzLleWbeWXAoqR6r5bmjgMIvPdC5HLCqju9liwpVboWKKG2D
y1O7gOzQqnCL50mGu6lG0/VrtoCSjCBzf1y/E5QJa5Cu38zABH9He3IGuv7YVADApFnoi+VIXbfm
rIYkLBQhvjR1k1hyFdaSBw9w0+SgwxXuF86t1oMmjQeUA9GJFn9zkO8j7oetbFgx7kmFy+azGyDc
JVhe7gYfNlRcmQKgLt+ks2vgn6UtpXG1SKyl898nyODW88RER2xFJExV1Nkac04KEuI+MRbUZKJh
7mHVCcLTe0bRnfw2Dwi4sX8ocSqhO+P9BPiwZuCmz9ZdiYsnfJakr2rxTvGWLvdOx16rn51QSv1t
X/HK3CtY0dOV8ZQWXcHeCrEh4WXSItUOmBlLyaOh85+DHz402LAS4MLDByQJgbPrpP68HInlK+5l
rInLo7u8tijnLAwQB7k1zw0XMzooG7oJUY3AZDQlkQgmu3aGBI5wxcb2ayIlLfc3zsMx3+iohvJF
+YQHhOxar9JMwqpeKBoGquM9IFVWoeS6sx4Xf1dB6iTPOFgEby64JZQB/o3fZuSjFCVQQ+1DmyAy
DUvLEvJt08Ke2bxBjk2btDEYseZwefkZOVcgzrOdQSELv1HdAq2HCBZDFkdT2fBft+hW3VZyCMXm
VT1YblYBynAKR4CD/KfCi1V1r1BsSFDj5COSj1/q0rWJL8m3OHxUTAg3/MvAzmCCkct75t85158D
7EGFgmIVko/ITwUMfCc0IkWNkzA+tQtmyFyqQIM1M40dJt+xvN4bJWQO6zE4A+iHR8I7DnhNpPRq
1ZsvkJoseIjxpWnV7/eTmrKR9yRP65rtNehOwlNvxAcjbh7W7dmBhO3OvqEkvNwkptD8wnMSt+rA
tv2xlgGPnVx8mi+UWy7+FyAFTrw/2ierRZq6B0zU0l3HTlssycyM9b/CM93uXCb1fY6Ysz3EXa0Y
1gp1dFQhpzi8HiCgP2cO7mZT7qJaJ7+xwm43lSlvmY0NPi+/IYgbH/7/eT4QwmYQ3H++zDPBrtWh
DQ+E4hGwLKM7ftG9bfmDo/+AqC2DdDI+NCpz5qo2zkxs1XD2aG+Fc8V9z8XUf+J6/C5uQxOMOsoT
vYFitNKw9ZXQSwn+KlJb0EVIaooG76bIIM9MZ3UdJk+VdNBdRiehR4GJANF+Bo38aKnhSNbSmZ55
HnhQiuBh/qNJ0aTwrNd2Nbdgbt2IWQ4/pOTINtovqRrI5VWJqW2ROH+0mtf4MXti1gr3ehfvjfI8
6O4tflDkhE6k0OikIXHIqe1OmP3uNgWLfhNDcReY0Sz9tXXmyijKSGVndLK+npvWZlnfafIYtS5+
dkXvUvWbWFduLV3Et2Sb8jSHejQKnX7c+t+62G1W+fbjjTNNOF651pJE8yUdsHCVs8JvbwLahfuh
45Yq/LOyeFqp6vNI9G1XQubXBQZS2ggNXjUOifB8wJ4MoAyyZEWMvXOXj2RFATalFckuk7szJ15n
CP5OQPISfiPiC0/Zno38NiL4Aw+J3mK1tkU2iNqziLetMjK83O5YRFahJbbXmdjnfvxFxNvkOMd2
QMKzCuYOOAFwbDTGLXCTuCNbho0U/vfeIWmRa8Vo1kHAgxCOI+/nZMP4Hr/bb6xpwP2iXpvgv8k5
dpXO9VrCB7zwFao7E4R2DYx2rDhJLjtu1JDjE2gIJZEoLKF1nNId/+tKIxzEcaxlf8xq3Hv1KNSO
kDjEFdgKRstUpVx7aLW5vce3DJ/5Q3NcqMArZ+rCS6Pp4dCSJfYeTeMhXyzvjeduKUr1mgmYK/sB
M+C6rB6+x0jt7YAfH0dXdaepjuXUoaHxRb/lXDB0D/ct5YkdWh3fln+Ao+LH8KnytBvYkOAxFtZ2
raxun6csC8HHKV7md8/V0MRtxukJz52Mowd4sn6hdiaALDLjCI4MgT8c4pjq5wL5ZLe0XVG6sVaO
XPDQbumdIdY7aijOBwIhzTxff7lweDYNq04fmimQCDXWGxVR3BasvxOIirP13TEr4pdNETiFo/iH
HPLXpvN/zgCwZc7hNHYn/et6pwxoTmhEbDPCdjIjR/H961sDpQkdFHJO4+08swmc3jy9k0CM46UD
/fUk40d/P0PQ2QI3RScUK+eEIh9ORdNzDsDNorSuxbvztGHHV6AtxfteQgBFFzJjEdxIzhBs/07m
epH9GpwKHBcra4U4K0g6IhJQ3baNC7ASOqYNmUNBi8cBwkZz0dKkLN3LMoQ48TW03t5GB2djlZhp
MuOlpGLeBNtoz8SyDfG3dr6RMy9yOx6KExV/opZUHOnKdsBpt8R+seTMiw0j4cCdNupRlZ2OWqAY
MhZimt3d0H98GVY/QpW6l8FWcKph+G8MsB5On1LySbsFkNf9Gt+Fq3iWoi3uhUVLw03mQCCR46qQ
Q8K8oR3Ki/2wHKawqwqv2x0OH3hjALTvyZwW7TZjOPzjRIh7nzoIB5jLhXVP4UavjsBT1iSCVafc
R8JVuH2VkRY1LzROY4hYssKkeOuicOWXsDEQWTwSeRHql0V2YgjhctDgvf99196BSFv/8PMVUspN
JPhAYMM66c8I9E+LBwLSu0iQiNiWMdAiGUJKXT0ldQ4heNPhWU3dVhKMXH+g47imH7jx2O0kbsWb
1is7ZTxvDN99Hh6DzxtFy20+uimxOQ5bDrNtdEOSFOKTSquosq0jWK1c24JGfis3CREBG5djQKQ6
AKmtl5zBMfUUe8yeGurCoRSHHfmph7bEdSyabBwnVlHzkeWdi3BnOfzoYXNTiXmOYtxeqFPHsIM5
zD5eCgz2+VHp4r7zGX0ClSrEFv6hAzfH/JDwbt9IZ/eED036Jlp53saE27KLUcR35FSIHwCOTzZv
yVzFiblc3+1suVGqZQVJn7ZKR5HRq1EVkGSo1ryaa9XsL5cV4leOu/ts+vdLlY2z9ejFM0jBzsDw
7RolpHV3glwcdpgQYYwd2h30lwH/nxeHTPirBRaoakDGNHN72+XjUFCOqQgplFeJ7xgNAfOqYsAK
wMRJ2DZpRbeJ3iY0qGbFrtzYNCDjxwKEI0rEtGhf9ne6CqsjSa9IGW+mSfJJK7Ls7rRgXW6WG/Vk
DY3rrcCDvOyZNf7khdKw1lGXhOK73HxeySV+M31pNnnujgxjE23Nmvgykj0bfI6wNdmVOfVJZHf5
K70Gu/+LfepMsvEHCNL/c6ydPpwBczl+b54AD8sWF3L2H72Es0Ur9aJMd1XRiHHZNCogP59I8tHf
wkDEsbtaO7pzco65Jd6HDs9/q9oAFiJdANBDlnBpxWjdeb1f9nAj7CFWJQULH5uJCoHL89CYdAf4
3fmK8AAUsZTGDwKJgpZBCTkO2oXClLVnIm4hA+xwrfH0GBU3YmpH4WHG0/HUJ4sR45AtJbmyheOF
XX3Q11Ph1Rvo9eNAvWl7OdLAv/1nDNIs4NA9cW7Xj1eTS/FKStrtAtBodmlUO7PelSjfyZU2Pv3O
e7wmqbBQelVTX9JeOZ1B+VpT/YkxOyHRGJ9DUEI3W+3IVidDsHO2Q2QJkRmgh44eBpNMRwHBU9BG
Bd5Ey9pWCqm+Yr4AShps7UDeo/VLLIaEGS1kwcT0Hgtmx7AvoeTGT4CPATHBGB3ebcrPw7vZzO5U
s022tZMqwDLqRkQUzVxnZ6qML0t1g3HK/LsdFa4pdR9VGY2Soy+1N0nuh/AEJ79x7Xemat5QRjWc
6uaRJcTxGXEi69aYgL6hbNsNnXh3MPygfiM3qaqkkKxThb1Yx1mDTG6rsghaN7t7b7bHexARLEcZ
sAZl2STvvn0DEMP8mjdrYtldEZAHiJRj0jxVUXyxG3n74V706MNAnQ4UlkBLEQkSIKI/aOWXX62R
f7iqnC+VFp4mab8L0I4iX3M4kPTlpkiWRCUDH5qgjQ3cDGNsZUTcByYFYaxn/sl9FWoRkGimdhas
NIkv76joKEr6allMTxSL/z8GW2DhmtssAmrNdXxBkqOvMGpFgYKW5zQs9p9cEou8HztMowRkXkWg
VPw6JqnRwwuXOYuTs61VCgkcZiJdVPT1oMIs8uRDQZSiv7f3AGfEdGtz6hnkApXyMcrchpheBgkq
z50XtNeDVvIx6LXwWSPcETpOw/fkOUravHa99gkRrlzywEY9V/KhK5FONs41w3h9Vh7pzGoIbDeg
78oIul7bFqU2Z8eXxZ4y/WxGbgb/qorh+SknMw/Se9gqA0t3LYIZEZnUDyVReoSrYP3RO1npS+Ro
cPDO/is8OXKEsrpP+ltCGskkvaHC87rKLaIh1FStYDMGPOIh7TBoi+78KqXlc1CyMiCQZIzeFxBU
RiGZ4+0u0r9nYGrT4nBj74llCoEf2C5+pyVY3Bd/4AKS1ioMUvhsJXB+PQ35BxYzQmTHDkOg1XyW
RR17MSFGrTHdQN9Ut3os90X2WDOx3/aofBDSKyHE6scgx6/B0QWxQ9DBT6/61o81rkEmC9VfYhaG
gQY6VKhuZ+1QC+rfl0f6ik6vA48O6RWyfkG8XJXsXBOKK6XbA7bXWBnqs9xxepNsiY7WQSbjieUB
h5yHKIuq39ePUh55NXWe9065NumSh3bl+lYG+mi7Pzb5i5eLbFRbxu8+ONdOC1alqkPkHUGbreWN
cGCmso+ulwyk7cPaY1hxKne/kjgY1D/pB9cRXSxcWURwREYxYGAOvNVh6i3vC0ksljfInyjhsTHE
jgifvKra9+ZXT8n/U3lJ5w1okMi68ioGsONiqmkHuR7/BQdN7ZRjV/oweEDPtZXfBnEDCXWBksXN
T0+GqebmlYIYgHCbVf98gUKlHI56V9J7j84rem/jG3CZqwHIniPKOHF7l8YXUI3di+4q/WwkspvI
OLexYi7EkGUEZTq7iNb+9kNUTWTAD18gIGz1LT2Cex+f850xVeYKNe6h4zbLdSOSpBvXe3tQXbFK
ges0I6KGe41iUpZ5VSOfaULDUs0eNF8hw8kr8s5Al9ENhyD/Fl3yM6v7BQwmBkvxoTJtSY8ffOEy
OZlYauMeLC/GLga1YaurL3B/3r3y+DnY2nMy2mYZX8B7Ht44TKb4C3iwTfE1rLppHuYzu4nmpBm2
d5dKWE7dc9f+BEMOuUMOxtCvj9G5UY7lYOP5ePe8o6wdM0r1YyeTIqOWF9CkdZAPwirFx1TnV2L5
2nPLsxufKMeKvbxHIuz0wocZlOss3NJo19VOp/dDN8At3GSTha2ng8en2gNvdfShvjDcFgaMaRXB
eG2N0NYRrB3jKgtm82N2HyUxeuveQxEwA0IlMXxAOHByU9Eml+wnAQ+yQyp1r7fEvpzG9jJXkYFo
H5K7nLK3bgN+WDhJ+rolGHGC5CvENiJkhAIs5EHqBlhH16pWQTYkAaULLHMK1v5GSZ3bpzCqRv7T
u2o0Tt08Mmsmbu7JPLftY0MKqz3cq8i4X41yyqEf3rkSFCb4eqQSWRk+XYULjlCZ3ZLbbsxJoCOV
l+WqRgPmq6QCSydi3VXdo0H7yrZXIFZMQNG3I+5mla6LCwd3iS51VHTtSI1dZp9iJQNZ+I854Z0/
ioEpx43bYJJDr/7cAehLPtR1mW31d5+h+tQDyeIgKg/mXCubYmK6Ang4r8MoGpQGbg7tEvia5VNm
E1xpz1VBLVgPP5XZRzrofnmbnP1wPeAdJueaFHYiXUcUUD8Ja/YUB6QxQrDjN/oBeVn9JISjmtt4
N4/91ccsAC1wGhFXYa+/LUAQoShMnwtzaJVHm9g9jIDExV32+Bsqff///rhZTPfB5jzsgLImXGO/
ZLAL+3HcM3h2n0z37SWujajsq1u9o2Xlm7z5tWE6Z7kaHlJINCRd+aA1xZERLeCuCj5X+3bPDlJV
rfRdGWustF863OIMTPHlwBZKKpzDH8+wahPZ9OdypZmDtclH14WSeHDAYKr8LFONom3q8VgffYuP
LfeD9nI25ykdtJ0WTP2eaMetySQ/ZFYwEXtY2/DfrvUtfBZGdt6/mrdv98pXsGWDEs4rcAmUls4z
t6T0n/oJ0pOaM587R6wJD48CUb3QYI97barAM32fJhLA3+fMaRIqBnXp6VK7Uxaoz524A2/GOwHO
1VAeO29MB0KQGkYNkl7pbcLpS1tmT/6lvjgoF3jso5cRvE9L8Zr/sK5bjsFvHogVYV4ZAg3rQJFR
NHK7jCno0uLoRGTwBbWBjvVWZG3cwyLSX3vufaVqOmAmKyJA6DmeEJKupPTxZMNOQAPHhNkx+BCN
4ZvQqnwJ0LXV3Ha4RyCb7vv5gv8MCAB88gQXCBBuR4kbSDrPj+KALMMeV13mi+SOnUtM3OKSSKEt
FTrgV2BxmOTASur4A2IlZvq+CUIntPRBqT4wjBer7aHETjGsOaqyWmCfSFc99uyfAhLmeinfx5aw
oIUaPfcsMF8LTFEF6OT52c1JLkQpj60vYkNGir4kWAAZRy0p5Y99ctgupYHmpqlxRQgivlGpuKO/
qo8h6p88vMwmUR8JGSaS/HPfkm6JuWzCdxwfJVwA0n2actzBGz1uEohUrNnCJFF/taE4Bm6Qzb4D
auJzyqPBlmxghNyeVwQkQF+xy19zqZ2E06cbh4He76QFYYn17POVhieRvyLCnanTXqEVUehNjuaj
52ZBz8/jrrjBnZY7a0OcgVuNEPSXbuTD3LAvrxxRQmfkBV10/iZvgNpyP8xTs4LysZLxAwwzCKIS
42Cc/WkPqyfflqMFruyJu7cBGbKeFc/ZOOqkr8N/NqyFRIZdn75ghzNbGHcF89+23zoisanCxl0+
FNY/Cpvv+AAoCcIrQNCGWNukz1axnBCaN6DJzdcsf5vJ3VXn7R43h6OrzMu9eZBtO4LfBFZu+OwK
KQQhOmbWo9USZsmLKBKfLFuAnok/a/7KGVCenAATugO2sWCV5LF4xlVzJ+c6jwJ02iZ8Yqlg5vCg
eB31V7hWzEgLmZzxuuwls6LFo0Cv7DJ4TUbYLRlUdNUHUbN5YzFCU8ppzO++5RCdrq0sob4cgDne
8YDs4vFKbYaehjlbiUe7+atb2ndhO/a8tyd18kjRW8uh3S7cS4w66uzpj4kB6b4pnJZzD5arp8Np
aa1T+z9FldWiOb4A3eaL7uVCXmH5M3s5lj6LQjPYZ0znf7C/7BvsJvfZwu0TyVyGMejjPw65BpoI
7MISea/Gw8yddbZ4WQicxNUZvY2LxAvabg5qWwThaWa8/f4a634elnWrBk+tbEG7+fpwnzsuaa4D
hIzSUzW/Bi4IyV/FAJeKVKoZ9pVr1KLW/91I0L0kKXhPjTtBJ6Xsb31h0VqQeLp/JtZBJR1BVrDD
y+z6TvH9OL+8F5SLXLI1tOUloZjclPNGLyxFAlJDsIg675Gjc2KC0Z9S4ESzM6AXG/r7BL7SP1YF
2QLglCzKOye6ltrMXvVQYaS/ZpcdB+QeCqUANwWovV7gQhRrdBr+CTatFt9YceGMohlqgYCQZRAd
MmuQwKcKFGWAUfgWWWTC/yyj9lbAYTScKss2BaQOL9led4tqdeDhSV1ZF3/Kv0vEox6YZ95yteXS
kuEWsUydXEJliyL68rKtpvgeBSiJqdDNAEQxtJriTGZzDmZGcYc3jZp5j0H1lUwAaI5zTj/ZJIuh
wMlgTf70v+DHS7Pzpis30jXaAvDoAvl0jytyITrBNrGhivug5OvxElq55TP61PO/fE+BtzspPEAp
liks5nOP1ptogAAAnqlLZcdIjRrliiL4NtRcBIF8wE0ChVywRxeFlU7fAoCc1KIoGDq5LNePe7sf
XIMm77LMg7M6aQtngo8/IcR9w0AfupwKggxBlWhuv3oktSOBs46iZvxMP8FQuz0pDgutW7sn8W8g
Lu2S6RCoiLviKI73/a9k8eVonl3elGtsFh5e8+RJBEzSnxP5sguZTu0uWR+iymjvMxPjv8PQmxLN
XhoNzEa/hhdk/Zx5YpGQJW9NayieE63RINOqpW0DT/zoHggf5OnhEsTxRV5s6ipJQbUSZNU/Ts9r
XBhiV1R0EIQ6Mkasl7AfsSwT9TcQVSns74vyBjXAbApyvIeM+cohsRwxH9V396NzoChcbUFEvw9x
q99V17xWIjiVWtjObLr9TXzPo3jq/qnevLwbuhWiUaGfC3xzBA5RN0zk1zTjlD5ABKS9fnOR7l6p
QOZvwPhhoznABHx9C/4hi1IMlocQWiF6HOSfV1G1Eh//txQl3+p5MGD7w314MQF9IY8fNySnGyJb
0tWW60ghtdFxWtxaLsxdlnZgket0ZWlLO0AN+GZAXZmFcjtpj1vkGoFMXwPduACF8FCJxHwUbuqN
NpKzWe/gZv3ZPgi4ZIm0RN6Rl/+y2S1tcmaObNVOSdfAwXCWcxoLxkDQ9KUSRnjnypp462cSUO+s
TiQ+8dXsF9QhQFku0kENmO76XqX4cC9vgA8E1c4zViPKHdfTj79BHeDR+R4JMoVNPYXQX6dAY2KB
lzQVRm2nj/mfTKmVO2QAkwKsTTwfclWzpSOfcKFJ8G2+g1DU0VsVALdy21LzuHC2qIyLx1Ud55ag
7acl5zyjSgf4y8cAMIMkZA6+nsjj067YvgMUoqd4UPhXDafOCoTijN21Pc8emCP64fDcYmYv3u74
ZCDXAvOsGoDd7f1oCkABA2J4Z+htcENz4L9gzSXu5ZbkYTMNjZRfWiMTAJyh1CuippPSdcXQTpTt
m+uQlkWPZgkGn9JH65Di/qFu081lhEvFUT1cQVN0cCNlgrk299deN9PtBPeV9sdAjrMdCSXKFYIw
XzkPUhVED7VwwkKoqr7RuW/PWGzUQKm9VU3JDD0IJDiZGM+Pt3L8lJHhPDVUe/HA0GO7fYYU33nj
o0PKqZUp52hlyqwgOPJI6SgI2BHC0VC7mVSCXGclPrBsGFo4Ryy8QZGq1onQhymZo6nQTwjGd70t
Hy5RFLAO8tTU4pqC/4X0naVY2Bwupp1OZ8J0iKDQT6+sGfF2eYbxAIrBLEC3q2N03zlP+KZWk5Fy
AsmHgV9vvN3P6bYXUmNzTmALAWnUY50JZHN8laIZn9k8CvxmXHRRFXTZ0XYLbXXEQsESD0ePvwtL
Ctdb2Gg5AIndESaGqhgPu6HT68QvZrh3EZv/d1t+/2Q+U7n/5qwL/lDtu+gpRHBlV1/FOkZ5tRQD
az5cmU3ith+ZYh+1Kc/SOEEkKaJKDqqgDlIxKaK/ySluRS5PSjysDBMQRrbXPE8XToNJ9sWdbXmw
VsCAu/XqfIB/Y3JyMgChUUY8VznBHSKHz4kE8tVXGxQSp4Rbd6UMiUc7lQhuNPmBS4JoCLBC865S
fDH27Fx/fy9khAClacKSLz9Tq93Vswm8BZLbPxBXNEYv/mAuXmKYEn3ER0Z3uuaFZbIryUyaAReO
sqGeAydZ8tBaj8OPO9hEClF9290S9xePZJSPLTeGfOMCPGT1hJ/sA4MDz+FfCI91jVr9uDA0enRs
6S2dG9zH6U91wTm8ESPyy0ZKxGEzvznphnNcwWlw8/ctqgI9DnG1LEcn601gFn4wTVfxwBZ3dy2Q
Gwjb9hRRRJ/VYxzZ0jlk+qbm27HCIclcdT3gTliPv3vXsUfkrXMY4KtkF7YjMFrGwEVYcih/NXyJ
CE0zY1BJjNgulakioVNKzmzXBJs7tm8Dlm3bA5hTTDUP4yV6F3gtMEcDJqIiQf0eRpL5hVnOfqb/
bqZqGU1JQ3T1Slm3U9l/2dJn66R6wE/mBu6ff7ssAdaTn6hFSx1ayAekhqz3kNlx6r4sjcoHdBI8
IY8cjd9o2bS5Y7L7ITCwRiLcEWcV15r1t+iFWuPTM1DOsQLoCyqrDqCGazizapeXcOrbZZCFuJTc
6ULP5ui59uyvmaydUb0QLszU2mUmhYbECGKhKFdVRoyEvKriJ1qCil8ImSJuflYH3QVl2YSRbIiu
b/UmQOmpRHD0eQkDIGXkOGIlHSiyIehLtvisGPB03JAromG+m/PssuKsdvv1wdjmJ8kCUGjj3rYa
jTGBTEez4YzyBMLUwwseZI35dtn3yQgg6L27BBaBZ5k/wiVU/4x5eZ7R523U++x2T9fQi31dwUvo
X+jrB+yrI2AmkDZW1SNwJ7U2qaz4X3swbDeUhQ0VUAhBIakxe+6s+U1dLdevtrK2mLqdVpERVAE1
PWQcCIQgXGFUCA2my+k/9bTVn+TbcY+ERbVMt3a8RgDgcN2SCF4jQhd7QVZf5KZqq+DnwJDMlO5t
jaQA26zN3Mcsp1pCOoCgRFHPIcsnL6LD5yU6+bHMfdsveVsFv/WhSocxzvOUKTTxpChvGPMjHtsI
2dT4In61wCPLGD7hjAOhK3sr8dSqpusNq7CkeLrw1cQou166KE+dKzztqqIlKrn9DJjKgn2tOgzS
TlWSxGxixFd72Bx5C2/FCuM6J+QNUP6VMp68Ldm2f3BrGsH4ZQ+uPYypzHC2tx9lukRHZLWtVQ3t
g0Cm4zOV9a7ajTCI88Pcs2f8oL0yPllfJyJGpEK5vCPppK9pIIBFWCTyaziPBaBJoBSWpUPi/Lu0
Yg1kdQv4L77X/44OzY9A6sp2z8Lcou5eBUGTFqxdMFxQmEDQvPtFc5cURFiSmmyfwbkMQZs3FDuc
d6zYn2mYstm5S5zqznSDVjzY24UPHlXzAo2uhdmad4YiqNHmHKA4q8w5FbNRdePyV3Tj27I4LC/V
v13B3igXiYiYRdhZMcE9isa6Tveq8hzruLbFyBQoL2md9Y5JNKlDwREw1EFJ4vozfetrDR4RrbzK
oeYKRCToQ9WtpVcc3PKkWgD8jEu/xa1kZOCC2XVwJvTkkLhY6SYAkRYYg2cdbYFPETRLerkm0K0Y
sRZaVcgh8/q6L9K8v96DZubmmDJkqn8BB2xCU/dZIWK+bP8zRH9TfVmrEyxx24qinmMI/WuRAg5V
Cn+fh2Pc4DUC+2autT2nXXZbAiPqg35hPGA43NDD43FFfRwECdMng2ucGUVjHGYofYbfJeDQ5dcd
JuGBQFFo+gWhq0bYzVxbTaG4x/5+bGc6f5N5sIqhuChPM8jV74Gdvfc2ZSZEQLYVlgF2nZZIOySg
wnQl5p55E6N8DWOUCT3I1MisgeikeQvmLDLXdPtd346hq5pkRMfdykgiCWQm+V2vjzzLWpNKR5by
oKmnAQmQx8QIB7DuFOu580Z2HNQHU6DbE6EPSTqjIJXr+lhSXQuaZmgX83rsWU4Hqmjco3oAyAy6
WOVFdhfqkjqf2EYfNIggHGyrE8DcB09ZzNguiQWKy9z9UeHZXX+18WYa8B5CEtclNLUuYxMQaMrU
whxL41ZAnrhWDfpoW3EKCzjrwRnK0SGVSplkZJGs2/YIHGrpR9WiArlwMPTyOTY6AKuXov45iA9S
2QrgfLcVwnG3duP8K143HhAKAdd39YrVPr1dXmOPBrho2cye4YZXCBjxHQzz2Ub7FpuoVkMCog2h
4sKNrwi77Fyz8RRpvrKbk4EXBFkEJc2uvPlvjXPF+r10kKIo3rMpPGAr0yLYQS3eQIz2qR2ksxQr
iPPOV9zFESX47ymNm7wKPfRN4PZtltUwCYOh3vlQNuqbJhCPxMGliedL4BW2NKlHTmcE8Dw3I4+5
iZ+4T3uw6gJgcaQgfcFN+oX2Xn0UcNt1ItChHj5Ynl/ak6StseBUeEBTMh93Q3Tks+qQPgh8O2Hf
xZLMsJwr1eBMFptV3CDg54rybQFkKGUzzXIWfOaSzXdvXrLAyWzFK9UXDJ3orMV21KLt/ABrvvrj
JRIBhlhUbLCjfwV2rhEkcMtx24VC9PkW3moa4wmR7yrFwu6gdYmLGKb1MOzHhohUHO8kP3wz0UmQ
x64fBnOgdFNKUwzYuYbvac5R88C/J4QSM09CUHsZn06UTNzsGqLRByP91kLRM6TOm+Ob+ma/IEaS
QmBe29WqnEiXhPevWlPZKb49b24E9kwMp25Md5ZXG8374e+Sf9V6nQIDCTuAC96iuuLbeomuowcL
dVSvet0xv3oVsWl2imZkm8jUzwiWpLEygTqT+5n1BZsMjVYsyvD1lrl0uZp4LDTT4pFtB2GFWH9a
6JwEH7S+WOxZgj4vpDCWiDI/ABJquSQqV2LZmg7ImIH1oezf2WUl/OPmWLLY2xtmAFcxuM9H8mxc
tC7QxIJd6UAE0xXSHEBQnsbcCvDsii54uMe3b+unDTiDXl3e/WL4dAbgOrD/6NYLeUG6N5kC2IBJ
gK4CLKOYtAHor5hcFhO4T7NR9I0R7i9N/KVu9DjlrtAZf+U23OdCrJX8AYyzJKgJ0s2vCYyD7TFm
Ny9rcKXbV2QupLgophnsN2TYToC/cDXwEFhkOUacpgn2rmz/CPUz0/ib8zqxSqjM/y1RVvPfEzKM
C8ZDO7jiR8feHd2Q4bplusRHyDiucG06dz6AwjvOJSzqzj0bW6hRuTaZ3fzLOwnLACFLNw4kzpQU
0wzT4QdN5GQEWXFisItu6HQBIYI2SXmyL9gQwOFzKww21avDKZ7lPWT01Xo0uwkEWN1u8x+HpEKa
n9xOwqXBCk0zdbtuK02Vs290+OhIjFnjeWenoc4ndNKIOFqbWOPhsdgevvDf2bZWx5iI5X41acyf
p2v6KuCMQhI4alupLjRnUZycX1gxx6QySQubx880J9vIiVzz3D7yJibEvMKS8lyg+AZn3RufF+Hv
ti3wBUuPF+ctKvOZnThriIFFU491XMi1wr1oyLbw/lBmiOBdCg1FV+uY8avvuz85c3lyxMvp1+SU
bduDDy875nyjSYmG+/tBEpPCCUUp7TyaRKgTusOpbrJ2Lcxyv/TqDpPURWiKtN+ks1ni/dPfL4j1
hwjRu/pUhap/r6AkscLfaGyoNLEW+SQuyNyWoopTsNKRDyXMakdbvVPMdwO69DDq7MVGI1c5+SEd
6lWlFFenIJvI6e2k0vGXiZuBeInLUQ1gllIK1Qy873ZQJGosoWeSxlMxxZVUPfDy9tE5kr+mKp2S
kPfWXOTfOkAhIQ+18vFWy2DHiw9LicoZpyun9Z8ZAP43YeP3a8D+MXs7KSlhEM9JjsHO/mTZxGWa
YN868sMp/MEeUdkXaiQ4+Y9W5aaSudHqEr5uAlgRQAjbvjfNs0E+EKi37OTjHuY2TnGMgYyqhbkk
dONMI0CeKaXBZLz1bM0et2A+Ajw9+xPBARPkEkX65sgi1HqPTYxWqrqz52VeuZWRf+QsFFU2RVNu
HeDqsp8i/wPKEZy2sRCoBJOBKO6uarvyQCCeZ46Pn4Csau99oh7zlHdhPlCnfrx85wWjgzrSetTE
21kdEZ3Rbc+w1xOtL0dnaHPx/vr1Bq2zWNsvpIjyi2nNZh28uzSw0W91s4qubX1DEgIct6kvIXRd
X8NizJoE+E+Z84KKHf25npiRtTnpqlevSGYa28F9Ox0JKanNiq/b1oLwygTKLA7DPGfFRtj67knL
xrzKjTFlxNPa40sUX+FqcOXBbw+NeCBjzDysU6Heb38vOqJ/UeXTBt3UXyng/AwAzY0pLJI20b/2
JeyBW1gkWiU/C6x6+M5a9bqYrnDJIXEMny9nR/J3ny2fDYYKs8Sj84/bmegPYowHYpGP8UqHc5sY
Q4llOUQ8ycS6d2Bv28B003DLld1zIAy1rSfKQ5AKdPu5FCnPf+imuZoCjvPxGEbPGOimXx8Gq7Mt
qCQ5yBn41iBOFZlipPWMipKhrErKgwYmO3sNiWopxRskCdpQHGAuI4dU1iSLePFRqKfPOuR1lDqQ
1c+c/p+vz96BBdDaXUohlLZW0Zv0q/KgcWj5IJb+T24rKY09EJnNJTUYJNNZBWNGnAnBrW10CFrE
7RchOb8RN3eUbV6Jbyq3LnoK/iJBdxCXvBl6XaLheNm8qgdkr/qdr0cE/BarFO0DbmBwCq6FVYLp
FMcUON/y6mz5vTIC6LaNBHisqkMCH4SZKJJ+/pT0ZQYn2r6YDFyP/v1H33unC54Zgvq+DuVE/KyF
mVfQNPQR2tYhruBjH0sXmG+RMuHZDQb5kits3iKHICEsYz4/Lkg+RMyTjt/GGeEy+uKOe2c7QXI6
GaaXVLGZnUzOr4BmYAkJ2VdKizN9BnaZRnYnBDaWkqH8dgs6bagcrWRS5AOQFnYxRgoAYlJJJTwj
PJt5qO5pQA5R7jv8cxT+P0r+X8WKRxxLZmlhcoFawzQqoPJbtcmmgM1qRGKzqWFj6TKxnKpWMlE/
EIsG9i4k2rNxASUz1cy3zCjWnh9XT+h7vpPfvM/GULp/9+wEO8VSk6vgbvRebnCLKN5bnhV2/v4v
zJo5XRWyh28WBBYLf6H3G+I/G73n7a0RzWj23iSlfuGpBB1rAGxfHXgx7gxJ27gwnlWFHiuiFM7L
FaWEFIjtWj+tRZru0sVCJV7x+LciFhXmiHzyPbi+1wTUcPZLeR/eqasRNJgbmAmXKj9GIY6JZyM8
8vcvgG3GbhMIlX6owwqIMlyxe/Q0foYW0d96qh/IKLB2bXJc2oWH16p+WCz9Vm+JAj77kRHhftb6
vluoJeoEsh0fLmAqrfKTmnb9yeKBDA9wDebGNIctAgQ49TM8IlvFAcxKjgZhvvo31CEY6rDFPWMo
eUU7sJjer5w4U6R6klb2YpOGHazAkCXVwXXiy2DV4nWSApRhvc5yF64RBPRmGj1ozemaTe1hXxBP
UhUGM4dMzbfH+Sxc6cPUMNO6WiVeieVQIiIfMmbaEFMN0EKjVKB5hhhe9J9Qdzae9faIScNWvHJB
eefUyBcmMUm08rN6fANhze7xpuKABNxLNgbcSb6F5T8lsV2EDihc0rBXvvo8HDrTIm4E2XAqM8Rd
desnIHQeogrYPWcPjR/k90JuSOpeP104kI77YYiLhQsp8OWfOxcV3lf2LvNdqPqA6wwADuQPD1/m
N14l3lFXDhGS37bgLKgShRn2PRdFV13PtZ5+4yXTbL3dBiyW0NK6fSHAUYc9CZZq30QBQqTFbsbj
Q9EHW9AjvqYaHdxYUbGA7V60+F/Xzm0nsxohGyjQrbIJvrj0qFoMYpuBj2LqROi7qPuiv06dxdsO
UIne95L2a16BfYQtbvwvXHqsly7L+0yFDzA2zM6gxj57VWfNneZirfJfCd4Lsw0qejOn12D4lrmq
pm+lDQ+ZtnRHWICGRhb/6bneh5rETFunIEJcjYk0hN5bJ4jxwG4uZZs+zcOLg5sVKBPSZ0TUAmYq
1eFgeGqdiTz0mILOeb6b13FYr/3LVjh3BDmpxvlFyjFZ/HsogIUSdIQfPHbTJCftHWmee/stBd9u
ut6B3mQRl9F8P5Ec7l2Iz4fpatpp30KUB/b0IvVDmHE7x2335ctIAR3FU1Vn/8FZtwB6iL1LgLQ/
CawKmcXv7PPKuOm1VWIPu2ui6ZvKTJyqNRcvHp6l94tP11XK8Iospx8dY40teri4rlEtaj//a4+H
f8Pym0lDG7VmgCfOOaHhAA3oFlrWzsGszxi/XqlN/9slcuVyQmBT9q49RIz8VYmzAP2IKnk0bCEW
IjxKBWBHl4+0AVSYRoFZD4gZKWsKepaGg3cGTaIJXDbQzhtsDBAD1b/wG9N49dHtlzvFP+nnEdD8
LAphE7iJrG9soaWlukZKf6AqUkW2OD3MgYTVsshyehlju6jvaeUfhxilHuEuQVJNkuMzCPZ/dRso
ZLQXz1DG0jd/uUoYqGfj/AiwAWw136j0Z9p1zf1r+W9BvHuw5FuQUVuxjf8uFv+5azWfNZSwlrGR
59F7z/2GUvvYxp2B5liJLCxtOQ+Oep0R7ltogR3fbc3gwXNJmPH0w5rQvZjaIhYBJGmCyjVtlUo5
ZxwukpMI5h/R7UWv3isHZ+mWdZTQzZr311hOVTL7R+PZBT4zfo3expQw84np1hTdMYVGMpaMtrnD
+sgP31OnxL2jZe+QBdRrTjhgZiuttbLPFxLAnDNmMgc/olkz5+6c1AMEY4IilP/CkZXnQSzefJDb
9DglQB6ES2I1Hvw0jHQcpjDvdIxdHyEmV+2xY7FX5mvi7OF5JCR+z+4wDEnBJZ8DKWHFBJY7dCGP
e8ryFgFYiMllffwJSR2wGh6uuBa2neduhcl7yKQAABlhevl+BT3cDyMErmVJvJyb2zJEEMiEKEcJ
+ReccdQzEqIKXSOmDKghdAHst9ClAVtM3oENXeI3nk9jl9SknAm93sBqq4NlYxVSk7ppA3HPr9eH
cBofZRGPAXjGNiizGQhGI/kfKOekbgJDiroHCZiG56PHl9RttejwFTSaGdJYnLFc1bgm5Z3fux91
VLQuL/C34ncxYnlUV2ZAHjutnKUdD/iitV1wmWdMjgT8FZ+V/sg4C5bwiPBVSuuKDSm0XbxxtTAl
Z7jLITOJyo1xqdaMOFlbuC/3iOYh4QRzXGU7pQ+d4xfZddbHSTnbGP1jlKoLky5mLiSN9Vg7KK8J
RL3yvHyVHNzd5eJW883hmgdUQDggcahMZylxJlTn+i2KaLCddujfZ98OT/IOV2tvS0gtG9b7BFl2
UUUpr7K+A1PKR/xUCIq2drsqDR8wfqyHfa4xAAMFsoEgP7A81YXgqM6+Rk3ID+NDhWbI6yA91Zm+
smlDJNyFnUXHqq5sZwbtyCiKbYz170BtAh7g1Q8IYD3nnnwnC9hosItdr+iNSSqGXxapNzSbIGJm
qo2C+yU256mF/8SdOwNe8zy0K0OGvZ48Tvd6JeUpMU5ycnLWXbieXVX2KTG03XCdNc01QfhUKXIv
u1nNMsY26pdM6L+3mTtSE+i1sC5Z2joiMzreuicgRkqSMV4Sqx0lQOJMekE0nbKqoGBlT38IrzGM
OhZ4j1rjvm+AV2/Zxz6jwhO1XyLxAKI1Or6oYJCpSC5MuhCbv0eBU9+FJ0dS/mq/rl5TE3lHtDdI
Sww2YgpLrche1fIjT5kMkHucakxhu7fS3nKheQiZzjxo35M1uCeOz2PGaoR/xLvUibF7X1TZ1Zu4
V9NY9xfRSFyg2aLfDzET+dOvyVFmjwz+EHgZ9fJzTlgZmKlwrTx3Cnr/PclQ0CsvLf0oOwSlHsYq
ZW96KEAC051iWLgcVNYeHxhCkGkTTz6qfvPrrflesIOf0YAiHTetr0igBo64gMmJl6t2WP8td66F
di41Y/sNjZGvYm31JXg7NrxxFRmKqHAag3sCkVTjKC6aAd8qwTlyC5ojo4qVwoQkl6hDxSM71ON/
vWI1Ux/cNft3p2fk+qwfGGo8EtyPK4UY1EefK6azEFMUMM9pWi4KPbBRqrBLi9K8jDAErRr1iO28
KEz3BpGkREYL8bFPcUEu9gSgQEksL0eFRoORccslqMUOAdJPLlgjjLXtTkSDT8TIXnV+GHaIxwdT
rzUY5IvKSCg+P5+G2kkU6YDuG9d0YcRCS/HBqzPfQ6Zburee/dZEUrsZy+DEqGrelr4Tpus+pguk
aE4v6IkMLR/JtEZ568spV5VFXIlayR2Xa/MYMS84NvtgVZduXqxGUrX43kU3hHmxaoEC3xrJ13Nm
Eeb9hPjeObbW0I3zGlyl3l1hbYOgB/bFl7wDh5pI9DikQHXKrG0dJLmtSgoLOgKT6069MS+6hnhE
g0S/JidCtpXJj7I+KhaAFSR1Bxsn9DJmn3/D0QU9nXH/yyf7juZGtu8oLGJN7YtaIh7n+uzIZS3o
uSDduzb61x1yTMMVdhDRyBVIiSx1Eua8lxNqRDacBj7YLn48VP2h2HeNWPQbqCUwCCFHv4G0ud4G
8hXWjDNf+9iLMg/BGAd2pqsEZxZBWjJy08APz0HFUYMBn5KLHiabbqmechQ+s/+8dgepc4s3y22a
YEAcvjpmROobYk9mup+ayWUzkTZsVqaj8GK76dy/2ajDhTMErNtu4LJY4dj5EdP8QQBHOpzl7DMr
rEqCRA6N5OaAagjVLg+nk0RieXmkRNshr6R8bHgPYmEAEVQ2l8S3+OZKKN6o8oNw9UJcWEgxqGIF
f400ozdTHBYe+L5P1ZP+tOZpUHASQDzmTYQqy1z8zafSlQ8dVWYY/UTt0Tkj3kilbBomXLLqVZRP
iVyaZ9kX3BY/qIXE3nFQbyAMOJCK6R/5QSf2t+/23AIEIrhEMf8juK8eHE2WuCfHkxYu8UcbwEGf
0HIwYwBlIC2RctYmv1E1pQws/jb+UeOevblXy/27RW21VNk/juTXipSJThbvQY0b2CSA7oTqEpSj
hFu2td1B9kIqoMIH5hW/CnjGMymwIURlSsRGhTVgKF63MS76zH79gg2NIGxVeB4+YYybvUFpNvZq
CL/Ylv+osSsqxy92X+NURsEy5CTveD+BlX515ZoN9dy67TUTSbd6GYv6abYGAxP4KYhKsM2OJvFK
privd09w182BkxxaElOhtgixu5Nudi3NC4p+ZMnq0ZtGJ5AakeAP42DdvvxgsOspfI7K+PTg2/l/
2vu9zrH0vsJff8B1c4Xrz9B6kkfIFzQg142tiHodnOP03FOHlvMlwgf8K2qOHOQfHZWgyiZEnKTj
IWk06xEaTBMlKL8OF08SVLBmxhNplX/fLH1JZIU4uN5BxjKnO6VCjf88do8gEQqC3pxOsABx40AT
mnbue6Wi6stICkMe9/tofj3DN6uJB5n8JJLI9Etv88plBw3mIX8m/uAt/BWhOZEb9PEPt8BV3Y6x
4PW2wkQnudZGiagmB+NMxm3lc7O7b2u2o54cF4hssJj3GHNNLvfvwtMTZpUVED/gzBQZnUprsGyl
rtFh+S+SSC1Jv0kwOzEhYYTmk01WSI5poEQ3De0hdPvm3wdjiF24kVrEWsI7DG/GeML+o8yrWvFX
d1X+f7MuOp/vdHHNDoOrzlEuBQkqHapPpEFQChyI389Qv3XLULNTlJ4VviIXpCX8bhpg/sr1WQ43
kYHdHNUtPA28nNoRCjQOpq7jnBAM72Vzd5cUTS9U7cAquuA2x5WGPZd+yiE7orAp+V8ScCFCeus5
XGgylWbu2Brx7zGWcUnvGafkIoPwie/mLNl6lWDo38oc3ZSXfxhKg+ZGFMTAVzZE2x3Og8FdCJtp
H/SAyDAHQnYy4tLFTGii4TigsKyuXaYi6B+T3ZFm9n77gXbJUjtrUpj/oKpK0UKyQ/O6rkMGHrMo
IJ2kNrWTwhVfuDscp/tji8V/YPyE6DXTR+e0MmD2egh68GT9fJk9vbwebjeWG/FP3ujiGsFkKgcm
3zcQZspeI+9qw1rk6Lt7R6Va5LJovluh/EksDN+hEdZknp8PUKL7oPgJh2U80K1uXUI+UvPJje65
CW34phjzmOgxYUwBLCEgu8KdfR+FLTFkE/dhoMEFfR059ccF0EMxT7LyO4c6jvlAX3sfvBTIU0ja
787hPx8RGzWAv1qVG5BfGm2cv4TuitHlYBVbz1Cs7K1Zp76xtBbGfxaLBZv29s3uX8D+osuAYP4X
jZfV+RtjR3wZyNgrEHr8KD6IBOHval4b4XK4vCuhCGWcAlcjMKM/yLFjYpusV++nVOR9BKZUKPAo
d2Opld3Gchov14up1zwgHkbAWCQ+8PPB9NUTJ7VCMl4h0HcUvD94nC0Ye+t2tIA/cLIe8cR9hDmh
u+TwljFuFBSYR5loaEaBTICFEXQ00fg/mB/PIuzl9QLwkWnPxyB277cWZb24Qf6yr+zpVzYqjCQD
xJlhusKRAzHrhxF4rF+RdVAcNBiFQcqLDell9OQE8xVBlpgaSiSnvs+pyKCf91UDOr0z1MXlHydb
4b0FAETssy/osy4rBMgjaQTL98Kx180+XV4+sUSfkQIZQYv8dS//7p93A01sokmcvm3sOKdXQgrc
BNzok0b27s1ePrZA/9bW/U7NIvroqoNsR2evrZj1VnStLIwQoAl/Zx8i2flb9Vuvgw0XpuCX0Lx7
A4mNf0UpjcQgRjjXMkF0gX0xlha27nwRPG6Mg9gq5ZR/+KFCXDpX5YpfhOXMpeOa+FCPtuPjHR09
YPaKhHDyimaKFlIvRaBuLfHwXPyLUZ1k5gBJexMN6bNlZYmb2f+cs3NrwaB0LY1Joa+mIRirnjF3
o91Q+mjZ2SkKT4daSHyAECRosRKiUoczGTfI9JKvDv7lxNh5RubBNeXz8DeA88U5El3mjN+4wz9O
kwL/fjdLKAYmK5cIlxot0BhscX4zQveIto45z21j23bQrfQnUFllSee6DhSzOXWxMU40rHyhTV9N
Nim5h4p+nYCGK3zGtT19yibAryIyJ7qDcHWH1nAJh5Fy00LF8nClhf3cZYcufBcK3ard28b3W4hw
oWUjRiPNIyZwR5QCWY8fRn97B/Pv8dPm35HkT3XpsClrokqg7TeEIo66pe9fvQE0zMN7acHL+O1m
TwbQYLy7xCh/G8z3TZkPi50PcW7dUlccxT8o7lAONLdFjwsUnHHSivuTM82oaiBd6L3ZbGzSC+DL
7aBrwtLwyJi9xvq2JFS4aSjw9wm2AcVENMUrzl91fQYLjwrSQ6SGZFc19gvpUwSZ8PIE90YVqex5
87wWaFxIxlm9woAh7hZQGgH3VljcIVz5Z2Cpis5Mq1iDViyySOX8IRws7R/qESUnjZqhBN7THjak
rjlvHFSADYwz/n0QdC4GjyxXQuFa8qb0fkkbpIp6/E7D2hSOoW65lqwfaxy0kmJb8tu64FIOs1b9
91ynofAQHjEmWQaCv+eE5+Zf3lkq6xcmqhKLDD/WRPYXqxpmprLhKcwgLL0tZmQ4hb1cC3fk3Wyt
06eNJ/gNjn0mAprmgjubNbYeW+YxyD1LM+Jlt/wW3scTcTvq9e9VCiENgdSY35NN3KySDKDP/ZDX
V8KXRoCj2Nq6UdfyPajexSchhHH7Ke85tZX/e2bcZQB1yXGjIpdO75xZsfuFD6JbkKQBetmEitap
tG+BvHEy+sXIdXCkeyKpgdHLnMQOOgWXkAUakgpbQCtfrU6WmqWzShtVQmf2bADda/jdcQ2DRhbz
SK8sZ/mYsl61T2QC0GMw5Bzm9iWk9B0jIzPZDGP8VRVslmKm5YBXy+B+cVitQOoQISfoMPp09hA/
aF6D575dTrifbEn6Ix4i6ZOWRzf4WSiLdqOy2wJQuVk9LzTnaDUdht0NIPLgaX6wR4Ia6UwDuAz/
R/uL/GGaR5qFlxqh/gNOTCrVEiijvhxNTC/le/IUQokFLURf3G2Oef4022STetZT53F+JVmDcZJ9
0lSGTfPu+XDOZDx4KCTV1ZsdvIGle1JXQn6TfC6zCnrZU7eDUWcaTcyD11Bhcd1JddkFlSwp+jIF
7eOcPi+MkveuHUm2cxJoZr5FHHpyFpnIOGqNplb3Y4vvV7zdBCrEFBhDtJOfLTwwLSW1/8156uuY
8ssE2HX7ggpA+Bhi4C1iQPYyaxL5ReL2qxMeKMp/kgm7ksD56T9aMt35DgBWZcTjm7Kbai87SNz/
Dw6Gx+xaLQlN4UCn8rj3F8gOoFyA3mJtUXIqRryTDXdQ3J67HDNWhzVmUiD7u0f6VgPFBd5Kn8Qr
suzOW45EtCKAzHgPSlQf9vkHzX0t4jWGSdbNN+ANMy+/UbtHhiui34PVQwhmOkDzTDDQWwAvOxP/
+Tpb+JJ2uUGDD8UF5qprggK+afgrW4Eqwb5oX2hYmH1f4QwJpzmp6EtP1qC8msnXtWXylH1Zj09w
7G/+zYCtKirCRYstozbV5s+RsMKjBamkEWjgrsGffqF00bmpxfnDqTxEHHif1/ssZbetKkpIfLiI
7S1Gnn3SB9tbA937q+otdudaczbvTzVjFtTKQ+Tcgw4esa/8x3+zNXaDFlXaf5AYbgI+UUr40W0F
awhPq9WB/Xk9boJFF7tzPRO0WWK7ZVYqlOqxbH37yRq2F4yfH/uN7aOT6/EZHEVZPzDrjf+UGtuZ
LKrMITYzUvS7axE3sw7MQO7kg0o7K4VXsrbTMoS/Z/BVLIxaP9G+ybZzookwxcYyzHldr1RwtC5a
VR+336IJg5i27THNZjmWyj95vLYxBmUEyQq+XEH5tC9sMqXIyw/ppI9BZLHu93DIOHoNGNhbPns9
mSxJxEQthCWTsmAn5hWPQfEXlnYcEKvansRFIIKe3MCUpzF5OO6jOe/y1uYqMY4L6xEJr/SOzZNx
NhTH5UMLttpHRW0gwIbRNO1a40NU8Zr1bXZ+puiTLQIYFvFU5fFXMpHhQHhgXJ+coiZPmsnaRYMa
MB8/Ia8FUajEMxnjzcrsml+ycZKvP5Nh6A5IIahFdkyS7a2yb+hfFBjaRkK7wTHBhDVk1In7kp3y
gyXEcTHXA95aryMk83X50yG+R8Ime5WURQf4FmlfEJLFp77AC9CcfpCsRcEhwn9+pslOi0x4KPbC
KbIqFGdoIxSKxlpDSBf/8nyleAhMfGh1LaQyIjDGWtBs0zGHj3F+cJCiuQK4awRoDwuTWmYfXHph
Zvt6lzdhHjv2K6lKncpHMKOrl9XSoyb5seCKd9t140/dyQo4aeJ5co7uo4d/Tl9fu6fhIvvUYFbh
SYjivrgcL5GGZajs0lb/4IwAELPnnKNOSZUvsicYVh9PCVgIDFfn8e0Qfn1vQ+1K9T5c3UMEubCq
7VcgD7Pk3TOQDPytDnudM7+bIShGerc7Z21PVkz4KzwFrP8XsB4TZwvOlHRS4PNt5GWb3i7tNeRM
Jm6XGvwdobmodBJ4nBb10wffEy5GSqMXqEoLIwdjlNdDr/ZS6dnFu1JeRBo/VB+8IvjTaa0hGADC
sNeMo+5VT3Shxk45BcoJUfFtrXDPGANOCyCOWMRakmTWSp99NEhEZxAE7OXI8MPCXphkEh9lUxl/
mcU/nuT6573pQeNqMlVQlDxpC5RtLaonR4a4HrA+g5/ljuk2KeBk4vpBYxjeJBd5Vzi2TNS28QsO
kwnffDd3YPYbx5PZc+UaawhttT7uDJDCchjaRpnUBFzwWRPfxslXE2adWDYBVxC1YzjToNGLSc6v
f4juUrGu4Ehc8TME06djJahq7sy1oTFh/Gs0dgsTKFhwk0+zpq7Pv3aeifb6eEtstaYMbl65Nl84
FR1Wm13oswaxh3b/V0mmnEj87oVrSBT/YfaZWovkgtFcfzY1/5MAhb+2IB+hyF7U46OFoZm8HxOQ
WRgyez1IHNGpq8oaO+2fLadGYe9DUZxzFn0otigcE/4B7wB5gtm3ixi+ffny1yaXaEZNDGeL0khw
Ez3A+cww6p5sQwTzvBaS0dKbukHYowIyyeGYTQnStpTWhp8Ly4g3Ps7zG3CnSR2kgb9vew1q9LA5
A4E3J85vVqvLda7M7MpCDwFAnAkG5PdKPI0tyYhr/4DWKfKFBpxMFw4/68Q00W9aZvlrr5UdHvv7
lGPyeqG4BB8c2qvpPBBJSFJbjO0lRPkLpaF9ZOTsNnk3NJl2T0wdUXp+zOxms0liUVdh2JBgCtu4
bJI6XhNUeP6lHIsiVDvV9a6pTd6IDaq9DCtb/lCAqfDdTxinvvbeQuZjCsHWX7srj57y2xF83SPl
sUZzfsCNRr6GepwbVdwfkYfQo1Oj3csUh3LU7uS5FQZtklnZzqOrH2B/nDBP4iAGKavMZI3T6L46
QTIN2ZVoHWyD9cg6eK9sFiDP1nAz9CJxsRa4WgEXUH8O8GlhQRQg5tItseNtHEVUmkXRak3UoDBe
joDS5W3vzSxvlEA2hhhXWMcOQj2yhbZgb2Ygkn5v8kf5ptZK0mvqvY1qXB0THt0JzlorkyDbcJRP
YSBRMFMW/RqA5LYSE6IYtZmf7MGE+LiQeu1U4n1WOMorYQf3WGCGYiD5SeEqg0DPDn8Cw1eI2YjB
i5XHeVu0zo9IwlbZ4MQQ01hhGmKDK1IUrORCPvvYY0NIsvp5xqXhaRFYpe7AUnIzPst8RAH8svRZ
Dg7Nk90mC5WP3k5XbzlkUl3MXT1//GqWXbMOdrYvRTegwydirkO6iOv1eOxGNETJh/8mMgHwnCKJ
clI82NLxPAEcvasCwHwn4xIMIx+E0QKUKRG/eEQvOatoMFyGrAnr+/N7h2a6yzY/inTiYehc83lr
BfnMZ2fuD2Cka8VSBYjD2n196hHgwjh4ATNAXxfZt+XDq/G9u0Lh7T8dynq0m35S+/8S3tgoW+Db
67hZL2osmSFvZWkwZvZP0oRZ2q9zn8KL7doGMI7xzgFpcQ7XKWtDxsPwRkfRdHLSskZqbgMlTQxk
4x7tyAXsWmuZgvb4Cis8QXKilNPJg/7elsYTj/eg/wFU7jHr9YfLlK06I2b5aTFEcg8CohlEpoQy
u2QSMEKqW0QukEThnBxbLYoYS262n2AnYkskmrQA+BJ8BnI6DAdaWv4IGoO1WzPzJozQw+CKKN7b
GtcxUg/y0I6WiiWIPv16vp8J6fHg33wyWJSRdqXALT00krmfsVrQ4wWVYZW05ZL4HdUUwGlpociJ
pBGsZXb5yC7Bx1bAwP8oJVa2pz3DV6ij8hyVNeEjURDUCko/mABfsqPmG2kAFVPxt1gvdIG11Upq
rNIha7NScHRx1iComwO+cH/bFIxf6ojUJLWWgZpKYOUf0VwdKd+odP4HvEjSbIDrONi3GSQ6vSmx
jVJML26ME4z6rWqkZVOV3DgnXeej7HXCg6oARm9OZcAhHnG/r788E7M2S2pNWwzX+T2AOOigabJ+
j//0k6mZY6Del8tWQZzzMxKAZrO4eG4OJ5cBVMPl39x6AicdQBAFVgpAcYGB991GOuULB3Yyg0+h
EXAPrdzAbra4+AR8xXjuPa+wwbu8n4OO2tx9DE3QZhB+W25P6xFgnfQE7r7ec9GW6w9uPWKkw73A
deNZjUAWDnFjS2cO2y9r+ekMBQ8S3UnVcUPT81uulwkFd27b33X+0rDdW3mkY9yCUSefDMvsmFOA
pMjgeNXZhB12dJX4mhToGBP5jdxXAHZ2gVid+TmAf5fJZSiCd2i55gDWkvy//2gomTAGkXBa4eTM
FDe2A/srKsnHJjD7x6XSfEurzY9EkFW5kMNd3RgKFA7dKh46n1srbdTGrJqtBZRgoj7oPJvKbx4P
AIhUU9BRerYjn996BQ6CiJg7O19uYS3avQoq6pRmAGKiLTT/U+1TZXC8AYSZPl07Z2KXyjKmOefv
CvVWcqWBUjvWKNEnUVa6ZCbdDkB4XxCm/1TcZQbh9Z6H8JNzO3W53HjR4PEAy9Fyu3TN7dfvea2h
RyfCO+36zFKPaPbiEaVgAwLtJCK+CUMJbtxRQP8yJqp2OTKAxB6s+DfYwUMR11RpdkhCGBCwa2SB
ltTQXcUfJPHK3S7bMeo5amBM4RXT1+RWV4AhY2HcA0N9D9HIKgZPYwQsr/Rj9KX+HJUy7unCAX+f
QZ9ymjnLQ4DGBuu4mMZ+/tH3zN2qZNG4y1QzO6jE7mIxu1GOuy7D7X+FcLr/jkGLDmnTWibJhTbd
tL3dHkIcPHZJWF/ysnlwlMosmD76GHaXoMrqmy3bmsuvbm2grN7huBQRJfU2HjHOawieeAhWeVOO
h923YWYlIyX/V0avSPHyTKlea9FdnyVU5Lmd/WaXg8UXyr5Q7HZJ0NZEiun3mvFWWHthPaQIWyqg
Q36ZBUHma5pHUS/DrPzD1OUk4l83nB/jdj/BEWIpsaQ84Cd5fvc0sviAgGgbdab5mrR/DBL1/mft
TaZ7eQbO1fnk+pRs7D6W6AOtcXWg1EYjEz5xJIXtoiYX+wq6Y3EgUdTl0438KboSZk3OuYFiI7Pl
Dq6DO0UTWfHVQmgy5Uo48hCRDNov8XKEjjfabxzW/olQg6AJ3+rxzREeIuT6n98EEij3Ci/mXRTa
nG6ipzerc/bRfYThwifGWH/9ns4PqX5HVePqvpZ5B4QACEYwGk/w7lKInOw4eIWlehs8xCbX7lAS
o7FBePO+NOPt7uemdLi2RzKpQkvxIbAeY5ywx8ZYhNMLkyrz+BQBmtLrttZKeYgui3+foiGC8S/j
JRJqJFUCwj+FennZKLNYaZOxtHDdISLJXRDqOfR+J6rN63AXyHpPF2xca95RK9QaPVZMY+HVm/v7
MHK02dnwL77rPVfNhjCm5aZL4VV5gpSLK1FQBCoFuxRJrO5orsobCQ2SDQ0FCiysJMsAC9gogOcL
KU/sBJS5ZmDscC7blVu37hzs5/GKkOc/C+qLVE7CmTr5eYOPpd0iOfYriOTiA1wtA68UKMtQjBoN
mkE5IM8RpXzlNGNt5NxwdtCkjbyad8z7SnLuKgI8EEIg1L4x493TPt7pYvEBnqE4lUYA48xngAGw
PZOxw40eZSOFv90QvP8XI27Q8KK6OfEUSj7mXEt0y6RJ++DSYSPt6ZO5vjs8d23naZE9ico28WPh
k99jI5zoPJJlGzROZDUXIKfgp1HsxNduocdvmn1ICAxiZYG5GkEcgGEljX3O9lNLXR/KEpIaYJp+
MfHzcQqAInFpQSTLO/9OqLaw3aCtaFtmzNcnWIlw0K3xoqkWrfk4ofEH7UT0NuL3pUIjEMjzCXto
uy+QwPGlPTgFaDE0g0AO7CPWxZWbX4mhmZ/QkpS4MvExXE3Zge9ti8K2Za0ixXgZVZEtb+pVGP1Q
g75dLeKGYqW1A1ZEnhlKyfqHr3iTyr//fU5rIat6Ze76qzEmFrrY9+5z+76CZ7T984LVC4ebiL2W
VlTaSBXZUAaITPRKPPm7suJLZPj65MpH2PSBVD4pEi1qQetzraP64XjdAhMq4y+6aQ56/Qa2FamD
h7uWmViBwN3O/c7E/YUlDkKC5VWEe78yoGFkDsuux90ZyL7XR5n+RkswE6sl01VJ52MNkQOmDgTt
kIvp7B4sG7vi/hllulJcMhN/lQphauLgMAlY9Ef6GhPJAN8dSuT9/igRBIz46OJK0RDpfI6Jul80
e+CgpQHdZnApt6mPoAz9yMWvoiC8+8nSeFHtmaq29tw9Upiaws64jzfMIqpw5OegTt/vJZR7wHDi
cxYGZaJY/NIHWQsiLH7+jM1+YLOOOYFOlyfb+p4P9w3M/PO82HfyUazA5nDHSnwX+rQZ8ywePvlT
ihqIYaZwyy1ExMWKxVzPSFhhQGTKK8Zf1qqz0fFOLkxEITxMIL5bZ38m2NxZGvncGG+vfacLAtbp
AZpuzZlHM0mC8WRmJwkbD2S+jkWmxFjVmc85j76hN084lHkpktPqbMEaHAzRNsLVIJ/m8pev7SIo
v2tAmSJqQGyHkJ9xaraQYwP6Dti9GxHmeCLLJSWnnCZ4AcovCFszxdedyf+MEC/gnQBquyhE/q/j
CZdmkvt7HgulWvugMYN0duDXjtUVj+hV8hKmwdBL0J6ukUUxR59N4CfxeHyGe0zGZsidpOPXl/Qt
B5X9l6XdAFwmSlWFvMbb1sP6EcYrDEv+nZVqmNYavC7Rfh3WEsZWEaz908Q2h2FppCBdFfl+Z2s+
jmvcGHd/GaxIIV4jwOWHeiNG1Vu6UO1SzfbaLD+XfX98DRmR78fVf3G1YORrWnry43strfmiZAqP
ieFuk9nXeRKxBVmycwdUo/AMUV5XulqfFCTBmW0DSIWkTa5fc81EKXEH8l2ueEEq35gQoRxoWbct
9V4ZjKYOIUoZyYrfDWodZd4lPkc8mcOcDcDY7C0m6lZs7AHzXEzUyZK6XRr13fA2I6UYBUnAlSnA
Hzsk1myf/m67jrYNhFtBu41Vc5eKZNvt1ySk59BAgxkGufL8CrB4jWklmGuSO+h9mfLdkw22vJYm
FyhDEd5kDc7enlZSrIX1gq4p5EH/2m/gOlsIynI2We3Xy3gDDKzHK1Mti0TcJSciXrsTsOIY36qT
g8GyFnPxF1nPF665b5gmKYnkrOPi/ml25m/TyuFLD5ZlL8+KOLI6zHDa7Fmjggzo/DbiAguMXOdI
tw42trm0MIt62BXyrYYOThfiQN7Q9NI8UXVwlOPAGRK6fLX7jug5enf6ax1EOWGLCbGZbdtE9b6c
LdHMtUYazw6gGAmmDO2pFcx/HL65ErI3gOMArk92sgK1vlmVSdb64DUnBoUpr6/uoZtW2EUbnzY5
8y4UykfStXgSr1pTjx9eLaM7MNJu/Pz/jfjACz7JIaknAo61zXghryCodd2ASNNzQNf3WCRYBrjt
fc02zE5v/+y7IpTVGH560eEXtXQhg6+BQGMmhndj4UOo2xxivsaxWP7JBHM98UBqGG7rtPLg9vZm
QN/YfPXCp097egu/MssGPpkWV+OSn9GyluV2iRrKQE/ECnnm6d9LucF0WtPOaDtDUpuMGajY0+02
HWNSJSFdA5z3KMcXFV1xT4CiggkK/gt7LMD/zz8tDgfyrz41cQeCb5UNvzXBHhzptMTTTsymZxWA
dzs3TZnvOwg03rEFuaxhGYmQI/jN1XbvrXSoceAYpodqJ/2KI5tFLt/dpDMVccv7a4KOHG6+Dln8
6fKZWtgjBp8MckRqnSaLCdQaYVP1kE1imQAAN08wsDUNoWfhQZ5gYOugM/O+iQ4f5nHltRl+OG73
h68wFPXL9Nd/CiCn+OqDTmECxcWaMnWo+j0aGb8BybCHX2/olnzsQDftCJxUJrysIjD+/z/2pWAv
Xwmt3pAYmgmMAzmIfeXKWBGgtG3X8LulJxIiw+0aH6CHBdbm6laUoqeyhkHMuchYYh9/gWMI5C0V
4jlHsmT6E3WaCQ6kHtOd2bPFtS65CUqiY1dNx4rta/gaTZRDWrhZF+G3F0h0aytnpcRQifZl1r5J
bWr9trt+73jqGQvjEvmi3fo2wjePcn+hZLDmFZJUhu20mIe1TWDIlV1/RIV+LvBge2Pco0PAH3Bp
EGP1SiJcWrY0CR3B9VE8AvaRE2xQP0bi6NvbMfflQUFqLfiTK2A5aUCgfpET7PW6P5loNGAVMeYT
8C0nfxKEzjUyZkHKXSzwjBVA8qiUn9i2ekrYDme/PxH9aO0cgtTnaUfQOQc57mC+REKz24IwZTrC
jY2eSI5qJSvNQzbU+a3vgHxeA/dYlgjmEpxqMRwRtlNt2Hk9lET+59MJrKz7DD5SrWEv6AbXlT3C
goLQWi9p5CvqDDWCRdYOxSTUf9r6ir0be4uj39n0/pIonNOmJs6OxQKIKb71tGYSAobKZhqwCCrh
Wft1An0PcVDXmRirsnpZnMv+r79nbijQP93FsNnsb8LmoD8KbPOivMC2OyKhU6x9K5Q4IxbD0/TH
CGE1Bj7K2SBiw5e77Hq7hZD5ilrdB/MxJjAZV95PfvzPA+u8o13qmg1G2He7k2gWirei/9mXeNL7
qnpOm8HshfGk6K9whOjaoIfdPgQkhhPa7/C1ydWSXfg/xatw6UpTSRvS51l+hk3uGY8FuVrIpkSZ
DD2WU9HvMFqzaeBpIYUwy67+3aJ1rVC6/zxstph0fBAA8eqNhOen4joOBO9D+99MlNZ8jSQyAyON
sQD/pbuR8+2PaUpql+KdX3Q//8drPoftBjSnM8iofYtoGDFkgLgn04y3W2uJfykdfQMYQXrOoR8X
vB82n2FRkPe70vi+AI+ED9HYwIjHhrRFXtmsXLtZixut/L0gRrzA74W4SbL5hg2fu+t2GrzLehvt
1cCtbLhu7YTsgJIOuiRa3TeyXJB7zqBa6RYKtzpzdsc9dqYP4v0g5lnju39RRhbsRU7yTTPLE4AR
g2YILMo1uMJtLm9zAc5lNNl1NGdzg+xHWtgu5n/nr4cXRB8NHgk3fQ7ytqHcjNDVjPKk0zV30YHQ
1MpzhuYCpGHBi7Mm+gYe9T5TEWcu0muwk3kTTs6Y3SN/iUNmcJHwYREh6BJco+QoGhmV43Cv4ScL
9MCP8Nza6ECL5tcrUMBtIMi3tzXvjRDCqkZZ+Oly+buDek07Rah8SwTgnVMDw3F0ZQwIw+By55eM
z8+QspMtLvvOIDlJDqMIK6rFG09VLjF+pwfkq8KdVpxM/4LJTeJVfYCdTQRDlhDF8sVGUxG7Qhei
kgQu7z7G2/FNRa8go2ugfgQMyKWRTPd5Rh2TkLPasnpc1bgrjzXx5xhoRxwSm4hT+4L9SXHc/1oW
TrmY1vTXvjduxrYSWYY9oYfqsBxk5FNtBrtIjHczqucfjNK86R0FIZcBp5y4URfH0EbNVInXUXDr
ohfTweqhvBPaNZORpaIfvc9wro+aNIA3q2CQdJ8H63Zu9HRKF6Hts5gaNPfliHi7hJUECVjxAkW6
n4nKM8Qb1W3bVH6r2akxFqFc3TQT11tY18Y5Hy/2deQUx2FE6sT9h/i9DeutjO83TgqOOWmUSbET
FqKEC0gAGcjurRT/y9KzsiH5jflnhUlKfA9ROl6La3l6gvg91mLvb9MybDcAbhwadQYz8xx6za4q
XcnpgktUu/4IAaFUQYVLhjvCTtKE31N92wYLpygPq5ApckiAQzdKQEk7gogos/Un9tCRUfG5JJqQ
Rc09R/zjvsA1GHfEh8v+RA83k3rbKc+gJ1LhQx/jQX1Jla0YrFJSWPYRmWpQh1jvHUH7CiJyExOY
Hqr6waJPbfZILR68VTk3/Yqq2FTtAtPOOtoWQTIFoX2EvDt/EKWWVRkffXprVFqmudHCNMjW1hKX
Qfhp17P/LwdP0hbmncK5N1DNCk97Shc+/n7TAq9/xPJ6mZjmF13KoLsPSnE/sp9uWYVKxNTx5aI+
tgSIqLWgQfuJd7TOQasWB8daGD77ixqqY4wDBX2eyQWN1P0QgaeItMgMymQPQDPzrSxJO6FU2LCB
gs+CHTWnYWG4lPJQfWx39WBX4dAIN8Kn2BHnNNjOiWY/o4O3yHn+yiE+3212ZZwmwdefHEADfQlz
zea+KF74+2IA97qVmwawDoKJNMKiVGHnRN1fABlwwFurHPjeCIKTzH/Ws4d4bZXsqGYMxbCsWRZ2
Y6uyPaJn6yu3icnKPidPPkcl66Ib9BQ+G88MxhJifPzacxG/Tizu5L1NK9iCq2dWA7JK0Rq4oEbu
l1PKZzt+FcLXQv11r3cTCpMVBGdoavIg/D4PR+WAdtQ8t0Yw7oImwzRTGUUzzZvl2ywL1Ao9CXrX
CuUSqkYvc6v8tXG6TC/2gnr3wRpMmYaVk5oM3h3sbjPGKaOo7N9Aup1VHpUsfREfYtV7csx4hXqi
Aj2A9Gc2C0Q42q07PBYDakY/BWRPpMOkEXB/iMhQZe+ln+GeI3CXd2JsSVvee4rWaoOGhn+sa3of
eA1O2opfYg7uqtGuFTtaRT/e3g+27NtBFLrYS2Y+i5v8fEidYk5xEhD8qJHOsOdDS6OabeU9V1ml
yqh5bVRmx4q/sOOHyhci4IQBA1hIs/nqyd3BlE2wKGXlAF2W/cDaX5iITocdelNMUL5aMxKyOFZG
r0t8icXKupKvGqQdQtFGZ0gISCpmI1W5mh/aW55o8kd1uNHMwHn4wibhRFUfgdB7dn6c31rETYdP
njmmweV7mZn9LiM/yI3UF7TZuK2HsAFT4WVs99xDH+mV9KYIPgWD+FYEn0tYDvu99EL4gXnyREE+
wlz6MCVmHndarssHr8rSzU4ezlAzZ0aPU+bKiGw5lW9Hrlewcg25YC0p3bGAZ0xiKQL3m87s2QqI
ZAVOZYQui86CvdN4u5qCZI3LCZoZCVNMRJ+oDKO0CKZCFbK8eZZR/g7gKtril2+k/SCBqm0I32+H
HJgzQ3qxLWMCND4F34gvYCMutucPofG1ixsXSZxaPb81YLFzp60LYJVMdsAdtY3Jo++KIqJqxpQK
nwkErlMOJxDi/vWl9qb4024jNwQqx4FjBcvVDhB9MDhBkK3WqZuwPpdUDGyb0vpnanH5wpMG9vej
UemU+qza3BVkuDo69EI6fIAXD6lfrkl/6NX3Ak0kMgEUuiAIvRm8FkriSkrCvg+l3ep6mQPo8beO
HYxzymwZwKL12WhChQMhJrBLopRWq4N3sgnCa9pi2PvaaPKVAG/ikH83HTjlY8vurVtOCzuNX6tw
OBCiH4oDanddD342q4UDKQ5LCN6e3MWPQ9GMDBUi2xnCujTJ/2fB9bknmoANDVJFKPz2lO98uf7O
OZ/ta8WMm4jSDnky49WMy0hGEEf2jSzw1IcFpHv0R0Ar4XfyqPUbof90Zy3kwIiCbEHzd4ce+aD9
30RGd5LF4J3QLxBdYX658j0yjnTHTfoMc36OAdVGw17AjmghRAGKvTBsjr1noocwsV2QJXLO46zU
07geRdCldwlKmkbEMrdJiOAdCKq82MnoAZTKeL5FJ4aowzPkKfNrj99BC+U3K0C5c/zqSZucTEUn
wX8wmbm5rPHyEwgZkTGa6JipExSdAO1gq4h7FUwbNDU0DVIJrjr3XPUz5Z9cbNoMSqCGVvIzZLCs
3E8Mg1xa9mhHy18zARCnaIrTtFhjAjGPGao9Xhui5QK/pfEffr0LCK1glRdcQBkLtjn1irwUyOpo
Mbi8NOYd2FQoxJcdiJ22SZ4jhg4iXyVBbpEWMLeE44fOVkE9KWlaZApCBw+Y2eMzSp3GmvwKHpKS
pyu+Wn4mxtfD+aOndiM/KPWsVVtHDqIx/lmXvpuUKb1o3+M8iEHkhFVB+SKUg3FwNfsMBBVRQTZm
chb9iQmJkJLfiaQu6dXDPoX56sfhEXC7/2OrMpb+JznKFQvaX7B8Ceue8lsjC2f4ZvmlhEe8O1qj
IKixx8vmsvUWNgvBWjiCFvD1hUvsdGgdB8Q/Q7JD1ScAllP1sDqc7TPsTy/mkp50GG1KdOe6kFJo
bBYpiZCPBchmQ9NpL1tF2FW6FEESMSPJ3DH6bCgK8cFivikmMx06VXPQ7mrukCuZX31Hsx5vKFRi
1kfKiiSikIOB4Zh9t5ImmqDVn3VBi26wCmi/FDopaHyZyNW/XTn09ZKnUtnrjjE23xwoW3dM/vC4
4vFSTr8zxch2d9heegEMPWOKSZBn45jXvTnm3OqvYG1Wjr346sL6K2Zn++BbpDBNQGW0xZYaqQsY
deFKeuRibXFttg8GSk6UYyFaXCrqkaPgYVjMkuwo9reh70J2W6S0ah1dNMHanVXFvJ+AKX1O77kQ
39kv5lwTGrWbjFb1qJrU9YsE3++bdyvGEWWskEP9OcRKTOymIx4n6nxk/dUDaIi1AiARuqWDaJEC
aXqRwViNOvkktbdaltSrAPiS92uShEJn2e+3yGZHJSJhkYoomDLFfvmissi8tAwAnNrAH6nGpVil
LQx/bT6XMGhSpaYS6SUJJy+zQDTRDHrebXAGC0D/Nnys9lOxq3/UzV719JpcU5w49IzxBADZ+Kp0
ZcPCGLvW+CqjMquA4CdWOFaalDddP4TuAQE3y6umotXqbP1jYh8XBwp1UiupwVchzKoRFLbZ1tro
4NGQ75pE9d4zfb3/lKfNH+fKrC8awzGG/p2QU2FNGREUClKjMzrf0FvrdGVqySaB6FmPYnTQkR7V
uY2yqH7SIeu3bc9KiHe6lNTAQMtcbbNrDQYMKScaFQkkH6YvPAigs4WyOoDM+sX350xg7J2N+Opu
e6HVBft0x1GelXQapyVS8Uzii/n8XB53spx+RsX3TGyFfYK2Oe4COxNAAOfDqNLctaHlaqFTHsLf
Vm37kF1N9Q/o+L5t8Ji6aepL604nvMDgSM0wmQXIqpNYxtpu7elQ/btLZhnn3j+M8Ien5+93urcn
PJCoIqce7ChjMW6Szfh7jeWMf7m99ddoxho29agX3UxIyvjt1eAK2mq7jCiCqsVjAFYkdInSHJSD
HDbir/sIUZ/BTqfBwMX1LMXnKEvCUAJ/+TW/xVKp6bh6PMmXP6Sv0gx1zw8QKakN5yCl/PNMfe6z
3nCofJhteYwvRDZMzLlwIYLMqzYufxyOzLZSIfEopvFrg48ZwcHJkRbVJ95YThH0AQImCAu0NaLg
UDihlHjMeyeZ5KUwilzyzHOKu8WYxz8lvNtC7/NJ1M2/zNyBbFeRhjg9mDNYfq6RhoGQTGJYQeMp
wsEize/qREBXM1gi/UE3SkEnff8Z06SyJQV2kAsCuWCdy7yROy/obqutu6T21C57eAJkDIp1EnzG
4eq9PG5fRcbjLbZAOH2agfT1I8WXcyql/READRWepdb00OGl7seBd/xuyzHA8TGavG64S3InuTAI
2jLHFTn6H6M+nWEba83F0mcIUQvs9EOXiT++run6hDVQlkbH16nBIFXQzotUNZIQxDtVHTi+Novi
A6ls7yG03X3DxYFIYJ2cDan5+7m5lp37r/l9s2c3WZ0cEp8YOoHWXJEm8WjprbKaUFrB4njPR0Bd
qdmi2QFWoxWfLO6xfoVt1JE+oq6HC0dtc7C0S69fTZtSi/U2Dhni2GfvS1KvZG4P3+0dNJt0Scd9
VgH9ldlHhqfjzKFyAKaGqR/Hj+V8HSMt4OxRJd9Pon3+4tEeFg3tMJl7ZQ5fpbJ0RlljKx6ehmnF
Grh81eVeDjEMgLLUJ1wtITKdIQXcR6ZnfUdlVBqKUPDbPfAsv5F/IUiZcYMJW9r3kidYSHUfV9HU
Hf9OKobyLJNGmBXfucaCdjjRw5ZW1Kcw9QZZdgmZhmpuffN2/2IR3/DtzspBLwIaTsAvupe06IHJ
DPdqTAeimpLrcqzF4b7getW0mRAh5Myh74HMdTR757m75PeaHk2JXEF4Ci5VnC0P4hupFkNrTmsI
Wz4F7+v6pmQSn27W2u9qgfagJUR1NQh0tTcB568rlWxBt76i4Br9kf77enqtjMef2somS0QXMULl
Bfyn9H1aQGsJKKcgkQarJdJwSKte+FaPwjQTyjps+cRSkWKNNqvp1eH8WgKUEFTtNtb6U4n9JJfO
tvJI4+urkw28IPxh8IXxOKrv/umkF67WWacXTuKVdxN6A3DloPHDbWF7RpDFsO44cMTcF8EuKs7k
31BjsgiyPOa3F7QIW5EAv8s17GYAuEKGdEmyohPJH9sBA0vPWfC2YxTuQjoJuQXJTTAwxR6AMlMZ
k9fahSwqdsks/cJzXYiPuhARHK2GbU4rqII3UMM9OUlM1lM3AP4/NcHlVC2CtmR5q11i58w7OBVr
HpPH2bgksqHVft7K9VsdBGIU2HNk7cWBm6FboPmyaunTdlIWaNfFg86WqtzUPnF7XSkytmIL20Ct
QuuDD6Z/A9vtmcKORWeevPMFe7eo9+AB9tWBOeSDy90mLj5PWVneFRYKLdm4glMmvE93Hb/xO0QH
6pdTllYQNEkf5Mg1wqP6PZJVlno093OnIEC6g9x40/cyE5MimqXDXaIBvqJEOd6Zm4udjtNpU9JS
WoMARbKqXQA8kYnrMy8xwccb7xuc2lR2CvRIEuPlON+W9MtorWLou89XBvvMUXpOAWxaQMn+Yqom
BspANCFf+IF70LVWoA1ovGUxRTVhd4uzBUS0dW9kzSN05xqKhe16CYjGn/82qmHMgRZmlXL8Q0MO
e128PXXMGGQ/mCwbsjNZCC3gmDj2a0Olgnk3KLiX5hjL//nbJBeLKVSKNdJcGUL22GmZlsZvLj5S
E8JLPURRvEcTuWrtDphxlyfbHkxlAtlLmYkXSbvOIH3bOZVNEKNxGen7wldzC2TfoovGJdcN8blm
jGMHHZdphl1hrUFmB6SbrHQvHBI2hsiQ8ie2iBugFz6nppF7923b4AJDs9s4f3j6/PEhc+OQA0RX
QF1ox+15refRMlbPKwsqsiVZZncYxo/Qs9KEf1ApTP8oY+Ijjdl4zXyQCETxjlrJtxZV3neCtaJ+
76p7yrJywv2rnFkGK5V1eZ5xkZodZUlVw/SJbNAHfF+BTvyuQNRvCZra94nGh6d8XmqzVSiWD0zE
36pUp0nTGtPBR4od7Jatm2c1VuYCyPOxWIkqvm7SXNmXtlIdTpOXZQWW4IUxXC3xGGVTWkOMJ0CL
OFE3+A86txnzQdYq4WyOUvbxUSOyQYbHks/p97ksqip67SuCaUViClgtIe1X0DO2BqxM6mDrZGah
CS01RZ3Hb8icVDj6hGny+pV4zHklEDFE6U1vrQyEk8FFNvGlK1N15zDyFPyIBYEHNPjGOaKuEFbW
mrHkCByuAhy88GEoqXH4RQz+ocXx7v/J+wYVUqLXrTwJ9t2v9iqEnHl5Q/hM7Qd0uRyBFH882SK6
E2Rvf44E5eeiY/gHVqailSFm+DRBg0kHM5VVHUxqprN6HkaVcWtprMa42wQR7f45+M5NWE3eEilW
MD5FLAFW3sQqHDox3k9gJsSJJDubfHGoWBBbvGsk9rgNcoGgNkpDB6SXYLkOcTZGiCg9sBaBsaSx
rVvd+AdW8zeDAXX6aEipQacEk2tGV8fOXsakdRlvDQ9Jbf4cFcj0VNPcrkUBYFHJWH+y+UDCP4Lc
ANjipZtIxfFTg4HMl2KcemsmEnMFd0WwzCLdLgw+zx148jaWyCpLI3C/S3iWOKWIa5Iiq/RwPIB7
nkr8U9UOHJFnCJvSz3hcsirYea73pu7PZi03m6oESU0Hog4OC1Ph4XH2Q1H9TivTwI2QGzdX30EA
wRQip6Wb5aYR+acqpCcvONv5GCQ/4etZlNZKjjv5/q2+4WSw+/1U50OzZzI48IsAiJJSnQTASmoa
O5Rvmqwm0Hz67bfnod9H+mXmddTVjzWiDsCf7TssrM7cwrP9bVoA1jGCdjb6R3mZ0oYxBj7rOsHM
p4NcE93q4M8NoCcc//fxazSqTwoR0K14j+JNWtfRb0GcgK+rhKcG/N3E/XGwxVkLlaVxtSONE2UJ
7R1eHIaRZYjA9MUn3ajFp3rYpp1aYcoWgkD4hguDvQjopv7nQJAKakxd6lz28opnuBxX5uDinOOq
0ao5Dqp5QuWDLvS3bA69zE0oMXPtZEWZJUbTHEymKZxOuH4X0TEiyD1JDVmuBhXI+M+O/2x9Wx+E
L8XiTRRcG58PfD/5w+lYrIdAheqRBDllZzTC88sr1e8AouGPa4k/+hIea2JNuvAwJX0fomx7ijjr
XLxwDCJUXuOeBLFTEGV9VIa+Y2TFaLSCal70iTbmxDAgSEe07xyam4oQu4FnvcaCeHoh+ezRLoMJ
evh/GM2QJVHs/cv1CAx0k7CWvy/WnDhSNLWNTcUW2Rg5KfBeUERXcfRLoZQ1R/vs9POYbn9Txl2K
ANMCU/BhGq9QzCGL/QVQTFUC1zacoqDx3YmHHCBR1IePMsP6MJHU31gS+eAkt4f4XnQq6eUL0zPI
drDkUdrmoC8aBXlJ2IfHHpcjc+nBbfckKVDszly28KBJQHg84rIbH/7AwohEGSn1re4cgYfsinyj
Nk5pr+OQfG9D0GPvLhZxtpY2ViiqqWS56onk5ZHRuMan4KYQnkMjuf+HB9GvdiIe1B0PYn47WAhv
WxSCJF/FTUUdKdURpexgT6CMzfuJRnbTcMKNtdcUtVloN3/DKYSH+6IvALn/oms/EkcGQIk3t4GB
d0HwkGMH0KOTUFN7363GCDaZd2KQIbYe8C+61+Seu6JkBjY9yEKHeMSH9LHzLlgxhN6N1IKHKmnz
1ZsjB/RiYRgpyWroKx3qVDEasZG4DUo6TMMB+PVB0PqkRmcHafDYnDSF3nxph6osb8wVLThFM4Yc
oYvh1eei1x0wI+Dx2m39Uvs1JmUUD96OUTHYbzoWEC6dimfdOrh4tBR0cHk8A0zyJqjJlAKAuv7H
9venETFhstJNK/7Zzx+TVIgs2rUBqY4aSEut+cm8/jWxhp7TTnPYOuXVV0zsTbjcvMiPjcB3Xa96
/amDjBY+4p0lrlHwUAkilpZAL7Pl/sLrFldQOgGuNDLk9M/Te9vFifctSwdoNr30F6YJCCGGHKIB
ayFW5hEZ13iFAXqP/TdcwH3ZvPbi4urnmo+hK+rYAo0dsA7dzyK2ye2GpQyf8s1c3YbC1W9zjNSM
iPQn4aCeMcjUNwFySdQ65qPIF1o1G2VZtJXmA02rMyGEe23icsKjaBeI+LYshJGomvVvW6a8ro/d
HCU02VMJ7qPW4iKZImg381vfs7vfVVfE2r2YceEDYoC2hvhVEgxHUMSEzYofslvFZjfL7ck2TjQ3
txEVTsp+mItxDs/gmbVuSpBHr2VwLhcDQVsnR2ChNFJfTuhZLqQmGF0atZcu1OPK2JbiU2UQPN9+
37hWUL5cmDFrPf59S7tcSa7VSNkMo87PfRAAQbQ6STa/Xto3+DUVAmrtYFMQphUuE0Dgeyela6kT
OUV/A4ZUF24/vALx3DqsbEv2AORAABfJUcCMc7PSPFvCh3fVYe7gjbTakuJr6KjeH1dtZRXSOI7X
ZgnYfKYxDhcb1R9Yo4BAvUWjz3cOlmn1/iWNrg5AmCuct5xkrG3r0EgWPnWH0Lf1sYw1UqEumo5C
gRkKp5U0FxSUhyXfMiv7U7yeakkozgAnNcogWMDJmk7jBnhIJdyMBbFMbZois2OujlewVQyCKtSU
TT1tLQTK/yZpJ+Mxew/1vuRRybAEnDdk/7wuJNgLOFQbl+8Bs+JkmbXMQ0VTjdHO0VPNVlSyZO09
ORfJ/URc+cquNJCx/0VJWYLBE5fHThivIHd5ZLkB2xF42aWEAS1Pxvvx19DqjcMoEBOzffDLZII6
HMMFU93Ca2Bok9wvq1C5bfYgmxAP7+A2uA8uK6Hx7U0KBZ+xSdPTRN028UzfyxWpWq2lZ0g5CK35
IoXLgSQmrmM6Z2IQOPTGK7GZlK286WckIppZ2hLu1yoCTLHx6K4/2j4zLzisnFvJf5ndYco4FHiz
ZAIfpaBgP+sK9NzeKGeZJCuaHhb0fzD0/aaJChdHu9cDu8BCeBG21BId3kYDJmGppGVWtX2ogPcs
MXj6XGNlQch0pIu5YOaD9DRaY14nHPM329dKDYTOuqBMcdgtezQWJGfXrjtqqOZ3LFWlke9Ddd8x
n6T85lHtoOzSoc9KUcuyeLnR7/jKklqFnungcF6G3svZm5iTFCRfBPcxNBZh0vH/x8JYNlI4LD97
MORv6TR8m7zOWp+L8r24rww5ZzZM2kTD7CxZCYqBwtTLs1V0Y9pLsrKntIvgbHqVy+GOl9p1Ld0J
nYG5Y8ckT+CLbO83/cmnLIL7G35FSCJGKrz5FteGw9cZrXZRxCG+25CPixzKM4/pkqsjwqQ0M1G8
gF5ZlhtnxFukDagYMEUvPIJUARxooribODTSeNNn7SwzKVIIMaUpEHb/uTRDFZjRCd1Sp4KYMwV4
iuE7zjS6QEHg3l5sH8bVUOGIJjLdQs0x4/aCVmUF0LlWcVg2qFlqzoVuvXgZBGBBCVVbtBTUQ1Tf
3ZOyUZYYVUNDmdVFkYQoHVKLmBTCQOjOz9HR40D39GmYqBDWn7vxjF7YukE7ZYCesGMPHuaBJHi1
h6PO6X2leSBMYEZ2WSagx2W/llUOszX8sANnn+3AWzVdH2W37WA5XYSPZcxwPyHd7Ye2D596m76o
LTUTb0hVjG+huKSHJYwZYT50gP5s2/QN6DWF6Pwfa3rXxe8wHQLD4KY7xxfcNiszmFuw649hLLjY
6kH7nBIKAmInxk1zRVmB3gEtII9HZye9crc7/crn6IJBbjib3f1FiIpChy3qoVRWlnGHuc690req
JHj/OSfRk5QERZeX16OmSJGnFGuSvYlRCK7hf/reaOjfvaDk2ZisUeizKBGMpvLg9LE9V6g4DbgY
cIcaRRh85ktc1Hizvv6qg/jqvy7il8xj3wpQ4ZA+82hmqTOp+wmlZ3EKEkmx9fDeSvRejYVBhhXb
VnynMjMtJQlVBpxWLemWtXodbUf5nQ17clAz2UXAASmthOgPpxPM92OPwa6sAR119nBN8xpWgAbc
P6G7EQcMYWFnYeMLObIZUa8aydsYD+qTKBOX9++xSFD7ul2o3DD7nXFs0YGkYIbT9FYrqm8xCYSW
JeH60DXmuWuxdZuAETexcEdU4A5dBzVTZ1krwr2vVnwBT+Q02BKCCI97wGjePuQSz+QP5FV2Jn+9
5iN4YGLa/XQwfgPwDpwEtBdpPjl4kcSnkakjLH4Dpg9AA2o2hr/EwktxA54eX5iCzDf6/d7E22mR
h8XsrvoLxtWcHBef/j/ZcPM7rpbaKUTxNXgoeuoJRSPNhW3oYqyh8mNKXwGto8SmxTl6gqEgrn4h
rjEuKz9KZV0I3gYvNbH7RcB1mYsoQ/NspkZ6mGiVlMPOfy1J6GQtGCMzDtdAB3QsHw5ONSvn+P5L
728tJurvrcA1ixfGl8SmO/DcjPM5XlnV2koYIKIMKzk7QNcRu1z99t/JtYHgClaq6RX20RwBuycw
AQrLH8MejgrPrMtlCnUFrsn4lqnWqk6c9wxZd13Jt47sEmbfhnrzT84E4SDJOCMI7ihEOw+7eltW
eGndbD6Ew50NsJ4B5D1J5pcDKUYIu26rsZtxMOCw7dTF07DCoQJVM9PZj6GO6DfrALthVrGr3Vgk
KivBj/9gwPGKWsK8Q+OIXOSkJFjmfLjURs5qWDcXYU2I/BiGEPhi+a+EKhfFU9WsI9SI0Fctpcc+
t4M+aR+G46ccj6+Bsot0do2DyYzN3295xkVxb9lRWNYlF7o5syi5t33ueqtkFFJvd0UFu/+/zpYv
M54yUv/wG4SM5SX3G3q2R2u0PjLu8XlKjRf9f3z7gVDela6ke+M5HOIAhrVBl4yFXJ0pM4LiOu05
RrmI4dnEDeVBexuNGNwC0qxqUYa39VFrqCjcO3K5a5WjdTvleuKsTN+DMLNUbgofgBaAohhspVRZ
VyeZKIqPkapXH2frbhFnZuWIIxWmUr/WiEj/xpxafanc0F1acztom6yD4cfEOZJsiCqq3Flxifb+
Zr0edHDP7iMEhXeJju3RWZPN6aMVPodx+JwoH1eaA1UEdTFB9vdJSjlRfkQitAjrInRNs+4DckLT
Q51zVeXj8DrdFjibGahSYfJDqOddK2P78b1DJ7e+P9moYHYqMpGmVcoYFNSBFKlFXxYT0yTRngcs
QtLQ0YaBGBaLdTuaFklcLq5EDzgo71rGN9RdXrl82Ofni9/ZvoG5PseWjCt7X2ESkSpJLunplv6m
f07di/hItsNKubvMrRYH3JByJF68d/MZ61caasAKxhUPXdt3UK9M1iQiOiF4XTPPz/cqlovI8Uoo
ScTo/ggRsHrLqW+RcssZaG47D7RDAIxLQhTmgRpl+zTiulgWpmzDTMS9aJQxCZjMVUISvTNmQ5Ni
YffFnDoa1/sw5kqyywQx5+IkJof9e2dv4IZWOHlNe982165agP6ySoSbAz2ilefglrTMXTBEdKWn
mn4ZryDDuIv3t4OY0MHXByz3vx+Loqtpv0AANcQCFjkDevGxv+ehh/rJhXFdhWfVNCAiEvPSUFIY
gN85UXiM92yWmutmSrqOYfc5yo//atuWovQS0OROlZCj5JVYoF8HY/9at8P0vQ3Ckvw4qnP2cteQ
9+unTvGr9oTwkIEQuS6Cyr5V/l3a8qfbvsaVJuZHBiDmYS3Tfu+eFUbfz/0WYeBN+KroX8QCYwyH
R/jxOnWeuym/nP4DMWb3qslOMv6G1q6hKO05QXiwzddWtVzhTRUQ1KGCoqiDhAAJVgWjbScK5w34
5RsJKDDig8CRXmKit1vO4yHmV10hUD0WiC2xX7vqYJ3aie7FKdBNdaQTmTorM5t9glNADa3cRKol
r+DQ/gwjZVIx6qhjMt3L/t72+TrldeXfb+owmSEBvOTY5EuTM6G+ec77t0rKiIcxNKAFbTuWD5Nl
RIFvbcNLJzrreeEqafzhP+0eAiZlgJrFKt6QSWkCgcwJplA1rnpgmUjIgDOvVEYkj19QsaTx715x
ewDVVL8l9bjgEO4mXg2H8eH8lrgESEpfKSAIQaqbzhua4ePTKQgEmPQXCsnB7mu41nWP/xz23Z3j
dLJnlGIr0aL8rw7jJf5uqGVyQtMm3ihBRjlIBan6ub7+JYh78K++Y6OA2T6AWTjbC/b/IZ2lSUMj
3kWDGZRFj201tbOzeuGLRIz6rhzvpdV5CjqTy/Wu4sBLjC0avoK88MGJVYr539/VtKJpUyWSAarM
SJluUSNtlzEb7+AEnRTuQVpPETq/nH55PolJDk9Y80i3nH13PsyU1dROHTB/kufKx7rwCDbqn6ZI
POgOV2/WATIl+VF4PohfJ8bcRs5fmuCVSPIsoqsSy+5RNHarG1V8K/7hxdQMH5YnvkG6d1vY+Pcj
GywzWUjH2TKgE514fOdQ1NjQMHHn7bEr3rTSWIjY7+BfpR3YB/62BvBVzeFF+gv2I0i2TqpEuxZ1
p3zUt7zDVFk7CfjAbKjV+hCgPjKONbjIXetB5C7StXbr92bknoGZz9rRLU6f+9deYo+lrfX7mUCF
4xXG1XN8c3cJ+7wEeRBwO83Becma9YnwJEJ5qNTv3E4WlrQ1M6k3xgF4ZE4DBaWGVhVBAWaGoR2p
j++K3eHR1y3pLDAPOxtDu2DH8hfSopbREeypIp/ymVtDm2Upa2/3fqaNQL7IGKG2/0GKyYEFvf5k
jAwRBiRe5PAxina55Or3eoq6XFNp+X/BKtZa+CAOhXzE3+kL54Ss3AtGrTmMMDDMal+iUmYQxhqI
QJJWFHp3F7oHEB0ghWHnzqsGKzfUqaLtZCXeMwW0ar1zRfM4K0GkixOfIotww9ke4mMeNxRFfpvQ
1discX+Y495Bih0P8+O/IKiiRXT9D+SZ0tR5jL1QE0S00vJSlo2Z6ZfuFqY3dKmrg58q9grlyTi8
P1dLt/WA3pYES+NyiZOh5TnxeTq/m8ppeAjl+G3HIimChN85h5fk8w8wViejvW9U1AhR55yZku5n
Rq1HaYAX1TfQHQ73CWqf9l4e9oAGT+JFfzsQG2zD03QNDiYEsCjnsraojLOMZcw/Fd5o6Ehjsv5I
3uYSvQnY4cerzrFpgHqZwLBIBPhHy9AuRC6UEXT6GlesWrl58XvmvYFoq6mmanEYboV39FUQ9Q7I
6G1bygP8UgYqRexqzXx9LVMa+PJe3pSQLlHb6Pvbz3r93mpfR5BX2qaWupHhOyHoYD891Z1rkNWK
NkJr8AV4RfSPNx59aPJZ6OR86XRyb2leQakFtIVURei9rYWkXtGDkipKmmWj2G5qNP6kpvH+yK+D
v2Fhcd0Wd5YLGbfmLFl5pv9N/hgK0rY+l//mjqWcI9iNlX9j3QMUI9ReHxXSgnHrFYN2zz4D5Ufl
LTZItQtBxMloyOKzc0C08jKhMtRKbECP2RQAdcl4Z5gEORRMjUwEa24KmvJerRGuemwvwnS6x1yQ
CaIGMCULdP0I0NL9dRHkhKQs39OTk99BNzPiLEybTp5EO6rBGby2Xy9YSChZ6tw2vCslHEtS+n34
n3yn+1bBQoufOWtK+ReHtzYAdE66c29pZ2haDGSjpP1qvvqABrG6iHZYWxS5NyhMTVvK/0+3CDQp
MBknFg2Mcd2QqA4o6r8Fa6FQLVHihIOdu/v/hKGpPFFOJXjiG5/o75R2X4wLdzJDd+0Tu0aLiHbz
YGWEJeIuXAeL+7bvmptr0Z5K4fC/6yDzbFgqoQ8mffhDM1De8IPg0WWJAEhMWMVvkYIBydKvjEFV
NuatkrlQJQE3/kNQ6btpf7vgI51B4QWGyQF3DzeXCR6GZTPIp1tzuNWIUc2q9PYVAvVAeEDIH/Gf
vP8lUQOC6KkOTQ8GelQQt9AdCNNPTZJE/nggdORgZQkbru/8ggwW+lY16WYD3Mpryw6LK9g98kXN
JAbhv9NVHgkBz6GQ0Hb5pT0h82EQ/qbY1HWsKUFDcfMC53wy3WHnhVDet+LOP5TMcdhGs+bK1ftH
TSqXZD1A9J06czmYM7ilMaLiFCqGz+Bb18OIJog6lK6GE/kFwuiIMsfG8Efyp32/m3Nf4pvv4Qbj
T1Fg0J6bY/YLhj7eKJffUtp2q0QnJu985fXHXVO7EQAQ7suUBYh2SDZ7ZQrtFYniN1hJPXJal0W7
aEVIorj9XfBUb0srQGkLdR5/HyR44aJrh8WUMBKHQrbuxlNXsDIYwNXhuf9hGZ61xqFiR/S2ZPSB
46nHoyKukVzIz4E3KF0tcPl/Sx+YZT9b66Dnd3wYvtMtWPPpTiQRrnG9QjIv+6jHfO+2/ECrkM5a
+CQqlIvI7Z243N4KXLngfskW3uCUD9xTip9MyQHnTUwy05P0eNlG9Vmqthf1OPhOjnJi1WDU3sNv
zCMIaYm02FrtsyR4+aeqJl4Jg+XEszyddb/qygGacB+3YbdtGmJgIyrsMpKnvSSYj77q6Ssb28Te
QSG/neQL0x7kkhVC6aXGZnQ4XCx8GRy7/mR5151XDevUowVOo9WSI8z0S3kF5KGrvJBA6ZtLk0WE
V7ljjiV9GX2bUjOVbUI4ok0LOBcBuQfvfhcLNmDiDMAbPYJ/PCwsRHrxbKV1IlG3gVb6vvbm/p20
zTnwlM0pWMdQS5llzD7kKn8cAD3IXvjQYglqGt+gJfAH8OEerHwjW3YfGLPIvlqjU/HsoXdkUvTV
eQEzVpd0Td4QobM5raPRRKmZQp3Pjp5wG2R6eojnOVrjQdiR2TXkXXT6ATWSNe2aEM04z8iP04/w
zKdRZ0uvCgre7LOjrIr5CsEksFq5lAN9oMM79Qv9N8QiqhIzaWagcWzVCnEqHHmqnFCOvOvfcB/9
Z6PskvlC+uHQxz+KJwpQV1iInEK7dt+jIkGcxFM7eDLhlpr/q9POXqXBTx71yHyHgVWw8LTErSly
L8oik3EUV0O1AZKMs6GmSDs0F/X2UiJfrZTwwurCQyWU9yBjgP5sIZfZOFDo7nlO7masJHKDeOqo
PdYC7I8SZtgMHmN1Yd7WCadrkkqZHS3DZtAV7oRBdyRAB5rtITx6CRBbtvmT1eNnnN3at4EAJPqi
DWHUMEy72L0hJjcZ/2nGx8dtctHorJa6LPIaZDrE9S8uL9rEC7BVqvTwvWw+xQyak7a5s4uXvZOp
yvkGaHbS9/ArjqfpsNJ6EQsy7YnR+A9NBL0cX3SLUfx2G1gDIFK0n4HYUsVVV8eFrwq7xCB+xdjf
3N2WXY6ycSADj5HG3ER0yejitonXlkqOOQf1IogSEi9PPRpx+PTPP61r0G+i6JaIseT0heoxV0oY
OuNlpVajLmccTcbNPIQLyeS580GZb3kLhsMMZl0fHLlS16ZpcrLyXcfgKVAo8G/hI5A7SLF0rb04
CmNVJHdGKieypBNwkyB9blF0zxEhff0N/EonddUUEKlBcEc2uqGotQffh+Gxs7kFmrtkQmgMgrMq
eLJXtU0kSzXzK2ENAhTnT51lZ8kwsYOA8b0cMXyXkVq3od/8sw69GneiDKjFLfqEHxBvD4k+Rq8n
hSQENCLsWADzrUZmcBi/TM85baWSGM9Ip46znNChO6hIB+EPhcgzitOodyB+BU/ENsl4W9lLh39P
mpU3FDefpVsrL1kJqHWUzk5Tk5c6GIAbscg55ieBds74Zhr3RUEOID0Cp5bHuvMS8zXVslZssghi
IX9iaVaUXSlj6pxHOiS5MWVfdNZZQ0BI+c22TnqZ7A4a6qZNdXcUJdKWWVx3UzaebJzOBlLsLsj4
custlehr2dwWO5oTrHdNkONKbwQagHsZJP46iI+Y9NRGcxVz7/VEYyBVI+kWDP4KVksZ5rR4NbOa
rCWqNc/QeGPrjDkkBNxhw1WduPfENPly0g9fgFmyn6iNYp/rUqvXePcuqnam51bZgcmdDnfHY5Lt
GZ82xUmVc3Zn0kP5HvOAgpsmEamqLaqjPb0sWTbIGDEei9uLgl7MYac/hC/J3HH4mPjfPjz97zqr
jUsmXDnIT+G7U9tMiKSrKEdTVabLpbdesXebzdvdBwmZOy9i8MLaGvrlv36bT+X/3IBLFNGJkLM6
qY9f0KJAmSRQuFYsKSv0C4IVkGunVar0uye+AekooJ6SBHpGmYFy2GdKWdm36arC+/5TLs2MrDm1
QcR96bBjQ+LlZ90QfQno4+E6mNr4E2cNtOh4C93lARhMIhDsyuIDal++1RnzFfY3wFipyzGSL0XL
j0nldNK06oRLH0BgnAnfxqg9jjRm4vYa9qG9+ZRMY38Kh7xYqwjKc91kfcWOb24I1iN5KrILQFF7
fdebao1Yozo2YglZdIZafIMw1I2JNT0/ykhDKyV1TVrmqBJab27teYBn0bdRvKgKGv+tJ9ZC3DRN
nBgvHxJeXS65McHdfHuy+lc2ja9M845hgxqM842ffguMrUUtSSROlj+G3HB9KgOZT+t3qcfwkmTq
f1PSI+WC5cBCSacVWY+T2znFUeqzEq2DDcrdbTHtv7NeNlTbM+3HxE4cq21FGtQ9vdXmekkLR7Q+
Ro2fvQqRfKQ91wLQEvQ543wXybflQW23alAt79csHuYPwSrw4z2aCWRJDuvZBuDQ5w42xYApmj+a
SWlPapIAHoA6/Bgdtyk6Fhb7hKEbUHP1f8k8WFVeuTIYpkwt4oHyLxjORPoXl1TNhSoogJxjFAv+
mElOvehPu7jMcSKNmfUcXZoOYQvksn2RiMj+Xhq/Bmf8epHWzHrZeVVQv8Cl39gVopdnPxTV/WDn
d8/UzEAs7YbAddekuFCVKAjHps7+KWh2esZEvyrRu9ZhKEm9g6BGBG1yE9gI8HrGjzUEUySsYA3g
YhlbFXmg+lvRykFepyjYUvD2/DeVx3lmkyPa07MnP4kBalMGMr3XUcX2PkuR/0/eucrLiQNgdOwN
2/cg0N2Qkvx492qW9lw37bdYeqBeDlQnTKtGcIPNS0LiFaV9JCrPelWOLtQDrH6MyhQGcbFYXU7Z
GPQs6kjo8eq93jDwCfMdeIJa/MQjXQS5nzd9hWcDmHXCm1ITEiZbREc5cZgLxaw9dCuP6hKIlwqu
wVdMcAhV7A2/miIZZ1H5SmjrcCeOWdwb+hOrejoWrKvPIjKpcIkJeDh1Nwj7mFyoDBhcBirvAKws
hJC4ccvIwGsc43TetqE51QDgJJ3kq4U5MXPc2vHceZk6TWnVODgK87/w2trzQBvpp9dj6xXroh87
vbHuWB2luRJmxSa13FuukqeRIF51AAiffCNgIwDfPzn9OG6HbdniZb26Kh97ehSFg72H8rUnOaEC
/7+DaeYare9SHw+SZ7P3sh3yevszeQv17BsC9fvUrwOjgrxqRzNvYh7iAn+7VHQL92fB+GRiPOX+
QxfX/iz9cvAeNVmjoRy+0345/PJkgc0jl+USpdHMfBfP6B0UnXzHXHoew40XfI4k2Sf6WuPHIIPG
WWiKx9RUTSNdlNarnKww4n7kZ2ETBrLQ5vPSueNLGb/ogIIt8ueOLFfOawERnRGufcjOQfQXzRcB
k3Wd/giIRnkj31dfQuDMC57bNe8r8P0LwLs3hiLLXpK06x/ENbabPQTiVg1QOJg54BKRSGlLyflA
blPUV+xJ+GG2X4ynYL9RMaXNG2wLcTvbZu2CY+wWO0UeIqPVDcs12MI9s0NgJSsRJIASBfMPHifz
qNY0fwfzAw9YaFrLblTxBoFh+5uycSTP8QQZOoAnwg+X/dxsixtK36VmrpzY8lt/AbtotKerBzEi
02UgFSRb+9khq3VdTSBLaBVFpk402WPy3VtvY0F+ln/T/iDuG8Bs1+x6BK6E+G7OOXa+v8CpXg7L
zQTP0kECimNcQNvA32qzxOWBrhz+4A47xB8X1FN3UZeg/xU7DIcaK3tEzGfRGsokuUynVW/0qD4u
Ew14kZzjfBmGOVoOwB7uGp8Y8Dz3Ln9J1sOjY5FEI7lBrNxCqbLgiPXdKF1TAPc1D3KqdHU62W9m
0cyYNmcIY5CHLuB823o4XzSAHKrLyqMa7c0t/6D3srdzW+MayT4iH34Fw0bbDQcfkXlDirvpO/UP
einEorgWdap6xNHekFUSakdn3pLeK/kuQJGLZBn7DPLJjIRn9IIu/QXdtuTv1quqADMgf7xpyADa
rV5oykiCGIc8gxhQs/Q2dcpYLDApjr5/yzYpV6f7aOhx8LfJGlYxLzUHS3P1uCaX7xoMkUNcD+AL
jfgcXxuq0RR2AKhxsfGE2nSC6kpWjSY9891xeezWNtHkbASoIxDLhhFOPhBUV+1NC6DssDZ4jfHo
vlnGTUOEorUZq7w00xj++LXWUMo8UmXIiKYenFYaTiuMoappyDc9ydVgaH27EbtJaNPb5A9oDFLQ
zgLeKxiJZ8dig418f8NroIzKEH0N0HPTu3VWgufYZ88guWc5Xw+Y2TPJP+nj6nMSATFdDBtHzSYp
uKOjvHZx9YoNm12SS5QncbyE4WK1u0rPABcLZZXo3Ao0AA+WnIsplSExBGO9xWoJ6YSylSMHesQd
razdNYp1YPtG+zT3lJcf2GTPvkur7MCI8uHrqQ/EIdAorz7rRvBObq6s77Z7T67jFp7PZ30/TRxf
IoRlWQ7f84EEx7IBmXWERx3FFzQWJSBUKT6k3zGIHq5OfMRhZMqp4120JdN+tNvnkaa7IyzSQ9Xl
6BQl09iR5kG1ALiupG2OdTqiCS6GoHZ1mscLDnyz2ZkNzMy/X1Vl2mHIDvy8Te2ryAECeXE5pFgh
1FZ6t9kuC7l9t20mdMaA2iMT3GYzs1rt6B/ppWb8ujLCsOEhnv8SXeOIjfdOEwmtdfMy7Ff3ADvs
W3qUgEbfmlYRmh2wUuibDCObaDuRZppz7Jkeyzc+Ro8PEvN9ZryrPsyrR10WSL2b93sa8gQETAB0
8fwEnXK3pp0xZhyfjhLbeFHRuTQ15xSArq7nd5pjVl+8rdlg2CFlgPQ9jyu9Nc8R/9YPEJG/Waks
VJADUlD9yBIQyXLLdoIz/Auqt86de0T8YRTJBl+JNOm9fOqrb11+28s43dfY6aSJqLvl/4AaHty0
o7HJpkxp5FT9dlInCRsZqoaGMOji+CiPkCHwA56afR5EstuzpS78uKAMgrpsl7Eg51gpDT3BZm+o
Jec0mmNk+PyF21f0PJ1DjChpYnvoudCdbv/8aW95nLlRow0EQHtAjugm6od3cQQhGVUOL9ZS+qWn
MGwFiOKRzxVsH8D2AZgqpjt9vUmeqaoquZOddaO44bmqiL1Ntx7GGSzNf/i+iz6jrGd5rBLnTd4F
b/OU6jR8tcav24S1Aez3eHfV4rGPIGsrNUlBMrO6AhKkJwWcDuCojL9U/N2FiXDIDwAFCLCAWL6V
nu/ck/GYJqCtghaK2cOJWgFax55U1EqaotnshZTjomFBzH+rNE8HDLzWdptnJtO2BEz9//8AoSMP
TPs8RRJW1TE0lkDQhAaB0P93B0vqf+r69YAPhvHuap9z1//RDVmC/3QGeX8l0gTX/kdtpNv2Nqr1
AOwMRG+Wi3cq/6AakhKk3KrgVgJRNsLFt8SJAudd6yRBsQu2N8ag3ZXNfiYbCS7uWZBOAUdsZWGQ
BLOY2oO0XduTEPrNe/cgk94y4WtZSlPJzVzDv+aL69kZzJUqn+P6f9ktkDKTwmDcqiC5WrOqlJMm
qWTbVlUsLM8/dN5pzGzbW/9KvrctwWWZJ1yBzEcMUCJfHbGGuc5OjWU5HZU3Hqqvm5W7EKlwBSkv
EmNPq/jAaCrme0VoMkyizOVY8C/whiFjFSyWcNDoyLC7upt3m+Pe6XJpPjPhiKxtKdfWTksFbpcn
S2XJ8nfDiYZ6762Dlmxwy5RAVM7PXYl8e89SHK70kcPiiuAS23zxNfGr8XCwWmaV0ZZI+VriKSev
yP8gB9a9HsrBHRDbMBegZ4pfzsVZTJ90QgQQn697XV1l2d6ofDNBDEbYBSeiTosKOLuFQWZzzwwg
NGSlzWprkNqTfpCvDbvpMjgUtl4zGU36zAuvmXT0aOtqVg3OS0I/rBdurrimUcfHO4BoH7Bplafe
kDjdsuOFNQDNjVIrB87MqVrXkiuF1tkj/pD8f/nw3jD+kUeYmI76NJnAnM2ZXIZmm12xDScjdqzc
qPHPaWOrb/DyJyt7ahD9Rnvn/W9D8MbXmYcoeicEj15cAxstk5CbHhr9K/oBxNNoVg3W1O+zM0tO
qSlESniXPfAPOMoKtKrgIu4zvdis/a8jdPK3OJDDzhVC1yyYCNrYGu8OrCrCb4BkekUKl62Ho7mJ
fmWQO4Ak7APdKiN0Ls7OaXpuJjwww4BwrC5egmZlZ2Ciy/uJ8FlClX80SIGAp16LH2C+DPq+hGYN
3a/js4kYITL1NwbO1eQeW0xflnh/zd9+QBEw3Nwn4ueqNrGP3bbv0EHGbybLhRt8ImHJuoHUw8r9
bfJ8D1AOz3KlWhKH0enuNxKsPt9bm2Rf8YzPcfsp3NdlXH0nLLLDpnYAaMuoN92LNxzlGtl/Q79U
O7CbDjGBJlZ+GiPz6kIAvWG6wBn/IBoJt3Ml0NP4cMF1FOoEwwQ7bQjdrIWOUTkKplrOLoIpUuLd
bvm0/efMIi7xE9WCS5CCYUkBsbYrPmaBsXuCvkROZTxjoaZ4gMKmupGYvl/3AnKCepnKjAnuutc6
dFHdwANjSbg1VKQbFoaD3SRhrn3UGAH/Hn+hUsh/sFksa0YzJpXb98UGZEAwi5JVEVcFXK8vHhan
SxmHvBg/OuNGCQRXEWfOHkwjCigdP2nZPLAftnD6XynErfRSQPTtN7I1mAv50vxC5hg4g0NWLHEP
7bOkg+OSxpM5VXN0JDGwrYWswIlzsrtvgXOIn85IR0ScsawzTPAEaYdrm6oGqTsJSqaQxaoYurQ1
BmKsC0FT7F1QATwgrmJvVzWaVVsMUt+BlxR16oXSm++Hw92MA2Bc4I54xhO0YlJurnr5wyaSQjYn
dEmp57Vfv1U6otw8kLOFeA/eV/QC617EiTZKAyBt3lRhGYzh5HzYSnpLO4wPBZG+uJsl9SIkRjqu
sZAjCaNaJDT6bK2VVDtVjK9aTr+ehpLZ1BViKcxf6Ls/m65NbU5b1TSxvmGSrq0D2oYBgKMVrRMD
MwMf3oQ7gJ6hdSvcWDxZoYIitnlM9fqnfovWr69uZkOFr+mXEOLrlDWuKoR/Rk8FC91oQWKO4k3/
wW9z3AJ7huaCPIULuca3w3NUqe+PLm9k8ar+NQtQYGSqSfphzYxJxmCFCBL9eYcD8dffb1tF7fOI
tgOtzSW7glckjO6z/beaWEwci3pLHxSeR5VRca3sczbJo3CCReP3kumWkpLv5255618JujFVAUTY
FkgW6yYerQKjSkCLdYP0ByVlByfb4C4E3w34Q9jfjNX1PgJP5fbrNrlnUTtDtOBhCDykHO5M+sdo
1ckFwgSKFYsSds2+dhUY+KQRm6IdsUNN8qI9aLVwzCPemBiExJlVQlkOrbrbqAb1GCmmkNgno1Cz
pCttaLJQJDz/k5t9uqYSXWUjK0APxfpTuW99rSrNNmzSJ55E95itB59H1Cf+y1r3wRhdb2xxgiiX
UeW210UM4aZVkVsRy/hFqI6ETqmizS9u4jTsB8NoxAjPEBk1N89im6W5e29eQJcK0f2bNLDjRslc
VNVEGCnWJa+DFLDMOKVki3W6MoJmj0s02uwweaOUJo4WVe9dlBqp+GbsbPiP9NfgtsI0gRWcYAIh
QkYtj0JnQgq2/otcQddMH9Ydte/s75KnaImOajmxgwftfEgTdl7i/qGSrnutW3FK42LMaVX+Igqy
6VjQd7HX8MUlzEqdeG9cIQHFsOI+fRwDPMkLAhY6SZ6X+NWrV9HtFg2z9RCfJF5y9gtCwQKry9BT
XUFyHND149ul1Knhlkcp8G5htRX3g/KxCoKPhrNuQmco2jQNO8pPFRlQtCVk2Z78apZyfrqhVk9Q
7GmklUX+svuqjhjbeNdyGHH8+r/Qan+RbeF5IEgCbl6a4Gc9PJ7eXo3fE1zsnieCFhJedgoIq/SR
DLO514QhBsqbOVxPaJTwADc1HrzU4T3ybtYw4H4w2HdHKSfIxRV2JZqY7T5znxT40xCaRjShMwOT
GIBx1oxEz4vgkcyzUD6zTUZULzY5+EJ5mKz2Iisgj5Q2Ie6xm0RY3zN9U8IKqfMvZciMW5wB6fGu
A+F+56/Dx9fB5uT/uP6Mm1YUKoqvuR5yRsLq6wbcVgPqjsAz8trCpuwI7wZ1JRG5qGOyh+OFF+XV
4h9CRsZqxlDh5J6PWRr6AelW+RvktymF+z24NHUo57s0XDyg08OyMPokTieG3tTC1duNUq9hqEa0
6bMlY51/qj4Qw0iWtQ8ANmg72aeDBvR+juj52/9ISyx5PPUqx3HP+1R+rSGjhJA3OHfF2iJFgRQb
T59SFm1SlYjw0HfGAs4irFVVfOcA50JnPm2MlVKaMo/UPXoWT+nTRMW9ND8YbHUW5YZ+SrFaguAV
xT7A3jdakPd4qX369adcfFtG4vu3PlZzxhFsZElh03e4fXsD4aFeHX7BE02fJ8hfHw6jvupUpI/8
oxloplPgimQTMq7aYw9xqF901A8QqbXNinBJ4I+oj7eljxVnnOlnPDSlA2HVZeLCh510RrPCzrxT
aF3puruTieaS/1DYmMy3DGmm08SX3EFZDYPyXcjhZQbkzLoCRyVyNhbvW1M8sHEj5xqQiS0HSn1M
DD5Pwl+CFbLgA6ybghnJd3fPkoP+CSSqvtE+WOgUeCqx7rUPPnFhcL1PUYLF91SGAhjrJF8AsYcL
9V2x0vFhHUfstAVjdBru4qJ+P/h31xhZb4y2Saan8bWKuSMysO/2XZQe/NcMrlz5As5DJIun8GDZ
80rpTbi+XJ9/LzzWgoyEuUqyvtI9JIspCV/Q3m2aYAsxihJ5Xb5RcPnoUzt3+ud1RnL1l2O71AhP
nyiihNVcrkU6N8oLScfRuxOGx8P5dadRuxKwqe+8CY6Y9HGDHpOiq3niXZOudrqAHQ52LLPss0Q5
E1pFGAJF/MGJBQfiUb5sx5CIE6zRg+hjCkAoeKPLMJFHPowWLhNw76JFBZfqSdeEVg1BlSafkYcl
WNorSBUPhN23E5lkd+aAI8zh0S9iOe04LMlWGhq3onnpW8MUdDAPgYX07zCZvIvv7LHMn6PuupQP
GKS56M1zkSu1ub4yG37S9gy8CqiWcHViyyTg2BJ9J8Pus7MUBZXnoe66VnzarUY86yjEJ0781ZGG
8kpwyQjoXR73tTw2B1RTzWx1Eefvzl3l6JsHl6QUS/Cx/Pnj856HLJq3I0PT1/u5ZacLeyxZgTl8
DD0mXyhizbIt3V4cBj50FiorWQpYlj1rVg7h618gejNGhH9TsJClaS//ExqCO6Weq82xqdKQcRc3
YV+cc1MbmA+7I3e9zAJSEfI3WVEp1hKYvBvSEBwm7cRfyx96guGAEcANwRUY/gS2OcfL9r1ctFhC
J07hSOHda+6Xhhgg1f55JIbqOAf3r2ahTMYJNcWk6FtRLc08Irrs1xiOQgYjayAYcxAur6m7v8lS
U/5eEOspHcx86qTDzi/yAj2qssBAYU6i6cBPmR8BLo6x0aEm6fZcuaVZTY3kEFaoavgQxbXcrnGW
VRyDyJq6xCyN6NaBBqWX+RNPmKhHTyEULTiH10JUBA+i8mw+yxQ/blIsoOFR1v0oeb1zFmCb4+K2
gP5B8Y91kXbGYqzlP7Ehy8td8VuADUnwmTdRmpeNaCVO6uk1a3sXuNnw8X2wZsolvLtqfN+QUVJf
dmCRODEWLGbzc2WTaEFLUHyr1RAnS5yNBarUyGm0r8hfAP+c+uj13WUbypJJf/ZFRgTbwddajjCx
wDfL0KaPZJD7wH3LIlvyA53zvKmRY+nrze2+dlKWJc9SzhjbDElkF9X0kHkxbceSYaKwxYWQKntQ
ro7clWWmUi4VdjFd+5vykOtJvtkBDu2iD9+4e6V9dkqRNoWpFP9ZQw3IzBESpInPrCjHXWnKCylc
r0BG4Uc7FMBqJQxFpdwtCLvjb/duxuCYwyJwHAXVZet3FF6CxxYCcGbbG5aEimoFbJyU2ULmMCHB
qrWZUmih+Okrsgf7bIrWWqgX2scSmcwd0AV1n0xfqV6/yWE6oOEd0HqbOpRY18q4ITTE35lWOt2E
FKtVk/DGMoBWXQltenMfoJ0M/cX5rMASCAIg5L3qLLEVQUKm4HdjC4Wygma7gbZeWBzK9ZpV3Tl1
xwzd/Vp064QNAKgyfBTl4SmfqIE2pxzO8q9ZVfh649Z2d2W7cVu6ghZzgw5urFjP70t05bGgMVHs
+yRiXUgx9fEsTypX6wK0oXZRCzoAG1wQTOswF98Bmh/yrnc0Sc05WBk+/39yNsNExLw3Miij3ldP
RaT3TJb4g53P1O/Z3QzQTfVIgbe3circggZlDZap4Vk4U8ADBlCWcH5Sda5gGaVvm6hXtye45vLZ
ouXXxZ+/vgUjwXg1d1NW6JsqKl2+sKxTSkeFcvY0JGqubAMCFpaLCHxbpAiw1oybh1g14QneX3Uu
cd5mQJr+rSaso+sqDAvV+a9DKsWvZ1vxqzyXdeTD1PYP9G5iPqAkTuTnb2PpoFz4+o8aSdu3ZMF/
+clZ+9Xm5b6PdXZCa9x1eTvCNLIv/apO4E9/3rAsboa/oD5Oz8wkVjKZ3tsMy28gLp9q3dciKg5B
U7t3qS6EjyUYGM+N+2QKaXeD6nbDIymu2pL6jduxNQTdoXI6YtKMGQ39zUeerwKUb5yR80eTNCkG
/YTKJ0XaGgFPFSq2ey6lKk1SgRs4LDlHs/IzO/SpDh2rk6RQIZ1XJ91V6/wDYiHfC0eevXKviDES
4XnYdxpQKdFxIfgO8tLdVna5Y1f2yz80zxXzxgQytTlfx5O/DaFk9+vV+cOMIAjuIz/ZI2QoaWiz
u71YuHAsGbHC7xp0DBnw+BM7u6yUJPYYvm2VvCmsmhkzQxdnk//A4HLGYbn5yURY0qmybv/4rT/z
K7NHCVtFZ+IlznoI6O9XuQ5mapKD1PWE1S7JJNfzVYeYkX2mz0yqiPaDYpzWwFlq3iMd1/IgyKm7
sv170WCfljJQKXUmJAhy1fX/kb6lN4P4Zu602eUaX6kO8IgPICE9IEOeSJCLbI7AUfp5QO5TbZ7j
+ED7P+z+g+vXy0KeklAe2q2L9ue3BKYRyTnCzqcExlcMUMreO56N2cPuAaHgN2bj+qvtAlIRlSXG
fip1tnU5CCXZWp54pbsLU1PDhBk+CXmM9jsEtnMKK8CnvL148Q0K+WoGREh4ArcGqpGhRN8jiLcC
ZiRZHe4J9zxKnUG48sPHEuE4AEODARb8wxatmWVDKlX6X/bW1UMskqcuuyevy7gpY9F6uNQ2qIEZ
lnvP0duQplHNJe53j6VfIvPL956bw5AZRIVI+xBdEjaMA00FWKizrQJ3kM2li1OJHMJkTzkjjuQT
Yl++fm3s87ucL0vUQZ+Rsc3KmKqFwA9R/MgrqsssDOB3Pk+yM6BJygEwBVYyCn5nYrwp77Wh/OA8
DHorhddBPaVqINV4raIXfXC78UgPMZHsUOuE7/9m2VH64X2wyd2zl0LxL9fmpC0YfzlCJBrU2OJM
c9tVjGu4UIAwq2EviE+uVMSIFzit8CJVkeOMdHQQkC3cT/LN1XROjiDmXdRmwxvETz+EecFnTNQV
8UWNB44XkP7NFv+CUoTcrNRHtDt7B8iQfE7OyB5Xgclmhw0iB5TSSW1gJNd8ipIkwehessTDRGDs
m4Y7wJK4sCw+fmMxXpmsZF+km5z1i+gf0ko+n6M81Kt+wxRb4DrxjpzLh4O6PsPXztJfcFtWvugz
vY9kl3XExKoKWYRsZAYMqaDxRbz34lWMFwVy4CkEjX3Te9r1qgxg8UhtpW1zdmwe3n0alOSiIF7S
ciPoZo+4EbJLsfCHKa4GMxtVCP/LKBtQ561godFFN1hzFqm7aADs4MPOU1TNImZ1jVxCiaD0/7ag
xuksCjTnFu2EF2d9xz/U2CwgS0BdDKyyWJt0Xi8xTj4hU8LprE2VlQ/fh3n9E1ivDq+9c1JiHtW0
11wkpaZQqYBgIu/ALuNDUtvGiBM0ncOljsENK02kIY/sEaK6HvsDA1gCKvcRclT9OPYXMT5z8PPp
2QzWeZIIXz8yxR0QjsIEKYQRAe+pnGCmofxyKkvvwGJJExK1FtHtnTDMXkAiLTkVdrYrDMOY+g/j
Idb/MS9W9QHI9CC8RuADrBui13MqGe8Q1BoJrOKDUgGPqZnCz5RLWR87uPDyeA/pQz3UH/8KHDxh
7t5tDgbTCwmOV+nl8nlra4TcUu80PSTspVOvV2EWNKI4TfSeKCZyLyDHFvTteaFoz/OeIc/ffs1l
HmayvRoGN5iAz6GiVx0zGZolerog5mwQ2ukGjOloHeiMYnJ36uova3ncVc+BHb9Dm7AEmrZYY0Gz
1dv6gdufD53wFid3aiQ8hK3Xya/xrc0cviGJToSNs1Pt/mterWfbWDdocyTXmxI5rVX1g3/4kOVm
QULU/6/Yov5xykb4UFfX2NVnNvQ2g/7r+3gy8QsR5OzzS4TinI6r2z7umBx4dAxs6y7yAqXCGl6y
6bMjG+tw3ZJjyT3jaZs5RzhWcp/k1UJvnbN1TMuUcSujVCl50Qlt9WTMDVL1yhuaW/NIp/4c1rLd
5ANut3XmcKMmq5x0MJM1E+5ql1p3tN3d4oVnRRfyzw9JvqH+KR36Y+otmLzkxNEFKgtg51jaoUWj
ArzkXr+HSgs585Ejv1ZNDcIKwD8CcHFtfRMTPET3zvnteIHUJVpPTgXsLhmwnMivVPMs8aVGDT4t
Z9OsQQoa3bI37aBqn1J72Nta0dBUQgIWhGCfofogekjD97kYbFzqQ/WXloVtLt3Q2T5VFio3xkzy
/3QQ9MRUqbjuLKV/Zz/PbM/phhFnhPpzD2rQfHkYv420QXH02b4QfrWi2TMX1MNTGbiLIR+hsMFz
cdiZ5ZodLnoMqsKNSZ9tHdvBv1uAYlmStSTUXOr5ZGqlvomu7dSnK3RcVOIMJcQJYDDpDnbd5gOU
m5J9BzzrL2QGrIEGa2akMbHxCPB1BPei+LA2Kz53s79XYITyohFuJRDhPmT7imh6iFq5pCeY1vuu
hqzzhLZl7iPNLU/L1fF05AdPpQIiX9z3ID6ZPJEc3IKZbV7z81Wxs/ReA62L1k7VoVU+qtnPGpFG
26l3SU3xcrsbaW9wTk1bjwhxv2hX0ff8J6ahWy3CzrR/BMGjdP+jXKA8Uo0xceJVMkUbkvU/CEPs
wtWYGGsGHyqQ7h1qg3OC+ElZmkKYY6mPgJPR+uf3qxLmQMkt8ZcJtSXZMcb+LSROIHtiTEWqzk5G
qmSCUWLC/INUYVN+b+R1SXoMV/I5Sf+mVKs8hwJ9xt0+rnqsWNZ9cfUWkouaSjRw19ZkJjmY+twg
TrjjFASTdzwJ5F/82ttTzeqUa0qb39y9KtNKgkunrLIPoKt7aM2IBfBF5GRnilCQlcpw6Sh+hTfj
vxC8sbmPYvP13AzoeyCcfyQV4JqVKljDosPcdNfipLacxtipfQKm4zLa7OwzMk8ijbmJRl/TI8bc
mn8s2X0O2LmcAeBvgerNNc5E8pnwnPU/nLRWwg8rr7z4GF6ZeFTxfncbvbT+am3g26ewRuFMNSyh
vJmJriR9Ml4iUE7RAXyamo7MazMN8Sm3ySHSm8xV+W4mkKck430Cg9rdRz8Jt0kSLS4PjK1b7nJC
gl6S7wqm9TYjYZv6aJyk94hljiyaFf9J2gZR6QkK1krUH7s+0BWEKyUczHv2zaLjX6/wD2rru/aw
C6oqX+hJhs5yQgw85wiCO9nYPdbgPVNCClmK5Cg+wHTNMmUWMdk38daA+8hRkfvgdST4kapM7i0j
nPk3PWU24mO5/LElF1GPgDqW0hnd6qvbCzRUjg/74CwPtb8sjscErsB3WFnSEfw0xqu+UVgvqagf
ZUjVrG7iC0iYTvGfsHOBmiSTLe+F1x82PO/0zw75Z07xWZIYSLS/HFfwqSt+BKLubulXfLcxR2Ib
oF+d4WMu6c//bhgK12VeM+K5fPVFZo66I7Obrh7ctxv1Au5r7arUCL5elb5Cgrv6sCbOgYd/K2Tz
kaWLG8BXLjgB4QokqLCU3mPbUr3YOVW9X7Jk1qTNk7ORtv7AlOBSNDAuPf0vLREZJF1He30Ty1Om
9hLlAocBwUDxqfECdtUqEP9dwuHiIoyiK+jRMdnE/1rrDZOJFnAfk3HlUSBJn9al3xqOAOpZPA1D
0VhzcUSOx0scYz/gtZEOk3Ka6PPYsp7soHLDREWl9plILVodf9qy1X8zAZ6bdEwOt+08HpqzMWt2
bf2eEWY7LkfNSTmoUaNJuEFHxRRVk96xm+u8qrcAaztwOEldp6mh3leImfWmrxqF37sf3rI+S1rr
Ba09LzxgD1QQmI1fQ9FCgyBAHE+taG8j29SwfdWeAZmdP/CJclnxzP0B/PWnfBcF4dFr1AL2awEL
tNY+fcLVoqTTKVLjUfLwFNgi4QFFIDFYtpGd6Y0/4SVTDivQ1xPhiX3fHeVyAT2LRzo9gzEHuu5f
urdMpTOQyKR3EOPgGJUqdjmBZ5H3vNoPXh1T8cBR2xnodSjkASePLEjJQcFl1Jl6g1kLJvxj5RoW
NlhxNSaGPjJdQ8qLGKUcLvJMZgzxv3er4M/bEyh8eL/XRzLhMlTkQUmtIw5UVEc36uutEfrzu1v+
D9ZL2nFc65dF1qnAI6dvQbU9sS5PMFWogVvZ4h5ROHOqqSpIoNf9rT6TdRBrpmKOjQ0mAFsTssDc
Gm7IesSiqhYqjf0zouH4jt569KyAxyvlCBWTMYNQbukkG/+KCzxqZmqEu5T13m/sHZdV4mv/mxU6
eR/hk3udXzYrc2sNZoG8P/LP0+DCZpZiQNVCgPXZ2BQ3DBTwSFehoiad732Q63A+21cC/hZVrwf0
bjSPbeacLy/oq8ipRso0v3vlos3dWeFjS+ELoU1KpO3btZKYHMur+osn5P2IawIb9wYEcHPP128H
4rs+UV3aCQxYeOqhe/vyd7Pwy71CAtlKzwGwdlOlDjNz6dBxNj8y/Bofb14aWpq9GTWXkKrvdYsP
eRsnVs++kQI4+MqpnHR0VHpJtKB0051jn5cox4xkC8elDmNtypeuIYvGG56BfTcl3rAVZLxuUAA7
fk0b/WxwBIgYo544HI/qF7LR0nYbrqQ2JG7+SqEHXgbDKtul40VGvCA6VKHhHIe1IAzQE5GsgMcr
qz5e/FbEhfrJP4bnLVZfy1okQJYNk+V+tXLoBoTdMgFvTG2/MbztPfAp4go3RssDm+TQe38yQaKn
4IDbgJYuo40FcAw9DTCBvm8lfU9XN1rFzN5vLrTyrPaA/ttfuSHaGuipn5JCX8wfNTQ8C5nPo+ZS
JIUMyGtBrVIt0PpUSvu93b4LBUO9aCHQsTB4f7/PMtvb25H4yKxI+eoA+GWoDD41f5Ly5uSXo0jX
KnqBVUtG1uavTEHpfQGAjqoAUqdYtyJofb43PMsD9NIaWSrRNLV3s0q/NQL5/FAcXfQ+GQFRq7jG
TiAQB3tujHekyFwAKNHP5AoWx/FiHnsblftL9/taucIUcVGRZJOfkxce8BlTgHuZl6D/meo5g7k6
ZIiE93xWsNzc056Y3y7gWliCa/t2oioA/IMUuv+IXWNVzpWK9e3oFCgBBGAiozz0UeF0tyjnJw4v
nlDi7uDDFrw32/FR+LUP/EIBfC9SdzFZPh1TM+mUHkvUC5kXsbAONnDvpcMOCNle0iDx4gfq3OHP
MWEVLsvdu9ycOtuXkc4C7NxYjhFw/to8Ly8ryhqp20et5eVMP9lIoBKlE9bik2UPDHmpqxEFdJFt
egnAjn6i/UtIN7v+t6t/FDeroseLTUxGbr1p4DNyt71x4q0MxHrIP1GiSS4GcnlwA2K+uGaQ+uEc
24l7QGxsmmmz59DzINIO36uH1M0ag+VFmPlKI1RIMmWTeJcyKlt1nTvYgJmB6AcrEZcV8UFti/ka
l4OhrqFmhDHSn4jyg77xF4Y+E5XGE0S1xRCs9F9136w6fyaCJ129hU3Z8Lk/JKCOKgY96u7YPvR1
5kjduZI1K0tn38MgYBdhmWpHY/aXxzT7QLN6rrTs3Iecck4J4OJtm8i8kAhtcefHlEdLcmrIWUP1
j4XPMKEqw4lu1Hhq9Kn79ij2YirT9mG+K5md3ehR1Uqk6U+oUXiPvCTqT4yGaMarKapjPAb0Swqs
uHLN0XWcLu+wddC0Hr/G6l6SYiOov9i/rSya/IIEBnfZbML7VJIz9on0U3nZNrf6CMkhe2jShGUs
Z1CeMj+6pcca+aiNyxynQYoIvA0LeLAMWmP4Zme8V4eR9NMj1YqlZb41uO5JTOgBT5V+nl/zVblv
CXsiCeuhMJiR0U9f4zKb+yvVm7sQlNjLooMVKGe/q+Vekndgc4ww3SvSHXsJpbUQZzOQuqNR3VYR
YEqpzFQpVJkYE9gPLCKIJhugOKivwvxr1Ljr83iM3SHm7/kXHXmVKRSGRjVjDfI5RYkbR3RwTPUy
GFMvzIPu29Tz6t/liphI1FRtsZhYYVj4z1ao3cp5SqnaUzXR/ASWqswIFmQ4SQu82ce53GpkFv4H
ERZsCb8Z3+cmj1gGP+hZ7BHCrDEsiZ+kLR2Ga73yUm8Jm5msn8eKqJ7sS6Ts6AvuABwqjiHiU5vY
4YScLGgMeVQQ8YX+7THFGXd0SVC1j+YxEgQcM+Wb8i2OSTmRj6VTYH4oWnfeUiShc8uv/q8/FgT/
q+IdmKjylrO4wgVfvYjdyZM9NAPFVTOJQAqYlQQf6sGJ7iwB1ih25ZzzwuwTLEgEHG0mj7nZqyEk
ldgroJa5ajfr+dnIlplo5iOm53iHQQRYfilqswdPjJW1EU2+qkLAb6dgqtZap8dLfeNcUcpZDUuU
pCMlOOCmzBY8pi6gv3sGeGOi4ZgPQupSKtb7bQjdLeKfgJ9W/DiXc0QNQMpabDMbJQfHMS/bpoav
KaqAnPCGJKsas1Zo/hBGYcJUWCCpALe43UBeFr1D5D4Sgsd/ezn37UcA+32xPMk0rfGcE4yz/Q5e
8aoaqpfF9wh8eLbT05dSs1yVa+midyaqLIwYyUUlosBB8HFzr8bqfQUe4Lz5J3w/hWxd1Ybghnop
Gh7JMFq2FzOSgTTCXvh8duYOPJQs3NoX9uqbVBycyFNQye4MSn3zCe6XyJmhG988uspS8ubiGCQ5
kXOPeQ7DTw/IaAR0cYCL7+vFKYoG4M80QzzYocWxiSTvWzo2vOpxr9Gc5t080cDtYy2f41IrPXrA
Cb1xFpDa4moSWGu9usVJEr27ahm7uEGnykCL5X7JJ9WnL4JkEaGw3wHdTnUYCpsTS6jaeWHK0/Y2
WaIvUySDZgoHillv35GodIphurod4YKlOdDhszChevtLqyH7yq3F8yy7z+FCdNbAiU63VkNYsFl1
EWbYS4SkwVci3XlUInuUm6Q2dajPkGZTDL14ylH2Rgf+rmo3ZhJaqArB3l8U1Lmsu5KGHv2Lo6dd
XfEiPnFCrp0X0oxuPY07P/mDFqSqKvJxARtS88uVmemwvib+ZQRWvrDLDHbq4hUztH2bHj4b6BKf
Hb++P5Ei/3lfp1nPRZWMant/pddYUuQHUE616xHKxTOhc5WW6s0qpanNtaphtVjuDk1VCKI43g5r
GO4E7eOIFAPaQWlB34zq2bnreMZfjVp+YoRXzicuNI94Iw8kSD3QFQjHUEQj66Lwvc/XccJcjuai
vvspPbhaB9j9NEslOimO7Q4b9klD7H9jaGRjTY/QBfZrGupVsKSbzMpbBlqMCoZ0n622u10DU5zg
aIsoK5WrjtfwOaqwCD2A45gQBJCJjCtYOe+fRp/+CHx3+F5uyliubuXTtfc3G4Ct9Kz24sQ7HRQG
Gpr8MXLFzzCFN/35sjH6Kem7952D7bw8Pjv4RrnRrZ64pjzqAu7BWes+s28I+76ClrE5htrtWwpN
onN8J5dsz6drwjVjx1tGgbhAi7Nkg143bSZE05HdBV4L5gIRKQErcr6ve0d8lMqqUBKoADmU9H14
7bwdj0BUZ6Oh3reOYf/YlW9iTr+2SdHpkGO51btOkWodY8VDYokDsz13jS30TZz+v+X1NB/Bxl9v
S5FxodarDZYT0REZTt2aE4KMxc8iUiApspft4BjSSMh1kavaG4E9X/h7n+NO+5pVnUvFerI4Xtk6
zepJfL4gVBSTsDEJ/I3zeT6S+k7UgNcQsbVmsSGtepP+nElNSq8iyLQF1Kz8jSJtapQUIJ+v1wf9
++RNYDYXAJ6DtNIMOpneqgXPC40MRuZjOUKHpuALMc49dh8DHl23LpQIXma27BEpB097996PUTP/
Izr53JW8v3As/6dr5YpdPUzySbaTNaOFVG8CEwCZa04VqkjPQxjP7HQrNCiT90O0aWtCVphj6p9t
EFGutNMXLUmT3xS8+NYFO0FbwEelpWSTZGt/pzH0BEPyIzkG1tFX997jgzm1eWgujZ0OyCIVvXAQ
JwfAKPv6Yz0nvxpKbuqQvooMS/oMaDtPODkofZdSbEFy6w8LZmLc0/dtmWje18s4HaC+TWwPoBAo
BQq9+IjTjrB5T6ZTpkOk0n14j+saevkjeifyT04nDV0zzBryrtc1S7EuOHdGwGlTWjq7o2ADMq6/
nbZPW35G0X6HJHzm3WB1j4fUhvTxUHBvATop+jc2lXFmCMagy9FvJyPApE/2+Dqg2xsSTot6go24
y2PPn5YQh88WraueVQ8yGSzbBoc7QRJPX0k44m9G0qlfs9B1FcMkhKM/nLK90DlbiYCUFcLOxunT
r+g8cipwC/29fx+J8wnZBm78AtZqJmWMXiHlygE640zKeGvY/sCq5GRYI0MTUyekw2//7INl6Nbg
MJAoFXx4W3F24RL3B2I/mQkxGV/CdS5GeHOQ+jGQuLgts4lYAsXts47PWDwhNiP3qlDZV5vrecYv
0creM4p0buVXi+8iyT86KUPFtMWaa6XZI33oWO5tZBOnEcxGjFhHCkFDf3BtZEElvYFPTB4kpzSi
NhM93u/MxVudKN9n5Zb9dHtAvFnTEW0ZWp6dL2dAKkb5fca65uuAURtR1BLBgXpcvJmK/8SpHa62
gS0zUxp8ztpbu6QiSdpWgay4RO2XxsyeWOJwDOGh5HypfdOOZ7+vLnNXdwiFeE+ArK5TnOAStiEw
EktzY7v6kJOm0AI279lmVXOej1t2R1U9iBxB29dyVwtdSiRB3lG+FCf6vLTD20vMAEkaVRWy0Ebs
1JDlzyDZ76AjErNf4X6fYQm2klYe3UOKwyfpsxUHOfVlu2FsidxaZos8OEHDdfzPqtJsJ1vwZX1b
iP6BPeUKb/waL2ojPcZdwBRWUHJ66zbf8PtoioaQJ3ZD9tNveYbvVtF4Tc3qm6HGnUD6d6hMCtOa
GOJb/vPPUj5fOgaJ4u97bh8JcUXoIWuM13Yw4hFSI3XZxSCr+fXapL7mWQijC7Fw7PSkJCXh9z7D
UXf4iS4eYqEt7QsmeiuPXx8VrH/eq6Bcdz0RjfAldT6XdYOaT0M+znGYK5ySivByCKsquKAkGMgP
SX/JPWTzknapLRyvf0QoFinYc+rq08P2StcuIk5H3Yym4LGZ3yQL+NWzKsKb/DlPrQzGPFm42m/7
H281R+pPu25dRte8evizjX0taBfE8xwASIUPAqRwt5x6XG1tb0Q9/dOCrS40Q2IJI+mnBzDy3Q5M
4DlgJGjN7iqfFEc3vxaLHz5fF9EggAQY6U/VOltyiW1TM3yZ0cwbzFkaLvFgyyGYPm/zA+Tb9mbO
qe0sl3KpXy70Lg2f4xxxTXvkx6nVSIjhaFtUDF+NYoznkWOsu4asxByax7aNcJqUz/XxCQzzoGNn
8XKzEGS9B4y8a70aPGg8hqI6FKBsO9pwUGgvSnvziwTMRs+C5JXr0+h/BP8Flk3dTo8WOSekF0RJ
jVKs9dJow9FA+nNLNY5BHcNbevNPa8awt53FQN7fFoLQADxz8loaePZhT1yUZh7TizvdiR+sfNc6
/b9IUVFYisBRzBe8e5rAnsSfmHJfk8ZOEznnweowS5ojPlNGis2Kjfk8Eu+ilmfwDnYAeUk2JIgh
2fsuoNQdbgLeZOdv7ShADeVQtqQw9fnOwYW1vqwrInWQwX7lBsPyIUOdMyCO/ChtqxlRETo3IH5/
SCJq/OfG0GjP4o56HTnNkG6jn73Q03KPhXUgI0EsxuzBqDUd1Jntgwikj6z4urJx0GjEIx91iRex
HjICdsVcvfEGJe/4WiewJ4krvAgw8GLn/N756+o3uoFo2uQ0u22+HkUURJaAv0sOw+Y8zNwtEdHu
26/PlN5yusUfQxSBI6nOg53fT+vKpjZedAqrEgNtDdLZp45K0qUx5L8fsi0HZYYhYQYx9C2pGf9t
zqSjUo+THxFT9J3AXTw70EU1YNEvmlO8H2dhQFq9Nc5zlQW2YdnicFD0K4jX1CE+DRWDxnRdvaQ2
UhyzV8BCfsf0tV/LMdRtavNmK/Q96ytqMUsfZ3IRnAiN3u+4W6iiw7CXmPFLJ0LRAIIgOkpjVVOL
cKd6ankxcmfq3XBD1J/eATdbvHSdAwv2RshPWoEVIInuUmrgJUy4o4sO3rGDWRzhKtaryzHnycXF
jgy5Oi5HLCV1bupoEJ9ffrGdf8L0MiaDtrgXTIiVkI0zUG7bGhgAMi/6BsWAUt9MD5dpQxOhwZkx
uTfbC34+gI/XBdMEQFyaKbmeKIa8pf9kKHU40m7P3q5r3y9MepZjA9PmBjCjpwVevHzmq/IQ7Hb0
tMdyvZJcz8VwOdC1YNQriha2koBkAQ73vWjgKWLlmXG2MP6bjFwHbVNaxvQrb2mgsL9fxFI8U5TT
Xv4u8XBxgI4BiQtfxdk1SYH28lrVaZkDMexvHzPm4/bGXhPrimYg8H26QC2izS+ufwWArdp+HRyI
+ZtpXyCs85nP5XYy+v5Vua43oF82eGKGShpOR9FsQWTExuCj1VmZVlnH1jQdX4yVop1gTNVrk1mG
OhsN+WHeWrWvfr0/tqan8PjnHo/CIZSDsaCZz39mW2Bz8IsKORnj27y+TVEXC4WDzLwkip1aYz7f
d1wnsrVJ/f4ACpEvGEcja0dRser0VEXgu1cDY5LAq++mp9mg5bkaNfn5iOsfAOiRFk3ubc8kD7qX
7zdzuPxTCyk33+0jxL1wR60KrhKs5jXLRqdcubyJG6P8XtRGgFa8nbIhF4fN64R0LmfxaieX/YkJ
bjz5WPokOVOWUPEf1anGJOn9QEP+i79twBE6pKiFjLMCdO1tVvGj3BqcGaAl1419diPGYu/LYzC3
p4HFMRcfLdkT/1Wbwa/pHUqcJsQCz1UcJMF4tIQitqrU3zTq//v3GPTlIBK9lruHDsVP4IkE5dob
O2YrvIbF0Qz8Lzh1+UxibPMrY8e4aHlpSY5r7AI/mLxtkiZLvMr4KAx5zO3H/rDs2Abo14rk1+6c
rWjuGO5sblCtyHGfZQQzC6x35vLuwu1X+aIjzyAgVC0DS2bdNDOcS8P0DIIGa+qwiwBVKjyK/0Pi
vehUcQrw6gThsyDPPgiQl5sJ9Ief4VR26jHGfhBU/ECDUPEMER0fuGbK7mhoKqa3YEmhfbpyGUe9
wI/T2dBCEKi8GhtI6Pd12XeAV7WtQtIQ3/vaFRKpCPnDOnfGe1bTZiHuY9WUWvm+qn0d0Eu9hh/f
uH2S16MFcOKc3tm7PSOXVyNSsKAW3cGF5+aVjbKH7FLo8lnTkzVBFEQCNfdZ18FqoL65lDS5ittB
UMKJlCsEouVaG2opGXttu0kvJ9OSz9nxc3UkePyqiOwMPIr4tZRVh014CeN72uCs6gBdp7Yx+iuq
XX3ec857r5n3puPf3P5/j0z4loByut7pytg7Cd7ONL/ZhKrul7+ktFj1v0bkAHqHvI4E2ZNrpJpa
ro6HX5AK+bJm1gHvYRJFLCti6oYcjkKUPEvITWtoNOHL+gpy1bzGApw0IQMQiunzy6EPb9XvMru+
pLVpT2SRaKtpePASfitTeY3ieiSZNzH+vU7xJCBZNmedUXtrp7crdW/qBsq9QenlDo6NiU7TrGpA
65qxWfcFw0xpnCnsGExgHwpaJuE3fgzspgMOgOeojRvlHMCPlS7BA5/pXr7LYAmVlYXF30I5BsuL
zv0PiqYvkXbEvUfD6E9HyVr98yLRaXoWy1l3OOw9ictXVxNAHQY8PqwGYT8WEQqcT5n01UYAVSQ0
zRdeswWIFRwp8po5sjxMbBc5fTvT4svrmYaY+y3FmK8scpgR27nMKzqGQ+D0zGrf4L72WCNqRIg6
SFnWkiBF3nobrjVUM1jUIZOloOsr0mtvCtpn00iph3uCs+ad5V8lAhz3RSeBzShOLfnv6Toyw0p9
x2jy93ANAJzbphAR4FXsEgrwPgPilwMuR80A7UjuqRgC2Us4+cVO/jkyksuwiHnjfgegMXwk11DD
GE5oteqlwkiQLMSbVb3WjFOtw7hGesjoNYGMSqwlnbbzvfhcdJfdRkNcLxHj1mTbp1h0zk3Ml6jV
IS3iHjzoQM9gA9zQGiz7AYtOsigaYwzXCslAQ3/K8mr4nBI+h7nWGfenCqu0O/+p+wNfs4OMaEgp
p/gjqoxjDQHWAdMDKL/gEyIcYWXtMPYAIvydwtYMUdCszdOKdKx5b1czcPS80ooJzskPECGwiAJW
xS7lUWIScbpGENFYNXtgWjmWZvsi70TMsn1yJVZXIxYJi0Wmnt7LCc3vTwQ5N7FOZoQGLp+BvVhc
pHLhAYFNlzrFhl6lDRaqwpOj/dRyu+VhDyrBQ7T2dscLXFQsAg4GM1qlnGrb9mVpLGibqJobE1t3
DCVqUBcnOU2WSeK13HqyUJGmGQs9/JDoozB6yUFjUbHqbkKM3zf4HhSBxVMQY2BixVdjGPuWcrUz
am5Nfi8tvFEuMBOQDnb1wqUli7Wxn4xtcLDByXoou0PxpK1+fhMvsQXWSc+ue9ZcSaeeS5KCho9G
ARZOrxNiUawdA/fwLPGFcMLVx8LnYMchmjQV8UX5RWF7P/CziArwzPYwGgI3zq/QNvNGS/JA6NbZ
JQZfc0eKuT29YTCHpTM3nLxcCBynEgJIEDWjTzeCWPfI0HJfBee+dTyiKHaBTPxQPMVpNRAzCJ3K
NM3d26ghlTV7NGTXhdVFt7JUVX3BSAt3bG1kr7GrZW/+9kWapS4+h/GCdyrJooqVr2chSpOBQ0Fg
bZDz/mgyixoVySXLKUH8pjxIagZBPhu9mu1I6z23BYxYHaVfVAABteIZT9+aSlPiFbiUSxtEH1Xm
UczD94SfjAdH2jR4bVcEqSblf0VVafkksvhjBdKFQsvUxMsfMAvVMEWSjMUYxf5Acjn40jtn5w6K
yxPUhQLmz3LzXqfTaw3XYuyoYze43TNqy0ODq31thZqe4lRY0z7f6R6uqs01wTJ/zSQZcMTHrDZ5
HtFgjLVpOrmafj32OOmNY+/7D4UWjdVcki1yQ8sKoVqe7YA33HKMzdHpGYdsj761s+ayn5889s0Q
SCnxY/h216jt8xu8nDb3hsVfKw04t4lg5MEJGUkxBcMctr6dMaPhZZGuA11ELNcg57jZpNlpRpf2
wpS9g6pFU63Yz0f6QxjqWJF3kDIXx9t+MVL8beUeBc/jNQqbSmkMahDjNyN6NRQWDQ7lXapB9kzl
fwbk3bYNqIJuhf3teTKpnueYJj7z2Pn7iToDYM0LNwqnBfX/CtqWVaH7s+P7SQHGZg8kbDo14TiP
kajJuOrNs8BpaLQNafPv8jtDBilQeYRUlaHJsWS/f0UC1OyZQrqGle3c94cxFHzPXyT2GnOX4U9L
1iPC+H/fIs+z8dm5V+nvHzXIV/pKKhi2usK1HUu92Tb36RNaYzlGXrS4XGEGMbFOVZ6KJaTjSoxz
ZfvIcuhjvG6sku5ccm67FEDU/4ug0+MoOuGi0PfTDjOHIqEERqPBzDmOCW7pPKTWur/tZ9TyYODZ
ZYNUKTkO/q+NGTHTur+JFxXFPNUj/RpRvWYYNhJyoe4SpgcCDKCnesawNH5W0o3Xy81Ed8OcIiv0
5IA/xJ/jEBhsErgrnmSlSPbvjsTSarQozgYOOjWWExV+XcY3hdeJHdaug2zdtWecsCVyDRmTR0HD
iw4MSFFBVcbEBVKKXLegiigNTr4T5I99X7oPvRM6BEpIQhIc794oA4GvEf4+hlcImR/QHfHTzOeV
/Gy59ZIBKIpmg3MZTMKsfPiMe3HQ8uSxU4J03wub+mv9kuvxqFcZmF3pTQ19569lX9VfnVpUYGsQ
GXAMEQjttx6/3HXY0gu1W55dANytina6kRfxcVhOA+EfsgCx0/77YjWEsiSn6QPULdTBY3dKuQfm
LP0Jo3hSomOnxUK5ejIMs35WjooprW01tAww/ppPqY+Y8BUrLfq2BlHe1Y+b1lEm4LN7TTNwQQN1
zzvKfOAwpfyHcHlFuUAyp1BZ46hiBdfB0xFdrjg0uxgOI3HNfQ78f/9nl/CN5JiJa5IFP24eKI+X
Zau7H27NaKUVK3gG9tnXUihgb1pDxeFwmovr8YMUQDOD3N74+QIvfBcBUYifPkQ4Jva2ybUZ3tcg
TtCvWfEWmmCE6enR1WnogZOOYCXCWpsOv4q4rG07njtkVlNySAcqM0GnjacRqn6kTqHmZvb/h0yy
v2O4ffkV5puQAyzPiZyfxvlCJmY0sYxFLIjCDWPnbJkdE7gOr4LDp1TyyeA0doBg2aklHpBWPGjZ
2WjX7OmDlh7+qog+oCdog1Jp3rz3kd3fy4MKsIRXJCoBs1cuM2Pb3wEvgujpK4o2cQ2NFpk8MNcX
AfU1DRCLKezzqw6c17apwMV03pFCa04166o5lRsg3egoYs/2kNkBkEynaf8/+cVWmqS4YNtK8r/3
MjCtUwc8ceXBBn27l0tA6YKz34REYFOEYYcd5aiPY9pUmX1rKu8gRsok5GoayvHQKlbhKERKAF1O
JnTn6TiMhufAl/MzcF/NhrtBP1I7v8ciM13K6cyxLelsK3lqVteB5BW0DRyQdcgBwBVdVuOwWzA9
n8jVhb7X3o0dMgd2lfjQlt5Q0I272QIkUZdWIQhOw5sVrBsjWA2mHoRQ0BOWYeMFQnNJC12Yt1mU
oCIZNy1/KTFTUo3sjamWIFH1DItcAMNZCNMVh6vuDBL+CJhxbrXjpwPjiuhrqqAMbkcKFmTqnF80
bzIX5Gm9yiAvxar6Z6iYHWVTTcaSGuHbrVy5i9ogeRDZr+5AC4oagl/IyTIaFs/7FIslYYYAqJOK
BTnzQrKEg0pLtjJR5nRuCR527as8pLqF4tKx7ECbGqO4Datkp4i4uAIQHwRafwJCKXSjbabIiQ4o
C2HcKI8MO2hM+/5pTyFMF8/MK6rn00nzIB73BurQAxrmmkOEvuotWurI4Tj8lQ+pce3I82s9qKl/
FjH9MXNPV83osTIwwVg7RwqZzZHulJpZyMyNjwc2KRyuGlA3STMht4eNeUHy/LbGA1ZhiFLhlC0J
37oOHOpvLXvk1ilvtZakowzH2UrO8whcC4DYlZcB5Mf0I2DIIrE4r/Dvu3mlYjTs/DPJNdfvOxsG
6gwDgBR7krnze2cTVvbLnR3Y8U/jND4l7qLspYKWOrI1wHp1uBoPbkiN5v3at8iQNSld5LuzHST0
aMDXJl7nt0lzQifXbBzxY2mBmS0w+NFRMzVLyodo+34aXULY7/6JX8Eexdm/nCx8cDUsPgwSqkQz
nZgcOOB2NPIosmtrAZPy8e12ZMj+3QhGFBo7XHAHIeF00blY/lXJdF54ezt5tYw3h0tK809my4KI
1Yw+uVmGdzA3PLGhwgiFBSOJNKVeys8wkGo+N0UxXPId2PWyA3/7szLVdiLn3ylf6PDkbKnZ9lbC
MkohNnviD5sQanpqTWfc2NUM8Te5rXvAoGrQhkabnVL02XSUPEmh8HKok9H8pxKv4NwPz53Mmq2A
+SGViReHW+gYwvSLPyNtvumfajMlj/+UAYKI3DWUZAzTHMg0lfw87oqP8mRRKhkGgRA5QnfDU9pu
UjiAlObjh9q+oBbTFAxWBmTo5t9Dq4BS0fiycjIqNp9TMsZr/Xj+gtZygMmtJIzEhy/qtSGNBCFL
+gSkuB+CHsCMfWfqu8BPxHOFClgrh5fGk9jGbx6350RKqkB2cOfiC8rAC6LCofLK1gWWkAM+d6OO
dAvCu0XJoN0j+fFGjE71oY6TjHMNr6Oa0wuTaSZhjORKDHAGDQ+j0HiscaTxLvUqwMXgdXM+f5Oc
SkuaK/JITH+yb8bMwq1Fn2eFqvAoQ+3G1iz0L3KEYIKu6vJhIg5Ldk8OCIWvBojH426FnUY4oUPO
N0T62tLQZlOLn11wWb0FcAMCJiGpUJlca8gfVORhBjDVbz17+2N56c7SVlLdy4AVqCDGvq3OhfYB
aJxTYrrJoObpRx/m6vJeF2Y++TY0VGKSVLgHT4xzlKZMHEXHsZklQyHOeJntJH99DB4ykrOfMURJ
OTd7foW/eLh7ykPu81DvqCZuD+f4bWJ3rWsnaiKTbD8f+eZhi4ZCFXtkYRSO/kt8afWF0syTC03b
ULAG/5+I71Eon9G8KkZILNC88+uRgtDTYw35Twv6VrVjI6j6mZY0gpMy8Pc53TvzB9t/3svEvWkZ
/akzZ/OgLbQtttVzo2YpiWe38fUyS+CH3RLhqlEuEp3zYXYmiMJCauPVgi3HMQY7NbAojpSr7skZ
8ZqupDfwUgArHVJlD7yhNxw4471nuBBCWdeqs1UjhE6ErxRJoXbXKT0KoDKrqQSIsqHaCrIhAurF
h4oSYSwl8CKrOX1BRXd4YZmGAd4jSDhUkj+wm3D9+L/1JUgW5msaZlTtqGxcoL0pkXthLQJBP8aV
gouJv5D9wv9b92GZW5fPVm3VFB1KkAGubZ1gC3kLnxwS9AfIua2S6sxFaCZj6IqpF/PEsgLcgwsj
devZl+CzB1cniQR3lfiZ6e+njUhGM/vZ5wjlslGyfZzUEZltt/kEAZyGQEn2XwBhVKn7gQ97fkMc
BrAonm5F2+beqt6x9I3/KhKztaIoQOZwbCWhC8ev69G7sbyXGmRkHZdgK3HBxgl9e26yf0qCQz2K
AzcizD9HfP1AoOa5cI+6cmRS5L0knLip9+B+BnJ8m1xhdXAMAcLyaeUAKT9KO8dRVAXejG968ko0
qgrY75MFl+u6buu12wVXlbxbY0Q/ocNwC57jyQjYijeTbSOF9h5JsZljf5hJ6jYFej3Pga8uISAN
Y4PjV2d/qSApvl43iwxJVoXlDnRIlQsJwAHH2UhFr7QCgm2Pfoj76VgOjFjt3zaECDD4bApQ2JnR
DXQZythl8WazMeOH/9qYIMzsFfWGzvMk8nESPMuaWnF8G/s54zTibgDns6Nv4HBYWWmjS3TuK0hn
9J1fKKaImtDYTDbtpYQP7ir+EliXvYpcmzM5KFkmt6vwM/V1Bs/g9SJbodN2Nv6obtOHNMGD/zuO
yXLRgGkwCvBpVDEtnHgguL1K/Qswb4si+rnDjkQq14vE7sM8oyziwXodPwss80Mv+tGosFNc/9+J
4+iHFV9fa5XL4VzcwmSXeXquQkw3b0N1WxKxKwsI1FpeIUD32tZfmossLIqkYFyLnZb2jkUMpGmg
jmULMpzzST+Lg3emjE894NKYW9NxKUgKn7we2QkNJW+MzEBGjTqk/WPCXx5sKxf/h0BqXMxXw34g
5VWgRraJ4y0WOt8TnjzdF2+rU37MrS9PoPmAA1Q+QSAFD4MMRWkBMcnOSbVEJPVmqlTqFwgvdn7y
GW3pn7MrPpGNK3cy6HiPOiEVM4WNsExYxgO2ms45meigqvB0pq223yoqtkJroLhyXjImSL8RpsgF
QybXN+UiOcCYDmRMRZaZj9uzLGGFJ1ndJhCqx9woOxivNqFH+LfwV9XY0omrLamltYXRNZnu6Y0F
UsXkYIDQvcACO6LGNWyC7itkA+PnhMs66aDLsCmBXUsYteMDrmpsUtKhi1m+prIHQNbmfemPctdi
YEXMCGmzfyfrnLaBal/b8a2KCAvmxpNm6SsEGW7yC2yb1YJJtri1XSt69wzrD7sSqrbuZ0qafe4j
vKlAgJlrH2QS8FENWoMKcSO1lJFPr1EfesTjYqCCI/NpNjG8KlkeSEiMxcEFjb/i9571IlREMihD
jD62iuXYV/b9TlswsTnP8V6/VtBeA7gNAlHBJPPKr+tFnCPYlIfMiWFpogFxvoFSJUIkL0vbZvpm
1Uw5vF0jKmfSZhrFlKi2M51huaumwc/aw6VWuLbtTQeh/7ZG+EvsO57Mb2kR9VkK4FXhuRzd1lQH
gunq/w+lHkOJJ92v9cLp7JCSG0gvec4zXXixt6GkpgCWCVEGwbjkSnz13r41xysmzclIvj9iMojp
W9udhaZhgTSq9apEAtC7lWahUON0LLSBSlf1IKdVaED+wr65uPhaUgxWTcjmrHSIMdkcfIxzWPA3
+8am0h7NiNz9uvQUuP2qk/98nxNCI463pt3frO2bVDftyZoWuwUL6e5DwA8BGYDbUmLFpeK+TqK9
bA7jD958jxo2b13bhrwVnhr+nld7SgYPCeoClUGUsugwOg74m09WuUzIJLc5Junj6ifKf4l0VXdA
xpKqy8m2W9deMjy44u2owxL96NS9lKUzeEysV4HQR+zqvwu4236NEFnJ9CmHjPHPOjDA8S6IRUFx
l6XYWOhNueb+XC86APatKa2VZHWcKG8ql2IpoYNcEZ3c2hSyW5LqKtDvkO8k/LIy+GCS5pv45D9q
YpILmEs6PywPANPqo3a5VlZTcsi8v+sPJxhEXPfnFSZRXj8x72Mia+lZ3gMdaanDXAVKIGqzI+JJ
7///3Z8WH/HOCmJajYizN6QJ58+nGPGUiIzAS6j3gQ+QwALLRWb4xUDPSCPReQrnKq9xlITnBUn0
WsI0VMaqXFxoHnkQGHEqd/3/E1UeJ4nlslM109cGyAOxNTXFqiTk2lO7RXwXrHzqmD11ZGqC0yhf
R4ethTNQAvTq6aqx+qDuF55GnxFK8Q1YG0UA2oYg3Zp1XAbn62gTTBZFHkZiOqVcO6LVl6p46N0J
3rsxq4WiXnwJDQZgvZTV2/1hN+zXeH04mXjIZ8wYlxxD9sS8gRwiXndBLy6nSKbZDP6ckn35k87v
4uCkUOLvvw0MmvIK1BA21na/24EylxLu5A1m6e/MBtnIu5mXCPbsZBqG17JpO7/koopO53IEKMqR
dllM2shfXZpb//wTIbZOzuO0vxvIqLtihYQcow9AygvD0gn0+tant7dpO1jIHE/5KT1AweULJXAE
GaAKwjDeXKU6JKCgPY1MNkIpEH/7xLaqiBAZrAPNDWzl1LoxpbKh/zsVM2fuKg1jClfPViT0ULnq
GAvRvC2D6X4vZ5BZgAu9wSFtlZEmX778OdjFc61C3GFcIpJDFOz+lAo/Mw94TabTQ9hH7PXQM3uG
FRXvVI0iRG1egsie4vlJ3MPm+RegSTQBJuUALGrUlEpCYnXGB00PKdyfKpwwDCKTb04rpsp2cNnl
x0gKSj+vbby6RYWCyRpSSSjDG3cVDefCsNh7c5GQs4ejCrex3gJmlXfSuTiRF94++iY0NmjVQLWf
iuPYTiEU0ZEV2bAq6yfnXQx9PtjLg+kTKQa0RGNA0KAsQLCCVb4VfF+nIT8cTESWjtEIiq0pZqoY
582V9jbTwFUzH7lFq3nZCO5w7BN+1LC1ReFAPjpeRP7r5kwHkKgx+0WUZ8ofI3RwqyJjX4MK+GPr
p+aQ9T+6fEh+avJpGzOrTRQBwk3jL+UyAT4hforgB1hdOkwuxymhNw4ZJbXYl2FVBDPifj0hFkAd
/9esZ38bTMIYGDJCyp0KWt5Wu7KAPAbm4YwxhNOi/fmxsJtzSJoE0cydYBNLBSYZCzD6A6fQI6+7
NI49kUXoLBSSqfu5tNgTJTFjhnFp9bwfWt8PVcoCafBGgKq9J+ueaTCSUbtDoUv2pxNkORvQ3CGm
/FKvHcdfm4KZCJu8nVj5FGMSKJtEmbTa11hxwg4VX5CvOhZv9kaPT2JE3pRQx0zF+nKP9LzYKX1a
EmffbumogLrH6SA1nr+/7tNd19ZepT3fg/VOEbhIEPG/8z6HHR3cord9SBAFw+lWpDijxPJsAHmY
hbm8iWQkf7MSf+zg5nK43rm0g4YOmEziGu83HXQ0VOqdSkGtzHC3m6bzVFSvUCmC5Kc8gxNCJVbp
6ND90L1MvtOScm/3uPe4NxCumpHyaqciMkaHO97kn4J2cPtK5ynNVkhQDQdRs79ZW4lNY3V457XW
zxrmT1gHV2MmaczxlLQCNFoTbUfOfE2yWqEZ3VjKVaTy4/NxPQ8pii+1xC0bdyA9A0UGWD6QVdi2
FuvxjQ4DTUkSavbaQfYScImcegDMP1rAFGu3SaLsJ9BKDe+fGDUvVFaUEcX355XAHmKxL9iBI/TV
Gy8+DwTQFDc7aJ/lRhmzsw/6HJlj9Yis0MwLaIkt8oWpQzbvl7UTf4Gh8ajpb2G2S4WhrqVGaAJy
hOxqMc/7IYiSMd1Ma4h5ANFAciPxsvvSYOfbhDegMhmdA+fEu+WPzoaAwLdpJJ4Zckr3RffKy8+n
6RAznvVJR+VhtNFYezrLpfcaG/IJMM9d/lIw9SyFDiTN3SS99wRArvVwF5xKgYBGf3cbn2PPZkQ3
qWaAGrDnn6DOJy2HiyPOQvLvByPBMYkAozH21HHFOWyu5VjNOXeEfxSzFOx+gl9kzHo+zRJpRJ9e
C8Dc9FPdRxUPm6mS2WSO1mhGdyKA1ClNDO5t6d2jP6fxhv4iTPh7x++csK65Oy2WIztRbFn00Pfg
pBI9rMSHxnio6q68mzpMSHk+C7nzvY4DSOi4h1oFi6bs1RZym8gLNTMjjA2OFBY1fx4bu3PgoKcE
Xk+6MOVBEsr3NVqdwFnDnJlIlFW/WIQ6lI4uAssxRQ9N9uCzCYOzokomyW7rxzn+CIXaTIXVcjsE
4NKGitsvbyskd5Bf2JKCwBUuKTlOED2WIkgjj068QxMi+E6TzgrLxJSC63VhfS0ekZUd90Is6r1F
AysC8zgnbIWx3P8ewKQeQ0freyLrF1iApvMuzCmEySzrHiy/oAHbM+Bvbuw3LR4I8SipM/6z7xw0
KGrA7AyqfQFawuXpnpR+ysZZF8jGNQFvAtucQ1xULDBJDmWVuptlID7Dpo7meJemvtwPKjtC+vSk
SHLEtdMR57MwA2D9LlgYNBhIIpo5ArhdDy1w9mKQeT29sfkhkA6Wu8meJgv9HXhaXsfb2YNTbDie
8tb2CLlmQRoeWIQI9YU3OXuXWbuRAEyWPZ6IhUm+fhhD74wxaV/AQsSlR2daq1uDxGhkdV+OyFCf
XOJmi5GSi/AkHbYBo747dTXBiYuijHHwh1+2CQ97/95g86OWFql3kuJPYkRGD3l8eQ/PB1JAWHoc
uI7keWhYCEAslkeOvVxucx1S/3d3Z3VisIzSoIIReLZyP8/iWEXPLAqNIGQZnnFkNMYTMqrBzD9o
FfJpMDZiKX+BbE3nceQC/WMngEQi+m0g3mxT5jgWafC+oGmnv/L7OHWWz84uqT+/wMzl9cwr4UmT
6MA8E3hKzrJ9kOyWG2LH3fbYy3FTJayPdKoTRjQQO9UAiLnY/ZAidMQjn6YellxdRdOvgR7IWxog
CRlNkQSI8lBxoGllZqs9urhUaEmihKVWpsj7a58KrqvFRWtPwnY0eEVQtoxhdhcxREyFzCvldSo8
As6JMHu8QS7A0QSC//73HpsfFkWKbY+1z7jeXxc6Lj+P15BpRrTOww/qvFoQuqCQa+BPNzRwrz0M
qwl3WDZbnDjbYzYGmRxJLVRJFIorqD4rgZavufTvKZPtKvn/ay89cJUw7GmaW7TsrKR3skRDfp+e
0xQN+bFSpLbfe4qJ2iZErxO2b+b31RA1HapLCdMNBI6gBpyCDc7dgqSw35i7hXj5e9gOKhfyOcMb
bBcWHBFDHIhIyd9J2x3q9pLhCkto3Scqy8VpDwrT0ML9yYqxq0zCLNGYqNrczctHH24Q8CURk5f/
YWBqlssE1EmOs6BNe6eVjGQWNM94FrQebytn9tjESIkpl0UMPHTxJcseHOmI0xkxVaaOyIB3Hihw
2SUKl78ZML3VEr6rej0SyEMGiQgFLKJM3r2/d/dXEwbnojs2fGIE730ahsCGuArE6Yg+I7nx6ZnB
uOHDM4CHVnTvTE/LqaNUH87nDWl76GWGGpsRuY6+vqLULFw0vDXYWnb0EZMVURMB4Iy95wsVXfqP
eZoktBg0WCNfFaVZywuKHIIgGwtNRDZxsfFrAJAgZhyh7jOkQIAJqJhUaaXlScRK77k60IZ5pIkh
kq1WAOr8ytq2EO8RWEl2hAL2bXaMyn4zm0KnB9JIEApHlqGjZ7eG1kTmfVlU6uDJBiftCbkNh+yl
AoWicnJN+92jhTXQGj4SKZTu57K+e+KYGrAAhMYE8bAp7OolMtGjSKWQVOiVoLIUWhvlX6fTc7zZ
nX2u5XN0AXdrvaimlzXmWjk9O9q65JbKNyBoOY5wuqnsUSoS1Cx5Sc5WbOXMaR2kPjkb/kvDCVHf
m/SlD4KqsyC9bJqIB8yberaUQsgIvzPgsGcDraNjXd2muLM9gJBCosC984bcH3UG3kKDPLcMnQ9q
5hOPq2B1sphNSsYulS2icIACePYGYyy8Wr9r4wBxy0GuDcW/pdpaocEW8hJwnIrsb2WAKXNuL9Nk
qCklqsSEkCDKLUtyzbH2nDnilNvsmcAEk8rsY8zdph2E9l8czMVSnrl8w8GAnnmm+Oi68/MEG67W
TfrIT+4PhQ6iursia7+/KsiSk9is3Sol4le70/HHjSGwU20MPQrGjpYpj3w3GEOzdjV25bnZ4swF
rcLXJCnd/Ui/k+VwMZq6ELC+AFFDO5lQRFhBUNVv4YjLQdYiJjLx5bMwlWlVzrO4M3aFanR+mKvI
Ug1nTMZfdlhEHCp3YN/q2K6peHWiy0SXEAX4XNMkV8b5tTzR6iwbyUos0O1yvnQKQBysWmg50ozg
fstBQTox+O59fIGtzHcy1Se0aP9z1CUzJKO0m2/UboMDGT73BjxReCnUY4iJnPJVz1ezY44Bi0AG
g667zvgEOeMEepVYU5SX8k3HxyQWu78fXSDb8a+s/rngBDuICiVeBLZ7RO1GzzRZx/bkq+SbCO7U
U9Gisgf6yzj+A59fE+3Z1uu1pgbSv57376bIGxaRtfVBV5e69Kv3142z550Ci7mVPLSQWpttsyES
kRyST74Bqwd6CzQ/djxk+M9MVwWjgY0MiFD3ZLHcRu40Q35vAYpwlNAhW/KF2gq2wHLtCnztnZca
kzWIJkZ7SjZJ6L9oYCZLObGU2zZMM7VoqOuekJUiGcexdoTMcmgIOlWIazZn6bdWJIP7NIDteMvE
7GqlBLf4tcTIXgGhXztgU8A3b/E94RVC7M6TBHicAV1/OFTJFNdkJP57ppCXYHuGT0lD9dbSB66Y
EbQHD46i09c1SX11GK4oHt+PYDdwTyhwgrdPpDmfXSXHAR/MZbDzG+/ury/Kxn662+KDTsnWnbIa
eV8xyRdflCA7BY01t3EezUZNr5ctgBf9AHjiqdlZDNOC0MpkAv07dheYhmT6fNr4ZwP0eiQKa12I
MJLNCu5fTCokS9ZFd4jDJ4u6ntBb9zdc4JtqaHvRen1mSvFId09n1pNgeaBKYl/n13/j+Q2LCTyj
Im7hSrHhBGcjeHe34Ae67hfcxPF2JO1xc8p5tGBqdUKtO74IOXc7Q0ee8OkHhajlrPrSNoiyXn3j
L59UK+n3M5dlABW58WDXlnZvzSzUw1+KdMfo5kawZ+FMjHDfchKtnklA3N6rEtoiiaGahkolb897
bvUFPPOvMufUroR9/aFH4s9lwY3J9Z+JN7c0o5fCNlWyimj9ATFyvcyloFgqlq91W+61Og1joUFN
AiKVfWWS8Iy7EuZGx796n/QLtZnAvwReR98YYqaBpCZztDGluz8zdv278hrS012aQ5US1/b56Tgy
9FrMccuBnV61o1OL4gvkcxDs7jkgze/mXy2ZtSEbxnzTBP4J/X7T6ud/q7gy6IonIfpPfzqLZfVN
6l76U3ZMGUjwph8Y8OOzbOzUnxlcE50rjn+tc8CrbFbH90TvUe6Ow2x3y5uV6AUd7AMeg24PU639
3mB+lJSYiB4yADbEGtpM7lgul89OWmUK3f+L0gapaRoI+7Q1SFX/1uMmNd40DkUVl2mXO62jSplD
PP9r5mzuyXkSoiJGRlqVdxxp95z/GKUfqly/0bG04MO1sxiEoMLAoNG8cGSRdnVZD1V+xjQtaP4D
ZUb4JiMwNDTkJXEMqpY7PrpKHzvFrCidCPYzPRCTQt7dHgI8me3FqB3kFn5Ns4uKjboRlWPC0pU5
gxuHO7cTkMVGS0Td2swFKpB24WD1WETrYlp57heVePWALuo2XZR0XfOy3Q7PI1CXsQA9zoM74MCi
Hxh55Kn8HqeH7oriPmEMk/w3pS59y45cb8snb86XAqHjluU/5lWvtmJr+3bhl5taFMffdK5PnsPc
d1lFbbfAFpHFZYnYJVCA0ii1UOMXgCeTZBnALRRzt6Z0oDbHLGO7szVvskLmyto2NiLZL/SkzPvn
JHCUgHU5+U2Cm84jopwzZdUUX14ORNDCfu1hrWx0me++VZGS/d32Y42VraetLMNfdQozPkT1dlyv
T1KwSHi3kUG6zNaX7oJXblnnOggDv5HmB3zc9iYR+wMXW+VarBMZe6WLF/nNb6z8mXKdfZLz+d+g
xskgONfPmry1rKur8qnyoghZzMoTa1re31qklZrUpB+G/b6sav9+/YrECc1CvuL6cAk61IMPevka
Fu2MuVWbmUfbvluVFfXwUQtSm25MFnaKvaDAScwG0hVpLW1e/2XctRfiJ3gaBUM0Tatvn8xsTbmo
I3Rq2Io7xqIwNSfocmkEVQuG4otHVLJJXQO5WuCEI04pFNPfKzzlCkyxfbQJ2DCK2nvD/ywEq2Dk
doul3JYTHaLmjcqb0DrSRAOV8egRcjjXdTX5cGz/H7MAF2N6ljfNDrhKOT1Rrc/+pq45hFlN20hu
/xMjDQSspFF2uvgdGZOE7JI9HvY5Z6sk+ID9ozIxDgCnuDTGI60gSO1k2C9EITS+WAT+Ivg0gZyi
gm9t/PHz9k0zINHzWD8OR8maF47rxwlVELGEWRcEDzb0HLup9IIbN8FeECZ0kfjAvFfOcuy1Y4O7
V3PqHdzGfYfwJ3ZlJ6xSxj0GaWdJ+9wx/agSNoF4bRGBKTdclkJYUL/AjsRaRU9sdW4RfJl6QHQc
CNjVM1D2Q4YSc+SpqkGH3xEEZRcDr4IiyCeMjwW4Nf+mMWT0A5Vz5tlvDvSDmaMA/UhBKKmN33Hr
mB6ziPVjqgkL7ELUvEtlYntcvJ43mCnIEN/cl0SkQt4ucHRIbcCZ1JyNUf4z1mB4RK+BdCAv4oQ6
KQ427phUi7GdnQIv+FBtwmSnjsNvBkhuQthxaKPxaJk/j7cHPU0CgKuIvB8KcUp4Cp0IlvRtx98T
kD8mkhmgdjRs4rRcgph3j7yLlvJPM26OvYfhHN6IDWZ6KGAJuV9xAPPHKV1QgLxM73Q5bQQAQpcK
44ovAsD9m7nozRS5tUJFPWgmbQOu3uZ0XYpU3MtSqwg4BIo+MXKovKl1rJ+QeV8DTCl7m9kysgD2
Xs2ZGov7z9C1tLixa1GU2SfmrDCGsc6suXEXNsYbgBx69n5oflcNDSltrHfb6QVfIOW5whsHzTG5
n4kKgUxshn/c4ltr/wZCqsmAihk+VXw9qnc7+54DjnXzr6xjLVtb3d04H17fNo8Ddl7Wejjw6HXI
e1qOkYTbz975mYZBI8bHztVtVN8etS/iLN8IPBQh0eYtc6/2PXzRX8tgTf0UQMEBGy915VPrKqbw
il8D/eyOw/R3YJzSAKnHOR4lX77cNBKwCGvZE6s4hla2gXIgbJZoIiYCWb7APaqL+dnhOExhCDHX
MrTc9237+2LW+TNordGvVvcUdafJbAomXsKBOcQ2eyZEdoWO777so/UICXDku0LM+/93DLRNBhfI
xRZcsy91JvyB7oxdVVLEah4EtfqsfmDglOZLwNIR0Un+Shi45UE1UGoaLqfGD4f1DAITJYi1Ftsf
3K2SY5i71q0uNv+c07yk8s4Mfly0dhifb4quxy9PNJlMX0e/SXfVe0c3aiM4tpr/IUPE/UmwjkKS
GJraW8kPhcdmND5Cezwaw2wRYpnSWtL4S6f3EhfFM9I9OKIcc548oj/OsNeST3GZBYjzuAI7b92B
zMe93vBqnXlR7radgjsJ0JKb61yJfS44I1/n9fRcxyfzXFOFfuZ2rCGNzHavk6y2DKfyjOlmElF/
YFneeKzStlm+KtjFcZ84trE5d2ST+bXfR8MiNSObA6SgQZEeX7IJGJUc8TQ/lHCRgtGvLPm6/prb
WzeLGhJOwVc6gHiFdLciP69I7PtXCjdTYhke1omAQZbk0nZlOUFy0RMFvRy8UAem+rh5tzGbZQBw
P1eSp5q94j6krhZu9LEX+NjGTW/bbku/K934GNzadNRmRPZY91M3YN8rg4D+XOZL9oZbqjSIuXhK
SClvYIQ2ms4vHA6/fpBNRx0LXOlMTiBv3oqdEGgTE5M5Jt5SgFAZpuICWyuf+kpb7y++eeSZByZP
RM9b9iooYyHnYJF7XYPY2HUiVgH+QnJ0XWOQmhfbmFojxAx6VbjNBo1GRH09aaLaGMEiS1VJumZo
P0mmObgXStvGq1nxwOqnNJWuzBly380yWPFVbRf6qZYaYdfO4TzVFU9Tkho3mKNoYgPcfesU6hTz
J7JskJnvuPwoL9CO5sX6fEXSwPoSiM598xSEaNVKxZM3ZD9iYNqHhU8oMhYYnCa4K/CNczae3WR6
4AO1+OMrJt2aU6ZtL2KrPwwZJ6XRLZikETwuM4TasUPAd2otTMNMRPAFuFYTmgptUtrA67tiamKa
/poKliHxBhQQ/eKJy1UG5nliJmltzf91vNkT0/ws5k0EX4CJFhU9XihcG5hd9sTwh/gkTT1JQRdu
nF4/30/KB+ljUUYHCAXWeSm9Fy7GzjM7pYGBhqybZq8+aowZWDVQgZs8xh96Lud5QaBM+lmcvSJ1
pW+9M0n8I1oxHbe2UZrXI5Ix9UOupCnsVulpEnVaHXBxiI4OLcLT/ynl1rJkXkN6cgK1V9vXjIvW
KFOB9MoUAIgs0B41+F5t5IZLow1v5WPgPCpui2eQ2bRdFPNoSMFqVS1XVZ+7phukncWXbjfn8aNI
1X2DXWJHfL1Nb1e6Q66TQsvNj1d4d3iP4Q9SSXLomFTQpwP/fzQFw37cELGRsQtPRXEhl3ce27Mu
hj8b6vYvOxpBe0YajFKB25gZbynHwK8lV2Jhf/A2zrC/juKHL1d6/mziHeNKuZjfNacVwAUsuBJM
hgSQFAAZ7dAGoD5rpsQRgNtrnMbPYQhwFO0X3V7HAEskeBvH2jATaBE+u7jmDKX2SN1gwiTS8G8u
CyacJGiIeN0prHg8/EZRYBeP87CFp8tEx4zZ2rClqFGCau0gAE7whGlTdSFEyvCwXyVbdh4qZKEf
E2q55wm87aeRVQjtt/Z5B5gCatQNRG1VMWP9L54Qdywl75rbBMtdRAW7aBdQEP8yXl3F2gldETBc
5+rmnNLDtcwHve3xZRnZVG1bFZD72g3ZL+pwN5AdcPfO3GDMjkisLsaUl3oSxn8wH3NVmnOe1f8O
vGfqE5FJmxgai4gMs9WtAt8CGxsWOEmaKtp6itFg4lbkFaMKtO+YmJqt+9xq86/BDYeg+rkged75
uSLHQNi02SCZSHoMQuJ8bBRHPCX0kRkjte5ixfcEaZiekeZ5sMxCk8ckhccw0KfoVes43niesEs9
XMxOu1dlnS+bUFTNB28JMCfkF9rk0tKp/dlP4CqCom/L+XbX17/S5URCiY/7SKj2QZXP6em77i4Q
j8NuEZriwcw5GRIdIQdAavoFamf9ruISBz4cEgZY1hu20/eVWQRA6Ozll3tEnyG+XWwqa4ntvYtk
oz2wbjiHBCnAcUKBNPISeKSbr7QiJWU+o1GJ6qSi09ezGQuU+m/yPx/VbQBdr4ynZwl+GIV0tejP
3NiUf8ydjjPGbkp1Prp23dlm73SyJrUam+NvWcfQs2qGF1ORKt+p14+C3muwWeGu/qc2gXtKI+pM
+Zo6TFp9HdSRZsSWHPB0QgfhPPn4CizJE545OLFzyu+H7Vg5kVAKgI00hT7zpCwHMPpgTiRvL4WO
9aqZMROVgMhbJ9ep3E+59wOMfZXYXsb2TnmXHZPbZ7mDIApqrvB+vDPBpzKKecPznauG8Ppf8306
edEeiLBAZo1+IJ+xQ57CYXzza4Z1dX6RCTFBDz5pJOdtozCj8pYqhykeNv5GqgTfCngg4qyoodiy
GI+H0U7WqsnS3m6L1FtlYWrcCO6fINWe6RxadaBO9XPxDryHs9OcVNxWQLNnXDeKQGmnolynx9lK
UekkXL1A1ftwv1c34Dm+or5wux9YalUqn4oXu5VjblDjKjebmPJ7l26hFI/J31Jzizvxo3Cl5ugI
juNXi09YvA/XRWMDwpNWWTREBXefIVHfDQ3ggpf3w5akll4LSyuCkBgxMysbsgynjw0s1CiZlrNF
f4AB7n2K5NUZABNb2FJqbtsBlJW7dvQV2UiymgR/ihGEvE3Xwk6qTKaRJNaztFdykCL46lUwhioY
muJgRCNpln2grFAhAwMHv8s7sxg1ZxpERqKNDnBwF4dvH7xJc9UQDqBrW6N3WDMKTEXTpEolYjxY
YWGNrWE6wG3eCfYmXtb6kARicIbMh7nTmTBDxH0hZXh4PrVITKTTT8CbSF736wv+ror5CM80Eg1y
FBhHpG9ZjautgjecIIhypl75L2mT9IODsPPVYmQOPYgKczd8JEGlXhOyLN1Xo7NgU3sez0dY58kP
YDrZy2HmmMnWzz0ScRk62XobJMACFmaZZY8JaH1NcSZwpXr7obuVI3TTy3ta8AHhE5H5ThoSkgLn
zy/GgwDe056VzUP2N759tMX8L5QM/2ZSaoyhVKPMptYD/UDzt77lkVJ5WqsY/qpLfCM4bQfst/36
bYciQP1ma4HeohaFJkfbnEPCOE+UiBywgQduuweDulNCzNwJKu8EhqM1wfZrew4sSGeNNgmV0sqq
l3sKGFySRce68GbHIvTt1RCBBBFynmLjbJ4xTEn6x3VbPDD7EFC5aKeCSLpeRcPVby6KhVXR4x5o
dhOi2WEP+wWlwM/i3WWzecp0ZMeI8ha2CPxjF/kLo5sG3P8mB0PuQGdCitLs1cyW4Zb7GJsMU5Ow
rIJgBRHlubYFHrC0SRVZWbY9vyiMuhoRO92WPFuwZIc4oU28Tfa/xRkto9Z12t0Br1BumPMCpRU8
Q3w8mQj4QWZEvImMA7cr+wH2pKCDuN+tGe2AWAojbO6IRrhmLmXVx/cykWML8R/n9DjTGQ83NV0o
wDzSmCmXaXufp2gNZbWDfhXw/Tx02XIg5j6II5Y+4IJxqUlsAr145lQ0gGsGDsx8GXquSEgnZRjT
rxlSSqOKXgGythbDiGf5yVmp7ycwJTsbbxFaMDSEmONgQEmEMfryVO8YDrqA+rWnaqwwecZO6DbV
T4CYXkNYTSRd/6JwCNkGUgUAjAHJZNFbctb16YjFKc8ITWl4AgprFE/yzuUi3xW402UHewlPjotu
Y148F6jF2o1XQ6WBgwZ4Dodh+0y+aizFjB9fUjbSSihyVxv3Zz7UEY+NhYpYb373JIbzJ6ndRxQ/
b0ut8kh6zKRnPCGY8PHaEWiFAwfISms7eRf8AwzIv6xA4OjDAuZ4nHDhSj3Tg5iX/r8mjLjHBFve
InE15qo7T7uw4RJAr67rkkCvfRjZ5BLyg2MXLc03SV9aws3PUzUJtsvOJ+taegdnzWjcG0uIlQlB
vm1mpZ2HngY4T4gl/OKSO5xI7D6BQK9aJEt5pO6UWB5AIooMwpUFpmBf+L9NvLSjzXwrfGp4AmjB
TxDqnay3ChzOC/f10/c38kcJA45fMAq4eOfNyrVyJ0bemgbh9+1D3vjvlpkjnLLFutyd+EB+a7to
OxJ1DJldhY2L4QiISKxC2JvQ14nXP6wP2Sl5R0E1h/Wy+LL+XRJFvRnyjkjsJL+CwCmi4aX4rOHW
bEL6yqP66rB4QV2sjbNQdV+Ppzf0cRxnWwYp778puj1yt8AKiE7gufZYJJsi1FYukFM0OpYxU7Os
2/MjUYe6s6keH8vYz2n+RjrDcedBonEcE19NcAvuABGDdeDNo2t1Eg/oLGjtkWqfmyEoHQMn7D24
Cn5EX6EVhD37gvRQfLcyXc03ZCO1jif5Ge9+jobNRum6CKg5TpLdYoEhCGqb+EALn6muyBjm0JHh
4JDzxqLSVYRLWlfcwmZbr/dO8tY+vkpT2vK1h8rc4IyM9td/fQTzrh1+I7RbkXPINLJuSi4oURrA
5tThorqSbb6cAF6z1p6wQi/KN/MAEj/QSQBkfEFYxc42kMNlaKGIy0P/NcRoRcaeKmAmZvL/AUwj
oqqzQAaMYCFgpImMNqoEuti5VkcSxAfIJAtjowWRNIFiZZ78Q34oMWVaJH+8JoKEeXCvBIFKTiAl
Un+GunmhyJEYNcVFbvm4ImsbC9bu7R0DhhJiD1T3GAhQ3M/3f5wGngc4iFwmiP8S2aFSo9BqfGqB
wjBboIJ8S59GBVQ5yrVDipw4k1zf4M/XsnTwBq6bNUKhUtwSZIgoC9VcIqHSPpg+CTf6ekgPfSbc
gKJ2DW0T0rZa1pwaFcl17FaIPq9I9HL7KVnFdl/KykNl5HbCUkxBN3U+WfFHtfVUzCgNF5THK058
AiEs1c+S9E5BP6+XhU6tpYwZK0VIU9AJqRMhPPj9SlOTRXFkaLe82FaUMn+/UfqHbR4MMVBeUY+z
AfG6ZCnHxmU8WY2+pNjslFAo6Rw1YRsM1e+c81tm0Amfdp1zX/gFnoRQb61eObK4BrllGC2/DCKg
gqOfbIV+642TaQFMrIHlntrRdvImrKJFiGVHfHCQ9FcXtWLn1d78BDSPJ8e/slXgmHfG4HaHpWsk
TFpvU6E/IIKnzsHBXLhpHWQ6mzNBOGUZP652EZqGuztrbUW8c1NnfiHQ/sl9rKNc7bI0nytB20pI
HxEIi7hsJS7o02hJnm/nvF8Ben+c4652tEgQ0EoGIv2NsZwxrQyrpisJ7EJIX8j/hmfJV97CPoLv
KbuFtCh1lF5gaMGe7HyQcAm6vlZB8tFIsV1c57B5DFRrHifXxojfFig6h/a0CqsvgyMtAFEBlRRO
l4fojJ1v92yAsZO0npCNKSggyQ5cO3ojeSzFuUqW9OueKO92cEf74XGfr7RVSqW/CkGg2XTcDpph
+L6INIgVGN+mm5UQfvSDfd2b6Y+WCsY0cScvW0vjpAJS6YoLQwogktLwuA6f+kputRCoFEk2+rti
76Nr1xW6FTBaUYOMM+NKxMdEgqTAhQ+MeuTAg/+JfEXgzLy+CypMrGCNN8n/+ywjTXKkLOHB1IjD
1j2ZQsSJeUdAZ9q6LM6I3an5Beeu80hff62HltBsW4IHdDbhLY//GLk7JLNVE4Em5y0HsS3ujXeU
st0S6cp7Qq7OOZvdI7irfbYuKreF5N64N9EOlb42mXLMfCP/pfBC5KY5KjkbdRQ1VDfLq6RoEgDo
Kl9j9OD5dd6lZSJHA5thn3zig8wXIZiTtHZuahsQanuIb46vvWBCiEMyorVKhLrh47qxI2MB2rm8
kxkrEhTQXJ+klToCRLcSq03IeBzUhG0YG5/xc5xzcd5pIc6LCPLy7zNvJxr2p3YDnBfmxtXMzpo4
R9hHVzWFt6HIQK2EHorUIckANiBIDwxICvpB6zDmjVZyMiKpZTdQS6/bUe2NIpC5KNqqyNbsSFlg
rYVw9PDUzKSfJqLVAr8L4WubZC/JqSEKaHOgMTP4GINdXcI4f66M/S7tbOyGn9UVWif9ypW/XBJw
4AF5t8rVK+ZlL/eYaH2pcxyr1noJLnF0Gzyztp35d/XU5Vmv4L07eJN3O2skJzc9nP2erGyLgQYb
RbK0B78N9iAsxT96ktD+QFCKmPBf00VYkDfuZsMlD254YVqZ4rxbYTZlgS2/ChPfyFkaKk5+hFg4
ubKcTXpiuOR+cP4dwklJyLuREbRgRgzSmmdEC3rPpBa5tLvUdqGc/WZCAQrdx28AU9gBHzhBnXtm
OyqEjHUIY1KMTc9+r3+6NQo8BfhzWeT1v7P4FHaDzJ7nYm2wUZ4PArKHiGmrbErlhlstjXPwN1UK
XkcXbaC0uJy1WoZt0xaKbhVemjRcZ8xQ33iqdrluuyCJotzfyisAB3xtPfifZwXjIx5rx+6CYizl
q3HssldsI+Pbdr4GwicnkZmh7sWrcgv2X+Ms4eCUk6c5CYslSwbIDQOJx4o6pFG4d6AKRxFG4QD8
P5LWMP3aFlEnuoYJWNi3aIyYURitqzoSVn19eSPN38S9nEEOytNEtfpLLTfc+ECw0MM/G/rciQUf
GLTfovzwC7vCPcR18OdpKLA3oH5sfiT9IqSue4BxZ+ry6clJLrnXdmRSSe5ak91DcEqqrO4O3S88
9S/OMLyw49bWk7fBGYtnIyioxVlglMmVZPGxXtlwSTbyD6L6lfAjXw40wf+4TdQHHR//U7lfx5BA
8YPRuwAIZaBBseInqHaYtmYd+a03a3HHcYGbCzaXx4UdadMHSMAyLkam6P9wIjV0dBCwHMARfdeP
pSlKVlbj/bWoZvPXFY705TdU4R1Z8UgpOg9p6qciObGwmznO0/A0i5ZhdBJu1lzndcT68GUoDUiz
ZDaGrt9V69+8ZrWKhHkqO4fRkQfDOH2GqqcnxZLX4A0eSk84WfnMZelCP/qJW/koqYk+bGyly5FV
5O/0rwp+ArZjGhYM60Aez3sEJbcmZKe48hK8eI+IEQoZ+uLbg5l9QtJKdEvkaw3Pasq1pjX7FyXT
ZxSezR6cBneXm7f0DJy36adPPTN709msWB0cJ2nPTCPF28wFSI1Drmvgd6ikzcYbL1V7jIWT0F0h
3DBW/pNRBcYzr1l1lr8EBHYmVsOM4BqOi/ac9Y8k6VLi4H1u21FjVwAhG8qAHB7ZlHH8HJFEsfJ4
y/h5ZU+gbNoXKHRRfJiApCkznlx1gE2MyihvUbEBc8kItfdfSX5ltBSIkLbSArMA6h6YknpoCn5R
zDjFaF+3Qvi6Ajy6mgzBnNAewaD5LY094sOKGu0qHCrsKjp7xmzeqUCdDpDS41plOG1b1FBN7p4m
JpwyBfgCtTWjpK1DCYCKFoBjeaPjIlJYkVzt4qGd7JZltUbiRkNf/IS1vX7lF4VdvZaxBwamCkKh
DMfpbaqdjBBu5IcQuTbtQ/Pq6jSmw9z2E5+ZCXacu2PYP58Fgf8kdqMQPGNbX4AF/dau0osmNk8w
kwzmmKRHowvZV7414rKNDhKz/7c79U/w9nj71c+HR4esmh+DcK6zXISv5XxL2kbLWw2U2v6JgGY2
CZldCpa3buMXdP0RIDGWIDoc6BzKOwumtkXT8UltkPqzHUm2NjBbNaruvKnxQtg/1HMQHvbUcTdv
ovTF/buKp0dd5fqGnLOIwQ9/wpXiyh0uAN8vJKXd1RdWoyJt8l9Lrl54W0BbqSWRSocS+qDBtJ/y
TJ63uPu1E0nwVqasWZp8K+JfU09P6K+3cf1Iu7IC5oQ1vVVabCw3TVY0PhkVbbEJEClIVeny57Eu
Gj8cr1JrPbNiCDCf3qA57w6FaFNTV9r/FlBHNLLm42BSoz/gHz2tMBoAeo/phqtBBhQ3KtssIYZ8
6e5gs0wv64GMqYG7/QB5cpA0bweXpZJ28emRtCM6XAEWadu6Z//KTVPP8ZWTNloIfoEHwfNFuhAi
ivhRBm0c9X3OaRAQWp4y4uEuYaOy+wMie5MOGLkvNHdefzuTV0r3+TkFp/qiQ80kIKIkUi2jm63I
Dt3i1fM8b8IclluZFMxGgYa7JcymvkeHJicnix4DnvNZulALCeAEHLZmN6Bzpxuuz5XGiDIremJ2
pUMttTO1Sm04O2c0BclrFUVxSnd7max9lusROJL6LIpXJgJUNX5wtVsJ+ZObcVv8pXQ7pGWv1/1f
MId9B4CCI56ZMNZxPOOXXEyAY2L1hXG1r52Pw65jjseXCnaiyfREa8aOGK4Z7XnyQhhSjza98Yuq
7OMdBOADSdUSJwvb0CxPROmb4n1KpZzbNxsJk2JQMlhbrp+/+WgQ2u81Jeyou34I2ma7p5TlyMVh
IMIZo5TEmJTJnzJMVmFdlDglWdLvNFxxjqtjz0rh+moTjj6erUgGwwXuzXe+T2HJNJIKFJwPLRtR
RjrxASTM7yTvnuLePbz831g9Q4BvWSf5u8SuEaHXvBTVmwEHiMUCVRzuROyXiZmTSLJ0fg5hV31y
QlPC5HOlqV8jzFBVg5BVjIkTG03Y9nUa9ZCLyKJyfxNqxKxqkHN7SpWWsZtnDCOFc1G8cO3BmGjk
VdVv5TYFv52VA4uzeVGZwrWQNaFuznEDrG9TJvUqIKo4QDs3dP7lIpfuNWfFO7kBuMBzYpxPDdvS
Ek3iyT6Ycaru+HZhtCa6Lc8RyGa5QMiCG9AgNyWZnmPMp0GsD/qqR3+JUHqceqWfUZxunRGtZEmo
mVdBRqh2X/Jvudvwo/zYRf3ypDrGCuQXy3sxQIV0XmwbtJZfy4YbBkj408/xNQKCYgjfclsx2TvC
fqtrKWGDdexlntskN/xlQpH6eae0PqyydkvspaM0gion4Kx4P8MWN3WOuaGwyl/Sj9UVwk/VLoYn
olgEzmfhU7yV25N3emN8ByECb3wJzJDGjRIC/YygnmQUwpZkFZ2PtWhNtuxYZKmUZQN1MrLTl/Hv
SzthuqUIIs8lWzmf6QyNeBFRW4+2EWyIPrPukJ/ZEIw/13A5AqsgeYPpshfmZ7Ty9+m+Y9W6JXap
+i6vREHLo0yFXzHh75qH+s6qpnQEe6ZZLGqpHcEi14AZM29lZb9UiUvzGTbZOgSSqUdluoJ9MOUT
aIx9XPh8zpBN9LOtVfNWWuz/BSVOTxFtXwCiPAdN1TybTZQS2gEbMdHVthbeshKvATtwZfuBsl55
m7cDswqRpfRt5xuD/Q/NOmusI+1Zrh+l29Zu3A5XXtJEd7hB/YIHRqqSzm/Z8M6GeIeJN+mqO87P
eaENjvAmgiSpA5Po/aRX78242CvOfXNWyhndmMLWYGDZpwS3wKUnicHXXsOtawfdRx8E3nu6u2/l
Zqfe+xkD427/77XPSz1KSxGYfLzGJrFcTWUpnr2HrSbyul6RGXIe0qPdkZ5/UpkplQQrPPIHEcFs
XqTXZ/2azd/1KhovMbfWkanOzJUPp7sYgDFHu8lQlMb6ceJGl0nvaRqhoT0DOxiMOZj4FK4wN9N0
MS8BMes/fRZsrtf+qzoFhMlKrg7T1JuQiL/lEPKxRXX573sfkbysXM0ErvgKG4lJvcXBS4Wlap4j
R0N7V4VXVjbHCTKjgGULfWWEeLTSc6UV4Bjd8aKxGLKaCe3vytqW/YvVGxcvYIyvgjL9rG/LM25I
vPQawO+I3+FzZyqwScJgbUdYrp6+s8GBF0OQgTaxh3XmlpV4b3UWqjnHAx1X2WoBzGqLN43wC4zE
Px77vWC4dKTS2yTGAmDPbLPC15+YewYk6II9NtqxLZCUzGHMXU9UsWbAdvet58Yxk41NYVrze3Cr
3EX5nRDga1JrLaIEN4zdxmN4Aa1KFZfnZBaGW/VFnq1SOlXNPJbZrikdDmSIEB/WimBvownfkznr
sFWCwUS1KRJ9W0Wv3fVQ5shb85JqkRs/MsoJKB/1jhSjS6hPoKfpYQYiPAAYQELTQRHA7CAUEG/W
g3wcvII4IbhkYi3pbtW9xLJDhcIw1298so0kDDuJY4BD1Aeuev8ZQagWcitRL8exfTkzkeKuyq46
egfMMgiGhrJJnIw4CfdAKBkSQLiZzZS/Q57B1zYnnXi0+omjcs9ZlrWq2mV2G8JErJAhNYt822Nn
Q02dmtm3PHaPjlbvrA7hJLCBhSSoeGcnjsQyCDsNqdBAiIHmd6d1/MZgyknxRRGUgsJEnWsxdQZU
0aEjgdao7G9x5+BSVVZKkkMLuxdmPtE1UszJOC88PXnGdh56tsAVaTWXZwjIKduTCwjRyquvtIVz
mP8/jY71ML7duCpFdP9G2nEW30PAvo6ecb4hqtHwUFy4eiet+xmEXF8D93hlwDJvTTTadJcXqaIv
yYAfDAC8ckOp2g5Cpvc8xMJZECopiv244L31f7E9hELgCxFNs19EyEFX4XwZeTkKIsA0rQV3N3je
eUGY7TjIB1F7tiZSWZYfQEgJ80dk2gTNp31DN3nhR1zZ55pR06Htg2WBcFKrd6Bk3xPBZ6tcSDS0
pfPzzIHR8Rqv+vqKld9xaMK26iWKgzMlTaEo8I5xxiRvSh0llIzFPt4CPSWhWJU6M5XoCzykUb31
KLPVGo01NasjK5LCAHnayLJ9WU6fxR5uwIn58cP5JHA1yoX/lKJvR1hyb6fsUewrvj4/goBsm+HO
znAaJpTgM2uEheqeBSvXXcZSjpnGXIHF7meM8VlynewbIo8L0gRR9DEhR1nMHXvj+bc5Qo358giN
g0pRcIf08SSkaFiVIwp8j+VHuvXUGVqwJe0ovyDZY9Zx++yU58ERE4E7ivlE2EeSCxvzQKsBD2CA
GN0KmGG/IH5atUUF3YVVSiYoVfRfRuanKv/do/oWp+haQX/bmFIQCjFdtRLExbT7m8iIvxSnoijU
CCVLCJcyJI+q4BWl3ZRdOcdNtwgrL8kXKXzASqjjr5fwNU+hdx6AVnkAGxf9ITWiodZRvojb/l5w
i1nDnVLD1CSasemONMfWaoLObX9jQKWYCCY6h4tAdfw+B6CATjUo0lH7lOhupsXY/IfcNErBTHGL
EDXXAYZnKN+Oub/Dx43LNz3ZK/pAOWXzdAi6PAtbncBiprdtm6P6J2VS9DLjEHfG6uV13ucm5qt8
PAtYbM5Lq10sssynZ4OZ/RFcIbu4n/ovNpD4yCzzzW9rNqogSf/TCrBhz/lQWToRb/b4zjmnvUqH
GK/XikwTZOzyMcopsD/KktgttgZA6yxBfw0DKzCeVes9llOU/p1Uqle5BVEorMYAE/MN4Wa0d6wE
qwyDYa7ndTuRTTK9tdqRz8ovtIJXRNhwf5X70A+h4AZb0twVQ0HTJgMXhA7W/1YszzTRHFwldupq
6OfXISca/HsZK7KRtYnA12Os+wxHcT3EtihcXh723JJAkjQ/9uMgKaYl5LmXZB1iXz6D84wzqm01
Z8sUp3jXW8Z4bk/jnKozVrGVfwoee7P8dODP0UHDDRY68tlzkAczD8YDTyoML5N8WGbSpDF1uwCL
smQ2CmJMBu/l7hRz8gEMeYefamUAAidqNxiMYmx0QnIu8lW52CQ8+NDd7QohwbGc6as5sFhSNArV
CtJryjBO9I2w/UAPcOWlPNp4BXjlwSNZCpb2A0lhE3Y+/k33+F43GYD+fld8E6Qa6fjga1lFVNTW
5eU0PWehLQI8yD78S/cK+XdmLHUlILhXHObZj9+mcfQGlgo6Jw3EGsDyP8P+hmg4twiMtjKGNxDS
voG0Ijgd5L2ui9PHfZrwRgvjbznCL1AJ8juF/mjJ0ivR5l+KfSKaQO2DfXLLHeZ+lJtajBXOfntl
jQG4YQq7bEdsyOONbcowLMNhxEw/wWJ8vnrdgGHVAxMXoha5Zn2lAqm8rWyatrJokbbFTWFybPfN
6OjNIi0FGOgATh0ivJpSC82IdBQTH2zygsSBom0DVR6dUY1i7+LyQF3P4/rbkoigA5b2yXHYqK0A
gPGiqf3TUJ26ocEDARoa6k0Xc43moC1XFQc0RiV+67XrJcLp6jlW4rfStr9N7JItNXlI0VIoJ/VG
xz3178lKTfixN8Bn2DxMmF88iYAPnd6vkKiuCLa/2uZKZ5caMMVgaqMlaOPWwaEnQD5SHtCDzO9V
4iu/vvvNaGhsGDCns+06jbnpI6QA1SEIyu2vNuQU6IuW18jeNyzHyrFe2w2lREM5ggJihAZhGHNX
gF+HR7LeqGbK1ZWGYH6/NT2EYm7FykIhdIDquJ8iOHrJHXQSvrh4Cp1dmz9U2kEtGsDLbAbBUPfS
PtTLdYbhCC7OsrsUJG0DDI4IyszJMZQOHsQTd+8NVPpnB5BMq0pgEouZ+TpiRWgzGNTTTZog+hqU
8BFajT4untZOfHeB5JSYaojA7/ztnyoOtyAcgBgb79ZM+oPE/DbKp1E6UxhbCSlkILs18mCRfBzV
qOvpVnzYvLJZRK4MkExDdEcbC3qDXL/OWjyTLntt4dVCQ/N11X26M++N4vI6qp+wAuF77Gqr0eTp
45kEuUKIipUcbW56StsoIIaL2/vbZUvj95bocROskf0w5PQiC2/qczhbJLj0PWHIFOqcyPRwr8vQ
KS/wzkT5C5oI/mYebSTQRhRwojgEHIL0VDfq2+6W0KPYmGX5Cdv5P281SRbjgOuGaJgs1aAarAhW
MQYtaYO4APbNdDXmwQkSJQCDKWlYvqB8BOdzSdPnFNAjdMp0r12MGxzhkhXrwjNCM+H5VFh9y2WG
Hm/v+7FLHIkvHysyR4o6QMKuaNQP2vrZ+dL+ngRq5ZwEfua2su2OaYW0UobEwA0TkhsIT2ITYDcD
8lfFS3OGNGvQ+LV8mrAV0zhXiqEN2nbaPPqXbqJdcS1giUnNa4b3AEAp/mZb0FiovssK64cY0Iu0
7wZ0HbMSFxEn2hDlxeCFb0fAS2YuMkzjtV+TXLRTFNUsuz2FZSpaH2hjLTp+2F3BD4kYD5GD09Ur
H/mw5n3iOpyrrOtzXryd2c0o51j+yLDOi1qSuf1yvJwf2pH/SNS7MaOV1IXDDJXw85pZWURVmwx6
6cvgJNJ0rq12cPvclWmDFXdxXY5N+uOlByjrss5yUgnOAT+fFmoZxmbqrRYXZtaRp82kWYRwDksT
+E9QEC0+0rIlWiJBp10sntAfddSMraoQ+KCBnmK1hUKqchlBB4VmpNtp+w2KNmRxRI/rozr9aE3i
HB0503zIiaQOfrO7ShyrBrRyLybFIrpd5/82MI7O9TRSqnXDzDRqUs2ZZXI9uus66aIPhim2vy7x
OsbGQSBaA9q8MAMGyYogP8QB8xbTBzQG4MlH/MfRic45M74kv/50GGFq47XYtT8zq0eDUws0krIE
/xSF/S30Xz7N+sDuZ77t/5Bob3L4q6cg3i/abB3pezTUzpen9PX7vJz5UdY2zjj2eFZ/lvXtIs+0
vx1dMV3xN27cWyURQxwxtbfnQB+FPphPZhlWyx78Bj29p08X9k1lJ2bIZBPKquJ0wo6yyrI/H9qu
MVFff9YYEbRS8/8gVcnPSy+z9SWXWZX6X220jTha99w+vf1FZSw0PJXEqMKhjG6zKekZvZVN2WcG
Gs+6rUXFKPgRwWs5n/zGqwF2IqsgAFTu2idRZ/Gi5/mnHzOMhZBjHQRbYCgqklK6FwInOLFJRUQ/
HKdKl5ONi0pgue1u2izDBA/SYMeLEvNw8f0gN5+Zg7JT1VfK7f7RLoFGPPuLo0Vb7womk+9yruQS
NkQqdKdgSenUKQfYZ0SnZUoBYfWuTPac96dumCf1Y3oizEXobRjC0vRr3DkKPXYETxe+ZOXb2K7H
w261q8/9w98/FwuT/KCFC+yPdJWh3CKSUgeAIAkw0EeFkjuQwMNgEtEgJpa1XpytDaloMmZeyc8g
s/QIZ0SdfH/j6URaUEwOW+aYETChgC60Ev4umlQvYCd+0AQGMTUWIrJrD3ZLYBB3TLddkWOQruj9
j4jgItx+UuZZxWywQcxxLESOAWtY7IQEjCTx4o2DREZV10bkL6IHa63aqTTeikOdJYrb/REyErcW
tnpvSsZohXVu9eRyDUXgO4UYf+W+a+8m7FTeNaVljgb7HSPDOHYXI2/CEWuhLBt34YWi/nJTHB7P
mutLgjskccLg3fHRmYFkq8uHpRg0Re38qqRhv/aKmh/Rs9cyGXXT5SptNxcZjecPDmMTbmvGvdE5
Bw7R+cvDTEdwQxHZLlY0qi+ovp7dLZZ0AXulgfs03bpmEYsIpo5QRDYoG/suihCJxbP3BJrUEF1j
PGSuIOIbDi6A6hTxLJf98yv98yin5VjPJf5lddFSe8tLuuQNuppmYQCloUCwIWfnTlUkTbrgaJR7
xj+4GQv1xO4fOOfkPX0bL4r/+yuqHuDqDaYLmoH2DWltejS9t4mk3kY7oeUU7fhH6zmQ2OXxtmYh
/gqmhaW7G7UtOLaLxDQc0aTOI13oNnyRE3BYzJe4pv0NbWnOBAMK8kbMK5UhuuwLW4d+5B/mgBKV
3sQnFQwxXcOP/gv2SocYSNBwUl8w+YJW3PnhtX13zGHx5eyYyiAgeSmuHENF0lbaXJizw9ihq1M7
CSc7VhZ4bpBjepkWuHmakWODuUfUF+9vCfL/CX0YxZh+kLv64m1Rlu2Sib1Bi/oLCtpFMgkrMBYD
LHAW60H85/Dino3k0vWGeNlhRKcSbF7eF3++/s0RvJAKZWD0aebSzuo7LaUX0EZ0Ea2LBysoqny7
Y5RhrdGCpe/HwdGST4udzn1/d7wyHbMtZcb3x3KMS6xI+eWXNriXYWwhpoFcEdl5BTES8buZN3Sa
9fkfNmZDutqFqjowlgXJmr3y/JvzTAVVNZeXdZ29W9hgENNaNF5QCYS41PLy01US0opaEsqLBb+j
K82Q+ybj/bu+y0UMI5+HFuevIndfbYz6WC0TJRYMho5bk0JGemPzyuleOrvRjHMv9Duri3DNZg7d
XgbjVujBLw81hIG/WZNegctNNxbv4Tbnik4G33Fz5Y9GdFLnWezOyHDkKnpuLF1XWEzzlEaUM/rr
xVDvbyhPlF1rJCPwmNsYZTHEFPw0je933Of0qf0EOSAblCt86NKABCJiXPdBMJbs+42TYjvI7JC1
S0c+IC3hnl3F2xMdXfLJxEWpg60bYXjSMaAbFB7lPWouUMmw0HbPSfM492AvjBXphMcCJiZuPrnm
/F1a1Q/DqBR5wJ7OvSH/BV4b9bF7wr4PHvTsa4c86DByKJjTr6ZMCD/mKW49MMq/vTGZN7KCI2f+
JksNs8z37W6sxMkMJ8Cet4JmBbMsltcUjLrGqFi6VnoekTN8fXIp6YtNZbA3WjeUkcrV8Hts5rNv
zWtsb2xsoe852ziCbrQMEFvku4IHAjI6TBnK4mqrN593BxxtNnI2Q8pAFeluBXobQOKhgYTiqYL8
yiTLN2toXllPyCAvci2y1m1Ta/+/e5udBt6m8a58qXr2c5mdGiNwVqyaAqfPDqvgFWN4rcpARB5q
EONfUO9trkNOpxVEXZU3ib5XWHWvhSIn/CsgjWYGVEdPhoTUwZFhj5djxk0+RrDtpu9a2+DGOlaz
6mKEhPZpQRMLUw1A9gnSqcMoUvllG0wpMlnVPSMSeMllmzwJcVKQzXK1OZCShRMckUaG+vk6WvuK
/F6zn5wNTl/ufGJ8YXxS9kotCNoXsdoEBKHjpb8RrXO+A//H+DCubDstPJ6jEDNv36sGz3ORUGuR
qJXEZRlDCK5J8sKC84/IbwWfiId1s6ef8KQ/8vFwPkiJE/ZkJtKmiRF0kyc/4mYMybqamYndiOVN
g1jmnu528/qjw/BA1ciVygyBztcXdNvpEiYJBDnhMpY574AdwhtDoDT1LjTR32M3a57M9G7G5HNO
5x/jyYTvkGX+CsR5FBnpKCuo98RuarzwMMJKCAQ/gV7tMwjMGlZRwYC6PImIzJDBbov4gQ/lvlYm
I9MoOKZUUJUeMEoGsTr1oHtyuyxov2vj4E9n/LYy4fAwWpI9aRuFAUIygMUJSyr+GYOaTjeyQZL0
YzV5bGTfChhrrs05Zbbw8i91n06QYPDp67Gf/+XgKZtUHcagirpzkeZmPzff0T75Fzimq+HbiIj3
sdG7p+l8DYLvFv+VO++MWBDnixY/2VIv01hRp7CpGtrnqw+WVxguF+K/kGnD31qQNuloo6DljmBZ
WqIdcsVwG761KmEZpHublPoHKXVo4Rkc50rSbgWvr1rDhjAysaKsSO4A7ySHKVMAca0RIIVlH58H
8pPkB22VSiJ21xHWrf89q9TaBbkKkeYEIGDj6zTZYHob8cirbEtRbsSkivlivfWa6lvexHt94qd7
0Y9fb37V98AEvNJvP+J9JoS650+6p9HEjoMlJifFSA8h8Xbwyz77XSI9j3YOc4ePLDa4YRdyIKud
xp+bra6qJ+ck2/YyJllYeR0Nww5ZjWfNlC2sRfEDxVBnfTdEDJwfpsP73JAk0HE92gzKA1xZ6G3Z
7W8V2XSdDfdh2oRl2bdZC7jhTAPdSApM3Ui5iHl2Ko+RXyGz89zaUdLVDb585a7RQmEjQeR4y9Pj
riG6Kd1dgQooCFSKbKLi6Y9FIwlE+AeLpMbWz9yJFX49OfE9r6HSmq4RJLwRGoVwNCkKxdRLOgQC
XyMcgAe78r9uPy7H5SDTe4EbgAw+xawKsl+aadyWBnviEXu9jzedvwlDFmMFHQBAIOYBXJVRS/pu
qDStbyiQah9k0bLOqjVM9LegMZe74aArY+pibghtk31OWomjanxT8PKCu/D+LfDevpC1/tBdf1uk
AEthLHYGM9VKw2+LfzBKfigDPI0H6c6crcUnWGMmM5LJxSIcibH7eVVggTFT+xzzvxq6VANzoZn9
31DSHzt1pLXegcARosyP8wyWj00gpfHDsn1ZaAO37Mu7Db5cYp8W5QXYl8pEJRdbwGis1t1RkTFe
YdSmQntwhd3uZU6rHYbAj1wE4MB32NRrjuTO9vDPxDz0pnXzYv861qWoyXQmHxCged9KzucBG2uR
arr7v0JqkTnVm5CttGB6tFyc8IfbHvwa5PSGAgH8lQsu0SVhvUeyUZn1y2Z8I3nPjSHRH8fPBOhW
otKlN/CBuE3npvLhebln/nr1oodgwuTi0ewYaPEqpzkhrJizLLcURQspQpiAi/XWCionEIoJymVp
siDzWaj0sDsmxn/gEbZqT6dvScV95LDrb5Vtsk0L5R9emPdD6WBHJ6gGiy5rfNWsuyx5Rujp06Oy
a0TfVZ0yP3I7sRo7MnUEqfU2mASdLiM1s6U07XBePNf2cPvo9gUKeB/tBtyIzTBEKbCAFb8y3IUo
c/BtMy2w0Cn64CzkTy+XfuXLcZjc+QL4YiOg0cJ227aFteJNoX0s6CB4UmBSp29eIDCLSGGkkoXn
DXRr7kPqEkVodeZ3ymTvjpOL/WPJEO9O3yx6U9fWh2J5YpEIALvPRfqSUFl2zFsDZBd8inNfZTz/
rqsKAREU9Q3tx0fgF0O9VOw85g+VFHVUu7kwtls/fjpqDdmiVgd3vVAfAkGI5DRZRZkN241AAKKO
5+tZMVVvoS+Z5Ar5QmoNhQS9fRG4W5ip4I3eRv3WejMJe8hTmlTVYYFSKsfVwNnxTR+AjGZEAP9m
DHnZlkVlB0gaXl5CvecevrP254d+3L5L6ng694jpHHMZLCbQnxJ1HghK9Wyn39NKc2tUYtoKP9ic
7uuJ8auK1nIWPLTv6FpcXFmXJOpl4hLOOOcMVxvt9lOflJP+JKgLZLYImaGnzxAR2h+W8ghqKORK
ty34AIGks3cIPnPaYiZVnONlnxrxAWMG0cAr3vwO9rOWySd5Pzi9Lu71tgxZGpZsTSEiLASAtOj0
bLtVHLRmMXyIAwfronGe3G+kNLBIxp8Buh/Dgv1iOEyIITRtMiD1yCjj5GgcIQMdrM+fLqZ12mh+
yr59hT57sUMfNPGUVKPTALcbcKzDuv05hK7lqtAUQ7KlL2btuvOaf7iJtX6cTI4PzMXR9iZ6Zg7+
H/jM57pFVeW3KVu2KtrXyNL3XtV/XXwwIICDGRMN/4w/vsWjXhrOtJe3itAWixJ6j5uCRIZVRnHK
uGdnhOCipdgg6VdOFPiJPeLoe/MvUGGq7Rasug2/iMheoWMelqUgQuXiaOgyjBhSkRrF/f4ekDYR
6MbyydiKIRCqt9B/09WbAHZvmZcP2DTmQoc1DNG1xo7NlAWbvUUBgDstnhQ5ecNzcVsivbsIu8JD
LEmjMR7rt/mfDMHiLKHV2oYVsX0RY0s7Ph0pwny2hbaxL4fs/DB3SuYyZpxqUn90A2yQkjeLPuMI
ihcmPGxom4nYUmJpighHVKBtfOaP2EAuVm5kDAg3eCJQg5f2NZpeJSaifeEv77oJKdyP6FkaVigR
vHrOix0pUgoWfp8xkxsZgGwk4Qyfof7oqLKBS5uwleXdCoxCS1BvII7ulEq3dM89V/FIvao/hO08
aeBop8OYTMfSjzzsHCMqiLEJhtr3E32R5GSDwG+0zi3+teU5KbXsC+CJlndxGUi46A44dUeOAWr9
7OSYfudb5OAMHM8BgSsxmHhow8elmJ72x9gYGGMfWEPTXo4uQWCn5xB67o1DzLXfR7f3Rb05XSZS
y2xIme0eaysQPwyHz6sZ1jr1YsrsRI7VjuJ7XGacAdeEq00uGvUqiZ4hvp+0A3GN6xPHZg+Ifl4H
Eu3SAQH/iTlNqgqzRtPhPFUUB0sXpG2kAiY9AcMc4VS76piKNOGVA4EtXkZal4lcd8DmVTqEZgjm
RPuB+Wbl8ZqLG4bJ37QgG5c5XltU4gmCV0anFEAbRjWHrTyWb7+YlGE8eP7h+zlheS71UxBTeAn0
2oMaEltXCQYBmgKfmnEZcuAJGrQoIgNxC6W0jr8RuwQemVEXM6rtnY23DhUTkuS62QIUloU6h+cp
MmvGZCnrGl3D2UE7sh/9MPBB3IXJ7C1hyE/SACcn/jfXOQHGpQe4jZ7RMLf1QySvFvva0q6wInn+
BdQKOobnLRFWGFCm27g6KTfA6p4Wk4EodRKk8VfmKfBaQci8KTX6h+gmp3PPFPg145fd1/IFGIuS
I99vL0WOUx+OTEQFrkqLtzAXlniLQ2KI7ePhYobHtUj3FNHFBkFIVLeITwjcOMxnn9UyxmARXlpI
x6Fdx4NZ1DkddMVtVBq/Mg6/8DDkpXo9Zbuynu8DRv2N2edvvDz6N7vxU7lnSVgQLOwtb9ePD9Jz
M6OrzAkKv0JrZADrrBvt0BgLbUpfCYtDdEaytptmNnj30oU+god4d7Q8BifpeVM8dT//GgkuTJTS
Jams8jlTV2kP4x6fDt/TMm50ORtmjRWmvX2RjAI6853K/JfyZ9pcz28gCE6iSrAr2zreEZG8DR6F
U5xJR7EnHekTDKBzPriNTd7yPdDZioX7o1Vtl/k/zpzd4F+dWKu10+PPPzGjRa28Vi/+lfjQq6iS
nR85OhFsFuE2KzzeSvSmmd2Qfe8lR4F2D8wuOkN2LVM5FUq2uLKU0hSwfHCcrtaInf0An3iekdqE
MeQFpLuo7tum+LXyKVplULgVGXurLt2myuW4dHcd//JnS4CHr4XSMlc+1GqEU0joMdEYdYsrW2Xt
AKp2U17QODTkVEhTbOExvsPGtFCgsxaC+G26ytSjiaqenpP/QKKida+t4zssgnrSnPTKJ7f+7wis
y3Hgt9KSMGMhvsNQBhnLs94Bz4skc38IVYhCmrVbEkOzRMyLitt40i0SO1bOmpkY5cgeA1JIOxab
sfituuClY4AmU0iBLEIRSw/zZnqFp6Sl5UDu5Zb4NoojXUoqFmwi88DXzVqyO188mIowswX8q5oC
r3NS8Md3Nni1/BWHNOR67hDlfgxewKJrxAi78RYcfQgPy2fOSLekag6uhk4SxBnDqkzdcxLopX/b
OH1WOtyYy4FUlZGFc+0bOoDlP1SiNoPfxSMWnFFGasMN4suFTBNVtHweZ8u4FvmhQtp0MNzIqb6m
Fi4KU7IW+rLae83Kboy188XBoTt/CnKjyOFuSbLEIu6pzk2YRPpWhgmed5Y0skaaOp5xvm0sfE86
DMLJ+cky91qpFrAwN6jK1/tbPSu+v87OJjCDKyYmV1GEaefIH4X+60fI+EknzTcRsf0DfLTPj1cg
TZsrCXAYesCIvZ/6/K4u9OXcXvnCF/ViDAQbPZOAfQg0UcOjPxtdrKJhUvSbFVWIeI/d9wG++8Zv
PIIHMw+IY76LheU/UFGFu+uA6sdRMylPtC50O2tclyESwz7rkwYqLQsSs+kUaPD6AxQG3L5OWRg/
BReNMWUzQNTjXzhl1cgdLDtbppVG8h9BxVeKILVnVRoHKAo6GOglkcf5I4GmkaUXrvpUuvZqJifE
MEWHl7/dZRb9reWgHUu3NhlYPb2/auDh7NYvFt2QV2Gp2G3KY0BcKxIlxtczXmjd3GzX4Lizm9OO
Ov0GCJONZ0CcAHmIfvQ/ziadAjxqkr8Poh1uYDIjI94XMDIHtAyOTnT1b0JZUnU+hGB/d5FD0pcx
pvyq6L9kk9NVnMVF6JddCwsnOE6U9vfj+nV2CIEZ389rfbGIkvbhIJ5soObuwsP4mIJx7cwLs74q
xHd12KEA1A4N25b1GHlN6uAt9llFFMtbwaZBi6IhIMC2wEc6fv5QXdmPCuVDFYiuSJs68HIGeR9v
7GJiP6gZmPSkMstM2qXFooOtg0/3u6z0cDJCTx4TcOKxM9K7Pq466z0ABT2smQAZHdT8IwamO0LD
ap37mJ05YuSlgNOoRYPHXYfru0+IHC7HqWs+SdRnuy1FQHYYtSM7s6jpNd0i+h0QTocCQNMlT97+
zkZxRgrNl5QsSJak3Lwqf9TZwMdsDzNQomVEun86feMl/f07rig9rrBzDPsKoAJHADaJMRJiibkx
/uld3vDu5jjmM4U5zIRTBgP/aXOTth9gzetriguYV4WRSSwj2jtstuc3fR4G5p26w6NWQkpoZ7b5
RiC2pySdblsbrr5esTSOffofIiJRf4f4OP9LI+afHX3YxqN16R7PqSrJyJm9zR287VGqFbLfq1gd
bWlU38dvqgbv/7SIP99zls1Ru+q+1Qfl7Cd10Igl7hALrQXgu2Z0Fzu/8rLT7Nj2VdfNoM1JRXF+
VvAbITSOsBV6Mr5Yflbn5H3AGwlixvbENWjthTSOiyqkTEKV0WMbv96JSN9n08OMqj7otYME4H/6
E5Wk8dKzXbc2eZNjEwXysqDUfIXVLLn9r23Vi427Zcabck3cNGKRElBLoYN8Ao14JNcwpT+nbpye
LBr+ZeJlaM95Ni6BXO9vrgpSTkK+AmKUnGEtWRZQ20eDsUtjUR9O1nrG2iX9QD5vl0jIKvG3u+Hy
JoSxgQkZnfZBZkdUwUArssBuR+e7moiJrhraCWbqld3Ju0Gp63lYQtgxtyl/ixPP5fPWZI++blKp
JnFkdYi809oTjoTwpd1V+a5/CtSaZZvweZcCXHKqYf8Cqku8NBXLIWQp9ui+k43t7vMfEwrTVf6b
fxrHKY4dTrTQ97Em6rff/RAD92S8CE99/zSYqpRCpob0IrTBKJYn7frb5FmHleVfy+XHW6zCbNRO
Aybv53pnCFF5I013RNWoK4D+w9zFaOuNQ3lXnsN3jzBxVDLxubnfyo3XvzjQO2qkrB+ZT4N9e7Pb
oU8kuEKVfv2c0rsay6LjoSbJqTMYgovdSX1GoVAeXn0wX1q9H7iMV4OQO2HX2aAqGfL4AMCh2XxI
2W/eCj9xr/ZjlTbLbW9VulhVsOPFjP5GZFJvtlQl3uvU4YOv5NF6IY9rtok2FawAhodyCSKLkj1v
o5Tt7c91YzOrVI/MguIx3EuD7fRV5P4VVa5XaKrIK1nhQRDE8asOe/eSzSddK4QhDe02uEcKxdKn
juUNYm/HwjcSEU1Ha/BJFdrj2sB6KZaHmlw+timWWwIuM48bZI3XmR/rXhxF7iiYp0Ys1IajAF0T
KuTKeOJRtpuW2f3lhT100HJT9kbsW0JHCGiUzZrPOTsPAQW5RYOCvm5w+so06V6TN06QAcckqb0/
es3psNb+S0V6NCWQV/syttfhvYxvXzVJqpLnfQ0C82vQvDQx72dtjC9ToRZaW+susCMjJ3CWEpKu
QlOiBd8AcHdDIRLvEt9iPSGS1EJ3PUggAm4bhIKmW/zWDEd3515u07Dx9Sk7dUFmGpIGfOPSMC0Y
97dTgvCIEe8vcVMS4IyhfAHgerC00xAeBH+Kd7Md7c9u0JK2jeraMmV0Ahm/gVJ70u8sCg3GS2Gu
YYsnZvAR3LKowxmsnPf1fV9HBXCFyOVjxdmKGikWAWqKJDKW0u/YMctj8mvb17/0NHWlRV+DIwi4
YgZdDg/yp0nRmEWVdyicsVPXso8JnlGcGPAQHpSpcG8LxcJOvjGg/ncOR9DD219qRjdnB4T+DiKi
NsBR8ule2mLRl2zf91gdEUsDv8IadGsvSu7n2en7P7vRU9Q2w15lPMgY12aZPFFjx9IcSAQw43uv
HXps+FRDTNmglOcdZKDeflCQ3oOMrQNdZYTQQpwtkR4r98W+d8PHDakGW7y3H7gcgSJYOptEJsWM
8nwt9RxJhSetV6mAhX+FEqOK7XGygvAYsZqYGm4wCXgG2aRXa/WOXfTZpdNqK6PMjprclgTymFOk
Ew7QGKDvNBZLkjBv2cck2W11yLkXcmrWoq8rS+2wjUMzq0S3fu5HM48cCOHeZMYVrx83QxAkmVRN
T4NAn1RlKxXjmrW5U5GD6AW/vWm34+TDVTIbx+rHhkjX9CG5/oMdwyi/J9UR1FYMl7q1AGvJkI0/
wYY50klByZ4yyrtd6mN2NY8fXl+y2WJA6eH+xji1cOJJSaxzTAnAjUi5bWtO7CpmKXCo05dviP5T
LVJOXfwYfdxr9LgoOWuIiTttR1Jhysz2SFtnr6FcpUoXckbqEJiQaOe+D4HrERDhFQnqA8IKD22Z
BT3mp5IQEXs8psAZ6Em+XP72bnpPMy0Wq12oqh14iG072hPJyiDftRUyZA5vIri2CxCdT5xrINQK
5p4KaarlCvwu/IegqIjdOeHNzmYg3wJ2nUCUUHtjTdkBCRR1gMalA4AI+VtDoHNlIXNtAvrfiLp8
kfpIlr8ZgQiRiu6X0NWlJ9Y9pCTP4t1cVDnKRYhq4UFP0BUaeMCYa1yJeZSXaPywE1arOUoF+zcl
jsNrfwVAXJJQ8vpSOtpin8+RSAHzkdeDp+UjqA6MmWibvZTAGI5IHXvD10gpjRwm8p6mi60fgWR8
4uZ3XCkQWI//HGGAisCPFfu+skPfLKthzIjf9E+MjPhDusgRzgVpMMxej8UT0vixJwn5G5XivntU
jzlu0gMto+mHjaRrYQiFcsrbR3tXhMENdf00qjCtStf/w35Af+92oM9u4eCqBOYZ6xZ9kN/OHQsb
kJFCgKMLSH/r34iNJ9igNJWDM6Re+KXu8ylTZ3vqjMTJr5Q1OvulzOaiS/y2MRXpjkTLstZtT3cc
1XXsvwXIKF4HHCspxh9PlbibMpgKltbnuyMm46H7EeQuDyfv1FeHmCSK1s/acpejL/YfUI30ht3h
o/Bz3BIsRvy92qshmenWZ8zazVtHR8C99Niz8irEvnlKJkTnZEhnpD/rAQS/L6Uc6TQomFWUxctB
hR5i2Jt16HqvEHqBNr/JiMY7ZKt0akFDrMxRK2DtIm/67cv+Q4Frg/X5nzV+oiZPE6V35lKddsXf
MEjQkmG81XzfCGtD2sPOYZ0Odvwd8j7kzAZ/y21/b5H0mgOV6yta9XAq2J+UzyFvpVPHLioFbds8
IC023hbYQmR+PkuXCCQ+9lm8FkMvhi1nRMkyI1dj0If8vhSd9c7Ip5vZf0GSyZZxG66mLgtFHaH8
tz53pu+mHvDewY6zfT8NmvYJgT7F1oolot+SUbcayAeMbq/QFqN7t3UzJBsN9svt3McnOpH4Vs20
TKAWHaaekz40nSM3PkU75/eazBFIY6ubj9NrPvBlzKvNOuh50B8yrCqxS0ukOPB62OWx3wY25LBb
frPk7myWoYFkUElIV6215+4OhsIncYPRKwYzOJgnUkEygOfFWPIhDifs9r7BeK2XF12gvopnnvvd
Uci2hR5jh9WKL/vWSIw4GExxzLZQh3L7bv6q4xGF8yDStZerqybaiByaUg1D2uGVksYu0+ecQrEG
FW6PG/JFOl9WUZ4ab2M2lb6DSnh9BSlU7jmv0u9sNo1rQBcQG/8+9ZQpZVhnPrakX0UxdBeKlAfn
QKjIXQ5PrrQtH0nio24XQdfO99eiHMwQtTmdnAMdwBR6I8NgYj3hqPRSESHJgVnKr4ZweVySU+VO
LlEUJKvIB1q+hSjFewb0ho1pou4q+UrjBOym+81cpFFk7fvUYAyYKDU/DcOcBxvIAlDW1+LC/24e
0bN+0Ht0VASJx8vO8nMwiXYIzZmYy/MACa+CV/L/IpcNoVxoTG0DWxlhEIEv6765H3/9oQaQ5I01
mqKk20RVxBk/AtSpU4v/gDiCJV6a6POkQlZkjCgycp9KxMni2Q9fNx4n4yYcTFdW4c7D4RrDyB2H
YriQajO1XCYmb2KiKy+a4zYgB2HlmMXMe5iDEFB+oXYzJb5rYwR24vbyTfrhsxgPZ1X+oS1HbOHy
McT2V7kPe8rOj7jgaF82xMUGSA0Yo3XYIgoWAM58UJyiHngEYU3u8OYcrOHmegWyt6qa4FTAz85c
QAMovac64YdI3PaBPYubHep7zDwReX0HGjVzEneHmcnsFBFHlP/VuNH3r1rCSwQbagjV62vd3JnN
MqFfMfH+tj3FeTFbUhZBRz+MYDtr0+gl2etOxg2AC+JOr/t9ewMWUK+pfUNvMISwBgnblt2lTUaj
8cNm9K59QfaHXxrpYDAmfOCiRsDw08/Boi4ieNE8cg326y7OxJKiNxum58sF4Eb+fZUABxsTRYUT
KKmRaO+xfPCS8lY+cyp/ApqizqBiCvsyltyvxvtvmzYrIA893So5zOrVmRk9SDgfyu/Ecz45MPJr
2CT1hbN73NeR59nOKxz4bq/psdUftwVR8N0WqYQKsv0pPewg9aUV9MZ58FkDlx1kSEz8jHYgFzqF
EwMLxzyJHy/3DJYP2DDNJYwqLF+k8bldDQYAGdKsjL5DulDSlNbOeH/uLr5foGgYgaNnAvTPd0cy
ZlA2ffNKJa9QzVIKt8v4/LNLnUgnYhLNa/SDR6dtoGAOvXlY9mgVS2n95s6fM32AzikWLtrt4bMI
cOzwexqdYXIWW90wK3Of7FN4j4nlFrJMdzm8AA1JnMsqTwKxsC54wQkIBtk4BMnd54tyt7Z49VhE
mNiNeI/SQLe8tJHx9+3xtHiHGb7evZ7Xc1lb24kNzuHV3xYR6J1jr9DRb+VJDNQVaV2ARuZn03xC
Zu6tk1Z+uvigY7TNWXn/RGm4mR2P1lYR0Q3/0a5AcKOtPMRIkkQ0/TSQvY5238HGxUgmlHvnuYpA
OwqHZy+aCKcQ1w8SljDiFqsr8RNj1JXCJ3930fFKH4A43EOQsDwdzMfRLREpaVPbc5V4/gatruyd
vacD7RjAy1XK7KZrduttF3gLRsBNA7hlvvZc5lglQZN00LuxX5ZA6AmHhw2SNnU4FOemu/K6u2hU
O2T9wHLvPl1TwaDcNZcmXmeNZ0Bx3+9W1iKXnWX1MllArSonBZ7WzxXNdm8EiCdEZXQ6f7D+iWQ7
cfqcXVRsSEa9qGeFia5OYaGjwjcuemcZ+fGvR+tzHlEehVNc0Bo+fLSl2+9XoNv5VNocOjKCsSQj
rf6flaKDcnTNF82k4urD9/Rekvduw/ANOeoEFnsdQezPV7ziQmRlLSl/lC7EhgggbHcaij72NcBF
btCu85xVxMHSVQq4dtzQ15sgvC/7c5/LNzJQrjoMZgTzt61okEx0kvmQBgV54kifOPqd4W/O97wV
GB9oopQbcQ9r/4BnPxhgaqUw4ySdlo19rhmZOMY1/VVk7PKDHF1A7QfPtcM3OyTBJl8DU/TNg32l
eMEhW4jmm5ZrRMqCX30VHde7xjFYtp0/tY+cgx4kXmcFGtZVnikC8FgHosToLY+P/H93jaHzpe36
C1C9JZMW6yk4yNg/QZuFhdfzTFS00GIDuIJolrU0Gm2S0uxdL6HlV8JBxCcUFzs5+UQeFwhZNpGr
0zNK7JwpHsFqUbXCG2OYpTL3L8dUAUPAFQDV8pxald3NS7JhUJFy4imSTYoJLRUCUpThoUwJlaB7
rvivcPqNKkAuzERmfbpN2LdYQg95jF7DsXiS9Fq709ivva8L94cZabX7TazatIdOKFZMRlf8Uan6
xoDp4FZo6hWQvrHWlZ2w7QYYfB6yr9KrLWhC9nK0ET31Gdi7bdoI9Y/SVNIE371F1RcDVu9iCvfX
95rPnZJA7qlE9Qvu6ewmqEn9GlRQvr/37qwLnnGLlRKiBcuGsD3bRvtTGuYR1uJ5xXf4vzpWP76/
gLVovz+Wr16PGZUAmxc9YFxPxSyf9fLHZ7tvPORVGjHBxGWDTcs6Ev94A70u6x9T4T2I4wDlUdmi
bu/goDpAnazdMF+CWl5x+0jLxDejABcAo1L8+SlOrMvgqxn4ncIOQ/FJgr8/6b8CofJ7nU8pfvrs
dXVkoN1xHwOB6MerFLSKNCkOY24WP7I2VLjRnZl8L4pbRDMIHMMXEIG/7lAiCcXlCaD9koHBfZF8
ttaWNjrB4yQCH93XdGduV6MaNz1K4QIQjuBQjunwLotGAxpD5tx+neFdk/gPJ+Xpl81XLU5yWchg
RczpFE5xcic4yF9t83s0N+zI8kPl5tU1aY9SCEHwqYeR3Qvod57w+CDLhP3HQ2ttxWFzG/0ctdYI
6spgbz4JJaeVtPY3dGUDJXQ91T2kBv04XNEWE0Gu7xDlgj7kLnxhGDu406GO8BHkoeCLBNX+Ra81
H+SsMptLIV6kAO4hIttgfADaTI5tWDUV2EFveM/rZZOHcBEdvDbjWOHTlh7NxQMsB9xWCHynikEv
CMD6rOzsXNUsTuBVtSs1udbLAmxDoBIxwRnWVqo+GLzGI0sSplAcu7uo56sEJwRKVVHoKxtyj875
BIvLdigQ9uXcwvo7sdDZfdqRG1kjiVcGgEhoqb/W56u+cCBBbrVXMsqXSU/TtAdniE0ZzcxeUW07
gpmmduwOnB/sg9Htya0Z+QUnY5LYUqrks28juPbjMx/hlCNHvD2FG6tBTJ8eL/0fe596FXeRFpgQ
vhKgHiaVF6R/EgcCgwIdnMOMUr3J9Oly2+YxdoC52d4VtBZGvkvi9Uo+J766DnKHca25amunC/XX
LVZuRH1fY0AnDh3H1NRQ48l7SSwALUtYKHQ0nZQbUDl7RXbRusjrABl3ARtYZICB0ubd7tppPWk5
gt9OQQjh2dO6r/3BKYr0/E/VfweJwzA21xeduOSfIJV9N8MGTwf4miPVSnvSkAOUux8+A00dnjjA
YLhKIGaneVaMdMMIl4RbN9kiYf0xhp7MVuEiy1LeiDOJXRjpOnR8m/338qcdXBpembfdGfrIJaqJ
jBykdzSbW42ssH4Ggadav6o95lUc24Z2QM39yvnTBqdbCSeDiC55Xlt5qpXKwpqT4t0FFYL2w+/3
XkqYOl1Yly00DwdjFQd5WJGTHb15QyPFVc7nRmT0SgcuV5JftTgNw11QLaUeQOov+UGeSoIRtua2
nLwRLjU5hrdTBThFGfCBYJP7m3ck/WZw7c5kgpFpdu13KedxiILSL+zAWIf+M6cUiauVY2tL6ene
y531wem+vpsrjDJelbq2ppRmXNUOtciCwXvnZRvfS2Ze1wkCPGK0bYIWss/eEIoZeYhq6AV4dRDG
j67Qr+OONWP19jummVK9KzTt7U4YjTwVe/b5S6vj+H/ovsUhdohaUiaXtZAks0vm6HnwCtLfA+xA
O5O7XQ+OlrkTiC47CL0dJ6aNpwnKhIzkiAOY9U3an2YFJGtTFGzrcGl7N6D/Yhhd0qVtYFEljJ/w
x2RbtZpJCEKQXTICuQ2H5p2lnWqtpSyMwegzPVKbGSCT6pMlVswoKwmk/puiOJEbuJzLYnxKSEaW
nJZdesi2P2IHOcq5En6nmhjAnei6wf0YjBLKCr2GqbyKypBoJAuBMp7GmLaJiOXezgLUoL426xgw
m2+J0jM3Evn+1DCf6u5ofpecC52ZhaAT4k9a4FYOV3aROin0dOt1exFEkEkGxIY9CGjlOfkGWRpk
jNn3Y6C54UeFVs+BD9+iO3El3S9CCGj/xKL3/fsLldl06eboxeS9Eb4eXDdQ2dcafMZvxbROYHKL
QRSwUIy5QtYhkIwAYRdPKpOgiS45IkcCBVjWG42Xuztll4ORc18raLf2XBWwqXnOcVX0/T0wwRKH
oDpFvO88K5xXQIVCsSLdqqHzSS1FT8AAiLGudmTBzxiQVypkkPe9OGjpQbPjtV6X6qGbKWZykHlV
4YTzE+QYzTTWypH227NzmFPiVNAoTjvxmI01Z/9rvBbtUSY7on5EcIWwSzMnTeF0Sl1t0OyHY8Zh
yFRfxjhvF7MKi16k58dsaKAf0sLXs03Ne7deAPDJGaiQFbCVMrqprjFK4QLyMpoivPFOyPJKqfC7
RMeixdOcTvnHV6l2eTDKgiTRcfQUt5R9RVYUOOj4LF7KFa8dmn9LrlVm0drql+2FTUCouvGlsAkE
AFl98lKTr0PiitiPDm0Mwr3xLw7owwvhEXF0IlNimPGt1Dmp+d8ZURZZ5VhOKCZxGD4gpY/qQNh+
o1bp0cibywFUC+PpqZCbUjwa5WADUDJkKDHmW7gEhApfsy3IhvJbD2cLvUCejITh+T98asGnatb9
mny5ruub7Uzw0WnI1ssmbkgCUc9BsGH2IbGMy5VH7du3xZmfEY0r40p94koRIH4QpQFWSMaKdXf3
ygN5ePcIEbJEnXZPcFFUJ7KC5alMYSexX77DtvIREkyHkkx8ALGOf19dFW4dNmdm+evbDP1E1wik
1oXuOExMqi9Hb3aiRS2JFjGVIugXIwz3XPhqozquovfntdfr/NAksmJKXkl4Nv/VzmA+TdZIolX5
1//C1LxnnyzVojpGKM67xUJFcmTLp4HuhFuhtxFW0GOi44VYppwkxRx0gpnnPTo3KVG0g9JJajNX
dNdEBG/GAWr33feyCfH0QZEhbi7NFRaPnw4BiEOLFEcUQB/vPI+lnWp9FLuuydgQw7VNHOIpVG7L
K6HkX3ihq9GZsFYI9jS1FQgYzcohER3lgmYPBvb4I2EVQQcI08OWE5343cBeDHjmzN4npQuUY0Ae
mKKpchnpbEMwnIsYgQPLx1bmI64/qLh2zHktWFMbTTEJMww1tj64uFA3l41myUIS3v/Aoz7edSnu
XovIwxHa0TNHkcqmRcCmGtD2vIwuas3iS1PZJM5UbHDtcmAdFV3oIdaeNJSRLxCW//yOS5lUZJF2
JYTt01npyXlDybhAb9U4UqYOJcwX+GgTGOA2Zg7iGNzMgWSzp6n10reFMN5H/cnSUc0vUjLSGOmn
uJnR4fx/l+YiDxL97z/6NHBcWoafIv0Cc31VZZa5HhP9nByEMXcqFRtgJLOd32mGHrPjk73TtRPG
6DqVZsAzDyRy5HKuOpn2yQyFxWREX+HS70YhKAoikWbKubZ75vnGLO4J70fB7JIClQBg9x4SBmgV
20Ck1lgLD3PqoYacAk/hvzF6p6cRspiOmiTEC7TfUN46zoS7L+G05X3G8DehCEfbXW9tca+gOCzh
pafa+bdmvMlzKz87CzLttEEzEarGypfB50NbAsxHuNWzAzDAKaq6KfY8yccahv4aEhhQZjCBSN1E
PESttxTkogoDXkReLFBhRykmmpwnFBxJ5Y39XcgUoDuD8Q9UnYEr7ep7PedEplKJcqNrrBharDRu
jkv6gNVPXL64q/WI2NHvcuA+Ev62UVWPqvh8VhAbZP9FravXgjuaHFk/Gx0Dt7NqV8Zpl0NXGeKi
u2SsYZRQc5t7YaQDbe9Qtmw1BT1ywGWTotXi0DVP9XGa277yrAQ40UmxgfEqU/Ix24BPWnINcpLZ
KPsOI9PBeCFQ1+ldw79aCUlPUw37ACsw80g9Umh0Zbx+aATu5Ffc6NbA2BGxtQbKBhpf1JAR5nvN
K3+XZUjEHC/LbwZ4PQU2GmXUs6uitKRRFzrpE6rb0TOqKHZLCtuCft2kkHkjYoo+xFdd9UE4Ggn3
2jFtypCtlEUePCQCw9HuaAczKZhUIALz2F0zcnEY4rTIylmf5mKGVbKaGtmzOlOwTMz1xhLJKDJY
RWmHUtExlqznEdcpxe2w6bnh9ZloOXlv4e/jj3Iqix838iLdKHLwjUMZ7Vre4XQ4kDWJrBlYX/5B
UUu8H0awlCp4OCyKoTw9g5TnOXFAWyIGWxinsoxDnFluUadnWyLiELB5eumInPboaDRHIyFnOLvQ
PfPeuMmcEhF3KTZx3XD8JNXpQUZrCxhgac0RtxSfXQHyDcRwhUQSx0hCkU67TP0YTuEnO5FH9u+r
IHMYjMSulDFlYB8t1PGL66FlFQkyTcEbGhb4RDzbRDtTPdJ5wbco/jqFTt2P520fM/HY2vgUVODM
FRKxfwOFUo0MgeFQNxsXbmWnQ1FW1gECdNBae/wezv1yi3szN83S8hj1DuHCOzXjgRAgsINxWzFI
PU1uvP41sO5KeNi5HvmIZYxiJy1mXfxsb0bSUsFK8L6DMug0jcIiAQOdATD+RsPI2Hi5bjoLNH4Y
K+csHZn2ZKGDMFfGpPie7sgPWKyDKIwY6SvNkMVfldF5Kq0GHX6je7DZnvY65V1tdJsqDbGsTCry
cnJW1vhrnqQLOsg/DhVKN3kVNxBV7yPMaNt/nzCZgJUaNEAGJCgaZgKP4DnpBR4C6onsu3V1lXc2
lFhGVLbYWOB+Ak0IY9pcODOYpVOU32QEL3/BtaryexZuHChe2gFW/nk9lSV/I7SiOJ8N46kZPyRP
meY0a3lvyhfI30ayFBObnlMuMf3P/8PvQpjEsrIktv/nS+Ihz28P5qfB1lSrMtPJh8JlJeZWKIVk
EJqxdJDcXBudK9KVSJit18apjK0VEfT7m3/0Am0Vl2p/xviIlDQ0XWek6iMyssWzsS4b/xG/EkIb
AWtPY3WfaoiYZp3J/XAsmJe0ENVd0dl8BojSB/uAjUMribb8IBJh7VW2oJU/TD+rNmjHUraHpwvp
7qkG6+PoE/2LSJIXL/xDWTXiHF6u1jsezlTcfYh8MF7QY1BxTC8Yz5LKs68lgaUkTaZe+TeSUe51
zARCzlitdiE4cLlxwETFKI7RteTtb5Fvw8OUFQtLKRCcQqWxX2ZLJ0TIwGHq1q//iYPvSo87ng0n
jA5/tv+Frghm1H3q7gpx1EtX6W4EfB3UtJE9geL1TlXYq6K7Q7G63ayatcZNlthKD+TAJjA7IkPH
SOhpJ96GQ32FieOc8Hl9ahRii6k3MaTZKViQhyb0kl+vGIUH1fC3fVvnoMqRGiAMjfGDFUHZj1u3
NEqGvFTl/0kiMS6zuxlNq6zecvxMHdU5m/QVKBbg783zF1yodPrylpWHQbHX+Ne5JcrCrEnsQXaf
Owoj4iP7MKSZG4rfa68Kz1APqlynrK4FjgL8KZyl6d6tDxQBzNoqOuigTrrzmStk3a0GaL7N3A1E
l7GdCNo662YnwX7GUcOrFMtDc6p9EKyFbZl0PiymH5ubbXmKZhvr32Pgr177ycgriBw8NDvNkm6C
ozzcsnV+BHt3QGWA/kkaqQXAD/SJoQPOFwBKV6NKhXaCOimuTIBm6Lnou73qJgY1jJEPbQQMpol+
6GCyrdSOiAf657roJZuB3SAt95os/vfix+L6COfnkFIYm20LuJDytErwXs1OBpRkjr6rI+LdBWTx
DNuJ0LGc9wy/HCKrniA+xZijW6Z2BFb9HkZZZBQcCwrG6074L4x8YL5Ai251uhEZKA6b3NJ04P7K
+R8+ngUXBz9fDkgFLtKvCv92nXH3H6u1L1npCeiY4m22pR5M1TuylUkdLdxuKB/ZEaP0XZoBkYhR
zm14HCm7EhKBXZMRSRsfaVRv0teUz+P7hQqY725JTs2EBYxEssjHB4WiDfb+eh8Etp+hV309Pfb7
EfZL06Pv8wJVnQDW1lVYkzkfPYSjvADZQliFHj4FDy7kOoNLKV9pf4BCnOQ1xkDR0668qY7/WMpq
brhblVpti2HW5TkYi+DFRFqvxjxeNn7HiTlETEfisglcKXZbNRJbKkR2IwmZYLNzyr9t8S3iZIzV
mJHp8vWFtjz9ZELKwdjvaAtAEaOfuBGwOH+mW8mConnCZD1TsKlymaSzKTCLOVeztYxPHqAz+DbB
l3i7KKY5jVLS9TULLn61gmnGG4QAsRE1362fmZd0KzA/G8Ij55CFlsemt1Z5nLWz7MpNUxPZeqtB
asBN638WyLdjqUWoX+/GvwhRKlutzRRZPoGRIMjCkio6iov774Q7sLwOD9DvoJLliQkRTZqtYoo7
7+9oHdXc6V7Jg9YB9RRwZ2wnqolkxiiKDc05BDU9NPxiuqRigddm7bMqESqLCPo9X71MzeIGSEo8
cuVJPE46MICIzygollrLgmiTnEc565G6EiG0VgF3TesC40jKPfrd9PZMoy3msfUga2V2zuOjb2OY
YLV6LfkovBwXfkNaKHU7W6h7tLv2o7NP7bTDl84rnR1owE8KrE3G3PaOHeO9B+8Gsh23lE3oYz+E
7ppXbH/BV1hnKkXULNUO3k0eWqbapoNfC6EZA0rrhCXVW+ZSYe7VEd9SNdJrkJU++VkO/2P1J1wk
r5pBqL7OLotXHWKQT8mpUfVfDX0BoltwU7IvUPYJXqqDbDyWNsh36MHgkIrYl15MIHjHWH2MDF+P
CjTo2ONc5ib1un/NLRp1TjsLOUQ4FLUgpysxA4gyPph4L9L/kmAO0N0qvRYaUaRdDfrEjgA9k54A
E8xgzzGmCqKSuD1Q0EC/13brMsGudZxBeKyMNHukJAARv7jtrqL+2xgCO7sSZPAJvOacZUDkoSS8
ZwLbwWtjKI0dXLxQcojwAW9l0kwUgpNRkz7cCFQF78QOOMTVscVIOuy09RP0B93C1+VxEJtIitcM
sBqWzdLzpP8+WxbWF1iDz6CsHoPcCchX4z/RHmSognAyX+pSxPmwdifW8cmGs+IdPuMwp79NuoGp
xGYGLFPnfQLdj76fIEQ/6oc10kHXnBSVFRCDu/jOeO+VwyCwKdB11DcAGOSa0Atc7lDJJqXsUhrI
rij2OPA7ngeRp1OrYTBxoQ3nwhGtVTeysShqWIEJ7mkCEMKFdT5U/gvuZRJedkGnNpY+Yx24t1UM
TlnEGXFXK9/N0cVwijN6GYbuSy1KeuK8RLWZPiLJrHBO3+PYZJxNpzn41fu3pS3Cg/uDMnp8pg7H
l0BzaUP9onD6lHnJeYRjtJ7KLCpPMi3VzYAmO6sfjyDH243dXGykfxbRYBLZ74O5ky32zGikG8d8
YPUIiIymd1qcRzNXQf/a+tzej9/FUfmezrFdGETj34zr9TGMzeJxrFnXh96PvAN89waY2szxFl/T
VdeuSZxmibgbBo2tDUAgSuhxiSbfG39r3JWx28b8+c6dn1CxIl3idkDsT7GPCKgjBukY2Yupv7QF
yrcjqSfWNRyYFf0MM3TtzTR8sSJ2d4864SwAhw5yn1x6FO+C9kSkJQSTLLuZshgL8casY0P75wsi
LNdWP4DO8qxgdmC9fNr7XJ9nqUkmJJE6DFCUYgaiRecviIpDK0hatQTBLWvc3oYZdrwrAl8zHnan
X7/Em6W9VkpYPVWC6pM5IH/JbAS6nhDzmdDLS0B9kQpbYfJm+o8j+POlB3WUBd3oHp/c0tCUlxYB
sBf3B1cVPCfWKDme/Dtv8som7QOdipJsJY+/QhzHkeKGaBY69TRdmgKabTYZNLxCDfK8Ik9ksArb
Ews4bwHFbrHUZQa3dx+NGBUow7yuVjUVgk3Fq6K0eEmqYzB/r+1FqFJLeGUXuLOyxCqPgqrvRb/X
UuGBUccq5O0ZljJpQ1enfi4nMiR6AS5MqoZky0FI78udIDmuN8dDmXliwRjRjo2NPLiumorpR2JD
WRX1jRvK6QHQGDQ0+m+5kMm/M5bdx8i1J4AJpgQX/vizdNoSdxf2x1H5qqF2ERJsmJGoQInEIpkl
BWqmamycjSswxhKMkf6l7rdpESJ3/8bnHGqA2VnQ1Rg28MKhDAAoRa+9GIXd5DpvrgfRmt+QzuTB
sDQsFkOlYWdqt8nfTOu8Yh5c+XyljWJLv8LuG+6pGX5SmP8ISWB5ZYn31PNQWf0xzmnRJijtFbFP
CI4tsNX9giaHe+igIJt+HjXu2r1aG3US6JnrbfvdDCVb7x5XF7pHgXf5zSbPhGiq7+2wWc6MB1yH
Z4pthUoIKWC8i2WKLoFVGenbMIvBK/22fACNStdmFBoPsoZSt6uxtyyx1K2nTQr1sPUzAiqBMU1T
A4YQ7nFDKTiKqA7o49eJBqlF2q77GZ5YxDa1Ebj9tyEv9mcEpILZr8cgT1+2sFJWi5tvbjbpahge
MfRQdOE1JgpH2CU2re/4vcJ8Zgzm4viYiUhxU1CHo5b30/FjODZ4ZsyjL1DJr3YW+pa18GQgQgjZ
eL9UqVme+dsWO+HUmTy94YCNCOpKpV+ci8/ohyGt6GDqCK2ZCN3Ii2PFnkOMk2pYOLlbUPv70o4N
rnec6V/J2wBOuhOLNeXFUNKMoCZ3vfsmGJjBcYV0PPcySbOuOoZiDaskmS4xoR0ddJ5J6WuLGuXg
rKs4iP/Mb+yFjlmEHBMo22sB92+5yErAmBmZ0lYarwy58PzdS/vDhZPZLtlRtMGhPXZ1RIcsmQZV
4lUU1U7mq2Ea+mqp7GOLjoOB7ZdGJJqjB6USPNwdwAz30YZcSjaiBEhaTaHHxzZ3ExQ+sqb0d8GK
wC1qUJBO+dp4Kyhpoc2kaZhTOy4jOmYJFGRmoG0/XOseEIhxfeE2zKTElHiuHE3qVnZ2CzXiaGOr
CcbbrqIMRO6M6Az/52fMOsTH8lizj4IO9BIkwiPaGNq/ce9N/SR1WzKcUts2VhtgMwL43kXaIBLk
ihH84oLFZdxVGaGFmmXmhdHc1Kd6mF5Lncn3Xif0T8pNmK+Abxuwx6s7NmXkMjlIC3FPYeuYLK0v
6GV9mZAU2GONigH4rjB9FnM244aAyAF1MSGI8Ize1Hr9VdJ0u78hsbfgxOQh++Bg1gtVvxnYK45n
gD4C5nFWGeHbD+C+iDFVQiSWl2ceR3pDuRFLwXydaS63zWqZvk3wZwAopf52noFEP+5pIxrKM0vY
QDagPeZWedCFQNuqOgviNWssoYnEQXFpluJ/5517zKPK/5rWgO5Y8BcAzyW0u5T7ByVkVsW3jHBu
W8mfanaERvONvCnEd+HuMQPZo1cM0eYxzEbxB7IvsEQeh2cxa0kK6MPuRqgMePSN87DUxgEXJrN9
RerPei+/idgGfsWsBefS9xu2Y4LyFJ8ikbU9QwEVVCb7Ewd99BFNxsj4rppERL8jcwPPFlGVu8AH
ojwWTJ4Sj4cHz66am7cFeYc6mN16mRA6H5tbHy60YFxdksi5TUL0RVN46hRTq4GV47YXqCVJv/ez
YTyTYiuZpOoKos7kwYdFV3rctHjEJP8gbzKjLXk9u4ZY+6GBVM4mgQJeokk8HYdJMmvNWF0GjGJQ
vBtye0zPGEdoQRRRRf+2bPTr1ci7BhtsEWFcbYtMtCjfQ1rrIKUN83edF4JP9/msDm3rgwNBPy/C
a6AxWK/mtucgMJpDEukcCjaFOqr8PpkgfZLpckgYxvnLVVg1EexVYmUJ+FebHb2D6IxIbcpIa7wS
h8soMkWQKIwpK8VqujmkVq8mIJ/HZhdTZSGWpkmOYKlNEWZd6syMi7mi0cYPDOllsKkRsgpLjYLT
QOoSix6YmHCvI6/d/6BIbfMp0JC+LfKOMtph+p36eboIBwmQrEiqmJgR+mdHQWoi+GEkR5xIbpEo
USPwK2NBQWTmYE+irVCkXgoKVn79NDyj/0C+HgfzSjbIDQzAPmVR2MSBxQHloNCRwvIYrVJ0vVXH
cEO6rGTADbrWNAuehPpewNqTb+6DtXGkmbucnDrtoU3FFk6uJJugu/lY0xGX5oxWLflmi9iLehXF
Aav1/KAG+xeWBbVAB+dgwf/0nZYKMKfnWfHw0i8BDrfJZ062eyVr04sID1GCjDys1gazv5bPlveR
1VzRAjTZwRLWKKzdcgXPpMn/jfqFSBMuAJCMOmshV/FqoToT8Fh/Df3RKHFh4swApQ8AR8leWLdC
FKcR2+1/s2hkWmFrhRKEmgjwRWxITPPTDA1T4m1AEP5sFS+n3dZ70qRjmhJGfE5PEKcLbxJ/wJlo
+ejtHy+CV60ITUqR4ClRT1qxQuXffl2IzO1iligK4vWrmrqEkpLCMsz02A8sn2vs7uvpUWgwVDrr
PTSAfpeHlc2cJdGv9T0rUx1b5J3ZNhLEq4ZaF8NpXUThU0F4bhaiN09yfuZkgU7F94IShYfu7+xY
h7Vb+QjMZPKxqs4+oD0NaK/z33+xML8I5pcYfQU9XbWnU5odTU9iEz5rlm6y7hc9J1+QOYFaYN4O
Agema4w5wym+KE+GwIS/8DPZ9DZyajhY6hw8+h/Swdtfv3BdOsgLxqfUNd8tGIXwrqlFBaFSBEPT
IF+ErVeShHwLjvgeHsLuH2OX2mRbIdxG0KOQmlDFdYcZiAiBplMetQYyt0K+zQ/cjJcmzRGCTUvB
DJuzhQQ1QTBrLyZ/QR1194Z2UOep4FFsqzIx4ZRILnj94G2SwC4OEQsfzXqXuIg4YTCZ+6UCjTsB
5Q6Vtx5zuvn58q/zE11tUxEGZYiqG7acmxXFWMLjdJ+qMxkVacyCSZjhE4Fi5Y2lFrAcjUFS6fm3
WvtroUcMOm9EdIxQPlIlH6t/WjULxg+0unMqx4eYObyECtYS3BiGs5tX+GCLNwrbUVvsRUn8R2/2
19DYaR+fhIqG1iKlxR9NF99EoZdxX0i5KxvVkn8EK7i01uKXICZKnMHefTNMAZFYcy1/Bos+FNxi
FwNaFlI5Ds14jI1C3munYacXFPBKUE+A8qiuHEDrZS7HJLovET2roRUBRqSHEWYOy56sOhnLE22x
eFt1FrZg7jx4RV4PzPzWFtt7TLuXtS9mFn9hdBqwWFGCeFlPOUOvlKDmozMT0YCfmgyK5MuZT/cD
K3pv2CsCN8Gh6NYdAgIT6J9erzNh6S3np3gMcE8Pm6Yo41bc/qUfac+hzB6r9K2QwGsumCtWdNcs
cCSJm7Nnc2wl1B4Tkr125muYFAxyO6q6FjSa9QSSk5a5LQW76pujERBNYw9PXqcbYaU9eF1Ue5U8
TZnKmvGu8TElUBM3isJBgAQzr7BXY0B6tQ1JtfL7L7R9tC+LKZQ+q12A50uEloOiQt8bOmuJb3Ci
8+W5liL7Kn5YOnz8d5Qoh98cjEDuY5o3hNn84MF9RTx2AvROZ9fVFN+uXr7qMlJJFRnk1cjDxZYR
Eb8S0eDeQLI9GPcu0yv6+vF0kkHVi5b3NGPqzHl7rCASGVLpaT41vzaM/zQG38zwVWdGPj1+69ir
5KQhGOIuDt0CFK4sizKXHshLDTLxlTt5BkdOza7ztOk4M0vyhldhdkplUTB7ga0JeouwYJ0e78Oa
PARl9JaVWMeFx9jsW3D3z/EtgpcpwYF6IBHotl54gu+6ns4RMANIYYzPgW3GusD5bGgnYh0Ly37D
dU8qBzSPLQrEG0o7G4jXMc4ipV6Bg+ej+srtLFtOE2RFscHCbx2I+kJbZSnxr0adQYEvE3EM8azs
WdXZXcFtuNfLyf5WOUxedA3fp6DCwYit2cFvftl7WCHpx2sJBd6PTC6vt6nPhIIT8CrvE/bFlN7f
5eEvREO4hy4L9b0/5PsKuXgo5/UkjlYmIdequTGDXfAp2YjIZZUB+fVdPAQguCfjetc7FBWNHcSx
yRG9KmwH1K78OO1ikt97J+Ny7lx4O4OX48bbJYRTLo5v04fXdt0Jrd7HeSqgHo5hrSKuqPcDQZxS
NF/X7/afxpv4G6w02vUXqBr7KxbDPbwFNuW97L7uy34Gs9CUdMFNNwDmtyY1yppkwcDJwcI9Tpkn
sAP2oSbM3K315xtemwQdQEUoA1tTrrDft747M90VqZXWsqB2c27gWs3+dAU8SNSi55OA6vZub8HS
/cs6fSWGOb1mo7sVP0wxsmGqhv6PqRjhL1fWFhXbuTGt7VSlPXuGUA5H81eHj0x34PpKxbRqbXic
bhgwsmBlI5oBSBFC8slgTTdAbRsu+s/pZyoLBPrAtmqDYY6219/Ru3pIe1HyAD8beyErpwlCuBOz
lNPBCzWkpUhnZPlcL/ytD5a5urOY6DADX7Pj4XpkjMSJM+TGZtoPc++cfV486vVFOk92/yZa1NMG
CrfYEnLQvtzWHlK/5VpnbfcOBGR0mE1vp6M9Y2CuEUVnYwipbjJD3AuJZj3GMal7OD4B94RZ2dAG
awdEVWNh1DtvVLpIZr4rpNMxMGS5K4/DfMzt1dxUlbkLs34yARl7XEfrdSn/97t7IzNz8M06gQVm
Ae90jFAJCvG9D/PSS6HOYsEYs3gvRkiw/iD7xeqQpsSono3sj4WC7NRlnR8K9LaAinRR38CHjckU
KXA85+tLoerxkmsarW82bfp7Aub6hfC88fxK4GavhO2via0jOuYhzgKBZhU8Oyw2PfhLIVkh0o8l
uvanUXlPhhFap7RPglwwlMh5N8PjBVyNX+J04klu+wyWwPT/fcozyW+nNMaZQbkwFgmXL7BWR438
tZydhyR5p4mW4h6lcCm5WEKEzu94XNkVHHE6Xu1XlIOUwkDoVup3y4kWGl1Vlf5DSjo5mp8GpTBf
2/TZ19KHmhETj7JvMfwOEPKk+0mozBlSsTqsYSc98jXuZoJmXFt0HEEOPQ7Eb+eeRueyckUnoyqV
4P4pd3pVJZ6839tmvA6O2a2CHg5oXNFXowsQMjY/tJmpoltCg/itUW28KimZJEdha8SEIpQ9ipzB
0Im0cOAiFzSXBJl5e5a3l2SjjUFaKo2+j8+l243A8G1JEmimS+wOM/bFI1sGdMJPflE6OjLBBKHC
7apZTaSWkr/gWDEqsTck020sW1NL+myYfktHIXGeAYHn0vtzPXMsNO/N99qFYYiZJyNpMwJNyAPV
EoTTUkwxV5CNkHXd82LouH8Xmfn7PJ7GPuir1EWGLeI1PigqCl/1PqOvFNAkbKeL47lsS5mvxLv6
HxtzNv1Hu+NRkzIuNP8E55KCajc+Z7nXoaFeyTa6LfqapYfZcYKnoIj9ZmkZWQqNSnoj7zGasNU5
Ur8uW2EbcRX9gyt7akMtUSXrmng+rLBsVyUBd5N2bRiZzM2i2F2I9hPAeRMb0B0wJ07or47gez0J
qHchL3TLOgSva4MULQEPYAgS9C7XIC4suHFwcIx8viD2GbUmsYVHEYO5iI9vPB/Guhamsav/oW6g
OgYBb62Q97rO/CpLKAp4xkjThtEc2+WJK8yB5sj39ixxumCE+s6XlAd8B4VODZ9qBvHhEDS8nBI/
iWZq4yTKiXBogBNX+zZjLc0z8PMRlxGoxpIIcfdC+5p6IGneaL22Lt5KssJr6je5SHROrkb7AVJe
UGijKOvXulaoFsc8YBXytipTJuLvGQhCyqyhRCEa93eteX76Z/AuniMrKithO73CZGrSUTjdDzAy
CXr8++feqxXa0iMdBb/VfpR6wHBMVGlne7DWbmRUvNgfEIRNs2hEtFE/ZipPwf8Erotus9uWKo15
+pYs6nk+Zzj28CPg8wZzvn3cANqLqLwqw6Ju0saedS4rPLoZcxT8x4cGy+PL3ObstRaWsztQkrhN
7cu7jlTzbNTaQwEIL+WCXlwFIvHpz9yg/qNScXaIUlnV6YrN0XvK5V3SmQLd74mjwQyQNjboV1D0
k/RG53Sudpaq1Ic9EQbwCCQtPreAx1NYB4ylD+II1RBWVQl5HV3pH/AjBO1WMW2IGpIFVNwzw+Wk
4709l7fIKDbx7PwTZg7aNDJFmVq7b/Wjs9YfaIB62xCkdREbV4Zj5X0pqn3LezDz+jlxOBG8Yp15
WgxQNZd40Q209n3KQfJjYmjaetOSHYQmz1aKSsCzKfJMvT/Z1M2+wgBKAlL2s8QnatDMdS/6O1S9
7ooNDXan96QgVIn3ridFoOz9FtqC/IT8KWbVTA9uzOdl7uMNWfRihyU5hMt2eHw5CyHlJ4J2JROS
8ESYnyl7atyOMOVaJpAPXwGXPuCJLj6lWXV1k8mG/P6B4xCP+dyAihIswv2TACOHOODIQ8yKzeK+
iqFaYAshPkT7FszGMNyxDlQH4B1nw6DHcKGoHPrxjAD9UqngURUQ/g2eXCvFAiIB8o/tywfbTt9p
OByTBlv/6Bt8oRErrQEH68CsVCLbdwShDcZC3QSWYMDCbdoOt/tMMavuxdAqeESn7CUi6I+gpH0o
B0eKo0SPsRSXfX9l9DPANxLpKx33K2YtXLY9f5W0veg+/SgTcRmjtCM/QTZwpaov+aDbrzm7nsB1
Sg2BTd+OJtcAf2J2IU52nkeTHh54yJ0yQTdl+/3wS5AcFgRQCrvJcD2bj7++gtSNazXrovxmHrzQ
OQWVAWzHFb5+T4m0nu55chNEqGw28STy1sMS5SNqhHUt9o3MUkKp826xA6JiEPO5sr+0A9ymbdhY
UtAksbvXOeFYomL1Ihbl9WHReG0AtzI23OdZTztBPzT15It2aDyIwAurpf40IkLoF+ad2z8WRPZt
ux37ZeOTDLEXuKLZPLvnAtxfwhAmj0grcPaD6qdkhN6dpXIPORZ002KK/wRyvgYqlowSAQniaUHH
4F1L2DyfUFyY3CH804WSv2+pUaUkSPSv2s96Wc8Cx5BDPVj2nFHa1dHMAcsBrzctybIzUIypTeFD
ppmsZWu5SjjhOPa+uRbMV2usasOjY4Ftg8zQ66+hH9SpF4AqTBi0FZHEYoxb8ne9/Gcee3za45ua
o+A2b/h6OISdz6USosoD5dHbT+ORAJtBmkWQk25KTW4ld4knd1xjDevo0JGAHhdcQnR2vXFygB/s
FGtFy4PiI/3pAJLUjKgfovEkoI9x4mEF8upJqyxDFqv3Bg3KY7pkmtlDeBW4iQFNFakdVGuEJPG/
sZu5c2UhVJpBeBTW31/WLrPqS8xXxcI2VJ4UvCSAgBCtgg/78MmqbxPpC2tnsv8fHk8hDuvE8Pyr
nG8mOstyVqJPPCS20LPw20DWhSaYA5pGaItwApD+4R7gUn9U8F2kEy/UXVeu/TMJMHdhs2KvWppS
3cGQxNfPXSFbuJpBGL5TbFrkxiFEIMNrdT0cSjMlc2lSq7hnJwncG+ION7izQuHzSAM7EPU96XTx
HhD4d8pySFt87WRw73AhJArRWSoCYhM+vUu2bBjKfzr3hhCW1SDBnpHEtIse/vTGAWJoAXD0iAH3
pc5WBM4GOszb1KvMAdNxBV7L67Hx27vdfB01fQpe4xzLExY0+lQcLzacJurDcLWpdVlfifL/fbSw
PBy2NchqDTttl23peb/p0tBsNcSFJoC66ibhccf8elrIOgHjBs/dPZRFa8Cye8GStigXV/F1W2Td
zeQBHM89zlO2c/sQTPoYgqwb6OvpbEzxsaOdtatWLlVXmNA3uzdkpXPk9EIJFsmoR+YlhgJhCBXR
r/moFxotyy9+w1wkeFBiIDEJUAmIpdLDD0jq2wSIqp3bKV1uT3BnOMLlaezYNFAIlfB5ESWSKRbu
znL6263QhdbeOvKqxq9nvMvpMyxUgWdhLJlkneDiRIpGglY+4RvkkpjDPIYtAPRl36rRTIzvS2i5
I+NEN/KW8WMobzSNKY/kL/HCwuvArAe4VjG5xrDwle1kV8+7uIVQyy8IaxQVe8DOoa+utVxh8xQh
FRg0GBug+IwgDBfuFqRhIWyVXr5oRnPVzwGQPTgbHlXpQC1qaJIO1yDkEFQaEBFsql5yv/qCrXAq
9+IMYU+iYmdbCRa8Df1cUqUhct++sQYrqXnD/NvB3w51D8z/2hO1HrD5KWS6uNG5iaY4Qsf4+mUt
pxmgsx2Y1Kw2ZWvchW1VgVHrb7NS0oi9zAA8kQymJXSd4IL8mFEm892rhXJdFHEA9tkEI1mzy9ak
IUB6yfqTNEtTXsETw0fYKD7WsqdduwK4v9mdlqLVsHKhk9FY00CuzY8OeRMYZK73dtKNwNM8vuYi
NVYSEpbDcdxnubjP8abu1lxTG54tNR9a+UxHemtHifCJxvrJNKfC7qIgKxnxESlMRU/R/C6npgw7
v4HfDADVn3Il0F+uBsJufio3DJNszRlJQVblwRwfUM7USJJHhXjsOJKvHX6ZXDMdBh1RwVenSUDk
BJGPvyrjMMVEBR/n3+TtkqNgZy58rSi56QZmJY8QELGzjLsaK+P4N+0VRAz+kMVeq3pGNucrQjQo
++o1+/q/ZoaChgB17RspiqoBRHiKJGDqLiNbD8rFcds12rsvk4AkBjkCBSvtnSJNR+WtOoD9Bbor
wED+Fgs1pwbmesTgCtZ1zMISHR05j3njyKuC8toR5y1IkZ/fDiGhfA8VxpN9zIZpz7jfkY3z/HwX
PNOL+yw/BOGEj1Aj034ZI1DYVeKNsgjG32fBEoYUsz7jKccGcd9Sb7VLCs77y0xu9doToFnETbHl
9Rw6ivVLJRGZ0vKG0jtN8k4UxK84YPnZE8xcbJcByZmCtrHCFpnkf7lTmVfmQPSiO3KS19xavOq2
Xj1C3iS0a/CZC/JpKuAqzqrHrjgzuY7O8MKG7Gmg8qYiFhAJoUJdZhNWtjJ+ghrk1HEdECl/8S1l
TLvuBrDhU1HQ4LbyX/ZPUq6qyLrQy4cVtIeTSVs/lOYLZZQ7zyz12+AMuPy9nA/VnKkOMfWolSC0
4cXPHsNi747cAWKZ0hbzVZSp7CTG/JooW3296jCyV82PORZUZP1eH+j9Mr8bVNPfyxCZX8MKIzKR
qm+M5TXuARPgihZB2+NppPZcZO/KkbiBeYaQJEtF/HegsjOVXhOnYc0Lh/eNgOYcVqAvh+ip+Mwk
os6kUQ3UhqUsERVdrCcFte0Wd+nr2m6LQTUzbw1b8etASm50Ckb70i6iE6qDcivozyuo3W9xiClY
MOh0b3Fl3qBQ4WI15fH/H923SILYQD5bZO5Eg/0f0P1eOHjtK5IYOB2lQWnnVQUMZZ1Hh6IT1ge/
2UNFOHLIlTwcM1GMj4+WuAHEcc230t4ELkZ6E+CYxnvX5uceXTyt/13o6gutXw1BiU6r/hiOXwlq
eOhPv6bPVBG42TalWPudChyO1deSMtilyCdyN4kGr/rxejRz8j6PtX1qJ7NL+Vyi2GD3H1ebWfZk
1eeyH2xMFVIuLudRSsdCP/282fjNjqbEK7fJaQFzvrvij6fQ66Dk8fFpHh2I9hf28nCf2AlU6Z+c
7EudjwYxd64mU/D7Tars6/X1yGA9m7XqLYRif60tql/9s90efcar1vHPHB4GaJDUMFLns6MQ54e5
cCiCA1aDbYCW24HRixevm+Bc/xN7bXDUkn7jo6/i6dBz8J0I5nG8/IXGVcYJgvVFAkrcKvU7VhaW
quWxxDvV1DAWf/8ULYCrkxbOJN3HjSxdo/7iLuFHVGpZB1J6Nvnso2Z7DZQpL0tw7bhTLqtuQdJU
lwoin8AP6sxmOEHp+wbBe9W2fiWpP6JNzOPrR+MXSb6Ps8hrW+SXf6Z5qQBQ24PAV7psBt5XUun4
VSnFF1H5CTxg+Yzbo1MBWG0kQWRC359/Hjux/NwW0fz4ATk67BZq3ION1Z8z8hevOniGPNgrzOrJ
am4MDLFm0xxZhoC4qTtXla/it4u1ORNJgNtqEbkwyohaPH7STYEPia0OV1BLMfCIYltstKrxMNFp
wS2x8hfPSiVmzNwrE3KTHHG7J11CHmVi6t2QCRdOakN6Ug88PjzmD7CdAgpUJBhinzxKkKouPSoq
XcwcWJ03ET+31XgoYZ7EKj5IxKDF+ozj8rzkPfU39uTRT/m5ccgzYotd2d4LV4/efOj3wM2tze1b
INPBHfjMCMmCM3VcIncLU9yXpqaRQwtPw7u22O4CgPX3IGVbIrl2/Rqviqel68/nVQYOn8bsHqT9
l4r3qORihx9RHU4SlZAxqDxW9bCSsiM4EoHZaEMmJqrLndkCBAAz1U4KMnr5f0ITiketl2hQhoWm
z+/lDhN7xoFZ1uLX6szwcQ9Wx0XXpyhv5X0pZk2cInHoTRg7xaU7P+S5uIX43QxFNu8/ZUzTadou
1XoD+NRTMiXl8JFqhgt/ZZi/vPhPhVIYayTix5GnYYvxFifzn2//Dd3kNGofKOoddJbTRTg3MB2h
2h1HXKq77dXQ5/wq6Qmfn3TY9SYajUMS9o0aM3TwA0IHJBCec3zGYjYgxh31VT4Ogh+E6c3i8bAM
O7o/Dg0cMUOTFetQUZhZwLnR/iE1pXa645mphSIIWNu7dpEMfEZkUq7pHCkb3KniFlUKkJE0OS86
sZqo7+smhJDt4Oh5cf+xI9YN2za+mW7dj0hLZC5ilSoDSULzxfOS7eIGx2WXTd25OiZwJq7dX98+
cqzmUsLpvr4KD9SW6VgyTJJaSlo8O8fQrY7OQXy8JZAES4F1ZUHJ7DtLSkvRhXbBPER5PjVZhjhn
HRDoGx5dRCTCZE1WvjoPQa0FPFxziVgr1a5Xb/+2UlCYQ9H8btTHHHltf5s0hZv35Na7Bm5qG66J
Jh0F/XEMzb87Re/U7wYMZKfmhS6j9sQhbS7oDwXX4nzgW7QeFlF8a8Y4+HjkDnj+KlzUqyjUeB/h
DUfpd4Yu+ucloA20XbDZnYo+dZj+G42reLY7yqlItcap+IKgF8WVOZtFsJHxGL720o/DxP8r9pRb
F85NnR1+UuqYP2GqkGwqMltP2gM0u75yHCOel6oaRDhhKxSxuCcdaXlve893YceA4Uxmi3+46kDS
qVepMk3KNAuN7JNwyRWhiYZmdX1+r9SOQpfULhR3NhZDvhIBL82KvnCq9Q546PMsYT5dcch7zXWB
8VTtTmL8JUWnuc8ARkKBenVwVXtd2yurMr1JxUjYGY+IlzhmcJgauMGqs8lTWZHw2ckiqFC3+AZa
HIKxOBw+M3XIbG0VYrPDSSVKnmzyBpKjlIdwxOQn1um0K/tXxMr0f/nXLTMWq9S/bsknO6E4ik3b
+Bq1iAeRP0a/ExDuwO+sTqeW6gVoPm/Fgb+VVTNGNRlhCC+rq1WaMQL5ds7mOCZGRq5tnCFnR9SH
kJA7NReoE3G1J8g4LwqozIIVzJNqCVmsMBjdojp23K/k3IbZwsmFD7CEPT2HY+yrovtS2P0bueS0
KVF9DYj2DTpI3RmTvRBiOKrQyZEbde+IWwzLr8mqdEv4kEzLz3TVLe9peRkxKijH19fACkQEeGxO
DLzNIfMG77tcZ6U2tBGkZsiMxAAwW3SMwORlNP4djoC0siUC4yVqArbW41uO4/uXBy8fFxxjGZNy
l0YglcOxVeOngXtcBHpQW5PDPFXjgmzUUV54jT09jhEXC5iwyBKCoUa/Ix90lfMiYXtHIXNl4v0e
oaOedWDM1XwShDxloyXGHeEQrBvrr08tVfTwjp6lNCjgz0TQOpsjJFFCptpIVhyqA0GSDZACGWBn
xQDhzWGb7LVVRzP1xMvKMnB7Kx2Hn37dMqSsO9ARu2dEz0Wke+z/+QB04TnKT+71xqQqO1XLKU+d
uj49iwtD4HuJSXGyWinre3R3fBoMZVXwAeR8L/T5vJy+rKgJwZJAc7hRTt4WxWrT8dqEOrYk3WAf
VWO1k4nUjpwuj+KqUEKwPStdfIS1d0jva07kEUH3C7qOfzYSBJvepQ5kFH9ZF7FbkyMKG9Gp28XY
N62POtlY1NlWRqLoBwJg3Y8l7tZkQGf20bmaP+QV/qpt2ZGh7uh5e8azni62WFy8F7zQL+8Ona6P
oVIKg2qqVod0LiQk2hTWpZv/poskbSs9rKLOyhvMarV6k1OkbPRgn9RWwVemz0EBWYIkyPBs9OcI
ulxqooV7zU4rmivKow203BOOm8ZKqqBpeAnztrTSrlSnqBNR6vXd+wiukh6uf0qUqljYW+Fifl3v
jYu98g8zU2uflJZDUeRDs5uTwGk4Hhoap2RNrR++pf4FDMgDZeppcj6ZaL1iwB0Amtt4vh7fW8Wo
R5plJdopoTds1seypli8QokQ74vjuEyqd6TDf5ZGl6H3gvrXnwoSbhaEDBDdJdczZ1uZHQyAMhxP
W1+Kj5Jdy97hprb0jI4YHur7fHLB8Pez10aPAhdmHdHnYdKGNr9oc7kBWx3n7RHUL0soKscr8WiG
kIsgQAkPsTacjaMWQ3IhqeJLi6pCVMnmLr15MVhWMAofx7WT0R64gsXPyQaCFe9+ksTc3iRH+/Ur
tVYNEzQC26n1fLVgPiUYCepNMFdcU3Q53u2yYCHYM+jwj2v1gt50Kxc8ei8jPJKRj1CNOsUIdujH
ZP6FQpikZg5ucJ7HEJg26GIlW/R1ui31OmXZYxhRkwv3Gbm28Ub81CaBQ2ftfFNoIp8GYZWG2K9s
nBxYTX47BXxLMQTApuwiPWtqglJZNJXXDFbL80Dxvq5yy2uCgmrNkgmEUpDKaCRYO1yF3dYEFnyW
Da8umeF+zoWdvMGloPDuxiACo9NFdj12B5okXZp0QbZgC2YMrnFmJIcbMy/yOMxfGLZ9pPDxwCsJ
aSQXGIgufPd3Vn0rdhZUW96O4A04n9u66tYFYL4ARLGBo4utbKckTntOYMPwOaTs6JuskkiOf8YM
P6TJW9V7tRAKQ7l1/V1DVXAGftQVtLbdVbTycBCIPLfe9LqeGi7MxbFW2ofQEGa2D6yEvzoy2th3
P9SqF/cHQXSc2/xei2M1zB+Xx+v9Rq1WoQiKu6aCdPiIA6o3kYh78LqlcIn2fZf4Wht3RmQcsMG4
6MkX/cJs8BJSOSGWRzj+1suB8sZ+m8qnc/Y1dDkkPaSIOEY9/Mu5j6j1g2kmFMzTUOyO7Lgd23Wb
S0adKNeqaZzR8F7XkYL+O7rvbGhmuxUXEaP2id1/v8bugImz/oCqvdTACGoSj+owsm+g5xC9lKO3
8Tu94oPRzr+87q1Ps8Ic/c74o8j3F6IG4nn+Sd98LUtdEEyOdA/oe2H6W+4y7aYcEylphiJmSZhf
OwfVWngEYNsyRGGWYa3I1qhIBD+SGHXoetl+ykqgqpVzd3RHWGOaAMUNxSeXrYbEShsNN6dnw91M
vXsYqOIWefA0wOSvodLGUZz5UAIaD8qc5U5eoK3Q6mPVSA2GuxJIe243lhFzwkiWPMhojMxA8oyJ
7aMTZJMbeVJ3yvdACSYlzAA1/nrLxwFcStPyvqTISZCvXe/T3NtU4jbBc+Od2adCxKF6lKSOPuln
xdqhMI4931GyYpo1bjp+NqJxODsIs0Tp5fWrq+zh3EMLbfq9i0xrlnoITpDvl2kpeWqp4BDxX5L7
ewQMdoBMvJeidfAdE6RNZASCFJ/4QEi7+5gNIlbqssm2CQH3j+vQtBZtv/M/3TSGb/GL+szDCK5Q
asiv1HEtlOgtwCFlMU8x7MxGUzw2+XM0scSCyzIcIMzfZfZA971reRJM5Y1YtOfj7wlcfORZq7cZ
8uIjFww1D2i4/j2gjdov4cmMQzIycWAZHxo6uZf1LrOzN8jipuPIjgmBWs3s0Wht1dwywc4CiveY
vVSqkeTfydrncQd95077crXPqhBl9UEVs9WIYkCwHRKEzEt+CBXyDjr4lF4pnBws/FBwOzkhQTou
Qlg1CTabfKknDcPz77+SaPbsiyaJHRWKF/BzPZ18GRm0cS1+jJ/mHYuMsRIV8F01A6uDnuyzACsh
HO6v4HM69x78P12x+dwV4Kt21Y+97pvGAvLW2k7BkJyvvmqOvI9TQ5BWoaw78frArRwFiazqn2mm
pz5ZHuwnIlsqAxvVpX0L2YHp3KK3jqzT4DQ9ctQQET5VcULd8PWVrN51HH3Y4RL/IdjK3DLeMfPA
L7ZzU5Uhn1qd1TUJuNMR8Mz0I8UBHS78G4KcRKxOeiS0aYg/vcyX+JSfAonSt5HLOvhfMPU3GHvG
QGs2BlzP5Bg7rtMkm2a+E0I6+Yr76ov2DsXvlJemcjNjVXRd+YVeZyr5ePSPZnqLnNSz4xDbGFOA
llBBlVffYv7Jl5uAoaG6PO61ICUM0vNQnVj8N3/iAeJpXUQhnxCDzNQt5+1fk4cEgFREaiaVRi8w
BjO6KV9d/Y6gZFRN1Oqy7tLmzneCWngInrasR855ouL30kTg6KGLt21omf/E7eZY9VpCkYsBKW5x
PGosThOkaZKUhtMpR3PP6zSxUtbdekCPXNMBtmXym2z3StDTmi7DrdxgJ2RmTuE6/C4A50uWNzwm
LIgg8mZ3FSh89KuYqUR3gKqyHBCkCkntdOQfzxRHDWDY3wZF6xD8yKDPEh9rp3Ybx2fC7XJF+Vyz
EUMIMmrUxGpUrwBJ+MHhQn8pOAXBizpuVoS9xkfQfxLhWj9W1A1T4Orh0iN5Jkd05GHgxrXEbZ+q
Ia0XNW6BZkUakj95Z4ieyJs43YePckUXMKjUkD7qtuUa4thdei8mLdzgs3B6CGAtBoYUGFp4xjn+
SiDH4kOvtSqRbb4NszEQ9ByaMuequF8+5xSPHW74pLYUD07l2XH0Ru9MjG6NxG2I4okqPajLLigl
N8yUwkndJHE2w1BXgD3FZrlyvLJ86PPTEls9eD+wEiuQPA+b7zSTOYUV551EOE1h5qbdby2ny1A5
lCU6sNvWH1B2yng8rGC+Is7zGYh29Wmolo29eLmcbcHGmB+YqWrKIPzd8k6l4QaImazDId+7Hljc
H1Wnip/uFlrZxwh7Et/f23hQLZLyazATs7kxxRf5299MkOLd3a8rQdk5Sr+FMPxLbUIxz7YInu5H
VCYMWAdI/rBsIAuB8FB4kaS2pHNPm58yvb46UA1eexflFwnYegUdGcXo5z+IxN46Mu9L3drOBOMO
8LNZ9eyx4ESu8NBSsVXjjXM9+Ood65l1+fH/1oiLwp3Jbr/uvcgLnQHoE/0WECEVbfl5bbLJ4/J+
BGECpnJBtUMy6iz1YugyH/Mu7nYYZAQMsv2Srig6B0jtkW200iGUcq15axsNAxb0IulfOiOnOwZp
QxdFlJHiJ//cbvEtRUInTTUenPube9lBscobdUNZ/wy8l00UDyC21prKwnIZrEjs13lcNKKBwohz
GEaR4gm1takwS4o8F5r9MIP8pOwScxRfPXCuG24LJrcSFRmhH8CETmGI2AiPrkNZEqxwJ2CfJn9w
o8rKI3N8UxqPQz0XVoJcJcK6JdWDOtjX6pRFxkzNnvhLlnJ2bbHy0wYc0eWl11O/8orv6HVslIbQ
iktr7/zP9Rjn+KEA7vncouDIgLkEq0b1sxLRqRkTh/tX1sb2KhY1FEnZlkADok2AYqR+Q4MpX3NT
kk195W5C90hS0iRnTUaRwq/ehZIs48sFH+CyMPV5n2ae5JPPSX+2weKlCgQKw093oHAfpNB13pN0
99WhG5yyqkYO5xxaB/e6YcGufIVyeRPLzTwsHsM4Ri06Dvn7RKKKVicSblBFoN9busjMpUAEkUnh
AaEkVSu3dBKVnk2kzCpcD9UOhpf8OXknw/DDTuMEXpBawj0LfOm3nK0O9I62e9GKOM661iUbsHY4
FXHQwW4VLLfAVm7OlY/Vj4MFMWueO4y20HhPO9Z1uVeTJDewdKKmiiQczY+d7h8EpjHQ82EfL9Dl
P6TCO9yrOQ3t/XJV8oIlzdi8po46C7JnwwJ2RRxs+wm9VYMCt1b+bVLh4rI8D01L6ujDQ0coZhtN
WaNGvXrwNeYx6/m+Ms+WXP59KhSCBZek/klEFDTyvi5rpS3XWg0Y+Quc0UsHJB9QTX2yZiKoqXWl
eCliYg8h+a5uk/0lwdh3xREPD74jUC5kWT7Xk1IWQ9zCAUdWCA52UOrga+1gLebpVjRAUVaeVcUf
UJqREpt7TZQsZx0/gt3cWcy0ZOJQZPqgcKlFFEXy8sbUaOQ35+IcLb5aPj2IR/GAKo0wwA4i0ehc
zOKsqYCtKic5HVrSsx2kBJcUUD6lGRZbmk1Jmlnta5IojF6NDFPRvLCivzqwQmEprGBSkC8A+aJz
m94CFE1b5Yo0nMifMjml9VsxUtR1iczD6QsaaFghX3F30sJIHIuasmPr4J/XecIemDvP0t3zE7LB
nDDlACSEwZx0mgh2VGSGndQgjAIMc50Y89I3WMv8B/wrnswtwetjaeiZ1WwvqsCmUUxaGHxAL5LC
0oeswCTMIDU8kPJ6oHNJvCKt4QIw7XIIKFl9ql5gccgD1yLmbJXSsq32QHMzL2NW93z9lxkuGJf3
rnpqxcsop1hW1J/o2RwoA1bOkThPQMsUSXT7D5C0cJd2CwPvnbcRwHROgg7NvNPbjt7q7v4tpxqg
tCm8odpRPFG/6I6MIBJ4dm9lykYw3HPV2NFRnamO2pRCSfbSmYQtD1FwzQ7XRSQ9U8uwDHgtyqyP
2OV0PFqcGDYZQ0eMcHq6mmdx9zg/6LMA71C5KQ1mrDOhzK/JyE7t/wiwrDyhquLz128pNrH1WIVt
ILxeeIZ0SbB+CcTpVgcfxgLq1jcaowPHD+dgvrL9z5LakoOr0DHIhHqCYwr43SNDWdz+XWjtZh8l
wI3k96SnuFMeSbjuklXSiR8bF0D+zuoS90CFkeQVMASywE+bGNZGkvbvfbFYEZ0IHvt+TFxhqjZQ
enyNXZ5DJMszCG8dmU3aB7O+AoQCIOw+g7oQdOB6iLE+0//6zT7Ga0O0uR396xZO84Xc3qwOaiQ2
HCshF214fHjh4CKEhBmt3ApHVIT4CLXsX3+yRdoIuFjGZh8VNzvj/f6BXGhlopyXOXntCs2rTBjY
M7PRh5hVBDBtPGir40XQF6jiNqLhj4CkWdv/K5h383QVpdeSGUTk8jkmjC+IgcVou4BrcmV6/0ik
B3K22umqcvBCxiwbYZFQmKsR5iPr/hmUzqr6xqc6X5sOnYGFyiYBkRoWc8Ku4kmj/+jQ40d4u6st
R02hIrjwibvHtJta8ifiJ349jPON3y8/4HwC3Jbk507WPoQS7brdU+xF3LmQhGbTVWstvgxa9HhV
+yBUF7oWP51uJoBqSWQTiEGw+hWwoRGlm541sbkzUf4B2Atb6/5QD4cly3b1cJ+6AoBiCYhTGskT
QHwhRnzJFTmj6lfwL4zbgiIbTCRMIvyOYk0wTJVMsoxkJ+6/p+o8DhMrsdWwEvVXhmHstOb9e/mP
WknyRXtyL+6ZjmEnTSL1VjYIrhwLSZrzdJPooBT3d6ZrxnX6nWFKW06M76s5I4aF+fV3lrFjRntO
bFiqetRY/L74GAo3PDrsI6keL/Mo5ml9O+8ch2bwO6YF4CAWB5pqsrjRcz01XfvJWQ+2x52shHJv
T8Rr9yD1ae9AB5xaySqOsJfQokKWM9cx4xjyYlU+EyeXEJCfKQKtuXCWPXWN7+fcnTdBEy71dQrC
LaNyY0BZrmbh62a6WNbAtXxNRctfoeNIfUBy0EcV4eXV1XG8MhXAuixSVq6RoCUi6PA7m2JxbKsk
nzY2TzrKNGAALuF7eFDsVVRQhGWa9tBClO/Jo6lEPZPSN6We/6gCPoNuwqyeVFSRA0DjvTAgaKST
si6p2KrfobzjOzgWZCRkekH7epMQNarwYrYqOOI4zzljfJcfLkRd5fjpVGMB94gr7R1nHlXUMaRk
WAIVs5J4zKQHPIMO3yU3J+HyJYzd4ZOGZFoM0v/BuMbrAXTlPzx4t6F7E/NJSnJTkS4n/EfGUbON
DXtdmzlMKasOJ4uYkS4r8lm1K0YdONux6UWUrq2k0B1brhELPvPp1qk8qmekeO0+hcuZEptEqJNf
u6QiJ6BeL/mdbAubJqmIgDfCWQ0+3w6iWZH2iQVjlNKfEkv7R2INw9+HTOdz+JAIiL1fhV3JZSv9
5LiJd6F16McvYRkH13/zY7IpoFqs4tRE6sxHf+Ef+Aqv14T57JnHvfpeu9laHd0AmB4G9k5TQKD/
jjCXoNkztD9kmXte1rPYx7HGUUb4O/9z7tdJiuukvAjxnjZVN7V4NY8Z7aSWyO64HLn51SumjrB3
69Zdwzzy5TxdhYutziKexAiX3nI2p/qQkOf8pskjSH13WrtboS6CRiteZZqgdBwCLlzLR8TjLpBr
KIwZm9pRo0FfZJTD00XrVGrnRYiF9pRTcsrUSttrqGCwI1rTGrFMKzFETEwxorS1DO94XGwBosg1
QhtpnYjfEmYFLjlHcAYpiTcqcHYlbhltwGRJ9dlIdAsbzOo64m9/KiSBoqlr0S5zqjieycTMVdHz
LQmHCIoto/rwq7ivDY9eOxfYBGJqHI2qQjWWbvEBCYkYkyWt3Sft2kQvJRAdO7bSbvYnnpS2+a8O
cNGhdylc0MKLrPwBM4qs91F6/hpuQpFCpvM6AAvRPK54H3LUn9Oo9A9mHMK0Fmmzw+DtpoEZqGHm
8hEXsHA5MYvSZDWr7OCjiZ+2sgX6qxpOTPd+wdHt4OA2LLgRev/LiAtgSTD/vfM6g0R1TyYxCVPq
6uyXC8QIkX7hHuh5WnfRip/7cS/pwPymDhDP9rBqqNyUnNDA4o149Rxm0fb4Jf6JL6xqCLsaTCcX
r7v/rQALaid8CC+LbqEWlrUin0XhPWNPiCT6q/887oWZHeIobHtFV7Xc9ovEEBqCLw2fA/RFxXa2
ozOkgJJoTxtEavCv8r2X2Yk9xMDXklAMHhnVIAUAY1uAvRUSDXeZaJG9w5q3zFdtFMMxYi7evbP0
V3xtjRoMBaz6fN+UrKv/AipQsD5dgUVncFgQjNOfy3gea2QZ3QFsuKwtrh644bUMn08AFCHz8EZ7
iQm2JAVLfHmjLh+dnVKCB4dF6UFhVuyXNrAaIUZ+rSmfg3kNuc+Zqc2CjcZkn/0JO66kdfIui2Bc
KjUCkmiJTXD0U2Bx/PdijqRCyq1PaWHRUvP6c5FCuN4IXWwLjZVJM2EnByMeydh3xcYuddRPzEWb
O/SchE49b2n1HYLljDKJA3EP/8YJ51BLxbGrj5QXEF4WbRc30aat3dCj9UxomYoqw20u43+XKawz
ATsyG/osQQw1N1dYptNDiijQOk6cLeCv5XkHirepmlhfrdoKhiaE1v1sFArBLmD1SWsItHPCjUd3
9NMUddRrrulVfmLQTTT1PtPVwzeabgxAmhZDQo49rHHbsv02FJ0JaJjIqm8KLZAj3ycur/VjPvTA
wVoJ0mUjAeZP+1ds4VSfs1aCNOX9t/CsFQ9ASxuMhMeNRhyU22cl3O/vSrhx5Ph1JY2CT/qyvBQ4
63ZtQWGQf99ka23BWjSTjIsS3ROH7owU/WclLnAX9Mf0lv/0F+S+cWRw3P0SvVaC/NSLe5ZfuIxE
0zjM1DmPm0LoARLp+U2nVkguwp0hdwbVj0rZD4+iHcq0VYo8C3xsbUhHxxJ32VIZLcR2EBfufdt5
q9hCPuET9BA1FwiOwpECvn4n0lLnsHIloU9r+jSPAwLCQ4EhLj/EjT9NVQuTJpAbuFJJxSqZKYhj
3KVydQ2FFZXGqt6JaLrg9xpx8ygKTQq46nZjVLb3KATV8AhAxr6YPiKVlU9ow/mJi/HOEE8ZxmJi
+MG3fFwGXrR9vM8M/S1vo1NWHdtGoHay+092UlyZ5KNwknIW3H56CLlerccFKfS4FxDJrciwe2kb
1iA/V30bomaztDNMH4n/9IhBjAhC73NvTmro7cgRE61Vwzq3H6XuS4ieiEVFmd3gGjwoBcrPCprw
gU4edLz/xxg2We6OHdP2INGLAKKe0i1za6zhNHDgIhzrzje5pkHWopX8e/Nxl1acW7nE+tHe+iDT
3QTIp4mvKmf5tiFQX8GldWXCPSwlXo+bOWmfnchwwHFPMBS3varG0Jqu3+BfjfrDtx/cMiFcWn+T
qJ7q3mNPBm3uTt3wZIBOT49bdzpwbiRWjt2Wi3u1NhJtexSHQTRWL4p5aMDKhCLOfIpquCX/MLC7
625yki9BXp7HIGr4Ho9nOGlGxaQQT4ZqY7gJhUtS4zoXwj5WYd/BucUtRX9WriYX9X9xQ/mj9jhp
xOpspDGEiqfAnzuys+38hxgaipaC/QRmVuoiZ+GZ4lAKJ6COdOdcLDGkbdkct1aATBTXBYDhk+F0
2EttZdTQDZ1sb5OtecAk/s0rNb6qKq6NcsIn8f2M1YYEgrWAquNsZB/GSrOolo+lf4CKFjodFDy4
uXGZ+pAyrI6TTsHNs3+5Q4IW0nwok6HHOLzROLswXUtdXDxwVKhwfQoLddC3HpXMCCC0+rHsq93d
JMPgpoQqe2gTrxOqT3G2ywdDnPDd5qaT8Y0RJyXMJ+4PkKlTg0wzczC03qwowz933ZFPyjjrazHK
W5roGeSS9DAdJ67wUAnZL2eG9AK72vY7igHVkZ2VzGtpc9SgYJ1f7P67PblpdjD/4/OBkRJ9/z5J
I+jTxTMBJ4uy9deJT/636LJMdzZVppZL/W2uopSjePfFu0M3+Hb37ZXcDg5KFPaUatjkewDLPpL4
VSnegRa31o52kQKr4l7HIusUAdWWL0TpbHLwsUYTVRfj3vhtp3kPu8XStrX5xG5wivZxQg2Z1guy
94M2FEoi0EuBKsRWp2v8QLfSVWnmzJRcQJNePjTAG2e8pFMvgQi2Wq9POqYErwtFJvP7nfXueVd/
ZlS+1PAXYtrijgnWCzMLXmwzIY4LNLaMLvmIqLbgk1BZ0hmV4lS6/txoMZj6QEuuHj2QknSmuCeO
I0ci0tv/Fzn7KlxzWVgFA1+SmOLFPIXjse8vzNAwNd7Q/bgDXRfmYxrbRSeIjLDw/vem8txonbqV
BO2o8bv9tTVSAK9doBHAfKoG+RIUuN3Beg4oGxMTijGPU6tBT+y8CjWnJxK3pin6X1q30FVIGwi2
ZMpp1SObNlGvzL91gl2qg+gk/RRU4Zd067knLvU5aiwlV8cY/le11WwQvsHWwbPMitUAAqBBTrwX
tzYbnHQXIYPkQa1kDeRCWdlnu+bPACPCnDIJE5d2anWUlYdM6WmKhfkc5Nfuu/NQ/+qqGZb5rbTz
DLGp+ZXSe8lxrfCf4vEjCa45ZJYXlPhA++q69y2f+wUVmwYGLJPleox4jn6kjRPwUOsZk4rdNtui
UatDJEDtRFa65ZbIw+GS0muoYBxhXXbgAJbw+qIOM65ySlP+ANFYQGWbCisaHc7rVUYyVPNAN401
8N7y6oHDnsdxh0A8co5pAdLeieKaveUcVrCuz9KNotpQS8ACYgaxhq1/XJIivG8XyXpcqX7p8ZCG
2Q4Z6AT4EiNCW4oPH6jjPAPHoPw2mueDtNveYG4wmQTnYu55EiqOQG1hkPw2T/0oMZhxvYt58lfI
4GNe1fpEBwJFvsh8apvjcoe3vDIlYZtk7wQzKyvYpC2/yEAsHvqQvtNGfgEqe5k/GcKh0LJU1mqs
gFunTlyvy/ozJAKhaLTZO9uPKYzv/rbBmYA9ah78k3WuYilSkK7y0FYWfKOqFri2SkXbc5IT5ryc
+al8j1hbefbTUNQUksbSZWQiuE1ehqfHqkiLIJVoTnE7OI3wW/GtMqawIPwfm28wHaKK7p48Rmf1
WmnMkeJtLBu09lCPnfY+LOPbwl54Qc7dl19U4ir4iTXuXmM/aslbzlDYn99HVDHbSgQSdYEdpj3/
2eVkF1cUEFaOfolsISobXHYfx305lD2vBGKnl9DYMywCzn7mAGzYHpl2PGPpPvQFBPb8K6Zjo+Gb
XbphH5j5YAPWYP4eDFMBCoEcnOOliQ36qr8LLTNDGhOJSWvWiiF2Y6cF6KF7D48Pf+813sgSmx7o
ZiSvwLo4GOk2oFejtygWOiELSx5j92cD01VP51nb/h5bhw6ZCS+epAD5x54vBrquZ60n0LGxyPRc
qhD8+t3D/DNCtTLbEQmYMBf0f3e1BW/iOuSfMQeQvsxqTQXKD1vswFgFrzpnqtocGxiiDvfQYVkU
l9KFlmxUHEAtbUzsOnI8OyHEda2OgSDT4GBRRWrf+YimqP4RX5wB+7VelvFwwrFqlxtO4b0kGe78
TfT1MkPRO4Vf1Z5mYbuq+5WLztp0uweEUNRBTKDt4RnMu/UF9UGcJFFyt6tB/y9PoPXwDMa1xRqp
3mqqojqcsG+4ZajJ3535ciX89oi9ouxzv0+rBgE6vPsw26gMAKE22AZ+gscSzb0VFtku0THRthdN
raGcl2P0nRp05HBW4uOsc01is9rxxRCLw7dMMlh+x6TFC0zThYruIW6PwwxravReltSR5vpin0ih
HJAC3hDnc1qz3DO2EV5wClwJ5GTh8lHZ8PqdMQ8NHhnhVowgi0rThHvZxlIkLfxWyx0/mKreQbBa
/DAew6VyXY4qDNT/h4j54ZK4ToA6txX2z9zBumFS8OqXflY8WENmXBiz9qPfMXeLtESM62gNSXvZ
SH9HQLNhfSiufbQ30cLw8kxxBUzTg0JdCXam5fTqqzcQatJmddeouX3rz5PF/h0yVh9QZHtq92s7
AgYGGaGnMLnRS3a9yU5et5herWf10rOz9qyfmnx36biyrM54aI0YJwvTS4jWVh0R7JT+PBPouuJ+
PexycCvGMqUmP/HWDUwKVvqSput0ZWdqI/SZdCRWFU+xYwb2NCOaGv46Jaf2x8GeiJTOg5AvUNNZ
ROBOaICRMM4ut4jgRFnfS0coWQMYWC54FF4QokWTRSA8W2IpmF93JynChf2bTFaCqQfWbEyhmzuf
OEK5t4tYONsMu7/Wk3SBDuhrHrv31ijvOz+FSGhzyXJzbBCZxbWWMy91oJAqQE32n0pnYxVhfl1G
uj1S/tGYIQ27R0blpDompPYUGHqMEeY5gE0nrr5mse566wPCG8vb/h5yMqOxNZ5LI5vl3Ffsq7MP
KK0Kf7RnbFFdXotRf7zPSuSPBBW6zgW0cpvSCM7e4WLQT24RrcS5Go55jx0+GEagyKX3h1kj/dV1
z5iQbxSHc1mmYVxiJuMheu4z646EFXYcD2qIKVaXD1BKnmhRZuZVyldUbvMGtf4UyXxP8mwInPZi
+xQztwX6zpgBfVoTQfmgMNJbvaUvZKNSWcrJJFTCGxV/eqmDzMdvqNPbrHqUZBWdTHCySsaJoKEl
56k92hd90ni/KYcGooJsjoaW0RIMZ7Ar8rpOGLfqAMe+qpcWuGLH2nQZOhlnzJ6aodsjzdUV9Xvq
M7du1tiu7l6P3l6Pw/YwVzrhTtcVzPrHIhZhs6LozSFG1FEin7zFVfzIysvoe38LdcwyNiBtSnw/
/XLQOi/oO2p7uQTNyDcqBtJI6dYeWeuWUL6JZEFBG19/qeZA3iQtInTP8IBBWTMDvT1qtA4Jz3ov
z5mYAhZ+rj1mZuDuOAMMMv4ysdzJbNtLHa+uMDDBRHbByd8P6VnvMVyeWHdYLlG7i69aSeYt8Him
fCBbn41DywmDP3TPGwRMhJ00oBXiqzMOVfVEhEm612voNIJfkDmr34II6Yi0SRZw5nbtPg7vgXzu
cr/TSeWObbSJdgLQkFD0GzcgAXCelZ/peQCNpAG5ohoSoVInqNHKgknDCUPQI2MnHU0tkXeLA0Lg
PhdATjNZ8HKkxOfowMYRzqOnchRZq0U2IFg5D+tIrIexNv4XTGHRiSeev2kmtlCs6F4/VRz+LKTf
KN91C/wE0Of3i4P2CsBesuTR1+APnXXAzldJRYi7rd21aLqgvA/LF467fmIjwSs1gLOEFDLFY8KO
bFhpuJ8qVp0Qe+2TRlUauHsu1hsBUUDe+bRba8Z3N4kDCkvWLeAYHZWrIpMcUHGE6sQS/bx/FT+d
13fnzv4TbC3NUBVv8n4eENr5pb8ZkFRxxykN8FXgoaNRIoWRNvRQpEpxDBskrQn+MXBL9DKaxGGe
X6qEKPzTHGzMXuhlzvMeT8FfrHu+aysFQxeajmUDpYU9lDIqY3eWWT744fMdMXxtuXRXEuswyiHu
ulNmbjGbJ1e93E7viiNOgz9b0Xr/tN+NPBSL6tJFnmPr4/ieFTK4EI1Fu6YgTYDzPq2SatwbguYY
uo1GAzH15QfV3xkrCWXaYYOphhQkAu8N5gc/KMwdyUZZ8Tjd4pQez756UDwA8VdYpNTrQt1JXBkQ
PC0QbB5GeY9O1RqnV/UTbk+mT7TQNEVRYhBip7Z+tMwsLmSLtO72XKJ4ghIYi18r1OrDqE75TE91
J7/l3QpZs5/Cjkstvrdu76T5Xyb78nJ5avOYbYXvR/kImAxP/I6rHwiMMla33l/FIS9soqM++0Oh
epoGPEKyFMblreRZvkpqHBp9ZKtHgZ7kJrbLZKp1gPkZ7LA3mBSk0mRJxqT1aETGQT3DjacETpZM
4nD1VnMYVTQv+1opqnwOLmuY2abLBrnBqBK8/yF4rLaAiafCDamVyL9snBRech+Kt9g5cQjlXX6/
jIlcNATEESUQUKU2bDhEfqf/js+8YsoyaTmg6maqgYEm9amn+rJ3gcd9Ro+KzLUZLq+BVavUGQO+
T24Xdb9Sac/Ba9kcrrOnHHPuHK2iLa/mLYk/oB2H8tgtUqyjjcbbdOOvVEcyskuvtBUu249lL5fm
y6sy9H0Boijo+HPlWPyyEaHTbGGxsiViuIEr2i4KNbHWcFKT429B07lYm5tixDnUhoIS8D9+63ip
Zj5h4vMtC8WZAXIdf9n/3CIKuyU4bRr1Ve2pqwq077zthMO3/exjffefNLTdBFqAYI40pNO6dOfV
XXZbkUVad3fiwVmcVl3vYxmDgCL+3sP++n/Wn4KZfBq+ka0//a1TIB/tZXpIYvmwtab8f/yF6Of3
uOaBLBEU+2DU8c2RuaPzZ0vQgpg/JcEuzLObALIliZomtDl+yRkDLAydNr94Qr2VQG6pGTyVFdHE
sYKN5XCi3tk1yfIRZ6bnwlWPveVC1akUSPGBipesnA9V71w7T0VF2645x8Q+oMlh+UQmlW5vl9FG
ZfpfvnT1Kpe+adJntqcff5IX9NO85gCrUM1spRknCN46tBbUtyhbxq05GIo4G4RDPRyNJS3mgn/8
afyhus+GKF8sZx+7rPk4Fi4HYewlW44WscSPWiNrTRKA/LHLZtj9sn12H0qkHbhR+HMenLZ6Ktie
1qICLkOvYF1Lhkg61F6n6Ui+l7odhLfghbXWhXXtPiXwgKBXOaVR47kZk2Qbfa9RhfM7q27tU6z9
r9pAoR9Qrs8+gPqjoPn6AssV/PyVUqYihuhkXbZWUbeDhQ6LJwKvu9jhr1aaQcZGe1Uzf2R5voWm
cSTl9VzhrfImNwaZmlM7KU6weDEtcCQA+gGL9TZ+7U6+yR1cwyeiE9gnoSaLOdRupS6YzqzaIBcN
mVqoZ7mycdcrxuDySjKUcHxoRlPQozd5KgfYRvqpXYxlnjYZp0hdNjV4QPqnlgiuv4b0BWtZEgvi
cItFx5j1FpCss+4WkdZUidKoEkDclrFORulTv17T9Wz26ptuOC4mC4SPjzUhKS35NxpS9oi57kwe
tYkJivx2Rh1MKQyyUhJ2MriSn+jBFr4Gq38UUEPonqMp/MFB8Pmugq3vhcwOULBgVfirMqL3LMue
Ud4wpqHrnAWDeZBHAY5OYZmlTwCGWwS0umxNGKWsf62rdxyBAfOgCCGXp6orNlGjWUfOrn2Oubik
KgxmZiypnc3LvhZFKc4rWuDjMP7FiTR1OFbnYVvc3kupS0e4S718VKMCidGKC/+gj0E+uMSOIagY
GKxhVARaavdY0ALem8ghcFK1pUT8PyMK4TmDMZEi6+cPbmwOyCGEOfKp/Z2+oRHaehtxfRhGW1lG
K/WdUh9TVDpaJ2hn68uW1OgPhEYpOoDedLMFR1A/farT7FxKS2VDE23SAAf7ByeAQbqeZhU87Jcz
Cxt3zr2OocCyKkozubVL1mQYpTRrkYb8vV1yJEDB+5V1oPB8Pi2lIgMq+ghkrM9gNSwd69OoalSE
Q9pKuH+AfgyjirjvS16Gjvil5KlII7cGUf0yomIMe+eN/xqot7qtuVHSahTzltYsOwVFggD2zT0s
FCi5ftYNBRcEA060vk3ia6vQYFBzFbXwUY3WVGs9t/FkhBew8OQkoPATSpaImFoZ1ODVUgMQ7zs9
IeC3sWwO/MTR2akMA6AQZjMkRCHl57BBePOP9gQO+RaXbPDPom1UN3flE03AAGmKUWM/mQ486bCm
mE7wNd4s4xqkpQVNG8/e1cV6PF9ishQwxjSZb/GrYgYQ0QdpbDCp1IfYP2btE09OLdMZCCSoKn6G
OMfnwIGfM9qa0terUVqKANzAE+Wbyoa07NvP30vwUU1WYFS+hEafNQ5/GY4gzLljKqDe01fenoNo
bMSKnse4VPDTZxFRcSDnZUOtbV9aciIqtCTJ737YnMpnXy9T77qVjlK1s6qdcRUftA9Hzar0Cknt
3DFrVYaYQY1Fe6b98eKT6hfpBjjEy8o+2B+uwbEDX1Ccrie3EkoFT6fuNWwMJNtqdt83sQROWUji
/lE0/dcDO86WwHaEtQmMVcrMkdTFGiBDvgCn8NxYYCcdhFwaDG+z0caTj0bb88lG+RmrqMbC68j3
aKhjoZNos4eC6m0ehH4xR3O0lLkhSlNUkzKP0ZAfGRnqNNaZBftjSTkYi9z/YqlmFzji4Y/M2p9R
fckvpmqDIHCQ3a5xA8TQu7D5AQjkbUgydrVxuuyE4glPnoYycRkHTaKCLPDgw6NF7S82s527dI2k
DkLS/ODe0DOPZcDknTMo9VFkhb08WTmMu4FlY4KAkm1qepaUiPXLoN6xcNf6ZK2akN8cseFBTeNt
GG1KPsi5mfVaDphT1KMOCQis7EFfeMterbFGwbN1rlGA2Ldlq1QsaciG5Fm+YndiJx9ewZOvbnJy
nRGSUm7aoM3CJzB9wPAT7nP4OcUtds8V1VrgGRle0+IIIH/Jn+0aSlgSt37ZNZ8U4CAxHQ4SZNed
Gs2g3eMTg5xlDPg0Ld6fU5/09jqXPw59V6hWmOC86ztAIa+TGqJwW8/BE3TjURInHHpx0CFJ1Nwr
RbgK35B65lfljXQdjoMoHbLqw1YmtmT0AwdSLfusAwjlVwBgdhd0dyzvspSjIpsWtvdVrJnQjuup
h/zoNaZe1rDqiObZ7rIzM3tcdy4HQaZVf+QarRlBxiRFbpFbEUZ6coU65i1bEBSrZf+M5OQSf0xW
lX0lt4xPaoLUHkHVZAMkLiDao/FUSM8HemNcl+PrV5C8fzmk1mquJu639DwnH5h48dkXKAiEf9OO
yb1Q1/5KcWL0ez0shqzBxXWAqGEWmAqwKlSb5GePUo652WL9cie3i7uyMo/dLfW+gyZR4mPniE2m
bZ4PiN3JawYNkt/ZEQuA4lAW4ZBF+q8jGx5GCk9lde7ANL6wPMhLyJ3s16pcd4BaDYmQ0mWsumWh
Uc95/nNdg5B816233fjAIx/KImBj097ikrCszkBzRCIHa8MGZbliSFtljZw1MjoDiK2wa/e2+EUd
jTcsi2CbaB/sQEeu41OR5t30uev8QwQjCSH9Fi+XQ40Fjd+ZH+ivuDLikfH3JicYveh5WR+Ci4Ql
ZmBojr3kF6w20GiZKm/t28DKO4OvKV9NMyoUGLMp/8lw7uHddaEaki7Mf5YmcX0hEywE0EA1MvSF
h2XWzPg2IznatVZd4v2o2kPgvHCSDxM+Tz25pnhx9qiNVyZUY5cY2hobwVzRTIxs5+yi7zKvme+P
50HokgJm0lZ6PP7ToCjqN0/JBnZRkPdMeXXfBT7cy9mVgJ3+wdcEosWBpL/DLXXk+bQrscM41KUX
2WwKyDmTiPFeUgaETRRLRvAvjHNOKTxL1FWM5QGgioJ9pDnuD0SG/CJ8qbmbtagkbKgOylIhigQ3
iFIh078jxBvTEQOYyG0MM/d5hngRK2ddQMF536kSlnkkZpcIquT4V0RyH79uDt0k/d5fgH8R/MOp
zDvrXGCixCGu0d+lhf+CeTIwNdFas9bMD/yu97c3aOlgQIJYopOEZFA3OBMvZNYD8j6AmHBJzxST
lx2zPKHyeYg101rqKa80HMbhr1Z1uIhEXOdV69p4KX2TO8arKLlcuTzKGtWQEmrYi+bAKkZwRX3C
39yGXuS/ZaPF9wIo6SIRbD+1L1zthOHRNtnjkFKGSOJgRQZIpG6bIsIO3cHIZRsFD+5VtL7SkkX2
YewofC5bboUp3O6IfWhtwOxIwOVxQcIKMaLewcl+S4ujsXRb41T7wTUy3/InoIAmQe6jdUQaZkkF
WXX1wgdDvQMH1xkxiYh15CDQ6Xv7dCX1Q799Qsczz3at8YljS3CEjfn1c4wIM4ygbrlOY8RZrfaX
/0d08Q/3qfqLElprsHqem+IOlxNIBIA8eHfD2hvgE2WyMs7s9mKs4WX+ZQtaNDVitOG4mZYj2V4S
ac/YOnDurvBLKTUnUVKsulJ4L8OA4mhmWQJVE2nKIMj+RoUAY4jmy+BDFo8CR9KuIQmUpngb4yHz
j26qRGKTaJH7LWTAnDeC2Leez4emRd01BA3/Fo3d1vyQcPgoDbChG9xBnN7u0V5U/8CftQMmZamn
/nJsbohhjYt7cDdMw9TKMNywwYmwiQH0KI2LARLVRF0KNAEJZd8PDYB3+j6wj1/c6Ea9qB5KF4GV
QDvWZZv/9mQ7bbj3EcR72K0paQG0s1qYz44xxHyvTBFLL7wMXL0fqnYSXRWoGd7V52g2UdcRraCx
b+yZ1G+Hplweo2LJV767TzYtmbuWp/gkoJqI+HWdJunWHDi5Zk+sJRdwjpG4C+3TyxWNFmNf7xf7
Mr90B8pvzkzEhhUNvDcxSSqTrYuDQ4bcK0C0AH+f8BdBactIgCGfhv6OJeuZuWNZ6a6hhlmr4yOc
NiDyyZ7kaiAlE21sCJWx1G+bCeG+WDnDBqtgpOrUOP8WKxzeyHbvWg91vkj7kfOm2okT2sJ7GomV
Zlh2AHfkAHNRJkEJ1dTCJo3lOBDeLxwOCDPNWv4Dtndxaxad3QAJ1QohtmWQpyHsQc/sn553q5NX
9oI6iyHxAWbCYnWEuOtMYscYMq5W1t0WPU4kNOc7QoG7+qj/Uv6aauQX2Rt3V/JVv7oqTK26BxgB
8o7cRkgjOlNlrA46DT9BbEo0EoSFgozSMHkVFg5nSXUda9D8Drn63DDhopMjXmqcmTfCek1dsL18
PQ8IsydbaRbXRFbzuOIemXY/cVl/IOwZcDCMgo82+GY7PrasJOCdF8fbXROhxOAFZ/FxqejylfiR
3K9M2P3ePIY5U4Ee2474IJumBc5ZrcPflR2KybtN3himXfQbdrvzkIf9jc/N/H7pGdmVYrWADV8S
EZ0ICqopmmuU/ssl8BsAYm5RZYkpsjBmpOyFZ0RqwPf/hvj92DLp1JFlGW0YG67ONqjuzdPQl70s
fIb7nZeOiycFQ4FN8OdSWoMUJ7pWwTAH5bcN71wAElXZSzlycA6ntQ2BSgN47Zo5FN8O7v0qvjR2
7qsHxq8hG3l/GIEPxWuT+JR3pzXk6U2C32ivIf0rw0x78ZV6OGUMwLwWD9TTV6CwabUP9s4K93w5
W8U5OGswP1fthnTI6RctFg91zD8JSWhN2XZ80jjH+e9dCeYWRlYM8/RKNkWjuRqDALP4ZcwzBhjg
b1Z4IDZSUcRPcPRdNyfof3lCVWGrQ8VhecLKTbyORj6JHSYClxekJHnMwNJXj4oDFTFShbHbt7Xn
feEOUB2Ntv8cjxEBd/1OMOI6/PZsOyCWH0ZLlbjxe9FE6pT7fUkIK3QPKeCff8adDYlZLzvjAeg7
Sny8c6gdpihrG8qehKfes15634HSvbKNPVIpZl+PiXz17rIMu4PMlNKka8iJL4iE02N0fFZJZApL
0LGOaO+bvp0do+uTRzqHLAcwb8VYG8+gz7fD5BhohBRyjvbXlmPAJVEeQU72eWHiv1nJbI4dtoZJ
MxKDWIOflMnWLpB424cI2ik2jWwmGM4HdxgkePIe6j0svX48hDUk0an5cCIr9LfnbBUhpfuq7/2X
ryMeW1Tm41VqV5EE8WpOaqjFGUD2YoEvWho3O6xZ+DEOfxA0gjLmPKyYcZGa8Z9JACg++MjlkjH6
b4Fn1BzLP3HsJr/o7uzLEgeQG3hAyPzqrBCEptuJjbMon6rLHWEMrTrcIecQDJuLMk+uf1xi3tA5
KaRiuVM15peWOAeBRq4w2n15Fpzj3M46YkjtJNhJ52FBY6QoBr89SPzAqbGPCzbKeEQlq2ix165x
jjUJQJ627A9IgCkZrmsYlQxYaxlDnNgOoy76RUufBC6k0xlhBc2gAAykTdm4ypoekVmSK75Doc8l
+ACOtWiL2v3h/geRSreRicgQaZWXnkd+wyixVzsTaVaKlkXxWyn848GEjOeplSMSojr2wTPyEzBu
+C1fDsPmPtDf+VTSmuRmGb/2EDVydJN1+H646fjNjXFSTFcijsJvd5aNOdaJY6xlLxFSroUg9uvb
TM9gK+JzCjIBYETDY6/juL+vJPaL2XrPo3WjJNFiLpGS4nA+vXz+5EsIFxvjMaoenEsoRpJ+bjJH
woSQbkqvL4w67N/I5t1G6DwSrXhjKJAUmCt5nop2GuHEDxNyDVezjhp3PgnpSsAivY+0fcqYW+k4
R5zFaPEzGAaQCnoq+6/FTZ6KVqIoV89bJaZw8KkNsAdxTIGmsmC7oJhAPOBHdn9iMxQXElWwvs6J
jJuV1KwEIKHl+z9L6lHHG3dZKfaSLijIe0dfBFDE22lqbo434SLe4BiyCfb6BTDyGgGMDB/8GxKC
5q15Zj/cOR6KUVPhEztLT3P7SR9HIHGbvx01Ejv+C8wgHL3qrbJriF2acNkuojz0wgYQc7ns0Mrr
qeCHZUL1E7+kj2jaXb7Dg8FQNnHoI0GfaCawFBUsy/ecq0tRE/s7Da8PZwyIMwxjSfP/hnjxnyKE
SPwwWA53UsjxnfFth7gQUWlQRkuui/WjtpPM3tK8+sM61M0V+CA1QeR9XLZVX7H7DwYq9oqkzeaH
l0ua9PTM6pF7xG8gHVWLRoqWuCUOXFEZ+uGlY83QqqQ6WUACcob5IjBY27kIXPR6LgyDGlo4GaxI
NgBjguMRmTg6tDgfod2GihIFLS7Pg3A++4x7S9UTkfGc8ITCGgQak2VzuHO1qIvKQrpNmLzieADz
0GFfTmt218zt+XgpVlXsOG2wB1GeAbKXwJ+Kp0nJ1Me2Ln59oMp++z8q0ZOt7dbjt5FOKGlN9ZKX
SGXoUff2sP4L/qoVjwdCd2eG8DuG58JUlIihomoPyApZyNBXHb8kG3zo9D533CJ4qDsH7BWyK3DV
fY7jPvgqdPw4y+Bo9JuXgV14EfxqrJRFMjnzd2Hld7qvmlhAeOsEAFOeXwxWFgES+lX6rFvzu+6H
R6M4srXXtpp5dKZgoX6dfpvBS3e60mtp+QeFv+/GnlnT1DFIEMTNY77AyyGEL0JATeJsb0tXmkD9
IAThK6/Q6okW7WLOSp1u8nUhrhljyqFwixdvSQ9hOmFMTUuSGXZmcgZoY/hbUeVi0bZccfzNArG6
gOAOUko9QiWpqqRudqDUhgTf4HDdanNs1oEXMRGyCcbwqXEvGn05WFsF2kWYGkxPDdLJzV1HjuwG
qftJ7qNYt6bIiazDOWNRHSQ9coLYKG3fdVFgKoHdAA0YOOeVasklkAAx9hJz7zWOzIpzZhAGmrcl
+y3s0uivtRYiJJvi8lZOL4xae7Dv8MCD/vCicCFlLgn71ASW/hmuqeuwwWg45z2n4vtp1rvBHD1B
bZqfesulYyUwNi630qWPTYijZMvZV/eRzUC0YcL/xFvugNufeF8eeUN8Q3R6gfVeglF48B0pGsoy
WLWUUq49lTA/jWfGhNfPlRuhk1bG3UKg61nUK/hDE7FpBQZ0kMadXcL7oI4+DdaQu7E05b1gj048
OuSzdKbkufvG3IQdiutSEEAOw31QUzII+OrinsK2L75ZENZTkmzIyoGHPBRMyztbzbaVN2dwK8j7
bjvIPcyY7YC2uiGgXO3pH2HyRA9gfIXOwUoD4+FuVtBpm3OKm7Kp41sNs+cgWcdUGR2PWwbuRDvi
v97YDOdmE1pVARKjB0RH87Hs8EDrxsHseluxQRqZllTbg7NQyRV9CjCOKc4C9iCJIFFEjki9EAIO
jTvo4z8czt7hL3ZpTTePSNn90FkzTyxIdSJuRXetLUBmEqDPValO5x8P5vLpqYSVZSzCp4SVDsx4
52/FdwT+D2vaciC7n/kU7pDeZeDNmMnREzO8ws/ZozZPL5oH84gY/tecdXSO+hYSQkQ+gkhAj+TO
ydUjRm8ZXejH4+gPGTScGxxLyYuOFgFlqRHQSdvUfumL0An6k4m36J8M2E+LdG25+H1t0+/dL8Vf
l2atMVAPHkWWrZoJ9mCgdFlagGyv6yibqeAWyT2CrL+xewpbKlu7+g+Ih51Zfcv7ySVmHeQQb6jE
k3RFhFxJUmN2NXN8otjohtCu4J7oy5IjDTeRss90e60dwItKfmsHIIsNxzh7umWsv6Yv0A4h0myL
90tD8g0sPu5v+j/T117k6vdH/QU9lrs1LWAbitykwSCbPpHmELOmy1xv3LSPgBXSaryxinNkKfeB
mSose58nF5lnbkpjoirJ2NzqI9HROSozsf2FRWnEhKqJG6FBMAreXxT+UohtkslOVL80HY2SQz2W
H6BEVaVS8Rl7uazbeOiLf4mb6vi8r8C4sQPjNn+6Bc6NNjZwFiD6h7yGciFQt5/vM+qcUmlFaXGD
HHFqcqeClfXTFFH7KBDrVry8wo1YUta+wp+uQAVxtJlXU5W1TgNDGMz5+qC2BV38bFZhe0f9Sa94
IEbXJCYq8HpbOksxQP1FpXC6msXDu73iAumqqa0Q2rM3jGDJaWuVAwR3UTdfvo073PEFCzxE0sKz
xu1y0hfQ9aETb0XEK3ipzoQmbbrcaMkvfOuZqinYdl8SxfC0P47vaWs+ZkLz4hhrscKWyOWkhkiL
ZDEw/v3JC+gZdT4dpwRWD/31+ffhxfYGjIQecCgnO0WLGutZiG1yu19dFpmr7aujP5TOimuqYaKg
Ectxep1djyMN+eXnXNszUkbDL28TeQp9bakS/vBhAzWqKiMH1MShPGupp1QAPPKJeqIgX8zwcQVC
vLZTQxapzgdHWz8ywEUEXSaVefLcjz8889IbAYctRm4JnuBUV3BgaeY8pByqVwtlqXrIV3Ag/cWo
cZWqis6HBBcPbYeyb5opeCNWPDBEdIJxkD6IzjvrmymyTbgz68QWI0LXfBZ/xf2zG/EJYhbXmNbs
GND7pf/Fvcv/f/+UOKabYnJYk5nZfiNAxlR1VWRUyI2GAWpmg7JAzPyrMw1beCUIx21taE68aafz
rcN3tcjduJMVwKvhpPB5giEMY5R7/q7zyI+3kBwgOSeFLRv6+WRvZxwrVkMD//ZUMivwqKiWZUuR
JLYCJ2oCm/bTy3j84rJNFNmR5BUPumAUEJHnXEhTeKjDql+V0veQlbMvpVN+yjVyXYRPzkkAyEM/
8VDHS7K7R2f4eTevl6/N04NT0D6uu0KWKTuEMFpjfz0iJZNpyPnOuA0BsCwWtyAsS+bTvkH6XptL
g+IV4Ofd2lkP7OyKtW/y5BnS8g1Je19K4S2FF5KICZHV5IeXS3/xzImZ4iM94/U7BPWE6LeLXxgM
H6LykMTontodTkDZvigTSyHH8lfoeS3LKgHDh6di2BmL2XVYYXZLC61B99r9lGqlE5oCP83Y2z/I
lYkQlmWvCdImhWdjiESPAZY8ApqwzJnOc7AmFwObX3f8RIDGVQBy5asmtIuQYePJM9NAfIOq84LM
7oq/UUSOwOK1Pmqg0JpZ3Z5rGOzg0/SQyzz13m6b5ufHdfu/ruI1N+/JEnPypQRtimzYJrqtfdND
+2k3zv+TXUmKzVxQHdCFOcNwM+iLRx8b/wS5ECPeOhq4dtpeMxSAomYAmrTp5+J9XWK3KTdaGEbf
u+ewN4nKuN0MPk0TyFtNEMD0Cu6RNfd/unSoIV5yx+ejo/Q0Mk5s1pjHOo9pkBk7Rjf1anAvpMg5
W1obOxtogYFAdJ4YXKhW8NJrPC3s4y9AngExkz9+ppynWCv/xDT4yb1mzKpYBt2WHs3F60ienlWA
khswttMEm2/uZAFWukfKmxl176juC8pRplJMLagzMhYyvmsoLg1rpmPYRrLK1lIAMaDNQqwWzqdw
zdA2Op/5ard02GPYf3lmPTI9C7J+aPLxJxjPLy2u41Cf8+JPcHuV6RMZZAVIMWc3AMdn8NgD6BAa
KbtfGQolZ2YNE+83YqBPw+Spj9XnyCjMIDW5WJLKfdBqlkwPX9A0A+j0D21fMZ8VsZOOUnWvBkIB
wYiny+T+sD1ZWXGdhDewOn58CedTXi9AWw1Mtr3Uy9+n/aM4RC9ah/1RxiozyahkNxxV+VsyxOuL
8BccuarLqDAPjrVXOXIjFBZk8UAUSujzfuTuW0hsDoV2tKJedaDyE2SPYWHjEbVNozeS8y9qX0OD
3Sv1IixNx2EqLPi+es7+a13swVGYnroCsk7WQwK3ip35N3i2DnwL4KoSgCRm/9QizXbRJYIHRu6+
y0UovuWX/nYiup3viV93f1CIUQWIDdcNStBKwEH4aULdD+jRCuh4j/FplZopFzGicbLmHyufArv6
mdazXjjoEx61NjwsbWZ0utjGi8tFpjfWCGWQ3KKSCMpGARNbO/wPkATrM563SlOiL3OZnTSJPvlS
JcFfAuLCzK9NUONeqyngp/Nhw8Ez+zzU0QhHmwxGL5ADvDHQYXADdmrwei+pUFSCPe80YIOJ9O80
9DIdoGldmbza+o8uBkYAXMwoPfm/pMSXgC6Qm8j1Z3HrZR6BuGdQfDhD54aZ3c3yLGLBd+pX/4PM
JWK+GhSCLm5O1vCvwmFjB7VOQsj+HbRdsfPT1RqKJA8+jTth3lhVocWZ7uTv/8ZyphI+FgQzS9TO
tGcwiNEkzKcldRgnBJGiuZKPbJdNIQvL8O2fK67y381j7e0N1noNz30wLmbuaKQMR6x0jJXwMaO2
P6TBM4AvUhh/XLDuSF1qtDPilWlSpx4/DQgX2eaU5ms01F3Br9CyRdnTv6Yc/REnroGPcjNLgKfD
3GOqB4hjqsH80UbhL33scN2K7soAjfYaZcwL6QnUKAsh1ddRvaOC15XOxLXhZ3YIAf3jzWJuXyHX
TqTR/mbICO4zxZsWacreFm+jmSgcMASW7fLk8Hs/QuTos3AJ89h4uBNrdqK8Ab1PKfsgasvg2nB+
QeVJCHmimWV1IHb5LyODpPbcj3P+xEdCqgdU13eipwP1SLqp9XIZGIErTILmXCyS+ewjlpP3Qyl6
O7B79KrjLSzHw0w1eZftXXmy9GiuoMMb/gm9Kk3XGZTgZrOc6shrII2DumELmbSKMQsHuaXZ90pN
lwNFN5uaBVmyyGcYZ/WK3tQY+9/WYxQZWZdcbCLjB6YMCCar+Yg6myrFoedAIRNmeSAT0cvRxBG/
wWfIB9mqnz2SPze49uxJ0aUXh35LwFQLTN24/Xyebs2UeIpWu9B/8QQ4iSoTalCVaEP35XnAYRLT
JNDK+tYXl3qmzaYo+pYRVkBv4LSypYDM/FqCWUGaaC9GmBre6KV5uLGnMs7cBkmYxq9mllRC5izb
mmiWxB/NVncliAUa9gKYmMLeCDvSW7UtgfFC2Isl5mKZigkO7+fTO0G58OLk5fAMV1Vu5o8Q2ztU
R644af5voaEU8yycgs1oqCvwtaumInX+lnaNhlDLdEmM5QhGHzipOndmw7r1SlzZwGSoSFiec58G
zIEWn/0JoX651fHu/1LliSyxvk3uxfpZ6Qn7ETKe8PQb8BxYu+g5ukJ88nX61b2Jcrcidg7HOeJO
OzcOAMBU3yw/CcQ4eV8uIeWG0atTg1XusoOIpmYffXLDp0xz9do3p/0MkXnlv6sr9sfD3XBrNMt9
B2JQhqQD+ESRIi4icQMMMLNdWAHUuGtbGQCdVdvhbs0ie1CWyTqYftEPYITar26V192aIQMhxFc3
wpzw1i2Pvnxf1fxSAYB5gL0aVZ9vJNY3MmPlHXG7VIXE2Z4Bg1kQeqjjEFdJ3pfFqBvVBUjt32YX
EKtxsYZJNJ15bbdJH3KTT42Jhnti9cEuGyogYsnKKrE3gbw2T3bhYAyuXgochiTgrdt1efmX5ral
SYBnZ1mp2ihkumofT3aLZwUEFrDohqIAhh0ZrUjkMKDVGBylY9rGRQNJvLbeknIr3P58pS3mpXI1
ldIgBHmzxUmKWeI+0f20XM1XFRWFGaMzFaOxsJcq365yRBW77sf/13HGdBtrXJqjySTGB5+Uj5vk
tRbByJQVjfCtTnw2Frd7XzBGomNjw5I1Odq/nCc+1AMmZXXcqF+Nq0qFyRCkGDBlGscnuvwefrIO
l6CrkcDnsqlg7yaeZ1qLRZIWlB091wNYwCVgy7Z4t+F9YuQDtlW4q+Rot8FA0u3qFO52HoQ5Q1Ug
/BVsexX+z9A86Rj1q5r4+vBKlSUKS0MCtQk3Dpy0GJGhofas8dY//e4qTMntFInEqNR6TDKZvVYf
5hIrT7cMGAp1KZEGluls6q9YW8CrrhWv+BJFangppRY/lArgyVoChGHabAWs1QtYQ2LSZWm+5iQf
ludOangXsfR6F9PIdfS94eFbJEFpUq0I5hFp0aCgw7Aihl9jpNaCGk3AaLqsyuae1frSfUTXBJyq
KBEL8AhUC7JmeNJCMwZGrVXxKlS2qN/q+lYkMZYabe63EyWoAr4oDfxxNS18qmAQKp//I2RsMrw3
yeUEkjwBidPpCqRyO0YQ2LLSIB8Zl11FJvhSjCzdoTJlXT3IkqgIjRQ/pujZDLVzv0XkCywxHP7Q
XOL6gnTpwZg/5qaQ1LlfIcsfrWisTG9OdYu5bll78SaWBqedOkyecz+wRect4xQCL3t/WkYwjJVc
SrAT/ddJgtQFNh/oXx2015OajI+fE0FhWLMZ1JwJxgsSpz7gMmPMOPkx5nv5AcrOyj2jcAKa8d48
blo75O8EBjgO3oFi8j095UDGbyeHBlHRWbEbTxPvFW/I4jcmlTN8RKH+4kb4CQt7Zn8sP71DSWEw
pvniqu1pRKi7EorHIU5glMxnHyNotvNnD9Gx7xs1nZjzLL73rGaaYP2ECRrWOT4NKvTwjPGu2qXl
z6MOblBetDg0PvtrRGEgiLsFItni4+B7083tZbpeKO/Isr2+vnVljsfRolNFIceUDqJfPss0UwSe
PE8M8CPAPMx6ORMAtEAKAj9wjF6fgg2LUGY+pG5Kxy1QT2mqnynvk8VSxE+Dgw2C5w82Bgnp95QG
XmQMHd4cpGTv/qfne9JCv7I1t/UEO+oHaV0rLyrkj1cfdy/E7VidXtbGk5H1rt1NBkrDTGNYUM71
zldwjYdh869HVEVAhAwxOzIHAe89no+XL/b473KKytdFejPC33APX2PrKMPwxqK47hMNwg9G4Jy2
Xd3tGMvRoRLprznJpBCVNPTbpXPnWzsaw2G389GV8JzXAMs5XK8f9Yj5drgc0teZPgzOuM6dySAj
Xaq1wPX/mXim0S5Xk3PbTsg5Ga16GP93SY30zlGcvvdFgneyFS/MaClFQxTveE/ClJq8IQ5HOfDh
TaVin+nC4BJherB5mOYg+Kjfzdj+Wmi3v/J6HChDex7K4yDuw+WnfzO81/bKpjCKPJTKdyJnNWNq
R6DXLhLlX9Pmt1bbb+OoSc3L/VS1cYbEJ9o2z3L2kcA5k14ncDpokgeHcQm0OZq8Q61No9nVxtKw
iIs/hFOI9wu9k0inf2Qhc0Zi01Y+TkKqIvPahMBnEl8Ea+NVZnKXAoTlKJR5sOxx3D0d0Dnvm3e6
hS4baGkRUZRCQmzCeP7l2OtpEYIMIkh13rXA9i6OdxUtEyVQK9rAfCkDtNjDhTEFBDTxZpr03ByT
EVa7XNjHlYHuirVz3yTlurLbZvGLr2UJmctvzNKR8hIiLoHkpcZujh/3ocF2pgF5ycP2aXSnT/v5
dQo8W6Yw4kAl0/5n4fnn1Hy43bWcC68B/CztDQOcrXTiKwAQBFJGWqRHW4j9yBh3RCePk4TOuWSb
yzCbf3sOusUTxnpmOX2cE+c+ZF2bLJ4VsZmmpTvccsoHADKTehkl/cG4y1EtP7FRVBBbFXZF4BRY
dGOGg777Pigm0fl+p/nT+FogWDix2thG4UlQJq7YlNnusf/z24EmQedEmLHgZ68EiJwtzK48gA9M
dzrn4LFttgARaYEkkjlsImk7KFxUg4dVotEtHhhqQMC/uerB/csZ8TMNs75iukmieUVP5RiQ5xNF
LDgpeFsNdiv9LwmU8z6MPyTNM36fLWLvgIOOFEpLbYClP4s51q1zoMtPWrDfJxvIJN8YgI6AhAbA
SfUBnEgoSyhyZAMSgn31X3R05xi2jpnHETS3vH/sK1KmxRUvZgTWgk5v+KqGzhaZPh72KRZ+rnaX
woPxW8FNiZJsQ9E3N0PHRxUjRPRV0Iz/mwHKjjS+rXN69NI9rucchSfX31pQnebuvYtPqGZIu3gV
RKBN3LEOnyJjJwJKGjC73Ye0W8WYU7k1Stp0Hh1PE/4o8ZwzA2R5Zbmb9/5wAK1R/avk5kG3lcSA
Gts5mZ6uvv7zHKN83XteCwowxNCdNDDNPQIFehz5dA7r+PeYn5GPWd4r0CUCbOGRml9H3nQ3Gxxv
Rrl4wywlIeswwLmiNHxVna9E35as6vhcuDg7eOjFCzzSQUJmByLnYFHL3iVvylDnUBSH/mvGlmu2
EBK7yiyJGrAHHNngXDwqh8TeLu6wnOaRrL8WAMHmtX6/kCsj/Gq4qd3m0mHZ18Eagy5phlWgxQON
ShFhIaEuhQgcBUd1kKWpQpZRIZCVd7a2jvaRAbTWtJ8OAKq9V9hhJkLqq/0ByfbE6jpepQ+A7dpf
puhadBuIiiYkfA4XS3nMhGjeqKztKaII4K+fDuqvwmqsyLe8hL3orY6NRlFpw4j5/osQ6CWSXwCU
riQxvc7oYfp8HecewfBla7guimsyO/4dh+bjPCcptZ2tTIvpdOElUYkqJzw18SU+RcoCdIeCBekG
j68eelWhiFjijVifmeuD97LPAVB9MDab5ljsM17rr0m7VWYpMRHXWXE2wkBoN+xx0tKWPOUT4Cn6
k7TB01J1L5n70JEEEEIMO0svujL4fMz1vychBVrg7AQOxVfl/BFQpWoGfwxvbx8Ltu4o3CsnbSnr
898kidTv0F/lsOl0QrggC4J9fbh4bFAabxc2yf8XxN8Qj/dRgg/IF9uxOvGPamL9oROY/7rsHf04
uRms7SwNKusmI8Dxo2McQrUlgb5EI26ZGQnSmvy8Tsd0V59Ozu3cI9h6CY0cFXUv3VozmJk8T6eM
CmQLAdFbNj/Cw55c/U7Dh8rT0ZWzjnmhhJRozxGhXR4QfgpQ/nUrWxPC8if0bbPWQWakx/vVqxxm
1PAbVOgRrwvDa4RORpfnBJVtD2SvaXmxwUXhdIsgukUEdQ/kFJb2bqPOxXF86c7zQT68+UQVHM3g
eaZWpJbze6gB5mwYr7oBpc1vIlB6ROS/keCC/bo+NAQRyGtdUx0xuLAreR05ZoZVUIUZxhmTAO+6
Op2gMNiTPvMK9nl0XQqy2ohVTO2be/LJ3c52CKJcMa2MkRldjhdH9gmeME3A1ZKa9gFmgVGn67Sd
Mxfluagijl1dZxboH0HU3ytTJW/kK8GMObV86Uzqs5o5N8AX1cGLrpJ461jHb724irJU1KdVRbAT
cVqPWC7r8Q8AHIQrIJb11w3xcvil42vBzM6Xt4oL99BIihTaEw0jYoaWhCgGizC8iEO0Fo8sNt0W
8JfjuBl5VuFGBAwsJzvlxwUG+DeY8TWsXl1LDVPUhDuRrugOI+oOlm/NTTquROLbLSC/6EZDEbik
pcS9/YbHMSPvKp/xajBqMVWam4USteAVXDz02JrEwGlFk1GC48XoUkI77cO53SSfz0TS3LnEhi6O
1tEPYEDRZC0aDEB4LEW0pce+2nL0Qwths3b9Ar5fCn0NE5c//Ojhvpd3qEW4XaiGTmIpQZEfylPA
1ZQ8C4/8HDfZrjr9cwf2UxBAGVwg3yaJKSVVGJKznvaxlH1T1UcLdikud29b0dPWXLwZSXr9OYrJ
w3/1j8xgtIp3awx25aQrasgcUAmYNYEjeSWxCw1xzptmZj7t4Ckr1R8wJGXRD+ehHtdf+5c+J+ek
ItqAFNpkJn2zpiOjYcYAzTTX82hnKpGkdt3qlzCsIL6Gc5usV4hyXU21K1ZyYVV1AhCgfDMx00aB
KLN+sJJ6vPaXOImhD+nWuPb26L/PoasfRtfV5uJ/irhlb2yoBwZtyF0DLVWxbnZRvWDVeBQB6ofV
zdq6bvU45rNwcYwDcpALBTz1rYzeoiKBwsB6Y/WugLovxnS5xbVQsERqCImXf5Q/yKmblIEnB0bw
dScBI8KcTtYe4/JeSGmfcZxHQHzNXuo4HF/Fi4HTkst3Vw0VmtVXkRyl54zY8CQcZZqrpBEXm4te
b/e2qoj53VRE3LlpiU+A1DkWkdJHTPDI2PeVUZeWqPI8mQsTVzeMu3oyzsfBNRsHfohefCTDFfgA
pSXqMY3jrbFl8FtySzxwIYHGM5dShXCkrVPaUfE/lvUk++ElRM3HFNSrWgN6B7eSz7ncdGBlrbFp
1utul2JPxy8Y9lCDTHM0x55PkvKUI15G5cDZwYSrzQ5Hbb02TigvDIYjBa9lWkY03SG5nYLPSijN
yoTrYfzlQ+usdmwCVaRHzw59yXl44X0pq5+lMjLwgE03e2ptpjawSKeBdBlt8J73ltKXov4yU+k0
7w1fp1+L66FAjFdiFW1NMDo5AZZqvgc3NQi1ffpILEv56u7U2mxR6ke3AefaTJ1isGxS2xeH9Shx
jYdwh6vuq0H0yk+yr/u5UY8fuwi0HSUYM+sG/vZ9nhtjfGcUS9arX+NuHhAbFhGzmx6UlO1PBLNj
xqO5D07pKpDVx4blbHrIIliTcPVpU3tY1ifrbdOnrf//XX4ZJiMOs23oYnUS73JU9PxevYa4I7Tb
879jXQwpvlE4gVtqE2bsuGbMBBXqxKbD8QTC2g6v/K0pYNZf2h7vRJmCdctgSspYYMq3Y5C1vH6E
B3Wt0bmtV7yWCpHLTa45GJGhAstMztfWJkfm43/dSYdS2xb9WDrayIbQ9XHAhkWcAYNugerFP+Zs
aHnpz5rNnX7iw1E6JWyfwfID92MG4keE+4bjrIbAyok/noVjMNlNay8dxzwFmqaVaqncrmA8mxTQ
S6JPjZ0uuZnHPqsx8QIIe9Qa2soooFBr9vHVZ1aIk0V35wpzed02vUeiQsNihdFNJB6H51c2E5v9
2tG4/lT8AGBiJJVoIvltlgsMKUdPp687AARLJKqU/X92FlCk+Y9Yki3M2Ur9nGWi0vgZZfkmqT7u
OHLyS9KDWRIloyLepDtzArwNLkhyuYPJorFOMs3lcaY0GpzrhMTdyjHLma8zPp/Dl97RHai7TOpe
9B8GH4u+PIA9rkFkoCkW8uF1pRr8l4CS5J9XCwKeq/3wRANrBo9QS7hqtRRTCSVweIEiZIdZGZDH
znNvcp/EF6dXn30UZi7MVey4vYjM4hWnVqu5TKabNGph5WtHTLc6d6UEgVhxswRC4It+os/8Dwbe
TvFbSoEfunk27Mla9IUMCjvWOiFw+m0Ro1GRQpRsQKOuZ+uyvFh3vGAmtjY9jfPj/Dw2RnI0Q1Of
+fRd4BMgfkGK8s2ev3NEqABj43440VjelqXgJuxUveTfPp7Jcy7bZcrOWROELRxOJXeUWwaOh0LY
N6kucIcUcpsHRt673lQaBuDhfwgDSskHK+qYYhfw9oLl1gDRlm+V1/knK6CCfc0dzJOH8XD791g8
BpZr29ykCH3l2mlhpfJ3A4/PSsZ+DYu4BfvEWcvfDjh3zDkn0Jcirdu1urTB5C+0bk+dBATVuRem
qHhutaY/QIP8g4UDsiBRXTpp21oK6tv+IZfCgJifP/ZHmBUlJ1baEPwxmPFbkDe/pmRl2Tce3ZGE
gaELcS9TH0PlD917Kkiy2F+sq4iEFVev3eW6QJflmC3tI8nxDxV9OotN77ePF3PKs4p+w8ywDZyQ
a4Dlu5FFB/CpKf6wf8bD+CQzP1nXq8MWl0QQTYIfi5xLoaoYo9H3WKXDlHcOkkL2qghBtZNhVozK
EZGsG83rrSxoH02k/t3W2nsrVvQtGO2LWFxOSS5evXrcjcaGqvEwS1aLpaO3BsX8K6YDfof1DlaR
raOTgLfBe+Xvf71cDb1xn8J5pPlW2T7v0M/PTnubkkwCh1Y0HJ8Cji53V8xn7YbJR7wU57HPIJu9
jV42OGTGmf+D4pMDYnRNiU+/s0+EaZAavhWU55PHqSYv3jutGLjofItdmsu8Ru4v1KixGFsHpUmb
KukeiFt2oi03WMMTX85zngqW9ZlqK3UD38SMcwZLzAaY1tsNKYrPHJ+1v3cpaIY0uICkWi3ltpB8
keG1ywkvJDWEysqVt7WCuur02VVxubyE5GTdobzdNCKdanfSBIO6rUn9agR+u55CarYoiB9WwlBe
+FgREZ4WpKp0qoZypGzrIKszKZFgk7FbfCrb2LK8roca7lxDXbISPpO21cbd2hYXF+PWNtuDLh3s
gR5X7sOXCcFOfXpkfPkS6jW2GFAjOiC4h6b25MWHwH+SUYW5SMrhBolvvfk5vQd67GOTtK14Dyx+
bn0R4BI3dvRLmyoMPypIV6FYlycRekk8WvWZxFiVFB3K5pg+c3tswU6f2ygTQ6AdOR3d6D9EdrCi
0Kop7lFx05rTU8j+ofOfUM4eSwtLIjQEAF6dghiqaTzlesgtb57562OYDUvUPtZg8HkdP4/f7HyZ
Rf7LRS7tCl8YmWrluWEdqGithghIfx62J91ZQt9y29LGWiWIGFohgFpf40wvDXVVQLHyUjnXYGQ5
TIK4t2ZpSec41dTE2WwjEvwmKd86e2I9v0+dyehudwst2kX51BUihtNvV3SH+okCvbCPW86ts9mY
jN5bgSZqdu+GeoZFHtafLGT/fLpggv8cLJYh22vKcOG5niWTufiRhRcIguVqcFGcup6qj4JHKIbv
agnQ1KnEZ6sUhpTAnkH8wKFFiAc/U30ppDx0veyp0msJXD8lY8S3pdRxDZ7YL073dL0lHSOP5v5I
i8mrGMq++Hg/QrG7CEcsmIFeQhQkbZN1sqyj0lMRqVMEjaPiCPhk0CZ3CEehiu7NZOr7LLfMBpHQ
fsSEWJbpE5C1qxnugnDdpyrtKryY0P93Lsk0NgZWeYKpyEnUQfYix9PPBsb0XC6hm8GHfJH1TJZh
ArX3C63w4h1Hb6+sixXqaCaLDOP9ewqxTecfOafjAZcyK82gnWlS8D8h+spIFh5xo7WDyIXG+YSt
Wv6R0+/q3F/fbnDeTu2zhVSpntldQxUYyPAotdtLK8MituNCdUmDbgZw7JroXw7YIWpTsEBHeOUz
hkmfWes1pflSMVi6j31XvjSsljsXaLPJzQS4hUPQgHSivCMrOVO4JCOIN2CWgaKus0sbMyWvLFxm
VOVgwCEaOnIZXlOKZhBbE92grMq9L71BWlEijMzon20EiMybO2QZVAhwkfc2GEdrqvlsp729DxMA
KAxJwNkpooCjffn6OX22jHz8p2ZVq4YuzEdqFz4oARz1o1HiC+xShK1Bk7sMRjmI8/rJVzELniko
ryTkoePKR0qsq93qRkJRaDAGSu6ZJHcRxMcXrv0jDtriFNSqHq77dEqtU6V7HzNvc/sqZjmQ7e21
nTb4DzPEUkM7Jbxou7MaurmQoBJxlks87K02QOjdc3e0h36v5wScDK0cqCFUPAGkRe33tAHe5YLl
AdgyHNYfmheLpwet9ieWhNbMSViORTb5pOURETahuBA3k7f34Y1b6K6ZNYPMBTUYX0sIudZAcQNd
JWEYRZmukmFI42j+A4PDY7X4fLa/SUtRPWMn/gMSgN4LTGJLrvf28tzFPmkh/5b6X8qQkd111A8U
pB+K0iJwNCRd3lu6Y6oA5H7k2nVEqeoBkkULs/+O5VBNf6+KIHtiD8blVMVX5NyAyBVPfbIFd1Xg
nqzcU3aMkqSVNf7B268YF/71OZIUXpjKctaMZVOT4xzzDdw9WarBKcwwOl11YOHGdzncn8n54r77
v+NQUSHC8NkVACRLdg7xgOq1Hkghxou/GfTVkNVUEZ9BUxJRSTecZzkA6TN/ozOO/4hsjXN/X1ew
i+1j5bGslez3OCfnMXD/o8500LfBtntdzq1msPhS3wllpMCNL0bpI/jSowjfex2jbSGPrrr0NPhJ
xHK75fWxjNEA98IgMLiDxzzblWVb0oGOjBON36qYpqi/NmuCsHZUBYLkMD2ArAZgZo+J4EU8CLS3
C9hM5SJ9VhiivBsrsFDyDyP7Zsp2sN4TUaPdUgp+3rNp7Ln9zBxrhhJ/a5LJ2V0Mmimpjyj4qs64
wt+HVIGIu5JrdzpYjIRNPp+93YhE9Rb+1JRk8lRMjahg53Cs+aeN1w9ODNYg8jvyFX04ofq5Q4CH
7kb8pFFqDArQGMYdtV3ELqrLPNzqnIeMGJU82KSzKyiPTbkO/fPFWAwdDrU5JJqmtMysChkKKyb/
KRvDBZjoLkroFWDB/LP92ZLy/K6P85feRid/PBRqfRDmp/p8991r5opXEYgEvORtAQUinb/TaN8b
Nlc1imsdP9xB0Fs7CgdgRzoQPQGyXa9pYvVoBCB6UKjb+jM8qqgbiq038ELxkN0mQyDr5q+lobIo
CSPDd1IDg1ZDVoCNmbCQ8h7viCP2knoASY8fBNzIdwcW/Hj2MU/U1NWIMVaRGqNL8yWUF6ulAvYm
auB4Zg66cjTjRp8gUFS9YSQc1SmcE9ReB7/wVo4ODboTqp8Jb+SzerInIyX32qRJrgJdbvla43ZZ
GtW7QwgvIUwR8lVhvBDAtYa0ejykj5bvc7GH9kLrmyybpnAC+bdDA6QO3dB9VhbifbiiJeTgqCQg
zoMLijvxRHQ/KuY7tkikGgeLQij4kCWNyDuLgnobStjEQ2VQ/oipfwBLSvbbX1N9DGIAu1/7IB6n
8HMvbtn7afryjixU5WQcITYaTWZmI/8scj0Fp1ndadMsYVx9LDk629O7VDnbSnVUOf7w6UDVP3MT
9niCArHqofuvjUe1qI9du5BrM0Idq936gGL+x7GNAoHWJO90FvFu63QMMb8zy93XuK0lC4YXcnD5
bwRkEscXYcANa28zaJqz/IY5LstlNxRHVn1zlSSE8f2NbJdtcdpdwZB51iyxZjkXpwonJFfRBA08
JYZgE+N3Cz2xnT0n//9hQEX7swArCXsr3iqi+nhAb5UkFHP5RQE8811Vpm7eAIUXstZ+Gn8+J13Q
Ygqu3Oa/Yn41aH2agAsV7RWVhfObRWM99DL2Ni6gkA0OY3IxGrt8wipfIIm8wMGZ8LJEYHUf93yW
n4Fd+usGIvnyId3YxaTfLONRcpxgBBVKFYAflIQvghZFuVb1bfG0+V3DaDRLom9l6UpK2SGV5ubD
g3l66G15YtIbDMtiSB57mf1gEzq54CB4dQCiyu52NLwUFCYlc4h1yy7UdnRtjn1uuGjvq3qEac3F
gNqpMoEB0J5qKGBDiwh2+BZtSPASlh5DgarZEwUx8whpe+vAVl6ifkKb7sMfNFoJIiNjrziCHvU9
Wr5CXpcP6qgYcFeS0GuyytUtmYga+vwtA6P0Ef4azcUi8C4H+pM3qqPuY690wtHx0Q9cCDQyQEue
YWvEYK3mUUnqwSKliLrPUqlzXTnuyvSormF3wTKs2UITu9slrC1v1xiD0OhgGJKJPo9W2wGeT3JG
PdNoNE24xkyJOZ41Xl214lR/pc2QDds6YZOy/anlcLacYRfQbJcWp7JKxwXJmjlZDvc8eIPmA+iC
496Tp3PIClTuBQb1CTw+tz+qz2TAZF1vDqiaUAVriIHCBoKUz/utB4QdWbJWajsh3ZQjVfL8aBcX
7STk7MWTGfOq01sZmdK10yK04gTrNNwc/NC7Vd8Ny5He4YB0Bzx1XCwg+XjIpKN8hG5ZkJOZxxr+
XJ/NeBxmEtGucgWytg05Ky80GFWDL150rKqfmNCMUWOUBe4lP4tLtTnVErZOQtVTtgrz3EVWlsfV
c/6vsInXYN9iVk/05Weg5sfMxZXGZUxUa86vtbtBLllgm5bKI444Pte7b5b0MiA4dSlb3UsSNy6o
AQdFeRdoQFuWGEDrfO5QXD/QXLE1SXxiTmjtwtckfr8OE4WsxsQl43VdEREJMMASFQUd+Tibd7Oc
Yz9bXy/kQ5+DP6YlXoqElrXNnQgFJ2FjC4yTrV6n8YFZtvgwMDNwiQ4/2bDNyGT2Ky+TFTRZedZN
h/O6xQ/p9MsbUamZ/r1gYP1MROFTZWwsPQFO5oQtbOKYBapbOqihMFQbLCCIuc9DDXXbVyqzewaE
pE3nq2pYJHxQIFohpU858Hx5Y0SPZyFZTIVolKsJA0oHd76BsW4+Flk0uIMJzWNJpy1sQocH2f9E
1CxTZ42FN9eqTsIM0rM4j9FcltpH3KN71lsJREkQucJxPMTp278irlU7z+Sim38qtI1lTeNIuFjS
xg9R0i8CU6vfsf4KTTbyPG/yxOSQLKmFDY7gVDs5KoyXxpowA73QvUmakVfIf5F2mmVYg7FWTYUr
CycIrngjWMFUzYNAVd81ndXFcT6k64rbxUe0DbyCQNChp+4TqcZbtos0VQ0BbA4jPJADh79wRKSE
43Qk31jRo2FpSSjbAzqwm9Vo1qDmjwwNnxzKLZ6ynFUTeA+cjbdp31TkW0pL0JnDKh08H1QHJ8b6
ucutZz6B+lb5FLfbRlrExbMLGEPu61IhzPObLNxedbyxkrqgijlIlrFqNw9EQ9f130UTbO6LW6kT
fWpp9iOloBrQnqN2PEJZvc0pS1t/lGCKhUAkIs9EB5ZaJAzgGPE7arqcFG9ySuJ/Nj8RE1H+v/sW
CXVwNGbCqEyI9pMin5rGugV3ZhWWbnX61qK+gRfptLK8YeBN8y0zhhDg6w0A7hnsKictEh7Yp6+a
qcx81CJrydQR/Q32qmKwjZD/leDEvfTtf25y9ts4pQn+p8/dltKvhcXxbNvEyxUmF1PwwRnwK5dj
j8INdok1pgHMj6Y2BsrU+h9PQv2whUpDlFE7iAxH/iZ8QzOtEyF93l/b/s0KXdAVcMRY0oPQey64
4Tz4EtYicOnM2Xn+XSzpK2iMD9vFjnP/yun5VyQ3xew/5X7jYfElSYrPU5K7G0w7czQaA0L/czQr
RvLNYrbiSwKWWyjCWOwg1oXnhG8knj6AMtXMvNXXPXKnMylvVIxuZhtolsmsUQgim0VyKtfLxn7P
4JNeiySAaltt8oEBSMqxIyXKribxDw9d+scuSMhylFFhaS6gp6+02gU2G7rzRPW9BXYX7k7hlYAd
6mrqwuQaIE+Ruaw1qmKYKZ5Qn3Qpoupa/yUwPqB+7rxJoPCHrF4btJVQ94JZSz6F/eYUWp4od+CY
kDntVDVDbzcbSPbWLnWLZ42wYyRsaWYqs52B3pn7Obv7/5O1W4jV8AUAYGNzEoOKpTL+ywOSfmGF
Hp7F1f+KrmB+EQkLHX6/hPdveDo066cLbWD5jRKI22sIc4LTXMd3JqMcQk29+kk+uhdI8mYf5nvd
zVYxzaLLl7uC1JXIb9T+l/1rzABcIBE9DG494o5pOK9waIEVhA2HB341UmGB5ztB4E3mXdbOevaB
DhMSQYTIePOIC33/ZO6EN2m9qbBEoKWbCM5/01SnTubGsRGtLBXxrvEzRALTj6e0PDzZFpBiaIdF
KgPBs+cu3DNBvBvNhtENq1QcUNEFYftFK5eh1fHIGXgi7CqB27gNGonI+en0PgzFEU2lvp8J1RD8
Igx0r5A4+Svh/Ojl6UFJ28AhpbWCht6U/fuILkvF0VCI4m8GOnnsND0HVnD2/Eu1VzxZHCdnj/Qn
VE+2yM5lnVprhPgSDqDNiPoSsKvzDMp4zpTYPI6wla8PMHbdBBs2Gu6XifoEsnp8XOkgUh2PCRnp
YfFfCn9/nrYZ62drPI0QhZhGgt2gujbsH0rNEFV7oYnR5xm6bFMmCycCJb6IFS2VPSfxIqeow11T
xCFWua1bfoVoWH6xkeOV+m8Ncb5kQuVSoVeiGN0J1TkQq2K0w6mYN87GD9J8zeIplB7wmwW+GfZM
Prs00YxYkaNKzubymN/cBbjvQogD9sbdzbwAkAwKWDsJcvVO1V1PF/nK50jyGjHjHYjVWmu52lpF
byyf12PYuepGiZeHQCMOHHsmpAIixd/Hd9VtUdreoEQhg3asFVa84FTAKpc+RWNlQfvFlW/HHkEr
KEm/V84G/YSezhfvcCv5/aazr+lTlgOLLn+87F1rZxI1vXEOvUwyIzh7r3EmvueFKobW2OCEBNbk
jkIZtO15ENPV8pkUsYdUzrv5NniYMZH4l1GDo53z9zBC6p1dM9QGbENWvs+Z9wGu4PlTOGzCgTZ5
z+caJdtk510ASrFJFw0MbL4AHnkuKMsYH1v8fePI1TjAuQMkePJG+BYFJnXQJfM/1YyUb4f9DDgD
RaQ2yJyPiLzhRJ84LuGL0dESsH3IUcZD9CYz/+QNEHpt9CZ8NM9J0bS5lm9OuZH32T5M1luWtDi5
ShPl4zlx4mlDdkt0+KmjkB2c4olohCvfOu/kg0FQKp4qSZijuSvzv1Z2LWxTz3slg7lCd9i1EjiO
SdmA7yWL5MtUjk/Hh1ZQ0dJjlU9CyDGR614PZn/B5TIAyEijdQuTWNNnPsfXaKX1iHJdc3eAdqbQ
Sj2y+NrzZlEvDvddoBb+t1XnApFhCfrylLZHZ96p6Ek73rqgNMCaUaVB4VUdaC7qSb50YgijmInG
0Bsovgykk/72T27EcG7SQ+0x0AK+777pd28t7bAhNRfs9pXBoYwOLL/BCFqUQQgxqPN5t9k/p9u+
JnCgf1ej2YN6qbIEvbwzgPQweVs5iFtxX4GqGr36bfwLBJIu0Y2Q/yF91FqbMetG5AWjRqdVPXo3
HaK50ON0S7CBgHFN65jfIfyBVIGtzwJCpDBh7WV/69OANZ14ZrjczcBEg05OZ9aQkezdD8CB6S+1
NMk6MUQYST57WasXdeSzViVi5fmPwpGPVauUWIc+hA37dOQEALgEpg3SwKSyunXr4ChsBNhqKbUG
EPLumlSIrWqRRStMW0Mvcf6PM+0y14RNNCZRYDkKppXr/zSaUjXm2MTAb86Ag89lAEgBlrFQ/mRo
u5oIvYB9dvg6/D5AgugsZdZR8L3vpj9LTX3ASO4QnAkNVjpfR5l0eXDA3e1K3bbs9W2sdowTc4jt
H+FmZCFzJqcaiSNHXa2N2YKYkFz4sT9o48G6xy34v97xo2PVnVGCYcP2L82jRenNjJbbWqbLwzhl
nxDNp4MCH3k4H8yRRGfaRcE1Vy1slyl9AsvtxNdXuihTCdx2Lcb3vXm1ZUmXwL/wprFmfruLqhob
zCsSw1vs9kDcTmCg2l5lmbx0D/AxZOoJAAdYm4pdI983r9n3Z/BYFfVy8bg0wmDZgwz5YgKWZFjz
HsTk8Ja1m2Po51U5c9ga/tf1tA+UTalyxwNbYvU68OqiRe8LV5alaK3IqQG+wRUsQgk41SlGBf9a
CCsVadySwxYOkRDL4uHY5efIfPmnDsw9zHD4dWApMK6Ya5p9uUxqLYlzcRjL4H8qN6xd8Te+htZJ
L8ToTSnsjavSRQ0ShSwu/0Z/cCtFGWw4MZAyaLDpDrmBlnDuOY3W7PA/g/ZNDWDtC8C5UhrPfKKc
G2r4i+8zJYSV/d257gAacx6mhmICUVRzkTGh4vSoAYqDveHDyruV4ZMBUMabSMM23TjYKr3PhgPs
sFiA6pNJjCVbiyrIvkPl6nxFGrSZ823bNh2GyZEoJ51Dp6eKOqyxEC9f7oi82O/w9UPYXJoVKfXQ
X4EWrExKKd8MycTZZK7ibChUpp5C6ZBjsrsoiGaDtzUY6vvw5RlBGPdtWtTsEGpf1V+aREVdHzPj
p2f7ZMYDHibCVX2b3FVRBivcMixgeWG1V0+m4MMgyR99sxjkKprohrAeaGc9SQWxw1ahbU/DgESO
gzp7K0/Ik1vU3+vKn9Be0t3KNSxNdQXgar3VkiOAoAkr8QyrrntD/b5xjtn90/oDvJhjEn2OSaDP
EWSTSqCcNy78Bh3m8RC00sAwvVGFInKslr8Yh3KQnL5qwv5psOsiOJqehErTMsxcMP8NqquVzqAE
4vrHG+ZLmYT2LKI3hwlWqDyljUiEA7NJGySF3IvO4n4ESOjW3PuXnX9O+9sg3xg11qwzmvFiTTFL
FRoE99i1NDhYhyWzybt3TZu7wSgHAJ/YAKV9W7ASH/Nj+wbQqH171DVk9S12SjEW/whBtjiR5B9A
cE+Nn431OOndQoXPh248h2bXcdNV4tKcpplcZ/k8G/jJYf6R/x2DH24J5du5LY6t+QrB2ybiIU/Q
7TZJ6LAw+jJm/wNCMQX9uLaSSrp3n9ZwlASdlAwpqEbkr1D1o+auBitvLX2mfnac1W5TrXlKc3gX
iliaBcxj5rTZ5kXcvNNn562oH5IKhr64oAtvO32n4ik99W411RpVEbuBRlHHnJI4QEzwMtW+uLWk
3DRPmGUS98OgX35UZ+SBphPMJjOfLaf9ZWN99ca40ZwfEe0BzuQbep1j7aJDv+AGl3d+fhdmb9yK
0f6a7VSbh44wnQJK7Yq9MKDSpbgfRoA2HnGcZhqoSTOgJqbD76mUU2Ww+YL4z35d1gBeL2yemmux
YIhETQiBZt3wy9qAh50B7CzfDTOhGJeNQJZQw6A2OWe+ww69A1AjSWgz0Qisg40SseHRpqHdkztJ
b4mqyDvGtDhN8Y4iHYghJca19ewvH3+T6uOqsqAZRB65oIINO36YT2UDWsy3gpGTMESwBcx2/AE/
1TD97rncYuArGGeaLc+fFjxA3OJBbG7qw2pRsrrOyLomNuQCMATAiKNhVkj9bUxKKlKkiV8Cxd+o
v9o7YpjPqDuUERuvUkokd72cIyrDVg7Xu4d3mVhYVcnZLM/g+UmrWut1hjRu+7/fh4XrSTVSSDJT
8dr6QF3GjCp6T0ZHU7vVQWowq1JW2duYjtHeueZcnCYGlogivArI+qXhvyfVIvLR4Km9KfYtNDCP
3J1vpiTsSiYacRuZuI8Fbz9Zf2lzSRNIr37khQYjOrxbQpnzccuWkhaQeHszvJLiP//jRQdVjWgQ
MTFIadGxajnBEDVt3Nph7L9dSYUKZRHv+1qucRnMHTd0wL6zt2MW+cM1gltAm0AFUK+hEpGZuGNH
/VCA/wM/lPZYvNF560ZPXcCehwcvszrwHV42XYFgaOYQelmUKCHe47Fb8to2jiBW2G9j+v8FKJeF
Cej3PmAjUTq3jRZ6NXE31ssTBx3MQBPaW7Xvs6MOknwEPAOwVUG4CBEZnpywxjRBSv8fjWstIFa7
tAigwgBuvNSfupB6hHuraEXdZMxDxQOrhTUbINlrBjbP3IthElTv2pr17IfWplf4kDWRxFvRtZ+Q
/yxpwlZTnpMsrhoyyRp/ApZfdJRc7LG9eSVc/2ytJqt+9TX1G2IUuA7ohncvMONT5dol4JR6UX68
KRyg7DV/g+BzE8NI0Fx7kn/9NbL07rLq2Dn70wMrT0odKcFwioP7SkwU/jajawwjqVPmKtobzqjk
srxdeYCKCzOctZ6cCmL/kNxjhIOY4NPczrbTq2L/o8JGOhJWw4cntWOHp2nwZHUYNC0ZxfnSW7Nu
MZKpQvwSVs/wpNp1ZzCnQrc6tfsvxkBQaSPGIbSA8T7HgY8cFpRORhvCMZBvUsxkNumXuLn6+Bxl
vXoGvioW0BvQNl379sA2I+SPJJwlDY8UtX2WE0STJnFT+spY/M+OOvoBQgEGfp/ntTXIvImbVWfg
4OQff3nML1jJuVGqS/vPCxP5vaD8TSKj3XF/z2f3o9SlVPpRHmPXQC7kuFqnxzYsZLArokcf0HJ+
IQsJik74jsMDGoXgBHGfSUvOb7t+6go030THp/4/nn7Z+ClJeEdsC0X3lfX9U844mbAY1JGUu5Z3
f62lKdxwmWkNxcWiPrrp2s2NiHYwJ00TUaj6tH9F7qrCxMwZdMPQA++Eye5DBySoIzxZ7ZOSpfK/
483H/5ydx3K9GJYcOP5eb6W6Ue1Jh9Sjas2KILL9wR41rbyU5mfrn9c7ZWYcfG2cLNq+ldtGrilL
+7PvD12hUUppodY1u3NsFkntPNFrv6fYol+2/LpMwhX5f710wx9EjpCyB0Qwp52v72t1u8IQqZkt
T/6mRNLu+KD9n6C3mLghg556dNrwkyrnhQNXA3ymj+CFX+Oo0SJz2Q+hKwmUgyg+G1xE3i316Hi8
xAhW4vMDo4qsxHupUzRtA7eONBECsd59UM3iC3++EnU0GJGxOG7a6b7UnQbH7Z/PIWakQ6Ncx91j
V/rjNtjxXDXR2NYRQkiul+PQggBy4xvuK9Zh3ILuIFFYgf0fT++wp6rsbXTYdSmctitZoN2ul+3T
0F2N5dYPpT5gdI3QqV2c7G2KK4pibU1OXJbsPZsV6DI791cv2LglzIpbUcwc8eJaw6Lqa0KbHVm9
GVIeS99cSfkc7+LWHu9WnRdzOja9uefEzR8ibj7A7H1CRbvzUQUp0KyIeTjPoxW475pnQUc+QfbL
FsUKCKJh8VGMbA9BSOjCKGgZtHYsThXySNzhz1yKbs4tv/kltp8QaEpCWNj6FRm7XiAVJjiM5w+D
kS23aAUft++D+zKqOyvl6pijoXyRJzXmUZTAezsXdLqzI5PVOeU3/b7iUYw7j5H+yfZ4NeFnWTfo
XadHJNuvHFEWk+oL0e6Y3no1Obz3SYgMsUCiWqTh75yDTBGbTL1sjNSBhzzzXQ8RQEIQDOYZC/78
W+I0MBamc+6823dAUE8Lfy0wi2g4wXvmKids57ZBIx956y5CTLsng7I/rvC7VDF0VVO9FoXt/B0W
bX1LmEK9YNp43dkO8izrbwcF4krJ3utIPU7w3encZQOQ5fXdp4XH4t2/oFd3iczbL3HGwClNXvYd
QS5DzjqYGPVqnMrQFQBDMIPjAwIHmpBGv6LZPpH4kTDEwXl2YFu2/6re7v4wIx8IWpEuf+dn+weR
zeZSwxtmpg0Rw5AwxhdwWQQRYv4RhgxatulXt3TzhcD7J0l/iDT6t1qLEggI5Kkf+uNHCNQV8wt5
U8Zra2eRR/jXKFueF6yqOAWnkmyrHUXLmzj7Cho/BgQflB83iZa2tk1Pty1ZCwEyfwUVyfw/PEcv
imvlETYwVrBMlvEfelrnUbT8mlK2uJ6R2gzPFPrnjLyVL4o5m63isQ728meIriarenEnzG3Cx+9o
VdqjiZK9OQFwWgGe7lWxua+00KP4QLX9Y1R3zv864gZu9PG3GTGX5s7MFSGcLQdrgoeotJC1Y05r
R8J6DmQRiGXB1RUNBhtXgWFg13W0N+Rjqiuf3oIwT5Th7/wW8V2R1B/z1ojwQS2RDoTGOB8QejCO
ao7daUORLafBdeEFF9uVFnY9NoRaB7wlySvH/66HhdPSE/xdYbqbHOijTQduwthiw1cVZSORm+dR
DC5pcEevpNPEcNrzuagPJ0zGzJ6bQwX3vP1K8SKKXHyDBBfVbdwFIA6wLGjny4q/yKthUbzfUC9R
9xe6W6BnFq9NQZj3V+ow9Vk0qR6ZHeOuEgNSagkHA3tBP6qulLGEmX3sPKZ0vVQd8HfWysEb9Kvr
iK05exx8agiEmQxhX2ID82iqU7q5CU7sGGe49Ej4uQPbF/7Kk3RVV+koaKYMOpTjKBJeZVwigNTA
HUsOcRdU/6ZmHNd+vSFJbd5W/OkF5UMHB0D/GmYQ1BfislYfhqMQXvbhOvLXM6N6PTCf490tkGZ3
RiXR7XCMYIKZ9bySZ7Edhs/zIbEdiqo/kQj+MGYV8kuuf2OPGaBkiG46xHrTkflDWdcT+MAfxJjs
z9OI+P9YH5i+O+U5BX0IEXyLNB13JL/3QIZDcG8tYbWbYujaw/lqaccqIHr15jmn14jeeRuzGZ+g
Ni263tZC+EZ+iprR2FY96/cgBJn1E8FRLA67DOWhYbLSygSGgzWZR1JCIl10Ec+6h2+Jk8hE1X/c
cnfNX76Lzl/lxivH3GZVEVVgitd0/De2GsJVXdGXfI+zJBcMGWhLFO0kWr6E80nNle3kwBGzMB62
Mopv1nSqSawSFEXnSLUcGdr+U33Dmsu0FV1adRSMboqcV7y+MsYqSHzkN3vw14268WQgNq1MobaT
DJCS5Ot05TNgfsP9uebAEhJFna/hhdhPPFyt08+bJMQ7UvzvT1/jzxx0dUTCWevlBenC6mgH6RFp
7oBlRmKYRtj968x7mZ0M0UMT0C7zUSxsJj37jw339lu0VKrnCMSRyjoUwPWWtviWN8/9LW/h8hoK
eDhoi8/Ty6AhjD2hlx0niKjAaPmQFK0GoB5O4u49SPTfk8VOLpO2iykM5EvPSGlO/16/cHnHcC0E
YnJazcFZnUFAb9UJgxZw2ejFcO+isjz21JgGf/LUMFFzsE1JXjxfyTnbQYN+rj/Znvlle/JYeuY0
8x9pagxS4IaMlsgWH+FP7S0ELRC6/bBmRfJZjWLgrLCEICGLvCrhKCYB7YdG5CqPHxSWojQ2UCQS
AUMxH2yR9ixtd6gfPCj7wvC0lCx9v7YIe6YJvnFF6kzFJQC/i5Ob/dgRuC89+fddotqICmfwaQQl
yQjtSZ26UrgY9IXvM0d3QTSGNUbyDXUaepFjWXI/V1n7aKutSG8THDBedNzBMrweZDURLBfAhc2c
uBKbcOKSKIg9NHowWiy/8cJsJOzFI7J8auM00fFmKhRzr/G2DSpI3Nr/+0vhI2Nsw0WvPKnyAJvJ
Bsuq1TJ1BhXIpkegp6zyGonR0uPEAbKhePEH1hUvquRjBEgxV581vDCR55E/GHv+bzb3lpq6KNxQ
TUqkvYiVW1/IzkHh1FvXfpKMwhwjUEugvDt1iCBGk1b7BwoTFX/wego9MfRfOn+EzzzdyjGTzMWz
3OKq+WnVbfZZ6jatrUuOunFkFI9wpPQt/65YSM2mihVgOlQvyn05DkLViaEmYUJuxBgChUmay23V
FbjXj+XcxDu2vv3QAGBNMD1FACMCk2VPV6+kGrUZr84E+6iyzN2QtadOpbQolaFubCahbGqhZdh0
tlYRtF7Zk5BXfUpCNlVbK/Dj4Cu6qPZVzjfRO2HT6J4MNRNx7hcBm87m6VKU/M9tTVgvc0XzvsSU
0PD0cbGJtlY2qxlWCKjV2uy75CSJXhVnDg6YlZo4VdnxeIurhduHI/unxBHd0ZfdQXgB41yRYIY6
Zww/wnrW9zDHP3vWuLQLOFBa/bGlIl3CPzvrPXf6XvlPUF9p2YZ4G30zKZTDZBe7iIa2pk5DYlk6
fQrTYev4Tr2X2eWvkYMRaWRO90hFJmFkeV9yqEo9ft7aVpJwxR8SLC3jy9QXayKWU1FgmO3J6XoK
3Fkh8AWnL2J4sLVyK28etRs14XsckjjpzpyfzJwfTu/X0U3ZwTOyAUvCwGrvO+hmTaWZrg9WGnwb
nx994/6oFoeEUcy0IL4oFRHa4AakypNBp4Mgw5G3Np0o/szDZQLNY2UGQTSjEsqHOBoPyF83nFdf
p5PxLYMY5Pvih22xeKJc2cksywtT2jHQq4qjlPNa5eb4b8I4NLcS3X8+W3WLak+CoCKXn6jSb1kq
Dn2UoWW/gi0NREDHbIqR76kU40Hq8l0j7uteBKz2Friuq57XIAI5TF3GdnFjfWTORng0rCfLAVeD
kYmsonIrFjMokKeOKmQHu0kVPLQC6kWvBxGd4yBuiTtx9DuRyJi+uquwGLN+YdOnepAzVl7ME7eh
kcB7LhLIHkzrsR41C4tGsb3KiNqnluE4w26FY17AghH7dfy9WDyPBFFT22S839ltocdpTAQajXMn
hTaTGpKKX7eJL4ULjW+kzTW3G4Z22vL4Jhokc8BJjfUF32uCILsBMwNWN+YDY7B5gKhvTlSGSi/w
v2y93aN2HOlfzdBuiCcC+pm4TROxoGVFLlMPOqcFdqn2VHHUFBHDWkxyDXDr12ciPqiP62lzoaAA
1fJZ8jBn0/vxZyz+WK4a34YoqAhRA64ja0dcZxIXi8pqvkmilcqsfSmN+a1kO4BCErb0F+39hX6m
jn7c5cI4B40cmE5YacrBA3nRdHEe4lX9O1xSU52VelO5rKRgUUfUrAoNQWYRM35z9s/FT+5W0o1k
z0gX0LV05veh6uPNQlqgl46BZDjWIGIph6Y98m+kAW5DgFVOEuR/ib0MszRrBoxAhgi++DfGvFbN
DPbLVcMl3ya5bE241cSK9JYVKBqcVjmcd4+GCIsASw2NbFzJ7ACqhowD7Li24Q/vQseMkY1fOBRW
vyrDC4GGd8jOl+orx/GG2yW9zOoh+AHG700RWGqNAOXOSshAkw/tcOxlPLFQb+r43/mdlFjnGEg3
+pgtRqfHzB5eGeH+kaEwPoYjQQ4c/xzGBMd+4Tc3kIBbSsL/z1xJCHLbXS6Do6VWeV56GWppUkLA
g8XPFr7+lqbJCbL79oFfe71sM7s9Opc5cV0MSY1RAcmmNLXJUPvT9Ne2dtPbsXh8n5s69LcqOjB2
CXZcUJxYABdU9297xri+C+uMrzkU/sCI7hvHrjWqN9hyHnfmIWH3o4VrL45jIPFyvtI/Vaa6ze24
sM90StNu03DYMbRv7fMk8f28/3IAur7rmSXjDWAnM0ezexSLvNLRzevEGnUb6ly009P3RBmmJfaP
+MopUgPw89N88EWvq+SKjlM4YC+4avdm4l7YWWKRjfbKTxLFHvI6b7K/ZKEsiD7bv5UEU9kxD3Il
7JV13mpQWKXNzWQRhEf8ZV7XPTTZ3gOnF/rRPrYAZhH+JTI+fJI92xo5TMWptGok5zz0cOxpdEpV
y83CDiiCFBZDw0bAY+8jEb6SSz071zVd0IhyqFi2fZFP+Jt2LprrugbcgMQCqWPXoFWg3DcbOnrF
cRj6ZHGF0H5kknEuM6m2QKl0zfe890bz/+CwhVMHMQBBJYntLmf+LsVD6TpK9A71kRhAUbsvbMuS
8pMrE5F+V+KligSJp9VWRCupkSx1zytX2r1qJSADBw3Ym5mkRuTknlS0KSvMaQuPky8gQfLqLS2a
tF5GqyTwtmdSYtRUtUYdIp2ihPVZkEeZzkfUbXXJ9FFN62ZC+WOrynnMDpu6vB4sJa4yPzXczsIf
WAsuGkdeM7w9eS0XRjqHWSNTPcFoiLKMjQAHxGmdmTmGqJcx+avUVwb4Wl8DjzCqGjAkhbhQVs0h
ZNpb7qPO5WvbWVCXFCehQ3CB7PBnPXbE5DOMLWNyUhKbxn/uJX66wuj2NBGQN6Ox+w7DirIvbWjY
JNM/ioqpqOy/IBJRQ+DOPpikW+ywiEtWXvZyMmqAfcEHiLrqdvosK6AhL3E+A38lA6B8MROcvh1E
wWY918rwz190y7dESIqr9kdcpzhttkbR7nkNd+pinHNj/x5ntsSANZXNN0QpQ5PRVFDL8SWVjZaq
F0Fttg8HaqUBik9p0E71Jy97tk8N7iFlkMaeCiNaNab0TNmSxuECs/x8QyXP6zpppP7F5s7q/B/K
aE9Gjv97j0T7gummfAI6tAPF8gwnt07ZezKuaPhq2BUZyPJ0CNJq+J6uDq07gPIOw6rVO41LL3Zh
ZqvbjY8xKJe9nA+L4dChKNlIrZjCSyRGBlFnWggjMFjzE37gIIxSvosdSMzItiiJ2KvHVGZp8pqe
88lD3MCA1mE9ZSdeaH7CgFDNr5zTecUl7eBsH/cZv3OrzwViq1A5b0zR8SWmICVqSqMNWyMwcXzP
vqlV2BCWvCbLGUXlve8uCGSz3SBIUGL/woBK0z9FHWzIH+QSYNEcW3BzHXbfIHCb2dR3AngGVH3b
MdmvzwVuF3q38f+O8Nlspq5lBxbpchlj89E05974Jri0Kl7LmVC2ReGWin9aYi+Aggf3gSej2tgB
brtZCLpxDnTlWHH+Pak8jYySww1Ot6/uAIqXOfSlTsDl5kI9qveesLgVlF/QVGAOz6fXhJZrbHx/
JdamTyGnPMOgS4DeU2oVUZT1FPV7YO4ZQrS/2zT0Z9GkjR1GdeNqjEIxPdy7zfzsYwPpacPme6fw
Hc/k/D9EmhR+RUn+Xw5Rn3RDtF9G+nC7J04jx2SnUdpADR4MzAOviFL9B6IBcK6BI+ENnAWnMs5y
y1D3yotUKutquDS7A8ZyFl9h9mijytU4/GxwyXJ4z/yI9Ln3j9CT++FZC770ErEGJqWa+hgRhZiJ
uoME9ZrRJH3Vq0JJ7ujsYMDvaEYEzSRmbU0OmE6GsZ6HL/Dm3ySJhJiIivv/X0Ya/v8DEEqd7nVa
V91zF39m1N0TFguZtFpOcvswa4xJnngZ6k0Tt+a3v04w3HZb3LZDzVJWtbQhdQIJNaxbc/mjGuvf
zaoW0p2cCOy6g7d7wwHoEDL71tJrW6TX2DmXWYi9WRggoTPpoV/jNpPpiWmGQxnypneFwvYxwGPQ
91Cbmp+r4ewaBCVLh0wYrZP0A3gczuJTiv5WyuIan8UVwYYx4qWNBrvNUkb8HxyiFZsMtIIfWG9a
k3iZD0yqAN+i4dxhrZ+5CZynQ9QfxzZeOk0FKPRkfLFeD0m2+sOnD70qdfxpWwPqHsQk6CkYjZIg
bxPtbO0j4Rm8HtM3yH8d6Uzs/xgfyZm7fA2Q2O22NovW2r5HyBh5sSg9WJsBuScPXwzLIOLmwSV8
kLcxAzwY3ahqzQ+WOVpr4zHPh6qgKk/Th0l+/zSRKgGdjVFOu4F9FccD8SxLf/zJ0db7l5ASAqbh
BqQKXWuQU1ALOHXTR2+FysYgksRHP9p7QrdhZ7+AHRQgDpz49tAoUTzIkrsaB0keNhdrvOb/33Fm
3MCWUTzwSOnaOKBENIo//UMCVdiw4UggI+hOeN//VGd1yQNonsFPKgR4kGwc8BhvOGxMFxrrLm4a
gBiSPzp1n8zpCYAz698fegdhu6XwWl5aBJmWHMMXcg8kuVCEdHOsqPAEQE3pATnrpyRlXWFtQVYx
o3Z+3iTfq0e+5SzRXEWd5nZllbwrXZc+/wIdIjYfe0f/XQJqWVxprS0dJhh6Hm0uczQub+gkM/Z5
V6lcMYG+IoasAe3Yci/3piHpMbhE0TaXX0d9Bbhhb9CdbLM+ad1Pc7JHkJfEGQarRXbILt4LaLo0
8hlRD+Swov79aksEDKZyoj+r4FnAoqijT5dR9pKPcoxhGF5gJ+wucY05ewKvzWK3q3kBtvR2P63Q
M1d7z5ETm0cZO1B+prjWeq+/m3a/qlUJFeNnnsE8syR5Upak3nZEQlB1lfEmO+wArfnliCeEFPWI
iCntYHAoUm+nnhoz0p5LIYvbzG7DxVBhL301WBTCiBqrQno4wqehxk4tYNV7qh/wtRZz4SK4Xvc1
o/ofFuN/Z+Px2gRF7NcDR5eStCqvX3+CG3U5l4vWaJqQO1SQcRi/UxJPX8r1sLpQ/sutxk/HbyMA
fQ9hiAPckxzi7EBTioh8TC8++zOlJMMVdkRYIqIl/sfBRfWQ2rQVvsPewLCFnAwq4O3slA2gpd8r
KNiZoq9gy5n028KFPzlZydh+mgwK2Mz6gvs+k4oEDWTqrQzNfw7izyBNpJRJgiB57PSKYbfrd2Bm
LHvY2p+AwjWOujW7zD0fXHAsHgJqR2HCaLbbHVaVsDasjvxufRoX75XXhfiIvqaOy4gtGR6dam2v
YJ0OfUdVNw1UOuMm0JPr9fuyhTXCBbvoSpE2XuPz9IInAGUjlSJb+QH9QF0rpIbe0atvAqAiSQNY
MQ7XzwCcnQZdjbZbqkx6IuDrARDqbDIE4zd9mTJlE4knutuAGzOSHi1d1TOJA4/yyDig8v83Shzn
0Az9KvAETsL0Xps9D30ux0wWTIVpVZQ5tNN163Uv08uldRFP6Giu19eOA5vmJeGbPsTBjiKcjz+1
fvpkxX507MJu7yajoVjnOCvpDjl2i4TjbGh94PDj0O55mLTF2gUTLwZlQTdWccssBHMdCMTSOczQ
X9o/JvvTgEhMjaa/oxjfaUjJ1xCAbMExaQjUhMz0PI8jmaLERP6MvVjllw8roRWsRKr0RZZIJzIz
4g+QJLOXvCWU76JdcnzhhNWYdI2Qe+f00AM8KISy4gEKQQZYBINFbV7cE4nqVlL9qRRsfJsTzDWd
n3d/YSf2xYmFqf61gLkuwFPJhbQoLWvr+WAKrvkZ1RWQgKaaTbgPTTpyo2RHmIBW3HL4uonfCHV5
kNyqy+9+wRMx2p1TnDhU+2WeZZSPrv9f9eZqdZuZjVoacInxYxWPoXJ2glRpkL7QX4WD1r5LVj3d
5Ax43ty+jHcEA1xM2EkscxcxnM1JUDvgh3U0KR3ZEC3PTpwJG8EYjr6dJmyybApTa0pOdsbbo9pT
LluA/IqlwtX0Wv+LiA2VtF1bBZNUJAUJP4O2gYkGIyycHLN6pgyS58ZUZaAjyUN7OdkdhEOsoWoI
Yvzv+VOn+O++Phlh/BFP5i32YPWPcWWhlmFjV61jMhwW8LL3Mic5kl2Cmdpj76kl7UBUCOhnYm8r
/r7D4nZjYJ8Dsq/a0K1WQuJgCsNV39mgIRAiOBS+QOX7ajeigQVGo1owOmCdP3ltFPROnGsNmDul
MG9kcrziWnXa0L+3tXh+FH0fUOtlEO0QWeSajDo9shl9Q165ryWKgX0CH3UyC11VPdbWuvEIXDTt
MeYQd7Ns3l7JMTkgInQe/NqY3EQR+omNjRyiGoF483db5qawUs5hxme6Gk578Y0JR4aU8XwiCJ/N
I+iQodHFYu14QHJkoZyIP84DtDm2qs+NiDEOUvnDIrvtsZ26j97hXDjMBqhGzq7ZOfHJAaQTL+NE
GcOq5BN+MbGUchlVCX90IQ4rlAx2XnIoGGcM/K831LKC3VKxBhsCkONmNlCEL15IFx8OaC4sccRl
wkdQhoZNMBXGseTNzd8mt+B5A02rWQF2F87nHUCqLteRGR6imgyTd5EI8aqrd4C2/cdYSBRzgjuU
0LbDtprWqNtcEy5e/f/ADDrruzy6BuNI5nmWO1RyhUol5Sg0b34z0T17luYsE28+eSBzbLmMvAdP
wt9FZstlAhbRs/M1H+rkwrl3IsWZaovCkJ4CJYo8ZI2YfRzxR8yM/VAhCimtNxa8NIbcQDXL3gjr
/Upjz7kETC/bZB1UBbgVtCUU5L+H8+IlOgJ1MaVP9TiPp/Wr5RFsue4372LYqeasTHy8syNrR+L7
VphgO+JtjY0SV3F+EIatbAQfBXH6GwlOVeouNk/MzdP+iZHIuTVHRlgor5g52k0Bm4jzy/L5CA+K
4u6c4BeUMB9QxOC/+g4+HwVSk+914oSf0llRX9WLx0gqzUCepZoHaJ0zEGBQwSgKwvF/LOgwyt/P
u7MG2MAJLWrLEORhGT2J///VxkbWwPZfMu8MiodJ7Sa+fNg0G1ecKhcFHYhEp3KnBTWA5h7wXzmC
x73gPkynFhS5ULuerS6+3hkjMdmGaSRNJHsrZzSwZ4V2QqgeT8r0TDirI/ozF0N/GdTuWg8Q36X2
ddffaCKNe0y9/PLMbE3hbUdOJT/Qw8Bdg1s7CJdK8+7UpTaEuM8+HHeMbzpZZhxyKo1laZ9VkDx/
So4E5tiFHmQNACOUQTI4FuEacEuCnTlTLeHj1BzROLi24rRkBLl4o6evv/ALoba5F5bJ0pT+UXd0
HdhCXNQ5Tj1hpWj8xx/jBbIcYCJm5sKZgTJN1/tFomDkM8B1GorxatnvjRmHi2/1Fo8Nn12rVIRJ
hz54OXhUscT2ETzdQh19P+6A1KVxo+y9OCAl5kmM+U0GhzFqVUCQxpFveMD3wQ1L9MD6FbRR+Ipa
PGu5+CKjvr7AG6YxjReqXjY4DyFH7nDxopxFwcUEwlp1Y0LnMe0zlYrmGU65VyhxNq/2zMfhhks7
8F/BHeuqysZ8RHldXux7JGgi7usz4IVVD/4R0D4uqKW70wDUqzOD27qFRF3fo76uzMtgy4yBSKPK
HxhTY9YokYxqM4vdyqlOo9aFOr+3Z3w7A9zvYvBNyxx85rCzAmaL7f5F5A3hWq87R+EqZP7Gc/Pd
GpYE4OGaVVn5G7pD6deqqh+odlJVA6cd2QUSp2ZEBfCfbe41ZE9I28VXTr4n/VhR9tzxEQGbMmaQ
M5RQUNL+JEp8nTl9KuEPc8lyqm+8z1+7+2tWrVBffWcSqpg+qnm6QsueV/betnSW/NE6PH3PeF1O
tfXp9WOGgyR6sOOHbepz8Oj+jVxarct3Tx/KsK/CoBWKpDOPLyweixhpQ6iIYIgZfLxAGHVojZgN
BuNIr3QLvv9BAPwji3n6v03slGZqzrMUTJppFRwIQvyJDXeGbz3jQbqWJ0cb97WPpmqwkVMpyk7J
w7PC9BuQbdPT7DVWeUKCVlBIUhf/0YTbSGKVWM0ICpUnAdkwH9iVwSJ9rGm+BBb4EgaZcs0NjfZQ
cStCMQYFhw+YMqyO0vpua+L0Cip0QTdybUVYYv8kZ9edn728z7xRPK4yVywD+tmT/likdCHAT5gi
OStzHfmSXqHlXMn4FJxlC0QD71rFABTMxXA4b4+qOu/zgtFCz+A1/q00OnpZbl8FjDPTkY+05N8n
tbAAO038PXYcU6VJVm3A2VDtiASQjEn77ahihTCh8++l8DfHcMta0QLZuNF8h0UWsavYzuL2rM1D
ElV0eErMHayAnS8v5KYDAvWWQf96tmHOH/2Ado0QgeZ4qELk6Lo+IKS5bpIBtIvV6PaJDsACoWOU
NLzfGnnA4pLdyCVKboGJ9lIhMQggk7pyLUIA5PUfCWWofBXnDkcvyYcwORLDMxDBU3yxpLq8qZlU
q8AsQf4pNODaWmjsdevhKmcAw5RTr0dqhXf9l5glI8DezxH8Y4DPVwrdzMOQI1jwup9bICiU6KLi
uwAo2uFBH3CuY7+c2HPO3oK5px9n3hth9TiV8gORI+eneAFlc7GAoWmPWxXnnOph27owN/4vlmnd
yNAgykt/icN7tP83qXguHFsUM5hQfX+QHfSWDiEXV45ZBkfCi0baux2K9AXYhohRZz9FqK86/P5n
MCyfNBTQYDIex1MpuaRLNL7WHdyPjACmm7hviZHyWRDHGwxXMZLUeHX3t8L18hbmVAJvkkW8mgJ2
Vjc9GaGwXjeSb7cAHDd8YaYdcuXGQEs5ITWUXVR2gP9pYC1hs1pUNHIE9phkX8RVqhdgFcpyd+sg
2iqGnhMN5YZgw+d/oEzpiWHjHkjSYKK8A29UP46Ob8KZSHPuTHne0RQbOWQ6HaqvLBSJ5Cufp+Ww
jw8y2qgdLAtniOpJ6FO2a3nBwwrYTpIFtiS4zntCHCreBYlg53PqL9Sh5lG37gGiL4qpkUK8o0l+
SjZLpeMKFDDiot1Oas5i0DV5nkU48AkUdY2QJz7Ge63tZp189tFk9od8TqB5wS8IZG5CaPXQREZz
nmCk3x5wl/BaJw9xKQS8bj1rOvVJCMIc5WHrHrMwbveAqAWnFUG6P9CzPe8d+mBtaqLn5xTEAgOV
pPcDYS4hPNv7I1RUYLA/q9mCTXlIHSdKHZ3HJSOtwei8mZCufX86F3NOx7C5WMsvf0tOV2jEu1hE
9/k567aS1LsVA5vB0wSHz4n5m5C3kPs8XFNu6HyV/2ycRLioVUCvotnPJoL0vP0rnVhgkljh8YuV
Xisq3fMATZuV3hr1q2F8Cp0j/AsWdxK4zPugwxMOhmBRELu8YDe3p76YtsbAR5MQhZYYzze8082/
bGQINkfg1d1gct/tJ5BH2PqMux9jN7YNV3u0b/vXDkH2huFkG2l+IQTr0lS3443cHzwdtpSSSekt
/NCgrnkrqhZcbqM5PnxHfu+ot+nNLvRtIaY3VCTMILWtXJS9BugLfaBj6kJCMXA2r+o79jYSfoox
eTgmLIn7zdKFvSWP40mTRxbpjqqIBBdmNdEHlPtAiZOFLX3sRCNkTUvHqT/0K3DFNsOCspvI4VFI
wjCMv+Buxe9UYXYfCtnD9MIoSkRYmMt379W9ibxN49/0QIpY1YCn6cGJ3sI+zOjvvGb8Fal8qAi/
puEtM5xrn1uOXQBYU0/fmdbl3SfIx22DphumqRxIYzd2ubS28fRsOf6+poDFbAEku0CatLUXBWMT
KH9vQjdUIhnn+oSdC+fvHuctlfFuEYhZ99UkJcU6Ky1B+yzZ3IP/CKFluq/4Bh2i7JAespJHbCKP
DnPO4bbvn6iqxyuB3P9x8d/g4WQIq8D3fw53g9FjOvIrspeAAyijLbdV1y+KrC5qeaUilP5AJGSI
IgdXcoJ+XdJTu+De8DgM1Ui8TShF+fJI5G0NFmZHduAvHnbB3tb0qh5yuyCaWGjNnD3vhM5boOYb
5swCYz+R988BcQQ4Pra7laPBmwaCTfIzNQ7zZeOawvx3J1UZloRTqrTfxJSFeNR92gucEynr7sNX
skZIPalupug7qZclG8RJwwcSxGm9PUSg2pw/zMI+TEeeTs4rGjQi4Hs4oepnKwNY6FAwj8tdi0f1
CaA4YV4HPLNCcxNDL6gxp0Ggv7SdTo0O2RzZwb4RHgFLPOHJopHEDRi30H6SYe9mSC99zYbBCYdz
9RH3GAfPmPjAfCEzSWcTy+I+YodbSsFRsbPWwwveK4CVYU86yYiQ+ujxWumuUh+8rmNdD0CqdrIS
6v5CRwZd7e6/XfLq5k7SgLTVZNcRiDeBWaTUZGKG04TVdb8KvfysKtedzkBQzrYcWinkndXhpsrI
PPwI9papVs+1YVjuycNjyuSjng5S1q88YbZyAS2VIHQsbEDm6P6qHl1ySTxGsDD4/zhC9fQUcLV6
BZSaDItYgDckbQ6x8G7MHRoBRKb7jk4jUbuSerYQ7qu8WO9nP+BPFDFk9Ypx4nrzWEMSIfG4EBtH
RTwGabE3awhjnG7efiuAXTlURw4+UQ6Jpr9YecgXXZP0ffK+/4/2qxvbD/dzsxa9pka/fAr4NdU4
FthFkt47F8mnWIYDkFZkf5e7q0mONmuVZ6pyl5LZ7KJpW1hKFxDhWdJYkn5ngZ5lCQYbPpznTB4J
8JT+jVuOQHDyTuVinnU5vOwvFmHf18i6R8bYxALDYWae5vNWoAdz3zd/hnD82tH2k3Cls9jtu9rd
fMj8aIN2bPackxUOKwbumuXGpcbnxw6atVyvhXVqRepNC/UoFvSRZLGBZtnO/peYjuT8AyBqq4Jo
wafE3t+DPaZt05RZM0XtJ2u1ioPHkxHXA6JA3FwWqqy+jCB8X5eKj8aEBZd2ElOb5v1dvIfGxlHk
XhgBr7C9fehiDOHG4sCbs9STf9S9c9EZB+N0WiMIhcdB/CT/m0qImqAoKyRvv5Krc4hwUiy0sVPo
MUmVCpoeY/Sc289oky9zG+tXMagfseo0HI9NaCEncMKLOTUoPzpBKkWizDFtGjWk1fVCVHyVauG5
vKOCKlmpbRPbitfQeWwPQcsZHdOr65o8AKDxtsKNQQdMqd3p6r9S1P3pygg8xePI0tU5/pt2EdqD
gmGQQ9KTfEz/3kzwYWalqT9qCHVtT0bYQFrr8oUr1fxOKGG5XAkrJIi1hiIUkbeFj5DZtb728vut
wfHHWR5cEaN1EzVIj28hsFRcjCWkk5B1QKy06kopbdSz9Ud4BN8jt3VprywjUI2q+A708JEmo7O/
1JriD/MeuuIw/PUMhq8S3gyh4nkA2EuKT4U3G5UkInhFoECNhn9YCV4WKs/bcE5DoxGbtQS1GgQQ
NS8anGRdw2tz25ZghfB9q2BPz37dx2Adve67+W04Gcswn1HkoPV6pLgKcsvGoefMmIK87+bvNV8u
NOeeUr7o/rAareEErp1ZhfowbkXIuf3M0dPdIEpNheCdbvP6hpwcDNtBCZF+EG20KYyUNrkmjvJ7
8xBm4gjOymK8fHDwftmdZ/NVPZiwQWxOdFru7FV2tKq6NX2mibgidLmBbl/rlzSPT4ZSgGQyvYvu
xgo6o7jzMdWdbXbnBMJQz+gykCdjwn7z+FF4EUPFedPZYm7Ef74sDipuZVq/FzcvNhPKSBiw3WLF
1qR748uax8UJjaOZpZd0zrORC42NaSskiFPZOBG6B/aZC02C1oBy+S4m39nIxEJzBwakNKg5NOhA
nyHHTedim63Mqs+6bVg4sVzol9dPz9suEMoppqpmmXVGnSx61jX6JTp59YvtCogNogy/ICWqTbvr
O2QV/6Vq3ONnQrgyFApaZvNxejsh9DioSGbRGhelD+Dg8z4pGRUWTHY9FmsziudkEiuSPdSPN93U
Tq8Oi1U/AQXg3mshX7k++ApNy3qH9NAPvXq4XIocNW4+xir7A0Sy1xpJFEV3bIUN+FrWR1Cl8eUc
6K9LKG3FhEmvRNzT0dpWgoxGoECimgQT5vYmCGENF2hOSm+CkAAJWbeyHICiWSzmd6Estve8FAi2
6949g10iKxWGseug9YXF/roqmKIxpJim5jVFG0++i50sYuJcVaFiLXMvpQtMrk+Vg1WW5yB7N6mD
Z+DQcCfCl5vcYREcw1dmBU7CYyzHxoS3GPFvImNoDkJ3x4DSVJwQcDSQuo1vCCVChQkGOjKsm9eJ
j4kfS6SkiIT3YTYC1PTo5McguKJzgw9vqqZKF54q4XKpBAfsxPrNfGvjGzssQU7kzyQUo6rF78yx
y1QL2FtJV1QrK/Ad4G7hTFMVXzvoTEzYIUNp0NUiHAR8QLAb6IoZjKuZNSEDpLtzktlb87gSNHF/
h4LkL0lGNPfy0wJekGL33G+t7if4wmog6hgEzHRBjrWWuXRgjNHQKk627itsO4L3wxlDMeRX72IE
tKo4UqaKFuXK7Xmxv20/TAF2bsjPmoWTJZ86REk5Wz+MK7f2XuNNwhysMIjj3d9eFcw+KdilRRTb
e+t7qIx6BX/pRG8HE++z1x+j5hjs3IsG1SH50hEDFhKTnweNVBBs159GY2Q/NtLAEPKSXSy+ba0u
70cykESVbUhq5rk2yRF48mu9V+Fzy7y9nSOJz4Hv+IsqKy8UQlIQPr2DqSbmlw38n3ByhDS1cVxi
Mg+K5sfN690L1po2kjLrKGVN5M0gLo7wV5VxTCMiB1rEe/vaV6rYZNnr3L7apaCec2Ct4wE2fX8K
KwNN59LK0Pp3JAKCxZxL5lL3vIlm5WaT2511bbJp/cNb7JZuSfwpxBbkhmzEKBNTyLGPTzrTttnI
VSlJM9N4ljvh8+vFF0cyEWU1DxpkcPhtjEyS+MPr7LsTa3a0+ka8Ost2skYFpEF3weiVS/unYf44
Gn7pcGTKCpz14sykx+a06S1Ucv8+bj6s01+aEZmTO1ka5K8dJkwN+wn078yEwkiRnVBBRcJqmo2V
fyqUMzi+y6tFDX/DTedavTEsMrKrBtxJIOkZREw8x5Tqm1lAKocZH5J4qQe6CFsmZe0U9fkARLKE
6L7iANNEAZ1inroIN5IxN5jqlDPL4+HIa5rCdiDsenuny5enJtY55Pop5ilrC1nUsZSAJk+jPJCK
f6lByKc9tuLbLjJe0qOyPIAEbF4k3uUAOEKkZ5qYK3aCJWy251R5TtJkEBHhZD74ZOvKKZoTYIjR
9Wa0RgzgeOo8LnoOnygLsuGNWmaFKWE04hHe4y4RZt13xlU0Pd6vgcO4CKYp/kI1wdaua27GITO6
bJD3UMWj8gyCwnya+QnXccKbg5C71US+YTtQ3wIpHcOvrQ/3j2+UXCFICu7D1c2XDbqGOi/4nv1Q
Xl6u+T1nRaAWxCr7bJUAg2NgvXmdHFqULA7/RL2S8c1Rk4soO1NDG4mU76tN7sob1+YCO2UWN53E
6TZtMJ9bJu438RN7zsPqbc8hJ7l9GuBlUyjXKBLZbat6xaGxIFJsUp1uF99GhgU1poaXxSXzLMN3
f9Dw4u71e6l4WEGmSA8T9ScW/ybCfEL+F/KnT/ym8Pdw0fyKxQY5gWGrKVNgZLb5TPkfuTMVV4X7
pjMl+u7T3R/cHCYZcBE+zJvFmmkChwOhTwzrNuU3tfp5Z6W3U9j9gwVwun3j3BKfnSLiE4j7MDud
lTM+iaAyMKPV1MvmQqoiRGgVlaDS+m6FCyZDpVzX5+liRxsXXHUeXqsME6AS32uSqrpGidiWqj3H
bMqnXm87LcrvVXu4badGig/5SccF7nlNgfeBfWV2dorh2YVX5WNwJ4ZnZ87uinBumcOFwreZEZd6
uS2pXW/qZOYIRTdiO3qIO9P9/ogxHTNIE6RhFWhzNaW4i5ME5AOEcxsXwfgv/5gNZbBs820NWD/d
KD6tlbNTNhYhG8akPXI4UsxH9d2bWOoDhSIlNOlpDyU14VRDgLD0k/E8zxVosK7DpABK0iJrmGDt
MTqRpnFt5WgnRZZfXuRLQg0sFM9R6BZPi1DgTzwmU9sXppdA2xXskfbQ5A0RZieD8+Xn48wUmiZe
0Ne+YzfLTuVSbvwCyBqmxmdsn/yXuu14MXdYTEiXg/hC4azG0eggfc5lunVHWZcLx38T5fbmHFGW
5nVDE+5r+TeF4WqZt7x5bezcdxbHFsgvK+YRmGDwyP4EFHJIdT6vwx/IxtTevwUCNuK2ZfZZ9cPo
1AqKY6nF5SQU3wRfm3RbKKsnkMGiLqcKxFqeo2iVBmhmCSeMFyduSPjyZQHCwqaInDEUMnsb2Fmy
Lyp1e/KwH3C7CD1P9112qkSJalF2SinePRIanYtwNs9OM/mESTLoibae21yloEGTz3v5yFBB5On5
Q2PiaKgQTu9T+LFIUheDDe1TxVDAhXQ32/8R2NhjYL1YijRz4GgWFjknvaewxG8vHXvPUsGszvVS
E7CJzmuusktaFPyDU4JS3fjsNl3XqLXpAtMpOxDaMODkVJzmmUXO75N9yobR7ZMa+NmacMNHHYNP
T6MK+amKYOn3tI01WhNRmfX9idMfzCldqRyB6uRpvoW/n56TTR9swqJRPDg9NjBQkWDxcKNQ815o
NaG7dHMbnIXIdfy+YAz2iKN6m8kjzys0dGCJ0cV8XXp8O/4Xpl6lHbFPIFYw7ySDCQcYhiaH6BVb
PPqDuOetM38woq+JyLncNvO1zjvIown8cIDGTBViPIuWyEaIq2lpEsCwkuhx1P2xtNbkar3nOoUW
VmAxWh93e8kkPqDNiV3Z77UI9G6OkQkS3ARfLZbbZKfWVCctXC4OnNO1NBHekUdPRxvqBw1tk6wk
E3lMzCcr7PpNn4CbEMNYlYKg5u46FrZs5vwCuwdjbGm6MUNDHpydx7lnb0rvfdHmjehUfpbDiteX
Gfx8PRUo6iVFddn8WBjyHY6DDRAWxXcqH/dLhTaXbNJUjSvqb59i1LgIW562jIQVINMBFAM/1kPR
XZdTEbq3FSKNHKeVOBbQHuKL2Z6MhlL9kR68qnaaH7cegvznMQT/Qok1ZmAx4k5/ICE0R/GN9u9V
CjHbJRZLUWGNwNxgGFuRzEWjzD+eIcBsg19nFh70Br1qEn4sHZcKaijOAGMZU83QeynlIZXMOpEO
L45gMXig6JZ09xmteeyM+xh5aHSl9jg1u6Q7iB68Oa2T1Mcvlpk1S50cQZXwzfBjuXC5tQnatGET
hAZLwKFf1oocUsJXqNPMp2XBDYDZi/XGhqsdfY5N4qNxXYuT3CUQIx925h0aRcLbzIqlqXL5pJh/
BTE8X17bskO385R57z9P09y6yprYEavptOkWohPXWI65JhbDnQpo7VcaMiSMk+Q5iozBJZw7mZ37
n9GsmdHUnjjDUnGwYB9JDoLL3vT4r86AgzXfwTPgenxiToj0osbpUbDc3SAcYQwXNoaF26lXNfaR
H+JBah3h+OQKdKRGlEzcd2csZDbS1PwnYUFof6vl/xmaN5TWpFAOrUNnYnWSeOA/FotAq0XyrASl
DfHAP4zvMrDP743j10aIfB4LQA9UcWVa29e4hx900U8u6PLwC0KBwFE8j23TaomwhR5Zpb6fTHwN
GWySIUzAHwdLzf12It+SUMAC/Y8sQ73QFy2s4jd3rn2BRyqz/4vN4HPEN8mW0f1Sxh9+YoJolZXw
TcyKcPYILGFdqZktNfX5Nk53HMd2TP/GA77otBsat3bVJ55nVrP8Eb3Nsb1iKPiJypxcNQHid3cP
+S7wZuH5wvuugz54JJGfpMHewOvqIj7bRDaO04GNV9KLDG8sMrbe1P4RWNjbag+hKX828G/xSpaf
HM34M67l9WpOd+4LKPJSt7wBGX1RS+X2jJ21U7G+ZGiMvKq06WOsBMtH0a38guh+omBg0oseKvWX
kXPTi6HZKut3AzVPQUoLWgvP0WxQd64FveHn4XuHgvTaz7hg/YCX16/CbfTv/gSM5yZtuGSys3eB
nGT67dzNYFscl55yx4WiV6iaOePmVMSL+f+hqENE2DePEv0KIOhGGvfF2FkwPsETNFezAMh+y1Yr
/WJHX55ONU3JgQiPE0dQoVO1Pdyw9CTsnQTPuoSgsKHI+ooY27e8eC9zqAehAph69GWjqC6q6d+1
Bd6Y6+2fLaQg8WUd5VHW3aaGxklK69/8AQqDO42SHiLgRJtM99VGo7CWKmb7fTnxxPZtMg9+LvHq
cklUlzHPBghs+GWdx6MLpmGJRt0xYLSivsyk59bH0kzYhCVSII7tKhu8RnSq55wLMZ0ZYNpABGa7
yqQeA4QqOesc7V8gLf6HrUA/xzzMnJAO5cXOglxy8SrvKGNtfhM9fnpB4xT0pn5LaT8u85j4tvbB
Sed+qGTvyiv+kdoS/4FRm7EnnGUO2KptA9VORDmF6X8hJa3SvaJ1l4Jhc5A2fHVPuAzZ66aL1No0
nj/TbYDVYPzUEJ+GkFP2Rtr0/BfDmU1bR7G1EjU7wvygyN7VfL3p7reI709WtJtR48DIidTXCQAB
ltBZSOvdQFU/kPMFaYKWm1+/5Zmka87rTV/O9l1k8XBI4OgDvcBxPF7bQ37w8GvNvEDt+DStQP7F
1Z9cEK2iP/0Gkhv5x47ttyvsQQZqVLV23hzUcRAFvrrBgVRV3j/k3GfnpfSirGSTSvGi4dF19yXS
x32vbX5VNxHF3NQVgq/fRkKTefMYCwqwSgI0XEA0aGA7W/kCOXpLIL/8MTsuv+loDsAL9SFt9PLZ
hMqjLSrTDGKTl1D54ymQ8IXBBBy23Pq8VXAez0fFba09SNj76jINxvLo3wEQHXNvjjEtSm01IL1Z
7ifjbXiPcYmZINYxMul1bpdqRhdy8UpfRlcJqYJ4YoWQOE0juidmxuudz4kXU9UluKJbfSG8aBkl
gzn2KPgNtkvJRU965yh4vRUBn4FIboiAk3w1LleYWZUlqk1yLKjn5EzaYxSrVzCff+EneuB3vYDt
tCJnfq1fY7IuNRKnXy8U8yhOjhbiJZTGGPLZ5Y1oSidrV+DHbBLROgb+Po9HkPeUh8hB46mBoAcn
q2TDD23dwrSTelrp9zRywnMGPFRvZWQISvAU/cVVpGq80DDEw7qzhT5HmiaYAeAfDnecMmefJHYZ
Ch6L5+WCRYvu63EALbdboQ2EGQwSF9zMXCjpwmEUCawZX8WH6+Qy7rmkq/+6JGwO6/LTIxkKhZ88
SqTYZxjxtRqKmjqI6/Ec6Hnrv07SV0E/3fI/xColYxcp4P3/vo6wz5VZ2VeWchicb2o2bPg2JFZC
NpRTxfrBdPXckelrfnlLHzZ10Ne4IKGrGHW+IGi//vjD9QnngO3BK+BP9d2DJXdTPWmupwVbIpBh
pgBcR0G4wCYeD/RkTsIXKsYi+hzNolcgG6L+v6BVz0vRSV0brfATCnkWjfJX9wUP1drr/nL1L+Xm
hlzuLnlW6ZeLH1ld29o9D4VnXxIWyMV0tDo8n3CnuKN38EBSc0Bszg0+3dksXnPCxA0OesfnngC7
tKw9GKAe9ukyCG8rI+mtCYtl7sQybe7Ifz+O0Gegr5ifK78JGUkKHV1haIZvl9iYbzPUR68UveXY
iI1N+zcQmZ4EAqTV1pNYrYDjDmFuays4+wIbwIDiYRgxlMlUh3wFbXIorIg7OIX9A1pNX/GudDvh
URERllYZ0Wh0rY3mwCGmo248D3DsmcF3Dz07D4YRC3BHjyPmc8yrLmrBvAPd18CgqwDpKcHtcm/R
jJQSLRtIWvO1OfcHdr8zV7T+edNEST45pw7+SVD0MUXUsCVcwbYuMi0X06EGTs77JSboRuxFkiZ3
f6AfVv43TTlBaKJ27BlguXQ7IJlHcB9AOrKrplsDJ71bQCV6Kicif0g1F5GO4zJ2zVhk2ewFm4E1
y1jmGoj1wHSkXeywTOcxUveUPFJefCc96gvci0Oh0kQACv9P94mRLkIgGK+5AUfNzq7Cp0fX7CFF
xb/gxEBisdLSsIcaFLCa6FufRYrtGW3q6rB8Smj/qrh6wEibrecGrfa7ardLU3TxyUE5taIXqbiU
wRfJtjjPCEWiYDK7ZIfBYR5zBVX0Q0Xzw3xtDq7nRsuWZo5AwMyv/8kEJSupVl8RaVVkYFoizF3S
zc+50oJnej9CbNyvfMUu/TEEnPJi7U1PCQ4Hx8PD90Lo0Ha+K+0ZCh08n0LPnKky/wnOQqUTkVH7
uNiLu8pLhuTrD5WXr7v7aI2fUZZTkMsYcac6/pbuWXQvCpxx6uu6ps/71IT8gfachdwGuuRrNl2a
Jw/rGMyYQ7CURdEbJ5lBmbJZ3v3RK39Ys+DpEKl25K3mb18kB8QEiKammnKimdDF7Gzi9vKCpzER
Jbn6uBafKWQNWDCYiCwCqgSCRyn8uv/FG0uTSGLQW53Lmzz3YX/KuevX5xcJSJm2DDEL0OeXXKoo
Npm8wXABkcNVD7bFBa9s0A3cx+egECVXIMoi2dGdeLEcsSCcWOKc7lt0Zvl+5dlA7RdYwJRrkK9+
GmxGSccBjqIrbHeWByfBmudfpZMa0LO/cZA8fzOQ/hhANdvGM/zJNsydYdvuV81zxILr41oE73xo
s29cbHjYXy/ItYp9IusxsDpjkm9C9eiMGNigKEvD8JrsUJ2ZabVaiC4O6M5USs5LLitisCpyxySW
d/iBbAOvno2v+WF2Unhw1e/LU1wIDqPq9HaeUrh289NtF3KjycK67zwVPnWAF9e73UjwowpWn0v4
ufyUmfif92nGfNgIaxrW8g06/gErjfh2Tc/5ZXlCeHvb6iotIUmWARWyPRpW4EWOXzlw0XnCOVq7
Qd9Y9wpmTsevIuPYbvu7BVzr/92A7fkB48N526QoWdqMEnS2K8CRS02BGu5EdlXJ2cmPBWx5J/7t
Te1+v1gmmzQ2JXkWdudRALOnWHQXLUYdo775JQxHcl0gQJLJNjp+u2zIxCo5m+6Metjtnfc90UU5
PtEau5WV9aG/ChJ+H4mMo5IbP5ZzVU89ky5j381GzKERNQ1699kVNTZyVszko0jvZPdcmtLVxtWr
Od5DNfFcGGOMaZY55KDkHqGmDzjrlKqBbCok8/IYG0cjZT23ICx4YAIgIiPqX9mRw5QSFX8bh1SP
SYLPlvZJAEox4qapnQvkqMd8OVssQ/stGiqWjX1zjwxzcUUnCBCo7GXH/hxCtP8DNolWKxtCvRFF
OO+/EzVOxl1AbuiJgUk2BDGrflYS7o7+hzK+hPatooch0aCLyqWEhfZebeQCryAAK2GXLlqgs721
L3VBosnRPs17gLwTbc9uhqad7gc29UjwPe7wlDNii7q2ft6Y/ui1zr5wNkcfcSJTAFkUOkFJcQxJ
xz4BLGYE9aZIXT4O9Yon5xEpMYkR2z+H/l/YNgjX3DAI7hcP6XIh6sSJU8JsFDRyOvcG3qB5BYKg
QVYu8frHs2/VvqG7ozWv6Jdumzkc98wiy5uFRfFSpsStncWdp2hOb6cmvX4iS7YLtT+oqjIv1iSB
kxlV1TSPP2x1FNgIK/eYhAn6+c4u+2sZ/G2J30nxLmVucfOzdJG7UxRnFFOEq/OZlQIYanJpOtzb
0E/OWM2lJ+TrINRb9fMeDP8LSm6GTT5GVGco9jqU7wWEOV0amDDPaJXUyQX+Nvei4d/wWHRqjGwA
SQj0P78OgBuGXmpd//BfX7zcFGDva3Z2LL0c/OLIHPvn+WdcawQARUfXv9cihUeGgHFlSE8fbAdL
QDXp6BPUyJFSEMxwv37QbEQU6KrPOp1+1sPEguHWUZLbJ4Z9hnGqXXxhtHb70raeokzgrR3fUusv
giIKyf1tXrt7WtRFIJHCD9oAawq+Q58MYy0FO8bantw2pOBE6k04vVScH8C+miVsowIMYqGN9XyM
HzCZ68Ti5OEJ9eL79Z35AWLG/nfWwXka9p8Z0xFU+qDOUMlm+sqiXe6utlvCuCIh/9mnkViQyGsH
06qTIxGCkWzHil4uBorojmx6/4kIKy2SHUhowrhT88kKIbYygsj9djszKFYj7DCd3YuMYe8rg7vN
A0le4wq6/ICO7F4DRIiEJC6mv/jki43pUZhe6QBXJIg4JYBpiGDSsBRr5PSbRSOWnntzt3L62AtH
E+zRcyIJu2EwO4h68vvZqmmxCsMos6MnZp7eAy1ebsBpWX30+lnHqNK+yY1kK9lHV9BSvjOFOE8q
g10mVzzx3zdUeO31pQ+EQ9A0dgvJPXJTz6vLlW1+z4v5/AOraH/GxLTHE/Oj7xhdmzlaYI6J8dAV
y8NzqKkmZwI8gS9KRM580D+2LlUxQSy/zPcjg4SjXzzjE4fZS16s3lMC6NzjZ5GFWRZCfo9Mlcmi
8wb4Rv/ep6xEXmEmHSl4jvx8nJf+QkwYcfqvqmDnq67yFhdyZLYbJQPqR/IL5J5gFzKhAgslavzB
AihIsphv7B8MeVGk3CA+bmJzlXufExPAHjWJRS/6EavfLXwx50rDnPgjTonwG8K8IbSwjINDixFU
T+W/ldEOqrij3cyZsIVCOZ23F4HjHrz7b2UolcjH12ir7F7wN1a+/CUI6SWKZwuiiFc/qdj21Dry
gR4LLikKv+RUnZzAkdm8sAWf1l7IV4GBVMr0kHrERlpnNDU4ZJX6Ud5XZHPnbVOied5vBO0+QTyi
NDgBCkk5+vlCgieL1F+NHhgCc7CIZphY9n1/XwRnzmT6RG2Jk9H0yszHeHDtHrPsrRD/9lFO5LHb
j5Y/g4YsqyBhRc3o/llUH8/WbsXCy0qVvl2D7FPvlo3DPb59R+OdV38/vM/bXVdulgXVU44INpfa
jQiGzwVOBKfxbz4KgALh6amPv748LQweV3VWoXpGuOzKBRBBpx+Pz3qN45CANChzX9RA8RqO1yJL
FuLoL9fP9EytpP7cClhIXXC6V338XIiRt2I85pi8sQGqvq2rPffnSvDlRjA3deWxnpVwiYfz+z1x
ACgPVCtutH9gFxYlHZoKpFT1S1DPTagG1KaWMO9BEeJXoYQWNMABccVn9+XxD20/aPgHrSUr3QB+
Jbnv1aO3gGmHDvRt7WRLXlwBOaHSlthEmzAokvUaziZZVPI4CxirB5w/mbyNO0WzqK5eR2qoyMx5
P21c4B75a46AnSEckfFciV2KUUpb6vQ1dAWhvOgKPCtoi2zIAvYrwPQU6vwa+lVAlfO+Xe137XKZ
eWNPOI0bE93drqPkX4ioOla4P/axsN6gjZkO5WoLq1eeu4MP3KARWuYxPsRv0YPbNamlXHnQy8vl
Sgyv3XyuC29ev45f29PQGHM20LY4wkKSjN40i24NTyfwekYXVq/3goo1vAASofCL1i+bqgEiBvFt
6ZEf56SfqP6nprHAqFzWYxg7OZ5o/H71sNPS+IsEM5vbMLmhqJJfCwgj0z/Qb3TlmmGnZDaXu7s2
sKLQHGk9Fyv/+PEiMDvkhX/5he7bKE+/epMmZyI7tlOzUPoz2dOvRZV2kXUTwd4vZ0QT2kYStF5a
4eoyWZ7nkf0Z1iU5ypcqNXqmnAB8j81ob8d24LL+s19ZcOiYmopCxGFDkpEOKJ84qAv88BrEvC6S
wYshVMqteSCdk85dduK2Y64pPWD1XPwE0qrqlqpcNSK2NpU/r4MC9B9d3E87wZ4KnVN3jQIlehSn
JU/zyUdR3+9gvgyBBFpJuwxuPCCcNuGtW3UI8OaIX1/T+C2eSCGXtv8I+OGbUeUf9KGBL/xCNSg6
6wcGnWsf5XyfcRxns6S334KVY8KQ8tFE6SJ81hj+6VjN4W2PCXvN3SmVRna//8XjhxyRSDZrOr9S
wv1QWXvNDIxoojEp5QNQcxt0b74Y81z4rwY1t8urJCD33X/AzhoWyYTyNxd1K40cgYAXwCg7UTUq
En+Rf2566RWIAfe/kNaESG13SgTmCIQMJ/DdYZYHiwQRuPsA1IvMMng/r9BbUigLrHOYy+Ws9JVJ
OMWA1SvLMAd0LDE37eHpwk5tzIQCxUDc8htMeSwIAVpLSt2sgXGNPQ4hLZigIzxiZEcoC0e9bBtz
7Q8i4EMVD/k1C2VEUCParINbqDSl716Upg6ek5TLXtrigEuk2xe0GR7h1KD1ayf+jXetz3LgRh33
FsT8H/AP2nZq1Cs1xcFD5/nGCSXZzpfNK4XdaWPrGwSvjmdTdqz55OUNfzKSUUAwtbWrl1tXh0Wd
Dg7DXZJQ+s/TD8NE9VU6T1NvFLE54ATunWZJd84axt2QIFzLdcteMktfP3UBvsWOogFfSW7qGIcw
s+jmhaxxBp9NpMrEF9QcVI+mIryAD0ilTW/nNB4gV66wsWwxbi4H3S/UU9hPvwcirZjH4NC9+GIF
xMHpQVrnvA5hI96xJ46MJ75B840OXZhKoqX3jaRI16zuGqnHP1eK6gA9jchZCyvsahWCDk0NPwz6
1ep62XYJpRygd8Rb3mCYAfw81Afp3QG+TtffW9VyT5ijQwVinFoFzbHbWh3KsTkhEh1YEEcv401L
ZcC7cUBn5nW/k5cbiR7AWpqkhdHAOxCI4tFcJdDrHChCGMmzlai8lmhcl1tPZpYkVb6NS4LGrtSz
ibwB155GH1y7oQI2yBzKN+qhtl3upLOLTpmZsWfrIf8DxPxsJP749laivzI2EtStu6k51uRviDLK
ah1Fl4j9jO8nvjjh8xyc0aSa5nYfBzXZshPKCgl+T3IENEBPWD2SMsFLzNoy4GgKi55IFpTn+xsv
fAW1Noa6u/j8TLzpbpp5Yz2mA9egZb+rro8Lf96wvAEePtZgdL2Oa0ElMl1FZwvksmUqfr0ITVNG
GdcuAk6vQ3dluqb9n3iiXPoaEgtVDN1yHnMhEeojIqv102uKjJCvu57mV/ZlRFSnt+2LFMvwMyjO
0VoAGLlwBXLx9orIhHjMyPXkZlETp9IRvO8RKyoubLMl9dWZyQ5lmMj6cyHMe7EhHXrlL6fJhDer
iuwcEa/A0N3107rtROErpS+Tj5JeqNN3zOvMKUesvNc3z/bobHusGOpEzOvH1HPCtEP7gTf8A+vR
GhxP0AsX+oQ8zUwjoP7zpsmT8hQEu0jE6RhZcW6h3bPnMCX/KrRotheDzyNSCHo8NE5umbjD0PRT
lkHy3HLvxB7iMBdHCmXhFpLuvhoNlElDkJpzMou5jxKDKCe56PIvRISlTI1Eu2+gh1TTOyPwIM2j
SzKdHfQpBwaQaXD4dysloTmFgC01b+d93vNvaLczxoVOECivJYubQaddqh7uwoBotzOUmS4tHYt4
klE6Kx+SXQwlCAJO1I2g5B2W0wE3grR343perLkRv/4I3V8HtUB1s4ZYl+e2B522UzzCn0CXVJ+1
BGrg8KoKnx+5nM4Xcrnh4Bbiz1dUCGcaGza7/ywCHy49RQ9wXaapKcmJ4oZzxUccVuEjeXw36I3b
/NMNhEYnSMia/QaccNYuY4HwEavcs7IiZKrwPlFmmQIzLWsByLUDSR4rKE2ObA7A+tfqcD6RgnPD
naBFxtFBWyXAPO8q4HqiHMUGNSDHxviO5JZyponz9m/jaM/Z5VqAfi99s7l0syODDPc5OI5d2Gap
ZJT3nrb2o+8TB5flRjXGCNDhaLAednbOfUloTcyzC7TpTVxT93bYl5G7wEXBUa8lWRiEOTxmNqYu
T/ME7Ay44ZH5LmQuicP+2rUY1Yzxu4nPM5yH7yb2qc6rdZp7MpVp93F4J3XBQgVgV7HQC8xWwo0x
ljPxt5N9aQwAHoT3gkx+QKk2nqmMaQnuop7mQzEsjVlhNqu6YrS66ukduiiXUYlTQiqN9wVm0Y6+
tQdQJShOmsO9eWewS2kUsGtICYVAQ8x/1kGBDB0sI4PtV/YQi1Wo43waPm5YM/CU+RRwub9avgmK
Wsw/BM5+5DksFPOzoZoVNfAbqEfYaYkOF4IEDSKbPEp+i/xrit5E30S7AXqryqXk0nxYZi/jE2KK
TglQuPUv0UfQqFsBYSxIprMEsx6UyeIZ9aaWglWZM8v/4gz8WjYNSJqBWUW+cgmv5yRTVd/XMUhM
8QJsB7wGEisrUMxfEYjlq/i2o5mJ39ahEywOx4Yh0gYOEL7AB7pGKC4eSaH4nV0QwUZdmQtEVlL5
NWhCdbLZ5SbxoXt9VZ6jYQSE/NR1Igystw8nTbkAl4i+w+pnuqm7HasMYdOMgWGIa7Pq9Gcc0j01
owPMoSH40r+muX5vI2d2fLyWva0iviyWZQPLca0spOWPs2sfaXmcloW/nAGfOt/q5M9WOyTnGk/K
pSaNULp510nZboA0t2zNgErcucZPh9kNPRxSnVZFXrZ7APZH8rzQDG7HiNi0Agg2s5Gdvqe9/b/h
HAp1S6DzP+GYYGfZTS9sU+QK3x7EO2u4bnwM+dVK5+WTacTaR59dHnvNPgRhdkHov4/6iIYNOrCn
sFdMHq9psTGWqseOYGogI7u01CenMNJDIzbZqeVAzaELKmlk30cmtRZgVPIXtDEal+oPoVAWWuw/
Fm9oEDpEiCbhZXwa9ROWPqQJP7CBS5SgL0mokzj12Ct6TGffuqqHLvoQv9L6AoNdd8iK9JSXGl8v
UXPTdZIH/N9L6YLEfwjHxDW8tnlObW6zvZrxVxIoYO6lyYR4vKiE4/h5hmMkI+r7B17Wi7whzNK/
v4nEor40NoHpEBTUqnpsvmYowLJ2oCUPL82boSuHxSLvYiDpptKOWf2MOkzRq/8aSTAIhVAPsaX6
i7CHouQ+dTFq6mw2jcU/KGJh6VdNY2iElEq+uY9oMtBxq0pCdNKji3ktTyldydXjRQrTh4hfks1f
PcXxpHpUqIXGx2UGjdf/du8Do2g8Iylns75tAR+FMx3Rfgd0Q5GX9p+GS0q7oLZLKBwjAGmM3vIx
d0A5hmuiW4dw4hflJmJmu5xU+Ukio09jULL11SEq9gtwOBqP8MyLNe6bIf8yvXlTKMLwN+IB+TYT
Xi8tzTpNjUGBk6Q8mO6hNczWiNqswMkyhUl16M/ufkKwv2YrUHdDPNXkcI+ef9k7u1XL96Yq0Nm6
UhtaEP6b4lbwO5+zCyZfvpTu7eoApWM5Mb6ICwzuwIoeNg0v4QP1DRMLPLHvzO1bTTv4OO+ChU7V
pSr2fakRXUs8RE43hdif+xLnnefL8TQmgKH+RowmZaSQTOBeP8APDZowA/ql2W0xCAHpbJ1Tf+Zf
fTW8VVAdK7QIjlyVv1muy1WGHMIVOQMJ+pEMHWjRZ5d0KZYsOOE82GldMGu5iJxHGEC/VErHBeyv
wymc3hgzLlbj7wluzftoG3qhRHcgP00biNNkgb83TZuiAZ3aYbJUplF4kTOV1mUHTD7hupCshtrH
nD3nDRzS2azhDT6Hnb1CBVB4ozIB45J9LDBxbH3JdEauLBfTlqJFk6cXwqmZqpsXjbTXZXnGrliG
XPSapPZsNUwncoKPCTj1QCBMrY1A5GV+O2j5z9KZCOLKx8RXSGny6LMaOV4DJmc+MHkx/m/vQm6g
sitdGr46U2/ORkMRaKd+/1o4yDhkOyLali5wDAB9vjfWaVtyOtwh4GVHynQBMU2K1VvWTGsarmmS
aZ3838BtMs1UOy+EsqJEY1ShkX+fOKNRVHPAzw863iZRWRypOMzXdivybY4+ZejEJK7acq6rtWi3
/yM/dSgKpGYHf/GiuC2kY5/OTbHCbZkDlcwYUNtrz8K7JGD8JlfhnSbMsb/32wi8JWlp08cebm1j
obmZSuE/i79WmtJbfl+RyM4xWCtKd668M/6LZMrsRoXhtGogo3ixfM+Sg4KhYnSrZ7apf/l0IneB
LSjbnoIXVF+YvsJKsHSeccop4VU3BjTitWESlIfIlSZE/+qEYOY02vt+P8tIln94kjsE+kg9hlf0
tz0RrEXpLa5jhyMn8abG41NlDUKH3qz7/H/jgnIDWA1UqnVWwwmquP7BOB8qDJBy9rN7rIXuTp1O
RekxZaW+VymcZuQb2ZH8Hfgw05zq//IjL57Q/fu+0MNtRQiGJ7OnKeoNmdzpWlTQwEsYo9w045MU
5qrOiR3oFaBP+mkwsidBm+5Vg7UuB8Idk/Wwxb4IsLINEYp3DBVEPVtLSqczncE18XV8jWaSsoXr
WgALY4mu3HTdYP2hZ0PZlpteHQdtDwMAGma1W0dI7lw3aFnXHp4R6OOAorbnWygyFlk1s2NgKKnH
8FnUCodJJj8DA+Q4W3w7LmC1uZqsXkql98coZWOG/Aqn/HRR9bzS2XnRixxudUzmuqvw4iDmNBB0
7pKyjJaffR8yY0qTHNBNBc3TGGYw0g6HRl7WP+jZ1S8tU7I4Q7te79IvvR7FmaoPNk7rGw65HB3j
l0pLJLvwTEM4fUxvJLvwAH24SJQ5Y1XDpjPK3myy9bgOz9mPlmNnRYX1ukh3dodKdJm4LLn2gP5s
KNgLh4QD6NFwAcDmthYragZspVsjOuILBLWBVj6JI/TjuTcTr7D5cVrXkL2Xri15wfEXJ3bNJeCs
/HC5uNe2IUWsTv0VoYJ3Dtx1JDip7MQZQ5/H0b6kM3+csQ4VBhRwcB8PWTJliCjVFo8kPm7XuMCI
2G/tGekgpK1al0k8MazWmwY4crVrK1x9Dmhu8inmrJkfkMf/VSkL4Gwkyk6bu5gnhMBAFuRVyUkU
9tn4SRz7vLSrL2W1gpv6TuD/YZz3HyO5wf4M7JDZn2wad/hlc8sga7BvU6SW1LiiwZidmZ5eccYB
BfQQ0iVCe+z/83gLPpXy/noFHxCJ0hHUcdDgSw/+6UzZh2bFWqgDicJ1jCJuBvo4d7A8khD5gENm
yofNKtLrdPDcI+8WcL+rIJMGaMHpDO/Ks/sUO8O9XHLFdLKy3KViK5rpCRnP1uDlUy51e+Bmu9sC
tVC4wA2geZ3j8L97ltQRG5A6E9Mv8/jeaOZZCXQpLVVlooqXtkdKmcUW9reP+2dwEaffCIwTgy/F
U0E46X5lsHOHy8XrkQTnBDx4Nc2KZjSxjW8fmEznmuJmX2EAQw80tIbZjGFmv2y0xBd2Fee1ZOuh
JadIaugSijiLjc8zI0gxSapfdvk5+eOHGl5SY/Or9TV/2mNlrgZ0IA44S4XjE0OD1nGkcl9TVmoc
e0Xi+xIBQlcB7Cd0CByGzQfsuwx5D4cUvwW+T4c4E5l18QG0jXCQcVkzHZThKyIOGDSgiY2x5xNU
cxELJo2hUqPClnocBFispp1xWFeryO8RCy2t3TgOF4c++Jx/fUpcK972IsKIYbpi0KvOvWCPutsd
lcBaXwl2CNbtlnoR3p4Mr9U0x7R6MSG9JRG4Ia5Ijnrfun9AGDodKZcCckL+A69WMmypdUxUCr6A
YT+x0FIhv8Fk2GyGZz9Fpsap3oRWShU/2oMzJCvqpjrC6zwwhLyDF6UgscliO6e3Abrm7MzR0zKM
QnG+bdXQcbthBbkju/JvmMm/eJ9L1arMQqQc9aPY1HVrhbV+mNBaf2PqerCcWEI9BPmCxdB8sWpM
7jLVpjwc46HrMNYiDdg3VGPDTteolN9/lA4a2ncz4y96Str8zr0n7JGLikjaFSVoKpcWcgl6TBFu
VaQuBTg55TkLcF5lAMC9XSuNCfdylEs3d0u1IFqq5E8AOUydBvZvLt0yfjaecXpebgZjg78YZsky
3DnSZ6bgPZS7ViCmaiehXFqJA0TwlZ1g83z0P6XB1R+8eq2csM8TWPJbVvzRlMeiKRD25Zt9OAu7
YpVlEb+lsqVZnoX5IqiMm/AJ+bx9hcDVOrLyJkQDiRZAwLFCg2Sz5ZmvnHOhPKj2mhnXAYsw+Yq7
jykQQqTuteF/CwlcM5sDkvYNlvxWATGULSe5zjP7sROIX5dV7dq+OjMh+2DjRMQM/RuFV4RUsdva
o6yKNrfSlsfNB2BP/IWpe7o11eyfwS6N7qYpBBbXDSn5H5+29C3HVx0lPsysOZwl1CZ1YiuiXsvy
zUuF7gcoQNoWVS72pB3iZQ6SLUN478U+Cm54fpagLWLe3sJ5gxLT6p51i/tIuZ6tFPM7c4LaEI58
yXwy8qs6HV+TVxHD2zdzP7i/82GHBfyIhqehSlfcNHKEeKDPc4xxUg4wEu281qJyy94siAmMssdd
tzmqA/GDB9ZxhBu0wqcO8fQZ2EYsIHQ9AdvxMBq4j3r+jW7S/AQ1cMo1maCvM5YyuNQEMucPLOuQ
kjfmxxAbbWCCHv+EKgCNW6oZCSh1kdMuqzWHbIeWrDgE7j0W314kkHYJroGw5hPMoyYo0wkOP2LD
2myNWJfMDeDFc7dNFeXXnT6EoG+5BE3NdilyMa+K6D7J06fCQY4MNdWoeK1G7WAdJMY49coBP7v9
khIogfegHnExqfv1xsnnztWNt7EQbeUeWbtNDLczoJMv6i1YlipmRJXdENb1vM+dILxmB2dd0RzR
zT2yGxp3qDLKbNxUhfxK6v8kajHrqpMAVyKUeVOVmV54pe57T/7Bk29yCG5OhGkFPs+1ZVSSf+GM
EMxUi6/IhUQxaupyqIx90BnyAQlfAmwFmt+J6vOzLpECdESfTkHyHSZBuPBIsAWlDoUVEo/MRjpi
f/h3CJuBnYXHVoLo+0Vm6pLrlGN7YKRENabBx+nqQacejW8QmPmaHmcj2GKVwLGfm2WeRRaEs00I
9zBjayYSnjlMoaYynskQclJG1Wq719ve/R1/gDQjNo3zbRNsPO8MwJ9w3b238UGu490HuOubwodj
Sr5nc5INd46YjWmTxtEEHtQ4T0Haq9XnM8eckY1BNrAgI+/liE89fPyW0nBk53SAibP1MMrYMs3U
zD0dYJLno29NrFHCgROjvOkfGc0A4ct5hwRYL0hNkhtjQAU2CZX23IL8FBV3cRPkcUvnlii0C+lX
Ji88mZ7SViDJrEcvhcXZl5ZBAtHYu2QHlvD1LgG46SfzQY6HI4pdVjO0mzqkK5zNbrtZgzvKWK2F
WwOxrYlPHI4bAkdDzY/p+HnXwNJADC1EuZ3GfpSpJyWRjItTVUxXdmABraWf1KaOxM2w5cWZwkwZ
T8Jd0Oy5dWiwwrwnULDk3GLAxMuawHCYuNHpIB6+5dz2+cm7gb4d8epsBR1jN9zFGOcFEetEAi6U
4E91RGvg+GREp3ffYNHfyBXeoBwlUW77W+sgHGHBtWplthSGF7OaV+dyspcqn14gBTc2+RM8m+of
SH7YTgj+VVW/FGJ/Yuc2prM/WcR1weOm/9MjtBPh56YXaxT01fS+WYDPr8AKk645tHGhzdIZuGx+
pEdfD28ift4zBPYwb5V41UdcKJw4FNamEOjopAyC1FRggzdIzVPTa1SttbapaAUHoYbeg/Dc/Toy
0tmWByP25BGbv8y4xlIJMwn166faqfkrivzkeYH0PGurLXz+VODuhEBNhQT7nE/P4nYu6J0RVfe4
lBG22mdJfs1nhs9e7D+PcH/z9HpczVzMAu15tefup4JaUhkm0udpQLgt+TwqYx3yXxFQxljpX9PQ
AJCiWPIxkYpzLO/7ZbNtkSgXK8gBzxwbBT7lEp1VFtA7+3iiREzp18nRzbxli1YTrQjnID/sANdY
kW5hMa7UY2BJJU/6ElgUxaWjRpD0GJ/mqfrmd6WY49voFEYuJJDIKkiW0FqoSKRrmT7+wh4VA+vV
NG3yl0Wq6e+hkdiKa/zU3tH02KHFr7JETwAAWEZ1Ztai6Vpg93AmMCOOqLh7S1dRDSx7kOwwXTqI
ZvKyaqIgsanA2kK8NJt7RysDmXxzuyfX+LcMmrf6Eg2uf3FLby0LfLRD8+wLtqrFbBwFv7eZTMmR
B+XzV+PXXKnt+sKwJdQ/5PJO6WJEI0YR71xmreEG+utLy5tDxEf7jFSxBAYfrJXbz/tTi+FHGpwy
8Gbz1eL6t4z9FY9MQnkycDclvsOcQ+FyA8ktM/GmqCpCItJdaa7vLHy5WgFAy3IhmbfNG7AYJ4T7
s2YUEQbnu2gx6yK6bcmq1fbVfdf7JaC0KhI5n7N9HjN7kk4ET9rYPrdumrqsbbR2URIqO1tt2JZO
I0qmLiz0RW0oSFmTWtZQW7gYJRHqDMiWznHV9ST2BBM+pdKaYu4aLJoKHBLBSEN5stNdKTemjk+0
cb+UflNmuZfAzjhB0+KU+1kjWJ73zxwwtr0u9Ud3e2GIgU0jZgs0lh2u9wlJOh6uGHsgJczflmNE
baUS6PcIRaSRutpTKS6XPGRVv5OulEO8God6hFdJB1myVMWKA+k3Pk36p0CH87zc9FjVf/7bIY/B
BMMXXLPPxXJafW4HQnKBYX+Y75wY577L8xcF7oSFMZFCio+Az+LBdGoJxm78gyyK/CDxnUnj1wZ8
vIFx1QBRZCGu/PBaxp1LVhIP8mFbA7itA33envrTdQJRIAj1vhN4YdQXrC6vgyJ6a2l2iuUONSt3
JAwU2mRs7rIOJhG7kaJlY6Ha23IyAVQ8aL33aGeW48/ZkhziTDNAFLXvC1trJSi/5d9buNBt1bTW
z6Dd1sY9LRZufv1GB38NLDNE57wJ8lyewJ3lWgdPDmYl/p96jdpgqn0nM+eOhTKLgTK9Mek9y0Pa
DdLEkWyu+FcGDuo6jTGlqANpxNqNmBv232WKxdfVBqRK9/xnnBXoDjbrbb0P2N9w492z6GfbKYjJ
VH/6OyOaJ7jhQh7mdCrfp0k/XZmC1yCjk6bLyutJ8W3RW+U2IZG2NtBE+Cwx5yfpkHiY/utUaM1Y
g+VQtIKsz+ir8WTscZ0ewsx0g9RdrLT70Si1ZQOB0eFkl4hSPr4Y6M08hBh2Mn5zWMexMNebWJWj
HjALpzmLibJ6qENtodUus9c5bftqgfNtoq4sguzAqXnPlC0XLPu9BJ5vi0DoMHdIpKWDkrQeJR/V
Y01lgqlx9Euf24kj3NrlcwaeoIzr1Pni6nkl+urVmaPyoZbO626PpyVJe973u7iCCRg1mZ3Qxnb7
PPZmCVXPOgLdRJfQP7wJhJqsSrP3WS3mQttg3bpweWjT1mhWYXZA75ukQaZmoJOaSMsxc0JltsX6
rlmniNWcQuZ8hdJs7BFhPre54SA3FZdrdNagGHj5xuk5JCMqKBE8gR4zU0r0kVkfUsBEr5ytmhVv
3kkvQy2boZSeNILdIWsoZ+fbhCuhU29amn1+8eN5qIaq948GRNdOQqRIf/rk+ppY2U/OyqNoxH2G
lEddgi+YO74owPizrkkzg8jo5ahdReHzmDCHMRNzNIUCiRJ2Zw62eJzc2d1Jgw4ZsuIchVqtLg4q
u+WTWlaF1A0Tu/fMOQGZRoI8JtrTozvVPqJJLTmoxOD3UoX/V6G62X1Y40npK8hM4Q7qqA/7gMlV
dBry5r6jnfjtudspdqPm8bYCS/lQk3zADU77kJRnOQ4TxAsPJb3Pzh5YEo5QppfwER+grrJcm0Iu
/I7j64GDK3yGFDJWKVuhxtXwjZNe+zjZB5KEJdo+fhNbxS01PxSpGWzbbld3dgXvIsxMZJJpkYex
87nDwIGB4nZ5w/rH9W3j9+QtdeLQhFg1H0viafn5wCQidzZu+6xQEv/LGXZ89WOuC9RJJIZO/jVL
xpGcak0rwHbNIRDaKP5bPBoGFUxoob3HE7q2aIWUch4R+ElsMAYEoxsnClDh4jNuuaZmp/1bCgFk
jsHRFxSOmVv1QvIXPpXpf54cQnGyCZRtR4I4W60uS5Y6HEp35bayqpqCtBks7enkhaHygj9NAnyA
6dV4i/fvHVJle9Yj5TQxGTlKucPZXtVVbmbBfB96YzvKpzp2Lr4fQoK39bxlfPjs/DsTFCrkITw5
Yc/XcSgYHOcppF9T2QTbb+M9KNQ5Sakp8wzZLv5dhkrI4YeiwJhQMvCz9eE+7/7RJu7ohP7ZxUhZ
52bllXZDRs2GfTpJaeisGNqjwMzor99/7NyADeZRe9f8Ftv/CDT6NScTxWA1CZeVbHUIbvRT6UY2
6rXBcJ8yPutJbFcsdOXWUYDqBsuFCXiAGn9o3B/iK/GXMDmB8FeqU9euaBNq54jTrg7yenFL7vTa
nW4zLqOc3/nTKz5LiT/ji/ZgYvNtkFo6wM00iuvGG2jC6oPIqFDRTzYdWkMoCKDCXqIAaJM7kzA9
YJAUZX8Z5YgwCb7kNxDE+U8x7dH1g06Y0ooV9Rw/JPdht8hgZkR4dI8aB0XFZWdRNcqv9LECVaR2
vaF57EZIqm1xOY8GMCC9YtR76Sadru0L33H1C9Io75NoqiYZynCPfNv4kFFsOGvdRKDoi82yJ3sC
chP2JZNc/m68KJDIOeXQdwQdDVWN0Fz0hTdCbnMbWo35kkpDmv0d4e9AVBhDUV49SUE/4K0Tra9v
T362xi5dDD7wcs2cqVYu5p2DiiwgXcetmBN1v1Xkbi8YOcxYV4CgEKlFgn7nO7V8lZqtUZtJp1RE
kJ8Xe8HdgQ9Dz+DT+uOCKf52oRKQ2+n5gEDaHZ6z+FsfVwhaYIoAK+SxB7vjBE+zOTsfN0slrSeT
CI9b71ofNM93iMKMLolBAbW0OGoThirj8215SsTOdOiUXpJX8coYGWJcZjLSG2t+tssWvIwl+n09
KKs9dy9WUcdGeDLqsp8CIlhhZO3rw/CmNU45LVhtZGOzMAtz0XwMAINRIGAiIktB47Rcd/yYThzb
+eapu5IcNh8iAdcJG4bS37c0cwgiauCNifeHfU79yKlMYSsxiECwkwaDI9Xhe/rSB8xh/pc/OJBJ
7ynJeOsf78frJtZKx/XUTPpC1LvV6z4ZInT2nZ+UV5JXA7xlb+gvtzceeNKBZd4L1qBwN1pz3gKB
Doo3+Jgpakxv8df+IsGb+GY3oeZ9SvZKF3ex7cfSB1hTtTxCHcytN9R888D8XGd8mUUlWbrNSUB5
av1XHIU7kdOTw0GSk7Vg0U5TeXwqK0VNK4We9ghf8xcGxOfMZlRQl2PzRffYMt5L0ey3CDa65h+N
zSYcsZmbSmohSryqQAFGWyQAJX9Kl7/aQrx9k3+cJf9d7K4AqT1c+44nLyAUEP8e1OPmqqFYqZf1
PaLvI6hlO/G/GiLGqN9aPBHsRvwXtJbDncpvLEE9gQG85vYuZAFYyVchcDCZl5ZG/VnIZXh0suyx
cW6pi6xYCB7JSfYns+xWkZzJ4It2zQbnEPWszx3pWxNkxrRmNH9zco0sp1lTReAL54THFKUSBnLT
eY3eFyBrs1ZTAPaLt6yyJH71htQmtwGDQ6VPkz4AJ+kIyrN2esWkOvOxSKlnOoiASgyPsVDFZjzB
MvrFjhYIwFIxorhbMGq6pyFGaYHcYjKL8fWVFP7xMMEIxnRKMqMVfxgTTx+KVNYC4haE23GSKyYH
E9Xma3V8PD7HVFuJLRbz+VtfGwIFjc9RyTHHyQk/lY35mosGJLzIp3yPbX2Z4t0PDPM4lnJOnu7g
LRFJtIGwf3aKoeubGbFmM5sZb7j1xQPaIUHJRE6a8/psuqBCIKrHJLebZydvn4HXpxslv4hNYAX3
6AGwNs4Xvo5XDse8FAp25mDlWE6NLGDZvQXMPrQNzZHSpXJXW5nY5ZeDol874MrLiDKqXDZipATZ
1Ps6geKlUSglfadE74DTIKZZXd1GpOURZrJGHzXpYGAWWSK25Xxeq8XLpY83Gim2msLk5jdrx7vG
hUxKF2eOCk6TPFhJahP4sc1AWY8BHrO0DTWWoef5eJaaffThVHqBO53bbNcyk+yrs8hVbNb76Xqa
/K0vUYtMwwftpTQ2N4VFafBTPiwKZHlt/8JzBPeftCS/iCt0UOkc87A4XCKpqIzcxunK64wAP+TA
Es6RxzWfkM2L7kJOUBxMZthL3odxOQ7kucFE2g2l2GZBiMgzB0X8hJ5gAvtpf616cLRhqnTIP7Cb
sp3Vpysd7K+OkWGPPGL+ua5uum2EYzhD/4FIy9wSDdOMcXeEpAlN0e/+yHSzOGk4lW3yCDaB7Bbb
InNDlYlmGhvZCeiNv9vroEn0LqZwODbn02pE6UqrvO+/VIfUlve0gLsgK5KmcpYdDktzVSzD/tah
mBJgLK2swmEsdOjjV/XLX4r19MkLnMrIll7Qo2vZ4CJEO54pgTfd4JTv6bh/jmWHRtyZ3zcu14Ay
g0NNp/4tbgfM1mRl84VpLuDaQFHQt5ikK7z9Z+H5/RSnEXAJ5AkPSTh9Ok3DpadZOVI1majHRXlN
60KWiZqEobZzpxe0TQcMujr7lZdWhMRx3ycARD572NNVJZvkbo9CtIzMTROQpY84YOGd/WGW/I8b
RZ048p730B6mdNhviui9e/IL0sa/fSnLpymFHsktfNo23h0lkzqhVdCHRMpMcShSzf4Uy5yLzAbR
mBflmGXHTlSbUVl4l2L/3uj64W+CMQo+B0PyTWaBYwSlUE8o3+TGmhkLIJx1kuJgKFkY+hEp3xJR
aeHzeM4vxhMLmkN1MUnJxGbRic89QTTnKtWjKc8Zb/kf519/Ckne6Yd1WHhBZqe4Yr2NMb1P1L4j
3QtmyP53UNG4djVGMYwqN6NFj5HcvRZGH5yXqxrLazT9UELlUcoLuj6OtofYdWtEQnbG1LFOF5X9
TQxUOLB+gUzpVej4l6pkYjB7xLt/WVcmg1gVXOD9A8TTSVXkkpdtu0B5XoiHTflFN0ZF3PhJCV/l
cdejMmBbsFqILYR1Dyzs2E4taZ0DypkgGjSQB1bbDaN/LE15a+apevxFkDdEWUyQVOhGpsWp57Gk
0Dv/K049GZvVBOsrASil5DAHc64YzHMXjU9k/KPIbxMhtjucYUK2i1u4PJ7wbU17AQ9qcDa+1L7O
say6vqzqmWGbTvmrOTW0gOce1pf50VtEZ+584/ZsFdbw2zk1KXUkqV44j4xDjOo2mJFXbVU0mT2N
ed4MdbAJsFQn0WgDGjzteEEtkdJfWxIZOeko+YWkdrXHX9jo6WqJDVtojxTbux01Z/0Zre4SwKkt
atDwaRzZbX2bGutpGgo1vG/5Kf6zgI9/TySV066Y5BA0WqyEURyZR8yHBcsHqvWDR4xLGu/t/Ron
mkuP6Pzc4rzb56fSVC6ZzJ7rdLpXaWGweu3Z/sp0hCZJoKg+/SbRE518iQ0H9P6+f4rF4cK6VlL3
H5DxU8ver8N9OGTZbALcI0DcJ1SoB5xAz+/NN2H8psg6d1ALFXExBLMcqrCDn+rMrWUSbyXOUONq
/1orVQoRofR/EmFDzMOISW3aXuULV9241mPGvuDNXghaUjqQDOXKHHxcl4ciu0sLjwV5OFQZDYgX
tED2DXRPDf4aOWWNQqYqGNYjs5dZiPOE7WbwKdUPqBwyFtxdQwEIShPUyEgx4+3IVVPumIkpTfih
vSItb01hmrglUKvCLTPSNmZuz3+J6s/jwG36WYi1IyoOA0JW4zzJo4Fkt4RtOWDbXuk3XiSyqMTc
L/rjyHq6q+XYQcmeV1zFHBGGYS334Xm3GA2bFAMIM1PR8f2EYTYUBCmlJshg/BpYqFuAxVdMfUKV
a/tCYSdn3I7jIC6120lhcyFuXDadRiPdo7LVWkMIdvjNSj1mkCpy/0tlV2rNkXs+NTOHQ+H159kU
vyjVC0xaNjdu2rF+0BDex22xn/eAgK9JsDGyQ7OMmh7EMJCc8eh5/GcOCv9QizObigAnP/EWn6a7
bGDDXiTpmK246bzNnpvh99im09wc3E1wXw53RpCJ3gUa3S2LzJpvRRQYTzyYahS4MS5ubKibz8Pn
Caa58wd2op9oWjMP/e7kg6zQH7+0e9T45eC+71gIikeBKPW8q7RFDsRjeb7QvNIhx0RcDyrOVM8q
RkjAH4ytFz/Bs94KXJgF0uc2OOZvEDgSvLZ45QebWUL+FbECoSfpYtKqKfSOMS+4X2I5VGa0EXHf
EMYHliJMIc586mPG0avsdpZxMzrKZk03udTlxRTMKQWxlywLg8glNlQSDD6olmdlWF7XPI48a164
s4W54DcqUr3aS7vgD+tXv+77URqyZCW9uSlBl5QUWBtq5EZuO0XxGEN+yfOjKZZYZwGoTTqgclZ6
+EB7Jmdf6pL/ruPA6ROYFzPWylmsSOwtDK3eQPYXc08mtKn7rGEhuxcaUbBn+47+0KV6sbuMV1fB
nJg8s6DZHSLw+b+GSnR1uzGkCV6KnNeZ8ByL6yVyAgmdhq4FBV5yp+iL1egcySrB07rY+2AT2Jym
OrYkr7Ngq1wp4L6214JRqu7Il2mnoI2KBV/KfKfLN1AieUgjFDIR15HVCapEo7eXijcuTbDvSWdn
qUIKld9GCusO3x0rQaiBuf172Qq0q+LVFW12wcMScKLFcbMPNXsyaBjbOIR+A7dO1E9MtilxwqmY
RQbvwNj9AW4PCy6vXTaG4WwYcwq3ss4MDl6akh9BngSJSaLIQZn38yKs1ibjAvrqhVme0AZOEHYG
uqg2VawEei0WH+uiC8rPcJu9JrzwMzKDrHu2+m3UkLHSFXh0z55qi4nVT04Q9uks9DNQ2a6g5G4M
YI+ofmzrh3in+yMRBia+/br1qc4YCM8oYO11zQYwJtI2KkGVTQaF0GwJ9TSqltgkylIzCc7RCa7I
jqbgUgb8VN8dpsVoM4Dc8pcKu6KeV1fT7VImqsDIhME94irDnPzFqQYe8JKmlZB2CbMyG8OGAcDV
uMYPw0IVRmkOMTQY7iINpRpIGFtAcXyQ941UslK1k+xGxmqRHS3NTSToJGckzihuD2fywjQz/HRJ
fEGOV3VLScq2EHbvBinWkeDFUWK/cCMWOflv03vD7GqtSIJ0F4ALtl9ir0ef+N1XHtOf/wLj45qf
ptHfT0xMe62grg+YyaDRU+qj+pmITrqzVwSGTlnzdJA0wSLWdCjlL1uTzF4mes54lZtie+oD8VvI
b6NeIyXqL/KfSrf07wCxHHIoD4sOZoP3HEIZKgI9c17DauNmIqAb4fsc5DHu7yQ7C6016kEvgcQI
tmbeRl2DhLXZSw7LAKIJzEkUyPW8mVoVU3gNJyguujNdrLoXiBevfzZ3KMOJzbw+GrE3SvXeYJj5
LjnHWFDHzz0qAwCwVIFW+k5y4upnxjOOy0CA9I4Zhi+VuxjUaFvsfwhgVYy9yUaGWt9VPvjo03Ao
s4aZnSrHn+Mm4u+jqW6yWt9W3v/uj9+o1ZWxzYpNv6MkItvyX9BZqplt+nUgkrqVsM72rdbKi01r
sB4SLEm+6woces+PoPC6/zu9HTgxpViREL/Wj/LF+6ZpiCsN1M+nh/wk3/yYsTRlWWbPuMwtop/e
HCWXrHRkVW4+YkwqtVBU5JRgowB1EfapbGFGOVJlQcWetuMcZWR9SS2MFnRRLh6vjKBzr5hq/kIG
SJq73xwHoBzdrRelX+5m/ZY14/dhEH119XKvaqAxZ39htE77HyV/u3uu2jUzhbQHw37qwEMAcu8U
BR3xYtkEuA94vBMEkWTecZ1tofUzK6WXjmx+kNEp6OtlqoTdstbjEekDtIrewnH1O1euu6Zu6BoX
xtdcjJpltX268wFjiGiA2libLEkOYB1yzumvc0PLEuUlPAak0csmTWy5BOaFuMfjezg+LFZoAMoY
6gh+qPBdMeWu6ZLSW3zZ5xU+3HWNulEosooOfZNEemaxrGLRSNlsoqnR0Ymnyq8uQQxvlpa4BATt
SB4J7rKhjKsKTcCRTgxEQIpxnAkagFCUK3JdxWPvVGHHlg7i7Ca76gvUbs/oRFD7aUJZ8vjWikZR
fG1oLX+wC2knwawb6Y267CfcWCaC8H9DEG4zQAfnviCnhs5oF57+jIpzYTY6KeRwIPUeZ6ETi/ts
Euuib3T7wQOXyFxVHIlK93nchwOtuaI/MQJbZeQswqA+TlJwPS4wsQHYZduuTbbPF95EvoJiMyjr
eIlXVCroAJz9AsBqHjcnhZE+x6EP4JPnvDVpP6gi6a1QJ6i4xK5Up2DNAGVix9aVOmHMMCkL2jcO
uXE0tKibO6ZWVD69O93qbmj2GZEenoxV6ma7jiFagqFLV8ti27BaD/DdIxo0c5mmCFOcISGIMOi7
BUjbnlsJGYPZKxn1P4//9FbxWnBDn/AKnv2djIJyZQrs40wbL4LgKJVEeW6DXKzfDVb35E/WIOnp
R2w7QHqwbcy4mG7E1vq2MLOUJl1AF1pu/orfTfMBUYROj86YN6S0X09XnEYlxw/awW06Vkro15BH
Vur70IM3R8yi9voiko1jFIrBUtvmC+M8M2WcBHrxHU1W5afd4zXXJOxaSl1Z3xMzCckDBP7Mypz0
UcdM6lcPXIbolUqB8nk2YJ6pUrJEAxeyB7JBskqllPvTrGr1Bcckq8RG8yHGb5HIuBbEdIZVVN1R
2foQmKSPpDMq+8/IyzWsL7pymw6sEgAs3FKeEk1FJUb2ok0+2dndeALX4+3wpHPeZXKMI9FozXhy
zBYzwbq4ETUoMPHdIOhmuq1RG2GEvLL/GU1RctrDI5f+XHMO1zbDUCn19O43QEaUlKtSjeeqdyex
+P4TwmtGhaNJlXy026M8ORY3j7BGcOBbAIK58k2bVWS3nHiXumtC/5UZAOSdUhS7C/l/8jbXwx+W
cgGXG62id7Mhm25NjWWMY2VLiDq0wCz/jgn0BCjZYeTDK4HIIBagaB6FgR695jrXoD4v7SAIGHWn
Jg8JqdKNDy72d4nKQXXuI/J6F5rEnOmqgZM228lZLpMR87/mJyoXaPG99k3vLvJ39emyuZ3m+uuM
RQ6KLojNYpoXT1WC6IEdLR3oFfNm/DoLFb1GDf6kS4/S0osDuCX1e4naCi2D7djPMuKTmWXvNd2W
x5Z8wVRXF79MR0+K9Xyt807Yi/22TM+e8vZetZrLILeGE95sG+Js19NaVrRb8l1qYAJm4VlH5c2W
d0SXL2VGYa83EIqIoTY5fjq9aYVcpjfXLCUblm4bVMV9mFE+uZ/TliT/L2J06bfoPs0wjM4SINdJ
QK2KkWz6pL1LJGyQwG3JBxm1eMYZfYXRlWnsgvoeGCvYBwQTSKaVack1OH8KtRdfg6kgyQlaMioO
0rsAJvfbcEcgEL99g2CkHN4rDF/EdmEPZWxjwlAZrqc+LBrHJTYQbJQrLU3B1v71vEt3c7i3Dn+0
kKgC6iKfAeTc7imDqDrERQk0ye9DzG7UUvpT9HF9+BdiQgLX9L96zjv04gWyZ3zlfmnV2vgReQxC
Qzwa5Epg2o5QEIWXRCpUSPIWYMIoSZl1N1YvQ8NHySh8Ylh3iswoJ1YsUKSiklV8PgmkEN0VckTG
BGNuF4PXhKD6p9Q8rn0YC/jH0lGzXgn8cp2V10anaN5Xdq7NhEpMJgxzk09woTEpxXxwt4hl7gDu
sYrdxYrOLD6Pp9fY5zBtKJml1Ezfwo4vXey0SbFxbPLy6Hq37gc/FIrkcMCkQGg8r5c3kploq8a6
DG9bfpC5I9boPwKNX+GbF8DI5AINDUBB99sfr/eraOBJOIIHf0IfQxYDiFPV2LniChx2UOf34Ef4
itDvMzOCZ1kT5dha9p5V0e472n881RXHTI5DJRjsFx+pGk4FlXQAB7wm3NGFUAVzh8lWAGBwsaBw
ieA5f88KDkjH4zoNy65rC3ORwV03oUaeGx8/VzeAZUXJDG6OPP1SYhTpUMmsE6H/eC9psp6Y5rRQ
jnizVsMIqI6QEV5JSbwGOEnOk/XmSZyTcsSu649g5ZcQVX3gs5ge72Yd/2E3RQX3z5+8kCktVdqL
sxry4Ok/KrhozORbSuQM7TMVtxWZ+Z1rG0kB4vFKQ+zINKrWNb5rsIDSK95YlP5a3j5TwFcf5Ydh
QJzi5tvFGZLsZu5OEvBgWo6/JgjZBqDYNugYMblPgbM+8xj8mY0KDHszO7XFtCgGUby2ZJvtyFrg
f6/WhYXCF1IUOPffVjQkBAzYDi/5t2m3epOPCYSehbBqewH4zmvV9i/RtkVLkNjlAz1CdAJj1pvU
TMZ53p1A4QHU0oSuwWHAZT9gBItcewevWDDM44Ra0KOZ7BYohHtEfuQlZcwsvmS1HBrTSEIbjBWa
K6JWv6gvkyGpOVbMWG/zOXcB+m/RwNjJaF7hXJs+mbdWuuKuq917XDxbGreHyAcHS8nbX/O93TQ2
7KJ5g0oWFJg4Wo3oP/pIND1pWP5lSFierXLnkR1YfAOw5Sg2RlSaHonuEIYOINB3KbBRCsS439Vp
uxemMOi8iptGOAJaVwL12KBUScZRNgEn1ngGw4erd9W0OlyJLK/LudrJvzKmZRJYb+4t9zf/8Fy0
MbkDv89WI3Y77GtOE+WKhCDMGLo2FEtguiIQQCLJbg1NkSz5DQaMzxw+2ipY2U8rBp8ELP8pCzPq
MNh4mVxIoOeq+Xo5lB/2+iq10rhaa3eUrlb+kWUvg59GjvFXK6TmrTrDLN43DHXxDt5jRDu6g3eX
2ZZzFdXMnj7F6YAfxJjnaD+McKwfAqLosdA+aZH3KweecX+ebmLP9FcAhvzmxl6zWiR2lQFTdahQ
pmcQrbNM7yzWmFXYUxk/smn2ICqmoTvkK2sP24USvC+77Xl+ZDKIxVgqUKP9eVWZNSayrWAc6l3T
xClldQ5CwLiJe/FHrKsd4hFuJ5R4dd2QDa6zGu/nINl4OpICHSQ/hhWeQpfEMK+5fpw7A0G1e53S
IztCkNCox3vJG7RHCKu07Lb00wFhOxt+4b7b8FRjPLYA3s7qG1TyE8EtzZS653p16qFFrfk7rX2l
sTgz82NmN/LwGYGjCQYcN2Y0NNJ5jH8MoQn2mxLEVnsT6P6MkMPSD5ymuxtY7uZ45Rx1+WwyuExl
vU1ZqZpcSBova9sfeqVYB46HNIancvOf/gdGCEGD6kzDH8knFeXiB7al5mr4hYRkDf7j01yBfSxS
TjTNA13lgmgkf2VSL4Ypy2HV8GeYl/MDg0aGnVC9CS2w1mrQx2L2sxm7iWgkDcXyKNzHrQ7sFKXs
ZAOZ3dR3d58byvirKosIlITZ15T2dN2JIGlT8YN3lhfWT0WMvwnp2cSOiQit9T3vnc7v1KQ/kkJH
BJ6IS6VDGJ0lqMBksb4P9CyMfK782UQVzRi3Xs9rFbePKbVbFJA+OlrfjS2ogE1kIz0qWiOZwodC
l/mwOba5Sddr1hq7VD67SKif52bGIV3PNBEkB1TSjN2R3PM+KbQDksICBQfyPj22HiwUckTXw0Ge
JHOttnn+GwgYYfjSnVK6dKyIi9W92wWIl0nDl9TK/Bt7NFhh2+uGtllqNT7J2Nsnoux9af4xBYyV
W9ew0+sChB7wBiIL9lmrJZ7J+QX+NbNes2mZEaJrtOb5UjZeGBfPTEQBFjid38oZrCzr7DMXGqTv
mu3PPr+q8AVoIpKy7Iu3PGxaDIAY7v+uX29ahAYpzIl3myzVz+GAQ8igrCJ21Ttfe9GUnyk6B3Au
vkp68ns2LFb8NyIHIlZpyrf4mhA3QkRZfR/KyZWz5Mewl/dIyFVEcrxbtTDmzX03rB5UQSALynJi
0rQKvThMboPZxcNLneg0VDWkVGEyHlc6mgLV7N/jIzkQ8nCDjh6DBg25lrL8a6P6Q6AqhWsJw7bf
r8MzU8bSvJAA8I2Fr1Knk/2DNBt/kPZRYjxpRSEawWAVesdvCzyNvlmmdMfAZu2faSh6tumLt7Lb
4y6uwn2Q4EdDxPXRz+wBiq0H38NuM7xYwOwnkXdcpCyImZvoywdqVahUiDoJ3BSzc4Ucvvr4+gWH
DApU56DWIf+EM5fs879La3sgh+nh5j6p6f4glMwjqIT5dYqUfxjoDkiFixzk53YvckVm4c/es2kP
nVd+Xe6rL9ixPdiSdajk88261xNmxR802DafgIs1yibdW9rI3FBYZngJCZR2wtUMpLQbsOZxtI15
M5fgVJtykTS2xA3iqD2+hSkRGKURPJm2FGraeTiom6UdTDqxmTzU4oxO2TVCFZWrBT1WfA+Lt3fc
gdk5OsH6o9Z0XFyaf75mVAMhpoRzfueECLJXOz94u9xEOcBno2kTgj7h23s0b4U9OSevriafLM9V
jk8AteiRgaYGQghp+sKDSHuoM9ZuADIQebs70uyrbqF2yqqImdt9gpMfO/YgTIdhfNHpj9gegI19
WjQnTbNKc5jC22h9ntfKxE6q/oj5TVO+IE6jNOchvzuAIoXQdifZiHsmw9TCNGf4q/WP/vr5CbwZ
L/8HfGdpKKlqs/5Xeoz74wYWorSJutJ+3hWurVN99/O7+BdPyR0q+EALjqNMttPYICs5u88e9dte
mCgJpV/ZDVLgsf6ugFh5YPkKYDx9+wh84KB0gaSPjz2RULjApUmQCHRlmzrV3pykz+gfVTkIKKlo
c48flPCw7HTwyCKARsOE6iQcvg1cEQz97Tp80Hvaul0SKWd2U2ORuBrHvxFIa/xBVRmKnorjEuhb
dO8jnZK0SRz4BG8fZaw2roEbQqO5h3YlRHUGXLJyP0dRcaY0wTmVQ8AmkkOKtnBPVp19csC6O6Wp
cLCgDgODjscxqsdEOcfvviy44BFwk7v43SbvkOPgGn27DRI4KnJfDguQXbVxezoVJCEaQwpXZxAU
WzYofRaO1nmjHK2S7vtxHFkm8z6LuNa0xMtVkOPZFl8peLAy3gFHqgcW1fLNH7l/dNMopwv+XYgB
tU5mz3FiBj0hYVYU2YZv4LLAL3+SB1UQ/RWuTmB61UP1rMgHmS1aHlrnkPcRoni6cHUFnj4KhfPi
OnvOQ8wB8a8guRbqdEVAKaWbiVucC3DhPBGhRJR9OcupX+EvfKAjbx6FcePKPg65kpzV2YLKkF8f
JbMeIAPXcfN9pNYai9O2JxOSyS+6aHamLElzUaqGlfSKcUKW8RCvFHVQbKqGzwslVG6oIwlzGTpv
a+uk2qP0nBG9k1asBT7NKUBbvfa7FY6PYs1QVXaxb0KuA8sBpZ0378eJG947o+y4tPcJTiTqVS3d
k/ws4qZyGAgueiw6XdNMpQ3T/cUb0bZCZP7LueeAqc/QqPqpLgk623yVyYa/qgzLawmovoCO03DY
AD98Pmys0jBgSkbpLTQoiRQwHORYp7yach81xok0jX/GU+VIrbZu4OMmI2j2102LLsT4I+y7DI7J
2G+SU+YnApB6Ah18WKcFjRS4JQ+I0C8XYNQGKyO3y5SgV1C7BZ8uBH/+VVXaRLkcSz2O/NEdaJqa
R6j4OlX9+5ZWUirNjjqu6aHHhsL8TPsr6FAMHVrNc1VBJHNhz0JRAAW4d2Y/wS2nPWj4d7AvJRkh
sEm1GUnmVoUgevM82SGF6S/eVhdKJ/M3fsThyexAfZgvCw6ej6m8Fw+uUP2I16eh2LlIvu+L993q
OAPie0u0tt1x7XQ+uK2BxTQhRdfBImeK1C8JqZ/nhnshpLMgR4YK6VVz6Jyja8CaOxI7O7SMfDiZ
bD1fvRBeqx6HRBb+2FJKzMVAT7y/xCT7W2c0hYN6ISL6XPe8ORKllIqgo+D5xuPWWZqxd0PiIWNo
2TIruyJEE8zLa0y+bJKQYio/wQUrqm9e3uKYO/re5yRCLTq1L37/msmvk3306NlGz34MiPgVP7er
NJMyDnTKMcfFqQLmacU9ytuEU2epfbRCXsL5HQ+hKNCDgowcysUo2GiSIVjkoPXFs9Bw6Yb/gULa
OJFPeVgWk3DIaQZV83Cm9/TON8+srjsQfa4vs7M0Vg/tXbAp+1Vt07kM8336mX5vl8ffX3T3R6aP
Pzx910MEwbIdNmCbUfTSJiIh163ZV6W3qzIwrYynm3YznBJMW6W6/Cd/UpfbqSc70c/VCCFOtmX4
IDAs2etukrD+Rfl/WE725SOJTqolS/9aMwlDZlIMaCAAY8Yi/Z97VTKuPaQ31D7Gd6gEdACtcUqt
fxqdhR3280v5UXLxGLFbN9n3fhNZwTC+CeUXRY8CdJuP9slTX66fluNC1jJbYAqw16peYTmu7Rnv
vvyzit4PmPl1+8cjsmwCCgyNpU1HoBm1lKVIWqyAnCskSl2pe0+McmicPcnejwA8vm4W2zqhY1R2
0Qck7AurTAp+SIKfeWJn2nX5MyB0jfiIhjQORIXw7BJ3eV3z0d8WAdgpCw4aZW7dZfJxWwx1m9g5
VlE6uN6eBkq9oqlHxLgFY2MJSm4XxkrgnuVd/u8a033lzQnsnC9XI5DgUbutY/byJjikLdP2Fd4M
mbGPLth+IscpirsLQ7oGJKDeaDMJh8qlnVtDGxrGE/CunpU02coOLUk2E9iQTaBx1XK0LlzD4mur
dHgvoxolNixVLWqJEzzL+afVLhksUlYjZh4C1rLPyAV/Eh0vYkWqavK/leL7K25xUzMtMM5o9BLZ
fw4Hxy/G/9URoOanGxMwqOXNIHLYhwKY+ixEXTO6nWTL/PcSI03yLLvTTB3ty2eTjgnq3HCJO3yN
MWPnquJPEU96HESiEBcRcZWDLkB0GuajOsTWuzQUtuQR/hudc5GkeYouizYhWByq3zjw+fyH8m/R
xbowkeXllwwgVMeM3zApyeoPz0FjtJN5wGw8+V3f1i92bAuh86JVEkOtCdTlinNgNlGxCsxx/x5L
7ZhfzoMVbFo2Adnai7juroZixU2W1rFfQKcyt1t/6d5V/TCDkLZX8Y0MhHXvke/geV39pTyvyUkB
Mv436PbYOH7wQ5Z+YBmbKGRrngyQbfjLsedgTukdNvwYKLU6KpO0blO3X/+J6oizPWvybLxmHYTb
MVOH44TUR3dx+Oi/SWoNSEIk9JYit3Ya4Q3qh9VMvjUEH80iZg39xNQBddjmPgjti7gERrbi4hWD
0docqS4OdM1dcKl2bdq6xbwkVN/v/DQ2iiKf/9gQAMRkBmF9INNf0FjkMg5qEKIMER5rk6Htvfa4
hADYkBOgySB2nN0VBj/jZgKDlrh1v4yRZ/NH0Dv9XdNS7fzvBaqwrkVAL6Lpbb2lQtEI4DrLK1bd
sxobpTCrS6wZ5mrkDisgXVdT36H+dmLGj6Fw8tGeg8U8YtiT6+HDXNsaY0y38garZLtfj+oxSTWZ
rsOEdsW0W3ZiwBkUBX/v0MruYJlyXiVDS8JNEo8Tvt5UvCNgBDLubsO8oFXkNBplU3vMy+1C9rma
Gwcncc8ZcPcuUNsyhdTGHNNMq9igZXkoSXznNBSpRZfoLZocn/iq1ez6VQ6EsJLKiT969uvZHoq0
oM9SJve1L/kR7VQjN9t4jTFbMcUZ4T/cffIDhtgeDVYLCV7lK1qgLYlZYZZXQniiu1EKkv3RG2Oj
Fv62jIP18dzhqXwOF5RDzfVDL8N9sZY4AKiIB0Dx2UvSCcwRA2QENKENgEm8wWNbbZHmYK0uLjWw
r3gmfWMD8VefRLMUN3jX0yzG/r2O784jYdhgtzuwJsqRVETsFiAklFmHYrg1FGu1sgZ7QHzGSfJb
ZaC7tTxLdv9BQdwbGwN0rV4aMwvUJfwhAhz3RWztBIlE9YxIPVh4+7XCi4tJTC8+3fxAFwwJF6cR
VRgiUQDKP/eWxTC0PsKL7WlH8hTwqDmUU1v2o+ev4gJ9NonranmyJ5sHXef6LBO1266OkIztt90a
Y13xrYbBQCElToyieTBK5KRASokCSfhqd9qQ4b5bdnJ6GEzmDJVgG/0AY30h4YhgCCns23CyVFja
XBu0HWRz45/bWDg+ZyTPQiVnOY29MJHpEqq6I83Evx/r8Y6eA+3dBlfME4VK9e3KtgrOwU5PkQyl
ZbuuAOqor9f+DVK8FPRXtba0mopRD84F9pFsrgw/BjxTB9s2NsH1KIHSgnHkh3ATUOz9diCCxWma
G4WqopFySEXNXHp/+FYnfZ3jkTdEIHdonoT5MmoaUqXvwWGOSTUKtbOBfTsxpJxqBJKfJZb6Mld5
bstm+dIY//wda5K5BmevCdSfr/54LFjA3kmygxqmtaeFZhgRYCPRM1vmf1TW4WN7A6qoKwzk664b
2A6lByps8ZTW6bZbsCSuHpef6fVfsKqusqY01Ra5xNUnyuEz1LanjORCpHjZWghnTiiuvlDpcHRg
pa6t0RtRVh5R28rQtVqfyDJpCbIYehFImBetYjGpb+EeuRaUW1L9KORY6eqmhrGXpwnT2VrQoTpx
iZY+SEMNyk6hjekz2iupyve+QeD2crwtpwWqaAdS3dfl9uS7l6UyimMDMe/kxrShykA6Rz5Bz/dj
hl8sZ0WDQ73RTvbBOoDpNIIbmQ2JFP5Lo0YRdACdshn0vkm6d525LxUpPk1a+pB+G46vXdcADFnk
IbCqD39ZS9XmAZLQNRclCaPKqRA3D+xW9kW/THMINbJ/n9L6PtiM7sLpv+bc37Ik+sVc3srCRY9o
N0AjHfFtip48L9KFWJA/ki7XJHCL1JSNr38OlLN/isf/5j5Xqp1YqgKUQjyPKLEEKv3iAKlE3XSZ
J+2Kyj2LXEXY+eoqTAPa4wOXp3OkztZtB7KKZjjYbJ5O0nqZbULn3f4NHnelshN6Ekh1o9Ppsc3L
MEBmzZ+8hE8FLwZjdomKbP+dolQQxEPoNiwVtlque66xPBg707OpVMrWAGz2bnS5pLR96IW/+FY1
r6y84cRxfOw04SVwHJvPIguzyeqz4KN6ae6BGWxj+GvlqL1I4cFbACC96v5hHxTGrBH3EgWZUdk1
K3EX4Bw+22SCb3zdTUBFThFgmJkj+W2qtb8YKIYAZd/BtpBG7Acs5LKL66kmhKsqiDfVLzPBRlvJ
Y/5IvBU+GuQOSN+ujdQ4zX/5MCTRcONHWfNa4jhqJvP9GnQ6ZfUq8P2A8FlSBYSrsWsRzRrC9sTO
t8C7KEpk1vfVp4HriyVcXm1dSzYeYgkab5Fu6OdBk4ySkGqF0ZkI7f6BN9IxzwOeBotcsah1M1Ob
iNhFp+yzbD9hixYY594IaNcfg0IKM+bvnIitwSERF9j49yCxLazAv8XCkJmT8hPpTJNiflFKGVnc
TL0fQzOGyTWifB9LdVBOwx7KybeP4UZy6305nHTqWShVOqcWQ8+HzfB0xhdzeqeYPRCrkAbqwxPm
J5IkxyJH9o/X0EPIDBld8rWo2FlCnuOb1axqLgaiWFuyT/fDnWX3L2KGyDlIBkiVWlnG0+JovcPE
eMaNLaFAFgL7lU09/pbp3IVuLahx1J46/1chcTGOsvF2GoYKRZVOo4MV7l5tyFz7+cLTIwWETTYw
hAQM30AldIo0WBWyHRjw1OpgS/N62b7T9Xy35R7VS8qB1tp4jaZ6jeDcN5WvNrjkNlfraDU5sVFD
gPJyTLmyrZxe2zMWZT2v3HqWVH1uFTmGyCQrvmZD6nUFZlQ8p98J0PRrtmsGTdBdSqStqQvMms0t
ES+NIw/FsHoq0ey2yafPLJVRAPCRFkFQnbZzQEEIsA/rXEA/FFx3E/AjDFvORTQ7l7OaZ2vkjaxq
z6KQ4fHj1LBf5+D0DIL9WCTnvrEAJ7zU7aH0Uc1dx8CohdHB2t3QmVZeiaO/TE5p2SV3EZfolndc
jroj8/O4U/eR2CuOHY/kxGPquNbPi3rUCDX0JG3D4i2OImB6y3aHhUFWsD9f+dpmLImTakMeCtUE
JzcJg0B+ZCJvpqA9vEZaAqHz5zDDLukdXPkFEP02ihAhiz27bRxqD8bFemXijPsQBKs/uFg/+i79
BFtcDpaxUPmzG9WM5QhNpi4pk1VrGZT7NZSA2l3kU+tv4Sam6Ksj0dStVY/H75ZYY+9QBUMXNEVU
fBrKe8n1jqzNeToWSEmCkG0s/SoJe8lpte3KqnO10IgRIePSmP5Ooa9ayMDQYBveLsaquMZ8e9GM
aXcf1kZ7E+cuFkX3FmJ4+rj7q9nqXKjTCC7opMrbnb3clNMHcMC0+/eJG3nQvtLFuchYFQ5mqIqZ
gpI54wZ1w/4citd/3LbWuJsfNRLLQbeyX/aEYjbtpb0Vsg1YwuRt839kwISEI03hXugykwaLy/vq
se1vXT9BGrXViYVNmenMwv9XyzoTCGTz0wq2XKTO3u3t+5QWETGJ5r+WNVVZWPr/AM+Td3cCr7P8
QYISjQHtxmxpiYxaOwHaJdMu976VdMUcU1gSl/0xFbbbzvrrUKOGKaYogldeKNfqxHvVKjjgV2UU
D7iDv4X+OC0VHvnH3qIYGkQ+kHTAlg/O26wdtR8pcz2kNcehB0qlapBlIjtxOCh49efLhA1RQ9cL
dI7qCJYB/+k82sU+p0oAxm7MQasedPfctNpUPHg0GVixwrGhgBqZ082RHdjJMEC4EVx1okfOy4or
zq2NkeX4maC/B/jTfFVcRqpO7cW9uiqjzJhlw/bXR8DD2/fV7kSzfdPpKF+KJqfQa4Q8QZrDUncK
Y1X+1uOmC01rzqEDcGBXREXGJ2XNCEwctJLuuiz6kBqStj1D55ga5jRyyrTul3Or6jyiz29QTgqF
F4w0sq7T2RosBqJ0jp06nbZm43d3CRy9ymXVXJe8FONnMxoVpnizl2MFW5c6e5uqGQ1dsrw/uzuq
iV2YC7mD+b4kY6jlW/s9U/cCj+jsvyTb7Si8LaWZNKmHT+BDHIWELbtlaTbQLGWfx9sxf4NCETLe
lO7vYIcUzpAZhgk+GiC61nKKMFesAlnppaD7v0aGSu7dzSqdWNxQBXI1MlulvHGSPkorhYmPujFC
6o7CoZXc0zLEwlAZh8WiiaArH3qKJd3pbtXGkXOfAsfyUIkozSZN5LDkRVs4j4ltEJQc8i8S5agn
5RvQ39z5xfm62RzfP+3i6hpzwqtaC6Jt4WtA9uh+OfsKb3/MGNYMHohZjpjpFNRH0BOt1YhiGzkL
n/xPVqczd6zR0h8/jPrImLmtc4yV1Ym2Xk5BbWF1mlYQuUvl9EinpEMQzo+yw0BfNbDqXoTzjkXt
tv93v9A0mmCfiG546/SwbgKmU81AF5eOWnPuAYobxSQwJejzRvQcpQxEnf6yCiEdTFLtHxvQT9si
7+WfL1KGG7aRauV85cp6TL1EhhxvgdbBbhSB/FqJCQ7T/dPXR+9EmKcWUOdY6YpBMr9zOJJATm0o
Usl9e0b7GzQa7NrytgS9FcmWcMF/IBovHFr55FnrzryMEK/oW60y+eKBlY9UAJUwfCNXwymFHj0W
Aepoi1QH4kxiJg4HbgJGuDCy3ZkoNBatHKCGxhNRzu87qS5sR/Qqpm7ZC0dZLdxpn+ORUc0RIBET
7Z8PbMrIJoOSN+hPc5HNY3z2Cfjb9bL4y3/LUyuNBAeD2XmA2vpsbvaA/yXeXxERMpT6d9f73ZoU
cK0ugB+edK3s9WpzRi5nxIvWVMAmRia4f6xuBD6g6jmzWXX3md4LoplAyFajlspRMlGd57ZDJBRk
kkHAY4NTIAXj06IHdsJ0n065LT6c6zhfOaatyt5/78dPvfpkPmUp54JH3qouJq3Kq9oWZUGb8UM5
cU7pI2pfq1J+nrLA8PQMpnNuKNu/auBSnDTzEYKcYhHaiPINbJt903O3fAiuUwQog2cVCAsGBsB4
2kkcfH2GooMi8ykM/kFlDziAFaUgbt1a5akL8rHPsryYanaAkELMPlz3rW5s96j3k9sz4j9XvKWG
pYWod94rIvyws0k8kjkZoVu2LiIVVH9idHtN6YnSeG+9L0yFLoXkcU+a2O77uax6P0OrCnbM2U+2
TIEGmk0VA+LuhUEqIbKo6eszPja35VUpV0677ZSX1+othtNS/VxkfLY0HCrSt3SXE4VJtocLgiXn
FtYaGL4aOBiiaPdVELuTFJrVCzOaAJ3JzeUF7VohoQVgZQjAgLdO9bF44FneJDQ8KWvaGuXNMa+I
BzhklSol1AwWEDrgiiIXlgm+Hk85Uw/EkpLhjjiVKlI1HG9lcNhgSV89bO7RJ0jr9ZTDwmHizUSF
Q01MxEl1blRaat6BP7SeqqeBklknfXy/ww/GBc3K2Kww/7DrWsJ2iblQU8IvoTmq9WChv4U5DiEh
a8iB9/Ep/tcJWbBfAvTIC3XUUJde2y6ZElT27sWOZdAp5W2Q+/TIiOzDfJfFVwrOQTQROlqNsHod
r1+NXlioB3hHvJJZ5nEAdqu4YjEtkrYNsr8EZrnlhkgRLlMX7IvahfXsZTOva236RNcB3xFG+E1y
EcvcKnVeShpv3/f0M3y6jsbHVc+XCgAse+Id3mKTVNhsCjcYm6IsWtFJkSlf+krViYwcOgOGtqah
UL7ZNQyiE5N4vLpd3mv8Z1LODwPdfVlpKUFHDcb1lf+mekJK09cLO5RKlhKx9eb4B3MUDawnAdtr
W4gFtKaKxFa/USLUjZoSxW1rVRYay2gIjTxDodwjEYyNHtYTG/ebH0t0r5SWhbAOAfC5ir1fz01l
WwuUMMF9hKmIawi7VtQypq9FhIKZJgqfjlM8yv12wgzueaZihEDQgPXIsXnPb/WH6UugcH1XE55s
ucQzyjAnUFxE+qdLzbw1MgWoP2hlzGWSdlSUIr50V14p7BaMKoPo2enAMWJcNR69lwpZmZ0kTMH5
C/ZhKzzEfV+f3M3W3IyvRANUbVu/snFylfxuuRxZ4/8cAfh82aBNZU0Dkh+6jsYGezMvXSN0skTB
Jz6jH6NAnRMIGbXCv2L450aPyUeY58bhsyF2q2C0dqdMQzlSp9A77Kd6Za/rs2665YDzKKJW+8Gg
Xn8DqJ7jQoDeTQ1ccQ/Mm9DR0ZY2+fP/7zQ4ERvFVaOQX1kfpW2qa9B40Qcl6IEJmn4n/a25XOd0
+brwh7hCg+zzmeCEEhbtw+xcZM6yZ6YtkdzDaw/nuVcAZiFz0idUvEjcWKviUyrTu/Fr4O/DqSAK
0KEwsvdWZMFmjuzS20kldDOQdsInMn1Ohj1ayP87zoR+c1cGSkfgdKVKZ1R4ktj00z/gTMwbKbp3
g51nhDqncNCwsOU+d9/oQAH0lvnGONNi1PyGJvk4C8ZRYwyylUB9YKyWS+NTkEpW03Z0r7jNoDfy
MNtL2nCXUH40peFv66KT5Ul5VC8sJ6GYW2uQYFf2sj82BixxwL66I3gjE2x679a9GZcueJC4rZIB
5+Hs3BlwtKIY32U4zpEcwNJyAawaaY8cnckDNxJXQObRm24jwLFQx2Ub7UB/Ui5J6lXRCmWaXSjH
iPlrT9fvXJuM4SvlW6m8GVEc1h+dnsSERxRR8wqzM81906wPIvKGlJirCxexzhc1Zmqlbgc5ThuG
tnkIbltuxRkyJPBr+pfcAW7cx9mdmpEUS27bO5DHmOpfOz43JuyaX3JIv8700uQkUSn6DNj6R05J
nMNP2n6xDH34e+1k2lhB8+QY6txBbUYmmUn+L0M2c0podkcC+AtwWl4Hnpr3fwkzw6ymEnj401f8
XMd/U0mq07lwZq3NYxgF1Vfd5oo0gBFKtLsKCsBUWOb0hDqjSJKHoN5FtRyIU4ju5QHp6uoFulNi
ieBzTFPJmdE26n9Qx72CxprnBlwMA1KK2uJuHTDxqSijWQe/EQ7ZStgqemKOl5tbbC4aTngdqXka
dQap21xnKRkskuOdui7b6wkAoRZIicwLkSDOfrs7rOeGJQ+gDYf4Z5ozhWMEw07i+h4Wny+eo59R
+Qxe/ZN/3Wpt3OrMCH0urgNMTRtMvm9E+88nyOLVrl7FjsmJMKXOiqgOAX7J3G0It8zo2bPy6Dgs
fVG34ymuWg4HI36GHz0VTqfQWBCV1B9J7qYYX51p6tVrppFPSUoj3gSiXs10gwpoEzmNKmLigu5h
QNye5rUHRemtjD7y12HkPyCvFsgyTgwCqvOZhUfyq8RHHA96oCl0NZKYo/gwlpE2xWWmOMvVlU/o
zXfsuai9cDvtrMzFhTbnvRKTuscfJCGvj5JOI/WU8ET7ZVzAzH78doXlRS99oGfRpS2M5wi0w0u1
zXRdq74xyJdrKleX2cbZ7+3Se8Y045vqrj8Z1Okbc7BY67OJ4P4Hc4bNkrF9+L30NZp8lD0jefy1
xYlOrBf1vwZy8+018DYjUt17Ek/NmaVraDDMeB2rZN07Hf2QJAD8VzMGNnepfmopluRlTXwpo7hH
hEr4jQVk45y4GlawVnIvEjJ5pFXQnrE1xIc/xQWj4kaOo+zv3y/z3r7dRU1wwfvDpvtQSfwjSpGM
zIdeyNpcYB9ZBDPU2pHyShIuAcTCglrEIwKNTDfhDH7/1bFZH0TS43iorpvDHu4zffrfegymkZx4
59lVro3sCYOvcpRy/Fp7/O7CzEfzgRpQ0izl1n15zhQOniB6a43uj0sHDEV6ve7+Ne6ClYv6wtFv
6hNjogr4UAUuq7/j4gjJrpGSm4UztRnew6RL3cojzLN6AAl01NusabeDe9w9LGL8G/8+up86N0YO
6Khzp07bvAITSsEis6VugnvfuqxWeHNJUU8a41ZxGrOos1+jYw/bpWCUJyk2KYtWTWrhYRUNXUwn
WSv3VLZzR6aYk1p82xT7UT/Hj9EvvzKigoBVb7sWDSxHL5VsqTYkTuUomcP/GJIfsZE+LUEbCu+b
g/zN3lcziXLKZFod6JtAJGoePocseTtYA5BGx0HY6RdrPY5QxKYuPlwdpWGe6t2rO+ib+l4FwoXt
bhGKTBfPrl0nosfJ6FIHJvojNKqn952K4lxqQeGxWNHZ/M6gmWJKfAQ+sPNwsxlJQAIl3zTY9R2m
A2+r7wV1TjcPbASCsMCyksfThBpok8Yj13S3vgZHDX6Yt+TEyydO+SS83pf8N9vLuR/shYJbgTyw
7vMMi+Tk5g9gi8JgsVOIUtF8QP/8Zs8kcg7dLXF03T26lviGwiMFuzCmhZLu8RcqalBtNOihboOF
RaHhVFkod3GsUfqn02ZhD46WgqEHqpvHwwhCJpt4c85+NxvfIeXDd12Etaiu+BJdAOIyGBbgsglB
Prm5hprvkrllYpjc0juvVdMgyy8BBN4oym+L7oNDL7m+UwJuuxfQ3oXaWuUbB/I43DGJ344xyOdC
9V+yAkWYJu8fNw15USKxBO9qnMBsWnTCVONzzlzsKR+yKHlQqqJ1toebnCJAshWD6fihxJhhaRHV
/8BBa57DibM/FaRCntchb5OgYHlJyWIaF06sU1TbvHGbSsyo5jCuG3rfDuHkIIJPWyD1YUX+BecW
KY5MsvEncLAzO4QaJdqMk0OP3cJZ64063c32AGOtPUT8wD1h0+1ib8h1RNzEF68yJqEzD+qdArty
bDQzm30sIAtQpsALMhSd0lAm+j3M/GJN8gBJcdKSF0is/G6JrNZm3VuXIKx2eXInrj6brDPCHL67
+2UOUErksXyZ41EwO8aj0bHw7JMNHvXoyS7iaD4HP3waRKy9nZCkohKCMON0RB+sbgzB4t1Blcld
9OLSewj43rWzhUMpzEPrpFb6t/BkqPUDPkrwfuwJu/lTKO85CTTBT57IwtMpWdkHbPgMuLqrHBxc
TUQl0nXGj9xzT3C/Noy0RGKVa/JgoNCz4WVXTg0j3O9uUk0eN4L8LtYpcXI0igsO3s+juzQQXv1A
Rb6H8wA5iVZ0h6pO33fHTjMAKJ3mfUDwpDICWLBlh6Blp6dbX6J6ejaQm0dlOqVQS6fL+J0z9L5T
zCFdeidxRaarS2+oiUfTroTxx4WrFk5e80x9W0H+YEavCzj7HlY8dV9uyFKX9m/04nP2cpbuu9dR
fofSrTtVnWZ+gj03UwoCH1Q9HuNe5qQlfwMPzleoZ8VqlU0dfbqUKIEgfxoN7cTMO4w2vv8NcRN4
kE6+3Q6FR+9nrveM3bC5N8EMNQhirjMHj6sbkRGOHxEYOJXKDkxkxkQV8FJXI+HaHVMnJd8tdD/C
jajosUlVQhZedjI8ZYVGNXZEphh+7Lruk4MJq4yODvgsHtQsgdbP5zYBR2Ew3b23siashM5Nx2Eq
RZHCAXljhM0H103BaYxTF5Gl6kLld1TgO5shqRmiFUYZ/NJ7JL7z3EXph3rvm67UysvKdm7bDzF9
K67hj2TqcGqKJpJedExp+eSDkQmZy6sbn/+jDTo8G1qPZqBjRQceA8gms7/OG5cN4VpZ9Mpotf2B
65me1w0KYA1srSV2LUfsCtAFHT4TwIQVd+oRt4tFbmoHBxDHAoKXcg4LRgo/zsHDsaxnQ3rmj36V
bNiDBR6qifZmaAqoEVk4KXGZRJ/5NiGhhqTv97xzxIykns6kbsaHDTaDfQAd3Yyumg9DON0ZanuJ
Ux9Uzws130t7OfSrwhlKjyJuZ1CFyC4eqUTbt0q2u5ymYzENY3QQBezjIkCeZ+EfiUOKNjXCj90c
+ENRZQsHQpg+BFKRBzgc9qihSBqtBaitbYJuVQzonYYLfK/WmMe/OTnynyNwT+0GNix0ypru3MU1
So0o+G25ex+IpDEwdIq1ddE1qJ2nPgGu9r6jzgWzr32SmXqFApy7nUkcgnpBV8jql85VSXR72Dwj
MikJFIcIKuO2555/VHcLuYXC5BEIMYrRnDLJCkotgexSRWYXzKslrwmOIIBq8tT9gHgaS1FlAlzA
bmuOqq/vz6p3iim4Uoj5DHOdnooOpSpM25MQaK1mm4HyC3cz1i4oUGgRdFZ4EU01nr15WL5llJpK
kpz/IZGHfZAOAhkIyHhCaWiPPoUzk6gRS2s6BVRF8qjj4ldjqOGJEbcqLxtb2UKMyfVLFEGUZGGU
W7ihz7VnTG/7Oy92UNBYa94h1PW95MmLqaXtdjbGVWV/+R2C8tSBWCUsnEaDaItvW9SPrTcm3Tcf
W0UB9YAvuLj1P5rvneZOqfLeJC7DLs92k43RA45Yr6gUKLp04z/YcDU3MdBEzCMhpxoDvxFOyqbz
dPx7QMQLY5CRwCeKnHZZR6/NWHP6czrmy3slF7Hzh/1HsJnwWQOCpDFP+y53V4MOdWnx1omT+RyY
Tx5XN/kmztNBt0RxprI4uE+TJaWWkt4gGEHpG+E6hBw3IiWMJJqqTBcJ6b8DXhoxd31mwY7eCwrb
6FlKCgXid8YTncXYE+op/jgpqNCKDjeVaDpWfF2J3AG3CFtg+UdgmmZ+f1pB4irXiRNp75+hNV4X
3ZZm/SGKyxViERRHlIOBfM+7eAYNX9ow7iJdZjupgOp+fmp5tw1irbv1YoA9unMBeBOaySDsHeLy
14Di0yog0PP0ytcqz2qPnJwkENqot0w52wu3XvUwdLp+8b1bZmmySLhs0FWbNmBu2IZn2lAYNWZ7
ampJp8pQmJB7oeAbCiB5lbV8C2ycSGY3QdvJ5p+rrOT6jVnASeewhOiM/gcIFXVUyd8oBzayZTSH
WtjBKV/OgTototYM/z7iGHzp7Z7EiB+jcIqH3EneO7kp3rY1gjFZbs0h48RgAHBZEY6jKY/EI4xe
ri6fFyIZqT2fR8ISJhoRAqeR/HkOIlgDRhvZOoMqcYCN1Fuu/cmWDMDMvttDb/2OwRfJx9GzkRBt
cgLlugqiHw1v55OQNSWKHIXq4xj93N2daNMB3qgm+GaRt/DIE2QOH3RrdrIUIrbW6cCMCHhLub6E
RQZn9OhBeT1Yo2UvGupYpelIIygFrLiHuzZTmuyNYCU+Ykyz2WKSoZs2yRiemKo6pslt5QamyQ57
T5VV3REZfiUa7URad2lGzXObR5QFegPJR7ozrK8NPx2+WT2UwdUHKymIkwS/vNq0y9rxFYf1CaJP
XfsCJSUFz7fr16ow4aFCaie8rUXcTlePF8hE+93+mRWsCUzmI+EUBRiU09GXWac/E3M+YTXygXCw
tRnks3De46qQT/AzFn/z9G/GZIkY8NAa9PxyVkI4zBDaBuWeCJqa6xYEhpW8vfGrPOpgDU53Bp1X
EZWIkRFJjcKyvEJeGVIHi6m+wklx7mRTeqOOVGRUXghudnDdDv44XYKEyLFb0grTel3Nzm7zEU09
oopP10txja41rpdyK36gQRoL/50FxiL7h0jjSJXmv+lnBzeKqBAPSyxKQvN/dBbycQdDhxWrFG2n
Qct9dy+54Hxhq9wX4o6VtJME+OMMGh76F7mPGwWstEXs9ipvWlB083lPjhnVgwRv/h0rOilY6kY3
6SIKCSV9GD2yGKIRHVlMktSobpg8mh+P3fc/X9TLnPQkX2kmfbJtquxkbW9PkJqxXuQ6Q6e+mC0L
XR7ijZjS8L2VP05bvI5ifjw8c/8Zj5WnzyVx7b7GGqKnznF+yJcHX2VpZ3NrgtNNihXs6cudvgc9
tQbzfg0/KkmJdYiwqzHGXkup7CeDijF/fzOrRouxeBMp/BzLa9mRqVZlHUtrtdUdtLvGQbHM7Nj4
R0Z1KEYWTKPvobG61wys1xV6KMjjcE9gSYr+ZG4CR/vUtcGTyIkxeqcmeN0zrpNbEM+J71iL6auB
Gdr0L6/lXGBt2Q4iDSlxCj9nU9yg/BzSK1o5of/ycQayc8LomNLefdRHzik6tCkkIAzccds+vivR
w8j2srFjtqiyOiv3GcNWiQ3Whh41LDpG7QxvxKqtQ4MBogwhQ1h34L+wj5euQ+jMj/kzppHZ2+hp
UyHbRkmJYoKeBzdsjjZkuOOTph1fLWfhe8s95z+Q5RubtJiM7rEScJqVdK7HycXZDWm3v9VcfT4t
w9tHz+eHS2YKcV0yB/9iILwaWixmV94+0iSXhLo7cjmzJ7dapa9S03xyQroZ2LOGZROY1JCNlVvk
O/whZg/dY/njoFJUe8dBXSEykZ+Iyp54BFIcd7a3XBgGFLbtcY0gDV1P65EC8MQQIdI72eEUyMVf
VO+VKpV3UL2GqmjtlIfGHVZ8hFkjV3dV3usbcGhGkSooimkHWHGQjRx5gj/+QpMb6uHpb+ariH+x
e+YgsnM/TB4opgc1DbZk1tqG3jj9fLUDJO9ceWjrNE6v1/SU431HYMy4Z0JGA5isXj5r258vRzrs
HvEKeimhZskC1E0MWc21C3UtnkG9P/Kme/WV+jjE/zZzG5rh2W6h5q0tGOqFAW7HSB9xzRNZWI8a
m9Tb7xjqcF2plINF5qHsHVJMom3wctEKE1oqJp28Gh9sg8/YJV355itbw8w4BFKR/DmIiiAN0E9M
ALk1VpAWKBEFzMUT6Ry7/rTtub/56v936md1JJXxxMfxE5QhEIKLNKL+zMov2+yrQTBVdkzu0CGa
l9aggSe/rKhTOLGZ35sHbARbaHoEmrt0EIYM0Z0X255drymDzXI6ysuXj4/xqThpqPQlM37G64qt
SK6Q+Z1FA6e2oLt8Um3Lub6nz1xoKjqulW1qL24CZ4coQt7j4qKFjhDHRUJM66fzJvigPoenCQGp
Z/TTR6ZWJaMerlwAC5BKvlSUzMpr4cqhKd/U5Qd3iE0EwFCSof2z56JWK0bSSV8McXIeY5N3IIx3
KSnXF7WJaY2XIxeDUhgFfbaH+LDOsHkq0ZBX8jS50jKjIL57kTMVWs2sH8cwCtboRZ9O+0fLC9s5
bWs6U7kijEYijIJWlj5c03TdMk1NuFCHmKMNFIjUwRknsG1L1s7xhV6V08EUqVKXP67I76Ob3esx
yKv6nU2nCHz65bXeqPasYW092dpkzMZWgnFQ1UupYJnDTuqOqrfbHYsVgSbiO0uPkIq+iGk1QpKc
2HmFHTTuOQD7sXSuuKBENMagb4o8tjv/TIsF7VpeUspf7oBNI6mL6h2CK7orRUoZk46jjzLUBQd9
kycnjuMkRA1Mp68Q3Dpus9vsZ2/r57RZZEr06imr04d6UXnyV8B8F2RBtNdnEtihHFqK1CYYeZBl
0pAc7vEYjdNJUWXXZT+DKpn6SsI1ZpXwTS0gtRC/EXBsWR4ZKX28PIwJD+fDxVP7Is4lNukbzn+W
IUNdU7Qheth8RzPtkmg9ctPaSBRfF7ziD2s9LkpDz2vgbaY5oTYIpkeEE0HZII5YZOsDmUc9JJjq
apU9mEkjfEtKqln01/SRuADjMdtVm+wuMRJqgdHNrHI8XfwsNRzsbSq+E3xm38MwQzWFLDFp745b
H4NRb7dxtM7TRCdkxhIXOd8NHNJevcSAuDulX6DcPmj513DZcUQIExy/OpqqI+J06sieoxsTc0X2
Y/0DihtAh/fS5h1ttmC6FrtlS3OSDnWZqF6pT8pyehQwL+Zu5iNmRCW4k7u93hJmpVyIK5BkjzGG
jaWn9PQMYJBScZLgojjKn97/Dismq7kdoA4cwwYBHDHMOLX4wNWKexvsGEwSpi5QHUvm3+lg5C2o
GnaNlZbn83mrEh6oSyunfeTF2+VUSPQvHrSAkk2lLD68ZNIPpv6EWiuasYewQKA3wlVqglG+oK+a
GAo/jz30OUb8ythA7HdbP1ompcyMrytNF1JLuP2dfVUaFs/W0UitRjL8JztAN5shP8s2lBf0B/P/
CPzSjDqbM+82/NwXG/BCdXSqdwPqXDuLEOYkd4NZLVz1lE05z1cSFfj2CieAHrUhekO7xSV4qZ1k
znpqQaTrSFHRwFRERGWQ+P+Ynp1mAXZxJ6J8BINnO5Gi+ZBu5uosn9pqIPWpi1HGYP2a9U/KUn8e
Nu5yGvifZd8AZCTobVZZDmAejPZGo5FIyYFERqafZ5v+dzsg+aI+wfLW/Z6Xwle+B3vpA4vRetrx
+WzPLwVgXaDbRZtbpeii9ZkQ+0pRrK3O85iOToWAuQfRLtS64dutIJabWEE9MZnPAODCmPmOVX4O
tgRV35hYDe22xRfJrag2PkJklhivtSMnxTWWxhUKxAcAdH9IH7LXrjfVkfTDppN3qofPAVMMJj8F
YcBcs2NTlCDw5UQblsnikAlMPNQ0zpsNZalELAMjHpSFrXLT4v9tj1JRU5jWm6rZQLb8kt+/bfkc
ny7/9iBO3ZBkUiFD9gZ2CZqGnhAhQb0Bdojx1XTy5UrN57qGw/ds5S6eET0R852wNsvdQBave1/0
84Lg8eCnCGercDvtAdUtW9/8YrvWd4BSn3yHR/XAsuNKlGgaCNRrcu2XjwBkNltBwo/nDRatFJGR
1N8yz5bia+AGWOX0xv9up2GOQMXvWcnIayl3/MFIZf6HjWK4e8l1YtOosf+yBu1O76qk+DWLOZ05
k292Qr5H8Ari4lR2Dt1W3O9ose6698Qd6uj7hNLGtTftPv06nZqqonhjkiG7pXTOlLGJV52OOB/A
xhMgyNYXnSOWNoQf4wwkgKhxCfJpxZlo4evm4TF0AoXUcVnvELiY6lCedDqo7GQ+Ua2YnQHFhtEs
Fy8r06n/vL7rhKoBQuAReovAt3F3ZgyjEnf3h90cgupFAQiKcibEXiYT3uyb5BiqTyp0B3cgpoDJ
5iAATZvU0e4lKQkuCQYYLIVJpBZ/YZPibUHbeL5k+g5d5plkDWUAww7Ergh2dtqOCemQT8T5xmVj
pc0FzvEB2gCgyY7B0Qzdd3795ueWKBoJFu6UiauoBrAkGq+sMhIc8MoJw7ROD/asDRYl8N8DS9Fr
lb+HjkXdRyviPwRkLoNq/7rR4fv/BycunsK+rYvuLe9jH4poDt4DZC3CBuo8KTJHXwyYDAv0jPRK
txtTzteO1CnzMvs9Edl+IRDK+IZotT+HH7ndyq5vFJXSd5u39pAP8sLi699cuy2UmRHH7b10JlZl
8T7hMkRX0RDcUl+jpr2k4m7S4c7CR+gtMhH1Vz3dNYiOmAp9GdT0RRLxvTc+d10bjcvCN2bUFpPn
430yC9aY7JXekil0Nr2PkcrXXW083UTNaMzx8F8Ywrpp/zVniDEExyvtr+y7m2iyUnjpWuGAhths
xOfwfRsI2SJHx66vogNf5e9tjyDAZaPyhROCu5bL+UexCf1JiaUwiyiYsAWTasXasr7sSQR9Qw2E
Mhs2oda/G8n517K6HWnDxu2Q41mPI8pgKksB6AGPExaGe1fe+EPvHoEZW0z7jSNbw8fqTjFICC/d
EEaNG5Rv/KufAGgvfhExxajFg6hUMofAzah7PLz55haQZah5cdw8AFLKj5AyIlDLdsT6cbQVMHjG
731yGPDGgV711UsgkU325OOXtGVW6+5qb7/Gp0BPJdou9xetv22lLPCwaD/WHV94GxCAnc/JkfWe
xmPmLhdZWGvhygKfnorZ94Xn4VSslpoFe9Zo44iRpYkS0mljl0KXBUHs5tu/RqhLifrTaXe3f4jP
Ls6kPqwJE3emKcueG83sNNkiCwhG1E08XvOQ/CSTHkYBlNnsjATuqef+fjUEWplI5rJnhyx5x4rO
Ijxjvz5vnnRNC3hUCz990bWH6hqOWLqXDrzHQqxiw0Tb7R8RsadVLw0NqvGSwCVnA9e9kRDm6HfB
L/FfUTyoFj8vgFAocpCiImW4qNCB7IG7BONIqZGabdczIlXpZt6qtth/JS6mLZ71y1IUSISMWh6r
2ifPW63lsaqlJ40k+sbH1ta0sJ7dZsdvdwiNPWrhSs8HV9WJHNpniO0xZcyJKSFI+J2kDtpxaKZ6
omX8bLfKcfg/mfR5WFbapv3a5zXGFjkO5fLwziXq1gHAy5oGx3Vuxvqdoz6ixr5kbue3H5lr/0aM
PmEbgzs8sUtGTizV+VOTrea6RMLwNI798TOZiAENSXKiTHXEtumUa0nM0BSf+nVBuvJDcreWlG+X
IyIcuoUm55Wg6iLwCuj/NTHPNZH8V+w0AwPptru/L/2vySUl23EzAOm1v2SSNGJHOYBEYFFhExRm
vM+6d9trkHFx+Cdt5yQRsmFFHWcYBB6iKgoCPJf4QEq21BmWT53bcrCwpxJgBMbXEHoV9NdnPCw6
nRJUdMTjBsmkfwuZbPqH7I9PELrO3kd855eyhF4MDp3nB5XhsSCuzgq5fXzz4/B34fLaYsByFA/i
VyGugrpP8/bUIGhqsYBdgt64L3wrEEKWEX5ogi9fIq6jzp4pgDxJU6qEo+0VHMWuZ30Ob4iXzegZ
yytK91ijAprFgQji5LkgDfaBHHMW3/LslycIQ5l6c3c5h5S9T8zktEnl8ytxse0/mdPiBiTVzldg
tiFNiudiLi0qsHC/HY+8ck75ZC3rtCO6bFXn7H3e8nqF54zU+n6rvVy55pePiwBPMFG3eCA72Pif
0AiIvK5d0WM+t5na7BgL6wGr1rKpdeuV9sG43tlFBRBeAG9JkrB/A/Fs0sk3ZE5x0KQ+1cK7qz6S
Yg5LPx0WzlB2WC+r7EBzfpjT0J/aulARMgHSbwuPVg0Y9L1q6JvO5G+Q/Tk7nfVylBEUqNxIxGnO
4ddWfIuiiea0CDK2iS4qGyT1+NOiM/GZGM0+LknVvovguLL1/WpJbPlctG52+e+Sg5oRrs1oWAbh
8f5mUX0Dq8KOtKyU8+x4OzZYX+N2vwflQPAgeVoBaFkzcBAVDMEe91I9Q6a/gYWlvKYAaTxBGVGD
rYH3HLCLo1zcJoF4AaUVSufAx7bGbuOMhzdTBm6I7Ngrsx0VcTr6B0Lq9t3pxEz+QR+AGlV3zBYJ
WoSQMkEeq1C8PgE1vc1sZHUn1NgpQTnzu1tKh1qxRI6iTv6f+UJsqSuIW5GgTbZqyJX7kPyRex2x
3m7XA1fW9OL2mYC7fACdWuws18VLYq/O1eg/So7s34JGEBeyWCI2O5fcC0oKDVTxGCETDQe7G7RJ
6r9SMma27GqT3+2KtR/WH7s0wCNpKIaP2D0jP3Ke92l1eEL4gSgOlAJLDpIDRJGAtKRvCy9VmpzI
69HSdRL5ciCXcWamMa+xPkbmm0407uvbK5a+6ZNDaMAvMP+KHSBbEWiQ2SiXtbC+y+9dtZ65iWYx
mF7iRmDG6doU1/vrJMUK9iuvW3rWE8Z+h6o3BuNqR5aMQtc3/YaP5VcnYkTWcfZdNxCgA8xOIofY
LoHQ7YFxKZia0RH5TUigReipqplWZAqW+3E1Hj3m4zorUbLGIV7XVzAsJMId5/FrqzvN5UddhuD5
VB6JnC0RnAUpV96KcQIyVjgQYq6aVtX62XKlwlzRCrb+px6CXjKW448PSfqasvyzp/b48MWtR6RV
1UfmlaBpDMxV5Ix5WGCM+9F+GMymDJkn3QvlYuRA2C+OlA5b2zFTBL3nfTM3zyAQX3ZlMy2LOy8T
+W7W/j2zX/1d848Toi726GOXZIW/F+rndZoqFPFH+VPJkgKYExAwyoNx9om5U+ceI5VIzfdOsPnu
7rfCNmumWdW4RSdEvqPufdvKSqdGB0m9d0VF0QyfWq+0wA82dz4+bWmLqjy5XRb5K5wEimVpF1qh
VaUPHVwK+mVB+t3HVTKHET+n2Zf28FogsvuhANSp5rZUGhgjFxZr2cbNVBkS8B+DFF1GlzktkwLN
VxKWl5KjsyS/za7X8gi0OVAmTb13/sqMbX2/aft/+PNEyNpWUzWxheTVZ5QBAGp+veeV38Liiamc
+3VyDA95BseShFp31pXIjMgkxqQKQA4d59tBoA4YoAkVWRis/WC6leRuJtGUVaX1xfpW6mqxtdKt
1tW3/JAKjjO+8GuCuFJOBUA7VW4oIF1u4az2Ym4Pv6HWdjGwvUNbhtCIEOlLwqvJ4SFdb29YdkBk
BtBDB3M0kaAeaLi80khf4dQnBJqYlpf0DHaE5vPBmb1WBEkX5or+qqZzxxfCjzygdRKnxe+O3idb
7JqNR7etNhv7cjazMx65Q23+u9TIl1icVikYZ3vhjQL/ML9f+96RQVhaDvYQyjLIAKe+qxgP73pi
KpsUD0msAGGep1Jnl5AmZhY6RvTXVQM0wiulOcxzV0sAnN39/7diP8GX9Cq7CVmhZoSjDQ/PoitI
n1Jx+cX9G91DSlpDFXrpWSidyWKE9LbnF1bvvzYwhzPnWSAGmBNVR28DmkA6tj6aBOAX4TfxfLXz
VtPH29+UtAcqfUFIjT/zScSSjdMAtooiS/JkIshYzYLyK5sFwlJAuJAEjELrB2rMih/ml8/F4O+2
ADSQJHrENMJ2vwmf609mT1/ZR9Bw3rBehV2NIqGw/dEh7AM0mIOvl832ismskCA5q0+0mYtAgaIo
H/b2xTw1kedeUVUjxIMAu26nwMyD3WFxLz2JIhAGT0vWM8Ml0rL9BGC0DG51Nf+bItGBqKY6cl0W
B+Rt9In0bcsAGLb/njMtJ1FaLh5TMg+IL1QqGH8KxAju98ja/ovo3r6/fJfDOdX6SxCTMcz86xHz
IX9Mh1oImHhVTy8ZkWa+O4srXFaiQuP5npwptaEaZA5nM0dJVupZszgS1C6TVc+uvh9EQXSf7dwK
KEEnFIhzMIZsmqJZ7ZqmBKA1VIwUvVvEjYGbcLXw4Bn7Fpaa7fXrLL42g1QwCYfWMR0/rolAMBl7
l0RRPMkCtFCsFD2p1Ney/7qxtjV9AzKW8xky55YtcEex/sREZO6p3QpliyGSULrKxLu7gAbaVKBq
XcRXt11wrcAwpOJ8i1L9Id0hOcYEJUz+e5nSkbr49HJInHrGP2K0jEOV2RJIhMibmC0jJENupRo+
WTGNWxpHN/KeWL3NBOkKemhBsFXc+uDwBZ8ptIWNToCe3eHx6aZWLWBmcK63WEN2R7tC52p3n3yG
s/iCS0HJ7bZ1C8zBEx9L8iUtm7hVpAkPtfbshc3R0yiEVUUWnEH6VCgyHCQRWSnIRnM//CdcFimU
sBLY9Ypk1VGxAYF372HJtyUxzW1VG11fOfoKf1w4Edgay2FokxUTJef7kVcQLF59Q2Zo4aBowRAH
j1qsCWMpCMUliPF45c7t/Y7lGmgiX365OaKGPraqU9wbSG8IMLNG/t1fiPqnHhejVwK4bXgXNDmE
MzqEsXQIZbcUBKJcuoI+eocjXvcld4rJGcROrf80KIgGhXGl1D25bJeIW+siq3N3XwYLYPP84P0N
Y35RhLrydlP2t49J4bD1gcUzVioDC8wLxCX4sE1s8EwS5mq3pG3u9qJJZzbT5BYFCbCSqKbBZR3q
/dmGIBu/M5RVyFTRtnumUR1DMHhkwVK9AIrLXG9QPLLnp1xxz0EDcI9GIO9/sc1gTxMPrE6jmgkI
ZINIZaHLZgLx0rSxse4pj+hc2iTek7EaIvFkv4vPYcuDr+ncNunIEVRPgAxlieJ9hENEzRFPRgsg
bz6NtmElEZmR14Ydy+NivrGueXaP9RH0VYoLtNsSIveVFf7+94Em23L9F9vzVGpIQRNRVF2QgKrx
zxuFICD+9dnC0I4Wq7gocA3hSIDFeyznUkwKfBupUw39sj61/evZbfA9fFkxdt+6btmo9H3HYn01
S17q+75xO+VaupO8d1q6s1wrEFh8c1AIAWv3QCJ0AV5D6nlSJm2MJWNqWbxFjEIqa9aH4R3NBTzn
3XnCG47bH/xfMQ8adzrt6P/DweD0t7aF0jCoXSTZ1j3ff8rEpp2qwsKLuwZFnXJv9QLqcRwylrZx
Wr2JHnfuwLT7CHdd+ZeWEXod0vqsRFR/PBYtF+PsknisE3qVL6s8NcxS+t5b94yolxW+OlvrtBDP
AjC77yWPTlHrk2lFZtntc5f8DPgp28lGjtb9ERSl1bKlFn9iheZcGCPosZMpc7aGP9lxy33/5jMb
FRzazWPOj/B9ktglLQmY7PIvi7UZppLnavSGuuX9umuSz6GOfA/sET7dObj/Vzt2c4R1eHQqCrxn
51quTM2MTqw44FGDxoYVa3l8s5G3Fdy90I+IL3Pm4meXj+OBNtfA8P2n++TrFnp0U6tl0AZIeZ6h
dMqKut2V+Ep0ApBZEnfmkEet8P+H0YJmYeLIR7Bo5G2yrdfXMlKs06erS8wZF81dHE1CQvcDQCyM
+un8y2v8NQUYnUe5LZ99m6F1m9LmXE+SpRoXn4h3I6+rKBeee5uiVfh0B6HxAX2xzR7tTRTI8jRq
Vlz8lsZ5FUAkjiaVV4Xs/eDxC/LZ2kBgWFLfZ3hOlknDoYVACRUVihd5n4BMPqdtBbbL1Iv0yL5G
MMS70XNjBGMXIFos2ExFeoWESQJzJEKW4lq8556mCkDreVwJJtH3CDHwBMMB7FnqglIia57IIHFu
IQ2ZxldPfpLBOfhAyVB2D1HaZGZx0qMIwOiKwImlf50xRj6/oddoGNzirbJHL5tId6zZLi5EXDCf
xEMdQpyEldAkrqpiyGR0qXPZFz40s/9LqfzGLRbfhyTtHfO5wZmqUL8V7vq8n3St01l/z30jj6m0
1Ax4q6E53Zr8AyhHqPuGlMVYb1sMA9XfMxeLEbw4QiD46ug3jMpz4DfIaFU8EkIQwSD83W1/VWnf
/Fi1wdhJzBRXUfK/f5qo1yXcUFzmzYrUFwlV2h3qhQ617vqhKIXhCva4322YMLZ4kfRmnYji7xEL
CO3uYjXDqf+wrYJnnUENK+yG8M4GtDJ5+DMeP6P5rHlxBkJ30xp+pZZDdf48PzE9BF1xk85j917e
4tnDNhtksBP1dwSXgTAFMCoBvYygw8eSxzCMKOERowqtjncRcQFuOwLsi+hXQ4AB09uYN4IdIMTi
4sWLodsq7AKY8pOYk9X3x17UEfBWJrT6AsD0vcZR6o6c7EWskWMwqYJtG+d/LLd7QhDcyW+zelGn
U9LEVzQEXf8/eptiwz0lE6cW7JVT2i+88cA/r63sUHmGvK8U8di+KL/J1gfeVfYBhGEV6ZafkPqG
R/GXKTpW6XTKWfxWgoDgWApmG32BrNlC9MT7urchOIiSUdphCL1dNUr39Guc0Nnp6rVD2xqKVeOF
KELT0MHa0hntBINwTy/wUw2OQMdqA892SBOZqWa9POfav+vjqOYFWCHPzwulZtFMEb6GHWZWCL6d
KtrKnmOJB3aXUsfoBzh7EnUnJtUiJp12kkp7kmaSGctanNuo09xogHbwm7L2RbgCUHTX+thgNjio
6PJ6PKf9fkbbF8/dqzpWqg5j/LidiSSXmF19rsdPtdF+dJaTQmQmK6jW/B7o6o7I1uJQmmei2cua
rNnCii4OiM6XX9SYCG6f1jHC04oAn4y+0E72jctjxWmL/2bcWfsa8UbMY/5v2ev8sAG8KYtMJf1c
mHaN/+7GxS6/7Zch6G6Y07q3CsW4+lnGZWQjC2ThiYXa6qpidMlm2jRDMmsENX1izTmdWEOr1hB4
NlWHoTVE12Th0/j+fYTI67R+/IbfgspWJBqlnu5hU0sgDy47fwB8gLFoyslRVNgc/V7QZIuZz8dH
cbvWGfzF5J8IFSxCcnzkBwg8SgymA+5CcRPnJLFx2uPW/i1vMg3+1qrX3o2/ZiB0rWsRr2HzkicY
s9NMgb/vp6ieq1Ib0QbabDRuN2raTE/ousqtG+k+xplNuqaa/QJXI06BwwRhTKlTiRKzdUhYIzIY
31V40/17/Yy7dXxvWeUuT9C4jeGpQYEkjl8o7c/lv35rexloHw7dUjpCGyKGXFpjixl1ne+1K+gf
ytJOnbZ/0A/y9h+fTvmOlNmB2Bl4P2nA1LLTaLBEqlRY/9YwVRxQO7GBRk/pJsR+O4eBQYzUUVYZ
HgHng9ipuxbiz92QmIGn/VTtBcdnzIuLAiP+W4/OmUUjEiCVcHh6/TGz2PV7Jjj4r00pWXgsg5cd
UaFD6t4ZsxIzEwQiBD0tk8HiaG2ajJv/JiqW2F04pMwPH4a7si6jn6xuT23fFFK+cvVRhSn8wLgn
mwq9QZxZEvHjl0fo7jRahGs4z0ZRofo/zALEO3AYd1JOsCzjDwC69gvh6BMbcbvFTO+2rhRvqYiQ
UAydDzS309GaZbDHT2xxDwecw2fNryd9LkZITgE9k6tkQsiPmuKAUgaHlOcweD+o+kqu/LonnE9T
94buUrjV0f66siEG6/ad/A8h20OovIYJ1ZbDW2ekgA35uu42n8lKtMPuwUw61v8u0KbX8AI1qMHJ
TvR0S/M/zUDEPQwj1sRsc46xEjkcGgg9KWTEcKlpipMnb2KLCo3ZTfAMB4EAYWyRhEieDb7b5VJh
IWo/VItHSpjwf/f5EDdwCZH8ukot6+aP1+podDrNElt8s0DiVoyxpfJfui2WmRX8IGmoifB3XtU2
sHJoqogAuD5lZqxn8ODiPOuTkKhdYejCze/hJgFauXDFR22OgW6jfNeqzg9VBVsviWncv7VA2fX3
PsfhSZDA8h7dem/hCwkWAWxcJXufEeHoFRlbGnX8AVHZqVH/27agq7K2CA/28p+Qm/8xRiDoa9lt
togQMvlCw5H/sXuBPEWHm8IPm6t/M8M+eKiGQleRIgUcJlA7rwvpWd3IKLVtxG8Q4t5Wio9GP92z
B0RuSHpqdv8YDjs1y9a4KhC4Bo9fZ7FchE69Sv7A3tPe16oDRAMJLtMaC10XXEyQA+66M6/AxN1E
GokWCaDtnoJ3Dt9KsG93AIXuc/lxbzEKrW4W7/9v4xj/PS3cGDI0f3oE/NSlNqfpblMrEsE/Ph+o
UxKW7D0k4OBq/G9z8+XS1qNQTQOafQTGAbh2WKk7OIDqlapEQpZQmEDR2LCtOOsInUKjNbyUID8e
WX7JsLTrPH8hbwCIHAOPdjNqbZhlC6CzPIdErl+qQ7CJLlZ3azO+Z+MX+Oz8oE7QA4QB77DFb3l0
oKf8c/7mhZUQbQxKFgfgOZOBaL5s61dH3f6NQ3OJQTk1KLU6PAk9EXnNCDTnHgNq/+T1R4LucGPh
XL9Wv2xGJMjmJe/HH8DF06TDrWEMMFvLUunybJIfzjhtGkN1SFd1B5+VyRQevVCpWWhoN6JXtqLz
f1jqWJTp9xV52y1DlzMT62cYFzRSUNbUSLeTIqTSCe48+N8fJkLhQsR3EHF41dwmuosApmY0otEG
G9XyDe18RbfogOU9VXLodv3bkyXSiCbyF/0YMTb+d6EiT5jZJRr718WqaEa64nvkiQPoBPgr0tBT
6ICzPeEXOR2oZUMSH78eh27H/p/k2hikO2R99Kxhpm1vlMe0G+dsCbeBNtdX955YKG0FPcUEgT3P
xpSa1rF40XRZe+wNNIX/SbuhsxRx/iKmYfK+v3w+Iu9LmUv9cOJr0hoAK0VwX+3kRmgHbKMt8F6g
40N8EpdWwIVy4NkRwyHipIZf0ZBXeGdevxkuEgDRZldWbqA/xvfdh4tGD5LTD+/vxPLnAqgCBrkO
X0Np8QfmBin3VLoWTLwuCmJ3FlQdpaksgnJyl2lo3IEK9H959vC9qeMukgd2u7qzKbY99ZjnH6TE
IdgtoQt/hMu96GHpjqP/XFs8dQLskKigJY3Do3UaqlUTYIn2t+GGC/yctnBjCnrKtG1YFMr1LpY4
TgKKRZKsMTDAKG5LvbAsMJqURngVfo8uorHHJKliy1y+w8kqfdZtU55WMiN8Xt2ZabyeIuvuc4kk
eV3Z6VQIuxXb1bQqPPBesggQG54UiJ3JRYiwUXj+lMG3EWuhvSPN9zv05jSYwmoV1SCM6HHRlrw9
AwmADCRF6kiCmVS/NzfzE55r8dXrVUamYmFxMJAfNt2ohxW2K9cQRUn8iqJFJZ11MJf6g0ZwW9OG
XkTdYos2SXfs4GyktYUdCWeBGCC1imfHXwmr325/Fkw3jswvqd1S9v6wlMJcO5/n2YuJJAVjxY6h
T0mybpY1QTJU6x/kxvLnk76urDN9XV4JmGsgWfJqNISVp9tUKDpY+lMMii2glZiQmT5A5s3uDk4Q
cr1QxtEbPuDvKJHxUurWjQPvkOBjkGu3rIHzSLLX/0uZ5y8yNzDEgVUzXxoY6PyZEsmUDH48UFl5
OsL3+Etze/fTgAQdOxWcRd7XGBWcRff0mo4Qr0QXt6HFjE04BMYwn00fWbgmv/xfhGq/bWVn+CVA
mwJlhw+BYFNOQCU1sOBJAue+ec62xKL4MAN4/4MjSoVDaqLew1Tug6WH+u9kDwdq3yMGsYx1Kse6
s6EDs1Q6jx0LyIGWvQk4SphgNaErw3j7/7hPIDF+C0xUUkpyLbHIkwXwR0XbzdE/0JdUwtD1wBMK
NcimXmBhegh/++yRRuB5BJZXdabsJqeHoRTlLM+xMEQUHkPMPELVNua3W9/eoRQjVSCkF9D9XBWn
lFSOpLfev0z6231OYe2gRCqCi8amD5IDvAPgEu1nlsKdaYOVmUSIA/fNDiFDbTBSNE51QpcLXnJy
MmKchA7EN9+Pz0/Da0JoutrIHfZ4O7qZ+Uu8mj93sKhG3xIGmxMfovdT8KnuxGn6VNbA2dtJKg32
/ynuCstxYeyHN/jCWswGxp5qGdoQSlLI8WE8FUAgWvHq5B2+zoQF34j+9ZjpiJDFblSbo6cRSJpD
T34wqILrW0L921b9mOLAfskjErxwa9vflOgSjCTZTiPq/gMbL0hAIxBEafENyvg9xJjE9WswsN5M
Rf1e6oFs0FUjzGOwrgiMEZ+S7pvDbNIT1DoTOTC6+B/EyxdR2gxUbAuGFA+RTq4nJXCjfhABhgPn
s9KRWX2djCEskAByyKc53q8L0cec0dbupfQkV9zc++LK7Tiu18nS39v+wd1fKbKbpkwuSIgMSNzA
4bqJVNpuuZqSxVSAwVMkNCEjwGsFuShb4+lnBDHCQ0LlD6uRQdtd4mjqfH2/KZcGfUYhVGmNqcev
mMcEROaFP8tawwcOHf3F3kwssGOJnDSHomXkf3B4B/hBl2Y+uwm27kO8p21JxHtCavHeLvPgsOAy
Jw1LR7An+oQt4GCgqyK89ld6dgvCO7zNBw0fyMd/S9me7Bj46meFXVFNdidOSFX2dRx8tPGsbHRR
2dse4iotMgQjPtJ5Exxvfl0ZHWT4dmJJ38CcoKF2Yc+L3pFMGoAMOY6HtVc3rzLeeY3cJP19l7Ks
e8rBm6tHPyAL9gbdIC9XOmKFCijhnimwPezvRK3u2CbEbifxIrBt1Fbe7mEg2GDEG1cBeqpdWrpR
2VIFdUF13ZVbZIxAQcDS39+MKOlSi4QHoCGTC7EuG1xJ7LovvCghBCzYVJIW+2ucE+qF6H/Tj7yx
ZeIOWHfiDT7curMSx5d/fntONFfTSY5WgI3fQZdf+HrePNtpWYCT6JRBCgqDH/Pro1pISyR9sopx
XNEOTzmSRC7HfrVyJHNumTNzqEaH4cuRktdkvY7/AXOYKoI0iaiZ0mdyE91Z5cZPJOWav8EsSqgt
BzB+LP9SrT/8fHHTRjGByHbDXS3/E1aK/PUlHSXkH+yOusvW+XeBa5iVuKNLwA2vK1UCzt1Gp0cX
hmmEAsYBKsI5mBqd34dY4wJh/qxvKKJCBNTmEVi2kVg1sXHmW0rMGvVO4b+8mvCwomiZ1vCpEsKz
cOBi44kj2l5rnXlZXgCwMgJ76LxwN76LvDLfhB/39fsX1U+rtoJ4SiwvvKiVqcTbm/R3mjrvEVyk
4ASpq+zBpxBZAc9UVmMkQT8Pbr62vXjrM221IC7xnHQPMT2xrJMLkKIwVZQxQxSANtDDWNCFw1AF
1teO/STisoQqAlo2li2GOw7c3OoSCEt95Sis7+AZOtMMf+gp59k0NY7tbcDFuKsdIoDHbEPz+5eq
F6ML+idzbRKiLo410M08aHeE8GnWNJLkqqx/WdBmg4wHePbcqLAcxIEmjHOQqMIXXZZbGf3AZpQC
W7AaAFsqLRwjzZzFJbOHQGcDzEKLFCM3zjmdWByW6UPTJvqtyT8loj7kgiXaENLm0axnslxEzmbo
mM3n6Ny3pmmh8oiTluDXxsDpOKvJbIyWEdkfhmWxdnGf4a016pJZIfmyYhiAR8yDl75LPP5sQ4Xc
08YvqX/IfkT0f9Dl1XMKxmbrNVcULVUDOB+ZPLkCPNf2EgfxQOb+VY4R6YWoIaxHYNgR8atSGQjr
4y3dDE0sjvlD4urHVPm1IA9AiqKNWd9lBvF1N7S5liNO67/XcxhPiHuxyyzlDVtY4pKOJxoHdlLE
zY+9H5eVQnMHwltSBiIKSp9YQoKdjyEqWs9XchweFJf4FNpxMuAvlEbzFvy+KpwpnCzPZsu/V94e
z9EVRZdJvuDxa2kWgCr/6sEX00KpxezCSndVNT5A5INUTbG4E6AaJfh/taer0nUWrLG9IlD7oLy9
kMC7HdVlBtjdXcM7Qm7hW+5YbVJCYZH0AMdIEcgzytv2gDef/ZQgy6QcdM6Uw8gamYuSoueuzp5G
+ktKV6tdWeITQsNzj2qkta3Gq1lqXKqGsnvO+40tvl645kiCCP52XHmhZ7CAzlZPxXjuzAvfENrm
f2pdXa8Af+LeLYjMPRWAClKApxJLKWjCYDOa5zdul1+sUDhc/E6mNiwSCwWLt+KU0cggMInKaCMq
ls/mt/rVYSWcSYUBFJB2w8xt4SNfX3E7MShSfeAD4VcnfB4dM2O7asQjRujksXJ5Bsqh1sm1THdV
6Ik+0o/31Y8/+Q/xrJSw/ew7JX0khfByYWN4i95Vk43fDI4+aiYxB2BTqS81jh5hbVNTGvkg2Iqo
jG41AbGAtTYTWeNkpncY1Rx8NUMf/wBoAvR/2z2QMhKnYUmoWxcT6vZTMc93Jq23DrXaHjmxKtbV
eC8xxipnv5ZQHpYeF2psiV7cg1Vhufo4QAfE1PL5wfewp/9ZuvHqZBMQL0Sh+aTFAQM5iISpOKKr
5DBO0ayZkpuY2owyb0dVPdo4mib41irdROag79ac8YdxQYoyRJ4MPhRdBPk6m9Q9zYVbVMAWINsr
ZMj/ZhlejViREjXS8k4quv8RYncPcgOPB7wkTV+tJk9G/cQFpC1EDTJFKqrQqAv2amMPdZxvOKBM
zon5QbQgYqhgRq/8LdwddSY8L/bBDVzx1x1IIB509bno/oj6L9nr1fUIhhnXrK534/DGWRTs9O2m
YtuwE+TuvAaW/5nCqvTrmUrMUhDDu/KBZ58tuCk7uS7KOUqvjqw5hkUPVDFL5EKH0Krk7jsoo+8v
kFwDEC6BSAL5orzEt7069xzWNHQ2mr8vdozvRoDcOz+xv3/GlutoJ0uxlrW0AZa1gntLG0LhTL4C
rm+W29xk2IB10VOSWf0/pRrnKhn0/EplAOmOd3o0zMR4jc0jWsLlwN7pdX4O7J2tzOAUGuGMLbFH
ty1L57AW+iM+L0WyE+KY5YHRralXHmsa3dezB2hYEVFBVE4+iRj2iUahh5F2z1Bth8HBH+LZUYpF
q/owoXMtA271cJmqrDRmye9Q31fUHMJc59gYp0xGENtfaurhCSZT6RfzuSW/UGaQeOyh0M/GW3qD
SCZlUdHHwKMnK+qUjisazSd2HmU3Z3SDQUO71ghz6dACnvNrslvA/OJuM6GYzo/Qrere1Uig+xIE
4IFa58B3n6Pnr/3AoNEbT3avuMwFRVARNBpQIZwouDjUZ5n0yMcgUqkU47xJvWvJQjPabU3+0yp6
tPio3cBfwKBjq3h9SABpzLAzH2y/0rbPUvRolkYHm87FM7VXNnVonmBSsS+hsSyHzRWHWd/tmYp7
Ig1SEydpiRQavQFowjI0WbxM/YCo7TIC14oTYDYycQLNoKEGbkbEuXuy1V5s3jrwxRWeThqEpCFA
T5mvyzlJmk3PN6E3vUKH2lk9/8oPz5YROyxNVWsesXEzEVxbd7YJkf6572WbjnVvWPeRhgRyyDcB
IhVtEGtGwkkKkJ7+50CrtV4OPiWnPF56/W4WrHIjI5IbgxNiAv2dbIodC4n6uolG8UjvEPgZTkWI
VdXrIbKPYLrBAWtDyIpdQgvoIlyPVODdmskAiTH0O3I5PbF+/EtujnIqqwzSekL+injGLyyNj9SI
bi+LOJ7GnxjiW3FbbUy86ZQKFD4aD5f95oag4C2eB+kfx76VGV6sXxYThPxJxELhCnj5kGQnf2Lr
IfCr7BGupEwPPzrIKoeYaaYvYLSGrXX8cLmTtMuL5kfEBvcpSPSajHHikzVzzpUIXi+2pxGyujMU
dzSypzX8JW6kxOhEJKxHUZrlhpdO3Nr0Ll2/aB3+AmrhJRkDdGEhab4AAvxcjjeOq7zWh/1knb7J
yJSCbaSZry1Vfr+Pj1JOHbLxpnQQ513SIznkDsws+XW3ynwnr70/hDmQUuPVsNiNUXQo03JchOuY
b9WlJFhJi6xesfw4CmgrOuXm+3ZECt4GHeogfku+AcAgX6/7UtQqBE0wVwucmRkH8VPKkMKNIR2A
Xd9DWDd/Gkhh0QUewTkaaipmHKxIVbBmrIya9/NrOdTjTC1pQz0xUTJBNI1VWzVKoQLu2y6dvIRx
948xEo/GZyRICbMw0sXWW4jSUdquSeQiOOXBJonPfFESD4Q036TyxjPYpql0oMgq+IwD3up3syQM
rIg+NswzCn4rYFGOhLbEj9sEOiCSLzKGgCfOEZaEtw3bBSZcHgYAmibV2sGnFGOBqJ3U1sxocRE0
WrHS3C3t9EIlHvpTTneiLnoyrf6msX4jMpJHlk+ELqMaIAGF7oVXdW3sUTFcIdhp8R7heq21rOn+
4Lm+Q/LM1W7+VkluFEy6K0EAxOQ6g2ppdHT8pf4qgSOKl9mgzEhAjPJ3tMOCpLa2qGmRLuNZBcZg
EDkjLXArJ2xqyfGFULBFO7LAXUY9bQ5pDCONKYkTS9vjSK8U5yHHl0ksa7NGAs/0FpiSpsnqA9wi
nu9smPO+Y6Kzptzj4WZQN4Qh0O5vNI2SMJCHc8kY5Kvy3qTNhknOGbGZugKOH1BlE54lE+hTwbaA
Da5U3726RNI2mIJutE63EsHp5u4D+Qg8BkfmlQY0Tnivyegerj1+HsQ0TXf2m3rpVFCV21XPSfPN
JqC/65RttRzJepy8uP9mzwzYqpU+OWUo9cmlKrtRv7fNDMonKXeNkWJPlcTV8ci/f9DaDBC2fGTz
Ete3Zh7HDhTIePGg2dHh7bbmYSDLow13N0rm9fP/P9c1+l+ak3CdanX4ycwXhLUF7RX40p0jNt4v
DgwVxqnfD/AHAeDd/CzohluR/b/4em1IFZjyBXbUvThn69aL9NYK5IsNTdfVveOp4KctEtogT7Y5
25kmMpMZc7bhJXWR10lzRaJ8kWJeLZBagV6rfzLUys/yo54X36ZCL+tV2A0RPUisXzdQzJyJ4LSY
BL72LoPDtLNPC8QXGcO3VZQgN0tOUdC1XCaS8hjuHOzWIqkhbDrwsQe84EyX2skrp/APzgD7EXlo
0/VNB5xy0YTiO52Q+C81mInd8Df+959S9ijrT7bnvzHfDZ999vLMCIOeXUGUahimFcTs1y4RiOna
po1ckukI0qn4ISMAQkccCdo62BdpSijVqaQ/1S3PYWa4vurB2WFFFGQjxJIoB3Q7rI74zcYbyK4t
9ceWIwe13kwidesGsUVeMa0Ws7lw5JEP9ePIjWu5ZkY9XZ5OPm2XaLib1kjruT8IzE3tdlGOMyNj
aH7KBLc6fsfAjO85qFHvA0H8U5ZIUSBbbb5qkkPK775a0FrtStFXHkzt0J1595bxPFR9TacnMrpJ
VvOJzTqX2DSh7cphwRdqLy9XsXA3yspXY/aiQ0dRf26oxdI1EP0powWrtuTKLtZW34hF2xpIOuta
/bvz0HITpFwnPL93ctiDcCswOlOzhYCjFH6X4EcDDTr0u7EVa7G2v3qUZS6BT7CdiyDW0hEt+Kdy
DirBVrhsqXfkeYmM836ErVp9oWRoHVj20uMBbjbElKILWS/vTvToVQ630f8Bvzp2MZgvMSXLZgtX
uHxuo4lamWRb7BfTX5jQPuERGPVeeTbD8eujIUO9hyPBl6QcOBLOu61DO5b3L+3EghmxvccsuzHG
hztqTyYgasS8p/9MlAYgWnvYy3O2Zfh2Ch0pHTit3zNURXbTG3pwtCploiT64W8Kcf/ohIh1Mk6s
6IAXpHClnp/dlMb/V41Aelqu5JbtRLO00pCAcHg3G1w6MBvPFw0GAenHnVIkjgEbXLsnofofnKOr
Ooe98ocVV51VwzzJ+/Zs4FneTUs7luedPEFAi/cOiA2OZCjoIwbvzdDVxdd9QY9fgaRqQmaOiQOw
hez9jpzF+KmmddD34PraPWYcZ4WMSGLx96tC4DXkU5WJGZia4uoQxe77RARxLtsMc+rl8vcJSi2M
Pe4+XV2lv0ayAUe3qpwnBZG7pmaWlczHUOk7By0Sf+LzaV+BtmYqQWR1H0Y36pLnENylm99juwGW
3ecqifEefAAQLCVoLWVEXPx+uUeBT2DG+Ow2J+l2ASyv+pju/13niozPuyRpLJeuOQwVwLi2w9wH
Oi2H2Wyk61r2gLC3ixI3ccbW8CqZCH2M21uVbQN2PTCeBSWUFeUlqnJefpcKaNOdQxwhTmtzxKP1
e2OvRmwhRlsf3dn2iSa/rUyamA8Qghd8DGd5z4aMsei0J5mrHmoedb7ufiiImYyK3y+7Hr8J2KHp
UYnzFlZbRqIVVqWxmcOVHpiJxR0QJKh6An5z1ZDqYOyAjiYKu8b8jNR3ngo5BTcGsUZJW2msiotx
7nL6HXRY29TGmN2cGvbl4jlVDtOMaMm2ZO7adWnADM/f3dBr03wLLqiInWeXbQH516J9FUSRBx/E
DVrUskRRpudboWy82AmEKetgkz5sk9imTBwKMy32OAIeDueo2LnKC8SDJNv011xk75eW8hyfF/J8
TRo0SVZRhMlT2WRxQA67Kdd3jRaYKgZQkZjsjeUioH18FWCEKccn4xPsqKNJJagsvmbXrYTUw7ZL
HLTk4f4aJeuxMBEwa4h6XLyi5aWNPIqCs6Iod6r5+iMo7SCQEYB+TzOJLGRopEU8bBntMnNgjwwM
dh5ptN0h2ss5Y1dBC5Kzbe+mUK8Z4lvzH/czuEd76UGJy4kPitb/36oddyBgetYtYqL1MQUnQ42h
nJMZyO7OL2Snj0IADkG1Ofhfy7mz7gZc592YCcE/Pn2d76NRmwSNPS2d4K1TJ51oTSK0FukakVle
8sRmEasUPJYZ45kZpcaVzAnitH4GI/TYUKWLrIxdf4HMZrc2xOj/El4ZlbwrlBnpT1FJZFH2Ck34
oRRVeKl5TT6h7CIpO8lZtgp6L/iFHqII2AZLf8o1gVjHq42I3V1BmARthP5k5gt7lmUY3YqlC/vR
XLlUEt7JsAFMPdX9URv7wTooFZ+DRI5jbO3qdnm3ZvvS+sZo4+BHU4muQciK6VCFrBI2DG8YUJzk
F88BjRgTM8M+zS1DE55kYVlHbRK7D2ODzzLga3lOndOFAn6X01jKpM+KjKYjKl74U+TLrs3NLBWH
/emKMvQckUIQZ0Tr5xSE/t/rbbUSuzxJoXfn3LDiSVV73X1icOumolIWxZtTFVqzpWniSmT/w9Rf
h8c8kiQSu+8s5Yq+skL69ohmQuBfnR4aVGDd77D9whq//9slwFB0HICagDTeaw1AyfLIQc9U+FlN
vEpcBhwD+SdjNRGVIuu8a9O/DE6gCosbZDrT0gypKY7Iyo/Yz3VTxAxFOt9/mAIp9RFABUY2DDX4
DwNr+7iWIQcFHVQKf7yMOIl1X6RzmEZ6W0MHCYM9VieKYYpgSKgmtn3n8FJ3oysKskScmKMdrjq6
HA7ijhfZasLUnQpy3tfNNTEoqj9/KqIQdRlv7yjqgRbNAaE5pgW2fShV7IaB5JSlPeVoYTJRfeXs
3iPWbPKyeY03ks91iyWY80rGfmFvVuLWe6X4Rea04Vk1C7a4kZa4DlECPjrSuabZcqJUl9dECxKM
Z1vm44YZ7FSAe8aUkEwJns8WPZBHwPLvdJRYCv3b2nJG3o9UcVob5XbIlZseDFZW1XEX5RwGBbsM
EqdNQf8kUdkFMKVjWNdL/YB0BO1gO9OkqbRMCP8DgLXok030+bYPp2zLF5Z/OKeihN7U+XyDVEqu
DDM+6KCa2z8NhGtQrgv0m8Y9zA5HyXWUTNTaID1lE3TPDRf5oqHGJtXtJi4zR17iziU6n2ApPre7
uIUnPVEZtlmYJwE62vQOOX84tQAz4K/cyYkaXFOWLHXRGyTFJ21L0w+n0SZVYXpLykpJCNreYMZ7
ujPAYqjIOh8qJmQ8jhJn4tViejbjM3tHYYpwRQaCS4tOtLwD3b5mkr+6Am2aMDjrckylEa/WbI4K
fdjV9rISziPwTs7DPjnnaZaueCQ6k+K69pFRspn323BMfpDNIqCNIZYmdfRFbVQy2Dhr/vMxdvzu
8a7Cp9m6sCFD/po6SHjnk6XvozjKIgi0yalmAKaPK6FqKSkPnrKqnRNp4/gp/XwvdT1M4i5wOPL2
Mf83eALmaEMHLXe3bbHfkD/vlbwOx7ybxQ/iaO6InTtU2Xt3yHeUm4BIJgO53Ld8ps+xeCEPIxfr
Q+p70KrOxW0piWaUO5KDq6iVb2KoV2ALoEFAiVKQ1AGHA4GMLYQnw6gtgLC0uXvwPpiRdhyKF8Tx
0m+zXVZhWMVf28s9Ueut4zk5LuirTy5HVevjdEnfwGDhwpLtPSXOb6JuWwScg0qgitxD6lj8nKVu
TAkn2/0b8hswdLzV5n/RzAcLX7X1X8kro9OvsS9K70GGhbHnFvkRPtWeSaG2X+7pBJcKQPGIm4h/
yDXMH87WHSiwCLLLh0b+3U7Pkdg0wbwR27DweFf+mIBh77PMjpn8ObU3YoPm8ZVQ0qsKcAo/Q85Z
jlT+cdQR18RS+zoHmPLw9sqVqf16KHGbPVAZNktWnvSoeNfzlzKElKMAdYY/LruRVXlXzEOOvnLE
jvinj/NP32lZBknSx/3qdk94gn3HHD+sXObnZk7EWYnaeiuBpqMJJWAnhE7xLVrsGc3aEYWKxmbW
fq6Wh7B62370CDbnwv19l4wOPEnkiE96gZWNFswmrulsUisq+VXwnSwH/t46oY3bMqe0jv/fDP0s
g1LtPvd8nRk+UDwpBKf1ivO9Pz7/DhwRroo0t1icIJ8RJWlw3XBDIKe2EX2t9Fyo5GwYfI4zwj0T
36vLS5B1ZlKQB4zDJLsn7B5Nz5helnXQsd6E31OV8Rm94rO/B5L5WCj86pZ4Ej/s6K8995HqHGvj
mEhQgteZyOsGpcredVbFgJL/DQSEcWnersi224TFayfdGSMyniexz8rnA9HduuYXCZyAlNE0QZrw
PEuHZTVXNoOst7NyyejvLMQS4FVjjzK1z0ofULo3taOm5sdTyhvfovwXKG2RvelpXrC0qYXyvdn6
I0Rglu5szWRc/QEH3nkCkxUq6njpdq81TcoN+3lsWyXveD9XmFKADlO2WzmCRhmxxVryOzCeFlv9
k2OL96q8oPHdEytytTT4Nu7yuzP+U6VqL1eHAdVf6QEarQw9R/fn60k46AciPGWTP/yv4LskDInM
67YA3Qt1msflCzCbbgIFlJdTdwNuJwRV7mxforGPPWy9TbRPfCZquG80xIXJrk0OnZxS+rD08o2T
P4al7aL2CDWL7fYcTdI8xOOlkyW1GXJaUidHzEvWNvjU/LAXPbC5EqDGeKjcTVbRUMOhU74zMEiW
iUj2kSVVJHYhq4L/F1saIPeH66i90IUzUSQ/C9WIesc8tH/TNd+JbygFzDFsEKKSTLPGqLxOXdyF
uAw8FkDRfsA4yv3D2GrQKuCyWm0RbqQ7gfFc/DlHUx3/fwsoHMLRuvicPV3+sHUZFlP0RoCutER3
EzD/9hgnSbKfvAnUEwtEGQ7sc/GjQYvTzqbSwLGh7B45xvaDwAb7h/qqCrLMlhJBIT2XOd2+O9dB
AByVZA27y4eZJGEy7jt/Tw9VKh2qZ0If/8T2unvXaqyQO/uouMOYsnB/oa/FdmFh/O5SkPMO9uwm
U9ks0n8iSAq1I/mrwJW+YFuozifPVU9FW53rRj3S3T4kIfnfPiNizhFr6nP6fUrdIyf+eGODW2iX
+r5dxhh/BJdC0BuP1peLyzVquFNVDms08eJ4nY1u8xWtivkbTcMdrCCyKQ4+PNkELhMdMJIzOq6t
UH1fJAy4PUj16+gOIUo+ePRzK9hBCar3wF8DedYTTk+dD5WD7le9gI0+OcBkYgTYXqmG/QUwlR57
rQReCh11Bt/xYRP8RLB/OOjPgoV0k46sbKcplHZkNOzEOEP+M1p2NqaeXAZoPDqrLIdtTOvdKLXO
bQgeJawaMmI18Aa3YO2FLnBZ4925qD9+oxDm7Qox1ErNm9dKQDqDUOLxoenZYCT2Mkq78gx1+AzV
M958c4YAVDUM8u9DO0Ca9wo2wq2SEWBTLocafGHw+rqP5Bx9+cH5AqC/PF7ccaZ+5V29VQTWAMiA
oF9Zf+2r+G4TeXhaLnooa31fqJ8datWSNOLnt1swaoqK8Swda9SVb15/BkTPPeYfDGQXUl/Q2TL3
atQz9iIre5yszdsU5cIZIyECODIdcS3JB3RAivPTGw+aKZJ1OBJjTUW/Kw1tdykmJYHil96wQOHW
k6E+IX/2CwJs4cjR2cK/aK9EUDBL3f5YzPc6f3w49qO2zbGPw7Vdh5zsqIcQAtQthuaK3NeBW3oE
3/d3qh7IJ+ue2dCKer8I2tEuoDGH2b37iX3cHELdpPf1q2+i6XBxOuLNna0C0h080YBG8KXsKH/A
Lzk5eAdUgg10niZ7L4ZzCJmsjHVud91DU8pYF6l3bSALUR07QZZXWQ0R1fs+Zj6IVJNqnqShOoKI
QK84giWIouHl8qrR0gqy2Rgo2aGQny6uGZSHWLScaW0RoTRf7A6KtYVTRGvhqA6pyez8E3cdAT7u
1Ynl/KG9dTbEDJAU8zzFqBxcbXrJPNee4HfEg+ZUiyDXB0g8SvclhBKp4Q2bWw3PPtU2Fd/R7ngp
zxwccl94I7+YOS3zIKIIPUkUsGigZ24IJqnMXg4kKkqXswL+074mItw4WTIcEvrKP2+JzXgl8O3/
TVmpGep+q9OxW1fBqGflmSXM0GQW2zoh1l9c+Ln7Ae2Ixg/636PgI7mk0kztS59QmIM+jx8O4lQi
Q8LHvWDcUu8iM/8M70Oa5eIswY3KRRft/UpkMk92LQ/1jJvyp/x6DJq2heNGqtXkklqTpO1HCmce
6twSA/tLwouVWU+C8cxCitUiovx4izOgL5K0Z3S6AKcnjl+mCKXHhSECurbepfWM/TtvY90WgKwe
HgpcQTPzmAfLPYDEqmxrg80LPVJNmtti9YS81qGvyFiIwwUcyo95kgsO4QdkDdhsCgvAvP+rSOCx
ucpa5FmV3OZivGUsadDHzgD7CUd6DGy9Mt8qo+9SDW7YhH2zcjSiKzvqqtiQOh7oSHwaeiZL8no9
4qGQ5WoE1/u03ryEIuC9+4jOMvjd7bTP1yquIOZSWrRCsS6o4j21X6pZURYQ23zzOknt7W583IO7
U4VVo7vXOTOQ2MqQSeiMLamqRzlTKnJAKza/129W0v7ITawLEnXkVbd4JCRBoTRDjr8Gd8FgnXJ9
wBeGeO88fj5CfNcb8XGGySZZPJGd1t0WqflrPoqgNi7nyxfU4IYG/wVx32K35CeLq/4HEKCj3/wp
cNCMs5gkPF/gzm7+I5fc/4onDQ7Wk137T44PZKYtoXMW6k5arCFzVca3l3Si4gJ9RaFB/HDJC7rG
rZjRpzTls2o/YT3AYN+71uObdJlhut9l0I3fdXcCW1kHHvQrhqYF8ZHziPTkMd2FKzUXt9mBlDUB
WdlHoRe2D1A9EqGaabh52WKN+SvR9nYbaAOgoJTYHR1MkcosLFHHXr0zBc7FA/O6pK/J5T+CWwkA
5swXhgr80htHZ0w+tPjbyAuQeGbuPrKSt8LSnFaQeCb6NgCe/XvPD/Pa7mbNytIZb06zGvGa6xT+
JUvgIEoA1iJY/43z3vdDEq51E34/5kA2LrkOnnuara7Qj5BSAwYNZB8mAOVymBLbgtEj9g5Vwa7w
5vKHpZGtHAK/vquE8wCRQ7yg0BP6919F9cC89vFnwFeLO1SC30mghWfjm9mZq/Ofs/5U9CEobNt6
bsehZX2v4JC7bauwOamTxD+6e6K8r5aup+I0aE+bDcUracMh8YN2myfNw+CKZ1WIrwUwf0xJiEO7
RYapkpaivXwmuG5mHeKATRgD/Fi4zp0+2WlL6Pd0cuk+qPBqvARVM04qrDQ3s1rsD/uRtwGZxT3C
M4+aRbxzkVMoIB9bPtAMweNljv/zTfMTNndbOukYyu8KSUcT+ji1zBdJIgkGOlPp0mhnFIZ9KX9F
nns/1aQSdE6540wdYAAOejmi1ZWHg/eSkWANGif9jNz1tXiyd4kAaQfkAfypwhWu7bKXEyB20nTR
PEEQVyRjqVKKXjpz64LY1GBNj+j37Uf6PfxDqsebtAczyE37aNTe4NpVbeefRmFtyKKCfp/leK/q
ia3jCR6RZtntqmImfTzZGk4jcOYBQpHZLhCQeKdJskkhkwXC2+pB972gjtT9SgyH7JIuX87CBPep
2jihyQe4Sj78ZkkCfnj6OckFVvyY+0yPIbUJeL2I26IjHRqOq2GxRm3zIHbtlk9MKUtkzuq5gSU/
+Xk5TrIOhQZnA/P/yd+7JMBYWjL/0vp527xfKpDQtdQ3I+zDsD2FUTxM7bhdM8nUFk30bOve5fDp
vGxqbJP370xPFk+X4A2noWs3bXy5R5jlgzfbdyOD2wFqSPW5Nb370V0ivTEQfuVXvracvzMVD4vV
tnAV+8Z2UIAIP4rZmEH8+jPEMsgodrFsGwW4ryRq/yLC/Pk1eDO6oEnVd485noTgO3NVsKbEgFs0
7gdmjm1/WC0MizVC8ccFHA0Xs9ZwR806et1N7nc3btTzGv+ugwm26GKpQ4R5zPigO31AUMftVjBL
NKwk8duarAct1dBr5pYYGdmCyeO34UuefX6qRudqosYpvDst6PS4j0Eak9M9PAcXuAu5t4L0p3Rf
y5tIhiHuK6m4qHHXks0ZKU70NLgfYMp/6z2++Dvn+8uwTKApQWqoXtJo6tIvEJbqh/Z6vwe8Es4r
DGsrkv1shYnL2OyBTrkCZArMlOOetDWOHGEn5lSRoMz40JS7/hktE3R9d8XOrbJFR/dzVZOgpDNa
OZut7KE8Up8LdrnGlRWZpCu6z91l6qEEyGtV2E1JVN5wVIhC8+DJnUn7TYh6I9y9ZFhZtbSIV3Nm
sNp5ejk4EnO1U1c1ReXYW1bFncl/tt45QuTEOI7SH9H8Me3c1y1WOZfsdadvijaUdDGRGTHIsqb6
JWIW26hpB7sG7f1hoE/onwSbXxMLYuM1gwo75+wTb3SY2+cuRjuXDvXh/qYfwY59ifXm254rcRKk
DCOx01XDKVDq8J8I+2eACY4lL80HoKCCfdiUyx6N8EniegJAM1FmWLzbkYw6a9ZtNZeWn8brnL8Q
cnmPGcxuBlwCjeg+N6QlM7ZQjiMvMCE///5LF/SATf3T10Sd/WpoWM1EPXDmYTd0OkEV/S81rfPc
hg7PqiVCDZ1ZbY/Qx6yZHPc4KkxsTI+hJhhbH6cBE5Guxdyi+6wTTRsyrVQuxurd7HzLjYXLPX6Z
+zrujzRfZV0jGBKxk8LZTQEeeP2cH62QCwRIqnNSwbwriUBBz+WeavjH4bycOzh/XVqXUgT8xmnb
gm8vWxrZFFng18dScyrrd9dQbK6PU6qVMr0/fKPdAopGkSglyLf1WEqgqXyqwEHH3eMLMXFWPT70
B+nwcr4IanDw/LCCLtkyl5Bka3kueRqkRxVoTRbbLrBypuCkDa5MT155p3mkIdfAsfIn/ML29bKo
Rx+xImYbVn2YrYT28fKzJMdxGe5nSX8RjSDp2E4f2fque9pennHJdHKF42jSIiWtQw4lvtR5SCaG
0LwEcLid0fEfwMHTc1pXFYQEOPqK27oex3rP0O87AQHoR3Kiqz9bogEHc7qz3oe4WPmVOnNcJte2
gZjn+uWd73SZ4u6MCq9U+1mO4H9XOsBuMvo76hlpKNbbF4xjlfuXfEvxyTWvUPwgWpZe0ZZAOV3t
R1hgQns1H2Qu0CZG4q5yQBEBVFgqD0mCPTz+NBmbaZ2yKyWyjyZwTXp0PoycwetdAL/1I6+WHd3K
r1G2gecK8+u4IdsZm7Vqo5d2DeI+39vlYA4akMEdsnCWoOUdCWihFAhzHCvWBoOgm++LagEjxG0Z
RVrZ0HFEiHACXVwhXRKP7BwSRLRmD8V7kqDZvMib3JIUX64D3V89Umt3kH3fSRtIONkrsVmU93iz
KSyDCa3Xxw8bElg0N1PxRIPWCeirbKuOcf1i59L1HBJBgJmDDii56c0xsN0En0VOZnZHrpOhl77Z
pcVDspztVFoeImV6YPehxGZz37fEsw05MzLavtpnlqCjBs8ALKLwJOB+EG1cxnD0FEeQwC8xLGAa
OvwAddl0hx1aeu4cRavptqwrNNPQ/KaF6igUU23cYxLIyDLWMqBUBpNuwvnmCpFXTyGbmswNKkkq
XUVd6xWfDpHm6UWAX130n9/V1EnCrhnSY29ef2AIXAaTCt0IvQ0potab+Cb2zqcTm1mkNrGWsuDm
kBkus4hmdQFEQfM4ebyi72dyHPNxk/6Qa5uYPjDze1hTefibBDrUvZJEuZAH+UKJUM1tMIZZiJIN
E+d1MKtIbxPgXkajL63Q8PdQgWR4bGl4F93uKcHA3pZj5hQiAb+mrIG0gKDi3PBqcM0GDpT9DUXQ
uULBqBFy6hwuQeVPpv55H7Nej3645DFIMDfrmhK7f67jaX+oihjdg3UVS5zuyvqIKv9b6tfVHNc1
GplwK2tQwQ5wlhsSoFowG2s50hlsxXYW1HRZuqC1JoL4xSQ7c1y4JcDQhIh05MvOEx54DB54EI0V
Z2BKRTGN31GrwpDDkx0Q6j43Z9d7yua6sYt6WMIs6EzUSZNCPVf/Pkxu4NktXkltQbrqMTe8hNys
v1noJSksLuXJV+H5+bOYIr3Ep8JcTs85HPiGSquSSHBNodzL4Qm3PjfFF2pfiUKj0c/B+ZKD7I+X
jNsl1O1x0BzAtn/Amqn67KFazdDHbYpPH86iUQPbuWyOxSuyBphYgWGpzcgLvOwMou636hqgeoiW
aJAoUY5mxuc6rTgiyGxBpfaN0GYN0fHrQOZD3Nf2gFIS5/4mSOu3SGg29BVnDwQbwTI2i1bzLG2f
dl0+KzTeYSFgkkVdSJefPNXOEpxkLn5TXTPPBpi8i4NbBP9UK7PsWH0P19E8YbHb6h9MED0ByW19
A3PCPvQvkrQkMevB2P1gR304Z9XY/3B1MSVihFudzDQ/I/DlUPXrOU1UcC08X3Jm0uym/zNxvtrR
cOHGJYmcGKNctAZ45Kv8M9CsCOV3HPfF9fNrOwbt4NmFbUsRgJ6xhQQW7zkruQgbtwDlP3muVQ7P
F4I5ZTPxsUIPNAVQLK0omN7Nocpmot59DOgRPS5VG+AN6GnRh1EVMueWzOPivfvBvbq3YtA7WR3+
ONlmhnfLIeTUdarUVRJrp7OHOjCTgwLfVgCH79hoioNfUhnTzRmQW4Ls6dAnoX5dRXGxMzyx8M03
lmfe1COVYB0amjl5+5mrqr7Jf84eXp7f+elNeWpW9Ma8nEYsbz/xjGhYVVY/bGXfm1SIQaX8/bJQ
DjNCLu/D0uMbbG+t2/K9KCZuOAJBYOtXK7MXRHB4ftFTS/tEX4NFL0DcdD4zKu8qH87fSq+60B3o
WW5g2ykcg193dQVxlqpTmHfOMetQy+3EEw6nFnJuJT+44Z38GTI8l4KQMc3OeS2s8gg2kJGvtQCt
cmK/lyATdOaQ+wI8RgcivWsfSy0k+vQuTp5M2XHqqpc6fFFvsrwsP3n11x8r4zC3E8ne/x5yX7jF
u9ro6VYsjjvT7HG/QuRWDO+qQcynqHXDd/R0PkMI/h+UHZ/cfWNWb1adkEJCbeCq+zcF2G5uhbaB
OlciquPbcw0upZFJrKuyvDHpMR1bOPCfADWkeRt/Ie4AF+lKlYC2SLs6EPAeLN57hAxCVy15SciC
+wgsC77hiy+hhsCiTL6YqwDf7xAKcHQJA3z3iJuQpO0kyG426hddfQvJAKMgM/NzmDnQjF0ovBwS
8sr5AiBZjlqCNpLc1GZBWlJobN1y9UL6ROFtGqpd0nFbqa3qc733stqB/fYPAJR9MLoavjhJZrWe
yuq7d+LlPdlwGwq6+0r4KE8kQ/Y4od+DuW8mwh2R2GOL8z0u4w0dhWB4zNzl0NdPKFJ2SMWxpNfb
W6yMMGKViSFuJFkUdGNLx7YlHWIy8LBG9yWANjVDLJ6wcQGrkqcGy1habnhKfxlndj0zGUPbAjps
CegG+H87HDLyy07+lC0bnBPihUr72xNLvt7Or5lqdKeRVWw8BEnwZa2CoD7ZTSUkO7gmf00YL9NV
SgAEsp5SYVy0Iqfhj07TIkxTJSNZg2uIwQYUNTS7hpVPnT+/O3R/gkpN1HGzpK+2tD8qGfgC6tpv
8cfu7b/5i4Irl6Ms3Noo95dZQf1ioHTtwuuls1tW1lFTUXgamu8rAvYUW4gUWrRsLtVScrOVOEIf
UBcjHYrqV3uMQOSLnlZi8YxmRKFSb1jkD2coEnNYYYD03vzD+Z5b4isHW/LttzNmHFLxFGQneSrX
RIqzAG/2PwD5pp5QaRUBe36YSPabj6VrpMMAeG4TYZ1ZAfwkoJfse+IPTHu8On9z/sBIkoWfMgcU
MWpKtw4b2TSyAjqQ/Ft3ed53GKRHp4KVrQxw758GTxit6rHhWd/AKEdpNzUOERFvkg91ypWcj6el
lmCla5PrgXhJ7uibFNeNZNgY7s3Uv2kY8UgNIgiL7KL9PZjEj54BiMSNTfpR20mi5+dExaeyHeb8
5ENuiNmtkCRj1uVLGIpevH+0M0cl2r3xQqWhTWISf+v9pjBdkqoMHX5n0laMjLBNkQfsDWkDdB1l
ckStaBX08Q7CUODp/n9vujdXbTMZ3qwCjwGCwB7oii7hutoEwNwdUdYs2FkJvObX+C6XGZsCR0cr
WPnT2S4tGLPNYhpKKJj5LlE/u51/n688zj31dCPR8lJzHLMAfgtXCWM3Z82I/N7/3k79R/9IqWKp
tMPiRvlThgV2Y5DrKedD0LdHQrOi8dYqgrGwf8xZ9sCt+rp1Rn8qmlQa67+7TcFC24v64KJpv+Tu
M2fsRrtnftTL7rsiM9ol2FlhU6q0wvEfwYpvn7Z+NJMFgPykOyW2vmFvzOL4vCPwcliHkNGrrGnv
r8mc1EIkAMFgLBDiWkQr/u5FRiZrxGNAxtvf9Ut8w9hto9S5QqFdHfqbIQPCwywmCO5/66yCxZ4W
YzxLQ/WurRnafgtbujS8vugA2TWZDrF5Be41PXikkDNvxiMNYg8GsoXehPlqUc3b7BjwG+SxsR6I
A6SEm1X+XhH/wfORXuyC3zu7FSOep/1fCj4PqEdkF944A0DSV6zDxVwlsVvaFT2QY2huO4mni+jH
YF3Ei7cFzrXNrbS/bE/1rJcdh0dIJPmSFIE9JRgLxWH+jBow15B5zFID72/Y8LvFaYWNSEefquMp
VgvspAU/ybElZRiRiWwKBvdmDLHrV+SpLKcvSnDKvvZhtEvY3irVhGy4fIt5GOVrvLMUp2wcWz2s
06+JA2PrRkMlrlYzTkW0HvEGySZEKuYOkUYmisntA7WjApFK5ppGk3FMuSBeLMnvRHAbf2Xws0Ok
Xlpj//BfA9uJ63V5LnEIUCc8go8GFlXiYz9oI/ncho+tkETlfI6OMsoJe7Rqu/M75UULZW8NhCOK
F5ql1VgTiUQIolji47QTyYYK9bp8S5kiYLrjWz5cCvkjYlxlw5zCnRJAZOBiu2Wk3O27vXCohKWy
W9DDQIPFRrSgnN+ZsgmR2PvYawT1JjNdeX0xZ8AbF6g7rZ0srr5bELF/cgKLsnr+dtlLf4Ooxr7X
X2zjs2xeKLObHj4LHua+vOEvNcOuei5yzlG6e3NjZjMC9stL/ZpIBBexJGSioqMRmW3/H8cUY6fS
bRemVrersjtL7ZUDBk79+M/8rhMmVG6PZ94Yh7ZWOhZRqH6HmCDbIlerEBoDb427TLZAsfQFkq01
TcszbqJ+A0A8vAtauvAmr3qwqynQZna+K3pg/vJmPb6+rQvVVpXSVi0buorzJuGMX+bpzY9RHtOH
sDnUVjS/tUe4aJe29F6QX1+3tPHcJwmnPL+do/mLdor3a2Ywgk8+rqeC0PIEKylzq2i8zu4xr65p
JMr8v7rZTfSQbAedKmIxCl3kFy9OKlTnHpHAw27p00e4ChdIxSXoKp2XZe2SgLCkxEYRbswQGYz4
CNaM9bAN5lkxlET5lE+nD2y8KVfD2+sl/PQ/eqRLMy8QF2hcg7UzgLRioXXof6m564qmG6QH+uL+
0tZXDZjzo1QliGKMtH902bxZeXLUj7DaSx7Z2mK4UPMBGpHgHZBaYMWQOPCVMNhtd5hd1Cn/cU0A
QyrvwSuV6CnNjf0eOri5NkG3hrKr9oeTekWj+4TqZFVXWEwitMmif2YmRt6m/pEl0U083q0xV/aX
STJMDRki9jIBHquh573jTf80eM6+LJCZ9Lqp25pV/zfxzjz0IpFpBWwxW+GBjhnPjvCEDRlaGmYZ
UPDM2G/zph576CO5IfcO21sNOxO4Q4XN5ffPACRE1iTonzl3IUQRlnrFn1WEUFGkHZKv2c9R79ID
bgfDFrg9FXykp1ndgol+n+1mPrUBSWljXyn7JboXh1Sah5i3tUcpVYmXWSE1DrxKmtumOe/V/GVo
+cxE/4RqbmRKN2r8nMxgy2XYgSoiTynGlHRepxoISXAD39IF7iuSXthDvwtmYAyQKjqMaRvNxVC3
GNU/Fd9aNTr8e0jNiq2+TdSiYwi/4ybk27WSiavc9T9To6doQokXfVh1mP5Op6qIxaQZHAvt0+6P
1BqQZJiQieiMCgLcVAJ4tmB0+0JQ0rXPsmkY+76wvvsgry9pt2tv8pXNtAKyAptKDqp5+Yq/is6E
huVtVvq+9O9gmv76HGK8PS/gUrzITmCKc0WsRxouWBSaRI6+0DPnFKcIFBQpbYTkn9r6tBYNob8s
1h/eaEMw+N920PDuPxnFkEa5YGChcYlOdFoNAceEOrjPGAJ+RrmwLABUJroTwVdhg3ZvGKsYz19p
47vJc5lkI5xerX9ldLhCGiofQaRh46vIZK0n/jfK8iAjn6PbGQT5zcrX9Vqcjcrn8aAwM+tWqLco
tSHHnZvXvvwObgBrcySDtuEsddOJr4x3M8wgUT3FgcXzX2QS32DygboQy/b91E6MnBNaxJA468Ye
2C+VvlyxjvLip6l8mk2mjP0Jc5tY8LEDoL1O8iBIzfpH2By3IEtRS1qtmPEEEXTFc+XZiGHNCV99
VTozSomOiF6O+ceaBh1HQkLWcFtpMDlf+NFg6i01RilCN5QvVFYvTmlGHXZ6+Z8spK+bPNJG7m9a
RAKCmrS/O0KkG7wlntG1OFreuAcGF7wUs9wb0HzxJSeq+9ObAAH/FuHsQliRIoK5pMcDKkEKLblr
hGTD4yGLNRBHqJaWy8Wug2/rcbFq1y5OVyCRerUIKCNuLPP1gVY6fXFWcMvVL48Ht+3mKxePdrWI
xscftmZ1Yj3iNpGQaxpkXwrHp600iEbqqfnUu+6SrwP4eekVBl/Y+b4VY+9jh2dAtXthwenZyyj/
2rq1C3tiMZbRCBc2/yjz1rMxgY8Qzi1yilHg9y151nbIs6avTxhy8vLPRdH2l5UknSpZo/93syK8
GCSlLgFi9Vx2hNRib+lDo3ECvKMEbaAY2vaIOWGt64YSRMoK5Hg70zRiOWaYsJMdW7KS2eOVIdsd
n1/Qt4Zuh/SQiKeAiemNCYwICGeCYGPq+Wt/b+tFRR60idR5OKGqr8Jk2J7Cz5AZWEQDOpo+XH4Z
sJmLLS8Zjz536o3kpx3yUJZHq7gYb/hjBghErnhhPIiodGmcu96+fAKZhGC/QvAFb/t9TP3hQpRG
M7+AbicR3qRXSMPHiomxwCqXtui4MZviI6KnPo8r0GI7UC/s73hB5IuzthknOlXoJwgpSjhVNYAU
IS0QlQuju3k8IOC3MBZGvAFvuHFpJ84cbm32M0Tyjbkc5UE0IWFnWY5i5WiPWEGi0JI5EAK/1FOk
HIiMI/OkY+MZtG4axT3L5Aa3+3uXikd0TbksMlvITy2E7Cbxe3EdTf/cUCFAYQ7TMLxvtoBZKnDS
LgGp27ub3siAYBW3pPiT82cgaM+PMvZ5dSBZXWZBrAM7F32qlOW/bPBOBakkZoInuTqyURgEe0Fp
E5VeS2+p7G5s2U+YDkMxffRsSewEupb5kZQYHVbsY8KnOXUhs9NSQgDvccV3YS+cf5UcRxcHk1IY
G3fYs8oXko+sGzNMUxJ2wGr6XLE8YlaZDROpZWq7qlTIzf1obS984nr8gFFMvd5VserPaFXBCZ9G
IAYIgQBqZ8eF2h2r3qRS2uQdhpmp3EteHFGeY59fn4WZnRCIwqOFV9JcLgB5rY1k5P2cE8zk69+Q
D9p22uUFyELtmAE7FrtOMKoSo4kN5iSQ1K/XU8wKhO/skJXAkyKgrUYvpaxN83UshFBu7MJkPLTf
/4bD85ZMSN6NjW9jXVNLn8FdzjMujaaPJA/Hn/Y2dicAYhRRygw1dkY5fkukGVEDzhIBIGJ/w6sT
UR+Ylm4uVdsCOk5zh+S0Fh63R3KSJxZ7EAXIhSDPL0C89HMNOUs1EsIFgBNjZZDtYSg5kbI7JfPn
xjOOPa6Xw5fM1GVndBdEv/rjH+Wp3UWk8u/4/ss9HA25oOnR3jxWTK52Rx7NQ0MXX6LVchIQ5/gz
IifY5TE+e36U0LLT58y+JLywtKaGjd30OMgSdVh1IzJai76opqxYYy9lklJI5PXeJ1PLVyH24rrT
tLW9kEoyII9nS25XCdfPr+of+gudPRQsz2bTOBRxwXJRuivY5fMz7kHPa4XdO59tGZ0Cr/AFYw5l
H7AOp+55UzRj6cKkL0d82fFOM2Sm21MV+8gbp5O+gV5ndVIrR/eNK3BCVdpMCa2E9YB9a1IcGn7P
FSct57EAR1S/nU1PUns7agSKOHZw+VxiLH5NQEugqK2PwrnOiCe7v4eAVCPyb/54HGxnncoqzqF9
DtJcrniMDl9urNnSiqSrBMcfaw219MLXkzzv5L0Shmz56hqNKpCoNXjOgXX8O7auyAjLMSt0Nfv6
OibAHoTt6l593ZcjdFzJ6PaiXKEperKe/esrABJuVcpnrxchmY4O1JOfqwYCu7I5NngZsFWSx9fn
O8/vFAUdC/hscWXnp+lcD9zm9NtriyB+6MJG879vh8qsW9i9pSgjv74TrVwSd/EhVCn6q7TrYjGT
QXtMtB/0AtmwuWiLBq4nvFDFyYc3HHbbGzOuGxzuQJkpmL5l13TIIwd/1nn4GpgCr2OpeLPeyriD
8UNQADeLI+eS8726Egr3+KXqOPleU4a4FJhcuZJqLO7ECp3cDWJX2rWCNE7tBp/oBKj4UYgE73DM
geJbKILLMWT2cUSxqieaBfpd+ixzPSskiH9DypyRoetl1GPMqIKXIrOeKLoeM05bUhD2wo/dboXb
PUp9W6QlFPf0fShaYoS97J/hOT5pk/fdFT4KN6fTcga6mfgrofmj3MEk4U9SxRV8znLXbbLKLl8L
VUzCnl4Fg+o2MkvFjNxTRxUvF23HshOBsgXuZ2PrHdINVikS4bPjhf1kOHCcQ0mgOC6upjCYrR7T
BKUwbtrRKMcTVXlgJDiLofP1YEpz9k+Z+nu83dT7UCyrbMOtykIh67RyVSSMv+7BjddCvy+hdw5E
8/x+t3hRx0QFMzzzJ6xB53SCTKoI334+w1H0BT5kfIFV3pNZx+s2WThkFrccxcuyLzgzjZMYXgAG
FcyGDWGSF7sdgWcOxmbD7mki60CSUVZQCs3VdtW1pBwQdF3irgh2OS6jbsDPTpZ8HSGQUywWZv+J
5MemGlDhyM4k93+1UlwPQre1FE7lhs2Qmc4beQtSMIjJiazpbcr1aPUjR3oWBwsaH784+BRJ/fd+
jROcv4FOMtQ9vQNLbbBB1r96w6tqXpqLLAxo+w3yP5X0ixuzVen07i/CWU8DwoXVmki1f6SitShO
AA8pARDc8NpjJ5ujv2PZX3hYoHNlhkNMKwJ2TPpWDrXek0sqCS13vZ8IzHkm60KxFmtz4aSeCLqQ
ktvW4Y/gmjQHU7rfRUM8dFzhR2gsHCSEdDd/vwSsAWIOiqurMJjfMaBUnNAV7xBTd/O//aREiHdC
MEt3z3pnbIdhihsy/FmGyIgeSA55SQJoIKY976c12oaBL/Ogp8a0LTqHP7MLVmDxbPAtZjOpBWdb
N3KAli0tn8IFWYY1GMnGJSATWoWfneDeIMAoBAgkqCVwBJMIHhn5ZYTG2ZAYizgFLZGzQyyef8Gq
PFQMKCp9aWXEvk9K8azEjvEscaZBTUyD0Iuuq3TB/glzMeJxwOIkl9dI3pSaqqEYrJ/xIpkAtlHI
dm5AzO2pZjm1ZuS/5ktiL3I/I3YYoyDIOmVMpERSOEzdC9J1MDFZHOLZtActeaIPtMOh7tIrmi34
5lwouL0rElPQCcoFWckKl+XZHvTNFaptf3z81CQ9Q0eCVXHL/p82J1n9CTMnL5SLjqD98tBLwEPB
rSh02RyMdCJf8xQoaf0KN1X9M+XgCPZ+V5/zbNpZpDMbjow8romTTe6bR9CgfEuHVS7D4K1z9SeP
gS7BTKeirBGo6Guj0+7oFqqTgSt7d+mnKdsuNBMkF9Zc9/nNx5+xjmUiTha0Ms2WeNR3bThYdlVT
D4wHG7aDLnr94vSTRXuts0e9KxTBJYXUxNBk1XHKWYCIWBu4yDO6+1z48o6D4xFW1ng5GDzjOVNp
GNxS0IqH4kX1xsYAWatQ5Q/FsfeDkNKmobSgIk7s0x1gEQQjv2vCgfxrfUZfRAsf8rHzOQHV7sU9
SaRhzFgmQuHOVMXg4DoS3I09sSAMIQPk+0BssODZ1/V323ekN2kPqOd9h8fwffXXGuhcgDby6Vt4
9V5vZlQhFhKaAOM/jwewbK/rXRO/QsDIwnqeOfRHGoU4XHLp+voGSC8At35Ceq9ZKrlk3yDo6lVr
ks5VQy4aXDlJzCYpxQCazPtL+6pFyx8NSGszPJrMu0WQZ9F1yOZxdC2XUWQ0fwp8QvU1VI38yFgl
a4s/CCsZ3OUKw6LLPU3t11qtFvM3CrzbH47AKVolieEgOIAxg794yyVUrr3Y0xtQVK+MrkUmhinK
cMmL3zgZiqJuAsI8dZly0ZG/bGFP0IHeMQqYkY1pxow6p4yWgTQyqP4GO/XR607T1bbhk2XsFAwP
VjwricWMgKCf52ZoQi+SuzoKyvcAkvrHgK7KVGKG+U4+d+K2BkNbTfz3lZmu/bqbzcZREVgZHsCM
YQI7+Dt67h6o3/YrpzHaneogkkYZqQ3CjSCxkp4bcctaQmiTFf7RgCW4pBcLAguJX58YoThEcTGm
eXmu84tT0zPkC3zSpE+OPOF8CLrBwH0lNaCW+TGdZHY6t7oiXBoe35Uy2c3HTkKy1T1E/P1nCW+S
HRS732rsTrAC9OqsSqZ16t3AiOFxOLqUTZz8JSAdSVJdwUpEoWLXQ14swGLVGCJRT9X/3nO+cGwX
3Deyw3x76Sb9dQOmG0q+ekLrA5bZ/3hv6We9kvFUdQ9jG+UJSy0W+Kg/FvPXC6HY/bDqz+ZLakPz
7cIOJcplC/lk3LZqcoQJM8uBQUXr4IEuGAecCau46gIEMSCtsc4h14ob1MCl9jvYSrvD/w/Q46Al
+ZaGT/Nb+25zsys+wDciTJj1RJJFnJ75cLYqdMa2ZYUDn2P/mB+84wq6aoW5TdDFBJ7okywBTr7W
oxjDccEIc0LSMHBGe2zQbdIZEylpP1Fdiedr9DqpTcX68gwkzw2HiLFt0zAncR4M6ThQY2tVm2k5
Z1CmpJeaxeZixnAeiujaProZbuGdztFBFIIlZbzJCryyB0tzAvbnsdMR29PCzQEbW5Q4bhj8ifRl
4Ye2HX8/1efXIwItRFrnU5uLJsAsHngikEb0azYtAIq1KZbs0YerZltzE5YrkE/WOnYKHppy1SEg
mxgMjVA7WM3SXzqUb+p7nb5LkLqO1VQ4fP72uBSoUkAEDNRYXnoMYbIjc/vDuRq5Z2vq/WnoLL9K
S/tAj0izZXlXz+LEPg1NqAfjXIpkL7jCZYkk0hrcKMO8fU1nPykwufuvvn+rqlmBx3yjA0MdXq9P
YMY6er0lC+6SqUZ+oMirQCp143ClHVzQdLdsK0X3VnvmAjiFv5+NPyPS7nY9OP32zIyEJ+jeF+Wi
VMqwLb1bc2Iy4619kNedAY3mmF0fGwQkAVLcw5X/JHmyEFRY3uoFw9aKAmW5DzQUgJGtxSUI/ztb
agd8HBFewARIy6SxVR8t9u01l/N1ZFjWXxUoqUtAGfm7KBT4Ztxz3D5L0Ck+b440CxwvjRA+Cj6x
v1Dcdyq8a+6AfHV0gSdkVVVdaXqbDvJPjCVdHRokZRGMTLALG6dD4qNm0OF7NQN3IZNjLyuGBVnL
WU6JlqkWMBCLxMqeq38JhIIN2GCKhWiptbli5P2bZwM6N2jpWocVPt4/oe8Olok126gfrc9Ysd8N
R0F3Wy5N3HjJo1mM9YTBYvGcGwiEcS+5OR1YG1G+rCFcNfFzhiy5iF8i9aD3UevEAe8ppF9VLfCR
X9HwocUS9dkMqC8CTm/CznuXRwmHOAEj2SRjhZqkIJcdoeCQmJGzee3vgjIyAvKhHNuqFmG7SwQH
LIkiGKOhoZcLc4MG3BmA4ajWafl99ZXOimZp/ouh+wMFI0JSiLbQFUQ2Vn8e6+qpM0pnLUbvJYJY
jPtBbxLQRNCdoU6Tv57K/bOQB55Qem9cQy/dZ7mkugeqCPTCZ4E7l4WvRZ3kOcu2j0Go5RAtGDg7
eqm+jWDrTOdK41lBUzzbGMrruYPdJkNo6KBcUIaUy4fY+CLXt69DiLBCzIbQfJzurAnr4r35BNsP
NCwOuOHPvqMiZOlaqpdz0SbuOiuayM21qUhzg5qT1YqxRVG83KIKAnD0A65EzuQm0ttZSgL+Ovh9
p8muc/lqL7K1mM8xogAUiqpYr+c7nHCMV/ayt5xbkP9xY72IrOSI3nxiOohX59gP/TW6Ai+1tx1h
7ubWYOXxCHssyxJslBzhql3gEDlX6ydv4gqQs5hMNBKPd9DMYCVV6l1wNypZ20hRPgrv4F3Hgh1V
Ri93NTjdUDWLgv3Q8UTERyHjoEr18yMXXgbF1LJq30OdFo7PiCsI5Bk4jrcQX8ttdIpdfJMuLfi7
sgR4WZT3qvZTzcXkWIs34tXwgxXLrsLkl3x3HkkPsl9GAao8wtfOMbhscpoS/knTcMeB9zQlwCSQ
bPIHASHclQqKUwlqYWKQbnRAMPse5As9sgy9rDVdE5bBA1jfF1nEq7yFF693D761RfssUFKOXfSj
qoDoDJjeNVOas4ifLouIYMpvrd7A7NdlyYQsNCvYOaU8xKWeNPu1lVQwx6gUY/Oo4OTnAzE153H9
IMOPO16d3fO0fdAKYxKofgysEphswRQAI6+X1HzIMHOJj/m3APNpJJyAEo1gEfRDAt5nCBs/U6vC
82lmhmHswgeEXINDbTBGvEdr5Nv26AH1pgQHrTiM2W2hbJ9GMewIrsMZDqRsQgAt7j9Ky4OP8MLr
FG6giZJVyCJwXJnpIFug+s+C9gKYhVMpKGXPOQP1s74JKy4mS+W7sCDYP0kV5m2LcEOgvOwrsJo6
iEOoJLPf6mRFkXBBnxCkTjgIN5ZmbdUZI8Ysdcsm2MACoDdgk0HVLkTJlUV7Wv+CeTI47OGRdNR/
y1C6+PIknWrpwoq2/4EzuQb3ukB0IyYBtuIxTbj4luXZ5pWVxJH6/3FJ9tELOMANCUeq7e9Yt3Rh
1I1nvxN47uJ37vuN9A+CpApNtLUhBRsfmx1zOqtesUSLxULMD16MqQackVkXEfvU5kL1pjEdMCi9
iiWnlDlxxIaZWfl6q+jZbhzBsJERqRphD1j14ZoJDOophQzVtHlLXsPgjBOaIdkBuw6cLMei28he
1p/RvdymJVnj20EuhJ1uUDdKNawFDc+82DqMW2mXhmEGAEP/dty220wBTSwA2MTwILObY02whvRH
Y6/NLAOjGxUDU/sMOXaYwIHYXh21ps54VGJLxQ/lHRaF+13J+ZPSoIg5fpGS33+zkXLNiV2093PJ
h5yGsTfGlJJuWhXttT4vhczZVI4TUrgrtrEpi7qNOBuhWLWwCEITh7oWozgl56fD+sHx6r9B6e1e
r9f685WnCJAwAIm2xbpNJWX6WVeurl50ZEFHIoRLP1md7mn6aUtNKVs40I8OAjI2LX41WITNpwRm
PYg2WGpbDxR7t1y6yKQyW9+wbZra8/OPEM0BkHFug0IZf6PjPyqygQI6iL9JIrhXrRRSS9AfgGVh
t1McocRe7foqnkLQ5CZZYMIf17v8dLEbCFPdwXTZSgXE7RFs/pxMhAeMlYgcU45bE4m+yRhJLPzW
Ojq6PO2yvPJetnm7mRd/5Yzsl2bfKFKVzv+eYAec+0fL/Pm87Km5k71f4M9zQmtQF9waZkXHuxJO
55xcx60ehrQX0FxUPatAswsY2kBORDsjNCg0rCFxKrEAwqhe5g6Qn6gI7SCxTpzim7uCesDeBKgJ
0uxub16mezatjhjPt7VvJEeC+68CRLiSvajt2q5BvRlbM8aFTU4x4vTGExbdZH+wNixZzYym7HyB
u89GegkmAGxT9SGDdfOZTM+ssB7ZXBdvwoy1sMa2tQkYa0iAsJWhiXcW+zBK5oHzgJywKbwaHOBI
obyHoO+gqeC2Gliwe0jkIQ4i7jwz1SMcRoIMT4QHResbCcrjrutQRL76Fx0/O7iJVK5J/p6xcR8q
RVGOLhXS7XKxILVZx4SERCg72Z0p099ERSUzMXXl1z6fthTEvAMTefxZ+m6ZelyFIC7cC0oNRV4R
JraLOGGRosU+3GEu/R2xIZkS0XGQBAQlQ9wKfmPSvBxzYNQAfpxrs05akC6Pbekz/JdQziBAqAaR
7BpackbmJD3C5iUn/YS04tIhga/7DI/n9Rpm8mx8ula0SBlLLCKZDQDZwGkcKjhMdhyYksX4vX7M
a6oLWQMtwljbjpCpf9E8heTjim8JcWVyuiMJhlD/tCCiYkjM3gg/kOdXFLI10XQJsakKeA4PDNbo
uT4r34NCzipAikOBvWtpt0/k+giM4+48tR8c9aTrC/snOAQxmDpNYLkH9YHNleopn2t0+PiGWKrm
3xfJ1ZJrEI2a2jCIg5aUL6DAEOk2M9fkr20yBnunGUD7l5dKd0v4V025Ilsn3PISpl179PwO0hkc
tpAc5yQdZ+COQS/TQXzAEVpiUox1KdP847yYpIqEa4Jv2bfDtAvW9t0nUuZ8z1pn5PRykXOJ7gjp
pKLNgYgu01NDrmgtzfIXwu2cs8z4k+JgfmzcuW4NiE3g2u6IMdv2UcQR9dhfcVMH8A82Jw68lTpf
ZNOcZdsPU9Vskss0S28+5VDA74GlWyIR2YntLHYs1h9tSQxBgkFQXVEHNZu0tI9PSY/u/bz8rFlj
CRiEYFyOuONcoqsVd18sMOf4lj+u/kmFuqYQKz+bYpyppnPl5Z58Gggj4wVCOUJEQj80STk8izbK
dvqPEFQNJMK4prP1RsOcrX2zRxQa08QqLkgpG1Pl+5OvUSgsFaF8MA7z/EIdCk9j7bC1LbKVm2bS
eYtndkDgF6C6/kgoqzyMcZTEzcCBhTzMPlDK1h18TgkQDB3HGvKJeL6Up2Sno6pQVHBlOn+aT78N
9XFJpMpsSLo3mnEnfnwuyI8KpQtdm0l2IQmjLzjxwMjZM3F3eE1rvmmDftuw8DTNGEBaGM0UqKuj
7oH+Y3VEWt4RRhMkG/b7WkBnKYpvFJlqBHG2/FmeQVASQ2/j7DkS88iGikURuu9YJHbIRpUr07w8
s1K0AxjuPbRbEDGoCF0ParwLAbalqiGiJdIJX6972Sr8+nRIQbS9wq7++QdT32fwDBu1QKhm/zYz
SrnqB30Zft/7kJDHyAxZJGJaIEbHAYPrCB9MTMNEuF3/iCNWLY6mFFTDOcVQ/YIQBYF6gY7zabsc
LPFp+G6c/gHgQkNWPzDDDJHLi1IWph0WhiJ6I/Env5WE1U2ASL9goglHiR1agfL2OELs8BPaG/Xf
PvWis3lgP7wz7+YEDrKHJzHAXiBZcXgtqRchixXXVyvtvzryL8rsbatPBS3gmkNcvzkacJTgaXVD
3P7s0ptpMstlnum4XaoYcElGXF/7zwiCClgpSH45XiKvWuKmZdjH6a5kQF86/emcNJIOJD/pjaDd
g0JrO5i8dyyAuAUMvQ4+JnD8co009ieAi8TpbYelmH/0NLL1OXBvimNSy3ZT/wSu9MbdcZiNXIpX
IvbeQAdxqe/MfEGD7Grswuos5vz7VYRG3BHwIVgq+K4NbKxCCcpb7UqcpJ35w7cmtvqB1Wtv3PD+
KmIma3KZOMMI4SXCXZdDWHEZz2DRrNLk5iAL2cG+1EqUNko19wSMlSDm5HBVBeDOm9x6eJatcvxw
TJUgCfsPsdi+MKoVRSwKEtQC1S0kDJ55jDsYSg3qjFFinOR6VYsbDofao1LurNKlmFMTpla/UOcR
s1bWPwJDM+9NTWU4tnyOKlh5x4VdRikTYMQfCNrVXJreK8GzxzaEhWIljd0RZYETZi1YcZwazk0Z
rvpNcFMxhYHvJaDY5GDpLSEvI55UFg1x/HC1ND3hwO+Bqa1+9lHr/2ld5EvMVyHPIaFv8ZafjB9g
34W5RmJqyWceGD8v4LDF4aoovwPTNZTd+JY2Ax7qjPkpK5nBuJmKqlsRFPWOXAVSSve19ij2wQzk
Yst47jNT2AKy4x7iV08rR+rkZdrxKd1w2CgiGg+aLxnYdqUuIgAphtBx4MVRU45hJHwiVR0I0813
GmsEFdNDBCBe1k5loDcEvqWTsWCC4TagLJ0z+lq2IBeACOj68Vbl/Nxi/mPT7Bk/tSLJ2LtmGpyW
Bcpa6s/pywVLqy13YgK2/lb0a9KTGqHml1DDaiqW86wM2Jd9Z60CxSY0POQzIShQn0OfgOv2nVP7
rgY7Y+LJrX8+10Ml3YftR/uZ9Akwemphvxl++Z6KkdXeODfHCz6fliF2YnHEOm83DOgmGJI6Zfob
rM2jhuzn4SyQ/IVa8IthLcOhwrUhKedBT40yf/kDx3HBOZUTJBXVMFa8N9wtRb2AAe/Itws0yBJ3
RCp21eeaAjkfmJUekQDHKVJi+JNCJFhGnd7a7VYWlM7gKwag1mwQQq5jBCz2JkkjmphZ+6ZvNq5Y
EYzr3y+WyCVzW+Ng6aqabCfYMr7kY+wKhDoL3h6PYmHm6r/QH80JrMLX0FFi5UJ98F0oqzs8CT3q
WIfdZu6SC8YWUIsquDUnawPETzGnqeGhFoIzvg8iMIvdu1/2WG8UG+0duW0D3FWW6bIo/8Yyt5CQ
S1n1AvrFhpBWBbrtq4SubPHNSxIUQH9W8eRh7q9RQ6zKG/L+Lru7vBgVOsKBBv8iXr1jSt+cWqhi
E/+9uQKm4KhfCVcAKGQvT89NmrKkaqBN9tQ1x2nh6ruMCMAFN85QuZVW5eyGTTMwObyro+ad0/vK
TiYzSS1YtHi8XlaKkuyTl0TmPLxgAMCkocORhFpvkOHGiKGlcIl+857WbbxXbIhxDEdDi3lGeW12
yY1yOqZgjdr7LFiVsLmEgtgIYsYgiOLtuw8+jEVC+GfBquucJuQ+qeHVs3QEtzf6+yZZ1xL3vOAZ
V5kgG42xYtRs6xgSMUybJsfBBD1fXu6G/Y+JAiUxKOkJSXQL3YgNy1k5upEbZ+f/u/q2y5uqSRF8
lZYhvRsN01t7hjvlP2rYAR66OYA1paWhTEq5WfSjjzGxWUl2BlTZwDFO91Q7B9NYpvBs0bP30V1z
jcKKrQFw3SFp+J3LLXB3QGWHuPgCySAXZOM848nc4ovOE7RofpA6Vu82jVENtdcLg9jM6tyfNylE
CYzHEQD3fdKXfGcrM87/YDbL7gnuT9W8SaUHFCPaakVsQwAbLWWvJieIfZmmBrGTS6ZED3KYEcRm
8O+G/1UhtWBB7M+8O0QNGcSgowj9pYTD0y4Wg+u9OtQhopFDrPAwnSnsBoM18KOy9UeJra5ujbqH
kQ1pp6sMho6AnWKcKZghrXE/iGMIqnw4ZK3nqRBgYp1mSmcrxJHezO/lkclCdA+Mvpj//XVoqHWC
+RpcVcr7sNTGwzFE1exxTXH0DHSRDYq86GzwaBYyYagT8qbgsWHThd+Avsd3JYgTrbGHIW0trewJ
V6Bff7DFnt3Q+KfgjB6x0r9PA6VY51McUljCgWRUmECZCnro8O2frJTQtlOBnKkuhGA3TtXAash0
QEVORbTq3h9sSZbTa8ySvXTEjz5GBToEpjrtLLsfuH1/Dtff+DpS0vWp7KHVrN+ypPkiqKmQQW2Y
GMrxqThAPHALEot5/e9KA1mNBduIs0tn40d0idyU8zwyDog5MEDZEjTnk+3liXcJwcDxnA8fGdst
u68PG29nWZakw2Cs0j1ozef0iNGd/0ke8cracaaYuSuKvGGQrkBLdo1Q74DpRz/RQ68U1zhz9K+v
qtvbDmlsJWk2us4hhYsxbFcR7Byww47B8DPWS5rcltPWSeFU3P9eLlwDbbThfdGKHA0l6ybx1rOw
GH8SrPgA2Jd32pXgG9TaMvjetCVp/mi5uk81Itias+NFddiqdwfHyS9i682+ZQXg7Hj7a57QXQc1
yrfao3p5EckYEAU1l2HtNh7DtZP0j7XPPRvVei/XVMfd3Z6qfjqO198rtA+yaJLibzC9hMhlmaHh
Odwo0rpGknDdWFUyo2KZPM0gKVjSy3S+tOTb6bXZduedqqch0XyvlDGf4ks3YTyrJjIFIiY1VUV5
UWHutaNhfQTqXGksaJ6v4QPAWp404nx7YmE6JFbqcL+z4yCNdwLpig7Ed9X3d3CMOcvLDXZDhh4c
PVz+S14/FAnTpK7Tk2xgz8bIYFIQlHVwPaI9Vnyt46tWMTqE4COtLkW8rZYT3VEXQ518chnWpjuZ
g5WL/3q8jVebWKozkYjHMR3YtrYr69kk/fX+KC0RA5PbXpMPAO4Z7g/fS2MvzT662+BaB02B6AJs
MtJURanIZMctR3/6DOerLYR/V+1Sa0HOeGlS67eF9CeGRqrfkJ+BCsmLpruBiUXp3eraCEvOwcSG
YxbVcoKaPPi363e0Az80u2PA7m186vVZ2DS3zDWS2bEpd1IaxXcvXLSflqnGoRyJVfNeg8UfqtgE
WEohpHWPPaGFFTw3pAQTFb1843XnSgwV5dJSsdCZvinqZi9YMM1FIM73p27es1iFOMxjouwk/2Ou
9GaJNH4bBqFFWuU6TduX9i/gUUg9pKubx/3cujtNdg02xMehE+d4krc9Oaihy9Js+1QNC93o1jM1
AQJRBIvzNNTNdnM8KnlJgdWYRdZDYqzj9WpvYmxbAAEAf0T0URI1c1VEKqvTVkU2V43eM+TwWFK8
+ISZzGxMIJ1zsg91GaxDqSXEkQXnk45eedsVnJFoPttYqCkN4v0vYqQj0JGgyKwGdLSkyX8wTJq4
WIHWjHp0uavqX8pCqVXYMEXoNkQLHZuty9Uw95In0Pd9ejo0PB+Ox0T8JtdnUAb4rIl31e4Ge/Ie
088B9wdmhBpOgu30kGZhswq1CUEw0G6iPBAPV2YuRPv6QxJuVawvDluG7J9AQ0+kegmh9Kqm2Cgc
KTaX9oYIohJwAuqTIxArKjPYdW7dugxZZJ39wam5M3GXBHY8QVDahZ6zjhvVrLlcSea8ToQN5wk0
+LYbnv6gzvLaplVHag94ynTxfHPZboWaJfRiHSsbHkJ5nJ68BzGz/u+CJmBySyhz6NRtCPbo3giY
FcG3GGj/F0KdC8PyQBdXjx/5a4pLkHzvuXiNajfwG6mJCizAE2Qj4OmhyAunTxfdH9jMHidIgdlY
MbdTaAzqi1q9IMFYJo+aqbhTsiZ/3gSZvXNHZKDuPNWEzghIXb6iWZzG61MuCfZPslAGnS9XSv1V
0TNq48tks/f62mvFi9xUgZKXnuYNjw6kn5quSjIvQF5tQ2TvS22A2y9CqVYjjAp7Z/6n3E300reV
mpu0ezhNOmTOf2RGUnFCv4MbngptDjARLtaBgrUl+B/ifra/7mjvt+E7mhGIcQowGun7IX+gvjJ2
+MlRc0Eg5BEbA2BqarwyCyH1+ozBaMwu2+4dVRlEL7GBuiwvn1awJPsCLL1Wb2CIgfRg+NjfUTG1
IQnVKjRBVpaR7/WAiXNZveKx09M8/vK0TnXiFkS0GbvyD/5goaHrjGt0rhCKIc8gb3uFI9U/+Dx+
bERGjOF8gEr5oQ48SimQRBSm2zPnSkh0GRIw37bWGl2PtgYEcbQB8ovAUaiU74zuQeMYVckktynJ
h/LSjF077Qe5kIrvJoRxpBVx+wcvFyCKdvXCYlAO1e933kDuJHBZLyBadK+sZya8RYm8K5NhBdjq
PaYeOeIbt3yMk+IjyCrvCrfUW7IE106asqvV7a9/me96tcZKLkZxGhFnM3L0SsWVjsl4TDsheQc+
7FGCUZvEAm9ej9CTZ0/GSCLRdwoDFRMfs2zEFigvE0cN1gMELwR/RH0dC5HhHDgaFkbx7Xk9idc/
oGbv5JbN4b8RKyg8/7H/BrVhscJRxzznVjNlXXkT/WmnlNUZeZTbX9OFQdph7s4R2iMwsvD38qsX
S/T5+fxG7IuER/MQqJ2Uo4Tc3Um28MnH3uL1RUs2IMoOWiIzaYyxE7W7rhULvfm303E/HTEQRtSW
k4qwnuxq1EEfULuxqPPvoVkHIL7wjCKXajYBWvT56yBFrIikzTdyMb1A3s+VomJuejsVPuobV0aX
DAHCW/67kAc6kWouoN33EfSmzfPhZqQoJZNPWr20b2oFPXSwDvMAz4PkhnhfdfvnW1/89kKzAPHa
4hUQeWn0mR6UEj7CY1HeJHw410rzh+oRST+m7DxqH1H9o35SXFLOoD2vWXB20nyWHV17UxshoTYV
q48yR/byh4znKcz+nd5NgdliLKUa8KhRLbrdLeRw/zpvBtOUGK0rw505LAvMKznOB+ykIcQZq+TF
XvKdv2/w1Brll8TpcOsyX7fHFovEepFvoP2Erx3pjqhxjZm689P0jmZtWrnBPLzcjrQOoRegm+RN
lsmmgFykJyRowtyjNVtq3hDRgKjxnrz57VH78W6y7LYHZwNGfacDhdMJDrlWf9WZ2qTCZnd2IZEM
ytc2jPZPmcf4bWZ5+PnY9KZPkRdWYzzzND8rFjDZ94iXe7+hOdxtZSc+tLgYUMQ1+UsXrzM/ZgVj
DVbiYQl5kJgIWiIGZXeT+gq8IuejdgVOq2iR3EAz0XktScaPUmCh4ds0417OeCuJTkqBS3F+CVXo
gHWRCACRAEKjVhBTVXuUfyTRf6pjia3AOEAFuQ8qr5S76zYjJlIdbrfwI04TY1Lw36L30XOeTjtp
NGlAXsyFTfcl+wCBdX0QeFmv7s/YCmnrRPsUtdQsYqtaZ0FnNzR4VdQUWNBf0ZoMbZhxnRc5kgeL
5x6tqjvTl0b/VoWqyrRUBvQrpyscu0noWKprLXxPHOoS25uouOJv09SF8zzjqPfv7JJEb6sKKxAa
6fJOwZZDcdPicE8Y4XymNQh1xtOUqkpSyXNS0B+Hu7GSoECK/7pRJvxv3dtGP8K7S7BvUP/9nfYw
LNKNlhLukcLhU2khTHHTn3UmJcCY/N40P1VY/489xpDSGUksh+RzAb7X6wR8lPu/uNJQTUPqWKeo
FXIr9DcnHvxFm4a+J7zEEeXmpcbzfvrND4wTVguYyOFZ1KAC2Z9MPcehdCfMje3bEiRMZG3PKl4o
0LgEar7avEBQcBb+V+sUY0MjnQclz+Fkr1MwrXkq+kMWHewQ7egpmIDud1sBgdNemIfLSVShkXyW
NSFo2/dmtSrswME5lqdNvvbff8PcIHNL4eK+InmYFxNgeaFgNd/cm1zXaJ5lvADDS1uDzIPX+7DX
vpHEaaNP2y03aOzPPKOV5m/QFcuwK6GPzuPEjCGUQi7emHsp4EXQ3ZMM6GhvGHOIUnM3u8dAwwuL
bSRfs/QxZIkeM8TEmsB0VOZyUwGOYFvX9MI/h99vQO5xZ+OVwNk8Qn6NALtQdbunX4TzN186u4kE
iCflo6hf86qDe9UaTdvxcY7IiNoBAQz4981XGOCHo4MZ7FdtIBEqdULrH5eBP6fftLDMoj+wMvwz
EM/RfTod7bU0cKWPDDXEBDKKQ6hTJ/2CpXUTHAZYvWdVRpMBklZIRnSMc4SZroTJzr0dMOurBoli
HHgC81Hc36l3MObtWkHPInmkN6fKOAAZLcmPHYJLHE11DY0Kr5BBcBIUM6UQFskw1+/iQbA2ura5
uFb7kKcNhoxBblQuEMCmN275h232gA3j1wPVds8pmqFSGpaGEGQbvrhmO8rJ11soYpJY4KvbXmNk
mLNrca6N/FvhZ/I7BPs+o5xOrXkcJzuSAIIFV1f4VaKf6MXlrIhi/6N3GgXes0kVlaju730BOCuq
TLVKro1caJ6oDom8oE80tCYB4juyvkQodaF892Fi4P0PvEw/iqwoh6HiKj8FlBLvm6MLT7sJ9x7/
k1/D2BnVqpSU4OrQvncEKnN0i8wYmHdwgpBZKNYbmlRSqMhaCLYi+cUiEkYVRARGFs8nuREYiij8
z3UEyFuLe7fDcSdBVR+G8R4vkk6hV7jOpHCRFX9CDsY+zv9KtbI4AfmS1+FDKQqReCFkekK4pjVa
ak+dNWFd67o3aIrE6yByi9YIKZdCDI/QNZW+zwbv46b5CnvV136BKZzJMg6GDNC4nJSs6G3WVbpy
MaVVh4TqNWFihpFip+vg9QS1INR7kdZeI6+T3OvUQt2gvUXOr0BShkNK/kS6NnbthChigadCQ2GT
r8r1QV3sVh3IEhtB2mJiZRkZnkYaohG0Y8vuhCI1eEXTUk9wbyQRlxbGa1oXv0Rt8LBSCVgg59Dy
rr42cKZ37J6lOlJIrBfdz+vTQC9aDHONOr0oGxt9IuNruGiUoESOskXOX3nyruhUBgyzeX6g3xMC
hV4gX/tYnQrId9/KWPFbbrFjwbH/6jykLbZtlXeCtnXrfRMF2xADMRjiLKBbjHe0BTRifgsZ87kQ
EBXJ65igOvs5Gj28mi07vCz9YevnlN2UCniQCumCtIH03z/t95of5W/Q+D7R4x+vseS3NBh3ts3y
wunZ4/vO2cDVnun3EmdzR4wvgmsCiJmw9JQB9QrEe4PPdZPw2+oLW9kaRe3DmxRNCwUa0YIbFUOZ
jZL1Licj4tMtxspry21GyLGH/jb1rNvOD2+Mjeopy+pLIremE7eNbUP8KGyVM+qdrsGhiOiZ8g/d
OJR9Xg1Q53gD4rhY5EWbDqblxHk1XRUN8pHg7v95W/w0MCNtqMkDRIh10poKdUFbqh1cwZKym6tU
NRawrWwW+IQDqUZrpDeuFJMsxiWLsHWsrsiIVxUncgRbUzIWIpAwtIp71sjfhf3TQ5crZEd4Y0DW
wqIotaUai6WfJWiSUwX4etsb6Znd4EUUo7SUoFmGOyE4YP7BTsIiose8Mr5pbF5Eh+UiZYiF3D7Y
5NbYLYbTosrPpIDH6P51QeGqYNtW/ldINj89pS+HHZuKajqAdMbjExouIBdiMHk/EWCkUTvt+PWU
xF5LX9KD2C1kM4oQQ7KcjJAT3dYz3cyj+HTyV8QeYXz9LVbuI/ZC9k0PJuWB+uiTsxdpoatVhxB1
LS/pnSoG2/KE0GUTYbw5RJn3e3Ra40QQHAzAjMMnLHhtlqndcx9Q5fkhuabYDy7SIXA5QDw+ppy7
vrSGsd+2SfP7Fca98GIGmho7gYsYfRU7AmDRB7+D11Br+9XFxU48/iZJ412GN86La9M25wn5rdVm
9SQ5rwJJ0O7DXmzTmuOyBUJiTSnrjY0Zv+KmqHDef2JK/qG0GcNRiV6RHCjvN7rLL8YWXoKI4pSx
2XYTgRlY+3HrlDHeJ+81C9DhLKzWikcYEdjkB36Fiu++ejsvOY73fu8u+mz9OIK8g+Nd/0r8KA3g
LhvFiL9SHWX9aNpOml4kmdDTeHHIG5TcZdDtBbGK4aU1tHN7g0N+3eYyMCJquUiGSCF6Po8fSLeL
lsWruA8zNqylhan/QZQq70qYYJUx2eJ2PzL5iCVLsLngpB6ZllbnaQasaxakh6PfEA6ynW/sxHs+
CsfrtNixArD4iRZLmGO239MaB46x5H8gS7IDiYTK/dxVHfI4PvrpfXmtOzWUFyIn9hw8/73JjAsw
iIAjimyK0sWSGM3bOHUFTrOU8pCQSGf70Ys/IXft7CCe3dlE5zfNOC+mU0SFicbisc4BbxHQ9SoM
ruXfVmJ7OfdGH2Sw4CXycXQz+YOjoPndn5PjyHgOnRDkJS+AHLxFND4ujYeCjuO3x2+SsyfmhQrH
mriosDaCjsQ6EErT4on2Uki2x7fvXeSvKoIfAptB18UTIK8RVXBSNXfFZ/Uet6dIx2QJLYFYQyle
kpmt6BATwFBjFXggoZSaTMCrr8EGX5F5XhORLa6EuC4UZQFRl7eArvTEGs0wx5H7pKhgYUW8cHUx
3QKem0CzDIhbvTiOR3a5dXSNwlRtccrSef+GbLQJtIxxUz+ACm/Uulp5Dlpm/Eae397j2NXTtOgj
nNiZ7Q1oyKw8+JYAQYHrN2dcNCCCVLC2Hqy61ilGADwk+icsqWFQIBS7Mk2JK0g9TPQwX2v+ZaQm
WglDBjnXqsXiuTFSBREcDsw6u2T1xIHSYlbFK5Eexe/Hg5nYEX3UlXFB5+0rysUEO8zu3iLNiv/F
Wv1pMuMGNXL1KHpoXKQrMshhIikqvV4JfQcyyPU6imE+vNEZ9xqITp03ghISEPEHs3oUvtlTbhRH
+k72jQuCGAjITD/nFk0KgNt6M9OkKvyp1uJdwNa9UvdeGB43Bq6xQK0LjtEzfMk/2WpukRirXhdx
0y7F9wCXlsfAi6xmIqR+khTI42SPiMmYQwFIq3AnmjplaZLDGPm7iFLdzGCFg3BCCgne7GZvgrhc
YZY9xu8e0l1Eb8MlJlphUOq9c0zyewXnG+g8ZZA7MBIlCGDBDD7ksTOsthhosx3aNZVhitFBwHKO
aElTI6C3waOgmq+0kQaO9/5LTpW7lKS7xhIex02SArYlAvdDfX1VBMR5wb2RMkf3kbA6zLqNLKIp
KiJb9ue/+Wv7+6+4i7dc7QeePl+V4CmNCUsDPiMc8iw/BDO/gbhkNRIrtRp6JT2Hro6qEh0pEeer
AqNKCqzsu81QEs8piAycoAXgvZoe5C+EYXvtdI5mVUfAvchG2vSvludBk1rCZeAdOUSANaZE2tvF
8UfNw5xIOd71RfAz9YCGbp55+iWBjGz34BbwKUrDObxow/+mqyRfYYcUEqJ/eFTntstN3pZsjTrx
I9sqmDj603hp2qFRCEVqNeCWZlMiU9XWkQRJYlRlWW1/le9//5HeOkdomrCIETaAVahgMtSQIk5Z
/pHWF0jZmAgjoOSrNDnp7U90ngczwdeyNoELINDCscgAPZ1mU0Lb5ES68xy4q8oC1BkqBk1Q2GsK
1U7iNitLbP0WasCnSuaLUt3yBn8WkVTGtAifs76RQLMUdQg+saM/2UWrBnUVMKVEiOIwLDkfBxlc
Wp2dXkjzDBug/G+F2+D5TRw2oHi1ZZ6ui9HlWtn5TCi/LjSsdeip2l9zjzsiM0yHcm42zMDZVOaP
tZnFa+VB6+OyWAa1QlMJkE+lhiWwxd19xN1m9A7AOfjCteL81kHw44qESFDuIOTN1lc0MRlERE8a
oq+UvLI2BNIvqEolaMGirC2hKxfPRiFPyKO6bu7BXA5VDR7877K9ErAUec2FdPb3U1r/7ckMsMLA
T+wdyz4JLz6CIPXTFxDWfaSRqvO4Znz6++1P9txKbvrO1ghkxVn+5A3k+1msTLe9Mfy/N32a8fZ+
ljyE2xr8zfvxXzATK7dvs+CCc+7X+tCvdI6/AIqYq4T9iqQ2M5OeswEdL/gv0Lczt1vC2fk2KEsf
qf6Pp/5OO/D99ElhJ/hIZ8/KONRWFOxHEqkpg5bFnmiSZV3vsRUr91NGVV8QVQgtylfQzL45YHV2
bFnA3nCdcnl/pB0MzgSD91AAi2gcHGLLaAIC3KF5nQbT8+CK967RJffuZTe6hfVdMXSibHBr0S1r
kJL/R3IbcTSoDCWSo1wzs/8dfnaAMIh1NugbBE8Cp4zG7pSPy4SmVg0W65kHxsLibV/a8/l4iz0I
qV9Ea4AKBy8r6PcTnCmxqURrkCzCd2WdKxWvyYwROaXTBG6ZuEwUxwAybBajuJSOITseQlC/tp5k
TK13bfd6eclyWW92VRed5EAL+em5Z65wm9YWeSY7M5K5SosEP2oxGOB3OoTlNhZUfdUjA5+JhFEp
GO8yDh90Y4ywoRZcaiFV9d2njYg+6NUlNCrH0TKrG54qWscD0Lxct5sqsbuhtd7yF9kgDU1XSmEH
rAjd5nOS0A4x26nqsYg2dKOyQvLWa3Yi35BHUsKwjlzSWyrL1Gh9g+VZDs7j4azyQtB78ndTNtQY
n7yF+G0FObLsLbWzD8JgAbpcaO2prFI5MT8NsW1DmHESAUGAkzT/mqvnwYWeIgd9Y+rE6S+Pd62Q
7TRmpufqCWgpnkCv4OCAVwwoI1vcDzoVkpQH1IYqp11Uy6KNeTcGRChEM7hAK0pcHYIlF0vrKkgC
VdraEZBwsSzlQ+WuDLQwOwQWhOZNUs8fDQk4B2+/MOCsp4ZurImJaQOQ+fDAaTuXGQmWHn9aGEKv
eWzVWPXOursTn8GjkUAtrygH23HP7ecwRpJ7XPPiTPOEjVX7xn2YDIVie0avod/kcxVbKH60h4Uz
cboUHB0735Ktub7lIn6GFr8D2QjGqutNqivYZA6H3IDmgkzx297qrG3mwSJ8gIK0WYBq4vX30NOx
vNCzTqCZjdiaHxSEIe4wgoT9tFluN0nQFndZ73dHUpU1V/zQrbGR8wcNoGeW3/tu/U7Q5/KmjVCr
8Wge4jBbuL7Jj7I61M+btcMn/IjZp51t2KJgH3BB62mE+icM30BYlavjcyFnBMf48cj5FPpb3wHI
r1X8Z+uv6Yhnte8pfpMXW4orHKJClrQO1wR1LRs6eSqZjjO3vLPd1dHY8/iKMrQQ+uS4sXbsiFCm
g9RCO/tKAECjKOODarIlzQqRyXbNzxRaq5rFhZJkA03ixyvyutcgzQLWPWJXKihkUE8YWNwcYGQY
/MDUkcqjzPZfOM4smyS00ormG42PIRyk4WO+vitI4y25D9cudk/jseOB1Ys6qeNM0Y5mZbFAjzlZ
+NCh9rvuSswkOprGXtp1auo00h1EXTT3C6cX6+ZwzVcMFzQ1HrbYUlsKMtz6S4E60iBp7wVptMhj
JNmBFoz201k30BuuHl0upwJgEe5kFbH01UfgplecyLEcZUT/x3TvbHfJCk17cq/18cbH2Fxcebm7
coj4g2EUzVLQV8A7Ehmwhhp55kz0b6xmazaYlOy8aiDdClnCN6/E0KvMDQHST7fTuhONyFxpqaWH
Xi8LRS6G61GgycbeKuRhzSjnW8KLY+0qL0uTkco+donNNC8n5dBOxQ1/+dONtZTZFbxc3P7OI0jR
4/QGmEq/xvTNx1NZy+S198cHEtv2H0GCTeANqZrAsdvkF20Ve2BUJYyg3HTkdL8thN/Dq3zaEtrq
Vub7n+bJbKoBHMGIe7CiNt2JRbur+kIPjhlP5Pcjzmi4awHvWce4Q287MPj+ch5PWiYa0AQTmOfD
cZBT17pfdL39EBzt1rgRw6oS1E89TyyjfOeflJWPaHQUogFCOi/s15I7tdCyts5RQg69ityXUAD/
VVSDny4t9H1FbakFR97Ons+VlgERuOmCqEjywdl/hxQhjoQtYbTApEnItHAYHZct5GgE3K2t7Bsq
KBkMF0pl945K0LmTGixtoeRU3GMHso67F1AZBHTwHKCm637cf01/IEL6oP4iDY3HrKZIycY9mk8e
eE+6cR4TBmV5prHlKkq8k59VQ1XwTNehG5VV1r9G7VoCo0YQkG6kOaw0zQ8IvEr+hyewdXrvv0qM
w6+oVEoXuWLAw/eily3y7geEWMKwsMgqLnuPT7ZGy7Q3TD0mBCfhotGN/TuB4g/xyAm/3Sunr3jf
JDN919CaBuLt37MPXJuKUZ1iM5hRdiEy/Lh0Ch1rqwMwinhSjqpvC8w1RY1sZaWEk6ADtD4yu3Cv
6Eq1ja9m5cArK3W1ppPFU/VFEDBgkyPC6fnuN98UJYGWvRKq3zpZXY1lqJmnZ4oFyH0zMIGqr00k
HEewXq2YedpgbW/DrGkcrrWFs/1FV/bFlaPUUfib01aPI6nvHs7QL+FAzgd/mccYoui2gAfH/mqG
b5h/dp1zjBS0rSasSlyH+Fg81/U+MC4wMWH9hSOgxDOGtD3drQr33BxsKeZYVsr18CCOhYJzPyYL
0GbmLzsmkGU7mYh19diaOobZdO2q0vcVnhTmT+HOAsupDnZhyQBOEcf+BgA8H852Z5tvlmzIQvKl
DquUSf6OuExp3UDGK/pLKxF3qNPxfBg+6vg9Q8CjLVE37qoFxkaNvW1hCqYFyLbz2U66RqB29aLL
DQPah3SEMWFPrvyRTPUsypEJOcqc3VCYA9pMG8Tg2uFrRCJ3pwqPAy3kbHwUfbvCZlhbiyG28JsI
i8MVAsoNuRc5zyW1vdXrkwStHSs7QCTCU3XezBXrlot2TRIdItl5x0TaZ9YobpJmTSAj3Hk5bj56
VJtk4ilgpdBkGF3LbZ4UDBWGInBQ58bN4tSprcJA0UATem74VwDxKASrjDRYeS4xIASTbL9a1oNQ
8jHUm0LqwruYV6fQA8PnzWX6PPx7U2h5oQEzFS/BP64BTl9gjUwdwQgWOJ7lkYJn/1VkoleAlaw4
u9xdbS05FriaBKTIIl6CjwnpOr2h+2oATSecLbQTYY4tje8RBKwOL+Sj5nx5azICP35cgUyEXmgi
Nconfimi4QJINhm8d1Rd+ZLrskryWl6FWKM8k6LdU/oyNa0QGVSZ3yUxFkVtKG+b2L1XT8D7Y4qq
ZmofRJnYhDoBf5mN5IEAApJqL8Un1PLBYX4X88zSbCO9QhY4FgZ19hNOHkB+NXAn6b1RZde37c5H
iGAEJ/241rI104q0rGXf8BGCUgITChpQO9kxx6qVvNApscdByW6QtqcoHf7ETNCVuW6gR1eg3wC4
TxFntDt++BlD1hrAEC6olPHWBEXC/lk8jHsyRK39xmRceEiEbj0sVjxWyRWjWVx2/YrdwH8FEPQK
mkhLfWruKTAuZsANVeI3UIikL3gGkp2GrAEUoUz7QrsKzXF9J6sipsusgLzoroCWx3w07QuOt5P1
3ei4TYCRMEsXQBty1LD4V7EKvBUJv/qmccn7LHK8crl1SQ9iRwRT4AGgkJqOMHyNjcoTC2xE2O1S
aeca7r6jP75nHLO61HVKBdxDtUsWg4BSW3pXxsLCZ0z2wJpt3C3bNPsPTEd/vbJji9SnruiC7mjE
G3T0FKO3Toe6t/52Vr4JtMpGFa3CoNHDG15HXP/ObNVADBRmN63+n3UyojieF/s3VwSobaYTvTrt
cJMOyx7L61h0cbAanKXH1xRrajPX6PYHerf5/QrJTA3iRHAoZMoHZp2MQd3VaITVvPGGNWkGuvXo
kjHoSJ/x01pIXSAfke/J0qdDQoMVCLr7b0ipxUcIxjWc1s7quDw2zeQWvOdiL4hzbOm+Hat6BspQ
D+ebZf9ihKJRiR1smRK/rimmVqnO3JfWnJ1CS/U8V/Dx2CtOgj0ODudN8wHWM0HCg+Y/lNsUlH1u
KO/reJTGSFmMcEjAth/BqQyDw9m2mh4EfilDeG/nWiYf6i3oTmAXLIQZgZLu9JhYSTI/wL1qofbL
DTRyCOtPpa49QaEHU3aTVhX82xU4WFZWo61wrgUKHfow1fV4ODqh5AWVtiHlWcX6Fu3msjaOM8Lt
uJe7NUkvGXg4T/beV4Hpmcs5Uoj7bKLUDUZK5XHtQvOcuMmslbSokppJg1PCd2w29JJhw/LokAbb
W8b1992tU5ue74wyfvCeX6u3FHbPxQyb0cFASp0de9E7gKFwpJ1ZryUTsylrJwrYHSg7pFSKNtFW
VpY1OYVOOeBgxpNphQEmsgSeHv04Ed5ruUqhIWdd0vHDYxhg7M+L4q/0pLRngPWUrqqrVJDvf5kZ
/4uV6HSXuVLMBpIZI0568hr9fTPvbAR8c1Eue4FdoGzmpbMOo/WSvEo00lrCoP0Qmjy38xKSAhN2
DFGGGJzCvaHmlKenrUNYylxiKpiyMdwcjJXm+aQf9km81J2anF/E0qxM9cLz9TK3YS4GXbUtZjaL
y+BfJ/3BozDx6qFSTOaRLbW4/UJTSpmzIBySF9qriuyiDPAIALHux2Z/yHJOAwWhXGMvfU3ynPIS
UY9GVBbwg1fX3QSwjNOZ6dBNyTt5DhPrCPGFKMFBq8ROI596nzZg9M2FxZHhNEJ/k2K8XIP14Oon
OSEZ3d3YfmVoeXmmVfUyv9qAC+w14ribvjfJrpL3SevZnjYd70lT2+GzXtobx2SMTdgb+klYdMpN
cv8tEWSE4iOBVdAW5Y1exYG6+ZtJbHa4bV1MBq9CWDIbPNNdN0hTv/W9iOpx4y208r2p91j3ALt2
LOBHz76X55SFZ+g9VfzbB46j/l/mOAcCyjOsbGkOG194JuVHcYKjYA5KKLW60ArrBkiLDGbb3Tly
rrF0HOZDR4DKdHdU1vUbGDCc26i7c94FnxItuEBrtp2ZDelkNdrvCpcnuCKtUPZwZOUiKker57AE
j6z1RC7vGKDzI0t4apzXPmTV+SYmEEb3FeX+yWcJZQ08PCWInzLn7/GFV9Y9XqaaogOXlO2i7T5W
Ovqdpx3qwXbRsDDyTUczuSdgCMXZyf4mpa9NFTDJlNa3pfbNnArudMjJsqtyS0U6zBs2ic2xfF8f
mTkE03Ko36Ns8HmLeLNIfvB8/Vta0eW3TT1cYpU/llFBvh5nJSuxtS47vTUs/y2DZnPguc5rOxT5
my8l9cxCa76elmbY8xiUmFxA4vyWI0vd++gyWyQ/cIODJVXKFcLvyaaftsR6CXqa865lIEBdvpl5
31FPWem/6CNg7wRFxmTiW94gDVeY/HmlZmdTMKYk3IKt5QXb+3iIzV8ud9vTr5qxAhBpOtfcEqSx
2iWnEs92chzpg0+j969i4NWkkrMBB6C/lRKI6BAzEgvFJL13jXaxt61hs6mKCKMNXbreGvmH//k6
63lju2WFRkWR2jmsD2aEUsTvNMB1pihwFdH2YMmeHgt1bLtd5kOmm0Op8bJoa5dsVSkzxLEZCHCL
ZwosJXP4p9286vWd2ZWconKxWkPqkIKgTJc4YNKK+fnCk6kMp0A2ofmyc4HSG+eLMLWnv6f3TlGt
V1/U5dCoU3upSL+eW81H8y8oYylPbRr2BHbEniiEYnLttet3oYjcbEKC6eCaoZ1qffIZlAi9AVT0
5I2Fff0vPH1IHPWfDhWw6jdowGoZvwVjcBQLMi1E3lnp3nbMn2/4Cf2Vu30opY2vrETM4xcNCMrE
GYcmK32zmzPL9bYE74SLJF5eVbdr9cheOdcnhA4WvS8fbwI8T4d1pCVH0RYABeuTDjiH/mVYlYS1
Htl/TvUPw4ZwqIQbPEBX+cjP/GbAKurdxjYpWWQntdnnXsT4YWEGaCIdsc6E3I+8hHVUpKDrA2b7
MyWL69itNly+QwQcf3NFpFrtYm1gUBuHv9HIXI7cA9jYU8Sirrx3Zb7NV1BFkdIUrfbRBxLFZfYe
hJpVFmYVsfq7YOPp+AJFF1E7NI3QAsGjYQZg90XU717FYSZsXjihVGqL3xNIoXFb2TYwLwXszlx5
e0pRjT/KBb1NtN/Pq+9r1yqZ96hj3mJ9bO2Sb3SJjvbEFmdG7t5i/ZtMNH6SbqFA5PPgNV4IutGy
ZT0E2G7dNNzSuh0UqXP0zwFuSwIIz3bdCTpE0nBZCNSXvNgIflABT0x8c7oPN1SanuyUd+HJBrpT
AVoAWQh0tqYg/kRoOQu7NQK+qBr2wzN6Sz167F3c+L18l9qkeVCmWIdYeyef7P+CAX2y3XzgDH9e
4e8vMEc2CdO5Ri7cKBNrdt9TQVXDhfgfcZYrnAP6nzfnzJHoCj6MfQuZwjPriXjOusS+7ErajDI9
S918e8zvHR/hc0sRkXEUv66WKsshQe31qcnhUjMcmYzMVNQsTPSLUuQW6YAAVn/kza4AdN1WZ4Ve
8OKG7D2EYuMbZrkxq1o0eLy1X1LzpToAIdEcGEaNDLAcx/AUW+GP1ni1kS2lVe60+ZNOTXqBwrd4
vmfk69uNXXxf8SljfcoL9mk2d4qGywS1bsLA/u6fO30yf5PAGRdkK+NvBqdxOp0lWQxnBQS/Sxi2
XVpFInzLhLpAnFQO3qbjNR7bNvGTBcgRSk6RpLAGI5rXJtkYeFr+9n+md9aYjPejw/fA4P98mK/a
PfMLq00INlUppU6U0iFsRWpkrlt1LVDvWv87DZZ6sBqjwcXT2uImTwGc6U4muV7A/DS/4bGcMZFd
NbqRWXWDIUaeqhNJ3igwa5jU1jrvn80lPzOhgdcKKVLI39GluVTw/TCxLky299sTvfAIyowFdHoK
dqxMSOri0aCXl3vdo0GS2CcJp4lg6qBMazIYe17PD537l0UC5dLdmk6qG3a6j4GgR90fpMffs+8u
1tUeBbdDHnbX3NDPq3ygI/MrMwlA5X1YF7U1E4CB1J8X22eoK9kiFxbmvFq0SBdUVHAnvuachvpt
13RdTJAftCdSxiYi0qnjhuseOwegEI+W891qAos460l5fB8dI3E4cGMo5c8oZgLfrATH5KJwtXxf
lmBPHvzXWsqMvt9Jkc2zYK3jnfR9msrtpLu5EcDxAIdMht47Q21TFe34NqCoTuMaxNsvlqm73ugH
ieb2KVGgQkHMd2tD2w46nXgbx0N4Ds8qg09A7iUt9m45EyBh6EbrNwsLGP2DK+yxa5kWM4M96kTF
PTDerYQvli7VkPEo6S6y/BTjVeXE9ppiMuRBY4AcYjHBw63VX8LoGwO3/LJbCHnZATGtnqooFQUT
woaW+mfjPnB7v8nmQg/2iNF+4s+a5ShseTH1cb3f6CA2djZpPkm3Mz2eElyhi9b1Z5CC24uy03Hz
jgwy3FfLM5oQE3dk9zf3eaM0AYqDmk9zc/7ms9Cb7hU//hpfQnx3opqfe4eKH7IVh67ciyp8MBJF
rfP3f9pTTknLcYJpCAsLPW+XFgC0bDEFVc9vVCr+jRfAEgj2TPlpBX8VjHCYRJbFWrqoDqPfsOXS
cGi2qH1b0F6FWd/mk3sSErF2+8p++LFCZ42z1uDsvyj/1RL4XbqaEZ5JMEbqs+kHslDgEDjy2pB1
qcU/Ys8Z/z71FohJxeE4VgSsMfy3A9z3eZ5zxsNANTOjEGCJ0qpZ0zGjUJ0AZRMPbYMd1J6IPxjW
KVOfNUVcPDdCMvPfa9od+9Hr965eQiormfReQjAz1q8FWzRos1WSqajnxBwgQSGfXx0byW7OnaSK
Uz7tIiAbAdfuXcYBWCMxpcoFqI2vRV8Sdj8Dt0Eyi7EeeojZZLEGkPd8inEJzCXjECwSsz7didwo
ClcY7aMFrX/hrbJdU1Ukn08DqQerY7N62MXAybID/1tZpUB8gy7AnEIf68aZc7NIaL1vV4nP9eb+
IgBxondpcd7FjypO1VoNrJMzrC6WocYSokIUNqY9hbOjWzRciJ7Hnq32tKf90GoNt95ty3+kZnY8
QH1P+yBerjkF41yWtp1WqailOdIxH+etKIQQt7omNZLcbq8rXRnwrtL2i/dxK0J8zVkr3flFCkac
ZmahHQecCLPBCLFCCUvS4sbdkJUDiDxLo2W61JwVii5Lp3vNN3JB52FBRc8hQF6+Dh7AEsvYafj7
a5xGqHrlPdOcrZA0TOI71PML8vTDtRgfWx4jKGtMfSZOGM/8zqXKePSTm4yYiOECPaL/gSE5+p73
KoX9gwvJQ5wnNs/fuKKFxMda+AR5dvRXunghxKKpdQiOU6TTDaEwXAVKvUKaGsH8OtVO8f2gj3ij
7PvXVVXKMyOrCTDJN3q5Eil1Okatw1cDC55oJwwVNLJA8wtR2wMcvNOTj/mUSBTRLbrIfGF25wTu
5CmLX//teamxzRoZ4fH040vBJywfOKgyDBsb47CpC3CjzxxsN1IuxV3+Y1LtctC0II+Qe1fFDTvM
TqfEB9J8xE8jNk2go7Zb8s0SVRD951vIbIAB+zoF2keaIPttzovQbtxM9X3/LPhjJUgBAOJxS4YD
VqRMRGunLeZEoelXC0gOKL/KYbO7gAWHffNlap+PQmIZb9kTDxhe3nglVIQgj5CZMH8ubKRdpCBJ
Qh9v8iLOqUlFr4SUUSLlYtj8kiwqAoDfYL9VyNb1/1SQK9MMy9KHSK+BU/Grhx4HC6y61e3QQ+wv
o6T+3NVHK5+TcTKEVYmW5KMRsGHlvSEvImVhJLYBlfJSDNo1NhFsmGKzolY1cXil8+TtvMmg4LTb
ZAfBh/lSCcilxUcr4K2ssZdW/f4Bs5RJs5JFDM88PZErVHxeLYB+XiQY+xyONKH3RAZPYeU2gips
MoPdq29UEDhan7rVm7x8hj/0I3qiueb2w8KB1y6Rb6Vk6eljo6S7d/pNSZtiQnDXzzO7EFHXGzEz
oW9ULi2tPdjpK8JGnIL7ZAGwSwKGT/zxXPLhXI0+NkIfRdWnSoPfwRsbG9rh2mT5rVC2UBxkVKFX
xhUn4QP543rUeRxGT5OFKYLYzQ9RGMR2iXUsIWzTI3D5f7ABQWcmonJMIWtWOnHRhZp869qAFFG2
fnNlUKUtLMF62+xIh4RMLEwEP980JnWDuy0+wn922spMli1QiU1vLcDwThjVViqajrXSsyFwNNdN
kZ1VuFxpZTDG21iZFfIboG/7TlS8iURAOogMkbdcpg/k0sfDNMLwjs3DII/+2CyqjmW9nuBkBjns
TsYWlsRzMtUELqxDY7CeSgc+KsB801OkM78HaocS9Ud7BhGrfOqD6t39g65xeCCcmydz9X9rWWLY
39klGJ4+zmf2vjSpnvznl13DBeJkmtft7oIlMBjF0NbfAyXylBmNL5SUbL3VDqbb3CDabebR7gBU
audy7XLVCL+svqN8pwpZzfs2MAsiGGlLvgYs6ghKetjYevYbyfJGoS5SbZ4VTtBDxtqftGCR5YrB
vkpGH5Dzhj4vkNfC2/r/aKm/TQvFvxTUhgBjyq6GJOlnkfRZRjhOXMsTyFQBjLQrIYgEn5hspPc+
6S/d8VLwn3vfM2p9bEuTphjnYna3SLBAfwwuU5t3NGLvehCgC4vfKA065hPwCMur9gb08HjRglQm
QP5gWS3TEcHcWhlldSWrVfEYuJm4WnJEBin3uyzQjq7FiKFGvUY+u0+THdfcoApXPPcX/AP13u44
xHjJhmUsQObbIEGpdvwxCDkr8vkQBELdNUuyyJOBxHe4teE/WeaYW23G6uYIL5McjUzcok93tRwU
pEKAJ6TGMSWnB/n7sO7jSwhttJ9Gew1+f+ZKQKbrU2bqTo5darmSRqzZaJkrLnVqNjd/kVXwCUCB
qn4z/mkakH+H1mDV8tROC5TKf7FLb+z41Wn9Ao5pex6VAZpxqJ9/G8l0Zs1KpJMtGMLCwCNgmqTl
PJqmRRIvdBK3G8N2iKiW3Uq8IE6FoVXw/0Pwv5s0IUKmoQuXsbaMp59qjZ6UVdZm+jdC36vebtVx
oF4kOHx/k6JLRovU7Oud33ECkogBNK942wIhfJT6pP3Ixy08Su9pwrOUrlYhS8eIu1Y9ttv5U5wy
KjOooGArAIvGr3yG4qIi1kLnbe5jJvPYWXHGfZsqZwbiICo9bJzAsJtrVfjXURK1JMzTwJfVCSsb
svRFw0KMDcYoF1kN7SnSFhnpXuCp9Asz0UATB0kebrqE5xYQBQxsPcpbIPKen2RtM7DlMn+/hgtO
2FkkKN8K1YbagbVlt4X8mbRzPxmGAARwXdlzymXm+yetVvx/uy9qayfI48pwAlbDFkGs6usRAPwZ
uw+Rcgbr6Q+3HXea2pGbzt/JIhS5Q9+ZmJys2Okgto/TVRlNLdr0J49e79mQLfyDGfVwrdI06Tnb
+Xs7g2S+JcUsblDby4UKzfWRUbhGNIjeT9MJGqlSvJCiiC7kGHS/emet4cQ2nQib/F962EAgPIU+
I0/MmTW/oWAOS5D5R87xU9NusXtmuP/3x3IhcgeeBMdBp4agA7KHu6GmAoydpg7oOjzYMeaK4f1j
xYosnEt2PifqopUnex5WPlmOh2ut3Po8EKRkOU0vXNM5/BbboU5SZBLnBys8TowA/So5v6gJr4v4
qQgwJ77IZzWL3v2xqQ9Ft0xAmTnX4YzDgqR8WHewuDGirGovJ3Xo4jn75/8wMxI+Mw/izutzplXx
cQXXwhkBEUi//98ug8YOwf4YT63MuEqNO89QzIwHqjD93O7wqVFHIHbuCrEv9Y5LDY9yoPUsfVZG
cD8Uv8fBf4CO2l8cnJbcnU83aoB3UWx8ucqvWgC1sp9+rwJfjtxfzQwn7FCI+haiMYqDYv1ncbce
veyXirBbxOBqKR3sjkCxVBA5vEUljpjaYs2dIBt3BpxKpuT+fg7c26EbJwGl46mSQyLWKNckW12r
G31zMAnxGYU30RXI20Cttln4M9PV6pVKzZRZSq5YCaugQvUA4wsRzJi0/XiMKHmjTDi9TAMKN6og
hB7ljiR4Lf86+Lg+5mS7Ss7ne9nvybm+ICkvAdlZeC9/t2hh2c/U7IqZqM/JVgJm8J5VOhXIFTqQ
pFPZeFgPkHlUfpHiLMqbYMZPZlP1FsG1i0O7T2FKWlGqdJCy7K7wUeQPddgEpu1O/XhKf+74yXrW
w4Hq2fyuWg2KYUeYp31HvkSXtzM9H9o/1g3dutQMSr3HrcgIlLWbvFoU06ZKYLs5XEyFI9ZEOWur
LRjyde6D6jPXyVcUSmzKDz9gS8w67A1L416qvFUfQlcVY894eRkuo+dByZlbR/Skh/egP6k/ezrC
tyITMNinY37dVjGFq8FbarMz80Ep+sTyTsnxrFi+ZmKKgthx9jhnjTf5BwlB1/vABAPL+0OxTLcw
ZMPze4t7B77cPHFVt4XpURl15hiThVPqtoG0/wr0tyvysqOxHiSDg8FX/AhWeqtgEtN0SI736edX
3LApeG6w1Ne5tKMJj939LHAUAnFhD54gSSK0BCtmdXVUjMJWcEO0A7NNG+11vXACPz890TOMTdZp
A1WobSQ1Eljx9q0z6wMScOMmsqy302IXDUoZBHg9nVxaoJwP8mWkJHBYImXoFrABopiSSPjJuSQs
YbV6Xwr5k2n9TmNszfsS3S2InaBuVa7NhvIKUydBedcL8ynKdP32ZktQ/lTU4NhWewg5KkvxHcdf
XKQlAsRrx1GjimQcFYEDoTX+i+S7GTNJD2LDg29lSrP7dn1VvLVy5eA/1gwk3s9McE1kanxX9cvn
iyrb3OBSnJqt658rnKWg1x1PakACJfrzbLScJhLVVLvNWm2DNEBA2fzRl2vOEvkYoFpId6fdALuI
lVzY8l/vU/nc1KJGFfpNeIu3kyFDbXQLAZ0tTsaoveQk9q0Sd3bBICKu7d4SwNM53Bxor5i/URWW
6hTLu+G+yV0Y6u4zzTUaCsO/9bLqpQW5/mSAl4nsBnHAVs+p0EH2FF2s2Q0qjn6cvmlCd6mBkaNh
hVWRYTOiUt9N1JRcNybljwQ+qpYZnOnAKroJru5Wq7uetqEd4b8+xZv09KsUQsQNKw48cMDn8aL1
UWSfhOKNB+v562eWBPS0b9oPAC3GJnS+1ge/4Wgptw+tHHJs/uFfrYsHXeRm69f7P6CkbFKgRJPR
C2gWxLIQmt0zPJ2NH/RxPrQpcScb7UqITcPxjgtBnXzwj3NrViikInfcLhFappUMNz5/Lh+AHuAV
QmxN/UUyqIh0l6cX/Z7JsRifkCOpt2N7bmoW/QzTK+26R+8In1yH32SUr/POV6XoFuiafRg+pb/e
M/DOF2xWL+YWdY3HYewG/LXMj3K62d2HcTSo36tFFDTA73yHjKn3sh43iGxt2okIgDUUndxT45zy
As5/Omce3LCTe+SdFTsUhQMnEtHRqW2WdKgjxuXfKPA8h4ZbKi7q33bpwKiRa0tN9e/yjMxr+NAz
xIEdX8qFaT0Syuc8mcmFz6YFggdy49gWemxsIP2E+8i0jEX39pfeaMgxoeB/3sMIgZl6Qs5UwfIr
aaF3qBVj3wGnktg2RT0g14yOX3WzuBpOE7gR1Ckps6QAeOQK/cADpl9AQ8B0M2ikN2SMGnFOfoub
6mnUIltOCXt+8dN12XSSLXLyucCdpE/CbfGxNNuP+y/klUwVAnePI+w77VGqJl16R/GC/RRQBcNj
ylYC8dC5PH8f7Eyuw0HtjR5piqUYR4MMNyTflNrsy0NANYVUmjwQbpJ12trSxjLOWrZyf/AOVI8Z
uPuJlzOrD57Qkg+Vj2kHtZKK0DwjAw9YJ0IdqY7Dlk4NHtt8czGQzImNnivaldX9gxdgkJGN/RHH
Iowox1exdepscwwQaMFwdcR8DZ4qsufrKk45lZURwJ7XoediIUxF/AOHn8XZ9v/6IhyqouQ2Uj4b
OdeQlTbB2PlauTcP5LI740WdA7B11KLIp4wC7DfNcTNtBvzH/vid1OIwFyyYUTCUoMCLxDch8qZ9
4UXMbu92DYvJtNZrHj+f1dgwL0Z1xsiIP5jUFEJ89Bx35P8l2PWqNvfCiw53q1sW0RAtf9WKXuP8
YuaQUbPjkYErq+KP7hwvYZ+aqWLd6biVloWFugcrK2JN8QXL3iinoIlg/qHXq2yNj7RWJMdfXlxL
bskkMNni/P/h6RliJRLYCjRNAfOQBv52KiQAnTVm0jZrT8XTU25W4DW9U6xmutk6FZA9kDgj2Nyz
MiYkA7Qjz1J8hMg5is52iISxPNg4xa/65fP/TBRGO34QlGAx72hAMSl+/N+0YwYTmrimgmGf0Pvd
uxdB3vPZ4UvxagPttYRRALXlLdaCI5j9hvaWjvJ0MPxy3t5WsECi0WBMF5maF2jKSeClprZPqSA4
9DhPdxYhkgpRiqrCNvNXGB6GB4SqaKrzUTYN33HhKUm70aqgaB0HjjfyuljLnP1xIvgYyRAaLPIU
QMKON19afvd6BkDFNPOWrBlL+vTv/PQNIzSzTOeh5yp8Rm1QTxtWv4TOCyJCWK/yD7bISl0NRwBa
bRfTEWbHP5OzrGh0yRliN3hpRF4kmL7CPn5gIpXpiM3vhx0mpBURiFbsuqtSPrZCNM0Z1FgJJhyv
3k8OG8B4qXxTWMpKdIJYVRHoIxkeVDUvJ3AM4iQKhi9ZGnE2yPHCArXa8rNdlTECUwAx2mo9EWnA
CsI23Rpl/JYbjJkvL/vRsTONKynxi/yyRnMkCCtV8vCJxX88ts5T9/kvUYfWpl5Rd6hfVJioD7xS
vYpzJVZp1rw37dHKXA/DVwEzM3cYbTTFRHAzUIocl1rEsjDH48N0g9mOjAjCIrSfqjavkd0rWSyK
MKlD5jZA7GdQQwN5p6WK6QmsnBFIfyxg2WrxL84exHN1U5o5qpecWZ6ixVgLnAKyP5OQK0ArFlpI
QXHmA3u/bgT8p8wCF6bo9yXwGg0XkCy4Kecq3mb+F/NNZI8CiLkmLNyrfVjt13t7K7kmh7QS5Ysa
XR/whY5Bh3n/7u+WvgvpdrKeTMS88mRWs/PAl10GDh4/8exwtxoTn0V0mSILSUNNwskkI5eKt8lI
nnTJeSYQ8N7rQOG2EEYEVWHRlGLBi87GBROE0dryJxGKXt5byNCN25rL+4YO7sNFu/D5wOysWhan
qTX0r1rlHfODBxgxVqHpR8u/osFcoaVgbs+/0z6JzHrylvo3v6QJwqOnGuTqisZPCz2yYwAWn4gj
Cy2GSt1szAekRAYWHDdeBIZYMvN5dxEWlOpT8TJ/D9ygZoCYNn/dXMZrwLy4u/CBLOctBzzrJFGy
3w506FC5z6sHGQU2g7jdNHA3zlUleiUFUQb2R9Nwt6SUkubDYaWHtxvBI0Wwp90rMh0QH7eS2EKo
AxWgWZUrkuAFAgPtdWji3whLxe1N22uoc0WuTZXUJhkODtxihvv9CZgMo71irfiW/kIoMS309oeD
JBAoh9BrcytYr8/QxRld6jTFWgKXVA9NX70vgXWpQHorrHaXM987iFH5O3AE0eekI2DEemiVKO/C
f2K9ZVvTNyFlAjYmupWZf9xI8k3g98IJG3MkJRUL2ILqL9uteXPUoaqGY3FkArVFdEbeCwqKaUqD
GNbjwUk7RvjywPIGyk/6V+jlFiqE1XEiuCHvvYyHwbMiw216NnlcB/c5RapF3r2pCk8N8HOgaYw1
7RpkprUPpU6ac48IzX1R+IwdrsMTdmBP9SfTLd0oWGeHb3bNbfV+KEofIhv9qyESVYxHnUM4lo1+
MvTXuff/hh2Zr2nahDFKcnt+p+6gstfiGVPy0yztZxzSD6ypAy8MLGXULvvJkm09SE8x74HPcdLM
dPzmwLKzFZzpFsYKur2Br/pLpQg4yRUbonD01IShEAnso46CYTUuaCYlX+MxRHdC6r/fkk9r81r6
AzD9L7KPfMV0BtlyP3SnEYlJvRrvNW1e9Ga0ZYd27f9WVn6m5Kj5xVrk1mxOIECCO+tVOe/1wsJZ
Uz9UNW2s4KjMwZZxtFxtZJDzHum0VvKj6734OYm1mWAWsmpcC+1GQ5aJ/LUSbhF0uQ/uAdsz46OL
H8FTN8ZviTCu+xTffv0WhwZiR4K1xU33EFJsHZ0kC9aMw0h5YxX38wXZQ7AgEjShGte3X/yvjWlT
8tNL7YQZiK0IPS4GbAr1LGjKcba4b601XjthwqOX9vAAe0FSVF3qobpHKJz4r7NjWvlsxQytpKFa
lsE/lFtVlimg/5Nh2UdQZr0DxZpCZh7yhlavp83jLD9cNNic8jytyI03ByebAHl/97u8ZPLTAml+
G9YsbMHGlPDS4jVy/kcivkPf413pDUum9BWOFZv7CS7CHG15awU5QpxkK9+GHugL9A0W8r+kmWMf
kZojGuP4IjZcNV+2wr14s791wDDacROlZiFcwhJerAbjx3SBobJfC5UVmGhn6dhY4JIdi+5o/kH6
TtQODm2Zuv21cnften8AC56oEbCDKRhb8zkkMUZAHtm6bRSUnvRS+SUaOxt7h43UZXp733FpoM8S
iRpMFlgpQN8lRQ524wT9PUIhQb/3BkKrjYlDP/OdIBk8bf7+6hQeo9pP9heKR8lS9eVMDkxOxgxL
PRq9lgbpixphewecJVIlif5moX8/QA8f7rj7bYp3YsE0i51/w7JL7BZeo+uKtDinfJQOUNsAA1+9
SEGEj4zYv/aDJ8WPMjT8DXMkFJYH/dzJbPt8JvQd9ZXCSfKb6QmYqnRy3U3nG+5hr7JQkDRnyJIH
fAgiXImS4ZLIRGXF/VLNv8dbBOSHt7tExfonVZWnYJywLuF/GOXnTsfYgX/XH5zPP28J/rLs18Vg
xC1gMT42fwACndy6Jr+DoY6X4XxSOdi2SfsIUrhgIuC1psWfneM/9PQQTRbDAJcfpW74sCG4zozO
Z7km0CZmEmdWqkb2HeCwmZTZdQbkBm/nmoNAvSPfS1cNUQ0AIGBWgkr2Rfr/Qou5RjI2QkALDsfY
lZ5fOwVP8AT8nRdSpSfkwKqloD93vj+ph5107UJQUHGInz95hsaaupmDWO4fLyhzNoQeFW9Hgik4
EGuQjYeuz6k/QDPJmK+4zphowcKMfKEhNk0rWxX2wv91oXfIVg8y5uXSYFavBEmivY1RSqoQJTwQ
Dsb9CljlhVcTAduFVIh91bC4IJ1k2nQ8nRFWlmY3BUqTQZEPEbqfMQGzbpgIXSBRH5evYKROJjHi
9/b06rCw8UWwohtE4CBi2nysBNuMCfoihbogH8cZI6cvIIsXT+NbQ0T5PujGhmTEOirjp/W8yjUa
g11FulJ79Vhr0H7NgFmLYVUKxA9pslSB4qvGoXsNOPzLx+IiZjtTP4IUmXskj0Xwh72+0wsXFNay
c6jIXuReB7p4N8AsO09jI9Z2P5Q6XV8cqZCQQlmwLP+k38A06sxQKTCACJm0cymPVdgbgYQyUMso
HWu+N4bVS2ocyoK1uWn/C5CC872lPl+lW/nFAGxteIG4TWXnrwykZHzITxN09kqwxQ7UHO85Hb1V
pyfAcJoA/YzMv6Bxi7Tol5IrunF9xMKCF26Gfgv3RTBfovzBCpFbe1LXwg+9Q+LvYM8yysfshomT
aeFGSD5HopgaGPB7lYfSbWohp/2cImQDI+r3b8w39A4Hn8ovMlsqmkVx6LmyikrWXjiJ0D+ZKkk9
BzIAz0+ytbEKuDYcACtwnL87j+MeF3PyHY5bbuh7ZuIfRQBrEGNMLHqDIiFX6X4S80Hozxrp5WWJ
W+xBy8KU3wvZfaSoAaFPunrIzQtNpVfw8lmPy5GcIWbzDbt3HbYeOWl4MFDJ9XDtwnoFFpsjmaYm
uY8oVLPK+835ZJYN1zlTJvon+2huAuaK2iw3tNH8whIG+zSdIjczflQdY02GzvNQSJPs4RvKQU8l
guzccv5P2V2Ovfruj82fyjCxNWjc/P4xZhNwM+YsKfbfxWzEcV2KsecP4FxsHtQH2wCCxsf3B4PV
ho7rrTeSKkjkRdSg/8XHSfjpO0jzYzhZozESAo4bEf+FpUUClzghklH+hLLvPs6c1wB10DO03Clm
Kfx2+rgBHzL6XIcGgNhkyZjgsxdoIAS2AFfHUI+nFQMt555p5LVse/zsjWQ0O2q7g42AQXIAuO+O
z3SNjPfx3PEdrNt1JrZTepFYNGbAZmSh2Nao0RJiNhrmBw7O2eiU/fk7oHoRA57IcUFG3eDj/Uoy
NG4KQ9GRp5hbkeSYOqRALNzoKrKS+5Xs4ieWkuXYPpO9FTvT0Yw/Xu26vZLkw6bZvspI+XEL8gil
u+XCIgevquIs7iR9mWqYMgXAvwqAdgpDQ07RoUAI0rWaXlpSuYO6p8i7plFWUoKVKyRisOp4+4Dg
P8CAY7CyT6IRyAS0Di5/OBPb8Jh/SOUpXE4JmfiU+i3IsB70lp9Mu5OybUXBPmuqK1aaeRFXhcCY
1HcIufyX5fp8MqFb+S3GbQ3V7TTg7fAYhyZl9IOIOdqCNGO0fCYarWCOLfe/DaVZ0uwwUD3LYQAc
VMgiwkVKJHukcLjpnOpeYMR3ghIaeU/y8oCuLcGEVHpDUjVETxPK4a87eeOjz4rhrb9fDisO0vRk
ti2xqbQJ1+ew6ws010RnjJH7iewfADrQQ2m3+vlzGRHb5/frWziLa9nV/foClIXzMFAhG3lUBeo5
PYJrLmM6Caw+GyqsNcxs60xtLlr8i3SXkMan6287oVV+JNsjQK7AxdltIO7RHeNCid2hG9azWEUa
V7Q4AkvcECLpg8qUvRv+Z6c/FB/ELCxfyMBC/ITfBnxxYZhigC3gzzhJ5Yv2Io0MKOH3PENAUchX
Q6DyMPqBlrhZf4g6gq1Vl360RmysY7lKfM4FHieW0qZT8pByqYa0XjCUWEoqNmgnsjsPUDvYDuFB
1eP6HScLQ81UEKKHNs9jmVwW378NWr34UYo1IxUrZspw73GRAl03gxE0tgJN1TmJJv7yc5tld4hf
NJ/OS4C0g1KjfU1lX2PEEsIcAT40aITmfaA8scJoMy5nbyN/QpGCwZkj9kbT+ZLaA0WumiHv4fBq
G2ZX4mufYle2M04642q5PmL/9Qc+t47fq8VnVkcYeeJyQezYhItpjrTRFhxJFgd6Os0YJx57dcib
pDwZDMG69bcQ56r+IhHjGFDC4DnphOENuFDYShitvq4vU0r/FFqlBvcbbOhrAu4uI/n+vufX4LZ0
wK5qq45VBmHXSe1mUKlP2t64T3ANU7xBsgFBTBRA8fSgzbdSIlAZHmMJgj89DL0m2RV8d1OepKNn
V371lMzhWf4FaHMMN7nlXlVoUxYhVM6w6vb/fsI7L6HNJ/YZnvjlnMzR0CV0Dpr98c/5w1qE0syk
yrIW5RBIaA6hpGBrRwBmzPNBqjXC4Uq2t46RB0M5pJze8TRqStO6GIwJEx4qQPo+dck82bJLKohU
pvqpLqBftbqtJzYswb6Fo9uZaHvm31fWAZptg+GdsJYLFZRuFd95H6U/IiCB21OJjAYQfv4b5brb
Pp08oytOkxBFmGXCvfsA3wrhyNfH30+Q1kPSv0/siPgAyoK9FaO/J0Kwpk8MhSdlytKwc/Y9QIqf
njnohh/JdRPKYysnYZZDNp1MLNP6Y40If5OZYiJCNP7n/sUcnbdKJCy+itWItAtmqmjsxZu4UKrI
SpJC5BLrnLqClECj4ntMdoZhzEb4rFNGmhzJZ3dT6iv+33RafeeKyvjYmLwc8HFP+wfGdOGb5895
HE7oZSCfxDk/CBwqcaLq0c0zAI1JFXO1+O3f1503CdHNDHIQPSDdIDsoueC637lrB1GaG4Ha7utI
7LLiC12pn7r7af5/zOVifv8CgOWJVDazBLDXgaaVlKop3irS0bKVJWRVypbHYKn7FpjSa36f44l7
+FvJFPoJqBbTbtdkTveKF36oyHd2ZbQiegYJbLvewKnregrkXB+A74oKJsEDgUIH2sKC7LBJiymi
U1Esv16Kg/wZrsPotgz/EMxV+U1IhdArSNRDpoMPM+xRXddNV1X163+HzHkiabGmzqmQKOz1Z86s
ODS7R4fP4MgmJwyIM8d0tyyVpV86AvCWvM+DYEPDw6sqHEf7lgWl2nPUX+yeimvGdZodvTc2lQAx
YN4URbNBEYOMIYUvjbsDfCFmn++BECQ6KXSl7Tq2xQrZA5QBL+gAinwi3PC46m0ub1JnlIRW1DGt
yzBs60mn80jMbys8DF4e4tMyAgOmJlhJl4VlGBfC+8wapptG2t4C+KJqhn+R/QCYXOpijSLrQhJv
6ZmPS5nKulPqh9Ej748XS9gGTNn0G1KZ1aNOhvuEvNy/wveoHB7zFc2o1GKag1zD4ej5WMgJJwfH
VWSjAmxKmrJub/waDNOTpniTZF5r5BvDsS6tCprrbk5XG6IxqSGklyvNYD9Eek2nfQXLJyY9wuNe
234nEqmKOtYRVIgO+MaJ14VEhAMrQ0w+QwoYwVH/mrvq6VpQ8aTXkYcyMSSc483ueObdreCtKu9u
ud7t2+97+vJ+MMOuB96JlyTySHO5pT7Xjt2cChoE5GsXOVMfo7scl6tFbFvRGZZ9u/3R1GhV5yvD
8W1vDHdVLbAGvEvJb+Evj1UtiLf5vngZQYojVOLOLcHuqZthIamHP0fCoStpjLMJ732Hr3NZmY+a
f1/xSOaCrNuHu5TlSTFmLrM+S0SNoQ2/BDXVN/IaC+GS0YeIq0eZU0doADR++tkesSTz9avCnBWc
FyL2UmO8a1H21BcSPdRj4jz6lrWdEyIg09NYfpQbzyEH432wLxeoRjPg3WB5+tJScDOVogqhsVyo
bYffTzYMlWn0rUM+njZ38ZX5NbC9KEQEhpaOieWSuZO+JCE+FoF6N2Tris7ogU2J+OcmJ6iUcUIy
/EpssW8yDXD+jfcoiEu2HfJRloeVcH3hFdUwq3OKJT/qbvkcmdrxOZYS2S5OsH/bzrpmGtoYMx8t
XYQwtQ/9Q/1qp2iVytxhsMtWNXgCf7+mLZ1NjczI9twKV3T2FKs5zB/2p6yfLIZr4ARaT4AVFMq7
qwX5lrM73dNVai+vL0+3M5XgSYNUvgThTHtEDCwo2xTtTKnH2IwlF8Ir8rUcqs2NfSpppYtxoqfn
4cdTYrlHG/Hu6QO7nv/Z3FoH6ympg+mIoyA1BSpsDsItjvk9CdmYfmlRngMpwhD7+Ec7VLl+Vq8o
PBrPIbg63Ym3CpAc9jufsvZ9TvfMl1v9WnGKMgNDADxZYEBtWDYeECfdioBnXxMs8h7rCCADAQLr
oYwbaGMDCnn0ZW3U9igOeHs9gYHe4c/XaHHfuuDwKLD12Eh9sz2uo2FgT2LL869OoN8tDk9Sjq69
P5sMg9O437bggABDx7AV3iFJzPOc+MJDiYcC2Plyrfe9td6+zt/iTNejoNx3nhVTIoy1XgWtSGZ/
uEsgQVRWP9gxRB3K1cE5WvVdO9yntWxlG5HiFF9AbtTvP3YdDdA361vU4jSGWlWXbX8YbpYY878f
qA07OE0Lt3r9w6WoE+0UDSX+qI8RWFVarbZbm8unwwGJ8rJ4oRUaL9jcUMHYNjzu9FBghNwtf4Ct
Pb5XFmY4MnapwZDRPEwS1Fpbo39qMohFLfXggsLOS6IU0zm2LGRT9y9H1/bYxDHpPasfVuxa3+o0
H0HPNEyAWhcOgJVIpeqQFaOp2lrh7mhpJWFSycHTfmywAjjaYPe3uaReXwc2PHOf7z6XfXsW6fFd
s3NYQ0Bu6okZQaA5UxnTbRoGwzlmXok3geOqzL/G4Md4LqBX7jGshcr9SHztLPWgNgKK9zBFvqop
8tEU7tMiJulVrvnZ3kiDhOXKzO8OAlavUHX1tF8ZwN+NFltVPiKK1xBYXhrfDE2LziPhVO/3McFN
wgmBm+AWIGzR+TdtQM2tOsYpDmdigz7Q3lLtMUycW/BJSQaaU24rVKOTLvnLN/QxTQzpp7NwiYh1
0Za6pknNUBEHmlAQx75OemkkDVS0cFuyaa77bxl/wTloh0BOXRpq9eghbSFLFutm8gmO7sPHgsN/
bPfq/FgCkAtqQWD439WHIhc8Ov3FDAo5T4TdjChVIwNDbDFP9v0dBKwnYqXuJSGFt/UYgiGqrGKr
eSaQQkTTmn/GIFHY9ybm3IQURks9mj9cdEkHwuhKKbBLnKw7392ujbBnuKkfRyAH8FQ3iaQ9XQBP
0EARX7srViDWYOOlHp0DxBV2HEbkl/zEWn6NYO3advh64UYOgzZIhDw0lbNO9SM5Em4PRXZ0EWSI
3pJIyAXO7oWl22ztQHB9B56dwUVOx3NDaB2JvWOEBsMKrbD9GCSQ58o3aO0xm8/XKhZn8cbFRT/e
vixduSO/qJzh9tBLqYaaea6GCa6+ZqbE4vxU5O8wtikl5NRNpww23DZ3TKVS9yaU13rHCBF6rq2c
WpyEZfLOl1D2GMosr3bGncW7b6zxSsbJsdflsAUa0IEjJTvnf/oUfct4hESOd5yt7TAdz3Iop0cg
HgdYY/qNENCHZHOpD5KOfoszbH3j4OoM09VnmjgjR/09Dqr8LycHejuP7CEU5zE/kOOJ5BP6f2P3
SqSs76yrvX/lQnDosaOQCNSdpbpEGNwxpzPBKfSsADw50cRfgCXqSbrz0GnN6gRT7AMldDlV8Z6s
SwAV/wfcdpTQTgVN0wZ3PqtEgdxAmYxqMT5zTOEESXauAhTerk6qT3z8SCCqiZyH2cbKZtxq0VY/
ikTIXe3usryQHMKKEme9+pW/ulcsLoy+GiPrBe7j0qtf4jIeA3e8NKwM5/c7sjVM3FhB0tUHhh1d
CNmuBwu0u2INBYK/M63PDK6LIUCgNFKrOc7mRldE+v6jpHiy/dD2iwwbjpFkQFaXIGEHtDBu3ODD
wtqXDsaQGHO/uFoZIdt8uGjHyPbj+H1W6W6SGGMz32h6AYTPrF7VGPpd43FFiA/qiRlvT7N6sCYS
/N/qsXz2aFQDeIogh6O8FIhYNT6BUB+z22mLlG2ACHzXKYpAxxZH0K1aaCUOp9Pm4UqQZPX8tDBV
vanB8Cdeq/1Pd5zTk0iXKeoiUh57871f3NET9NbvaMsNEJeUtpVmsd8ZPe6WboMaaH3yS3tSV1j/
qFP1j/NQiYDUZgtnn3WMuJcz6GUlb9vQtXAv3npyigvubKog4mGtcHPrwpk0fCebYW0tbx7CtIb9
jqvgcXUyd9r3uThA/9xG2vWUrw/Ou3+A9gqsQ9qsHGyU6exXHBuD3VEL8J8Gawr9P45T/Ki84luZ
RgPZNSMJGW/bH+e96kpxmzOrqoprPUwCZNYwiNWuFPpe76ZkW8I8qFGc7OG5ZIjf0Kq/Hn0BSl6s
8oi0F4eomE40SIxVlUeyD5vWl0fuXEZvFtDCw6Wz27uTKFjUThMBB9NJUCbciGvOEPFw/bcP2qft
nihCgLpq9AUf+MSUqQJrm3doXD7ZxhR8SY74xxUBRokV6uPSQj0H0byLrNzNdAAdjdBvASxkErT/
8w1ANjXmAEoNKvUe1q8jVHAWTZsnayfXky7eFwoxo8eziSQebljKyolv7Kn0zTL4yY4gCS1dp+lD
roRpGIpqBQ/1WmZTU9+ZvfxNKaWBtG13lGcjKYv02BUreXMvr2gOCs77V87HfpF5DAXJJIau/Maj
eMYRo5R99SYyECt8ZIkskUcfKGP3oevxtnGWx7YeOJGiaqOQuRSDRAeUjML/gPAiuEtmxm3b55DJ
hPPscCEpCWMCLE+h/rZVeoK3tkq7cZoDe0y13dpdA6BRKmPqCLJM0PD4YmeLgD8QvrOXFQ9QvYBe
lUd+MJa5mqHRYowOV2CaHe2vkB2uDB/3hL8ffiiteO5BG3zjHiD8xJMcjcPr2klymhLqEW+7F+Ln
Omo/k51qZeV+V8B4n4r5ePPSJLIU66Wbmox9wG+MzVLYckj+kc4+wwjxF3NDdUf/pDMUUQ1aTze1
LKlzQ7eSuaQIycJvyCBvEuuecxXPWUdihLymU6iNwWzMdA2fPbb0p0rzxR7XPJux+G2Ozk6laSwz
JbwRHiN1OjqQB7fwnmLhpBn9xn6VollUTJisqsN0VzxeRr1Jv4sZrAzbaJrviTI0JLoWh8n44n0X
ZkGJvbJAB/bBvXKHl2lEW1kNqReNRjdxVq5rNun8d2xMSryU3aQT1P3RsAJB5hgxQdmU443JRlpC
EkVL2Pj3dLAb7Fp4LkLdewV1Oi4K1+5xaATrRYcyXUguJqAwPK1vQcwmRcusyuDlDXCLnrRpyLtt
dpCGrHz3mu3p/t19SKRowd97nYtkrr9GSW6bBgX2By9ga+iOxH6VSWIRZI33RoBqCzPCRbmAkpUv
O4dNNab65IMcO54SG8yRIaA2q13Yoywp9oHQrL4Hncb2kMtwqvGBBWQ0ak5nOL9CNZAWlRP3bdev
pGFWZ/R1tQBoNcUwViFla3KDsbnD4g94m8UnclJC+cqZNPUfOAx7mTR41O8AQF6P+xkipPyr6b30
Y1PkEit/gpcSlucBBX0gBph53QlI26rRjbsMXx8UIt+jvyxS+31DocSa19UGhOoSNURsW/eugmXr
VWtxfCaVRP+wtjYkH9+22jRhcRwt8jtE8EKUQz5yignYbEh0PB8oNuvMrtSxtX1bi5T+Gfq7CgQQ
nqv2O+gt1bvqpGi855pc77j0MBwCYQbBRf1RKu7pWIlEpQ7UVRFg0/qzOYrggujVFqL1dyXI2r6h
magGY2GkCmzMUn2qO7TC5h1vHY1tdzHVcL/cDxyENi7mtxpS6/NWTcSKz/lO+E8UImRpK2hWswI0
NvqQ76VekJQ9nuEBDr4nj/uu5eWcGRiehHKl1mA1dJaT3lzll/CIhzNtHwLlJlvponUVseiJH7ii
WoFPTh0vSFVOTqbRWabUQUwdi+0gUviDdAVpxC4DxTi/bvPDwb55ZvyjDS9nuteupvyefeyGGtCp
ffo3RPvGcgdOkon5pbkLN9dK0etwYiwkv0zUP+5FZoC6tP/HPMvmiSHCadyzCvS9q1CBfoXhaThr
u9lECvYA8KC2boRVW6A4x0rXAemcKrEyMni1c85vK6K80hx5OjAvCzp1gjRL7cK13XVP9NBgT7zP
bn+idA+schKun8QEiJ58iemloeokfuX9igQc5nxUgE9ig7uiKYsgGObd52RBdhJLF9sbZb+tpZgY
dX059FkLFKIGkM5LOZVrc/dbnf3YDmziPrVQVHcFEnKMMpaFMdkSedcymD9uPSLN6qyoC5IoTAW9
XAWX28BfM+9oyStRe1u7kMiQf12w/NFmi2N7YG8FUwWN4zWvDIZNe8uzOKdx/JIwmAIqYIR5Egb8
w//mukKHjehEDDnTvAJZC9DGP3dEucaEqYAjsf1hi+LdrowNNfNc253Ca6U78hI8jcUTs827z8ZO
UABMxsprEFc/Wy0XmxUqZVG+ohMgr8h5VVq1k2dSKjWxj9tVQj4CuHbJxy7W6HkSGXwwf3cHS/0i
wwP5UBKTLgS04fzSAb3bfB5hQKowesWZAyBj8oHuYPSTmm+FiVh/MqubSufKsO28k8VSVgEsUmkb
b9PIRPYTsXG4YzYWsnkalloWiuonNJnS2Qnt+nliIjHNndbjFdidBPcmrPYJ6bcGEzJ9Xqb3f0zd
PNf9TM9GDm3mp+VsWQ6cQIyQoTiEXm11rYUAmo1dsyfCnZVrn9oNwkKp8swOt4jvefCiziNKivvL
j1TtyS+tJNDTl23loJ/DxT+Iyu5VqWEqw/N4h7cN4L1LhOcjg5mlUvJBCXuBBhXdbFEShW80IO7N
Kz8wa6gWe3zTF06u+eqlZiDdp2JMr740Jzm1nBANprJjHSLE0JNAztXpPvkO+2THEyrNOq0AcXJC
kRcr4kOJbIdj8uNAu69MCvA7BmVjiwM0IxiyRFRTISdGCQdEEQS9oDg6H0LH2G7OnHQah5zfuJMM
BGEUgrgmyfbkr3SNTdbXOiejoqLVpFnS9dDwTQAzZEZit0dnKKms6QkSvSIt5T92JA8Je0rHysln
Ah3s8QOedPIkt4PVq7RGo6vIho8A47xgR0Arl72AbILkEbrxOure3KZd37/M4Jtbc+ALf5F1p6p8
ryOTbd600Qj8+EIDzpniJ16kz+2rpOUPf0gZINf3lypu+zHOTJiWyygYFtUilbeBfLjC+Vtf31o7
9xXhF86Sw4peQqaGs4IlyQXN8s86vD5fKDO9gkYawZnymMzJ45dqyu/8KJMKKd63du1l0+QanFrB
dEXYcDvadcCunXWDuRVRhFruuBfessbYHgZDxocKCSaQr0K/yeeRnUXu083lig5AoUyY5V8iDVan
e/fkvPNlclJ3ftaFdw0f7cDsIWttQvDB6B2KOd+6eM75PsIUSrqfYHBX0PBwaXCtbEiqipdmT+M1
HZszigvU/eEd9F1a8iS8U7mAP60HPZvGD6drJ4Y8WDMmpoLHfg34mJx9foXrRgVU+yAaQx36r/eg
30fbbY0iqgx92y+fpNOkeBKZRRPfAKhatpI3eczhcKmNK7FZ8kAmWk5fxdIwAE+k6ulBbgnGeFTu
HLEsY6uvz2OFpIAz18HmKgxX6bdEPm+KVg5YVPYnL7RzJmcHJrYkNgcU5t6Icgiyww8dOPT2fLg8
FfSbnfodPFnFuSrZttiadW6NJRNkCsr09hTBN7yomHRNpyPxKnYSwxK/ILbmxoGa+n0l6XvyA9vc
MFKZK1CY+vLql9ObjGJoXnpmSeM2P4dHmmp/zk0wHPtfpUa3hrRGJ885OLNUNYrw6PCBNjHdLzv+
K2YC2Neeyqcq3feBLhE+LvxRfZuqXzbCyBhpFzHdkLHw6NihNLpol4cQzBR2XgrtsAVngIirrl2V
4lt1aSXrEK8nyWAIvhknzROiC/P0XJ996cV6GWDqqhgdG0nJyoWaWeWfGsjtTJYvNhbhn8Ax1QIx
rxrShV7wsGfHaUV0S1rRsYcdMiXrBIzPikeZiCeo5vjPN+5wXTcpUs0Jyb5seiVaMCtFFM6NeUAv
EY/Ssx++ZwnoHVarw4iRFrrsicp/akpfTQAokg9PzHNdgSGJAbHXLe8ZEWIhpcKa8dBdU31wUA4p
IeraJxTUdQwBgozCOYDwKeDNeOmqxKI1NSO1Rhp4YljRWdPavIMkQtDkb6icg7Ts7PUuRdXBjRbs
lg3dvVz5Rx+91rfhv3DTTcF77qk5jmydkMljNmhvTEjQtteh8dytfAOIsmQcdTspRvRlntZWSjgI
q2zGAeNjVyG8gPCdEk1KWL1VIkk1H23UqHPNIWelydEW1X/kmMDNp5MhJLRTymDj1PiBBT6WMHFe
ordJOdATt1uU5z+zrEdar6Uet9eRvtAXNANK0vrB0wtHsR1BQlMJdsUF1B/nP7pebEsHMmVu1FlJ
DrRxldKkg6Y4eX2qunGkcycx3x0zeJqN6XRym+yerOVnAZbHhpC83N6PAXROT6GysVpJ9bM9vSTc
GuGwJz0GGydvYhsiRifzjWcOkts8U7JjCMKSnzcvf62bi1JMs0UAO+ONBo/pb2/F8y+avWuHH6rE
Oz8dhL/bMKu90Y7H3/Jjl+XdqqzB0XGcu/iEmASo1yQ5+qT/mBqqBtYAurdRD/IhFUgH0zYGayIn
uVB5km/K2TnGGV32DWELit/vxGWg5iDem6/wz8o8jtxVQgHUInxuj4isoONS0+dIWIHJwNegWlma
F5GqEJzAyxoRutklAbwfx3uKgt3mBak7ogu3bcC6zLKgXHKDVUi2nRk3BE1Z6p3AmPF1fsbbkU3v
9ofW6SitDiyO+rxxUbtVEYl33dPBw3KQuATReZ5kKQQVjbq9CWZ4lHnsCgJ0WXjdYkw+IfGibska
gtvgnA7bu8ADJ/Z7gv3w2o3e//lpqwRc3a+NXxOWb8BKO6POCtZ6lnXE8vXZRuvUgSCyIrX4R52P
f+oWcAsN/hj3qVNeb18ToavB/NUYPGoIOuVJB0qLR0l+vG0vKyHT1J6qQdx3K5OpzUOZrdyvROxP
3/kFHrjktVngKZaz1Ook03W7WiQLeR9e102ZD0We6qhcXQlxIEPJ4mXquDtm9r/qWBN0lmhPcoCr
aie+luiRpaJ1twBLztzpakM8YP30/Ut9lWkuYRaY5Tk7exgHHsXtjE+Zbzc7nBEWvheOiuRmtoU7
aIThy70nMsSrMr2wqux+h8Qi/AUCWF4gkXAP3JGQ45sVZS/mRWRQGCzEqHqDtQ/t5rd2ucwUBaij
USUaXn2SCg9csRGjm8ccresJEq2J0lW/uVcNGBo2E+UiWM4W4kf6ZtAgNesWW5HGrBaT840Ytmwb
4SiVIg/wK2821GxVYS2FBsr47fJTtde56dGERFCNQw4AQOGwCNxfW9d/qf8fa7wmvkZrexLj3oF2
mQEivumBTOUvIhvAA5yj2iPJyVO48HgyhnakdSMMCffofpfVf+11FA0RBX7yb7TRtROMvMNk4l5D
WnszgtNmktPEZ7bYyDhh0Ks87pBMvXj6/nMIgs+1y5AWEZ8p45BrJK/hg3Gqexw5bThg0gQkvY39
cCn9TR1e58hoI9fj+0gbbf5Akzr40BFOmHSywMCjndtoWVXeR4kiYOmJtqnSnlCAWK/g2kcGZ8NF
ADF3eG2XmDF1Rmb12f1W4XOz3F5YkMf6copq0TAxC1vUwGikHQaOD8axDMDWndTgtle7WiwJY3Eb
qEkOyOBolo68/mYLm0RcKAGxchVmepM1p7upnG8rdQR6qJY9qeXZZm70YEBGXsty30/XGAgY+EDZ
8PSvpeUrXLsykVsREs6Zp/G+4aI4Yt7h03EuAM1CXXOs4/DTduTWHWaugMTlPqjSzCZqvSu5CKnH
62ngTTt4Pz8xzlozqO1NnEG057kWFmoRukc2Rs3OWYKVIy+tV/JRbGsaSP3M0uwEsyIsEzctbZBY
BqfFRsXcTHGCFk1KsYI4iYij5wbNlzfa/wNrt+L+wWnq+aR9x0SNaleonb18Z/TR1b18XI0eD7vC
YhjyTgWkGBV/O2C/3HUDdJdGU5deipe60YdPpz90TtlVBW1CjWD0tVkEMMmSXJJC43yUW+gK5gXf
qD9p8lqN+Pd+Q0uXTQ9FpJ221NtnmADvAmcv77BRippPycpjtYe9QOG5ITWTWQEej7DbUfC4LMq5
dPZVAGpVdPb7JoS11L3i/XIdlAudhNm4yEqyA8wkGpvFezn84XoNCNVUy3oJb02jl1uKVrPHw9zn
HoFFx+CNJUUzhVEr4B4XEVLDvhjX7zHYf83ljU96U7sVyOyYKwelXekwgrS/RrUME8UbfGrtAOIh
nz/wpYSxlPo5eozUH5x/cSDyXXF336p3+8CwZ4OMrbDXBnHpPrbWg7LveMlSR4AclmJgdHUMyk6Q
GuvEc9uIyDhewTT/fHg9UwMS/Rv0JPg0RcoCRD/qXM+YXsGDcBGs4krygX6C+mBtz29dJ452kXD8
ZwC4Q9WZ/M0jDlepBi3Gv+buBx/GQq1f4CJOTTyN1aLo4cAX9ibxopBZ+GjBHq6UWlp4bGbZIUyD
HBNn5dEuHSC7cq+K4JDhdTWtqigDUQCPGA+nWBxpXaZrtayz1PZmNkBm+zMb4onRCRikxAhHba5Z
j5Otl81+Pb570vUWHTu0J7zKpaAoSXlQNWTLtPs0xqhPYNbCaANqoMLjLWZcs0LbQPRTVPWuGJq6
4XkJ83PKG7hdDieAGd/5x6OO8nBP+wUpxRB8sv9GVKP8OBLdy+eJpHyf4vmRhrDVTIXG3OGLHmUl
pQFAkO6qpk5lmzSLmG7VEOcPuIexLlDj4K2B5WvnEQ/LcDvkKLvv/D2p7q3AxvKqCgjb52MX88rH
+lREVu6FH5gfROjSyA6fpS2QeFtR9Xnp41yVawM+Vu1LRc4d+n9wUwh4ajwHBQ9AbrYWvrXAUdt8
nzqxjwjPBBcER+Mfo/isCM7WTOStnhqagfUfBI29Thc1/SQGKj8e0BE20SGE1aYFsME/3Gzmek4M
glPIUGtZd18pNwj7Euhr3323mIkP7kru20VPwx8YDNx0ba09PiHzgvtMUjkfYZ6jF728XaUlYExx
lrCobuJsK4hi8VsYBXWwJ3hP79QKlmufyEmDMn/a9OrrgWSU9xeXyEmXMwkvF3JHaEJAg+9aMVlV
2Z7Mjwh4f3G3qz6059AFNXXVin7pEcvT75pInm5Psfti+iU5lOL/sEyq35xbjj4q9DgPgy8tAIcT
oPht+qO2EFCGzf6HPDLY80oLcsYjz/YzI4aRGmEhX5o2F0ke9W7zvWOjMDqLbRgcWyZaxlF+7wn9
2ZqSUH7zRbK9G/Bshmyok1tTS/wC5BnvGwyDbkxn7rtBFzmbW1PA3OS/Iglc0xGpL3pLMweMwrpe
6HEhJCtum93LQN1ZxXU0FAakl6n4pZOEZ3E828uRzxLEHQ8AR0Au4AzwNXWix/f3fENm+P/cSkZI
vngtGjkm67qfrfCwkz4ZiPo3Fsa8IYwdPDnbAimbjx8zJfSi3J9Rba833pLxw5JdFdSwzZoJ+WJQ
Is9HXO5Iq+GMeaImHK9IwTJt7zkjZ9ddKzhcgsXGdl0MOM5plzLwi7+c26w48EaglB7i9ksrsnHS
JFbML2XuNWyfStMbALqLRiNHIMPKiXeHxIiTPHbYUjU2EfYJiDzeBZGURLeHmCRhJNbyjNqPE3dP
nzDpQt4iR7MWCTED6sjwfZdEYz8GfBHhIoOCx4WxYs8o0T8ZyxO5oAOg5KMh+B4T6oAHLdQosnIo
da7jT99sKSnIWIpTu/0LtAVCtVsjOMaasnR3Jr6gu+Rx28vmO7PgydWPkDd4cXWF4AdO60V+rkTC
ji/SXuL2Y6MG7l6TqjFb9vNLik8cvq/sIM38qq2emPGx9n0twu/LCxTH2UpoLba6C6Lo8IYpsp8n
TM+GJvC/XpJc4Sus1hZ2jEKlugruTWnlXR7TOxUGqV4OtVkYv54ppR38wXGh1hV6LjCsXWrNtxC6
+wig8+1hr075PgtIl06KkoQBx6Jh0KKgdGk6S3MqjMtNrLpbDm6A3J38aInjQLcSsejQCmzvzhaH
mBAkHHwfGN+vN/poptn9/7d0P58HUpoPbukfPEmOUm+Kr64LJ3g0KB5jjP4OEhx9gUOpKjTNHB1L
yYMgiE46aM7PotU3RkjDni/vKeTfAYM3awEwhmzCEKn4IoIMEkoBU9UoEYjbFVFmtyJWsB8PaSs3
sMQ2G3wlq4hpx1kHBnx4UX1ozDb5rknkIka7CDnEBGES29Dud6Ifcl5DzZ3b8iCVomOYS3XvXaro
P8C+/VmgUreICNWSVo2oS2z6NL4MBkqQ6DDsZcz+n6eFep+kiQyu/fkKisJxMcoELkveHtIJr+s4
R+ekd6NZmyuH6FPELoQqrq3YeXL/Eh+/i4//a67v72pRk/mbE+t3EohoBpQd8SPrwttsLx1lICAZ
v+sjGFdFvrTtCjG5hWXRsw5pIEGHGvz2XorImngjHhTeJ0hx2gQ3ONfh/GbjK9DDqgJHCml9HUnL
9uI31r7iEMbRjXI/aqrbDCmqu/kQILUQNvCX8HGg6dUIYaDXxBBnDcT0ZnnIf08OXuNDgVhpu0tw
O6IdaJ4cSdeJurNKW44cycVhOlDfqzhadq7RWv8Qls5JLe94mXmZvzjtkcTlTRWh2Suvk65jFkJA
y1DAWMPhLhYRe7lWygSvSpptTVp0ARxAy/7K6O8zrOcIU6vgYBmXQrXDpGcwlFoIYJxQhEoemKJq
KJoMSmkYwQrwAjm25FfxwbVXLjtLHv/AjBlXdPPjFvngyPMLmNaTjsaxXTUjbjV+XmJAajCPvbfn
uht2JCxTm4LkhcCieVcQZRrOXVnb2BXSLT583cdZAsY65+leVtzqWHhzUnHK1dAIKa1FA4nO23Qk
pfHXF4pbyvmq2+w3LmjRNdLVrv7QVVvc332VW2DdaOBXj0rHz19MU3LR2lWwuYjXYYBlBDdu8+dP
7JL38ukW62bwyUWQzCRNDWq/jMSHu08s6bv7l6ctYoExVXT+uKTjxktTsW1VBFakYAr9CXmpBph9
vtMs3lVO6o8UdEEXXPaZWI1yGne87BJXA83G4ghc3MMbEVFV2a62SvV3b4Yk+tF10Wtje2Ei+fS0
wmj/DNuSJdrEZC9fK5H4eP2ossoj7m3Zaa70o4Y3BYBlxPzwHq9aMEtLj2WlcxOflokWuQSQMwjM
xfoPybHVVw+E4/h9QMdjqYBZ+VPZXn+0zz1vIUyjceobMrc8pSfpdW7bKM6Dd6Xk7JOu/YheCr7D
bSiVuZYICBjwzHAnvIWKrAWzOLYWHheIaDK8vVxJFYZjF1FrY107+iQmfbaqRuLMUVNjoQ+pjkNj
e2l39jih9aU0x95GD9UTBdkutfEuUw1uf2C2HgR8KsGibWUA37Spf6SdU1cs3djXCLaa504aiyvx
UwCPX5QybFlXgX1dr7Gf4KetXw7yCLGstOAc7KYTaCAyT8byYupElCJIDRzQ9D4gN+Aw3l8tK/KM
645ceolxiYt8fLwdvrNTdm3OH0lhFiD+f5un50Kc3Z250jNt8lbf6u7dYu7DNnzE3HFkk7NDYKZX
dLDmloEdiQI2cc3FNN+umo/RgSZTO+BkWHu4Xg1D+UQu+tja9XxD3OR6GvEKSjWFYIEtT9+9hi5E
92QsYFPzPl7209KSb946dyQcjbR35DvZvTTuJKcrAckgrcJZ9DR+jf2jfcTfhcev9KXQuEumFdS3
Rt7AbRNRlS5C6SQNo2Z1W6qvDMG85QGOHgMwJ4yGaZ+U7LwGemj89Xd4c35d9T6eameQK8y8yjln
a038HFXpPee+Da8yFiu10mylG+IZ1YBE/SbAlXGPozu1uiBVpY+4rAjJrH2fqzNsGoIYkDMVRak3
13OLg1qs7B2FKtFEXeh0Ua0adrwv5EZPc/6y1heOxU1fj/q8uiPtzzbuB9uinqoUzSighQ0FBNb5
/qdT7tDk2ELWnE6CzfE2XRqwP3Pd3WdCPEzT4h6D5Tx8Eb75g+nl4vgBd/gIf4Ilt8Ib61xqeL6A
pMSRA7Z0wfIGNVfsBOm3L3mTCLwUvEAlCsGn/c9um9DZNX+lCUWjAqyFJmQP2n67tPOytnI7hZgr
sM3RrFuiN5VTMoYuv/TrJL3J32Ms//T+vBGvE11fXUr7LiJfBnxm8McvIcYkPbHzRohzx5OB4Hfr
QyFeeyGLDaezxkUWjqQSXdOQAvOIFx0vTmEbC7KQTTdvZuG+e/AAsXc8fx8xU7HnZG0DqfzmNtyJ
MTWNVPFGEZcrB+he28dWzfAQl7JJ5nfMVGoQDIJEz4bc497Wix4liFzTUsTsRVgKI1Z1YM63LVcv
HVuXBzQeAO+2B7NRIKr4t2/jJr2AL8YYLoFXZ+NQ7oL2xz96ANOz/792zCNsJliN0Qqz82pPkDBa
W46FYCXpndJmHFo0nWImgFH/88EUUy2A2dn5CdYeXd8neHV4XTqxqbyqpr3bsqcensDnfJMRaSbS
qhyAV+oAzGcKVBPtr4jMm76iMPTRa6NgMqg/Tr1IBbtdFYpCG+SM1CqN3dfkQy85fYZElR1pxdLh
1LGiZgihZNAp/VDWNQwe5yJi4R37xHErmJ9HEzctNNdb9YRpluImNpBGTNhKhIboJgYoLeGhLdCH
khAUTXwT9QdzhUVkElQamBSoujnu9sNWyeYAndvUuwBoR5+w0g9pOzsv6PXWMd5sRHePY4jd8rJB
XbT8PiTkGjZqyt3rBeGKScaFj3VYUJV48IglJfoQ9UOTWZuLOcw71MU6sW5PZQfru5UD8v286lVf
HZMBvqp6riPwYfsvo0wHGwSHDj2lEHHoYvSvIgzA8+GaSmqOzh7lkUG+lUEAQI0G8dfly3EZMhu/
2Z2xuLjB5VRiBZyk52/znjpeGzDxweTXz+et4AUUmjaBVKmxjw82DMNFfQEJff/KrxcOH2/HLUuV
vpiWt/X+DJJohI2Aojf+0vdOx7isIQiSGfFMGpb/TF9hLfoPSg72usyOxmGyei4P9xu4BxU374tB
WT/PD76DCEmn/zwaQOEGQA//SAEGUGomlBVBEHpM15r9gGSF9BtQtUYwNpQjxxCUE13MVnBuXtdU
apaLsKQTKYH7yWMiJBvXEFrc0zSfZNis3SUpfcyYVvsInJBE6bj3dOJ9IsibADID+he9aNwtHez8
K0UI6y/W2oXWRJZXv6pdS4oi+FVF7J4GGZU70FZ8EkWK57gB3MsWC/u8zrbyA5OM+oIJXFuv+Ua7
6OAj6JAtbHaWxUViiKFZDgC8pIPORgFiKPJ/7VfJeM8LZy3P4fgXwOXCWpNkr1G9muJEncBEt0Fz
keLl7hdbUXiXn9o4jguKQg2hFS/7LtlMYAMfFA48N5vJSoe9kTb5B2mRpfTG2mQmxAxyuXEGySgh
BLc+2xwu21ZVWhfrbwND6PLl2y2icOE+5iqz5AxZ1ZhX6bIiWO4FOD1KobIUVkwJFfZvvETHX7jl
c5tRfVE3ExmyzuqrSOpqMjxn6Ngv3BcHjxjTCUDzRR8nGPsX5KNd3KYVycxoGwbO8CrqbVjy14nF
2E3PcDu9VT0eAo6R/i249655EuCv9lu8JiMH1dT/Cc3lzO3hrzSevnjnUrs2hlN0xz6qqnA4U7EB
RKV5te1WBBZYh8MqfFlyQ9uWUjkFTyfT+6S34FIazkLbE4JHnFrrtr5Cc0MDxESxY6iJ9aZM7lXd
1bgMdzTjdUFIKyT2qJhI2O5sdCMXkc9MbKqp6kw7+lR//pFNCYGk0Zw1JsbxtVhTVpr26TxrXguM
KkJA9BqDVIvABb9fcVLt8yP4kp9arvytbqzKIeCXM+XgtK9ACYlGGKmFsofjn6RuSJPdCzQlFU5g
fB+lToI1ZJpwWRFMOYHFo0v/6Okj4Qr1dk8/MvbSErwcVlm6RAC/SNDmHR/JgjC+MOx787A0Flf0
YbDUDfGQwlH5l0HndjhPqLZIA4ok2TwXmNv83diNoGGd/SUnrpqDpzsPGQG/lvX7P2bUQj+LvsZE
766KZqNdvi+nmbkN7Pc8xfaBsqz9khrqhuHL7lzX1t4SWup6miy48fND3nocgcXyzeXM3+3U5EZB
vZfK85yWziAFcO637AzzYnVQlJ2YHMUTlCZMBbqw/da7RAD8SdICaPORai05i14b3DEIKKukdK7q
a53eUDNlriXITeEvfovrYLMuR+tf9sR+kOyP6fYtKqAVFC412tIJ8tvoDXdVqPHtv3na01FSqEHd
C7pCXWBGcksrnF4sPT5R6TfsIW98Uhu3eV2PW++Phi6rUZSe5BUY6XYeB6Phlz5O9ySBdnhzlUnK
jonuUGMjPYCeF8iWYophWXStkknejgmeOR5TxKZJPuw70nS/FU50f9opb30ySyLulS+t1jnXho9S
ncwWijETzaP63DksyHDpS+9xyQ5wMa2DnKCFSPuX8bwGKgiZFGEkMf4cPBJtEPL0xL+SUL2L354u
c1GngiB0JwZyBF41iJj25QGMvDRTnXQfPhDfNdvA9VvOYdea9jRoTTcEdqeDj2VzgpFU054MIsud
upqLtYt95S3vrz6KrwU4uCnNvGCPXLD6athFACuYuaQImRZJvqSyL/XR3/QKdfL2QIAnlOefc7Hw
+9vqkE2152et6jeDEGdWo/xg2gs4Wu2QWcGXIqbqI8rjYWXK7MIFOWOFHIQSTsDrxT6NeIsX3Xqw
s8Ytkvcf9byN5O2/joNTPcsD09j5ND6wgLFdve6yolfrjMgKhnZ+ZxVJjMyPlUX2QG+rapA7O/ot
bYqFj/e76M1/FnCpJYBOXe+0sN8Gvk+qsetj0r+mTdorav5Az0AtJuvRWx49qO4wiZYKNV5WhS6a
bDs/f1lewDRdNb5WOKuahBSR/+NcllQiOn4/Rp7W8c0go3ASwztAVS4noUFs69x0JlnSMSzpN2qU
FINdpf6PqyeIW/COtDPYCInJu3x6+oqcy+w8FGoP7IV48ADNhlsDVa/UpAkZ+GPowgrt5hzuP6bJ
NV+05//w6C4J/vmz6Ztxn6fJW4IEg2AWEynjVxGHChKVcngb0Bz1V1PS5Xt9DQrK61hfopNvR6P4
3fWF0493z+i48CE+5mkQJlfpE0fJBW7uIbtYSgWkq50niiII83wASGSZIFSLB1fqGpBVC5hh0ego
PvRjW4jWoQNSwSganSf1mal99BYZtSGRebt5C+FbsjeRQUwsUwlHBg4ooibienZ94uc9Xgxj55jb
n2lDimeVEpyfdoBcsgCqsHMlzUT4dFGWiLAsRZ++2IVDOO9r0/WDHXZ3ydxhAt1U0U6RkqKFnP/l
nTbFPws7Dfvs8oSaxD2AtSu/Fnp7wWISIBXHdLGSBAniEluWOt1nwkASou7WrgiMJzoF9m3PMZg4
hvjchC+N7tvfQAhvRbGDzJ2LsErvlJrH9nt5/fuOs9bSvu5Adra7+4B7mVW5yfGpvJ2QpMpG4f7E
lHz9uZyMx5sPYif0ij3ILfAuR7VMHUmlDyyg/DbxI61dYMsj1oOeI9MMrou0/QUVlCxlPVjTDyY4
xlSNTL97Mc4wsfxQ7jawYz8eH3aRPQZGpfXxpIrSePq1XONKipOWeJWX/Xp3iqlnsnWh81AUyLZy
4lE4T/MJWAENL1TzRqtX2FqAKPU853xQj6dMmpcfesKWdErQwgluZDndfvTaYBotIWprukXv8YUJ
qzkb7l1JL+eHR8CnGKqFSjooggAy4ZOle4/XhYOtifP/Jz7Y6WobaT5OqPBIXXkJTadnWZ45oXRD
3zT2o9riKvtjKXGQwd70/bc2CugIaCRTe4gWzeHJD5dICTjRrKZxj9qd3kwrqvzGOV49+p1OapOF
iBijnsQx1oL1RqiuU7TpetRqerjI3TqM1rAYP55Y9T0p6crlpw9kYnr9Mguzmnj4dUtgN9ZLZOyx
wwrsBS5lB+Jtvv//tg5OflMRFfvl28iq64AFS4ORrfRcusndmavBSlThzq+3NM5NeHk72c7vAA6j
xNzbEAoTGt3+sYdgAI+4Oi9cJVicXjJ2m7ZBZAMccYER4T2hQ6+M7LwJuTOljfmntWQRZUwxS+2c
krA2Tfgdas5ttlwP3pJxuz5P1RyY5E6UcHnbtvY5BFNkwee178ENE2fjxANo/SricB5SnMhHAVEz
dJK+pSoF+9Yz24Sr4rbDo3Hg1nLmdklBY+B72cHv0sxwKXeIU6hRnWFR899C5I0z7JjESB/GU4Nx
YPzZ0WdxR6SP18wId5d/Nx+dyzknss94TBSa4tw3RlEGDkaL576iP8pfS7zWi9A/XS3yr5kN9736
rm959yyfqJkv8XefO/L6EqD9EZfSETYWkP16CcEIVi93IhQ4ThFYaFvSyAG2cqJB133yC2GmPiKI
c7XYDG6tg7Jsmu7ai6v3t8DKli1QuoT3Ph2NfOKodQixN3zEA0dCXGKBo6VFvWi0LuDf6lkjhYfD
8tiXWFdvpN4S5nL9zUQi98YXSdGTEPmVpO7a/H+Y+sFjrsa35mn5vnEn9++dLy42X7JElfNQBZEa
zocSoOwqoQBjMTS57PXwMX1rd3x61wIEX89/nwxyGiwYQRx8j+UDrlhf4Gut1LkzvZIDcmgfksCe
FmOjJoglNQRrUKuhxYp0HYAoHU9sM7rib0rkJAy03R+bIbpNdKztrwo8QczXRkJYAI+kEQ9irm0M
Czmj/QxU2fv0DODVF3UHPeSolY2sMRokUjXn3tangPzThoPdIdRlwUdQXuPQRqouX4E8JUuR92VU
77XTXnVzWzEs2D1e0cqK12K3TMwqgLkufXBecZ4tqs/d4bl0MhouPihKiyWUed/EVG3vQAcTo18z
HGqGRfQLUHGyZh01x+PDnVDV3GDDpcVjxsfcSmHxK9WJhBrOTcaFnDVRUlJ0YE8hY9cqwxbWeVXK
d2Di83RZM0c3M4dNoKEvTS74alBPedmwK9hET2h591Jn4qZyqL3TuJFwQbkeoPz+77yAW+nqzWye
IsqF0GHZFZK1Vsx5+UJNjHIDQKtcHlsC6XFxtFyao9gT62dyu9jAxhTOLfNakezfkntsLAfUdF8J
3er4y7236r7JJcKHNd8lN7yedDYQ7BOTvJSAar6QRUo3FDoaQujjvrTYyHuvhFy8vATIHXfm4/vI
aeTrsIvZ75cNBBV8jtrAWcHZ8rpxDmPIk5it78FX/pfqv6m4TZTK24GOv6onSExUWit5AVH5FlLh
zZ2vrakAQqi3jS8j/7CAOQCxnXALrKdrrMm6xzJ3ueuAPVd5y9z1j5feleL6WzmdjKu/Zsj8NsRE
zc/HXzFczkAB9OrONrHU4QF9biAIfjpYWWONChzyHq7C1MahkM5nypcSrbod2pNOCiaqaJM75fYC
LsQlAVuEEbmHiE+MU2splC/qhS3VudCytGnWQHASST/j6gOnjZlof3qLEikgynueBwgn3bGG8XbX
6KTbKQUjstuAwzhFALlwVBkOByhzvhAOVGfHtGKJl+BCvSVyZdvhspzgy35RVyhaBNXlSJCsl844
mzDpTZUes+Q9ft6pKCxXgw7dqo+rx9DTtVfX3X3YBvbXMQ+PXwPgdOm2a8RspvIC7YdyouVLUBJd
7q4n7ZkdtkTR1sTwYqI8KK1mDUPsSWou+Tt29HsKg0ZcU381y8KJlN8crtOd9HRqq0iqzhs5UyRB
UFGFjqlB2Pm0u2QL2aP+mhCYOh45Y1FHRWYqEAF1WkjrdJXJ0lCDMAkoToM2p+pQjbnbe2NqohHS
vC5JVVBVdLjGg4DFVPIYbTJytoDSR+6nHYFkm7FWSFLcqIVek9PmN/ejpWu861FxXu9WUIEBwx8e
2EEBhPNq/qkhiE768tP/E4ruQ7w0pt4HL8kkPjfP/SToiXcPmYMoNo1GZTIghjlamlRpq5ativj+
h/xczSodmkSSi2yG+JW1p2M6tUvFNeVS9LFSKCfqqmf9buBfjjRlfN5YQtCKJqlBEWqWdcNfZmO8
gYuq2bsz07KR8DtxO9KVP8JeXoLmVyPrL41AcKs9jp7Vlq/Y/AuAqY4rA9ng8cZtt6QLQiMfwfvt
Sq3PP31HK8IunA7j9O4e14D3Gbyj/PRQxIxHlB/86ctqBT2iUqfI3zQMcur7FGLI47qmGwnggd7P
t9ROERhINAv/3YSHnq0M/09kauthpdhMhoQ7L+VfuGiRFvUd/hMdvDsWhD6sEf1fWG0J54OG+ptA
vHcaaNZsQHXMoCOtFvGuu0n4Nr3daeCP86FzIzHw+mfHcK0dx2HfuzsFfQlunjKu5aPL5r6K7sNR
THpFY07m2zFeopJm9mR9L2YqolMScwT5wj8iJLf+qit2D9pN529qcBTB2lYEP7a8aCaQDfk0mHE5
wwrc2dxVfg95h/6VmgHfrVlYkEvfPuYVdqJ73MY/tjGczYzj6S2vtj7c3UXm1Hs8xBW/gtupWk9c
YRcl93JfLURzgnlWwOzmsbBUl9GV3HAVkRTn1/sfiifjotLh+oeTXyq4KilTWF/oxqRlrYR9BEuZ
OOYYiGrLifVkqnp62vXroAsJFHjYIyv0CBl12h0jEh0j/qwvDNCD+tywWWiY3XQE6GA6LMqXKhWc
e8tYBMu0EMf5mLMfxntcutXZ91pL7P/wS6mWfnR3NdDmIz3WORmt4SQBevDzqADK1uawenZN50HU
jruGxuhXTq7C7hoEoQG0bqdtV3hcmdo8LbGJ8YiwOL/wI6BfzqZqqGV8sNBtEFs5C1FIHno3haR+
ArZeZdOtAZU5stNRk6NCCUI0F4T+7JPFjwl8od5JIVEM+JxiTHYL/UqyhokvOYvb5DpxcNjy2k7s
YXNuPp/a46yNpzclpsss5N8OvFluHBFWbK0AawugEaa9PmSR/fKvAmx0ns7UMeyRJrk6ibDkUpMM
ujCwpuso1WJE7j4clRmNcCAUWYl9NY4/yBIhw6KjJxDzCfpQgXsck2uKA+2Bpo8NWMrvlQ/fqQE3
3MwuTCtAhcb4/VabhBnKVsR8+k6SR9TYIVDJGHda59TBS3I4A51Q+aQ7oYLxBCcz2615zlkgTYcq
czbirPnau5c64TNp7tQIjkA0svUHN2eOdaT6MllmVCf2ErOvItCaR+xZY4yjuzPMrgTUF+g/6Lz6
Q7YAJV2W7bWhZwIdWxv+8H6FRyTXCYcOwNETwOFuPA8WJamGEUY5+wlUexWxCYIiAgEKKplD6247
Nmwg7tQPjez76qyv+fZXHDG5mHeMUM87wbCUKIro088afsfB3k+7a57vIdEwUd5UHtiibGN/aTz+
2wSSvsIirRasc2oxOBYXeog9dyTBi66B7EKzkVILULgnh4jtrNIZHqxRkJJ73jzVJGUmQwTUIKIS
EInDLWubDEGXvuL2Mw7pX96Pr77iXYVDWhBIzMRJf1VMsrJXrrOzYVaEZQCGHcMtIgLRPQB/YsF2
Vpnb9l5FBIjjoKVtMdp+hoR2CuyhdzHD+AIH0z1HHmhzV65G3vt5FYdCoAHaD0tHGWxiNIrZNwtc
3LVJi75yKk3+rkJEME3g4FZbIWtqJuMVIYwEl31me1eyepFTW+gG97jdQN1UrzO7Ir5rYFHVFCrw
Z6yf/EoB5nT8eTdOlFPLbfpYT3ZS4WVEol5zYfTuxhMhpJnDIQYJ4rpsrx9U6PZapT8UJxr/STMV
gKPzF8JQ7+MkuZVcB/4/sQARlgJgoO19iJSb3jLSacDBXzIfti4Vx2Z9qE+IVHCOxXZLBzmI/et6
Y1SRnASVRenRAtZJDY1XhIrbw0TK672oYL3V/Ayv/NWbSKM1QqHPdK9I3JlnWvSQTxpbyZsXIj9L
UvVOy9bWdf/AcmWLFIYHCyl1Mojkos0Zf5LYlhoj66Ruf+M5TCZDqZZl9dzim6J+NNwyZwawa00N
0cKH1oyFJVeTcmr7CpKpLtz11MD92rYnEDVI+dAUM6uJHHgRI4pilI8GUowgenwCz+Y/rzEsiL9O
Xr8KBMY4g08+2NKbGGY2ww8j3f7cQEwS1Msj3ZcgXgFcJnLPpyv/xfjF48UOOruIVHT5xYejDNyo
HhNB+fPP5f1eSfHhpfSlxXB8p7MuukfTy3uNbWCACw5rkVx8h/9qycz6RHSYaVCV6uhB5AssD/Dv
M75CfjG9ackOOREAnaV+Vqrpldpmx+/CEm6FpIY/HDhTFD/fdFBgdpbcj7ZNI44ksddOJRDIuBeJ
waqtPMZyTqOERf21aUupS7cm+n4EIHK2L/d3SR0aEUJvJznMKMtvnH7pI21ZZpH5Mq7+O73VkXWF
Tx564Kid+Y8PdHVtISYxiCeBKOJepwhG1jmrHnCszGJgiNdhM8CO8sqRFbMUDLXtPMB0AHSdtmkR
v98S8oVD1c4Ucgd+SN5psrlLJEvywOKQ+m6G6+whN+Z88xvJT4/7VtaBHdntt+bxE1MkpjpZivuM
Zuo2kpQAUnefk3Zvcz+FWJNnK18WEO3bsdPXZ3XDEyQ43uqH557jvapvHo4JicLrJ80GPh9JHO/W
BX+Ls5yCKvHTaULD+sfBwBcSxhdWh6qsji3wbFkXgpIO/FwZRhx3un1UgdUgaBrZOf1LaWiNwsPL
9qQw3XJgg6S1f3TAnGZhrGw8Dr8yunEhdHJXRxQXJZgY/ggE3FTqBHzImQrgrwecatA+axOLTswB
SUJkxuV2Le91grUNFg1I2RUvGHxy+65kl/A3Vq1G1GYhVNE/D45YwOxuPCDq+5WCzuLGdW4LBH57
jUP0zFPQgMtFhY1UBC1U+UJPsgMEfHic+i+xq7PYjwWAJVWuMf47G9IEGsAQ9Y8gwlfXeACWPLXW
+LSuYVe7fTt5RBqY67lGlfVw7AfcpzLzaKC2bxF+00Zyz/NEFJZhW1tAgP3c8MefFYUgoQzJaIJ2
PMPwTqgZtwJdaoQaEDUYAFJEwCp57DAgq2uw26y/mnMbFb2Aup9Ah1wx6nwz/r3IWWacokrlvZpl
/vR7ZhPRMwkteume6kfxCj9a3i02uJzF3H4PZoft8+HTYeC7GI80qnyhcPvfSCUGizZSvjXwBnn/
2rPfEBd1fr9CQKp+KkBj+DvsDTL4eVn2xQuUqkwb/W2Czd8d2+GAWMJsQGk4Mhk1W1qPs1UVBA6T
PcKojoQmUWd9vp7wnzdBaGsTOkXLN9DEy6uvwxPWGQJhpQqKZ/iDd9Xfw5kKy2OgoSBRAQPq1ZuQ
0nWOQrkwMjNDpdMttUh0xnaTy4V4LAmlvjOlnUg9sQhU8hSmhCuJ4Wzu04tt+TD505XAqocWRB5I
kIPjmz81j+ua9hblVzy41Szx8TDCPay428wqyMiEG20CzYtIUuzM1HRozjoQktEZaxZ96awJBCpC
oDA9YzGl91ojlCkgPzX4pYvct7sdSi7UNz/5JIz+CRbIvUyJCq1QGP2ky57XUf0nXJjYgtaEdI4a
jGL9hO71TJc//IM9WpW8vRC+QNpZ5ofHKwKQ28ms6QLgTm5EfRbGfBJcMzBlg7Oz30MZIenD6TWI
LdVGRJFgugiBmhyWlUv+ZH7QIzPuNDvHvgVLSwMV4SL6yKIUuOSQgDl3rcQ5OfvHgy2SdwVWlgan
J88wlKE/pg2PyQcVOSJ+wqHZJiKEIxGbeRNmjH+qVms2gJOjlCUi9krgJG/+FsMnkRFLfS0rR2WL
xl6wzD560lg60iTPlIBZ6K4Ku+Ng9Al/YxPCmv+kcBNA1xuLzH4HCYG13v27ghzTuYXG1IDTsn7M
OB6ioQsK2zuEyTCZ01l+fJiOo35S1qbU4v3V6ZmNbprIHp7NwtS8TPaYhTXUY5Qi2HYEx8Vt8sIH
an8iJuQNP/zAmlZseuxZgdbw163ZvfrtMTtezYVT0ccThnWpIA4AyeE+GDhc3adRjZB+WjN9bw1/
fq20/zbvQ0xDkTP/UY1EGxTbLqniieOkDp8cgYREMPLU9yKUyegTj45slpTKesSSmT1VRj1mQXOy
TbaA1uVY4LWvIFdy4otvpPGCTeg0Wu9pmyuqmQIxZNHYx6xpXb4PbZN7AwDDFfjaaTcjTdcsy2+p
aeYsz+5l3o39jOu5JBNS1tG00yOdJ0VJqa3SLJnqIl8GiU03mrj1Z2UeTJUxSo71+TRcMgtgA9b4
Dwd1FVrVplLprAQEowFXKpUULfNR741DcHAUd6cE1Tsf/fY/ess+DznnzmEWNIvGLZDCEoSuRLS7
DbiZpXWpVMHoHnOLwsFwG7/oaHuwauOLfD3MBmsHi5frO7BuAn6IUke9kzQgTq5Ms4Giay5Z0LYF
1qVanviMPdF9Fwgr0Lh1pM46xLDawGGqquyJTkb+yq7Fmyi71Hv+zdkKCZxci8jf+5ZWE2GAb6gw
dmu8Lve3+R2yW5uMrrT9BQZBWdgWAwYJVlPncPkqciItjURZLfop6r2esaDnI7ez4ycMVJ3MBsiB
05W0SNd4wDa94PE6XdcEil0RIuNeVp45ppfUVeg2NvjEKx9KzrUIKnjL4X0QsdJn75GG+X1mLNhq
kL24s1JxEbHK4HMpfxBOqypm2cPMKDgrLteRoGlvADFchIeGXE+5THLu+GWGtMpWmT1X6pzi+wtE
l2UMutNJfXaqr+Ay5y2uRQlhAJy0O71q7JcvT9UPSujoSGh/v9ogPPSWth8tqHKjXCKYHEFTjLZn
ROQc25cABBYmZ4TkX9JeF2kmtmR6AF0fOtfB6WXZlhBiyTi3miPqFE/uoNmeUIRt7ZPG+d6jjz8D
CwNJvaQc096q00wuWBUJzJU1WI2xuXjJIH34DXy58+YRlClON/mBQysN51F/qk8DijZEgqvRxl3Q
30cvAe5RbiXwJpDc0d26m2fBOVA/DbHw6ZBgMPQOTzD4hd6iUijFb4msMRYeBBOn9oKCNuMI/Smx
o1dSBbnVprKnokx9ar+ivnLjh/eq1pQF4bkyhtGCBme7nZYtxL/m1to7c4bOLGTh/+fFLBd5N/gH
LRtMwvP3G29U0CIIRj+pfQQdbZGGbfNAPwwGy9qt7vV7CXm7Yn7lnXXN1gpAEEin74yY9uSityKR
ESoUquv+6R38YRcvcQ2l39ieToGxgDtmMYoNSyasA1pG1MZgbOQAV1USG9p695ZhZz+zhdDX11fm
Mh+yi4L4uSElTRHnLVhNr5t8I5yjJSJnF+7oxayS+oddMuiO6OG2g6HhmJxoa1uZkMtsuGGQscov
XGX+jcNS/UuQYgBRUr++bR1ljNCQeAl2v6tC/LRWQjvekzzTomZjuvJYv3GEL7VanQwvK2IyM8fz
vBik7FZ7Aq8ylQ2zEPSAJVr2Vxe5bfPYyd0FAyUR5GtIDzcAV1OQdVN14nKIuuQ7mzrkOplS48EG
DPDejwHfBz+dfD6LNVv507ewggSG3fJtaePM2MgQ6UiauiOkMi/hi6WlpSBqXz7DDLI0wJXsVtoh
ifsY33MRgEI6dgyIs7gNolQChM9FcXEMBkvM5ogKowkQmRTC6AiLKpkIoN/Xu+BTJKxAlgfmDlDQ
XOMFl0uYJmRlqJyCM6v8ok5KNTBjWrQGHyblmaQYJ6E4EJ81Fp+AYwbRKGOGR8r/lp15osyyjmX5
DKSX+Z8hQEh/jyTu5h1wDAmH2thKWTH+zTyl99z6ov6/R/J753zJLZkLeR/ciX2qC7no195d068F
s5wBOZuzsA65RCmC6V3wlgrsM2ukwNhQudw1mvjUk3Cp3eKKM5JbuuRqCNhzaBJh7Hpe1EX907Rd
3cxk7ezfvQednbDEGoZwq8CGOp0KqlaERwCk9G6BWII1B6c1w5OhrTZ1nIV77wzW6AtFc27GlbQL
FEHMOAlCydWqC+CDcTHBgvuiFSx9i2FZ4me+UnC5N1ma3E1/uzxiiR5UraIVpKMeVnLfqFOrG2m6
HrKa2m7pX0VvzkXE6dHOP8PwjRJWbXkL8SCsXMGk9jyYNLsc0QwWjO8omCWXG0ur0yExAkcHJhgz
qbLmc3G85yT9J6AiU67/4H3rbwv5o8umy6ugJE+LqgM5WKwKB461goHks1okQI6qG7KI1aAJYh4U
9DVAiniLmkOOPHcEpnAPfSSR3W23vcJOAcyP5kI9MI459gjvDvEFnVsbKIMdkve8S4X/UWnfzq1Z
2fT2v9CtbBgQgfhE/AcGNEto/RCJ1aorVeiJA2VGpn20t7yOH6/gqL33RXqFqITbZARHllPF1PCG
stu0KkCptzlVSmnVQOiQ+V5p0I3N+fPMxztgr5Uit2cciuocDyyxfgJISZYIzPTfwcCXgqaW5jsX
mt8gj8o1vV3PUtys3OqDdATAFmpx/EYmCGLs8EbfgbYy2OxHYBjxe8lZY0rytSuuBlgeA2lz312Z
k0z6JicZoXYEHV3feU2GteyUZMoZXU1vj6y6oadmS9NXuSkT77eRyo6irHoOHTYcNhM5MZd0A0rD
k5kEx2WL2jBzP3DlqV4hA9W+tSinMGWB54Ba1L3nUkxpK0aLHyySc8zOX37zvtMG0kCqYRoLmE/9
+tfXW/kWV6jEcNTMlC20DQtNLWP9Ym3FW3q9sz3XiT5nE3w8TOFbEAHhahx9lnDc1EXa7RyxjnSS
Ak1j5ZReTYqcIGQspXWKa5ICmNFGXnU2xbFOnebud2OF4Xe5gSNuw+4MMGpdCbiwAjWEjkXMu9Xe
vtTsoqfGhkXUTxYuQUHnLOIV5/1igp4qeMVGPJrcl0Mzh0hDtfspI+UhWidPgZPJSzreaGgfgGGh
GYsquikRBC78DRFFE3CoiG/fcRJoyesLss1D3TDCnhLPK//oglFCnqPh4/REKCkg1bnUu6E+uO63
RIByi/JXucv32QygdfjQ54x+V2IVAwLZ64bg3Lq5ajOTv7Hhmrfb6yrpQAfeZ9DYwyLzoaL2yzaK
zPkLgY/2J+qu0vM5Yl3r/IrNCTWVdvdvOGXnAzPTZgLONMMqrkUVBPOKA2M/owIywD791GykuX+l
voiReo/i4P+NuChFOI9KdslHJluAWmOZx/YMt9vrCR+aTjNsEj7/KQdAe0tIK8mzKgj3xgX5Yikt
K98zv+aFR/gziuZYVDuPd+YCoUyWHI9i0esI4CJ72aQhngs4fC3JDNcYUpngRp5MhzyINQqIKm0H
mZ2AGeskTr/AyPVlMEYSTp4Lkp3W5jrq06dhg9kvPh5h9ZnPs88Ao+6uZoYQevHfTeoqHe4DdD0z
9WPFfj0VZFFYGiPF9qxWJqOINsrkYzwO11lV3NS8bmTbNVXCIfAL1W2O6lvmToj8QimV7+V0/sms
HQrHfpiH2z4bdFdBYqQA+cyYaUYmniKZWvuFujxuzeUzMyqs8N+j4xxEWmNag+5LioycGZD8AF+y
4eVwH+vel5KXrTW165Y5HlI4UD3C+SqYLVrCu/YvJ6uYWe6XCZhKo/75bgTpoZEqFmBr4I4bwyc4
lMEDIrPF/7WVQ3Tq0JlT6um5cJKX/0KMMOph+lQyvtXq+MDD/XoyeFvaJg4Far9z3H9ptiQUFeFX
cEy3CZEUdi8SoUm7q33Via6ud/dCxuxA7Ng1kKi2ENayeU7YeVfMy7GKxrrj9L5u4lmKsk/WJKIV
V3M/7iheY9ZWCwB3ALs7qjbSfyYD2bsp2FCq1P+YHQjTRdUNuWx6WtTg4XFo3HgGg/jXZ6dO949y
DEK3Bje+YAv5KaLLprPW9WthWQxitQsrWlY7KaV8pqlJiMDKvWgg1T/X8RQ2+RgtXu1L8FCy/9Jg
8lC4LV9TQxGASZYT0iuSu3iyH1RqleDb5m/nP7w33o201j4toPKtSk7m5FkA1jcF+cWI2GiivCFv
53MgbiBwPTDi50lXRN8pG1PWv9AuhPWr2rugRyA1HZ0pfjYrxjBL5oJlfcr4rxHQO21DiPpes4xf
ZP74qoxVoIMDYDCKjA60/dN5EJx+FQ4iORgAqYjo8selNMkgZtIgv1aWq7Jc2M3tCAAGMEys/x7N
MbUFJi8R6+/JLBsSQ8/yNE0h2oAERpgqkiaDkDJT0B83OOqX22F1hucNKBN7YYb3dYZf6JlNq/XR
SdHZkGq3mtaZh09lQ03fLyVpO042t3h0Ha3GpGEPeOm+lmG9CB+GdWZSOycUZAcZ7pk7ukl1zxFd
l0cmn3AIhvGgLE3HoM0kNpIf3WxXB9qQzPbDA5PsKxvbpu3h6TqTIhXgr65uDSRDr9xn5HHRFtex
w1DfyoauuQD6uUYGhynf+ZwrxLPDixHZwoqOwskXmCu5vb7xSTrof36QiPswTnyArfiH2vp0bcHn
GksSm3J/AhojURCaNDtgogKv4QmnU4vIja/Jw29qVW+cZO8cs/2lWsJ6pRhLJG4HN6NojDQ8xQmW
dG4ZWSqmFuysXMui+vVCV4vkhkBawY2uftzKpS1heB7sijcId4TQ2pWlbcOHV4zijFuZM3vmkre7
wEtGPkzIIbFTeB7pCVJp8bsSX7Eb9dw/vYqoZh0WjLja6ecaG9Na3K/GhzWj4mKu56N+14gick15
OjOcV/v7Fk780DWeLZ8vmzvsQQK5iYnbeKb4lt5iZfnixCNYva+oAtnlOWCSz2wOW3d8T0cgHUMc
csjYPHDHcldfbI8OLkxCO2RXnNBKjnRK5H+u9OfKcif4Tr28vl/1hWcespvHAojfYxo1qlGTmu8D
VTBUjxoPT3lZ6wWC7jyHcS6uhBTiX5OGi1u4JoQBlvYr+m0FLFQR3XKLzl1dRc098b7KQ+f3+ta+
KfH7Fv28hd20R87+ub3EL/GhZJQKRvU24Ylq7fU6ZpTOasEqxbDPfiCCGyN7gKVqwUaF+kH4R+c/
zMUStscOxHwGtDfNdgdXXgzb3IldDLpSrBN23gpqC4DHoBYqJ8i7YUjQfjAYZ/WV6fnadocG1oTR
4jVllxWkLH3EJTv25y5Ua7mE8HTsT7Kg/SLtqwLyZIAAtyllbSgGPULSKxi42Ih/s6+drBD3Ofuk
A6JT/cdW+Jb8P7hkgB0+reO5nso7zl5NbBFyIdtWChlmiLdycWVojs2WO51Dk5YKLfcmp2fTKQlZ
KraA+1+zV1BEfg5ATkz6pZD3OYdQKqG8xKGwf4UPXqPok+2cSWTM//DmU88wpgEqckM9+F78x7S4
lDoOjyCqSSFPdKuUjzgQKShVSC4lLJStlc3dZW7w8I9yETyTmkkQcviuGquffRi/NsmQIiEVzWaq
JnB/zEWAKsFJPPEOOnbzgSbRBSw+L4bnX4zwCoNTWXgPyXtrTRuoOiHkxx43X5+/0478LSGhdyud
Q6u8+FnlMHKQqTlsDhcaeVl7WYI1j7dJyRkB8rmpXcQOihtOiFtrM5K0mIXIPWw41Bg8vdU0q2Gl
HN9VxwGnXEFv2HQxde5HCYyxqsyHvFBsRNRzm59unyPLDipNP8PcJYAaU3LxKhAkBjosIKPWIlRu
EiSgtqiFOiEV8IrEvls+yeyhY8j69g47S1D9Rk6rymx6QDKyBQM1+2Mkdfa7wq0bZDfJgVbnRXmb
J//kgqgc8SUROQ5y0S6WLvq5M95SiYgEjO9pqxe4YuniWqaT2k5UJDPEjdOz6gGyVRcbPgNySxZK
rLTlxKJZT3HnJ4Wz14ru6nrcZH/OaDgad7FWIsOBkh6YIKoJzAXWFaN7XloW5CiR1XbOgfjeRh56
sMJAFYS/Mk1smeDQk7b84YL/yVfCxPIfmyhqstqUTg5yWhsZMzqc+tjn53QrdFu4B8ObGbBPzgT4
BrxqvzexZJXjL6s/YKVTaTkIcAQW2BgzlIiBTF4UDw218up4Z/EBcoHgGjQ78pga3jodm6ijdxBe
5n+mfDgn3KlvdsfHMmqDa0E3/m1UEnxOSNn+pMAhwBYiOrz1wkhm+qQ09i+RICmFkovnUFaS1aaT
a0Gs+KBZm3gsvED+0RqnLuonmYcChN3pmMbdC1e1yEINLGAkqXh6I0p2A012+XQjtN+6a0LSS+d+
ZjnrWtjEbVaJN47Bbxx3xT92KcTFngYalsKWtI3OdvIAdrQkdcw3Izl7waqZbAp3RDQRUMLko5Pp
a0rCs3iQ0j+HRYK3bVGYsCM9C7Ligdm2vlp2zcW0u6lrv9pS88Co3+DcDyPc6dYj5CYvN7Dk3qPd
a525+uppni3K8bNqMclKhmA/tLV0i6e6vUi5U6p96nJW0Zu4Ja3KuOI7PSdlj/NFM/CXwy7boxb/
LtrvWbtQrPhKkL52QEJlZo5USGxfyQEDfGF78QdjJp0mVjfq1PxjvcRpiJ4ohaLqWjUfVm0CEP0I
9M2+vdi3KBMC+I4OIWmrb9+lNlTAPzUlPlhV6ICpV/vfhGvSrbb69u/4A+jF/lu+h7TFFR7pw99v
jyin80W/wzzWC/ymtBxqXF+9mFc2gGM2q8VkyoiwqNVwMAMc1pO630uWHNNC1HU5RCmYCqNSWM2b
NEf8ljxUgCOIvnmiO0ftUwUZtI2P038x+HZQGnL4i3+XZHy8ITmeiDGK/lDUo8hAtQVB2cq0cCzG
F7NqImWA2RBGSMYXjG7T7JTQrYtNXRbhDQdLghlfvHa9vghlf54nEWuih6nbqdNF5rLgRdPwPeGp
W3gJbI64cA1qkVEm72kJrqlygTL3qXUW0K/gRxQ6H4gNWcRmQTs3YDrTMgHs0he4CPikF3GjhOPX
97iSDbo2kSYdt1qlVL5Lohs472HgBttxpMvh+tqdD/Oied82PY3jNn7o6fO4sgRrSrVoE9s7aCwN
OHuwJpVDLxJKL9V65fUTVS5wSAbq9ZA2bhDdG/qrl1VkY0YLoynrOdKRRx3LZGLo1YjAC5qm6q22
/z1pIkrAH3Gvee9W2neAaoCJjDy0s5xn+ux3IGwpu987/1fi+jkc+96R4d+SSIniujtLsKbvGGeI
Mv/6LSniDpqVH+brRzPrOh7q0lT9MUgeTigVNkzrEwIb2gOAbqoFTqidk3bVnHsEV7FgnYNlZj9g
XV+8jL3i0aYeJeJGpvQLEg52TuNCFPt2RqQKdQa4ujfyOR+tvbpK6ZmcGgRU3NAQQlyANaSdhu2o
WcrPjPthXb7ga+7mlAVLyqLxRXQltM2yagE4quehxuIq/Wk2ntszLoWID5YL+1pG2XnT9JM5J1Fd
IKfbdmcJhrf+gYTopboY/NT8v5SRH5GjIprPk30HqtfGkVXF8xxuwrMYjH8SmbtwvCTk15hMAlxN
y82HIiNh9Un8KTRDpCatKefwou3+QvhYWxYuiSlKt6EfklipuKIlIzels3eWvO1AjXfD0EUEfLAo
cxqfR8xHk0jBnFmKjfefHmq1LgQQpeKLOZxWfQBNqvmfcLogo4xvi4l4GGJfjgYSk5p6AnxwuTLO
fC/qd3aJwLO8d9rA1Dta+6fKX4NTSvLkmoUXJWcqxis/LwvU6+RE/MP4y80wrIvS/aY7/TJ1t1k/
H88iEtfHjhQmSrHcG7Sl+86wkOrYDDty3wU2ZgYXqMyJpPa8x47dtLQ8hHdlqG1F4bhx78S/dpRs
e3+cluF0G1Ti0dR78b8JtXKw+ZqyUv16IxDdeyO9QEhksa+wcDyDCeIHK88r/6/8anESrJoWpM1K
sHQwcWtZ8lqbDJuwTgh1yVZcnigVtk5mgcbK0oEGP71eYJhKfcgaRJzI3F7Ch/qm9wIvu8brSeP9
RD7D+IECkQ881t6wXiNMe8P6o6iTIJYCf7XSPb+V5xCA93Lmt/Gn7AaH6JOlbHhUVhb+V7gY+uZ6
uldipeq3e+hOz4G9xacWiI199hZZyheM2m0pushrzuQVOcnlW/zezAuI0GmN3YLe9LKctCRNbTgW
5DiZNaODzOSYYHSGAUFTX6g8TR8vEueo813d09S/YaAmc3SLoBCF3l3UkW9yhnjOQ/3ozA+7M6b5
dX7daO+mvb3v8T/XD+lGjpzEuDt7PAqMPLrfZoghY0HtccQIFpRP3FADmNrwzbQERfAQAW3yRumV
W2kduowK53utywXaYke0RQdSxJ8Y9B5xqnPmS2Ycluecg9AhgHAxK7zB5jQpfalEtuPa3O0Dz71F
t0qi3AxT+x6klR3y2oB8/VGytOz2muSMzyabs7DgIfYBk8EN5UFIE1fjaF+pjmRLH5L3moAQX8oc
Kr8n3qF4uo5xGMOdIVh47GyK97mEaF5xSMB+/RI16cC0FYqZ0fP7E8LunBGbJTSYbiKXAbyZHaa3
Vu/LBdAyzXdzW0TnqdAoaXaNMGOND5Y5dN6MUZg51rhnz3JLDw7VNpIhnaX7FNO7Ibxh9E+aLiEg
2gvsus509ZJmQfqz2U+4UwmKZnVXEftrpJgb+gE2TbgpBhl8F78+5uSOgUDXLp7YrpMnXlZYYSVr
iREQPYbDGYLamSCa42I7OmntsQWr8p2UpHaQx7P11KRT7YujvSDj0zr8ERjnwqGxM2tb3WR4QNxU
yyW+Rp7iMzRF2xtRljQH96iBbp52evLiUfASFDaUND2YGbuuIBpxhIFbP0P4YyoN72SEgQxNlN3x
OEcvN9AiNObhprWPqOi8zBW3PlM4ooU3DaupEZC9CbGX60vgz5b/BDKszk3aWgt93NqsOeIF312I
hLVeqlllLUNvim7CLHvJf4sefV1xoGWFNiE5tFDEWG7lF2aYzFqyZAXo9idA7ysbdrU3ZobjHy5d
oYji8AdBqv91IVIN4hdqx8psCH7mRsEGJ60gZ8vY78Q3oldF3hTCgrrd2LD5Zq3Nd/5ee5GGgT8I
zx2U/DoWvyhn3P39EnhnPxhnLwbaChMmmi43LvHs6/QmFOErnk5QLR5mRBmw3bF7oCl03mPLNwg+
JftDdYD7sSNQfamRqSVTePN4sl6mnx2GvKG7CTT6XkMMF6NCQg8//c7qcCPTaL2c3te8hqdG1tA+
eXOqTRS+oK5vjz3Bbv6fFVnRHfJh53SzB30TS4pYGV7swTYWP7CFeUu4Zx2UUnZYeJsi+OoFiVxF
UD13EZsGrP64W3cHQWEf6FrroqlwXxosBCA9MrRr3twMeSkEH/306jier2s5xNIteYQ0leBLosqz
9gmz2E/adjY7YkOzJ5MXhYTZOZUs8z/L9cFjJTkGgLEVNRkgqEy9rxebYSjozRo6HMrm583mAeun
ecALWkOSxErL91zn5qSQyqSODo7/QU9hzY8QKCl0DzWEmTdWimE/IsEd9ubFFmrxVsQXJ6QzgK+n
xAP7mIY3L2wHFY0bnEY6ovvvzZdcmHhg+iYCMZ1pzqhXhguUaej6HmhnUniuU6Tmg1EZoqUJY5MR
UkzDwaBDarVwjCF3i5Oj8tuFzJ9zH5s53MsDSA4kkcfxGQgeSrzsL7bvrLSXh0EQLuiYUD65iL7F
JeT5he3XvFGxMw1c7YbVkSlGfhUJ0cNs3QmbymZzDJ5W74fBpJ8eC+M5k+ySTMwVKW0AqtkygGOf
PF2Ggf3O9ObNngqEoYhwriZJ8Zmf4qkyW2xwcKdGSGypWpbsKwK8sp3Y65A6iRV3hKfTlHPxWp2v
i7EhIELEEMNv8omR3kmcPs0PDLrir5+hCagk01LmLe8DYshY+CzXDSAr+e1EphzMrRxHKKaWR7lq
QedfjB5ONTAdv7tNauoWa8y7puIlayiIysrml4zJpFFKoyODxsdpJugBWducN9s1JGEyH5noZnQI
k2PY69/STf2dRJelPA6RHv8G+I0JImH39YrfOtvrxpujKreZAikvUmumbqoH5k3hyIgYiO90hFG3
LA+J5VWUA0J9UDBT5T+WFJlWRQtf90VHSUoNshnph2syB5qsleJiXQFImPt4g7vDpQBo0GS3Ew1H
zXlI2At8hXyI4SpyCqSji3Fu2R3qTN8dhgfE53p3z/GzONOqzTFi6QdlJ4s1Erc3ZM++6soSAVTV
d8mmoKwGxUcrZStFKf2UjuHLk4sEtfaU+QKelmR+mWGjubPBDwqXy8hqJQgmajC5hy8jT9yvmUyc
x6Ky5rtGufWmvMTYtUHG8YKEly7qpbVr3+OyGTDZt38aw0Dw5NX3BXa5mGTFGPAM18qw+By028wH
9Qwy77qq6M1RcDgXfe66K/al2jE9XTxwhPkGbC8STy2KBt4ajC8edseQSVuv5IhUk1V4Rr04t9h9
vYGpsaX0FXRRSsDIWI4bXAAXjaenJZxEE0h4sXOS+w8+nDNzH5ed1X0Gj5mbmb1voc0MDJWubmlB
evnPlJsYvtJ8yJ1rD4PuT2P9iXt6qj1DZDeo2fcwc77TGQpmFwPSlJXkfFmdLsCVdvEndOb4rUlp
ieE6S8dNJ0m9jaiCvC6fPu/xGNnZlLdu/rK0Jhpuld3cwCuR02SXVxuRfkKz96IOUKa+fBP2HA9J
mPYt0lQ1MddNSwoWMSsIRDnhYinSPns1snE/fJSm8NB3MgWxmHhdU9iSAQ3XziPS0vLC92JTRM/I
otwwUF721PzHVS0/eYmhrAcn5Gvhj7v3RpYbHIITUfuJh34BRhvCi7izBHHUZe2XJUvK95aR6JgA
W0MiypZsec1Ds52fOZa1ziebXvCzXM75mtfsLHLmIS3XvyryaSqrqlbK0kwDFRam18S9c8mKLQHX
OoIFfIeyj3RxN0a7+Y4OlPJxIV67l9Vu5qDoDONzD0dRhvW3w+xBcyieLda3Iv6ikNWA5HAmwATT
u1pCyuM/ZfujnC/NqMs3hRMhuEcRiFq2KQZhs+mHWaoLKrm6zutkzZs1qIijwzptVCi1Frue6THU
NaeSZFm7mGts2CFhewQaL0Hq/jUKtGanm2MN7n7FG9CfzLpH1lN/kIQwh3MgVbum8n54hDHawkjS
EV6qsPYxaCWo/7TV7g4CYs+xdnX3DoYyYFPvrUdRPkT7KMk3LDQ8l51Lt4OKTwfkN8k8z6RUwylD
Ls/YH00OVm71z6G5SIO0BhHQkT6vtubaZASZs+T76zU/bGjhSdJir2WnQnVQPg7APWDXKM22z6AS
KPFLzHB+rDOsLxM2s//CE1OJxaoBdpwVZfICvcg3ztqjsg4b/YFuENrY46ZXT/eI69X73vs7lZBn
TGNPWt35O8nxP6eWHE21adAcOweJ/mtpO0OLueQI3tQhzp3X7FLOaqEQEBxuO7RTThGCcaVh10ih
QCtequH48Wd7JoB+Sn9KZ3B0qUHjM3wuufH98yrr+l/1INh377Xovrgj2wPetYA0FFp8FuGnndw5
VcwtnLKlWumnvtXxz1/3p6YNlMa2lzP3w7Vw3ZVl+KRBuDlPPZjbZ18t1YHwvFJfFaHFmBHa27I2
VTQ5gx/ZcWkIvcUj4cIwb6oz3UIALsjWi1D3RuTtLvxOJI3zSGZ2qMD0ZmFZdYnR/e4kRDwUi1Bo
wAu0yG2v3LHznyMWqz7ieObhjhTzpIcFD7bREqH0OG9/qjHrA6aQVHlcuTIs5btcgOCaxYEs4mFk
9ALTwRZQD12iq226CLzwJ49mqOHOqS1+mKg1l6TAFJfS9JVbPqE+tGdaaeaaDgu2TWrdjm1OFwmZ
LvYGJW6IfNkwKTfxg5SJtwU2dFHkKQvIwGj2xqlRZojCduXhKxodTZ8yQwf011ylPw0wxET6sVaA
omk0CHE7YSiXjd45CCtIce2bWGtbt9jp/qak8u8rusXqB9eEcf3fkjKtIjdIxHVkinCdFZblTejU
BeTwEudB5K86hEP1Arx3PZTnR5yCty26cFz8zq7hzyWSXH9x1vJ2saTFEfLxrzHleyG0SzwHr8k7
b+05tYuf719CowwI2S+vbQif/x863nthFLzRroXINTTtkBXKkYKIrL6KKtt8NQQO6KEa9if6EDxQ
Us1hY6BMJy44RXZ1+0gcZltoixYU8ZPwqT3oCVOD9oAFGkhpgAIonXzIE3ujq4np6YUGsSdpOLs0
ISNoOnvLFQXU/UREjvRqtN349DN4FWR+b6Ut0SSwq50IJFwTv/s/qsdVz4MGgrbfjKaGpUEItHX0
ya+cH9hrSNYRfv9fPiKaFDS+bhOAaX1jJ8Dou0h741TWp8MdgAGYI9Sds/bePQM2QTOf/FS75gTT
lNQE3SoqF57b/30TG4vdCDZ2LJUhsyNFzAuwC/67p21/VNFZ8FxhIIkh+qpKtShIQgALMU8Fl5jP
K9YQl4WSZzCU+HyJwiprSMxo7sKA2hvP3h1k9mp74fUmw4a9RRowJH4cU2HfxlHvWisE4J0ijVN7
aIO+YeVv870sXgrOrb/eTQe9j4lveoTqrILoe0KWjEXFJyddONJkiPwzSp9lZX5UFri9zKQcKKVt
XLAf8n5FYt4bi8z6lODVsLzgttBX7q25SWyf5R/quFSff9GQMYmi2Gz0wF7M9FKbdjoUocI5u1lB
3ML7nl70Cu6/jimm48nC8HDH+sM/7IbwGS9kU/PG/IR+ugQL7wMjr/3/hF0M8C2ehAdPL/N0eCkB
2vs6W0kWzSpRpVjyQBbRYN8YWecZPHHmZwrFz13ag3HkW3HD4PjUUUePDWA1K7uTNSi1F9RMRaiv
ymUaLk8b4Agfl8cK4pZvj+1S42SPgMf/D9f7QLKWXQSgwhCz9Pa9VinpiwJWPw7F5eFSLtzdiA9k
zcb8e09gqcQUTVcHwWmvnpqT+2WvaT9FllIVnlq5IA17FZ4/uezhVnJhbg9z7MgtfBIgiePG20ax
5ptnmLIhNs9X7O1sFGHUrYu0ag0s0MKFc3Ioab9B9HLcY/I5x2FRVJY6/2YtIOKC0kVuS9atyF4T
7B5V91pc9FQ/flFS6EY1rVb7/LuL5bjiIeT7a+ifab2lpRcSlFWIcplGoubNVzPD6rHMsc9p2RPj
c7/0+a05nAL8q9MFcxQV8HK45l0WDVxSdGkpAK9BD3wVkQ01N9PLmqQTC2Rv9tbpjw2nnsMIiuVR
A8KKUbiolJnq3wx+ig+z4GsJy1pKdypDL9Dv1PJ/dJ56LBNvoqXVyxpCF6Jox+jaSkeFa5XQjQhl
JUOAhg60u4GrnCEAviAupslTW7N7ifSHVR/0RGQp85e78gladPJsjgLHiFTEe1qPb5jryRfIGq7z
mK0wSJFFW6r0XaxFBEPMz60yHSCWwJIRlUY6io1/wCqyUuuTCpgLOmmNHYNcK3F0z/z9ljvywdy9
0j3znwQYvvRpzhBC1wdfzCSiPxx8zgLKJOYSs7BsJToU9KzQOJdO2W14qa9ftIATPOrVYUWwHam8
3EHy3fmf2v6eRN6LGpr3NqBAhTAnK/CUjzSlis8TJj1NyynPJMG9ZPT90+TLKYnN3PtP7fQTJPem
1/yCuZLG5/rHBYmp3D1RZcFAlJAXzDJgBVweDFe7A0aRfcdeFCvNrE9DIBm9odO7aRsm2AMYn44j
f06jtrYBQr/6fsq/h9yd31Ciz6ZS6A52XdEgsQ2pMu9cP/MNt+4LD1kvWyp+bYqq53Yf6xtmGyXd
R9GVb2/kDSw5Sd7YJaRjysH4E2VhTKVMZUHx2fbZVWQP7ClWj0spkVIVvj/jHUdmM0M0wtDvjvqF
y1NPtj4Vge7/h3FfSS6kL5FumbEPPdyQUTt8wXH8i3uTAV+vhHRwgzkOh7RWEo2cIas+FdEFupT1
LQIlqZEfagJMietYmvjhJaWzXHYszUNuI8EXXzeafs4yy+jJhEUaWxnnVRBEI9EbSMVFVBXuZXcQ
wISVZxBD6eJs/5cPSTVRxSsUpCTCBPRcaIqIhVAsZnnvxDcl6LD54Aa/scixyNEu4a0cEE1Gby5Z
bl0RbQM/A5SCaYyFzKeju2FDwPUAhlWkYLhSaHhigwxTbjAI8q3/81x4oTC4UOXfTkqwYULc+Zoj
558UKcVYmRxH+quNknzG5RBm4I1u8vELEx0XtxrqAN3xqDy4Nsh+Moc1kgWsbvvc7cXWo5NXxdSk
amO7FjtgX036ir60KEsGcGqSswgzgD4NYQCm7B6pybxdnZB7bm9k3EMtvmjGukkENgf5/NLkZicy
X47bW/G6Nc7x2a2I3Ot+J137UiIRkm471LG76eEQVe3Dsr5PS5X8taYfCluCcgMP5jbf+LDDtmG+
VhmvcyIqWiviGdSgwDS9mwhm9rHKyy0G2hKWr98Xird500XF1Lka5+vZHxhBAXTyaDg9mqNGP+f5
gDReAazh+QheW3lfyzgdYovZrdc/9Afva1GmGlFrKycxuSxiIEMXSxNMcR5OZr5wUpfptugQ3mSS
BCC73xbGGCvPhmPcf6YK8sKJJnUht0vu0D8lYiUIxv7+EnehHBfqV/nTwp2hTKW3pZMBYCbdzmtk
8e9Fdet+7a3wlM6UNP0P/bNwxO3BBkOZKA2moteiNtJG2Cwa2v+6mLDVPXQEpxB43VNlsrtJKkBs
rzZCd9HyqHfkrFMtmiqmYYkWmZchhe2t+FrrDfhGXGBs0FojZKmmC5E9Y30vuFIOALsGPXKFEgNY
X4t5wfL1jAi7dxjWUrrh6pCPvTO2kQwdw8S5U7M9pAOnu6cHpa7AXd6I/TJFfr3RzNRjnp+KuPKV
/Mm+RBuapPu8j+DEleYchLI0hNRVQoUjuMzHRdk9e/JXhX91FSAD5PPNnbBWPKzLO/xp4rxizagS
OeDf4m5QJ+KSv2A+1x0/epH3XXJT+VdE+VXNXK3gYU9thCgyMe5LWn5tP8ysbg+0wPB+3uypfTtd
4tHCtViOfRFvSp+EJHSolO6HBoBeAObeVVQ55U3SLYcBfPw4I916MG8lpIx8WOUyYZ5YYLjncg4e
fUQsSgAUyyxk95SmAZZAUzT7FKWCyTMxOVBYcCJcFEBPt/yKVGr+xX0UuEOky+32fsxCx8brdbYG
cOizG1nbkr77pUYovTIOq7/r9boLA4tcS4Hbz0VDw8kU/R13dWVBKjvJ9jw71DUzl6dt3zSkTI45
qx0+aiNk5Dy1DY4xO5qAA3qR3oqymkg8A2nxf6XHYK18ftsuDCuHqP+w4uU/49qkFcC+qcuhcgVd
79pvx9NQjIX+mXvboNCBA2lRgFhuo5cAXduu9Puz0MN5VcJNUP98SKwncjVySUigDYHbYw4/3Mzq
mcWC6mwOeOJTsBGsbktmrm06Q4fW6Zx9y7Y6HN6cs/IIRG/k8sRDPsQpw/hiWoyqEu91QOtdEE4G
ZbemlM3rn98vpidWHKrBzN7Zsv3JatsbqX/DIkFQ3Zrbo+WiHLf69XVO59hztcryATwUcHlG74Pe
04z78JE8Fc6lumCPi92dfBUI2lTyKXz5Et6LXHvUOeE9CFq+wxQInwxGinGBehoJ/iPG2mE6fcvQ
yGYPiU5AL5nuPN15OHxVJOI/KV1q58UP1HtuhLirFNtvDEx4oi4dtViwZE7T1HnaSBpOEQMJHL6r
N7LBoip8UA4sKu/XjoacbPGvMPhEvwNbIlvtf6gmD6F53l74JPs7IApq/JIwYBTVrwXRcl9SNEAP
M8qbv5jkhmuZ/BKcVMKEa+4BoY8aF7976gHBI1a4b1LSVGHxR+J1WrFqA0uc+CJVw1kpXCTfQJuw
+U703WNjiBI7SWUt3o96fdQLUnxzBmdE3OmItHB/WofsSFTRTK/ag8+mxKMo5XMI7uPcEGw9Wvx4
lFCh9OtiEYt1SbnVDKAosvPvHf1WiTy0hT2+sK5evzNmjyl1CKrtgs4Zfy0s+v9/ny1bMPvtDAhE
Lu31oHre3WKTA51pfhlPD5yijhPF+9WnaEu5MT5WkMasDDsccxBuYTmRUM3Yh6XLk4s6l1lQjoNc
Awv0NGQKHNZckInZw49p96q+vug6DEmVL1RMLyLH76rNp75B6BWKWxLK4/PIukiAuY0htDmJrKCt
Xtf2HJB6bUmQ+DH8RT2AAqNDgqHBSaNA4XZ0bnvPP9iTbyVX780adxgsntv0JZ0uNmOMnOadbMUZ
piVfZ0/wrTpD7Clh8oAAxPk8or3v7jiQzR0KKx4Eb16grNlSK3U/lqRcdw+xK0kT6eiyvVYzgc+P
l4OoG91aHGr3VpTXvJyOcDDj7R7WsBJL3AkmskKDSde+YN+BWFJ8ZKj4KzVdf0pMoss6Hk4Fdxyq
2XHTjVvtnoimj64JCCmfZd5wPBZdKCIjUDqR8e9Bjedqvx2DLLs+SI21wx/RopSpcZ8mBiwuxQx1
0uuN3ijveYO7saebV1Xhme11BeEh6FbtjPhlz5lY53TH84lwW+RTa2ogR8JAWz/Z7NSFrAkjvBVN
9usN4cw6RIthddpdkeoJrOszwtDdj6hDYlvivELkRNcXnE5H+5epmWnPKYsC5Onn9Bx7Q7NCfVrh
ANwrgyxF3aOjw4fabv0K6s0GOEWAzZ6SmxZz7W2tLbZL/4G81lNqd3Lya1Q/EJFcqm2tP9hQFwx4
H5gFU73a8G7ux/CIRpICgwJLUooyB1g6CH75Wv6VRqNE5pIvLxYYnTwIaljsN00m/9CFTrZwio/q
CCH4ewT/XNbbA+FM9z/XzswCryYGFIOLkNS1pt0TteLepiyKl0SKtdBuLCbGWZM4aIhPsG8fcrWg
wkc3A8gYoXAMo11HX7xg30r+qf6udw7p1o9uiSPSJenOfvSFqWSk0A2M6p0TF2iXg1/tkpRoLyzS
LuX9OHVmutCcixN7iaFHhW14DnAIfUoMTlZsL42gZLpQ3qpkzFPJdAa+94UefVY6q4rOgdKhNlza
psWXVFiyIBCmKnNes4YNCuv7LU4/T1ID3TH52TLVLK3QyCOyzDzDFpDJNbyitMLbsrmGqKRM4pjq
wtCY7EGKxNIByA7NW3HNJIlWSGSkDhMVsD1Yfq3KrXH6/ACsOuPKcSEY9z72OOsIQxFepf8cPnc+
HyXfNBwxBq7VpEWgyB8g6sUIMz/ZJ6ZA6A56x7cbQlcu8hYNhIw5O6h4r7JfZqoP2zOqs2J1IE8G
mTXj4L57oG8s8j8Dsp8cTwbMLdSenNLCPOg1+69e8eDVj9tlRtr6rdmeKqTJ/9iXS0EYAGAwAQ1L
JqU3vtWvORjboR/Nxx8MWsF2SJYETG19ps3PqN1gOwPpxJf6kNUz3Znhve0Y1OuzyTmqSmJ9q+Rc
eFdNLJ4zp5N2Tfr4Q8HN/fMF/f36UnSuy06NwO0DsLco7fOpbN16MYcYdYAJA4wUhynbCtcio9Nm
qKCdXtekaO9YTFRQebsuZ0yAcLsmJOdqmp9pEORFyaCWlMISsV1sorgTv0qzAnxpgHd6YfYCrIGI
rQrle98MupKDiNS42SCksbRVPHp1Dr7ikWuw3hvps0BkGlGUzTY74cADeXow4ngDsQIRcYwr4aae
8RI8ATOl1wurhTA+gNIGJwms9uYswkyNN6E/aeMTVcN+FZkAq1tRD6EP5zdopFObfpMMzKZR8Fh+
aBdqP9oijLVjMLcqhO4if2RL/YH1uUNSipRzU6nIdJJmhTDKbuq0ujbGl9nxQWP6sX5KrlPmZUkV
f10RPxA6bODzie+Jj6SbnXTDXP7UgIXhQvkxlC5IAK8wO3pCZqX/2quRRs3wvZziHoxwmqF0DS9L
I5OvoSZUL4sf4RUcaNgWRLuUi7AEEtulKBSYVVpzj0na3idpTuutkEtb58Cvp0IMKEQOE5QqA9hu
UPGkAVCSfkTkAbdB4m+MzCvyk3dhbT6/aEB9q4D7kjZgJRtqV+W18YbseIGLjxeBpNniy6SkArkG
yV5AJkRxIla4gUFe7pX21nsV2tcWubFIG7cp/sunz4LyDhk+VEA3SlWTBlXaSfvFI7yOUtHdFpyk
DKR5C9/VKdzIY4Rtq5HywTo0J31kaFPoaVbTs7D1KT7vqAeepH1wipFGnbP3YGcKgE/KmwaC9tbQ
n+jjct/ZJjn/YQ9oDMelEjzHJw47yf6VGD9k7FehGUEXdNcWcdbx/FCG+Qq7/d0rrovISSpPtURP
2cIh2d4/3paW8o3F4XzK6x+W2ONr3KuXsBYVcosgylBWJXliwo2RJe96+qZsx7pFrfaEn4MPNC3T
+a477KYgeTZ4RigQHxnXx/P5M5zHiXwT5y5T7Dyo3FT8ylmfYn9TT96LRMykXpmBxqq0yjT0uHxS
SP3bqE4Iywe7zuFVKPNm0433tG9ZkqwNB+gBWGVnLwry7SFRQWxKjicvN23LakVGfik/5X7yF1ZQ
7qFG31nbxx26EzRI+rDca+ovH7PzYpPvmFffCval6nkV1cPxLFIbR+nILAwcSQeZXxisiP5z/4E9
mEuABsrEg/zVd07tzkmD9GCNlLpNNzsBZXKJAqiUahuD9RDsWTvOnafXfqEgobLwe4gNKGZ+XjFa
CBGN43r9gNUDUxP11ygypY3CTM2flNh5NIKhUQA3JHgDy1PTPJnKI9XvdFgZSi9cIv61OU/EUngy
YewfvqmcWiI6LWFX1esKCYkuLLYoVg9Jza8pqmcVVIKlUJ1fY1X2f7IxSVErCLzFKHbUDSDZAnPP
0o646Re5F5UAFxYK4LAVzuPhD7lUrTPpX/NueOQq2/hUItg9qZxyWnNzaF8DHfgVsR3wxrAIlGBw
TRS82T1wJtnn03+OTamv9B8crZNtKINehg9kzzo6v6ZwJLCKDTqWXKc63Ye4lpPhTTG5nw9VThfs
uXLxxiMJYsZ7jZd1UpfJUvVg46gyMZX4N2RQ2kT2mlJU7ga7oSaFLZRI4nZ3TSIXIZlRzp9fYAxC
emSOn3olywQYFtLwN6DZy3Wux1G6MkNpz+TmYWhnW1dLpu1ksPAqLm2dRokcvpIlqPChvDf/PgHt
QD2imUcsjqVFm4kQ0B+BCQDRelatdtESBpEDO3OFvzexU6yeiqdELC3ap7w4EGZe1UGovZbgeqJk
WONZL9GX5JnMF6+f4PWviLLNPStgsVklpii1nZr6fUBCzfGEbrZi8UX9E3wJ/r+l2t913GNxQtGq
WfM68fNbV4fKeCC9wEipYmst1xj0yZkcKsW6qQh3Lmv5/is79jJIIfSblRic2nh7ERl7BoQwOdIk
B8H7xhJ8vMavbk3tkIwawCe8iaxmWHZznLZw5Ih4IIuEqpPd1WV7yjkEeCLgKrpV4V0v5v3jY84m
6yakQdMRm4b9GfGnTsKLYmWvCcbXSzXdl+cxTwCDRU9nXwIh4VnqVRAvQ5s9OuLso9vyn9NY+hFf
KNHSLJOI/oSlHPjcVcTI76K/LnjFfArY42x9T+uIYiiGVrL8af7KL1tn8NgM65mLhtGeiG9xegv/
RgMdLZic180qJzjYQo6CcTnhwCTuE42JU8Jti0nRJ1C6bjipnJZcNv4NLL0f9v7UIwBRv3bEkjE7
vSsSIR/YzoYihqX7TkVxFWIYU9mCl1yERwB42nBijM1V7yBfVlsCNRLadrFJnDUOOHjplrxhViO9
zX/OtS5Fk+qKhWqz6QJ6NaBufpETcRVlxIPPKAvlxLPthb6BK3zZtc8Iu+gGjNNuEH6zHxNCmJaq
DM2XZGhQKMR1DtiRkhnel7T4CqpZxDJyb8bwSGbT8W6vZ/ErsOkt6h/guTi0yNcUuZPQ+A58nq2l
/0fmZ111EulSlaPZOLT9z1LYejveodza2oJBkfFcF4PBJWd5h7ZLu3rtCiJGRN16SrVxYXq1iMuU
1qmj8pLyqHEr/A061rD7MHel2OOQZt50BCiNgqGxOBRg9s8l0MshwRUPBSAxJQu7rEMmQKG8YK6M
taM120r3IkOwO8SHk8YtphM22do9TfwDNRNdqYbNehZWU3QdkPjgaxn253d1NktuvmWIIb2dPHdq
DX1MwIDbyL9bHunA75H1dVw0HgwkLLhFGdg52um3xJrJ4ivOWGYbx98/v4yffzjwJ54WwR0FJx55
Uu/KuVqlkOmaz+2lrwIEs5AVq1KU/rihdo+8BxO7UzVY98eAkdWoiDOqy6rAiHWEkp2XWBPuwtH+
H6+zQ/nPU7ePdPyIKucsfNsQAs95n6e3obbc4Mdskqn8XNc7A0rFKIqlx1B+uN9HBl3as1dVw83b
oaeRmL050MbUFc9dx5cR+xDKaciLQEIFufbrXLsCfyDoWa7a3w05Ws1AxyZPPlNo/GhKi1GVqq+b
Fl4Bn/SzAAsEOICRpIn3srEKlziO62iQ+srHodBHySjKxYYZGOGSu4HTcsTIizPs1vu9YLfiXtI+
Wr92Vx3kroMficZlkZGSt6va9BIZ+Vo4e+QbDJzpK1EjxJLHXjD3WvJPGWNCLQexkyL5YVBu6FU4
cgxIUvPyinOvPMR4A3AWyBwYTPzqWxm6XBWlOeiA569WNTFmX17GqwkrdhuyJ2oIrdDPKuC87J5m
O8B79PmLqjuf8D+gRuEYwYhgprheL9aSpfajIKLE78+C4j9gGvCWZgPLru8lQATQHRS2y5/JcYZH
kvOAnRQg0AMTzq5YgVtjc8hji7BNB/UdNH+5/w3i3Esu9uE9bZG+GFUtHWUhV/aQ4Mt6x86Ro4th
L73E7oe5zBzhckl7jNER8Q2Mrzespmjmu3KxFUf6bRG/WAOquMZZVLaF5CtBKwKbk4TpGokt4nnU
nP+4UGZPHZ5+ogh4KG0em/fLON1/IiFUK+6G0M0rYX3fJHFFXrpxfxU8aomXWoroNAkXPQVOIfjo
gD2JFDJhKXrc80guB28ccX9OnTaHS9sm+UDx64NIW+9WQoUpdhUFM9D72Nd12EP0Uiqi5yezckrS
3RsSyoaMO1tsK+oIbwvV+OFluAbKOAiCndo4j9qWbMnooH74r8b1dGh+jaedahofoN8V+e7YDrI5
5/BbuY52Kex9p0YqPY1AxjRT4yOxUezuMYk8xbf/bjMGZRPhDNh5Kkfmd+iWrFpTx2FDG+4+N0xF
3d3lz8oRnGc0Vp5Q6FWeluiPrACN+PIykpPvTsHaeR0wcUMJgAHdBNyvokp0+Z1UjZvvBM1odeon
Qg4w5mY5ysuEB3VdCBNGGHycotNwOHR0wEcjjNzlj2sX2L4/P2cApczcVSpNKTXKEnLPrWiG7t0X
yc5BWi+GbxMqtZk3Zoi8llYrwzpgQaFgHu9jTkgPzLf6cy9cANslDj3VQgtZl0iqLhmRpTPBRDCt
Hpho8kmkzDbDby6dFCfu2SPnn2TpP0EOh7Rg69Mbs7CM6t3vN9kv6fmfIQQOj0j2M6tmFDad9QNQ
PsAGpjfUmG3Zc21uJ7a+jo+drwasD2G42IJKK4eTBKmp7v++YzxfwQuGGmddELPBAN8nTpyqqQxo
hIiSOuz9yYClInGqkBi3nokjL0GhLNzZ0xYVpjFfJ9yHBzcE9PYzk9RfNMTaqPQmAUjU+eTmhCk6
aJTCmuo+KRPPYtWgOs2ycqRjfbNRxCPW1yWDGFf64IAF3hFSvTDTGCc0cWL+s3r6B87UOGF7APG8
Q4kL6+FRG9kHrN8qMojw/+3E/ruLxTBindKKZN4Os0vqIIIMPjjK2fMO39TPuo2pdyErvjJB5cZj
lihDLna3SYSgvnxrTl3jRIwLO4c4vALUVO24fzxcFfECwl/1yaRimIgQZBomT6Ye9xQAPfqz5XUh
lgdGylXO8cPNvqn2asWzDdsl+Un/34N+HbFjAKz6V4RnbctzWeo3R3L2577QClYi6GKSNBgTm+GK
VKOHZu2OSVjBVbKxCxbRa3ycY24gYwRJJ/OcjkK6vX2cmeLzelRdJ+PEyWDYR0dyws2dTyxm1J7g
5qFUj+xZtb8Ul5TT+R4/Erp1AN8iovoTx/0VgaAqO2nZItXF318Onuam8d6zxk64ejrPzZEdP8SC
sw/8GuViMsVlGQpAG6L3YZos1HqWPs2pF9y4sBL6xe7P9O3+i9XIt5aMOXuF5gT4mjEBgRek2wpk
N+vaNOFDR7Z1lyd9JZ/sDh6dKMHzmCEE3/0yYjau46h7EikjGNT8tc3P7upHU5VpU4LEvraQbSL3
h/9aQpIhHr/uFIjndm7MKh6qhvouBMJR2lOsWHPDOkcPKWSvyDCxWgo0pUnErfKt8rEL65NA7der
nwF+sYZsGsh7GQbfZa+itRpeXe7bVLy+R90nPY4y+wY1F8LaDnpJmQdIiTnfmkXigeJ6Y/E0IBv9
Jh/bALGCSx+ugT0N7oZ545Qy1JXwjs+0qjuMHXLkbgwrhZa4/qKebN10qemVNOSUfa4T1+aEB/9A
2Y8Zt4/FWTWNNxKgIeTPriPG34vNrXhac9vPeT1tid6WEGUDr1uFgOht51KxqPdzEEsHCfU1bxwq
AGX8WxqM8u7+0dxMEfIcWaOpOeQXEp9F4HX9Yw9jYsTUfWz/8njn0ofPQgmbQpj0wM9VkZI79R1s
QbcCYWcWk6qNBa+gDNNKXXhnJrPVUTz5EMOQmNJwb4GMLJDTy15bQVnVKaSc42aN1Ogn4Oms2fTQ
aE6fgxmDToWnxddvHm0fJqQp2ZJyPGJSPGYpHfSTcpNDCMBTf5w/gp6hXJjeU+yt9/Nu5V86rNhF
ikMEmRrvwITg9R5fF90EjGGngMi0pFVbFaGFixiS1m7481SqqPSqwr6+pTHDskN5YfPcrdqiO4zs
uCWy3w7+C9M9/MesCQXyO2YijgWU8a68RBiaXyso7jSMf/Dxcr3UmS91tPrt6NndDYsO/abLaPik
MRB0XYD46OnQYL9D8KgC9Pr8tpT62iUo7j5QR0R8ySrsrzbq+lIh/lTpfkMaolqgwYIwcUICz4e7
Aw2OjUUyzKjQKvXYijQrhqS42hF9YsauHSElhlaDRn154JpELjIGl7RDOSc9WXxm3QC33MqiQSIA
d4HDrUCPp4lzrr858REc8yPhRWoL1YT9X5BPS7HcRv1TPDbfVbP5jPxygAdGpoCBg26EDqGsOtxw
YjM7k/qoTgWPD1CHMcJvafkMQpqhvuuNmQqzZm18YplKnHy3lXoWaUF8lnqBI1V8xVNFUUs2oRhe
F0X1RAIRasQdQ07gCh+v4YkMiKh4AhmD91v7ylXcfgkVsTiY2OjsxMIqJXqYM/YbDrtE800F+yJo
Q9PrZ4aVeqpGgvnTsTrSMjUk1Q6O3oGnPE1C4WdRiFCOq/TQzP97pmGNtkuNYyY4Dz5rYDPHaGVg
1snkwZOfenAsYhO9TNBS6q2T5kVng0ILohR1+5aC0UJgssHJSqyuIJWqdK7oJDYlvJPbX2reLJhc
2Xs2yumj+RPMW5et50ZDYuSGw+UywGHv2wLepq8rdo75qsAg96LBbthE84NUM/pst9Kxdd0Ct+bw
l4mwGdvyADhZ8gMOnAqWKDYMZtJB0+uL39MZuF4lJQJj5mMXjE0g5f/0Q6YFzjBqPHNPll1/nH0Q
SRZE5ka900ZMpiudFITUY3lgBjK6WdVwKTC3wJt0qDj3d0/UQwoGKH/z18uCt7GQ1M4ibG90arfJ
sPrbAi+FH9lY6xZsmRvD+Z4mhtDViiQYcSymDmGw104idhEEER4u7ZdxBr0ibpjvhCPAwN1wu9LN
kOE4QQ3K9PD2Ekye6d2ZED+KlnTXndqNJkXnUUaHIjQzFrjG31uZ9UsJN0DQOJolOqSHcKFIvV//
LTegtKzexQgArU0NrRsUwn7lwipALAFXv47e21nBZP46hXp1LQ1zznqhm4+9g0KxhnhvFAwn3Wxn
H17o14wfBE1Y+pFViRkUkhEuGHFu1gVyAH0x0FCAZahQApCHY9/kUSho564latem7hLH/n79OKkU
v9V2HYWscxSXGpZwCZ8BHKCawqruW3RJVBrWzVfSLesxwuM2I/Jbtdmc2vsAeZX4vtAnticIMTUK
SjQXWGmLmAdYfMVPk+DLgzlkpDAUZYatwEo/iJccmZmlYLhxIf9E8Kt65DCMUhJHRpLNU9gDHNC+
11vRe2Ibalr3nxvTe07jtdKbTfelV44MNFzW2wk8EfNyi5k1OktCJchBYe/u/o1BVF0jmGiJHm3V
OVjyQo9gGPuQGeUW0Q0M+iNGkd8H3dPEGxKsFRDmtodGhR0JGRaljj1HLXlEKOrPXZJTrSUCQlvB
j9HgQ1AhrusPHzOXSO7x/EovXYGF37gIXCDUd+aVlErNdw6/R3G2RNHa3dYiUVSLYgKPX8UApog8
Fu0EDWLVhQ5XOgtsxmsqJ3k96eEUmbiLG91NXfvdfoDUJVa4tu008FDokCuvm/js6wJDLGExL+V6
PgfRm0QLftXqovu6YbAQJlafTPuE3zV8W63NhdE2TGzUeS/vX138h2V99rvO+p0v0B5pCA+jFIbe
XQ+BAzCEncLbPLbS5hNEeOcp3uijW8hBqCZQy8RnUWXj+mb9togc2PEh3Bo0FqABHcP21hkSbUu0
KI7RNZvMLzX1JxDo9paFkBb3YBSnpbTeiUluMyeqoHG8qRB2kWzqm3EBAb8Pyez5aMAYZEcOJ7+M
5aODR/iPSvswZ6npAJvhUllOFNK/4xSuoAbH3vt5J74Na+2k2zXOHr+fLEOzK+ICraJwftL57rVC
lQSHYNgwUMtVd3oH1E8HyL4JNODaxNuaO+pGNnzuIhBFA7OHEThwJcawFD79Kux3PWMXSEN3g1uU
SasbnPpheO4tJziNEcRLXYFgv63V3UF/y3FttJ3umCnixXDvHKTvROWkwoRCvrtpoC1uSSNyO1P7
X0GoyuEBix0QRJqGGtNDHE+FNF4kjOE3YoykJNZEcF0gNZMuPkeyua9rfmTBiiEAcYb6LSe9asBI
0rWHIB0LUeOufHsCwFGX8jBHmAvDX4ZVQB9jrEj/WF1wFdR6TQt2ZTAYfN6H6GSJJppuBVQALDEJ
7s+tfkAnrjb9w51MzlR2J3z6qLv8otp5twzeDBbJhrF9KBnbgYHVlBc/A9vj4d5kd1DnZfb7jJOr
oV1nSkEJeoJB+f7w7vGaHkowWmqC0FQHj8cIoY367NHx4EjhNkanb1GKoU5b3dNgX5pL+JfkIvls
p8DDROYBf1yDWYrVKHPsthKcnPc9uCDK4IobMBXP/1p346UP6XXVBP0VOe+ioc3B/M0OHt/62ZDY
EOrsqhLEuPCuOBm5aqlEQwyYAyW0mHitJdaoAVKlIXnFHgR/7ZHH2LKV44UbIBkhLUWb/tTCBnzA
+y/NzKACghRW+0oC+bxPl6mYZjg0mdj7flPPZT8MbzeQot/gocm454AFIcNkrDKU01jdj1Ho571D
sujbkV3xyuKvisavwSLANaVxOoPHcU8PZelIsLtkWkN447FuGxJCasWN8rahwTxpqRjlLYLbX2H9
EQ55mxYJvYpQPiVqfyreYwzSyOjuCZoYt6DtkqCeyql1E89zNmApQuqhSGYApZoGvmlh0QKdc8Yj
wZultKlyvQUchzzPvspkFr5PIWu1w2T+Z3CDxNQWbVHOKTV85u6hcNQk0bXPGKPEyPYRfKChTg7E
tklDW+SpaompBztihdnapkP5QpPnIG69ek6MOpEIV50G5LtlvDWBxN+mQYhfslG6NVezbqh3czoL
cVfIT7YznusZscM8bdhSSEbDCnuEPzviR3KucGzvxsavEC6LXxGhOM7H4YNEygEE8PLCXRqM8rOc
Spyt8nuFwQQtiWBPzlK9x3b4CnUFocoaRsbWtA2ovJMMPIwUm14aS2g9qcK635ojtn+8dHMlNELv
TmWAj0F7mQBd2CdG/la+xUhRGSRp2Q7DLAceeAlAa75XUYqsSlku0KI3vLhcXvUoQ/an5aRPIpqb
OYPZbHHY/trzdhRSLX34mT0B2vnstGdE1YIxL/SKxeVTvtGdxPJMshLo9Cm7FrLXw9qzx/x6M+vq
DwnE1L2NOYZQOBL1uJ7xiAoScaMNYhG/tNXpfPfWR8uNHRzZ5KkRw3RRncBKNJS9GmyC7XweyJ36
uQrQuK0vgeY44Rz5SbrpMeNyRywhlSvkzZM+hUknGmh+z5L+pbXrU0j0RFVTnfWatIyDrm8tfhqu
CIuiWmfT9c4voUxSrCJ8JKWh4rtae7NFpgaSdxbdVL45zB7fvb20yQqbJzYvlk2LjeD2mnW5TN0z
BR1M/ltJiZM7QQ6unO2wYA6qjTnOUl21KAViW6KXQLewDES6txsU130RCzYOHSb8tQHOvBC/da+o
hR8y/A86N5ncIyzIlMaV9/Bq/7F5R0pvBG8eDWRM8mqJ360Tp/GpBrekExg/GYlgGqhe66QgSjVB
upZWJtNCsst4s3TywmtC9SeAWE5RGuWfuCe+jt2joMWVAcfz7vjXlmLfyiOZivQlG4RpYLlpaI+E
oCczseUgjGCX1RVj7mpkbm6ZOGCSSWtoocG92zlSm+P70LkD+R70EDkbspeTOX8sB1TJwM1QeLI7
JR5N/ws4l3cdVQGHYYiPPBHwcutPS3IMfCQc4OuGe9y25UQr124AlnsyNCFmgdB1TXPQ6bzezFzo
caaCEW47m9MvXACzFFYpNOQ6OPDMZr9vRXRwls3ShD4wKSY07VhduwZ58dhey0MnTa8sujymCIpl
1bPVTA49JZAnOJB5bQzYHahId7fkXVIYShKhb4RAEDKPZIJFLucEd8ieCLxjpRUQSwlNJS+Yjou2
fQd0SUgnfxHU6gg30ccJIo53KknRDcNSgqv2z5r4MFiDzw6QVkE6CXQ1cIhVEVnXXgEstYD8IoEW
mToVkLicVhHHd5txmpjrk8BdUcb2r4bQZpjDPtncxwwHmLxCOug/In8pPuoVIuwUOJAj+okGpg4s
MuDyQLkvoiEwwFzfPY3SHJlK+/ocvpdw0Z8DgoPsPCBM8yOg1ZQwEQWvaEgO4Sl3/A6BrrwUpspR
rmkJZqCg1Z0dFVUkFzSkRD/FN9VAqzCaQsk0qQGq6ByPVa3egRwBemD3p6knTjj1tuXNn2bzdS5F
u4XxOxU2jZXdIQC0iZl0qhHPA+DVQ0D/BZOlddXTaBl/vUCM7bD/u+d+H1F6xzVAKWUwiR1xcdnJ
GPoZeLD1RRLZQc5CCVaKUNfkeX3p/sCzErmtIhvvfjTICTnqGESkOIO7lqhh4kSLGXzs34Cw0708
KEfYWm6xOP7lBlCmLdjoSpPmTBrX+8affBCg9J0W0egfk2p+HXcAWrZmhkQCzjcg+OcRsoWOApoX
FJTeiCUXT3PNVQ4njNCEnuUYXtZAmLoujHmD2ZrnJrASdtAweOophkGFnEyDMljLT+X7S2jFyDE6
r3JBWHkg1hEBdzfAqJEX3iy0rbbKbE6wNsk4wFreCuTtAehwYsRy3clkRkMk5yCmKEPUV91InDzZ
pn4f79Y5hWvF19p+kJ9HD0br6KB7zwbDHZlFOS+dMKBZFh03MPjC2ystB7v1+2D0uDBeSY83u8OQ
nNWInIi+gkfwaihMSFIuMRz65XM4h7rv+P9LILnWlEQ3ZzyavhA32iC13Y25uLHrQLKrwakjpXW0
Z92olA8sYqZ+qF/eronmn/O3tS0hQ9AD3715xTEqlaDOkazPZlvXS4edwV6MZV/dM4LK5s8CTkmk
v8M6SKMUCfpEuwPY9p+SST7AWhbqdUWyRi6t7yrcGqP8PMJv5/bX4iCDlA7NEwhpE8FDl9p4JpiF
tgP75cOxiYNR3COPtV93jegQkf5XuYgLKpe8mJQZ2LBZ0zAdJZLpBvK/9lQJ7Da5nNlkwfBYLnil
WKyQNQOT+tFlmQr7yc5r/6S8omegAQXKFM9N4OnVtavQJLYme4g8KApn5xZGMq8nBw7/X+aGJi1Q
o876V2D3EEbZ5TCPWXrq1GoVfVV7HdR3Yc68QHpdGpwV2IgCLGl5Uvt+MxC7Y7RgKbSpDRrw8koC
04W+ud8OYn7vpqhqVEOplC5PcWsuK72/mbt1eyhdEvoO4NtojfaMnI4ABqca+XnI2lqUtUEFJiZz
UKBNycpZu4oKem0RJkUGKHgV0L30YuVdCll/XmJWYO7lNoFbMcEUiCHz4wYAURHp74ozF7LG8DvE
MdKHnZ460Id2HZsDqzBvpV7VM0Fc1/JyAg37SBuZM7EJ+SMZR3Gbf6s3XXL2occr8bdBFpsZdDrx
Ti07PWxeTjKy4NNYx2aASwLzj8/QMaZksY3uU4BlDr7x5XRjiUQcxNIWmGWWLtvERby6oQ1tyI0v
E/NDB/Pdpqowkwp3v3elC+5rROy6xOPQvljhi8sNiR9ga1PyGcRb6h0tjjdssq7WD++8Sd3gKlYt
LVklXiqfwrDzUsmCpiFjlVwenKoJP3G+2tRSrgXGkApYu7k8aLJ9/grzUwxLBlS8/HZ9TJrtF5Xw
mq7roITRC7WnTMKM+Sl/3OaGWC2xT7luehvF29YEGQ5LUZSdUIDtss64z6YZigA6bQOqLPjh5mL4
6D4GFvccv6vl6Tc0CtPD05PvSsGhFCxBIcNoS36GImW+ZKe3kgXayjxiDxZ11XQXhRIOwSfCXhB5
G8xrcHUYepYUjmVt+u1PuypFYPzCocFPyIUcEzVL4uO1KL7pz1euIonvfJHfsbycPtAZjQ9n5wuw
ZVPhg+SoZqQ4Uj1nEsRch0dkjdYxfh1jmWqYNFu5JDXdvsI9OHMkGJytw3dCNqzMYiM5f+OcEfXg
7TiFzyMjO6oK+2a77L2A/ZDw61hHEno9Znk3L6ti9Vvstenvvz8J2lf2H6hOt+MXuea3z0AcKDsw
06v0OB9fg2Qlc1xB9hEHj/zslu76gzuG47ND/ZVdSe2Dh+rjnu6MuF6r8ccSbSDhjCMR09J5R25T
6eYnYeYgFQDWZK/tKSNojq7xM2JXoauD7Nj7NHKuMa37dgfRbjoDw8gz1pSRZ4v6C5s3ShjYZayn
gxAbSBwgE5e3ZI5/dP5fuQic1x/yAQc+XknPSHV/UlZD0sWYvH2Dc/doGUyJPngTpan+bdBm5SHN
rkxQoNE1lXiiPJU0eVJieNm7PRgjEAG3Kw2O7/PNBXCcUxxESugXeUomuNa3nPb5yQUOaZD3cWNK
OKWEOiJmHxqvBWfH8KFxog61h2pxEsKhfwCQux1L/z+t/Piotm5fIsRBw/Vt/Q5HcGJAI74aPLqx
muiDIu0SG6X8KI6agYuSz12HTi/81ixJQEqxaCNO8wSstBxjGDOVFH+BKivnCj6tLrlKbnpoRLlm
jpciRTkOAP3KBKoFFkdPLpNV0t9HYoQTm4cxILKqbnhsNt9kxtSH9XQFNTo1ZXiwwK2EUaycMfWI
2SoVcbPAY0T246OhvlANf9q/kOspViY1Gq6KEWFcQ5KeExF6CbUrnfep07MEp+oBZuvXb5OGv1SC
vr/IOPKNSD9UHZRNmjRbzE/cPUXUozBLPo+DhuYdAzNR3t/WiEZLNnrBlZZP6BhavXuuec8Vvn2S
kK6o+/5juVwhi5KIwti6319wRIbk9Lzd+2Ay7c8s1fPxNvYIzB+/xcLdbBSWSxy21QXPu7iOLQaf
xlJF9FesfPmTqkXTVTdyEmmnKTf+NOWwpvE6qzfzJfq3P5YV8eE1Z1JE8oq864u+FHI6B3I8Oqoq
yeN/oT2Bo5F+2YigP9YYE2h2xBnJoP6lw0rxDlyCGUzLH2ttkleGVD013WsTXa5nYprjl+HanuJq
4KzjPoYCd6fl+6W/faSO17bDIuPa5sGbi7hP8lmPINT+WOs/UVPLmyC1PkeqHS16qi67kIDoDds7
L0u1q3SMDC74oZBf4yqBHs0DtKl2tbB/uuyEqybItOGUoXSqlAklZczgJ9o9l5vfUuOl2WHyB5PG
lV5YEGuSj8xhiCkjmvpH5DYwE5xh/h2JTldsrr2OgMRALNpbtfJC9i0Jrjye41hLY7w7wTSzzzZa
YE8mpiY/KRZ17+zAPbkd0kG/cP9t02oHPMFZBonag5RRWvpaTutKsBmSI4R1fYK3gDNQH7cWGxdd
DDZUWB8nVNEblzlJ1Iu2mhJ72kfGRptcWvRnaiaGKpsKO2c5tNtTz/dFE229WzRrTsy24kFInT4b
Zv//9DlTJIAhP8l9qPwoGCWt62XagvagYV/bwa4B7GlGgw7rNTtWey6ETwv4HT4PLIFirjgkplgD
Kj0Bpc5xyQtF3nZxhiPM2/gz+QzKOgJpyBxRTzpG5B1QdsbQlSjq+IHExe8Lptu7ZULP02KnwuH2
NeB5TeWXzNzItSe5HhwmyU8pyFQZEJtNxWyQDqlMRXyZLo3XF15jQ0eNJQtP+DuqVd2b43n/4VsW
2Y9v/WnE5yLKzsRU9ngBfDxB5YhL66MKHmH56gHM6t2d4jsyDGMUjXDXj/PKweshuyWwXvyfvNz6
SXLF9ffdD+WSNT4sI6/Cf1XFOUlgEsThB3gOvGzVRzYOdFN7GLs1h85B3YmQefSUzg91y6evIH4Y
Wm3eW6ODKsj+kUzIYLCIGJrDiwEd2e6dr1U/rYlrHDxmAW6P7buSY4cSfmY4G4XBuHkj/+1atG6N
7P/y6pZAKklybN9gwr514U9dFYzd5//8tBRzEznbaarYz3A85qrT3bx1wB5CVSDL6kPuq954fKcZ
j5R8JCsNMsOvcU4SPWWaIX4pNm36xACuz+Fuc0QZBQlgPHFpRxvGgeT/e31bzJRMJLCiQ8fkJq32
Brn1J/k8DtMOBMEvThFBFmkd+863tdIMiTwuG3Yyw1tsJcacZWE1/WojEoMj5IdOz7lgAwzt9zME
RnV2000MIQ8CH1aFb1AEgZkY6rb8VZSycWf8/+Vz65d2xMtlr3rgmUmttwZsg3S7aa3eQ/hN4Udz
WwdygrCQIFYEfI3TSVo4rNVfa4RRSTMdBjuDX5F5ZZYmg5seNvXQuUPmoct5a0fQUjD5NxU+gxhr
Fr97R6c4aUhFnNEOdiAIvdkIGy1/oBPmVHxh4dzy1522bdMQz0ASg9iFkC5oAPRF+TobrPsXFiHp
RqK2DInG8eCLfUti/0K22NeRdk92/wN1ZOebwMQBIgLHpPI1/Z2viFSXqrOoh3JmQ2UTp3U+2hI6
mSfSVV738DuyumC0m2g4MzCv38QsSvxhETJMdBfhd5/eW7aHRAs28jUk5c5Z21ImS8iKD5N3Dv7A
p6F2I9WsYjmP/D3jjUf43o6vnhQHwYMJwb0nh6+/fVJlNOrM/bpvPJ6krZDqkHEPLkA31dldrmVL
bibh3p2deZzKQTM61dKRNP5bGtJQv94PIFWBV0CNrASPr42mmYIDb7zD98QtFD78YzvoqmclBDfK
0tqDmYLCkmeTLZJyCx1rAD2ePTDE2NXdHeIVbZUlKSIctBRq8iPZHonL73wyx+4URWuD82UNxSKc
dYTYreuBYdj9zW91SiJIe6t4juyYtHbkAdxiW8NJZRoB0WSu8nSYAftEzyud8lCg6dKJFNaKTvmz
nYL3I5M4zYFXp5+D4tFVXY1wo6nxHe2t5C2vwUZI/l7XXz9pJB6lq9zLbfBHl98TxZpDBUL/TgHV
yvaPFZmVcHMg8r7Ot/0xQl+5YJxDAPPXM0uNCX+1qj22vreP18Th0VRD8FnBGQEfqr23xBrM/R0J
bjizpIAs+e6rtQKcyOv4rnjPuOKdgZn2TCawcIlf/Ht7rQYtkBZ72jwEs/ivE+Zt/+7SXTeUNbMT
UKTys0892AW5L/2/2XjHVZ8wF2tCjnCwT9/PZH0MdScMNc2oSh48ocPfJ09Y5rPGy/ssgxJXt2/C
9v8cDPbL0AmQSSsHCeRrK+64Wq9XvWbI+aVLQb5gNQPG3qDFWv41Ks8pyGfY7hpeVjOmWL22j2+Y
AT3vk6i9hZIvE4NWq9R4pKhFGCc68TcWtrpvGC3eqkia3Q3Dj5DVTsvMbi+qGZRxCMxOzFJLqwaz
PoC2MR/yXL4DVqlKkPj1TIuhhshqM78ao5+ACU2IdiAuUFCNM6NZ0OAjdT637AmlZfk/agr0KSO3
lRTNFZhIbXXMHWWJ5Jh/Yj9/4YaEUGggdGTPtHIAZ+j+SttMSEX1kEQIucA2s2J9k1d4upEjG0XW
dItjtMCYWgkghL/s2WplT1LnXheqXKNfqY1MEB1xI4bove1LVUG5Lm23bgLS9VtM5TQNePZ6to5u
g0fTsbf+ItGiAcx4LBue9tWanIbeTbeYExxROiGk5lk4MIUeSW0bOaDOLlqLW51wVSDOXDYUaA6K
M1P3DKoxwuFURXx3rd2KOBwRim+4lMzZUK9CMWndz1/AcItt1xb0rDR5IFR+4uFZJE12D0sgxJBw
PjHxzT4tOf+6YK4J/zI6bxAG9/nOskTh3os5tyiqyvmiR/Cmir2NpjAv50ZFWVk19lH/4gNvszgA
vbCT1vOudWW35qkcbElRJ91vmO+M/z21I1HFYBKNNHR+imEv2eCMZPESsYlX4uqL+FN+DEj2xuf4
8q2E+GT5KWH27Hut1hxDj6Fxmg9gVkN31Ruw8r0vszWmKKpl85GMn5oj8j7m6yzIMqLLKjbYN31Y
cWVJrO6Bp31I3nFtQ/N+29lElinxImkMg0jKA6463y0sxN4lP+nFuEWGTV+f6o4z82px2HkdgnFV
BRfrqcuJSzUY7DyhV8uC69TFBfIP9FUtELeBaYupjCu1qP432fuTFyqeo4HRssaF0XWwFl1sc58O
dIljW/mVFjmbilIQyBmRfdLKgBQNFHgt30vczLnze5/SfagfzdOOISUMMWxoaSwVpLWMV1kiRfyS
euwRPDjv2XvZ6anYaFv6N57fONCh6Xcb3nKpexHqCrFGa+sw19S+xfA/bu7xDCL1mrHPo8zetthY
kXDksjIiCIN1ylQMHXDMJer25Tmguq46Yxq0W8MyIjz31H+mjgDot+0RphmnebKg7KzgA3Neqkz4
04LDH9rzTh+I/7FEanJwA1F4A0jR9vcbLDjzGChYrBrPEf4IyroJPYurmN/XQFQH+mpLE+aDeiNZ
NbGQ496Khet+UDR6Ggw1RF2kOzPJtoGrY+3ZaMeF/NL6r5I2Bq/fhEiAsjCvvxRE3eAXlGYSlfJ1
Z0NlSe8N69sBKdcorzJffbA1xAeaMnNE3GDH5JtujGMk4yN7IcQiuEqFYEnipBwcWYoCAbe9jA/P
OWkwzEQUfoah1zzL6ji4rLJfUL+l7KQNvLJmQi+jE8P3wEt57pjCglLKDfa/qk48tt60LKUp0v8c
SG1AYSGUzkHoFTjPrjMIP0XvrD1wlSFpEjpugx8h8wcIXLHrvmHxGahroHqC/YH3DuvFZGkVbWPu
/FEsjqzwadec45Hu5KW+hVMxVrkHim93FzhOCqCHRvpqKvnfoIaYz5+lIUiZorNLnhwo2VlBzosF
NFUZJpieLRNLMuvxAviwfMHyifg411fvSa+msBSed1OMRgZFi14YAqBoKTekjaaWPIdgGXRlaLlD
8ohrv2WW45dLQp1dFFsJQaiAoIdgTaffmDFEScEdk7QzLiXu+CJt27xWRmwL1c++ZNnKhIp8X+hU
pwNbwUD9WVhm69UCB4RMqH16fPin2hQv+bqDrutcXTnQgPITFcDyPGyRQV9z3KFDjNH1IDOJn4Mo
oqerpAMn2F802t7+tgt6GCdUkQnSkvJxbY4Sa01+xpRmhllmMbfaJzAygmcyCYZcILgDIZHmmO41
ZC7A0+Yd3dFqwdR0PMUAJzvLXXIwPitxLXPlu4CtQWEoxUKUpcvynp6W466TqW1pqYofTQtJeh7V
PHWt7kCELkR/5B0OQ5tIHrrRlX8nvjeYZVJhh/XUyZ3VlBVg4iVqkGggKMbgGmQ6pHHTjsPjJS17
TiRuTDuVG6+Ex05r/KTvqs5BaVyJaxEHtRwwY9Dkw/xcblZi4u+YLglDHdXaOhTeOG9Ebx2QMEeT
2b+CSACzgLbxC1eyzuilYLszmLyTv6nL8SBumHsxbABEEcgnx+XmIBGvSgoI9q0YUjiTXz7eb41r
GoMnMdGrDqaS8KCi0oqsGl+mlKRLw1bGr7VA/tEx1tM0qt1Xropu/RnHNImb3D5ULCm3z+WQ0o0G
wXmOSODX/nwYA/k4sDdKZcdcCJXGGgt92i2c5PkwDkbgDe/BLxkw8Ps9iTQ73jeYlaPqL7QRCpkV
hX+QKS7bndcJsMqJDbTYl+xLMEyFYtMsCorHJoKFDpV+v9Y6ROFk0UWmjItdsCNl+Nb/iFzrWmFP
vEu2T1grnZHsXVgpXWanYNBm05aos57lW7CPKAoPzcdYn6X5ruaZ+inPM14S5bRgvW/2jpyAVIHV
RCx6szIqBd1f0LOQK+j3f6cucNdNxX20rvLvmjkMV94QYY35ycTWCNroRaCfbEFPFtUtwT0WMmKC
uRD1tUAD4HfAX9OlMwCOIYOOcN4sZ/u1xRCBO0Zc/zfXJ3CsQgi/+RSIsW1qky+eLHXOW4XE95r3
NdN8aFg6HrW1pXtiobv9JT/B2AxkmKqG1f5VDRtXWvdqdOge3NTrMT5CIuYLWKjsjXgknxmbtWJ3
fwmxFoLACsDS87SFuyZqTnjEVKR78FltidazVPGfscH52x0Tdm0kI5qxNPqGpAWo+vk9hlxCqpwj
MeamLYQ9uhIV9IjnLsJrKzEBwxCtF5HVZwZAQy+WqY5BbMm4YTbDvcDSclBZPtGa+9B9zvEtVwri
lDr+Gx+dFVU5r+iVXzT0SRSGm/DdbWql76w2tRE/Q97Xs5PpNpMSzhGtL+e+oFed6viSjmHYSIJa
XyCXxZIAM2z/J+3m1B9MjP79WgfjL9FXBdIOgC8s66vjNc14W2urMKxCC9mg83+EMFRf9dEx5ljP
Hb+m+OvEJ4SwMAW0hHtCF1oi5rhUoWrh0Av8NRCuAyKKjjex3ILVXCpJa0NLPNeuCeKU+KXL6LOR
ECcAvO7gNpmL8/ZYAVjzTt9CegmsEn67DrghChNNn1WgDyXCn0KiNcdRKkwCPgu/sF/HHldf9rFE
z7A319h5tMVRngu5Nclb/iR1vnnGKAu5RhPE2sUfvth4ODeN5rRQQNdZ5DX57XAEBQ8nzK42r8GU
EL8MqUOaBUMJteE+NuI/agxUzlHWDaST7k2Rg6Gq/TQAXcn2dJMbZ/9koCM2P2i/zNoG+Im7QHsP
WXR381S0eJDbRceYCWmUgL/TLVDJpjqT9gIONThBpnObj81ICA0yZnUNp50xI1rdin9Ir0NUD/DR
3rzEedBtvehW01fDyKBLKN93aXUmfJkosDRUs4f+BfmZeJZTsPbNx9JlOuRnCmQQXo/1iYFMU4fq
UjvYhg85yG5wpCw41X8aMLJQW32L2ahcXgpAsmZclsRgQR9XMQ7pyBPkcEZV7v0tymnKfCDdDJn0
0nX5cnJCywx27zbXeL9sNgBi166XrErtQTb+2++fEtFS2UumE/10op/X+Js2U0oAFespCD0UI3VM
WRfktuBl1mKHLoS7oAnPkTtliQz68DMNYYQTcwV4QNwqKb2nC0Qldb7a3KSZgiQvabFkVggH7xPK
GfHI9tqLpNCojOS3pNZN/Jv7z+FzPHo1q4jU0+I6lFOjgZzZNA8RUHxBtTBniMSINHVJUz612KHk
OOi62m8oLtauiEf/0HkEf6XDd9SQJ5gefeTnADQP0kFmOX0KPu61/vfkBHOF8zczhg1QPYzcBl1m
Xf8iXMuzcxhnNVBTHJVREMUJR1IlW8ie+BIzP2AiuiIMli2pCQVW0lZvwCym4iJCiDNQY56Eg+PQ
+mWPdJcqSPs/VBUQRklMm1AowEo/uOUsgO1iDtd6QIyagUqGaGK3GVCuXqbET06MG+Xbs+7Zn/bP
OH5lbNMlJYXxyESNe+QCmQ2ZHSlO7UgN34KifIbc+aBynvjYhWWGaCf5AF32ZDMqnoCBMOHb7a24
JlQKaNYCJMuCl6eXXLlsUg5UpfxwbybvxjFsoh7Fod08nm5WU6UP4ifkUXSPRxAAY1Yq+W1SLTjL
x2XwbJ8vsrlf9UpVm8JKhuAVMnWDcRT0XE52jhT2wa09Z1HF+spDLZszSg/AImLvZf7yV1Glr9RJ
7MqJI/dLfOnJbuXlwnuCS29TKOmTSNCj+rEsg6NBGc8NkMIY/7863wPbum+OhlPVLShVQOgyO4yh
hepP1plnJv62yQE5vzVDzYhTbM8WP6vM7ZBi71SJoMTACtFsrkufrejqIW3/Luyg6pqGLjrOr2Cv
oJy4TAfDdTfKowpnqYjmdzlrj7Jn+/qR/b4Og4wXwxu8piVdfqXg9un3bDXu0qw0cKFBcZxPe2iL
bW3yLRQ2QRPu8kMTLQ6ptS9IcIAi5RZdQUdwn7+5Sl4+vAjpUXQ8mRT/NYmex3qyJUshmyN0e/s2
9tHGiOfhFtc0J3v6kLOs7X7IooU3UcED7zgoMYq3YP1d5MYRvuDjQF9y0J6rbkhHNE/KdalRWUvT
8t2SNW+eGlifANwakK2cTRSuA39BQBm7dvQMzRL99Pu6Qt8lLwr6M4MNQ9/SI9tyD6sEGJbmCv1m
RWhPEKmwjApFMBjt3aDPl/IjtkZZiDEvCr4kUfu+YsPXqt0w9P1BqI0oaaDo+s/nDofd7k4pRXYN
sK7R2q4IiWDLf8IuHA1bSvd1g7XzhP8oT9vj/KG9Knv1gEMwNEzh3XEJAdssKhuzY0r1oOks65/Q
ntXNvIRLbdDRMWdqMgZkePHcWT90vZVdVuLrUOiuSsFgdpLd1xepvg2gkNhbC4puYFuho7/1poyx
SsKFT9g9+cZQRgKwfMs/Mf6PZPs0G9d6TewLAEb88dNH2mP0qKda3cS+/U1WhJZD6rRbCroB0Nw2
FbUV26nFOg7gSGP2pwXkuNqEazP8DMxFWKYjQ25BRjJc8wOV7FXdZiT/2TNko75k5aP7A2ZD17fy
sfIA4NmnGG8fUJ0iBdGRlvgH95iT1M3cDQ0P0L+fzZ4c4BFbMO1G1DSHtdubZYEA1XFqnOEZtg5u
Ca5nNB6oxJ4snxXklg3CZUcyAjHE6aslv8t2SXfd5WVXz72gQWjq3W3yRRZh37GTBrAN6sDxOjwA
RIxk7t3B4KcHriPuHZ9U4M4iaaeYon7nDw1CffwWunLPx9QqeOVxKxEfP9ZQmZLThjgravF2b+er
ZKblzDKG3qLeTPwlCNzBsGPWdFtovA4CIqXyhRURGsyBmcF462XEIRaa+p9/L6UuICKq5y1IZ6Md
hUeZh54A6oNEDMro83lzbkjOXEfMh1gN34aOXoaKfolawfnMmNi0g0/VVjPmQYGCaKy+F49B9sDX
Gv90VILNRdKEz+qwM+Pegr3pCPB2j1aBIj6ofFuu8LLYB8pns3d68NAZ1MAJBgbNJTTDycwQ78Fo
6sgf17W3nWTI4cYGqafSFKmks2n+ksZaF2E68w2aPRuVR255BO0xe3z5/mH1fwcyrGV6VtUJcR13
razmrUUwaX+0IbQo1bsONlB0MWNwQHiOE0+IMkIe0wF0OrRUFjvNAEa6fS/7kre+wWCNYC2kYZ90
Herum/xEjQcJLA6vECQKxJBARceqOucY3dUw1aJ7be+ex+FADS0M5dCRyGLbmsFfncvAjQMrCBXN
RT2xT8+Z5OzRESTKJPg+Myo/pHAMOPnlGL19irrtmDshF0TzRXVePmesGJeetkdLrYT08TPr2g5a
UBU/S181G2YhiQWKt3CjZVOvRqOPTnynerWnsUXQFgg12Obp5f1SOEL8p5VeJZ9T/JiG8F/Dey/K
QpyVliqX9tgvu+hkVDj3JDg4J7BaA8gMxokrQz4qRFYzdVGCCeRmT3qI/GlbIFe/7EO6WQMqMPDp
3Qs0Wvk15nCMv5CTYoWkJR3vcmrG9fC/pw/SszQztxfpR4/3m7GXOIULeFTmdIl3hM3IAmRxz4Xc
HI1uTb70db+i9ak3K5CjeLz3UfVZ/g8f+h6eKmQSROoev6n4s58Q/YiDc6UYaggJ3Y4SknKrzFJ8
Joe1F7JpM+So3DvF3l1TTymAvfqHdCyDYmkHS0RZ7q2M27xqvWAy7g09hU0cmCanJlihLZcHloF/
/xrtuxYGUASchGIrvpHWpUjOPkhvFJZX9nhbNdmCsq2Jy9lx7cWC+La1nrxAipZfIYprah+ssIrd
t4r2Ta7CF1ZxDNrsgqZWJ9XUF/3Fl1EWJ0vPzX+53TQSZh7+3A+FeKfhGPO+oWBQ+hElLkrKnu+4
e+0RKpT4bZDgqYGXUp60azDuvgJI4lZ0iegUeD8HvGgpLvLzjWYkNUcNCB07ch/ZyOlMiGNydXhi
416Y73JVoJZAIRQkELY6K0WMCP/JwjoqKeLC7BacUJkaWbRlc2TzrXjm7CxlvgsYOZtHelnX/uHb
ASefGc5NdBd1N8YxhPYUcmSwW24yf579mu4AXTmZKa82rOS3AHFhT/xf61yMqcTxo3SRRyrMIJMV
fc7OegqKhASKu4c8Nwgc5R0mhfvI1DBO+mMCk5QB8iCauDjVnGhv376W0uVlOs4oCUj9xnF9kfT5
y9PeYkI8TooEI5Mzz24cOsMZ7vrQNmUTR1nFQPUVlx5DywTTH7oQRZDuaf1icWHWIcrxt7PeprVt
0iUTymKXfkUF5aYxkvUpnAC/b/C+dU6euLhiAK106zv6BDjQXarCNLU04rnwPqeANjxaBi2AAKdt
HO1vQ9baqmczXo85XTwVJPT7Vd3RfudirrRFvUsBeZM9GQIFYmiwJsZtnnnJ4DiFgdv3S4cec3aN
DnFpHvgvDiV1ixa/dSU5bUjPIcYssOhgdboslTXTkt5YMG3uZlT1NlktB/+25OWZ0rc3nd7UISkH
NBT1IAfufBEp6LlvxYxAvbJmThZETuQjVv4Z7ouxPVrS92U/UsyNr17p1L20Dbj/GBwVSr3gytMh
OQdT4CY8gkleMz5lWBZAUkz5ZU5z9dcwspTwl2p3Xi0jGZT/FYMEqq2cHutPP2clrpG2LWDp1jDG
OJeF9CjK8Cc7QHknxQnXuqvaA4Yh3LEyiMduN2Dtcy4tgN8UAZN0rtDeJGU3gp9VQ4Yvr0E34Pf1
p2JX6tMSs/9aAZVDNn+N1QpyjbcRW5a/5/Wxhxh0XKRx95fYHG2DtYKuNYUmQD9LhHxrN4UM6nh2
2oBNerdgPmEVt/Op7zF55Y5uk+IpYpgbZYnBWwFICgQ1mU3e7N01P/joT34gcABqZE31WpHkIMg5
whSEN72cmyjptEymLmaFasqak2Sxy/02lfdi7mTzrFPg4/sctJMUvzdItf1zRYH931OprrzVHXKl
cRG6TKGeeA5WHzMpjb5wTe30BXRkBdFDSKyHuxRzFlQLwcj9NzRWmpzKkoSDfL4txqRKTbiKfj1t
TdB6WiHq2aw76AJqsBeRbR62sZyY8bP+siQJ9bL6CPXqpgAbSIiKM3+FQcgF1sXZIW72/B4ChUFA
DNa74saggv5sTb7kozKokDC9UgCh8wWhPR9GDmo+Da+m0PgHUnV2kVxpZE1TepL6b678ScHSd97m
qXxYU7H2wwDGzlHB2lqR7Hvlrw0IItt7tKuiY916E4WAS5LnIoaq1yTTIAH9ryipiiLJRVJBjxgM
wk7g1MGxF90necEveeVVeofiLKK5YupGKjexeCSqzyBL5XHfG0IyiQ7o8Ezdaa7Fo2cqehM043PC
2X/VoVTuFVctBoI7emQ1ZUY4me5sgSV2inngPCTd4yD2/JP0oAEm8DdbnW8MZCYVwNHV53lE2GH9
69dcxkErFhQueGBATDaoiqdMh/FbY9aJMxTrcaEqcNRYsswbesIJIaspepAkR3OhQmFROUzG0wqz
PxsO1WN/22jugLojldPvaNY5gSh5abD5cNxL4HStgpyj5yH5qCiZF7Cz8JJjazhtVlKF/Atlhk5Y
uODm3khxurU4ke4F8dFVNBRPzxHOR7r5/FcLpWjyoKU/pm6PAsb9T653sdmTSeTu81NuRqrq7QdP
n9sdz7WGPk+U8o7QOfAlPvgFxdOh7YM6UACOhwHweNyjp4b029NaRoZf/J3OGuNXpNEY5/Wmrtno
DmMvDoQHoceVPWQA672qo1dyqRGS+prA/ynneSQz+lRWWixyyTsoIC+g6V34xc5YDhJz672IJSGK
4T9DXg+DFmjyMaWIFgcjLqXGr0KIPMwpArNBY/HrXLz/vViqFsLN5+RjXGOvMmTnwMQAFnpACd1d
KvHIJ2v1OAGteEtctRG63xmOhz6HsQOc+yQkJgs+JAZPFBChFolfovm3/41TYt3fNLS34jV2TFL0
j4GTxxw36216V77CnWZ3g5H/FFN0nFY20un8e+xEdaEp5aJpa5m4N1ZqBq+XV4jV5+WdG/eWKWE6
5SYXkHjDGNNiYwvE7Ui4atVwv2rmuJOW7344/0iQpIKkxHtxBgy0MzjIkXpiaFTSJHepY9VzRQ+Q
soRRF6h8zpXgHcgyudt9B6O/9S+ha5OjEMjhDJBi6btMgkW+YnMAhKIr8BFf3TRamoJRU2vKYxGR
/T5lpxfprJEmQIcFJVk1Yv7lmj8eiot0VL9JHv1A7gqFfo6NAalQP6pyx7FTvZcLoRutBMhnxVMa
YleaqqzaRzorp0MFd0P1VvWZFwl+czCfS4qKFTN32VBxvDhcycM7tix83FffUdTf2zk/rr2MhU1a
egS2az6ycwQctl8pXEQ2OmxpkN6B/eNjDcPNzVbBzQmzjtiTdhK3vMbrvO7D1Dxr7is7YJBdk+lY
yjPrLKXyeRPh69oudwQg/a9QTo0df/j+r6vRdrybfRgZctnnwpMWU525j2VGp785Hkq0jtFf4qHw
CcZyiC4tFFZPOh++JtpcGwYqitUXj7V7jvzc0OSOd9azwgDsC0g1HGjVq/lDtg7LiIIFBNGxKrB+
31aRGQuIfZdkMGIsU0kA71gcf7gOaP5A9pINtolwdqSt3BNwAxXwRih0sSiSEU/VjC4p7JIxB84u
71+FKzsSfT6tm7JlwQWAtmBqJeKsYU40gnCUYjVM1mziI+FLnOPSQAUBKsAoN8Qmel7oiYBW1E3y
Mn4XqfwUJy91oX8NesDApNEYXEUBPZKm8vV2uQDP4QvlUMDwk+A2MZCk4+9adgkaWZQ1L3jw00VE
+xED23G1/9DSa9fTCTK20Q/yiUI7/FvF07lDZt3qjzK+2iMlHV9VmApmToz/e+4NnfF7iKvxFan8
uq7F36msbZLyOkoyzkG95z5OtPl77x+4k0yYhGm/bbU6vxK4KWvdtMKmz9fH2HkXZB6WSrqBlKS1
0dUi5eaaX94fUracyv5mCMEnQVfWzIKwzrBn6M97gZBdh6nV0YXMfMLDRvUz8eZs5eeNqyR3Qb2J
s5J7Vs7wjTrg3KotfzEPLqHO9+d4nVKyc29O/drODJVkToLND8k5uuGrKYDlAHh5OH4vTw5mZFkk
v9EuZLqUUOKyp26ugYhxY4p9ccAfwW2OBYoXxVSrlvQpvr24lWlr/iod9jN1svdZqwlencOJ3/Vn
VCEeto8c0XkmlSQMZJG0uIgOsItUbKHwmTvVzs9DDEiMZWJSyzPpgLworbyD+/hN+i3rheMyCjgz
WozgIvTFd2cA/wn36f75tFEoQMjF064WWlppn0TOHNc46BPnUqj0fHPvc+YkiXCvrxhMI9SbYIGZ
pbEUeeC8M/2DPvd/VuZwnhVsJSAj9/NcnVle1AEBNjDCqVCN1Xh6IzW5dRDJwEHvNh4BgQUzsKjk
ccdFdO9+DNra0Y2Xto8CnmYkPCwhp7SDwyusookFsUgWJGEPdVgcP/L49/SQIKVWZpwA5xAliOfG
Uwt4Ye4Mnk1uol12DYLzcHjgAVilGYyUImVZmxKDwj96rlSf0e+dzA4ZosOZl3GITX3V1Ff7Vwu/
tbc91TMs7O74SKTbG+zZdLHaGD1x9x0MCytXREEphYwDCcR8sSX0T9c5FTQm53EBeP+xnT0MbnWA
SSv3IpizEKJcc12mV+Qlz2NXY/a65b6SM8i0JkMEpPkoMQm1ZfiBg46kAlCIJHgvsSB2DDNbBvJ1
bPNFOCXuI4ZEIjeLtVszpA/AZgPxt4zvjW6Pe0Z6l6BHKQO8aDUyMiatGAszGgoxcQbPKiKgvrKA
fQaCgkvv2LVDsvT9BnOJd/8BRywGIu+ykJ1iogvRkq7gWSNZE3zP+tl9GqnBw/Gwnl1I/cFOrPca
mvXiKI+ZO4tlKtuHvsBUlfOKUUCgOKqqfhczrJk0A4q6hv4NoHBc6JsONfEF/R834T0fv7r4lMQs
VcSag4hzj9Tf04pQMmjEgWFP8iOPEAj9I+NB3k48P9ALdIQ0GZONexWRDRXrEECBJbz7c5PpHGep
wQRTNNCBOIOlHICGMwK8LygmtThal3blt88KqPc2mEwYfijO7ppMh06EGvXqHeN/baUeGHZ5pY3K
FFiN98eVYJKNxEy1x1XBItBmury02TlvYQcrWCZ08XbDxeNSD1OuyUwiAX+wefl1of+0I1Nxuljs
v+Le4VwQO3eenWbpfr6VjNLX7UL1PhGXcwOuUyD3umSdHPyvDLzkKA7ENRjPYFbfN5TDHKUTRmBa
TDsVUjZYoDqEAVRqJmxMO6NuIiPzHpCeggT+Ut4p4aFgEFxQNHnTiiz6HK8XN4FZue3xI83lKDM3
I39Msw69ri9j2Rwjov3LY7BXOzoRnA6U67oem394V/qF+I8HOEBUsiJpBJI5UPxDrM9nlAhdg9V9
e+0BQUMwc7kDz4b5Q62XU6zSD9VjxANRKvlJAds/NSliuMySDxpAckhR/PXrDw0Pkh2a8SyZkI1a
y+M8+1Hj4T0YXXTWtni1P1W0+yHRIvHq4IirEBzUTuIbkWgNRQPS5p5yxcIpBV9uR9c4uoU7tCgq
aCC8tOCz/1AmDWeO5I6mbk3ZcM+/MY9vIYXm9LFsEkHKRER4XO8MjlDlraaT/VBbs1KQ9scaEdsr
fU4zTcK98ogzv2JMqm13J/DkLlpjTz993Zv50cSmKxyDPWjv+ET5oUrB9XPhO9f9o6nfF6Ilu1Lq
xcpyw8Ei7RBmf2gXZUMlj7Axc8Dv9yFZl8hj4wWKPrgfAMPoIEX8YbhS8lNKM4C29/emhmQ1CPTh
+DCqNVdiA9PJ5DqHZLfmjPq01N0dVJTEWT29alAxPH6hYTqXqEd3maFoBi8QCtdC7rBzf86DGaVV
kYf1TxqYoia8B98nMUKNTheDTX5DDrHFbCx9EJTkP2k6nl4FU1jv8xhD6C/JA0np/V3g2KQAWfym
VWtl3rT0GMJOlpeLaBrJ8Sy1mjlmUq6lCBE7mn/ZDqJQP4FfwKSXR6QLWOjdUjtuszu4c6fFziJR
rnO3BTWejWlp/flEKDQPxGtSKX0uVtimjQXjK1+jIJhwci0ZCdzyVpIRdlqyEr2tRXnuxAhRjpAR
L2uVqDwe2LvOeZ6pdMIaVZrQD7PieFk4R6bYJYRze2ClpIjUwYNo8EAvJDfNtmmGKw5k/HNcxCMO
V4JW3VVSnfZcUvqUjOdsQVOyI7I3HxdsszoPl93K/g7qzIgaCMt/bwA8erD0lt01plYi/HxAzUbt
X8RgXPfp3BSkmpJw8mSaafFcvO86FUEPfKhxIe+Lyw2b4GrISuN+Co9zEryqTHkUztp2uhLnjTKc
/8dff337C810nqj2iXFXaUy5JSYLmDw/2g8LguFwVXX1BYAN8rxEBIAUSVbXNFHBPliNu4Dw5/GU
rSokflLvNH6Vz02hyeldCJqBtEq+Zxx2xJWHnTQ4c5YZ9dtoT6blLP6JOOwK70GeRMX6994C9qV+
8RhvXrIiVAUqLEYiE6rn9+fHHgLBHhj0XtAlD/1Ix41JonmojZurdaEdnol7UfZwKv/n2x8g6DSB
Mp3bCxZU6Y2AJcBkTb1rlSbHeDOuFedhGW7L8ACbikxZGXoDzfksxZwLWtWW+Nhqh8PHn9S3i5F2
JgrJjj4HAPOGqdDVBigHvmD4x68xIYnA0QbXn1r5zn1HNEg45+FzQtzerIpTgJvdWBjVNXN1A4gu
P+SliNUm81agTInbkFfv2cKaRAVvcpCIsS2wbp+IpjlrkTtipcSPYrT/LaGWb8UyT8sQZV13y0Ba
HmGmcJmEgh2+m+9EfgBO81Z2oH1RQ43VdIz6Jut+sl4xMnZFF3MUfgSQVTA7/rBz5Zf+AGWnHYaR
dtZFf2uak/TdUp74eDJd3qjz5VS/d79oQ0sh+tfFAEg7YFzbZQnnoavK33v68QVCxF2/AziwWgzU
YF+5j7xhg6lGkkH3BUZL5tWNzLmJ7P+YTtjtqJiuw9Y8doTv2N/HYs7CPj8RX8ma6Qh+VCwbqfeQ
V9iiDVXhAtJSZuHYibt6sCu57hMsuGxBQdKqR3WEV/QEecAl6QNNKx65yM/Ud5/im7UrzOULrFFQ
/CO0AiSC1diXJw030lxJpdjoy1rfdFl+qVzt9xnxgKrgAHOb3HVGfdMGJDNr4JXLfKY40fVqO8zJ
HDPfa/+zX+md1Q4jVXvmSOTInKnJFQThc2GOqndczUBT8wPbhSgrYpZzVEFJjym6Ylm436Oc/dZi
6CePnFpd2vZJ2ZMvjaRFVX/v+nN4bOp9252I6XlTJ9jaJvbd7W63T1QpGkaI03Nnn3qd0URqxpQv
LgqDrclZBZ+3QmaDVmWgAhiXjnN7GhseC1nkGPN57cTqsGHrDBCWKldhNVOEgGSejm9bErvJ/iDO
xMgabMa8ooX8N6srNxXeLAcyPvhxaT2uOJVZN7YlJzPXjjYjAQjhz6qDHXscZ6XNL675k6vff9ax
hOsoTWPJowPLKe2TTH7i7GvtK7F921qQOFS2Oxo11w4v4IHp/MgzQn4gAR1zgYEjLPwrAwHdwEaD
JFsfNNIaBcmFYjLfmJ5QCik5wOEPHFjrD129ojvgy9hAEmTyXC07rqCOX9yGRiXqgi7TUiR4Eafo
t4BRfRQCyjgmngExwrdCURcEUxvUvPdUV+smyl7jYGwTmcTtDmOBD7S5g9ei1ZNa1WT7pEn0mASQ
5vEHs+s78XbUn9Iuytt+6WsudpiGbsDtSf0eIfbucz0BfdKAuHEKiaBkfJxvCbMI8HMp97H+J9Rv
NquLKSz92K6FNhA3td4T8oBsH9blk9GhZraBoRGALKTqMqv2v3dgIabvAM4VDiXFIOAxDowvere+
veKUgZSrBxpysszzoGo9bpr2/U18C+e7NrCWvBDUujIErHrcL6iZo6cOZ8FHi1PDD1O8ZfUZoxqs
buWUiJ6jdQveFtpZUxW4OtP9OeuCKR2HaH+tbZrAkJWXlXihmrMU8o/zjdsEhKwAcZL/tLKpHVJs
/HDsYyrfXts95XD2yTlQsgq8OCQ7A5smI3+HPie5oVWeVj2+kzYXj5bMdDEK+nk4fg9UC9+34P3z
Ot4OHJSeWjkiIiE8qWPxXOKtq/p9y4wv4/RZG9ejGWTdoossvTjYErlK71wqrVcGffdG5cFmKopU
3emGCuNBnnKnU3mEvUgrOtHPVnFqX+/yDclSxdXVhF+hxZkkWvH/RA8WqZB+m1ImoI340NAT5+LW
zlb39y6JoeJ+phmFaJcsDb7Tordh2AMFSeUdpbzPoDb5K2+XCf4Wdk7TOpVVLEw6tdyDTJby37Li
awfQGYZj0mDSMCKN85v0KFWt145EBT2ArZ1PNRY28CpSeHiZhV3TCINeYUGzWgC1Ddva5qqvKbKJ
TRleK4HDRGf21tJEpAXgGEFgzSp9WcOmDdPJyura/E20iPktjmVPJfmyPvKQvNuguwvzIXAdvdUe
NUKkQJUocy4nSEGFZZqStRF8re2KEof+RzOwMw9ysxZhcXoN4h9HAKmofiGlTCA6l8C0bsel6q9+
AuLfGphMGuAdez9P9+T220MV0cbJralfsCF5kSw+inA15zd+yTK2rk76p6VAdOuruaVd7+87sIFf
Fm8QR4eOLR+a9Xqe+Qj2xM/YwFEennXLFv7O254Zvkt7HIF2xnxMxlabGCUUVfEXJBgH+o3QzJGU
DNdg07ZZsidaZRAwvG6htQuHkeR+6Yu272bvXjIYdCyoCBKrt9BTwklgVtle1JnhqZXX0bFxXC2y
I0ukPm3FI0ACZ+sVJKcitwKFHGNNSbp5kLRolMY3zwCJesWE1QsX5xM5UboXfZ4wPTWRW3XzmkuK
KjpLGzEaUYihGlwt+n0UufJhYt9L9mCvFhqCF9uqqP4B0GlgiHg4dq6GKhkLlvsQGBdxBR/ZKIGn
2Pzt4yFdWjAw0gL1alQfYLffstPIxQiEKEE9zdPeqyEef87zC6D0Y8yqQETBUEHTBcP+J4SG0jdb
cQwBvg9Uh3LA1a+nuTIPqy6KEeLLZS5/53uWBBfBCtsfH3jMYFUjsjaJ0cyw8l4AR0f6x9ywccWL
g7EGkt1S3FqlNvOVKYt4ENjO62j5cXyjRMOGbglUPOENO3Lq9oIX7IZtAN9q04KVtJIR8pa1DDgV
Toet9yferPIolXhq+qM0l/DgADvUDI/BR0zYy/lb7AI7URp0k3B0iP/4wKJtlf7GEK3y/vuoH48g
bqoY0ZsH/Vwi3dalLJn4WMKD5CLytOiJbZXmEwBll1tbLpbv01UwQ9G5tnAP/KD34v7/7sZC+/y3
phnWvTaE/7c79u12FKcP0UGGVGuxXNJfdP/bQRK5iivCYO2ECpVYCW8lRdsf3jDqmoVjII53gJoW
C4PLjB3cjQCCXE0igypAd2q4hLiseeHjzQac/PN4DkC4nFM+eeDnzx+r0zv8Y3Q+Wc/Xqzw9HT8E
u+WaRozXC6cvSms5ZXQJR2XqtDdTZSwz0WQewpPLXKaNxXhQx785SBcc6dyqH2OEf+Bb6KSV7qOn
qOKB5rR/Lnk/NQTDF59m+t2WmOP2BI4skrK5SigXZQo/NQD4NIfG4/jhQ5TWYphSIg1c2hZ2H6BF
8s2m+Vh1ZmynY5VaDw8P4QuEktktCsuvTwGjz8A0Nbf0hqEPg4mHjeJIgWZeWyQxDwlXjiqRdStd
X+ZVaeclxsfbSwkyFQIpJ9YvAHW8bxbTvX6aoEdXRr6P4ZKJ+MvQOHE1Pe37NjdWhfXdeONepaRz
2U2a3rLWc8Kh6OGmcnVnYiwKKVRVlk5MMovBGd/dXIReouHBoeoDtlRcY2Igo/vMkx/hWaoxQk/8
3+40akL9ABBg2D03PVyD9dLsdV28A9dQBhS+pwWdJoQPk3sw1ql3VB8iib+m4bqntbOJ+BLQuVK/
yxilDwRW2dmnFOcNNoGd0DpHj2b1tkmLuMrNOwP4OThJtLS9UjZO+LgfQciWFFxDzwyzIVFohHAN
iidHk450FnAuUm0G8pMP/LF2cBBtq1xc25IQCzHA2C+3Moxn6wc4Wop+BVCcY9hUKJVD9PfbEirE
lfyI/upssqXGRuACvQd1GY3mfkniLks3QaU/6g6RYgwrdZhOq4POqIlaAOnfhXjSBc5MUJ3ieWjz
IkEW66LYyZmYhtroak8NXp1t3AE962j978FdeMzrKEBq5p1l+aRHBVCX5NFyDEz9L78pHu280uFz
3C4K+GUgh2qwWt4EHU+Fmd5lniw31m1f6oD8z03iF5wQi0mxvxnwiBvYGWEbS4v+pn0mrg/VxJza
RceuefeLUvzMtO/kz7NpoOUUPRVlmHwHzGQJxbbCkjkIKeULqWTRpu8DNZ6Gi2KuCcZVKDEWfrtP
AgJIerJTY9E6dNTth1Vf1n6gvypBPrxh08ddDEFPVmfh0Nk34SurlaGM+RYmr5YLEPUHa/pfGC4G
MZl5/avhH1tRkeJhAREE4VxE/m+//oje6Ft7AivsK7WWWk+VdhMpEvwq3cak125xFnzRVwHwK1dR
NMLjMCNdrR4hkbadu6RmiYt6O1JDu0KhkGQ5DOXC9uUoPY8IPhcvaePcNl5wbN6GFnob7Ni+oFDv
7USw/hYBlGgPL83xdR4R8In4l886YYHZAqUWBQh+rhjbnj6QB0YLmzhuXEc/LWznIxOOBtsZ4y1S
awlO5ULJddsIgrCoOmHuX7uO1BC5j1a0rySHycC8daFHJ+WCcy1ab9UZ3NvLjUfYqJiFlMrg3/Au
3mRxd/2ag0KVj5+NJvQIWR8JIU2Cn3q9TmnOetxjRlHmJu7mIZ3SrZXPG/4E6DaXfE/cK7zIEKB7
djczQIdhe4WqdO6u9944+z4JUzAO198j04dmC24rVJ2rhvskx50mUk0h5xhuUnkBPxPA5LqpAt+m
hecGqkOZV/tXj/hp202d2W/73W1PMrt/7vQOHJ1h3FHwzPn0DQo95dR+hg30cxJwj7s1fkxg4Kun
+D/WDoyxN8j05U0RUJXikOphtCutabNGwU931Xyc+rlbFj5haPIkT+mlBIscXfev9C1kdozfk7s0
XBWlHRcYYTUxAXnLNJmnWlr/MNV2QO9UlHkVfJuz6JncN533VppvGIsAukOC1KEmmwrVQhiFufOA
a/KTb4D31J1yEceVqSaQ/DymAJIndYXZLvOP8/9w3teXLQr58Q8E/cZnlHracoxyyEWTCpqIKjhB
KbXf+k3subd6XVGaftmVNXOPBd842eCtsop8gjwikEmIXup4ZPtbDGSHgByO2HPMkZwbvL3cUZdv
rdonQ3zFK/v0M9+9h3oloFk9wRdkpBmDmdjaYMJ/w5fP0UsX3SVSnVyKHcQRSC2BdqBz1cUKSgqV
K6vFHLstkzMjAzGEW+SJyeB89NUcQHfMHR3HJJPM3wnJpseY0k+mkC270urp62ktn8IhTxdIsIuf
5eV70iDhDZFwP14kCgWpmvIyQjA4cV1nVJ+04hHFy0JLrWVW6YdJJCV58oyvlKE+xKqSWVKubOFC
dg6opTpynirxSneaqxXR5lHncUmRD9BA7tt6QzRcgVjznOZur2G+6M/dwaIg/dHzA1EN5M/j8Fz0
ATFcq1vdDMOpCPH5UOPpLnDrcKv1fqFW9A+BG6sj/L5qy5hSfJ8yUSN6gYzRo+fg0zRh/ZmzrBgS
cNe0L2A2Ro/9zWkTG9/oD2vo/QxWGM/IqR0R9KyPZwGM6WSaI2Cu8jGRSgYs4Z8CRYRHITxWbnD1
kteWaOJaiCA7ttSkY2Yp+MHazaVOqiP83uGII2tkvbEL7jlUPxT8CDW2yxqKjDCfGoxu/Ok3x5+/
iUUGltJFGuHjWLhoj/67CSva68evPwaiu1PNGXbVeUiuagZX91Tdq+8Xz2jTtGMk3uU/cTRBmcxR
QnSwNGbqjlZ8Q+6IY/hW5bkBFlEEjOH4AW33N5mX4usl1pdHb+V6KDTBGMXKyCKbQ8PoVmrq0rMj
MWpo8HE/HvKcXttTahVHjzEElNke29dnZjWkKqzyYgKzg7p7kBGT7LwTnz8eAZO3wGjA8/XnJHPB
iKRH2rQM0W0u3moBLer1GSi0m2zKyZVwapJ/gxA/A4JSH3NV/Ne4EYq4iPPe00u2RVR6PWt0TP0Z
bX/g2w28RcbYScQ+G96ytH06fMs2+gax8cgFiQ4GxFEAylXq6ojFQt7lDFTjQijVhhCMdRIecK0e
L6IFMhQA31tx3p8lWq3ez9LHPPO1Bxkdx0/XY6ief6JUiRhxyo7oIWm1FJVMB7Ux3z27+DPfM/Cv
krln1dyyimxVPk1r/77xJhZtgGvTBl680CTkUbZlgWIX7SWajOKTwSVX77z46SqcLM2N/ar3KYQ+
MaWBbi3/OHntchvbiencYYcaqVAsU9OAUAOTdCTIaByVIQdE+93mOYaNYCMJzVKMvbpWiRO5vnKJ
eOYIbOA4N04ZHE3HI0GJyxQEpbGgw1FZvwamHXZc3k7NYc22SOGDe7VvXTChC+N8JONuUPGvItJu
Vm/REEcbKk4XRUx+WI4tqCuW/TMLiD2PCMRsmt7ZbiuDlWi5SCWL2OjQYGWbXCJd4cxKjqIU/VCN
cLlDCLcE9dpuBMWwLsmXW2vkK1SHCRti/uDqBRnaxCReBTTpggbUaMu10HsJpLCeiIEd90m2475x
Oy9+xSRo9zX3Ux3kFjGuSI98WrzdwiTv6mHj66HTm4qgbJpp1HAnoGcu0zGCzx17mGm0AHxrGU/m
7YU2T5Km1auSOexzO2WZmKHpx+LSDf1nJwRxq0GrY9s+cmmyR7PeVXVI4DoGIdR5JoJTfV6LA31z
RPc4uc3Ga22nc6TVPvDNzG/eCFsUgKKxDG9ziP5eAAo5myoKzHoX3o7B+bqWGX7YMnsoU/4kYUGD
aFrcwqVhFs79tWDkdEhTVzLZqJszQIIU1jGJlRQr8XS2qisAi2r2HZVTsQjA4G3fTxycuLym4FAX
nnr4BG8LuZzB9b9BqgQ6MG2aPmMF3Qco+sLHT2zB9YD7HnxlFrt3O3XPYR8+/0h1yuS+7AE3X6Nr
DHjt25n8v+kfOOcAF3e+5Qo3GLmxdrtzGF28QzneEXHKfq0GayNnU7IHFnoTL0rv1gPa+Ah+0QKk
W5ST4EKMuZlhiBqOeHW15ZJekv57Kc96VK/J/Xahpq1ErznEQqZ55Apji239l3bCGmCDdppSeS+J
QzuvSatKDovajN0Tolp+6qVZLBN1CMLlIsKMtf0lPEWBzYWHjutbybn4R0yKnFpVPAWr7ykyDTp9
2FUZQ5QpVifJ87VwTPT3FSaEre4OoO0oJzrgesdzRtJvt1eqkiu3FjGGPb0Mxc/cvBZFEoerYO09
41C+l0i24+axMi3MLzlWMtVhAEO720le6fFT6b5Vf6Luc2MWy5nSBimjgh0Lw5CngdgeVOfEac9W
V7uG0aQZlAgmYfcNxi2mbYEJHSzLrdr6Sov40LHYqP6YgjahSDYMiHjHvcmHb9bEVndK0sSl1dR6
YIThxfhL3pxrNIxJ5hSG9sFZI72aF7ElIny1vV+k84Mq/mmwVgk7ZEoO/iu2uqWVEP4rvDY58jEV
GZo1NhhvacOMYUVI7sMT7EHGX4Dc3yi03xV6vV+Sjtlx8O7OT+hjPBobABvDUpFVsxyYcI5lJbsN
D4TxBrddVfgDhz8ByzDZXbHV2Njm7YC91Gc9s1JfMCMl73UL8JocYDYzQxrySAsOmRLTGzfJ9C5F
7hzNPYGnC0/GRuP/dWtoRIvCMwRLx2OohwHtLk9MYVD5+jD2aerwnqOwmsuK1I9wHmZ0+J3tAhHD
frHGr8FQJMlNLZjUVvmPmSGfRLYwoPTwWfPWd0oD6NV3HAfBvzguQIzZOsSsyVHxWt1ela1MwQ8C
Fw3HkgTMIa+4FRHGh+GzwSkdhGrDbXBU7gBLL47wrQtZV4EcLDDcM1HByAUk3EOX1O2UvucW/p+H
M0A8niWSfnoazsfq2ZRKb49VKNX0D6Pc6ieYYWk3+E/MZNrZIyxhwZY7F1f6nZQuSwgNI/ZJOtJQ
7N2ObXLSKdelspCsqTyozi7JhColQ3/+zCrKgNO0igcW1E6JhTCKLmyzd8NhUposdxs1TV35sGb+
Od1RQNCP3KU6pgsyNhdAa0vREhnrH8aTvtiz1KUGPmBtBLuwvFZO8ZfwMUX64bEczdH+GEwgJO7H
p/+RHxw5btwWichMC9q5b6j7JJAFYcfA/vZWqVtTtFFG3eYBOdNKMqjVQRJhzhK7M4WFRn+BDDLX
AGtrVHJxmq38wcbq7Hx3w0npipTVg/rTmm+HyDycfhjZjZUZdhDtQ9NOf0OsdRFFiHRO2vsC2qOh
5VQRVNZxJehzsvfORhuOj039rjRCH5na2cewIY9hVExbs1d6xUz9NVEnG81ijMTo0+2PmS/7mR3+
EswbF2GZsTnQ5n34V4IcVZaYndwuSdZ+u3VxDy8YtzdYB35DaMzdLENyyWDcKpWhSfonYCTfeKdd
97ABhJWZEoqlL8mb/VkfMdR1eCQENHN+ad5Sm9mYesQONIVQHqosKeHiTn1Ekz0t16yHUZYh/Im9
2U1NhTn8Nag6+W+eESc1OGQtmvgML2446YXiAxQQ1REBy1xS01P3SPQp8v+2eW5tbXQxfB6LZdAN
F11D/4JNIFr2fXvY+LMuTHpJjaD4adP/bE8dHmsPaIkutmGrpOaWZkw9QadZQAyIsVTnLwqWwCYq
AqqbMw4+BQM1WPFuve8wkBEDrZQNTk4yUIiP/I+gyiA8j31lGwZKYAFEK3iBmBdrCVDki01dkWGw
+itsx+i8VYk1kcIsT+rmN38hvDomIUucL6i6OwhgEdGdrboL7bkhBdDLlFdi8BUQ6ZSuzkhfDFG/
YBkVJvXOEGoPhRwfWf+sDflPUKGmFiFHCn4I2pigwu+6HmdqnXEmaQk3f60q5yRGcW5XEScWLsaB
EjtSnix+/MXFBSGdbUxzxjsFPAFz+F/pdws0jKwTPsf7nP+2zAJeeMpK93w6EG8NtcFjL8xORX5x
NHtmari73ACuV63rZtWxaxstgjliQ4kugdELw7rkn7dq47YGNM2n0rWgp2TnWeqafrdMR8Ar6PK8
z1RO3zlmbB7ZD9VkMfdud/gopUDjWWs/qiHL9lyzTYpEdQmzgJMLMnPy+cy59Kc1qCUcAriQjriv
rEAyWrS+0Ps0cfOGF0k/dYH/mpz/4bFzVg9Uw30uUtVjpY4xPo34yPcEweLnRfd3/yTpFbjkef+5
+b2VPVnhDWvzt4iInszyAltz53+P8nwIcoF99qCT3GR56sSinQRifUTFMJFnnOsqFm1Q8tFqle75
S9vE2e8Kzyz0tpGZ62th4KZMny5hPs1T3qXz+3NxYemWaR6ul298xPM5UvnPBbnx2bo2vZrUQbaY
WjyMljuhO9UGFu3ZIOTTRnwWOjAr6wHQOiSzJajqI40mjMApNlneyp0OfZGsbVpzeGL0SxmnrTFb
y80cGltKXWiaKx8Iy760I4WAlijOYWQVSONuwoy4EuaQP46pTLzNI8+6wk0xDWCGNXElZ+Dpp8vQ
BxeAEXoDxphmCD6Sts5Dnn6CHUFSgT28+Ajw2RtUXThGAEK58M3tdi6xsI+QuxwVaOrRZf4Z2SVY
c4pnlRJZ1VpkzSOC6eWuam7YKHnZTkKHLXBga68vzESeimm/yciu4r+F3C2LncXKnPVSjEON2/8/
LOs70+zaQQiWvPW+WZYbqD7RL/71L8XA/S3PicUdr3OgXoK8c/o4gFp/DwU3EfI/3Voct9bA8TR3
osA0WqnedmIEYhWy2IbUumAVR4CJDfHYLWBhHm1rHZxaSYK2v1VLzNqvdiN1ammdMzS7JikvsQnz
8V9CcsJrsx3m55e/r+p1pxknaubzlo8LRI+vLQRkOaKuIoVe+xHpYWE+U4D7u+2Qnbpu97tOHyZ9
Th/2Ko9PNVvUf5em1uQ7hqhOENPRSh1qdlljkH1qXSFMbPO1/vCQkMsw6kXuABUBcfpcKOUj0Ag7
1bdyvKagud4rMbXRPiCOi+IBU5nqbNaS2FB15X2EfGtroJh3e5DOv+a8YJSjQFdF1SqbV92dgZcE
zK1qa7MCZWLtjzI7pbWsFfoCo13+g6O4NVowf47DFy9SBJdFtxnSr8VeRO/L/vBdAWeBDIJRE0Ys
8mSRaEu+j/ISmwuxUZJGcbGMciA1hNWyLMhwa4RtpTW8GWps+dDLKzUsUJZJVQ9ORLwkX1Y7f9vA
NEqqY2SSbO14qimJcmb5DcXyq32edGx1fwrjuXD9/Sgh/i1YpbyuhP1zE3MWs323paptMX6+MC06
6uahBeb1QJI7XRhgj4y6LOqTxeeZstBpAHLhzzrxtbJrT7n3cHB9EBirtz+1m00GUsCMEW9rUpMP
JRINtFxiEa8kSYzHwa7iPSWGPuL5uXH8GA1bw9jN5ju/eWMwr5CFTmD3+/ObZig1/uO+x1m3rhyK
cmcD4pNE+qLTnNxWRtDAgMG5RLM9kkt9gXkKW42MpJnXX7W8A1wD67TKNke+lzP2Z7j19WGMH0in
vxUp40t1XHNocoKcvKfpsCmZ9IvUDnkq1Aw2rK64diw2hZWNWm/zCk9TNOvdfrD1zXKZ8W31jvNc
CoI/zXhRcmduTmlMP05fhiM2Bk7ogstgEm4lIptWZzASG+nEugXanZMk83Qb+r2iz+RWWHNpmJgQ
tu1mEi1fjTrpLqvCReVwhtqyyp2jQWRYwW2eAESPitalq2NB9SdkiCeAzijUiirpQiJphpkAYUg3
LmtGrngLDjhdpEP7KeCWNf81niwNPkbiJ6QGIMt1YcGgLYiFNaE2w7gs0J2YUe0dcZygR0pLkR97
3fv9NGL/7i827PFdwY7PEBYKJdi5HXrbnyLvRC+FKGVcW5VNrXfADJ3Gc3DMwDV1Vt8G1/FdO7FA
fQYXP/hyRZHQIirv3Ac19uWJWPpTOsxprS6U5wx880mtpBDPLNfC6HpZYAVqFns62GJUWWKFnpWN
EGT99OJuhQoV0KfpZ/qAx7QZQoOykiZm/evXKgtm2Rk9kOGDelI5KYHdcwRRmHFg3FrHHLHZzY/F
TxYwmhIwJ9+Qz2FEeiSi9GwpurLG1flwM7frLvErmIRRBBxgajo/JOvTDhh5ibE8Pm4DEKWiJG/t
MAdyLaHAnMQgeDpncrO+HAzMYizf1Peg3JsKYKYu9YByYCQdWpZvcvCSnxUDF38fE2Gx4GTG4Ev+
+A0sBTbn7RFrfikHraSl53ZrDGzQiH5vwIs07bIYIAL3v7fWz1jN9gMR7Dc7JqDvFU0zSGh4UBL2
Fs44GcYvTmb93MfQaZ7olvzopamewp6JUW9EwOkGfndz1KHfUCqW6E00x3vi48MZu+Qj/fIZ/I8I
H4Uww+6xVGhFuVV+s/AwDYJhS/fDXOINYQ2XLIp2b61TCNkuRj1ogdlcSBirPkTIS96FgyypDJ8F
wCidEQWwJiE+aggmwlVC7ECYwOmULkC4p7LnUTwG4xTg2rlXMo4e/5wrUfjfR29X25VAy6XHIShw
CYqEHqkfQbjqDTCb8DI617uCJUR8XE1YygI9KSH96YpZ4ARRKNQSp5AVk6myFvEcowC9tetRaTER
twq6cFnkNq5PvWYoiJI3gj/64rqkGHP1aACGh+qH5W1n7NeiXqau+M/VhSCncWzLPigHDZA5lgbq
HdadB9ekiYMOYgKX5VhXloSVIRb+tcnWVi9IqQleRWkkYs7h6U+gxzjIcaLVXW6ugs1HcIv5rlNM
rZRRejt+6fUzo6E3w/CpjqLBoMRLG2T/O1qyeyqQo+LSAQp+hO76+1PSWRpHPB3WlcR1AtbjGaFL
owh3BdPD76l6qBGXkULWbEZxY5kxZf7Nr3RR/Ti4iFuo+OHpA+Mmpipe0P7fD+HQAeUsnxVmG0tg
Z+hzN4ozrx2VgKXWa7fPkmzLAXXDrSN2oXAK2nTVXA9chc39ANs55905L1F5x5oj20GjU+lPCyzz
A4McjEP6nLS6Ec9fh/+yZblW8OCeEmmUJVVTDD4gk6bth/a8UkCbhYJDAnxE86Dwi2bE+KTrMPci
RfoSYF1vv3cfNSUnr53PaI+Ma8y1rr8X0or6AbkF3BsBOaNZA+oBi4EcIGa2kMLc45mcUZQC1/uz
D4b1UjrxUed+5LjxbF39ZvNGNUZROpKwPnjXEvL3Pb3qm8cJwYHWQpxioO3hwwFVeJTNhpXTpBlG
Dq/ULWtHGBUnIbfL6KC8nl8+wwcE5HzhVClprCdxmXOidIOp5JZI6bA4kwuSLtwaSgYt2/nUWWsB
pA1KUK/I8iU/RDw53wgagnc9CAyQ+N78vDjdekohahyiHPT2KyacpZgjELdIuSpTvBuGFwNCvJEp
PGVsNoYEQnIztAe09u3ObE5Fv5mJgf5ksCp1DYo40Nlx31IHizQVGxN7GRCEdtcDuckljlOZ+sIn
EkU0xC2sVm2UQfWZ1uahsfFCUc/fDHFsvH/V1j/I9+BgNF9CoYD+6EEOUmjIRQDD2+Iu0w5GqMYx
i9kLkXH4M8abke6AgesMKoLtBUsoZKLXBrwW8fXGJZVl2RCaQ1Tk+DkK6HeDEL1YpWfOyKG9beRQ
edKp2AH6PwzqoKiMReIRo2irD2pMFdIKMTwj8y45Tp43efiKphTrm+j7JPVDQ6N4wnmgRYIMGNZ+
9ZiVXAHVVhG0+o6cbzmeFjv731dlPBRMZ8fGqqPQmyKLU5QcFroROR7yPnO8gJrKKSV3gxdXdJ7P
JYSpfhGILtWCjgVXQPgbYmk4ycw39BWnOK2h6iVJvlnNH3f11g/dhpMR6uvSKuZitjxAh5wC50s9
bLzVwnVLbbp2NyDTnix1FthjSK0tiGTH1Hs2Hs5S8tCKglfoj/J8bHFiXRDmiNsq4huAj+F4CYuy
S8GfMFxKzpZa/DmdXTGAFpwMriES6qYKPlPqiTJtu58IJAjGnGV1ARHDNjadNR1erFq4TIziVeKP
p+NpahQPFMSrrayr8hC+LOxgYlfY+lRxlg/D2awBvcm+uKtC0xL7OzIcVpmHJW6d8ISM/lrkXnqp
zA8xVTyMV8ObNkJft9l5M2xTPZAPzSu99br1GjVc9hrIABxeH4RZ8iHJLUjmIMUfeR8MHOg5dv/U
9EiVkN4AHjQCkuoJy8slgxG/G+kw98YhhrK2XfXY2uNiaSRiBIlBarMPkJtqwWZYJPMBaS/8MNz6
2yf820QHKT+a9/LWuarnnzO5ROhgZ/NqTzww/PzmoIZFI2WZUK3m6xGqEEPc4qninKPCPC/8zeMu
aLRPZNMhtKQQuhVlFiV6wF4bregXI8NK0u3+o3UWNv8RYtstTF7gkIblMr41TcXJnhoEMCfCRA10
MF6Qra/atLdLp6tHh6tyckweZX8YFqK5umLSohEE3APE+Z8TdR6kgqme3vZtN4nkSkAP9VhlQpVW
IeM2XHKQEQIOngXSOl1F15Ga9lU209D83XGSdEfn2J5dkC4wVeg5Lvh3/WtmQijSRxSQU7iIWUUs
s8nvJersYCoMOXZeEoeWIGPMUnmDj6hHnj1JUA2yuCFGamFf/pQNI6gcZ5lc5HvI3+zy06Xx2RQm
TJoRMTpHAOFtKQrpMW6btIxk9aV920MUQx1pjtgGELxiJHfPqZ2XblnsK4Wt/Hmo8sg5oMrVFB9y
NIQN97bHuQMyxSV6ysCngRzqaB1j82UFvzHKY8ZlIjlvSzb/5UX0edNw+SWt0OnGIwIg+D4tnvvM
iwhLtZwwEaFbujOhyN8qPwLHKcrvkGnugIHoU2j8oChdTFN7iVgLexW1VQUjT3cpOPvyP9uqtrNr
vDy92grLjQrODj6bRzften5XiUsmRzhWr+WZ0hPMiZZxE//wbApGgtUbqYg23ojhwdu51IaN2kBv
CYsQTGFnan6cqBLIMDTJiiDcBPbpmtvC/rqlgGNZdyqCgTeCKrRQpnil6yBJkURniV1jKgp+TVEY
DXW4NxHEyKdaBR9RCvN8W8ZQREJMt5fS4rM7zYOaK/98XkXo3GLUswK94o16qzByRNeCYzd9HbHF
FV0yphn+XL64ENZwAoChdArNtyhZkhKVd85JPF1ue4KjUHE06LsTMpaaY3omoGpxVGZXy/9jSbJC
PpWmxcG/asJOw1qNE9wCBl3bYCmx20s8tfs67N1IvjmZ26RWFqM9CIDUt4nXNOQmwSMqk4n3xcdi
8R97GBP30PqUMohKLDrrJ7DTiDiW9APmz7DvrmNAKq6ZwDZXcwYklP1nKWMIX1Ecf/a6OK03i9da
kFCws3bLTGHv4Lq5wJhFwGHq1ZU7aP+gQPSKeoLm7ajqlCMmltETfO/vH8iTx/r0XOEMSAWI7E0i
9ImKJkUerqkj0GkrKhmm1HW6xFbV76unu5ZimKedmwkHQN4STHu+BvvVDZqaxBRp34CFnla1UYGo
YuewwwYKEWDAhiHTomc6QWWPTR7QZ79GLgmXWN3R4Bk9nNxH6P8WfHjlIFUcXcv+HHzJTtfEkvye
NvoE+WWEIn6o0+LXGUx2wKo/fJsEttnpCB2mQlNKa/XJkOwFMlMChUE2JRhOhmroUXtLivofnadU
6BYWgEc6UIp7RuuZgiPASTLaT15HMMQVcGYlWwCnmQiqrFyLjMGCAIB/G2tTP/3mQyoYrTcwukq4
JH6DF8ngbinT+j3aC2sdLzJUpnK4b4LK7200G9rXxBmwwVNpQ6kKSRXPa2ednTjpQPb/1gvOxjg8
P5GGOqqbHSlfSmd19U/lwScwr6H7oqwUJTKliX/YV1VuIe6wp7iufB3COzFJC2V9KLUTKRbAbaCC
dxSCL23jKgvD65+1vgvurMhR46UTyQylQpeB2PWmPDtfd2MTCO/oKrL8e+JnPKiNUirp6VqM3FyY
Jvug9enR9rIYuWIIdcV3fLS+4eR1u8juYXSAKwslJ8trG2Qt7uVfSiRIK7iOnLM2UplFWxhUXGXc
kxdrZJj+NEMJ17Xqp6GKCaXOWvtO80yQcTO3xEK8HJpZizywUbk1B7jiwF+4jZfOAYEPeJAd8ZZv
2v1lBErMPUyq86vNCpCX52/ekeSdrNOHJMNN3qsxsDOBsjipIGiTIJtC/I35iyLkAfP6Bsvqg9eJ
1LTArZGhtEkvvD1u299tpuc5tKZjJm8ike8h2GpNr3AlAdpp1E4E1hVjkW1FHxWFp0BDaoVU7Uec
jUEpqbLJ+ItvGjHnA1rp7OhAY1YkmPsMm4Nqoh5R1wFYmbrp357AtNY9MwgnFP89a1y5KeTNzNPd
YY001LoTVPfR7LKmsvSdFhTqxAiMlrS+i+RpWsOs++6YTQvWsGkAiOhjYdfLPlpOrN0qWO/QbMVy
O8NzHsrKpZ7KB+Wom30FH6QeHic9psSG+E1SEHlZ1v1pdiii6+JNprM5b4qP9/FwkjCefyJcrXyZ
eKCy7FND6lyvDua+/lXnoJEIbeBqonwHKMFl5QrM31kjcJWc7m3PMbB9HlPhBnlk8HccTE0JOsWB
U97Zz+9vkpZby9CbT16HCgZITMblXnln0ESZcofmMqIc7YFCd4CuKtp39J8em+Kj1cGK35DL1MtM
f1rx+Ea0PPPLaYKT7Hw8xSZJNDuyz1jLVyUG0XWu0vFfN9q6RFathJoxX7WR/nT+g7ny50jkB+8f
U/RXZg0lANnZUkWhMqsrXK/HCO23xOk1Jw9UtO4hpu/Pu+I3OuekbZ2XjwFhAeb+wmh2CVxnSM2h
Lk/VPsSgzNG52j04GIo8A9eJc4NLNoEfmtv9wqXy4cU74CdK+xSRO8JQ1LZ6YSsynQWJToUHj8am
JnIo9LYDkGSA/K9DRUt12uXfou62EiQb/nJ0kSpwSCx0kFJf+i9FfxQl2zHy8dTTNXCIiRwMUhM6
qWO5ikxlb7+g++q3oBsHZzw4sD6Of+B+ITvN4gDk6BM/gsbeL8uTgLKJV6oYIOdA/Ei5ZdNjOePW
br/oZVXtknHDtj2c/J+V/8IbWCoGIt1luNJJLp1Md1rWE2adB3NeARdj3v+/TPqx0STQsfMBNCY5
cwA6z+WUVXN1h746oAkIpfjkZ6RUGLeP9fQ1pbXxyFUtSKRcRwvZUXhWVblhgIM0Bpvgx6sdBPXJ
+lSJcmQal274TFNFPTQ2EjpafrWwWhkQjap7ebl75nrQchsq+XSYfPqUjTcuhkFjXkerClzo6adp
JqZd9zdazcqpsBfjG2CFKr4EKWjoez7VQY8AWlqo2pGp0/bEH3PObn7WLY0vZdOYgDOFlMyobPJa
GK30T1qmcajffuDf9OVLbm+Qd8dZF3uW6xf7QNgnrLDNKwv1OCwK2l6hdDyPTN2EGDl50MRNly4f
diOZQwIUbFE2hV8DKmK4+nHXJIQ2Pc/s1PhYdc4s4ZuH8Btu/58WUw7qNxnAes97Tz1AduUHRAeE
uPRGwfcI2273C/nfgFlQjfO24NUnebmRbRuVqXJd2k/fAGIo+yLLrDRydLNstnicGhDitEx10hz7
s5TKuG6NRohtYkFeBqsg3i/ZaqnKj1cWRaGR70CUYabc7kTWmPt1hosRaAPHXWGWATnD2SIXunCY
h57BR3y8w6v/QM+H99az9ZLljP9yBWOKAcZEawrCJipkkXw7MrPHZ/Om3OvHsa2x6eaV9l1yEYwd
1k+JKV3ofnqbOr/yX4xDwBJkI+yBGziVChGLv2rQ5vfwyUY/M/Ycg3HyuPJrWfGPsodqjMpPxC8o
o/uJFgzehdR6qhb4ZzrKydknaQhnRRTh1GwA2SUjwBLufC3WPlCssXNnVHAO3P8/MTqnXmW+oWfq
54lLPyqi4Lo7e7vY1h82CbKokCOQdLA8BBzOYWwTDmmH9JCV8IDwL7h1D14jptMIMpN3fVO1torP
Sf/LxwvJbFPAqFr17Vyb4L6IRYiVcfqBDPohXfLbrXTPpi0O3fxqBTXmsWN6Aoo412BJpUK69ZsQ
PJvyVsaRGbun1tfL954FFxc8DIHa2F/DLKhwjA4hmZfKst2CfTqTTvR2rRvv8FerSGwQr1mgR1OG
HDlwaaCVmEBdSvK4FqKF2bLgFSVonM1RrsAdYN6EyX/gpwgl+qT5kIzJ3tZ5Edi5BnlRmCNDplhR
lADdppqlJR4CUJRjDFO3jmjpAIKhYxllyKn2mCTPTHRdiRL0cbjV/XUOJH0QehoxAqAEpUszIBtz
xFxBg6uIFPvHrWQQT6Pxf/OmbK/FtQeQMLifvMPE3QCq43Cop+8p9aWOIbL4KI6ISswoy/o6FIf6
2nevcdJFjAx8F92ADCEmvD/W6LMSAbI5zX22CseRVNlWfs6bPeer7afgNWBCCDpgZUZeLLzVjKai
l9KrXYI/WAVPlUlNzOrrGxtfeXfYt4k/PpulyIQcJoKH51dk+evdjPdj8j6G/gRgyHEMUblEmyGk
9vVq/mdLVQONrRQPPIy3rGf9aeKFxd4gM6v/vu+U7IVvPfXIAb3U17nKB4XnGdDX2TBGIQcajEvW
VvHArymywCkuDEmLT4cgjaoOc4yXJG2FN8XBW23UGtgdksgIdHnnon9RrMhzq8LoN1CkZfaRNEmQ
PI33i3CuUtsiVxUa8IYXRdlWun9yCOKdjuJ0CHv6Vuxh/a5AFNAGJ3vIKznB9phA92EDZh5y3Jew
7j7z3bKxXclGW7Ej41vBH3C4Op897siUR/fGR+mmDQOqogHd9a7LOmq967IgU6DGUWplidBqxsUY
1/rgBV0uTEfG6O4Z+2QI9nLiZX16ZiaqOQd12tfbcyASG4Zva9wxRFtygjqhUM0CAz8U+pH4THtr
u6Tn53/7rf5zZBJs0QZIe7RpWgsvgH83SirtASJA3Y4BXpTYqQeJ6KKTz7IVvSKW4js38N8Wta7R
xH69MRBGizyDLchLJNm3AEf8YzyvAlKVZ37LyF8LwWD4mUMwnEJuUza9rUrA4UBfb4zF4fnDWSi5
LLbdD4u8gUbOJ+upJWEPTVfSQkgRTR0w/qHPPWTW5whnzOSfzcPuYSVn/Nw+ousjm/K3NEGydJqJ
CrtyEcniEVErYWf6f2G2k3fCloTIF+NhkVLlte1yesTT3AulpnPC3/qhvuWu85QWSnpm+H4uz3xi
iKsK0tCMO/Wi+/BW0MxCwed3q46SHbTV6ni9LTTn9/5ehUiyICx2QuANVeZTspI92LiD1ouP/LSv
XOdRC3aEEUT9TKoYFISvNi+ZDJb7f47SOmNi/RocgBrLP0XltduJcGsE2j140C8UjT9gRFZqaKoC
1WwtVciGs/EPB3n8wBIuZJjPnWQ1vl8SUe/XHUBgF3CC06sNQeAeEDEmhxZQTkTxmikG1MoIENt4
ke+zj+fkSTtTND0qeZMWhz3DVaMCKOiZWrpr24q77S376gm49E5hphkkPH4zQ1hf89hB6b7T+rQ0
/sIsxkmp+nTuvx4g5v3hZasjUzoImGDWkPqkIJe8coqman8ZBabWh5vTCEFg0UTeZP/mSF2JHfWe
UxDa7jVe6+PoQPcJ19cWh0nK1r5OPolWVs108boyuDFunRCNXOLIoTCW0yNcVXGXvF9/IJac6t+I
PdwjsLJOThS2gNbE15k+kZU3X7EBJ2cip9bSzE405+j8cVTz6wG11oG1+BWTIvvHOsLqQ20924AJ
zyr/hxo0wmS12oXHyd9xVsKIpRB+T99gMldWlkUoVC8h1vcxLlEUDxMyqfHZqFbfE7p9+dm8egik
ImQOK8Qqhm7mO2HYXpSWNaKYzz56Skq4EiafGD06i+/Kokkjz+JYnX914T/R+sedUzbZIoEhSUgX
cFKgmxGGwiTrUWxhi89EJEob9lQJQGvjkMr+Aa0830MEFBVY8IKNeLE2QOBX6OkrWQi6hqpiV1B3
OuoBmE7IKdnhfqGfPD3QYp7cvk0REPG9O1t5Aa0NUdlDW3a2oUSaEESM97zrDM09cwF+esUd9MG8
OfHhEaXFxIheNmeJmIrqh/XMZm2JTk6m8yUzDt3Qzx1ePLkw9qItJ3wp+o+ryBdPk/vZyaP9bfad
FlAtRumuubVjrN2SpfMHgW2RdnGUWCgNyYOlDH56IcPIlYMUYhV5LJttTa4JcvL2xLHn9p8hJ2IE
9Ti4wCXFf1fseg5rjNmjeQtXLnHyRJpPc2iPXqJLyJMrKshhDBqmlxenRU2q1WjmffXR7Y33tvvG
M8prWvHhberEMBGfsS2C4BQD3eKLaLVvHKfgFhfDqkFlXYu9JdsY8jpFdiBzckKi/tvQo1n1YX46
4NwKvyCJxdyEhonHCuf+pj6fpefDxigsRU3Gp0ltKcv9bd1rAK6Fk6/b93PRuDdt5tc4rodumlXn
YW4uwejo/liDCBnzWGk8cXLUHPJ3FBGZMcoWeIU4OV6NH3GwQ9SfkGSqbFdar6n7F2oNUk2lkEIL
v8xjLZ3kjZLaWiCVW9JFnI9G6X6xI9v/aKt89ckTssdTvCpFqRi6vSjeBP8q2w05Yjb+pxr7UVJV
Gk7Jtwlzv0gu4BNwfPFogrL9x7ZCdtqK9Uui8g7tlnUHudjzjul7wenLPGKu7zYEI8Gydx1j3jWq
WLh2GZUcmKrgFkKHwAbpoPmopBhigf7kiVQ/vkDvJKaGBPrlVs8jSdAk8qzRQ3D1tq9YmsE/oSfF
ywc5O+i8IQnB/OjJR/Ko6rxLGlGIEW3+gNyoZdcIRG+Ar6Ts+O+uWieB3Mw9nKQ6mFeSM6CeT3fg
zrlBXx6NqSL8hUHPPzzOPfVDHEuGvKR433degG3kg5jZPpeTQqFa3Ccj02TI+KSIi/2bTx5CgUc9
02HWhWaU9LacSBJX0Vz/B6lyBamMn9Xqm4ZfxXnXDfr/eps25bgV/BS2iZP1bArsshjaZeHfqoEw
P4Ws5+VSnq7k4fWCk5TKJj2EDfJYvg48krJsLrBnSBj3bcuOx0uRab7cQj1NIH1OdS+/M2MlmTn+
Ckdw0iubILbgAd2JzRiVRzSpqgyK94MCKVHMMyBty2yv9bLX5b8AJvWtR76mvvkVrGbYD7dEX5ZD
XFXl+KzRMjSBKoyyn1JoE5UgB8KbcWH1uOXS0z2Ht3n5rZ9RrIA6ZToh2ubGPcDm2Fek11iViAPy
OAKX5LGd+qr3CCOw4WIrh5t9SfFfYhkmthpwdVcD2WGU6yaqRx8mzsvSiD6iEuw27HhDymz7P7a7
Jz0OODyxLJDd2GFbnRXvBs4Gwbb2B/KG6GTAjvIfYiJhVIeX3MYNyvE+6TBzbaNFCR1mPE1XB69l
QJVQtbIemT8W4+8hckCQGVVajdikF8ZVFr8SIkXR20v2RNkiiBcx08eWAujpuo7+YqDfo2ZYytRw
aiKo0dLoIv4O19yQlugW9YvwyWKQ7cC2tlvXf1ssKuyWPQJeO6vKm1bdKW/fZT1txEiznsxEs1z1
77nl9thF+hh5ijNxOLuYIwexfW5PQ14agGkCHHC8QLQfJsAbOBj2QijMVjljW8i9tyZVXAzdFjai
+DIw5XI34aLq5ic681Za0/XlZtlQHDFFUC2rf72wVwrlg5ZSR57VEPxlKnU7LyGNsUaLf7fN41YD
ZuYsrznXuWAiUfYvhbaM1ZPHUHOqR8JBY9t+nxEnGVcPRzipgkdCTcD9XMkau2APYdD6/UPSsDhz
Bn+LKMFnXODDIgFJie+8tY5GxxPy4B9l+0+HFf6Nl+yN9HsicUn9JtDvq6MEgFCPxNESuDTSNwea
CgbOve/mWkrCzcp7PlsBtSIyRhjqNJV/xw9AB4WxKH25HF9OJoyG54yfF9bTlboz5//hIno71QS4
Rcq6z3a2CMy0PLNo9LB/zGY0F3Qkced377j4zduPGThQAWLvzexbyHJgSUTl9qGfocZFasgfwXGr
H0b3/HK2YHYTzX0A11SA5PkPcXCmx2V9tn2QqQnW6vtbC5Bnnr9Y/H7iTlXL90TCYT349S8RtzCz
WbMPc8ensV0tdVSUygmYItYDiouY3dLkpQhkEWatk3vBxYo/aeqrf34rSzZiq6935y47axVD99lU
GebOxGVTCUi8RLUaCKB1r4LYQHagvh42qLNW5tTQxOzfXYUlNKE6Qc3vFm3gDPHbhevSfd+HWsR7
pIsuQYKZMgJN+Qmw2bA2tGkWvVXCdxcT/ugGroGS757RbFH1DKfeJ+wSmoWWXzk2qudl3DHk02uN
BMjc9hRcFQK8HmIvgkeQKYJK/24n1FdUXRR1QLRXRy2mRKpUUoKb7GbmCf2wILMdWnZONgGqrgCh
jaurm2dmKO5u7A7gu9akEz9om+7DLwxzCyzPjQ2ra9f+Ls/nPnWTAcXw2kjtGMZkKatNUP9PHU52
Il3igFYNWLFt0sIKIs4kpfUdPCbfdC9oG9tiJtP+L6KOqIrQL0egrZNPRUDD0JGDZeBZ1+8rRkxA
ffzKDxF11LrmmdRBKY03AgS0Afp4NFAvuqZC/8evu9D2bdMQBuOqSJdCKP8yk1HA5nDkMIlyavxi
4UI2n4I59f3aVCZlLG7sIjqCMCa07y7JT0jkc+dsUUicQIPloeM75dtNhzkEprVIE2TFTkoMtpDv
afpgKYJrYifecc1MmlTm++3cw6rJGaJQ6a4M330yTL5JA9cTMdorahRFccLMd2O7DsBp6H+anzcZ
n1TkHeL2E2LPwzn8mmuhoj77kZwBs9zEeKj+rQb0bWv5vCZOE9FVMISIoJwuniqq15XlXqJz5HKI
hWMdJ/U/hGsM5bX61X5T3wJORcKV6lJxreNmAKwL2Yfw0J0rFXz0dlmzLRJcYnMvANY9VWlTX4sV
drvNNJu7Fb/t3KeX7Im/cm+YdmkG9Boj/I8M+MHnx3PN3O6YpGUd1hS234g/G9CdXPVQTIQpgqqG
KyttgiEqeRUar4AzeWCBhJIvKUh0CycIWiZJ8C1VHEYwTpZdwA2S3deTGXSnLSTJkeVqqcq1a6Pe
lfIFP8D3FxbhK1G63IMsq5dLGN2C9jiNCDw4iQi/EjDtp8dqKh38QDux9siGzoiQaAgrakxsgB07
mrJPMyyKPxXJUf6l4DPA+oMMpLnPR0ZamkHCUctWjRvi6K7tHJSApYkhDaE0dBWsC3bCv76oc32f
9UT1Xi9HZ65gMN8rUzM/qgJPHkL0nWwWwU8sF6OHyMKKlxK2SeIWkIm/tGuooAFLNQ69twecVYRl
ePYd4yt1iJQ7rOyu3sZXlMwwopG5EhZVC53xBSEGGWiScciI/YACfeOPRDfdbrI1NyKgQpe4LQGo
yGaEorCnvdUe/zMHtXBe2ryo2vQoAX0+WIZTcH8nONnDuyCyDu0efK5+pABLvdJNkiyH308IvQLX
s+mpXJZ3C247rRCgXMVcRCMTBcOfTXNJIZkicyl/oTFyJXerYbmwkPa7d1T0armHUky7tcyaKprU
3FwH/ws5OR01R9PBXXPONPiwRu8H4YXnveHN56zVeGUnJAWCnixoK9X9m/LWY935A0CbXL6Zf037
pwr5Hqe50A3r3/dlmV2EDnnBVawiAD3a9PzhmZRjg1JkFcJkO5DWcacM2Tw1pbARnfwB/iJS4I7K
Tm8J6bFikycepPXwvmjd02nDmXA74HK03nt1czJuoW8oAHGPuzQqCA3WnwxwLL1PxjVt9xLNdA9W
PJZcp4lU3meIBFD9iWREKuUFSHdxKVJsVZAyr/qpT20XsdCHUbII8azzcjzxTFstQRhDArgvgxdO
vW6asZkJMytsvHM3WT1nD2MEN+muyDegjBWnBfhkyHi9B3gcmsadGOId31P8cCI05ORjRxrK8Eij
rqpcY4b4qzOGkcLc47TQqYkqiuoWK5h3NIqeZJt0nGaNdUIErY8R/SnjY1LK+RLTZ8xYMNwS0QYC
BffQifhNFrW9O3beDR9WuJUeDEs0bhdy9eKQ88LVSzClE8aRzs4Fmn+3Xsj9KHs57ol8+H3pgLfa
vw/2QEX83BYM7i7OoK5QQV/+e6D8cPvQUAbDAspy65g6FEKqqYzrmfp2ee6hge73F6AD8SUlus9H
bnoTSNZm1goT6C07FK4rsTOadry9md1tgo9gLB8OgBI7GBLIj5TpvFCNWlT+eDY/UOB50e8PzKqw
IZuBwjcUXTGZ7hNIHLzWAMvrxIoiZFgco2BesG6dYqHMM6hb9suDojRCoqK139rmrE2vtOQONMRE
jLBKMg1eFhMcDslVRGFHaRP+Y262fBjU8FdOShJpcp2sbUZIMFFxpUl/aki6RbezipKxNovHTDXn
YeFE++aRlBsOdaVQTT5a0O2mvmAk4OaW+o4VgJmbxfCF5hHXQI93MSeV4KmHfO7w0mGQCmwmGKdP
fmLpWQ2Vo8qQq3Ob9o9E8bLC1FVWUDSLJi8/q2QVBTzap2Y5L4qWfc8JQ6jmiv0KAKrDffK8+gP/
jaBIknuyW8ap6PjRu6T9GVrMvzvAaaAWVLekbaIIl0Cn3PY1JUdNo2Yd+BoEt8xFLWUMtDEhQyZD
xZoGpNzbkCECNDWVL1jojXpf4Ei2OZv48t2Xs15NjLNtNo2HHOpsXzqzLDFICIN7KAujSpFo8tI0
QLRw1KZU3plJtaJiPHbvHXDMCHoUNEMAa3OtNqroH42mTIeAhSRK57+0HkR67+N8oWOiSsvOn5ew
R7tiZ9JtfCKAUhdory7P1LdiA+Rwe04zA6m8ZVE09I9nhyqI1sva6BIwh2r6dY3/lTXi1m/xbBnC
fGFn+qtg3p0XXUUfdYDdafK/EYwScaczeG73LBfqebR12OD4V/NNjmGnxseg44J7mOdSobi89odO
JkukYI1hvhbrPM+0RhfXxlAkPMgokECvLQ9aJcOD/AuzkESMZp/PC/CLaFhKBq8lWz1pDR+F4tAw
19S4BgER5o+cAg4dj/St1C8WGpJPNtdCvRdms4VHyNpstvAJ8/CUj+3oyrtTX7dww/P6nV4MS1NV
dMRfh0zwKlj/b4tioXcVZr+f+cU8Y+cSvAzUie20NaOAnquFC+IpviIl8jv6O/56vVAdZYCXiTsi
22AMlYVkh4jiDVDbqiyjXctPzNDixVXJW4DFXx6XicHnA4mPvGcUJw+hIt6ZN3atlvKPFnkbPhkm
MmxMFKX1REUfVV+mW/P2Kd/O+VH0v7Sk4T3xNVbZoBPPxcmx5KN2dbmz5zzHoAOjXUhiEmdBVCjW
tq/q1SEBmOFb6PAFraTYgFtuf1aolp6+hr7XFq8R895vUxfm7DY4t6K6hr4NbpFvW35jC+bBJJRd
WO53FEZtAQ4Mddi3AcLhvE97/vStLbb9Hg4kBUlBRGlbPCoIJ8a6GxtwVjeONKNW6jn4Gb6tEM1H
7raaB1OSHJsoJyaUWQl1C0YPbDUrSddbTjoUl1xFz81MIvvqtjhiLgTzLeqGCWk/E8T7YEU7DP7T
7+LACG7veVo3KbTfY3GuN9jNPaBbG4DlV0J6lfC5aKr6h69FhSzh/L1nU2BI4LbcAyG/hNzUap0M
jgRSAJ+p55xlIVB5wbWEIZrz+iNJ9fNpAVJx2xTp1z7Ko1eba86K1/7aLNeVI3l9KPeIC3qPTZ0G
MtXK1SD5p5xm1xgC59YNor2UD4gQBz/P8sz2h6a1O/EbpNpaQuZEANSTlB2D7TYTyB59TJTaXvQP
MCpMrxxAJDNByAKrT2764B8FyS9LVLE6N4uwTD8mjBQ/5og5pgI4AidMBd3YETQG2JYhkG6yGDO4
mLFSo1LZCdPFnYy3+6Re8lTJzRJwM3nuwOnCUs5s9H4BPeXKNz3hPTFrPbZt1L5NgRlt0VE38l1m
Z8kq1RCNuo2hvWbagiG4m21HnYw2h3pHWpf/qv85Xj0ki0W/viLAXYgAkffHFuLOZCxu3rxStxNs
qi/cpUDte8XFif5eaq28ssXhUBK/9bde8k38SEE0WbGIMaVz4Lq1Zn07N18fp+gtFztHAw5TF57E
kO9oZNxAnsdbcPT8jD00bSyFhibueYo5x7ypg+kaoPhXNbxc2PWk1l9RGgbgrVkWjfSnxRXQ8Ecq
+FQF8wJ2D+17BZ2qE1skn5yca5gYMIBVXc98TyJFOEOwqi4PUXX1mfIPQs3EVTfhEXP+t0fXGULd
RHcch32LcxpZfLzpFatCQTKbSBp4efq9ShBkshsMooSgdPPov1QEgD9uMlho8ir38VZZa3jKO/Jm
t73fO9swnAIClICaI5WwF7jJod0o3H2ndarhxRIuKV4U5BjzUOghIPcr6232Nei4zWpRzLlKYhY0
ekf8aaX014KKNTJ/V1fWbBe2iWZL/AfL5XqvM/v+yZy9GJsfrOijOs0lozItmhtAEQcXtHjHhs39
khclvYsLdGkCNbREnRxWUvEaGjh7yShACG+R6evZaHQg20taedva3SKfs86tN3+BOi+30JUWkJsh
3ywSg9khEBiYbMBxiaL9krMLkB9eS1M48nlaWfccHyOvgZhLnUfahEc5ARMz2X4y8+hJAowsh7Lf
W8VWU24/KJDQ6RWGo+bYC+gZVMec/We2bgpZLAko3HCBYfiiHHz2duPT+3XeKw5uwfmFOCw6IFjq
bEyvREK33Q8r6FWWSpWG5f3JwegFVhgMINyxPi9mJMxxsKTInSpUTAbOxdHerGv5w/aMIx2y1vGe
UF2Ik1cLH/6r8J3nCDN4AR/VpuJR8bqKqNT7oibuo2dHCXzkf6t/nGZo/MKbg1yRV/jB8wQf79OO
xo32uJ52k0lQ1d3Vst1swg2JCHyrOhnL3/qSSk+WVz97LFCSU7NXASAZ69OcWxJ9jKbPZi1abY4Q
o86HXTzpLxfELcxMsApajWDEMKawuewkdOwPi+0/d7X21DKD9h1oNcs1qeXN/gWVmatSFzJEAPyh
w4NG9qVU9dRsESjgGDHXDNnUBLsr3SgzT5w1uEbCUOVqXnEjOWt9anVviRx0HHEv6R5GmXVhpLLG
ExoNBX3njgjKXMzoYWc1S6OVP/kuweHdKpcVIoji/nTpRCqe3uEXCVjvSvndRaT05GhuufTZ7v2O
h67CdtD1r2ORF6xdnSXfa1fOKHlpGpsswwVVbTucyCOuv9AZh5dIBLE4UekqZTmWmy9iEHULj7jn
1FveA3t8jIsPCmHJeI/aKsP8kcuRA6MGOXOgoX87RBN3rJdiEWduvlhc0dIqTkO51tQ7aisx/Qpy
kV42tkiz0seXrMQzCpyWqDAV59mPGqPAOqMTpDsN64cVZMVwjs5FE+MlzNHXAicd/3FhNXD10XYZ
ywZ3uVtqZ20wjydFf6VnVS3m1sZX9ug6jhfPgEZ6RImE+nfYbE0iXaAc5RGrEnAjV7kNe/8TYahl
zZKoZt3FBVVFfC0kP5iPt8IozDbBBSwIx6HK2u809VM0+RfDrag+twJgD/baQUHBo1rpl/+43sL6
FNntGsnpV3BmTYeX6NoLN6fuCnnz5Q46XNNvnlb5dy0NwVd3u1jrqCJW4l4FXFAN46yeTfm0CLm1
Fjd23UBchHC1uXFQy8/ilbH5wfJ/FAm77kvATw/kpSFfxBNWwkUIO5QBzUqiz0NSZ12BfyYu3B2w
P2/yZ4ZwUMhm/rYQqUqksZPGpkal2ax8BHZQPSUwh643WsqIPu+S6xcRn2tTEyoNd2Vc7sZdzzRJ
dbnl677ffTsenFK/HPefxerX9ruyJDOgKgjir45Vw7xYO32hXENSlHQeHld/3wBrfOJExVmt0VW8
SENufmaVUa6xBgEIaLBqp+Kg7R3nmazKkw8Db7VH/m0tamS6ENffYCO5sB+tZxFrm3QZS3qR0+3v
i88MoXyOAlBB8sFxMf0sP9QtH3T5M1D/BO+7Y0hEzmGRr0ZRNyI6IPUfoaQbFDNQxtJi7Knzqaea
wG61nVZ1puvqUI6hPkiJYiUq4Pkf81jwVwRYeJZRysikJU4JV7c/EBrAHd/gcmVSf0Btx7Fj0Ktp
zwcjI0Naw5j+bGSkf6PfaRai7XfeYf/uK917O6Es5ycZK+WOq1QLKZarpQ+mMnvhesQrfNGchplT
9E48mHPkHR4DiZyt0bEbcgKZcN0J7psgEdGdMkrKCa2vRW8lTHxsUv1ljoSuYqmBaPU1NiHgrWKu
WdQRE0D2d6JinI67J08b3bWKVxsl8N6EmGkCV3rtZN7QOZDTyZgkuo7SncEKFoQB7jMkhBSxhU9m
Fs10ajThI8gQXV6Gxu2zz6DN9Hwac4JD71LYZvgvipRLUSDjKLbLyD1CeNW6m1FFf3jNnrcEabwG
brl1BQV/FFHAPBoofioyvWdpLT9QR0YhlZaUVXwAacEhi43VqNIcYtyG+PePAW+LIziW0MZM7uee
i7c+jIPPVvto4LY8RqRMowTqJqOXlq6QMAcQsaeArQR0y9zVX0QO4vMrPUWJQVCu3xO7dJUg8Rsz
UT8VMDad11h0stTh9WrqZ2MY4ND+9v9s2IxmhkxiNVffCHsCtZFp6Lm5wRIlXzPlryhhevh13eLW
k6a4QmCIw5ljVLloR22HyOXWO8d5/+y5BaZYQ1xueA7iEdYCVZQJLHw1VZXLAVvWf2DuxxCg9gel
Qb6KTApBqZXQ0qnMLBzChVMpjjo79g93NFR0+0trztSzccZZZrvF2tifMon+4csSfQ8OhCH1uI7x
TqLqLbduoqF/pV9sdpCFZdqyjEJe2XtkmtgTA3oujhWYHKdCI2soHMnidN9LFFFFWmtSvVrx3OuT
zAeHcMEJFDh1266Yz51aT5W+gRyzI0mLC4GfuLKfmAxpompOkqMPM1Qk46auL3zZc8UAaseeyWpy
OzeVsOAxuyh5hRMZYEIh4ZT/HyrM4/oX+PnLniRbIQWNQyeSQGaKPu1T1gMdMeDenN3gTQB/ysv5
LlAI/EDzV7aoI/1tF99nHQO7RNtRXt7nbyQj1soOkSJbj6awjnzbxRHoJPNfec+EKSY/SXWgc4P2
9ZCGbKQopYtIgwmIeWlEx68XZ6fmW0pgJ4QILQ/L7bY0FSAMpIIj0avLsqOq6Ge3NIfm38tLN9ML
3RIAbaXHqo/P/SPto2kaQCVhTi/S6R9cWwaembGqtgffBgwUAHC4IM/6FODbQ16i9qllGM+qOykw
Pr1n8t5/55rwd9whytZ05Fl3V9mWifAMA18W28HBz03YhriK8wWZW1nXyqMUH9Hep+T0qKBnxiIc
0vSnqzp/064bZgea5OFfk5paOmnNxf5B3uT/SKEkCmjYQ3OeiV5vUONVYOHz8ir8gMKu4CTcDU8v
4dp3l+mspDgAdbZaaxGqTVaBYtR6MMen2YBYy5Xu8z0i9JXoFTNFIBgsdauknwjcUlKSLSLIhP1z
cBP09XTeq6Czf0ck+vu2CxmowgiXloqOy4s4mfWELHQSDQKtYCe9b0d3k0GHwAGnt3SujSqFfP/g
pOFWOvRoXZjdazXCfogkmCSkcS47Ls/MYGkVYzNBPqB1afjuz+QWRlLAgwimd2xRYun2/x5sqGA+
9YBx7FgOL15ozpYXH7Akuz7d0c65KyLlo1KisaBNZWsy4rcNo+NDlrQjWTm0i8VEP+Yix5qsF9S5
qvtuBffPuVluatsiTPnWFJsQJ/1SqBwzvx92p3vrARgnD/T22y1XkX7VbWLR/06nnPjh0qSw+79S
SKeTSBeFN4mo3oijH06ljavHrIBwZybbbizzbfKN7LwGu2kep1Lg11oTqNLiDViKRTKN4AXibtuq
ysCf54vKtH5KbeE38UPCV7aeYxakO9OfB/GX6wuDWknAg0gZY3CNIaHKB/1/9HHMdnIzdQPA7vTq
cVPZAOH2UhwuPLLg2CUbVKeWWvxiK8abwqh/RzVvobEQz65vesvNn+tcVwH41hpX8BRscNjdF0hj
tW7zVU5BgsXGbzAmxG3+50WwCrPlO7abU5dvZQoO6+0Fbhl430KniVC8bzLdwBMsz6L2eCPBD/Ra
1PoXbAMpphOaas91gXNokOtHyd3GWA5zbiPvMZ32aEYEPoUEjNR9+NPA4DWrEiGUrz1PgtdlwVRc
hPYPewj1vsuXbUmf1vHY/PFlLciMfmmVNDj9YdhewtnWNEyR1Kh3zQtAMAdRfL/iemPjpEuFKobe
aOo/2l7YvGHcXZE9Tpe5o4QL4Hu5Pbc/47PbGAkQ3BAgvEIUvG5VvnRz6BXhaLTw/sqzUQYxlxQa
lFSNMbJKHyb/tI2JQrx1k8pAwV7bupFTaY3macLLewQ+sZKcAw1Dn9rW7tNV5ZRoqKT3fYB83UPv
dWZb3+PqTYZivlKInmqkpwGKesi1tfH7LaXiaXyVORSKIoDi/PCSV9oUuJsRw6oFKEe0ghbdlqHM
ojkLaAh3d1mtZoAFBNgh4cOAxBcg473tfeaRYZY/62lRot+p6XzMQLrdAWIMFeMOPjgf5GTVz8U3
AExsSWTynA+9yIWaQyklNGom3A+ZCeypUU42kaIq4XlpT2SQRFKNwZkUaee+YGZXNRghkt2R+Nu/
qguVD/lBc0iZ79FFuO+OYZZZEZW66nDGjcE/+5gJzNo21QBbXCU8Rbwe9L1RcEzhEN1FSi9Ru5hd
Zyd0xAFIf7Yhlc0UoM78EWeY/VSJB4MG3BWgTr7Uu1+DYXp7qIzJu/iaGylDsES4/EERv1UUL/ny
hXYtChSyi9oQpFoeASM7sIFD6ewoI4jn7YffM7iQF5HpGpt98uK0rAle6IvlyknJaDtIg2SQ6uRj
E++08SYN9lcuetIgVebRwUKU44lL0LHLZAWVvNXOzwj8rrpzDqGjDctc8u2dujM8CFDbbzEzPuef
emGySeGVTadPVFttBOxwtsLdPMVMd1+JF/Dx2RlA6GFHAS2GwMJzR3ztxL6sId+01fhB6iZJ36f/
Z1vJech0NXDkR1vfvpYd3+biInCpW6oEaaVkWGd01SNZwF0KtFxuFpBOHJnIH9YXvYffX0Bv8v3W
vgcua7R8vMrfj9cev+kDRyosvr16B1yN+GnADIvZ9upmDufTS7gM+S0qJAWiFdjrUiGAWI+jjinM
K2GJYp4Gnw7hRLsuJ9+8zGjmt9ekG2/Rz8zAfd92lQ4F+zLpU7SvFpjGiF+gYL20QG/BiBvfbJRp
7GHilgPDJfS6nQA1yRYdMZinfB6aRHRhVnok6KcM5Law5Teea2TGjQw5YxGBsgW4ACjlWqR7liZt
dHYscAqZihBLqMEi3ZCitjJKf86kzZrOSoD0YFTw00nRm2FI3a8N2gLo9wJL8KpEThv7AUNL4rgf
Us2EASnkZMGs6o885qwExh86KJLFn0mToMQcySZeX/odC3vQv6k4GMsIp3cQYexlAM2veDmWz5hT
Kqk5DgJXcr6dtHWEfC1wJeLR5M4Do23htWLGEM9VJWzLZJl3iSvCekBBwD1DSTz0qZE1xn5RtRKA
MczBCUCp3/wybLKQ1DW9gY6KJdHeCKYzuP6Le6hryxsdDANxR5QhANwa3hg8yNgbvEObXvp0oUY9
jpdPN8vu/D8dQRXsTZCydDi/+vP4ryOLVFeKj3qCvSOHloVmGnWLrCi7dbQSWOiWoRs8B+HKplH+
/vJ7Yb0Yo0qbkDHYGGL+5E46U8BSZr2z7XXngwRrzo15o/0xrnpT/jmG+fHxkX7rzZzYkeS827dZ
jMFI4NU3zpHlxou6Qma0WYI3O1rx9aWx8KoQeyggQwQWQUNpyKvX0jADyL1H1dfp6/Yv+eEnv/hz
F1iWBDb2UhjopmMCFf6+NEu90hIxYpbGI7pPR2a/Wp3/9HrG37Dy4wuBpLyerZkTrlmDO9FoLQpz
ycXQfiUFidVZjAcw4TkX1Vx1RFztbtkcTbYp0h7SFmA7CxtHgKUGKwCP/7SSFJuslwtZDYxKCRaQ
i5vlf2nLfhU8siJmhlyRZuvheRrhVNcXNf9v/agziW0F8p0XllxRiaU6Wzlp6fUijUoUUtx28tbm
/V6V8UqAdQeZ2GTDEk10TBuAw/xlVBNgHGyl/UCkBO2SsR5ZqTLyc4hhF84Kk+lXr904+/ygUbDu
ylbvAqWDcACYMUeavX5J0ZWvHxeFSBxuSPR1Pfga/yYZzZu2u6yLr9DW5xFcoT9YSSeAT32KXHu4
T+jKJy0DSd7ZEQVkIbbW4sM5Xa6JOqxwJnUzadFM4bn4IjZMDPsdVB/JfnKj4qsjfGu/7h8ZZY0U
2mX5KTMqdkiTna8apV9145+JzNQ2mCNBibqeJMSAEYseRuczz7BhHondRutrGzEUf45muurNUXqj
wsrznQoJ87NW1S+0xN43FNvZLs4ZTu66QS40kCS8Qsdmbwekg+HPg6Se3lj9er+/a7Et0n5ob72/
nxEEJNX3NAmRK4T/z39EbrNtbDHKwPcs3SQGjikFCnN/NYs0doaDg2+itYM5i0VobUqeIc6dE5IS
NS0Er6ywqdzVetzPKjmpk4sm1jpriEWHVw8K4raK4bal0NfSfRLSbXmM6xPi/+Rt33FzwxAqyxdR
5VJI6AOw2iALjTMRnvOZ68of+jnDObgp/+Pl9H9yhGEHF1ZwYAmsU2EF73zC5io/9EflGkAvkiVX
oNW7Xbzpp2y85oh3xm177+NYvpYss2sL7Sn4p46xy9WukR4D/EFlScg3YsLJBT+ByUspcaOTnTAH
SU7S2NqHC1KetdFWlPyWfeYZ8l9B5BxxzPWZ3TXA6EHsPyC5rqgzaC1GlCQzJbfhCk3wXH7t02ND
vr5EneIJlNDYcuIodXeVJs2mrAuWEDeCyHvdPozyHDMH1tdLJHxs6XxA7PPo8cNy09U1f0xWk7hZ
fhaCjSuJ/YsiGm7hoUSzNe8KrHjcuLegP90IjWWkwP4cTT24WyN9yv1JMmcJXFiOZagYiqxC2U2B
DY315YyiuuHV+lVbR2SKAzzKt68bgxcJU6e5PTcYj6S4thbVwvCZ02RtCr/Af5PLGxhN6C8PuAkY
qzL1+bKLWOIT5IPozIbSo7OUbkVkvwmOKNVAZVQa+GatdubHy/OsUKf29AJsqw/gwoLA9HPbpB+D
uHbTkuYkVKDmof1Q+ULPRG3ctXj2aWZIAdDdW6rNvJXQtNKr02zXdQvHUIhh/hZv8mdq13tLRRBW
nWU6gkrY+GgNyNj2OIkUs7g/a2SSmgN8gjwSSwOqpIQP9RzcZxHzceclLPEhGULwPKR1wkYAYng7
IMAGrtXnpLY+09y+HorKO4kCy03jzLPuMkUxB2C4t5IMlZjMPtlvJ+Dl0tuFWtCpLCel/v1OAjLp
EPMQz6JI+ZO4DAInGLnqWrDPst5UYIwWz5PL+3VxOfrLrROVDsY6Ae9f7RZAvhM0Z6CFhDLbX7F3
4ZRKM7Mui9aGtqZb06zKwe77rzg507W+sn9VOyb9W20Hdm3mEIfsl6O7F/+tK5IqWLaYhMHJTguk
ypJQdHH1GMbVz9G5IyaKFXOoupvQ7ofPCNmHyL4CVAefvjieA1K10ygSQTMGQxhKxfF2GwO9aoLD
Q+/ePFgSEWiZxZJGPFharFsB8Hr41y80UnsDcKf5UaYqnShbyNSfRDKviwCOqUzfxrVVrTkYAuMu
Bc24ctY+ONsosYiexdDLoq97PHTW8YOyoMi2Oj+2MGQm7ce9bBoJsN3NfsafASA28wpo64LKwzm8
9Ktf6n43iq2CTJnW+AhtkbE7dnQen3WyqIhP8NmmeUBYg2HVGIwJJ1UQgkTndJcZD7k0kT9oDy+E
kIiSQ+o/h5UlK1fKU2XBNS/5kByzigG6Y5K3Iiw2Z6vg76Rh2wsO0cXY7PTbbHUnQT0e7dGwZ4eO
fCiXf2P7OpHR20dZ0fm/GDj0krmSruVlZwtkV6FwixnGFG4V8Xb/EjhC0Eq4RC4Tfsf/3rQjzA2Z
IdsqMtmB01ceZTbDQUfW13X1aBF00uVT5QaoMhcAiv0RUmfn/mJAEczHw9ZaBwd/BjlUCB/4Ljnf
d456TNWzzvUc4KU+m2AE+3ulKE6cONVSBMiqJMNPvO16YrGVNF2siOvIfC/YW2e9YtoaCgjVkEhg
I9tFojsFiz2vtkjLN/RYDRzn9Xvo0OnCd00XmtX7YGlBjzvknTJ4VUaV8KUiFMj/gPdNpG900sGg
BvH8bLNYsHLAJkdfBmpy+LZ/TliuFQM1ui/m/JLxQ/OArR5lAURXCRdI+ER1UUg6bzDbDERkjstO
Kb3D0hKjeKwpVGd2sEUwjsFwan/N0lf7oo6XA+gYWbwguODgZwz2Uzt4P2Ni+zgupLKCf90dHsjq
pquyvbDf5tO0dGSDtbFA3G/NGmBgC/QNtFpLOoVEgkMsGl8AEU3QOHYztXTCB2EX4SWg3Y9Qj3Y3
hawBHAnoWnkwfLUf486MrgZOYcyRIvcG9m2ib7I5eZyv5YD0xe+PQUYDo5jtwawRuFiwlLqcfB0t
0CWkJHNuCLbLXnVATmavfI1YKuUGy54wjvkI3deHDSfpScrRvC14SZ6B8Ua18112lm8ugduGKmaA
vIOKizSpaQS25UisDajxoFoElny6FBegxml7b/3Ekr3D+0KJfunB2ipPyN3riyj2I6jpaIQLBKNb
UOVSzJpdIB49kKZpl88F+CbHqnrgIZkH7L/I+qfL3qK0+jOX9dHohiTVQUsIsGw5s+caXO2Oik/X
ydbDVKooHJ1GggmrMrnVVx5H20SIDt5gXMje8XQWnsA8KVjy4a1uUSPC2fqmKzEGhHe6IhFxAVlU
dS063SN+O+El1iHOTs99GLOjAYm3R0g39YNadPFZzOTb8xXJmR0Rh+2tCMr2+P3MY2RzSIzbD/80
flyWTEZGKyBwGpPc5j8zDVS5M1jMQd3wHsKqzUh5fBYwJw7W8oUffgKVZ8YS1CZsT02eEPz8zAP8
J6bQ5AMSkRugyGguVDuSRLsq4X3wT8qztXUPTpB1T2OHOgsYOI4zPD0DDBmgP/L5zcslDoP9wpVf
PabQf0JK7/mIijCYZcGAfM8TeveyPfRT1+Iku94nP5nwwVM3rfEu04HA3Ct0DHO/HcNGR9c6kSrw
fKOxlTsnwV84kD41gWWgkG5r+0x1+wkcsUhiCYjmYeho23B9pufDrDBlPBlhaWMzDvO98d9XphVS
Pg5VxB49NAOUDM5+oEXIBR1tGOjuKcVnRzRmm7AzGb5FefZcbjGOYla5OHSpCpmqDXH2J40YD7HA
vKsiWlLDCvowvJq+IUOBeS7icouJoJfK2WWpfGybRBmuev6u9R46drVYTJY/8i5TaMNlLfNy3hIn
y0NGwSwxAHOAWAW6uWqw1Izk3aKjl/htj2DeLNsWv+e4kDUMcHeMkCm0GKMcRqEDupmghBO5X6tu
4Re1PtXpMwVAK5+ePV5yFxZQGlARukbaQw208NNuxA/VpaeVZlBLiVaVdNW+Unigt2Tc6NSs+N5h
RrBTgX6Rv+6r5F54A0G7G97ZPU2+KN+ZU1yzk74PUtJHHOoJEhq8D1NOvAVaBNw7IFk4AqpPk/7m
N4R6Gmc1v3zss0b9fCiAbI3t3ool9BELN4o1VaCQMTeWlP738Gc33KMxKODOPayGi/dHpl01OcKK
gcLFif2CBkU6EjpyU/5QhxEAYBGGtFcDJTacDLNhhE4KS4ixv1qd5cYJTWPjsWVF+R2veBah/ZYH
9yp1GGB/uHCykjt0qHGsJNVbm2WXp+0Z2sAYprkJ+xk0IgPbTgHh1cIKI9Tbfsw2aHm6zHEXxM1I
kuDSh5DIlC1e5SPVLaDSKxVvsqHjxLBaSI2s5QYdtFgCBf25+VBfZdCy2x2TwveXlRXlik/M9AJ2
iFF++TFxbWQVG88RfOlNePSKSdLDqX5AaHi8uzM19ajK/8nqw6/TUBFpWlHYyBS9yfOS9+uDVN5O
FrJAlm7bqBzwfxQxFnCEUraDXI5se+5qM3vvIEcI55krcXvfcWziHTQqPDMN8GoH31aFbrxONOw1
RN4fodbxKR5e2sHnxIs6AnC6lVdlMWQ7g78VysYDgQ1bL4jhZbn1HyiTNGZqzXErLDw3/ydcrDdz
1cjsFgM6Fi4t9hcWXfDWDbkWFqBVm9pDM9LP/Kql4+lPSGStYUJH/qanyH31tFg8Rng10VIAXMQj
ZCuq3qUTbbp4A2tev7psT2Pwi8C7NCHLLE00/HNWuMX+7MZ70EF5eDpF8VxbF3x8HNSoFKyx0EME
umejaNRnM40GsOa1w5JhYBgIi66fre8OO4n8qiAh6Vuig8YZ8tMhdK/uGNjzDQoupr8AwTnb2LP3
wMJQ/piCTz4siQNTn/W7eMI0M41pgn9Amw8PJvqHJYiUlS5z0qxP02JmM2JHQKsqDLM2+XXOfroj
SwAPsuibaFuMHTsmAPbNbUJiHmZRYZGZrLey23E3to3JsW0qaqnzLAXPT0UVvtJh+Mt2nL5SDW1j
k3JXXPo2ds+Ug2czUs3yIwIU927TZwMY3aeEE8D4ZKEf1UqmN+YA38kEJayjVostGRyfkIxw5wht
jRRAeS2upCQAMOWeiH2a3bJahnZpVMM1HAzo06/tlfc0WPk6pau7TQ4Y6NHEqvvp7h4lcIqLQ1fA
K9Ggt2HYYIvaLzyBHNCn624c595HS9sO1pIbx+NWJW4vyaejS1acE2uor/FL8VbV05IDLYHhgh/b
FtrdSYXv25iO8rxoKHOm6uVHeFNjw3GrOsHXUF6wvNnn1LZt8//aBjdr+IWq87h4dviXhjntLyvZ
rMNu/rKFH8elMMZSBsOLRh8wpfRyWzpRMQozXktpQszrzPcldkVgHTq5EjC9yUsoPBY3JjBxBAV/
haRW9cDW2WWpF6CQhUmHI6WjW2Uj1XA/HfH1nh8460VXjBwbk7WNyG0H9Mx45k9MDnumYTmQBjDH
Gj2xWBIZiplInI2RSoGqseIJpDqYrWPaGADZSB2eatCyxpKwTvP58w8/hSXviKgp8Eici0eYzdTm
DwrGooBx8WzIy5RZNwzBBpNbueFHMApy8d9/UmpmJ7ZygFSSmhlWyl4Bsk47zbAWyVSFC8o6MfTT
NRS2D/zyG+OCSO0XjB2Nm/IGR2Ne8RSUxN7gti1O7/d1FkeB7T9jxqAlccxkfKgDPatosyGKuJpY
ibS/N0S5j+hRm08slYxqI7BsFJbcdAVDgQQDp5tx/2ZJp6hbbZLHRStaks4I4j5LfsCKcvp9F0uC
Z7aP5dTjC9VZX7PTB67fyUFFJydwPNLvRlswBL1Uwfh537Ve0/PLYELJFcpRoZ5wPDPHJ7DKWh0o
o1InZQIV9rfqNos34aV+9LFDp6dvE9S6hRKyHaY5Oxe193uikIa69sugZvpsl2+w+qbwYqN3NJVk
4lK2CPFSEc1qIyzsf+3nrcr+2RsXz9Un6kxB9bk3cM0/YGOz9bGN+3BEA+ZQTQ6YtaO4C3NE4dfs
yhs3bL2NIcOIbTSncQyMY7LWK0zRDaFkbjyiQjhdT09Yll8i1g3Xtxa+MWeIGuwV5E3w6dfhGKcX
G2hvtETu5vZNMt6LKJhJp38Aii3NufrxDis7llPnU+QSF3DKzh6zf1qNFJUhQb0bWvlWLrH/YbRu
Vg8QsQ0bsGvKgcIZKgWuhk6vBC64wLygYaG8/VL3WwDqjyMhgzS/DLhoIEE9P4+9kZ0+SlhsYFtU
77GhoCg38EI18hefAadpCOeKajElfCcw1yYYqYY+f2SIyfM079O73439QD3JGykH7+MfDVk+YtSQ
rB3k9ZA9Y44ezrS64dhJiQtA37OWgVLdPBVTgM2m2adTDbI3V5F6g7XfAWDUVIfy0a1i3UReWgTu
QwbpBgwt2ZhoYjKtO5ADiPOBccTLbxwP30wagLlBxocHmk7YAlUUQE2T3hVLEMdLgvWy/pdDjzxL
VYFrF4GUYREFtI0R659qAWU/i6By40syvqMgOeK27ogaWW5KqWHn2L0Nn4mg4JS+SCuPGxdYtF5I
zWpiHG8ZrEaViLw4UrzmnFH3CuMuwpUUQXZep8TiKIbrjGowjv/j7RXS7vkJqfpin3fcD0DoLNmr
K83euur/ZVYXZFS4g/tWeRKdNEscGtWl4LW+/yMjnkLghFxx3C6+dnYFgBDbPw+jaBIQgqlLyy5I
evJ481vpFiHh4ysB82EykYAxr9U9fSUJAVZWAGM8EYHi74SpcUJ3MhZEVRe3BynnEM9bSaYTManT
MT/dcJ3eizoYdljtMn9JwwKWpjpWP2FMfonWKpXHxoDy/YvnEshlHJJRfW9+vfk/po0Jm/+HhExu
2KN904/AaZ69CS7uT1rjM9U2y0Kr1SxANoqLd45wAUE83ye8W+jYX/1WwN1TCdiMsu/xM7jzX3ru
Um1cTywwGNJshyXWJguIt1PI+sd1VRdIanIPKNrM1cSmPvHtMsvvw+NjX0oE9rSpiPxAevMsRZYX
57zTpiOm4qHzm3+kwk+zPLb2ADiT+posaXTcIWpXIyozOvJ+luY6LYlUJEtIqtC6riiLbuLzwBth
C9sPRxQOQe2bTeZneCui3d3wjsJ5SXKdhIGTOxyDqHopbbf+jizDAq2nBrj0aFaV5t2WB5LiV9CF
hcwDtpmPZtlNLaT8RMMk1Iue52rAwjymOOwhGQs+FraY3qTXr+scGpWZdA6mhkbJnbG+Uj0lS9uC
ZFZbZJwtelR5tgE/TJ8YO1kjygUXLfvxrhJFZVISUZUizmZwlAqlmjG7j2ZT86CBrvAcrl4SVZCq
+9qs+NrrGGMYW+aQQzXO7dAU44ygLYHF8TE3qAsDfyFKXTqXn2Gdx3J0/0Mwj9UhrykCKu1O3OCC
FIg+RgLNp5OxF19jBAOSIrOmv2HJjeAiE17w2SuW3kw0qxbqM5SAmARqeZx3xspOGBBDkCLPUxDJ
BMnCTwMBYvZfC337BpT1082n2TqDPwZp1/zb4h+MO/arlnDwDydhOPZBY+fch8vcTK1anQBERvrR
Q6hEgPLBaO75+JuWZ2tAZfvdIQgCaAjfth0+VpFVx/If5pdKuilmTDCW/nFdTe6i0mJQKuHUck5W
HBKQBK9L7xhybuTArVm6LInhRwsR9Urxz2ujOboBA0isjEZA6Oa2kctZM9EPdIwMTF8pMWXRn7oQ
nAfCqs8K7WSlkCmiYrcmTvOvXB/euMCyLJgPkZO3xrhYUa2zIkwAUWJpVeiAzm5+RYvGBmijuGWt
cm62VX032aQAsxnP5dhVIxGJI2ZL7jIRNAyTITh32Bmc7Mt2D51j0f4nMpnj0GedKUDjiMuk/ZG/
Nh9rXVUlled3J+4taR1YKJmV/yXnAVpEncJnWP7C0EQvv8A8kxoOdG2NUtB7gb9E/mwzNf3NmxFc
eeNA2Pwv63iBuQ4WSaBhPJZDLKbGYG40adWgGClWIN/idmp5E4pcB9QQTsh3yVCj1FyAREp47zy6
AfEGIfkh4ned/yVhR2ckXeQESfp2anuVo+/1XQh2CP2Kv+FAqqCcSFmqvVyb0Hfr3CVYDp+Uo/O0
XFXdhxPJh8I5JOuuo8h7mgZr6QjhdGO8FTCorfRTKz2GrCGiVyQ5m4325fjrM/rOnSg469fZfO/a
+zOIyQZ/oq19nMFtTLL2NZEjO9CN3bzNnv5GbOuq2/AFrDWmFhsyhQ+cyEjcjDOn97T4DMfIl6Rl
Wi+FfnlqjRNN9/5+IeTLjLjfy9rEak7RTxcg3mJUvOB7t/bPlkRdmX2UkwaggQh7HiyPWUqKhzhW
hVY3wVAv1hCyeQ7FfrplWmLBOxZLsLX1P8x+rM5UhF/SLgUembcIGY4DUssoygRaxHvrauO4IMyc
8RVJMujWIsdIIXJ/hWrTXOGXscHADLrl5x+xqZhTfbdGkFWmqn8Ovh6a0OuuRIVyLuIAzfo9RKP6
wwRC+sfO5p0DrY32if0gTMHUjktuhG6uVkVvIfvco1w7xWPs74uoQIAPOR9ACtq2wo1hjZJVMumu
RctOFfjZ3R3FZexKu0Q5crdTTl1+hcXzqlqolggrXTeJqhZktTCjlryEiTGZ4dXlcxnCsvUBJ34h
jBie3OAnSDISuLxKXU24RqFm0kB6/nCHRT1cd9TTxsGOnQAH2nnLablcdEf3C2R4rv/zgwKggzS/
Odo26benAeOe+ACo5O5Q3l0pcGFv9f994644ClsVCks5MtMF69rUeOqycdZ8jR1y2t4+3/zZuMil
ceukWAg8UrTy0FVyrs4CDcte3IEBl51D0aDbqOKdhVtkXS6+c2N77aK4O3AviCmOemRHuwa9QzYY
hoRcyNon0OkWAZk8ssZgK35ye4dX/q9gDd79YRcDmc21S4HXModXMVyz8Z5EBzqGt/3TIO9z8qeM
hTLhpuXhO6nkyHSyTZJW64TFBhm5GAObFhkbHzb0lGoKB/XOci8xMDfnh3tdY5rR6QSe1JsytWIi
QO3c2CA0HEX984LaolZZK9Pc/2/XRQaYL+UlhHPOFLz5qdmHlY4pR4NrksHzEVAVbt6D8NXSis6r
9Z/7FSCAAWDLmDMPGwsgqtTb4viapsuIjnQg6Z7+Alc18sXJe+7aCz59tRQIDq0qWu9n1gitWViJ
uJoR27lUPLBwKXT0OdgBXBTC4tFXOz9KwGi30cPvc0MLU0achxeuPxlCiUojuwN7mC2g2cfPGQuk
WmpQr0dtr/6d8zrfhm9m294i/UuaY45tnvQ/FaX66Su6X4cagPm8/M16TN6fYBe25gz5lMBV7UHP
iH8oONkMpMdki5+EdxD6FInGLsCiNpH3C5HWxyxPH+bKkqsppdloV7SDFvwsCggLQED1qb0ELuzY
dYGrejzim24hR2Sq5ErBziQ+gsgdpALgmg6dYTpYPSdS58wsJHeBesq4VEfhwL+kH8HsliC+R+bj
b3AaWv64bZhbMXhueUULTSP7FqZJQonu1HxNSedhC7qQjs2iPcJDq5xKtKargO39F31lDkcMEA4s
euRqxxgLazZeZYKc3Z0Gt+ecklqIGj7/T73EUDq0yi+AnxMEqj5C6BtGy3mPBgCKW2nfZG10M3pM
3c4mYzpMoXbYtSq0288GV+3lr570eJTEqralEmSTMKV9VD5IttTwlhwY3ha2uka6pyHObRF1tYIF
jQzVeNP9ks3FJkwwx6fJadDt/O5IYO2Z8O/F0mURgIfMUKbtt7xPotTu7lsEndFyc6kYSfQf+yfB
ep9DubqHv4uMrlIhaYwU4nkawQaNV9RqLTfQ8Kc3RtUioGz+ngZy2aE2ZqOpSkUFXYPkaDj+2vqA
Dy1abNGvGDKYKoZe8G2EWLwqKpSTs+TWH8i4mwNn/y7hz6l37C+tfZrTTbRUsNz1nzusdCy2lLC8
bEtEtP+XmHYBSuYraO+jPdpzdtTQxxzff1cK/J2pRC5r6yerNm4ma9lC14WbakhccPfr4ML9O6Nx
e4vtQlcyCETSi30YLfgEMXZBwWd2IOYBxk7UEFu1jhrFbip5uX50bAgIzsL46ald47B8DABbm9WV
8IPZvsi9dCPn7E45P6b1iSRPkdqxLN/8EmZpgTRVwa/7hu2lY0pKEfvN/cPwvzRRualQdcV+fgJS
pJW+qpMQWhSM1DkAHvlK5/AMi+LqLY9xJFt2Ee+Nrb0KYK5ZV4toS1DpdFVmYu6U7jidbqafSiUw
A1a23DCi+CJqu226HBKcgsO5oTP6ZkR76fQoFBV1ctM6r0Yv68rcxdKwKY92O5RX8F2zPhfbS3/f
YQjcNdYlF4/+xzHZhDsMLN7T3BJo+lLANI1RpBZiXrDUPByEq55EEyUOurfK5RoP59vo8HthBiTJ
oLbvBhi2jTDA3wOm+YZBMdb4/AuQ/DfexBzFjOFyK/7/+pibb+sdCkEdL/2Mo8/dsl0HXxOYVYmu
6VXQaKVku+90w+qLndErFtJuxC6CXvs3StwDFFTL6Xt+DKXL0+1XEZCu3k8/g+KGIdsgVHa7TuJi
cAJqn9gPRNOlEbb+UzCstpZgH+g1ylQvNiSBTRz9gXoGIfwxh3CUnyVYwRXMVEs8TRkw//lRaTRR
A13iXeq4+57bRhIQ+At8ATWMPiN8mb6tLjZ2tYf5KGliLW5umSNPhAV50kHg5cC4YAgLeLr1z8m4
EHL7YCuRIyWu7grQMJ/pxUXvhQQVjySJ5QL5D7j+fHCqyCxJM2B7y8eeHmqnZW/ivWXPmq5I5rgN
vhVCVIOhwPQfPfZD/tAujqxQ2tgpGyfhoxTqs9y2plnwHmlmUjgl5kJmXf7N2VbQvk1oRuL0BRMs
2UmB9nuhb396jtQxFrx/XAjbJ7jix1CcUpVBOZxKSwEyy5O8ORAXGwPb2dkx/+Gqczogpn4erI/A
5PPMFk65UtjOtjb78mhL4sut8wuuKMjK0wJgjppl9wDwL4PGjK6rrVoWAhsnrbkIUIKSeQGr9lrr
3U8gJQDqXl70v5Rx0ZMZ8o4n8yWv2WJC9PT86Gntwgnc2qBAEDf33Y0/WBVjE2ilLq6KitaLx3Jo
njp9iNWrnwmfwrQ67MCOMgGs34IATBagW+vdrcV+lC6RH3q+Qe8dv954TvvNNbIOPQzHD9SQRWnV
21ajapcurvVv5e7st/I8DT812lZaeLygajIqciXUj3/Bczivtvz1wi8LHAnbgWZfuHuvDGOqYeVW
x5dc2s2AvNkyBZ7A+EhspnDtiHLa71umsRgZ7+UFAtB4WDqvyBLQzrI0gv8v5kOU6jowQz98NNli
N+Tbt0zu7Xy9Q9b/uYfr0g1Uoq8mAaF4UcoFlAOJC9IeAPZgn9QzKtlIJ8SH/AZBn87G3MWv7dCb
374BbF/PKvjXJMPGB7ry+HGlhonPgg59X8vNkKHXHJiaIK5sZwgfd2FTkl1nDEM1cnJgwuCLBPT5
QWKQEIVMyROwrKvGn0xr8cMyvVV0q6BpW6bLC3Kx/cTfegDMRaSARTwzZck0XMdzC7AVkMmUXpih
m5GOvimhYqpEPfpp+7UdFzk8xF6gQ6hbTqxRmW+1G77lOoYAMhcasLMPLSEkB8wx2gBRoIVZXita
U4IS8rDaZq9hxkpdPVJikoFl5xQkAqhMwiabhf2F+ZHACgLutUqT2o94Hmg29uWmEHc0TWuUTgWv
xQBAyNtsvQlOhoPL3VYMsvDeF2q15H3n/Y3GR865c5K7dLcWqqwnM54r+2781DjqLwRu5o5ach5c
d5LDNwo2Qc/4za4C22uqhNs/Ft0fEATycqi80NDGWRqwLM9ivPTh99LyeoWD7g1qNJaiyJAsmzvl
Mo+1H71nDtOATRVvn22E1aq3Jp362WNHEq8ib3WQ2UUGAjU375VgD7QyNj6zspY+/Uhh6Y4IpLov
bAhq/fVRLaJa//AIIZQBX/2utkD0HOX2ySHt5dLwtdMTZ6JTfxiIAfLOwItpIXLcWPGspTyXmFrq
1Jfugkvp8bJRYzbqc3HSDeXcvZCHFQBnpRNOWN9NcPCaNi0CultXN/IZtXVMWoZ0sLY0DUGe8nSC
d7fsgu8wr/KPEmvH/gjE48fzjdhVM8YnzOvgB3CYqlRSAwCMDqDHGAK8xrdCesaKgK0cuz5c+NEu
EwsMbmUUJDJnXb/IuaqF3A6Wkl/ryuo4n7Nx8/YNLSP8J+RVwUyawjcIP81K78Y6KoBvlomNf7Tl
CuCl//6l4JYtE8VK+kzreoOUgiErrnoMD7RpUei9zaX5bE/05JabrCrZ1fvqSxyuaXY+KoNlb1/G
VdNi+RJe0V2xtukRB9G9e3QquoUH8iiPAwsjeMruZsWvm7W5wt5pKAoXTN1RKVhtbgfzMzBxtnmq
g08g4cCPvlDBqjr8HGXvW+JybqSGW3vOufvLP+K+nx/k5TaZ9FMEzGga4ll9rQUrhC7aNlkkZElT
veyfu5gtUZ8c95gd2zw7JBT9u21dhTknCC935QRFgPJfAcpGcbJzcRL1kHO+OE62grGYZknBxKTS
g6/uIy/9AlqVIa2SIsc2uaFOgh7AksMNfPu1L60jbnAQSUUhoTjqw0uBrz/XU6OO9KVa5RwJfv8y
4g8W1AoR6gMZ4QXIp9gIjrz2zG0aWnJGO83ut+5C0g2xbVaREE/gFfNz39haXEXJG2VOks4G6iYR
XgvlrP9H6lIJ53kQWBXLjtb8UTXRZYdMzzPx7Nmp80QPKy4j4Q4ARC1wfYdj9AUj3xYzfMIUtBQP
tmfnYfMb7SQOSbA2d7oEywe2qC6DJ59rHAhUJQyE3RfiWQ19ZjY+NGBFqYJrqc1s6kUvmKiXOhV/
Raxpn9OVWDFDyKSS5KE2M/s9d79wcNO+i2iIVI1aHCBJqtxlDRSU6CiYHVWJrv8mtd9/OYelnK2Y
DV1ORa/PIh5iPVBO+OQ8zuQSsfLJmbmTGbmRCji8YxCW80J3lyHBMuRN8KuXbq85E/9zMyCcLAOo
podZ0aHzkI9QLPhruVRLyk/JMGnA5aqUyjkI3oJT1GwfkJdU2F3MdCSA4NZ5crhSx0GQmEjTSSN3
3xjCNGuGqW+Atg8jiqiBe9DeRzBMiMfkoMrICS15JGqBNxydaxeTCVD8d3HShSFHS3WxKTdEWe1o
wUag9aCKCVEPlNBW2CVCZEPwnON0U+xAJckZRhGihGDlEWt0Td5ZMq26Hv2aV+zOdJ006qowvGpx
vk92soBv6hNf4ys3tDvsNFzZQRHHUOPez+CfC/GNTOhIN+pXkvRHz1IMSl3s+5/SK02ENnMjOtZv
q5BPiE0TWE5eWzHhzXWooG/v8e/CpXsXIeBpUcK+VPcjK3vUs2GbSA3BpXZSxMLk5JZUeG2EWMcM
5tBbkRhfyb8gutfI9lwLfZ95rxbdXqabFYiPfLZFK+rNuNP4d3FXEuhOtag2vvJGQFwn4ZI5sRZQ
F0bWvsn9mZcO6EoQPPrsYS4iCQRgDRQKq2+UPjF31rGssrYozfRW9R/BqlA+17H1QjkGfOTVKrh0
lB2TsCQPFkwgAuCZCgKVkltl7RawYzSj+V8YCRSsfuce6n/BXYQPxfQXyjvyOptCd6nsMritEPvi
CojZ0mfPFeFKjBSs2vOdJFVIAkTDe+FbdG78NU/9jROL0D2Bm2Wj10KQjF00JuTMyboCf7EtSZXw
VQInpqX9c63bndD3PhHETCTF3RHdRWexSXHHhBnJzTae3KSD9g1hOdTv4s3fUVryQLklIPk/tPIB
dFOY+3W3mCHgmBvPf4iQFSXysjVTuMN78/+1GgR19xvfFDqSbAWQFAJ2UR2QMPYzgpftgFAa3eJl
DWMsclKnZQqr6hEdySkXr6Js48QVthRHe6WGzDmFbiB0b4uORBMFrknqQvsW4HvQ14cYDUmahyfs
QpHMxjZZsUz9mi/1MT0jf3JdVpMyUDclZae6M5NIhbvcF5C1dY9RfhznM5j09rgoQpNJ9ftynn1w
pHyIItmB8mCquRkkpx98mOPPEJSd1GOXpMtiYuvmChHVAQCsPbjZZ8tSQnUHGXHxZFRevmbozZvL
1GjuyUkWh2cNiGpXovYeIqfxuypA1BjPxDa6ytZqkLHIP8tCb6lCzcSZEprVqo6ry3KhT+uYZy5/
s0/igmZoLfJFMRNiW2g5LtiFRTNAheHtbVi7E2evCQMDb9/HnngJBxmnlx7pjMh3AdebQmxvoeMN
kDxROwhb/T49RpaJmXlD9ruM38woaTXLwPbw669uW5meM4GjZQ4qkXW+6JZ4z/FaqTc/D5wD8BU4
2oD4YYYDyaQgvspRRlhGAfqD1Cu0Tq0k0FOjEOupWo8UvEAMQiyho16gbMXi089th0ZR+ucKzT6z
q3NFG3QlPYByLNzuPMfLj/kk8QGxfg1Q0I+1amHcLeXAOlI7VXn1zrIfBPFA1Wz9xnkpWdDHpD2J
9IiP26psXY0j5MIgMJVPEEEWez1eK2gAL9JNRJCueoNxe11mU8jNuYNdRbYQLkWdBAFEv97gIJ7q
Rz5QXFeHC7TW3jzBNOVHWdYPlYn0/JPHeQJLfSTzWFUrThSxzkeeSsfC8hSe47mkIdxSEybqt8wM
kCu7y6uZrx1rAEIVF0bPCdelfBn/OSrP7JPvvsvcMhHMSSqJSLJz7F2r1+jRaKN/4oFGhwXBWZIp
DE2Vx+AGm+qvSzvekpFVngqNGGaGfOMfaEFg/5YA+L4cWMLOWHPn3GfS9d+jHNo56HT/6aHhLFac
GODF3kj4Q7boZhfrVhldHE8HeYMh48DR+wp2P5pg4QvNHtGpUC60BUNbGmTiE0MVAV1x9WLuU3o1
gynOIGIj2hA6GJUsJ4sXPnjg3aSaPvtIcUc1aODlbzbu3p31cFH+MNzxovfUkPbFXO2dqIZd26vm
hHeZhi/le/T5rBq9EMpT7RVXMvengxFSvaca5PiGGxNiYcLaL1qAfPbTbtZkx6c1cQMXQqt7cZrz
5qfLAFZl/dB/6hyhLB2oOYc3f3hkHK3Dm+s7iLUiA8olf0TML+F8F/wwht86V/Nr90Gq8Fva9zuZ
2tB3ATPfX14a1M8neD6iRDQC67wxh2EpAep52CfgWVIOQvBoqfoNedm2AA/q9RRxb85eBabpMjWb
peiUBGANTmzIHnxXd0OzbjnIQAHTOgvcMowWiTKiU6uylp7g8z1lanvbbjK5x50MnIc/hsHlYAWg
DlsW13oSgTLs3ObUlcHm+rv5ya8Wl8aRpDrTgBurgdqvyJ0jyb3uTg8CGU79tNbHoBzBrOzdgL5Y
NG33zkZ34uDHdJBO3X/WugBfKA/YViUZIOV1lZ8sDQSm1Qehvyxj+Gig7StTlSEtxwvhPbLmRar4
5kF8KoPeEwRO4MmD3e0YxSE9y46eh3dDWiO5K43Fdu41MvTyTVyjB29EY+rr/7PyG+dq5ba3RSt8
Ml2Rxb+gS6rZseXSKlR+7DlKZkMECQIgCrqpAs4LpbMUc3kitYBD7wX8s/qWqkbyqjdgXJfBYgUC
GdiL/VV6rwqp7Xkar8em9qBmeJ8afBpuNOy5NwwjAZtexnVO7vmLzeWn/fzc/qlhgmBCMooJ+m4r
+g3MBJBVsPvumVhez4Ot4MBgJxzhQtM4V+63N6D2lcZLNmlqQd/QCMT+8HGd9WeC4urV5WvAhbq0
6v49TS1v7T9cKwLwJ63vS0ZQetmvXvbC32dIy2b/KHlzgcOj8Z7mF6jXyJN2Jls4YyL+ByNL2uHJ
Yspb760Ve5bz4nb+3F9+vCxZH0BJ1cuYzQeb/zfjqSpY4p0RpNu8EI6Ox2qbGaWQA1jhmKCPSzOi
SLAMUHQgWxcbXVQUIQ5KJK1CSyxWS2wnJBPBPJ18hj1uQpjHXIvT/uXr1cPwp6Y8vIaijuYmnHKr
Q56p7vZb/rKk+2zpTbIewp2t+q6QQA5FHltwWR1fy2wUdYSBRS6ZEaLkZNzv6I5vQYLfVjYrfC6W
7GQQ0mcDBZyegMSweSe6rAgW+3eeD3LgUbfEm1Ysd/YZb/j1oDLqBJ0Go/nIfz2mF+mAVNFK4Amq
3AX6P/IBuRioXLBJAO1AQPBHCtb2tWPKbpfBiaowzoTFEq8ql7NKV2cVXWiFnS5cSwy8q3xAf0rX
C0gE+TA5NrbAbF26q6y8C/wNgz/VvwbPuDtfIkzT2oPAmDUZkmvroW+DmsehDinKsd2+3+kLTObT
iTArwY1h9LYMEC1NVZkJ1plhj6VEW8oR0xspnf7lmLH6FpwO6YDjK64t+zG9zdp919jpJMAzDvl4
FWfpkqIECrRdmhyIczCiOvr5Vkmg1SZXJzIRYa7xcEfH1Hm6S2ccMHiZba3ngiO1U56q3DnbvkpW
11pQb1vVHgVoHGgSn50ArPVnlbYKbR/cNZoJYVw8VkzsVMms+EWG4oPO6ENJdGRah3ZBfxWZKHut
WtXiLwcL84WnVuWS6jC3N19y+boNhOBOFTJz3lHdd3ehVGy9Hxq5U0D/y7eLYxzFYU3yaxq4tscd
phX0b73OMRuIyybYj0E1iUx3n2SXon3IuCdPF5O/5/MqJ5/u6TX/kY42raT1z2bKnZWHnL1gmIwW
J96K0yJYlEmkQ4rmPYWkXP3QqPTxIWvQ9neFyHZ9OWRc6IOgtCwbSzQcFM4qL6foqRbpGdtBNijE
ND3dxAJfrIvNjEidoooosntgPs/hEIQpp4g2P4KiMIEJEKHipXbt0NUAVegdKdjkV8lTn4FRqWfZ
iSdPxjIls89pAXZdxQLdXSqEWtaKhk14gESrX2sX8Xrky9yCWFKd0tsxcvKQzFbO6ejklo08g6Xx
njIn/q9Rioek/+X4363ia1fR4V7xZY/09Uh2JuuOHoMc4Z+of2b+6H9QVbkOx6H7m31dxzyY4EHS
LKbd2wHPbNdoXdJLGJD0ULloBFGGH5FDlXac+nF5cm9HYEd/McgcF9FuPH618mXwcPOMuv+AGbpO
hHmcwVyx1PAlVF67eirbBedn8KakH5In0r/Dcsvu6t8WVsT9NntzC6kWza0QvvGKjgHRk8Qsci6w
DHW+v0W/8HdcITbByi8K4AmRXKUu8esdhqxKbr3t7kxOT2LBgABo87/ehgpPqr/JOcLupUxbCPsC
MTWGTHWI7rU76n+jetWg9Nekj670RFb1hPatzvCOG8fzCH5n5fQNBbTLjmqmHnmVTtLYdqcDEJ8y
TSzmTBNvSwt+airuzkC99bmCrcAlxRs2kByxxMnjAqgxbh+KP3KZmMGyQ3UeVowyASzUMElLQyMF
IgjgsjoHY7iP6lV6UIRR3bsHNsPjcoTnOqFTi5KL1tZWdFkncsPyFBw/AkcsgOSVVhK/A3+XugOH
3r3x0rzMlgq+Wet0C0UR13vRM47BdAXYlxnirpcf4pgYY831vmeRXlqj2xJRQoU+jqKdtf7mmF3I
Rof619y6gAZYJHX7XoMzVQkZl7wJdfOyF+DoEu1jP9cGhOG6eFMPoczOQf8rPCkM70rSGKLtjsCk
rm4Ca7rsx1W8liQf5JfNBiswTQmqt4gPwcjO5S/tCP7Wpnnv+lXJe0vqeuUeHpifdb30cGbEa71h
Ka8RAsYtIx+0RSeju+nexNRyI2dRQOCeLwCXyPCcGU6pcJ2UGkRWIbFWmo1NKMufvQwETMC4VzGB
USNbBfJuKi/iBH0JPfNE7Pw/vss8balp95AgdWkOjFO7jz1MmI93E2jFrTpz4m84jKafYpqoONvA
Zq+BF1zUqb21pO8RU0Wkly23OWwgQU41x2Sdw2bhLFbnUH/gRhRWYBuxxh37/51zqsp4UrY4YvsL
C20wkXzQzlRxZTlQsfW/4etImCOj0FPfKYno9N4HvvJHoNIpTSpbG/GBXP4GmNJxDk2qczyvSE5k
cXx336J7QgvemJg0jsTzRL8D+woYOkqwL4Doa8FCY7I+hXU8yLZvnGf/ock+CvtNpsCn2o/quQqO
cS5X+OypeSMDXB/zwTH9BHowEHHzsbDDWqlmKsZ0oa1AjpBdL5pQaAtVej6/XfCkgYSUcYmOYYGj
KT50IG2KwSNZsmyxRNd3OiTSK2BjJjsZ2FpspGMyXa2a3GRMU38FmeNAw0stkaHPgItpqWJywcyO
3od5Sg3ZuFmtJxYaac+njxTutCcEMAHEFRTfr3EokPdaQomw3kKSRIoDJgnpqg2R0M4QFV620Dmo
VprqV37BNKXHs0Mgj0YIM/KG0u3VUkxBps9ugJUe9SRxH4/6LZskNXceil28Bdo8Lx1kagXS6AnS
XlCFQAsJTuAzhXsNTDdej9c5xaCdxskWHiSPwO6rq9w62kPH8D0dLGAsRPdP+ZDT3fesDBQ9609s
7k7xDe6HblleCu9F2rgb/nm7zY/I946XeY5bGjJiDcUHLbVW0DgGGUEX/n10SbLFWxChbTW1EZS1
k5woTx57iPcgVSItTQlEDmUUZldP6XiAG1u3gvYnqyjkYn7yWD9yVubm/xP2Vlo9N2dA0ujDOMuE
8b8hLj3V7AEloDxg7U3zx2ZvPYHfA6NR2vJeE/7aivN1Qe0ZYWrNWTDvlX31HZbxSlswNH2E7Jsl
EoERLWf/8DBXE/fOO/GgGJXTCv0BfyjCnv2M8yyBkl1rmT5PSqh+/NO4z0MOBQbH4LZnFTzls0A9
J7zqTGTlT0dLUuw4b9k6kBfTGuoPJ+GzOrOqHhJiJ7vDLdnsyOHJAsYP9avTeMEym/+4l1ljTNFB
612uukMsRdTeJFcsw6vehTSOkGHqpJXaDpZ9uiFvz8vv6q52vWNPl3LKcl+4U95mbdqnSQd/xrmP
SJ7syvrRGHNOHN25G7AwM1v1aOSjwhqDPhXso8v74c4MftrZe64qfMS58d/ZNxnoOIbfjtkHRRac
cT5gSWPLZp7LbiB2D/BTbHSm9os684T/Ce3B1XfBDtf1ZSKTqzU73Q2o68/4l25RpXPtxb+BKrTr
vGJfabUFlqCr8+7DQWkaUFH765HUzEtpsFVP0/pl8cGCXtclxyiExfJHedOC9jFjv/qI4dN4EsDp
Fx7z4it7SbVEOCm4XEJsj9Mt7CVYrh4sR/mwACJRpYGj014CHOXv2jkeY05jyeGDm6gUaHHwZ0DX
tjsXVMjVPMcDGHcjYlG9cIQEsrF4DTTzoFQ3j8OqhMSzNmMaOprMiMGD+kigum/avMAAP7kcSUEq
RIZ+EuZ1srAdIrrMtxGtq4ErkOn7XdTXBgRdVbNiFLeGu8tpWcbe/pApDYEDYQv5ylXjHCPBZKOO
jlrooBYnm0XoW3PxQqDppK8knQprsQYco+zAyYmERKvJkQEY4/3shckHLt3eb6G8EtV3OedyPq3d
8mW+o3tcEbgS3ZMh8yadh5NsXg69DcuVUlzWPsyYSoNxklQZ0fkSYcVP9FrMIEfoVOrbOl+3k9vt
LynFYAD7QgyCCL1HSixrAix3LmPk3wPuZeVBelYE3OBXu5Z+j0z4SIWpfBu4NBImRwPhq4RSKZxr
dqKgo7Lef/iWrLFlPcYyTtZ3gX+WMxYFkmTBk+HMURGJR8hFhiVUGyZLm8vkkl7b6nEhUBSW+6HZ
fOlYBuM46NRg6tW6zT0wQHrPnvi6vzEi9zXBR0+a4YlC3HoEfHwwxsjgC57a8HajRT2qZRo0kXeA
Jk/mPf5vIYmN6DtEnK1csHMkeG3XDRvYVZfFe1EsTLun5BaZ6If4idMTjBeexKA4muWqf+w/RFKT
3Dsmd9TJzdL7c1n884QcDrQuXOBCftUT4egGgsYjG3AErBrcYGQpFJNAOGtok7I6f5wph5r/aU35
FRjVy5aQPk03jZp9yMLXbiNaRrrv5IRVdM8p/6p66LRV+KdX3aFG3axxToWMfmMVn2y+FV/9v0Ps
n6bbcOkEgkB9UMFQzI90d4QJeIKQmSPMshEjn0dnaJVm2D1nAijKYR/RaaXO7mRMUpJvKw5E/Em1
4OfJsCGSYmqnSkLIJGGL0hL2iuTaJtWGNqRLwV4N99RZMOLBGS0fpv3mxGpVDvXtSE+uMWp9ow5f
+WMu4g+0vg1qWDN1hEKmrOTG5CDJ7BC1orGn1dNjHDI/Gu8xeV7WhJe4noHSNAlK4wLYrnAR7Fe8
UW4e+HYhbuusizviVT0ZmasGDWB6wdWcrG6TzzoLbsf9N8TINq0W8VDXlKXWj9DiVQp+ziEtt+Ti
CqZyyjb636Fb1nYSYtftvqV0s8wlzm+GEEGdhK2Dtpt5W+ZB9qX7ojkwfrPZ9qd1EaVJkbFESeBh
rh3WRQVsE2wUfTNYfp/7FW49C5GGnQGiM7TdSDIK1jn494E6xvU7cqn8CmZ7XaZC8HF7AvmIwkjh
VWC7VF6zv93ObHsPSSzE3eHpdLXreszcTbcgyBCDTrLDz5cw3rOrf0DSyhi/fEtzPOhlKEu2vQ6p
hystRvPPZMs2mqqGDtbS+ivX31xiZv6v0Kngf/4LWahkGaTlyQUklWfGqtpAcp/VCeZtINOFvQ6i
AY+PUaKXu0krGecPbLyFMBZkoidIcJJU9BVfYyyOHnyEGoQPnqf66d16YFa2zKeLtFV0SaDfkEfS
s8aB/EwKuK3muNnTHI9fgmWhij+WPiOiQLXHOy6Qj3sSe802EdRqSOf854q+vC0DTi2E9OnK2j0G
adqI8MqaFPK8SO15CeuakArc+3nF7phbfpBDYm+HER03G/QcxaYkaxHhZ4tjLEm7lEzl6QuqMJk8
p5O8DQwy7TeXkuYL9d8Fx5wFLpDuJH8mWfTIECoxWQAGX2o37Kn1XdfsciAk24vmw8Hj9/H/4J1x
Q9DhBmoYMzxJnEagXWmjvSoX8S5ahl7IAkPYjXiEmB/qoWzO+UOTaPUVkMLuuJ7zHUZIvXIC9W41
TDLdD0mKxBfHpUotYfYLQ84VUEJTLuJqPNtbTWlpMSsP4YkFeyvG9Swz5JIJe9Akxj+kovQseSDR
8/c/bRSmIpiNJLy5G/zMQkXqCeHWrS0jye2qRf9tDWw1wiilE0lf1cXd4MeocKRMV4HZTICi+k2l
53kjVZoXqVpfrS1YmQXnOIB4l69BVtavfzEv0xknX1nBCnNclSIgyAbuumlFsiAcVV/T+buNurxp
Bno31LoOiEJkJHXsbebyX2jXHL9KIHrX+uxpRDnecNdszgxJNXXRmCh+hrRM4AnrLacWqkV79jNc
VaDzbRPjODrx7RrQRY0HU7GM3cSUA45wm/91mp0eit4QGMPOgxAMUCMjOwGTBY7Bw7e5A+SVZ8Eg
ytz62jxo5hDQzKuz1KnSONQYA8oyNL++hATa6SspvNNLKO78LcnqhWK6qKXL52ShJcUbBxn3RYfe
2By7pK9bI23aGFbZ433tyUjoSy8Mdsp/NEpGctP7gfLSd590BIHRlxZA/Wqy7QnjYu/PYBMk41Qw
45cEKqD7yKJ/3eIifEUli2kG3ShGVuyPsdvA94m/5BDu4PFzDIk0IKH/yMksKuDboXigP0gTIPHV
w4+QREFKCMyTJOoGMETDQDfoFZ3vWnL6C1p2VlIULIgsz8ErphG5IhT3LFff9p2lKy+BmQ942G4H
JHLyBeAbC7UoyxpU248JKF4MfGOcI1R3pdYNz3GRh4tm9uDxF6gTk9EPwE3CIDXl9w+kwBQo1kj6
vD0KrDFwR7St6qt9+QX5nuC96FVnpzCn9xO7yseu/jB68wZ0od4rkefOVQvWFBSJXn3nXckWRPXA
9rQtwlLnqLqZ8wBn5bXg1VKaXrhfTUG8Ri9SjePYiDEU7ST2/qiRKy9mXm+fLMJ+7p/ragO78mWZ
gR6ufrzCR87h3TNiZX2N1YeR4hxj23MWdvfQM7riZlc1Is36tz44+FCZwz3cl2ksFOZ4FeO2jhvn
i9BL8ES0axGPdUvuQU+PfdPSmws8hzJZ+0sAM10w3M4xE4v7FUW/eYtTsMidZC0JT7iD5fgS/e5G
O5nD6B3tiIHDlYWOb9i9q9ME9GS/AaJtR24n+mo88FufqT4Ql5+/B5RG5c9fvZ4iFtFOwKjPbqCi
HWcXRqOB2Oj34gu/dCUTCH9i87qMhzywpa/6Uie7IwA6M0LkEI775iq64CrUMUUDnK8VK3YSLyO0
4l/9lFVCkEGjO7rZF78vVh/Jr8pu2i6EB4lbohvzujx++w3yORVaVgV0AG7myXJkc3nTDc8iUfYV
tTCjzJM5I1wnYrivE8+ejuT3PbTFksxLx1ca+VZH90wCnVfTZ6LPKqRMPnY9UfxxGZTaggmLQuvP
XV0o7OIWEl9RLFU/PdpDi/jHWO22xOCkUsUs79g47SfUrukTgJ8+bm3ISxTqsAsIyubYojrQjDq5
sZg+5L/5I11ggxAxdtFQehJ4F/osNLPJx9eQob+xKs8OUYQqCyBdnoDvkr6RgK0aMCn6plCEIcdX
0n2hdsU5sXG6ZVi38rdHoShS5ZpYW5+SplE8m+LJHir4Pe60ibePzAbMTCSn+j4iaQlclaozZ0qM
6yqsgz+K6lwZuHmcOwSuqtf2AGBpQ6YHjFgfP54BRnL50KTd9lL43lixmNSA3a27izmrEIZU0DlA
Qd+gMx5IaFNXn9MzVH4ZiTFZP4fuYU9PwRLyZKu4gAiaMeNnBji7uCvBzXIJRA6AzREaNyDINkmL
VK1G8bAaOdbM8USnJ+o2vyyrPajf6KZbrGyZkyYX8tPSZgxUCfquHHrMCTzra1Va32xUKlhdGx3z
usD2BAcjwoaeoWeb2vv7UzbbDP9ohamjQFj1yfNJrPBuI5t5xJQHPlYDCWijtuH03ULPxLuzS4GV
PQeWzJAr1eP0xkpr/4PiPzkjYsMjphxz6Bn+8ZK7Z7vopnfgov3nywwvMoi07ENxzWUnGL9GnU5Q
I4aWJ+L/vv7rlUivTjAzRjU3u25rAnf5ICKKQiNI1SBDjByHidD7I2GnxPIer6BCLlsp3XxvIs2z
SfcHbL57gD7NJpE9Yn3Dy2OIBPMedeb8Hc/LMJQPfzwT8hXWxMoy5keu9HUqVQ3S4BtG10461FFa
bSfocFVdwTVe9LJbua8GAHJsICtoOB6Yh6eoqAbOh8E3RnYY278MDWGjuA+7zqP3HItfwNFx7gaQ
6a0xpDblvI53VKfKdmMFh1/n2iWSqzDNjUeeaU9v6iPTS3SCKRfyjgczAoL8lsmhqPi4APbu/phG
iBOg78NyL7OkY+RaFaay6LVhmH4AT+XiUZf/iJZarxQPA1+A2m7K+biB1HlOE+zAq5xIrOoPG/kg
hiF+unFpzzZH0HbZldDMB6nDdi7WrI/956uNrikKb/zBnHdsjZosy0dSbp/sSyXaOfi0RkEsLSL5
GurknpFuNNwx7w5DFD4B0UIHZOPlCh8EE43n69G8DQyYVnon7BhNX4DeULc0Kuyc+C4Wb9BhzHKZ
Vx7WuQBSs2+rb0JpMGhsu9gqS7Jhbo2RaQZXz2UHiE9LP8dDA95xJdsKVimWU3Gynjv51p95UfMw
AKjnUpZ58pV+er/J0rPOjS/dgNud0CLStzwpsap8ufMwKEMfQoSmndymVj5o4w3kIDLJ1QDYbdab
Wgf44ECZliXJ2gX1lUMypSDKqonc+oJ6XVMDmMMFaVM7gdb3oSEUJpgfmTAAiqMT9KzFui/21jmb
5dytsoRbVjtRd0BUs+zJo2bf4rQw/0VSK4qwK/cmgwdv8fT+9W8O39JmsgwYIrfd8Z1dyr5EcXaO
tNZKuD8Z8vPwI4id4efzyZhdMDUR+shP56fY3LVcab5vB47fWU6L6DsmXfBwJu2N5KY2KibIiXpy
vR5+Cxs0ntlCtQUVEsDcqYxyJZgJNCMvEcdP9uf5xf6YjL4bmKpGjtrg2zRcr/ae2IABO1Bo7EdE
onePjzokIZDBx6hg6bUxiyMw1fR1RPlyi+N8NoL0URvetip7dO7kdISvBpkVIoOqjIPJFgha1+Ly
5Nmnvdox9+9JtJdLjy1wiXh5ReafLcOH9NfjDxy2PiIMgVKr9sq6h+2eC/pRFqX3IvCC/R2NvhFs
A+hNZHbo5kdb7GXSPHbnlykHOLJmXE9YjbTQdrJTZFrE9p7Rk+IFJfwlvmzoKlnISah9bVuiURzT
oDXsFCgGV3rzfisVZLfy9ovUGdkaR896urI7AgFy/+0bH3l82ezIN/+ajgVg05XlG0mgOa9by0e2
QzMtYQGhNPlVADsukkxmh55UTpJO+DL6V8NE+jb/IzEWK3Plzek9WX7Awm7MyEgNHCbv5O53JZBN
oyGSE3KiDGsFqj3Dh3DJu6Cb9d2iAPls8Zz06EMgYjVUGZ5sDOTsTqkj/H+SSSzem28Mi+ihEqUI
Apm6y5LCthWWv2kNPx5CseFixvZAXKsdK5PCyIwX0pr4jl1xShb75SIk6VkxPLXgFTEwP6n1X311
tr2naXYjKwc30OeV2Z8nOmk42Rj4w3NMhov4Wftn5cKx+oF1m3EB5eu/bd4PSaAYW8C90LcpT0HE
VwUvmrjZE4Tx1o/AVdcMEgwa5Re5LbGufDXcEwxnhbkrTo8pGjXxzMw7M7MfwvQ8e+vLdMStj7NW
1iyfbxZy81TJNZ8sPjbwRl7uYgGkNNzeDw2o6R7UJYjLFlEdA5zJrEjNx5J1SxJ7LrWvQ4WPRf2w
VFX35a23VH5kuB2JPqP0/SK9S+Lc2zj7zkU04gIMjNe9PopIoKW2XwkWpfWWMfnNrsVx/3417tya
vpFL9OP0LoRGsGBnhYt4M2Y/DPSub6zTgqoGNe9GlBMmHatUGYAQz2H84VKwECCWAInSPr2G7vzQ
nXbX1Uut6nMmXK2RG/Y4e5zi51MasoZrorjroqYVBWr0KqQmTFBpTEQDn9zlpQgE0Uex/N6NPUzB
544KWQJ27OTeLY67vOC0b7FnfsAfcj4aJUF4JF9hdsutJXkKso9YAO1kswmv3UTKx3oYv1fLj6lI
HhRJzZkCfJ/LdCX7q4Fo7mtks5/BkIaJbOapCF414ONKIOLIOU2aLibErP0IBJG1lx4rhScyH/5b
3/Bs++/aAa12snTiJ+lsvrrcbvdfdWtMRElTI8TZZHa51xNb8eQniLV0LScj7MYQdaau6tmI1uhm
9XJ/aEgI/QDttiFVK8TDNerbHzVU6oCHzzYwjkTR0VG+TZ0oJWq9WzjoIMtjqkjNjaEiJKkmq3kl
HOiYRXwS1ErryUOEF+s4mv2cPB7NUuOwCCfNBS+wft9EIulEuJ8VxoHGZbUx1H7BmXHOSIVs2s/1
sM4onzW7WsHFdzEz6n8oS/LazGlPUX+yLG1Aa6EtOnUhq1ottau63fEtaPPFUwEInUfwr1L4sI+8
quUXlkWINUF0Zcf+UafZjViqx78PSGzT51v0PI4CywoSarQLInb0nYeEqEjT0FxVcAsHf9NB26Kk
XvQPcqMvYIA6/meEiUp+RHL9GRO6PoA05HhyxTNwYpnhP0ZCTk1Pg5Kw195PcCcQWn5t6S3DAsnB
tgdcLZHd26ZGcp6abzjBv8OSuvSAk4veTVx9xBF4fSgEq9lPXxzSGhaEebe4/VqFSGMvh79nEoHM
5MJTVcPiSYKZWafV2UJcCv+vtoZTXPLfoLRMTfQNmZTvQzuCYaFqEvD3YG0nlhwVnWoxUziHIUi0
duF8/NsM8jqik33uSheFQ2xjT2w9FRPDBTBRhMlygg7OpNy/WVSqYArxlcCaweSKjcE16h4Blhxc
j6KtUmX6TBKv172ZeVRjD1mgGcVsripVzlj64Afr68Uj+g+TJgc39d1T584B2QtW/91YRPbgO01c
QWV95ghuxY5jP/+0HGvUg+1noIcTjrNFfad5Qajpf+oRQArUb5sLf+cCs14j98auim977dQzF+d5
+Qgd+kC34t1cMh6nJBlvQWSEYVMhm8kzjFT7kcyQZPe3CeeK6ohpsLjytobO3bgwCkt2H1XG5rgA
C7snXzxm/f4CjfGA+/d85dOMb3/xbWNX4oRAvXwQ6S+ITR1Y5S5xL+Q1jL1fQ/tCbxQm12lDd+rT
J/JX/e9+dR2u3W/34pliezsDDe/VqVdeUA+jvRYMpolXG8iUCCOvNsp0L7JyVW+lkr2hprqwiCvX
LtiMv7Zeuvs0vzKFVkkwW+F6INq8fQYJBcsurImDq178Q8QHk+6iHI5Kq1gwS+CnGkbyjWcqtis2
aU3MWhGkoM01F7VBcKCHF8F+dw1hY5irSO/WyeGLgeQNK72EkDyFsfFGnTR8h1GzvfseMhrfEHrP
Ox4k9ZIAXOQMtDZmCulX2AO8nQfiC0odKXvtrC8nzLIWbuRH/4bRBLW1IokLQL397oVbSVFzlm82
scGdPBYEJAkQh//AegaBvqoeyC3FwS5th+fw193LKKkQEMgP1VLSSUGoEfos7i5PiDrNyIG9wDkP
o4AcTaGaV97AD4gvOx+R9bmaiqldRU8mnaWAm7SX8e2hH1R+Sl1BgvdzcTE6YeuvhnG4mxqPPjMU
4U6pVfovV5kWqU7E4R6csC+MzJDfq9z53H9oDz0VnJdJtC2vwIHnpazYizIGbcjgNgO/RRLmVded
vI4+2oAEGSSHrR548dKy+9nkLQXdUAKQMEH93bQBfPO68uLiNUE8lsG4dYDvyATsTFnqiN1qLcXN
0Qz74/oDL/Xs7fzyzMc6zcn6Bn96Gnmv3MkrUfIjU9smjhab5iDP+jej0unGJspDjm/Jzipv11m/
A3QI9VMHedNMCx7s1BXD1HLtiO/jvsdqw1+OpTb4rq6Jccpaeng/xTt2YEpIYYR7e3fcvmXcqSgg
6/IsP4/Rcl50OySpPuti1z6CJ2/gesxjmuj68NCbhG8nVgvy9rWsYr8qrQvg3y3Wj48jZQCb8IMK
3wjNmSCcD/btAsRLuMviZaX3Rgw5T75udnhVMKe3ti2kEV+OuiwmpgOQzPVN2jNutypDnfmjHKoW
CBz7hZofLkLuLli6ou9k3rfZclA32hGZU1e4Eujl+RxQyhH+J9QylK+X9+cVytmBnBP8OQluGDkQ
/wIld36Vj1TCURjuBgeKhvk+nNpsjE9TjIi+5K94XVJZ1VAOY7PZ0wl9MF3TRMGsmnxr6WA7PvJ1
t0//ANL8LFDFyp5Cr3rHp4Kvmz4HlYQYtFlzzikxhPjWOklsJMSD+qPdQZLaIVX1tJTbiIscd+49
rHKus6UuE4iYewmBqoCH8G6Ur2OIaHGPEcsuSqOkuEgGe2Qf80yLbiz342/8Jp+t4u6PMWUcqzhT
jdIzYC19Q6qAntrA8vKjiopTjuvlwLJ3GLLrwy3K++t1RtgXH0Jx0B7AsNGksi9+nr4jBJmwG34v
Gv3XX38XJqZgZxnPWYJzc/mhjlOUK6ts7hqAoHzvDsCWsXbRQEqn64i1+LvUfyfG3GcRMPK4hNy+
n7IyjdaaImd40XERnB/bnkUtkB5DOyTtRRr27kD3dgg2LBtcPFF2reRfoc87vBOJjpeMu1RrRR4I
abLYF2p9RUJCZJAZgEVOixttr8954gFfjEmwasaqYk5pqBaA4nRunhF8lIdbrTR1r68FGClhy7hE
ghYHA/fuHn8tRrbooq20F64zBhxhkkUFfgWtnCiB2I/xRPT9xHkn7jjXI+GFkX5NUdK4LHe+vjpu
dYxKABvWu2/hEtxYozA5EAaryH/E4r9D8P1nBSks8B1CL17l3x4T7phiOhznIDRp0WItOv1kmis5
gv7hjfYzMSKtFx/4C22GQSfhmPXs3H2c4UxCLS5ejWAzaTSjqd7EPwcQ+Gf3RzefHQiAZS/1X80O
/S2b0CR12sSsk4551qo9+eU8PdFf8lZsq1P22hXgOhVcOiORCZax5iFN8be7Tjzgw5WUm1k4OqSS
hECYGau3ooP2T14crczr6Pd4KwUfy37IUpIY6yaStzHxxQ2ND9ZhR0GeGc2sZQQsdHpv44ElCoY/
4l56nXEo/NmXnnj4I5ngyqWLLfdZmcsPO2vmiBkPX4nYmK7H9er3Ft2d+MIeqArm0qft2tJ0y19p
Md6csFT9JDTcPGHobj5lpUK/kLqqmePaCf+nsIN1mHkXvoQsxVgTqPhHUAsY3z9f9yOF4WJKarE7
VnMWj/oDdmHlW+0Z+tWljJ3RTScel5D0I4t+8kyzzLtNfPiwcu9IkmHITJ3KcofwD+d5y6Ml02cX
lAMjG2pQh6sVriioOJjNE41WN/ngb1gfRlSG5sIKmdySVHaR/Dcoo62f8d/tbCAAJzspk/vPK/FU
+tXz4PK7VGrhek7STyIn+MY00TjQztwmg4RDKQbAE50085JMGPplhiNCTOSK1764hwGp3Imtc07T
Jt1a6hcseVf6gVNJaaEP4I4W6BCrWsNePjZFhdUC4uRMxOm9HrFiuN+jrkan8+x6AmhKD+7eHk+a
+SHebL3yXptTeY38HqjqUyKBhAns0ZD4kNNOFTkO808+Djpc/r+iu3/0O+1sbjbAC3WfXGFub2tv
3UsiZYpNGz7VCiWbDmtfvwOEfy65NPXTp9B5euo6Iez8PnUzUsJwv/0JrXnwTPn+ejYbh6MC4I2b
zUObKmSox9odvV6h9NmHc7GEbhs5MVAbStblpqicExpnwmEkUq0QJecNiQ64a9dXyTYjwucdO3Pf
R1LzSJqiEScSb89hE/kNQ54u9e+I+rDozDFDFf2W8DBoxKr0B4AvvXE2PB/V6bMDIBJQlCOXaUjj
4DV8XUQPJlQe55RJK1uF5s/P27DV31bHTqfShQnDerJAdghVM68l8McAVhN5F/idO13xwgzlQNvG
bLHmoMUvx6UFslGD5wLvkjRiZGFRvGVS1QSsted926cPDLElxudaHytY7YTP+6JB7GVFoCSqVOaZ
FuEjW5UyZkdINQ8Oop7MGDSwVW1G6bDxZL6kdxXrBWTnL73FYz2c5n+SnsT2dSyINwQXj8TBNoxR
odLwZyhp7dgINonsLgn7SfH7sizgHGKbbOLNfIUmP2GyVa7V5EJg0/wNheZ+9oa+lxifi35lNoGR
pxkDTT+4NWKiGjLdk95cuDCfFMlGj8s4aZB9v0lrXCmfkZCJX+0enPAHNF3LU1DweAPjzP/5p4Ur
KZC+deFJqNVvAuAKxfQROU5WKRS7Y0lPBZXNf+RgNXH3ONeGOevlRlA0aZ6MfvedI7xbHvPt7Qm4
lKAkZK4B1n0+7FQoZGB7U2NCCsL4L38+Z20Jkk3SJG0l/DuvvbDnUt9dqDZCAviEyXvMz6BywwEw
VBgwXpkHC8IKpF2NISqKm44ZRkoex9lK31fwB4b6OKxah+E9McT/YHOeP7uKrlmyBsPLMi39fi9I
4YgPI7vZZXtsxze9TZbUUSiH4l0DQKzxRyUsW/0VT6j9R4wcMb48pEAwMVyKQqbRCx2+jHdWdMHC
U8wRd5/DReZcVL0qHlVGKqYRpy3+5IKhSgYc1vKZ599M41NXO3vno4JCzhMm1Ixw7u4QBF2EM6h5
I6w2kuL8Fr3TgCbDiepDjVf97UJ8pydotjK76MvdFEsLBbbrJzJwpEHWsDk6T21jHW49YYJ6qRmO
eUZ8ttELTXwL5KzhHhiu3d8UIJ5xGvWI9ofJ9ojX1m/8/NbRt581t6EmhIKxv0qagPFHkm0MZOYe
/F/HpAQgV3u0KILKiZwT+ddAP2ZDWkEb32V+rjkDuhs4x2+HI66aJs7hr3hCX5IYon3PD2/q+Qre
rFBMzDZvkmPnig0xwxCH/3WbPc2WAs0CfDaafHfV1w4cvOLcVN38v6Xj6OFX4ebzG5KAGrtU1d4l
zZhgOtWkjmws7PW4oaFdC+aMW27OSm4blThqkdibrvsvtTkDz9DVcFZe8bFnwttf3828UmIMZABL
nMxbGjg3gWAzYj+wBAaXryUtOdQhctJGHqrhdZAvJyltGdG7e5kb9L+16+oiq7e2QwDxFmzY+cYU
qSO7YMR6HKetUn4G+jkGcvA4S07NRfPTkF9FSumVT/1DHEkhwyM9u+D8JB21dKf2AZLGtMxvmKeJ
QCS1pv+6geVNFtq2CkYZKcBoJBa8bZzn/Chcm/LgEGuVuHhKxcxFxTlGHSoC+5z9yrxzkBsmyQlK
tpMVU6DpeulMe2rfY3+w6G7I24s0NTdYa3iIMg60pMO1LzOoAXYwaLa5ttpXnb8EhiU2pmkAyaoI
adU1hhdbxC6jdSlXJITeI8xCYrtjq1Sz6tWU3PmVpHCZYqDTojHbcnCHzYsQCHIiDx/S+0biep35
WyiYkEfp/20afT3vRK6qkWLqhp8FpEtwK9glSEGXV/tSMQGsTRERWpO1I0akFY6QudX9jav4eSN7
WGrmudQt8t3fjROIXhjJ6mnHHrauKqrTBkbi43dUKLjmU7si4duLEVkte8Dd6asQEpfGygWHtIh7
CHNwaMGFwvG0jsKjth9B7rMV1q00UvydDeDBeFGIQZFo/Jgu0gzCs3k6hP47MNL5NaEaqBo6kItu
UyKQUI5Lyg7ftvkGG/EZ0BZ3PSwJIB/HOwWNZFmAZP0qqjqHCbaZvILBj+Rm5Ca6J3lcfXay19Wb
s3hbAGvKjBkYYuQWjtUoSgh4abNrynlhqyZrEyWiNpTBpEwn061IBAgulQmeQhPcdYlR3vvV6u8r
12oZGKJeXqvOaUjEDUnlzOVZrCrEVa6bx7kqEPvuB+97tH5sDbGkBhPS5z+krO9Lplt3hNustOaF
Avp3P3JPzDpJAQm7dXUMFIbbph3mrh6HUPFUpoFZWbjhwanXnuA2ti+c8cJOBIoQQc/6ZWK7PBG1
StrUGfBfiYYVLW7A1r8kqJ4e3d/lgDYklFvbJ+gRVmDq2Uc7qKJ5oRfcPKRvgP38XuNMzI8IJD8L
ragJ1BsIJqu9c8mSfOvwQZHCS1u/I7O9Gj3ym2aVhI2jaYvdjG1cGyIhy7Iknz/5TNtwuIqec20U
sRqu/oU31nA1Kdt/XfFMuJCGKj4ntaR+h6BriGeziaXDxS6IsRQipBOk9zeNJEGYSRZdsOoO27rI
MuAm3gYZhURIjm5M86kw2JAJo/1I1uNaPpQUrg6JG/6yPufcTEzcicJhwaBQ2qXnrCeEWY9eSWST
umJ9Nhl2W2zCe/LFwm70AexwAON42rrnybCMtiyz5Zu3llyElXgnBmZZAze0AA7nDYTkqwXv2+xv
Bj/4s8OW2X5RRGqUoBCRzP3CAnC4L4SIzm0nHOQNPcap2qngpn+JlpZWyJZZPE9mEtHZ8mb0otes
/HVhHAka4ASeG2ZOmM1fWXl43yAAZp6BelmEZCmHNBgQx1IFwzLxSwHANa9FMFeesUKeiCa49vqR
AlTpY6rGLpLhpEYGE6XZjmn172MIQEPRYc6+N9vJJVDtH/7pPG0DoDlfVEuBmWs6NuDBzygTK1sn
r/NTc701c8n/Y4FqSr88CdeqXq2XOs35iX0I9whgFLMU1MZM1ljxq87yHFETsYZDSNCMxDAve/Md
EhDNcbMjPSg3kkRtY3kOSNbW7ToeMRxiU3vT37cnBprUFb6EO392TjUqYVm4gjkvGXkD6YpD2d+0
OnW1xw0KcKFtPXNqz0ugzIL2p/zBK1dPn9LSLgQyisSUhVJTB0zRiww0RozCq45+GAckJvCS35F3
eEi7+fgetC7+LHtnUVXlxNt5KQjQNcb9Z0ZzkAvQShJTwPoU5qHkOAyyarnd6++3r0GOkt8xAaKU
ft5SrkHkNCWUSrnUwxRkcZrh5I4WETl1WAyNYaet+6bkwVN9ZD90mpc8EUjeDXun9dsd7THr3V0n
SGhzebNO8GNvtfQ0S6POtBOv6S26QtwxfRkLEODeFtatX539UICSfrEX7OSVL6M5671adY5oEJD2
4TYN23PqxFeXqj4bDa5N9ELoo+74BdxrNWsQBlXUZir9io3Td8iep9eiKggXwvcl3Gqg2wlryMoR
xKehrRGNXjMPVMci0tkRvKMs4ITJndU+F8+qIlZr5fPwa9rWetPSYNcvP1S77qiJtvxX4YsjEC6+
k/jMtII3ieZYJnxdDARsr7SHQaUxni3ZbkRmuDGvt99Z4cilZH/+IZB+WB418MjKBGHfB9EJ7Paq
iCXm5TScv7Evy59jLR3nKwSK902UFePVgBYvBKdO2Y2wsAHiRH0QVnKOol9O8VfcvzuBDoaU9Z2V
rgu22omf/iyfAWqwSPttbSODJSZ0XxSiiXIWWmv4kb+lgjjOAXqPDeFhbCaFbbq7ZKA5Pc6fJFFc
LnpxxfTD4U9sw0a/bHBTJGKhbbro7RsQ46KtuK1x728nARZKuhy4/hP5rUsD4Y8FFZRIk/jQcWgB
sWvATHVctci8a52poZ3kYR47kvDzqT/ZMi/3PtY7gskEDJBXmu1mB2JJgc6OcFJBqiEl2QgIylO8
lMisny9Ee2Xtq4JxMASfqUhUCbV4vot23ksQmjn25SX633Z/MG3WR3jHcRsoOUjzhWESGr/ynx7t
rTfAkplLrJC0VyINucuLINAL0r1v7NlZMzk2eXPAPDpMvM0dTJBNoRpxGxt0KwqKpN7ofbO5oTEj
BIA4HdtC01YlaTUxBU90o0TGcU+L58H19l0maMLmYr3+/kqVh5oHl0RNmDR7Eqz39fiiUoOIBfia
IONl9USzOELLUp3Fm8IXrMUNM8CZcGu3OYoeoSjzBP41q7QwuwsF2e3hu/RXxyzLYdtK+qsXtudv
cV64+5deGr0gVMs0M5zpNKkfigSnwOH1ZHhXbXFReYAhdYqH6LAl11DAr2psWRzFQJF8Djip5qju
NS+Re0hcsTD/xsVXLtlHkFzIGPPWTAw9yjs6Vkjp1z1zTn5B+PF2Ajuv3XGJa12w5+K+UHJu925x
D+k0AZF5NDC+05p4y1xnOZm4tO+YEYHx1lSWZFFB+AKb6PzXzirDcuFyaRArDN4IWcxp4ass+/lq
eI4qgHpwAyTUWEpDGyEFgDuBseCNm1515rGVdJNI8VexdWUA2rs/beT9Nbe3oue9gmyX5l3aACFm
p0pFfS7OTJnlRXxghgSGrBUNYm8FawKb2RXh1VQUCkE3KgV4/zyCA3nhseT/EnzgThMrUdz38Kor
0mbo+HeDLGkdL52gIqYrcOzreXxqdhIUAywt/4F1Zkcz9gAIwRd4txEJ1x+lMV6L9pMvsXfbl7NZ
MC7Z5swvsYvW1IpD0E5DcDA55xW9+t1+Zmmlwz8mt/GOyIHE2d7SH6OTmq7uQ9QB0tmHrZFSZbrg
qBH8cWAFac1CJEenl+yd/XeHCUZtQBzAVkAlAu4KWSF1NkDJoe2t/HCP9TLxjQaH/XrbdlYdCZMu
f2rQ5nuDmbxVRBOgIzM6HiDQfaQk+34zVeiqiv7MZlJ25y89zrEDwUqi9lfegvaQZGbQFOqglpEu
EXgOIZS6qCwUVlC6mZqKbwcMZYwsPuy6skzNS2+E7b+NIPzGc8+XKQc7/5Kw/2l30uCfnxGB5mYN
qzMfDB37swXmAfyNnTc0z5TVuuAEDFvyl3ku0aMB/QBD3KZi4aVR8PYhf7iIVtMgcuWV+W+OoCVe
Uez02kF/RJjZiJP13Sl1GUIvcTdxtKdUscT23WYlGOpH6amwC3mYKHqmB21ZlhvpXvgwsSsLrn7F
FaaTewWO9LmXuSQwsyAjH2dQUsKqQetJaRSoxOzvyDUwh3EaamGVmHHtYTyEDddu7rbSlceppu2g
NGaOUPM048jH7qJhPhJHKiczBR9AmpcuBrCbDcbqw9k7+TnyX8syrHdRJDYMS3uehT9hwk083KMO
Uf5cuYY0JJoXOj3gYmtfr0QZD5OIozoHFmKp2Pp8XcJIqlaipG7Xm53wqrj5m7Age857hGfJgxqs
j4LIZxhcuR36P5kQNXmJrUxdM32tH5NKELcCUru8/DQ90g4mNCiBGhvFkbt7U43NbbPbIIqDSB1N
E8HgaaoaKj+KZPuaNIQOsN5JogMO7+ppfpZwuOSbXnn/EtBm78h99SA5mzUsD7vvyob8wvZaFq36
VtwBgxoku9OgSP1Y1QeTqaI6VY9AeeCQrdL1mW4eSMSLjVjY22Et692WyAJzUC4Zb7zSGFJ1S6mk
vBGwDKzHAVURdhonp06naJnawVaC8S6J9n2qq5NNgx6kZ4YR3IKg26a8I8rSH/BQDTvpMi/n7QE3
CQOTqdXoVrE3lw2FN0cup5oy/UrVOvBphCYe5QxUAPL4M0SSe05oPfIy0YeP1uyqGIqmR/SCD24O
1xCJ20mOFLf96bxOIHLWpHa3+wQXpGEQtQQAMBbhimogGXRIVp0xKHPO80YR3DcxJL8bZnXkFJg6
rlsfDU/CPaYarU4JTlUsXgzpJkdiFtBMPuMh7JUdR0scU7EWfCkGj53p0aeTbnJiIcxcQw4KZ6Nm
RlIq8skM7qNORpjq+ASAaNwgx8AUGJpI8SIr/J3oTc2JhB4dzINKAaK02buFKdeO+T1oE5orpLqT
W3ODAWufYhGO8+srh4JyI4memYL2h1yrZhDm+xV6XSn3bBQb5xD5DnGUvdYptw7TFbEqVMVJ6eq3
6dtfu8Pg45GTuNBJwEw4PWgdlrw7dHJYq0foX5xexvn4JR98s9/pbBm0aw84RK4x7pSRdzxPKFeE
6pBfau2p5eCU2lIU8bCopJG9HcPIq5D90b1Yt6ZOPWLriiEU4UiGD/w17vgZX8BH4vNXZDHm/G7B
RrcZ6/zhgp2qFdVHRJAUqtGVkSaC+9I8f/DlWOrLswTelRbdOC0DSgVPIm6tabD2IeCreQ3Jrjgl
+8hNPdcjUOjyXFiVXm5zrTxe0YbRGDc9acoLkx50BEdNq6rjNywLBGQj8LBqAVhRIsNJAke9kNCs
ReQC5FoRMf0dWWvWy53dYVYf7oVzG0m52nqtfIj1iWnR1pFUCqnHFuQIzBdXMa2PHWJfbfeGBmat
cjtRPF2YHrPkZPkqBwKZ4o6y7UopQkOyYB1i34ZuUMPuShVkkEgGzLeRp9nqsoT+piBJ+AEUFRrq
yRwE+j2s6FVpquw+87OXYOBid12gIQ8wh3yNvYyFeLUSQXtvbanpj7rJaHJUpGd8KjqrfKlxh3F0
as8uYDN5qc02PlTVBwTJqjj5NGbOK+qlhIIPrHTcrRtGV2PsxfH/Wa7yYai7BiT8SinWjrNPOB8m
mtLtp4Cc3IwcruScM96IOW2aeAKerVIRwvo3gwDYMyByVC8NfesAfIeudDwmLgE9wVCpl/AogXR5
Kt23DQZijrMp6vKxo4EVLrcKIPn5haWNwYPhZFDpA2ezrdnxR58LWbUd+ORmPsMch2zmJ1gh2MSo
ZRc3ShpCjzzrjaC1xpro4Opv9gV4S16c3DASvieAbk4dDdyjdRf3v1vYOJhPxkVreD4uAYC1awG9
QIkxjNK5x5JNLyDqbuERHiXKJSrHpVgND0Yn3xwTOIa7cJqU1hrWFYJZxb3mWFxN1khjQlrqSbIk
m2uhuQ8qWizn/b9HHGX0SE694upQVi76DfdQv5pw1Gm7sBTDlWM0gAMErz2c2/blrAPdFVxcIlS5
N1l5MeZeV9TvODEo67Ay60V7jfWb6WbCvw5zGK/zAXqD0IEWA9ES5tCqR+EBzktljycoeRfJbq3T
Fr4wy2+ktbDdV0ROgYNZ0zTzu2MYpyfgonbMQLj+LJkoxgF6ctH+h9fvy/XzyIfknUWgtG8Tu3/z
mkl6BQVc2TyEPgzFE50qRkJXg1lL5TjK3IW/KeckWt/8RcT8A3SOkyEbDbmZgZoxucEyrXTcvHN3
JHQe0ePwCguKNknlf1fCF3f0WkkKIj/GGfBRwY1O/cGqXMvqv45fSgCih4K6Z6gB3OuBFzJ4L4z2
s2zFF5HMynThDRz+rshnM9BJrCWDehbrU5Vrr2gD78ViUgF6XDk64NN/ddfcmdwNwa+6mulKq/Vd
dA9evl1cjoLK7d3IVZdHZvTiwyGGhEuS0URBQ3HuSlgFZSKZnbw+2to8ohdqr4vaycY3+02jwXIH
OA9m3JustcoUmDmMHA8I7mN2IFtsIs1rCGLqSNR0hiL06a0PAkwmdD6pTiovrdEsbNwIo49EVrYk
Fol+GmOIas09BlFEm880+gCOpDUrCicnlTp7oTYI9SnnB5hgKTrxkKsgPqyf+liYH2Fe9jqwjR1v
KbfQnTT88sYID3DZgv2zR2Z7+CA3i+sBGZBf9V8wS9fll6V6+JzquUeV4fmqgMfZW0k92D7BUF+F
lEBdN9mS1ImGx29+u4FRenEut+hkEN/BCBvOmK4edn1y0Jo5a54RUW6nr+cglqE217vcxzjVQ+zm
afpiXEp0eKYjn/5TpZiRnRyCpUsMkuus/Hmcq7ZariQ0G+bR205gWI5MwSlSqYeI39kJMKbvIiX+
9EP/Vp4JJvGoNhhH4BazEVOJr6UIYCUuuv62/TbDAZyI7kf05I29rIagcYf9ppJRmBQr5DJ0JKby
tSxbc3NlnDTeS/H6YDicWmkN+Zt+gbeAy+vMCbDcMU4XORToNE6lxfQiO5aGe9mvv4VGPlapYR5i
W3JhLKiEH5un4iS6M9xUcFEviyCFeYH/OAl7MctHByb+33Mqt9LYzK+sAzP0tAuxFOeCbq7d06Dg
wpN+K7gL12c15u2P+KJcRVKGeUoJvNqFOtZmJzyLXxnd+81MpTTBsS6wh9IB/CIbHqymHFOrsrr8
K33aoCNoNxmud2cr1U8ymYu/xUTRXzYF12CTNfhteyvvtQajUHQfolv5IzcFjfwUJ3nO8gbmIQN+
R6Ve4b3vhNwlffqN0GlqqtmlmCtwFJsoqQYPiXM18TIc/HRQwubbmiGpVIvI1pJFlahhM9vJMcCR
0PRe/LzRHg1Rm4i4Vwp6pI/qOMjwjpkhdLpzE9cbN2RK6NzayLAajlK3Y0UpYaK0BlpwkRrq8KjB
N58zw43ePkR9AqakqBLThSEkhp8Wehs/VL0CCqHSFuWRVjCMA+UQlqShl3CvvDHbYTNunln9Xzhl
tLYnKypo82FuurJKECF6im7wfN9wKYVBwAyhGnFG8giWv4PXZqLNwC8/Qta113Cok2rbBOV/oW/c
8WNc9ziU+KoJ1hQkuFEWZsNH1tiyEF3cgrc7EvbDwTGvdc8z/pv3DFNSS+d4rURfdnB89KfwJbNn
YLKyGvRtE3tGKaKtbsBSqbMQ3dxjyyvIp+1kxFvVGYM1CqQdU1zkIu7blwZNy6kHmnZCHsNLhTtT
4dyUnawLFuSE8LPsExtWQO3HZBCtvj8X7/wUUzFYRHCeWkEtPmqxvXcF5zc1fJQ0L/KgZd023nGQ
3oiPsOP+ex71s/3pI+SOUDZwhMY46LT5r8ufl6rf164NbNhaRmEVVxzAQGmUHLDIrwj87aTthD0P
C8YrDi6c2GiGXVbgHrsKaNvqqwOBKDuqdF/WgflQF3sC5HdlFFcSklp+iPUVeYjmuh319ncAoPjx
3os24mnf9HaR1ggWpP38KYP/BPcHkJyb7dyhBWasLIEKG/NGlJRSfmEJ+mSVxn0XY0gI4zcAlc5p
nrcIQkJpLY9NAxh+keFcwYFntfWgo9MMixTrBrPTLWmJ+AqeHj25BqdnTvvsN+6NbOu8h7FKtHWt
kzmaQT1zfL8JYH6gi8+dtfayRFVh3nvPS5oC1YOtnJJY2pPGAdgBue8QIaAEF5ZRXmbv9pTDxFYL
OkwhGRP3WF882o0vOFjpIYQaOHgGBBMPdlerqGa0prPXN9DP5bQapAI2HEYDzbrQabrZ8U73I0Nx
9qSZ0zBm7FXCOOCQhHsXkrXR4ZRpgGX7QknZ00ZPLVRWN0q67X+IgUWHjAmoVWJQ0gWeQ+EnXytG
bicFfNbUUsRC0O9jU2UQXfM2TqFHQIN09GPfijAy3egcgAohrxgG2vmexXB3zmGuLVMW6bTJ0WVk
VtgTNR0fV4ss9rCqErJBwpFMN3X+DLCCUt7yfnEZNNOnwnjvoVY5QJCNVCvPt4/rUFHPCKrtNfjE
trZ7n1JxNcddTyO3YFBCi0kBm01OCJdlJ1ItnqaHJp+stgZsfH8cj8o4OT8nsygcDAHgFLz0lPkY
ZGtpyZG+JNUEk6ataJ24TllGVcDkcOsI1H5kCX1kx2ioe7axuqbgltirzqakBb1Lzn6t79qpEX/c
Qp4zXUwQDuElWc8oI4EE6OGpwQ8bbw7zjRJrLRsOlxodKts++8/juieygkoVR2vjd1s0kWQOiKHU
nWAik25VkBW8uPzjDeFTOn5IuUm4a7LdTEMrddTASUJ1IZqzSElIf2Et1HCVVOvOdVEplINePc1o
aEMzSasvkRB6zXR3ZSha5L6twBEyn/TxLiy3/z0y4zFv000edVL8ggL/wqSZ5PB5sbLVPLHbTsj6
0h4UgHDYlSfHEEMuHpw/kpKn7InTIKD+t2dJV+O45tQpyEsHSULYplYUIy9UQkTi9RfL1D4B/MK4
URmeSlRsFabVY2zwCDKSGf6bn2bAJo81F0wvI1P0mOhBafUGfFl5O5KWrMTbiDVNr5Z4Jj0Nj7L9
vh10HrolwblnNLLWynOGW0KUGsc64SN/arrig6w2wlmW6gb9S9j0fTMcM1FYDVfytpAMrRPgTHTq
WIx02S3Oum4wYk14AllUbknMnH7Wsst2GY2oxbpVeug26/XzvDFKkQOp8OMSLP1PuMY54oZJQPoa
qjzGCmCT4SAK/dNjUnN8lEh+VZ2NdW6EUvYFUAQ0Jl1CGfEY5NKHs2g+byhc9RJMp2huGt9lqyO4
TDMQH9AXGxc29a5yTfRYb/lgT47I4rIM+uf/eT76qVZW7NJCkZwdi1k1r7t1FxQ6y1BZyzsYrHre
N2Zq/CKgKEybHPKCDayqfhEN0wUjqPcOHwlCnE8cO9+GWPibW/yfsfzNRvz68iRWFMON/BJwRvg3
Xw4v1L6R7aML94s9rcUeizL0opLCKTJxQyNZeF0v/oZj3sZs7zWS63Vr8yELjD7eO3tJpkrvHUEa
mVLbHDEqebKKc9px62p/NRA0yblnQMjzSIUCeDrscQ4Wi5IAmtwJ8nQzcFRKUmsRk0YB7FKowMyX
WpHT0zhNbXhLR44/y+xIefZClg2lmzdBm7f4dHWS2J3BvipZpi+JJi31GIBWmduZoGkeamsjxEdi
LcS2wSO2as9nxOBvCDalWIPenGUqp9x86ruzz8r7OArXeLIwBdNnUy/PLonV7ui8refb/JxxjVdl
z5tGZQIbdPgRthTYAZeIyQgjs/0aT0GKOUUGSNND90F6VSK3hn/SahbFDyFembt48fcXdLWqz1/Q
7l0E3150wcpJZGm0Tzqq6WxQEpYoj20EkLrLSymTQm0jIAK7YMsJoZU7bJM+OOcNgDC/wYz3Y+Lr
21nM9kRlvAiZuTRRy7rQGZHARwJajkxWTwWBe+0G+e7qg2xFLXeI8s4sxaXI1RAMOlsuWz8hyOOJ
PSt88ToN3hI1aw2HzToJcIG7i2bp1+H7AeqEgNNw8v1WlnMhKQF1hlrqxfnvIPYheG9iKu9XDtmY
LEiHHAr6n5VGAgqnm9QwXOX/M7RhtHr5hbfZoS4RI+mTaiJie3JVf0dPs+iKs/uiYqVttIDk9KP7
KakhMn/+bozSLwlFGj2ebVpe3DgW9JRJl79kl3zCBqXh4+YK3QUoTMXtkAlD7BB6TQVgOmaX49MG
TkQvxhOHvZZPdHaHJhfXypR6Ha6vpHIgmVpXu3UmhNUjl6QuX4L2arw1u8ryZlnm0Dz5qBJqvyHZ
rrnjUm67CW1A4rYykHkP9OUB6FSdZ5EZCK/hw2EOxVbBZj5CadMGs0PWL/G8iioTHW4JcxROaDZE
D2ZKRk1bckj4EJV7p/HZ9w9rLNPCXEyuUUi7GS8EWmBL9QzsLvoqMhr+ua7qkj0fj+3hkdmTsSw+
pTxTfD/b3Y1cYNMXeAsVJ75OspJ+kA7fQCY0BKawWX0TWIEgd4VUONm+IS+VPxy9oqN9zuqkNRBU
a/gkY1f4pgz0zqzqoQIsglwCAWuxfJgC7SGy7RZauCiASO4SjFOTUDUnUuArDpyhJPOTnnlDsNC4
HCtQ+dr4HTXoNbiMAuU9ljNGccNnTX3l/4cJQJbQI1qSxOYLH5JjAft6irdcJ1bfzVhcW1zaoQzR
TnI7Kk5FKIIIIdzmQq2uYeKaq91dJCDj6St/xaql5oTYKhPpCq49+SZw+DQeEUbWtl1KozxmR42a
6VvSi94eJ5AwnzLolN9pa3dmyeV8DWjd/VlDyaT6NO0ipa1yj7ro4Lg4/9GOHqcQUH3jbI8qgsvw
vLnBcLYzIfZ93UXeQwTPiKQPlQtt2aO0UudlaskQljzahB9eHCaZJTUhtssHe6Dv+rMz6gs3J8Za
5h7SWoemJfInJ/qsaHJCYeGdIoz5pNSe1H1TW78rRMXEpxuU+XQC8GjlQp8ocsfW6jat8itcED6F
+WcrXBh679S18pM/wiOds4qxFMO9MkoM/gZTyuJ0UjuzQwn72XqCzc7eZLWGFFqOdSb5NnjB5mYX
jHV7GKHpLklouahlcR8eQ3tLLAHGvmkAoX77DiViUETzdrZvkGJilL4/5CN9JJxtkp5gjoXXZgSR
BRZNvfxfRO0GQW1SXPDAeLXIN8zYmKlY6bd5YX+5m5NnWSOkJFVXefzH2GFsl+fgO5S1gufa4R6l
7qQFp09n7juLTMtyoVyfWn6EnY0FcpYInx/rMRu8KubKEepahlbwKEOXchBKyve7/Pj7VWUpKH6K
rD0/IkgNC3dWBdieivhiarIyLPqo42Mkxbfj9k/R3kbkODH4oHaJZWEasIEqP14Yv/9NAV+x2jjg
JiygFl61ftQd6ZKMlGjSA/MLZFgNMXHXrBrF/Lar7sG4+xDGYKcR9UUROpQkDCDJIIRY2NpQPa88
1ED7ADzsgFiEU5IW/+f1ozJe7bDVWAoKgZ/RqgfoGSkpiKFaD34kVhPRWj6DOvaiLDEYjW0m8yIQ
ELD4FwV3zv1HLoYxku9BXA8OS7feaT6gFnyYodeU6eTno3EASalrqNZ+4LcSQ2MoBeyMLlZid6B7
Kz7AjXj96oJJD8p7H72RLWJz1pKYpKzmxjXaTwzXmDe30LmekQFtHOSOmFHXtBEVtvKTuLvu8UmS
9XJ7g8PO/YT7oY6/yBobRyFuAz1H8OTmDcySq0KlrDQjiPbvAVLSgyxKv1s0rX3d1NAliEl6PIBf
G/t99nxPS8HsqHn+1CdHWjmuo8mFQMDwXeBiV4qZ93kguaPDihUBZOWnmkI35rIRQRNiAvrM8FK/
UCRaDMDSzh+uu8IW9wrvbYuXsnLCIxJaHKyZKCgh3e2jTv2yKcjiS8RVBHXKfJG2ZzymlznDl9Nt
OUprRy9F3x1djk3orLJHSr/uCM/PFGvBqVqnDRRGRCYZfZpFqJjufwJQ8nXRRdwDCOxz+II7oE8e
JVh28LC3gMuhJDWL1C/jF6n0Fp00a70T1pxkulmBeCoRkJZgXbqmX1lLSE4lzJ55VZdNdCZ5ulpT
raly7h/7KcHY7pajVqATha3L5+PTDqfG/QfBcbjZowqxqugFA6R4k4UEOSm2VODBAsa84glL0KHx
HxopD9oeim4CEJsCm/68zc772DtsVyKSBCpamA85nWvKSR9bl+rZvWJynKbpeQiUuY++T8pQxbpt
EPDxsT9bTq/7UidJYH05qSobCmskr0Re4pp+TBHZ7WHAg97U/PIaqnNb9cpGEFJ5Z6vzhCzRaeBZ
wyknq3r5l00IeW7F8yl08/LbkTshdHcQuJMuWz5DGQkiHUz0F7fHmIwodf0Yxydy55vjiIlfg2Qm
urg/xCLAXagiv/Ov1SWxXKNwaHpFdz6014k9FGdOHs/qZeYsPn18Vew8/zHVDNypOSz4tC14kRtl
xyMX2RhYRYW9gVzTlb5TimBEaDedCG9wM5GsdL2Gq2E1gKfMFYSM6BeE/EehXBVzCHHpwEWw2SOL
YyZ2koHsCTuqwrXXBV9e+No1fpLlefLCHjolVhpLS47OCMdK/jutbIYg69IAnuwxbFYPFuyOUoxt
4xBcIYNoLuVMT5mj7skF0xNDyv2uAWExECN0jWvZBxhbC6d8FHwyD+FsvsqXWzyotu6VKC0tn7YV
A6AzP4LP1Je+Guz2KU7iG58fM9HeGO+IwojUiUlSaHKWjX4wWUH5bvoO62r8hrpzLqnbQ03djEPH
3EWsZBCdvD4zENeulG54zf0/vFjI76I7xbnImlMu6fJvQRKq7+6mdfboPgW54o1MKpoD/+WDg9kh
KmAWgwueFcXpdBP6nPp/uNKOnwwJfs7gaikbvQ8UZ/lNL6S/BTW0jWyi+6mssekfeCDRcfRGBAEK
Pk6uZRSyeK4naTaUOcbmyU1h6Yu/EukNJWsLeOZaOKuWfW2N03Y5AcXO263ukksz9akQjDazW/zC
jjPE1sdEpXcyaI+4ohsWweRbjdaJwoql0Tj9dUMDw6L0OvEoyQMlmf5W+SZ1kHVSGf+kfB1GuKXc
oQcFDvXNDeRiO+HGzNXo9VRsJuD2Gjle65WsYVe8/W1KOQQ108+cgINOY5umtrLqEgJym88W+5ei
uwym1RpENUxKWvVPlI5V8WoHL3+zX1tb7FRo7/AeJTnHSrmapTgYzQjxesuEe7k0/L6g+QDspGda
IBHlkEodpVc/ww98HkpGvD5GObZTzVW6BvRt9Qxrn6mMypddWUvNs5m/sWKOFZAi8HlhGQrvo3eR
aiv42xPxkovAMiyyci9Vn3w669lq20QW2yxV6CDVzz+4aCsXLlwxSJnn21lyopWUkB85t6u7fZUD
KIphHSD3SX4JUQ2WE0b57sZZAIjXGyW5DsBiZKIyKLr1jDRdjJ4eW2v2mCjinbKcfT6CxUMjMef2
l+Knbmsypkv7WkP0JGfZ+M2B8F015XJz65pJ5FC5WjaZWyY6M4l+rsKyh/RR0DXsadymOeu3fcLY
QbHUE8UtUKzS+8NWN7GBJ/eNw2W3VdV7VmMUU/MEubz5/B161Y/Ut7a+EvpslDTw8SpfmCmMMNay
3A4pFYhXeuDJ1Dd8xWYy6PrBps1tPUd3++eSy0RDhZznLzOYqq25ZdIAcjzoNE/UhY8haG1blVtd
zWS/tqw+sa2TCp8riQd81e16K1W7dCap1fZo4mm72kDgL0/QGP43Vm9x5HrXpxIs82l6gmurzoGu
8lV4ICYoMO1lO9AxZk5BYJJ6Fwnf3WToQTGxLu4QDnhJK2FcRqinv4xtOvVDRGN8l4Wk35QQgMp6
E8SkUui8wcQ31u2qx8OXigJk55GfyXPkfdf+EwQu1+zmTgX00nzXIYokjw8wkAeKQjPxDX3Jn+6N
Gx2QPftkfj2wxzfL0H91kt4V0USSPffmEcbkaOLwwFars7J2CNBAvI1QcpFtn1eAYjj1PN5lTjyY
mKQNUo6KoyF6gwAius/e0MrpxPgEyoZsrxmibGxnO1f8CBx++twYC3Z68gajYeu+gLG0RYwbzfP6
HBaZnPuYajSxffzge83aVKLxxpYnSrauwZCd4pL9BzsQC3OShmmMhhOFCf2yQYDrfwcHQx9A2HAM
FRq8n41eGWRe7mxuPU8u6da4Ym8+dhIF1gnvNljDmwxGKj2mye+JjiWq5KhsU2SCYUMo7DSj6jBw
/KEV8LLfMuy4zaCMvDRtOZYiHwmm4Nef/S/LtTtDyziHbOxPdzbf+6CIOf8tB1O9/L1FIxANC7pl
KsdQwtGH2F0zOT7qJgoNxUSAAN4Ckut1IIhN5o33Zzwj32GyIPHZqE6lBQ1WNn2rSt8NqsJP+ZV+
Ry0z63vNH9C3na1NicHJNwaBC8p1aSWFHyn4TWb3ImC+JvM8ydL+RO4nlPT6QmkbjaufdySfizv/
lwb3HtbPQj/tCUE+zMH7t2yxWsQ7rkqF5CNkU0mQMrH7NZFKJOqSR+oZhcSdpTY33XXCHZ1pHo+g
pOcucrNy1HciWVbt+DMeJG/a/LB4+Js12ZybMGL7dGfi7aXjG7JhFKiJsXhrFnYtUvAY7MWBq427
K78GCmqEB2jle6pqN33t288TIWo0tTdzKa8MtopUhAlPk7IuVfkqj1BP8/M3Z7ZpAkSaseQOBVX6
tqV8lXJY/8/kQ09LU6cXF8e33dKzNwnWjpR39+fvzGwprhWSzsQHd61suXO69mxx357VXZ1sZFrN
64Ps8SVCqzX9kUd2AQ0lBBhk88jQ3eh7DSEjcOgoREvczNmtEO6/84KRMyUc+M2rX4I6QhuMol9J
7DCGICPJl09Be9zqr3010usrMuQzewCQpxXXdrLHsNcJuasEWD1/HJHsoW59xa5kNZe/y1rVJYwN
f3fwDh+rO80yYsitXzy0fCPudrrUidsnDODZQ7Te+G2MyKLT0aOsPshvnjziYdc40osNkWZLyjD/
H6qRHLWfyDZDTrm88cEkS1t4eeQ/rmiAU1rQxwbSh3xwlNiULjg1eVV4VHMWJ8Gr8otEmwAOxV4V
urdpKsOu6lxxpbk7u7AzJfVa5zdFyOOP7mOWS1fWK8SBlTsDMVLhw1asi8QrZHGjROdDMFs470WT
macIVrIU9fkxUfdNTG6083TR7CCw4C2EgycoOJXOyxZfyiqt1BjwP+NcXtr8Ea1m/y4q+s/56dz8
c/3aTXjGpdnSx8BPLKCYo30lCY/dkHsJ8/FEyCVz+CWWhHy93YKNkjFK4qffS5TkqXhasW3THbI8
Qo3Zd/QCWaxY1bY4Zopsjy2c7E2gPwPCm7ZBrm4JcJwWXw21FGzgWRrZfKETlyRSwSyKaKbr6HyX
cOVdczlLgDFo2Vxa3w48IfLhClFR2fSFgZ2kyFS7r30ucGO6ZTh7WGnNeKhBT6LoNlqlLIJYWe+M
cULazTnq82cQ1TlwyWiyuLVySRYWX5OglFRPcgtcuOO/Ore5DuQHknecLXNjKhYymTm/o87N/NpH
+BYDox/Dh7L7rz1sBj4Jz77LEhYMSXRWTb4KjUnxsjW9mccj8HPcoBPve/VGuTiHRpCV9I/bz2Rg
XJw4vxAXC97vDqP0BfCFRy5C7yDuqEMeLZMnHa7sMC9G2Qi/5G9UP1Gr5MtUJ9KYM98pkhNWNJ/7
FyfAKAKioyV5ZDi7qQm/bXkwPzRWLIeC4T0/DNTZ7f/mS8on95N0LykcFxKhJnWchKhfjx0NvJFL
zlXnTg2Nk8wth9Ke1c+1sOJ+QdzMow0jwpBJ4vGqjMDzOLzRsp30gwz/6EH8qmjIFGVWrzxuwU3m
9X59MtYxAQOaXepui5NZmD0OKEC2YLiAIS7U68esyUCQsExx2YzTrXElV+zFtDNqzUz6Sfh36+fk
CERAGENJ/OpESYif/YT6yJ6AvULx0opPo5O6SzssTsksz1A7MCnmjCoBVVmBGxIhF4S1gpTWabA5
A9qqGQTbbhwVauRi3w/apiNT0LNvRT8hmQk2Fp87gkfV61qbEyeuKhckVwNpv9FDPtbP/uvAVVHa
T3fZOeDNbd2xv2PdMj7u2H4myR6htB5CDl/9NjQyvgU1BFEBs6s0fclLOSFWyFBHoHjN8RmDsDAM
wS8K0lkrP8N4i8nQ/YhqM7P4gv0Fo3nE9Wj9hJP5UYv1I7kC4d32jtylr1Ko0k4nKBudlCQsVI1P
JoxY6YgIhKuu+HCFssQj4ePjpmAmFEZGx26/eb4oi7sKCSGRxj259lJipwBOP6CdJaj246uLUyqn
fCN6XWW5q3wILZWVPW08Vj9MLU3QTmNgo26xBrBohOqwquKsEk/EqC6jLb6OUKlKaox5KMBncTNl
BspLWa9VpAGIH/hQkbQ6IEP66kMy91TRSJPhupTUoaiOC07OGQKHLnn/Z/pUtwe/ubcCNIfHZNbY
Px/cQLLDhn1jjixP9PBRt63Agmx6WeGBXUnP4ssOlu/6SpoXdAa0j9bnJWroM7obPMq7uue0Vgxp
2p435W3zbnmpNlX4T3Onbend0OVqTrgnt68Io8ILDZRvmupR3ErGilubr/ZTK6+cn953wCFVb0HA
x4jSYVzKmbnGXl7iVN53c0jK0I0PE8BHsUpcEbt3wxr12yuAXymsjnR1o9m0qp82SHooADQ4EHSx
Z1BalXPIFGwc0cR5oLQhgeQmdfTND0hd2rnjWS531bvrgM/oPr6EzAiG+BzcrdJ9BUnuVhfZ/efh
6nj805mQKuicbGlO/Gu1nleFqehBT+pWyWAitU79Qu5w8ppgBYYgQDHwC/GILWr+9k85pIZTg/Sc
UChk2gmsZRWZQRiV1D1fAmVXrBM6JW99V+6oXseC5A37GTLTPevQWRasDxy/tjOrAfxokQNxZEhJ
AJxpBpHoZTx4Hfv8fCzBhqs5DinROD/GAIeqyGaY9ns5pAYXFxnxd/8a3CbcgvSTC3AvxkuukaJz
MBKK31DAkiTug4piVXjm9Q7aPiOl0v6rZhpuLnciqEpOMkI+ATPeNEK3iDLlpYe8abB5KvIdMI8M
Hxf0LFF7QSKZRg0t+RDL6W7Q09Gj7+SxncNZWW1tTMAh9mMxj0RnMC7Fd95B6+MGbXAx9bH6wWdo
SzlEcec+G9alGtHXvHjUSrhmRyYo9blC9cLFKn/H8Gu/9p2rKWP7EUgH7N/AgfIhwbBvYICtZ+GS
VYOxQEE2w0uw5+b01TgpIGWl5xlpKN4d3dRV30VhV3qBLWTnnNN3uDyEWQ2/mDzTJNMZOisNDc/J
5FEUM6uuDV07kpzH9FDHHxZcMVg1AcFR7kc+aR4nIeRvLCzy3SPiUTn5bu7IY8P5bWeQInZXlkE8
UFTGC8JEZVKdn0BHTdmn+AsrHpr1E4J+pWCo2HawCY9PxNsTYJDR5I6gEWVwdfoc4RHrjPw6igBf
mc4RBU5bPflZqYUKHiQcYJRGzauNd71q6tqZZ7YdpqlAGQWI8oV7uYmvKKepBFUA96zT9Dp24ziB
oeHIWjCDkfTUOTMdxqatYf2oEZ2JHFVNaQA2t92Sds/Gkgj9Q287vcrwfcXzyKptGGgKd6FPedkf
GE4iJa7BAvx+tVy6zpybB0w2YXmt4E2ID1Qe0kAaOArFuaWFWqNwrD0tsy2t76TNSrmjengPSZCe
rOXAVOQSem183WB9v3ehlTga7SIDJ1o3wiZznEDwyQRAGXAF/IDOUnE+lu1MwEJSesaJc/PG659g
R0UV6I4nDX8Lsh6fX+3Y5T0rsBlxYvFb35qsPrrGvSg5RojIMn/h72vB8ipbk8ccamRPLry/wBfL
ziGJabjgSDqWt61Bo/A1dYQ97Ej1KNIxnRWG/hVIvqQarur2UyTrw6+tgraniYrrn0qqI3VKZL4g
0gbO3VOqXBIXLvRJCKVdQRfTpcSCS2P3Z/5CBPykZBdKDgjk2rVRywq9O8h+8dgpOwF1VSc1Xeef
dX1CuLDCWyPyL39CiR5pwhRAU7a2rlidDczRRtgBQeZHW6tJQp4C8ymcLDel9xmvEMaOCQFRgyKl
Rtz1yOtwk26IFc7vhqfRt34wXZnYgmSq4eJ/VmumdVE5wNpn2qO/qII3bT/ipKBAx1TUGYD6/n9Z
rIeGNb6KMDr0kW86O4KvQGlmPzdSVuLw+1jdBgKsIxauloooQIU7SkckrBbIztDw5PZnxt1vKeyS
IGdD15Edt0Pq3hmZsawxE9GXbhN8psszVdU/VXABlxNdifyJeEE/KTymXhxOVbolXB0GOKT0uA9Z
wb2CpyXazIFgPn6okw7g9/EwvaSWONymu9/EgebpIjSjLhPPPtW+nk7NGnO2kC/9lZwq/Noz6UpO
4nfT9/mnSPkE8WiVleKMTeVgEkh9ZDie91DwWtN7NgHigyhiyP8lpDGfxTlAtmMWgH7cSRzWzWB8
MQq15MxgKhqOb86sMrUXR5+Z5UGEeLiTKb9RC13rmpFGUYQrOCbW1Vt3UifDZQFxdvvPNGf1ydDF
gZ2i32ZlnyTtuW6+xxNSVuOJlBiyfPkJ5VaI6dmEySE1lsllLbK8cxokEOwUwUryEOyKydt7F4Rq
NN2SKuzOca1dXWRIX4c6n7T2uGW/RmJXWaqHrxbcOfokpHY+4i1RXp2ZcyzOvpMjVc8b67cyjIAO
IHBEk/Z106AEhYB1nUNY8eJGMoTQxArRLRTnFlw8IYOF6LIdVHVWqRAlyALgi+5ZErUbd/3KF6tj
8f6ynud7jXE/UVHtNP9TjRhEfy3XezSiaKsWvXtLGg4K+onCSBAT40bzkMRMuy6hFlLx3ZwSnfDa
Akp8uX/K5vDEw5n5xulisuQLfaikI8oYMIm/i6unQeaJFBV1A95SIilJdjTAdwDmDKNswL5NajH9
j/z5xxSSWL7+owR+KY36HLg1054Ig6kKnXqqYc6ZXo10o9WGbcsDZ1L+XFcy+lyLEJ1YpyuULUQh
OzQfHx8BMIZ0d40LLE/KGAbJpWjlDcDgdkxjijcsWhw2zRTVcoa4TNIeoMXaX2V1M7rEcFJ43GTP
9r3WoZ01oiTOdmAosAK0+Kp/xViC0Bn66B1NffceZ6L/z+rXj8a48Gm7bQgNbsd/4C/aIvlvFkSU
/nI+rHD7PFxk2LqjNFRWDV3enI17dx746NZdVhbV2JsKJS+Ht5Rmw1fX0n0oyw++ug77YY1wlGl/
7g7u86wiz8ZvOdSa+uJP5S0/yNMIu+fGzyPObkZoRs4Q5pVEEzFjhQr1Tgqfq8BVSKgrab8CbFJd
c0iJ8V7b6rSpWGC1qGWeXFxf+HZZfMYXNm2NaeLekjoJYp99fFG0tqALPdudxW/S0F3UjeS+8HWZ
YeoDPD1rEQVuGqDM8W4kdzJeDONueHM7Ssc6B9hxtdaQV8uvfUFD7E/vtbjpu3J1AwiUfe5hDP8Y
cXfANPCALNjayWGLPVHDB/p2aliJRvWgAhBDBZ2Sp05elZ1WeVyCK0/E1q1TqhkZcIiE9IX0Keup
P/0lezxyJzNyOCOSr6WpKbNe9bXud5rwS4HknnVNSMZmM6bPSbLrB7Z/DxxBmDm2wyvyrNOXw5q3
IgcmuUQaOhwKPrFXrIEOdtPyATrO7RCbXeth8K2jR7mCDRgrGtw4MKjwsjn73PZVWxXhTGMdpX5y
P8VuXk6nzPm2ZFsq3o8lZtukcOPzrWVnaJheTytNF5Y7GyrJBj0HvU9v03UE1HPFcjiYW8PorNhX
W2FNNCenSDXLH9fiMmxYgVg34kyHnYJROSskJBJ5kvojdrUKEqbhPHWsnPTPxG0T7B9UGsG8DTA8
uc3SJ7XYtetOgnCWQRLwNFLZwyZ2I6VnEIVyj7/h9fpNaLg3DkxiwNtpdR/JEXNwQ//aZAxL+SwJ
0PdqoHC4RbLLiVZh4xF2Sa1ISxg5EdWXFKNXibisH6uuFBCSzLxiOVNmhPVxsdLRhP+GU9BwL46H
5FgpxlJEXM2VyYOPYhN/38/sYF9B98xl55koDQVzZflRItjETJRnx43NcdQTjiCyiuLBDgZ0Nbba
hM5vYQTUznXKt+cnToNXhaGDhF/pmrrjAZshXGd+ceV83/nz+3Vq1pUNBS8y/wiOdikUvEla06Lj
RdAlk5gPS+TcpsxgsB6xypdFwCDHj/UgZKOA4q+NIhfleIGgEkrqfLokoSTg34V+UuaEu+MVDHY7
wVrnGsorTRRTGm6IsPq4dEu3j7yZuXJIh/QzkKAbFIsSyOi0SZHv93fRYs5E13p1eV8SAsmgd3fD
S8IQUAInLIlwYthXMQXbd9XU/MQRGI1kA5wiDSN+N6uFtsBt5G/tmEtAmcaW6VPLLf2vx3yly4k+
IUCECviHJFcvYkqNZhW9dUIYzOdHjfsmEfKzQZAITwigg5Ds/j04w3aIwPuZw3K6JdDrOj6C9hg1
6vwqf63usV9PKLAjFvP6c/iUHGiPjG5aoi5jS9ul2Y/qSGerYxE5lbkouMe4XVrVFyVMLzAjvQb3
6B+Fp/aKeNCGntlpIC3NesL2V97vUGtqZ51GZKlxvXxxG8XJePz1dvJGTzHSuelcbdRyWaJZy1Rm
srhufyMAdV6SulXE9EyWAgAvbLMEZ/C7uvGBqcFcnrOYxMfQgu2qG6OHNPCzafmxKoMDAIx4lKO4
2Fhy8mKFYzKUWFwfdxTFVkEQQcrk3C3Sq0a8Vo4Qe1uBC0Isws1DdtO/Fo3LW9Y8MGPGINXSgaQB
kTRwoNXoNXeFZcoRzxu+o6YgcxYeNQy72uMYTWVzE8/WxAG1lGcsRSXo2Vt9EuKGpH23n2Wf7G+V
pZ2oXHqv95b100DGy/ygChQ8BNc6LaSTLmjVBG7ooaWyonz3TZxEqX5fsSGszrltBpJ10qVbUigY
WYPzislAhzSYZERC0Jt+LwfoPHjOtiG0XlkVzP9kIIsAv5FbRTldYHAf814tamXjm+Vv/HSOuxZc
BRSj2dt13IN9yzQ1kXcZ/MtvwLKLbp+mt2r5/o9CxS4wSYuKUp0mk5aP826XGGTBQ5z9+YgqmYK2
NA/MuiehoGHJkFD+TYApOxjUU1MVxGXvk5a96uIkOARubGmP5JDJzk3tG2u/ePx+i3RPjXD9eo7y
mTAm9bITnVsCwiIM8/nvBglBSxFFD3hgaHnT3446qUR7hkS/G39iGdpaG3s+7ibWHg1UImK0WrDT
nVNaKCwc2+RxUcRAh2HaqNZvU5hP+VnbpCipuXQDoogHUixqTmK2lZBxPetGIsD19sN5MnDPF/OO
WWwCQ4x+LydqmV/66TLCS1LE0l3fnhUfkLlv/Os0VZWWNgAHhiVwiAzxX9sNICM2Twc6qLldVRkz
nI0VniOD2aGtU+uKJ6nMSo5cJxtWxUOF/XV5iKyJMS/cKwVNCi5SpbLsrcve7tDlyD11sqBK/o7R
sZFQFDfnGToTnAOJYpSKZIJzdNQx07De0vLSI+33W0txCRA5X3bPiVzYMpXlQ7hB5q1LCJbHBupV
kfTfh36T0crTJijMnHN9uRaKtpClYxdUj2p6qq/SjtasBOe+BIAHfFbUpAPCQc3rLhuVLMcDK4NG
jNAG6EMjTjAi+DkMGXGa9S/cdklUVT3GoT7uZXl8EkMhgEW/sHyJw0LcL7nmMNyvKAb9Q61uJ9cB
1uvYzws5khtybRboVFRca6LC2JnruTcbglZc+vRyfPG2Uxhy8Xp9CVspukgATiKaeD+tplQk0Xyh
4AoAikG2zlVIHRM+AFD9wJRdgikth8yd0V9C6Oq1vhon0R5ATPVyYFmQaNbjFY8ABJ0x157gUewu
7ctXeeT5zP19t4xBTr41nymxRPzP7Dt1nDhcD8cXRWMJYmV1YutrvYHEbHNKZVg2hwmPnfMSV7ch
3tGZalHyz02v6CPFODYU2THB4ED0v6KoV5f6UYLSNVVajKHbdwh4l/62A+VP3edkkrr5QQeZl/Qq
3Hb0CiyZV0YjLQdfjIHh9oQn93mkgvZTdAF8zHMVJK70TQ/ClxbTjTC6L8EX/rBJ78IVDstbe+TB
AFkmHnVsPQdxwfx36nj3YoOBZFDGpSlS6zskrObf6abXnDdOGzMgimvIJV31oTjvOO36D3lwdHTD
mQcAfjm2Ge2qCOnE3s/SGLPP2ertNDR0GajMtI7TmaPnlykgfgIAnsOl8oA1oTY1lcbxGovwCFs6
RQE9ORRtnCECphmkFaAba4ApC6a2lIWNF5l7PNR2aaK5HQtcdeYznnJIN2heW7QPd+RwddO7ZvfB
Sx8HSd/YgQ1THhf/g6N1f41g3SUPP38OesXSjryEhPLzJ3bbC/ueRySIBdp9noP4KxQBomblcmgJ
8ArRra4QNHzb02h1RFz6b3J1vL3d/H4wlfAvFPT5lJ3Jpbr6gnz042OOKi2F3QnU/Abh0WqOjU4U
+VJal4b0l+TpxJJ8GA18N4ilHpvqZdveIICJ6LDnHg4hihlnWfYObEINzEehTRWOPvFoMQD0eG4A
Vv4/QE+eJjiHVDdULwT1pm4Jl1sIvAx0MMbw/cZnDJanIcAulnXFCtqv8qq22d/lk2tE191HI9rw
N+LAtGWR048aejwjlUCNzkYBZTuNYzSe1qmZr2IxxFfUImchuwqd6HePm1HREOKTgMZWOKk6wu1T
IZE4lI+sPqS1PNNaWT2KQbrWbctfWnM9q98jnCsHh5yGWuux8Ph1t6q3Aqjg3FkcSHFhRKAFyN95
TiMaWRQ0TJoGFKYHaerAOdZHZ1o7mahD9a6cc/O4yONj5VoBVLr4pIVVfOPCmqk+T714ELm1BREn
3fW8r6Eq7pSrWIl/cikkjmIZZlHELRQiOAvDa/bZY2KJntmS7YarkSMR6wymgziY62N/35UrNONG
Yn1SzdJ6lYQwAqKw7OtZBS/r6MeYhCPfMxkYs16fjVeB1icRffKWEeDpQlHMzgYM+qrHfb999/Wq
3JkxXJzKZccrZ8d0t98piLb2w9RWMceNrk2Eq7zz5mqUni9a+xoUPMgtM13RubLZhPxZMJZSq9mQ
8KxKgLFMPxAvyFsv17cGd+rlDUpEXKTYdZA2JGSfP30dspt8DxPojEYxdGZbHzPiroaxcenact34
NuvFVnwy9Vwq2JQ/NNwb/PFiIQtl9g1Ocl20X8UotedwQp4sOTrdPqUF+G88KzI3Fxg5ZbayAeEA
hSAXzRrtIGWr3cPUgNzOP+zbwXMVkAhirjxaWkNzTOIN8ypen8iw4Fb/exY7A3tUvtRM6M01GklT
S47KrTAwBRnSskFqlGe3ohrLwDIRvNA99aIOuEd6U9EF2iWz+GM9I4XpqomJiOElVfeRmRwQqJRC
wPOaVkukhGuyFKoPqLabKecilpi7HL0469JfUZwGpmosP3OXx8h4y9qXsKvEMKtlx6NJXbZc+KMN
v1depNI8x4CuOyHDjcfNdn/R96cNfBUepjiuDvrd74hJ9sSkff7aXCSSQSE5CzTTL6O5b0Tl177B
YSizBEegyh3ZtR2Nev3/wlnBFxysCVB5OxBqE7NCkp/WCeQYZatkQMkNCv8Y58n/D4gzKfzll2xR
Q5JbYUSvY7BuIcOZR+oCK0Xy6UunUJSBkK9yhxVdmzJ0AiUYaxyRxraWbolAhrB1MbbQ4/P/jDKi
FdkRHfhR58K98Xt1xI1IC9TsZLwL5+/AZMlmpnWzQou94osPuY3qpo2C0DxrFV83K8UZwG6QCdD7
HMsnvduzyD+XT7PEWjhghc/3ILlWQRc7yuOjRJNZLNHXGDWREEmvvIiENnFCyYRWSjRUT+pkSiLN
S1/T2GSn466dbrc2RasALB7/0yu6iuYH7FgkQUzEaf3ZbLnV+6ydWaXW4qAtMzZrxyEQph2O6LK2
RK4J7i994DXBRTnYzM4X//sL4fpyrR1wCvMBq5ZXqXcu617NpWLzWlbMhyKCKA5DjSDipJf/FK7z
+WCrXLE42ZDZaDfuIfJWXZELLX0j8PW7rxrrQ+96SqhA+9MJwkVTHMrBqWeGUE6o7rT8ha7YR/WL
6Sr3yCJ9fk7tM0WHT0cdVfXungJN6w8mN/qNKofWxKx2jCWp1Mur+zrEC+DP0k1D0pZeiJSvuWBo
9vjn6ZKAzVNgVVmYkA4JM+lHYj2zIo8/pmnFnleIjlyO9PdElIboiSfVHNLFvDc4xD4KNZ5y+QQs
A570omUy8Brse+TmOWTxbqwRW7Y7hspcoEwsOHH+1Hl8BU+VSyNylCXJBsZX2BIbW79x8Cftqzyy
3eH2rY0HgIRqN0jAyL5D7Yw009m3Z2Gfy0J7GexJwfIh+2ow6BXbcw0Yr3y36C0ZcGFiUeYtJMg8
xbE3OifHIqTkK0o7lzKZVosIqAE0SkM+Vzdl1NcwjwKFLPlPr4tDKNvytGYgtcv4rjaZt0yAIrt6
w/h+0KLfnMbLdVEkmK1v40gNsOd3Ad4A/FzLlP6W/yqu5yKzbav6jRFiNqPPmdTcehtD9QchAa7C
0h/TskJKUSYNMfFZopJVNH0sBgpkaL78EPczo365PooSkNnI6TG2A9DLKOPcjPRAo9te7MckMt58
EaHqSa+4k2M9XAxYArCCfAwof2Uu9qqR4CtHOSjtgSqMrjFy2IEpdAMlzm2ItpXjMnnXXd/F68XV
I54Tg8kp9EASA9o6z7TlTfpkv+HSge1bc9ArnqnLLnwMtDQf/GyNLlTJ+/MbpNhu6nQEevaHMs1t
8/eQGPcQx6hyRbHyn49PYNaBVpqu3iJq+sQhUZPZ1mEyK+Cj7X42OAAPNL2W8RTjgfMbuYOX2Pf+
XjfpNRbJamDKCnhqRx5KKmN2Iq+O4uqr9Qj0pK7RjYHubV60W1yYEnkjR1K0WYVswDZ/RWs2gpdt
X+y3ITJuOa1RaEmlq/Sh6wY2fF3N6S29vgIWZkvK0ZTE37rRJ56F8iBwVhalG1k77p2yPubx2urs
TKObk2YNpPP3mCdFafWf6UDuNII5WOm4CF70qj4MLTQDwGcqOwl/jmkhM6DvwbMvyNwA8YWW9wpI
t8ZaukyV3NhWksNu4+CV3OfFMHwzEnJLDPRvINDVDGZrsC9ROc+UR0RJwyFJ2iqYfUZUEPNI7g7m
up9Abhuh4i+UaHBnLT8a6Z9Bd2eGjYiA81k26V5MJ/SDcKX2MxbJyqcQNh5d6Lp+vae6M0BMF7O/
VoyNQsp+lT3m1nlXDWz6VYgocUThbv2sXbq2+0CTrscNgoeXW9SsHD7nqMq9ffjwVZXsJNpLE07T
SqVT9F+rkQ3SLcgk99TWqS6m6wUljSP7BjBHPRKzE9Knmep/yG7D5NR81fo9Ma4Cy/A3Q+JROZp9
PqMX102r3PMGn9YLF1GhTC0CW2rJG2rrH6E+AjTxOjSeHA1Bf1dt1b7C5UHDoumS6lWbPa8W1zRJ
S7duGGBMwc0ax7LJr/xe39whZMkFrw37UN61IynTfE6OlDcr2Yw3ixD8zWIHaxr21TVSPgYEbndR
qV7ZNo0q32tHKQ7UXTxuvMbzPYXHwrZ48O3HGPjnViDSWOY0zSJOyD2msw6fIeDhL/ILg2LFBXV9
fglrRUf0IaqVQ4uISWwSS8SkVNI7HeuMyFwUFNqKGpfnys2wuGFDvuMveQlZ3BeWXjeSTZ9ohezl
nnM7BLTjqC0B9CDBlRTrrt1rRjVnp4GDbnGZh4lmGW0IKe8mRaTc6QPvDv3J3BVplGLAPbjBnekc
YjD1Sv7Q/eMGv7OXe9XlX3z8OqbjIw31kPVicTMDqb49srxZDQc1bTZFeAHZrdIQ2lbeXfKtEe/V
l4x1KQv2Wlqo3Qf9DBO4L0LZr+eaQvAybjm/fGyH5+zNdZz1RN/S62xTKGoewbI5b3AbA+13RJJl
QEXHokcH9lv28hj4d9gQdKbe09QZ3HXoX8vrNqhaPa/TXi9Ux1O9p9rpNI82CIExEKlT5GRMGuEy
zDS296aqCXfmune0WJ84gsoh8DlZujeHIqUUEGTmM63zrPIPUZLTL1ocSW96x8Xfufmvh8XUfudz
9AWHgXPbdl8C64kldzcl9U7RuclwX8x61/8NGGfxp8B8/1GwVQQbhSjKheZlFmD9vwhpMrpxUQph
c5FK6vdRFHWf09SDTngQDuLbMkobkCGTx7Zj/Nl9k7l0Nf6TK5YKa5GTYZqiQOVMtq/SRvVPokEd
HYLWDQcxn3EL2p6iv3JOk7OVsTmJfnCxTpPTyVyy1EPZ1NyrXYWAd13cH5y9Slg0khd+BEDSt0nY
qYhYwBRB4gT5KM0wYfgJykf+5DpEKuVclYVJ56cfFJzRAt+aDER+ha+vBWTeCDGMJL5LUd5WY9GW
D685d4bRhCLawtAtD6IO/TA6tCNYDe9mZ8dx3FCxzZXhJq6fh1mVXIMpj9d7xG+e+2SqXFl17PFA
Gg2OBno+Um5GAUHjpjjtblz18wvj4m8sHoDiYdbKalfKqAkPW3DbyNg8U5J/MOPUXcCvSQm3bDuB
V7lCg6zSbD7QOC73uwyEdf+recMSdQW4V8QwSaQn6NYAzhEeb8wJmfGOvzriiK7mkVVFIe9qJ/sI
JzoLnDIVtJBTxF11BYV0WTyRBkrAuw7bmYr+n9XjFjFlcosRWntFF3V7WXUIJiLdkF0P8aa6wITp
r+rq0Udo+QTV+LYOJAVmJEQDhASNnVGIU5VYt3RhbHlY3GKiAouf8+5qiyD6MpYGWc52Hya0s3Bn
c1M74cfMZNQVtA3wYWVJVQ9PrWxqWM8Pl2e/DIoPL1fTbomYOhMlRjIVaU9mMKCWH8uD/tvI6J5U
JjCSQfsl+/Tl7JfEz7jRbs/LAHq8pPo1psr0HpSUx4YImkP240I6QN5iEObuvqMUs/BWGLFr3ans
+WDidH/j8QD0kDe5fQ5HYbAYm1oMC+3xGDm6HdkUR0TnyThhIQr9cs7xtnBD4OCx3ej8KW12EX0O
znZ/FNCoPrW+8efIumelMfUABtkNfnNic+IMvjpBaLrwIIBOW/RCbafh3eADaYL1C04CkFohapfL
5n+2IpDl0cUuU2DGdB6w9sWHSrEBNimwp2IrPMsrS85K41eac2sP6NgBgj7wJnEw+lsPLHIGNhua
NpTy/yfupAqL1r9TCYFa2Sw7aHBoFvsfp6AZeFJfJO5C22j/KcOqw73rziJmjFnBwL6dhVGHuAoT
RIaPM8SI+qV7kuYIqwSnxNvLlSDm/TvMOQUYcQ8k+8NqmcrUAaTyMcnRwldUi+qcHR4RRNYcfdxF
fogP4IVHNpw2Rj85EUhsfmEF9UfJMK4lCFLfdaqvHcaN3bj5rJbrcYaCTboHvpHELUckalxDmAbF
t/U9vY7oFi3Hh4JmJqhf5N3Y9brAwG2MofmUqpVneyXxvDMrcY0jU/YMCLq9O0xnbHHPMD+GsNjZ
hNtwk3iKeQzQPiMKB9/mgmF3hegUWVTS6ts0EXEbU0NCS6qbr9QtBHchAiQMR+M2G6pHi6YSbslh
WZ9PlqtkfXPZdRLzj7XqIGxH4X00vKn2DKPc4M4sBMLj/qo/cXvHXaIg2cTLwD6UWn06zoho6NbG
v0aAxOal0VxSBmS7JfVIoi9/OULGkgKXt04XQVAuiJyGz1+YUIHWZmJoppcFmxGrJgXOUjFhbVyV
7kjsTdIS1y7KWperrLxGjOIh7qInSlA/ZUUkAaMDleQu6VLCXrvQ4ALRMPctJJRasieQmNbdQCgx
eyuQJr7WSIGLnkk2T2IKTmIBRm9SimwQBkDgZbKDpWW/qtDR7XU0+KeDp7+QV1tyot1xQF1jKEXF
M46WSq8ARMEXcOiDxKBNYd/73F+fxJ9sIXl8XIzpQXKUpbHnwlkwRawWRMLQapoikFS6pUN75Chn
RfOe4fD9Th/ej+58JnDgSen3WrCwKfAlugzs/nFwuL5VPj6m8HPTuIDFn+WZDYUgPJmMpGmWb+A8
w62edwIgQFTD32HRwCAC5LQSolAOmeLSN1faQNhA5Zh9WujTaWof1L59tkurP/i7fbP1lKLth4VX
i72T7AvTghjByFXnq53zx1F+MOkmVXoybCl4tKukrnuQRsXmxVwPLcAURab/8zq2hDFApecOE0Gk
1ZEPl1j519mRfn83tWXFuSA9Zg0rVIJJ970YuJp+wm5qrcOPTFVMdWg58/RP098ow0vj5L3thK6K
1all4jb2H60Io9wEHDdM2scjgmyhFxDvyyy69g1wg8OmR5pFmhX6GgdW2NKbxT3F81mGfX/mU+fr
S9C76hwQhf0EqA/ts9RqIWtimfHNONqm0Uy6b6n6ueotpO40ySA9qSHSecXt+MaS3vyBUGjxgkfb
Lbdr0A6Ln+jZuII1UWH22kO0/a9/c+QgWvmy5lFwu0/dShLcJgJv8y4yNIOf0sPCNupqHUGMz7Jc
Afz7f+X9kLNiM+MEBiqNQnvPQHba2JvAllahZgiZqWjnjDFHj+az2pW2jWjloT+6ESbpk+Ajjb4s
iKlBgifxlJYg82jOZeqetkwihBGdkp/6LAPu1+Snmt+Epi/IHWKRtRIliNNczr0g7SMKIKSmiO3I
6/AR03FPhiCtGfGQUsoGzjY4n1jHx1CxA0kxruusLkyNhNXw8CYr6PSIhNY0Ezz7fsgS6UvnQsxN
Vv+N6KdmuP+bjLyVVSiEnJl2GN6aEJykLDQjCjzVmonTuK38yYgvfJ+PNxnUIzI5z94mlgYp2DYb
FlH6aiFOPcoFMiRGeI5BbVWVkc8qZ3YfW5aRg6P0OSlyH9WOxmEBjws+Yo7nKTt/gbU0tRnl71wK
E9Yc27XUHfxE1rwfHDGsMJdhvntSdj8tgrFyrnX7b16i1njlMTUPdfMZrhWxQQLzjhNa7I36C1Io
LIX9vj1mrLO33vljNPGywQK1qPZVHhnjAVfbnCL5Lw87zDhlCZKZd+HZClcCDQFWs6S8mq/RPOuY
iDi49S/PfUHdPp7fXjpIWe2LhK/REU7X6IDF4RNM75lnfUNqjxRaJpFa/ss/iRbLYBmdtubNtxcB
87sdDTlw+0K2btGj0Yq5moX8Uy19edd0aXIz2flqB2Df1o7xcAQFNSu7JRFsiA7htagsIikY1dY0
/s752aCUMeqkeHXRPHWCL6B4JS07M527hVptvAfx8YLV+MYP+60/mLt1SD1Su+Jznq/M3Gvx+22L
89xC/BPh+LIPk2cadHlCNVfEpyfS9pgiVE2GWYHS0jxdq/GIAhe/n3RY4F/qCrrkyqQyiOmjvthB
brGqRtn+Ub7mCM6EUbl+dNy4S1nGLA3Ezd+EtGj77vqAqTw+7WjrDHxRXRUl2j0oa7LMZR1HIulg
2Q+zkbc8UXgManYcbxICBd9v5eQblOdoPCDzjbzupIUDpF3kGWJ4Ek4gFM554svP0O+HLQiGx+p0
6Ywb0uTkCSQYTF/nsC4H1WuPR9sKALoXzSmek6ih/ufgCzRVhMezdRasPJ5FpQDmixHcNLNvB6b5
RZvE/cV5jFiqYmy1BX/Tjyqd9km1uRa81T3dvBgKffqfNLFDfE+zsZyVeUczCQoStMr85trxchs6
UmY5vemLwxOGS8POXJ2sYRxN+iraDXwxL0kVeWkeLeGxV6Qo+r2wE4c/aLP/0Su2CiiCf34YUwHK
lb3k4WG0TpeVvRUuKU/VF/NLtucCMdPP9RYW1jmIq2p0tivz2ezoRSPtjPsI4Q5X/bvD2I2oprmq
qZCXzkC8CkusX0pJGmcaeiX6wLPVVDWwCZNhcYxUEZLk4L5CPegt8a7tLr/MTnYmOkthnLAuwBpq
UkfW3wFygpw1162BmNgdXyalCJgXC3mJ7fVuo6I0FNfdStH11DX3mqQfO7neBn2j3BTR8nGF8gGT
VTDj8Iq6HwDEr2ZSx/UoKRWHmgtqsafWEhQmkkBonX7pW1kcyrnNINr4LteKw75BD2+MN7E6/Pw7
BaIhU/Cv/n2mol/mno7iYu21u/6l9Ie+wENO6R3TDrHzJZbEzmJYE13pawAPJ6hWCx2fjaZ7rGib
oNsR1xufAYkXJ1KpuWU/HtytLk64+68H9xgzMw85YvrfQ9hj243SANV5U3D25PP1xCM1ixBKK61n
MN/T7BP1yFVjJa7v0l54mzfUjp9htyz40uwsXG6fzaqnNujPV3qt2Kc387VXbZ/WoHSUDJdD9SJN
sLGVr0vnIFRz242XhMKYhJSpC16hTkCTxAaeqDLltb57MgACBynDTykbji8hN/utONjujvpPJIg/
inc1MxgtmplYWfs0zALpQ9ZdqhbHq/t48vd6yIV2rAzUkqwku8EoMhP7ORill+fDDc6KllH+iQMd
W38RUCACFHhyDOet4967nGFtZJK1kZxVZMuXmzA4H5Cs/DViw4mW3SeBHkVNFVrvUzcj+eHmeAHx
uYTgz3wApJ2qHhquHQYyu4qk1yEFsDrAw8pCKF6s9pZSz/p3pomTjdw8jsQ8Sri8MtNGWhO6Rjmg
d6vW4E6EpfsL5bz5BaAkB2YkBhEgf1p+37Gg2BVsANqcY9bWBih2Xu6ko8u9y3n9P6oPHGBldscc
SQI6jjfOUJcJXBeHS/i2xuGGzpAKZdwxCfRi7t1soyDFN9OvEsxCfiQ/HOniiAJundCGVJcj63+I
d74Rm8ySB4jTHzJMu8mMxcf2VpuuUxjE3TaxB2IiALNZC2zVeRx+NxamS2g0tTmG7qjRL3YErJ5z
JdBU+2enEyQWmAkr1Xob9Kqcv9ERH5y160L2NNFSCcOmaEGE3vGiI265VRRMrhvUh0h8UV9uHa2F
gBYt+cA6WksrAKrU2AAr/jkNJMZ4sugcO4zCdVKkRpIXq/0rbNifOrkbSwBkEeHBEu0AQLLYK/bc
+35BkE4TuEck39aOXFMQB4UX9nDfuX6STxhIWcXWjmUG1kpl1Q/pr0H5mjvILEPpi4rdFoKnVH86
xObTNjxhYJ7Vj08KydOqxcOQZ6EgcqsQh2calHNHSY5+tVRT6hRpSfrvkEoKjG0egNyEO5L9S5rj
w1yK6yMdO1VPPNVCR9m48A79Ng6yqKB/oJC708hkHw8qOTg/BPjlMxpp4uniHSyakVYXzDa3Iw9b
F9g56x39cpJefxerBQFbcsS2M9kksHAh03XxF18Skkwptcv10YJlsdUmeyo475jrV/XmGNqBeSch
Trq4EJ+7YrkKUPqO27UgHQGuN/cp9HCqHW2ilRuBsKKswBJQDLpzSDsXo0z5JnnwCnv3IrAycjaP
p6GdkYtg1Z8NqB3s8sLX4CxkVv5L4WDWPMM7Th2tQUyb1elqxXyaSAlr4WbKSanmiEC7Qonq3vRX
zh1BrIChA05xZWKdLbIVKngtGaFu2/tv8WJS6qr82b3+JLrU83d6icKS1wRABNDwb7BVEj/al3Ev
UPEOPlz14QOSLrE2E1oY6yCoOGpuMDtmDlQa5V6j8yhdI6pGyBXzYqdcTeC3iaaOkkf+mRcNPyJR
fNbyQs24fga9cKDPiacG9sSNBi7+ARh7yUGwSuS5ccFDo4a8FBS589LMc9Lkoy16Hz03pzbC6d3S
qzKZjwWjnqeheXKL6AIRVJLQMKkvoxMq2YG0WAPtBfJVOYBJ3OKwWzWJ4GqOJZjkst2/DKBF5wSN
2iIfKrPBQZTMeSSbWd2wrrau0QzVFcY1uwxCIS5gXDCd1JeMD02St6DQpG3HpqfcsPOcNulWJz1m
uj3UAI0HkeAb2yOBczPJFaefZbwrAxzWAAA8DV8brs359mdjE8c7924Su1kadCv1BJ3oNwiVG9M+
TKOXwmk9YQnBz3B9cZPKM73eLow8Ec2kZ8w7OoUxEuYEWxVcUPxSSQbbrLZsln4R9G5P7e5jW8XC
YxbrOXEkVxysXC343haHfJyCXTUHqJXkxaO/OLe4Hd1veXuXx+nzdL3/cPDlLnpQFb+Kun4BrOq/
/Hy8dk0OBJF2zL7kWBaKTiZ6PbLPiFdWXuPoQ8Mda4pNi1WYqAYsyC3D1jsLeNAkZFWbKZhvo0TE
bRELpgGHwqnMIh5dF/Y3w1byYLTBNNEgF7KcrPfvuDldFgvRi/CvFx9zruA20u7Blr+k7pW1EyvM
MRLkgmwE1pKyY33JjnOiXnDtz5556I75+LKeWXn7nR+aianasvPL6l5DbY7h/nD8ouTY7Ya1bPOv
UYu25MwOMOJ1O8NZXizGKploUq9eTlEQZPght4suNDWG2W4V/kCawVIxEHBsqE/NINzTkiXdFYuz
yVQwfCK1/br3O7/DT20oQ2r0p/lUXc+cHyeXscjKP2DpnyNML1wYWJDXUuQ0haqjNM1/gtKlT0q+
cWYskAqjYCdAfy8O0o10zrnA3h4e6GLBsB/Mzlo069LZXbebE++T3D1DoVsXJv+R2J35jJKxokAk
5F/jfjYnA/hQusrA3kOQ/S2Z/GfIq2bzLObf10QobuYWA4i5/nScKWM5IdwXfRZVaPVigPQa8m8X
C6SQXktg0MY5G4o8ZIUpZaJw3xh42hMqDpZnUb17+3BUdmhEf9chGCkvf+kxpKnR80e0+EoksZU4
5fVu4ZPMUGD9cVQXaPLJpOt8pN1Yyp3wZXKES1mA/8D3wCAn8lBPOjYA6kG4NOqfQGV3iajTKOQw
NpR7jDlrKxIZkqirda/FbjEdRtjIl3Dz2A08MfcwwhCCNqkrWLJ5fox1KtS2p5b6mDjF8noAJC3K
7fTQSZTJ8iSjMcQwifmxsUKRWsademfrXelpWuSqOJ4Cllj8ziZzCiZG4Bb5BW6ommCZEiuUjgqC
Pj4zmVQ3Myl6IL+cFFkXXyYskn7NKaf0+1W3nOTytH7glXQmIwvGIdvPGaR+EeSofPXAa53Sgu7b
LXgQ4BbpMr9xE1VSjyVXM/id7Q+nwP4dGkjsbd/vLw1onThVczOebrN+DMe8f15VoMIoKX34ee56
g+A+hIHO8oUr2kWAJDJsMDlFSXnmxhJ+xV1Ie1OUodcd5144efkENAruHB41m494CxXCWWE2Gz4s
/OI1lIVSqTxM75ZXVNN2924oTGTxrnnx/RfhcdEBkrtOl9B/zmpzW/ixdQ8Z4pnE6C/RSoeI0ZtP
G12IKVGjsnaXPpegTBR1oyi+7/a44RIZGi4Kho7Dz7wK0ti0RoAD+cVJwhmdFwUdnaw6pwEK19FI
P9qX33GjWWp6QP3GfIN3ZmKrFWKrzb1AM8FGnQtZlYFOMjXqnVO6SAMCoKg+Et5Oymjkl43rIoPd
FVeKtm4WzzNMvB6S7BaLjx1Vw1Ey6HhcCRz4ES0jXBRU6a6ikFf+zIqGE/sy1GdYV3ImI6OvOiUa
7u48cj8hnUR/dRPFjEN4jzd+OCna3JU66ZsGh0ahSK8bFwrvzL8czTVfpGbxJPlpcKTSoXxLjeFc
85P9tM/dZEmH3CgOFAAfgwP81YKkyMwrAuWptz1ifdQaWoNOGF8C+b7fM/Fz7WrWa1SvbC6Wq/wM
34BSc4Of3gKQVI7tbQz3WljG1Hj+n+3bPMZgo92F+wNXJGHUFl9IyWJ8UImhTxTgr/QHPLJvXX+G
utmp6PXyjRPGNl/0xJndCkZDLx/hmAD9gCg5CIUbeXnSS7Xpon4J4MeEbWcexpatF/4/zwLtEy9T
ts/wDt0vk2mHLSiOKkNe8JLpzM0nkYQsSwmX/UigbeaNGuuvlgRiWtDS0enkrNgWnhZu9H+lretg
EGtyM1I8AmV3t99zoGsNYwuO20LepHBRoV3SjZCZWUKlnbSQ0D4N4zBjmkOhPR9BE/VV3LDuo2sE
dZz8RVDzgB2sYcUJDjd5LAMc7DB1C+xRFji5lUuA/YDaaPnNmepkyXAH+meSfB0eUAoy9WhEN18Y
0Hec7kHGAi5QVG7oACvNp/95zBPQvPock85YUBf1Kyrpnwc8NOefwXEEHKtQ4gAWEKmLn+Vh15tz
bgLqB93+VohwChGUUUVilNO02FyYJYWp4IzbeNtbJ29wwnEQJF6Q/PXas/J+ZrhnG4JfyyRx212u
7HKvlUCdxb94PsEURWy02FHzdkp0aZlDz0LJ9t/L5evnbgrId7p2gmk3FQNskXU3IfU9YJRwgQBV
6agmTHnTYDGw5S3eCqeoS+3G4tkUh4fVPvOvUOjf5il79ZS1Xi+VaBVKftsg66ctmzc3OZgqZ92k
BbTzpn2GSdURZNbXLd3kwuqFPSeO8t5LkOXADaQLhuLlfXPbHrtyuZEaLZggDFtZsdUfCFwm7V0x
I8JFD3SeoDWG8I2gFn1PgOvxD7becUu4R7lrveI6VJNd6QgN7gUWyTF3ONXbZe2oLbpJe3HVyy2B
/Oc/Qo7XFIl+4NEaudKwaNg9iaVhW/B/5WkYX3tvZd3T5psVFJgk23RysxoszASgKl6BU8+0OZ/2
CopPQQIUJ3VLySw55swan44YChorRW204XJ8GZYHl8cwc2XYBeVnfTEfdMGrrar5EuYNdbIf37OG
Z2uPwG454nMXQkD7xEfbXT1JscMDHnRXw1aO4G5Lp0hHSwgGdUJk6w+PbPQA6mz6qW6MKOY+5apB
jnl3xLcfMW0nFjJeiE14OfBQ4r4nDjS6dItTizzJZN34iouwwNeCc7EALoyKn6XH+Y7owzY95o7U
oxA/ZiLETaX7dRLwflbBTdGuO5HtjLNZF7Py1W8xbHF7eyBzmAP4kMQtdxDTRPXv2Z140c+kr4qZ
kXni0f1yPfBoZxXWCHMoYIvKIAibegals9kzpT/7M63KhYdI3zZ3nqQGHI9Jha6tTnEVb1ci2ZOZ
aSX5CTLPY5tKB3uKN1b9/QEthp6fawJ7wgX2b5MWhyu7OsmK2bP3lQGINqPXnV+UaYSMr4zi5Jh+
jCfN59UNOQk1MWFUN7m03kU2sHowxXNND7sWWxv5oeMSoo1SQg9v253zue9UE96mY9/HvSiGw/Fw
wDW+Hf35lGMf+vABbW6FKf2knT5vv4uz1R2O47Zr3GXM4bBmTQrww3nhn8266T8msPsJ/KpxhMJj
J2oHBqrqfoqLvsyD6gxHFy+EggeyU1CdjMHw0i5S7CSCtZQCDc6yhYXBCj4XJKOhoLwh3Gpgn5SQ
IH8ICd2wF19uUiqxUvWP3kmWuCsNo3Opdueqhk/5zbHOI4lVFiO3ufUhb4XAaX8DMIIJLfLQX/ZR
9uLBrEjxJNiLjOX9UGREj6Oj7SXR+YIzGw0/ZfnHQvyI6TGX0ggmJCowcJidT9/Ay+I32m8yEsKZ
9IniYUj1ZNhVi7Q2fIU5lBJohM7b9T+eyFH0DteL6rloWSmMAzYwak0nJ4HN0vhk3lFCDcwj0vzv
fLM2L1jIfOURQibACZ63KQSy9NIFwMsgOdGoAzokv1VEbHFfpfo/wK1+gNnJZbtSTY+L+gqerK49
nKp+ZXdSWh6OQETXRduRqGw8GauS3Y1HKqf0xeRwukvy3Hh3kwLhglD1YQ/eqQbu3TtM4TGhoytL
Y4tM1bXj1vRBBO3Vykb7Jh+mcYIU9Eh4RKytrp5YIX0TGRpvPupGVk5UGvDJ8F69KZ9OsX0aWmXC
ZOI2N3gH8y4L/YBPHJiqdpzsEfdYy+b88dQxpcXHqZoHRfCsgYgv53iBvlIJxCcP7DPzykiNbk+0
NpqK/wEw/B+1lOUpoRnsjSx5+hHh49xByax0nswH8s0bMWByaquQbsEN0LnUo/maQjadt9EwOjN/
+9zAyWchrVSmjfO2tMK2PGv9H8QMMXSYb1aUIANWxTavf+ZSWtOGNUuiIwipud5lXfrH+suuWtmd
WJUVoVFsLY9Hb3OmlHvc2xCvexQ4ILzTYyJ1T+tTGaTk7Nsq4i9nftn56doyn9Eex1dSeas3rDiS
aRZT4DK9tN4yFhYYiVIS8/LGH4P1mpy9mCAZ1Rdk5OisPItQa4ZmfObEfaFP7CbCQtX9DrPexacL
r9IfacwM1TK6nVz3c5XCsZYVyXogJUUzbWoT6uH5M/34R0jLMKz61Xc1mO9Ve6sweZcBXlXtwOGB
b2pCOMucEwUx8hHyQcjVA0p6HXvp8mshlVzhBN7Jtn/nq2051CAITk9BikxzqSIHF7vkjc4NFAl0
BEkZ5qwLnSGbgK4TU6g0cadcC1zmwNC6LGJR/fMLrsexK1Twk8VzmCUbLg7boQ8JeseZo4LBPvwQ
AgyBxJ/JwH0GIyUsMKXBg+4pxsC1RP/DUCMjrF4MCLluLI+HMT+8LagGDAJYBIlBm4nu0fp1S1ek
xRlphwaXXBeNcCVinJQD59xKO9R5qLbQ9e8mC773Gf8StVxp2ZBMYaQcGt5WQfCeQ4LYKJX8UJ6x
fRIhzRGZNx7WPFmss4PR36lUk8awKbp+oUvCiAxhA+Rz++nneqRwldXfJUEHRBtsV3WMdUi65mR5
Xr9I3bxO+mo0gp8+OrMV2zbTrr4Hn0Ob5HURkhPIa0UqUTOyeJG9aEXRPERp0JBRZ4Y/8+Hs8Jwv
yMW3fKHaSS+QYGxZrsXYFmr1C+yLn2g93Brgp0B+VQeJTU6khDPXK37wnWD3rjQNegdLjFGfWFsu
2Q5HxbjfTctdnUANDdgZ8VVUA/DFEi3F1vB97baR1/EBbo30jzofE1F8o3L8UYnYW82XfiLC9W/o
n1Sq1F4WUDY08tFr3MKf1oQvqbcCrL5ByoeY2l2DN+SHet7Ed4jCHA+qIPJpVGVNBzVTb7SY/GbI
xd6KBkhsZ7ndvwP7MulRdiAwKhx8I+VS1OJcvJLnIsg+2c5EcKP6kUBId/QDQEGs1cSc2+oFY1Ek
827tbAMixD/1ospNvppyqzCumJI+38Gxl9j8cF7WEWRc67biRKB7009uBlKMnvsueiDxRcefh+Ox
gJi5wiOjUAXQf0WstGQfxvn6hX05owB12wNrV8CIw8MraXyFrxlnfTLXAfEbrxzR2jZJ7cqK9P+s
/2T/tazF7S5iAPhUN8rz0Xd8IKusEnjHzyhPE7kWgMhWzW5GP/Hz/AVCFRuK+W8ZZyZSOg/YMSeN
vfIX+kovIpMGzKAmfQ7IyTto3h7+si86PqcZ+Q154cWVrRKmkjZincu3ao/oovkhahSPj4nwO+i/
eQPwViY8VtO+PDkDdN4fe5TmX5/vjQ4DDtVNvmubDorS3Qpskn7+9xG7dIsJtZbzLIdHcbxbi0pF
ic7jU9ce4Ii+Km4RVDpOHWK0v66JcshyiPvYgbbwOUgJSee6DkqIrD3JsictnDgPh7TOqQGGu07L
G/EO3NpzAkVRIq82DosNpzJpoAWSt5FXy7BJcdknBo8Uczw5LJlOjqS9gzmHmdZD9+TUjR7jRicL
sCk4RLhD50XwdrwdfC7b2HjvM0dtweYCQtyTXTipTDFUYMgAmTRZ8W1gAMTONTimmeQ9SBizKM09
TZUShB/yxaIIRWDTKWNojIPwRVEIhesezuNGRC9/YZeuKQjqqa2xSRat10QELJ5t4EyGfEwdfXs3
xhMCUyraIwFkgda/oBYTN4GfQjqckCVix+8HD9tgMw6AFI8jMppgDVIoIvC38fuSbQkBzdIlnnBv
P4gLtA6AQ7UGoQyjgQHRz5hJItGmiG+LUdxerWOptzsB8SvFB9dOtZ7K0Xg8V/pcj3gThQRd7xe6
a6U20st2og3TfYvBRIvgWgCZSj/g0QgmVLjdZQhhFoufKTkzeIU8WtaqiBmpe8sK71cFIreZ7rk0
wf/0m5yynd4P7wXbYsK0wIPPaYhu2UdjlUtx1Bs+FS25f9zHNQuqV2gChjwp95lcSqiN0QIZ/I9D
D1V9d2RGEqFrTJPGIKA/lEZhsfRxnlM/YrOJA+4W0rHCHcICsygD8jAJciA5HLY+zRo6wNSY0DnN
6Npm/L4hf/2x/jCsC/UBEmVGp1DmY7BhoAuvmnsTWANf29JjOLaaluDavFUVhsIUPQZztQvy3iJx
KA6k/iPl3s/VZ7DmXFkp1NrrEEfrl4yKxCoc3JpY6fS3FswoUcoYjkJ0rClXmjJ4GY2U4bEfZTH8
ubpFULIz73id/O7nMp9WOz13MAP2+yw2I+BPx9SRt5EvJjaf3rbEGZFP16P358Y9+BGym0A7euiD
L5g3nqUYlUeFVAC/FT3UtzKMPKhdwi43tzoVoSrL6l+XGOL497HG4Fd7kkQAyUkfJB08O04F1n42
9/JIdc1CCXBrTytp+9w0XaSsmukxM22cauvk4qD6xKTqyQYgeM2/oJOFom8QRlUnsSuyVso2LS1l
lToSLlgmalSv8GYTqRmclQcgoaSTOpQtYvWQXQYsYb4RYpitI90yAHCcWrUxvU1ghR+5s/h9AoqZ
ePIkUEXIYPH7SuS1P1vikDIkVL8x9KEk3+WjtWvGX5hNaEyI06GHzE+SlsTkhl4xrlYPeN74NbNI
vHAz1ZYAac6EWecf10DZk6+1ua8Iyk2FMofuqu3hJD52Bd0EHehKqMtABU+G2tphexPiD4s3cX25
Hj+z17ie/W3QUcXR4mXFPBifxfqx2ZPjzDlShNoMw8OzFHtmV8cu8DYGorweSrh/wVNbGKE7EDOu
S6klUsYO5GkyHCkpQMFzgcYIZlWuI295oHAmF46TCKLCY6BZI6g19OKP0+4c+JFM6l95JlXVgfYJ
qSTvw/P9UHj/OdEepuezaUbUrYpARva2QuQUncCHFNaTh40f848E+NuWT5v7H8+qb8iPGA3ZEFpu
ynJ5AsQcAZN8bS7eJ5jTSKZRgIm9Uuvzq+jAZagsshrfnVuJ49ZyG3eA4f/oQdNbZySre//EytJQ
OnphtcAiv3j9om4GJAtU6z49jNjgH5Oe8JlxJO9FQJklbRMm60HOlAskVgw0BdvNOLsnS8kYM6/d
AW5C/uYyoIB1ZI7DKRbqOS0QKB5fCB3G7JWEqK0QTaseX0RFrqTLFuaSC5i3d5hIxdv4mmgbG/am
nAYo6WawmMHNHVFS9b1gIJq+rkpxfhP+HfNbFRmuvbJkwS3b+HsdAHkM7cLPN5wPhl5wdswx6Dis
sKnEZASBCSnMPpJ7VGh3vAtHaqfJKF+Y9n+isikHHOCL0OooBwzfihkpRKJaqTVsL8AytvzYDYky
JziW3h2kDHFWl5MA8V71aNXFQPFZkmOC2HWCYZG+GNJlLrGrU9nsUppuPppt/pl9LEEWLs4YUy7w
+ro+XOHY5oo+eFHjg21z92K27KoeDptpUe4Q4R5qf6I3g/lyFQwRB8IShhRyxcB6snGooiOIYu/V
wJwFthch3R8MDBZEDOJi/XNFOsg6NGmg8Tw6SR0W3Nx63Rm0dD6CIxL6Sgs1LlWQLM19V29yn29F
w7anYP0DbtAKcX0AD2fGXSdfWkLlN7oE2QWY5CGa9BE/P4edThcY678800LVITGGNiDwqQY7CWKM
TFIsDiofO/Sbb/mc5Ytho2nQ0l7fViBS9D1QOGGlwTkEwQQH5OOtW36jVM7/M1GIzsvI0qv1ccu3
y+D5UrXm4X0Ei+x/bEzZOA5bmsXgn94mM2dzjNfaVCLESpiXx5e+Dw2XpxBNcLPQqSEfx57s10Xa
1bqRjxkwppMPS3GZgC9kst+hqXVNFq1IaeYg2GM+c11fClqHZ9Z1LbZTjNkFKZaoQyUIjwcWwzeM
whJ+N9gE1JK1OsLu4+4gX2sfTqixlVdPKZEMduqsu9zNEEg1nmLAAkP35hGNyzznHNKP3GhyDgLt
mmmmw5ZIpiMKXhC7GQWKr3sB0eXkqkz9h/wVeJSAItw9f8YhuWEPpgLLyLcgwBRTjQcu9XGwNojn
x/VpOm13Lc8jz3cWWTX5sw7rJW65oc5nyIeeV8ev1SVfmrrj5weSVwqjl1cb+xe8Omq80KtUXMJ7
e7aiUcs3jLN4D8P4gzZxNCkhK1IGasrKf5ZHqnHXYpP3WFmlLWK8mGREDswnbgNSywJyRaa20iUl
PtOcUBM6J4AL73lFfYiXTNrklwskhLRVgiAQRy9RmUkds3MhBfCqVvhRDdTiOaHo4qijTv/ICHhV
o43gbxxnhIf1qGcYRfyt3uNKQ7RvZdGKWa7QulDyk32o+RByssaUH0shtnLj3UTb3HVr98xAW1O8
+PFD44tGlgM8u2+mJoRZRT+WUaenxIHnRKiqjzJZiCBn57MhWT8EKU9dfPxCliCHsMFXzqrjMKvB
vnss4p1Lone21lJuDQkC5NjXI6ijQ2kBwPalLDd4o6/J/O4PSNYL8oCmamI+PlvCcBVWYDjvvbjg
DU/s7TdRXuasmkyumydyYV9k0SQ3kDLSsXMYGNMxRZtFoFtyZZHv82NIE0lb49PT6IzHM4Acdj2j
ZxZXv0hF1SnaHtI8Xf7waszB5lwDhU7kGAmSfhyF/1/rsC+6/tYCIaHSeN2ENQuUQbthhtHTB851
CaQGF9C6RBhYrrlDjhLRMNmvOAB4ZXeSvfQ9LIpgaTjN7DlMkzIiBTzk8+od/HkUSokWjftoJggk
jPrIdgOII217Hv3Ych3ZuDLFBDlKuWrtJwxoIM+p9okvAKf4P3wfqwueQBi1GMhrs5iNTz9IKf5o
+CPX6aClGSrt3kMBbVSmXDdcxez+NXSVwOQtE9wgEBVkf01ciP8MV27achuriOTyuFw7ablvmhBB
ao2VkxFk3UMgh9MjV28GpxarfhtDEQuSVUL3aUNBwED4jcDiBTNpiEXmkdon4zRsXb2v2jjSOQi/
GtPtH6bOEE2K4jKeeKv26aV84Y9IOO3Oi0Fhx3Qh5GT0OH0M29Q5Y4TUPYuzGkfEgDf3MgIc4t6g
S6zrjzb3ROEp6w7iH7wImxdRYhhwo4fCUdXV4lmib6EwokljpPk6mp2ya/ALNIiXXQMoHYgLXPCp
iziUef1FoxIqN24mmuJB7uA1NMsorwzs/qh8f7RiXUUvRxj4/Yi/5zicZ99mBjprxbBjbtkHs1N1
QlruCS18nPO2kfGHIrj2Dwz0xQrd1+BZnozUI9n5g4CTrCScflM8V7dB7VMDtkOLgl96cuH/XGBM
DCTlsrFLOh12ubWlQWuW6uZkaZc2w8YVmLmFvy99kRc7b9OKMWiigM0e9iAvvmZhSIWCEGrXyQs6
rt+VKj4BBE3GMr5fk3lXC6SY+iS9TZdwJwfws9kOENnFKDy2kmBHprY+1TbIbAxyLdyUQNGqNP6m
M9zZwyBh/0CxBuIkNKQ9ErdLzB2uCiQqg/YttzwVANFnyuTrJHtvuZnI97MmQdm8V0h28oo9ssqt
Ri5mETqcVFkSZWMNMvsDC7OtxU69xA+m4PkfmIUIRLrGm084M9EZ21RldW/igxn611jUD+oBkH3J
smEVHVT5D8WhXeArZVFWefUS5IboYNlTpsLZnoaulFofsWtPKRMDgs+lGoGpDsoa+ttQQVAYyZWD
LG9v7oDJqlKQJ3zXLzstLPwzINfZYrNI1poTRQNn61P3cdoqiGjcHUO/lhxiSoJYvbiZlQosJSlO
tjgSpN2wQ98Ekqz9245WK9ucAqMiau/X5tC9pn868bzuXcADrzgdAcgHq+mqdDzRGq7mON5kDebE
vHGD8oCAy8C/dLHMkectyu+1bTBsWNjE62UcMukrwK7UFgdmkK39bebNFKOyjteMjV+ZnQ7+nyHQ
XW5CF8bnaAqjGDXFpHuRjalXY4KPZIZiPB7TiQZxQz83x0i09pur87AWiX/ubItfyq9Y/kX6ss3G
GqsW0s/Ptb+JZ36HPgBomFWuW1dLnG6cUc+UifL+wZurGJjy51gYtdt81FLY7XyMSJqJU59hy4OT
mx58k3E1d/hA01QVut68RSZ80CECNLRRCzJkRobt+pFWxwEETwPXJyQN45rH7T20B0wRSOUhdDHr
/Oc4Bn55BvmMdCMnb54UvJMD1tbMZJeYjxfBOrMzRtVUUHSD6GXP00WrGVGvhWzZ6ktE1kp6AJ3t
nUMWUbW1nxl6N+TkCOMr+5OmTyQehODOxg2LWictcE+zXZL57AaOYwcAnu3yNU+LdW1kGpD1nohV
lsP+tsDd+WPzP2F4sM0daaak/Q+Sc5Oenhvr3FjwE2aDLBRG/qf+hNapnlbfsZ3L89lMU4mtou9j
Ftzm+NJ4ETd4wtcKx2TvUcrTMNzsmPFYehpNZT2fgN/wKXX8VEitYexfgZJ0/WDuRZ0e2aIRYGzd
Mwa0Jya346fW/VjzWInbAEqiv5P4CQtWEnYG52fQ3MC3QRz00foAHhMhAZ4UwH4/2TRG0eXR1JGB
tLqHcd+DtYGzyyRi13ORESRcpStsFwEn73m1EE8U4HA4hJSJhgvBl8Ghxsm1xSV4fmGuWBWADhQg
g3SB3hU+zL6RYJMCIJUGa5f5KvaQFiDm0PA2hyHbNDjqZTtOghzuZ5pqqBVJsCPh1bm9/JS4icxI
2RdU+6Vm3dHB3iIuk9+GIQIY0NIyTGubfmFCccuI8m9yAjLUBrRQEtJ3kuCxZ5pXfOzRjK3ApmNE
KuKTCLBbB0teIKe+RezCkO39KgRJR+o8A/y6YKIfnZOi/Lse+yC6MS/8PwzoZ2nzzeDFV+vA26k1
bnp+ADLTQVSzH2OXwVqjrBbgxllXXzLrkuokMRA8Aa+ScGSNr8Jf8la7TpfAPuvC3ZzFyLtdN1y+
x0tKdBHyeNIF7K4lpOtyZ23M8JwYSGxsxBOQuS0F4g5jOiSlF1zhZpO+7sdu2I/eSx8rBpcKFcTO
WGTbgRbvwZJOWsPmWcW9J+Hbwy9YO9G3jlxY7Ne6xkNOP6fE522FpCcIhGZstzj+d/jYgXu0V2zL
s//yFMkGyY5N84W72Wc3UyQXZTQyGPHYyG09wNHucKuOEFEAhnNZOtcGNDpDRpPcHijjwnWe5XN+
YgMP+QgmI+ErBCHHVB3xlbU5lRhdIfJJguSCByhZturgk40l4NlLRLBQ3WwwCuAXQc83Box4sQ5f
zzo2AbmoKqwhmh07tlhfXs8BgukybVlEvf1rY6EVm/zyq4/qWN1nNVBCh0udlZGlR1+h5BGUHL3D
8la+tym4Usq80sKt9+lWXwcDI9028CE8jIga+nrL6qRcpMTrmqsWgc+EBy2xC3Qu/8LDqYIi+PsF
HcFdFtbYi55zxJUvXmgwS7lk5lN9rLpjfEJ+srh5eDLqO1vv8V8Kw5sdE+g3hAG24pYFqMwIyu+c
8fsn2mws5b68ZrM75+u6OwqUOO7DbWMhyjnSsTKatPvvxhEl9Q71MRlIqw+2Rw4BAxkYui6KXcNs
9mwluzbDI/S+7ftaWBFADyKnPc1kTkkJ5RDyyAKIbfqDqiBBSXMJ2u7/q/3M++RNf76nm7hmF4nJ
VEMiSjS35sb1uWCV2+f8SiW/5Gp590pov553WB7K33OkX7CJN0AKNHxh/r23YFRpyd/M9R8tOdzZ
88oI9lze6qv4jAxsht+tD3mgQ6IvbH1WgDOEUiHhAnyW4eaL1Y/eulVpsM3ztEFkFoZSvEQYX9wT
7CKy/dVJ4KeSv/nfD22hl/M0XCBjSYm0i1dmj09N7ZiJB4uE6N/Ke5BKzc8VGInt4xac6+UXcSiK
MDJgKxmV0pYa/joFD7NVzQD+zCJVxHq3ALcZD2zuP2fVoBycUF84ozNqRtQL75dAv5nCIGFpRtO0
BsOGEyrkjfjh/ArvRR6yhPVksDBBpWlbTNrt8AuW68TkaDqXdCqEoso9XWrBYziTF9Er5eCxcZu0
g6zutVuiMNygWNkPaW4VWmYzHZErxWyJmg93VipQ9hcIAviyt45YQaetY7qBhvK5mS9Yhn2TTDvG
qtm8gRdCmiA2nPXHPpXPynn/LlCyRRyiycnn8TWzx1IRmJI4uwdH+eJ/TOQDf3Vk8R+ZbN4dKleb
8lVgT6kyY6ROUt+qW9zDpZz3zjFh/H9GhQNuioVqGAtULAAq8bjo+5QTQNVeCgomzVnLWndzwoC2
K3Jw7vXDJNWcGSt4DUVbRpsYGUSJm3xVRvR6StvgQ47c5s4NOwBLeIJtRNqt1YwcVnl4H2w2cyy2
2/RK8PAThnB0U8l5ngV5wJPi1+vMt3E7isWR3XfgSe8JmXSEfcJm1kcBAe5/u0LkvZDj1DWZH+TL
mmHGFH7YkBxwO3PTAuxv+0RPEZbT8p4baK/wmrIVoJ3tw8jqrMObY6/Bmq8W+f2x01+R0rCwog/9
mQYmB/nA9ZGvDNVJocbWngIc8HPWSkkI4UehYQcAqyWztBASJq8QPpMY8LlXSIj7xtOFw16DYFto
hoYOh1qbQ/DrdH4PbgfvukqnluqSMyinBW18MJA42gBFWKZoISxNkV+y27AisB6vF8KfnDIf3ECx
dkjETOGBGXBehbfC83kwASeiR10BY/JlIijtt/Bs6XP0CZsBy0w9OojIB766MlZPgSChfTWxk6nx
x5nPKOVNZxMRuboLu7tdNO1dPH2wun1ajfV4cqM0dDf72FBHlBtjW0qUaiWnLRL7sbACKnQjS1A5
Cj/64U6VH83LKAbXvKNwyZGPoDe3cyMcu2+tQRxjXkkZ7krE734DcVwR6rFFq213dyg12jp1g64U
CgFuoB2TtcU3n+wyQC5Bo2hqdeUuwiFweO+3aSzg9dh/fkg8ULysfUjDFi7LmFyiel+EWgMuSbeZ
26HGXlKQia00/yEt1+IrC5iYD3fahGoCqDVaQ0tIiATKmXh6nakiz+j1QYvrAoEoD8Tc9uFjJmQN
G6h22HwLbcli3pfsGSlCR99dZ0OmDtBw7Y0bLdJWGIVLiXhF8yjGIPr9IGLnIUJBZ6brRK3ClmcU
E2AXh/FMES6X3cCHcuuugh1WGJ7bUL9eRwuZzl3wppZTRepo5Www7a2ZWA6NPLRLXJykLIOWSRDZ
NBxwkZKA7shH4TLcSBnJHYzlMu4ualtVzMGUbP9F2jAMzGYv7CkzbRY3Hyt/9szrlRM1uo5NpsYp
1YeP4T1trBwtVf+PTvr7jWO3YPaJAVf/bG9UczV3eSVEPHdFhwr4UE6IHJKDurs75p1MFhdXHkTh
tq0xEzQa9MOP79yllVUc7S7XrXtbrtpDvv/A69rikRF2v/+EWHrdHU3tM8etAf3VqFaJLykTXTbY
c1CzH2vpfkhGMSJCZdeYRQ6ZA8B8OBMDK8JaCCHPnlTw9Q/EbxPAX+DlF6al/MGmczSKE/+qc8en
GV2I7mbGsU3F8ekQEbBJX7yDL8U44vVbRwkJjco7Qq9VybvPcS/ZtCqwccJrJvKQN6EkpvZiy+gt
InjyKeJXxz4VEyIk66B5VGChRGXZe3Rco3JJlKiSqTBdOfNnNNSEyur7u1SkDErskv/H+YaR1d5E
Fn+eJNaQbXRxWy9Ln2GZD6zAYQIH4/Vr085uKqhAi0DKLB3d057MlOgbTqFAWgetYanOBRrEHv/4
KecprCa+RCsNK6U9D9wmr3cR12XDCfHPH21o/CDE+cZzcrJQAf0nVRw1wsUdSDzQNRUgEcWGZ9xy
SyZVsIMtZ2UXbiNZjNymM5QNvjeWZ9yesCGPrIxPmTCYkfUaZseKPigUzf09Bww/ls/sHnIP/gqI
LoiCMCZlLkIY7W5avqjBB0tI9flb5iYYkchwi4NS+8DsWy6G75JH86vMrh/f880FKDvjflZVAz/2
fzj85Hq7lF36Pf4JAzXkEQbumrltQ+dxvXDQBywvYgofxvDS1pwWqJuK42GnrljIXhwBGMSpX6rl
nGBBEenmrjB0mjnqAsofaMNZbzAqoklef6bDrtYwawBLG/QymTWQBZlr+XwYk5b/ejfcjjCe8X3K
pjYpfp6hRAHdX7Bd9wXB/ghuwpWDsSQdtMn8q0JftO6ecCopaVu06kMgUFlG6gV4uruIK2pz6JmP
Aw3aXXvIrcFwi/K75TFhVH7XJapyRLhzI1H4lLVVWDURJ/5EKj2PJwkAhyvGubKUD3EijqTrhO25
4/2CMoOfXgmNuJbp5waXcQ/OiSkvva3f7D9/5g7oZ4Th0b2vy43Z4WB4JVxSp8tm74wK8iS8f7AF
t9X70ot92j8GZJxqSdxcRUZHMQyUej62ALvUy1YjxFF95MZP9uE4ry6pj5y5y3QrjMyFvyreX+F5
MzT0aKALSPWUSZ1vDN/TIAtC8VWcQyKpDabKxo00bKhJgK2UcyZTaaYBW2YlkYnwejJ95gjy2RpZ
WkZviVKDixGm2ydlc8tC15AB+aJrBDo+5k2UD/W/LrAqrYwXfX3Zd27qoDK6mv1O3JwPShTLR+U6
qM8TpuDLb00tde01qPElApNTjsR3elwgMI+3exc6JM6n9Dxlic56xySSPScowEzAWe05Vo9qsJRs
UTXLf7LfSQOiZD4IEn0W/ZVi3iCo9xcyKiWTUYHD4MJZw+Twi6G2KF2ySaTX9ZtuyZyrdGfb+qnx
s18FKyj8g+gU+JRlcT3QiFJV3DUwv55UKoOKTP4hf7W0189M9enVOgBn9TQb9kmLo7E8HYKq1fM2
VzNndK9oVSQ47FPOdMbzHvdwriM73YxTUKdS1ryOh8GhmQCxbitdgueL8UseANKba/UPYbzF7way
j1z7aDDaJb7JRQ0bm7mD6VGxItqmFkmtcOUBls+XmaZpm6SnVz1brCPFZjeNZELCbIlC1IEkM7Bx
oB8ijvStDGIEnHKsqJnnQM1cr7QQ6OhTjLXFmysuni79fGK2lzvzqIh815KKKJW3fnGO72wkXkHc
YIoD3VwqIVcgMmIEdiOUrGlhKNaoN/2Oqzs3bLguj9tm1Gkg+Uybowwd5nyeqiNpPpnCiHCgVOI2
uzz9DO8RYvnXbTg6NYb2inp40h23c3qk/LYSI0i/IMqYeYTkSnR87ZY6mxg0Q6nSvamKt6cBzKdG
/O1eIpj1fhiAOmsTmOK3ejl5jDnOYdx/LXyIWTKB+JbrmtCPUkV86/1quO13QwfDcK3vC/hHmp3j
4ZILHsF9MA72s+UXAPay4HTggAJTFPiXbb2pcteZBuDfCOGMUavLFPeJGwr3PlXZZptP1OHecelt
w/V27Yr2WThGFlZAsuBjxkoGrs+NdMqFpvwlF+lQwWWZLdCZebBNSJj8SCcMih9sYK7TA4u7sRMm
qqQxvfEb+f94k7bn7KUys3s/oufAnM8GwKTrX1sLxwnsNOeatCCUiR7x7xorB+LI/jczoVn92E2B
GrLVEbBeiy2QC6iEZrBv9CbxU1BQyYT9MEAF3gztD+6/E17d2cxt9RARFKpVf4hwTdDb4uqVifvE
mDtC4+0QBGerH3Ltj0w9+fpoFDJxxLDaqPVroLTGvcBwMIb6sv3ARTLRl7Bgh70rFkCRofdggFvj
VnQYCG2kOMsJjcUhrh3JNmtNB8SEL7LR6Tve/Ok+WPWrZ1aoEngyide5NtJVSf5s0yyAXZuNuyEp
jjsHN9ShMgoU9hwZnhtQauFkjq+XV+AGFSjpXcJQCH+6n34fM7agyS4ojxKw8bkNBIrtLADHyFlP
xJkGMdXp4ddw3oxZE8skj1ISR8wDUirckQ0Te4Z7lDuEvpXnmXNYrNvL6V/uN40qZ0XSCjQ0P/hT
tHVuNJxqRH8Uj2Qh7o+xCXinWSE4yGXylAGlZDnGnON71Kootp2CYdD0xa2QCwdsjHjgl1caLI69
baizoBb/xYZIBjoEl0Lp3XxadxT85hSITUYDYRZxUM5uH0n7r0oXOaBLzCxfYZXgGb9Pzldfay9Y
Y/88y6GA+miSJO5CmCsP0hb0JUwTNHP4wegtuVXei+uZ5eM+Mvmpp3rHAbTofGCn6tIPbOu9JtOH
5Vw7XLLvAe6JShj8k1FnGQHVdvSH2Vb43dAebNBk8uQRYVsphBZaa+AfFv7MYfpYil9kK2YiGvIy
S7aU1j4gSAzI4zHjFj09ONGP8y60VdAitXpdw9x0aJd7qc1O+SjDHPwu5A5wcuKjdNW3AnAxfQkc
HX9H74VomLa88e47OQCYi8dtA3hXa9Ca74dwPEIETN6G8fp1MBkwuJq9NiCnNERuupWRur5v0EkF
JcjgH4JNwCf/+1A0ZEw07IlVSVamkR+wtZaFhjSXBRHiuylCgXN3+4qlFN9CwiBMUvWujQBgtQ1+
GsTCglSJjOV6e0xuRUuVGkyTPLUG4aAa4DXTiS+r6Li/0zIESPMKIpYpYZCCofHdvOzBUyslI2x/
lw40409OooA+uapS357TBQrEsM5dHUIgNEkTIMBCkOFjBv0nH63GfEWwQJRfN3Ml8RW8vLGoaUOh
Lu2x9GAprlglSmQ1A8KSDpl6nmMAoGyPx6OvtNDXshFRFPaed6DJAIeLJASDUskYS9RMbnuCwID8
QMmpC6b7XovAgKo3WxAR6pzw15VgSegJ5Ys4KpfYgPxglGzfGAlqUW0db7r4wopUOE/SnBj3Huw2
jlUM3yneiyaiQeZREDm79+qhw+59ZOcxqi5oPfdGKzcdjc8iFR4E5frE8sSEWsCSUhltbTfMNsfw
/RkSSfYrZfesPWSWGkX43RZaXaVA2aTzRY0c2oFExyLxeZx/BwWVoWiY0a9nhzqcjg28LvL9QaPH
INsL1kVRW6jcssVdCsedGeQBg6ycVAGAfVc/LjqUc9kUPA/pRILw8cWYdAXP0AYlGEs972dr7AAj
ZV6mwmqsRho8M9DofdHnPk7NEZYjBrO4xPkEV7Y50QmWryHQ/kFnmX+pUWZdsFVWjE3JU7ndwq1F
LyZUvzzAML1ruMBSpUmHwTQduMXOOdAXFIlr5uIL94vUmHMHDIVdA6QlDdbusg6+hMNGTE6XRO4L
aVkUcHMLfNxLuUpYNQrsZ6yhOsY7ntjCzYUBn51E6+IIcnC5PRUxzxuy+TuxPpqTpli83RafScym
qJQXnj9WWNBtjvrabVaUUHA2YFsmlAWZta+DCvb3yc0XZOOjurNRD6i23Bt2ckFQCY3QMr5AI746
JH8HXXwhtS+nG7G3ZXTRQciY2Gk7KfuRTQi4NQafMqqNeYQWksMxkwDoZA1yUOru2qHn4B8EUrU5
jJEaCbl25tlsHz2ZyYgyz1NlzdI3o+wuvqBFZtNcuVYYNMvCYtlj7pruZO1/KKE3dQqxuf0PdiPa
HZE8TWDWZ0/sE/lmY7PTkY4SVXQTnyRWJ0qR7izchRRiLVKtCk5trKfnw860F1ikfFUPYhtIyJxT
gIk5gmub7QvQeC2KWiqoNk0ocmGeVqUTTYNo8RXRJ9utnESMewX0UWnnObc6uqlYIuT4NNgkV1Ce
g1uCYxZrPmKrkMv4TsrzTqQQmEwaK5at5N5yAjTnr6bIk4Qzi6F+DSHarxxuaciFl5Wig8R4VLDm
Iba67NnNBFfNhxjPPfQjxqHKUDIo19KgzMPkVX82Q3ccKbZ/OtV2NMoN4HQle6aoQGyN6KYYBsC0
zsPk2e3vefdR7vT8Ff16cPMXbq+COMBDWo2WFyZj3f5zliDeOKIQEP4CroHTGo5mhNl56wLeB1c2
ZY5AvugPvQbbfDMnDBYjJCI9Qm7fUJbrbIzb9kxN74hBxLUJj77vz7Org9e7jKsWHeqpuj02k//F
YQ+z+9tn/S/jtGkJ2gpc2a5nZkkdIJmvA4Sa9Hes4CT5MbCt6PZ3Hd3MrdlRr7zAikQfJ4KEcd3G
gaEJWd3MWP3VxkE+RFdaImzxsklgbtGpVnM1e6kthTaIeFw68a7JxN5ilRnSjz7cvFuN823LQRMW
+zjKXc0FnMwutyUv8mhnqDHNwvCyNeVaXoSV1zjYRyqVI6pCtoRACAdLzrlaFqZ950lrRE2DqVFY
QwyoEYVtH37z5OuJrvqCXTbazXHAnndM+9eO1aH0Nl2HufOsAgRqVLROwOBxXP55pBcOudTaKPm0
viRyB76WcKBMf3lCjHBK20g17alkxbCKPd4hy5t6TbKaksQsxTGkgwsCnOWsUhsXvHDOzuXiHGxf
4HURysM2ByAqyz1g8zbc8FfTsE/XsyW6dYB6rxDwgXJVm1LfJSRGwtnNGH2j8zAmmXOORRT6D/fD
oj653Bw/6UjOCSiRxnBcoZ5VCFOHiiZ5OYkI1aXu5sUgrE2yZbCbjsmMKtGLTSwKhR+/bnXyT4G8
ZzroTV+slyrDlq29v8EojdImGuCkgJ7Czu/DU4QwKo+pI2T6b5ejARYmtdebOTTkfyc+7u7Yt6Ub
Vs5aY9dBtncjlnqEdtBAXtU8dswDeqb5bIVlkCEbkS7ungE6xsr0C+inRRH5KomprgqTXzUk5RGC
EF+4758yKqyQ1emQsxhINHDdpYLni0MoNfGKobdY7dhABAN51EPc6M0GdGdp3nKHdnSkQRb6KX/L
Xw6gSAczQwkg3jtvVxryLMzFYYZ3i2H4wotyG7EvIbV5lWQiI0mNRXFFy6abqZjQvI2QNf4/tDBg
Bt+XVjmA9ZEgcuWtsXitlIVeLM4Ov4rs0w5rz/o8T/Myw71+4fMxusRK424C0PQImMX6HXq3SgOW
75E9ce19T4mGNk4W9876efmf+pTuo7gwFEN9F8kjl5XHVUQY18MmApnqa323LmG9QxlSPlF2KXak
QnHtsnDHF0VL13ZiJh/cMmxqAs9qQmIL5KA7fR2VDLC6k60kjG5dDhax4avg6rYcz4bGJs9xXleD
7aDjXkGv8nuC1OEe/KffpY0GGtyuyJ+Dx6PbDOjE93nUq/eIVq6rNupclxe5nFQgYW2jhyJtkDm+
5bvkPoDskOcYVPXA4iB2rlqoblSQNAtZw2/qeOfdlmseKYexKlOrrP+zsTjfh+P8Fak4L/oYcmkB
2fbTw8WtVYtTflJb1xXs0M5CuZYVNX15tt0zDw2ICA1FF8z82Jy7IjjMJGwnCGemGJHlC0cR/DdG
8ye3qHp5MEnVuveI6ziFlSG/OrGFmOrVbE60sEA0goFdcTrIfn9wnj1ZFXgQtW2Xf73vbMApw3MD
LCyxCWlqMB5sHWpYuHaoTNcqwsvnfasXgHx8Fsa4qEfpCeHnAhgn+ZJjESYOVZvPLdKqC3Pr/5SM
LbDEYMu6hbmkEGlu+2mhZHe4BzK0bVNNjcb/h14ccjrK7QQXKnPA8xeUPh8EUEaKnFUZvN6Gwoup
+yNG3KjVCzG10+Yttz/DZzSto3R35uWch/LXE5wpyw2kgIjjFIhLaHoQewE2XQIRPDQfD7TU791J
j0PGSB8Ws268i2fOSjXXaMNNtV0rrohc5RayqYoI/03sgTS+xSSyd7lwRb+bJT2AcNjiYgt7qKvu
eRlihlsTzzVr4QcwXBzFitbe8W2TEhHkxE+3KyPQwcYCb9OybRCTN1qhdYxHhrsmbqo+H7UzyjLj
jnwEcVWfnYosrGNEibdbjClTpWRSOChFg3y5YR6ld9Z9Ziw/rPe7+1uYYNls7Ub7c5Ka3ZeEOCpw
YDO7ct9t+aMxwpsjy5I43p0s8CGbdp9pl7U7MjvSIJ+YdhfIm5ZkY8hOZrnPtSHnHROScBWXSEGp
NytNH3b0S3GMaYr8UAiorYZfpxLhY958MIRqWo5XLWEry375B55zyHHetm4rYj/7DqogcSWzlKBa
SqmOnd4LyGm7410AGUlyCi4cBr0E4CB9IauLv+fZ2vDvFbe2yO0DYG6dHGVHg3YtitVorGAD2mje
jPMGm+3gU1uBfkVlwT171BEK27k90EyQMETwQ/B//xvyOK1QWyMw0maN9XHjihSpFi8Hr+k/U0Vz
hwNpm3FjLUQQX5eP87jfH430WbTwziXyuCgfR5jZQ4JVWr8oqAsMhzMb7/BECXkewOQugZV7wjoq
xvRITl4U6PFMWzDF6ThpRZMfLAArIQSRTJZTBst+IiFlM50jl9FOiEb88nXkZaJ0cBM0EpoBJdV2
51xggEdP6XsZvb7YuptsUz3Lc226VgYmw5W7K5aZOaPjea+RaD0F0ZPxUo2xniRNGRHj9wtnLRRJ
go2F2j6tcTxDgbeZqvWGiPcWK18DJ2ZnrXXGRJn2g7rxflCFibpPrrm/MP+ktSiHCJoMMlj8WcWz
vxvb8d2GFvNs/vnJVb6HAhp118xvYX9sqPTiR+kOrnET9jdc8OJA4G+P9t4zdJN+iMvK11hefYIo
VG2nHdhYQyE/QAIVVszEm+3708B4Ic2A22XY2//SyIh/Snb61S4gvZktEro1IbVO/eihhtqqX1na
K7injizEc1iCGy51+cLnY5oWSSyfiFkbZ8G/rWYJtNioGZLGVBoothKgb18WR7gZ2b2RAhLGmuMG
5Au5vPqtufwFlBNRj/U2hgzdVa3zhFRmlpwwjI0XYshGDJBUWAhxVcoIb6RYfpzWDmJvbTNEubI2
ECd1z8VWFQpDFxblveZkLJQJOgxm9FnhG9X0bbzqa0B6qAEsY6Wl6RA1fd/ArJpwW2/I5ElJVZWh
IcmxzmRgLTeVfUltC4Ps0nj5bZjfsp7WPmy1E3v9VAATaF8gilgv3gzLEfrTYimkKM3tGiVJ8Spg
jof/J4R4NcYXA+srBgN5uEWDIAcebglEpi8m6cx6aCwpVSIspDXyWmdC3gK0pGY4Ff6TVT6KK2Im
LQ7kfU0Jj09ggB1EKPtJdkN3PlJzKfyLsdFUzcnE0APqCuCETwEQwQdZLQdNQfArPcwB68izH/sR
5ta/8tXTM52bjdMdi88cYH8KLRFltKbj1DUbiqY8cDWY39niVo+6Ay1d4v5+XpEzLrCKIqXTOIOp
wTSA970eWlyqFjzsp/W4cTqvinqMrp9/80IJAV7qVTcZBN5l1GAzvJtBCP7g+WGWzkOUd87AsJ17
HCsfPLANiqMiIkznm1ocTvtFOlVtp4O2yfGdYQK3H23DfNKkN/Xfqxz6pkCTkl/EIxYQBn8ScRvq
MSVOg1UgRqgVBLX4EUhEaMWJPopNfp0UkyWQG0twgMfW2WgDW7/oLdDaFXDuXjOiAXWUpnRlnN7P
bmPrDI4Mh/hyc8STs2cvwMDXHPpEBbBQl+FuQ3Z6l7BvGQ4lgu5lQZbZxiNiKnBOQvX2EdNQshIG
XWNl7YvFYyIbCEiS5/Ahx4b6VH+wYmj3t2RvpEHHRqGJqJSZ7RA+6kVZlyvqobRs8tYGdcSe6D+5
V75Qo0HAAfI1BaWsuiEfh4abkkdq76vPD+jqrIsDVXJSsQGhROVrBVJCi1CAljCV93XUD4o5IXQB
2aaXiuEcE89bOl4pXXyG/+xdE62g8AVzV6Gt9uxVePJN108IcuitMGUDV6A1/Mx+FxyznizOLTcu
JbLm3qfwZcFrA+37FjdUfGTkQNqCfalVP5jqJTCooAxtNM1x+GPffXSi3E7U/G+bl4g/ROQc/IQT
ImuoQLplrTyO6LphvkZkvt3gNOb94bOchQR/tK3OiqvY9wiWtWUzSC+ofLGTuq6wCIHH5r4cVHuR
B8jgqP8vCfjPF61WGjBagdMOY/B7w+kXQ6hBKycY3u6L9XVYcaUzFlUsw3kStxX26uKfzZ2NFZ1M
hAocnp6fcytGFsEGP5WeSrl0F5DYCi0CgmX3wrjR97FRd/muNZ3f+WgDbhlsMXNzSBVztiIFQyOT
WGssIaQ7UKUN6rAbLKItUo+JlE5UqGDxzxjXZwxcG056jZ5HyZrJjDKOVzYWXSshQ4cBRCVtxs5z
/Ahz20sO0ATLutA3Qgt94l+hkgPoVva2J+1D2soi0qwKBXH8zfpwT6AZh6d1LPp1EWlKLIf/ZZhG
I9q5Jd5BDvCJ+/UW1ddToPjO28iS7zQdeHneP39SjXPojNUNBuvQ+WdiXgnN6tpyxn7vaKwie2MM
+6wODzZGGqEGHGCGDDHiKV8EqsKgZJQARGRAAlWdUhwNbkEzzfImj1+4IAOXpt/lQ4XWZQQeB4RQ
Ls5CKdXpokCW3X7VxL5sDrmg/4K0hQ2DW7w/GYmcsezQr9Zfv6hu688v5gpjaOEs75a2fye88745
7/A6K1ZUViZ7ALOnoqHuY6QFSqWesmiV/7d2rESm31ebQDf+i+t67l1kVGPia5XupoxApqOxuxDz
xmCtTXXAfulQqhJSgKCejzqC7w8cMsiOj+tSkJKNa7uO5GZTL27dpdY5cpjgnMuCPntZ+qWR1thX
ypD/hDhHZA5e8UZI5DsQjY8Qv4stzk48YzM5unT8FXvq8R1qtGzvKv/DK8cMOVMkFSy1srYm2Z7I
xSntplyc8eCnxI/8PI8K+fCX3q2jqSQl3TlVRHt0w+IRGhhaLBVxiK+41TR91Y246O3JMhq44D0T
uTmAPqcdpxvt67v1n9opeJ3f0TzPb4JPER2CxS8O5god6K/D97JjyeDX9+UsJq7rYXo1zDzW6tcA
KCICGiCJnyHACUaSDXL77rznau9y0NZOQjMLMMySnagMc9Fgw671q/Be4SyqOA8MD5aDl9oGy6o0
/y76EGmkwKMd+mIRSvMl/86oEfwmyXvZB3aMIIZ2lxUigiOrD7BlQc+cdVdUifasXikGGDbULdKv
5KjSRvD/7NanOIGDvc4n1+zMxz1TO7/L2e1Rgk0rwBODw2sqX3BNwU/F3S2C+SAvFY6Lo4iKYK5i
lHhFlPrFQJ4WAGuES9r2RkgDz0eFlv9Pg/QY2Tue52pkWn1AdTdLefC/dwXYPF8PvPQOHDJHa5IZ
cxtjzSIgBtuHGepJ6rK5oNsFYLvIn3FL7Dcg0RLDrFbvLMbOx2kdiFRMeBsVsKuaHLRu6SvgmATX
XK9ENGNreURLBgfMDqmnnZ89yjLlSriKmYmNh3HbNS5eOoYPmWaMoscr9s21I4RV2bqg2eaKXkQB
8u4xXtVjAkeDYDxsNL0nn3v85+0H+xT58u3ot8tkh+AAseAynn8wQV1/h3SD9N/A+MWF25OxP4J4
/PJRK6r0D6RiFdxU7Eh/m74BJYoLu56nyuOndtxUxoEApRxuBlXfZeHyH0ouacnDvBcoomrQBJvj
d+StBMLoArittVOAfJOkFxN+0mRPaZknrGhN6XayaF1sjqkldhEhlA2tguqFZteoSR4UEn1PUzCQ
CzzeYMH2U/J4XuWNJC+/Wl5McU0Qr7uJSc48bcPHQnA9ze5RQ0PdpJBEPUJLxKfCBvb0ePAZjGj1
FHoa+dSl7uKbW8Pe7FoTO91R88JHEMLCjlmm4iO+nBv0duhAQHgnGgVKXwWdUwntGZLAIjyMiT7I
mkY4rXSbTCoFpZRmohE/kyvDpLaqhLcGOKCYo0I4wEZRXb/ldLhFhF3x0DW3ryUA8hfzLSOvNXvX
/0SzDkXY6AVv0V6AcPNUXyxHdiRHkckj8cSIb1p862PzYG1smjC2lO0xmQgFR/2PgMvPw8KY5STg
whKnbOWaMfFVDP+VVJ32enqKZY1wCEAo7BkSdpRSl02FN6paRf5A9zwSbI2jCFRKhiuxBjQagxgW
We9YlWWgDHCBexgHNpfusxnT2bUwz8BzpprUcyZBLljh4u+DNnxPxjpAc19CoDE9nrtaFy+cqIfS
PBsP2NnUF73Q1AZeALPUkueuXDA3qdKOFHlLDO2EQxKDAzfnV/hp87zOK7PHxa8xv+IJ/UrNNUmm
pKznGPOcO2mZ7hxpBlXI+V9JWJHrFkBBZ8+bM0VhR8cIIXwV943Q9lNl8/3p2csBOLCNgJO0v2VB
jts0Ove9PsPQ4R1zusaqgJzuuY4qmDKKbcyLXZ1UtoALJW+2fSvoCVYz71A5pY/C6RtL6LcflgOv
kiI8DrMJ2DyRc/TbTPvRPZF4kNxqw29YMXUxvi5Vr8nfMX6gq1Y35nj2MFGZ1b5M7NdHo0V6FjgZ
qGSknFBeDl8fInHtcgoj/iYNJbsmxPaWt/vx3srHedc1ia8OvpMZMhRuC2krIqdHmR/uLikd0Gm6
ThNMzmMPNtn53DNb7Y729sJOtFva+zDb0FdRwcyXNodTZkJumu/2ZHl+vmPs+Yx5jm4abdMhEBqZ
T6xMvVIYTp8k67DzKYizOEzLnWhQI39RM5AcbEtoyoJ3DI7joPnqKOibjxl/uQ1W6sezhOeTYNwV
g26PEVOCpEq0b6S8Aj1V/xWS1vzdfb9EhAO0MY9shKmM+26yQu8ibRT4yh3LPOGiOzn2hZRRb7Y+
ftBEZU3x6wqp0w7Zo2bb9a1naYZeaAVeyrcP6aOaYmhoPR/hygPKVVmOdr7AlVdjRzyM/tVxQzK7
Wuyw6KyMFhQvKDs3q2KUx9cCmehkLrFJYj+VBZl3+bN3yGO2jlysgY+cuLb4elJwAGK0qWUZ+w23
FuOm+EQOXyZ9Y18g8IdGffkG2xroDpyZ7APDGNXYn5DVwtx04MmlBDBTbYlbk8dfaPj7Fnl/E2fO
TWEusgmAZ9d/mzm5Tr3VNZJBIX4+GM96PMeQ2wLmowrqTVuE2tJDeHU1zSjNzjoDMWdokey9HFBE
MDWEMD0RvGmHX9h1aZWQ++GErdsuWrz0jBylq2nMTdZ5118gvvcYWOsnvFrgvk+gss/4QZY05h1N
jGumK9ws+pxj60UkClDyxoYm0DRla3YB9zJDt+kiSx/HGsExxU8qIind5Y+sdsLRKjGr01BHIyj5
7Cdgs/MzKyCnsHd0GmJQY+/4nq92NJ9M203nvVzNrwwS5hcgTeb/N0fY0LdLBgs2RNQ2xXNoDKVF
YP3CMIRcF456yBXQ9fjOO5Vk/NbElV5pwVYeGJ4yaVmCoyhwrx9qv/s2Qqd0Uzy+UFuzhTP1KYMh
qImU66EqdTegY+76vHF6XuafP9ue3oZA5JUUnYXvDQaL89/IKN9SLIiI9ufFrtBsmdykeevvvYqA
rX/Kl+9RPEx4mtK4W2OESzgM9e+PVjTfTRz+PzgKRL3vR1XvP84OVbvGhOmOU5rgVV06vfZRLmUQ
801Occ5q3Lq6tDDzXWej7Nu0AkuTlQL6GUzkeLRBYgV/1SRWVXAISH6NGozpsdEfz+NqMD3voKGm
B+OTnx7v4/FAm9ihRlfyQHuJzZRG3retxgHe4TzH2n3b7FkRSuLzOwvbfjSqEZFbajliKZG/vHLU
/KybbTJjlnB3B/73B45mS0U2JpeLYCVacjr7anNoy+HCHEMkscoYTpxE+0Sw0BnWtuf6PHIVr+LD
3SdvP9DkbBDDNxkfN4+B0kcIF0Cp4BJ4zMZRrXHtSefriONhL8N0M0/AbQ+cHLc9IPHUx9sOn2UT
Dpq/i72xPNHzI4nowRem1/KFxFIesGXtObSXUeMQhmIuRUMmf5QbL4wQYUqMclIX447FL2E4rbcT
hZOl/PFu3oi21/gOSsgjjU5eMOEwtw9PeSBBnUxSXYIyNwljgCymzTiBRZ1dCnVf1cZRGaFQ1GY+
ZOOTCPozd3pY6w952XW8qciaiOorRf4OfFGSSvkH83rCfYgHBOFk8cbll+BdzhCTt4fr80cjkyLz
2Lzt58m17SPlLpN4uTW1RUPfnoRWaoR+FD/JNcWUKVyAOQYCLKGyiiGsKW8ysob8ZGVPwdWmYQ8X
TvRJ4C+EdQE8QfqXVbjTDbgnswctF9Fg+QYBd1/y7DwhwpMyjEdtAxHjNAQenPYBWvN6bi6jb9ot
Z8MnXy+WBlpEJNrdFf0iZENMQ7uba/cNf3mgB81WmdJ5BY2NktqrQTnisSRt8b1F3u9cQDzjfyrQ
amVxw2qCobYNchepLUfBk91/WedvxNfZxJ0Pi8R3AgLCplAmwyre1GF7n8p4mA9L9NH8eMu/QL4z
JiVy2wpqnCCGSbb5MdlZQieoEIV6fGHOaVZ8liAVi8HuVA4HoHac91JtFRg2Cm3eV1fcPTyDKdAt
i9fLpJOAj8VcEY7T9BMf9rtK7WJruRDJ8udtMVOXroZ8qtkhjxzT5w4se7DSXCNwGGM/vyVzrr+a
dLHpuZXfVlePvP3fZlTJGE7Ob/yv/KJiD9gzrQairXyhu7wnCoVM47vO767eZbIRaTHIuI6BiU9P
GLCmoKIdC4Ywk/6lfif2PKTbUJO0BXQ6zw6HQJu8VGKjw4hL+1ycL0LmGcUt/wUiFM75rdRz+QfR
UBLt8pV9ivGpn/qRGU0W28lxFmcybwjmH7PQ9LgW6HS3EOBS0UF2aNbijDley4eUdjWc9Zc62jU1
30j7wh5yRmowLdR8GNAWN9ZJ78ArYcGNjkfFgEAifZs6CxcEIbhnsSbTY+SyP3VG9dD1UEaLJkw8
Yf+72TAgktSVqP4zJIpeoo/CJxnnvTrp+DaZupJrmZm3EcB/5rrdVdnacvHWxKXCcxewVM2Hnfqa
dLGeHXyJdqHsuG8uHPHEQ5N5HBwEi0UqDHT32fRJR4aop9YaSZY25oJ0IAjjQb3RGEGyo4GlXVFJ
I9gb8xRjdwvePZubvEeXJdJ1QkJsXGTNXXunf8oswYHeonj0HRTppA8JOoqUxEbetjh761EZBRxC
JhpbwlAupJktvtgn7TdQq9RKRsxlYNpmKslWKxrj223B+Is19BPnx6M1Pw+Ln/zziOrojOxbXnWj
/ThD/cgBXn1zHuz5fC4ALl62xl3H+FTRL6e6b7PPT8hXSnUzSv5SNm4c6wezTsyzqz6OmRvC+JT1
YymlGdefyF/HWdAmkeLW7OXUomr8UPyHuifcj4FCSEdXyYcqa3TDXfHQdo6bOGb4MPhuJ5B4CbCS
LU1BRaEsKCuxEMnxj7gSGLX5fbGtvRLEaI4HYK0JCBANulBkmxtqKQ4t/v4CZbF+ZnYytLMtBbtd
sduAMXO2EB+bBXLi8KoCRdJDmeMcEGzkf3Garcq8OSR1pSBwoL59QghVlA0OWF64+Sn+/tmC7ifd
MsPjqoV0tmqD0ucYfxvM2sjkDg+ViyzOyqXZV8aW13xwccof41PF1UHbimF/78NCByDGH8KcZumv
lr992DYAvrJLIckfACzun9LPutG1TVJ/RbysLFVaw2DQs4ab17hF2C400e1EHErFoHZHEK2NfF+c
nmIzRD6PjNilGeoU94x79UMZa7R56dHFCH5xnJAGGxxXJ9+GSzPj39CSg3EFru1K9YZ7h2bKQgzx
iQm4RNUKPixPdA8FDmjMgMbbbAmPKJGVAAlw3Adwt7GXXkITGVfgv/ihJFX6ZDyvMbGfuTXPrf6b
qZSRqEKtW1MlJErSL+jR/L1dzOuiSAE21GB7OVqQ8cV3Ix27DSN1mtphPOdcETBDrML4s/s/ndfs
XFU/AOt3VSZ3gzzIcYVNmCSSuIMz38qBeo56MLoMnpa0GNbk8Ha86rcQnhsPhRcqSuNeT85dGrnP
42PmkNowokIrkGY2DoIMIhWaj9iAXv3ijssvw4nmM14455CDUbgE2LuopuS3petFKAgbhp5RHLCQ
zC6ilQ/6uY9FL31rLHQcyy9FRHi5magSHvfPH4x+X52NxQHQOBSKWYzOfBuc6zKJM+xqlmAw92HO
RRZ53BaEdguCIlwiOqBMgUnl6iQjAIcCsvl/lQttQNhza4OgsqbyistMyCC0ERWpHKR9rAv9FgXv
Wh/ue9AFzuNEzpAuxdEJyxq8Tbt4wu4r8K3yTCj96qxc4rzEfNEkjQsDZsIkLX+Ft7lYj9cMF/wn
/z+puWGTcMa694boI/l0VLjGsAHK6OHE5UCiU1ssUbelnkb/T2fjxsla8VlBVQK4MIKBTPmDnrKh
hu9bQsxH/OF31NDxqNKAH8tiMlAqK/wifDsFAkpa/RpcZr2Gz24aR0RB+91G5pyADEqXqTMhgErp
pjT60sfsT2KE67CXS/UhL2yyKfZ2XIodYFJcNhD6doI4SurrUqXu7/1p2oB0F4p9309xk6+ooM7Y
83pQ08IIXBXKwW4qykxPgBZPpFcKVEagbbKHEtiV2H92GVa7jFB+iy+BQ38FUb/y7FG9pkyyVcUi
/bGPDxDrE9YK/n7sZ4Tg9UxIyxzT8gMDDhgpetzslffzHMO4TSLW60QjtY6TcSP6iB9ye9/0lPdz
/xu8u1sR1kmcEbhVFagJRtdHMNXRyYtbV38JgOIUAtx40KiMEAiB9/hKVgg9Lv4tUuKhVcKccQUo
rCwSeGMLGbevdCjwX6drgRaCUnGvy3lxPQaijZElXNe2iqhLNUioPXxyU4H1//CLuDFalgGcAvOh
TJdn3H9CJgntHi3I8GQ58s8z+K+L+oGvE0o1JF5DStJHF5wc7+KUj2IIBi4qaZd7UvCYRr8TmLZc
8F+/8lcjRovKwJTsWBZiRfG+6DwYIQYqEkoZqiW2bE6DVFi+2FomRzo+vc9LG89hK5yGJ2RkZUop
WpLWHE8+oi5NeBFXKjgwFJh+OhAlK6Jt/IQMorMcxLI3KCfhGryEi21t2Tp8tdlBPX51GLndNrrs
+oOQhunzsjCp+sroZDXzeKCOkHLF38hkZS0YLm7VdzcWX5yyQz1WHOrTaH93+7Lzqo0QMR1522rQ
I5uZ6eXYAEJs6XWSceILh6wacp0PIznTe7a5OnOozP+8LFWNKx4Domqg2KgzmHMrPpxbmJivONxM
EvpLoLS8ob7ej/hZDRqAFAtCxftcfwWBWdMq8CCaiM/P4jaj+mPM9mzJFs0DQ6yBuFGXNVFBUDi3
PO57JC/l3lDOmX682eAUoQJLq1Yw7y19EXBl6lZfZSYnBipoGpSHE5ZGxk5d87j/Iq1P4fnl/Afp
BbgFOgPugDiLqSPrDIb4mKNVWFzUzo2NBt/rhyp2fu/4SqekkqqO0im9XBuZ6cx1srgHb2tc1a/9
ZIlYtMPVAMnBvOKlCojv0O5rA+InDpNVLBFrq/u2twe6xYC9IzgvKZZOsmC79S1sYGl0NFn3SAPQ
u1AacI7OFqHgAhpXwVQKqlHsr17jAo7M4eWyiUETqUTjb6nZzSyyGDbh9ncPmLpP+wsNxdiiqXHb
bT2oE72NUHU2cliiRVmU+RUo3R2Wt0gN43uaCcxLYahhqi1jMWLZN6ptzZZbJnuJIsLGMvHEN9Dr
MFvsfs3+wtTq0Kt5vQ7faWNDJSR2+4q0gfOjfLAKyd27blvDJsRtvFGHqAbifw9Q3YbyAHr6V92S
xxwUQ1zcAPy16nFNcZKSkLd7wTaZNkt8IrEOhWeo2xCzpxfNMTfcuzcySq9EfWSyhC5hrQQ+D7Fu
46LJNOSzocsxTJukn/BUuCaZzYKm422WPMfAiE02SCrH1UwiwMVFUQxMLlwb0xGBF31mokyPpgJ/
WTwpLmRydfUJ5roAh/foOs5Y9ZNPfuyrziDwor9XlZASkLOYYe+CpHtl5sF5aDdUL7B2ABK6qtMD
B5jwxU7I50a5Rq1LGyEcO8DAE+ocADPyl1HIt71AdeD7NaB9Lj2liqsIasjJ7kTdRQ2Ez1PMeKP2
rDLRFiSZTx5EpWs5ovlZk8ix6HmatH7+2Qq5DisDE3AT+G8HyZoU3BwxIRzFUikBa0N9U3MwFtaN
qu5u7vqkOLitlZ9e6altM9ICB34s0FAaCTag8hsE2EE7FTqbioJr73z1KMo63QQBbDI1s3Q4lcz4
G1PnX9ClPJeIUPVK/FMPSK5Pyo3gmqLIjoEzC0xY2lbN4AEfc51OkRfVXhk+WTYMp69G/zytmOtL
hAfCWRouoMOouqEaPHAvh1cqQii65vwkPfn7ofRrF0sLxUumQnWi4atboCJseHxFUUt1YeD21KJ7
9W+cZJuqsoYuq3NpROtzED+1iDlXxb9ySjMFLx+9BkiG8e03kXDFEpGnmHswFRD6BKY2p9BVEuXs
dDACFTHWPlaQ6GR0W9HX50sZ8pjdsC71JdU5FrnkDNBpSTCbHqN7PHuX3cJg6icKHeJScHaZ/vUT
92YwBB7x7lD5eTcoAyMoj8U+TRMuVNTWEqy9InL2tHQQle9MHOir9yWQWFxLHeZ4TGEFck3Ds4rW
MGSYm71w7eSW76Hwj/RB6EJXGaS+knMRtF8sys8dr7PaBzpU1569yzGdbTx/cGL0wkVnVP7nKHHc
E2xafp+dhF5++UCoYSxAqXYS/llt2h5bIJfsGZaBDbHCYEktNsx0D/YeP1kGA5zpVz2GejSgg7CR
Z17W549PV5tfYjK0glWSOBVZigru7JE5V67Hw/mZGxKyFMdDmypmm5ODHwJar52RTQtUL0o141pI
KBNjp4djCZ9Tz5vWMguWD8rsOPqv5A90rKpHS24W+EFYknj30yD0KiKC3ww04txe0lMF4pBK/tWi
82XZobCZy5rNMBTRArxVKHPJzqQe75z1oq0AtcCz7boEvGgi89e50KOONq01WJRjvktoH4Nkyx+T
Tw16GgEc2pWMnmeS3rZXL3Pvom0ySvLWp/NFboiEb7Zkkl8v6VHxWI1tOZGpapRkhuPlbAeKuhOu
qHla1lgnffCOmy7JeZOY3py0e6W47p5lku/Q4ZbYU2XmABZ1NxprmZ4QK6cwqolP2JdiubqzEPn5
vlnyXvvTa1LriNY+CfYM9DrAx+Lm3LUW9t09BZ8+nXPcVRmqPMtoA8a5dtUnYdz/e98adYUz8mj1
rmeT3t/1xmHX9zskMrgGMWDIGVq7pOMR3Me74IPAJBxnioOsydvLaOcLljCKum3QjXlvVDZSDhrI
bCIFVz8eZqephrtDHyktFeY+zdmC1iv6zPFs1V+NLup5w+0nZckuyPZAU45+H9DnOb+yGl2x9J04
Tlo2H69nInOxlZVKTRtJlRr6i3nMZXtD5ZcQDXVZjO7PhZPY29jqH9PJqJaEWlgVQR1lVQEMQ6Bt
hPHBuVWGM1ca/KaCTkbrMP4Vu/Gkgzr1Qm+5gVYGl31AoPa2ePh1c34DWkNtACJ8PbZSZqwxqgpv
5wMT1MUxxa+onn0AHJhQNIoeUjEcXv7gNzPZwzT8+Nu+zZoC/DBTu38+VuybuSzefc+dKdYUUCTD
0vbM6p9J9+5jE5u6YMSgzH2IHfJ6HEhwjCxO5y/gMaMuIxD0FEpYhDZJj546OCxyXEo67/DJajJM
F/CM70wCje7A7f7rMY/UniTawlspoYWUO2TloYWBsSHtlKwbPXDsj5P9rl+3zx+hkVcgWZBH9A8r
n1sVSldj/c1/LrrdQEavhia6PSp1tcnYq4fT7FoMKsP+Ho9r2hF1bFY+v7g8VFSmD9UnKmOchczL
+0cqFkaAyx4LaCpRJHyQhHi3DnEksR48rTTHyVskUWfo8dhiowsjoGdKR/mbuomXakPQjg8F60ip
Uzl8DC/uDrMSutJzw4cpj8LKdGw4b3DPJgsjDu4pJ4bYmK0mOwWhJAc9OnS+DX2mPpctATgkkUpQ
AZSgSlvXio+GhEBN1BLuVhE+7uZfy9TvmMmGmGV88AKcOS7pj2ry+xGZu3+BZd4C82CJx3R4FzGI
8cOaRYQZuU+vNMoJ70SVIE/RXJa7rs0ga+rUqap5DH94KQaUYHDeqsqb9nhqyFXC85vCjdKvj3bT
CHAUZ1fH6ThQw6pPZISjvon9K/gcchA4Gl2yZXmHmeOcsYPlYl8At/3bgpu1vJjdgfcj1SnAKMkr
rSNh6aZwWa0P8SAyKqSt8ZerTJ0poiM/zwOgMFFDcm3wOasORgQFPMAbk6S7LX4yq9eI4TiQl9qW
zz7lbCssONVJC9e/XdlvoLGgWWChXFTWQASdc0Kvn6esfIRhCaRZp9yhk4yMa566HN4rzxecZtJl
edRwTRFbIfA6RRPDtBXW5N90+8f5smJTiIUKYM52ieK6Kgr7yD/Fdlgh2JufoyMiKZK3vODL1oYN
1lFhrMxKXjJH85x/jG00mQExE8vMCXMdpcpJIeFCe6XIYrM5Rb3SJbtXlcFIdMwHSGVso7jjrcD7
T2Z8cIz+KRrpBYQlkUPDfFbfaOSiNOcfbhhjVexJQ5yibyCdHIc49k0BD22prQW7HwgQMX3WPcg1
f773dnU0vGKjcr0heYqfs4cKz8Id9wFZeelC5Dr+T5rmY4vBR5eQ8L+2Mk89YScZa6mU0aDHTemf
6w/vCzSDUoMJciXooajsfg33VAa+PGqbMJJfvwRhfqwaumvFfLdKrTzJoWGSMBAYolTjcnsucwwU
vtdglA1GTE+Q9GnGcLGMjCWKylhk1ZkvWVP/P0nBVXpM+551B1avCRhbHP3VYYh+3x271DddISs5
KnbXMfgAiwXOqMcFe+j1c0Ya+QB/wW/G/u897oiOMerzuCEr9KhQ5YBnGIXIILtPOZaQGK2uDPAO
iaRR03Vr7xSP3l24r/ujFmCLUgVaZHnWatwFvkXaqTFvdcE7z0tg5jUafa6xes+ZgIRaTjJ7X9cQ
aQVi3yKzS2CgFLMDGR8dPdsM8bBCU1AHuuvX6dl/SXvBJH+a9TpQUut01PY5b0TGcEcS6Du806Sl
5v/ijtbUYBIWcFWxnz5cTcgp4m2dgIYYt9B7/joqMfcE/sO5t1sV2Bud75MSko4auMRjtRtGKSWF
xnwg0ym+u7IpfB+jb8E+5yr/ysDnOBfS4gbVZMdHZle7Hh5lIJzDANd84udtnz2WwlyNg0lx0LMk
m4BV07Ndxr6YADP8tgMJ9N9yrUGGWHHuGcbNQ4CaFCEAOO4oB2AyCbOorCnKfFjxZSZw+WPD9CfX
mQQNt+kJaq3bEaVh3gb56ydN6UhgxNh1vuSVt59jQcpnKCVYyK9xwfd6uDQRkE1QFpoEC42CSHT5
XHTbv22eS+dCizbSOlFaB9rkSM1c70Qzd53e6KUP0gpDm2BasTKz8Tg7GduX4ST1Saqx5QOpGoCR
tyxtrLzPNiyrLDXBWkynYxwj/AI2B3RSXQtsuYxgz0B+oeeB/sVL9aoqZfdKxLwbHnQPDkXO8owK
6HX0tQuS6ikQRL47keyQYR/aQuYvdrFgvKIjj2WKSOz65kymFWfhOShkl/GB5sCjET0j9L0BedVX
jAx4H7e+xZD9wdkl4dBcL4LsSpQ/M5stkWSQ/76GdDMCtxGE6ty13WX7Jm5mNGEr5Lu9b9c73ZZJ
W2YErMMYfHf5IlU5rtnX9bCyzbw96Dh45bAZCR5jNdZdf2sxDzkrkKCqqQjtEc5Osa1bgDZbxlLz
dHb7nKCNEfIw4UjSOTq0drXsA6E2IwcYSRwRRyRcKLgWR8Mxhk4m9xj4dSbSeXB9lI6AXS3i2dpo
w5VtZpWANxHDefhZlzWvYGqbDwabHmKL0fa7Yf7huCIt4jlO6zkhCqNgAxyHXL9oZPCGI2IOIzxJ
r0c9vEsI7YKrKU+FPgAvLb9wedqVtRTQ9IfSoB6dYK9+xm9ige+11j0HisJIm3gUSRes03tyPNBI
eax3ZRvKudIE+hXAyc/PBqBO81iTJH4+Y2f9K2RdZBHFVVN2Xm04o5dnSDvwa0ikuo87cqD48z8l
dQrzJow64Yf/A6dBFzWkryij9+LvYfmuVcXFjvuS3Brnjiuo4t09CfNNcfXGg+q5dH+CY4bg6vli
3Vqqz+5JEEBQ3EJaqrXjtGyLUe3a0HXSpOFbqkwK1vb622/xdb3PenxTcWj1ZaEhONhu/Mm9Imrn
hJyOko5ULZN9uOBfsSz35JlviJq25joFwY4VKm+IpjCMGjy2QOF/U9BuAHsjWoIZldAfx7gQph+X
Jpva7peAmdkXoncmaxB314RGCdLM16Ydmi/aAbkY9SDx1YiWoeqRC+JdNRnqtoetR19N+FS6HWPr
cyEqB+x8qfFqJ647EBpRW4xQ1+vbpX0arqwclIypxSav3VOExYmupIWCL5LZRLdqR/iSn/lUUIrN
5WcJpYfXcSWgtPVnV4SpSejVICSSd1MS2czMpAyKvYOLtdX73nkI0ecA3Ni11Fu/5uCF87mMCqYq
7q2hg79OVR6m4PRpnBkjm85rVOKjc1c8RubVZo7H+KQcmPEPMe5T4FsKa5inJzeprSeV+whZwBJP
zadBubCDWpyY6+bQrINFUNfP+VhKdyfJOkz83y6Ftn8TpHvh4uXkgEBba4J4U3Ts9D1s7drLkzED
3rGsOcs9E/W+LywTRhxE8AjBCLKd7fGfNtpkEpfdsOiWBKAa6nfuQYjCB3kiFjArQO0xRtB7DqDY
yTL5EMpEFFFw1iXW9O4O0AWayPRbkIKyrBtp1Ixfz/GCzXLzVp202naAHbIPV8iK56TKgB5wCSIo
IBBarprrRx/cf2GI8o2zXI6joTrc+rSB9f1GDWMF/gByY/oxjBS2MxfPn+K4v0hLP6h0UG56Lp5S
bfMSl63d20yWe0A2A57LC94LzXCagvul/78LJQeAh2XvWnaHsk5TYDE/dgjM61vRfmj6UPB/TG0/
XwTAqFJwjCSSWXeeupxo/e0MeIdlWatcqDAFkExPLtK1UH/7hJyJjp3TJROZsJYF2DyqMznKRCKX
C0GFuyHMLP5/MsaeHApZMdXd7tGzMqFv+1HAhRjAL5HXYslimdxLXRymWATDlFGKukByHIhODITs
R+65/8cseYvwTsFC5NnHmGggnJNTdjZb0wWFbjKS+vqJT6ByjpJDsP0hLUahO0M9ED+JzxTFRucO
ttn+x4Iy25XEqsGrsRQPHmy4H5xvkJS63giXq/zpgJo6puxbZ++p37cbXd7Oqpvq1bRyLDedbvZK
pqP+Li/pCVJnP0ZTcB7nLlIWDQ1j55IK2M2vdcK1C4u4UsuUxt7odY9QvO5ZprGU6p3OxyoEdFf8
aFAUbMuwsCyWt6pW3KMoNS31miK7d2TWZdgXOrlb/Sywad76Su6BADzLFa1IAwaAW0wnxU5JVuvw
RWntdLabRaCU2JH7O6Fo2CZHv5AMO5gIEUWtyC6iabffdqD09zxjcpM1pIipd1OMdqvbvBgvHM2M
IAg5fjKPGYvXJAudhZ2d2/EbSbsC4K8JOfazDXxY119an7MjH6TxxFk2kGgRY5p9GzwYJX9ZwgwM
MF6AGO+brvKsvFfuWBGvHXmbDbkmKXjY8UxLP0ocYU2EJerqKztSIUNbrcyaXA4lZw2NqUQPGhrj
XG7cZhWXQ8iuYS6UhytjZd/qHxt/0chpZMFk1TaXJDFsGeen0tmaOKQXh+0edyLLujFbklaccs9R
kHwZX2w4LmcTlFF8Vwcjc11tXufuSadOIc95nN75kOutDGyQimUaCMA3aUdnYSOa7NERdtvYyUdr
hMV0YFeiGwM4fXyVL+0fB6FU2zZSgg99LTwh3oxE1PCWsPICYH+Scy6sdnm9Qs+R+CbJEXXe4Enx
cduCAk8JYgLyeOh76BKrWIxJjsPfOqJJu3lTJ//eHrEu7YQLguw0S5CR4zJZD8SVZRTxtcPQHcn9
ZNoOEeqMXaEGM+f63M8ESHUBopFu7SCuEDh4wm5ztt63H3tKQJsebzhak1q67gDPuTOX7BxwgJqZ
cDWceT/X/bRk8/UK0Nry9q8CQDwdlsrkM+I51F8jBdLI1bBJb8R3eG0Tm0UkMZKTQd258UWxdj0W
s893+BXdRUHZe8+DC6erpk0W225I89jCr/pJJ0QVSBdAuEtWPi+kaKoDpoeqgWSKHJGmSHwpsZyA
3ZSqN3d4JUQZSJhT9XZvGXjbu5mQWX/AsZXVmmqFyxDx1ZFqZLYVl/Y4lmLN7rFySQXJIjGtkF3D
tZSJ5KKljFHKWiZ8+oIjCBQp0HWrYy1HwrmFPAeVzTucn/rWKg92HUBOGNBHiPBOXM5fDUJV+P2T
7lkAnchlPg+OgHafYoTF2wsv8KqRdKhVtgzuHQ4sEufizoQKhzzmMNJGnSGA4UbIScpuKPRtJxrK
hDeTXBv6a/L1L+yHo9rASh1b2Z06u9juhMVjgk1VOMICeyfpPuDKtSv6S4+uOmEfroJ4gsmkah1U
i/Vwz0BM6Xd+w25oSU7jFemQo2614ytfba/Bas/DzyiS8XXt1UIkmmM4MEHdvHlteMc6tCIT+EWm
+w+lsvMLbZuZSFfLhHo4/kXLB1xDYOzBQEb8iePAH/K+YlwgBDsjNqt2nbaQxjw3KHCnIYXen4w7
ctGG/10okSFYEXsvBqULSOqduGiMOBCFFkfksXBm2dFzykSUHBnDMWfDmN1c09TkUbdDfGPwLlNs
b8AfDChnW766VdWgAoZQviS3edVLX9c8yQXNZ69tx58GdSVVjdJbzN9fj6sG1CDg8J80kGCbdETh
3Ts5AqwegepS2dfrwQ10H/VDuGqRSJw+DZYtfC+XTyzspKWO8AF2UjowO7XvURM8ekF5r4npKzk9
+slAmviseDLkKD4uaZxxgkkI/GnUwoM+QJVX1eYUfT2blHKYY0hCk1gMbFfFjqkg5PlOfgTwqq9j
amrQTVvA2IK+KiAY3q8490qIQeCOmrypZ8C+VJt8FrVxsszQBttnuRzehQo893efctSnz+2L6q4J
CMh5QhhNWT9y0OqTzZKJtXwVKfKfyfgFU3rIgR0stOdQFfTWtHZe0+px0WI4hKTuDU2teLgGUBa9
NjBtlVBfhz3haFz1CGoax0amNhXGgayvYcoCMBTjSRtTnQvFpqixsSy8Ah2UI1ta7F9dzi+JcmWT
gKzmHBanqRPQMDADbuNylT8t7NYQlRlch9cCJZnqmIWAj58pOMbbOGTQ4UqYJBmIf7Ue9GZ8sJ5g
TxZsHrNcku1W0yXEPTxCUFVIuAkVVlXXdmNvu0L0xnswJbQbwqL4PuVT4wS7kmEbY1VrBTaFcvOD
m+iiA0kEe0IQ/5lYGO7KaN/eFEkc/pM/ARozuG41cb670jGAGQlRUpSNLhuO7+LHaOjz/HuMQmpo
qsvV2wpYko4ZRRjZqh7tRmmN18YV+Ia3WZ6iYzd0+mF2+n56hzCvKpHfR9oIwInd2v/nGiEjY0MR
19FqZQcmN+dZNGgE2nCXJd31ujzQWFj1C3Hvar5SI4wgY00FaNriNhPRm5jquXXFhi/8NkKvnJMX
epeNe7tQ1Dpf4gklF52QlB+UqaDrrFp/WYfkEbeWHTLIEAfk2Bb4rpBD8fLcAVTijRZePFIWo/tH
zd+GUQHh8gSujHwldxMoNhF6EgiMiOeCvu1l0sym2Pn9GW9H9/D8lLgTzD/ItOphYvpomyY9L14b
jPRyikk3uKOe6m6eleL6ZiKJDANMAzEix6Z7AarQYHp8ZGSi2n85UxNcMhpM44cQ3J4Q2MWLoefQ
PYnbDMLY8gH+I3s1cDitjgblbCWLuQguax2GHIPptk9uEEbEfxdfDCDaOy7yv8FzNfSVu0nXQ3Y3
KkKtkxQihmKX9Ox8X2xCLNf1oM78/vRrVbNIgNV6lyO00r0UDQQUzj8DHmZru1KiS59t1TAMvzb1
DsUzgsWmI9BCEVg0gMh4Gi0igaa0O82+PNcpvnueQVhp/DZZV7XVWyv4ba0VhA6pPph8lx8q9zwh
qfzvll3Kz25/UDONiWi966EzyQMPjpPOMMz4qDypOpk1E1tEZzNRtgnmSVu9DHJs6IeLyDsvECxR
awi4KZCzIx0rdOgs8gsrTJdN8Kpyvff2OSv0cdOJmOny9WkGYKmHGxneHQEKRinQZuI22oXHy+MR
Wzdg+6soppX7VwuYRth/YgU1BwVCGifSdNQIi0jUX6q3HIFNWBTlhQo7+M9z/FE4oJVp784hAETh
nGyaxqKsd3n8hXL2JZlSenzL8xZerMbyfXmUnjp7YaNhZaqsmCqJTwq/2gK7+fZhCbxELUzJkFEj
EsvQ9xSu3yqv04fjLeY5P6VoFKv4zgVsgMgcUEy4ozOui/xN8v31QkzbhBzOYOP4C4neGDvbt9s+
qN/tFfmj4et00IhSK6YMmNySAAQexGzax9bcYURWAo/H2X9i9UtXUODZNuq+zPxoUiFGVryzsrwJ
R5AQz8Yneuvka/KJFBrJ2W+tmlJAYti7sqAhlMcoPeYgL2jzw72iRJl6gga8dnbue+vAMKidgmtm
dMzXjwEt1eTcN+ug1NNVQKcond++6aNdoq7xuLd8QOkf29L7DqQn3nW9AR+oO2SU4I4ZPCbGmZ5K
ch6JdcW+2U9lbMBtFaxzufppVksktu16ySVpajwjug5U9Ctta2wAbXz32va+khktz3GDtXPcIMU8
rxeVj1flm3C/r2PG/EqlKgQke9FV/GG95ikK/OBz3j1mtmpNNLknK/svgU+yi7BxeQd+0QZjR+Mc
xtjfJOT2racXZyOCmgoA7Jw1pnUwWR2N3rQy0dAFEe6BwQoN4HOOOglS8rs9/vPsawJ84gbjetto
GvlUvPWDE7xP0ANstRYF6oR5kb2KQxLZw6X2BJoYS2m/3OpcQZK7m2+Hx92ZwLUlJfI9Hl0SC9dX
sh8HROt6gDipCxbBxrv+imQ36wFIvBqL0Ch/WGFxHbP3L6/A63/YEcqQl66v/v/hLaTe8mzumtpE
iIIdUccyjMtIfoB7UiYU8fHUDPMA/VwHDIQhxxbA2Ve5w9JcmS1PzEKzYjzaIcFb6gb61jdGZywH
f2uL7Dxp5I6T/pMlrqjiCZ0F6PCGuAHuBPxrDazQV1I6rOOsVcmnKnU4Jcx/beKLgVzggsMPYbdm
Ja86Z7cEl7inL5qmFY0jp5wErUT+tUrb10CoihfgFyeiKRDnOQZyOkmP+xkSK3qyOGvkQlBLGl8v
SPBxucutwrKjSwRv042euoc5UKYcku6jmyolk7QaX5K9vx6QnhJL2YMsU6MWYL2Rf+HrX5pf/ZoN
8PSx/204gFGIiJ2RGWBed6EIGMz3SpLOZYYuRedUoozxaDbtU+mAWqr67McX1SvvM3wnzJX8Ko2h
Hig7533UWWYgfynD+uo7UokIYtnjyJNdarQTmFSDfBqMLBjiRFVeFYeR/bF5Gj7+JAq74P5qHIqj
gNAxxkNtLEwNU0JJq5Nn+Qxt7mkhnc3PogMIJA5wb0qlcom3QvnsHk+89qBvGYue3EtHjTg4r1S3
U/8CnswOlBUGSq52m7MuaiZqv3YQTqoufHUPV3WzB+NAScVpdKcjPh3oDWKPuhp7FxmH3EcubrNJ
0Pp06HOpy678fdJISEFHks3KLCX4BHxVtcyQ0qjW/5XvGDeLJ09ETrjGu5JUCW5uPUsOpOxlVC2P
JAO7Hcm4dZkdONzD40hyAgZcMWiLJtGExBrlw+YKU11+PEOcJE0iR9by47NYT9xZXIm/HO6AsnF+
fR3rQb5vPzapoGw3bRGXZLVAjgLEZ+28Sfs6s2cnNGMwM4RJaIFtNbSATo7F2ztz/DhLkVgIQ1FI
TUqSi66lpsGW6Ur6Wdl6HU7VScuG5Z/oZ59tCh0MOzeCedMkHZazHm7n3Eg86oKpiuIvu5DsRz4f
snrsloe21s675gbQUGYI1M3nAmBXlzihDo1/BLFjs//vDqHtMcuMy8Kj8dEJHVjXbKS4P8Gx6YHA
unUq2YiUYX8/L1z2ALS0HD0hsz61Fpsnv7DPeKCuiq23/d/IEK+TS6tQiUbrhccI11bTizs8LYuR
K+vv+GoTJQw7+LvPynFo3wU5gnOLyQixRjOAQXbLq5spjX05w0FDeTeocA60FBdoNeBrZ3JbfNC9
sekhSt1OY5upk/nrT1LRNG3tihzXyAlswXIElYrJaZgCxcSRvT+bDXGfrZQDyGkvGI1a6k2+9gOn
NUb2OyTbgQg8dVBWoZG0V7Gn0chxOExwU1LHisj1mAvIV0x0AslRxBP7g5E8+pnbJSMmQpBKE9CP
RYB82Eepcas0toeVVRG3lhdn+NmHOptvAnCeIWC6ePfHP6Az3N+uMQhoYVkx+Q9+NcnAGisOIo5T
yTm09aYSgoKWXaUqD5LuxWkBBTxSxqSQTdEUuMoj9vmtrBxCR/aw4lOjPY/+S6jWGPq1QIPSJZeq
R5PpR05QsdFy0BtxpXxo07sKnw04FJitaP8MQcasPJ1muBSS7zDWYXDf1teDBjFQRCPuREpdY1WN
sIVU3HHKJ7fvA235qpnP8S4ETQphFZKBpfy22XGkPiloblbtjdJ3Vep6RmHHo5MvHh1LmFXAU4TD
Ofi9QF+qYrbVvLROQhPCQsuZKTmTyy0LnOaHyHE/luoF6FxtAC2ufE87tH7sYHL1YtsBirdG5cTf
T0qOn0a6A2arM6ncfscm8Sit1f4PrRbh5m97KUsbA5paHWsdbaB/Hvr01SmTTVqFK4aosEuGep2K
us50rlVckPQKcokPG1iKcASSadquQfAfoqja+nXYbSzKUlZ0jCfE3cZsp3eHSuE8BbR2IfIJTuWT
mYRhubJ5A92/i6VKP76mE4IYyzc8ZdFi5EYstE/Tt97h0eTxvXarUzhLSJCQeRC69vZdsofPFKG6
fZFIQz1+OA5Uz4J/vTjohzRexYg7U+S5hqcR2QviGjWj0g5/T4iWHylU6X7Dc2TOCclzuIcUWNg2
dogopeilOVuaB7Ixrzob4KixswYLsCLyfRe/F3iMP0Z5FB+xw6EWrH7Avtbv2GS5NS6zCe6/f7CI
V5sF693FZT6w2GEbzv6U0cjRGXG8GymsWmFok272Gjj5JpTTrbvwvZB9FrAwMLIt6nbavk/LPxZI
KIdQJ1k5WTkq4N72uZNjaGJvtTjAr0pw1TsIaoS1jQZU375MjCeOM0nvPVe3pid0Gw/Y7xW7EHbC
jPzJknUwMCDArfoxI08Y7UzDLKCgWSwgZygb34uCZKHFxu1ORAZ1gyiFPtxumUiILQiBjuyeitPY
mlu+SIYOhyHuhewxKFS6dZIEcBZLNv4gifz0AsQxcIseiVMaozSkKznbST5+TWlCZg0oz1etJiME
iw+d8V8DSD8QWwh3cubj0lTPWbxgpgjH9vK1tW9Bjh7MruY4kF/4j3nx6vBIawvo+CjiTNKvc0UC
r7ols/capUFEsUM3wOHy85Yt9JhO5fvXEk8lsRk07VDeqlpVeopcBy41/6jhctjVuyU/nrhtD0Ax
BNs2d96whTbXcvIzx9+RZg9EYKDWk3yAPuUcSqpb9MrtzEhUe2ay0Y989W+qZrUnkrC4MLTeXxJF
cw5Nv+Z2ege6OOj+WNYeH5eqv3KpVK18/z3yvciRAdsNxCXAMDNXNZ1DJTxyK/egEuArrAwTmHZl
7Jwjm3WEUws30lPBL6ZVcdhPTBvfN1x3CzShlAQuLffu2jSWKnjqBclogeZjie908JfN6IjheQZc
5GPQZU9kG0WDR8l9LtUMMnCjxEdgIv7ZgV9rUoW0P9P1OoOeQ6dFDkztzk4NJ6vEdEp/mPXru4Wp
0QMyn3xInDh/csGNxsgelbjK1NaPja/cH0NuNH92Ak6sJ/WjpPQoiavJ3bDa9fAY8Eg+J0M4aMHq
hle8LIbuKRlO4csAKrxF34gXZADMOmsi2M59Ca/0jEzMcOIw2f6CFVzAGSiq//9iM426Uy+pIy0i
+vu7xME/tAFKfP7s0jC70AeuIIjR/4f+Z//MNVH7KAyQUrUEUnIE15hFaTul/oyJLeT8YTEjgEmy
i/XFMZV8n+pJlZUzCRgs/tCkYbvCp/NKRdELqZ59UUWi2tMd5H+pr90pmTiFMMGarINb+x7JyEwI
s/vzZDYQKk/XFnmNYHwLCPtys988pjVhPCLbbM35PjhAJMxwqWYZ0doGxJfYaVDB/NE0fPO9KRuC
fVXn9jNbOMQGXmh7zhG67vEe30S3+Qo9hqKeHfQ1wCc1gQQjG/zpnDssi0Rtj43Dibe+tE4aRsAM
H/drfd3fixL6zeITv14FM2iuVgrnNORUpn0E/v0Jfb040fuZAAlDasCPbdVGftJYY3RZ9nBjf+d7
cX0r8G8IVzt3qkE2f5nkCyjUCraUvXRNlqvQsCG8mail+x/hAiGv2xJegw2Fih0dc4/mkDOmNC6d
exp7iH5n2KIISFa5ykQQdP148cmCup8/sIBOcqoWcGvv31/Yp7qGXeWs8ySnWsv9GCBn2B7pLz6z
vxZC4j4j94diPCTNcxBhAVrJUr3V/KxXPN4oldYj9IWhswkoaIkoTKQPJOL6wqP69oBkS4YDLjST
ylIZrG6DW1iaLFd/rvvbJam4yROCFPfI7kKXqvqwPeBJmdKiKJatQGicwM3XsiM+Ok+Ha12dQUuQ
fgb5mP96ef1MI7rCfeeF3UAB4sVLVHOvE30Rc+1/etu4jb3fkOLS1N6FIikiYSwASOh3U+rPNVxi
6nQjlAOuwPTncVm+/9gkVCdJWm1mwZ+hk11yKIxVEFENKEDQLakbPg7HB8gBTojqbu47LYPM+bvf
qb/EHtN5Fk0kMpAtnfxAMUdJg3U4rGegGrqNLhZHxL8O5aF3qAR/l0xrE26AczDSGfEOfDej5d4M
qhlznJ5LTMcjl/ZjzqrW6jFJ9OdW8Jl/J+S6RJmEr5hO+Wm55Az7qWsqk+OnG1Z2xjnFjROLNNsU
bg1DAN8w5Cw6nJPRjdhz93UzITMMxbKSKYBEu5XOfxne5Kma4VKFBQA1K0UOHqp3BKsrlwZ+ZeBG
zTGQW8JK2gt4xI9jtoo7fc83hx4kBowlsmpxmWTZ6GpdDKxJd8L2H+tXp/dX5wia2R+xZe0Uovsr
ppj776XgQVOSOaUPAPUI2laZLUba9i3DIf35Hmzgm7zR0v3T1b7/qg84QyLnUIvYdzb4iYqJqViv
ZG2dThvUayNEDH+oFnzwI6KMUg0CJ5C1Lr/dCFrMedXyDlCzADwOh1IQNE6rT61UV09cmhmuEXvL
PV60Y9N+H+GNSrdgSl9m9gKmzbfPV0fyEyZpvV3pqKXdyGWuoMdU9tqt54ZInQy6u0FBi4J8lzUH
eUsfelEK7nnNDvA5yanvNVZi+0ZQ2IRZNoXcuPa4DhbJefsniO44ALM5jCJtoB/5rWGAx0cjhAGB
cnt2ol6RKUz1g8fuCMfgyl8bRdd5Rg4PFH29s0G3EQxxUNRjZR9xd6syLSeTpS7ceZ/xtqmp0tcq
mKPJBrxXIh7uzH21MgaJdeHyOjIpWgtcaaLLcnUAxBmiCfJ1587It1fHGtmlGpCNxAYM6afqmVo7
w1L3/kql1tHNpOqnTf0qk7bmZfDu2CGHomXNr41RlVPtO2LdiqHxess9OYeD6DrIn8qQMuS2ipom
hgnt8WR5f0oB39l1zG/kmV2tQ0LkjAB911N+mwwhIRjjRv7neFlEDjnS09fsvWiD4zdMaJuGO2TF
4b5zJZMKWqXstg+GUsrQu5KyzWy7FcYebC0rkSE8jp2n8JwqmI9NpYyXHPxeAZSBWQg9sYQTvRam
feq3mt1oZLcrG98IT4vqsaHgn6wdfnTTyizczNSiCq+SorOLjEm+b2pO/ORRfhadBkoMnzT6We90
X3c9ZGwohIK+t36rO+OGTIQ9v463nwVnUMIaMc+rPwT0l04WhZzducBsIbJilHRelbtrJ9zVP7S1
dyQn8KwGL7H2bWCLS+bLfywQ1sW7htpSYBRBviq0i3iZ87nvJcB41gnWjxNGZZnjafwkS9xw6kF0
VVaqez+gJM1uLOraSB+HxsMxgKM0vsavWwM3x08SPfTbbW7Jvfj53LubwciLS4R0AU/yVZUrNHqL
ior/t1K5QDVVAzsKa8j4HNnk+Mr1oUiVI5VSCNhUhP2TCEK4AFmaS+7XJaDCUTYwoIvCzEshfJCQ
2uL6sQbRY1iHKEq4+X79l/s5LaahVulx0J5Q896SIQBvPSmJXc2Dp2RIF+h8/7gNntTm/epcmgv9
mmIHLxaEAeUBoxdEHw5CA/MyWARrRYdAjbVWFcyPcLAMLvDCUt3ziJUne9P2ATsUq5s3HCM7NUs8
np0sTTVhczKvl+29hX3ENNChF5TFVva0qkyHjWH5U1nq/rEnlEFYRT8JQoyZGDgGizojj+wJbvVP
wyDyR9S8thssU3NpidhDT+zOmGl8FVrnP8co9PznfZmp+gJh1sbxWS3rGY+7MWDoEliZ4zqdIGfn
LRvRBRhX0hwdWKj+RIx3PWmUtxdSZtoDZ+ZfQ7GsxyC4vGYwy//vfAiz7R7yV9p5lWy+TTMByDTt
E+7wSZCZIlTuFgE/ppOefLx7zXg9iyvtTICE9zdzwEHuOEEU5UFGUjat1Q77JQMJXmlMcJt7spKt
5Q0mfDeOyJzeqFcMO0+foMUmf37W9T9eLENCSCbnYHDjvVvkf2Bb0o/BXOa7sdMN0tdwxSkoH7VV
0Vv/HPXVF+1qw1ZwWpN+iEtjoKHcTImyj8SWaGnaOg0sviagMpogk05oXwqchC+7Lck4UNIoDP9c
Inzft8ZnQ+oKY1xgMFwNDd+I7+LgMvhn4FXuXFYr316pMWb52iC+zrOwUk3CpwMSTUgDFEKRle+Z
dRywbm/0sNnXQzVkreLef2d7N04ok/732B5mPdHbp9LOJ9hi7b0uTxIHP7O0xN2Hs5+j7Y0Z+PFG
fIi5GcQJ5R/jf82Ex/Z/XOxTHpCofHD+bgQCI7adqDGAFnRMyPp0GlAVQXWB334qsiRcESxSB9R2
G/Xda0z/nBCi7ClsDwAc4SbtPbfuGFlBCxlM5sl4lL6aty8hJSz9ZBiLcj6ows6EgNjKLW/ncRxE
n4nD9aDnP7RWEkXXAKnFCWENNOidl8CwkHmrByJ4huTvepbUaYiaCYuxayQH0ig12KxiKwK77Wit
6NyBNjmwBLiax5l4tdWMwJb264RDu0DuFjEwzOP5R4Fj/YjBGQFntqmrI3DdubNPS4Y25DrJuLEC
Y4tmkCZM5jm94SDA6hg03We4XhhcOPN1Sf+J/QUDxuxX8P3MigUuyotBsiusk+U+fHuB3cA2ImJx
e5daZa0EK48lrmEogQ77ovAKMBXcleNNE9+mvzHQR+Jm5JlGq3nQMQ+wqDkVMYYzIaIaKFtvSNps
AyClyY+2unz43rX5V+PzitzRxpT4Ss4cisZijYWneq9KYovQjuGL3rNvFUz5fN8bnhUr6wArAGpS
Uts+CiBmIDuy2s4YGULkNdfdvyGJS2NJq8eJQJRBl530wyW+xLoqUwyqA7Ek9BWEilEUczs+VSVg
pl2tNBm9WeXs+aiAJGxrdqB5dzEhDB3JIFT0270dM/7IhJK/sugCBWuA97V3pYo35sjNTHQIj2H3
2/8D3XG5iU0lcO8MYnK7VoCmcwP7aV7DYJuuDPlaxl86DaESClvl9Ht3nvhzigCoucMHluxbj55/
axpSH5ZjCNiTZwf/6HjwJawE2DGQeRUT8HGgvtrAhlIc6aEjtXBHouMX+8asXghKW35Gb6VTwJTF
GfzM9XHmeHrYkfIheepkuPrECUXVJw8+SatRe/55JgRZmV0tzIBQ8X3uY7+7Y6BGcc+DtcQpb89i
2zCwkipBE+nP0d3OBIImA8h/S1vXV/hiNd0xlec9QAG4DaBkSlIIP8TVO6+j61/30hewbDn3B0U2
Y6qX2xgpvEX4dOAXQexFJ3QZFegVWCFiRHdRNTFviS3vfVP5yIuHwoMhfUxlx7fBJVIEW82rYJ2m
KYLnXvwA87IQjUogEDX7GpCm1XPzaBOJO/nNZh7XYenQ4Fa7uFvyW+0qIO73sAPASFuOQwiz2D9o
rYIhAsTr2DOqY4NBGjc4HvSfTP6czZKJYoYeHoDyc4qM2/zU3boNH5IZfCvc1iXkn9mDLd0Q/ALD
43XHL1MR9NareTe2F73u65Asf3ItJfFOlCv6+G+laUf7/PKKGfpRzbDqQfgdMnR/TUGR4FKNOrl9
+ZTvZbYMy7hWHfHl3MT2q+Qa0+GFSB24txp6wbioqApRc9seKvptGYhrKZyKAP0zSiNYcCJ2OV8q
J0ZTG4W1Y4Te0xuyfsanI9hLTR0847decNY6czTjgsZR4sVi7ZmePF0WrJvgdpxhliKkuHMSl9D+
6RYSleHcQXC1USlxxmw1OrZEO3chhEImVFNK/uckcr505+JwObxcaZIrjDyFmmMNv2fTGmuKUlUR
ctiKIqXzQLY74jKtYJL4f5fX6B+0i8Ce2+7GTGctDv7SM9wl5Z24/0+M5BNE1ISXVLe/lDn0GNhB
op9R4p64io4T3le5+sFxvTq+8kHDvSyyIEuCLO85F7ndOX1D7LU4WHbRGODWQytML25j94d5lmwj
V7I/DjSUN6X2I4BpQfLOs9/rMkuiVope4ngiHRKVQPV+UlEVaO8chPGhdQV90wGGMotl1NSPFKiZ
IIH5xwTFHB8II66KBNz0QyLuqHQ4g7Y7UadPAcKgHxv2IwVs0P2BthMpDz1KVUSsu4oterL6+Xjy
dZJOquGIWe9EAy+Rrx39E7qH76qf/ibB4xVe/2aT6Yc/2Ci5d8fRWjzIjwrx1IH1XkMG/gA1W0WJ
BYVXPeLlo3afg0XTJp87rf8LXYt5F1Rzxdv91aML7zgMV7GZCoGu/1cJ6edM9ASAJhf8D684aiUQ
AHmqtUS8tieFrtoKGCcyf2qWHWp5bOS59Ai+yrAE+z0jI3uQ/egQAij9Xv3KyoAq9UyZki1H0xGY
EOFdQ4E6GJdLE67LhEdy/AERxS5iQLQMTWPoCD9iKqs/KdUL5aoFr5CU9Qy9m71XKiFSJJVvYQV3
h/6mYp2l5g9Vk8M8o5Klx+u7rHidEsQqILW2SSqJCLlsjZ2aijqK7PeXj1RLOitstHT55Itc/dLi
lW6TGY/788T0f05RtGE7r9Z5TUQ5AyY2mKVGnJj0RkJJE2L9PPIl5B6/AJqTsy0xz7KK6yPorRb4
yUmCSmQ5Wnl7AcNqLCqTFqcPxpa4l+pGo6vuIPwc1XrukAglVnSrjfYBKvlpM81r43jPpCIjECiS
f2diOH45s5IVQYhPIFSBnYp06oJRkVtKTLFp2r6wdSfEtOAg1ca/kT7cBBJFAoQMiLgo3mGqt1+p
pAeiUxQOkErTTBl0PK3Ae13NQr3UJh9nCT+8ezAqDakLfjBwbAA8+JPvNlvif9DSkYZ1Yh0E0fgv
Ieik3HW8waqGXF8ODUc4m3GXpybiHr7v5/V1e9uNytKcWaaZieAOR2DqHSLgILIwVNW/JVhoJcHI
Tz0so2MXnZMps5ldgzQc4byQ79J3KkhNzHnM/umyTqgwLmCEPELD3pFI+9xJo7LaeuC9tXubq/xl
C3ZCIgRp32j0ajavy9v+sQePcPvYGSU88qwAd6sutTJKJ0wIJItdytBInCBTTDYl02vzEvdTa9ls
wgg23CusGcfdx0AyMo9CGUx1UcFu/YeYXkaV7UQMJ3A1S2K2sSbY2iu6NSLcCtnWKWaaxZzP0E6J
mEbCfT/6X9boXvFtP/kQTtMpSeQoe4SiSNBOuaBFiuU49wlnmZRAsjH7jdCPqukFzR3KMvUJTzS1
/dgNcddKBy7h0D3q5zA0GDyfcO0MG0mY6XdrFr/svp1DJj30YvwKT5cMTUvzpIvsD8xvp0/TkJH5
vaeVWwbFHQiH3C5/nLkt9DrbshJDz7WF6Kry2hMzJCiRQcb8A/kHGmW1xwiBKIOfRpeQ56R1XS5L
kRpAnySJpJM9+wYRopHClpEiiZdPsiDRjUaRX90Gl9zhr+gFjP8iD/zXd2LhUZ0+0mK3/VP2I1w+
HtTZ25e/Ws9hv/ATu3Jllicmsk6J/mt86R8VwuFSyPZQrNxf0b9aI5Zw/v9fu7rdvKe5YUp6hTH7
udETJ7MvMb+XhBDIcix8a+Nd24UZYLPFHdY/X7ZPgrvV+uEz+4Az5FfAIRaroIANxEYjHuvbh8XG
39G2PQ9EBpTksOROw1VPfBH6+3NO6DYVBtUxZPTOK7z7OyZb1yB7IXX84nNeF5GKqBaTFvxarAoD
/g0Mk4mx+zroQVO3BABEAUtcSncYt4BgIH100tBnH/O9ngU99Sody1MMvtXAjcnUnIF1aEc0B4nN
sC/nMScZHeXsOSC8/NmEP7lau5BuNwMBzb5leooA7UIak3ho7SworcYXk2CPKoV/U78eysvtjseW
8Ldu2KI0rrIUmJD42FCYDPJLzLnSd9f5IPnk1v690BnRPo2ZJ794GAnG5MQcg6aqHFPEGQF7ZWpW
WoTNSW7uanGXuLljjVowYc1pwPoymDj4lJ2ba6jZw4LS9/xPGH0SU/mq+yvIQgs5JzMQ81RWPAb6
+lV0qYU4Cf4L+ABK2AJlbjIhif/PnWJwXewnuWKHgbDdqkR/xIZmuB0LELQfwkfScqEX9QR+TgH0
KdxFpVOgRWi1abqRbf6mEaZouRL9CYHF64N/cK0A7qtN7CF2Dqx5Dctz7Ztq6GTrb8tCPtj0zQyz
GApXY/nz1JIlaadQqcGS7ZxvGYdl/D7IyIuwcMcOD0AZgtdbZ740WIKDwaxG3kswoFa/61oajOLX
6HbHXhoZHzP9jBy9rtav6D726nHa9kdKpEr2pkdT27sFS2TwUwSZ/mYx4pCYbMAWhX5Kv/80uXCr
I5YM0sWAWoNjstYjPkGxJ0+4xjXCECoDgyQvR+KzrTsvSG4wQbz53nbZjXw95PzveScfwwTdtYhB
iM/cJNb/JKSSwG0tcraR4gnuEXjIFDgjVZkJkmncjb7sP0oZuQNnxzRbQv4K+XDRUumrWsgokhGi
QLLhU5TtB0auE/A7JRKR5N/ktFUZyumEe5XF4qaV9lZIPWyoAUBw4ucdFOrMtrGMMXHgvvlvOS5U
Ylu8FQOqOj6sqo3jmdzSrbD6vn3dTZ+ZqDQcNJLDt7uCQwPm1T0cz1/3fbSUQ/dB76fAnmyRLFKM
w6QJs9Sh3Bg+pZuquBgthnb81N0pnF8bmSO3urxyJn7sFrnz7g8d/LbWHMlXUtkGtLMT8o7P4EpN
5U6BsmYSQEnmIWRGjWUz2Wpfnfil0hxxllVXgUjSe3miUvuBTQwixIjtgMhqp4NjoPePDqhYAoZB
XPP6wrRKqK6MgaAZKfWjVxl7cnJdpDiev3eA9UYPwJazVi/F39RaSEDGIWY2EqzAzFhXly6x/MbB
HYRFq5UPGEejKf9DnBsqol7IP6dcCxiqe6wv9VuoaXOlDSHZBSQ+0ePRLEKFhDpTYjKOmvUpScq7
L1dVHibKg1dQH9yc3Yt3elbcEJvEkobFJHOnkCHJZQnOuZuGr3QFm5bkxPYk4yTrVS78G4l+WoQZ
8v8xELbxa4v8uQ4zD2ouRy9uA4OoyVVGwIEWSRIVa5eTL55rME6THJ4RimxpDO8QG01gN4LGIN51
Duv7HXmAAgc/MV7xRt5scvDTbOBCZEDeFqYeNdg7xDnU+BaT18JCoD5kD6AjR4RFO9WAGXNozXI+
11XjD/PI+c/WCvQBUOaEtrzvaYrCu4K9MDLpfNBV3MCoHfIdlPll23Gr4tDwsDE4tRu1j9eI76hb
1ZBWih5ACUgtklj2Ux4Ce2YPHKbnE+r1q3/30v1zePWFYTo+fVl3t6K/Xc0F0oINKzs75YscSppl
0eCQEw5XUkjrexpYUVWDNtlzrZDl6WUpjIayMiTEiMyNcfsNnRh+JF8g3VRi3wboApzRpGgT5dBZ
Yc11FqcchxoIGGyfFmc0YIN/bDXm+CtW4iz6fFm2FPHzdKGBp9OcOuTL1S51tLoKXwCUD9Dcpmez
z8Glq62csR1M8sYDeBicg5OMYZjA3hU6U2H+yLUEM+R08QlxJtYxj1YRJHPt+97OlpIrqmKKL8aA
1BLm9dEgxXh1oyriC99rgRh3mdaZ1oVNSJm3Y67scwql/phdINbtFtolOiSQaTIfBTwUtVTy4nhg
3XDRQ0qo4yCA6pKsdxDo30E0uXXpjshBWJb1tVKDqde8OZyGWfOz4s+C57PIfegZ/ph0DS2/Z18+
HOPaUJKKP5SF80Nc4wDtFjePx+o8TXW6Vrf760oyQzK7K6JuTqGVjVitpK8pfuB4aNqtHIfDC//j
/Ce4SIoazbWcKU5ZA4ZssZvV6yw7YIPz7NTrSTzJMRLCU5F2exwW15GzC2ghq+3oijH71sESUgo7
/+nbUwI8prDxjsgGUOoyVhgn4YFJKwFdahhDXgpphwUCVh8k3ZbMVR03oka58N2hY1NCElpESkiV
kfVpIAYkerEba7oXV8hNTsgdL6V4kMJ8bXBiaSjSbIeZ9Z4ysjpp6sQ55GWOJ/ip378QXyZrTAPK
Evv6op5Ct/cnmytrA5W1nQI8wVE5f75wU3CCpWmU9jaWpeaFldlHkguM7hKBZwy4WKdrJMJ7NkkS
7mXlt+zlae9y2e+8rfppFwVbEhaV8tip+AoMrHvbz8eSCg/4u5ONtAgoWRI6znAz9yI3y/pykec+
7+39/cREteONneErbMT1W9cWKK5qQnnJDfMrNcNTRLD/4TGGeU0PMZFQpXDaRot+vqF6mbhyEmKS
hatMTDv9mZ6vLye2Dh+7VxWHDLeVc+jO6PZbgVrRVmH5ZThy5M5Z4GsX75T4XJQRZDInhO8jc7sB
R7nQ2bpziV+z9XkBaTEgIhZUVkTftG5boMZN4CrTtUh/KVxGmlTMHlRr1Kr9NXeTWx1aXyptHOLR
ilPfrlZcxNXzhii0hkRZlK0yFPwXi7/mj7wxkhzPse+iSpeJyt3363GNM3KFQeXSyOEqM0KXrZCp
DJRYzF8KL4Pvt4c4F7h1kEmbqiG6uhZQ/IN2wKa5AoAtlGlsb6RlRdi49MprlbivLuOZi6pEQg1E
VJw0dhQSVLOYZEsvzjU93L8+orY4gHq/Wju3E1z80qPLmnOVBV1IQZ0oinWd5Wgxf62WOMD0j2cT
HpdeX/amGPEkCGo1Wqo/2FMgjPBhb+nm4fNHJ2OpT0VvIkQ4kajOuzR5JY1LOQ1xp7SQDSSs+/h3
6Ln7/T3WJ3eAIDMWW7qBB6FazZLgZ6oPAXptHsVEMBCD19Fh8gyVOA48c6fNIrbYMyRaImYcxTSu
dbAY2p5IdwG8AJ4HSNUzGazAeLfKiPIcIHl/ntTNsWjarTopC7u8ywWZv5VM3kMrBC+P7FmFzdkp
TMdCKC5+Dkg/QEodrJkkMKkm0hpsRZYbTvTJKpqGPZT98IYuroOajEAYMSz4tx4LY9EEJzwGbZYV
yJq2F8FGmz+RlT6WcImlxRFYOFfkaNyAULb38tQdCC/L5ZbedXBcnC2lVCl9VbDc5mnSlwWELXU9
+Ml3FnIK2Ooc+w5IN0HiiPxNlwDnq3oGFM6YINaCYstGDEvscS1WwNABRO8HajM4/SaGGeTHPdIu
VULNbrDmuIJnuaDOva+RAwbnobywsV19mG5MYpb9cSZlIDDTpo5WNDAFmo84ULAONFlkuKV0ntp0
HTJBnexC6dDFMCgHdyK0iuKsCXDzEq/TznCr4cnel9c6D7jp2GeKXUdAWdORCC824pzRjxNGLcdX
2KRV2BmWtWrIr1Qszc6h3B1MY91S83CsFvzY7o0GqjKZeIzVnvGJMdvZzXGDEYhDOSy2uS3Fip2J
UlE6CJw+M/+J5tZRdFcz46HODLd4wrYZJIWf3yhcVrMZI2DvhrMNZjwevyh3tgYU41C7RLICwkNE
c415yYIN7JThxblxG6QvNbW0XgB1gzwzF2OM8mkUsctLcn/Fgi4HeiD3wpa//3+s59FVDxIba8b1
7Em7Fju9dTH/0JSB8inothXtEWVb8UwJgznmzkSTU0eci9fQwTwRWbKvJhhioGLGfbCe5tK9jAun
43kALdX0YGeyF6j4f/XKrJKivxzrN6rex2vb9EjCGXeBzaYLwBqWAxOWbOm6CJsPzmWmTLgBZQSv
SdDR/jQZG8qX5bXoexPvHEZ+/JI/rs6nrST2SPq1x8yMSepiAddAq9LQuss/KGwAoKAUh9GAsXKv
q9mw3V7d65T90AI3U+GchvUTd+bIK+XsEVfXwC2KORHI70+kekwgA/f6usz0MS7N/nJ07uwuMQ+6
NeKYIvdSTPRtSHnO/+zmHGdNj9RdN52iPNLu6+JAmg+1UCOW9UApsFKzEsjgTDV7AOgw0rOZk1Cv
mHUxeyrjLMAr0AW5XgKmoLBXbekuOLSbNdlw8nYPyAUCNs5y6949bgB6SMplVbEJXQbo22Lq8FQV
PiTQArl9hDKMC6xPKkoH0EIouUCK0Wn4tvrucV7lw8MgfS60Zli9psLVi+O4Nn0DcLmkNjwejZpY
bWB4WffL1qNA569ruHOLdY1dQo7CuAqSywKMdrzVKbxEZnNUxE1JMA9nrwpSKhI70h4FKLn0C5lN
YGtFRIt6aTf81IeMG0dey66TlW7H/7y/CulFz3LjLQQwVi8ZIjsLoZb2JkrvCEPY3lg94qnz30CD
kpQ/y3wVvyVN4cuc26+fY7yQPrBZRGUqEimp4FZL/2wzPfgp68yUyxex9Qdts5bLqb7XU0Xt4e2n
/i9ZXfBnDVj4SV8yyNAQZB/adg398xPuDUwPh2ENO2jEjhoJ7nYiHk3Tnu9nXFifqfQ0fEGBzTWy
AJiTIltmf7Jsy1GYjGb/z5A7gqI4lD72jsqHOHC1MDWZCt4Y2wp96ELHs0EP0RtQuFHyUo1N4Bq8
SGJer1Qfyd5vzPD0tXf1dxxs9JYCMB0pAg2IsL58YBV+f554adFuyZ87bR1bFMUBCspljQi6mZWa
caH5+nHS5UKuR1lLGrzS6iujwSnLEJrUe1tH1/mNj/tgfqt1dByNeCWKP5PgcX0MwAD6u+HdAvGH
hQlG9Qjjj9KL8MtnVOrNBWkoqAeagU6M2BZADJoDWBS8dgKKDtSxDdNm2FPJbbXtY0xjE1eEyIeR
xYS9k8et0ydzT/nZ6xVp3NopmiMHXce9GQvWSeIdIgXZD8Bm1Od4yNPlr4Ocsyz5FBzr1hzZrth/
+TXxtSEjuTNpDcX6JBpaRSHMgmIU4cr8lgbOD5fxtXOiHIkF+dN4XIT8yzYHk/obb0U+vR/LJd2d
/6d0BIrJ7KPqZjZDrUtSgFOmepN42Ea08hd5wepMiahsjY9PpJJGotwKDJWr7SHbmIWDtoe/JkfR
6VNxXw76F/wLFOux5jbpjqjRh/NWRZbzmiJWqetqtt4fAofWrNRp9XX8XqG7WMFu5SwNYbNgmC7b
4CfBeJO++ctIEXR2BSRdRUaMrgszcOxd/wDV2jzNlwDn+eBcF3o9e2/MOSyCTqqEP/hUz6fRZLxV
40fTTNQg3x70asVTHcXYVCo4cdYYHL60i7s/JVWJNTk/9Mu7nM5zR+eohO+U4QC6qeTwmHo78/jY
dlWE2xF7NuHcGFJYz45ur48/XWN6MOIWDFQgjTLcvfh4S/JO0nOUDeRr5qOrRSPHp/+PFovOqXZr
rU6pQqnDcfXjtbJcbxkiju+bNlvVoIjld5BUzXx6a4MVAyNcfdsGkLPcbnjHBgCF5mpoRmt8GUrK
EY/FGU4/HM+hHZf8XAisWYdVHZgIDdDyEPbHyZwLszHEW0iRgvOVvj2V3vYpHnnGC7eEBeDgicak
7YlV5ZDy0za6w7MpJgwsbb0Lw+z1YjD97eHQtFiLvyrjKVeM/PiZOH6Bvtr0d1q2GwQHYNBRW7Li
CPfoXEjs4S8WZDkijtRlWbNlGdmktcNcrh+UNCYakx0hPSg6pjMu/XfYG35zxBXA1AkbV+sb1UBh
LxQtY9QKHf1XAB9H1mS3YW1NgPgIQzfnIk7qEBDSQrpcPSwLxBtG3/iCghVZfSNVTbqRVJ/IYXnU
ydXCGo0KVtFHC5jlR05HTyO4ii4TcmEDmJVA9mh3I0SGRJ+V5HoV+gcQ7Z1IEHSufZkFeZj+SxA6
/84agnXI4qGuCRlsGDKvGOzWdTxh/BX5MRKUG3TGxEotuYZWXfNY/fmmrxMjEtnQq+HgnVV/Ere3
Ulcg3TXtaRmjVEApDK9fnaTv7M7n+YGoYXa/TYBINqOIsnhcZDmAahL/9Iou3LiNKJPUPqkXdeTl
w5d2QpEV9s5UcWaoV2p7T+eE1QVt6QvmsxFLrr5zsFrNYU4KfMXWGCt5+X98S82N/TkQ79x2nw+q
Q4uI3/HRyczixxv75R+TWAzpPWGyc4M6QJCt/VVHzocozgn091U6kfN4/qZVuA3yYS1PxMl3X1zr
6KepqrbP1BQDroB/y9gnE5gOPNyDeqNbp3s5dtmLq2iWXPdfPsIimZe8IATnZjkmGhRVsRAnSqCO
elzB/QbHkQsXzCj9MPDAMP//k6o+vvi2aFqhOMfAdZHmOglu7D1vk9+FakaZL3m9tYlSwDHHbagG
eVqRi0wpSwouXN87oTrIH4M2diTRSqvwdRReBbhWqBD4I7neWQCG85il7JwNVSyl+KmYi7Q85KDe
crj47rBjn9TJVZCTvSNdbOP7wnZaQwZsloBbDn9AS6JiDedO+FI+0P9mhwBrwz3YqIXssyfVlBuq
XhYXT+caKhVjqpOu5pDMWdoeCnsWDO1BdF+c0Q7SMs0jiRhwYzidFyrY9DmFCn8oAoZfxXU6eK2Q
/Uf9I92Q5LUVf5kLFgx6lF1oo8a4Ua3+xtw5a7sdUnYmXdyw5y0+Vj+hP7psjlcE5lHGVQgvEGbr
MjU/UVVVVpovnS/oAWnyKVLJMlwsgTMlN2aj0c/3s0zT6Zop/UOPE6o4NjxA8NGa2zgHcI1gYn+L
DyeibCb3Wwl7MovijDvGzl+nVnJBt7sUt/gaxc1CURs1AQaCJ/KOU9cmnDbBgXztqYtTdjZRZ/O3
pp31S8l1TzGC1z6uLvbrMS6e3MJE0+wf5WQz9Hg0HOyqhYUF6mCNzbi29CC9Ndq4frwC/OnZernh
B4JAUvto4EG+4CUwAExhdYzFWDSyDa+vjiAC5gcp0PQTQnJQNTZPyCs2ANvlEFEHyaObSPPqDtS7
wHC29YO3A2AKrish5OtFIs9DBVXoVVGBKvYfRyzhrnrrPwUVNmxMMre2KhwGudegLYDTEmsW9APo
dx4zWaJEfHNeNC5uJoou1AHzUBi8OsOmmZnX/bK3LKfCdYiqAuCGz+381qp8OPN0vaSwcBe2kUZk
kwRNZJmmEQGQf5S8B9fPYGSKMvPanpwq77NjuyJKuw+L/LhOWf3h4JybMN4c+gmJcqevnfWddypw
MQ4aiIAnhL173MZD9CUJWiEdQd6Supq07Rwh0KStKvIkarxi3xwNN6Ry74HAW/OLJMR4uyGhFcF8
Ui3wECQ634ef/nvDcMO+rRnhr/D0nkE0rFypTn+4HiomH66WPn2BI2nCvCUVX/X5PzRjV+iTAnhP
Rqw3EfCdfDhSDe7mb84E32lGz+7A16uA1yxwGfs8I/RN0xSf0tHcosMs7EhPTw2K19YAGxjf8lT4
rhdWOC64+lmaftqekaELEQ1Kl10SUiwskQnJskZ8kQCdsNQL+k9j7Hn0zuZxkAXB7+AUPt7LQ/ma
r7lq9Dt8YpuTTQsgz77ogZtg98pe35Nf2YsHnCpGj+zPWq8TSm7GWimT6Az/Q/qOZqQzn63kTarW
ALVWybgW9mhAl5cj7u0Ky/H63dJhBpZEUgJRuc9iyjepUJvli1FokSgE2PulRMoeX2RjCxJMX2yG
1Pmbwezo3zv2XwrV6FTmLVn0Q5dvu6bGSxghukhYZl0CLTiZO6u+F4pBfyIwyWYI2ibZh2XCwlJo
lMgZdGy/J3dGAv5pA7yRw4glVybobFSv+SOsfMyN4CsITqH7HU4ffKSEtKdsrvQK/JPIgopcPvlb
slsRGocyb4HK1XEleu3liddH60wt6rm/PdmTibbMwZKeBsvAbpJBFtGpd1Emt7WAfeT6jDjlj5AC
D6k7R80+/3z6iQBBCkLEFmCD4ZEO4zocRBke/FmkKlAJeV4/qfLgtCPc1ngQB8Sg36b0iDnRPIR7
NxfqiZsS3puPAOfyDU8Im6V/3AC7O4/yNToq+aTCHrJ2L6vzOslOxA2mjgEDKCP+P7F205ILyfkD
tRf0GCxI/QTr0nOnR6daSCgGMQNVvE6qepIGnCIrP83E1UE/5wKOO+sfQzbSAxRUiLvs/o6VFwKC
em0hxSDAwWXQtFy1+JfGvasYPukBHalndIOG6P+N3QkBIAbnqTtLFMHHgy8QderIngkAxYk/rcJ2
2ObWrGiNB1NNd4uTife9KqXtv0W7YfZMuBe91Dymq5EroPXvrwsuujqkwLEaLUbr791CGkf7GKbH
Ne7BzdsN0rThhLN9K7rmAloH18wJ9GnndUOtvu5jaVA5yuI/lG6pQowMBe4UzTUp3j+RLYiGZuw2
5+8vsj/EtROo67ktFfOToM5+rMOTcngMub7+z0qazphrhMSKgzx3PHfQr0zGOWStIZEDy03Eyppc
gp//rE+IvcDkN+Djhr2RasSXQ0GE4IV0l2nrO9wikO0PJn6TyOrYA/Z17UXvfKtByfd55BWoicRS
Ooo1nAkY/TzcZfZLKhAFYj2zh4xSeMoQAIgyPWJIAgsjvDVeS7aOqxKfZTZdvGvnKoy8yG5aCuQ1
8/Kiv2FvrRZYBg1mDCW1lsWSUzwVBb8PbHZlUjy3utGLWKqXa51s/7Z0l8Ng5ezFCYBKao3oOCWe
H8GzCj/363MLe8O/AClmSxQE0JyYQGAWKT1csyZUSmLgMiNg0c94lkip86A2Ds8UpfKAyn0Ixilz
o/pTD9MZB1quS1pN74EvihhgUEfygnvzkNXZ3H9naTqghG7tdJgzPotPooF7rEFJF+rBNH8xVKEl
GXOTzxJDeM1OUjsMR/wykPbl5sml9oVXyth4naxdnOR0U6kDnaEomJWMPyGWiOgOiOZrBJDRJ+yG
ZTHPq5K3bzcJLr6E/8wM0GnwAvl6b7wTuPbX86JE11a7jypQ1Q1jDoQmmc4XMl0BlMFnc4wFPMj7
drnJfaQyvo0M3siB0R9SvdSDCQxj1OazYmD8mHla4/3WnZGM1I4I3FJKcpibErnNd2Sfd553Isrm
UHHAyP8LRrWe1uD5ysE6ITq0QBVUYb3dZPjK6L7Dx1fjrG275Z5j9vvF+xvZhsLv46fcRaYOdIaB
IH2nwOy71qbvPqHX3M+KS/oN25n/rvwlAOB4pMAIbNjOuL5Fr7ELpNiCxgI8ktn53TCZRlgdjcJN
AhwLjD51TEPaztqQUlqe+aQCb9oPpu6DNZZ20QBm7wAz/SOnuKMkcij/zMuvmdykKNt3YyNFVPXO
lDcitaYKQKKTRBs4etu5H3jyVIJhwIEMVH4BiLxkX94MfKsH95QWB/2igLuqB3un7KPqvMws4WSw
ANcchXQCSJiBJEC0yLxXKAitKHHm/LJ5f62n5tORHIUBfIPF72p2v7jKraG+cJKl/grce81CRkBI
ZUEMszhgEGQS9rqzoVZCAGA2/HkpXk9sS4KnI8t5eyg48r8YQlo5gyy2zzpswYd9CyXdmWLPGbEV
3PWwSdf1EiZSoUxSrMu1b//LBUApPDafH2BLVX8/EH4nNogy0AfLUHeHvqknSLs5Zpr0Ngkq0Qd+
Zs628/KG8DJ0r39ZwEaESstR0V0dgYO0GyBGjYLrH6BRFYqq+89L+yk86iSs/qGeU0xcQsRC8/jG
OUi+Kx3oQdJaKvqvpM1phzFN9/OFxvHSWeE4DHAoEbLsCVROFbwkMvUNPoy+X8hBcDTvKL8/Qr56
xpQS1kN2CAiKk4BKM8OiofRow0GXr0jmA/k2v4Q5ZHC5q3dxxH5U1/1ltn+/ZVpd6lxEMJjm+it4
ijPSH1K53SCtSs1d/VWhGR7gVKPwbjlpr1TVeKehcdsup9mprMFNCdUmCCZT92ROxc/+Q9iIiXvz
U0XAGaptLmsYtTYa7hlLLFi3K1yPrFtUNjus09PwAAI3d2cU8YZ8VHCoq38ycNDjkmRVbE/BgcSq
aV9MYMUoAPeD/ZrA1DIDlcRR+/VDUQ721DiNzQOaoA89CdfvaoSwbcjCr6au9H8Mer+oZ/Jskcdr
Qq/LGIji2vL4YuEfqRM/skFGONpOXkkMXpgGxMbl/gOIvRo0aTXy5s0UHuD4SrHy7311lweFAqA3
v2TEU37KNyaKO5PMu+jGfQWtVdtxRY4DH0fa0IAFEd+4AqTLuqsRfBAb+PJ1m52FSvlAI5GVt5gE
y5S16zTwlC7xTJ60l9mf4hb3EpzIIjp2bl3VepWPyiIOj0Izl4q+TqYIhdNOCsUzEcEef1YZK7oE
jHX1dpEdHOVVNpvjN9PCihIFSk1wsP+mGS6UdAJf9odV0diVMD19fbvgjux22bDqLonNe4lSJKCo
/ic83VocesBNpQ5oq9z120yyhPaLJ9C1WGg12It+hESB+oMU8qFd9hszaYesNlvEuiNcq5Z71qSL
33mdPGnqIlaeMjPJKqp13cHRpx8B4e37ZOdByKKAhNjSZ+RsrDu3UghCp+RhqIri/Xe691MqjW2e
ccMvSDWP8B32ONUs4zTnhg+Idp/PG0K9o6/RW8SQJt8j1jChFdGolYb5Yp1ByggKkWYjkDz9E9zu
KJsx8TrbtFUGFV5ZeabXheOkhPgy6ADdJhL96hhIKnJfx3aFjYPpE/fbc3pj4956Lu2BeEdlhTcf
IM9FbCiVEzyyuATAulw1SMA7kBe7dKSfJrw/x4BJQCBOGeO4oE+k/Vy+T4WYnZsCST2lDpi8w/Pq
TnDY94o0GEp/5SuF8k17ZDmONEk+QgSTWi33Cng4DZOsuKF5X5m665FbQ/hCoyrC4gaIHYzKy7aW
GOtDMvgpuC7SGanpP898tcMfo5hcGx6y3/XyHKcg4f3k1mdULsdGUG5QyyrN/AqTZRPMOz92Mbt3
SvuFrjG12lRc96smLyVE9g/w08cs8iBz4bV8U4WJZUjNEIFa2HLMwIXW+RhF8lJj/RfZiW4nCJCF
fPC24MLPD+8Ru1OGTi0KNKcHb4yciPIHYQpxOReplfKgOjJtkAQOvLUz/DzHiPoQZOXuzhLpzx+p
w1RHGZzD7r0RJigIg5TgGEWOTraHD9xU5dTgmibz5KQgs0t4SdZW8WyM9mhuuPxg2/hJD5aPqo0I
PzRCuSFVkrJaTvCnc8vpKe5ygk/MwwZGOwQ9KSYOvKvZXNeyTEWsdW/iGYPqM2Z2abq924xFO5Iq
7+euJyfF+PGtCi+7JBhKVBxOumRD8UDci/MCRgTH9r+DadcglgaWu9LrYZSmycDnZcvDnySycN38
9r+/0pQkgKfQxpXyXpcrenlTGkwttENJHBZ60YY/2PExhXjQW98yhS7xyzPLIKL6SGL/PNrTY1tz
Trt7GDnrHiKDjjOLL0+NMgE0YME5gDFEf3185nA0rksDtaK8N4mCgfLH8Wmq9nsfaMaVtIjbjHsp
zC+QJ/UHmq/wpo9B+TfdH4aaP2Ya8E+mGN4hUMomHVWLyc9GWnjYILmQaEYLYy4dQNbYWiMrQN64
nGz7ooE4jwiD7N2ymgy6Jvd+B1O/FS4+L7aohPNY2COE2pn0COtjM2cR1iw+JnHWjZpp/3qDihs4
T6OUGdD2tPwPYJ7KuNAKepfcBxfSqkBj2N3HJidE4KxxqhpxMRtGIkOls7iDYchVkDZEE8daOod2
pwA+UpCMt8xvZT+e731ZRGTqtWN3B25zxyTsuSqjlcFxeozLkmZDarNKBxany63JEXrqe5hvi5lT
5LQjx/+HHXndl7FYxsXKFdPelab5DRelJlUKvEBUStlRIGi66KRz4PojqhIAAEOEnXfaATSD9+sc
+CYrIzVDK8t24il7WQan0cqNzzI3mVarchbUBYihqb2k9YFc0fsrXIZb57axiw6BDX6c0TFE3xut
/unJy/qmdRshA93hwH5cbgUYKEGd7Viki9D2b9PB57KoOKjzz3LvykiieLMnnoqPnLSDAOLwWOhD
C0dWi4xvR6B0SFVfGJ7DzbXDET9/Pq090XvrTjKGigHqXBLf7Nsf+geEPx95t/b4atob23qsK9TA
SZxNhN+0FjWDLVXEJyE8RDTvDq9sMn1MfPYJhKy8bFhW54syiHPCEMH2bXxqbL/z0fndY6rCogmy
68CCN7B8Wxf1wb6di0nWsJ8EEg15G5jzN+NLOh+0rBHx3sNIU7LVCH6YHoUn2Wr6zvltpceRP8Js
ATJPj54Q/Kdp+8hrlOhNAbaz5snbKeeDYDVuDaWfMkZ8dNkb1e3/+MjiK0/T8y7gGtfoqtI1/3pO
xM84u7VsdSHeAMkHnfBOoNqB5nFClEFiwdFuCbj1CwWiofzVDF0iHdve41FcJvf3X4L+EwHzBzdT
D1QBV5WgJr44xuEwOsblsZstQG5mNht4SRPE8rfIcbGvd52J/BMC7CQPbasBxnrsxsdibD2A9dAn
KTjekbR5HmoxfdmDd/o/FFX7uXfzpT64Y/scOlEyr5OYMg1gRWkhdqFIE3hl+ozqPmdud43L/B5f
JCHXJsukQetuqe80zzZj66EQZMsB/7uk+/FghxvG1LuJxr6BD/FptDy2jMKU5dwuDrmujI5uJlxL
1eDEGBQG4IFK4FIj3xeFExYBaU25U2IBZq6O2Xzqi/ujOkvn2S+6cPm+tg/X2IA2IFBUE9pALEnB
6MSBmaiV0NF1gd+lteztszhtw/hXoYCk5jBKuZsfEXNm86fJODTKlKWta4tDoy0zl646JosQgwdH
yA+CCuLC7IiBnenUXP5Gf/oKVgE0RF8pfq0VD2pQxBxhlXZjAwo7Tevfn+j8bZQDlNzFykuFCjiM
oaWLpX2tQ+1SAu+WmLXP0h2gNszgA/UwsIq1OosoCmRiqnIsYebqwwqekxn/hjn5D28HgnXp44NL
0Wl4AE8IfGvOVA/MvW3caNvl5Pz4C/A6SbBwe8+MZgRhV5u5p+ryeeAWnpIBSN7dmpircitA5jIR
n83xikb2fKgXd0h4+nqx9nj+ZAe9dlWka3pW8vq5NWe8cRmNYHG9Aas4Gh2fZ/omZh7Xb76ssn84
CIu6fU8qQIcoi+q4ac66hluH7kq0uexuUC5wOZshsGhU7h4O+O0fiHyUeRVdzx3DXVTBL/20w51u
p2TFNZC/OpL/5fAhCQ17hq6KHCajQUzK0I7CRFqttbHq6ESoO/Y+DQQU67kCERWYzE3q2InaXRDN
S6yFCMA6S6W7C6fOE1gzS7HtDWorjDLb1fadkrWunMHEglh3NTvm+K4QWay/PENCM5FcgA02az9h
SvuWiGevCV8PnHIAgKAGlJ4dS6TIbSqNkgfS+bi7U1BdHbzsnF0w5WPjb06CUXGDgE3nxyowy4ic
oyxgOs7ag5+yblM3ezeFXDxebEHM/GDnf7y5orepSsh0+ySHc8MmJUkjLqxhlxSo2V4BKpwS43Yv
CiP5KoLIQ5TlLz4Ubwed58+UbJqYs9l4zVRQYvVgsEJ4fmEaihGw/a7OjNqnE66Vk8QgfyANDHPy
tEGkt4WNhspIN/v7O1V0LEq0wxG3lCb0Pq1Ot3qxjiHXCSnhZbrcJRzYH7X9IssSG10J9X+rEvYs
HtTagyxsr91yMjK4+TYSgcKWEhQbO4j0/Moagz7QYSqsazXusYRUxg9TGu7Luuj6xd5ItK/XzIMJ
hVhIvJ1Oq0ept3+ncYKy2Sp5fKuwbX5FQ1SOm0dvSnRD6ZQ3KJR2VrA8PiYflYH349IacA7G9G/o
ZVLcfuuKSsBO4b0VWlDMHhiv5wyCODvMt/6jXUTVzR08LuRX9uv6kmsODCo4pGPLeed4GzdfoJUy
jty+KTzN+EnNrFvXYKVVMAn1i+z2wbbBerJl+1G6AQUgtuE/En7MZ3cq2ZQ4WiBRzj7cNACSJhq5
nv8X9oKQonRvAHaC2Zdo5KEaNXyVSawA1q8w9to1NNwNjAKaRz/ji0AeSyJoxBQkarmHosQK7poc
IoMyh6y5lI7nIsoYjsKUzypuxdmQfgHQOR9mT12wKVo2++LzAzxxGpL19m6FljZEJLqT6pGXifqs
Xq6NVgWk9ldQ3HGABfSgw8V+ECsSoFBMUnz8M6Lnq+j1rVyhsRjlqgGd4w1jPf+OFRpvPVpK45XS
CxEKEzfuPLzvp2V0c2JQuyGceY9yqHefrPn91Hm2TJnIieMKQww7r0jwPtto5xzu2X76fWYOKQwD
Zt0kQgkIctzrx+02OyIM+cShZ/F4sPZ0lkgqnU1SxZFrQJH/b3H5rzpmjFAMSJjIZnlpBh/iPIEe
Je3KoXdZE80Ro56vw6Yxszw3VwKapyyYeMvQSm0A6ZBz5PIkpjV9KmwI9ASvyR0ipEvfoeQkWjQT
gdRe0N5ayeWqS9WrDC3bJ7GLDXhSopY07BxRyAp3B3pw2vhgYMFDuOwd3mKzomCgY4bWZHl359iE
KHGF/GkM9nAsUOoeUAxfpcOh3IGVsGi/2as2Th4JQPjk1faH9eLObVsS47IhYUIPwD/N5xs+IT8Y
DDyr2aCCRooQohLJqnujMXchwhIv8BoVeiLs/hpFD5hclDxMP+BXVUZ6gh3ZjtQgQJAaUnMg7s6M
yhJxnVLsNMayqKHWHBwFZ1l7q7tzFA+bB6jDFdEv/sRu/w7od0lsXkTZAX5OsRA6htcUbM8WJD+D
loqtPjnlWHm4jUhRk9jKkX+XAVLnxU9j/IhZvRK7RwNeqMdfj7c+QCZSIW0dG3dug0a5OxeDnyTw
P9IVxJyxbqyBsg0WiK1UqHIqAZNX5hJ/lwfBZFplLxf1Tn+56PI/Cvz86hc4HuULvvBdhij5Dre1
/4YgrOy1EegdK/I8svyAY3WrvClxeZrVX/eiG1MaXbVlmmyHQtzAePgZsgX95lsKKxaQyHDX/HBk
M8DqYkKSx+4N5a8fc01alx3JDNUYD5CGYvWY9UDU+ZTHxRhMgDZQDSpeAPAwQ+SNqfQCk9uNnZVR
GVfdxhWXFbbzVzU/JYVv7y1Iu/veBTUCv8+WdS6knJ7ami6GXBeiBWllve3DWql3V1qKUyxlP7o+
lFARGdXnsN3Ky459xXFr7srxWV5zDxrWRnP4TtbXruEtBwaYieVixA253zJfbukuNZ3xckKVdnU7
+7NHYd9oKw8Z5Njv3fuxRA81GjAMJAPu3dqtRzpWpt31tbfDlWTuACHsQt/FCOZT3/hpnJKkt9aq
YHIzi68Aot9rAsWi/3AKIq+biCoImLn9aoJHEYPX8Rg5eF92qRKaNONL4Ijx2RJKMGQBln8uhqQz
Wj2KUanHj2yZk0OrqZeop7bEEhbEwVT2EdU4pcZ5T3JN8yWDOfraA0k0QHKiBHQPZxtGyTPlDTXy
pu0dLgLYAbzTGQZhzaj1Dio0RXAS00oSEgu9tlu4eL02Co55iV7jWl03V9msz4JtD15qKELi4pfF
eqmmCN5U7j7Zp7o0g9xXtVgjJoaLyusqTqDLjq1VpDr/abtpyPI+bgjzH0TVmQoo/IUYsIyZf/Rr
F4JUQGxWUQCIFAa2iTBreiu+DMjIxFtgX66SWhnDjZF7okfTekmBNZNTW0aJGi6Rz1I8Ndoxb2pf
taLATSurKSHyVJzCz+Zv9816TOAF1IkdNNU+5N//WhIXgh+JcRBRTrP6UC4tYgSdUA8FV5MRE7ji
r86i0rRgeHdA6B1htffJEhbYaFOwRPTPSN7mts/QoOp8ZLI1uJeL7OG1/nIcOlQ4gRC4EevSyf75
6MN8zeVk4JJVw/QJch/03qAiv2oaxAHhB1VTeDve8Y1dirrjFX5VL0OiaxDhwtkeLlZv0RnVK+6k
EtnCCpTRqbmTa0w4fSt3rA7/PlvOV6B2bfriavD8D2McBzN+BdJFWghOXsW3ARAAs6gWv5O9NKBi
qSxIRxH2koQIE61FDEWa6bMf6yRYeaB92vezbJlNI+hAlJSoI76bTtIsQHRQ7rJEJbriilZqz/Yv
Uz+/EKXWGDMH4EgDcbqCAd9HVvOFSL3PS1PuIcAgTNBNDllIel1bUrMIZQoS/qELdLcGj9P6pCz0
JH/r2I4AMNZC+g2qHfTnwQSj0AUU/7FeecA09f/hRwXBsSBjAmBS0nOImq/MkkkovAM7mTT3FsKw
IE8DjyFe3VwEgrsbBLDOWg78l4KwyoPxCcpekE//gsLI/5Tyd7VCDKhPvtyiMtVRODpy8kXMX6h5
Pf0PuGZ3qPbAUz5SYO2vD+UxlAaptvpOguqEUjNP643g8y41I0w7Bk3u3uj1Du2rcqExAy3mCmZi
co9tvbxDE6e2jG6Cky0M2Npbhcsg5Elct1jQp7bjYPkerdNeTfLBln7ORwHO0Gs7Asg6fuxvbj3R
LMQmVcZNYWvucE78kwMqWtsEMj4UftTMuz5AViQXCL5ACdP9MAEGs7GxP73wobeXdHXwd6cojQeo
K2Lb9FyQs0WN2uK/z1LTlA4M2sfWUlUwxU8svDJTUtJ49pcOOY8BzBYaHzjFYVvD7aMx5rogzLID
aPFi4ihZIVYFDRQ9E2gEx9jcDvGFOGvtuBJF+P68x+UBEVJgccDmb2nt7VlPGTYaoGBsqmszN854
0uXqq6/Dv5tb+USEdkwQwYIpgityE9kgm5E2UmBrQEFyg2iq5qLOCd9DYmSuJ17Dp+B7aPKIk+LE
rPKIeexYC/mL78dWJ1Q6QwJp0Hr1LD1inW0NZHm0OvEwhJJN956JB5oKdUnRZ6onZN1HEpFYwc6G
PtdnYDYCCfxygg9w95WQSmNKab3TFciz7+rr0rfTUrecMq4Nl53knDehzxzkvaCNjsaGA1/8nWLk
2UV/mQ+S2StRwSXji92fLg8xcFMY+4ghyGfDVIhS9lZpT8F7Cgs654Tn1ldHKcjgKmkvsWxB9Dv/
3jlqz72czBkfc6OEErTJGjQmejIYPCZnnAtykQMb60FGdCKppHMTE+MNANl1dEzA2qkJv/jEZkYE
nNCaj3t6DpeFxSSbRNwZRlNalur9K8HwlxKaQrzsRF2pOnakRSi+czqxVirOdlHO4jk0k7WbK634
GXMFJFPr/O1MtoUCcqviNRBi8eRUpEAXPg0BbdJV+oMXeTI+waP8FsatRlcVxPZFgXDIiP5mBoZY
W70uzOypAjq+DaXWY6DZg1EFfmoe6HX2NDoaoUa3rGMI+HR/LooTcHgtSNNg9Mu8dKoqkFKiybcX
WgyuphxCrK5hcryuMmsdgfir6lSPS2mZaFu1bPPKghYw3hXsALO5TnKWZls9Rvh6Knu7FsgMT4qM
fPHTDXi5MnKSzprBHsIcQg0ESfM90EQhkhKXgICDZwogtAn2PDe2WQA/CgxzusIve6nQiHOBii4W
08ehtvmQXSh0gW1u9Ql36VD9OgojyD/rwLjVu0ZnXqyulewsZK1qPDKRr68VUmLUednU2m98kmyx
3G3J93BEH62ecFgkJ0TxC4BN9G7LKITK5P4f9oOQXZeFREsQLSoTgzgGzF/oCWjR5qp0tw80uybq
qdpKK9eSpLaQCyWe8FH45Aq7s8zE2/vusu7MHFflXNcziWnzFjdV5xaucVNa0KmpbLbC103Svhay
7PblkwVTRbJCJ6CZ3zsQLr09Pd3H7p8PhBYbcjsT5hWn69NdKQfos1TZngdkiSXuGu/GSnWTY6zD
UxnD3LxaHaSLB9XkZKMzs6nG81plUaviagIXr00W2llbidYmPewzQJ0bHTwyJ6vwxBrlLKSSsniu
IAzK83kZP3BDBG+x8nd++GF2egiYGyOjYt85OJdANLWHfxjWlVkkp5adEFV4J3/c54m0v0uKDLC6
/eP3r+BAFePP5up/JuNpISAMp5WRMW/v/6lCCEcbiZIa9KYSKGA1SM6q42mel82tfZo2anBBwy5a
sut5JIZE4AlPIfKKXYbJobdP6yZO2qUUiv57jHuWgrLsTT/6oQBcHnambh+Gjb9UbTrjr8oLPkGF
SyE9OjuTTmY9+NAfVdt4MNErkhKuPqEukTEQ0+Om6ZW5gzpWUoonfdQsCuyGShAREf31UpgSYwA3
lkSUSwq1GAg7H3cYtMHhQNDJeEF0zdyfL+C7HuJxFsPipLs9Zq291gavhJkUu6D8Fty6iFdF9PNk
kqFEBk1LgFIgeQr9uUJ4Wb72i71XTsFbUSRdX2ilet2NS9WEeybv/dvApApbKG2GUYBSwdyRYcwK
cnezLlPXwVg6id8giedVRPEnSVbBxrmVguNLG1GKUtdVSNM1sgxMZgHv19tJ7qi07B4M0ODPII+j
XFukcbxJnjJ79XC1AzZmF8SyKTgVeilhIpRh9cnhO4mIQux6ESXgCqKLdzTqvUa0kDEG0qdXM3eh
M60VjQ2jCzFLZsQ4wXsBfmn2ppKEa9VWJjCV2oWB2gTymidIbmdmRNdOhP8X7tFlQWRHsw+FN3RM
JnaCS/YZaYsgDugq6UmTxRP/PmKCCTKRtEdJ1HMcAie6It8nUR3ShjdTFcj1bRch3Sw0roFvWEGJ
n9mXvvih7O4iXYNGY+U6J/6Nf7dQypKqJe9o0ebm/TnEnAu0+pIfRqxi18e/PASSQKsCuvhT9l0+
9/xhmpBtlysXgqodt3fiHJD/brvCk+WCWthq/V6ZksiqbeH4uTIGOvBmLWv9zBfdonTKlq/IeHtu
xKq2cMNBhy+6rs+wyynBAo75V3mPljN1tEc+vpLtx7miWEjxFlFTZ1Qn0l8n6QYZF78m0ncQQS2+
4ZFJ/CEQu9f0ZaRk13XSKIrtxTkjb2N+X97RNssVDrfXxKY8lnYiw1z+L/cOyTGePQckepC6Q9Ba
5d7pbPb1g06qzs84cVQFCOgWQyTI6ozyzRY8y8pqjW8MPGzvCAhq1r2UUEjBsGfxgL8CtZJaiJ4k
pQ5kRYOL41okT6uS12a634Bt7OgzhH9kV1HqwSGTXpItjq7btRqSSbBGzlmEBi1wc+rOsCkh3lM8
BhIlJBgfQDqK6IOmwgfSyw5QxvHeqsek1X8VxwVZOPxUj7/7t/TdghR66N2mLvBAlcQgA97H4JWS
Ss85Adci9GTei5eKkbWVAVbDEzVJ280FyP0L5vFLxxCYjkVV4PuXzpLxRZNQgQLuWj9r+HV9yzyn
78XLh3gaOhLu8E9XvYllo2HVAP07xo3J6X9PCUSh/BCRtTvnkzXtYQkXfbx5KuzlScqXk+hIiZWo
Hk+KcmKnzdxYjSD3YUZwdPAWUOOTdmBsPgBQlXipfewW5cKuHwm6h765EcPexQxhzxGbSCtbPXMF
UkI9jSXMvMYgmduIKdebzQyyRcswNdsRArDfYFrdQbQBMffnx0TSRhBnJtyJ3hjrzyQruvB34qQj
Go/ZRYm9EGyB14AjO88VsH8a2QEYY2ynqk8YRKLM1JlkLMuNULL/fgbCIL0Ji0xQHQHSwAN/nmYt
4dy1Pn5Is6ZGkIvVbuWdSKubVWHsbI2/JB/T0+KjAAJoT6J8uvnCPeYweP6jvGDuFFEhpIKL5T/X
my8+dOIAM98XZVlt/iLAvFHyz2TsblvwnuWSJBvWtkSz89wLAgr6FsEyyCXL5zL655Y6n1qpEg1c
Bd3E+wlfqsrH4KsfOV20mloqK6U6VYjsGTPEpbOvogxb+E46/wCGZ9vOROhTiXHPBcRcWVds7TWO
8Dx9EYhlqR3KzIrp4u+Bpc/js7elobPvgEVDqB49vwi4remUPQp9lsinAJXbpc6yfwbZkiWNLAaf
Fk8zML+M9T10nRxEy75vdyDtIYCFkMn/2Yq4u6Bovw9ffbmuw7CrbBrXd7sVrgaIztVyLNjAe6Lv
Jn5Vg7z9gFuV4xHkKSlJnnoL8v0KqsmJhpboDDCLr2Nr+YA9UqxbBE40WH69DzhaJo9rm7krmeSp
ZZAE7V/itC6gXEn6pkXTBajIuYl6jrRjQjsdPKpWIWq8wgvlHJSaBdjM2a+A0IFnOjbKIltABJw7
yWm/SoWbMS4P56FEjyGWUjaiwPuW0HFdypMQ+fK9VOQsaJ789uGeclpXwkx4OrHiwMJfNRj6UIwy
iAt2e+/ABDy7Tiv8EbtjWl6ZJBfbDnmzmsK50OW365K4hNge2DaYu2f5Qw4KkJpyyzA813Bhl/VQ
VnUOnyFhpkHhqmyLW3HOL0MssgEnsEoX+zdubc8ulCBG2ZJ0dp+5e/jDO2ivGv4kdjY6PiP9H2EJ
vdclFcvoah8d2amYnPyx697w2jetv18+MMe7Htsd72RwLd4HH6jzXS3pi7ymXmOlx2zXIWnPotuh
XRfZjDRqONt7PwpzJjqSJyngB7D/ed016ATaePXCY3TtKfhWJXQuRPtR1Im1rkZuDlv+F83G5DlN
35XZSOn6UfEhubnIRm6Qz6R4jLjA+mGlWaOYFvNpocxoDy3Gw0l2OH8ziJSFyY7qchzMoXeQP5P5
iFz8Gk7ilKxVtp23tE89g8XnW/4RBSFBFsPW9sEHpBAX77/7JE3gp2Y8CAeRqBpOaWqR5hDunTZ+
21e7zCjUTzUl394mWh2eoM0R8Nw/C7TuimBhL0Ud0kSiDz+S4EYQnJQOwcRZJq9px6+LfcQlIpoT
vjQtIv6kjJhczjnN9BMF/5TtRFIZEWvqpVOm2T7nBdfnELmuZf/qmRSticVmNwwjRkX5IKDpRPsw
1ujtwuUBaRpOMi3W+awg7a76Fkj9RpvCrMkr+J4ItG8mlQdQV/tWb3Fd9tqQF2ADuePflmZIaBBV
h8ygnzA3KVjbWbQ9boJvNLF5okXLOKjWApXB0wK8cYm4+4i+kUk+Qq6QR9+uPvlXeL11G0DenZmp
ZC2mZ0NofG4LwyLZ7Dbxlis1F/A+blgeoN3N4bVtj+M0OZm5t5w28MD1ArBYiZ26yerAKgpQcRQN
9554wx7lvcvzSK5RJsxUX7rxPVT3ANgQ1LRNaJrwBlUUXvO2vi2L42lCu/XtzxsOwyQ+cBS8BaJm
1t05PCQbZLI7iL8Uw09+2SXtAohARdS2xcDYReJde0OfPjDuH1qdliRtCKU0E1PgPJgICBJD5T+n
dSBA10w7ZTKkpNq5E2ljqZ1jVl/b9z42qyN5nYgPFK2nYbE+uYduooniY+kvairmxVayMhj4JhHO
MQr77b6q7/KpO2zDPnpZfalSVKTajYuZNiCXJw42WbqateCGsVp5UNc/Lj70wjj89myDTlmE9Xjj
SdiheC7HyCyu7vCi62D/h73a2JfGkgVAPx0yFmIJkYc9N1eCTS1M1fMFKc4+WJhGmEvavIZJyckW
q5xv6mPikvo9dcnecuVfG+4LKFDF7EOtji1ULFE64pjrf7JssRQA/o92IAK9M9IhGHGmJlLDU0Ur
HrAVXJ62SPCUe1btIVCKUsWHO01EUAzB/KDkkZh1k+PV4uF7BHpQSoXxh/2IsOOU0yLZvH1Zunmr
m/aFHuMQcVmHQBwMqKdQ3XQc/V7/9YG6jGm/Uar2XLgEMEG9n1MGRDPj9vej42lnx+TR8chrkzm0
Gue2dvslJ/uu1kEARo8xSQ9OgfmuATN6TNRqCgShAPQ5iiE+255RwzWMLfyIqPr3iQ7aus5ctaDG
kA1XkRPljlIpAyyz8vRPHvuEQhlywysJ/W2CkozIZt3OkHPzlPC591EL/lp0U8o0yKulIOUhF4hQ
zwyE8+paziONgr88Ga0Hww02w15dpP/V5QvIGQLcDqtOuWNndXn2/XcK/JayFYUmPhzuz0TyqPt2
gBwA6l+x2KYu6LuejGb+k24ssXliC+/Y2DVLAsF7HqmSLktSAcd6vytsD9ylxvhp0ycc/FYXsP5C
TuD3sKNXz5Cppxv6exO1iG832wAjwBg+ubFdhadlRMvnqBCsJaYTK06u23ThurCuvpUWpBTxth2V
LpSORHimU4g+WZBbacIIdXGwAK7vr7dvC+/2xioqFYoVg6KdhBvfuq/KD2VCXPd11UcHRNrNyf1+
rPWLPyPhkeFuZgTUNli/Rga3npUQcz5HgIWK95/KCtk15pNlSCV2Gcd0AcdkafTD05g9vTXtk1pI
VCOp/rfZsSxpqAy4YU0a8KnMp+Vpi29mfyP5I3dZWtn4IXp1UICwfiUkaG2XJScOGvbzguhpmJPZ
obdyMTHdD/X9OMPhNogjba4e4QwdvIvIiKgKLlhRUueQUSFhTnKMtfcPr8UWVV+FGJykz2qjowgW
K+SBORJt+siRXYuKkGpcc3G1kxc0jnwavMPdis8yf7CDq0no+tos+N9DpScMVFfwFwwJhWDWWfKb
Gkt1rnrbb2a12Ud+sLgOE6Bo7Ap6lOG4czNB1of0jidn7wfoTw9KObu5hMYQp+/OmZ6upN70Ua2H
H2l+heEBLBF9SngMyNSM3iMnuOCeK3l35KBEFKAXmfyO1yc+7t1tjTBvlXyQfPICCFMyB04n02mV
tPMPohFDY1yrtkT2lnqRUuUcUK30BiLhxH9+B2XBjYkuyPs0oNL0KP6wDImdr5OuQ4rqhYGmV+kD
SjYTQpHKuBKF3ttsiSMpDh5wvOJeGgOqs844X7gJV/04m8/s7xoNEpqBsEb0xAS14F85UCdBNfyx
jPoZ5iu8lsnrDZNX+rYb/dMVrVyhEjP8GR3DeS39jrkXhy0LutjSzht6Z8ViQ9AKjf8XITcv9ve2
lFpWjA3ty2L6CqT025npoqUvyUC6xf/AljZ9A59We6gf7/irVO2d6LK9ieWYr6taiUnuXL8CyLO2
/+dA92nLoRiTisU289uCZwwFnNTbF+ycmmh8qVOEz5ZeXSJtdkDIFPw8lrZoRe4RNhRy/KjsPsRJ
qSqtJCCisCBVqxTRVHWlY59BINNJms3nI3i/1UNlWl5RUZD2Ta5EPYEcdLDc0FtTvwSTCQEGRnLV
PBPFF1BbHTN79lN+drIRJmgzLkhHhZqwSpNA/YgSHP5m5Dl8sfAP9VUiZhS+AhtPmsOrtLZ9X+2Y
fBN4zdXjZ1XWP+jRyjdYr8UTQRRwcUSpfB8tVAFh/dQnSO0inmR22Jwdh+PyzPBzT27N/3H8D1SW
1MUvj/QAossh6V3tp5R6xQRAhrZtV1OBR1VvP77F1AIQ0HSv6BiFYjaxfdXZ0njeb8LrmTKRn5fX
QIunCAwemv4WJm4vt3tml9YTpw03/PD+9RxhvyJDDj0a/zrpTdSfkbuLz4aotXBNN8NazcbJB0fn
fOPJ7hyuVWaXiheQdSxwx1MeRoenxH55wOKVzPLjtBlQ6CC08dwSuoWAU+9k4esW9+1I6qn8zVh/
lEvwDGHsjDpm0AqYNzRF9p2YDW//hcrCDuzcr+5DqspRTek8BJKejc5z62WeXVpjW/UANbGvgDM0
bhfeOiCfuR2FRqHNuXahh1pPAsxhsl99QiaIuoOFqvG3bmTwg8E4wHN+SiT8tKAQmRJutG9QcIZC
HNYnsplXcmpXLLhkgefM7x4bF8Vd49jgO1sASd7NlBon/+Gk/D0kqhUXEDWoaZi0vqA6yR/+8cds
kXrOrTY4PFnEBSdqmMluCP3KyHRKSqWRjGDLVNBpkKCNZDGhDu4cLd6h+HIliVe3fBkdKa0r2zYf
4IcJqAmryOUCuApSjycLPL3ldfgnh5DdGJINtpoSMX13zpkwLZGezgSmx6bn4ms/fOfupGAnaIrP
l7/cL2SuCgzD2dF4J//2UluG93/QFDd4hVeBG137kr7SkIapNFGihNLfIcOZWjUJwP93gz9sQQhV
6Y4BaXZqE6cZ3BOf2hUcgEKFbZWQmNeLDO5AtZQdcrUSirW4jsmcvr98eNgPmDN73brorRWzEMwU
EKZCxJk0tiqmZ1dg/bftV+JXvscC+84YWNijArKkWDde1FTMKcnH62C0pQ9YPYoy4haVGkzOG7wz
n9/aDFOWJUt/BSqTDdtKYVboyok1mj69TsIPs4G2aTkwbmoseEKAIggJGb8dydPDBDWW3h/41zy8
I+4uelpHzl81WZHP49W4ZvanJ5a7YyVqWlyP7t/kSY/6od+FVTnvZ/uFeGSx2ldiiQPAsS/FI/oz
iLsRpiPZHHkJHsjwrQYvvPn4/padizHJeXZrYaXHZYiFFD4zjD5O7e+dJO0v9V71G2SmD1QyHyHe
k/Y4P95fIAT2OkJd6c6gHSVYhWRgr2vvsJWWiRypLEgkK3xN+AILUHCMRZFYv+cMmlTsNFvo/OJB
25hgtZ27mIzhid89baIK3LXvQGzuHi0fEC6yo4xzEDVq1HqGv6H9MqnjVUwFQSSgMk1zZ+YUt+Sf
vDTeg1s8vK4jkARz3HxrLeUSgsgjV75TP4TsN+UfLo+6JYaojgRaC5pgqK28fHkZEq5VYKVeSqkM
yZEX8E1cj0QShdD0XWNb3HmbaI1+NOENzs0tJs0Vo5SFzujnEA9GJMVcqscSr5v/dRslJ9jthSqy
5kF8t08JYedqdM05FfurF0XDVoWZ4OrYtw/xudCMEBWLzuByoXCF4n7PR3GkcydwSfSVaEeE2AEF
PvghMCW3DCa7IHiaJmFFUz5h7H8I1UrJcfvpU2OF2HxNSYxEMA76V6rPgVf7S4uKDLBI4CiKC33k
6FaO91WnjOmA3d97lkqkIZYITXX6K/L42BKU/gf3lt20aJc27Zgaf3WbVX1UFB5p3NGBnWf5QsVH
Dq9Kt+qsUoHEiLEr8jaA3lEAGodLNqN8C18EXtXvQxSQym0CyLBkJJ4eDePZJSaf78WoaLvloVkq
1+hTVczH+3HBp0bBhbFyhjf2+s1ItnJ1N4bUvbCrRi1EIiEKs6fz5I/sNqTI99MxJ2orsTPz5LO8
N/XLAkSIyu/vIsbLwOXHrJz4iMtfOWDIAUgHTkiDhMPtkdwRv6K7BMLR+lNoKSo8xg/SxSOaaJwq
GglxuFF8e0HxBp1I7dYZGVsQzhXKo9Z/C/HizYtvFq/vwCenIHhDJ+pctTlk07qGY7h08DZy4tOx
s5fFt31bf8H6CCGOwddoh1ZpYkWkHRYEEKylAoQO8gbpglEdCWv+/FamASTfeMFG1SiEq3EXNwnL
7m5mxMp3ssfuMlT1f1urbD9RFQ6Amng+8E61do1uNmFbNpBqEdmiA6z/K0c4QdkwDRGlhykTfIVm
Y06hSoIeAuYaUjZ1CVjjXkC7UMQLBBoI1u2rXZmtBtCMRS11M+lsX32XtIPTLzEa0sk43AsY69iM
ASmhL9II0KfBA4OPRVtS3chwOqKk1pyJchesABNeGQ7hQyRa/5xhuV4W/3lAWfCjzM2popznAl4j
JTsSUa1rsvL1ewnuICFkfpHSkK7SqRs3Y5qM8cZEWkzczpYxpIeDys7bpxIFFeLD2Cv7lLUE9lFt
G/ddXzaGo2I3Rho3xjkdo5bYqBSwisYfl8z81Kp8gwJVFWLZvWYiWrNub8n0sQcRNxn8prf8hYhq
J+Ebe4WivIQ3ToW+JvL0wLLe/K/gVJ8ZL1c1NRS1RGUrVmxzvj51XLv5gc3/x940Y9p9+CKJ9snd
exyeTycPl1V+IxdAAe+hk3nsFprK2uI1zyHwrBipxzEOtOVOTGCv4COLgQ1bAw73dp84rZLyw796
B+SSb+nlgR1ItpizXGUZhSFHEv1yaOnKDl6/wuDEJsleohXAQw+NqpQ4c0E5Ek3pt4pFb82M/ehg
XnJipHNR3NSB29lBwABvlcrYERa7SY9OiQZzPMFfb4MhZ+U0LUf2gATj+oTXURC3SdRIfVq/3+9n
+d/vfT+fWuZsyUQTnOA+fascy37oc4PDxogC+3YOtYBhLzB++QepZvzwR6ILO2hh1ZePJgJ+gjUS
EMP5hkYzrtzYV3Ki4XAywgm7FaoxyP37nfUlNmywdtNTCWiUW5yIq7UmSPFWGEVwZYV1ESOi1TLe
l7MZ+8WB54uifAjjN5DokotQJcQI2BWFqslT5jNkML4qsrKMDDuxK+1qW35ar+O7r7oBF+IBOG06
ecxvqbphDwsnvf0QzlGpe6huV2op3IiyRxsNSch4pvTchOd7FWwVFTANcuFko5/GaddlTMYPdDTT
nGtFNodEfS8HviwEKQ1c4KZJTa2JX3kT+f7x0azzfhqoG8N8FPOzeMsEJWAoR8zs0+5mGEJ8N/tQ
T4fakL4TKKuT9trEwoVh1rFsr2I3tNL6hchKLtTyEN0JhEmg0w7lGO8FoOie27TGKXNMRdELztHa
T1F9lXxCFo9b4F2ocU07Q0BcphogWBfghd+TnQLHkBTdEZaDIHoQCoVinKyh8GZNtooErS+V4EW+
vnrKBbOPdCjbyLdMAu3h/zHcbQ7UfqFBZBCSXWtwRsW3F9BufNfy7ErVqZodetBniLLUu3+LWjbt
fgp6C4XKyPjCACX49/uYnHBPmTS3Lji7k2DZCJXYamA4KxR5fhMpRCA57DnScKkp9aP6+dp9WmX9
tyvpBE8gHRu4tmsKTQw1yYomagl8H7GWspTIyZaheL510690SAU2TDUW/ju4gXKCUdBzdyajkhdN
t0+6NypYQiy11AuFJjrqlL8oUexj1pQuLSoLxYioE813X40bvqccIMTbqvYGDWun/K9yFcp50eVa
5f+MKWe0UfMBa32KFGSu+SIki7RTx1fZttGZ08fRa1YOXLRp+VmCEWfZZiI9AdVKqasJQYVDbIpN
Qv7xtM59ue+NzdEvW5QZRXYiy2aCQEpfh2uZFnZ+dNvxebUmhACOLGur9LFX1/ICLfozLDuvyUiQ
RIC52B5G6cc+5nE141iyqvPQ3sBIljrHekKIBbEJNFMzIdd6RvrKl++2QmqtqEIE3xUKgAt5M4Gi
Id7Uq43sE1eVtfBx16axS1b19gxV6qPxUH+FSuz+Wp62CauDp4ghprxYHohVkgBCA7GjxTpgAW0g
UjC6Nyg1lmDhuAf6fd/r7E7H7B+ZLn/8oHzRpsER9JfMV1ES9CDgKUXI4inH/d6oh9YWyKWXK0Nv
LjYMvpVuL3wYfd7nkWxZJzxyVeiFzUL6p6gHrkwPBjOOIBESCnWiXABKCxXtxI4WBndXQhqB/NMg
4EM1WOi9eBjy/jGtCSZU+0hMBy2z7ihCMV/yspwE14I7Cqf+h2qcrrHmvyCPaHPdYQAXl3Gmd4IP
2kXYeGdoMPBcZauad1z+EQsmDWxaK/yloa8Vt8hdOR+IQxMA0G8lhDUBo9QvIJ8z725WAQZ8btvQ
YvarQJyK8UGrLFx5pnVL5QybAZ75o4XJRh29/Cp9KKW4UCgKrGyEKauGXrlpCVnG+opi3aMluShd
c8Yk35m55Y1qDSO3+7QZakyLsWC9r4qzjK6bTDDs3ghQt0vTVhbcyiMNXUjmkKvMyrJsWWwVqD2d
yGJNuP2WDwVE8RnZYNY3IyjMv0roWtjl2Q3HYGTJkvzcu9qzc8aZUT5hErop9R733jMEFZkZVHeR
fi2IDqnIqFnF6pXD39Zwxy8nhIdMABRwmOPG1auTeDpvSooivrTHU7iIVAloGJtVOLbzeCCNkkyh
cQlCmM6pO0/52phELoxN7j8X6yxeBwoBUDrlg2SQTUG4hNGzqeocf8/A9EATMj4jNi7cn4672uUW
7hEIDLAZZIHvvvlt5OdP3q0eIQ8i3oEZA27Y94TDcLgwk773XuXmYssmlOu8qZXzxiGtDPiCXIi0
To75FQ2ke8g1RZ6q6+kTvbn8aAW4gcxM8xZkTiUQkmOeDSvR6nVJHebsGQtRqNXNuq4jfDmkMCGb
F22tkCog5gnw6Ltx2IBfB8eHFm84ixPA0v56wQdZHw6bzT3DSbXHym6crrLm7v3A5rF5z6NSM5cf
6zycwWhB0xtrVNyQ1na/8BXRYLnA5r+2ek0v8A5YY2jS5aoaXwA9RgP8SQut5iNAE7hqoJaGQPPb
nkwzquRvtIzld1zLqs6uGJJp3jpLBU7/ycc7BvrFQyyUR3xZ1VHJDezw4UvZ3W5GbU/Qm2ceue8i
Yy4pO47D30JMxGQpzhWh67cXPyQYxBeepsEBK5xoPS9w23OHLWNEhsL7Fepmz+Izbt3suESaPt8G
GUNRbySQIWvau+nJ6wNyoMdT14y4Vlj+q8//8CZXJQyO+cknEt2cAu8rjRB7w/PwpuMaglxKAE6/
vJiV0BHo8xp8ars+Xj8I5ix8qyB7Qg/8sBSJj+LfgFSgsnHieFDwgqiW0QghaYjpvquxAGlXfLHc
JHmNG+eZcunaRY79qSg1+NBIR8xgG1TC+p0FyFcR9XE3snOCILoCrSt2mqrZLoYzmQK6GSzVJN9n
zM2kfce73/EICsgVYFs+D3cUcqar8V8xJo6cgjjt5j5fGM8iK8TGfQbzwhoSOCnPh+VyKh78HrWa
hRExzRV2FfYivKnlUn8bkrIrNCuQTq8BXVez8caBygfUJJZPWfyjO1cMf5Ta9Hz4yPPpx3x/m1NJ
L3qpg3PJUxuzPlRqo3+/e3P5neoIYwPr5JYR8bPqiZbADwi30h2py/75PWkfJErut59v7Qfj9itQ
L5pchxS7KMIU01qqU7Gcy2cslDHxUF9KHqZqdT6oC+goRNczIbh9jfTmdABAnNmAyQZXtvhT6S5P
sRpXuzep7JKLLuccja89gjaFnDzZcwIbP042EPdGJfqpIB3+TMFQzIokLcC7FyWC2iZhrwZogoXY
0imCyzIf+xG6NbaPXHwfgkL0v/A7BML6AjLYstXMb7BBCaIDvMM5PLt8IUQQRZlJqcm4Pel9Vk8v
9J1YAeV51RYoJ8+dIqmg4MQJsA5vgRPwDhigeMw/ryZha9VBuKJtpoKb5QMmxTbmNpK8Hn2YkxNC
LpHo+glveRfdEDFiBZ7uJrrt59vCoow74EA6lj4iM3V0BeuCunwF8eYNtq/pnJACLHKpM3DGAwy7
PWmp6CG21X4q6NMJSj8zWHEfabB+roI+cEBYBT1d9rhLUZPRdXtpKvhZ/YS7hJvcS0aipHTPyc0x
6T1eD2Yi6eAORxBz37dH15WVOkRY6u0MCpZHU1QdeJ3GuEWG7r76gUD1U5VVGsK6dtqInAb7MOmu
rHNmTNOLEBsKJs2j5F9NEBRzH06oj3uVclLrjpd3TEWYCMsiphBp08W7BD8b73cbXidouY717NRb
s4Lu0E5FuKxJyEjhlnSfFJDUlKxTvAmXWQs7sTT+ADuKWjWDBgWR2Gkq/Q3qWCXWATyTe/9OHIIK
QjGjAsjJfShh1OJqCyujGKgITeAbBY4CP6d6YE6DD9NK4M0MsFxvesfLRToiArI3A/1ivrGl2pmd
mvdatjV6EPNC/6vPBCYiAGMzi8FJf/t+irvC+zQ8XGIlCweamjYp/6MtTKs/y8xB/TDkfGctyHoq
G288qkauF4KybVIQwc+BtSZwlyD9BxqFjsQPqn2fYPpLNbebwc9yJD1dutKs9oUWkcte1kCCdALs
lfN5qfLHhXvqkH6emBe2pVtgutmGJsOOrM5i3vTYC0YXDZTbv8z7aqfJoyPOkrFiMMWrgkSZL/UU
t1FNBd1XRZxNoq1rxzJlkfJ7xU+gKzPcbKqBFVIyt7UPk3snwHPa3EhRyjDhVNtxjOsUINijry2C
hzy35Gh2VIoT8cmj70fr8iKxJtv8aeMWllPRN9lakX50O7fhHwpNDgIkJqvgncH6dw3SjMrZbCRb
Fj08rPfSQy7T2wZhnZOBd7FvPZyWQ3rw03mP8qYy0tKwCyN8+oxnZbf5s/znh/yxTQFQ15Pws1Xq
q41U2eJOBNqoAupLFOcU+GT4dFUC3mM5bx2fY8EtSpXuWtxih38rv/FpA8YKSAIrqMxgaNh1Cc+e
VoVZTCQPS+VdmWp3Gl4sONIJF5kyj7dM+wnxvLEfJ5Dyrd9z38whBX3XauxCD6619lOkswDzj5yW
EpzrK/gKYayp2zLGuIJp00k2nfMpjB6zVafP2I+C6U17gYker/7svYf+kVNtfdsnZPUVj4spiVjw
0PqFjz/bBTZ8M6IYWuBND9b1kLxu+zz2Ul6ht9F0mU0HtYz6muqT/101FBOxDARPmoLokVeEAu1U
0hLroOxLXjxBQaMW52k3uHni8Hd9xzd0nwByzOT9DID1CBTSXlP+z/7vkF8uXvPeGNdluwJrEOQ0
RV66neBZ0Jn0wHtCsnNRECojrKki29MUUlgCTTWJW90sX/Af9vfhOye9UvVVQkMbFuF/szjoEwe4
vOT4Exepz/Cis1qjaJ9mZg0OEG3r14w4CM0qTmTLJnsVIOpstd8ZNhskC363UpOLY+QpgZ/YZrKk
FKQYcav5/mLP1Y+NW6CG1Fo6tmb5fBBMz8coVKA8g/h+sIWwKysJlqjai5pNIsrqkL1eXwFenNjq
E/FwMb2n4RViXdCWk73a/aLV31jdN3rpvE0krFpA45ItVMI2WjZiTkSPD/YydlQV9JoTxrQdPGBF
o22Pxja3bggRWN/9YK1dLGCxcRdfOJNzct7+EMoBqo5X+dmdsxrW3+XN+xoa7xxGI/ofFH90FwJX
fyqj3/cIINqAPfzBoljdmTab1KzPTjn+g2hchjYZEBJmAABdx5D/dX44FNRL9qBi4P2QWrwyvMdj
vE9m1Z3BcO0eQlhDfmKslOFFA3I/1YRe0J8lCbLeMJkY4/yb8qKBTpvJhP4H+NJrySCNd/tWqOd7
678mfuHReDxKl5BVH7PWF+dFN/UWIQZLRyto4CUyQlO2EkELo1+X+tPPo/vsIbGCVrnJqQtZje1i
UmOSvS9PUqu1cOEjGlAVvq2IMpal/AwCo5MNNB0bjggKd4AomF74V+Xe2DzPSa7Oo1v5/DXZUQ9d
JEN2AExJZWPUgYcTTknv9JTm5wEIj5BkmdDq4Ob+PRoNP43HJW79+V/GEcFqiOiAG0asvR+WTdeY
n7RlmCm11GMZejPDzYeK3CXL/EllnHCHi2kSSTElXBir7dYPquyHWN2ExNzG4Iu9AHsuwGuT7q27
iS2h4Jih5AxJHbPSOg9cPqdwsaZCPFmeLh+1OGo5GEm2jdS82zDX9eUmlcOJKkMcvciCLYXnq8cD
OmoIJrZ25fznI+1JyfT72MXU3u6qjaJBbQX8DBIaGuHed/3uMjyXkp4d/GHg6vATEXUEZb4wi6cc
DKNyD3SiqWSjiOu6w41kYTL/Ec1kUFFz8EQNRqhsvYdqnltPUpd4G0icu8MYlywTBXkyFlxO+F0M
eyFkEP4F+QPemkAbvy0zxADCz+IJxyiuzn+cdh3htTQkjq1wWxC1PcKYs/sK1z2cEx8LIX7QdlSk
0j2Cy7FItcEWxI3MrU0kVFfWPycGx0ZZxK3j+BtzjbNPrAyGB6uSCkGbPMazXoEV28WsZBCU2br6
Rv1A8wgZDQfCkncUjz7SCfk2/rMsd0sdQMFXNie7/YsT8CYM3LdJJMH1LRtnUdK4x0t44nEQErLq
Hh8oms+nL5bE3Y4CCAY9RJU4zvqFw2F+CqibB5R/XRZoq2RRHRRRgjwqIPsvoOnCOK2mkkuXSWcJ
o9qaM4U3UFKTaAr2K3q04Ckgaxvbd7MBsmWVnHdKCcDBgxHu9wylMemOy1FzQlM+AJy0tdWjxlT/
CIC3ZJBeUJU3YlsVln5NR3JQxX0sXEDA8JxBJ4oB7jkmxQWEDFNKDfuleItNzxY9Fia26/DUFfxW
SHOKqwfMfLMZiyd+552yvU4V2jgE73KAYboFkBD93VcnY9L4c/YaqSRZx5Zgro5xLWONDVz3PVtR
v3N3i236ZFWVKvq8Eh5tuJt14FbonOjiA9ok/k58tZJqOXU2GqhNjWXJVqe/1A/IxcVrZQiQmQtw
zkrkxmXEp5bxd9jcXwUUaLPjymXJFR/2VPka5A1KUkzbyvDGdVLLOWkBlNfCAonzo0WDe2W5WqTw
lOKsKYVcbIzPZNU0NAiO0slGJc4PCZTGoc4MfzrzNgNl5VwGsvRTTP864T9keQpsxlOcL4bK2xto
hnN2dZJgUqYyTVNuYnsNBOcl6qs5PmqVn0Ek//b8thqUYsCKk37hdT2bU5HaA81lldGD84C5P7aS
7YwqJX8bWW+QRbaeqqIkkkdxv+H099MD8KywdvfLEnqfkyA9QeEtOmVJa5lLhGhbJ74v4B5IFbRW
4W2Y9dWiThFmhPamJ2LTZJrLVFLkEzo5j5lOkI3DOOFa+bY481iA3ZhzMYsuiu/pSpmEome6Nj3d
uwqkKl9HbNoC6SHAmlSNpMpmyqAQQbRbYitRm3yI28dIwws8QbNoSK8CXrG0SsuPKknt5kMVD8Dw
syiIiC6LXQ7oOoxbQN4a5TBM1U76hHfk3XSlEUB5PFfjgfG7Zj97GZL/Q/1w7cO5ClaHfZxFzr4U
1esB2pocFwZvFa9mKJnRdkzAU8coqXXV9ttIVW0JlcHJBPjNajCe1r7BGLkcJu6nQhuVQif+SXA2
deCFIdwqNQ8H2KYmeV1Ha2LuUvn8gXLsdXeBOzqK0ZbsJ/99vb0u5Uuuha1zDItIp0A1rfsyQK4k
wJHa3XF85flGqqa4xleviwN8IgSxrTSjzMKbUfvDqJqa1EzJ+gUHwY+LP6IxAymPoSj5SOeWuy0W
CjI4V8uQzleImaYoKCJs6hlFyzpKkK30oUgGAwCC3aPIGu8VIQ0zxgklOwzz44q+6sqATPg04KJB
bDothmTcLVh3oCbpIiKgmB7xkfw5KhdLv7EokIwMR8/WafM+q4h7YOx2BIstD6TwZ3JDNJW8zV5X
M0aa+t6T8NUZo12ErhPaTob5v1Nut1FoXkfnHRyghrCWUtDfu/lHvXcfZdzq9+UPC26+u4rEPkfp
XLPEAY4lhVkPCS+g4BchcldBgmLdzURRrZGVDQWGv2zV2pc/I3ZDkZN+j3WIfth5u0wCYD5eNhG1
RDDK4xeJEjTISvWwexq6Sn2AaJZA/XRSDL8fU0m4zLVjrJNW6n7lIwQ7kqhLteD9YygHUw0BVrCm
KktJcz4Ytjaj9oTP1F2x1L4IkqZUz4I7PgrHt2ybkdVeev+Nk/EmX7TCZBpuwaR2MpZsPjGkJb5r
qglGkKdzcS/VIJN+GFeTT8/stCi9IpAN2JjFMJqExcWqRrSF6ZfouE/lOXw1qg0m+msAvh3g113R
LQO3YoD3XIcsVJFKJumy3eYdYVkMcxHpvqtz1E29xzkP+L3zDZoLdh+H9CF5RUv2t3tjDcggYzzk
pBBah4ATHm1nGYMVIiRFsIDFAssq9MCrAOuQLJpw/5irIW483+OzgqXtXOijli9Q4I9x0bhhxyvv
BnDerM+krhLqdIwSp6VqV4lkcPeBC1n+vMPdcsYmfFKen8kXqkXPbNfZ+JrJRRHCg2Qk3juWdYv2
hCJL4c7ZC0aQjj4lAGKBXF/pzAVQFtqbv6PY1oVL/yjegCYoFHKsNF/LqW3jm6GxJI0lbDfbs9F4
6RsRJiPLd4Zo+mtf53kH/rkBPEVwd4QJscPrJMN0jLyR/DuKQFTIv3r3uj2Sa1kbVy0R/BKzZShw
pAIZQnMf46erNhuQtGzr65Ay6aeoFGOwz2uIaPcpX/uzp7fk45IxZw0J0DwyCRkJUCnflRu4ujdv
ce1I3PEPmMaADVx/mRzX/il98QnQx4RJa4VUKnSnC4wDorgZH+X4IbI2+KXlq8zCWq4et98K56XS
+WG0S3sbpxn/uIEI0M4v0DQ3TcCjYflNSaCU2yErZFK4z1KWbBEiFrSXAgApfDAuRrZq7dGV6LZQ
16XZ3IBDRijksYcNSQBnjsP9YotqqtxS26AWmlXy9XAEMRyTT2QkMb4NablG+bR7i8c+5jmdjYDE
X6/xdy2Saw/eaYe1nLGYtXsNYpxESAzLqC/xl1nzUSBR6HJbaXHVY0hcbJxZV8fIukkt0zjCCoWJ
Y4/1qIkRbZGEkvL/NUDn7xl4XbUzKXv+8x1HvDJrqNxnKumRsUIKKm1/A81uVXhYyYWhXh/2UyKA
OB4ne5Wf+9GX2tvd0HIAOUAXTZmBgEUL0gM2n3j06kW8DONx8jSGDcrzwx4sm47rpY8vgzXaPqXJ
dnRAOlTitYl5x5xlVzRQa05RXdggL6ibeTMDrmfQr8LjaacrA0lKutXkgy6RYhARpDDHkP4muz3o
9FcTfnRx3YCb+/HtjO0/68miRHOE8TUNPfVNZHhwRB+o0fOXz6NzqLLMBVdrxX+3X1oz+wniv0ay
9Nr+93zZzguCjiBh1fb2GgaTDOI2ylIPA0PvHThKH0H1BvM5xck35S1ivxk736P2DGMkAVbCs8ky
tgzyyQxfCUdwnKQLT/luLlwHuH5YpRjysUtjqdSzltwbLbwIQGJXXPi8ba5ZezetT6IDhB9slnQ/
OFkPa+XLWWQL+HTsLOmYFBwuj8dLjMYRkYNhUEwFgOuUe4BzNs8gmc4KG6Ofm8ZbiDEKGP2TVzn2
EP4Vh4OJC0++0ZEP1UH2uuaJdDvjn0t5dVsrxmxattU0t2r/9wzFHBFoQWNtdNIT64DW7Un0eqO5
mP+y9qNsWkO3REx5UfcqAXCCzfYy8EgKGX41A1HKJYIdzV86yEBPTJyVe+St1/NpPDC9pt72m792
CevfBtcfvLJHbKam+MjG8PjZ5lfkUzpffH/wqW5Ouy5B30O70Ir92mxli6Wx2ZntBBLFjgYe49ce
JT/0JQHvKvnxY78HxNl2pn4xrjnGhH0Oy1icHh3PL0MPIecrjrqhpUeoi+QN/mrB8sQNcxXqOf07
1L5T/0Jpz2bn68CDSuxsKlML5IhC5megH5mRTBIOMcD94CXwlVWC57ELZwkBvLy2uQDW2kEAqDky
yLU695lkgKLbf7hprYXfBs/rsiAQcIiukL0+ZkmnRiN8IpxnO8u+fF1OzRHIr/4i/kkg0R57lMBC
nNfqd6yfUjBGCof3PqkjDFLcKxR6pzcVoFW91EqFXuP5Dz9cHo17HV8jrexmgAW9bvf/BxWc5Ctw
HTYf5iHokqDFLdGOu3nqM/cTvmcWNq6qobaFa0pUAz7v81qSo0Bsbl93TShfBojKmso4Zj+bdhK8
Gjf/7D6Awy3S87dM2vNH5hrczpbOm2zUyEKtUjW7WqicaPU5qFJs23o292VqGx2Hi0YoagvO28dN
0qCI1v/epJHu172jmmjYMbY5ZeuzY8RjWj6IEgmgxb69BYxVCus84LcJb8NmGbAs9krnDKuTX4FN
IvOZzm48n7kCWAF1t4vE+6T6P4q8ij06NbqsUzd7oGMCXajwKLD8E9dKYyW65mT+CX4y5/+Y8MtU
5jn4kS+9YvyV6BPabbSs52s9JlTjTzr/Lso/HFHHMMJLUIRhCXrYz+vlOuVmqmV0vwA3W/zy3ta4
7FMWSyQ/8qWcA0ArHXYuJBOc4GhY2eq0Z58D7W8JMSBq2JiRUaK973jQ875VcIYmOKjGWNHGVfdc
zc/ywCJo/qwvP3Xzp2c9HH7G76AW3yrraQt+5ilXQL8zX0vCN12y5Jmi525UdV7YoHDqeM2jNpGM
I3Aa3KDU111Rug6tCBHgxR64qN+YJpaLL6XNebE1IRdUTS5z0qfZOmypHEOoiAke3iHC+0OoqjZ1
X7mItJ1Gjhzi5+OJfA8Upp99meBnRAKyNKc3snJQ8J1wSAABvKjt7rrzW5IZI4WkQQNmvVSBRNaN
01J4nVONuoPZgRjFsZ9rvGaTdSD55YE27YQB3h8H0noez9hko9ljtmFHhtZvh4mClGwLps4LWDTo
5so7DwMc5Bw2f2V4hKNUTK20rOex9a8NZG8sXc4D+lxwqKd89e62QVWac1MwPR29y5yvsxAByn+s
DA5jdrSzbB+tv0pil4uzrSfc1ePyV9+c7QEdJCobpCl/ZLU0y/mGgXfS5Oy5aG2wZFQxmYmCHb4f
10Xd+d8LXeF0zLnI5Fz5aBtTeBQySF4h10ASXmE/j8jk6vF291vrc/OzHbJXdPGOX1uAumHu3Cl9
FPifWAwbDmo6zY4GqRBdxMa3YykoVdIDTn1n9TjYo88iueU2BjQIHjRGKGL78QMsKc0FYRE1sBwz
mnJKAP2u/zvWOQa5kJZ0Vyxk2SJHqzf6OKnZDUzzgW3ZwfbAykoPKYGE2UWozL1cERaI93zd6Kms
Z5qCzv/Tb3YWw2Blc1psEUnOSaWxPKGV7wu9km5sIPb4Cacb6+HfEw6OaKDPyB7zkV8QSNRPi3v9
cqBEmf7LncJLNwTOCUQDhKB38akkUIeWpQi30qLZzT+sFNa1fHLhKY0wkQe1cXb6CvJ8AVy1koft
1Yr00ZxMcDbgC7qscoy8UoQc6RzLcXryA09huY7TDw9Z2E6xRD1dn1K7dYi/k2QIWOwHKoU2Av8H
EChntJ/dpN/tr5SSzC2zbnYobP1cy620fIZMR8qWho7Sg5RAPq+SP5KErDZ5YNPn0EMbMBJZMqWp
0vgxEbkMuQr5zf/e8Ja0rAu9BbtUkqqvfGjFqANvo0+4fb4s1cO/hixphU05Ywx4uPbjiN+I2Uw9
DifWwya4a75qv7BDBI+T9KnKouWuXA2Wu2uaQu+KfGKzv9ZSYTVmN7xVsEx4YHEeCrZJeuPgembs
1vtkpfyWcbhlc/4pJ/JMzVe3JNzhgtb0z77ViESCKyVmYE/X59ONQxpaVwv0G2nqlXTBZzDDg83d
vCgsi+Z1eKbipIQKz6rVLVNsaB9YwvsmdBBAGMkiqeFN4i3YrtJNWAs8APbZgOLp2cjrLA3jRLRQ
V+cNSKtwKZsBnzvvoh+mgQK/BDh+xDomUDqjY4KFrJANQneijNr5fFLe7tfRngJ8qKXt69LDUrYm
oB/5pOW5jl1UWx4I8EgiTI1YqqJehMe0eUv8f1kPXMmy+Vvy9jD7l4sMVj5dVMcy6Y6gt2UJbKvV
tj6DlDlpcIXthFfJ69ZTomxDc+5RlSODDJQHisUyCsxH/D0dQbHWB9qP1kmF9qEnPqiy5De3Wv6q
b4v4BmfF51YPmvTBGpgviyeqzMQLQZLY/44k7/nZgPTYcq9yL/n1Qt31ZlHtZm+WG2ol58hlv1JQ
QNcoFXdzrWc+i1hznty65VPZQslcrF3kykjeeqs2uHDB+JUtVa8xOrCDS5J7+BABo8zMmSQsa9wO
l18ClVaW/57zaKvojIZb2a5EpSAvc29gPUio3ULNGvoXUtZGFQyrRYfcatqtCdN7K98rEGyxFpm7
uavTRs3JOXgBeHMwSLWC6PrdYy/yZE2yP6LbO+RguPbFhIzeJ2dlMLwTktVyjylMi0XUxnfL4ILT
h8qY27FhSuystRSh0V8M/dL+2wLtalBH+O8We8gTJsTtBAGV0+4ppwLrCFSNOgke4IZ2OtEJAwy5
CdrhaegSK9gqDDJd1C2DifU4CHubMl7RzLZF7T5/qNtdO1dtLEmXhh+SQ+JCBPVNGpfCIEvlPq56
lJNUS69AhJOt9duFxY8CuZlxbk+svD09VYczKN7lrh1sJflxYm/iXmJeE8Mn2ksV/PmIiqscZWa2
tAzJtV/4BB3k68MbxO8/vhg/IIJn1gHxpi+fTKsd+O5qdxmlmMGPuAFNPESm21l1/McQ04PjLccc
Co4v8EGbV8RbuyFus0ElBz4LrkE5aPhc4HncAGO8ydjTgteOsPaMDZxH7kH6M02GWpxiasJZxsuK
moYR5TaEqPYGq7c+UWZZK4gPUWga5RqMLwUd02EmjWC/pd0biSPIHD8yRs2JQfPV9NxxSsJ8xoVY
yunHCSSeG97jdawNor15AcKBzWiYNSBf1AIDcsFxlIrxEOh96sgHeFooL/LDScsBoQ1QD8UId1Ik
hlJnDaHg1cgwN1VSEKwvlFkzUVtzzD+Gk8Ulr/f2WSSv7rq/5Kp0gRpQ4RKfjBLNNfWCvCA9nXLt
HJtynCkgbe5e0T/6vfraR2KjQEHaxg/d3qjzvk2w9bsvwEmNOYnCGizchSj+j5bzkXqgXCAZGe0Y
20RZVFL7RKWcvz+TfbpnLR77CATK4uVLBVsOUcMkrR9Mh2jSAdwVEdLriFxtzGY689tLmGXvGqPZ
KxG5kBYWlwPwK0SPQ3AmqHrV9IZN9fjtwBR1fnrXRRN7gPvQl/uy9+LM2XFPSEFgDp0aGbyw71PJ
FiJ91BZG0MsYiFHeY+DOVatm5iXHW0Oi8OvaUIJGKLOBUNENUEsrHhuT700ry1Q1u3/ajPAkIXPc
gp4xb/Bfu6BTDY7erJCNaPjlmvDQOsBl31KoPyJzcIskr1bKTKQMg+gCtkWXr4VepZH3mYxjdxTF
hoCJaiMS9skJVyyHcXOXw4bWremT8rTneqPSUGPOjpFhRUNbdkNSscI8hiiXIlelsFqflfQYYCPz
bU3bz5qLOw/R3NPXPhsUvAWv7yqJZiPdqYuE7dLUy0V1r6CeuR3/nHgtVma6Y+hQwtEFO5ugiRaV
XfEE1kOhmwZ6dU0WgYCDg3M8O3Tl5p6oyk1jQQrPCNSzmCko4i+Jydahk7MgW2Q/5EmmGTPh55ns
Wx78SmTcwEcJcbYZC9joHbxMMq7NHA7jRWVwMbcDZU7BGGei11PEuufqc0GLTOPqnDArd8G+UGyU
446YxJf8p85kBie1pVMr68VKfPecfd5salDX5la217SHb9kwE4Q8G9LBmtP7lC3On/lbDrxbNdAS
6jZX/CKlHlxPQ7tFNM9+XndqZ/nxCIEpZwD1zmkmFUKn3F5RCoijeLvZDhw6Xysmtdi7G/z89SHV
WGCs9A0TEjcnWC1f3BCQfQk1PsSzYresu+rtfwdV3yDteKfWbDdPPn5R80JW1hp9oh7XMGQBvHsm
9H/jNcajAnsc1z7c6tuFQwvUjxMDJqNeb5fKNuioxPtUYv/2OXgE5z1agESx26EmrEmG9JmSmioo
cIoSVPAFjzk4ATpucO53B0ztukErgqsWNE7WmXBpvAxVGjsefpE/Lv+XH3mnJwh5f1osN7C+khhD
9l/u6+tlgMQ4R40jmxYdzwP3Rg2X+xFdX02QMImXzH7VQAePG59K3RmG475IYZlIxBDYkvAN7xCL
TwdEE99AOo4xjkZZW9Pw7vleQ5mNcxNa0S+YK7kmRQDEC3ls8USFpFTn5OQHK573cjFLmMJQ2igW
8eMRv81x9u4CGLhT/sCXco0dYMGoFWqZrngv+UrApiJgkQrAboPvczIaKyLqeohy/vgw1eQicU6U
4V/0bS1W0HDRrSq+zQI2TnS9yjCa74a3Q97oaJtPsj4MOH+eXO3p5R5gt2U8V0LhqBa9LYphTunt
20/pBh74Zd6kzCgsUVj4KJWjgt2AyDeNhEoF4zcB9r2ndJtvPB97/Orog3wBiDkuIuVqu9ksMPhi
5bgWPpUnx3DUDA0z/0NI2BQjZMA+kXbG+lisc7u5g6Oo1wlCKKaSbZh4bf+a8J71h9f9yktWD3yL
rsSSv7U0DSA+Y3v6VRQUwAp9t0R7EvpxYpNkZcmus2Y4KbccKe5Hqc8USafZqcO+K/b86VKnLzl+
cPM2p8pU9zBT9kqUFdm34QTzv8ECy5eeky5VMd84xoYEwFsPBrWfMMI8/x2cNMxBC8hZHPXJZcJx
e9hpvUrRRtM+OwD0/UypWHnEJrPb0DyIR+PSnx+/cJzZou3whx3HARvvSa5qOcpKX+XxMAtKv7u2
HC2vqA2sM38F1J9zCX7Z92ew8hKXKgo60LUjknKN+s2hxWFniiJgt9Aa3i/7ACiKujDSLLnosh1i
dkr6VAsQaV23Q0RxWMQdik5KiM2WdnYGmuSKkAQ8g633egn3jkSNqx7n3TKtjvjClb4kPPwRZsXs
hVTdXPJhd/pyywIAL9R/xPkgjbfWrkC9QQ9S7RTitEo3MUMVsqBVQ3SQFqxP+yLofF/6h6cVLdGP
hMsbOZrOI71zj+7m8EOLTLDn1wTRQV7Hf8tlWiaKtn9DRKjlZJM0q54dS6eXc/gQWMPMLKEjJbgG
l88ZZeJtWq4bdfFP2iSpAD/C1qQ/pjPDh9NJH91KQ42G3zqNi2otc+DvtUdk/SbZ9mKYMXsz41JA
RqStmCYs2Gyb6SW3pkQm8cuWJiM3kF3tXGlBfmRRkfvkVM1qfllMWF1hyh52ABlhaW1xdQnXpPKO
AOpexh0sKatI0vw/ftT5hS+h1/HFuu194BYJtiR6Wam42USnh/8DKE596thsQlh+RAGrc7eLUbtl
67vX+cMGH6TPXnCtvdPQ31CnlpSryU5zFdj7fVjq30Ukva+V+93npt8A9oSUtLPEu4KhLMoQ8y6q
zz7WUSmdqyINJZVGmL09DYhIKOoBswiMFEXATIIlBML0M4zPIK8mfp5xqkezyy2DppV7HHOy5WR0
H7ZWxYcN59eoEmxU+3PH1EAn/o4uhxcKNF2aot4tOTBdPmherCxtoqEKh4bJ68/91dvdSxF69st7
GAH14Bg5xVS73JlDlm2+PYwnv3DNze2g2PS/F6YPBn9G0CJHX753wSFWv1mmtBrfyAsf9C1ZIqWl
18Gf4g21vqrj07QdgzBhmXaahKvSnOInQfpUHyDi59lRmnqAawamdTMS4iGzTStwEO99tPIDOhm4
J7uRV13XttD+2OGH9hHXPi8VciIw0u7hYB0c/7HJhkI2wIsr6/7pdL4nDjhb2AH84IiBIggBalT3
OFWrB+VKSbqSxMqTO73F7Az+zwO/TFUM54rokcgM1v/O4DIl8svG54MSXKEt7QDq8lFIzWzTfxZI
FA+D8SXStucwNMbfcmDmLHeSsl60twreUXMUuO2Uivakx2nSu3IORqFTqz/5Dd/CRWFR4P7tDB3X
XpJP3AeU5YAAmalSPw5BC5/6dQComMZIjLlxqVgwvSP+ZNpUZBDtkIsUGoI1DcJU2CRjzqizmrWY
nWkvirH+YwHPgNZeAYcxSRa2jPASxXncbvNB2IFlX/+6Q6N2omyyartU4ywOjYtqglvcfWbsO6mk
UocbM/H9HuAFprnTLa2Yyh0PcVaejH+ij/CzPS8kz4ppmB5zac1Vjmr1ZEMamIjdTsG1Y+Mn1jzC
tR5vVdNqPn/7YP+C2YyTXu1H5JHlNcK+h/AghqBPZHZ//2bkUsBPehDEBmfxHuzQ12KKUNlKO8P7
bZH6b8BOw+VAit00d2sTMU786RxPr+9Fp6eRtz+US8n48Hahfg0CzIWlBDAHIA44OZmyhVY5rqoM
3+7o2mP3cojHVtIbHlLZP0wBWe0e7qZE3iIUXqXPiz+s0eFXc76hGNZ2C/Gi8jYme4oKKLvj2cZN
X5ruwq2cPjVnnejIXDCWjFkSkyxcMsCR8E/4DkK8dZOCt+JDpbUcV7uIoT0z6hrJNY+xES7rPg5+
ANQl+4AwnQ0BvyD92NskH14oBgCcZss8l00w462mSB52cizVmN1CudWBbaJ2qK03TD6nLdff5iXH
AA+vWK2Fb78MSx+AyRqh49YKqHr2KhBpQpZkdi2Os+cUZrokiYjdanEvptZaQ5dVcP5740LBROIG
tuMCipcdSZwR2/eXAnhiGgQRKBagWEjGp1HowoY5Pt8kkykFwCgiW+x98V5J9IfZsY1twjWlp2OB
pM4sxm9tQXRVAM9bSGf+gJhLXUXhSyMXdWfge/TNAKlzLXvia7TZgSGfKd/U4Kde4IZV3r/CV1zy
C8MsEMoY827MhzdmdmHIiGmNuo4VLrXnoyzTtNx5l6PSGVX0QVEUnG4IAXbj9+o9QSxGYUGNyqeO
kd1yLPkW610NVGPEutuZFMaRNtiGpuXHCLRVzpxzs3Ot/c/yK/sAmHShw4wwvcTET8NX5lhy/kvo
fta0SCUk5GOoTBxqkQ+HGb1OpmeEWajLNGkaW2y53KWAzlydyebuVfAHjYwe8TE8a39LBRdemNba
PW8Z1cGjhRnerL4Rrm99ASR9wZhzeaONXxuPmiDF3EaWfV1ffkoSwiN9ZitpBShlB7Ez7BnoWLdx
DpTp14cYD+464Id6fnR/qMYV2IRDcihsbmQfFPR/hECI0urssaV/F/sUYB+QkL96MmLoh9vZxziU
dcIExbRFktJ+s3NvMsls0JhO3gcsvr8QglPiv0JAbguQXknePynNMAaHYRppjyxzkU1d2QGa+hSa
XA2lBdWrkHiY3jlsCUzfRQulAxe7wrdYlz5kL7zKiqM53AyhBRbRYbkCIH2gPSsFp2vaWpDEZKNh
JKl3OoSiDLN6uMWn2aZJgxOqACEM1kLhi7blT+ehGLUTLPzYQ7L3Mj5fFDiOJmw9aCmoLQKqilzr
3lFnoFIgY36lsjMNfV0buH7cJ+Mkl02Dky9NgaVg8t6AQykNcqDpbq5bMcdzlXQuqsBiX1kDw8RG
NAq871VjGLQKRvhAuFBemciRGgFG+eoTDex0UXMy+9EYDrSi/yKcWylNIeU6YINaUU9m9eLE2hO4
YSRJifsDE+mQkk+tsLWqMOwJZoPnxoTRelI2DsReWMYZH+tHC9e/j9upjzyCEQZxc6/sx2D5d611
dWe8LHIyYO4Afbz4xGLhZiOrZeFA0/T25ZjXWKYKV7vXDMbEF4dXz6pCMTSRFyqzm618Wg/qfx4e
JgClueoQE5ephp8bxtsQG9Tc6uT47S9LkoDZQ+lWYZWnmZ8cWXLchF4TxxGOKko0JK+Eib2YxWqV
WZ8hsPr1PoIKQUEtF/CEi6q2qOcYM30TuSqI8gfGi96Yj0Kt+9K6hcwePzqEAxiT5h/u+/GANnfl
sZrTHy7JqqDlOFhgQTKMvk5Il+hjgJQte0IrFCXGJ7r8Fy1xpGeEVv+uGlMjsEb6KFQDGnt+8FKF
nWQVljJltEUlAKTJ+5daaQYYJNgbjY3KB7GfXXnQvblKXDjZcmp1EHU/KPnOeEZer5XMrc/jpVeD
Sq8qbKRWwYnkB2iJJx/meASDBN31mcX4eBnoxqwAt3rRH4iCjqKMlY+CFp/ayAMkpYmz8udKrrpE
KYTflezoTxInDTBtsnB6kDPzYgXTnUZT1xZ8ag2pp0nMxEruGohBARMSk31G1eOkrK0DVDeEGr9K
OJjrN2ivbg2ogFdPHkYhmAlHoeESK7tLWuyCwka5mLTKPKEbg3gsu4hf/LpOHI4pXCSIJ25pO6vB
NJ7KYT/hOFqI9O4JuOXzBpeVWlQSyBTxzvE3lZseXP56odI9T6Vo0UbtH1VHF40leOeGjIoHYvcX
kGRQr5QT5xWEDqzjXt12zQlTehprVeDsnoSrprk9SB84iPJh9dwKGryXfvM7pVFc8YJwv7r/JEIi
ehqcz6itzhhhFYniz0Q1E/NaAzMDg0CheQdUapz729DM38aKFyqpuwLUlRI4qoxJHFgnC838JA6G
/UbZFW0d4KSKaT9AuAL3FGC9+zD/aeTO15SdTQ3fwjpwYTJiIEKw5pP1mXDzKRgBhqlezDVnt+Rt
ryvmbZx8AY6TGXxMK7mKflvMGIyMayb2RsxeuZ477sI+O4imPmr095c8kvv9ajy9UKyM7reCS6xq
CzLoEHI2nIqJteQZdm3yb0Jywvt8GM42WXHjM8Q5PSfq9gNuET8ZvCcQuINCOHJgCckgZkZAXEXs
ALZmUnVUJmzIKAMCRNkBniTtwUiQS+2N0SCoHO7oHKn1sB5Hx5rdDym9YodYNaayMy7Rzp48TE0m
p/nxKjjPYQUpH9ssVz+PZSSfnLAse0UTTKBMcRaSV+A/Pz78T6gGoZNnWCXGUeK+MOCU5sNwJN3Z
hQKQ4qqWeU836yrOwGJdYUQYcSvdDF4g+Js0H4hkGY7h7QiW4Bh2ODQ552phYyPayZuLcqPa6ZD3
1mfThcj2b3TsOLLBIqkNMJ63+dYs8fGtClAEmcGGkbE0jqAszfCZbzHCvAxc73If75MgJsDUYe94
G0ADHKTr3uQ85OBD1i4dkIm0vpf07t4o6zOnL0Qwam3d+lHi+NZX6YLozTX7YmXDHEa1azvT2Pmr
miabC2IAK1jDsJVdLQoyxDKwt1KlTFEJAhcP0gdVLJYvY4gtSGvVavtbAtrWCom9+tZjaalmiFVq
N6Re6P0az0MwM4i5n0hJGcQzHpFoWND5rgpabZErIRgQh2pf6yyh415a0SYlJkg6pRe1WSx8Hq42
Kzwg1Aa4sR1D+Wb1UDuFKVnrKcULoDPWMGXVtjL1Kh7jeGOu55kutcuzcGmoK/eupZSBu4XvI3q4
ZRaCwV27+ejb+YNMjZTekMdoXgBQ3rBwTdY0v5Fs6+MbrKPimIavjUyxLS9V9ePTXaQ8GqUsDhsk
JcMxF/ILCmlCLYbrhQppUMeDPDAxjPATY7x2GbpyRdhGNftEWCH6Ed4DZyDBf89OgaymRiqN7tBo
pd+8zBOAEkUwhD2KiV187tEhFvohV4TiyjcDkQQSTfQhPN0buPt0KLpz9romi2o91NpGpOaVZTHX
YxOGTCc98aYcaCaMgNv+NmYAX+YDXQla/UbVouJbalJoHe/EF6J0XHz73mJJgz6Vqni6wZZvXWLt
LQK0FUf/U9arFmkuJrXIxzBAkmHBYMKify0PSVr6js6NodoGpnkc5QPQ48llWLuMYkmehu7PyXFM
sT1MveryjRSDlrDVfWiArFa203nKq/outvMy1fsTNWh58jzTc81xmm6Vptod0O5+2CF0cP6/ss2l
NHSSRey2uOb7xRtNp99+T7jjzmgdmHBLNsCvOqjjzupOt7OjQlUfJSOuLGvPGeWXrjRZQIUIecZ8
nBUGoSYcZldysCwA7bJOzjZkY4+rWvaMnd/fg7v9XdPzsehEbeaPLcmn3cqEOdNrSK3wqm0pXgsv
tWYfywEiygvAwbHmOG556oACVxWf35qg8dNzNFANVmkNuxLUO0iLHrOLc0+FsdHjAJyxqylw5ohH
gVezwwFw1DWKrkoERrHqe17qsZjP21nnjmbmIaxr/ExSOMBmSeBBj0QyLHQ6Ai2cCe6LXCVmBUrS
KhKCFLOvJsAjXHe7knuL2S2ibrKDbRFDhrgd3eIuDaZ9cqtGpzK3Eu9401MQCXUY84ho8Cm9qY1b
9AsAs4QfRal37cE5CrJuADsUjAuJNyZijC0thKvPevreyhXQeH8Ot1OtqEteESiryz0N6Aeyrqf0
5qVzxm78eNh2tvu5kPzoIqms5qhfagGCtu8L6brDIKg30rAASEcOCmF0+YqQL/8MEStGE/TKD2Ul
RGgpSLRc1/gx0ei6x2FVZdjP92omRGSQYoU7vbZOfEN4of4gfo3OsJJrf4QaW/bFkLJ7MfLNhR9g
hCyWuR/lambwMlkwrJa8LUEo6gvfu4cwbCPJQurlAbNZOeEYoj2vFijStvFdCwqKRj2O6rWn8X9b
cQFp54AlKXF2DYNtuLFyM+Od+hiLFx6KrzB9KRP+JP4c4rqKJlhXGRjCIzQI/3GnKwJPRP71bcGX
x6N7JElGjikZWZrvJ0xJ9PxBkZgM3UsMoG5lXnf7k1DLjtHgj+IAr/Rh6GyPKb35jgKGRI1b5M60
mVeZHjXdbtF62aUWPrrLM7RE9CGAxr6H/sct0tOCunUaLxHraEkdfFsCHHD1E3/YVp7XHEhkMOpD
EXP77Dezy06+ifmZPO6eBlC86h+umHqwWmO7ZKF9215iM5TQiOwhM3+54NWn6V8vx0e2ZbjxTVyg
8fero+UcFOcgMfiWjQ3LhzpUr4K9v/8RyumznTPiXa0ZFgY9i8QPy6Ii5mtpnEYct6msjA2ppCk1
hV3sDmrWt2qM7V0ie8ZvcEg6inkpJOdeEKvE6NXgVeEUCDkppL7IvIZR5LhfxMTv2SP3vC87qI2I
sRFOQNJ01grXiUMs2Zfej+hg1ZhOE3M5Pg9/bI2kvVjH9hzcTlErbVnTDBEgOlOOD65E6ouMhs7K
nx0VymWQ42EMs+2iYuFp8w1eMZE48ZuOTosl+Mkk+N0lUzzCAfMv/URGrcr47oJAawowPyBi3VEJ
ZItTOKaThGw/tCOm56cWEdgNTq5w0T7lIf/tXH8gcwKLJMp+tDwgoFxue0IEXQ8o+yCoi6IHzszA
LTRJVPYDGL39s9N6BdVDTloxWHoBp3Vnak/3eWLUerVauBuqfFCDhmCOp2dJt00hRFFepnqhD90u
Y9KdeXvSdWWdNFwYzyzUwcCmBk/somJL51xBznMVaQUTiqUXNAjLjIGhAm0QPJOfLsEryealIsWw
y4zcbxW01CxP6hJYJHmi5lQ7Ig+t1pz0UY3OJLTt78Q/q686s9i0ASTjNw09BGIQOCE8ALFJ6nU5
CzYFt3t4PxO1e8Vn5gYoyW8oQHTWI2QAXDDCQ+R5+oop+b477YSVP6NfXvF+Mq72VW5kdPgPtmWP
wR+i/awJUVlimFN3E1tspnSiNpSVUiR8/clzdTABa07KBh7hPawWaucqBvIP+YpaOJ39VnpO/vhN
VRQsCqbAdnEa3r6/FDwP8QHwLHEqzbeNmTiqP/kmtuIkIcifcROFjs7gPZY+Wfdf2AtjjRx4Ohg7
cn/45vc0iqu/IQf/w8QJUwku0KGQBmgfVCjHjiOVCS3GnZPrpgYD7TqfRpdm1lhoeK6yr0t/bYaG
ANNGI+5N/D+tD+48unFFITjJUr2GG4MnvxnizwOPr5SAWe5CSumrwCoRDSGf8Z+8FbRUc/a0EdJN
bAiGgV+DGphux6MSeV7WUbuZ9q8uyOgrK/VQM0u9FfRVcvWcvrOKYBOuj+Fx2zdtP2Yfq1CFsnAg
cFRl0KgFxaMXF0JvOPvdE1shBov+0C6oPxkIKzNtMttCv7OgTzwdN4d6Nb0sAMIYmROfE4rd0SN4
qsHrRyZFetrpFQjDMBORVQy581xMaMkCk5oTX+GMaZEehMuNNcrx1Odx5Bj9Dx/m77WI7Vn7XSw1
i49X//ZxSzDhlimQNyx7DwpxJDCFajvgL45CiSLLInmMfOMtzbjsP482y1/dmHgo83fW2yY9z0fx
O774a1ylRPB0umA/JV9JPpmA+cH99ayHrIdUxxQLrn9E7pE1Pb3Odv+174iAYB7AxraUai/3yeTG
aVLoZe3ARLVG0kRWTsXGDK87SYnSACuC3lwX/mMBjw7OKMECOl+yiTKrKQO95X7rukME6U/mT5Cw
tpnf30K2d7XOGb2o1OdbsqA2t7tLY6lsdhmGYdeCRKovQCuY/0HVBeQaqD3Gd5OupGjhC3navavP
sB1U65HII4//6u/AgLTdU4MF/v1vA7c/eAhBo4/UM0B2LcQ1x/XSfoJ1B70VbJ32craBUuCjnPvn
2FhOXjjnqzo2IDKqJ1X9IY5W5BEI2CvnMDf4efUmsR9KqnyomE9VGROs6SiyZE/y5fyCmQolDR1G
9499NHq4p84W1P0E5iiu0YVdBLFkT8bvToEXbQ2N1LrKFJK9NuJmqYcPVxgKUPXv17zD1ErM2myn
fC9TKi5JUtwGL6m3vmDffZARYFck4J/DVWaSFsnJMbPGV9/TBev16eAECaj0AJPynDa/B6Sdwxuq
73a7lActU+9IHFgQ3yWRw7AXe4yx+5fR3D4XwuZL3MApsFfyNK9pc8mjXsXKrazEcFLNqzlyBj7w
BnYs9pt/XSaWPflJMTssfIqRmrijmX8Fb4pu6v+npTbY70RSkXpSwpysFrWI4np4vnJdxuXwMmfU
ArRYNeHU3COr7GPstADGjSik+xKEzHsHIMk0YdvkJN5uJKTcEMkKKlytusWwDjqc8sA2Bo5a5PJa
/NEiuXpVmjpoh+JS9Bzy7poxV5ilAnPVKj35J5YwQ6dwOFOn1+oTB0Fq8ylE4qbN20Y06iQF02HM
91mNxDfoD33Sr7TC4if1a1Auri/qDOTKDGHHi/Vx9KjvqexoJ4ni+cFhMPMxkJCgoZTYx7E/OzbJ
0nFSb8G1nzVGM+m07hm8eEsxqH+9VP38/1Ix15iODl8xzTd5grDK7pcPgZCXH7tTOuKDBR92ZgbS
b/OBSnBDe3ifV1IM6du+3VPt8dyNn6Uph8s9i8/XHniAWu8Gm804DPpBJts/Bo4v1dhgafDsDgPk
nukgJPIkrUnfSdwB6QyHgkRmIfPIGiyTNnrEZpTpAQySLyGICbefnkabUePjWmY/pkmCKNjc0kAc
zXwmHoOr/sHgNLJw3F0Fr48d01Z42J8dkhbW3jJac1RjESe9Fihc9pTQ/L1TH1+ck+/sQOm+s4X0
X2BnI+OJWFspigsMd8012W59lgwyOPTgjLKB7iv7TVtCJ5rZ5EO34PWWyVyBmzUHe1xm6RCrDxGI
UAf2/pav/MlJD+B4hCUhbNEILewG3FmusbeDOZl4NYMCbi+mYO1wyUVhzp2vSmVP1tM7gcU3B5gi
26x/nHrtxvKiZEOG3aOJEzgSmPEwMUXOCyJ331VTQKfuhWTq0CeMgJlhJLnmcwKw6BBabHEqHwfw
eCbB5W9Gmj/cmF0K/MzA++jT4J8t09bj1Ie4wA142gwm7srQBTHicLFZbk2FHQNtomnESDxUX+TZ
WFy5NK6piiJ7VCSkxnG77KUEyparpDH72aDjUDOdm4k6/5q4kHb7KP8j7A3fpNSYS76EmsQckUiu
yek1O2P/oDJUGQorIM/UnTx8Q37LcRMAhDY/GfTajIUlPdwyFR+3oRMDCKSUCDo6YDE064d5Zmsc
wOpJ/iZuJZH+rMf4tph5dSm0I69nzdDnkqKaZx6iylkvrYzpb2yZYP1l9UHB0m/H3W9R3CAt0p1s
Wax6/beqNs05MH3SnfU2yg+qsYKsm0LbOu+3pkdKplQJ/UiWC0Ca19bDzkJzpZ79iDqh/q0osnqc
VN/MyT4XQm0pNDDLSL9Npl0ToLQcfbSsmWo8l7FPmEtxb6D/rKtN0Ne0+uu8eDsvYXP1djNqDDin
fZaHW0su6Bw1ObnuG/g40kvKtESGtWjesQRBnsASzZ0bqvK87ob7EA5RJjrCIpdJlCa3IxqxE21K
/gf9XXds3Sw6ywsvSJYNZFu/6/10uPupR1CzPHEQZFDou4WYsxj5I3Dwjde+xmPm+LF3byxnnk/u
XJ2frv1twb9z2LDFRS2IHnR8m1pBjDpEus4BJOttXfPGxeEMRW2kjBjot9w6O59T+Pk2qKfVqFrj
D995tv79tBh8zur1p/1QV3LVuqKcNHiVcrWAbLuMs8FwjfHslmKIZVFhUOWt2/cEt21jPsNL6By+
sPuN87PH/VCDcF87NHJIFRTs37ZGKEpbs7C2WD6TIe+wW7VDiNuGMAmf8GxcX84H5t8dcdz1Heoz
RrGT5rkGbtMv+KeEqMsWGKuMpSXzIs1zKe2Zo+y1uEERulWgt/bNEMJeQxYn7uD05gPlC9CIKrfT
AVD0ZRNHMkf+/D4ZDiP6/YZtesiHYpQusyZ9K1ZV4ImvnTSX7uF2lX42E9CYu43kXkHit0RsZCRt
iEIU9VscfZEz3RHslWFY3hQh0yvVDVAfX4GTjiUNqyE7N+WLJQNfSUM7SDhMe76NriPbItdslDm4
D3Bn42ySdtjfPtz9RYQvIaJqUGdI4h99Bpt8lxH7VhV0ofZjhc/5AuXvhBfU2mX0Px+YTE5l2Gq3
9KquwHghnYP/CvSiUir25o7shAJZIy3z5LJbg0UbiMac9lCNl8yFQ93fsqiNEj/Aw2S7yPYkp7/9
/PEvCEGNioNdn9xjviLdUYTdFyDOi+A+QiQn1tD0hyBXrSJF6olmyKv0o8coY2HLeTcPLss+p59s
fAd2kCI6YVnb5dDrAW1Lq+fUbcWmQF6S8ErhGNFxtEp21Fa4Jz+oQljXpDk08dgceuryabsNF55z
eiZHqhQWIV59OqZadaZ4CYgSfWd7GfhSwVbAfU5h0vCr9bXfDuNYK4yZ9XG4Ro0R7t/QpqdNDuuI
LQ4z1nXRsuZl/GHXTyk7tP4B5Wv5fQ4cjGe6V5ZDvmhu+GfzgAzwdqOXdVlQfT9Jf1EY7BsUjWmI
Csa2GHssS+YbAhE2TH0XkzpwYHhgH08DU5CnF/yk8XHNkWodpacI3HDyMe0j40tj3rjK7/l77g0i
a7SqElTaDRRsTgkQ6EuYW3iLEEHcYxQfRNWISkgq7Tat2mOWGSI09MSYjm2PveExPz7Rch2E+qf5
oyADQm2XApjrrNAjVAgHKR4r5ZZM34VGWfYRNiHcc7Ee8Rev64OXmjWp36TZwPs4C0zpJOzF2R9/
nZF/OSklAuOTE5vFKCAMEjFPT9c7HGiBoLdRJX+xJ4UGVKNJhu2HX7ltR/XSV9Br/d30aG8zdYfQ
Z5hIcSr67pgRAHSrspGu1YnGFH/g78eh7d3jr8dLaqN8AMoPscoX2Jxq5p9zpte/AVMYChqDnm24
KS2KCTyaaFXHDLt0IZ139MJXegTLdLeLHGt23Nvt5+zpXSnd9GusxOifRSpa80k9tzuCakKXnakZ
VqZLHtOvz3Yt5at7WdO7idfhl2c3WdtbtNJAGCTHVm3hZKaq6l4Vb+nuE/xY1pZoVRVhwsb+3KBh
EmzZUgiRZcOaTBswcQQ5KTWDTe549lpzX3kCSEURQXmSrg+gkOlBqJ5+tECXchLtUkWKAbauOtAy
UMbqX4LJL/Sm/6+g9e0tOTeBQ7dHrDFWNtLZerFjAVEk1Ip8bCNlvEwbCEThLUfMoUV/iS6JdOsi
r94oeUQ6djfauiczW/14vXZ00D5+Z/3C9NSRr9ZiMpEgyU70BV8dGpYG/Xr9jv//6HQVdhzWP7Dz
LX4wfBdjuRR9VvOmEIfJd0kTfYFcYgTpmGIsUuawR1w6o+qEhH+9I+BCjDhDOI75oKAYWr2FRsol
L7vU50Q1oXn3WjCyx7s+5tUSV/ZuieF6jXIA+W9TEXGFIE09hzBtPp6nwqEggJp43Oh74aXzMGmr
lQ8aKP2QqU+1lrYESZfTVJZTGc+U7/VPSayB60eided7rr1AE+RYrsF2lF+CFcjMxgTHFmVzQpdH
vCRgGRXlSEb+zxCI0DitJXM7JJTU0kxjJR/yUoiIrqs07PIMhABo5gL3rQn5MTKm65nu+kQGxhpk
4FUIeu7/18kNp9NN0YVKJ7zsSfH9CckvlvW6AwiJpNlYEmAIEtKWEjjZe5kyDM4hvsGx6MxrVeJE
Gvn3os/PLY3hFf+0adULq3QItKOCkFI7vDkAvrj7ebY3mwlXA6so2FEYVhCznC7eQgf0oZqe/m1b
Jubwa0FVwCg/s7NmOzRKc8mzh2+9yt9vK/0QvKMJ7YBh50iLfwt06ySQhHQZQbItRvdaVemoyBKK
JA7df+VlGCv0Yi+BWF1tqe9jF1nt1cYznE2ShWp2KzmwJDnLMhgZ8Akrl1skNhOZbvWgk1TRETw7
04UbpRRHgMwsHi3sh9Pnr5PNMpuaToWQ6gq4nD3e1E4jc61Ith3wDPr7XzLJfHKC5RRS+yGxubWA
QEQjR1iacEkgTGYS25OQek095IbElV0yFo3r5umtWBwpc84OJ9uvvdCvkIABWn7yRV9EsOa5NiS+
f/sZsY/tQ+eib0gYSLIb0yzaXREPaMw9z9hAiv4EgPkKXBhMF5LGRkIPpcqgpU99u3534H5X6O1Z
MbqRK+hrk46f3f/6X6J/HOHQ007FcHcmH9E1mjTi8OCxMQsweG0oPrfUhTlLjQLmhti4GE+8t1qy
37vfKu4QTflDCWt3Hrh2bpJo64i2Ori9GuZHCSF397TIhNpQPrIxiLs+/l4FakYM967nbPpXnFDk
BIG7cfFEZiqEnDfbcJ6jcYQS9baafIFucvJzPTjdGA5zsc+69LlX6y1W2KAspEDDo0UEMKKuH/D8
KQgXivTtQORkLmsSso/slYbRk5XBr9zWl2K4VfvCdV8LwQAfgDGkMFt1ntZoEQVUVwVkeVGIH89A
07fxaenBnx0Y6cn6Quq/ZacpOqfRyU1g+cgm0ZPm9ArBYJOTujBRxvCpMnapcgh1jk3+BNVnYz6e
D1PZbGRTI4nFgbr4Kn98qbNo5GPymDI21IsJAx0PN3fJO1coOa+wcgXip7Jl8TKz55KZ9+l6eSu+
DjS+RJHpOf0DRE582vZwXS2DD4uRvGT128EAYcPgEBSmhUObtSlRUBaRS6UNgSNnAbz1n1hCaIWg
99Mvc9uiKPEdAnkMro5Qps5lOfhbnbmvvNtUtcQZAA54k37x8q48NGZUCX1nn+pJPHw5j2zbxGfz
kRCOuX4KaulzgyxJgzQI1CZEqC9kAfWsWmAzemLFxjKhmyVD7gLgceNKhTKveu+PiYi2nmUcg7Qd
QVRoRw+3fktn5Vyj6u3oKIlED/7732Izl3c7S7lwaeh2AL3bwnhSwHevR2HwDYdHyAzoxV6BmT9J
s8kXbF52s9sqslsq8EUP5pKe6U67u89DELMETrNRF96xVFx6KmkCC5Xcw0KbVKnHVUI2ScKkaspe
ajDgE0ogZCpowxmB5h+YiNey+HCj/ybrTWU8b8QKmJ2DIIsQ1oMrnHFMjIGuEoEtKvBvXg5yOLOA
rTFNyh43ZmjdGX5j9if0SuKMRjQlyDamJ0jI4EUt0bMBiERbOYPqukE17ms6MDnZdT4S6LNLILiA
f15mgcnO07hZIukJciRy8tpkpmHudIFC2QpH8vb+IZzjEdcE3PdWztfJ36JQ/+VHr3UklGhl1Gio
LM6mCgh/KuL9aCK1eZs3zMD4/t1Qpm1aPmf0rjIRRLfEiYtTst/OjxzQ9yV8rul7heMn1rPJujek
G38xAwXzTd+Yxjdb+RyA1FG/EBBcJR4vvJhT7lSi0Zm5u6SCV95IKffJwZYAGG7WxQpY+HR4doJd
2Gt7r8xW4B/uUevLMoAuOLR14akco6QH5Mmgh3dGyeRlavvORM8UWrj4G5SAlZzz9FJ7MK8Z7dbR
KW1CfGEz0/j9NnBL5z+gl+RDxVVERzC4DLcwMFaM6OJafeT+FFY3ufsoel7ZHas29hHuBUj/at6u
wzc0X7sTWdlJZT8cpaH5Awtnng4P8Hu86rZupBZ+5qV5GFCP7eSBOtPzqp4bGXhSIjmCpSpha0wd
9m+dNzOIuYthDmX+8cCi3dJIxq2DrqOhOmPofrU1fYmCGmn4mKi9UX0mJWWLHIhAo+afFtqCXNd7
99y/j+VP/8ich4Ocqvrh3884bZ9z8H9UWMvCTCUXGFQsnXHdesXSO1lbnWYAo10HI3JuiQxbiozM
RRtzq7GYpvyb9HxuGMAdAGVEINWO+wmo2rh9nb2j9e25E2cA7/xhP3qkwspYswPShnQNQHQlS6pL
vYEFBEwbs85rLztepB7Qfm4twb/xP3UnO1kWcLP4ZySclCjse4Rjr7afr4JMQxqkz/6092LNF+pu
mYd3v7HB214XK96n+PvB8yU/cKosWrf+L1YmC1/WYjwhTbwHHOIK82qGSeHOw1wILLEHVd+vOQuh
cYcNiJvPGuR+yUiIh60v1IsHkD7XxCDpq+57BzVgEZKaLgJ/xkx9YCVVoXITki7IVA+BiIIEfVXw
iQhDCWZlA/g3qyuI5tBawZhOqTF4Oi8ZgetnxUX4x42LjNKdmqb6eTUIVlN8dxWgx4omuivKzjsF
8ETxttsFIyrlKmZw3iiOVa2hhsMdqZxnn3/m9JxHgKOl8bsR2AxnZeSl4RGkTfvPIgmtP4qjTgND
/MmTu2H5+pAls+LzqeN+vMOH3Gq1zFaGJ4Y5M1sXIzdk4iLPjAgyD+NxvHc/RUum9k2mTUMFkbn9
z7v6KL7ePmX9xC8Nvs/Wz1JN/qOAms+jkWd3aCPSezHDAdOvIw0OvrWNLX7DTnkzs+KUqSvCZF98
0NQ58w0GsxgBZ7xOBZ7FroTf57fe8iTEusrR4bZzSpT8Lwj0jj1i++Tv5EmVV2QnEB01A2HSOsfu
YZcVo5nsYmv3Uy9ze6IyvPzigyuqjvqZEvKPdmL7iJ0pRqUgfciCX8YMMKL/yCNOKmTKGuj4xQ+e
lpdppfApEBss+MX/LajluCDXGN+v0Bo22H2OStH++18Whsw4wgVB3faOoHRTg+9EBJihQjLnEwx7
622ggnI9lYnwCwaTUGsTHYIL9z1V63WuK5sytTTghlUj8NYY2pUDzpwrlIRz/g3aVCLiDa6Hb70M
BC4xttGMDmoMzS61ncSlBaBc0+6wMarzFb9zbUgqflfkepfE9k9odQYmcNhyJwitmgtR3GUZrYjt
4W0vLSmed0gZbxQSBa1kbT73e6kIlNeEWTl1td/yV4ip8uy+0XD+9ZOIpJF7sONbq6iSfVUQi81K
CL7oug5hsB3u88790Bh2D19rl1Kry7V+REHemwnXqb0/txZbcBqnCtrCHq66GI2prJe6oUsjwkQx
Ip1daHqANmpQpU4ezv/D+ASQOYLFDRfFQyZKamcTdK9/6ry0tgECiMpuR98u6NC2tQ0PFekysOvd
8eB+lsX0gbhoRh6GvrbkBxDgCumzDtV2bBwVoVZja8RuDh/MucdbcGTtrQZRarQi94oeNQeYB1US
iEaZUDFQlGByYZ4q8KYbCocRdwx4ze6ByPN9MEll7lBlMm4/mCJdPuzLwLv6iJSIDatHLZ35tsJN
CqcMxOcA7JJZGj7n3AmYpUKnGSwPGPKMm+egondJebmpsOIECC14IL++81DuOWZrNL9br/YlXutC
eSrkKiToWXarTLYweFOLzTYfmxubH+cJQuMsvIoljPvNh2bhHy9h7eThA96UVbttePWI3Tz3Y+cA
0KY0x5D028Bjd9q3S2Y74Ruwwyq9qga4/XUAMNUj8M7bMjd2DQ3xP3jXMMRoBPoPh3rBQixyI1b+
ThiLldwJnIn69HVP1uRpQs4BoBtUcxRc49OzGr09m2tbq+6CnZl0fO7XfTDNys3W1ZITjrwsvN3s
TrdQij5uhzQbDI1AzRAI67QKUt3PBmZ9/ldzjERzEI1sQ6iNE8W41QXy2N46+E3ARpceQZt+y5vt
voj5pWc4T9Hf9jtPRtxHX6BkghCQRpv8rgS1XdT86cFHyxeagVbx62KSRGrkd/rB370NxMhCOh8M
ABazkZbMqxwyhWRjyj2VvMhBTtskdAEoNMOKXafVU323gmvGsVioi7S9Mg8PI+5iAmxnBa4hdUag
EtHyBQn7lxzUT/bSwviWJmAkvRsuBiUDbojjkky6JfJropJAeXa1tuXYu3fqezs4fMX1kKx+wDIX
Q5p9elEYRS1Jck35Y5DwHgn6Gkm2weaLtS2vpRL0K50yiwWBaUSa58VbQXnTJvTnWJx2FgrJFVjg
eqRyvefSiC0OJYHJjjhYAVaXkcPa8PiXZcRVLAOt/EwK2ZL7ykK/vHz+4uMVPHp/2kE5GonTqv1R
8XG3pKiT+6QlPbVaf+XMDoiQE4DofSVe1dFDhxZgirNe9kj1Ckl4xyI3FAJaleHkq4PBsVkeNhZe
wuMcbPnV53crrPiukj6zGIPDcZ0sWZpb81KpVwtjdh5oZyc7SmauOaV5AaRs1gC97kXen2gF2B9U
8w0kHciMlLVtPY0P1+sHFEmgDsBLkOKi4D/PtwC7/58DpTQ5XTjoCVP5dADQLCV6f0DRC1n/Hf4U
CJsNRkhgUr30v9ioGIbueVvlR3yGfbtqTplZ7xbJ+TBkEEhRgdEXR9F0GWoMx6WqcVeaSUuvaGX9
sJlZr8nzo/AuUQqYxexYo+22vp0gIYzQLQ2MQTEP/xXILyTNWR6wOUVPWEBIgWr3HBjkC+a6gfM7
KL7iC8j3b7Y75Dnkgp+Emt/2s1txV0BO2wn/ExYcmzX5UydcuXzWJoP9hLekxF3lX9lU6YiMklDM
HX//NT2nHOdc8VlM9C0xlU7zLAFtyJXcNxS23oDPZLO8h7NPGHtkPyBsI8hDVzLnNBAA1Wt6IbSJ
N72tFdO0GBF8W9K6JG4l9nif1Bgux32KqP8uvHSGnu+SkA8FMs/yTi55MQeTcJZB54xfR6oRtUQB
GN2kkMjFCIMaI4gsdj8wHgBmIEzeM/+92sr9ZU2bC5MwBpLyb5rN2wZTiyJJEDRs9vdJYUhHeMSa
nj2Vfx8X/iX+8GLVv+nqATIHo4B/JbNphX9kbNDWqpTlaj68ArfZP/ov1hx5Wfsczn2A9MMr1slP
ykQyhw/LaBoZDF2SDQnCg3fbQgyXLG1WKsC/6+SGxU1v4Gi0727wMIeao2Zf5aHF0ur8fg+Ul5Y9
C2tC6sbDjspYQf99axU6/N6FesQzlsTjr9AHqpOeRMGMhUzk6ZiMFfpH6iQYYYdfVwmOs52/N+4s
hzLMJSdIS6wu1RYVl66wXoIv/Btkk/4TSbJYn1B2K2ZgGyI8fJGdsRAoc7MydmugSC/vD9DXGhhn
wanLuth/HCjZPUKWdmJ4u8ZzhQf8Z8U2DX4F3Lr9HvLteIKt3C2psUFGZlR1sqG0A9KVYpQn64oJ
HmMpUgnXHIcWyDhPerhd9SWVPLmvVIPEimdU1nocV/OWmAcOr8etD8QyLJzNHEFqABE0baTQstJJ
PB2QSqUUHcTgto7BibJNEedN7aXYPeMaobmDtG6eOrn3tuuTSrLIu+okfcz1SZISwAVsGh+JFZUg
8iOzAgEr5Pkx/vYstXrcjU43eb6BvIOMZkDgQJ4LJ9BmtEJmcZk/fckNwRG3dH1i22azCoTaj9tQ
wvjC3s0ZB4JbMillf/kYoTNOO5Ba3eybc9LSTj+ClOcUxKxQb8wq5Kd+N2UAzZ8gmFmuXzipZTy/
q7x0JfpIKvYeM6UuOmDgNoFmvFJtwVBNjn+jyQCJrcKpijf1lW2ipxs2g6ra3bvhmgooX5pgvmbw
0xxdTjzh/2otVHti2WbAt1jbnwd/sc7l7C4iDGLDqcRg3Z3H3kGSYc0dDrF/b0CqVW5yl7OrKm+I
vB0dFfb99KLlDLVnkDKv+8yDdmHSqXf6kzvG5oRqQn00HP9lyjpdlFIo4sIeYoKy34NNiI9JDOLX
bY2V6YtvPeiactURU5CnOvZziuK5bnJiLLkvIM/8nDG+FI9I2ErydDZhoS4R9/H+GJ/7x/J8luSP
kKlCb3rHZe/izxPL7HVjK2VEMpib59456NRteMvJgeVljj5PVn2dxpc2cyVOX4nzmB4g2NMT9fRG
1LLBWAklZUfekoIVfvM05u9lIofY/WmlRbXPCoF0FvoQFCL9HCODy5V0wx3bDixeY/yzL0jUi/ds
AjZv4N2MQVu4uABulmVYqX0p4eu0DTGyRV8aiLr9cBvQtCaIQ8wh/m6vmfipphpBHq1XJ0iSaTjP
KX5YKyvHIVLhP+AhMpGMJzDMtFjQ6rPDFxkwl03B8qqvH9T30HHf+Vg/QEfRXhJMSLNnLbSCDC7u
nhPH7rbK6+ZWHbolxq+zcQpviTgAAq1nhYuBjOVfQ2zH7qNHVFZPcCy0/mnhsKfwb167oqVfByl1
ewOXHIjPmwoFxPOXtcuDAf8c8Vbx0P0F/snbqCzqJntitaCEpLeb3CDHpUX7otctC3weAShVpGVb
Y7MSq1lbK0ZCjMvYgK980ZVYh5jkdBlkK/G/wYrSXhiOeGCXl/GwtKLx/68GRChLH5S6tiMrdy/V
GcWpF727pVHIo13MDBCY1i4gxDuLoNz+bCPFsqBqv7Qx2vlrcysaa0D1qSdbmplyCv+ET9FUHFD/
OzhEa7CuGpmW43B94lKVE8ftikfm+/ziIF12OpukRiwmK0A5yVKb/g3bZrcCcWmoDjw3vCLQj8O+
tjxAAClN94xUefywkHr/cFMmMsknMr+TTgybrkO33G8ef6F7jITSDhNfg5SJyuMNoZuQd7Z1P5Kq
CxE9eJ/hwRmeHYIvyU7P0yDUcFOzLdjyWQETR0BNBBlHcxUZOwbElX6y+yBe34P5f8eKTynqcj/j
HB9U1zK6MwtTbyqpmK2xBIBCvh8M8NGiNMgKNc6XKtsgA5w/fzIoAbce+jyglITJgqDoDURcm6kD
r6FMs8ZDi75ikSc/SeQCSQwihxiCiOKNQp5myqOm39En6vHP5CbTrByAKnIx9EZ0wYU/nAGaA+VC
hA0/yNgL90uIrj7RHw7yIOSyvo9DUk/4nTzcZwxUmGJlwxV2o965+bcAbl58jq1Es0n1lUXq2V1h
IQVtZob0khx+HM40v2JeD+cSa0OR9Wt+qXI98ROhdH/0XMgVN0mpXd/U7hHA4hWQtt/p7Cn0CXG+
fbjg5quct8bXuxbgayO3/LS3TzxkQoXaaXUXZGR5Z1u/au+IkKfLQmMVYfonbsFVN8ketpSe6LZ8
bVn+EF+UDDXeMONq9I9vAaHUdDxgdifJR8FJpKoAXfURzT0ZFpeSxlnkltKk+ydkhngH0gGk11Vh
gNNHe3dPeY6XTDmiRc7jsxiSnt3MwEX9zPS1G9Y0t/7QArkGpxaxTKub6HDZ0JM/8sX9XJeOMfcT
/5DuAJs+5pKzDoJQRQnYi/fRsbWXYPpqu7i2dVIO0TIRmYZVMKaOb3FtwMY9uUu/RWvSAnDeLhko
8L86Oymr1cyoY8kp2Lli8dzlFHk66qDAVQs5cBVnZtZZkFnGZY9YfsQG+uNMmTjzFZP0dENzsZa3
JsgwbBRpZHhWVrKknzkgJHKclHpj2Bw4bSf+AXce/2p6+a5QgWOhcXXMKbbFxpt8s54Ki6xAOv8k
37o1x7WyjnPmtmmDXzNvxTWTSh8rgnuXujdt8OGBR5jEjmOG7gFpr/mPEYlPQFwX1BvW4rg4I9AI
ttNxVmel0vl+5HX/EGaUvYa71sRxfpG/Nr90SNQhoc20WURFCxH2F+EeCZY5iZVg9Yx44dkqz12k
WY1BifXikZJLbVZ9aSw5BU4HSpexNXKXjseVfePu4TfEgJ8UU/GWuaPAEna3SZ+2DU8OVP2do9Q7
Xl40dvqWDaP+kCZFkdMllmn040EboBdGSQL8KnSMkbAQAT9/T8nxjxU6DlKk4QmAUNOtdlklAzpM
riSMI7NjGW0ddPRCyL4ZIBmxcE8vsJmJS4nDez5DyNlXGGhhu7bXTBFHrGZ0Vswm7so1agKoY1Wj
0UyRfZtNb8z/4mOOMVo/yyO6zqP/q3nigSDZDiu2r47nvyWE7+AyJzHmn5sJuuHw91wNxoxJUFP8
QdM3frJ2jVgf0e/q7amEDhqAWeDJ2Y1oa0vWmTPRj1eWg+irOLUz5o0zPFQtJsFILBUZCG7cvj6r
1DCBtqPe1pIat712pW/YNDfPbXFuSipGXgXTmMIzTiEOxjssCnZ5p5IPvBodz2vB7T/M2x4PUiWk
jargm0oH+YkbJm3/+1q/nwiNQPU4PSsYBJCTiFdfiUKPRGwcOchi9eQHOBlssrhKNCRpMTrVF2cG
ciHUK/lHGHSUjuqFBGiPDaeEsXngxGimwuJY3mSTAcUJvxoeA3MXlxZ+RDStBM30MVL8KVOaLrS8
Oq0Cdvr2trGS3mtNaWXzCnOrEnGwwgFfuLVMiWd5IFHmv49c25KNJsfo42peCgvufwnMrjrwfnUC
4+qpnWvvC9GUt0wiYyGMRlHjA3FqM0o5zhUn9Ft2pYTBbPzj47ClsyNyT3JcH9tyYlj3SXhbM6TP
wvfh0Azx1Ht/BMrMx8YrlYTjtGGafzJb5ypME3MEuAYdlS4f4Ct7KR5Gx+pGerKApNP249igaGcz
0CgXr1T99agXun44RaT0KT7o/1x+REZdLDmISurmpXwBmj361l4KAK15kSXB/WMRg8auKwv69Vuu
VdlNyUAgvxY4bIO3PdN/+ksvN8BUzPTjk4K7sctP+VCpnGomz33ngDVZyrsozYzeAuX7QzTaySnh
1bNKFASaXlxf2N8FMOqEwcooh5avD48tOOyu+5QqRRUnussPLCbuFPA8UXmYsgTS4si9H5ipr6qe
q7774B2xl853pvYy9yg1H86P7az6Z7Yw4XRamj2g3cHnxHCesZXlpFAlRqgFforsSiCZOqIRNeB4
d32fuxHKlyghxpGPVP/cdfxjFRsHy0MAYQKNTqXXQJWN0HT5VDEbJtlEKi63+gTs0NRA3wM8yPOY
Rx/LC5z06ggIQ9EPrdTjlcSIGD3OGSEMGM5DNqFciYTxM99emXrJy593JBS8D14DlSsYyNELd2od
4iiLe0qKKnDE+t/zCTmcgTgRO23naJeP/Jd1nsd7Nc7LVv+rkbQsLaU0xV0mIUJ1FKGHBKD3AnZT
vVCgZrPFf+tPH7ZbpDIIsah4ylq+VAhwAkrH0KzhWDeYJ7BBZ/POxakYIegj4xVpWP4HuwEFtn16
HJrsgWuY40jh57DIwUcE+1rtM6EGIPBKHJ2c8IvZSClFZhvdosqJ9nIZYRq4B1kVJoUu6CbOGfhF
VS1KhEcOLd3jlahKn2X4mEkB4Q9fhAfYB/uoMjboR0X4Lq/evK8egb2DjepAF8oQi8vq/rxzjBEt
lVAvVr4u9eFFW0AkPqp4KgwZWDssEECapquI7latY1kb4SrDrredn5Fe7Ni6sbUUjkGcb+rM1WIU
QCO+OEw+xWl974RwsUvlKhvdLM8+pffpvwxlrhYOX4LvFkF7r6+r7oJMelExjMQKt28UyRL1Pttc
YaRGo0zCcQ+LhuxTIKt22vrLJ+Lsjbnyq1Ipize4RjitNmh5yEqap1tMppYDRaF/3wGHd42awIZ1
ozh48qlXrSWXoLiBIodEHj41UusxC2AXa4dD8Jk0N/B7PNg5b1v6jYReVSm9zZcaT58Q+tV7bvmi
d4jZkT/w9TpUwa4wFaKv5G2EzmZMiyLiLZsd3T+K1WNWK61NCpizUqOeuFm3aqEMBLsUpuGMxkf+
5uATCCrmOW/dSnSFFvMNxvBeLUy5XOpch0+cLK6VxgzCQOOwGx8X5IxiQ1jO1x6AEofFI/ZaN6SW
JG3uKSVRkzfvp5+IYrWTu1k2irZjY9/KxtqN5Ek35kxknezH1kbqQDlfZ8LnWNk4ABVrELLg0Frg
Kb+XDKFhoUGzLUmtbJUjlpIqGRvH8fRpSdIK/19GUiBJ6/MEjNNiGfOf7hwM2T3/m2MZJTra9Y8U
p4kK0lm7+UJ3BZEx6vC8LAVFqMZ7R0yy4hLUG45In5B272KEcbqhlU6QxOCIoXLPEqRZ6js7tDrV
FMiYV3jgFHeyjvaK8mDG7Tm7/GCdRti8DIAcbewolx2L3tLKoRrvW1QRmApYxt00Q12iWnbYqKR9
2KjqoM7ZYZzSDiJEGfkf6vHoWOvSYhXytKZcl/JAO2ctGa1SF8uU3ZuWPlJCIWWa2rYOUMwkYmF+
GN/W+ZIiRVPdwLvqMuNnC/Vebj3eiGTyB85MR1G5jGj+M2Xv68Fg0mMPJRYJ8N82oJPMpZHEtsZJ
VQ5H0/NQzeZVYVTP6UY35IbHY4w2q0jiRdmdvmHp3sKYdv1Hiytf531KUsZ9MzsXNQSD+hxLAH0x
DlXg9cIIFNXSPCw9hdE1szDt3FeM4irc9uWniiXAioJOTxf39HW56LPq6gnhoKMPaVM49b1PsGkX
HaSeKKnVLXgaiMC1DUaVUKn2EVDv5cefXz97pTfiaUkt47lSFWo8OFVKWQVEu604Pyv5vrR14BnE
dtixlmbZcWtVsp7UQvtMJjW8czVRHUCVCFcWRf6PA9ymco1V8mKvHLtXr7FVQ7sCWFv9amElEMFq
6UYgrrUl2wpS5y2IC8TQa8SF5ztErgsd981fyF8ddBs47FIqfB2lXJuWKn8CC8llNCSdUxuzd9GK
t3cGzqM0bGk/ZLJbMtmUwEPKmF6cD0qFKnCOlXkHt4T/dMJVHg0ZFsXQq/VOpqa86a3304ZPp+92
G2xYwT9Urw9d0mgvghylqZzFGPGImTyxz63AQI81UR9nNPueTwMupuXIWio+5o1nHphmrNInWr38
Pj91fUruBPEZzRQMfnrxXY/gBD4yJSHNIkffTDOZ3upUuyXLIezjMpBk3ujZ8D5kIFXABrQcSeah
sKa7piUEFY2x0SSVIiC+cG9dxtJFkMdV22euQRhqc8Q/4/RnFVPTn8r//pUIliQq3JiBgjQIyDfn
ftYzkOaZcJGdvMP2hNmps47mDPuM+kninz6rH3/IIUnyajUOXXp4cz7o89cLatzIFhzYvcHPJ0hh
G1C6VUT+EgG01vWkPu1DLix9FXaN5UJqPby22Q3AalM3+lq8PLvMNVPOM+jcNl1+1atsua/g3XSd
1DiOYlA/Lryz+dzuRh4Amn6RCz2DFISla2tl0/Vq2WfOplOZEjRaMwzxa1oISlZCTfoYEmjPi5hf
jF+w8nQxsiS9Br2ihLD/z+2sviboGtg/FiO9HYFWd7aGo2q0w5rFZjWdJC9+yWiiW1V1V/pB9jaT
J3JmV5Haz3S9VI3oRKMzoObvTIFla6xKBTW2AEVP3V3sOV381y9eEOOp2TeDlEt4ZDInfekPtoJg
7dXCX7eZ9ZZbxOBfL/8tUQfnXB1nfj4bwOgtzJi/nHfi2MPgNg0dRAkQz6EGp5BkntScjGMjaL/i
4JL4DVCJzbQYbsAG7jn5B4VVT7cTV3zhb2wzGdnMxR1rb2zwkwVfrKTbLpdHUS/xOc/w1s54uApT
5gKlKdduYdSJgP3Pm8Xf7WMnegMtPMM3bc0o0l7YPEmYN32QvvYzouBet+Tb9V0Vspg5CXFIyGpc
XJLyDTuTE0euxsoJPos5UD9cyW8z3FG8Ac7O/sZ22pkNt8nL90Ct4Kp9YIsglcSbB7H2x5ebX5E8
HBKZzCrRU7Ys5QXjsYxCuR3kVF8ciZqvlLcqcZyR4DfFvEGm1syssjG5BEBIVQgoo1pX4O7DS1Sm
hnlgV4H7WBpuyOvZm8LcQGxfiBQpeSymWfIJyev/fzwb2xG1Usvg5xQ9uz8vKlg/CBZUVjXK3hhk
+40CsrqztsGn1U1LPew87yulrhr+Gp3zPSgIOG9iCVL9ssaXN7soZhPyp5MvMIQ4RXqyp4ByeIUW
bOAdogSSlwFP31e9Q6vxYZczSWzKvyK1y6y0secvaUQAQ+ehvBk63acmXwalToC983Aq4Fn0bmEz
rhnq2YTg6cvaaqcl0p/F5VqBYwrjSNqiojIL/q9QKgZtGCrA04t0TjGmqukAMeUDicBz6tyR/VEo
VhZES7TsuabXyAp39UqaBePljl0I56UV4k1+5n9LI+ew4ade/IKUON7Gz71g+RyPzDPhtRcjix+g
lz6zt9hwi760EWptKm3+0TWh0Lc9CkwpOkYINDYS/el/NtoXWSsiPrsp3OneQ82nUe7PxrI69Gjj
g/q5C03GCiltwMg54mbNYCdCJs/R7RYTy0USOowr0vYQ1mLbk0pnY3pcjYtn7E0/dpfGUXBYjb77
E38Khu5SVmFswNwPiVnhsmBNr+yCOxu1ZMe3H0uZ4R0a9/2vF83K2pKPiK830ymoPN0Tphp509bw
Rrajzoi0N432l7DuNuloHWbpSpupZ2KsDje/SoLCiBdfYCHF96SdbcFpO+sVEzjz3NotsAAi05HQ
XtEcSZOvqn4iDFHl+rTzkAPH/mQxBgy8Fy/OZnm3iPGfSidKN0TA/Ah4oP2RZTPGfAKJ16UxpOUu
sWUVyYJ7y3igMO70AVAwVF0uy9i074yHO3Qocz/s9PCxUrXOaveHwVuu/zBXd+Lp3ck/DH51m+g+
JXDouPq+a2WVscQAg6V0n3XI8qVCanK4hGSSiovYJDZrBGZbFkqe31eibiyF2p6zLkZPC++rmlma
2DYbcjk1Lsx7idnAtCtKN7Gh2FhObI+fgjYSOYRenRJDvU+9mdkFD66igGUfAOIaZtBP1PC/MLft
pw3C1MebsnpB79RXaL9DFIT1ouXHAL7atSBdZ71YHSnSvTUzshLq+c1tTCgM8s8AI60WJAmGjq2V
yQ2TF6HiH7SAgIF4kD3vzks1O3ViFvAZM88xNF2YZTlftekOUdAbXrb+9AGxTvJkg0K9v4i+QToH
gxx1rxwqiFmE1HBCHz2In9dl5hjExWYOjlfnD2x/3TPjxnNPSQYXjJdFIUaEaAsGDfrKs1Jq0zbQ
oBQBAnme5lkGp4oAk/dXBXcE+gbuAQiIx4yIDwt/cDL9Dsl+T33R/sRBdnabPkwwBfZP6T1BqJlh
xLtNC7Wb4ynRJnksClzhVM/+3bi0Cr00Yz8cMgbA2O0uV2utWAAnC0YtyyO3l2ukyts6rKGvxrWj
6uSyO95si62HEF0Rn1grObixnw0fA7ilunUxr1r91Aya/WNIp71HqL+HSb/kNHKDNJ2q8YVTuWjd
9gCBGRVCZoRqI+DdSC+ldicKR7jLwYhHhG/mzFspaOge6OdRzM1VcAdmDfgG37S4yuLSSnIL0ig9
7zKTNzo1JffJQg7Y9O3xmdOKexgprykxNTJN29i17DrPjrU6yJ8huRwWrJVeSj03VX6lwrAYB9AL
s4Bf2HqtkDzU70N/Wvj7JJutUgeOToBsoopyTr2eBvvymUVqr/3o2yW0R7Bs533sgZegCi1APXLF
kefMqf7jTaI2mue4rchmFxn4u6KrqF2x2On8zhh4x15+Tf7LjYfKoPIFb5OPkoDXSCVfWgubUF2q
6f0pG+3cekUAozrqCzodx3Q+6IJZd/Hn5dOBUoaKteZTvILXAbWnfJu+DAivA3z/8nKbptSFMLjE
k0M8Pf8t8aZqEcRQVGnTlRT4HH1ll1/8n27pG3TboHLlwBukmBBxOFlID5tYaouBOM6YaG98PDTU
lmKC1PaFrVd89TZT2yWRo9cIYKLR937gPadeWFFYHkZ23rRaY7bNXCNPfVlDomZihQ8Czymq456M
JHLcXwb2teYB4P4U8apMF0kwvRmU4YaHm9REjeFGceuq2J5MCkxopiPD9J/gkOgEcXkmCs4T/v0W
rxedyL6Bymm4mbI5ydxkOsH6MyrZy8O9HQC6nYHMmPi++kTK7+Xc/b69CLYfgcYVf6YjOEW0fog8
hauKSqmiVF4U2L/VA7lqSPChCrMZ7pMBf3PqHD6ymlOC0vOfDPjwbXKvqTQSk+fO/1UJeEl8hiw/
pdNWTm2R6krwim+4B9e4BNq6scx5loLsMGT8ljx4Je9uTxmsVqUpQ/G3yb80LA+2uIfZ4DKmb4x0
Bvpo9RXYUKaaYGUxWJBQDk/WpemP5hVIYQ8AyLaaocy4cHLb0HCE5Amhtf1cXe7/iLHVdoZOWovN
xUqMt49WBagmNsSr/sV1eJUhVEQ4KFCb0eg9DDsVn6HuPMK2lXo9EvD8NQ/rBM40Oe3xo8/5v3Rj
hO5WWdoJeZ+niZHrpAkUqzNrAxwOvbu/qAQCNWSJbmbez7iDCfWa2hNZzeT6UDDKQgerLEMva6cv
4dF7x9XKwJ+In8xKmzuVvIzlKdf2OUWIKDwvRQNMDoxvS18zpSrjfcTJTkMuo2tAWHSLmcfy3iFV
DGwYaQWIf5P2+yaqsFqTdjkCHaPTYbxixWHvWgDLyHkxUQAXP15vJuMCSrdIGcGkSBRIDF4xBr/P
5xYAtpgWM3sVYcPXW0MBllFNth2EMhJ2xzOI7GczR96L53QS91Hl3Mbu6eDyuX/KfxKvo90cJYoN
xtyZheO0ZWtJm08N8bKcWolq1DuUFmfHO+fS0ZTY3f/OG6EzPffzZRmOuPE7Xc8SSulI8PKuhw81
hBeW0dKrOzwAAMdbOcid976FWGLZy3pqp7B8HcIPdWJzbiZFeXLWxebWAzm74X3FhQTJVZuO4tu/
lX9gN41iulK93Zq3GmMf+V9NL9Gi953u3K4wK7TgASR7DfqTzDKi3t9QL0cikuucYqZVTbMPjzKY
AEzxAyAlnWlmVlLG5mtxU51CzkL6E0jXd8PPAXM56mbU0aJEJGGvlZlJ1nrDUF+4W8Y3fp/XEplB
Us/PEnUNhRJ8ubKheG+tJfPv8nvOxGxstPG2x/sd4Dzgg72GzeE4tVzZ2DNSrFl5OgwgI7+/DKf8
hcRVcIZLs5QVGoUD9GNxmNnglL5M1QblnqFQAEXlT6qxyHo7lUhonqGmOlmjcScaQl9G1OISWc+k
ggy/SiAbGoseMFog8AebXtbexnhMA3v4YBhL9h2JMgSYTfxOQd5DE++An5k2DdqK1FPiMjrooFLP
OwZhGP4xay0CtHZvva65qOAh0QsvnFXslmAuVdMQLJkZTJI7/rGmgTGQeJg+QyJJyx0WswbicCAT
q92x3ulmnI/Huh2Q4EzJ2D3H/tZvlxmaVX5Mypv82PGpUUV7wggQjpLJTWtUX304uupdAZjrbHB7
5NRM/EOxGxkerwpGUBCQLphnl+qsD/xb7UnFx3hyz89KJekw0RQJcY/a4CuKBry1qvMbQLI1TvuK
HV0OFEIQ+K0uEkmtCsqZ+n0vZlV30Y6L319O0VSyfHzA9O7zkqqbHJhjx+86bHFtYlu5LCLCSmXv
tv1RAUPDFCscfVXCCV+sZba91Z3JlcGkNiSJfwASg2lUEZsIRcpRBoQqYKFskXuoAglvUNzCN6KC
MaABahA4pENiPVY1noBuMXrBVd/3NnvRut0CLrs+EkJeSpDA0Zk2c2SWWPMQMHXmEsplAwmwPEh7
vejfP20nv9M9MjLacR9Upfg4DQQTtsnVMHmVhpLW4LSvz0Tfcs0QJxQvpuUd+u9W6FppITAWDHGl
AzRw1WwTMsKXHdYN6YazD4kECV5YEhSDP+Oc70qMzJNTZM5SsuF/k/MqqyUfG3VR5YLPaqwJ/hQV
fxEQ4GyJBSbolz2u4OhU7s1eonQ9J1N3wgjdL71qRKsrtxHcM/1Z952gSzAko9V1K8/9b8VHXbrH
x4A/oSkU6xS93P5RDFqsUdHOf31HLbiKAIMHIa4HoWMyAGjQzMJ3ABqglqSR/RGKRyqcDFrPfJnC
0fHW3Bu5mieNbAUJjddJ6odWp+N0HnPxRqyVrv1XTHBac47BODCTpveOxQDa3hsZdNz6jgXXobya
nQm/kfA8J0ROd9Epdv8JxfvvyazOw9piXKfMIBQBNRvn8moAubw5It22ubjdfGJZ7X9IzqBHeddA
eSVSCtx4pX8H2a/ejSb7Zn1HyNiFZZQ4BaBbm0Ex8QQ/ZhFPYWNtvbThsHmsQWANid+g+ID9bm7C
75k4T7N4STJ+ju87kKlu8TfZWHm1cRI+gm4AWWQzLPKJjKY4GHtoTvDT6qGPWJrprHuFltBaKH+D
cXGd90yfpy7m3KqZBm6SsWD5B/8Uz0eoPcVtR6ES2QAYiTMzcOFjkG6Reuxj6JGDbf8EEIBLVjuO
/RrWJA/6v8zNhsN5flUobKQp7wEl4Vi2yEeBQbQANTwL0/qPc4otpWhskJ3JFkYhx//YEMi7XHfa
YnAkuq9S7e8fU8iXxm6JQX5Urc3PjVsmx5sJ6VrwYIfR7/u0eolGxcg6+QI3UDrYZUG4jsMYFZ6i
QoIYl9k1bPnw5DaRQ3Rt284cqFulJC1QHQ6C17ZXe4G/deZaw/asBwa+DHPEnE7J/3LqgkLX1JbH
LHpm98g3splrv2Dvf3O2bCBUl6ufbIb2EdEj0w0L+cu8BTXx4oLHmVCTbn+FT/kwMyvjkP5ai1GG
kYcoYzdRDdtI26r8krSPEUQBLCckt9KYbzAV2BPByf7oKTOlgnZa3Y9ALL9CxXGkLJKCNoKRO11c
Zw7ttTqq8WbHVsWWD31tqqYC96M73QjfY1wWnGjE6P7SMEzxSJmUBqacGjeWLicdLiP3atC489yj
4SZm9KCDztcpQuWp5FeNYFPj1ngyv0sPLCO3fw7CuKzSo57aGps9oBSnJOyt5vRYbaqsZ6kFP4uQ
qrvoh+v1JqxnE42KbSi66oNtNdEzzO2LgkrU1ACeQlW8YuP9DbJuJj5si2jcF+E4Q0OWfHVBm1MB
3MaRaddgzPnTLqR7ZVUcoxxiJfSqFadzPE6dEAvo6EhWbO5mwxptvqxJJ8Jupt4RN53O0Vb02J6K
IjfYsxFhKc+lJnpY61Pyh8CpvchA+iqzekHtSkd06udpMCLxa5QHig6BU8kDOanhQz7LJZqZmBiZ
dhgrOKBZZov2TD1qN9HYhMyFWw1veLUaT1QP/ZnLeZ/ESp8bjRc2ukebDeU5cJKrINqHgBo3q0qh
JdEanuImuVfVmFcLG7PBhwojADEXy8LcUzcPcBOXesGskP0nX77DP7OO0iXP9VZrNdoE1S/jvqOS
rrRzzaICo9Q6Pg9JfQD6Ymu7a2oYjTPkRwfLQ8J2lHuu23DwbjJ8BL4DlAS1pozwylceeYCfa2/G
4B4sQO3xYSx7JSaeAgjEjUyYHXvgbti5N2GQmz79Mu7UutYxFTkxD8cue/63fHUbYACokZEDzBZp
KIdCRX6bMtx5Wrm/V8baA8pbEy32d+7qcYn47RsAaOs17AmWDz4wO2HWWQ0N0Kk54V4guXl4nuU2
Vd7s5psT32RW56c59wKnnQG1HtJ8nU7aS69mD62pz1WlDz0oNalBtnH7MTeeXG/d+B47ZCZqPP1i
vmlE/FfseZ0dbvO+HTqqy7p0frn9zdCPHeTVf8Ogzqbg19pd2xNqhSMge3AqSR9rLCXAAn0rclxP
HtmFNDdTpZ+FihT7A9zQbrBnbqGdw1UhGWPiypZyR17p+AZl65jlWCAAqOSg2RIWa5MlJfkPOUgj
dff+xcUvH3KXTO2sNhREp8DPJqTKBa0tfkS2PIGteS6Y+3S03JWj4alK6qHrFeqD+hcu7v1UOSJK
OrPNcs1Eb+6QmA7C1KeE84eQDd4veYw7k3jIzQXNcZOEfd7jS2TnxoXHa+HXHzuPIO9iBHPjpZc+
PiMOT7Zt1iKbxecgwh1nTsm/wtkNydTNJepHOJLoplIoGzjkJ2f3pQOvkq54/vM6PXlcgFwwzf/B
5OXjKBW7or0y15Qrhgf8ImaC8YTLnoIb+LP+wSAj6JcxOIFLyfy6AI06t+aN80coyCdugbquf18y
7SmweIcj8O3/Vy0glhwflaTm35dhz8thcusR2o/VD2DIJLX5lRjShcdoO0UZGn8J0CvlHLtuHNq9
A1SYwJcJNvaJM96XLNkyyJuylp+FB1qnj9KjFKyTPn+uRJKbcOAyGhxE1bVTXLWtWP+P02q/Bvin
WDMgMb7S5gvhXeMdR7WEzaxkc2WBt75DJoKZLo3uwb7B+q1IoxsnBwfVQjtNhQwPkkfdilAG9UFP
yoBLuiKjazRyTTnQVqDTF1LxcS25Z4RXqwpLqQGbD4AncdDYkjGBr4rEzldazhiIMP2ykv90iLIa
qia4v+/eYoj7WaHote+AQ/sU5rGEZi8cClcmI5jcwlucCblgAn75bK/texZWtY27rjbdbGmAk4oa
klTJCqDdtACEuiv5p3J7enRe89Dp+mJXzRz9/cLAiWJ03oVPKvrR/J/qM/824nnZZoytDuhYI+Ef
uPXXHOvYHJBXsMbWnkoTXhnkjm4Td4It4Q8s5J/yTGnNtFuEd5xEMtsc2e/slT0IhrZAjUZYKfHS
er7O0tw7KdZr67HdSc09Zud2fl2Q5xSYkPo2CtGmn74Vq1sx7RBKWCWxWVeATDhiUusVXhUp7zSD
rzjvjimPlTR2NregRCys+UZUX/zdOh/UBKIfYMBqPHaFGucx7J/fGwzY4obITSMy6dHR9t8K9hE8
h7TTJA64HlD7Bq27d1QTnnviFhVy4crGKo/dJr3nPHtu6Lo5mTMWcjpV6jWY/tRc4eOXSBjaQ144
20i//YBSRU/junrKdV5P+sPwN4qKbMBEbiE9FMIarrU/yUOyMSWbjeIKh1ICVI1LH5b76Xp+yhib
JcwZHtCijal7JRLs2e4vEqT8BIN7vkNkZaj1IQEJ0qXhsZMzufMbY8YyllmUoOstnIPAoC1d3cdk
x5oShqaczsnrdtkchEXD5ayXnWIBYRctlAiwafQ5NIE0UGY7jC8W7nC5tCBwpjCobziTqO0PKOV3
Se9j062GcQI0yQCYr8cIgnIUEubwcZ0igdyZ2Pn2bKxqfpi5clhlO2AolWOnE9V4/wPAkWughbqd
Z3fk9HmXF5JCbqKx4Li28p84ywEWwf6KbsnhLyPDz6Z8z21/7iBv9FBaeTLmU58uaqR7pXDs8VwD
YEiVRr3C1DOKVRznEWe4r9IhyvAth8clte5OYoJsZe9+UVRgNNgyW8rubHwtsL632X7w602P2RZT
qeF9xb4a7DYfPnc6xsMxII/qXMWrHF4nj3H5m+R6WBrUXeL4i4Y38fAuBZv9uVZ89GIY+taOFN8+
uthAFZ9WnjkUvb5TTIAVp4SSfCZIiXMgPBxytw6Kkr4CnePBOHQpKIusi/Oz3yJ30C9veCWt3lUq
RZL8N5BnCxUNTaMQtXJ2IUVglHEoZnMBYGAZoN13wF/FtG+1jCz0IsbaBqZJfe2W7jLWm7LoUZK1
C1hjbTfmfosaaCqaxtZUK5s6qo4SInWiHQ0GF7VOzcnlOg+sKS+RI6/LO14fvZqINRsA6Fb0QOix
Y3LSnGKGWcEE7kcRe3psJPvn3U9esEC+drfpueCIzlYVJhYQRAztKa2MHsFFURotB1b7j4LzSMfM
gGIQvfyWPxQNu1cfpddf10AMQgerjYebMikan5fJVyGdSgdY0oI2jIfNfY0nRr2YGSTxrhtu1/lK
08tgX3mX9/NKzwz1P/xH4ym5GprB/fshdJqbwIBT5DMwvOJl4dnrZvO/hP6Ehf43pq89flNtP18R
0t/RHfLRkcr1zqR3dEXn6nc4zJt04NOb8WYkJ2GrGLxwQmUr316T4Dj20cVN/B/L4KCJNt5FmZsL
UUCc+LIOf61ouGvPPwYHQS4H9N9DEGvZs+m6dbWpCPX1AHW+6iGpS3FL4R2VTAs/A1xNp/a1adTN
1OEuDYGrXD9gV+OHHZfVJpHXlFJteN0JNJkg7ayk9N3b7WxZUG4FXAiAA9XdjsSSxvy8wzZQK5wX
sZdMBe8FL6UgEj4bpE3UvNn1qXy2K7YVE5QgyTb7VQhExq/i32EEdHsEaG1nPT6/GBoxbsbLD1AM
Xjc8M7KrMxIxnMOwLneg7jKl1Y6yXPAyK4pGpXuH18Fe7Jny9j60VfdrM63e0x0C5mR/MLB+juIt
d55jRvk+Jbl35AI/tVWY6wb1SSAnCDpnw/1s+zOd88xer/kVNWUHgZkFuHEsgTXRgzmuXuVvoGBa
JFvO6LjzEbg9HCNVqLMNCXxU66Xq0Yknx5gD9L2ZjHkmT4xCD+IWINB/qAfI3ELWXmtGsa7kqMcQ
XrXpDi/8MtTz98+ATMkP2Pb/JMKAer6jchhs/5U8JL/7rApq385ARXk8qpsUoQgZMWMNNd4Df8Ae
1Xcxno8fXeBfxzYSlgN4Q2V0+M3pnQLNmMgJZ+liQu6IlN620kdhG7V2NGZVXZdPYleN4gWJdN7b
TsI+twhlm54Fqei+Hh1Ou176kLF/WYNTzCoMP7RONcUlKL3gA0AuwCys8ULejXtW+kv4YaNDAFZP
Ug6BPVGvLbvVbU8xEOHW5di+2fobttYgpe0fzVSJDCZ7UywJ/MHpkNISpd5qUeIBOsxsytlfrxmy
/O38vPhZ1W/mLA2Z7wBaQyMaACj/bt1jMRQ4Wd4+vCBTKfKBZj8BoQSFcT1nKZ6q1+9jMth0aeaA
/aG67JrPcWUmR9A/k9Ankn+TvA9BorBoMS15hZz55l+k43v9D7Y2gOtelUgqptSTBVEs49HgZ8jK
8a4YDgqES42oMHwOjhKWa18Igt7A6YiZaGz5FteRbE/u9ahIM4HXKfECprf9RDYVxzapVW4LS4eI
HCeOMmd6tysV8NgvSwJIvQAXujMUpcDSQdY0c+wpOSD+gNVh7k4g/7N2Hihbh7NmQVqv286hlixa
S6UN9Ey9dnDUA4z2uwrSXTJVwWEXcYtx7kTBxJiDgyZ/c9pCivS5+Ntkgvjuf6RN/ukLUkEAn/OC
RAu8sy5QNT7VeCsOFoVW7lAyzrynx6DtKGyo2Zs7qBNmBJ12QmjZnmD0PBLwGQGQB+LeYY9ZPfTe
PNcC9CQH51XxAdQBcREA7tMFD4nKV8rNYBevwsDMRfDMydcIYzc/RHQosU/6hTOhNSik+7itIxpt
e309nOjalgbkss5YTzi5XZ5upr/7ZjWTmZKBr8/DFKUsyKM6fBY+sSCPkXkI6lqxIIlDkPj8tNnd
84XtfPr+2PPTukBiKTQE+gekaUQKPncHGn4IKvSp1P6cjsGTyB5uV4cuTf/5S1cQNRfAEAdGsw/B
DM2q1G+ptX5VjYWuf7dW1yMEQZEzsnQt0f1wCrzRAY+/unwhFGEw+u5UP7YmfDO/zkAQTsVGHQjH
EoHxKwFWmBg+GHMM/tGMETUO+/kAnPzsB70PZ4Wz6aAx8LuDAZFhkR3upw/HNgtVhTqjA2Yycwuw
pa3MJIhLLklO/maiL3P5upyF6VC8+aWwxjXlV9GS1YwGpPKVchtMLanjpInyT10WwToPSGIQAoEs
zn2+rkQUWcJHspR6rNfZegEjDsvay9XbDSejpfy25lMDlDM026mv7eTfN65jHsHUTo04yX9LWz/R
r+KnGkJkDYfIFpzjJ08mOhAN9qAwOycL6I84AM6St88y6+i2jm1Zh3qSSQJUz5vEzyjdzoJG0r7E
0k99kPT1mYr/oBBkf2u3tv0a55xwrcavWDT2YnXduIna4tviP9EHylNh6vywdm0czvJb3u/gl/Rz
tczxs5+y3XXYtZyKnGAVYt16L2gpGDuMgJtm4Vg6FAQBwcOSbYT3I9noWmXVS3NvoMEtiO6s/0zJ
XQbiAPOfeDhTQ+u81RmjPGlambrkR82jHRw2aDN9AwdppVJQBhhq3v6t7G5LsDV7rBwil6IcEF4d
TMIGGjHMjJm4Ee7PralpY6sPuYu8nEsVlpYvUNcylBXxGTaGJVfOJYKz+KwgWa+5Abh5yEvQfZdB
miLd5RZeehQMjI91/0VujS1u83+lbjeMkAKEYhEq8UQzJnCLS9fKiL1dYqbAiD7BxPI9O1CQXmdX
hwERQyZ0SnCqD+Wzbb5PdkvntVHCVWl/QXJuJitvRxJeIRbBBPXEdb64ahTRwRIwG70sQeYG+6Hp
LtXPJ2E16R1gqGsbKMXA8i03Rq57kvsY6LqQF+gGK67uf3WWcNKfptjbfdpQdJewPNbAu4UWQAex
xuxi8Cvll25ZqseDvnvnVQqBwvEFwcVAsYegdo9FeNATD9aruvgW6Z6VTiFQ2IPTrQy9ZDAgkV7v
+rN16RJ7/Mtt21OaoIVK48UAQiqZ17H4UhvxmCBIgkLQjPAdePgyXX+x1sEGwyhq1KOGytixzdd0
2phKGECSnW62t1L5KTUSFY/pYdOhyhKN95varrPswYB8Us9vsVOyYmrNyjmhcgi7aKcxtUl0e2r+
G1BWzbVC9oeMGZEdFPFj0lpxkezJkyZmadXb7RPkAe+26h2QdQk7jUxdNjJmNuljeftwQOCn9u59
AB/a1NfJb64IrlApFwHgYBOTYV5W8kRzYsvUL60edT3pEYEhkapsC2kVfBIBPs+3i80ZcXey1AAJ
ckwgrNs9qJaZavjyteXmik+oiXM9pBZ5UZPtxWp5tv1ag/g8w6bvDuy6kRv4ro+FxxXrzbS57Bfb
jEVlMny9HHpGoRrZADMFSoP1BSL4JW11YaZQKZFDmpdlmYkz+NyqXFtC+86MMblgMZb2CyqrGSnY
1IwpIPjzZo9zfwisHqispGMLjZqgNzFjegC/C8y/w/spz4JPStS7iqQZkSBD9BfZHi0q1pgBuZI8
ITSsnjVxJZ5lX3Gl9bsS4dA7jy0UQb6K7VeIcg68+QAbKtbejYMfYbJMBtgccj6exiBUIgflcXMD
8Ou8mtIhAgASd96izSKe/msTQmoR6Nir9Ms01e6i6bHTWq7wL56ZxbxoYrC1k54yue5Cmk8JHVja
QIEqbT+kwaehTMAfdLw2w9MOLnLyopS5oCS5yEAF66lm0IIK505DCQmX611SLAj68U34PvVg7u2I
jG15UGCjt4U9cyYq3aabzQ9CjNDW1C1VAFt4az5RAwz+llSGwzQdWgpx3t43IxVd647Fak9rPlcy
9ms0v5BoqZF4qm0chw4tZcvirOmUC4rjj8RI+ZwHTDAeTbm5FLB7EybWhf1Cn5i9I9nhOrqPD/qp
GtMcW0RIbInfV4fxJISczetuLiUoUpwOaZ5EA0CFfoBtM0xtiHyTbYlsudIJYidnJWgkFgueOcJ4
tbtTiYF8Vk4S1U25OBzT8ESCNTb7AHt2dCukZ3Q076+18d6AVM+BmKzWc2YkN/Cg7hyUiDs42fV1
jMo01QZHS0t4tvqVm6L/azqpWK0kRpzHW807uVFPu91Z8yHrUD1AhUaRwFvks/p1bRljNHCt9fJ+
Zn5RR8obFlE9KP/eijHDK9aqK6lcgVnrdZv7FDPQMVgS9HS8a9OIFaXQcNy6NF4gJG/bro0PuRlJ
StaaSzHNL4hW+rAogEI03uNQM6yNKKlGgFfO4PB3peAwL8aat3V7BC3K9GlNj4LdScDyeeGcJSEL
8dgK8hwAOz7jGHyQuMBbOc8W/wD5DSQvUqdmOUs7on6CaU9nbdWbK5JrV0JoFtTqgVVZcaKL9Z5b
NjUUPzc8hBVYRyXFOQRhgnKjLFvaLU0Ea05oI2/g8meHLM4xQFB0cMLqzPwIn9MZcGJIdMSdH2im
bDbSd6zPTqfokWZapIWfOsmiVva+VGp2MjgAbFAZhtUN9E1pqVedlpV6MAiLLTDTkMB+Tat8xn81
am1NArD6iYCOEMEMaDAg2crckwMgo/ofrlCho0JGInNvcjnkVW6zxDHk3Rsg5wGYsHDEtYlL5fVf
uvWiqNGC58gNhvVJtdTwlyrrKMIL5tG5psUsouAGG/n0+P2HCNobIFzeKtWjZ85VFcZGZM/zfOOy
rgwYbB2eh5GXWUe5LbG+a9BBj8La4JkW+QFLKeiLGC0ghX+l/4feY9v4BIHkMOOugWdXRbt4xSLb
r14RTmet7UogCD4hqGvOpGJ+BWQs+AimRvttTIgoM6DRCSI+DzkEb4EzPOeEmqqPr3j5bOYcT0oB
Se+d0QRVG5yLwcbjPBaQhSDW5tCcp6MdAewSHTrVBIW4BkJp5HMmNMl5piETTHi1+T0gyQreKq+a
7C7ibm66QLVqEK0lQ5QNpXYFqveXrXMrA5lPojhqFSYJ9z320mXfTROvEL63Vb1ZjFp44pRX2XvL
IJ+kUlPnG9yr/Bt0ItTnOSyEZvgyklbp8lUWIiPsjHE1NFdZW6xrLaYEoc2/fEIMmKvejtzYriZk
PV/2qX8wUEhsy/k1Sx3CF9Mjn22EnU4AxTvDWz112LZsCVZG6hWlFOtmhk5QM7piCNJPeDypXjcx
KI37qTkcqwjx6ZBZ8DJo+4T1M3+Wado87L8k+1OZt0xdOf5iBZD4ZgKghBZjOx081O4bSrxHSMwU
s11OI0OJHnQMsUcF0AQnDyRcOJsO2VU3bWvrBK4nL5kw8bwiJmk12Tr/nv3E/oBOGdosXxqEsH03
Xq/t9f7EQGnyNH/aiAHyqnSP1Gsp2+B/jvUI8Fw4vUF3M1HsTRb5yTEwBw5fLm7LKKGMvBIrLCmW
o9QvgK4gSVx+vd10PT9y+4YZQmMJfmcqim5tZ8CeJVGP704so/8+vw3pZJvFCAV6RHaq2N1dkaDw
lgKn8Mu/8b42OFw7oOHqmIwBCiACu/LXka61LDoCfCPzZQ+2JBMGKoNAwdpxxWhJ4yPFVR8qQJSd
xE/4pI8Mq7F6RzHn/DqJaPf9Y0Y+D98ji4BF5VtOxDeEPL/9IxTrqHB8FjtgeN+YzDuTI62KNhvT
XjC7OaO+KsFCoP8xgInbSy4speLFC5fgj21Smu6AGO6k3it4JH7IwtFYk0zEhvOWIQe1r/f93cZX
dVLcqeWx5gO6JqPTNYoqTNbQE+426ylRPMUQ8H9JmOqFtlaM/cTi8YrTcDsetRu8lTr3nPC8BDmO
82AnAHrIWW6lJw1KbzE8Vcab5KpsolTwK+sqLZqfQXNNiBVKWJ/rvgo7jqH94OQ7ZSY+b/tulcLE
E9mUAHmgxNSF/eXaBote0CJPWR4owRT1b7aR1o74Nz0HQtGOkH4WVF+zXZ/orNP46DEmVbiRFhGd
rSQDuqCBEB2alBzaH6N5oxEcUv60uUYzTzeYfjIn3jQQeK/zMdkOWzMyes/lNEy72RhW8HjiYdYu
HOVMFGc8snO6dYCycveMyT5bfC/p6alqBEQVmZd/YS+OQFXodYO7GNiFOg5D/sNtHymIQatD9pDO
h4RBxLt7JfsNIULlxuB8HMho+N5IfZ5RUESewXxBmtpYtHQumOeGpdjDHFw4k1rWIrH/dOQVC7Or
rZTVhcuhkv7S1tT+Jj8vChoSAPGmd0Fdrr242x4W2cOjPtC7YR7NJzUd4OpNWDd0jcmD7W/+O6G2
0jAw7plura0008YgrzohtPUN5qWUmzbim6Sy53ilbAW6oYr/pkcKGziyFlJkW1NpXK/P1uUMO9Pp
H3wferEeYmCM+jwblbaicoMvpp1gTN5E+i3a+T+dHEhvxdOOnPAT/yUYGKS36RLpGL0MWMtZqm0l
k8f2fRLldBVmQf3qpnoJZcfYUfFjByrMVjL5G/5S3Cfele+Lt0dCFFd8QdRrUEkMrlrMToZ8BZmk
iot8/Q1tgHYjdjXhTe43h6d13YxjCrndMu54tO5LotuLQTxttgyXnYZPAG/DsaHWCcXqifR6N6Ep
woTwUtw8+5p4S6DiheZhKeZPBgdXf5oIirZBZROwDzngb82jayteVyYQGCOKo+WaKabD5JGg82at
tAJwfCwXnLBKPdxtGHq+l95s76k2CIad8owMidusyLw3iECMSUtfcq2xCj7efriJLTR/e3Vwu26I
KiERkauY6A6QM2IHfyxaC4djaQeQValXP6l4EtYd9/5Dl0eGZsKgeYYwMfY5VD9K/DQB93wugh54
NU95remlonKsv4KxQ9mjvlnOO02aozXYt9yiZBAWphu4nj0nsyxL9QunnqLyyHOQrwq2UfKxOHsi
TLbuf2CBVPnZneOaA8D48iRYtRwv2G09jahK6hZoJzQD0M3DE76HPUMxdINWg7HaV1YzQM3BQqfp
kEeHW4SfYk8UB9sPNs+9m+oy2pr7bGT2a+8fUUlJkPXQjsRHiy3NyJYZsJV3g0qQ6ilCCh73wxYu
luRo4Z36Vna7rVGbOQL2xMKSdnvASZqjCFQF+bFDoXpcTbCDN8eAHhFoAJHXQ7j8v5czruqO7opG
NTD60GK0h+8FwgUggJeRmb2wsidWa9x1pO7bQZ4O5L2aYoWONsDZkIy/B4PBZQtGIR216nvvbeEl
hVyrcyqDufOBXCCmgtXxmP5H6RhDOC747eFjaK3o2ZY92Hf4q9dtDvlAL3ObwmDuR9VHYp8g3FXd
Jy3UTNLSBDVe5mk3h5TTZa5aAdkCKfD1d7B/Lq3ZHwb4e62xwuMtz0uiKdp2bttHaKkNPwObL/WN
BAnOE5BWE4VyZ4MpzNk6Uk3in4eN4KMOEB31UhyFbEMielaK0SVoCAb8DYdZGlmUMfUTAdeOC/gN
0Zaz+wIYuDlIXV+LJSumReQ0pMyFp53zVcFzyklzFEgmwCPRRp56lhXu3aB0Yf9pUrELss/MKEi7
PjBYk19ssxKE/VM3gXu2FBQQSjMnpXGXxkEt9EUNjACN8Yq+9vChI+bO4qvRPzoXWA/DfcSnGFln
YSw6OBWUUA7Q3ncb+mPRCOL6V32vxDMuj1LYMVfdxL3J8BFQN/vHDYbR0PHAVQbqaSPFG8C2mHfR
kUadnuFTv0N3/h/deZS63tY2R+2krHh6WAAHsWEUGoLde5MzvnSIk2oLiVqlD5dBnX+HjWNENsOl
OrWiCgmMHvTO7Yy7Cb/O3hYVDDvTOQbkXhjyDeOBvEhwDWjCSTdcrX7NgYeAdi4mh5ASXdp5IaMA
oUimc1OPIvBU9IfhRIFzDaZEBR6ZsVQgp8FFyVHnHvYXRMvI7jNbFYCMyvI4Fc1GqYQmCHMQroAv
R/cdUjDcub6Kw0WLj13JOC4wBqn22ijYqEP26uKGZFAi2At9Lvj1s/Ta0AmNz+PbQHC1MyvQNKWT
xS2YQRYSgBXO9VTGJ+8nMAvjfUoouiyPlmaqJwQ7AKGNhWKPLV1oE4e2XuxjT1h63j/TKBlYqSlX
zYteTBzPjkiaP71PRev8GyaMCjdvhP4MpI9wm66739zaMcgE85Syk2zwtO+eiqlXk4y0Ek2FoRPj
3/9/x0dkHwxRWzOzfszKIlJdhq008CymCUV0U3BQmwlJLODjWwDigw4LdRx0aIxZuqwYRwkkGC7k
4crC+hlVKlwwZU6C7q7TFa1LphKE3i7HvukFU1/2bEtIOVVXcC+C2yeGrR9h7a2ODolDfIxf13UR
5nwKEbqgXqNLAXTZcp6z0jPnuyFIh6PEWqHVC+9mmItLkfPPorAtIgIoSXsYU0Pyz0P+PE8nRdA1
Ml8Ftc+PLAp65aCnvD6v2NqTGJTzvYm4zXus8OS7vBCzZdziqMTSRIGYl6VaMSQR+DTVLLbBuA28
f66IQpK2yqR1wqT//voIZMq+n1BPWlD7csZzrxUxsJlgp6vFMAKYYnDy9IzdQ9pjPnQLvZQ1bX5v
f7+sZq1Fue9ZJKiKnIoeMzhSsAtkd+1YM/E/CRHKOLDmhidUOJ3na76e01iOcVeFHC/xz49PFkWo
kK5c3xAnGadXLicL8opLiliF9hP4LK5bQbwYiOiglfe7zP3uardf3HqK7vxnX9u1Yhg3Vm9GjMY/
K3KW9VT9M2+hM8e2JFtRlwYH2y2jzy97AJa4Q2HwPuN/Sw9Z8fzC8uYZPBntafVESNTnUxmxWfH+
BtKZMGRcUc1kdB5NqozK7nbd5IRIlcyqWCCJDFDs7x96hzwMOhzVX9ioqod8F12Vb5kBxJfiWa3A
wbBGgBdV6v5d0TQG2o7ZTwQ1Ecr3ocXXkHsk4fyjrzysGzaoOuBxLYuDcOrUioY6gPYJHdM12STu
XqlX7FsLxL6Fxyuv2C3bsadhEvGNXLNDxoD+qJA4n0StQzMIRI/fl6liQ/yk8IA5AcA38ffh0KRh
UD7aQLSXIm81IKSClj5b9KHbK2JmrOMcZbf4AX3lWeNltKF4Un4T/jpvbqTK4sXARe0H6JmUsYT0
4cHDaFWoNtQjafjELW2epFauEbhCWCaTZ8FlF1bE1XdT9fzs1G3R8vSldtD/GkJ1Xyz+8OZspYBf
U0xB9B7k9b5M0IBelPg4G5kX4TPo9XbHoMamSv/LJ+UA99iNbPth8itp7momoUf9N0k3XPrR4/2h
3F+E5QivpGxbCgWIXXgY15KG4FMIDUxaW7VvvUp91iZRfgJDexRK6TFzVnOtiLnzcClQ6pCKCaV1
VHcHvlswgfQOilq5XT7AJHVPj7IsWud5XB+m0zqb5Rv0E7Z3HYTnkrzXE4djfBALr1uqf21h49Tk
CSCdO845XyTPs3PUGrQYTjaEihdA5ss9N/RLWIeftzf0agT9922wbue+Vo5bIcU8Tr3kuBY3tYf5
QHz6H5JrFskmMD23gZ6F8WINv56Ycjx3V+sUopu6i8/12DYYA3V+uuqRv8thVC0uugsRFo5jfqBo
hsoboSRnMzP4KlwtJ3CqtxjNcVqB6dvTyEiLUHiD5I+32wdjetqxzmmTh1uJTxbo4Fnp6ySqc0B+
avmATHHLCI3ug6l4MiRR2Qp+bd+plHSam57GOb4XyvaY2XvEhNkt6cQMsw53qS7uASVWD+vqRCgo
9o3jnvrb4ojKANjLw+d9u/oU2kSStJPE3tmxmp8D0MEm70ZzO/IKIYKqhGqENO2RjYMlXE+DUzuy
H/fbwVQO92FIf5O4/uB6KGHMTIH6fLOqMZFoMwQvF7o93zSZkHHpd+GGi0YOre1r5W6Yu2rhAKUQ
v1xa4sbVsJZ5IiZWwyBdAuJZWS/BfqopYvDaWoAjym+UWlm9HaJYMt4wLpMHhgJ+1g6eEm+j9Ei7
yaO4gQbDtTO2xgVwYhB0tWxf1+DVhk/Zqj7cUKoucVV8mp3oBcVG0sfHo7jGce0PtuHb/2MrpIDq
5Ah+kgKIcZW8D6+PyKb0L7HxsYSW98kpHfilzFjZ2VWMHHnl6SMjLP2M6KoCphQgb5f6KE2ckmHJ
N3FlRcsVbU9RlWind9nFqyEVikAwcWf0JmL5+YtB/UxGc0pYzhCqETqXz0l95SlXPNUKMLW7RH+b
/IfuMZLAM/GMgvTZZdExVvgQTb3sUVmzK1l3BChVI1OKwMHI8hHQqwBzPhIW6frXvUZYoDuzw3W9
hBDt84Gn31RxLnEUL3U8DNGPufmWsinMsEH7R7xc/TWKFRxbtJuuxOmO9B8E3t+4QwFwKSZ0FnQk
1aJFuKspws0OWsaeE58VpBfI2pBX6AfYNxYuWWfouPvl4ueIKLd9EMvfAZSA4Qf92BXkhQFCAAyx
q5p5bEfmlEKibFEBQniu0C2lqLETiFX/wllMGZG3yCZrm2t/KnSOslWTASuXhJI5lzrElk+aasU4
3xg+0ZsNrA2AK52jEgyI2x0qRxQZVr7uTyCEMyDGI8XmNuZZSKTeL9fJK4N0GeilzIy9zi5wraGm
fsvmpiUaTA56bRiy+SseFhCqPr+bgfT0TmnwMRZyb2uUfqznq8WxfBEjluvZMeLu9gFhKfyK8GZq
mnuc3JQMTNcUKuoJOAU8vo7pbZXvP2fI9mTtGCHBh3LnEBsPlrD3yzyGSVGIhYk84szNZ4WpzdUA
8ZpsZaoF8lNbOl/s2FjUNddKaL118w16xFzHGLR0mtv/y2KkRmUfDB3WbO+R6nftmg7O2rd+qcDD
OXy5ZbH2PdRRLZEz2c4K7zhqmBj+PxBiYORQHP4uquJVAMkaFR9WDmhDhqzRJmwRyCDtWNwVkf+J
dKDjE7qvl/IOmYngFOP5mPjpdPRaH2HDukpZvNdWB6RqlpdVMomx4tsAqfVMdMqZ1PNO62BgoHHR
QRA1szADALx2iDNWlRzKuVxLtaX0Gb9aVOb5QD1T/s5XT/w6H/x1DBNS07MpHOc25HqNoODVPjqO
SkF5qb7glX6p18NmJINzk7eGAFnNeSxH/xAND7IW3gSngQIkn8BSsfiDET/Zx0RP0jqQq0E+VvEs
bpX0utgUNEbAKGDlRVbRuxnEeVeMnkJvbU20VrwRSd/HgSjB8UK6her2xlgEztTWjk0mYwBwZu04
MuXwOLykwKYwIN5NWLpHrm34hElKHV/cSs7KJmdrEJh47URoINlYFbhURp1hGX8CMWUIw+1+v28E
6mfSAThAF98W8JwAOYj2imsvIiQL1tsYH0iqGuMZUx7ty5QZ6iJ7+kGyCzVZDicetNbBvskgmiNN
AuW5bXW3g2xMQfqbyPHIcx1vRMVim4jCtoA7wVxUL84vTJJ8/z1d7zt08TLYFojAK43a7JVDRw/F
F0LNNR2VWmI7DgJmXW/OuCkom7u4TiBfWt+T5VqdJVe2KrTdHPZ164VYE1iJp+7qXmDfWBSEUuqn
lSUXIEppLcrxjas9xXfMydbkW8oHmWcBgK8r1ikqphlN7KFpbjz4aO1XLpdsqyk39cvgjhr3tg1p
eGNtVvOyMshgW1XiBmpt89cdx2Qlgv6UCArT5TsrQCk9v8VAXGn1xJgY4rs8PqtgXp8ITWlTj2X4
ird02r1uqqb3eiay0YCNo3QlLXc2Nlj2zXaXODCDi1DiVvqTr/+/uxKE+1AWs3GN3MG1JRXI2atZ
oVrVt9fttwqOursF3ByXRjZulYrYTizplTJDpfmUqJJiNy+E3sME3vLmOzWjNPva7kumNUCjeiM6
nhEvM/pHMi+Skd799xTSjDsXBrDkmZQHKcrp8I7g1gIIn7gTWP9LJWSKkQEJHQjVtSRMdv6iHzkv
O0VALvBdopesW7oZz/PKZ7dOnqMnU8IVYmGYh0waGywjuZoUH+5FCaO3Tceo8yZh/lJzKyUT+eTM
6oBd/L+rctBZlFcLb++JQcOmQ9qAmKu371nSz5miP9iRWoCRk6Ew0rxK66AmtK6gCi4sqKf6uLLv
kBOe5ptcUjDNbw3eqZiNEkzKwlPPELEKkkcslzCZJCTECTFTToXdP6K+okwnnE+q6iPN1zpXJG1+
SpYHiB28ZtVi2jJxva08cffrdHP3COI68Ypr/lyHGi0aOnewj608cdKPLe7NIvy0seRX9sox1b3t
kfBZvTI9IMdzRZ8sADgHv8uimoVIkdrHVt+DTHOBgLCa97u/CFYYAbQyDfgwfzpf2zC3lePoXiHg
ikjpH+vaw+LOq5gryoeEvRslT/Gyhw5IJthbZ+oXbK0l1rENXG65B4FJsy4JaiYXoYVitAyImQeI
Nqeu+PQ2CmItgZAKBq6q1Sx6DtOIuYdsD7x1aCVPhrjdKOB/AoSee/RvARXy1Hjs4EhWecadR8Pd
F0HtAhffOShmw4xwh4hhvocvSivIkw6wJUYvOCpr4xKfYIM//mMFbXZ/6Merv0ZCx3t6EOU33930
gaotSoWth5mGgt53ba1G87AhOU53jEY1jZC2U1X1BxPLBB8PHQSzLvJIBkdLNCg/OdFWoYHQfPlt
mf9Mo/2zqcHAV8aPy3J0PCQI8v5Fv/6BcQjaeYYshdDlCgUeJx9cktDM+BxtsIKYAzVlp9e1RO4e
KKRZFW7Ysf0uj7oubqbP8rKSuwRHTZQEVUE9ugZMyGNHv0ddi/Ikc5BzG1Q9kyLEFkCa5HmDU7QH
tEsMVb4UKEACYzqrTc9ker8NUsv0hRfqv1A2wdOtJMBjlWwQedr90On8jZ97oBBjilfEMleI5S0K
6hcOCBN4B3uYpCOXUBf8JWDgqdEjbXrC4x9cncwsS94s6N5LOgcI82VxF9tWzW6ymJVzytMRDjzW
INNC+pHZ/XIMPkNWyvVE1EDo/UxkgRW4fMO3SIElR7qSM1W40/HYo8FFyV9P+s1c0drgzGHTdDPw
qtOwAt9/TrJCszgNkJfuGiEyz0g/1is6kOCIDajRhbQo5z2Cr9TvKDTrn8Cv0bEVRZo4QKBc+re8
YFrxt0kSTfOk9OXVWx2ExoOtRfpke3/x/LRrEUgSE7ilujHIwCfBcYaiJmxXIdybmo0JCsKvxo/b
HQz4UbZxG5Fsb0VTf57a1fM2DKAGmODZ8o/6oSBIwnDl/yV9/yg/ju53C0/uGBYMcDGd5DAkD/vg
9XJvhy2F+szW1Qqh4xpmKYwZ/C82vn4mvcIzHriZNDQ4AjPqhg9b7hKu1m1i0k2ShLzf3V+3Ouhn
mtDuKrzRv3O7iDoPYKotPyoOSjEGob1XbcvAGejBVpX0IZQdQeiZfUi4+ACn4ofIwyWro8AO2TbB
ZtxiCY5lpFV/bD4zUyHN2ItcouT7+fDv8K2OzK14TKxxAt1J3Ycz3RXPCsdhX+UIX5P5gmm87mX6
Jm2Wyg5n/Ff8KxMQX1BfaTWfEJtZnNZBU+TdFsB3mH81raJwLxX9Cv3jIX/XhJCA+/R+NBLGIzbL
u2gZ3u98NOTrkKqryBQLkZUGN42QAbqxFl6dT1ePIY04WhtZMpH5QA5b7Ul+YYN3EpgDjkWNcG0i
G83gLB/ZGdRP5qUOq/JXWJxpnflY3iEdiYQ6a0E3iCrw8qEqmZnl/Ag3zEU5NY4l2VaFGCD/ZvYm
C4gLl4GVeQ4YkzVm7B8bFgto2DZBHPg5dFwbRA+v9HPoiWrTBd0TjVb2Y9Ht2WZkPevUomFidhuj
LfibTPTZNi2BTvtgaEGBOzPoMC+owGTGzsb1PzsRKdLYXUlr8FzeG7g4Ud0OsMRb8LeanS366m6W
Ab20RuYqnsaw3X6Y1wB/euAijVRg8wLAf3V48F1HO3SAm4AwKG3x6duA0h6Bqp6gju3+wnv4mjs8
3gsfJgOiMh3FKloMY2epbDdIoUnOzXG3WQ4MKN298wkznRD2JhvzxdSTtAEngpt4Ksv4hVUZurqb
5HIhYLSpV1+JefbVExqiLyyIU+6Z/A2U/oCxqwV2XIQu9CRa1HiO1KhGl80ry/D3+bXbgg4b2vvD
U2rANLOVyLDZBKEGmH+e2t+eAFW1vQQKMFxxlixZeSJ+E4LyAfP1KQrh+tD/YlwhfdjDjcfia5Fb
4f+Gqu1qP3SfaCcWAqvi+DY8DoX/M5UYI2l290MQGSd9Je0qjFT72su0zvWour221UZqolHv/vDl
sbGaHyA9eTCx7p69BLP73RvIld9jyw39WSAPZaeJ1aHLsSvBHjqlw1++FMrcBX4ZwfnR2Efxyz/a
2T1EIqU3adovto6LU3O4UJ4x9CSZ1YkDSC8RwAl9ubkqxGUuXA36UKc/KNjAebCKNedA9AlPpRQu
8ULYze881zsnAgck757/rPE+X2XmhzHfYFBDHCutI6MWZp1IN2pzGPK4JCfAVEB+GXcIPCbUNxwM
7DKK6YuicWlLVcJOExl28JrP6kBESFRRLhC30cY30fzK92kHzCFD6BOD+N70YSg2w2YjtbITuC/f
WLO/e0+DTg4O5u7sQ++4Q7G4NOOb3rzp5xtL9Z8kcD6P4NAyC9ASXPPRBE7fZbvyjfyHW19+k5L9
9cAKfbau0MSS4n3rrCw3U3picRH4xDU+PtqneTdGrBWpNaPyY6Havl27084NocxCNl/J6d6VcGMi
osuJIcv3Lc52IpbQuemPThBdU/dmzZJ/o3SYQOGN3aN5YiBS0O1xzYClc9yZ+cqLi9KuKfPZS0gg
SrcozIEcLMsnD+BhOuRAoWrY/RPUHb3xWabINdcMd48FOVm7kjIdGRz8Qq3vqwAaAEpnBD1xkcc0
Lp7MRZ2P6/Gs6CwfG9BQbrZujGbA7QffwWBxydc7PfsyoqlsR2TwOFb3206/s3I3+fGbpxKvDKEs
FOsJ0wprQohV5xT3dq4dxj4xHdftFomtOIzYao0fKuF6AyYNnLcjt5Zh+9uk1OdirFDllqnkzjRS
b3C/pvPpSidS0KB5D0D9ZQbi4IEIuOwCu24yjsDaSbziSzjy0l25ULGmw6cm0PRIWfXCpat+fCKh
PeDz0qr2DQ73NZkjX+dpQXfo7WvKLObCPcZEr7WBGxCgHT2HsrvgkJtR/WA33MhVmSMQ8Rzj3R1i
xr12wv3KoYZiLpHBhw51TNxwjycrBKBmiOERPWebD+C5DDLFa+pZG0ErlfTCgpFU/Ft1ecrKfGN1
Zy/GJaFDPKck5I1jPzGCbYYwhLom3WvRd0uQINthLU/HlGApprfSncZ1ZrQqV7H9/zxUkbGpY40K
mOkhXBGgMyluIeTiGdm8DE+uW3UN6lvpOjH2mpqdxZrwQF291EmZw/guSvcYWVO8gX7CQCl/VmkR
z7f+oarb1ktxM2eT+fk1TKlfZ0iTcYSLtPGBS90ek8Otl24P90i4KVG10Sf7N+t79g9W0ogVDxl7
rStPyy9Gi/Hs1LfGZdDfy/fZ0Tv/zM5U4bu6aG8nc2uyJK9AVcby3zdweNcGMa86k01AcvOCLo3t
hmyxGetzlMjNYO8Fuv5XEJpgcr004RUETL18zVww00Bi0AyAi0BsAzTTteHaELegllxB7lpumWTG
X/o2D9I+Td3maYuzHmexsRzkv2hT0UHEYGTPXaeUQAWEPVaaXUBU8VC+H/pbHq4QZhIgGhB6+mH8
d63gJVXo3jooMFoSNOCyamEL96oz0bze+QKTcvTgmApGGa/RkHee+tzl6mwww1paigwGGVkprqAe
6Ke74LxA7l0UL0Al384v9ct9sPsWP7JuU02NceA3TOV+DIfsVZTNMFhGgorTCakp1Pcw8B0xSBme
o93G0dUn0TPia63boAUEqMbYPPomzp62v1x+xFqvlY5mcskaX2GW01T1rn6EUzx/Jk3q4GPgq2lk
BR7SUsN4EgvMRg6agxbz4n0vE/JaddEU3eKr2y+LQrXTMjcJZDZ9zVutx6yxp0N3oNWfMOYujWxJ
Dq6FzanjJD7bMIK5NOUSrFxtmPN1KTp/SeTh41TyxOpgfxsy94+ZUADTpRJDm4DY839hJhQhViNm
N3lvQuj8MazsM4zcAv5CiYqUBKdYUpus2wasYE23CXmhtQHFzd/d15QVPaFdgobHy59RU1PQM9kD
anuIpRqeHr2J0IvRqsGEMLswBrk18bnWparP9BC/rd6KS4/Z+mB8yzMgpQt3n7GaRbvB3h6N1bpq
tmIUDZmReUJOI0nakdYhimapFH/mZoR6Zq+lsmCwl6zYVrYpLhzrlm3Hz1KQG2Ljj6MuDZVKgl8U
YtpOh0zS5UMpaBQ09CclM0ynxycLMSKoaRk9aubb9eulLXCs4g9f5mUFiYFXiiXcvXeB8Am2ROgk
uhuc1zPpcwg+U1QW9WkN+L4MCS5oggDdARsyp6VBIdEyyfYkDTnNI7ZLsCDqOvS3++o5k5bGiiM+
m2/gOdC1QA+C1Yq46SBpJOQYmScub58jmZW2CWshABE6P5n+FIub6Grb7jFxBxOqumGJsZSht5TP
Vd4/5rLxHazUZj4VtSGtlccCow4pmmVfgks0wk2xlkvaBfJ50wZ2Vgki2YSujBQ7DV2eV/4CBnE6
9L3/uybi4FpO7FM0SbctGDJoQq4Jd4rmJkO9kDw8cl8b1Q/+8EkmgUz7iMY7Imk9eTgIMaytpx6H
+JF/r6BJ3seTiD/jNnwH1vsfbkM9eEnzQIbbfpw5EyFghlo6OuJCOb9iXqckyzox42no1MCUYD5D
yUA0CA1k6t4zgHUY8yjdxFrtOq5lM7wSSBLg2pm/mD011MXnwxUwpFuoR88Yaq8lMrgxfFdJc9lz
1dSVwfAx8rny5qSuV0l4gTTs1s2D4PF28FV0ToCSuZBrcnyqgbp/reoa/uvExLeVLOEto2LJDi10
dR2X1ZxxKyQ5nVcc/fDkhk/z8r9qENUg0YO8rVAdyoHqzdobnoUuoXspIIPGUczt3/6h/KTlx0K3
06RA49w5G9884RCNDKIKj7BrMrc0ZDiE8JoEWAQpcdiXL0q0BHOxGHx6FDRygzQLLC77Y5qUmE0j
gxIj7q6WXdPAG8vK9fPN28ifJLSGSo3vNvBVxT8PiS92pJJfmt3+ODQZsUk6XFPe3HXXJqECNM9X
qvEKwG9GnCXhkkN30e4Fx4gVuRaFcyzKoMaSsN2whb4HgNOLa0luQsBcfbP1CCFiK9klIEKAtIGl
SXvn89JIg598Thr8IvFUf2gi4VuMKZ6ODwM0d7W/eyoh3ycGFREi5kzmmdxFpBg0npKDUsbQjOha
0+diMtgLW3VYNd2SYaDc78X5hAwDmehZ4rCPV5qaSe3WMN/+ysRb9IvBR6MfrG5G7tjmoRKZOonX
yLFSdtE6+xXi6YdogeO7By+oesWynuplnLH9PsGbOGsgLf0FC74xibr3O+aLAsVnoTaXx5L1FHd+
CVszE7ouVde4NRRsBaYyZFUjHihRqzL11h+8epfURCZyHp+41e6MPLx3pWv0AQ7srU+C8kUNc6ro
IMdxpmDORiBTd/Hiyk36JF/oGV/pDM/PaQCtpNIxnL20V+gb1SsIniHsugCI8Bkz/r6LQM6dshyk
bxvrsQsBBGIWJmYTdBMbicwpowk4AKtcHeppVtcKiYFGIfQDr+6FYw5Zj/QxsCOIfVJ7jWRwkAo/
mXd9glHKCBB/SdD/Pb8trlHUV+VtLkJ5jBj2TuPEgMINg6UAXcOSkvWB/dIulIikGIkMBCNuxaNG
iRrCnS1y8dtepaGxS95ICdlxHIAhh63YY9i/cWT/fEKmbGWquSuX65B1d8MNVzqL+J3lO0k/K9rg
gX30ovaL2EVQfrlBbspXL64w7suHlrFreipclMXP0Pjdaa5CjpsKVbEKz2mDux6cWcp40kNfaxmv
XistVV8Mf9uBjLl4Ui4k0cIeTDVYMVyZpXuuutUU+TLHaWu0LK3iKfIp2JWfOeL4dxljbGXqct28
qFnyH/RhkFRk79SS1kzZqbh4e/dh+sHYzompM85Nk5FZg9BMK1IbuEIrwjqLUTmPOSSD9b1ONjUt
9wuL1t1KEkbwuiWFKdMIV6q7/quINIkrBiINcVUmU2r6PRZyjS8X6WGvbjFttoSD1iKd9tgq+Erk
7DK/yW76HoKxo9F7cIYg9OhKY7kTcAgNInEJAxJAZiB11z48e/BXFmSUS79M9ji792AMTZq1yslR
yjS53iCpsbSwHCp3PbkCgSuMPq0T/tlvYjozWV04kaUv2k41TzvKPmOXoU2itufMbbf3AsETXqKV
GpI9hZ907JkDC/Ngf3z7pxSoiEXjErwtrwAFqHwH7jlGqhQoIKH6DfJ2qd3c3gfnykYr1qNYaGaA
11MqXulY4sjBd7tjXaG8p8WoinfpNfITkACuDPvOyO7eh9dnsnoobVqVy0eLA+w/W4ekwTSZJXpc
tOtOjY6Mkx7Vxc+VFgO98vRjvraya2h1HFPwjDC1Ulg1tx2mfbvNLKzdwpeGszy8oJaqBLA30Rut
ZgV8M7kTvyPFF/g5BM4DHDqY4WWPS8EJa2ciZORy+uJNGDEMp2e1zZhgkebCyF1w+H17WfJmojqm
x+qyv2omURam0ll1mYWanvQe7QPjcOhgGFJ9+eFM7BRzVJptdydA2R3C3dmOSLZniE7QFXTpzp1e
eQIvlUvbKmkOIVs6cqkYvpjbTRf6gMUKLIMyNHVABwifUMDJWUkteIjmpaW16OZLGeL/d82V01FC
UCjakrOY8wjDa+zGQLvU988x7wV2SwElAmIjhU5Oxe0svynVQbvn4+ueICIYoMUL1bja9ZO9MhYg
A0UpU7DxzISp3tUJE86reqlUaNJ2FTDpoTJFIsK+2A2f6pc+VRMy2lKE8OH9gtiEH2OK5tTfpqKz
q+If8cTK7PkSw5+ucOPG4h84yhsU70NbapwHsJcag47/14P3y7cTGQWv3pMyJmNUrPiCu03FIR3/
eyzCSV6R9VPFP84Ds23L7dgeldI0vZ1yEM1T/1CdUpBYHBYl97pHcPaOC/xQ4pFyeTEuAXnEiW9D
TjsczqJM5tSvIFAG1KgY9SqxaxoVe1LklbfKJyyE5lNG6xy/BDmGK7paZqvxitXl24jD7O+9OS/U
X2Jh043haoo4S4Gr6oZxTGXC+7t5ATKoHhge//Bzy+KX9eG6Nz54WiEHp+7j6T5VGa5trP1WlLbO
UJjKQrO3l/ImlYk0g5K/E8jAuKYXmB04ohLRLRBCUyxdIdttd8vsw8C6c2gMeAVwpTTWAka3sjGd
s1vH0IN+6RvbE2e8hLBujaH0SlhwdOxAua0rcZAfEZiGbJFpO+VeP3dwrYETk/8HdkBJMZGSPGTv
pBZ6C19Oc6PMu7O7zMbzpxMyOIrwkc1543Ju6EoOtVzWtqxamyzEqg5oQe/MAVij2Q4jb/hYFTNM
/3EWtLm8uQs1owtBayT+UppaEM6Z9A+xvnMod7UXP5kf9bJVZDxx49lwaKXps2eH2azbDKHX8nCP
cVBZmtYODE5tSpQouPmUuyaKIZxLSnAHtz8pOZC1fE/JkdTep67sR/5T2tA8NbhYXkUInp+x9l9Y
sVkYdESXXg/Ix4ECpyHXUPFH2IWka6j+leE2ws635RSl2FGXRGSvwfmTyy0/SrjO6d7t55W1uzfP
yp85dqTTyy0IKg3abfXbhcVJk/hGAO7+WsebUWy6X2alDLFTxYn7KjzOfMXk/u+X5sPz1nv5E7OA
wd7erq1dY9YnbU1tZrEswpF49XmZVYEQPrR0+RU9pWRCgxNMIsiyxf+yi4f9wSwmrlt0TSe81dF8
iOubRFqzwwYFhWr/x5KhRouinkzPZpSqcLd/WRb+7XbqaHlBio4EZ7PPgOGDK3nqoWtfPy2t4d7i
TXB4DDT0t0YZ5v/eZnYfWiF9kKwmKb+FT4ZWbGjGItDTTJskKNGTmdyYwhk23kmvVTnGiJlBcUoe
EbNqtM16KXUYe5smDTb2l01CBaoyGBLFWvWNVzeerW5wiDcjHGejlHrVk95lEBtU5XJpsrjr3k4N
+9n8rZxYxEM2aRokCICMjeV1ViqVvmCcq02Xl2ptNdUs2mWAiVq4uz8q6HYl/5RSVVdRcA45RmPA
u/iqBQd5RVujZpng+TuvyegKA1oXoB/OeDmapwVYggymWx1kfmy6v/MQJVsozIICYcPtztHt1xLW
2lTmLN/TnNPACHGGcDpiNeUZOKPBcJxFeS4h8GeyPeGPyS8Siv1OLYcNc76zuv2zU0aOQUggd4sL
e1sDKjzmEh7b+GduiVrnp/WdYyGZIsJCWhLD7ZO1IbXD6oDzHoupm5JfR+rynFVaxQtcjBcKyF47
DuxpbqJ4BUdaExO8iKATOf0JxSOPLGeLJrBH9Mk5xxqm8GHzJCT6iBb4fcxy7biaLemOFbwPcPcz
z1Y/F1s7gltoAfVnzys74AMg/wqRpPuPWj/BgQkrAa3QjLtSwMo+DDb8b18ul+FuZPQ5AJbrlvst
ZTIx0/AFCLNLEYhjFAEplYd20R8L0RRcoI2MmAmrX4mi/AJfysIp+TwM9F0ogAiC4RftzKhvICv1
RkLzcjl7iTTe+ZD/USm9QJp77WPXCSlCXQPsXzaAxifF6c3hYcNSscreZzgff6EB3teZCtPJdJaS
X4qE9niOlqrwc3F3a70pA6xe3g9l1zYUKD4WOYkBl9qyoOvxf156lb/QfibYlQDRBG61Kbp6I0KQ
98RQv7EKWEG/0VFc+bMLbAP6yZR5QRYKDC4e2XCDFEJgBiRUiY5D3yuz3acad2SygO+kLuRsoaT3
HNSYWoE0gRPqbjbOpHmV/sLzgqBdXRQgJo5ubwOJ9ZCCAwwAgO0ldU3PYrxdDhqNZWH90m/2yre4
oEls64sytYxr2tyh2vRGFPZM85eItZsC/jM1kNWFBNM+7kIQgDRqjBN7bn/E77dJExITwiZwLCAr
5QBcvhPfnyX0XF9xg07vEEmx0AicLntHpwtEKBRgflugrbZWRFU9aLDpeQOvtMfpfJxr9rA1lhSu
RHOD13txTtKjyfqeK/tY421ocx66ibxT0Mn/psaDaLLy4i/nr1dHYHtZlOox6+/4hYyZeQv2yjsX
tcpiAKsrY1DE/DdlEi/N/g449fgCPXcWhHOGH6JQo5zhuhW6WwJa238bjx2IlFH0HhmbC5zx1yy4
STQBJVZir6W5rX0Rt1006yr6BdvLqgS1T4U6GJtPFOO7q9xtk5qLwV1U1MUJZ03qgfbylGpUqZQF
dL+urnoDMsjYjPFZi/0/D7rXJiIkQ5twUe1J+Rn7E0M6D3flEBdM1i45bQpPDnYcJbD9WLCBCDmL
VryN4MnVfcLhWx0wCVhbL15YQjdnFy4lyUeDaaZP7zqUKxhI1Vs+MOLwuiTujJl8FlOM85rOXFIw
zHQ55rvMwe3CKA0KSXjpZGNVv3OpKHNZcgNH+EpECTZkK529Qn8EAyHw4yD06E9E2DroXp/bnJVr
AzNQq7zecYrBd2ZqDYgIFT3Lr83jsGFSOSaoUCMEaIoW+EvjB87KUuaODaEjbLjbL6k/p/qCK1Pm
gYU4j7/PM6RwD/rPo/iRuJ8Jy21wcjtJ66pDqEJZ4/iKCIqgsGPPfkGA8YlGIlzpcSo+8ZuUm/wh
Q4zn5QTYNMbe2574Gr2KuF+3Xs0BSYGCnRUeplNAdlpWr7s2JNIzo7RXMvdhIjRp0Yt61L10qV+H
k+Jpy6t1kdm5x7kcwifgl91xKc+FkcGkKCoCPvtM5bEJZfbZ0Zu3+4PbkmCB17cvrpVuNT1ebYLv
KbUmTAbD4qufIcPDra0JysTOIufPBtp9FC/YuwxvcSLyua1nLg2cqtk2MfIb3cuYeDwiW3MFtNBh
P4sPNDC9YvQJqUlwaBh62hOIstLfRsZNEIRwGdeXyrpdRxKkxCHN7w0f8yMEoNtQylRr6i+hAyBI
AVRd1/KypzdbcMR6TN1r2eICcM621oqbNC33aLdt7ImjBlN2CiHwwgiFmxJ1YLJVOASOkDj1OSWv
37cglSLTMH66pqg83oKC7S1HR9ShMInrgSWLS+g+YI0+7qY255lsz/zLSE0vqy/lIN6P3123Dz6M
ZGUHb8F/JLBLJdqqi5xAiW408IV/X0pe24FGSTAYfACB0y1H1rySNSMBuY9b95I49k8RuV9/HBfI
Cs6dTf6FnAMRJ8Wd3NGrRnV+4y6mGWnCtovafTgs/+WLeOtkJz6oIsXYQUMNGg0mUSUsIpr0ELg1
WJUE1Nr93p9XDEvI74+U5LLuPZ4CxkOAdRxDOAiGwN7O6yV93/VI1eCGMlgxMliRrRzZ2mc/IIi4
mMvhwhx6+qsbGWjHOhwdI3qUl9PNtfGSAdB8bHeoP1QDbkLPj74n22MpGL0o4OFUwnIJBSHeQJga
Qg/9rdFf0zZLORunf+jo8zf34iWw6Eoh8IFo04FusznhXTQHf/4uw8ilJE4NpEGx2RhUl5zIzS0r
2eQU1PX7DoiOQlCyHixyS/Chv6JkWvvHjrd9K09jbcOsT6pEMHwiRsGTurroksOKxWUCSWbnyErl
k6GeHWHx3Uxa7aj4BMUAjovfQi+g/345fL0O6tVjl/X667JoZNcsZB43oFBif0Tk+vxYhsHJMLFA
2cJFp34E8+T37kdmUIka7iviyc3fdo2HpqMrA2fuAVHr1rSunqSvKuiPACnfzKOjV4xg/n7e4EHL
gK48OaTCHgOuK9IglVAqHwl9npr0l4bqyGfJbXMzZlybObjKw9OCJlDIVemXcSU3Icm84uwxJkyP
Q42dIvpSQZqe3PoqCNMvsAdQR5cl3EoeWyWVZ2Y+Py2AA+/u8Npdpc6hTwRqfEbG8wPBxYawXG+Y
x6Q0sh/6fkEgOmMZX1QjCGRM0dnaKIklmN4b1qDznjyRIjmZpmfxVvUiUpyBNopEqTGlt22uQ26Y
gJuwYVaTx7/MIkBvsMOXJGfcgcCbAyEnxxKoCOL+KLaXezJAq+fMwyZFujDCtMtoCA4AbOdzF/Zn
4vhufiNkVSGzWh7K76qNkTvrzpS+X+GSuLCMSe7PWlztfwcl+aj4BpNzxoPAi+uxU556lTKCOT1T
tHuccek/fxSlhxsHl3MH8dc4tOvkBwhj6tmdfs0Hk9q4q59n2njpHHlcdLvkziMEk3GRjVkJ3ZUT
7bdMe74Hb5aYgnmDdDGS3+AQO5e8peBWi/4sE/HnBRNROsAB6uG5+q9f+bfiqZhbgShxmiKS2g6x
JJxrcuDip5jAUJRSWLzdcG/haTNBlNP1BiLqVNgQjVeHe8TolPZKyyAglg2wIi3th0OickwvztIf
BQAC8ph1LglQpT9L3ycacO/z+AO2Z0neaY8H4LdG6DFUmy/D+TJ1FKk+QJet4rVIzUxxHlN8jUTv
bbJXBz2DmR3UzIzyyLDLIxp+SSJvhlFpPvfJQpcmVGEzI2bUuFqIG1pcf6rsZzztqwTlyKvOmGRc
4HXE6oq9RhEe4+Ul9hjy5KjR0Bccl0LoQ6uDye9tklkPfIAQWqZ3oB4wg8EIvW1BDemXlwnzYb1J
l4ErZIpVuYXT48bmdYM4791lPrC8qyDo6LPHNKOI0dfQal0a9ozJvy9e9motP/Mc1Ff4GlhHqq3d
0GjWIGf5grLbnQrIJRkHdJroxmGdt38AuxwO7vXYBuWC4NoOGm6P6xaxeA8LVwjVCwaDllFnjUkE
F0UpclNzcVLVioRrvvmrG3mFzVa570zQaIr+RDUSmyXX/tPtuuW4QXRQGu306TChPJHq/fP2hopr
9uyLqGlFeSOxFYAfrTRXrx0/Yd+95z1F7Dm56A5r3b1KKA12n3tVoy5DI4onP3LPTPrQi23axy+Y
FSg9aPT+ygF0+idVTCwQrgW0fWibuLZkS3SdL24KOrKIYMB1TQ1mxbvZVghjFO1R/272AVZmeIp0
Ih7PwEEBBd/xpd6TXmrYN+tVjgzfRDQJsslwWaeQxJSVBxyi9i95y/Xeg9iVuYKdqNN3FpCKRpde
9DTn6wiQpBvYgPvDUJ4M5KCuW4+4h9mH8n3RoPjM55087uvbKs934upaCkLF6uis12ne+Q2zUTS4
FeGfz3mxnIMKr2j6PrjMiBOYyItZM6X2cU6AKhvZbV+yzmBaoA3N7wFFsxl34P8DLnPWzyioF6Ai
/TuxoLtfE7cK2gRTOCDRJIqfygvH/0Tq9y+4ySKW3hDH2ezGQb6KaEuTQbvzq4BVp1XR8dcaTwvO
V3WyWbGFq9MYr+OjgTCZvlPln3INW/ZKE5wlxFWu1InDohz4906wvuqS00rCNIOzQ2PMvmubeMw/
KFamtye1F10r2mmPJPGTLgi4F21lT1Pt08aV9L0SjEAB551X2HPU0vHpJVCrNknvYDAvLmYdIjd0
fV5xUIaukKA+jdWVd6zpAY2i0pMf4sgyKAbV3SydKOYRRzk6shxaD+z9l2RhWwCU+mWohjIJrkTg
7o/+Hid8CzDdqOIn0MkUyxLkV/U9DWXPeMHf5gGXSW/zZfTremyJJC4eHiPKSGjlTf6f6B6Heo8n
Kqdqj/WcNfegHpdwSAvlb5QRVCKuawsHwBSstdI40lFISwbLtjD5OJZJCfaJXwG29hJf1WYfrkOv
JMYGTLu7MoeflFB+qLbHgnMHbN5v3e7rw44AllzyY5ZQukrYLGYl4cayvpW4zqi6jLUC2hZsChHS
ZMQu1vTN0yFXdLmMGlTRZT1bsBEre3J4+lC0Dychl0rakj+duc2+W+lMeUc/klCk/GkQMlpBq8oe
m8t5uotCc8aq4BW8Tk9t7hed/NjXRPX5/5HEIDQdndDdwWlsexl8B72kO90xYwWv9GO9vqc0W37Y
I7eLxi82Rpu3ZYC7bvZJpzXeEZLJZadVihlYFtN43l01R87xuG8p4g2YNshryQ/a2QQPgJZrDvmi
44S8CqB1LvEVaa18jPVTkr3QpMlBneNG1818tfndMzAWysbv7p7VW1CF9sK5FnX67UaJhZBy45fp
FzWeKvkOutExEKZqbeXsYI2PvZ+FRwF61xJ8gKTAEaAZbnNXMzPrCQv1BOPyrrqGUvfmyux/ms+P
cWJsqG9YAuq20LLK3n3ictSWbTkw+LxEqVtj75BNCYcdvTdLqoGijB5w9QH9Ht2HlDkF1af+VI/V
f2yVfTw9HWP+Eg8D+Ev+yg7ENzwH8Umq0wPdH7wSM8UxPUOxPZlmmD0XSM1AKqO9cWCNsFIA+hJN
CXsWX3+XnI6Xo4KfiRJ+35ZyYQxr5LNVt2tHaqhmJRhf6zsL3SBBF42mRr+80oP7V8US17W+hnBx
hk3V38kQVysU5IIGshNeR7iZpY2wIWJe2NcXvx30Cou2gs8v0OerFKRgY+YzxFknqQXHQJ8K5HBg
sNQjck/8DtvhR8Pf3PJe30YQGV0tugaflT0+DvpAr0zylxFTjlkq3Y1mdaMHeYazUHsSsebHGXvN
8FweIX3/hYER/RR7lcnXe2+SJyDxWlL3IO+zmD2urCDbiJZGpTL8YUheyTV0CBqrFm/XquLzt+Gh
yu9fu4+AXH08lhgex+bMLtObcMOQmZrr3EIajCwirhj/h0Hrtld4Am7yeIDqaMA1AO5eXCA4Q+zn
O4W9eVAztYLfwWSvLniVFSUuArpLIzaScI7uxZpdy1u/U1zdK6lgPgBGHsU06OKl7zQweI2vX1zQ
I2E+mPiFSKQewP6/w8xi2Evg2tvWCC7njW2cMHES8aMXfOi3esGQQ2I0McTvA1jxeIjlTx7z8LXf
KCj9Xfd3KfPUmdzTnkUSZiwf9bas4LmyWWuq9MfrR1aA9sYAu1yif2yNXagSe2dqTUypNP/PpYtF
qEK2QqX7AgX2IgBIcj4yUe/S4GVxAp3vMiaDvUpS7e2dwWurvX4aumU025Adx91ZQ/gabRANsvZm
Kcwfr5pujVJhX7x3JV9QiZQXOyBQH1H3S6bks48yWbiXuXuBCwTXI0H+gbZJ7p4AZTyBATKMq7iO
O4ekITUcsPQDerC6SQwUoz2AapCq1n8sxEjMmLQD10noxokScXzNWlKFhduWEb24lnoSfRNIthp3
giEcpuIXxEk1CHCr8Sg0zt71+ZkbtYKlnY40Oxp7q7UQkuFe6v1LZXTyGbmCNvaSVCUX7pUyp2qY
u92ByovVKtj2xdkdD28E3R/FvAY4UTOj+ptp8RyeBKGsqUPIiS0tCUyoa/Ke+w3cRYCjj4KdCxG8
rZlVKKRvRlSE7wEFIoc9yqD0WJw3Q0BzKOSZrg2onmgs5nhLkep42MJZwCug3Osda8Iz2eGMtCGv
Q2FIC7e7T1VldZ4xhQZHEJEQSKzWjCHbQl44gZztLAa9octF7HtMGmtRQLwfM4Pu3b/ZPn5nLWfW
Z3A+RJ37Ab/QkwEX7qJIB6RCdKMrkFVe0tng21RFN6OMXuwlL2Dr6BZwCq8zaSFLcVNGWFd0nmNE
YDF3Ld9bg54scRGAwuL6lJDw/z6+/Om+2W9B+FoUodW4XmtNcRSPE5a0fy/a1WtZFUy8ksNcidPs
Qzto5GTotl6ZFI7xH5b76ftaB7SRTulvrTOuddRm3827iHz7COvpQgDIKhA4GuHUiN/UjtLMhQw5
8Ohxcpd2LPe5CNgfZ81+2ksuDrr2r9I+HhLYIUgxLhA61pFBTlG40/SdHi7wG/fQPXBEG4ffErDz
NW1JEQubgpMBgqOHZH9vfJQysZMyJt0SX2m0OWyOLoE3/od4VoHGfzhQzcPJLBrIg1XIKVvsifUL
TiUNIhTiA3VecrBaRCIstk2wvFgrXdJgVK/+cvv/jtFxNPuYO6OxtBBjbUEo1lZvpK3/p26OVU3z
btW7vCjg9nfAkIyFbDE7ALV5XKj0FMo8hOs3YdOtpMHHLbJz6UlZUpbPbyiMJJDnvdsfQWqkA16W
+DIXHDPp1lkxW0cbvzSMquXrr4XT+0I1IurMxBrLFmt9DndZrULiCpSqHSDrdzruWA1YKHpHe8Ww
KVLs8FYMuyQxxIBiW3hEIy02zFbsRrsB/OuwwljK5zeonGCFG2Nrjw7mNx6bukxNTt+wscR1dA4B
R3ghyJmRK0Zm3qcqB7VHdLSmKYuI8uuKO6FrHdO2ekZt5q/E4JAChVN06/L5nxR8x4TrU14BBUq/
WtGP61VozA4z86cGYFrsHPctksg1vcF2yPrQ+wVJbZ/MUkI56qD1K+IbTF/SblpKc4SBKHGtwSZf
3L3eKujczACA5XQRBWtNWi/Yv7lVG21SeHpGy8fOCZsphZmWCAKX5ZE2WvrcHIHtnC1NYNckjxXK
b117xiCDKHcuZj6hbGQWiY0SnR/EbYzey8iNBdpd2j6WPwmzAq46HCTx0Q9DsWW8pPC4fyjzr+4+
/28T1hli2o7Q9JbSZkEfV1QmDRUrgpv4HXknB5hxSq4slEbXDBIY/+YaD0B7h/dbeMkIxbnZvain
+e7byfv3+YR1bqVJgGJiEpsuIb1O/S7weGGKZyDCO/j1DL+SeMJZC1wTMyJW6lYxxOitPTyIdgvs
mMRg2fwqRu7vGIdXtEMEPkeWD3qZAqfnd2EH8uaT6ZbaCh12VeZ66CXen49varKj0r16QMMMsFp3
jBCQ41h8JNBZYIhtIuZF0GdZmdeARWNniPipO0rLD1pXTAZbMPF7Hevtpu3dZCvO3FHndCPi0y5t
IIOBD+q1bG/LuXynnhQLY/PHGMh+vVd77SiHM7GeqhGnt/HP9g94pSrxjnQDxWOjgEyl9crV4Bhn
5dBJgFnWvvqo5Z+Qug9GvgUmgJUEyj8k/i3sAUHZhcFelwK1KMiQxRhMC+j0ZXyR5VF67e/QkJQr
qnAENxEYLEnR44If5UDdziYaOlGU/52iTHb3CdkEVDpVTPR1vYXAoSTh1e0ePvIVDGH1a2eZFukY
m9BqQqA1JcJBWqZsnRQ0TjH8HjciU7AfPSB6kZfbbckf90+bOy9VqBhVQI/VPqkI9OGNjeW0G+Fi
BrXy/9aGsxS9X4qwl9BRMSVCMwMvcpdPJonEZJWxTj51mpqrbo4jBpNO+57fkLlsDcdKvWssXzfE
ouGBO41royppowKkgOjpluaikhuoA9a3xqtyWuaZDJkTyjq+jCbrUOuCuImaFSKawxNpKNQIB6Zp
H513sj6/mY4juR0rFCbVR966hnIdZUZ8zE8aoosstIJNdLCqhlbRY2CKN7zciQbW3FX5QbbcAxuK
Zv6KPVsaDauujKDz9mFX0YgCZFnw5JHpUIw6DeYpYGpg2RDH4+rSxiqF4jBFF1t1Z3j/fAeMzl69
hHnJz5FzXqD1eJj1xTKjoVkR30qJlAxOaFcIdFLBZDAKmu++mZwnCuVHBpwv3h8mISgS6BW23o1+
AnuCbI2w2My4wulO3TuZeyeXWo7WVyYnIbFy4CSIe7DphTU0Zo0D5DXs86wll53/AvRnJb6WJFVk
r7ssQQy7RxeRBPrlphiPBaST+licwFMrCu4IKqf4bc6Ia673YaChc3gyAQBQv1t9XEgd0ThMdAvP
WOuRuZBu/AHGER9IyMUKD98Rmw232bLvFjxg4Bxb2HNxH/iptd3ohJR5SNAHYSDfFDF1zg/mxXbQ
Ob14I7Vh7u8wrsegpCCaDi5kzqoEi2JbDHPXJrjAJrxDmXaz1yBE/rY4PlPKW2tuqwNJIXHKK+mR
/2IgcGixuHGUVInPAokxcd8cqgK/s/B9oVBOrRxVZjiAGNtPetCWsFsxUh+tHuuNL64FXwOEhFly
W7qWZcvmy3XKUXmBZLm6/vUBXcgbM01KhI5CLaAXf9OetXgUf/OFZQWi9BZx70Xg0ifMAUuBbuoe
E7e36VK5o0Wm/L5IyzQ+uDWf3zHqthYBLjbLgvH4/4bX8nRsVUY0uTxYUwb7weLFCR+heQgqssor
pz/IBnO8Bv21PcpDU3I2hZjY2RG39vOOJWT5lcaEGT+pMEkFLx7b4soiAk6plQ6NqNemneOJNNWf
UgyqNuak0q53UqFBpw5YkN19IT9cwMCGduO+UVkemGUFg5GcW6JEfPdp/K/K92tomOGBCFL+1g0I
1KguQ228Ril/+cMopcEQsF9819d+ExmfrUb6rUEpgQ+NKHXQw2YhKXff6JpyDZO9CwqQ1vcxZQJr
b1F3z93fTBXDdDIoS49LbiKj3+udEUIunqzkrxbWuPX199K/6gUjqWka2Yv7D0uYIIOuhDb6Yi3k
rZiCyWSGnbOff1KIvb04C02/IaCqkyiQ0oA2FXNGRSI+091NKeVY6OOXh3sGhm1HelgoyHWYz1XU
+R0fzyaJDb+550o03Yj1yq8BGtPdLpvZGaYIK49pPiDY/0cSHeZaMTSij8sVRg3vewEAnZM7G39P
TCeNmnGhEvo7l8TGK0JLU6hF0AXvqwJaw+RdJ2jJgSwxzkZio1rBkBCEfIk7dWSM8LfRlBGWtP2A
s3yQzYAPYLr4C5fzeKbYM9oRPtPiYuHSVIfKnxl7uSXxRfj9jYa1VOukjjwnnDCjfGEvJuXswKUD
X6WBpIZHTpb4SyJ+1HMtyP4zKRvtw8WyuoRQIYpuN4KQVTSEjvMU3Vqo634MqSVIs8bhRtZCYTab
9V9UPVUECEjEjprVcthaG5nIRLd+DZWreEV6tfFGtr/sC5pC6+9UI712Qb/d/f/+6f1KRzzsMPtg
zqfathceEx1WkayUt64MBaNKTX6837dF4JrIosboOtDWBMkRYmVESTsKMDhKRzvFSi8dViBBv1Vk
V0T0SdrywWmfgizb1G+8LwlXCCzNWVgdTkwODOb21jGKO7uD6sNX3f50YT3mPhbS3bIVEBOhlvjB
tTzZ+FIc7MpHYnx0nWGV36Uv4OMUXzCr1suJBX9ZVNf5Mh/E0Mica86T9v7CTiap/Bk73o6kIBjg
4MNiW4CvustILeeCBhYO49TY0NuRyB4/XhPFqd3vNOnSg7Y6ROc90F65XJl11e+mDCZ0w442sREi
jidjZZtf0rqlmtY44lc36p7oZnt8I/fPEjZr7Dj8ALM+t31RmvnDXtcHcrju7/ZIPnDTK8jtjYoG
SfGIh3hmAMdCSbOlnF4EWp/2lAbKjAIcVP5U7U6d/AcrisSrbUGi5sWoJeD/k+bc6nE7xeKLGeVi
4RXZN+ZzDm07EX8S+zG+E3+D3wSvwIC6PqCbiCncae3C3IywjFGYKGEtiV3SCreOvL5DOkFXbIBU
YmEs8eia0JsHWMAl41zVrqA7uk0NfdR2TZcjG011Gihs+CXorKKEWSrsakJVLAG8TJw5tYcPF8lf
HYql1cvgyGY6gNDfLJgWm8S8e7A4FPtdsm1P4K2X64GoAFhGriZev0X2yFbycvADxReJK/v79euf
gZNH3O3o8ig2DEF7pLv2a6StLvRelowVPaXUiiJ+oKkZf1/+M8Jx+MT150coZoGbkomPukCCUQJN
nsP0yOCz35glCZECqla8QlwB2BaSd06cp5otUSXUQWK68NFWghYtCn0Kk0FqqPP27CoHoczCLA5/
pLXkxJjoLjqNVbbmvVaWBvMWUz1HABh9hQx3CPmSauCcXLQbn+P5mIVhGQYsRqANw5o6UPahqCKI
JZOy2EcqbI5fRLbseseLSxVMeU03p7DmZMhP+z25fWAKHJt2hNUnzkZv37QtwIfxvwasTjh8N7ax
nXp0HPIm0Hse8L49S39AL6qQ/YjTqv/d8aqNnLx+s4CPIFZmqXnFJ5+4LAJcrOPno5zHuGVwufQB
+bm41O6pdBK7hHP4jtPf1FiGSH/yD0SjGm8/4WA8upfhDo6NeCgG0viw/WPpY8LWw3kCtxu/uWrh
RkwNdEa1hTB5TYrdN97TDxznEORT4KevpWVAYAB89BX4Svw4oAc8G6rt3mA6U9e3bJ4Az+/tBNl1
txbyxO0lddw1LV5Yr5rqVDqQ55LmC6aFv2lFYWEkqm0nKC+04+biDlRDUHHqZK8i6Epzz2W/FHvI
5OvL4y5gHheqheKOnKuP6tk6mTgjGsvDK3NdxBh0FU4Ya3y4aR5Psxzu+2AL1CoxpB3gLrA9obOd
4sz1p+Sj7DFndycuM29BFr40yAmcSnkW+c2+wjhdZEffI+fbDHGyyadiBNSh47nyaTP1Dgr1Wp4w
5QTfKZnGog2Ze3nqSfe+PoING8zKOP6Gg2BQbOP1LmqOI5Fea5t7ld68WqRcmnQK0PhcCGU7qNmS
5lEB+UR83x+PyzT/8BZlGcpK11QtX6tO1Forj9hCpagJjR2h8V32S8pzcC0SoeL20d+zk7iLcjzL
u4rDlpl6aCh6FznXs3vklTV0mrt4/bb/iHsD+HFYfKq4MP0YqSe50mzk1wfolsmXqWlHrOYkRqTB
SCEQSbMvYoXi/xATWm/c0D0UUnvLzh79/yqLUbZrC5Lqzs5YfKzJtNseZFWGkVuP+qJFnqFVS5g/
lhM60sw8Yn4IDMZG/f/Bivsl8MAwUM3VDADKvw2oDjpuNb66viM5H6v0fZUd1Edx4SE0I4iFGCGj
mezRal5TyIBvZrWY1p1TQ29BCFqxy+Hc1ZdNsqrtxi3BmnIfZku1SupKUKS7NDNnDQtag0uzWiGG
eseFVE+hDM8OwOcHkgVpHcXw6TgBjQv6L4M6GVQaSjsN4pYUK+Yr3BadD0RzFVhExILbht3I7s7R
ylCfpRo0kTwz/WTEu0QV23uQ4oAFV5YFQI6rpcsUdzLZYaMtHQ0Qjk1pZhDGaHpwR0+Ch/64/T0c
XB+WdPzqRzMOLknRvz323GBbnV+/nEKE/883TPpBlqqKh4vZPKyFZLspTOQuJyPEY4sBWl3WCbZs
jUZMBJ5vOZ2v1seuL+Az79/xGdhR7tPAcfjpyq4fTwtR2Suk8yfNTXhawyKnW9HkPxol9kGbven9
9XzGj8Hj264JPs+h7BvOVhA15iMPHc7K3yZ1EZT9dJq4kdz2VehmUtyAlxKhTXjayInqJCceHRqT
meSDERZLz1gQYYLNPxPNS/45nZ55hat+EH7tDpd7jKd6/aR5saSEJTNDhipTFsJpk/SuZQGjTsoL
JG90aIWXYDZ/cQkRpk0ufKAm5Gvu/sHdHAvv4Z1hotP7OcpbTdne4zaxgXlfUGitACk4fHYidb98
GgvEDRx2Eb54chnqV0NgTq4C4chsgID7COuS3LMYAjI7cq+CRBKiYfzJ3VhpTUPXcBnrFfxNshMG
t9fWiLz7wPBj/HTYDadsmjSqoBdC/AI6MQsJa8yYUfEcK5Y6IWagYz2fRlxRx+S1L631+ffeUb6A
2Aua8ourJpIHSWxRoCCe9DWzLh/6i9KdgIa//TmJvQg8pWwHU06sQOJN7Yutu5DNAiIodKbKYJqx
rd5ja9gJ0CtNDQTOuf03Fzt9lGUCJSHPBjnBx2wh7oraAKsch8mJwabUbnUr00M/+fQ4z0YlU+Ur
NkxlCgSvZB6ZGTDsJCVp3f6mxEqdoE9N6CL3qIf6hYPZfs93tFlqmb/8A2ortdXj9GvaOraCXzWo
O7TW3DvBAbhO/HHFnl1S9ZCgcwdbt/LDowqGIt8KZPkbTMznNvBDs+yN2b1zBZHI+0ZsLClHvS1G
EdJ2A5Mj8tgXiExA/kCYGCMg0XNeU9fzR0qH7rsaOGNG6uVAYl+Exgo0y1MOzqsCPR14xzOE3F8h
/7Irli6Zk3Lb4VXHzpINqRR5wr9DMnvEDrmd4qRBtV4NURq+m6yRIZr1yeEwQS2t/OF5ju5Owprl
D7h8RusAg7ohWvs5IG/aAU/G3flKrhHjhPb4nf9j+ikBfNPbJur6P7vqtYLGG3N4rc28BUcQ2AwQ
LOGRbvybGuhQRVU1DbvdEuLSf6ujjzhQbFYBJkVQ2EHFmdNADY46yP8fTrTd67x9nuUOvtx7bwA+
pHVyPs0RnZ0+eC4YDma+WsomRmfoKU7fmvcHY9g0wLrjJAZpQNxU6j9fOWnBotQPZvMKVlKKBtSL
aqj+LlJuNigFJUp8/q2IMAWxeApds4OkxZH34G8inIwiiWPJpq3v+vgyTT6+55fiXVlOrcb4B/jJ
ykJ3fwVzJD8fenOi6HKhojW1Lhaw0D1Vpi4tMnfWSnTXt96HKnia0A+sXb7KzHJigx+b/nRJ+04h
/aKFCsV/m+UhtWU66V2xV/Gw6lv6lWYR5Mbbwcd91KWqtpFwU24MK6vVXoYfmlimFRItRDslequF
GxxddXPr5zMC27pR/LU7ojWsBe9014udEcaodqtYYXE29heqkGecQFIxYpkFfwIAaCPiD+xy5tWt
boIuYQTJcakwAVFAPuGv3yjv2gCdrOv/kbwiCoCHC2C/BxrBmQ8TKYihgqt39omyTG3gbHKxmKJ0
a7Yp5E4HbPR9V4MLajSJn9+w/++UV4K+2XuNrzU1zeqcX4xem1FMSkaZ5Zm/u12At0eSUSdyZNrT
xq/7wXii3bBcUaIwQQ+92g1AFR8jZ6io2lRYxi/QkMsqgsIIeTyZCGNXf6QO5qkw11nkA5rkgRkP
js2o4JoQ/XAtvRJ4D9XE1pU6SulUZ+9RzToS54eEDYtbvx9cJwXF9Fqf9sDLtu+XgpNEb7geMpc5
9glHws4rcy+8Ioint7My9BBY+hObP5YN29mEwFQvEzaZm6wdoC8gaL7hM7/Ur2OQMECY/8XHRrdq
ARDh1rQL+jz/of9pCXk0D7JRLmxvTm90E6Z2mur7ALLmwYe2ReRy9YBTcZC7ML/MwHwYjs0cufnD
7Ot82mivwJFlHujTJTwY59b0der9+jZLy9Z8DMbO01l/pIxIasHlRJAvEjInRWODDjxHtpL/+/GJ
dtMHb107dHbX42x6TainZPlZVHFEAwwbigTE8GzmT1RgYqJze7KM/9ejT9Vy/UTEeXEbuzRkXyap
GOGvnO/tv6ckSeeAP8Qm+onrhucEP/PTQFoyTQZ7a/F6KMA9FjCn54P9V+DurgrMMIDCkG2BzHXZ
JvkTmtVswq4eqJSK3K2EBhV69bnrm/tEr/b/fGGxnwgu21tPQOE91ht+lD6mXqaL4YgdmXhCiqfe
bQUsyzRh8p+Wr5USrHio281aGg2phY8YH+kFZzTBYDUuZeSuhBn22k3VAqxKkY/PYRSEnOm+5qrS
3iL+DJ3FiIldWowj+tHnOKsfPdq8G8m4GtKjj5t0dacb5Ky8cBqhF+V8Cg05UhfcOXozvK3D+DVC
HxSYbCEVrz9lunWgGT2cRHYu83lZwX8kbcozwov9UOhJVqM5Zs8wTKPOKLCkRNdj54yZNupTwONE
RlX77sivAKLw7slHTLDWtz7zATVJHphdVhgXrvRdPlGq/oOeSRfbgH8VcSSNA8U7WxplAsxEQcKV
UH3uFRI/Vux1+i3Pgk+GKdlUphjBpMaHqwOOv/akU5LVxpPlWoaLq9VDgkacDeNk8RVkw0GsHur6
YhJ/FuGyGAJe18pzI1/5gvQRZgnpT1jdvEGBfXTHUHip/j7AHgr+dzA5O2dVhBz+Kzan/jW0g8o5
QVfe83Bw+bsgiorYUg2qYfTrekkr6/fu77eqWYh3Djj8UrNF15DkauGku/5ZSyZzQwleKBLsK4TY
dz0Ny7BHWaM9cMW52lctB89fSHK/meYG8kJnA4c8HcqEmb0j1wwbZPj9XGkvyI3dHKm7rO5EFMJG
oibDyGT95UeE5KbEYJ5wkyQf36s9bj0A9zwIyJiKoyiieQLDCZdLd6vujU4lmsyOvSlvhuNoTxZw
R8sCgVwv6xF9EyW5q9GSNDAO6bEcC/DjT1X7GuZGW7vK/4uaN1qMTDk1jeNBVOnYuQ/wOArSSg9K
PhhSl0zRAgd7SSkQQfIQgsE63Jiuhh488PB/y5XNMQc6wJzqi28DMJiB/P4uXw4gByspimILFm7Q
o/thMf/A/TMliJBV2O6Y1TOJm+L6OrLRltDrsUeNHf6bXxYmU1aiE4XMguuB+6nivt5eGV/CJTZR
LM0LHiPPnjpmJbHlwZja7XWgGdzekhMzWeykdC9zvkmJ6yH+sArH4xcj11deCuBUulWr0ox5+ut8
yAfCkWf+2FRi1xJApKXOn16HNTFMp+8Vu3Q7ja37XBJoTil3de/TWHXks22dG2kXbddxot9cVU6m
8fFBwrUtHO+0yy1agAkg2zUQaVlmVWBEB8B23hmiGo9iKmle1sQLFBVprfgV5NfAuFE4/f5lhQ2I
g9t/iNHlwVa7+PIHbyElzel3bbSOLQ8W6eAOiRNgomIM3Z8D9erqPB7dcnLz5s/dGvnSLtdPp4vq
rk+nvRVs33TzUB/7wLY8svWcn8JkxcF+sP/3vItSs+xhVCuIlBFuLkECAWINg0UDamcPmGzLT63Z
jG8tsedyyOTIOkPYERgeftyAjtO2GtNMbyUlKjof2OJbTc+Zd0j8IrEKsjU8OgUTAxKb+j6uX6x+
GudWZ7S46/7O6QPubXtNqGOxkKQmwb9vfK7RfB8zNA87nxv+EFNrtkd1lDlnJ+LsWZPusNEd2BAH
mgJgGjxbm0twpmR2UJK109/8ez/u5UX8FGFdUbIUcvkINKSnvq7vrDzw1wS93uT3cMmkfs0ZXR3Z
N+QooAODjHaq7VCc2+RUtPyqr9jyaSv4usObV0e95KqZv9ohpkp9LAEZ/uhFAH4OffiG+3Dj5OwB
o+buRNXnjE+aAWzcNjfaxcq19p3gu3ELTXTRcxnX7P/X8E2+IUKWHoFy04GzRIV3X3axLRyaf2Tj
gPlYwlBmi+Tg2wVQaygsygEBGUvq1CqpbBLN7k1cQjYZWj0lpnFkccUBbq0tJ4IUsfYpnqxx0t7G
gDA+qBZs7lFP0l4GSXHomtZmzsbepHu1DfpGpq6U7zbONBO0jKN2t5YNrPN7wQplZGMo5F7+U6aU
dJWgJNbDdr0P+cI+grYaPlZHUYi8vFrG0lPu8VCMe/732G/ZM6n0YpO7aqQ0VBGCZ7+hJGkwM/7B
V+KvRjgzwDkVyCprITIm4C3Q1exvm/LEBqNbuAB2Fggno8Q5nvHtgODIKiY89/5+SWSt8sO5R6nd
PKOgs4g7jxtH4OhRM/9mHelGKvVadxVw1CaiyT520MqxCyRw+qIL0W23CrF1u0EQQRpXCHo1+3Yl
G3etxOeOcUxUyp1pLVGRZEYEYE/A+Cq8AhNcYdDK++YVXeWTe/ju3y5v8kwhn1I2l2WF+5hzA1c2
OzMud9ZrgcEd4IFI2Exhw7D8ADloYXW65wAcBCvl9UE0ReDosPhx2EbY6fS6W8XSofCPRD1k9j1w
xAdXxMy3aVF+fCNMNvaCKExtjhbBsQqk0C5NYyTizNfox8z3jtrhFaodo6dNXvS/IM/OENL4lfl1
th38PkVjxCLP7A9NqcavwsqmdVJIICL0+vs+cua6UJ0Y7muSNA8C/LonqZZlhCOBsH8Skx9pvzQX
IHRJEswqaTJr/xRyV2ZMy4uYBuPA+nQEy/AmGY2OEQ8UK1z2wVeNRkAaV0lSD+xF7ut/MGGlgtlH
VqzgYfi83koBBd6uoDEbH//QJI0yWUxErkJDN9lNrFoQLEEBteSPIHWxJD3/SY8HRC9ubxD5dUCF
JR6W3fttUOZ2yRdQ0J20Sn++EPZbP1w5kmGNmXmhdqL+Wfno3ODgUjjnQjTcUH47op3l2sCq9RWm
0LV3xpOqJ35fjWnUv4AwTYgijH4vjyHMOa2qOjlI1v4a+TWhkc9VWlO2jyI64Byem+mk6Xu/rTLV
fqF9XaqLDlyTA0QriMvHrsVsSV0YdqvdCXjV7xaVL7gYyZAdtNc1EU9meAIVNXDyAGeLOXLS0ODs
4etxkKYcccTveh7Cr3EvLRYZHoDATkHUAvgLBwFeQF27uWE5D5OoL7It1WwDL9USF0FTHHq250u8
2nbv+N6pRlJLxN7eOiFrvt1ZEj0VdpZG6l+vDNkBr+ugGW+5cSxmrXO2mOgiVBzk6rx8Eb/Ih1dE
BFzd2baltSQJajZik6G9D5i87uF9dS9in7AtSTYGgMtLzJZBUZqhqHoe4DNbAG2XLi3TYX41dUVJ
d45oR5GpHKvg2oQXKZKvNNPbBsasLWyp/MjlwtAdYmrGBF3lyMvAXZuZRs7bMexFEAd9m/HQFyue
zS2WJaVY1wk5nsNDtLOoMovk+6PUqA0Dc2ClIidKXx4nwOhQWQ923ymtPw0TwyDJUekdamJIT/zd
lAFGGk9QdA0uYWAgijOCzEdCgBvAG4kC/vTSNgLehWAz27dMkx0lCiSpNCd7ROMyH+X5Srk36ZNw
Mdl8yQpIacmBUsDr/RvaAOmMMHYkMLakWxJ1cgcXOKFFC8HP7aMjdTfytg3PzRhjK/4OCkUCKH7Y
AjiMU7cmQMHAeImp/0mkv9KouLt2d7Y+QnXui/KwicOumJW4q+ESzk9YAIxiS2rVwOr5nF5ITE30
qypeNXTqjwh9iE6qwkXz3seRuz9xxkMy/OsLTks3qX1IgGN5tHBkv+J1r9dDx62RZVkgFewIq6NF
zMNUNAJ0VwMRYHXiksBH8zQcxoiFfbYItA5hC8SStV+12HbmNPNh+snTuhRN6VDGlSRMD38eu7gY
/ftjoqnhOI3E8me+0yRDyxbwOlsF7m04SchHv2VzECsPdShe+JEMAAELofn7ElnVAcw9hA+5qhvT
JJSZAvoYH+HiV9BTOTuNeWyeC14UApBWgqQrwTTIwEkJrRuvAhKHaKAIl3BFdRhGgBM08S4Q6ECN
7Dpmjk8PJc52zKEvKas8Hlpr6FA6STPWDlOIAL/WLuOOKZ1JSxgH8+kvBQmg2rBiHz1u2jqnngH9
stEq6HzsE/7uUh4bD4bBbRBwXXnox5TRKxGGAFLyR6ETBD5OH2gyhPcXqrSB5t/VQDDl1Y7b+3GB
MCbeY4ZA6eZXxjOkRwnPaYF6xmQtV6zlEl1FMexBgtooGH/jQ+aZbNzOJZWK5QGl5O1H9/38q7bf
lbtT0dsnTrmKgtw4W1qpYH8VF823W1sHx0bjhtUeezpGX8CtctAveCbfs44wiFI1Wq8QTbJLtk2n
TWYxY/mJBGH4KFWkJXvzvFQoOEEUnX6wNXFoFTWdZxKH2nSGNZiKmql8W8wDRIa6zuQmzb/PLw6Q
hs/mQVDl3Wc+ySM1qTQBUh4xlFfAckNgwkXSK9wDGivvsFXK0o5NMYzcZfghW5WIaz3BmX5u/uvg
r5cJ3PMarEVohK8Zoguo2cET8uWx2G42SrcTSHbGhw/o9qL8xaeKTwnwIaXiisSRjT4BDENOwdK6
WuhGvxP3fMNQljWsGaK3Iyu55IbhxwKO5kehQcWqyitAFAM0Px+jkgEL9o3ETBtjrQbmz7fxgqF6
YxLNfcDuuZHjS2Obn1pya1psw6DE/L802ARJa+lQlkocgFAfBYrYEnFIJ7Uh+MSzNTIIM16KWDEj
BNcFmlgnRT9Du9zQDA2gwQFsLOR6bNB6U8GIRtoWwXUvEv6U+BOBYQ8xAB2XY9hQvANSbMRrWBsa
eKOCgiFGi2Mu3mwIIdUnpil5fG9xJOZYCvI4jRj8Tz9YywcJHJrXVxGdweVIuFiajswpC3cPJFAJ
JK+/JW/th8pXU20jsJhfPrpqSuc4zlIL2iNx0ee30cBuBmBB6agxS4xSqwjzMl9B6oDK7HEX4Er+
pP+QCd1+pnKfy2IEx/EVQ4mZJuWiLkwX1/jjN9zyr2wAtQKLQo2wP8v2mYykYnG4d0HZjeUWl4+x
/FxliWOnyghDZn5eDiG/GTJlFblZ9vsOnyUjOx1G3jWhKRPFgqKXZl7RQjKw9Hw5hXeRqwz1lraj
pUcHK0twW9hhAkDCyif3p4j8MLxoksFscKL38KLAjqY1fLSUA5ZI4WAgzLYWR8GxTFgTSQR8n2g4
wpW23W16/SKJZtG3GqnlU4K44BU4VxtUGSDpLStKLoKzERGfSVzW+tn26O+Wn4VUTnzwg+MyHePE
tTHVnH+o/3g+rFo+clzdDIM72UO9knX91C7v1gOAl8EYGl2+YGf3mbpMkuPm0PG59B+EhE1gFvzk
CymJ3HGPSm1LyPHB3MKSD91X0WNHXKY3kMUOZgUcfQllYYYnGlEg974o5AfHJNCJ8KE27KoPHxHi
e6zBHOmQL+nznZHnIJn4S4Ea3HV3S9nOdAqil7L0wAwi9RRlB7D+XOl6qswwPRlO3rT9opeFeVvX
Ak8bJQ3KyUHiaZhYa5wxJcmSpob7uJ8EApNzX6TvotyxDkZNqIJM4K1OVeEo+SSbTzw1Yz8Vahsx
2wR2U36GvyoEpyuyxaoW0qHgbuo4PX5zw+ic8MQhJVkOHBdDsxy2euxSTiLVoYDe+5sZFwj+0wNw
agnTJUbmnrn1BXOtxdWiY3vXPvqHVm+wTpLvHUHS5RVrDFi9ku4rRlyTmmdmfXs2RfERRZAgzXmT
pOy/GREuj2AjAdwKl5bJ7YTwvfZEek1+5ckB09Io5REwfwbfZQM83UV823denqMv0VUyJAvRIezd
c1sCkBUsEloZDJfxSz9faRzfrCsJpeQKBARCSNx+XTRnfVJFIQ6KpNM05cTZ9lq0LF0W1OfKtkF7
H3cgRa/fDaiSupG4AqTUMfHFbHD9qQQQQr3cbTapheC8scZZmcyf/3H6AynYOuSk/gpJXvTTRbh9
BJNOP6LUYb8FbpE5Klqbom6qf3tWQrC1u2v51ffyUOz1r1A3hOSEbRkuVGHcBS/VFl2HNmGBOwbI
p+wWlM5PZL9RTftX5vg7OqI/UPS3z0UgskrSgpkVj9wA7HCiNaDedKw5vAuKgN2IXuDwYr0y2+lw
qvgJaH2HgjwF8qjvKAF1ZMCycON+22PNSIk5aKLFcdLE9qbufHV7rVV3F6QNEjUo0GgeSnFZL08i
zuZHg2IYuVbcdCDt7fKsE9YTzVdkY30QfeQ2FtCKSY8uNZGv6Ty4aLwo/w03vkn+TajfOf+Rq6NS
MeR2sYl48er5cikadS7xpiZ7qw1kq8GDnlrm27sWIfbCzXKn1dibRvr1KPaGV1xoliUVTE5+Awjy
KuIT4a1h1Wps6osRUdAiAixC53Fkfvq0q/aurEtbWcaGSQVJ8v2+CPqaqS6r8/1ka+l60ChlK1gA
Bd+TuY6fibDMxctwzrsWPEraM8GFEoWoiSKoTmQrw1jJcazJdUfP7sdffBhqzPkkp/Npk3gCAPvo
4DkD204wlJcUbesQNXxSitODQTCYKI7GjrRvYCSzmaWvfGC3jmFPphr3MgPekxWLw+5nY0NxX4+S
5go5T1TfBT9AxmLy8A5Y4tdEbk90m0oCPLETnnJaXc+ivBrlaQxajOZKIE1DnM+Xf/xaalFbdIwl
LPA5xVOJTdyb22SVSitrwdIPIWMCqWUEalhjwVzXOksJuYPWUkM27v/u/+BptLh89oYEURm3ePjo
mA/C5DCpIxG3yQmjwQ8myfQePMT5TBocmApfEuO370A4KIhyRcc+LjJR4FLJwfc4B19FnAD9dAnM
gLwfgxx+qnHv2sU90+Q1SQDCw07f+SSM9vg3SOMHz01qMK9R8e+TE6yEvYN8M3lHvS/TzseJXOic
unR4bpr6lM6oBP3oBYz94K9cdzC7xYBV19E/ySP0o/6znsMBxAJFCKIdRwTgRfKsW2HzadHG5Hgx
vij9QCYxJ5VNqI8TWbDRBSbOi7fkJz4+CevxJYK6opYMD6m5dI1GIZ5A8GDCBzw3wk2OIKWTJSwe
bbJ3UFoiF5UVGTKcfcGuojYcf/vsfd1l0cIvlInl0Q7jAJ9E36l4WutAOR+Pe794N2vxP74VblNZ
bjWuSLvf7F58yivwYjb2O4PSS7m+joTA/Ssgbt8qa6S6yCIoUok0JDYH6N9m7Xl2GaRinBHKzml+
ptTo+/1ZE2VP5Ygqq/NoSEal+TpSvCq8cz2JulUbzaAYwpuEzjt8HTcNt+EV8s6Yc781XiNkxKJe
iT6+daPaSIsPSz0kFc9+4wxp/ACUOhFIlFQ5q9oEyZU767Q4XMSJNHXtDPaCTmu1k3LEjyFGVVHV
qvk4WU4qAC3vc2rRp4u9bXA5C6nwxMqrJOcjiBacOkhS+WYY+ChVLCquNykvhrq6wktmlVtcFa1+
EoOZNOTa558+oAJdYc71/qkMEWjfhG3DVXrpjCMetu//zje24bvkxSYSt88KFedXuin+WZ/6GPVB
87SYZKftt9n14KW3difMofz8jwMPQXA9glql3Ny6poNa2PdQWgHrjB9rB36lmx8KxIBUutjg322n
RlxnnMNxTmB6K8HTf4aE0WZx9Rf//681t7mTIOag+mK9w9VWVkL7ws52wZggHFVBrG7k7JDspxkq
tVNijG1tbZsTIugSfveZq3oYrUVAkV1pUKCR7+Z1+cN7pqhCDXrpn7giHDe5iLR2l/d8W1UgpOz7
LxTh0UxtW8zFZx1DxEqICF0svVwcWZxD/VthqibRXsufcjaLk0KGcllXHpRNKnRKAgjeS+C/sujl
5PGRZTc+aaVvhmWtkgZvUB+rhPKV4pwPr3RAbeJCcoElaljIHvK7/DvqEK4O5cFgAqPnY9CZgUEF
bntFSxmWAvy40BuWuXvWXEKVvZdm1TlhwzEaXIt/YAzTfTUd5d1vIREDFw87LJnBpm3h8D+1qiIk
x9+qx5WCdTM+4TFxktEr2FohHr1qqyA+D6T/hhA0g7/HRoNHW20UNQylHmG2k0D/vw8aBVTuYVPq
rGQ3BaisIGQknOtC36kKEMqYQnAFEdNQdF9X8gT/Yy6H+BmBpl6JzHucvSCUqSxrrv3mWollnLPw
uURjg75NoC7zwCz91aui7ZDqhaqA5a9qoCAmpzZ5Y7rWFAuDL2Bd9nIBFjtERUrFbZsO7dSl+IY0
X63HBv7YE/aG/umetL6x+feDgY9ITDb6iTGlOfmBMhw3zOMQCySsdhn3Ru4r9rz5rsUFwPUJHrP2
zH/gpvMwI0B8xGDx6PQdXVzqA0CYkbqXyQs6mVvg0j1UyhGKtwhcxOx/rveydX02bTwQX6HBv67h
Qlhjm29Wl22OFeQR8nLjoZ7Cca3BqW5cBs+PVyd16cQpi3t2y8LWkhvZxnuoSzAZ0yOBcniLM6Nv
3cj1MP1b1UBocYyNPr8gy3QlR7U6LJcfYVbHtu1DXTPsU6f81AFXZisvbsHrNMDMdgGMRKq6EBR/
Ujs1YdPGF159dVtFew+O2GRi47LsEFCSxI5E1fWNvj0GIrsP740wJ0RlVUjpnkgD3dJcIuaPeD+E
L/f1gq8OR/NleEtM08F9t9NnOgKorER1PNTFSTcG9H1e76zV13GScbsDpoUyyPgJY1A+TJYv2xGQ
qyM092om2o80fwOoOqDhjmDYLq3aNtaiV5iHCQGvZz94MPx2hStLqXwbBAPkvw1IOloAD2g9fTU+
kL51Q2DBJRn3LHnG7FOYvhmjYP8jR1isJkLSmsLcDnVUULNw5n7LsxqKJt39+ExFzizMh01GGYUB
CxM10HYRAxalSMul6oD0O00IrfJo+f6KSbwfNvTS27zrT3G7GMXCRq6ext5L1pBzzAtFajHgiA6h
1XM9BfwRNthT+v0e58eTd1/Gd97MIT8LwYTyUvQGRgiSq6uNpVIbNY/iml6u81g0keE8k8lCjoyc
V2A608Df4Ps+zCec+IWYcCUIR6aP66CZPfy+Cnj1F4vC9HrO13u5agXHOo14g9R6ikMjXQp4JXfD
rfXYCKbFnsBgGoI3uu0W0vGDxrwMWM0pOeT7IobEVb0qZOE03Zb1gglq+H/WnM1PUWsiF/RU3Wqr
7OzMbZKmoRpqgRvv+OMqoSeK0MVOfJbRzThLJv4AGodGXvsWL4as77cssRHuTVDi4TUuVAm4gHF+
c4Zsb2PPOBZu8YB4aReRVhlMUVTvvHmsuGoWWKgA/ZzY/kGUw2mJnNmFlBGqW3WYvNiVW4ZSk6Ax
jhjlrIr2mr4ar5aJlx/ztANkSuvByy6n8Dbs2AVRW6Jf/bkqzwWyWwmR0sbW/uqk47bemialyCFo
zrQcA0doKWGzGF6Zx1cssgtzgbHQvfhxhwEomfUavyc/z+10LLqLi2C90ve4857g74p3V0wt51KG
pSUts4oPmRefAE1VibP0i+Rvx/kzEGRLwkYV75nBjLe5fap8iuCKsRmBjqS8J186LV55sVXW4+fZ
vCtp2lFl4CXunBW7t7oWqWWAzyZUb8bp9w+l8mqWH78XCUyzsfSkq5+khgiJ9VKCBQvka40tYGzY
vrUluLUz7Vz401a3Q81ITrfUgu4ItS2xK/bmUuuUEjwoldemfBlmeydtDB5HHee72XE90VW7pIek
MfhGE6OtsOt+tNVwslq6QJW8zWTioq67nn4cnpSHyZNLPk8TQ+Ihp/G86/+bysJB5fgvd1XNcgVY
Is8oZDqY24vljCSKzYPSdpPmBFmJ/owx1eR4TOqa6OnkESw/spmMPxF1iJwTzL/Ob0f8OpCqHuYk
locGRajdCPDUYZKZXHsKo5GLoBEa+mANtWbC2zfryI1tWR87O8wZBKlEVwoh5n895Dx6oLDjq6Xx
FWLU2HFOrgaxWgmXRRZHoag93YtzAeNZ+ml1QUxFwk2I1rUGSwEHjYE/if7sglIbjU0mNdEQTwEQ
+EZM3SUcspDjJy6dz/CCJaeL76sWqhLyGn4Q/AnL19q02ah+gmavBD45qyHCC8/m+mth7vrAGR8R
3ItzYA8/jDnTTOIAz8xnbsxi7Ynk2/mBH0c8Nc1jt0IwE5JNksI18WLVJztvZ8sJszaHMQKjE8VJ
z07rszHMSMaSB0YGVT+ev74CoOtK/BYwy6WLnuYgiawfisSIis2kseEF1r0w/o6QguqTd6g2WSl2
cU6fVsm4Y9BSvvnNAED7AJOLAWNVnPHezNtORXC5XOyD+sLjfcWfSvOrXrK7WJl9Y2euUUkKJTye
CpPFLpVA2a8A5fNINABgoSur3JrvzuudCeTMdNw4+xpccoS8fB/ugXyrii2fbU/f3E21rhUDAsFh
+qD4fNAQ22BT46MVQwq2fZ/p3J4hjlX4SGtsE5rA3fV85Lu3MgHn6zalc/1J7W2hwNJj3fAuJLFP
czYbH2MgozJqSmRkU8RXPyrnkrZJQVE6QDGdecF/PR6H9THiT4BjihB8XO1PoIW8x/Zy7z3Z94dD
5dohas5HK6jQqx9uF7SNdFXjxWoNjSmpmoawF0N3dDD509/DPrQewuWmne7Dfr+8+NSVZBwLnq9N
b8kpXn9WZ/QIQtYzSgmb5WviSonpWQbYkY4KFEX6S/KbBOihR324orVWzRX0n25Gd1cdBfhweyhc
4UaURmKHhAkCvpGYCqPDXh1p2v/AphYiOQjkyZMfFsOYMz3dCUQa9RO9xb/yrMbQcS4YDfC4mEtF
LaIr2cm8ZXZJQ3QF/vNVeZu4yaEH8eCyTv3q2XpIKabYkCdbYAg+zl1gk6OMLCSLBLG/hholTDK/
EOAge8aaoObkay0dsVrzSoWoPt08i9x3eOE8Bt9CNzDVWEw+X+VFam/BdhEgz8qGvNgm8Wfgi8Hk
pbFElViubkMpPcpOr6UijXefRh4n3ELKusoYOh+qAxFv09pa5RGHTBeHSG/j//XXPEa5PLZKsaEl
fQHtZ/ETGDZeaFloamotYYztbZw8qHcpSLYNrUiwlxoEvX0X34LGd6bmgLlpJ/Jjjb6ZzqK3kuYA
UXYO+tRJUsW5Cd6qUHYs/yr+dUrq0irL0Sh64vxGLG/8Tkv2samWh1d3h7XivwGOKMifGzkTUzDc
sS8Fd8uZDlIe9agZTtxtpGudNUobQpF7cLna9aBlE1drBNTYBkukTrKAuSjKakwx/uYXHJRn6ESD
GlDl09UX13bEh9466+Tv4OqSE4kBQFbltKgfJIYI0Kr+OF2/bCJWawTrzQ+OfssqWdSrxWGcw5I4
R5I9q0TUm/ervl+wAU+MoG4enWzpp+ub8dH5v6DD/gTlrgqVq3HYe73o6VBGAifaP4tysCAs1tyN
d6QuhCORpO8C9LRKyF4vcP6JhabXxG7K6jQ1JtwDhoFxdPKtlo4kyxxsr7avTMvDdOJzC3tkrLty
Xn0q9hhGjNWHZCJ4hKX+/RRrk8DdV4IWN1MSCklR4m10vbDmwWYCd51KAN7glFvlzdO4hsKATisX
3JkaLrzyLc7D3bE3ndQm0HW1unz9xfzSVcZbsunpbQmAgbP27ROX/fMtyw+Sr6F9piioJKTkUjrq
OnxGYGRH6oajy2OsXNmyXJ8BsUA0C+ATwp/ZAu9Vg+/Uc8Ocf6B+4d/K3BHj7ksUqMGTEZeioIhe
DJNC8LJW8NXWytXI9clD5SUsG71jOSbzRJHN38QX9/nWAtGp0/GfxkJwYjkCEnIlzU+kppJsde9B
m3/mqPSk3DLPyEhL2YUYOVNLV2v3+vQftNWvR2T03PY2BDjAG35SMBC/IFqbTMtMJ/4+IAT23BRx
hOBXFxTG2psejImkFNISQtVKmpYORBMTKB7XAVVHlvXJCyxiGu2kEVRwSj0/r9exo/IoJ5H+4/Fr
AheNVeSKzcaJsxmfkEMb1PFm11d53hNUBv7ss3bDSrwoAN6ESgKwtRow7+eSXzWykIwgL2bcUvO0
QL+GtuhSZag9cCzY24oE7mdZaQ/RBesP7KX0EQhYY138wZluR6He2z5/3zQfCJmYXaMCdW45qDzz
bGrqWUX3ogOEoHSWY0HCcd9YAunJn72f214NNR9Kx2WRPMoitEPiC8iFBypzDqmZkedh6BcWjveX
9isJBRUSebx4q46x8ztrLWDzRBDdEXtpybiPsq7RUzmtQ/RncwEAK3OOX2TeQbhU7C4Z4BDQEB2o
CZcfiPXekaAdWZ6Xym8lxwm8eT+auBA3Mj8uLtPhWKC1WHEabJEfjxQQR1hv8JCZhjTwQJ3AFlYI
OhpYbpFK2Jc4rPR7+B7X6AOd9ei8wwfsady8a1GLaI0Y29pVL2hVRlGKiBB5vi82tFgqdCZNzAG/
xWxQzCUkCN6E6DqM/OYFDDoaNbkwH7hdYOv2lH0uDoq7lpXKu07VV2w+tSGveQlgZEt+3FDBXV7+
//rs2SxsHEkve/RiuI5jlE847EDdda5aOWPCILkyJCY2LFz/zBZAtuKiz1S4hGZzNvEP/kiexi/s
54f08NZgMcjOt3Q/i7QUAG3P7vGAakVTHJ5owzzpxLRyapSQDjVgpPlXudJtpwXef/fU0ar/Obsf
PRxARDCc1G0RVbGUw8Vxtx/xC85YHTw61UQ0uf+zZ0eHJ8tM+fmCF/68MXalzvl+j1TIkBOfqlK3
uMAib+On9cmAUTacCWfdNKhVZUFhNM5p5gtZ+i7JJfYDHfe5a0q3nWTMtDFJZPFmnwNXgEcPMlnf
FLyjs/P2o5f0q/HluSke30EKvzswMSxCXbfUgCZTijoqMivWlT0KTPP1DaLfrkdNqGyldr37By7t
2Cp1vb0lVYjG1ObEDXV5iYd9BLCBs6kBwqGmJGQlQP50gXydU4v6ivL7yYBB9slmMMNPqf1ktd/c
tcq2k43OofnHpeWEQHGnqrqK7Tk4LBPvtA5Vcm5zLzWhr01Bi0EaMJZVoGXdFf4PoouOzFIBqo/q
X3lrrZY1JniMcLRYiitkJ8zd6fyH2XnWqs1MK6uU4TCXgB3UWf1em1courXMs5+OpS+LjlBh80pC
vIIVabcO6jJqBlSIRU221U3nCghQxFrpVwXc2sAAS0IIAtkG4xh8WE1xxU+aYunkFbVwMWpfS5q+
GYwnisnj8P+NGs3IuvPH6qJ8+YXJgFcngS9VxPKXMAOPL2s5n/DFRdNSmh4FhinFMxWfx6TnDFiK
SHJo8LmtL8Ssz5SkpEWbjczqutSbTulDd5mT9y0M3/hJRnu1qGPaJaWoKDJBQ7ButYCYg+FwixkL
iltObQ0e0+rzmKftgFDLCVrqnvxSEDx1so3zjQDzBiAXc7x2MdkZDFF4XyaRj4PhNCSV6xAE4/1m
a1iERZ8VwG240ujPZBhTjiES0T2TfnwGt5Ag8vbKFrYZfHhDvX8fLo8qi/f0nZLBr6cUWGO/p0W9
8+Zs2VPfRMnCKXN/DMyTiW26xes3SdhRoC3MFmZJC7G3dolFlZqjIq9mP8PKJMyCMIo1BdERTmrm
HdsTFYAmKbmqq5lhajaWC/4dIhhg15AqngiHTxzcwFEgw8KGS8tKbei+z9La8nYEVYVVLKdv7lZ6
ymc8ECnnablgwzi6l3lpNJYwKc0G6+2IpbKrtkyzUjNif9VcTfON85dcEOtO8HL6pMaag53SYs+3
83Wr1lr37+AM1zjq1I7mA1iGnAHg7mC5wnwL5AI0H5NXuPM5mQV4WdLLHgmEXv8QNP0XDGKYCQlQ
M/txaUhkLfoPx5OGecLGuF7biJSYw/6yMhbWSFT8agEFWfJceDyfCsYbdMBQn393+Kz6MM/LmsBr
lJhDWsTkzGCySIxS84j3PTkIy2eXEDZ5qZCOdbPsboGVdaVzXvqbj8foBCX1gAtppzANME4dUgpY
4KvRA+5560xwoo0Kv91Fqz/E+zpNFy5MhLAbJBeV7YdJ0yTc7xuxXnR/h23DbJTkz9o+QoHuc/yl
r9Kc5cUHWdmcq5qSCh3fMAnLVjk7LhHwdqglJbCXaqiwpRcEq+BiEEr2QfghicRvVoCekJzQ2HpS
OVFIhucWq+L5GtnP3I1mx5JdPAWSayY+fQokPmcMKBsyg4l7aHo7FeWD73Y8FiMOrzBKQIAbxzsv
cOPghNZHsnkCGRuEf3w8A2cOGplECQza18QNY+oWJ0PzzCnCLfDfQH7d3qMeG7cU/rlztsbFzgTV
yD57KTpkhMC7ir1J3TkhHU5NW3tx/C8hkc0NMcFSHnqPCWxdvwm7aZvDxxNEe76rRd3vItiMV4yz
Dsas3+pr8xovZA4ScbMR0vFBIk2CfHYLztahctTvYld6APuBZbxPDrNL2f71fbeNTZTSuBq5VWpE
QC9gzIKWo27fMF7TJr+M7JYT1a/5WQeulktwlykkKuc9c8Q8MCUQlGg8Jabun6/2mIsK9GuJBhQP
uwYDM7kScIP3BVPg6Zz+mu0u8AnetqvCNbPK+ox7NRzxZMXr59Nn07S9WfyUiYl8rM4QBt7bX2a6
9Y/Zr79NPyOrGfm9Mi6XluEZFDLdM9UXiAh54r9glduHn15Tig4ZeWg+BOBghpabh97Agr1FIwZe
41D+Oeg4K0k0XsNDZHJWeKGRY3TsFiWZEYohRZT3JUa+QhFQ7Z/4k+8frI+2O6nCrSudjYaxaRfn
qXrrV6RpeNmAEcDsFZXTKrcrViEvjU0KUe3iAjm+ccPfJNRExJmwmUfnEdpBm5rPobslFf/DAoxr
vv2ItWWdY/XRn9SX65GTbyS+Y7Gw0SSrqAM9LyzDFMmAuoZ10GKsTOxJAJ/KFZpOFZ8DB80OlPly
VMhPUy9WQHWwmrFKg7ddS5FfgB0+85PFYB78sACUExEt5qVqv09PtCcDB+TkgrPvrpSx6/0cSEec
RR5XAh4KJzZGCvaYa7pJs+zv64dm9wZ21dHGX1RxknoXgyKMBs0b/Y+NbqkVV4ffiFatlsHs0wjn
MmHbz01RAefwDyEREqXz98Ug1mUlFLRbN+0gKppLOr1Cd3Os5+kDOf8yy9IH4oa66acThBIcgja1
Ckv9iVow0LZ3NMySL0DyWt3XjaeshbTWtHH5BIBb2ktrCzK/u25ay1RFEMpQ2SQNH7lkJPIWzwCL
yfUGqf9pQ81cZl/we7d/Fs90qdUXwinl3r5kAlihedi6opkMeABaWiqZIjHO39vzlHdQajFB5uIZ
bqbxaJr2zIA65U4FPc9rQ2kbuX6ukZ1VVKRCFajyJQIBWUFJsO6wGRBsDsLqX86+vy2BvVVLHAWN
mzWl7V52R+hGug/30lwPbOSTmt0K2a+yr3BS4XbhdhmJcaoZzhmJzE0CD25agk7SRey/TdMzl4be
iKrb99wg8G7YXRll9UqHVkHAUBLP4lDlqOjqom9gEBdf497IiKqEaacZQ4dloDwWdtVDZKp9bOmQ
+qq0lMMWMv1mElLsfH5WNOZbbETP6umCIur0FUBZkFvGkTUZ6kwY087LWviYglMKuSEuZuIsQcaT
R/OGZksadGtbl17+uBEtk8/NpiRYTZ8yqfj+PJ55/FelMgABp0PMmTk7ppw1NAtk/4G4P5Oqul08
c5H3xFDRQe4LpMU4kgTXNBUSVwB82HsjSQ0tzta/zzN345qG8L7OpIK0xAs4E6Lm4fINPsBC7Lz9
k3hn8vKPJYxhfYPEvht6ewE+0RI7wnEWyDadVryb4erezK3nQuGIIym7Gf7HagFyx9RdS0aycDPf
v7FvX4JsfZUsegOU6aeywPbf11B05bNABrmUdPylS8WcT8muSsLbhLQzj+ukaVCVTDyAfLaYaRms
RDzxCCy2+Kr+kELRPjHCydgjRlShuy/cZY1WvjKqz1+PVrdvkx4i8Qm8vTXs1zK4+yqX84CbVoU1
/2Uk++R7+F1mx5lFlMkroQXp8FcNwnx7+2hjyNfhPsXyQ324Q3/P9b2ZorM2jafUFKxXPgL4IesV
lp0+7u7B9b+laFu4wyo5JJJrVn+LLdC6YaERMvtCqcggrShfgbOy9kMP7w7HWOPVP4kXRJ2QOiw6
9X2y4/oiEqWwBYPpDaSImCcXvDUKugvm40Oyt87TFOHjV/GZHd42aL22PoIjziJugozDW3MfyH22
rYIg+2iWRVmEq7pEMJ6DXYDEP4lJShRjiK5wWzgw8+USqkFgC+O7liE8K/Wym54ssrwDFsdeLeAD
ZoVy5FJOgUuKeuEI5qFoxHLYXbqQ21QHQcJV7vX+8xUyi52SALx6BbaQB1jyrYuplwIwNVAT6c+/
VFVr56y7AkRYK/vBB+upZKFXWsAxCE5RRiLWq1shigPrNFPeL8xf2JvySLOxv/chhndGbilR8AP/
JDKlTlK2ZTWPH9ldQRgkDHj7Ee89HdEet7tMkj+q8iRGDIoi/ZLgYrcKwadjebjcn39gjycivGSo
DF1RnKJPLtXl+fS0bvRtcve2UZ36xtXh/Lmcj1TNL3yVhVxHbS+z3CeoRwhwzkfE5IC5c8NezmfW
D3JP8iWSsT0HUN7OH7krnH/m8Jo7r/qJ2NZEtwGmhJHbT4RjMh26s4UKF3tymcSncWRwTLXhy2g2
I1MUZt7GaU7Om4xevt0KQnv0JCx/6eLVbPUkwPRaP+awO4e1OZfsx9zrz+3O3iqrkEKP3rxN8/dP
OXCr7USgSs/K/rG0czYGIGX8FS/QTCpTx1Lj7/OLognBx1xzKxUcQaKg0jeSOBk8IwQejWYdoLEQ
QCG9SLPdQVwamZQinaNf47zt2cLGFXFr7fAYA2d4kee2Nv5+7239uuBh6LT6f1eD2FEK/lNGPeZp
7odyMcwfILnfoXUEHRT0thKVrZK4LzVm1ziH+4wvCMRwyqPxjuPD2KGt6DPib9hwEUsJdLyCXm8/
4ysD79t9VsaohsRczp7keF44lyeZZhYZJI/FeT+5oKHZ2IcGnZyUU/mGXi3dBDMLEjLvhcpmG9Qc
/NhcasSIVWv/A6QFh6t3TsWr1dSZpKU2elZ9uzbjPCEFkcaGSjWjV1FFcQQFSf5MjjjBzknvsH0c
emAi5SqW5K55ie4S5rTIpWwdH/7XAu8uQI7sOXpAWqOMxUJ7ogR6plTU1BXeHDpVt7+8/D2Hx7ER
UoJrbPk5xZBRgAH3fDl1HodTujJdS0S7nNUU3WGRCSUGXGeF7ehxzifXp76wgwx6Lc+WLUX6ja+J
xy+LtV3IPoyedCuURwL1MHNZI0qj/LpOLvDgYL3SGlDzUiePSFEVKw9M9YuAkl1tOra8zausVLMH
TdwnYxjWfdKoj3HswNMW+YvkBr8cEU+orvnnXptt5hNaSzxn3ro4sOSPmcs/JOCsd7hHgJD6I5tX
/EBi7uKwAcEhmJQmVKpYoAOGOkaO0F/0Cx6RiO7K7N4pC/DoiV0NrQu0kytvxqDfr/fDKL9Jw+kh
/t3M9sWvhDkK0Tzleuoc4Mj0TtGieIF1KXFx9RuetxwjL1vbqHeRU/KAocmdSmOsWp3HAc3js90G
DRaboiOjaIA1CoQI4OLNViVdbHD4kzre680CgHTL4GbD2DjCEDcwoFpHPp6TPejG/nneoMh3fCY+
wWWEvdwWaMzsYUXJ5qnE2ZovmbMyjTexuTQWJIpXxftBWBGjR2JTdBj2OtHO8tCR/iR2AdCZXtA5
VlrMBrC++gtG0+NGtnXFR1LuEuk96y88ZLuzGfd1W37YXZS4XlL6Mo4il4U9WV0bJ3Se5q4cS2Tj
nvnXcfdaIzfF2fGKdU4e6M+6i9iTg2A7OKwOqPw7BW9umhbFH6uJwvC5CLpkEodD1LDKZ1iyT3qo
KzM7wwL/9taQjldE53tskC7TT+5BXCkmT2VP6uryEWX76P/rlLPZOiimAtQy7WeGPS1dArFCuWKw
/Tz1aaZSOL8J/DUkDOkoVXBiY8Og8utirKrmIx2x014NCIYJA/lSyVY6pEEJjpJu7K2jbHVs1Crf
shq6IA3QJT7QxTFTAV2uFew1ziIPcHjPH5eUZeq7RhQVJPQa7sex7JFBcbV4HpD1dGGIV7yjxZtC
FVUxf/UE1js0irQ6fMhuq5eN6vSEKwYe1cpbXQ/UuuAO9TG0/k6so0OcT1IY2pQPYPX0IXTIDTU6
yNe3yw59SA0KCtmH+T8ZzwpPbBaQKZYpgPYswJnTrQPXUbnnQ/3Ax+X+dzdNvaJbl7KezLa9583L
QdtgHQ3lc8p/fB+E6bkAWm2+yAwDkuUVz54HEZ6Md8rV6Y7k4T+twgnOaIL5tgti+kxhISYfBKfC
w0vLaMA0jriEkPBWD2I95RMPT7FcAXEzts8FIBaMDhJas4hcfSsrCHliwuuT0J+YHdEqUhNCQdAG
tSb121SQsIFrBJds4Rigpt8N94dfysBLGFHSFbU+pvdm5/GsBz84CtsCXjqaQCQvgdGs7a2g+/d2
+/qACrQaNAXpwFCPs0O3nYb114KrbN49LWgZyoUKktEiveTDBRdYC04c4lY/dm2aAoc/zD6wZIqv
IpNq9NT5u2YBunFfdIHj0o2pOipMtcWx82mITmqefKcUT/ct89GAkYucyrL35w0RqEbzJ3uqb9My
/YAIwzwYXN/67xVsQFPlVXilNEQJdysyCOOz6I2OBFzRN06KRA8UcR/wg1xEcQ+4FGctI7eGyLS5
fj9MloLVNAFo2nTFqCqhwjazj2fhwxwXokeKzSEd5xdyB2mMeantUL4sauEB0f/jfBixF8v+i5i5
uY2rEh3dGjmPTjucbQUyW+gE4sFuxYW+PU3ywlvJ126+QA2C+cp8Vu4Ylqj4/uIpfsVis1mzTP44
cz2gmJqzcazhjaU0wc9jeq8uTfQpZU5CrbHzi4kxzOuVLZvupq2yZM3afCrMbY2pGEheh1VdvvMC
iXFNt/fERT9L5BglsQcjdiRsbiq4+InFcjnmqWn4/VBXew1pNLXh2sKPmJsGkJ83+T9ITtflDb3o
hHoQoPScbH5+9HBgLQ507j77fPrqQ9XsimXcRnv+UE1ScJpqOdapxqplT/k+pYd3bmYspZMshpCV
zV8Qi1Ze8i0h890f8dape4QddjfNR4bxM20mGk9gbEl3GDkua0nrzyxzLVkN5UFxqmM6WL8HeX49
3Kg25/4JoH2nc31hfMd4c9nNAr7ZD9AXlHHKGxrcSvWf52Z0H1HU8OpTcxgOJViiHbAR6DTl26dD
YIELQj9HSEPU2W2S4vCASm4V8tS0bbE2b/BuUjA8PBYe3+YCg2bNAeVVk0ZnqX0YskrQrlIJQrki
xgyhxaCsSD9tYi87gp76/+UnY/TQKo+YEoD8VKedgx4FiqF2h5MJp09K2eB/zCrtQIRduyVG3a2t
YFsfKgUdYK57xsVtBnOJmrAsrnXlbBR/jCbyatxYcIpdA8qLQA7BoB3KSUNTU9lo+uDICuKuJLjV
kETNoc21tFIlJuH8Ltav8+HGvmw4T/6ctWupDio/xxowzbQK5D44OhWV3jn8k/A0osOZcFO1cxJg
AsMB/5lhyFHtBIiLrLc1NKxu+YZhVhQ010M2N2ZPm5SFt3ugy2gbbuH5p0UkCy3uR9sOD4XiIyga
C6ztHOG7071DeqC59RdujE4RRZp3KPHCnEUlkfAIhwrKGna3Eg9MOj762FjqHb5Q9N1aViTrTRGg
wa/Sv3dy0RRjgCUfXXiz9CCwU1JpG0vSTsuSZFyVN5Z5ffxgIjxR9kI9laANaWXQX7KrU1slE4j2
EkpZprGWryap4FH/PC8FITVMOkZH4WFb5cAvBTbnGhvexsVU+ID1hcuXMkgJCiuE823OxloCLJJe
IZyJfW2RRuVyjsPP6NU+MRRRaESGhcwEdUh+hwoxyO3S97tKeXJmIwXfmcehSyh8Pxy97lRBNc5s
XICkdlFGM+DXoF/684qO9atrgDD9zp9d0i+pulKsSMsac9TShMIjD1cDht0IHw3dgdh4Myvt2nIE
LeyehFhEIVRT3YjMi3lnE9CPbmMn3iq5H4343ppaKZDHtN2va7xDRTh/zQJfYBcYtlUM/HXCeJhB
RmfDo4DwbjU7pA6eGqGqCCVJVi41y4IPNspPN8ItQAAuQVNwgj0W9D8yanZbfhOHGzWFdgz07o4+
ASBSOGf+EkVU9kcuubZ/7iShgN9ep9C1M0m87nCr9LWcSIrCAFCjlX5BvkgKNV+jSCsi5PBvq1Em
zaXB9O2iVvCM2tdZcTe2mUuIFBGSP7M+DDRAWk/Uk+nKPF/A7pnNn/7gAhCz4jSsjbeybL7kAAso
Rjkd4k+u4d47BJqFUK+/XdUWZFhMcu/OaLVmcvxjTug7AiUyR1qT38wxlsc09lISWYCt/IElAhdV
UZHKgSa0ULy7wZ1Kx5HvrTeMrpR8xEORTDEaDVCN+tSQ++ZnPLp60tw4zue9iQe/NB0YT/CeZWDK
CAFhWyr/ikINOaSG3/PODb8ZcLsZW+LRzLAIRaR8jQADxxQJRH57gaPoO/u95D2+oK9KU/byyjoQ
o7/dSN+mSgQyWce8dmsYvjMlccyOvUPpKpQgHajxwBMlH3hEL2f2mzauqrd7IgmdyiSTkda8jvFb
/+v22gLisl6d8c99qTcBMw4wQIEsUnfv6PsM9JwfgCHugLGL4E7T7x+HIRFf9RpEMP+vRMBCJOsw
3GNvNppxo6f9/3KeH6xAJBauC+5taI2GbRpfN827HRclGX12px+lnmp7ZgCbVz8SXbSYPXT29CEu
4eW70nKBoHBIOVqLyAoUFX7lv1FgzWkJKqnilbn9wRmmeLO4vSGS0/lKAYvW3eo0FVzCqFBJA3CC
e1wZOnmWH858EMbtsk2LiGgTiMsFcCW6SbfeI5ZxpHsGgQZ0dW2qgeV5jqt2WdkKNwhTCYfS1CJA
tA8Yon7TGS60X2hrt60vOIiiN6YlFkhG08AcerrytMfKKygVdS7Js1Z7GqKCky0y0I6T6TOzWIG+
y/L198IimEPthM9SQIbYk1/yiJokZVjS6NwGmRNMniIQQcSD8jV7owSEfvwevyi6jdCae6wBDtIV
ZOR/owUMnvjvOR2yVJOtcvnZbxZqPiqjHvLPnK2xa9WIsnWAEGYAdbhm82CWixQveFu07r3FM0/c
Hovzp5pwC1dQXRZHEKiZVDy3WtfFixu0hSzsY1YdRNYIJIUCXWvTUCRMbhDFfC6DVc3vQP09s88j
tMm+K891SoqVyVmXeHWVRybqBAfTmoI07Gnix9LYxUnZEgVTX+IGtDhn2TUQRCOkpxzxAnvJds56
Ba8sLH0s5oHsGmNRducYi6FM/8E8/KUrJSpT4kHnntyW1kx1Hu3Zn5AqPx28m7m0b3eDP8/Ps+7O
vDLTWxYEKxuz9Knc1m5TOigjJZsprt7RR/a1/cxJIm0ujqOFwzmfWRNfXA/In4y3ofVlHWOaU5SI
jDBR1ldwLHewPEBeaZswCiWTNz0nYk1tOuvabQlW9oxpmfJ4xBxaMqoIBnbg3+GuAsITiZpp/0jh
dGBqksXdxOvPgg7XFWoMMU/jSHY04dAFWkyDmYBvbeGDKmvWdggC5hl0IjsyBic/95KDZ5VeEeby
GulpRbUgz/803PFVXperkRPKkll0SkcPK0RrfGe4/qaLK5XYO9+jG8bQUiLfbPEqlARJQNX31Wco
73unXtJnuSrJcXi2bjSOiAVMIbL5vEuTC/ZUaePtL6asZdgNsYL7NxWVJ9hInQs9T7d4zEYrqUGW
uWUrIQ6t7FfWQSyULzkF8I5mcxvuuT42weG6sGMU7HsvOtOBS/ovYvVDWbWwz+ePNn3kTqD++/pC
/apDsFKiqzRspQyjAQEkEHEixc4IvuTmy3vnmiRgnJWR7Gy/Guy0IyTehz4VT3T/1OdhfR+TEeiN
ShiIwzMGkYFoj0gRLppw4N6Ug9q8NcT0QASk1RiiH6ySyLGq5JIdiqWUhQ2+g8DaejrVKAMBoRBl
tfTt6quADW6gG1jBB8wDG1bdDf5uDJCz8RWHc+mud0z9dc609XYSGX3If4ZGs3dRlWX+XkeSeRdk
DuBleFoc6QOyCo6nwaH9HHHvjJ2uEgZLG05FZNRE1g/n1XUYABVMjJex58P0xFgMzJocpqLLg2hb
s9VNy5+NvtkYZGavIYswiAAGsIls2SBXrDOvnpFIK1gTVTWzE0HrmymrJuFGAxFAhFSBWsb0GEZg
Tik5yTxam462LtZo4rAafr0XP1XGMiU2ZNqFp+qJzxC0JTer4QgCh1ZhSfVrzv9sj6h50i5I4Bkx
Jzzu2ha5o5B17YlNQ7mdmjRTRvUA/dKpIr1z13E8+GMhDOPv4XvWLG64qILalgiNGpYoIuYjkr5W
L+lVuug7N3BGBes+01dwfa6ZsBcONpY/GiC/+eQ/3/NeGScDhHkr0ASnjlNXqHdnEWEYmZJHNLTq
TjednTcTobJPbTIYpk9NnHaSRjCogWBAVAkpQuDYWC/PrRCkf8+Qmr87k6lAwcrCGAbest00h4RF
BnKXRBg1l7zJN7NwQeuMlHKDfA8eqaG4YcZegE8dAaemLMjhe3i0ypfmtwXcBb8OMH0VoAD5HX5k
U/tEv86BQkB0YD0inwcsFMFut+hC3edWDxCK/xxf4foQrij6xTr+rX+haY1A9wbEegV5alJsaaME
zBPfq5hQA2juF610sU6cvC0E7SX+DkWQGb4MyobaWQVBcFlbe3gZND6nCJ+/aSx6kFRg1PUjDrzA
NoQRWlDeevubWQQKKiI5wEPmJffqX5sDMC8kViLoYRQCWvWHxUIcsXS5Ou8ttrPaFzeLjpp2W65W
g+wTngBloWHv6M41tRSt1Zci3Q6W6coHR6Q7Wb+TQ+JX6mqd1opEIMH8I4qlGiqEzBNvwgi9Q6Uk
lB5U+14f9PMUAKLBQOCBX38vzgZORvD35ftmNvlTwuWRj8+B5d+uEZdcMnMC/vaMzg5V7z1zYbkp
nueC6pn3YNPnSi0P/mhsZeqMyHzXU5mlxGZGAINpOx/68t7oUHuX7+cQ5VUAZpIuObGel7b3mtRk
L4uywYGLc7gQ3iHihPqlGUgLELda9NI2L3VlMkX7LrY6FxjD1y2HxDA2siZhTshSjlzSWlzWmr1L
H/8/NAFgWdw4kBIxMC4Em9zwvVroewvMvW0GZ75NeZnSFeEvZcVqbQrD7B6Be6cbS3WpfvS+qsPC
P3RGNJWcWtWVrQzpsKcdYB2ni4754yepBAn/PSGrT8ANtnGsZ83hy7pmdCccH3yQlnvCH61W9uDn
sqelYy21yssjm874Ry/Rh/VfPFpjMurL9fHbAI4pa1e3hs/kihZJgGlNny/xPy+Kl6xXzgMeJqVq
TLWaCb0Clj2eDHYOasiVWzX1nQBTbDQg8zKdbQK5vUXXZF4b7vEh26nCfCAXNah80qpzu+rGES2T
daAVErSqzyTYqdpno8qJB+Mrn2TO8oRDPaMuLob2il1Ix08YzAABEYKIo8hFIgwtE0gN8o479N2i
Ft1t4cHHWtt+I1Olf69KfjUtX55+CAgrtRtP3ScjBM/l1o7ZNW0r3Ww4VSOFaCaCPog7tBUSvMhK
2dhM00Kl6/T8Waz3PL04us2rlxGbo54mBkpFMZFKDEbA1MbeM2pmKi71C/ZZqZI3jEK6d9uUf/Ve
RqDzXyenS4OfUc+/S7Y7PE8NI56afgpHktKs5j43GX/yvxJECPAHUNTTK7nh+e8Pefd3vMbMSQds
77wlxiXtePf+JUfu39lXr/aSmQSD6f1LR4fzYVB1i8DR8n9lrqqsDaqCg96b2EHQKDe6NiRarPON
HyDF6FmOQpY+iUDX+sC29d6w/jR/UVlLtGxpu2to9+rSAZS3ylWaQ9uIEJZchykVnh5g/nU8T2QV
e9rhTPw8j5fxwOpOtx1qCJpmJc9Dpy2iZyN0du3u+/kIqmoh+VkQ9MfXKIWrkq0ATgYeqYCRRCqM
ZCmk7uDRKxrlCdblm5Eb5ftrfonm07YjtNQsXYnHPa9JwM2dz2yZF8MCzPytKPSF4NZ0nlvHmdlY
5fI58tsBBFt+K8WHYhRHZ4yAz4a9DQxAAo5jZJHfZeHtPkZ3QSfNWoeOZE9j4U5uAx//zSt5IpKD
+QIWMtzLPqzkRn5Z9RSjVtJEE+F5/rHeXdFlRvcejitGT5VzcORA4L7NJDj9ThxnnBwAGBD024EV
mbqN749XHC4a3Jqi0G/bzVFU794XwE/3FcjaK/ZEPK5TLPZyz5fGU5pHgN2zRtwES7PsFwHTH6mw
DsybBn5Ma5sW9UZ8bOUOK284x88RrX+ZYXwaCkR7Rqiv8PjNwXmxKL8JyUQnjR9KYAKILFTRCMmq
QvVZj1AB5bDBT0a+KQ2jRYo2NycWylXNXR3oe75rJYp7L9IZvWTfAatvOdxbvjaP5Quvm9Jnyhak
EeYfK4jHYbev3+35pTB6L0ztQ4NiroF8iN11PCUwNR04/9APJjKZubfPH38W7cNNfW/Eu42zc+7u
PZ0mBvD1ag5wL5IKF5pCsKEzKFsQU0r+AeQXXBXLjD/hvstZ4U/wo9mlzHLk9w+yLO8IY/ZPlyLe
G4a6fVR6bxJL9I0JY96FC2Cd/OXN3E1JBtrawokPzsCIKMTchw9ZgZtem7CvqeHTAhq+SfbJuTJ+
sKmDMnBEpHaCgnBIKOQ8tmRaUEqsBpr62VTd5YIiwHWNfB7Tkd0yNMkKP+V+gM9MlIZMCiN2R5Bq
ZOauOkDiWkXwks5jLbgEE6p1saEL3Q8IYIE0mzdOf5ZXrtIxcReaLKczSymsR4w9IEimMUQC8mtQ
FhXu3FZqIL2skS1URpqJ7/KiFxHXIxzSYR6Dj5TizHNLQmYRuJCdcNannXMZ2f9N7yh4mq3cb3wr
JrhKBIkzLmKKXTif5HLRJbTzBjlieowGxH7fK5DPPAnGi6iH3GomLI6ZCQfJP6Ml1uXtCRe9ch4e
6reSpwN3j5P6Kh+VRC4LkgIeGji2hOp1KLz/XqkClxbege0saOuYiHqzUAlaBV2lwUMpdos3vdSN
fYuK3bVRCClsnjraUFhPasz2+3Gmg5c0661DqCZRYe5GKFddQv9s3ED9FQ6YGA3XnhCDg/Qen7Wz
7PsnkAz5ptVnL1wrzvY8W9+9qgdvGnPxCq8zM17ZtwfXOKwEvHdqI3flm0uJ0IQ0BFg2jV15x1NE
mTCRmPBWH7Gn6xJvYHaXACYYlDWtgP72FAs51C6ABzNvejEIbiBk4nTG4WF5FGdCA9H7V90rCQWC
bALOiVGvDPVXD7jZmYSTMUi0GKbsO5SYYSa+LGiF1kIXE1sVejHq+aU/x+C9cUxLlcT0G4ahLVxQ
MIIY9wI4FU4Ngk02mI6f6k8SlQRn0HNBa+1Hb0VAjOrKGr+RbSTlNVCZUHvSPxJ48O+Sq8DML3tG
F3V5f/nKZuHMSVObPMsUsMLX9dNKeQcmZddyHenryVmXrW8g5VBClVqEW9lKE+jtUbc/n7C40nCe
GbYylRqZxPkGtuYLCqUJqoOR1coyQ8gHHzXe4wTy3N+SO/eWQ+nFgMmMRyG+TB8hF8Y5QM4BfD5Z
YCdAfRNNMbCiF8rCECm5vGkPBPwGt5LWp4OW2rN/0wCeMo+2T9ksfHswev89UHZb+o2diNF7ZGcU
OM0QaOYI3eJewjUdnNb8u+BknhUDv3dcETQy1D8fX2xmUkoFFbb4+gROH+/Hd2U9HxW9qmVHfNwR
2j2XFDeTdJh7MQli4Fq/LY5HEblbm30D+fCAifeHbBEeX+NnAZqeQIKJbnHsr9Bb1GTCTMYaC30a
7kqwHOf159fKrqDWuq8AzYkWL4QBBSp8YM3XSuttZF6MdN60ThfinJ9e8fD3me1W3mKbc71FZfLT
lY47+W49Ij49SL0yqe8Nq5UIgE7vH5x/jUsw3AyzanNsrBM3lGZ1eG1uWIU6IH4AIxsfk0aPNJK8
xPyCYGHFh9CdyEy1d97H75lbvZyyYCOenl98kIYKC1m0QLSiBVctqZI/hte+gkq8CUqCC8v4AlNU
iJKIlIBlBNHThDEEd3gDTq2Ufg89vhLDRRXVVRgG2mqrYhT9HJMhl3L2kZ0xjgmZj87qJvn14G5W
nypmMukc9yrokkeSb2UAT8fWzazX4q/XENwCsfXueeA9taI1XqeSNn1DuDzwPqKEsqUMyGdmXUB/
xNWdLr9TDvKasbYY73/rcnWOkeiDR9oEwXldkvMpl70a71odkAwY2sDZufWfnsrL6UC3kUCvOS9y
l60MjTv/JlOF5VNAhdknokKc6msQx2f8kTwO0T+Y44gqDC02lQQE4H5iajlcRoDcoMASthVwezYL
+SqEQfeL6mm7K13H4u7w1Csu5abe0nJUS4p7tV1ldJn8Gt5ZRBbWpOWXpg0l27ZYRXRNKWfCRm0/
FNzx+0gd6aoxTq4rlcPo4kEdSJZ1jtC5IvfS3XXAL0c4FvH/im4pGrXUx06la0LMxOwMOs2fvpAU
+GJKTWykw5siRtZclsvFCQTwiT91+izCkGFmchJWcRVMG7e9LzM67WMvJfdEgwj3xZAZju4tk+gj
niywbWzWM6SQHFlIwQjpuKjJe+6K6Y9eMBQR6mtAaOUs/S1m2RSuS4zg6TKyEsL/pYRoAB6h0Tp5
mte+YfZvaBwKzYhE7rXhTFlK5iCSC90HF0Z2+Hn+cp+dUx9k9gRwK7Bo/xXfVq7CdS0UlJ2PGX2F
uv2lrN6QcmVYBbbhCx+4jnuWC5Rgk+ezeONxAWWI7+GmB2x67opFMGFhVeeOxSPcrx/Ubq5jPU9A
9P1xqir8WtrrPEGo4drp+n+ImmaNISG3TXIzYBeisffT7hBfQGZO94Vha3AbCBObBJLuATVLsTiE
kka2NDhm+9uLqpEBeip07ZXyZmpqkZyu5iOSxacgalwXPpcaf8qZ/iXKXIny0tjp07TEJedH1rnV
T99Opo2TUfnl2j3+Zie4DqRuEs9dXHyS16kA5Vd4xbsoHFRa56SYb8nPOYACe+misTkQsnnVFa0M
0IKyiB0gRuedfxynoQ5jndD5fwk3fikPNf/g078Ub1f0945dZEfBWIrNFq0FXKIImkv813YXx8FW
Y648qoe7NwTt9DwwD0bHTTpfgF0KqGT++PtCWUrSI6+azVVKVe2O2MQPLOszKE/1dhk5FqjYOimX
PVmqR7MMJyz+pRRV8Ll1oi282eU3ZpN6gcB5I5eKygYUugJHxOlANcCmodHvz6NtLQy5ZukCF0ii
t7tK7jJwdOZQoHn3C1rmAPK3f8T5OHHs0fB5XVpa6ZLwnAe6E1R9psSZRWNz/PYwCPQcdxayLB9j
QJqkz8qI3sII+CRjFIse23ttZi2XKW8d3lqnnMej7x2OKug1HBJA6hwP+mqEjO1zOQ5vKQKzoh1U
Y6vE2wn8TTVwi6xGNDfKvS8KAHShqh9LNdt9C5eBgr/A95noM77F06MT1GodHUwYjPTghvZpmsGw
+fJT4SkuhBSr2qFdpx38599VwYnKFx/H7ZzK9qkQ2UdoDEuM13fVqorFxis21MRqbmDHy1U3W/Mn
23qTZrOOhRAwae0pf2bAjF8uqa0VuK75vVGEGE+Hy895rKWavPUbstyIzoxzigbbnFfzSEJlF71t
lEPZl2xBmBZ1amYI8nb3KPGc/i4XZXq/x8BpkO//fvgHKevmdS1+wOR1ZxjCOarBMOTdVeJyMpi2
u5DxlRFIdDjFZGWflYpltdrFr+ofcc2wjltjBgn7acOk0p3N8dv6HIVqa+nAFeGvRoRZhiGgXTB1
29VjY6BgIvhqTlnDornkvU5g2dcrj/ZUPGry+ovtp9zERGQK/2Aa3GpBZI9MXuElkcInycwLco6i
5tG2DlhiPGEtxgD4/Pr79GU6PjdGM8w3LdgzaUxG0Bm3anF5Q74puvVoG9zSzqPfj5Mj2stMS5dt
4tfVg64v5anFYZXGdFid0e2nFzxNNKrY7NnoWFhcaES2jIl6yyaTQ0KrYAsUZCg5IObLkXlCSpau
1hZVODcw5w6gjk7L7durmYVk0yFTo4GdvME4fOtecZjQ6iAgrhIIC78PKqwVLB7t4oCho7JvMGUz
BO1HhqK3MYY6Hi3cpYO7wdrvqCriN3WAZqbiA/gXQdkoxSvqRPl0Ha1r0kTFVVXhT/7rt5EIe9MB
7vnXS8pjZITHjb0UNK7SRijVlc6ymrebw9gmy6/1YunRznyMu1t8kCIjVvH2ykPC8+fasDU2mCWv
RovRgIKkkr+320sfAW6i7y37G0l0jcYMWYBTQ/VeeqQteVJSX8jTa+HA2VhABT0c18fhFpO0Q0Lg
t7wwyKFm+O4iDnRoVR1IKMfsNy4BpYPQRKRvVhaBLahhr4uU2yan+XiqzbzKIHU0bjczRDe3XIxg
5S/CmIWhq1T98sd2PjEvV74U/2qfURYFkXWsf3LqswmbUh0mN3ggNHVfSG6lRxETKlJULJ6/JZ72
ko0tq3CabR0p9DxRWrCvuVW6mryTrsdTcGLO1IH2ZPrdMn9T3DWe0APkKj3mwuLLYykcO46Coa7h
FVfi+YyN+BYM1Yxld3YdOFR9FyTHIMxkxG/BEQIN0VY6/xBqQB3vOJnJdDJJHT4SruIjaUY5ejUa
2TMAAx2izLgu+yKmfoWNGPUKRcByQYtIJIPWSV6tS3WKCjnThgvXKx2vzOO2PGnu4LbSgpZrNxwT
dErAExrBxJrTKlV00peHT48AVGcMVXSaYMX8fDfj+JEAOttiwTwD4wQvxLufSI6Kzwjm5A8OW7vP
7DSAoZ2CeEgNzJjO3fTmyBOe//MR1YRphNykyE8PFRLw4MVkwJuW8z/3dIqeH0pKJtAn4k+shtp3
4vU/pD71Qie4hNqS+hDarcp6Mf7leJD3/r+RFvw1m19peRSRAiuEqj3YIIBs9p3nbj0wfhJ65JgT
vkdzfavgfAho8e84puzY3JsjafHmXhRsIu5KcjTBoaa7x6SgnQbNNZZGiRGAtjKE7Q3w2WNIOaDU
KHe40lZYsQx52KNO7aAkDDZEq5V/KWzVR23FydV5SLBGyi2dG7/ZcLY6sRCqTcYSg3+l9bLLJ9wV
JpoV4wKs1gGl0qdRPf9y+TPfQ7YAPk17JtYGTCRFVmU0eqpO5kLWPRsM88UxtQQCUM32CwMbaZDE
HJ20n2d+DZ8/dqn6do5dhjQstWjvqcRNy8zSJZ9CW5fX9mywyc7/nKlOohCB9qdg3OMQzmHidxlc
jtmkVHivZ+1XfnFnnH1uiCdnqbg3wH0/PrTDmJmxSwM73ZOWrvMCakteu5zz+yl1dnKTILB+2YCZ
0xBU1RS8vFBSGRUlaDt61r5lESSgKs5RAlPSHp9E642T5RzX7jaPV2/yeHdXOIBGeMqGWfz4IFLa
gBPF7CZj4MKyCq+fE53XfiigzhJWQweuIIxsUxUvAT3ExzfkSOttuJuEjVyqABIEhChKCh0L+GNU
LvUbSSucIOLCHtKp+seGwnh/dB8SW/qyLG8vuI/WT89JK3MF/nQjR3Tr5ZhVMOms3Y8UMcQcXQs7
T/qEX4JrRrVTzxaegAJ7b42SFe3fRxHkABa2MwrIpxzTBJ9xRhgrXkiiKeRG0imXnd92TG0MvG+A
a2hJ3mYKAZTP/bN0/OJv/BaKwGRA7IZlfriuIhfYLN1xTpjmrRxcNPKg91vxcsjdH6BVsrtqS/ES
yzZhsC5JPhUhqBieMbJFXNJ7SqYRBRQmWSLADQvwRdFIUvuB9lgrlwS6mhJeMwBSQluvrw1GPgad
Ne6A6h9GdryTDG00ZZaNsLt2uMsiOeKCR627952hLuANiWHT+1wPhkXdWGfLmP0s+dyZH2bQEW8l
xrLt7qKqiO+IDbunubrXfgFQVQjazLH3kSe6MvukrT7/27S6635tEjwk6JzLQHRHZ/g2RfVBPgNb
1FCRVusnwF0wzWvZSqLtNpVcdtWoKYfjaeikxithV8wMohBuTOibrhe1/4/5miafIho3EPZ7rAuY
sU0V6pxjspnwMcTIvL+HNlp/H9OgqF83UKX6cYqAndQbzEoUZmJwAxxqoL7+/yj7kHLLBPgBdZ4A
C+xf5vmmCfxTMDKe24Q/yWT2czcuXt/nxSmpsN/LbpDo7ZEmu/dzqyjfLODhvsU/s/pJ4jkMZ8Gq
x4oqsAEwgP9lpTySZpqPg89XAk5no9Ow2RzbhFQPruVz2Ek+Q8phRG/TTdPEq7Om7HQwqRV5BIpc
2EJPvoXmhbblOP/xx8vrgKzbYDIwqGwxn5cRhC1E7iB2zZ9xxc3wvkB/8eHEgZRH8IN4gTZMkRi6
BJsV8XhrEgXEznkCcdDm4KyYZNzWN1pY/S+zzd3S4TnnNHRUDottCYu7Ayr2mXUncdcnBRVK0Zr+
bLUrv9gARDfh+Vgz5Ceob9GJJkFuQLGhXJIabau5BdY5md3/krB4XgSeOyCT9hQ4OnkBtLx8ONvd
/1cQyfnCqAJT/wuiJ38qv3UsMVYmAkV1pWgUYc8pe2p+l2n2SBJ8inVx0TVBCaE+Th1t48460Q5m
ql7K14k88vqFVfq1Q6ZVJc9Y3zhu6OHsSCkgydV7gswW6dSDPTQRad6A3Gt1CecY7iTAqWLX2gqE
DiXcNqWmsj0qGKvbf4MoHoruZI+gWYVUlE+dGbIjoxsj11Quw/UCKka/Tr82vp93To3JTsjz8iwE
ahfa59IgSpAZg48wXDSLT9wFuxP2+1QiQFp9WWorzjAOmyYXGus/K36YZjoSkEvzAfWyX621NFcy
6cN34ENSQ9P1VPTuIkiCbsyOfMZy2Xxl9rmgwwRdfo4rDp/hLMG9MfXIVJ0yUJeODKJSnbPZUDoD
RjLrMkmw/pyny8uuOI5EJtT9A7NVsxztUNO+fWwLea9wD6PCEjksGrLLvfTiLDx1tlya3z+iBins
rihaGI/5KQ/d+LPfs0m74KdrYBXN9Hcux4bLBj22QlwVTMayzT/Tt4fgEDip+E3ph+tsTIF8sQV0
lAHKFmiQpfZZPtpHsSdy+qjNF98Q8KK0AqB9NvEnVJt3qGpJFHHEVq1wqsmBuRDazpwhcNk54tXu
DNvcQtzNkiuonCBRWDR9nY14le1j0mBNUj3+B99EdJgfJD4+D/fAYb/00FgUS9+hw9fOXLX/7NaE
3r66RJF2JSBv1hgQrvMaw8q5SDYhmwYMyJuRkclY6STHsNragDvWfAbDoJ/uNl1LBvK4ZhEzm05Y
bzHagYt9y5HrazMwTpkixs96f5S2N7Pw8UKQ82ExOTZLCk01N4xBdf0JiCQIYKRKEDH0pOII7txM
JblvZImCId1pWdrLK+VqeD35HW8geUSyuHW8refUhbbiTfTYVLf0H0y7PYKzjuW9fWCZ8t1j6Kw0
870K1cD3/fEVMjkC05hhuQ8KcrzqsDrFnOf+UYwviJjSDtExpSX1Nn6UyflnxE/EkLBCnVRadgAp
WkmL6guCquA8zCvhnZIljyJHqnRa6CwPzE5GAGuR4lBmmoqhBgIJqij9s5IxdMZqwWnglSUR41gY
nm2CKgUsqV8WCUPRHPupUGNCmVZKHohJjtJCV090jk1T4Wasf2/3a+2EnE09uRB0x4K3zqSl2oIj
txKc3O5tC8yoS114462tOMWtflGgrowpF1L53z6VZejdvVhZu8TRU5VpHDNHf4UoZmGTmkXc4rEs
Yf/y+EyiNFLXckCRpfb97ArhcleygZNROSyTOlkhTG0e6B1meiVfhlQZ52lbY3lb4rS7r84+AgKg
ees3VurwGiMatWlE1JaOSOJR7He+5oVIctBtImBPN8BU8ecojJftMIM4wgZ00CVqMoxz+g3yYsUY
xJ+OuaZoV/pC8h8vyXyynsB9t/JLU3xQy3aWq87Jo8rO9mhvJlqIGRo7eKvoaJM7Xl9lbcRjkmjJ
ArCJM796rKWR114F2Sk7dFdRdYIDbRUzpB8M6GnoiB5pS2tMVp9vSCJR95Dt7cZIwdvY987V0jzA
ajSXrChy+mG2UJTTd6pNKXLaNxMPAjDfh9kvn/GJju/3SdpWSnufbOTzU+vfJHecYzPQ+YNKgjh7
C6p83dzHvcrPCDOYuTcSayB5Ej2uMmFQzwDdxUycVbih1brOaYORBQh7c/WCroGSZnMlEqW9rckE
8zJdXWZMiHU0IeMNECR44xynZ6Y/WgZccgAe66LeagLeAjVAlDVbtZXq3PCRkd3GR2YHDrzVFvIV
B0hUQ/SxXiJzMakITnbdiTDHaC64fvPXsnAfc2sVSlYU1A38HqQqbO93BtCjC3FDCfkWxIHWqtlu
3ioJ2mAPioNESxpAOXl9MXjrWU00HnWGdr0KxjKkyemBN1tPoUkkk5O7ueipVztfTqpGA1W+lupS
60JLFnq/PAEYKidcQwq6B+Tq5/2StTzS7bWeUObD/zJD1D1xCfI44wZPwPjNDx79lgy06qMOPpx0
rJnP+iJDUS5A2rC+pT+8M6F50qEWyrwKBdBRiLYdqA+mgRsU24nS/7jvrY3m2yfkEHODXYrrkX6h
texViVKUNgz7UZCAka6y0Znox7S45bEadIBv1NnAb9hLY+JtXDU3Suj1x9ItYKC9xSjCyTSrcwfo
+LgcDbsDtILPTK7YtjWBiS7TuiaVtXrH/RbnwoVsEr8MrcSXJQgbDQJd2TROlBC31mhux95LgnFx
tv2pWhilspfCMR0MAW0MQDvSD45rK6LOePBb2cO1AXx5YgtYsum6SxmHfD4OP+V9DkfzDBdjhr03
oaIWq41aznlY5nxfe+hFGy+nDnCceZjEq8PWjfV6/bAy7fgv1CWH+U94QbXsaGhr8SV3bBc4zqrY
ZRm48CZcSWRMA0mhlVAwTDj10UnRD99345AYmE7p22vTtbZJ4oODlZWVWDiHkb4ObrgkXYFx9Ma1
dtOt3zIcZQp3+lpwYeIryE0C1LlvkKXi1JMchWchnAtdWiFyfnnNqsmS1SJnrAnbeuSXnNkJgsfg
awSrSdTcjBs48rRH+dENdvpaZnPs+qpqww/rHy3OsVi9Y+Im4wNkPqiCpxjUog1O5dp1ZDrjtjha
xNsP4DiEplB6LWilfKZeeC8mGtbxdiyqJym6SlkJabnlWDDGZ0U3Sk5mfanZtNfcVPuYdI7dOSgJ
OUix/dvGsz5ZjDZmxcXHuZXXh0sJ8gRwEkYufaptdguU704NBPd6Z+X3i7WNI5ZJm3J3DQ2Vc39B
AAfNqMRBSCOjiSicJQPGPFqgeR50e64Q9sfMn0G9IjOEPTWlqfmpbtuS+St9E9BcW4z45xEasFD8
u2zmLNR7vRytnMAPAiuTFdselCL8GR8jY31r4p8dSSl0KIFmm8jM3q+orQO+HT16e9OQ1w4zkXMc
3uMVG3sKuUvpEGEdFeXJ/LHgYCIv3ENSS+p5RTNxX+G9k4zFGQX05Q6OBNI9BzQ9rRn6L2ELKg/M
AgTUvtgAvVInUHq0SPJxFCWTRT1eEDuIap/bCFNApjzwUB7UQnaXXmMwNyGCymytNDYBHzIMflsf
KxLln1XdjYLhc4O3oiIckbsKk+eTPfny///qBpDfqh5t3mc1Iw3suis3Twftr3KxTDhPDXoOZtIk
OzC+JEOuogQzaapL3XNihkrdVdAD2WZ+UERT/wBHD3Ae5uu2wVUDBB+Qu9ip0WNhCrWlH+erMe8R
grYJOUEShbvT36fZcUK/ZIiHSA+nqLieu3kzROfPX21sBjPPYixF7ihRmxjOYkJP4rSOv7AfbFCV
Xiwujnq+AD3hrhOgiBSVe0NxHsCkHCqMVuNdFmWMo6THe/5vA9FXrML9AlbPcZAE4HTJRAvNEFH2
8O2AojSqJDuaDeK8JYmdsLITA7H9UYaELUGxs9gFqJFtD5FcCTAq3+drI0KVxsfuUUBHmMbfODUU
o0i4lR6rV4xKYvuVUkmw3EneffSmrizv2fI402czOgJS4teO+sNy22rtSUbS2qtw2ETFn4xhYkaw
v8gO5vXx0tgeOTJrQ+7oOgaAHI2wea0BzHcr5W5TfBUQQVX6pU5iT7LDScQ0G1oKhEAVKXSYGVEU
i/gR/cb8NLheWt74khej5fdUnceH3xs4LTJ7CR9eoijyOD7XlsvwjeP0ib3mbtZoDaN2FFHIkJ9/
3ptqcXhiP7Mr1Fwl0F2s+i9aYcNz2YU8pWSYg7sESCIQn9CBV2ymk0dFoInxqfJhTchzLGRT311H
6R6nT2SVL/LVmgW5/+tTDxxP1UXt2dDQYLRLllcTlkYBufYWt0AG62TPl8+HqQZmGgXFYipSZZ1n
6msWrxA9fjwK1z4EuHFQPtZGe4njhwko978j5wFSkLGgZ0p5voFdJctU1TS7U5ZjtHn64uVRzerg
LwyVuSejTxDombtM0RnHLZ+PxgOLB19w2lywjDIEACoa/bD/l3VSE83+nUd2iMWetfBhp7f2TC3k
//RmLKmAlX35h7TrUvuLwHEkBcyVRK+imqo7HKmaWmjn0EDN0iO+v4e8qzthP9YuZo6hM3Ofk92P
XWn3G0kKbTBx7jAylTgR62DTGzdmZGPlMGO2gQhVUzP9zl6WdLvL8FHOvE4zo+ekYsqzK06Z59/I
3at8PwFWlsE/Mjom1aFCMRPMyqUiU0VZHxZ4UUFQbt18HJxXkVMg1oPbsUQAhl0G70Df+fdkB9z+
9okw704mVv9QkacTrP0VLRUVbofVrJyH6JbCVy1MASWzO+uy7wIIWp/+Yqu2YFkK5sXjHhtD82hH
0lsmEvwRg4wU63rL19BGueQG59pitT9aD6MzuimAOVeOtUVSIEaGuUf2EstMYE/NrM81WY+IXR84
PU7P5TcbQKf/R+HL96SrWys8cSJXxRqzBzI3mf6I3CaXTLxwyaw4Scr8ndgwl6JASZKasLMJjmys
j9wG4ghnja+UKrq1fil/x03Rc+DvVL7AQ0A7zwe7wCsBQ1HGx9byqV4PQufmW03H8In6wruwUIKu
2VLdO4i5mYo48EULAltmR6vkhB5kDmeIR63/hcd4+zz4OLfE/2uU25zKEOL9GH9yOjz/aT/dgupT
2F5rh87cADrR1hIBg97q4Rr6wvi6QEuvkXF/LOJShgAG0dxPQBd/b1HcqZKuo0SmqRlFtyZWnd1Y
pKdX/gz6FxSC5iOtVUuQbNgHYrzD3MaEScYydDXC4Rl+R2yRF2G81om/iX8KPTL7KHScTjPu5VpN
i825rDrv8pOH0qG6o/4R/7PdZmCl0HBTglOfQJypD+b5dnJtJIAOfVEbwLNIOpQge9iFG49c6XyL
LBJWlQxnjyPzUbzpAtRDGifizG9e7gPAqGCuq6KMSabnBA92xoOQ/utEkNND32oMB16vsRfnAL4C
GxdNfz0QtqhvGzvpl7I3/q54NDOudOql5l+5PXO/YP2LG7mvCrWswvXGwJZBXtY8E3RmE8Rv7OYH
YE2YOQnKCM32+CzUxoGdkVVSsIqwa7sklVzsO03Il+nCo6a0g9XvQLbFWIWvUK7d/Zb6O12GJ9st
U3dkfZbefm1181rg9iV0lIrJM+uPY5yViVOVDbHmKIhZ0nRtejKQiMZViGkRQodu/sEuF/NaYEH5
9MEYCIy+Pph1qeTp1PVhg0b9pC6z7j30PnLlNSlOAra7XmAvCruPMmf1/ehNiT9hxp4YJnLwnJJx
YTiFZN3St7gzJInQ/FHNNzXOvj7qtR+dimemMmke5gh/xedhbpgxsLdzmeb1faovgG15nYNkE/HH
ld3Av8TZK10ftCiZFzW2iyPNfB/+VyIiLb2CY8qKjUesQEppczmeregWi16KqXeui0BaM1ydn2w9
/MXZAUivGsnsChVDia2wKdFn9BmAH83aqJWtLW09ItTg/SDuvrVI5vKbT0TX053bIQVd148HsjxP
Pl4a0RSh49suzoYCSi5QzG/TnWU7MBRLIg4pNqIwXv0JdImc1OupADreHFSf53VHg+Z0lwlS+VYf
7Z3jY9SJKqs79KoZIePeWArB/q0NmZVPnbo7FtuwweIri6T6E1NvCFCkTuohf4WfwJqfaKnwb3oJ
yTIt/6oHMySaDxt6p5jTu3tcQ9HCwQwSfEKRdEuEtIZ9FsCrdx5/OcWELvYYqUlhEX+2tm5+nsfb
pCadez61InkcaYaaNB33WuW9JAXxHCu/iP2+nvWvNJxfl89sWzU9pTcMziRdLZPvIdFuBPLFHuJb
Xhmbp4Hh6DvvvZBngy2ePdMVotX4HavzNeFrgI9vysrYLOhx1GnuDfEMC5Z8SCn5hoaBZcnu8BAy
M0Blhx78hw5Sh2yjLHlgPqODC8HVOXv9rryjCKbWoRilhk1SsKEsaVExUN+1VO29dLNysoURtU7t
ehAXpGxOM1vCk1NBMPMRzVoUE2pKpKs4Ok7w2ei1EYVRIkRMd3frp098pI4PmetJnmq06vl6gRlK
4IMcOOtkNZjQ1qe1kLbkkc9dGebSNIkK7AfH5SnQ7ivXjF2aVevDUuS+K8XLpi/fereg87Pi5zxV
RlSSdpsPZn3PYNm48PV59ltccpRHCbbJSe7xWtn3VeX7BPE8y/b1E1/phKzh+N8VQgNSJwMxqqk7
pHX54bzkfybOPQj7DxEhBF3nmVRrdCup01lTY0MavJ8wmLBuomgzg3Z3RBwqEll/CwsYD0CcmT0I
SDq6bDwoPykPBawsH/pgfVGhIWHx1MmlnTu3sA5bWcckADz/a6gjKWGiaVhaqKZHumyHYfaRNR3M
bzvgWjp1BA5ePjIcSHmln33XBvIZjC5gIjcRAjuwaVw/4jTxMTYCfSuhD6LcaLFbmYHlHxK4Zfee
w266Ccsj1rttXzEhVH+lh0x7BAfPwsiXOTYjpsJ0TzsZgAiD6ODh8Eqq/d6/yiuY7AW0e4h6TlAX
tEXYB+1jsGN5s9V33h8/c5fUo1LcVLoKcgvtApTM2Pfm49b0dFyLAQ2a/GKaIKTg6ywiocBq1IpP
tHitIG0pWYuYyo6/DO+OmebCOdC46p+4rQIbt2HSPspA5IvZNDVJxapU5mBWzuvwVqNeuCSiM39x
t2iZeUYu4SnbQ8/g0v3Aafi5CRI8C4mDaTbkob3XJBnZv9iAujX2C4EuTzOYk60+woavWUPgbdNY
b4CtGI/7m2NSeSnhykB2XuP3NVPjNUyff0C5hmK4jYTXov7Y4HygZhlUni03/MrUvsn3Qgdu/h91
XkAPjhDsYND+htrzPepRCTRmS0y0ieGevArgVc0CG/pNynPvESgocas3DZkdTugl7QJb+JSZ4aib
uvL3XwBRNu9Gi+AJq4U76pphuVFbYQ6J2rKw9j8FnDVR2qsrQz3wex1Pp12Rfc9ucMnXfVbXesJ4
Ai5K493K1lxf2Pu1tRH3VRV3FKg95DDOTlEgTcrnl+U+I6th8GPdzvIFAtBgJgKMkUQ/pU8N7FH0
5psOIrNKJJd/zLpAgUolgSw0gjh77bxYPyR5DWGYOl73o1uEcLUHPGv1GMTlBPebwvcEpazEwdGk
80YFeKMLcVBR+VHn5+M/PjgOdRa+hvpENWWv639QXZc6cDgxnhU8ohWMmRJMm8XEIA0xxFNAlfsM
X8qlimXmd5GO+sMAUTzYunl8R6oxsC6tOT2wo/uEspD8IQR2yVYiDgBWHh8Hy5Ng0SRAqhhSN5c5
Z0Bb9FDps8ZvaO6ohnkVdLbQNEbh/VRE4t7gPAtb1tQseAFY3qIYxDv5h2Pe3w/9P2y+4sE0aRdc
xXpf20FZ/Co4afeDcSuxWsXafnPB/E329YXahBClpo4wVDbp8Mnq2z3MiqL0SGzcc0uMkKCw/B4H
rpTeB2s7tXbwGnL4d7B9ZtxTUBYrjHI+MUGRYdC+nHbGgfZHLKwVy4Qd2rR2Hb6b4gGGLV3oXJc+
mlBXxMx7RXolDBAmvPUZx1zLIMq/w6fM6JqGc+2AedWtM9jC5Lm/hJimv+m5qQPsUv5mrFB8JaLR
TxVFBe5V/HW+EHmZAamp9d7Y9Yl7uwpqs4VNKMKNYuEWPCDZY2zazszQGN4eGIgPhHjyQIWEhLNv
hTgF0bYSxrKD3siPQ+aOp+rdIb+WhwFEmVP3w2U6VVYGgdSwv2tTqHTV7kQnCYFNPaFjzbwIopSe
/kfXdOVaVd9dub4N5vgDw0aUUPVB/MdK2ti2UYApnbSJR/WE8y4wVq5sTN5zkpbkjieawosZclhm
/4hJnbSXRd2a6wVTw/DKl/sqKKGgpL+lfZjXZvUei9PhAoAeztX7UOCHsXnWfDI2mw0pUPIZg6ae
fa2SAk9ZC1/K5R0N3fnIzwfy/5+l5xX1/Gz22bJ+Qx/9EJGVvtEzCKS2Nyvo2aySWKy/bMHvdx8z
WsqLZZhhSyMBs49pNQlhoIcrX+EtrYNZQWMlGwhBMKAyV9Z9dV1zN8T8T1IvN9A6gbuibgZzXA2n
WQF0OMt2QqLmg/6umnavN74Zb8OHY5PZmuNnO8yU1BDt0/mc1nntn2HdpvsYlBPgCVlUTrn1fJib
NhRksGz3Tm1g1xk7GQguV5EYoYu3k/R7pvIFcF6bS4adoMfLxyXFJQxHLG9AP9pfIJdEORM62UIO
dct2xxASJakJ7NwnS3OBv/IX+l04nfnSm20eJ1D4p8YLPRBkbriILRzh2SKlcA0cpJ42w4jdgzg3
WUlAWoA/zrwIc/2wGZE0tp8244FK1AQ8TX+YyaNsA57GtIXT/AWDllM7Jl4OQd/mXwqnQOPrG21V
BxU+8Hf+5G6WwIHltVb4YUBp816yuQgki+9ievYwTS8xY466ZcBUa7Fwu8mD5uSS2lozjyUQtfNG
LZ+JbztI0NLWaPKxN/blPbGasU9dPW3ewysh6ya+6ajJv3bJmyETx8P9sWsHKjdwvADBWeOWhJWt
2bvKoGpUTv6YXiDnVCvrwgM4KUJf4vAIPNwiTwZ2EaCR9Cq/BHvBXGicKymIbE9qEUr9hKLzIjRP
20dNj5KASf9xmNYyMjrh4bUz0iGpXvMCONmlbpNb6t1tDUzvuw3dAbqaU9VuFp1RxH+L58+LiU7H
VE9XBKW3s3AiMt7vNsLU3L0xaS15G40KRo52gm1TD/sq1IJzseZ8JXPeiid+DjAQ4FeDmz8bJCCv
qWQ2CCfkMrbkX5ehhgMPLqDdSwMNZ31mNGOc5tAWRt96nwtjXWEMl81C7ZwdR0y+wyUpjycIHpOS
ZEmpFupASZGuf+fdSwb3z+kBwJIHsL1JgaxTLeRafEyCQPjSs7tJbckRWFNqNOseRpn8ryGpEwN5
mNbJTLDLfNFHc9IvjUjhDSm6rmP3fh6mnCa7QZYScKmCotpG7vGPMq/RLa4uS0+CrZfv/GTslxb4
gA8S7HpnMRYuOx5AsHVN5a/1EQhgI120x5ksYPZotmFxAi8TBCEICdEhF+4b4yhaSpreI5uvFvbS
FqTA6ZugD2rJ8zXghoeofkd4VFXMXeA4u79gR5z/PQZxi03TKkuHIKYm6tUCmAZE1f5BJ2cwEdsD
FaehsA6Mtvgw1TcQaCH/PQKPdsaE9rIUuTMMONa750gWVc6AHifDg6TL/hKDMiVdwhtusfLAhbht
KyjhdKu92QsFAzU2inzreQjjPsjDKCwdpv638+a15TA82GKwxQtwGNBAfXbnBQRHqjq1qBKLTQIK
VDvDn4j+N3mPFhE8JALt+ee/sESEf6XnyeqP8zLpeg3E2pTDCe68HYt9MzDSPRWBYXOguwFuQu9u
duTFnjcOycyBtjgq7z4EM6yAIv+ozXNaMQe59Gl7BLByUfbVb+khtmuxDiAMcTyBr263nI0tSax8
RNdvcYbcbMCoR/nelz0Eup0zBnHhdKPcQ91CnsCl7rZxIA09wHYZtzeMZJ1i/rj6vAdI2vITCH7c
gRlYpQxXWY6ypEFubAihOv0zqAzdV3IpvXKrJDqDKEln+ZhERUdrteJA0DiwpjxSl5OiqT9kla+8
/DsdAMXTyEt2ZE9hSp8bzPHUAADfeqirnhkgkLXF0tolKQSk/eRplUE5MUeIgHbU0LyjMjy2t7Jc
JWV/kEvyvGolGoGf35H7PO4P2pF79Uzw+B3UVkVTtAhEg8zaY+rQ+6kEsftjKtLMhIVR6QjTEExV
WoF2ElNNLjbPpDyMovUgmoprpuVbAUT0XED98CWhteb1vCWPeFz7VUJ3+Ytamq7d6FIF0IHJgINk
vD55OAqVq5QDu0fByFqjMYlkIpZvR2kqvhgNfuIm9264UW3GSl5qa6KnPr4YUVCl76RnMRYYro6w
aA7V1EsOKBA4fwRvXM+WPD15NBI3g49bW6kuULRs1+XbkE5dADb5D5IorsAf6Cqpgaa1htpJxfm9
2HysHuQMZQHQcjtmHaekadi6CSIM2CKkWULRMgSmzpPGgYYqS3/ls5yG6uxqNEX/rmMqsz2SCN7Z
RkXnENkeKV0hrN1cPqe7K6rfL1ckSQUGFA4+AdwDnj0XKjoyPTKEDXguyna1Orh1cfaDb1oarQ0y
R3zT4tVEf9QwNC0PmDElNyZM1pZQZk8AaQNVakNgIwfqan+w18KwBALKammiApPfbmiTHzW73wM5
lLIPSnQUinVKJmLRypAfY05Rm7pzZewx7MvWITLNoYjReUzO3THd8Nalv3vNWQK98MXyaT205srD
CSfYdGGzDd5NFWf4r9+7WkEkEwTm9CbO/X4m0habeTGf10kRSAMOj72tFJAPsSFUcEp47snbQOyY
zMYLCHV0BbWEDE7qW3cQ5X8drgOYVrH1S75BgvWvC6kV1hcUkypFbD2hcyMSb6EGq+//91hE5eT7
SZOQYnRQHaE5JO1oZlr1EIh3ET3uXLz3Rg2NRDgkba8IpO0Ynre7+vQzITgjYgcLUZu5cdj3QUpB
PkF4E8BScpzWmNWu0j4J0iqtL3gp35s57XiFiaWK1xGex/DxY56ZkUDImRdwXLD17GM6BFHj/v9a
/mqCVLyZs/623Aok9/4pwBrYcLiPvRJKgPBuP+5di+Jw7HWvDOjPvTbHEpmoU/6Vy3csxpcGyFhM
w7cpC9pevpAAGBumawxfx9qh93yZ/e0dR/bV6no2n7FX4cpc5qXHndMMpcE6Ivci5S8LLbcb540n
AX2wKXByJBNJumPTnfma8QRWtKCHllEltgupY8A1Lxkr3X189TqZA6/uyudy747fQ+6mECbiA3eq
EYYxOce7Vwm6bCiNvLkFkQtZrYYNP5z9u4OPTUYNebv4VqJGEP/bVKi1/K78BEVp3j74kz/aX9H+
IFGjzkCKShkVUMrom1EaifdpmKEGI1aC64GwlZN5qv68njGYSSqB+w7g9dmA1kRUgocZanAsuQIt
9AdxpVErqMbhJi05k0Z8C3H1IZ2WpZHNHYf7RLwIld3nT8d6QSKRq1DfMTpblLuoSAw1FYutjQKk
VkY/66lCEFvcLyLx5gDtLfIorzFuxBEVgGucG6ivT4nvbjL9ZNKvMBs8GpvsQ2xrtxeVDWsjuQqH
40Gv5lEOf0jIEs63+cXJiRhsxoox9dZEz9BTEjSJxaielqSXaTfbg8RLfzfs8UJ9Vec5lOpBl9rd
fQCKKOYSAB8XP6JO5bLFMvOAoi+xZOUa6z0AZxTdyeodktInfk3y9aFOSNNvf7FsVPdJ4wFENMSI
oDslZ47O5uscGGVm15I79OSAz/TpsTEoiy8VcT75rlwuGkY4mzl9n1qttJMDiiAoH59lUykgLmlf
NQx3hlVzmYH2YHNNjL58d2M3k5mtUjYtKQIy/9wWKIbR7ESVo8h9xp3PfznoD7fWWw0NVoqbRlNO
OVFj7IdZxmJ7E9Xmn3QcjkpcLRMdVGREB8h4vGhErZKzxanhx7qDLXl7J+aPOahqEu9utyo2RGbg
gZszeGcRJzB/lhDLMp+FmfB0ZP7M+bUg9gl8lBUQzwCwSFxFH8wkgmbRkCo+h74l3sWOlSKd5NUK
mZMbRmzzWEfwCTQt0TslF+fZzGBlYF9DFhPgpB2xK+nuEFQqeZK1Z71p3wNpA9mdV9sFrdpszzca
G1DCRIIOomCBn3ubHWJMgWzjTUTqfwLzMi0iM8zjBwi/ISoNBB1apcj6Dd0Cpz35yvva5Hg80xzt
xuLsQt0Em2Ha6N4OTfSy+qvgJaY082qJXKHj5C82R7G/6pO3mAoIT59J8Hk37RsLyAcmTKl4MzPw
5XaiRWDllj3hRY9zGLG2XYot5+0ZQDXZJPUi94ejIEWXRkxzCaUKliCn2pEepn3Xmy5VW+ReGFKh
FUNitgbcA1gLobuJhNiP0iAdqJJ1bgFRyJO9ZqiPSGNf5ULM5ugftxnRtqhW9Kywm0jNaYytgpgU
l0pgV+XgRLgs5QqCZquII+Zjy4H3l4J1TGhPxLy3Ro3qHUTF0ec7HAWOFw+RQ60x3eR2q5E6SXEw
MKdEYVIepFOpZL8XerDzIZ2GQ+Xu3DfAs+MBPdY80CvcoFf6KrosrpWn0bbDQcz0OR/MOx6e8moo
IPCnHM1Vm3dXWw34Vahe09DtgoWC8fG2W14df0Un09sY5c3AUYF2PFdV0CnLfsy6/SMHP7y9fPe0
lHY0euYeBaQU7jFyulsTEarI7t8PbDg1M9fHcQ9p7yVWqChxAf6q9z9+inYdt3pVxf9yqfGrP6GC
HIdM04nRphB0HccqsQZx1JyegWgNIpl0U2kvIXFuCwSpb5i8iHtfw1N6OJRU7L8I23Zkce9U7uAI
6AvtchSfoE6Rs/ekCb7N1ecr16k3KduvEw0ahuFKhFE1gJwXkIDw1NnZWh+McZwTxYMjRqFRAmch
azZ62pvatCtcQgnp9KRk+vYpfgmDF8ojs6gzSXtpjOpdoMmXqrHiQScSngZhgLgyemfql5EcYdR2
wslFZuK1eaqaevt/qyF/arVRHk23eIec1F5Ov59JRwnsE4onaOauzS+cA9UQQ0cmPrTif/3Fscur
6Xa8npjF5V3P5Y1asihq46IPZK4BYzC5raCMrCBffa4cx/pOuiWJIWNFJq7F3LCdtEZjRSUMzoVb
Tzd8ZqyBNOoLQzDLjwOlpSkgd6F0dkrEVieB2Bxn8ebvhqpUl/Iviu93SytAU3fS0C2IRUEVrw2Z
vDMmq2gaMEMUZqoVqLwz736OPMpXM8z/OeQEHbs7lDMSg8Gkmi44Rvx5IK+KpvxCYAq0myK4RdIV
4W8gzAOjoJnDrncWPaJ9TRuG2tI+Y7SI3UhprMAVTzDK5IvA9+Pls/PdMRTNUv20l6A1DesRUgZx
nZcvQRqudbzP4wD/wzSG7KPyZM5EnofnDnaMzi1FyM49/aC6GxIYUSG7QZrxQNohC7QuqFpTq8zg
AkGq9Objx9Z9fr6CVMK0rEm2JkmWT9i42+EGwQfTg6G42u13StwlQWruEto2CAMHcYf7PoxwoWOQ
4tixJGdliEbpYHG1JCKUJxdduqBhLRpYmT2SZvP+bzXA5i0e/DDXlN69ZDv1g9DsDJJzMKOTOzWM
07aewDhXFRlolEXIkxB0aiyqz3w4aQay/FDHCkyi5jqi5klhdc5JX/B8x3pk8OkBt/MFIweb+was
dU5+BVtk0oL9TmiQzzJ7hw6ccw7JxAdYn/ru36gKZlpVlyszIoEdHPPKg03tXSkpSu7cejuzHDZG
nYxiKsExGfuHRfGPJCH4aEo3OIWdYKCtZmM7EgSxX+SdDEjCehPDjtTLl70dZXYdmgvTatnsXSG9
5vqyH+3ardbynKYQVAPW+tkFGIBxmUdv3ec5TBnSsrBM0yxTBP8aDXCbA/R19Vk8S63WsaV8kif8
Hc0sqjLzg9A610SY8vJwd0WDa0VBKk1yDU9xSTK8VDcRawezi5Vp3EhOxgLoI3y+33EK4gd2Em/Y
4t4qV7zhPgct+4mArwz10FBMQ4i1AZvaC23tEjKEZPCQT9PTcW7TLosgrxWn6nWnXtj9KpTqOZSL
8QJBSyQy2qNDg397lmReLAacyxb4sE0OxVLZX6RhO0YFB8bdaBneZ95RbGNmeRVXQLE/jAQ1WJCE
v2R7hD8toH8DGVU9eD5rEqKyBw1Qqr+cEB7/uPNgLfChpgLWwj7wQy5efN3lHEmkD7Y+PoMcOgN6
zI59NAkB0WsrGbvD/CQ343xYFSKRdoCb1LObNJIAymrfSQ6aDxiiL4upYno1whS/GKNn4SXV0XQt
HuSi0LesK6Y+PBmnrxegMwv9R1YsWqgYpnezbd0clyQExorjIpVY/bkcpOuDBOZDAFtAd7OAWhXY
PQfvnc1alf5Sag8OETRxDKweqqnhoJ1U3jqjAR2rCueR3frADOa8rsYUaNrLt1HmW7K7XhgLGr4G
oO4BaDHWGwf8JPoY2J3x7PVdtT/fzYOlVXXKd32I6OwE/e9BuTo9FqX/YPtVWIlRkL96vS4EqjJt
f+Uan8r+MbQONQnj6f/FbpsxZ/Bt/v8kfiwp2UOrcMpGGa0grvTzMQarZV5LuSyhbIluIViuw6Vn
GqSaNcva6FWUHHhKC9Botltdmgd22np3gwUqfJGnbQbgPBY9ybsAAQ5rgf/xbJ8ptz7AgYCNXnyP
nzkNmmrvvkxlTnVLkwoYZAst0Rc3PCBHqXsk6zXTwYSrCON2Z5JqL1sSA++vEBiqmYQQ2pmzDSmI
RQVeXAG2EhC/nqMkV82K12XiXxHX5KrTWHxUkHl0E+8xbDdZgB4khLF0B5aXFz7mpH2vKnMUWt7r
W3i+Z0aR8932lW6a6t4R4sRtUSOQcvJvQRX2Nnj5KuwKj6jYY5Cvwytm4q5HXdIGRa/8F6mTxsCc
IbYgg9KzKkLc54KD1oSY5I+5ZKfndjHvxOB4ZaqcvMKRCe20MvMV5oIBEevsZzh5fbHqLywXVeFw
FJ7Rns2zLFbYg3tZC20p8k/YaJonRVO0m+fM3+kbVhpmS3lO483rjUvFyU/z7Ym866mE0SJ60lB+
4X8FkuVWOdNdlb2VH97X9vPfcHrIlsYjWh71wrqb5iALi3BNOw29wKKSaxQAWzumT8CUOdJ7mi9F
08W9sLKWJHostGTQaMQoqrKeaF1WLPvKoC4B/2RyIKXm1++f2YGu1p72hJrQrVJz526YvdWhccRn
eSyxiqTD7kxc+AXByu4e3gZLK+Uz7z5hn+74NPstVnSYkMEwBCVIDKSYM6SOjvlSOgHK3XONsEId
KqX9iPRbCUnD3c8KEQfuFZvCyx9EMnTgTsl51kyF2IAzyKllUIXXeSK9Esi0DRRMl+/uFA8beotB
o5XKKT0GTwvVibDh4DFEI1zEIyIKbN96MXVVdHdEBJXGw+Mz7ECMSDsmmxQ2vE+MHHrpJWMOAIzf
HZi7JkmmpJ+DcisF7U737vh0/SeI6VVmBfp0/LIRZCw3GtRjH4wExNYIEpT8jcE6gajUozBlbmr/
NQwiLpfi4mvI5MpP5KGmqrWhrBETfy0a7JUrtKILdpM9K0eFfZriraPp5/zfEVCwk/R1957wPTIE
esf2vmrQwgtiETHpXDF5QaiB2grGMdxTPezFIwsIFlOEhpq1tiCs0BsbDr335esNR22Bcb54a3Qd
lCy7M0HjdK/Yw9tHRM47QmboyAISNwOLqjq3nDEKfenp6KJZWcTkJ91Px2zJjrLN0+GERdnfYGPS
agmSC2zipEh8iRPw16rge3NStZKBV1ohmTRbB1popU9Qgqaj1sgWDhOfZy8lwyQoJDvP0vfkpVEV
sQlVmmnksYUvEUox93zNRsrpq7pF0IMkpXC9/i8RB5VIjQsSsIWKYC3npOWWZGoe1oB6MgB+GO7C
W6ncLCm74pYbG+K0l05YWd+7FUFTXGLqmQy0wQ1qblERsBLwT+gBb3zJQPDi8Dc4A8pQ3uNmpRg1
VY7hrHEDcsyCQa53YY6X2KGREpMpIPO5vcVqc0WcVcJNOYzNuflQCKqjZFJnTtStK7TlpfisuKul
gqb3w5Um1W4TNeO3gC77xjAYDYgPiNFG7F0u3Md7Ez1GHKFtyiMlC2dFBZW+VxTGzLx/T1kSXNsP
nbDWx9nvTVXl2ambRyaQrHZuvkSOc+NnZOTZJweJX6WDeYqZOFwzijNXAM2ueA8aY+ssN0ovK1Gp
OF6tIt/m8pcQ+E5hYtTRqs5NJOVqlfK8P+chLBwR20Tenb0go1EDQAnmHC2svU1dHuhXGkCLRRHc
xkzkxrk/PiWKlDuEHKZ2AC0bVP7tM2pvFfhXTTOKfMDmu7dkJTHB63VpGb3zmQW+qEw88HFzf0BN
7gHoHOiBerl7kyEsRdmya4M4NBfSshVOPsDAKkxhhvRd4ZnOtr1DpJzBmrqM5d5PLEazWRmKed6x
O+lO0ITLyeeppwx5eJIn1UneXPFVikyRlMr6be4vz7WLzy8Q7kOyMxz7jJN7Q0VrmjyKJ4VJ3T85
l8yZNxUkjkVvh6Td2YpnPLAylkXH4iSkA7Pc8uNim8tcub7pzDAx+YuTC1ksOml3ItxDyj3qqUdn
SAfnVt91C3X1QkvOHOvX3wXbYZXn6YGf7wMoou5Tw0JlnNrq14jNRtVy2W7qte84MoRSJtsD8t/x
K3H7R90QQ0Hlqm6V9DjuV91wsUMqukFND2m7n6rgK2ar0sdeAk/63xdFi86izlKXKOxDBEOplUn6
hGndROiPGRZF9tlu/vdRoQ/p+Vv1aSsb4GEI2ezlBOAZbB7u+qt8wW1JgMIa2m8oNKrVqjxxfPi9
fM4MIL7xlKPUvXU0gERUO2PyaAec+7Z5QDzPh8L1n0TNvXkQ8z6ZMb/O5zjb0W4rXEE5zZc4ItXt
PIkn7nw1H/TMxMefp3rEENQ5q3CQEhWW60LJ8A2yg7MjVSD6xrNjFr1+EB8t1vgU8U3Aj3ji45JP
DYaK+LuBrbq+6La3xvsVGKBUhfIDsp7tkrhhUUUk+WsxyIsaZ6Xw7i27ftt3NttXXdsm2xHZ+PZE
npHkzYifDAUKNVz3gxCNWt7HBcvzaRLm8Jy5bBt9jJK7g9SgqWvk67eETKbhl5uCJfo9XYwNII6o
aoroJAbzuOKlyPs///1VQyLelWxDnqJyqbsOjIm0hsTAqWQ2DdfbVj+HAsh6cK5e8wIPnlXjC2eO
JgYrteXHFsgVKAiDppluEWG1mJzG7Q4lLhCsclPdDvowXsPQmXoVk2KnNM5pzQx/hvK8s2oxPOFJ
7AAIrAoK8he7I2HuPwcuxe3JXgsePCe5Hbzut/MCUzf4P5uLOQ6Vm58v4od6l0+44ffjfzy2jpC9
EDB3NXAXb9uPths64lnPTAiXxsjh66puoxEs39psGZdG1FK+3fP6TORG2Gj1R//EdfwJjqK4JFeI
0Y+tCE5ucltn77bdNt4RCFGRqBbfhN0d8JL8o1m7a7xHOOFjtYd5NN90oHWPwTz+luDw7xlueLtJ
SsqYXvXgThDDwnZQG6H/R1qYIsTXtWh9MPTtU7X9b/51EWtEhdccJvQPESVt3PGIRSMnPpXPNOV2
+AsqhljKPUP0HDgPmWqZIoou8pp4MZ7qUOuAS/rttKToJLHDOfkXrRjLF7Pl78/Ljgm9YqHspRme
AS1NJNgrCgVEe9H/eyCanGfAdHVV3rRr3Ou08g9BRWKFcDQGgdtHyliA4VMm20MoYRkrF6d3NlyT
sqfDp3TjiGdtdIOMCq1qAFnS/GMYV3MBXLMDAwrYhMtUnlgTTo1JHHnWpEy27qG05YPX8CLeLBJz
AeBAPSoDMjNxq+tTYhogdOt9ikwewYHIRPjODx15v0o7wypRhzpDeTKRylglMXFePawUrRm/lTw0
qlMpVLDEQMZa77YqDmQFV1VByMmnIpPb0/Ee419OyVDbwpR0J5dne0pnqDMe0TycyJNsSwViPz3e
ypSy0kd9pDxStGtuKwGS/k1sav68u2ksjZ7MN317EQQw5Cwu8srxXUY1PymxMFtGTBVPQBKyA95w
i97Difrcl4ZngjhRjLvrs++JK1/wOkOWB1sj+sgFdGnMs5kZAJ/T0EVVRiiUXyTHIrpII4yth+M3
rGd7IT08ZPxzZJ3WjCLBjTwwkgB3Jf1eKoHHbhdbMTrvVJzBk/CkkBOajmJOyyAmv6X23hmdgiNF
U+heIgWFW7M/JKC4c8QmC+2Rlv02PAMv0Mq2IpfdRQ/uA3rAnylO+k3gDXOa6F3U1pFc6CzbHxaw
ouTD6ruosF4zT0tfecaIz9znCY7WDsT1ksQ9UVQYXrnSj4fCkq56K9jx+jq4WoIyKN84wGV79FpA
CYCIvv95HaylGSB2jt5gqOj3/wr9BvY4fGo71cT6m2qns9oorNwhIeHzJgcTSou3dpBnQcm0pp62
ySNxrcZLiNSs5Yo7xJS5BaApms5HpB4ZLFjXk/Dxz53yEiTQTMO1LVNke6KU7cYPGuiMVq+3Y/4L
AfR07HyL7vwbTFGMYFCK+Cdv4DFFbCi4ijRB9wKsFpFp4rD4aJJU0GvMEgqWSKE1E/liPwokHyO0
WEhtzTSIDhIQgzdg96Qyj3NCFRHHb+kGnnbEkgt1ynw3OMUvwRbRv2AQxzF7rvZO9RQ55Zvr05ha
sPRucEQB/+jYYrWjhzA3aWJiTDj6IObYgf0TYS6t+mtsX/3U2GVtzldMEQegKPTk19lQSmHpIcUo
uxPlsn6F+jXljJAFeUrPIZ8nRjudPQO+O3lRtXi73nGKCvdAuocsgFxtY9QHlVYcVbzSrfWbjTUC
rtF0PMRYuqjIu+2nDLIgV1RrIW7GthBBOgM12CQ8D39UwtiUzYARbG0ZFfPrPXVCRORbYqMhDWpW
48t6gFABQBuNf77QCXl5Cr7JXhOQ4hrUpu9h9xZajZc9ivoXcFfzvcUv2K/QPiXGmYqP8Znk9t5j
cZcivAAxq+BkiBEoSQthJf64t6rcP29W7LcLXHc7NCz/aXAb9Mv3gHMHtJQzbsWGdvsKcJG2Qp7H
V7lARkBU3r+Hlr3yzlXT6xs3wv67wM/1BDNXeTr1xoT+OBegJZRM9WjrDWJJvSeG7QoZGm+VZP+a
fRk4sSiqsaTAWZgT6syBJsqe4MrHKlgPFNRmuS8PRAq6SA6hDsFgp9FC5osNFhgicZQjEwNdksEE
6dVTTt2gr5cfaRF4Pkv5szX/0kn4Bj13nOVvxtMLdGO9WU7YcbcINPBUYCqQsPwiKy9beJqce8mj
nawXmYOlIjiTxoUeZvLfHQ1BO0FS/AJYTfL0zi8BJRKuUrG64m+kEepEmHhx7xpWHp1Kx5u7ROcV
vDsNyMe33GZJH4bFuvCQJHvFFlFgvc+SeFtYAQrwAJZDn7GGf3Oyn/RzCpR832OUoRpwamb4SR8+
Vg0qI8tZx9xz1lkHo/U+nsWeKsUmIn2CNtwwMMJmu52CM+qAOKxcBeCYcyURxMwFdRwrhlKAlklN
rWuqiS38cHsksosv4FRD7i8Gsx/yzmMbnD65ow9OtUaC6TDrWV3JYNJLfRcL0yBT/tbcpYsb3ZTG
xOyZMrVWKV3DiJj2WwzHPAUr7E1dvNRhlsdpmF1hggloJGZUrCrupQiVt04IgJKstER2drjjvnTM
+kYfTsQ1EGDEIpw9oNyUciN3WcCl7lIkw7ZRuAniSm6n3AEn0S6J/ov6mgzNfIKEwX6PT8oLNnYK
eNmwVg/u6ePki0bX20fmqu1x1WhTIW+w5w9WLgRZozrOBYftUsuM/nuFi36oN3vvK2g8+4zOeimC
mUUyuNhw5h5ZHjctbcSOGprbcWehwUhTYukw1nHftHXd8cB+kEl/oi2ofabCemRLA+iddgVdmL0y
6VkvEta3SomAW5MERvPW6p4IberNwRPuA9mYGPXGsmr4epM+39nkxxlz6+I0lytMqhIawvGvWpU+
EpiOIE3aueMfen88shlOYvoUuiFdp99KqQfTZ3TsdGlAEHd/io1kHe42Df09FY93Ou+qu6Sko9WQ
GqVtCvh4NSZXDifwjMzzrwjPqCOsCKMjjPsm8LL70iLSHvHikho5cqlJKA4tjYZslSJvPGg/ZZI7
KsVd6FkGogCJ95pxGbFQaTKdu9kCFoYBYl7PoZeE1oIxXhZQ68sXOCPBZlzPG0DNcyHOlKT10Y4R
tBxMoSZ075DL1xeuV6jffX5Cl0FPdnEC/19jDgjV1fKcUkxIhd+FAWdLlH1vNUmEJ+pIFoC+iem2
Iy6KiMQ1+9qldOxg851NYpWB7XY7HLWxNYOVVfgNr7tv6WwIbpr9yThlkT+7KzeFYU0bVfOTN8D/
7gKJu0Zcm6ecmiEE+p9KDYeIDJjnPBsqqNC59QZ2dJeutqM+AQxZUj0DYCCVVApbpi9OhWCtGuY/
Bq5LXA8PMBOziMqVVugVawbFcY/vGtUMoQ3zRrE1ntK01tEcFatmELpj9nTo0h4XKlwc/Acyz+aZ
Kg/c4YqOQJ2oBFmcGfXxbHCl7fatplJM0oQsD3hHNjzFzIvf8r1EP/CEejsaQz3u1M9naUd9Lrxu
7ku94vMZHJm6J0expl4/eTlnRl1UFe31nTKBaCpJmjJuA1tTTP06dep99JLf7YGGPixEfbqpC/nL
Mho8onn6dRmqOSzKi3QSrYxgNTIUGhR/ZVZfFRkG710ZroIDcKlmRfq6Rf1G+XnGweuIq30gPQwV
6WlGePVQ4opXFAcx1QBCQuXv3AwY/q9IWgfcd2M5QQ4Q/rrawLePbATWcAQXXUX8UDoEcBHiXSIf
7cbeXOt950/4nwHFEendEjmjIzt3d+kZ/FMvoLMuw+ifZBKdqgjERIrgJgPKTwX4LNSRoxN+4Gg4
bnBnAOdgWyw0kohTeXyzM7ankjSJO4NmPqLc0YjFBfJ9REgNYm/Nr46UTBenrqINzOXsaipjQ4jQ
xhB84XfFS4TY6Uc3qr4LsLKuexCEcZC2n0aB1ONUxe1glGTQcMLssgvDA/qoUWwRg9L25efhuP5Y
v3eV51PCz+VCuvOCH2D+NBtT7X8XgDe+EkYkGvAmrUKX6vHLmS8U/gbLnno6f0NBmVd3FCbJAprb
GkS4ku3Tp4hNNYZS4cJ8mLtsoRGvu4eqq4yIGQ+UAkB7M7Bnebi+V4UtgMImtY5H82UlDyy6JnUZ
O6eAYEsU0lip/OyhbDcMp+EjEWH89sUoFPhdZgYt5FOWE9eogThgpP9tlVnbGF8+5bxublhyC1Dv
kIflFIDjbRaA+NWaJ6VhbMHmhUl6wp1ox4CdNt4sCCOjsBM10vovPitKArP0dcVJDpLnranuoIx1
cKk2DvsxrZsjw4mRp3X34JXswoxLiK0y0FhikyiD9BK+Vvz4XTCcOjqCdHgTbIvlNDHObxnyACrQ
klj+WJ/BHqUeUosv31LnyqqKwrRqeL2jkockUlrcCV4Mtphd+pbinf/siNi8dLCiCVzExvU7j8wm
RZM7LFX2Yrk6xNTTDmQeXLcEe3QafjctcOGb/LUvlPnTNbrJk2b/j9ZIMNPaOyi0jTlKpCYdz+3Z
6XToFDjaIdO2263MN+pY+DlUHqFHvZkNrevdi+ZTvwcsTtMg6oah7ivF1oz8LOck5003pbZcAXKe
9m2f5CjPRd/iDv69RU/GYi3ZSnn0s96GqcnQWDs/JkripGl78+qNaxSD44VkCRQUu4puHY6oH8Xs
15Faa9yIK6QB5DSCBozG2vDDewmQnVaHxS2+DhuQ9BkktBM9SYxoiU3dgZk58iv96FcXSoytePxK
rNN1Pbz5L2wbBcazXLmFJ0UVg4lWFLsnFWpPdCmbyRVWSbXnDtsiBsU4RY0iRNYjHOcOI8V3CZpH
MgaNdPmskP+sriTDGMcS3oczWJzNPUYURqJkLUSmVf6inxBqqfmSp+mM2YEKaWLNTiS/qtyXqa2h
e0wNc1xxnzvlJoq4ePybCDbPaJTJe/FehviPKILu92q2a9JTeMld0LFKsXAKxcFcXuOVAptV2HFe
UCbmas/vZw1PaIdYfGWB79aLfsjk3uIdBwyp9MT2ETLPfy7qGLYeLhUxjaR+TRnr+E1eRoZb9OHa
C7wdjyUPvLl46SNMNWhf2jC28/L82N/fOPOD6ckUezjoQTqvGcEr5Vny1Aa9TbPJaljekz+wHDXL
JNzz3gYTiMgfSg6TdsruPvSQHqIQdkXL0CSDAbv/0SfMl7cB1dSMaNC6JxmhSQqs5X/yoOylOfOm
8GxYx6FvQic07BsnqH3VJrhxsidvNZSQ1Qxurpgl/GE72p1avG+odzWcz1ZA0OnA4lGFTr8nTmCe
Th+j/v4MHAHJt9nPzWpFhuQT4KEel6ojHlI19mfsskFSLjqQRKcaGOV1zt/5gI4Vc9cUxngU+WEl
b5iWZyf7Ix5lTFLdC/RyUsvDpNLMgwL+kxo8OCv5kViZyyUl5f7fyclsdBjo8+EzI5le/3rWMwO9
mkZhhoT71nhHCFaguTO3cYP4jWubvku0WpjxKb58M1D/9vvx++LyoLPqfy6URGlg640o7O4MoNso
3aeD5f1+vvY3XQGt4KGOe+0yVmq5OvpPTp4cmkCJO2P2Tjqha8E/BduqZKVH3dkTv2oyx3FfVQYR
FGTp7gA59naJjsbGQ8LF0XpuGa056lYtGU39+drgLffTeNr25M8buDVhFff29OCVDk+Kp0OhglbV
ptwquYWzgljquYfN1B5EvM3Mjpk/vfLWci/JL1SHaZeimcrycNTuum9FVrVyNI7OkpMRtNonLRnn
ZI0HF7yqqw43CB7Tt4XOG5sFpEJ50Lb11fihVT2KdptuT8TYTiVPDfOSdiJQISSfMLDldukAfRjC
bLOgkN1TSjrkcBofI2YLGV/ANNhlEkZIDfWN+XowF66hhWMG9DY/+l9K2xAyroLPNMpuhZFTivuR
wfz1F5htr1DK6mEfwfFt7lnNMPRrs5OZk+LLxUAE0bcCg/kqZpUrGtZKbmxG0Z8J8v/ovoJ2L+LO
vDIA2dvht6M7oecwdX2dY0gj1i7P1VPPXusAPlIIEo2dW94gG3ntEF0g5ku1WCjbAwhdOxCGIEJF
N4u+ABjVmnKwTz951eoFmzFfQvuPUVqF/MOJRwW8LU9osaUrHKR7wNm1isshkKRJECGEbaljhY5d
+2y7DwrV41WFKF47mN3AMzWz/Du8+Hk17Sz2DDWsyq+SUSDoxJHxO7YgEVJr5nC3FRcLRVFa7P7r
xNag790mso27zDcZxHCrSJyvFWD+FWNUpXI0VNLl8rHdLycO/SzX61CTChWDXR/OmLVJbpsi+Wi1
Ja4LmSIK6q53cT0IiCWbA6qhrStadxNRrCzgsFMHbA/8Jfbus8yNheIXo7j14MP2pY8X/2VIum/O
u3A3e3nItcERm+0OhY6zFYMGKrktrrHFwT2/Bg2gjkFvhDf5yodnpZ/ZPIayaimlyZg8qrLet2ev
TuoQDXxu4T4jaOjbrVH+N7jW19oJxEcRyLe5l6KFsdBEK1fgFZGfLstaSJ1YBoyTBo3otMBI4CFJ
L5ZoaEMAGuhSqpPji0KFw8uFW1QEX1hWE11Z2ZKfgdwTN/vt4tdNRmKycmDY5LqhSjtVND2EFfIG
kKdD8tovwSl6+J0uGIsohqs51vP4H+AwF/yU7lzhwbjHfAheBn8JCaSH9/Qzz+761OL00h+IzIRe
d5NochvFvrSujdDMkzGUoCIJBcVCICNyCWf9vIc8xnqJUYU4/d1gfihMYLDWdmDvy8XnniKqpQVV
StL3ovb1zYs4zSTrxovTmu4ZTZ3oPEbW7yMx3oC2ItVcnuJoWn9I8epkAogIcn5Rw4JR/i3Ihpay
4wNyxFezywMHDKCnV753HqLAkKTPPx+X6nFy4AUn94C17lQ5QQ6y5hpBe+iuvfsDpaG2IEmikUy9
YzSyQre6WmaDf0hnx+7EJrpqjUEc6cZfnTI7gaTIx+nS2bE3B9dhg4tLCacf52xTbE57h1i/E7vM
Dk7Jyv2LFTdgbQ51O9cdwGvhYbKi1oByRlY+nCRaEly1smGpUwRVwy+Rka68ST1fiFyFdeE69KYb
hawb2EI8EMjmkMQ+DM07TSBmWydTAPSsLbgMFikmx0A/91h8PkNEOQSnMRWfr9bjXkmwk3TddbrB
urcD1MBfqbGGLJ5ZM7l/MAwhvXOQExpV5/rrTj7t/+bR+5hbGgoeH40kL3S6yYUZxA7dECEjGckf
0ne7TCaCuO1oT5ef280vO7tcYzm8ezlDXQofaHhgPLkAQwEjZSaPgmSY/304CA/z0BeSBTrTfx4D
qZaP2Tfwel4Gmjkyb67b5/G9h3qVV/WOv2+/p/TDP/RWfWHAS5YpapkuuyOhxK6z8bS3DAT9yIQK
dkaeEnGjbyDR/12aV9ZemkWdVABVjHXO91JOW+D8MB9MIVjoXDn/1KxoEbPLDgi3xmSOS6F/AbOE
F3N8tzWIBvP7MyAPk8z5ZqHEgl5SJFtmW+/x/svO9XZxKvTmQfLdUiFhr44w7Vd9SxrZ5Dfe7EnZ
SaDvFZIms7T0zGkfk32708O5nHeZ3AB0yF17QdMwD66et7XvCEra7V3QyRaOaZHYt1MQlbssHPKf
yEMXq/l+jbMkdGiz0pi6S3+K9xyeRxAmLKesWNw24b4r1stg/HczMuaGDyT8LgIYwlmZ3L/AYHuK
yfb0zKKfHQFvtYB6wWU2o3UjYXTaS3DvqUXDHqrtN95ML1s1ZrJKN9DLhLu4yH8WkDN4umMCD7oh
BYMolUkkXvDjdsbYJbn9/JB84muglolL2am9/ms+s6moNcGqtlLlPKxqX1HcQGTfaEAehPXY39DG
5kQkjiz7qPkyPUS32Z99Lu7pJCZ7cOdR7bk+XnVSl2el6CkZxfqS1+h1P5/15XH49UuIiqIG5xId
8PN7q30lq3WJdr/9bO7jVNhDpKNl2ciR0W+xZDSqw0SKUR8iQAR3Q6laK8TQGwgqli5xg/yNpRFZ
H8Gf6I1W9xztIqLmyDKOG/BPgXDfa3a/BG7y2CZi93ggFX91r1mrd51VQu7PJ2MulB9sJzDVlrZ6
0fglD8B8sbOeNlXsOZ/fG+JHQ+/8s9y7aGxqxaNMBN9OFWejwj0cRI+Gil5I5v0IBaVbmMtZMbQL
YLTUzLSnGaVwX96+olvR81ijc8CSEGaldNDecgVQ/2Q5BeUTJ6PEVQU9V8q/Qjr6SfMAUF7T6l51
yH85xPVecf+rzeYykoq686hv3F7TBEb6BxgJnjWViR2LeiZDXsZfCsyXWI5jOIYXpCyHU3o0KwbC
DbNw9hPuIYWCrB3K888wqSmmRYPIMLSRiKYcU8VMmkqAEEycYiAC+NqBD97vCyS+/f6Xx3h+ekZC
9welJFPfsTFkIJNZ1CXzFesYTXOuUNYk8fwr1SNyAoeONAlXU67XNTml6UtuKB5Zo8jIp9U+g/wT
Jf5iTHUo1I1NlWW/rHPtONn2RG20RvESdxjcTMtMWT8UsLb1PnR9MuaB+qKVtzfL844PXZMdpkUh
bhgbcS10NV0UgK+eI1pMQAIi03hinc0ziYH8gRIjDkT65JtrX6GJH7T7Leaci8P4oSD31V21EVOj
3I97pAyiOQkWfNuJlmPz72pOHh1O8JB+nfnJSvw8qpqv+j9vXAYiKOFDZ+AX37562xsfxC9OMdGp
/GlqdN/VwWFnvm/vyW94Lsn9r9KIsdH8EtqHZH4i/w+lmUYmuqgl2D4F4PP0rCd8v+HBRHO+dMg1
3ulKoCh8SXwM+9+7EjIL/2pKFmRZ4BTo8bl8b7Pyb8n1XhxMlf4vntkkYuoYMk/sJYgiBDQhhFWS
aQgvtaqMS/4SZs8zAhlI1N7WaRPJqUF+2IkBhh2QjlKsTJVvT1vDM/LHw2YH1oI/C2O3ru/+0VhV
Yb2DkBbDI9itWF9WbdiclxYMq8oN1YRIalGbN5qFaqkdz5Hu735INykrh9L6RffiXUly/M8ySQgF
neJdzcDM+JPZsehQGPTJecAm0BWXAF5lBXSnmVVRNhraOF40T7/wIQfZU9fp3MAt3IY3QE/8yefY
8KCwbZqpOmwQRaolG+z3AEdilDGyKRgfvDAlXOC/9NArg6kYT+hBPt1EI0s6vSel/7MGABWpzY0u
55db2halyYLjUdIH6rVHF70F3RXTGrePBdvQVwKf2CEGRSf3/q929bOLkyt8hOwkT+YD6JUMQnZa
6oXMfQxZf+mVXQYTlPHxB6PGx0hnlEqNGK6H8jtpaPXC/7L9vgE/jSXz2eLpPG9xYyUH8rAiaXHe
+LlahN1/rAk/g2LohKmkWnh5xD6hSjU55kNEgLR2KGccrBG28obLm5zmhR0VzCgJGS/0xCTd9P1H
Hz0k0uqtXmZF7BeDB+NaCMIj8OeFDNEb6X+Pm3mct0I1Jnxqx4RzPIIYOh4/jbea1G3aLKiJUzwR
gj5JUfSZ/jgj77eHDuA+LkMMi4Rpmyul+G5A+VfStVVBHL/eHEI9nIlgVfyQYn12ZVXWwl5+UHgv
jJoj3t4fxCuAyzIgkxPA0W6/OGiuo7Rnh1EqS627rkuQRUx4Qq+c4ekbU6qBwf0ztt4IpAEEiGMt
K/j1OgHX6jCj9OhbSXJ4i8PCboZGa6DVWbUH4Da15imC2UGaxvWi5/MWDIRN/7sV3qvvc+VnqKjy
k68UzKq6eLIc/Oma/O5dhT2Pt5T8NKRcIkvYvj5pT2cfcRGHjhmOwTh/VJJY2upQ9Whbbc3KNGp4
dx2xpj9iv0hHDoOq2UXnEf6RUkziF3yRjx0sr72Nl8M7BDRdl/TGoAKeGAPn6A2KrdNjUWZ61tet
czR0mVPX3rCw+J99sd6IwW50QlWn2BpOytypLdeQgilLybHjZ4X5rc3UZRhczj9jfpC5CWAC5yzy
aflaPNJAxFkeeaPvkTeZwpDxOiuu6NCN9qa9LEctsSSPaTkk+DlGYojMKH7NQgtDuBlrhpwjBs2g
eVac6u/S9nSLfvLu2IDjUxNMihB3DOWxrR2qzLQ0v8RJT6+vRYjDJl51QinXJuJROmLyzMzaPkON
eZbi9pNi1vVMShoOW9wdtdOIjBfTTYSyYMdFXt3x9MrMdzaZifPQd0YDvFi99NbsvGn7x+ZxKO8T
R+8pVXixVM63BUbdySYhmlT6AHQzxYSLRF39Bn3WT+NNkA2Lh2+Nz/NLB6dHAGzClO5NqnrXGjYj
zSqYeCIbqx8GkLEcBfNKx6xdH0Rts4qk6fCUX6a9DCeoE5IfbvQXJwCBXZTRuHQzp9s9eYR4g3uK
TmL1nnfqwzC0zk3oeE47Ga8owbz/0KFEgiOCKwxXMkHP2AiFd/0/fzPaKcxp4dAzCxhE57I4JxSb
2IIcJbZzvQNK1H36OR7g3WUDXVW30aRs7FuXS44I5s+JDdBOon2MoN1AMZQcp4Mu2ImH/EtQ0Dqj
yQCkj3mfvofabwL+ohh73DiJ6QbiTZP2uKhZoq6/Kjrukm7snBofPDUrTgYiOq/o3EYWqTiLgpRb
Lav291d9J3DRra+Lj9miNRP1Zr1HknVD240nNjoADRenLcpy/1S2NVPF/jYyJPbCJlKLbfRGSnpQ
IgXKTrbFRv6xG0JVI8ce5AkPk9jcDdnBX5D6cjNlhmhadjobOzrB4/pNrTTOW1kybUrmyiM9SN+D
k8kzR+q6cFvvyZw8+8lPQpIj/IKJpZQUJOuZ9BKgYkbIjA9oUZEiD6PKOC0cIBhudxPBNskvhM3n
o8RlJ0MBWV3N4MJWXr+EbVXbxnzvrdzd4Gppoa+xUSpU03o/2u5aeSHH6SAER5Y5lX0NCvkkt9zN
/wQLb2EIO2ti6r5bGcP/6DNYFBbe4lGKgmo6F59mNPDu1LmYF7rW+wwEVJLYAnL8oWw+DxAwqz0u
w0PfG90LViJI1b2Ga9VOo1OmISYhCkfN8fvnSATNQu/8SR7992I3a5VUFS3KF2lE52kTe+fa1yzZ
y6ByjcHOKo9aLzRpWchEQqnTNMPJm4VfUFjEz0qyHp9WqCRUjiCdPJyfeEUpB4Tk7wJX02dPTUa+
uxX14wSIK/gpDhwAQArI92CETnkdDLzvoqoe2TE9rPQKEvrT2lvoqzCNVrb4E+fyfDBQCwllPGEi
6r+71ug8qqxs4PYbk1vzuC/8TJ+YM3nXtbkxCLcr+DKC8yfBKTTcFrKFKF1fmtzOUb0htT9oDD4i
ZKwsWIfGMeBQKO//9dBqDUYguUm1tlpNodxXdHV8mfGIR6EiHj5C0oEV/hfpdNOWN4FALz+tEwDO
Go6VQ0o3dA3cz2no69sVQ5WMTMwJlzEopXRLRhoa8MdP7yav8vshwJ1CV7ehs28d7ZdYQs+WO7UF
+XoM6J3jwh+2x66xG3NO1FEUCFH3v6yny47CB3bBARk7W6VO2/bqQHb+0NVlTQ0haPNYKg5QAbo9
mU9Ous37APK7SKDde8MHo6z9CMiu6rB+O60Xn7LdmWbd8TkVl7+afD8gm5Qi9YgX73lXZudQxfDe
cMpZNyL5CINuA1qcQGa3pp4r7DltA2rD2nxpJhn7PyMt14d/4agnkdtgDn1BFyYnE+DLCy2LtbOF
lWcvKvHdgeMJqQRU9d8U1F9Lffk0QEGis9P9N0G8aNe9yXbEZZhgiPkdWX2gyZ/mTBDX5tAutkld
yKenHcooHZDIk2GHLPk8zjZvZL8/LALvEsOvwb4DnKDF82mHg/CiGWqqyy6YA2rpfOTyZvFxrtx6
m1NbAlNpyLppXPTL32SV5zDdCCfhbHmVC85fSVAxdV7+sHjr27qOsC2+6kN5uHHfveUgb42XL1o4
grFNINxj9VIwY3af178Y5LbZ+7ngwNn2+8FbpmxfeEG9sd+26DRHi3pe+JhKgO9sgz/3LNbu8AT6
sya7TTkT5UNaucQLN7l9ApFIXfKrQmp3b2lODZc7s0nkT1sA8xhCpe7bGOZgNZU0x0TOk9+P7lRM
keRCfZaPZ7M58+84sKx/4v/VucBynXv4ji6Q/X3K/QvdhsCBlZtBq4Lv+DE9KwX2pKSerYcaVQhp
Xp1tmyMX2ep8vphl4DSinZqE3kGlwpv+MlckBQVgHF6Q2pUQM8/BTSf8dLoa2uymumIUiQLxuYE7
qZ9M3ttUVr4NmwOZTa5mZNIPY2GJ4l+ICXaFTjBNTOTYonNndUYl6bqr3V3qU6FYKsDKBTAqn7Nc
y9VMbpF1xMUKTuI6ASCDi2hpYT2/P824LF0gryPMy4/saS4AGsQQZw/pv0EzB2WvXHexlUq5R9ZT
9TKaHQcMrHsVRfcGMg3YE7bjYoPAvTNzfud/hSFNZWlXA7InQU6j84jieUwREh2IZfOlgsi2ZvgV
SjukkE2+YBp2Sj0uIwWxPwFDN9150FJf8IINu59Inimn6qFrle7kt/fQZ8906SC+u7vx7vC/mVFK
EzbVNSU2d1YQVsM3RXW/zpQG1f8/a/PVFk9qhT3aHGvEFBKJD5+uyLyvqMuNf16RxhgncDr/BRHu
Diiv8t8V2IRUT9SC4IrfaoZBd6mHe/8puuwmgB9scXgrirkzdxWOu1Q7EV2l1cQKm7YxtnfOapJa
7icgzCWVlC2pVV2WJxC/txadecmMpGm8rD+M7hfXnIq+6mW4fRjgxKiDTFdQ6d5zRcDp962z1vh1
0nD1pnP7mldT2gURJdrO16S7j8wBXS9RMmGsALJfHmTnIb85B6d/b3uw+g51nolgwU/VpLOnYLoT
OtIcgyfrkZeg8aRcwlkmhpDxfY88MJFuQ4hDgPFQYUSIL5Pqsx+Gz3nCPYC60Ju3bSTaXNsp5zZo
2w+A2IjAdu4BfwpYl7U6OtyAX5Aac8rmFbFofktC04btr0TQTRxL34ass3wleRXZB5ngRjNcUzHG
P7RgV7L/N0RiuD8OWJrgL2Yf57OibdIrMw+HiPCWGnvJsxruVowTQs1M9ZbXw6vwrJZWjZmABotP
VY89TVQepcR+TcmDkCGfiIiTvoddTd+Y6rE1fWSxW/2s3/90bFHDzjI5PPRw1MO5cMn9+TZsrHlH
FP/IegGsqVsNG2CW9lXzUt/r98xXOy80WKBySe+ReavJ89JJDt3mkjY2/5ZvHIg/B+TFhNixkq9B
TFMU44RFq/hsonRyjc8W0qUldy8dfG920nQYvabQnX+fLu0XXxYUiLhjMs9TIZRkILdDoHM9yeJ3
8YsrRTmt0MQ8LXbnEtKLm15871GUolVa3syYmAcvz/7nuvp6V8BDQeMCWPfc6gRcqJHrXTYBqInp
ZRKV+y24PcO63aatlazX+SadrKN4kO272w4YYu7vINKkSJSm6isn1WXxMZ0SzuEhoWAmMkAxATA5
skTHqEgbgnwlVBl7Umxkp/RuircT950VmkKmExYwaCz4siLOYmvY+Qgvlgbiwtg/asNCbBbp9KYq
6s3k3jj0xPP/K+lvWlQyNZxj1qqTlmA8VuvIPraXZc3F8MtL5vJhvZs8N/vLbK1DaLvTahxtNxsz
K6dcq7Nf5ZoviQkRnrjV5ZrzAYc7G7Vd4M2pmi9y2Boz0X4Dg4qCySvT/+cJkc8YMZEuq2+oal6W
bY3SUQnJRI3GEfWC5t65hvFG6KL+jasgcPx+tjC7iFGK34CvEJ92/4lud/x4bsGqFeRkz/iosSFG
ZUsapSL+7myu2O7bHIAdKCd9a4Lb4Jm+dHDCDTpgM+XtFps1xlN4T99xeXFaWzTAO5KiFY4+CT3e
MfswxcXgU22hjPNtrwzrBn8WWJKeNGTEvzku07Trrjgmh1SGagrOCTQ8i5tt+zuyugJBAtKzVxoq
bFBQZ/9U5b5lB5XaCeiT1MvRYSN/ci4zThWgMi2bLqoaJiN+6d/cZyINLEWzhJx7GUb/54Gg5kEy
/X8ziZXS7wDmRp2+teuWjpCeR11aYX75xXsQ2DBIbBmFDeEjkQkBneFsuYjhPwMdQtcUIwXtDfgU
7+RuYKr9dgrC7YqZGIMXTdyr9BviUG0/PeT0yGG/Yu3qixosNpb8itfvkmEv9Orvy/tKC11UeMmJ
WeAxU6T5jmgc/ythH6/7CJqfg+8SPnaoqmnUWN6pTEJFfKlrNqjIF/5/9708w/Hzf7Pxrbrxwgid
WL5BJwdhGJUNidDowQRRTEiiVriXESn1CNoHkDGM8PEDGFy5k/IY4dyjCKwMP7dat/wgHWdkeBQI
9ZlegF+8zLNnYHOVw1tYBMo+Crj7s76zdsfMw+7f72Sd49tScVWhFiXzo7xEu5iHmD4mDgcBXfJ6
CvbSl4sSOcYG8o6Ic9TOeXxS2M/3P+JfLsnQo3WyUwdUwk5bYasmwHk9p7ZJF87zbmN8dwUuyq/a
YzF02i1V6sqzTTofzPz3V5BiCGNtoDkeQH8M0BkqLyMTEHs+pjzgyuFlKIbql4yE7CtJi5yMxxA2
RY0lgfOGwJn6MUjGZMQnJzrPgHfUECRyL1R0mPe9UsjVKoen882XS3fNWTq5e9KoapyuDCDAqwXF
sNqFgghwWxV4hX62N6RBNk01IcIMyCFKVRwnDJO1XSAJgPRFF/wpJC32SHjZZoRGYHcE+hgF3xm2
O5K1oKMNHpI54/0wAgkCv1g7e+ZJH/Nx0tpRoTEleZQLCWRsmAGyKdpAavYLX0IQz1covxeMD2wB
U2/AT2+walP1lvGKflOJ2aovCLp+7iuWqsZQwW4liGEmkqxihwJx7A9KNojnmd384MVouJwDFTYj
qzA2XRIMwq7Du3p1vyoVXLlQx3yWItU+B/ZzkLtB9zW9s7hmwCMSnt9HUrzUO03ajy2ZbXxaE+BG
izQPjLzllfvvKReuTMwlW+8D7W+1B0vWisXQawwBhvRl7O+FlvDdVY80ck9IYo9IwKjXzjOmyclu
hLzfTa/DkHJyvmHN+v72EtjFopujyBb41ajItt3lw4ezxFrZf1EBW5t4/vGOb/XVAmIiB3xPsAK2
Rmy69DfjHrzQPtm7xB3UT0mx7xk7X1zMuaH9pxzvWo5Wo78PqmnJR4PR8cjO87e0Ryg5eshpVdJ7
Uoid9pRUMoz5DNi/DipJXbl4crHoT4Xa5cb+8iSJdRdQAbsDWv9OKlyN6x8Dy2N9D54D+QfTtV2G
YfI0dK9EXYphAePxi4vy2h+4M/XZXUd3vEUtqhGi6ELyjGRn8TYX+rqqJnyx524TPRKAr+Mzqhop
Ob9CdxcqGdaDK8fDQgn3WxPYIXAoaENtTkzyPT0EuJlc9MeiLSpF2QSCMoBIwu15AUEcHPJNKLoK
fS0SqUnYbK1ydZ5TChY2+MCB20LQyYoXi98EY/hf45i48bNpIRxQl02uhogrSnlZC3w75FozxCsQ
MlqditLQXzDMMyt/SEOEZNC+Pk3MGwhKgzWRx5NAd/YPZwW7K4e0RO5T8wnIhjcXD1GZIrYqPTJX
8OHnA0j12vKZuVrRV37cl+dyakrTRSA6MLLhmA6d006bEGbqCJmeCqT+yT5TzmxvXIGP9kFJb5hO
9PH0n/LdvLHSpJJuEISfH2lBadynPgRwM5TdK30dkVpIxX2UcDUJbuQTnaRq2lHovjIRO5VfL36m
VSzXXUG52n/s2lkFlLUVz9PrZNUUkJh5bYhtu0ylBJp9CHUfah8tR6MsgMN6De2hEpffReJqxVl4
jgwXI6g/0kS/7iaaRF+CYYEUY49SRCbubJ6QXFfqcF+PHDNsR2254TUfBjf8/LDvT2MVg0S7ZFrW
q9QZssYIiGXSxhdwS/VC9t5wTIKRlWvAeFycmQGshTKYM/O5y94wEI2X+2C2pTmTc1uPK9bRipfs
ukR4bNsjFcDmVigCJqBXLfG+mKLLGgDwy9Mk1ZoPtAg8vC/mezGpMGlEuwpuDUY6NG0mWfSCpXvq
yoHrREJg7FmtbYUNKk+3DyM578+EJvVZSBpGGENhaaVCS+tejadib7EF92aCAuD3qKmckyh/FQB4
MOm9wV/VhuaWrawbYyfnZ1D5t6Dyhsl87IupyJ5l+IcpOZtFp2aDGGXqzE3eKqTMQaOqbjwZQW7E
fIoBXEGnMLdE0mfmyraolGS9sXPG6EZ40RCmneYY8gZ493QKa30nVC6pj0h8cG8ynBJ/OcIAFM8d
elNle26tt/M8ZEqLYejnhWACDBi/IkQwhqIjUjat/krnpmOYNM/9FwpoQJBO1P//IznGI25fNHwr
9UPH94fTD4xsgvAlbSczkF5TUWWrrkmWzTVdsmTSQrRAuoCgf0dq5njZ3DPHZsb/odPAxA+WwDZE
TDcGDIFknuDbLrxEAV2Y4nkvqZefm6aUB9+r5gHo351ZTHDqe5U863xtPTtjuLt6Zk8T+vbkTn7B
F1UUKsBcxtwDLv2Kua76HtHzoIWlwkB3A5k2UM3t7RUcXiTi47GDiE2WfGug/DCCx+Xhwp8cJkxl
rS5BpwVzQ02CTLzgpmsacpWfMJZ+ncN4OVzADYyYBDzwS/tdnROOCmuxw/HwAhHERi/uipKDHX1P
EJxm736PAvHudwgPbm3959AYQqXWkBqmBD/Cy+8ZiuVKxTivjFdddnu+erGtUPSgv2xog+xQDhZH
YYfaeNyHhFGkurlV6doO4mPjJNQqAht1iBHxCTfpCRW6vw1Wm/7S/TrvRrb9a5gfz7pRUcJYe5vg
X7NsRBfxu4M46K1nZ9B7IBbj4P9iHL8HwvDFfpQ65C/3eNELmZBWqiTwFOjBBa0jOnTpiwNnmlyx
kxPQueADn8qEE7URJFdZ0Zo4cpg64/BBq0egf54yM548s8x9nZZmuDlvy5z1RSbpzWOPSxgQRB6S
JcX9AeAkjED3lirXy1ZnukA8KbCZK33fQqKPN6HtEwRLFDtf/H2OZM3MT9zmokFks9W6zI/wjOev
cp4bUTGHzsU+c2T2KaMSZyxLj4vEELQOUYlFFjJMpj/bonc8D4/uGeYIYL+4WgJLqMpsl3ctMpIG
4zIhNBgMmxzUzOJLh87+leG2cl5hxD0XG1vHQYobBjN7be+2uawkEfnI9VX5zXazmRN855Ueh73o
eft3bWbIdjOTWwpv+Ue4b28lwNfxkiQPf5zQb4a4iBTWMuVzGV6ZLKC7I3KMA5wxggTSdEq4tlFW
EJzAQN60rKpykJHR2B2ZCOs21OG/4do7rtkFE7u1KijP0asnATGZyMUvzzUT49cjm7VDRrnpwCmQ
QUIo4r1vUYti3r1XyZGUuVUXYTSS1ZG2PDh1LzLpsm84JyO3dXwqN6NEXQwqcG5ie0usdZIQh4D0
54FHHUmZ0a3pm0gmuM0ZZw71yvRwpIAHkZra6uxtJdvZIpljLhG1I0eAtjkwyBm6sXjsfLc/meY+
Qp+w/yXJMdRWn4YleuMUYk8egdBGdTNKI4oUiG4acCyPTVpP57rr3lGLAj1zJTgaRxwk8XS3lL7Z
Th+CtmCBNIykf/ZOgkuJ4DqXJveJABaTZTTX7luMz7ocHx+2ZOqPYEtpQeBucqJoexgzQ+1y7qOX
ll/OAOMUyZowIp2ZPsi9af7QbRqGsbq6FAfWE9pWJTN9tbbxU1AqKZG5xJ1b9VUiyqS/i0Vn13pc
5w2awV4dwIZRelcNYybdIwIHlJTC9CBqfkIAe3mdhyfvmpzZKTd+ebTUZ4/uo4nbOZE71hvK6aZi
lhiOexlIEbyLMSzWCKZrkjC9ONSvr4N+DqSqYxE1zzyA1Kr3t720Gga3NJsU+SlKrG4CLW2mQLHv
PIM+I0go6vhgGN9EsW1MpKqh2OjJVIbmJ/k2Fw0ffK33DcmPwQkod3N26baB41i5ESbvmojSXdhe
8zJpNhEQhF175BHQy/JeaYqalLgtcrbHwMysSUZsryEywuXtemRFJ/ul7kpzaPidKqmMIBzVOln+
FDC2U2+haku37fXcYjcS+VghjTrKYjmg0Gf7vxvzBETkaqbvfBTFIYEpzoK2f6GmJDgT3EP9VLLk
d/0T8IYPma8+vvr5ThSW/ahdr9+X8zeiIecG619+xxjhwNMou03qVwJgI2WQNpALjr2BcCG35Pwv
q8sUApg6Bg/Mj9iBWOjCkApUzT98wDOKiBqAPLJCBjhtor+Gi00dCuKPRtlC00bKFEzqkYHvu8jB
57JjGt/YBp7RyiYt78B4zkaooiNrarcAUE+TctRvpDstU3nERdvMITiiM2Uq6H9snKRPtdujbhMG
2eddARFp+vlaxWxo+O43Ot6QpgkSV6nFTBa5HWbWp+SBHFO2qXaGZioiIA1CqzXwKqqs4WdAfwf1
JeLW7phbCyLnNg5EVg4V9FTJpzGRUFWHcj9QH3SICCJPrkcbUBb11hvM2mgH1l0Jsdo7AiiPj8c0
mqWEgoWnWlWEUfsxSDfR6rz//485MlgAS2lhjEHmDBxWXS44QNIEK6vl30uOyYHzfHUKy9o9KSPq
yoO+wRMaxbz/wboW/zbrsr/q4d4jKiFLdd206Xa5YR6MWPYTyOjJX2ofdkhgL90+OguPPAgoAiWR
UrmyDiBgFQECny5iMscRkr/jbnJJptG35YkKotaveTsbs5h/2atAQSAJrBIKADAyoa33mll1KJ6e
NrFWTiRcHj4CH0V/Zbo58BJWzq+sh0+1+J5SBNit7eJnlGAOen9GbnrbXUMQa4E9G6NBVqDpYbRR
Bl8jmBxCAJV2OLvX/xu2oDUhNCXSfoZ35GoKMsJv/QaD7kq/tV3tOJvkXOaoV8TxSf7MPah2NIv3
+krSWpEruEo94mwt5jqYp9HvTlQZ2bt2jdIoDytKoY477vfuw06znTkQSYQTVsudyHr20OYvWQKx
ra1ShK3J83+wC2Zv4MVI8lRymNEChv6DTCi8bhVUUV3mC74ymRrEAgNS1jhxa9lWD07RuH3mNrOO
wCB418uli779HoCWzu7Q8rE5HNsB3ZGrG20Lxl4mUQDSK/L4ywc70M6O+vbcMUMhyEiNX0stvG5/
/XRryHdVJ0q8ozB+jusgJ9OSPSCGQNHa+qKhND2moQrEKYgvLVWAcP+zuIXHwVn3Fdgmqh2MdZjL
PftHmNW6ttoIusUEE7RXRCEWp1Dk9qpBMmIJ/e0Ahc5xPURQzIfsIcu1QZBFYMmNWHNNnt1axuuP
I+BC0kC1yW8BPMHGWjvSp+i3dghQErj5nzKSbbIiUf7ELbWNHFr9xlKhfa1rNqrTdW4BFl1e2cCq
cVgVWNZxFdW9TKHfxQgn7uWw6R/aulszlvsFZujM7WLTOHGpYmq87eBCZarFyX4No9BVOPNv8nsv
GUxhxUegYV0VHKPdOQsXbSN1oc5MCKmFZQikQ8/uqu96dzyo1Pmk3lsb6dYyhC6aWFoFydD69LU8
Rl47oq6EszEQyp8KyJpIHn8TNAeI+KK7/1uWcGWpHzaf8NxcagGL+YOkfrB6iueRHN3YbdDvAaD0
ji3ZL4ffXnJnyBsHT/qJVv32mqlthlt99wpmWLyLMrzN9wh7/KAA89tvByBi+3ySWS8gYrQLlCsr
efnMz8/B11ApOSCkeJDgsx0R1yTN49iv0xVdEb5X3tFc+pRbDmCYmQ9Ho/YimWCJKpfLCq6sqWmw
iq7eiJeDrzbcu19q6MJXRD90Fouj5X4u4C96a7bmDW0gxFJ5dfkts9bwk+iCI1jXNPzZlNfgXJsH
Mqxz9XPRMNFPvmx9L4xCEMGx0oBxdzv7muq/+Fgt2FTvYaWOkXXTVd5Et2v3et/srq+U566Z+3hl
6XJgRIGkpphV+kDs3csL3NQCozod//v+rpOUKdVnPVQTR89Q6ENXdri5cxmVOvA7OXv9cP2GjL/B
2k5ssHeMNwNIktKpntKG+MsL6PFAxZJo+FORorWUwilE/S8D4T++3ccb+36Zx+BU04fFA+dhK4tG
MuF8ai7F6IVWQezLsrs00LESNZK8Qie5UETiRENQb1p5bZJoJt03HkTbngOYjSFWBTzF0sFR+5s5
IWE7aZXCj4wyaVqPzCoyTjWcQThiKp0B6uWhxN8NOoSHAWnO70hz9/4JixI/OphQJDypISE/c5uE
gEB5IAKenHEV/o9klwZhckqcZAfFlyLhtTAC5XIN1HSWVH+1DcniPlcOUugQKmriz5YjKQPl+0Qr
ylJ4Bx/5sCyq2JHK9AFzeG40I0idqbpJrYr2MiW3Se70zVwH2X9SMhH49TyOBZDHb/7G59uBp5vT
aMKARWScmBIEQ3BYW4HUfaxo5fFlDoyY02CX81RPKcziqyLUmkFcHgbEXgNneja3utAFhT+rQi72
RDJM0/y4qqzzBt2NMv3VnWgWOxtM8yMn2YHOTET8t5TocpNdOy5QCnbHkJ5Vk78nVr9jZCEpbTys
0weN7p/NtT/xLii97yR1QwOhe+9J6AYEMzzaPD6pdRxBFPVtRljOFiyVY6LAbBfSO9trMtbtXSND
jVBcBQI6ESTT1TNssGJ5keNib2iU+m+XywG7WDkyAdycSSpvy9X3T37BGKcSgnSNnzr0nlbsbTBS
5/q9oCtvVEtLXr2dLAVmJ8bQFBVhB6V8bwNwbrwkyNvU5SLiYKC/q7uYc9pocamKKNWM1U48TR0Z
DLopxkzqmlPwptfeFKUmCy+9hO7/r4Hnu+FUfsp2nBz4yteDQlkjAyTIHOW0rJj/zivIj99b8ez1
iJUt8eSsv1BxYpyxB2KiNVU415u0uO8nHs3KQjeaY4L1kULzAk+e3wm/3kGvH3sLWw105vKYASfq
mwlEEccDLiaDzEx0jBEoJ5xR8E1N9SJxsHwaIAGvQlRoIBl4fD43eZ8/HnhujmwGwjPMex4a82AZ
3yzGWdxTGrh0S32Cwk7SbB/dWqVRn/k3AgVqK0qxP5V/lgGgwnax0o3gyCa/SOsGAcKq6/L8gxuX
zW26jH+AivMjSyG5MoghKEGmlxOAvAppqyb1aY1vUFaD76IsjCPu7j3RvLZTVlAGoUGrKfNiSb2m
Hk+OJMF5SLRSwzvVYTeRGP2SVKz5dTsrsoOfxGNi+TVCff4CVSUKvvXz9Op5Lu6RAj/JxniR3ghT
GC0Z95HabzgGUYtc8sB2e83q0kUTo3bw6yZTfYHVAXBYiqOFtl51Mt/EdkKff6Ls4cGJkpfx3V/b
nYR2+CzNe9BLeSFzVBaFc0WzsWCdwhC2m17p17m2wpxKD3SOgQFbz7PYI0J2mJAameq6T3EnkW+M
eJ0Fp+ePkQYUpugfDd2B49P1CCnv9piTvwurOhuJygnIsOZMe99rRtnZgf1NtwyukC49BhxiLEvl
+e9P1pPYg3Z5e8Ob4imbFCc/bHNk3HPl78rx+KzfYRzJ6PUgdeOJZRvjXpIC1x0Fxz7X3Dfu5KTT
X5tb5oeWXwBSf2Rna+nR/cPiHujIt9c17MpN3GUWuxMEI2zGXcEDWaysxu76GBegPmBwieDU4G1Y
trydH3Om5gqZcDCXtfZWLKHAIn7LGTfrWGIy5N72SngAmqkwveMgH9cfnW3+crNhpB+2rcWer5IR
HntLOMsMjGVWTvL9z6L2ntHrC/q2ew4adSidAfHRVwp+xOD+pC4LEf232FDUmLgMqWHR/MiKDiU1
Fh9cZQAuyvEnfgGT2FkStk6QkHg1ABDoW9EKd25EEem8WNgDGTHGDIEKNzussM2oc89U2I+GHObx
1mmgTJJQGbCFyw9yXWvrFf4QW6yvgV6TTVCro/Er7v9ptvjsEL6i8+H2pHkPVJ7FdOdmh2kLkU6T
in29mJbzyKQWFCoxQJc1AZD79oZeuA1Q3ws1QLBWTG4hXpfgGObk8/0K4Cg9S+6OD1fgJzXjk8fK
hZtKs8I+9AIUm/6G6Mm0aQtR7m5iXLBp1FaUdH/Cjs6671mkl1D2fksQ9ShdBdRoQQRpkJpgVvMi
6s2seuw2y0v3EZWqkg8ziM4pZv0ibxNgecrT5heUnYNP0CEhb6ynaQ0/57O0eXsSGYekmLJJzdY2
2yBEdWLQIbtWhGXB7aiswPT88x2WwqU/R8oaKprjg7PLXB9Rg0PEQT3Grhcq3j7Op65yU08RU8JY
pY1Osrxj+qMCCRmPaFh287Cnp96dmmPMBi1m2I/x+iOfWxyPe6KofN4GzpQSMM4OIXJ0vFcAIpNR
JHNxGITrswT6CexUrAkfvZxaNwoTYgZojXJoVDEnLDPSuTvs1efabfjP+4OQVb0NluCRTah+oyaE
kCZ+JZcl7uSvFze4om26h9giigyVrik+RZRI9ChI9kBQz0k54yzECtXFEL49QpNQNmCUYkNpZauB
Ya1t+dfX/YERT0KDN/quQZ7OXs5oRfVZJYkhr6sWG7kfFUzM0kPXo1tGqZAaUuJbQkryOBCtX0g3
OBkvKztr9RuvrUhnlz1t+23NjM5yhukOdOwv0KExr11WhJfn+O9RTrUI1IvYy/gee98KC+FFRdXC
URgHvmPHJjxZA1ZrFpzrOtDX2QPjpoQCzfC1DDk47aDPLWgqoueo7ySoY1fE+qHRrA2seGL/yd8B
g0BQGnBsI/3+qH8S/3vvTP4tcfDq1oY9uuR/fnmrmROD0SMTVtYFAZ0FPk2ho8t28W3ZRfU3xrR/
D7oXglPTBwRafhjVdwNAtNnMrQ0NE5Dk6Q5szVjDhqxaF26pCUrEmwdd8aZaYptcJduOR/wnoL5r
1JEGL5z2rEmQiCjjRgUL/H08I5r1GimmLZFxDWq4z/C017DRVx90PaGbhqx5KjyMj9+mimEzxwZh
iIvMZdwXBSxFnSdA1qAvlJ9MezHdizAG7g0G4xG8ThI6xZLlVgrmYk8bETVa6bE0Qtd/OUXfWD3w
X1mLr+DJQl0lx2hSMGhupdpBJnrXXg//+bCg/9FiuICmlZqq7NioKmtEFncw0FbT38FHs72EtvJQ
Lr8ApW9GdQ2DSe6VHWcUErPTD29YqupaiyU8jZOFAynRk0b48qYuxH3B1aAZyjRv8QRtOt4zBN39
Ag4sHnzZqjZ6X60gox5Dr4XLV4/P+gAI8GKQ6EUfoBpsCRJKhAJMNsCkKFfFf7e6CqwaGHA809T4
BTbiVCp6RGL7GfQq7O90C8EZbjEwFtqDrDesNC2vopXlIyPbJzQ+gFXW9EICPSElIRoB25QE90hw
EyPXwSsyf0QmgAJ3wBfCUet2KwPrsBovUT7TUQEJC1SG/ALsATy/Lhk2L/X1KzEmWYQGYKHMulU+
P6cxk1iCryb6A2NbSnq2k1o8OTZ4qxHRU3OoZ2YFH0l3avXxo78ZyxWdcoJqi449ulxD4zaoODMW
gW9L7FImNbD1rDfX951YVTa8ca70t+Xl3uLMNiNnpE40rBzvW16tQWeV0GgpmSrO6vhCeipACMKm
l9D9yfIM0jgAxiQ8mfjnM0ba3Fbe/CCZmffyFGygJq6Vbz2ebHsk1rn+pEd02gaSOwuMiGDlZao+
QDVA0lIJiaj7dHay5YiCtUOBvcxg5R+yBG617k4MGWKFOsAVSSJFxoFz9ZWZGXYULH+6a3SMTWmf
1RPK6DM06NDy/J9RhMA0kY9fzFys8ucs4Wq1UBZf3dLAiF52qNbW1lxejsWzyI/0dtJ44TRGIGpW
uNB/3sUkfXW3L8J/ziAgqQit3qq4VuiYiFMXADNLO0VTNFNs+FaO2suxjx17o1tsTupwolTXrDtC
d0kRulg6cxPV2pjwQyVgAj2oBgZiqcZoZgBxXLspxW0j0zgfK0FTW2U8fOBJsRlksQj7or/V7oe/
rW/Jbhq250UW7pcKr2fG3Q7EsUyT0CHCmhRI4MENLZGU6NfAu2f2RirOisoayUozHMAFW2QHBM33
oJmg+Wo7BSxA65gsZdZNXHDGD4gz68kni3sVJT4Kk6NXdohf2kr7ZfbN+sgJYURGYtbbcIMA4ON7
qQxTb+Napy5mGLFLU/BcROaEhxEEreQSHHWVW1y1SeUiAZ5zagi67OMkHh3xtPRKFYRMHDjS0bmX
A8gZWPDMgPuUHg7UduPKzQvwwJUb3VJ8s5MVbK6yg3OKgSw2O1Zwg5Mhw1hOmudO3SdDfpTYYyAL
c7x5HKBeWjM4HypDZxneUUjaWm9KFRMDSn2dAfKwNB1KAklJT/LevWoMuQ1d9riUpE7MoUrB7xGC
x9EBJ96hkANqNrNBJQV7DrGkSjUjCyI4+GuldaOsXOuMnR5fkzBFtrcRROtGYM1MK8rseCh5x5XD
Qc4u5bU7H+OIgbFCvWqoKt1OPgRVQkTbuqvTrYViIRGBNx6pzMhpTqM7X9AtjIr/ZebcVYuVWiCi
JYgEP8d9LdcgZ/IYIdBQZDQySEzYD42M/bVVNLIIJtg/F6L2drnsMTEDj8fxBviQvbr6KZ83Totr
xOPzaT0QT13DBIEbi/Lok2Vzn6Wj2PxwXAN8XcaGBytOWYVz8T4fv/tGUNLOXeYDpYUEnrRDBitg
F98/McFj8NedGS0mSsDyQU37czofX6uQl7+KybcYX23iD/g7ofJxM0F2K1w/XKz8Hl1//wF/lgpB
SROmCtEjITYhxQOA0SGHpl2mHlmwiUXwdGCVTNLSWPwOdgTc0ysnb5uSHWj5EcwpCKK2KX5OX0/r
cb+cDZR8WrErKViamM153pM9xgeag4+tVpTjhNU0O1m9Qvhc4Zt7HeNnf4v2Hy/Lq1e/e8CtOCCO
s96ZN3tHC1XO/9sBuabdIHZiAuSupJMaNHVEYbpmH2Dajd/TBOu3qQQwaQY3jiRo3zFuIdvGSnHi
OcWtlD+Rw4OH6ihH2q0CyGjTFS1cqpx/zAt2AH2LPURZ8Xc0LOqCqYXplJiBxoM+OIzG2/BeJ4dM
2U/5aBIAo/GbZ+3wloXWlaQl9xcBksvUo5ZiW9C8mToLd93cweY6kAFdMMZxe+pVJom30vpN0UZ3
HP6uvl7TbdAumsXpkPjUw6uoMGqJC8wa0ZRl8N2k1OFn6ouKXHfFf7aR5I7mz4Qv//zeNblTsoAx
y/yrBss5y6KNoKZ+HRiIHzBV4x+1vZASXqU0yChyWOb3z0cX4Xqjg5RdhLAW598H6Bz7DkpeW2S4
u7n4MbDfAheVf1iOpmircOMrvZWcrFUNExwLkJN5TVzxk1jiM10Cf3sVFItyQw/dIQ5VJ1OqFt+E
mvHjX9IXmfHBoAAm391ybsmDAlvWmRNfFtAxpUNguYW2tM4iz6AIV6mcGde4RfjngU/KPANbhWK9
MT8KOZjr2nVZhNdGgTDJCNmq4qBYG93ZkRNJEWyorAUe8615+NpTpwzEZgmNEAb/8B44cYtzLkEx
9KCUvH3tGyMM+YdKa9zkbuBEzAB10PZrO/JcN1Z+H8pXkKkbbNYrjvNx1LnmwsFGmmyxXIwsScZ6
oegUSLX+avnB7+pbbVSzV0dCc0zk9ezo/mAO9BYxmqWZxKKNy/FQ/c9b7J+DfdzR5PXI3ryLQ6at
o8j+OLU5flhX1wk05vx+dubXJ11CzN9PEkPNCPm9e35og9qihJlLhoKrosxK4K7emSAGOxYeKjax
9aWY72bAvwZQX5RJ1vEd4fxR8nP/2nodYQUXrNnO0FUGwT7Rjt8WDbNnds32cd8/rTlveupz1sI4
jb21Ex/ZD+kXjxTdQmSeO+lZQkI4c0Grd+ZzauTuQX5N2zz0SKp2MmP0q0XUmQelAUtfVhRMkGAJ
Mi346A6UaRaHtA9G6SVzTyr6CMltXdxEP+Zv/LGwv8AsRsoMStEjml94GpcIdbAckhZy7AHkhVgj
NG01RZPMvhBGq0eLv4MdSrU3PrGRhDPOS1Yi/X2JBFRPZ4PLr4VM3CNE5p15TNLQWm55PKgZbgxO
UvsmxrC2lOr9wJ2G4lvfFCk7C7i63eLCKxWzuE23KIAOYn9NC2ig7y44+eDP9oyzgBxyv0UifCAW
D4Hcc5hH9wtjhPwjUpJWhS9EYpTBJ4FZWBOqiP3DMfHXZGwDgITGd4HeGFKsfVSo50mhjrfjhABc
wjBgpYYy57mT6Xp+p/l3A6GD+euVGAQoRGd8qYzN2VM0bn1XxLnVx6Eekz1ltpA99Xp9Uzl7MRB6
+P52IGVNuL1UMaODVI/G/zaElmqu6kEnQ6DnViEaMJmhy+pafetS0xikkJ4CptxjyImkGW+KMnwl
DUXIKYuKQFcxlwYZOcWus2++8lSWFQJ3hxoWZFFjIFXDWboqKoyebxKKbHmZjb46dFiykDrPXitP
XS3p8ywW0suLII6lUo3EMd+wiFQjl1s60AVqCP83PNeX+NBz3Dvyuk4nU0yJR0nWOAHJ7KcHnDq8
/g/HbUIPs09pAEgDiJll55Wem4/GOKpBvHSKMNLEyDWI4FhJ8ncXU1Y3bCHUdP/pchYF91+cVZzq
q3Rnlhy714Mg+BnMcXfJe7/8RKouatNmDMs21c70E6mDNEs1LFEmhr414gUH/GXKdrY7dSDcdACr
mYyyJZ4eJ3JedD3K6oHYuzEJZIHpbdmHklec9RLka4EQQhyl1YHMXXkhaXuHEnQOlECvn8BMX0dr
x6Toi/U7sJ7nWxHLDrT/kN+A+BYwPwu6eMRC8iHM5RSFcggg86phHGAdSdGsvK2IbUWgoEnBvfYI
z6EL3DwzIC2e6tn3pQv10LXJYMtU0baLpHZ1vg1mcHX5/y6PCJcxeIILVpButpPQznHWhQP1SQZ5
8NCBhuV8qijscEUiHuAUzPsTiznV8u0vDQL3nmJRjPgaeICB0OWSHY1bQJhq3uXlCYtLgaxCa7vo
9ojzJYuV+PP5KWGa/hnAIfRug6Yfhs5xYuQShg07u629Ll9REIYyO/CedvwRmx9fWLchBslDBdYC
xf8y2zVUyScDtiRgw5SivrhRnwEsvUO44NJ1oJnavTMcp9+VZlgx2Fhnc2D0b7m837NRtLZIZF1T
GHPN011bkJdRJuq2ro9J8obkZ4Yd3PsjjOt0Gsy/nDA0Lk3Js6bKyQe9RveptMfDSqOrgaWOIWUe
RJnCso0TpcayibMVg7/gMA5dhhqmDR/nhxh36s+gRpTUiUL5Metj4ZAzSniw9XjRsVpRVL4+W8pL
qL1hdiHgev1cjm9vFCLK48cvntwqSDVCjOcdV0GMbV+1YVwnrrhIFuqW1ST72aF/KxmTldScmZt2
1l0WviiyqTyYnB82nR/X/L8owTcsMcpV5YcU3mcCrN7gypMEQKb92buP/JSTAgyHEWT7QoXtf3Kc
ZfPx2l4UK7D0zgajgAAlmcSauc4VhYdRmvrZB2G37CnGAgrhDCwiBfUVYPcC0LXW3mgo1qYKpSJ5
xTFXMsxr6faCGJuyqeuqZr3tEg6NFMrQIQSye4lqwZCJX3Z9N6Jjw7oTdKT9IfFF8vUE/XrLGuI4
T4GN6IeVuX+lg2dmFriygDz7MWZDhJzbxFxy3DW9vBCuvpU6lYZSzeKXl2vgyVeY0wxGCClpGP6F
ebblI8vcg/r+lT33A3A/V7rA8ECHVs9e46OSFspHlI8L4cOxfV9LVxpxMY6mrJMNlacVEe8LiRcG
7eaNsfCuDhq1leYWt7qCpKrUJp1X/KVv64oatHj5LC+XjT2rudovClVSglFt5PtLDDlIap+ElX3F
hz9FqPUgQ14mzdw/kdtTw/nuWxqR7zNH/f0TAN83W972jZOkvpTb3dG9s0wVLjA8e3RCMhZkeVfc
18LXguWD7j8KSdvjbVRFWbIrOGVjXtAIzKwGO/ZBwRW2p3atKQ9cmbfv3VoQORR1Tq3PJtpokuKA
vZif4UcrmqwvZ8IywzG1T6s6vnG+mFT75hbDW3a+4Sc/JKvBGjkD+wB8/WfsRkJJJOBT5BTO+UV2
DA5xysA0Mu4ZqCUBHvAcGg+AsjIy5YKby9kujYHPq9rNdHdq0eLqJXJEvdpPuMyvfEc8Vj/Sr0A+
SVPx5XBJU8G9s0vUkI05fSSTOlVE5ntyfTmkMNUZzLYad/9IqP37rkOA93C6uRUoQgkH1jshB312
pYkOkVPeM+DOVkWq+x1xOnEk42MkLVuruWTZzGEW1sQ02XQpXQKTee59VeQ94Dtx+LsUZ+UB0iJm
I6JqAyuf6GhiccrCuISskGF/eUFs86U6na33EWcl03GGSiq6TAfxyFtA1PTWi5kd7JCpg8OF3HRQ
oc5NFPH9rmUZU9QtQR4Bysfuhy8mG31SzhxI8rknJWYKvHhabCws76KH2l1arjpSLwX+958IuXaT
3IwzcW0/k8O+wfKU3Kgv6ADt1vrG8GqlnZcnH08h+8FMbS+GcIyfdo+3Z/M2jWhUfr4N7jz0BLPW
/pS9OxxHO9XdXGvB3b3YyfJMDYDYDWEvPzzY2Aoo95pxj6w+sor9bG7LSSxtLiTPaYwuT367h0jk
GfSIOVQp3oNv7aJ7pBSJD8UdEnS0Id99hLalJPyxu+FfD9q2bJXDIhFYElNB5Lw5fjsoDO5SBrFK
lPk+igU6c7ZrqK5qIa4JD53mfdtq87a7iHpRpCw9QIP6VAdtz8VvQ1dN0+RQmGIqFfvRFoWjRdko
tRGeFj7zE9YVKfpuqbn/XNbeq/F+JMad+RTK5uyHmLyB6rmv9x77yJvGw3lun3Q4RwR5h+zflXnS
g8m6b3BMMmCJFGd363UcNq4qlu1vvmyXSPNs5qr23GVkZlpDvzbyrDTPIoydWRZ/ffcOyFBgdHnB
JPK0WaE2LtGx22CyDu9D1Sc96CY7q8+dDq3tvtDK9LP//hqX6pwzR014hayZOK/dHcRJ9hhXGS61
S6xAca8UWzM7ancai8fgMCZlaC2bAqhjkxdynQiA7eZdmvi/kcgDGIe9E/KpWUgIz68Uf4a9o2uM
euTWPZCo2abBNjV2XDdM4oO8um31pQhAsgQ2/slNwfWX3TkEaZMa2EuWhzmy96atMaZPfqHzNXUT
SlOMA0jyu5lHj8G+E8jRimk5t2VB+o7rk4aisxbQvDV7Qa45i7eSurhxNg5GRAic/cSX6DKXl8FU
iA/SdUOE+7c0SobONxLlGWqywLlzoEbIKWVBFmvcTIqpDh1uMjqLckuULU4Apkm9rRei7mVpYvSj
nOQquzBalWbzSAyboIfgzp5rfzaEjK99M5oDerTSIOfE9zTkOyoJW81CD0SHHAMTES4YPK94UprN
pqP8Yrl46Yb3aAc2/oqNzKDn7usIAj7+vRy4Vkvgex3OAVnetWZvuOgAr60byQENJu0jcY0ulgFY
r0QPbv5bcLhsX3x8YtktcbWm8Iurhoa1Pz6OZmrHQTSwyDzO3ww0ZZIWSZaoaYtZg7+24zQ+Oc7s
LNnVq/z9Ge2kkG4qPZZrJ66to7IHrYRDVtNzxm5ZQJ4eLUDyGcwG8ah98LcleGGt+n8DNzVNl5sB
Z1WqLqpKkQnxJqV7MMYbVlSqpezcTu7G0/J9YFFJoZNez98vAXIQojmIM0/OaOVE8tsMhc0r+5if
2lKOQ46s2XhgUbcqnlFOMktNWaO4VvHD6d6UgeWDkTkFSyJ47hZJeH2ioLce8bdSfTBMAfy712/9
zn38FfYgoWOF3mQtaeYGyf10F/YoT/SgPneOCNV1h+G/2kY+nXowzLUEcXsSBCswC6rm6u0NhSK2
Jv4fc7FOg+Zq0A+ekvhnUk1PgQBAhbb7BU3178GNRsO0E8T0BspLNwFQrwJPZqFp7gEB5hN5ZA2i
ZRCFScxldPlnXuHmKEfnFzlvbVuvJYmFfdV4NUbziZY31uMGbC+o2Orcy+aPFp8/GdGN0lTQq7MD
QMsCvlhS2SnUiGrAlhjUCv70TcGaLMQuCFJo1zGQqyZ92BHsvpZUszsUR3R+HpnF1uNDoq9sTdXg
UPFQzi0UR8ihQtlHmUPSFpeWzS5Uu6IpnmoyobP/M50blxNR5dN1SUVm4X/p25zOgFw8RZzbjW+O
8A/AjW9KQVSdm2Pojfm2/OGohHxQ4lukkGLAP996Ru/1ySK7NIPlFu/ixn+UCnS/rr4Sja2x5cWD
KM9N95KWRwfjHJugafX/MjtsD8AaTFI60AI5wFImycQT8Mkbkb+EBasa4AVC6cUUtHtQUHu35InT
KrZIyNR3ucZAloypWI+Bykeky7qRU29sJf3zWLPkOV5RqWvIZsyyKPKixxALDYwvqeIwrHWASNYd
W83VyFigbXs4KO+rsXnx78ijRbC4Aa6NTvJ1rTKJpwKcxvlaZSznkvFOG059bLbT8Y2iYXxdy9CZ
rtHYT9wxfSQDgM/D4yKvj/r8P+4m5rWyDEe3S2s1DHLIcuS+yrK4kcdxhKWk4HSqmDWKJjj6t8D/
KD19icDabcghS1FHm9CNxtfYiD/d1vlbibOWWGH9ZoZh4QdkbFNKEDbtVdiTp0sEEe985HxZ6QWJ
MJMX9+8BA7irF/FJhk/UPWbz8xc4whSUOQhWfaw4w+0m9kqpqtcgIhyT2rIOadwr2Pg/TokrMOE0
vovN4wwQK7uuY6uGi7lOJfy8mw33QXoFcM+bDqPTbXw8XLrK4swjNdX4SlLfOw0cuBFqS23rykzW
FmdeS4a06qtGkQDAq3oa8IGQX6i7xinyF2EfHy0QZA0KVffNyhHF3FPhhi+MWYzsu1fo/FOrBWCO
In5IpwkfFruTx+MguAI6D755GDRYZS10iHeg0hwMTmOMQWpN5/dM/WfBVGCK0wKMe75Y2dicHedC
RN1ueiZU0N7kM3EEfr0Pbf8H74QsVhHU2yrbBNj1WAVPz4qpwYAmEPHrh7oOsFvk/Ccfkc9UldwS
8IgpLpMFyytGRrRjBLCPSLMqgbQwc4c+0Q7Cn6SB/y+XTTBsv098VkpiWik2hhmo4rMIz/ejmRBO
YICDtodh32znr6/ithD1zjh0Qn38EJdRlRz8hMS+NTVqfWi/Q1jEGJ+Z80b/ouGMycXgzbNI3sKJ
LM+3f8l6PgQTqj1TzP2Mqzit9sDS68eL3vH07Pd5CI8ZLql4sroK8FfvxjcMINTn1Gg22fU8vg+9
/hFfbeGN1VczCQHd8l+HmIrqDUv97PArraFWjWvsUCC21kKsCSOfQKRG726M4MQSg3T423JWcS0T
hUgYU1L6nomvGBVlBRcs/ZAhm7FuO4I7y7VDHj0eWv/+QxdFdZ42ZrVrRP3Zlapt+30i0gYPrrxu
7hsxdtmbbgZtfz/x+I8S6lSjBNwb1xl9W3yTQIhXwHDhPDLLs8aWm4G9pszj2NJeHBBuivnJlokA
rIhjmVCwarOYL+aJczLun8w8x7xNGH5AMKSqnjKRf8ZZlROFa8SDC4V6K8GDGkKnLsREvmT4BVLd
0LqqzIe09cbLnO7mUk8RqPek0aCqfCf6yA2DwH6jSxFgSCvEcp6qYwiF8a7FuN1IialG7Eao4yEc
znX7s0Q9qicBAGi55/nAvw1GU8C75RuzINajKkofr7CmdYGsj3aeEPcxwkDBACHLqZg+hTm1kU41
5/HrjIfbJaDF9qne1wp5GJMBiRmD2mMWmwHnZlbUFy0X+MwWoE7te1yKr/lSC8TSpAqVR/v5BwnF
2xhE9FHenC6hFlnI9O0kehgxOuRug/UStLvsSJjAxcMRIrnMgAw2jER52ShaikdWZvriSrP14BiQ
PWTr54LNr2SlWbc50+7wy+nnPHrAByy7arzVhyqltw2p/A6pMxnPP+DnXA7P1JydlChrOAJUa13G
6835IjmxLeaVOI3/xFgU+YksHsO6HLYkewVKZ6P+SKJOlHnUFBn4T+KdEZDX5jzDncYIAysqPT3O
gpBGwZBgKQs0RemQnJzwgs/yP2+DrN5IFS6kYdU+ZTwTn5OXfO4jy0CEaLxXboio5KNMKMBo/Y/E
C1QgOE3u9vdRABDdftIMrlKpu6b8/Oa7+uPIuIWsIDp5sqdqAOo/H3eWQ7Ci4y5/Xd6P4owFV8Ch
BsK/XsTtC09R8JIyfrmNy1B60KSdwPZ3woiN/ZQz+RZDqYnANWlD8iSBHhzmxW280LOFP4gFe+Yl
nmRda0qRhtw3OBu/I+W2/eq9/WXvZ8FdUssao1/K9oQudi4iRL2N2oiCuMd4PhxA+b4ww2HC21Ue
z9szKGdsW/7HhdYLoT3IPlK8mfEdPuNxA5hHHvkGI/nrdU8/aoGR5OeBPXg9rmGJLVTEdUiLQZrQ
vq9OFc2c37GnVnVEJ+SQWQU+rV8rJMd6d5iCdAEOH3y0Y1awUkBaGE6EDs26AevY2RlY0p+cQxmC
QGa0VwUA4IaYjhSXi0mb74GXUKLQW9kp3NaiJ+++evb0r49+q4o3tFB+s4Im+x/DPzjA4bIEw8Pi
J7dRtsLN/nwGYkHtWhnvFYcMzVY9bBPohNB/euEvCzHaClks7Rt9R2buc3ctDx+JYcyXQOnLuqqB
Arg8aB33gdj7oHgaWtWLoHgZu+Nz+AwX/4NscZkLDVs3FKmFU6D3I/OPy+7hR9YiUfWQcIA+S1wa
MVbxykFQyDXb3fSNSfxhOSG7XbOaUMZ6ABP86acZJ7ZWxy/Bb152OTnDsyz5nJGUlXeMLKEnvX0k
znyhMg+kmoh7xnmxelIJvCTIjleiZNwncz8xoxoj4n+1l7wvjYMVC7SnV1s2RvSGDJPg2yNCKhco
Y8PDkd3lMNh2fZtgWPgi9elBkK0OYmbWNekmQLDEQCheOLrTCGtFBQ+Z5XtQ6ShZpf0O7wdwCX0K
/P0vTbVbobRJWeQ5EcUI7/L3v5w2Tqp68A3GA2AbX/x7MOzi8JceTyzFuoKXp+YpaXQ52wkC+qZF
3qAzGnblOp7A7sne4mjbUTJNs/3jwBLh574W78Nh+VfIAbMd+0W5kEKlquV8rgMNACXam0xN/XUE
5/HnBpuSrwcJfIt9CfWWKg18ybf/fdNOF16WwZi/tiu9FCT8mwENjm3Rqc9BQeN/5qjxgybmVgN8
ROn1OK2F2c1pPwPasPCVFNdnrG1RLUiIA56nqmUVKXp+iWvzKd7iVK745OBGZgvMoc/cci327AtK
OI2HtrDyZ1zIyDGQCO0OfRVLzc+34GmQlzdC1jFuSPiHcSYYCPbhpUsRmDNX/GR9VjRMQcx+YrvA
t/XxI0i521LpNnrYWedjA+xp6wD1F5QBaIVqJ/ZEuT4VtkczBedSZJYNcbI6GN3g8upZQHtPzBBt
KOYl9aDrFkFe11AmNMhzlme3/6iYEjFYPLFZUsAjps1H3bdKALbl9kSm745n4l7FFN35g0L5qNmI
dFFBYx0eansVwi6omZ/waKKXgioutmDhGbIbp/XuhcEMn///u4ayoxyOR610B3Y/jtba/ZKEz3PP
V5L6kkTGTMTfY5w8s/wt4mLRZ8OgXqxZ2iH+eD8Un7ItzNTtojhRHPnZMcBabiVUo3sQCG22xdbU
HWC5qn+7+zBUQJpfCFsNRHuBv144eZNRyqRboEOfNzPnPd0iJkz0sjNITdxOVpZULtK8i7CSrdI8
POxjee5w8/Uo6BZrjevN9Z+qdy9d/dwLOD6gJEtS0u+D4czDfXRjdyjXqDBxJqFX5nLR2CpSRKH8
o+jYhNtOvhdl56Eh1m/6klEPRxzkwkb9F+hJAshdBNtX/MXiZzDa0kE3Lvtkbe129wl0Em64Ybqm
/9QMNm9iWro2yiDUEMkButeo/uH2huXZVVbT0tVxbF94XSnr66eHtyEt9HbSM2yI0Vd3XKvLD8Wp
n5FDk0bAq9WZ+ThUxJh3hKvb8IQLq9uLB7HMDTpmH6jJTSyaXKYhNHvVOA2wLiOulOFCF2A6Bjs5
nVpKOOxzXOt89JoKwcPLSX+uWQGbaf0C8jrARjbesaXifCuMeV5gBEKwYQn5fJb0ZG2nVMUqDHDF
P5zLkwBDHzldcdIdItdZUm8gQQFk1s6nIrOPdXGWWzL9dM7GHLDXKFumOuVYb5wub9KcWWBVElRa
mKdVcEYGO0XmEQ9mzZrwpzxVwu5QajlyWRcZ35fm7vF+CwrWct2Z0u1fbRD4oEcn2uwQT9AhbhCQ
Jb/XxJTqaS0f8P/+my/NMoQ2wIR0Zf4UmKvwGmo80mksV7nw53VrG3q/FWLg2IOEO3JdOnhNKWPr
Xtbh6EdWL65reRxDGoX5YXAykBveAlDRld65moUzSB0UmgS0zmg4m8oSNA38yFyfTKkFFXShaRAx
WsbPZMspcQzdh6DsFqcZEdgv+0Dz/Ba6ky9TxjDVBr2y+24/llfSYzot8hKzGHQlLMz2ojg6FhJj
3XiEo7s9T5Kv7N5hZk1Xgiajl4H4g2Yz4C10RaLfwPd76zJrX1uGMwRO/ZrlE7ThEP6N7UotWPyZ
p6psOvNAS8lEKFOLVGo47+8h78VkOzsueC8FdA3wzeRqd8X5+qbasExBIMfEKFbyFnxcpoFKyr39
wWX0yzS+n/ZNY9YRYqVyQHnWeulyZO+NTzJp/Nzk+qRg3RlcG6443NmzGx50YvhVVwpXm9d07TJM
Yt7YusKlKun3bVBtUyWCgUZO+RJWdtorqHpvNwyM7xRUK0ZdeA/osmCccNrG7m4x9jeFcLft4+1T
4x0zghIg5MA1AvFJ6X3dKpphxHAgnRWMPFY6DwPSbEhqf/b2+0wdqm7vygYX9QIxLg/Ma33kAeSs
Suhhky3TxDbRUZyuHhmYBoO5ABh4SmXemAkACEIrK+P7/rk4Y6UmdvmcG44gBlvCJ6AI5QyO/cax
Qw+bwdTR4D4yBKx2pgUigNSM7LtRTJeaxMK/YvRotifykTIbiFTpGomTe6nAwlLwBQtti4M00Sge
Y2wlh/WuyqYvw7U8QhU4bBHM3mn/+XCKyoG1Zv8yHnhh0kgtJtyghlWDR0KxLhXZeTBGuyNJPyEv
cH3NL0YYs5/BKbbNTsSkEuIGU2BQi7ysDNcRlMikr1nVPwQrDVPRLBF9Q+9OZYEKrgZ+4mLiSIcN
soHjjWqQs3HyQo895/0D4+ZADcdx1Mn3G7abFy+q5sK9Yrl0rsIN5dNtcpOIXkSSkaIgYQwZhnUM
a5TmXddqLfSjaxy88m603s5+V3+dYJLqjtY37Pf5rK/Mt76GBlUvqZtYxujd96obTzsMnyStt9gs
6tSMEPefHYSNe/lhrxc/PpwMkwC6LWTn/BQJ1pLRftam+RNbCiSd7vGOTREnEHqAGUlDWVtG4GdK
eq8zsx9zYKnTkAW9eb5vRg6sKaeqabFZG6phpk32QFJm3Y+4NSD2raMcZEi8/oysLIPUs4b/O9wh
Nvh8pYXqvt0er1OU3NP7hL1MMMephu3XxOOorYPkmce2vC7Hdas8cK0jYCvwHV+1bgZ6nIM6sjvP
ahDNL6iPRNVeLHdOMG1E019maDYR5YWHoVstItMLbHk3i6q+r6jtpYc1dWxoFDeCFWIUzAthOu2w
PXJ4E9aPKsIrhr8oK19DI34yIu0w2GHisAevrJ/v3bP9UED+mU3D6z2omrkQmceRJGDNpoT4r15n
MbzySbxlip+NqdzEvELSBZ7fgBPQ/FcV1iviGHHD3qNWLHC08nvymJLhuAiH8NV6je0HNOPAWP4O
725LWs10bvOH5pbfzDOi0j13HPjnEu1J/mvgemdJTQE2nkSfyDY45VWs9v0sDt7k7tg/CtyykpCu
lISXK9O1oegNFnIX5p2m1vH/wPtv9+ZArDGOimMrgfvb7NzMug/cDXOYpXemXHXMxiCZsqnCuN4M
JY7Mn/EW4QCio5/N6H0b8J4DwGy0YgYDwutOiC1xVIpkHSyJ0ofADZkJlF2G+EO/kaDpaNvpTyvM
9OAyeBWkLb0oKe3mYXFLTDtJcUGtWadOWYKkWniI4dOdSFzW83f/xAahPlqereL+0wnRXwPF2nlo
yRzVFrJy4KvpZjns1KfEurGdx6di1hzssbpqHsPzXYcNEqoTIWxTF1PTWFpaGPZhBd+RTRr2bZXD
r7BJNfJdCN1pQzwZqfJ0mhDwKi7mjpVvKt3B+gn0v07MwrUOhZZCd7pT8GIXPMMAsxwFQBxDN9Qz
VeO8ovy8Ky/mksQ8OSBFVT6A29DaTvjIEzd7ojZHw/LWp5flAE1tzB4mnIw2VIMYoK985tfcSz9k
hJt7WAPol5sI3FJlONzVmBtbwVVd2PdeGqnG3sUBZFOXv4gMGZ8Pdpkm37QQv9WdXAx7/2ZpEEND
j2nudNFI02t3a7ec9MHbhAm3dJcgTvS8StVpuHONsn/1GaN1zGKPqTbQaRJKyWA/1Qc/SwQmrXO5
LJXEROX/mIPP5RH28NpwPqtn1kQ1jXBy1+R+1lxaaetXnC27HuPdsWgVV3VaWOvvivhDNzSsI0Y0
EpV88+Z3MB6PudINQJQWu+fJKJ6HjvJDknYtCbAsAikIOmGCSJk/QyWP//bQAtuJ8nrlJ3bvuFxm
yhS8RXua2Df5MxGADyn1s2N1LZzs5o5jyiM9VzaFw91qUS/jFlSzkycN0pARH5W7UJA80dK7iOPK
9rL4bmKjA8UpV5lTHsruHdZ77vHCLF7eGH04k8hLQM8Lo+hn+kuR4FxNQFsrWfATgN36BlUWjVNP
rvPG3Wf/Mo6AT7s9y4MUx5GvH33vh0U8aGgLTIkp5k3o82LhdVsaS41o+tgtZIxZfxAXDq/ayto1
3wyOu42PZ0ETarKR6l01cLZkC0TrY/YnQNbPOmsjZCd1Lne7sQvtxhiIZ0VqC2auMaQOJPY0LQla
nQE7xr+qYWZ2mMPKmi9aghMXMmqB/M/c6Z3BKiPuKpR2mOtTcV27EotCHIQDmrnMKHxP2YhCPWaH
7es/MRDasXd19oDoQNP2pfhEhG00ndcOLOP6CG94GrSlaGJcmypKHNIHxpaQ66gtWgmU4B+9lCnk
ZnvfFKn83Y6fkUI8usl5pG+JGBDpfMb+CkGiv/uZUEBlJPhcmOSmb2bRi3DwLGs3LcSYc2wrS/a8
pp9wOVmEIRcA0gQaIIX1Yv5WMU7fACQTU0Mrr+klmY+JAjhVtlu6LmxhGMZDhhBXCYes/44Q/rD8
yL0m1k9tsN+kK2u6RWOgmzEYCe4Ww9mGkEq73Oi7JHulB2xdxc8BA4qLc+/aE+ZWc4JTlB7lhp3V
MP/1YdaGxF9ALOSPwMGfwZVcdHJuberlO6sDVOJDzedm36Jkg4b92bfZ47U6QNlsFHS7Df2DDPDc
mtbNz+TGKHYG4qjGv50nakBcebAnXOXwLMt1DHZLolaiGQ16JhmcqwLniDiFVt0tzq7RS+5kFEy0
DBqjsrT6S0p2ktreZVeomH6O6bnu6h0R85WU33nk/0RVWoYnb0OyYE93na38ZOYbsAGEAeHvHL3r
DDDxv3/e4HKvpRCBX/SeFNZU6dJejsMq7vekvCCQ4MtOQAZvk/KEQ9BEHOcasM2I6zJy/HryvI8Z
yvP70D8TddCO6NdGNBGjWvm3ua0FS6CiIFtOpjpMRT9u9JSnMDaBIgRMlYQ2vgdZ3blJ+epwVgLo
AmrfqF+Z7bpCcBXZsEHVAz2ldde6s3I8vG52HU5R3rFDV8tIrUT58kSo3ryoDUP2aofDif3gplXt
2GBMujCpw8YOVKx3cCFSh2mzEiwGr4kB8YveIibzfMNdXdBDAwNzNWS/g33JfL0EPpDt8rDSLwLy
NPpVru6a1mvaaeBtD1NgCI2vCYt7YCNGuCFBYqEUIW4lzTF9xNDCRIsQd9SM4vyJOM8lZucx08eZ
zX5BVJhaUJJp5VfbSRF2PSNfdQzQ8769jtdXN6Orcs/7iqM4/KbDJ9MLdUiU7WH8venOCJCVEP4R
BbBpmJbB21rKnYxQAciToQs25gTWP+/YSFGsmmJlweHYmd6XsU2hDiEmiMqNYCRPnSlX84s+71i1
tLuKkyNnDOnvANCzl4NqUQNffc+THH2/ixyPpBf3awhZXGO9zk1DF6v+HQA/cppY7ruREJ1jzx/s
HdDJrdSwOUzjqhv/JtbXQ61ufSWhnnFfauVo1p8SmRWpsvVhZjpR1xoZ7GDO6e1lX285rB+GTCfC
2Hhp1cpwMBzPQY2Oc4azIxcxZg9C6LiF3xe3ljGTqLaA9Y6i0zChWdDFALjaA9T6i+7KLKmYMbMO
JfGXfwHFaJC0XuYS/J1W9aQi3e88nhKoVz0emFFTDgG1FsNVO5M/iFhvlpea9qF81AingZpL09Of
dsy5oHscy060nqapoEFNvB2IcgXZkBVdn5aN+7sdf5eH50XW9BJZAaKKsTGLBEgp1DStnRRQe3RZ
M9rtGmbXT8cdUKroJWC4b6ReKj+GF8uVfWQ+xqbacaorvuUKUp312JXTjmKXmfgPFK4hlp9nH1ZS
fhbwXIHqyG0whvAy2qyetqSpIyi59qZg7ZLAsZJ72pWc2lzgpkp0+MbpoFYTKymNAu6ZtLu2TmM6
MN53thxsDnzwO0m+xUUs/tNtVj34cfxkhXus51fdHreT8x8LhzaEnhlcK3tzqsNXFeAjHDXN46XN
netMCrz90CKAi5z3mVbY2h5y8Po6n1FMFOBJSM3YJ4PYAf/k9hOxu6RsqZln51W7jAObixunhuYO
I6PKo2TAnMgErjgODnjv+vd/CfiQxPcyf3G4pU2tHVeVcsJ8JK0F3RsUXKPblj7bHcsLICcxz1gs
iQyL4q1+iXYRdWIe4BspSli22UVPhNBtkMkz8xUlwHVwvSD8qXwKr6vtparfqQxMxBlVbKTCbqu5
23iFOjZw4BjaXQt5wC2uXR/58E+8sqhpHaOe/EQqP9rUtxOXM1TlN6ZnoNIUOyTIGKZbnD3JOE6f
/iQY/YgH79fCkyg1cNtZBAv4dlMMPJkUrw5hAtDGKQoDPpT77CG5GKfWuNEH3DAUMbh8DFQvSJrG
dox2eIDwSFXXO+zeQdUNuRHByIbUtP0WSVm0UD4XkNlgYjzx0+3SSSKlRAetZGUpfGslYyA0Z84n
SUkG6cl/ZhGov6jUC7oEynK6IVUxgh5/94wJKnO8+f/jTSsplf0XV5Pg+xkeDcaviwmpaD/sreJk
ac3ucfhWIEB2DTy14ahhVVIzz4sigO+sUeCxyhvbuOdLe0WWmlrw7vZqrGnDa1/WskNsw9ijiFQP
GN0tvkQKyPdC02/iaTYKEcfbyWiSC4CB7Qf/eXee+MDPMKl6Emn7NYTnp3C0RYMCtSp3brWAGfFo
IYVe31cxSa0uLBp1AvYdiWdFBYAciSi/IAUt1QIzBdXIkriy/TJr9FdkBSJ9WxyB46/35E2tIRRM
Gby4oL7FcaM4h1DTsJpy0C180MmhrN6maHP+9rzOxNHLIWe8mjl8POfCJ2p3RDi6wSkaJsZZh+dj
3GgwkCKpOa7Lcle57u1KS3tBj+1zHFIH4D+vj66LRyrxIrYC1jPaeH4HFekI+UNDIi0w1r7L2/ls
jtmDuybmZruAOH69UFdLjMe7exZKZ7JI9XQzfd5ApHe1iYnnNb3mzxvlfJUYD7rTSipZSq2uyHY3
jhSSsbADcHoIyybFzy7APcEik5JiSZ9xSzgAymhjVur5fdx5yWSaSpt8hebW+Jjq/bQrb+LT7z60
3TaN/Dilhpe0ZPCNVDfodHFCCHatCdwKEVeqE1fxxYcuAOz/AavCERMC9PpIM5g8+a/b0VDCqFrq
2H2FGqe8439JuQX1zfyGmHOywvyaYVNaB7HlQ/oRpqOTKUkDzKfE43FPAmsQdKaKs81wbKC3lxUL
S5mUMehZvB5s5U1dJDy4gzMSDzrz+Ln8lHui/77pQhKorzwGNWlLSEX5EJEHQGI2d1MFAcbFD6T3
rwEDRvk7ZlBQRSMe9eftWHu/v2cqcoM4EP9zi0wC8Kp3HlLxtntiC5cMjXKl1SR8XPqzjRHNMQBr
+12+M2iKyZyf6BSX1MMPHRcCC/A3q3mdXxv6hyUFG5/y1ktlV+y0zHI1fKK/8U5myK75nf2/j+FQ
jE0OwNtD1NEVq44suYA7uGOSiHnWC0xOpQco0qVSHhwolNM6Ysu1cpV0h4jwEx2DoNoRxcklrXud
/7UIln0cVBL5+gOEPc2t3Git5SELdWqyKBIqdtuDK4+24ZoCy12pYv5DHmFS6C+FmPp7M94Go6/F
LIkjKEdnqNAUs7IJHRTwwycC8+r8X24vtagqv6FzQdpAolPe8V0Hnp6zjgUoeaxyMun5E/Rg1MBB
RjnFmPrL6Le0AJUqeG9KJhZGONcydCEqQ/XVh2+9WuJOxtTksBAHM2QLQ4u9yYJysjUhSRex+RMV
awSURzhrKHT1ltQGHhQjquuz6YGQFaXgLphAyBTgFqrk7N3o6M4IL6GhGVKmcW3EAsOlcMmVW0B6
ku7Zec7PrPVy4CxWmzYzmgXi2AWdvcTjcDBC6lWvydLD+UEeqCMmK8+9w1ddej7hMI/0OLQsnTP4
w59F6rvavBjUztrDD7MQKk+O25qHIXk3UarP4M+/a4tR6MGLeIP7NZWaNl/9l4GKJ3b1YRWL8UNc
rMLrexPkFHodiDPWb90VSASg22CnXCFutpE+o9whV5ynZVIZQ/is15zfZMbUJWtc9ZfNHJhwJ73i
rptKq3IYv0gv3xjETT7xamJjbxpr73yOoXBxpzt6MGgbX4XELYJuhGca23MaQkBFi9Cs7aVIPCPe
k9kSnnzlBLwc/vy1h/5dpt3mYj/Gl12WbDpuQmdvgiEUFySQQLcQ++Mi1GRW5lOnHrZz9ZqVVLxN
rYj3e7d1qieaUjBJs7qRTYoSyIEItRj+AlLa0LspKDEf+MXHWuyRdjK50e0QMz6E7B7VzVzwCaiZ
EuRWZI5ZissFYYNLtBRUiE1bu5dfV+/5+AOOVY78mp4cm/RWlyp/qAyun0xF1LGDVs22Rpddm82r
+J1AdGsXPsEkZ1jPICg+wYLnqoaibhn7wnuPzokilDYh9v158mB+GvQdwQ3m7RDuN982klT51bnk
46gz+1QD1LRpSIUPMc5tHw2kihEZleeP2rQ0ZhEI0Lye3iRSPWIxnZjRGB/gDR/Xs1RRI2Jjd+5s
DgecTAHRHjJmQwyHXP74vUv3C/t4uq6ba/FdHHdv4NEpxP6eg1nEE2IJu+uuJSsKwe3ySa6NUb22
AribMxvehSM5wW0TpGK2e5rTwlhB0aU++fGiV38Xx+L65xjGpAamKSixYDx+TzBp4XviwDwobUr/
5YAmR5zeY8ad/dsbkeTX+6DDVsxLNih4EK0rgJ2HH69mbHda5Q7OlhajECnCPCkbA61gU8qL8MS7
xW010GQQOqoM8A5Sv9xCHXAJetOjzMWaXfUSsleCNUHAnL14cbd35Cud9cSxPI9rvRSpijXyAizV
2FhH4GSTKKFBU4b5EVbAI9yDNoPmEFTtlvJD29g09o87+zd3GxKaJDObxzx1fvgRfxE0UC3hJQPb
gVqO6mF5pn5QCEgdBpgtXL1tbMUaLj3cXuK9oNG+p76eQMuF5/5ChONS2VS5/lRp99ZQoP0bbDaZ
j7FSNFPBcbm1vfI66VWETHGS3mxFVfWMG+G5MhHTi8Ftn/lntOYvnvvF2hdqCQbT4zGD1/yZ0Mfl
ieLKkjtoTGtC1PP3oBqvjkDi8FTHs2uiM7MQDzWkq/l9DN0r2GEUnQa3+75oHdd+bGnRL+1k71QJ
emJRYY6IOAH+oQ32/2WfpBffGqRFHIVLRVewiKeuyFTIdaBXSo1hbdptsEFd6DJbjh9lx87io1gm
1ruDY4RwXh6mOgWuh+hchsPdjdDfGulvjuAyjS4vBo/jyhBS3I6qcv7QS+DRkqSxKFuwCezVU0pc
mblG3VOvS2Sk9HqnvBJVsioNrjX7N3pODfdYAullZhNON3StMuGhohnBRGV+J2QKFjPt7vV8GcKn
GWOhG9Yl99DurOW6AqmKPvNmVDlYmQr7cScvqLyLaFceWbfTkaJd7X/z3SFDZvk+y0luXYAAdLtu
uL5zwNOEu/noBUbblEJnNl1Etf8E++NpN0JE9AXCP1aooqL2WHGsXcwNScoB5YXr0YhHeVKLcVZn
3X/2PKDOJa20np8zmQwm3xyKXLz7OSH7LHHLZCEDe43vtmNDiaXHmW//XbU+81Vq8nKIbKvNa3Ex
SvbvgWP4YWjzIhrf6qpG74h+a44weBQKBpPhcGvntcwqDXjJM2LzUCq72sVPukNwDoC2xYT1iZrD
O3zZtuKmK3oyJgmwPFtF3/gx+sZfwAN3Q2nzF/bnGtO2XGSpxUpN4vCzK2CM4wt9Flxokv5yRHoR
ew8ubkVkSkCWPGXLk4jR4LOURcj7bimdQ8tqwY+W/YwgVs3kHIXQ+wPNGYmgduWD0yaKegCa6QiX
q4JRG130QlLUe68JQbyBOoIkV2YDcLX9rPDlCPNo3bWOHa3KpPe2cRp/MGH7wV+56SnSCMIvZNRp
38/CYy4QoNRQTUglwgK5lkG0TTYsik5Nwo1DXdVed/2dnPV0DZpkYE6Gr0NmCTBAHTWmkSErt5Dt
BV/HPV13zy4OirVqXCJU4fXh4GP2dPxe2Hz5HT3lWVPYfNOstxgRhJ5P+lgFm69phgZdWSH3/Rmc
jPIjhp5gYXULEg7WoyjZCZlx1fqhTG2E1MWLku8PuwKIskoB21BmppQkNpQt78lrF6hP9NMz7Ebf
VqHvMGds/00sJ7sJStk7hVOHvM2P+gMiXVUJ242BSYygsUxkHQbVsWd+/Rnf+tWi8cpOv7FcU4kn
maKzgsXBUtQMZ43fGe9DuRBlB5IQKxfrvzQEbOrG2do8yyxvTFNUyaCRDr86YAJwZvfCV+WhAjSI
Sb9i35ll1lO6BNwbQTjvU1D5ae7dMYhlbH8xMeGe7KZgWwKYqCZiDkxtB2woBm+WgZX6J+hFwx0S
vVYfQc4VDzvkNPQzOUvMJYnYEgKECbmL3pC1W27SEE+jvAfoqpqf5dAv5rpW/bvNvTx/jX7OuL5P
q6YXhdxxWZDKr91tNHicdc/U1gPg6ugYVIMTDT8sa75v911r5ODEWWmNMPjpkcKzIvSkFH0B9XWL
3mzywruh5AX4gIog+J5FAf8m4+hQ8MRMULmFergX7vqKrL279HBNJB94uMSk3+WtIKJcmtSWu7Gv
vNYOE5h2UoF+7n0ueC01KQUTCXumgfxz0ZBd6wNLu1d2TJSa5IHk3R7fSQq7ECITN9CDPbTgRykI
MHecw2YpRKSR9rh/TWwu6Y9FloeXr7jEfObCRGwrO5bDmqm+tRnrqG4C+TC24wcsdBAcTvo4pU4z
1JZztF+G55wDO/izBXqjNiD2AXcZ/5PtNRDdwUks6ZKw29s4kifQSc9vDfLtzn2IjRIgGM99dwPx
5WPK/iK53Pjil/r0IQAB3rS5VOR9pDexUzVWJNtfOdRpJ78xrSKG2VlSxVdpdog7qyjq/uoeCC22
0g7gyqILsut+LBXTdz/rf+zJZ2Ta7uFprcp8bKU5k773H7BPZgAoLbavUmEqvGpQrko8H7MVXJC/
ZxAWP8z8pEm2prLLqIQDVMMaNA65jc0C75AtAzgPKEj/e5UCCZAr1in3JtVQa5DyZ4L4th1XmhTD
OVQylmZ7yl8B6yg2Di3CFzL+oo2lZdwKXxmzHX5hrUXT1N4OwJbIURNccR9TSC9x0S9MIE2luPV0
hQi8YZAxBVwbcp4yiXc3rW+p63eUiTgHxrPOXAyIbalo2e3TqXTMAs/5dQ3vmlzS7d+wbTU5bMcK
tXhFUwryp8AyGh25nXK8Mc2t1x87acmfnlNOqFRu3UXf5oan1t3TZiNC29/BFcGXzh62fyG8wO3S
NDa02HV48zsPM/DucOqMokT0BrUGN/404hCZ0T9ICpQ07Eg2C8Nw70Giba6cYKr32z2VU1Odn1XV
Zzg4ngS2idmjkbisGkifxvME08YwOuntyo8HWA9XfDt2cDLRuRH4BvW44/RyTah9HpaqjNXVw+f5
TI+mDErE1FsSneEUDuKrGd3BnKyxRMePeLbls/J1T/Q1bUvEl+xwy86T0UYMUZc7KCnVcJB6HM60
NcezfxTppqKvgEDg2GJVZ5RIvsBUikNUNwDS1/OpTfF7pm1WKfifrricVKznDhW4Q5YKUV1x7Rnr
LHdVRxTiXo0cgY0qicr9SoNsCBsnmGJHXTlSqeWXZNHGXD2V42lwk81KDR154dEO+VwvKbRWXM+0
sKh0d1hkleBo9RB47VC20ehK3bjgmxe8KFuOUChbhx3mIBPcEThw3pduvuel/pkTZLdhYMfaWKkv
cVPU1U687vpX9RXjSlf8Nkbnm6QhzhsjaUNVDCGA0UIuDym3PU0wAx8B6nja6BojYbG8B3gofkmx
L1m4xJSdZa8SM1lWyc6lnEmJwHsD3eanLN0q3XSO/uw7kyMJHI+Mo7mVq1XZySS85YzsJx0mrpu2
zXdcKp/CM/sfRVkiHtPebfC/qRViVBcdGBmSw+Y3hfEUzABsfsqNrl3t2jRF+RnFppp+RiDKx+Sa
Sw/upON7wBbjV+t7o5IMijyQ0kx4OfyCEvCgf6RNB5diN8TW3s7EAc5hLvI7s7NWNoiV5TSAxI4R
oAD2kUmJ7nJvv+pSiRwchtRukZ362Fekgh1o3aOq0mi0CxWJFQ2INe/XAejvVyeIdttJmMJLVrQU
gOr7EKjuGAEqHrAaWiSa9fiAb8lPd8tdc+d+yPL20qwmAjkBU7z3L4Oynja+hYeVAn1mMLHOhKj6
WC8yb0UxFf49uDCLzPCTEtvOYjPT1UiRM1Nzv0DHFXN9vwu72luafvsHy0GKvi1WFfpiBhqKsTzV
b4HZBh293Y80Ql4gmDaH5mpL3RvDFSMK7vUGPBimWWjpVkZGaBG3cQm/7KGNk3MxOpAkz+McUV53
Eis4WerxJ9xupgeCGR85MeXapw2fYrQFUffeDbNuJTVUGUxPezbygL6zcsPMfav5GZtqb2XLp5FO
5UDIo2K9KH5w1hsL2GVz++44KhwZRTTgCkpWt7ZxbwdJggsQHgj1FO7391rnPEazvStFR8ppfw+H
GnKyqemZs5aT2hdX0j8sMcyq00b5yr1u2s1S4UOojmYu6CgZ+QH/yO9dxjhqTVh2tvXEuTjKlxkv
UiKBjqYSh2uv6a6CqJ0erihpx5E22FBTxqNr0izvnIJGajLNdC38Dbmdqgy0MpS/705FXRfhAEjP
ZQao6ZKpif0DeuDWKMVmdRsFzArmagGSHWDBPk/Lagfn7GkKqkHYiLGjYkRiDlwg9f7eLUWuICfw
R/JTMQI1jILfs+CSme0ZkMHCPsE9tuPM/HPcEfQY5HDNCDyenvjTvmnPklsIeuBLkQWF6UEahM1K
GGErf085Mbs36tCScMRfNv4ZzOQPBcfwQbACemyRvy6GhvafZGCnoBJ2qHS38xZuS0zFX3Y1IQKg
x+0SsAdtqzDr5rJnf81o4+wkSCHWzZ8I4eR0BwtpqNpQT70P97lTa9kYw2AMwrC6Ea9XSMCMrCTL
Hw9504r6tM04flLs3qciCtwZHANvxc3hG0urUhiPgUkzjspFQi9Y6yhRzQGFXfM+sYCaeY/ShNk/
EahWF4RGUIyuEr6UPY0TDR1BNFwbW54ViEqnLaxmT10hHW1SZta3H+49EesGaMYp7cZCrmT7asHT
WjtLu//gvYVaXxaPWLZZAvb+vr+yBllOOlnpKs0G+RNwXe/pNOSke/77DeGYzZ4gVhG8caHUaOis
VJoLX3hGBZIsx4AD9tzU38qrysZi+76Z/jVK+V4ZPYTypVy38NQav8YQJWAKorx5vDdRKCEfM9sG
KKAPR2HdYnjdcjLEukSAN65Y58odOohK1vtOsH2Pa87Y6s1+FUBk4H/4eVeE1OpXTmYs6ufTZnK+
P5UaagYu8CHfAtO8JeizrCs11C9Kfu2S9aDmxvLzSYi+WxxE2ZGoMY1i4I8Vj9v+GWzFFVmJVqla
sK+Bm8UGm94XCoSVAoaqhEub2daVF2SJF+oo0l78+EM8VXmoL3i+0Ioj2WS5scJlYeGpIVZ37b0X
g9TsTG9pmy9AdoOwZhzxIows3AkjPwfkShWnCobBy5F0aeg23uBv1YO+TpurknpNQCs0tbElBDvW
woRxJlGjcEPKxqgG8VZolLwgTu1RsV/i5Qc2wbsMgfDiWogL7bEQsfAB/WA9qmsA7fZJwbS87OIo
NkTyXnI50SOGsegFPQz+DSQXIDDJq/vjI1xRTNE2VoZMTnEdw/KsF59djRJh1x8N085K0Mv0wGO0
hpo6Er8irhHi1NtpAJOT5L5riBNSHoJtFlctaKnfKK44RFjRTAR/IY8G4Sq03L64kF84wNEdLQMc
oXc/GetzgZY0lnyuosh2DnaJT4KXL9Bg/BF8Sg26thilxdbmoSlbwgU/Z+o21E48LhhGPG3+QO8O
/zyG99utkMF1efl3mvK85vfg1GecomvxCqMvmrA4wpTIR8jsx7/H2JZtDWJHYK1+SCo4OxzTU5Lq
/1rcVz6PWDIyIM9GUrcp2fl4dhAAauPodOaeG2DYipaP0IzPGDTyD+LR+ZFa2rwXPjG7C4vuGxK+
BvFdUiq1NHDAKk/daPbOPbqtCfpktJUZmwlK9VKtRlec4YYsMDSDzo5kFIc7A6Cwr2cCPb/w7c3m
cvcufbKsEJ9iPZ9s27S/qhBllspmM9y/cGmuSMcTEVU71bbPEa10nJbYeQeEccYcfraoqXFQfnvY
fqOly+9pElmbPTbqJSmrxujp7uk9DbDWhtDetP7XopZuvhtR43gRQWmTBZqGYdAh4253FkKAWjg6
C2LH3S14BwUa+qtjwv41lBxMF1oxjvL4OfQhwIkIEY+HOP+eapCWnWCEJMH5jbQQyqr24ctwx9nw
HqOuCZk3qvCTNRi0etwoxDych+LL4+CeY1gkv5DikPdKD7Nn+lgwOumnaFltxwdDrf9jIN7jUaQb
dRHTznxoZUD/YxDOxN1GCwm5o5hEyqNPN0Ao+qi74rN89bQ23vXb1Lo9uB6s3/4rKaKsoqdzVrRf
/++Dh7pzJOVvslCVcJxg/GhRt46zV9RltD0101FeT868IC8/Ov7wENwKc4/xS7mFkUdvwKeQ5RRe
6B9tDTDDmd74y3+q7rowLbpz9ShOz0sH4F0qgqAvUzFZyNaO3AaPnBKSatlbOTaQlzaVKqVulFmM
8qa/1v521lgoc9q3p/VNHhxx7CDIobO51b65xbJZzfFw/vnAwPxdegG+8ERGeGec4PoUp/LHG1Vh
+/7rFM2B4EZqn35MaZfDFqXZT+IRWJHYEoRhSJKiVI2/PlDTNZ38ugu2xD0fLaY7dlRw8vhN45gD
CBwVqIZKDYLbfvUCcqjEYzNxA0b6iS9pH1J8e9stq52kiuz7i49BGLxT3Bn6R7v0kUEvYXpa/CbN
/PLyz6MWk++ShAoPstr+Uc0cEChZ8gpg8yZIFPPEsLf/whIBN1G9qjoQO0DuQNb1KfA3zTvc3gjx
N5wnnxfh7eKDETSn0Er7KKODZnncoJFeuqnniNizdXj6WWxI1WyYVYaAW1rvJCMFa0ibcSMjQxN1
BvuF5uXEa7VHr8lKbkYS6j2y8csKJ4gB36K3kfvWnTsR9lBK3uzc6PNyNV7F4xTfFSRZRPKd1Zfi
wk3Zqfqlptl9aly2ZsX+eAMGYOv0PRw4JzH0ix7gVHiqc2rumaqwIP6HaaL3Nc5yQ9qMoryJJ+5l
usMxlJitTuWHuHgQtTkrXZYGM18ODvGTVgNkQXxNMXDwmC/bwR4F3i/91pCp6LBCIgynbHiPuF6e
5z00LwshdrKltLp4Ioj8+KdvLIJtcMpMojasOBzaW/VHPJaXqRfsv25HACkpzkH8k3mV1lJDmN0z
jTwtw0+GApCsMmKx3gqzP+0trzgPEykHtmkNBDwNDtJQ81969m5D0ULQwuu+AVlRLAj615gqGz/1
+cuB4+g87fN0x6CoJGIHq9QNJ0ELktCjDNhv74lJv3Bbd20MPJRpHBptHVLRDgVA4NThCqo8Fl1F
iMdPT5cB3jQ7us0oEPQsKsnKKibthkYvoK8XnFaCHIscUSMwLzWg+9iup4nSw3mYrwdi4tK/TdVe
xI1bWhQ/4Flcl1h5z6o+2fFcvo/4sbvfpr84bFpjuAr1ddMSNL7W2HDSd0jRQ0e2fsJYa22aMF08
MeTR33ntPQ/iSh5D3bsvl4aXq47xv0wNWS4fBjMqMtQkQGlf7AVes5pmQ8VrFTIXDtcwiTRGd4J6
4cyb4Me7vzAMsYesjKjztEWpk4LxizihrTktzON8ybVbXptOtCiwHxIDxSqYuXRLxRwMW64JiSP/
ko968Gt+ID7arqRin+OAcNmaBKjdFl26QUvlgDaTClAyrN4UsOOuz7sHNTraLiiU0DyrV1OKw+My
1f1KN71DPciQ5dNLPiXXDncUtVtcTvt+TPorD6ZNgrq9fYurwwyJrwDD+a7EGiyAk2EtZeghKjnr
BkWE2dzc+N/celjHpC8xUJd48sQ3QGRND2G/oPQx6MJQ4kwcE1fIGN4OZXBWG+JR+7FGwMqlqc8f
QpY28AVcB60WST0IcNtbu4lL3La8zHpsqjKJZWODo93eO4XjhL+Gd29WBR66eUhHYzK45nt9315F
PoKGHS3E05jW5wF9ksqVXO/7W0PgA8sJGxLhZadnmGgKsAu/OJ62y2ET74B6PjeVH1PcXFbCXlC9
bcykISKPuAOrHVC9nlf46YMJ+VMYG2HKONR/qw5ja8nZ2uEa3Jc4rrUPZWksuowCSazrS2Y5Fp7d
ss0zUH1YtmmVYLmzg1JFK4QG5gjfWrMbHrY5mUjMDwFu+sdwCkFK8s7ZK5V7axnr2IhNgIc6RmIt
IWPqFmM/ERDFe//Wo7kjZj3QvcOMt14e2PgcMBhU5WEAc2174IL2fjZ0fn1VYV9UHoh2P3FNrFac
TMlHOBkhtcVy3hemMnR8Q08Da9HiaE30HmxB8mUBvTtqss1PEhTM1io2VjwWQ6+Flw+4qhZjazRt
/+Hsgi2Vm47nsu8RcBo3Fitc2Us0D4qN9l7YqcdeDrV6dJndDHPnSxzTq7PU/2SmUcTmvKP0E65v
BU/dW8dVsxDkbRLicX4btOUYZ3ThQc+gJkx8iH/NvC4FzTcBFYKg7uGDFzPpyImUKO3NV7RAp6EV
p1sUTYXnq1Oni35wKJkBlG1z2yuGeuBjBBxqZ1g50IbcANAbn+2JnAx8yidsBM+PXY5q9rVkFxwP
ObEudzUyxvxX5cnMWoMlpfiOmcYblh4ky6YvDKu2PSMdq2pnFBlGkIThzZnPuK+ghTtVv5xqfRU1
IxVN0kh0QgGpU8X9uxtpZecIVaTPAAPj+r5qh2A7KVgGECKplp+1wp714aUG/Cheu2Kzzs0K9+Un
spRwReKFI5cAoiEzwLwCfH6xuiZL1yESh79a9k68rMp8sInZmyjhDogpO0paap1ngFA4ELGxFzt6
JKZ/8BI6AmyJaQXic6jCXQvJZtkPZhzlj3TEWMN2S9JTndEye05PIMfP8fJA9v5wIK+nYHgsCULj
PWEx+pRlTL6wRCvS6fy26eqYapEkstDj8FzfJnPHlfQuyxPlOtchEPOTqEWsaaCpOQQBf/eAHFi0
q3B4QIuOqJoRs17vd7bXxgM+CcYyyd9CSBGg1+MYSZgozg4uHivHbwtOjbapynqUz/qTjnWNf15H
YOyhTAYYg8QSgXiNn5dZWna97eQgoFyCImR1IxqUHnXHiEx8jOwWJFt3f1Y0eZBwHBSfdvubLjn2
rzdultLeMzb2AXdEcXBP4X7qOfxf9QNKyUoNGOnxrGhjupxfxYFch5kFEdu/vSwi5TQJIWj9QgNN
uU6CH7C0i85QgT0c6QRX+PsnnBrNmyoMkAd8i7IX9UjlonIKSvQI2KKlKOx3af0mGNlPYNLbEbfY
Hm0MMYhn6XzBsXopQiZ1kGUuRtwzC9MlZRxWmE8pRjjuElmG4H/lKnynKiJpzgiRHn/nj2XoAL1k
vKRo0ka0fHPcPITLjaeamTPcfKKG8sW1HpvmfWxh8fvzwXHcSKxgParhIpvQW2weLz6nl5LLW7Sg
4PoBg4Kn33cpgCbTnHbvpWegMstn9NCUkmdJgHwoKRNkrFgq1VrSVu/kU8eKb7hk4oYAeGJ1GHRW
eV8gdcPS3U09KD3If+yUQ4ynC3RA06/8K+PpX/JwPwMhLQB0oKee1s/T4Lc6sTb0cYVsVbOL4TUL
kBX3T2TPVMDzveAPEfnVmUlhNoZxLALeMWFEAbvUiZ4vvbVh4nerVmuJiNZwC5/mUnlN8YIxxJUK
OTrYHUe0ElAPHfNpVr2CelF7D5w7UFbQT1WEjoSRyf4713OzGxmMWTWO3NrE6RtNkGNtqQ3DpeiG
gpOjZXDIVect/E2qe9R48/5MFPN4Vue897Q/TK69ELzBTJFJbksg6XT4Bz/dMht+yomntGBhQCUZ
MWDydIBCjm9XALhB74Wq5+NaxCuePtUsAlG6yGqsrBancOQu/dhvOBDqcEFsJPzXC7wNYGtivUVV
RRbQTwSNYihoLEnpkVr0ctTMuEJ5JWYM/9ErO43su2fXuakJdkx/Q9iALBAAUUDt8/Bh56KxMwai
5mSOIGVkg5tF1ifJ8dBAhc9I1McheaoXp/nrapFFCosqCE7lYdvEt7jgU6OtKxhOu9aQwsRo3mYB
RJhezeSdd4bMULYuSMoki1wfcJh9thuFLy9mjMTVWtwD9Vwqj9jUqBhoP+8KvBfmXWdRS1j785UO
LHQYiVCR5xA/bzFPEJZ1x47/ogc0cU9i69h8psAwAquzP4buNhbHu7fyfIPsAYDWP2qqL3anX2+d
tNQuSjoHca/m8V87PphBnNu6t4UThJH29YHuB8cEoEqa9TOqtP3YIBFBwjosIXzbjYe1P/KRMrV9
FUxAHy4eBxQsyfPL/JR4/muvl2t46rFSGYJG2lomGmzG5qtU/8jAVxyuNXlcWgmIY6wvahdTNu67
+G7QEEnj+r8d9jAhQSl/U/sv3me0baiF7ZREFA/6uJv2P/snAC4JfwOCFQz3k8TqF82ayGq2xLMb
hzO2erXR+CugbWoPivnvX5Apxv1zPCeKfXi7KPLeYbM8tvNitW1i0jkTUjEEUEaated4fCvdK12P
Ry/acSWeWdmWAdPcdp6bNhWkwOLCMwkpsZFU1dWAKiVFEZ+rrOKkgbqbf2cdzCAwWfcw6twMBI1S
hxAUT2z7qu4E8/HfTV/9specIkeVcoLAwY88la9/ykvZ2oRvYbNrDNqXGfnd/Wrnk42KGwVBo+BI
BJFQVfuTPElrOy1nSRJdjC83Bmrdo/n9EW72UwqepE/OxSYvXmKNnrO5l01A40flzGrDPY9vwpRc
GjZd4NAniahPQofpgQ31ibJaJdl+w3RqBjuck4gWf7ptfwvfFw9A/jH6NHqsptAGQthxPq8+rvae
Ktofot6+VWgcCsSYjHSsSq8hZsilQRo1QonoZE/YbyU7F5fNlpKn7udEGyh2TLOtOV0I17yFh/5o
3J2lXl+Xf4Bfco6VPw0pwE3fO2bccQDaOMeqg5kC+v2VgOA/AhVyPtLVEoarHhQ9y05PGL4CQMkW
6nE/D5Y8TnZj0XrHhu4lcN5TLBzLRwgGN1jUlplBEOtJE4U9T5IJkrrk0aGY4CRgdihvDskQYnr1
39uqn34hcLadz5mOgqpf6PfIroiEkcNeYGJnKOts6aXOLVQf+ayNHE45H3zCSzdx+9lAIpMar9CE
PC1ueBaqQBtzUgMOZEPqyFFAnnt4HdqPrCWehoOwVpnX8JMOAd4AcJFn+wzFM8sB7H+0hhNVgSuK
T6W0t/KjMi74g8F7UbTDzZryNBzp2m6m8gCrevg6aiiA2gu9/BSTeU9C/BDfd9fiyavXREw5IlOm
1D4DX/OTuLTHzNc+iZMDN7nQ6EroXgksiyaGQpT8Pxj3Y3zZXBlVNyav5ca/nKyrRk9kPVNJf9s9
9F1ftkmYUVRuPEEAGYSZGFAec0CfSlMMZyo6fzOqizC8zYcXwzpTSbroD9WJEZpX/Ll6wyVHKK/h
2FD9mxy9+/I2stldEVG0pUFnFHJciw5UFe4jcTsMSL/33XSsEc76MlcqNju3QTBEEhFgVsIZw4sb
aYme7gHDDiaiFz/BAunHu3igpY1hQ1rqamg3uVOT78OcgzkVwz+eoyt6itp+XPdnxgV9JvcGLsX2
y1v9+IOMqdKA/Q+3+InHe+9jfl3rBQA4NA7m0z9ep/baz/TrcatS5kYJX111n94OU7yV/9o+wS4i
mSidX2kOCRHWt/Lcy3AZ0mWhpuU2/8flG7DyI68W3uhxcEEhohptBt3JI1Ct7gctJhN8wls3S0e3
1zj1moYr+e3/3S1pNbuAkAaDjpQULVn92Ogvoq7cPRNeMbzQt72UPCb3jrYJ/nA4Wa618rZfQUG/
kVCVpSWZzUmCWxbvQ7WXy3o3UW9iGWSlVH5Fo8NIcU+UFgsmHUfZPQ5DIgFoGd/3HMTmpgKlQjoF
JdSCn1UZFo3bRakNQ3gQje29LagcfaxjxMVhGs6qIGf/rCtUi0faVlcXvEr5RL4rEOgOj7PCD1yB
6rVfktnAZEKjABnEFC2n+S6BDjoozJP/Gvxl3EC5Sp+S8T4fCWbVjn6XLQvNcLJ6bH/9nJo7r+Cp
Lh79tQnceBWaAi/tEo8Xebi4v5wZ6lbHFFMet/csIPFCaAYGwDVkzQpbpaa4UzD4rLdfTPmKtXgL
ddm74pZyASaSYCbP+0t7ZpwDrqxjFXJAZIPygu3YLRwuXs1N22VFmOZwkP/7i6WuJAQgmaq6/CRQ
OgjxClYwsGRY4uRKfex0GuFV4eeHH0cxL8oqOST1wRNfsLMJbTCj3eFJpTK5QZm3pKhNK2mZ9JmW
wPI2apGXytgpYP9+eWCxbgQljjILIvaZ25Slye+vkK3O4D2kymq1L3UbaoBT92/EXQWx9WVTDzo6
EtTIMG53LZ310OavhFWbfZh6HKfH4lgMyJgYZ3wTD0k5CxjS8pS2RsBu0n5tDgrSQbsnjE1d5llh
vIKpOTnezboir2eD5bzt4Bq6r4ko+ilQrvqQUniGv77fqTrZS+0zspovZqOE1t6dql5uFW9QeRyg
sCdwi3okUUGz3wQUc5bIPvqwGVxl6zFZ3Hg/asMbSzWJhcJ2YuYjOnhxKcZQB9Vhvw1mrhJM7laf
4V1k1X6MtvTFXApMqQC8E2aOUQnoI+pXE+rkfy1XzmTnWP50otJ3oBNDAiNbNJ/AA6rVohG0Hycf
2kLadiI24+JD1xqjL0Jw+eK0wv9ajk6JKBUFPs+AIlPSHNbHIxgE+GfqxP14uvSfUv588VI/w09C
uVFj5h01p6MsMkylCLtPuXzJfjPCmbQbWv9eF2/MRDTTHguGrCVxCgxdfdXnEvmmvNezI7MLPQ/6
MCN1iaqZJsfsd0O18ePHouSmdvXAbEZfuDhMtSXaUvx1sXmUvpJnQZ7HSMgqHrBWZXE6yULFLgoq
jtLazouQwJdNxEvatsYSzpry/Cga3AAMJyW98x/91M1DsKxoDrNDoB7892gQOCojfHE6fuKG1u7A
KqYsfMcUdd8lWs5eanoyV65K6Xhnmr+I4CTbEoPTTmTzXwnS219PrsJ9wa9uQa52AJPjmCOSHj2I
pUvLL7ScEKN8iXg/CzoGxk5OyoHZgCuaD4B0i7sh//tH+zGFqkJegjwPreCJkMQ+DpPP7XG4VCRH
In2OBKJp2lbRPcT4iTTHcWd4v/ceLnE2/V14ujkRuVeBZHTWVKTTwb1jnGB2BcrXpbROXiDsHN7O
izC/jnSA4YAGRN57upuQdisD6wD6hF8MNX6ELSA8nQhxbPeGP0e44qZvo0YIuh9YWT+h5e0X55+h
tUYXnaOnIIg/LDDqFebUmBGYHbKOjN6tcrZjNV5T0eeuGC/U5A+bamzAM3ZxTZtG4wUINfTtKtM3
XLI9Q5hJC1KohCdsani+uUB5GFJWxk2SofuW5JdkjljMF6IUYzdYG8zEv/TGAT6XwTjDvYkObK3K
j3WIvA/G0FXRjAqIZecPogTJRAmxwClattB5BFWCbKlhcS/HEaVdFvIoUJ6RsoU1PlNdQg36xcoN
f6G/vl3SDGc6I7G+Oyzjy12Ma8jtGWStA1IktmdL54bzxZMGdXJzmecKIDCY4HIeT8c5ZDAzfGb5
P+0Ke8g2YqUyBjXXHhekj6zKDBnOf8jWiKAwSObVjaiL8OcuJNZj1AKwBBnzkdyuOYSntnCM7Oux
VO/8aB86bXvvq/mZbXvv15cbIQZKY7tJzwgJNm599/ILZLXiBgjMUDqivbdI5YHMisFTJtzda7I4
v9iTe4/k0m7e5u+oZa4uU8xx2h3KUhaqrOWEHmRznbeA8M7s8PiOJiEzt/0+jhslsim9iRYjv3Be
3xa4FQYNlGgy2UtL7ySZ5Jz7CeUV+IBTum7Cw8uIQt8oc8Wu/pFvyUCE+BA8xRHsF+QWBDHjUxl4
ndroRg7sOcGU88av1KsFpa1zTYuXGg2+hSN1/n8AAwrR5T8gpVGb7UI5F0rIc9Ptcp3ulaYzI/JH
bhHi4m7kFBkYfp2j9S1nubaVlaJjNpcWq83HbmcpwNZcuwdGPQsia7/HzaVHE0WR9CYXCkzgicRx
GCfPypQvzGMNxy1pUaAsgOGPlh+Fk9Cz02cJzFWCz6hjb1LscC9JLfV2//1dwCRhLscmi0BENpU1
M8kHe+Vh0bZloy4gjF5nARj7s9kG3EtYlXqoJ5+h5dAFHhj/t/OAf2ujaAokRo0QZKPKsEhGWddC
TcmSbsvzB9ewq13oGpkhsfWTwLQnTL7/P/czwP42RibbPnnRtkI2wC6vDqY+IG/t9uqvrERE0jMw
Qd1AUjYA3E00+Cn7VY4YvTuel04iX68gxHAsdZtbbpAIVqbVvlwVCAezP3FD7xdSgfc0lSkiPuPE
qDNDNabM+S6h9uAtABgOGj+c6FsESfwKSDfueBFY4tJi1zfnXKQF5lLDiEyv9tdt9AptVXxIW/z0
q39PLHFx8FunwH/mzRZHM+54VzbuZ7AfDDWlAT35xHckiN4in96dn7yn6kQ1hFPJhT6xNJdJv/NM
94+8Btmi9DIxe8gBu1guoyEOz3bhQUpn/PmBSHnSxO12J410VDrVff4EFHI3nIcaVvzb1y311Mi0
AIqExPZY4kH4hkWQNKyZA0knqpfd2lZpKL1eyqGWsKGXC+BpGnz88CSk3Nh/b3Tu1ANYjkQToBcf
2OqEydRwvQ/fLr4pYkyQ3l0CL4GUH38Hlk3/3TTHBvjnc39bEUi1Hof9pX4eE9dUH8p1JKcNbKaM
v3BoEyI36ypBvdorWMuaxfzZA2DQeE4/FR+cZxxiwK9kUcaFUAyRa1zv8cSkzgBX67iMbJUyEhxI
Yxh4Jm2UeiZNMeKD/J3kxeFY37WfTb1h0Lw51wj4kU2+O1uxPrCovfU3eGrJFYEhw2Q0CFLkngw+
PGbJcp29D2Mm9P3/V9PrbSvXQy50AsVAUikvlOVUl5nYtQsPVsgE5YOktXywpcJ7Xfi6kmbddm7z
53q3CVnqK1/2/P2r/XytD9HrWxjsQ8VgFnB2K54cp8q5w9CtXmJ5UTZ/dVytZKb2HsdvHRk11lqx
7c3x5m37mXoGfNtXBo2lV77LJ9GhwGbCApn7QQZJSv0GwGjga5jULgKOuaVedRHPrZ6StI6ESEpT
d/8ndCnmx+JbOwVgtP+qNyepQL4GE5CSakgTSbW75c027rJap2Q5UVLvKTDm809dGlirOTL5C/9k
Z2CuQ/VQ8+FTAGzWmIws9ofqiAeykNbLVZq8G0hzSNFnO36YigmqxqWxMv5b//1sWGXnkJJ32gRa
K0OsQt98mhqnwsSw1MiNmgCclsnnClerKiN1BuEIpFBS/6o2v/3518aYyc9TGdaEBE4XunzbE8f5
+KcqI5CttQyVNcyd6Uq4gcTSs1t5Q8Y2GOkABsmtEZ5/0ZzXYdLcqlRFqIRiUHR/cze4WrwBIGJ+
r+mdU7j8IBVWroCVfOvsX2a2Q7AVIMTviDyiityiwxadTP8fXakIgoUPxyNdKcX9/8wlfhyLrrSh
dANtXMnLwt9zZtEQBDnXf0EGKztMCeJQAFHXzQPzgno0aE2pzDRL6gm8eMG5FkaFSQ2E4R4YJZpD
IUTW97j+h+745m8mbbARgpYUrOYH8ZbDrnAs+V+eVAx/y2IF4u+A/6loENq2yA2vtXcpTv+jQQYa
8pHCssPZV0ahtWP6lrNPUS7LlJL64aaNXIE2DmENFYgScObwpNgnF92tT0xHWlEXrReg8jb58jcA
HSBiwR6F8YKFyU+iJICfuxhJb99+zWr/ZjHwU8QSSrBaJVueKRcnDSqRQCXGS01jnIB47MueDsHw
+C2lVzYzB7jJuSrgCOq09BkiF0OysYyx28Ew4CvWtdhJ+n6IgYljUbhpJcVROwf5mGu8crrhHwqp
g+jkr4/mpOcjfzV5kLKbFkvAJO8fDq4EnB/sub6AVzBBiO1Tor4vEQyThas5ih3O8QbLRccRF7ke
KjvniI0RK8SoORASh47twXY8DwcHzydSm/2g/LkpZmPkQKkr/KX4UgvzBJvtDYJK/dQCA91zTZ/0
WvbHGDmSpOVo7z83ljVxTgogkpHHPTbXV0artnblvxFgutU6lwcN85MRFY27kEVj7MeXtOjP7EyP
HoCoXQPkVoWAfn5QyXaaNxH51uhncu7KqjGOvDErZ+3FmnBe6xH7L8v4Z2/SAN4zNZdnGdb+guvK
2U5FQTkAdRXnBPzVhFsYURM0cQdA0ESbT5qLTMzxdJeGR0h0DuUVQ03w4YAELoYaidoNycpHSZZw
VzDWCZhFEXhQOSa7Y2qtgxjbs/73bQXBd3bFa0FS6aVmqygeZBUq/jUtNDhHRbwDbCVhIyI8T3aU
r6TTz6cvzUSjN4QBTCwOWwyEqnQM76btXdExCtLEi53R5Q+pojN0lyZLyJOcX8mfbCM3vWS8/iSb
1V+CifYz3m9Y8vd2IrSdqEbYXgqag3ONliV1/1GBFI5iZQ6KOWqpMIj58zPWQN1jxIJ4q6PfmGBO
B8t/f33CrRHR9DjpEIYsvlzghpTZubpXGkgou2DjQRzq9KYfcA6gcAM3j/xA62fNNhi/tOHdHUUl
SF4rDWJ6HGLrf7S6AC3U4KEFe7pGw14WeFB5YRowLaX6VAoSSk5SCrCBp4m4hZqBtsc/4cI4055M
dXsYqjknrU4RhtpgAVG79s0unJyTg+Tr6F27JJu6uuBAPFR2Ba3ZjckATqgORHW/wlBU1vkSfs6k
jhr6AFmiIXoZPfr1Fh7WpVb0BEXR2e1Sc3uEzhqonk+bTuSUKGZQ+C0V2B34QF/OSidQyJo81EJ0
TbNP++193V0EWbmByFvueifJVrfXlImWkyppgA1CKrX58FmwHUm/7szCBvc3SXEqcje708tqXxm2
tn5nS069174rCncRH/1I3qSn9v+1uv4AtrbY7w+bzBbzHe3A+w6j6Jh8FZ6y70uaIaoesv5jZRtH
i1jselgQiJtNYhj/FZs/Pp6x5gdRfZRy2XcDxICoFlJsX7xvnMt7oA4QkVpC6YrcCedH8thCit0A
rEpv0Cu8ejh9DZJwcn4mf2yyvNmNBGsSDDMiG7ABUK00IGUjIlOFEK2Q7O7fei58GzIrPX592TMo
itOfla15V9YP/ybHZQgFL7E2EGMlfIl8ctO97ArZ/TJrDTZ97D/5eJYYam80bbLsFGrLqYN6Zx2h
yKZ36bTESqxMrkkB9lkjG2EXLFutJMKPTIn0Zw3osVwHR5Rvag0SL9nd1LHJETtXuNIIW5Ua0j6u
XWeKj+RuTcVJCHh1zc7VG6NI09lqHv76a0zTOAKlKIrIMnxwdf9Rb6PH+QBbpI/Pg2EXGJsIvf1w
OP+jK3Khpg9YJTmsKGBRRmbrKRLhrrayHuC26WegySjykFqx8iR0v2Azcp1L0BMdx0tvfoOmYHBq
80IJ4P3o/ioyqIPPq40ygcA1qU3Ti/yMcKo8B0fwfZ4/FhguA37Ppw0WiOGhvFjRchsVEUEVbXml
Uyuac13j5m3HakJaZRPOO+1jCtVZWpJmXpy2gTjOLQxsDu8odT0uusJ7lpc9MjSObUiy60h9r0b3
zbqgllM23BVrIGNd7zMxp7LvGWFCmg8L2w4+2jSTSAhoqzH035ZxhLuR8XGmpXQwWcGBhD2fOk4h
gB5GJ2AS+K+oeudaFoXu7eZIN4G75888QTso2WmWRXTU5tIGmWlQj2A1smNzqIcVgld1xtAcjFQY
FHl8ezmniwpz6zOLxAKe/gxyHjtJksyG6eUfOoJzGPpwDYTUykkgIHLVs2IxLny8mLgmSQJfoguM
6lBJX3ogxc6yMgEebxZJqDWaDfBllD9YGadiC0NIVG7VRAF5oBTOhx0eig6VOZf+R9e+TDtAHfAJ
9B86u9TYDANIaWyXbyQxQ8g9bUEs9HPpE57Zoh6Wfh7fepqlQI/VFFylB38l6sPF9dEdJywMRJwI
qteyx36JLhIiJNkerktpEK1SPZKQzOfXFZcH03EjCi+rpYSBXwdMo6qqjhuQO5u4YxfsvSRLybQ9
dXSmClcrgi23kKYiZSPeZMwOftxaKTzpWNHUWt8iDRS9bhZPV0uMQCpBPtCFPlpshy5wtD+B4uMW
Hzsg8vyj2c3Vtf+cEXaXreuVjMolwa3ANseftmDS0cHv330vLoswJB8Sl3WZabtAoiu9WwbmLKGo
yo1R0NupjLdBFBiVpI8H8bbbpK2IvKHTEg86JaSh9gmOajgltnTyzaHnpLV/IQAyMeiUfQypeN64
Nx0nxtPW4rKu44OGHu5RRJxxl17B+Nqi2tiAptKbskjhCdU1KRLXXCj/LRx9A7KZr+gs93chLBbd
pC6UXGm/GEbgqyNb4qOeiWCkMkY6Cn+JTLYewlsJpxPOBbonDTqbQ/GX9XUp251xDpAvazUIyG7c
t4kfSL1fjdCQhkoNKLESRl9wxBa/YW+VCr0y4snxryaYUrcvn3AawB5InRzI3YziwWDgmE3hCWyY
kfs4Hfe2iyaWhn+NtjW0F4aJgHvRSfCeKnNDPtdlKxrBeqKTLLZgz8YBNXD2Owy6et/byQXf2jrE
J8MG2pMR1UXcmAW5tJqgkl53qAp53IsdVBIBLp0bybBIdNdrTklptSqYQOPCxO/Mc+vpeYLJUC/k
0EIDHBzG3rpDxIbDNxbUmqUWxh8F76wyf88R76P8Ue0DM7YxytnaypdsqShqLTvxIywEO9kHG+uE
qUXldd9Kt4zH2N+DYulFO/MeLSthbhjnPx0X0xze/ggo6UNUjs/3Ri1IFzi5WwwUPuN1SZPlsnw5
OA3tEknlwHUtoDIfvwZ0i0sK5MKTny+lLn24hjmRtCoiIlIfRu/i58sXeN/QRvsiDjWqMs4QLXAo
AXY2hmZUq77OSgYA/EVbWLzKWTKhUpZrTOxaWit6HeJK00bTOl7V2EIJ3HAV2dG28csxg91STfHW
v47Y/XUI/9k9daEPCLFGIUXhfBo0daaP+7rju6cHeTTYcPHGlWCvjIYsFjrgzPrms12Gc/pI3edF
mh/41QaLJZ3QKBDHAexZ3zX47Psq0z2D76yfGMYQ1Qhe9gGAAjILlAciAXGM+1ADnOEYSd6rOUho
A041CpoHL//qZF4Ll1/56qzIgzA/oGAahXfk1wG3xg/SPPzbtgB8iYQDT/pXCS2HyZHsPiY9DUjW
Eg5C8smFyStF4GCGtqq1VU9AiQtNbKLsUHE7Rv1aY7x5UzXtlpX25pKjsCarMGmDcU59UMIiYlLH
JKJ8BFJ7hA5bMsVYtWb1vvc+x8XAky6e/9xHsGSbxdcecaAlC03aS99G7yW7FsAxBsvBQzKejKPD
eeNWVc5uqIp2r0mChRrh6MPC3s5vhp/ysiW4ejo2fFxxJQSLc5g8QF+l1zI9axFoHypbTDjZvTRt
ASnaAjJfrCZtSMm4I6ZpXDPJEZbWu3Wp2gcMoukR/p7NsKT9onEwkvCd7nCormGgIAQaiZQm1TE5
9u8QPMgcCewieJIkf31z+Ptooa+Ir8GfRAYMuwW4Gvmj4QuQSHIkXCZ7OnRcBRWL812vzwlKQfR7
p093t6aYJAX5bmgEHkW7WxbF+y1qCBsgYIwfOfWcPiuD65a4j+ZuLNvFmbnhj1HOU1hYgxEZuMeJ
0i+dzXuQN6o5vYxjU1Zn12CmEkzMGpxYCWqXAOJs+GwDaBFMW72ka/BejrtZr0K5a4N9zCwruhnZ
UnqptWi7SuBuxFmgbAUyhPXYKUtcXAJL15RYQyuo4L6bokMfHwUF0iYBx/tCr1jjqHc6E8JCwTrk
4ObhNETNc98KAEORrypos+LCXBxQ2Gy1HbqKJhdYmCRCUh4Ce7Qg9gl6C/EDqIcwuwzqp4OELaUR
8zfCwRPY9YtInv0tweq2wJeqzxlprA6DKMuz3hcLzrl+PJKX3Zcl2sdSR0Tcd646MASVWrSgsoDj
fxEd0m5C4pSL3l/NpRTR31BQCJb8oNgDElCg/yE3qj7jEFLX3UD7RIs4yyUtf3qyCxjH9jujLMdx
jb1Rv//P2llrNtTE859YzQhn0fnGRAaB2AXs4+t9pOxEGO2164cb2G3CY317JX4uZ4dR+oYEvOig
pMR3i7s71LfhfxUtqEaR9orCy9qDoqSs2YO/x5ig6zC+Vk0hCcI3BAVLP+9I+HDlTPx+vLxhTHPW
f/tcrJX7OtiRIQM0gR5on0UqkbYCBZYKFIlFPluN97SJhJDSrnD1lor55YJ0kswgt5ZxgZTNSz89
EYlWX60TkhpWQGIXGzAQ5iPFszM3gtb1cEseSB1b/BQBr3pMlKc3NZ8tDymJ9LGMkhyYXlG+4B97
ziP8PTM6ckIuCEh+njtX5ZCBQZS9UhcelqyYkZ/OEEYGxS8uFih2MMRHCFIqx+idoixT6gMC8D6h
IJTeVkKN52Osw17HkCoXywNdxnI0vEHPsrH2cAUpToZQ1CTQgrCd8vKtZp1iYiPxnAAYVxc3dwdv
XsjqdvKT0U/Q5TbxnvEZO1J+18oGz8AMpg4kln5A7OqhinJEYC1i0vpKmOyZ1u7Fwhmpw9MbhdP4
3YZ0k7eyxZPIfRUAeaKBQnvO4fG5mMvwOpQsBoq4iW54li9xWGL+O+7zAEu8A5Lx03JMc4pOObBV
nva3evrnqN4FQGEuJRdJ+K6RrejbK8GfLA2niiPfvZpcXGdkaFKVy7DVRH7/+fgKDW5ucw3f944N
7QumR7TwkNIfQdthCxbqgpwcbn/o7NMIEPrisjibh9CxiUu+L4ktGLXfnSXLCunps+wFpXM9BnX5
jYXi49GsMwLEGm/Cj4M3NNu4l2+RxMzyA0ljryPrJN35NS/aY5kUV6mXJIfQZtBcIqjdNmAzlqiT
ByWli2qQWJFabtckRR3iqqdgDnGakDsD25GPfIXCO2gZsTQjXl34IuUMekIRzP8Oa0AweE5GJwo0
VulfxweXVsrPDq0A6yLPfbqU36OBx21MJNHsQmsy2RzwgckWLgvS47/rDeRuYxYCqRJiS2X87LHk
ry5xWvb2VXzH2wHO0rDKHeqK2jlb1FRgKPTwY67lsqIf3Fn6yc+vn3SnG8uYh4p81cbF8GDT21qv
pgkJtFd/DGDq2h+hfqaZZalpUQQsTSHS3tMobAiTnahNlCFiXF6NUzdSkkADv2v1VEadhA+ea9Ie
U67eLgLFuN2Thic2Vz9gx78ecfYmJfvSU3XiPqInjcG1WxkBpIINp/OH6T12M8X1lPL7xO3WaA/D
LqvsqBxPTifZ65ncGV0MlLWfUasDhh1EyAj8Mi+/OlAhObnDebsCfPEhUPfFOIvSxpOvoAYPdNRI
kAUjjKzfxx8CHTcLjCF3/A1la2XYxfm6/BBgTMtXI9BBn8IyoDnKAmb8WxkUAfmVtVp0A+QdgmEs
SMFSTPoixObtbcX+rIz76KI8KYL6iPMzrCU0cTK+xqVArPliaXTtUXvRoNhK0Xz+VIOImD8CViWC
6gaDxXFPnvVmu5UpFUCMGl8F08L44j429w8y0u71Z2hPsrWULqIZV+b7VD5r3W0bys74eTi7o+cX
zP07r6kyFPmnp9HEcoWIV3JppzkVEAHs82REcvvjjqyiJ9RJMWb/sKVI+Zfm6Vde3enM4IbmP9fJ
fVgh/MKzowdEKS4cTSlUzhj1aXLpC4my5SMOIvvn+0HszrPT9fL3C7B8cQTbo8CotOl/WSwpJeY1
+OTy+di3NN/sqm5XhMDqAWTfweg2BMF3IqwTGkn/31jgB5vZJXKM2EzO6c6pC2A0xrFe30b01CbB
/QgBJwYM/RTFt+kqqg/j5jcsMjh78sJSob20MdnLrtYTgtSwKMRFOwx0ET5dGjOfnrnocEZra5th
e/FSQqVHFOA579yCzBjNU/TpqAEEAmLB6Jq0Sdgra//D+oX/XVSBqXBZ4XIqpZVz2vWZvYDNC/gh
r0oOI51JxllWhpSLEP3unLRHBZ710GcazUmlXeVGWXk//31SJNzc58pKLfA3yMoFqnwf13tP/Qoy
uOOm/NeubgHXobIq9ULcNBeAY3N5aEOMtLzSzQZEaFgduH8juiop3XAzitWQPmBjE4e5SjcbrV+i
3K2xVP0v5+TaqoStinMo+yfr1pWZ8Bnw+Lwa7xSxq+AfccGShOUrN13tmnFMD2gr9Fss7R7jOzlA
CkQjg1ZJEit0VgLfvYVEUWchlF5gmukqd9duJbxqw4dWAAVwlBGr15Xet85Hq32mejo/dlJ5IJAh
3e2C09iGgy6oFPj662EIv0WqB1/Tz9Mf0krAYgR6j207Jy3UMKDQPwh6pKjHJCwDCNZ1bb10u2RW
Ef2B1kznRVWv1WSd8+uJ2WD+HvmcNT8k4Tn2+UsQllAJQUWp3dzrYXNMt4MnU2mF4zq6xfX2C3sJ
7Q+PY3hUvO91Nu473/p9zbva148jttPlH9MeLcEbCmzikAl8trWA7jlowHhkLGqs7N3s7ySu9yM1
aDyCoCHpip5lF3wRKJOdBji+sFAQ9Ad5uyuHFqG0TXeLofObpOqniuFxApz0FH/bVZfxxg9HtJjA
r9KPZbnDWkwnRkhOsRLBeGZ3EPwbIoT1YYoIxi7VH3IQK+vwBKt1T2ErxHZigR4m9YGgAs0GWgzs
vzGM+5lQ6Piym+J6w7V3PeUksFoxZb6077NP0+AZbuiOG/6v7GuAqzAd0WNWGorz6tvsVNAykmbK
0g3t/fQMvhD75p+HH5Kxh569mOf/MWzQ0TdSEunR0C7lZs57lbHWaUtfjx2gHChSqYZt50unKGjD
lvJ5Iu3JdzQjcdZKDeijp/6P5b5edsJjYDHsuekaErraZ7K2/lZ4tdinttY0+2FHpvoHQ7UONbJG
y7fg2B+a3xFAtnBCl0b9JhkrCTkVVDyDk0gwuYrTI8RgLmGLici7xvQY637upAP3vGZa/hm3Gdu6
klbpo8ibv6TsLAke0BATxQfEbSGqRn7raXRuox2p3SMKtV9ZO5jKRdpaNSZtA7w7Jgq2BA3hgGml
CO/+RRSeG2OV1GU+jatvk7QdNM1/k9J9bR3UL8XaD190rlv7gQ5KCv8k8w47IOVXR3ZQtIpH8c8k
xJOIBXo+ADZt9m5Wkzibys9vGpiCGZHuknGdV/kuUncXoxAtPaJAvvx9J5PwmRjyaOjlBAca5+C7
L3Hzo+gYmkgk/n+OlOVqhGGfNW67Pe5iviTZ01gaRzLHkVc31FkZmCPI4VKQ5B6Yf1iG2FtCquTP
hnCS0+k4jSxUBHTzSWM44v9945F4vV7kRYbB1CS6RPbCryOjk+DADtzQfEHw/nZkIS1uGvRPh0UO
VtoGpGhyXkS0nZ7/jou63aBmeC/Wq9q1YpCsFOznmaLihvsUBom9WNtYXQqUngKP/KIonhGZ6AAD
aGLkJxJBqG3WkKJuyA0RCpiTO9GGlcJDSWJ1Z4ByVEMcavpmqHQFyWa+yHI52bnVR9qqMB0nJqrX
Sl8rxGMVqQg4TyXcLR41Oq+k1aP4rwQdsgBRMWT0TuGZTWrfaqnAIvHQU2yewHwxozmLdJsi37JJ
ElkgOJSsqujS986afhmVX4wTntgbMMwW8gUUEAzSU7HDRrwMBI4H5HcYlgVWaFefMVJq8GKEzrla
a9S6KtLYFgIeBB36xiOi12yRzpQPhDW3jOYO3/ALJyaaFszOxgomNv0+j/hKQr46EechWtJAtxx4
p5zo3POXb2yv03EDcILvDFWtHV3NI/y2d5ov9KrB7pFueiFnjrNKaNg8W5fMI/OQB/38L1y5Z9T2
hy0Lgp/sY7RwCs3D/Z0aVUabtIF23lMqT3fjxUW/4ms5j1k3T5Sumxr5X7XzHbPnsm+YqW7D0gp1
2tW8PRLzgXOH7lKzxxYUpigLOdFjlKntkS5UciXJm0lsv72MdD9eLhPgmUjQK/2i65qHgaQB307h
YdREdkcXmSwDo6fTFU66GxaKsTEhsOEzOSdk0Ej+sVaH4jF+s+EKdGG73LndDAq7Xb870kFoKdiV
EJc2yjAUhGEH4Cyk+Rbv+dfO+Buq2JLhqzoXsN0rByqzCO7LWCj13Qmy9ydXs6ZO+ldX3hdqxPsN
5im+NhgFKz3auPm4W4AD5OYBjc4+tx3nPdFtUCURajZHF3ur+PUKQqDS3YaLjHxpd7MAcdovUtIy
PpBbNZDbOEAL1WWea9SUz+M/QZw3b5O6JGG8/EdMf+/eR7F5rn4cG6p8VWK8UTdIgXJp3I23EOK2
t1w1Vas2wU2H6aW+zC0ABUMpz6FAHSomMXva3rm70Fw6lX2RcnEl1k2rsOks6nr84r3XOb7HPG8Z
LD6pQB19OkJqtBTUrOC9b2fGI3iE8pzU7tB42yoTyXd+WumiF690XBtntEx764y1y9WJD1+dWVzJ
AinPZUo57OIvNsJf1HMIHu3TW70sdNsuxF1jsVGPN3Wo9FoBRS7yVsANYK+YYmSypiwAEDge3ITO
Ght2RGm52HxYEmm2fo4Jhy9zoED70QTcNdMm5pov51mXBC0s0Pix/CCNgW9rewTyF5lH+vnc9OGR
ClMVJyGd7LI93CGGt+6F99Dmx5CkaLki2wCJauCUp4jNsTTiB28MZCYzxGO9UTYfUif8pk94qmVf
4mlBi/bqEG5K1UMF2tUCjmJXLVBTirbvbYF7T2/Y8tIy7UKZdSdhzL6Cj0tPKvQKA1EIqpIoo17v
DYR5E7n5ptR2KsqOnZeLwqaTvpJNtUGIn0tGJQq1Pwq89cwP5lMNp9aoyHtJWrd3OZoagwRrOvbk
7/miMPX7CSZ+xjRIapnOpXEtz8Qk1gG6KcsWO8YZi4xyG5qSX7HtN6kzkKAIoGeSeoG59YJsXy2R
68QLH3CtQeA6rgqVuan+fnCVYJYtzMymdVU8P/bUdReZunbHGkH0hfoajVnfj+tGqupKijHyDu54
TivGob1goFwpPFQO/KxJBEfZ3j2+S9+dqTbhycn3bmR4YI1QAwNP2+XnHLdYXLMJnqqxGrh+NtsX
8VLF5zc40wz22sRYtIoGjjdWpD+BfqE5C7gUL7LUf9MlA7nRSmp9flc/tq9es9uUyB3yBxZzEJ7h
6OKWFcIttaBz1yb1W1o35fBS647c2ENW0UGl+tyKm6oFkn6Xr5AxmE4724JE3HMGn9kNHowXpgJ/
lJUo6lZACUaHuWefwXsm3NB87UxLYJ213YZTWjkruSIZ1SFg+lCL2zEopIt09sWLSq701gTuSO13
lCF5AKiEfbBwzqVVT29lNh4pQRclVPkycK6877K5yPFpXGEbj8fIa3w58kdvGqzaxlPhK9CFYJrg
XcwYDhbjM+GgGwL45uEHleuysO4uALAE+pkob+aVkOJCH5CUuuNtx3D5Ft7Pe0Fa/cut+qOU8dFU
m1i7OiVP8vusq+mn5MirOztas5ZFDTRZMG2u/3swtiJKgKsK9Ksel+nHC2/FnmQbIInlIV+DcWWo
lIYs64Eygn9gQwFv4AYbmPZawR1P16rhw9G/DwLSsm1iUvBN2WNxG3zJ4pyZ/Hwg/FFdj04DcDDI
UnFh81XHeXDLa2VleZ18f/XbVHILyh/9NynNoxjHJZldS8vBgF+kdPKAiQ6jS25luOric8ih2kQJ
JvbE8ufQxb9xy50+FAb2eJpEQYOZSHt4vcBl1axOm0Nb11hZSB0SoHiCHpbjptt4BeISbL0K/CaO
pXzl1ejgMunRl1W96eb0Mn3mHp9ZavuPtehj2sMF9CZtDn24AA43uga3o8owr0n5L5wqKTFRkuox
TyR3+gYLu7Qz1h7oA3ssmUwtvXSEqO4aAb5qRCmXK6DMpYVvveUhZ4fJRviUtgLAjJw3vPxrYZ+y
c4vDp07h/EpuVXP45vsWS2CvgqMmAy6YAV0pKDFrwTVWV3Q/x6fyqEFk929RRn/XbhGXLP4Y5rbE
ioEoWEDrCNTrqGjRgKIkc2QdFLqTjEG5i+ljfSSJuAYflR+xSdHe78PYBodgSHX3ljZyKSsgcgAc
fIZRRjPr82k9Mo5+Z/lVjvp+3ep99QXrPB6GrXmjLYHcXUNaaDwA3h5ExqCun5Dznxmw5gPtf6HH
13P0aHs6/0cNaV23q1JU0Y6SIbCi80BgL6hqrJmn5RdPMZ0d0wXTH/a3UuVHI6j9l2l1cAWS2uwO
fQ405wR5dnUFwcof0TgLqOGtC1YaFMCAMtR0Xq0/TtOKgWYbHjpm9hfUV4HrCXrHShIJXw93PXG3
okkLzID6RE61ZowSb87mKuQ0XCqLxz9Dv+7vZy5Hj1/ZiakpwLnMFjmhZOTZ//PdtSyNfdvm5H17
lfm/R9vBYvOztusnj1IjCgm8n+i6eHI2MpqMAtFQRNBpqdfzPuCXrzOzfiMjbgc2AM75ETASS2fb
/WqujcX8H5Wn/KY+t2+0t1h7MDVCxEElzuFkGpByGS5xNcW+tdp6OclER7sM6e/IK7ujG8aMGLdX
o/5ujFcIyqCacszmTbMNNrAPMOkbyuMpCR829U6WYTzmp2gELEksifgccggpcQRznnzsHfMSHnBj
Pl6OOi9hy4Afcckh8mz4iqE4Js3mRokoPjaYFQD+sXELko5Rxi1wJOluqzT92ooeJDuqQSYj9d2q
uTJjdF6/ocTKXBgtTZkSxla9EAK3NntwuNh9+rzG+3nO0/rX+JgQayZnMH6ZjYsq/Fm0aOtMQNJ0
xF9IsP/ezpsgGkiVPpQdUXEgcWZdGlYyv8jkGIAHvj21HpQFp5dxf++rreoKBqQRlqEix0v9UV6s
njLhQgzB6+pl4sWSXI9l2+AolwFs3jOpdhgo7N2s2cA+bGCAvJ5U7cdroamHEtJo4sUK1sb5hGin
FeJMphpnDszvPaL5Kelgizmrgy6Oa838qEchbgAt8Sq6wDzUMsQRlBy5nr4VinFWz+PTFSjsx1ID
yeYUP5Pa0gpsuOpMQ1+2TB/3m6W69+F+1d1HLmagBjUT3+nIePikVvTG+u6ZIxcO63twi+J1zf7Y
4qLMJ2Sb+oJOjPZAcKcvUHYvTBtIxSXpKDp2T6LwxwFdri06P8njIVa1KV//jDdqPYTslJ+2z6Gj
FiztfFEHtR6NI53RR30kt1d83u9zElI1+U6Yrm3L1gWglIj6IKUiqtBeuTz49y74YCC6wpjBrNgH
/5MKdpjRHJ7nhUrpH+j5BBJgF4t2/SnoueWaVrE6gztqeYR19V2qR8kWPLtEGddGf0J+8pSXLAwo
hycAsBK6OEXIjvW6L4cg5VteMfdztJuJXbFeFhXDOu74/iQveHpl1OHLKGWHoFeXE+H2cZ3FpwN8
HvH+tQkoiKUFeSsZPWwSKopixv22tO/+KBrS54p9dnpk1FJ/jO1khaou5N5V+HjUbTAxnQs3aXOj
lhcTc7k6dQQjrE/LBdxOUH+BCtpNBfigk4NLAwMOx9CBGHPp9YYjzfBw0Bl+LaFvGdwiz9xKA6Tu
N5KPyRddVT8NbzxaLre/08x3X6rawkQTxbHO1Vj9S2HuHqIToAGe5IatDoZI6WnDC1Gg7vH5hWG1
l9EhSGzQAt1LtW4On0MOuMsjVF0oItAvw+JILk7dbcI8KR1I1jr1mc3TQQaotUHTVE8Iw1EByhH1
M/WfN9wWkFKRUt5jGM/bnws6Hytph/i2s4sqc4Ys9DO10zrm88QCg2RI1dmJ0fjQ8lsreMbYcb1q
oN4lpAf9YWk8dWCIA39Zw2bDLIEouTqNUjHQbi+5EgyJJWl+sUxuuuvf+0j61FlFn+zrgyehJuyH
xxUj8bRnUzh/VccMjS6eMej3ifw6OXK8EEz2bXZz/5KFESeE7YVoz9Z1tI3pZE636KKJ/QPB7gY+
VmZqb1E+36javMJTCQ9XoHiMBe2iXQtr6OtIILxxtJ3Hurb6Xj4rZrg2zIxk6olvMu2Jd3oWbypS
qSBKsas497a5THGr+H+kBN0DfoL1GwYis4nghmNWeJCN874R+2cDltz6Zo0ha7sz/hA/Pt417k+y
daQrj1uKA1ryhM7njjr242j6U75yXgcRIo3pTgh+5L4MmwiUDd5Bv6w4s05relvgfmLG1fzeoNO5
8dumgMmzl7YIPAHaaqUVDGva6aXuoW/waWvowwKN5xjfoRPcPrNOsFyOvFFcnLECbNnDZO0Wx4Ls
KdslUVzvUSrYg/JL/ccixN9805P3Xa5qhypaXx70R3huudzuROK5LU05eIkWylpBtoMY2w/YcVYB
5+RUbrWWJCEdctuBCmKMIlBP1BmiDS/EF2ZSbZgYaeVUA3uReYn12oj1a2pxd4F2qSBQzg7iUAZJ
xD8dC3LmtCg5GiKIe5krmlrkkQKqBAke2p4Jyq9fzaYGcd7yZslC8tH5EIQdcannbDRU+CYzi7G4
ZBl7U9X7gObWC5TQRrz8fDeHOZ5brmYzXhXsIWkVN4f0t9izCV2Z+YWEeR8WeG/i4jWsD4ALxMJi
W+Y3wsplNirgpzh8XFBmG4WMOywwY8un5Mz3otEYFln6gajIlRowArEth9+GAsHKRg7PvLPaTJys
C2h1IhBMj+NMtDQJ9ieBRHC8UTn43cB2wgpPERmUkEIR7jWdQjJb0739QAx8IUNUpes1eHP+6VXQ
NkFlKjSmJbd5+rP6xltQqu4MFVL8UEbuuTMPwIunw60yFcPRmtVk8PDXlBMf5P56eJXh52+MoKUj
MXUW5YMwNsO7yX93Tkd+156KTNhuUsRGtGpUJWbm/cCSjcwGMlMBvPFSikUT+H1T+/rquarCnqR4
/3YztD5ESGQSZfua9GmwxKCkvyaUTivLcxvnOxnmX7Wj8Gj2rr2S5jf/E2u3N3kGKEQKcMCKd8Az
rHZHyMj0Cs1waW2c+bSONy37jiM2D2psv0vrbQXKEjq4jKZ6PuGnnmST/rR3OkJ+vJh/oDPHYU4m
R1wn/qnmp3voiybxfcOBltV3avf0RbZ17gY9fXXFcVsLTJZDQJrV9SYRziShQJaZgFhF9aw6wAOH
tbUP90at5enqj20Pm8kvAN4loIJ36Np3rB60SLDkguWE0CQVOwULpeFnVdQ3NBrgYdrdmQHsilJf
LHpfouel6AE+r1n7u4gl5Y6hT/pXErzVZk8UFQk5MaZwcpvOTrnjGQAG97A9S0GtgCXiHEL72HGF
+pMWgfg6T1Q0fiPWcFrVy9WhOQTwggRJ37cGQ897nUP8tRKWyx5u3F14DoP5AFlThew2x1FlAHaA
T8lHqf4xMlMG50ntHKPdl6Bx3OvRiyJrRMwBvmOyZhaVzJ8c2GC+K9WM1kvCo2PqBQlk6NG+6Hza
v8xzfGAPU/zrfipqMQg9xrqmOyX6h2u5pb3AMW+4gB7dcTHoKEYF9QhQY6LcCAEXLuR3tlyQMYzA
R2nVID8BkjONugEgXZTJiacWqhWDGBV6xTuOFTtBQ85ubZRky93dyHa9MGhGTuBE8dR/cMOAWoOV
XHkKGHKEP4wIr+eA7cTZOc4de5i7A9Q5ugbl/cenTlliCqqN8fMcgTH80UPP9fScLiALt0ulxpNr
LATyJouGsNbTS29W4zaUcIpxz+Ky3FVwPDjPHnUu9v3lTg6bB1axCuXmx7ABMZm/Nk2e6E5tOUv6
MLHmc/51MyaACuJytqmLX5suOQxTMuAEa6UBVj1NHb+tsj8nOG54qiqt3UiUwcDjAJrKF/rLnPZu
JWKiH6CxxUkN06oKdaOES+v3Wp3aS3zZxqAN8fe9ccJvAwwzx8H7KRPDGmPVWJu3tgLQkDBo/vxl
CsUxJz8/NSMYEjuL5vsvhNCLN8RwMfsuwJdtS5H2ZAJNxitkJ8l9VFNW6fu6acj2ApcVFEQjSJaX
9zP/8J3Oo2ytnPyBwzL9efKhGEePR2cK3M8x5uHLr3kWyiuFMWSsOiSKz5Mx4fwMtouu9J9AcIhw
VBfFNBsqyLSmj0pcnSElOgMForf9Pba+ybyEQXy0bJKVvDQV6F4tntxDSWcMIqcIA0Yl/7W6zLlx
dKwh0pJVBUFVcexPmLZwlSkQpN4AavzRFfUKmXEkkyHkl0MCcC8xcYJ/2JYC2xwbQS4pesd+gIMK
vz9OQel19TmNK4tDJVBmCA0ZNmqzDZcnZaftl24AnM/0BZFWKbKsP2vsI1RhbZalu1qT12nlJw0B
wpuKAC3AduxNnQVpmT1lI6PAV4vDc6rayRMvSJlcK/BV45rJ416JlyXMQTymGBE/RJ6vo31koggZ
9ihv+/1q8mVm/5da8ZZ06rBEymOlKHIn9hdHEv6K+1XbvQDlBNXuwII2xs79ykMGTP1BcmYxfj6N
/5XRDqn3YU0+K8E+g4lH665mGoHx2B8rg+M2A7Cao/UCrGQCj11p2uD2R6v/LxKu5j7OCbRmTMbG
QI13GjHSI0QM+FK+0cQ6RwkvihGf8vzeVZ8diJTM/OGuQQQVbKeLP6L2l+j8UqFsYCfLgLVgDuwj
5IpCl19szOC/bAxlZQeSFd6Crvw/OGj32CavZc6ug/fsRfERzFnqdnsOhmo0y6yoTHU/BPyxi5x1
R9wm2kOWU0/+3uNKKIEwyw2yV3iR61a/ftHLMnEDesuSCYYIznnPOC7RGFO/EPrfCiZhotvx5Z6W
x6YxJAPx0jVz/tbeu+WVSnwDImZFu9UMlGS1hYO1GVfsatzzHSEWkP5JFg8/9XtufnG1g1yUqxCd
uCgpVtJyvyaaBbNLNqlo1UauFXxyVZTnVsZSoU4Q86n2g3p1gTjDJXhpp5CkO9iX0lM3xkKoFWty
lGMM9pLbXHjH51mJRTi12TqK21MYdUE3IujiczqkeyOnBJezdrlc2YgVh+YtP4yhbANtcxovTItK
N0SDfviUIye0ABh0ectzKrnDkjQtfKj4PuENPmdgmJMUhWvMUWFgweaNnvot8DsvHZ1BK84pIrb3
Z2ggpW9PkCgVK3vLZck0MV2eGFjdz0MvaFX2ZIwO0+DywQeB02VRslV8wtsttgEZqmJx4r9mxckr
G2TYjDWG17jNxfmwWJ9gdgHer2ujh8Wj8hvFM+VfevXCoh1u/Rfr4KzQdKpF0LZQunKX+u/h3uAD
+mZWstNO8OkD/tTPxYfQVEsLAGLekvsM4HAx/jZjCAp38KbwuPHPysKMh4x4LvZiAVA+YN7VooDd
P/yD3yn8yqrV7xDW+2dUfIjLxEa3DYXH8Uli4sgN7wiFVsS6n8Q4y3uhWu2zlIs3Bs1445zHzAU9
kQVF1gqxeTigHhOYFxFxrJqb0NCnJJSwpQpMCvap/dXfgFTBX4YiCKiBAiPH3Ff/CAV8YnN7EKl8
DOPmwXc7xhVdJYfmh5rv5l0VDDDhA/bXWPvNg63Ht0KuT3pwejRRwTTZ1jzY3iIZ57yaTiaxFVJF
zKZTk1YfDvTvb7cNJEgi6zYLEz8SyCgEiVRYGZbsiBPzIQPDmY6R/Vbc5iSvI3trWZwNA5r8WbGk
CXdkWFNm+xHaQGq/WCR7hmczPCj9tyxR2cbuHCBmuQNLdIft7wZj/P6WNP/If5fHbgQJSr9+BsyO
4l/+3pG3hcp08naYkjrheXDUBl6LxohmjOCdMf2GVw2PkM1y5OSllWCZJup3YQXZpPaPrta8Z0GA
Kwxuje9hVFWcYbc9zrDsP/qnl2345Cu8xR4xzEktjSUPJFGWDB2bn97Kj9Z0Bu/THeNtYCdAFRso
1E3u9IchxTddFW/v/W5Yg3FrTJbCSdQx/wY97XvNK0OSm3q7w14wycIcFDqPHGTko9jbO/CJzWb9
ZALhI9pJu/lBZx2NAtFoMWRlrjQBABf/pWgXyYG2A+gsqNcoXZ8EVs5Dm2OFCUTIhRjbPoMxKnBe
WRn0EDOfzIDhXzcLjjT7wzkJZ8G8eLEbL3H4/eo0CPW+m8dB9xR7waGlSBduPSVPpb6zL7btETzl
cGvEw4DSGVpDKPZckLUjEn0lw8VrN7pXYY1wFC1sk3HOI1efzSvcqYsZrSVcTSfG7cB8Swwrs2Cz
2J46+gF6Zwg04hebTSzsTOT2Jq/wggTEv+6JfuAsfBfQz7uWCkaK/Xd0rERuGFcmQH5JKVB4RLr0
CO76/Vvv8Rwu3f9uJljOiHq6K0Ulwur/OL64AT616LeqTBLX+ruBYBHhtLo4KCPxPyOjGtJuJkPd
KJmHaC03kFi9bza8ZQ5OQcJ5DkorDw/Yws7i3zvLeBtFCIozVezaTU3GHpGne2Oy7YooBQZQWaGB
vjln8aNunrdaRFuPCuMvL5U0zz2jsMGW6b1tJ7R3B42vab76A675Tzxusl4H2PrW3IT9haN5nIYn
LO+pxZXy2z7Nk6dzamcXkBSiRTKmF+G087EuVKnEG9v9PgAT2EyHQmBJLKqDsd71xFP+PYxcCnCL
o4AUGW1bh3d7b2pHMD1GBIvnfRdkJoz4ooeYuyn68doHuVT+y1nf9H+YkOum9OOY/DTF35GZG/uP
d0PQy2yWxzHd9rrcXOfecwO0Vg7oskltPoM8mNRMJdbbtgKs7IGz6BVJpdm/lBw3XHrmCF0Qdoh9
rTTurpUAVTH0c2jzhJ3BnMDIwynPcUYJZoKYHZvsoca8GoZ+SPks7XU9nAVfus+WkqUCl8UP6aYE
cw2cL846pIatFdI9LxkObnDgG1H7LQvX4js0sQI6v6yiiNGg0HoMrkP6SrZqdDhpyrM7VKg6m3cj
M9MoEs3Rl+RxkMrQPpdH0HGT8Z5jGwy/mMWa4G9Caibx3+8Ioz647VnjhgVUi7jM1e2X9n9AApy7
6/2RRnThsu9k+OxFGqecsWKQs9+3482IAk8Rd7Ep8+BmfZz7bn82a7Cp9/G5jtwNJ+tWCUI3k3q7
L5YtWN57iNcuUpNaxa3qlW/YDJom1JzVDfd02I9zZX808U/Y6V2HE4Hv5kPPqHVGA5Ebdk3UUmxc
5JTIneRDIHiF+W2k1mRda4ODsSRu26AFU61hiyEx2eT7hB/lrcJ4CLIKNqNT0zuBOt4IvMamhMSO
vkA5vhjyh0dTWnrBqmJoR6vhq4B3HTuI/Oa1e+eI16rEEJhwh+I6hUGKFsWfSTmJ/5hHCH1Mf3i5
1yRDc2kwZwGAhevlLODhGxGxdg6b4EmOkZG/q7VAmpNunY0w6wa9hJGkac3Pv7PpxTfk8kcU+3OV
Jk1vm1Sd+XzG+C35m9epHiMIlZTIOQy4/7b/VKDYYJbOh3/IjWs2axiSvyGJD/YAnaRowMXLWoZj
JbNhZcZmAVQmtioXu+ZeTyNuN9gBXpAHpSgJ377K19Bg3H4ExNxBRSOw8+hZwTf16x/wOuNWrjoM
71mNb7oewGzwMoe6EKh7vBDvojaEiDoq7HrfM05ZS1hf81yVvjxm6HJSRn53I4jLUr8+RhIEFj4x
RiA/W4flimPewQusvou/A6/mvGjZuZnSiCmxtZR7ykdsfFCVQl7dz9ISRX+v+ne7hHTJ5/lmeGNn
9e5gf09ye8SndoLP/h8I8ySEM7jKawDL2V8dZliP54MK9FpGlTC5ifKpQw2OgHnJm+MhptBpBsc3
QGOuu1zQ6HBTJ0Ujl5qzLWqHTthFhfN/CLe0WIY0pggZh6e1sSDjEL7Cv7JCOEt/knjVCdwyeDNU
k/MQWeTWoXXb5mU9rflV/0wySUxYTsKP6Xp+wdmBBPIyGMLO91Xfg3JT00JjNsi4mwedubsespry
Evx4w8DZoyKN0rTFql6hiwlFerKv+Vl5O18PtnJ/sNy3DimtsnKpCVJ95t2V7E5hciOmBkELY73i
/lyADmKEKqMeOIuv6wTXZPUKm2R+6eVZNBcwArr+Uf7zS03qTmhxnRSUMjWGiX9afs47hIopVokJ
NxdpguA1hnu/Eo0lyq0j6uswfk6ueVd30BzRUFXsbALLRwFsE3TYIPvSysyajZz6IDbDn4LPT8uX
ewLrt6zZnHaHS9sD3vKnK1ZQ2R9DrRZm5VYxZIyrC5YAjB1pamnrNcRJb04R4i/7H2yt88xBKdfF
NOzHyJgI0Gwj9I4rfCHOMCkEUeEPlcCi9nfAp4aqFjO8DNs+hNBw8FsgtlIWkrwhQxA0H+oZNiGE
gEX7SBUMVopphPOS+cIqnoTbIzvBmFKsIvHrpTLqyjXn54pas/MrGh68IjSUuNRw4VFLA7vTd3kf
MDreI49D7ytBLaqtgzg1yn6PqgYg68l+m3wS2Z3MFlJhLGQO+55pytRCo9UtkJP80ihfGOwvhDO7
RO4mYCw5PiWPDlsbPVrJ/UV16FMg+x78gA6/RJUAWLBSfwMBPKyqDmCV465EafsWcVIugPswmJy4
ixfiVCrHOKf+gi3lwzd4scTkJCfC6ufaCP9p5TvDyUJMDabZbVFlIYYwViAuGe/LA++L6iai13HO
lfF4oEdzXxvLojpaoWt/eEWnC19YuPsvExcq8AtYGgcHZV+35gvjHt17OxU8xgipffapYPNNGV5Y
047C5JThDp0Jxu8A+DQjimC3fx2uso6iWTZxnw603SI+ERP42W3y0u6fZ5gfm2IyT6iXZH4gRa67
S9Rqm9Yces/Tt2KNHoxmbYEXo1LkV811aC1ZChUnNhicuaLt3ct8u385ZCyYo6O9vuIj3Xnilck+
8Q2C8HsJ6jOEhXjR6i1lqDqqf77pFudGuK+EkMXW1Yft52IWW5ahZeXc+EWJmQR7xoLtHXaQ3soT
j4psQGvrf9TpMbQHcaxbFTrr9K42Ay9v9BFprHJdiX0QC0+eXIrsCP6mE5ffwjx7KIwlMIwolfPa
EM2bMVvisU6zks/5VNOZq6e/T0GPVMvFYQmzoTt66H9JUeKe3zeyTZYn3EsTw0qgTkhzrkVhc5u+
ByWyDAa8EPa2l6541WwBo83a/63lLWpdpRmPoc7AxoEdTjr5lm48moedyytYd8KvRtN4vdIWYWMc
pTCXiq9UdOOxKPmGg/fdqGaKIHgMpPlyAtJkP0PdW5+VrjfH+IIRvQsmw6u727UoQ+6K+FrpmjAE
DAdNo5+Ks2ahF3od8zyYDJkAFcpvMzYla89h72H9v7bOQpfxPWV3OsbAA9iXiBdzZRY2bYW7pVwI
2Y0uK6ogUoeB5360WP1Y/v61lJBbZ7WhLXGubcRwbgOBzm81vv9iqESjsVJWVCyOJeY9sb+9zvB1
QUNqlOTAPOoY2HmNd5kbGNDU+VmZ0lV2UJT9gX7PpkS0rEGEZfvAEG6KG5zpMv8Zcf3VacM3REjP
qDvvECTEvN+lq98MZywuBV8gD2kL3MZte1d3Tg+gnFpGmyBkCzHoldQrsIS9pyeI/m4Y3nI7//K7
aYw2E40BQem4+7kOny8k+pAyzq6mTMaro7SsF3GBsk1i5xFt8NmC+VfTILKDF6wZBO+m9ERx6lak
r9prqAKI6A8BYddTvyhKmGk+Si0+ueFVDsQ7lMZSvDBzMb2hRmSLlLdYU4iZS3f83LvDwu/enEyB
B2kL2Bz7+MkMlIH95u0fAfRmLabftUd+zxdozpmlb5g1b5x1/4aSatWS+yUs+VxJLLin3m0IRA/Z
S3oh8tRbJDSXlqeb4OIRTSwxoZMypOTukl/o6nOzzoYSPRQXEztRMQQi4JDYdpjPjFWCRSkLsFpt
Y/Ztj1K2Ff9rq4OXl5y57+YEYxqkZMaVD69sj6JTrT1W0Z2MjDs+Ms5dVgwhQOrJVs7jYv1aNTyp
jIRYZTzzxotKahTHPuS8pplwQP4S/cudk0kjxVdYM7/28zUVUgRMkF6WvBBqN8ecJngjGeUL8xwS
TSPbQYcErEBvLwA40Qgihhks/HyhM2NZ7TSJ6fE2m4r/8w3lNwqe/eSmHxvJ5Wd34+ahWNgOxLqJ
68sOTaHknYam/PDcCKRodYJ0MYrCyijSXG76P2YzUksadLygZg8NdivaMUr0cJB+0MynE80tbCLd
fmGqlrLCZUvItnkbsptWRSVLOehtjq1X2/9XuY7e+Lj+BrPqNwc+iE0oLuvTCvKiAFWO2/zDuIWR
hG+Sb8S7MGGiPFICSsALSqz8+b2feKF11yIRul8VXxzuaRMiL7KX6SR/P2scnv3ERmUqgJx6oPfz
YbbLMwundv+g0QZsQgk1ZGYYevt0eslZCOw2+ev6vi2RRDGvmjtzjunho5D9hJnkbqWW/WBGwhnx
8D2B1wS3mMCBxJfl9eKhsmTRupuewfnqHaMv79q9xW1q429+OPykgY9j3IBeG/4THyg9oPj4YYtL
qog0fNjcPvnbFIVDrRRdHL1UUnz7dlcRadZLAZD0gK7VZwfWFPgQbDrX11BXMD06Ezfl4NryqZn+
AsVtrWSrM/NnGUrP7DVLcboTj4f4s9BXDcf5LJ+hKq4X6oDzUPo6n4xx/FuGOFX5ui8WOwG3VOdg
z1oyDhkHCH/cliKYH9dLB1HDNQ6klqQj4N2tlWzzDy2C26aiXrWdyrSdQxcGW06sadRZLJXA3XkS
Vcb5+dP3Kq5+fk7iTYQrMlQme/4JWpsZW6PjYqj0+NNaahSLZzHQ3Yj91x3DSTUsBWYZ34ezKtYt
KW/WFwdoPsiLm6xZR4ZKrB6wqKQi00N+Je6Rx5xe/MSQVUYFYFio/CXNrulCjG1+HMT7dK/cM2N5
odmjVklriO6ICUkryxTstHa6te2Tu68sYIdz/yK6Q5UNqCHnry7LT7pyBjZcODxR6x0zl0PslqOA
GE5nDC+Lsp1tzkYpZXt66PZhM4j9HuNzZAY+yWyUUnPUrTBM7/LyEBexVJxrSnzHKAdscrCWwvRF
uJfI0gMrHWzm5qLRQDJPiUgQurgcZkbhsUf0xk6Go+gzXytDhnXc4Y7MJxzD1RertngoMRpWhwqI
Sjic+dCaLtpRqw1/FuzE0RP5iQj3o5LkyZIEvxOQDSNjkehEmRnC/l33buzI9bH0Ey20IBF0Aszi
+jyVEQd8o1uK92YfceLrEwWurrmDeL4JkOTz/zkwg0m0ylYYYj0CUmkPKdGAxsVL5k7tXYHzPJGs
KhFcazsKAHUHUjvidGAIeOizKlUd5GT3X5vKH5RfVgkhEr/zr6DRDsOmwVg0Pdl7yHS3uVFo0xms
krVXjONHsA8ZtBpDrxu1M6Xy4CNPfjHSNXkjxFGy9FYzPpxA5lEqNSvIVLg3J5A7U/Mb5ciFotN1
46tGYLwk5FIjMk4hz6AtOP8mzCR/ic0yq1WGX+Lae0siuT61zCfgspop/GbJj0iGLPsHHqYzTihq
yHSMeZ4ExtMc5F5OgCEi3DHvsUAMamE7xIB63vTeGFuS5JbbWORxW7buedWoAjxewrwr1kPxFiPI
GDSgET5y2kCDjMy2fvOsJMcWaQW0NU94kvnJ4Ok1IcZ9cxRIAvx29RiDfnZOq2aZYl6iqDhoD7de
v4whRDqxhEO2/bsR3JnQ0ErrUPBq3Sc2Q76fTyQ/XYdVTmqJ5M2n+ygQZLlWoirRkbRFXZwFsbvE
ve731KFe2gkAlisUa8jVYKDUmhcJniCntLrdtte5uSxn4D+N/WepNtxMtRcuoGF8GiPqjv02WIHh
oSMELp0W4NkAote3JVpkL0XVJlDN8zNTpC537WFquM39Jvr5SDHjhJRZuDTu23/rmE1OI0+bMp2k
1a4GuiVhp9Lai4JJNo0jwcCoFrmPgmuZ4znaEpHE7g+m6V2v/2zDpv19qc+MzF9Ukhp9lrChA5Lf
bOeTatgH1RW17zKULLEW5F+xOsGerrXKzk+Gfe3MFS/jjfAN9QAPXTQi6qyQfof31RyOKvrIhjbv
FufAZ+d+gIEp8Py8oLdDgThCay118griPFjxN4dEWeGZNNczeBFzZeb5plr1vZp9iHLXakqlZuO4
kQgr7xPOs+lZaq3GfaA3y1b0fQdJJYrVw2FN0NnfYbvHVwmNg9d7/TTEwGFr5Ys/5mnqtmc8HbIp
OpTvmq7EN6JE9g9q/VQDSaTmWMRCDPOAp7Pqxj0q/WRhEcuQncHtc/MdoL7F8sgHDeNQK6Kce0Py
txqm74PNcGRJcsuO7fYsJQrvwHtN8Jr4TPRLkqCcSR3lyA5kWo5/nI7L+bQmu688XPoWOWLq9fCi
U2uhLu6yqz8liEaSk1QMgtQ5SKNugqlGbyESly/DpAgOUMfZ0TJqQIYQMag0bXKBf0wNFydxPkgF
njAtlleCzIVfu1N30FiimpKJoh4crM+ActEzwm2XjKoZ6G5v1CU+6TQEZ8l7bXOnZ2Q7eIYLdoPs
5yFSFFYgWTaAPuhXVSy2xEKhKrrjUQaMC26eE/gIg8pM868oAeghOTxzslXhqjJMm8H1rpOWJiiz
osXBM4syUrS2ccRHdIF+ixmucdzBDnr1FyQdAF3X5EcqyN9DXWkPEduS1QbmPQADSheMAQj0ZBFh
PGC3E3ErhfOKkF4gWLPeVBXcVUsEINHEKlMOrEJKjy165ZkeJfFY8tD/qwHQRq3eGnKzDdmCSJM2
XcMSoh/2xaXfWX2xwknP4VfC1JnIyB7Qm06wzg/HfJAYxMXrPUAzleOyHmJm2cnTsdKKRItI/jAs
r5byKsf30SRcUNbjk4xvNJVCAaPrynYUiLP9r9TwfQvXviLsc1+XBNZS6Qf+/bWXz+mBR1MDgZat
/+j0267H7WN18PEfnR+PsCXuD53cudBC4+7VC/yLYnJRm5lwi7VpAvEb8WpDCqXP902p5klph4Jq
OozGOd/gmargpVJWlQu7Lmzz5/bDUk2k6iD7jARSoiEQFoab+gqORu93oZjHpBjaWUuvBfMh/ZhB
wf5spHqNdgRmdC0myVODwBLaA7tRfu8/w5uuxVET2B0SSLoh0DZgVZwMm3KgEQmc0G39VTelmRwT
yfGUfwtqSTVPRZSW4P8KPIs6KaqRuO4ShIufxMFohiq/9uv8Y9W4dUxowEgn1NnVRGK22ALAPeF1
pLUk31JztpbrafzWsxqNb5U4wBH5yLHhw8m6k8kc3kI2G09Mg+mf01V0IaAc9+ztA8s37IDsGl8p
q6z82HBzMPjr2D275jgizOMKAJHLQcSGamziPjMQ701lIn8l0/doRekFi85y3mlf0koh1L1d4pTd
paB2Vx6HjlrW1oMbRxUhyxT9NlwPe+EC1skntR3WynuU/6vPT3TYNHp3Gi+JlFnIyznsPLuXJhta
dlTrdMOmOxW05fd+OJybhWJUhCWovVXv4iW4u0kaDWn4aOndCEBfThq8W5rz3saEs9UL5cyYOiy/
2PM+JMDFD0As/4zqNChqzx4OGou0vvgOAZ8/aFC7yzGBi5N2qisdzjLEe/c1xtll/3mnBpk0mnaE
2OdTT9uXuuuhOTN3ixhFs+n4f6/ufZOoK8ofLAM5VTU8iBnBN4Yi2mbiyUojnGCm/T3563xCpIB5
GJbb5xnVqAC/j+VEqdAm4nF4tpTYKl5k1an9uqfy+dCRs6IHIoDWTTmCyLlr4Au4DQdiNTUt72yE
YhaTVu5liRWnB/iqEo7HNXUMUu7rdus2Jdf2W3KSPdJ2thGR0bcYXIcWc1Fp8O1BDGp36ienaGmI
0m9saWh4ldoiD91kh6dbpGPBZryXtySP0aV69vlIEAzY0LOwMZCBJ0jlRfkS2xhKm7yHHbnSwlr9
V7R6BFimk6ZV3ig/P1xLW5+63ti+3OExiTYcP/smo1ycyV0m2NGt48EQnZUn0bs0GaaRa9prqhza
BmunlxMyff4zCsnZ7y5Wa+W2FVwnA0qEiB27Vi1lr5stk8QqHKmlY8GjB+acEFZs4G2ZxXz4SdR1
Be9Jf0+YCPneKTVzV4/KnNyzQ31W5M5BiNrNQ3rGDd9Xi8QlxT40HWPnWtSWjTUin4X9m40JUHQc
lhP9tWN3ENMlRgoQHxrvQVyC3QSOuae2yK6dqr9r2Wp4wMoEbpgNfzULg+CC+n634lrmuYGFqkNh
FMPqgb0hlFzQ8WjY3lKmrGz7MuFKQvUiuJZdqvuq4WQonugNNNQ0jTLlQL1DDoidOaPpks0oMko8
yUXEEe7796b4pg9/XWgRK3erOEUBB9psFZJLAvWuWniWS+QgEMzExJGLCktauRI26QyfsjDC/J4f
LjLerxm1HOTrpoWx5i0EI0Z//bW8xpmMXIkdftKe2N/0B7ETNAJ8kAx5KiW335hvQ3Ttb/OdGXzz
TkXZEi6arLsltnjYLDv04dUSoWr2tjG5D+j+s1HXTBwA9IhGkhfOacNCEfw28L6NFdHdNGLUmtNq
dsXDvuFFgHoe3XKJY9qy5JyHYyGUmsVHR4ci+NFhfXg+qyxhGVGsruoPqLVTK2qrsfu04FPmvW2J
ZKBvRo8x13tGoYF3T16YR8FQuzdfkZpzPHWktLazDCotVgi9LzENOKUEcWM/Wl8AeJsCUMWe/CXr
A/6P+apIrxpIuh3mQc1nLPNz+y0vxlv2gdCbEuL+Ga0J924jeYYUQV6JDFRmEUeEjNG4OYCwISIq
oHHQrdoKvgvTr2/oTE12+GV2q3TJfUpXljBHDDl8RgiWid8uV+YOALms/GoiMxX7r59knQjHBB17
WsEjHcNGXqzFvwla5cptiHUm2wU2uczkVles43HOXLwO2VWiEleCyFI+p2Qbj5J+8ceXanZE2VLQ
p7FNjEOX/l5JnJ0NxdZHSVWmEexEtpktJH0ZG2EbQW5SYZOhHKN3dPyoMh+qCl0d102ZOeBydd+b
dCFYN78x2nDA4RvtYQtn9/bFRmJcjyeZ6XD9gRzqZ/RZGwthqXitgJvL9wMrnIbHHfhEqO0O+kzZ
t4FyQFz9MhG3JlQpkaSV1m8AgGeWaKInjA13caC4nA9LTrFbH70KtTFg6h7WkZdgJKSfMR/OblK5
sxWe9eZipmbgpWXxTK68zBaDyB3vTkN71aM03unkNlafgjMM+XD99Y86CrWBRC5898ejOaBLQcN7
+1twQCGhrtx/lDM/ipoQByqyoesXJZl4auyzqS2r4TYtaO7SM5Ipys7W0jwwRA28JBdyHH3iS0qx
jjC2OgBLzyJp2QnkUF2u40zTYGRVZ+7AIVvWvIkNaVMrLU5BOt39TdM1GnR/kXEjIAj5av/BHvFs
Zwx0GRqMAQvK7mWqXpdP4UmR/4sUjweGCeVBInIgndxo2NrFdf9SKtiXztfyYKNM1v9FLjgb/lj3
pHmEmG0hUF6WN5TED1PYDPzGpfWjnlTM0N7FI3tl/V03WPZNO5JfzuL+xyhSg4rpv/xV0Nh+ITRH
UCYARVBQ8+qxD7uPtXxxTQ5FYvAjQLy0M4alEPlPW/ilkh8H7+/VXunMMroZpiWnfupeT73g/zip
PtEnlSLkXZyzieJRy4t9qOm8jrVY7mSd4zn9ViiuMDqXA3FR3IDDrcUhYZu5XQe4WMi0OGiz46bZ
GlNx6tjoe5HLqSz9G6FuEpJAC6x7pFV+HTEeRGLDb1jkD4PYcmV4FVo0NzAaKtS2CAFBDOod93Sp
HUMMrljbLFeSUfyyk/iMgwEbj2/rE//Al+XsHxLFLjskKf2b8ctvTezMzVva2E56NKFpmGZC4hIa
XIllzg/vUo2P/cdUNtGfnMzyTJEmqwcP28Tq7Q6f/ixXmEe/amOkYlhwHShaBk3ZkBHJ/nvl4SE3
nAxusNTGwsNjUH1j73fOOrPBxJYprA9Vc1Choqm06Ms1GrSKrAfq4oCk5TVj5I4GfnRvdRA5q94P
tqv7eiTvwnl54avey5ALTVoPQ9wh71izaXyl1pO2YuNqt9vJmiNZCUYHsWHS/fgbKpzhQSMNO6Lo
yVlW5NIVm8B2Lzj5FGrYnOZRMmT6sWNHJ61yyde5rZpLBWmyXS0tHEDe2d0Tyy7TjeEJeWonD4kU
hUmyrPDEs5XbN9PBfEjY/imSZgPiujbR71LduwLILLzWTPmRWlBPunezh41qKi+xPbrNCuxTA0Jf
LE/mE/D1IY/h5CIg9JgOmGEIcOLvR9o6LsbeT1qyHwGOZ/5BZQF7EnaCQvvAICiRKqugKs1QL0VA
R4Nu4+Uen1zjN9L8MnLtwuOCVgUqKxwHgjHoOCXDcm3nrP1bBU69PZ8WvimDcY7UGJ5Q10KRnFyX
lG/wCciC2Kv61ek2J6qXT+T2P2Va2Q3OXJnKMBSw37QV0WlRYuyJcYlTH5j3mQV8nNUdARnMz4yV
GHjqTxBPFRp2FkjnWRWj2Yr1C8p0XuJ6BE9scQA/o2eMFZZNjIkqKgzMdbG5Gg4c0YnOklga/Dpl
tf41AJ9v6vK8xK0h2Z0MsQoFsCVVJoK6o7uCGDNxOa8S2eGFKcskI2l6tJ6kun8D4BP2odLBLtBO
i/JkmtEOksc3wqaAOcERklXSe6eTjwMKSKpNpnM7nARlpvop+wCJMcAi85PbJ8fVny4Tr3sOsaIB
piDvpoHGQ6NRJBuSRzfDcZJAUXKYDSfvFKNrzaVNiOq/pZYOrdfBie89R8lj59/gayeRw9VR1Xpx
vNcNbX3voTdBGvcDnmVgaHGXI0QHr6wMJXCyU+/pBxcGruOz33SaoPHUHNBrTn3GF2YRdL3+ErCe
LDJ9j740CUmq4JL2MsXk9Z+9CrJQt66UyRInqBQTcVyEYzybNuAWE+nPRICiw+4fQvPX2mJ8pWVX
vq6c+PfyYJyOzge+72yMcU0I0vIHsLTNhqcTpIGG/UaE1Emgq8k9tBT64PUtBdDXDT1/B36FU3px
LDy9nyYL3OC1MjP4EV3cJoMmMU5O3e5NeBR2IDk5nkbZFVmrQt2qJ9N4WrPL7GXv7USHQuPOo6zT
oZpcRzL7lxOgVqlrxIBVN8K8xP26CpzaEkdeC3VC/VgxX7k5bbLTkZRBAtJ8VhyBN1RUPDRyqI0I
AGZFqo5YnJ2mPdaXDoY9heFmONRC/0rCQ+JBaai9KUxfQon24VeFL3V8Q0yivPJcWx8L1grp8y4+
oz0AdGBC9huVSH+99PdXgjmhHRuh8hCtUWRdOLTvgWD8rf9PcmrFkzjrpaIOdhZDDVX9Fi3E+5ex
e32Y1Rns2IUrj8nyP7f1u+ZZ37GHz2gH80ipEtnsCE8bflTCFNPzfWdlXVKwUNVUJEeaS8y4a58j
b6FONXK+a7dZlClIobb4uE8WnRht3hVDIC42J33Su+iwPaUehHT+Ph7GL0vCg4wTzXRif1Qc6Vav
NBZ6rYUZG5SxUXS88bG6kjJXRFVlciIfndYSTSCgLjKHOfOUUP60eC1gGICPiBhvYdGxo2GJCdjH
FTNJ/UAfm1b4crSGA50yu/FUj6Datm3L7pecR5hxtRa7vApDQ2H/nw4vl39IAhMSeZVpn0lk0jFh
rwH84H/6lIconuqYm4WrZZ1jTz/glYviUXmuDHZ/HHv6Q3n0EqpKO+aCSojQzWwd1Q27vnpb1TKx
zn983yVh4sLbrjdRdFk7CVRTzxK0zPPFb1+6+A4Uk5ZnMGANePb3+QSFie6WatMffkA0d/kx+2ke
FM64NTeqVTP81Bqtc1YlFKiYz4ZG3gGOKsuss4nZ0mbrAFoCcdZV1/iYx+TP5gnllKp1P8jm8qZj
YtQG3eGNy21XW4vr7JvPGVC/ikQR8z80KZNDMC5Nb+3aNlTBpI2lKmpEDj6KEQ7i3119wo9anHFK
t2cqiBzDKuuNgjYy6f9DVwJItuNZEkOr+9GYuaigOO8N7AKalRGljVEY5caAW6HsO3nXPgjx7m4n
vxtnKgpIeNMYTEFS9MOOKRnEj1rdeO/Ida79Mnv2YzO9IZm4QePsyEToH4X+VezZCtzoxxZXmwQg
3g4+azSXgClO9sj5dXquqHhlQd9bTeahNoxFMtOOeeZpCMTiP7xaoyJP5q4+TFKUb2e0VIjA6HTJ
Oo3JPzNWYtcXMRzkD+2z6zRMuPCweCTI4UR5Cylx2igovtv3IFBZUOJaDRkriJ2MOJCLe6JuaKZf
bspSpb6OnwVljrkJh2rZV8kEZ3Arpnn8S+p/ezMedXnIlsDgTHpqc0NBbiOsluiWldlCtxdb8cVP
9XXbypSosJM13EkScX49/DMeVyFqdfDwx1p14mMO8AMfPLsd4QoPNtCdb949oZKZV2bKsKpNBKfL
Gd1wsoPOBgDN5pVNdcp2+1Z/GHrEHhWdsKzz6TKlFe4RTiBKAVh9vXApHzr/1Lw3aV3CWQeJrXK5
vsJg18+BSXajsLs55+ZdLmyS7eqM26Zx/1Mn+PJHV2SiPGKPmBmRK3FXKHw8lf2PY3bKu/+YtsrV
JbDlGmoJCtONxXNyETNcQFdsqeRiGlzRddjgQvsR1e1J177tDsLMNTtvvSLpi0Ui2OLG9wePWLyN
+psNr6gRo6rQW48mLBamCqtq1kDq40LB+Vy7j69Fo4AX0mDU3XxBPnyvL/BnnYgclARBW+6PxkF0
ztE3QCJ4ydp2iEv5PthHx5FQsJDeePVrrzGCeuAu2X9jjX4m/tlu9hE/Q97riLqAouWm3oXaUX56
sUP1WACooOnDttfvuZbAVDdaZIgdXwltuziu0BwuwiE2AOdZAVTDh+XgFw2RWjCMpZd5DTzhQJbh
1pEhiJuMHqUqNJCJL3yeuIdBW6J+Yk/VeWfE/CFblXE/u/1OQZFJfDodFzdZ31UHqhCj2761yJft
b2WjmMyJmetpiL0wdkGsmspz6VZK4eKsQSmOLx3XUNZ9V2loIyZO71Wegn2+EX3YgnhzHLidyysr
PshWx1ecMXCMzYO+nCKGa7q4r3B+EOfGJTcCehwugRq3aRnZci6Wzl4IU2g5aVKGsBIm3W1pKiio
nKS/Qhnwm9Wri8RLeOyKznZT2W9E8/ngjABR9TfK0ntraOf4jcbx6UgmSFzhI/sN3nxxxSGA7p1d
VhKdu07f5Q00fpYRDOoRtPDC1/fkJCDy0JtSOjFz79GUH0jL4HUj4EqeSpoiPd/7ciskNrJevuce
EgIxVAuJQ8k7H23AjqYwX2lJlO2/XBFovZmWRXdI5Xa2wAsUAX5WUYqHZWi+FeXXM3yJg3jjj+WL
lvjAlI6wCLzIzR4HaismTG67Ilq+DgZ2vJgJwJsSrpLItGjCSEVADZJ8t6Bqg8xUX5Z8WVrh629C
2T0N0qHmgWRHoNUjYjt5V3X2H/ScolblVE1gjWSciuXCfv77KAvgodk4q4defs3cqL9FniuCXM16
JTYL+fji8vw48dplW7uOeE/yvzwJIsN0svk+ZiXtRQf0sURnz/i5TEDy4V+k3ARnvLZmvXIv2LOn
THmzliLy4Mb4Ecx+9K/fQ/5HQ0GH59biyagRIda8k/aSfl+Ojyw6pqp5TSYkuczp9Dp3QDITOKfy
fLckAMvbTDdPYkh9YA2YuOp5htwt05voFqNollHC56gjhWydL7Fr8bo9edUrdXy+FoFvcB4U6oeJ
No5L5+n9IzA4UTcESeKY7dXbMDR/QCpGMO6RZ+4ejxSKfHH1jDKjdqytd+Y7970Ih9aYPUW86qsp
aJAK0V0ScpiKrEp8KH/bLlKWNHB7N0yfaGOuGgpM9HO0CzvUC3CFlGBizlJ7xxO343h3c36Vxa/y
VAr4vag2T6Bo5fTdL/EPY0PP6vrjyiV9FxJSayIKZRsoyBonYAMhHl3zjU+2HkfHkWxkDT+6j6yd
xYFJLgFaLsYkKqIGOgVDH2dojLJW8Glma6L3uvGh8mxrFwem5MhCkGRQmkIYqL047gOK904HOeiO
G8YPfIej57GdT28+SWtsITx2dRHC7ftOXQ3X6eJO2Zchxk6vQr00BnZVqApSKLfz+zd4aPlQ2Bm/
QsQpdRIv3opc0kthR3CHH5G0nU2aFZYGq5bahMTW+O+wZ/nhfrNOg1fTy0Ep/qyHPikPVPb+5dle
d8cInCYH8u6boJgO0lA48MuHWDug35qOPn5i2CPy7L1m5FeKUYP/ywEPVFuHPXUah+FTdChqRr+L
s1y3+MHZNEst1VL174a8h+JvNqJKRfECwUhG4fOnJM4BjxOyXLPN6sCNSuKRDmORpIhqI2ScHnjG
TVwtdCJHDu6mgCEPh+vzKrseCLpkNoMYHd3SJI4JbfmibGMVwKYL52pnw8QaK0N6M+RtumhqfmnS
uYlFgQXYOqqB+ty6Tl3pXa62XrKzyUsLLjwlO/4Wof7M/4GLqc5oaVByMt3B9ja7+vOGr31+isPD
YLg3v1v8e9EH1k4pWtz3UhFOM0WXPODKJEhQcggFsNWM41NPSOyCwZAUJWKneVfV3oZ9/TwMM+Ro
UoE2lOlJTN/S/E/AT7pgKGZB7ghkhIidUj5wCfYMBiu67hv18e8TS1v/9ER2sn0+1k56IZGNBex4
fYSfn499F8ing+pwKTXLat1AY5Adge0G3ocMGJcwOEJYSFR+1rljhN0Ip12mo01P7q5nH72TsZKd
3wFhS8HjSi47x0TkaS6nFhH7u64/E96lwmFF6mYC1GbSpvVOglYfArGBlxuqvD2W2aLkkZ3Zs9RZ
AtrhfVcd+2O6xYkd2INMdtaBii8zkSZYZ5ozhGfF1R58yrDl/BvO3S5ibVKomO8uyE5gWyBscE2u
0booGac6XxfwbHYy3S509HHeu98Kfnsx3EFy9f9OPgn00CEV/YUa/7I9ev7e5lvlyarRaeCvmYjc
EUucTQmYciNW+nQ7d16eqwaZs3bhBB6SfDXfG2zQ2yUkFyUmZTBmha2x+fcKEIt8wZ9nL6FL9Rg0
u5eLEJHLvxgtnbn81S7L1lzGru8gMwzGgcvY8qABJYXjnb/bLF+OBSpx6gxrrbOpKadbZJfSGQk2
uVeXkJodCUzYmrqoz9e4rEX32ASz38lIfcF+iAnMavcGStiyoRTmz/bwTtF6lTHpyOlNiPzyWbp7
Y1YM7y57Rp0iJu3Jnza0hWeyWkULMtnqTkYzTaauIb/p3fSAkJ+5E1WV1NJjL2agQsaZM5FR6k4u
LQAj9lgiCPOUEYf/OVGtKhN9ekw4kUPKXLAKNndclmNzZC6yNYZqFWuZLCQBkA80YsCZD1x8Bf0A
P/NFOzTJJiRkatMxo3OSBMm/5zj7fK3OvDg+tEkdL8Cmz7UImPd7NeYk+SDuHSp4ZhA0KeRu2pUZ
c1sdS5zywkDDf1Qdvb+BPbccZCkNMCG/NaFbiOxOk2t/3pp+k2YLP9u38ZGe4EYxV5GNkbZxzQiT
fBNmBdAlMx9IpBIxzwCHHIIj0jGOi9SnJcJ32+OqinSD8SXbZBzTdga9NIBTn89LOWl3J5v+8o1R
yVWE4uVYmFK9r9IxoysFOsHKAmk1nqszoeCIvs/00nbUwbQhj2pZcR4FnmHe//Jkx0ietI23uFBy
ejJa8Pvro+WEN+EYqxxJDNGs3NDbzNk8B5sGZr6LHNKB4jAPE/vf6BouriveoiYJrPdbj4eka1/1
4hiye7xSXxJy+7Hl2fs47U/QqYiN8JC+JgI32fDEfwdyuVnmhyYo2Wmep9uRS7uoiUiQavv8yUPt
xsHFwYl0XV1AzI0cnWQ1MKxhpUXj6/xe12hFAF1IaglVJZowt6snHT51bGC/FWtjNSzfPPI6Wx/k
S8Y2q8u5ALRYqyiiXNmw7L1OCGW9Z4FzMlWnMlfJG1TEqvhsOiKPivxhphenG+LhpJyC4Rb842eD
Sm/46dIn+Ytk41mvsifPgLeZUzulWBaT24WvvvJIBSqQZPaBHF3znZ7hZmPiLabcojc60SPNIsHC
pO7XJvwc8+IxXISXzrSYNbEqRswUQk9fmJHIUpc2OYGwJdU2aF4GiyAGzMftDUwIS/ByrHug0t0E
ST0MdLZxbgcfgRkx+iDCbwlMn8cNnzVssPhOgz0rMaO1ie6RXDmC4vDBNFH3GHa2MCBpOBFAA1kf
+Be+hXRoXq1zQdhbGIgV+L7yyFFU/dY0+MCxfltSQEuNqWGZKNLa3561/mR617QdMsFdb9qAwZ1F
gkoF1QmDWL2p0mb7PHAbHL8ufhM1fJRs8lG0LUOzRq3/ynI5sLLzD/LTP0mT2aW8bFtROLAL0nRo
EWKwnHGoPNwNwPTOQ31tW+HTOjzULIEpNfLHJtktf8qV89SdmlYfu7gvBoQwZLrpNT6pBECQ4GkR
VBHSqw/b7kP9FYWjCtPIithVSJ4cfSO0jfv0h6PAvLQmONw1Alyr0DbghVmlpO9J753/aEFO3d17
eKBHPLQXURFFwq46I7TQuohZ4+ArxH7vkCfQ6Pd+7+3CuWmvhbKHiQ2fUtt1jgMaLZKFP+E/NAjQ
UJlNlgw9byN0fqUOqV1MFDj5K9hyysD+Z7NtsUCXYmzEdy6NQdJfiGy3Z+PIlEuYIoPcgq4ksNiO
gDa8b+2fHgbjv06+Di9Bsm8OUsTO/c1NyiF5algNK8svjbhl9P75CHDg+tuEcfl1oMkeNk2HChfn
SG6x0R7mpqGHrxNlhTMV62XpK3fDdQO2Z++QIOcFw6SD+FBLfmag6QgE6wD1ZTh/skwn4Mp9i6z8
RN4HXL6UXa7cZEgMP4tT8cloO4JlaSq76FFEOuYhPK9cWXmwU0fDbL2ZbiDQEnhWzQMAdLOhIQ3j
3PiW/yp+sVUNyMwYgcoIjCPdAiSi9kiug1GshdU2gZ8tXKU50EBrwXNjC6sEJVNcUDXzNz1jZhJ8
9eO1oD7DJZxzreIY6o2JR9nYvhiPVAL2311iygoW9106X3xL0IkhthZkimNIEqE19WDij/QOdkEm
0HX2024kydlJ1JrBo/b4LWNSGAXTj4hEIhOwu9Pv7l+tCbmukq5B16G09gL9Ei0TH8qZiR1jla5S
jCB0FLcuc1NW/umnfq/S8mua2miQ7gEscv8/f5HRlMRF+VfskX46Dhw9p7b2DM4/AwcFaVfYLz0X
LS44LUjOrf2r0BQQb4wGiglONpmT5pKgZGICsZnHA4GVPWFh6ojn+aU8/fxE2/l+V51tWw4JpFAP
VWdR4mWS6dT8G80NV5erVRnmj+5IDLfVILa6DEXUQZ8K25mc5Dmc9afrTjJ8B2Xeca21tFpBOmK7
XyqxWuIPJ3r6O/JI3rbwO0a+vs57kZbc5910kvnOTccNmSq4/QZe4UMzeRU+2XzQMrep8quDFjSa
xoxjudviFz12ZEUAVvi7ZYMD1bttRWwtI1WNK7GXgZ7yAEgFkcbdElzu92MYllOwyA0vvsPsPPcF
KV22jv71PNGW5nfgrFP5BsKafy6/kSsox0bVlQLSXak3dNQWSsbfi8000CIJVdxvK0yKXpEf9df7
BZ/NXZqNBKWpHVvAdbyvERiN7ZjRAjnSPo4PWxepmdxpS4A+e6cu/mrYF3SFI7qaSwjvsqjWOpO6
R3efGrU1un/SyluD9xlOfLjvxnB00hoD203mM8TgaNjwx1R24j/AOBASYr/25h6jOcp78INQYI7j
258G/v2uLurwszcLvZIvhjNUEA8iQUiu2IL4sWfa9wCX3QFZcN0k48QV02+zQWXFKkZzXCWZjBh1
pBI2kHyx/dgRWuS8VRvjN7uBP1jpUA2H1sqaqwVGaWBU+MIvxdUnj8ck6VRo6apbbIpYzWCEkPOW
+Pdd8aX9FJF48tQn1jBz3BM5NFHhmFocXSBBary+fq74zoi4PcUOFPQIM4Pdm70giOK34nxUaqb8
z62Hy9MAoD3qtacPx3MRCs8Jv4cpj/LjfYkMBDpLRkKpeSoWVIv33oRFQWoSrIg7njbtCto22iD2
a8YwJ/U1sLVsLAbkrDImg7aLB2TEuIo6WkycENzL2wUpnz2Nq/N1J/UKKHKZnoeeAo9IW+kPZN8j
Chm4l6TgYnraXxNYf7Fh4ZaEIHDqlU8tu4N8m7PGnZkzrYfvQpUsDbOZGamDL2YHevjNmKUWtgaz
e7fQAaf6972cO+Ym30lxUfUrHQ9oITrjetrXLo5jbkcKIEzigRxLUlAHB1MJ7Uli2VBR6z1iwbTv
aDZ8plCKfVh77D5uAHoSIkqvhiWx/Tl2aacKjPGFFCzLYT5+oSzC4/rpJhAnP+lQbrLODaAnbfuD
drtNHVY9YMPN5gr3bV2CfAuf2J12dKH78KLqRDJXSShT4FV4USN3+9wXi95fy4uJGCC9Vw0j73S0
WsUHJg/0BLIy148CXR16gdkR9XvAL2fK4gbIcDDKWuU+Ad6nxRjVMy5d9HKAloiacRnLu72X6fsN
sv3ZQ4bnRsAMNsk2c20AbUWhXF4j1G03d+szm45rs0g/aWiPIXwD5/0eekL2URKaMlIilFtt6hnQ
V1aObK+83r9rvuuuURw2JfGLM6c+4pcYmL7M1ZD8mAQawRU0rVI4WO/P8vvVnkBjzh2z1mAwSnk1
d0V8ZrdjK7+ggDUli00WFvrHRcASYl2UarYPfT+FbHI7LnPngB5vtkagelbYXaZIANVcxco5WXvw
b8JkaLc71S6yd1awfm6iXxo+ATNwPiwejyHpwDV21lNqGOXcNZZEMLtB9nm6VtgcpHwUY+8YPZXY
nrTxSHf4tV4pkapL5qwmnR6+CfEX08Wlh6eqrgQ3enBHkGGCK9Sq3eMURUpjC2wCfef2G/uBZRNH
DkRv5B0fA5eFxqH5QlN/q3m9kNG60wW5y5ULUX7BGK/Gt2IydVhJObC5Q6hoq4NFGrYqkBTks9hR
0gOxc6/1OkKPd68BZMQeHwDuUFkZsVrnMU+Yo3+CdKVzKX0OQVVHMx3AFYzU/DOgOmf6PM7yw8nV
AdF1nOKdz+nKr+LKElKBVYQgx98Oh3nvPVrSCf8wlQ55XTHkfdfhDM/SEedIXfWipaQt/dAWTgJF
OBwC0caizpZpbVSxKNWZyfFzJfxRnSfsyb856gdKmd22XLxN7CR02/dWxgCwXoqQK7SkUl+paYv6
1LSI4YDLlKd841CJqLktvynzZEDrJGTYJMXPHeKYyL/VcVHmTAGM7mHqaJn693M1HL0in5lIreY0
KJxrODs5Fhr5RyG5NLEQksbeAGC0+nCdyX1pTvoNht6cuympX82nxk6aZ43ZNySaqwz5opRfmVgS
6PsSSBlSQ2h7u+sPmdUOVoseTBH46v3hFMic+rIerwHU8gIqWPNGNVbZSwD0vafGKvhp/7jP25t0
1eV6D/TLkEyM36gDsy1wgGYjxjgcpCm5a+ksfRsVPuL0u9BA1rOH99ntfWpMfFz5opGctAIozFXi
uKx0W3BPccXAN3HTkKyd4wKAVAWSBtN8Cui+6ULd/nLxB5zATZk/ZxNO3KiN+eJSesS3xq18NXk3
9aXq2lX/nWg4E9oAPzoFDLyiBZ9Ir/+t1Vc8+BKusuHPfQEoLLgI4hoow2Y0Wd9DLpj/KDjPafBt
vcXisCD7JOsS4LY4ATi2KVo95YXlFY15bEFdf9O/+eXdkccfdDzG3Y3xTTvyOHNmuYdTggtr9jwE
qNHtnJlMh9q9ly/94EDzBAschtK65AHvUdJE3DwzFFr4w1vEHUUYAKTPQuHs9Kvt7umbnWWKzTJ2
T6rMgpb1wbJHODP4rnwtetWj9d8KftH9SBZbV73Gbn3WnGLgp754DpLcpeXXcE6O8/qbX84mR/My
jstWWgJ+aCbSPil6LFvmawSg6zAM+9TdzMgNEbIU1sv9YRwSlmbD5HBb4Tw/v6dJnoN+ugmX4En8
+kmMtYt/36EULQaaRoJVYS4aI4LPhCH0cgCi4tHrNuF+zgC55gNVB5sGmVYyXkpzStZcvQt+d40z
n5+FxhXkTzG1Rkq7lKfh66UuM69Y8Wb9+rQyydp9ZvlflOUScyHWiIMg/Kxg/cSEL9tNfbowTHTg
7nwnh5De2cKUFRDwSdWYijTDwY9qaRdP0e1N44xQVqlXOHABR5EQ6lK13t9IzaG9ZGyXbdZdMAUb
u0pJMnxV3agwfX41/J8/OacdBdTXuM7H0S/b3CRuDxfxclbGq17E1oLrySJn6PRiKxehFFT8xebK
LyHmsad10y5X8/VXxywnDG0g0SXnHMD4PNRYi4p04amQ1m+fgDtAmgJk+xROwkkNtyo5oTjJergV
SS22AfOIxeM+AbDG50FZeNZZ6DlDAjBNEPZDKnAU9PGC3EjO5sYlvAf+P3rAh2vHw4ORFFEQXbsJ
l/K6UiGmX8lNFB69UAcfV6si3YsvTh1fsobLsbCJ5CmgRgwlA32i95sIWxA6HiOH5JBj4XdZb6Sz
kLfpDlMk1flcm3aT7iEPbUdA9PiJ9YfcfEyj+fmiJOKgj9P1m2Woo+6AsxQPF4ChfuQybFTme4NJ
fNaQjYBcl1vu53tQ1NWqIkac+VhwzdP5Iuws0dyLaKVfai1qGGpGWZeYC0urQ1VncL+mFT9zSaff
bgh61FvkbQYzazbPA0iJuixgUHECN1H/VuyUvHv6qzpF0w6vnJ7NRhpiJ+I8t8FW3xKwsRAv8J75
pl9VmMq4ZFHSXnbBFs5a6NXWtNmV+4qSWfTFZ0TFoeSateuEQKj1Mz156OcNxuOtQDzFSPPAMf7k
2MPrUebHYGYSRYt9IrbxFeExB8A2aEq4Jf+yOwBeS9faztkb93GJaxqGEL9YOvM5aZN1g1YO0XtY
2ZZo6pxcE3Ae/ccyNjTlUpm9+4MvoIeAM9bIUpfwIj4CqVIZK91c5nx4M/JtBlnxg9zRJxVEOy+A
wAQI1ObAkyjoMF7BaV/NDTYZJGUw2OtlWSNPffZkBIZch780huYwHwg7b5fyguDN/QDUPaTUtaGs
V8ybb3/m20EGHSnv1Jh78J//DhuRb0jXsuHQTiT8pmYSnc2Aq1aPwIhR8w2bZgiE0KTwZi/G1orc
lnZDmr/U8CdUtIHetTWGUU64dF5y4Y32vG/x5+81olM3BeI3W4B5kQwWXLy3RzgXRFQ8O9cguSQT
D+ROVnR7uQGsMaU4jILsqoA/YggmBa8vaZnQoDtMCEGBZLJ5aoVkvDutWWBZirIll/ttA7qA4IqO
h8X8V8oJodCn3MumzZnWe/k/fH5B6z5j+9bnSo3+Jr87YhvYnNcpgnCn9rS4S9X8hIJld664BjhL
2wCWsr5zEkhFtRzBIC+xigpN/R7YeDzqj0uj49vtDkzndclO35McxiMnNfab7v1Rc4VJO+N0MSGc
gwbbzrfsEdl9EtxDP/AC9pQIiimB5Oj61H0Q1i0QXuLV+KykZqXbckYJG7xImLHj0lj8fa0JCXRZ
/iZc3MFc7VkdsEbNEjYDvvLb0VNFnK4/8unbzMyfPNcIbQoty1xM/cHxaPxFI1yHCzd3/Snvpg4H
5V+cWhkbd2FFYssTgTM+vo8yO1tunRsKXO/AD0JIF56RvXETGdYf/3z214oOG9y8LbN2rKdbudnX
4NOr+7s3YFvT4GzancV5xGXvaq6R0ObZ/f20IIp/G3MH6aB84SiDxPAhGAks9zMCKCx/V0Kvc40a
WnRcGuVm9k8Usifb6Bk9Aw+TTOSyyx4LsGFJGrdGJOP87Wb0CDHBU3upEUMAkp41fmaZoHBjecH8
fwIotJbnaWoP/ii1Mhs8IgaReaZiTfRC1oFbroDzGWfr80Wtfc7qb0Va0O1Pv/dOIHluWVVyuZ4e
isqnv/TV8dyJ5ZVI+M7/fENN+uQk1BYjCGhJfck1nSxcbKIygHsWUhjQw0mMPkeKGzBIrIfIL2rL
IbnSgOEag9CUt/tJbpsezWgRAkvw7GUXhgzc94zeQAucICWRUdRTTLG7yL7tUcemSTxtN1WQStYO
Qpj9aRjQ+c03vqAx2Ab6wTj7JRtaWON63KjR8EjqCGhdjXEHi9l1KwnZPZC4ZOrQUXhgmVdmJDeN
it9RqJ5lMTg79nSRsJ09Ec/lJgGnHUuin2M1PefHR+zbHlZUvlkt35O4lr64OVvmnr6/Ga7ur/tx
imVmKTMiDhY4hx4GI2MHAZiE9vExsZ2n1Uru6DZkEkRvrq21EdEvHJRJvEmnXacLtEd7KxInq81S
OKJKBKTXAGhijzlYdFjYD2lHbbiMm0DZFQwhRdikdeN9Qcx2/9GjRaI7g72VeJR4y5zJ+wM4MXNl
SUtNiGtwzQyUpm78qmvYdPXMpyl+nQ/FLZD8H7aNbbGPOj08x9Sg3+RkPZpXAy4KcRAChX/jSSFd
EKkLi2Dmy2tXiGBDSh51bYUsqcxTFRxqM914Tcjle9dExYweKmhxX8GQFBkkazWYDZCGpYZv+Owd
zJaPGRh+VWCmreIn1wAEivTFvwchTe1bEg57WOhbjcocqoBcH2lGuY8GN1zPv52bjbAEDdNteB4M
IMLpSYbdWHF2VAKvOu9WeKw/HNOOaj2BWpfEBIYjzQxaDj/SpF5cvA7iCkVEXm1lTQK1wCVAm5oz
yrE3GQD1iyVx3tyPugcc4t/b4EVd7lVR5SFeh4/PF3JWgn6TKZIcA1/JkurpiDqZp2GBh09awMZr
4M8xcqL8uHEzyrAPEQ5imjAPasTOHso1rMoKIui2Z42H6WCXgHyJmddivnndpPobvaTUlAqw8PRw
mP3l1+y2TVUohPxsCRx3oaO/VKIRd9L40g2vV8eb3KbvvpeVxFaBpFQcZCQOQFX8shzXNQDmzSmM
3tWE+/VOUhCgJNzsKV8KXM/6LBTugVTyUP2/3OOLySp0htkwyAcwb/Evu7Sln4ZfIJ2MYeX9Y1i1
QpnOBjNeD84EzeHciw1Z1BuO0oWDt/ARZ8t/oadDxiiwDzpwuKjwco6pBErlzAC/QC/se6juiw1F
C9i2AlinB0waAUgCB1p1hFxNHhTGYRqVvOpLsnprA2tSU1Maw4C/aGaDmsm7Za8eSPQAxJ9tsLfy
BEy+3aCVco2TdhqZcC5y0fJE8AxyoQfkze59s8r4F7fG0F1RH5m3ISTXr83fMI26frybBxNRHlyo
8Z76rBeoQ/PryKG67xQfndb6z6JX0u1tJT50gE5+ZYhl1cpF4X8p7MtcUvtRZKB4McvM/5y4dcE2
/XHVAbE5KxNguJRGEpTjlXVKKT90pljv+LCt9giuyBu80eWksNNSF/ua4PcXzGOQD6XhOuCIol9l
ewMvb3FxI4U7Wm2nXgbkLayhYi4lX63YW4m7M587Ydv/3oyZXfpUbSGZTYz6e/NxurfTJHrc7YlC
nfFguzpIR1W2pRFNhN03GHV4xMEXaAe8WO/M/mTvohtc7PB5z9jL3MR6RZjT/zfTHWuhQ9vx7AXh
Q1EFK/hQMBWxFbQ3dat42Kdd/qe/GzzyeyzdVgwv2DQd/LmTPw1O9xo0JA4+zrjvON5rNlbC0PHY
CkwR496R24PFBZ3jsAO/pa58xnSgfUsZf4cePAz+hiPgolFxbAc3EyZMQOTrldiNzVbVX8410cX2
LucWqEJz+jj0cl5Qx6sC9P5SimOgK+O4uurP7OIKXEW2CBf2KS32/zAhLMvo+t/1jYmndReBfHKD
wXRLVWarq8p/KOjCiCBiFCTX0dVdVQuwEYCVPz2g1MQy4ObHh+mvsuIr/KBMOR4Oq9XbzsSDU2mf
O0nEhwTYYN3gbGlabD6w+b6M4muRz6uAWqXFkypW4NSZP8XHUNX2Ci0JexeWcGaI1YVP215AJ8Pt
D2Nlz8SERQ78sAJYdLgTotSmT6jWbLUSjLHo/Us32vbWv4jilUQHh+8DlqBh+7FNUqRcCQNZ1Me7
P+HdvYQ6dYFkXkhALfe9rS7yDLdgFGINu8ajJX1JsXBw9nHkOgdk0+nnnl8AxAWCssIAR9p5ob84
Aph2lHvSVySPKac0e1ohVKcu9aHXQbnfYHnBPqP766M+5cFFHelcT3ShWimgVQ6PqO2Gr4xlyV+P
qyy8AvIiKS2mvL+97ds1spa2MSrBKmhJFZ+jNHc2KzCqNCGeP2gjqeMxscZjJ+pVMUZr92yYQaXj
eQ8xafjTk05Obp2KmkaOC0TXEhLSxtajR+0y6bQGDLQI7AbYg4QUMfWjq5kk7ZkwRZ7cNuJJUBhU
LY21tVmVWkkfe+0f+GG3SL3uZqBtgHu3DM0YtxtXp6L0sCEack4WZWR3cF7fx34WyrZsKOO61Xw8
NzCZ1cZMEpnCtfVlha5tA8IhM6RwyfVlxzkvRkzZQ/5V+ApR1KSnttQRJkTRpJTZoGLFDARjnxZw
ixI8VTSxafaX/XKSnFnBfcWCVeCOwoj+vRAZ1s4RpLARjZ09ajAAK4oeR9JdzUz8Uwj7Xg3SH2+4
Q3G5YzBJ5agossNhABznujuqfc3SdDugLwbsq1Yog8uqKvTuwuhvcy8rZ8TC0Ozg8V5eW+zdOd1p
OVdpeHhIBTV/VcH6X9B/eg4uu76ZtIqMTqEdEKkNdKU0DoVW5xWdV64Th6jEyXgXBswoQ8gdh+Ap
1RdW+bFh2q3tunRwhVKfQPX/6PWv61nh2t3jsW+A0LMu19R9IqV01l9k0x0tiHbPXRiXfxu2C6ff
1Vx329hGfYxuthAr3QtBYKbVoJtNnsrEqhW7AscyHB4bDPkCFPgC2GxRD2b2pxDv4K9pDHVnRHht
fIIOHP5A1oegRpSkbHn4xiN/ZAlRzinw2LL0McbdI9dyqFcYRZ3spHCCdFR/B5tB0Dk0v2CNgu/8
52o+XbvwYxH+IK4QaAGT0TILBezsnbomM2T6nmfGs9cKPuOBjRnGD+hNQ9kHH7awLQKmOo9L9fvs
7wz8E4a9/fx1fnceVI6RKlmYrgEriuR+yVCrvTZR47XLN8tleHrNdSkvCQ+capvSS43xm12/d2js
lNSa9ePshYCfqfgykraCzGD3B187vq1t3Z2WshZ5JMp+ve917J2FTzqNkiSgNxGf6xlYDQXEaKDO
gVW4LucvqTYzRoY6vNF9GOscdbHWkWmAefDO5XysXal+QLVfJx4lR7mZpqiEwgXUy7A2SxYlRvAU
K4NXwT/4fKRk5JWvAbBPE09vpQam6HK+kTz4JvYA96TYq3KRcJNLsaAEcQSMrPKNMVffMertzdu+
2VTzPEm03VXpTbqV9/jXlbt7lBqWSr4DIZe1S3fmLr6ujasg+ZQOJdu56OGmSeOjwrFiKqXT+Jpf
9PHYC4oqpLybIfM47P3CAobhPyQluxeSqFCKtN41PUvNknw2+FK/bGj6HfWwZcmGB+rOv7mj9Dc8
leJGW2stnIJY/IxAGVjywTBVqehsEUrOWXaBE+KnEG66zBfPAPmtqIGKlguycQNx6D0mnjVmToz1
K+anVF51KcB732l1cRzk7365wOQFG0weXzbJ6BnvHduX7oNrl+m9IeSW1+nHb2l7HxV/nv8oFh5T
mAZJ+TOp83FrDg3sM+DrLUu9AWi+W6IeOBpnW1L3PhoCwzXiGdA+2gFz0lJwp+aGktlDZEboxUG3
5tDgCvDktc76dvvQkFaWo1gcllil82+Ze+l+SlkenSZpDo95+X9FmZ5wzQZfq7M2v/0zey23UOjx
1dR0Mt1vsbbG+pFUu0P0PULUw60yvysJwmW3sNAmsaPq+rlQPzEI6nRc0nxznGthUGBk3HcOToBr
1r7hfhEIc+sxcvxfPajv7Hnh/acwIcftGKR0TYnln1FT5m3qB8Ywhjn3IMY3LsN7JIjIQZIXKVOR
eWHMz8KSWmANy2vCgALh6KvodDJW4gmsI4/GWSwIzLV+QqMyovk3I78JHo+w8jtHv2UL2ImLeAqo
MCMsSJI4Ta4lFYrw+Hasl06vPhxmI6ProSwfdR4vcoPlerMyhCDyZWzICpuSsprKm8oTd/nLO9+J
/nDkHMFeSRogV2OQaMyEYtK+Exg1zV9xp3kVecisyCM+U6pYEQ0lGGadvqCxS2sp/kFaOg7Kz/gv
1BC2QeXEBDnQElX44kD7P7V3+YnilGpe4x1Znn2HS6nXloC++1GMMYDKMffNXI0Ezh+5v+32cHB1
NdyZPkD5+uxTqavVNJ/BDOof+YY/CBurlZuVtFiBUdX9hMG/Ret2KV/DYkDlKlcyf5jpu9m1JjWx
K6oU2mEzlZhCnjavb8gANwqnxtFP5jDd1jtSaUfXLGSaHVNSNeF2KZA9Iwks9/mV8PFinIg9OZcY
lhy/O3iFXuCRPiTfNnNbhnc4XdO4bkbRWoPbSaUnkKJh1hRDjJ2TO3Sur0DoxTzfH14LNLjjLIGr
31iMIjP4uDjgGsq9rD+UqQc/qi3n8E1X+EBaSGLrNYNdta3ZehxeE4uZkO2Z846KwMjiRw4yo6j5
jwSH4h3ockdTFDWL7kIQRPIqFMEzSJEK+8SF6RnkOfrhbXXDPdFNqWQpM8Y+PhFE2X4SXMyFCnUB
2mEE8L3yel5glozLZM1Nb63R2kMeej9wy2EKnC5LAsk4luU049SKmnLnf1uHvqGcdTuhiVF0w8iX
Ftmwb+Ha021sk9LAZG9hBtCkdRnXpf5cZJzYd7Okxozbrl5mX3B4g2FMBvRrU/fPoMaGhiXbM4rJ
P/qS8vDKN9iYU08/VZWTyBFhp2lW2X0ZhoQECH0g1PPi1QCYDTRq/iEvKRWjdT5lpeLjy4JdZBCD
/wrxOoI3ua+ZTAACULKGd3/P5axc5lFoIlQFic6ndOZhSt2Gh8+NyNHBZOPa5ljHqUfQZHSdZb8j
ZjBhjD4d0Ox9pEIWD0PRyjdoh552hcziaaHivRRYBMY+CA/5X5E7eQLRy2xRqUHMGm6ErI/4byLO
XQssVwR2cxudPFkxhN0t1MalGNpuOU/oyARAYBUzPPeofKDcGfUlYoWuWlH4MbsqAoiOaI3YIoXI
bwP6QJBSCqgg9YqLEkrPBmVVAO08pMKBUBO/bXHn+1+Arymn87txoIX5K4qGdzUB3kZ7uLXSFPaI
pouM4/7W/90NV0vzHs2J5r2guNFZumFwiivNfentdWWrw1zkNLwWv0xfD6ktaTa3GzeAMLLNOzVt
YaJ9UOeS/+ZfdZHbUeb40YPTjSm8dvn4k75aHc9qZbpIAT8/JUSd2YmVddyixVcJ3XjYEhGdSg5h
6yeAV2iI3v/h+GS1G9XE8OHQGud1vMgS117TyVB284BRWhJk5mC7Brr1Y2PUOlDsmE+crWuQUfLM
RYBGtxU5AWSKDcVlAK5hSV79+CiuS2yG2yrzyD32vMs50jJ9qsmpv7lemeETBHqA9k3g3ELtMp6b
RLcZEPtirBnVKevPiMpTgnNc1OYnjJqt4tcXYue6FmkP1qtlHzvKD3rrx4w4B0UnT2pMPuz1SlJC
CQlyZ42Sy+g68x/Igqt7ntkQj9aGsCwjGhn6gDs2qVtq6tibhTByGSJt3h/d6DU7oZzmOg//GJB+
cFUiYXcxgPw/7EQgjgXZeVCTdgxdkhNX1GX/227rUCKwaen1rhrmQSyo2dkOj8jKTaE/Ccvv5plI
C0VuNllkm945WqODwbLNc354O2+rioMUb30VjUh3mrrQb1YLLX/C1ze4b51kTcw/gg1Jd1IJMQGq
L/Jb1+j17y6yS4uy9md3xbwkOajadRuC2VlKO4FBw+7nloHmdT1Uwc8JqOaYwG65Hd6IAPphGlhF
iOuITEhyhpL4Sxiq/zBHTNzKBGeiJPIloQ3ihUnL+rQD5fwydYZSC7PEUpRz9j008nzTyUaYDfYJ
ph1kBoGGl3aVZ9qAclSMRkwtUjYUlR+JQztXtSa+0z8sjE1qXpY+xWOK5DUYXU5q9lnOQLGDShRr
0Tu0MQ6/z1P2NcyTLxvpiT4D0AN61cN5NtYG03sEUWJ+zhyMq/CiEqXQyrDv9dbz4vG5Dj+OW93B
/CwcFhXxGTrNpEqvzvO/0gDM3oTFx7CsT9cPiMUmin83Th8KXUUgO1fehl+eZvurEppcGnZUlgaa
kvSKvb9dKQC+ZaMTQdHtj7N2FmfJygRveiQpAWIgs+Jj/sDLFqLCyt5U6QMw1nmHk+wjrEGw8QZG
BsAcTPh/lwd1Fmmo0s1FX6P1S/6N8m70XCubbF8lts/vQjZFChGAC7HkMKiCGUkoQLUzuCJMwDU+
1Zl/zKEOGhbkigEYfLHZG+rJPCs5ZrP/m3HFuqAV5ttz3yQawxpArGjFoCWv8zPXT22OFWgAd3nI
+2huNqyLEzIR8jqG3mgrxuAWwIt6JzyiR5CxmLzitvYvQXFJMVWXWWnhtAZcBD4Ci+K0Uzp8PDKc
Zr3StWV8BdkSPObWZVY6qy82oNIsx9y9jIeXh+sSwnlI2yC88fCSZUedUO319EpvnqUb6F3Yu6yg
7TDs1QWwiv3GDNu0TdsNRv93RAM4GHtCTmqMoG5GApXSQjbY6PpEDfO+ZZ+/JVka/N2ZtSLLXmEk
XIvtNHkqQAO0aXRlSnZIIgmYW7P8YMaBlQx5diC0qAeQJzyj9BAMQ7nNp/MJKuAh0iHVVPirgLcy
3WfmotIfE5Ld/Q7NpcGAbKn7cw6T84fO27WP+GBvyiSMITFWBhqp40tHf75dvRT8EhiSUFubsOmE
Yb69tsrelUIE7STFLGnmhE/0cs9rImy3aFGWaUmgtub8Li7vdD4MQXgy9KhCJ+OTEUUMNtoU3tiI
ofDe8l0qZDemGL/OAkGwUE1pq+hYz3q1zzn868xKHX3I96FHd9So0kzcwdBIz/7QxFOHHA01oN0z
+ECNE1F+pKXv9Vl9pYRVwbyoe64y34y9rs3AEAtDCbMhVmERvRC5w/bEUWuNk/SxTAq2usGfnL5b
kx9f80OJolwQSCysKXTuqF3lPRJlcHvSbKUBWmVg1bI+yziZh/NRzYbjXkJZb6IX3826D3s98Sjq
nmfNmMHK40aGezgFaQ8cRbg5IoX+LTghR/ve8JgN/e3lzbAfFB4NdTAWNsvFqPxPXbO35nNdM3B3
AZwYAi7U+njZgUPeHifVasZ4Rtg3s5CY4HWKcloB8LMvELjLxfW/ooQP/C/d6QGY0ajzu15zNKI6
ciEvmFGxN10ZEQTg23uBRASK6k494zWt5v4iUweTwlIyXQcXygCkApGHaT7c3Cos3Zx0cA2/FDsb
p8yib4Mr57QghQspolg7Fci+ugZyKnZQzGlqS/xT8d7oqepNufeQtW6qLbHidaYQHyyj4neL3aUX
wiTQkwGdSOT/13aaiw+zvolt3loIA1vT1M4XQzfnlMCKUBuoNJ2GL55rdM44lAESpoe8jtsZfRoU
dLO76mDyDoCk7loaIBlFdw0hViFAloPnvIx9VGVReBjYa3u9eWN5k9+tuOMspcOH1UNI68dc0gWf
KGWkQOoONYhcOB+6AyUGO8OvhEHNaB+y0xfW+dcss+l0So4Ga0NU6wYakiQvQbpD4bQr7CJuSH9c
9v1X45/SwBW8QEoADaFqxifYkrWZLK4DVlEWug1p9ObiMCo+hzYXVqRKcPbES8PNLjqXREd3hNl8
+vlN9XNapw3/sru846S6YkOpO1f7i1IYZP0rrokDni9l8vTKWuDvB+J0THP3Paur1rWDvQFILEIl
UIUwsQ12sgr5E7MhYx0hvUVDON2jtIho4or2ExNFEGU79Efbt4NqfsbYVY1oeaBwwc40XhzXuhjL
eCSC9erU7nGZqQE8VEVQTt8nTATDk4N4WuQPNNZ0Cv3PW6LOkyTMq7EGCBZA1nXXOcRsRhZn1kwV
vkKlMV3UYFjqCFzuMemH9QIZLChLTDulHax8pPMHpaXZuwM3hxWgIYwBquU/U1Y5C8vL9JPYHv/+
jSYGGIzPqjmlCUPhk5dootfQkurFo0gAJuxvu/qd563/vKUadfvnHoga2Mf7yr1GD8EJYv7PTJUv
qoxfSAvqLINTEf1aXGkey2vFYhlC9auiXOD9YvWarZz88yLoL93OgIBLQaz9dqFh4f5LojQqCKEC
tMjPfOzI0Jx8mJ1EPOd5FXVAa2gJXXQeMCtkH9GVAE7gQ8ZcurzzikK6FEqz02nLh0FLVs/9jDVF
66pGOEhMXqw+hfKinNaQRhjwy7/uEIRGVTNRcXj+/LtXfUTgRSy9kOCWHnYPatscDwfRqy2/CiKj
+vRc7bM6WleWEAjqYxeZIKthsNymp6cuBPWvlQUqQ+qZUSGDPXGpFK6DuqbFC5CaYNzILh6Nouvo
lYkhapD6125KCiS1ARRr9LCIweHxkjrBUrg5ZbpjlnaSnbUN3nLydt+ZAtZebbk2JwF6lK+nsnTt
hKFYXMEcwmd57nucmvoNvqEiLNa7z56+y3tmKe6pAIrq3rVxuY56Rsw//kFpGmvmGXzZxVfNZRg9
BH2nNDjhUUaSww9tLZVFgsCQ8C85vf4VYWowwzTUfGz/3k1zak48ZNs7Df9B111ZnuVTQQKB66wR
rh1TUfsoyHJPWLqKBCET+Jhaqhw6Kz2ESnfi47M9mG6jCycgOUUXPa1dYkDyRkorm33HF+3kLjFn
PTdxhxFfu3e69629A2FU4BviTdtKpLyxsvu1OpUL1RKUzHyV8+mhpNUlUYKKjNgboAIHxZdiOV2T
FLQ/qR3W1wGwQM/y+XHZ4HuraXYaz4EzxoCvQAX/+CzhhrFqJ1qpXOpEDDn+Mm8c9vesHhVz84v2
XK3b/rioB3YPZ/8G4qWjP4OODbOOGVPoX55iZgjsT5yVxSw7dQ+5Jlii6hAcVn2pQPcFAV+Kfjrx
iuSxjyuX7ts21Kv55ESMx+slquXhzPnuVR9XHoqnHgCNc+MH/CTSUXKupYUtzH9/jXrDPPh4gOXX
rwReGcvC374ekG5xxK0/4e9wQH5uAKMm3osDcJuJ/FQSR4dd69hUB3romzJH4jnAw+pcuVwBf9lG
yfx5/6eIM8AC9//CT4Y1sNHYGPHpQqjzjYrgemEcfKGiq5ARqE5N2kUSn1CpAnHzeC624oHXPU+5
QCvuPoM00XqucEoCW2yZkCzdLZhey9RfnkYXnKJLjg6c7/5VUNy2CAvI9mdZ/Hc0fyAt2x/z1NIq
+R2MhKikUSZOzHEelUvUwbdn2U5uAEWvwGB88r8LOkuV2gH/rSzdCRJ3GSOXmeFro1MeGINJfMYI
uuEsFafcRkyJy8P9bOle2jDieBqIFEBZVdY75ktBc5MpFkEWdpqpnVHvFXeg5l9+1I7ExsxiMraV
/Dqd5pL6k4ikXEIm7NmUv+lQw68wCKUXmi1h0h0mNRgaYKd2S0CIPI5ZgLSLpNx2+yZDG4p3dlSb
lsNvmt9721AFArIWULXGUWO6k+hXmyaY1uEO4ht23Y5XocoHMLoQ45adMNEBNj3Av+BeIFREGeKK
ik38aroZCIufdGIkIunlC3HfQHjeFeVe+AH6i4xAlhsBc6Ng2mrTkYlN1/JVnbFe6l52AJ86Jjey
ymLIybDl8IU0Toxf5MChI4JHsdd/Cu93geVvoprF5djL+rig+c2sOMYszASZ6iNshiZgQwBcWLrQ
ffQxtf2eJt5I464/03OEZ5Dgl+9hujtU6KC5hitg7ot9CT3U0TcQd6tbHxB15taJ4BIxqJZmkj9m
ypGLwog6bLW/T3TULl5AiubSN0kHaqARdawBa9Nb4zro0T1bAQ1m89/YrHF+vRJE8GxXffogQ5pz
YVUOpDRVtSkAe5nLaME3YhvqQxdhYxRA3PYVtrcstBEP7iNTzN8t/OTIiyoNJtLBPnsyz0J/Rv1m
Ptn/YOAezbdfGTSR1SZoh6mCAsO+XSQqgkj8izGvP2RHrlOZiNJ3I4aJr/FkYqM4tgxPtnblKryL
4BY10clKyPsAoQ06RXuLGhlaRKT0YjpEEAzOcGRgScf5CsSYwdfNnRNVdSDoCHr9uDQR1EqKyFrE
DySBwY38Ra3fkbnri6TX6IIedIHi3q/5Q3YYmObnnW/OfwCDXNzUemRXhHFOW+RNE3eT12cDdfax
gz0DZgbv20dZ0FNYMDQqusDVvcx8SyNPpBJLsEEbYTXEdtHjBgmqXlTuZukrtHxmBDCpfCDRPw/j
6LZpQKJcnH56cBUv9ZlrfaNdfeT8Uc1v/ZUjRFsyD8/ZX0Je5pkQY5p31kflWvGna/ikLEXJDTRC
MSN1MZso6QajbZhcM49fRxtlV4TAPS7YoON8n0kzGKwUxzOMyHVtU2sEc8Q9oYpqzFch11BxDFjc
RqXcTu44D7Ey5H7JcZu5JBGHjcAVpwoeqzTLNwTy76Q8/kSsInJcr/VBCX7EKpJA24Ahi4HSwJNx
KbLs9pVXzU6ZiiLO6jaiJ7eMSE3dJYacS+6UrtZs7VBpsYP3NSoP8ZjJHJWIHEwhxUdk/gjPuHMJ
BwdyoGBmlQAd0Am3jj9bo8+Q8qEdJFS6MrJIfV0NPSOrGFJBlLxrlLqGJ6J7bYRvRoz/wsQPmNf7
RLTYWWOPml7itKbF3IpKe2+XedetZiEWxFSxLHKObIPhGBaFDaiq9AEptVrXpnDBPRy3OdapwPL9
ru98ViH+sK1Fxzb3GF4d5MUL8KO1pJEluhxE99gqj0f/rHwkRsBm2i5XnZENabwLPH5aaMoID1/C
Aq6jEiaPS8u1cBmw5QVcy7s8UIVHl2I1/bnBtCbXz+wwihLyz+GclFr6Y2/XQoHMaWq/5f5Sbqcr
Gzpn3pGRvKEsuqBgQol98hIg9kGXpXRdnI1T8gZ5nvdmYjXxU3ViIwMEKzXR4HRzqMHM0LzYFLDc
lAgzYkvIhoWrkYi2yHn5u59P4gABPiPM5/HWospa3u/Sa8YcnNqbzrRB7AcBS7VpNUthF2Zj6cnk
90W/PEpwUrrc/ItH8czsVKC1whBz30t5/lgoZcTo0GQgN8ND6dEvX5yzd7+RvEk3lcpgUKiSF4RX
bi07jd+socoIWLMVnxhtNXnNmq3C5Iws8OXe7JWZs/Xb/mH/UWL9vcu5GuuJS1n5w9cOgv66Xh/T
rmLh+qYukVHq5AUFOKnaWBVvZemZaaDhBH8JzZ47B7uy9N+P75Id5tWUI9W7YlwKgTQ0nR3h+B7W
oy3SAyQGb6o/lJEly823dQ5XXBkMiJJRwYRk9ARoC8yR2hYmsoAjEhimXlS6ziyc0FcxdFqMme7T
2zV+IggwaXTBJA3lSMaYYuSQ8Ug1v89KIY4xeKIWxvP/TJScyWmpPYBxb+Rg/e6K591shoEyO5ny
b6DzoMs2tfrxJCEvM2IxRnnHSaBCWFNyVobJgyYGy4OiiUMLs/DYgsiIG0bNYTZ4m73061t6Iw5l
BScC6o+p8NvUkHwnV6CGRZqRQ9D73pHml7mOHc0xJKBHVva9sS7o0Qdd+4dvOUjaFsM/fBPV7F54
YqlzArluaMfD7iAO0tAlTexJeEhX//TaXCfHS3i6I+5S1e3EzyqV3wWDZOsMhwbdMJ3C2Mwey6tp
u8YslOWZpUR6yhCyV2HhBK8dRROn0pAt/sXRGDvKn8NQQkwleyNmYI/NfTpUOjRwlE2NcrNB6kSs
t1rCRKGapdqfWXDTbgp6kRTQjMfOeI9wsJKON5e6ilFasxZ4pI2X9hZ1WoPAfx/hxLQ/1dW0Ni6q
vEt9dSlNdIok8gNXNR0ulrCi9Bq+PwPiEMi1+QAnJ2PyKNyqK7B+rR888rWJ+7GAuweAxby6o71O
oS8vLbtMfZkMIg0yt6JGW1ryQb6BJTTyMe3ubvLF9vhkNCJzvBCifbQdqHwX2ULWMH/wfGC+ie9p
G0G6K/yTbzIolGbhGhm4PhqsyvvOOSDftgG6bSTWCxDI3ilHjzlkJtAB1ZYpEbRQDE8ucnof2iPJ
OAIIdHo9vebUZOt52c8tXwDPKvOAf8j1424OkZCd//wCdvWLKWEF/2+X2mswCFR6OKOVAEn27D/p
mISQKZ14BLAxgtJdYyjB+PLxMQBBt8Do0C7bcfM/Gz0rDSxoXxPGVZ1e3GogYRfYqbeD9t+EnOHh
OJo124M35hU3ZNK33ObMdGow3jPWe0RkEE7Y0toI6HeGofTwnFGXjuB3QrEsZ0fA+mJEx2iXwWIQ
Vfp+u+ux3xP3V/RFw3yXtWdMbW2jm0jmyF17qTb3vRgleedIT6Ke1JPS4ph+FMPXtUUMGdF7nI8Y
j9w82N/kNI7WdYnZsXUmfL7qTOxn0+Suv4KXTPLyqJK2ljTvvtVn7uLBgczLaqVT5kZ3Yg8V3LJ3
bNLNhZ2hjkZO7wS+BjWKzHywLtVRLq0hXQTAxcjHSliBEQzFtHVeYEwsantthyTtfbk1yBTkEitK
eX297Ok5wLspU7/3Yu066EXsVfs1nb24k31VykobY22MCM2OKvbxlbF0UB8pkpoWnwiFAwpKwG3V
3quqVbXzJr4vfAIQXe0hCHpNzzyD6xIJoLpsN0g6IJ3leHcc72XZI06EBYRQmEROcinMvTeSiYQs
NWIBlunTNg7YJXzKZyIWkjTrkGYwW8SNohTXRgqHjcCQ1IeFdSeiRsBvvnt2GJh0C+HEh/Axm8+2
cdNC993i7QhZH02iJtuaPpumOhdkYh+70D4Ukm2jnLnfTWp+8N9uiOvz9zDXBsmlhT/gDDcU/Pnz
u0no/iiY2N2PEnBj72SmSK66Z5G2bDS+w2gO7yVnwHp6e5Kmd/YW+hWn0YgRaz3GtK4LIjb2ksg2
CZxCacTXciv2ASb+s4A3Gr3w6SUM9W4rDgzBMFlMHPkaFmj/0pU+SQFXBfxq0wKWm+kWAlbMV+50
+8qyOlAr6r0MJbf3o6XNSTbImra7txC67ECv7EPgVZ4qDkwu6QcYW3uNXLAxrVRuvl/jRmQC/431
XME4c7BNKtvYkjdHymTq2WnOFpb0JqD7MxbHvhlj2ylpduqKkYPBTl0kcrP8HjLahy3BbL5sg7hf
NIBRbu8es4tUH4eTaVu0v3nPrrNv934uGJbcsvS5HypelfZ5vg742w9qnAeP0uS3b2NCht6zm0Nv
SEeMcg1attwJE8lntWlHL4iwqBhp/xfmp0vcujs+BIKvekWMjHkI+aofFzsw82CLwTp2sCLyJfxO
k1+U7GyrAzb747SETXeFJGeSqEZiWgh2IPSa4MWjPr6eM0hoGPg0SG1fv4Gj8cO435Fpx6pvc47d
c9eoIbDpB+V/bv2GJII4I+fUfVvyOC13B0HzeoJvbR0oJKBdJj9wMa7J1sqy45BSjCmkgOfKl7Kd
beY5GTM7TUYJ+ArSIbN8MopPCf4won0Oekc7iQ/q7ZnygrpxWvcz8wQr/xVeoINEv86Pw1P+VQP2
+NtYOspHUvO7lfWWNKHy/KgHZogtq61ImYg4FPucFvmblsiJzhaitfv8gEo///2wZnCBpqdQltq9
g1TDBusoxu97gPtf8/KvhO4IrbJccNkMAQ/xXRZijK7enRAVhp5GcUEnznfVs7ata/JAbn56Tt5I
x4a6SXjEFE4DMhpAMXPJB9MClQpMd13z3/Pgd1493w2Lhb+wrLlXVM303T4wAOhCNLmgSqPYXAxd
OyDCSv/S3Wus4kvD0tADHthkDbYPoFDt5TYbePOCv6JlQ8NqHi2pJLGshNQAp5Wb7LdbhxnmQIHo
ZY+niw+MXGsrRYEWgN2ta33Rxm5waNWPUduyOhdEeoVVAOQtjmDvmmAdsHCgH8MBdW6OcE0lH8qx
IJ+KzuLGDL54hBcQ1HA5zsolAAHTpcxGGrgVZZrOaQqHCVgdNu7MmoPtvFIMBV1XQdJ3hHPq4hV6
HTH6ySbC0mPkJdpnwbRZ0dtY7TBfVJB6KzOvroLy7pm+vDfC6g07QHIxYoboi0LYBIjiLtXV+o/Q
FHrM9VppiZtarNZzJUfNVmfWGH2PPJ6aZs+QjmSmQBLlbzyMXgiAgQeJTtm3l0qj0HjNXDzYq1J9
uYJGYw5bLN3htL/sHr6rgmOOuyQlCP+avujliCRY3kXT3k/TjnQurykexOphYGAU9loXU3MnUzqL
p9kK0z+0rhgzHLsmWtXFxfArWBeX8CLdyulXsI8RRREjZYs/0NFdTLAdrtk8GaYtP+vNd2T4uM0y
6eqm/fS0xUioXbwMyCv9najyGOfWc3Mqzsu0Wx45qlU+f3rtJqDjFkZ89XaD1yAj3q82RMemoSif
gU7V52dSP7YOyAADVhaPizbBprBdADGzdWFzzPuGK8EAefmK+i1JP5h7RGApQlvW00ItvWfuwmpl
ayI1ZoiaHBAn8n0ZZwSKORSpS/jknj8HbLgHRwrdMc+265OxakRR/wL58bmvs36CX9vdW7k5lepd
vM4wAyZA0atYpUzLIUjLghiCw7H/ifvjPLDEn7FnLsAAo0/4W20NRCUNYeZIx2wb2+v2Go3RO2Wv
uq9td4iBUWQRF8s7+LC+qIKC+lIyJPv4tHNHqN+Jrv6mgvW5M5RJUbej87cPUZtCB4exeG0BeTax
0efo3vrJCWh/hsWm5P1oAKehMNZu4xhXc6GYUn7tshHRAMB1/Kw4Md/DemFgiRcUJkXtoWct3UWx
OCCMTsH2fOEu4HEqKeFQ0YEr7/k2EsalxPxCMgY5uUUy3/821mSx5rfwXWVu1HTPmdNOcoDhQ3Cw
5jYRyopQNr4/l/YpI7+tvZFHC4ssOVfwoz6YnuaIKWbkNiVYg1qY3WYP1ryTsEwA7zWrfxTCR1oE
Qj444lkNpBzmnIO0hx/VF/sPsbDtVXV98J6rSq2IzGwgZYAxtrc4t9hZhAFQODtxR0pPspaj6HL0
fI1satHMilDq90W1kLI41jNoSRHzcBhyuW0aYyCzZap6Krm69xGjf/ngYGlMQvoxFdl/k7XXsjkD
/HiPMuKF11b+L29dWUgZoZ78g6VtHOYCsPJ7biLAwwXfGaKfBPX873Bfre3ZSaJdJYT3JVA7Td7C
Ekl4nNcOIpWU6kluUusW92qzS5hLT8fU25MQ/NYCTpSIGYxBxt/Z89GXw0DndELkPtOjU+xPeclU
pgHS7VApth800f4hYLOz3hGKzNF+sske+CIkP2fxoGxLJtnMh3PDWIgk3M7TFOa/NtGRLn8gQ1rk
jHRjg7Hf7Bk19hFSyFeSiZNrHyfVvlaGroiV+KnXztCvKLlPnY3MgAy5NagUs2zlteRZBcqo31ly
ploWRCezyXjXX1plpWHvmbWow8NS9uSYAu/3h1bar7kClpFkmlx6Qb1wzjDv3/nWzJGk/wXLTEsP
yCu8jpvU/n53ggQeFv/ApOEMgJhEgyLA8Dsbb8TaaQuaTTaEk1JKdrlr8dbThzwMpET0I2qSEew4
JJ6VbpIum1SaFvK/oFis46nTyGqc0r0dWU+58zfHQ/mjWdl4mkkFFMT+Su/xYrMWjqaLIWmaHZrt
DBmKXRFEu5foi1RPOMT9bov65sCY3qmXb4ifCdyjgW2YXGZaku0UupfLqL+Hy/x20A0COyvS3QZM
7m3rRqpjBJT1HHCIDh/Uz4IGk8EMC/ExJj0yKUDTEX9j624IPjm37bOpBhqOW0L4wNVHBOvJz0vQ
IkHSlxYOXmRzMo6TN3tPXvfGVYP0/vU7mq3siMGfVNlGjLtqq3nBDe5+82Kz2DaA5jCRuWnepzQT
U2erVgPah50YqbSE66STsqXG6sONUXmS3zHf2R08mosIhJcud5XNnFBn5dwDRStWzo33bMS1WHWs
jN/Dx1N7paWvE+j/EofbGUfaN/j4FElbTG9SSF0j/PBz8iU/SAYwvCF2o8jSkDSOi+kNcYZ2qn8S
7JLCRimKKro25g61oUhwYLxepOUBMTHAyb2dqBPLBZ2vkNjpZ4N1vBbKKJNrvA13WeGWHvmk4/CM
9r+gqCND+/JrLobIdqAokDB9NaQlTGa/WDs/cRZD+4VIFJnqF2zs25Xrxbk19uVVFllGP9+kBVtS
+haQqZGJC1QuaUmoqTygeT5FDZiD50lknxHMUJpNsm9HLMgVxzyiCX1mpOvJBo8SVJu/Zt6X0C95
2IatMXlp7LZDjqCr18EFv1OWYz0MQ1/NGgShj/RhRTieYSIgVfB7rgFSUxlu5AZftAYBQEnd0LTe
Xwfn5qfsL7a/7lQsBiRrdurdxKe1FNNDgXIL/9KINQSDYr9FNb84S0ZaUAsAoigaYmcYPgrGO4Gx
v0fczKuXPDv2b+Rp8oofeYissKFLD904he0L4RTdG5OUIXtOY9ndOm6zeHGPGPDE7c7vYD+Y9cz2
EaYw+ZyboZjeaeq+9ahrAUqXWIv3X1tAq64axNkY4cp4w+jtZLH303QC4uvAjeHhcyI87RgKtMOA
QhjShMIaZFqcMeWcLLPwW+BqUSof4pL716LnNbFLZH4JybfaEy0q9QMrZrfu7urpxSjFnzyhJjBw
5aFUZIk7F+yPhcJIGXQFx4SWHt/uhvXRYVnsueOLk9RTx3t9AC1sLsisnjcQoewXtHF1/nEaS89v
iuXDkerWW7YH2Mm/HlLotGZo3ORm4qSZdkQMYsjpfYJblSb0pkD8GnnZzAHGDWU1gPr7bZhvdQ8N
O8MBWgQZEdBNJlINlrdNSWIg8MYH/HrUmYqOSBgDml+Q04f+b1WTVXl0vhfyIlIBdSnBUYYAIrf6
DQadSiWmAk2Lz5QvCkZTGpIkljkrz0RavwirI3m75JrdYNDPXVAAY7XXLbHujJrh9+4BzvryEncf
hFsfm6vFfD8toiTPowA8nIo3aklub1doNHijfQfF9HDlWxTI/YC9Q/cb+xWT5aEtqthMfc+vyksw
gwHn/wqRbKNiVDqZ6Hw3tk/96PW1jMUnK660oCu+BujfEwqGPU7cffTR3WVzE2AzGecTCXKm+fzs
WBFP7HTBJS3ySco81xirjBoIfuyXxq9ctq9MMDlf3ylfYK4AmQ5tOmJ6h4m0HV6bTqLN+vhXDzpS
uPMWfl/XyB15lDe26jioc6v7/hfMmo+yEPkvUI/xTk0IqaLb01yY1PwPI7i61iU8jWr85a8cGy1A
da4OALMzReTgWFnE9r0nnOyl28jWFDHiIMJJLJ4ZIhRehFKUAIgSsBndu7Z6dhXX5fxiMZkaS26J
UaGO3QgLQ/xXbuxiBvLYhtWBpSQXGaRTC5xo3yyit4wzjWU7HSnMF7MJubfnFVPY6sK0UAb04KWB
CpiR56pVcRiZx2TSGekBRMWqn9WkIVY+MT+HEqJWVh/yioQynP0DrU8JyRa15Yxl1ZgdOF4Kmc2G
Z1QPP/4OBOEKI/7KbFmHyZOKAbSBNvcckGN8FxVwaTw3i1lNDq7ukdtVESYU3eTReMc+UJucOyvf
aCuT3a6+IEOFmr7Iy38yudtPSz960i7I+X6ZPRiEhOM3h84WLLPgnzFjl5vJ7jVMAu5kFMl+IsBU
vJQGdzl6oGtpTdHdTzGAAIVINzwLit6jNP+5txm+5rYq0myNjo8RqnyZx58JalMm79uIRa6wzMWy
YAMUVL6g6NY94pjU/dzIrJY/Jkg25nBYHfriUrA+ki0rC+13eDLVLIYRQ6KwiIdjZLBDQFlfE1JZ
J2ffPj6/1Za+6nIetXrofpDB9TbhH07DW547GvTnwp/4kX+LrQLkJZdulzx1y0I6ZMOJoXm3q/8e
BzY/yG9U+c73nfwzfsTK13ZmenK5XRrSqXUeZHJsDb480gaHrYoYy0WHYb9rymne+/1g4fR5SPO4
QvovWnQDAMR1ouUmFDgRP7jBWLbXbOdYJopln80qKllKsIBprNlOaga7zRWu3ZagYMmkNPHhA9Ht
rMXLO4b4DpXgCvdjjKnWs9ytLhpfo9LXE5FSvRcEZYecYQOtU/bimx513wLwlSQLXyUbVyNqodox
MT+XGYpX4GVIdra6V5ZBWefY8VoSCKT3w+Oc/CH04IOPVrTXqrgeZy4r84cD3G0V55t/QbayBoUJ
oGA7TpuwGpu7P3AQFtiP1LdaCmCzi9560SjJ/M9cIUuOn3AXBXxcz1xmhAdFB6zqjR1hIrrhp+au
c6Z7fRNAKMJXYsf2LW+CbZ07ybxcgjvX14P2pGNpU0vYxuh77QfFYPB1vgEDaI33dmRMWV1u3OU/
7tdUGLkZSk9WsR78QgDZVZtX2aGlAluYv8pvTquYWtdyKfnnNTPdSZiyKQr78qSfBqBh8gJjUC6t
240bYxOU+5TT3qCV5V7oOdw37oEbk5/wQF2DzpT+27R565t9Rh5nNnq2UHJmZ8jBYsVN5kgnmLlK
8+wYDavoet++Cak1EZl0vS1PwW9l0v/ScjUykXkrwz0/mg6I5KyRdO8Uqnn3tICtRQGqFoY6pq79
vr4bIr2FVmre8NO4FWwIIbNCenQa9yax0bCnyJb7+0R4LW3DdrYiZ/iE9jsLURhwyRowr5JpTejs
Fxt8bFWjmcrxyHFR6VBPE0+rLjaDURMQoSn71Cz2FVI5eycyisKD5J3AIpsj8ZQH2HcbkibhRKtT
btUSicUdj6yQwQGcZX9zs9B5Mq0ou4JLzwwDs7FdY32p/37JTZDzT7wmpHWGtJd8wmRZ5OIsIjJ3
X2wrYNR0QEblUrXKY+V4I1gla47dhd9bmAoQ790TUblilM/zmBH0U71Lc3GJ0lRKJHFQOMe5BhQb
ZJtha7eNNMdUGqyJ1vZJXSBF2xAqCJYLAGM7GuEkO78D36hnBL7CLCLTMRZzcTIF62ry4rQ/Iegt
Z3FFIaf5tVPhJjQPCRO7Ni5Yr02XO5v1O2Yi2e5Z6vCAQDmNappZly7FEjAZAcfAnh4D36mJ82ro
eM2+ITeyNwoIvFneZSsS7XoSf7/OMLTEFTFmkx4qzoOqgNVlI5O+0bHkjC6OMYul3MK/4/T3mXC0
7jyv+PVdfYpmUTSX6O4o/rIx68xLZrmYuiv25wHXp5oIVxnIjukmB74zp3L72j39TmBmFKN/3wfe
fA55gsQ/d9AsksaRnk83Z7RPO3y73X/cdV/AtLNHpL3OXfp4eY0D7ybTsFY4I6u1z1qtO0mcsQH4
OxFsDMNgS+LVIBcSAOeKY5NBUV+5qyNciKKv5lQlOuTGDDABNZnchrsT2Yj17S8IbOflhBaTgWXn
WBF1sX4BmdDaSi+T4yZBKNlVhUbxduoChuL+5NF9EMbMPN9xZVCjAg/Hs1vjNnlrEjNUV1BpwA5f
W3h0Q4E9MZ37oiRZnnbMIX+eYeHDrx4FajzNPkdorFTugKtmzpw1McvTYSFI3zPSfbS2NwlbJN05
6rBw6agv32xA8MSCfZd/IWfSD9oC1D/pT3gAb6nYkq5aJNfW7YKAZxJQS2ooRkHIRjnLa3IF1Ory
lPemGEeV7wAARYDvPr+sQVCKKsDVWr5jTGJMY1ilfgZ1oMOyfv4Rrftig+a3aPO6WABf5Mu2E0N1
Wep4+SBZnugiJKgATLrolOwf9dPMIU2sYM+XSfo2mYlOgXMruX6LqBdNE++LlHPuEojSBFwHUDri
ohPyTjCakm/tIMomKbw8pQ6INqR0B+ZmY3ESUvmfxbliqhHW/AVdXQ/xyelDUvlhYBmA1lQXINz/
Q+Ng1Vdpgh77s1FWkmvD6yASpB/0xhkdwO8SyKqg3aTIKI+k2SCRxbYL4X/UQZ2UYFr/vI6UOBKi
quzsKQv+zBJyexShSkQfeVD+VaQH3tOncxBzLlaXTmM0WzFjFkWb+gU+G73Lyzd9ZvGjY41godEV
pzQrUZOMwgZhxTMRSbeDf06QxF4XFFcPah8jmm2ceUqtiJ57slfyWAE7lSvfzZkjL310i8AXZcnO
ntRpvRpnwMV71rUdYiJV2esu2zYeYkBCdiGOOQsovytcB7pZOb/LhBpuDnu4UlrJSen+dcOWJRM3
W/D+owdlGHyHXnFRjmwPAQe6pZ+sBSmH0b/WQLvB8oe99pNt3XDKKrNwxBTRRMGmBvJd8hp71qn8
poAjbzD2ajvSgtrnc2hBAWawG74WPQvBK0zh/wCEOWcDvv8vsu+dt/gVOvIyDhvJBJoys12O3Hd6
FQ9YUBUQBiBGbTPzQD9xEq5z9fdd4z/O4cWMs2J+iGpUWNr+MOYwr5Smk5ZvUXn+znMe+un1gUqS
NJTQrnMNag4qLAKOw508SDX+6n8QrnSE5gS2nk3rc1qfJSxifE4SN+hLmEd2Uwc9faSiUAkeei3U
36zNzioxPUZ0iIlcbUW68v/CJw7V91M1u/0hz3zzBKAuvqc+LcXmxV6t9YS14rt/QM0DP0AFMjmw
PGBQuqUnK1VPwyZsyTB/lO3khZ5Qg2dNMGWP5Q5O+RWAD4+RTUXWLb7k7Alpl+eTXhb9Yk4hv1FF
KBrs6J0YZL29J45Hyni0hN/kbOdlbAmltU14pTUpZJR67UXURBo8SMZqaxhpWwaLy77rYhrbif5X
/Ue0FUvdnimznF945WzBlCar59fNDVH+/hEfXge7OKj308SVaGnFOmG2Wl1KBW6LmGxQeMGOGxb7
fgqVfMaaeaFpR7w90q7sMeYCjNG5yjT6eqLvXjnD7EQZlMAS8LVHLz8LkUUHRVm6KA1kS6jIt4Fe
fJpugYpvcDVKBQ68UtpsAkB+ykBljM8XZqdI9fTDNIo5vYn91pBVD6XIAnDbTYgILr00ppZHfCmD
R6/4rKeKFS3ijiukvBiUyVcNcjE9BJhqZR3ZJSGuseHEwNxBeALRncPtK1ucEWBDXMO5X/w7Rdqf
YuiVjkC2IQFAGTe4fo6tFEI1AJMNSY66MQhRgdgitJ706CmzQROlq7U4qpYiLEv/zj36IQqhEbrL
NmTS17pKGudsn+RoBuFDkwpoaTFwoJg0707nfjVljSm2o1EGXp/3YBssrQpC82qn3kRqYhjYI2cw
aGynRsc/NOgzM3zl+SwqYCCU6HCGGKKQNnM9mFBfzP0uB25eMJPnB8LQzYCikI2tUMldAXqCNGsL
ICab/8QXgHF1vj3zGKsDA3l7KpznNkQ2yC4InUnEmC6rl5CUK62wbCXwGwDpF5rIinMV9dfVKOLV
pIVDqIWBI2nx6A3VNWXRn1A6ZcqCYAnW8ez8Ap1vmAgv6gxHXamVqiVPK9WMW+xcGOxd1OWUEtrU
YQnmA85MDLlXGAklxoqRlFHUkxLLRuUzzZiFoqfqMfzn8CXfWH3UJzXLoeX5ZPRl4Fa51GpnhcXx
U1nwSaH/5MlxvhTz9KeS8mzdO2MuDBo/dIJtXJ9RlhVaCbaqTDL38ZDYb5LWikZ7ajBrPPHcAVBZ
w0X7zro6U+5F8xIbPjZ31+aIfdG/6isNsPZu8V7/wrFPTVojjx4Mo3+1bLir/fwqzarCxnY9Xvw3
qaihhTdhNoG5YYAo2KX4AcEl5Y6F0ent7Glj7AWf1fkc+zW8UN6zZuv8f9tSkK6XjfyChW1ZzwhZ
2tLpKJ3Mm9o9iEapqaDCmcyQdji62dAo5byFFGqkALi8vcygedQ/mFF+onC1T10m6T8UR3AjxFpb
Qu3JyMN6hpJ674IdgaofAIcGaLlcarWJdYnDdEt49kS/hkuLbyQ2pZqRsVx2FhpBN7kUPkybDZQ0
4eRquSfl5rQrwTUPk7gemFIRjxb5U9vthnSyoJadyLBGcMhBA1/cgq8FKwJFhsw/xqT0QS0uw7T4
F+arNn3zRst+H3QcRJBdJLp3cVhmwMczmz0jsTFXe050snk/msDq3FVpz2OY8TbeQ6WUE+4HPV/S
TaKbaE7qYxhvJW1eqsl7Z48SEIMps1dXDlKwrEv4TqqASSwsUtA6jWvXK60hiYbCh9NDl+IkmWjv
NjcpgjI3sMCyKM7vUqne+dkmxf75MD5oxh9bp8OtznLfPnKDSz/3DRXA6aR0AhCEesomiGUrmPRY
XuWLXpDyGNTiVuv5acV2y1KtktDDNYmSKb+dwiRIgFeeToVLNxRkBMwvvTTkUQ7cXnUciat/LjQ9
pSAMwl+PK2Sm+1SSkyVrhuJtOU+lMi1mhyHDcq0wJJT79GUXuaWxf6k8dZUnpl7iDbDZ+nEMroOB
14tQkAZOfSpw8/ss/3eSx5YcsmzL0AtLMWlpWMk7ASAJTgrbNTzyctNB5OMvXBKAEFm7pJb2SmCD
Ns408hSXw110PDKmRvAMMF7/Lv/WqZMUwDLmwj4KuRpEuLGY5StsA/dZlD+J0Wrjv5E0bAa36x/z
ZPLUjxeipSdco/utWFo/S5646ZNQuUk0RUUKn6WWLnqQ62sgAYxUrb3T6/XIGi6NXhpdJjruER26
cexxnPHWIHHm2yw9A6e0d8MpUQI3xkemUJoNso40t6B2Ze74kFVN+mzQ5q3W6L6F6qYUkC6S/0dX
Cw9n5dgHhWzq4qegTsKkF8EnO4CGtjiuwNix94wWixt58nxnMap+tqO+TjnGB4O2eGlArPX29dIA
b7WsmOOCsnHpOjVlo+o6zekTvigCr3hb3W+x0bMpnWrfU2idr1+7A4Be8JXcej9gXxFzV+EVWZpO
ngQfa4nD7zhqclby8pQRplu2m9bd2hgriBukq7sodq1naqHqpCMGsHWm3fABoGIwvH1xZYk1nygI
hCIpE9K6QqmlobRicYS+dp0CDbRAWKwGiZlx8Mu3n4x5EURBs2DPEGg/CWA1pwhPflt2FfYmlm62
xRaRAYMoZsKXq9pW/WhqCY84g+BhrArJrGLE5fXWznOX+HZKRkEVKF3iy0qx7j+J4/Z/Z2QM4z0v
PW3uy0Y85h450meNCVk88MyLKZh8Ete+aUKMWal2QYeXpnTDYiAJogIcayZUOcnXRE1Bf3n/j7Vn
yqZ64AemvuQ9KR4uYj6L/wbWbF6WLaoi5kdJg7vWmwYJya1UXr7rvk7jUJ3bfO+B8hVPKwdyjLlY
Ne9zEZOwR0Pamzn/39jBnOKfD6brv6SEOPmyT6lPlpN871TebB6XekvuJvhScytXx8xQl9jsARlp
U0tdIC3ubnvcTLssw5Ge4peBANJEvHt1g6lT9zJy85qxfK19JiaNON6wmiZNFJmqzhbeY9Be9E2k
BrWZPUzAL6wtWdVe46UNRoxDzbagyXDVxTVB4XWw7oMW+P/FICWVjNLEQRFd/ikaN7qDmFGSqcHD
VFEdBCx15qEC1FYp6qSBWNWmGtIXD+RVrWp1V23/xrRDto06B/wkDYyBvMhoPuuw7ROgwY5CLtug
FjABDmNoqVJDdRfJHIc55XL5dgR9yh45ccIVjfIDTZ0C1J21lBc19rB11OJUw1ODO1eoE/BS0SkJ
h/BNVjC5313u6sfEXViunH7XCT3gdx6UKu19N+bAldbHEWXDZFn3G3LKXSjDmRt5Z4mfz3NnKiz0
XGNyav91nODzk7uPOuAsJ1KlSB13GEXuwnzv4B/NeIB6M8JHtcNWg517GeJfMISApsSaK2Nw1vaX
i5gxwQZaUdmmNxUyyrjNSjTkoYEqmwrTh2GpDT82YVsAPf8MOnW/4HYQxMf0i6YORUVzGRKvh6tU
6kjrUpUtQEMVN6YTpchZ21Wx5Xd3ivDPsYHK4Rw1jWkbcmFSOSkh9gcFyL43EP0HkVyW0AvBJE60
anFJXP+pkUdm213HHncSfhkFWL7AB67MM0qNcJXXBH4jRgCXK9zBks58QqrEYh4s7fNNZq/An3j/
gSOg8D10xXpBTatXeXwRcTAMDCx8iyu1vQK62prfFoPbreXeV+rseyWrRY3jzQAN2bb2f4pw3aYy
xcUQRId+K/Jo/k/Fsz4T08te3uBB5ZB1fYS8yim1i736DhgNXvOi5KUl53dL59kx/8iAHrI7auXP
67YxXpZ3vGzxicRCkE5kPA9mS2YVMEbyI7smizRNVfuihxA1r827T/L+n90ZA4O7OKXzpkAY5Zqi
wFPdb2RX8GI5kRFvjiV4LNQRJGLRuXEsQ4Dzg7VEUHzJEBPnEaxC4Mkc+4REGq6y2qnyZiyoUTSF
qrjXZ2zdMQa5uIZpT1U2fSqJalVLFsgTE9g1AIH0lpkEvurtUSbDdshPHiJ+iZLBkekVrgJPX7ZB
p9m00uwQO2msxJ/xODID59qahRvcNufHehYwSOuTodI22rpJSeYdOZ/URtZ7yW30BuR+XTjrAbC8
hEzF+4QqMO7mMZ2FVrU1jWLTsJB/ClKd6loc22dgIRNYGfFKZJE9lzU5/GtOKFPyETBHc69y8AIE
80mXuXAoj/noZOfGKShXb3cMNBN603phhMfOMEn5YRBu8d0RYKFGe5JF67Zxoxs/yks/Aw2TZFkF
ZDoatlst1mMpprZoPxYuqPixTlM/0H5ny3/uI3k1usDs1nM3YgG1iLgQQLqJj5yuZzVyJ1b1+m24
OBXqLmFPxyuQwbkQXDaSJ+GrxNZJhmEmeNq3IHx6mpg/Lytul1TKMpDh1dpLsz/0YkzgUKtO16as
7KexeWsXWHvpIo1wcm80zHhTC5LmK2LdoSX0QV3YjSl0beMJZb2WdIsByG43PpJQRpZbN88/5WIJ
4KSSBndCYDG+kvM0S07yn+ortvwx4ycbtAr7e4zcUUBaoRAEhroYf5zvUqDWR6DES6WI/RgWdPwf
Bp1/SZlVqLwNd2Wdg1aSCpdUV3zL7mk36iXYUHI1/GY6HdFOW6ENJT2YiSRQSlf0aDvyJhYZ7k3M
XAT91ISNFMUuo7wNz4MpCGGqlBCumwBbYeg3tQhcAwClvD1wrAe4oNdJA1M1AI/ue0wo/mz4AfzH
v9WLNTMGaTSSaYqHljEwnjuIH5v3rW8+h7IfFJ8zqCtZlEZNj9eQ5HJc5Qea0S7tkr8QO6otcW5F
Lv0t06yBrdPkwDhDt0Y9iyqIZCDpvyXJ9k2B6CqUL7FUMjZ2s4SoxBATobHYvvVhvrGn4tpPGTag
JMMwhEU6bQHwxVAc6PaPxKppLEjCrP+FYJxHDVNoNOYj6KjdRGK5kJlmv2fyZTOYZnOBReKheycL
cIXIuJOQT7QGL+GApTkl0ZtsJrGuCNz+qT45O9XG2qYiFFp/iPR+nsbgEMd/SxdXkOPjH5lAJcGQ
x1RgLWkzA9ETidrRMGCbh9EGrbhCFQXyq5IxSxNyvjHZ5e7qp+d3EVk+TDyewpGwOCl6Go1I2mdx
XCyjl1/8KkMovEZSBE3ibDAaSbprYdRe73bt+f2ZykZNlT1AYaG3pumDFKnSLJIiE89lB2lNHQCt
Ll6YnxjMGZ6yzrBy97O/zY27ifQMufWiSaK2MWUcNZKf2mx1pneG+YeGigO+X22GFq3uR+ccCIDV
Uzc5SBEPETvekk4UxY1vja52rdFG03qZeqxBHxSx6BJ10JQu2WBVOV5xIWls01CgjYXSpXYLW8dd
1VQQnjXvtenNusJq5yl0q61FpCyRj6h7vdw5x0BXA8Q9NfQ/G6WEQd+NPX3IxOajPIkAEMGlgHVi
TCvPNZ0QY3HbNWz6hR025TdWnlyd7/oERZaNyqq6DMSaj4x7fVdfFsFwwG06UyfMdjxekMbYzWfv
+qk5GfqGqfunw6GHtFWquGr2pq/Qg/XrafLhgSdp2SdLFf2Ld1mLbO3Erenu8oV+VtBHyKbUst5e
w9xCNUN7Nq6CJjNFbKq3Atx2sf1uwAfgP7yhax8vKfjtaFys4vzId/BUV6k7pKCXo6fylda/rdFT
c46J/WJZjUqRTTQ6935aliqumXr1a++ac1D9/TL/KEaTCG2AkQ6dogmrzQyfvCcMKlwyCd+cwc5m
9aEh2YLeF1x+sXEq01SPUAknPM/yQVb6Y8biAvi9LxlaYNrGrfZDEKwSD/+Xr0Zb2KApQ0UtP35E
zewvSb7KzDUJW1Y+B3+/SziTX6UlbbQgl9HAwREaC1TBCj0AEPHArziMWtsOTK5VlZc7kDovLxL+
oZhyVBGGD5DzjMGLn1EC9KKz3t3Onp1xqJYGu7hMrLtFkv9lBVChhr+y+FAOFTuXaobZ+uI9v3Gl
aNWr9tVazgN6CrUTwQvFaryHV4aqFjT9A9FZ35zsJPNGJx+kUFP8ZM8yuRoxod4UWgLK7OYjg3m7
7mdmwDYLEeggq5u3Z7rU0sggG1RZ/FpUS8tCyS0BW2hQpJDYXvOYqb0Q2eHFFahi5OWcejcL+mmh
vhye6GbjQncRGZBJUg+CCXmRRAv3iogb0p23ss1jAQ2pP6aYMmTl75tDd1YhYUa2In+7oCaUfUdl
KbxS5XUoJhAdSdD6tVSVWSzNIDM01mWvZgv9xHZUJYettFeeAmqfN5WKEWqJbgAgFY2VpwzddA4B
MTiRk96UGKc9bqdkP/IivXDqjb/WjGhJt7gWAWh0Mmg/9LgnURgBBf4dHPSFO1kskhrveBohAakY
loNP+kzp1jpsh8nIN6raYvLOWNDHOvz/fwdz9/8sX5BU3lG8IV2WDKmnaVxNLJxdkIyMYYcDD5MG
ch5RjAcHS3wMr7CssvIJnFIjgYNegvHkPev3A42KMQuvRYfEdeKeHZlsUaBWps8yUofPYnAKYEuA
BUgAGKQ+ZNEHhGRqd1HBT6mLcJOw/P9WGdczjcdTWP6Jk62RVDgKnKBJ+in38TTYMrUaOElhp1oN
nSP/psM5+BWA0hpLG99lZchqL4eey55P5pphF8ypWy87fowzMCqC95UP0YtaXrXmXUr2K484jAb6
C5LTdwiRYfa1IpcKWKn/K+SHp+xbjFE3Ofw5jyNXooJMN2GgcW3SZxh3Bc/NMBldW+ixdSPHPKij
bBDMUHJdlZ4I/u9GlR42MgnCoE665UKoXVtW3GNlw0cjdlKptiZHJlBKQSNBwzkv/E+1jO3/QvnD
LTDAPle5mzU8A5aMns52Z+HrYswbbkY+naCKYI2wDfxhR62vRgydPpGRxosE5PE5Wd5G+cQNkP69
9NcOHBiqoqRfIDCXAafn+j2l/tBXBJ6MVmpbRNfEOJIOjb9K/FIFYHQ5kQnkXuWJRV0aCgf3yZ2i
gMZNkvI2GjlnxD7GkBqP+RJQ5N1bmLoT9rQEwpYNrDe3WOEc5jIWOu4eujtVnm+kYIzoJ6ua7cDw
EWOimhAIBt1vSTguJmoeO/m0GJzwNYjsxXv9lVj9i9hgYOrfroC0xMB6gGvBmBuYa5yO1/SbGaLE
z9Vrf7VdQOcK5bXIl45bsMDjaQqjmaN0dRjzkSpSfes6315d/obFud53JeUEkKa2Y2pnUsYjonqD
QDbbnZ+etJwC7Fa5YDbD38OxOMIrQ2ESTvUbuiUaNmEfVUiR8BvOcdigE7y2Eoykxf5vzuH7Nj5L
nNb/VLp8ENKfZWcrFnBSTUwVcHUBknGi254FOKLI3ZV+QEHyOuLy9QBlJ/+Z2OlO1XfkvCOSOt7L
lBXQfVD7nDSleKqH9qcDFxJn4WVZdVBV8acnV9L9y7TiSEWuFMLKZGBXoxSYhrxHpqlIvVcurpiZ
zHZviiEohkU/CWlrmy7S0CXhry/m+ckBUXDB0iEUmD/5N+CHWWe4PdFG27kbeuzumEYLsZzmrWWi
bqfoQd3H7q8wJLNPpRydfteP72Q/WqTzfPjp6rR0i3wnaMEjohD/MUFwEPJlYD3qsoGzSWIIryDk
Gn1n29X7c3uy+NJ5lXzFr5mMfmY+GChhAQc7UU+77nF34k62TFn4/6zUUwLTPTZ1TN0BRR4cOV02
Ig24NoKgVDvEkp4kAjs0aCil+6pdpA01iB4V4ataCHiTpQ/C+rYK3Yai/rWdzKJpt3VDirXUHrno
+GXrx9NPPLJAAEkC3ytvCvVml+rTqSuWi6vhv8Xyz821FJguiv01syD6Lk+2p4FCtHIB9Ezb6Ywo
S3wn0wghO/L5HF+hq3olEPbDCrZGk9Mo1kMDg0n0DR2qYXWmHsWfcJI7JxjVVeBt/g4QKNOXFZMb
wcsxq5SYrih7WeIoEvF5InTDBbv6jWqWdbUVc89lI2yQyKxnqeJzxT2TkgFJlBF1cJpDeqkEE6lk
5xVbqgjX3ZFEw61+DPM7141OC7kcGKlxZQlIM1nQxj+AFr2be5W4tdXzGoMWalLdUXc71YzuXmbn
GnyNKiKqIJx1KsEeTZfONnjwNKwyy+R8MFu3grtIB5lVzqhPJqrzz206nVQyxxa7Cr+5BW8lvU5j
DVej40TczJqIE768/UF12M9WPSooy/vMqho0KdDAlSG7KM68Z+pjjWmIi97R2B//Sk/o+w05E8/I
I4kXJYZlwO8F3tNlDkeC6L+eEFOfbLG1h7XwQlm7VCG//w6DZ31VSVxoy7Lg1s9G7BUrHwELGpju
I09ZGroPbwFHXdpvMiTC+6sM/6bfKabkInxJoT6d51WgNkywlN30H0tbZucgvfN4uEC0A0zJwMiI
vZAl1xK2zCvrfcZvn96ChBOUxjssVNBqoBirfBQiZdCEIUTCz3jlluTqrraxZMYl4tGqmHCtNGxq
mvb5SoKHKSOEfziecMBtzgb8ZcJPBs7UmLadvZSBXlIXWvqN5Gc+HCGcJAwQIRDQ5L3tNWZ6phY7
X3fdNLrEamzbxDb0s3j9DQkUWrFRa+6w26N2USV3GVP9DXA1ri4UFAZDGwQBL21nrB2QBQqsllzm
0nw0JDDl0paLrx60ruLnA39O2kNSTZV3pqm62RTlx3jz9ELe9+nPJ6jO5RBjwi6pzSHjlwrkMdqW
FaJBzspM3NizIRwrPGaiA9P+rVvEtW4RQIe87y5SCmsMrOnYQn9wihFxD3ZvLojznza+uTnYvyc3
2keTZE1haAj3Hkuqc3gD+PCRCwdC7RbozTW1QcTTqu3IZQqEejtuojGiuCFkfRZKX8UVPBeahziL
PLYbCZ9MMdf/EVa3o/c3QRJdrZpLj5G3S3xBYuDtyoyp/ZQzteYChdali7Q5pjVCtA808gQg318+
wXPnVhubQFpQAZjLWlLKvnMcgOBAjQTTAEx7OhNMbeFstXUaG6FUOIX2dlFPB3hUK1ehF89xlEpp
6VFPDgXqC3p4RflpTjq2rg6QxvR2xP8rJ0wX2gQAz8RAUhyg4igfRFRB/qW6tIAYMjbLCP+NKAhS
TXGKGGTuF/T8X04WymeZzDeIi7GUbeDoOh4q+YPPOAUZzLQsTEuzbtOQfSM0xjbXctmoL5j3rHIh
OJ2pzbbgFbWt2FbTOpJmMUM2t6GXsqSp6E03wRT915RmDGniv0bkArEUpjuH8LMfq+xoB9T6n+wS
dTNt4d9z8H7T6uIKrP1dQG2WtQZQ8MjretFIPPuxWhXOa0sr1enkmg5AlmshLHCU0eKZKkxLCwPn
nwkd1zvvGBrpfvT48C0fEKudAJdpcKG04tnN3nryqXjM562d58IDmh83huYKicvNr1AZ7rJF5rnc
ISCDjDFgGWYtWSyKqVaJCOP0jXMslBZWdDGfzIof1t5MBshaRpecoig+UPL+UABXwf0eWE+TvHT2
sm1Afxh0MVkAQ9D04Lp1+nEUCJHT0o19WIvOaxeYXiZIZMT/NWIoIb0laD9HRg4sEXsK0BXa0Eje
yE+woY3t7C1QnCCclIVl495ni1cIJcMue1SWqEHPVW0y9pUHk2pKUJwq7XxCcvG7qsqV8lCOUbeA
wiKCezjlxKSdREjZPT4VazSdB5psf2hOqTRXS0w0wjF/fRcoGu23MHuwz8iCpkpzS9v2nmO2cpht
pdFdoeTolFqYHVKO8H9brSH9tjMMctDSWDNe8Sjde026wVHWE9sZb6OiG0SF0kI4DsYuDaD93SQU
zSuOym9OS+WEdMk8Hth1Jt0NdeRZfNEE4BzY3kPAr/XNqDSdE6wY123hhrvkvwy7sj3e1pxXPOe8
RCMuaM7RNn6ZFlfoM+Tix/ms1XS7Hwd4XYfwcFk/wL0u2+4WYbfCakd6urlcozQiOuD7TBYv2UlP
T0xr/0o/S4IDisXM7pkRozmcWw3/+VnIZr9XBteDUg9ui079OWyDyly1jQcY8EtpIQA2iEgKT9ph
9AUmbcXe9FkvozOmEGP6ohpFk5AURzT41Mr4UVo/Sb7YhZcbA/7KpJV1s1KuLypgUMgW948rmVHQ
xb444/7VO2a7HJMQ8hXzaAimCdGf2uyXitL2A5RmN3tN3tfUKjSBkHYxluFRmWXRxGTRjS03yO6z
Tf6GclYG/8xsdlOjelPDXUGTNpqPg4ztsL2CtjVBHAzVrjzPAB4LOsXJcnoHjKuyBMYSEBT/8kti
lVRPJOjF0PP/DrBRD64QflHHURUy1qIXAwEkG2g0yYuct90FW2gXvRBTCbxKxCnJ/wBtIcX3xsoJ
5qVxzlSiIhDRJdbwB4hkdXtg8rAeKQZ7GnhrrXHCdT3KdjjkFrQKpQIHdWblaqiXQyPq5HRzgtFX
4HTi1d3NQQaJ53hms5D53jsS5Ylq7uf5j3szTDe7l9UQMGCoDtszj3/uZ3RrK1QfX+E7MSEbO7+K
e3YZ7X48QQFjAYN3Ny34zn4FXtd4Bt37ALck/6SDLlnRntkRwSJwaXGI2lXoqP5alb46OZjOfPfd
eWRujSAf+9HoWGXeSyxra2/tWai8XjInOCGexJtDZXncFxHn+1u33vxAw6WmMJ7xee4d2nyZ1IHA
7Ak0Z1dWvploBuo2sUbmCQn9sgPcxc1Bgz7XarPgX12YH9x7Be+1H71RRhZk4B4CAbOw/CmFv33u
dkT+xebbbOhw4Rk+PNykmiMPZpY4bnYcwywrdiH5g4Byu/W1Bemsf+TGcZv3kZd3P6vr82j66byE
dy9ZxjNug64VsQ+lVFw0RptW7/VMmU8cqdtFZlXOo+o5eKUUf19z616OutrZ101V6pv9nRq2VPU3
L1h5d9Hn3MIbi9bB7R4rzjd1JBcuWuF0JNlMc8ZyXICxlrRe7cYLhn6KWexLFS00xWVZxeeO/yhX
DaRY7H9FjfXwd7kEf2S0LFdLQAR5wfNA/WlGdgN7jZj5t0xwL6KtFHzBVpR+MIQGWXv/Dsbi1EMu
qi/6R5vD9LnAPiwmmr6YWTgrp0wgzHMd0RFB8fSxpbcYmGhvQhjvGzP6r2U1cgDlRObMDZp7P4g9
d93oalyAxC6mf6VanWRGDUnliW0GlZxYZ0LSS1Mwgw0390r16wkZr6oHEEdYGgVfqE+3stKpLJP7
H/GK3hnZS/zcOTAYSN0Y/hBYe9uIT5cfXPDeeDlVDbCtWRNR0XbFCFT8EoU9STTsr9h72dUTxsIF
hKWKWEDI6Kli35vspkrb61BYO4IowUtem3LYg851QiwZCM82WJdRykDER/Wl9Nf8TXo0v4p0QP09
0AAGhlpqLFTXV6TUXw+NXaFb/+lyQD9K1JeZ2CNvfq5vTMMCyTGgEhaizRoeujH0wfTO6qZH8q+0
bLeYwUprznApqRtD3qjJmZU9EGkpYuhgokLMw3iqz3AqTDqnW9sgW8oIlLmTmyTMqcAqECqHB7VP
u2XVYCR+s1GYcZwhPTI/zqX+/jsddmuU3BJQ7WryeNlOf4apfeHvWqS1AULHL8mClduzzNjYxnUt
JsP8e132dm320hGlx7pNBeWnBn2+lrdus3oPiJvXywUpfoi6XwHEajS2w04bgGMkPEgsYlE/qNdb
zup7z1xfPj71RTE71yf/q4ewxf+7qYEB8Qiqct8JO9Y21S7ZqsZ6TVBh1Y6xm9iLkHh4GThyqwD5
j65yVipbFHPaXn5DtGrFsF2C7g6wdnT+jwHodalpzSzkoCw6gLZyF9MGE+oHONYW6JSAxpSPKQc3
ARegGtySGKuod5h3kcB3PpnILOnIjEsXWT5zfOdlKbfw1QSRkp+XVjEmGGnxPW1icCkGO1IvEFpT
zJ2xucv0tjqdz/WVSPPW0pm/coJQnWbusKGD1rIvoQXLYTnlmXn8BsWv1vvwwxNompsVPvcs+yW2
/PrLHX9t9zpGUeTsHaEvuk1edS3lrWoR84hM7RCo0VfdAbRAEhFXavQT+BArCI6m+qudLHuziB2+
SpZLCSufwY3RRF3GUxYjJQ/80zSzBLaT+javaHgapxaCzoJHG61vBCCNK/wZUvIDFN1oHrnm3gac
0GbBcrFaXJhkaTzQ+2vL232i95uvnc+UVcidIX/Daue9Au2sXAgVqhI/54E34xk9Tiab7JAkIC72
f79KZWGs3YgCAU/OI3F6cJy/3rK3Lf4D21Ec1vFrRzKD98XUHoZBAhu24wmdS7DyTSG/dPExq0Vk
U8zlXeZ39AT6I3t07A+TuT3mri/NwFYkLRh9gEfrXk3TaUacKydCmJ7TAI7jtBPdwqltJjiLJ/Kd
etrtKeewswARt1o89f8tRJU54YlHjZHBHpQ7UFZPpK7vhpxGOh1CZmRwVpPsEQHWmaH2CHNJ445C
K2WBmry8zUKtt9iDC7HzDpUMj+4uvQAwX97DoJEU8AMmO/ereMv2afZ/KNMnRU3W8k64/Flcj5AE
/Lo0RySRcu5uXt+H2ZCoYA8K9lqGNZuNFJxXGfn6Sx1xSwNJGlKzQNBs90dJKbkZz179QIbv72aB
M3xdURlRH4h7raWbTrO6mRwlnmAcXzEkjamWjy++VODMN4BtAyioxVldwT7gFWzyav5v0Do4G5tW
G5aNZlN62gOKWOaye5330jFjrdcn+/8/N02SK9S0K9BzJBiZZD/n420Lq/vGbnVIV6DqYy4WSs8P
NSRhoXghmdFftX61e31wJhsIQ8L+gvZ7Wu6uCQkcpfs6b6zVLCUkhaVAkT/X22hQ5MSHc9mNjWIt
KqKV9qoeL4of+6uXo8zkEz4TPYsJPrCgIVX7KrXBtFiLOqZePfV36YoZYe4/M74DX0DuzQdqUbru
ns4+2i4VWz8wTIDTNusZnRIEYiQpvYyggmmVbxm/xxUyWwqSms4wlta/wW/vItQV2wUJ4WVg2beW
yOCVObVHtG5AyRzyzCEpzAWMBzRG+X2Zi4fZbzMGMwVyDa8chf0w4AiEpIHfB1Kks3AnsjMiswlU
kRpHmP2S/d/ehSs/ypfsGTQnOXfXBTsISyrPIFPbkhoyAqWbWbOhBwDBREIjZRG0fnzuIgdcRne9
3jCj0FoL3cHm4zxkuKRb4aut+Jr79E1ZKtOqwJgfVoBByi8e4dMx/lJivrM+pMXzXcvlIQi8ldlK
UDdA4hVGG8Tx29V8xghm8A+WnmMxDZ0/JEolptyMiFqX5nPugYSpm6NwCFqLhjgNE7vkj9pOHdqP
o/6TsZb7MDuJka+krBtfcNZHGRCOKD/6vBfCQzdkwafn3fh5moALkuGUNJ8hzzzMp9b0AjPtdgSj
ZfEGLdkloUQsfnFozf2NpKyO6fOVDJaZzvXHbmwITMxqMXN+3HqMQ/ZQZMjD4S86aoz3XjfGcM9Y
fLr1ggwsvVKIVQCg69WVFIQ9fT+gDnE0IIEWZ7SXRaPKKU6z5XXG0BrhJRJG/LmrKrVoMALSnxl+
b9p60bunnZfHx4jbJfxZJfBNuWi49pCUfaSTE3i3Cju1nKb18umAmh/fGc0x44pIist+RMz94NX0
N0QZi5UMf+A2ZIywB5UWvUk9c8ZdvL0F4OuYMYHlPbQEzgFsBRCHQNuCi1afQEiz6oHq5YLpc0Yx
tAPtT/KBPxWqVDGrQj1ck/4EGa9h95oa+4xvEzqcxd29JSuw9/oNvEw4SO9QNgCJgTQO1W0j9sRl
wUKTxa1XUTLxw25feBZ+U7cAtgWlMLpLRjtemXDWN3h4rs78XvvLD7c2G1dI8P16XbkY5gpFGLXa
0PomNRDnCF59Q+D2U84Rc4tr/q79jefkAzyy/LELqZXpFYSsMdXxmAmTQp0Bb8+MnZv8TXMGYPaQ
ol3pmG/somjVxR0+GkmQKoGVSJ7pjRknq0fS8MMwTPnGSjRlWaPh273NN1yiCquov0FD+r7GUg2a
Mp0i9U0kHnpj9edAnv4Mb/MqxdvHtiBvrfhALeFY3fhblrIiuRi069oURnFMocifbT9fAhKoT4On
4fUy7h2E8vtZezyI1eH1H/BTwSURVQWsZqe/Nb5FaAMCl3rNyfnYZk7moV1DauLu3Y+44gPz7FRx
xI+O9YLVQ1M3utH/eIEPqV9ApmuiAx21axAYb/399ZBWcyC1VJemxCWDDpuwwxMQdj8j+zV/Vdd8
ABf9b+QGfjF0DEkh/4ujWLsKTibGOoRJFtOWXiDg8UvWYScultxzTTAUsRIgCT9uA/hB47ptFPKB
Nj35yD5D8XIO//odurXN77R1gwSrm+B8rqo4H/Ww5q/rnyO7g4OUgCvKrjru5ptMuV/yJB6LiSn6
aAntVWq9EDKqGCfuUpiYMd+c/YbiMzaSdy+bWugpRmZZwgltjBGDDmT2tSOkl7XKj6sCyXKFa63E
B5luDWr/5BW56GM6DiuWpZSUaH2m1eU6TahgNBc+eA+IK0l/ZvYJ1KqLzuCRCZDcZ2e74tShitHb
/uWDxq/lD66SsPIIKPVUvyju8F76mv1eCfHCJFjOXefiz1V5DUwlCRChOqNZ+BSk3gFa6qxzUkCG
hhPfJaXj2r9y20+MG3/15eoYUJJtYBnE85KKCglq9sH4FQkNOumMdTv4/ppzJ9CutZOilijhNPoK
lyz4PhJVhhg/BJbL/6VUy10QXrQwNJUHsnEkbBGklK5stQENju65WMPMpzafwcpYuDgBKXmgUZds
NKK9kJe3yJK7dc0ebC4ne6xzOH+2u7d6z5HV7CMKx0kMVX26qbKt/qcfJHp30ghBSQ2r6jvXxSMk
DK0RQ3qKaX8YVtSd0m0+warq7WIGt4MTxSDAh/ELxG1bueIK1feA9/XQXZOMYvYgslPxDq3lvq/C
VUePLcM4q6yZbomGpQMV32UXspVCHfeto4pUrjclXMqgtF39opLw2z5viQJex3HzZC+4a/UUnULL
s0VxrL4HKdf40cGbfj/i89Du/EgWOGp1fhNKsvjNJm6tHTU8SGzSxRbLK+hLKOdI/raWth38jhxZ
OWwSqnXiQ5e405oN5ZcvYi35NGkgH2MVj2EUNd/ll51+mVESV5Mo6nrHUDwUz0Z6v11ROnjxWQ4a
1hyGAh41/zQnZItnApGZP+MUev6EsJWbES+cSbtOdNmY3TMcPECsMfoZa++ip5usT0Cs9eYJ1hN7
daaIHAPuc1TI4P3ZiW9K6wzlDHyVvr3mHYaudcl617WNyLFpgUjDibWFgoO+EiQkltE52lHDhVDQ
v9ID+RBcPD7wdREIwCRyPoitHunq6wqHVUl51mrRoYQJz28jCprEPKMxWWZNfVoFhNiQETbJRE+2
0pYDB977RG2ZWqI97jXPWi+Fq3Idhqn+agMlSNFfG+D2ppoEoOkRwUeUnt1QowtRWlzfmonlbUlI
aRUSyLSLM8WfhVT75wLvQ18K19mFVN20CiENJqrqX/v6UVAz6niGMrtKIVP9X6oF6fQlruw5qwXN
jLAS67qUkmqGnF2kbZnK3FGzdwlczrygcap5eeDQGn5wm0733a2ANgCFI9HGiFJck9UeOI9cYavF
URgdhYdDVouQSlUGI49WTtC873NHZZ8LAI2cW64rxQn8k5gEY9uAaBw9CnRQMuo+WOqwA8JNvvGV
8Wt8ZET7o0gs8Wq/1/p0VAfpyUeZU1bDu5dckGKaNtskAzHto43H/mVXyeToMg4rzTD6di+ST1zm
AUGiZRD2MQiVb9NRKaiIIS4jaezzKt2tegVsc187w+ES6zyMCdr7kpwbK8TMQPAHyCPmRizOjQFa
sx/Laay6ZdNeVUqvFg7GtS6KP5Y692PFaTgrsDGrav2gAH4DMiWsU/QaVgmYD78/s91xbzsT5cM0
HqD0kfqKdBe7Y0R/C0GgzMonHJVtAcK4E91PoJyg90CewIM+K/PtnrRenQWNMIk9cFcDv0Iiwyij
wJLfMnmNrnAHuc7ERSqo2Uqrf3A6ZkTWXgTSnbbEXpcZWIeoEuIRb2h9IeE6l1EA1Stke41oTmw/
OmG12+t7rvogtOjcJe8ohFgDpQOml1tAr+qh0cLF0uGNl9SkbFF4kaZzwkZ39B+277LDOLT1LhR0
0Hw9JI6oKQeYJjWI5Yxh04Mq0Fueg3OnQt5nukv5jSgetlVTAjmWS8K6V0vq3FWjzOpKv3bwx6MA
HyF/UkIJ1AYEwE1/EagDBP70/djxT5ANgkBJ5UdhQvAwtjw0XK+yGhVk2iWwT0I6A+0uTWhRoa6k
o+kGVNF/LVo7W9g/y3QMa31BcPl/WNv0ZxwDhEA30d6x37YnhzvKAOmg3LUoEpJuIVdp5Ud0PisA
tw9MfBxU8Zoj1nYk/ri5/jeyOAgJJ82jxoPjdygomudzRGulFtkL44U0AXXtBLqWTXayiS3t/GPH
xX/72BGCjXppAtsa2158Re7S0/AJBMvwu0i6i6i5Z7xJil/zZSgzLCG1V1DHbO87O/7dKEsa3RkN
7DMviBcfp2U0wR1coaBomC6MTjHonKl42PaU8qoxfYlOiNkbbBWGn80pwOoxohrep0WXWIUKVgca
R/P5ExVdfMxRR33+cPDRC8BfGqZfCmPk3+DGkH8NLdEjb+hcyjCUtkF7CSdRyAV8F1ihDR7nkJwC
xNmCzYvxXKQMXxaFZ3Cz0vkd3miZwqcR8kfAtGDrzbCecZOEm9+a1OARde+KcNcA3oU0IDi8OTsC
rVklE460k6fvo7XWiYQ2cyOX3LPhFn/JEXoA9Km0bM9VTLh/SOJA+di0dcBJQkam/qiFmgUkiUeP
fjcpwga+wlZetkmSOGNp1EiPVXPQN7lV6kCc+fvFfguaDSE+7aTYdV2wHXL6o96VUq7RPZueoTS3
QDHR/TQvgCZjElUu06zUT5pLCzRg0+J954/3zXaqI7bq99J6VG7bFdd0xUmAnmHFD8dby3J2N8Eh
GOZMFjtdWFV3Cko0ozfrw0ZKLtiF3bNt0rr8Vgk4xzAme4BHYAiRF3Y3tx9e5qmgJCYy/8i8iMJR
cyKb22UZRmeE5PqI2XNDC0jZV3jBof9fMTieBhB5yEV3jn/fBQYXDGoFO/OGxLA4LaxCCtUsue5L
kflgiThur0t8xQxP+olRcaTs3h8TvOqj4244DnxDDP3+KUatuNG60Qn0EvX28Kxbr4GIKFjY/rGr
ViT0Wgsdu1ZlllzKg4dkIuF4Cu0KsyU9/iNUWjDaiepK5oB9RIP77LGwWjMovjsqLrFRjLmlk+hd
rZlSWIb76eEcbVITBBgnUogG7BbaHcixkxXcy8C4WeB38DNJFz5xmaI10glpLsTo+a3qnHYflcm5
RmWVGmCDb2daPe7nDTDLkej/FCFpmcCX2K06p9w9mb3QgB5GLmFjk6nTUeSL5qCkvEt6dso6x0WJ
eMMifIwffRnx9rKGPmE0G1WmvTHIJteptCmKLcB+Nd1f1dtlAJvxgwOiBsZ5BoM52YxS481eP2xu
7CAhESUr46m5xlD4JtOn6ZIXjeFDvqpH09JUrLxdZmBLIgtOTIrapKY0VZl3t/iRQ8NVdaDYTaNu
Cj+HQJ+8h/REVfCsg69pETNTLC2og+bEql0nGoWVCmfkq0Yqd9T49XpqAzFSvGJxne/lJ1uNhvA9
pebessQ8kIXzNGYEGgnKq5oihp98StsNYdnRMdVUgQJL9xM7FYvmTdU2QMOV8h4y2AJk2CTfo79i
3sgoFKqVNN17/QMpGeMA3ciR+EZIft/3z4H2NjHTjkILUuNoyFdbPODdqIrY7DWxIG7kkfC2kcB+
11sOtV+bWWdOSsA4VlawhSnBmgSn3NkhMTPJMKgaok963hK53gfD2RdMwrnBN4Bq48tW//LW6xlJ
jHGftug+tF262ZcSY2PKupl/+7geebVFZ9b0xvpWfu5WyNXyNsUDhbAv4ff+dH1BYmflR2cCt0S6
+W/bRuAv9H7f5PPsKkQVmDHdzESmSPm6+KPniIAmXI0xP0rZQS3R2CtSwlXmgC6GUJOjCAFTxY5w
HXmWYN55sERwJCjdeZ0EVyxfjl+EUvht7+UB81r1X3uH/YTmMIqDzOBohwQZWm2uR/9dUNx4MEIA
kHIRoXRS+TuFYMnH+JE456HPIpWQYpCp8enh/r/gFOtcp0NJmjA727EnvTbgxCNp31E7rQsD5ZPE
HjDJ9aRnfQFoWSZFTaImgub6aZafa0X5lkOSy6DBPy9pEX+HJeef0iFhBBcUBx7u4n4cbe5D3bsa
1enUOc829EW6plEy0kv0XAhGQ/gl9TcJKJasMC8TCVagpxM2Phe9+RozzpsoK008sga2msFoM53n
yVxQMnVZrrp+6+S24Rl0FpNzIeDAzFsG7lbg/mLtVOTjKT1bnxD+LQ9DljwaXMa3N87cxexPplY3
VHLX5CR8ofqG5LKEANs81y5+Sn5vIeUr3cp9/ig+i6ix6393vYa7Xrybti/RToaYW5neyGdLXoNV
USOZlhFgXymb6+ftlbpPDmKdl1deDTNSiiC28zze1m6XZ4S3SP6/2aQPERPZKRUnJqtZYLeWD5kz
wjtkBs+zEConBRfZeZgO/cG4gNiMyxziSp51pm7wT7V1W/UOkeHVADHJZ8Bnxpfb/P1Q/MNR6vz1
SCzW9HxsaLFK2WI/usVxxcxXrTJTOooDUxIHzbpy7A83WmVFb+PdAkJlqRTCe0Ga2CReh/mdSSn3
n8wSjvI/NsSlZevZ5Eacp0LNsIhP82H10WqhnbMryflW+ik2mrpnL6SayZYq9iUdy47Zermh43Sm
LLFPcbiI3Hzfb1XimnkMEOtuDbwEqJwc1YdEKN2uW71bmcRE70jJ0+x4Gp9TYOyJVmf6xlTOZhJG
wnoixv/ZV00C10G2QfDaJZsUExxbl++b6KC2wWKVTPSkUJKg06czrhA8obEuZQNv98qG2FhKs2F8
OGldU1JSjO1lAnTW+fnU3T8xOV33nAWl4VanY85UzufJNeEUUA4TVh1YSjGCZPnrsZ+8c4kVZ1Hk
BcaIK2A4URhlV5wH40sRLqAbv8rzaKjwDeccKoesj5NHBilypn4z3IizGSDqSSeXl3gKQsXwtixm
2BMusJJx21vFOloDO7rSvX36zPxpWYaE0XNfafKa1wd1Xqsh6d4pn7FwOLJQQsIKIh2qC4pddagy
PoDkKC2/Pi0fAJPFKiXNXcroEQMXP6iQZZOB79b97BZCXSEKlVlazLsbzPoLTrFX70A8QBGGOrXC
9L0x1vx7BiAkiV+8hnSwnrtowwvwPswZLcMPFyYGdVD7acvqEzW+3yaFeRgCi2sJ65oZEOapTQMN
te52u8ZjyOZH8INhzjMc2Ex93QfawlpVKl2wcZYHiyziV/damwkiLxdEuGCWeaQYqtgCPWn5B5nw
chrOmK7qffPNNDJYeM0AP0LK7QXqd1opSb+g/sV3jfMG3AL3jmM5IC/M3mJISwNLsg+b9DGsyAMl
kiZrs7N+ntQdII44XQe6Zk6Sb3AQscurrrXgQsoQXjQHCkORFs7ximriGzxTFywWu0NBykjs00kt
LDdW5jv3liAnWZPjdp0OkM4m/rPMQwW9HRmWmydAonCc2vTq6JCKrhMyLEQr/NrnoQ+l7LovmBkd
bJtVBG929cG01XPBzODjm6pqAJWx27/3ugOU8qenicG6B/Qq04PR7YzbjNIMJB5VZyMrQaM48Pdh
/8HtbW3t0I8Dxk/QznUIGnRUx18x+K/JUI4xkhr2RZKPwTLn+a+PVxNVRgstQ5ZqEWlVivU9ItCy
qREAZCSRZ4fSxckpj6ODFIhBzUKKyFaAlEjkBhE+78f0md+kgnH3wfTKoMoHkvG8XzBG3WMh1IVe
noRRPa3ZFuxfcF3U6GaIUARjKGtyZIvvd2XHq+W7rJ7DEaBPBF0zILJmW7UhszGSrIuslIy+H7Y7
6+QXdyvfrr91lAsthzgMrLTEx/0aGmCNda35ZthDRtqBbE3BZgvh9j7yITRegYPas9fA19Ah1rbU
yHafIQmDmOwF8RSRbku+JIZCQWITY2OhXusamTdpupfuCwjnULAhIcSzC3HidWgUCCLqYdinwDbJ
euBlGC5WHt2Xc+fx1FwXZZ80OKbYlQCEgTjeeg4oh4CAw4gnN7KEGzqgI2Vrt0K6evmZc40zAZrC
BzG4rKHUa9PJ2YVAFZRv8tlb21/w/YhMMVe/BuVEPBxhN8yobERg2nDdjDG8dgMbpZ3/UaZUqgtM
K1YKyekxXyN39LFgRaZLaTaUNO2ufETB1DZXQKyzV4ot4ADX4MGwm1+FKHp6LVZstHDcJIJlRW6J
cOoHlXhVcZd3zbDzKQuBniyG/3cLFEPCoep1XthdxZBg1nUfUjmUazoYo091T7mFDEgq2tVx6rYA
XS9TWN0wbGKiSOqb/KWDj8L8YgDf313jefRMh+vUQbHsMtx/JmmroqdZNE+7ZNFuxg8CR9CsT4we
14TnnZlkbEYcSFEgD2sjEK1vrTYu7878MLYTGrbpzfzmr1SrVihpWlI1Fv06rEaQOyuOBMnixsHX
rJQcA7IogFvgzsaBnPQAn2weGNdyC7cHoX5YDPc/m03PsmdDE7czMCc18s0Ey3Is9PIJzjo2XJee
NPRS1z9MLz4TTtXwf6CMUmPdurMuM5QX6KwsjIm6+2yRZ0zJCl0VQCMTTbBABdVx3eC0j+y1Dyje
2B5s8IB1yNE9FCPIg58SdAB7y+2sqJ8lY3TQnE2Rq9dBWJ3r6Wsvq/tC5iZmmkT9QU+b4LbgLp7C
bsd7sQ4+prf43ohe5y6QJan+59EVywkC2Ns+PMMWH2Sc8SVTWW6hPqkuinPsuwzIRbFiNERJMEbh
frgBZz3/mtiV/+Uy3+x2frwI5RjMvSd5YTeSE6TFFpghK5es3ktFMOXFrNkZdTjJ23DHMOdCivBh
RVa0/PN6nEhZMqxu6x8NvMfPs5MY1aQXPEkiU1A2gnEZqpGsG4R+1Pfk3fSD9B7+5YyHQhFIvkrU
UaifsutNhaYKHvhytKtZTsTsWOnLz0sa3vLd5+WjaGpIXf/AEWyQoH3lm0UW/4hV4KbTYxbkngij
XKBNFeRiUEsiJJ2qM9w3JdiMiqKDWowy+jsfNbCbH0tmyzc3n7gUiyhLXaeljD0oRgxNnP9/m/+g
urmUoqSHWDhrODlEoCT2JTkf5by4A94mWcTo+pr+8Iau2cI9bzd5Q+zLRnvX1sedZBonPZyNtQS3
EOvE/t9boxuTyurSN76XUf9IdAy7QuKC8v8LQRLpV+Oj/lxDxtCvEGq0tvmnFb4Rj+oKifyw350s
PpvGL1gywrxZXd4r5m72f+0128h6GO3IOQJINUFCEXaBdYPnbAy9ts2BRM7LqZjp0R5AH2vE97Rs
Is9GEwo/bXt0hrMv3Q8R6bAsYmcvhPNLbk4wkInasOSNDSBL2jW1wWxKESXpQAUHnN4OqxTGzOqk
NMVBQ110Wo4W9/NENjJFHxZbZLvXD/4Rv9dZJdPJlgqIIst5xIL/chTsRnAP0sJ/TEFhW6Z3UvTU
aPyQW1aWdd82fvjqr6cb4qqLhyJKv/9Pv6FmQdT/+7wZh+G7lW0Pem4Vz4qNxEK411LXJGDyD1rU
PYhS9+aZEF9QHSJGm+4W9efWW8PWabZbd2ISa10mLn5+lVsyl2lpp2lhQac+YBvv7YeF+2pYZBWY
v1z6tFH9uZ3gFSMT8TQuWOvvaUaVNGAaeY74ASE55zX1UvAmoBK7U6N8wMTrxxGfn3QJY1sIYCky
wKDrecd5SlNgVj27m4SGSMl5ThPmBqRDVwJ97TJMhDv2u8TmEIjPz3O0fUiGvFj9jo0YkN1ukuCj
FzHtRM5vTJN4KjHCql0hklG6+RFQkTddt+bFpM1UBgV3k1sNkmV4F4vZDzOHBR0W50qWNtW5M2+k
6t+D/dJOToNmbzv/h85I71g3vMsdF6DowdAcRr2OcK3bq6zXktnOTAot/fagpQpTJa3UcuI94oDn
ZWjZgp7ThT7PK9TtTlLSwVSDES4Wa8N5fCClOC3xa9ewjIX5tiipu2/2eOjxEwgWL9QkgHWwdqFl
SGke6crO24CKdO1AraaRRTydf4byJ9Qsf1+bFDIfmR49Q7i1IYf6oKsaxapZkC4Aubur8f/tPo1f
3FUKBNBla10fzTvn1sfpTjhTiRsyv+E4jTklAxIHjQVKqxSEs5SWTnNZOCZ1f4+WNgXo6XvrIv+K
iT3ad0ge5DrG7Iw7+m3ZsDTrP+vWAywWX6srHpoeHwlW7cTikX137nmD1DkK4by80qFLBXQe7UFv
AUWEanX1REUPMKCuSNbrui5MFYp24et2bGNZruwXJJ2dzKV5E+izt1+itdOmDgJrYzsXcqUhBe9a
SJK3sb4Tw5W1vSEebZxvkoi4zm0ATIamZRb1hWs2Vgiy6VhIYcYiAWWjYh/OJgWevkcAB4EcewBc
a4pjhHuLN6XOuol+OLTeZhNK8AH533yYoGFBl7M03ExTirugpOZr2LHYsi9cxWQX9DVRZMm3t1R+
9QAyAIFPpLYeKGdf8W/WLSQMrTaQvepdMAXy8x8cz97dcFm7m245rfxqzpFbRzvPsphT/8xGiEt2
sQ7Gn1gfZ4QX5G5Eu8lhw75/uP+JGb1FawpomGsctNgo+SqV9bfJAFPnUFfKXhufrJJkAREirDQa
9lXAtQaT7sCE6AetF+nZEnFMLmzpFlSPJRayyj3lle6VV9MDS7P7sPGrKZPiCOCiv4aThjj4rPDB
x/7+pYCzZlOniG7/wlp1dsj2zrJ2Ucy1uRSvYPdoxisseXYibJ5OUUrI8IhpkbXSaj2usndb883K
xT/tm5Kw5LVxq+CJyZjPVimCt78WZ5z5CfDWdIigSztFOles5DrX6A9CZAzPynJdTXHnlgJ8zlzY
N7TMSKtTlN+sxy3gdwheIzUQWtdiNJXe2F1sz8FKIW2JqiDCFLnra6MDVsc2IFHAByEUkoN0sr8P
WEyhJrb2o073ru9EVQuuu+kVDMZaBIgYsr3H10pVVWjLY2XEP1Eenxr1jCE3ZeoC7kSowPI49Eli
26m7q/cuwUrwiXjPd/DULcYbz+iqpo8TZlG+/DAmWP2jGj7o01tYCD2tZu/L6wVFxhaF9zqrH5R2
ELmsVBOvrK6cDp9nix2UkWkG63WSlG2sRIqRu3fxl0z+n3qh+9bHurt6Cv9CwRdxjt/mWwEC/64x
Acl02AMxZqLG4XXhL97bltNgMoIQLeBw4coVfw64Eit6wV+VWeISenNHxdtglwoRIX4BanIrL0KG
yBZpj4rC8++DpXH3Jz+LPXEX7/w2DqNFEoWWN9ppiojZVXI1c5VAL3CHQdVoeD6kUDU0678hiWnt
4HqZkbh/h5i0L1658E+Siij9Hcl0laX/Dbn2wbzwYgmT+K2vyKEz9DmVX0PYShr0btLnrQqZdmLv
IrmIkiTvSu4BuFJs+rWgZhvnH8y0wcf9BkmNbjnLoXUO8NsoMf+b143avXyJl+Syh+jzZyNt80S0
OKwLyFijj5WXMfN+r4g/8v865+93YmdueRnNGV13Ib5a2NEbsONovIjsIEYo3PPllasdo65UqyTn
8G1V0a0u+IQzbg9KpXPd9ZXjSvJKTEg6qPhuN10PYibvPXyvPvD61UwkPB+CEEqFptQf57wM5kEt
fQ7/43iG4GMp/3MG53gRgQ9TURP5wJLXifLYQCs4aO5AFGewfJ9OG36PIvBgJKtOWzrONzkVw56a
PavxktCKoh4yeGZfAwE4M3z9ughHuZIOY418qtNOEfbc1/EOz1XMKd+JKLt7BaBOAO0MxHVZP2H9
8U60G2U1Ygt41iVTFuTFQItEqnMy+uAfWZDbULWF/hufRFItO4PjFAnSE67G2vdCFaqhhmmWDgdg
hxcCSr4aZ1JPVyWbQ8hXGI9sNZki2J9RNgzDDLjkkfDQOrIA2dmq/ofQeDm7btLAWUFY8dWd4vkF
SowXY5svpkhO3mdVTfl/Y9FHtMkxBSWvLzx56jtkDamAl1W86zitcLc1QsBkhR4+V8eWvR4uOI3h
QVUxUqewRQ2XAz7gJ32FSb+EHV0cMx6RRhWpUHOfy5C9w03HBVK3NRIk5+9cWq+CRdWc3C06Fza6
DdgiJKfpM6DLUoxyvSF4Vj2WfLumKX40ddKHmjZcIcQetXLm7sKobDd8CWYhjgxXbThDEpbZ3dEx
iQis18oRHbCnP17PLAElzG5jNJlrly0hB8vsU1Nu2Nj0rdqwNT1VX0TYBq7LICntOSxjWblkxKER
TABcD4xe3Ro7hrmfDHymwxBi539Q2cu/2WW+u+okFgSVMRC/hvNXUrnEBjwuO5Ag58Y0XgQXFAvr
1RzTZQ2g9Ho+bNH0KKMaBdmMWOq7EQBX95tHtkOKx3VZR/4RipHOZ1NdLI6YRLF8stq+Qkj8vhs1
ayIF5R2cKX4u7QatwVln15o0JnTC83x6yl6iV+2OAwigiPHA7aRWxUxv/nUA4ZizRXa+RHNKXic5
uvsc+BoRe8T+FAcJjxQWmeWZZhoV9DSPrPOL2fXdxEG+09ZS8rPZ49mQuM3xJ+dEWdg37+xIGa3p
opjFWgvq1p+HAt4NmZAzxA/6pbfJDg3U86jnS3XkRMaIMa5ilP54AwpTcDdjqMynUTm7NNficBm7
UCf3JuXNLP5cw8SfucSqEZP6G5NcKAQQagwrBOu7asWeBi7de6c/2ToR9SogbCR1jWj7eGVxZgl5
tZxil4s+DEqpGS3Pa5jcPv5mBvXwJj/k0V+UbO+VO+2Kpua3oiOUUNd6aJJMlsD+0VMcn3oPFDJ2
8rl5ra+WdlT2uYMI98snED7m0S1DK5iLQoWr4J9MsACL4X5D69725oDdvoIwgLxvdInxotSBaLDe
8IjAgPnnX67K7cYWnmZXD77qt4BC9sy/Lf/LQ5JKEU1N/JSfPiy24htwoKXtVI2tfxfWz/h/xE0B
BQobezT8XJcAVWqd4tDsb/bUkeM2rfXjVUoYM8dQP1Nk3ubaoOC8wSoGsZlYl9DFx9oX/BriB7pA
PfunSZl1eXjJM+jBpk3f+dv2S4XzzgOAKUuo4y4wiScP7DhGj1BnMvp2GCTPLQLQujPTTashDKhd
NXY0BpwXSnRBYnXI7x0Xj1vIk/kmm6cO8BKY4Jw6Wma9eMOMhRmnW4au5XiaeVf82G9a/Td3q8gG
/wXyaWHa3o5+kJOFt/2b1P03nPgkik2zDTrZsjcWn+OH6bkMsbIBtYtNYrQIJbaQFgVVGsZJZHA/
LiCZU5NFQwKzq0j6gpBf8oVPY6CqsQXRZJ0oyU9ZwcCfZJNVtpQ2BojUc1x2TYtEpWsVsi7U2dqK
5IjvV+7sdxYuXuYwWzubb+Eb493gMW9Hfxg95EO00RREodhVRDS7/9aX0TgQ9DTLnJQsWJ99twMR
HmlUdQtTlHEkXbofrrrlw0TEZ1sZJEnqI2xESXkK0UQ9bW4EdvNYDsXtqca5UkuSl86+5IlRBbKP
PttK+OUT9UyMSCvGpB01PpQSXtHeh1IKi6nD9P/NdorVvp7EdpPbHPtRoCA4sLToD8dsUm1/ax5q
OH320nizF9BGx9FYvmDlgBzKsxWWBzl3Vf6Q/wvxQGujRz/iDHICCU6mgSQx0Q50zl87gD+Tm4XO
0OsvmAbJKSlKWJJ4B7zmHeAuOXNkX9YQf+fRqTIIdf3FEcbkCpKIwCjCAJQBe/5Yn1gmhJbQbv9+
jltfxDwy2Sbr2zw2WSV2m/zMMZLaM3dlCIVKtpIxdfHwu8zHE6EciUYIuVguVUqYp79oElvTfk4X
hmpHtdOatebdCPZPtd13ycZklvFke2XsVfYPvM68XHkuBX9MeUv+PZfe1Kw9E5vbpWMK7DAlUL+B
AAZ8lu1I3pwRKxtt61A+WgxV+QMNioEsnT1TykxVlGRfIsG3m+R7txNP14vV16efD4NlVA4v2JyA
5p8w4imFxd7i6MV6c2gQDY8+sGDTIb8EYHj6a7eTuww6vJuGPy+HbtARtVc7Yag3UbKOwz2eGf4R
wwb9vNH6xvjJLiN/tGt/aRrtZjhScKR3AOQBM7PHOYbUpT9AP1NzQ+lr6wt2kDbW0rF1HvTYKUeK
/0PyM7tY7u0YKWpCCMMiIBWaxewRfOM+vn/QqDbmcWNKIXm5OghgsIVLwH3yHcDsJspqE4pWXCG4
FY13i4XAh3XR8SpLx4lZmRu7id6j6odebyEhqmTdDsFT77zSRa1YGbagQoNGpLGBdhkM1Am0MueW
596yWMYl0QXJ8USIQdG7/mlrlV2/fZvpH9UHsfMQ/+URjPKlptDCaBEctqcHXzL/y+RWqKFXc9WD
MBBV6541fpyjqCd7sts9tI+xb9wI9w0XwFjJDI6SYw8c6a+Nn+ThriCNTj069QZpEmav9B6qKaoy
8JtzLgGITK7fSf913cLLqD5eT2NbPM00Pd6sfidsEFXwRxKaF5PrOmrH/snb9KaONi9njjfEVVPO
dfQTNAHXAH/yS8uIMEiRCK6qNNksrjHTU+PRyt95NmwkQrSJ4p4ChVN4ARYMwENupljcuO5QgcdJ
Rv97hxijw855DuK3dxJbum5Ey+c3vv6EhN2sxCOwSnHEwmugpxGuv4IUvx6MdZP/a8atgiVnAX8N
bXtMCaAEul9OjEYPJosxgsxWluX2m6NaoPqD2etOKQHA7DPwwg4+oNvDpJ52e4kXCpwU4go8CLqW
BanwrR0fCDLnfhFwtVDG5h9YGZfuUR23BA980zk2y4YfDW2j0OSgXhz8kLxx7ZecEdWW7DgSEt5F
YpgSzg1FJNQwrz1OJhOqYoRojrcn+y1gu8+22Mv/gXY6Fimv4hdrplPc/Uaq8FS/8ahYIj2b4udM
EWFLRLyc5huvnZZHNZA9uB/3arA4nxwCADlXDlq8/GwvsgxmXlv/p6mvjalrbuPyNMfyZz72/5rI
9T2xnB2YpeIit5vHQG4ZnM2B6i0ZQMKMRM+a0P1Im+bKF8IH6NyJldAvJ9OTlJfC5VlTSN5ejLzR
+YIaHjLdlRfzw00AASdk8WRddFghyJuJmQ6lGjINQ4C10wk1h8Dgsyt7QX4OA+VnCGdhwsuS9hL0
lN8Dc1zTFinMguQ8Ys6Okfyash4hbMvmT9/bZ2hLbRqCmQzZepT2fbC4C+JLTyioU3CGHToB028H
IAwAzBU8ivMaF3/Uoaa1Z+QjtDGLfsmi0OljPsXRDGaRBNzn1+8UtvfNIyZf5P2yujfaWwtmbqmG
94qXw2KKg5U3LP1eJAD1wdanbFhuU3lwkKLm4/V3RPFgzlHjWPLnVtV0eVixYh7qlSsn47zQk2Lf
moOQjU3FQK1qPHvPldxAYeo81KFDpBUprza/8YFDAjq+iKQnyhuMyN7mMrJrgnezuqK63CoJ9jSP
90gzYlnmYalide5GxFqEsbkoz1oq+14vsgQo7Mhln2N2JcL8DQn/46lRH/FuNKLvBJkP5cRdMyug
d7kwlvqNBei4Otb/jDtV9CxVql47u+nvgaQ2Y64Tr4cL9RGXt3IVVIrZLmPf7AllpVq3m4IsMLfp
Lp8naJsrB9PTy22M745EciK1DzZdzzTNnDrJznoSPhFCcGs09f8MS+uTo/0hsevRQ9BnkzZ7pXla
TL//pQCXrhHbDl5n1uw0DHujXUjuZh2yFniZj37ktUfs5PDvBZILBzIsEnptJ7mLQFwfifNHbUnw
GN+f1I0Wta0PJEBDkdgur4w5pz1T6jVuN/0qSYoFRe4gYIp4E/zb2cZlW7huZG1GG6kCFGVSNsCF
H2YJKcZnH8ZY15KE5x6h7OJ5tizxEqvlaTDmScwNDNcLA2b9lqrdPEUu8gYO+JXifjueibPCug9c
XKgDaMBPFFqTyTOly0HMC5Bvzwbyre4cpindbYFBwnE8dGfxQw1RZZaBSTgrtDuD1B/CdH0OsTpc
EV8HWZmQBzj80rxTR9kCWAQUbIuCR6PR/UWyj2M5XTum0xVdZ8ukaR1lUH9yp/S9yQz+KaHGt8Au
7aKneOoQoBC0ptxVuyBmuhW2n1dq6sPMCdxEBOSSRglXk9qr4bsndtGlgtoEt0t70XCAidY/VH4z
MR2WipV6Mn2SpkUhfujPQjtvOHbfNj3nYXs9BTgr/naaot0B3EwKB+IUJnBAciGFuc6QeNCyhqHa
ounIJeqRwDxeFAsuDRmgXXzdUtltywJWzoycOF6CfBot7LXtfxDJkC8qm7omfT1KA7G6QM7euwzW
rp7r/2RaEWwaS1bbh7YTw3+NBLU3uFuiKNifGII9IHTvLgDWKHqJ/2jzoD9mXjMr68WRgFSsk3Ws
WCE4W4Caype1EPvCLE7RW5k0qgZB482sJTHmKO0gZbmzsRjBRWzzEF11+u/kcOgK2k/FdsXBgVWD
9uEfjmno4VrRzEXiSOktwTdgi4uoWAYB7aOBDcmluHaEpRhwPRRY6mbOzC+JQTmeR0Gyn+SBWTZh
NoO91IQyDLtpWpqXh9cWMj1BR7rFAIgSZD8gbvi4xFZeneDnVN/4xPcyH6QvDCB7ObI9hLQAtIXk
6vF+8BgqHpNq05h3c6h777Pv2K5vFxIkkrJCtBtqnxIv7QUs0qjFYDp2H3XDIUdrQPzmnsC5A6tw
QpIKk/r8jJnxO9pLS9o9aWKOHLAsOzdepB4dIuiWDDLyRqeZpTwW+u+vH0M2Uuj+VhCYgBlx5DD6
CEfuIgPWyBgWPrvm4c4H2L3WqV0JxiNXkbibEyP4GWp8OGxYXMfOTcjT2Lxptx95rSqIFWl37gyU
YMEwig49kSsd59B47IhUWHvP7ItUo48QvIfzp30h9rmkl3j8ObbqwwSqDsx7Tdk9+Qi/gvpUItMS
7w2lNuL1qmEqoIlIrmVM3U46+nyc3kh8uHnt8vYfzX1NvuFls6fFDIj6V9Zb4CyKRFCux3dOPCQl
1vWAQZMXUfMAgJLt1BGzqELy0Q+Y1olgA+/TCPcgVVUpTIjlOvf1vMzRpqRn/rSxzby8gSw8FW6I
emSczb9shGHN4t/FzdP8YL0UoMmTT4pyecZT64/D0AxKYIn+cdqe50PLTe0MLox1v/YpJsXgQRY4
tyVM7oFZcdO2k6smzX/VmLK2lSVcZz5uBb+GyU6lLtYbqLbdspiaGQs0MMjgCzdmEwKrO56twWK/
e2t32FhkKTWN4xYVL9s7c4Y36DAqV3WU5trHiMox1IkBXSnm9jQZI6QMmh3u50UfeNi+V6MobXLs
pXUaGX1c5FiP75IztbPhvboqdQlFjGqoD2wyIoC6++P0j2WNwWErW66GcP/T8jXmVX7GaKkBmPu8
DTJOpXqIPEPTh7HY0C0MIknu5n6nq0qpExJKjwZ2zii5oPjwnSPBGGA8ZXRIeRhCXtdLkhyYklM9
WwuzXcJ6xye4EhESRGxWdn+NclvUp3hTeyRBHiz7g9nvEED8wa/wsdoVlvRUx3PgoylpHLhYf+dA
EwtW6c9rZ0a4G97sbvHD+a2Dq+eSXriMPRyze3UHP639S61Cv+bulHHUWLqi/3Rys8PKFONSzpVY
GIhXduajPlSLqrAKPo40/ZrSd4Y1xA+QUUbr9rnm8OCw+GREPuc4eA7RREbGqaw5wSQxNWeNRXwB
AS5dryZKsIXo2XIwYMSRApinzre28bgAoRRhTxyobiEO8DVovxgE9bmo6Sp5sqcaZxyRBOxTgBFd
R7zfOj29OIdsguECLdhFefUoMnhmgugCN17WTUbDEj87jbDRflE3ICFqhcNi5NcBn/slqv5AuTgd
S9/mpo+Ta7lmPU7DFhrvOokU3ZNRbC87hdZwJ0LQvBFomDtqU4qquIs+DJyZKDlbgIHZjJ7+l/RV
GHsJ9vkYvCqtDwF8h6gzmCRTN47gDpRkROMHc19ZjHWcxQIpNI+eaK/tm9Tm2hKJD4jp6sBUq3iU
ub/1d9xpIeUHTA1iMw1uXjy+AnRRLO8z3Z+xyWQxrIVks7vl6m8WXT88bG3Ex//VtvSelCH1UXa9
ASnvrvcWjnRluSuIZWldsuhKRJ7G80f4gtVMqqQlqrYrVNJtQBYeD+PteqTVckoFVhs64cKoL2XO
LK1iCXpSeJmQU8pIN+2waR4XKYDwi81TGOwfxebxF6mSIrAmbPYDPfawN/1Buad4sidTofF0WZAj
26pZLwCtgUIzjtv90p9Q6oLQPETyOlXEshJR8yQwuGOMx3GOjKub3FWKJgFY842wfKaKzVKhhe2o
zbgFrkEpPjp7Kslu7c/pV/qMUGsT4MPyRS/ZOc0HEpJtWn6NL6doGhBpNpX3AwiNdl/Dga551eRc
VDpdZ8tGZzIk4SmvoA2tOAA7Rc6WootwFIZSW8JLAEfatBRASSBmeuBnkpnIFURYu5u34rQikvdX
VCLK2vxHipXaJ5Srx/3Vs2iPGy9GgfXFvg9ILXOrQTOW/AmQHOI2te84i1Xt7hSMn0qhr0Xwdb+u
Di9+xlOPm0WRiXrWqt1cXxzJ75y2Jjl+EiUAlLVcvdd/GGe4ha4UcpvesgKPA/MVPTo9InTYHoJ+
lbQAiagruK1NlthEcX/DygFgIASMK+Wot89Y6TaGwrimEPlkl+8rU9X4wSH3gTryEBwE5xmIbl5I
A6Kwh8GKemCM5Vo0IjKry1Dx4uQvHHhXKFt3wy73vvWCPxcFmoNfnYUIg+0+nAth4kRYm7pH89rT
dF0tVILXqvbsjwYhT7FoAKnpEi0PGdUNVuFlm2PkQ8hK70a+ovYc+8lQ7p1jDjjISa19FicLMB1/
5AUmp8XJbOEJ6GnRxJKjj+zwcUVlYbzdlmMUPIP0oN4xjsOaBWI7yS6e/nEDDaKVJmocI7ZyvQGw
i4i9PizYCtLM2/emDopf3xaC1euIwPmDqiDWva1I4Dzceop318Z4SWdA/1suH2MK/wlVYoAQ2fM/
MO2xSVmd2LHZjHSwyIKL9HiZtRqqXBtaZdxEToUsV1i7HC7QoKfpLxHlrGE7Q65wz9WwRvRTtgUQ
mhsV+0G5Dnmi9cM8AaBHfEgjx/T8VAq1i1hzbzrXk7U17CudQA55elA8WuLVzJ4wz00K9ogdFmpv
Jm2yBTU/C8+MdFm+cVn4x/1d4eoh7L47lqNiM04hJe/HA7eSRAixb6SANXy7bZeqVdJ4hlnbRX/U
3S22wSHeTSfOTH1stMnUlDe707QEipltoTabIJAiUywggstewCDiYQLIjlxIjqdQUsYJoGVdQggp
GYGNS+m3lspgiNBVYy1Ch310hB0Yjfl5odHeQ5nTKubm9bfL+yKXDzZHIfuXhI1NGA6h3p7ZBDWA
jcQWLWJPJhq9/lmBzkSiQm/6LFVFgL22z/TecYfrDrCdsFMkULbFT7u90Ss8KPqXLp1UY7Vlhn3Y
ifWuZGMlEMhx1+NiStkC+pRFXb39cKrp912oik3LSll49w5vFDfg1vt/N/v9Vc/mpzzKHSmrJ0yS
uSxjcOxVxkXtGTIhE1VjB5lpy+SLUtTpj/VfbfreJ49oZO1eKvR3WxIL6/0gu8BrxqUnOgIWiFnM
3VxvYJue2cM1D8TLIkh4YKYYCuzpe8Hfl//+KUPPuUTd5V9XQEAa+HhyKrrmTp98sPpGkViDZxsh
epwpyfIB8wDorsR7PbzTYkUdDniuFUBTZdngcFRhgLFgNu3voX1mwi3G0emC+yPuizdyg9SBXP0+
D8XsRkcOXUx4ImpIs4H+2Bkr5pqGqU6iuEZvc2gXdfKCbSQ4RbGyFRf3usWvs8KGzMR8UALvbWGx
/TYZIwIYGfI9b6h0R+/nuwBNXZtFrrT7VjkDH/ESMljZVN7eILh8Zsz9UFr9pibavsGn793b1nEq
KTXeUjmtbScH1/UxvGvcpNiQeyGsupBY1h19tmrD5jiBNbIz6O3ecIO8JqsYF/CzzsB/PUmMz1BE
3aLbOCSh+5umhftc6JvftRUkzDyqlEtCB7KI6GsDOxgxMwqzaSXxLzRGl18x90aTfDrjnyee7o9k
hjYGx1pmXXNyjeBC8EmHHsehEzdqX31o/ryRRcsy9a8hrAr1iOWPTmKEttFNFCNL5rSJdeVxYAW+
qLbSDWWNyq7Mrcb8JAETf96NzJf0qcRiR7EU0I0KVyOTZZUamj9v/K82zPPJPEjzrtYXLCdTWiMs
9f+El1BrKmbr0u7t1yMqW6CqOXrJrcFz8oeUJGKcXi+Y9D/QU92cOL1mx4PMlxH6QxVK2w6s8bQw
UN1EnUM/oqtbLxUbw5fZzrmTjRBqsz16MqQBfc85z+dUVB+0amU3hvmKEouP+u3OaDzoRFTHWhU2
aTTdSBtBN9Lp3ksJB2KiSkO4AYpu78A6LoHvqF2O2qy7Pt87I/SptROg7tDz0hKZastJScctx1U3
op58pREF5qaH2OIbPVYt0tVPosJtTa8JAEUxYMHbyKA8UeUzvTDblNprIyIatxbxVnRJpde/5KXZ
XpqJannVwLu1DCI7wHP33Z8rzwVMV1TUM6xs+LXb+iAxLdQ9L9pe9LQhqyuFIgueR3LVy1yzfzgc
wDA36PIuKfvV3OlGP3RRQdU4efTBNyuo1dNOzPs/K0G0mOmvK0fEDHAWkTMTiW9Cl02Nt0UNKBpA
llhtgpkGoTLQo3N/pCGXTjty/h/eJAuinNRveImoQK4z+WOl4kYFDwWrHL1ySS3uONDiAUFgKxZs
dCkyX28AmfVG4koePJqBCr+DNlH7bh+1dJQYxfDHOTJv6z/TROu7YHLBdPWIsNUihmLA6fMV6pj9
oT4LKtr44VcUSTuqwXA1TpVP6uiGV7dcjcl+BTOLi+UDRYeS/ctmw/QrPN20pxivh2jkVSAKnZYo
NfOEaE0Dbnv3WGt7Q80z8hBy9rHL3T6LnKlicO29mwZ8OQB5Wn+u4cPYwOVOGiebPn1qwJ+EoAXY
EVzHYu5yz2Awwnbf13e4W9BYO3InZ1x7JwHOJB60oxP3WwE94BAF/r1V90SISaSCop37xYcx3HKa
bHp99ieiRuk5Cibmd3VPHxNVlPBlAI7943gaVA49oPd2VDcc+PT8ISzBUPxGaZ0Tz7kraR+Vs/ZB
x/UtznwKvJ3gtdE7QvrgNIW+6KM0h6GQSgIUfa0clucC02BAVFzp0M2zobK1zWxvP7iBoyVKr79B
n6A4MSdFnQLiZbnFQCBa2hDJue8zOe/Yv95to0Ef6pfO+iWr3wd8JWsGn718NmUYI/BP1pkZzRjo
M04hQf4+WO9jy8sIrzdomyeOgwoa0Wz6qODnpte9/44DXn9G8hEihkAbH6tLkOsOraYZHcQK+kNq
WSZZgcJabkBEU+63gs6rF+zhfKih5ocpMuJciR11WG797eFRaehYdqU69DYdCzWyZXJuaxtLQf67
e63quOn2DkJ5UL6owQLJYdKnYXL3pSxbj4ZFtvOk3r56JpPLxztNlbVW3QcYpB6ajQnetWn0s43t
TN+66SRnh50UHPxy45KA+xWsgU2o5aFmy9BYcF9/O0T8vzg1RgvDIxd/Bz7wNYrVvFCJ5iDWRRSL
T+zqlklT8pNNdTSWQ9BJs3+NZtYoza3JvArl4TwF6fqLBK9iKk2A329+/iUp3/ThxsoFDvT6jQ7o
cCIYgqkg8WoDtSwX3v6uefH11lodABWFEiCFPnVaO67mwyKY3ZUYohJX9/a+B1jqd3poI4u2NydL
85+V+TWVUKglqNcuPlniArvzwVIwRLthRYz41s7fWWSJq50HLUuDcwMl937walHVLQNEVm8PJXAC
yUfAjK9jNNPx9hKdYC9r7S5Ozdviaz8lNmVzcggFFg7cfAIaXVsmOHyYYb71Kfm+QWGGmhk5GGOF
mO/cZfPerzzVyIFzTX53nD8hBqEB2LCJacmVW0lBkQeo9etiB2fNFV2hQA0rqmNORh2fWhpFaqIp
5CwCsou+baV1uPZbuxEMGVOqI1afiZL5pH9r2Ys5yOyp/+ZmocH3TSzd90sph6UNm17NguGL7+tZ
2C2eVzio4p2UQz9yYOZBKO1i3V+JAh6zv131aswgi2b3+HWfnhFehmim0e4U+tCCsTjFk3pneuy4
G8t52t+OyCElbqO864oQO5TuS+YusmLajr081+K8Zx9/wOh2X5FDU2EAUdlHzAg3nmPl81sKMTmY
bBd41NCzzTluV1KTxPw8+Hm79RMZV9rY1r/OIP7AqKiCi/pnmBcy3zcDfx50So/xKaVpLZskaUCp
NzYlYleTw6ltbPu4wEEvZiFqQh4fyiHJG6wtBqZDLHO4EVoYVCqeMFT7TK8X3DSMZsV/ps5aUlJP
SzJZA6/HlFG0wY7HZKWgyhYR4uoYbraGxIIvXpN8C0YgYszdeLYAL2IzegSdYbzVs1BI4H9RSUnL
Uw3vf0GL2LOx7pbyPdZjCjXs5vaia0KVJfTfY/r29epBeUPZ0t7W5z95gEOLP75G7vJzzoG66p6r
5/eowXPvBLw9zj4UqylomTVFJY08km29hi85+91qikiWbWUnUHpo2Pbar+hjaRErbiXnRL2nzuYR
jw9BnXLQs8ZtvbBmiQcM0gH1bRQ4FouzWS1wHsl3JJrquzXvMuWZLmnqDfA7ze+Y3Cs0fygxUQ06
tjlIKygEtIprHBQAwd7UoS1yNR7G3f1bM9oPeFyNl993FJ0xtZKXWxmJPq6gbw5KZ7FURFP2XOQs
KaumxVO76EML5fnYQ9Bz4rTKaKa62YOJbZMQ8KFcQJuIbyNnjKLA20r5Sx7byyGPV5DO0fy3Ix5V
CXbWoSwBc3Qi+RGVytl2eOw/LWbvtL2y3ILw592S8EVETdalyWyzy46YWCeT/Q9IIgVkmB1+Fn84
kT9DArSlcJyv1BS9e/Eiw7VOXERzDhQi4ufjnlrzvEN/mmAJWDnA9vmZ7/8tYhviJyM7j1zoHM60
8xqu0Ic4KZKyQ+SOxonFWdjz8jEAUpd3KxouVc7OFIhCIoWKFu+Ddqg4Cy6JHxtb/cwbPcecGP3L
Eek9iCdL+cvfIyQwUaKw0xtPVdvazwuk3DjBO8377a1KMQ9SGghRWMEwbxpsnDouptlevr/P2h9W
DCm+vhfitn/bGXx4r9KUjM3zgF8mCsNQkNZUBEMODUbrCH0fLjcrR/3IM6SANKNPq0bQv18KSRiT
3qxUMAARwmsTLuY7oI6G+jlT4QJC0Bbv2uJ43gv0FXVaGTU9qejVKmeiPcX/9yXYDV2Mea3NeaNU
qobQm6bvT2UO6j4vUFIkXQObG4N/bxGUhHn91CWsXaNwa1QvAEYVfZXCtWttER50WjNVTvGpdPhO
ooS5StIvj/c/avFkr6eKGof8W+Nt2Ehnwu938SvElKu2Zztia8kt0EKNIx4u3zl24uBHMV4fIviv
QjUeo93ItxPJ+P+lSZcWRUNvQo7PHoUBXmUI/KHCcleEsXoiVXC5hKlhtPC6fjHaQdd6IyG3B/fN
C4LLmRN4w0/IFDBcsY4SlCsJUcZeM+FL2Fgi35ebhJeXEhYhmTCE0nzS95KEVCkjq98Vqqf7ULuH
2J3LWwZ0y2DE7ntMO1we5kp7z6uapvUW51rMuwXeOeaikY+xt6Mm7sybMZ5e6Rm93cg8rlQlPHMG
6pj9i1n5oHLNzBG6rlJZSAq7W40P86DSdzsq54ssix8al9FK04MCoQQ0vWd4EqRgGWb94Rw740DF
QYHx00KSJ8g5Kps4J3WsvkFnd4yj8P+hC9oLxMVoaYHh0x+k9dSi7NEWZ1cdbFbs6efw6CCT/FH7
sC4+uYr1xoY3Abnx129YYGv9bpafet/bppKmKoMkUYVYDUuc3WXNCIFSUpO9dFzEXebbQe3ZOn78
dZBz+bulsmnWfZA3jjWPHTlZlNdj/nSUwO0kpnmFxpnHPIvvpLCKcJ8GBvAjfpoDWefDSgh/Xyvu
oPnpOo5or8zjj0qkAux7ns6CBvca4XDMx4b4uTQmBdmHwwLe+LC1A9pjQMIZuKLzpjBU81tPjRno
1vHbiS/53LBbaawhzoDeQCv0WbRVV2PkRY9OTWwYtggWAztWJmOFkiMoqPgW6W1CT36GI/903Y/d
p26+p7LYAI59kM7OzgMzJ0MGAOkkNi/6yAP8p/ARhtZsQLiyO4GJxEnlgCJlS1FvdhmHcxlKr5DL
TLoU72h8VoE6QOOwUJxxBQU5V7U3c3XAFPr7k0MfBhjrwh5+12HFjUQZtE6D+FZqY7SYtKluGRkM
CSQ67bvZ2W+nz5XDfJgbLNIQkVqyU8uh2EeKyH2Ht5OliOmHHRUkAm7CsE3CKIJVHs4ISUctjr4r
pHrp1lkaxhYo3H0pl+ixKtxaAJy5klzFB4Mq2is0k7JtakfkdbjZz54kC59jCBhWRjlcw7C6NpJk
STm5Z6C4xu2OXwPxx5siUrKbIqvUSd5B2F3RpcMxorq1GY5IqFgCQORS44tXdvmVbRinYuLwuo+w
lpEUR4c1cxT2sKICuJ95ttinPt+P2M1M6dqNPwfUulRz1cx/2UIdWHXXF1ShPBaytd7PPAr6cauA
+hss6dwAZjkhh0XuBBA+ggvAccnG6Berjquev3683pAL9vEE2czPHd+egXdTr4T14ELZFICA4lW/
0PO9cMIL/fKntF6yDMcC+XIe4EJtSJvyIztPMvAB0pzodN0jwiPPzeOt2b5mLN+JlS9L76Jju1N0
nKcS2UshB7FcxG8XVrhVkGiZL6/7rUtO13KcSAPpLiMyv9h+1HAtgyj3IT4hPYktKQ1SWDGHW9vp
8iQGbgIv1bUULzFikXlEgIQ85sjVkLw4NobwnXLSeBgPs4/rpcl9V1WLTCkGZMXrpGDiTjTpLg8z
o/13xmLIuGudibWYSRmVICPodBDK6afu/dtZRB03JH8c5zPQkciYPy5XfmH8GsHOQzeFbdgwAaMh
uK0P6JFpd0IfyJb4pYzLeSR6/bjv6ciy+WOsL5j2VuBmKUWzXOuxnLsmVLfF45CCBl53SklcIupK
nx9Dakte1aw+pkFtA/5ubVAJgEtCGQHwXFlrutLu4SvIr6wlMqZtDztG42kc+Hhb0Pb3UEAdcqw0
03rQR+vM+BXxGvTYMQLJ8tlR0saWbEqEUWetqqW9HN7wxwYWdX5IQ8Hr2HALziOGsCkJV28T3woI
eWq/IizUwHylUWAOLh2Rip79U2dlSd9JLNq7DMspbmqUrfsSbcteijFmZqIjUVl+d+6SnpqX6qBI
qySB7PuJBmk6LtTFCza6Zjk7zgCN0h0YLLFibO7K7uEAsBT+kccXqnQekCSJ5P4JIKaMTFGaH6Sr
HkvMsuIAE3jaJMPrs6L5eRyLFfRv/r9fGvtYbggK0L/6HdzyUSBeYEpRVwNbsp7f74Uwy9wLK33W
7ezWPRvJtPmFz4Bh9vZrAE0QGhzNWbavwkrsetFIlx1S+tE5DCNTyrIZu2IL8PcZEYbzjMYydgOI
fbxYCGJHSjB8DDAowxZErCP4CsG93PY3SYmHgWvRoaF3N8QuR22+LHqggQAdeP5vSfDkHNcOTcAb
JWGAQegcxqsae7IAdYiICP5/hj4ZnhrDNZWSS67BuvCQk4G4/4hl0G208oFcCuszFFI95JsCVPOO
hJCSuOZH3AMynJLwI/3GfzgsQR+sYIt5cndD2CyuPSQFbR/OR+tgLPPcw/HbwVcp8tLvPmCEps0x
Fae85/yQiByg86EfoLnkZPIALgtvkAvntv01vHfvvhdTZSazSusLR91UUTDiYvwcNySDwdDUv87o
gmVb4k0DVkZYjzn5kTAX77/hNOqickHeEit9Q+ebq2WPq2k6csLJrhPfJpw2Xk4VyhpdBL560HtF
oY5KvL4Xu/e8i/L41rZZJswRZEsOaySamfZHJ+LWl+lq2SiQQjGeR4ynQLdJdJRdRiRq+ezTOmA9
aUDKhEhtEvDUWGgOpiGVDsqST74m5BV1kGBf6w1iIx5FN9genpUvxX/nI9edMDVerko7VVBfWymk
+wwXzg/EQ0opB5gHKSfjWjfAuY96UjDSwn7WHXSm6Xxh3JrHLHweiN8SWfJkSEE01C+FUCQMjSZX
CM9kIs+rJ8BWH5jFBe4TZyfe/SQcfNMKNeS3Ydi5y8zQFv2QcKnl9r2oM8enDsMyuQZclSiGweX9
Y8UpVQiZzFtK26AcCEBWlc+K5qkyc8z+AR7xg66g+kJVuF1W4uXZi9FHyrxTcclZk3+1FjMZF+He
pCYZYYHFONKASAFdVQEOJObaUa04l2oLojQM2F8xFTEigjstp4pc1+0ZgL5lfaHVIs682CkuME1Q
ts0jUBGH8FNBm9gKB7yOsw8E/9ZgZaI9wlLuoDS0U7gGc0zYeSBccFxGXEAvfhlhy42sDou1g9MF
wtGxUhp74B3+DUCgJRKBF4LZlIqm55wkFIG3pqLN5uS3cffvZuH/f+BAO8lLZMX0hm1n+SZe9/8A
ZKPocxpVgpKJkc0O7RlOTiNOdEU2jrXnjwHzB/4FoFkKKNoJHWnwAlnA9N9UX8q7Xr2LPkq4VvAa
uY1ceumFO2hZ+FCq7nibxoZSVJxxL7Jnrscw1KfhKBPfhFCsv4+V7sxIMegDUBL8CiGPAoG9OTjm
VI9e2eQGtKoxylU6LzTPltv/qAtANx1Q3cr3craDkbAVGShYX6Mz1Rzcyr4cu5a1w7x7YSW3zjwW
zGLrZMaDWJu2kJrR3edqLfFnWQcBn1rF4Cchvg4P4SZrXKfP8/YJR0C6D2zqLz2ILSGAUzapLqoP
q2N4I5o3foHOpiW4wpfdsEJN514MIE4hLc+3pURTVRf3HFlayrIz7w6P5ghGU3j7YuXnuCa6eji7
i91ibmWaupK8w4KfGigmC1BXxYLInkwWmLUcQOSbmL3zetmdxJoVApeNngPGH8VD9Lz1039SbI1H
IjN5q5y+agiEzoKELe8IZygyf9Mfdt/XpO+U54HV8txDwjqbXtFmVlhqPATAggkt8/5Iur/BwkgT
w0TiyAiGfnWUiRtYAjaSF7iBb/4riaOinY8QrcJxtgyId9GoW4TUNtOiuH18BCXnqiQ/0rv7m326
L+/0861tFI5ztzD9HdBBqKt4vqn377jaVicAjSG6HyFkbMQrBID+uRb6X4M0IvlUG4iQQAZmKBj+
StzyBFBaL1rm8KE1UjdprZ0ZkVVz5256Pd9DLPwMpV5EGWFPn1x9sn+tO0PWpGDD/GyE/DWMdaFa
a4ezbzdLCd91LswrWnKbV+tbr73FMrJA9dJ4EOKy6/lsWCEWYZO0SK6wGGRdTSZykhBPZrNxOnGg
x8uvFD2TNUrf5+iSO8O5eyQAb2oCeiFsfwkSU0lYOWCqc5muKbOspgkHLdhY/FpxY3mtW2pjaPuH
iyzHyO5SLn9U+ZKtqPkX1xCCve+PqCdFQwqO/75e6LMKhvcYHY8HuiR8RDoSkkmEiUpHoicvbWVW
PfOTXNBxBK/NUCG1gbAJC1zuT1mbmG/appeTaSHo7jN32C0KBjiXDmJby+TGGL1n882GyxunS/Wd
43IpDLO0qnbjgPY3DXPyL0Ym+WpRH8OaOMpijG/NJBSTJ/yiSvzwkJ6yxtJ1TXLK9OkJ2QSoPCVh
Qs4uRnHtUVytJaOZGMHQVqA8rWmRiSczvZO7UZW42YeuAj8bmUGpuHGfpFnC3WTeVGDb09gixtSR
VBeVD8Z4rL22Elld5Zke195mN5y+rekGIz+tRk5R1kmknYwkOBDE5KRjzg6+Y625eoJa1X0C4GUO
CNHGVF8GEilrpZI/Z5DwowqjpuW30TKiP/7WAIOFIF/Px07aZcY31//5WZf77s2XwJjqzOaC2mHR
Jf/Ds4xcH14pjtJbHtE4fxIahhe9nSTWDHl0lP6c5erIAaN6hP2Ki0wjRkjMbGTI/EZ4jlZcjF1k
LohZumWIU3KgeNi6MXpOwakwJSjnEKQsUvwg85986kGVeHx8vCDvnFBPh37HSGttlEjTBQ0nb/lv
CBh3LuY5jdkSfDIIQGTJcSCPgV9wdKsMtDVBopIgbXJ/4SbKUGtm9QxY8U2FDooWQsTaZNFxeux7
Rji5vU7kBtQFJlYVlLK38CtFlcuGMQI10Hw+SsJJkqTtDCIQLA1kxlQbSyEEwWFWkkEBKTXmZ/7C
btIT2eIMxna+zPfVEGwU/I1FvZ0wA/8p5+ef36nIoscBBJ7pEk0Oe4A4eqF4rzwMcIG2Nj6i9ELA
h6wzfZ0yrqXcfKXPAQ9tUgmxKr3oWLzmXKbassHPhsvnKb5fg7WS7xfnYQDgZt5F4G7FsulHqLXq
0ggIjB5EyUEsC6OtYOxKQInYJiGU2lVe4Q54+8BtGFGR2LJTBuAOH9x4Lok+dlrMUSt3cSo1PoGp
QPGZ14xMprpTz2vKLgIi6DbQbCfRd7SRkc4yULeBRwG2Vj4Mc485IDT6WAtz/zdl+uOjvBHx5uoK
AFMEBCgt9t7pjTCnpkwl8PHHoa5+agLG8XyaoyycSZShxD11N4T656/9l1KWFVpiiIIDt9FdtKk2
IEFcdoa/QgCjaM0sBtMZ0W5KgM7EsuGfK4Sffws1PTsEcOT8wEJGhUM4IX5c2nAJ0APcR3k6KMqg
akd+Ae2wqyXyDxR6wgpejPBS3vQrzIsPKs8sc4c6+WTKIcyS8sl5HZZSIcETPxcUURxlhLIazkZ/
8FN+HZg/Zm7qkWJ/qvPXjrLVKhs+ty1Z/rF0RYKkbXYVu4f+LRpa/ML65HI86fPHVECV8fMIx38e
bTN6ytb1aUcLLWLd3mUxD/3qMafG4JgiFB3CXgfKUzpJ0egm5TE1rQwkVruejiNejTnOwPIW0XwU
EoPiDh08kncfoboxbJRXtmCgLiYeSpiwYr172A9Yg3WNTqxzJPaltbPR7/hFgcwEGxI0f5dqYm6x
QSyCd7Z6WTxovFntS+iihGdjWlp9C6bI0TlRD2rPIHxqpYJkPVzf3mTWaDhQ2cMEwcTiavTjRoq5
n+un9kXa552mJDqBscfooUqmn4X/VWpnJRelgF997r1RbATxEWyWOfbQPGw1jiUjJ0y8iIuLMAun
xwES+aWHtqZ2/ypJ6x3JFfymRAYbqG3u86QHqttC3C62IyYOYyYHYcU875uVls0sBWqPPpgEYQtO
oIymhXjwy1lEuNdDMud7JvQqSMvFrTY8mMgA0ulb3nXl6LtvR2saz+3AKGhDS2Yeu+OanRiNy5EY
lurOZPTo8myvAom/d1XAbBg6GkOfvvjI36fGO0s+fIei220PIp/IhO74SC7TGfI0zkO3ecpTjLJn
XGRZAEopKL2gq7TADk0XxgiI/g5B9nkuIT7+jD4DUBriMFzyPI2+HJ5ud5WrrPtUBEQg6JhK/l4h
YsvqyhQrTz2PHtSfFDgeJfrx//e4zv2sIKt9EZeiFAYqdCIoxsx+Y7MUlRoLrghj7u+u3eYCQqE/
GvjJXF75DDKWWM7at9oO31K4dbeZnSLmHj/H4HhZGudf1Y9oDoBLqSUWw2EwnS6V0OXiL1sq+JPY
GYrnvS0DCVfWvQyWJmLGjMBWJSrjCgojwq9YQwdkJ0+fsJIO5qJzjhMIogGeZS73c+FtARIS+eZ8
rEgeICwJDH4Kyh1rRSsfbp6BMYftsrkQBW8mX6jJVOJIA1FbHSTCRKY/I/F7lY001DJUKN5fKzkh
xKSE+xbWbVDotgz7Ttxp7xEkDfyjA5HF1ArtcZPIIAd/1G89o1o4i7ElVVHxfasc5wYvvfvWMdOg
vU7sJnzsNd4fsZVRtdU6ZhkxLG0VgXZFI8m9bjx5YPhlcAIxnKhG6axF8UWyB5jpBIVCWxqHFyAR
Fs5BQQGt8/DBEfPMTR6KaTyOVXKJBURnoNm0Ii8jhPHW3QT3v7woWLGhTf2GsELh34mUHN46Sn/c
Gi+I+X7PzkI1CZYfrrw0X8poewJBSyCtwUg3uVfJhkiLM+7bs2EjpV8VCtyekryNX9A/OdRtx15g
mBj54HzCX2Qo4Z5zf7TVXLTD4foYLOOIj0Wames5xF4GipCU8aT8EotLTGULwQGIIy/wCjp1cgJI
csHjvytNt4NrJd18Oq1XwxgE4k/Xt91fPKwkgOjpd+Vh1oW2vpfd4m2DQJmWXEmbMJAvnG5uBq04
0yxxKtp6+mocFCH5wRCWXJdB14PxcEXAGf4z28NDf6UB6FJcv41RP1OYieQKJ/KkaPRLSJtbSlJw
WokQmOYVif305qXmsUB4pnEDa139silaz9WJmCUYLmBVbhfG6z7kq3ERehZrMDW2/OV2VNi4F1Fu
AQmWv2eJ/kSPnweELd3cUbxPYN/sPJdPqB1BUMSGKoG6CQgbNAr4mkXbS6gGjI7ATXoYoRSDWtOY
iqfIT38EyGJYAeBOjyB9LNxcIhAaP3+/pgeV9Nnb3Iv47RmZJZdEL5dXyHaaRPwx7tEKwko1sfvZ
Bh+qTJcnfP4zVxu6FHilbbqmZoZjyddOf8JQzHmiwPOxJUmClaa+9yu5rMgCOXYXDC9qJI8H14sC
YOl16l/qwuLPCcyDDWivGBo/SprOLlFWi0gKAtuYwKdOcH9/h8t7oFUnTqnokPjYl+5leh7FZhcD
egvsZyMWIBsu/KJ1hGy0w9Z2VX3ekfV4tgDvYP507eYYvjTR7OiOUDP2okUeCJ5OJcGfEIkeDK1f
thqs2N0tbPV4oB4n712TEvlm6HHVJztRAPzidGAlDrfGBfEipTlM270BI4+BXPyG8EiAEnJCylcz
uJjq9Aw2LzVab7l6+NNS9ZMhA6Or0QCFhKHtmDpDu2NTXF7ILhm+rFfyK1/xG+lSG4+7XBtgkrPa
itMEX4KnV04hw2g1AS2Krt2s+I2AkP3F8YdGMIThHaPyql98Qdq5DqXN7kgd/jDArvhYMr+cpu9C
ZUo6INFaIR9pGbm4dAs38k+eBPh4aqeQDK+7wQqKRvfoxp0L7N/NqslfKoxm5lXFzojndbQ/uGQL
ZzuO7VPYykn31pqREseh6cKC5svaKDvlwtJVcXlPb9E+NrmJRw3/0ZBqeJ2neGO97MKAe20MxiSI
yiBpbQCB7GQs5FxJ7YOUvgbn0rYfyNnbTPLsYDfSYI3FDRJLFViSTblK/f1IJDJTZdgD2dlOZdTF
Ef3aAX5+oZNMx5Pk4H28xq+yLNbMCrgAWrLI6Cl+8lQciReoW0fTeuEVuVwXIk+XD+INyRUQ9n8T
TZ+0hRKrrNvXBuZFzSPWNie6ZYACF8WLroIC4RoVQ/ZqUiLB8vXYVAcl3es9sdQjv7ahToIoZw0l
mg8QiCFgRoB5Levu5t8vWfl2Rz7unG4p/u9GO0QTVWnsaJOGbdyCxNAoJg+/Gt0SQETVC1lty/JG
kKOH7di0RUh34WGw8NJKS2KZ0/gfGyF2oeNqcyW1pS3WF/Cjy/cUrwyVAjk9qhYkd7ms5FNwq3xV
nBPOBTuNQ6TOqah6uuQCt7tcdO/4JwYN7WUXFKTOf7Y1Ao0/KKNXULrbPpPcDHJ+bXKw3JSr9x10
NBwXfefPMifFJoxLy3RJYl6UiReNhnyyshLHjfDQhu4b1z/vNSPGmoqiK8oPmZPu0Tf9Q9LNSOLW
eA2aXtYL6GoCZB9GHuaZEn187ieeqtqPq3kdfyPUzuD4LykKQ3CBvXriKFxpaBOxrxqlWb5eLdY3
mePsuzbT7muieQuNJLr+acPM0AtOhGOBqKXVaMIiCqoe3Q/0ZVUVjMs6xF+PJaOBkA+G2Ivn9SXM
A/s1SCFamwoQQraOao7QR4wrOkaHCROKYQvo5NNtj8siSapTqQ5fSNTGI7U6dDgJIpnqnHaQ/xIT
MLqgB2gsuvrIX7s4wShiVkZHjzQzj9oz8XNWAaBJ7oNRD/XhMufNELIUHOg5hCGbgUbpQ1prL6qU
JOJ4z70CAs6njb0l6jeg8qwTuj6XqI6iBF6s7baaVMtH5QznU5S2FYKBVOC1uWJdFDqlw86F4A1f
OGKe9fZO5Ni1G36KKkB7SWLJ2347LpyxHdAbCXqAYy9Bt5ldT6/lHh0PELxp7KX1AjrG+LbifQVW
1I+HwWTnSQTkcRVl7vUuhoaH4LmVVupDWJJYplK+RLgFpqTuKNs0BDDZ8qecfGTpjekUUv6yNSin
i68e3eryHb/4FZbVw3se4bD5+ClNX8b08g4KWC4gtJaelbcK64Tsqw10Nbk9qtERT/XzxywTpMtF
VYvPqlx3sDCIM0nSynUIHLssgef8tY+LujMUrKF0F2lwzySagu9n5/NI6m1TMpUVOSDA5pnpPIdq
aXJQVr18/oheb+M5JwWa3aiqDtUFA5aEJZglhMOqqFunD84zImZ8OLdrGx2macVYlP/Mpoafu1Ix
varL1+quT6VjNY3ZqmePytvHC65NPLRT0BHckXJSel/fh/053E4g+kRkMLnEEAaorP6Kb9fI+VB8
iaw0b6/97QWeQ3PHY9zdcOoWfUlMa0MNVVpmGAE+agG7th0X7yg9V/19Mu9Fiymqza5Ezub1JOVR
bFRUI/fP4HdlXhXWnrEUKgTSss8NdHX0BR9O7mJn7pESmcbG8dr0Y04l7HObAq7W+YmW/UbjB/5i
2Amdw7gJwW41cRfJ+vmMCxDG8teEa1N/gIZkLQ5XKv2uyxbrZxYEtL7FQUJ7dzPDk4WSKYEEMkld
V2Aas4/nMM8lHBB4cyl5Vh6IF/zVAaNAs9idJdfq4du/v9z29UjbeyCEu8bZ73CGzzRJp5DwRO9M
yaoeaWkhsoIQan5U11EaAE7RJbSxjQ3hLncIOCazERCWmDehyjfti4/ovX3h84DXREJEbiudEJ3T
x1FL7fz4HprKk2jAknNX8UjeNy/uLikUOFrkAJCkystwxSljvWQ9ULZeNTcoFD+l2Wv0bmDPOisO
QmkqOkxO2SX5NFNvYA99uVg5WvdWnGMWjMdKDBRGh4qJoLDtub4ibDtITvVozzLz5sG5johauqbz
ILLbm6+mjFGtfnXOPSft7rpFMREfSZsredWf9b3TI1EuNbH0wkjpoTXf8Xewv6wf6CbnaPXKa5f2
zstdHdf1ohPrn5mmLrk+4NXphE4/7L7ZRWzUC5U4ryLJhXTkjtP2IOUz8htAz8yACtrrs4NsPw/H
3uoP19tB/vfAZ5//ou78HeGZsdjA+G9P8BHRmTWS2G8IkEq/lLZwy68a4niniQBWHWPj1hpjDAQ/
4vmGMEPOwj/BdU+xokCJ4efYDLQaTnv2HkyzluDXebbh12uRM17JgAGR1tYKFkwCMMNb6lGOxCJI
Ve+PhnOLgWOJHdyVNC3KgicdLy4+petUBuouDN89v19qZlpf36OePK3r5EGuxNqsjdYy2HJxMRTv
lNPDcTqubkH4n9mOb70FtoygEp1TNjpfYxPmDZ6Gv7G0HEtubdmaTCoayYd10jsO6GKCb4RHcvzd
WxwVZS8yg7kXBaiIhLubDPAzeh5eQnqxFQcA0eqNkDzGVo7GZyhASuCTruuD1wOOnu66M2pQwduu
SiEu9Ga5KB0EZRw6k+N/h6XjNfhuzokqCUtoBdDgc0W6HC3TKnYpYsGz0oz4Vta7OURCSJY3nxRG
PbQYwM62/6pR03VNQnfIqjoB8K8c/3muvrSIUYyOrvbl1e6onIN8++LojA1LktkSWUiqOjYlq/ux
WfcyIeDACo/AbDO2kMdtqufNAjXuKV18ByI8SDB9/C89yvVwvC6LFu/9NboX879TWsN3XnXyy8p7
Xf0lIZan73zqBABtaSev4R42ABW5LZso4w3srIrMIfdyn3f4GJHXGmWvOpluhYLoIO+KsEXUoSEC
vtrnXciw1lHhOtGXFWb/fES0CK8HzKIueokNvefC8jEryWJKBrngZ9WRCMUWn4tNpDXYo5BKbeC3
olwmsM5f09Y+BswV6hfB7UdlJcA3WF0rUx3pMQtMixSEzTz0C3hQpB7r5Bc11/f44UMV2xSRyIOv
rUy+74+Ygi4CjEPdz28Fs9q4ZkF2glvHQfMY3qLfc72pUH5jpxfGoUWLiMP9NuUfx2RI0y6YtoLP
YlfwQF79pcmZztGGfcaovPhSjUm1u3bEl33HW2tcb5l4iyYKcnyrJcjjlIjUQE11WNpfnse1z437
ReyvbY/ZtsC7izdkqUzCmsHTNOEWpoS3hg9SfGkZpdNyfAjHV53q/v8ErOPcfmigC5tAKqJFLasJ
xrgr0NruyJBqJMufKr2m22orZrAkvykhIInJvxH68oadqp2Q7ndMZ+ob9lcHfvetT8Mef0KF6rwk
DlmfR5USuVStABLJByY8QB7cetFx6CK+Nm04ywH6yZdOaBEzluRrJ6iDgVr1XMjZ73xJiozaysj4
22keHH43q0FTNbMq8Zq3KaoPoLIIfzEDNgs/Xf350hV9JVgaY58Ulnvi/7IBTeucGFk55lGW9IZv
nHvy1rrhsVgKmIK4crIBGt7rH67FBxspEJkfha8iH662pdHxDU0126+7gJMwqzQMRaNNdHJGzf8Q
zryCaN3xOacm2zQlNsqA1zI7rlAGqBmMTL0LDYvX/e/hEqSWM/kS+GuqyQCOW6Cwj9qPUktLxMY+
C64ebWfBsVTCjg7wZsEOrXzVReyfOSkEQgl/9s6BQU2+ey4/lcluWIXJIzkkoYaUpg4Fzo3I4lvk
Sn0VrsO4F1qXp+X8e+2tLGwipfPQzg5gpTKl0rGOFMN4osmAvX48tIdcuqw/WFz5ZU8j+rQBtJct
drgkbusyQHIVk7H+dLJwmnlwHg7jEFv/+8poxGKFvHna0ESGbIQnqdcoRHDo+WaclmDkYSP/CRnb
DHZNNlwQ/+Gg4HmIe+kfimyRdYQBVAF8yNhYteyjxuux6zlhV0UKxQnPVjYLLZDCthwle0WcAWAC
plwmlK5T2hS6Mbp+5FTYH2xJCO9Q5caFTEwhdksPHk4YJxoYIt9VCnIN78yvPNOexC729YzyCqW6
Cj1WWZmU1xl7KgS0ONAwPYGpD99uupwzN2+5UBc49Dhnu59XsQjL8WPpUimH90Y/DS3c237+81TV
25W1pVCL2liXI4Y5ePvFs1jkp8Rb/idCZMrW9DCKgEprGz9jLCz1JDX4pE33tmBGkr+SFHIHH/rg
JrDbKx0aZWOSxAfz2EyCm81m7mN2qFSecN8Tn1s/Hu7i3/aTLXOXnHvg6TXH+K9850b/LyXwOcTq
sgtC0Vi/n9bUaUHUfdjmZ+FXIlbU/m0kNvphdveMlST/6gyLpHMreKjXo1Ms6viIcaLKVA3Jlj2Y
HbFxYGIz5Wkg4Tb04laI1Ye3oODKJqYWNWXFr2u5ZYB7t752eyHP2+ic83RnueljXLl9siX0VhDL
N3eu1dxJ/8WXqnuRMimL49jA8vCw35X6IVNdj3OPUKlAz5moMwZ55TJmKtoE2MSrJ70Y+dDB/VyP
40X1DfQWe5bjMqR6FzckSkolDMBJYZqx8r9PcQUxkjs5x+n6pBLsqiksEKxNAdk07PfcHbZwalhK
HAyJtQuPYFIzGgHDBZl0bSJchBITKK9gdxbw3OJFafIIbxGr/C+8Y2EHo53SBf/5kiwxPVozm78V
fRzzGOURQKLajG4J3V6hgZhff//xLPXm8yQpeHCqj9ISTKXzpTEGe/ZV/uDFPzEy6ns80tfjEvx4
kwEWi7RTrEqPyYisCd0m0DyLT8WtvRZq2F4oLSWpEqvL4oi8Gt7v4x/6/Stux9j2GOSV6bJKfJsX
Z3WVmiLjbE197c2End+c4zU9KZE8JUVrfLnOiskuF0zXOV49Yf+XHEVw3dYirZk5DIU4i9Lb6MAF
J0rbda8qVKIpPIryUzXmadxZjNWTpuqzeH4y4oBAQ0FNyw9+2jVfaYRSlwzlwbdtdhzk3CB80GvK
8EbozTwMLAggdh5OEpw2d4RNZvlmi3aua7WcpXJ1OgeGlKQ6ChH5XnwC8ODJTG2+3d94FlG9ZYo7
dyOSrFG93NH4k3T2EB2z1wldSLIjJ2b4ad30/Kf1yx7gc7+iXdajdMklGmzqqh8wmEUgNp+/DMku
MS2jYzDObc6Fl7bRZTfrNy5WRFgykzjK+pv95UWFp2gVUOb9/8OwlXMYytu8rPYYkDBSWn5b5IvM
x2VjqO1muqmT7d7BSRrxqSxbgFOwmaOt63Usd+p4nOc42SeNrzdr+07BBtbv2ta75O0l6ra2wHhh
kwCukM+V8jKbNoSJiXTRd8LJiUFLCihor+qWkZnmIpzGfDa2OQZF5lWjSRdljeAYx9v/OxLvfZ0q
j0x/oCKNdyQt7YnQm18jdgcMzjUvsHl50Mji/VG1JgfcZWY4Fx9oTNEI81tSi5gVjwG9f9YdZ7My
9K+Q8l5kge7VgKwS95Wi8HKaCNfPGuIThACWThozJ8MU0tW+FcT+3Pkf3URR3JK+g7xzJJm1ffww
dm1+u8Teih7KefV2fmKIvRcWYt7AIS072O2MKVldKTQc61UBcX5fOTCHHxarKTSk910+WcbH0EM1
srHU4sy5dCZ+FpfxVbYX3KE3vHcB15Lq2VUKHVRF99QSI552uBbAngZEgwzPddMMZM/cO3k/KmNQ
RYdwBYHriEsckWZGIzu6SXZUA5XlbliO1oAiSFUYi7X4Sr5Y/Aj8rn55n9PP7DvlMqb5VPXJlEHS
Ndzl4EyFpxG0lw0lJs088OY9CENeUVE2//7EDlvzB7HvVaJ9Oa7xrRSZE6MygGhwgDZw0N0F9d+3
zdneD5EKtI5xuZUS/jCKbW/Mx6LKSAeSUv2ynJKXbl5wOcRaQzGv7f1QAlVr3QElghzqLPxSt4v4
5OdVOOFxDLAuv6N/eqY9LVaWGu1tnNz9Y3Owei1qgqPqk+WzGeACTIWSC+N9bIFZZtdlRQ3AfLbC
wK+p4wpodjVc626SqhHqmzTLyFTo1KxgKT+D27w0L8rSvU2exAxunP5V539YjpcEqXU5HT4qeiCq
96eZ2ojyvAnyuLsPdUepfPAfxL1Z4t94YVWzGNMOZFXvRzl+U9DgsPwrfN+qSz81QYpQ8Im5cR4S
UTZDm4q9yFKq9+u8KZXS45vpimImcCEZ/TTpyD7dvck4s884qS3oY1acFeDxdRRGthjjTgEZs0q7
xlSm8nqY8e9j/LXZy/IYaavY+Bf567xY1HZXfxK6ZHfz/UN8QBb2AsHG01yYnSU91+fO/7NIruej
xKpdQdiujMeIAFBYXvcxaEa2MJbAqd+oXxb6Ydu7I9EXG1rji1kerIXuXJ0FUHf02q1RKnW+KHtf
M8zADEjFWtkTgtcKSRW56Q9icqDKsIXfLxcCvXy/1yMehCZA76HcLUSzL2vd+SrNsAF6O0L/PxSa
VUXdSgXA9Y/4jgVEMaw8kJyHCSCdAkTdMoz8M+UenjrRCrPo5zgZbi3j/6u5NPyJbD6b+zRjnHDA
Is3GVftNpi1Dut6dtK7M844wV0tTA35wxVw02oCJBFu3k0sFYyWVf/flGN+TavFUhdCr2YwtqtRZ
vNrckPFXYJYRMkR9V5yLCd7dJJc0PI9RhpvqSmW2Ahe0yxTpXG9MKXs9WTrJh5CaEgdDs43ErBiJ
3U1O1Vhbjwjpmahjqj7pgrereBZHqtFscOfWB8z3v0zjgvR5sOoLR1IW5XYhWn9bFlSKdB+t+4Br
2grVGgwXGGlOVhuZqgJKC5rUndfq5S4GtyZeaqlqWXjy9dEdRcK/TdNiS8tE4rr1S4QWJumBvDNf
ZPievAyLJoM+KvZoTMgjSotlqghVa8qKBKoHptFpliQ0XrxYByRFtrv4/DTo9iXyxw47z3+SCC+b
5s1uOeo9od1gGEYeh9oJvYMFnQxCvbt+ERqqgrzGlC0r5DOnIFXfnsNojqae1EZntxZEpMPANY89
Gp8aybfUxdYNzMTzJnh44jYDqGR8RePevod6r5C6rthSpOfmTAghmwdkP4Xyqq84suXEJqjPIH/2
XcnLGPGaTajNX405+VlycUsfz+CfnvBrHI5cBXm1QWC3Pq9UMT76HWq0eGvqet1Dfr7enh+u4Hw6
QHU8bbq+hhA7xYjdhm4O6B+WtV4KP47M8BoPt3ZgGiVQ3iF4Bj9rhMIc9TCPwNPpapBGKnBJFYTd
iqqKyU3IohKvQD888d8PyHBFqPD+2SEIR2IkKNmV3dxXWH5F1754tocy9CsaL9wMzt2BpVVPF6G7
RrxF67ywXVPoUKMPFr9jfpSNxkEVXWCgc9b94D4cPNKL5CXx44140haQbwCFPEBCetqjgEi/UR5I
mnSspJGUI00092ecG5LyC4bl5TfUTaqvMQ+HMxDiOIsughwhPD71ogA1X42TqhItg2pv+lKiliOQ
FWeolYQttt6lvSUDPuhafXxHXgUQaWF199uwDKfqru5nEvgX8knk+txpHszsK1PxVogeKQ+0dnxG
GqmYmIOYDsCT1v4KGx0nP9Ilz1kiqNtiGnH0dsIov1WXmaEFOkeun5nQfRQIBZwitIIUOx91+Adv
YFVThaX4Ne0FoRGSyz2WjEq60bd8wPHYu4ncT4/fQ/IJssYIwBykA8JUkWFZW6zzU1qYzaFHl73P
TXXdW8iGJMHOgOSPTWC2FhAmpf3AxdkoWqzCbfojPUP4axGo/sGctbFw8sibOG/5srCBCPppBDFL
4+OJiRzENPor8rsmEdUdNxs3lupIvtZ9O24uUfDVTg9eR/lt5TxueLDxtpAPg+I2zBe9b876wZzh
9e0+qQb3goIOGlFW0kKbtIadn0rkLev3u/v6nj1DV8nFWsIyeUwucoeRAsHudsvLNcm4mc0OCaD8
64X+Dx7RKIEm/UrjtMlsYCzn02FYt/F4Jazxi2ME1P5el06Xci8raAEZhsqP42mAYsyAqCLuukm4
nfDL01yKOYquq6Za9uNf1Y2DmHnqCgFH7JniXcgrUDzNw5S/ZVNHT8hViRazYaX9sXzGdIu7P0ou
r2AMrrJBmJhVYlvzDzSp5IW4RKA1HhDA13T3KD3GsaVLgWgU/iVb/8/I9tu7ZNg3nQbarWAubJx6
KVYuPWJo/sA6TKZc6zLTzReVyGEr1wdCTT0SUSnbsqyXSxCXt2muAZezUQVaBAbEFehbQKqfYTKQ
2fQHMZuhKXPBB44Ei4mpDenifk7g5uwwdqHIhZkDuk7b2HsNDgEEiyiK8h5/nZllgxC42l35TKYi
kluO+23fFMRsrnmUKkxKiyt45KHXgnSosABJHDbSIumMWr1uZUBkLpjgmx2vwbGy8auTqaqn36ki
zBh1HjjrgUXAn5buRnbWnlHca6HvpUTmChXlYH25BNBTchxXsjMrqzMKpOFixifa/jEdI0nj4kqQ
hJ4wBjETnmY1oQKFdPHkNSw6fJ6eObdYaNjC1RexH5Ze6+/1k3s933laXyQVGkGItD1wttOdZZlw
zvfI88BugoKjttIDICEuMF+P266W9NJaGv6HnXE2TRlZfl5sMDl2mlZRBxjv1y6NZI4qW54IUVgu
gkAllF0WpG3jfCzJmf5SeQ8zSrrOV4y9OHiowS6hzKRM1fZ+k5yRJR0j8MF1AMO0A3dyLO9rNplv
NrgbYBFTFvy8fXvNGFef9YQva9PUOttASyydtmctH1wSXnEbJBKF8gm4VSPqK4j5jvcMMNRtqvdE
gEjsrscZ8z42OKNn6nvqBFZVFbR68gElHS83J1d1RTQMZnOMiSwwuBBWFMS+q8dtmMz7kA3Ac8Qs
3Nb1WfJzesMSkWKAXI61nAEFmxzd3SYxEOkZ1G4G0YqLeZWIHKNlExHSMH8dY5+bHcYu+DXjvT8J
6eLcaGrc9DApGLRW497WhuT1ibJEs44E08ewf+TM1+Zuu58EhJ8ybq9gNtNOW/fxv+WsqFkdZaWk
yzEwK5mjynv26PmjqXnecPei4HeHylVPoldGK89Ys+fp2HTv5sYqLQch8jXGp4jlTW9O18F/1Wid
B3lA8cn8TgAycNBjaSzj+XXzcX2vbnDmvLARGgGzNFjqHKYDfEkoHCaEuRui2sFFnGK8tMSWfnTP
On2QSFdAAjfEMhjsmzl1QmYCJFNV76s65MPtvTqqFCIpHpBq2ES7c1AXE6Nh58Oacq3wcQ1WUyBx
peHT9GK05IYZm94Xx8J/sBucJIAlEUfMvcZQGmTA8Pgxn3vZQJbLekIqZdsEjhso6VQ4ltJNMO4o
bIdcMSqTDPnh+s9Q5VjF4JDVXcghCb1o8nIOyH8lbGn+6AlwIuAwP2tZJMBnG8PyZaLM16EyKJus
V6F7/dj+DjMcqFGVop30GjQB8tL1eSwFH/ABDdzAy7vOV/Bo0Ph78GWedpqQKDjMZpCBnTZouDca
Aa0aSy78S2pzJe22IWY77uIArWrQPqk3zERfQbQHg82B9VvhrjuXznuuIFz9EfNAnH/V9H0T9okX
nw1iwjHCZj2NiHhU/ygRxC6zbCpJAvnR6UM5clIi67aU8w1jkJFFtsraPtLRGU0frv9Bf5apY7CK
lKaXG1Exp3hs3Q0EbwKiPPs0WQR5LCiet+EkPaSN5sGGwjn9tN9KSOeM32JxUir/SkqvxAqUzCeh
ZPWho76rOEvc6BNuYZ3S7nKzDMMdnslnbz/T9QqYoWQEsyxCNt445sfI8iUc+NlcdLZc8lWpAY41
Fm8L+C2htK4qdYXu7h/C2hMK6CapTLPwHT4Y7FuLwxOSrth8mCO5hWiQy0xc1ue020i4pA9xQROi
By1pnPwyYN7qVm9PY5qcte3Cl7YbQOA3d2bxK8LltTDm3G9lCMSOUs19L/u0RCDTCWnQ3+cG4E0d
tC8tS4HztNcVXRMNH8UhhYzvGysi4cm02Mk4IC6KIWhC0soFq899AJO1yxI5yI3TRgcoNCjehYpH
Is6Av3GJdUJWSQ4c9XMJlh8XiiOj9zLfyl4gKQ5RNqg+hsEBXyRkDnIWZydMvdw6EEP3GVqRKQ1J
tfaMT8U/HkqhZQsPwiUBK0iSHITJLW2MbHprqCNIDgzL+MQ7BElAzNqsSmc8V9rlE4GMoqKhCSMZ
5HpyidvKDWtuQIfYM1PmAiYPlBFd2zjQ6ovOSfKrKR6pahMKy/SCNVkoX5BhpIs28ikKJb19RCKk
qzZUFN/VHSsqL0m+aGzCgrrcNZNTtmqM09A0pVYEyp5H0R/8nZowT5oRslSJ7FsQQIKIg6Ohp50N
0pNpda8OP6DiT5k/1YcEDGsVIpBxm90bhyEQMinrs73QrEumaTZd7VpUx8L7v1RMtH1eE6qm4gbQ
kucF3FipvWf76xTh1851lZRNrYW82yRXN3x9ja4Nax1mOz20VpFfDIPQQWikclGKBUN7vD0rF2TK
zPsHi3gOx7g9NZFaStullkCr2mIdQVjtOsVE+thyCuJAEOCSjw1wZUdYvrIkrGI1wRtcVvY3k6qm
VLmssJdPBMBRTzznzJ0Oy0YaHCmM/Vczbkuq8DfF9G+Mu5zcI4KGmidJe+WUtlxHjGUiYDzwi+VL
t5XNk//pPxJjn+bjsj64oYiNhNkJnWnqOGdjCoyAaTrHdmCetyuJQ5LC7ouc1pnShHM2Fbo2O5Ed
Qj7JMn+frrTVBtXNRsU52gfLbfAtJ2lZyzxA7pAu5YEJJl3JUJry++SaMd+L2RByri4BnJCgDPCD
+16HkkD3mXfhpr8DSf3dgUFpwjaZQoJLpFr1R1T2OSJRPjZOD3LuQBSuNqGSyj6enAdeqzDiDJM0
6pQe6/WokfX8EhjPf/YUf103JmpJ4TWds1RI17q1yv9oAvMP6opi4LQJedo5tj3gmZsy8YA9UMrn
u4+ve38770BW3E3kF8TcblKMNJINx4WCLQz/DAbCFq7CKRykE/+jucw7pT9ue+jQjvRglnj30eeK
SEpTjSpWy2ymG6ODIuavdVrGlpsvuMByRwLmnow6j1gDEKY6Pn0ScE1cqO0BTzL7T4XSyT6weiHv
g3vqDrTPcezMBSBY0ineTWNkg1NM7g4OxVGMqJPdROjTX5JcIEgCe75PkXbagIsO4g1n0BPAdgRn
EEcx9gCZiaFxZEl3GSJJGVfmOwH0VjrNfjR9/15OQE5pePVysmQLHZ+v9ckWpdEMO0gL4OKfqAgZ
RPavufM7zauRFhgDBMoUEbcWkXCtO6KEog8P1IRV62uWZ4IxxRNGddt9Qms80T413Ce8R7dHHiOi
zcYr2IdDPr6d80hv1Zym238EiZ0fbviQDTHTmlb77uZMZ7qSmXnYX+cbeXAi+EKAyC01SlkIZcnT
+MRcv6eH5el6+dfuC0W4VASRLh8FBunkw7ofZb945jmLPKsc2aBuIOWwpsA3y6oPrAPaoMPrvLjJ
LxZal3mpoU+q+WQv5i6LpTIPNtoPqrHzcrO5Kxkr7oNK3VGz1gzu+iViT+9fwQdK1iCHhQ9+lwhj
FQPN5m2XC/Y26K1xcboeqz4vNqpj/j7AobNeF2py752rANyWLNKwrh40R3At7Z9z3ydaugCmciSg
I+SV20eIYZxjsdPOQmGbW0S69cpfgCUhy/BBpCSDxvkUN38/YSJQdY3IBsB5k/Qy0TyLhA6o98fG
bWHKsBTisC0ueutHnvsKP8IAKLv/4063xAbRMYGV2U4RheGdZrVcTVIfdBO5a9GRd9Efc24Sn4Jb
+yT54ewAkTMLAWTHMfxoZ79UNGK2Btn1sPgWJTcR43zwD4R8C06qOnphW6O1c32K3JcpBoFLoqNY
2SFfl/VVeUtSHOkKVDtPwlPk0Mv+X4CWF6th4Wb7soBZXYWEy0+M03vpYISbBLhtns8PU4Yc0kKd
XrbkMvVhCrRxbrEpbiwyZOnvi3TrtibZ8RhkuCzTUP2++xSH4/rx4KxaDw9R7qtCVU6m6AenGUO4
N3YAeZ3goEKV98Pa1lHCaZJyGbEtweo7b/NgXcaJ2LRxrbces+Mfob9s2HEvTdGYoy3gWqQGKvk6
os6OanIVgA5Ji/IJKzRvtjMsS6RD5dcfclm2hfoZSqpyqe9+qsrZ3lBoPss1b44l+mz00VWcsfC0
PLQYUqIhDJttlFS8cSIm6ypVm9mMMUESO8XAkHc+dzWjO7Po0NxooXTCX1V/oa8AtUTXn5cKI9E0
fhYFukt3KJ2AUaGeVWAVUvkKzbpp/QCX5DSRRtqmr9uCai8VK+f071DDjUXbrtRGYAPVYJvdjLY9
OmSuEHiCUbtzo1yqH2EmrtavWrW2E/bCXSA/O5AY0XsHfa8Gs5PRb3a+pX+as4/LtIBPYle2iuB5
m0VXwjeTQmd/HBWuMDB5Ig+pv43JnyoBylwHgG7xxAUBmImftmNU3b4DYJzW0E0LruArc/rux1UJ
aSa/z7LbOm8h1BbRyS7Psycqa5BLBI0NFy3IfcjOyxLo89hq3y7+DlOd2ZiKxxNWOjjbrtbGW1NV
vQRYZBhSTHED0rHOtutzFJnjnoimIL1+rowRlrCREB6nqPbyfUd2pX4icmjKcBq52p/IFd3c4nto
miWKex/enNCuW2GmENQEAxv9G9WAw2y7uLaikZab3MikYJifakK9/nvDiQb0F5cwCfJKV2MqClkH
/WN3khC0rHe1xYrjaQaRG1/vnRPiJbhEV42nVTHo28FGaxUb3dyfJVlkWVPin/Jjq1qJNW/c+DLp
MZMW7YX+T9rHJi9rvymEXoykykycQQYE+9SkQ11Ig3BYMWAdWXRDb8AURG1sWdUb2qAauZpUaq8Q
Glo2W6qCjwcqoKhNupZw/iKFRQi78R843fhPhZLKs9hBpiTsr7HLfDdfQQgsxzViFMKBHSoEzrgH
QxKX3bUMPl57xAb2RP8qcFt1Q+vK52Si/Ox9wZPTRwFb1sNLm4pbC01D3GWpjFhCIBFo2ixVRwmS
mXROVeWHmwp1IROImJ9vdxcztbT/JzLRXV8XwZY0qGJHcXgKAOkEmwEEq+OAiTtGHKFMaC+Mnj7X
H/E9JoSGxgnAHHp6L+mMWT3wJkF+M6HDs6vcdVJdjlqcqAJhxeX7Qf7AWarfoB/IGDTfEPlIQP8/
Syxb9D7WOOMK5/ab7aw6Jkx7RHlhI8aAxpIra8a0Qlg8nd05FPGYq81a2L7pmjj5gb2JABSvfei2
w0mCLOLzFz4tvtcLZZjHwClN8rhaDJOnCLRdGbSylkgADhA/oduRwVtYGeaJsfvuH//Hvoc8Iqga
AOnT6eObW9xFmXslp/U4a0ij0C+TU5TbPsuajpIVLWdMLje2Nd89ZPPMu78JdPPaRS8psWzXXpks
y/XUIfFicGr+IS0uLGvnRMqEDX61jcJMon+dYlPQL1z0wb/240XgGGIxqGSe8XH7TREYAW/Tiz3/
Aap2TftWWaWrdHrOiaZUYAD5tFUxOZ5UMtsHfF6fT5ZX0t0Az94gEXUsVC67d8A9UX8MiGzT9MGV
yAcDCFHrQBFvKm7xuK23uYpMJhF2nqQCwO6+XCtWIs1CIcdA/aTLts+zdtlHTEwLjznRnrKFYlnE
8au+LSaN9Ma8NDYPCqcTtD9iJjJsIz6Tbn5gIp70Vt0UlZw94Hj66KRHZ413hekfwutoJZZiLTnP
iM6GhKWwkeV3XoeveRPNp78LeWnvyyE7DS3zDrNCaEzaEIvB9Ae16pdEBUy/xVobycQA9jhq/OPg
bCOPHCtHZjenoPfi2RrOL2tpN+7TfpeLLd2fSyKzY2YyqKvj09g71gK9TyOlu7ZM+gtIszIsCx+N
e4cqdUcjZWxIctpaeao/RcIfkCXgcxWjbkzCFjk8wH2K+IRzG67v+phTzqirvOpv3JoTRb1ZJmSY
g4fJHCWbvuq//oBd+sPIZpP+ZKqyhB5crmgaaOwzba+D3eEuqx++j1m/oCYGyhC4Mim8Hk+/Z05K
MCNOYEhq7cWrthoVqooc8pU2WzRgV/NY2RlQc9L/rivmXw/JEixyIK4RdXyQKZ4jjavFC8AiJzMN
EO9xECCt11Nz0mX1gln+exeg8e5pDy3EKCALBTbMZ3nwZwyjuCXroFxVfDIU0mgt+FpwY+oQGm9r
6v+bSvkmlUdtRxKSNOiOqV7JjtCipeiqIKam27Xqf/hhsznr8T4sx+LUvw/OCA5/ncoSI7rguwXA
mJvbXBsTEDJSpZTmwnVZiRhwH7d5mPTb/h8Rl3BMbd7oI1YAlKU5ApjMxhCCrfdYvRGzwcoYZpS+
qSdqF0wYnWKK+ZQW16kR865NV/ZMp73xNaOyt0kMMfFuKSRuacDgUtFgqtabVmjGySsbmhTntnqx
xHgN3NycmeJXizCoD61295MoHC+JmAliWLfE+VyFX5WGd2ZDYJvkCFVisxdqpOajEI97u7eDduFp
w19Ns6UI3O5a8RmRQn76OvEWLvLQOUAxLQ/8I7UJMATvLo5JdpBcOOjoNMN0eo4wYbuEnk31dNIb
HnveVgZ2K9m66PkINA6KF3o0QxFb+i6ILmBCUgbyA5dUaJKjwml/eoBD8ceEpC2qMOoL1XaxrG7Z
KvC/JlFWU6EWSqYxB0tTwARXZj+sjv5bM/WXUF0SMZYDdBp/Tu/MHQx8VRTz1yVfYSPIMpNz9/zC
z6zSCMQHSJm3mkiBURpA7Tm9qpU+OdlB9O0TYsjgps8Juqtas1WflK1KrEoYkCup7U9s7lqxngK3
JTCV4rzjs/SQnWcLXaUwODRY0Ct5qRk0XDkizKOreDbns0OSIll3Rq+yPW+FUZs7FLpOh4B9U2Ap
9s3RsxRqy7pp3zkBXQHbgfNBnenptuaWxS8NmIX8vdgXC6S6MDnsXLYpqBCtSNHSmxHoCLTVeKi4
bXHrWLB7+3jXwGWW+2s7rAt3MFr4K5YWa9Ssv33yvoEaTA6RrHTkuodo3KuA4jYFYROAf8sdJe7Z
CuFu2HfBV8qkl5+h6pDrg8F/VMrFctrk3snWq8YpZYuIOcby7TsJ8s4bapBJTtaxFwF1rKQzBvxA
yQwJi/Tm85FJDdo7m7aXZPvHAA8Nz5s7yIRo1ESHARnwMdYok3IwlFqKPiG+zBjHkJ/16x2d6PEV
IhynUtcHol0NVE4u2el/zrCgrYmtIGBM7ZCgmDrFjIg/0ICV2NHm3NBhcvE5yUPrd2qsNqQlEtI0
LDoVM4iSNkWM2Y7q0GWBUwDjYGwZKQeANcTIUnKhICjjTtiLymLZABjM5K5VOO6w8Fx1lNG4O6zc
QhyE1uQKcIMEu/5NZ6y0EjzlCfij784Lh/daQn+4gGybxaEImM6WA4v7mpjuPxyieo7oxs+5zIfV
CiVa9YKFXHDvOPvJh5SYvZaR2RqviEYbYK4x6ujo3pMDpvNVwRzvsG6jTXzBv8eQrUXERbILxY9h
U+3I8y0PMo1OWdlm6v76XjZWMayAmDg+ySqNA4ES9Jk3MOtzFGtDiFnofbnTOrsQ5iHypUYF/kwg
6YTPfFQziDCkxIrI90jBwSGaQW5EDnZmTB0POGpMsiq46ANOFbBLD/uprGtGFU3jdpWTPhksip9U
YduOxP5jDZqad9nqHaYGT85grXw7kkWeioxrrBUIZMAOIryJAcaqgPNZ2KuB6Z5EQeEae+zNgebN
r9p+qRd6o4JiAC5GGSoEakR7u+eciwNNNAEigLagTSYcYV1eB9VhW5SpLJpv3eUOIUO2Af3D0C0Z
ooSjXB5IbR5gw38gJaqnl9Fos2HrEXoCy0OexEVe2JV4D1Gdk2L2fi0ioPpQiDymXxhAsI954EjX
FpHS6pbgBGuDYE4Xr5T9YeknolX8vVNlyV+2mlWBeuWPCrsX3ZxW1/XwyYlpL971VoRYzZQDE6xe
vRg7WAy7gxhck10D232CRLn0cwT+vxj6O/OG5MpichnGwy9RFt7cvmAah//2rfSladlVOJILmD2V
Y/c5bdw4jxBZKW0hinHdAOywgLJTNLVryHStw1P79ERgFrC/zmObYv6RzmGc4YNoChAVHrv5tkG/
QuI2GP+t0JoFuDA3i1itpRFdUABWDvmPU0UBx4gH2CFXzudgUWyIKAY+V0+El2DQv6HeBCNyGiFt
yPyJ6/9PWunMWUaQLyQTc3F7g6NvRd39vWoxSTcD6ahzcLlwk0qilpc2bSmTvLnbvTSSCC5XAPUd
+GTsxmsMCnE3C+sM00/vkIiL/cekzmjlgEu6zJh6zwHWt5w+YIHzqYrDlD+GiLI0V7vKB4lpjnLO
H5m1IXI9ziUpAW2HIlLPZ6uHz054LHrEfK0J1ap1pE0uH/BwYoTqjLsjk8XQJ0H/kgv/oQJxz77G
AYSvRMHVx/9IAFDs9OThl2A703gw4Z1aVws04adaw7DrquRepNLT7tW+NvYA8dEfzvbyqVsX2BDB
2iVk9uq/V15SmMnt9ZXBhr7woxUxpN6i/TN+WExiM6UF/JhRobXRf1j8J5P1ZSalX80xr73mk5B9
6pbRY2hRjoryxuqfH7nl/Z8rXDQmdh0mAL/dGvIuA3Z8Id0s2ev0T8rXaERLEGdz7HMjkN7r7HeL
blFMN13UfmDbjGqcTZrabVIZwI4Fp1YYa1oWD2ZzeffKT0gnRb4mPE7hMBmnpr1mSYMSjHDpc/sA
74yH/q3+3KqG7xiAB4fRWjSb/h/Fd5d9ri3jHoQzm44jQaN2SEmU+vZWzalJtDkAcL71DuiBj6dZ
lJ1xURBXuigba/NQGhPaxRGRR9blYlJSODKMboP08w5HMZcpI/9OJ0zwMTUp3YRDDZBPqIMKgrba
luce4VDhrBD/jfyi4b49q9EydARLiVxqv/tpNyW6vkUhkVGkNXE1snAJctjaPCGrDa6xVfO3/dAv
Dnm0CjEQWlwC2JNjZhXDM2qW34AV3SI/n7o9RIQzf2Jvs2I2ceiT69JaIqFzSGxLuR/Et/fwXZTR
pGKTNUaPPey5rDsxjPGybMuvhH9JIPfwQhJlycIT2T5hhZH9h20bEar7fNBNH5RgH+iU1ZIzQAiW
7ouPiIUtWhE9QfAcVgdk/lkJzh89DRZmxhFu/RWYNKo33WZsAINjd/l8nkroiZmDijQSJXiDr4SS
rwzGMkRHxskTsrdDjH+QmNA4G1x3nN2eSkMR61OBPIZEulzeR4kNq3T2J+BonffT0IsvRH8MCSjH
Y6K4/3LG3DNyKH5CDY4OQ15jDVxa3ivsqfvaiprUrq+5iL0TVXmbR93MWXaIhHOuvhPE5uXERFWH
A6hSeWpd8X9AxwSPQnh/BgoNs8i4Z4ki3UQjdEMqzQ/6gpRyIzPkgTSxNEgk3We96OmBRGfYpmll
XLseyxg3d4o7OL3EWR+YDtf2zxBvvvdvVp6/XhXqenVqv1GZxgE/8rZBWhtJ0gyaD6cgF2/tSAAn
E6/pkkoazsocWs0RucAXH4CfiNV849RM8+gNTzY71zA50u+nfSpIT0aYb390RRDIpO7rW+ifcKQc
EFYdp3MH0X8+0DsVs9zKqqP6zlcSoSS3ptbu4JWXUmvFlI4hgb+qywmIeVR51hMBd9w/lhlk8Atp
CRc6HxrXFlmSOGTbqOYPhl+4Qt3M5chlqTJWU/U8K4APwdrYXYs+k2fg1XUv8r+p8iLhYH+yrWEw
NlMI3dJxG44twzv1p9HKzS6SgZvIGFiI5JGrzjq2oCIZ+MRifZduOzY5396ORUwUnA7m9Nkq5OWL
AiUSrJ4VrLsd6kjdwuT1J6cjD38RPLQil77tMYXCxLeFLck/P0dSpwa2FGr/XCYav0MIDrfEW57F
a1WbBtCYz/Sc9R7z54sifJhq7KSwSYvVqeCuGYD/xAIdpXXHdw+KWDlrm/f4bb58DGWZGiFWMC5v
x1PipebRPvxRo7ESYEMk5XaNkoOu2Ih4hEaz1OyMzhzQCJM5Se0BjdyNxg/U49WkcHD9r70QzQdZ
sysDRJdGq3+frXcNBTn5IXmLl8cdI3LufpgtzoId6dJUvnD94xMoA6qLauyQ9G52zRezY545HLFu
gFKEtzRln4fup312ESZQacXa3/Qt9JMoHbNdk9g4R1mLVLR2hw+N1IFRvUGxv1aFaRLnsvbWAeMs
aN17AOGOqohFrXXQSPa2LYrleU/8PLOyfno/uXAn3cuJdGOCnXY7xtg6UHfquXjni0U+OyAB9/ue
O1oI3c1UlibVZcW1KlC3jBr+K95DHbHJZMKZGkv0UkHKYSlt2o4n2zqrnI4wIxlXPnEP9TVNQlGT
iTBgooRZW53HxjBIKK1m37oKSrnM5uy4hYAxjm104PCjFJdE0aFHxBTdtEgeqTJNC9G411pjML3l
VCplD7eOEPToNxVw2PxSaLMCjHwqoGAjvBws901qaX06EEtWhLYHtjrGlY5NFASPBtIQIiYkFLLS
41jURNl36B6O3OZyO31E52uHbk2+0KYTXFnDhPpW8elvGCpwEGYzRIZQASOkiDdX0m8FFgw5TIni
KKK0EOLsgEf8zNKpxn4GmGtXjw68IATFHmqJUqrLaKOo0ulqcYGxsmaYu64JfqpBgyplX27pBWLy
I0YOtiTo+TSSkF+l5/0B2LVOmF7vyO/q2reaaKmj/RJtS+XgZPEYDTE4HaKh16hln/NuFNVkoUY8
3cJyZ8ONiPCxAQCucHsbzPxrDFDZpN3P7DaogDQKsyEzJ7lTwe2176iYzLzBPOHKQWrcNPLydxG9
TTRw6UIADYMupqtPQhAE3kUoP5JerXbmcwPnf9i5QszmJBT1rPCtzYmg8RSnmWT2Noa9iRJU7RR5
jTRRTYTTeNq9gaDr+8f6Ex+5bs6peE9cY0iS3JorPGpoaY6qV7MS8TmGqqptDHgGvr50n5gdR53N
EXWsI9BidYnZMwPlBaV2ohSLZhanRVgP1bxQwI7HYfM6rE0wtDgl2gklLc6u/sOuvmUYVpol41r2
tCx4owehauTM/Lshr92s3ocMKNjiqk7KM+YF8kpQKCe8BEPKD5xMoN7O6h5oydm5mr2sAztLxfzI
bKBzZ/FS1jrOFIcuP8E701K8Pev/fpS56bhMFSbhTvo4QWsoLdj8PBvButD+XMmHtIeaMy6t8Qda
UdFHMH+ibL0vjR2456EaM2c0RuuFC4vUzYD9V0BTRDGqN2xhkrVF3qzB6RfOHWh4rQcOco5KoZ6z
P5B/BUe1pYyOPW4jkjHaKrFmZuE+fPrwrxRtEtHhgpof0yFqgy7ArD47/1txenIxnK6XfR2dW96r
GRWO/AsOxGTnPUvogcddnY5mUDadQ70euKNDnioudehRNPZavz8EUjWWS8VBFIYwCc17XoCE32bz
+oOwXHrhrHHS7kV/0od1woYnpqTLE0QS5rNOwPxg9AWGKfhcXDlyuXM9SuWAYs6zEIE3KdMmoOfg
D5U5ibrtv1kQfj0JpPttP2GRgfa8Gte1nOO3Uses2BCbbjMafROUBiVWagSBrkV0aD54nPMK4jaC
oILK4QeElDJJqQtb+pLdGMnFrpYZbVx+AsMAFS3lETWzCO0T+Awr5EFrhPFPnAm9AG1F9Xb0NWYY
dM3qoBy0bqXsu4vcPcrO+qZD5L298SD+VbLWmmXiYaoXDZ9IT2M6qw1f72uczq2bJPeF60F+hudM
+s2g+pd+1JS+7aFdJTNm7TIyUsyAZsr5odWKj4+yLEIEG6jKFnjShfQ0anj62mIyMeBrSQy00iKK
gZLG7M5N4ZWFdIg2lEiOQQ6KjWqM210a+D6ZhrvxQ5CsxpyVa/lqPhloVC3O0W8xvgcrTTHtSlOb
zHXb+d3TDxTM27VTtlAIelKBcQF+Fppaz/5YfycYYYGiPslSqVwYo12PnOMhN6+09Cph35jvOwPN
K4CG0ulEBGG64LLMDOzNKdN8ix2+exL6FIR31UzUTFjEzeaVFLk8cJ1dHzoUK6HSJVtq8mssa1zO
dqwWRDmTnSuVPK6vCEHrp7I2KRx2aVCkYLf2B8tAuEWLYxhx2ui8b5obkN8bSq6j1bZq5V6LYQEy
jHa5VHw5PIvOAUtXyFURC9K05cCS/qt8x2IAUcBL+vCN+G6mLpM5n9XFANrRF+QqJdE/3xUBXtOj
SI7iEmXCcMCRwV0eb32p+BXSPVpsWluI1MxdvON9UJmu6E6WZtBWaS6mi9uUckw2wUqjf/36Qt6q
rPrelZnAH8OoG4Nx3C3CA2scm2GEyJ91xfiK/ZdN81nvWMPrCPw0HRXYQGUoXXIRaFkGg57FnpNM
2vZ3uaahdWcpUeBxiQIqY7KHqYWZ6xwRRvICum+j2QXx6fQ47sA2Ot4bzLOhndlZxfVHKf0kolRw
RLQKuBgkWwu0hmV6Q5PKCpWd1pZj8e20gq/7w5ZNyd6k3TauzEvqdBouqIi7k3Ljyg6FThq065IP
BAHdkQOywSz5CMmlwmT7BGewJfmrB1KNiMvP0qnxjVdJ62uLv23Wwxp1SVD7BE1CrxixViNG8+GP
c08lNBSzZC6gF5Pg0VdIOBVm9r4gDtl778Ra3NdrCZ3NzZoxGAjl/h7uzOzxFSIvw57eFV+Lrh/t
kggh9a3rjz7gLGCvjZuxChTu20ECKuX/QBdzd4H5tskNOJrJDNidgVwgoQPb5ktCxNB+/dS9318W
uJeQMF7CGmSKhR0UH0FzUXO/jmZB4o8KosmQh4riCzg1yXuJWgts+UCg6dDd4l8uIKuImwG9xIL+
iaPHLUjXnPrHL9x3KtAugJbv205Ue1piqG/1k9uYcHWqeKedOuAJHDDjGPU0MAUU4ADzaY33l6ao
lrlqYJoo2puSXkTKDQ8gj2ijHqOVIyBmKReH6tFqMsiKDNOAJ7JaIiV+/Lhyui4MoqgM/SSAddoM
hgo1/jbjIKHspI8BVBJrfMasr8/C9kKQsY5V1XTuioTX4eN72VzYZTuw6MrFvWdaNu+rrgtFgxtc
MMtv+jgyTBV7wTCYZv/Rd6JTAEXkj+a9aY+K89oIWerDufTHEzAcqJRXitotH7kD8ZR4Qd0Phdrz
+J2qoMsPm7BBkXVDSJlk2kk4cjOlzozr5P5BUqCWBP2zHZPrWfvo5JynVGM4uIcOzwbNtxtYMD2/
Dp71u98MOL96HpLXMMlSdEnA1N5urcuzCPah/mfQolpIvk2UkpzFQ/4kXR0YJm3DOT6T8LmeJbNl
dNnTCa4NgOxiqUvXZPOt8rudEYrkzNHthoTPtiBZU3vpcq5bRPZBy98L8Rbd9w1V+oTr8nHC21V8
77eSgUzHYfaKwvAqXRqDv6TAkKnyPz6OCMVgnlKpZexh+JvtiTn3kkX7b4zQITsQEjPqQTFVhf2T
+OULWoNLno/PB+r3S9zEXwV7zCGz7tF7JKLFmGH8VGR0zNoK3mxmcMBWl7ixqdZtYgBARwWXWsmL
pireEOR5fwkRpfTVa92iOO0IsaP7OJXiDEaG+snRiBuqxrIq74graaMWdiXUN2U1BkcaOZjFeUSQ
/42cRYz0oEIx8sZtCF0eU6Rgmgh0MEPPfbNamRQUFoZg3k4J3u6mSGhtTAjKPUO6723hMGixeI4I
IZeRz8oHmJ1PYr2VCJ7ujlVbFSbcsU2QYkPogLa7LKIoUd6bG0w0QWu1VpgyF9Qy36jAZ1TlkvgK
kzHYWPasOQi2rXvfLkaKFHtZnyhEV0dacYayAFsKwCPTrXZOR7DBkjQ43kBCaQBt/bqpPXQivHkL
NMqYMyg+Mo4CA3mbsEKysWjQ6luQEBAuDlEGtoEvRR714XsEhyIKke/u2+h5F1Jttx+hW6eS81aq
dOJVsC/YC68X/bD//lOSRr2vQK7YFcXEUT8r6i8qMun8wqI6kSr+JEpgx2TyxSOvLNLUocYH9ZxW
oIYgFgec1/GkqYlnKeya+Sh7/gtwVv5z1WttcDENL9C4Eb8LsS7Hqp+gN26iKIdGuciPynPSPSjF
kO1QFjPNjwLOTzGyKHNUwU3X2/8MFhStDAPFRiIe/NbSZk+dSNDxeglkc3mqLSszKsOCMDtTs2YA
lBQumT33LaHZNdjq6GcB3sAfluz3aGQRy6pGRTgQotUAKlTZ6HJk5fs9W/KLP4PueBp/SycEEuHH
EFQOM/aAgF+9Vb608nF4AKybGCePUfESauoKqoa9nvA0UT7S5u6olC5wBLtn7FE2TR1pgbXYX7Qf
vCp/rr3tS3l9lZCxj6TaYiUlqkezCEZkd29pPRGgYUq+TzAJLWb3FOvZ3G6f/wHZnl/biNJu+h9y
F5YeG8FJRyEewM35go64ugnIRINuYMWPuKFSKSG1E8cqnfNKm4J5VYZiinlXvvCtRMjRfmQO5oiC
WsB4kULPG/oRuXQvHemqLGw7veph113AVc5CDCn7poV2Pz8zu5pbwrZrcwL6Ny07zaHw34JeiH+I
3Sc7lm8J6iV8gIXAZ4wGJUX3V6t1AbNo0J4pyBM7WiBPBvi/oAWml/aO7aFcgkAnbtOWrbpL3kTl
TUOPblx0x8OqbXJ9nKCR44Qvpl9EEdkxfj4f1uwaK0RPbJwLiSeNOC1xVrr3KfvVeaT5MDRM/mq8
4nDZA3EaOBPp3OfaENY34TsC2/ctdyGJ+0S8JkpgrRmkgG9cKky5ez6mUqY/Fxl9g19FZkdd1K8C
kSgWrlLWMedRlKlfl+jDfZfGGiZkTSgJ0/4b6ejypSDu/7Ru0d/TxjlRmwMovwHTpSup1ERyRswO
LQlDIIiY7mrvdNWsQFdFs9J1qkVdAX893OMzBA+MIYWkuXsVOPg5K/Cu83vs5rjB/SR0JeLtz3Vx
UzrjpThvKG3S089zNCYfzt+MTr0yLdbhXphjqtbCPrYU8UmR5fy/q6j3IA+AvUnAxX3hnNMPf2oa
Lxi5n8Af+uA0M6nkgpxMvIGnkeTu9FNF2dQFsF6WIZhjS2rlypz1h2qxqAUHY/2esyAsjfjgu1Zh
Rv/CdpLkf3zxecQ3Ppbi1pK7iQydYZQ/WiRJmAGqZ5LmsEc6xZ8/LdP7yPqqbskQr2mbD81/hgUL
96y0Twuh2tw+1Tk4lMgCSs5I3/ZlORUz4ho6Q/CugGZeFNfewyLtSfKWsLb+VfH6EfIZcN+9jb1p
ci2eKWPji5+AUysvwEyO5WRIT26DdeLuTEQ4lPVkVDCibWgNxpMRgGpu7FLdwroA56ecjL+U08cG
rmcgjtMyir+YEMVim0+K5fQAC8oyBmEWSkTwxzwyq8breQHJIz2CVdPvJzOA9/Y92jwuuPL+AOXe
1zr9hj8GORGVz7MN6d/zkZIkz5WVDdaeR5UAZ1I/EENzsz8BSIScx1nSavzPcmsOPP9bFu/LTlHD
xP5iffJrCpf0A6+hxKtfSON0burfvCK5TO2/ueue+XYnf9H2TV735uFJnQVSlit/FT3AHmGwgShi
tVl6jDgLatPgSWYPOXOxaQJcRGqDvTXFL3ETc2IvpN+Mlx1qAipxbBSzXdARNYW7tKda9OoP2pCf
fncpAFNjzeTIfzpiOb59IM7fM+wt4dH7gsquW+Nhc4NZWmSoYNgsrb4so+ieklyIyF2gLnr4zaNY
+9Xw52IXB2QMrvIelwEJdWfCdwydQn1yR2riMVoRMoHGWHR8gTJ4u4JQ66CPUKFrJwqBrjDR9QxL
71YkVN+apLBRW6Q0AWpaisvkfsxyu6qK4DcykMSbbx/iM0uhJvXijWrNqw0sbymenYT/DpM6ZbfM
LT1FatlkCq8hpRvE2qFql/IO2uaw9RGXajTBlBhyeByBphDj52FIEo6Kt6hWZ3iPOOnuXQGhxGqt
TE9hR+U6DeGYSokbnK84pSmuqPvpOxQIXfLElQ3sNpN2hC0QSeIT33T2/iW9bxT1OGYjdp00KQ5T
4sve7eVI1twcjf8Gs/vuIHJ4uwpQGePFw/EDcNYSuEWQL094InulfYlZDwqLJjY/E7RothLAehYR
xGUyzEnce2IC9FWgz3Fbat+IxZgydIo62KggirkaLAP837MM2L+NZGoa6BahVZ6KLkqZCU9P98sH
e13O5f7d7dDbjm0A4QIe7Ix8oheY4pyqNb//g7/P8k6EPATtHeZamRHbiXWYn+a61tAy6aTlZb4V
dgfDsknFgl+MuF8I0yo1L/uoH1hdHTYAxr4secZVW9AVKwb8GEq1bTBlcASwI0QH0YB26Q5gHr+C
/ZBDCuXJpDVQ68MHOtmE6D0SGwwEw+nT9V1o1iMuVAgfVb+hFc2Qo77x/fBhiAcmDFokbc/Zmehh
V/Mxg7xKNGRxyZTPHy5CWpYFa2dAOyIq1IddWdqvVh0tswqZZxFORK9g15mtSL8gGCKtB676LBQW
759eRStCZ69q3FGjCqE2f5IA/a8Zsrc1zwhQlNij5Hc1mLjMNbiiQIfqMIiX0RJGgXI9swAsW5vZ
y+WjCnCIPT2NMgnycwFSe6cm1IwZZYMSN3Fkq4kaqfW9qkadmNBjp19UarW/pXkgl98/fe5e0Bmx
ZsjmcBnxPLD8ClXBZdpXjK8kZHMXKcIGoCP7aUMtY5ypPuwYCtHmDaIl2qhElreOFoqMQdGHt2LZ
0br41swSeowj3NX3IRWbnEn5ZdX004Y5RWKMgrpGQSdjGEj+GR1JMdWBRDWEHtTnmDiMrKGoCBZe
qUY11bsaOQyoM9WSQTTWMjN3Wa/ZYLZy5lmae5IoYoGTw3qVlFPh5AbxyMjNw+dp5om2tFVsbJYX
y8bB99m8uNWmhUo9NC6z7G77S3XBXCc886fhLabTHoBhHASy0SeuCCxtFgFEUwXtBX33c5mmdrGR
S7omO6XTN0A1ggArqAvoP1Vks62LS6LhWXljJkqDDqKt1Wu2aIKZSW3v+DbYTRGD4CjdxPT7TZu5
YIN7SEKzcKZuaJ6gV4Ep9uP38cPq6ZbLFkBtiXTDpbibZ8uGXMQpUCkuSzIuE9mmEta04yyGEu94
C5daIutW7owCtFb5VhKOC4XiouLEt5q6l7P6+bj5tpJ0Q42ycC015dbp8qn7N5+ijD0bxdZ7creZ
XI6ZpEsnFzIsUlD0s9tYaw6zUCARL/mcw9Hue2gDhalmTOUJTd3tHRF9ggZzEV3jG+nzYhBOx7w+
Kdm63hVh/TjshF227lIQJqCXltHzLCtD7wykuYzYDloHm8rmOatlNkv0SvyyBNkMXBsNaRE9ZKMK
AEyhyw/YPtt4xViV+q0GZaef06n6b3e82pfCDhoaXpHgpDLezBN4xxdtvL8/8hMzbU6q0fc9b1mB
msU9QAM0/99fU9CX1qhGkDTnDKYI7KRQt8WwsWaebS7ZgM6khgbYvYtXlYjPp7THdD3suuYQ1X+X
LSa7UQqpWskVJ/WfZ5eKUjLxtZuFFtbBQPgXHDZOuoWzN4N6O568A9nmH+8Ue+PRnUS5pBA0Spi3
2pZy3IoYx0R/ZRSLCa4WBazRdUx/d2lBz9B57HxkmzzKN46nuIy1UlQhXVQXMPv1/oJv5T+2UUVz
6Uh5KO2iDTiLh10jQEMmt5y53ckpVTRQymZvqXMxJ01kfmo7THrxWdduUvs/4kwzZDyFvR8iit0L
B2/JqNDCkIvZcKxJ35Tblz7ELxZyYmiA4ms+AWPbEdaKXLhgnyGmbl1pz1pX6oaJFrKmkSZKeYiC
cf94Y+LA3PzQTrLMhHEfBw/bYQ1SCvZgJmyelkDUlGJbx9mXtz4ZU4zLI2qTBiHYfThoPypPEqXo
wvM752Kj1EC7Em92MkdCLK9dtpKDAv0VFwPfuPjDk/EJ5s5rfBmcLRn8pwKMc0kI+Z/8HM/d2Are
rrgqeTDjGTQv4Bsa7Bb/OY1xwsvNdIuNRD+cXD8I4qwFs/tBRP7h0+dAE3k74DzwmaLhNz1tJOud
h9/wzwiCzMz6kCqslU1EtS653GHivbJ5KvHzoca7iWQxhwZVq6cs33ME00igFs5jNt18rNY/cnTm
+ivThD8ajUJd9uSZrBXY4GBsXPAXi5eBkJwf6bjEjMnEVKfo9RfHp5tKZGZUZ3fXo293DzCvGHE/
R98Hl7af3PXAGsNvmAJfweLqtnk7TcbvcjIjxcWwQ8KC/+U2IUakoPHBAaAe+oX3SbFyovEUzp5v
mVShuQ/Yaz13p1KCJVO94nl+mCXUJ3OrySXbgV8tHbckEIksoioOB+fyi0kvAfcl9Pbp8jdtfttc
RtHxQokpqR7ii3UWFbWn3Jo56btF94Fedf584jX27ihSEWo9jAP4ArMmeA9XE21JlhIGmA86U31D
ugWKTxsf9t86NOByNslTTS8UIhiO+0GtOpzVNKpHVfneDo0pVFO7HMaJWf7NzD/7z/5TPE3le6f8
T+wwD1Htfbn2hsiFk865xNDHVdFBZrV+DdL1aotsixfiXaM0cJ7fl9aMhLV70oNRLRd+0D6BZ/Oh
+6nr/o0yp2DJyABPX5gtA9/UUdld/ahWrQMW8PJPMg7vR9zemqRGZUw8u1AXMjEjpLlde/P+zedU
8+6wqG7Krmv2MGNn0cjelmAxbZrA4ZuZw4xcaOY+tz7g9PTk7bruwgoqcXW+CKhmFLUq6Wdlc5L6
mSudWbxPwpKVm6/uueev02Bj7+owhu/qZTWCdCdoe98KliQx21GAmYTTllrDh0A9EDs1cE2GTjQu
7JeiGW2Op+1DqXTHL4cFeelJZPm1HV9uOBx+n6/brtpD43fOv3RX5iQTfQv6Mi/wWZFTMgKJtjRH
l1kyAk2Sa073LzUV/AgsBCnBsG1soPWuf2IJ+rdVpYkHtbFpau+eoShCM8+eRuJxo425tUgM4hfj
Rx9zks4eerocsDmUfYnAm2WZKYpuNoZIJB/imBEIcNmLJPq0jeIv4uFQGYKsl1mhblPEYVFXZqFn
VtrbGJayPsV6M+Pt5Q4JXw5gsZcSMmT1OPDA2v5mx5hTdPwquUoIeQ84ljJmaaWbsM2n9d9HjzNI
mJR28b4Cwiu0Dnxcg1rn9iuSVzxWT7GAm6iyRygu73YOKTIoFM8Jnrn9Bs7nO///kvR0iJNtOa4c
eVk5kLxFrJVC5/+eRJgwkXgf95YMzvx9W0bK2g3wArNw7+RMkLDgG1qI24/n0vMjHUe3bZ5FfTMw
8KX6mxCuKJUih1P+jQnYVEaRXWVh0TST6ncJf2NIr7KFjPjx4Yhh9UnsnpxqEweP3MnVYzf+YRGC
mPV/ITdLjllFXEH9OFJgPy7bMJmYkaxgCTV6KBjO4lV+CnwSbLZLSEGwlRjKlIDvlCSP5tPw5g1N
UCyYttaNqns/g15nzDYo9orWLjKTxSBWIUQjdRbRsuFb+KObZLvhx/rJyTKoK/GI2nsPOHht6fdm
wHNoP4ZX3+ZlGtCKPdu25/io4Z3SCDAfXMff55B63XLVsR+Q/VzjoG0yz1TyC/gh0xHcL7hzkJXr
trYbPqAZbmnOD/K4bqjaG60ePNdS6Rxj6unDoBAiBZ5U7MNBsrZIMxx0/ZmXYcd+HzJXRHLS0gj5
7UlePNkOECAipTc9I3kQ2jhyb7Nm7YdkQWLqDb0bQCIBAGEOXc+ZDOXsmuzT2XROWw2aHcjmVlJS
tk0otTiHi6KvIyDlnxu38SGt82iKGnYjbBQQvqulDMqlf4Ca3bjOCpJ34EGIfe6XF5y3DXx6I4Fb
ouymnXUCoX+t2TS1Xm2MCx52XF5UKQH7PZCjdHnbATsFicMnn5mBeQ3S7x0/Y0TtC40wyiGNLo1V
Vq35vnAquxWPGmIY8phgtrokS18/191ioGw3ycHCPVEathcPDdSPB/4H7N0XY5Wj5d1yElOiuiVD
AQ0MQUvQvtsnt0Znh0ueILTJf1BGl971kTUs8SZjVEjHV4Kpdi+SgOWQv7nvXUPMqq1z/QkEJBeP
64tH0hzLNgb149UqX7yaPQfnWYTsJtm9SHYK3t5cgFvdVC348gnnMQNLVS5xi80ZWSUB4/LyhpxD
H1kgq+eo8jB1f/I1Mdr3n3zYpuGf6+29Jfg3UhQwLjNgHb6vjrF4K7R/2lM8Hrpka+xUd/3H8uN7
EwjGHy6xzYIe0drKrAdEvnFdk6qgkQF0m+5I/p0E3Fr7ib3sDrMp+UIMIGGbgj1MRdzay1AyjBvF
49IIGFgjhKp+aS6QnWNuOuc7Ff9EkDYzd85YqVRaepI9XslSSuWZR7dLIaTJjO0UtRFbH8V8/9iz
2qzKvUNb3POjHYe2h9jVCLCePTb5doK2jKRp3BleP1g/w6pTXAlM/jjait3DZGJbtTjjxlDpnXud
f/dWO2zxX1+qNqGNO0FfXJzpcMGatxGCoPVji1X+PVPLaT0qLuwt6XnZKzONHjaOQfzu8dzURrEV
0U4poYVZdGBewylvTfq9agGtHky05sqpEao7yOppIh1IVAKkzuPrr1reUICKJactIFVZ37U0EuKe
XLZZ4pgqLeUJGREInlirYH6h3sawrESir/A7zECCYBlpKbKArJPmlG+W+RWnNHMoL3cyjtNG0N/9
sLgKyOczUc45AyC5EJF+AncHJ6SAiu0MTpcwwnBN9eF6vb1kopKk6Rg8Lrfeiyo91MD+HmPQltfY
1jRvWZOQwTHXQnVU3USxrIG67OOqlUEMlqw7HIKNBKWDqfKMPHyn4o9ZriN7KsGjeWeH2mOejSG3
GkjJylFsZMPYBUcjiF2A21jKTX9oW7+qyVLtJPADkwD3AMgagV8jx5A0he1fDXyqj7s2S/xBttpG
2UZTmRTcnvdost27+u9MsB+CUuZMUpvVCBNNJTs77Ijv3oWtGzRL0fzEjR0kkiwZl2DPJ81GcHwS
Q7Wei0xpQLJnsd5MzUArsFmFdUwKE4MFPy0NEFd7VsNpnC96WSU1UzUCV/pMy0n7KT/fTQNDj8v+
3+sNg7yQ2EYhLyVknHHj3/naObBrPAhWBn2oVkLDivSlU55fu0mn0AScZ8jt3zzfPxl36Wne3F5T
GmPm3EuPsaMgoXtFYh0s/mtzsREJsw/dJOmPVFTcOr4jZgHL6GCKR6ZgElSU4BLNl5T9xM8iuecJ
nWrCVfst9F7np5tRYgJZ4JTuFHeRqxpujFI+3ndcbpAGWn4/MrMOjUwQlE4Shess6RlX3hsYB2AA
3tFFWy5ZmAhQZgwMb8GqvdlprINAcbdD7XA8IKSk94IT38GZh+82yhYwzob8gTt9gtkJYGLzukWe
B7anqNTU2IWf3BPXT9dHhPkpNIISGCs3xKqoS+heKgF9VBnJkxEBm28h/g5ZLFJvwm+eZVbia0wM
0QX7xSfSrjZIYB6/kf/R9QEPc4+6invElixTNaW+GskEMjMSSBDjWvRaZEwDeDGMOyUn2w82B+ve
dO4oBTCaNBHmY/okL1ukjg6JjE/M8WTNbB2c3X6sQnZ6T4LNzzba4G9HEb5pTJdfHqNquS00e90q
RoSjBdyYhsdyVm/xQIXUS2LumKFMhTNGLp3s1NAIFUjIFLSpNaqZl65cL3h9CyOJwqJSzWO999+P
C6ozFnPtms1IwmHR6vm1PlblAck8Ui3Jh1tcYMwToHNfKj8rHB/QTIpQXoBUaQwdITokVTXaDzvR
PIx3bEm/XobzC/gGLx1NEfm4+vP0xFj5le8Y/raupciasuUahRJUPecZV4BszKY6S4dPFU+0Il3u
+9N+32cZy+vw1SYK2ZgySKkju2v4HUn03flK8LGCEETHvh+7hizjHN4kilKMIwSjzMtbfkB/YJmL
SNtBNHiE8K1RlFOKVy4L9cA7SGTLZm1IHdmLotNt4Cj97oBkgVjQQ7ecnxs78ibOlVzO+IwqKtDo
Kw+HL2w4VxH/xnNiL4makrLtN+lDg4GYki9UBhSRfN/MuHgCvw2aGoJIaWnF7b62d0u47Qc6ukQM
EJOJ31RAWG6iJidUSdvFGV7tasqMLdG5pHOaVHpLGc6gwJqNxB8cA9v6CcUHEJvcOsmpsbR5KiH+
49hUTmM40OsTX86ArqDGOhJsEwJjHqOM3w9bq2H4EUGJDH3QBEQABOT9NDcHsNVjYN5D2k3wQ2Dz
zDlbHIKEkcc6sHehyiECDsWfD1x22pONf8kVDWGtXOl1KtYkcDWIekfscJG8RhKNh0knhxL1Bt4n
CwPdUN/yy0SQwmBdsZjZ1IhhORfc1rT4z5ebmK1NxJFvEN/LR3GoQzhiMR4KTIq2WBZOcK+y899O
wCi0zbnHKj76yiaxp0tgnSNPb2MZYKQD6h7ZWtvJtKdMdHkCtoo7F9vlS9YHfjJ9mPJtSYoyVIfS
VL73q1LMmw8c3R59bboMksaEjZb/2rj6Qu0BVcD6BHi+vkUs2jkWLMONHBnbtKlygapGr1r4DTbA
qU8o3H8lvjXkJXdoTY9yGmwqJwAIUCDVoEMKyMggLvrHLtO7KjA0TSk3FdfgyZWcgqzmDvet0dcd
wHMre204xLXziuou5ODKzWbh7LIOdJIi//I1iXFTCFbD32rP8INIQQhs78QofpWDVA/yf87RYVfA
1S8B8ftVKk+CIg4d3Vn7ZiZdvufIedzvk0iK9E1SOxHklXfBVtlh2Jt+AjTa/meuTqrVIIslpF0X
4qjABjyTkMOU4Mircj2RCyHNEzFKNMke7EuchEt3YuDFWZvZpP9ydeso/g+FVgaNykzda1S8VBhS
qA4QueAjAUMMusL1xSvrdBtfvP6QJ9BWdFjBy/0L2ovxAwHoCm1x1QAJ50ccjOZZNb9Xs3GqVAGQ
l5fPmARFiEdZIzwVaHzgahYJKlxbVGc43codNhhGA45YK6K7v0kUzJzcq7M12hH1wfMBt2/XUdDw
uA3mFi86C7gFtBIAUS5BJMcWrYXyfXPBdzNl5IEulu/h8h4iLSmF/jgZVMsXIkz6Y2nUA5sbgrWu
MMQ0DrLcEsKI9KygC6/GeqPLi88Ks3g5y53GkMV7Zmd1dQmr3RoFecgNBbLldJszftzkqBxvdIQ5
4Hy7j1ptP91oQitP9eICQb3KXsFt5s+8TKtT3uiKQ7cWkUuQLfh4IXtzCk/hCn3Ilf27zeSMvwLx
sJ6mzW1SGcNk2LdAd0JJWeRkFN6HKprpNumtTXj6Erf446kJYbKNicS9Uarq7DnRPRAsZOu5Is4V
xVvux9lnQIXPINktE3x8OGne0a28cTDWIuBEGX8puh7R5pRPNoxuO5ORZEdFF8Ar2rf72JM/8r/I
3WSBcmCBRditbaOMS3opCi9xH/7433P8Opp7Ps2gsF6xA6LsxCk2YIBci0160cZ67O665c0UHdxI
2f97deK+7ugbYHxX8u+VLzsFrXa+6xkgmNTxww0sni0XnXNkWriZ4tEFIv6KIbx9Tc3is3u27Ito
ywAGp3iFizigC2sSGAKdWJI3BmuasE4knYM0cTZwwRaiuGpqhTKZN7lFDCMur9AhPaQVZf2Wx8RS
X6Tpwt4DbHiwFZZEsIqvlGUuIqzQv9htCjtBb2JGrbCILcflF7jpbNwXT0NsU2GpDbuJg0RZmmK5
TyzUNsSw3cSpjz9bNstHqjHSHnNe0dx/pTF7Dtxyyr6rholI7qgTBoAomxepNhyx+CVBApuY6rgf
vkRsQAk+480xy7QrHqaWxQ+9G/uYz0S2AC2+QIgSLL8AgHuBzR3j2htert28OF11g5MSh9Xl6CQ0
bTldgT8IM7A1NSUQZs2vz/JU+rvZM3QqKpLdnHe1VcwntK0n7GL0JCFsrvG96YGsBFTKsVet/mRH
IcS3wAIXQWdQwPtm/nSvV7Sb/SK5hkM08tozO/vZ/VDpN0TWGTgY+rnTj3lny6puGQ0KvGLZ5PId
HfkOoQVdhdnc+Sz7QnFqb3o9/ANlOai7tx07uxCoMCHWt/pVGfW6Q7r3Pj0PWvg+rrx9LRdjuTJO
LegX/31bagGMoVszXbz13A+uiNNUTEvTtG2ibPSIN0L9vK9x0ZNvwc1+MA/EuR3dL0Z+9MHovRgD
lSbdKdA4QCtGEBA1rMo7KVxBFQqcmEwHwCpLugwWX/HhaStRUXsa5V2DcxFfbMDoT9UNvci26F4O
86MGvMwpyypIR9E/pMW+mEL4HXBDhS7iMd+YSDdqv8s/6QDFfULBZ+CeSMBHGPxx038qzKxXJtkC
aLHlRnQ847wOJm6qnLoWkKHSUSRJtPayehNPu48axk/fiD5CxyvbRKYXT1xsXFC+KNMSaoAgLPin
Yt2y3jXg0KG18yh/AsPvkS/1UiOpB4leDZKv8ikoHaCVkdSmnlNMwCZxkvUeA0JeVkWbpgS1d9Sm
jxNoT5Y07oXdEMGS5fqUWk8J98a3QxrebUupwUNYS+kW4qoiG0Zo9l7qjJl5om/IsApb+BeZ/mif
a76TkPHE2PxY9Zl99FqAZUFTRbNzGlHssgF+YS9onbKW/1tUNQSPkXebClEa9l+1LRRTsgOBO1MP
4c8DF34GzfwyczJjWx3XNeWpTyT98g1MOa8iyo3y7z/HTbrDB0olLtnoYk/rqRrtNxr4jh3QAPDH
CJWWwsKIrFN+QMrZG8x4tih1rkbLFQO5yPd3EeCWrHD5CGEwm1cs1+x9Txo+orwN/6ObPZv/MH7T
oGvaxmho40dnCVjrHhQSPiuzLgC98nHy07ZnjiWdnsY5ziTIjRCBeQGDDN0XTjm3Evvu3JTRc7dg
LmO13ZeqHH1KyePfUoVqVSttW+yitN8hL/dhA1Kmpp5moz3gqyqqlNr+l0sIOqsvZqMLjxAxGt2N
X95N+/qjS8FjKTzZ3S3Yp0uNrcjoS8IWWFTCsBL1qD2LOyPjIrzRHTRsL9QekfoSq0DeBLw2MabM
3J8fZ1dbaCNz7SJFgGVd4xurAdhlHGq26RALxVZlNCTLvLtpVu5YNQ2jSf7B7cZlfNDU6paPIP0s
EBpvc1NEE948RNCH8/uDOj9oVZ9pQ7F/l10u3kavw37S8uMHZVHsWFcV/u3h1+7V8FPwfOgezEW/
f3H6reUhQZtPVdYHaHF4wZ6L3ZGOThCCRIUq5K8YX30mAQA22HGHrvOr/k7sBsXdHPAi08Okqmen
SDW0G+lRuURXGQTOUHVpIevT/Qb6P8owdQJwkVBAqEfdyuEPiuNLAfv4Kk45n1ae5eCr1YQXS1ib
k6RGhoirmbsjvLdjkIYWOIr656MT5VC2i9vqQkpDArSSGzfIsnQZpBvGLIXNleeH05z1CcoBJPFF
WV31v/3VHgDHnHEzQheDQtLpJCyKnxDipJgnc/et2/U9CDwMz9KOrLUfegICNMpIUzKFcclACM+2
kQ4tLj71cZZasolpnaji9zYdQXqkaKx8XucUkI6jqh2Kkek+kn7q3E2yTljbHa8YhQ80A/htjIQj
on+dklG2Bi3HJnBLc2mpILBDkV7WqNMXZMKDk8NoBEO76TpM3unWE02KFcet4A2KBPFn+8OxCKK/
1Bpc0i8+Jz5zpzQvZNtqSfdLvyEh8jggfs3kylvMhEdeMx/Xb4geaHhSANJu5MAr5pVslsHTs0vx
1r6etf6rv9lIQbw264mU+g0iFwsruxX8UVp2whHIp4zjccRnej0Q0gyF5o5StFDpeTLsYTcMIqAp
C2NwGaHNpRsVsJju0TBysn44w/q3yLHlFTGWQGr4uUTYUMWVsJ3+3cxiRnXY/mbdS26bVENXb/SB
SyHTdJMQPXZc7arfflDzW0APJVygAkZ2gWeKxykyAtxXezQUpDRx6VsFtPje+4zRwtHYGl4wz/Kt
lQqbjD2h4uGpzJgfTpc6onUKMSDGxVs2bbiHvVCpeIQwmwiJ1xA+oQyPkk66VWCAhDotdYjkx7CM
r9qcWDaSRg8W6lrAxgWXgGhSBHwQiCZ/ViI7LuVbzDPt7UTLDM8Gd3d6ySSkhFNN1AFRXZcneyWV
23tKwNDanqJXnAh85DOwhE+WDlSzSgeX8IgT+oZXLgDXdHzjuL/VTrZ/QY0RHiKQKP2qQUAmm3U+
2uKyOBnLtZ3FsCYsSXjshH6vp9JwS22l7BxHWeBctEMKou6SbD1kgiOOm8hrP+rD3QxSBvNoCyv6
P7L7IdJVnofbaFQ5YJ/UTIXSBpRcSYtjTVf3sVY8aIjz0fNJs1JDEMT15+czsevL3SHpWJMunKxz
1AlPaF/KxbUE9XdheeLw2X4Rpb+FbxRxc4sK86+yz2lB8dQGC8Oeb8q3GUGxOfwPiIDbtMb8xN4x
9MD9UWQ7SlVfFl6wRNLdRTVcKaTg6nVFzZONzCbJ1u/uJZtdaboIIhY3rjfq2Pqy1qOa08dFclds
lmcso6lw7GwvQIMvkSXXctVBEgCLnP5rYlDvQTqdecaxqXks00Us1iZu4gQZ7aqeUb4UtHzclJXK
vfQM2Ch9HpKRGP81sowKP5a7SBJg76MTeX+lg2wfxAUztpeYE3u1sv9kEpdgS1jNAtZuaxeIqFwz
JLYizOgwsUqKhbryfOxV54ns8YQcj9WzsIGUc1YHOCIolyHbp1F3sxTKU4tbnHJHSXuWVxfzuT9X
E9yRJICHiLXbJz9sPi+A4SnWTzm8RTNK7kHSk2tQ2closCw8j2BkU4XZxZ6E2dvwrOe9KhT/mPjj
UQTnYiY7euF0QrhI/CIASVCqXMI10WmQYBl2xauAdWT9yWVEQI8Sj01X+LyCZUTgUCOPxo08MOsy
ZFKagelTw2ADOBvJNpfrTq9pBPtKkNfBRFePRk93Tbtf/Vdg0orbN+e+kv91mywkyKVZ5rc0Mgnr
0/UiMiRMQ8IFcrqxrXPclbhI0+x9i0ZI4SeB0pRCx4XF7CIOw3us3nBnUAqAdVKd0oNPdShBqbHH
lK6J0F9XRnK8rbrpZuQhiI3FnDBih+36+JBGqC4GBk7Q/EYH8rSHfv7j8CS2HVy96DYUBOhBFdkl
3Kkz+27rhaHMwCJs/OmLkOJOmPKYEjVicqaQFJJyOx3qAlOObPvZ445aep8qiSHx/T35qFazD3mZ
8GhtOP1hO4fdElk7hBdKfvDPuYgnHWvgrWZalZNweCVin0qM2yoEqyTU6yQ1omuqAtCBqOoKf56u
3l5qjDn0PgdgIZIN+kVe1vuWA/fETnUjYPkspqwEhAriWghsbeXX/YKV4RVLs5oPwJ8mG1uHMzzU
TvoIx3xAT0SsB/eyXDG26BZVuDpBgkB1VjM6VtxEJo6AI3ZTkVR2+iDBQ0a+tTzCK3hzk7TqD+j3
AYgBldW39FMAEa03lf5z05kjSY2cfdebUEtUgtJgrRCkk238Ceohkv06UbP27MuRZHgbA+Y+yGY/
UKRzc5c4fSYYdDSnEDzFtz1C+HRHpJJ2K0IVKkug8oojSaylOebAsDStlMYNwyyK8bLzddRw6Gzx
O7iNEWaCLjv+k806TqHcmYdDmIpQ+r1f4ErDaMQ8pMHIsVMVhogfBkW9XxlR59ocuai65A5sx/pz
kj9EzmHmLwC9+Wei734DA43MF2+FSmNVJ3Bejv5Tk+swV23fGVqthxJhD84p8I2tW750MPzq3hQd
/Hq5l7V1Qf249iOJVRXcIq4siByVu0AYABC2Hr2EOL1ceqvKhitRsntgrtvGud1ZdWBPhzoonm40
h83FiUDL+XR6Zut1h/RjFh7qtLmiIz4xJFF+G+BFtPA0Hx5KlB1wFcGI6LISnsItXsjZ+fORsWtJ
J8xc6GUTd9H3xBNRNHipEjgUTCAfbfS3K02WDgTKmhNWtSdhj3ysDnp3KUwdpCoVUk+9gamnh99X
G4KtNzT8eUs6wRIjXwKKX0i3fwfk2vc1EO2y8RvGjueAyryfn/JEhkvuUuwtekQ0S5kzhcyvui6g
GWJtsQuWEEc/P6Mhvbp2jH21fXu6unCOvh7WGSIMxB1UVKOlgnneVWmNjnUrLSIJ7XCmIXgwAMcx
D5fH8Uvp9ddRsmSzQKZhJupDX1uweqfN6Wg6iFsz4V1+ZfXqI9x6bJWloZybPC/wgz73n3X6/qYl
JwFDJ2J2Q/FS454nzMrUKM89BKBfzb1U+xwMdjYnTSYfAy6mcTiVCJPkXL1j5DNRcA2fYlPK6NXg
djPI9aCkEO5HQ7UIa0jmYKjxsOcKsm/qd+pv59a4FbbfgdrhuxQbgRpBdmdQZwQTWCur2CLtNOi5
7+pBLejvEUocdNz+JF8y0XCkohzCcMQET/7bitFtbqFPLawlWQraZgIT5fwIYpCjWNZq5jBpfqVX
ge7WDeUdnkYPFAqxTVtYOQkQq85F8UKcSOEMReu6TF6DM9Qdwh6x6S/d0yH30d5SgOUWITTWf5ut
2GhEAJslyFEpEUMdrpO0P+oKHjweu8UzmU42nmoXtHwvMk0rCIfwhF5wkF4wQBNuXFTYMZlih84I
LRz9JEkx14EG+vy7Hal5ErMJ7TOxW4vWXKH79hzqZ6r8GTKzLmnVdVPOGfNtyAFMM64YSicrgM+3
Le2542RwWpChw1aEyMYeD2XcSypiZHpRCOv49GBEyK5DY6YGLZIIp56+yh8KWqW2s7cRWvgI3Jbg
r+rGbZRgoo7jvsJkC3fitZZ6p1QuhVIC4xtR1sul8i/ha/51qCZDca2gr9WBMG1XBMj+j555k95F
Bla4PDrsMpMnC/MEyH6njgWiC02teI/iF2Ddw8g2Q28YcVttm5QJexELrCv7zMGeRSvTbOHfSBFw
o8XmAVj/g8dI2+CmMf7Hg4a2J/WXWv6bG/bd8TGoxAAU+v8G1gOlORrQ5sHGb3/wqmmVNaMiXm75
iTtr4kwEzfYhgd7BHk6vg+gieJPLUI3hzRTT/adOEC1968g3R6DX6N9XVADhMyhez07BOvB+totQ
aGXSkdNFPhr9QMbWTgi//iNlnJ/HbcpaRNIHOYIxXT4dUUMsVO1rFdQdO+DR4EeeAUu6V5U4i3cy
E8jDEUzT+ArC4C08fjKBqDaX0c8k2WIFJhvRo/UBryXOilfRevdQexThglEEgUEMjEgyZNCsK+xq
u3yW2IgtQf3UMoXqzhA7ZHjshiIjfMyDDlmIKP7qUqHNlSoL5wH7UpYAwxDzAW4uBmjQ7K8qbw1E
EoxiLgvyihVqm4bLHXIQ7P/8QH7h3qVYUlylCD9DM8+6H2+DUjq2TuFvu/4iWLPpuZ30MUyzrkY1
p8N/hxoVtnw7NQlXaWAnjyDhRfK01BWJdZTC2wBm9SmkNcoY1RMssCfpQKA5vWkf6PjLR23QBwqK
fS6l/mqtrvCtbC4Y7e1TNi6K4nJWWsabXEgw37u2V2GHYhDT3C9va/SmTAM+uTklghwNYlWmg3NV
5TkNJMuRWJkrqSAQhoY/JFi8LSdWlV877dFhUSidFP7btKtV4U4tceMjD8VjcBMpDQjuZugJ3Jyo
+ToraQxvNuChu5JarAGocmGOqmSdD9yKfkBzh8zPKvbkGWUqK7BUCl1TPvBJZYUUylvy9PkgMq+8
LmehURnaj9L6d7/CidEBHSapuzUfMcSF+LxkXKGvdRqaRDlEKbpBS1NVDssuKGZSwFlNZ/kUUGaZ
acTYahW4maGqFvcULNz6Oh5RinwgUQV0Fd/PumFeLACUTFhFtyuEb6xbSl1CaLEljILeH4OGuK2s
3uDxcAhjc1r1aA3UBoUCzR5Py3Lod1rVh4Oz3xs0ymCcOJgcw7DKtcYgkgmM1NfodSSyr2rHw62n
Q+gd53Rt8bGedkshszcCYxmTKcW2FmOelOcoiLJY9dvNNx9xnbZC38GqDoqfjnhvQDbcMUrc9IDi
nUaBQiO1VwBIUBwf0dkfqOcaRjG9MvgcexgUUTe1BPXrtuGj1jfTvlQ3DfiUpkRYu1SfmNZXf9nB
oic+mN53oBViNWlMlH+oFAFXAfLxXnc4lAf5i0wlLZcoaErL4f+P9Sovh/mbB3WXFub3WGRsc4qa
yk3ZOj+A+LdWyPNd4cP7dhTJ1jVUDsnsKx6MQzcU9TXgacN/7ibkOs37IxplZEd4O2nlzhAYEQtQ
RjJBwLa/NWP68w0ze/XWNHN1x1TEEKy1/zxBw4yjK8jQH/et8xKE6Gpx0YOvD/JXTaWqHnzAMbkd
PPb89oJC9YPoFOAv5LCmzktq8kY6toT6P3YLz7e1EiXDS6taLFp/X41dqpzaoiOXuLEOuo5xKRqT
fQPXpfIT06IvTZKuUwKzyHiIAWZMNxe83Vg2A6vo61eXG/3nSZbmVmEJSY6blZ+T7GUrAJestwun
hSxSnq4y9bxxu95/GMvlwBQogMsB0kxbAXRDVKj+wkF1r9nDXsLeJN3AUSwzOYpUQwPG5/GvynsP
oESAAICJrHE9zT6Ys1JDDWWYizJIyjlAEeaoaIZi9eUux6VxUzL1uIyvWdm+6tcWt8mk0kastdT7
4IoUmzSMCZ7BTAXD9vDxxTSSLLFrM/CHpT9qrrqns1Tm9V9/s7KQqWCuwNl28eGqc+N+DmiPOhBu
ikMaKXOfyc+JQBP0O0zzN+Brl7pOGcmvHQwzhkntLQN92QlMQ9yr8FoYzy3HDT0a22TYJI7jSsIo
VHhRw+yUz4+NnIrMadHSfp7xoE/6fP19/MwsbNIVJFK8erheuYP8riRI9pTzfxqUStqsPwoSfous
wrGfz8V0ByWJa/v6/eh7AzeukyzQgOslRTTZOIIOneEYKNS3U7hp2HFctOTOREsyRMvfidmKZwuk
zF2W+LJzR5ggnJF8f5xKXDCYoVN7wjl5+FZjjZGuc1AdNxytEZ5nqepNP1Cq1LNNZFjXk5UbpZj2
N5H6Ry+WHzRA0zn6SUlPmNXQW6ixUBvKxB5OoLHq8Pol6Ed6qHYTnRYPna2RdS2nkBEGw0Fkxd4i
UelzAhaiNGXPIYSj2MByF1oxZPv8yrbvuH7bu9+2fX5YWqQIE5IDrnEFUfp8Dzb7p4SebLhvR7xG
WJg9+IsAthJFSftBKtB5EbZzrhNetAg+JZnepBLnTFL5p8GR9Js9b4yfZ7MWzcELUwry4kMg6VTW
ZWxwOBk3BK7/xALyNnSXkux7UiKmElLdA8kG+G0Z1KRnpdCRkZYxSxkeilyNpxSMheQPhB0lRCTH
YdL+Gh7OUJzMwvTW/MAm/LKUDqf/6IdWg3zgQd01+NImBJTRG2G/ExE+OjQ02tNdpXy7l/oS0Aoo
M+dLiDae6ZlZNr3SduseJN1MsBrdMRy6WhV86d/34vszFpP0NkcHqKCicuigNgNWBN/BKXyQFSNT
PRIT/BVwV/Xi1XiAt3dWXu9ASSjm/os925yE93w5JKkQxcwOYI6MIDX6AaIfqj40d3l7ssxFm09R
3S3ivWACTbx4eyR+jOMTp2nRTkq4x0+P8+A1d9wCBq15d1+tr47SHpR9zylh/z00myixYm4aTLie
WboZThdfCIRwZHxrq6ksOlEAcR7O6LNdCRLch9YboE2AjtwOJDlt0L5p/5QmDdnM2AY0iT5T7mV/
mSDjMvGfANKHUR9MDaNVYMIi9sJZxRm8/+atTP3d/pa/eMp0OX4KCQcxglA29I/BNo+u25T/Seer
tj2obE+4PXE50w0upyiGuhmrzWJHxtAoWKUnEwHN6ILPXP9I+dU9oJwJ2XIKLAA+bmgqA2/jggCy
X6PgvaMaYBmEIBXgIlKOOOGF+cJxjf7dihLOuRNtrHkknCtNVaG/HTD5pnyUOCBqRhUwZMmYqkqF
1xbCsK8w5cxCvaZI5plmNLN2YKoVDxW5lhjKz1NaRaZS05b7HzNaoxzJEAkeOcAK+HTfA7ut0m2I
gICf6XQo/Km4OjnPB4my6hHqHyEdD1zduLJdoCIIRV2b4Ma1IIlljGeSdPTeRd3iaiG5vQrQu2Gq
wPWzKdZPogdTZ5VP5P0x5iw7OHEgBuQF40KGJDJyycqFFcS8gzqYGvp+Eu2YWtAAVeNtwuIPCwqw
cBOqRPWq2VncauVinEfxloRHJ7epfznEl4C5HL/HLbGY6VcSR/okFuErr9vqBoR8CkoQm4eHk/+M
9kFaHT4qRy5gAforZ7j/fcV5ZCJFU5ea37v94MeIIYddCanem7oVz554o9MqH+oQxq3lReMAhxo0
O76rvONvtwxLRrGclm5Cmsemaxa5tAPegMBAnbYqP84a9VuJ8MnDwFcLIyZGk/Y0fMIrFxa77OhW
Mxm4JN+ie7f2lJztlys3r2KVxmSdenIkBz1ymxAiyZ8JurhLD9pK+fxqzgDcGKWZA8XtaXfKroeD
rmRafBFA0TLy8s2RyisNMHAHYaoSUdi1QDFJ+O/RJFGUnXlfBGXIqt5Tb5yQLpEBVp8mWWjPjsVZ
D56cIPAT2UmTiEpzj84UpU92uOcekx8V69n8t8Lijbkz7RB8y7+z5lOFyUXJEuBuybESqe6AoATf
PX/c7IoKiZRXJNEHnvEYRlFss2dwZwgetsI0tFsbgD5GFBFz2XJspM+6nbzvh/Z210H/gywJPVAL
Rjb/g5lZxaFGY2wyDCEixJdaIR9oBJrr23x2a9TtOwg5L/ug3nPdmFjzojb6ANm1zkn5EntKhrse
EEi1U5stQhT/HcWSK5OsnMKtY2Qu5WqHpTu+zNbXD6jS88xz2MmN2Qua0SIt4/n61KVxZXVjfmmA
J7rM30rmolJgTE903R0Av/9vEdXGNIdHgnPN74Oow96x4mi/REtgFSLCxwR95msf0+taUrrGB0TU
W3fSvM6LcB5PWAeH1o2788R5W5/tfFzuUbqPft/OJj0U8swr8xjBrCg6yQRhql7E6wJzXqkFMl9+
xZsMtWTqkfRvCytZPlqYcahOnwzf7TD/mzPZj6h83ywCyRYbWWamf1SFm+U9VFNI1gEAh1gu6vuW
cXkE8NXZWSa6ukCEEu9H+ogXSYxr6iA+2B+vvlqO8wNUJPOA0av7vXWeBjXUULTd4bgyycPugI0+
XwHnHm+/V8FzJUyHaJNfAPe1sqHYTKm5vZUbue1xdDdgjjRqRjs6G26orO6zBICP7D78KMJiFDwj
8oqlDE3F/OqllxLBEcnoX8M8ih4PvrO6JwTF6XT/ClH6flweh+f9om6MbEXiV9bbF+jEZiRoUFq6
hWegxWOqKUp9KRIsexesulRqom1DuPnbs+g3Vy5Lz2ImsBj0niiV7fJrCpl5RoSh7NbldR9ARvr4
t20vvzY/5Rtp7FlshPynfK/ffQ9hMSS4jInhIEyXNbgHI2S171tvkDHpl8EY4e0ztJ80vRwyzBDe
LOBDrTPjSnkxOXsLaI2GIKIeOPhzZEamZcy8VhKxW24NhiQV+TNAbKfsKg/rObKrb+ucRvPTTHA6
HkOUf7m7OC1TTBQENcxk8UqsNvzpcTSJ6CB91nIMhBITrNlSkF9H1BE9Ir3iM9Tv2XyN6G2oFBQV
NeoaYbtaziekn902Ro1HReFXHTlRlOLbzEi6FbIqLaext8SdFP0F3FBp5htP/XJ9jG7QvPoK+nQM
7txeEdzjw9mI/0CPM8Aap2eO3QVt4NuudfZKf0UYIGJUS+q3QHNsymEx3383/CkraRkhmCrGD4xw
cmSGxbXGAWNm4/jNwqDi7L9oCU/NqPYMO4tbsF+rX7AkVSqs0FCfIDPWUsHbfl9NZqhXtS/+wpZ7
j8RAyb6Afqf4N9AFGvsGPdzMp/iGItPotZii3mbNs67HODIxi2axxKfnayDpWYKpHQWLOpp+x8uk
cx3BJTaZtzuAgS0g03xXaFVoLzylFmzoZAa7TvBVnpx2q3rAcgDfuB9zP6GtthLcl2TWxQd5Yq9I
gsk7mtBr0K8MMFObzJentG5smGjsOpZ+++f5OE78fNfYI7jqOiZyhstiufC35eADS0m+ZF4559ky
1b8iIa1e9vaXBvA0I/1klIIgSsdvU16aQoz+0JgrZuNFvZpJf+DvOM5iaMG6ukx3eSnTc52y2tgV
nRyYeSmCfLirGccViPnkK5Bg9jS4Cz/hpDenDvyny8MLkKwdJWH2yfhqO6wuhV10EXU11BNHWqgp
PDW3MgeYHn6odQBlGil/Dr3IO5FbG9wK/XoIDJg0zFx1zpe3BQWmZAV8dg0I82GqF052nLQKK67f
J1CsYgtP265m5SgVNyBNFJuyrlFgfiucPRXk1spO7gmdU0A69Z6KnCLiA8FrfEeyv1BxoWPCuNEt
GevjPZQ1mw+8KtuusojomjqUIqZcu2S9KDViTkJ3v0pgo1lknmIkVzUOBAbBUHaDq/8YXNb1a/FK
FwtK1UE6pGWhK29Z7WGa/AhTZ11FyoXVnywkSoTaCt0+z5rGjKHvXlcdZ/oiY86e15Iy167eCQJu
qknoX1DbQPAfg0/V9kDvgJ1pxlZNMTzXyxiVXP33AtGJsZG/atMFM5dr7rIupzBZB3CyRNYHhn2B
aSXBVCOT6BwOXSBKlH1fbfRm+fXGGXpzNaEEiKtkMOST15w0Zcg/DXdCcX6QwcIbQOmITk6bLoCY
TBEGFRt7SdxPnifCrXKgogX14uJaXdHs63JnCUdl4URz3tHQr70IRKSk6PO5/p1jF5xlxFz7B92d
reOdqjdS1d0Aotf7TGYwOP+uzqqKVstOGvR2mkcAJJnZ/RgYbQfKqd1fOhu+1LtqjG+6lToHKqsv
tYfN+g4od54/M516HxmxRsoJhy4lfSuHgpPnpZmOF/HwJMmEojVDk48kpXOkQq358lkB4YdWiWDA
hCi7tMuDVuxyskkDAWdCw2uoMunPSQjXqDJZyvz3BD1PLetqR+EtFWH9kkIoCxUP+g5FXKgD7BB9
xSneNHPjh1XNupdesvcak/ag2lC6jIqFzCiMiHgkcAWnPEPtgxPaxcySEVmngVGBDyIA1cgBvHJr
VzLLA/b2vUz0W5CnPWlx0ErlY0vaaaWBF/S+o4s7pPWXZT/mS8rdstHmmrMT+5E7zqJZXXVorj+c
CBun4LGZeZhe54b2Zh7YcacEZPip1QRrZnz4EL8jG4/qfo9XDmxBh94vpe8GqR5wXA9NYSV904KH
LvLvtIoDLQoMcI7k2pzlXc72aCtFwYAMy18kLIErLSVmi1/PieeyrpeafZdK6sNrUuREp+RmjyiR
qHmJaERSIXMKKWXsJn6w0tGNSri4T07+cQAJRWe98qCTp3Ee71dUcbgBVnCksCO0Nh8EMakceTE7
EHLQz3pRYaU1CuVVf4rqnFwMbkY/Zm0pthemKlfJy3s7kFvAlEfsakfS88TffmvR8VGMSSTV34ic
9RYDKTtLWLGSyr4PdR6soNm3OVTWgI2yTFnQvhchRnn1fk2Et2yOidQLjmwulEK44nigp9dgrj81
0Jx+Lu7wcs/V9xW8uBUDKERRv11jTs31rhj44V2rOQbcXVCQxRfMT2mLsqvHJbU04spoDTlyc1QA
mvuOS1iR498xaJUyKhiK67uVgUhCxiGQOPUIl9oE2xDG3uClEECRU0Chgc9A1oUWWXsp/AL6vax2
g7RLXD4meYscBEwlK3XUqBkq8zbTXbooPHWUW+kRGXbAAm2pISYksdK4I/fBLcs3DfrococcWato
3JlQC49uLch+7tF47Nsz2IundMlFpuua4qA4VdYJwXUFP6cDULAde6vvHBrSD7Xpx6CPaW4jzXt3
7STgXsLEJqIZOQmp51J6ET5XsbH3lmIhmdsdm7LEt7XYVKDjgihWvzJxuj5QuIa8cedgNrx9Z7KX
x5uUNjhYUGoA0zPjN4Wt3evW40ewB93cjOmQgKOFarka0V45jWn8LXBij993F3joCTS0RGzVjYaD
15j+aqw+YD3EyIgjsfndTk3Ge4Coyg7aZoMWPh0H5uFYOTsaeVazT9FcHDGP6DCUbV9lAIIDaGVI
w7SuG1bb8PPr77vuq3GaQCF7X/qofYkek3uoH4xk79PRdbAKeiyoSXWBKXCgHFsu/wp9wUCvt/H+
jWg1JKAP6QYoEyyP0pGJGiOaAIBaRY9GdmfHfFiTN8ngzlOIJVaaxy1M64ImcwUG3Ky4i3VqhuEc
bwjr96phHM7GrGBLLuk3I6Dsdkp6iPNq2l7Pu1EluCp3AP+bVRe0OCCyPOHLKRvRBq7YcvqdXhig
rbhTqD+U015EVX3qAgi75We0uQHKn93SpY/M0K06jBxJQZC/YSTVQFccgDU8G8xcGOtinjX1oHih
fekoS5RlE1/OCV2OV6QkGmY6/gUibXyyUnsd9QVR+x8SfcMwm6DXJQk6HA24pXYODT9IyhTGNiv+
yOWesutYDliMF0r9rI3kYqcFirMn3cKd/WPIJMLZvl432kAdvlUcm1cugJxw8zuWHBjo15UL1dSP
CLmFpuVbvnbNTeLWXfDVI7XacMTWNC0eBuL7ne0kl9f+TaPoNyqCgo29aMnXc860wh1yQ5Qm+xbG
44kKNobaTKBRZKE/r+slgmc90akqUoIWrAh6+DR2N+tRKRjivFg8wwH2Zg6f7lJgBXXrf/KQoNZD
wha6UoHU4kkUe+AunIAHTFA0AHRrGoO38IOqDYLHhaAZ8afjpwJLuxQNuelR/d1sx6laDMYW3FLp
QRJ4ZS8hwNKWR20GUaASzLPO4MgG8SB5W3Sc5hS9Wqhbr9WFgzfyJkHNhB9xJYqErJsCC20Kxi0z
yQgRDnMQo99T+b9SGGHlVXge1t1z6/E0aburSAjiNgfXe6XHl40X97M+dnUWVHFEPqOvwmtvle4N
cCC/fcUX1bolrTgdFqmrMg/dWLXtgRc6SQZF0Ox22ODqaQnEIHQBmbIuw/RVQMsnI77FkL1paojb
W0YeX6Dw1673HMMM2VQvQWXeXpGsO0uw3fgRXUhRUEgENKAuXF2z9W3R/l+1X6OekB2LfgxN90Zd
cSDs25POD0ySL8BRnSFbjVHyUo6N0ZYpUStWjrJ2sUZxhWYSm/nMw5/opWTvdYRo0ndYtlGf05qx
wd+NmEUZWRxHOMO1RnVQHZvLep8Co1uDT1N7QylP42Y6MtDnDVzyyd9W0h1JWut6LghC7jzqIu2a
JeLNfdCy/e1ckj7oAIcUJT5dRCut2sqm/lL1TEcn5wepICJZVEsrwvIkxJEYZ/i+0dxbMO7RNEtI
iCUJ7qGKg+ez3xE2K3ev52VIouNRB1enPxQh5GwFziDRM3fSPgsy6zvmHl+2xsirosNz3PMHrFKM
d6NyMNZzjEYWjZrf9X1TGlz0CQJNnQiH/4ZKADw8HCkKZ+J3SCujkZd8Hqj7tiMMu4Xsqm43SpPc
yxXQbqnjPpJImyyVUmijVxzoiWoRF0fhzVKCa9Or+f7k0CHb7krNO/jN2ynLQlkbhFGDVcWitc5E
esXmi0kprLhgpnARldEnUc1nj/FxifdoFaTHzBoK5JvrhHnT+94eeo6y3beQ9Gr+UBrDj2kB7lYI
TH6cK3SSSJ/5lqD3SnH4smdcSb74mMndjn4mX+ByZrBNbJC1TbXrPF7fLQuaj0BiTe4bMhPatiiQ
KNWvSa7dQn7hjJQnVtm5+lTIqHcYCcadvYXKM2bJXwiEDlLxQMZDqXjGAgO4f/twvUQ7PjAnOeg8
9h7Y3LOvMYCkTrq+8CVG94uu5Gazilqzjl5MxY+Fj/UIiJzrqCIBB6rNbrrSDGOfDNwkkLzlPGMu
HaPz1qqElgJcdaqFgGtTPtrMUGrJM3ty0H9Uz4XAeWyvzPJR9Q6KUsMsPyrd9Dze5/aVEB3PDmtO
e04ueJLTZpOusSWVhvyi/U2sFOLyRg9RJEQ6V1VIl/5YVsmNBh9BMoWXqe1+v8/2iAQgzxDcF/I8
qtq21HqpcowS4whS3jK0m+8esun4Ag/t5VLs4YN8o2iJ94TO1VzpzHRAJfCmGULnMQ+jGxrW4bJ1
dbt4Z7H7MYX0xMqrM5ody6uxiwSkbFxf729GPX3sADSIU4yYwsEl/duJ3Mu0MnubkeMmNOdEM/aK
xE7R5a8tkn+AsyS4esQJwMjRJJld5CSVufmbu0S1M+fB7AxEU0sNu4ohI5M4RfUmQ6zA3paXf804
4+BRmPilEUhEeZPQ+LA5DwnK6BCPNWrIREvq6F/NcFfepPrUHsx3CYmQqtsoVV9is/bLyplwwIUg
xmMRijEi+LhD3hTVMLYoYIrBeNeVXylx1xAYrqGePAep/6hQ/dEfiDO6y3BA1RbQZLTaG/EJkTrC
DNGKedC6E1C02WPg3OWmqONg+tVK8O/nQZLGyMHxGwSFXww+kYwV9V6DqZpSP3O1yLHE5B+WWKNl
N/+zHYtApp22D8Bjinjx8p04gPor8ElPzMZSeENuEwZ/bnSpbhtuYSx81oomtRdgrptpTiwydPgX
R5/n0j/sg0GdWCE7qws+S59OR1piqTrJ3UNuhUZSbetZ2vl5TvvrAGVYmTQVb0ReHMx3IVcxxmUr
2gpn9TtsIycqnEdYv4BRFBQsigfGC4affsK+UW0ec6lvBuR5v5h6dzADCaKhffGUSg8Jv56IZ25q
jmm7PK61lea5m/yrIK9P6tHUeEvosaYlDXkVzgYvxlqMqvzUu8zOQxdoaJzTwxdK7pf+3JoeT8On
VdkQ1jXh6lkik7zHEZHUDeeYaiyV8CqMbQZyrhc9hBJevRbzze1omKhd1k6gFGBFpJE6n1Ir/Z7I
I8x8pmvchqxNniUw7R7zLM9ScK7V9sPebPG61gTOkvrhVWKcWQi7rSW8w8svqtz7s/tbNMTzsKa2
2/NVLuAHdKMWVHucvRegTD5kJv371CoK9fmQ2/nfVTVHF5hRfBbxMEgXG3r23KxSuae08o/WaoA9
3XR55F1XrFqrwRr2bm3bFih/pYPCWzj5J4eq+dVHSqTNh1a1OE52D3xEk1ww92pfteL0UINPr1XY
RUdhtr3u7hmp/XPNzhGebu8rPKZbvzwDIWad1/Lf90tcNIeqfBXQrIH9fFdJlGHXADebHEstsB/6
ViaBWg1PZfiT7UtmObHq4IPf8E2j8NG66SG/tb1/WLzh8dK2dUBSGAK7WQyQkpMqz+Cib5tgSDcM
6JQO6fZVdzGDuOWAeolqbf1RU0Bhm/3zIMrIj1IoyIXJhBNeNwkLw8iOWuK5NRhnOtete4j71RSf
rCtl40djpKTFaP6RY/AFsdPnLDX3zlgCvJv1Epvxvm2GOjzRtCA8R05Oju901jPcbL8KX3juI7NV
qgHjOFsQq/wAMa9zM+XyU3bOvWnDJN3P01z1SDMTdF5WISGYMWKsIZovjZ+wLvK4yt3w98xE5Srx
ZHgNKP1ZwrBfjsi5TWMiYgYlhgLT3RHDDcSNVMgS1bLxNjnJqJOl0JnDCJK9qeB2vaXEwJxJ5gKL
ZAcM1J3lPLMQmi5BRHmB+ALoYRlPH/wuFsO4HjsNUT+A59p97pbToyBmwkyX+0eMvOoOI9nQl/BT
tK28usDlC/wMSLsZKE7HrsgQApfL1RwMIaYZtt1Bf+ESUp/JxV6QWpi7kALTWpfiVoFm8qxT5pZb
0ISPhVI2MVMb0a+XC/BgJsj6T2f3Tho+8TJS3zerh2oFvXA8W0C+L9jPrX/pMuQBiLG3SXWM5KZM
WorADzQaLYkem/vxi03B1Q4yuosSQ5wnGM+fRHtNBxsOOv3SnHG2/1HdfmruM2L2ZyoyWC2PyZDH
eUCSLaffvUvok1dGGKNjcIM0KFaLNRTzMuIScdfdYpnfZcbRh2BxIbqySNpgwiHL/mhxGfUbGLsh
mEyXaHFK+5j0USLy6kFEZF5KDX1I4obNO4W60DgJ7iJ63gnIzCg20yDYKbwGejBYb9Ngt6G9odNi
qKCVssBmocs5pjqFC1gZ5p+ns+c7OpKc+vJUbjDmrYSqxuTwP1Q3skZrvyinXqzO3QWSl7+nmEbQ
3jG5bOYlPH/1FHruMpgoXfYEe6PgS4fdkw/Ni/xKKobLuIjNFHq2nz7sUSADpznf8JfAsHoECenJ
+JlzaKIzOsioE3g2IimC+sMIxTrjmUFVLkWYhcLEhVTC7B/BkpW1CRcVozxSt8Td5nWDh1r55vIy
JREyjhV4YwNVpYnfSiTQAk059dVv6ePiDff7TSejghUGPDIfTvTahGP82ABhQnvqpC4L+3XBfbgp
XG2ffpyxfHvthYjoSUGl9P3XSwwTQ6xcxpsqwAOJGQ6hcD+hQBPz5ybQhN390Lsig0UWquIKaq3X
4LI5GEHVrKtKlpCE+3r0PzEhrtWyJcWlBAduuYcoeR+Bhc3q+lZR948HVFrnA8Lj01ixYGKtyrsn
Kd9sT2xUSwpzRBL6399UDv/SueJUq0XES+FzwkyDkNUgCLJFSaLHRkPqHrEAhB5lHCrxYf2TXind
DOzKVm3wZlGfJvk+ZDNNRi7rgt+UCzLyGhucXZJBTHLjQan/EkrIsQv3Twcg6VX0dZeejqwXccQ/
3KI4SyhUDy15Dv7kAFL+z9nuhjNbEaEXK58S4hI2wmlGbGbtKLzIew5Q8ENtP21sMJ6ieE2uhUdP
88/03rE305SrF1v05is7/7MzWQXuEmUGmxVX2aGz70rSN9iAPDzYSytQDaUdxzujGyw+CDbVu6G/
upEElQ9I6zGg514NqHov4yKpy8n8+JNxX9u4QALxeDs5yCkz8gWVchHJM2TUWNxPJNebaPBGCaet
8ie1jiuKdxcZ5xO7ZGbYWTBScp4wdL8qco29UEWq3YphtaXadU7w65rIejIIvhpABDbvqeoM+x7M
5ICMapGaOXO9FoZbwgSILJUoND3s0KyfwWpe8K1vHUWdXRtZ0lorGSWfWNS3/o6o9hv1wpiy1aep
b6hXMyT9aw0k8lgTJP4mPBEbmEwjil7Qr09imsW24jojyuHoeIoxeIuVyCfgCLkFSzrYwBx63DJS
XaJw6TJ+dbFhqUNVlKxKphb23xUJudQotaK8l1V00s+DRNiP/SbTpAs7Pd/8QBvNKiR4WWNIkkPs
p7u6Fkt2QR26E/fZOglLurrauhv1N4/2fv5c0SN+Cqpn6LY2LKCUDRZz/v4sD8OfzjBF2ito2FS/
kV9JTB2KBsx1uKFyx6S3PSFArfDVe/mYwvWB9rxndfBVnUIdaXIrnExf/Zqgre53qtAc70jb1QJ8
oSQEhjSLug/5xhQSHaG8kPWzA72M8BhLfaSgboCcq6NMgYwFFZLNFrQ3bfgknT0dTLBpwz4ZYAnJ
r1+GjBAqrJkqt6XcUon7bGO4KQOlI7M1KAbkBq3RbJ5O48xLlQ+L+khWHlDWGkKGojTga4Nun/t5
nD+uz7pMzuBSNU8Y3gdIW6U0pUpHWWL1xvUq7Yml8VYuWw3WngiHqnU/uT0GIqgHz+Xn56famNv2
/PJ+P72Ay6r0l+JqvUa93Rw97/Z4bF7QQ9ntVPsBKJhjFp5HeAgRf0iO7RvJQw/O951p3zPjrjXD
+CXbNMfWI7naYnIuw7h9ta/9zDh9gtLt5GldRgMhkurjUWl2t73QszRK/tDrQaYX4t0iXahfYVT8
jGoOZQnNfAl45mGdtJc2FGHUMlCqFgEz7w83hU+C3JwotFT+dHt6GrXxIIKxSL9xiAjFP2Bk8qDn
iuY8Ig6yFHoQmSalwTkTX3H5yLApfaFF0IEGjYONmpNCpBNlgES4g3v5dBf/Nqzp7nIyEGbbtQvT
7baQkZPAy4d92saKZUcsZxA7R5ahYwRBd1oLeGtZo5sdSFokuYg/9bY4kjsRcP0Sifr8x//LaFSm
NCHIkJ1tbg/yRsIDL51TVHTqi9wVxnqvOGnS5WLk5oiVZDzUGhFhxoPmx2kwnCUWY2L7mOGb4x3Q
uhNvlfGI9EBV26If6xOkODBPVUPyOniv+TYBo4wXD/U1k3tsNZHX89boOggBPIxh/ECSdb+zb6KD
zpMfe/wsQ66kFJGCBsh1l9Zdm1hkv3Ka+6WMxZ1B5m5OhpsPondPkiJgctsBYPk1Vso7gmM+y/ng
DaxTFZfAjL/MR2OFyaUkcnV+tF71xYNcxKQDS+TdXxCYibCw0EmEt+aaDOZPOwjCABQjVREYKzd+
3bjwXu0uc2Ek92yqlRa87NwsfQk2UIj9vBh+7a1OW4ooA7Ju8+v3jhO4rdyS9s+bQpEVJOcEm6U9
qIzC+9UF53L8DGSPmgJ9vkbTZRsrq4iTqVcG/XC76yZI1kjW1h8nw8xXKW4Co/qEsJmRQIvbEPbn
+Qv4lBCWNCBm67iiZfvV3Sd3Q2zT9nDOddjtlyceKdgRFGKYUeHStvxwixCbNAp0/vdoMR3xBwDy
RK6lqknMQWNzqo9fwSyD3LLA+roxlMQS51eU2HKBtXlxAXZj65Vc2XtE7Q9CmJ/SIuyQJMtP75io
/e2Ly0ItIvz3jMkvyH7sU8Zm67J4KwQNLv0oa7cJ6D3QMeKsp6Neo5m41EeSBHB84gmWe8Cb6oiJ
Mpk57EeEHKewnFzBr1CoaR2Cyvsv2QSxN6tMJiEdVXH/rmE/JcmOTeF1kuzkkTJy1RqsmYlKWDPY
9HPPse3kw7MLUN951tJD4Towoy+P3Hia+9zaw6yJ7NlNVhr85G2vvgDpNch+pD6gmW1niHCjbPXn
TZbVfFuNg5OI8jk/VpFk6klBUlO7PtRVQWS1OMC5Xo3Drlali5cRuCAbhm8xO/QDHZQw4/95O5VA
HoIcjql8fwGx2So9Ltn69q9T2RqAV8kYt577GAYQDOY9thnvU+7sX5XPJnFPRziRYc4i0IfhjU8v
RUViHH9atB4vnH4m9KJgU3MlyiYCfJ1ZatZnzO2YEVaIDpnHMcx+qS4Y6H08teTvC90a2TGPvRKJ
ohXEyZZtmV1euZKFSME4TG2lhPBpso/1h+kja15iqFzg92MqwsPmF482XxuV96+ve1ai1xYbZ3ZY
OaDYd8RCASPJwc3llJehXhKXyoc0D7Cyy6OZlMuO/F/H933m+uufdHiiWCRMeGDI3v+HzkDxHuqg
dbS0TyjkmE3SQoIfcSW2MVKSgvRcCbFzLKW4DvDGuQHB1RXq+NIST5fijM0B+6HLYLiqqEZyqRgW
sabwYHqPOCjmGcHj4D+7SF0Gb46bx3b5prGmB6PeQgAPfO67RuoZsYUGfXMOj3zE7XqU8hosgPYw
s0hvT5HnSyKc0Iccss5LoEK12BxbJ8M4OpjQCeJatNqtBMee2ccBh6cEyztnk9s/bKzV6plOoEXi
763Oc5aQia4Np7uz038y/QzSl46lVSWV4yx9jU3IWkmkg6z3d6qyK6tQqzzlT52aDTUcAitk84cu
X+jqP9ulZeJbR9NT2hQRQB1vM69hW7lcF4xybbI9lKcLrWyp2ntlxbPffuAtWJLc7dPLM+RBRmr/
8TyvbKXq++zbXV7KqrYoVkfAg19c3b0c25hO8S2nKT3tJp9uEuUHCZ9NrpMGuu/FnaIARyLQLZ5D
ikoPE1EgI5sUS4IbusZWSzkphHQGWy1a2EmCYlP82S1MJpLIH39/s56UV8rwwCgkI8yvVr1lEQ5U
OGyOwBURv8qHeya2ZBwKnS2pjh0j6JaU5UpOospWfJoAYB/tNOFJ8iuMTnbnrls1Lb6VWHl9j3Xv
YJ0Jk+VZ2g0El/b4d0eOqw0DlcDn75QvoSlNZ+9sO20hrYjFHqO+pk41CT1xn9SmHxV7n3M6S6zx
fbMeeViaKghYApw1X7XaknYtVmBr7R2l+U2zY3meDQ6fCt2MgS34pKJuUPoH2BIiid3iG4MD+cQI
esN5/O6OtRvyNe4uGnIw2286k1OPTE7MhkcOImbzjwAJ9GoVb2Jx3RbIhyRaowexBT4EW+9gLswM
/veCGLG+xeTsXdQaboge6y2/EFQMTv8fLeglmQ0Qds5WsV6EH73kYd9zfmwqaHw+oNAuwDaoYBm1
3Vw/EyS9IENpiNJ6Y0UCSzmPQlIO4ANxYD5QdSgpFwzsoHL0UaMARXSkFsFrG7MkDLNzTP+c4wl+
X9DA0sF83YFY2Hy3WNcEv2ulJkXG6POQveuxzwC+sZ4ddPZ4iclZk7GnPy2Bkze8zml0ZKNyDPi9
uDiewkpHCuOy2aklyn26CkuGPJrlAEyWDiERIvyZ+QVMQqEvkwgC77Vo+zVOa6ncf638ihfpLcts
MlrtWpCutAsyVpvEDUwfCu0i0r02qTJPOuc6sz4e4Xfwy6Yc0y3m8hD2tXS5iDc0C7k2vBifesFP
ypi6XtNWJ/WX5oHIhW1rfbrOfVqVKCIDWmSFA1z49PeQHEHrQxThY1XKlOI1k/kB2rKjZ8rsKIfW
ldykljJqDI0G5mMP+dNsd99pTlTgGhFOWc1L2aX/xrPcKzrLYwF2itMXv23xVenTa25Dir/DDUNa
8LzIWcmBPcApBJUXZrRPuz44NC5xmtRZ00qOhr1hCtuOYWczSqLc6Bsa3mVOwizkQ8FBsx3+zEEZ
+KtvSADr4cWYvQ4544YQlTVctAhvB8ulZtpdZQshBAP4kZhWZmVj2wkefv/A/hYm4mzfOI6LFOq8
qFx87DUX0CiyOmgNNBMPNHTb7SrRS+7FKQZl9jTHKPLDNvoxkK+SCSEQ3kWp4gYcWTkJW6KuF8Fj
0qLJRfSQ1VdWrsZ1raPd639ZeGEscJ4RSJ0tRdyyekUfr973OhSaztWDVwSahgj70KF2b4oBm/mi
rWm3CM5sqIFFPYrpZUi5Xaw3LPoS2rvJ81nDPqMTdLGDdV7gbPQNPpDbxRhojX16IWpJNNVwi4TT
g2/cCkA8n571ydC9Yv5bkPLxvuMTzmBgY8vvLZqY3VgbvBFZH5uogalrM2lSB55bGi2OAZ0TDebj
ItYT24UoTdMMhwbmc6veL2QeBBL+7kKk44lc72lClmT1I3Huc8C64Cy2IuszbtbOjQTkcu7yWKJ+
108Q0VMa+/dT9QhBy04GtHz4/cwNT9Sc3RV/kJ0GPAaBTEEJFOHCy1vDd9mTbUntea9tj2/WZl2v
Zo6b4jeYz5UnfO51kcDGSgtVzPZkxzoybHmmJMxn2GqX07HMz2zx0YGUekwkF7A7iQ/f25jwk8Qq
S5FA/+sXzLlpBPtbhf5hIXAoLAwlujJmdvgi0MFq46NNa7dfkE7JHzBQ9ki4rBtiPWXegAfHvuqv
1hvpbKNyFbMxeIGYV4kUf0c+tjveLigzvuFLwNOs3Aw16+1t6hhW051gmAc9WRAARltonM0BZqOu
pVJVfFkr8lRU3zgn/oQYVUOpNf1nnuubOhYvj8iJzgYfwppdFc+tVsf0IBPGIjwCo4IINbvZfD1/
bl/hcH0+ozZlbSP0eQzINEZtlSf7ENEfaUNbKT+K6En1C1SdqQeZd/vsPL42bT2cHQamBPljUoST
ZTIKjWHGls6sUrKaWkSDV7mbL0mI8BThnn84RiCRXs6hxOFVBm+tmKfFwpMD20iIDTR8sEhE1rP4
ydnF5JzxftJuUVNsQvzFTDa5E3zf+UL5EKq7R82uht2KMeue4+m3PUwCK7szDvfwAR3eeZtYNBvq
m5JnVTsB+uosiAXWrBjO4Gz8WowlEx4APkhJozDOmNOzN4XquKsP61shNwXzSnTduyNgVoQE5oqJ
pqy9Y2RIRfDCUdOcDaVjmClPM5u+n3DHaTMsuFuQbviZ/dubQTSGfJAhi3n2bIICz5ZJ5aST/pHH
O5rmP96Tj2VSpXBYL7NFa4gZ2UHrWnC35LDGQ4RF4EzjLN4tz0lIoFMCPZCPXvVyH2sl7bhPw/f9
LiJ2d9xaWws5/EcPpw1/GHY/tIMvJvqOHjLM0C1TSuiCs7IR2ov8pty/wQYWsHtBp//je3P9WD0r
HFFSM2HEU302YmgkG/sSYwORRDKsqf4z0ncXkvkvvCiyA4SKJvB0Yjb9Fas/Cg7NQg4sGPfmPd6J
NPPRVT60ImyYLW6VSqX0cggVJwUWnIbRz0wPIQ98umFhDJJrsEB+BJO1YS8W6UOsgVVZcF15VezN
Vh32a9VEx/tNtPU0vxMjaGm7JJ1v5LPRSCSXtwWAhzBOClpvySJOdZH49IM7+P7WvCqaQbXJF1Pd
oS3UK00BY/3kMwJBRBk/aGH4yZfGoo2zUk4NWgfcRi2glWRzLCCx+eOhwcgJcKmNIDaNnxFlI2+S
GI9hncS7fMCo2+GayyMjRVbWtvdqIEMoGsG8rsDApX8nIBSA8aD4iiPkq/W7RhkdwpKhWi7kbTwo
Kh/bvGMOSjcWbHK5SPC2B0tUdFySNiB+8EMGsitPasCN2l8tBGleZIIqxWgTMxLgfRj+8LK/aLB1
ELQtEx0D4cv2BasBLJnJzgTHIjddmW+GZ56JQVfkvmkz61OT63blX6KZWf7eb1Zc1UjMCWOkCp/y
rM3YdZfjE5Kx/c0U4LlWRntsjulYwik1GEu40ujoABVigAz8pSapSxsK5wUHv1y/HW6wMhQHQX5D
nZ+Iz9+sZ+vued+IPR8NHPNgaoGgmSoHvHqvzKgZGm1dXL2pqVtqLA4wEUicRA99f5SveLFur4l9
NSJxJPDyDUAGMxTZU+8veK1/X7Jkc0EtS5vB5xmlCaBFyVa1uL6IErc/gtEhYNZxbunDXDqyfg0q
Xy8ucDN/XvBP1GyMEm1/4zO+g6fgCPuAFh+olQzGTNfgVfJt11qV8UrR+sD9mz0qJq3tElDbJvAT
KTi5zhhnc5lVxAJF7OHrtG5hyoQqQFujjqdhsVZyKcbaBrw29klss1/WVhBGibdQ8/jc0XDLlL+I
VWu+/UG2vhEEolkzpPlvgLqbf1UNxW1M6jg9X0cb6kt048ug9uP0KwP3fjmYero61NnwBQQrtirl
+QawL2g6U7QMGgbqclTu0LvRTO84OelHW9MhuYZskFHE3Uo1z3VKGG+U0Gpok+AveTUxTNm0a3e6
5PqyBqNA1JzEVae3oAHuUo7QxXeBUN00U32zL0SmrPkF+2NzcbM6Krn+b0HaYyY7bgQTsN+tIYQw
0zaNbBjy5lWS//PGwqcDhNCC/ea+2vEyVFsXJF8i1ae37gYkqBKd3nNW/chaD86SBmGYmnMg1NXC
9kIVYKqcZxjNURzfc18wXLpkPkZ5yD7P/HcwBrsJCc7NBluu56XJEjMTSF4QV2ApJrm1BK5Z3aGo
PEXhU1/Ohbdwxurqqx0xo0eXGDnw3OuAdOFu4pq5i6l0PJKKqWqJ9uL77gP8TdAAhCnd1exYdKof
LHjIka38BcbYKbokTVLFRwjwmYrOZREYnKSowM7IiBBZJ4sp1qKhdUI/hVbQQhWVoqt2ktwNBuHA
mFtCtbxmqNB9el7KUmIjT8ae/ZgOg8U3ERZ8G+323O7Zgiweqv+80vzQgDGJIOz5AxsvITxzcYGR
lxy0eV8P+M+efCQnRcIjdrCAadoKAvdXZQqujxBdkXu4jE4uKl56kCGHf9Jr44hE1x5Z9kqnWn5j
ER2GuwNy0hHec6YRzE4lA3YU0R77F26cENBinmiq8/yElZNcWtwurIv+ewl3hHrrK5oV5YWUO+gu
KGDxdHioSUzJfK8GJuo9KT2P6OLRi9kZ4LKOuKrWOHqidcbLTi354VWXt0QNJYbUCTb1oJkcwKQx
cQ+IxndMJgNUgyr1XHBpkBSGuhk7JpmjCwnfSFi59sI3DXtOkBRkaBIXZgtU2DH4qufoUuOAJ4Kp
411CO/ETdZbua38ABeg8f97bKfn+lAxMfTxLu5QsSeVvCbeh3VTmN1ENRtwCZvg1I0Nv3Q8ElUD4
PY0GN/DdTpfiYRha8vf2U6ysZtZjEuVrH1NL0ZqyJmEfpLYU6+2Q5hrz2TJ6BjqPkgzm54UqIxsO
FcAmiUqnfwx2TfcASxr5czP0LZvTbHaJFd+qJ0cEo2LSdlRkojA65Zv7HAQpv58MVK0W4EOJFoTo
UVR8km6NACQ2QK6eWI4HLADzcZuiDs+JSXSxe9rvDjdNOBHKyK+aaW22CEqo4SEkl49uwdjGfAev
5jDnvfelyzW4iYLwVOIuEIyEhiSfdxr9qukblEdZCBcy2Zk9LSmp+tvnUKYj/XMIbFXHz+nIt9pq
6nYemDvzGKXyvBCzPtbTCGpg1b9dWBw5FC6hd/kL4Rc23Mtk/6yggGz39/7drF9AeyDqMzc7/bKv
VYTvLJXPTDbiiV4/zS0eJS1/o/x+KjewOt0pFbjM7bWe57oVqANuFYX4w8Dh9x/n4Zy2wJx7VjI4
j6bHMcCKzkSnohR3nFHURjVGTZMIz9WLVYxQTP5ePFsydzaegbuEyHcQvZmAWpAURM3y/zcXrc51
80X/fgVNdEduYi1/6aDCs0UJcxEsADJFfey2XLRDOIAiV2BYexAv4mNUfAMd74Hm19ZfNd7j+3vo
GL4ds3UrMRRrJI2/TCfHUs49rIVHfWkqyJTU+pcETjQBCXvG+w2BT+JGgEAZbCj100TZp+iNhZS8
tRDSq2DEJNYm+SJ7FC8il4RnRnhbuXdjHfiU7MGHPmXxX5ouM+VLC1GY5wBrqguOjDhPU3Qa8dN9
3V6pBLn5pyVMBQrs/10KCEU2WenowzxHveS+RBFmW9IzQ5JzsZMNq5hMJEH3GztjVCp4QK2qp6C2
IPtaxlRAiu66zv7gvo4/ahiWmuqteAjE+toDxad/HKICUnjWL0qigCcOiHCDqaZv7KII6OiyVYs7
9YQE29dpVi7Tu7QLzwNCSt+bQB43OyYfXixpm5Ycj1oHN07lRoGV8zIoH1+yu0MEs7xpilUtCDIG
wQNXgmX/TfXsudxCEkqTMC4x2Gj3l4CdJRxiuCu5fwnq2mwGblI75P/GmL4rdg+4AcvEG6F6IiGa
L4TAFGrakopq/iZczPcAfiKShdFWo95U/RfgtDUVL0Yc0xmO/Nl1iO80wY3NXKqqvxkiK4ddpmT1
qaC7qy8457NzEHRDtYXQ2yc52CiEf9L8cai+PyKZGAlcuXNS4FnbmeWKGKlzAy8E0aumtl9V2II1
PTgxL0D4e1g6YloPaduqhQdcXiGGaYBCPes72Ug4uW2zMJY31T3MFjjUfnDpzYFxF6JP/R9GHOYm
pOPbuu14ykoCeJdrLz8dkmUt/rJWVlc8uPeDphLaPNDcFUnGxssIfOgLHvwrGdcVf1FYweL1SnJp
aE5EEEJEkoxkSK3mO/u7AnwycSAllGFTD9H/czkPvgjyprZm/6ieEnAIIdn+TRRPXuOExIUyQ2r0
KP9iY9PKd5DilcbReerct9uLoCrfM7VMXtCrrLofRTCMYnDUgfDEdoqQJwntZrlO4XmjkuYF/Z+0
khlLxM6psqDS3vyJMHVq3z/ri2ba7kSSAAuuSJDCAMTaI4SZY4W+J5Qyu7qtKn/r3tTrXwd1SOsY
X249oy8J0stgq8eCmPphU49D8Ci68xGfIsRf+7DZRYQLjnEtxpliQeLWxTfysArFgjFNFYcAU5t8
pPFmkXbmyFiYyRC8m/67VgQ/MPs1rp4JpoiKSYlTqismp7Kmnjer33g9EV85Tczi2/dhJo3SUYTo
rm0JLax+DX7mcUiNv4t6WN5hGnXildAnENt0slswXfv5NvQCBjAo23mEjxPALH2aRIjCKQsGAV81
JxZdpOWCZDatP4vOGnQRMREqrTV7JMNCD6Zu5zg36r087idUmT9kx7nS22xEbMDVQBT9fLQIWZjl
JCfR+V3rIMoHDLLSOoSviNfKWcRqiYVpdIuvQkDvomLB7Mu1WEi5QEvQ4kREZlzTjxjgMMuZfwW4
bn878pB+x4NZCDQdvCnMxzvDXQhP4Rl8kTf24Ud6forzdc7R51I1ov1VuBBa3EQlb4LoKKAqmP8X
HED1cb8cZ1NMO2tDGrRmRmZ0uYLxXYYlT6WCx41lDqNZpbiXtHK6hrZ7/9X0Ou3qVOxwjAtScbfV
ePTCppEleWTSMbUmPn5Y0GAtMMQE7MSYY3rHCT5SdbIu3InVfCOaZ/p3VcmOGVNSykIU5HTv3pbY
8Nt0B3AZ06MnT3Oh2Jlv+chQaOvb7nVbG+99kIeut8tfQxnbMxyr7hhE3G0hHEcgWyAwDsOn+p+d
/a3G9lUIr/WEUvTUNI4KdoIQ1KPiC6AF8IJlFD6DPBuLdMVyqbHKvwtNgcLlmQkEOFzYQBxXPkRQ
UwB/EN8fiKwXe+TUjLGUSqezFsReTfOuqAOLiJJ64QOHUM9tIbt0BI+0Qo12Z2y/K+NFlL3rQP0A
/k7CEfbCpzWbLwW/2AEGE5NFLqB2UXTSQXHE7OU3jFk8R+BL9vQP9k+PKeQR9n+pTEMUsilWqLnT
pLCnYcOWP7wq4gbbGRonkWJPI78Y4YvtRtUSmrmjsij3OY6Qu8xpU0HBeyTRASHXzYe0aUZ/gzOv
j8Oxv86wksF3OSvlVq0J2tzvFJIH9zQeMol7eZrT/ASNgMg3AHXfs65SCp+D1bojAm6mh2g0PXSb
EYuyW8nSe+Ma/eRwIHFqoKusAlqfMPQwy4yN47/jSIxkkryQu05OCnKBZMyVJMCoaVKA5LX1g6DB
mQ1PbeHlj/nhD2mosRCd0gk/c5bRCOvAm9WQh0owsbQ93/L7JOg1nrmNeD38ZUxxh+o9OscAiEAY
7w8Dco/L+Rp6QTw6Twy337SsWSY4UMeCz3cGvfOuaTvbu8DKfNJUGYmXj0LmNRrDnk9Zb87uv+ZY
+aAbkjdDDKdIda7w48vJsZu2NyUCfHK/ngOgxqs2zB2HLCKFE9ngA17fmbG/8mjz74CeREzwxgj4
u1pYPoCqI20laXMYfc8JQ+LI7D4kGOSrGTd4YeZdGpLdefQ7E9AhQIB3GNUWWWgFvHmV3NzIx/8I
Vp4dBeSagwvH7XSPnr6fOrZQTo9tsyZIdbzNvVSB6rKjs/DhI3bjJwAk9fjBoDGI6hi2glM+89Kh
Ajx6CNT3JFsg/X22o23TbaeJZRs1Xp6RuzmXinZYiLdmBuxqqs+WeOO3FX63VxK+qcgJdwhJuiFt
9/B6qy2EIYYRd49BQ4HzcNJpZnNEWWHbxFITneTdLTcsJANKNFH0lcH6ol/Xfa42B5GRx4U3qJQY
e8pYpek/CdTwUtleCKepWAuCeAWx6rqI4ccUigm4Efy8kGB5UX/FE8CO3Yb7dakfquSgmCQDCEfG
0MFkKADyeWL+jYRmeTwIRspcq33qvXLsNM9NuOnDzoMkfRfVCOpSc6Gn7u/MPsBu85lT6+xbQC3o
1RO9GyI4DXuIhyDYS0ueOPGyiYnMZIs0sb5OwIvtmu4vVKUAPpCnsdlE3agbFu0H1AV5S32UciL2
RGJgo4kTLtTOUOsw3P+tneHlHnMa9i5ax8IpzfwCjsClu4z76WX4phYZlhIFgyGdFBcNNfYSPdqa
U7zY8fCyJM0SHpxiC7/vViAfBFmBVqB/zlAFKp0iQhvWBn941K6fI8KKOeL3/DlyWM6GkqOa9gID
EwgSGolM4YgUo5EYenAWT8ByJ60AlH5fZloR9wyKBC6Fh8kFja7kd7DFc7QkyIACCS+vFfSzQBN+
ixjOXYrsJWEuQ23OakwFRCTVJUmDrLlKF+WbG+/DjosjIG8aXpwn2KH02LNucwPJ0aKFIM4aqp7H
CQcfrAi/0ZV1iYyvZRzjyOMn3cozvdn999juTInXcRTtGU154pMWtSUBlWdCWuoIGNVvx1RqihD8
ckzsTQv5i1x8Z+gbNZRqvNj7wTdcSH4Zs4cCOqK51cLzQk4+TRJsw43CpKwL/e56t/glVPWtOPnM
2SawDU7XhIHPe2GqUd/s3BWufj/aaDoGJJYJN6ipgoS9j4MAEc3WVY4Plz+8tixyEcLIqguAdnFQ
NhjmqduTqPBzmuOcHW+7AWxVAOa4mCwIm/7CNHpyrwbAVIssfNn0doNMbvVvajXAmpjaQ6oCV8jB
tDskGpaV7Tlh/6BrNtranMVam0MBLRrr2GyQLYAIVuskDs5byKAMD4pkb9fIuMV+z39kGBwlI2ol
+TBdcqgNLZ4h41GrabzJGtZLDBpNQjsZfo/522fVUpr1jcXTIRFgYxViwX4YOm24x05lYaayJtaO
lIPeNvb5x8Pjq9VwmKPJTD2epleftGOnsT85BYLsHfLzMKV/Tw5LrLS4NZASgUXNiaTmr3w+pHtm
jm17hI3sUi5YKYuBqh01Rvb5mKWcsPEkYxk6umxk6cqMp2woy7QqDputraogb7yooQKPKPUoRilO
9MSeT7BiQYjk6k5j/+j/RlRl7WHGMi+TUz2dbpV/vdlbLsu/R2/kez0oZ8ew3BSlDGj5u+Zkw+If
/s0gTl9JDmE7VMjs73s3GGAZtX0ZBD1JLTKJOslCF0ALDnOEe/T66jy1OzPJKAH/iyNtCFNouq6o
LI7TkvZKk8LpI4Oh2BH5EKw8U8AOu7sE8w2mWjefXiF0jE5awQXF9GNN7otMZng9cybuwTaSc292
pN4D6fGMAmyzPzmLWJjsZj8buMlG4wr7SV6cioJLFR0E1dPyPVFBggzY684J/5MKGqR1byAgDhew
f5QiiSXH6hgl7krq2JN61HmcPP3elS7Kn/+Y1qcSst+EYTcv3Ff/0M/nHlDXcKCLoFaff956Jnq0
Wz899R+1HGi0FuP/UzqZComFMcrHP89aqDpXSuWnAHy3hZNakMZDmsfNoQ83Hxi3SB9RgIk1IcNJ
+0w8g4udPOgTIAcqasLcRq7DqP6aFB8eL15rAvnUcfr2a0tDyS1aencks42XmnRRsDK5RTFnkquf
XMxbmOdUOGRdQIzv0BKg9pruP0ulNaqqa4NaKxIEejZinwR3nM8IBkA5wWRWX47inP+mO/vxZzhc
5VpcHm6J8qdDwe6be41HJ9FbxKNvkiZBxH1xS2s738szcVI+S1blNR5Yc27qGgIyk3cQziiiWS10
fhQ6JwjuUAXUcwpnHiq7dPsxMnMHB+inw//h7T0Os4PLe9jB13u8NmUHZjiTGVZmCjn+Cr9EBZ2N
OSh8c547kn2RfR/XAnlUlBS1UmvnDicf4hnR51gBpYsSD0+eN222CEvhQC3KnGO+GFTiu1xtqDAh
Im2Ga9K1To0+VSQord9ZsVxyQTbD+Q5/nUekdbGODCuWaTPN3BZYga95DXhdmsMPE6cdYHFiDqu5
vvaau1gEb/ZcPP5U/wnHrp41Svk8dwaPw9IDCgBcAy79tPJna3vNsAJ/vABP3CW+OqbhLtOdjgbM
7XimdIZc7HeWnMHhcScsajhmQvHvj0EQRe4ER4xcCF5lRxxnn2AVtdiiV1qkjrMRjcHJsJXPqof0
22L5rTGMikNL0At2Jz6yrx5UE3PWTuaAdAhlVSKVkh8O+YbLE8kb5zOEo6rSQc96gkjqMrk1eJiD
EK5eRTde0e6rj2gKGPX+1IYyXGipchmLP930XeFBgxuBAES0plKMofeWv14uflXVCs7l6htCAFt9
7pLY8qCKQ7GJ5xqIqTHEwrrrEtDYA6hDNIWOJhpmjprBDIha6rfrr1C//Bn3OATlqj9kFkv4n19T
dSAYsvRF0FHGdDC2DYTR7bCYV4qbo73TiJ01T9RyYFoJHwA7BSoVzl7x6nxn3yrDksCbwl1XkFzS
y7tW6+drGstqYcu17WcpUvD1nybMs4/hEWZG8rdcbmPeoaBLhRU/TqvHiSvdj6UKPXsi9yODe/z2
nFZb7Bmy3YsQ3Hcu7+Ub5LVprUDz41+c6ZksAm95jdyWSLw8vy+FRjUdOcnE3mkn8HApc79rbOpz
THL3NwZ1v07Y4LFCPT8+LbvgW7KtRQbM8cuag1GgM4VhgpukCA9nuz34mj2K9UdaZKkmgW1y9KHU
M+ijCsS18y9IIjuqWNI2naKtAbPyNz62JLSajNbfv82IamfVjQt3PI+wV3o/bC7+ZBEzp1d6gYuD
/L2RLdATeqXqK030PdAiE+ApoNnsepNWv01gRHCKfGJ3e3TMpmj56gH5RV9Niu75RMiuaWntYsAa
45GEYpygQGrzvRCne73Az+CZzYTsTc4V3NTR1Qi0sY9Y6DHYHESu3tYpiUBGPBAUyS8xoMt5kP8C
brCrO1J9oFG79XWtQS4bs5B8hkrPyU5xVW+EtrpblQyC/uq2IXimN9RCnH0XKAjkgLmZrmHNixGV
Ms2W0x9xo6FxXzvmPN45NUpgsMwkwCU3JcaXMFa5K0Cuueco1ZUbcKgRJWpmPfh0/FaIK70QhTYS
vQjvaKw4beo22mcIaValKbxvxdQEotzDuzH6fseGSn4CCoZ4oJEl8IIN6Aa1aRSctLS1LIAy2ZBz
pvIOmVVUykxgYiD4BePSgouL2YhBAwaYRgXee5RsTZQ/tIdX4gM/k2NPcvMlsr/Kz41Ui5pg7dmK
zeeG4kJAtB+NhA3+KZ9T/4tVs1jcNiubr8HxHSgDuN+vb+MBcoKqb54uf56XRUJXg+Ev4oh2J+lx
mW0DIDi97NJsrJX717AtRRjL24R9XHroDC1Z95zsmdKEvLVayrWO4LCmkvHP6qf1pXNnjZUpTbIv
8GrlI2J3szzQA4LEj61HAhMyzj0R6gVrmC/0x1KMpU5prITuXlSIGdSNd/A8GaxGgtDxmFoPqbO5
EfMoq90fzdZoj/ACZz/N8Pv3ftMQ023He8xTxvaZL6A0NRXNH5uiwQlacI9Rli7XSVEG9xfx1hIU
RtqFPxNhThzPPFKRkLJYV6y2tFm0cwrZ0WV//mDmDP0rJ3MaVl9ZmwM7mIMdDHVt4MQen/vvzoXX
r212yHls091DZs7X9u4XTNJU7JxaVRHenjp27NK3dTmtSn6wudgwKMWBl77XAsupv/1dwRtWYDQa
mmY7pLsCDNjfzxxLinKCREqT8KaOhyulPsFIA6iKOE470qqQbObKwsUrGkpcxrH1eMi5+buuhIBt
3OwK95+MEyrwndHniBtVxwW0f1rIb0SxtxTS6ENH1W5CbkrrLjvLY79BB41V/gzJU1K48yX+4/Dn
rifRkkUiZ8aAp4hzfW8FHp46YN4tN1CYbq9hn9zWcIG5qGKA/Wdw6XEl1uHpYZcalAG3HJgM2fHe
D6rajk9eLvtRX7M+4lk/BjdpC/zOjs1++uGURq36bu0CRxRvJMuqXO3tcL29gZk4SpkTG1mG1euW
YCt9dCy7Gd4j5by/iLbnevn8FGxhB9puPplhh0q10Q+z/SXaZGgwuh/J2zdOvD9u4fOMIBFy8k0O
qCuusc5RR37L5MxtVoA2kwgy8osu7JQSapdx4POLxOtZUFLktoacbsbqIplM35LwSXMYLfssNwzc
RraLrBzXGNO3wtoTZuqzGTBBa59F7Gs+UWK68+c9FaAJcKnAKLTgxN0cN6F3/+sRDV60xZHzYUvj
4FOKvpNw6nlhQAQM0CzvZl06rITUUgM6mNgR9O9GDlceJsVNnbvoOpWj/87f0Now1wV1jr7ktZlg
Px/eW4n/jjqaBCF7rrnOQRB6H5G1erkwvmnFWe+ERyKXS/ynEgpygkPDbYGrIFitpwarpggXOvN4
kjMFjcKaAAw8F/XhzabO/Y4qL52Jg8gSlnjGeHi6Az90aMjwQtXl9T6vJmqzPdM0saE1oSmZIimc
4WPiwamcGAQx9wiL+9sDGsciFVxlZRyL4FoCxtIRCauWzBA3s3teD7X7M7yy/PKFEp5X8GS/u1Op
J/kK2sCB6ybtevvpOEmOy7HVmurYAm8jW9sX4zoiPGszGJGxsx8/UX0ztv3b5/apgCtCJuj/j1X9
yWVZWoyTcs4Nfoxp6DD+jrqKENUfrAvliulwqDfxqcj4zsxEsrcY9heSohojPKaplEd0ooCvWQEW
Exx/x75VK1+M0lDaOznzhOr3iJGrgJcSyQiWp0Bb0IhrOLi1O5ghVFF4ejdW+239SXznaWYPK0qs
Y7TiLmZK0YwQhGkpwCDBBOKpilfMJMCePPiwulnv09uKT0/o4Jq7p7rRfJq00NNLb/Z/F+QcMSaN
AvSVmS/sXiXyWgilbZ6DnM0oqFFidSP/yeUWbY5Ele+KVJoYcJBtJFOja05roFnOa0D+AJ1zey25
4E3rZ7MH9FTxojfk1suhuNH8KzYNC8BvZ/frmh5vQhYsVDjn8o0zEN/hfiTTaKLXQIQ6YppLHAUt
ddjA/cEq1XcQJ7U1/1jOHZQbkVOnGwfeo+2QRgeVO7LLHked6h1m3agOkTvw1jLk29+F+HPGHJ46
6eODSCYc5gdfLGqHeUm/jvO/EfWgfVtTg0AxHugmMLh7iViFvl0mxi8WTzFUKfJGHmBCJVpGC87j
gMif3Mw8pBlSRkruoBnM/hHreGqPWdQrNEkM2+BzCQJ2M98sYjcw0/l6vtJhhNtRc9Kl2BjZPWQM
dYOV/LXdLO0FkrFEfbdXou6qGUzGM16oojoMEUb8tH+oeaq8aZsPhKMPL0x2O6VOKRFCsmj9qb1/
DebsYrBP8Upw0Udpa35LsQEa9Zqdg1Bijdow9VGjXZpTFZT25PGA7d8sJGubB9Q1Vyd+JgQsYp3g
5+EDCILzVy8bsWgk7dzczeSb4QasNIF3zSADC6oUwEIIThq2ZjKfYDul+DeQ/RXol08TzqAF9Cq/
9eOT+RzoC5JaMGK+iN1ackREdJG2YEFaIg3JL0LVtwIYyWqPFXeee8NAgHgFqTkZ8VTnio3TgVUx
n7TMDPuGR2t7sVwcSS+/q9xUQfduMXDOXUwjW8qvuucy2rp510HhK1TNL1aShRG1mhJjD343PiF+
XkrXPpkACDUrK1aE+u1TwWtjRNv7TazA93IuHWErbBGvUABBO+PJ9QD3Z4IPxEZ8vCjyasCMxlmV
5iP1BFwfBUgI0TBIYXUKRlT+RoLjRZha4M0kZrRaBRUqmEhTQzlk/9ezxACxlcfGSLM9HJ7h0Ake
VkTV1Z8yKpMgAcSBxypPzXt9zQ4B7E5c4lZAXBNOWdig9sC1kRRvMzJWI3SFY2xybGR3UAIGf6Ej
EQrASjvEVk0C81ShVzQ9Jqf+2ecLiuSHVoCIoNgQrIuUrjMuuibyoHP7B62ZGTIEkWaX5/FtPRpo
t6ZIlIaAyr+lwE4vyCxP33D0E0h3K7YFDpB8MNTkGA/mqPl2db3v7EgmRNMDOMPO4r7/tr1FCQcQ
YGU1eq4KM6aBx2XMblWIbpmzqIZSQrLbFDOB+lBpo7wxdkDF1O0gPaTdqrLTJ+AfqbcS+A4WIrKq
Uw+vnm4wq7fcFO6woNam4K2l8CZ2vVMgENJKT5e6q1ODj/EYiRafWzas2Mw0gkAicbFkoB9dd6pB
v4SyTA6niO+J6Mwuczz0HwQUNkJpu+auXmLNBcnxhbbKc/gSDa8WhsugHQxu9Qffw9CWGjXZ9rfX
/lwkIsNi4sJud79bVnb1E1x7rMjFSNmZoUfgcFeQUqR3ZwLedHLlJqXkroE98DUDzvQXXss0oceK
ifult4QWQBL5gNJ14zdh9MLa3EaHz4s00rZE3M5L0yl9JXoF6OG3SwY0I5T3e1Ve4i1kQdURFaVJ
EFluXnVyY0de2cH9KGZLAZS0ASBvu/Wndncl4Q66+7uyj0qXjp7258XucCnGO8UbdR1VUsBD9oy5
A/fVYNys1rF47ywVAyZWJdBo2hqvhTHRsWonXxKX+6Hy2oV5JedQeKhzRms6Ut0oLQvbIomIRcYa
dmGXH1MslKl6LzmcLrFB/7P/4oCp65iLznZpWeeYrbAp0AEkUm1aoFKBCuONS51JnsYRam/OUXNB
Cne62mpyqkPMNxZjmVbsvg29Tke2nVrrB31gXt3swVanGkIM+m204iiti1pOr9OijGxtQ9Oov0SR
EjPZLpKcnkCdQV4ZyLYN3p2wFyaXWESu9hxLDloMkg3Kc9M9W73H/clW/+uox6oV4t8id3U3BGxs
v+hGCESULN4IQiB7IR5oiJ8B4gnx0qZ1tEIr+7gJqCNW4V16x03ngKyx40FseNm2IdOhq00dHmaE
YuC8RnxT2T9FXX7e2vmE3An7OZhKTarr6KT2AMcWyuIRPYnji6mSPNP8gcx4gPJGloV+/ay3yZb7
VC780f5T+RD4G0Kof7LjrvGEryXAim4vlVHeSJd81Nl4JDprQhA2mrFzRYDDezeu7hHr5N7+//7F
YSvqPUNy7h7dNfm7shMoA7nNmMaVZP2gRiMQgwhXSiZdzCrFvrHQxsZJiT3OV9dPNZP32rry45WC
XBcV1Lug1i4MHEfYnPMmVYAAznrXVyrl/ABs+r/zIyGZv2codoA8YR2j54f4b62d7azYPz2xIL/A
DRHiz0Ap3rzmnDZjYMSPOzxjcaSeJ6VFcqR/DcehIMa5vs1cnOaYfMWejg/enwvGSABnV00OYaIG
DurA3Ich+q7bynLSMzwTQvjkzPMGaD59mt7nmbravr0mne7nIIgrpgCHIjF0h6rveLavk/ssHqL5
c+rxXA8GBHnCpdzja6KDVvrASW4rqIvQew+0i4ha2t05N7HAu4ZBTi2S6B5MR6WirlcfDNIVsuQM
yDHn7jEHMjrWg++8EJK5LLe4D+aju0f2GkoEMQUWpwLqyuy3PO2UY0EY2YH3IqXT8fhahj6BUBs1
LYFvHVhiVUGeh25dSCdl059eYXWqqDbb/zs+bErhZMWpmw5FR+CI31I+w+lbgq2xyvXWCdAI20gi
YtLWHDXYBI593rlCRHUsW96Sf3xETuYOvldwxpn4jMoMl6o84gGAb4oHQFygbFj3yKbdB5PjXfQh
vaZO+OXIH7b4ePA9E6r2amGnCiJEQ3qo2jcT2OLGFRYTRkzvf/FUM+M72g0lVSA9mhfhNTeM1BHY
lEECSYw2G/ULytGxWCGgBR7iRxQvELpn4Bfl6WetGg76/hAAOoU1Jn2RuFBuG75T/dDQ/QPjuuaP
bR5BD/2tNmuJjHg2gb6iEbBKKwkKlRTfNa7pwYyJ4LZlKgiEuDGaQ4CpUkylWCcucAkSxYeVgOfd
K5/fiD1AWxDl4lWcJx/2dqUL7FVzA+CllSIsNEVC/w/l1ZDnvlOdWgZ52nf+dKPRyRIZcChTt/2/
Tm+7cpWBkvxHTP3FnzQKNyK/ExEGxtPQAEijdwdj5c8WcyLaai0CogaALhgVDFG4XiBMr1dd91w8
il3KAcqNcvcxUJI9j2JvTL9Cws6cYzVsUg+Jgv9pKQptqF/s9mUhrP4noWAP4cvIKhrGyBJ1rVYQ
WMhVl8p4wG0QQPvyymaZdOU9E3clMudC+KN5941G3c4BW85y6ih/A2GVzAkngV0lOw4rr2ug27ps
7i/DncPKljZs6o5oZDYLnickMCWG36l3mdOelKoYtzi2RbfY2kF14E72PDSpS5BnBRJZMtERVbGC
Z0FReQa2+rdtHNLehey5suq3xnFqdCBht9owKHDajcvkAVU4BxXU+A88NjDZsKLB0Ezwlpj8jmoD
Xw3ptqJPkdTQRw831g5lJzMZb40G2kYyEjhiJGshLQOKAQFvZ1WMZ+iUxgoJ0SzzwkyBSQAuOpv7
PTedTlkpBwB9F+EmLrGayJnJ3FADlbXvnJYewmK5O4zAOzcYIFlAEMztWC6xv7lhomQis79qDLME
KSoMH3/srke5oaj3KHS0+6cnZp3tbRlM5PsmjbmHF3/SWGlYkkk2+qAQxOoSY0JxnEAxJ5IP4PT/
HpFIawR32zF3qVhxUF8HTeNdulLCSOA9Y0LouFXrXU6IDEX027+bavRjleKdfgNihZYYYUIKR48A
qUWoReH3/u93fdZyGjOPsnQEkUMxzST2zve8lqnx4m07bqv3wMzhCxRoYk9V4DMLbQ+oAvdrQBzV
vUIpwdxqHs9xkOVyTY2//RbSTnuahtsZMOhhnxCqFA73jmzp5brxRtZqP6D3IO1VVutkpcTxQxvQ
5jaGp+F4tQyOvgxKk7t2IsvHRdIKbpZ6m9eHg287FTsMafV14LxEBG4v8otKJ7zXG4UFdBmeiprP
05ZOcbmHJ7GXrzwFr0RVb+QMPWDVy9p3Cne9WcmIDE9JNm5bmKSHyizitdJ9EjL6F7rDjQt2BCAn
46X9B+BJng7DGPqeGRsCZa5OFszBQkLJvIcg8fUBLzeYeNmSbDbcioDS8E4bFfKYxnUv2Lewq7Ac
ho2FoP/8UUSX5BAABWPt8lBq9AH+7bzzII4bXyKJR4yh2RXw3sAslwFNGN9RCkCtuoezlfdv/bcw
WtIUavJLt53R3FlRzw4/bjx6l+mEZIlUb1cocWr4XzHiho4smWY4oF0ojWXdIRS10IS0RYaEwbVz
k3zhCtP47KMqjsJOfcqByT1vTUVSUVtUh3hXDB5QMwsy20Qsc8WqWOqmr2CDAo6s+tQp0FmJpoBJ
2jFafT8k9ZdvsBlJ/nbLj0inRjSLVGrcgB8fKhRtZXiLs8lp7wtuqP8mffXpq20j6yXkib+Z7UVo
4tTaDTlDqq+skF5/0qpezlUdvLYKP3d5KuK4MqovU1HleNaMhj9io7Pujp3mLTdFRhD2JtxqY/vk
Cr6voV+31aIlVbPqGEIU/YbPUlnCwpyLVmDUjk7Xa01hc6iiFkIqXNWKFoty3AdzC6SqaQGMLsCc
lvXPKXV60s6Ci8i1T3IqR18G/X9S7RlLZeJBBEDuwwToPQPl1YJhLGgXUPCQAE7k1gv5pOpNg43/
5zuSDvLde4+VijR8QBRXFm1NyJJ0i8Vo1nQORfy2oOvXTC+5bHkACBcROu+7wX+ijieHjHhfFo1a
wcinVZ0oeWgIi52+gy3hZFuXL05R3D2zJVk9UIXDpfarfJ1GgLk+kAc6XrtsiPgPA8DpYNxzKsX2
NPqtQMvu5J3RB1eu67ZPT+3CXxDPIe3UmvzuWZfPiWDqW6H+ApiYSpe54mVcpcDEckZJlG1COYNK
D7cEFVS4ygbMyqMgAzS5F/K8crlcO4rQ7LvTPTtdXlLQpXJ6T6EJ7V2UE9m5GiKT4JLG8/ZgZFU4
GDc3LRgumOdQuKsbXGYV2514lJciRDNAJQdRRIsOjI4uHXM37+tnsIEUBbdNUgYF0lG0+bskkAJb
5Uc1iQDfcpc9cmkyOEjY2B40A/zOGdMUNTqd8XrTw+TI/Nm3cXgXNN8mUpjXa1F8oypvVTse0920
22Hq28QSTeN1i2hBjyvxw0HMKgkd3dbDpadVQjmbHw5rLYTDDKfu9rbtJltX7JCXJwMMtbb5X5v+
0VaPkP7ezQLb9TFS2vfRLo2HwxZjttp5LkS+OhykX5PVKQLGbahTol+QCSf19rGkBPy3RaGIX87u
S0BudEIZgBlwzkt+NGekVJlyBFkCqcM8W3Zh9A6p5ASGX/e7UVWPeOTWkf6OTZtca4l5PkTBSQFs
lQHVDIZnGyRpWcNQXaUkore030ZawRtJpCENUSNxFm7GZRjvKK8cxaKRXE3chCMGHcpOL1LkC6UY
atN3hLHlLt7ltOiTaqIE/hdjLws0VmgBdsPJNfZiy86iNjjsl1//sHStR4OnnjzMlO9OPjpwkuJL
3pWxOI2Ud3xPMzuBgRLemzNPwkBwqKH/kvgTsUEF2JBD6e63OqQkBhEWb9xkl8cvlSyDUrDIts/X
dQ5kFpqQ3ABQI/Lzlx0C4tp6S9NHVG6e/niQPNsxSwrTRbY2uKUJRDlaKuAYxJgplBNO5b410QHW
uqWWBlDZIS87WYhiYXK+Ied9nRL35fWzp+lUP4EnD8nMdkdfx3C4tojrP57Y08b7KFsKBbOQLtQM
70tjVghjOpZC6UTRmHbryK18v8VhGgKQisYyPVgYe3C7NvU+yzAFHM0lOo8ZtUiFPG7OuivruE7m
rmlIBuaeEOdSNZzZ2gUjZV5SOhWcyuovVVAU8LkFQWnWvUJh+Z5iP/2XZ4XbSeGtAHVD20nc7ULz
VQylzggPZaIapIz2EHPeEvyOqRbIpV8G9RptPNEbJBM3iPtNS9vswtrbB1PO5FbAMxCG4d1dXNQD
3UdrC3KazLSC2OqvGdDcvNWgphX3Ru0HV4JR+BvXsYKa8i47GD3UUt41zGB7Tv6QctY2ukwuwWaM
YLoCg/RCgACOc704PJHa7/K7Esbk9LzU2bX8bFMLn9ebVTSwE8RxVKd4Y3xXJh/9TuCOMpAr4J0f
iM6nqfHAuvmwCUCW1gDh8nDUczHYfmZnJ/4Bcemd7yB6H+Besxaz5uuHe66viDd+HiK6Vx943k/i
JaAipIvhPOnUKSjf1dYTa3jisH6cA1QXuUw+QDd9Q7tnjBeki3eDrM8uW5nLzZx/1E5f+FvLKzBW
EqqA8FVFCm1iN4eHgObqO9wLnHEa7mRHEg9kzlkD1rdUTmvb3Z+sT+BDHSSFZnLxpGV8AGwakfVh
sDcmnWPpN9FoxqYnw72smdVt1ZHscOSC04YLbyL842rnuMpY7mqrwaqMQAcW9F8uUPxdvhWXaZAv
e+zLkqOmW7fw6LyXnkAOjp5vI48azi2BELWq2n28eEzC6yOqujeKh2GRyhAvMr8Ve+rEb4Lo9R4z
pfbu+K4ykRDbSR12Hja0uhTYkdrvEfQ6vKc6t32TuGEYkos2JOUdRXWtEXWthtRCXdH6ZMeJ9bxO
93THTElbLCcCzvwOt1GCSVc9CB8wal75k9cOoMX/3gIq/zRT8C8fTCEmr8OlWdUBtUvWqlyQBPgD
CqfXcv/nHV6DqgPhKB1db0sbRq/j79gCh2w1UnbGoPE+rYiDIenXghrQKjDlULBIegMewqoIdtbX
9YMU/VsJMQEHbNdDWPF8oSfC45BKwa7l1vkjlkX3RuRTwVRA7XCsJtPZFhfGWqocprcz8mN8y0uK
G6yYbvRIDgaKhbICRvsW+xPT8wRRAVMC0Y5XzHFt9lF5KgLr6ogMRz3+2wyKZC3En4yWV8J8f4iR
NVnBfPgFzy1GYzRaT+Y+9K59ROWoWy3zBQfKx25xQV7e+feC1lYxYlKPBHsXkkDOFdkrqkqRm7HS
Hh9do9B4Zn06Th1NR9bqNXYxGDYnG4vx8Ic0jolXR7494OvXqNQDmRvlk4CLhQV1kKDGxIVphmHB
cKgVWRz8indtM+L6LDPosv2ObIZdT2Nj+NY8pOmW9GRx2umLCdnV7HX9z4AozTYHyEztloX9qtyq
HWqlnikvp2byUXgHaL+EiKcr/UWFCYR21lQ/lXEHPw3l1gb2phowJD6fC8SIqa0bvnvAb243bg/S
wcQLLrJTgetvYvcflFxWFphuo3wNXCF2aTu2tTqtLIZfQqw8NY3cgkNuFa4BRXvyO7Qj2hZLCCt9
XPbOQ/gCGo8IT/JH0EIsFmYDEmi6qDX8UC1gi8mrkD6trujR6nFBGXsd9AUiDFyyi+cFNxyeoSXQ
pWy8O8v1GNA9GmfXhgpbZPLC16+21jQYkyP70Xmaiv+krqsBocaEktEIWN8h9r6FVcAIBBo2TX9N
24bk6kuSPld5Gv+Xcp3RALySzzn9qRYxJWe2WW5iNn8RBoNpDe+T89q4Qk8RnHZ6anj070CSPYwP
MPl6vR46t6QUE8EZizBF774ORu5T0TORM+bbz2na53XqEdtYgl+SEWNRUunTdcbTEArFyh5u1FwW
cSJTO5D9TMO3y8E5EXcIa4AlwyfRCECUyVcwLuqwiSxvweK+jkbELfWTqurnBV0IXJ+9JMAlkv37
QSPNgdN5H+1bP2jzG3qKnNUwSJrqRicOABxxz42mAqZZ+k1nidTjTekeHNvsQ4La6plFKyzE6a+s
ayJvwzhEVHT8ca6bJSZtVBrUY5CvILjCyIFp6Mg1XmAXdf4QV6KrphrNUtrAL8ZhlEoJRjOpk3wX
6Azv6UO2ZvY0Hj0PrnNET2Ko6ApyFlwfC2WEgOLYB7xsNQ+YuRYyVoDyw8+raQA1L/GK0KLVFdiA
nYDVey5Z5qhIcl+B7wQhGEFyAKocabFhPHOGE2LYyKFT7Mqp9fl/D/In2TW04EdtsxXSUqH7ovon
DyxN1dJtHsZWxDlaveoitUdTp+bz0WMSoXlSCr3XiCH2nUZxaOxm9jL5XOl6fMMNwPbbxKYCCJzc
1Hl4jGXGoqXyTH0z0A0qltcCjEBmW3iUOWbLMp52he5V5iDM9r7vSFrQoUFV6AaSKMcZDs9vRxLu
SyaiMmkSxS56T6O4zR7zaa2f9PUn6qYbB91LLGVxDeKkZBdxoCQgLNlwBRkRkIVsq8tkxBPmQk2j
mgf76Q2xBfY7FfpKhY/iR2cV2t4Oupft/eqYMJIIIZRfEHQ2NkVFC/X01mNkw7Vv5DT9axnwxnv1
MzfpzA2EzE7L0C94lbrE9yVwMOmJtuWGqXJoEA3jip0cRwECf12aHD6sAyGDjXIuPYMZ+5gxWJCv
VN5U0RPSn/VYnJAEtaclv39M3GqrgMVUF0jbjFQifKxrRw/DZ/UqNFnKBfWyl5/lJuxTaXCJNO3N
egKn9pRhr41dTepNH/U82XG7lFNm4im0JTq2ucl0bCz2YKlg+H5K2X5cNEfBtY8omTQfKUCEml2x
dST/J/uJIamiezt/7tslHvzGIPbSCkmd8zQeVGjyoWkTtrTetZTTWA7cJw/puvP31RjWYZtrTnWW
4m+8Li1cNOdEK04Vaq5GUq560ux5EyvS0t6dwCmjOUge/8ftGjJm2pj9/6CDzduMJr91DE2Ewt4M
pRGvlo2idGJgyVt3YPsLNFTvZJAxUPNH5+IoUWvt9egULwHcap+CzvbhmWtraBNTp6wBNTFs5HK7
a9CffyF7QYIXlWrPJW1xTcIK266nvUlQex8CDcGSrej6hBhdhUrvoyqvuTouLgKaANBerlAtffPJ
doEogcIa6C7Lug3AsWEUhZ9QW1A6cMk6db8YACO/NR2iRpKHP1Yje7Gj0Horhl+1apJHhU9/jZcU
/Zx5EUkLgBixJ/XB/Os2ysU6zwCbKW6xVAVkKZTD5awduY2QlcEu3UcxDLdVFP/Do4iNpFTxlTsj
CJwGcgR9yjcKdm9TrzgwgRmvFgTalEdlQ2VqmAr6XIstrQjrjp73+A2loM8dx2XIbYmHXTgXp6qG
qgs4sAVt74h1ZyBLqxnbpd1yollgjIwNimhyxQuLDhhqpt0YEK6LDDSe5ctVCrSxxVbAKl9MBsAt
397+wswFDmgHW/HuM2ETbgdIxyeJywSEpfNmC6QSKMztkl58MgTvlO87FL0x4p8T0MWaSKzB9F/G
6NKBWCYeAnWCQZiiI5kSSpujTrkxpp2gmr1Zs+1ZfISxBXZCMDLfGNRLmPyLq14kxMirUMWr5TO1
c8tK+QTeaPPOiybxRhspwtCB5WIjXTReznM3FNsa3RqKOAuMrKAmBdmMS/s9cz1SE+KfZSd7a9MY
dJ15JC/GPUwbaQOD9so+mgcy3GeizjNYWOp6ucYwiJQYBDe9npAZfbXC2cERpbGupOybFE+3wXAd
qGAmng14G2qE9M6wOBvMuIKOBxBd1weP5n9rd0ubjiQEDTl+9SZ4t2u7nWdcpjB0VxGHg5xoAzb3
TdBWlHDNrY7LMdJ5j8/XraIcPswgFwGxrWdtzj7/9KGAT1CTQvlwkii9r1H/dXo17pBgS8K08TbU
F5/25QSvzNe5W17cznktFQFj4J/lObJUpSbr1LixpFQFnc56rByb2eXVlge+2iyhFLfovdy0x3G2
FDWS061x3Omxr1VQkK2CZqs4QrqrW6Jn3KX3U+dB+a6r6goD0w87ULqdamm3+I/0fLcyOGksHlY6
fS4G9aPpq2XtFJKFzotCXik0fp7MmUGPEHjb2cIZ1sGdq5JOBU57XTXvUIHRG+ukm72ipHhtvOia
aGowrSttXL88OepmLwKt0II5SiFBZ5j4kDD3wBgqdh6bF/Kwdu8Zrbzf9TmhPDdz8mNq3Q1e+10Z
nw4rPak5PPzrsq5Rga7Ec8HlvVqdtqulNWL8dNOurJP97KUjGkKIF2Lt0Ovq5WrYXgqmKKZH21Dw
J0/e4M3hRMmGdvbv03VKuBuYktVwh5AvmiBD6U1ranJwzA1hE9UEgC/lMmd/ihPFdx3VW4P5UiKf
oq6wsd8mBPsRevKasWv1Dtuk6lgFoBNzSZFliyPUz+NxSIr878CcmJLpTpqK2Sft4Y15fLyY3OR1
G7ZsK6kJXI+ZMhvps95dslcJnOz3FrCLexPn/7bexyj6yLU0f+sPImcrELBK75SEdKTfmJoKs+37
4I6U/TbuUxg538kOV6QxN5asgkICwJvPw+SUlejsQjXfaxOyzMwpCuDzDHb06lEMkb1TG/Z2Qp2A
0Z5oKWWP0GGvg368Wmx3HUzes5WQ6amgWOZKv7czpatiXVNcuELHmu0ZEJvlY08OeUcEfIDH6E/w
63QlHb5K2YbymJHFamQkbYzRyoBBSEmVtRUJ6G1B4BIoTKDqILkuNes2G1GyQQvE5O8YpgSkITZF
cRVgg6s/Uyb4BTQdb9HbMDVeu55yNX9cmZO8P0/OQaqlTFdwBKaG0MZLJSkzl+ADtZiKOh3Iuluv
CQzWjxwrRbIV52GSwSOg+YCNJwkaKrhE3DjrNbhp54zbLnytCA0fdOxsRQG81EJsUE1tRmtszwYl
s+YGZwK5SpCHSQnU0yTr8audrVErSQfLAOEkHlThSKgENABSZeqfFB6bOhLpq1H20uruyL/yQqOz
vQvkFWMxEpa3sUTuI4jiwmHfOetAcf9hgB09pCbdBeHl9+LxKFiJnJLJOYMZgbu/jzfDZeuxFJnG
LU6LdjRFAQJiJZmde4bXRi0JZpo7wA3cSjAFWPkpoJutybDo27I5jycewnhcjaVXgEBzkT9R5JSV
sbED44nhshNV5/FpdIwvzGj5azJ2rYxhJDUQ8pDjQpaEU/mwqDqnYyYZ4+k+/NmW0PmE5oueWajL
3o42si9bFsa4VOQOOsn2R1IYoDO3lPtU5X9g050ZfpUlAEHAC1UwKrL1oYuwVbcO1940LTCSKQEe
8UXF9E02j8ZtRqZ5jV2qgAeuIZ1gLY4BUGDDLgIhWuXYZqGCqF/waSLpnmnzt8MaFDMDl40ad2vP
eFxAfXXgidJQ2PR6rXdRFnrLpfb9sXhVYw4A2nZZK4b283ONXlfM7dqV0WDaQf/R3c5s1ud+LKai
6r3AM4WnvMSS7lbYrDkvIdNqMNRbVtkxH0NwSlP5v/ZkfAKobZHorXT9eicOo9Xk80FpWSNcZQxL
gCbLezQhLX9+4N+VhkqFyH7ZNVZYHds+ofyAmAfzc6ZGJ856HzqV8xMDStcXj7mHm6Utyy92pNeW
hnXYxGNadTWJnQ2E2Mn0Tp2kpHdD3NFsJB734iGWMicW6OdwI1rcDypNvTX1MuUrimA8QAnNDZUH
xZ56XzACAkcvdnShLoC28M1x9Jda9xLRUC/LfpGDEZAtv99+p0EF7VuQ+cVKEW44/CEBF1KGEpfP
StZyOaEBIU2n9kQb0P7jiKJsv23/LpxY5p43JzVd7JJxYx/PJ0JXLvoK6UItRBIyfq3ZgbU1vTag
w3dkuBFxX7cFae+65WItK95oD6qbNRbYWyU18YM8ogZSuVbC2egVyjZjjOy1MrhJxYFvugePIBbN
akbz2rN7eQax9EfvzDwVOqb5ksGtUTKiNLw91T862XS/EUmnq7eP4esJZSZhsa3hWmr4DFtExWub
BYKdBOZis/8whlrBlL3c7+PJbmohxBO7ELuGPn7jRiloUeGaUIUeO6uFCLWqW+GFZ9Eq1is+457A
yXnpDYsYxReotcxHfohzebEl4/I/84sVcUAGL2I8beVnzPCCBQ/yxJnt1zueXzVc+MZj/M7a4FRL
w/Pn29oJ2+Y0s9PDH7SKdf39jo/JBztZFA/FsInYRTY6T5eJnu6sv1EblHCxiWsXJTfQMQt3OSTQ
DR3cQDvJuI/XYd46mFu3g+hO9cpJpCYONBu3YtGznYBuycyXGnuz20AuGuyXTfpthaH6l6dg+Mdw
b2t2buLpx2e1OxWs/2M5iEMk4jfQ2Ao4rhf231TofuUkQFRijFqGX7NtOCsOCDW18yItRxZIWwrE
4ZFmBz/ELRk8v6i50ooa5yUlUzleoBXXigqTKbpT3fWkUqTjqKhIsUwYWSD4sPgPFHLOOqpU42Ej
FNzOwrjjZz6SXNJpmDsPh6PuS0cHwSjvHu0FpUzXX2gh8suryHeTaYMs7O+OPangDfM8MNTiHEWU
LS3qiD1eN56PplOkf6vgt4bMBf9bz/p+Vp74cttzy6J8tvA/Vx00lIoexXJ0rFpD6J+urUWaXiTk
0Z+fSIs2vIQ5INp9gnq+elYjvdRVGu5PKWsO4CPpGnzcptV2rd6Gjo76d4A84UPHVErF3BsM2+3a
x+BMqOBvxdpxWNmyzppuLBgCAqrfJQ6quNElurzonBiANe+8DsyZFO0lg58B5g0ZABDRv66hwB+E
BQvagAIerMW64PlEAKb0PFFP7o9OXG4JhHqCA/eDlGQcunH+cHweVhENK5+2dAwYpMruIXufcRKv
VC/RO8rQf2Qyf9x6pA+J1T/cVANinrUJH/vnzDv1Q9JDwUJ0AZ9lV7eYpCpWXSfk/I3UPl0LdIK1
gozCUVQ4hR+HNl7Bq7I2gYfN9kVbxjNDPiNLqoGEC32gex3204VrPrwbwEhltqmgj0kJdg+Iz+G3
Q0nmwyhJLFGz3V3+Bv0GJVrjY3RKKkQasPp/GUXdj/vSdN9/issw/J+DpX56QLRuMNYEByZ+ktcS
jzX/L8s+9lE2Cti3gD75oxAgIU4nTD608OaOzbLWbwphgz2GLSk5xaEjCZ+ASuZOQ3v9TUNyXAIZ
ZPHmlTpld3fSADm9MoV+XcD4qJ+fdrLvbbGVL82p+1rvLZm4YeQVLRQgw4FLHxZbIgBp5A2vxXwN
8pCvdvK/kV+0erRKgMhhLuDC13Yrp4QkMNexB4HHj79LFNN0Wo0cpOUHlfCyOn/6NDoWNfo2Az4n
20Wl0j1qfusqmnvSWnxXrQhdr1r1NJ/chlrYAifXs2aqah/N/Xbn4UT1E0AK6TNN4oix3GmFN9Or
WyyM3tMg4SXVEKvUwhU79vUEEjDnVM9t8TBKrm2LXyIzStXEh32VX5FrRSbFq4BFckiJvLz2/tan
4+I1pt1JIPyOp76vO6RL4mV+3OG9FrwpKjn//9WTVbOFyTYqpm5N+5AfYTgsRR5eIhHOaW1iGvBx
tUmSP39KeZfjAIRneXOn2jV/iWHhCJg31CEhGGeNiccTwSprgZv3rcK65QT4sZOKQHrSjGSVB4Yd
6qQXQC3PHYT2F2zWEcwzxM6IAGQKPmWq2s451eqxNdZw7d/4YNWdS6I0LPa/IVd74igNEAciSC9+
tpgT239j6zYHUP4iF3Lw+sRZ2F4uVEUpEVa1DBN19hO1HRemtOZo4MKnEW3yuwt3lrpNnBBlIt+1
cj57DqIEBGTL9Os36JdEUUKi7AEcindZHCwKHnIk+Lb4gJ2KwOrE1Lfv1Ci0Vi5H3pM57KKfiEmj
v+oF0l+EchOCqjZV/oSdd9bo4MlwS78Mbz0qpyAwD1m0lOhpmvuzAJwuXgeLAt26VcP1dSyCtOwe
z9u944X/xlHO3C3MvMazgzz5GYIYAhlfsKaEUvUf89gFQmx6tUAQPhnkntlkWLktnjgWOKq8tBuR
4BWeYvR5EuVpprnt385xS7LWIvJb/8xY0xk8iAqPRxAeTaNL9RwdF5+4NRBZd0f3dLXxZ+usniqJ
7X0LQqxZftLMjCse3zV70jATGa3az8MaTtsob/lr/TpbBWpiy6iauKcDRwRXfE2cjShhr3wvWHbI
F9wLb5s4X2DSVpClLzzaOGYFcEi8KOkG4H1YNf7v6MI1JeCsUllqCYnhkmOBIN/LwUZPUocxkiFG
TrsbJnwRXFDl7Zx+If0HT0csnd8yK/r6ebMBLCliBfNiafKzMyf2xPYvNg6sHVpZ2/OnbznYbTqC
83EXKX57GoAKERi6fX+w9N8k0r3zSvEIrkVGJ3icRKcYMzSOLAF7nGcYdN+1emSOyDnI1TdJJq15
LM3BdbUzcWmxpm58y3Qyx6aLHTi+9fuLJwgrnDcLUMzL6mjwxe8qe44qWRkQssa0MZ3JgsYfhYHd
RT5XBfOOft0tvhpxIenPpqgePmn0qczuqje6KT8JbvcY0I/oxvr7y850FEZ9TIgyTR9OSAlOFlWX
AW8BfAo6jCEY+ZNZ31B3Hg2r/3jRFBRSJf3s8oiw38Mf0X0d3fZBGPXT3NNyaNycMqG2q0mEs27d
Ge5dG2gZ9Fi9DgN5ZZ8vwI2mW5+NwYiFx2ixRrFgUdalxkPhhhMnsNdKPv2BrWgC8jSNpIZEYBMR
80Ns7AMqwpUI3ZMgtaDA81OvvnmKWNsvTYMDru325fiI/RTXTFXD6ml+B/QquqiHpUHe0enEMn4I
tDVZzEMhll2eiAeQl97XBWbxC2ZGLUaLzOq1fzgabHI9oBQjodS9DVXUrzZRTn3D4kbNLDjEV1/D
CeLucW0UF62kYXUCLV9Pq7KRRXADzkHzU9cOo5CptHlAu+sDgq6HkIBPlZlAQMYuzVMm6LRNHfUm
lFwB3jicT089XmZB7a0U4g8Db6Ql9+ybqGNwu5+2NwpBi5OL26juUwUgl263yNGbR6EW1q5m9qiN
2sjxuhn9HvTU1b/JmufGHoYwQmRDOX4263sy4jicag397wuKLZbifYlT32dauxF8D62FOLZZJlnK
1P58RPcJx5gT6fdD4OCzjhYPRXTm6DSRuyIfO20PB+lJFKxPZN2kolncEGBX7TzYFRuguBBd7flk
+LLTIKiD6aSRU18JKutyriMEob62eMx/6r9LnXIN6cPk409w0InVyLqW4yzHHSCE25IubLysOsVk
P8hCfq7x1ALH8w4WLDIMn7Z64WFEndN2c4mt2MNP4/Fo3/WP1qb9cdr0GsNpIVt1HjZjZCUACFOg
U0diDqJLRcssqRPXx90vWnyC3kRFkylTaHYFUkzm/UCEG8bnoGY0PVkWaJxOHNKO0+v0dnuYVt1e
xViNLsz4E0s85Fmp6nU8IWlSUMEUz/fBxpQNAw/FwFtAcOgFwodJndiCwDJOmlmAxHd/eXwQzZCm
yt0Wk58JXyBL8KJI0jln+JGerEtAgSCqzEpP/xJ8XbHUq/InlLCXHFiWSWgQWvTN+aMdsoBqk3Dm
Gu8SgOqslxhyfIVik/9UNZUDO87RujRTKmziD0ROEqmmfVvb/+TGaf2GciB0zjK0Sg5XLZjr+Hjp
5GkwfxzX9d7+nBxU1pDy8rVF7d2h4RnRg66y4Mi4Hl151YhwCiXfW/1GU4aJ0e4lxViiVmbLZwAP
Glps7x7I7GsH9zA0k15i0G9Kf5hjxrbFqVkeBBA3ySB/cjY45fTfuZuhyUdYcf3jnUS3Is+lSVbb
CFPbOQYiRsf/XOMBvHQDM8sAh34nZpfjZMQb8AbeORkMhpm67VcyPcapFZIjZjO4cQEPmbQqER00
xNmsasxZc31osmdZAogUAex/7jdVb1IV4+HC1csR29Jg3O2YegjHuMRycC9H72Ym+n3fV5nQzG/j
OHrSll83WpcFG6OjvtTHNdUss21fiwlZELtU10dOMY1ZRcjT8PciqJ7xr23C0KsNbmnfaV3lEFia
fpIgiRJjjzafb/uTFi3QY9t80ua8Xc8k7y+VwjWG5TZOFm2oQv5Zdl7Wl6j18urjXwGrMjkD7B2n
J8XI20Yw4QZnZgUqgQcBmYQEuPmcDIFh81m1XES4SyxBL3eZwBkztSrGnmffg5Lpq1jwZda+IiM7
9zuHn+9lj/b2pKQmtxtMu/g1p5u2I5eYL6Oj14j7qq4T3FufWJ1AaJBjyTdnHrTMr5VHps5ZdqR3
d1Ry2QyAfHXV8I4CO6ksNTIkJeQV09+LUCxYR88i7hePrLHQzoZybs8U12kGxVyEGxwv1unWrqRS
eymdznJ7g7ujOWvOx5m/WGlIDWcRLji6qsiR925QTUrM9gI7JfxKjd6YnqT9iM3JisUDdzNTB7w9
axXapt7TOiuoMdeC47sQgGKJ6gxis6Dcp/OmMLvKllIOfteXMTH3ybCjshz6y8+hUTbwPd7TpIr5
O6e3d9DDzAVIo5EnsryyX0I0gQEyKXWjNuowbbJifiZxY8EIEyfzgOWzvao/0R731d+qUnK7hjD9
q1hsVkiPcRoAaw/7d6Alt5gn92qZhLixEkee3hACE1xY0/7wK7yMq7rjjCRhFABhdTYh7NsIKdM9
KVMFz+66tb/KlLB5BrfE2JaEfPGmx3xqiJbIlfDGyUKiWDdjFRoY5q8RETl01LZzSRkuYnVlwq2E
jIznthmB/Au6JVA5cbfromlu4eGfARtEIzbn3oZJ8ZCban5s+bN88thpih7wuYlrldW6fZZtEK7z
bV7IhBIDkTURi+gT+B2/BftwlIFeImb9CCvD3uMTJJYhyKSZ361HZ5jVAJ12BFY99SpK5j00zeos
UY6l1JTsVIhpipY/QsxojZuhved4rEYUVS3bKOtw4CHy+ALOBiUDMwmFyY3FYS7V19JLKl+17s4C
o7vBM3eKYSQy6Rykl3AAUjG7DpMgpcZGDkFD8Jd5MObf/t5cyIG14UJzBlc87+YBcCvHTe8tVYBC
CxnPMS2iowXVf62GN44u2q/TDS6+rL6f2skimdOEXRyhCN4J+gA4a2MaYTJ25jJhH9K2JaHNYij8
zlCiMioVt3WVWrocQIQnQHK3zlv6pZtusqBOzvZ7KpIy9q+naPRZ+epKPvNPe1MK16L5jVfUVrJF
FufJKTmt0ZBHs5KzlBsS9M8JERJb8zH3I9ahxO2Ml7V3+yejR3CIjPpJzI8gtvzdGIYLczgmCWLw
BpydAuQrTOS99XX8kgnmhqjppLVxTfvoxLLzsyMG7hXPdYFCNzbJ2dx4I1x1QcfZ6so6wIqJFWNy
mq6pLKxiGSK67mktdfEf1mmJ9nRRRSLbAAFrtv+Vm495k66dscoEoMaaFERIR5FDw/lxzGVO5j3X
TGqBz16QBljJ40Qhd5ZTosTbM/Zbl/PyM/9L5FyoyjDac5aSz3zMN8JhxLJF6+V+wEyMZW/wVRJW
/YcxTF7XxrvDfF6+kFBu3N/rq4twLOVgIgmjDoWTZNJvNe430PIXxhskgJDFKxEDlQHkALyrVpp+
Qc6XrGQvbCbUXS0XZVGX/lPHVBiKD1vcVzw3KHLwGRSw92IzaQC4WxHxVqSZA5lm9qGag9RGFVZM
SSaK/3AdVP22l9WYSROFz1jdCpzV66ZW7uDTGA/b0TtyhzIyl8evn4HQ79rbM/u2xSC8cr8TQm2K
jyerrB5gB3I9RpIstgB1fC1DfJhUiZNKzB/INWDUsu9CdAW5vzgtuLWCBtJOMNl2D6O3oaPT1URL
0qXTLS3JLCwOX8d3Lbuin6SToWkyblnlAi1TKcJ/rK/Msv7wOmve2jjU1LyWoRjzSsNA9uMpz+AA
iyLUx1QO04jNGztrBw4GpoAOFA9lLB1uiYP3+KMk7BqfpD7a3pNn71JlW+wh6wfkk44Lsg5jsAMQ
FPWSs3hwmHfUcR7ptblaj/Pbhdsu5Sf5xVlzI1ChxDF/uhRr3w0F5O4L+BnyWdZPveo7NyODH5DI
PRgqAx5e/d9HAoAx4uWJqTlBpiY7lrIt1YQx6W1ATyFPEHoEqNYa99A2HPwJMOqkuANqzRnoCXTa
LsvJ4VAxr6KPTDjaOzQZoJeCpTQhs9DtiSlLNoC2bjVj4NuiJpYjxR6CGGltJpR4RN92H6v53w0B
EjeE+nDF5WIuWqKW2Vp3zHOQvxJYjV9nkvmYtXce2b9KYG2MCgp99V6jC4BhlQ0lFwhqzcgTZlCr
w0y6H2ii1cV/BAqCIePbYgIhGjjZA40le3NJ1ZGkzYMZLnarmzHN5TgHNK/B1kCMxks7F2zjfQq/
l/zujmV6QmOsgaPZ+rswhqm1Ww8eLGmzaGaSWJXodGue19zUf9MgYzwbOhoi8gvOLj+QU18lwF5x
7Ez9HX2RNo8N4IPfqOuKmvKlAUAJrOpIlGrM46bDHT535WE+jh+O9PmxwHj/4hEnvYl1vSEsEahz
CCy6HwXN7QOAgo+0TB7TTsrAtKUnEKQA6l5Lcq4ZS5RwRRrHsnzAelmT5NM9vJFhAT4RYoVVlpGl
HqYno2WI8fMTlFgI3Czt7fKiu1xEMmb5qLiE+aU8Yo/cOgHJMDQFmvxSJ0GfSr1H4S/X5Q7DZFzw
j41nBVtl6E0ByJ6J0HjA1TNLwRdXuMfFIE1i/4i4IUVnPpQ5IH0Ng+qkSud1SduD/kQu2NlEdim2
XDX7AwSzLQD1CrzkxTSFR1QfY0grG1nnEXI86DrjZ0bcFMCC1yy+g60OaKlxYwMQIJC8saP0oSLt
Hc8GPewp+SBS5cE6EG7W5OyMr5jqaRpSifVxsQS1qv5DfHvg58tG0eOvypqEKfAXPLSCQqaqCOQk
e+/o1HuJnJVzbdh4AMss4yGcGGYyFlffN10dukyzlhVGKDCkE1OF25o0cyMpHKGGBMSFrDh/znSG
MYL6KbUidag03BZSEQXjWGdTgbsfq4lsR2hTlKm89j9I2WnFcxWXU3UrMGhYs6mu0IiVpWwUdMBY
BRiLq4laz/pXU0RW/QTgIrO4Fp3SeLTIZuqR04e5l/ceKzJN2TNCSfP+YRW/PcaVLEGB3wSi75fb
Mq6kOAiBWlSn3g3atLe9BZ0yv/c0poNkH1MFYzRKvPHiDHymog0Z8Me8/m9+BMOP2f45Swb9FV9k
W7xPJ4kR0gkkbjnAdRID0dJH/oNUn/Y7mcvi5I6RXacC1wI6J4zYksIiL4/TEw1GQIdkNAjmCqGB
jy8IfRel0lM5NNZ9K19cctbnTvvBrSl2qT5uyDSQbnoYmnVHLcSQ7TOrYNT90cy2ydtf9N+HmGQu
DY2qoM4OnWNL4lhC00FKx+/m2oUDp/KgGxVy0PEFkLhcdbbBYh9+WndkIBmo0cmqtP5nqgVbj4BE
cU0owr/rm4eQ4JU8yHb4HMxbl86nMxnzPAsrXRT7YGdRdI3k/QthKlD85kXUjbJBDvzHr47simnE
JkUCJlWyPArQWPEusmor9SNslhCYyxmSSKOsTNqlf/nRpgrUV5djd+IebuN/vU1RAZLJEG12eC2g
ZUB83Ep8qWGU8wU8WS+n0EW1eCG4KCDVd2+uIwPJ7NJJU4kTLhkV0abgoLjTXu4L81T8/tMI7YAs
9Guf3YUzpoLagdDkGBRW0/2vtnLEPtrJu+NvLJq7x6AEymq02ySkgWwIqXLHkSLQCekT4M7uA7wG
Z62xVXOiLv6HquXXVdu6RFJ0YcZNnXI9XsDhpVHe0BHAw793S0xDx51Z+uASTLQ15srY1Op+YfX8
gPkCI9tIJWy981E94s+qBDn0MBcdQRiwTmbpxmfnUt1MbpVIsgVcvSB5AvJLqksZr+iFuLo31F+P
pCP2I9F8mYBMb/N7oNlCoc7XfUdL3M/lahr1vhbYtwPwxbaSev0UYhzYiIyPNSqGrGQoOcvjK6Qy
UJ2RV3g8EdSN2nQ3m28brXNmlYC4fee5AgCypE39KqLAUWLIB9LqilA0NGnrdeULtoUtVD2ubPTo
I1IYBHSjtuV/B4/d2E+tmw8TQSnR9ztZr/N708tcF2CVrE/YF17rYghaUAjuMqSOwYrk5yJ7VQtf
xgSiHETRLiwRX7YQybf78K+uY4nBU2AxhkTnxK6ssephG7Do+mA6bsQj6r2047qbQYPFWi6MCqr4
cKkpVlBCYfPJnbraY0xETVc/0oQ9LR8Kh/5AaRR9ilxM3ULimmJnEkwDKtunXplRfBUcd7rEHgi1
4t7VkW/RCjOQJQ9J2zMfGKeSl9VcHvaoBDLMVtK/3sqhIMX4xJLzuHa8LhOnvZEER+7+7Lhw1DfE
AlDXpHRKgeP1geilqnN8HrAaQydVHVwVpy3IDmoPKOAXSqXvM6fAt3YfF6xjgXoTKGe5MDlUgIrE
BbF473EMAYLroQonvWIRilzeJORV4pUaa+JGAYYyf8RZ22BGsmcXckXMN8nzQe2+ReWeWigAEki0
avTGXYqccFvgU0satd6I/G8VOslgfDhAzjXYE9GGDA2WfZU4ETMuq9ZC892gyxeR5Icsw/Az5dB7
/Kuvpx97tFvQG5l58jNjybSpbrkLu4h3F3Lk3IapBtYjWSzgXfWuynOk9ELY/G/4wa1vtK4BIxT0
aLeWhNr1T2ug/SnFG4WaRjG75OCeAHKOtXeuVoTcLXThUWq9A/iwdBX9RVwvC30DkNRuN9S13k0m
1M+Wgjq+mo4R5vU3h1yIxqc6kjkhIXLuu77lXHH6p82+dTOf/4De8iMlyf2Ey6QSuT+HiV8onWM9
pue6Vc12qDIpu6RdagLfiKvVZ7Y/StxgwH+jmjLlWtSMGnKulCQ3VXKI14JaHn0L1NW+KUfWjA2K
g/uuQ1/UiXcf1byG89PbCMx5tefC90ykf52O8sRrt9D4D6TaZhxieIOR3nhGN/MQ/HVCbA+gTkp/
HSvZubyvJRb0ulOP4uRxz3Bk9/HR6Wi2lS5LkAgyp2HGcqNXuM3xcBS7yIpGDuI9/iieo3VQg701
etI21xaxN4VyoHc4npKgJYpfsuiZ9XAzugOtZP77kUxXaVvE28e8TSmvQkxr73DAA+IS7SQ+vcK5
Ay1pIelOlcvb+ECK9x6pFTswJ8kpfr4HDm5Lvv543WHtVV42bp9SqB1tYF68yaCrhHqnpCSmshvX
d6ZbTeTkr3BMcLX2PlFZrBmymG0lsR4/IH/MKgjccO7+uWZ/cxG+JlhPJln6bbpqKr7XZC20Jazk
C64F1EpJGmmQQzonahv818Bma3bFcv/dTOXk3XDndLHiSmRhhE2nekEUJjKZEHb3BS/WH90DFPww
eJ+pbwXtvtODotmwNrt+0qE/crkygt4KdWNLQMQMTOpnX+kNTmbFy46deQxzSkzbCGocTtRrAzU1
zZ8mH9oad4A3UYUKwIQAJbAbwsT1HGJwv6AB1bNuKAT+2EnOOKW2VJssT2G6Vs6E/gTlAbTHijlI
2AhFisoPKmBE3craDHH783rMPPMfn53qQEc5dPPSSYoSPI0Eb5C6A3JOLh7N78JFs45lzZLaBsZy
6ui/txex1jG6k4TxOG6PvqpCYamKUHjwbmlEUJFnv2oSXadXjUPIc3H7AUOb+bWc9rZk/Lb1oVB6
Y5o6gZt3jFFolYhVVVOaYMYR1Ehvz64R2Y9ozu3upn0mBeua3aXOQV0mBhdBMsiHQTXSG97bqYOA
w0fKkBWtEv3v55ghCXb6eoYG7KqKGDO6JwQD/pTPcrkcniJIgn1aKJ5ZGuZpi3pKIj1FC82rSnxh
wgT05ACin1Ei9Qzt6jW90D3hl18yDooBPMXhM5gldecypxBvkrKl1nUKMlQ/ZLTuBXOB5nXdvNS0
yQjUBx/PAZyxoGVbC1OZ1dXopc2uPKSgKrXzU2So0PwdicErZEoU4tgOhtPwHTqFfVso3g+2ZW1T
V4RCpRqbEhco3cq25yVnxzBpz8bC88mRKWppTMRn+TXYVzwR0MMnPAk33lilqUy7nO8JoRbnu1GS
ljuyJoys+YHdYBOGkOW+v0CxCGf++kdmuHJl3K1oYe+3TUNBGm/Ss+H+/IPvm6sUPQXzAo84+2fe
sYqOSc0O1SjLKXAGV86PQcYWU2CViTkjpgSm2i6TR3tDSq/uygIiyKjOXG8v0DfgJ8XxedOIn/LV
fiaJ24jOfvpYcdYNvjOYoAwmKQ32XYHzgXFlFce67meh/1kM8Ve7ySIjyuOTn6Ad2LIazjsCOjIA
FeLxM8QGIlsVmCamb3oQOWrDpqR9LnwcEtIuEkADPlCaO6Bkg0OU59s4tQNQg01WZcyK3DtmiC+T
Lu1K+bGYbdVw/ORzV/Rke4UraHsGpjbakW8KmW5jfP5wBKtrjjfoBVnf3jD4RencUL0EDJetgA6Z
ykg/MiDZwhQXZasC2mv8SI/NLl+frAVZ5zMH1tWoaTdaB95FBwsnAxxltphp4mLrjLAkd6my7ejL
USXxGVWvwpglSfluUz10TTy42z0Vz/yvG0IL/L8S07ldDC5jWAretZYsQYaQG9CHtnslWWeVwTJU
xJ5sVrAmTqLvxgan7iJPblITvUZIUfsWdCdZ/5uRL05PmtCnTOav9ohZKZvGYQvy2tBTJo5GK5Hc
skWWfoeiPwtQIyriUmOx0CPkEbIZHHX4jG8IhifT3fHyNiu63gkB1SLE2rLLnEQ7zJo0fs4LaH8Z
OE5g7R2OFH1PRAKNcbzlJ5kvKbySQEmbtz01iCUZc9L4puoKtCbRrH+p3KoDLviyKVVWRhbhaPrT
Y6SF1azoBOFcPCuUWL2iKC+9QdCDVRrv5gR1JFFVYlV5maMHoz63LKcXeNZdKBpyoy8uNYyi2jKB
gJxQwoNeDgggCe8XAjOJc3kklabw+mvoFd60WSA60Ra4K9XKh/tcYgRb7XLJXMuWXhVqH7BpdfyV
8lgmEuX8uBb8sR8M30vcQ8SHdi22XHIJfKmHp2qcnkAFxzC9ULrW11Uzjm1KXPAQU6Ln/xswgBYR
yIMUkpULfzFUaJf1vXsmQbQ/0V7qcMOU2I3X8gqIf/gWzCsdcDMZPPt7mxHp7xcycGEz7K4uVcR2
chxJZDArRUY8OAPCHzFKtggalaOj5bSlBwmrxsRTgVjfN9MauJW/QUJgPM80KasiFKGDyxcDk8lc
TMhkTILE3ZwGsoBAPRUMLCkNtgaPtEHlv7905i6dlIvoSMDnqNCrDl2OtHqsHAwSAG1x39FIeW1P
Iazau231udhan57MZkS9x5zon2FtL5k+IH90Za4IlGGSbc8/r0JbRgkdGy4O4hUI22zFrkzxDWjn
mvZvJQSjYZRVz5DSb4vTN7XDQbSBauRZo+8H5UP/pbCfn4BbzZPOJVsstdOYq4OUCGy2riB1afTQ
1iJXIcxrTOnleJvXx0AOthTSLHQ7icrUlDlbn+T2PT+BbbjhVehk4zjrzl1CU74NBb629uvVSUss
HMzTlkvJxq59VtKhif5lcAyKykOlYCnPDkoc/JaSo4HCH77LgGUpcdrKmfDVAwv7ByPH+3R2088x
TqaQrTgkuoPEe4ToXeHDtOa5O6+uIZS1YaowmyOkdKnslUAhbYFqyaWGqfcaMAlhg4E1CCHxN5jD
thLofuHKGwNLdaxTdNGIpo2hchws6QV0M+UF8tw+ZFXZg/x8y86198Eqo5ALb5/DS8dMwlCQqN4t
i9LuFCgLmJamOJf7N39wtIzSDyT+0mzNgeEUB0DvsJEsrzmJadZZw6wyngA6fgGijmpoiyn8JLNv
HTxBYrDLHevuhQdEESAYL70g/7sIBY6uHDOVPyO/m4xDoxQw9TeB9onbAn2QDU1RSs+B1Z8FqDiL
KqEJQYp9injcdBYDLy+wXuhSD10NAyCgc5cWkzYFz6ucCtGa1VoGAY1BJiDFGulijWi51xtWcUjV
Kpyz2z9pNLURLwHHRUki09RIbo8SV0ZDsKnQUB84rVB8Q5JiTvrDXnj8nQK+btgvp0/LcBYvUf/W
0oNi7j57S3J9N2rfTuxBqPzV7GCrrtNEHIVbmyUCo3QOQ5qCNaJ+34kvgrIVWjSSiKL3XbEF0Tf7
+Ej864TlFPbjtyAG855XbGFI1cgFZsQibqkra+xKLUMsFP8t34Wu2uww66ioxgmHL52zM26z05Wz
mQhPQdd4GrwKb//Hho91XH9qNp3BChxC9Bd3dH2wluYcEFHftPMaXeQCH5boLUu4igLi2oNUNJAe
+8/fFGsQr0avs/4vzVH7EtIMeCzIxEvRM3M9w00Q7qKO6J4p1VzqgGcaaSiYW/DCY3Iht5mxLNSD
EI0aMnDeaCxe/Z1NZzkN6w3HVb0b3Jlc1mDxXWHzzS5wOKl0Tp6P0qvDfQ7PVrDDG5jTZBOaVEK2
1JXcEiOsRN7wO6Y4iDgWk1O8Zjms5DUhWUFZvwCDpZXtZoMBTBZu3HjomtCsdq6I3r4oC/X8Y120
/QtDXY61fslycxhRhoKTzKSEsdEHNsnCF4+JM8nnvEp+sy4wzlZnKoPfUGhPakN08wNLtMwwWKmW
IQKoMh2q1pSWTqJdSTsuilhSGsvfGVrDoY2TDLo37/fZAB5SBcR9ApC4cHB/KDWwLxByPITVScgO
nKQasm0msOCOIMY6touhzJaWVZabvdhD6yH1bmzGCK/VQ7WsYZ9ft1Ghz4VaptgSImMlTgCqslji
WLMy5bGLnv5h07LLStLq8ahnwbWnGQHVNF3Sk4bTJwau1r4fjf+4noyDGbm5mtJuGUZAtKQ9Pimo
UA9xB1RpsKkNNXNHJqRpnGLavmuQYv+lpdhCeVAzRcznfGb9fjtdMNqQHBZUEW+GsaNPIwL989q0
uEsPZJflMtcFo2Ffh9YB/83fa6z9+FXNL2sBjjmAY7DPxpv4BXuYNMHivTvguQkk7FuttksZdmZD
d0/zj+UowUKT8sIylaym5E3BOQzTJy7pdO70lv9YVkRqli9dfq180s1njgfXxF+lSvrGcGTSCLjH
rAwhDNCjHTdB0D5/ISAJFqfT487rv3EXo7aWxs4KthG7r+YUDtxWjZM3YwU4cOvyuv+38umY5y6R
IMFijHPdhSXOy2JWXWwpgdnmB9VZG1FrXN62dFSdwtTYPgz0eOE2YTuQmwb7SYBzNrMcLsA5Kg0c
dpT5UQnZNHGD5+SvsZZC1srcLnjdPS2/fP6o+MDaEw69YLe47Gt/EzaQLMwM2Vexu1fM+70+IYwx
LhfXYDhoce2yYTnY4TjXV9hprqe72YnIruIA9WeFrR7f/NTa0QBXqqLSTPOY7JyPtz8gCEQ6A7ui
/dfizWh544PwWMz0wdCirO9ZY+nrXKZUGI8OLvbvELlyUqhqJvx5grW8Fpzp2CBBfcJxYNZx1phh
GYQ3Sb6JM10Q+WzKBI8vSEkA60Ud1JXzxYeVguN0RfMeq0PNyElVIOLzXLNnrWs0byWA4B7PN9v1
FIyBQUGAk5/2O/NtzYLjo7g0P84nbjEPNYdLTl3zp7ffFWgtaVBcoWOTyHGgMtVgjpZga8ums2pL
/6rcEZHJFyKZNj5f170/JJEdPKMMdJ2EwAOHgLemhBf+wkT0I1TSlWwDGJanQ1mfAAAES/nHNr3R
5Uduxs2+43rOkkIW/dbAy+pwr5ejnq+VM0QHK7ogQlvu8cF20q/xJXxCHF0clp5MljYkpoxyT71s
uIMm19gxLu2Cqc+MqQ5Z9no7GqV7d0xM2+RqWlwnhC12pJ50TviqX44OX14zodchN3xAP1SaAoLm
IzMRT7SymVll8PuxyvxqSvMkQMtHKH8+XbNMXdlBJzFiNv3h5jAhQrQ0CuOUEVOLHGptAgNiY/0W
nFU1h7uqnSjv3x+nivtNIh99KmYvNpmk1rx3tb3HrY9L1ajmx6k32AbUxLO21nwd4tnYs/Xk7BoR
dm3HW6yOHV21OjoSp5yTsmLQ/msIaJcop9NnaqL1DnOI6y6EOghIvgKG1kYG+ewcw8T8AAABTMWH
OO6GW9zYL9hQPOMs4qjhv+0pN/+w79OWsR8wreNXkek1YQ7mPNh1qgakVsLG4PyK4XbBS2VIXWuP
YiG37yCHWCfJDBukLeRke0XZGsFhsoZUOTOzqC2uy55iANGB2YgzJhpWWqSiPEtxWzmY+TxyQ9U7
SRa8OSjdiZOoibqwQmcoRDa6KZOHYZvxiR/6oH3NAr1/2DsV4WvubJYdsotExfeEIv+I63F8DuNX
m4PmB5wrpPzLrPCaQ7qNbZRmGHgtOdyXYPMQZrvvqVwoTUYGhZsSuW9i3MGlbRPRG52vP7BGL1xQ
oFkbv2kC0zhWvjU2GJO/P/ZvgWYt+2MxxQrbobYtvFzZblfM6FRKXLHZE+LSoTxzx2ofVlYEjkMa
N9KzvhXzUavtNOAEmXif3Z1XQRvb/z5fSZj+tqb/O4b2KjVfjBOa4cU3A6/StekHZx6KWATU+VlS
fPB00N+/egr16MFI3m6HBSQfj2OY7Bxo9TMGxG6Rz+JormPeZKreA94hYdcbV/e3JRdDueJ83aGQ
IFDqjeH7zmf5XC+grTW4mSsgOcPeH8qU37C/Oq3kexKIYHQ0nnImzWEH6BQGpKTcYLagrxj17Nb1
8DNcyzYNdHPBfrtwh67zUOBjYXcXvWJyiu7aqxmsL5rEfx1l7IvvxTSZ73ecYle4nlH/6ovFOBaj
2XkwvGrGoMQtmX5ASsWUkU0BTjKU6y2weOeYb0/qsQDflMUfVNS0apGOP0ZVyyJ9ZeeUa/VAjbXo
POgoFDnBHzaEFWlHUECOJsBQTU+txdXHY5H1Oo8Pg5+y10Cyv7hL2ijzOfeEBIPk5n+TouNKjudT
jUle/S7oTfBpMYzK7vhrqqOFI9FeucjajA8SAOmS0aicIt14Hie6BGq91yD4+bGJH86aDYexe0Ea
i6WUICGYf/wk9Y9/P9ZosTVSLMjX9/hkzipCK7xthlneqpScp/XKoioRgxVe0i0G8vlUpb75L5yj
ZIVmHhhgoYRqVcgaX1FkwNsvoeBdJfpczImPon0Wr1jvTkJuVO9GcwNsQ3Yxa2f0D6XL4eIeXGPU
cIW/dXGN6qp+/W3kJ2mB3NzgdvhuzYZqqPzzByrOOD2iwCSr3mLhMtmrALE/DiW13Twn5MPEEz0u
c9myBDmt8MjNbspe01y22R7f6JgzO9PDwu5pLz8pMdIYcAxemIKgG4UvtUGzvcLONB+NpZQ+DE1v
+7WcenOrYQo5kHwXqpy67lrZCU6Ni0+jUyip6zn0XmB29oGxqXCq8KAgMwKbvn/+r5ay4pB3aKbm
neu+a0m3Er+MvA9p4AGl2qCWOo5rCmBqds7yGwKSH1sXTUIGG/w1Fkgw5A85GkCNQVebQ1Jur6+U
1H212hk+4kB2HkpdxlIu+FqghR1VGeZZUpESSnR/8Sm14D67PkZx15+EnEmSYEWQ6h9xkFwrOP4I
m9pRivOmH00Jl1i8T7vgFfi+rgOpJwhZCHhFoxFSKJpsEpow3pf1jo7VBJWyoY9yuYFpzog6Bv6/
JnSBndVfFj7bDY5pHu942nmKbreLYakIw/0L618HyOIfvYUGbES/4MX5jeIHvba1z9WsYgxyBcVE
5VhOYPRDR5FR47ML11Wkt4Wi7aCv8BoJBtlVZD08VyIvV4eEJLZUkz2FK74RcGk7pvdK8LVwQ6dI
r86gSCM6ZeQYyrxV3ajp7XExg11zzjA5zBPX2AGUurgL1G8ut9banQTXj6U42OpKiLzOY+M33zN3
FjQwxDCqtZQORNfog+ftiWeRssWZ/v91hMf7RVpjHEqwLg/NNEnVUtEYwP2AuqqKz7JUopY+ls2D
zeW4PzkN/VOkhnVkd+WqrV/00aesPBk3BjWcSlS23XnN8CkZUiTZfm/ZdZ8MvRKTnkI/x+WAl1Rq
Pd8FbyHEZS7WBE78uh2akMj5513l06IBpKDxs8rwcaY46VLy+h0MDFBb/rKaeyDXxEKrTvyw+irH
jO+VMMo/su1W/Xrmmdiq+QZL+blI033yxJNSI5htf3ltGEqovO6oXKGiyAz/IgrOYkZ/3ufItZ7P
Q5eDChU9AwVEEiVi8DUN4rQcMQ/xriL2fHQ7yEGJEBUGx62wHAekfEURHwkJ3Ib4bfAb7Mp6YyUQ
sLJgqaS6plJsfj7eK7uCLl47suUlMlA7dPNXnA4lMR20KG00ew/ZotW2Tv7iK0ZrI6IeyUO9JnVU
9qatDJWWW0t1VJgoLYLX5xjShBAvLvfPy7fCmuhJzNPV5klTu5bjWnr8LqXyezh6MZd42W1R+WP1
iBtEiSciXBvMm0DFuStLT1SPtuSgXbbxexUtvfmAl6NFmG3GrSq5HPRmaqkeJ/WEKmuAjdWNmo5V
ZRCAARc9ADHp6zvUgf/zF9p56JPhWUd1TsKDo4hqFCTRySlZIkyevuWYBZDhzU1Y+YCqou207a1O
HDhs6STEF2EkOjkOgIVUF0DXY3mNx873bbjRCA8oYVdizOFH/F1A5Tx2DrmHo61Wal/dupif1+Ya
lyiJD+8VTJ1IhMdmX7yfsqXgapQlJK0elm9kHJyXCiqGfFrD4wsAsqWzpW2pjKDPzhdWXVQxjMDQ
9AZGbGJsscreZvxhSuRLRw7uBOzSGU8tdf3zxGJjd1xEKzANiO0HSn52gWaiGDwb33PI7b2tJZ8a
3Yw6nMVW5LOQ99LZpG7R6xo2F1I7jGObx9o+pDB9LBoOZgmC61k/aawLBmXpcqA4J5lwzvEJqI52
MgItpbgNiy11EfeGyO/M3irDz5+AMHLQ2vhc0GkNTArDU5HNz5b0ZKIyfhOn8BXOh9tdXoj5J91g
wQ4M4oBEsafwju69X07DZsxlCuuENA7NG+SgclykNTGIO95MDz5sMF1oJ29q77Y22tejyyjE8pI1
9hC4YPeqmuuhbjh0thUQqgy3GnbGYw9TkmvdBvo3KvNZXuaEfwC4l37RZydIuZ6LgB8bME+wl90p
ISxQ3RkfFveDU2mGMZjkxA88iJJHKZlPT5T6dIL0D87ZCwGKictYJRSiP006OaT5fbuestO1cWvb
OeD6zZX4WqZr2Zt2SAWGA3/fn1dxIuwIKlovPOBeMwTzZxnyBSSRJMQ6S0irkTuXEJHAT59aC7F3
vwCWX485KB+U2eGgReXkxStXs5km8Q6FXMD0O3q/z3NdxZ3HpYb4VmOQj5CkU9/42mxWT/oPY0sB
zuwZLE70I37xMduHC8EqsOHOR+F1MORXaqfzV8XAHKleZUxgGdKmQ6QqLF5/A2SCVCXR+PUH6b5A
KRq2IQN7j0CLZLzfQWt+pWAshjISM98nrrIsAjUZWPF/PNAOQCrHQ6U8XXQyE22unpFQHRWuq3Fa
e/WDt4i4BLALz2lwAPdbZjrUSL3mWsMUh07QXW2ehxCAHCvfpPAmK+s9rZhcvmO0/f9z01HZ58yZ
3n81ACZQf4+p73Hc4M7i1JOcYMryBnRR2Pa3wWl8ImZPYAqi9+1qR1au9nhjj8bW11CQhtuHeQg0
YN6jv7tyRpOSXn0W9lmoNQQr1e1LjBzh6h+Qqq1w0vz0UTbK1y/rAtNrVmILo1D06xF6Spc2AU1g
ONlA4G3bM8ixRS2GUkbuBHMVmGrJ8n6EheG1GfR17I1vBpWl+zCDNUEPBP6pMksEtYhuEU90A3E3
j0QzPvnxu7Y/ob6sJYa50OTa31bvEv2fcg6KXFl+4+HtCQr70x5iPTK00L4oPb5dbnzSY4XZVeJN
oKUs/Bpn4nmxjnHdwNsXDIia387m9Lo47xa4kLgoA605FMcPoX+7Yl5m995OEDfKfZUnzWpeAIYh
reiUOE+VjtHGYSlvAN60YmfN2+oLCcbpYRhOs0m9gOQHUMyAIh6sybpmD7hxgVbHROlY1obJQo7E
ENA27aJzLMosinP6qmu0s3IQ8w0BYmwxEdEzA5DXCKY3VUkScVmEA/5ptitpfbxHprq097hK5WrX
06n+zBOIMR4Eq1duvy5YldswMAti6F15p0fZKZozvEM1ijrI1SZD3/Tj9tGP9OePeX4iRtkU8m50
9T2y/TaaPl9r9W5Do0yNhCdV9r7141VlahTRA1YPhSJ2+b6wIbbvRANcJeGzsJwhuUDwLuCo3pQM
q9+PNcsUGifrKCaA4OH9Cjs2u1QbVKMz4RO6JIiyLyTo3F7E9P7ykfitPjLMT7z48VDG2MYr+FzQ
OxkajUXsZW4/lfS5WkkZdIyrvxbPtFNoQ80TydtJT352XE4BUQcjaHJg19W14m73928SjWFETy54
DK+VM/HBjuJjUJtkmUMAd/8k2C0I9QoizjipiLzkHNSo/gze9M99aOgyFXFCgLgjlI7dE33mWoi3
pZRzIscqgdctA9bbHDujRAUPlewiThJjsQha9VzuW79KsnxKo+7pj6SlUtiJ/VSFYwux/aOCOpip
AUprw6nLMIWrlAOGr5r4r32kjT7LbQ5zjqu9lBri3m2+89s8BWfCnXcUf1Qn2xvr2rRsnCXxbD7n
mtqp5pRo81lgb1Kw/TdNDzqbOtkxcgVO+t+u1e7OvPITvDNz+kJHhrsA24gZfWn45KCK2aLSDboh
Uq2ndajFc6LfkLmh2r0AVm1RLdAMsYQwVQW1QjAWcZCY+YwbJCXISOlMy55MGgr/CD+kmPayLYEK
c+SOWWXPOzV5i7BjOzMlzsEQLdV6ZVfJQrGMg2m8gTU6xdeb3nehrpMr3HQhsKWFYYKGAh8pnPWt
IXEORu/ft7b3RXYWIj/vHjRA7aiOnVTgtCpxT8G2qICMCtz05BuXjSGB991MqMQF5cJp6MlOH7n+
bocHLQ1Nq3ZjAj4TWfOZTvq81giCtZrdMXAS+3X/64ROKbMZn9ShfxGlraE0vnOLwQVaEh2A1OId
CcJo9vRNE1/dQwPNB5UzldgnYii4/Yq6QnXI3nMHFao77BcWDpNrefdXw8wztTkn+NdmxU6lPLB4
bpf2uVtN9KGXRHBNbymcVWGhnsjEss9U9hYGkpD3ryqyq447ejbdbZOigM3yvIS5NKFOCiu1ZJ2P
CfP2QnF2UrvUzz8dsKyg//3DLkiSZLckJ888D1QFpv9O4p1qswODZbV9j6+uKvODJlBuktWA/Du6
fFuqJYcOnFtZC587J/aHFJNiBd1Qs8jWu4S3Pk+sc2OLKoiLlEoU3oAjDrymVSfo1/3LLP2K6FVA
poRoIb7vuQx/LyYnrzfZ5GWpxxaA03dYXxY8HFn48Kug5oyrNKU0D4vARYtJdnwvVKYwaf4Jdw3C
pT29Oy7ysfhHfwXoRGUAnp0DWpAUcE2D3vK4hMga6sMkuiv3troCjzI/j6zcY8k7rNn7YozdDhBn
lc68ZTa3nX7b82mxmyG/pWep2d978BYkhg9LdY7LbEf6RLtV6ww1VrsFDY/PZs4usL9PvWoBiM8Z
pU344EVsV9H0Jb8DLxGo9LD+hjxnyXNUKe9favUlw6Lj8+03osj7/bz7IBgBYK02wAWbSiHZOJjb
+I8SOK5bMHDReK8bobHK7OdZN9FTKukYuAKT/QsG6Ys175fDy74mMdOxE22c3wxNI2+q7KdBhERt
cY0nJah82Ag2RHF8iNl3zOvj/YuaHrrZ0oNwzlzq8tb+UVLSWrylHRM45vmpxkqg2ywYfs/CV3Nf
8Rp+48DlQS+sqPECiep46/tJdy2ZKCraC6NeV0J2H/aA3t9lP/jgoFopMafNUNWBVHK62g4m3bAx
cutQm/C4dRUNHwRkhnx5HBh6S4FlbvJ5eX6jS8XqXiDyxjAblZyZ2WygNY+RHE4jAgNFWv9QdUz4
Wc45ZZoAOJn4nEDrLq2lyz1/yE12HmpjSeLnnBdeK3ebmeLEeP/SJV1Tt79xMIMk2EOHwrxTw/ew
yIBklhF4zVu/6KbOOBh35w5EiCHBapaTtQZri6tNlVG6JrFwXF6UvpxZmf/LEFFpFw48N1cOUQXJ
S06sb0gJ5tOwuWCeQNj8z9o0Q/RjgevmYfy4544xGV1jU+ypm8SiEVRq3IaanUwFoMcpN4Wq5xoV
MXwW+BFevNkZOZqbYiJ+YCZUHUfvFNZE8eq84I5kqK6fh1SH2UIvsYt2nnpZwUPYFRfwz8PWYoyC
+znT2te30l2sZkZd7CFdvkKcAIloEeJlUtbw8cSW1Rg2DGVYf3yEAjxuznys1Mu55sikGCCILmOo
QUYL6ZiBXOKU92kMcQ104iZjPQO0GJ9qi9zPmP1BSp1HY6DRjoP3lyaabFm8JYe4xtObyS7BrBxw
EZX30CtmShGTC820tnyUpUuXfGRv/QbNExIxxEjAM1/ViPbU1kThx6d5Iqs8qtiRkKy9Hb9YLZzH
PV4+yRq+syIDcw5wlQc82SInhL0jkblLEm4IFOJDFntjjCcqkzVGcbA8pSyioK3TTAkk9ajiVluJ
8cbmb5jJU1/vUM1nTsAtSoQ9oOWSvqG9A+pfYfED5Tzs2sTEKJoG+g/U7XCOsZe4GEu7DsgJSEh/
eHLo2zcFn67hepPiUmTTbSCDPc0Bax8UVzWRVwl7kDz67u6maAFeLrBFT9d+7vGZJZLZP2nbTNYY
3jXkyr9xO3Jzc/JozDXUrkUk8Rn01ZdzuI23KBkPpzv4CFh8c1SoQinl+RRRPK5GoWzy3POQ/4jp
JX7hsXBYeZAtIRVCa448T84dGEkWF9P6qdAaYuKqHVNi0JF1/2d8xWtbDwpnBiA/NKWYns1GykCe
veW+Qtd0RNOc5+9wixtOsZwenuCclcgsqIwatjncKdbs/BI/s/qh85a1q8Iwtekide41PAvt4o/+
km4K56ZicMpApkLpYFhINmNCdmoklzed5tOLRv2CYuFRPS2c8id3y+/FrQFM9l64DDTLQUYQr2sQ
GkKh/kQfjcgNcDUG3k3O80Bobj9/cERqF7yVjZYHdZSF/yR7RW9JI83pAAiwYAAn46kAEhEyuhzQ
Q4dZta4erp7zWjd9gqXurr4ZnJteEgRzGH0AIPmdPN1O3tyDhNjJVQ6Kumod1XqETLUrvnfyQp30
xyqfhSZCInl7cmUGIIjzISP+HexV6/4jknlBwYZiU/68NsMjxuNqGrZPEZihG2/bRuywvdcwaRaf
a3TuPMvwAQQXpRLfolbxNbgs1OLZvId3iStv82boOt+4FM95ZAi+d9I5Reht/Zdl0hyWG27voDe8
dDhuGNFvFFn6xZgjbdB3w4DGvc/gF0zLYwfGNpL3vp8N/wVnns57uEj+S+AdqzzPVw3ZTGLuQRkF
y5zdCNBeEKm6U92lS2lQmPfaQdaTK3rpfXCDzGyRiNPFWV+GE3l6h6A4jBW95gIGh3bhT/Yqx+IV
U5+Pf9izLVyXDKh+mK0A2LCRJww247gu4wZjKSKetSjGFBKGQ4k3xnuNbVn5vu5QkXvorxgqezzB
lCUr4F/PUWCb1CA8Ms8DQl7OQAcG95onOTvlzc0YXml/PSWXfv1TLOg81KcQyulLUUcR4QQBrZBQ
LOLC7hY2hCF/LCPSKhx0VyILQCbjSXn8/70a5TZkE6eGj7LwcvERgeCa0pUQqRBQVx13GLo2TNrf
iBFDEiRtxmzHnhWBwP4uiLaa7kJavzVZ6JZB2qsxtOW5GOig3chluqEkwGYCVeo2aRCAHQ9qyxV4
FgMn53HR2cKqEa3d+tVLDuLYUcX+03tN/T1o9H4Xdl7veL6VRMwPmYHCtAPzDl1zGeHMAxDXp8/i
y3y0LhYPZRJatWC5MxAZuUnLCyPyNETVr5JCG3cC2fUaOgzl9mddYWzZa1PPa+iPr6CQxFUeqdGr
kuHpFr7VCW6QfiBx9A3NKo/iKilTKgqeUJQaauEymRzyvGEjrfuGF+tsLSl/vnKOmPdCxJnXHFOl
4KVX3+yhzH+ZdOEyW1UivNIkzZuhpFbVyaYqyNqYyBd8pEvVPT4GBfcG1ohS9eERpn406evpoPbF
Actr6YnVyQVeeA/pgUCyv7ytkwcRmQXggvvGGhg5x+5tUbvgVHx3YZyiNFDEeUtRGMwj2ocMMKbu
KHbJBwyxq5Ob8OCbXhGecwGswW2XbbTBe59Oo/1Q1YzOsXHLEn30+eCsAamFGNzF5lyFg4kmGbAU
VjPp5fsZl0ujlY5qYtSj8K33FUFVyHVhKhsN3WsGTcBQsvTG5t8vx+zB/q0Nl3/952C6WM/x5zSe
1MEErs/WY3gcnEx6q0z1ZtKmo2vXoR0b/e9HsYd7H9rgbuN/OB2Rtcu7NYg5IcpDiJaTWCDr9Byz
sUS4hixsk0HZHRbzFDJhfBC2HUSJi+moDZYw7YZLlay+3xqAtmMQwJZUrRbUdkb6e7O4bh9cxJ4E
lCiXpHcn8ET+AD5hm2beWk8loLeNkYo05caGAGPIz1hLzP+mE9y6D6oVw1RZKRYVod/mZF4koCW0
05elSOvhfSlW/Oh5no1o0ZzRkThFnxBDhSs+DOXki2mY56jlDMjV1bL3iVFflDfMBPRquOnEfl3d
5gu55jNK2fMdS2pt5bsGNkCNNhPs5w69s+kvPWZCDSmygMxYOAHuAFvJYYE9TcXAydyhrtUFeFyC
xKQ/Ayx5d1JcOC0lFOuCbPyaJc2gzqLHprk/sAbHngBfyu8dFaRVZ1n0Uk0wsaCMkHant0cmAblg
e4WrFOGDOKgBdaRzvDM4eb7UA2F6sSesqCgAWoPgbq42rPWGW3+m+KflroDLwKoYB8CsYRbjzeg9
VpCDSIKZkKk4Jaf59Yxv4gSvXlX4nGcEwruvIvtROCoUBPBfkC/SOHciyWNsuYu6+wOJlrMYTf/n
HL/CasTx//xWkmMGLAjVG68Ma88iDmIXBPtCt/URnWaOeKZUePXtyXqm96B1qCIh6V5HPGpE8ANF
0+6APu1sqh2jRTgoCEwQhNgGbGJZNJk2id0faBxYlHxli3O4F5xJvRdjFzzrPXVlOTQ4NitfTj4U
2iFY2j01ypBaYhwYKYC76WrmI61zksrLsKronQWvILpSnX9xoX0BblYjegZydLlcOYI6/ruDI266
WRnHVSJPsVTvrR5j23j9Dcs3n4PqKNMyfo14S6gEBZcLujNaAOD320HmzPnZXnV/abM/9cq5UI3G
EgpitBl/An9Wo60i0/dJ59tJXWyG7dhRLALALPp9sO59RA1iUR0uPJCTruUm95vZ6r+C9npCCOAs
ShGI7PtxK9KEc627qZ6+eqtfz3s4ulHEdeC5CRBRhZHgBtPbbMjMkGaPa9ZLrahE34zjiieunURo
GOVzTzZ/ouTeVcBNwz9C7GMYZjx0yfrd0TY4CNiOY5/DOmEcYz4SOkVTQQ0d/khFPwhoAp2ZgJkP
0PpCrSGqg7CBozD1rw21P91xo8Ap/AHd8RzgRIvJeVUz2NKC0M3pSniUFkFjj6lJkkne1MIU9gd/
FtR70CwjIAFGYo0rjMFgOzToMhmmCW1r73S3kqqxBDZKE3xpH/pzD/ZOW1KeZHST023kwnZoJH3H
3nQ3XWUq0mE63lHEpz9c3UgZ9tq3oI5z0w4E++iU+EiI/HTo53RwaELpjQ2xhqOnhiVz3M3ZLgYe
kn/i9J23CIajCquKDLhNBv/0Z4ipOe47dDqVx3+CLMC5iCd6t90cYSdPCIyaLTtfI3eOP/QnK/Ez
EAu8ECT5gERZ6U69B9+GXKZUcMqnH3bTgTjqevSjFltlSA3VH64lCN+TlSagDjjPPobY5YkHcOi9
7IZbsa+7RIdlZkWki6ZJji++2Uwmzk3EGZu54KR3R4oj+7cULKpbEfN0oy6t2rC9/0sdWyWmJaKu
/NKnaLH8Y7oz3azotZAEvTMnAi3sg0Bn98sS0ID92ugWu33ax04aUWemjftfaNduu6v3ylT5tuK5
xCGrR7oXOPuJ/1yPJi+a2RlLCd/UlT4X4ig4UgcFjQev4n4NmvC4Xs0ZxX7P0rZruadkAIQ+0I4N
N4tDV0mYDvFItGgCKcCNEv3etzUw5t7f1K/AtiiUwmODJebWRfJTUDLAAXM2Y8cF0p0wZ5EDyPq9
ynrIPmOZ8E737CAkY/WM6EKsfqHQx5AkUVpUfR+Kovr/myjoAf+7CcHaxK89seEXRspkIuPc6tVq
kaL546JfFC4GLCpfyyjq+/EDvj1Ez04GqovQjS4Iq6sjaT3u3V6Tg/3uDPW6ZDgOeqgSvqWeZPZg
GmfPoZ0ZMHgCIpsKrGgN6wPpCoKEhFLSWCQRZ3Az387Azmx44fALrWbHSmE7Okor366RkSWInEeY
q+oQ2weLlqJ63mJQuKHX1wv0bGpzfVCTVNSMtLOl+RhaicFQQAkkZHtVadXjMyqi8tFgMW2X8X8U
b4rHUB3QJHW28MbFsX7xf7nUXinAA0N7Ojgl44A5xvahSHEakpZnVkSkIrtduLGqlzfvzFgC8FYA
AFQ2vsvJ+ZQOy49sEA1FePBwt8uBK3gNvoGNW/KWbugn2YJfeZerAThC5uC/UMTG3I/r0/ka3gq5
0yHY2xav9+2fdHFPg6K0LU1WPMM7Y0nuEK6GhAEiiYy1rnIqfydmVJOL8KIvBfn8rq7c97maUKIt
YZD4Ur4bEbH5fE4IcI1wbNb4BWVmvFJVr9hzCboELDNdmrKAZ8M7fj0giglMXP4hzXTQ0PtTw88L
NhCQVSN917n6Qri0tsTDRq9RqoN8VJTHuuB0n00bgKGnIwhB0vLcfiudMsHTGBfGjYTAtsdnqVRi
1hB5q2zo244KEgN4QlQZzP5E0WHU2ryMFADRffTaRJ6P+Dq7otj19haaDU3F3jrbHT3K8vAAcIC7
r7JZLJ4H7c2hh8aCDiEx4vxT9T5lugz3cKiOGM4Uy6674uzxCk/SY60yzin+GcICQFFdHv2AvUgz
K7hBfYFghioE0kZs11i7mSly8qkeZa4XPgoAZ5MjMTmtsSUx5z7X+906GWCPCkL5qF7T+oUgWhx3
gH5KPBeFwxx9r/k25mhPVZ07wQ5PYwm851LrevDKHraJmnqKLJNqBtzELIu9a5yrv/JORnepskD8
su1Vlpsgxwkn+SrdYFgGypnjcPF0ojJdb383OpHl3wkzSJjScvJ0yBuMh+FL24ySkQoTtFIrk5T4
2qJQ907TO4DAxl5kWYwjmv0amNtYOp+t3VqUK7lOiizRWuOrEzd4JGP5M/QNDBPrV7csenJjbsbc
eCGjP3lb5o5jJgOpvDRE0+EZeT8WuwtWo4rK9HnTQtsnJuf04rxBy9K/Pa4uGEgRDDTWLm09WwOd
JYRxXEg3Vm24mYBX4lmDM9pxzMlCpa7fu/D6/RFX6lzLqZSL2b52HkJMm3eSiDh55Rnb32PHsBsV
SbHh04W5f3OwubmuBidXRnNUlT9nmL0Dss9TZtO0MoNMckq17qK9m2bTuYq6IxV6X94uyuFUORGq
90nAKp4MyLmYavc+LMu7LXwp3TWIp9nITP1pi2l9hkmeiMDACgGMD1yqJoVECj1m0g2OmkBAax+g
xDg5amX36EOLYAvzPFd44TCldiTNCO/F6XcsU25E6VSH1XfB4AjOcq3RXtk9lVcWdr7O8goWHrMc
e+LCG5g0LchW1rqVde+Z3KAO/90eT2UyKENW+CCq/whgE5mUGdtq+okreKnC0EYDrh4LPNP3fedC
kjoTfzO1LyUfwlllfBJwpT5sk7JOm4LZEEd1+EuAe8kz1xyLymrFSRvxJcv0zZl1nu8LZXKVc6bd
+VpQeFXiKxn8gJeLOIJa+T4AIwWYByo1RXKdcO5WLhu+fRVU+eA7m6L2j/pXx4jtRWutZ2Dtk194
fYC2qiFxL0UrGpFBPij2w2oILnJBsYiwy9VHGqMvbuERb1rAmj5wpzvH8uRCOYrf7GNDjdB+8jv8
dMCfqDufg8oU58FVuUX9m7N/CBHTTvylxFlYGIH0p4O11aYE994GHY3o4+pTqw6JXRNmJtkHMgwF
I1gWqEepSE2R3KbYYtDoa059LLWwWRIRRR9BzMD+txQyJ6eoQZPqBWaAUTHHycCO7MtYqr11s8sw
2OjW43EZKwU30nYqtLSquaf+0ID3yLkS7FW2GmqQr3fZGLC208iMPNEdNJ59NwLNOXASEQofhC9c
vznZb6mGO9KdjT5wa0n2ShrZVQdEYS4y5K6dtdkfTulKkwzEoNaPGlYCvptFQoObwSyKbDq6Pydk
wsnX4mAjkdf4ZcOk37RitCsuHCIUvWTAvwZd+ZDZXEqeAnzyu7rIe8UfZDK1jg1YpzveTp2XjgdP
P6a38S/2dOVckAL0iK6ibcetFt0danBCTbrpPme6zZT0VWAeFhnw7UQ7Qo4VrapuDZq7gIQ0+1/Y
uWVaudV2n5ZvD3RMesJ4AUyXzB5oN7bc/zqPWXFZzO5tj3d/7v0Y4r1Y6dt5I9075AdTKCmPwjcd
Wyj+XnOOtD6ekcCBOEoYi4PSvaWZ8lKqZEDIGaXtmHyzrYRabS2r2uCXpP2Bj2TwOMdFoVI1/FdC
C5694gorpOlj1UBqXST/5ya2C3hqR5NEvrNdgkffqIssG6CD2WA28MEsFp90nefSyMrmldMFpTfI
OMIBklVSqN5W/5Y1gMgPsky6rT8cFFzX3wXhLnCeKgn0zpD4nv71CptVWDzwCqo5eHPl4InZ/Uj/
LkJB5kRfwXV33mMPpPYbjWIW6Ljy3kGzJ9oblw1/6OJ9+AgdWmMVoLmE/hrhGNUw/MOQY2H+W/oj
YlDS6HWvJ4Mb5/xpQuUPD4kJK3WgrBBpWAGdqVNxmqbyFvjsThg5reAVzrUTUpwaI6BfYOCRQ9w2
r2V78QMXzuEAWAOiJVderiEWat9fTrcBLk/QgAsHqrlVQF9M5yqhMH+++GBUMFC2qVho0/y6h61F
W4rI/8zgQmWTcPZwdQbkalbBQj/bGKy9DmZzPHJ5jfOGUJnXfBsW+cSgZY2AyeegZmWkWYTZUjHS
hCPDSRzzWgfT/V75B2YcCkasCwDHQYv+wdVHV49FTzJ9MuiHFWH5zgNzgUSLXjxlIyG9M+3MZQEp
gLEaCbjFNrz52qsWbEnYNn5Q2rNj+5U+vjecOVKx7bL64vJMRrRj6BZj6DsY0dv5WpruDVhx9FTx
NWPUZ/dMPMhUObB6/YZMSJISmuIxhTNS6Fe6pEk0hdtTHmK9dqBoGqpSQWHYNJRUjA5V3j0Y7y29
7KMexqAU0Bo2F7D0O8MJqyFNB03GLY+50HBbHwIoSvqZs72F1TIpKT8Be4Turf4ueKuxLbkjhje/
ASpW2Z4vFShQTdXmAqpUOacIcV7A0ZKiUrX7TNXdjkoGXa/pvlrK+3Ysb7HM5zItvH/7vTL+zMbq
pLtVHVohG7XOelt6UGBFX3lwf7U7kX9ftWOq2LLItpiiIVvm2QjZmQ75/MoSZSzrwtztjpBI7wtJ
rxfGXL+5YAk/IypRIWSzycGPEXbeT7FTMCPj/O3fLSGsZsreCg8jsoY6QFBbQUkS1RiiGLDDtXtJ
7swpRpyuVoT8xSxkPdV8utuenzQrcTqrPbyrVMwJLM2jOUkgUxGLcy3R9m+QIztoKql34Od2NQ0H
43oP1JkqWO6CjWaJ7vVaQpLKzaxD6h2Jaivpe1qt9lOlbRpCs25jePVi8CsXG6HHhXvtIpY7oNlg
1RE/TxG/A0T/TxZUZJRygMke/Q0XbloIGqbGnU1YYOdtQBPotX86T+owo1P+8AoWGklkSD5fHIlo
Wa/cuGyLlcEcN3phhyHEQUu6nFID7EOBGQrxXNI87tzsTcEOgLQDvuCWSIgMZ64spYIV7d1nJkyu
BcltXHEa28F3joaNzglD0kb7fjlVwjLvxmi+BXTjps4GWOki34TzCypmLrqLRN/jUxI8Rl0PqOYl
h/vbCR3cV3PNy4rkqKM9yhQiGDu+Bxjh2fou1eMdP2jjH3g8Q5n59NfNdryYAQRxgOc5TeRJ8+JX
FYBI5JScU8Fl7aGBTo/DMuCScWEEY3LT0WJv2/SOfnEkVaRU0I0VGP6/JoysUDU6ajec87Zf/KtD
15vK8k1raEUEP0JQaoR0D6vmnn9QXU9jokm8xjmJZxAYwLI8+infG9QBwCkHTfI4o9E7YPo5VygP
NjO2WjbD2PlRMJE9Suvs6p8ddqi/KkW1x1z/1jZHO/lYg1IuznZnGbeAufdVKEZOKrEBWcnmPPq4
sa3ubjCgjmz0a49MO2TnYRP88GgsNGtKaC9Hvk47Lk2uNVLorRYOi4OdN3I0EYnNqqals66YKB1x
cTLZWhi1BoDE2Cd4Owe+pimX6OK5IfSHwz/Uv6VUY40YO96VOFwBNyW1vx94fAm64JyQc/IMC9fT
V9NHQQghN7csy0kJzJVkYsXwwb9XMS9NQTpR5xdNGIgkkltMstRcdGn5OERz7/dRGtUF3RXite0P
QhVhwjp90wTNM+4DKcUxMjEx/bcehJmQnh3SDX0BgBBpgtLSoJXPm8Vb274L1PLjQXq0y2tA6E+V
jxBf3B2jxXSyIy1Ej/JBcb7LDvqvHS0YiTklCgCp47UiDU1Pao/IUq3RaKIBO4Qbcz8YfA+7xasw
lS3UKGukFGcnuwTq1Yh3jWYcKZeFSc+Xx5lizLh2oADunCOupr9bGd6Gd0VnNnVmTCPNRx3F6CvT
ySAcg3mz90O+fzH7IWR7OdEjyIJjh5nk93B5hNK2ftHsJJ0QYC4PHG/hnJ3znZbvfjtDyJq5Aui9
gqjC5VZJ1bOS5/YU0LerYXeoXVpoVBSRK4jXs1ikEhLyFFkNIPzFSWXBoW1ttDQSY4PYjeoKbq6X
wjbRqcIfoXPQYWok1AEiR42TnYEpz3LCgfgFEeCs9hTnQeK5+yTh9V95BrzxD/KZS4mgtd4iTqCl
ElF+s2PpupWl5amSLXsQqq6zdE0i0N7a439ZtmdT+ghbS71F+sT0+Cf7ZVFaoQzjSGvy3GaAzfhw
EdVnMdVMjeLrOdJQvGLHEqQE+WONfBhakt2ZRnzpAFnqAqsYLHNs7FD3TdsLQO65tbOSPgufp3pR
glb0FemNXD5dTUsw8GHQA/bM913N5bvJgrfgUA0cxwi4sFyBpQ2BkYvlTvDpT44IVX4UDfTs62g0
hwJVLPf2q1KnVX/gvfjDL0iETUaNQnQUXFOQM+sc9ZijxTNvgTrWhx7eRpTKJA5/1Tkx9jSFq/S5
9Hp5ka45PCbflUAJs9GcYAPJ/LB5EOqW5/qbxguhwUQ/JjkwmznhyKfmV6sb5f0n+MIA3s23+5I6
tk5V8KV+pNRGbCHP7fD9MObmXf5ki7qKzB8Wd4OaZZA8H+8qLKJVGArmujOIrAKJkxXfPGJBsXEm
BC+/bsMthbpLpP53fIUerzlghbnMpQLGxp5kQfvvZ8SdVj1o7L3wHB4niVzpe0iJOvq44vCikOL8
bBu5WhmR82wJXt21Y1fJsaGT+MMs+8FGsq1okoKrVCyBmNQ1U58GHQCX+XsNhUTMdBOOwQ7lG6uf
+9G+Qh7GUFIRoquH+QrUYrHm4OA1wZtau8tjxuq3xv/w9E0PwRe+WIFupvEcR5Zwz7vYp0ZxhH5z
aGKJuPc9s1VjVzfrrxx5oUq8vSdWHmjEKGQrAJImDWBWG131sTEeeIWBOZTHbW3IeyXANfyjswHn
ZOeXhyjXamrtUuklMyXZekX65l8Z6lrl7Teb+YIl+oRwHXoHaffnQhcz4bV3rC5IFEQIOk1TJTGW
EAOXcy8MY2o0uHto34MRDfw7uNL47r/z6FvfbITPg7kI+Y5H2WYn2Hob1OQxevi2tX4VdtLUxcGS
IYtd+xCJKRAdh53lqz4qUOrIF5zwKefVPL1/W7yn5bH5opec0eh+BLdGRiFK4zLaLrXtMIB2ZXXs
FiwLhxlpiYLNEGASwVDu5kVUXsFPgAytjWbwoducJjxeBrK1HHGoTGnaKsXq90WkfwgJ+Rl5qUaf
0uyYYXCfxq0XDFENOWwD5LKQpci7iesqTMzuPHB6+JTmhtCqsF7P2MS/fK7+CYUS5PjSorVOeSKm
v/RZjWBa02OjL9vvz5kvE4/dATyO0FJTSImN2fZWClYeAQeQ1i6Ox6p0qb6qOsB9IssVjgKLBigU
wCuIK7MBk3ipdn+p73Am1iU6BNl1WJgNQ55VgU1Ise1NAbWpseYj3FDVlSj6OFE+gtfIuaAJe/GY
WU3ULAVlUDX0TrePUd/u1iJMSskIG1jP1qV3DYV5lCa/aTjYVyRTOmdk+/PqCs28uW9q12GU4Esv
d/3jZlhZ4nEuE85zl+bETGZfRJbfJH6+1Uj1qnG1Ris1ka2uwZotzLpvjjTljbIv8WoZTEv2mziN
EXvurQb+5veJUN3BUGklRe5secM4sH0Yice0MxisrvicHiDWD5gW3UwQjMLUEx9e1uTeV/WWtDwm
8ZZZOGj271PEj0F0JDhtqsfA8LJm1mlIHzaD8r8Vo1AEak+7gBT4ba1Jky+rfjcaiFA1ZttNJqNb
6tSIsGzb5WE4j9cOJRzmzTcNDblNS5CCD724AlxhzWoRg/deSJ6xcuharASM+nbRduzuLj34CGBa
vai9s88JAI5QkMiFtG9l0JuGOD1Tm5HTaO+Md/mSPwKt6pj/O/cT2X7exWxkxTFYyKxf3UKi/9Nz
TQ603WCPOla2DDlPcEC7wuOs8VPq/rcDPA6gvzY5eoH0yXmEZ9y1Rvt4AaG8+pvSo4H1orihf8ng
DhdTlK9TdKlMHiWJEOfOP9IZu9m0jzGhWh64qS2CKNHzH5LbDT6/X7fjigdDuon1iGXkmO6Whfg9
BmUIfh+pX8ESEQGUa71NU35KV538G1Z6TNAxmPbB3ifJMBFwWEK9qM1ZO0lnpjjTOeCBicaak9Lm
OpQPt1eDk4J4v0PR0PF3UhsbCXf2HbY1kBuj6MLzWy3ATc7/u0cDl6U0OFY7IHsC+hocjePWY97X
ES+SGJxI5kN6cQEpsQR3GRYpkJG2Shc0vpKUgBwnZ3Er+2H1HbVrshOHsKzChQ7CKb2CwEpnhVpZ
6W08CHeo57Xde5R8LuszuX0md8uQ2MhOF1xg1+JWWHnIl7bkbQXqYVyAhPs8rlmjDMMEYc4/Umb0
2FsTYnhbrS824I/igQD9qY1MBMzx1feE+gXUKAQftyzx4OTM59stZ8oQ8MDYunb2ynWQhMui/qxC
PKfzx0EdJlpm1uRcFwdgKCDFZEmwpZ5K8wJXN/JLNF1IZhRaDhaQKq5E+QjFbcaL7bXbYYjWUzzY
SxFcoMPM71ZwOK7qn4SSfZm5fyy6XcKTnKCy8k1r6FvZbgxAxanBxTtIElACp8vL9U0x2QnBfhrw
qQl88e+d6o/Ad5zVSWfQqVwaBEGCSIzGHmdPoo0DpSa4N22onibim85XMlbSDtDBprkeIDg5/LV4
6DCWSUVSbAl8Eh6b+4zdFYE7XCRKoGNXavRJtH81dstxWWFRdDXN7125y1n+zRS0rKQJsDiXLvt7
xbPjSeR6G8194qjRhoBKOfrEXng8O/ApEKndp2ala57U8uzPjvkYiS6gawR89QxmMYd+Yh6keils
ZEhKS+Zp4Z/fbqAZkhE07qZvfXz/HeG+DyCYrsaafiAiVAU8519VNVWuun7f5EfUBiY9fwVr3e2g
2EpSbae5UaJIAmbGpEqvvFl5oMha3hWDOTsJpciCtPkrJ/qMbWEn0+8SlZR09s3gTO/QW/wJuHrh
HuZ+lo+IkDrmYjDzERgQhPn5X0nzM3jxLrfJbKVx+KFnMlKyVoIqWyAqsdypRp91iRjr3+SSvKsc
k0dayiDqJ11Wti4V1TA26odOSsy1qbQKnZZXUUn9y4roCRrekrMRgZ/PaQI7QIRiwsWeMYVZIh3d
lVgSnKAPkKKf3yM8b7Y+q0gJM0K+0I3sx0TVZTs5ajrXJhDkYHa5eliNd1sdt/mPaAY4eYSeDSlS
Q2GQarixtgm5ztYF2qQ+iJipBQJtrqVV7IYemN05yvw0yetBdTVmVKyW+R335yiqbjYdpgdGj6Ru
Js74X+hGccuc8v5bOqPJmBO8v/tUrH6dXvQKe2EloeIfwMrnrbQA0YojWg246xYG/SeBNqkWfZna
0k4LBKUEFNNKxX4VKzpWKmYRo+HiBGUWwO9iBehhED0wji9RHUcYCOuV9loNev0vPqUFUXRU4+eW
38Sh4C8Y+cEFuySYbLuOnd9Y+ol5tRm+HrPnJ+QugH/naUDRaxYbwUXeq2aYhHuWSIfN5T6+yjqH
fyAAEPbOEBoYApw8ZS0j7YH1BKxQqusd7LNx1jL8yYqw/GWQi4BzIyLcaxV8ray0nopkxD2HfKb1
dIb88NRPOMilWR7wrYpsfrTcxvRUw42zNTQOiWFBNOZboWcV/7sDePOFIWBa7vThYxLc/49putfq
IGhERAAa3Al+cE4GswSvbPlXfNNNDYD6ffpSj5/ApLwS3msey/qdqpOChy+pmphYt8dwTGkntRIX
fWKXC23xfyMZ3G/O0yn3G6VAXjhgshDTuAe55JJhUmun69rYqXCskGvmuhZXiQCRg/FYtpOorFo2
kbObez53ru23LZpM/4pMVyR9lNJPmq+No39Xc4s5aVQhuYQ3+O7I48OMZlbJwEb6hPBBNVkEkmDS
Ayi3KxFju+S0JzwwqMeKDTtCjuInmbOMhSxRtyUkSQSm4Pc1mJkBB6zgMro9W9VzC9lCzvhmXBtM
/aJT7Uqn99K1vJv5A7bw8ePXkijZ6KV6C6zADqdyR4H0gZEDZQ0GCA3wLCCcP/QkiD4sZeFc3xuC
hmkx9/T495Gwg+Kr5O/tfszHIcezi3moU7dl0ac8MRNiaWwgS5cFb/M8/RjdqgI21wt65g0r1g9A
xhW4xBtMF5TyLQzNVdPdYRz9gOuQP7+40zOBLriT0LTyUIYSW9uP1ng0/hF0GZJ73eeG9Zz4q3ef
OkYIVyG7MO/3Jep+ZHjUmNccKw3FDFdYuacaXjYkSGJxPv76aw/n7UNI52TcWrEM7NdspC2iw4vv
WY9Qr42Nq2ecE+eIVWTGRMBchYPkpNoiomWRzo2QY7OImAEqp9Rw0kgI6LA9iBznGptjQ3MXkXop
bV1ClvgL1v62OAtuY3ceIwo2k092YozuHLuS361OkpFrt1AdwQutP69ridQg/9acubwb/utAX0AO
0172sPMEn/CqvkbpRQ6va7mG1jeqsOrB5wtCSOJ3Onr89vhzvaHQdu/3xKOb5LRM5YHhJJNcVRp0
+HepOK1Q9x9gtyNzMlVPUyfNjHuFt/0GB7B2ac4HslMJxpVkUWa0DFYJOgn8W52LCYJj/VEGIx5q
T4RNIIjoR2zFMuaHPx50PtJc19W4zcVanQ25PBgCSYVoeZFPpoL+s4q4sb0JeRBXtf1TD2epZFWK
YkFchJ4uYeE5iZS3sVM9inQC5+4oCvnLBSKndOW6VJ97zIfZpCc3/eQLexfTHQn0jbuVL2hLFaRZ
0H1k3ExyJGbIQfvGhvOA07TpJ8utqPrB4JeH6s9a+vE9Tkam27D+/KPfDi2KaFGhzlKD37IIlnIc
qThBDnQcivhsWZTyWjG+V+ExMwAAURkxytA4V9PJQMeURjqVRPZU21GrvvsEfNxivyQI6wI+kS86
qyiQgZtxZ2NPN0OvfJg2gl1L8RzRJg9mZNWWmq5+DtSq30jXAWcktG8FzIHGWNGx/YpT7PXnSRTl
kzdx98nA+LS8c1qlCcb3XlSOZiGT2Ymk6cbA5I+PfWNYub2ukv/OTakz/DLGVKlhmeLtbBUz2ain
+59YA+iQlAxOZp2yYt9QggAc+e6HYnbVLFMbAenjVHtz3x49qkCGpixWTeTXqHKanuDOD3t6+1Kw
Ms0UsPqprI85jcyOWZsgjJsL1OXkd+yUjrjGUHwSQ9J2pm0vcsCWe//xxAYI+mH2akLONwT7dLeZ
FuIyudKu0Sioy6xMjQzzcRgUj6Y4v8QfvA8pSrvINnHQFNNN5u8pViz4ikLDPhAiI8o48g9Ak15P
YaFG2tlTjE/koZgbijm0w35JN+/7mqYgIx0wl4cHnnOID2BJstKEBlz8u11a6i8BbZpXK7kRIhgj
nfUIw8nzhBfTpT0eUgBEedDPR4ztLPF9/P4n7i2G0WkHmQoC9r0BiMYGHygzXYsFo/vQPCIyO1pK
B+X3Ou0smejmP5isLplW5QnRuTiq8ZJ5r14jArLJWjJwinOQJKwhoW9ky6Ko8/sXxMeHqCrmT/T6
JLfEQ1k/VcIuyO67NAwiW0Hfi7Na2/l2LqtRDdSPP0M7kaLXPMWmSK7k7waOUYTbC79mJoy/YFyV
dZaVvoRo0XmV/XoMPosKaWc4K7dQoduZ3svaGGNEIFKy+K8uyF8izU9bYABLrAdgCXTno2uGJz9A
ai+9MPhyBdUxyVbge/qNuQhMNutA7VL5y418/8mDUBRGysxprUJ5n/+TafK5Ha8fNrUcVrpZ7dmd
vgcHc6f/tXuZJJeoBVEHhcRuUiJBTuAj7q4Lkhpuce8O79HsDCJfsnYqpj9nRLoK+QRwflPkZu8N
ITe6U0tsMirfi6S/K53jvVpGkEt4ujq9i1Akb+cpbv6Fb6aJReHYaY6v9XMKQxGWtvpiJ7KwdBHk
Gox8VaUNxEO9dpm+Itd6XRweoy7R+ew4hMKt2vTgT2X059TTZEiUqVrgJY5evdEo1Fq7vo1pHaGv
9ca8gHqP8Vn3LJG2gc6fMaoqyiqEKp8x0WzcEE3hID9QT1vbZzrlJUcuJxRNA3T3clKJ09t3M4Gf
ujGJE1PCTaF+oCwN8EIqEE1qAKwNqNlIynDJ4bhj88jdGHRR78zmQVvMhWB4LeHmiOt6pfXRl5C0
xYTcH3l6EG8gFGl/cJ8PtqUF/pQZFqzp2A5c8cn0Y90eg713ynpGF1rNQtLDPyTHfpDFhIViUG+5
YP+I8vasvACqP8JC2hWMbxvi+lPsfRS8FCLHHeG2VnDdlFVahDTVf6J9H8agQcXozMOgdUvb3TdD
f+3wsRMxvuM2NnZwvr0uiwHbkvBimm15MP/hG6XOese4/wd5KFMFOw/dmc+lEYIDRSQLDqRnUk2k
30ssmEzZD6AjZSox8lvHpuu8HRO630suXI0VzdVwu+iAuc9Yp3wfFfMKfNWdRrjQLB3CLUuweLP6
MQ1qhLtqIIa4bmjKMXzY7iQ0DJkYHYekZXuom00R19HcqDtIWLh/EnuhoPEm0hvevlw4XBZMzmt3
u8S+Rta0wDUAyoEkuqRVrdGmvNvQFxk6N+mGBb4FOQR2sNmujOpnhnVxKjcWI9pEgdKlx7Oot9m/
/3IBYFQksHaj1xcrJHbIqAZ1tLa2873HK7xQbuozxP0rtky590t1ZauW9q7heG4FkKCzlXkMAfYY
fvEkrUrFOhbD29Vbfuvphm0060yCU7FUiQmYTLXaPERqic2SXFyU4+dnjzKhiuWTqYM/gy+dU8R7
mKaqRPOjJu9uXrusN4wJKqaPvGCdcPuqdABX0O2eE3U8tM4stQ+KGs+fD6Tn0vEVMkbzv4ONRwXs
EuzWf3Ij9dfqCopYfvaYFKuaacG31E5/uLdI9MyZ83RYdSZGAU6KRrBzY5giMR6Yu5Vrjsf3Rz1x
1utuQ2Qds0+LvdAuKUZ6m8yt92EJqVHNt/3JdUNCU4NxCB/0YWc02uPVBbi7L+IgrCcm6XR/2xGT
mwi7m7ZIH94Zi9q3Pl3wWxerTXSIkTDmlDUVQLXZF/z0uYVz6IhQp3BU/vEywd2YO2PMLPAkUdv5
NkgROsnNa6sgMQcXnWKoRZsG0VVw62PN9DqG4HDqu2qK1XWjD8Apku1FOgi34fhnBz51EZlKS7Cg
Te1Kyj/ri5OWFkaPCVoujnZn6A/zTSAcCdDqoS7L3Z0kQfghM7qwLK+Jr411Ml0SEj0m5h+RTdAU
qfsVz2WThfLL1tRQ9r3p0kPf+NCDVxN+D2u1hdKNW7yxAyI778SQ5xpxjUHuasTPi4oqw9oZWAHx
/AmzbmpQpA2fzZMmStFRJ7EaKhJZde/JRC+iFhGIft2iQhXuIXZJowqnKPbzo5W1eYUvLSg27JPZ
w5lQ6pF3sdvhMDBTsYZUaau21MMYjkRv5A0udRcCmgUk5WM/a5x8TzK409/tKW955ZpTps6H+myh
KkMbGPuKpWiMzTq5UvI1AcFuq7NGLd7DyXl9Yjc7hPcZW5p0NqBGvMGo+YeT8kV/z4JlmswUxy/N
KC8fnslL/MACtbpxSqml2/MNWd1z35eWD4oKAPP2xEc4OWsp5chNrviXsMf3c6eAQemR9wJUY1il
TaU6xvf0XGvNmbbk3bvhuIhV0L6gilIuuF74bY/KKH/3LW5zVF+P4ptCeRGKQIERSaax+kX2dt5U
JbmszVp97MVUmC4wX4XDJJSkWZm9dBuAIP4/qZlnzk1kIU8HAXCfbeqFCbM7SXwT0QTIzC7dZxWK
VWX5hM/Msb1CgK5kic9ZLBiY9P/qV+3n1yUPamZkMtQtsx4LRKpDGy69aC/MWdeJZCKj0Uz7gqBc
O3aB7fXwPcxISUxLY2hCihZyXZpYE6C/nxq5YzwWoJcGubGOH033HMAX2BimMG1QKBaCWpRol+66
aqKH97cbJv2hxoScHdafK6K5/tqNt7NOWc3QswELwZPmuwyio4qqccFOodkYmUJTeGZrmupOlKAB
JLFjyZGWMHZOLGlqI4K8qAAEZd9HW+08MMcF79l2jsCn17OligT9ImzvAkC+4lmuljEbFn8xVDpZ
uMEkeSUYK4fkQNJYF+MfzufS1YIcMzbVYYcsOCeszTlz3DahGS6EqAOfhDtcEr6QxjNXOaHcoorY
ZdAy44S7bGjTpn4xPOvGLlaYknD5YUMMzWwW17LdHc57ncYRESSN+bJ2PTf4NQcaT4O57RlQUYJ6
jj03cNCh5owem8QIxZuhYTln0l39Cn4L+lGFFzx2y41m9WLk7t9lOHhypDKjpXudSvNmjmhR5j6t
1EtEZPz2U2uu8DayTGu5fS0uHK4VFhx1AVk24ZKxvKPe/xc9ple8F2gkclhqmZVbBdQfNGY0VRZ9
NxXx/8J7eEyHwtTXfkA7bHlPElXJdcuZ4Oh2Kc9x+wZa+PQmSH8X1B41MVSrOsNyioMqV/Sq0LV+
m0fyOaYCLAvU+6q/T/xSGbcLdcRsjnUpwnLigNmL1ZTJYN4bnwzPDsb6daHxFvuPwTrtI3C47IzB
L1xRjdXFcxVwlX4plnUmanaJxxKfwyZ4qku65bk5FYANLqwGAM0hCFWf58e0vwpCky4TWUXKlTrh
9MnHPE/GxV/+LFat97d+8ZbXuBZwUucm7IFNfEIEVwtoLno1MPIxOycS18mPFHg6R9W+La795zTk
uzojeLfnRRBcE3wfWmmaKgb9dClJkjpadLd4SUqUNa92dxi11etrTejab8pat2LUvfPp8VEnBQVP
I5kHoP1gTuRmMzFt5p7gbcYxuYuZNbzVc/90UcrMnvorr6CpiYKyKSttJq9RwBAeoM+rvYIUfsMG
63VuAn+Oh5pmXuPYFXKUW/wYQi7iwR+UG0Jc9XjQLGnMBwHnJ0eAbwTph1kHKQrqRndOFX6CIvGs
q9XKyq2HbAb432MjY/A/svwefS/2g18d4lsrCulGeMCEXEATeLhrNTTv/DJdXXINVoItL8WvgIQw
KRynWAcdcjDmAJqFn78DfBQIheMvwulXhZVhST7JhPu9uh9zhUJ/gKeK9CoQUH30+78YpSo5lNIM
bPN5/jlxGfVr6eqmTQj6qIcpFgNmBbbwA5w9ie3Q6NE9go9BihMGJkYz9DrxVaIutyDQzQVsfREf
QvfCEPWlaKTgn6kNz69xT2Sa2JjRZnq2l4zZ5AES6YWk87LZLvyDpolzqt1DEAh9ysGi3FtpF8dh
oDIt7WadHxYYd0TdO3BCQ4A91KQn9DiPdvhL2kcIE1x9Ks1U/ps3lxZoCzT8NAN/KPkUWZa8C9xh
0Z1YthKzEx7mPBGE6V5E7E9kr7J/2USNijD58AaUE7r2ifb3iKJEI4Tqfyat8+DBP+TLpV4cj6sZ
KmyD9aFlHJMgYLlmPy/tnL8aOo0cOWv3po9uItXFM+k75P/fWR+hUppyk9XDyEf2c8JG/eb3u214
ui2lz9ECULpVq2XdgZAYForAH1nqiNcwf+FwwLlfNp3VWpfwz8LG6whfjCcVelgzYlPxQgVpX+WW
w5fVkpevjbR7oppLwfBCdMcmTAc0fPkDpqI0uYlPCqXOxpxM0WME3MG4nT/HVGDtIWzfKwmkBApO
9zwIRhVJ1t3LzPCVxYG3sQUt5QpkxxcS+Gi/YSN1nTM5tDuSP/9phz31Roz9/t4lq7TkHYi6e1Xj
Y9Epoj7J24YJ4zTYOnMwmFj3kPCGVQGaxkv2UOkncFTcTYhWissuo+dDJtfaNL+L+SZLgSYUth8U
b5ESwcCwDVXGU4ApFV3N7w0OgiA8kI7ohtVa0+ZYEEfg7vCo6tzLy7toICUI/QtNduO2CYzwmuPY
fJ1l1QFMBtnpCwRxIZRld0Rte6M0CYhFO8mPrpxt/tO6/0MCafslohUORzx5tgXyQirUxE+vq5d3
mFDGKd5kWDycl3/yFj0ygcxPTcPMreG+dd/BR07Y4yM7sekUPt1Z7bmEv++EAXX/+yMk0NECYDxx
XePDUfWvzNZRKHsQ4FxdxPKqEX8ERCNgzZYNmkZoYSYYZ95GqoY16M0pOwGqeKj5Pr8tKi/Yqyli
Y+1skQRM/70QW9rzJep89nf0bN9NgBcYTiAIhhvSKMM11atcKo5LJAJ0bnRevpENJee4J8+OR5KD
gB4d9K7WT7oVzOFy0yx58Y09HexUd3qcAmLGJoq+Ai4wPKbZ+eG+SPF0N3QmOfUBZHNi2mvyKKzC
0TvWs/2qeT+4ku3tZ2+KRZsft35z3Rkw7cyzt3NDk5wTqRCPG5G7/Z4mTPWOpWB1ekpeGNU3y/Wj
jzcCHpXWpVq9/CukndZgezbK24BXbtmrAx4QuaknzjkATYbTXhtM6kG0IW92WxKUCckdiPoW3lPN
MgixhpOVlzvZkBLZ5J41NzgNI00s9ZYt525QQFif5tr7+XkSASJR4UCrdBWz1O0vhXB/0CIbmKHx
yWH6ueYHth50AmCUQAxkJBMHsYzQds1m+Zz8YPouygJBn+dmAHY20YUMaZZ4g0QCFGkHYYu/Nn8n
rjNYDkpPVqRG9PHcWkwEzSHmWLbSB5g3Ywmo249sxJ2dbD+VGvmeW+cvEK4hISu8ybNVVn9+K4Zw
r0YqHmYYhneqSHSHZPiQ23ObqVNQc+3I6EjHWTaIGcAWIaKADl/dnS6El4T9+p7mnXMA5AWKDl5V
V/pXkjmPhFzwzb8JvCuEW4rAqxOiojMLJpSDp2SxDo3nKPZYXrZ9oiD3cbGRgeKL6wK2/5qEWerR
3uH+OTip4qQZM6G087itrr9NV6+2cUWIGvxoCPow3w64a62CytLnlJVuuzFn21lbPSQAvqjpdLFb
FfBDA8u2/r6MlC0cx1zwWnee0WTXIx6QQf+lJAd9M5Cxb5styB7naxdQHavA/E80gonZPH3eIlXy
+yVmM/bx8B9tmL4vZ5tXLFeoHhUawBZa8marmDKaXXt7BDi6iTTnqckpzv8q2+nN6BI5AAiRtsyK
36aiF6zwp9yOiDWxJR4J2dx4yh9w8rFG0Qb1zRCcpc3qitNzPw25ZM+g2Zfhs03iwGQk4KE0j2Ih
URyYzY2WakSYAQqFUSw2JNwki1iNjodZn92NNpAUzo3uv/8mhUdOldb0QTTXBKXzEimJ2P28f+OT
3d0XkQ8Pypg2a5QYHgUo2boj/BRq3AgYSSjWgBA3FYGpnvSWTeihPbBoWEumXzZsYleeK7LbdDwM
snoS5y+eFTJBBFj74VUAq00i2wcWoGyijkk1Wug9t1ET7uf+nlenYRsIkorwQZw4JucCfbKETuqB
N2kEf91kJTriRpCxAgG+JAjxnKtkfItbl7nfWW36g8Q8k5VeYmnTjR5yFtWEIp4KrrE+axMU4Gue
lL6wCKMQy9Yxaq++gMGwd2zETH6BChz4nA8fYuJw+TQJO9bsW7aL+jM1Vn30PxVtzh2kQe3YVcG2
qeQI9Ocnu1TlCFk3QQGrqmna5i0LHHDPgbiqGG2Hwzk0IR26bQcgLqBslQXlNxrSUmk7A1OoRmUg
dH5+qWAbZK+Ddv4tLt0HPSEt3hPPg5bqSWxQ2aVEsU1wF7+TpLbqsXE8osiQbed7e+lekD89weJP
qLYbDIvSDwxX/Nvt2J/8haCdnFSEICieN1mw8mOgYGW+g5O5R0o+9eTdqyPLtZe3F1huxz2hEWvB
1K0D7E6YyTNIcZfKjp99dfJUbXQ92SCxewtcylw/StLKSIHp1q1FgYyIbPjKhHf53qb9BkpkEVD+
oUKbbFvJEa+ZW6zqgV4AnZ0NZODkMoXnp/JfVjtK0T8pzc5+XHu8w/KryVRO0N5zdi1GRTet/Uvx
xKqIMf23dkGnXg2Da2mu60RGzb0PEY2/fhisj6KXcpdH2KBgWb6pspIp/CYUbsLQpCc3o70G7/u1
Jrv/gDgfwiVwJLgSt5iPycoUKfrIyid0h6hgvYbOc6FYsEPMnrI6QzPZ22AnU+OVZ2X9j+WkL/tW
cm5pNrFeTJUa9SOGp8cnUF9usvtdvuWbM+A5byXgmRW8LjygtUFydGaXKoa7VA2UFlLYNbfSGxi7
1RV5W2V3ItDQtc5JjQrdUaqPKvHJ05xkEPld7yg3FLZuD/g/7igZfqH2kOVppbD55aTaaQVHCzNZ
2nMMJcTQjwsEVsu9FivuhaxzXq6t+I4l1rP6TYh6wBYB4tEW6nf+ftAwHWYm0P79IEdwpoKFErlS
KWdLfD+/M6MVw55dO6kfjuStpupzlb6c7g8CiX1S0w50SmekqyLFaddtulsMILyfaqTKulmOVZE8
qKQOrKdod+RcK8321FjSKZLkMVXK8SLw9XLNlwAq+lulMjes1FVh5JCVlrSQgLwMeVHzmH0559B5
b0GJiTdAHTlZcjkfmkcrDxoXr9nKQYiUqPcLbtPtjdLw52Y2rVBtSvh6mKD8J5Mw4JebOBxyg8bx
2xFvQYGHN4Y9U0EC14r+sJfIdjkl44FfM3dIwIY2CF8WHlCl7FWZHkLbxz6A2XM3tqNSpx1YFSBm
tiiP+g0uWEJP4QfhrhuK+TeQdpEBGU0mt9o4ws5sm24o2jRPjYwf4gNZbLlOWbOwh714nBC5anvO
7J+BQp9Wz9Sr22hWTw9z5LAirEUeusxQCRi06DIzqK/HFy/HWu/DMziLndSAVB7wvdy2R3cS0yuX
6UVFfhCEx5Av0qcqIC+velFUfxmLjw+vYYLjAQKW3eL1K9Hu1Ysp4PowkqC8luBRq9tbmP0Zo+fe
QQjIh4C+YdFj275B44yiNFF2TPhjAocxesUQAb+pp8ELosYTmUfx6LPcVA73qSMOl2ILi8wgT2HY
k7zPW6P54NOzDq8djMWsoqCxrUjjaPpUbTZwrJud8Y4BBxq1v3St2VzTsroIctuaNKhIELl1r4xn
rhbqaO2tmwge5ez9EW370qrc7mq1brICLEu7fQZuM+Y/dC7sv5brjV8LjIADn6CitYR4Zdr5yc9M
UqE/TWzWlWkPQJWgq9I5/438qMX0uSo0hNaLe41m98yo6Au2vg4FRq5uNS4LfSK5hdRo8QcTZiQl
HpeMxBknooimuTjJJVP4VaDTJcmF8117hT3w/cDN+1MuUIhsBidjtB+8HtO+e55kCRg3jpbXPoGJ
DAPPvGG+FMQmVf2pgtwQtEf1wKEeqtb2zbcwe0lfCgiQ2iTrR6rQq4GkqfyA3DnnpXCybXnroB+l
LDyZPK8ZVTLo9oPf3X4ZzwUytgnBbK8AMpQ/4lNs1LdTQeLBWrJpeN7oZlshwDE9TxdkL5ggKv2T
/EdaO1zBM89YWB1QXpxjC4ZAHKxAp4IDqGRZRVfpHQTHjsTrgRKPif6jdxYRPjr1l9J4fL5HPr9Y
pDBFiaksp0CnHfGPTjenNEDLoPHi0GLTGY2qTxQx/61JNVJNFXMq5NLsVQwtHDTlnKpXwlKZRh2I
KUKtTNOj7lS0XwlNItsd3/m3sP8u8DymSdFv5qIuRqv/VAQd+oGqJDPRiV2z0OPLx3AIpC8JrMdg
f/tYuGlwKBiKYeNyxmuJ7OVuxDZUKhjzWtU8bmjKG4fR7lIMX78Mml2w7k4E6YvzU3zCKHnHzC3U
Ri8/efgq1NR7qWba2d8qj/sxjknOwlwtZD47knxA2/yQctjivxl+UfiiAVhKJbjZRY9DAp2iTbP7
7ITjXs2gMxy4yIqxmvvLZoY/2M+8e1cQfpdQ2gtJDI2U2FVzll4Sad37C1dqpcAiuV60yrYnLSUC
5x6g7TSM4YXgJTnNbq0F2vVNjqvJ71pm1+GKCphYSknZf5a8DM/xp/giqGbcNKNBOoWXxg5Be6/a
yLpBcZ0XokDlqAkeTpdxM+YDj/6Ixsr47R5qEtwnIFbJNu7dOnEWHjXFUy/XlB8FqOY/fLuVYVCy
5hator+Su5FJuzZcP8SJFjUhJKJLe+HD3pMlc0B+zGdtlRmXL7UTn/auOZhEgUglM8aodqoRwUoJ
loL+IdA3iqW5YznP3pRONTPj4/bY4OlGnhcjyLSDH95ObUijABr/1Zd8HrtIgFD2g1o4581GYlBj
dXJ9TTk5X/9WlXT0pgWjuOBEQn/xck87mwDFWBwKm7W8Fahfo2V+P2xiaDqzAUKxrtVjMW2ogEf5
RXUtwJzp8dV+Bke1SI8sEtmsaD08dA2CFyBXJt0ZRcUorB6scw5618QW+9NHEHYIHBR8gKRR9Wvi
Irfxcdb26NFjTZBcETY1AxX4zZ0FZLmhX0RkBkOYEXGrGv1sPvc84q8hyGa6BgFakFpJn41veb2K
V+IrZRwCbr2sbgfiIqAmvwasKApDV3M8DDdQM75NjRNWJd0T7aL9j6L3ABrmKg8oYeBSqgE49TvD
AoUkl+bs+Vaw/PVZzLsn2VhArT+Z4aysu2aoQ0IYBPUbVOTrq6fSrdRG+5TDPujVrr4rTGWJ5YeP
OQEhLdg3Bk3tJ5oRRbIbZ6Ai3fMxQDhbScn6AgqLEc4wo05dw+Aa/uPCipuzy8NEIJ4TF92Jwsnh
HFHzE+mRvE5piKqVPfEU/tB7kwN3Mgvyyf6jpFWgTTbpuccsAEp0phFRCT3sdZSjwnuruGZ1GVOv
2YE5QHqQ9bPzZW8K6YoKP5G27j62QmKKKbIMyJjF6JqxKGvm5lb75e5TaOwh4m+Mi3qtAbDp41AB
jOBnjMkOcppiYETo+yPI1ugLxRLW3K6vIs6dNmBpZElvXWSzBhc8jnhJA52jAS6lwubr35QZf/Er
gm7n3t+dehKZF2Vj1fnzJzr6ta0HFVmSE8YX85V4+ZhGyXMTTTJLh1vw9H6sINF0c/isJtaZeoDV
rETWWWEXbxheR1xn53S1jGFU0QcplkXiCZQWOrHlN1qN3U3DGeG4ZEEI5fYaym7oWbANwFnxUVBQ
jvUTAUZ7Lo1HLIiHDL8hZBpAIIE45vkg3xNTdwSxndrWRP9HMywp0olwsCBaOO0SMRemQQpIzqn5
xdoRtofhI366EX0cAnF4Zt8PXvU8RvKUxQvW09U1R553tIc3umW/GATl63Ct2BlXIaNyPdnPAqwc
mLQyJZueq7LfJw6aHTezmjRZmsCBcbkg0qX6UbP7KVV8AkzjwHsTH3TuBmOqe6QPhC3OnxfI5/12
bkfGV/xz1R7D3TeiYaYBTpJQmdjc2PuIe1eize3GP2HF1eGGuqYcv1vqTelrJbRSeMnPgEXKhJeB
XAfy++wrkbccTp/4dy9hmnjdUC+fq52s6FU8pBmMoEgnCVM6QkNlmHdeP7AzAIiyzjU9VyVA+6OP
gPUYE7a+vyfpL1JPjII579pLE+HdXvkGgMpR8jxeH8Lrzy1JTdqLgjB39VfJdwsVbHhh+LcTVV7V
298DZvLb/GKiaPYbAvHpPdtjJZiK8lC2ttc+dE1iLtXOOuw0CLzLiiLORyYAs1UxWaw3Md2gC4HP
aiEOvKLzVBV9bzPcPErEU9FJl6zgibBsELYDYwwiUlS6Or9CtaKl/KzbjeFGINgq4ZLEvI8yKJAf
+/G+bhhPa9uBWZJzqfbe6jFNdP0Es9bnun3WunDobpvZ90VkkVdTzcER36nwrCSqZ+lp2MpLuRgQ
Hy6mbthAGEdzjG7Tks452Pft3YZ1XKFYRsIMlTlLRB0BNA9+W75SqJTxCuOtQvKHOlHluRmoW4Nx
R9YAb2VxBUujBoLUQM76Z377lf1xFGgaELgm2feDX3Y4QHeXjZEXmQLn+9UQPPR8kNJ1oqpjk9Q+
IiqSVR5JP8xlVX+EQ/ihyQffdBGn1qiHbZghdABzzu/z1p7SFijO/LdV+45JxdmpjxO7RsPeYO11
kk/wPLfcobk13Rjn65KwRCLEr5zfuSEqfhkFR8gYpLVGMJqQ8cLhGzfhXclCU6x5qT6guaQYWZGH
6l+tT3BdkQOqOABEeDzX6zJsDVv9l4XxFhYAXR/qUReORTp7aGcEQ1nHPdtZr5OTyyV4lD0hfk7u
pvDlYo3Hm+us0U+gxuoKEUXTedF60F4eZIUds2uiSdJ68oV33QlifQnfFz3IP2WYPOlnZE63X803
AF4JCG6nqM8iWTIzrVAqYE++NtGOKvysGZ8EEiUVdCBcXCTZuHxKb6HnICHCGCSaKcveMwM9X4zq
LUGXvo2FimbDpZFVxvNTWduFUFot8Rf54rxfacgs5JzVAO4l+lRud8zZI/PT/cLVSScCI01ZI5Ng
dWW7a1GwU5CKe2b1ol5ARNYZtef1ieVOOw3tc6rxGh7m1ZSHVPHabtSQ9oS75eSTUTKF8HpCrL3m
LaU0LXgf07QPkf3Gb0nH7iBGDB5NTQf6wBQ5gec9Bttzuu2NNqcJJme/kzDwJ137lc3JUy7QzLYr
pOQeotoG0OuQM945jIixw/NAQ/NTqEKUGFKfIboxoIV7fIKRd+j8u5a8LocaIJERtBoYLAapgHNu
eMi1KqbyMSPxSw8/JN/1oPqlcGpUqfiGXPj9OdBs3JOREZ48iNezL22RXW9fL1TN770Zornjajfj
1xctnh4v98GvSPO/RSpDi0yZaNRUCtMJ4OHzUQ7aBvMhSSFHwicC8W4lQDNngaOeo1Y3Jm9AmF0P
GWdtg3/UAgLRe2Ar7xTwsrCXRJFPB188HrMCLHHkZYlGgyiOmpGEvgEQj7U9A6N1MtG3EpyCqMgT
cr/G4X7l/i05GxiWbKGGCmpRFOElPc9aZZXCJc0AC+CwjU7JHdda0r3nQ0IFQrH1n8pgHs0Kd50q
TlM8dTVCHQ3PgCdgcVaTrc1bRH4zqt4jiu1/P3Z4opjKLKBm0+opeJq8dXFZSgFsYJyoPS2NNj9j
NDFt0J2C7rAalXhauoiLjpSn0rrOo6AWSEEHbBjRC7uNCtKFIC7Q4GSPo8iVQGNQc4OBs0F6ti5A
Sgohn9FmU+NKgjw01Q17RuME/j2ril24ese7YJEdl2mOdCKnXJ8G+jzDgf5wNO2MiKoAP1na1CVI
KyJT67yuOanC9EIiP5Wjio+t+UV43qNaFGMhTIR51og5TdvlRggz690Ng0d3ot3veK9rVjSLY9tD
KZrMppUWNIsIDY8fuIK6V0YohTTtf82Dyn6yH71+cxGCVauR6r5s83kl6CUFXslq5v4sqWK0m86D
lwcgXnqhG5lXSZRb1PO697kPo8/1pd4eEh12XuwCOYpTQWZiHZLD7mnTG9ZeLSTHEr8cLrZpBOja
rLqkgTSW2vGFRyS8QMNncFCXklBliFnd/6FI2m3ov53Wl6ghMyUsK+l3VL+iI2F+H39kRepQYCM+
MW1tWYO3yWUHaZQXYK1zY8EQAy9UboJP9XDu4c0xYjB0pgNyxzdBPi5fI6VlzV3Ec4O6iBXeeZhw
l55bzsn/Et26P/hk4H6Ou7iQBXc52dm9hgPi3eZNWWy+maiUq+07tIz23qieSrxCNDZ55lKH4gK7
4ZP3BnmpyP2przG1P9ZO/Im/MaenwUflvOhwz5jjAuOGs+/Zwassco4JJ17xqJV3ocQKuILtyapi
uaApxDG8MYhiCRv8WyFvSzE2g6JjPN6QRZOiod1FZ525SEMueibr0ix+Jb3zOwS6upbkKVHEEkHi
w0KFTAKFSytgmvm++D++bYiyzafhrL3FstREaYzoL5vsaksT7kfIVSbBIf1rc0xsJKdfVTrIxIK3
PYXS8JxOGpJjJO0jwczUjhNd22ujbbKtOkeGWysegJfWhUDeOMIW5zkUZDIHhoqQvucZuNdp2G5z
TgOltbGuiJSoX4whXvhOg5xuciY+3ASbzoGIxHIqz0YRTH5nR+CN/Rpd3ugM1IGZIqSyXXQBcewZ
98e+Rx2DoWItT7kalJKpdfTas4mR5s5EhMiBRpi7AO6ZKehibFsa5TvGkYyNqUdkXaCfnh4h42Tl
5DqtiujXPyjz9L6bzwgTPTTO30gPNUOt7FodSH+MvS3AzooWGrIJGqoUYUE1ovDFsMEuLf5bepXU
2boUnvwjuwQjEc9M5SR+FFU+ADoLMizsybLJSyMmfEmvdAbCnK0yJcRlUTcvov9ovtsXnZkJ4hpG
bcgWYq/PUdfSmOKjKsTGBwWme2d/f3thFbmLdbCM2QQBKBPdvATCYt0GA3JxfEOBREzaCiTXPMdk
3YcVUDkJcfZ+YgqL800JooSnGJgvgSH742cA6ESOVfZXookSY4aDGp4OjvLcsHTPk2TIpXGtcXBl
Dnb5YIdtP33Hd6bXKsbgjaAqVdTHwu1YZPrIZ73vnFOAY2gP/ZvXp4HIkiCuIpHQlRWqNiOVLBgu
c6kkeYYPPZVkozl+EH4VbxObDFjEZ+HxjyvEqyRiJ9UguK2G5t3jvaUonEdKF1H1OAD2DWVksnKx
6FICsEtAP/zwxQVeLCWWZx6dU14n7Ghu7HPmYGltm8A9QRCix482QlpxVv0ddwFZPwdh9Ob1TcGC
0M7XDqfGKF3SOufKQxy1Dza8ed7g/Io1DO6SKTPfj77OtvMwbZpext/dgSYq584Hn6yH588Ptn9i
cYF8zr0s09/Gf7cq9+HhCoXqprx4qXqMyVCkxsqSmAJja4Ix0SWr2KGEZmAQZsw8vftoHo0qljle
9Sx+X2z0tK/DmbYFqyl17xWO7ZJwRRgBmDe/3yjBCyoPU3NwzixMpXFIoBGs5HZ9OcUGPtGiuHbb
IJWVkVETJu1LqhUQgbaZAKeJQah2LBpXgN0w9eC/ZTJuPbQyglQmZR1XpItCmRVj0DcrySw2Ojz1
z1MdUOq5D/zQASWXsYC7i8TioJ50wacyy+Aot0El3W5www8a5FHmfQnePWq741DxzmlE2BnJud81
vpAW6jlvcMbvp2cbkXswFLqbdLW+VD1YrUYEdzKzZP2zqECL5AcoyK7AN/Lu9OOxADqP2NRg1x1b
RgMEoRZyRWOVixHAUauFvF7UOnn90DGnKJJ0PFXy32+N0Dvt1/ekOWIaqqcFMrBEKGVcwDWXXI/3
eziSB9syybY1rOKmHBhus9Ar4BaDqDJGpiVBFytc9sWw8rTGch9poZRnnARKAJDc3ujBlGPpWg3Z
LjnDfz5bcuc6kcip0YoqovXp51WNhRtB9mDjnVC9G09bfVLWf72wHY6yyW2Lk6T+eXBikQ7AaUl2
k8HI7v8MJfkFaUUB9odSuOKkoKwEXlbcN47j5hOUqnb0bg+rzs9l2wJUrvVYPN+MBDwP5BggI2xS
fcvXvA8gmZtbX5oL2ByYoJ9MrT7zXK4QX+FPcM9XdbIOkKTgtVg6Vw4vC58zBhou0x6Ut/B8FlJk
PzeLgrPNay8Wps/OLpfPHbqTKrWoIbFqcSrSGa+RtdqforHnr7VUXCrtMmvNN3Djq5KbKtXkpY4I
98oeLW4T3sEBFrvVZYOziExS3goXwkrkRL2ZbqmvK37quGnVRw5ClbZsVF3SErpKcMhjkC4p37Px
lTQSt0f+20ixbSlZS2uzR/7hQOyAofc7XniJmsQo1G06hfOaLvHhpH7IKSKoiwc5Ev6adn9BtDON
n1y9ipADVz8M1m0BJq94Jm9Al/SklhXHc9EWL9jRfDndS5JfCCQu1bzt35xrirSxb4TyFTAccL5U
2nBCUfAmCbeqxxB+g+tOgOjaW4szd9Exwpbo/9kwhnvHCDOaaIxCyFr7HVhQrxJPZtQjZGlHfd0m
JojE/e36dlQx59kOyrFi+K3qVk+mzWPm7i6LhAz7fZRQRfy2BdVUEmcbCxXHm4f/hzYpbY6swLr6
5T8CBPZmbi61pzRD2+fNcNXpRtZQBBy8YCfQQAyZEZO/f3ynjOFI6abgKAiZM3Y9/xplGCXlTOJq
6CZJsWZa6jmUh2FUFLh9KufU0vB+DHTI8wP7wv9QMLR1pdHKmpyZTM8CsgDbKhAokcgDe3UsNtP8
+hfxPu/IUU4SzFlx61Aw6D8Uy3wy2hEXiGe4YwFS6COaMmsLYcJRfqMsLAlIpS8H1CXWey/5P/dZ
m38e1pQLR+vN33WXsuAD0FD8y34RfTRrVphAw2rJ4nbHoldZhhQVYIC6IKb0gp5ni2ETnBzpPJny
aVljIMPfppYt6twT9kRt0iU2XOIMXUr3cg1nza4730EBff5cqscxa7P2FPnhLM1z+JIX0UDh72S7
aykctL0CHYCq0gifA+1UG/0aLD+RqfTov1bCPeP3SGsP4+NqddNl/nIH6LEO2oCu2BB9856JRlVv
IRgkU90f8Q7LUEUhj9KiAyFqQdB3s/DgBo54hIf5bIO1GhjgpOxIWRBt9qzTJq5Jn4x3NBfprdX2
L805crOHAAA9hHMVrCJ9Vn7wFaWcFmMUlXW4YAvSWs1bHOH7hDwe2MWUs6gp8xfCaSMYYAojbsqG
bpnjOzAmdK4mSgqdqnHtE3BYODNkN9zgilsbL1T73uojBDw8ZN0R1pa6DXD6pbO8GH/FEfAqNH6l
E9+7UT2T7X7XQZbnq0nk6A68O+svMWbFKOsQymsSwTlweNOen2H5n0qwe3KxH5ItMGu6p1SDdm/Z
8BmnCKqLoWRwFZLkOv5z0VdarbAZZmB4UcBr8vOyealMqB1Blb5DdlXxZcAJtAnh+1xGnKLnnn7m
DYRH9P1atwBnzxL/arZjOJuNY3dfIM30Ai6b03gtgOatbgRy7s65g+oXF41FnrRV6R0qWo8flosC
IjgVYPgMZpMF2mSgPlTVpSmp5Rv2DFn+UYVo2Dzpk5mPy43Eb+4PVgErz7hA/8jjnAJ6fVzBhcsd
EGA4PdVIbxuZm5SXhBtnKULKrcs9/4NCTOaDIWiOQiHcSq2OJlu2v2fUH0NL7TN5YUiOn/jYisyn
MgpMvwdS+P9EinhI8Ll5CkwnpS+F0c47eLnYahkna6GTbneP9o+I2aiPA+x4dgkdZ79+7o8GiROV
OSeqcd1DHvljuEz47zmfbBGRlt5rKqUqL0Vd3sO2h2cz4PtKPbWY4YRXOg7dfClNnfFBfmLH03hO
sAmyLPmvS5/BnyNtVQrYwGMXe8sPATx/Tjqu9fc1G1MCz5mZUzj1xalqn7kTmiSMTIQjym7rNxZn
YjwErH1vW/b2U5uFMal+p4/STRgCSjscsz0dcwWDvX/PIkw67kaMQTZ4Hfpn/IRA54zpCB5Pydl6
NPjwnpTNd/XE0bnGMz9ylUm64WCrEs+mi6kkqRmds+zXYoFDrBpI7T2E5iRqhXZ+F29xYoNzmdzz
slMuNny3AYC0NAxvINkbSFH73VBRbVezgNU4GDkUgC2wDLe4fg/F5uQaUuittov2HwDImyhQxY8Z
Umef+eIZ2w7UAnd02DiqFVQ6t44RLR/kFheIkAJ8NAI+Lh5DdoRak1PveG9AQIKBc48bn0pH4Mr4
8hnQ473YxsIZusbCFM2/mB+YDslZq5mRjLyIU4bmjGS6e7cmYKXg91zsteH76n4xbQkHOuJ0j8QQ
bcCanhuKdi+CKE/YnbjXL8tB8N8XA5bwP9zvmJoMITXKv6ScPBpTvRUR+jEZg+jCh4opaVXZPstT
+uKlYiJ/Qy15w5gJd+uzg4ZovKYlM6FmZEsxgBPl4tRN8qoJkSDprVVfrKfkJLmUPu7HD6LihvV4
yDQmZp010Mp62bZkR39a36hxELwizzw1p2vTyhf0w0IWSsBbS2RpV8AjvO6QcaDZ8uWYu5P6CnnC
HgxxDr5puso3Sw6VoNa4zmuq+UN5uNo25vU1OdnwRftzJGFg8WvT1vaBy4KRx9IQauJo4KP1dp2h
ZO+jIF0r9XtcMilA/SPr+iSrvpZj57Z6RLWOH+fK9hbPYD1cq6lYiF3uU3WXmxbcIr1NVN+O1eKe
3hdv0j8rVwuB3mzdX9yU3ii/U9htNcIb+9N5wdtHhJB/ZtltEeoOpRt/bS+0jQofr85XAAYKOLhf
MNiXYYOqL+0CnticQS/LwXlkHLbE3mzfoP5yBfc5HYkojnqDxuD7uMFhLGpnPmuVTiwnB9rQaH2t
0tEIgje7DF1MilN54yXUkiCUElF/iCPoqDv9MzJgcbzecFbSH7JgbN2NYqXeYL0svCDxOJMByKBN
sSkEwYmcrYoeFiHcoO/oDNCCx52Wzm/cF8M6nQuOCrE3eRQZQQDKe7GM4IhYbaoEZIqgPhQSnq4E
fYHAtPMLe8cd04geg3379hm0sSjlIoJwC9pc5v5uVLc+RSRHHRPfuG2fdMNd11qCduDDygN4zHCN
GWrHC/IN9t/HlDJO3G25cP1g5Q9ItxtPTnyCQWucIUbQpDGQTo0DjuZQNCzmELmugcx0aGKzrT7B
BOzZp+/stH6Cex+2QNGxqx0k9VkRVVR+jlDWyQhM/dhmEMzeevv7eeQFcpwTuBiPcCIpxUQWcBsP
dG0FOl00VJ6xk81mQbGIydmVYIEogBOkqjFVq+nKv+ys2bVjC1wBLIsO2xkn6DwZZeR01ut0vuEN
uDmHQlGWHuAs82Yr2zn0Ot+TuFW1rJebjr/2io+zSyLSpNh9wNoqYNC9Yrhpi1QFh6bU0tp1eZn9
lBk1uGNYTB8QSw01Mc26lGQgYq6LA0tkkyd/nEIk3xrEfhzuP+Tp1dhBtBRtPRRjHERF2O8lPz/Z
g2fDeILL+XwNYO6q/bZlelopttfrPUdGCfbZ7yWRdUqNtSu4pcKN3xQQWC51Iyy8avJvQ54lkSH2
jy17i/0rElBZp8bXqP/0ZPXqa427JkvgqNr93HVZsONYDRXvEB6Y4iL5HVskV/AgfHAwbbIQM4VB
N2u/u6c0EIRf7bwcw1eci8WR1nkkOS5dOAZ/oXqwxzaL13TtabDZkT83dVQ1UMHG+7SUcz3jc9jU
22+ZWWZAz+N9ZJE/+xEYONszwzS/yyJCH0n2UNQhe1FWMVj6rDuY3J86Jx8rXDw9PkXSQNbDIGjA
G6hOYGZMJHnNvEg1JBx819ACXqXbaNvPgWVtLsQABrd3GC15qZmg8g9JMuBnOIGYaJ10S7rO189R
Qjd2e2UY6wHoPK38nwIgejh5biru5vHncCefTtXGj44s1MJocGVsyfp5THCfVM5ibwnvuXrx0+v4
NFSFfdz06EL9eIiFenk+OZqsMWAMB5Ykz4OINr08fG5hgz2p9Q7qVQvhBTMpB5L+OUakQP6jDbam
RqglagaRn38PM3m9urCtOISNNA/XVJx5H9tkVC7B5ZOJtK3OtNZEzKtuWB9uy95AU2mgAtEwLS6b
tmjjfxLE8dV2RJjicC6CLUrqQsJydvSr3t/laNoaKa5YUUuoMMFO9jAphfyFsS+s1fXIQumeKUSd
HTy4a+fqVEFLRTF3jlnzqJn9AlMvIFA36JPChXqFZJHAgX8m1cxhcfhgWf/h/NI0OrzgwpTc7Jdu
+2wzNnVssahROUt2z05BYnK0umyIkiUJ16wZ9Xg0ylQ2M0uN95+/ibq6vjTr3Eii/o3wueGm4mDU
YctiFB+eVdNT9Dsc8rEyhv3iiPzEoushiq4EE46D4kSjyk3oW/89brQorEtk2FVjPQr4VNhrZiu6
zaMD3LKC2J8lz2LKGjmIi5C7d2wbJRqmW0aeJzWk9Rc8G3MEyYVdUEejtvIcXDbO6gaafuxok2Fl
XKRytO7Wm0/LAhoVv6eSpSeIMwNVasyPd/GSACL/k1NAFajpNcX/mPBRNdzcO4MCUpSeyZ363iax
GgFxAFiDIAnykyAsXwdEtf9uOZHb2rvrJ7feaXw40i06J+R+7mQuTF8r6zYZgaCtY5lKK00tILL+
ilqYjsDqOmJoMVeo90tnu7Mtd1uX4ElNcgkKKwAAecjgruZJ/q369OH6olimIzgaSYNgiZuBp4er
MlI+a1TRdzGYPYIRctDHaKXkXcmddSIEPP++3In3vFXMk3JiMHeVT7M+gYggpfZgLSSHW0PSSdXO
H4it8yU6F9CTgjrgv0GJwKKwEKyxTVCZYOz92xNzmW/qkJAfTPgfI4tmPdkefELCsKMC23hmcYb7
xnd2WWyo8VmSAFdMnuxxtifIZ1tsC9lerU3pGBnUMEfgACmkk2QMwLoVw6FJrDV9O4MT3VIFnC1M
Sfaq6sEvqyT1q2sqF7CrcUJklf1cSqIXuGkW3IuQgEyTEetpYt1T5h4fM/7yPPSDV0UP5gPk+jaq
Q5s/CAni9lt80VAoMM1EKLwj8ju7Yojvl7wiw0vltFFnl0leKM+pkFpWYo5PvaivhwjPmOCeLqhb
GGohsaUI+/vvMooCeheRZVQNDuv7ZwXkm7fP6ly8WcKO3ib90hoI117rFsRzTd5viHPab3Mh2i0n
kXgncg3Gk2nFRKYGHB0oTdcE0kYotgmZdfSkbusrtkrJ8bHtunLjosN6l8RHb3fdZ8uRwbKUBx6+
BX/8zz3ufjWuJy9RKOQv2/oQmf9Jjjl8QyoMZ64IcIrTrT9Hh5khp2pL0S5e3xhxbNgKcuWoCxS2
UwrkpYP4Zek4OPynMK99OO5u0iTTSAATQ/8D+9bzl4Ei0YETxkW9CJk3fVBgBNa8n+2b8TcmBHJP
voEwW5qD/ev2X621ePIerjsJWJojrHDsnVHSnQj/S0cvIRUxglHa9tvOvLN+IsqSe3Y/2CI8miAl
PsC/fAPH1++lt0EzxapDOERzdLGsomX23h8pzDM7e6myBYbD0gbgztzWaNiJZyQnV8rOTrLHMrwG
3wRoz2Xyew9AzDET2AiCKdJBB/wzUUCu4aX2pdFfEOkjRSqrytT4bfM8eKIIrPpTYGVaUA8A8/E9
Z1D1AOFJIzAlJyvGgY5X/dqYkzlAzEq7zbFyU/JwMxFVs4qOC/aeIin1Qi3qCcPMMWyFqoPWj0Dh
KFGf7Gvwuup+VEozc9OQTbmONG/FzGkNszBiWtKQFf2riN4I5CZdSWmxghhn1U6XPF2TfZL5UBMv
G9QbFeyd9StlG1vm4o/fQbQXjGDGpF3oPdoEpiYBFD21BqTcxOwRjl1806tP1Nhl2Hh9xAKoe462
rWX7mKc4jmiB3/2Dw8U6h6CXuXgqVfFxLpQmBGXjMmf0zva0xGH5NKpjWMvq22rhb+tniBrd7LHk
HB32ODCqpfVNd4TLhXIyhytl9L5yYkIRvBl1ZaqcBLASUHnTJVarJj4vQVi/p88LOS5G9KbQU+h6
6vOLVYNAVGM/43BLoraMXLFXnYO5YWPxotVyvEheevnjG03j2iA4sDYfAIxXzVOcYXnjYFfgRM3g
X2l20wt6NJBP9qLy/iYeP9iTm4snLUeUFoxCoEFhQu5t9fqx3AQ/yM6ny+ICUj1F1HwHJ12yT9jx
wN3hDrsEkcMgmJ6OK4FRTd6c0zZJhgonKxZayerDOftDY06f8dRRD4GrcscT94lJrvhtZ2ll4yOy
mz5iDXUosTV5x5Y+hoBTMv1exi0J8MIzqjuWfox7V0RxWTrO6nBAIh2HfjIx9miw/sskOchtHHrw
NnysWBAp2RAw/JupsQpK6EerZr+32X51DQHGbNAgIoQvBwkHHFli8X/I/Ez5fwpl9AyeDQIHHrL3
YYWgp/nmKrVY+eVa9Z24fjCeODOkv7XeTFEA55RkHAXRwQRnfhU4oR7nq//Mb77OUscH2JfrfiYA
7Av51yRIs29q5cgxKMXdqLvADBLie4xGnRBHmhad8Le7qeBae3GDo07OQyTgUiEvczaKeAXFG3L9
6D0BxkCERdQYyZ+RTQGwIBccs8vCmif8Nngpt4cnyGqpyGqL9gj95qEhGCNMO6HWe7PKibqnsWgO
5ipDUPJ7f148zm/YYZu1vlUHB7srB0PyGJu4gdJ8fzTdYQvFu9R14XopH9Q9pO4G2+s3pYGyAKlk
p6WIrrK58yC7tRbtibTeRu7zb8Fs3CKUYVhQNVVxFSV8du7VkaXg91wODc+s6U6+h2O4J1R2Wb7l
+W0l4ezdlKn4HlOWt53Qlx0u7osNgYUgsraJEF97EIMbBR4JYmAuq7ur3FprVvuLw3/Kl2T0sjy+
HCgmh+3XHIHoXmYWG703pVgk+p6Tj49iQivga+bQ8LkC4mrvIe0EDUZPAoWt48qZFik40YK8Uj4j
fA2P4c7tMYX4eWk7tUWGEz2o6z9hZydw4PhZVRquHcRBKUKz72fPYxf3L9jyGZjx786rhH71Kzmi
ZF6XFTiaZyzgNH7Z8iSVI0zjijJQhHvvY6jtZkaZkGqunskCrC/VCGas0kmUjU2t3BDm7ePPXav7
S3A7LoPpB0wBnn4wYY0vGUpdqGk/2/FJa2X4j3tgl3FsAmxzrXyoyLrTtTucHhoz/uROpBtOZa1i
dQhDby9B3o2mBSz+vGpYmwQuMWc02Nby/CVg4l/FYgSCbv0EtbSc6ILPrQluQON6IkpBXnz3oJwW
8dqZzMZfzk2U4FAvUHSsXlVe2UO3I/xaojPSxq6+pCyiiqkZUmAQzzwm8xToa9L1tgT//rZUoV+x
uaXwsEeqV8X3ZAuxtXGf0ExXozRHuwPuPY/C8t6XteJquiTnpBKSbm7h4EOByWdQWf3M46sd+Hbl
MtgCJD15QeBaMVp1ger8ylmt7erAZ4LoAT8NTplainQPs0lgs7TJaTgNYGEGeC9PBGxj7vrJCsta
VXyu7GWbMxNZJlJXMtqru+T2mzXakadvR/+t8cM9d/Y9gXdmAiG1lOWPAXIq7eaMG/464MXzdr0i
3M9xEPjDJzPP8O50gR2eR8GGTFje987c1CoLzlYRDT9rVAzvqYsbVjFsVsuXCzCZcxXz9IxT06oT
DdWMmJdupZHfMkBiRhXaK+B/ZmLidg+/mmhcrS67yr4kwhoelKGV1uGXn+rdWIhRUTJhs/As/+Fl
RGEryrfrPm7pWEUbcrn4JlflC/oO4wcRlaRU5yEKTHcy+zWKii+OsFydgxxLPd0d5fzuZrDlB5+s
Y7ezravqTPF/IsgvG3Z+R/4Dakwf8rMM9VWHOF00uOoU6ZAtjQ3xJtgl869K3rHbyCgCp5tsYo6x
+my4xrTKBrd+TwCBFHy3gcJg96g66NJ4ycdyR34Z5ixc2sHGFZXxPp58PUCyCKSsOuoXSXFpzaq0
TTecZ1fcVZ8x17i29m2mtpwdtXQ3X1LRyPkfPSi0fzf8pODP8dG6cJ5p8JE7KBWE7a+JtrvdRobL
05gaWwxu4Q2x51DjtKilXqHt+VW0eSNtRSmT2qRNsfxnUr+QzGplwKhQGFRl2j0R4DKtcKd4naYK
mFpcOEq/QBU6uSLR+2oQAA4wnt43aa3HNuB6Hxpd0rRzHWo1lDum+XDbe0i/3KGzTadlLgiJv5W0
Y3FASgmTav6NQH/5XmHMPyvExrKZZd+1YoJWL4Lkz8rBohySlO9okK02KLcQEO1fc5S2HE4WLr+b
kNwMPbhdNm/SV8bRIweJVie6cwQxMh7zweBH1Zt4QlF9WID5EbU+FX1OtWy/VnMG2U6AoFOn6YQ2
VwKNctKg2HDL8N3RjALDQIUrdyySi5GZKBbBRy09fnyBIjJ33ml/wU4dnHco8AC70akDBtb9Fgah
sb6Ch48d/7yOVJJeTV6aRKyn5ltCWcgzzieMJZD4FzcoavgsMnr7y8WcKbrrKVq+d4y8g3O9gGME
ErTl+M4wchuLQiu/OSlfFbrifE54qwr4RAOSOpRaVkoMMcZoXtOQ9TmCd0b7WViOmFrXvOqiRxCn
cSUrBcEvoshFhje+1mOYzrTr3t2XuqeRMs6zcmJbnEHbKH0njgoOO/yAwy3MCS/iQbm1LmAojMfh
Bc19JLm+3QGrImz1/dQM42T3mB1ZPv3Eri8clCH+fSANeIs+e6+iPGcxzqwNRtdSIomIKRU2Jpm8
ssFXCGuLaVd0cI8RdJek/jh9IPMgOY0qGqSyEBUkwtl4JDb/Yf9czSItIbn5HnTpa4tueNi9tyS/
2AByuZ1MlUuXBYH0huCQRm7Lhj+xIwqNUImScz7J5aNqf6j2g+hvZUxGK4+jTVh4Ep52UjgYSGlw
5tNTOFvZtJCvIEyk8Fpnfcz9UqBPiKwA98u7NZR6cPej3jVTaqZdehBcK5u+8Fb5bgxHOKY3q78W
Cb382WPN0bws/OPUxj359MGt6sW1t8sOWhOtxOX/AxlMjQlHH88nMhfVeXQNAvd1REXoIOp01IHo
WA28qjUv/rxHnptxINaWz9f5Y3nUv5Y1cDMuRIH9UY6dHV+GsbfDcvtd0EoMGW43A6GYw0iQlI5y
Zcr0/nGMfeL+82mi23CwNkf9kadqB9/82ijBkCpLp115rwZ0jslbrxHClVh+Hj+lfoehp6qD2X1p
xmW+kJxBRwEn4QvVZ48QOWMLihR004j25dLXwsXbW5eyzsxcCQqbh+7ZE8HzYRO2cvR6g0cI5YXp
2bPuA1P2za9iZt5MbBXhiO2KtW5cfPxHlQXI3Z60Kbcc3rtGVyer18sctxWWndejkKpY3uFdbSQU
rmL2yo8mnOgQWDqrUvrScQoUnqBU9SXoeMVTQMcpACMAeGIj4OYFIa9oKwiRvK4UtLYpnt/muYS9
44AIhEyNL10yLQ44o7ETgqmcnqOHI0ka12tToT8xa9xvX+uJydO2VGfRcenwOqb+r/bSsxPhrKhe
HBdLTn0XjiJD8P1YmTYHm8ZxjPQQHspAXwCJOXddFhS6QupnfaNWuEMlggjsHxhzLbR2cw59Z8AI
js1QfvkhIoK0z20/LUrq9nnOoHRQ+2pjL4XKTLxnAyHd3z/bDA0NcALpsg0vs7AQtLzzRpGwQkOk
u9MKsVcy0Ppno1vv/dIzMzRX6YFhqziJJZ54iZXyWG0effkuv0YJX2oUWDtCS6El/qh6Xk1g8nDl
ukrOKTKqSd73dZZab79lQgay8uO6O5hDryU15rj1iPrY+FkOsudy+ZoOzRxcA7AFrqVMFkyKIEvT
p9CiHFj/yyL+CCmfTylBO+NrsAngc/al71MfFCI1HAt+hZRp/q3PZQeL0I2++pZCQStxY4tavd8O
EKgOCQw9nLbV/OWKStrABROuLsz9zvNxaZMhhYEvEqa2BLSqdYtTsG0fLNSbVKJAfpHpA4vNmVPQ
xtHex44OJCne9jfNASAVYY3QlZ0txphxb897jEYZ03z/GePOsqzijsrbxYU2a3oaxZS66l1/9ajE
4MtX9gPgUZGLTL3z69bI0atWCZC8fHohzFv2F7lTSasfPa+J0IG+WsBkin8Ei2KFbBiV7pVn1pWj
NTFggDmGoWzDku3zx9W/p8E1v+JAASwzlkqxlfEMcYBJeqRLv9IPApCAf1vwUFavuCrD1fXU68z0
MLrMvOfz17yXuQjZA1jYlrTCUbqsimxSs+eckNazUocZt7vE4+DIBJP/kt+o6NjZTUzPpbLKXZGP
N9AyUaUXGSvtBQqXdIn8MI+5rtp1P+878XldndWCWF2ux6FbQd8/M1BbTkpLxzQWTGVh4XX5ju0a
ILeT/Dt6PZWCDvsAZk/ejbrzZ3vLc868Zm5PrKa9AYm547EiqO2Znc4vddSjKZZmvkY6cgtGTfO2
xgvcwATd+L9Y0TTauuIiUDQjbM/qufUFU/D0tA5QZX2gCqK2pDmzHGtMsJi70qdZC5jHr7kIJQOx
411WnJgjahsK0puDcsxYzz32MiBI0unVHS2JSu+PCU33Cg1nR+QK/5YY15NafDSqUYIuie9gkVLj
W+Iq4rHQBYhzKg86kITLE6L6DywmxGDOKwWM9lztoI/O4CmyR3ACVbR2Ph0PNvC+mc65XoPceDrS
JCU8Was/grNYzpXrvnjkV6NTP78gd0pCcJS7r3OIdCTdxHG4qcBuEGIG51GBrAXrB2jA0p+hlT1s
P9v7ROUJoOh5i1KRGI5VrOx86vtKfdErdcvIlQ5CF9wa3qqiW0/lf5osRCvGi22MaS1L+R51N9LN
pkROUFBx8xg/puc1pYOb5J+e2OIKvVVRaixVfTQfYDOUvPbG5DtP4M5bA/PgnV0ow4yTFkiN020i
HLj1/8Q5qthC/8rHJJgnIlQvje0fzZNB7fuQRheNTN4zqQptkolX/NFPzuvN4nyHYRCX/xeTeh6A
zzXILz9Q7bdBJ0nlhQxT4knTFj0L2nxRLHInoXgjqBpBKpkc30kPXxzt5fSV3eN1L4U1oBwCUwyJ
9etbZmPmF/tod6DM+7q1VXLfPsKOABG54BvC1AmUfnZb6j8zlt5VYLxdj3s1Pv3jJqqdj3Vm5bn3
iVNhm2P+f/lgJxNhHo3K4GLLKe1mRODf3KElUudVkqxbNUh7BAp3TAryMqQZzmtv9dHGMvTOp56q
EEcArYiUs9PNmpHd6T7ZlLE79z1lgsAuKBuVHj6ajK15zzZ0AykOusBcYvIH+6k9zXIUJFhxmUP+
kuAo0ie+sZsZYIiZqhOQBxBIDGkINvlAqjmdkuCYiv4hlyNen3UfRpZCCSM8Y5eSolkl7Q3gybla
HHDoe5Ck3pKNYMHMzDGszDW1aufpf/E5UmkURfnMQSt3jMDwrvtvwEUPa4x9k8JvdKAsjH2qAIY+
h5rgaYeHo7ZzVG80i26JYLJw7lLU4TjYIej1VlBli1s4hvSyAVg5fSejdf1xZH6Uh2LaMPfk5d82
eass3oHDgehlILVGHdbkUUA43H/HP0BC2Zkw/sN3DxyvdNLKDdCOtMZe9VXb/x5zgE9xnRFlGDhi
69BTdAVpE5/K9rpnjR4rjscNmrgroVswvteZ5pQDAyaxmDwZcSKxQ1Mi3eDVw2/48Q5obQZJDYXP
kx0n2Jo6N0M2PsMgL5rVOwXhCwghNiHN2+5DY9nis0SMrXrkitu0Zmn6NVUzn6HbL4RYgxMrCOhR
n1li9RWudwOCAWfgWRS6fd9OAlsIGboO+uhGs5pbj6UUMoWm36VJeZttBl/F8H7OEy2HBhkgahps
4mUawX5NeDI/FMUO6lcyhleNQQ9PR/R5P72qk0u2FrA4vRlKCh2QCVZM4/0kVqt8PNamnR+luCcR
+0BVGag8ye5mHKwF8iCE9oCM52NNC8vm8i9hRbHctlOamElR/XwthtsVGz1XPsZf6sRgQyU1a/tN
glatdhVeJ+KsUiylNQuzd9XCYWDtqvk3NDbQ6tbfz5xd6IQCzbSLDneq3obPm8ACwJOP3CBwOD5o
J3K1Jpugk30yL0LY8KCn4qOo5hS7XIFwj5gDC3VEiUThVsiIAooxRqw+cxK/wSwddgN+9pMKMDgd
dkF1EuCdAsT+gzPejKPV3godXSiWPtaPtIWB53JSI8nMsxOUGzdZzSstvhjX40IXrYWehuLUBNWu
IgamxWYZSrtJEKKzvFaTxeFpFzE/Ij2JVCVQGlGuqwGC0jt245cUkBVsIooWWt77Q/UP+g00XSUb
cD7ZzPYsMrM23NUz5WuzdFngEppg1V6wHHJn011b4B01eBDh3AmVazJgGS1U4pPCp7G0YwUmPkb8
fSskEmDIb+evKOXaVRwK8n084+7/qJUjmKRc/Ll/lrUcGeGfui92tO1pFnYLBhNXUFOKmKjdARCH
xF2hcqpe6FV4w9rW5Rh0c/MdsvlwU7AZ7MpeGZPGCTc5u/LR7XqurbE32qppOwaUxMZRImKwuSU1
CtYywu8QC6lSFsf8b+8ab/0Q8hRFvvBBBBez4YYk8lm3QKNqsX6JJPNseFExcNcxjNHka0Z8jHVU
18ikw0DK3T+fjisYZKxCWqdL6DK6abVBzgUWfvLL10r3dbgMUKXbGMOQmQ7+sWhKjutH+HBVyUWL
E1v5v5I5nGX5KIQzt3Q19dXYnTYpBmg5Gt1W5e+brnIb+SMpxRucS0I/eebP+WyGBM1yzFCbmwxk
Z/llOj1YWJ1vFgFecSo+8LRCdivoJ3SAskVtvPKcR/AYI6CcjNIGNE6v3FM2QqxacxNtHNczouSR
Xufgn6QwgMItd0HU4INX5kzryDc6u7ufxYqFW9BdCgvwFI0cpr5LyfQ2acTe86PemTSGrU5lFbv9
wSoNoUanJAR3SichwzkXEb11zjmo6iRV/r6AyQ/1h7Up2mveH4SWBZ4uD1W3/4bybAc6CBNJaAfd
/bPMijLjpqOt+mrIlnSXK3KLxZcN7Wqs37YapKao+2vFVLsgSLYAXRCWTa+MYnCbtFjz9xtL3j+g
hN8lxkPHXn3uDtqo57K1u0cwCxyKgCAVKji/zPFuEuYcLggAa6CrzfP8b6a3v3mmGTn88FSdU6HB
JM1kF42rcwgfPvAhe824O9n7HMIYjgdx9pSYdUUkaGI368X+bLv2GpwulKk5/TWQG3Etb7ZLAVFa
j3lqNmoG90W60//da+UN0UWG+Pe9yZfDyCSgxTBqgFSB/ol7gpYJkAey0GP/J0LM4Kffq1bo3rgd
T5hlAT7Xum5HmblxUxDYTsMM3LJYb6PnNV11p0F5tSLoCJDxCdMwd9FJTI1iSelqssYo8+l2bLI5
owsixSbb1dDE/4i6hpUtTOImvVfxNh/psbbUk5dPXGWFN4X82pM13J6ODUExb4mHU354tU/LzLV0
85Cqp6t3JhYWN3dI0wYE6uJ5pXEdgEfn7yVPqJZnCYFC6d4ekSS5a2F6ad9eBbY+jKcdPj473EdM
r38pRQrWesLu2akuxmZ+ce3LJDKLQ2Ou7U6pUxCwsWKigCVFq+n1lI0Tjdjf9dlJeUq1mAc8jtaV
2Yr9K5kcOVGRoEWTpEn9tNxuv8XnCJxaxq7sxMhR2TKmCcAHTyn+w5EKwMHdy3lrS3mzijPiQHCk
gBZhHD/RBncnbRyiJcyZdlts9LYK/ZxbdOLORlECOvyF7BOVSHcVOCGvVaXm1kCJqQyhWj2PYU1Y
XDiB0WUNrD7zg2XVizdsdAslFQIqqn14LqlcBONShC/h/oUKU9kLpPDmx+OXB1tdCUIx+hAB9L2g
Kp/F4XKir33vn5izQKXahuKfz+fU7SJDADU/b9qrW0kiaWgBrr1FgulJS0gJX2025SUDKijJSh6A
BXInVDJPM2P0akiS53cWVgwerCC1sIbuEmZ+4tmfpeF/+xAEAVGt7mHEo9ZqZov2ocFaKmAc6HMv
L/vXUoHW6q5nxzAX5goSIoqlhveOv62RCL30CnKq2FB7OvyX8v0GOmhwtW75I6r3whVcFSXc95QY
csp0j90JO1xfq3aEKyMZOAxEgLEqCHv2NSlmBz5mVLTxMWiu6WCtjgOlBlYzSKnrPRvjpKUFSPPr
8H2EutQRiBOBBPNU3XR3T3ZaktI58rS6eL8ckJOBSqB34vsKU482nbbXS4e2fOW/BlToP3Yygcjs
8Wsi3lZD6B8AdPyRHnATBYcEUcySVHxm/HP51bzrPJlOYtRG6Sch/YWvfkwHB4+9nW7hXYKROxPs
Y622IHnWWBA1xJiuLE7HN2z8oYSrpNfZ3JTUqdbXxTyjBprsgxOJ8zin7jqg+MEHFnbdheX9gYLe
OcVa7NJRX56il/24h9q8M0GJZz3G0tTU2XQSSv8qMWmbdA+Z6NTzS8crc+EUwfgrRjYeSQhHa+fx
N7/4Rofrs1yYuTufZ3aaHn/qRuqmeu5cxqD2xssFZgii/HWD1hcV5h14ZAwWxrAru8HuVYxGV9Pb
xGaryjT3dBHOaNExXSLBX0H1xM+YnWt0EUre2GKpigjBX9GBA+MzMYuqDTKEyIASRxDC+NKK8S+h
vsdXSrlGxQLY9kBA6DW76rLWCVsw1LyT+uvmDBhfOgKxrErYKUsTuAjh/Ob86UTgN+ZeMgMFcXFX
zBy8veQFqg7xwRHlc/QKKePF/kMjstiSVfIIYz8ed8p/vmXrU5Z0WQt50fYfzVs5mt7w5+CqslHU
Yx20n+lQbiNWOnLETmkdYtAtVcEIH3ZCuR3UyYsA6pAgcOq7N1qdLgDxehSrqO+bsoKygL91jKTT
21M7g8Lztj+9w3ycGuXGMrkKZb54zRMu4xwt32Pwo5q5Cjo6uZlRLtzsojQJtyn2p+ei+TpWdLsP
Sccmb0BXgv3WkgXy6Y1XQIS+iP1G5iaABOjP3l7lTV2Gaz4HLpwfOJp7y0xqDN0AmLWwSUgWQrE3
7ObeKzh3oMCpYnjJO8QRGNM6E3fhXxekA4S2DYqQK8lOzMTItl4pj/4YuOTnm4EgOcVwu3/mLsRu
p+fpt+Yw7UeWPRTFoHGgWWo7ga5K9LBtjlSpNAXl33YSRaZwAQxXWeGkUPFIEXUZgDfjX/MJUgcX
c63ZwqKOtB+CeAbeXn8ehuymWAlDYo/yvXuOSrIDusvF0ONx8PKtiVo8gHs76DfWh7KIVgWoTfF+
padPkvpR6HKlY86/0ycfIlBSJU25DFZkSjQvH8pmN4zz6eDyIoVKHH4PhsbXpHuSwK2O0QvXpF2z
vXSxzVVXK6emYYRSYx3pzXYBptk5IITdCFm/pjzfz7zHv6wJ2ZjAmwgg0jJ7+0yrlTcLLVKN68sM
D/UTNGYiR5nluiGFPrG2SHwGvwuyEE1oqol8z5mGVRJ0kW/q/OT7Uv+JyWRWCadLdp0i9KUWUOQy
FPd8tvYbyQrskmnAv2AZsGLnehZh7XH67pSo7kd9VH+Tbe7OZuqjKnhDb7sKyZC0puRmINgwks+/
5LfwDQ3fYC0njrak7C3HwBCpLLbpnlBOHbEPCcs/UUbLxyEd8aDDGXyuJ2XlczSobJ7/KPiMpb/5
ziDBfmQiZogNA9c2x8j59XrA+4l2mO1BstUSGvs3AgdT1BugEP42RY/nGPvQ24AcjgxabykKgbEg
M69+18njmEdu1+DlwWW59ptjjrm4p9fLj1Koayq8QmqU/za51ZZIYwa/7po04Q1Ls2z36pSRVvNC
6jwVM1JVtAVQNGq06mo3/ozGbzZFGJcsjZ/p0m19akmhB8JVnTlfmIUxuaQWoBI4L+FksbCNVReF
LJ77bzf1dlXkLus8nmLkL5PkB/9gDBNKSNOMw5bdqOamCGWFESjjRkx8kv0E7M/P5lAcN6XvAprA
a0h/VSZNn659NRD5pnZLkvqfXOCpRAANvB40zgcsxKRHcM3VQ0Y+aXpmNihWfnG+eouVCYRm+Xm+
mXBHFrAsLKd38mRyF8DyWDdVLjHUC4UadLgT7iILLgWk2f2vdl2hFuvmUw6aIkpfhHU+z2mjpu3q
b6FBolLc8eki0VKzTqgKS15hr7U7mVcK0TQWkgewcYftszOJflKSt8XXkvuUR4rN0P4uGLXMjhDA
UCXQr7Qx08wPHknQv9dRuRlOeYyXm0vdLCiRoRhnp4bBD1+p7p7JuU6/c58Dap3FetDrXdqYAcYJ
thf/YzFTHkfuvpVcj4aoZ4RF0tHpqBOLN+wQEixZ/oIYKYE1V5D42jwlHFaku/cVBpVOV5d+dPP5
6ro4MjFMRIUpRviPyuHzWNNcVqbfcBHNg2+N2ea+19kgFI083eLGPT5jIG9o64NT2gizcvVs4HcD
EHbNXm5dwdpLV5wL9Kd/jD87rzEc3l/rcwjANDCt3alOBUAgW9OwW5t6Y4PBUu3vwQj2R4p4//ng
ovjgGkBEUXo4OUBlamzz/d63ref71BC7IXfpTd3SqMUB6hYXbggq8W5DHVFAaMPZtrUJgKSlcZAf
BllYDdOcktym/KYvxwnE7SuBGe/B69o3D+IrDC6Oqex37tpgpq8O4nsP+zc9GUeSB/YWOkjDBu0E
OmC2fMCaRQEht5Hufs1TWoYvKz2lbeC8vM4P5uz0HvRAq8p7eYHjqs2oFlMb+uYHmbM4C27fnU3e
1OCif4MX/bC8cr3Yil0QcSDdqIx+NJZ6FyQYqg0CRDM9AYTKlel6CaAGCvC3iSD+o0E/BgjV84Ca
rfJNxuODmM7qHV5wDhU7dWG3qzQAuMfL1TjD7wLGsM4pHXT3uehKFwkEHFrSXC8Tio0czI0KTAEI
01+RymTcNSUpBiVQrTosjsYbJ/0iYTFmKyty9zCXCre+sAIn0VA2UEDZngAseAJv/0WApbluRqZo
NMouycxqKHqiZsWnk7QES/Br+d56lUbeoktPplsmNOqHPUkEP8oHtCT0xgcKe6FYSoPf7zkjG2pQ
2kzQ5RaQp7F1R9FJ3pl76/O0mYzEUmi8rRYcAkkG1Kzud9UjrH59nA/AM5lSvNdT9jnu9wd0JXQm
RyTM9vLltFp/WG9k6S07P1O1a2uN0LAprHZk9jjBQcs4iKd7OSVSRcGMxv454NvtjwvqjGqB0+r/
iYiL+q4wJzkxES6aIwyRk6R/GZO7Eb+MAAequpGG4advHfjI34ccxZw5vOEeY//mmPV4vH8HdBtW
aw3dF94IIE2Cwv6CAkJH6v4jY41aysTJ35KvIY89dPgr+VusHLXJlIKm1MQnWE7bmFAzJTMzseDe
ayIg2QN0USqELRvJwrP6dq1WxEYXpvIcPmpjf/NVzgH8a3UuSP9MhH0Iv2LsEjIq1PV1GrxRcOON
RGMr1KxeTspeFhOBhVY9+3Uk7ggnHF3fGNqX0WjzmwSFa7UfJBOwpx7xwdW1pqh20wFsAb6VkT13
pYRo63/YKifNsskGmn/8kTXatTiWrlFUROzKmWM5U7r5oC9hSrW4WHrfR0WwDuSaBKf8QYPRimGF
t1PuAkT4VJTGp5ZkzYKC2MFbplkfwceeOm8mcLT8rIQQ2pkF+8loUNrZ/PRJ33H+KjpZME6Bc2zg
0SMqfBLhZeaNhSTcVZx+/pc7ZGvK8WnyxA0LmaqvikFAvc5dxY7lBdNkShZPhLWJP8A/EKCR2Ywr
YUdubpr/fz/a6auJ7nN2WnAl+0vrM698QsWjtdmaFCw3LtnCE47jEYd63XRso/VKRsZJgMi4RSnx
cX1D2cGPQz6oV/QaoOwIspdV1QrGmvkbB6cskHr+RP5TGR2L1yefl9Gd8bpbW0sW7cZq9GEDbLBB
9I2vu6YLmGMkeJfSnvzsJ2DVMeLvaC+ArRcmunE+K4Mo3CFEUSlYG89M1MtQ+DYFUVtncP+t/2fF
X7+cxKi9OBqmoOSaGGMp+egcFox3GRz9o28u1XjMr8Wue4/HvnNwMkolEmlh6nVOwpBpJemc5b+v
IaFKtRL++NlCnj5lq7wmiptH/W0lWkIZyl9nwRx5t2ZF9iEk2A51dXzjFL7I7ys86zAHC2W87YET
rJ1OE+hUxsr4GiZzmfIMVKZCi1HuI+eDG4dBzsBEdAkGc4hl46dsa44QILIuwMF23FtAt92aqU6U
pJ2XvPr+W1f1QbXsDYXTtVsiIOzEE2+W9Kv/kEIR0yidhUrGwbz7RHNKQKAFlsEZ7psgFSa6w8Dr
oqYRXDLum+XBXe+ytoSKbYv6dcGcwqloR2xJtPak91lJ6VaxM2WMTxXsLTmGK7NSTCxlsnpLzlwy
oEQ9l/Cy4x7TfiqSko9N8xr7zoYSDXoLceAT1Z5WlIChFTi7pFhgkIVYDSj+of+yg+2RTOYS5yeb
NWuzuKD9DvjrkPSDMala0zaEUM/xkjhDnYF8yAvFYv9mwix4p+PoIc8ukwAqP8Zra4jkcuqUffMf
zzT4TVfGTlT/Az/JlY/NB4/O/K1iwCs6LPGZR/+foJKSRfEAHZQvxpQJwEej6sL70AjDyxDX2uQu
jNttnUgYjwr9hgrDZeQpOJOv0XmpeljKHJtCZ8enmCJa9bOSXAHP7rh6oHu+ghoemTreuNNHZKdE
qCk07BfyAVaP6bbKAVxqMrujHG69JfbiFh1tah6CImVq7eO3ynn8gek7SkWeMdC56P/1LqV1F825
jcKLwRYu1ps2To/Z9e3i0LXaGuwPTJCysAQJ76gdSVv482JVjnhBgZCnJGgij9yltOMIl/SNB0Y8
73nVc7yObpzc5qtQ6GZOjODE5B2zeotXMSTSTxts86utx45nwaYZcvB7Ik+x2E5m8xOuoqmOmlhj
V9vIuau5ypNpsGr59kN5hi5kjPIuv3m9ZVXTPTRDG7GiQoTLbTZZ44N5CfSBqkEdqCLnfClcfNb6
mLiecpZRAdomlYwpe3UJzcXm0LwWkMH+4RI7nDDcQfX3AngNGg0FqTbVMN00Rj029UwELKBe7lPL
R0spuS2sNOVjyaSIVwQp0LNg1zE5c/ahmIOdvc1GHNG3bZ0L8KvDbkqmmowDoqwVjbUM85A3htyY
jJ8fh+AVA6LGNUMxG5mBktRF1yC1/WaT+8UKfil2j8gpntSjY24qqJgavqizh9AFrEOWcZQ+asNn
OtKZEkQi1hBO1wUqGwdpXIQ/bnZHFkfbZTf8lyYCRyZ3WO4nKatkurFcqO/+5VG0yg8DgnEyYqTD
d63StAnYYFMmZhFKn7IijQm++vs4Ckwlyq3U2vq/ez2lBsyNUloi7GclyP8VMMXNE+zgK5s3zXMk
qy108fXW20PFqJRJqmcvLefGaGTqPHj4sQ6RH8u2GD7rknjesx2igy8JV0d9nGZB0gxHXf4XUGzM
xljvODHDF54BrWfl6VnC+F2toFDWH84IGUMW0ysF/x4vMfJup5+jy4OblcOoQVan1QXfdXanMrhM
57/myn2i+f7w35c4CxAoWWr8lCTjFyeXO0oLZGs5UKovZRDlNgRV1gM6jWdUBx46UaVg45mEMFYz
LMV+UjdxwXByGEEAmJJysHMxvXfEDNqLU6vypCVCRemBUFvbnHlO9R76xhcNZyHUYbbCCy0x/K01
eN//ZC08Ia2rTDfn990gtzuXabJdRCOSBptOxP0mYgwgtsrP5anR9OsxdzlRPPnFWQmhh/Widi4A
4HbcWUzauqGUGY3fdYc56PrX5qvrf3AEqJs+aC478UxkwGIFgYLKpUUMgf83U4b4vCt4qtVOGa/E
E5okH5bGDz4z1Mb8/OjKwVI0USCSkWXwljFb2QmeogZKi8cPBVQCZv0Qj5k+u+9zNADWtcgBfiOU
K93+xeQUm+KHGYb4quj7H8nkdl9MibvIFDP8fygL2hPze/lJDCO3UG0XpK6N34awvwOp3BDc9x8H
VbFS2sPvxrZCRMxjqgjDKLOiO70/RLL2sMqYspj3BNfq1m+tvkk7z3jsxV03O3aUqPj0e/annfES
ivxOpYhn4pIDt0xtwaILdUgFZxwSZzCC7XCsreSwQRNFc+d7CtAz3RQPJRbv9J8+ZNR14KjrHv/i
WhtI13MFfIUw02KWr/kcMwafaTLLPwEePNzj9CYGkE+3l2UuRgzTKOaFKUuFPlsce3ecV5DBlkS1
vhwqxM7FHfxXN7A0wkSXIzGgRGcreGI96m3DvX1TCQEobX0oB+MRJaPzCFIPfjAcACFhS5TPz8tP
Mjm8F4rdlHAd9MYgoPYmwO/NEoXSF3QiwLx5tSE41c9Uzw3yCAl/ZHVsBPSY/oLEEneQKmVdg14A
zTtvklQY6Yv3DfUHcyyah0+irpJz4NPuoNplcnvCbijRGnD0dEByONamu5LgqTT4mPMfh/rF6r5L
4xVaImkDwRUgUlcnTictd44ENeoG7+tlOIMZPtA5kLNAvSz5kwdRo96zj7dyOKlyXYi7vuix+4mA
n3qnseuL12Y/ano6o49dbk3TUNSLUaECkoHbGcmWKR+sTswPxr+iBkywYxTlvkKZiLx/d3hW5Zx1
fMPKBPdOpy5kNUboMnxqhUC24EWmcK+d1H64S4YGNG4SnAOYJ1+ljWOHlcp1JZjej9xiwfyvOYzv
JC0miiOjcEzHweWJjK8infCrnIbJFEzVP9OZ3U4P277XKq4F6pTIrlciusmfFQIcUdSMzwrLneUX
etMOeFlurTvrVF5aB0gb0EcSCrDyRGTx9vzY6PAD3gQogmnVzbWzhppb9piN1v8prtV40madGfi8
g7IFVWRBc2A1xygcuJ6VGK3VjzpW4s9BcnSKTYVCqYZZUmB0xvALmrwGd/ydnp6Wk8TuKO0mpxWT
TAGfONkAo238seoCKiTg+OajvFWAYums1VhvDkriHMLFqsBXkNCsXjNfOv+WoBzHzbUCPFBEyec2
Ito5H/lFRqgKTEWRV4Q5t0pHMNDXMjj2OehyGtnHTiJfIiForKTNDqeeEE4Rh6ZKpPaVF8EVueRH
AWajsR0M1/qpvqi/OikG34dcsUlbhCrxLbYkmSBP4qpccl8NkJKnWgTc8EKcNyaCgZbeermR3Vjh
tGdJga9n6U+g9QLN01Gv1ens+04wCIwlad0eOBjeV8vYSuluYoN8alWk7hE/PZqQfBYgQqxJuxFP
qB+BAfEnYFM6t0MdG9Y4/zM56WZqRd+5WPyf9I+UKQEeAysqPEk66ECtcP9Y6EgnjWgJAn8fn7bc
7xAA031n4yo+qCf6r99+KJElNZ2Z8pK7wIusDlENN/ku9pK6fwXoQcmOgVWbxx+xyiMoIMKN1+eo
NPpyvXVcfOEzPWbDmpohQhCkCmXd9K6W0nsKztMzDCB+BTJzJSnunyprvxc13gup99memwrBxXeK
kLFGB4yRexncFlT5IKzvoM5jR6cPuQAWDj3Ns5pkiTuR6jwlA6i2Erqhd+S1Sg+bYLkf+jaPb703
/+83DkQUbG1rWjh4DVWuMHZHBrrYC1G9Fu11mkk9CNUpBUM9A19k6dDMs0LHY5Nm0XJIDpk5qLqj
CJPtQACiN1uJzdbwtEt3TOoF2P/9hmBlUF30EbxfG4+aiXjp4vWL23rwqXYyR4YTaj4XvCQ06NFo
anEQVuwIkG/p56K9ddcb4qcjfBzbUxP++c2JFrGBW/+AHF7RdRCZ5J4nI6UlXyd+SKYJoyR59KaI
Hkzepx9O6GIBu56uMGkgQLP2CYbs59MEPplvTpmjNdgfagl4xsB4hJznuECR3o6NTIUHOIX7RQvJ
xstyzgxo7NvKWvPw3xNl2iMqiUMFb1oz1Bt+Sum3k4/EgN3K/mzM74C+e9Ub49PcXXiYWA57TzT8
VU+dC3zdkNB6DNtpEZG3ZOTLbz5F8WNUw6uWHX8ZteEPHU3Mp94SThMGJqfNA2iJ198ubmRecFhD
ht8gaqTXGKUatjJCOip2IpsAbSs11QJX9ATJvLk1BZaeV6hgrussswlBR5azuDlYLuKvNGqpATO2
u+26Ma4NehA8DctsQNGur22ChUruTjIkSBc3FHuiPkFPVwcjhQ2kV7AyiXlpaA/9MmLLIpqXinx5
WYfA21IPAP49Zp12KqMjUTwXrz0SkFR77hYYiWcJRAd9HF4AdxUoWUsY0KhtwhO/IJo9zeJs+OuS
SPRfW9s9/n3C8ILvmrWRA1+hd/7JBca3/FNyTP7KY+1FZiOZ7PaLIZ4FasbkBlGPzLxvJ8LoaA78
1mCu8vcMgPLlhE1uYd9Q0gpH7Il9egELt6lC/XtjmjzqF3l0NEvoGk/AqpheeHGGwSu47XIbQRZ6
Ar84d3kR2pImiKsGt3COF3YQN7Tg109RrV0dFf3PWVl+kewoOdR6ipXgdmaOxoYYdIVyv7FUfRF0
5l8tbt5DlARCtvM3Z3y8WUCy6eEOz8kJ4FYRlIZ311Mi4NhQYQ4Wm5DNtAIhBLhDhD1NGVfoLE1l
UvR3d97HtFY+P4vUAbfdtzleGKk5hnIp7kc3DvxXmhqjROOHmeELYfGs6rhtMLCQqfwuc8Wr0Z47
FXz6vcwOoiXgVexvfSlWJo7qD0IovrtcK9T5Jf10gYVD09tylp5aotThe1aD1aWesrJTK/re8r2l
v7p48laWWGDaWn7w76btOVrlPw0BSAdbngezH9JKSoHMqM0uauCeIyuvjchyBkWRaX634NuByn+s
MXxtyR6W6nxugQur7QLwVxHYaNuRyvxzF7niFHWX6UxOqZIfeSzB2P1zI13sSRbbJVdmgMIcBx0w
uVvdonjke55i0JXPZI3xpAidAHKIy32JYRgDNbPCx5EQANSLvFpwtNGvU8nKLilpGxcd2YLzEbT0
+ts5cm+8J/er+Zu47Au0ShzN5daS2LfGiE3wLcA20N06SMVmEQfxFNisERxLRPUm9XYcpfL6gv6Z
3kVBJz8LnVxTFJOJbC8BbgAE9L7VuYF6JnFpYWETgS/JGNVAB79+P8EWLCM6vzzw3qoaHZZMkSFQ
FB4QjD8x6rjBpcsKPShxQL/a7o9zImSv6OhlXFcufWDLUjATwi4SO314BcK++DccCXEzWdrz2Ztn
PHjDktYRO9ZvGtPHBVcXourElQByDR69r4jIFEXEbD8EPtuBhfHLbNFh0YrlojaouoiFGT7vJYaK
BFix+t/3lqacUsT7R3yR+chMfue9euvPkqczvwIyj0IG6Q9xOUZE2qR6aqiCo139lgJ0640b3KBE
w34PVpbpsBGSgvoUf3p3DXB3fnDfTVbBkKbjx1vuhN4+qrOQTk6SKzgSH/AQc7rc7BCNryDiTKSJ
g3MD9T4zlbIGNSUJ4+x+Fqfoufy5NEM9p7Hl54UbMkfTcBY3hUQNSQjKinwlp/lkavvebHwFgbAf
8391pLg98FpL1m/aLX4urqQrzgALKiPJ4k8lnJ3t8YP2iQc9m4pe10wLOc/3Kl1jVmODWIWo4+if
Ia2w9h+aqfnthtCsvYDzNo/huRQL433Xo9MCcFyu0od1CigDnWdRHNlrQxMG6Hbfo4/TUwDwTwsP
IzydR7mFIZ8W+9dkAGtwlFtrbUR8a4PLy/MnLx/q6vGXHcD+yC3JHTqKw6G9p/MNpq6ya/chmVar
hj+MJIPTnC3ldw9WXDGgA98aGEfumLYJIxO54rU4XPdCQBfK4VkDLCskyTa2xWYD7uLoRbnmkf3e
gJRkO14SP+4etiwDwTezZtPyc1jqWAoZwKCtODpeI851cG0KsbD/K4DS7EZkFept0pLi2KL+TfSt
IriCRltV5+dqyBE7vZOIzfQ3vfJrtyOY5e0tSwcg1friSriTgsf/OYke0AJhU8Gmwesw1RjqQyXz
GvUxLfUwvzID05IUojC+QI70ugihbrZ56WTgX79/vlbWnNsO6GEFvMDW7FbOxbLKVEvFjzowePlT
YLCk+jmkJxFAkteOhJpzP5MsvT8gzZcBMzxOZoAcrUqZUlStXX5tC7BA2PkJVadbaHLUK/JHrFSf
+h1v/kbncMGr827veV7xCw/neqVMiuzLMt0tarsXjDTSTOzD2V3YCYca8vHCp0GX7zNb0cG82NhI
Dul6CPvsJlcXVBQ0XQkM9bNDcOu8qPM2mrkn+qmU6HGWE44+A7FavWrKd4UX2QfJUGuDeeRzpch4
PRYYtG0GF72ZYztTRmOBzbm4p5yAKqokTpi2lURUS/betuR+z9nAKPV9XDZ8Bz4sxzXQP1ilDr6w
SfLOV6bUE73iNNde6GurrdefnCKlw15UQctESxSGhsk4smeYehdEKtfwC4F4rD+Xgiv+vH0g3c1U
zbuMyJsqAp2lngUt7KawHHIkciQevj+Ulr0JKZPWbxEDOHrM5ZEzGeGjB8t1J66/PSZ2RBAPR2Ns
7pAotaRMYnsTX3B+q8vZA3GYiibeEnpiIA2e9DxyK+pB/vbqZcQhxGBHfvScud80CG263ePf+F5R
VGBWoO09FMUyylE4jkFsP6139DFJI4vvXUEhMbi25ACRLvo8M9eKkgP07RJlznyFY4MNccTODgar
cI+GmVmdTq9yoJla1JV1UPVTd2U55683nV/k6pl5CNpqZxVpBwZBCcMVHQGLUkAb8T3Lx31336v1
cP0naEignAmlJsHEvdpzuDJ3RrvAUWlU0kL/1LGPkIH1Fq0iNuI5j6XW24tnWe3iSKZ3is5DzLia
1cXlXrnYTI4VgnpQRmB5ccGrHhy887aq3aeFWOkWzqRWx/Mfx9DT1CEOftU5tmv/MILUNPbjDdam
5LlJF0/kMtevVqsehrM4LG6GbR1BqEhz6iLDFjZlVaNDbPGc18XYQ7L3laUhQ74kafEAxqVGIo0t
/beMovknnJQR8qLL3bydNfkVguUbMincPmKTkjS2+YIKyW4WgmgVbKawJ8j7VbBdhSLHuCTATqmk
r+TgdxNu5aD8uzKFh6aNy5XvXwSf2hruVIb7i+QlaMjrRXDXTQHFgzusNx1pp2Uwcb4bOkbOiLJh
1wMZiYqFGzxd24ZjxGw2pWfVvPj4tUcQpRi+iPW/nwxprPeGgRViS/Svts8eayMva+O3eU9Sbm7B
FXit1KfOIWmtMu8al29ohHoyvmDM/VD3PS/UbEkPZqHq920MmJa7aQiCwX189dsD2vYuxC/8tOLN
ng+KoQIsubQXgMXhXIDdO8GEn60qtZB7lmSjwFMELa7qhnUrgrznhEB5pxosWr793fFu5copR95s
4oajuu82137PPrIBnFeTxMUKlIouPE0WFQZls1wtAZrleO0fp+6UpGnoADDXoDj5EWqNwi6sThNL
h+IF7FMuSWEzelUbylRN5N+kgBPxSyrPVIWEQZSuE0kPurnupsdSJteyFhhPN3iOlUS5Od9bYxdp
1OCYIZ4g0TEDzhczYpM3UW5QSxpThp5cykB4bkyfyhd0naPdj4tCK06obJIm5OpTMBvK8NGnDO8h
wD0ww4HgzDUa2fDFvkZ/y4ARV3jY7A/xrqSizBg1rLpdyx2eqeNCSIGNZs56T7JwwM3wo7gYRmWl
PKAa6LcUtBSszCqD7xc5a9rhUN1mDh50uefPHFkDl1pg0OXLs4tSfmvJZdawAtc6QimLau+L4KbA
FlHBlseDQlMaefMG2rJlOQHxVM3Ys3nJXm6QUKb4GQeoTz0gSkmHKw8GgLlDCVRt8bwkO3xvkHKn
We86P6hNM7vh610CDG2d0x6Zx0aq5S/uUC7wzmssQrKub24YizBF8DqhkjpD91x1LUvR7kf//HqQ
UzqvoCeoB79LsIRcXEaG6e0nS62ouM4SEMEZI+OhQC/g9QtRc71ttaPwnfiu9XEUi/HDd0Tm9ap8
cbg1lYM2Axkjra8VpVxepI/Cypx0mFK4R7SH5MhPUzRUcdCcgvJ5eBfVXGrw+TJXEGHWmvA5GbnL
y2J+fGOJof/GTcuBwGSg57rmv9utGH3RbfB29dKn6v5L3Tt/piysUwZzzgwQXjPw4Bwo6ZJStOgR
8BmoqZKX3fFcuAov95/2FYTqNLsLR/Qh8QSCEd/JsEER30buyS0M1xD+Z8qOVy/Yg2S5ciKzZH3+
TTQoY0hWZMadPRi6YzJ83fkJKtJW9oVg4sp7aYCwYxLkKxVXW/RZy5ln/gCvu5is1+7el3BGhVRN
5/gHPtj9EW044c32ufwW0tg3RHXWVqFqC6whSWCd42mtfSBkyG+yx4m3VNQnzlseIgzhlyfl48sz
gnpd5uvSj4DaI6x6mR2KVxhnusBBlYjcdHhmCQCDrDVGNJctYskWr31K6UZigxIplDg4P+lU6ZPG
UHvv1Y36wJWcYePhr7XtTRdSB+nqk5j+6jsi0xNx1ksfDwdukltyZo2s50kULMwDpIyFzAzvp5nz
e7y3gkwLMJvHycxgmg6rhwB3q93s6TnTOH7Fm/Z8wulSBTyNepZkPBNXCkf4CGdgdm/ScFgFJcBb
VR7MKzhbr+beJkGvZ92GsqcHX2LGlUvUqxVFRMqcB2TZtlzVW3nGaEj/6nDVURT2JYajZQVAzhno
nyH84UjULr/W4hrFdqKrHc2+MOKvsHrPGCwOxN3nfZirI4RB0LO28JNsPelwrIzNVZ2gIW3cq4pp
THUn3sy4To0BfcnDOeFI9s48w1jm+oTWcBLZtfqXOeCp8ST2Mt0mqjshIM9kPF8MdUDo/rtNvLy3
1fdTHbqScrbUcVFmriH60Wle1U529xBH9Zm5VbLs+JVtISeJ2m2xkP1bgu46Ne9L4bI5XPDxEgZ5
dJiL9z0HtV3J4ji1IsnntUi5WZd0zN7nbGR0oxrbsfvWDDMo4qfch79vm74nyy/PF/bMdIrDGyKS
DhB0IV7P9vUStf/wOMQabt3/BxQhizjJKlhrtiBj8Ryo+5dH1ENo5SNB0wfrGk40pV4Vo7+sgyTg
PMl4zAuKoHzZ7FOehvFb5S+2OavK05WNCpDartUx+d0L26GFrh5LoPwfriFoqtytnhtf0KehkbdM
Mk8SPJ4HMuDAb2Xt4dBGQ9foNqvp7OvX1aV3/9CKb8IBOw4ewfwFQdQRYJDjK70LhT3GoxHTh6Sp
HyG+4dmpXSUubZ+1ntjgJJaDt9MK/6/wiZH/0q2BpIzuzseTXnfwUbeAIBPpjDyTN7EdSt20R8ec
i5ijzC35ZHXtjzOxQLboBQLqrEKq8qzffSbwzkB5jkqDsoEyYPeqfn6IY8VM7rOaiJj1hD6GnwdC
7ub2VFlfC2Udog5yfKmsGOz6FZNQI+ETihCaaXXU0/n2V/DMccHn/XZns/+AoP1bJCuy3FrfKOTP
ieCzRDfLhuGLsbTACytTrUr/2+Dt5iXJtajCGMSBcNzHgf470ZdI4nu4VZr2faesCdiIbW8j6H2t
l/ZCnHKdfNMLs5MLSUW8HVOTIxO2Fmn+yOe4HVR9dZD45q52BkinFnRd1pqcEBZgrb3jf2dy7RnO
WxdxVeMTbbO6xSIg8EpgHEwnsuWgovF0QFwaJoncfmr+6Of49nyhF7DFNDeHgPCB0dDLdGaIbDEu
wA7bxlGkJR9tqQLzfrDQL0S1qV795y7JLhni+KDcnpXeYr8vEXr8SDjQHpYOwPscNXJkJefmX3n9
s7LkzKN8MtfoL4FQA+B5qEeaNR2ZaP0fKA16nGlKVYcvMRnASy8xg9Ob5+tZ/140wqKKYLl/ubZD
jf7YPt/NzRcGviCl8r62TGI1mY290JcmZyalWjttEj88dM3CXAg2HBCmUcP2t+kkhzSMz3cjbzCH
QAtoUsx+byvwa7KYunzfhJGkQcgOkRL66UCDvbuqhQRfZ+Aotac2+T49y+VlUiYc/aii17mDh6ZP
APaSWsNv7fQdx7vaEoMriMxjj50xz6BstVQH6oDNsh1SwLiCWzy4oz2YZCXe5ynVsnGpSgVeppRZ
r92lixDm4iSFhwZobCeBtoYC0Ev7ApgP3p/5H8Eh4T+35fyqXd29dN4fYAnzFYZva6fDh9JYK5hn
P8LPxOO5nKbE5BwD410oP5BzSexFVvyIYzgH/18rPczcxko4wRtk3yPrMq40GGEqNWDXtGCCHPeI
PEhr6wiTv4B+Q+iZn9JzxDzQE8XQe5bhpbkeEEsSa5s++rBfJ2/Ku8ZgIDGv/4u7MuDbkOFyaJiq
V6RwyGGFaYPlryD5xclCCFwFPVTvGudhPJLgSiefdgvkVcKVsQ9k36b02TcCSu9LkHO1f3RKIbPW
1Hmsar/z8ADQffFFGatD8+Am+pSW43/ImXliV79oP1tlXZo8KAyAGgXJ450Eoftb8r9Uis8L2MgJ
8JkT4SF7RltcAkxM6wzg2snL1AaRxiBblHUxWDRpFkBku845bgbiqxmb/Ns19UQxvW69Px9w+DF6
YuPfaisxG6DpT9jrWiv8whjTJyUqrONTAKJzYv1Gat8wvHwaxXTWo7v4mu4STmnOM9GAmJwqXV5K
cY8D0q4BHnIyuDUz5XpbQMesidDe7h07t6vUpDenIJBLvjBkGPSBChdng/wOxlPuQ7shMNvf+wwU
8HeCz4go/jtgF7Gby8cLXJ1aj3Dl98bkaOfq84iBIdZ3GUlDPpOSl4AZLPTVg5SyShiE0YwwOcLe
BNcRTs/JSg1SiF5XVqbLidYks02XpeaQWXuq0oHXNxZegCfEd3ffS3q/ujB5OXffPVTMJqz1il9t
mluwlpBew4/LvkCK/cMOcpp0zFCMGF4H5YVfqEIEg/8CbDqEaYfBVW6rdDhlsFGnfkOFTdP77Bnc
/0nuz7EMI7VX7dHdbrq2j0I+lOxc+8sytNzydUZs+VlErBx7ILEwZqIQRcVBHP/E6/9UIdJJvSIi
sKC+FZM1zJL21+uCMTVHr1cr5JF5fUTkBbodqpccQ2Sjc3dzssg3R0JVPgTvySY6tUr4vCIZpKeh
NpKXIMMqxNLtk3/emXPVHesiORrdg+VO+wLBzvwX8/aWIPzVklz099oBVQjC5KUUTMyh2t39Cr8u
9iVenRLdebOzy+WZAPRc26rPRD9vKV1iaKErIjgL6wVaeKVY3N+cXio/tWlaY4y428uUIGVsDh8W
kRNEUM7fJTtc5btIDr3H6fXr14+Be7zYrUEVDWDtRDaHaeap62bI+dGdCEQRjkpmrdmJBgBtWw4I
p8dvW2T9fe2gRghHgHMeJZJPdPfKIV5WxIGKkJdNIRCPcizv/tTRp/EqoSSdmPefTmXINrL9FhrC
4gcBTJN6Zd65N0i62AoCdHVwO+nZeGsho6tkR5+xWlW4PDjkAFHjlZl+WPev7q/B1UTbnVPNpmwk
IdXk1U9uFdzICWGmyHQO/C8z6A/jGibjVxho/z/pKkWWWYEz/y/fZF/hdOiEy3TgzLytaT3mhwr9
JvVGVdezcBpA+tM+YvTlZgKAa5h7H0lSvDdENKVKKrNdpMn19xC0tA9Xwb1h8gEYP8L/0DgvpQWp
MVntxi/hw36m8kV9KjXrbJPJV9qDiPE+Q6xHZenIz12U8yyJZUGxcvO/QCRDctSyO5kEkH0Fz8Vk
NZ/9Nm6Yp48f9004ktsPi9RI9/9DmANXGN/2Kbe93iBfQ2SXz06nON7joCbGrzd7yX7r5zGsZMF3
fWmVJK0JRa5vCjDREy1zkdXg9uJsAHX6eHIxZ/FufNZX8ZCLS8zOQ6XN6GlxmTCNGUPn6uzZXS3R
cthaIMp6JejGE6KQfoZWkIASIxTIc5RqjBgFo3sMvygTd4Fa90m/1gv8L+t/3arRmnXBXOdcQlt2
03dXyJbDk2R93Lmt2JngOamdbmP4JJ4I1ui1iz3dfxtnxV4iA22hj5orP4PyhnUlAX+dhp6r8Rm2
/mo7lAOWmHyywArwbxlnwBrRHAeg3ooz/1rzvB1DT3YFZLMfHzlmSCWyB7cakLzvUsdSi8vG9j4S
YvSXJynDX4r0Ay6posF12fYXqOpw9GuW1hKWNVMW4PrH4nd2cA3mfVvlJZ368dTI8hlNatqW2ODw
4D7CNrzPKeIyQHny2WtBNDeO0yMvCpUL9DVPHtwWzyQq6fQPio1FZ6XVXKbMrdS7OX2rQveq8tme
I2taOfm4s7Op/HG0VWfPoZa4NMxhsaVmskhKvQ+rkwM6j/zsA/fbvwcLhAIELJ4ic/GTFsyoj66/
NqZlZd8YDRro2/mZ6gFZwkO7LOXV8rEf8lpQcBKUUkDbtT0OloETdH6HS7AN/TShG4PnDZbpfRUY
S2vTW+lb4JizE4NllTkg5JNRIde+O7gdKhE1eaOiDhLaCGZ6CSvyt5rtlncHIf6HzySmkQfg039H
Uq8oV8DaEdC9665elkQvIcoHslzcKRdax2ei/CEQOEJnmMlJUtLPeHCovfJhUnPg4/s0BEZ1eByV
gELS+EEMAU5jy7IcDZfz6h5zmuTkU+5BPznkxWDIP1CgQp+KTENhFdb9T9YAxgibZtX360WXt1sN
cbaej4TTFvWBJ4Ss2rcz8TjGAhoIpLiUl/FTUejosOTV/QmSvSVOr6vIXrTAODM95Pjgijx0WYyI
ZDT611j+kNK40vd1aHHKk6kIZe3DArm4Y/PeL0F9WvAJwKW4gMv9IgEy1torywREvRjsgNcXcKC2
zYr3bji0N/tK/+ytj1KUgToeD/DUSA6SACEpln1eJlXk4KddCWPmtYbsEad0PbJFAenvzMOZtgUE
/tDB98PR/41Q+N0LEaz4IC58PrHpCCbDFz493UocOi8gI5ejGPhflttvuNgDzuB+L0APvhIZrzTn
Ir758B5jhHojdgnGqaJd1Xhvuqem0yOZRGWZDDMixLvgLtOcM3o/ucY7IWrL2NKIPA+XZCMNfFvg
Lh1SViKCUQ5aw2tOftzZjOiNWq+2V+2VUegjSTqW78ls/gcy2btpZ6hjMWPrJnvTRAp6XOKJg+p3
uMEi16V8sCWbEoQ3FxwR2ZtrV53nQRX8mmv+I8AdeHadZiaPQpSGWYfyBkth2RRmxJDbs8WZpHXe
lA2mpdaArIQ90H76MLtrXpsopZ3EcWoAdvEPY0XMRPBDNojstyJDmz/h6PaUBwgNR8JJpoNmO7m2
Es3jVlwwr1GZXZ6ENn+0xof3RKaHiOZK3lBBgtTbop0ErbU23yaY3wSzFpFptJm6A3QsfyWMu1Em
sNX9ze2QL9aiyHjlZ3rtm3PXKovhQjv5e0ImwxLhYIRnBgRMO3m248Ci5Nr77A2pp3w4UjJSyI6d
NrTjHkWMeNUxYjaVhUuu0QjubdX9LlqH3HfjE8br5bvkD9lSQyOzBGcdxDCiUVaj6GaQZC23kiem
++0aUHNqq5BYC50P5shcxUgyZn5/owyNqsNasiW+e/LuLQrjDn/YqTKbFvJX3MPVGvPsTaN3k7Pa
hrlZL7PKXWjZ56BhCZBQWzRciZc1y2KPYD4oqL167fTpGuNVsMdpiA61gxsP21WwLuqfu+ZOj3ap
PkjnRcdac/2gPNHxOd1v1eh66sj2F2W10SW73PG0zDKUDuqX4WEb7y6wUQZ0gvR0S9TFcbITHRQ4
SuWQFJWGBn0WsNqHZQfyLI87dWxSOJfYdDp2w0zg6tpiGY2Cl93ssMnP+IS/9o3gjBdnIM5WBkWM
+WbV0T/60HfEugNDVKZMxDeBmhcAKlIvSxn4MMTB3QW48TPzx5zgqn2cXRIzyrdz7OvnFOwx7Gwj
x1zB9ccv2vDOjzkqX3Z0LaZahDwt1TuvdFqsJYLHIvXqxRj6cgBEmcyr1QGvm4FyCViPUKBu76Oz
a2RiTM1g/Oly10vWoT2t/guHqjVxvDWtR5MzgY6rceRffmJ292rry8jNj+N5nsjW7unEGjT8i0Y+
h11gwI37BG3l94jm91icNl5F8QeqsFKXA7/5g1FHyrtpA7SeRvXGVB8xGr7KLYEP1MLIJUjLTMcf
yPi+d/QyVUAGu6G0CjOfKclSwUWzC+iIglfFOPUtJNZ1xs6YQPCtrGeuIW0yny85cPVOGrJLx6eh
121YkaaODdsojUK9KNEM3nGPFJl6qFrdXV9ma5m9Qh88NGT2hJJQT3sjLWZ++eEnbxb2FlNDpU8D
XSQ3rlo4FybHBHi5zxzv4RmYAaOQDi8Bi6mw/CMkLCoeVNY+Npjcu2B4h0L5z7sMqd0shc+xI9A0
jqDWmMufOepDlnAWAVivYX7VDMqudWdJ35iCh7P8dgIhaVLUpYkqeRTrAoUVhTaVDtzOJiLlQf4c
2DQBCNhkOGiiun12QeOhXrB5+ksOlRMt5sk/bN+3NrgvQLbhguM8kiQxP54wdq7hW/hdw4aZsgR5
sYyTo53hbFvUW8eGqJxQctP1bwnhQtzJPXS/Ei1xifqbO/uZZ97dxjk7qsP4k++6gdjmpMTJM7q1
Oxkl+i+CgkzZsHxzXFh4rFTB5xWYNQyvjctKNxq+/UWJ86pT9M+XmjTIzYSu9N6ELs/KCAmBgqvh
BaPnhmScd/aPf4n5nnjW7Qz0+LeJK2K7fzB7BVKGzqGmQw7bGOBt//JIYQvh796DHUlTbg5fBM8R
O+Av9G0y0ecZPqYOd8oz7/nRIpSIQ/vzfk2pd2qhkF0EDByv6fFabyazVctPq0lGMBJj30Ob6qhX
8O7xUdYm+6cFVlXm2T6o+g9JIFaem8cMykMaf4uTuL/o8TAhFAy0LV5dPPlPmi/VX+DKYvWG6MRY
2hgDWHrK4jvcSYQ+5P0GROA8kqkpjtuk1y/uXccmXFbeWd4HJkJ5mH3iDQDKOrRwzzWj/AeRQL+u
lAVEsb6No6kzI1goHX1FKExes3YPD4aDQab3dBq3F7lAkg1IXmTqgq5EhhgkRJq/rppnom2/uLYP
DfEDSRQn/66RbUtfo+IvGPGQun8tiH1Mxug+q0SeC8a57/BfIvTH7nOY0ysAdQaJ7Nt4C202nPfL
tXiXoPNlI2+Jfc5JRytnoB7nQp+FhQZK6Fu7IyHJrk6YQy7hQ/k/y74VkUEnuh0U5ZR7B9wpTgpW
3+toIblJKGZtD16O1ybljhF/kxA6kQfWTOq7M2R7H3o496CaiwIqYIZo2NOhutaPzR634OukmTSb
tlDCUQfVKyQ4IzwCUYfrc4tGfLYk/a9F3j41lzvLI9SY5DcF9/LCaOY1rV74q1wyUtdbnK5ARrNA
ErYAYtB6VQCKMEB8iLMSnwaqQN3CWNkoico4RPs13flfvIiJFhsFiM5CgGFLYIZDqArVrT0Wg6GZ
UEbzpHMNTU8AdVmWZvYr0LkBYJWke6dU3WuersGrFRWMhXVVZ+Gk0D+PrLNsmz4auunX28yRB+AR
Rrqd3QRGJ/KOdwmzNlG+T803VRal39RdBQLPYuRqmVeqpTZai5DlMz/Qh+Bf40wbkGYqf+DOB86y
uFMCtovfWA+0N0X6lL/OXStl4al+XWuRM4Pjpqb4avDwhe1/YWZCMmZ+QDiIprKKqc5Ev8u6yvGV
aNe1VFTjv7jxTBwgYvbXYm99iqsmF9ICyfEhaL/Urh5pFAE6rYipubx06fy8SXMdIOEhCWl8Nzs1
YDM8Bv3eiDlPtHjj1j7LFSgYhY1j8guFttAgOwZlfajjn63KTY1nPZEEO1BRfrjdUGqkgw74XHCQ
e7fVpUhgidWPl6RARqZ5PXfc6k2H2EwcBv6By0b+gCFNE2L1z5aJXi3RDUqdfcV8pp8+u7SlyoLp
G1yHkeABMeJgMw5eVxw+is4Wpauv9HFX6OPZWOBhlTzGydMCKF0EgPhbGXMZil3A/zVd6hMqJKp0
f4JxQpVgkl0bwN5c0vsbFg3GhLIMH3wdT/U5Io1SvldbIqdnhYYGFJ38skRcRzlBJllo5+DsmJ/d
BlHStqk8EM9L2CcKaRFobKhXGpu11CX4VxG/C9QTRiXaWEbgxNLCw9ZOjdYse0P03rmT5/sVJXzx
y/AEQz+NdwDWw9D0dQ/3wIQR5gPBhT/9KHya1c4r0EjKjkVc+/Kfdtz0h8CM3CuK1TebxN9bk8J4
hzLRZ7IPMx6MEez5D40UwSi5br5HsB3xneX7MMXJE1tM46IOMa9IVIhQv3Ci8frW6QKethTwwPNL
ERAs7ITfhG48ArB4IrLIaQfXjzjgBxcROdJTpd2vixoGd/45dQMqBQdXFeAy9nymB5g5MhAQcLGU
IxJTZCe+9Prx+4N04EuzVUYj0kwIKnWr41KAnxnCmeTplpsjfJxDPtodtEyuVMM2CVa63UlxG6jW
oOlySC3jsuJg0X8Xn7GN5RsAVfa6Jo1V4HGFzM/yFz5n9dwRhzU4XTMR+XowWaCHp9HYVgciLTeP
MtWmOGv5ojjG4MErq8EWDb4XXB+z/1+RhbQhGV93xaeQuZvkmsXg/Ro727zG2Gk7aQFmMQJZjK3b
wiUet6QEecPqqQLDCBkooVoC6vcdBye/rFRHfL/cM6fZvHGY9xe5W1OXnwxW8IZNO/vfLtb8WtQj
l/1HpDyfOxMzv4W0gmGcC0dyj5wKiajmQpSG0MZWGx5lan2EEWtMW2fU8k8esSFNscorqQXoKGnQ
Qrmplp1nRilcY0lhr1WiidrwVEl/JJXthbZg1cGTgjLHD+0ezZYfPlt4EwSKZNgnij99pY03hX09
fIXePmDS5QUjnoXvXu4z5Jkub9r0UtbNl7okXhTmBCKaEWngSBWSoGL28vRkvxnhZ6gRaRBzhWrS
QE9HjD215nflWbhZLOC3NIVNN+Cp09RazlxnvK8D8/LlPXoLcPB1J3YbXpYcIx2j3xqhjLF20DzV
+KusCvQWr6jvkOT4W68xv9tTy1Ec4fTui6Q9V4egjWujhx7FVORaKg6IrPx0xhFaC9KveUifGi/0
r9V9ZuIA01Kk1bzjgKVuGttfQxW9ukqzwqsAs+uzOnx5ot7/PX2kN7sXPWZ7ktRgoCtJt1ejAGaC
Tk9XqqYUjZDIr7Ci8gOjakT33baNjjYe7nL0XHQhXjJvEk7png2Oc8+sX8wQco1qg7GKa3725tb2
Ker5clclWOl3hzDWkyZxU2sDSgM5HhrcI4ONFhhc50sgHrpA5bQUMU3ptz3eNgGJyeuTzXRXdzvv
aXVBChlO1o9mGK2w3IAIft90fRaDniPgfmE02vKswWRXVL23dcGKbRQW5pVaSuLMYpS68UCmfdYi
bO5nFBQLZZl5qICAOlM77qP/U3tQ1D3ggXTBXxXqoCqmrYV+7kxGzFZl+Q0ES7hoKn+bVPyBIj2L
tuWuGnjV21IWXCxLEb4v77Lm84eqfo0EgovjQdUn/24yGDV3/8jtCvd9Tpkzw0CDuxLhKeUQfwxb
fyVyhzpevu0vd07WzzeLC6GOkeU8VkSe+ZZZPi8AkCLcOibRaPhm9k6/8dFPMNdzmPMpm5RzXkxf
Z/auq0nwUS7HvEx/J5OAemUGG3X05OHHmgUBqHSJ3JYmjQT0Pbi/W5ecGz1IIW1VsUf7Mt7Hz44c
jrKEs5WuHYXvIPe+pNyZYi7jlLB7ZRUm9KOImoDf6FhyVMT6C7v93lGVX7OFSA6bpx7gJ7qx7JBC
9OPUGSwxFJbd3CiModf3teZrrv20S/vZcVn6r3OHWZL/gYkT+WQI5H6vVs3cVODYGUJRM0C8gige
FEaOCYqRc57pmJs7h6EaqMdf2ZpZm60wp8orywc3qriqQP/ASjCVXdrE3KJrpUn7vb8wCkuJTIr+
T5Cmc3xeCalOkoqb5rJly0dGLcCX5JF5RGyrdePPkeAEgv14V5n0PwmY7Zc7OM4MxWsQkTZpUDS2
pPRN1GHkFnc7Xt2XzRXVf8k11P+V4k7FsPGiff55lmX4C4el4YrCI7MVBBqZSd3sYZy0lzgYDNNL
1sNGKsEhxvsbooOfixCJYQ1VwqWLxaZEL2HkInYce7M6L4vWTOPZxXMQ662I/86exgjESbhZEY58
p1aHyAxb1uvRC7JmVDkIC4/STqMTi3wXgwuX5lkaolfqIg7JZrpCZ1SNzOCIukaVudnx6VWyD3YU
Dt/0eu0JjdSwGqo2FE8BEGIQLTxdpZIOYLlzBNVDD12S++Vjj0zoq6/AUoj7X4K1SDdYlWMsdKuB
7vEzoEeLm7xHEa8MOPoogxxhi+0pF8BjdY3YZBZxuKYhWpW0k1sU/TfuCHgzN/X9bRy1Qq+KpHX9
NOZe+AuLYO0boC0HCMuC8lsRt9KshrKH/abLmICrsKeYai5CKUXc+2/HzRobsr09BeV12GebSQ9/
F/Uwk1im/0JpImfNb85r/ot1lYDgk82xcJgqmL9cHgrtbBrIBG7ZcDtTawXISlGvvVH1tuNNs3EY
9vnO3CD+Hwyh7oRtWA6V73aZFHmuqVm5hQLgk3mF6mRzWVcNoNMsXJ/6T+47kA0h9dy60bmNTpC1
fgJyJA7ikQMOJd5q4AQrgWOp/SzV+AbzG4VWl8TeaJ2lD08KalOFYQOMcFcLiKMMf0PVVrth1KQb
dOzYyN3kvqn6kbi3IIg+GulCqzAiCpocdxMTpW+mEnPTmT1BQiEyxyElx3yAzH8O/wCISzf5x75A
+Cc6fgoHAXBixKgn4sYKE/nfcKqhK94SjwzJJEdgqHdUv/DDPeLpYrGkjHHJAtQ/NdB180MJ4kEt
jdKRMFvM3wFyIxTIhKFuFCnXKBZDmxEs0PbvkR+5OzhxuFvCbJptZGW/WbXlLP27Qj7jc2967U2L
ZiUws4EjPxY4B+4c/dzvTftpwYqjiI4TjpUk1FYAQLkCMGwbqjf0D8Z8IpncIrVEBnjUkq1s1Nj5
1tW55cVqBMPg6mgWpgNdoSExDLrVfi054ObAwUbbgTYMYJk1rouk+VaIRsNZjU+4hM73r4uJJVH1
YdkyENr7uPnd1vKwGTiXJUudW+gDwAuHsoyOujfa37NwCkyJrbd8FrURM+V6+Wah+1tHspO61lNf
KOyx7xiqRBZlheDdAkCyTWEW8vs7khd26KVcue0KmJ0X8i5ysGI1FA6W2P1GHDGlL4KALQ7o10Sb
EPaXWdLRvWIb9zPb3XeFQeHuxYZodWPbTUxI+2/7KjAMlstdfSMbS1VLo+Fd8tVHDMR++qZ5G9al
2smbu0AQKMjAYosu0kKdX1kIrxQmS5SkKb29ZAH6Xu07nnbsKgTSeA7nGGw7/9eTnFp2POl9DPdb
OfaDvH3vQ2YPABI9mL0J1sAJYntcnJB6WA5KLh47phmzdyJidNq2SpJ2jmeIq2ZU/yhyTDhoV89W
kGoSjnjg1i8MsioJVSRPfPvTr7wAHJB/MUFhbLdhpePvKAiY4jMmXrYKJEyjna+NWRyc4n1S2aKQ
UBtyMsC8KQp/awRLObSIRD+sJGAFeuv1usM/227gOTMVrIZ8SnKGkeSA7/1K13M48EgmtUGzNdyG
XlF2/d2tojkR70mGocvQU93ysXNn4Sz20Oybezong6QGMc87W3IA3oSb0JWbi8WzkCb+vxdXpGQ/
/nGSJVLmAPPur9/7IPMBek7y0LqlWO2y8eyN8ZPJeF+URx0eBUE2fE06SKX9X2xkUUWWuVlsY+iI
Gqo7XQwBRj2sUJka2v0MPKLivMV6lrVJkDBkPTrNzwKF09rHoVtKTaSxa7enAGFSQO9epd5g0HcH
NtAzsf8z22skrWOhowruOv//a+lrzi3aLVAJeNdM0mzwMsvgodsUE5NZ4u0nfcyE+dNUWpmodB9W
ghCTMw6CXPo+blViFQv7zRK7e5JePUK6HwdZcds/JR6ZwE1ne+v71co9ngUON0h+4Ln0gQBjcJfh
GnyhPSznSL+O2CCuVHm/5PnkLJv18Tc9szRp1gWFTlJjxWgf+fflIxlEuoEKdXXCAxdEPQR7LIwy
ksYrAfWO0bM3qQQs31RuLoPKcpwacWT6esxeZOcSIZCbpX28V03F1Eor3Eu60xGkzFdC5Jbwz+BW
Uf6pDs+s1xu0AlhufrQ9GVuejRmCBdYt8FVRsCaacz4vLEd5ikg01RwsXntXAR46R9hVxnn667VP
ptzCH/C608ioxkiPUqyh3KQmfkxn7hMJqtQ2Who66omwrI2yEMDHfd0HDRykVbk2tCgFOVs7B8uX
zEgjaxu8MFotHKMNn7IQpp5yjUiHaa0HXlnxijtBdHawQIoHfmNj/bNAQAsKXvvdCky/Y8vr5soV
jmXDFfb3wUTMl3tgxx91oZHDzYzSeoJDPBdJGpROdiWvQ5Pnl0j5bX6+nbosTZo2tqJJTYKDG+5C
R7401skQHkfvt7IVDR+bSywjkcx831VceDl3legzCxWysNJvvoQVF52t5zyWNrbEh0+/N47SEHqW
cbZWvnZNYFg1IZ9/R4vBFTAHl2/aIw8kqUz3evcT0RJp2+F+lspB+PFO1hwsPI+xpLf1d5G8hCke
AmFlh8QG4uXpuy34uINoi0wfsU8D/UZ1IMUlkcc6hVTbEghqw3dXjb1iNTmcGMqsCLIUa26OS8UO
GkYERQSrlUAqfBKc+nybQ/7ktzJIWPCRF6mW7ISMrG9DtDuY/RqKVFDlw09YIKVqltC2HeUdjeZ3
xMH5xME2rnzgyV6Pd+KRDt5qP42Hrkmpg1qgVBgmMH01LoSpXn9wtuNg9gXLiM1oi7Iw3Zn/ejNx
LgPVnL6lvLVy9Hbzbyx83t29ZvFtlKym0GSuFf++8f7tVG/r2FaSLKXbSDS0WOZwKr0pXN75q/am
0Y+sqqVXVUjuZUZt9zvGmJg6aD10XEDdEQmqF7G0hOOsBee744JUwsJwRUFdFnn+lSx12eLuJ3Or
FOOYWLNLGbZeIVUkwvP6702h5FLQI/he4y08FtlRxMmm7rB2m8Rpj9nnSf8qCDHKZSs/iCXF5Iif
gYKiKkQ/7zMS6oBFZBHDuJ/GQXeyJLe3nauY9kQagcRaflZuRbTQR85r8MyAq0UlKF8jcmzDF4pp
HTvUg+JVL1LJjmBtwFihaeMBeIF4HHj5vpxFQN/0gkpeP3IZU1FW+BABTrMU9XEVPTLsYnVTOZ3v
ewTK/1/Gm1Y3ovz+G2C0+LKUUPoyIDsgidpiRbEfu9SBFSPFdFEE5FBySrl2dTX2f9GxJRcdvnAm
c2UcyuyVcQicz1bVMne9RIXwpBtHOax8dgWNqqhRHYGwWkOs49bgTugyvNPsp7+5ah/WRMt4HXHu
cEYzWV25N4lyvUzMTTT27326Qb68yKKThg6h7xP2iv1Tb7PsgVmltHX+W7SZI87ny3rb4DS6tm81
XW/3OcP5s/0MikQrKNDKk1N9NaTlpoCeCkmYzJI9Dxxvq2SLPExiUSDEmrLoy5DinjlcHbqiyoxL
pb/LnT4HU+DfczxcKWGFvfhdHHekD/fbvNssrf/WQ19EVIqTN0OV6dm2wQfULhj4RReCfZ9rWyuc
0PbuDHFeHj6hlgkZQyLuHphO1xVKQMIkuebRvQM/hPNmXMhPwoJFl88MMxXb7xpL9J1Y9mNSLcxs
OOj2/8NGzlmCjBBhmgiI3X61TMFmrocF/T8BFKD5Bn1iDbZvTHCXHhxW/4RO8DrQBLYDeyXqJSbP
Yc6pA2TFhFKgRF0tuGPtoN8APtiWPqFrSjN0/Acryp6F2xytR7MGhIx0F1AI9ukYaE6TTZrrnW7m
HD1W9eXEmGGJ2N9Ouh1Q1BRBxHb76sKE/cwLIID0WQ+w/yIEXi64xs6uoPaTO9QUrzJ49PTbvpEk
nLNOcPWX+EZ+8G7d3ZWnexvq0xKyfvFrYG31P5tYoTdk1R0yXTfgRTqeT/CxgpvDPevXxLLurnvg
/jueL35LqdKr7e3alrhiuj2DNoI/PPqFTceIhm0mwIjLVKHR6ek33EsVp2I9GI60/LzuVe3uo1uR
4We3F1XFSNqPU3KRwDc8HQnzdkIy7eGBdG6ucDUBlsv4ybb7JMjzbhlhNEgXl5hYmYRu3ljkBcRY
+/qQzHM+JXI9VK9tKWmWs10eEKe0k1yhM8HDI5s/qrCOlBDx4LepYWPDrwVO3XvOzvj5vmr8x7Ii
+hdDJ2vvgfm9coTfptiJkbuLaVTt++ZIFCIFBSRsMcAV3F2gckx7mO6Phab5lwyXhKtqgrhjQ0XI
oFlHkjzVI099EJLqzzeep4hDcsWi4YT3415DohoRH3f0HJ5XaEawnVdFicT3fjmpbpeT8M+K/w8S
7X+yJ37Ob9v1HL3GdhZSJ9ZTu4Hj8bfUFtbdiRSD+RnqHXNXQN7PMGD6xCvrE5MF5C8CT0uQ1ALL
ZwGAjMcVhdaruHe3dkAZxDiW2kuiIDCteFJnlFCLHO4JWOCw29uotge4QiktLxAR2SidbMxgOKld
1aMUVEF3g2k3qHkoF3Pv3rRsnSfhe6R+MIvYL55FBw/EnCPbTseX2AwSJSda8IwC33GDt7r1xyTS
oXWFN3/DvP+dn17KD5kyJx4UlJXLwJr1vSe7MZNmGTXXn6+vrsL/iM7GWlCFRUM2NE7M2lyMzrC5
t0PSRKnhc4KqgVw0tDvY+uITe8f8Y0CXARvXAhlltEMiPArE90ukwjdY3OXpM9kjUtzY15z0t+x1
I9gXnovzKrhBcEYi2bVXxcYxjzas7PNAbbKpaI3hcM8Pku/XsK8WpRK8kPJn7AmQUeBtglkmGJhN
7UKsAVsWvOit0oSsnA0AE8f7VZyyaS6XZQeL63nu0uoYyLC6kWmisvGjByTSlfB8EkysJcX0wnY0
n9cqFhCXMzgDejwYWOCA29UMGZKpxfEapqrJaJxKREFGYUStYaF5nMGa77VpPFDT0eR94xmbdvV1
na2vyVwYE16BOBimN9C8Oo63I68NsMBemX4u8yH2h1KWFij8i/eaJGUEXqwKmfxk6wKU3luiFeFn
WjZHNhBXMqUVFbDdrEEzRNXb3ILbYwxSw7HpZ5ueECfI2Dk3JE84OHAf/7T4d+HRBRmcYME0+Hsb
Ck8MCYK86WVp1yydqkhKpwaFIihOFZqdDNtTq/tPW/mPWQkqAXSZJ4ILpIpC6XOyprHSfBPNQhWk
rye7vtRCJ98QngUos8lbXh4aGRf3aV82WnIK0zbYkHYUQMOwkEGZSQF2vk4v0CFo2ZxtQPX2p6HJ
Fw7Z3QIpSApsds6MBFJlWmEdcxfPoamATp5ii7ubtx3czFRejqNsUla6/DI3hL1J/UxkJtMT+vDk
3fUTbtc6891sCbljq3QCoeitzhHoIThosToMJevx6eV30/1tnKyZGFsKUHl77g4Ia+MWFILIK7Bd
PBiyL0JqBHghWU/LWwGc9DPdLZSeKr1Sf6YXdOWMODf92v/MWtA4K6cWtK65M97VwYnoYTYo1DxN
l627a7txEUqmy0/Pdb85/Hi2Bwp1sKsdGA6rr8uJpspdtzZSN4StnZrJMP+BLKVcDSolT4+hYIc3
86j/rd9pECDyskz99atAE+TVnRBjglmzp4ixAh1EpvmfTYfV6LrOMLHria00MQu1dJFfpSL0FOIm
LrnWdj/XNhbGDblmMTnG8a/ZzZKZR80kxh7Gz6TcyOivMKT9UrsXm9GcdgSu6UFGviv8c1IBulRC
PdCot/novyPm0eR2bjQtHPqJYJiLtCXeX4ui9aMCaEOQBgWOPeWZwF1Z72tJUtG8XeQq6SYaLEcc
KetQL50HauwWkc0o8AZ5UBVFgr0BURLIxBTXcBz/Aalpar1A4YbSrA14X+sREmh0VQ3uYtsBY4Ai
uxB51IzT20yEXYTivc3wiwMIDD1CtEgvCM9W0fEs9ilNc896/b/SWRGFCdU3VOqU2eSDFuX54CVQ
Bkp3JXLXYtaTeOtAJW4MRAW9l2i3ww1h8etk6MHLLHpNh0qb2gsRb2H90nrNcm4dTfl6y485r15S
sM+jtwV9mCkeIFI5O4P/SKrjGBXj+ip9mEAHkBJqpccY3ox/Vo+++G240b5XsfDsYz6g0fKChKi5
u02pzuYOfENpell5c7DwELTQINCyYsZ54CvdIWNdLb10dpZAarQAuP3s0NVKmRgRxl2LiPJkyjag
Wimj5oC1aDP/KGnoGSjyetz7Vx+hYzqd7n42/wzlva457QZP/z+88VNvpsLyG7mHMf8Ar8eivVMv
gWSWCXYxtMQ0ufexnwaUtL5K3wfwXmaIrKnbKq03fY+CKl6QYnYMJFx0MLYU6Sd5uRC7AqX/HUdN
7PV/RI1a1Gf5EGVVwo2CXeR5UVL7oR2GBTt0S/YTiZ+BbSjk2nLP0BuHoML3pr01Ur6p3tzK+h6N
oTM5/F77je7YNpw7KJwIiowPxTz1l9xHI3miPoaKUJcmg6s0TJbm49q1jqjAb/1G17iZfc+MbUFD
nOv948BWmYNxLKAzg0L/s17sgSQZqI6y+g28PndRr4G9JJreFRQlFUTqPYBxosOo0Exd0FDk0B14
34z04HhvvKADZi/RvdsC1T7RlkASqgSijvTFhhI85S9WYNqz2GRvd27B3yBt2ZSE7weOOH5nNLqQ
iNY4v172jij5VS3IdtoQZv7604w6OjUbaojF9L2E6+WF2lMBYtQMO2V2ql+Vt2rA3U+HpcJA8Qeg
60zFjLSMUgbocoZRr4IXmghiEJiaRh5TIC4orqVBt3F4ZXVqS1x0EdUPaPeZmZ0gFYrb4BNrCiQW
Qr/a5kaX7tJ5WORmqGrkNbqfNsN8WESnOOuC1IU6zHQzjRSImBJeKfCDNyfOii4zqXtoYaGmWMTx
NgMtwQ0431ZGy0xUZb0wAYG9K97KHEGUo3Z0e8sbbLV0VOTc1E4k50P767XRVmwz8crtDjRjMeE0
5Ulzcp1nMxWsbCl35qXmfyqCzvW1ZpcWBsjpp1ixt0JfMNak+Yy1pvoMjTo5K4ovr8p1phhrlI2W
8ZNHBSgNJPaxsPd/N/YVBdM2KqZfgiwvMpRj1k75H7OkEL8MNlUKN22/1oirEywqqIPm5PhjAYpE
/vz1DHRblvOqvkXUoVITzyRAsOgkcJjqxBKWfsrvyCyaaFK8nQyNQXPOHmZaY0zhWdMCkIFDv/d3
HpGQaI0vC3c1pUPb5x+UX8ccav/dl6ejCsb3vN3aQlQ7lOTzy/YR1KzuyeG3R/eBHFycqgv5p42J
8j9IZQAgRT4HwrU5dZtmvUByAIt8DYRm8Ztun4iZiZJer2RjoTMBdnP9/l6ohP7DDkjXMwo3xXwY
oClnoF2OTJmaqiP+Jo7mI509mG04Tlyw6XPiQKHtQm8SqGWyUwloc+OWuw+qI5TGlWuvMMmiBmWb
aCBpJjHZfIjw8bsyNgglPSIgCemUzWY7YnNwrVV4Dd3WUckU0njtxm6UB0s4X/7Y8T2AhFPi+AXW
uz//PUUwDtlcwLk8yRhLNplH6UGVCUd7qCHKQ4CsHYU3nwZwj34ongnoNAet//mnP25h2/Q7oCIL
f5USVJDMdWufjj/Feeb+bPJvItBWzqbkT1+gZa5QEmfHjQzcPCRmjAPxfY6HiOHJ042Y8BGj3Juy
ZAc7uyk/eEv63LnLnB6+4nKCGLmXJSvNZSpJ/lnvM5/Xlr6soTZTXFS8xmoGoeBDCGzqFTFl0vky
774KpFxsTz8uovdb1uFNhw6uSzLI7RbGDSif9cbposUJAmfpHLBC8M9xLxR7kKg2mYAtIlXGlClJ
sD9uxxEQR2JclymhxEabuM3wOIqVqKSyc95Os04w018BW2BJcNN691MaPpmKLILrTohOVnFBbvY7
e2OwCGRLle22MU9jXK1UilbCYJjRDaZ3MsBJoXA7fLafIOMPLuCiDat2d6LHq2LJJSxHZGCWES4b
LuPCxBDS00wgJCM154HcrcmnPrjwZnj/FE0BL/dRw5ONkDqAwVQBoJq5zLWBuTY7ZW7bb52ZaKIz
kyChk+osgueONDaJa8b5Te2m0qpdQ3/2wnVDurGUOpbkeZTfjsUNv6s/IoLBzLaVafYusRGXFDD6
GJJn3YzL1wt8WHHoxCo3706Txu7Cpdgxdz1Uo3lINz7KkhfJt4NfVQgOoMhXDXOb+aE34fjul3vn
DMaxmAN5160bhGE4cqnaeq3CTtdK9KHW/BChJ8OppaeN+01ELkPyZN/wXgBA74YdorTx4t7uB5om
8PqMKpSXe0C7+u8A7AJY3fvqD61AaSvnNhb2QRklBgOzyc8I5LtZN2Z9f/wJ08xbh2NnE0TxE2uc
QbnXhHviPlUjf2aBqFgtGgHI65o8UHFqekGYtqjKDwu05USToYwmphRTOOuKxM9wFhMXryEXzRGv
IvUYGLzdWrhU1QSd6p1GnIQZ7LA7JCnCxq9Lpp0Ivj6qflaaGOtsvebfjRyuTm6/2boak8kp3Ad+
s5VyyMoBUhfiqA2PQAopKQF2cErxMOh+w8LC4DlXPGZ9NeoPl6mWVHz2S7zeczSQYs2iFyDiM1gg
BXra7SumrhHQwn0RkETU/iuuP+EmhNuMPMd5kWOqgHbySPBv+jxSK69dEcUMafOFROOIQKL57gwm
nD2P9GRGqoDL/wBBd7uZvDtf42INDOeyNaw/aQ4Pkw10M3Pthn+jZ+iGjOsesqB4B6GBMSntT5gN
gcZvR56wuWc0RMlJ5tkXf1Wxbp0CRJjDrD6JeoR9nTyVVgofnyjkqJh6JUi2i2/eQiKdg0LtAWiL
A2yhmvV9jk6Z+Al7/xZhaWDC5w4s3BHj8U2GcxRaIRagSxX4nbidiUcXMoF2Q+nlKjYSwB1RJzrE
xUBk6YmW1O8MJakuWvmpjYoP9Dprh/BmHOnhSdIbbhU5LA0nIk7qPSyJYeNpE9INCiI80qgRd04B
N3qXWWOiBpFGHJrFpAHF1RFx+2byujXqbcHUMpVnVOTKYHXZpfNk7rOotLIpZOhw7ZAeSwYSH3Dh
KtXikdl1Hf5u6bxQBiTw16eWsDkb9TFonP6F7+QrEPDk2m78S+re/q/Ua+DKM5mxzm0a0Na7ts+L
ePC20RwldoufAvXqdLf6ffvHqo4PPK/LIB/umanwDY/IepU1xTNDC+o+ZydhUR8h7mmFMTw1Xu10
KsN5edxDDvaZ2gI7pPTOnvhNgrwRDMpasm+2JTB3OWLGnE6adzs63dg1+1RrrZ8xuUgbg6ejeQN0
/n8he7YuSMVBz8P1WmOGQYo/etdPO4gPT8mA3brWL+254m88j4ZzvKvUYm61+DrLOkYqs1lFCiKp
IDXEUi4+/q3hAawvz8bGopMVE3GD1UpfMKmIvDY6u5NAXsfsDlI2VRyrtgeTZ1On/Bff/EL1ftlz
ADIqtdcrYQLiPzD36+NNSszF7cTpqGwSBbgrTC7BxsFpkWdLTjfDgsmMWDXI/oPDpzwtUc1FJAI3
kv7l3ydyIIxbSJHBytTETY/tNkbqyb0jbqEG/fcUFcDp8kBzDUNPEPsyQmLxh7EwbMbAly2EdfwG
+AD3Wj2fNe1kVGgEcoZpBbEjoLABqJTtR79XpsINkZaOqsLZEG1xDeEKO+QAUxty60qQn/ngHdB1
KdtIga6bgNM0YSxmbfo/4oW8lR9fQ9luifJfQqn8AFfqOzooArbRD7yb5866wRVn46al//OtGH1E
glrIia2iB/BSh138hXlljB10dqGAuVBEcd6MhkUJCCoeklO0ersfLqYMNn1RhpoM6mxRnkmpfNmB
kuLfb/abWNxeEKgmW7rjlTz2fJqKFxdkjlFDVrTY6MHjgRsxJ3mo2PcrhDLf4Np3L9NZVKNqv7sI
8BMgGKlMn2jUmmUeSmo6dBJOqrsl9eSF8IyHWR1JY8Y67ee4o3h3bWosG0rs7tfBn/z2jJFxR4kI
AUqQ8vM5uwjEvqNNu2wbNBSR2ZJ9SOxH4KmWiT6CLwDvCyYW8mnz4W1jWgAKuNtJPzjrv8QHQcFw
BoER+z9Ut+uTL+yL9TOLpf6iCWUvpooh6yP5BBsd00yxVfSe99UXf4+qBagp1oeM6yPuvgZhI1rD
RJb7Twj0MjuGZCpi9juv6p1xy/CD9KHfwyWqv1D7kagQ9dTdgloVIfH/VNhDDevpabQANLmReN4A
GU++rjepO76aI8ftGm/BF8dyfsEujTgc/5BnKRFeYJYtmKNaxmZyJYj+GqMOZ7XXYrSeEkUZs/0i
cLufI79Lmz250iGzuFCu4ufzbs86zwL0K0kh0DDkrhyHxQ4owqZAlSqNzBey8CK0AcmZXBB6luOu
tcKvn3PNX4VLaoosMSN5yFikU0kYVR1KpsAZphEE+192KrTS7xmmk8RIRVpyw0XOdI6Y1sbyS0jd
U0cHcFKcFdPezXEICnHAi/FA82LBWljsLfL0WdMHJJylUJl2hWheRQZPyQOH9Mm0/qCsEtqcOCAO
YtQ6NxZc/ZQ4RRIFVrKw1amcwl1ueWRbSXQPZp0tIxdMZ1NxZbUuRcpMWz6Gda+Fm8Y34PUw47pH
/eEGygd1sg+mx5UswVlERu9XQ4Qpzy5oV5Q5xfqRsHouqynEYI/3IYLRElfzgAwMMp9NBuhydEjw
fDPcvpkrcQDlZG3y6wc7DBN2VO8FlVqomYpcKvewjhGkr7Dow2klF5Pjmlrvj2DJfKusVrcUnXY5
CUqVCARg9rAfGULS47Vws0wWUbFBIAuss/EjNLtc7qtZkB48I9G4RKBAzxThbOeOlAtHK5sULq7w
gbTnEoZBkhSHy/Q6QNfDUJfNisZamXAlXRIuzzDOUYVu+Udskpg45s9inVhJtLstLXcRI/atB06t
P8TdU9HNf0qxhBW3f2FuJSeJqIhcF5bshn9pIcuJ5HJstPpOfei3safrzqODUPRZXhojrylEj5k1
QMXc/1y0xCQwnXKs0Z8xgSA5u/0OAfmH3/pLCiV3fYHo1vaacMijdHJQ14yqmdbznlCg2MG7aL7/
3+JbSDW00TxjPNcZ/s41r/AK9F0bhB8/IXBUhZZGpsvIsvVXU9+c4yAkO4mCTQlITR2bnMOXnbhe
db5oGaO6WTmoixU56M5SeF5FHeZu4BN8el9zhQOPubHajl86BSl9OaD4F3Kr+SLTuqwG1aSICleC
emwK1Ywz/xP/pG5Zo07/ob9OjxqDLf6NXKyN/cVhFOIxUFbnwl6M9ZnUyYr1WfahTtiuM0x8y9JF
niI0WeF6XwLXsMtUsq1k7rgc1Irb7hYFSa1ojZyD8/Ri9/BAJfoWNnbOu/5xaEvAQ34SBZ8Iz2oK
YAYp6qJavuXaDGSlWTzJ9ApAoyBZOK5ispOyzfLpNHVQ/V7pxbziKdXVpvy0/2Bhee2GAWLdM5bi
Tvm3DIe+hMvy+/kIVwYCj15wZmE0H07Q2LZOGABUsTcaA18viinskiBMkoUmPE7jLq1VCVj+Hc4F
GW8mKlDB69cwsgaVxlOAiEG6l/7W71HOumUCXxGyUOBAqpAo6LSuGPKpgeG1w1fF3Q+iSxJI+Wdj
QWzW4VIIaOOs4lsmgtpXOiaPCPzvwsVuAu+29Qs5Ekr8vCADhJUtVNOo34aXhLseKbST/gQ+XDRr
9rBeHIQj5jmqt4pvKl2AQck439qWy/ot1/DRtdgAwGKFGhWWuY/19+gS/gPZHlIniOGZtD0MHe7k
QBPN8A42tXdvRCrISVWTJRHniwoqXja50skEaEpTRbgY9OuQVEvsfXDWtKPqbp8Zi/wbi1kjj1O2
tLZpF2nrTj501EOlRw+qkW0iJvDKxNyFxo1kpcC513j6H7KdJeSnzqnP1nyDnQBiQQXvA4eLy2Z4
VXXbPWHTMgNlnhjyLauRv4CWLEszYN8JlzfX0ihSZDrUCzk7CV53k5iUh5gfnjG+BxPiiiNZpTah
OjusyzmhogmY15yPGCCPnYNOW7SrW2ACUTycWAYgidHuZHlNiBrQPKnj0jrFpyqcDWqOYVoL0Prm
TwIOl/huqcybYH11eHDJMmsbf5zT4+LQwQIAuUTyXgnliTmKtra9ZpcoAWuyDKMMJ/SMfyD/Mt4s
1AD0lY46TxugF8jO1OOqcqN66nPk309ghnwSqioy8xEXvLb/D9fZAfoRuT2i9xKVgy4vntg0ERbp
k0xvvTOhNnVGxIyVlcr0BN/TtS/UCfn2g0Ds0RnNZHOdMmZhSjsZn6FvmiDhk0ueFRGEDoKiqcF9
5IRGDHW58LjsD1VXzha7CzI/HbuLbWUbVj1ZCIrsDzMVgmeSwIjHQ0Q+cGiUuPjeNaZby3gh8hVz
Nby/2px5u9x3/JOE4jSViZlrOb3Bu8CYDSEm+YhE0tgiIvHtEiDWD22z4YT4+e3kprFdMXn05K1x
99KHXLx4vsLPUBLL7Uhe5CmNPyaLOSPfeZ4O5HSW5MRfY6qys1aXsy+m5GezEbzfD/OjLMZWLWvu
6Uj4VPs+/jxQfNinfIMw8qkWGJOa9DuOW35b1ErSVEueggWmDpvFzGN93pSIdVuxy4kSwSFdEUbK
g8Za0vB2ef22Ld11w+u+uCuGYL+maSNGiITkd1IOEAieN/mE4vQReC+Hz/zP6iArS3znbztC/8HG
DO5ZN2SGoImnG+3jsYKje4xnDK1DN3kH84zzjHB46PJyVPg+Au81LCevS72lTXx9JU+ZBhiXuX1g
yhL5fsEzNmM5VTzTccrWZwcX+XY4dFQqX/DILPTuBHZCAx00TMSq1T4LZqI/4NPj9HrFL9h4HT0A
z56FvWygpCPZiAzl2GBXzy4IsYRKfpr4dBsWpTA95obYypl9zyPQMRm5S1os5JzGH0mCcIQ5AaOO
VRuUg83ykiYQ6prtNYkjl3WFNb8ejeRRfvSUw4kr13pHSlXurpHf7xccsBBNynhW09n2XMg2s4IL
qqK5ymi5tTB6veG1bVi5zAtcaJ3EwrPpVCgV0cuJzVGTuJS1Wx/GpwKTmU5WeIVSKHR+Q3MiiKTt
x9czjFWknOxt5nsF+KEk+16FapgYsXQJ4pW/9Im/ccdLcJTdkfWC4nOh81HLWIZdB+rRWC6xiSI6
8N737CdL4zJ/H0FxKF4LVDSAQ1E1Va357IuWUNOvP1Mpy/wO+G9L5ax4llsmFDJg8XJsIqnmmqD4
uIfJxeMgW9IcAZsV2Uh1Cek8aE/nYeuSmdtGVozAc4OJ+xjwCaTyTNeQM2WolHr9nNM4rcE97t/A
7X46U6lOL0xvVEYSiTqNaW5DRQzMyTDe+nyq8Vcj/9AQoRegBb+5u9S5O9FX7TNtKVeESLIsL5ug
9gZxFdkJ278T7cBRs6zMdA/vwujLqnpb8Ex4e04mFkOAWBJXiI5TxAxFor5NR2XhR0dnRrLxpCTr
p0parbfesXcc6hxwkR9N56DdMCITU8ppceIm4aKqjqzcRZntXrDf9L4UDosS3CHq6kvivbCS/o8b
c+XYfPksdTq8XzdGbG0du/CZrYZ24Z/naHmM3QM1koWDnwWL/mf1yEDUZVGfMhyekpQV+zrSE0Qj
AGa5B7H6SACZpfIN7Af9usPiRmPbDSwH+MFYlHUtSr8bQhg4KJPdBufox490JaR64BjQLUvFUpPJ
W94SCMmNmw2C9lWREQxkPSdeL44SdIJspQMdAdB4g9O2xMo1ob5yxJ6DumqtuaTykfLe2v2eral1
f9KjZzSNYoswjAZErmWkQstPv/1il1rFgmAV3KJGT/8fe0OoilTl3vMWpYkZhhgVNmCCl/BCMOCS
owSJsKRxyvBOjmnLnHcL2ZQETR9j5EsoqYV3BhmRjVgWD4c6z/tG2fE+cl/HsvbpF28PZkxQ0raM
uNDivwFrZ/POQYaH5BOqG4mkSRhzRKilzS+Ew1KfRixLB/T9mbtGMrLgfSt0BZKC22388/b5wG3G
GIgT6LEsFELbFi71sm723InQJmliHxMwlJBgos8Nf0jxSKNK1Ij3PQ/DoWFqrkUG4M10Y9nVAgVF
BdCgEgjp0EH+59qN2A14v6cvq7Wq6lLfhoc2qc/WI6NapXpN19U90XW2J5AaIOR8ryiHB6Y34ZRz
kwus7wwGhNj1oHz1tWj1zRbsSJ89VQxiIrIU3Z6kx3rpFzO9hcYF8e7HvDcuyGw+uoz2b1MUO2YH
k85ZyunbfRg7PR4UbnkUdhEWETUXdyG0wrUoOOxT5rSfcpGmXZZFi5u9mrREFo2nMP0lAbGkLONZ
Y28OFXApf0glFmJesb5HIaj7R8WggEg5KrQEN7dI4LBmOcqiWei0gQ3zUmmLg3RTokOjgDrt38jS
bZ5lNd4YDO3PISrQwhnRjtx9cwphOXFJaaApcDg6GtCiS8MAOXQDljJuvFd/Ox/DM/bd/tVvZT4Z
mT64MW7PbOaDvAXDIkrfKdVtrmn262aNnvUWFxPEFWQqNIkg6dDas1dSY7QmKIvphJ5zdp1oKg+h
fqf/D21eMAw+NxjEUdwHROPJ48ht6RrZYj/87x12QP6R2MYiOkofphVtZh30q1Uv7R5B+GDKkf1D
5GjOk7URNQxBfdaa+oRDUMqna5NFZohe+A3w9WwHcA/QZNv/GLCBC2qnFyyZ/Zw8u8zYBYk1PJbi
6Mn040vNh/qSw9I7gRfB4pzlDi9cUeccGaj2YjkXG+YSuSQwiSQQT2roaynrqdCwoko4LnlKgQ3U
/X7/y2K+0M/c5Bs+bi6TKpT3/za6g0vNcX42Nl9JFzOwegJWaBgvP2fe8SYYPJ2TsgWqRWggrVWe
URkrrs+8aMYcWdcBUbsF+p9LSKRymvMBewbTeTP5uP407YDS+QXqCmaPfq0apsqt6+kz0Zz9beeP
unEM3t9/XZDzUe4gdZOG74PartyBGQTs0EX53FHYkjQTf1++2DZHqb3CsM7zcuWJDt1nxXFnthEJ
55WCwtoosdHryQYC7KhI8xwRk660qBQo0xE6395VjeJGgPYv9cMNfhDQH9bTBUZiPb/elCk/tpn0
o+cDqFbutoGKfaE0teeRT+9IAZmuNkY9jLaotGfcS0bgTtdM5pV6aN0Z33yKxnORqOZDd9ymZwN0
w8ITOUmOvHn+WJYq3LG9fspfXEkr5CEILbARSh6GX40s0AKzwP72gJhc3WCOZZgIBjXyCGiAe+gm
m9e4fksRiQ22OdFLLQOptV8tE9FgYw22KCScnymr/lGyoYUL3jlSKpEgJyF3Nu48qfFdimchoS7o
s8dPyGr0HSoEIV20jzcBsHwq8EAufKC4BlreD5A2+rXpdJunrZvWlxSDWI7kwONW/3P7tQ9onkAs
p5N1IwDOmffq70B2mtY0jnabu0QXjoMmxkh/5Ii4vHcJz+Mff21fXP20m8tsz7FBojGPSDsIywRH
WakhJmr9dyA9YrulTvukwNWXyIUIfx77oBRvvdxZdwSo/Ztm+sCV+ip84ksEPSGpubCYDJ+Mfgdo
3zeIRarZF/Xtnx1wEq38QhXPoYLWLSbnvU7ra0Od72KDA0WXMgNt6eIXGlyYHLKMUMSf9MNQEAOe
QRSqZ+CQvfwu4Kz8WH5R5+O0ozm7o4cd6J5lBC3JwlPb6CRZZzWFmDR5Z1UY3r6VbWPOT+oR0IBv
4FerppTes0ve0tpH301Zl/L+erbTf4YAViX3LBFI+FsGaSaPnzZAub1FqX+TPlxKTdjBduV5pmui
H/AHSleCRC4IPg0kgmeO852NAmggZ8LUK+E6yVtDXMkOfaJPn04HbgEWBTgvkkMUD9fTVY0hV3ul
cag1HH/Ud0qBBZ4l1sDcvb5uRrZgHmbSqSfDm9I4x6nZxgp9KSQJNWvNRl8GjMgZmcVptRcK6IjY
+dCpGkxZVxMSyLalauVjtbFD/Cv1a66b0wYp+Y9AZkveFX5jM2+YOm4l3IHiz1i6ry9HEYmjeEtd
GeM92ukHb+lLcHqWHbYhXViuOpmPW6YViEgP4ztF35fyQnd4NuY6Sx/FnGT9qWLdA2v3y+Rn7WKQ
IKt8UxUBXueHx1UB+z77ltpUQab3u0TdD3k1NgdKRmW1X4a2YqQJ7sN4ueoxoET1lZ/OYLB8vvpd
9cEOgWoZOeMeA04IPXbQTl1LD0Le2/TQ027t/rYzFM8YguSHC29rkBl7MEW0eHLxjp/7fZS8ppX7
JKgIojvTOFyTqwoUn8D8LiXIvbv7FF6Oh3SSAuy91hJQbIKr4BAuAdfSVOMh1vVH+FI4acl9woGW
ehbyxnUYBqhMEDlTks+MaoXE/iTLNtQO8fMhVK2+/zX52aAEGkFJybGPe+Xq6lOqDeUqFJuua0zB
GnQW6mYtIHLI5FuYehuM5qjcx0cJKvBBKallAnHmUHv+esiTzCySjCzojYd1B63M99YvRaTRHUc0
kM1Enx7qiX/zfP9csKI2DBZZYoeaFXpUh8o+M3cRt3ZeQ6EJdWwuN9kU7KEfbvExzSqdDDusmsec
WtHS+HKqrsrkhSXqnDeKAaUxVhMvEaZpyUGMObjjqx8nNSvaVgA++0+BXQ7WJr6QaBv6iTtmv5HG
nRfltbHpPwDQsMp7zPlnCixidvUzfgOTvDSx9256nCc8Mue2zXB7CLjex5rbxTFS1uK6T3FwxK2n
kwyJwZLlRpP/E99gnWAUJ/d8WXWgKfIDCn6YetiYWJNN+aksr2cAZ+mXgcD+yH84AMmwTRFpEivB
qidGR33eVzWKLzGVCgjrU0uua2XCVwCQpIvDUDfOT/9O76mLHvY9Wnm3c1XIgjz1oOwXe6O6nhve
xGgqzEhM8Vc31WMP5TYy8gz+ivAckN3lm/QztWlUQYLpiptLrBkbxVd+loPqWWUhKN6TZJMT6OBw
iBVEc2+TfV9EIphdFPlRnVw7/XHcaHIZERdl71Aci4RhDTcZv1FX1vREEouLhC/b95sUUx6+fP3r
86tXlJm1eM9cdC8han6P70BNIJEQSPyNY8OlRUQweuzt05ic/PmpQOsgTS7/ZpW0lwJjkdwaWCKd
x8bYjlOOqXU+GdlgN4abEhuvxpOpAQDAeo/N8uj2tFtI0a9/VgZ4fCYxJ5lfXy0U1p82xEGDzXCD
DxMR8RZJtiiWxZmmu3k6Gg2w3eBi0JwJMGrp4NWei6em9XJ08zyUInklWYsfgrYpfNJnwZR586Nq
YaIfNScqd/5jfE5yDKq5JfZqZu1jmntexWOJyWemkZoHX6obfAjQF5C4xUVcga6vhHLf0PEEC7S9
5G4rAv5+LH0ExsLKaaa7ngDQ4dBn5uiVPsd/yW2AxLZvd5U+qUA2u9dLZ2HwSMoac66/kdVL6eCz
VsRMwYeEK5EeklK6Fni8vGtYnRFNoqS6THqggTW1ROo7HX4/loNPmiZ2+6eh8Ygqy6oTY2RsWxc0
QEWHIHmJ7LMeJJn5W7s6FnWmltUMelaev/KEDfYKMgBExDBQYET8l/kchuokGgCtSVgn9+R5/hn4
l4gjms1vRP0CAsm2khQu3JxW7EHWadM382W6/rql799ZaCz4qQKEQyuIJiC1VlI9xZ77DEeZnfg5
cFu7RW18VfC2+u/pbQ6J8BsczOzQW1LZf0RIjgs/FTSQYcKvTR4LWmnFXFL9NNzAcxu6pwTsSlfa
ll6iPj8ytTHHqZsCpYqqPMKjglIY/EitGU1yugpR0mh2KJIgefm2XAm/QvKDT920zmymfwnCz5Fd
GD/PgB7ODuq2sWUrV07/70Ym61YPN+FncqzA1xn1f3Xkr46SdJs4Qaociyfhuo7BpCIFJDbbUfdQ
FY4V9BNSiYgAfxxk+STKrImRdEfAi0TswhqVK1fJKicYPn3BTkj1v3y5VMwXbo2KjqBKRik4Aln2
IaQJVUaJn2HX4DCgOMvc7RwRC6oHhRaTjIYNEz1VKgHclBwiloGgcdvqpUBPb1JQ4DLBHLANnki/
1hYxKShqFZsgO6FwTDpN7mwUW3rUepmSKE+DMGxyk/XRKYmFuYjyvo8H1nbmHzl7W00yA9StQZXb
3ekyuqHiaT6inHSJLPIFsoP6hveP+cajdSsaR3Yx+FyMBbqFQdQ2Id7L0CLwPJb62j7NjB0Tz915
kdSF/yEP07K21gd9drruGptgD+ciLjd0KfAh1VSA/Ovl3O/y73jyJXMFeGLoTWUR88KT73aFQbNa
cbGmwO0dyQFtrSFJ/sYxrkKAV1JhK4Oy6QGrq8ihsGLG9LM6pzqJul+Dp3+ltvUaIMY/eEi1Dkvt
SMsJ836u3cr7m5CwjfmbbyxTNIGnucHQgknDAzUb6xULhumfyOCyDuf/wxjlnonoGbffHJ7+UzH0
qM1+PH+B8grRjNdt2wNePTYV0N5pDwb0YbaPOygXXvagJrAGegUDHUtMPAz0IGnz/kt8Liie2yKa
VOq3geR+z4JpzEtrmi2X2S/M6/EIbvPqPtDfk75DoOkc0eVKuBqzZ541aSl9gL0MOV09ZqaunZpY
9ue9sC3m84wiYEB5Dq7KS014NtkwI2cXBgPq8mlu9j46fi6XLFamCrwzBi96shIzz9b0kBMf+Bkm
1fwZdzo/PzYTEMtTby7Yn7UWbkFPhJ9+rO1IZIUznh7NcEfWQV8AUv2oIsLZlC6OEvHvrE1oB6eb
dyrq83lo9Zpjmn39MPvqDnGLwW9fz1rTlhoYkNHx7VA+M5fJsaoYTMz691y19YN3NPkfhWWufb2u
ZGr6XK4d0lK59XvBKKw11vV9rkh1CoXcTBo9i81rbRKsRWKmEmVuD8PZGEX+zSk5j1jFvKHh2ney
ioh90ZLWYX8hYF29Mg6xChZWmoSad6UZDyULt5mdXXeSjJlAnpBsAdHh7wFLR1m9l0a/VIXB+VI2
RZUK4Hkh+O3FTV8Y1tYDxiq3IQBg9y+nTgJnCUQX3ATjXFIzWevHnAH7rzeFvfszc7XdjJax/JPL
aVPUlImAxF4zU8DbEhrFrgIrhGvb3rPxVlHCNKA4wk/U2+BdlQ8pI06lK52Z9Hdo/Wk0mVEY0z9s
shZzfMGGYwpbf4kUM48F7V/o0oHf0nUiEUNRUBnyRt+d3ZqiS6AEgSjxKDF8YxdYZZX3INsMc7md
LsLmydm0hakds6fAZWdMQ0AC60vLzbZ1YV0xiRa1X4Z4zW9YCBrT4+Yjb6PoOmkUrtNeV3sqRaSc
Q3L4LE52Zny3No20F/cOumVrrEjfShKFA8P38yGyuwXBEW0z717X/7jJthe8UpY3CLKqKtmKwEP/
/CFpz5NxQj59qO1VseO8IRFu7j6s25cPcRjE0OKb3LbLMa64aQTEEGMa/cWxPTsBD402Ica9idHE
k3XXzCIPTpocAPjTvgXAzp6BBTHuT4sHqIrb3/GN2SEYGh2I1HW6ydUFaLZfUV7hbSRkfY8ogX5O
DJm6PAKevW0qL9qI1Y1rnckk24KGbOfBRPw1/uo6aXBWk7fp9zmSYkplEwXS99OHX+O2uLeXzNDI
+XxQai/DRXpB05lC7kHJcGzrHaYMHZkYIupwQpmoP7tgvTiZoalZIizbFgml5E6wVW/Qx0xg69FE
VlIdDhsrrfhKRXglDwjFXJ5TmX3VCE0GAsyMp5u+EKjhlJDrLtH5Zzs7XXOz1BV5JZv8tqDfsDRJ
FkSEuMGCVwJqBMC8DlvVtMVfq25vZG35Oc4vpv34TGE+EPlgZwYTEmsyocMJmSdpiA8zZMkgu8jM
ZRu/hxqL7ikA983gqrxK4W/pn2zu5x+8NbOCwBg1bGieJXWETuhx6vDIa08XXXSyy5QI2Kq0xtTy
tOVITvNs3RXs/N9XUmVRJo8+P40MFFa4BExR4v0DO/fSl0aXX6h4R8HHECV6kwUjorp1f0KnmJL4
ujQEBVbQpwE7g8DdnwuKRPRvqfttnr8wTet+pPvA02o9IAKkCxbOX04wni97ekpvwb+4HaIpfkWQ
BWY22iLohtMRChTjwxKQEE6+xGwKdqlowfFvRInx6L5lwZAwDU7oBLJc4q03LOGaPaPqaNTpO38x
b/4In414vHp06Y/V5CBTFzXTZzgJpU6OdjOUQMuoSmCNL0XkHtnJvGu5dbXBZ+QoJE/YmL2Sc2Zb
ygM5NPkcBGsuMFNn4yMzugZkPNlXTyYfseN2DJ6W77Nw5nz8Ws+NdCYDx5ImlF2SBWHgY4RSH9Wf
z3Fx1sB92oaejx4PwzIfDz9PY24oxV4Vj9g8GhS81Ny/peqLoIRl37FRZACarD4g0NVLeBWLFM6A
gDBlbQfvhSmitT7RqIZLYOSQYxL5w0smhKvc1ZeQBL4WiKfHZfWcC81t4LKQ3w50VCDnUofaVe0B
GYcGJJXIXHdc1mIQJUNueWjpNuINN1W5Ye+N1b1EpR1DPfDX0l3cvS2812/SXwiREqNHUaZSZKVb
Upszcpx5dJYSnB66QRm0iHLTBUt1bFA7nFIgeChGSpcF2STSPNA3loCAmbNULY9pyMvKJm+9RVmR
klsr4MD6RpfEvPdszovz8f+F5hVVPEeCdeIQvJmd3p4JSvjTWZlaOJQfFVG8n69AmZGY9QdF3bMA
GmQ4cKEkzg1yn13h6sXIaXEpoTIpYy51n6rtJYaLnZIcaQZ422oHeUckjrPU1WkbBTwleVUuHbLH
/9oATEqt8jzMXXzPZw9WZ+ErLc9JAubN6MAjWJsRH8jVoEejGkyV7eBew4D8c9txbweyh7kNUQkx
aTvqug7UPA+a0epCUQ4zD7rCktamUsn8+y3mKxoZmXB3wQmsRuQazeaxSp4k/DVKnpwjSc4ObwpU
L3WJX+X68Am5SbEhonKztGbuy15DR7yNnUkLwuPkRYpo9vFxEAViGFh/tyIJBKgy3wlkrWZKK6Iz
08UMbqWmIlXZ8jhFjBEwwyEGpowntrx72EKVGZJS9b7O65W7sDCLyWKV4anhQvHpfZnfMstUbn0V
R/pKzajIJ9O7kxR8IcP+xL7yja5d0JZ6Uw6sMF8pFbRGDqjPyFbs8175oBOqw/OZQHDf7n7I+jGw
+nsq54JlF4fQC23wPJNIh/AOyNjGqmxEs+mQFf/RwPs2DNLvhGsMamGC6qA8Y/7FsvUOtHd3VWEU
ghg9JPFaOvP8oaBkRd/0bzQhBcElqW/nr3xl5awYIJO2cwEnEguUtVZ7d4PnFz41sfWpPt821AZo
3/yRrmM7x0RRa1y/1ls0gLhCq2Tyjpl1RJ/QEkMO6+c7lVoyQwMu53U9dRqLl0wqlZUqi71jzjC2
gGZCX8GiouJ1LQPQxPnKmi2WXwbKvkYpszmqft+4IjElQeUl9gH7PTWqtIlQpeZXtJGxcy/Zx5oi
itYCzLZE1vCHoD2T8jBxAguGqHvwPtyS5EgTXp083kTnJG8US9yq3uYojcJcvySkl0qwAi/QkKdg
Q7iZXA5V2T0rl0RyPrB5Oes+HCPo6r4INhBSpRWjkVTEUg+Z9njylsS3trdhI8AsMKVpBRcmQrcn
fI9SS5l946VLsGsh6vk7zmxuXm7lLK3Sk5vyEp5xqt0YxFaDEnATWGdDrJ68Io0FflqPofOX8ssH
c3bdEuFQXapttzGIAbz1puZm0tr9a1HpqKkLcWZXDAu1C+w59BWBVChTBqPAqCtGGPwDwOMyMZBf
bXtXJfqyT5r/ouhW5ZnFP411yJms6nzWjpemr5e07tZJbmOviXYSLc5pbPHQtw1VczWrJND9aOri
gAT5x4a+xx1y6Wh+JdwWhahnLLQlmahELYVz3rQ+4lLsru1r6AW+PmaA4F14y2bgRzAkz9MFsPM6
WzYsnLYvKB5Oay5aLR0XATrYLZHX2caMobk5WtAf/R4szKUYbjBYz1HdmtccfuobigzJweiAjRQu
9UntQXxkGp5oLYsmSOXbIAy2fchTmvFMzowGInqsIme7yguisYUACVBCCQhMYzpd+3Cc1QDIOFND
7vZeOaYP7LLVue/o59Awx9ky6mTIVHGhSDNKH+87Jded5jAdl0R/uhh4xGC/Jqvrje84FwrXkghd
ZoM/PrdamRQ8ZguN+pkFaxTKJ/mI3lEoRnpz1ad5Mdo2pkcAV9Ac7+701BYacRPNez3WBwr3TOTt
nadPDxCKghxW05EMIw0wb4oyOJn/6E19tjf2FHsHdmeD3lFsvifgA9M7HM1j+QoDB49PDj++nO/E
llGQhDz8cLjCdAyPpfOF2NXQ64qyJsD2DkFDEG0FujaMcT6pjnfzfITsTtPxPr+ZNxpXLswBKdL0
iFjEHgEk/tvxzMnYdETIox5jpNGkxCiY8GNCRsfwTinkBrbOj9RSJr12Ha0lzOgHp08WQSl3BA76
1aY5tg1hLYFOavsfy6hTXYaRBaATxPmzeGbFYB2hcJNNhhQ3XnFp8iKLp/LOK9tUcGOyBdH7bTN1
7ShqPCk9NP+M74hGMK2QlmBICqwdDfQbkEJaKzahVvJvHwIq3A2+alCHUxgy9U3s6gApHELn8/vm
fy+lHQdp3SPAl1hqAKkLX/QRjL5ZLOUEUtnmTT5QAUz7WAu6VMQHGug1BAOH21nVA/GmXelnrcpK
Fa4lhwj6QGWHPTcwUJLwjFAprVgnaB5T1mTT0WxbuHOh7B3H5bOnmvMwkkktdK7E0Iw7m7brks1Q
qsrnuFYTwaI9SJrdhOXAqalF+EB8dYVn84TmrqhsHQValNkeFM9rBR3kKMjJYKlInY9I8SgoTeOf
uis9mYVmp5nQeFBgaNzIH/6VEQfao1xdrjoJD9e2FBpg2f8phNCAEYaIAdcfkpv6HbJ0LCytp2H3
COVpg3jvjmdetzdjAieVnoqAekmrjgWt5DPkUW/v3VL6mw7jIsBJruVd+C+1RSXHZe51eftP9puG
+Jz/su0YKue2t2+/hHrGHAGK33R9UGGv6GVsTdbnSOU/xzH2YxckfwI3IBaNOIDhX3duZ6BeNt1W
fQZv4ZMl9mC/EP5InGX3jE0pe2ifwwrKyAGcSd3Jxah8SjcbR3bEQtiFgowl3xcac/l2TeVKDXxj
BFscBo7NsOVuIsfXROwJ0XaS/w7MlA9bweiNxNpPzlFomkHYXGIDSDMcXRm1nlOiAI9pDAvxrWUf
/SAGtW56fbgjL/kC5eEe1am2WzJIHf+RH0ma8Qo0imSrKGhTiEi63zHo2mkAa/CWl1OUmGCH7ehg
x0eeOthLGhBtbPXLngLwC2BeKhrdSUlqJQik4w0RUE81CVmA/PL14Lle6OsYQUoQelI7BXDynL0a
sNnNidwo34VIPXBnICkm1kE6DsQvcCn5Wq1zsmJz6WqvrTNFiHZC0c+urLha0qv+bIEDBBa+SOyG
E1bVoWYeRQXrMpqGc+0UrlcYHHnA/TngOGlQM5+lpNl1kHRP4fnA7VVDxGpFGDxYZzW7u9YaA/8+
oSj9Ue207eVB4dXhYeRMxGlC0ruvlleFRl9Y/YA0eGGgHQEoJm2mdXgMvUdC6y5ZIiCb1kORMS3h
5gIwSXGusxctXvBP3m6NH+EgmiuN4mxZPkj4Z3+9rJaXVNDEfP0qmikZLCzqQxD/Ph0Z6dhhqTfS
w+j2sTZ3V+Y80slGGxYF01AHAHeUhz8yjgftOSbVhL2sx8z6mycCXL5Mn7207uJbHQ3HmlDFy8Ek
xXUFleybPZtS96TpmmDllXmB0eb62ZpsxH9N+X04D7PFii9X+Xu6sn54YM7MpjE1cbVYPItq6iPy
ldsh42LCrf5dN4GTwbZYle3XFZlzZxynDJGCXOdXm5GMdI+tXRVbbnygEjP3dKL25cmyRDrPajim
ej6Q6H1JQwUcbFCut1hOwFnlMzHZY5Mnfkb7zZHchNiB6/CMpz8lUiO1xGY+aAEpd8S1pNJXNRnw
PV7b3B7XJ3Ra4Il5UCCxBQG0NTqnwbLt6z83v9PzwDj0QbPGebefQb/JNaYFNdDGiF4/xjFMUvqm
k0duxQ2xYJ/JEzO0PTspswM1tr+sa33mu6smyY/GmEaM/uujeol0Czbkl+6iRBwRx/MTcH55B5dl
R851g2Yh19mzkjE1uKdg/UvAgnjyEmWbekD6TwSpMfh/FYiT5M1y0VMv8G+etkydKc4zlHZg6QOX
kDS6HII94VDSpbRXTgq/o36dB+9W2kUvjjP6xGHkPMzJwAu40w0H8mv/FfCwpdzUmM1sreqe3A33
Xu4vHyM5OnSqg8vrYCG0YxPU/fnzKn1iWSgA1e2rHYCM5qrhcjp+tDi+Xfl2h2yYCSvhKLrB2uUB
iHmUQasFboNYBgqbQokN3JbCc50XLQoneq8MSpgk18xZ/fpv7QqmewBIRAExapanDr+sMFZOOjvZ
dFGmPSOLCbDR9AK7wtBMRfgMwtU+UVZczDTvtfxxu2NNGfX6pzrv5+z0Qtvn6eIApV+2K/XMOyO6
UhaRbtpwpK7WlwfF6AOVypmTWzL1qC6PEWAhUHvq0SQby6dOQDG0cb/iNU9zjaHAybF64ApeMdj1
TRjJehO9dQTjDeUoY4gb5679jEhXTX8OlxlMdHd7HQvF0Ie1KAKBzkc0BFBD02m8Wmpk9hx/uOac
Pl6zkPvA8nuNZ9oW+JXUgWscSvnwCjnsW87SMmO6PZDH8hY1lmWkHRV9Pnc2r2sI+YWHU15tLeSI
J6M3wLt92Tr+89ELa3pOjR/S/Ub2od1vYseU15b59dL4rkw1xC2ezE+hBWTkVlT+Y8oai87TlDlY
NMMxqMVIckaVEdrlFcidMeKp+fACSCK6ShxOFdEiGdzGSKX5l9K2FGjIXkjJFOA8/cM0eOLgDlmA
y3Z+ruC/yFKA3PUAVXJBE3KYBBvo2fFAK4A41yKPan8n7nKsJs4dS4K1jqfksFT1Lkflp6N6LfdH
nN/dpDxbuCTYO+d7SrBgiqYsyFPsBvkUwW8z13N1LP84ZeThC+fHroo2hmKOXUCt/v7tJDcEgTpQ
PMCWfN0ds0r/5OFnhI62sbRl74LcsEkPYQVKWRrMPHV0mrtwNkh95m5wUuKtqZyoGwpNr1PqFxGb
nwn+N9R5jJuYXJxBur/U01JQghUSZJxze/RryND7cWzUkGWc2DzsbhadD3WJtoKBSLAH10ZRs5jN
1XavE2Db2X8YbBGrXn3HAJnftzkY4IGN11OS4YDKzH+aMylYJ71/teGHvhSFWrs8fpML02uii/Uz
vWu9slC4+QQl2uBiepIB//ChC62HCstLuEY3dWODrfvx8fNs49KjBZAPP4tjibryuxz16n7z7pdP
PoBQBg7LZr9og9pLcb10NpVRynteQMY/xQKKXEMWmTfohEig9q8WS4wGUfba9ej46wXshLHH/dHY
mONHCSxg+0uZ/PUwqFDeZUOLq+3ztlFqvLzszi1iAYGHCYW7kpK9h79D3Bwa2lnKaVhsFEfAlvnn
dhWy0MZiiXc0kONP4myTGfrSaApkCDfXrCTwDycC8xPwi3xv2NMwvtagx+xTWNODYyuGD1HtxAUO
UUSp3bPI4RgRmIPoPVuVuUoR4+38Vo8PxupKyCDi+9UJrEVxHVVsC5CQ1Cv4RymO9CQlIeFaFSdv
mbQYb7I0Gnj7xlx3OXb36Db3Cgwm4HDbH8HzMHJVeqT7BPPsByrzwwSGXZX6g1hoRAYuitWWQeee
h0vuEi2YW7icvF7mFmSsSd9OnRHpb9E2NodGcy4lNguOelTWEWY89cMmyguWv9SpNADDxj4/XS/X
NGIsmrs5iLCYYdkzxJrLw+jY7x8luL4xSrsi3yV6Uh47EOV4Dg1ptdRW583mn/+7ZUCzcWBu+8Ru
0Un6qN8etmUhwW8AGJ3/XZY6KPLxNSds/f/VCosIIjTKUnK4XO0A+vnOeHSHf9ykDQDIzOCquTEj
DF+CFYVL51LB4lzMAsNH5zJR8oZsCv2/sK5rvVZN31kWwOu90kv4zuH/anfnYMfp4JbP4muCntlA
zd3ZX5Wi6MY1+uouHGoUhWaxxTFSMDkQ5d0UzvOAb8RCY5Bo2NVmuDbgRQX80+bB0goSad3oyx7y
03Ws8h2veaiVPLd5+TCKibUZs/CmnKxED2xToMJKRXVxNB3GugZXfwtXZoPgwKAbO61Qjm/PLgBx
tyKB1Jrh+F53cHT2HYQRF+7IDmD4AAXrUSkOBKGsgYeToUPkC6bqIMFb5GYad/2sH2/J5tcmprGb
wUgT6h+aYC3z0K/hH2t18dSvovd7LEsOOQopwNgt9nEWAtjva4a8OHVY6J2KfLLhRHhRjUvOlJgH
r8qG37GKsIkX/ASJ5BGvZLF8BK44RVcRyWS+Y6AE9lsYbaW2bsdlwcJ8H2RojT/mgz+aBGOrPUci
ydW+NCdxVdogKWNQZhgtXNP29qG+AjC0l/HUiMcy4kxeLVmtN7l8VP7VGv5buDtovGA3ovxXRcuD
wi8cXsxlu3j9I11yLc2Sc5vLh+Sfoy0uv7oPuKEKpgswRGOnHNT9ulC/7yvhUYSdrN16uMHGmIZW
CVY71Hft2MMkOOUdzJm2A8thZ6qqnm0og6fJHjcO2MAnORekgEltSZrS/eoBzaC6KkyvQinJyVo1
SBIudbkZWj2on6EHqZOsLQTajMrcQ2MIBqZQB75fFD0yWJLtILOSQzoN1Wmreu35AdgGF6TQSmHq
s/6ujWhypZcjbSuDwVlRB3awJOTXxNR20hSy10jWEMZd+uxoafyfq5DH+n1jcPikOF3hfx+73IA3
X8d3lt3onzK2Ebokv7fRq4DPL9k3wIu9UJilFW99U6FTjssxTlToWvxxIPv5I+HpErOjlHJxqm4e
F5Kb2FbAy4gg9fyFJlMLuo2sLhk9yJWHM1F8FyPEeqftngTMSTWQL3Nc/msXV25OaGQx6nM5QaIk
/i2XSy97fdxcNXuq1EteS22pLiOHYPXxSUW6FMV00ixXDN46lI9jYBX4or89S/y6pMd0yXBTUqVR
MAWux9dLFzhcglPCaJyuMkUwAsX1RLI/I2WiiIa3uwbeIJWiv7EYfL5NCxY44ZbqS+995LqUyzSx
8TfP0BIGU3cQ4UhXAIkU/Sn9Fw4/6s2DcCm9Kljh8uC859HyoUXoiEjAYEwO1b62ZXpDdRfRLNcA
+nXDeimItzrN0bucUFMMyJE2dPZzwYIxRlKte609msMFyWW0goP35Xa2OUr89+GyLtB+VNEQ+Ugn
GyFbBuv/Q+2NWj6ncEdjWskd5LGMekGHBDTSqH+OGE4dqJZYS4alfxeRAXYmHlL1lxIrPl64JySH
8hSg5VcPLi/B+yCAMwbb4JdEVFsFrebgJPo/HwpGMkXUC72HX+C1fTA0FmkJNuPB9kVHOjCtML8b
lq6l7MtGUsNPi6ypxjCkkYGuvnXuftjJ2sAMl3eq0WdYr214NBCTDxN/V436858undYAt3z9mXpC
hhOERXSmM7pS57JJt5+iotDpHF5hifiKV+Y92yeG5jjWBXSLwF8NmRimFa8JRCjy49DaXq6njHzH
HVtNyumewwaiwkRvcIw6tS31ZswZ0UGx6MqClBHtra0pauXf1ETpii35rwXGOtlYdcX7VL14H+xY
uc8djAVV6evL51FgUSVzYkPXMGiHhi7G+Jk1MB2tAy2P22MParzm5/KlqTTfNNKu6qWzfBRRRKSZ
mmWfULGLWJxHy/8wSuCu+HV9qan+VbHOdDE4lAJob0Mf0GicoFwm4veByip7sDQNRe+bMnEPJ4AP
y8UNEd+pIBeZAgpq9y/UCqZCQV0KMt8PMIyYK0Ix2CObgMHV0VB+GdqOvVimcYQswAIb6wv33OOQ
V6a3u/fCe3fWIASRBJ9nJc8Ycbw6Hd4cOk5xIjH+IaQhvRjGjgzb2dCH34nsk5lXtOqLVxxBLeik
fIEgELkKUkkCmJqG8ux5oAxZ6W2rJy64egEZKce+3R5Zw36gTbDfs8zTdAc3qfM2nNCn6EThLFK+
xidJXZ8QrnnUmgZ9ViQs94Klreb1UHdk8DtG75BN6tssJGb1pPKgd+XDBuEh34TsAH9EOMf8TSq5
f+ZPHlpJ/7IOJ4wxFHMt+3HPS+znd9uI6MJuwFAteITTzG980lnJV8xT7sbpAbSbH4+7Iu8X/rU5
baFbOoLdcbMkveuiRNfd8UjrXnH6H/7l9bmROeSyQYz78uchCwxdijvLS3hlb3JBK+rfuWBE6x9H
hher9dLWwVuMyNEteCJcg4a1Pwadgb+UUZ2xam8nT5psz+1ZdE0f1b/9KzWFHyuKCX6EVIzsrxW0
8mTsBFmYSX9o+vagiBbGWuJ4w+/gzpioS/lHds4fy7CkAq+BuYCVTtYBLKa1RvHeKK/HZZAw01u6
9K0vxq0nwrLdBAtYWnF3eKh9DYvL3ynWbX0Cbxs5T60wBZYrc4RxTcQ3xR0SHi6gkr2At0z7q3cl
IFciAiG4acF9/mTDtkkWxa/CsHfpc7inCJZUv7YlgNOmRVaTRyXFt4eg+/waX/cPOC6APkvXkDOo
SbBQEAyWLriwt2MlodeEPi8GWrRoyE9YRPmqH9Ex9D8hRojwvLS51a1y5hZQzVrNtm4sas5NMEnN
5Gao7dPRUoHWuQr3j0JlLpNgaA/03iMN6l0ofIxaMDX0TuskmjYGP9mSkCr782D9iBsLYPw8c0Ze
WW/sExLQ67xXDr0znJu/Pi7H4eDx+j9h8gZbpC1pKbS6tfxl9GB/wuslqyom2/Tlfnl9Kg8CZU+K
fS18DLmbhqogF3XgH6X9vqGdUvWe6UyuRg0OTChfZMmNVRQutWein3M30Wqsia1xRI3kG7fspebQ
jKq4HxU2UNxHgPX2sFaX9cpOVwGiRiP4zWC8CX2Vk5qbS1eurvZQiWBEWraKQCDga6CQjb5Deab5
i6vuLmrikZnaVxqj6lPU1MbGUTDcqPhi16bk5ZC8WFuUWfZE56sJCCnzZ1XJeZpMOSq39fnl8HyB
s/ooFHXXfF2yMKlMjijx+gI48QO7bhxXy+uh+9oamYsGMuWtPvZ51El7StGCHb7hdTUIhTQpgyS2
2K5LYCOhtpYy0wSdB09U7tibYZJrlTEXHrKOjoZlWm6LtPFMkdELXfuLxYX3Ym+7aUtSNLM+IR4i
U6lEDx/t0j4uDxPCB65N1mebk81lxkpqrRNG0Y7v4FZr+t5K4WBRY7UTAI7OhfSzF8cqjEC6PH2Z
KtVuG1APRy6RTX/jWgWC3fBmzFhZ2HTrKn/CbhM5L8XtzdGfouEzZhVXrVip18TEkxGoAq0/pwkY
m4vJlpC631FKjZiw3rCSBIE0c9TmhA2LbaZUwJjSWVonAwQwU4F48IKFFHIaP1RIltbPykti9a+Q
ZnzJRPtx0uS+lPE2vONbf15kYRH3Fozpk7ImAphP8VUwiqPy1ubOWFb59WsfSP5D2BL2Bset4PBc
0NutNWNNtNeglLNrb6b66MExtAkoW7dxlUWiJii9DlQAnZnePQexT5RcM/4CWkTFWUY/I63aMQXD
bVKR1dmiLl0LXElhduvewnNYtOcvOPtN4L6jxEEr2wvEnqy0/ppydng4FmD6Vl0HD2njbr3kpEDU
Jd/DcO80HPByDRpHMf+yZ7q/AqOnuDACSVAYNH/QLq4BEFaiWJXJvS880VWcALmPaXrsGs9NFPoT
G7ylF2ZC1w2OLKsU+Iyw+ggcQNngbHvztRdLwNQsAS7Yi+gw3MqyZ2va+GmWSNbH85tW0TH35Ekn
KOSSt/s5SuFPJcGYZ8jzBz67MqymX6VdM1PAjtM258yDe0+ZanRUjAI5gVs4OmcmUhs6hcNsBHaF
vmZ70h4AeBBqddeqDpjnH2eL+xomQ6fIZySi/tr/HrUgwQYOnXKG+mkJ9Kx2GauHKLYeGp2zPXV1
Jda8R9xGIJ1eUxLIcHU0iYAIg/vTu/f7uyVNiCRs1sNqKEkLIzY+8vCUld11S+qrJOK5e1n6Iyci
z+Wi9BruYGA9fssNRZXa8LX4ovwX9U2kxJyt74oY4sKiahcaNimx+QkJYdNeO09nNz4eylWCyxPg
xxviJ4WLCERSGKfVsSFAZ73KpU6b7lyTdqtQqka2+WXdIGPXTdzy3uzD3/keHhY214qg9GD83vuo
F8K7W9Li5spHMm9j7OyFMBXfGqt8l27Ik5gdz7hthzCGNSuiQJuC8w2UChh9R3NXpAZo68hzRFw/
LBg3ez+oIQKTF4Z1KElPDMURpf7m8OWyMnkxF520a5DRaeJeJOqUpiUOELU1LHYDlC4SkBKjtAdO
JQfxkE3zNnX/E754PVMMBA5YBYTlJLzjSx6dhP3WGlNc50vnx+EPDOdMNYcLbfC4AshjPV7/yqSC
MXmEaIW9YxlDfEVH3VWcO1U8fInyOfONlt870/mUs0+TlTOLtW+BbOacwKtQ3iYkgiic4kV+DPSP
S65XFj1QB3YlzRBJ7D8TK3xdkX4fzNgl2sKgHHXB1WvpBeAe/NSnK0TDmIvrzy5uN08FeYe8KYeC
2HwLM1FmudEgUtvw8Sp04tk9ov8oTXWYE7sAd8KesyjEMGwV2alea84p5oUBUHSgRxrz1ZkkAyh9
PPqfSHtn+7z4v0pyGQz3XIAPdfndW+8+rh7DQkk65qe5chlHcyFp7TfDwvJ2qBPf0s4OkL9o8uIy
MygtujNMMD6MS4x+jENHaUtIckMKsmElRAOHL1RmFa49+L4CLylH4jBL3xbo1ZySwTh5mDoGm983
lhTIlW0r8G/PzdNr28ysFjbbEmd8lK9u0GqKr6MbjA4i4CghO0N57IX6OUKfuAhKYlPC+N95hHIF
Zz9vhI96Axq/ei8S7q22j3S00jTUEV3BfM70fD3X43/s4K07Cq6Ne9BwdiziRW9LvEz+3qerNlXk
zJdCgVWD52SlPMLAhuxe8lceS6RjHQkNXgC4bxWptkM0UwyK6dUbmT2rv8Kt2xcjoveYJpUaOXlt
GBBQfhTeO/eaCrImkkfINTJMA2ucWl6cPfxRpc0wybXVnh1EHQh3xoTHU2tUmevLPODuHO53NgUH
NBc5Iitnmg78LBCc32xKnJfxfWtpeRZ+EF4NSupJnqwVXvnstrPCyeBGDB5A6HYYGeO6dXRfwdFU
sK3FqIkzD+1g5AooGdTLAHek4p7q5XdkaCGjhvEU1U5d9qXHXKgg+xMatrOZqRNWgcVCVT78gZ55
tgxGIsvzMCMYVGoMM/F2C5HTZFUyA+QPfqXq257GVUhLDn+yAtIYpm4f/lWZxzawvikwpomRh6fP
FHBcbAq53bv0At2dNU6rxBsASPEJrqsWQYgM0WAODIE7wv7jgD7+5Rl3fpCED0v6SZgkrz1k3MVl
iRITCl38u73lhThKF1MpG7JTJdaZlF+HfNpud2X68+r23NW4uIWJjmyNKy5XLofdl21A4GFaNCxF
oPS18tm4qUo6QBVSaA5COxORu22F6l+9An+63Zo1H3jFdC9oYkFCPByCmAUXOihQAQrJ4pR6KM/p
n0mMC5U45xQc+JC3oaGlP+9qxjbjw/QHl9lcWxzZ9uyZgImdCdPFy5kIAcGIOVnbOQZW1l6CO3WH
T5OVeLXzVWaWsUCfAp9sJtAaMip1p62R5g6Hwo9AZcEZ8kKAPNWbWTyw7PoKbCy5ZKEi+XsefJcs
uHvQyjaIPkKIJAPihNmxFdrIfueLYPZ0ogEeq2+t6qN1UJcaAWz25lHgEZPeOodzfsXnWztV2BBL
tn9TJHBhc56HBIG9hPnexu6AaW2MK5Ok9ixehJlpJsJxB6RqFIHYocXC6c2+jSkt1M62WeB/gSG/
qJBrsBnNpTVlFtiOGpD43RgXAUUELljknYvHTIvJ4Qtc+Jmpyoog2+iRH393JHF1rPvOnwo1rgAJ
IlE36MpLv7eaZkS8c9F/JUNsv1hO6CcY7rzDxvmiz5lBXaEAsCzWuP9kakDrXrdg36VKNChifx+J
dbkc9z6nVLiwiCtLP+zSa38auzQwjRbfv0LggnlpP0HsCXGfVq0LYlqdZuNgZ6K2zb0UBwdUQJYe
mq/k+fe7cqf3WtyoEgS4mAGgedF+unWjlzLgYbByD/6mMBIJK5+G0xNW2+Na+al3w3pOrShrbGhV
QY16QV5VVfbc/IVezl0yqHpw4YX9mavsmgYjJTR7hN/ftEFC/9fEsau8FS5FNbF8OTOeu1k4DkLE
Mjt7Rx17j+PGVFG5xFJQFZuu1j8kvJgUobxxXwCTCSPFamSnOdSca3WO0NeOA18XzZ9zDbqXRo3h
r1nNbnMdB4aZDq1lV3HXYNqquueey4xy105rpdidlH+rQ1vZnjIko+zRBOaM1gcKahN5zIFN15+w
eqIsL1SYZc6b4GoIgt6qeEskBjv1QprTeeAuNpXzr3e8DRXCXR/jxnUJpBlQzlSgbsdFNF37DEZt
mJPhFXnldMsM8RMlAe5cekeLin9qD6RQhyNOlpqOFRW+LfLbEGje7S/DNcbhIHBuKWESx3OGnk9Z
2UDo5BAEx8lULndfdYOWe6N23K/C4HV2jD7kxJ+1c0USgZoG+aNHRT9+UTRgaqo9xKuLNa6wFVPU
Gym7XedP/5d6vZ6KQTnl1zL6WyyYmIurvnJgW7j7Jh54tlLh9ehWZ8Gh4mWPyAYWsN2r7+T+Jsv7
tjkmI+WJNK/qJNDb2xnOaP/jnz1bll/+RJfh7rb917o8bmTzPM5NLY23WwM+ZzbzRo3h4zoLvk0v
FW/YY2s8xf0YYsZFvwASG5gxEpdJPmjHVCGSbWGSh/BOIPk6sLy5TZppSuVCoFRONzp+mzhWvhNK
yvzcRTpFjI9mW2SwBzGtOaKcGl/eC2ND5Iwi5ocKcWfweUZjW/ejH//2asKq8P5ro+oYJFI253oO
IYXtwgv3K3RQNZAYw3aJDzU+PjMHx/rVpdWsP2Er+yZ7/T/LTZaoP/LTSJgBbSzuMLpa/4zuFOOR
3rqSwCw2WYN31qLMjyrT36TC70OuZfsIc36LFs9IrEzB993BCfpX4tHQIzCunB9TytX9xw7xpH5Q
/sxIt4jxcoModt+YXVmqm515RGRLOSreLa26urEs2+gkav61k9U9275iBM0Mxq/h/OmMEbXAdZbS
SkNb28K6hc+Db6preBocasua6Brl5RmAdUwfHxjl3ay8TTUmcoNLhEU2FbsnBloQaHF8Dersy1ir
3akjvsMX7lnQGbh4h7HsQN+m0OLmpJXUFsMISNPfWn84poCraKrYDfK5gwit3SsWXwE06EZe1U6h
R1kZGT0n1ESnMDjJR1LQnoVFiWt61rSxYY/mixyMvz61VEY5++u+KDzeMWsI9UKWWGoKg3VvLsfv
q7wumZxtahfh1P2t9L6NEyBv5zg0gB5kRlMJLY9a1hxEz5e+VNl/3WJig0ZgjdROv/uZSsTvTj7j
DWYCD+ObAJ8tahoXbdFVPobzb5mJNZ7nl0xib9XHVMqNn5uhogFRRYnnmGvJHVL6cTuCd0v5jbQO
0o9upr5t1jnekXgLLoADn/rTOEAwObTW5f60x+/pTjm2RG3RGvjwz+G0Yy5fzlbn5HE/Q/n+Har0
I7kbVMO3K5H70HsAVcApPrvwBjIv7ju2z9SKEDUXHhotduBPwzVtQGjcaRyh3JWEHfw7owIucxH2
DcWWeJF9PtYxh2Lj8dFMb9eQbH2geMmjmtaBJzaG2gQfoxMboFvKI5FL9zd8PH9BY8okdySM4WTT
tabztUFTktI77huWjDHWWmMhH1fQY1QjXCEHWEcfWer691vebd3YomTuRCcdz9odiqmLmHCZpJIQ
em2G7JZsalO2WmLqxUoQsOM8JYVGFj8CVZRVopf0LSauuOxDkjkTaYYxY+CEQWk+/tIGTkCHofmu
q+HOGDwco/Vx1NJOrhDv09aLW3lchmsfkcuryE5B5R/4RIkE9eyXa7tI0lqzRWapwdCe7V9YV/L8
0EfvRKnbiYVSGhQy5NDV5i8W+Vtu8TJVE3cZYKlDzzJzqSGa7moZ1G6nwBqpn8mTfff2MyoPC5F0
FhGtEMl6h4LEBoMHoQIlhqpDoEEf7MMu27uYhqyuAx/IebDKQgG6FMFYgKRFoE0ub8kG80oe2gTk
PFo5D4UEyd1QPkgGLal8WPZkkRwx4bHx5+fTMNgMKuOLLpTu1Mzx26ftfZdtyGaT5v+9NZKy6O5k
ukYuUXrbuPHQ7KzR5Pf7ndRyjfGGkrtnFMtkyrUWItOSe1uHt8wkeNj1LZxDJCNkv4k8iPk5OL1F
Q0bCNvUSAEFLcvj0Lf3p7k+h5zc7TeUzXmVgjdNmEsYIlTxVo2M7p/00ONUDO+Yq2HHy7LhbJgW6
Nvj7D0eg4eAZoG4AgqZoFcW1T6dl7TJnYwCY2jSReGbTGvFMvpDvy1w94WeytaVefk/MqaKAa571
PN5u3Fd5Wd2h6G4z6xB2as7msMQJtaUPVKIQ/1clk0xQhDZStLYcPL0RvaQI/rTu2fii1kJZkuyP
c1jkwx+4kmSVv8JVPKEKvpLPg7uJneJb742HaIG4GNaPONnRc2Flwxsex1746XBnfZhOLOEzvQPN
K/j44ovKx+9R/xRSoEy3jO2bLm6JPePQlAmb1bmZtU7VYpuSrNmR2Ix/mFz5ot0U5CknJYwmu3pu
e1rp+HSndKf1le8VIzS81ptD+GoaBLllzZNqRAP5Qd/02nmdOSGcE2XQU8VpfqR+V+dy3Xt/UtCY
+ww5E5ezqXgaEJjRShXYxt71HnXOnGfHH8yCOTr3ZoGvb0POCuqrTNJpxp8/4HxWHvISoMdHjJSt
Pi+xCv4FqPMkCZpBgXsXrnaeCpMzKL6RFy5FgpgyunMGcWuyX1aukbNqMbfHB4GoBN0HPEhvdBqx
r29HP9IxOfFRrzInPV6eQJESgll3LAe+QImfSeuP3KMahrxK3IiUm4KBWwmnobQNR3T/bKVok+zJ
5NHpsPwbmaoRvAklX8uRY/ato4ALvNudNULG62d/ADWGbbG0tFAdOS+80Z+PMtGHds3I32PIng9B
Q4Vc8vQIEKYwnxm1v9i+/00zfBNXHd2DOjcNV9r4XfkpaSBBL5wULdDA4O9rteHKa6vZxIHOcuK4
BnD0U29W1fIiMr7h0SzK01aP8skYAvaaahTyFRsMPOUsz1w5/wv+20Hpo9AqSrbU8UsffyPdTsRh
Iqe0MzWVBb6gVK4JBjb23D9PXlrlJIekf518+HHD79Of+LFr+e/fwez+HcOSimzrK6JwDuKhn7FN
h0Y3G45g2KRA55OjcuujZGje7gVRX3ub7tvjCgtQtG6rPSGsLkDS0nuO7zwj7KMYRJb1U10pNl3V
d67RFEhaCi9PqBIY8DlHZg36frNfTDcKtYOPM4GUHr0MXiXc6xfGDdof7IOymBNCw1MGPeb/rPuf
W2nckCIPRWw06//DPG0HlJFJyEG0aYm5dhGJn3l0kAVG00vrMzEBjbCwDA1k8ALR9GJT2HvTNjNx
TYvHpcO5R+XNt/dD435E0vsB/VqnFBbF1ZEPg/xFS63xF+IkmT3/RtJ/8MGvIeE6sYJJC2VT0Riq
uKh55zqDAJZ4mMvuhKxFeY9k/Mgaf9WPetMTDaZjcWZcSEzN59kzdVNs9EG2yWYxsg5Q7P9JhGOH
cbKpx3CWEs3I5QYlI4effV7KLTpF9RQ0nSZXXrqluf+j4knDjqSUESdg3M6h8ZqUp2q4xwCa52gT
PLABn55ktJl6g+RkgvsWdxmHi6JJrqkLaJXRed0QF+T/83pmjAlLdAllTz1F2GAW2XrsEv/eaW7a
HJV3vlepMNwvgKVYYf2sMGNxWUXGA5NXqYA37duFnZUu221v4Q5aX19IApFZrtb2BKHxcx4CsClO
LXpa4PZR97lKh4MsOlNN1rzvjKC4n35gNIICWixqJCxDe9oMTlBr9aBM4ZJukTYF438YOFRboM5x
BA0VI9ZiNpPGUAUd3/jsaOGGtFiOhoc8+8eauBD2DTdiqwnj/b9OS/cTWGhXQkRrzmA9x+0r34T/
9i9wKaHRbQmaiCAfxWIwOUmXg9SuntnapNq3wleYvUtuxaJiWI+t0oxXqFm/3IW4E+TMUgrPglPQ
92wl0GpN5KnFdo9rQbrWLTsM9PU2dyxtE9bsvrRXkT3i7CSPV8nhkdd8v13DQiNaNn0Zw5iQyPOM
Of107hXyAgGETXpSwXAtI4KmvvHvtbbX75NaQw04/a30tjsnWLIzAo5SX1mNhxBwK6PO44uI4q7k
b28NwDuO6p2KqLzLP6FERz8RIBJlZFHfOlXHsIQSkx6NxpDeQaznNXCIlW3CgfEj6cm6g6GJyhrE
QvZcDK7LuZHQqL1sXHX7xmTtixynQ/inX6Y/ywrYE5C6A9yd4Llv3+S+3n2EJOrRf0YVUPsZG46Q
1LzzVxHwFEdLpnyf0yo7sJZrEPSya6PbMXXSH1Ts+Ms++pTtOR7nCko+u3Pni8kIrCVyRCSjQWwp
az6W7UUuTvs61ho8ccadiF21GYeicmHFd0SDAAMlra4aLATkvuZpidxN1/feUn/kw+1FtwX73sea
+PKWiE9xFhdIoghB1RAvy5pmDy2XYkr9anFQeZJTCNhunLm9ZyNk9TzdzTdgIrt6xtlJbcJ+iTAH
6s8uImDgMECeDNxtryTjiSpVSPI8tO0ryZgS/qpM7i96HP0SQgxAFtnKL/64kljalTNfZxhr4JUc
ZoKSQyp0Qpl3mVJd9fIuMcv0m1aROznSjpOEVkP9IWNS62uHY50iZ+60qNr3XYENqaN5F1umDyJO
C4TEVOr8eJZCx1Vygzj83OJOne2A87+UszBFnh8SVRJ6/3PtX+oIQPoL1LGykHg1Bw69IO8/IjIT
DGHtIHOUCppijjH0+7UrGoCxIoBm32hz5LkdcMIb8Von8l7uWjlf32rKfKkQWz98dqbdEkY+OCSq
FuOc56ofLMoTaA81YEVH5CX0NwyspV/e1xwaKn0euFrbA7NMHCMTrDvGx5YaGyqijw9Yj7MCf/H6
JF9APetOzmnW7rabLV5+ZASBzNHlZRYa1Op7xOZ96HSrjwVuJmzQoNPWVPR0FB4M+AQFZblUYIiR
/iJx7/THVml/PlCdHJmFXoVQVA6E616Dgd4HaHfsYUTf94fHkBTP76WavepShfB5u+zEFiLra3Og
mIEvozw6HH2wDMr2WNr2eOJLZ25K9Td6eKpV7/YCjfLz4h8piZNC2vuwJIsXCihA01P2SCYbIc76
hjLz0f3aMRov3TQUqcrQ/aUIJijtBmozbAzzdi0eI08056RbxttnWtNbMhaE9WZBErLPw5hpzaIN
JcADs6iMtISkVcXCoOWKb5nXXPPmsaOfOpOFqcv13V9CWzzezP0f9es4e31Ux4VtxmE07nomjIjn
j8qHOgQGk+nRAQqAt7sVXUK8ya+66bWHXhqRGNaZDeKHaOK+wm4wS3MvagR3glnBEJL796qrCGjX
SYp4FqgFMK3yhC1SK9Aq+tztM84HvsOe/dYRIMhAvELBSt/s4fPzV6FOficlMGkHyp7QTB3SKc4E
tV4idTcSjh1oW9Okb2+wNSzcuUyT5pa1LoH+mBP2n96nIBz+d9Jk+F1SMkyyOPi+o8BZJ+AL1QQ6
0g/euHuS1GR07xqVrJQogLtKzBPVJWYnjCmS89mrhDwidDbuntkxvJ170Tw5XYt41Fzr7akzHj50
Yvt7wSxhq+DJT59M/EqpME4n78AmRoBBZtikN4xVH5cJMcKW6k+QO/jOS3nD7+JSXVLAW5h3E/Jn
F1PKH0vWNNTw3Uo2QJp5ZFpEIo5HeR7MUuK0dWRo3mGQrD34+iIJ3JReitCH/OBAYEf9bPJNcCyZ
hogf8QScSBzn24Ajr9xCjPpbYlfdo4en8g8sv3nrkGsI1OxFJQNZdzyZOY1/Y3NqaHDST8UzE8N1
6Tq6zBvtVsovlP2sGcwD8QCh8+bHRsdMTJH70pkhhZqhtDtU6Ci+xURS7CcUoTe4H7pctV/OgTkq
46iY0WhYfVuMgLWCHgYiIoQ8Mcgsozfj2zPVQIuYvzN/MkizUCw033sXU5dPIqPtgkXK1xGISTf3
8ncZG+b7dsZhg04qp8oE+SY6haZECil9bH4RX1LpMu7lhCi+ZVcSK7EQZr5Mwo68Eqlbd2Yyz97r
6dRh02o4jWIO0NR4hcTvw9Jseh3BidSN4DIFs0yjDXupKrUYumxKvfmzjFxdTHNRvBUD2gDyquBJ
OvGrHVM/u+d0MTaF8nZ69mQRY111v/HsMhPVc233gZL3AOLDmzUWCd69+csTt1L/2bMrxtBTbQyQ
YYSW9ugPZzcn6MFq/W5fNLGOaSnZuN5ADG1M1xfBgHIp+iq3FpD9oFrRg1FEIGeaeMQfv5TIztVF
HGA13Y0Uoxsy7BhTPjWeG3l/BiTIoxZRMkdfmfnCGlX5OyweUS8HgwVO5tuMvkpBnTuXiHs0Gw82
ZbVsKjOuKeIE+PyvREH29cIZF2a0myaKWVrSaaLjTC9Zb7cFDUOhImREyvRhHcES1D8KnnnKpMP2
vpJJvAod96P3q8AGS/k2KvOzZ5C9j/6+F6HxajIyuNhZY3lSWJaEhwIazdJofxt7y3C1K3EoAZrB
XNFCTJsmZCTPj9Pz8SaJoKJRO+MTwlwJUvlzJi08FwYHXgaXMBIsC6nEqWpPxRbv/IOpl6GcIHHy
sSL3AYU4rg5gaAHXISF16m+ZWA+haFIDtjVCUY3L5Fy7wm7yxqQkEjfSY6uGi0lAO9bbt2IGvQyV
gpZEpYiTIsD2fI2tclOIRwK4raF8uQYq7WbsAgbwj7ta4/BId2mEKNTIpjg0/etVNVgQrSTb89ck
s2NizrnFFGDmaIwdxWmM/ue9T+EXKo6BQfPB0fffrdpHaE9FX879tICa9jfwYdjkgqIna4rovkr3
5TSN09E7yJxxACN1XSoWNFYtPekT6HW2Tdf+km+opi7iah5lAwUNhndGbj1mkBuycNMkOpxgHatQ
XkkYHSgEUUWsFOAPm/9ifnTAE9cckwCLKO0rV5hLXqc5DQsBygcEeHOZ0EdU1phQ75WK9oyP0IQr
QD5xMrxIznd69TkUFN5LmlECUeN/mKAHwAW8zejoly6Bt0YYIM8H7um18ElAEY4NZ6oWhC6KUX3E
Wj5jcYmZ/cOI+tp+y+qFe0GirPEKneYVpKNrWkSfV1Q4715HBdlpmaipsahftHbzm2/0Ga0+7CfC
j7aUMPJ5nQht/0EFbcmFgQstrMDLjJqf+ppfxime8uzhKBn/3m4IfcGkpy0p/toqSBrZ3kN3EBld
Kpz5fFxxNxmEtC16EJaB8idlqXYNBAZFO9ZmT+wflgFGlxUOy5WoC3wAodeB7rKFijxI+dEyLYIy
wmBd9O9eVlClkB77csTefG0fpRkMAIRMzZlaF/Nnn9qU1kWRuop35VNCO4D0AAN6/yy571g2vOc1
1hX9CiTreEc8bsyqUtVtbG/0KluHAtIwixiQhJ8QLImPscrEh98DpfRxRXGR/r+n7iM5In0P7HUw
KCWyGC6vt1hidKA1VicVIMKC6sSxF9J/sTTWVS34/xbbeB8xSERERDTAwuoPApDC+wNoaGR9YzfX
7/cUUmUANAqPl1feBJasoFeXo8EG+1pDrCARRTRzHpYtoUklByCxxY25VRIqFB8bWjec++oxdhvG
h+qoPC0AqRLURm1n2/vMPKrEiK96tYc1fNDZxbh1c++Kdu9pkqdT0Ep4Ym0AA4ax4bA7xyZIpZ3w
Dli3LSVztV9zmIFY1KhvNDe0u6EKWKvHb3ytNj1CZtGhQdZybgpr3Uc6xfC7PeRIDYUpehKMoD85
w9aR8+A9P2aMJcFM6cvW8P/J9xUqH/QlnzsM5nxcZBxcn7NeDueA6VXLwdyKWobn6mZrww+aYkFF
U2inULX7IgEO2/1GDHoPpxGvW+aI4qAhJDNsqvwGp5c5oFX4PgrdHjv4JDom0KNMdNCHobMkVJoc
M4cIGzRKMwaYbUJHn5nOzP/91Qj43RRaGWOdwOUeFrxguVywyPbzbt/VWWkFPiypQ5bNhrtDdofx
fBpPz6gYS7NoLYqjfPuDsLgDKqw2f8kOljRpYGyvLWpqxSXZ/j5cFKHM8eELCDYImrGc+naJQ0FQ
6P0b9R8PumcUG5GHz2DJqG1mug6y/giHTlD4TmQnvvGr+htM+A7UKYzMrpDtyApoRRZ4C2/HaXTr
drL0Cf/Ch5e1yUNU9YHObqxDBMAgOpdEDQqp9AalYveTlE20G1Kr0hnaZwm7OVrITsZeTVG30gOx
vP0TXsGh+VE+lp7qHmq4vB35ibSCA8QPDEFkVX0kXZNg55/p5AvNgbX6rbR1jOvVllsavqAuje6G
+t/hG5wqTeko88f5hrmcL5Mm3ZH/4Xh5ZnuhZD8nExl38U1Lh57VQCfYrMJd7/hGAhqbf7c2rUs2
JdoIApSV8G/Yz8iR+GjcbqtqlPwhpt8wrT3axWbslEPuorNsM+/6HVBkBhk/7QkytiTlArRpPJkk
6UGToha2dC91xm8LUYp/f64rqpPFqChzri1w15bpVH7yBDEaxlHPilhujGyR5wEPlTmOyLpEQxCj
8JR3lWDbyZKx90R7P8QdPHECLpksncT/+WJR+vXXd5r3Uz0l0akge5rCxTmGhCY62ReWmi4V8N+E
LJY2TPOFgJ48fdWE9rpLDhB/hredRFWcSSv5Uo9VjGt7koJAZ0VK6z6f0o2lRsz+LhC8/p1qhyg6
+SYJDgGJ7lvVvO7fk1Z9EIYBvVEueXNnNbNxn9OG/zvzJfTtXXKFnECV/5l0CwvwrLXWaRxUmq/y
KjIRKP8aGcG8umrF142EhLpm8QmM/IwO0mkw23sVLJOSSPuk1yzxyK8t+rZ0oZsOJVyWJ03a7XQa
3DVvZNPKvbxGyLUmUqdxcRqgJUnlxZtmNOijHsoUjx3E+dHTB1DKYzqcnv0e+XQtGyrF003CcAyV
V98cw6NXuV7w8poYdUOnDf66O9RH+SkqOtQ3fhW3JXPiE3cJ6ou0w7aVYbhWiU2grMc/Edaq7L69
UGOYhXdEyPMjQZVTOjD0NABtvQSHVm0RnEXSMzeZQ4Arrwv5P01cbI8FPFRcTPF376i0SkBMlnD0
76rU3Py1A3bPdl1JAKrvmzI4dPDWj38141jZdzyDwSuACKUaojvR736SgZPuA4OwXQo/f0m+5vPY
tX1ChHYthQvmwfsJ9qxS0xulMNrHvrHr7K1Fn0+NeMPaS5F6fFK8srQX1dGR5usNlI09oiTFAmz2
+x00A6kZiM2PR7FKw75yGE5dLmJuhxe0M/oHeN8e0Zn2SIx3VsInxG0vAVklthEK/I2YJK0GKECD
FDkkqDCy3950EbSdDFPEfZTf2H3jMdxoy+se4c2pSLE5NkT8tABtcRGx48NwytkB/yg/T9tRgvTt
1LSsYEECpdntTOVlzMiyPtJmbW33znGVM5qC0NXg7MFCGaau4kMncF6CEhPtKy5WpDXpI3OHtNA9
ODXOnRhqwfoiqlQm4QGNITuLlj0E1R3196gT63XAABS0HPzqIo551MkD/ee/jRkJStBFaOCuNitF
ViRfBC3KJEi2URM98X2c3xhO4Tw1bgszXL2/rBYKYMuqY4zNfTQxPUsCSo/JyNfzUpggEnWKu00a
FNi94WDTNCtcAnU7g5aaQRnKSTyujlGoj/uDGJrRZcOfSv42twKWegQL7kgMdekiNi3xa1/bwsz0
HQpydfA/KmlVS7uA6F/+/59CQbgVpt09SQbdMYZ/vsoxv2aub5bP87rgiL+5jE3oKfJmN9jTt+T5
TCSZfbcZiOPxjuZ6GpGukQuwThdxfUw4BTQmVyVauoA7nD0HB8gmHiQvGy6djWOwRdCgLWSzvogY
PEaeYXlw1ZiSXsmMkQd7B/iQP34EDCelfGTRUKjFtPaxERDmT1RGSc3rU5x+EbNCRMElFSJ/MEpt
bRy0n8HhVd4F/eLrVB0CJv+wE2TL7WXFvOIKTRr0575jrP+YOT1J+gSq8lPPtv9Pk1pYNasUyb5V
QoHdn6gdyZOCjGuH3c8iNRD8XbXJsv8itzYsHBqQZ1Hwguo5LY9ZCijI+f8sQVOzBHICqh4VV7Qi
ChjzGfSp3XzFh7po9S5NHDT8pdKCxGm6RMuLtHhcioCxABuakwwykC1eL1QAYdN6SPjNyJodEHYt
jj7jvtRL05H6BJG04goR2rL+4/pkYQg6sy0oL9x2riVdqPm95M/ybQV7sO6j98unmVlD2eh/yYQc
LkSB8Hdr182FMMigigpANnDg+ddKFY2nyEzw1isKh+YcoF4T7Ikxfau3wennxC2cG/pUo9yBUAGc
frMlRsTm5BVnMxIcTskeImVsYZ9HL+J8KDXmVdeOZJloe96FSdQ3sur7Bkh4ZEAZcOcqUAcNVq0S
X1QEYojabF7hK0wCaMNb8wvBg9LbdOwUoxQuzFFRHvS+tgU20ItOWywpqnAIgvBtqDet6RiZTGje
YfDOjYtoKTKurgptKAmzBUhbP+VMPRawd6kTK4n5yFm5VcOfUo9W1us63POLJbgqZ0BqP0sCdvoB
AD6VvYQNM41hm6LtwvySogNubx5eL8SLS7Ip0JYiXcgKg8lghyBytaxo9hU4SpWX8J1Gi2XLgj6l
tU67QfngbY6u5gi9mZkEXGDMS9PnDT6o4kw8Z3BBUHot0NO+pMZtMtf7qsbV0886FldPIvepTObc
t4QMTP/mbAyHWlnWuNbLKWkeWU+AYGLSNe3nepLWy5GQSfQxVravfbJwZjtriLFZTnfvT1j1oSt0
RpvKgT7QsKzIVvrhct2D4LaHx2cOPua/EIMKihf69X3fRbsuuRt3LVYRDIjMUVfaq2LYQtzMv3Xk
TqSxZf8f9Bamid1iDMACdhMJe5cHTvPCvP6AQbcOFQ5wyqGntHmUYmz4pALGnR+V0/3I29asp0Kx
mXV66N4qbNADwQ6Sqc0bjRpdgUuPxHZJUOVn2QQzQF6QM6nWxL/MTkYOGTJhAGui9IKzPlKui9Ci
Oodbg+36rIEsvo5rOyuInnM/bVeln/fDURreC4iklxl4dnjB6QfqTuqJRJtVE0UwwoaIjsWopMA4
WENBscT8P/hiJu0WZWYutagLyszBCvdfhmRhh0+3OPupUAGXAiRlU0GLhpWexAypVaPrSuQFf3/v
KMTQOiQjcZ+bwoSnvdvMiAUvykvPDOlA8q39e20v+8YRP815CCs7vQH535RE1JZBIxvOua4u19PD
lsvgRQiafZpJLxI0hXZDGhgrdpLLbEk6Qt+X72gS7DpGEIh7h7/6nSWRDgIuTpbDOa5UxLtJ8L40
ibN3jrZfBFCR5O97rpht2s5JVMMuLDPSI4yGbI2X+MKJFEDTxltvMLdO0UgjCTuSZFHLPcZVcSaK
rtWk1Uw0yQPidslmpE/Mw1YVVMd31LUdZrDTKruu7zELJ1b4K012E1sSmrI2HSgpjNnSPI2LqdYK
fO+L7PMqj7lYZV+I8PzuMIDXwhvcb1vHcZK8NgbbX+HbTSPhOMTA0pse9jvLhTMUdyylP5sWv95l
4xHD8dl11A8jU2s4tLr8KA59IXeAaWDlU+sCqVhXNWJpJvCN0fdKkypa8BQAsI+MwpI5QdYV+Nhx
1ghBnxxfwexjnAkmfCwdbqKhRJmZ2SuXa1ZA9mqXrUc3TiVLEeTgoVzfQaR+TYRkmVE/+PygFICH
ptmsSIr1ywJgSvonLnypI0TW9wTIPpM1TnVMxeyCJ57o/nCwUi74J9bc1XlRFNQ2PlLTLpfil1d6
7V+Z/BD1VBbcqRE+Zo/nUmBPOBbuB7DO5MuP5fB1wuXIEwI1372cYi2mk12oZSpYAdNXxsbunEdv
DSV8n/9ViYm4T2Og9080ksYcx3TRucsrESerp6lTws8Cn/c8G1CTfO2XdeMxm4X7lURN0rttZ63l
+VKfhaP8mxXblLT7VURd4GBAvAaD41+JJwShOMiJmx+thotsfxDi3UrwBizJ6rNOEo0EkvILHp9j
YbMkumYJPVVPmTMRoPzlQ9nuKBb4tyNMijpjFl5Aq4eeBCaFIXbpqvLN5caRG5FvHlM7Ej2Ro3Fi
ZD+/pSeRy9oa+eUgjg9gptePxhjntuyQId6SofsO2IhTRrokQyMFYuJjneuZJrtGkJtmqC6UiUMB
j1QopjT/FaxKBoJ+mOJqzwucQR5TI0Ra5/8clRBtMgwFBTVaIJ2YsLCH9Ki30ef/JLZfPUgdvhbv
NYbaFNT3XRJ9gAD4C6i1uPplgZC/E0wURzMDfJdTQh422yaegsM1++IyM0TisepcfEG+uzYtteAe
EVgZht8CsioeY7WZhpBh2uBUGTFOHI6qOuQuzsqXCQWhkaTbud2Yg9bbRcC7obmwyhJQ8ObgvFM8
VcqkQbS0WiMJr1Z/+viZiW8Z4i0SUixVSK8zvPwiMrQPGsZpT/tWkGArpw+ILh1OpObQb5TFXfqq
n85v3V2XEf1DohvpuxV8ntGE7FvsRpR6+XSrQjPEXxoY9PDk20Ov4I53cYvA0qBsIkFNxMI3FAcZ
LMqSalKwPwzF5qKwV04OAMozGaf0Zdz774dWJllTLnNS6yWP72fm9OCEk4BKy/vtlZYCyq1xpbKE
lrNo1LElV83isxmxUCuseLWCl4iPv6xBD2qLegoNu4jz2HhT3GMy8Zg6tPWGZKN3EJw5MHwQZIXz
6gGptMRMYO9JueSfNpTDI6mVhfwtaq3MT8TA2xrmt4eimNqVaBBr01h1OxPkFI9A2AWF35Qh4KSh
Kpbsy69M+Gtuu2Sa5ucowrEboj9A48c2U18jQknjzAWmt/dfArZ15EZPvhgvGvC6yqSTlZYGVEII
dnfeLdtQ2KolKKxuTp2bnU9pePNof1g66qo3AIsYmJ/swyaZ1cBY9uCWcMyLsqcaZloxBV3epwOF
XTdystkUH0zKO8RIkSSPif7WGyK51FqmHJlNXyZssqbxv81qAo1dkHwwSHgvBTYcu97VZwlkKAMk
zfoT9fPa4P6LDfyunJjaRRDaMGvp+mUdJZg53kiwHCX5GDui4Tqm6UBfEEgJsOYAgaxtxNYoIcgN
P796qowYU4Qx9yRLPWCzHHQropAYS8wl1gfXvPCFc04AVN4pC9A0DkemsTgOxMj7OEIl1R+mNEH4
qv89Sz7kUmyBFNAneQt1tBnlcN3SLFhuSsR+beIhll8RCmqezhyP5w6CjX942O2k35gqtk6ddBkT
iQeWndy1XIJwoJcZnjeYrxH2EGvMKkvtDTsKUl6h5EMp4/x9CPTKpS7F0OinIVuS9reRZ4pI+hzc
lIOpL3QEni9kJCFlpM5frke49PwHiHF9499kRihTy5cZPJ2zPIdCm+0nrmOzD1X66VK2ff8nPGTF
5juFCvzvh6rrnqrlpRNhpreWSvukFH2yX3q2L2VIWLBm27jzq3XwOgg5/qy88cOwBxJJiU6rwYsT
FIM1bj4XcuH7DNM1aEOjmw0M5i4iyix6BHyPbBzKGnp1GovLucyinqw2siPd+QmzoQ95ENWvsIyl
4ekC1bWEWqVLwtq6tlPL1ko0hIM3kbBmMNUu0AfdW8WiMA9UjeY8vQ/3BXNiPlNnS9aEr6SwXNWA
J4vCaqZgLsJKviiXRXBYWBXyvbPQUVzeymaiEP7Ifu2+XHhDlGRgOkHT3OM8mCuNc72b0boY3Yps
B/bj5yBNY1AKY9KOtdIIlhrGnG40uvKXALAmw5KwAZGHYvFJSuGEY93317fueVngiAMBfo+fYFsy
Xj6cLkTPfmk6iHnNLDvIp5QqcIVwLEHZjbD/fb1d22ulA90UGTrFcJmo3OfpBfxrfBv5I9lwLUvU
G9f6fDqDKdKjTHa7CNo96uEqv5Ax/MuF2ouOZOX5MKYeNWf3Y91xZkAXG8dyAq4tp9ksvNqIuECN
NIWjBQEbLUnu6gh0F7myLbVUZVBFOWik4Ilkez2mbZD3dRjeJD/Tymlp+JClxodpnAzGJZKn2oDa
3VuXB+QjCJ5ZrfCv/VmOVBGxUBlL4UWA/iS2Rh4kw2csxMU5F/CB1BLLAEWygEwBjlHOf5BlvKux
30SDk350TbV+rkCBft0bsxXlh+9/0ODhKure+BPRfPHyCDEnfMj6JlCDGx6hefYerLvvh4JcocHk
eW3HYSY/reOj9LNKTGyRAtOAih1exCjbTck1fZkPHsLBB9M+jjt/txHwORCei3Gza5iNp+cONnJ+
S1dRhYnL7xRFsBmZBDIy40+1hGddlXs/XN/vwI3vpUvGSqAvq0eJ8Tw6B0Qu60tH4d3b4BJZzkqc
3aDrwsus3Gg+WDi2mD0rCvpsvBJNPbHWsiW49J3EmABqd0OeMkJfCH8B9+QivPmOMVmoPScTjxe9
dlWqpbJqURgqm8SeDKK2iY99Z1nb2j6hOIM3eTV2cu9bCWJRpu+1mTcp9yWvMaMsfsgr1SB6yGKL
LkXP9ERonPTJLdG1ZyuUro9Ke1Fxk/UAn5StcFEzv49vZOEqz9wxVVc2x7QGT9fNE351F/EWls6p
2F+ujqkHdLL6j2WdH4l02Hf/3tGuCRo/MzZ0Ucpz91BQtFBFqx7mP962xWvztDPOTMh1Mo/GGZp8
PbgkdrFQ3J9Eaa/1PIcHRd+kREa6olC0SfPHctRM/i789vud/p/YS4lPdgVrajPUEWxXJcG+7R/Q
g+hsO/nx7eUvbYr4paH1f+a8E+61Q0YNR8e+ZjIUT8qVgVg0KXw7siBjtbeA3pE2mSd4mCEpXuJv
x1lKpVunl92C4SvddQ7+mk58735VjCy7Vn3ODkWY0yehSrcr92QvyQJ7/7VJsEpdQXrCDmN8jBAj
G8i8ACJzOeJYJKGoMujwmCoL/RU/PpmzmXz0JnDErjWTPvVhkbKzZ/tMUy+Qm+1CPtEVbESOc1jl
9UcmPql68MEPCvf9qnOh6tJHPcPAUw3ses+LwufHaFN/PhkyDquBM//gYKhi6NLFN04DMwbSlfzL
dcP3IUSii7I+qOeDHf9sXrCMjT+RiHuaVx8b0Z4yHL2YVvjCf6VDqY9QsWwO1ESH7uQSFRkim6tW
XHtC5JzNkAv6ymGXIpofWe81UEIW1T/Y8cImAJbhI4wG355eV6vkXjoUpuG9ydgRp1NgK8nqYXpl
8Ni/Sl3uDkLi4E8QmlgfR4+TvfFj5Ta9cf8d1BLeTKxLQ4njrimN4AoqMZVeXHjYcBDD8KCDBRaL
kL/k8vAPt0sW4xC0Hum/foF7ZSry3y68780J6wUZ5BXdYVDnBDx22zS5HG7bK6XGTzgxO9Gy0vV4
dEsasALf698QdxFBCOFamv9/5ukTy5+mQ8Fzj167kjJOMz+pgcVfD8liokHAajCgY/1Eqf2vabIC
qIiEHR9zN+MX+yHn44UXN3c7pOadML2hPt6EQPvtoVbXwWQXOsdklkNbLBTTqLt43ICtMSZn8/KE
JIGA+S3tbPiDcn1tGswu1i8aYsXOHx6fJ81y0700MXEgZ5EHP3N1+8eIEIIG+ahWs72z/O6Rq9lJ
b6Sn3DScv6pCro1q4gnm9xdfLEmsW3V77jKg8sOxujx3CsyZ8DRiZtGlZiuy0VyJ/dXVgRTnuXcq
uGktyR6itSAo/6mAMct41FmLdkD1PajRx1HaJRoWIEPUDMhkhcPgrTElnp8SuIRUKAdc1m+PZJIQ
o3M7XeaoYAMrTy8McILRWASCt0XVTHnIcmXe55jnH7s3yeUbKYzo82jEhKAmm4vXEuUYw8onqjuy
J77d/iOe//dusgHMSSEPKuOR04bYkmF76IliUbp8xuAeALD+t594NN5l9BBy+cxROtVw2ks9KUfV
YRFgfrYHMpRTlO3yrsFSapmTAfanja6okdhtk7OJ/wRbiuDydwF/ti+P89ERJHC+raOBsNqhnPgb
q1mPVvC3HHENZkGIiiV47KDvYSSv3cm5chLwbMH2qfNSCs5zaxtdVSwmsi2ZynQceu98N+EQuvqN
euknZcbZWPerpuopxybtun0XxHXXZKCusfmeav5wI+fR0JkiCkitWduHpjntAyodKMY+kcqDHes9
8vWi1JQrjwchU9+MHI8vqusVTxcBuiIiF+aeEUxg6HuV9upRIgDlVl+rgFqxpEPSMo4yz8kbSqYp
KVQbTcw9EAli8nUx/LxCuu8mVWjn8Q6ZOW3BKnHKGdPwyDKrUsPivwCE8nIuzdWjSGbZsUMsAOXs
yP64Ghl45oSWvpepW5acGizAs2K1zf78eteGCweqV4FdEK4WR63/ABy3JB+P9UueOeptWJqpXxTk
P/MnWeONC+3pVM/+/kwTEk0Kyx1WBt8XYyBE78Nooduy0yzBMTfe+NiTVVy76BY/LN+8PJotu4e3
Wgl9Z6qNXszqJYEPU5v+m8qmxKC5kCAp2JLb1VYFeYeUHuJMpgZwco/911C7/dO00RY4W837uuAU
GzIjjtgv2/16wpDnr0UNwwEJSm81ai+P2YPDehMdyYtX1WGoFuafNbMzYypTsmiy4pTmY4P/J331
QZ6fCUSoD15VTxui/Bt3BeJvbbJZP4gh2X6KAwbv380f47aoDihZq/H5Q+FClDswS+5K54r7suZW
zmOMRTM6AVm+sU4wJnie0tfQeaARHqjjlp0uUv83cQRp+t1iUXJpKwGXQzU8mZTaIxcca4qinCMJ
EzCU3OJnRdgx7MEqBphZGrMJDfrcLAybNXL+R8xWC4k0c/Hv0ti6wJ9/rNDBuqwzSlmGCfGsZmnz
HeteYkffx2xuSTAI8RQSf0zQvhszB+YiDBqDN4hxq9Aic0of6XfowgYnvGSpFMs/9VXTBS/wBVez
ttkff+VFJ+eC3nPd02xvUch1ZcwJzfwyWQemJdGNlf6FsRKNoRXazR3JGzv99+G4TtULuSQ5TwPX
FDg534fqjEeJRPpAUErGEmiTq7+OfJ18UFA1xB3XMKHs0bnRLQJhgLgqTTva3To4skAUOlE/qHR0
NufFiMHUhKYIuZ9fHzfu3gd9aL6xWn18K5FRpIEfiCDOw7YvcuoF0HSlv9KpTFjnlQTjokqwyttg
NqIYK8cxkpqJNBGy1LiW54BzUUAEKtHiag+4CVcFeYH6xCesCNNnKG3o3tM4+eVPoxNX/MFLxD4Y
XUxqeZRd32Roh5SoTT0azyvHdw8XmllybwPGoqNZGmkwX33kFnJijEkNLCfIvd4Pfb/YhSLhPC/6
mazKo4l3DxjwF6wOiLEP+mw+dWSJSxnGNaSLC/HnHlVauyeTtNMlkWNBP/6SE0rG1u5s5P7Bj3A+
n4UlWuQ567gOczJF/gOUUtrVavV35Kmbu7ekeBPT71vGfR8wXHvhdF5gdceQsHa6RsqUkqrufnkR
5fPp9NO+yHm/VC62wLrItcK0aN6Eyw9CCQBdsGTwPIXLD5S1rjE+xfGZPobBE80Yw0TdtVwlALhu
4kY0lP1BzIkfOya7uzq80shxwhTti/zu5yFSADoPajcmta/gS8cT70l0ZVrpSYyw1NPoqhjw4kWg
NQkGIN7Nk1L+1LUvwvPbFCHCX+rJ8I8Kz3c9upCOGSCRFgCGSB7UD1oicid1aPcW/UUSnd94swUy
7tSANdUNeE5WiZwxHHYSd03fPIQAKNFqBJ+rfa4EKsxBzrOHgrtr4eVRrjc1k1x8S7CvtJqZ9Laf
6CQ1MYXsTdA0OoT3jkAFflN7PvWaI2DW42E0SNH8HLG1HAFR1+ANnB29v0+P4AQDi0ifHZvlir87
BAKXSHb8GYihSQzwUtL8YMmLRNLbeGrjrRoI5G2/pW/la+yCg17W+dfPwcDyD/UFxUxaHPzvYdIh
TB6AdWWOvB3RVLmBBnEHC2rAtwHJI1zNobM451O9ttBguL73WwKaAiRRwkxB/FBqWOjfrthu0W1f
3VwBlaF0IYL4IpeUGw3rQnyMY27kwKiP1EDrE7iIZ6RD6MQv+hdFPisjTMOVL1xU1PQRMapaZNFo
6tYvSB9KXpSEKE1A7u+6dlRJMZ42mRAH9w3Z+aYnCwk+qqU0vwHEDbwZAqWOI9mpkhbh/HTQsba4
E4UC54Jp9vXY/WUhXOCDfcdVwqyDWJijoGlKmYz8VEBfW+6DcnlLQcAIINYs0wnnaq7Yn9kI3HvN
JAHph2GSQATwy5vEDsUhB76ROu36Yxe32KX1J4PmhpM9BxTvc+nuBgtbsV1103gLkU8tSLibbe+o
EiMSx83wCrdOKYJpxaGgVu3UGwmdGXNxV/wKWbKPfBxJnVkV4otAvtxUOnRlZ9vybnDs4bsWz03z
/wPYRRx04xRqdLQoonArxGn86/xAKRh5/jhW1hH5jmix2MtmCkfDiAYHTvXFPndyGoyDl9wQ1fxb
Q8j/mNnhhDtwADRN9XVXz/eXYnB/kGHqWid/JoR+902vCNcG0EAJmXVh3M7vLqF1dO+VK4+BAasG
V4hrYC4qEHfQF5qvVyOWf+PWoAPeQHHBrdY/Z/V3rjQ2Txda6AX6HjzHcCrGJRjtg/yXFG3dbzDa
6e3IuLV2NYS5JBSCeSFo42bKLqi/L+ixTTVGTqUCiW/uCglVGS8rNzxx57vKJ72lccjZU0T4R117
vkpfF5ysVxtCp8Wd7Yo4F3PWpvrTUFJg1N5h712rdG9fhm3YbWu5fEdl7yBrlFRpx7Am+3f/KQjS
ZkAmp9trI4w42XEdhYW3acT86CGyqXLrTW98F0T96gogX0ruU3rVJnOtCzytGCev/aV5+im/UyJZ
bjS0fRJ68/4BfGTqIRN2cU3Spckt4wBVR0v6mBdV8EIrynMZznxdSfnXhV7KvK7WQJNIyp9mNF5J
s7zT+992PRtZ/ikCyyNLdF/FcwxCRz2cWXEFyTiwleQpjpqAdFoj5KiVhFLNw4Jo8ESMY9Ifk6jP
rgzWrutX2Z9wTqKVfe5tjPMvB1TMBaEYWDOOA0SCOtqBU6NQHehAY437+7j9wdxCxaHDkvyktDv3
/Pezwj0tjihhOmGrXG4G0Usj1h2al9+VSA/85JlmMt/hhdSaO7g+R7G3lRVCCUlN21avWT4afbHk
xlrE3bMZ8n1Ce8382rf2a5COTEkwbMv53lwrT30/Y6c0eKP04I+3vex4dFVhlEluodGpWmg2wZC5
mF/kNoF8p5TifFu5nl2NhBHu3VrhSBtrUBKMQEqS86GYfVtwfsf0unFBmCYSTITh7M5q+MwYjRWA
mxXnhJkoB6uSSm7NukvCbfr8jz0jezRuB6jw7IgsEOvhjIjkm3ntrazDYJQ50WtVbybDkrJKmmmM
IrnWZtjbVE44dXTucbpPiK9+DKavg4wu3r7FgpO41+YbVC2PEN/SL9ZtawH5eowIUNqcQO6neHb7
2dUhHmNEah//lwysijGH63jCrXFkhE0huOKeHdgkznWZL4TBCG5hGpt07iZNrkB+PIiWU0Z4eXx3
vyP/1pUnFu+rKhFlSywRb1mnPnW4vSrGSTW/Ro9t+lO8sJqtaLEkF4/1RbcOUL4H7/fNdzPtwqnn
R40QVEZ5P7GFP2HyY5+Kl53ovYCuEpmYKw9gbP7S3ajq4U7qoLc3v2J5HCh/Waghw6hYSLYMeiw3
+WmVWaiAphCOZrR+4frBdiJIKUPW4B5arD6/j8rFtWvvi2pF0a8eqbswATRQbO4h003c+IL1n/5f
jibXiSKTVdcyzjzoiBIH7XHTDlc4niccSCXks95VEA91ae7TK1NFm+0c1X66x+vEvDPjmk3oWdbq
Xk7TaISkY38CFoX7VwG/sTki7fF1SmU3AmJqgTmSkNtfe31GdTJUUIsqAgqUNKm5K/Vw6G6XhBfI
/TCuQz5jGw+dHcg4C6OYMwC9vrhhyeE66rWfVKYVWYk8y+ySy2Oodnf8B1qcKxuNIzOZUmbSyacW
Exdwfl3xcpiqzoK7w66AEH3o4+8ppNK/W9JuB6hCaDwnLwPqzt+HVl3MEvGihLxbGOdgJAjRdLRC
JkS5/F8k/t+UHajJBgm22AwLQu6RsTv9Hffbg5tGMKc71JmTSWfLW1DYtSVAryj3fqR6q0E70PK9
BaA1oEeHEkEERvau2HdMEs1v1HBf3LAee6JO3TBOY3EfixOFsBP7L0scU4tw08JAnXaky0VjhNR0
HH06+cI5QIHRd4nTMpsI1jlTeicFeEtLLFvvhwmffvAht0jmU7s1xidDRw+vq6S+B5Qewo7UlDXW
3CQkad3ILbVdkFIdkmLxn/3rl8Vpibaa1TOJz2INZNRH+75xY4/UJ5FX3uLT+rLwF7DA4W2p/xGL
AX7HpyJUgkgB01djsIQ1TLUhj/GTmvoYL5KsS2LSxuYVpHH9nVspCDFSJyQ0YX29v/9IMemnYRCU
GNazJDAe4++xRUdLI+2Vk+0p2hXjqTkeDIIHvOHGCAt4FMyZv/605TFkc7BpVz9+sLMmIIcN1eVh
g4LrGy8/n+8uavCHDxODhy3yzKIgqq6NfI2WUQ2Tbmt7goadAxZZEPD8lJ4VmYSVqIdPiMrShkpb
euhwfdyaCGcrXUuEyg9ZasfMyh5i7Ns7C9Z1HcHv97AkahMVqkOtdUFisDdlQU9JYp/WkQ8B4och
pJFO4WFxPTOXlbQ7lIdYJ58Zx7OtI4yqEyKVyzdNsTAhpHJSr9XSjiCQLKe+VQ/v4D/FXdRuczkG
zZ9oUjfQfk5ktyAs4mR8nXyxsitG7OEayZlPxRJQoXdTVFVhAkuHyCbL8UQOIxydNf7MOI5YG23j
L/B1eQwefoQkhwynywMM9tqJ7tRaeirB01nvjk/s7h3Cyl7qPpIvWgePkz+pNVOqokE5s/xZ+P77
rxQ6Z0MWlA6JRPLSB/T545MYYK1XTA67tCZEj30Tm0kjEe7dZHyzOqZfySouJz1x4FWBcIYFf9vj
CIkwMO/tZaO07o48GkOQilh3vJ1Ip/pabTytB144bIGntMnqhQhB3+ICE+Vb02LCpEcAXbZj9laa
l7XkrpU9rNlIYwoU70vtU5xpmF/odspa2RsllkNrNzLcvhHjGy5NynEfDNZTNxEUIRQmJs5bkZOB
r54lGlQjMpzYS/HEvC1XWh6UUR7+Jr9gyxOuGFaN9NkCl6qYS+UBsfvLUGrpFdtTgW4jkADr18+0
TqjZ+eYFAcTUn4inJLHtmSHlC62EZ6700dpTlEBWAKwXRqmXKRe9N0oe6ZdGhS2f9m1+5vx7rPOJ
yxFkFAjOJ9kJKh/NGk7ppEtw7Y+pMyo7u15Min2E2roDwh8VHNMZ6Uo4r7xrMWOj1Omm7hcRHyEK
Js9F5mtlaldVCaJVgkJlYg1znBK8P4EiLM9Zxxhdae5EVa09pCvlYFo04RW9Z+j/IBggIBvWsERB
3afxKx9Px8F0TJMLBAZvBNiYmg/nKv9wxIj9eAEtDukDKGeeuxCxMLH/UFPbwqHPGtiLNkcl4FX4
99GK3Ft6NtLGmzr/SslXZ1dFbs4w/YpOk9xJRhknBLGCmYmUE4h5vWoi7fsOeYUETqbp3LK5C5Iz
35Sdho/XYhuIBoMmRM0Vhair/O5Cs5iBlOnbYSK1LRY+C4MZNUuEjS0Lybf68csskylDyYaYYCwP
yFnx0PQj0MYuNq4W4orvrFyAO2f6tBiI+tYrafCqE6IaDSTJ7o2Z1cL2CR9i77lSB49q066gPuOh
xbpMfFRlzdYJkCctRPW4CJrPDwdyM73HrApotNFh9H7HG187ZpPvWq/4u4jd9JFsQEN1Wv/LrfnO
39J7qB+06fpFoZYktuqL5ErWJk9EHU0qSsIVSkePwOSJ7sNx14BgftVAW/bbkuQXXxnezL3J7vfg
yjqRV3R4rsmE9aBiIgm8MHwCkh7jZwqcs27l47OZsnFuxh1c7KU3tA+V9xe9sK8RbPn8aE8hcGtk
3t8bCMSKS7pFnTWYVEj5jHVx44WJQrfy6Tyj4xIe5ZrI1MBrKt4zZcp5PjNqwGVgN4hDai9nu8tC
mjwbcyMRCZv8UUUzaS1Pa36fpU7K/A+YXbculsx74/5dA505esUbeS69WV5aUoQWuGY/KVf4iZf5
L0S+IpVmYYcYR7wJ48/RWhODaut29l/piXmxDFGNpuT+4IPwT5aJn/HbQxeWOnqi4Z88qofrodCx
Jo4ope/LEj/y5jFDvB/UxCjyIxnL0RgVk/jKURJppzHCPASk+kh+IYuGJBXR97jFxNbaqEMSqWHK
W0UnXAkTKDZxZoK92B8BWmPFNZfWwSZ9OLNxsUB55xX8OiA94YX8oZV4OgId2BX5+VRhz7XHCWJX
Vz9eko2NonHxXWULO/Yi3LRyEufi64BBVk6NsNFKzRwSW1IX/i98ihllKSvwzrC78Vvg7JuwJ5wu
eV8re6g25SwivhUK9SZ4B4cmrTNMz2uDc3qjlwDAv2ZjzhZjnUSdUmHCzNfXqG72r4LFGgkUgRo8
FUc4eB2OXcbLApcdvXqnc2Ok7hanZo8i9ynbibb/zYUUmg17xFpw7q8YQrX5ocRVzTjkP8UMl2gr
nxXty/XFyylJCT6xtNxYCMH55bDk2h7heS0ej0D1wqKK2VgbiX7COYe0iM+8PtRmAUsR7I59BIYD
ajngvOkv/SbkthHXQK6qV4F0/TPriPOO0tFJdEekPsF7mmt0aumfzzJPUiA2tzjRdrwIL7uqIZbP
CnWSSd43UFrWq7ltTcfYa5P7wBMGf/A2vBT3RMjLwKS2Eh7FtBWYtKcPgQMOQmDuuyGde9f0BWxC
hyIZCOTY8ny+fnT2Li1yfVjB889XDhfsGHz0NPE/w0YBPxAFxH0V6Od4Td5Znabuneb0syC957GF
Q4cZriQKOFYdINZ768YETkZMzx63P5ZXPGI7RQIcGU55YR01tPmJfsuJXbI6d4RA++5wpRE5FwPd
AC9t+KZeL3OpK4nPYvVPMVrXK1NhoCLj0e6eeOalzSjKbWYTJw1KNkl5y90PL9wp94LZKgd0Pnya
r1OVbY2zbErjQWJkxYLlbzCqrKLhNa1K/Py0kWmLOxKmajg/g3LFAk3i3y9ZIJcz9Tah75FQmV3t
SgKN6HPzTb28mCzhV4C94xrrzreY+sTbUvCCaZRe87uuOa9T/6mnNVJ5wm0vsfDwgn8FUQYp6Ry+
xsyqcE9QC/sJSgVGZxcpDV58+6pnfd7p4Q68SUSQSBeSGE1dC0pRkN+5hCjNmmxYXyNUMx8FEjbO
rEwDXT0Wf7YNo5pqkCOnlj0a+dd/2J/y84Jvxln5UHNaQxWHIWmgXr9AS/k+6b2irVNr9B1UR1GA
1N/5uoQEApN8sujkS3zA+jz1talAsmmEBU17nQnenoSvoUjnhkKwQby7IzMZZYWii2Cisn1opr5y
nOO+CzmhCcy5kc78o01sgYNHPZbgRCd1YJIZWc/lcdZJ2l5X+fPunH/xCrMSWTfFJMFgbtHBAViz
7EwQmGibt6jGUUf7qNJjqjFtfIZkcShQbWDrV+MBtT+Es0RW1PpBBCw7TL5FmPTw8I6YjVJbI2vm
YFwEEylEeHdBsFqB5DmgPMEUYtDGWFBWeAmw0wtLFG3tBbiYVMaHvryBQx7pTaJYen+FRhSgnR8p
gmxSNgcwv4ZHwwUBLtk1ZeeLl5KCt1mEE5ZKbJexHakV6QB5jSpAPRm8vEDb+G35CigSX7PeGiYW
s6QYoF2FnLDji6DZSgPiCRNqClfLCv9MTebDsvVYU2500HzTKoqFRZ6r7qFEF7TvGoeJgJ2G2tK1
LxOEtXRSTf+V49V6MdCut96DIAzqws0agG3tctxE1u/pifdDVzwMcmpHBOQt5rmQTg4UaPRtIPkw
ts40z/oQ45XxZYqdm1jO+IdoPAQu+lqKW23rlGkwbzaCeMfFEzzGHswXUzKLhhp6tbYi1WALSNDV
6/Po/l74wzniTBiYIY5g5Wob/X/dmE+He5da1WEF2ly3XUSPT/VMwG9vDaY9D1HYeGfP+yFBR4JT
ERbXmY8s6+hVj86ljklUl+C7yIlZpf7aP+JNK4W76UBEKucDD4auLI8vBFLt8in81QGYzm/M40pt
E74VPLPdBR9rQ30U2+Qc6S0iwnNHvKXz1IkUUOVsOGBegDJHV1zwr9qw3LDgq7ZYAem2nOVHAQyj
Qoy5A6J6gb30TG5hVg00YG5frl0L0TWiRzREHnfozIy6Gsm1BOLJIOlr2qm+KbuVjcJ/6+1PU/eW
qaqYu6FxKXoBwZXhbkDujuo8WWdXkd95zUCekVcYDeaSgglGrYx44iG2JYliGnoPy0FXU4dolND4
cwS7eSUcSYn5AMhRD4VeO1m8fdZyIQfkbmKiHlAJk1yb8NPnQJE3+Y6431M8OQ3ghI4cdu4TejCo
B30ULe5PTeovqsglCwYTI/eB7QEwVyxLNld7Aap7on/FfY1CUudlbgG6jK+f8wOlGPnCnnHKFdAY
gAbQDazHuTvH8jrROCyPayOmcOJnHIqhxPMyoCWbDi93doo+xaTo1L+ok5NMCwHbGbrWsVXLdUSZ
3D2e+ICdHoPZHt93jLP0Cm5X1I6Cbd0dqJ2pfFgABrS2uDZcRrqzU/nR2ASjanakHuh9b/j05NPc
GQcguhVvrpjDXsdp5s39jTzXXShDdC1G6Yh7A0y97lKQTZmN0EAH5WbfZdRhqkW6T82COqx9pxqC
o0p1+V+2N3/LfFDsY2Y/1sglt8GUIpuzdNNPjeWwWPV08ACD1X/RIrHVGCQksf52XC1u6tWOmTci
SzBt4z54n4jwiZU0EED6RCzcCBgD73uYeNka/g8R+lrZ7stpeIE+ZHxaKN/eHWXNwIINQmYAPo/k
rEoQ+EfkYgCxQ1Hb4jMpoJuQdDb+R1aYriO3Wxc+yqxGI7Up7jxIQth7JE+050jtQCQyqqoRK6Eu
DMeL8DiGTIccXaokQS+ANtEtVV0ymYQVfpXKH6R1FcT1eeQCWDiqgan97robMYJHhYQBWYR1kaPt
gNg8BYqfn0SMZ+/bRO2KWWTB9wA01g1cGtKWTAAYIhKS8eYm0Nj4NJTMsOtby976Q5f8w5h9Ge/p
BtajAnvF1qpkUEuZR7QuV/BuR0xJI0M5cIE0QndyVUFgARoiNEOk89Bc1V1sdQo7lcOwNNxqJ/zU
Sp+edtKm5DTX5g1SEu58DL+2yFMWY20FUoimY30M5vy89MrFjJiV9RHXY0McXvjTvfTW1iF2I3Ad
QxFLVbJU43z+0RR4sFinckwhxKShOVhQJrZXs6Dk19iZE0azRqIt8OdGhfNkQyp7gbu8lbi0Xjdf
ND1aTLDHIt/eI+xvI6LN9QA1wyYmWd3rRimjOKJQRHA38xblS93t3Zw33zh29gbggTFO6ddD/410
isvWawCrrNNt+hah7XX/1ngywKBPKjfixOSpAJjHPqIGwcxdJAeGmBwgXWXj0rx6gcSzcuGP1gaZ
2kXLOV/Vg+uHGU7iPPi8E66tY0OKveDz55ieShpxB8mvUiyP5JDF1OD7nLKp+BR4SrFxbz+gRXYV
xFEMR2LaxixoeyC5+gfY8FyVYKMlgnHqWxKPwZJPolX+ieqTiQ0GPYju+c2x4Vbl9hBJehMAYHFY
V2mhX0K9sz8Z962+H5pgKSRLt2r/O1EyIPJb9mXtN0Bq2ds5MnlDQeMttnE5hjlvqm46Qyv/iaop
gmSPC35qk7H9ZYNNC1Qhfsnd76a95lVnElP+VYEPOxOU5oTyANTW2MqH7Uh4H5gJzjHdwOqSL487
WmAsw6z27wvRvtcNS21lEemehGgG/UTv7q1RZBoWVC2atNDMh0+/+WDkUIPTYr0x6SPi6KMQvp3Q
OVAulwkDTgJ2kJnnHhMStVusPLcpBlW/GcX7IOjJM7QamMF0s3EjznLAUyRtAxfYXOy/YdDM5o0w
AZx/R1LLehmgyqOpaOsdO11oCMukdMMEjZvClMYubq3YoOYWpxXGmxop8ShSmpy+D5d4cB/BCLE4
bsO6eVa1Wy3KRvHskj1vL/h4PR1Pb3ig5zZ/cbDCID6YY7ztX4++qtaIL/kYbbH5UrCOKrglbVVk
GgH5DHRxqYLvroCbcDQF+d4x+O4ZmG2Rxss5+wC9cOEkHR5/XPyIC3r1CcYnhntR2Pii9Ron+XBx
jB3etJmQ+B4F4bzW63LfjbLwHqMa6WX2mrKUcpUau5OXvaNQKhwp5N59MAe0XmnrxOT9nq9qlzbB
UrMhtTFD2vFuYFY3vi2V+PuAG2an61qvMdTjZ+jnPlK4nGP4gB4Xm3ZF1z2tnblqPVkame5HCxLs
vmMdVJr9THUNWP0clkkX+3hQ0cYxO/o/SQM2Ejg2adrbGcPlqQQcc96L56gescD9+MZVFv9KnxEP
yhY5vJ1jCfApgzhrAxuZtTn4uxDfecDB4/UOsrsDMgy5dVL49R0l3gduuLr5His/21UhpbhzqcJ/
YmXZmrYcKFMigb2gif88P2m8tadfzekFm55eP4TZ3p4CBe9Zoj6BmJFTpSNyLXWhk1TBRdbDMhw9
GROoIqN2EzP5LoU10+Ubhdx4YYHoaIdU1EnkIfehESQophW4QwcpIEQKYGTR6rilfCTKbfY3ySQo
5er5QqAD2bPTagEudfFjbWKXOETracZ9D3a/4qLIl6tbhTaJ5Cj/aB+459/8C6kS7D6ey28Se5QX
d6kBFX6Obk5xt1Mvx0PZFwPS+Cf66e1J3eTxcxBexBv1GnO8T4+c0KTfl0M2KbKZmloHQ3crP6II
Lb38YfqdFQBllrsFP/AxBPwH7pBB4dyFeVFntjpdNEsXLJ3hqh2w9mrhPwJhCp8bQeoxeF2QkSCF
pDE23kld4qtphI+BRG3msrlyw54PYaLPSWrGCGtM+25KB8YvZ2JNAZZYtRhnC/ihHBLlJG9757Un
l8G58cLOBbhiiGegbBri+TWjhNzESFwOTEQwy15JbpZLxn/S/AHBiskQO23J0DEHohsw4TvHDQ0b
ESXBAOirSdwrNPhlWTCKqbMuDeCIw5qMFkZqkflIho2xoMdcheULDTOvR9w0DG1GUMeOMuzHmt6j
aaCjPo1AG7ywnkun5OpyifwoCuEh7IvYyRlomIY52mfzKEdh6/VdCBP7mOJZR1STzTro53EcmpLi
/XpEs16dJz0jUPGuDgqlV+GZjJN0CXGwKbhwbIa5dOdP4wmyBtzj1wfSb3T6M4NM5tAOK+Cwb9vy
IsHElkCqJ84rLA6iWNsBdaoKZUcb/sfG06+ob8n4ZwYHWR3glf8dN2Z2FCDpNQ8IqTzGxD6npHpo
V6JGwWv6J6j2tw/SFhAzLd1f7n0FrXJ3CnkdfAKLe8C8paINgp6e8Uj0U3PVjGci5xrrC4nbqk6i
q3fG0pqMhuSyJrHpNr/uAOjX8q10vltF2wEj7bt8kz/2DPzkkrXaxm3Fdgn9BK7lgkTRsjtmnDV3
U/ysZgRoAaTjssSvScwNhqEmFqtAV91hl+Mhl5Cfv3ONsCmPBwMXoUSqPrBmpVpJlFX0bQ7G6cmA
Vudk32U1S5oMKNL7pA0xukQygdrC7WQnG0RL9JOFC9lPbv3skOnYgPArgBsA+YXA+4oT6AqVzpZm
Lp3GAX4bJ5u3q8DO98T8xkflt/CVcNBzKi7+v6Km4CLDeoHyHtJkJ/mmjO7CTRFYgDPGZ+xCFPV5
2/iigco46CssCFGk/X9BIn0pc8xhKhnZ8vzgDIqnsQya1aAc7uXqxWlrEwWI//ON4FMSMJgClhBY
o8En+IiLgHh/orAjfmlCzhBwWXV0qAf5KqmZvhW3HgMcJUbv00nKyin7+yqJaEBN60R0y/M0g4Zl
Q3zL7hO2R1/NeVUI3sMxEO1qimu1xR71ctgCpi/uhM+YBfJD5Q66S235nZ8PXrCYXbzBS9UyOkWH
caw4iGpYRPGgG7cj6fySnY5LRlUjnLrh8JH9rumF6cBot0UqzCd0HALRCTE9qbvPGIv+fQNw4TNV
RrtfPyi3FP31T8SgEIn1v0N+/KtXnhQUE1+C44vf5pKIVYcnQCYHaEkN2uCNeIRFuzqQ1vArP1Pr
pU1RtbeWAy8oi4R+SzQKg1Kd5pCNkjHxLqqc0hu3VjOja+Q0dOuVO6xkdla8/X3VaHh7Ghlz9LmL
SqYb2vvBBmkD7RKcW7X3p8brekdrnO2izmxClp859tDDFfdIXgEZxsxgOVDACg679QXdBtvmr4vZ
TlBmvjhAUMEKD0ZQKS1I0peT/zigfPDdcFl177K6wVKnO7re8VqU6aCP0GM06ee8iAbd/524RNHG
EORMElwCYhD/gVCwVSWaXA9Qx1cJ3miHRxD0vk0kSxa8YwBdmEhFJP8ZfyyBWOgd2WMlJMfDLx76
jg83HB0uKZ+7DzXSK9em6vaIdl4UFwlOeov6xPDw1CQNLI7QPlHm7JivkEnU5ui6RV6Vf1V05UeO
yJGlFulUc2ZNk0orCJyRAZab7CVxJXS/RpcWhe5K20J0ta9t6j8o8puBYwCyIxbXz0YSOVXQY0Ul
tQB2V8zmhFLG6GIx0npv7z1QjaEOXLHkjFdVi6USQqiCtc+5XNdnylr9dzoakMR2NgWLHR2rfByc
Ftjz16r44YrPK4ArVrkVFsEInekZcDHQRpzS7QF5BP5qDEDZVWR4AWvHEeXdx0SzOegHr1o6+h1d
GymeJRmulID5hVxooD5v3us7qgmWgOMtxiEcpCIGGA/jrKivPggjOKRu4s+qRUhXc6SowvhjZRqq
DLYeKuF6jVTzAbdcnT2umxeVog5qSmFpREuZNoi4LOp37nn2JWjh7cWt/KPXIg4jozKTrCFonHG2
6ktoef5RbVAFgr2NYf2g3ecpTT5yzTz55E5Zj9+kviPIUi7tHL9Sa6Ktz96l+V/C0e/Uv5clVSzG
WT8VK/YB657aLfRLrtynx6sakKaKh2coe8qfoEDG/YQJ3I9ruLD/t3RmDkGUTkJMYvUgXLEdWx+b
KtSlImJHPCghZI0wGB8qUlptX4u9JOIix7J/vtNDXOLnwZY94Onagt3ONwpMuPc0BKi4PuaPJiFR
zX6lBpq/VAHuSvrG+5hapNGjeWiGhNVtL+6h9bxBm/aK/O9A0emUv5vCofFcnpt8qNI0A56e+NTc
rfQzk9xHNiWD3mOJ7ojbawao7eFAMWhsHpz3BIMZX62v6Rw7mL2HZ24GC1gu6t4qCXg34gydmkCR
ymcA84DkgC5m7CDTH4zKh/gCNh+wiTA0cX7im58IqE7IECgfRipBbI7kfTLnjpxeFYdm8qOD0kHj
eqyJgVWjZ2TKFqfaMo4W7hWGlVVWLdQsxxjT8xpcXeJ1hSQ9oFVhO6eWp3t7MOgqniFtIaisTl8x
Q4A+vyXx45i80sFGO/Y9R/DMlA0KanQ6vCanfXvaW0nCgufa8tL07m/aysUWZNlQvlgGGdM2DYss
QItqo18vYilSv9A7jl28iaSHGR4EfNlwyRaMlHIFlM/u/NYbC0wQifHO9tiIT6qJoMkEqtZI8wOD
H+d5FzpaDEvU+CHYPGXgCW6z82/iBNKL6ddYAprR48zKHvL+c1+00l+544TvtjsjKSacdIVVovlx
WTFiLV5KMqjPsRCc7kn4V4iypQsTO3BYPSs2lV6JbVZutd+nrr7ohFkFWschlU8PYMAKWJUfzoAz
vTeTopcl8neJcl2jrfrvSUqqUxq6jTflIw4WaqrwuhJ0CkFU5JwlaTnDBkVGuKcP1Yh2WnZ7rGuK
Va/GU+pujOWmCP+nQGnWBveGYQK56VBXDTrLwkCNkZ7gj2YQGxUK4jxq2dv5/r2Oj6ArTrKPrYDv
GPP+WMpaMz9NAEm0ErbOi0/u/fEUD+7qVkvmi64Ev/yjSTOLfbLMQMruu9jXXD5OVRsmLGycoQik
+LSL1kYx6orLStqbvGTGlYgCJOnZF22SP4tCPbpZrDdDZaiXPAhC4Ql4dZmQ+lIlibmgvoiVZfZG
QIljQyvmeG1jo56cQ6aDBAw91D+28smNCSwAgRMOT4iFtCJOTkbtThFeIjkwSUuHGnQR3Jp/+Woo
JYoIOL7PbWysBW5ST+AJub2A3nRNDMfcwF0GNvalU617rUf9t9ok7TJegBQOjmB+FvKHLXs9qHoQ
dQCgrEDUqomsjS2szwN3q5B1yNq9l95UaNIhwkvQEVqj0WzeFxNHdnlQCuwGxX1sX2rPwFNoFM0b
6FOjDsiKgVQxMbWLYTHhJxn318Dn52yso3orh3OKU/d6AdMDIOK4mG9l6bui+oAjSdrn1Vcu4Zne
zZl2oaoa4r/1GkPbxzg1NYV+g4jlCBM5Ih51n3Gair7q7xigd1Gm4h0wgFey5MiyGdHOQD8nPZQg
gr8u9UppXfR8CmPCkXJewk3p/yvSur8FkPT0676E0PwOKS+3A3GJE9uLt+t8JWb+3ebhzUrPiexK
Eax+pHcmpYrIJQiTd/IHf6hb2MHPgbzX74+713loqzP2dlWB6XytT0KYUflyvKnSy/DZ2EZ8tL58
6hNCcPfT3gIXEiukshiR8Tv8rDaq1MNP7jJaBO5hdfz3+Ty37PRNS7Go9XSbMWEUWFSSND+p3mm/
uAB2k7x7xvqKAXpQTE7lFhZLJZl5NaGSt+Kg8EPqcqMz0icDZF32UBuJcORr/rvsuTtcfayAgzN5
rIwvwFORdBjh4FFXbc+IZ9Rn3x6lmrWQDmUxr9Q7luJw7YUsrbdDLSEGn9oDZMRM9fr1uG7QS35b
+IcLFdJPEWE87egpH1MO1AbqBgNTxiYaHmsoAMpQDUEZPTiwZVEzJb2ev/2fVmPrVz2JFbF1Jj21
En8SsnRZvmuE+ALwDngr8BjUEKo0pTAYOL1l0Ur7vf8yWElhs0TQYciGUqzIJkomN2SdLpIQBjKo
KuXwA/CxBkXJJwMpN9x/6/xKpfh8mkuKirqZYyYo+VQs5W9EUESy4vrgdXQQOcgkFvHmVRw4PVHO
nfqkb8jHxBqgZcp/rmb6IUwnHEvYzMeG7Fz6onx51uK8psEmcYxsJKS7MJuDuXJTIAdctRbXd7tN
xPEFI+wfDJGeycBV5FHVP2pHYoocn6jlnysIpgpa1KA+isVLskcxWuyRDtl3eS3ORAa7YmKbACwN
JNstwxB6/7CK0vsbaMC/03+FGFgWQKa/waWt6ialArYYyrE6Yekt14zkt0wDmweOG9zkvC+EpUrI
XfI+WeJG2wUgQ/R1vGnJTlQZzrVv+n3LfCtYCBJBmZPSD6yrgvKUgPZlrokOgWv/c96saGAyYJbt
lzs7JL4STHgvQIUbCV44D861jMy0PNGOmmc9CefxiuiME+Y7IPiaFhvEjUs8QJMep1o6ES1aOPEN
27BaumIkk7fKa+k02afUuOZUdCAPL5oKGBYip0o5Ao87CT0J+2Qpd8JG+TUVUEZzALPCHGzN/K7V
p+5TW7zt6Wr7B/7AuRlvVLK2scrNolSh3clxAqVi9ZY4GzweU5kDaAe4hTzoO620dntvD0fiJp6Q
pqNUjD53OEZTRIr8xB0bpSXXtSARa35pDvR/ss1/nDRmjY86na6bwArSIwZ9e28smdrWybanDrMw
bpc3O64fOu2FRluYxxiwszaQQQBE47FR9v6pLKAupnP7LG/XDGeanPiCMqGxJo/FVIAX5+K7BIzw
Iss2qzJrDJqfdhBiNxPi+YmAL01uqFRLUapKUZSWg5uIME7R/z7aGUAr/BDiNBAb+1ZODR4prjeh
5hoN47pLXPpoJG7oVTKynefQVKojxRt6PbckMikpqV1Er+j52BBi2/xoEXF9ebxppfaHk5xKICtz
Vn6USHU6iK6wPs3HWRfG/ncKjDOoTyRLxfSh0S8nikuh+mdWCKWKLXzxLpVgRhFp4JtD8xkvyGkm
gSfct6BTuMjs4qxb+cS0ejYfsi0KxeKYOwEOPBX72ESMIvyLclg3iwp+D3VlVhg3vBpkm4PhbkcE
0JuLXp/UIe79hXcqR2Lv7yWJqRm0jpmjOQ/H1viEfo/TRjnl3d7nWLmdx9iLFjbaG0py5dQHYui4
IjaK1cfY3YCjFxXDT9RuqW5kLPH7QEmQgvm1iqu56f94ga9cpy02T/VRQ5KdlsuZmCI79onr3FIC
SZgVxJYKk/bU+VcnNbtlLQLhHiDFyM9W0lmWBFrjnV4KTMIT0VmNvOsyICp7eLyoIl0sgHY3HFrO
Nm8Op2XXM6GwYkbrEA1JqkANV2IVvpDa4r8LqNH4pciuMkg57+yByH/4UNC4soskJ7glHRcz2pe4
+uCrUJD3HZ1f8mPcw6QsD3DbpO7xo/MjrWSfy1bB/mTBMB9tFa9bvcM5hGrZTEcpWf1c4d8u0nMi
e/w5cW74XvBl3kSPSwp8S1agraf3ngIY/Lev9nZ0ECGyua0V++U6DaxTLw7Zytvfss078eXFOHus
RVYJKR98OoI3Bh8G5F9pLIVID4u7fjt4Z0Uk+sBCkIbZ+edMJlqcw+/6owkWrN61HPYLu+qcffbh
4+ajP6LCmo7ip//Hib4MqgrdyUNQtdC2wkwRAVDva9HMTHXSIDpDeL3Z4AVIOvxZQqAdYwPAd8AM
ISVZgQLk7Dl9FrZGd9tQSB7trooBl03cSVuMzRPL44U+kpTsM5vgAKfP5ZZ1qd45iwzAfYa1vq2o
IxhBVs+OszNJLofv5qLdDVswv13a1Qrq+0HiA0polmiOubQLPVlJYnS1wHUkEHXdOhgZ3UvRj5gn
njdnzwmbSf6rrTfU68rsD1WDO7MYuJjqOBTX/rc3D3RWfdb9Qe7WuvzHjjiMJmOhvAnvOXtBRJx7
/+qo5MLTxJ8i7y8tQ1IMbAxDQNq/R9tIxUpekJR924hSeF/use08tvqYFhdmSjJIdGSS6JOTbxgd
3whKXv4iJSteBVtxCVlYNVZvD2BPbVdld4QfCVNM6K/WQ6SiBzompN5zJ+GrlGdnpjY0eJHWDFQ3
ASdlAIXKgNQbvjw0qYZjOkar/go37D3aSN7QPOwCk/xC74JTaBHXtyp0A7udpBkqKnrbfz41TTdn
SOCMGMaOx9XMGJW6d2xAl+EXM5DQJOkMDfiHPSB+8pbiCZBgDdm6ESkRpfgTW4fRUrJRxYfzM8Ww
RV1hO6M/8MxH/x5gkozxmWGshgc/xhkxZB3FStbF8Rvt4/BEjvugtUQp7pYPBIP3jGTWHp4LpLNl
Z65wnjs0WAX+YMQzofcBcwwu2088dyjlUX9YdMSHw6WjF99y+nDEl1LAT1az/2aIE8PoLsVikZfK
RYgZNj+7NBsdUknIrOHJvdTVFJ5tJbSHIUTlVleYt57Ebht3AhtlRMnGywpOmpLMofv2RAnNrwOK
FwV66fRraEGRlWeV/V5CxieDTQr8FPJ7o07PwFXmXJJQuXj0ezjgEgIt8rtxWtuBw43UL0WfYhkJ
Hiau8lFgApKsfJ+yuS1FshWbbuNgqynS3AazszI9uGrNzoq36PCMzMHwwoLBSOEsoJbrPP/pB1PX
6L6o2giXr1Njk4GHaarlsbKIqdlaFGTcGmocghDOXBVaNXB99x3owWwQxRvyWDwMMAQTESFkLKHj
N8b3JzcrQLAkgJZcHW0YfIZvrczWP7lT2wsUhffeA1JhBF5A0bm83dTsvEsGAD8KyG0WIa7DFGrE
I5oaxUWuojqmh9KZVuyovmxxf6Ibn4YMuU7FYIzEuNL841MrdZIwKUVLtFJ42vcJePiJE17Iuk2H
qkPQR+LnK4Mri/zjlnxcHkJLSSXAyxvGrndgYCcMMgnazfKHVg999MyXT/oRHCVbOSRNE3NbdgSI
OaAgBNeEwk7ju4S+dWe7y6Ab2/M1T/agqxSXLDFJBNCbMLA8vPabfq1Y3fl/+HPv3jqReuVzP8JL
GzjPVPWJNqXshCms9Y5mMUlI5aN4lcgTkAF6vs09yYr04mC5Z9PPej+7FUYSo17A0LKup/kubAcb
MGhaxtUa7mmKpA8oPO7McP9uMydrDdQchC0iYSMrs+647TgpBq7cnwsdkZCBRfBSKiSUXUkXfYbR
Q12Uh6uib8eb18Bz3aj7r9GfLu+kmqW40FP7+56phpENsYO30otKxHgBmzTxwhP+mcW3iiKdVqLC
RnIe7hdwrBNTzQGMfqT02BfV6CtTNopyDzh+CS+kkc1z9atSa1jUEmSXDzyoecT/i3DWIbWNU1t2
Mxb+p19Bf/rjSuQh7WflF2bc+eh5w5eTbZLHQyLfQ19OSnjBP24Smlb2z8HYzAYFPggMz9hkHX3U
qloLlUR9vI3BbjNnEmf+CRpJrkXj+KaRCKGGyT6B2RAjOI37xNivUO/ml7VQKW8DL+mvqHwqvfgU
tW6ih/CitxDl/l53AV8Q2y09IvEJ/HiYn9nrCOAstLhcDiSJtBfKdA8qPXXpDxVlfqBZvuBCt8XC
nnaGhJOXFrrFHjX0iXDINpfQCyZXX+X3oE8qtUzJd21qP+BrYCV3Rt5rOttEgJJy+HOJkYz6kji4
kiWJYzGgdG1g8vyEPquqLoyVNvxBqbqonlSj1ybSP117y+x4MoFEEwoopcwpC3+nFNwT/yMX4zWu
SNieqQ7cV+xl86jDCvlxlJ51lBFL4TaZh60Rwuu62Dp6QBxNHKkHC2VIO37HzxYmmswjE1eEqhtp
QiFYpUUuZRD05PaGfuJBul9arxKTbW3oYRXkf7rceCp7Yf1DFVU8d7H9oZyYnvYA2j62Qgp8Er63
enxWwNXYna8BajdAW6Zt/6h8bGxFfRz7Ls7wjuw++UURtGAolAATfKXuepKpJ4KpTyWAqBMJaZlx
BrYfkkkN5zVUso7hlnCL7c1J+FjgOS6KSeBRtYjIwffOecKaPsL+qZ0O2HjNpaSgRbvRxwvSr6cn
91xucpbUd3sNtN370V6aLx56tg1fMGBhOnwT0SJ3H5tjKynExAs22ceHc7BR6UV5fBzC2JF2y7hs
1Gj1+QpPkR9ty8A3k5Yt28772mYwF+w5rx0t7woi7H6SvBQKjLP/NgIAyEIH6ON6kGzLLXZQgce5
g1pFHoR21uex7VJqCv7ywm+TX4NR3aCbYZkgpcky8BRpPK6F/EH8TTl+Fc9MiU+Gh6KtdfU7DaxF
+g3m5N1tjnZwRAquvY5K1XsI65Tce3QPji9D28lNfEaKHlHnhWLyX41HrVB06q2FPsM3S2JNEkD9
aoO8tTzTD81TxxM3pxCg3QRRlgaAPIjO7M9mMT5NLeE0Wn+RsrzXH9MgQz8Y6Ef8O+XCLvkS69m6
ESe7fWPcBVV87zjuCv3pg+XtEHsvtF9jCXMmvVT+N++SmiGQOMPQmvnXKzjUCkteN0Eu0Sagnm0o
CFwx+QjopVK13xQaCMXUIQhvB9P+Dx/smzHtveeV4KsuhULs0JOVA/YSv2vfAKcqj2tgZG6y4GBH
OihF2dkZyl5hnANcN0V3lg44FB98y/ioXKbaC/rPZEdR+CFoZx3mCrxpHFpOdrzJeEH18FpBNXAY
xnrZsfI4Pl+LKhpJiUkSiflJgDBcW5V0gdP727bQfm6UNyeRX/dXsAbDgR/H0Qrk4O1X/X1bfzZK
cZ/6fdiJU05OfANaeuabMrEiVgMAF4d+YfGxwwOguLd0ki1zDXrgywKKL8nNg+45qGpDatBYA6L0
tOaT7a5BZ/UDwFIemdHEYgZ6bfNvuwlecIgjm8D7VJR2Ke1Q068Q/Os6EhDIQDhGy5lRNR77Fl8S
wEOY6OstgwNYNQhycWFZvgdaeiS84JWdY3BtEPsoCGz9XwcBY4qnUARrQJiX07rOuiCg6HCZYHYU
+AiNhXPnL3NJ5pOALHpVeZZYKTqEajHdNFfOukzoe7enCoiH5V4QVTClaHFe306yB3WOrZF1Iopm
nQFcAvX4w/hmIKk7i3USRKkQEe3DQixNcvO9I79eJyKEVp3BXhEinRs3ZF00Ptc4g+OI0jdEu/JK
ev5zxW+bAGQetIy7XdOn4kuAxHjx0T8jBdOwXs+jyjZfZdo4wComxsekUBOZgiltAkR6BT4sjwW4
U2pGWAWq5e9I3YncevnwD4Wwwgg+SStSDuWbRzwKhIByfQ8tWfJqcHDAJOH/ZW6b/577Ax0/lqKb
BHxokysO5dPq5oxp6DbJdaMJQKJJZwr80+r2aOmcfSUI3JU/bcgdsc+eiwMpkGDXodc8gVAFzDWV
e9BGu9JlVmRe3O1cl92DafG5Yqo2Af8VEUHLNpjizRWl6a9WcLsWOpxO54H0Pd17QkSVAPpwNGQP
X8lOnIOllv0f0mR9fRzLb26oMY9xiq3HceFldP4njvAkzoTAjhyx0BTdi4A6bKU8PpcbwaDPflp2
0I+f0jHUdnCUSkvxMEpGOqKf6xWysJXpWX3U7rR3BWT2MjHtUNbw6wFaasKxH/aDryFe2QRb7j/X
F6e32mxaoEJKZg3fKeYk9gPLDhmjHXbIn7u3wKz8Le31SoPE73I51JvwJKLjp9O7zoXakaWIAByx
9VQNJ0stmaBa4TNtmRJjE2O+Kxac3wI4Z5HTh8ekZQrfiKnB3qxfsDh+LHaSjPsEi129eKBU2qYD
EzsJyeRDkSKN/60J7gWio4Q0qmLCB7V8lliy3Fpc7Vti4DnaUJAvSog6LxkGuUC9O5t5ygsEs5I6
EOKkXl8yWIJkfXfj+Cjwz2Xs25pTNQTfIl6aAOxOwwK425MbTjo3JY4LqqnKlD7GsTf/WiU9muSv
ZTSxVfv0LClMQylWoPnqphSg/6eODb0h6OWf5CqtqTKZrCt02SJGekqYy5K81o7LTcaArZPy4n6V
wQPR9sUOd87BvN1L4sHXRMkCU/BjcnghSoI/eoJ20vaQJAZjTTnH4bvsp4griZxwLyzKvi9/2iI9
P5/UnA0luX6gYStPbyIhihqPUmD44rftDS2jYpaDG9yGCp+AmWeVvx9yqaxw8qmOmNUZfHgnfttD
mF2qxe/5sNIfroGQ4veVZjWMehjSNSEGnGi5tNCmxZzspuVQKD8jNuYfU4Mnf8jbDNZ1aM3Qx64u
jnEZYDd9X3k+tvjcTSOtbRpu07Uoh1Gs09DBFW4ed7uXZfmIsRioPLB4g1GM8Ok25CvLzgO5CT6t
gs8tg0wmL3JNBus0nJeZSqnzuchCJHFKfnaWPehsac47ahsnhsiZYNl1/5S+yj+ShCdSLRujjeWj
tx7vcrWXyUGA2jYwZEDtDlLEW67Lf7V/LL1UcAZRbbuhQCqbD8mJbsNUxPropHFnHvcilgKxLNlK
pMsraP9rd6KslZoE++2VxfUbPp0nSS6T0BCJFkoElndkHf6jfGar0knx1p9l8kTh2NlfNOqfmKVf
qCbmaMEBn1/VzXKACpd1AcsZEfVsjZ/C9F/qHpATDnRb9iws0SAgCHmOCeYVaiMaZ+HI7ca2+JCC
ybeiLOG5Bw0/JNO9yMgDS8LqZZ46Tk2+MdKDQsbzi/v/uq3gUDhD/7Ytkza1Abcgg99kkp9Vp6l/
wCqzg/N3VKxSJRv/mNMeeJVdm1Qxmf9oyS0CQOqz03RyP/nnbsXQsSo8zFJy664OwBn9ubx3xtGu
lU7zRCT6yYHm7Y5LewAKN3Eo6tFpilNlRXWyZGupMfXxkpcZy3ffUMnRUVMT7IFxwM26dWAE3Ocg
rzcIsogw0SJVqBvGKZHlKtYDFSc2/XGsIxt48GfCo2pWb4QFiaAhJlncj+OggMQiN9Pt4uVzRA+k
m+iNYQUtc0VRtfZp8yOikXRe6POAaAQBai1h2rNn22aH8eXUbXqMTifSif6A9zg0tUDdrdcUqnK+
PheuFKd2FekSkRQITOJcuWxB0d6Ra+saMtMzW22MxdxghmrWbWNDj+G/OKG9OPabwsr9LQ3YA0dI
54OC1xzNKXkMNitBFMiXlZocnhTnKa9ch5PD+Qf+XtBT4tNOIM62qUNOnKLOyCPje2YaviBtId86
WgtCsAGbKnMra25Yz4KiFhzZ+B0PWs3q/Ix6WMtvQad8DelXH5kkVW1ULSzVgq33qvlLDFO4Wtzx
BLeLOtrGKvRkEl/jsC9U0YG5ShTbUs0874CSnzYNUhytrp2D4icbMef/MAHmz2UziCy53sYL2qNL
iMxxawq7iuxoOuC9ysAegjD4vzdtOmoGxza8ljgBFMM8ivT2tWbubgJHAh+8IhUrWTIxTOjLL89K
XHUzsfqZuRJa5LXXqJxwmS06N0PAhuCJucWLxW3eWKvF2wWGZ3IXPPkgnH6R87kjCBBu4btXPnCv
9gJuscmt9CrRZA8Zn3XqhXPLPEKGca099sFQqhxbVdFff6haAmAdkJYlQmhyQGjl/d8tpoU+dxMD
6HFMTJokmfoYTyWr4fmWh/G/zhoZncjwCr40JS/7KmjnmN6R5V2NH1Eaz/VPltX0mfKXDKEKwfZQ
Pv7TQM1/KPht/tWw79S1sK5EZCyu9Uxjg4hrnc+aS15aJIhA9wyCbxnJARE4zpzvEIFNSXuYzVb7
lTyr3xU3z7B3fGLKi1/6Q/wt7B7ffbSzi3bkFFu2YjcGWQlr4PMSHrW9i1JBthwVHVDRcM7hcKoV
TcjmmV/oulNb0T+5rZ0ciyASrm3qIviDLZgn0PZdKkDfwufGSR/BU1CIQajJwmWWgnTBBBeTn872
hx1e+Ynf5yOMyr4qN0gXIJpb1HRpoDlzc1aKU+pL/tl5dGJozpZPdgNtSbuGvKQ0gHpP+bNt0Woy
DMFaPqCsET0HuCfnkA+3x1MhGQTJGTW1+pKvFylnXS/XdPxk5rP2K8jJoGfPMitoLhr9MvBYoD16
827Ga7fPpfJPLFJgJxQXsbJRY/o+QKa0YPdNxsL5W/1I5q2K9BdjgHIYgJJwZXVhze3n/9/Gd0HO
2YeClWKepUIqxc8HgKJ+pTJkDV3p2Vy++PiolBhs7F0Ag0oWWxK5ZTTiKbxeIpUpJaj9vnpAkHce
k8Qoke+u6WlJHIkPHKJAVEFBsv58kCp48XutD6GpOz/ICMgT+mtkraGiAhupS/wii4ZeC2z+7Bk/
f4ccDh+Rx1i9GUdtpRNIoIuWCV5dGGcR0jIpFS5nHz5rlFyXFQZTb03KxDH+YtGbiZhSj6//fVx9
bk/pE8RUs1rZp5O3LcRWgH3T8rQOtFYD2x6XGAgsPJrPyfy6fNF7LG1/fde2jCXOxWYTMnwZRKSs
CIf53ViV+dY205CLfi2cVMPUsDrtB6P1C5jt/yET05OcHKS6pkMhY+nG93BPdtLS+6EXnK6Pw5mt
WaylZrhZIn2r+JFAwnHl2ttQMwaw1b9xord3XAif63eLhpk07VgC0dQvt1Asg9KjF0CremY5xg79
vGsMC2V5bFQqvg6Zq6X53Jq8Gm+MjS1l/NZqrHYzXN8chK0gETRtPXhaRy4gabLbPyRrlmbX6N6/
zhiK4D6rfcTGkkqd+18DVPvE1Lz3AZ2Bl6S/4POuGYjz9GkW82+Fnmk9Vk63dVBmI3Qh8VAXLy3X
KZz8rzaIizgOZBC2NFUWRhUk3l+WYdztytFWS7RWKtqPMleKrLi9j6M0niYQoeonxppHufy+1sEW
SgbiXrzBcvVHkuBUURqb4sljQUOiltHIk0o4zwz6t5CLIXdZt5Gk6oxizHrKidHjrUAG1s+2Zqy2
D7d+SUcLoAW/LLV1WsFABjUi6htQaIZYHchNZremHWsM+h9YOh1cBpLhZSnmh5ScX/u7HjYPJawi
DnF/Z48faPxg1Qn/fsHlN8P+LCyGp4hr0bYycOzT1j0kKod0Vrv7oNMr+cvWxiVRqvsDlKGYCWa4
pMEx6rs547MMKTsaDsw25OB6Ckx9Z71VUjat3XLlcUjMp/E4krHvhK+cezmASx8FhfcLHh/5psXp
UpFRlcOpGdkX9jkeZLVfJd7bCf8QPPwtr6GR6EsjnwZ8pSnGFAKePjH5b13r+BpxzTH91ksNpITw
hqFZwVhbgRmR1KtBcHD19375A51PEAEKhaB1cxnC2QKyzesxY8KGuvGUUfC8FD8U0tVrxrLW4y1G
EL2q/cRp21Mj8/l9vAmeb6L1ayF5xrl91TeGgp4JR3FIqOlworMb+PtheENof9Nej8zOoKEC8n0S
BWzGxC2BjlxvtuEw575w4p5BxnVynDjhSvJMipBOb7Y++OCTb27lQ20DBIEw1Xa1Sv2W7tfmk6Ci
ViRiKm3QPxQ7POaNS3dUH0Uabs2WMvnXGfK1oLdqDPaTw6uH4+VdasvAN4VXd7zZ6F86XLmlDacD
inU9p7N8D2pz0fnBBc1nZFlPh1P1EKsZ0eC/jy2619PQi6tRxrlcv14CDSNbIMwgvLJSK33KQMG+
F5Fqs2KBgqMe2HpqpRJ7jYg7LeSId12nOyitqTsu1MqoMZ4a9JkZBj6ZQQDT6CTNNz1XfhaUpCZh
GmDnu192uO6FdRr6TW0/KHHySD4C74qGB/DSDplw6x3QpqGPq/mspGyOgJupEkvU6MyEcGX0fELr
LAVJXSfmXeOxzixEDh76ejfvBYGSDB/CJwq+ENOgTswE6EvR4GoH6u3r7Rydc6F+SQxW9STdEE7h
0lSKSoChfit64RQpVFGLQqtROj0UbqMP2yTB3czmGIsryXXtKQEcgSpk5G50r+pGxg9LIBrKWE1/
ZHpyB1qCHHm4SL7rSXzJi8pmWscIknW9uV4X/NPdcATTVeCgEuHjAYwZcUbspRHR+zR5WiIljggY
mgqF0bmr5ocHmD+uxffnbjwkxZ5oJwosAKiw2bb38TBjCu3+i9HVjQAp9ocajJSOvzG62E1V5ct8
i60Ppc6uxc1jxG9SEavp1MQMvLIYsQe2hM6MNkLId08B+7kmyn/axiCBnN4LcR/biGYfG/smTwkg
k4pw0YFS0fnGywcJTLWbX1xkQet/HECpjBzGzcvOe5lfi6U9nqdtPsVVGZfPMbt79o0cjvAMAlUv
IYJmMIKRrFh2HtGsPJLmCTxX5FmE50LBq6U3kkrJ9ZD/Q9oZIEuz3pe5qUpYj+So1agANHYlAapp
W5ESs2h4zA1ZuMWW5ejaKejVyzCH6R3RIPxmMZdMM3TmCn4skMQ2IPflrtBEfHWDLExgB5EKTYPm
A6CRn5uryU54+ICLziWgEYI70zxiuTKE1VqQAS5zd1FQvkDJIwLUq9Ogpp5yuJF0ZGPWCD4joS7c
pzKXBd7kzCcz56Q6H3WR23/BKQ9MbH6yCD/JeM0E/kXu6ftPrAWK939BMrtNz1otmM+wbgGZWEsB
8rePH5J7ZtWFHkZx8uUdyegZBOSklA+QdPgJjQrf7bVkMk19TnrRIgFgCuJQViMJQ9TDY/5yqcEO
qMpCqgH+G4cblSTvD9zTaY/Z+Z42FcvPWGzJ6x0OJhLlr6556Eu/QXhT05Y2eP8FSQlNT4z93N7x
Gzla6Cb8yw3G86O9GAV6hAspN/GMFOSN1aa+PhVawcSEiP9pp/G+nYwaxpjKXOumXnX3GNl4Hb/D
R9eU6GCeBHuqVj+C7m9f2EAy/7wZuJYr2Twb56DSjA1GISB3wbCUgmQZBAjCdepwA5abPldhEoqy
8XB6UNDikiWi17qYSwaqO/7k8SfUy8oiGdayLduUNPszmpjgnofqhAbbgCZhnaeNmad+aqPYjI+V
HAQu1wvHyL7C3f3Kqd5rDaYnZsa+4GbU3KYrCR3rE3ST42kC00GBUAYqwWjFhECyjlam+Y/texG6
bvb87mt+bLaMTJ2Xg60GUQM3NK3u0m8cUfVbcewdxl2JNeocT/78tcfD+4A5jTIAdc0njjbqYqy9
0JD3lMXWn7TV5FAw5seyf7KdL2+v7yg/wwjKXA91GpdWwXAahtUI5nj4gRVHpghlzB3RArNdT0d6
BqL4yA+EWjnijRuo6N2SEtMPD1rQAjbnEBJBBhQpihPoBfcvva6XBJe/N1GGoGxFPDVnuA0s0DJL
MbHMcg6QDWkaxD1yZW8j6kM+3xXwi2ecmtUG/uMoXCiI7ozfGHx1zZhHIu7ztT/q8xzqhHnFTgsV
XaE70wlvwES9enYBJWjg6lOmrzanjOUgSd973EIRhcmH2FANycF3AvY76i3VY4FwJliIDVGIRQcq
x11l01zPtLoJoxHQPNH8PoI6ij24AMt6dw0a3DFRamyhckLI2SockeiQ24zV1VRu0k38OpMwhsdy
fdsUk9NsRB/avzb+hpTFWGWd4jyddZW2obWmNmLpPB3KuLi9Kn7b0tVe7jBXOxFzz7zbnCfD9UZr
iK7A58/4DyCU9JzAcjPlqvtf6DqufjXmKPQhgrO13djtynhIrKCLmHBaAD6sb9Pj90zzA+2hGHyJ
nrSDllCvorxrsE7k+7TSbkM7v2ndIlSq5NXQZTz/7RUPj9IBq387qTsKglEdcRK3dcPug5R43z+7
VomRLlDvgYNj9Sp185lFb7QHgv14mXUZk29E3hyrpsapWblQ9B6Ca3JKFxZP77ZkVlOfVuGwBNZ4
+BOwEJ4p9e3hsPsv3q0WkHAMQx57wENzQ6dHN6d04taJOtaccPw4SXjpwwrh1GyVaxadHQrvlb3u
GzIIcRjPAnkjTkUYySiFhM6n2o2D61P2RJjfTC9lMbBU8Wj9NzQ3JXTAsci+TB6CwSaW9PfkdmR5
mNYBwWPAxLCiazvzyMV4U2FdEinPP0fVw9PHIWeQKOp20bHjxQ3NIBwQzjtJqinLDkDaOZYnL/Yn
Wyp8gyckLvtSXODJitEZVAky8pUEuAkQnb4LBDSXCk4eSZIE+tjFyuFNoahex1uaOlOlVGQeBOQR
uhPVBH/pCZ0QYDZ2/1Xz+vBrqin6IykiItrbU3TPccad2nGMLl+uXC+E3lltWRfJsollQe9Vl9nA
ojvLkRdY5t3lQzA+b3T24/nJQm/VTsc4MVSW9ilOV049Uz0o+BrFHWp9ejkwxd9kIPOsPTq/LFtG
CrcAv/T94xoIpJ4tspwTi5t1rg9gW42UNlT+GoZDY8Xxtpkr8eVdbaLCrJ9OUDi6BEps6BRFl1ZD
be+DoNslszlPgABtR4SxEE6rhwdZ6lOTY9ctl6vnjhaUdklBB087pl9OGvoDdC3Zu2ZNEzn8qtGt
giOsNDLKsYEs38e4ngoE5sblb9IzF2Saf65mtj0oiUVfBetjuoRBJm4Pywn+6HlsqiDJS2im6CYF
vv8+Dqr2aIdw3iNE4wIH1kS1qbXhZJKl4PTZsF1gw5IIvL22SgfQ0ieJjiH88cllP7COMwuC3CQu
mh7yASsnUri0Sio1Mb2VhAYLe8/G/sSYbI7OqQbKith+P4XOicK8OS+GxfOoJn37sDPY50fGvdLv
pa7yLV773PmNjnms76/6OIDbEKX+go8ww3eHKtnKVOLo/2NYy/AIlD3Ou9UjP8uc9/OIq/aM050j
rqZOvtXb51D/VTf0PyHL8KZhLRCddqDYpN8MYVne7k7QJrW6aYxhZXjSDF1P4jrhYUVYvJzc6ijr
ofVN9CY4dC55Kb4QoB4BhWVa//8BLikt8zJGKuAOiW54vvk6EBcUgV1jiRAvxXv2iUz3RojXVrBa
cN9tn6yhvCyliIwFR3P+WiUKe/jUdn/lLGY+JWaqcWCTibIwSgGrSXeIMFJcv+oj2tWHngxRb1tR
xE/o+9vUpeUj+jIivtGZXHVM0bTfVzwxRijbZvgjkReXIE09TAPtEoWPZhp9XkCxCEOS2KsT6LFs
GejhFfjYoqz6kHuvFTKYTWVVdfm+4RwXrBc1YkifiuP7lGLzEMqxNeW8avDmUYwcKLJlX8891bF3
CwjvTzJbcqiNMR3sNp1ByqXvnCueYS9z5pEcrOtbl3BFG5S/E+EPngHDC7VQBoslv9yqB+IoYOzN
hRz/4/Y1ay9yVsfo6i911eZ/73riObxkXYbBTHvMfJ5fX8f/0UeG36oNsPxhXhQ345TbtnH4s1uY
E9ir52ss2YYLR7sIDIEXi4tiTjr8TgfmLUNHpcjNJUYelTUXEWBQSbMfz8L5P1pm9D7Z5TKLzfo0
+yy/Qi5IPRtgqMNpOh0fueg7c8ZdTdGJsSzkttbuqPBFkrTYfyyUQU2btaUcUVOw9xU3YBUCex7g
M48+Lwc/brRotk6IEKhaaaKqU8N/uryoyaXbnWAWCxWImPM0BT6Z48qdLvRmtIcWu5aSVTnqMHJ4
5Q4PykfhZSPEhwT5muWyR2z8cRsWc9qYaSzS8HdnAMgm+YTakvAqZ52yrf7a2D1SYrtZt1ivlUw0
U/0COR+q8iO0VaeEsRRMufFuSZwq4zrJT5bkoi1dgK37+zSPlHQ1vtQ1Zoc4id9m8aNQ1fUMjbeq
6xgBzdubKk3gRYbPJ6xSAXgMu0RebcMx6lw9dlTHP6MHY/D6diRyz2MyFEHr4Eiqdx7JKJs38I0f
IlvUik0PulD4pDQpZaCW1vqwtH5iEjOaF9SFS7hfFW7Zk99TLcL4HKsdSzJig9ihhspCx4C+Cwza
4rtr/M90ayco5/Nw+AOiowzvqwrb7CR1HUVIt8+c3oyzctD5sfNuiKQEIZDpFgO///kTs0MVFIZP
NFqRk69NOXwMYwYTtTZBUcBqU3dhSiJse9z+hs7xC1j7yKG4BR2FfDeCNcTcGhBkhReztwdBzoiY
FA23f+Vmqdx09z+AfRimVqCymnKzF5tIo1JCi4SaffNzGPZlnLiLIQ7CQjfTchtt0ayK9dbibF5F
thKXYUk8VG7PwcNhoI8KsyDQA609nq7XADb/LkdOnmGT55drQP0WBzARw+8u7kFM6wWWvUhQve+L
nZuMoFbwmpVwFBoZABx+3vaQyyxA4G1kwMz1MTgCNJlcdUsDARjJ8fQcOuNbcgSqne57336r2zQ1
USevNZY07LpwdX6/uQyay24DdCY1zr5OvJ5txAL+JM311sI37zdsrbd/tJxm23PRfKzoX4SyrNxn
OWcqhX5qWvSXsaWy9tD96+TcYEkxD2cG4eIQqV9a+XxCOyK2Fx07n6tThSIUSgqF6OY+OwkK3D89
t+ESe2/rFn23+2jANJR2smNZcQ1TQXC4/sTtg/MEFTjldghUbRZWaDSLDHJExyC3NNaFTCOzcsSh
YkjD3J+4kjbZ+EXVn78w5/a6Ies7cUdM0WfDl+1DlaoKIIkkBQwn7X2uygPVsAzTRxbP5kO/je09
BK4gFtU/ObFrZ3CWHD8e1zwA/PXvE3GHey/F1S2A/TjGJ5+7iZaOuZa5PXt/YkdEAdZUG61ykM6i
WovjS/qYVpqVmhm+0QnIRvazkL87TaXhyuSDLbxtUGDJJAxjvB1IDAylamyw4IPjadH8bf8MRBFK
xcmBE26vsRwnitb1BVAX5bZ1CTEujUO4OTFBNlMv46LqjwJlO3KgIz8dDtOh/VgAfDts2ipUWILA
etkqX+qVAYhja5MWlFPhkBrXPOsJlMEHG9lW4NSa7MUkrLrtBS1CH4j1xjb8iHXVg/U11FnglSF6
5Oq13uN1mCHrLs+sjON27MYaud2N9MHwn96syttGHpRUPYQRf7qltAuKOdOC6MFuMQkkcERv+woX
AuVSYIxMYsbps/CuHje0IUrRukoudowuQXpOHIu9i6HVqFnBAesAesujIqjn8fdxVaXmGpq9KHDd
F/F3wD7WcnHDWnFBAV4oKeNeoTuVnI4j054awOkEnnss9yta2j2S/I082Si7jSF8I+Lilv3nuvF+
fUHCiRe6vgtIr7qkj0n5K4x580MSZLp93awz5wubXSnYVcn/JOeoP4UpREZ3dHOZzOquLZifzu68
6R04lBPfFk94R8tz8/d9+ImLO/gPT8b1mazhhI0X3k+dgUq+rDghaDs9JXptwh+R4nC5bGHZvKjU
985onyRFoKCEUcbqQaTxgfX88tJ/137Oudsxgan8/D6rZ4iynE7V2/BosyTvN0+p0mQ6dBJSSHYD
8E3JJp7nDwFKe5taIQ34jNea5DG106o2VrclrYv5lz9VLSkvCw/OeNHkzUhofFnuS4sfzuOIN11q
dEQFG65QyoOD7ZIrqKqBYT8Gcx0HvVwPtw0KLt32zZwtd+1qXKbUvY6gvZWf1nTN4N/rmoYmvFBL
oX7D1E1nNIH2nfOCxI0wG3BxlbDszchP54kLvG3CvgfxqFEltEyxb9n8ZVZPdLutsyEzHmiVDN81
Trdqv/ox/FxiWuMY+nd4mX35J5Ga+9QDDow/4X41JB8c/4jspF0prFG/Dy1zjzbf3KDy/QxAnDkR
NRRq2LIicgoyserL6iB5Nl1DZxO/zUlkLOOqqpX3u4b1MEDLNpK5ssIieBPyA7xxs6keqLajVJuv
HnyUk6pLGylnTx5QmioKYctHG85KxcSFXWaffoUvG9Cxjt7oMzefz1tE+3YIILmaGk0DxNk9Mja7
UKvUs9DsRUqrCIrQcLAkTVCg26J9jBV+dJdm+oe4QazKCyxL81ngW0l+7XyTY1dOBUQWjhb87x2r
d6MHgNyJQBt7lm/qp/J3/J18B/zFWrjlVDqSsgq5toPS930jDbcl39fFSIV2NksmyFdE57szB8oP
rR28SpkjuuasOKZ+p9oKtevCJjp8f6f1ZiJQ65vZBPsxuQ3/5WIBneeP+uoOtaTbIG88IkE1KCJW
cvsjrn5SS+VnbGImbITU4xN2FznSya/1M8IkagWoVwyKaA86eP3hSmUD/8qyJqWopNQMfNZUESYK
hDa8Of/SGw267CT4p+Hce0ggE9qHTkEJr55ZyX9WPnYqqbyx+L74/odFs/x69GOzPZhk5tg5kWti
309NE7/1FkrHPam7u+sTq5+MlIKKmLavZDCQBZKjWXpCvWbVFNikhZlqIXp8P2LLrdkfCcHoyjYv
BvMP+eEyombhWOeYSGi/r1MPbNKkv9dout9eCPh/rn2mgrY1ZDANGSjklSEuEWK7dI4QZAtvGCOW
G/hruEemHVP3Fc4Oc05xxGtttbw/R4X/gB0Vyv/Qcgu6dhH7DIu7flbOORUpVzm8EaRzWt5ed3+h
wkshNQztsB3Wkja9Eb9usRIRCGGasHyRx1bKGuhc990Z00X0fOoljDbwSZ0JNS3VIMK2tQk3eFYE
fltLNVLc5RVmjUpUeiZiLkxyQbKAFCoduK91n+LHHTslU8q8Y0foVLDWkSTtojK9vDmYpYr4bYx5
rK3sNTOjx79wvRzjROrXTx4gOp4dA21b7QwBByqcuO/fhd4Pa4ffwtnQDpBB4A7KciFCbP+YrVh+
1lQscwWuMWnPWrEPgQFphjPVEUn76RTkEkB0U1MSBhXTvantQlh/a16YcbHUM8LWiBFysHx/G5vM
JxEudpG1vMUu2WzFo6QTWnk4EgKByHXJnA5C+U3q1cko70wClSGULtJ71/UkcDkf532R4LRHdcQM
sjcxo6vTH7dYDuwbkTo0NEMrOA9yoW9K6/zgVrDpR3Ik1wswYeHxn6xkCCtrrsc69s5Cgf7sRQeS
WjgViprNj5bwfFr9KmvBFOR0tXDR6Lm0qHI/3ldIHW5G2cvr3cWd8/lek9+6fkUheJLpqTk1rJqR
mAo06644BdKlibT8SLC7KVFmN6T4b4i7C5pWfFOrYRxEBHYCBfmphxv1jhu6kwvbrSVLTfJBO8Kd
KKJeOV72+kC8oestEamgwNnuG1I6xUMFvsWKwVWid6etz/ydqkyTb4Q7ZF/HMFLSc+9S8khjnYw6
+tcqY8Ztxc0O2OtvMAgXRqWglWEiRyRtUEHHsW31t8D6YuAKADH6DLB76HquibILDXokYSdeSKNP
GqMVD/BfMRSoysym4aI5vqJBueqqfjsD57nodrvpzOEqpdOqAMVP+dq5EXrvWrbkkos2vuv5TjFA
seryHj0jzGAgeTm9cu7g0g3qxAVXEAAu1sD7J5GhqKuFgaaZ5v6qSyKZECd8D4oC4ALn+DNKHI5l
7Vr6DQcbyGVEmLk4Pe4wvlrsr1kJ0aME2iqX+0d8eyISW6CvnsX3W/PMB9CqKQY51nh91+PeGNLG
AEB8/2aK8KwRZTFbqirWPmfYqs4Hc+hRLvsLCkJnZmYc6y88jRmAcOTj3ApK0tabl54z0Isxo1Zj
0VkbwPE29my98WLfan27redOGqw8v5/6Z1ldSU7fqOy25J/gJ3/7lOeDsNBqhmIghE0XdUlJ5LDE
DYVh4WWQYZXPqX1SpCdu8OSBWK+t5SgiaeQgNxSazKG2DAiWPhLq+VfPAyyi/mMneoM7IC45M6s2
TGTxDtrcMqk+f6oZlcTs7ctJxvA66Iuve6kQInSK9nzykMp4UH1+t68UlisW7TclZa9kkiGuGdJI
sbabqxf3wijb94lw1jm8Ax0GXGQJUXOt2qJWOdUgQYNmVqsXEl0YbCjmrGyy3QqjZ9DUiA2nGTXb
CjdRzalc+5yu2zK2N9r3zuGxdHZv1UK7x2cMWVaggYA2cGVsBfBGXikPBWKDgwkpBOx4egPOg8Fc
6g6K1ekt0W+A+4rMyeRFiHmBbiktVbJp8t22S+W4qLzwvZBNDo2HT9IVG7394FszYBAM+jIQifDC
qkIgDeWZol2Ehb7L0IUTz726WrT/21ut/hrhG8LqIbCqaLpIN0PFRA43ESN5D7iE1Kk17BaSgHiV
yDrL1l+tlkgL0CxrhBD5NhonAukKufgsZ9BPDYJYAKd4VF7YTMgp4j1elB6ajKfiqpCPzwywsJn0
SGmOdQjGAjehH31dqGtuYxzNiPd6vH9FTf9dMMLUBYkzuvXiIMkDQFfrvT2bgCGWd0OHgXiCvTKe
FLtCEtOHZzQ5zT2lIfIAVYzGuQ6vQ0jyovbjKDibath3liYzARVljJkQNsivoOMhg6aj33b8nhUJ
vIqUFnptBXBjDUMekARG7V9AUSuKKtoI3UafzpzIYAb1FKpK12xY2unSO243CZK6vDpUid2mAqCH
el/BJL7gOCai1xcSbX3BqBE4wPBDp/A2p18KaBD56S8sx1MeE68bVH46ue/QCyr8Zm4mGv55X44M
F5YbvtYNYl8U06ERwjyYxz0q9N9yzhaWphBwx6m0Ru1VbcfYEJ6IzAeGiyB4uiZmWPYvRm7VvBKY
i5Immx9As39e89Hpu64rz6l8CS3z8Fi5GGx31JH120/VlNItT8QqYHohiYn5HnIntOuH0uhj/KGv
gk17+LqralfSP0mX2xUDAn6KA407sRTQBSfK2EuUUXmTQF2xHgmGKQAm8uY+bNKosWN9OJXpHcMN
p/zI7wPrUy852rsK5byxrKAgwA7nezmE8lQK+25F3u34wgQOCvS4y9WsxmaeLlUKTLAyX+tF9DFr
4TnQUz072+b2yJ3bseojB6BrpflrBUk0DEyYb8ymGOzJpKMZhpa4x5kbs+0p0Vs5QO9LvgDIP5mj
8CWgW+8DuYiAlYPAcI2+qVV1lCjq/GAZnWocdLycrn6xLUa44DgxsYTtdtaMeC9cFdJk4296+HFu
XZuMf5d5VCbSnnO5J42v8kqjboL9pM+AkvYhsmm5sfv7Ipo6nHCoqzK78koqAip+nZWKxnKI91P+
U468CVi9zxXI3fB5MjGAr97Mg+J+TCQdlNOb7VcaqifT8GlvVRZgfqwdKAGgvrbtR+7JsgX/7/S6
aIDxxHF78lhJW30jOF/jVPMYT6K2VFe91bgPGOi7k/xoW3C0dWb2WFCE+KsjzeOoz+rprI0kuI/+
tl92ooTWP2d0KF5/zPT8r7gRYsxmXHqGti4uUUsMcK84djUUKjFcWlYMF2+rR6Ywva5nyg7F+DDa
Ap+YYGEovLIG7ccSBXOgB/SjyPCEZByAmZF+k7ZjuLEsk5KoU31V3wh5ASWfXuRBv8pTtFDHCyqQ
vIj1jXaxref8l1yeOygGDTq2Q/gtcMdNcsk+rJBL+v7hJ+5VZQQLHV3jBqNfBO2TC+1OhUci7mKG
eGQtLFD3e8YiRi2PrMgyptqYE/TohJMbORPnweBP7EA5eUyYc0LGJoqwgSOmTS0aujvJb7P5YbMw
yFr0+zW4KTNC6M9uXPLTZrlmO8a/gEkdZns+0XVlGTK71B8EDDzHmh2RWfeK+LNA4sYNgj1jmje1
Dg7um3jer5sXqnlSYVzx3yn1GBXjzUhI8fPYl48KgY9lIFhfVWzwzwaJmMnxtMjMAiN3k1jEZP23
ppxoH9N7voxhkolRwyShRIcHucO7bzQFRfMdO2l6x31CTogFeOzNRX+ejD+JM0qGsElbRRJPLdUk
WBysCkHPzD1Rn/ajkliS61ddA3P1j0j3ZEtTVXe5ZX3UyBI9BUkbdJnK0cs81WuME9bGwUih2UYH
ec4sV61hWVe2sWPB+2eCRjw7dJQhPIXrZ+tnzWK95ce37C7LiqpBHMzhwRgDV0AtAjYvtmidsVNg
UPFQqUSQ5zXgU62wTEhlzBOQ5WUVRFTDa63lmh54Jl/Gytv7eA+EbXX2iUVp+/FOaVHRlgRaTuwi
0Hi2T/4GPj6LDjQ+h+dQWAjipDJfOzL3rqCqnUOIBm38iLnq8pC867XmvDEPB5guClySZxaMyBGY
4Jdzmkx+4+i58q6tZlmPel3lM9UR3rE0qHvzHIGgDP4S6kEgeuJSoSYGqDVf4lgU9WNI56MW43SS
xv++SnvHJCBqjiK44p46vCReG6fSzXwnYyb73fUQ4yynOrudVDtl41uWpUONuN8AHojzF05QLbX/
s5SSIki/1DDJo1YtbfBrG/9gyY3H8MGXt8HPo5BR0QJdUjynwpDm6emSHVUuu7JmUmoZbpJ/k/Qr
/SwGNXbcMvIcObp3i+x046Gf1CiMLq1Z/Bya3SN4v+Ppf1KuIVLV3j3rUimL+lskX68Yj7pZex/R
8WkEv8TshaZl9sw2FQm91Ez0e0UTy0dwDhDt7Xbez18lA/eXBLDgWxh1gojhUwy7dsy519/15IJ9
Xq7KKKfowO0JF1Z9funqd7nA0ilh4Ilr/l47wumRKtg/nPS4fHwz+QB8M8G3jC+eDDVNsq3JefxH
G2ILtr+8Ex/Zro0jrGbQaGzcRQbcD8eAFTIMSPerktRUYTwEYfxVHqH/GUQiAdaqm33S6avc8DfB
ZjlGJFSzR8PbvR1P0aJIQyhvuV+XHnk89U/jubjXTyPcxeEC/mpHLGzTiBk0MT5nit5YQKLKHH58
ODgxUFUqN6Ro6KNzGZSFCHUfkxDewsd+TOfDhbWnIhvYsyeHzta7s8MQvPBzrAIjwSYO8GYpft7Z
GxOM7GZxDz7MqV6xxOmMfN9Pf5UbVbPXj5LzlU8XB1lbaUwMtzVVBQyfha/FrSrbUxX2b0pzd9ez
ay28qG4JBPEwdIXS1RiT33OVVJtMHyqihTFPfvOqJJeODKhUCrQw6xjhHijZO/f2GZTCVNKuIX0v
CCFVzD3URbyJ028V5d3n9IMkFnn3uFYOzLvoKQCTi6MLAXCoi+mYSUdkI8bWQjKehlY+dOsA6UiR
bKYqLm8VrqW0KQBZxEOApkCJQO4ZWic93Sjvx8YL721I4cPHGun4ET8kS8D9ZWXhGkwguudigROQ
JdIrwEO61I4Z0PjdHfUhllDj7hKEQ2/+8E+0zw1py6T/cIznYOmjibjjw7VRbTFRhI7NCJCc+Kfb
zkaFNE5xKsaEUlaMSaNir50BLZgLt75R17jh8KBiQbUuc+cPlbo2aP3lUlimob4ypWDVku14PyYD
Yzqh39wGBJxqF/8+fZth43AwIAXKIb/G1gfqUdUlSG02DqojktDW4OCs5OQBLlWGl9Xr7LORj9RL
cGvvXl18V1w4r/VUF62i1oVzQj885yywq1yOoblBWiwCmKQfB+zL5rviUzaMUEIAXgCM2G5Ao4Ex
wrdgV/ULeunng43XgEkCiGxiR5t2mN+ow7PqMv+9ClVgHmBPHbQWqGkqTtqEdEYR5dyCE2LuuhC0
1MogP4olggha7oOyGVrWo4ODf54tp5Brv8TtQpVXG6rOWzr/eeSzPMBRRb1HUUnyzqM6N+I+9avc
F2GZGyHycyutup0klSI41dBVYDq7ILsKUGZ08qhcmVjqrrlGaCtuXeGg3/zwCEFcWCeLeaOtr/fm
yUy0yF/ejn6CcjyI6YsOKGTwHSzlq85esLRIEFBIEO9J5cxXiNNd8OCsq14y6GeLL0FpUbLKwn1k
Y33DsUItdDV2AhB/d8q3S6cY3oicfOqiv2v8KW6Q8y37ZnJDdtFVnB5HUtYpDWCNwYMLAS1ODJV9
JQzS4hZ+UMlhS+GpXdp3NcDQpVuUhKUuUKylCFz5we5MG2XLyhVSjVVtweh9CTQkFxiTw0iWzMLX
uE03/bHoWudViRQ7GoeqfVDUEpqggYdahiWD0ts8LokRTVd3uwu3zJOC8N7rBJgQnv7OvtB7bQ7o
hneM0VEQiS9yWww6/E39kF9QVP8wiGiYV9fQJmlss/+z14PF9jtTeWxm2qWS8Ht0AAjdDQm+0RVq
Zr7KPnqQtZDY9W9RbyZiT//qF7+NQmW+YsmT8A1YO3GgNiEXPdMRTBZGcON5mjDdNkF+TpIajodL
20qY9hhMrrsOu6wAo6K4W5v5PBt9K18zOxI3fFXkZoBQo+3CsaG0yIkbxktQHHVx8gZt89unfoAK
QGdWqCdwDcAi3yzHYljDwqcPxh+AlBGUZY+7nbJ8KOeySe+5oGy9l61DvwbHNJgL9LhswQM18qcM
p0O4wyiS4Z3vtyn8wfFWiop3BIjFqxrs51oqHie7LEaguix0lQ+/d9rMUn2fg05K+AT91O8FtV/L
HY+yK9w87QhRTNl8pKxnR+7rZDLdEqQqrwZ20Q8hc5LlR8kdKfMk6Kj2u2g/eHc6t50DG/66g9Fr
FKmHbsH4gJP84wMU9AMdCoVU/eAmeBJRKhQ65K3aJ0Dzs7A262r7WanmAS0MGHT6fwTosiiGdIE+
Vl62KFH4z4IILN+a0PlFmfI1YWh0PdaZy9I/j4zHYLuIbzNnqqDeZ0SzFzrVmIuyErK0sQLmclcR
8d5IDV1EE58J1po4ZtHc5JB9W+Jrsu3nK070atZY47ppJoU2yK0HXYMQfHXIpnQDxbE9WAtzFKjK
7H25/WRd1tynPgUVgoHzXOMNVVCo3k3kQtjEDGvrdHGyac15Wv4i8A2xYl+tsop42Bb0RMxBpDtU
EU/J1iw5kBv6l4biBGymi7ZPs7KNNLOCcJaeNajiY/fxTEpXoITN7JciY2FVjSrrZLlCa9Q3sXWj
o1QTMrvCwOaZSBTMQaqpmBHvZI0pO4/pePQqwEWlHFgWp9HXjY2/oec+Z+RHYo1QfgMwmhKkGQ1W
0RebNowhh5qCwWZgW+YU5etpus0JZ36G6Vy6v6bgLymm/M67aKJrTW68GBYfRCnPVormz+FJ3B/Y
d/4YP917T75tspj8BJsOZZtpNE9fHNngEqjrH/IgboHjg+7A1E6SVlYi3hE8/BfG9usGAoTXl33O
pcpJqyTyUvKcvztUFJ4pTIfA7YZhT9/2+e8+KIbnxc4GWU8C+IzFsuYNmgQAdobvHMfG5azasKEr
+AmZnWoHdeS7j73rcy44XmppLDHcEBXlAmZo09ePc1qyTiSBwwGKQL+iM/8CPbgudbrm+0OUsaOR
56AunwTYeoq9HJ+j9pEOXvbNmekhLCl6MQ6Afw3WwMki5KjP0ip5uY4FuHmiQ6DgVzleazSk+BBv
OjGTLm5KRQJcBp0zpkaMULufZNnEiW1p+YV9Fy/iFEl0/QdZIgJfXqXVQ7AiO0FSsZxPhDSa6M7m
pn2dRL+0vsrAtiGrzu6Fds+uTglePrr1Yhvzm5PLN8yc+0GqC/VJIfRngFUZ8Y3x8lHSIdZTtMwL
JZ8BhzMk5h3PMybgr436/P/3FqxoGAqwXbLRJqep92CcDGuiZM6hvGw+AGOg+irv0GCNGGMiv24J
Qew6Kwajorqypgell7Syub9bUyWYpoKkT+kskA8WQzAMz65jfzjmka44yqr7l9z5PhoSsUamLOWc
0GYKBQyWf3O5jBA0FjFh6lTX2T07IHGkBbcozaEEIBfw83zWaDrIirOZrhP2Lku48VEAFmojQFBI
gB3KKGu1uonmKGvkhDGes8cGKAb9ID9DGauzBjRz+XLNc9y/+lox5R4tEdgEIjZ/ZhAHv9W84ukX
VL+2RcIiY6bR110ByPjIYiIqWZFPA6NLIaq9avrVytS/ZIf8QYYGbb+7a2kSV1bbdNVzDYXj8cSL
DiCVv8Y5HvxPmFoSUfgiCQ8se/ZiQWse3SFVmyrKSJ9xKxHb3KX9KyZNFeL8/kiijhSEtZzNapjr
goj75LV+chV/5ktS7lR/ukmjadi8dS7EF0l46xGLspANoVPzfR8n2wk1S0s+/IgZa/MKALO3p6bO
W8pzODVb9VZEKqe3/NtcMNrjWfldX9PLJp3MUC3uOitSixBhDyTdEbnMG8/wTygCb7eCQ19185pK
UsxpQkaGrx9MHrKR59xmmXgt5L214V0EYZwP2RKZYBmW/jrWXiZx+FRZluBwTfspBVs5jrXCytw8
x/ZeKLUKZ5OS4OXqsJhy1yxCQNva4ujLyCTvnTiYH6ag7JYRgv+cI5UteJ9tGOXhk7hLhBTLyZQg
Y3OykA3u/XskPkOX0EiK+bHyDU/p3C8pCMYOWeHkIzNkjHZ6YwGu3s2k03Qkwc2+zHCEDXdSWoJE
weMI+9QtcBhU+9N01bqilb0+5aRbSIjj5+KfAGQNI1O6Z2C25CLkawgaQpGFKfR2NckuvAZD6nlf
2+d8KZ4QqnopGzM7pPAImzuu+sdlQqk22B+boh0vuGgmRn5CDxLfmLWOYYLbs/NeYU6No575zN0h
3BQcpRquQQ10D27qGXdXZRtfwnAx0UTcZF1g+KgkLPdNnpd1uouFJb4jiJnqZpMkTokEWcQkYcvw
y1HcpICaVG5qE0TqF93ycJO7d0c29RAgkvVOXOQ+Mmo8BLCa8Sh8kKMMind/VdZ82K4y4AuLRxw6
7diljEh8uep/B70efYQ3bDoc/gm8UWlQe6QNrP//bj2lIvXXwnawWjk/pXTfQWvZPa/1NHPMwj4h
Sj6Q+asrKVh8xUoPdELC8h+df4YjtwwiVi4WKsD/1J/SyatRkuusQeQNFehqbnVWo0Q+NdpWZaSq
pdApQFi9EdLO9rY+N9IBVBUqDiU7KeH4pA7bQ/aOj44INWYP4KDyklG5YqwbTcFVLbs2cbQhK7jV
gsVhuBmlxOX/ZUjlI80hmBkuJcwFLfpL48NOExoq5yKFyc80ndwpZr/HArJsNYLRS5Z+kXRH+hfE
cPYzEUT4w6U66asviMZpPMnmxqOUx4urKMSwaa24sPlC8of14O6G8z11m+9IWHuPCayl/+q7lgdp
TUCX5qmP2PEiLnLRyDCkjzfm+jaxVDXLccI4A74QxZ1eQQZBf3neT6ZIy0/GDZCRMLdXRK8MiVgg
UWq+tH31s3pU6yqoSqEy6fhkeGVbxZCx9nJE5qZ7pxiosA2YJhmJhEEPDqJ/v1I//vl9/Isp2KsX
GcosWf59Q7csLT7PDLswGMsLfIBx2EQqjI8BoU2NnQfLxyWRS2M+ag/UbGJ+m8cCpKUv2r+MlV/5
RQZiNmZbGCWCc/bmhBmsSglFtPPo+oUyrtVmmsbdjtyUbyo53Wm5MO2GBDglVE/KRXquHBeO2aRM
dviXHUdTI5rfk19W9rYD+ZjZwy1ET19rAhoTei5PyReWN9KpVQNhnxQeQIqy1PjeDItXyiROrYQV
9Qexm2TZSxZsIp/hFaTYgXJ+CEp80Rd1uWWTSD1bgmeF4l+oLJ3sm6H/ML1pI2RDFCyFtSgwSgQT
w+iLkhreOCgz7PxcgcNFYjASNnxfSuq/672ya9HFCtafuRWI5VcxpLcQ5AmhWE1aFgpkX5mvs6oy
SDsyaNZa/W8rw1vd+ON0Q7Tea6++oJKjEhb2rk5ggHAbDRoUHYwKohq6I7UIiE4i/vp/TDHYNFQg
W6kRX+k6f7ibJsrTacMhWg/1JjQihwsIOmdKTzcH0OwHtIW7aAFiyBbTRMjw/Dol4L8Wc430GKWl
cLUKXdwXRCF6AHP1LzN7pRzWm45jTpkm4a4QwApG9nlgpyYQ6te4YGTpUXIt0huMcNekfig8nubw
fExZnFwgBVvCxDnXsIPSeraeGoc2WmReARxyfmslBeqJ3V0D6EjVTu4Y5vUBqIyqP6afhYIBtIuy
V1HOCNjYyqWNgJPiWEWSJ1aBhYa6sWL9W8C68lqZsj8kg03rvk8hjshbncqoYN6hvY1FhobJ42NU
xN4MaZe67H9qlceWnDRh51vTK6bZzxk4S7u30dCMC8x/eLTOaP26A6QwvZOXJHCXIem+IQ3thGXn
ZM+Y6qIt5do24SbMeOwBd4sP4/FisA+rY9/51dIHzX/hNTONrTDfGT+oF+VYGbe3rBEqapLniI9j
IRxC41Jbcpchn24BGz8Hx/sShNUpR18Jl+zbvft9vaE5Vj2cALuN5Dt+mVxQmc4/7qrnXWypqHoh
yKTI6wu4OoQcvoIvSqbnKp4FuiATzqssGqMW4QXcyb23rrptSR+OjI602t2lhN2w3SMccxajpT0A
4Z2EIESICICiLfgyKMPTqaSokl9XkFiRckK0y1vTQVgPvWGgFaPFnTFwiXDL8roUKiJjeM3+p9ds
USHbhDqQG1KX6NnuBSjy/rG9OK7Gqc5aVWIIAu0GPnuNEAiwJvysdT9VU9tbjOrpppoYpZQO0hdO
fNYA7uu16ZmXivLgXBhoQQIYL5PmGTOS5iCTHIjM8K+JlAC+PXID2XtcbtGpZpKSOutPuPlk5CPu
KjlbBjAxjLBz3Geol8wsqEctysmHalDoeFz6cM7v/F7jelgXTzl6xeZpQNWZO415RT8Ie1vOoIX7
4QA6NYTpTmZ3J9F3COUoa+LKTlFi5DL6Rgbt0jGBy8UET7hHMprYnJdzJh3BzsoNFPeMwJHu4/eX
h8T6+R8SRMDom0SfhJ+6RfdTFk56yjP2KjTHgEPLf19ZhXSUSIO9COrnrlsk3Jg6a91bpbv4VhKR
5CfevIh08VpKmEFGK/B556Ry6pn/k2X94Mz6n4eFxK5RsOm7+ueiYruYM1QnTVdUAclue2lsHItC
/INEKmom5kFfsDQtM8Y7yexT8hJrjmUFzsMKTLK+0yM1Y8jL49FqNEJFW6Xty81BC2w4yvdJwptV
j7inQPuhaTzim+HTouoZwK0z5S2JltTQzhrf28Cab5h/QS+g8uqKk/3ssUUdf8RHoIuNZDc+MDmg
e0hcpdocjPTWlhx3F2tdMOUSpzWhYfmYHY3KeU7KGAXfi8nVA+NLmZ5MVdnmjfiMnxucrYCbu1nq
5SKXkrfH5+By575qFdk8kLUtyp6x4VWengf6QTNiu1KydJQounOBdYFt+PE+6mUosaI/cjfcsUBT
tc/4KzUo145Faz/TLFGO13i9BdzlNlLgl2CpvXgDd8JeZSQ4C/Om+cSxBiSDPws/IM/dqzmnQhio
7bDn0U1XSznIcwjdJ2dsUtiX+mtbzUZS0ACQnDmTjKvRnk4AguxBudEkRaA1U+mSgNENSR0vFn5O
9rAvpu7lEEsU+tFJKj5iHwFqKDr/uhCN5D6rY2Um3esdTyh2ytN/6+HMjZJFua9PJnjFwSc/wN14
DxcgBdVV3038eVs4Dan0uYNWJmQkcbRtW3o9Rb2hi0xROD9JRuM9KhyzBsxUTN5wY+26pQ8Pb/Am
nEHTbeOcX0PVLnCxvypJNkIExPRuz1aT3D9ShAf9i3qAFxSLCmWM6UsP5ZFsPt1o32VDS56RgXNO
TFNXD2R431iG97WxFuHCUVRHXRuL0b78qROS4+au2NsHBPKs/w/SIzd2Dsq3ycDVv6folCOhlLdF
TIa0PRrh9AbBPaJiNCTV3aJEMHdus6u2IOA/fa5UdHNQg8GJR77ZV7V7qQWiqdy2heciptfkS477
sj95rLpYNEHSSsM75lYwpNel3HpOYSmDCVtjUYnxCz+nclkWBaQcRTVIGjM3ohlRQXJXhkpxI+/P
7L3BdBEjl7NJJpAiQMAmC1VT/pPBzO/f92s8bN1ro2XO89BtEpzMLSPv1dCO0yq9aA8h5CKnaNsR
vaJvL7nxBpO/keZ47SyukacR2Dki+pbQlFstLO5vnZ+25iaMws8572VQLE0GAae8NRnDU4ylEsYJ
EYraGHaPMD5p37TA6OHXZhdQHiAHC3hVKmT+YOdQfOJB9/buSX7fHqUWXYBbssnxCEFcEFGi/mSb
bgui2Cj9kWMSdZLLeLMvX3IbSmm7w9vM8OLbhuRm2CNph7JLFUsyK/y5Opxrq5wEEQpYLeK2I11a
p1FUSXg9MGAPpRVZ8k1/D2JR8UUn0GdI6GF4dgax2qjbvDCVTPK2m/0EbYiKVe+YGOWpxABnCeqj
begQ2TTXddoYNO1XhgDIaLYteiPiosQvDhQoDGZwKXrbg2B4W2drr1ccVS1ZQFAGA2IXHz7yBBCQ
aVKklbWOxcqoeTE+lXVjkU8TndSHEN/ditK2EUpFp/dvim7SY7DnxliokxLrGi3dLZYf2aniAVId
Dz5TS0KwCrt14DqYT0jJmlTFzFYfcagH6b1m4cQs4ULiGSmtVBE+7uFWzbFGS059NLh/s1TazKdq
TqG9zxqnPtmxGLkpQpx+MH0YL9jbEvxzjgfLuMQyCsmRmDNzxl8C/5dLeM0/9DXtBng0GjhSGKV6
V8c/cV3kNtO/XfW3KaJnrifpeHqK7lqR4Wpy/cl3Gn9ejmIcbtV3Ot4NU7B/ARWC7x/pDxja+y5n
i27EYMlo+JVEqkEKOggfq2jCoR7t5GrXa5gii9vN/pFkhAZWxnSzh4jDWZrKSDPOo73fTjm6dcdT
zwlpMFV1fihDc0wPpXKTSdJhcs6We/3DNbsMfg1b3IvhZo2cEZDQHNI/f/NTr3zUJ+T0UYf2mmeL
SQL/Z0SH5HY1p7H9l9jOoFQlr9B9zefpR0ZotYAGgLNnCeG8/TRdi4Fus3k4v+6XJ7Mh7Qxj3cRv
yyHopBIr1HcF8Rqp4ZcTirIsqajqQBebrLjC8oN/TU2PIkDhr9PoSGGkckNh5KBiIPZ7alwPi9Yb
wdvdNZyRwCRWqoiCvHiRZRMoROWFJcl0khBcF1jGmq2Y+nJJrXd53eI03LbVAnx28vjS1+XLAmJ/
egawrD/7O5VtmYRUyqwtKNBJBNfxD7MrIE1mImbg4mvKJ8KaFvT2NZzpvds//yoSzZftFdE8VDRQ
XNRhPzAdViHMETBEPwpz61xkdgufqHLrd4krDU/O4yvBkecau9kinzCjKn49/KFpxc5mOmJ2M+os
yrQryUwTDmIACViKrNB/My+hMc10i278LmWSP/LxHto8dEaCC5vYAWe3/TJ3FVZAcX79wZKbOYcl
+OiUzTXmxJR4bZzKMsKWpyja9t0D9SC/jsaJa7sFBcUOPPrQSYqOEEOgigH8hm1gQw4Tyk8Vu2t9
Qw5yvZbHgthH3aphkve0WpRmh2XGKA+G7xP12axzYsxEKNDni/9toYXSynRgcmZghEHXiDElKMFG
6Ue/ukBV/zK3kM4Et42fYDoChAue6TEs/F9Egcw93p0ZiFFvlZGqBV23BbiqbSckwM5brrjZewVZ
7+Y0g2/QxQibjolvSsudZg/8sQLF1x9pHkmJEbwOhZS0Javj5f8wkVcUvKMBcuZc6RQeCpDbEzej
JnnNm2EEarx1f3SmZb9nWv09YsI4XIQQvChR8S26wsgvVbfxUADf0t8jShGSa75CBxy69XN9mb4x
yKw8/mcjgRf3a5CQz4WDhhyaJZEJFOj3WrS2dVQ78sbb7V0pR7Mcop19vnpMwH48jNdb8f50/C3Y
CbQj623jzTQpf5QZZ1p3bPoi1VRkYWK93gp+k9n8p6wlseczVlwJZWx52v20Dc8mfaKUBG5EHySL
rOmqv5pR1DHp3Sbx+1gDXCj01ia0I+3VHqQXYKFfW4S0D2L75k4c6Rkjm2S+M2iYTaW9XxNgY3lR
N4QCEqY3oAFb5Mdrc4rJTzz+7KLOlAdaPBivZKRJWRuURezhlr90JRmyUJjMU7gkdcw698CNCImu
MSy9FBuGNSEIvULd0t3bhR3NIVBiv+/2LKCEtxyhRzQ4CJsVLrGa35dwUZSOe2NXzpPXX53iOjUy
0XRoJFhiz541mKImh+h7PntqUS9M0XtmWVBOtx2QtRxa2AXjCMxqOQzfjmmEZi5J++cl/9ne7/QH
fvXuTV5inxgFnd1jUp8Tx0INqhDPY9n3MuDhy8kSgUBLX1sDo0yWt2eKkQWOybUmPZVRjOK+u0l6
5ZdisRTqifsZkSs/jyhWZumn+2PhYcZcEIDlEoJru+erLTnFTEV+q+njlLFq9FxTcdK98uulRWSK
6R7DvyZdhkAsoOwhQkpHPM7qpY/+OCH1iYXojGkKuA42yG5A3JmhdMxO6gkw7G6grJY2buJkTeml
Wu2yiYu7Ka3BDgU2JtPJKGmgrR8jZrEQDDi0RLptSeOwWBObasWXtmzukMAy3J5/8+kPSJpqf7bm
KlSWAoOfS7KbH/bzhJD/wkLH3pmGLmvGQlhkvgZPdWmkZEvj2yqnCkkBcvUhQJccBfUFz0rQzI9m
NumgKcPXql0kGbjpT/hWcTEc815E6svvA3O+NKAxrdtaFneAT3ATzAUhsMG5AbSBGNUEEjmkgRX4
EMzgJGeaaAfN2errA7KE1Fu4ZRUovN/BRSANfmDkbzCVH47gkQV1soib/XIq+on0Jz7x8k3AY8A2
yXo2yZCN7k/2QML+ntjvjHJNM1RJbGSdLh0fMMbJqjNJ6+4TSf367bbCKoClEJNW8iNHq4AqnBn2
RsNx+iLJVjBEV+zogg9Sr3hYOr4N7ikSvmU4HlQBILKShKpwQjjcKKRGUhsDTmtDUJ86hEberLdV
IVZx6kdZW5X8Gz81KhAiLhqOYWTOSkMVFxndqoOo8vUXE9gGnZpBtKAyqMpjPBhWi1otGKZ8p9Yd
gJkS+wh9odS7G3/ik+mosEmjMfcZzrmZ/sAIncUCbT58J736fg+d6WaoGZQ+BwmEhm7MBIKq+dbQ
ra2hT75MnaK5JKC6218Mtxc1wz/TP53b9RmwUUjxlZszekI/RFBUVcpVv2bJ8ZOrUvbLZQzIxxoC
6wCLDhH0XjWEPkXqXrTiAAsP/daLtfWKex/VaoBqLwMTu9tApdsXmm2J8HhtAVg9jgSFeMgXNej5
BFr/WB3MbVts8VJ0ufgl3PxG/K1fC3nOjhCKJoR5k1AaJz2L0fyqfdF7zMY/KAQ65C3rajN+FBw/
xWgxbbR0Up6iaOt4eYoQnt0dLpufYAsBQgNyItVE2PH+dAWT1s7VVaxzAfo3rimR1CATOoH4dZFi
7OywIIUKghan/9q0B3rT9CTEdS1vb630Jf5jisBtF9H6PXVXy1ACFnyJ46dGMvqzamxO+faV+/zV
d8L9GohcuEKC7WLiL+j0gelcgtkMy0eGk+ZZusZZ4GBuR3eicfHmKx8CxIvEEHlgwBg/cTESe968
MDqN3yNJ9ZcI/69Dc7hhH3+5NphfUtacW2bnpRWM97ifCIx00OEGuRVSgBuxQXDqyeVTUkBxZ4Yi
84LoK2jpM3QJNvQ08cRzFpF0jdiLo557kY8wVta9fXSzl3ZlElu/6A5JLjQ2K/I5SoEQ7gGwte86
8ut2L40OWZVXm2GxPRebDH2178cMKIF4E7oWgeVF5aalg6XPSnWK4AFnfXxKF8wwOtpmkZm/J7cb
ANtIBc8amILtUMQPnHdIUY8tslv9fa58YHK3anRl7i37bk5Lqwa91WxzhCCXPW0QtA27B6Xl6gRh
DnOIB8RB6mZjjTELqgu059R16sszOM9c45wNCvOkkTEabsNqRTP+ex+HTzkeRjMqYbTSQHaI6tj7
JvRwoGUXZPYv1CxmF7e5aaZfONClFeYP9/SPoJsR2s8wdzvuhWfMTfZECzmTQ4/l77Qc3JIAdPpy
5g9B9VTAlNlyHu/SSgrnryOoRWvWS2QOC27fGk0w/DzqvOBiSsX6i2/pshWxUhjRR7Kp8AaHO1D4
y95Hck5VSI/5i3CZYaZ8P/OdMRK17/0V2tjzUrkuJsze974sqhrK7fW08FooO/f5P9cCbF2FmXN9
DAwCI09qayELpk68u6CDpx82FQSm5OO3fn83yB/ZRV6H4c1pDjHmDhhXsrpi73MC4QGlnyVQU+Ej
3Pcs1aDdwgA4tX8SyqINIQlmysgQ+yg+XzWKG0Li8Ma8xCCUvonwNbiR+zr3zrbh6i4C/53E9VSg
PbUfTorqsY+vgNsmm71h7DcFoJu84UP+SdtoItotlhlTnrjTaYMSHfF1P5IM310yZSoeSHt+u02E
e1P8tWHbLtopY5GKELWGAjj46J1kR2pye9aEDHVdoAiHfUdHPcO7UGtsIJaybGSmFfdjsT4w2ifp
WsCCricKK5ha2s7QQ06tJJk0T9pKZ3RKBeFWi6GXFrcm60J0OzhvBDaf7ydYGszdVcX2+3FR4vLV
7o9al/Hbc6u4iFxlV0bCRQ+kwZ+9BWoLqvohSFydRq4n6NhaEbztkWEXGOU5DabmQSMDAUfjFQR/
xb/nG10RCNpEJytfA0kH4hwxTJarME2+8w/FRbACYjSHH9weKAxA+gy/gnCMAmmrtPRfg3UkQqu7
UwrVLe6D+Cti5TMFNPRvNYMMTPS2mXcbVtDRo8jhn3TJnk9QapzKRmysRbc28Kmv+aWF9VpTBrbd
uEeB/7X/WZq4vTuU/BVOPw82d6fgiNMrxeOGMyY6HBZ/AbyVBXIvoHcttH5Rq/kNaP/NI+YCFF4w
NacdOuzG67+UX3UzfqeSrpZ7Ly3vC2WcZtZqFJf1bSvLxozMrqVUWK6H5tZpWDNs808djmhiu60h
tiK4m/hx+aZ0bGDx3dyGaHb/QNlRivKt/fK+aZCRNV1lZij+qk6H/k/zvNjYqJCxWVojPXalXFpy
BPCQ7aMCp04XsVMQAqYd9WuH+lGnb/Yk9I+jmJy/9cTWAkUgKaTBiK5AiJQwy1+tB/jndX7wh69G
miGCnA1FIRYcGcDZcXPdAy/GPGUXGphO1Ghfg3LiKBQBZM2sO1SvSRyiNHC/vH3YI5nCmE12QoGa
RDS5rNOyfkLx+C1JETb70x6ScX/ynz+HKkRZVQsneuK3zvEOGXyWfWo2o/PM+idjMS6zuksz/AOQ
XqTNTQzthweIZGw0ivN7epPLZJJb/GKyLS0sBdU7HlNFti76N2c/1/NMNDBimsC6WFW2AaCA6w4c
h98iaxhT+WxrxEBS3z3iTpAeptBKWpDGt6pzva6I+AsSttR7uBCeV/wBxUm9PP9jlJIEjNLNj/Jw
tlfJKNMoUlZxZPxamtdmFDAlVrURmy9v/wGFjSNVWayQGpHjfEx8JeZKZvaGLj6X70hyQSgyMB0f
P803C8ieCXBDt+s7YBspCQzAwOeYuVM2k9i3MeVZh/vWbqT5x5XjjToPiZv+LirSHwlw+KhbAFC3
Ge/xy2mqn0hE8oGMhJpcOhpARNpTR55NgR/gx2EOG1989rxmY58RyNGbb2hk4ziCZPUPdu7OW50N
ivWUI2PGtdGXoSqm80vXyF5X5yB7wB2hXAn0OVBXciigQUuF7BYggJdzAIYRr0SZ/EIVcSi2jHu7
K9WMBPsobf6Lx9tx01vt852tX/l4TORzTltLxdW7F5buE6DekIRywi/pdHN9ltzKe62m4MUHGf+W
rvBmHRglOe4hKcT2FNwC6nKaAr3gIePjAIuf5vnJIxmMpfKy2vPOTRkC+eAn69IwbRHzPB5FT8rS
HFnElUFc1twgAjiPkkSLfrFpGKExx+0WTmdUcnkD+ug/dF7r4s5U+H0tUWBFZaRBEx2Qm3/zZyoz
Keo/J8bcmfrg5DRNYYVtpa7ToH7HiMCFeopRGDQbT/381BTsza9f3Eb4zkNKH3WWKmGbajGeALOx
nQmgybI8MypAFqvopHZovU5gzRfxwqVBtgj2cKRAq/Jc9FRU7/LRwnf1QH27gv6RiyPNb1WNHMtj
+iC0tUg4Z+Hqs325D9IFcEZqvLbUUFtLpSz6KDTuTKxyqYhwfuOU4GLChRUPs3eF63McbvX/xENU
skbYtsH+9y0kpLl1Kl4hA+J1bp+TAxAQtv/tCFHXYXUxBUHcaIn6VtaKCkesEah9Yy9gh5lu9cSE
UzzBYTCuGkeAyBGMjRqt1P5XQ3NmGxTyM3CSRkWPV2ZTdpn1x0c/kjpDSpBKzYhwTBmdob0yRGRE
8iffK1p7BE7Z0AvoT389ytpomnkuGfN/tyfYG7QDfZ1HaF3ZQ9nuXwJW03ckTmV7wdCfWhixkV4C
BM5sZJuB6qXAP4DjHQZRUnU85OC4+D/8J4zkZJyUJSfV8WMwIoeNbiCFtLOytMGpuxRSHdF/g/ev
Fbixb9qv5jpu+Z2mjls/7gCb49BNyAAOYtDzqHOlkcBi2/VF1jkIQLNRPpSPgdHSvRA2BzDNiLGZ
/wplDlU4sIYCQPhD7gUux77Ul2fXnaFjN9HDMKO78kSVi1efyVFCGsNu+p1y35RflvMEUzyG8OHx
EvkiUv5GZfZFVdGJPsFH22QdImrcW7KxoNOFRBiajzgfYhdZItuE0NrlCPG+hG8gu/zrvrlElyDs
MUBc7DmjMONcFs681fsgvGey5brA33nNu3aK3ZJT/dLV4t7QZSNMA1wqacRXCjkV1THj4lkHRUbR
BEoSRn9LarfTX1GPBFCz1d79IdFuhxarwcZVgtpEmOkqSye8z0vGyuCFRYCadlfnE1GFsm0SXsT7
O9M9ZuM0lWRzGDFki0AjmbLfLPEyajiu+FawsMIvoyAfRUCpGb8CnQ7ZhXDLWyHpGVzUMBMcgGWK
nXlxb3T3OijaoWCbJVjNLbOrgrHeTlLNFvPYZq6wuae9r1Fh606cG2dl+Xy4E0pkaGTZyNyFAw35
r4LOVjD6MlKVppHuS1rD1Vos6tdH2lwipA9HJ7lv6ZijLDf4g+9AFw/9k/bTMnWWIvIvktYCZJN9
WWZaASkNVnVnpXP+uq1yOm5ryLrcnLayM6XI1lUYw84tYjxKLHexYBuXXByH6q9jtGnSx9Ix8FTq
rWbZBYrwT87tnrQXmp4i38YQqNaN1vWkqav3F4b0UBJmQM2G5z1JbDOnW2f05GJj74ysb3gdrrUu
5SDLc8zEtV3gKUV8H5fYSZepo7B1YXenuuY3KDnF+Q0Z9k75DtALF8vFg541a5fdqe3DiqruVccx
YIyGw75zp7QqI3n8IZBKENmZjbf5ZyOl/7x9ihM2qTKoS72R//gAooqqTFE4+jhX6BGymSixPQiO
bzRyKiAMPqZWpda0wTRl7CAEhXBA0ltHzGokzX2dpaXtsE3Vrx3EZQzjPyv4LTVWaR26HFklx67I
49EF2z/ebi1QPXNk6Dxp4VpDrWJ2IWI8Rk2eR/UJtEnno6qufTTb0S+Z7j6T5rL0CrPFdzkg7c09
IZFuIlh15Lh914Gj9x5LhoCm7PkDVZzb7oc2+1kDIno9YatEvNVk/qdGe1N9QYkIruPmLjZQxab7
AUpefMBR35/zfjVU61xDMrEr2ak8+QCa536f9al0AugYFBqygvfzOgZWwTcLh+TZYF2Eo9quDIxk
KotZxx6bAHXj74rEH8IV3R11bpKPrs82jKiTKs4F5jMxIf5nCY13Qqr3AIFY1dIwuX89+XXc/yhj
Cxf1+vc569h1mCp6MZoMVXODr92f68+iLJgemX3KbFKsN5R2+96TnwkfhGs4uk9cwXEQl/T25lL4
wE8SVboj1PJv63cl+dTwkF+TY4F6ypR7HQ/qiXztYsj1z1g6uBpjaw1/CSOntGJg4M0xpOWRVZl6
UAbs2ZZjB5Z9qeM7quaVYK8Efvmk8681RMSKZxEdGi7vBjmC3xBOh/9DsqvdWOabOsmBOrhNW956
fmAvQAWtDcLJ/wFxIBSbdyHbKQWwN9AbSpTMzP6I2MPc5gtFzZnOHK2cPCMnP0fJ9qhvTv0sAydH
KvUrMEOHH2fGfbzg8v499UlsTWlb5MoGjd9KppMvZf0iFsgl4HH6t0yduUhYJ7TqYYsmlRGc4Tx7
hiz8zRSMRwk/+w3iVznc4FPvPmabq0ZJLEOfGpQmwKkdS2HDneGuBNPBFHFcrVheNJIXkrWjLspZ
Zn1vpfppZ4Jx3vwRlEWI7MtTb5H7JXJMfk+W1WmwnVCbHZlAuASxkhAQmyBl4m3iOWNoBui+70Zm
CR8WBjC/GoPOV8MnS1a68OMYTdgrb5TSuJIl9u9p64vvdH7GmFN03Tno+eey3QkimbnotGKqHAM4
n3shMCJFN6AFwC9NVVjf95p2QAfUvBh7rJUp91Fx/+TJroyfuGWD8BKicPCrbaXqXd97autdGIc4
a72X9IsnOnbygq1xGX9Wdt6HgFzBmPh7DwCY5mFP0u00q0SBt7CnRiBSpCSh6n+G41d7GmSbl1TA
u060cBsT5pOAhrc6ztp9PnawHlyb28WSCwbsfNhEQrABKg/PH71yF8BcrnIQVplwL4J56Qwt5hiu
lbykh18ANzWKbeGRK5fXET+LSAaCPnqK6jxuIOQsh++9crRZhs/wSz0nT4aMLTp83DYnH4385Oe+
dX5yn8xESFGYUusN0gJFfls4wZ2G9HuHB/GUCcsoTc7ncGVi2bfH6Wrxss2DRxHmWuNCunn4w9Gz
hkQTFBUT1TqthOZhFQunP8D0onETpxgBI8aRHsDzCSgKZZYF8nMjUwoKebpMxZ38RtpH8imiZJ6C
omQNT0icyq6Mkk+B4HFSIhKJTodqiOVdPRSIWpzckdZxA1NiHWUUmBfBLpMfvdURa2OSRl888JFL
VhPYrnIo85nRcxo1WBKNqq3WtE1zCk8kw2QucSMrhMUoOvv4Ksc/BixRHtd+mfWaVYLJVQd4neo3
rUA3h9oWdMaM133ZiP7uCQ/hanJr9xaSOOs3KLj5yU1ZW7tZsdVSf53KjMqycrtfY+9c7L2R9DJP
dPhAWFvv2TgyL34QxrIRGQGFb8wXe8/kxsuRerB73GK/Jm/oq2Xt7nn1P2KAKA4X9dj+pak9glA1
AOYbAN0E/fV5tq7bO7HXt4lFZGNFN7QcVC3m5Sms49hkG8BjAW2j3v+v+DKLgTCple/lI+dIB3J+
eymCg1Cg4q0yaNvAmxkqvRrLRiHyHwAAYoFGklWGKzfel6UWzTgdCz28kL3hn1GG4dH8sNjaZbHY
NwnkNkFUqBgJEWQFjxaqTBZEuX2YcGZSzt2Pg9BgIbqReWqczPbIK/FWiPShkPUuU3aRVEIS5RBe
r6/7Fjy4gelUS1MDrhaSzSJqX7ABcqFoJJb/3qwPP9v1LejPQrFC2Uxnm5H1dsd49HOr96NYS2Mg
xlMbQQw58csOhyeZ8A2OUbCUlW+kpKhG//7BgF65kArEYwSja84Iu7RaYKIg3Y+ne7egzUMLDIgJ
2VpZOg6yFBLvXyvwLeuqZHrFtjfh5f6kg8tJ6Am+zlIozSa24YwNKSt4MxMy/xRAPJ6YOTT9+AXM
l5nQz+JImADMcT0W7KCXQrq1TPJSvGwMgf3OZMygKujbv+naCRBkxKUZ2iGk13Ai1tFqv343edfn
oMm0L1eqnSoHpuGlwqE8+hT4kb8/aNI//bRAIHoUVKzIrD6Vj0Ar5XW1Yd+skCDNg7xm5Nr+KM8K
uajytKmj66XqlaXQa1rYVbsAst79tss1aJKU//QXX2VuGlwBFQsI3nYX7PBd3Ny240sHo06yt8rj
rZlTNkp0V4uOttSm4YDzX8hxSz8qBGOm098GsGqAWBNUGsEGHoa9ZhwxkBKr9HPMl21B1s04JlDx
i5RbBysRiKmGO53WMR0snV3pONpFds2HWYCGbLpCA9Fs5sHJXmVlHHUDC1p/R3Lagr6dtBAj6f5Y
SPEBEf7kdfW7iBxglEOlnyR5CnOtGSy9u77mQW3bHQkuLdPwoAzTSX6J31U4XfKVjUHp4U/9y8Zb
5x8wKXgfOAHWRlLcC35bOmV+bACRNW9V/CU9Zbf8wpCvsGuemIekATAQkQwLVOrKJwdptBgiPAtT
I4UVxWF7vvwjM9BY3agZNQXkb+EqzjwXbIvF/s67KLJlpE0mJoqci/vFWQ+9cZzDU2M8CFp6wHzT
yZzTDeqUUIfkYnQTkdK8bGNJIP7TEmO/zjltA4A/UBQOIUkpWav5bDixlxIMkULryIBF/xnQcr/a
PmbjgJglQLLHH0USPq5vQKIyuRjZ6L4izPxLISB/sq47wbHTXGj3AF1ix5kCLel1KK8IUFEHRZvk
y7QyHySGhF0qyxREqKfGHzGVITsp7eIIW3Sds43l6wmUbwUerqlB/DygqiYMKtdUUcNHSaT6i8u3
Q5SZzJyKWKzqViQz4zSthendOkq8K1VEtb9fGTywcSI+j5yYywQGeeRgEKLONqNruMX5KRRbBrL6
UoxDlpa5SY+2k+fGnGS9QWDgymZnGdqX5evkQTAL7u969pWcxkD6eplqwv/kZWH19v9hzWnx0PIx
5Q8z7Rc/0tuMTCZ/Q2zVTMRSxLhM7TXTesBN25BCy4Ryf/ORz+ivjZZZcf96ZDIJLy/HCEUbXRvr
TZgHtn6vqUsRaYDWA8HLNL82Rx/Gq96WiXYYQq+d8F8oCCYWOuvzxIZYSgBLk57Omuq7nEZ+QJpi
qIJ4WZiKxy7/bZsyKG2HcaGw92ItTJGKvOhf6oVhMf//771Zev1404ONVcx4dSnj0FeAVZX54rnN
NJQbWq5ppkfKxyA1q5PzIxsAZAMlsnjcU6bYAioEYMXwTYlonC4qrvzCHRo0K5ZEL4tkSGG96OZC
11dvzqwjVzjW+ssvCNYt4PWA3XtVczVwV+F0u8I0E7RC2jq9SxE/mZeoVG6Qoyb6M21jcevlwAHC
VFw0SQT+nP4ISpBWOk0n5/HHkJk0Bq6yJR5qURx/GJNWOYUZDNIRfUREpaqZjpV/AlYfwnuJy28n
1KWOyEH8BVq9stY1XbtI4awg3Kw9glhR4wzQm9rmNluq7AgEmluaov6hx7rEqrvuIINaFGNpXsCS
kVbs+au0D31nNugz/1qXRNRxt1W1pehFmD39rHb2PcGIm9Esnt6xIc68DmR3Fp2v7EJmKRvfK7g9
dXiax5X97Sf3MbdxS+Xde2PVDiyl+9VOa1c1BHoFVIZEc/2dTshJ8Vcp6jCwJC2nbzRib9pE7LKR
sqOv/gxi80jjpcBwJA2MIAsa78J8QNkvo+5knqDzeoXlF0Cxttc/L0NB5m39gs4sPmz+I+MFj5jg
86OE0tmwL6GtdwuL1IGzd66/WSRYHzaMnaHstc3pYXP3YMW//oguEpJRQIXmilruVI6+MtEP5+W+
Epctc99t7Tf4bGlummPpHuc3gp3SOn081RpSAOqVzTeyYTXBUdpGObTdl2FUlg/m4MswZ3t2dPK7
X0VPs3dlvHtQWmS4y8KWoVjK2/mwgFp+4sQGEljq/fCKCtvN6giMQmiHkUL6mhlDnpkEdozRqzXe
eUGu1ES5xfU2FHc61KD2p7zj06vNuoAigt+o+BJ25+chnWVcKd9Pk0DFDA+Rl6S+XNy5YUHeBJmh
7+4+EZZ0xj7c9ItjxOZ9R4xSiwui//28QIzamRf9PmBy2iNQ4RMkDD5cf5NsArIinFF1eZ0ewTxE
GGTTWOhBTHYY8T+ax912MGvPooIPZWcrcoCpCWnrRGQjXZixc8+mRAelfxSdsk5wwy7fLbXjlQnz
DMzFlpGCoIJtnB+OiOl4ibX7P9Ak2+SVL50+1MMl4L+4bZ/SPa3Mlk1FH79iPF5rClq47BYyltPh
WMrXHHWqH8Y9Av2bABe8iDVJ6h/ZJQ3foQvH3S2dN8rs7YbVmknPjLcykyYViwgyYzCqGcWXiF9/
Le4hEOdz3xmcd1fAQIlPHUjngEBkPv9LvNzHlA1DQb0ho4Zugz7fsEb2yp8ydGKyuJRmHMgvm5LD
7L41OCnWwJjpDn+JOlnEYHAd/5g7sOpO/Gx7Ldc5S40tv5Ap63xlSRL/a9XDRVptw+bWnfZ8JMtk
ZJCeH/QVTNaF+5M60frQtY3Isl/k5VUeb4tRbXZb+MTvED5oXR9ny+j7voAl7PFXaiTXmE0IzhaR
BJbY7k2jHetoE1KzfLpEHPiJ8jTpgIOwZfX5ILtbrDkzd8T1wMAl1kS4adGSsKEABn6qIhB4d6dn
a/ESElK/ZVTMwtYSds76xguWgFQfWAWnVrthJTtsGSyV3AchhiV8h8/56vPuzoUKME5VXtsOVcIg
JDCjMULl5lSflhCif7gkdRG6wxfvF6G1RRFyZEqypLkIPxM+9gyljmK1xKcW0aWNq0OyD/nD70JK
Ld55aJ9sA+piKbrNQ5v8Fq8ztFRdWoe2w8ZIEUU3Xwijgl4tO+nmyddRVacFwzUtpBYU+CkMpVY+
XdoID/uH3xjqPAk7LMd+oPmiR29PB59Mlb5v8ITrMDC9GwFQMMe/vdqeCk1xlBsAava+lWCuBwJX
786mtMtdSQK9XY26BOTWgNvs0FHjkH4JvLXwt6rQh0sukK0qCfmF9Wm/0HGtsGTUbqWetad2NBWN
CNtPiJuZOZKhQWGc0ydn3IO9S36aHwoJuuacDF8pjVVxZv0oFuy1LqKP0StE5S7zcsQJJE0ML4O7
K0PY73wqRMV8jmI7bm4xAAWBAFZBGSO4OJf2oXHSIQSg4NMAP55qsWaUvphrEXHXbryvKDhEDGJb
EibY/cvYkapPo+8m2+klnxJ8H009Pf35sG7JhRClOfPnaDIwj37uSHzUcVzgcczcEkAGNxChE/S/
UYAD5+TdPaqyElawl7QopucYfi7k0vsJ9MBftZ2bxHEJPqhOCd5135nNEIqQxR1ab0GnYs3j5QSJ
7yil+mqHZqBoCFp+j+q0X5LV9lTHv1FDOPaxTNZUpsyC8fuEZtZZ4vi9Z6kTJ8oD5EIVoJ4cu4XF
L4EjLVoI0sslVlJY21a88wDil2s2SVkL/mqv0bYE2tWYk21cjxxfY5VRH+WwIVI0TEkW9DqIAW3H
jEhIpSzkjpl5KoyqJ8CBt5mQk580x0WNwxRg1lX20S5DKbyPc3bljSMMeNrrOfDR6boJtjvhIMYo
xWTmkMdiXUUqSaHIK5lJIxYaUt7u0sGypyE1d6bjZRHHwP9w+zrlEsfWxPynWrxMLuRdNk/Jc+42
n78kjr/WvZzuP7MjTCeK8YJZe6DcbeMmbFU+uivJyDf71xaN5YzZSiWNHdlzOXkxx/kGZA7WlqIL
wJ/3ufORYwU9V87F4PzPeG6D8HTfuNd+klqnlrl51LZdoP/aGh73hzMF/hw8/FC7lMDB6AIg5cvE
oelVYih6K1I/6YOq1SwsD40Q694TSvTTwNywnjpBlLZctXNwEB5duNmUUtYeyTp/bGLO2ST4yJCc
kpP5FefHEUXHAYgODb/GFHRQXi8Y+9NCKEXGJYjARHU4kERdNPDkAMi40lRCX1rgd1Bl+TsxJTnb
unOXACJvi3iZjC/C+6E4viZJnub5NgE0RHq09Q4GrdEG6M7ipEcwslJE/dcVTxMR1wJSnvjV0xQr
x98unkfsQKf8nv6g5yqTUc++yx0BTFIXmuO2zL2ZhnzAI9bY+jrlDo44kQJ6minhXEDxPktQc5Tf
xQg5ws7QjDKQ9TO4AaRbkK6DVayNgZ60DGR5uIO7yEPl9YlOsq66LFu/NpTIFctTAo7PExxrxM6A
uBX+0N3PSeHxeuHcNsNhhAbl5SPrUfhVVMMcBoa8Ka7vW2fpDp962VCuECiRXYCNOVzaf1e0ssy2
ehnj4yrK8OR1RkzOXEWZ/GyhLe7sK5MitFY2H2PJWnB+mwn8DcyP6EpAv7nw3k7iWsWSH0jJYTig
QDOe9W8TNd8guodjC0i4CqjPmrd2KoemzQoD6mf7MF0L404gY0q9Fbel2vaBdRLMTafDjanSn4mU
xNepMtWq2r51gNfO5AkY5e23aOmevXakOZzbNzmlEakIvwhmEP+fri/RK3f9VDBOZpbd6/ZYsN2x
7b7zqkkCKLUgXaXczlxHk0dWm9App/wcprc6U3pZz+p+7+0m91MWwWZpIai8Sf2zOEvGtQUNUd8j
6k8TmAXOlab2oWkETk2p91a6vXXkkMUvWDtRlSIeKRtS0Q/U1QsDuxdUWIWsPuL49MRJ54FIqPTI
w6qnNfPsRUfl9mc2SrYq+0Wi9ameUhKPjhXPDcY8bwuPo1nodojyYZsDmmVMVtstYhLji9RQJ3zd
pAZiZ8eo8zL2fM24ZT9dgiTD6v4wxDyJfkFkqsQspc3oD6rz3F09c0XLUj4F1+4WtwasvlhWaS5O
MyxxneCQLMQFfsMz4ksXb6SxSs3o4JEsSgH8jNq9ubT6o3L0qv3Tte3AqZJxqROxSSK4Ojxmdzzn
U2ORaiyGith0qS9nGb70duXNmvrOcCR8/kJlhvR55ZD1QmUIOU/K6VIO0hQScoH/99LbrRpmg5E+
xMw+Gqu0BS32PJ2LV2OmJx6r2KVvj/QfI0SBhEojIvclHzpF7X1Lnz3AnSSFUoCJdmiDE4OlwRoO
k1rECvPs3XT62RA9+cXvPexF7lfktzCMUyyfzIzyzf4q1S/S1fiI4+zMfqRRKy3LkC+9B4aEQ79M
Y6JtFwiZMAbe5Vq8ommyn0GpMNwG8aHH2zlaux3zsPbCXcZ76MZx8/g7AUUqzGgnZEtFyRdtqHVA
7lEsL0hI8BxJs9oXbv2fWs3V8EZ7DaU/NTFm4U1o0li6qaDoqeMEGG+CAcQ9GepkN1rXKHSxynto
BrLuTZ2I4fM5gprjmq/OlTPR68uYOVvtCRHhg/obtXrryiuCfuQV2uSz8YRWYwG+SOD35YD84FfY
XEe8jItvMbw0sfinM28WIaJW7zApc+dwMl1qY4gSUtuF0yx37Z5vOhGUNpEge4d+NCTZnUfM4sqS
EYndP7kQPQTMUddn+Cw0GnApkqacmzOa4wdUqPDN177LBPyFK7HO7ygm82VCN+pHhYuqfo1QrFUt
mwI58zIz3Yy9x1JtpdHMIWMYKdtpPwZj7X/xMPt3AGDCiUO9AH5U0YBQuyhvMt8NUooXvI+tDgok
NYm7UcgDxgQQpxBYZM1zi9DO3IhwCJBZyOJ8aUsS0dcZa/Ec43Wc4UiE6DEC8VMGX5eOzvgfziTP
65aCjxxev6VU+sZt952UkxvEpKfGA6I2w8yAidZZ6dinyXjQIG3QuEiSu13zXSHlccYbV/CMm/W9
6QriE0f4A3raUKgdRZ8ruZ99Fpiiui2QREeDGClBarwACd2IShigDsgeEwBZfrZRuXf0DUFKa5Hc
uT2X3Qg/JRxFH+xm45QRYjbvQ9NrRrkY1OqrK8b60y2wTbxmE1kOnk6RJ13eLH8EZyx1oPOBs/YV
xQ8ELw2ZzNQ4v20zrKyBK0p9z7rHJ5JDWJe8G1APV1u8+MzCBoq60gaAyNHxlW977meCOq5hGlyO
VFr80W5B2h4jp0GAhQytm/anl7hppzQTWRQv2ir+YR2uObkIm/x7VIYva/bQEtTd35/0u607JmJg
75ed26pIalSJRmmbmZGrbd5h87XETW8MkaKDKbfbW3yQkMYBqbjGSW3LUKqsnAo/IPl5G1eqRTxg
/6TWEEHPelGzQMKPcPMUxnFNIUL0P1ALx1qd0H3EOSDT+fqTpZGgUJFvcVsiE4mbSLqL/ApEhIqi
FGh4glu1QZFDTP4PfiiqZztTucwgB7hZQ6vdJNA/g+LgWgB5uLORAudVmyffxvu1qzAF0tw+vnsD
vyIU/Y96rPOovEtbmDjGleaJw2KGJmQmIs2q3x/t0WaFm1bF6mdm6gNtBeyRqPjy4bAguQWLm6iF
GXEMoqJ+N75SRDGfoM3mEtanrTcKsntA7JcKlN0pxbKkVnzrrdg84FHZK/eP654afus8ZTJ5hxBi
pXpfcOTsFKm7HMr2hXUdoNwyUwFrgrFrqGgicDzoBYfctO5/eaDplqwuDYPhdxQov2a5xUQay5MT
4GyHPGr7CoRhfI4swNmwO9BK8tWt2F09jNyujw9WlQe4VlktY7p6MwhBrTUH9x1oLbjg9zbH5IlK
ALzqNl18p3CxsNxCkR01mXH4WNSdPxtiU8n//ESHDliy6Jmwhdh52X+iC2grj1sIBx6kBF2VsWRi
hDKXVAjIeDk3DNWXaY1zdpBNracl07qIahDtFS0NEpqu5OhZtztayTIOxrRKvG/FC3eFUYR2WlN3
9GKMUN/rp1Nxw8HmdfKqzwbXVQd05rnvABVAlu/Vky3al3T2A7s9rQpG73YDSz6lrfNmZgOCMCMI
HiKWFr/ydWTXDVFz2AGKRr1N4UVqWjKK7o23hZetDYcrEz8A2Xo9E859XIK1tMWGrPEso7Vn2pZb
rLLn8vkQFqliGfjtKjsvC0OJHozmlAzHbiPPNgqagbAikavrQTHRDVklcwYrvsfUucSICgoPQ4kq
7Qn3jlZusJOCO2arhdeETzWb2MGx3hqYpi8J/ciLXou1Avwms+g8xp2bbsEiKUk6ThaBsq6ZnB9E
JXcxp2q2oE2uD330C/Ured2+JlvmhsNKwYiCTzAeOvefNkqgPtvWL8z7gWanNQ/ytbEhQEantuJo
eZeTnjkgnhRyeHf17mibQmbvIgabbFDc+J2pkjq2yjZq32P4+DD6XHsbYw6Kz9HZUT31uH0CSa9r
Hg6+iCi1bS1MCkBsHVpVMmg9XPTzYHfIZy3nYA8N4Y4dOC+wU26/Ckhsj2IjKzW4s1mN0as1tLzD
5RlPVfKy7dP/9xp7BFOuJQZF2OcbiJq3Kkekojts3ESFOzO6FcmcCBvahr5k1zGlDNxVOk5zPORq
5V6MzD2btzEZygcNX/LFRDWZJZoDtOXDg7urXVTL98+ASfA10h5OTcdLD0oG9hwzws9nPN3oOB2C
Y1WHAtiys0jtq3Frw3c/D9LdGZwVsBnOyA0OaVAE3dHziYD8rXp5Z0Jr1fDKTqJyq310VYu1rnq9
Y1JpusHtUbU2QSq4E5tsUceUBU3xTVBjp+ry9kABGkjaGW5gnWucU/ktoLDST76Jo1SQHIImZIhb
LeV8s6kWk9qDdcHmdDq/jn/0u05Yl7OHs0YSQ+wocweQXpq5mp1h98aCZQORwUW88CRQMSiw1HQv
WqH8T26DB86iBSN+1j7YPRdQoijRlznNAY+ApdlFgwKQAcDH9LuipeiDPeVn3i3tDUKHTs3nKeBZ
CnS8QxCXJrFaXxXWaTXY/qziFrCixfQe20ql2Yfeu4sYhtwMIjUbYanVWGdHbbXrKNUZpJDYOLkD
nbXSvRA5OAwTZLcl/3/BMcApfKnFzGt+4/SjO8mP7qQROU/IO+7rTfsDdqxcHrfYlUwg4bFWJxjq
oq4VO5XcHne8sbXCWjtZJpRgVexked+3NWwQIx7nLhJn0DHsYOiKe9cI+BIr8uTLdrPWziIQ+Iof
gjwvuL9x4oXWDxbmOcvHgyvbUocjtdE9R942N6ny04pXL4038LL/1vTgLMMdafIktMgXSTzMjFwZ
9TgyW5+SUB0swoRYHdDrGUCiK5CyP3WlrKSVxUNuCCzDU1vQtfBX9AuWmInF1j2Y99par2D659Rw
ryfTE80zn7KTbPTKq92g2H2PqYnK+euLFh/WiUjFE9dwreNOeFCW7CZe8Q+ZnbJvhdhTnZUXL/3B
YCnLBAHqi/kYBTF3PuY7XIZCGkghSYCAwYcIrKf4jlqrLm9hG2uYVNFFLuRkTwbstDp5E2jExMzd
wi2c+Wiibz7JHdmEU59/O6Oqq8cHy5HXguy25mgOFGLq8rV7EHgESG82s5bqop5zDSIJCb5d7Bu8
ZByumNf2LaaOC/siWQpFAC3/czXSEmNtwki2xI+XHSjlehl2kytX0K9ka+SmtBfKr51rbnUcSCK4
Fvz3m4gOJGTTgLi4EfBQuCCFg2EhlVchDaTyd3J7SdO08Ggmp/i+WpDVAZTTO524wCyDvzUFW7Z0
GvmmDqEoCPQBt1hz1y+MHySazIk400DCJ+P/pIA2lIrh86Nc1sWHpFzKqgAVEqYbfqYfgtAeQdfm
ZjyfCboRBLb/Fz7JeOGBHhWOZlI+WdAbdBVMdYEo+qBBMnHoHAcvAEbbo/1DrrRjbWvT29APkJmS
eyfwQCLmW7/+fc+oSstIHrhYzWo6x62YCOY7shrT8RNTq/LHNmxsIyr8MhbOUz4ZAxienv8zk2aU
leOu/l/urc0+8aMw/IhbvpimGuEcIacLwBnkwHaPKOtIQIbgegAoYGTzgy/nOgc9OorcEEC5naCW
DQ5PSW2xF9FY/Vwa4YE2caKC7Ym8K84LGF66Y95/YhohM3IVvBQXatsLU2pIV3H2Es1tj7qhVIBZ
shV+1W8d74ORV5F8vDYELM5VhUqNeeBRIf+Qi1Y3+PpdyWp8CLFCgirDIwPuW2cnMoxdpq209P4y
QS5SzELOe5m7BAwwaLuUocVWYf/bwdDkxSwLYeYfngxZZyXWlJgzsoVKosXSH8k3M2rC2i/TMsY6
qEv2gX2Iz+ZAB9IHHpM8ul436ZDb9tQ3f0C6RCDkt8dHDoEQzcga5P3O5RNy8zbcdvIVVbett6+n
SssgYhRP5D/hGUyKT8qoUjX45p4fjYF0eoOMPPaXdJ5euK5wuRkwz93aVVfs8g6OJVe5vzpEwL6J
TW0j/LyBViQWhcXODJ2tjEwnqvNjI0pIMhOLrY0LILP3i//DP+kbiwCouNeZtLtiDGZvKJpuIPV8
nt7KSZv5G1LV+JkyBTy9XuLPh1UO8VSfiYQfxjpLk7yuKmI9TBVc8zhlgE76BKWHsbOgBEanjQWh
TM8pz2Koe3ni3urCWo/43UscX8373FXhhdhbjinThriWv33h4+uycAbo7nHUq/mRTYXR5hX2vl4h
5JQg2tO19fHnoIw/PAHkPRw0LpOUXyLkBQWAi4iOsdvgPkr1Lv8cjjGxAph6vUT6LuymBuMgi7hg
LTZzWJhJEcC84qITjyq/k2LigeMp3WF0YNBlxBP8bSVs6sTpcuoPlCUghlWjv4ozPiH74VfPA69o
gJ2GFzHy1mjxlvjfzCG+8lzycP8Byy5dhIRtzA7wiVNBWuL9unREgHGaAVVgS51mNNAasBkV5Vck
8YDaJTywi/lj3vJZ/pWAKRK2o6izQrDg6kFi7Afxqq3U0kaFzpRUUGm18z9UjxIIPpYROyukBsCT
RyJ2IfVrsVIqavob8s6g8gXL1Aee/WSpUCCbey/Suk9zNlKPREXLG3fuc5FVbJKXq9arFeFX33tR
ilS1rDzSul5zXd5hYViVK4wYDD4Q2n5UJf8hX0WNYM5ff3AGr/B3dt5Llr3EBILTtlpZ2OGoXizG
gq1jjInqxY8XjxyMpo7+bOma+gOJxtSbjFaAuGRkAFqh28HqffOYPO7/sP/m/5QF1e8jrwX/laV/
FqMyF6wthZ3EfBadavlkS7z4FQiV2L2xvEScc9uF2xbDKnwTSSlxQQsssMKYpUEa0Qpnbn1Mp3y4
dK2fw/GyldeYlgQqvoMdWvDJuLJzSy69PC/CVQORU6pm4i3f80n283kQWrncG8T76Nan+y9uBvvL
c4gRmX8tzngmLRJNZPNCOdqYmVTDzE/k3C3MlSQ4NKoqR++LbRrt2TfxbY5dkgX+UKJ5pY2T3zjE
7GffQ4o3UGongKe8UwkC1ERQtQDG6839lXiZlbN5zUkh0rz3e0RYHxJuOarancG6fRIdnBhP8IsJ
xlgjGd8Uxala8OnPtJVFwAfYQVQ7jBLLDZj0M3d3Fn+Lot4Hj5m1PRxHjRDBiXBwFioLL4StGZzg
r0EnKz4C2KdW78k7FA63zdfcnHuDsTGdYNB7xXCDVL83wpIb9WGdCf2qI7yA7JhD2u431wIo4WKW
i0Xewu47OZDj01ZYDJNMQ/xM4QwQsR6v7HFdv+3rlgg292rj0fyc0kvsBslsWitduVwRcd2QOAoz
I0va82S+KRIB1/2oV2xR2kJzrN27WPPrBcFepu0aGhcyCLFl/k1OX4JPkFOSoxbaxCB7okX+JG4j
9FErckoqAgNHJFiE8DD/Uu5sITv3XFHvS0MeQA7eE7jUA09cLfEgVt9ToxGt6h4HjEimtrhZN9ha
IcoZldml5nOBJMANtwvNoCr34kPXo8jEOguG/TU8CgXDmUozJk5VJnUnbYB6I/CnqM56l+XUzpFh
UPx5W1ktUv68Cv8rBk/NN6FR1qFCpU5og2hTydsWFhjKKJUEQyEHvONa5zKKTGyLrIGbkYN9zhuJ
kBMD0Nk46tnQYaKMM1IrBwWEzVshFFENhUBBNWywEY8fdzfaRNWj0k8dFJAva3NV+Awo/+j4KHxX
jpdM0B3+H9AZchxS/7sLrxga7kj+yLzqQhBS91dmWrktX3oS2EGyAvWKnmv/rbl/myZv9D7/gE8X
QuX8ZoT19+YNyK2lvYkNoCHjgZL1DOGVAsfyV2YEuwQBuvOkJ2bweXFWCTHi1suBaxJBg0W3BHAz
zxmVwko9betbi8axnBOV4ZuVUXgGZ/9t+blStKhZ0V2jrAu/3awhHjboo5z355dUl2Xx63WqPyud
WC4k5jRx3L2NU3fdiXJaIPxXy+A5CtegA8efaci1GJfZjenJycK7ZGYg/I7ECrO5mxZ/hkklrxv9
xkUmXfAm565UR/kO6q5sk5w+HOFsRyinytbQPPkdTHwFIcKoqr0melWIovBDkgGSgQsJm2BvW8ja
cd5BJbBYDbKctQbXLH0Y/tZNu+R3qF34YKCHKGK/TXvlIeigGryn2nC8vcQHtp5G0D3PYk9EOXjC
W/g2QInpBpVdJxN8kUhKzcKYh7+UNKDErakzfPfd75BD4yhOELh4TIED1SkHAAKzSzKeiVRwcmMj
cx3RTJIM5ut1qp0afxZ4svzcS/GQiTfwm8T4YcxQYQg5YBOh6tncQr32mH41bblcJRs2W5t9ZKiJ
SR70bxX+oYlUxJBlJfFvwTgaYJ3W4bpSa+lvipx8A2jcR3eUyOyZ+x+ejuhGvw/0otVuycITuBDc
KF8TsfiUNCAkcBazuWagTAVIt+DKlEcQF5aNdllzdT0QdkJCDelrJ3NBEGzX9MKzaHBDkOs53zz3
yESiLlHrKjveJGziVeGsWLGz/iz9JMChmmf4+yY++Hcp8l7IZUrQRiRFokEDnGrto8zhPEjneUTh
EbO0tvXo/cKB9dI6P+QzYh+Dz8wLmLPca+u9CnpQo+1iOQtV5EzeN2EzlEsJeDM0tOOohJCnZjC0
E78dFngR+4gCxyxTOmCboENCO11TZqsa52Z7twW4W06sdaKLD6O4iFUQ72F2o+E6f/8cYyNpePo0
YRzbMW2Az3xqw/rKyspqqgINcf5T/nBbhStjLr1zOzXUJiYdqDJFz0umVkObVTYiGJNf1jCE4vHP
9q03WXxju4ZB5gSsaspK7LuLsD0hqYwCngWPTOIARd1mVw+7npn2/V5cLZA9kKI1uCw+pjr/AtEm
Ey4jnBHYkoLFJ36hCQmDFiAwqQPOQ1A9TjGk3auA2oIQ0zOt+0OjukbJ1SBP1a7jcBdqIGnfLO5d
/qBXkc5mUXoZ8qHYpSWUdv8gfJx9ajrmSYgC4lLVZ7eEQVKO1aEDexn6wFLGwE6w6YQBs0RYmmzj
sAlQtVT8pXPSkgx//QOh+CNOhs/NB5QsI8JkNytk9ClVHoXpRnY09BJ8Mpf5WL3y4SKOmqq9uVge
SaXnCBesjg9yuZOFnc9gquwUXZkc38P7Xo/9bOkDZlpIJyUoK630ri4io1mxiNXcfV0/ydqoKWDu
GpzQupw6md15FkRd2s8hfG5ZhwOYju8tJ4gTzcIMDAK6Pi8w5Ca1QSZNxM3bMum6UpHv1FAajeqZ
PP5UU35+mfsayEd9GPla0aIa+z9O2KAMvSBKakpS4WicY09BSXySZ1J4Rau2J4PZQw3241zC/5bv
78ay+h6ltlSVTB3L0iY8knJWoe5fZILEbrgYRgfi2vRgTL52CqjffTLN9u+qJrkg6D+qqwS7s5XC
TG+iMCJB+gxfWhgiN7pU9q9to4GzQxHrugvxRhtQVoQzlImEkR11lgAfre/Xy8evdfsigv4CovFv
oiyaOZ3+nzr6EhJi6SsQcY9JaZRzn1W8CcY5pvHnV5n5AbL8r1F505C+56CYf3U801pHt9QJbSFf
e/gkZSIF2mfBdOtwF29S+Z/ar8WkGUfWHVk7h2wbZ1CAvDc8mxFKz+5O8oLS4YApxWFgfg6o1+8Z
N0J54Vh1/NL4+1n+zcgcXf0+DG8FIJOgSA8eUoa/GSZquJKsQ0Jgkb0DhE5ewEnIeGKWuRIYXPSl
sb1fz1/iP5DlK7n19IA4Q62oVhuO+KgWJkBj1zYFiZECkaFSImERVOVhbUFTom93MBCg1x3SLcJM
DWkJZQ/okMFD29pGdWFc+8zFpBoGm2nxJmyOUfmtEJLDQJoG5hJ3kVTKkYO5HcCjWBJkAlBvYwAj
dNDrF8dvycM10xM8z3YJYwIDjmRvyRKO7NIwxsPY/acZru3lr39y8IqbOmylOQsZ+BMTdtDpfDPd
aepMYErCqsRThFimHMgfmNUj1k/lg6voaItomYsgKivblonglrz2HqzKd4NFfQowjEw6V3riBy64
mm35PZ2uuazOKaCGR+xV02j9pLIIx5oSo8dCDjSx1QIM07518P5kW2E+tNEdS1lYrJBowa+r7ISO
m4X3lpF8UGpDWRPog8pq/7UIk+MfC+P+dSVMBcOcjjnAuzUA5zl/LYozSTsmPmv0H3RIAQkHhwtT
OTbagM2siD2YBIHPc/UoaOO0UOnoqF6V7KrwnYgc7L4XIrkj/TXcSLH7rKjgpDo25InkxDOLPFD+
2vk7ahgjOoiPutJJADcHN/hiL9NsLAN06EKn920NumdN4D+e/Ppz9q/mRCgGoxUWomzRpYZtxUy9
DjhxQzXKYGdMUexBXH+hbZ8kSS2NLT1yseYnJId4+vBuQNzgpP9kNyLrPQ067XKdPCipnLvuXKlf
HbQvlU12ZF2zhDrtmd9U6e9i/jx2TWn0fNa7A/gozHXBBC7QT9oKA1XzLJRwRjNC4u8TwDiHtaJb
g3L6BjRTTNT2Og2kJ2U/ZSkt4pqlSyRzIc/WoW3e4vhOJqlkd12dV7x9mjymCEpHRxO0qx6QTGmb
eHBwiNA77APDsWWXzUMECfDea7HjMj2NX1/VCJIs371jOiQtY+QKbLOZEHM7029ko4khnMQ21D/n
vzjlIUMciLakBc/bFjzaGlGw6/7a4wfvyz9Tgou6hPjYLqJYTkMgk8d4bU8bNv5RfQsRTESBTofP
jfbm4q4CJpfNYz0BpXuxGdPGjQ8Mk4ONeIj6H5cxsZsTtGtv8IVi4nhCLBwkdfS+DRgG77DMkddy
GwiO28Sxe9TvspeA0mHtf6wuDziVjGwnYB2njDJ19fxgrloczYun6TduQDxKs4Onk6RVOkLLLs8C
Wx3CCuvq1mWLExJ0/8pNI1Og1lf08N663f8aCausyfuHSn0tyCLO4ETnhpXHQWJlEzz8y7oacWVh
Fazb4R57MUI3vDJ8fg4OeidOWDp3TlniGOeusBzGQD/6tCvfAgWIJprHMYS2Id4V5/pevd9E3DLK
xqsxmSs1fUJ6w6OCJzXERWY5TsJXnPgFkZhNU73E5kwiwW3v/umv368bbEEbpuzg5jFGVqspINY0
ngMSv5SxMnAJ1EuDIsOnbrfVUxp3nic5+p+ezBJTeJ8T6VgIP8HRM2JQNMBXKgC0po5kD4gl2cTy
W4l96ZGCBxfJF0cnaT7wHXt98IVE9mtsRwlRmTLRixPV3ahKLhu5yVIX/GPC9/Zao7PMNXvTxNBt
O2YAcfZzLYPlJoF5C3dYa2bz7gCD1nPN0nroR1HQwx9D1r1/Gns59R7tL+CuC+Hw6thdU4iGwE6J
AeKzngJUCjKz46pISdA+9JbORa/aTG4NGnEImRbJEA9XZjjrOfk1jnVYs6VnLcFYck515PaSt3k/
MuDgLWSPnWXtHMMNt9y/BFx3KUC5+9hd5AAWnxGqdpeh3LvJPGKdCGFHz2MiVpLfIhhVDmz//1qg
ue+f2z8ZRkYNt81i98nJE56J4oskpooBtdBMxbAD2FNO10LLP6X3X7SUyWjQi4doWWTFaJX3fNSa
o32gnyZW3eKpfu2AqKFGTK1JdFB/ljwV0ecJCOA57SM6DqaSe2jSc5qW6xgdn7KDfuCkk/NSrGnp
MFUYQ6a87cwB22hnr8lPdNjdWr8r+YyIDC7BlLiAZ+LTbaLnDcMN09WH5zhdiqieqmZcOvJyLwTj
ZAyYYLV/DrRC7Y42pbb/r2ojl3Rz195qg9glyUnK58N46SKqyGOwhtxthaaD4XoN5XMcVd65vjdx
uS5rN9dDPLJOxXJcGiojJ4ChryK1ixk9CgrcM/w/tTVdFfqVzDQH5UaS9rDwsAwDFfIgcx+Uurwb
OjRXu2YYT+gVY/imz+OtXZB3rg1m23gpTAE4rMvxVIOyfCVeMczOJokNA7mYdN6CxPJwDgnzJHE6
n4DFOqAaLdxJh8aNBLlXk145WgaxDzKfN3DxDKPd928dR/qG8zxAZBvIE+ZxfaorMcZGKAuw8WvA
OPmPqE1kfm6BrYJCqef0lmGEaGm46vDBa8n2xBK+MFx3Anq9YMTC7Dd9vkXHkECpBNquwZduKBCE
AwNAiEpX9oQE8cI5+Ry8rWquq59oC4XGkIRii9XLgYkmLKdwS60t15yAI8EX8L7Tcy5+OjmQiSrJ
dvRNjprTc5T2VFzcVULdYWbh8T6Hj8u/IrI1cvVXI4HfilXedf+iEe2S1CCkOgiefRjO9K0LH1jz
4pHbh7br/zpnaSuXatVldT4NM56Y7S6wYC+G50t9sCKK/83OFTy53a1n9mY80QDWK21Vx5P2129F
FzlpN8IEs+irMbUOBu0w7dtrI0s1r7weciz9QoPjefyTl45p7l2D6xYsCMqtHH/xrtRdXbkh9Z3q
NJTTpgAF/becEd17sGCpw3R35B7tJCHkAciwiAH9xBknusIl1RN0ABBI1LaglgN4CJOpG4PkIRxb
m/DyicxNB21T0pHcZApJEvLktBX2SI5dSHIqTo0sa3IUoYp+dmEKIIRFaOEuDiEGFgAs10X7XmIn
l04USQwEYUKJKzEK1KP1f6iAIaJNEE4zBnUKaY/PvSBgDpqtBD4loRzsXzWzymsJCM2vUgksSy5F
N/pjPrUYQSqbRT66ygqmQBa/jPsU39wpFnW63tWz/DKFTpwAfRoIv/0XMBpa/cFhyku18FcUuAY+
pR3afsAk9RrZuxZdu+gxOjZYP/okVR4KubvMmdqhQ1MwohSgXV2Xx4AX0vQO3b1uNNpS5WyU+Slw
YSIUeoz7rzJgkM9RRo8wCnyP79lYNz/nAfEh6+PLjZOGf8Pl8AYGMxRgXMAQj2MQvaBvilfXZVFu
lC/US/rU1yvF6bSVqf3ILo2OY10fAZDSmZa3KfbumxzOc26KHJCrlpzzMNtIbxDfz8p3AhgkJgGF
PBAoNcXsn5rJEOXowVWS5Cjj10BEw0/y6+20KhH4FG6Wdrr3gfaj0jytw2/unYZrL2Dcw1Iq36Kz
0EdVQBBPnMq52a/JArZpo7ONHta806iQpf5LuDLeYEEPu7QIZUXBfZkqIlFnky2XzgSRC4GB5/eH
pAyAPwv7UG2qM8z+IbGVLHVvJexzqgOc6ZUQpHh1RETOnpjcDGMZHXgNHZd6baKd8hmkW3y6lguj
7TLWFMjjrZIH+lGSpcNb9BiIvubP9uuX6s3Cg0Qu5g3RUfciK1jJTOJn9u7hAKN6n1g5WoWWirlV
K1/QxY2eJfcFnRpRsIvxzNZoJkSR+0Jh//tufFCjyqrF0nBY26haONIrxQcM5SwJY9KWJ8fiGDd9
6MBeFoIwGrqY9D2wRyyJRS8gV9HoGAElvL6rfG9thc5I9Ao2ruCLp86Ad2g7pFDDmUpO5j3118cU
xvV9OJG5GEFj/Uhq4ME0S+c9mQGysBjyTMtBEfn+RibRUOwK7u0KPxhFJAhN7x57anAp/Ay1U8q6
DELqEZPPIb8Oo9a4nS/kN5BLLOzs8OarZKwAQFUsqCeJedoPYk/sDBsKJwvJHH7ZGk/OgJVbxlZ6
TEHvFviH1AivvUHxTKruXDaa0jlQxkSxCXD6P8W1dLKIXJ5hZ0K3evfim2uf8q71e6utl9o4ppSa
STP1E5gl1RThjoVhcPp64VpT5gejmOr8MD33k/EYQ4wyTUyM+lAA8IFk0RlYl3w00EJkoGO75aNJ
pQ1pBSQ/gBRk0MWVzDbgMJRW8Z5e45TJmwAHfTF3dpCzdKBWfCEcTlf13ODMGZm9ypzvZV6muLLG
94SXhWoTtZVkBzp/0FktBaxOg7OQ/gdPd/gzahskSkl0IXgN5JbxSh5Ug43+7LgmN2kX0hW4Jv9n
Gh4kx4qDqEsngfriDYLMb6ky+Cd8zHThadbvSp146aIohZy1hYxm+n8chUrXDVIPEUwYFhEeknjL
XTk+07wBtI5Wu5I1TT3cq5LiHoGIy/RV1obFpsvPVGGjTePMo8JMSu89DvDslNYfOq2onPV4ntcx
DEQporm0fg/+LenRkarh3FcbD/GgXRLZrXFzFj/f2Clp61T1ehijxyXGfyWKGGgulmwRi5sEnrMm
u5VpaMTpSdpOJoioH/NoHiT2FYQw+uE40LFVLvnqbQunZqzbHaEPBwr3mBoJ+sK7cjuq5YlvuAeX
ClJWtrLnyV7/cF3/ABJkNqu/4xdNBragrl3JwPQYQDKMjzTEeTkbTjavJdx+hrsUNQx9nZaKiy4v
VPMfQnzhn31gRwCHlwc7BZuQtnANgyqraARncLxuIpxRnC5Rho7dtjYMr/ryCIbF+tP7rInjgIbm
xGWtzLAOeOtLZVWgBOd5PnybXruOewI9nU1RWpxWQkzK9f+n3TaN6EbCby/ZNeFy74CttDqhdcon
M2sPM/VpOJ4HKsZLg9cThHkxuU0UVuE5qxXsoE/TWYWj4RwgJ75ev05HE6Si+jWFfCAz1fLvoUrx
5o44L0fSYsysyqc5kkqSVxZU/IEhP94icuFKtHJaqiKmQJdUo//GJQc6u5v9pM1prYarqwEf+Sbq
GGyCzDPO5zNRgtRTdAQBnm7i55OPGLkRTIUa7Jqw8vue4ATtLh26jBqdgXazbMivglogddP6v+Zs
G35Py0LpfSh/G+h9r9Vszf7SqTbDtmyiO7lH1wjVWr2T1IpEfCmpGqeNVacJVvupWHEwnq2K/yRy
IGgAFRdV+usJKx4dl87829IhbRfBX1nRvN3yYYE1ykaCYDMMibM4xFVBZbz4HL2ZbepmcYo4voFZ
7KUycmBn8cFDHKGvOB3mqImTyy4GFmsiMCpaB8OmyOI4sNj1HeQ2Ij5bxrHdNX0JIFRi0RKD66vF
QA33QXcOiB/AI/agxEwLs5XbL8N+S1BE8EDDgr9+OIuQTSKbtV+f4FH1CVE6eNI3+vfJlJm1+ifr
RM20eXmOOWbtMIA4tFGqI7xusqQCWuWqNHfYktRap/BnPUmLI4zMFpyby0yQf/lit45/EZMvKWro
fJm1g2l3rKIP1TBdKNpiOkI19qZ+kMc0p/5WG/gU6lA1fpKJNk78tppw2MyGCf3yi3+UQaB+Zr48
9SrZ/C/krDKVo+Mu2ZE2byLOok3j9nV+A1LBQSIC/KxuB+I765zcy+chL2lV3YfVWC1xjmtBxg1U
TFEWThcyAqu4Pf/Bs0bE9sKJx8Ed7k0b4QJWvYT1qjXXqsF9d4BXny/D6Ti0cN8lsHmX6KWsHm+m
KhCGqf+CvkZtdMFW9MWtvb4nRjwNGECy+qv/Pn0MZ9qC62lw1baHAWb1uq9z6qGsy5mA4AwUpRtI
mRLKKQ4A9zN/wwyeAYIH2puH4ZYHYUy2gcka2THEwPCdsSypWOAYb855kdcqdbsrboeNMb5CpeoA
VUnwo0/Feh3awSOVx5afPetUawSZC9NT2iHxY5b9dIpooqdL4PZZkJ+NTfN4Q5ecxf+Xe7oZ64ct
oSiHPizvucjn7VPto/hBG24BTtCQzCvtYSiS17bbYFVEGsFWNPvPTYyISVHkRRmFBzppnlcts+Tf
eIvbB9gmDiDfHeiGwLKhgLPNiNmGNXOgAZTLR8E2n7NzRHY0EsSOP5kNvSC4c9+VQLKO21AX5Ww7
OkC1SwYPvyj8/x/4Gb3bEvT8ySPNDJu8E8j/e7I5AGP5JU2jgODj31IJV33yGYvPyTPIKHAP6Fov
qGqwRrvs8rBW91BXUNog0bsUZg84ALwJasH0lLc50sxq0ZeKY1xNy5B2D6bzC71DscEKbvQObDCg
Z/O2yNuxHn7kZYzFeVm2cRpZp8FdwctV5jSVmJhzRckyzh9FmlVPTLik7RXt4wDDAQH/+Lg2522d
zwV6aHXXDd7ssisQBbL9Z5YIDNM4rl4AFcUS0ET7NTX1P7m3cnLc+p0DRpqhzYby+2kqjaA9Yq2e
sRPFBmWvFaY2I/C2SRkGsANzmFCREBY+mdW/5rZOnVlUIZ+6dsRlpRdDEcvsCG22Qzd1yV/BdE1s
YRRwxbACffjUmKNC8ATIg5ojoh9SepNp6o8d5tLbaa2LABTqBvI+cXGHa7j922kWw+RddEkRD3QF
Ly++y1E0f+PcpL1n5Qk0GiZpsm/6v2Z3kURRbGA3LJAF17+fXeotT2JsrMJ9dArFaRxT5Zid4/E1
L9w903gfdLtkulXyJ7GVLESi/AdC/s8eMzoZ8rfUV8mK3nzoHNA28ln6MdWk5Uh3W2DaWHxAlvSU
6ckGclTdTdAlCl9rPpEw7FFcYrGFVj2YOYIshVKVTYTmbQ48vI8/SkMDdjlKq4wAeUTwLjWKsxn9
TcsPcRRi2MoiUBgXCzamqPsr88TptDlmyQbXcOjP9A5Cr9jPUfFD3nbh3VC53t07F+ZxdgoO/myd
HmsluXAGeYJIlxMi1aLlQ0HMDmtCcZI4NNkHMDiIa+hFCyWVd7SASQ7zRj9L0BwAIOOePrzpn5Zp
VzxQLEXtZlmZW2/nx2bEkZqbWAxZKeFYU991TKBwhFFzImGdwZEtZOLGJiY7i6YonCr4OX3Z8Kxw
tIRqFC5Oqz45T5nmb3/09nIAcs+k0H6L2V3mGbF1JBsAr4T+XmEjXv+7ZTTKwnGq67nvBGOG+WDJ
Mc/Yu5z7Wpfd8xVubQ1S6iTmonVGocI7wI9Znv0j+pZ3tDxmrQzDH+ak7P+hUvgwj3l4JY7IFn8a
uN9nI64/atalB10z/iLDGF2LCpxHC5HM7pvSRQGlmVq95CzfKiL1EKqoNkjOpDkR5hCINlJaG9lu
3pxwf7zOd8MmJEBZJNU+af+uHK0ZBsF3Hylj5Vq3DXeaswcMxjs6K7NGrqAMIVZ5Qdf2sXjqAh7B
+/9Cj+a4wcYQzoozxVtZhEFxjetwk4Nbg9UBuBVnqZY6WkxBa6B48MM4fDBllPf10ee9oYbMxRvJ
WI1hd3RJcqHlWC6LgGo5Q02nDFaQg3fb8Mfp6Dy5hBYVodqKIip9IgrCMzHuF/TnEqZuqy2rcLhy
lYweoB8I0leq72OY6sPsANTqWRlG18n2E/mR5jYi1SU0M8723WRv/j52ineW9yR8pJXe11QO7WA5
TPMnr+lDwS722KNNfqMDw3nV0ceTHspxhY2fSrKkTbWL0uIVBK2V6FqHpB+rQV2/onG6txmcgBow
lH009FeEGe6oOoK8c/lUM9Yi645vkULgx6+U+v7Wnmqd8lqAPTJFAnvkKQ+d/puq95hkYxiyDfg3
0Mhii9W6H6hLAVD49ePxvaoXL66p194Y98co5RY9MXHn1nzVKZzUvQBkSNwHPGcUaHEj16bCrINw
1ifFfRCxQaaSDvkgsRM1Zogsm160x1Sm0q2iH5TEWiG8LPM4SjkO1cDROFnEBPokYKT/gg3qDqQZ
Z63CkKBjdtka/K/FGPhUx8niJhp09J/8jkOXGJjGM9zt3WrDfh5e/mPWYu/LZcyrThHrozfuzfGN
Af+8TFOZTvFQZtEjZCy1tzC4qgQtgBBPQE8NMePBqukq4rDbgtxUXROgb9Y2wmXv5Q4t6i5w+8vH
z4tHj62fZQXk6AvjOwFLkE7ut8Ii3/HH5VwMB2NRzAgTTvtppC/ViXrNVzaljeiddAv5aJWPygji
phCOWP1l3KWFQ5ccpqbGstwQS6jEp50gIaeXMd94ii0wSAKR0wHF9Pens+yZf1cOzpENGWYK0A7T
YYBVrVZNb/o6Fq0eaDZ/tAJIDrcRYMxkWXKHbrSfxR1muRlHhqijnQvQlcM2U0LyaIUW1LodiJcx
yeX0Q49VH9C6DIjn2caQnBOsLIfGTLgh3hufsxBywBNg4/WUp+SW7RuJJOz5opnesEOacq+aUlVa
muxS/07vD53I726MIGW8GKqDSJ91bH1kgEYzmdw5pXyc2iB1xR9M0KKAn5Snw2427LqxdmFA8p+g
h5/adF+TR7t2YgbwkcWKi0QJNj9kQtkdqcfzIfV1XgbO70+TMewiOR/XYF7j1E8x0yer6P3fLU6z
7yvs6mGDRfYevZzl8aVPgik0Fvq8lK+JyAr8W6/LaXcjd2Pe6haMa8tcX2S5q3XbIxobpLbyyKSX
7hmbRBkpMinDKQ+KExllZPK2oewKC7SgRyQgtoktdsXoNr0fmaWH0mRpdEo003KGjHvQfazNY1/T
mixyzF3vgYItSqLLdExxYglBDrZK0QCdlb+L28WodsgYLiq4YlqYoM+LZvwWF7ZJKM8Lfr6cQV7s
7/p6EzuClbdx4txveK1tE5OVR6YAKH+iTCtC8XOx378JnAGvXUClbWyKZBUVcNNYPW5fzqR3Ersd
GEWSwB9QancMg7SID3hSBfHHSwuu4zBK6JuEmuqQb4FtMd39yAAchqwQt6NLGIgOisG6N3meDP6p
jG0tU2UydbMUO++2/fGpHgtHz52ME8t1Kiclq8fIDHVZSyNxm0C/UiCjXzcbEms+nQO4aATst4Ed
JELj/oCJMrei00KPSPeykqldbS8c2YHTywOrclT1XrzFxIDLTvm+Yksy7md+ki6O1/TRbvYAPwvq
CTF62wymRifuljYG8qd64POBlGAaZurtlsVuWJ/9C+C7di2zBaSIbJGHvs1gKYn70Dxpa7dmIk+Z
VQvzl8+Ed2dVgTy9dhOhPrJUt5dWKlgtrVeUlPYCGZO5JA3Kzwl8RqE2KjY7GOLRkqey5Jyv73Ly
aTxZVZa+SLIRRdDIGaMYE13Cd/ANjfcSetwwsajn72xQR4jVwt/TXxo+cvcEVyKWnB5Ew+WBN1eL
fp40onTFbg5eaK7yhsFWJ1Rfu6FuZfiujgj/+xzW9G/qvHblZPkaM1DdVZp8vJZZHkC4saj41its
aAXC0wXWKeBXbIKSgy1xLJLx3Tn6sEtx/oYp6tGwWz1GAC/8LF8fjs/a2+XGZFyLQh6Mt1SkXSLZ
EsHWtReX8r4SQomJCgFyg+YoiFB/NXqXaE3TfxBbi9CwpsY22X8F8sd3J/gv/Blb3DGyqERF6AVz
VZ36+egvjqsomUGzp+ZN5fGPHfP3AETebJxs0Rgk5vwRBmwyJvan8eWwUngBV95pDML9Z5AVcimg
I0fOVLxgTD6zFkxj8PwI2WmSn52GyeSPZihkTHv32FxC+g4vt6UAiPAa/XfwixEFqnBUldM7Wbko
RIAUnaoEObMCEsww/i7VwTzFghSl+2dOk+IXe9fOMPa213N4pAVTATbq0g6pCE7DyXmDTcHLTmuE
l+u+lYrtczHmPypfYFFHpxH8GUFkuXqQzuLw6vm/381gkkn5dL5Z9RmpW/6IL1MJ3mzYx3FQG4+W
JWyjnhvtyzdNcYtTrkS74pBOfmOLU+/6YcFc9pxYGvWUnwlbtj38ysFj5qsLl+dcRwJz+skthB/h
U7G0Q41ciD4gf+SdS31Db/Ndn/tbSQdPsoaiUy8Rca6ksJzdS2mea8cB1x45NJmlOGPM/gyYFrcG
2VUFRrWpYTgaVO5qTrPEwgOa0rP1HTEfiG+YWHgx3MkqXwXJfy84F6D1WOSXNrOwieGj3LfLGKKk
xKNW6F+an/zF1xx0Ivw1ILo2Gathgz79GDgkOcQZP3L6NVMNpbKu38K9rUJqGp9fEQONfXQ8iDCl
dbo1ZP4XOyD/5FAXKfXdjxlUQBd4iEUp+gdVOvxpLyyirmygLuHlCHVsEuf63c9tmzjImBFRLJHl
wqiZob3My976tcDQgcOrTPD1oQmEA70Xm41DnK+vqI7Oyrdex/TOnRn6N5Sp15RhsgXo8+2BTJK4
aFOH0C+Y9gED+rL/skQoh+jSj8JtbCcY+dPj3cw5ifBT2VwALWUo898kklw19PgqG4SwZdmxKth/
aN89tYAHxgN6nxAEUkxUPV/gUEfeWT9Mx9EKmgPE3T6475n0+0igiq+Lfk7TZY2WV69DBKuLCVpc
gtzbZMhIXGrjTivHQFePmrsm2Y+s7+u3cwK2XlROUNsggLVRf5ZJg3vOI/v25monC5b+JlcdKb1s
i64iKvBPYvvbiKjwGqAfL2y9VwbPAL7J6eSYoQ90k2Y/QC1t6E0QIxZ/oUSKSbFdS/QNUVVEvjFN
GOfMz8vAnJlVCwcFm0AKqKQzYZ1dnONwDvLvjrOlvAe+qwigJGmc7o7HjfyPPCrvYOS8xetcshPD
PWEAI45NWG0IwIXzWPh+YOl4tpT0j5hI7bb+lE9A0FT0dBSEq5Y/xgrf28+W8Q31NA/nV7UrKB1I
GJzjSvMm/szWW8p4Hx58kCeod+KmEYTTaJHfdzfxLr94ygKS74Sq0jG13XUI+wJweuKcrs4+5Lts
c3LLAbNlcU+XQIg0dlYcrEMAAx/otliUxZLmaY2B4/CJsvQvqphBVDvoaHkdRabx7ZnKt3DeZKAW
0lyPgkiEOqGWEHJSzRFaZiDKAlDGXLPapO+QGfCaZyGc8oi685g1v1No9VsLtf9Fk5fX6lWF28kD
WjVi8RqFdKi9ufCXESib0MjrJNrsvaRYmXn5q4N1Fm1yzg/cyqUrUwe697PY4MLv4M6R6/jqYpkA
vTXzxMdwyQiryVXJGqcoioizvOEQRRH7hKM0d7t6hkCYdpOpeK8lawMuLT2oFUIZkMZqo8md6P7e
Zbov17wCEaxC9DuWFDMMO2cznygudbtd9KsthLLxRyMy9KbHztUp/2RLQ38FkR/a7nrgFANMG7yn
w+7r/ULjkI1jIkqyUjLfm4ik2o9NWYbRSMR+Qgj+tMaoCzCPrEbCtf2JxPYhjNj6MbPvTzhGgjol
pz5agVMWQ06EwwZuulhfH8F5IceGZjhMJo38g+Zav/GVbXwAKoJFmBte+LRictoyqTYhLr9M78yd
y1kv4zMiIbGDcTrIWYKioMqmdqo55GwgYn5lBfbchDGcgK0Pn0a15IIaqJfbHA2Uk4HY2czjIbwt
LEAw3SodzyqsjohVRf9ux0KL6hytgUQ2BaeXhd0DoH6KNiMF7RI9vfIKR8HlUN7+yVUKJNAQ2I/V
IoobEqb1+G+X4S/VdY3D+0/pjX9Vf9agwfXfK2KHjOuPgj6trlVT47fA9PyTAeS154Z6SFoo0iYa
092rqokxkrwJz64yMcdr6qFvzEj9CPoFAW3K4Dn1nXAVJv4aUyqyvQQ8KwN8AHTT2KAqmWGpsUIc
0a398aM8AhtBf7eKBuDap3kOk53BlBO4bUrs6a3PYu49130Siev/3XVV6KfavHhNY1TD8kf4TpX8
f0nBwFvVuDhObht+xvPxU/hdpzaIADa1IvzzTQ+0ulBS1s7nh7YVkuXTO+h44kgGMA14g+YpcOSl
bOl7zPACqmNhGqTkiNFzhgWB/u4baUfer7JT02cq1spiW8elvv9j4NqdpdyKboSuyz2SDxy28zZL
eJC6ssO2f+CBHcNWjKn2Ved5URB0dutKBZIrvEnpdznPHxXHeOjVXYQzpuxq+SYmh+/C//TV7eIU
ZgoiQ4AZnmGi1vRwUccz4cFWtavxkTPWIFR1Fk7qv67BdU41SU3cDF1SEPKGq8bdUzoSFUT123m4
XKfFkwEr6klVm+EFNub0Arjol+e4FL+zLz+cd+y8sL/V83Td5HizS97CtN3GDHZDP3pl+GdVp//j
wsvrPefVVmflAAIwkBwnA33cnxXANoSbn4VMdYqT9d3WGYncjnjAGogaN6BsU7dCQIFR+PCPfwkB
XqCeYGHiV3gvzUHy16FJiDNz4J5FA5l7jOZn83aNLlJJrudL4FeZSAgzFzRQmdbEcNSDy9sQoDzS
K3UVJKJZM1XPK8MUHccZkp+29RTv2NB7rKFo2U+NfB0xa1PN9i/FLFulyj0FVMExh/IwNT81lgKO
qSJa8PzaWFrPUCvbEtCYdVBF29YDX2jnPPDdWLA3MZl+DXGqc04WFTxNKpNKoTAmAqT7SMPKl958
LBHAyRGStioRo3KTxUU4nTh5wK+aIG43O/afpIwcPkhArPYzICK+FkkUAP8/gl6ukwLPjDSu1LFc
MTEJN04WGpqBWjKQlR7ZtgNSps3VePVa7rQ9WNhl5l04dGlJSC+bR7hCZvKJRBXqaP1D/Irzvvhm
4UhBzcjlUfLb/Sq6E8+aIt/Lkp0eymKj3fmF3nX4OcGwP/uzWUT5QYxapbY4AkCE22fgJ+tqBR2r
bDnZq1eeB0JhdnePNcMYXberwi6GTj7ZuDTCFUYhHSrEvw8aEtOR5fgMKEs7I3+08j5hJ8tnaMPn
j1BzgKR5Yxf9XrqoJtf3nofiG98K+hfFKzUiBJJGWNJR3ijCBmdDeTmMnMo+C4UYXiNTaNfB5OUM
VPPk23CxaSGUuIZAqmecZqUOQugED9ZU8INhW6JtZfYOioAaBNH3nn0k61DZ5q0/E+H/3xsjo4h3
ghBhsk5WFk4uBij1IT8gT9Jg0FjJY7YwLXBvd07Aob6mLBdY+29xeX6MkNOEuv5enSLlRsr4rUj/
2Opgz3Q62qhTE5Jj9EOFpY3vwrgnVlEwz419W7qhjGPKaC9CIQDLTPWiCE+Mbn/RJUPiooYfg4Pq
zXFHM6XoAYQCE6LZ65KZAxkLqwEZRuf+WMDJV+NSw25qHIjVas2NmDc+1Ulvhjs6LJSkjO+miJiS
DhYz7yvmVfWBq0dQshqO5MADsZqYy5UIUTScLSbEyydlDedu1k0XCyprwbfsEG55sWhq3fjgfGMH
mqizES6Sv5X14cAFyMeSh7FM8PoXscBJ/1yBmoVdeG+gvsr5b64JdRRgTuchDIeiUunTPUjzuoHI
AzNewzNy2EY+v2pK+su5dUhJ+5l3jc5F5UJmj+wjUeXp0lQUWcfARVh7DKJi/tcf2hv8WRuznbm+
Ig5SIL/sCFMx0EJTMyP/iJ1I+RDIvsTfh8phJmCzR6eZILymU/12yjtrqe5EHocmiKuDddVOS7IO
VO751Z0ZIvIYfOufxsUHbWH/c9fKE13zeqzRImSRs5gdIkuMoJrg3kwSAq3c5SmnoivysA7YF+aZ
krfF5gp3kBf+cIm2dtUZ57sEto5LLHcQ1nROkC34iiQvfAOAfrYLclPZ9gA3IyBpRErzhHObvZSL
0EKBiHUrnuOykZWmQ9Bdd5NmSmZuaDbAU8EibRFmMzIhXFRqyXf3UG03DSHtSRQrZnk8uek2TFG8
hyt4Sx+C6ki3j0HIDfzY7TqgTkDbw9QSiY2DX2wSrwTDNcIh9293kbSOLMwfLGyk1Gv8TOY55cMa
MjQSvqu2SmcJJbJ7UEirgZhFfhkdWZLJMcVW2pcZ78pLmBRh1keCf+sX+Gyx/8feM97KRN8Xjd7g
3KUbdU4dtdnvYqcxHVF6fFJxbC1o1GyEZ5rvbSpU+rUXTmcClFsrPhN6YbinAgWcm/w8pDdWePbq
BgLm6QB8Ozth1hqQQKXuvy8PJvsIXxiUgURHy44+szlPv44aefnqfoeaQd5czA5d4vaMugh5rukd
LTnytUsbAYHEnUz2m+hoxGkxOBvd2/SOrKJUbSTEl8gF+SyaRy4dDeTx9rh48ZzPDLuParCYrIOr
2vjl5Fch4CNORLJJuatmYeu40oyOjduUo3/od0uvjXnCcPKC4CLhZcmilV5RSpTh1YcYiz0B/8eB
qMfgSRuqE20wyE47zgiEYgZQ8UG/5JjQWZ2bV2lGFCmzMs/CgcJGNQIc3/qYzjebxNsYaiLlJuks
IpWxjukzrSmSPbLqJrj7C6PzT0XBodbrQAYygT5p+5UaqY9g0Hs6MdKvhZHhyDQGRy1BaLx+42M1
VZunFRqQeu9/zTyF1Ds7sejVbG7K1fKvkD1RO+y6nSdq3qb4H3C1yy/iu1wL2hoJnTw9kbY55AJ3
Y8yU/WVs1t4fDvx73AZzwDW5WGxztHhc2r+Wx/59fKXTSouCQ7VJjDS9RfQ240+5+V4jn6wA1ROx
AURm8O5j7fsK8aVB3/DtqXD4+Udyt8yS5Zu6tQLjCqrveq6d0QBRFK3P5Ve7XWzgSjYtSHKX307t
HR8s1vJyVVn0Bhv2onTxcXJSATay0UAHbW95PM2FqhIbtol9Tub92UaCLpJKxCty/C0jlJFu+x/q
MdhlYNRuFdpl2t4ORFR4Wm1ZjFDuN9uKBYiexb8ipxw/H9uRI93awgD0EAsp88Os48edHLxE+7L2
qEC1lUhF5y5QWw2vbvS2uMLldGhU0y/FzmeQs/QRO3A1Ua5qIAPZ5soNulmTscaYtN7TYcaQy9qU
YJQTshUi5ltYFphMZeu7epKfL72iyKB26DD2ZexF4YfjeGyk0l4IffLn++tUluYf3fhJX7Ho/Hc+
tO2CGktIn9daUHonl+DoDw1X+jgiYlB25AeuRJVsVtCpTaZVfqYhodFo4jwVkjZrAaA57K19PFen
RRvV/EfvnWkr2jAlDW9EQIoD8sqflIuMzIKh4iDKpF+Ywx1q6q2qyWmVIG3DOj/cmz97TmvXZaV9
a9nxWkGfgm5qPL1Qt53EL7vHQ3ULrOXrS3OT5CMZa4FaDrkNjF1/AXMuqNWfXLu6L2i1tM+bfbrp
1eguBf9IvM8NJ4/r5mxE3FTjDgx0GyGKD7aNe9zVHZpeId8KL/SxaYGRfRX3Q97Wo+69Rz1YyXFg
VNKcAlubOKiKxeizRV0cdlAvOpDNfNcEMk+Ino3N1g+g5Rr/5Ux9q+QzcKy0k8kRmcumDXIrSvRK
jS12goac+KNM6VTUwtu2+tOfbEFiea8i47UAWu/jIeQHT7vm4OCghu12OIHH4qOASVDoz945PJHR
Jqg09A9qPMQqLmLtnGbSeJc3IPX5QBmX78ivm3ncKBUG2XwJs04OtMjMBbA/oGg8Wum121eea9sv
9u3FHhegvG23pO8NftERtJQgjjpjv2Uqb+55kvLXEG6cNxGsm1S9Ooruu2Sd/VadbD6Mqh7gUwc0
poQ9kK8mWDDJx5uF1qSLsbQb0AFY5+cSvYeSng4JpcXvWa9lqiQ/Kvat/1b5/4/2ZUf/DEx4nfTL
QywwURoyzdJ6pip5Vh+GAhVwFRNJvSiJA8KC9/hclqSNbQYgMhr90an1LW05cXuuMLKwlToLT1+f
6G/yRujK2yU71fUaOIyr8+a+dgfU0krhxhAVkdu/4yydedlL0+dx4pOWj2yPFz1eu88baqZ3Cxyk
OWo2JuRYhCwxHLjnNb+FNuvHxCHfWp6v6+a/4qzWaWmzqNYNnEksL1ZbrNDjR57QisxnRmEsjlX5
oGcDkFFMQRp7K0o9ERD+7i3VCXodbt1vyCblHefhKmACZc769jLOGWAwW8QzKfURHSf3jR7MmCOx
fIiKw5vnTB1roVTyb5WSdu4ioBEkT69DI0aiKPP+WEL9yAACbKNH76rDsncpDnzXL5UnJzuYgmMc
jAzOtT96TfE2j1IDAqj6nurAB0By4S0vraHTnoe6/5fMUsvSgSD25H+YqwRNKEafNpwz7qn7roke
16NJi6sSkgN1IFe1MaxeSOilmQ9URPOL97a4VzaVARY+fCrosMQHnGFWWs9KRYQeUa58jfgR/8K2
UJzTecMMS0frxR+QjoKdJ0bMen7lueE0EFbg5oHWH1qZkRgx+8iPdhTtRI5KKxxLN/nrSpICBQZF
vUeED9fsu5B65mT11kNNFITzmpOueeTRBBk01o0v68Jmi+AiF66swdvjSj9mBWQGOpqNGUNdXc2j
oI2GSRdJZ/riXKDaCuHc7CrUeoVxLXAPfmX0QFKrcqouG4lsiJ6KwWWK6unvLcW1Fl+5OwveiDSf
BddElJtXDyNugCMYDLNrV2RQvg9VaZyW3onitllx0BEzXNItoZjv2wYosUn4Nytme1q/TK2Lyviu
SrwUwzW7CabwYLERg1y4ZIya4pZiJ8ina5ybX4sipMSBa4IfEwm6LbAFvrbqztsE9el1eus2vcpr
UxIJkMYDsCgWgWeM7mQMz9uXEMjGZcAzeUXWtWFYphNA9Li7ZpQkqn+LNUkkb8/VngeflEABhvr7
ItDM3wY4kxAO+G7TIoBzqUwZR3EstJf53dl87Hyb5XDmvV6SZkyrABzkUTvgoMWHFuJh80muH+xP
4FNbcR2CldvYBQrPjK3kkA6D71gjyZXFSKw0WHUnFdyE8oVGOeGL4XtILNyBaQtAgTaeIHWb+nzg
xsA93zH3GFvQCEe56YvjKQkDX/CbceayjP5koZlCpzSppj1E85vgWtW8JgC2MiSm3DawmoKc+pyj
P98g7/OudjzNpI4RNaFc1uqKLfQk0uI+EKBkLirG6D3tEvmta5BWY+kaq+5wMdQlDlIOJsNicOFp
+gky0D0L+I0ITL1YULglafuBJu7x1aS3fiNBveAQC/EIpZv4bOIas/2Cx1ZycyHY8mdV/HodqYnI
EUFiq5m+LbnNqCpz7LZdc0X0KQ1u4j4535hpC3AumNQHk0wm3R4AUydyCfOXqgSBo3SyTy53Uo6s
J7IXOIoL8kZIbZ/gCsxuYRynrX83RE/9te8EB/+ARdfmZvHEgUBKLOKtLOM9xlbgkCy91CaeKtUM
BFGl+1ZUqkY2OZkXKMONKot2SpNahnfwSSd7VDsgCrpgLUUj4JRQYCgeCdt+H2nNdl2t3Vz4HB43
EerqdYJTH8WTozJA+pGIb1uqIQ6JMTsDYMddpQluGVJRauxgv0YsLFMGcNoo8YHDTxjlt2sDiqTH
Uh+ik+P8FPRMDv+oeX0Npvz1JJA2Zmp/vO7N6tF0EtFC37guVj022wEGWNRt9zq/M7zQN1W7aJ01
usufdgdTII7Mj/F0umB0ptFC4Ebz3JzroZd5Q7hU9sqE9xA8xzsSnQngC6nvQb9zKIouSlswCG7y
C3gcFHU/5R30E7X3uB2AHNWJxWpbHsIvcegNbKJAkFP6GWoLm2CEm/ob46lDBxR7cJ7GCHJCe3aY
tkIsPR777vT6fPu0k7YelrQoXsdlk6OqJjeLQ+TtAub/UML5TlLu56BJRZoM2maqGh+M/dyon1G2
zEcEmaFkyW3808s0xnkQV5wwajPeKD8GfoZcNLLhmeYdrqSdo6nRfT4sak+zDycc3BP7VHaWjoyK
LyZQKFcK9sVX7ioKNlPkMYact6ORv/XRlh6eLC5r+gq5VILHL7aJk7/r1N6SfxtIazWhiTZaHYHC
QKRH1UXKuNwqqdgAGJTCUFoS3Oj16vLqrxmbsMjvnBZx6TkdD1CFDyH8/JfVpVDbb6bKQnZp/q9M
Aah0q/54ozSrnrdC12UxL2qWiEWJ7eacEBjGqQcMXF8N4aTa2qTMsWZ+ETxa/S/0g3Oz96ad1RKy
03GmJ43n06Qup0LvXtBPRA9oAZHVoLyZpNHAPnlUBwWvSIB4PkEtaBP/vRH9ZkEKcv2+DZYO5zvx
EAnE/NMyOXB0UxjYCQmJAyo8p9BOdJ6ixJxZkLYJGVpAOuaSTzLOW3Oh+FYKD74bxobkrb2BDjyH
y8P8ilcQFOw9mSSzwZoOP1WD3PiLhfl7n8uxFW0RCnd61zYWRx2QZtvgx2olbGZ1PIaWwnFoDjng
yEf81qf6+n5FmVrZ9+eaEwoea1FBIerXGbrNCOhnlfF94x+ksW4Y77ws10PERyMN4TJYUqB6maSG
0erObSRBMw9KIDujn9JTdiiaWWBO+I2YtXS4YQXsVA4hlrIKm4M+DVmiJpiBop0rXLuhHu6tzlDY
QJz9VyOGL2lvdy4zl2/Z19pGLqq2O1TJUsfq2Q/BDcGyuIj0fmVK/rP4fNbv2JE/0l8EYI39RSfY
fKUsA9abr8MgQTn2i7udv3Q79zH1ReYTH1tK5W/XGAkxZib88x3YUGe7XeyaxOcVTP7Mz3N/xXsR
fSLir0laZ6WeX3+0REGUGqDtX/qjY4YuL882wNKaFyj+mUPrETBFaoIIovtQu+unQIAmXcMIg3wJ
CluJTL6zcIQnmCDoQnuSgqsj2sfoZP6XivMlshFap0ZGfmYLBIWQIZurWmdkYGD5Zlvk0tQb0Z25
tLaELgqpliYXiNDrCI4sqzsJlC4EC7Qq2ilkw9wTEuacySq7LUo/slyjwir8JAypKWgld6JkLfYs
kF+YrtMwwEX+ysLGrHUakrSOPF5PezpWz3c/bIchEO2bQij+B9SZ5axBNu7f3Rvo8j5el2BJQhTn
0tBfkOLetvlEpB75MIpdsEfdzKZG5u8Mppn2Yc+Z5pVd46kviCIIRLdtRRDnG4hWV599rxCGM3W3
xb7yJ2p0m3CJx8YPwKJTF4zSIPmK9XaEjRI4vsYPh4kC4i4rbceLMX/fvVeaFYFjyuE834k1tJdv
A8ncmp/4f+PIiy+6zBK/ebuuT5bPR05ACGLgonwaWGtPwVBLoAjkRejqqjo3jvv3jNvW/YdpmQaE
pVBnfmMVTvgkj8iqZbnsaXwhTLPp9k9G7S6x3tU5bErxUkoRQd1sOCQ+HubuwiC63iqvQ6Orz1p0
DedWEzmJzOdZD+kMokw5qPUF7px9vKipQPYaUibumDE8vvoMhxjbvpD7QWSU+0e8ycrfMcRsGl6o
a3tlN2M11o7BHXRLPiGt0+jrBQ489Nh0Z8m+mr6FMp9ODQHCwP/UbSY69VWdlxokgCKZEysvcPWy
5NLkYLKQ6OTGHyxajDM5ePMpQH+r++Esplm+awom6jE4lZomBzdoDSfVHW7/KPpdDDn4pVhwLlAn
arxivBXY5O0601JEVOTXn/km7Uy4VGRSddMD/tf8at9XyvIoNZmUK11QXaEcwc4ayBCSK3W+9Sth
ABKN91bc4L56qN/0SuNrn2UkOVlsCfsLSRyB9nt3Tg1BA8y2QkxwHpDNRip7h6lC9MFbUeFH27oy
M/smHeaV0Wb0E4TaIcYQRfyWflzDOcwucspi03Bs9qIcIiAHOfbYuxF1/7BsrN/SL4cv8YA5flvU
JRlfamuAGPbWyJIPM9egg6R8NCCnJrxg8IatxwZHcnhIf4TztoikiYusRVrleWCfeZw/IzCvKCmd
WQgx6eqmPaLQA0OI+nXDE/TfyIHyq9G2W7wx8942Xm3QWdHOQ1X9zwOmZxxNFq8gUXrHHV8GCOfV
NYme2FMUvfxWVsZ/pLf8vdoEwVIaBGPRCw6NN04T3FS2iGNlKjITcYad9R1MUETlJogAokPduaif
DEDsutkCmVN9EpPhxuz9rtPNAj3izfKLLMvKNH0KJWxY0W1DYGFXZt2bYb5U0VQ8NnjPDECm2qPi
ygovW6oRPekNbRO9bf53dvPxk28NWnip10Q+enuewcmUQssd729cl4bdBgqjQMoJQPSYclXx4FFT
Aao0X8cQkJhkKfjdu7xt7fBxEhGLnOR8c/8MMrRkwBVSBdTsHmLtHcldyJLQStnDJL6c9WmWtkzk
g+HRhFpxR+TgKtALWQl8bQVWFRjxT5BwbthR0aUPgp0qja0rtXmHJdjyuiPWRDA7iROCeLJUoHx2
EOEPDqD/6Iiov/mLfPhb/HP8c0wsHKCEphitDoPCq80cVIkSsZqQgHRcefVD1XztBjw5iXcCjVsx
KDfV32xLYT1lJAFZ3BqKTGYlrSOpXfw/NiHbBnlT0A6zBWBKHlsSBAIsovojl6jhX+ENX9BIH/0h
XYq7qe1WjA1AsQbm32tXZzwKvkiIdEUiqWSJV6xibsRuCs7HocMBiekQknC/C5oOuGsMPCbOMeRG
fIaEQW4276Intz5ITlCMB5oGqd9LwX8AGE7PW5LNSpsCmX1JnuoDhmzfnZSaKcWovyB3nj/FfH01
l1d5Z8FpCy1SWwEZIii2UyksyOkvXyEeBAYvSbNx8KO00yeTELnAATpgFM0w4wOTJLJDlIOOiAa8
AdbgBb9QRmzjuPS0Q0tVfxtoDRAD1R2QV/aJrqnSt1QAGWTFTOykH5am5tfzeF4GlirfYcoble2J
OqTIYqPSSwnJQsYhPMnpQAPmjcP3Wr1jHk5HlfYCHjnauGgDq+XgEwvPaofEQaBf+q15Hv8bFwPX
w9qqaljmaEcq8ZPhgvqx+DVqpXAGHfV6FBMr1r80JV7WmeFV0kuUSSV3pCpRiGP/DvrZh1XWK0Cn
o2KZLBlv7ZHLIM7ZKWONgNs7QZr+SeZIrO+kLfE9RUkBlLCrXtP5aDFQHq8Jv3Kkwn81d69od1XZ
n3UGWacRAFQcbcDZXCmQaQHUhC6SvSdnRySKv6QwgdrZWFnUY+N6hyEtaSq3bqbdy/tCd18UgPOV
t6GyZPe4Kl1ueRbTGNdb2+ntfWUqCwruZsiutE9PQo4pGU2OPR99Uu5ptmOA+A4/OyjyOvPHD4us
QcynNKC6xQ8fb6POetjXOJuwp01/oS1vS+vecfm1sBUPjHaVSR0vEWN2XU9xkfdoys7lszTLw2io
qVxcjOTaGIDS5/k1zhdaMxc3F920wwjhmUPSSFNqh2c4eeP1kbmElWYzUuiI9I1SZ6wQ9/EBH8f6
52X9s9TXUUV6xVQCZi2u+Yh2lv7CvHQchreS3nnG3jZBMqIJetrEc3I5X1tbGsDkSYY+kjEmC1lB
/M68iDyKBUwDxfmaYYgmKwcOj+L5Y9cxWxaYzxtYI2FuYWSz6pMuWcjivdxYs1moy252H5iZi5gH
+wCiONFjXaaP8Yal1u49LWkAt8UzzBGZee9+tm+pbjmIkfKUcdpSewDQs4pjV+PlOoT9MkXu+o56
G4nn6VARKkr0NNSFc0iohZjLjQWlT6/c2PgRWTQqi5dsHozuUEuv/inpQJTvXndLySK165oHLuQh
tAI+ePGXQfilLRf+kkZXeSVQ4fO/enjsqUykIOwRkbWZJuueRUAxJCchMtN1R8z2skJ3Cshgbejf
i1xPrG9W1q+tSrk0dQV1MBEvC8mkZHkX3ARplrlOOJHIr24xiO2YNzDPIp++PVctdgkLPLcOn4DC
B9xRY3ukmfV0GDVk0/en6UK/ymozVsR7q18PXwAeRYaPNJ5GOPwa0AX97oXtQYarMQe9e18Y4jdf
BL3A2yTHm4epfPJriAC6jjigccRgRPJyAGzErgbaX4hjgahzI8m0U3zZcp0O4xpKsW4GqrO6+bFK
rFXnuTq72og7cAEq3r5ag8Ps9KhcXzS0AEME53RJzJgAtfl2EaSeQ2LYEvjzJyNYl0ax6mL1Pi6Z
4X296UyhjTAyLTqd0HtthzZhHYJgRdwvvdEs47Zrs2QVgaykrdR1FfuxZTX4cgYms+pbB4ZRKUZ/
K/F2IH9x6XzmVSXtjG9WElK26Anw5yaW62fS8kDakAFI0PruKv6GzqnFvwJIALwEwegDDwL7Accu
EqLceP6DUNmDmXHqAjoDq/AlkYbtAwa2TD9mPLrJcuEHK4UJ4wOZnzMxVHqEQzXzaMLad21Y63mv
BQmoowGl3Up6SFFgrbXQ13KQC3ZUkvEV2dVWjiJnDMyCQQVAepNk9ORTbO1ReclGcM4gc6k4ntcM
YqUXEUqkLvgal9O+wD6ngyKUc/Cxfi3b3MtitXd9I056I7lcZ7N0hZk/eJ1DbjfaUzktEYv36oQG
f/P+nmUNAyPXjlteIPR2T/H+rwbt6kcsVnyxU5Yg3NORQHMn5Z+cCTBzNpQ3ZuOIvnqIM86mbN8n
wZNbOY2MDlVaZQ4ZbOUS1A9n2GL8dwjjEJi4sg8PN28+S4VK1M+loFJp45xV0b8clzIQDPs8vy4Y
8AszLEGiaLMKQGVj6cytB9x7K/g5pusT3Scag047YeFdNUsrCgz4xkZWLIGofRJtMlolFicHptwM
wXckBgF202K27dOLoQTju2N+bu73LqucYbNlQXWSAlBwkByGh7msSslN9a12Q1bKXL7g2ViA4OCM
AmcwaDqdGaeGzvzdez4+J2HoGYrYZQn/RVg/IrO/tkWV4ZCyS6sNUjzwXv3V+Qteo9FLL3Rxskdv
uQzsMVPpp+kFn9VctdbeqnBl7glYZvYD9JO6zuvLqtHqfs+GvtZk7xGW6Z5QY5/l5grRSm2AZJo1
WZ/a8UqP3ODz4cajuLIGvZovEoUVbGQmM7X2oZoIuLZ3dLGDrNMiz+3TXVmFA5Z3YL+WVc3SeGU4
tUcXD4z9iy1Cy1DygKGdtF66VqJ5At6atdy50wcAMMwblvW/KUrlMT/PwRFjx4CxMPtD5WXkIdci
3xn+H9b0SJ/PSwMR+ghYiGU+q2ENO7QaAo8DfUal9psoZxeESe0fr96gkuk/OJXIqw+3G7JvcSMG
S02L6VGBZsO21Z17vJPxyJm6AlrAHojpz8MaTFzMYDt7L7H1oXTtGJl61F52Zr0n/P1eQaxaq4da
1u9gec8U5iT0OLUVnJW5+QP5QqKozuj/1ocVwjZ4Nz3e/DBV8/G9j2d1qjEpAfRRF0DlBTVasenU
lHYNgkp+X4qynyAFvKp5M4uzBQlAFPIVkTbFbf+d+U1I0YPxeEiOeBL5T9NtpPMLvHSa0ATi1Uwu
09b+m0hPedPo+l9OQ6vW+7YiR6iD3vMPtHqiMzuNpoCCwCY/Gv6XSxHA0KUsnaXDjqMZzzo+A4ZV
n+mhkQW1dDrkaapHN2SuxA0VJhhLxgIdZLRRlZcXnny+2lbI2r50ToG7Yu3y5cpgdSrJFC8oC8jo
Io3u0UZ4K4/hEjwgbu3hf21Talq8GtxqVfJcITWwMaoSfTRvtdI2JxXNitX/5K065Rha+/O/78XD
XuGwkGpLM0JI4zjWGTM+cbH1AEnPzdpx/OYbGj9zjbRkoIzbBLta32uKWYmJal1KqiTjUJlXr00q
BonXFUoBuGIQS3xfA1LYNCYFCMZKvowiL4yTiX27A9WS3Clsy7W3UtmcXR+RqI01ev6ZJTjzz022
bR/JIWAO6TmcbAswZqcv3Yc/p0t4j5fcpc66R4ntijqZh7qzADoGnnqSh/8GpBSqb9TTBcJ6RMk4
Vxfyq6wQoskNf1lcJCOM3KKRqaF5Zrq6TJijwxX5TXC0K9TdpY0+Xw8HFExtyCLfGpVRSrtwYAth
Z74xZUpbX4HOX8huMiYhrnthyU+SrJ/FdeOnIT2/hAuPbdCvWNx68YB16NUBXIXrDq74g8WtIrmW
zQddnzk2GhJGmiX3aGm4ZpjKyYR4PmeeVr4Le4Xo1ZnYwrrTiWI81tAs5um+h4LfVuKzkWGwDO82
i8nROijaRu/MBXcYxabxZg0sZTjHJcQEzVjxvUL32a83OP9svF8Euz3KA1gPckMD5NbSQTkJssKu
cz/6ndo3ZvoRgiClw6g2EVK75ijif2vISkeXaZ6V7lwh5hNkwF9Dz4uGFKkHnASwIF0xOASp0n7U
hbclw5Sonb43leiv1+Oihp8rmpkhURG+xMfFypxnspdD8iiPhEtsUcg6LLt38FeTXnynLkH9o09L
c3MLGcJ7ypZBMkl2vUKTlb+ZMyZ7XNDRLWfKdGrrAGn68R/aQPwg+aGQSVimePkVrcvp/JCTZqUw
Nv+3jbjkRxeycd9YmfGDBpq7Hxv4MYt0505fulEX7R7IYBWDc6/cqCCyzjDJC6kQrNNBqtxyR8Bc
9pfp5tSr40L179RhdZbmNRqC02KqHM5w07FNqdOhWOtXHgtjssP7tiXgIYyYICeIA0403CKTC76c
OW5bz2m+wLyqfxU9ACtu29RHj47M6pYQXKmGMl94hLZqQiQ+HORkB6H1yMJy0pRqXN+LwG26dAYh
D3fLVsVUf9pZ6diaPkF4gTnKa6OWXRosNCs+aRG5bDwa5x+W0IgiE1fr4PxFmxK3SyDDugZpK1Dg
dDF0v1RKrGgnUPWZBqojsb+DFdAWmmxmy15lIZUK1eynbUyT0xKGV7M0muOb6IqWiaaaHQhc04nf
UrY7kaQW9VK/BJ605nPmXglh74gLd+dxmAQEVYwkEStOtc7P8Jw7PwdVRC2d4303fmv10FdSAvrL
3djFokC+iynykLwmv4I+aydUsFb9uERGQucZkBrDFnEa2Rn/vd/SgWF0vMYUWHd9DQCBibnsJWSa
F6QVdDVFubEFXZAqzx2SFD/skuCVAu4QujfMzRB4X9n4oe8lAPIbjY5JpMpDpoX9CVafmb9GR6Qx
v9AbmbORdexBY4KO1Yh5on7F9Rj1yHvpNJBlBQdx98/+kdA07MqFAUyqNaRWhb1y1M7QQFAsHGgx
QbQ5GFbJfW5D6mXNQ/B6YkmAqqbZQFJOJ1tlDoEEhvS8x1F3k1DS5yqBMTVuA4nlkr9vPIVApJ1t
AsU06hrvg0XR6+41q9fmG8nf9dz1J6mcx7HzHE1b4l8GY1ij/h0FITA9/SkZEJtCCsaMuFexDI0E
wGRoqgkihPcLrQfRcBxAwQsV9UWNOOCfadz8UAdfyFuAWN39pUo1fGNXdwMxyPloUnrdbMf0XMmM
fwZhvtrkhHD59bkfWVuRdVht37MKs4Vn1Ij62IEaTp6orDvDju1V2YGYzk8kxL9PO7UNZc/Ss/Ia
lwSHUUOf44fz0bMmxY+55vjHAlrH74gog16UHcILj+ayM8wD875fDA0uCq30oqhXS4QroL9DTxv3
4RfPKvI4gV0PGfZH7yvTO4JYLeOutuFydgT0QzpHNsOH/J4Wqg41Xhw9rvnnAC0MSnZOUAX+GU/m
M14j7XpB6JAoeH4kuQ8WnyZhPuLPNGEsetfw5e7oJAeKd0/FhTKGhJvQfOEirlb96n3WmpC2c96g
E37pTzRjXb+O82kq2nsZRsQEsY80/vCtkPlm3RlYt6Oj4Bt3S/80xYtigBWPao+K6uE9MBic3k6N
X+WltFj1eMFohLxW6tvYI3fYinAng3a5Ea8tyj6tOAc16+h83HflJOeMPDCvqbrApG6NfsVv8AEU
+/Sf9jiQgLq2Qdmh+/hK2kFjEz864ylj4q5hVoREBzNAPteUIdwkp18ijk71DORCWMl0hB0PEDmx
i++AclciERpK8FgDtv6LQ11an+pjLjnI0n5u+3r7UP27imBoS9dhmHRp23CYcSEPcM1HEjbeSG3O
oiuzU+y4zHuQUvBAWIYwPtN+x+60mr19by9yw6pSiSdgnZpRFuSp/xH03jAxU6wEVcsItPV876Qd
L3sJVp5Jz34W+eps5hQVyD/eoElh3jLCUJqZN3XmgXuN6IiUii0IK5sJDvf+nFJsrVK2vjnh31AE
C/lpHoeJVgbw41vQbXxMDKSYQGHb7NfE/JamDzh4GSb4PZlIxNTiEdKNEYorm8qACrIkSTXUnyew
quPAuFdKsUcof1LpIhVFxr3yu5lJ1Fq1rgpzaF85KZwUlng9eyVwkhLqBEe19RST+bbHCsUcw+Ww
OQKOdIRB0k9LDlBN0HAqEN+pjvweDW2x/pwMZgbIgQfutosa7Z3PqRheViWU+ACUwQN8AVvzK/gg
nULPD/6MKfWYxInIsiHTDukIMCmW3MQRzohkJLKzafpx4e7h4ssWuownBrcsF8cUq9m6WlY7AL85
mHgorJ8kBfwOCOWitoQfwS4KCYOwP9UzGpFZ3s9g0GnDhD143aZO5qTyUAJHe221uQ+rMqB4/OeD
AcubGcAIGwyxqmv7yJM3t6Y/wXY9elMs61a6m/B38fSAYKZrlwhl4KintM1+LBDi405wznL58e7r
isLlUDhlAS3BVDH0JgCzwo1nVfO+eLk+cfbQRB71c+OcjZ9EpZIj8St5JRL5a/FTCiW0NfDlL5Ud
trguRLikvVG9ppYs1o7/KOToftrUa1mGQujgcxYsvfxfI4h5PWUj3i0ZvSMtqpjOHHs5kZQMKQzn
uWOeR5tjXgDNhbWSk5QF5ibig/A+6H9sY/fD/kl7jQUwpjLDCA+/OQNZEyn6CGHzeKkbnjO6j1cI
y/S1lE6lNnl4W3P7j0AVLTJeeerrKKBQNLZ5GjGGRdAb0iWcKE9hj4R9znKHcEzCLsubF0AbD8rH
jYmBUNq3d6BIb+Xj7IzSMa61kQvirDoPu/aLw1DtJY+H97ejKlZwxYO9IH+/z9kE5HLrtshaTczS
61cEJx+/mM1gYIZYJjzP2qyHu3ytArzZrEYBVxqjYLXC4iaUfoehzzzuMGWqFwGsD89sngQfmK6h
EcvPh3QlwY/SgdOigxV3WOCCpinDShXsJhYwzpe3CwO17BHxh7i0pJTd0+3Jr3MzJPWa1xf0xWkb
on/prguQZf0HQrq7R8Z06AIApY4fEYgHqW1I4CrnK3TZ7s6tb8Dm3WN7QJn90/FyezWYPuMW8XVy
UkeeyUZlIh4igb2aXYDD+VT0L/kLX64Z4NaU7sGkyPhpry/4KfLfk3zjBxKQxoDLZIyevpQtdjMX
5stAa/XHMwTqVg4B6pIBqng07n0EaHSRIXQMj9Azfspi5pQOvyQ+Us0QciCxhhV3gprTWHOu2jMs
zx2SrnezCxz1zfp9yv7E2hnBp5hPfWbhM4/0J3FxTAbZ7xwCIt7uX6RObQqreJ4Xh66zNRdx+ziR
Jd+3ZZsOx5x+AsRoICCAM/JrlpQq68A9mKL5HhOtSFZY/0XvcKbVBFZdv/f/Ul/Ut2H7rLA1xfDd
qCyVt6DqHLzogQFZZl+qWj8SPXySIwZC1WaRd8uf9c4bEb/3iB9BUdh5IG7xm3YdktncWjVzIUTg
3pMB0GY+yQCKZwBYQOrnP0ChRh/SHjQQHnqYDf9l36Vmvs0axbFrvO81EYd2HO53ZNRUUPm3559W
KDezKofhf8FI6T/KlYJIBpa1fX3XIOrNVvpHiEfZR8n9Nn76taQrkCCxEZVRb2pgVoV3wNRM5sgq
u0iGfPDUt36ay3wM+5OW1kA4Avo31wGUN3E2t6Mm1pERXPvTJdbrKDRS6mWqIwFWmygvujzjXbOl
sBdPTPrHBY5gTs0sGNgYpITO2WhboOIr1QNTKlU5m+cMW2cHGZNz4Fe9ZZ1QTShoCAv1g+GHdO6b
hWESdokoOCqYLXFYWAKrbQ/QYhVmoHk03aY8uA4HuB2/2Lyb+cWy13bTRp9yDuWmYh/w+HkoKWzi
qJhTBFKFuAYaVw35YYfdm6L+VMlJxIkjNGa7V1vTQ05BBnPPwvjPV2t4AHXvXwg3e2VFVWW1p6r9
GbhE5nCVPIhCJ3uiCr7jAmAVDqBa+FUZ63cXX1bpT31Jq3cjXml+Ql2XvJT1VRrAxKt/P5Oezecd
ucIbQewUvgcuKHiuBXe7B7ZYfRDog9WHNs32YciN1w7+oObgjnb8tqGMEniWpZYL2FWIzxFgdsEr
1JE5C8QMMMXxuvE+PrmfiKmm7R9yg1G86V5fQkIECED7BBAlMtGlCfU7P7+242bg1p64IPS65GEU
wpPtLKtakoYs1q130Z6MUP37XFGRgDDSeeWqW4Z2U+sD3PqjZBxsB0JtC5Hi6PjL024EJM/D9pEd
wwXLmGdLsdtv92DpIXWJ25efBpbQpjdcUGSNBJktnjtILOcqkobw1tFjCLgwHPMY4ah/x0UgW0D9
nmNJA0k84Mk8dannhhwdSim1wXXRNw3UgR8+0U1zS3v0tvm4fan2Jjb0yrgvm0c+UkK6HzQeX/OX
uwMea9OWLkN9oKZJ7zb71txKdFbI/txpq8akVoGCQBR2zwIXbTneEoaXUrsQHGxoy9S5/9mZ6ZsQ
uqVNgIcD4rk1eGUfs7DACONKfaMlwJTwCv/sf78EKeuEQlmxKpgU0kquErqj1EodbVQfxIDeRddk
EAs7MOHo7sdgX0Iyj4WbDy0JZpuL23D1RjjlvQsf7nDRqmlXZvOqELOIAFAzCEKLAsDvEUcLnbjO
lpGJ7WKwuUNWBgperpbCKLsFEqk2g6nlhfLs0Yc5gleRXx0oYE/kau8MtRT9xHiEItXjN6RSaeoJ
2+w4FGydmqr6u7fTag+twvveqIMCCpmDl0cACgoDjRHsDjxw8zibAEkedDAWIqlFlMpbDiOgDLuB
9FyxPWWFWoihpF+5EM75BmIw8T5EQp5+a82kkAp7nmA2w2jjtEId0OHUUG4dQCScg4IW7H6l1/2d
dRqREiLR42TXVdAlHg1KnhoQP2PceaoBGiC3CiEgyQbBwleXX9BdgLOR/xjojqPvUjyMy5ROwH5/
fq49mWkylnElwz6iyj0gbRrtd2KXltVvTWXomxh+EUnXwrUrJHp4zGXOAqRunJVQBCMnIdKqit3l
cUmrvPY6+E2SSMwUxHMhn+KHKeMlsiCya8yRbCdWpDNQnMPSI6/Tl9+S3SZ9uvBRB3Jcq90oHsgD
WSFpEnpddOlOKQAGXCKOVjNuApy+uKB/654eIaiNRob7jeOUmzp4o2DPg+fc7qKJj/MsG09ApGyG
+r8cTZWfLzEOoQXRkU6MnJLAk9wyc1SLn3EzIvvyDETDCg6nxYfh1iBnEOTgoekpVPXb76biPYIH
vl5bxImdEZNWUX7kDS/C5024veVSfK6Y5zBZrUF5w7S5JxOKgzZLnbAFpFreM7FofplmWZvoVcde
hgLjz0FPZfRHvWqoZGARKgcukSmYYS7vNVl3MU7DEseyDPbRmj3eAOEQt8SzXo/53IyYJqCF9fHI
eGlIgR09GE61tntCdu6bGPUzmifZhyLfnb9ql0SYdbmpd+9O6LiBcoWV32b64CI/RCOqg9cc50yy
MwMiODoZkJ2N+sMySFvalEUKu+WEaiXDKTN/Zjw/qUwPExi35IJZCkYUxSMdbGEyvVSyclbQhSzV
70pmblPMG5hGrw628NSxma1JtM5O3NlNECGYAy+UjZuB0Na0S07b0qrGsRmh+jx/4K6EE7YDCDS8
HoUBu1lcGzXoYjggRg5ZfDnfEjSVJUl9ZUjHWXKtugDDZwjR/qI2wnFFFTrMixgAlIpxM/SnkTmx
bhooZQHC2RzTejE3GsbfsZlyVWmaQpwZFLeAggbIeaHce5C/2Kjv8wBUduriMymS1wMp+OaZ+LIA
zFt8UVav7RNGZHW9q+JQPd6oRRB/rfS7DS1ArVXx42gKEJZZDEcTBw0jmATrGl4mIUo+JJNy7xjB
21MTl5/ZAr4gCLDjy8SKyrHWGrVWoK0ttGswVCGs7cDvf+wtLXWGRiNL92rRHZWIfn9AaaYceFMk
HbRt92YTWXcfcdrFuaVnVX/CfX0VJVD5rfVxh1xd4bYOrxHbN52SUi7A9B+g8A8H0y+U+KecfG8O
lcE3xYyc5QjWUcFZCemxolbMj//8MveqRLdlxquEw/vsv7roYKZaLqDMcqUgFsbygTrhKJxJsYFw
xCXG6EqB0Ft6XjiS/DM5uK9TLw24xQYpp68qXgy3dc7LYZnB0khqKiixjFRBuog/zkb1Da1r1A9R
RFxo/W8EhIS1uE42d/u/7jWo9tNfADuO9nPy3e6R5ZN19GVFpcvrv6dB9hWONh4sCKULIzibdVM1
TxdoyGFr4ukhs7oiT6+QbAgS2NwIh/0sE4cb9AYZlIvxSiuzMBR7vLkxZ2/MSCYPRz+7ve30bbtT
c87qQE2lgECTi8ZsK3Yw4RrO/i/kzCk5sQGA+hB2A1fb6rG3iZA9JHCS4ugcI9OPdkUuAXd+/TgK
VwjRt4pThTYiSQSRp6EGiU2FHwR/DRO2HULjcAvLzsNnYKd+QNQEl21sjVvEsJFbAjf591d5tlsr
fIGSkDY3jkb1tLAX42EvcVnW87ukJCWdNRSUI9146fg1XJvBlbHFW1NFMZ8G5nn+IXxpnC5Rd9Hu
K6kafSI/f3J/NxofJ32SSho0zO+dlv+nGjQ7R6/gBv1X/Ujo2HG0bcRy02DcZdNyJZ3T6H2zFQse
rynMFMHAcNnipPzR6EJpD6mLGggtTcT/GrIoqkIk5eZKd4fsfj6c98ce3NbWvOd5UjviuOmnolUI
aACeZh41WKzGQBKkm+SfSCVzdzj5SbZVq0sZF2BEtqsq3X5aWThPHzE9Q1x65VuofkT1tXHKvsdC
QJY3685x0q0LyxUi84NP/SQgaaXjk2U9W88ine6aEJ2Lk68xLkzLHZVS9jmooYUxfa6HZrfzfSqq
CKizkdpEVDGhJCcfRYdafKWrk8rPEdMM70p3TPaZy2t6yuvJbP5VuOUoOcT0AGgcBN9wzBE/1PHz
BEahktPcdNVgeWJBc4tliV5WSt4FceUBakLszCdJsITB+KO+EnVdMmHwY+xqEzz3iHw6wmVCFFhd
GmJ1P/fHCIDHrRU2LzI2wrDW2RXIRMAd9yLSon5O6NZgbSIkc0UelZopQkAqyo0bSb7UgiTNUd8p
vpj8D7kpcaCHoZ+BrFFh/aK7eObMxTUMKcEt2Jg1Gz5c1F9CozJpqImi+OzkjZPMcEWFOp6hXfSd
TMZ9K0i2KDKp8vEKQgWuxuVk01+xFrTnF6Hk8fR0/OfdQE0w9T+fCIiwVd4TDiCgLxcGvjl1vs24
KPkktjdIKnvfkHrLQZLSXPoL3zP6XfuHRMBshUxcrLOMXdV1tozRYBiIW++OziCupeJn7N0rVFK/
gF0gmPhIEHfeJ709Zloi8TZ9ZnuMSGHSwbLq72LStFrHwPNNWVhPU8cAH3zIHSJwT/c39/wY0gDH
/tZX3eo23oFhkweviF5+y4M0nixKpv7B8un+oa9cvi4vkfOL+egfXbIhXr2Q1EvXL8f9KavFfoPr
NA60l0ymsxwZ6S53fq0uRXqgCE6JCfNPfGvx5YcwEqFy+uH1TO//M3C9G3wWLhpJlWor3XD4s+xx
8gzRHQ2YvXsBh7B9PdH7P5qIw2bQAgl2lvcww5xyvXFgBxILB2VYChozaLF/CGwr3185ae3TDnp+
67aYP1BA3tmhIYvznCZUo3ZLhgM1fWWGoah4RmWhTErpCsHTf7E5zMB6goQUIJJKUpmUgQJqKZ//
wEfIKobvDf/vjSzwQMFJUqS7JbFzSGZ37bCUMykbZlBEhGV0vgBjX5zwUWzJ8xCvvYq4D49dC0cU
Mi4aV3/uaJRvYFHoBa/DbbwLA+o5Mq0QCpjI+aH3xr97DTvSXdfAOCD++kRe8H8+s6JBzjL4LJMK
PCFcJH2zevl3MNYqL4hMbF6kuAmru7f6kVln1BEeF8Agl7NMkjgj7lsWw2fH7+7vv1abkXtoVRSW
iUKmHk1iwQdiLixFYGlgeLPe8aMuB5/Xdp331zzxn8X53qXGZba+OfuM0o4HiOVFMlzG4oBF2mik
/8Gbb+jwrNvh8uWoQgogJZ68D0zwSm2rcSP+UvJHnlfmYSYc1/xeNe3YyDZKsHoFtKRBpKTYFpkH
iy5GOZo58VBA27xka3mhvGiGxAHKWtYDpQOIDPJKBkLKJefwU7a1WgQxpAaNccvG3iiq2s+Y/xhy
By4IkyeI7lATx/6CoR1nNEVvsfiaMJA6XyPydp6lSQU9OgOUQlWx9QVvlYNKZcgFi/wwijygJens
7ndsvQWAhWyfBSXr9C5qi6x+3yLKqtcDuAcGSP3xQ33XAkAxtyHOgd/3g7D5eLAsnEVydA75b02E
LIk32O8ILU2XhbuEyjICtZtxSyOSK9L3wRJegWG9nzl5Cg3NhFD3J4fjj6/EBrUqcQ/esxXYJxTx
Tm48PSc7gQimPrkEa3UkhGQ+zzYHAwLaIqNtGi4THPXdzalgHBBESaRx189psFqav45GFd7T6DpQ
W6RxxNT8nudBlfxC4z/qED2ct2qjyoZojofW19k2s+iDu5vHeZ2BjgWBwAZcfL2gQolAmbK9NKdi
Kfnc62liOs9qctH9Y1ri1TeJ+gqjW+h+NjiTzLmtReJBR5zlcmWr8ep5NOJgbNACEw43xlDOnDw1
z2AIEZ9Iia1g/ADnkx1Vu/IpnEDZfMug6G+OgA17TY5VFYSJD0ZRb3G/eyebEZvixQD/8GRA46Gu
5J/gNC4IJaMYTN/UiuaoOB9YYXVBGj83OZQqU+oU+JrnGzJhQfd0i5rikp0SXv5I11hvTNZkU6eo
OszLDhhcuM6wImDIaSyz/nZqOqS5FsPwuumPxrfU0Q2nHQcASPObM/1VNBen+VMhikKoc30GarhZ
BfNpJNjo64ai9PcMgM9t+6y+l1nnu0aJ6QOXMSlfVoY8JtrSIZaOp/2ld017kPHCS/doSJAQSFES
LiTS6LFsdLCjkBN77PgrHW7f6Gf9XFI7kqepHM+MyvwBTXeR+kOtsU0QNKFP+f1MAsgirh+WoMUv
HdgDQu4ZYvNqVyC2+cnUpNQwHfRoNUqpLqWS8t6ui35s6c3h22I7wWwhcILuKX8uGmd49Axur86t
xOOmcl8rgKPVcsYpI6F/tBPxnKNcDjExHnYUvGAQfkTzYuG9YaEJtSRNghcbx7zl45e27f6XNCrH
cW1oMz5ntx3fUNaDK5YG1DuL0leQJLyTs2IIYaaAYzWAHtO574v/2xNekC6vaXr1o9wgLr+xdzvz
ixJ/BxB+6rGvQmNH5LuQZPkyMqk/ZtKEtJf/b9XPbdG53FjLhZs4YsrXEpQDHa2dVT55i0BdYAMx
4xjrB52W3LTAwd4YNQ1XiJL3L+OI+z/PAoy80sMGGQ4awKMqBk8ZCz2NztIBWpYvt3F/JdPSrPxs
YiuJwnuICFyc5JQm3//gjpzF9anYmk4UgtaXSS+TkuJVJLN47x5zZCYl8BSDJAGUVYD5FkNi1Ld9
HfX8/H/5ds2FJNJwIJ7Dkb8avwU7hEAdqq+GBlMdEjOja6bKS2Kxo0teWvlCWMEyQbJHM5lsvBP/
0gNjmMQykBQQfywjvmJ23CMX80sQT9KHk065cPGPAvcs84WrBpYfdZDJCAYYXo+vTo0p+xcV1JJH
zzJQEjPThMQgU1mdtm6JE6xTu+pvYL5C9EIHKKRKFsdjUR80PbNfUZQwDc40/LowLyaMTaBgcLEx
cvlcTnrs6N/tr85zEydq3Fi8Qgq0a1MzX+JCzkB094pTz+YtHQxZ+zWW9nABpRGZzlrmkX9xBqpF
+8IVd62qVJI23eVGj6T/RL1JD2Wr9MllG9KZpmnPPHUvKewlDvTZApLKut4E+DV63wH2ZQTuzIux
z+9AR+04sVKzxWyAPnCCKq7bMkvRQ11ubsJ8E43Z5J1VyKJgxw/NLODPc53UoFwStIH9chRZS5Dt
W736Ccqa7jpoHHHRy9/1gU7Mu6EDHp5LUGjflh6TBRaW9z78IqV9YwB5xDKJsOiSFUf7eRnWG93K
JCulsoGzPkX+LcDxv1dnf++8CRNmktpZ2B5S0FvuXuxYtN1Y7yHLz7BS9V7D42XkWHIwHmb+T/05
Q0Rvrso4f0zjDvoRHYrkWZzonJ7aSAGPTcDPb6QoMhJbrsfL4ChNBHmipfsUrcXo0S13TELHgbgh
kce56+BYKEjc6r4vdvi4o8syPjK8GlZ+k1cBwQbBdpTHqiPGL7knYDFwyOcqrDiZ6/rYp4lzCKBD
f+u/0XcPNMrZoJTBs6aQOnA/tEW/2MJ8+nR6XYs36F5h0rZZEx5GNQIh2Rc8khJsAWmNup+YFfel
0oC9zdWwiuC+P/LC59MOe37Wdqqo0hP24Sd6/+ypIdhft5aIjCN8m35oa0ObRNPtSsi5SYYN30Fv
A/PXnkgmOpa67h9/VJzJiteB1atunk7eXw+EffXABN26Rmv4dwP9WxrsOTKqFw0NalM0HttVZomk
/TWnz/R9Q5K+VM7ALpQbnMl/BhB3Ptyf/N29ZAoPFJiLyPkmEivhxPEbfYvBUQWkn6qibTRIaLT6
AtA9wyGCW8Xug00P7+djVimorN10vOXV4byj4mfdSjLkA09DwEtVsj/VblA8gP7uPzYS2tU4fuKR
3QVBQfxxhEhug7qXZbSH/8z87xMDNsHG+I0j7tFO81KPH8Mp7WFrS3XE43NHO6cklxSAbUVwlBjd
bXY5wxS9STlgJPyujdhR6W+G5nX5X9KqpAbNTQn72lzIyip6zP6UP4MgpHx8gKHSJRkdpPAmFxrq
3sZtUJLds20pk4AknkzhANo+DkEA7PSD+W5G4mbVYTgoX8Str0nDvb9cx0OTEChFev81wtKib+Wv
jZPH9FQ1y7De/aU+wuwj5PuWqA6TbtqVRFM8iI0V+7Q9SaEQUo5lzKBm37qhwtuXzJBjhK6uEb8C
CF6YbR2s6FVxkDeRZ/mPt1Sn0bcvpj1OvPIaWWwG0WYcohduB4LQXzb6rc0CCAQEPGezKOBjSMhv
ng4/l+6G9ZrlU5mXTukiXXDm2wU6l1bQhTzGNJlJGezNNwxFEf3OB/bzC7vG0AQgKKt+GjjyJQIx
GpFAXYUO+SocliIutBXIQcvWpqpNNhI82wJuoYc+7JOT9OrZP+DmTgaOqvC3oYlbKpnfnVjNtPXh
Eb1iVo2tGAplfXQZE7ZlbQFgAogDKUTQFerQ4YzWnnFCc8TF2AQ6kM6VtG0oteHACCkGEXZ4mB1U
aeHXZfpZ1AHFFE/Ckv/iCyzj1GjsO6/ZMVe6m9w+I6FTfKqTiW7YCKRt+l2sfvl1Zx6YUqc+djzv
Uvu3QvtbCppPbi92l2YkhgkAfjsZ/zKxnNaravrdfeHPdXbvoTCEqeXTX6mw4oct8r5+qXnOUe5P
m6Zpde12IOQMH7/P0QitRYSKVBHUne4+d5n8+9eAjnyXUfyNb3w0JA/LbFIm6JXq71jG02QrM4aY
8KtJXJKAqK4TnLfme0ZUOpK1W6tNhWlgjM7MaJpZH1c5/hhsr48B1dixqbYC5ZPpgFY7UuCBxA7h
B9fxv0niip/YVKOXQkE1qGQYCzarcLzXVcu8M3Pi7ad+PyIxeQnm/T1V5OMwKPjmdQGHpmkvT3Kx
1SRj7KHPEIFPwr4bhoNP06ee9eSo6KjYlC4E2SNq6mM4ERXv57gPoKo0VEE7MLK3r2PA4gW5LqIC
BUB9Z0NvZnqzntKSUuRjwvLVusi8w9/c8Azyuvm8WKhgLiYbM5PWY8xA3h4M5Er+YpjDHnVykmYk
oUhqYUHwXyxGMzMdtRCc2QEdCpGo85q+x5oPUjh+/3kEj/uE2BXvko1laBvyxOnmCn6EA4zIbJ47
4rm4F/4oMGhjcyb0nTOReeTnU9gIQUUztarN+0HnIVs8Og8rxKpvRsTF0HrcL9a+q7vuEg33C5j4
xzrMnz/Cn/BEPVzpX9l/jqt83WDXYwy2C2H3NA4EEkufgRnWsPJtDIUjqT+NbRq1MQLwRrmQnsip
sZJUXQm5fpKqA7zDtlBtNlEwytOgjUfi6Yveg+UujzzhqgbYTlZQ10JIXX8gVpogia4PGgklikdf
giV8ywyoWL2kCslPcnjPZmA7aFS/Vw9xb1hH8CqeJ5omDlz5Rrkouxzl8zQw92O/tqXhw6HJRIuU
os1yRvKdUaqd7qwtr3JTCl4f9yMolBFw6OFwwXhYQdeHoJTDfHkyHQT7smXZVs7ilPsPdwazuVbp
bJct9Yg9vGdglgiM9r/w5NAjmoIk4wXPj1Zd/4fGsAOhCEZxGqC1VyjREz6fK7uMO/GSZExXffde
R3qva0TlJiJ6kiFnbOEHuRSf/+jjJybsvQELfpMnNW7qeHL8sqd/0oeMjZu+pIWF5KRZSZs8uEh9
tb4cdEeycYoAm2QoyXb9FLS/6DIEuPEbuM5TtcR7ZUXtp3IaOjXRfK3X75aPt+VtX/XcM55U58np
szMshznXg5cyJJxyCdXpviC4s4m0MkvoEbeZo6zVzC+NouPnEUZ23ZaxQs3O5k4MR2WSXkCsoaiJ
stpOkszy82S8WaiwJBStchYrSnYlG78MQ5su0IG4TRPHmspwjZijTccbe66RsgmPh046JeWbx3E/
RipHIMgkP6Zk7Lqn0jmkcR4grJKig+Gc3Heb+qDBoPsxg0hXIku+0P2AeetmWRYPiUgMHVFOhD4G
xgPOZMDaWm0xQ7O5L62t3GuZ7Ptv1PsWnX3D0NN+O4YoeXuQfGI7SDhs/Wu+RYCsyMoIco+13mct
CxBSCGE2Ju2UjTMOa/6ZCfcEeyIqxPoJdZ1rSEwU0MaV41JjZoCea4NcL8HJth3xz7hUk53KhNZm
VPfgVyajqQFLfejbvWJV6gdAhxHPMHgVSsLholcxD7O2cr3L1HLTIBsG2PpdF+hHrH2SMYGxsw/X
QlVkdVOKOcEubztL6RZXybeNJnvwd31UOcClFhDDx4rq2ii+Y/GfCOhBnfvWbFI7hzFHtVFg6MSQ
nLSfH9qWovrh+hU0Llzr/woGHoZSm0UKza/f1hw9KFkA2tOiZ4pmYx/Zp2GQ4Uuuy4crUYlF7NO6
JOaFfi3r5f1MvzYepPo/Ojsn9kF5yoHezD6SDb+wIdivd+0MRyeEtM3Rvkoehk3FPk/B9p0A3Wrj
TJtMCmhk1lTGkySPRpikqlvAU4ZGheR1BFps/06Bx9xg6PWpKDG0cD+7bc5hhzSCDY9U3d1tTvxD
g1VvSXt9qASDX8VbwgtR9xqzVXKPuG9PWqrWfFFe/LlITj2e3ZZIHo2A+6WgNPSxCd+QGd0kqHO0
3epZuGcqKod0y+5JnVSTXlZ145PZvc3hUFtDLt3T8q9J61GdWl+YRLcdyh+ttOZPGLA2ti1pn7tU
7SlpP6eGgZcuYZa2ygeh6Gz6idIEr0yNvbzmIVhZGpo7BwjfjWRjCXxbe/jDcioTTsGc5j6tjHZ0
M8oBZT2Cmnmui8AnAcMOJUXUEWagyFD1+QtoZhRW7LVLaOd15mvWuY/ZK6wlaMlweqk1/nuBMcon
KN/Y0pvxNNAIVbfaQPrrvn/0D9BIMyuOLorHfTAVvv9sa8BSChfZhQ+4aIuGkQjdXI7IfUYZXq5T
FVhf2OD+JASDNzKr9KzuU7IWaXuuelRhguVaab1Zpfti+nIsWBqqDDuEoF9S9D5te70K7JG4z5HP
ti46HwXs4JVW88E5oG5lI8EDivv34+mmQY7PcFM6MlXWo0uhmYY2+aCwd+sAoqzZ1F2MRD0KWiCA
isM6gAD8qmydAlKrpft5oz9t4nBufNd2x4MuxoyYFHi74tYXMdWGQ9VTQeb3Mj7NmMAGJA0Bsmcq
LBzzmHL7hk+YZGp7v/vR1QGcwU81a3P/iz6mF2S4sGtzITyibrCVbz4ktbz7oknIymyzG1DbYK19
Pho/AuQfu7KgRAFd8RvmeCehTWc12nyuH3yPppRQ8uPSSK79AREZlOIOYR55fnJqHhBUU5KHRtxu
aqFG8AD1VVIau5TPGmIjwbjTTca+Ha9xwspZBqmj9ll9aXTahRXE+NYZgCSIcEcw0MUYqY9Q33qX
rnCLBP3puTumHYN/l5Tr5SwLQtcpRAhREeKYFh0+Sjhh4RIqGrCfeg+3Rznf3vtHaEGpNWkSnVYF
deqxNUJZHZCDJEO8E7LJ1rwxjnq2xT7nWvKBmwRjkDhkqsuuT926r7kF7aVCEnSMnY534gKQ5s03
cDf6q3wZTx1Vyl8QPWlArWaJY33xYDjdNGu+5SRoxLUSDAUC+5sps7ryd4KW5pvzyX+snGrlslOU
MaYiPseJnMRIULxptcUN1P8dA1vc20xueMHFgXMcqaghOGLiftBoO0hoycFoVTS1aZSm4gL/GoVi
6hoWVeRLKbZT17lEH0KfFDnhS0VmS6Q9IX/mlY77DIvibvYhpn5c0OO3cCY3hu/3FLnrZ1HDGJDq
gLZgJ9MmMnIrW3fXF0TXmxWYdclTuLzxmbi6MwJ/iySLNIHYP3ao2qbDdkbLXPlvsxT8wz9wjOcz
6L6veCFtIEFjFIVGbM0LrxtGKZ9U3CwV+izraEuDj9lLk10cr7/lrRFZY1xW70PYdTI1Rv7Fpcmt
7c/bRZ2IO/4GsrPXsQd5xQMR+cvrryE0sRhahkROQJMIRycWhbUg4sIbqlSWup960N8pb5jiu3rj
XtSDL6368StBrF2l1ab8iuFh/Sy60CFmEh5JSOi6mHbBLIU/ZFxwC/v/xYYQmn62HCTub7ADG46m
qJJ9jQJzKmtIqRs9oIe1JkwDRD4sdl3e3Ai5lk6OnwA0G18gRbWMCClINr8rYXcgoiA8VO7M19Ei
V4BHoeDUJgdwzFI+oIO4QxVN6dBzv5Xm+jd/9P0ddvNANFMHvSZwV7vbXhkQpP52hvpHSfd2CQb0
eoMoviOQUJXV5NoTXSW8mJNfnQwTZrlB+JHxVU7W6ZTI4exbPvmRdnMi+upq4gVsAmkbluXGOCjg
/3InuZe6BFt7fs631JmCpdDrZEosbZMEPU52/crxm1GJgSNElAa/iaXZG+svQbhIf+pefatDARkn
IX3H/AiibKdRWjpvEld/2Z/I+UwlAznTp9rMdVVQfgoxQM8V0glu497KCgKCEmbbpbgDcmD6bpEq
kvxg6FTldSGFlqRkcIe52vj8izVm2wXq+89WbRyIVqx7LznH6SvvKYdjyQh+ouqmOenanDzO6EZw
T9D7lVJ+5J+dzY+XhvCm1JuiRQvNDkTemQ49betrIDJMwPWijoTbwos0ZNhO9ad0vcsxZ1XY96d9
FydUUiAZk79DAcS2TgKcal2CJI8OAjB6/tBe6nA/z9j6pwe41ym/uu+p/DZWZU8ilrjReiBwtAXe
8YYyDj+urHDTMMqDUIToglmjDhkfSYZ2djsgxCg6T2AgdeM6p69cEq5bucbJxmo+N8PvD/qruP33
p46s5XpXFZ7lfX+D8TkK7C4cU8dIPXW2RQRphdgec/a/whbVT85r5fl4wQu6csxgtu9Q+tztm6EK
sfJI1OB7WFmpkfqWmD2QfkOp0hGb9eugk7N8SB3WiNPKvBdqlWtNbOj8iBRsQ3taUu/Uy9LdEJaS
7TPWn326e1LpnaWCnSQLLCjCbbQsR8tmsV5L2ZcgMRWb8aJBaghs+kpEDBOVdE8K6HGglTPLGCYz
p+0HR4KXlisBu4cI87oi+8fgBsg+E0VvpG2cQJ4kvGL2zri/DLAj4IfGue9PEmx2TKytDGUn2UD7
HAFp6kwUImuIAX11Gt+1TrPGVjffGPdWPYs86xHEwmlNhELrXaUqqK906hbH0j+DwXq1ObIZYmqQ
kLHE60t9BNVR2ennYQNo2wdSAwtMw1QyHidL/w0XaFno/e+1yqUrQNgkgaiiu6saKxmayhCckxL5
L+YFOtT44kQLYANticn92ldBnEZMZM+sH5qt1cHtr5DOTdQrNM96EZ9fgwXXF5CCKHKzWIRlREAg
XC8msgXHH3Pk2yMKEvl3A89bJRsw1BQLc7CBULJa0IIj7TrXkYM8dk+OSFD2ACqYyQMrUEf/rc6a
ggZ+QpxGtb+SOSswyZv8wYc2eGcLwbTFyWtcrfvBNTSagCvlNvhUMs3Sx0afZdRVCNuRWMaxgaEz
kBkK97NZ9fRtChsgPG5TM5+k14pauAU8QL3cq4ZS0SVS0PehP4PcXSl1ZXZda6Sr0UBonseqlMVn
RQxMBhU76/KtbyoPJTsQQ3H65l96iIZE0FLbvOEbq02g+crbVPoVBOJPkDK5PyDY2jeU2UPI2mFJ
0IpMUBG+iMAPHLfbAeNklg54CrJzffKJHlL58rNNOGy38a7sq3nuTvkYyBpALtX/htlfzs2UFOKe
yeV/u/xr0nIR7Lrf8t1mQ2UzSNg338QkcT8+Pyeq0B3otmnT4qd6wkhfRod5VZ/rwg1glGKvomse
8ZRO0bca9MoultDfg5zgFLFLu18pEExhcSnOtS1o1lErcnFLuciuOWjUKJb9/b6D+3ehqU9H1XdP
EerLUSU/eWjwqwZmSL/zzRKg4Y1/V9zAMbt2x1t2+89yq41T+r0FTTxDF7Kehc822lIrSxYuVnry
FyQSXg4hWdA+ZFRHKFSBFZ1m46+tjx/uZSxSXQCo0Ry68n+91dEESMS5heq4IZeGtKv7H0V+bzi5
umQkR1sAgB3bmghzLyoeJWslKR3IUerDSaU0gn5cGRFboxOpiarhQx/08mjrJ1AEnhx/eyZYI4a4
aT4yRErcFPfLjuhnvHK4qCyoYXwhs5YxRRSv+YLsY6LK2SLHDj1igYlThbjHdjH+5whptjiq1B/w
565uIPGQ0BfYATsqEWLayLoOHJwH0PolBcCGMQ52Awo68LVMwWRmNIVj93JuK9td2tfUENLBlM1G
bP2FBH+ZMisXm50+s4+d6Wk9yAi5+WZnjts4SAhjyKgId7gDDSPQyDItipM1Bzb4JIcU7Z48UJBR
M2C5esFBz521PxaMifugy+kV3mw5VxqFwimn3Ch7RKQDIxZS21TySie0pHkkAp673C9B6bOPMDrG
JZXotF8lC/C+5IraLbhLiJFuGWQiVMSjFW4J2O4w+YZX4RJbGwgGsRIzg9jI/iqiUiNW8f6GdrxJ
ytyIPIw8zYYccrA2/isansPM7uTIhEHGpFXNyQ2HiUN5+8B2KYBcU4fqDt0LCc9e0QiPpC8acnK+
wFva0Auh/t+8k5vvSDW7vJ+Ubz9v6PkX0GdblLhrdmFo6/IeIOTVPqnQOruyKhe8L51I9Ixl8GLj
SwNpFW9iDP1MUM7vPMnvXzFOVa6JgY/fbpp3wF4NDIFCII/EaGtch/415qk5CudW0gguide2d80Z
PstoYoRyQkiV3CjxpnwPOJFGYv0quc8ECkiv4z6uE078lp94NXlUlh06yqFcd9WhA6IXajKhVJD1
DZd+omOHF1ss3mmTaR6t8u6pANiwriM6zRTgmHW849ef1z+7URCO5iBhKuGylHJEPC4BTnto2V05
GoqaCksDFImALfFhekK+hoPlgXJ2r+ac33gyuY+P8Ydi2Lqz8oNqC+jQ7iq8x/0wqkvb/27DjMaa
eqMX+ntASjz2rp4QBBjiI3MbajZkiJoWsqVPUxXtqizZL770ohfM81S4FlEz+JjENM0WY3SouLMP
3YlwrJoSPOw/PyvXM1yDELrdYL32ZfoWQrYyep12NibcdWn4ZDqB9gsBOJ09+lICr+UVFK5rBQuH
R2nlKH68ENzM/w35OjlNfgVGxfrX3POhqY99cTHjZNyZHJIytQo0qgSr9cL6kVH5jf7h+ZT6YW78
SNKF+KZiB6Pdh8HyBE6Soc5nRNqmKLiFHGo+F6WF9fbKmdrIOP+i3nKOxPLb1bRfpP4zUKEJN4Xk
PYP0vPx8hlHdo5oohIqomxlOHLrnvdf6cZh5nW9HIe2vBh1mHZ/9eetrKonBKHUzuY16uN4HHzut
CWwFuITPhsD+VKF5/OAJTKs2m37pn8PtKnZxk+ujbDpk/ciA0ZqnqubN4XCFKbagEiJ531KzkiEX
eK14F4DIqizXk9aRotLf/pOOQ1LtBheRhjpp45PAw2XP0tzaspvxthaCtsV/lUv7x2jkp0F+QVUo
cDyRhR8Q5HFPLJTTXqMTijo2vG6bzejhshlF2GuZ2+LIC8hPSDrZ87OWP+RHhqZ1vqGe2SS6tddL
4mgBfBYOylvClSUe098lz/32Q0+ApanR0GPiCN9Ak25X/VFIRwJv30PaOzEiiYVd2fXuqzJlzNCK
fRJO+aXIx6be79zaYesJWFho2AoKBdpCsLT34dkiXa3XGvHKqfCVdB6wSG0leUJCk2/SSWJ8wQJ7
NSPATuX0KgZv2bXKKyGbmJg7EmAs2/ZwkAffuH60TN+PN8XwLVCcWFzBH7eQLZRq8D0vpEYDY8ZA
7SVbb5TFc/sjrq+5gZnuOMoeBCTN46z5HtLRNK+AoiUb/BmW8v4YX//VJimtV+uIdDOae++uGrZb
gdiUzYCrm3S0JOGLtHQyGI1I6/Gq9zQbGq+bXrjLUpxwuKlA25bOaSJ6yesTgpY66ESktqjkphzs
ElahDcGY0Y9WeEXmQdTQolUs8n/rrB0Dtkvd46ldEubtODqXmsWgvJ8AlWW5O6IxmyPE7nePuu0i
yqarqe752yV4dpeqJYOFIbxgLhufrdgqgfFEGClnHlMvBm+TVMJfcQ5jiQohQHKkY2wxNPOKDdFX
SUUUQqAuRjDYUVOExQkM+gb+Ch4oFi9N71On1gxf8jQDsjofM08baF2w4pZRgzAvnlM8bBWr6zpQ
YP/Yjj4F7siV/iFMbN9pAxB+D3aouB4EC4Rt//FgcYG2YH3HYOkgRz+h1QpK6utH7VqVxL/+2cDi
d0/c/6arFs+sfsmu3BQupvAcxqDeXRy1BkTdcc0SD11wetOIlbWLcyA8CWiyXs3QtgXyUo17hsPN
4J6c2y+3Gl54Q7aL+wA3eVGBKLwWDLu1f6AqIwgF/iCnJhkf8e86UIU6LTSJs2xrcQG1k3GopGMN
1m4yIbG3b1TVhd6eMpaX3AcfkEVYlW1hBan047/uOtegMV2BWiPZ5Kug3cy2bim08eMDCsPsuynn
lL/Df1lfxC/XdmlyNH4M+53kQQpBtRUUCToZfEPKohkrAE4OWcEnMy68EZH0XBYfnyCJ+aaebwyl
yAM+OhpxCU0mqQWuCzZTCsSSl0O+Ve62lLsPdPbDWDtYchOaV19RG2aMXlvocpFpFJ1Y5gegORw9
Z4ijNwtDOgCD3Rbg4F7FW9zLMUbtMF5ZFdSX1rG7SioIWgXTUTKZ0f1WPhYea0xPDwY7y6OkG8T+
75tuyp43wHWN4sJn7FS9dKGUwkKDH/xISeHMuGMIjjimKc8qCSmNADlVG7STJ8alT2AiFMJ57TDx
1NSLIlSOVeWrSbfcBuQtfm8PNHYX8nf0/w7H9eHngtskFdHDyUVrMnFdZc6OOhaQ32WE/8oQSVMu
mua9Z/nHsvUhRJG9XtYcLBz4bazZDurdfdWdtFQhrzJD0mNd97iIla5oOZPi6We0zmVPN0JU/WVm
RDCFadQMaaH0mY9znMrk9pbPb//5rUxPB29s0185VkZ6916Zn52sX260+aGIfqqznYWfmOIFCo3g
+LIZfMvvkmXb7K/ruqFf2YKtIfZQmxhkgorAyNmce0Tyh4bYKhyU8pG8ubsoNa2ecPcXMB+6zxu2
N2nWZlRJU1z6+3OmeBGv03UnxP9/+fL962qjQPdvNn1mrLJ6BdW65NS/4u85QM7abAi2iYb7DsQq
MFvmU1vHVpH2I4CbWkUq21vjmK7eKBrBlwSFiCF53o2gXHNQQc7Ieg81C7W5nJ+jyay3Ntbic1GA
3h48pCxzbC5F/FXZNZBQddHEjoqwZjx246USYUV4bAQ5L2nXF/iiki8xbemv75zaYRH7VQwJBK9C
KAWiVBSXKGFN+VxBcCcbBdxm5ZA6eptIthKupRP4za4CcL8PQOlhL42nQoI1IuML9ge4cUCYm/jg
2ZpTNtOny05HWaRCZITBMarykEbVk0DPIp4XK1jjZUooCdb5qnPHBkkmpE07rztwId3pQl+O9NM6
jtyUEMDQDFgEM1GCA5IkjDrDwW4IJ+5NO3TzktS6cfO6jxbwWkd5OixQaWxc6VJB0QXPumcQt+Q8
Tj55R0oyZ1lr74vjLrVaZxa+nsHoqVbViU/QGFhoTVH2SPhVqUlwc/QE7lsXuPMDzVU1C4ND90qA
WT/MTo5wy+yGoDyTsNc//SnXCJmMH2pTtTjpggyG+iI/HUrKXSweOLkNQL1uu7eTWsmi/C5zF3VA
yx2Lx/jWqcRwBR/zugmWl6LZAIrUGtEdsRGzC0TuWRv3ylxzI9X2gIUh1bY8nV4nNkEMtAxyL0TS
O2hwSUBBK1ely0xq5qoRlUv6gk3gvQbZLTjb8/hCXCb6xT5vGDjSnc1de0ZxNAfF4fl1tt1Yx+4K
SoIG5jl/4tWe4iHiG2JwRlXQL+89fFntY2W2vUbjk2MDw6qT5lrBqtYj+VcggJGKVB95caAv22a5
qSkR79Kqce4I+ct/GXACmp7JCCjPJS5ptd2mapd4IDn80eISO6rOY1R4K+/9wftFrRm85WDRMEuZ
qXyb2JTFNir/qTmjNz4Q3VGo6JlS1rXFKutgnphiTHZ+ONP1a86xS0SsymWu1ACdbckPFPSE5T0F
VXLi2RAxxdKQN/xDB+844PIP6qpqFNRz18B2TIhhtLQunU0lAZNwBLXLHSWH3JrgfammyZUfy5T7
YBjwIg/INJ+ostslkm3xgS3KptvZa6TQ+r0oose+pMUxXLodeog7PHCIF02SjprRrh8XnMldlKFh
bn5JLmZWNlNzQqd+ncpDCTr0GBtUTtcaS8dpF4juwOVbGb/3JPhMQ/mNUoCRkZmRqhp7rK+oQOmk
lnZ698vbePxSx56O2V/uAbxbG0LK5H3bifYfYthmskyYV8FwY/7A/RF5LP3vdS9WyGtCZ5cB7l+R
ii6+u0TSer4PRocycKPLojVh+E/p92N/+NYZsGfpucewI0olH6+A3UvbMb60QpebMHyPL6CH5xM4
Mt03V5f1ut4dGDhRElPIaIParMbAx1sKJmi7OkqfeZkLEmCgPnoJPqcVvr/eey0GalzzmHgUMW3J
v5EdT9xUn7F6VViLmJAypvCzU6HzxxdxMdqLgyRV5IZ4NMNgsiJX7Qae8xwVVdFD2zIHe5iG1053
BOTP4/vCx5IWnY1ifi8uYJ2Nk+PP/QPHr03I6oXW7VIDVPPPvuarxJqL+62s9P+XouiZxq9GXp5J
Z6MgVApnYFvVXN4VOLPSU9go3BuFZZoeclVD2EePGwy3FllOSp6kk4vYwbakJJFIOuEEbWUlezxP
5JaawDnZTFnu5RZ+MStaF7ehqQ2QewRsgcVIMW8bitp3qMez+HHn+6bhMr77HpmSWcMprOvAgHwv
AO4ikl0odFfs194MlAOqbef2out8cWigaduVhFeHrgV7GFkFdeAIHlLNC6pymp61fbzmPojUqR66
jO3jeHcEJk6WG7OAc+OtL4bFXnfUQfpfjsuNVMQ2h961cjiUEOMyfVvWhVLSkY1zupIfuhav0VvY
VcMofAhQU39p+01A+FlMnBpGuN7T61ekY5UgVozoAVhxU3qSCiQt9F5J5CQWVpqAUD104EbgaRu/
nv7pQVEa3Fj+X5pbLwUThLkmtMPQDuBO7prwqq7mV71WCeCfqraoYwVNRumumUmdZt1NnWycpkRe
Wlm5pw2GHUoB7119t3wRiHsQc6WrlxiOWSzRgu1XsGd9Xwi75KpMC4aPfEMhsM181Z+QOf5yx3P4
jSMxa53X7IiCEFR5aTUOSm8hqwX4TW6X7kQIM3HoAY6rxm3G9rKb2mGpSNCwaaT8t0QlLEtewzFV
5vETohYJBkS7zQmcu/vc7nXFbxtwG3dmlwNrU4JDMC0FbHdFBkCMHki0/MvimijJa/OPJJjjGIn3
vbkHvwWXnPj2+h6cCASeqO/ejyLK94gD0S3jcyI4lZGGSMk95zCA55XDRi0VY7G52jlyqCi2zvuR
eRDH+kcxef/ntV4VKSXfyHPklKF9R1qubgcM18Ue1cnQG1Pq5dqNgKpBNRIFfY2SHR+kjYtTyuKm
33Fgx7lKkzC2I7/IddGMTvnqKPmWfrNSIxMOeuYVdmEl+6sMfla97vEmfXXklpWAG2le5dqLp8a6
5vqzzVJk6AIMBBCeGJBcF1TG/Y37XUeQpQ0rMOV92KQ/wnDMT16wC2z3QnqMB2hF9IuKS9vm9ava
Nn4wHQ4SDnhreZ8Ft4W4i5C9LJTuiGfXEB3U1F0es53i/Y9F1aW32ExeMbz5dlvz1a9TLt8EYWJT
1gzQllRIrd0ebsAB4JKIMEwUnKOMlx3BNqf1nYczFgpFHP+cEr7ERfm90WWhpybXZUOSmJLSzXPs
8VQNQ8JmiaBOgsxOf7QqVQMYTRBlOoB4bdowHhz9ystyfn2j3POvMlxxB4eKtz/+MLFtpE2yNeuH
MgFveKnoMvE6CJZmeEuKgeyD5neDQVlXkrvOtQTDn+bzFvcfDiwxB6HRF5urENEpePY6fLUQW0zK
FHZCXmPt1qJLBnNHyeRtyTb+7KkfRJL5MPh2QhF57RPOfRueqavr3j8H+BfTC6/duO2ApTNDSBjs
84QlOhhzPOS7U5EXKmd/cRW92Y72vnDeeKwXzeP99nbIvFY3aQ2OJxHs1D3+/rpm/IMdJYiMw/Dl
Gsn/43gQkx95bOGtY6Y32qjejh6KFB4U4pfb5jP44zy+P7pMgev9/bWvNvpD0f/beYfSMMkuWihk
Uv7I/QujbUFKrjtj1aRuExdqb6HFRNAe92AOvEoJPduHayFYcrQbMPf/ryXqC/SCTcFPfyke6zz2
gRYkRt/cxrWyidxeJvZrMQ3psbBSpVOHsVRztNBSpf+zuqDDchZ851pmrV6TaWNdAwhkbGIm6VqY
S1cDrE4ZOAAeYDrtHgYYg6uNMhT/tjDBnPYiqff0gWwH8dvxd8oxKYmCTIn2y6ZLnm20tOZ3B/FS
YtTmS/oQOHTBPnD3jRpIiuz7EUzu2VIfZDIOZfsObRoar8VLGlBnDaPwFu/b10LgURDkAigHdPto
Evx6POI07BLbTKdvP+mJoAZ+z7zZ/35fmeNWsvFwpaB9M2uGggway5Md4kUSWVU3gz/359d8ocdt
MftNeU08V9r0lYA1b9Sg7mPheqSoajezAqfgxLEViNAZatqG6oBztmm1Y5dOk1tLT9z15mu8notN
cWZbguFRDgVHaezCgxwqR4dYQa92rgIfVOO3CTsFVg7g+JQ5aJZaQA7Vus9N4Yrc3kF+KAtWNdPQ
k4ZbDNKZxXcektnGWjEO/223GLRRFRZ5p1+HARuY9jYcsRIz1ZDko8N8eI9xU8Xudmim8pDZofra
/XPb8kcThQhPI9+z0E5Oc/0GiKbH15C43ui9xDZlnyMoE9Cun1FKgCz2N+Gef8mepsR9BC9bLWa+
NcQtXSanrihkoGDfESBnEP1yiyzTrZC/cUGj+iwD/Y0W2akMJkInKtc1CcPSbdAW24OiADFlfWaI
cMGIeR6O1Zi+sM7/Y6a2p6iOUF2ycIR+jCX9JfS0m8JAzunfnyKUa//mOiYYQKHaYp5IEtr++RS7
67Gqpp5AR3hUexTQ/I+mCmaJswGLiG0Zgiij3wb7sczLhSagBoouqcLDxHrg3eUNtjnj/Qe7aypY
LCpmKuTuNQB55AMSv2Jf8ZWzuyanY9BUIXh1+OxHWLDQJQ9o1AR7XVwdlf+0JTJZHbiLl6KMTMP9
UXFDSBrLPfG0/DYUScmFQyOAsCgqzpb8n213HUeB8nXs7q8X9ah9QgYjtrpRsKHPNblCoov7Ordh
CUbccs5+g+26GNDLnKi+IpIrpParnY16kYMKYlI+kfwSqzQqWjX1wdq+nhBYOwgsTEbaFWahcE7/
plL9SyPVwgaG4Q93eGp+MUyT7QGL4VnMad9x4k5nqmP970k+VSz2cPez1ZalT9hLwx5zBgAsH2vX
ksUgyvM0DfNsWgXTFPIxkBxBpgZ2vaEgTsvTWVUo4SxidAfIKUzqAin3BRRh58awIZWzqOdrdldM
jcD6No7o0qwnyVtYozTHtYnzRJZwnyOyXYVwiS0sEvBSL6gdHIuednnM8Hvay/TM+Y1UODghVj2P
4awVUFlI0jYlomCexmRoiHGqznfgiFDlodSLRzt1EUmDmAmfMMKPW0T5Mp6psyPa/j4qsVMGRd6C
dzFDcDDZ/WFXwP4qgPbUkplM1etKQcTE3fwmPJdBTUbH0RWthc4agphihWEoKqo7OL/0R9ajr15a
T//7aefWJVSXOG9UJVtMmKt0oiWeu5x1gKKQfoOLpZQvsXODjF9pUm54A/09bCB5FNTeTkI+IaIw
ZZBm4cGeNrBNzI5NCsypGuCvhNeS6tkfd8qNzEYCWj9OIZkNnbVmSI5Md1wTdlJGY+FQfW5aGDLR
e2HiwoqkkTCN82mZUHq+UXKhZZWJ3ux/N6Cmb0ahCkJnjifd7AeCDaYRIPtMjHYiH/FN6VR1E8wm
weu4znlKqZqEa9D9kZDK+ZTsH5LuHrJYKfyuKp7fsgxITHNzCoWwdL4/MXjJSmNigNRyQtooEGr4
zjjoFYytuwI7Y4oAL+66hQUvVpU1vCiEhJXpPJ0E9QOpkGUK1umMjWmL9cwfWt6Aa1zp0Xb9ncdg
iEJySiFQDz/uv6ryHe2+Y2bC7nC4WMm7Hw9KUbaV8gXj/H303nwl/lkTzNkr9q/KE9vYheNCyRSI
bF2YOYvpsZ7S9er/+V/yh8GAANS6Pv3I7+Ux+VslWhzUYPPDxkNQbHP9b7DhGLdNaY4hwXnvwUOx
qGCuHsl9Fm1JfuPKxx+YvKwgeeDqJ2u/MSQMXrIJ3iH2S/FVY/SxFNuQLsG2K8uSxae2fNzK3IrP
2BkHSAW3hlBRL62hTGVN+RE3vthTV+mYISABp/HbQNPMJ/fHZ36veEfttAT7WMevpaUc3R1LeKnH
/Jp0qLrbGxqUfkyab1uokAfYvg8J4swnWSl2QmM2WIoKNn3DetAzmKU+18hFu9c3WyEJXwk5RIvd
Qd6obCn0y6fjF4dUkq1C2YwoLXZBH4jiE5V24Ew/W3LifJZKSKxtm0YJho/wwTXC2dRjBkhqxoAF
e7AOFiZNuXtjw/LzrlfIEN8qFwo7zEikn7/mQvJQ31+Apr9nK9n4NK81+2ho5ylfcXl0IvtWZR02
Am4/qJ0Xn82zk8yd5eniAF3T12OZncKF0MCa8aaRLKmA0HPhbfqlXzc1+4sX4OhLYOJRdRCkgu8q
yjpmkClHmgMvrU3WI8XL+zFzPLCO1RirAXz4gG2GFsQfqfqECBxFPOhKqAYkSiJle2QrGCPAdTFQ
0VTy49+CNeHJQH/Rk9qLzwOTSCQNN561BOiz9kF8RqBd3R0qCs+gDjLkk1x5bjByvs4LPwWI8P8n
tpB8YqFmDKb0GtVlOzdlO+iz07fSf0SyKyOlm0Uj8I234AievBp7FfrV6z2LHu068EVEeZmilmKN
f/XTJmWeGZMMW4xYBj/zZXk8ypHLqjbJb8zFw7ES7ecLHkID58bEh7DvbLFoeZRepLL1s27w6VoZ
BQ3wUAWoJjoLmUSrIT6SJRSrAUm6LlVV8cwO9XZAkLdBGQvZS9MB67C/BbJnADbAYh3KvlBxqq2F
ewQiaM+yWG8zgK5g15ALmfC73s308NP9dMW6R++KgM5+Qa+AEg6ST6f0Ol23TSuBaGj/4MhtYgHx
V+f3SHebO3xu1dLaX84yRHBoq/uA5e1EpJBx4rXTxW2sjqzTRUZ6iqUXOGgadukdWJ7dy9c6vXP1
7y0i0pQ1WrK7/XuTJ4hUJLfD4pick1W3pV7A+VlEa02GDXCZAF+dMHILaV8r4YUEEOokgtOtNVzR
/44zrGBZ6aPzX5vrdntYQ/3y0Zycf7QqouymEQzhu0fOThkLg0UWNp2162CCaIF6pzSTTXFQYpyV
INTQLVxjh4MEdwGPya5ElA4XXZ1248QyP3FINWtvHC6LqzRBlQfmy3dODPAmENJi0hyFjrsXydyj
L2Djvnt4SEMjncNrDNVm4d8ZGiHboSn1X7NsTgaP0H6tegLHtrWPlw/4Fl0DEg2oe+Hn6vcM050E
JI0jDQNWnGrzqz2yPbzr/I/tgBoqhLJzFxudcNhxnM5GbvtxnyqQZYjC1poJzuvmhfXiYvqQy+GB
hebLgcabB0n3WHHkttsXU225lsFj46qQHvtfdgmaZxQt/EUiVBRh0lb2y2UbsVhFw0MTnv2q0xd8
73FyUtsZlHA/0p17QtWmZyVyM9xtWjJlYC72m9f9ujya0Ah/GvPsUEC4LJ2eB10eSLnPK4xgLPd9
AZWS0qcswmVXl0r3JAaXx/8JbcAJLevgdJJI5yD0g3juZWv90PpPFCVg0ofq+B4gR+MuW5U0aTQq
fhXzBk5KShHT7n7Nn1+sZYZiM2GfAK4yQurmdvBvBlFovtmv48I1oU4xSSjAQUoZ4WgRU0vcvWkg
KE6oV4sgI/+BwTColBINA1weJSSl6ovhSA94ViC9JifzbZ2hs85moiwGEV5Jn8cDK192ZbDtUGqp
KVKAzDqI4cvive2z39InuSeeFRkwXQN7fGc1Wi7trZFfscIVFooxLd7cyUEu6AVdGTMrKKHC16Eo
0nsyP2a4xlyxgEnig+PxlADk8Ze/AAIkgoKhxFmpv0Nfrza4VLcF1CNctJRFIKsdV+0ThJSQ7lMO
CivuQXNBkW+DVMSO43DpTWZN8G4LA8Zr04GM5diujg0qWZFDbNkHjq9F9z1fK1RZ+CT/s+igbouF
UMMahxCz4eU6plGyixlSffvayWlGw7yv/wNmexmmjFdGkvmkyhQGFeD14wud/pvoyQ+oOG3sCiiU
I3/N+znD++0kE62IUuxJHVuNHrrjDXQ1lSnNijjWcHkSJ+6E4lSJplX95vHQ73xy5YLFTsRP2uU/
+TRgMwBG0+lNiQX4WgI6DDNorTLgK0UBfi2kqM79BBc7yNFCoW1r5O+rZ/nHtTuciqg5E7jHWLeJ
00fYX1wflXWPS+8wZFp5eDqoNIDooXfCz2w1/nfUdmhWz9F3h7NTGk/3zm6UINXH/MmnE4AJT/sb
Yzw4Ra+SgvkDxKMzHA0PZOZo9asNpwcwiV8SDkkA0arN6Rr4K4Q+TcGuVNtL6e4ebYccOda3a7N+
GjCazv0Tp2Wim4AdoVDkkaA8PWZHEHGHxcApj3K8ytlws+gNDPkiGffuhp/EIOsyB1hDkVLrMwej
39m8N9ezXBOgBuLqtFGFI5XnfsS4QXZxO2MYeA5mndVBwoCDh2XTLiIWwCxHDyF27AgWGhNw0jzI
2Ms0KFZsEDwS2OjvI/LbgJRtlTWcy1McrFiCR+rvYWLe8jCD7z6yiAMVoUMSwDf0WElByPeOe9yp
bgTa4TcPp5ZPOgGWfsKkqcnbiiqlKfoTP4SnKir/2cZI5aX+CBXgxYVR8P1+ID9Ya8cb4iFtHpPC
sBjv/adS1Wbg/t4TvQ3valkUwHrfFp/MeGNkqR82kdv3kEBdaarNfonx8yUXxAnmHNJm0u9dWf0+
TJmUekkE9Lm+QtWi2pO5YKY06crLddvy6CTbad702s9MgUSEPMdMhzQ5wR0khq+Vq3uhqxO21o+F
gOtlzVKywyEpQlr4jpJXgLjQKc2wTT1EyPZISBLLd2LVnN0R4uPG6Q7RhxduKHAZs7tc5rs9/EDn
2fUYryw1CVB1/V2KGa60Vs/P3+4999+cupuCHBwDtJ0ml4gvzBdVZU/HWkcJlPCSGc5YNaUnrz64
//qf9yTD+4HlSlogpg4XSKV1K9bWQeHGiO9gUrNiqSIkJNxlnnpEXdfmWApUMxo6QZ2uiNdYIkeS
APo4597EbVAGEEvLdxcyYT5BsToJZOJKwQm79oaemO45UIMABLF+DNw9dmwQunODGBl4F8X4Q6yr
1qgFq9xvAsCNT4wTWGKs5psIyO/WYCF6A5WAL0BFIcwcalt7a+PjL1oW9i8BRwq0EK2bmvcWoyUI
F2IKb1lt0fsTVqDkRkAuHgegPYwE0tO6hbpZ4ZqJlPg+989sselU54oGaB88yLO17UfrspRqeS3S
hR56Q1QyqRXhiyjHbTYKBCKU/h8tciIlVOQe5q7VaFuj8d4/70+x6IfZDyRJZpfJsB62ihnb+vbU
BP5kM4+yIBjYwfWIVIz8wx0dL5+og0/NnwriWAUh/9Qj1CBZVL6ZSERZ8ITj47CdTdaZfwHwlU0d
LIjggHwBUoDOZGRrK0BVXswnB5ziMO9FVxya0YFmRkOid1Enusa8qAvunMyagu+v91x+RHLBLaGI
iWI0GMvk367nv+KxY6cfs0MU7gWllGevK3GV0tMVBp1sTulyRZZE8dQcNKN6EtD+aJyNYKTqyujI
vhdRaVc7mtL+fL8LTnE7RBdt+S+86/prXhnK/zTRHsJ4xbmCw68IO+TI+UTbR0QjpwOnAU+ZToos
mP/oPOM3roMymjFw5NX/L7R7T7r2nmbhzAe8c/rD5rjWAQ//VIejKxlH0byj2JSLxdaBinUpx6NC
Ke+lisNGdEuZcvIDQHUQXo6HDCY9tgqS7H5U1kHoSPp0q0JDg/H99okdyTQp4F2VxUlmSLLawqLD
DhJhd3L9bYSG7hM1gI7BJdItpnVZpwckBOGs6bX5n0re5U9FhQ4Y3F5C6oYe7YwKfeAW+0X4H83G
FVTtQnhnbsOGqrE1qc61hpqFZRN2OmeO9zHHArcd4R73ywzdEahZykAZaMx9CAkTkczV499TRE+w
ZIW8cJ3EszVgQ2cVbtnGtuHzOqYQdKX4LP6vptZ2CegBuKpJttSF98Zebk+Jna0gYj9QQKpUriio
x7rDDeOQ11ghJr8pmLtqP9vyFNzTSjPEWBnOQSqLKRwDfWzI+IJAS/pV4n3RTtK8TwKwdmelsCp5
BsCRbpoIGTg0W2BolAxxM89K7L4lIXgAjOtxpppLw9SvOeTKLPnM0U78m+Hae+uJz4zfnzG3CdpD
Mg3vxmvmLJ5YKhC/iYE1pZnZA9dd3zIgG+Iy3fHaWplQVv6PWoKlQWuoJybqEbV3sjJU15TK3DK8
l/sWMyr8VabB7FoMK5st4CcwUSmYr0rt/+RROGjuk8uPu5YZqgp9XN725RjFMUehboV0hnpuqLHZ
MA40N8BovfIU7FwfSy6bwF5280Z5sTG55voFVuU3Xau1Vo8rGkCS4EexPPXZzY4NWafIv0OfjAOJ
2L8YASn5uq/bw/GAZvMVBVwyoV/V/6Trztrm11CCxFqthxH74lM/+rFuIyHcir8tf+v0/Jjd8UH2
3U6Gjzmia5vOj/K2OA1B8Ju7YcEt1Fw9OZe0KjrX+dgtBdEL0+9gfZCcZunK4nwPWgSR78Ae0xqW
riO3lbbe7eaUFBIRGsQbZ8un5H+B83Jff2U5imFEx6O8xHP8vPnVKEDex9UlO3SOJsgZ6jbh1PdF
P+/mGOgRYPxYoCH48Kjexe+LsX7iA/LgG3tHG0mCMGKIKDSZ7aDaLgvO4gxAwDSm6pzm7dd6M+Zn
JLtnlcPv5XK7fwjl4t/u7JFkrMTvKv4V+7NfsxpoYOjrS6bscaeS7IvjdxUzt7a4f8dMcOW9dBv6
FW4HJb+6La6PnUtLjNaOsMHibwdoqVXgH1Z7AiMNOsjYkLKcRGk8cV4bA8dmYR2Aa0lMUe356FUZ
S/VzWmOz6DIYOr8Cig9szRvK/HG18NRJArtmL8J6piMW8PM9bA0NIFgKEg5aeDkhAl8T6AL/xgSY
p0nykpuuF4PxNnrQ8d6nDcNzt1nIsKnJS+5PVMg3qWbAwmKh44R6teCKwh2ZjE5NP6E2Sx9NkSfT
TMij2FIfLP42YRUTOaQm25mXucGuekikF6lRC9bvZytY5FTAoOzN/6RK9yWJyQGNZkFymrbhkcyx
lkTAzyyGSN1B0IwXt1qGx8ylFOOxMmLA/Kjvzqt7A2Ed4s3QpNHCVdpDhfSRw5dT8/lwqDCA89ND
GyyLE/85IiN0vwoZvc9rFqNe9LAdO63dN+3D4EcrH19glecSi6d1uTMBhvD/37Q03NOtJsozY9Pf
01DRO1BQKkMPBKvLapa6waQqB7zTMhAPsLHIL+tL9CA5v1w5+yDgToeD5L2FY7EYH0esNmLoAbUU
Tm7THexvSOOW+MtU/kajhlH8BLK6aD3h1emxcf+j4kPpNaaVIfQX0ESbsmQa6Y3bdl0Bc4K6I8WG
EjeJP7iNL27ownZLCOsEAgHF2C2cj+eZf69Oj96U/2PlQL3m2UjCpdibvlX5KenAE2eL8mYwwhXE
p8GuQ6zBu4AGqvgn0zZ9/uHX7jndqUStVBs4zBxS3MDMNWjyJUCN8+H9NOw8QbItswKzWnEgiQaU
thLCZa1GmuFxnOHETZZBPqweKpDGtGdOj8pcatwE7T0a9wEUXQKWMyhndbCyELdYCPCoaF4bW4qy
o9nOCNj4oDQWpQyk1soaN06xpVrcGyLSIvWe+g5/VcuoOlfcis8zU2eMgGy8ZrX0KH46wnE8mPi1
5YJ8AYIslCicMD3e0b4n0TcsFOZODEoqm0PrUuPyRHYRabfKa/kFBS0nQ5+McNukWovUsr1ol0uu
zvAl8eoYMFoZtcK34lE681Mt266lZ28sFWwY5ScfNjBxN2vOFY0i70gBtkkdA+ntfuvJMHVcDutW
Xx6AFPaP8nybFTAouuo+A7GD85O/nEkbEVE2tL4yjVMn4YwM7lEmB1AEwN74YpnLJyCRjlabnesu
Lb+2kMUw22Fz29DAP9f5ito6Y1GD/uE5RVO6SetAmp1VTMF0goQgCYrChZQ/0CKfw3xqnXATHyyr
D9Jl/7WfQOHjeUVhi88wudDPBf7De7iYTn7vqYeBrsxOYjy7e6+A5IWxHIt8AfiysiBJKmxJfwQh
nWx8QSVzBZ1LlnfDdE8o2hIuyNaHiLrLxpjRurPhLvejBs0DEA6QLSyuTM5OcT1Y3ctSaL9yUWGG
BruRo2+rDoC2+1MFNqg0WT9vIRGzhGPsTJE/ZA5RYfry4sZe+S6slYoNssnBV7TdvIwoyVWpCxHN
5weDciGvtqrWnwdzx/swqSuELL/f0FReRog2b3k2dJvhpCt3p85by1E21TZe/AoIiJ7Y7/mRSTCH
qHDp9LWcvw1uxGSSoluRvbCdRN9yVMEyFCFRdBJNCZogwkgp6C5ua25TpgVSDVhhnSOiWpZsV5mp
CiTPegp/ng8LnCK0jXpO5p/tFGWCZZCkDCej6UgN3CxQDvZfHQGtsdxsxLTeYNZstOvbGojNXCL1
4gXxLTqjFFMO23CsTn3HHbR9QtxPcONlWkE+QxtP4aV8R/3UziqxkGMWSVRLU3eIL2WbAx3E0yWt
fQ0jlOe8npEeB2Y6yvr9Lq03tvPvlQBHsXLrPB80HGLrWyZt7f5xu6oW2S1SsMQjTWcoMG7eJHOQ
GuKpxAwRAOv+T+DgtSrvESr4CKQCwwG0A1gR2lJVIJRHzq+/+x2mSfW+od9pNB3kilvMe4Yr6bW3
Tlx1EzlHDOwE+fiK+XYoVi4SyM8FHwpk8mw5GixsqUFM6LzxJsksMm8Po+12q4mO6SXfjjHU83NS
fgd92FPbGQJIOQ5Cxs7aDbF4ELQo4M9u9rJ1sS8eYlXTvSkXHKpGlUEUJqJgs6Ry0rl1nUyytpSi
dx4SyY8CYwB7SpziIU0OeNLLC5/U3nnMv2yrPwzYgSQQ/AET2V4dvfmhIWNzD/mKyN+uk2otr7ps
zHhwaXZxh8/+SKkI/RQrLEe2ba5OZJbDhpTIHErHlKJgAMEu4ThAeDd1UvGNiFJCwde101MQwIeD
wnc2XifJjwsjRela0MIPuMvoDyolB/nlrFfxolOWCRLiJqUEqEQC8AkCtPFo3js+4WNhUdlPAvP8
PpBE5DmroKC43ZHUy3E6BX40qAf97Z/wyDnT0Fk3wqvCczIXz7dgQZQViKp7VrAJ1vAUxhCb3LVW
EWFPcrJdPsWxJlKb3L9JYxfgurD0E201jgTjrAKbL4nuqXN9wHU2IMJWJ65fpudnioJCtAFno7E5
m1ZezQUnlNeaHkOG/Oj5R35/AIZ9ZTIKApeBg/U7UaQHrtNdrJzCbhpnjEcY840TRxhwuDDaeu53
HNcDIa7cp9xuReuY34eZyNn0Pg90CefjMNYjyEFE+cOC8mX5scsgterGVH3Y3low22Mmqqoh985A
VoF+7fz50x3h+oNtygmlPJJeXfVZ0Oli/CahEfcicLZfyGGMMtyL9pB2MHphhkjwqbkJTKCLFkCA
veufLaDsr66nWujr9XtlRV7rTVJWTgGRCmE1pZ9kjuBr8MaPx+jD3RtfuVfwzGIYkDRz66Vk5JMN
9iyDo6kqpo3atI0nGWgIeeqlx+rPKRth83irpEIx0wm0WrJDVASU7EBL8PvphubuI3g+a1GN0rlZ
h6Opjis64UfM8IX08rMhVAcCwc6bkAfcGWB4ZlgNPXVjsZoSNcend0Tk/q2ryLZsn6JHrBmy6lnc
hZys2nu7Eki5rg+P/WolGcaP4enVGRVBg4Nyp2owtVjAHF2bt+zaZixkgIA3Ngv3LAiCoVwf1Ynv
linWv+hqmpgvgT/gQHpDx0fs5juj2iFcrsOleuL8qTRdiKi8jjOaA8ZHVaH7khd33dh3tM+g6lmG
Gp6/xvGPo7Akh6DbZeyr8skDI30WeGUVTZf8YP1K2OzUHUDHc+ewRybuC/SwHTcohm5dDVMvkx50
lNDgqq821bVSvdhpVK3L4Xv8cEFrBlFNH+wn+dZSNC2aJTEju1l19ejGsWhia96eoSTFB6cLglfm
gn1XFIAg4ckTEv1kJVs/azUaB8b6ZZhKHGz7vnH53Yf1LOIj5OaYXVgXsaZqjWwFpMsc1/JPIhnB
/uS15fDQd+VcrVva02uNucjZF9UnTyEtQj025yl04mJg5S9gzWPOrvLDsUH3Cc3060AUHTJdq1Ub
bra5oRbByhK+TRAP3nkRjlNBzFB9KDOKOoF2Ic4lFPmtc5oxaqhUAwYxxqIUa6YmcqWfZBuGI++6
PRhibmmxIjK5MfNcr4vXPFUTzy5FYwQbVWlQx9t9c5BLaD++is8yrjiN0tzPDlXPVnwOS2/0UA5o
Q5MgEV+QXNe2wGnBjmsjNT4OHUgtEEDVsvV3nuHfZN9bw8spPaZeA+Vr0s1FhxwY9aeZZ4SUJVHJ
7pH3lq5FS2sNJuSD7YpK0jS23mROv26XyMeqbsBu6EzP5K+no+aj+9m6Qwgb2sS8S3sllRLbTsAL
6bAtAWsdP+ovG32Zbtx41looOJxlu0PfNSKm05nW+Pclt0ew7U0rs8QRPlZQKvVG3WzKVrErU6BL
dqNVpNfofPpICpy9fLpZHlxlex48C4pNG0rCLtrCZaIy86qG2klr/fc/hD1nGexSwGNjiDo/aES5
aHWr8isH4TDW2MSO0l6fSHKcEYfbF864Jzoen6mStG6pIotvUG9smuv6d6Nd8cK6DPsXpCz2WIJc
LOEuO3ffrVJODzQMpf/NUTHaZkjsiMfClnsXfji30nLkcEog1MIwFwhN5N+MuieT+UuVqqeAO6L9
wxPdT3doWPnSJrltRYL2Q2WmmdCwPC5F0cvALWzPhbyZGQCf6UwMhQ+JMBF6byt1uGa3sRjop+ll
oXrh9XOeCqbDKZ8+jiF0YZ8Afp6k4EtW7soj/4P/M5ja64L218YrYsDTf7WYMLw6AtLyaJ/uXO8V
o17ZQi/+goMwHha/9z1+jGpd1QzbQqCdyfmNkhMTXi1cMRv2SuoeOcFjPPk4Dei0hSceuk3TOeGW
Eu4V7Ibv8sMvSb0cbZNrkXj7D6hY67evBLqtuod1ZhfBq4k5ZZ1x00bdFvXqT1f/1f1wlUw2haZ4
VvYzaoUcluJ7P/hG++pyNwiTqSO8CXOpkFWJ9AOR1w4LGstwqqFDL3x1Z12UGVauVwnP2qG4lpPI
+0gSi/gJC18apl+y8FVVdftyApCc9rE6pR+w1AP5aejUkb9zk8O5ad2zvk0fUTIoRNoedd3ba0vK
2ZZ9QSMqywfnwBZWTwPxl4q2H7mUH9KKRKv499/+tfLDOBLhMW3gAFL9UgI192GmuwJq4Dh4s022
Mckyjtcc7wQ1MeEMuqX4zg6OJtutveLpuH+fnQInQ4FGTFjqB5+ChMXBNaUtMApuURJqlQDI4LF/
9L5sW/BuOp6W4FRudIta9xXHZRw2pno+UX44APY4xJaySmgvvpFNBnH59mSkTEIQZ7ndRGEfG20b
jdKGZ2qTbdOVvOe3JDs/6Xi7/29bcthUwraIHytrth+sebxvWX2gzZzGJZpAYjM/IdNTt97tSASW
8uZ7PR4cgIsD6PaYuhwKq5bbCm4alFpJ5CvUEiWceLORsLteLxOh7HDloIwW65K8z1IDYx8Vhmm9
q1f/1mgS595lhXM/5ViUib6of7FBBzmqEXITpNzthq6ME+x0lgb8+fE+FAuhUc/HY2RPiFhnN1wk
VZRzIMhGSr9cHFKdVT1aC+ddnHcRAVyvDcR//KlX2YrhbmjWO2j44qtvzGxqeQjG6+kAgbCyxXIE
bENG+mu68F03kljz3esmq9P7LNVKahIzmiD1OU46lGaMEXKFM3Tak6rrhggblcMibVtv1iTp6Eiu
MBsWZUKZlyYtJB8hNFqEU96AmiRKgti06fzBwGxNV5RmsS5zMJ2XlAXP/IREeeNVl2ixMeUokCna
5dVqrBUv3yRfnLIndbf+/3Zv7An6V2WBo2iKqiLcrOhF9uTDfmbL6V05iNVfTRRUMZV0FZUl+3CG
rruALHYSSabWCnm1IzUALrBNlNwaEhkvN+3D3Iz0GL16AMp24Z0PVxmZxJPtvxSo9fAJ7gY/Lp2g
YKxFq+vRZA0FsOJef0YLGAHcMMSgT8nI2N02IOI/DWeML0Kw7+WqacBMYj5NGTGTwwcid5HQ/1HG
XeBSM0A+0wjkhuZ5C3cyCKlIFb5Ifd0HsdfWE0yiov/zkcym09FYE6FEM7uw7GY5RZ5TU3jddPTF
ie1tQWM+GQAFGjMAYBX5OmTkUEAZx+qwXID+eVy4uYlc3QiPH6cL3rF0wNO98gOjlQux6K121c7u
uvarb5+U0a8lRYqNjfWnoYiw6Ql7s4e9CAADQul8UIr+oQWWlk+mpl2DunK5x2dfPJzDaWQZ6w7t
qGxNeuEbP08tcsBHGAOASMKMlKwuAdwO7JibfB4KT0s7s5OBzjRkVvGcl7VBatEm0bBqpEyJu5JE
Z9e9p3L3Qe56Gx+Bk3FaCRUQ3WCmy409s4St0GBkct1xMhwHFdPbQn6c6RmPrSK7dUumOKTmVV/w
Vg9j0m1dQ4wNMQ5IVxgCTy74rE9HuimWRtJjhnf2yrb4aQRLDMbwwialQAjq40dJEF6VJE9xfxnd
dwkr7qyq8IT4Hg0cjntcdasepV0IWTvWroAZKhGzNFW1SWRt8WQmM2s2aA2hGH3rQP+a7QI9T1mj
bg+rIbVD900uzWHQ5UwONUF1tzf5F3ddzBB74P6LQ1G2YzOCLpZIfB9XioNfDPfATC0sqd7lSbPy
QUo5sI+QWG5RL+nbCD+1lofYTtuQKnt3tTMDWqFCkmOATucrJtj06t1RmU98Cg+sop/q0n20PtMV
Gfmj7XwhENfeDcFozTWE/+cCOEdX52TaOZBtUMczcE4pO+HQs+F2e8GleC0Cs/ZUdGerHeLUk1Jy
rIfbchQ6Be/7u1D5EHxglpPk7tY95/lllJsHr0D5KB6rrX05idjXv8xu4OUWJzwJOzeacHMbOafZ
mdnA0TWt1KQ86ZSt8vfQM++M0lMNPNStS3H0T9mOEHzwhRcVcxJNRqqyxL6ljaWk4PoYVmwKAITo
ODzcIIJlwYJy9+cxOtTQlzu8nj+PY+5f68jo6hA3cVCoYJI8KGdmmMQuoJfxb0ApnPYDi6EIsMdu
kgn13TCdc/XYCsGu6czIzcB0Oe1XvmsvOC4iQT2P//z44aKqNL2u1d52M9P/wTulcnyhV0PVR7g8
eT4rQo2j+hijtnFRHklUeiEwSoD8l+PInPte9DUfOhgvBw3Nhgu1pyqtlpD1QqEyO/xSHPHxEmQr
b1tIBxoqqI0/ob8MUvSCdoi896UG6mg/lTgwsWb2nnWef0LE8wCL18sQMImOw649jssh9J5f8fP6
FujnOH1jK3S8gL1SjMcQoJOPzzH/Sg6k1UFH0wfZYlLJteZZWkEXNJxcw3IM52/FHpB/o4eArwx/
QsCVlymPpiDbM+jgx7BK1x1rqRjpoDKngWd9laqAHyW7FjT+2tKAQrag/DO+IlzjxLKLBzkl3/sh
yD0ea1jg/Y6DRGKaUU/zvzPu4frcGLxYTYKfLwwDOpeIW702pH50pB8s4PoZUAFqYUCZ7jpi7uQe
6+aZM6/AwNupuHzmmgmIt/ISRUiPjZTWcF0nB4r6a4yyQkDjGsLVy0f9hDMRogU/DmtpJIm0p7oE
aHGoM5g/ofdjOObOSCCJg8NDRR8mVkxcZ/TP54mJKcXlhEYw1Xa4U9cr7r+0cgEn+V8eLrSAjJBA
Vc+LPKfCg+P7YEx2QDQ6FbDQn10GhKv/+7v3VKH4BJGRjmw0ZQnb20skgH6ZHf7QAX9x/kjz/eUs
P5oM1yTLqCwTxuGdbxLSKYXR3YmfDU+ApBMJ3Bdq72aIYi21dMEqE+LPSI6z2DIOPdQMXmJwPK5m
00HxTLYNvdJOx7KHShxfmMlhd5Csi8LlsLah8zqDwDSHYXuoB7++u2ikLeRAf3kqLokXU2PXcEE9
5Mz5LtZprW9XKtQ7PPjO+ulp8NyxNkDLzf686VsC4nnoPa4XJMQS5jAdqKIyoFY33ZTe+wBxvAId
BqoobnDcqLdbkQwJsmc2XXQhyAtDy2xfdMy8dfp2a2zY0kVBKgKGStCpBbeSX1J7r+Xl1Nm7jNkn
4k/VJpubasEQgLlAoPc33XxSpvD8bbT3YdiAs2+mcxyBhuRxoCCkjZNVs3lhasZzQcE79n84qaW2
h5qidiGdumGn32xvwXLq+JChFxorfNGYPvRkrjQF/r0cqRisO6e5qBkHyflgdC5HCGhbvbhyB2w4
prk7IV1zWfCOQIuZiCNMPYP+YaChoOJGXzYruR6fxIpSyHl6S4awSMU31SXFmvX5iCRMO/A92UuH
DJaD4Ihccc1e5P7505+VXD4PHurQjV84p+2y5w4hjJYjy2m1jayq0BzZdb7yrc91Bbi61gup2Chl
z6Lvo9qBFYoWMdogJgFq68aK9/j3K2mBGtgvEup7qsYiQF+aCd1/FLc50wsFcqBqnOxsG8G50KaM
16SyEfg+o2PMWi/BcouYGMEqJdU7bm9asBH8NCCs+qoXxPusFNDfEonLV8zZB3bJ8jkp5PdkEYTu
oR82Lu6g3TpxxWsGweoYpZYwJNFmLqrO5+k71hU4865Iq845F9It9a4usEu80HbLNGZ9utYPSERA
kFjUHyJe5+UwMP326R1f2nmP6ou2zWiUX2Ldp1x29TP5gochYj2JIBjqFXXJksoyNuQp6ujAmCrD
rEs6sDafQX1Ve4ZJ6qjiljhRixc0OH5kEAE6YeUgdbItfiv6n8bSshbUW1EpN+GIlrfssgv1ahsx
btDlCspMKcvfabf48MP+pqQe+SRnzaBnCSRrJkH8+Whn8diyqJJH7bmCaBX8PHjICTMmyGn/jBqk
UAB/kEmbJsT0Ml8Nj7mh+waUbt9dtZNIoO2uCYsqh/62acrgWSDpKzxATp10hR5G2Y/cWDjM89NX
smQk9hiCsnwCvGwONnVEKnAx6enDH7v/d/9I3vOWbCostfYC8Ga+sAD+Zf1DfNd91jNgcMg7hDNI
zgIikcwZr51X31LuptECnuVFBgxd9EluLbW7a+T1FAUPXNkR3w0y8OUTORo7kCb8cwu4WDJ9qi4Y
luUHjLkTK/KDwYZ7CH2ZmN8YeBcqmJNRW2IvZOTpHXwT0Wx2tzH99G6otUUYp86j68TJ/Y2Xso23
1ZbJykYedDJW1BGlpHJ0Danb0/LLBDAHfimTjoRHwD6wTX7OH39Cd2Ijbn9M8EaI+LFtQ775hRDd
Dx++5l2vZlptBIX70owF7r14u2854FW/3GDOqLnl+1QBAjxoJWNn8FmqRUhTUtTX7PTkYXsjfXTm
IyZSgN7ayPjG/8NEzdPDZ9H96JPasT1xKenqHfdjRBLs9djUvnT25P04ryLRMWDTFR0vXLL2JkLv
+hACqaZh9P2xDA/3RmPhMkcI8x3HhCvwr0/vfJYfdJFW3vcuI6y+WFeKn647a5V2rWpSQD7gVXVh
rA7OixPkVyJjqdXAN0SMW8xhqIM0ioDp7/UzLTnnGaevS1uvLTbS0VpAUVrLzVc5RFhhEGSSkYOw
kv2jlqbzLpICVWN/LdIdxR5Jry1ZKglx4uibWA+RQkKNbOqynHsCQadIy/Vd0AHpavUDFIyTxIyP
b3+x0D4AEYFMrVMGpIU482yxGQiTXz3HXLFXa83PI3h+slXU3qATyxQcPEI8Bj1ewoz0mn2cHwVW
HAo118ROwHpAsAyfi0J9i7GrzHNBt7RF+Hiaec1HcFEqviMTGpk72SxVopEsSfBbNBIhfLULG7yj
/g9/TyVkqDHmgy2Qdq8mQY1xlq3FJb1OMApJ3qHyn8JU4EzhFR+zkT8Q9Uep2PqLfmlv4qU68OCt
Nnf7y7ZGO9yF+5okYwug9iG0L72kiW6Fe0r4O4DETtarbGSAS5u6poE1x/5EQCMQTzqMlbY7KD+b
BJude4kqihJT81egKwivY1BjlxKpckb3aGK9suAV2C0insEMOGPgGCKpGOubWL07b1PVMT/pGXIU
sHnzTsobGCBjwzPPctQGAOnqG7ReW5ewUkSabPeMOon3whMurt00pTmrcH6Cnpm9VFCJXg2jXpx4
xxBVSWOUM0+xQcJKmi648dN6JhmFaZ3+QERgdDlbmsBd1JiOH3dPheQniWEBbViZv8C7AiNcKAHh
psVSNUhDzUVtp/FVwRH29FO7Xmgtjjpr07P8AQmt0t1d3wuwxVGGa63LLjaL+ko4YOpGiyY+Lszo
T+zAJEFYFMrEgAg5gBKBIfZ/PwpfRke1J5f1zzv4vaJ78VsnT463keEp2qdRzR/GnAY62lgZdOAH
LZHhWHNaHXb+8uM9CUdw2f+j3lZ7POQH3wDKmL1bPCv1m8CThq4lFRicmGN7k2y4UtalIFJZ3P9O
t3ytifwuOEuYtWTWTG+5By9XU/w+/wKwxBsPcFesYbCaANgxrYOIohHSw3KE5h5t1usO5FNlUIgb
9faSB3UOTb2AaA675eL3dyrxCfB6XuzkmF77iiJLOD09/wI6YYHroRbuvE0YJ4CcvBqGWzdcWMvF
BfwDX8GtIfmihRuB2kfPu+RgkxkEkzTXnZNHTUOx5XZq6WMuPjrvng+G7u5t0yhzC+NtXYoU+Dtv
HkG1yqV+n2sCuYb3fKp3lSz5NWrEVfR/iBuI+Sgj2/JpW+GcQ2bFawYHO3bzwmzGSls6pxGHYBxp
qDmaUjzual39jhaEK/SHHIw0pWtlRlwRP345wxmM4SwXfOMt61HTLeuLtEoXc+g1JwYaADVOj9A1
cjsn/MYsbHVp48IKHbuWDweiU9Gk943HhdPiBuYqBrvQF7kZRQAtWZCKQfoSfREULzmcCyOO1Pet
vZnLHGw1mG5xiTIir4ekV61M7LgFcA2JQVj39XwujUBl8UHRiBhwu2+lMDSpzyobC6xlFMCFDyl3
yZZwO6KWUaVG5CS6TgH3Vt7V0Jbev7UbgTZqFgts+UHl8xF+jBzeIjC4UdXUpDgSQoiqhwGggnXD
vwZWop9I6mpIQtB6kZUAnopGdVbyaCJHKMGIAZnh2DW8nH9R4n1HYxQhWheOlp8BT6vlxI0c0fPv
esgXAQnLxgWZT3+2gpNEuPK8YexaJ1L+0xHY7pLRyfVI4GnpqHBrLH7MXAlTuf5OQnbfcO/+xsMH
j5791Wp5rnuefAoujrTRtipTdpzbn+ZmKF38twXnNpRYSuGJHGiK5W2aBCyzY50gY84vNINjAVm6
gvdJJooOntOzzkRopurHR12Ujc42R82dSn14B2dGb3fuzfPqc9pcTZbwlz2JKm1OGLm09DI3LIIl
0fgSponnHhc1ZdA1OvxHLAObHanLjDCHe57TUKPHe5k7oGILwFSpFYQqCFshYJvBZ6NmyMg0XSPN
TTN3MwSOadsfyy4qFYKawhC3N8y9yIztVrxT9P2hGkhO/oXk/+vJ+cIrgTeBF657W9mka/+tK2Nb
WsY6GpXzDeRUjZKfowz5NfEX53YKPFpZwUad4aBJIefBUjxPCV1I1dY1VERmV+vgwCIzL69kfQE2
SQc5FI+hq1wEZsaRBJ99oKnRV7nXFxnSaNTNJoEZGmKtlEe5P6jYQhjHgK1nmmZTcvxytGValH2R
YiTvH9Ik9f8EqkBs08FMQ7uuN7hBhpqFnZlb/QFmY77L71FWcYPlMqwZBs6WDjeJv461UghZMVGg
ZGr57CN2TJgAJ8C9UQoNcP5QFvEJxyajupGmn5ji2Ll2jiHdb2pOy3J01Q9bIehnX+yIlIdypzo6
SZ2Aqo5374JMMDcum2LHjEzqmQbDJd7DXyc1MeeFyyeIl1pV2xG4FbczmseF0eppLIe4gDnQwWNt
zShHtIEAlhmCC+enlyrUNPQo64Sd5f1DtBHicSjsqfNEYactMvr635PAtH3NXzGlcIvOdAJYQ5yE
MzebfSwz28k25qDDfyswYDFYWGCBYOvPeiJy/jhSqvjtcR7oEtcLNBsBbBV3k8mbE/Tl4l0RaYPp
KtqVnLG9VkOO/JXsjgfMpMAsHnTtcBifA+EHVzz5CYtNqhoeWldtx5J6lM1f2n8hPUJaQcwv9U6U
3GM+950ix214IrdO4Y4c07pd6uovms6MxHslVnHAtStUeLeniypSB7lca84VcxJaFF/lG6Iswfcp
msotf36V23engQ1uX9VKAg5w9Bo6ZGtpC7PmTsIztXNyIsyGHXsb7bpK2Z4Ktg9U9hu/IGolVS0G
zGIb2xV66/iZCjOTwn4swPQ+uD+D98uD8PH0otsFrXfxxFtkuDV0z4VjOWn9keZat62EwQ6NJPLo
v8mL6BNV/+ltFcyyQlCWITAzkUPGtsZrv2EfLfxt+0qcdHrqs9KGzggmLKwbPOmmxx2mkjIASloD
L7WS4APaJ10XryFnO0oQMB/V3bcepdEtcsLdgvObmJTSUycyS4hJ7ZQi+sWuiG3pmnhWOYT9tnr/
MosEkd3SG+d1IEORXOxGHNau6dd2zsTLq46d7FCY8eYAESkuBXkKdGqipST4uKdNwe2ETdIuCQmm
HrQqqvrYUf1ck+eZObZH3V6PidKsHfiiVPLogpGikzcSA9BEZ0E6ijZ1/DJOWL5q/Y2ac+Pz6HTs
Om6yVTZp9tCvPz7l2JvTZpT2D7HeeIFDeWSK4aCXpvxWxli2mKNkagyy1OnPWBsHp271TUtJ0JpW
6av5XnKDEZ5ZRpy3BB95p6Ic5bhWSGU8+kMexjcXs4M5mMwjvqJ25/sMabgdBLQtVIpeHCEEFEqN
bu6KHoHSg5u3yQ2u4DUn/3qtJokwdBndbo63H3D/z7piTC5qnvluF35w+shaOlkCfLpMmHxWjzJw
RrxWGISaDeEkwPj/fQP2nC3uiuae9cs6h0my08nCTlk5LoHVunlL5DhlUOs37YPMJ3niB19rKDaV
jl7UGLCxAIKg1p/ANux1ePREamxv+F3SJsszKICJ5/DcLG/bJkB1wGf3sOJ6cslUddGtrOJJPWfn
1+AlaHG66aXYLVsK3Nbk6fJp2n45GHkdLQy0xTrKgHkAZhv3yXwgSGqM4htOFAFTZmxdd1Rx3YmG
lEI/d4x8keNxECvWuMZH5uvEFY0xsr41ZgqYz6A6HNDlejhc2GbiihxdArpMQl5b17bBawhPae4O
CaV3sDmMttoyYyrMXbx+Adh3omoLtzuZKqt+w9hTtwoda6EruYZhA8aI+iWCYAXuehsk1azVh1i7
dU0bC6Sp6JqNhw6BEK8u8kSHyt1SWgIUmMLJ9kvC7h3Odp3dATccRJdyRuY7R7GwEyBwEuHdMTmN
IRjkUkSefwYWP9m/XS+cMeO+jijf2waqstUCh61P7MRhOoQdDqf1Q5R6wdFXwCJT6qgUcZGw6Dx/
TqJFBr5zCntXax8yfu1tggHYHQ5GFI9gkMLVjdSflc84uXTG6Z1oo2e/ZKmszGbwsO+p9fZRoAuF
eGj3j8/FGGshPbiOfwl0PcPmbe0CkLZ9yzsdGrPcIPdXod3cOLgAlp28/UhRPZek/bXcz1BOcTiq
mNdDry0V8b4SIVvFB9XvZ305uaK2F81MsbMKqqQK8BZmMZ8HyLl9pmFG90iUDbba/ojN7JgR8izR
LSmGQqbaKWWeTArbJ+dORsZmUqT5aSRyk9/xTzVYObHIHZBSDoUxVyPI1714Tk7cFfkK03FvtoVj
IwReYif5mSmvQYZJlzVS4F4ujw3gRY3VV+uLlQTGQnUITvPqy+CyiISnXjQ1qD6P3wbSj2dW6d6Z
Tttej6CAH9A5OY3olzU/Ja1zRYEfnXHb8KEUxxipZ72jKVxoBWWFERxcdfIogO6NgdIxECowY7AS
kajzZ453lfjqSzfMJsA9KX/sQ7EjcwdZDxn1xpv+IFXISgu3425QAuYV556CvxLxsRxrUUPNNw9a
BFvZLPVS4Wl2rr/J8680jpPq8cN/q1741/XOgPDJcuTrcWaYM7sAx2e1po3J0V8ybFx/hgsHqSUe
wSKDzTgO/2Gb+oWNvTAL/mrXoU9DMMXYaraDFFyiNvsWLFHOAYf0I0BPTU/st9/xgp7nvIHu/qQg
sDIJQPYqTi9htfwGyWFDxlfOEEIiXCelAdwWGbjcZ+zTWbURqUqTEOVuDW4QZDAb0FGCc3hLpdNs
5eQe58u3EWOBBvkuny8sCjgdzOyya66ID0iBnVC3VL6dp0fYM/diXo/wjca/XZCXmPxVaqXUQzpr
EWoIP8mZ9LeWD7JZm5SzKZkyvQ/7WaewhXmoQFFbomog7zpdnSEPFjuioIrISM/jA2P4hbHQgFul
MeNwzBJPhRXAplJtW+YdBQpjGFN0NiPePq7rzVXnqT/OF67hL+wXzP9jUv+C7Vqxl8qvGJu4nMtH
NztvRUfsWuNccoR1y3hjyi+GlhcrKL6VGdD+J0o4E3IoFetl4nK1DAg7QXmqidDFD/C3YA1+yadv
CWf3jdgSHT4AVzeihCjzkBISSL+KsLZLHOycw6yqJ+51l+scRztUXLgZXUPnTm0hPBTwElEXlaeH
njh349B2Rlsb2Yfulg8I4d95fpSV44itJ9umNnufK53KQaCZc29Iq2BGMlMdjgmfT7ssvLZcGRjr
rlc0E+YGYDMJfSJZb+0oFxL+I6+CK5M2ecCYnH0XkCQDXOWVSV1ABCWMvBojAu8ddlAJ3LhFWzlW
DwKYlmUAgapnC3HgqOOrQ51Fcppj/Q1vXe5jwYcPcosiGEcn6AETf2eGcdGRSsoE+LO/tmYkM8ON
z1yXJ0nVsiCII6zrUiBTH/6t7P9i2Mx7mhCN0C8mqJNWB8MA4brUfcH1JwTDhRGNxPyZYYBJBknc
WypPytC1dqWX0VkKc6Wckb9BKpEzgdfZbi292dC0Wyx7cTdq5JhO6MHmFRk16vsIqkIhQ7mc2ReT
gyziks7RsW1OdAIsZF6LkrXHWMh/uVW9fFu6HRtFIa/YEV8Zo+7EwoQVIN3tFkJa4dVprWXv+6Gt
9WjVqKXMOwWvw+UWfJd1evlqH2176PWB1aBvwxjmldcBqX4pMVujV+t79dQ0AvujZWLTXieuxTU0
s6N1G5sYsZ0V631tDaHt8de64dirAalZvcxdWx7ELIaASTX6BExbvPda1DM/jBEaZqiKbS4YE3an
2I+1mHv8jVeHsts38B4/60e3en0J1VTJiqA4jnidgK7kWdh1U4GAM6vcvohu0lVGIZ3qtEv1/Bst
lIHqe9N8bxVSVpjqUrYmi0UI2h5fBovZp4/cAnFZPcuzsNnyMPxQMCg0IcAOxbwaYXZZQUj+fiM3
yW0hqwJFOHc6DTXnSSK9Sd4BXPtdLoH7U5qTzExNMtPuiMwWuSHTLEsQ9OZOxV2Fk65wRratX8Y5
VetffQFhzq9Y+EGvPxMXd4LNHowpyLGP1YSMCZnlNXwowAhGBhYjvXnsApmGOPuVCmIqFRhADNkY
JsIfPU5ljLjHzeo5ueYiWt9y3RcKg2V6ET6WIMSxsRT7aILNYuuyVbgmh5SVBUEGEwjeBGZ1zpoH
Gih/zs5RN6zTvWzmxMd3XI5c2uCa7Gec0I+LrR8g1ihgvw3kDn8WEfDe+ZKjjpnrru0CqVqGZs8x
fg99MO2tEltX3hb3CC7xJ8SmmcmLWSTS/zxVYeAufJ4Cgi0zpfNpAe+pOStIqQ8FQPrzx9g8axXn
5fB8NGgd3LQ8/s7GBlZgBJ55/SeuQldvMe1qcD3eKrdWLfx2tp8VoJwmUL8nVpV7Zwa4gTucWebE
OgiLbNjIHbBIo9/0h3XlHmrcs2J9cfHqbjT3JJEqCL4DDLBO0oGH3n/tym8OgLSuZYHhC/nJELPN
nKqSAdlR1zYMuFrKBydlfycpCV9rI/0Au6cwxqnxr5Jr/JU+SqILogRskuqN05Dl8sZBxbRN2tvb
7Mv0kZSpCcHsUdX6eEI5KzZmegK8BKol95L84B9vKqOin+doisDgDhTA+uX7jTO5vSl600+y2ceE
CTqWTlDyFl7SMMN2WcRVjuqsWKh3Q8AM8Ib6QvI65ybk/1Beez0mx+1Snv0xs8JZbvkvwzaNDHwb
PnAxpQBNoK3e5Bb06nn82b9njDEQf80amBKU2Sy8j1/62QParDHTnH8N7/9QjaXGwM2aPiLKI3ID
Ra9knPP2fiEyC5LPs1WBOgkSWIXKfgddZO264PivDepB4zem7n/3o6V4UGQTQF0ZdzswpPML6093
0EJm9Ce+fSOwlYPYzTrGeEaY8S0Tmw/81dPZfPk6i5rbbyR+E0+z9Tbl4ePMvoTr79RwsP6w2lIE
8RLyhkhm5/Afu+lLuIDSbrFSBUcySiq/l+n/PFFKCSpO8+iQmD+oXmkfkgfwzdzQrwGH2oLSDekZ
SWnZ+mrHpx+WWkRs7rgNu24zhDypLmLqL2fF+gMHXGvQOY40IHTgjShkUfv/fi6rWtRqt9RZQiV3
FDcfODjjNkSIUxeTPhwiUXxdusi1zK4deb+hu98VxK+NLoUg5QWipBpKc0h2MjNu4O7+3PXqQ4Qi
RvjOf8JYpNSKnQZCMTmViz5J/jGuX2z0g+SpMc+CX/TtMsNM2OghMjoTOx6QH4GpR0Ti67eYnGd2
i0u07+5imOdmNjA0vZ5ah6B30sU8x24nndpi+PJZvPsIMhAaGeeJwePPxdOYxxWG8g903zyvO7g0
qY9aG3vQk+l4gwOSfQ/Yw0STsGjo2vouKOWn5xg09TrZySb/dNKwUe20stSgOQN6m8yVvBC/3dlR
WlDayBcV5qUY2haFDRz4r4MlWH++XQZ86qoQixlxfTNIjfburMuJ2qqRnTM5/mSx4BLib5uD0BSr
DJquTZgtHG4+J+wtDt7Kw/yuhAguSYuCfzRq0aGCHHN8ydtpK6EJndYGNs4Olvetx3ehOZQ1F0oY
5jsWmZqfUZwFnPE7/IpFngFSTRYzsQwTTHv/5zcdP04GenjRHM1n0szwMr7DujtYLHm10uAywpDc
e2LzCDfpqiV4OdjNClLJfiqiRS/rLlcwd5zEnXdtLsz3jS7Hm6hvmV3hm5F/UMpZL0EYMq/TLBag
2zFq8bjqNaAzxuw3QzGnoLW2ukN57DepuIrRT0vnu1OTgUT0Z5sfPHjyqySAwVPCsnXYJw/qRgAU
8CxqMbN29nSzfakVpcyNx9GI3wu/8Ff7wbmnfXfmYFjYEUtoFt/J9NZhUdP7TMukFTrHSd5eYSAS
Bm0XdcVSKCQjxNAz/98n59QWS0ZRjjUWKK7EXlxBnUUx71ZjlVqsenNXSaMBf8Y+Il1M23zVk9uv
VdXFf0Gnoyvf3K8dHhTJpsk/y0WU9mi4ZHnKIopBv8EE9SMsf7X5qSonsyO/+FkC9soRrC3WGmlz
eJAPqN30mLhVrQLOGIhMXayEgx4ZlAr65N84KDgM8yqizf9Bu1ZCGf3Kp9uGXYq+quQgM/nXD52s
uVkrWtJuT/adB0STIg99MjV0biHM9u30jESIiQ3W9zFG8KDDWoipmmXszkaEPXN3hthcvYl6qIzY
tvVHA2A0R/VZVqHg6KyMuugbPsSbVGwCkCVUhMIXg20PnXpnr4LvFsbp77m+1fLIEEhxDyJCiKE8
6FdIiAgx/L/Ro9CqfROarQtT4LRASWKFRy5RaY0KlkqFpHH1AamxS+6sVvfWXjU+9806hKV1nTgb
aSrn33hzgsuj9LGGTorGJ7oFUYWrNt1KlwLindvZsvmp79moCBBXJgFl+Q92YGMeS8S0T/PxYzC/
0p5zpAoj0Hm9lexYV1x3DcCVUbvp3lGYuniwUizJrXYCu/fA3LiqiAQj+ZzS8SazjrQH5tOgmaFN
TjZjVdAW1KQvA1TmdnYYxqbBJbVzUd/w7RqGV0nsTwX+WgwjnYvhP9rUSb5uf8mx4YbdUzujHNsW
iuEy5V+vnmPNqMZTiTUZrbKfioeWKjOG2VxfTrq+drpy+I1dLK410cVY/VTlxM1XQkNDE58HH1JF
ojQtH4lmX0pJLb6n+yovRyLHX3o4xMfRbLexibBZR/prCp6K7ebgdx4ZbiGRSHhl/Es9ecLcmenw
/p1J8ja25j2PS/oWWp6V5vGaePV49EwIS7Xk06M+S/r3h8ftdlb5yCKOm8Vs1eJpZyIU1zN+oQJ7
jQ9Slv+4a1S3MYGuipVeQVrf2EOWsfEeHvpNqzaa1XghTriksWdlilHx9TjGb8aUlF2rWFOY+byp
R1G45qmIi4ZgriaWdHMAYKP5/q+iFlgGVchBAqVqwuxkyiC+csFJ22Gb9Cww23wVtQOtyN9t6nYM
lmxmsdFUbG2+cVLDf+5DYk3wiiUmcmIw2nKU7i4ly43sl1qB/9xjHmMwI/HHDMVol+FdYc+sIYda
w7LVDBTpa9R+1BSjyUUAj5WbSRBknCqPOh5jNcaUx2NHDA/N5qFiQIltaEBfY9a8ayLTLLeHMyT/
KUWKL5oeNpA+YsNs5qgOw9UB/c2JBllopwy/UcxLXBVD+AWgemjd8jmeOcwXb1nH8xzpXYfssrc9
xjkhOxViBu7vJSuYGarH+diwz7G/JXLy5pL3NBssR0KzW9Vd4c4cxpKYvpmunTKzLno6U8EJdaja
KQXG/Z/rn9REk01vWyv8g0O9mA3EgFjfe9W+leQbA34GjF6UCs33GlL7MyA+98M9R8qzMhuwOm1m
14ny1EageQz++OKNs0zXSzGysLhywPbzC6G4EQW1eEztLdHKW/RVe4SiZFPG6qEObYAwYMQ5w1gz
FO3OL5Gvh0M8wRM2IkOvu+Qv6+UQl5lNiAofI4tT1GN+dSLrfaUJzdTzNUsFGgK1LWVRwnmnSHD7
qjTf+TfmigKQ1FUKwEqkbxYZG4DixAuEoYYX8jGcrfiLqM3w/4p4vHV4Jl4FKchlwO3aVBuE8Hrg
SuPseNlV/QNDooCqQrpLhsYr8+a+pTRkO7GDMGF1cgJ3ZtC2PrjOkN81zHbkWuucFbhRKDMoobdY
IQW3kqHJEy9YTa9WxnlpFn++hxbhx+PZodfAdKpDTnuDG2erIbh7CFUKAEZb1CU2BPLNLhBgSUCG
BdlTuFLhQNL1h9zFan+OHSnnprZpFfBdbopssxh4qpjBiSTlclfUC9aQTnbFv/Raxc9NoS7vGmlb
tHEniRdcB6AWleJ/kg1a7tg53QFZVFjn+Dkn5Qd6yxsu1a293XPVwXR97L1uoLlWnoWS/hY18qfT
EaEQGgQbTTW1tSGC1EaZmz2ineFEN4t4DXyWW6/TL5HPS2Ckk+UMvAAi7wwp/7sX/bs1RtWSbyp+
plBNSTbOmM7Tab+D0XGrVLfGwUn1KmYMQsfqVrbshB9cwkcZyIs71c1r4qBUuzNUwdPycvBj0O3B
xzuPtM/98/OsZL/VscoTbiqufBk9UCA3pwLWgnTeihEfVkzDN7WG/2nvJAswVD72yLTqHSz5taU4
K3ORQ2J+4qYLdjSQdzx/l0t5pvOuUL4D9pmYOCkPD8P9hFcVoWV2HKN75jDoDwOvuLznsyWB4O+s
1tp2pbQd6EYagTxUKbxMlteaV3Nj/RSdC5P0SYIeYnZCXv1RnC9s5xlVXns+8WZjgu8n/+wALSmh
zUfTo8toBz4uYfES8rEm8eJQKZ46fystw9SEL6OgoFN05o2LAgJymStUNF/YZSFUoc2yY/NjDRGO
6c8rZTyfl1pfB7aVXSLjZsF/vlGTf2VBvzaPhGbBurui6NcYlns+I5ZnQJwb+eaCvi5Eqad9Jf4a
4gMUz5HXJElCjbAByv1TA4+mQw1Ub7fWXp9ytu/rea1Vr1lUPIgEHWftkwe3mxpICJb2E4i/5ajP
SCCYt22LXC8Yw4ny9oW0FA94dQyzq2AKAYJHYaX2OY/tZf5aMzd+dL+aRwDHKAZreX1jpFqPRxZ3
XQdFibqo1WgcGy6XD1AQHYzO5FwB/djIB45OVVgBfXFS5vN6MeWKImTzxVTKRuE3BycFLbA8DCkB
sdt/iOxuhN+Bcya1BHMDOM4up+bNizo+ntXiIJ0RVo1KxcQNyXDdrMFTc3E46+gOV1rM69hHk25D
/0+RIhCl0J3QvaNNJbwHuIs49I52lyRWnmBJZg6yG58R7nylgQioNtQsacSqg532fTjQDFtbQTI6
djNbVPIo4DTvp3O89PONF3/5qLbZqfAEgSV3jeugttdklcZs6LqaeBJfskft9pxWtEozcyFlEhjE
D6iHnpn15cMPtLBUwCbLuIfnSe5xbZ/95kb6bdLmTrAbm5vW42fgPD6Dr3J6615/4IZD4aaObLNW
NrPuk9FuUiSo2dS7vl4ZjnsukXQ9eoRW6b0F3xsfdaB8n8ikzzJL+iJ0Q04wJ9/NY8UCmAv6zA+T
ls7UUxbdOsUPkTtMW4DrPRpvQYCuHgfClgm1SEc9DLPWRGDSJsHWHmAmkwpJnwM3BDcyvilOMNgd
KixTJOX6z8d5RO6YiFVWK/Dh+fjzi/At5I2nWrwP5XBKwHk0eBzETuIXjNtAalNvlMhHObzvTNoK
p9XjUye8pDAwm3B+ckMZ/NhIq1rIMBgEvsIIx9lmplznoq2VgcCQ5IIBk22iUCmT6tbTe40oJN10
bt20FFXuPFTM1olNudGinSpwcMK4jM6ICH6a2YRsgEfxOeFsfTeI2bMzLwkc18ABl+LUVdorovRI
CqYYQLp/EWH60ukjg/F0BJ9+T8ImJWf794CmXoDvCd/vhfRwRdTkmLoi7pRrSr4q3HyvOVADA6vj
Iy/PbTX1Pt4DxyfhKOXgMzrdmJ1PZcvr9vp/6qw+yq3GvuWxZNg5JBF+eecbshJDUy4SlT5Y8sRr
3BDmhyihzW6yXg6dxOPUNsERkxS/IMUpe8txliXFoPeg+jO1zvhuDb1uYQz+Ya0oq7A6RMXFAq49
+YOPNcmRuQR7x1yTcPDL8abM0p5CZqWBz5UOwn7vj0OHohef3Hgb3am/7Np3z8pzL1WHrUBMsulQ
90VGZZVC62x8rmnqnolmyZ5cWgQUySlnVCYhLBwItMnBltKvG/kSZ3jiZwkP4RcptAZUjPF3IbaP
2AKGi/Y4/9mZuTqulbpibzBZQO3V52r9E03R71or2T7CahcCg99bpa30ouc2CmKtIPSJTwPgTRPq
BY23CAJ7jaTRWi+a/rMZQB6EaIhK8BPNxPNRVpthwZDZ/IeHuwYVbsKX/6u1P6oHl7pBfUxo6fzP
ou6PjYMb42aYEB1YIEh2ZvBPZ7vfiw8FrOTB3VSIPilFiRWT6jvqex907GQVE4lStSoY9yzjl0MF
9RMo7PhkO+ewpmmazeENYOWPZ4vesoQOKTWD+bFtN2MRy3nZt91wpBHMpn3D5WhJtIRclGmeP2pU
0H/8OXNI6k/3bSXO2nDyLzG0NTV/nJRfMkk30kPBNUkVGhqxvN9vLihrEoZX5eB7vLYE3wdRceEn
qb+5F9TjgzktiPxcqH/Fp3+qTgqWLArR7uq9eI9dX1E0Yl0/s723ArhpR6dALjfUxHRfINhRVR5t
Yi94QP6zjxZb7F5h5T/9tzKNKKOrkTyAu4YiQ1UNOtAiklgkKGBeRGEEgVAIdc2UdVscnEczWIn8
TosuaPPopPWfJL8hwrf19SGtZuJ8bai6QT5fXXj4wRxRI0OMSiRsZFqhzKm26zQttT4k9GXr9uWf
5e3oyP83HGIQ07fZ/IR/I98nVnW/f5zNRhK1U1tRUW99c1iQ32tRX0G5ypt1eucI/7AVlJ22hsF7
AqNgH8y/HPC7hdYPiz9pU8jUrdhdT+4fQzwkBXX9FHU3w9CaIjokNJe0iwEMSMOy8ndK+6JM8iPW
SosfzNIj0b3yPz0RP1spaCIEnRHgYiIAGlkZUFd/tBYGhSEcsNE0qRjIywQBLCgVW+mESRpyDWGS
kKxnm/Ybp8RItdwNMKYAsStFR5ouSQ2s4rpGeNArrqQsny2UzY6PyIh96mmkOuGSaQkMNyPhseLz
fPrXTyRyZYB0Lri48RJ8VF/bonwXaQBlmOeSn7g2c5SRZ8k6FB79/RR9aWrigE9grxzQXOKzqlve
bemO0EnXgxkqExac/65jBjx81Iixmp4R4i9Lb75Ed52Ykdjp/Pu1+NOiMHUiivEm+rTUbqgqdWrY
VZagLU/Nl3R+XGIeYJS5riKI/xeyyag1SG4D/MeGMjFjZ7iz2n+2TZlVa29pZKcco/u81o/MckZc
a/v6GCk6ZDaMK4z2HP++S2rrOUNFkJbohD4QwJH2K6HM0ols1VD0cDPiLn4iVlpJfZaVkLIuXmK+
9DkT0G0QYIAz8fU4+xkewKtoi7MH0tpmATwkCWIRt9YEMldfUMFDqPjTiFbPqoFmjDab+T6eXDd1
2tQn1uRg3wctNg+mIRNO0DxUncxOprn5z8FTOqWZJcaeEuP6JPPCQ+tgH0J03gZzt0Y2RyuTGk/D
AWu6NtHRUz2uppKiB19rZ10dlRUvN+mRQFyNSjkXJs9wG4M0/psXq/RHUSY7ihcUiP6e789fqCdC
CLlH3zD2hL1KpvsKl2GWLPoIaB0CyjPkPjhuSjTVvVvMGD/jlqN6ROgY9TOn7DhU0wpOiX68N79J
qgy9ZGTzcLFnBOu9Ti1pAHq4tf7kjLtwDfh38OGVluwbPNjZWyxeg3gK51TyHHpZbV7RRfVECmCp
46ItikmjPz2FqZDX3XjczoDwIXLcjyLYxM19hEhPK/EvY3CI8VEAHzo2DitFaA03IHtCLKWYfXOh
QYEezzmEIOQwW5lckdrMg0htqxsXDVZ33+a+kWB1BYFDHBGt+c6uPGFae4PYk4OnaKmibWjZxo7I
YaeXOhBeNgBjRjFOmweq3L3ynfxbb3ZofMCQJnZi+mR0dUbbmxD5+qHlveFAifUqQ030/w7loxhN
JprJKhMpQ2YiAEZGgJtA+vjaCqofneMA/VEQrUKLp0ulxYP/mvIUbEGF7R1IT2s0IBlogefOZEOo
gbwcdgk47Q6dqSe9lJCVxMvsxMAVHdAr2YVyiP6SeGS4EEMMCQwg+kkGHHIi+MSTZ8cQA6P9e7e1
WDL/KU1tPiHmPfbdtHOF95v6FeqMBuWk51fH7EQ0GbUrQdtrTv+digOle/JTipRcMsuN4RLwYVHJ
4ytLp8ogKa0XgMKkZTdoRYJD7r0h3ylWZxpg+1a2HCW/kefWtPAE5ytaiHt7TJ8xSWAkxdVWK+5y
VYn/bmT8m6MgGE49/MVuiUmSR2p42YuCaK4OGrEgQYLsE7cc6hmkqQXrYaqCD/eSrzFj9CvC0WtB
ZXtJ4JpCX8/oNHh5a6nqj/Nfz3AO40U+iONikN2iglQtp9oDE+fxlpaeNKo6hQiuX6NzHlCOlNkV
lPOIX8MdKEAFU/rZ7A5YMQcKtx2Y1iN3zF5BWlJn95HafVTrRKCEebeekVj6rzROFl0ZDNB9DvAe
158bQrbMWjhLv9LD4TQ4c8ORW8Ek/KgHE3o24vnDWodWRRMSLC+gRa9NY+ngym9YVU/YVnVDWk7q
rjJ3BwVyDgeVaazEItNkobbg5DapPY1Nf3oeZ4L917m3F3LzaFYsZNozZQaC6C7yxnG2Vxm7wk7+
ZYDN2Ftwn/hZDNXWF4oeu3TvJQNwzpM5xtFgubLx7B332nluQRQ7CNM0EjmD8msgHIABGpLqTqPf
8mV6I9fQ+NkteATJnPO7hyALubNEFm+/Yz5zpkGigmg2BjLU5l+2J6oHXlO2jdh4BndfN+Z4Jhqp
/6L/Ev2yeQ07biWuwsqit+O2903FiQ67cgnAZfUq8ir1kTvEhv6EX7XcJUA/92eL9bY8VXNpgLl4
tYxij9PZqUkDTbpXmL7xgUBvTOPNihIlmRxTl/VGd/6P2QiHE8qoWp4ReIZcWopDqCw8zhaRqRnB
uPAITvG/w45ktb1l+ML6gk9gnBIe1PEOwJkGTVFCVNYnbWd8gzHoJQkt5WkdN2uvX0J2FHILm6tt
tlibXQwWN2AAdEyvkPsHCUxFPwvA2+xCP+C7MtWuIg7rlR6GPSPOKhNBkLKO1IywnM/ZCfX/JyCc
SVWvIKNR+/eF7OlZ4cOwEXbKImXPEACSZ+lU7IV/fLMWOq9rFFaLm7jsT5vAylNTrLiVghTXZtgJ
IYFyl7H85ZRd2SyOlQdtgvCTnTBclnLhIkdLTKBYQyjfr0vLI/2w66JapIb/y2AQ0vlEZLmNAzn3
tZ5Uu+Yt5qJWdbgKOEjBTLrjLrTyKbXX8r/1VTn0pyl0TfbNPkaTf1sYxaDlrNp2VcnUkdUhkoPk
iyi73nZdeJdSRbvE6dXSazLFRsarderDvA/uVuSe+VhyyHwyl/n2JU7Y9MH6dqqquycNyCsN+R9t
FG5Bm6ZrQN5oaiPNfGEVR4S2GKyXO7dPiTuEidg4I4QqHQw7EBWoJYX8pyFLZTiQ+udWrjzry4uh
GNf2tVNNIkHbcM6y0dEtsfftTMvIKl0gkzdTCfhtr4cO38Nb2b+Kdp3GBM+u2HOTc9ebBjwQ7ec8
g2xYqyFGnRlKzZAVXmjB3mEGPbj1yAPBy3v/rUv874V4eOGwhQpCHJhFIhMzGq+qyMKokmwUCga4
uCTXpH8rADQCbvtiX78clX6gP0dyS5Sd1snDn0xvVCkESI8gFzO2kGsyUO4nQmuSg+otmk0sK/xM
WgJfTEMm5V6YTeXJxCWbRVoAt/+2zRMN6Dj/vPaFtIGKlVBB+qpZhJgWoaEHLShO4sz1yRFfdbAn
gNTgpAvldbE5puZQ/QZrkAepBriJlpvDjS41s+jYKA5Ze0Hk/EnYpdSI48eh8uyDlJT3j5pNsJWl
fHzcXXYL3Hzz8x+buODttcDmN76Nxtn/QHPVSOCSi4L7TVQphHnbSV/gmZvFYvVhtuN8AN/DNUBu
IBgsj/oCrL9LPjGatq/Z0R/kue6GfEHIUE74Us6czc8HD+UH/8lFIsKW9i6cnEbwNpvej4Z6JZxy
DCaXaaSq5gdg3FoYUp4uFTK5r+YBGT0tZhk4NEqfecja9CMbFTBvlxZHejv0u/QXNiUWOVWKND32
hOsJHxKBtCJ7Wv1ml+nmv+kTWXHMBdGtr8NHwfcFBDU9PRkwK8sCsUPSrPpHxtPRzcHOZdM+pf/w
lhRr0eaJ0U8/33Ogkec1bvXZjuiFzCjA2AzRDijrA6HEkO4leyJrPYRk1W0icyKshWUaPp2UJy4G
lTvw9Zoydh0Rf1anMlcwokJmLZZlrUvaw7GXUn0Vjij4+M2OiqJ5OLrlY3JuyEvhnaR8pGqkMi80
4wpWiBUTXAGfwTYDnk/fcH2x9j7muo/AIHWxOCIXBwshZWGNZBNw+MKQYki78sSPwyXAN26mVpCB
9oJtkZ7TttuAP9MEMTjEobAntAY/CgLQo3YxNVVDuQoRCXTe2oWU3C9/Tf8xEFBexDZUT0zLhNCi
TdpAG8Pz3BgLh2Ans5AzwYXAZ0WxvGWXqhsk41KvmZyMrPy47Yn1JxVYflaIqaEqxioucjzObQd+
qQDA95yA3PvY5LMuetnNSlTlfGYKgjLJj8D7gayz8rQhTPvrdJEC3jvOjMlEfVzDCmqWK4BbIoRZ
WDZ4xnLS1eMv68z/s/FPTMSSGEGXvtsIv91+KWnwJ5do+nS33vj8VxI9WLeRtOnSCE41bY/3EB5v
FOQTsRaHzStIMXdUoZJgVcX7WlBXWbEBJOpeKGS+1Dq5f+/SIrtkQO/kunyTJjfbAil0/1n7JeRF
qkWEf4uJpk5WdXxAzAun99cCO6UMkqGU4INw1RklSpIpVHzMV1j2y2oDCUzMQ0of6mwBcmoKTRHo
kPaLwJxTpFFDsYpw8gUVyl650iiQyWOEZtcQTExYURxsqiVpuQkw4brTtYpZEjao8RET6c2C8tBk
/s7xcY4ZQVghDl9g5FHxplKl+jJXyny7YXSJi8434ss0nXseY6Ki6weo0JkLombpuVuGYc8P+GEu
9mNGQAHDhhF9qiQzvCeC0dDMUHZ3lv3I+CAyJ4mo4pWXS52rY6hrWKNHmCdZR5UayNirbOQdpQO9
tWMyVH8U2cgp8VA+yZvwI5efhaQ74PxWumoSber0OrMyK36i3zKqqmjjPlOsg+SRX5WjbwkgiSBF
rZrRUmGRdKRCJ1hHISUZnBUwOl+ngzU8iCjBZkpTWwnR+q5XB/AttVe0/XcSM79trzbH+8QDSIRi
MsR2oh3od9hyMxAmE2noCksI+pOLYuj8XhWnL+PbMyMd2J+AwL1XL86uJAVd+F7e4I4Ft1CuNCJ9
mKyVHQirOy1rqvMXkS05JC3JCT4fMFyICIkc2+qUXlnLRUtqIA0U6VSi7d5vnsT6HAytljBz4UW1
nZKhRHw6L4OtQvJrzkeYb5VK1l/OxS0ta5oqshmUHuskbbq1zFH9RFYjXLRKia+JkcaLK3a7pY3Q
xa92jlptdw/cizuzFRDcaLpWY/gH7X/Vxg0GZtIbN7RwvMCOtSHsH5FppZlEA3OTYAHi0clVe4Pg
3Nskh6U4UsM1PVFzUbnkuLeMWmPQhCcefr/SfdRfzkScioD/W/vGVrsb2P+eV8Sqo3f2tPI6JO/3
kYces1QqdMwygR0rjxokAFO5SjvkDgJYkKH7rue+CL+s2ZXjLl4Vk6Q3CkdiRzCIU8oWH3MsWOEd
oqQRxhszk/GLIBRRfzAwAN48Vkdhj3b4nTJcBwl+KTDSHiFtNfAITosYgoZhzbvZnWXsB3Z1eiox
DsGw750E9OlvNKD92yZejuAlJbPbaXfeJusV8pQb5u0Y/qZcUorzjdVIZLTU4OwRHZt0LScUmNc9
DAyq4tfefMvJJbPYNP5dyqpOd9UlF/ZNxTyC5u6VIHceI6vYf6d6AGSogxp8VTiGbAbn+2F6ToH9
tvDkdRsGv4CLOqCFufuRPl8Q4bmAnOLt/phoyLkET3nBB8TDted1Ihz6MFPWhId62rSSVsMVPKYP
suVN0okEvZY3Kt8LU9pTYQ1RhZGH8efumyH01gH8x/0j5IdmlaryLO997SCNrplP9X3KQV9EGJQ2
oWaYyZVj7PqBFgLltJa3uxYoRqtjPtuSX50w94mJaIfx+XWGdGdHlV/opXxa4ID0f6IUBM3ieTjE
r7Q5lrUgX33Kv+vPPY5Smm4yofd5+yt1JNR6WD+OPI5Gb7Ir092zTxAXkzM9YLAeKzElEinXaEmW
SpciJUly797eCOhwXb4GWobUPYB68vs8XQhBVhZNVvNyCsLmyjPdot/B0rsqDhxCJ2HY7IKuO89I
KnNoL+l8SSa66vBvw5pVyj1XJznJrTwhPnPkz4j8gmahxIVN/oEMMVvaKiODRJ502ndBEgi4WAeK
osQKLeV989X5VpqrYkElWYeLUZrg4xZbR92mZeuLnGMjKSe1wg74X81kxvquXm8Px42gtr3YVhH8
mxTXP7U7+8F/cOsF6g5Vnl6DKqJnUakVaCpAZzZZ/ImqlcyB1EeoAD3w8Ac40+jxYE9Qk2gdHvLd
thBQViPuiOWYSHjAvfQWLdZkWE5Q0OGU9CArFlQX3gnVxM4JnDUbi86dcD1M/W1ytBd7LtKWMMxU
S3/uIXYmsUrrvyVidV0nwC2OvNAfyJFODBg/mjXbs4oAyb6y4PBJ+RtxYG+7D27AgOOO0QQInpo5
4+zoklftK56QtnEK650Q29TkSRTpAbk5TIzAKGbtjjUNXsqXws+LedB6OPQlhkwTrO69gyAC2y95
Q8cTqVajaLv2AWz+GM5QM5c2/msnK2Z2eE+h2my/jnxAjp491CpeRSba69imgLYDSlSznOuFXZQu
x5HCPXg/fHb3TgSi1IjMDbX8ZEChSjfxoRIxj2VsJp5uTzWa7GYgH/um7AFi0ggBes+7zeEwD4nF
XKj/8WDY1QnrNEGBJHhi362kHOdgQQHP/pMavEZsUP1KP5tGpbWsSyCAPgb9ySj9jcV1pg+UUPW3
k4iWyvYHHLZhKp1/dwM1UNycj6nju468hynzuRr+W4EnJH4iOC8sMWbPslRk6NorxdrNlmGJG0G/
aEESKLsGa0l6Uq1Xgkj8uVzqTJN/+hd+AVZVJ/w00qMIQ+eB1jhO3Ru/j6lG3Bnc65hjuk9JQRsq
bESfUV81r8y1Zp6rzbdNeh6wg9yGmmtpy6+K822AbeK9BFKrh/LdFXMZgw8rku1VC22mZyI647Fn
FrYCUxqVDRbA33DbZQPUFg1YjvUZo+TFYrStA4uXs8vE1CmiuQ4u3AAmCFXrneg1efGq3eP+PdRp
tvm62vm5FaNIbEDOCvZlXvkria4nDjbOPaaF9IW+T8ObunHQDg7yhD9CNxTcOLQ12m0yTfKw42Ew
OuxPQ7ZSmwTCJ1X2kz29wC3eydAG0SeQTzxiDlLl8+zECxnhtWUt9boZDUXZWja5fy+2BQ7EMhrg
SAPShYiAqRuqvqjSL1ZoebQE3I8zANYiP5fmuEqKqEPMzjI0fFD7N5N7CJx5X3ocjs14oMh54rl5
hxjB7rQZwrd/Gb1zYU4AVTusbo3UDk4mWo90/8FF9W1cgAjHhdjAsw8S3yujwfCAfadxfDIALsam
HjazT52g6oUO+7QXGxCHIUPyNALrmm8QlFpOUOxfQfL/OTOTLTRJO3pU/x8yt1mlCwG9QfD+173+
0Hian/obqJZSbGX8m836ZUpurKizTNXljx2EXehHe1P4m6FR0L81el7/fcHXCXPEZn29P+nTnnFj
nvzjFcy9eYlmpE34p4mg709trm0lztt1lRgw/Dy/vQ05ifZA3lpX6aoonjX66yQiXpgXAzzO/HsD
hIq+8Q1c1m/86r1xFp1A5TrR1I62hjMuzQropGCsCyxeO4sz1Rsp41+UcEm/t9S3Eb/spwTH2aLv
/BMR2WBF7TsCKzWFGz4Flthv+udsONK2EfFI9PcwHVkkKPhnGtT7uLURvjRKieZv8CuF6X5QYvKw
NiOfxuaf6xDZGOcifBbSVBvZ7i7xoOxOKgah5w/X+ZmEBPKrdM/nXJ0jYwmmDX8cyojDNYs53ALI
jPsI4dqWvnYinTuVV7jQ/9MrKEbrKy3VXBzXtb51LN12E7u23Z/B4nfNYHWDkOSCU7YaIE0EhytY
emTgXF4GOkBrnHJ8ZBqlT0TMlPd09DgkFsoKvhXpBngf2R63pcSFSwV91bPrUyecy3Qk/ZiQP8fx
/C7PydEK2aquVViMnrKaYUkxbp3ldeq2y6v1zuqZgF04/h+6bojcrRrp4F6rNZlJdOBBmAE6eTd5
nMd+7plk1jNkkLn5QUzPSL5BFuVawiFWIq3qtsYiOZfu12g1xRUy51YX0pERFzQThQ8WfgirqvZs
GlTq5kVpicnwU38YiC1ny7bRmOvxN32wFl/Ek+iRlLgDYIvbStFLdNqQqt+wB5AAszvUTvSyl40v
vcQCNJfLKAKpKq1tn2r+ck6bNHY4/HCfTfpJZBlH57ImWumjP9E11Fu6cuCWIqccyaodhWusLM20
fansRLtMTZ2wicBv0vYpPYsRau4gJHmAk0aS28QP3JM9yff1aTUvECck27m3Y6PyjcEnFJhWFUn3
TjDBcnfZD4s5KFDJpmVBd9jE2u/7KgqTw0PG28qSnynmT4VEdzii1pcucd/Eq0qJN1eQktYiabTM
H9eeFalOG5s7Tftu1DRA+edN8REYtjALw615ATcwCSP6yOKqmTeZ9JG0qyDm/EV1js/hp7dCYsCn
2SySpxhq9cifWIECIHz+vG5SGeVfK0PLnQVKPHU0P/0gMoQ84BvBZub15AxqZwL55lSHHB6Rl4kL
2YRRE/+SwC7+zVpUWkEDBQpsm1EMBDtx3IJlfd3T/K1dWsHLb4V1UP+0YXKgsbf35SEEQi6JNUkl
CKwUj/yg2l4MV7KwI79JJNqGnWMguPm55S5t2XZd9ZOhkWH4MwPXibl/4CnI6oFuO382lTZU71yP
vxe7l2TSzLoIJ5lARml6DDYiuCqnAi7DYWOwyVbo08ZDI7vS3WKcugtyv/84Bt0YDPL1WSkMWY3F
JMYMW+WqiSUUDDSR3F0bz1rvyvuDX0EqcxTUlNh4DeWqR8f0/J4NWtP3opOo/7ibVU35PUM9E8/T
IuelFbbQFiD41pSHOQ8Ru9srccuoGW8ih9zUeM/Vvos1562LlQZT2EYd4tXyAskbRIpD++zBj/JP
Qz81v2oXNRlN0qA+9OQLqjbtj0HV7Vxe0q79DQuKi6JfXCtnz1WZ8qfDSmFwRZBSgbPPPAF8VZ4U
xj7UgbUJDR7nobovEjFaArBWLrmxINV8Nk/cZRT3JDRc1dpkx2WfT64J3wGxgwC0Aa/CB7eeQOu9
P5DWjh75Be+3oeyRnPli56Ao6PAPmvkRf2WD6Hty2F2px2r0k075FO9F6MRWyb9ziEHY327WDMwO
dJrE/+17NHW3G1MG0SzItkm0xaMyx2wWuJlbYapzf69O+J8JdtcoTv6LF9DYF51LEuZTch3agVWa
3tjUMFttFM+jbSwgv6XYdcW2M9wwyPc7HmTZ/A9SfzFL9OXxvmC2TqVrKTSadBn/rWCeMf908dpP
Z/wLIqLDvqtn/mw7E4cSBwLH0+qNTUgJONpjoKeAnJGIWUT96ZyhGLAk+zEAHi2nnjHZQBucs8gR
E2DfEz0zqGXLRlqTtLFSZBf9FFaAyUw1Rvkp51ADsy3nP5oaT3e0SKEZVk+0cROHoaXXwzWNi4AE
Wuzyd9x1ZN7hkpOYZLc8+b4bBO7T+LUDAwfOvKW9Z58+XykHPZfnMF4JYGUPUmlOUsTktDfl7oyI
HNMo844q2NF04Cvm/oqLhysjpqVRgs2eTj8b9tzhFEsQlnhsJ8thbNdb732t8MzMlyGGucm7oLU3
UXFHSBI7BfYXEXfChtKk3ZHqMlThd+O3aVR6v9jpWamA4bfDdIUtJw0cgGLmyo3LYIw4eULSToxn
iL2N+kcl34ofHaoeugfzMACLckwSOVbH3jvptvLGWlQtxMBtM9Enkht9i/dGKyEWLbsNacSD5C1N
3QX89gZyv/uZidKPPaGxqYvuMQp+AtIX8Gq00J+3I3kcQL1iYQyopmeYc7nzBy1IMX2YEd7NCMtE
rVPws8yzEJX5o5ENJSxGmkg6vbYGH787XqMpZop7rogiRXGPCBVgbevHANbUM6PXqbeZBtoO+1Hb
hApxVtfoaSPO1JbkT29f3ttRnwV2GflWysPVW9bH7fhTvPKrmjyjeOCgYsCHI8IYXOdNKrQBLP4y
MsKrJN2CV2ZGrciatHinlGwoANDXunBnp24sh/16Hhrk5axEnWO/jeX0oy80i5YzLA1yKNj9Bg9i
1FqXwOM8qNTufS23Y3dpsVdYpYUY2oqfv5wA9MV5NoxWrjNW1wBnn0kFyOyye7W5q0MtBeCNn1z+
nhj/WM7qRyeDKHFEieCFXCo0J88cgxpR+XG582WHP7eWVAxDROXNbnBxTZMI6GM68j98tUWl3ZGO
WnVn53SkX/WUryryPmz0AeH13Ar4Rvx5JGWW0T0mlwBb94R1TBF+sp5g4TfpyXnfsP9loIrnIRSh
HFdhHMum/gB3t5Th2f0CkAWAi0oMaH8QZObXr5S6RFeNVEorjhjAy7cDQq51sIL4Fqm3uIlqmD/Y
TqYsHyNNUm9QhN7S9dfjQL+w2b12L/LSStMiizKlRBKGu5bS+rFbUajRG5l0RVNlmz9nzQWHbYXv
g55dOyUwwQeUIN8sLKmJ8GnrFlpu1q+bS3mcbdgJxczNBzxZMCoci1FOuIye9XbTqnfds9HKBzEU
HFehiQKaRvEOR79TxJxudQ+5ST/CZC6562+3chsJ4Y9oV/lxywBbyYdG4XUKdwId3cdcC2L7+2Ag
5Jh7NY9epCWOF+Fg5AkAKB9kbttUYXe3a1o1duDhgmk3JunHbc4SJAPdBNrfMGjC9jeRqW0k5r/A
4P1ewO0N8ws0RULkYfDd5+JsRhbhcGXJqnNLNP05ca9Tx7JKc8UvY4KFYb6JR1ITkPVXg8Pitosh
1BcoG8U9xMRVve0ZLkDZUdrjxeQxO3UvzsSXxThM88OmFGUAipsA3yloQ8V/9pUYmPHRUEJrpOZj
JUseHv1rbQG/6YQiElTslwYn/Ne82bnO3yKnz7OspEOZ+wt2/9x9H7oTYC/BqmOrZvLJ1pdLgkT7
g5F2lqxvZZpT7CRDLjGJ++94dTKAmnk8ENf91EaSWDqb5aTZZ6QXs8EFQHUbbHn34/FDSN24/eVf
WJjgPyUaGxBcr0iMyGA5i8suyGpXVZvrMHUPUwkIohm88y++0m7jeug+LsyQKzrNpzjtwWExWT+1
2yU2mxqBdYsQjY9GpfKNRmdaYAgE+zbtAM8eWeOYFFhIuLJDoQd1GJHzOGh5CTIsJqcunDSm8p2q
y1wcgN5MauY4HoE7O/bJouzXKjR7zilj4TCh1Z/ZSgSiD7MjgjppMNqXwjyA4PvjgnfWgabR2QG6
fLv/5Ott6AF2GTGxjpKiN+Xe+Ytkw5y+xDtH1+WR7mmWLccLUKhBnEqHIvYIrylTmhSgAlHKq7zk
HKWjI/gC551d/xbLDNXc6y0oIA9hE6IP1BBBmg79DnyjWg1Z0EyCv3CctpgBteMf24NHFVgdhGRs
ZYSNeZ1lTBazz0xvAJndsbsJDBOU4EaYoyGxv4iLrUvoR7FcUJ0py1P2OsthGvPDIxjMp/h89jul
Q5TwMUUD+ReICKHrYeL9vhP7o7kuewi3Mi9znyNLbvpIDC4kjOGjGJBIQwPMAe+PF8A7LbTI+Tsh
gFd7dLNoTH2eHw1PofK/b/DQeTAhh0LpQfxfKKMEhU30R6OVDAeoviDrfitAdAw9wM7YJQqAgPb0
28IVHmUL/Cbp5zhNJGm8jEIrztw+7OWyU/v73QUIePDyJJ/UrBGDsiw/JLyo4HiS+kPodGOJYf3B
NkDlCrKgUNhptZ9TKSGjgn1iu/HR8iGRwpcBbTM9udUwLCNIoI2HD69gxQMBkJ+dmcrK1gETfsiG
r/Scs2wUkOooSwHyXFeMh6O2FUlu45/wilpsm4sRi3WqM6836sEdkZ+Mrkxca0JHE0Cd8451BUvd
Yu3okvLM2np1VUNyiNwZA17oKgj3WLavALStnbBM8PN0B7Q+cRZZSkl2KcDv6NQXc64DdtjRqpBN
PlJkMuP5ZppOrcTo66010fFfGCKt4NP5c905/GJmjNKZ/5IPijVmGVNYa3Fx7lHTGO6XoKwxFmd5
CKzwXuwjW/hGgI2uTzDzMHLHnWdwxLB8G53Xz7dzBg98P8ehTcnxHeFWdEWMuJwpKf2g0YrubRcZ
hHP8Slo3RXVDUXXjCoCPGcY48J9QQlUgR1qc9AZvElE6PyFcNAx/1Q8VH0uAPI9URuWu0qDcifbx
9H9jlUHHbKJX2X76hJ/1Ayb4X617hrcJVI6qNVGDyMK8eNs8WvWJFEkYdevWk49TBCopaG/9S/yA
Id7TWRK0u8u5TMpDA7y5D1DN/xe+OG80Ld2LvgzAoko6K0bTNMasosyVWoYh1jJzoCCLk6lGfdE3
8jtMIQjehpdXpwnIF86Z1HETvhHrIKJQtumnFTpRdxYiV7yk7byoyKFCd8+w85/i23t1Q9pZtnFn
ekntDQ4TmsG4eqpPLDcLiEM9lbHKgxSkeswcpbkiuAqL5Atc1qLU0LcLBg41vSZHBDzHfmVE0hZ3
FUnq82YHSf/FlatnA7d+wjnSbW13vy5H56mV0TKqzxo2CLev0KHeEZG4zKjPJKQisdD9RDoEgvMg
3s+gfHSrRVMfy+zcwejg3rJkn1iVZBnwaoUTaoNYs9z8Ifw4G0CB+BTabuOnQk8PqQF4NJUhNB1C
fg5q/VTf493yPtQM+TZTl8SMvLo7IEQmLQL9s3jaenGPQWYL9LUd5vm2B4o3O/JBbkbYsEW6HMQ6
MryWOT4YAOetegV2/9sfkpWxa0Zc9wO3OA/b3GBK3EesjOu3XNhBqakN0i7msu8wVN+OVdGrPMiO
y0xSVE/IGmxBfbN8zxrX8VTV1t/khTZfx2bpS6QCLfBJOMlYMOmdHYUgT6r/bbBo2qSaL73MBo+H
yRcbZtp6o0qnfWk/rEYwJp+RgwaDfTk7Fh8aLehEYL03cKltHY1SrYvB4SCcnDiCovoLotqQKhqh
jpEvEkszBQeJdHRIuT4YvI9X7gPtAtuJUj6mXrKPc6x+TlOCzNBJmnr6pbeB7BgtE1vFi3zefGqs
2oLaY247xrLSQvuajQoqJVpwNRnIfLfF46lM/mLlQZO3fMCIPP29hVZRVv+K+y+e0kGICJehjARe
r0aJkSXCScsOhWtkd5BK38Hw3s80MhvViKltfGZyEcUwqrH077GpErCbB5K+DczR7NT/fDcMnrh8
4PrK2heCZLdMf+CVQ5cqZICYoQ5jUNbnHRX889dC9ktKxwdelLWZQASoD+HXl5Xi6iBDmXS8m64j
Dr6i+ukd35StyxIo29rDvBHdftojy54TFj+j/2qxQv2s/24cYLBvXmppH+aG5g7+Az7mR8CzMvv1
OqIIQc3/yyRMJJnYSKDWcZ4IsMG01KOttv5cwFvC8bXw7mTqbI/Nx3VQqlPFvNcWln/76LBQvguD
uQewHR5GWsuILph56Y0J4s+KJmUq/gk9jHkaeZghm1dwG918omqi97UWgmqUBd5JSjKh7K8HWFIu
pC5TKrhcSpe2sR6+pf1XyrTw5+4521sp0d1D0JKN1Om7/nplA/zLYYxbnaakaT9pT+sd53MzOfJY
gnW7myJNzcQPh1JRM2EZ61SbXjVUdWTqFz5CfsmC7TTipxDlWeQG4BZZzKGLXpno3/pGhLxhm5ja
7a/qXSmGz4acSQX+7aw9mwBDiqFBVHm6sF3r2mGDivD75GVHs9BaD9f/qELwKZ+SWIEgI87h0gCC
onX5WYby5WYxtck1Tph/Lqcmm0clJjQy5DVyQGQhQskGk6JilHctzJNhITpjhAMr4YLha2VrWr10
pXmUw6QbwicYR8Z3mdWL5EDtrqYLY3SKnq9u5Wk+H7j2gFACX73V6kc13Nhcjacstj4g61Z2Mlcx
e7BmC0qZ2Je/CLv9jn87ETt0+RkKMNSd4AGZxv7GNv1hNQGAvbZucjjZV3WZDHOrMTQEXpTgxPuK
//KmxObmDfrbP0vF0IwbpCV1zNkfj1vD1okINnW/0zEKJ3T4/fRpUW4gPWeDCWfd2HuJcNMdOMaX
8JihyHEaPy8MTDsnO9xaLZq+SlgeAlc9/6/CFZmewiKmDZCCb4MuFtN97/2ozzc7pN68xVzk9ghC
+gyJc3F35n6hX+WsWGa4QG6sEu3KsCGs/18X14QJrDuP2UgZJuXApKLWPyYpA6taIrnDuAqJ69Gx
3WexC5CTBhmDzyuI1jgwF6OLTrXpRDO9EOQ0nyQWCyuSQEwLVJ4HLwIxXGViQyOvjc4nk5xtkLji
IHPrH4OQt6pNXKxuCP/hbIT831lpYX0Vwbv1lutnX/yJ5dHUNTVgCq387clG6v4N54IINNuVOIOm
VLQ6ZwXFX99D1j1cPBEtqTI7ASOSU/xx8+b4rfBkAEYn3LIKJSY0Y1vIwg0U3N9+Tw4mH3x8K/jO
A7IZr02SXtyN8dXSHKHouYojqb5nREOEnoeFmebTJfMbXR1CFW86FI/hGS6eyUEvCn5pA5+KXER/
PwJ2YtjlvrL78v51zfTg/RVgz3JVkaCz60DQmpfHO1W7ITqNXLMnGiUNaihHCNrbf2TkxEs8XBB8
mC3BHjmxeva+rCZBEMsAL9bfJ8y36ckuKfhXVC8SnnYxUEb1dtYYBGL6z7lIXlGcVa90FY3VgVM+
jA4LVh31avXP3l7lX3INq5O8nKBKdJ3kyZKbLTLcgMrL6b0Xvkc3SGQX6i5bMVSV2qvcGjeneKgi
9XqkNfwPaG6DDXrq0cdSL7+4OCX0D31mmUqZrcvR0D9uRHhzJzHKjumV6NvEv0FFAWZt7QA/hI6d
iMHFiQnGJgFYMwHu89F7GlgZ/T9C1+4FzGfVl3cS7yl79oVy75EgV3vN9foIOktsVCNhpGXRF8fx
sOfLG7qVvENwIILZEp0vDERhe7PgbnRsGUXili2BAKtI6i5ooXl3+c812DSgtPNRufjiqbL1FGMi
Xu+aPQN8YVmUF0K9YB48ukNMXEsxTk56ifH+dK7coaDcFzUcDkqka0QcnlwLZ/GUObTLLHjZ0xns
lmSmgHKWSs2D/Y0oFVZmWx26VDQFaRYjUjQHMwIm3+o7mCk5QFzBhlAGRIlWKgzx0q2xzpBPH2IT
ExSH4uFkbc7WjgW4mD6zWnyk+hxZF5KoP6XpgOJCpstJ1Jn1qB7iIHheDEThPRfxWEx8k6nUlcWV
RFPyPjDS7DK5z6OV3cZgYkXxuETcqdkiKO0v0j0CG/DOwq0ztWJsSbZiJbJ3mD87FQKgVKjngkSN
H9jdJTDRwAGXDzzDXaQD+rB7yluHPNSBBg6kjcq4N+zbzIfzAWz0hTFgnitG31ApX67QmeK8h3dV
3NdG8wW/cfhD6R6FNRYfiJSe82n97LnuEvqUwB8anINcdTIuSIpZeC1HZi1YvyRm6v3kbJgemSPT
Bwv0XEayPRUBH/Y+IMPQHir4mqGpiBwDqyGkfYTfyKKV4QpiID2nvZXmyLzeefqHHsuBI4bCWTah
ui6T2eoeCHgkxS1FlMJToETgkt5Ny23/NrDoK1cAPfuck7exsYhhh72dH+eFloUGJ2OTz7NWWcqZ
Sl4pcNm3Z2JoNLt2p0R9i/6DlstCOwNo7mBaUvIow19R3d7fEkv20JYFJPYPTco1ALV4IeHDvcvY
4GObkAkbXYPFf7o4l7uPSSa3vkFMPN6CoxetvRPA/ByXPhH1Wa8H+ZyRfzI8S4WswxLBU5MCAwkQ
9BLqmqMAr620HYfMphX1YCs7HE8ST1PilVT6BBXnuLlMIA2twEAnSWFwEo/R1KqM4XItg1Nzy7UL
Ea5YXxOauB7nUiv9QKmAGNCbrwiOo7QhAXapJRg4Cr1gvPJ/0B96RrxIuEDJV6fL4qVL1X4OMUaG
55lkg2jxIcVARneOW76Ft1y3lEKfCPaWeV42x6VcYcYIXQ3009mLISr+gY63NMZwLY4Yy4EaFx68
BM/KzrHM5xRRDizKBb4xViS5uBILmeNv5ln+fjKRu0obeaaAj4uVXgUAa8N96Wmsim4bY6fCP/XB
TQgQ4OUM5C0VtHtzmlpCBmn65A3efgEZ8ICq1cz8Iz8o6linH93DVO+Lo8svCUoWICrXnSzqfXB0
j/1RMHd6yjaZpKWNEzlf1LlRKGJC5udFU69yQZKTMoh06fN4Q4rL2mmXK6gQpkMOvdAfsnY59fD0
5PLLqqLbCLp0jQUCThJ2mxN342kRE1u86Ld377ZirmoVL7mEthM3J2mPwJmtILg/ypF5udP+axmo
fIQy70eiCPx5CSZsHqteiph00ESgA4rWH96c1owSIBLLWuOEq+TVzEYe1IXhRQi4eO+iwjgJjqNt
vSrGwLxOVkPq7ISjOwyaBfuYvGyKpoBPo5j+Z0PZvZ7d4IZx7jDXepO74ppYpkEcMobm0mPOXNNF
44q4P3Q3I/7bsmN+2W/2/MZXwK6VSvW5bIxhTgVHZyYDcVMxMyexUtzB4CkRsOFoC88XnDOTUNLa
Zd4exEU8oFhaKmkFGkVwgi6J32Iah1mTIa9yA1SNbx/7RVJ02UfQynHzC8arRuh0/jBNUFeTaaYl
oJGzdOZQWyUpwkn2VKWdAJRAee2kCcECf/j19rVp/UbCDf/OqUiVcIpVsODhJlFxrXfQH5S2+EeJ
m4FfCHi1ZQWZoFbA9Q0yrja6TODzrbWbpL5dWRzA93ipmQe33s3UfcZ04ycBPFkdgFAJt8rvo87U
YzC7130xKpkG6YLTBYAtaeWiiIZhnVmcrxu20VFQi77VQWpDmstCUUZyMqjchYUOC3SBxwZ3yeAS
TlIXMY+fq4KjdaIJp7OY4dYf5/f3ioTmqmsqCi7hboUwCPiQFTJ05749I1PfXZe1eTO/3CtEpHJP
GjitFMyyz2XwAgepX0xd7gem8M/9AHqiWNA7145nzZsLXywfuInDURAxXCqOgv+UaF/VWVlVT0Wg
a8vxiSYEleW1PTCYC1vYsJwSn5rtaeFEqAv3bU4D+iF3CC68teBNh6jlRXJyT+xstjgcXi5sbVZ/
IPekeTKBe14eQ6r1Bifs+tRyC4GYh2NgBryFtFLJgJZUSagpx6UkNd3q8iXwbOpok3/2VTQlP8Q6
QP+yzX4lQcFpDaskK7Bfkp6iQLBPs81dl3MzS2DvjjYhyw8RbvTIO9e2aiglHdGuVrJjyLkTuxsT
h79Co2lNjq8JXSQ4QKbwxcAjc2ZCrJOcd0Oc2JeGEWeUFjeNpo4ib8A3/L8GP4rHOZGAtlL6Y4yg
M9VlN92YlAgzqco2vf/89eTboF9bx2qesJelAPbSmeqaaNpX/UWvHcLGqw1wjsD1EhUB6aVEDecT
D1iAScMyEyzmkbh07n59NtPCyDh7thzVZsLBVEiGcdT6rZxUGpGbGLINzZ4xl9tC6/fXHNSkZtnC
qp80GcCQTYD/Sp8bQzZwXcpW2bK5DjrJeA9RkUgKCH8kp1U4sZIMoJ102ArxlPvgIkIu5D7VWbM2
kJ5/d/PKvE3rzdiGAS+GmkNrfmxbWJs5PU08iDr4voMZ9GgYp86lmmBL2y2bBObVYjCh7HOp0xzi
F3gdYpjX/+Hbww9BwxqbCIfD8oObnWdafZFY1wSIoTXOO/qpEEXCv+wQzmUB4Rl9E+0OrdajsiXQ
t4m0xQqDcWHqbqxt9ZHOQ/gtX1i7t4EN5OOvu/DHeYLEsz/2VF0WbASRipQVTjuak4AFhguXAc/B
HgnqjsKob+SP8rl1Lvj0nADQdHk8zZ7xYU5RZfU/V/KcUFXtgkx39K5ReMAuGRnZa293DCgXhlXF
tfje4tpqBkPHVVLei0ZX0uXbH5R8KzQWS604CB+CCHGcyMIhR3xOnfkS6KtcN+bmmV7ODIfK6Yu6
pTDzlxJmop9POjdkn2b1KwTc+R5vQAKhyKJNuIRDs6qgzko9QQ9bGOgrh+jL02I0MLwC86KWLzT2
gxZbR3JxFLK5gTjPmyRUz8o4b7YdOwkd4LS6hDEWEAv0hvkMwtqyUMDA/kUOZNKWjqFIQSErGXT5
DhBY+vuM4r4l8DxTk9Ht/hOy9cdh6ZMMBVSKlndAXLkDhJW1BWvFoQf9f31O/TmfhwaWVs/aQgoE
Wa/BLAp2bdX6es3KqkxZeLZW2O77mTxEXxuVgs8MfTimGa2hsc8nLCDyQtk50Ic2TJhuxaIvpyg7
z/jv0jKqcCmhulv1hVfL688GthjHs2YDsb0ONsRYveADFODSB2WeiPK+0qtOG45CBVTYcg1mOkfv
ejm1DRUmAFQNiG0YAUT8hg4nHrF+cxHO12NxRYx6cwJ6h5PZ1/3q61GxgAwvXNMYJQkQ/bUtZYPs
APfbS81eMsrN5dHbc+ydVboB7RBBcxdrjnkn1BR3c4m5e7yW/Yh5ViiD3FRXA+lZ0rVGmy+vl6r+
UWgf++U82lsWr2cgsMipUCyT38IYvtdFd2QOgeh0JX/a/INePDwRAG6cOh423AVeL9SjH9TgIrew
f702qVM7sRuWbjmICtaLjIGzdLToLE7BaAi+yzisG5OeeWeVk+fKZm+JEJiVbN5pcjW1/BIrih/Q
hGlZY8GXvWFDzZWNzoPUjorZZ1dAJfHlBWXJL64sEHk9LE9T5KWQKiKSp11B8rJ+rrWq/yQgmcOm
dc8rwEQTmfP3X10j2Ms0HD5wQzmxA/XMSWLUyXK6q/XIMVcEWdZHiQ7qKWu+2JJgqu0IXg15fzDQ
Op+uI1pmNMT28uxHjR7Ldqx2pjp8TxF8qeQLwMrrp0y7xCGNiMYprvfVPR64bYxhkI0jxC5YmqfF
+zOKU2TB3497culxJXK5CFW+lUrbMDWcY+bYQMwSnBdCnUnHr2mQvEsUqngatWGuigZyUkUW4bXz
ZU4szxHs8FVmKJhA2ViHR2hrDTEnX42S7zuDqLOazbmT6E0Qr/2BLMmMK8fSCJraDNrQ/r6fKjnm
H60D0UOqkBd/qnxEnmLc6l2lboAkcOpu0JHmxATZCX8eQFhQLKy/f7dwJWPb42T43b9IMAUN/zS1
zIS0DbxGhFbH1XWLKx8MP09SKRZ4Z6dHnADzeH8JIocmiEiOlupK63KSxsuVuJnhHi/qXJdilzq8
gisnEQt3sKr1GdYp1Mt9tNq5/SedNdnChALyrzNXkvqFKNGq0hEp2jduyy+lvfZsV7Iv3IWKigcx
3DnS0p7xXRHhbZjr2KPFgNaHts+IxqYEecn/6EZQfzB4qzc4am8i94mPIzvZmvcTeOdZxMhWJQsU
b/fyskZSgMCWFflHbb4u1vTT91xs+2tv0o6lsX0wwDnBIPRg/uCFq/ptD26sS88stl31rkzvuWyi
zZiTOYlkd8cswH2/eYPJtYm9qk5SU18QZ1PYvN4w6PDGN1/r13uUl6X+Mh7QbRTQ+6rg4lnYA0BT
HJui8lHVXX5nB2pDQp645wAKh5XJox13Uf1PJAcd6+hdjfMg4f55mgmwkiqd3DSFStrR7lAPKZim
gvFZAvpUTPdfgb5tc9/ukkZ4gvZHnnmqAnI9ryZoZir/u4ouQ28WE5g/OP+/Ug1SQ9bSXLeMnLDJ
I9EOcwrfx5pE76/P8jUhHBFzvX2TooI+cTwXPbWEopMhMoPjOzyCTtIpi6e0LxY6fw1yUfMtfECk
7XF1SfD8Up3rNGXQ9010x/PsLmQW1gcrDyV3KpzeIssL8mUWhqdBGB6fCVO0lFSg47gBcOwOnkrt
waGyC6xM0XmxmNrksqlyuubVv4fpnSsCK2ddjLnVncJtq59ljEEHvaDn2TM/01fWPUqIfwg6/D2T
LPwQ/9aVRe45iftbQAtu+iKDXmy3HYFuwXCbh5uiAFu3rXnexB/1mjMn/4GuQiCNYX92LAYcCWBo
76ky1WePjdAyXeAfbpdLAgLKx9ejjdKHP0DZ+T9gKNqE4+8fAKalL5xnGXrjcRMpuhGhg2cNhUT0
MtG9FTe7+x8oGqaplFwMBMnG+ms5cb6vc8FLK1PtUtSYiJT5hreXNnCmf9r9x7eSHX0Jy6KdlUFV
oX/ZtJqhJMxfXcao+uUX0PGWsrx7xzXHKFHLXKuxQ7Of5EHW+JN9K26M9qx3Q4zfZbP07UcG4GkC
A76AWh7xE0uMImoa72VANUlZ5HBCX+5IHJeMw1yzzgePqoIbK5qIfOFUl5dY+xSLRjeTxmsvOzMq
D2IVGSxwWWorsPafLMN52WxhKOWDVv2vFfIy0hOOV4T6L38nUSS49jY8gjofa+MuSmEbGnhS4Hlr
vx97ShA/17RXeZE0ZvfO3UOwjFJ9REAFJKUqZHJYnhaWWNP6ehBK0z/VxiTFpzpiFsdOKJbcgi/R
BUPO/6Ml+I6hJY+T1RE95V7P42WpQdtL4JcOQvXS7KUwnGGWLoAfjxG0WLCy83R46raKnGaFf5ED
rBgfAQe9MbENvbv+kgBJx+WR0G0W+VopX/t0Bps7IgGCA9qjCAKCfeTALY8+1uPjxtqiJSonOI9J
XJnYKYZSyUVOcWvc2rHHOy1UE8+YEEHUvyRD6BNEaHPjO8PRbt/yk6NYiEExKMfoJ7etnnU0k81H
SBOlPvpsF8EnIaNnCOCklsTgVvQiGX9hIFn/kieiwmfOc70v2U1kTXTneuhoWtcu3FcMkRFzT0W6
NHj2WSW0XHwsyQvoXMfVasm3eX3Ct6CslFw7g/qpaD8EBpZpNej/FQVTWjXepJsD9rz5QIjY9Ftt
PZQHB9TGVOBRX8naLIRDsQ5cmEoQUCrTfuYwNdHFVZigVaqw/jUZntwiFFRoslUTDXBTtUkLTctM
e0A9yxV5FHG34ZlI5ABojz3xbY1Q6yDBexig+K6/KIJfk2Y0RX2+EYUEHyYKQ2/3p2WzzMDs7Pr1
XwDbWyYuZT8rIqv3St3D8hutYpeFd+y0S5IeTrKSDR+/52Ja1JetBEO6QLNx4HW1mATNALPLKqkS
HD5sr8AKtQUaYxHvgPWcH/vUkNuEJafIMQDskBhpiP67dbrObQprv2NN4G2phHEizz7GO1DCPUNO
mXkFqERrfZNRU4iJbqjLjMyxh3EHfU3YXOv6YdA2yqA0bmFzdb+xBs/DSKnPR3aPSNW1qjQjjWGg
WwrUEu3X2h6/ohFoG+gjX0l6rvMYRJPlTfktLH2d+k87kOE4Afvv7gVqRmvabqGmkeigAeHwYWXc
5tecYN4kbmv/2FMk3k8Y+IxfkFF9wsud/f882sEm9Mm5Udb6/Ys/8PhWII+4o+jokZ6w8AWDfHNA
0YZ8+7SOXt9V2/OJPuTQbU3Oo9THbpVFi3HLlDcTBwhbrK+IW/il7kG0hG5SJK3JfBbLwhshIir0
JNUZEYOSkGSE7/IC6y/Qqwn3i0c/0DLDUIEimnjPv7JS1F7lm3Z9HYWoAdud9Q4F4SZMw482xLuz
tcbSu+G5FDlll1iWjMMRLRh/otivbrfKs0XpmizVFqqCH5BXKaNwGHYmDuwii4L3xnbHxtALya1R
rm0lrYIOZIsdSCnUz6rf7HzZtoxVbJ066ZGXk6JrhNV9AtvhyU3IyBra2soAKRLlMYYVgzSGeHzh
wUL8th+iLNYuXJd6qGA/uj5XuNZJ/sW6vgs5yB97aAonU6ocgjbJhfaUh5fa2DUx5lGnb+Thrsew
8q3I9/y0B2xhewMpVNv6dIyJJyi7hNu+AJTam9SX+f7RiA7NHEDcHf3cc5URKUmw4M9Bq6IAekjE
eK9f0dLEiyzkkMPxnehp88cD0V7MHjcAw0tQqbTA4I1F8DxOncIJHBwGtCKesV3kN6DPZLLuq5dr
g89baXu+8R+Aj17Rgat+FH5M1q7YpNZQZsVZtZaeucfeMoSZ6iqHHdduXhSWmYG+k+let53oVF6a
qlorQm1HJ8ycVYQ0xB1JH75dEbRKORoj37DtveCYo+Ro9TbeuSi11kv0MRulUGeqTwyGHJIVJ7+/
UqD9Lpu4WnQ0me9n3GMpgohuBs9Pp7ds6s+K16IOUYrRNZFnX1d8/OYWJhiVPiR6FtFDMRwXcUjI
q7afl+7O0E01bem0pTq55dz14JNX/uhLx4IJjAXgXB2L6RpCtgP5WlIvbYNjSb8SKqS+LYR+jpEb
NuIC25l16gOnFz2aMOKFj2D5DM0LOEKfli0WU52OC0j1vDBMRHBS/tmda9tQy5BUVIn2BJqXHyoc
obEfyreVH6IQIQKO/Pq/sRUjsVMTepa3KEWUdFDsunBCEPwXH2/KqqGrKD+n/UUamizCQla9mlpX
PG7brmp2EEVt8Z1G/16Wqb+ZRIo/6EKNh/LOswgwdI7JZa5NutxKO2HtciTmhlQV6DdXS6hDff0F
O/DlOAdKru21JRQ1KtuuzZL0+IveDjgBXcKi9xAo6QCb1cMMry1wY0KOcZKBf4wJzAekuwgXwRPI
3pXrYteAccCVBk/yXn2ebPssTgNUNZ2WWKqiJFPdgtdmJPsSWfyB4uHrmCqiZEkZPHW0eq1a+PMl
vOkBBOXMB/QN2XDHEKNm4u/fwZY22It7SAZ4IZ4DLcgAj6PLDzx70ugaJhj0zix2g18sF+IJd4p/
vUuUACyXnSlOczLtAXMrU98hAkLai9lnDNr2ovFOEbfzyxku5jL7dqn3281G+aFL4yg4kJG9yumE
Q+E6CzmSxW7YgTySebvW8Pld11r4zg9pvbL1UritMdbaABTA5R6xtGaX4/CBBPRxAd6ZGx8EjFMp
VwGF5XTW3qvCTEqkH5RjQZHw030azK7eqAJk+MNF0DU7Uye9tf8GERpHCPa9SzFZEqAeaiHqG8LV
HUg3DD8Oq6KoSnXEw/BqxKVb/0odDJZflfCnS1Zvw8TFymB+bUqKA61mfc+4cF6zD2ByxsQKYov4
IwLxIxgXooEJkabkUVkOBeXWt2Z/SNoj9tDkjpGwLqVgJUSmGfTK0UolrA9iF4IDY6QBTKVpzuGH
w8vQer1lvIPCp5U6UZlYGPo+M/ixRn30pg3UHRJvEeZBW/8DmF4QwEmslGUpbT0GYj4LqSxdYZYI
b1sO4b1dpNejDD+JhvmtBfYd2GDX+qKAjza9NXgOfAF99iUmIAfPgAMJx845pA7SfIuxFgDYMphI
4BSTZnT/5kLkIoBaiyZc+hZGp9LtMiSmD0c5w7Xfw7Y/cT2Aq4LGq2vAMOBnISNaQ2NyhX+5nkIQ
zl4gKM8v4+cIRpUddnuNIhsbAjHKH4j8s0Yg2j3UX3AteQ8xk84ktKBm9TOl/w9FbxXegEhjz0B8
DuaX9hiuW1NtmbBUjegUZnwEx45uTdIgtHs/hZPufF++ek9dRTayNM4+22SyqPEBZ3HNLf6426Zg
wr/KL3Khp1N3Mg7Dr6aS2YZt7Q+Wt3uCarVlEO5w6KRrex8eRyK4QdlOGgboCl25y0qSzGquLuPv
oXmsh+WomRmAc9kKOCNacJ3Js7rcQw0HxQIVOkSi7ZiEaCz4P0MRWRu3jZ3zcAuUFo4k3K//5giW
mBVA87TKv5cUDhXhZ2ejjNu3GYFPGn2WWeQW7O5JbTn3ImEHFYLPNl6aCut3XXombpNJpvaEmsWA
cu2HQ6O0icaZtB6gW0CGauRworjbqODWghXW2Tg/2Q/M+kELG7hVfxxr/DwNDA4LAXzjq6YXOiqg
VkVTF0H2oI/qFDtHWBoAjURGAK4BLORxV9d7v7D7CVkgxBR1bviMvqC549rkDKn2V1jxdbhtyw1w
cpN8cgYRMXys8WaYK91GJvu2k4DcUG+y3wGeZCiFKYINcse4Wu705bXoLo8mq51IictXAD/EI0l5
Q9InvBcqeU4EGTIQsGcofejnv9fV37oTMRsh2RuHNVckM38xsD7h8bRP9Tq7wx/B9BLGrw3T5/bW
pd+Y/amS+SIvN5spr//nBLNnADDVgnbnTVLAxNJJheDPZpvtAHNzcSif3foY71yHItz058TNO95d
viSD7gI07/nwc/D8sWHrsKqFmrRbsocgp/DgKmsH8leCgVvdeHWjxY9LSNBQdQyyIwUU+nyTlnGH
bptKh/AZiejdJRhYxkBR9CF4PohI/WF/yBkAQWUoFdaFJXq65X4I/CcRSLLyQFtXEwXgQYwCWIk6
wtlLSmkCX5z8gGlZcHTdaxT23FIKhpwrj2bv+VvF2QPr4UkLHx5YaDJJdsR+8e5bl00t923mdkYA
dsqn5+CuyHIsqm4NUJ1fBKg3ImGXh/lloSW0290OYcKtrCaD+5vue+mzXwghyWBkZvTy6dRT0UP/
fVss2yxUFiR+tzsROi61b78jQFcgjv+P/Vl3Brw1r5v8PvYORdof9v/dNBfRhlebkfRkFITtlMGO
VrxVbVYf7+KHJGrZ0FAQTdMRhvf61wOfpK/BioDhZnzO+fPu9qIx17Fm5f9knxsDkEthJgUzRog7
Awsh9guHDX9C7bsvk9+DCEevH6J8hCLAY5XHjBjyq0MdPIEuiY3ofiEyLbt8VwuZJ4uiUvgEjYYj
3TLPhxgyDDUbVEgQqBHKVRxqsSn4ham6ALMJ+s07InE360EXKq+YJKq4X7GPAa5xJpn5uVQv2B2C
ADtkWyAm/dD21Jgitdsb/nOW0i2o25v31p+DEwpqmVr1XtYMjr0r7U8z1xBYtam6AdLFiBoKfidh
xboq6XE1ED1GQCvnUW3+b/kmsgsprnJ6qNwgdclkrWNyZ+BiZDKHt0Ga3dlXTzpHvRKCZs3OVva6
cJeHi56pAqj1bpFzojTNmFiV0aP8pw3YrCPGQzjh7qf49A7nLirReQsCmrEN8lbX/7FTm4iJFzYD
iY2XRADbLpmXgMNSfCGRHuKngv3voEd99X1kCAr0ddY6zDAmyariFXB9VYBNY3SlgCJBTFKZghjj
fVMXL833+9V5BU6wtBVTeVtveAaqhp5/M6JIWu1IH2uqfQ6ORvRST46UP9KS/cVF6UJ/zXr8gUdt
6CaxH46/plclo8Pt+S4GFQPdxsxo5kmxbWpWDw4ZnRYfElI3kpjzZ8MipotI8FaBKVK6mgoRGMKG
BWvmN/M8zfDDMW600xtsceX1dIur7IoNHB8SeO0KLyBhXpzlrjDzRjTQLoL5I2zoFy8IFETrV1mv
B+caMJxYH6I7t1/x/EIclY8CMN6g+0qNFYxOBeqHAgs8OwNIIRm8gnEo4yHfZyHxC5rt4qUDrBM3
MPNwiA0/VlKjW1YlosrXTEeZO5ae6QRz30ylIZdZMLp2ozUayHg0/I3mu1EylchvRW4QhWjo/4Gl
PO9BIV9s76D+18RiRPTPWoi6VBUVdGzYHqz5qFYA5zcz3vszMBLI7h0bjlMGY4DwjfkuW/6mQyqI
+pTfAe0Rf7tga//lV0biqDRBM4Sn1q8yi9z3xGpA1c7s3lanxUDCfTpwOE2c+SlJjZLGwosvZ/Cm
nxxwrxmX4UtALxrZVyv783JzBcWbIJOPyoWkU2PnzY3Yzn1csIJ23QwJfcbd5gA8Tt0+URiUk5Jk
YNuTU6WMGxtZ3WYR6JWQY3S1A1IXa/7e1f2URPQwzxoX9gC7Y7UMhwWJ5KTE1Mx+zlge/fndtClX
yheGw/gYFq/ildCGzN82IdXVTH9isSThUEUJihncHqNRdExZkOPLPiha+vsgfG8hPTzj8WUNgYKD
XCiQnrU6+cyr6o92xE74J28MdrlP9jkyt2a9FZRGjcvUOc79oU1FokDxiaK+wANkdSngAMOMFC81
3ukpe8sLC9KZO5LXZ59DlJRCoPEG1KM2YcgCJlpj8hBCWI23w2Oq/4mM0ZL1qhLx0OIU6zQfSavi
hxI8h0ZRYJdXHoGwKAJ5/KtmNsxVYtgbx/rsal6J45kvAgQ4aNBUCJ3kLZAjnK3b2zUhBQwC+Xrp
FzaTTUr4AheFzvKBfWEa8jX0Fel0ywWJq8QsekobQmlY2YVhIiewllAxqe7SuRKOT1IWvunIp4wb
hnKJb4EIhG+Yj9c8l2HBFL9inZOVxP7048lXHtNWpmScuh56YnLCCFu2IPXT8fD6maVH6LbDgetI
HEteHjr/d8e3pcuDcU06k1mi1IDoGCMeKoVjkBxFCIbn1LGpMATEXSxQ75G0JEeMjPyvuQao4F4q
IOAcY2TTWnHYy96AaJP+v2mkq3/AxmSV1vp0nM2EJ1rIBh6mdfeNb48BO1xkcnomlV2f+69G/gDr
Gmbtxpl8ET/Fql9ZLrXoIHKQbLd6wRHUrxUeErcS9mk17EoC23HtEXHOTzxkPTaf4hj2a7netEQt
Ghh5D9i6x1q+iF7RBTsOVnONbopSNx+Qd6dBGVVjPgPDvkup2tIYgXS8v4vGOrcq524poPQOJTWo
tqJ48eqhk7pbJOteI+0yoQ/oUNzYIhDjci8gkk4pzEkDinJepbB2T0tlaOz0uCqQw1YqYOJrLEpZ
k9jPmbs1GsHZrG6v1QNBE5egWbFfDqHOi9s5mfE1l2GffkTz90oYwfRfTrLcVL8mSgIpm7ORxIlc
gmbhJ6cg23n5rdMNColNQFqVsG/iikHA/JXQf1g+XPBqePF26cjty+eCJWFCcvXOe4KaOdVBenf7
8NdUydFp/PuhNQDrRSBn70aoaOrM2FqrarJ6Nnwej5DcBgFQP0zZSNUa2NwFxjbAipgU+VNOVVaT
abQpqFTCOQhJutCmMjArmDGV0WcQQWi0ZPcd9HWdazkdJMxaVn3Kjg9cnpwhwrx83Rv/OLuY1Qws
5x1gB0vTT1XcUkHGMlHPaArDstJmAQZeipbf6IU0C6Qsuhyz31HLfwdHZt1V6jJ6wgHEUJyCJqnY
FYm9aYzzHMAgwbnw6FiffZ4IPIXQznU3aAgTKVWZjGwHa1H27xLPY//23ES514ztxFyOeKW2J62H
b/vdW80IyjuXnsLcStrnmgfrURQ15bmDnMPWLVvQSUQWe1sg9bLJIs7tjJk5jZNf0j8P5Imq7Y5A
hCwbbe3wM7LwqQsNJUQLyg3PuLWPWuN3+14cNAFhK2fqziroX6i0hnu/k4zvwH5eXsYPd+smW99+
SQwEyakbl7FdIiMUB5V82mXN0AqvjJ+bdRNoUqFEmSmy8KPuLqaLEnxS5R1kg6Bf3PQXl/vXQMLX
IVJHmM5yAVmD1ZSXi5AiK5yqLCCKxmHCGPTSwA3nMpxzLQsCbOl9a3SSNEeURM4/QwprxDg97KNO
wjCow6wOiuJqK/oYJxYr1lWMMY/t9O88lrzw9do8ue39bgVZoFg2km/EtLPy1/w8xE9CylLO4eAs
ajItMpOXsfpbH7DCTUXJu8nW4jO8JEO9FrJqn4dyO7QVb29gCt5uPHr5sOeYxq4KVuei3X1BmrXW
8s+FYq5pjQXXIRkWo/t6bPdQo7FDggkqocaXR9IoDAFycZ9ATbeWITOq4kQuvbk4utqCO5hEuu9r
3iPcU3ujU2GhhEdnGeVrJfZHeDS/b5QrsNY1MCLDMOlf+fnOwVzxFky65nr/LzvJQ7ug6LzCzzJ5
/qVF3tCBL8IQc4uGK95KoWZ1T8G3Sz4qQFIKf4fof/IfT12RPq2IPiCMHUxP11iwc/AqXPSwJ78F
8N9Z/EiLrruKrXhP2AFrYzqT4YOCjT7Sg73Q1mnhzpBsNVQ8pB8qR7/p3RmWeTONKOACjnQvfIIR
e5Aj+7s70vpxYBkmpsEE4nl3BBEwWqIAZ7cB0L2miNZNJGgeWT81/LFG4vC2mkHRJ9/VtE65MjGG
iJwra8yqcD7vFS+ASu6oUaZGmskXrBmzXl5OrKMIX7sCeU75oWCuVP2FBxekAm9T770awiwwIfje
UXJ5qEHND5NE0TJw+/PKPwvjrUhfskrRNg8mbRo33/Beh6gFzHcCu/6+3meu4WCIjlQn4EqDIQvj
8gRlNICP9VZTRDxxOe4IIyDf8vFUHfdnGmwtD9XzkPqTjZEnW+WCs8b6heFtO5AZG6OJk0Ko90it
5GZWH3w8s1xTTBVRiVX5zNsThdvO/c9w2LdLXT1snGlSlTkdEfmmVGvyEVdNxBylUqG95WzVenMF
DQFQJzJjgDQ70P8PQRkIr4J4nNiC2JfVytvC/tei2AGizP+c00a1y4dj9cF52OgKBS7oTBlWhGE4
NCl0h70m8qZF58s46P+9kNtfXqODP9MBYo+gawmtdW+z3aC/vUSJD/dTwuTYPdtbsp6l3Jqdc/R6
Yydrz0bDGdCdlhvyuwvgBWJRm3iqOnqUA3q2j877dGQ7VBik+qAb65SsLIFnW51ouqLRAwKklSJn
GHz5I7bXcNfbLwzgPgZpjtibdATNOvOw/b9zGVHUN8Vz/LhCdMnQHCeEYVzNYPMafce3YGrV55p/
nStIu2Jrbtd0jxhsAnkKuuJpFbuXFgcG4E1TQqcpu//pwATqJHXqyzrBzxJt5IwXJx6UngFB+V56
WFJIpsgbP2jrUAkcX9QoRPoLFnS1IFzsQ4Jn86170mOrQX+nSmmp1s9dHwkPRZpQqch+nwc7udBg
VU6VjNzyOzrVKTg87Gi7vKGnN8zsOFgwkPMbTx1MGbe5TD+FetFjaCbbcfdxhgUEtCdxO2tQMPxq
3lRDNKtCUE6S8uBMfggeSBUxkPu4OaZdObKt4uMVNBC+5nAMFWC7Pd2EzwcEbatOVXpfViaLkuBe
RLQKdTFyGR0y/rho9sarCdhlcYKNnd6Phi28I03j2cGNdvKyUI8zLtJNHFxn/XmswvFq1qenCcKx
LEdypUZ73p0JYc+elRaRbijYBvHuQvjOtX25Ejz7GdgHD0ZZUjw3GDAno1O7QUOneLAA4CpfrU+L
E/xfVLyR00yMEE9vulrOW//oeemltpJaORYq/c2k7BjY1dNqSIhyqE6R4zvTr1TU597EJ0BBP1oc
B0wgy4N73EKUgt0aocwpER9kuSBYtqSuvSDtN/hhtsxNozbqxH4QSdTgzYpIRG2UVQHGnuQXtTmk
NF+yBrinq7RMwY8R98Ts/Qgc7nax4YEJmfHNoPjp71Ginb7Pq59YeBRwZdExFzHWwZaqATXBJoRF
SvkEaF1upB9y5nU1FbpSrM0oy+NWhBvElIR/diCiSh37PBrYt/ro+EjtCSBv39I5ksh4ldUn176O
xnBDVTuFzvN2mUMlOc1+DGbUgX121uMXrXRbiUEb6lik/8uPqVPqHInlFfriQ0GSJX/0bkgPdnbs
k68FijEh1nh9yslwDeNJ+0/3dukXQ6Z0VpjPJ5LZM+CzrZKhgAwjGN9v7YQ6De+fsLVMrkOPcoJJ
/15YlhJXgE18So747qrLW7FdYcMf+cIbeuGwj9o/8Y0Nr10xDFUJLfV8zhXPE60oFX9AFgZ85fhF
GAQ340YNXH3FxJabHo2DzXEb0uwOGkd+nE/79Kjf8xwXJLeM6J3Z8uLxsR3YufFsnYe6tqb5Uu3a
xK58QqjtHbjIz9+pukBP16bHuH2QRVroRGEqQcTwKylgmBo9aLPxRXYYKy2QsKZXe1S38bQ8nr8i
X2zZufNHoui97mwB1Fs34DjImjkqaWaP527opEBhufLq3dkh/H+0VCog29lC6Ke14W/8UjbBDEFK
dQVHn/2daIqwxyHTfaouofizur/X/BOxMzAZ2cwZ9T/il01STvg6GBht14Ux+XOogvv5j6oy4KvO
gaH2NKps0feg4sJIJI10aZADfurlQsKyaufqw29rHO6QX2OzMDuMXw4Fl41sanV3C5x5ZEn+AxPG
3AZqreNAHz87ndfbq22flH7h4VeeSIakYUo7h2CaaCJzOx75B6pN08nBt7JMC/8yMOzrtlxyBCgL
pW1LoteX1WPZqzynegSpx4FSO1Y2usvVaVuEZ7qabT/QNzz/pQ+2MRZe4yRWTlX90YqA7jv06/iw
PjBV8ipAl+vngb2/IDHg3G1piGQG6I85WhCGnZUODZiB6ca9FaS2wspV7Cn9cQVPoXBKP5NhINTa
HDLyNhyY7b2nZcSprCzK90hZpgt+3sMxUIy5AP6TAPm5hBSYq7Ob4iRgPkUqxx1KgxRXydzfoAUJ
6c23HYngcWFKdaKZ1ODXwhAYu+c5K0kuA1LhE1kkF+UIMLDXt2+lrCS4Qe38APoNFsLzxXWZgd2p
K3C7M8S8WJyojQM5q6WSvdMkQrVg6BRLT1hcchkhJlWIOQpkEcklwZZtWpwLRj8b7x+GD5NkNKfz
0b+MyLtQeyr280nniNDL9lj4Y81EFiiTyfe/YqT4JmMfSdgQkAKy8iwW5czlB+nBh0XekS4IBEHc
hgMeuWk0q4l/KZNy+bWZIgnhaisOo6tR7l5ULa9ZHCmWp8npt2SDhdjjfy8d2ICNF2APcJ/h0/F3
iG4lJ+3efgQTmfrF7H3eW33KOcbRsogj8fYu+WSMo3pGa24Ki1omzQzJREXoiNzE0VcXJW42U0fC
bH0Y0JgHMwn2Tnt4MmVJjuZHnX9P1XwxRlj/N2+qUMng1tt3mmpNlUWzCQzcScWSKUR1oAmOqFKP
OnoxGnt1MzdVlkdXfjYxIotHnAa9JWOro9ztft6MWjib06q5uCfnDcikK8I2gyTNTA+ho8Gpo6iv
kl4+vLXDX8ekLQx2p3xgFuWjFTcb/BO+JD6IuMKU852FYIpfm771vJTXUpUX22LEr27oclMQN/fO
GPdfAL5Rqww78h/qVDIaqhj8IGBYk9ca0CGDJ+xR+nt6kRYc2SERau0lGDyowmlRS79Fe2yuVW1d
IUrOX8zQpK0/tPKSU5D+2ThjREPV5yy4c+KTK+kj6QQVgEW0/dy8DkLmAuUN8CT7iH4wePhF+vXW
xN0hFZqiuWkYCg0LXcpEfNWCTMDoDgPp7hNHE1Y8j6CRHJ6U2KbgDsm+a1iUyDErIffMWbutIMB2
blNm6FJyCV1IuoXoMwrlOPggYyIdhfapDb2/wZBeDCrggAVAI6DBBL8c5ImgcTSZAzBuSz0cgoLl
4zp3hf/Zj2furBaSNsr8LfrHNSyAewDqTeAneLb5qm/hUJ8IJkNWi98Mp+NoZUwp4YthnEmA05QE
QIdQF3GO5pUw7ngY/YyH2NrxW0r0aE+xYJhZ6g6XsQyvzTZEZDohHNfzlYdYQ1gWBw36lfngJvGB
ryEhA7uswOI5VeTti58w6IwZrReFw26NWAaA4Fvr4mQlZTWGnZAMgahe1wAAU9g6CRgBfyP3lkrg
Ble5kRcF9AAHg2/mOCEFT6ELtearoj76nScX2cNywOAHpbYEMdM0ZreQsUDNm7fsFvfBaJHl1iDV
16gq0/nhZG8l8xCdDjpqeI5xU9aWZK5dQjIWX87Aqklbn8lLRP0exCZjcinojPu/C8k7bbqysURD
0YhP9TdNCt4kAHrewn6exIpTLBZO4nlT9uZDWYQHyAqIRHveITObnhHwFkNOaVTglILMYr4GaMfL
GYgBQaD7nrQZc9ItHHzPPYWeTjtbjqVpSBdPr7J75jJsNwLq6ZfiamK0VxGmQ0qaD/KV36v5OxBK
rsax1svNEJxzyKExQHfDS6z3IUIS99um6Q17+drOOXTEqzT6Svf30hQ7ghThk5XJEsh+TzUBUQKl
TezzL10qkmRAxrt7Pzx1pyF8Jn8XetFfldbDInn/fD415rUyDKzFgCkE4ftPJkk5rMpRuwVGWZnD
sbNnBrfPs+cetQRV8Oas10gMhUSwvyOT4sgptYhPmv09NOCFWqkuMdVvdlZ7rC271uBAJaTA1Xka
6FexMkQ+oyz5eLiTVGCHr/+wHZZIqncefZMYutrSAw7B/FnQcaGRCTVosK+iXxhJMSeJ9xa/S3Vb
cyZzoPx7G4FrEU2tsMjov8BE2k6VJkLNIoZ+HDSqP7UlqvoFjes0pKnajLM7RSCmdDD4isARMovE
wlrYwxqG9LHAnWJKMiTKBlEzxE3E3ncYJfEeum/jl52RV+eIFluYAkWLERmE9Ylt3pM+BcX80kGi
/clFH8w6Sq0W8A2iRmf76Vk3AxbmrI9lyMHwZzYjhd7w8RT7Nt+0ElY2MYB16v/QAskUpTPSgxUh
eOoFR0PQ9Pq08wO5w6juytENx5z1EaDSO5mnIaGTWV8M1PbheHxxaZa35Jdn6uM7j0YhO1G/Tig6
vxAPc4ZzFXWe3gj0yjRWklRdLEaXEmViJlGa1LA2XRgEdvxWwcHq5lBN6h5LenegBZdPXHLyno94
pHizm/lBVD8jEt4uzEMgsYZQ1ZiNCVN5Q+x2NGSVpyPirhgXkIMOtepLBdJ/gmwveZvhJfNKamVP
/aKDLEHIVvHzgt7t2S85dhw5stt9lJorVEE8stNjZitG08kMbpzj8p5oJYmWrq+xhPIcJH+YO2wO
Wg9E0yOIJmJ2vVjwJ1HzgPSxmOBLRzUuMrRsTq0g5aHujqy2kX0FGsR3lYAn6ktxmwhKxhVt9v5x
VcTSgbT75IYtkfELmyd7q5w3ep1vSeI3SNJkt9bHzw8X/jAOhyYnvMvrR+qwsq/2T1VpAzl6z/jJ
Hd2pHRQqjoqulM7MuEngYBDkZdsZkm2R/tLl4YYKhcMrzefd3BQZSyjOkN3vLgKUS5AFxpTUOHld
c0k1Banplv7dGtu/AvD8mBb0/0euWprtm34nnNEjrBvHDZNTNY+IzK0YmJFLH5ZIdjVZcnFl5V9K
u8pnWmnuXZabTqwOWl6QEFkdMdDQKY/u1ve/pGYJcXpaBSzgvT4FbM2Vf0OBOnboxjd/yy8m2mjv
MZycsbWOnfa1ZDqo1ChfbcZszVJxB4bWIJ8DIeJMTFlt7CDDjopcAaU6tLhC07XLZi4KR9380DDX
nEK3CDtafXArm1OzPzcorMx98U66RiGYrfjWHJbPv6hcy0grMFDVEIX5cC/9rmNwOMYvlX633v0v
8bWPTCclBJ6VQBhQIiaMMKRFIH9eJxN/4x6ea192K5i1JGuDhSgx9hLlhqGJXbtZpbKbzDBKz23c
lcqmXddw/tPIf2RSyA95sl3Pagii6474KaiX1l9wsSAoqiobeSD74alhKX6tkFaFfYkmTC+WrfoS
8N3Ws7ePehWCVXeWv6G3SwjLysrOb+HaRovU89X0bzYGCUK3tK6rvKuVFQFk0+77omCB4FwLY+Zm
XJYIoDqA4J7PugJscBlaytAypSRViGQKdKITdOcSo/UUAtdnwFrtQDKKcczqTnoJmNbgwlH/qC6K
ovZkilhm8dtQibxcWBSYhjBM2bWQ4j9FaQpXJvLydjv+ArTVYUWEMiUpp8aqxSaCOIYe5uhcuZ58
nuNENW2CChuuFywcM9Ez6qixiW9X+J72Kt0PIJWGYNXaAZnkF239PwZHfRMFwESvuXC/2d2gtUkz
oTQly0X0pwZ54KsyeX84P9ZR/iOy60dOSlajTdGAHMjWlqdS6m9CDhUvIgq6SfBFxnfuZl3nImZ0
7igg1EblfR9WhrHPYLQ8BCnW2q5lO73F6ksfdpLwNQTNYgVh76lxUYXi/9m/sNJWPEq7O60/QpUd
IDQaAipHbJHSVvB85hAjSze+ODK+6tf2l0ork5/7cx5sdRXnyEmGOHL0WxqSEaOmSsZx+e2B1Jk0
ujxsA4zyfXeSfqUbpLsnXOOD/OmRNVC4izZhqgoLrpe0KFJqU1Y93QcHdEbvGZKgeL9zYHbjjvYE
6EuHQQ/+zfh4Jrr/DSz9HKZw3VyALKVyOTa5Z/OdYtDFckm5iJ/0z0rh96gpVCwwaBWLJltuphRv
HPw1FDaDklHc9izmcwxNcsG1KNEfFlg3mplPJs6imvpTEsOtOGHqTJZrL6ACVZELKO2cGmMxLlrF
osyhHtacRcq/7nJGE3c+rv+wmdLU9GKyEYOAho6wcl67C7/oUdGDWPFkPdYRzB7h2nNJWaw//wvj
jkhf8DYwJke++lcE9SlsMT1qPcWIRoFGu45vbRdQ6cdoBBo8DIjh8IcRa5T9SjwLhZVrCIinAR+R
DsB66C/3eEv7H0e4gwbPwUEAKF2+JPVgekPXzfnsJPAyrq4GVxjfcYXkIUOd9yj7aZI4Iru7tUmY
+c+cbqxaj/OH0f4ML69a3IIltAxmL8vRqtfZ0Vgr6d3h7S873AMayV0Q5sqkZi9AcPIALVKjCQZv
DI6jRt7+YT/DbU1R8M3kE2A7qEVLjNaa9PHisv75UHiC9mUtsf74LOKEc77am03dPs0zAY2OKof0
iLo59V/WuVIXRzBkHIEHzL7pXki50bqb2gxEvm8My2W4319sGzYJEauJh25E9iQQKMJEK9rkj9ez
fnpIB4+Oi6iO8R7YZ2mQdMvggjB0QmVvtx49xkkAFmTbQLZINV0QnGLY7sJc4UgKEYD9TByDeYn/
hveT8K8AHlEuuspowLogl9ST8JTlKzoB7dAkuXo/HEfcqjv+pIRuKMXcPmcyeesYU61xBfBfO8Rc
NY3kB1mfguwcLSUcLspu9N9Ow+kPOj52P4R7kmTrHeI8Gm74KSUoZYcjwYvqwIpb+041gSkAbLLA
+j1a64xrnjGzuwULGHu1z0ktxmaW2cqxw+A717hONC8y2mGPbKUrKyGx34iwyAOuX0Z28cq6JUbS
faBCOhRxnqg/rp4cVcGg0B8BU2nxVkv/vPfriysZ4+Imbg46+cNQaEk2X2WeUIqXuekib79Pj1VB
KbOze0SmJvTH225YBfYz4iDu1IFM6XM0wYGZp68xMwKsfIzgwAsz9sk3B27jXFYsTEC5nQijkvD6
ChhGByzuwdMlllruAfc/CbN5DoEclxKDkB6+eMEHprAy7lzRAAWQwYFs2WLNPzFwMiXA07vrPBNw
JYOZTKkV+DbUXlSN2r6ZQPWFJn8rBU0ZOUBEAWKu5pO+br0M72tCczB2OdWSukfhVynTGsQ15hPt
nGF2s9wHPf3H1HaL9u5KslwtJnFejnlPFuOGh41scoaih9hGm6wuZIgKx7VJikwr7i0RtTo8e3if
BtUaToUaxIkKn7QMLXGAp8HxuQmxsuOns9mpatBY2Vr6PKsKIDXFsPQSUmspxLjF8g8EN483qAuE
9W4z2rK2iJTgvXmsx+kZadWqsOScnIgG8/6u08YKMr6y6WjKKCcZpL/PySkuiZ3TZWAEY/0j872S
GXw6RnYvUeNXqJ/k2Iq2RY12sFBwUvZqjG4Tlohx4C9pDd1pS85wNxvgXXaF/EN9TDwVH3Kh7TGN
Jvv/ec3Fa0XvEMEl1sEf51h/kmbwW7JzIWAI7l0+/uuOtTqMU80m8NvoizflDUPWktMcmUrLRk9y
X58DhC0f28Ieh2V+tzKrdf3kmKW5MpSv/2B42SRMmL/Xlg6sfrbUKmckNMABoPz6KH2n6wZ1EY8K
YYRz8T/LDX6+Ui6KNnkyop3iJT7WlTymSbBG2lakoAbTms/ZP9aGijClS5SDlS3JaAWPaLyHAtZp
dsWgMyBwOhdDOCpSPcdHRneKEY0dLM+Y3dPv/9i99FS84w6q9JDF0z6yr2tACwYGyUUPkwVvXMfF
J7jbAyx3QD+xWYqxGfWMRXVnJr0Qy03Qn+GUgYnlZtG91kW+pixQDbucPub2t25G/afSSZS8YM8C
LXLVw/W/3iUyjQBxkLwh2x7jQfa/Ez9unWWhI9S/6QkPZiDXcs/7gmIKDwsDH1pAMxb5pxtFi1P6
xOLxRui5NZDR2JNdFlDkPNn7Cndn8VkKDE/mpvemBx4/P6xmmfihWkcixseBZaflWTa6orQoSkXz
FD8njXVCwZ6vKerdG3esKTaSAiclYrmxc8VrBCII1p/rJU1j594seJGnwkmc3qvT0ulnworUHhKL
lbm5dye7Z9t1CmkyBNVff7uuGbW2G0y0G2IvhigciLTxxX6O1MVJOpN/+bRmpQmIobqPmUfxF5bm
lHI95srQN2K38C5yW4pq6sFQx5nFK7aPtalF2S2LTXTkr386Xo1oVVK2yGh0vYCa60PZxGAWDEE/
0G+13xecRV2YkwMyl4AnRQGMsEYYIBWxzMQgs/Q8Il1FF7nTaNTnFupAee81sHij0aZi5zY+wW4m
meN3eOgRx8ZrQV8KSnYBzD1JNoPFh9qLzzo5XPdnPwCRRJBjnZCLKOTLDchaQQJ/UKniYAMQWg4r
nVk2fX2Rae3P3/Uiv2TlGVS/LtWHLXDr+dhz/zU6/niIV77dSNz5mfeHaQvDSDiinZaVRwWsTeKV
HB2qMpWYqJ60ticNj3u1csPO5pNDSS7W6USQAU3LRfN/bl9sRRE6GncT6jAHmPXUKMwK1WH48F3P
YuFw1N6UCjc2OCiz1mYVQBenwdcp0xhWXTONTm5vCWF10QwuMG1VXIPdvqtjkzJQFE5O1BE+t4xE
o4BBSzaxKYnHbo5KrfQUK87oTSp+Edw25JvlRnEy6gQkrLH3qykfuNOBq7zqHe6sop5GTHmGtwyC
u6X9178wvsKbT1rCwqp8P0xTUyGb52zZ2+VRjWSJDNvb3jPsIxzSCYemjp8GDiiJrMrrlFE/6apd
Tzi4Elpy7bZZ6cg7g5crDGfl8YeCBkMokF+vS/fucyHZro2C8ighTBVbNYnSi64phaI0PmOmiyDa
G+cidedKtoB/amZOFCOU4jax68XrvOSsN3EycXxIcCil20PBDLpGgVqEYXLC/QzlB+gFDbm/zLpy
/aHTPdkx9DRW4qQnQ8y9k1/hYh+7u474w2jBY0kWj2pFUdWrG7oDeuv0W06gTsOGprcRXEe0xX7J
fDpRZtgjl2sfIfbqsZm2CpMMwATKa/VqSRFRmMQ4Qtv8tu1+/OY9Naj2+34M3AR9i2tpmBFlHfYJ
ODxapsoIQpCFHHscDosOiedvGYoUrX//9+CR5Ey5etZgBv/tl6u64/6pF80F0ouGv7ZXbfiWoNrb
PEVEsY6b0kX99dI6TQh6mQCE+393UmiAELesMdkEBpriZuzdkvQu8JVcFB4gXFk6SrouGzXQhpfY
iKFkaFH40CIFFcem3Wh6PK+ATdI+0DxKSQ/YzorAqT7FQbG0sQcB+dULttwnGV4ceO5f3HepnzPK
2xw7vef6cvQYqlQwJtW2api25AHWylT20vDpOLrXVcVLnG2qCVmv8rFTyJhzJrBxducq9hE5Kr6N
EpbzzLvyB3x58/7SlBrXqZdY0FbItP5/kGJ3dSjrTLyNEH+bWzhkSQmAj5QmxrewR0ZydYxHN/J6
ZR4EdTNJgsDGqOgJWQ/OE2K3Ttw2/whGTZXjAfQ/xef7vK/Ezab5kqIqpTVVkdttNJiaewR+/LPw
iXE7rLCHRmhCwSlSN4wjeWSaRfsXYdn9EdNAQniJXr7N5Q7xzPKS0MXI0051FnjWrv7kyNSlvJE6
y1Rcti+lKntIn8gHKqGtPhYQiDkV4muxfipOzu0RO1lmV7rqh0uXJ8sGGHKAeFlVkgVK6JaRcsqb
UANQhMcyvUdmkll+26cYV94IpwjVdLebx2BFkeUrE6UMtVF8GiV3m7ZOhoTRUsaPfPBTNhByY1xZ
yfZ34knQw5oSgdqufOlbN/2F2i+1QjF54NnJzr4sD+rsjLysq3TJP7l9mzNrhsdHRhB9YhTGlWS7
x6VcLDHwr60+3R6ldmSSWhrVZrl2uJRBau5DDTuq7EJNFJbM+6XxLu8bgcU5cRhS4wyKYjguGVxf
OtA5yacrbEkuPf9BLvApCbAiSjRAvQ1lsGCYRzGog35w0kfursgIHnxP0786v4jRgIQJ9pb2v7iM
+VswdDMu3R1VqaWKzQnqBM+ZbRHiNOZ8WyXDLHeeiMY2wbBvIkNRbVe/jLCal+UM7MA9OGx4ZTWY
6TOvRKH7HvlncnTsBc0Dh7mdh7qrIF8xJ0RqVGBLNAu/ncIjiN+HIAC8G4b+0XeG/zDT/qw2IbvR
bmDqGuP0QYnlFyG2FDE3irloQbe3fFRcP3F6XWDPZqVGzM+Blm8DSdhShvLlcFIQG4xzxAXLQlLI
yLTo2TrusRP5nExcoXejLs+bdpdv7stlPj1qrPSwZa9REnZgViN6E8wjynxzjiTwlssnMXNDLYUU
hN+3+5g6EI63p9fk85rzf/8K+6IAuJ0QP6JNl4CJbq+/LpSzI0EmoBxvlZoCtmEohQRWmHFKCpUC
2Bbi9rGDfzUbp+1FGd1WdzGynyb+ioXeviLe6ziOeEegb1xUdmX20fxLJ4biNI4rHIgNEPudCQYJ
jhWSy5LUga1AvCRwVh7lprcn/+e1kfyKW1DmnMejOohoHIE10XZ2wbZuFbCMpDVXdnCaA7nFrjXI
RMKaAJTLvuEeb7wENfmvuOqTRBc5BYVz27pANq+kccCoCDxUlD3DktmRp0agSAKqkiSweyN9brt+
dhmzzxgXT8PFxvsOg9DgsztaWLPWV+QoPHzaDJ8L7nzfrAl7f1YMolcBwIJ/D6IjPfo1375qRyQ9
3HZOdcG23u2m8Hyxb8M32CzMKCKvmnXdSilLsJt7/F96oF7FmX4nioUWNzlMdhEKPmFatiP7AheY
WIQ2cX3HXnE2MJEYxDbOjCCngZUu/U3X0hcgnlXfiST3A9xkRXmUL3fM9WX15x1Y3bWIMRuHuRVc
6NOegLRMk83VMDx1hYuyodPmxRYxLb+OoWarP7nGIv+ewWTiCA1Pd4Pd4/Kv6ihZD2WD+L9Acilu
TFqRj9vCfPk0LdgCtV4wRpordxpCwe12SYRFi5SsanRofdlGOIDyudAjM0Y7SM88xuq5MTWHPVKg
6JVqGCpUYk/GNwMo+JEvmrHTlUvGc1aGpno4xVAOQm2fV6+Z96CXgP+P68ou7MD96XlNWkqk0fCP
8t/+pkSfTrjBFmNO77xcudWn7TJSmnTfe4UKuob01Z8XFrNgSOG7ZqXxdjtWK3n1J5Iw5lGM8Ww+
y5ciIpGA2ajGCFaGtStJsh37cHGZonVhTv2p2hB9/doVAcOrUBrUlXPmE6h7qbRaS4yzsTRkg06B
0IC2yhvyv2xRJ63ZujnkJEy+jMQ/iGSZD5GzkBfsXgclkjOTtLAA6O4t8GzTY+MKpqJDYDtYjr/e
z4wuqdtkK7AHKLzi7gDXwsRLVFkgnJR0O+yipCAja5FEHv5x/4YPAgsVmKEvJhTJIYfQTghTByt6
AsVpn4JwTZR8VRUVQ8FsfJKL0TkIQ2Ctp8B7fppC8hR98bDLt7IrKM1zop6QJ4V3Q2lByt9ET4b5
QIRrc5Gcst2+9J5/FQ9dTvk+Y4QutgeW2mCnQcIwH00pfDOFubys79wSroG1o99BOOTqXRFeGX2Y
xddvxA0OO6U6afrDysTpEun47hO+z6fuaX9hP9cbTN6/ng7l+PdQTERBXUfT0teqDZ3IwZf3RaEM
42QBa5CzmLRbMDxKCWdvY4jlqh0ZYuK6uh+pSX0kCmGdUXJSQkRk80osX3Th6LhJfz5ESXgI18kW
sEPfmMbOxk96eVZd8mRN9+FQlGSXp2Z50F7d5RUVlxjzVy3rxyYtRYChnWK3IAZWCqdNb4A+gXQs
2wSGMGB7dzcULZGPjxoyMy37xshIG+QJPAbnSer855pOdCqEvFADm/gv4i5z40FX/GbgM5w4jUnU
3a1RDTHNBjQAlFfQoZCUleC75LmnDOKZd75aJ2/5Ofg8FpS+SqhaygR6NAzWXggolUVfdy4RK4QU
ScgfZ0eZRgA1vSWVBqyZS6+vL9WsxUInEdQF1rJL3Q5RzAe+L7zwutJdshm1DQUVevIHQ4uwGAu6
VCAHNdj1dAVvosNKRzzjEryBljl2APIImdnIs+WXM04x2Z+90i1JHwI3pmXN23svQhXUrmFURZx8
+JZp4Dpm7x+ocl/HOZFeysTL8uiX67TC3Aq2dGQfsK7hS7TTsiLMi+e0dIBiZ1cWZyihIrfNTeeN
aUBqiRfbXchTGoOZZYLhBFe9YLMBgzsiOL9gLuMwXMbm040AwYygrqn/KTRY9ZyWhUcCUQse/EZA
f4ulv0Jb5R62HLG03L8CpWTiENk/PYI3r92ttTdPNG1kS8lkWSAqc2BlDqY7bJlRYiBYplCaNiOB
mpe66bdJr0hAEusqMqeSxnSXexsKd9BMmKYgzmBx0v4j2l7OA4tLFHYbCWvQKv2Ag0dF0kn1/cnn
/L+Ywqz4jXYG9v7AWeQD0PC2GTlzf7hqc9Umlj+rKZWcPkgaFYpJOWcPYChtbv39KNIhegw7abtA
U+P+EuaOmhPEvJcRtbPH62b5aJIn4sHqjp2tbkCHw6RJrTljh7pkTvJnta3ohqMsbRT7qCInOQxO
yp8n2mmOK5g3tteC+K1eCGQiciJmTxeihEOqw3g0s7Ib8FvI8WsF7bzy2bpAUTTZILgVJWjiF7og
9LCe/lwEGrIQDz2jzwxqMvqSk2mFFqcKkrevBdrZejJmTbMxytinOn1J3Xic7JBrFHaAQ8dXXbfw
0nHiTWPpKQURSOYpvZ13GNAJu1XFWlh3WBE2RaLd9b+1FdI6UqDS772gDCEdguORDaLsdnHP6hQ+
kfh7aZdUohaw0OcYL2TEF5LhXRbl/Zqdcgs5F5kV4WT9bTwfPatxIcegeXSSOsAIeMO5+duYJjYr
6aOLugStAwoJQjnDPAy/Pu0GOMp2Y8De504KNbjuMKt7ejs/W8nKDvpQxpqBe2py69+Y0Xtca9ZP
zBrEV40QbibptpwpnbPWxU5HwllqK4SgcuUVu0vLouVJ4WF6VIR+oDqv6a90DAx+h8RbGPGnH5xw
iO8Z2+VWYNtj3y8YRSgnKCfaN1kcEfKqvu3bQMXP4Fia2CCYpxxFKdSuZR2B6agtNDeUnkYF02WY
O78iZj20SgBxOcgozMtRl/Bhi/rfdgAao0q03lDF/EV+CysyCGT1QyyR+qEonAs1F3ITXyBGxY0N
GrcpW2LiN7/4HLBDw8m022IBCb2pHDW2ZxeKGn8NNyAEsd9hwsw+Lvv8FOWiXhUt6IcR9+K+i1Hy
oIcAJsEuYb+Ra2jkSZXqAL2sGsU8b80x4B8BE+Wv7M4ZGLLoxR4A4RdCezhMgGqwpr0Vn+XYDkR8
LwWpNg5jov/2lEeRMFjQHF8apSlcxes44bGYom6Qg0O8I5jTZbJSZ0IGFKs1w+zF2JVqag+/pBg6
9U5Cnciz+84fgNBoUtPtaW1K+6F3WBSsNeU8CHlTcrilm1JQpr+0uB4E4R5qv8nWeXcUWDZ9ycGf
OFP3XcYKosDelpPyuOzfymqBHzKhws8O/cDhoyFRCFOcRBcMzM3FDFV3HYLJPiqs4LYaxp9XP2jC
9ERzvVGW73Bbkxw7Cx1APN/M57pQGHKS5Io1vk8FsGj/MyMVtXn9PLUOP7N8WkyniV1pc3Ph4wi5
DTmDXjA+xTaK+dsjjvq6azfpbGdwpXF9HmP6XN3r4WEsRcv+c2EPkroEidG21BnowGoimfD7nW5F
G0mK36z5DNUuvZXgSSIdaIKryzPB36ROr4tHHgIk8F2FS+/6XE2j9kwNiw1thCnR42NQG//zjh6a
WecxvLhqh1yv3tj4xzX+RuqiIXzjfGnS3oGj+SRBsAy4yDDCHEm3trHZOA+3alBsugV3euevmMyz
qqja93yDPVFbwZSOiUjfbF1l1UuEKM+q9MJsLRLrpsCarzKXZL64g3khz+9d7Fo3TCp7Ypzl/0I7
9gj+5Biss50t5QwdM16x6Dk4POvpQbrX6bvyh8aNAjYJqUAIxobCY39byRVFm0pLAP9NA2SWNROp
PRZxMBmEhp0nRAqc4Vx9KAl1gANYXIwELpADAp3+vWWc5ICRZsuQ3L5LaukPxgPqSuquJIPJh4kx
oN/d9MCJjcTgU42oBwOr+o80aWbf9ZPCIcFjW45mJNfJf5UXI5WCHJGmT6froR9O7zPMBrmuF6Cu
YG6fwkARZkfX2FVF5vR7kbERweRmoswPyYuASzmV4MWig+2IjCN6GE/75mozxV3PI5S1Z4QCafzK
wY8VRfspc+K2lLJosKK5dd0sPVsoA7ZyY+nptvXNQOkOh/UYQDICMsyl9yVuKGWAOSV3dsx3yeCv
UKlURcyk2JSimzElpuk+HsBDExLt2KuiruisX9Qtgnzy1/P/28Poruf0vVrmK8dquNjlYuGlFSBu
wTR7dsHecXWWFbobOaUvjrKZM07vQJI41OvKvZ+IqO3MVKdH0kX7793fZ4C9PuAc/GOR+7BeOUES
vLLjASQRG1NgxB/1LEN9XXU1Ywslb1EEiTf7219MOhAI8wZ3zd0STSh5xuY0MgAeqBJN5GZ3gVrR
d+nx14+Is/uGh0M/uA8fDdVpv7gR+j0n4m9vw4v9B0uZU4kdj72LxnQfFCh2zaGmaLPDRuddwar0
qTXfVWjIds5H3wxsOJeKRgklsuCzusKaRzOAHTwnAtmcYWSO4PnSFj0YsP4uYkQx8v1FJbA+C2BS
uluO8dGVwhV3PEgpYKNmzKlXLUtGwttNzbw9b/Oy9tYv9orVJxjtFwFJlvQ+yAV15MK4z4G+7Myo
j+dvnMuhkO5pgKb6KvMqVW++WElONqQEAeOBGHN/U6j+T7IbItY40v2kwMMmVfPPHmqQzIHUHnDU
CuXotMaAY1C8yx0LpWZnOG9zJII7kEV7j8LZbcJSVM8Fhj+KYjtPpHKnoxhWr/i9FXwGZuGh7oiA
DjJh8OmfETz6/ssgKEr2niY9RZUAQ57U+UHkg6CTjsRPlxyhzhVrQb5lnNUDfnPBH/g0K8GI1Wm7
gJSKbDet4UEjuGiG2R4uL4ByK3WP+1lHdzbWbFYbg6q+cSVDGnmPzpSTACvuDRriBumosnLwgv+P
x9M+BC36emtmdOIHZvVZJk5kE9QP2dGaJidYWBJLvpa8DimLm2j+d6cQWgLkqMWpPRAQGD5ZGQ1j
2luyGo4gK8RTkl0+8L6k7qYB4acQ+2X1a9AbW0gz/lmyfEG6izcasV6B1Bt3JLvMuHRhItVuymLl
lbU2FHsGPQyP4pzcoAOHeYgf3QYwsHz1EI7FwjhaK7IKYobPacKiVk98amXPF6esgxJD0VvJFSY1
wSyYFQwyROJVAObe/FEY4NIo9ID2MVUPZSz/kh5N4xZ69dtdlrddw/t9VreK4jTCVDJSDI0iZQa1
7XsK9EF908il5QPZJL5KywrlCv779EquAt/WodYq2W9TV0C+waLZVtNRXFkYqJFElsKyB76NI3nx
h/2DtaGehB2nyu3+7VbFtKWd9vsKW11GQvU2b3Cmy8C6ZGdqTMbO+W4Sldwt74kK3aBx+wcPL4j2
ShMPabZ2AqoGItZ8Qp+if+DaYnohB5myfi3Zhyk26/Hiosa40o0sZwOeR5ma4jrIXfQh4toI/c/o
BMbzTh84M3WPe3aZZH6hQrcDKAs8+8zLIpsneuVzF7NFpwzUbg+sWfl7ftuZqjAWSXCw8IAR06JI
ilZqyCVyB8SHQ9FCfLtVw0dGQj2DVIZ6vcKLpZIUuwzNma9m7L7UxbMwtMWGnccLQVDncueRlr7z
bqARdE7EMjWKeM1bybXheHlEPqrVw6zK8FPGPy31d1Grd7YOjrrOLz0U5tgGV4yuGyYPUw6cAS4i
+4mA9spZl5881VLoI7Y5V3d3f6XsoL9yG9bt4huatadj7aMhLTEVcE+rsWC5TVKqRC/ToAVBDG4k
gcldljeZhgN0BdHC2EpvY3VpJCWSsmJEgoyiO4M/NwuKxUeYaep6WuN1/EsM2OtzJOoKqoda6iF7
cRMEo6TW0E8/VXJEnEv/6PycCVW3h6N0y9fZNdQhcio8OITosf9XYgB5gWldCstOm5e9N+B8WCHF
OhaaogRs1EWHhMYxixpQ7ONLiFUOtnpPAX+MH+DBiF1tXfl/R3MtgcfXk5H4WThwCLU9yKJnxqzc
RLemBceVa4ylJZqpd4TjXFjtXnp9bQt3TAKIz109yqCvujqRsy+QvU5bcpoaVRqsfocVAlXf5SNv
WjcLY33Wx85h38Yr97PofG0T+NXZoNaPqkuzJeaofhqerG1SjAh+SVpklVoMh1V53QWYHfVwAU4t
UmFEVi+isUNDVmlOZd2rD6MskPmArCwb6kmLX2WHx5Dl/Le50CTY+NMC+c5+pwiQSrXaBiU9+mxt
bLmi3eLjPJcvtrbso8GU7MjiExvNoNQHaMafAxmnUkoyU5khC7MAsE8NgLhqi4AMR8amsyIVWZHx
6Bv31i6EOZJ33xvlHSsbcrF1HWnqLb2K+Ar+DmhLMnf1fIrPyzZqIz72oEYLDM79JeN8wN//31gm
KK5oTSwugoxi/0yxmvA8Vu5UdcEZsZkud6E5Ckpm10MvjsM3cesUPPeqH31q0X8l8zUan3Z3FyYd
01GW/sYIDNrm9C9tA6votvPpBSTk9sHVM7hYTK+sz/IODE9R5vfGkfxVNmwkCWgflOVjsfGbrEAO
p9XdXn+gPprskZ2yGWdwft95muziYomqGLEfdcYFeRMH6oHWRKzyMmee01Sfrj3GIWjnlBGtM71+
DPGApifpBJOx7ur9K8U4c1Ccv5vRvYjB4nW5dQ6UWwuQI9lirtVOsNYi12QgS7uRhc4Sgf4fDBsn
mbN5WOJugsRW6wr128O8wXcTebmK7TEYAzU1ouVn2+iLtQtc2QI7myHYkmrKVmCpJaL9jN6coLB/
sk9ep3qjyskFitwMfw+Whv/8cjgW471LieYUP0M42wXrxlk6p4iYzxq4rYlqu/KKYKStyshdWqYM
0J3B3nTNsLco4Z5T0zXknfVkUJOA3jKOfrzxo1xiFQdtiH13IVrqkVwz0orscOrbvEvYEmB6B238
hh1OEHVpl4n/SX/4KCJANh1LLpsq+0LfnBlosKKk+bzlfKl08gyjnQ4HmiUs75nLERWBEp03HLdP
ob/96zTU4ty2L4msEGbhx8j7Awjg9PNVDWKDF4Oy1XNXFkurkdbFFyXSlRHbmSvxiWVXkyO2wnK6
JiSkcAFG1Lz+1fQoa1omo/4neywKwaIzw82ibDeB8zBiIb/zj5oBkhZlGJtujlpCqFxcsCoeyf15
4k/7/5wnfAc2ngTsduF+hnR32Q4l1gAf1BXKbsWbWtPg+HZauXVz9th06OgQ/lKvKSbkE9Trx6LC
gYfr1nX3Cv/h8O4FmrnQf6NI7D3ycDNzz9fR8zm5wK8CiAQ6p5cl9JmA1yQa8tvVRHDOKuvTT3jb
L2qq+1HhIwZO9ImtySVKoZLBvSpJ092IB1gpv2X4UGbz4ga0dCQtMmEdaZZ1QfiRjNam9EDq4OdS
GDtwDnBQw4k+7vdQACPpfMzZveQABTvWCQ734LbPGd1Gy8bf83eSbaDZxhpouXWA6HtmjiXR/JrE
GCzU8X5z6M2Z/35zlZT2XrkOl5yhVzEFgvqNd1E4+DSOyk3snGyr+JLkDGwE3m3/LVcXQbZiIUx9
WBojIn9EmR8AkJXyulS0CUxfgtDWd2VdTlEJLJNpQiLq3bfpUBlvhjPvWoHcb9nNmLHPl7HEKaYB
P+GBxLdip1gfiXaxQ5Eox2RsDNaKJno1MdOgcrHVjAnOuJE0kfXU0xG7XdGrEzFY1XCVoAh5uZae
wI8OXm3/QV14hkvULpNQ2S+8NSB6PirAtsF3MDodJ6gr/+NZ1VGljZjnxT5lkfgCOIpG1TDSKVel
Tqs8hmt+wgtz4bdacJun8kNAmZpNwwyNC2hfdFueQo5iZd6FLL5jI4deayAzBBWmzEEufyE3FuVD
LgodOwPDeZZLDWoo8Dop2bCSpc3vldCI31rVvqJOVGdrT/I324cLlaaBMGr+S8oHe4HOjytHrFeH
O33T54eZByVhfsoIPEDQsdTqoBJuU+z0k7LmCYNmqSfvyT64sO1HuADOF+/qUP8EM6lmNAuLvC3y
c1e3X7nyTvtU60iDcqRb6aeMUyM/YhMnDIKH4e729R0wmnGRWuF7CSoBZSV46Wfq55CndNWr6Epb
ntbEiDO/niqrb5ODf0OMso7P4eh/duJy2DYxGwa/N5N0lunajeMTaq2Hk1n+7qk8GNoSNky6x9TN
XVPB24Oh+cBwaSQWk8zdGlUr64Eqe4ojQ1/h/y0yxem5qgleuDSBRm6LQrRbAYcOmCo23Kr/Sfo1
Ong1BoNIPJoQb5zJHroISOgIL3m+mdI+ZwS2VwMElsaGTEmk1CdXJatFHJUDhK+c4RFof3/BlUbD
xMMZfzbD3gaoP55iQeKHqf3ueQgctvEeImsbn43Fw5cYV8dpBKtHWe1k5hc0b5SBHHL9yXj2lxe+
7JnSqOtFJUoZMCXynVPZg1EMEu/5I5eJjwCTjiVuXfXIgZEjRwCjKnYmxf5TRqt6baLD1QdbcIm0
xvlhIqesob+X7K/htUMGHSL2Q+TY5S7zHjNiiRPpA/i3DZRllwZkZ6u5FPn42tIgddTHSEIMLD5k
x9GSDBaWDx777jg4nld27g9cD9Myl2J/SgeOoNLAhXrOV5vVuHsKF4sDhtTdYqid/ykxxbh5JrBo
r/rGnt5hysCwV8Cp7Q+bgWHTFZauxpNZASnT6OgoIJ+VX24+Uh36gfeeKGxlSDL+JKIcRCJmeZmo
up5N56rGU0A8vppJJ8UAW4XscidT5nk0Bd8aviu9bjAE2qv8Z+kr30KtbA50zfE2FCbVkI+IWdOy
lktbkVUqbNwIF9YEUZVKsnUYgHOLJGtqQwVDEuYjXQWPOjh64FTSUHCUyOzzOWeDIOZRcDaWDGP+
HKEzhfLDIkaMDMIuoaEY7+4QodjVC7onVLMGMZoDMArO5DtD/pgoT9uPahFrsd4Z7trqx/rhPBRH
uKKGCPmsCYfV8kzkp6eRJYH5cMoOdWvsA033nc3rQYMWZA+HmBzUnw3k+GerCwW/Crb+JhOtuWUo
R2UQyFjKlJANuJL4nkHtFBSsFa2+m227OB25eDzrRk808EGmvBookh6G0FkC1qu+D30PUrTynZAY
2IBkoWbIfe0K/7zefrzyOBP30d5jyJrXubZUaOcG7je4G4x6OdMrU4Ave2wQRFOn1krD6ArkdqVP
tbqSPGt6gizlkUd4LVCFZj7ShZvkMIGindwSwFJv1SiAjdZxBt1wGcC215rw+beMAAZpVpLLwgsK
P9TXng1zeiQu8G+cbUEc40viBDFG88+MDus/N58663pfSGHY4Lwfmb8d7lk4IDJ8h72LQtOMurEG
jmqpM/t3WGmVdNddF1saDqSLDVJrIeqdjNrqKuBONaOt9JoNg1T+xI1LEzqRRFFHwioexElBeA/Z
IKeuAsFDlyG/DMqzymoDzJMuGWwW55t3BqaPZG/A5Oo7k+A4dZCaagXTfIjR0F7ZkZW4lcU3xHiJ
0zyTk4Jrfysyt4U7dtyBUNJbGQ8i+NfJOSZTedgWZAhxVlLMwQfbJL50EvuXQr0CYkOjJ9IdmZLz
QFNLXv3fo0oB65GkgcyXpzi61ou3vyNQFWakMT0XjAy6ctGmvkgZ8qZhnVvvwOZaRsmkkKFp0nqe
P8sS15S7SZk0jcrly/hjxZ2xuSEj8L7St8GagyJnWOgQXjvFnqc2FJcqg9JPaeZW2ew3vhREhxCF
l2MqYreLTX6vK/VPuBc/gU2j6Ry98y55uC0hjbGhcxu4ertLR0V90KZpYAO7NWCrZUF5TEbL9VP9
BtSFgLjW54QFtB18IHRDeNXMyoAXevkrHXQ5QK7BRWimK3p+Hr/iArADvvcyhPFOnwZejnRkTVPQ
AZ3VFFVG0MUHYCOFZJdNg+8YihoDm7LV8z3Wm9nZfNW552nfiHTpLygA/5YjcUJtZUzvGW4kYwXA
Jx9PeeO1fE312gYujB+7sfpg0zovckamY063t0R+T+Of+BNHbEg8+G80Xzd3FMpoU3MvPmtLYK0+
WOQatlvVL96EddFy95a31pA3PwOvEKKjXVe7CKGBI85Wp72EKSvYSxOEVXsRNALANQnuraCz/0V+
X7qtx259DSv7u+ch0iY65xh+mv+/RKHyzEyLMLqeAlk8pKbuuJ/dnsZ0Wxzjh71AoHmqcboiKacg
+u5l4Vtg2X9c2EZvESt3FRbMApZiJm+7JC1pFxO+AMpkyiMpN0M+3GQONSJmA5oUFhV1K87B3XKG
DF5Mi3d8Q+XjDPa/fPTaeWQ6U/4mL9OQEhrG8tudIQVhLw6va5uUFANKH2R6lRCEM8fR7ougfXX4
XOWw6UqgwpDSr5knZQvO/NIMwzcCaeb3UZeyCocd67L6soxmWE1oKrI7luE/ycmxti3T+OlD2tFl
VaV3176tUMcY+CmSQiqd5ukcia+//GQBmumy8CSLyP/aBLGFcVS0UQXf+UEMWmrQ2VuJ9WuSQ8gU
cW5uKex5c3XpYQIgqDgFKH2eoUOHIpHJuJvFIyEh76BluWsaLoo9L70cSgAIkyWS1QZyLgHZsXQh
7qQoQNPbyeAXQ1k0BZyZWS2CpSvlgbQmuAdeewwVq+Y/Yrh2v01lNDtmaed92+GDoA2CIs8sW/yS
f/uqpjJxhwNRsUKIJgYVAC/XrKBqcObgEbRB7WFqKM9xP9JcnXZHyHDNvCeDs+7YKFca6DRjtaMW
I3rT1gokWV/5R4DQXAyoSmtTdddNjZfSbxjSjppFGNPKLAsMN4Q3ymuiRjDHh4HdOL6UTK9zthtc
nDILtF/xtTK7fgQY7ZUjzqG4aJJmYX2ZYFFMUQtZS9N7mHdnvx0zDfyzc2JPdpidJEn6+7Gx7unb
0dtdK2LajwP/8W3PWcseFEdSBgBGTcD9uTsxevtoYX00gzcPJl+xupsMoRv+3tZa6KRtNS+A7Fnc
QFzeYU6rFU9eVwFN/qiUWa/+I03GsO9AdqfqFABOHB8XS2Dj1cbMsg0mvLzr7Cnzz25IiOBgsLFJ
xEWSbNcXfPMjV0/2or9AjZwe5GWver8MBnoJRGIK2jNW6LOd08efeBGOYEwTa32wG2WQYvs8dPSh
tUA25ZjVwNbaPSyCRtTmARST5jOMyxpyi+dVPkC2TKTkS4PkgMsIbA9NNKixVEl5V845ZxPTvKwZ
s/dIOsk/DHNNhSRUnQ4g3sk9w3lb31Q/4nxGoTczA/MjmB0gqw/TKdvwEpSWRj0vJGp7gsAcR7GR
dmOfiX608zA0P9x/xx2IIDG8GlFsktueaWAtO0lzUUCzw88tZQTWgXllWf3udcruAn8BoZS3wPZp
XNgjaGOLYKMfBV+tnFxyU6mdWdnP4i6DpL12ues5/abNS61YaCFfIxuEYhE536GH6a7Xuur6TKir
hIqBWShZ4clWkOle6qUzrysB7poYWMhKkCdh3h+us0PWxUTQ34jm94erIsArszl5fLm7rsIjyLQU
WnBDCM6anxSdeHnuzMTpimAeeze2uhCfuCskAiU+r12Rwef1ugl2EbFCg/HsVseEtMGRnRu2+e0k
i5Ncl/QaJv0bPzbzFjIEsVkdyOdDjyM3KhJEcrKQOvlwMTYsKjEooaF2/SOaSL9LasPegsDWC8sd
05cwgtKXNFlJvUEE6Kod10tDiW8/ubumhTCDzVosZTQERB8Lvhh5ETkdc5p4aqzKPeO3LJ2yWyle
dorE+7Dn8iliXTYtRMNZNzkBewq/4aNV5yksUpjP1pINNgEvA3EJqD81gBCcfTcY5+vs6lIacnze
+sP/emjDxzdxmPqc9Cq3wtoHLW9tDXcrouAr1HOvrZ+oQSfdJEOKCnVMmICyu1MrTOuGaTPLhCfy
FXQMbNeQSUQ3PWupvkVdv97q0RtBg8AJ1/gzTf9wz4Nac4Y/rE2dEimS7v+PlhQoKpJoKooadrnl
2Izr0LJ2vmCG6/pTPRqb3yVWoly3Ha5og73+RkngGPHeXyKPNmgbdBcZa7/kr9ArFfOSRbaBMp2v
BHx+oXTXzkpwR7G/W6YZrP2J2QkyMfgFT9pmFdhXDqWq0tFzIU/bVoc3VutRePKziZ5I7DrmNqLl
1zDOtwmhwH/HEPXnxD6M7wiL1UWcBZK5blLl4m96OsXM+PTH7mhe5AEmaBAB+GG5YGyuxcCgVeP1
Dp0/X27xdT6ysbZbYA+lbdbZUxns8cX5G4gsI6b4nYx19gQJEaWlEsUEEne5b6rNSKuWwHtNY/SI
vU8Y9GvFzkcAVUE7fFk0kHQIhl9UltdCzEBgMOGRoxeYwREl4t8PDub3hcnduUCbV0kiQblRF6r4
6hW1dlm4/y2lXBy1+LpqehIk85Bkpbi+aEyEhjzahXIDlNQWOg8/ugxYiva99h1WDULPDQ5skYIp
EDefnOL7NjllHS4uzRbJxTfsrdBaGDkCF4fKAu+rNopOEZOOgDWnqZjnTsk9vRQuPXkokG4S/CvB
8hWkSMJ/dYo3ZctZi++HcmfzDyFJnB7I8jBtdijb68Z/3jvlx+3v6UyJOkC8T10clYeyLuULn3vL
aCy/euhloumw/LIzf1/+2gsIu0+vlvBclIqeM8d2RYnntQevbiDL31QAvhGnKqC38XN4Av6OiSa/
G+snby9+ugliWXEB5H8/HgwowpIbk/JLp2mbLDJvSGUtxl+qRRRgRV4mBw42iIfTgcqCbMfENxyP
intuAnC2dkSNW8NjJ52wMVtpbVEDwE0jI77k6IZ5cy7k1yOI73LJ14OCLqrwvajls4tSXI4m+55E
FTe5RrCqTugL+sQow3IQ9t+TJkW7K5fTRVCmX6hVPNqeyHPCOayrlKVKHGGl7UYCn+NS0o2abuU5
WqOQbLBvW1syZDii3ekU/jHTHvBAWisVgkX27fzmk39yEPIZ8MNkMF+PoW6bxBHHYgUOqW3KE4uO
uJfii63iqMHNuP1RuEYHhUYsKj6JxfaQ0xFdB677n6+v5YQ87+dq7ecdRma4eaTozjFAqbt9ykKP
vTAey18ytQt+6IbkqV+5QtCrTr84CRgoe/GcwwtO4iuObM2BXX3T6WaR7YbKxercMGUwn0Fj9v/B
o0wirmNwuojIPE0d7/MM2hmzM9H2OK9y4gfJS8wJxv94yVOpTQiNY56g+wsNF5uizk79r0svxBPA
aU0Dn9eKS8CNVPBRS6s4WN5EdlzNSGIuj934fvtym9QHMpgJ72ksQDnNacXB87QxSMlJrHutOonY
b2aYzpolMQZ4kky7xDc9KtbK65U41sxnhCv6+XpNmZKxbrWctcbwE2kmsgWBQJ3F+KXqQT+D7uBz
AahC2n8qixM/3CveAKp93u19s8TNxcZnW2rex1FOkkRm1L2J6085FoRXcxIbXG/9JyhIa/k5wluf
030YImTldCI3nKcdS4aBQrl6lN91LulGwSG4R8Fc4PhTsrp8ZR4ZRX5fgiOcWorJyQnPFLpIYnCo
LBAkTzl/PoaTqUix4KSvXzDLuWz2dsxPK7yH4apxTf8ez68W3UOjnkGg0zenEss67fTjrttH5js9
fKEa2WMPZFaXeU3PP/zIk50HEw5MNnW5KvA7IUJrPcWo+s1ELUufZ6cqiuylrEv5nc5q671DgNOT
imi1MR3cUOudBsxoZjWE2Lr3VmZSW5N1HafrT0NUfr9jeH1bnM5qRaD+9yrJBybWZWtBtSwoOLIf
eeL3B0LUSYZXaFB3fS9Auhv41WvOuSYnQjnaMgcvUdqKVvJsH2alaOJYSXyz6YulZ+1iSa77Huso
G+tzasMe+wAG/JMfYRHbdihPMWyv9VWagToQf3EeaAUy6MfQh7uW6DweCibGTuPW51/kxFSbddlb
bjd8f+9fdgq/IcUgDEy8Vp/8ELg44BMzGb+QXIytJ50ITLRoN58WLxZtjySvI7KelvB3oP8cuaTq
HI8H+4wxBb2kWBN0QAuDUjZ6bwQJfPY+vxwVNNCHvTdnAEoYYgJMuMzWe+O4mTYJgnMljOUsItgN
uznUqgOX09bSG9d8xW7ifwRtw+/pvbZGxygHlDFYZxQNragNMeEI61muJSQ9ZOutAbeOR6plwrIg
5c4Y/c+E7+dZ1D6/qQNOMs/h0XKr5FZXbKSNPGwKQIUGDRJLZRTWEvvmg2gDjwqfSjjUTDWt3jNR
e4t8JYIMwGXw/y1C38HfpExXYehXsLBPAWz0X3LoDuo8dAl2iqZzzLfXSXFdJabju+prTKUOrjW7
RFh2YWlOR+LvJRu6oW6AV5Ks0T5U+XyUYmWbtjj7YCbNzr+DAqFDTA8sA20SpAB4qjYpkUVMQLqh
2k39eRLy4VxYkvqxrN+JYCZglG13LQtIsHXuuMm30qV8V1xg5BP9YlMJTprVFQiIYtG9/+Uz+i1Q
cE/INxCTQZJ52itWkj3xEjjl1lipoqSyBczCaPNAEWkYFpWc3Bcj3WFQo2suZ6CT+YobEG6Qyfv4
UonQEOrrT1RYeOecvlB1GTI9nKzDffeXTDnoisdzwt62G/KgginAjxcNflFFNHBwn4umKrnQAwD4
Tw5YEJj29sI8wSS2DE7KIaNY3BtZt1mvy82oxyr7CZ0s1V+xOuijrMgYQiEggXOQH81tEl67H52Z
hrk9+E/y0tJpF6D0xnw3Xf4ErLsjAHSHg5tt7q6D+6pr42k2d2EMZ3Z4jH/G3GAfgZ2mGah73Rsq
kEvm7YrJxqPYm46rKd2qADVLoCvSaRKrQA1yz482BepLc8RiVjAKFft0DV58H7LlKskFlEf9cOcq
x6lRqhnPl1T+y/wD5eUi6GUam5pKu/6HkTFAcFHuJpUE7+gXpr2K4mXI9Fk6n6mn4HtVa53pOsVy
BmL1zQ4oYv5W7QM5BGtpajqeKjzByzR0tzFcsuv8XRPTPq1LeCYIAIwFKnakvLVbh1XFfsPlssEq
kVQNwEyfvSDs4zHHQJywyIk9nCYE0I0/VouF15zrJ8e87pNpLoKpqCF8n2dKJKl7tee1bxrAfMmN
BOUCMgZkm5yjJy5e/qtt79WEv3Vfk7/EpvEbJnf1cdeAWnKpjaJmxYj1ov2sdBUUf9rbWsBXsxNB
aHsHYOCJ61uQ3H/KwJ9/47GYRVa6QPHw9ol7Q3dHNCSHqbl1OJeeIpe56KBz0JM/iGQfcBjRO6G9
Gp8x6YOF4i+zQsJY3cloP8uVkYUIIgah18BAXwRsPHVYVvRMtm3qIYFKZkxbBuAzsyqKDLimehYk
AYoDVVnYWESQ+6eYqMPfB3HrgW38Flec2SqnTZ7cy0Vgr/fFU6xjqLCfEa2U3LbEW5znHWpdpZcD
foKnJ5EXhMbjMdxQWwIM3zodYoLhkq/lHr/6Z2ehKP0sCkga00BZYrdIjoRHjetm6/gxaSV8QmLi
TIor08yAKJpzf29f60AtRRJMIRTA1wU1C2L1JSqsafanLd3p5mpUOCmL0uytktj6NKn+D4DHJaPE
yjtAGWHHr0CNaCOTlqtF7PBjO6aLBcShMewuRLAVH+/JZ9EEi4x84q5hQc9RNdwhZNtzUu5/OR7O
5JMxZwUIVBET3+V7r46R42y60lUs9IUBtxbUpsQ33DZly0CC6GyVbNTwuXvOd9vC2AuHzGCTIvek
f+dqrH41RKecd1RSl2B9yCa7R5fDWrr8c94bkSsyEgE6A2YyUtoYtmPj7ltWI2S9qNcUofhvholc
rrvgbMdYo8suHX8vkbfDqLSexy6fn6NZnpo4zUXtkq8C2tQf6wzRhvk1bKRyPO60aFIWNwzAnhSF
bVWjiKotNv/pq+QNSw3Wq5Ix9KNcVd7tVBqF3CeOggX9WVrAplxk/OXUqG2yoE2IUnMpHP/nnooP
EiOPFbFTG0WH88redt7hJxuLxLLlbbQZwd2sP6bHnNpL0TBAfxwwcEO8UZmb+/MsKK/WOcrxfhdn
QTEVtUWZdpJ43KDfCvdFSeI0dtCo9a8pZDSepZrTtXbvlrmyJAIxVjMF56f9Q65IkIAzou02nPe+
3fb+PdswMlYPJ8S3c7R8WqghPP1+HEP/8965ZIJBRN7MBhnf2jJsRS6LvDSsNBrkekN0ty+v79Oq
5rLbUSgE5uH2H67hqiOZxpjnkO9sPRGDTbrZ8g4th68aMa6n8LtluT2kdMdlxabHt0b1MzzTGCQY
nITUEbjTUZrwQS0S2ncXM1KWmBuMJgM+DyLll7cvdryGXkJdxGb6idFQeeZntJN2omWFKrGKF4Uv
XqV56PzBiGUnD6aUftBUHlN9RrHVC8htHU7NfzqMpG3d48cxv6wYlrbcUoa/ot+7HmnflQZO5x+S
g6UXjf98/IJ7OFA7pa4ARi/aoSGyXLXCLyjCzpV9Ywd08Sh0Fr4AxJggrY2jOVM3x1zwHtXTKFBe
EIS2lw4MDH4CRJxWlo1MgD9qK2MfXzfCUeELHrbvP+J6/00LWSBbMr4u12fitA3qvSVWO4aNy6To
hgSgKSnN2FqKwnGSQ2RKMNmguUL6bVmQH4HSolkXgCVqn5k6tNGn48qgUp13hNv8m+mcvrX7bSoF
BuFCo5dKiF+KpHzH+GE+y4oDY8vBabGNXTD3K96PofLzac62IHvGeQ+Zh1FIEvKE54s2nCQ1fTyN
kOMGXVfoNavQc/gB82A4pFzsq8+KIzpMxkWpXO30z7Qwwmcr+vT2F/nRgwUYVAZvENlNfWLD2CUF
ncHPOhFBnt8Sgc31j/Fk2zfmQ5/VDuEYeppwoDp8jyCkCUkp009mkm8Wq6Y8vyVdM9NEq90xkdhX
eLL19iKpuseNX4VPPvGQzz4Lw1CZYmJhHIxt2Y4NmzYzBQ+JhbGZh/reI9tjgOKAaUzz6xZ3MUkO
PXrmhqiuprS7athRIbemmMbZjlHFRn1smJVDCt51yQt5VyMr5PTAimytzMkFtGUR0ksmvWPPhlJ0
X1Jxk3EVRCfU00iUpZNESkkqnrDWhrbWWmjQcpfiTcxq8BaJSgJIyl/nMLd2Juzseir3nvzZEy/N
G6klL2OEeLbbvWzO8Ab8DGAay3JpEnZbmtaX/6lbwTiwMdlNBGpsy5kaplzVpeIel0q0RDvLBSvO
1FkFaABO3RmWY/HUq9O0ROzwMBJbFOp656L89kxu7toEWomZ9onQAm4HbEbNBhytLRPeU1Ersotw
pzbZOSGrxvaFLswlHOtGoZIcaRbrcvHnqIYtH9uLe8w1liIa8TMkFNtMk7O4YtN3Lu5cmhja3Jzo
gZfU+YuvimpvVSvQa/xr5iPgT+cwT2tzmnZzbXgF+QNEJS7VO/dGo4rfoXoFvqyURiktNP+TrWD2
KSXLEGJGwZrG20Iw9pg+nQggBLx+NwpH+2kQEYoLvoPzN2/gGjqVcehMgCm8IIvtFwWx9Xi73dWC
O+dz7QVRlcA6ClVU7BjEsGeWsTvvWol1onWRT0pZ+BqncjdkGCgZdC9oiSFDhmbf2C+CjEwVMz+J
UY9nWTjimB8aW8b5YI4cjVMx01h08zSLIAogCrsf5KWzz0OrMrhtHuA7UvZWJ3mLkyU+0h1fGW2A
4p6bmRGn6ik5X41Qor0ba/W04kYm9/0JXGXpgN/ETHUkMynkFmPlOSIBZk3rGvXCEEEkaZpzuWjW
bqrMgcXjrBNYzbN6x9FrKM35B6OT1BwdEPMRHoeqUOHDBzutija9retJSKPG3inXlpWctlr0Tlj2
460850mYWWLpSvFjnnwqB1a90IIhkUlmCPXj6wV3brzp7ukRvt4NlxCv7XEqpNYD9xRPT/a473H+
6uGJ3GtPoxlb6ySBDm0XEZc6XoO4Ciwu2XITQTC1aTmRHhEwnm85mw9IcVBnyHYBDNiXZy+Opvhj
bt1Jhn4qdg57R/ndRVQnzX0H3tgpvT5aIKPP4+mF2EHanz9iqNIcsEFRd/dmNuriZc5xXwyeU/vc
j1L+DTovqea475v6XQlW4xPvidSu1GuGDO5Dw9msJZf2L/TScY2rPZd4fJgAoNkXvh4u0MMB7E96
++v6Q/ywVK3BkRYAxuEM0kepI1Fb6+uT90ape1SJaAT0uroB0w5nXUJT65UAZILFOaF79yRiZPOd
up9Mt392X4o8rt3bL0S8Z8NLyzMYuJnLlWPzfXiWV0AdKDs3kHUh+vwxsGMiz/io249+Z9dsAJAC
kn6bpAu1ex7pPs/su9lkGh5FJFMoGUnNTPgxWy4Z73SlGE0tKlF07nAL7V+UHAo2SbWOOGRVE+CP
f9bsLUfXxDaM7kRN9KdhOpSTTnJoWhiXPb5zZp4E3D5vFKZNleJAwiK4QMBKIAwnmgL8CLDUm3qK
pq33KRG0lO/64g6mYoOgoW2Aiw4KXGbmqjyfxtvarFqjxF2JWaQ35L4fpjzpOtr6MuJAhH8lxhsL
I0dFJPXotR9cunx1hztpC0rhdTTYNCqp47WpdKvmu8RGXk3P7wIsWOaziaV/ee3P/IhvMAyLD9y6
Dle1/K60l9AG7v7X1m3iRqCEw3lBhy0okDdWVqvFd+Vo0TH8kVacg+mYRFgLdB03wzeii6zpPGaU
r1ACWOEY2tG2RjWjdR9tvkRPW8bXGdYU0uWO2P0gQ91WaOuIc/LAHu61fAnL2yDQhVHbEV1s/AeM
tU5+Q8rEwbVxaB4LblPJa4L19LpAiADSZwPgTl7xUZIkBF1AIh0T4H26x5JSCxgcRJqPPiq7JZw9
JpUfhd53lnHelaQiSsvngb9NS/JGrT5R365QjjjKDjLNZKk83LURQ8GCKmMrCjv02jheAduj0akr
1uQlg32ldnOqhIPOf/+lm93tJSHHoO6bPcgWGSCMV7SeR0ylWbn1XHrPX0Ei5AZyrCd8qmfdtrIG
CcuhFKhg5AVAp/d47mjtAyheCW0ISIdtH41LYNslSRu1SJVYBpDATnBfqPIZ++qDL2Ke4Hng2Hmm
e8kS5PBMjKnJ7E+nrUyYpW7bbF8VBZixWPxPHDzae3OGyiJHAO6bocokHzkw9U33UdTWu/SuW5Ko
0scIyqXK1NCNCjiVnPhzhSf0xlb7UsbEiIWbIntxUEo8uDPYd69rpSC3rP8xJil4V8wRscBDEbQl
4uK5qF+VjrBj5+PgaRoTZcLbIjlKtm31+1dVJyUoWEtwac0DGGeQT3oFEw55LmQm4+ZHPAcu/YxU
7uIyI/gtLfdR9h2InDyI+u1RUXk985/Xt3xgokT0yokPgXc55Ni+ZVrWczbT87Bsn1TYVx009tmf
bSjLX1pZ8DcBV8F1wiTGubtTfWkvoA01WWt0x0SYmkmdYYyrLleo/Yh591nkGddOMrhalopD4VcZ
Yr4RVO9P5Kg5CfOgYMFRZ2W66EruMDdpvrpeirCInFGdTHabMHNwmcOWg1dB0mT8LTXJ/NR7x2hB
A5Zj7mHr1DvV0BBySQYE1yHhetfxwFzPvdsHoRonpu3Xyw3COCGxFCCkdBcDXc+nQLJTap1Ev0yF
s+vV5Vr7SdR7BpZeUM743GBEdXUHGoRTZ42PbK/XcGH5Y8i9xv1aBIXcQ/l497dsD5Xe0cZ59PW5
FmIZgn6MbVwAmyEWZDCiiyZuMuhdndqsp9/CSSH43MCs2PN9a3DdTfKmBB3j0UNpN82ib9iWSvJS
7R7Zt1V7hTqol+HxMQP3608xh/IZvwrwTbbyaM0nEzi73dfuX0Ez/pR1lX5s6nZVaLHUAdfcC1Ux
uA2RhN4t1AZoKVxO+KntKaBwAnvx/BEGY0vVduZO4NlbFtgw5jC15HqLDO+mJqXTthaKSgAsqql+
oLYMi1rInJtceza8eGCtISnNFOHII8AwI6JtaK+8Djl5PILcEN7ItCXXIAZOx3tiFVcQCmg8bWDI
JiBE9HW7nvbhVuC5c4JJNV/CaX8iGN7VGW/uMGSiVHjoxAxFjV9JHpSbFBTsJlhqlyZjawbq7B+n
SJk9NINWoqfKmltgOcV7soUYQTsd9eAvivez7VR8DjwQ7cfHrGInL08/1+oupdIfs+C1EoQFJSEP
6Ttvc7SVIXCmTj5GLUSo0lHRJE+J9UOtMXo1pYDS8P+k3iLUznKlF/lf5s0CiYV1O2Q55Cu/oUK6
Lxfu3GU6TwNQ+EUOeIGyv2iDflQW8Da+Um/GVkGAUVf4MvoCjha89XL4VkJA5DAQDtVYRGYQ2vYZ
zYnX8Vv9TauqIf6VqrOAru09lUJnzaD7qlr+eEmF70+mJjn4s7cHSBSGmZp2Ihgq6fhuFmteuZcj
zSUTCUn87zEv9/QBRUkuO2mE0D4x4w6dJ5OBXEM2jxZPowiu3hAUxomzJ0kHgvvQK0cMQjrPaEaQ
at5U4NUcRIG60GMvg1WSSBwU+4CJl3GyuvEhyD/qYhlLXsDkkyJA3xqUME7Bs15uyodKbLSfUyUS
wuJCTumxk0Z/+pAq4EG9mSFa58d2rDOcJsNoQc3X7IP3KrczVllCMUzweH7qpaIZBuWZfhanQcxL
wv+0gkkWDWnud5qycpOSSRtwc5f+2eCkrMkN/3ANhlingev+y+PoiTdfszpVZzo0H3zhPrV4cwQp
fIGVuteShaD+m0AJkUS4oj/kSB0f7MJegCoECti+ZA6LjZyFoEKy6JWSED7/nWLM5drlxXwMkU4T
Ob1K1Wqok6dhaXsvY0EKZOvKRuATF7jnXjDPOZ3ilGf1dhWliphYLFzY5sw5BphxUbPqXTl2dcZB
6bUh+n28UDiWOMQ6YgyUGbGJzoMQXCYRyHeThUJMjCv0uy/amrS0pYS0xdVKjQxOqCb8Q55P/laT
WUybuBUE3j5ry91QXD4OHnyN8qO6tY7Ulp/DSbB8eYkJE4CaPHujVxs+WmCVzzeWtjccVq8Qk8hb
YlBojjcB5NwM7yaj8xkE1HirytCyfb6/BEZ2GfnVsxSvvja2ymKFXI1Fe10xWB7xsjuDWmtv1w10
VUkKFYqst+NWykk9kG25N+wPSgv/i+OscJiqDcTKdXV3XNtvoZHc37Ej8Ya0ZraRa+ZFPqVA/8qU
HadDX1O3XTDxjn3sSY4DLnskr6iuZdUU6dPSWjRsyJjfUIiGrhrN993ksyVqD5pBw3c91bJ3Dsfy
ZbSnI64VE7BQ0bI76zm3+umt3U28oNyVyziTtCTF2Mtf5xYbOi4Iwfnfw0ldKzSTgw62kl+zUKdl
CSisYmk6zYx19EcQDlS3Q8SGoO0WAd2kDYpHi3OIJtnCLTNhcLK34eTkzHPtKaV2ApK1oAD5SMFj
RcwOzfc4S82xcuroh6WtpLWs3ybzuAh7VqPTLcWe0lh1RnIjObrZs91KIPuAeWwejUjlFZFZxM20
WcLm2eWcfgP1uM9Px3Ho1jxH7QZicAwQC4j77miqUGnJDP2i16JXSMsMzG4uo0HAlYPRjZQXOvGq
IhDqVQGgRB6O9ac48qM/n2jgvjKkDqbNnsM6Zcw4o/YQcLMEiPUUKcp3m50WJnlLsfoA78SVI4UA
BHBsiG1Uw8pM4P95+tGY1lFRFzMKWd0I3w8ivq77FF3Cf8pLW3EYPOAVFO6k+O3H5iEfd/XmrCBT
waq2sAC97ngdPS4gyQ5SDgnAbItr0kspNfBXdK+6Vr8LH9L8pUOzk20lNkhHZj9w8nIlCe9DE20a
7pnJaz/OlW0+Adu5tRK3Xymd4QutQGMeIj3Dr3iQtfstStuFqfBjw/7YCkWlS9bFD1mzw1p8jqo5
J0YNus1thHDZy/LA9KhMANcVLm2xzC5zKSCLm2r9PkP17HIqVjp5+QWsdrG/fXKCV3PKqSaoj0RX
VBk1W/YN+jLhzzyGGyoyF0M7ZyKiH+L6TK9wq/qyfP6/wpgdNwWzQWhGBtF9EXsrtitm8RjiSEiG
I1KVoYte54jNc+p/vFOMi5v6kz44pxC4s+XqJMPvTtMr4oAIdMFnfxcPfWQqNpBd2GpDIV9mWMrR
Zl4eZthlXOcfqbyIBQ54Ht5AVpt3FPlllJU8DJ5+k4edciKEXcIyOJS6NVycwFLDOcAnTOB50dXP
zp0jI/4O20drkEnDOd+EjBIUFHrn6BcH7b8znFidHT4SlJB0511/E19yCYPfcJJrD9QmBgIF/SDP
HL1jQix/d3aHWADzalzrlDYgrJdq1z2C6MdcAWMU+6WPrg5lLdpQD59eGeiq9hRRu0waLiowpitG
1qmvlk97XvDUCALDXuFlYDKPVdRotH36b+6z4KSW6uoZ+i6ib4K1piGTeeld5Pji+6OuYHzIHFuQ
YCspaoVH+cOr3CMSDziDIJO6+7ZIkie3fhHVjeQmskXtkgAFsSj2kPM815LX5fVRTIkyDIvPQrs/
UYHd/9dnSBhWVf/cWrKL1DzveIvAITNTctC262SGi8gPRy00YhMGlK/IW2a3A10DaHfPAaHTm0I7
TpeCbmL1+WvkZ/H9wQ07RKHeMqkyUnXjm1lroZN0PTV+BnZNkOvO5wnC4pDhn6YgQjPeNS5ALzDB
cf3zE+Di5JGfTJ5evmSTnLsdKLVTXvae0gMIHwd4FYDYFYy7QosyFuDEC7xa/LV/tx77oJP/2enM
YVRBzcXPvyQISFIQad0uWwYSROYtnXO8gedT3Cb71HVXiaMVKN9HkIjYFNRfXbRtOZ6pl5d103NZ
MTlX6P59AvMozu9dwNOpbpIX6kbpc5fAkjKoojtV/1WV2iQ+A1X6+bpNyNyR7EKbhxvV6+/nrwty
fYRR0PnZePfB/42+IOXOux1al+g5jadKH7OOwor1U82/jQaeYzr8yBdfvoKUC+sBA8KrDb2WAT/G
O0jXPVAI1jukq2kT8N+Au7uzNYhdfLqggKnMMR289b3HWCU/bbUAxEAP7uA5FwvP3KjVy9s77sdu
BK7Tf1gXKwdTC0cmuzAnpYFETPNwnTjMiaZhBybsKmPW53It2wBi46aHQ5fTjyscfiGt4PIjVF8w
zO1pgQQDHh7SV+ERoeQ8LnV9/LvM5R9XjThiWF9WkdLfs+EW9JkT7VnikAGE61AJrTL6LdZ/hw07
rOtbMpYt/qDLpvcKt5+QQe5LqvmBU5zrYxzLMERS0woQJ+wrk9QPuce6uDkhQoVgX6wlKgHI66mV
CDMwyj+lIfkK22tUEIWQIUk65MlnKkH3RC4e9fh6AYP0Znnmtwab5H1y7aWIERSx4kg0dQzEDUav
ILunfqsaNMuxVmH0vpul8Slxdkfnn62JIm1NXsyOhDXkY7R0Xhqf7F29tr3GXP3H+cMKj5mpNWxA
CdKXXW2hM+Ms0ZG/XktPG1mnnveWPLa6kw13jDAo3wNfXjtsz7lzsRaKJraPLKquDu4oqZ2yqZLL
5aK7ZD1/oXB8nR9y+1Zl9xX8diefUZM7o3xhecyIavZOMycpV0GKtj4JHQ3UgxYT+iNcGuxwGtiN
5oZUtrJiZca+aXlj4ruSnFg5PSra//uZkRtA7PDxLUegXOHYW8nXSBR2xzFCPyVyDNAZkIHErbTf
UUn6JmM0dgHu8lCfxtJR5jvWYXEwKxcj/4pAMQ5mNQr1peqBTdtoS90RduyyVeCR3IT4SIlPrllL
XBaUTQdSrbNf9seCRWbOl7mkJDfleQlmzPrOvF8w3U4zay+2fOLacSzgOZu7XGRbcAFdUE5b1toP
Q0WE7flYlf/6HaiqqG/KHFlQUcLXnWAyPXsaAu8jDklujoL/LFEAzyPYr2cCqe8NDg86uyQNd2Ng
emtAGYxlikONWVHclWMSm98bLeiLW2dpIhyrXHfGamVmnvNHSGJtHNkfmaztEggRn/okxnNFJv6p
WhyF0mVJbRXd2PQGsPkzloNiszRwR/lRQ6Rkro/kUnl1pnv504ureUU5rxLaLfTaCU5nsNa3e/W6
8N+n+ey5XPOy6apYLf3SpZPDOKkn9TAHf/TEV7B/6Aii8WCvJtiwk94mh9alxdmJl2upRwXg4yQ8
JU+qvueSGGvTHwBB4nomZadjTCZPBS7/Rhtt2VRu/pd5wDhATJsfCZIrnsIjyKoMPT71AVwG50bY
VJ7h6NPRK/gBGQ85WaKU4KUXgEqHaah7UdJdC4Aa57B5nxCuu+uMkTi31gZ7ZI8QCSYOKGgMcYkW
JIvtM8rnz4nRvn2iI2I3eWFc2z1NkXCBNXH4OabVGOsdn1eDT4RGwCamPUJ52DIk2Jcw6Nw6OQbH
KnKBEP3G089rV6Wp8TRvWS3N/bYtxm2SZhjqURh6XhYamMzBmLHlzWdY4gb33tgJ6Q7dyy4rOqPu
E1MFdej/Tk8wNe4BYDVtMEjTCua0B63ubABaYYBi4ycjLuBbbLoY+z70ExRWMajv4Sf7kR6i9LHd
Av4VjcxrF3U+DnSvzKUzUmLIsYKkOLcLwekq2U6eaRp4ZE0ThGl9cmlOQ8AEhXPZu/T31LOZjHGl
tdledVsWVGz1oVUBfrJ3RNdJ8824+R4kl2aeaLgaWonLgWZsZ/RyvFuioz+RczWjNuyop6kc1HhV
iPPrUB33cRISQjVgRwKqGW8p3TGd9KB8jDwTV4t8wK8l+s4mmOhrppv8BioSLfoXGaJmIHOSXBgq
mmeG/FE6dVFj/rjqNuCgYwnxYtcSVSPNhfJPG1K4ChKIzGP8Kmme+xfaxjLuR+cNz42NAWfYOfVa
VWyNEb+OiLuvp1zIKhAHWVM2TTBQHQp9iLLF+HliTeHK2PMFuUiC8cG0Zuqnq5hxs7e2vVReLPRQ
moiVz1JamiLL/qvUSh2BhhazYgxo4z+bblyJat+BJZPsXX3AD07PHJBPdkdrlTkXLPmJijdEgDRq
7sVUkLio8snidlo13qQSRxR5oedaTKdQdmbQGWBT5+aFUtmYFyQqiFV9moY1eTiXwDXtznMkvQf7
hg+L6TC8vd8h9Lb9DQh4rjGKTLXI6AHxZnsTd+NIcFXUQvCrx5EH7wRPFsGSNK7gxViPKizO12O6
8rjvCGu42GAxZlyoQxvxMSNrvPWukQop38Iv0PE81tkscTyslrrfUWLR+jr++UXd5GkDZQ3x+ZRS
TfozTnOoritInDaOD3+X7SS20lTCAx/Ip2hnaBjSXxGvfvmZTOuJe5I8qbxjVa68cObwXK8eBNPm
JGr5AcqYqK0HpIR0eJi1TPaxfU2fPc5xvgjoDCNmodmTmYuIvmjs3pVqA6kdRN7wOkc5WIzfQ5Rl
SqJDf8dtXjG7Y7GY8Gqx4FB84lzfHKFadeUvpl8ZWSzTPRuPgn6xNjMuxtgpIQD/d+KhVFnFbNNt
jP2MdHx8sQjql3fwad8adIEvu1xZninLgNiVG7TWtFdMURuXK8sysL7jiAIT5QLQuoIGeL3IFlPX
ZQWjTWHMFwbCqGWAF3CzeOzGZFtLzbVHnlHhKfPqhS3w2GuClm6Xp6Pw3LQekM3/Q3AwbLLQ7T2c
jCg9yU2x5MnB01Wi8txdHcOkfwMmsNz0DqXe4fot1veo1OBCnYwimcpocxdyaqxhsYEsW7b40nnR
iAHhPd0KZ4fB3/SU/h7w2JJBtLVG0YACBUN++v3zEYWbqtUrJ6sjw70goL+LnUb9QrSlQq8qyh7b
WtEPXEkGtWO5QqrHiva0Rg6woGRXbqKvlP6RAZJm9RmLlkkIMpD5plJDxW4kOUSdtFnyzBE+uZQs
OeG6u1tfH+rj/EAY6cju9VzNkAhbeA6P1HR/RaXVMz8dwdxSMMcdxfCZlb1aTi+OhE3lrPnVoWur
WhJtHYDQQct7kzdSrdmwI8sHgTTHYS7ZsvkPv1VyLqLx/ALX8zbdwnViar6i6inD/EDK4CcXxCQD
whv2XQzuvK4RJaQ5dLVTRhwD4jjNwefEks1cZAn24jmEIJ+NnCtT+1i/l/yolKijKVw8dIxn8vFl
ZXthIuRr/9kYUseX0w0E8JXtS46lFAMIIpuRZSFjNR8cLTP5a+lVf90Pi5tTOrkFJ7iQmueWHs+E
xQTKQd6Y7+YIheJe3nzs59//anWX7JRyPyZYtafjQnYVBiOvgHz27vHbzAWyq6ukcIH4v2PpUrYe
gDtKhESGioNJhnSooVhixWrhfSd3GpOf9VzvLsYWluoihePWRCOm4cT74kGck+E+B/DvGLQ6316N
KoFeKUku4/pPJ3SU5Pp7Hlk0f7kbzW/wIPPiGk0N8S2buPB0dDmY7fvtQRBjWTQSUh3rkd7HJla3
7HCbGeO6OEcvSjXjsedWnPQPuCA+dalJxnmPXenSz1DQJFwzc++y0Lf/CBBu98G5OG7AmVawmg3Z
Gswzbg/oNIWSI4K85S3oY3noEMEZ+UWyPYx1v9SJ5coTw8GgiWs763gEcvmDRK6em0G4/K+pUHo5
BvIiF4qYmCC5d+uDi4hwn7iaUb4fI+2rAXpiyFzJ4dUpM3DKV9PewR+4rVC5Z/kX9PnDTmaVBNqS
WuIU36xVFpDHuzAjhzYhGppTqqRe0VDn0bNxIXSnpGqKVI5C1iIm4U+gk8aOVGIJp3oVU2keH+y4
7gETbdPkbucE/r9lgb2dIeFGLO1QGABjcKJRoun6Gs5QNrL2QDO8HkEMGLnywFnIQNRLOFHaFxIC
NlKobuQ419AL68mZcn3nZ4KTxqFfhU/1Zve99W7zO/SrM7zE3U4vG5z+Ukq0xZRO1XbthiVpqId4
4vEeOZ3Z7EYof0g5+0eG1M9SacQKHa49WcFht3vkAWpnX5D6QFzS29nCCnyJWiKCFRh7N3zykJIA
9aFCFDTy+a1hsWLdaRzM0FwWqSg8n7TGzWwvgShoq9zTvZh2lxeIlKiJSsKZE5/gv+Ho6/5FAap9
8u9b3I3tXu+BInxMttPuUnSZVBl2KsX8dE1xXotd7IglDSH9FtUx6rIw5Dn1MDXa/OhnjVleUw49
9jxOWc5s6eoe15yB1Tdqn5tXbaCe0CYvedzAra8tjuyyIA/pXC86Oc/AdpDBIMnRIvBYhpqvjS91
8I9gzPJsgYUKpfFlM3xvnBvN86WoE6AVZ0uZusWgPYMXGH5yGLfvKgNErRDibMIo1DokXEIGxFTg
GUjENQIZvsfHMJxxO0dBtD8NTC3L+TxLaf7TPMEUw5/dgX5YWQxvwKGKQQLjoBHdiRLB8rfbvTbS
aSuGIl+i8UEhUDbEa9bfcur8zmuJSTkjZ8QR+8CHjHlwHHV6C8F1mwElREziGGz1Tdrdls7gPHck
SDEwCELe8uq0MrfkIOIPrAsujWtLjxf0lF4mMtWP82r/WtKCGdZB3C16RJaTiE79KyhICZZW1FZa
jlLmYvunwO5dtZzrcpJ3qpWz8Y1oNyhr7X9LNnY95ncTkrCznlJCgE6zGy0K/P7jTvP7cDUh/Kb8
ZLtWpeZMtRZHKQvrG/4tPJ0vdc5N8Of7uJYVmYlllvXQN5grJofGswmNWHXOfTfTOdXXQCDaTInh
ByAr2aWfkzYhUQcLP3cuXIq+mfYXH53I+FzC2RL88Gu6iPggQIq1J+hm4aByxmvlDjK9Q8QvSRnP
EA2Vf3rEAOvLdJIto7roTW8DClukg4Z7bVUzKGEbH+riVN1TLN/9CM7NZmIk5sQUmzGa4nCM6WRR
uQLMemgs5Llpk53BADgVLHRiJMHtCy3TyyjOzIZYUxvNYLTzWqQlJFTr2u1eKdIWWgH9xu4P6p4H
2SsKis6E8MfvpV2jST7Z//atIc3xZzC6znTEnnfB+6HskVyH9M9YrQHJ1K/m6KN2aowoOyVdrffS
SgiY79Y4fhc2JLsmJ813mMPIRf08X0vOpoWbP8px/Zswxwzwvv5OAUBqYAOKNkmudV5BNDI/wSzC
KLup2HdMe/jgRQ86hE6TLKCDPgOXh6sAjOWE4X+0VRxxQfaajDh6EAT5ucLW1N/QUdxm9lHEHufc
rq5whiRhHi8yy6XXpORpJ0RyQB+xBG1KG3CqtJjeDXo8+NrfliY9zdP0FxCZiovC2iLroitzG7BS
ry7f3B90BSXdnGi9GjsCIKOuMPFd98kCbiCpBWMsUWr0eDVEyoIvFOouJCFMyEDmotVXzNb+g88q
7WowyQ4b7R0+Cf590+MewU0J0TbqzyuS20R8shCbTh79xQuaDIilfE1sq62epMg84ocNk/rxxvSh
1QX4S2hV09uxxCPS3d3ZHIwyNX8cg7ViLS/H1ehsEcJl9wmMdJBdB1Xyy6WTCAN98znvawmU7CpE
oP1H1ib8nDWKqj2wMPo77i+vtnX1WAsGcFXeyii4q8BlXUyfgfU+VIvd3ulPB4VGHcwFSU8XD9XL
57SsyIkVPNPwRt/dlEp6rxDoG/s4QdVeyLlJughV7EguDnfA1RDrj49w5U29TmTSCwKruZFATLQD
KRwK5A4ixQvWJvO1QhS1tri08QSwf2lDfVygtRK1NHe/yi35YFoBq4/XbXjWr1v+tsqzms7tavLO
Tg+VV4W9Nb06eViOa1pj9ij9mW5IMjwoBPzX+aOt3BE04k9Fftk1+D38u9d6PobJeDgm1Xli4MK4
3yUduCgFlUl5I8E4o6gtxanMYY3y5kLGtH2qgPA8vcvIJRWn5Fu2yjSN+ggMpLXF4qvp8ni9m4pz
OllKfc2VSjL9RBHPw+t23DJGSDf2GsXCNFd5Hdt0rFrnsW8CyaNtJTXeHyE75NsrNMwytBgR6iTR
8t45X/fHKUzNpS8exwuxR6IHEHI6hK1KrrRij9mkNbed23Yu6yw7xWYB+4rZMsbA/wLRE2q4DheH
NaF0kXshUomdajJSJV+K512wfg88h5KNL4FbnXof1svtUS6VTbXpQGT0xawnaOMB+ahWBkepkZvm
yNwstQKHOiF0KmzCL3jIyQMwuVDELYXlhkwXDqU4NvHJiF3HWCX3xwSI/1Po5kRDpg3I7D+Wag7c
5HhBjZIu2WrqCih1oCVweOwO1yC4Aj2/pnmD8Hpb2zxNs33sK2M5KpSgtbrP132+TUtYQb8/m6Fl
0PZ8Hb+mDE5YSKav2g5INspp6bKiLugzacP/Nte2RQF4YrQQxbeM26qcDlKMtWZxVVysoVi0ahNo
0Au8t+BBnfOidpj/ITWvVRUqfCv7Dydfa1T+ZvdM+bloTmVG8u2SsOg78kkq5zPilQPMU792r1pS
A1pTQkFf848SKBLDSunU4ObGJ50FIvRZX9g3QVT9/uUXqjXRQyTN+WzWRFY35XoZrM4MSbSkCiso
Z3ZC7TJCr6gD/131UX8gFgIby32r4xRWn2qgWzJboY9hRDFs1Qpu/BEi/752zeZMG1HC5JQp+1dr
j+erqlGRxO4r8fEPEbJ/TGbYum+h51zjldZhFXIXH3Kzc2pQ08EivCPkkwJ5IUn0i4iDiquSHjz6
UhcSPZtIn+ysk9G3Cf/NyqvWO+qXcOvzJjfrp8sQCW1IfKZIzAP+p7LItfpi25pw/Ko/t2L0U0KX
SzwcI5ApdTyYCJIn5UpgpkaJFRiifrsVsCwkRYS3M7OkWiQDB6kq2qsJkPAbcOVJQuSPsIPe4NWg
P5HStG+PqCgure6eg4sh3KhrLmor/VjaQ2zy/4IKyf+cRLgb5RO2BKzrICcfcTLFpbi9qVwmiQm+
nxx3PFteVE3v3GBURldpE9/6o3PYViITPNc1yw+jwwto1MUXKJwjVa6TMbwyn/Xr9NyGc3yndfUP
DANdDW4dKNhW3d0YVik54YKfcDjOejjeSQ+2nK/vzDaFC3TVg2RDP7W3sIL9A/wVE1WQU1nEsniS
WmFzymPvX6MtfiGaw7eEjxcBk/B417TOUWT3NmMwXdGNw8Rx4lyqqYkxYakAQa22Dg9HFD9fvowy
JZhgqitXkAn6QbeVILLuUPnlKUwAYus79VSmF0RTcFePREY/Dtk0m4Rg4PPKnoX7G6V5oeqbD37A
p8DDfJlHfRSFdlHtxh9TOBb8xNKTjI9mpqsWm3R1FRaUZRFmK19gs9CvjX0SIyCUZzNWsjW7hP+0
fYREypTRsUafZwoiwyxikc9JZ3H3DLW/+YK+fs4X2zwqorK0rDvFz7wGhI5Ukxnt7hEphKOczK5G
Iq5JYFYSqNlqV0Z60/sMWsFw0SxCX1hbImWRFnGuB7XOdkox+HNKOiX1Ff+dFu+3aKAzUuFXcAOh
b/cop81BvQm3AjsgaOJDgCOw4A7hGSAA6csJNVzamHdAb/eTrKhEPdjM6HO2qSA8LAkFmQM5LQp5
LY+eT/fGn+Wy1Y8eYSs340lbykkm4b9CsZfU2kqBBbtT74wXCst5N0zKLQr6d3ZQyTPCyKyatfva
lt3+2HOWS0kaG03IGUZbtxVMojIgw8NLGOsIsq/zBUWgSef6Ba7kMIXZPME93x3hlNSfzZEARlxx
W82/p72m1hONnIHcofGhgZLT/bWs2RCeC+hZRFNbmSd9WEo/YXLIe1YsmnNYAUr1NwEz/FEc2eSY
3/zNrDZbMPz1EFBP9mhlBA/gnulk9nwDXu6wp+ii0qfxMmfu5sWHUNfQ1UBn/N+pbTC8QvV3idAI
7WZ3LleEEoM9/A3nh4vVdhvNNdVeHTFozFC1rqNSyzljusEzQfu33EcU4ipNtRWq42J1EXcrbSOI
s071l7ef/eLCnCYnE1iaPbfvRTEBxVJVnZM0PrgrJV0RA1bW9yXFm024QMvfbgLUWWY9X0MLT/Em
NaflO81s1ErRFAjNuIEBf0pB5X1Dx0RQ8/fDILM6AtK6ijOTdYhh5rMatQUWZAeIIymfjQCC8f0w
rkgciPXj1jV8FzNBe89DL21g6vGX/vLFp8zI3aOXYN93NpCvcLi5gD4UYc3YQlUjrofIIlyfdNWW
ZFxxS9Outu4KXqKwpI/ZX+/RLbBGWplJrzsO9LicfMkoYXxD3iYpjNpXZMk016uE/5JPMrTBQWAU
8S7jrcwoD7ZY6qf+SJ//3IcIQ4US1AOOUt0Vrqb5qpQMuyNDkGbkdhG9gAfQM5muIFyFCYj975Rs
q1i/wbGZ/yrsR847gOkuotzu5pdnZ6lkfsVtxkfALxGkUWnpF/8DICCKD+sUq21ga1eWsUgyrDtU
mH1yXwvmF8TxiYGBu9fJWdShYFtxsCR9BdaNuEsFj/O4g+JB59zqEZ2kszRwKZghOgvxgWLbc036
pxYe8IrIXDoKhYvSEIkeVJMlk4NMBCU83xkI2s+voHZx8RBThyTPCBcBgr+Unss+MZReL96jna9R
2XrnnkNbE5Ea5BasZjKtxgv/SW0buzWC76CvnFxTU6qGJdu3SHm/hus6azRjAJKtl5jfbNp+NFcE
/Y25Nxzcrm93qJ7l6nebAMA9DF4nj/JS6LISqDNgOb2qnI+hXfzPrEAZHiN57HjlX6Z/oaY/N5SY
VUhJqlLMHNAZwWU2jM75Mc89kk/S6zkR9LYcRLf3gcbJXA+l6VxGZFKsn7DKvPlbSBmM4XDsd0EL
f3SmTna6gaXC6YERkYXN4Oty8FlvpMYeIXfgaMSQgBWBZNnNEXePzav+cKJTUn9qAA7c7Y9pz2+Y
Q8G32OzE2i+0uHD35bSnPmuePia0iiHSekQ1UMAco0/Er8aJvrRazVcpFAXxts1T5vae2taErcTs
3DlRVaseMN9RsHPpkdrIEjvGCj5/qXJgRsMcLeCfUWy5fBpy/WXJElIOng9uXbPIf7BvtI7JCGfQ
ZYRdgTM/Fgc1u3T8XGoHfpq6OGN84zS9LsQu2x1ZcE8DaZ2EiqzMrrOxKIVyJQMzklVq9axGOg7N
xcprZrxExJ/xakTJWvZ8bbGSqoZ5DLrKL6ju4oTz7BsGKaBrlXMFAPdHRLEncDf8tHCGIV/KHisP
ZInLC6J/pwyYgcjvBG9Q69BDyNF5d2CJu/tzmVkweLmbVPC+/VceB8jOcuRmieAa8XiYExLQ826T
OC9abzjVyIWUBT2QtLRCdpb7/CN2fHz32QS78jC0kar1Mhtd4SrkIa84MU7V90nv59J9HUhEZC/y
cqkgPPXlut7PdlHQ+a1xIg+DE1TSyxGOYnDSp2c9rkY/RNhgFmdPdtTfyvyVFfcSi1i4BtxfFr8m
y0txtld0e1fa4dtSw0Tr7fDpvQqAteUMWyvYGk869w+x76Xt/DBVdm12+gg84NFe7G6El+bRRJLu
txRd1s6IOs+hTtgy1bxSrz+bDG4E6eKCaZAdzUSK3jXJPd0EY2rmnZISjX4JgiqLMhfUkC97Pxju
q92D5x/NwdPTBFGc2QwncZNY1HbtdiFF2d3K3iB5K3M7/TaM3s1ao7AlEd8lXvPpiiqsq2i8XHrd
YOdUtxwivvVmrV0ATYgIlCwNo+s/FPEQdRR/hzUipJACUvDmbfmj5Hao4sxhI4IBjU243ALEQABG
k6hCvMQuRU0j/XELb8yK2NEEh8xtA6AWL8uLW70De3htmg/2Xr72VjsC9J5uNI/KG+fHhNSagq1N
tQlnQPZH7Tr9dW7Po23Himnxq17d/JSouFcaLO9UOBZXc7yXJ1IgUvM5hNzoH1UlZAUOyVP0Z1Jv
pluF4HhdOCVPWvxYgUnr+9KmKHdaIbdDQWcYsfUFkzWLsxjGeg+h7fzsqZTbSU/dYMxsWL8HDFIL
V/N0SOulHuE4sWDXk701Mrml5ju43iI2KhiafvmXq4XIXv7bydDmxMhJOTxvyy8uIIPcP9ax6LCQ
5HmIVA4LHXjxRyhKJ8wpRrOwGpOrRyo4NZhC1fmyiezcC95ne4wtf5iV/B6R7b3q6SMLRipuFmlS
xNi4WZQL+ItP472QspRwBI0YReh1QpmM6blBkJNb/jX+XfI9wrhSoUKv2xt+Ey6TNeNXvKSCGZoJ
XqEEMenaFZvEM88FEagVe10rFN17bvjqtXLN8VHGCoBCfKdqRks1AUf6wduS3AFhCl12iFx3GCR0
bzwdJYgSAzJY+VtEhLXaESX6fiSThK5jhBG0u9NtdcyRvhuqWOX6+Q6rF8zxpSa1qebbbrOE+0R2
G/MOpJjTYONKNYn25VvsV8Rc6vmV9Dg/Ghhh2bJVOXP1tWaU0NZjFhiorzvd8NfhohKS2BmKyg6w
6kJQ2hyBo804KPOQqqXkgT+y/ufj+mbTbQDNRG2AQd7Q3mpYTxOffWg+P+bR0F7RmyU7GBUeFHo2
4UeWRy+uO6OikKTligk2RAkxVBFB+m9HXMBv87/6BIsn9KeChE9ymddSbGAYuiqv3KVG0Lpp2u26
RLB2f6pvPoCZMmXqZb5zsEVTr+FkqRhGzr1Gj4Z00kcKGEhsyhCOJbpQ88XEJxmtDRGAi/oTxPV7
xtL2RRdVUgcoKB7GrxEutpoJE0xuJ28yvIOoYMkGQ6PJIt4Ghq5cJCmCjZuSGM2x5UASX5bZih+1
mT9xdXdJDh6dNRCD5CiEdoYhcPV7lDFoJH0b6B/uD7p+MfBDy26ZVqrVhR4r3aAXEmv4tt7HCNOk
jXsDLc+NjOQbdND3cmxm9c/fFG05KaJcu+w737ZCrW9O3cgoJ0UYzsrKpFzwfULaFGO2jb0g2PoN
3+9Io4+qbZNCYblpk/HRt94KjZsB/5DKEwFL74YxwKvUADBZFn925iIDZTqA8CJNha+pzGF4xCkv
DYBag/Np7m3axyszLqQOWQwM15Fn70M7VOdesp9sqPaejlXO/5dbQKgi7LCdx66GbbN2iWXxogRP
kNF8GJ3dSjJVKn8t+z1l5FyENuKdqAlMuqB3dEhT6vgI+Z+ViuhnDuOD21DxrAYXnXExoyN0fV23
/hkojn0jkqIZMmR6mie258Q06p0F/aYlGvB4IjYg7Hv67kYWQnaD/ozo0SYRgNy6BM/7v3Vpmqk7
L46A1HJ2vf+o7zx2CH44Goj8Cz+/JUXRyOosh0Q3JUXPBWhPgkqHacr6p5nR4z94bdTs0nSzJ7cK
WqKjhhfUOjAS7oGpE4LdkEFEBbCDo/EqmgUpEhhsDsp7YgHAyESTliVckHFqRtmYY0jdlEsGbAtW
PBRInGyX4v/6p+PLb2ZFqWim350XJ/b1VNJAMpmcnZFOSdPlM34Srx+SaQKdJfYaPJtECyo8KVhG
fPnuV/ai+Xm+mwsu5GLZcDU6KFZRowCtoBEIFS5nHGC/9grjZZ75eh2fskQuIoQCCE3ZHIqTSLkw
jlM+5GeK8chIVcsvbnTv2BlWwrpDa858K0UHJwWKFAS7bkwu9oZ9eyJbDGcXgHh20Y9SSR1fMa9P
/fLpQysGHop6ZIEKisf4S3MM1ZEOyU1a+Y/n6y7aHCHzMzz2eVJEIyZkKjfNbeKB/D98noJfcbYE
czit96P+hIjq7QRY+q4yyDACJRKq3IPolnxzQgt21tACXpHK68liupQW6oN5Gdi+HQl8ZA9NiVdd
8uCVHDVm6aFQGFKMyXBS3o7sX4klf5eUFvcj/DeOl89JXcBSmBzF9qCrzY5MHl0G9S2uyjRbSvGJ
9VZ3Azuz813khcfhJwmLVTuOG1rRlh5C1P3gpnR8t0l1jIOx/9PDG9wHLctfOf3v9UftBTyN8FQo
kwcPS/f5OzxGpYe/OtRL9eqhyq1S6psf2Nr3fWkcsojdWWC2MCKz2D5xOCIPoSa/G4Ko1IB88T5N
HQA0yLpias/wWisVdtpEsPtA7TVn9huvoPNpZfFKBaeXBGV4pn7xnGdGdaNQkxx7wbeTmMWJfD2u
CA/4A9WN/sfPVeGrWllBpZ2jxXd7YfuacVab+8eqE6tD25XRkS2bUQIfe5z2LhUbTsXbnR/G5H+O
7bSaEtWFcY3gCqlrx9iaERi5e19Ty5iXL+nN1rYu6ws6QljLguKsZkDEc3dziuHu9G8uyVNC5SK9
M5dK52+IY9WsSUPjMVzLV+51cpB+ChGsNCKcudg0dJK7cmcbxBlvAumTO8gnTKa05j5bWOUvjQ28
1qi8PuM+hS/Fz3LcOZj7ktfwY/+4wx1376+2y+/qz6TUftxj9OJSPD9WsBNd5wVB3t5oAjTauQ7q
IAP1asYRd/sifbNNeGcGznKrXVhON2vkmLDhPcqS8HT+DAXnx9JJDEB6UV43ai0UtnQ+OiSr9ILk
+/18LtDRdZMx620JvHfFQ5SDHs6M+/6K5tTxxXC8TzRRkO7I0e8AZrKMdt2cMTLoVZTPJJ+MzVvl
Gf5BW5w+a3xOi2+kpe5I4639fkiKcgTrwCvn+DbdzX+zGxBakQa12tpqjEoXAWY+GOD4ejt/KadW
R025PoRIkdtQgVl/1xqQWylcn94tH9wfzKGIoAxqEAKvflRbx1gNuZaOeFIPU4kveKNNme4e0GiF
0IUqaJ0vEgQb/AnLtVautqpA7nPi2llxq+z+Li1ccsAUpQgNY248mUnU3mkAELEPW47HrWuiKrIE
Vs5PPkiZywpivVwSs2aBYJeMmPJ1KfcpLSIjvWsr98lLZjc2hThkKpTiuFUGW/bDVGChiN1Jehly
ceJZZzt9hY8oTgn8uQXEH29xXjWRKb6GzXEHQkioEDujnTnotAtfiMnUf01iW74z2HPPWvmA77Ls
jFS+WyVm/bEkvtFjtlNMUut67uQGjp9PWFgKyp12QtLp857ikWHVA0h1eSAffFIOIJXCe3s9l+YS
+cFGjhMN+z33hWlbOqYaWrsjDFRF/StYhc7IWNal1Ks0BGEquum1bxRVQvQJEmIm4OP1UXfV0uJC
Bct/VytvylXujY0fYIPqKEvYKfzEIu/Xg5b5BVz2dCqkoB/o/wBoIY+uQ3/+u4mJzQeO0gi5ytb9
bLqZR2oOMKOM16Yfb7uVbhG8E9ijn7decPHj94pFuUk5lzAaQ+CG1JpjxqcXY1rvHxCZUsbH+zg/
UutU4i9aG/9VoG4aJ4SSLoggSdbdWsxAV9DTVrFIKk0KP5kg9OpP5BnC6RqiW+13KROgDhMDgQxy
EvCoF0zgnU/Qmm5norybu4aOyoWgzXfN5WoFqWWd3ecb4zEdwSxcEzvO5qnqfS+6uAek3fL+4LOR
RwTBI1Ulw+aLTK+gnH3pqe1LsdweghuJ5wgOacBdkXDu3SwxLAwg7IjL3R/W08nSUFNRftaWZS9E
wXy3cL5/EA7MfXF5oWXAGcR9CaINOtke/C/NgNUBPecRGoH3/KplJXPlKVp4EUh671WBgR1LXSQz
r4NGDIbYkMn4zrFTFqOnPi8LeXJ2nUYzYuW28pmC1knJnbOoEPmmeECvv8ki0OzcGsGBsY5qu/Fh
f6d07RaA1FEPkJWWtIX+X65ay7q1NvqznnybiBeaEqxksd+9e7CRTS9/iYVNhfLpSW2wf8BG4Ldb
C07MmZWNMtn4vslVR8hRRUt8x2QF4tiPkx1kiKT3zZuI9OJFIPwQHxkuWK24Mqt+tixT5sYyT/vK
kHW0fjJBhmsl6zwgshxhEEcAkTp0NjySB+pmBb72+pfKmnfLuhZu1Xc5v95GkpBwqPtwtM1/FoUT
BvyGWX1fzlTavmcXGqLdFDPkP8gdLBtaSqRbiNHxgDYUdlH2oeqqD5TaVam9kypgegZDfzmPS65N
koEgqBqOsqyJZeyQTd/EZP1b8/cNlj0vZODGcCmVTngOkqKNQv6N3v0UvSraSgirkkPsy5a+eHEW
4wCrtxo7p7nbw8PgVDYwvarvqw7gb0zvc2ab2BpL57TQmPpBM1sPUB4bdILDypo8+oR+4CmUx07W
otCL86+sxF28+cizEZaEkZOQlYjKXr0WktucQiLv+tHQ5N60cBJqGOxO1olfA9IijazArgqSPX6p
r77+Vor9QtFg9BCPoCF4aAIWtHWO2dct7MBobUlOdrcaFvYlxZczP3s6kvXZdAACFIFS6qjefx/m
laBoDGqfNlUE7HvyzoqENC6fgf3tTdI2KlsZPpXmZrfvOF4jQR3lO66LH59oBSvFt3/7ViKcAmc0
jQrtbHwZcsnKO42HVXPVcV3qgdCCGyyd8NK0vqQBKMUPpC4EfGI0lS9SQOq93rdjbFLuBccA3iGU
ozvSWBlws5YSSc2GUlNk5oYvt7KXIZuJ8/jvvCmGtWayCMf4nXQeI+xS8e0mHhnQVo8jweorWQio
HuSKn1c6LfGPbFR+vO3RkjG9sWS1SwkMkPA7lA7FVXvo815ahnBwd34pRLtCL52hB7HeryhTL+wT
SKo4yaCtwDn8ukkwBziIKvzI5ti3L+Cg23gkGDyEU2EpPoCfuAGBOOTgzO8tcB52vS44MzNJgDso
7wTjMmEgOHAQomMc5ksf1k2Re0topHOAIHeIKUWOlcT30UKSh7502FJIqNqA+4JByBZrmVe0dbKf
LlCqrRC4qJM4H4lE6AnpFAxCy6EVfFa5TTnvz5Hb/s+xW2EpCSTedNIWlW6yIK4vcDIsIYLzeNhT
2VRuKM3A9lHtkAQ3Lcft5zt87u3VMEeQyHJkgpBdYILMkccf5EMDSa6Kn7tv3FJ5uYuCvmC9t2f/
Fz15CN2A0Rf1MxBksLAcLoQzeBVeNQv3Kuf0EThgU7ejHu8Jhvh4YjOnFQbuY5IYW7tFPl3IKp1I
c43gUm2rpFTCZR7BeVJd41iRvi/IGlRDIgJpsqLKNkAujlsr/fsSNRpC73xx+uqjQ2NyyojmuJUC
cPxmihQ0OeOYILcSBGJycQFpRvhugsYqBlVpGBESviISWhJ+1I1WXn4bVel2cWeqMkdz/2YFatYu
BIA+66znubdaP7OWBc5qz7lfP3vBjGMLsdu9gSWUnXgnpe7vPAIlsxK7GnF0IUH77T7RwurHN8v8
dcm/RO2RL5F7IfJ/it8xA9JnsuEQjM9d+R9txn51BMBBrCY1PG1LNIEBVvP94PzO2ShU/f6ED6GD
cDtzLjgv9jWcjdf016lPtUY5c/FouM0PXOEazlpGyujIp3I1Q9DGQfBG2JmV+PA1ZAbSvjfaBfU3
nQeRrB19+SJnbMXEt7/1Hpm/17OA1jMSshwMZakyBa1aOI832qSVhMGYOIZIPn2EwwVIYGLfTOQ8
g2KFjFD+7xueckv7r+Ooch8MzWPUzvPw1eilrKA4E5usTyNFYH6VtkSj1YnnO783qdScOQDwzJME
qwfjfFATqpn4PGStMNDujyGXzMYsCbQ7I7ygkhmzj7x/nYuEGeFkMJ9q0CY5Cz4uLqYCQP7TjkN7
0/2QfmkBh2RgdcI6fJ1Q5C+RNDDc9WSEtEQ2dcK/4zWXv7sHxeeJi9TFvUhWbaBwg0owY+I6KACK
4d1S27vbW6vaqO/eJXFSTv9ysrTz+NA4xa211Ajz24a+s8QWYEkwEEllV1RJBc4diAm+y6rEfaPB
eXrfg+PqHvCc3UR6elHzyEwfWWLlSIUXMpSADMPwBJn1jjAZsXKUvh0J1CKWwrHm+0X5vWskj+qs
HaurmyOxCR1ci/m+9Wukq9Fr01aOrOwzXv/3qUR4JJLprdiH5S8+j42xzWFD8a5uuQ8Nm/b6bSNI
HlqkrrOuO0SLu5DR63F69ynaWCIdVF1xXC1Jr9+kjfub9rdm83rGppaWfLGx7lQ9Gjd1SHZvXgNB
wlo9xnsdtZ7aAlGPnfnTlLI2RNldFS2afnxoNdzQhnjlo5JRU+DmTwzYtLhtd1KxftwZSqDx/2Ih
ODeCdbE7xu4NewxZ2uwY6Eimx/vbXnT6zUsaYRKlonmBuey2MN/h7p9IX0uirrvYv4EwHIsOBlLg
mZvPGvE47CVt9uNiXmVNN2eYMK/JJvjf2+j2us05J5jajhPOpIXITuaFzo07+X0tLGI2qeHrICf8
nx3OgG206zrfNcbQRH4RlLNDCNTCMR9179YH0nfjSja05WePKPJMI5W3qNR1JFrvFxHxoJFy4a8V
5HB4bWdhGqa8518Jf+vJBCllvRMLTZHQU4NJgeI0D2+TZb55q5/gTnyH9F2NEETYeBrYEG1EOPJ0
W5TFq0EH3Ed5sb111YhTuYIT3ajnniuiL5KnRyf4E0i2PYXWUXjQUPLv8rY6Olz5pELC+j+chjHp
pMuK7A9PxvUCbX7riYobzGHcMCouBRLL2/W3axEDOuqvcg0u+oUNPdHo85N0pr8BYaHMiEvUPaPn
IJUFiA1ROylW1WMJvbgtjXzKK3VSy+1QyXMfJPOYdc/tlvf65DPpDmDITmLKHEQwhZuzjCeoqnpC
XVjEUxyX7VmnKe6fcz4Dfy3NHtuwrTY4UjRNWCNY7VLYeCog/WKB0VQKalwWomi+s+XPBysdhhXg
aLTXPuWC3ZQesljBm1CeyKjNtWDryqOW6mf5RrXrWew+K21GQj1q8NSShiFy/JArmpWc+2TSlv2F
f51dq2KwZD/J3uf8PakRhWzbUcBZCZFplYiqOONNy/8ikbvY2RIWgIjZlxd7jKCNzLG1zJMx0qne
ff5cbyoOTqmvAm/xgR4L9La2wNlK6hCGJmzOszFAuBe1slPIw+9XRkTMrhfSjKxHyQx98c8SlVl7
Ius5bxPNOXGMjQ2lw19KhxOZEeIaGP9KM2HfCLSF6SU50RuhzGFMcMmL7wuKAKeJ5Yf1HQJBx8b/
LWTI2GMywcU509ZWFfF/nH5r2A4264LQQHqAolXjIZhKNCuW0iUul2Tz2IBS/K+LXTlY9I0GEowy
fA6HgDU++KS7a46CbyiQZ2dHzqiiH3Kr0Rhm5pfO0AbyEwYVOOYkroFgUfv8teD66GK8xmanw6/T
yCL6tV+OH8tmbnSX6vb47v8HYKX57LqqUlfsu83QU29Tme95DqP7o5Ne3Z8ucadpW7kN5UlvfM6p
OYEPrvT+GhP67/HnGtgzsv6mtc+5p0My75aRKsi+RX1uQuQarYZiPqJ9Se42UUer+IlqjazpJRPU
7+0EevWqVPtQS+uj5UeLGIobNe5nsVBvzv6PdyHHF5jic/RDCScInmRHLfvYvKkhM36oKMgvzAyW
p1CDpxBD7NqviXkixVIE0SwiipXI8HqUdFXnyUxS4puP5spoQpVfuPQ0RSlh1EgOcZNhvzxA4wCY
LgRukQ5DY3Wc/YLlVU9w8DSinHdgLYKY0+n7X5awbMU0G1mHMUdfa7gKFmnkkMGwamtXEttaPwFY
EVIrC6eG55qL9LVtIPb7ot+88rtOJLNBMNVnGmcHKUi/jY9OcbmFkEnsMEPE0YZlhGWcMIY3aL85
AWX3S8l3K87a4ThGi6FaQjcNWaJ62vni4NLyHHXH+2GJOuCEeO1A1n/Ls1rq02+iU7jE33s4EyNV
gBPW9P0zefujC3ozraJfDwg/CfSDf9M0yHZtjAkBw/xooG1NJW1ze9ULDyPHXdOjS4smxmM7L60M
U3Ok47tmNUbhgGFoNhP+Ue1kWSf4A9gQYtJGVIfWfg0tlZ19bZHPjBjJ6Onz8rvR7PfVFCRR+STX
f3HrlAV0xDEkcPA+DIQJcMqhaRJHGGm99cEmJPFD0tdpPwjhuOpG/mUOGkhAh4oz+TR996Haab7T
ojdO55IvIf/8Sp1IN6C+xh2YK1KNiK20WB5u1GpaO9xxp09T8iK7qDuGkUORlmJIrt/feOWXhRqf
aI5Hun92qzdQBVgAuDnIsVP6S+jAhCr0R6zjiIhDnj6KrMT1Cuhrk2otf2i8IlJd7vE7+DO9QhC8
TnZuVgf/dBBSOh7VUWSXRkoiX07Z1DuOjODlTtgqtF+Q/XfHguKaCjs3gnHgxPMXYSVO2Vl0SULi
aVG2jTWDxYS8s2wPY0tayRVFwam+QJhZYtsSiTrnqDvFC/02QH0yTdJk9ysLg59ELT7jxC2y9KN5
lfTJbL8ZK6Wn9HY3qtHxF/A6IoPNkYe61/lXvPS6pUpGOB4M4EQcdVymQuR/Yx4kHrMC5PIQhPb7
/UrcVztv3QhKFyPkseZ8TtW9lfYQbyqiYk9CryP1hYcyXISKqzxclVMTntTRRcYMtXoQaj9ystcc
zhqZfrsH0f+deD4mcBqJoPbtRkP4jFhV/x39fABpunl+gnvniW/4c5hUWbWkzlEX0TW7VWvde/9I
aA7FmW89QkFBf6ZOTytxsl1DNoD/NxeZTUzwsugCw0zLh/utwWNfnnFpRzP8DKpuj9RU62D6IDV1
KlCmXOsltUfei4r/6LC0l7BA2SaIhp187hpw39o7j9BaQdEQkidPACbfoR0ZPoH0+2Bkp89luYHs
6jUuISuDurbl6O7zlpcAfMZDDHlfCn4EEnTbVAGIxftQRv4/KtFnaVMTR9YaYVk5h7SxG541ngNJ
HqcjpY5OpilExSTq3fJO611Dloi3R4v1aT/dwwvD9Cy12cjdM0X2SmbchMGv6vsqVnP0tJtGZlyj
dojugdaR5scPi7lscJshBhZXkyVXTrty6yZ+AFCR7CdrJkYq591y8jD/Q/3tZ37eUBgUtvzTHFqP
HnnQ+FHjGGCsE5aTDmHhMPd1G4eQ78FyHCnx69AvvC+XHdEkozo0I6hYlv2FmuGfGcWozjbw5BOa
sAN32oOwJRu1UNUi+WOt2oMdf0iIyvQdnZwj3RhdXW6q+BXqCgo0HJau5uCQS0G2RbL0QrrJqgBg
XFMWhE4yJff/TCaDlqkkmlURXHx6spCeawH4vRS+tGiSMUFdBxmghpIRjrGXL1M8TkUcFwa/OI6i
iR7AUZQ77oN2DGX0T3UnkqqG0dCjKrSrFv8WlVZw9oW0g/JQIMMtV5OM9WiuUTJmHG3cLeR8c8D5
FxfUEVi7QOa2mjgzHrbUuc7Ynntxr90Is8y1+P3Wi8+ZPuvfk7XBol8jH4G5615eY8fQfz8fi0JB
O9fSoKR6FnhOXCdEkbVD+t9vnP/QTosBxulev1MnYYvKC/jlwLwCfrvq17rvLasRGW3tUVTCEq9H
B6viBk4sbE4nkM9wBiPA4FWnm91KPxqdfDOqRrRLMEWRaSpuz2T0F+baWANWIAba6TRuH326JCKT
7Zx0clfp+loPLGe/l17vPpw+dXgQXkackRtjCiU+X/1+Oeb8iQdlswHcGodz06mv9nJVO6YWJOTd
opUa0U5ul9GGbo4qbMrM2ANd8IkfhUKqtzvvIKlsJuKudi3wSfxKgy/eQjpfhkNivzBQYXTusUE8
/tbO/Mpz8l4rxUVjEKZDmoDof7fdHZ/z2Fs9QaP0pzEs0ePiWR1ZCT+BKt9WvCBJOqrzHBlQb/ql
ee4Pijxf3jTaoHrJRcZQEiAgMSVf0hs5OQrEmv7HBp2KtB1LBHviJhW5PZK8fp+fc1gCcjsylb15
Nx0fLblFabvtqbBEoBWInsKqf/YB9VLRnwWBlMAgbylr9L1cdw9MSQBwKUpWODExuH1wsU6UHO9Y
aD/I6wB3pI73PsWuGx7cVQSk9JlaRehi1Rbv+7X4hJU90m1ZeclG25gZY7zsm26HROip+yBPQkIp
7ud4kFnnSkQ90or1x/AwxVWjsRuXbiO4qrClA09gKkb8A1SMYjlzA7XKR8jisso8FI4Nolfo6J9j
vkeV2sTDrmI0kVCCbiK2UkyaNipNRsUxAVF1XUwMvRSKGHaBUkKzrXRYONfNu6AiSZ175dW5UkNy
oXeSB4tM/96QDOPMnUMGMJQ/XI6GIMKNYVIcARxfidmkhncioSB2VZxlSe2SSNJa/jomf+StUTDq
Ytb3aRjdiCcOLsBx3DYOtyTV8waBc/j3VJPu+YT6pEPv0CDF6Hfz5NRjunEAgBG/1lyW1z82fvqY
FeAR+ru0M1VwjDChtfnwTqgpsqcvQYKbyVwRjafq4jabXCpxzH37S1jzMkN64+LkxFzsoLXVY8pw
IkioPt9C1eehQXXwO7EAgC7N5Ei7iK+i+HDSZdWKpcnOIqLwwm4FP1HFJ7q6Jx3GU92KFzWLcUGc
uGW/Y4MRBIQ3BOZKg+5TXeYTdMSxG6HqrEgREAoc6/bIFR0AoqH1pGbT32zYcFk7pZWEoHsf2tXS
22y+tQRpvEKTRNRRDQ6iibodF6JoArDJZeGNGDRAsWnfJM8W8d6ceI5lytgM97WE0Mx4STGm6Ebe
clCobKBnlCx3H5EXOcYFAtFf95GgCZPyQrIQzBWswlHS7M/JQklXpAPcZngPAK8Je71S2BYiNOyT
GsD2/hEx+RTpy3vX3f7KYKNJFiLXUElc0QVxYOBW4hSPsVLOLJOUZROeailno/ai6uFbdv6XPgaR
aBJLxLU7zmAq0/tuYx5Og9na26UNU2rHONpwrgOmYy0riM/z3EMHcOHXzghkFhVoHV0AhOY81Zi5
XemhLWOrTvCWTmHzMGaXtUHifdkFhwf5EOqFCUeJZp2FuxgR0qRlm/Z99IbrpzebH2s2LHksh3bW
jHUXENJiq1+VMYYIWtabBAJfBbDEcMWtu16Q9B1doHaHUoIYj5qKVpjllmD4hPQd8T8LkC2SNXWR
joWPmdcLWcbFqNFe/NYw1EbvCamwScCkDYRUexJW4JKP3wNBM4hbvlT0O8vsWVBIP4JkBb12GmIt
CLQTiQtD8/7K09HnAY6EBxXMvqHK8j/TNp8ik9Tgz1Hv1MEX6E4WtafCCIpf1Giwd0GdAic5IgID
ZOhbA9munKPxnGOJJc8oZaTGOoNANdjI24saC8H3tR3nxMvGPVRn3Y54DM5b9gvyTcUXv/6TzlSv
yRsR/0KElTXG9BUYiXajq7Dhig+WBnUshsSmlDv9fgcYITzM0+6oHKEIwbZMbon+BOqCzgOIqhNR
yUMVzWdQ3jHOB30/htI7XdPL0CdFwD8B9VnWzXx3KxWoaAVNBKYGJpedOjc+lWAqb3tAuGxfkrqf
Wzh2RSymmB/l3lPiXOtdOMb+gs3ssBzREwq/7Lb1frUPHbZIwJBFRbj5TYtOu0B63KpjNfx0/bVx
XEFFGq0KrLTLDJPFPMI0+b6M40MXV9YCRk85W1Ow7fvONijfCHnBCbLBua/LQGsryXWjiNe9YmYu
WbLJBARi3LWYUR+hsais+8GMP8+IkMsrGLoiVJm6JmaDsL5C8VGLfK/42M9Gy/VqqZAomzxgNS/l
oIZcsxXsl7/TcU7538bmiTm0dSmBto19N75iW1THlZkVR5gvXRYwYeyO209yp1OqvgRM7ag0mp3E
dQ5ut8qB4mWI9kyZmgTtMa1+4ceqdJ3oEkAh4Icd1MKQK1+MB1fCnNhQAvWwRLGWnTiiQGmCHgQO
rgYAlbbFx3LaZfmE6AK6+SUgx3DVaQ+xAJvzqkGUwwsRipOqH7oVYivxTQdQ3qGBwu5j2KepYBm1
YliOLwd4aQ5wjlC4GLX1TeH0xfPstb9lKm8E78HBnIKhdGmLJ932XVd97367a6N5p0RmJShhgq9O
dbaItTPWKZxhj3NK2j5gnQZM1OJXz1FvR1pw88PdAIW3MnrOBKnJybj7vC+sNkQuDgBlsH6CGV9h
JDMrmSDxbesfh2MptKGCI5jKDDRzi3dh56GHl1MgOkMLeMlX+FS+HTOCCqI0zAfA916REUbGgpKk
zu+I+2w5xoVVCqGFSO6xCzE980Ml6Qw78XQeJWKIURigD8EPuQIJZebslNJI2yUmB3dpfYdGWu/O
GiB8w5DaEw2nj2IMQDqVgq99k3JP1wwYoAgdu1L847Djb62GrUg/oOMn5Wr4MTVP8Ux1QuWJUgLr
5cRTckq9S5LQCRxRgNqzix8qzJjFmqPvtLp+saAmzVm8+tyfh3BhxnvPyT0S4/LLnVMh6sft8LXB
kKH0QhTQGZ4/cNToG7IalYIM0yyDEcrKrsvLd5VS0Cg0UPjXI667OcJMQzgpU5yD0Nse5HVoHfgy
D+mUHJn0tiqJkxTr3XbKuoA3f6cpJ8iVV0YgCQuYR7QZcl7CAOTzoWVcWSFXMpvdFE6OI0njZ2qG
jSNk6WmnGgSAnG2cGgJBNJE/QlhseR+fPDpwM+OOd31YQxAtTT1QrTo7h6+JUvEd/L7CvS8RjzfH
gt4IOnUJjAkUA/WeRN/FO/7NM9UPS+rh0CaubJRZ6ACh9EvjSFcNiMnHKLVgtZlUKsS8K94lcblG
w3o7mlJLSmvR9RRbWU5VcjvIYAgiPFndGnbzkBvanIVC75j2Jc7PoU1NMFJprgJaE7uByJiP+PMy
FNaDRt9pU9zpfpPnCzbgO9dqBBzVCLeMI734t+nUXgvFSh390o/vHFGFonXYRlkiLdid1mleLEp5
RlKIaULqLyB+Sf5fAIQNY0uHdZT28WmCE4yW/iDGI9V2SPSrEmRC6xgKa9vgbX67YtlhniASTTsO
pW2Cm0A9UAF7ybAZDzjbEVzyC2XqHRjcD8TtwuVFRTeFb+xxOpIZPhkT1a16XJrE2NiLMDR7DmQR
UeOcOXaN4fL16XVVKuruB+VWINvykIEhJ1o3x3KfHhin1+/j0KIi0kC4wWkptgezXwZs3ul2Mx5j
eps9l7prKthQTnMnh7YfGdy+HYHmwPQHPzWY3IlXq4vyZ7nfqbEGwE7mCjkfQSC2Ee5KL7v/JiKf
wfh8H2hHpyBjYEyCm/+j/vjkIzvrAWcbGERB9I9GnZwetKK5gcd/BwCIC3Tu+D5kf3FrnXb0Sirq
2Q2UtIRymM1ZRquwg2n3nQINvP0PeJUVr4ArYegTz7wKze+BpkZ3k5RKNq4CuCrnwXCuR/jF+cBh
9ONaFowESVefylO3pfZerdheTSkTIwU/w5M1cYWxO/bhuxUJLps9Tsm/kQk3V+qHCZdunIz403hD
Tl5ksMC8QYhF0HDL6obsz5uTXkzDUJJX62DFdAESApiKpLLKKEH9erjGcB9FuLE4kUh2merSF1R9
OiLYyrmrF3E8JwT8KmjJoOFxYwnDEPaPeolXoFg5Ya/mej2CwFVYMIS106ok6OaOt3gsoGLrOtfN
EuTmwqslDzvlUd9iPZOmi77uIIPTn3UX9qJ0fCR8Y3RnY8JIpOkOOQpBIYJW6KgE2Xni5jSsu+fP
htCOmJuLWGzz5g7NV74bzwqtpdbMWq41qMvjVWKIWne7U6m+VUocti5FXVQg4wks2yyDDkkhmQih
6r+ibeKElvDW1lmrwnM6kxWQLbXxyzU9OrpobfI2p5YlhJcmI/t8CrIhISVJjladVLfRMRfVoTXS
cvHpJuXOvsli72DfUu0+rjJw72c9ndob2iok+hjSDSfIJScfCNGtto9ZQrMCjOcx4vjMpg1uWvLX
WJwk1d8ob/n3nweqwsRupk2+5lDPUJBApoXiUmDJAVGQWPXrBVLy3+S/lbgY1a/tdatoURYVygeZ
hRqmLyytcx8ZfJXbRMZQ8aCpl8SUF27TbFW8nrYbP3f5nazL9M/VH8xfTEHmPoICMXcgFoIus9Hy
Vz/xmQFff0oJN63rtMR+36eTo/Y+Z2hlK+ZW2lwI+GxZ14Hlf1pF/A2eNhPrxsXvO64mKrl/eQIj
vuG6HQiWQDrxjzQOhRAfzti60oaIYgFNoWzxMWm+pkOHHFkw33V3WdOvmw4prABCvS4S2gczqhDJ
DokstirkpIP73ZGRzY85ZMGnMyzdEhX0bI+aQ1z/zxSABB7mRfLzxXkYCEbNCodRQsoVx3vn0qPB
moTye9bObT1w1qxcWekZmoyrK5GcaOCrILKmHq/9eGZzcafr0eDo2dF3HF7y4+8t3+tBjge3u+3A
zyaa52v6MvTFY5CJ5xTJjVmco9zcmeQN5ft5xg0++DulHLo/il+4YGTdzW4AGu8HNm60SzzDk1pL
EAhHC6lsI9XRrdWjmrqMxkmc4frwJGyrGGsF9w1mmRf5LyBRvXa8PHG8vxyanMSwpg6OKrdmtR+D
HdwdH2Dj2o6Gn2fdyIE1rJZrAq/fzxCVIpGsCB439E7XkkqT3EioAlgpwfmbhApr60bSQdmpQe5C
IjJplXiF0kmyikMiuca3KqkAfWBUxeiwYLAym6BY/1bbAyjsWyGu8WBYAK9dFTtvANWdTKN24kX9
hkaGtrnUVonx3lhjjrqgixsduc7M4fh0ufJ1W9NKxIofsjKbjTrdyylCm4bXeODMxiFp6Eofor3g
IYncaTT6kSnTrhv622mJz+pbu1ZQHBJOoQhjXLmsTbBk7mvmHw/aXjIKV/o31ANEgqS8RGHav/Qi
M705dG6vzOGEjkHolEQ9ZPF6EqGgrsYwLN6awDdNxEUGa+R+QVpZbXXRuLm+DqxuFNv8dXdrR+aF
qpZhidj9wKpx6N7Z/2YXFZbsCGhfNPBdnY0rTKD3YpJppF7HzyQtUpaScL70WTWhJuBovfQqLxkq
o5HNrTB9tCG7INKA2DitwIsw7kBWZ6k05k1YxQupRUxN8j0fctm2fit9le04PLE8z/qCBlerLTuu
d3H+QLtf2265bDSWtFUbdgK9PBDcBDZrUWyRthTD+JwMpVZMSU4Ix3v8iL4DSsFOpJW14FkWE4T5
OkKkXnX3vEUFp6AW4At2Sj1iNIxsCPVCKq20S2e6ysLTnxcFlxGuP8p8G12KCS+SfLm60Yj/3nnJ
7Zbi/w7HTYP/hsCwUPFMum8WFaFgnEh00aRU8VBPT7CK48cEHvDErSnFFMz9vNkpRsLkfoUYbpsB
cnbPjSJicGmBaZytCcoIblW3+3LxsE3Avh92t9WG1wSlgEwz+SjCoZP+ig8ImIn5e8aR7n1Pm1SB
0PNWiVMIGacs1CI/RH/tyu3Mw7KcpCeNQzrLcb7Ye12H1HFiOzPGO0RxPuYIgLbUY+OIJlrmPDZ5
WAlinkGF6zfOQ/3CmTC5L0OJVX0bpS/R+9zJeRy8ml51aWjhLPnEkX8y7UcpcJ1N7YAeL46PKqG1
Ib+Jp95BPU6j6G2d0g0g2UzI2Ldd1fr6Yfr44dJSmp9qaKszepyfjgWmnPZH+rJTWTY92w9jFvjz
abTfHcEJP0Q1zH/Sb00WzEk/Z0D+lM8geg8wmQiyMBrI7Gx3VjHyVVjkfk6Fl2vzd2HPN4FxJlYZ
hO+AVYpR99mNBm6xW6d7H47NWJHsEj5y8spK9c8GR5iSTL+puQPpnh9hTaOf0KGn2g7OL36IDxZq
ICsEbfsCHycODe4EEnS7iVvpurHza1FYTbkGIpefUX3tlmeorIcsDYZJLyUtLSc/NZY3WWVau02F
b0ksDtCvWhKPPLQn5BtNCmm8gZJEM9kEE22K1FJFJQC3DYL92EyW0prT7PhzN841CuzTgFGgHrj+
eb/tzM1P+7PznzwlKwUcQZgzZ3R1lpGsA/QS+G9EO5Ojp/PAX7tlvYyCh3sYBNA36NBXEg9CRFBu
YEUblBzVcZBZCHrBNV6xTlkqn0MGaQ9mL6KgRrsWG/oB1irYOTju+Wtsil2G93yhQx2h2z2xFx9L
LxmUlc3y4fpEGuHVaCJb3LeaLf8FhKC8GCDkb5BuE3/WVlW0Rix+H3dR4VFQtXFFKeyQLx3QSpFK
1JoJ//6XhZFHe/6ZZlLxPQuqGaf1mxqJKeL3pasf5PHpXMOeXuSniTiHq89YKylYJX30EANJxPX6
CudsPll6edyCnaqU2BHM9lA67nVv1wC+mAifN29WBDHAZVSQvCh8iu38yWYoluG95YdgQuVV89TI
7erIoz94+hnAVni3Lj60/UKQdET7ZuZOLOMZa4yOaFG9x7J/Eyzsf6/PL1vaItTDWM1HpdjcHIQv
bt8RfLHv9ObLhLyflaNtvd1SDLTmPDKIHWWhEncAJjuTr5AjKYqev1ThMHiqs8QNHJrkvFTZHMkq
bsuEi7+YqcP/jaXLTvKc8Xcbe978pFulS1Nd/ld2lQ1Mo5Ox9hyvGFN2W9ZdnTC8uhUiS9sn35e8
B15Hv/ZrRsyma/rNjImF00V6OwcZTAGAMRnhQksiKUPRsW7Z5BLCCr/nNUF+ZMVSAez07omrudxP
K38LdcwOMBOwsn3Dmm4ST9LM3/6xTjGZMYrozEylEyYEFbm1HbCupTZLPoaPGhEkbBxBIr8+4T4M
0Np4rRYehUIDvW5g2Fc6Sr7kCiLuOcUFI2gIkM0PL/3pcrlF9UCfkpiYDVhVvlt4r9/apoy3CCPl
xAzFj2G191C5RKYgMZxCtgeDmRi/vlZ6L5rw1nvZm0QUcPP6j66Zy/itvniLPVCimVkgXse6QP6W
eMPkNiVyNdYK5Dr46l+Y7EoyEgb6pPA+wKuu9pLv4y1GADZjLayLSNfBn3d6IZkpmLFz1ccVrS/n
aOZRUZB2Nij644V2YHnTjLTnvEXPdh6hfMxnLin/5h13L3c0SWZob6gBohWn7ghVo6mHuIQ2yivi
C1kj0oUHZz0qsEK2ruK6eND3CT73dv5BluY6xhvxvh1WcJIsl8eJLAmjqCiVXiaJPO4LK6UQ/d24
366SnPzwM/dlPxuJhQe0YYz8qceilBUKSz/MOyFDYTJljLic0YnSi2/Qhz6uRT7g4qOMfguhuevH
SkDo7+K4zDV6FxGefIZQtXbxMR+OGUImc8nekrvV8x8XKE1u+a+AF4pUCvUq8aYm4z1dz3aSI3kY
5qLG12439z9+tG2UoHxTKR3tpar8KrPjRsxG92z3Im2842Jz3iyB7F6xtMxGC8UC+Y91aHVkXojc
4ALzJ0H3V0VGAk0tdbRMvxabtuk4KHTEO1HWYkG+ihYBsGM5Zo8e7xCdktaXJsgQa/kq4L2ss/24
AhgRz7IJMXX6Af4tqdiGSJikCQGtApmVtPTgb1jlL8ypvWCi+kgyJ42i6ZManDc4DMvfOEW5llmc
K5/vq85Ec5uUW/VogoPauh0siOaRM8itlTszMufrbmOs2xN3YLkdhnK9Jh6ZaNsReTRmRJx2ibCA
vgXsmrt+2vl6laQTLc6ptP6XfS5sLXdp73Whv2i5/QIccBYMqQ3SAR31ABd0YnY1ta6eRxlvjx0X
bvTAVHdb8Ek+FOrQA9Lytx30fkHMUzuAXwUce9ui7/Zs5H6Ihkj9Bq43iuClPXqY/T+0JmPedZLP
E8bJ6D4aaN7uKByxKBO5Enk4aUitU8hWeHE+8UWW79X59jCX08WC7DkpwwG1Z4rYIWJDqgxKMB/Y
P1Ob8J20hHOQW77KsLUAlE0KSmr2UO/bZB6xIydNvay6U7SYd66yYPykSCUNsELzsk6k6Lyu2c8s
xTJMJ6JsbE6OSWiPkXypqeI74DLUrEJtxjDFGzHYDVQPI6c6m/XFYL/OaEkiDHpjK20zezw0ORRu
7OEVzfC3ybYqYqcvJWMV+Ko/+slzZJOMCpfma+c1Rpz1G34sEEfYt6qjoAsSjBSmbcuQDvQQbB/e
8u3Kz9rPdAUHFA9PBGSbUzfIAhhuuxNyeGbGTd2tWEyXXYl5Nlj6/EXxGRpElm2yC49ONR5OUve2
CqYEUlWP89rt2xXUjrO2mOuaR7pj4g1tfdwbl4N925Gc00QQrIzuunBxSNRZ1BlosEr2dGf5hKQZ
GkIFzylM+dgKJUqvsLMlL4DKj0SO0T/bcdKETtCsFbBn7UqXRhcCnmJJiVw3EIQGvu1lIqhw/D+y
d2Brvj3RR6FC/ebIgj6LOnVLzgzEhw+wOxAlnPpzl0PQ/n889TabbJW5RVb0QSc7sGc19HfG8ZHC
yLaMf1bq8uzLPIVqj2tGUBFf+m8hnCzE1K8BBCK9mtIRguCnEyRgCrayBrghCYqzzF1WLI0DL4oP
dRsEsXtyof2QudOirjsSDrlMPYlugSzjZtDxN8/hOUgVfczXrvAGuA+55bgXG1OMEM04NKmtHvZR
hc4dCciNrRjtzO70i7bkFrKIMmI5vKGZl4Ewp147+0LLW9zSl51TXmVLceKSpLYM98IPxk6kKXXG
ZoMVCRLM0LRpg5DiWWrIv8B0+XMau83eCE6doi6CcvZl1oCpRfDDeYqPrA4uaTiHt9GLvclS1q65
z5ZdQ21aVMqmpf6ZFRhNlcH8ATZz4RgbzL8XjHNQhepld6qrrRybWlpn0/+Jk0JRES7tOwDufvit
x6OIl/NqcGVaq+G1nwtm82cVX8pFjvCGmAgoec10pic5UrAuH9kE+KAfCM+v525yOsTErQz4itUU
lWto30zG6qY6xZ9BVDShE2Kcgx9g/pkZOg5LBd4ESkMy6K2LlLumBujDgd5F8+9h5wb0srkK1QF0
AWNwFg4lZi+umiTOavuwlBPQDBe72zXAP78EgYrx3jlwLL00C9HpgdErnFRjVSgkfkcr8UaAxrGs
CC4zTFlor9UTnrWXL9ANQNPYUIFh2E376LUjtongQ1vePKW3DEc33b38Lonn93UG/Od65RLeCnWI
H0Xv+lSQGojx+svMRwy5bef86Q+WtTW+C+mOtKGtuHocGW6fCdGjfpsXIRGQODVX4Oqe4Saqbjvq
PFK16AbJTRW68I1NB+Ilm2qmajI/dB3+KXP24k/uMOWGPc5WiYvduTfvYkVWy9xTRXUvas0j8k1o
JpTgpjV4Zn5ZdxunUFLIZs+sQIrlvMhNNfxe+ABAzQ4WIcWO29oy6x3ZEHCsIREs1H2kY/WwV0NM
dfx43cTwSYI1DlU80iDn/+QY/jnI7TK8g+EIyomTYvmXFo4JVfFWf7Xr6wN/wnM8pCkVVmwB+T8S
51X/I6r18H+/BvBagm9eiANEo6jdtMTiu2QNDpsS9GaMkUtNenwffUvNfA67cl9ar8BzN5qjpEFo
Z/p1G41NIsd5npIThxBdgwJ/dEdNk/nLp9nL4qhfAzfqqGfAkoeihPhiEt+uYW6rqE/7jsB8/Pcu
yA1DFN/nBoYw5CMDUb4BoEhrW2IPk96JVlTYihezrWHSST+abSknO/4J5e8n0aKkDD5fPIYa3S96
7znUeQiF5SAtAEjwEFGmfbXMCZucFvzCCHga8v8ABTWP2ffHm2mRey+50JEwXMGbeNY/tXqBj79P
C2bpEJz6MtmhFSuO8TKpIbOYdjgm76YvBGDZtrDwVW1V93mNrfnC5sZGBra2n+cxKhoRfkRDUGW5
Hzd4Wsj9Jap9didgjrd9YZh8YmpvQfMgn9siOTWjRDCvaaP6wK+T2UDLmy3Qqq7Dw5bcnjU8FX+S
Df9X+I0hoQCyMQp38bFMlGLQsghXqTvHTSde0vjIFJrHoKSQahbspjzreNc1SUW9ZhY0x979K0o/
DTOa/w6TwnB23K/aKBqawFBnAkIDJMx9CnlCe36QMQmggYGkgEQsUUI4QySdnDBjDyBsJmkAFwKl
CtGqqp9slJI7sTM/Y0jlDuUjUq5w/C2hDPIhImq4bNN+1QvQHCdu6/ulzccXrsZnXwsKw7vj0fKK
2wUWwmu8DIxaP5TSNFe7me21MfK8haa6XM2fOI5OtxAd9K8UgL29SOFuF9rmRyGNGM9baQ0X7PbR
WlckQzNGNUM2YoTx8YhNdw8mXH2o9urK6h9ft1bnmG1cKDUdZyatpxNq0T2/1d7vKx5T/StV6yve
oh4DYIeCUZe/dXWzOj0cANoK8QtiKzAvjr3jGSa2v8ykMhLMUbfVCIsz8F768hQni9tNZq0noNAT
D5qkVDPzdR5+ZJyyj5DnHZ9NKeVSkHHDzQ3bSovc226DYxHqJVsZQ2NWBXUEvS8gxdq8HiiJRe0E
FSjRJNcDEDguu/K+NK8hBYLhYl36a0BZMIJCzNoQLKFNaCEBSSwH6RBm/+xBZoKqs/8ZASYyXQoz
okkG5qvu0uWbTTLD5etZViBpNZytmCz6gVNTIOCpmjt8vOi+6PIIuVFsk6OdlAp3pP7JmYGBA1Aq
gdo0jSyWvteXqUdrZKgpRzjMDgEBROjtfxN07r1DvvtaE0jsEzMrJtfS9gEH47Lyrezr3Vr9aYIN
jY0mdK5d6yN6crobxueBgxm907lAlv2ZlR+IYlta7Y/RIGQjAN/ezlfLGWSoKQADv+Kbhdcj3gRl
4JjEXN/uHIauFwefpSfE5nLKmUAmoLrWeepgq/GAO3B0xRuosypWqLJMNRZjgaug1TBIadxmUWDA
ER5tYxGD3uduiQJh6cUGYQx8bkROmHNRLEkqsRlbl/6E2s/IEX+EUXsOfVSoJQeO+g6waZupgVRb
FF/bRJdrdvPPhBSAoQvTryBOZxmjgInasdEavTLJA1vBiZnqlZPo7IihLWhp6B173miMYdPAsKiM
clKgYXl7ujv4MsmPZueiIHN+TRwF1yWdEIS6oCCR/YHiUPr4Gb8dBOkIZFLhNdEsZu4eSPbphBH2
iO4pom1SHA8c3oSXlum3X04raFLEkz5h0oYDgikwFqYe5QYEqbsi+Gp9QmlvMGnTXq09t5srxBew
lXte0jkFg7j8UlhTz9Y736plV2eU2ckxL7ALbxnxaiv/d6RB1Q9Kr5JzVW0GRnraHxpRatZOewIY
Zt9EG8ZCTfrztLXe80vyKOdiALgYb7xm5Tmps4HB9k94an5+wFNmNf/Mc4wLdrmi5t/IuDNnXL6m
53aBI4cr6QASoPqS1qRBnLsyxYnTAQ//Cys5daslKvYUHhGZB/SThShPt/wpDRFhFD6DgUmHd389
abWZWLZ+PTpQm4OArBOPF7D+r+mk655LFL3hrlJcl26O0a6GiO1Az+6lgDHacZURwU6IgaDbxUXY
2Y7kobD+FV5RFH6YokOaEB8q8wRdOaBgFacfUF/Obm+g25I+WhQ3JHhB3RCYRFwgTXxLWx8B0H3N
CmKsMvZIMrfy+PVm0NNmR1nKb5a4HbIUu+Azt3ANdAj0GduGqMqSQk5pROonssjtBwehAMG7xdtD
9GKFYerJsBf9NDqRk6s+iIxK6wqv8IiAaxX6BL2l80NIkNQeKI3ivOImC+lFnyaLPcnwxbN0wcAV
UYzEJCG5v30laNxjTyqcEc64lUd6zooy8BoKBWfTEp+yO+Ncd6e91BNGrnFTIccBLIT6i/ER3++T
5I8NWYbg1j6mrgLikTeRK/cpK4KqKC7ocfnkxIA9UO4QdswvybUBZ1fzYxEp3l+ePlSYnLNXf5Az
3bgZdJ8buUHcVh6YJXlu87Dt5vAX8BJRWRdGYfTchJuQupO1kQJ6jjIUB7jClsW/0NZYZxsSrmO+
2Z1HyTRr8n317MUPC2RAFF8izipvuxIYIa7hKojIhLMCiB6QX8xZgShLKu3jt26s7eESgVTsnUj9
Awa+zNNAecbx7A8M9UDaJknPJpRpq7/+ONT8qV065h6tQ/zlT80KzE74v30VkO5MrB9J9TNns1MW
aIwgFAbrOy3cm0eFKzxItq9XHD8Cdo0UelNntdxRa2XJuJYe4nhNRb7m9CDMFlW1aPjUnsDBW0Xd
zf3z7g5l1gwxAieT8VuzOGg3AmNtxF/GQaKmL7tW00M/NjWd/R6VZXEoKg/UOJj9nVgo/qr4+CeC
26HmY6IFwfd9IxTJyl0qP33mrm/1joUCIFrADOPQ55DkyF945Xn9wgxws9KTXBOcUkTNkkcJs5kq
Qvt3BLI8+LRD8exC7xUBtSaJha38wLiJk3CTgVYOHccHuREEMRxdvXLR86kwAEMFgHvXo349TE+k
PKbRAK/AD9YzSGUjXohkh6KqGCdEke0kQ3gvamN7Av5K2q7m9wlmoP8uJOMGjjLWhrLvxCb2PcbM
Irq/eNuUKg7RO0lFnrDxzXoMDl7No0iUcpvIjQ9OwTQe7c1WVMNApzvllFgVMDzvUnTcz1ENrzrt
yEIpbPFoH76XO5sDm5TIbb89qYCEmosa2eLfNH6Wwu92pIkSlae8aJQ1HNJHFgRU+Ej1j8ku6jYM
QTINwXxjpsa91TMk+rBCI7Pq/jssez6+IsdCM+UXZ3T4QyYMC35s5mGN5Q8Gc9GWetDjn5hykcP8
15vnH8ehKCQTQQuhTSHnNPiAkLBQ9T0vilSnu+T5CyA+bpwymzDLd98tSHa5is3hzMG/3aP5Bigg
Jh27mcrRm0EiJEyLLhcAt4c32ckpVY3FUfPj/mXs+GV61DmP8pU7Cd52RcMXpRK8p9awfsqK60hV
Q7pD5v51l990BPsinaZqiKOCdxsfrI358+zi1BeVAPdXge8EQTIPMnPW/ZJTCgcMnQsbHnTEXRYi
tnV3ma55qa3q+HPcyBl6W5jmylu6xRSIX4l/UJKtyGCNj3sNS/VeANgqIONKqg5bYqQ6Rjf5Ei55
Fqwkk9W4fhyXNQx9XctF+dY0QQct9+w23meTB1HNi83hFFod6U9EoJgZTbhct4ZL+GyM/0GFV4m8
3jvhS5HdfTyWpxqYjmABXRrGl/w85s6LSHkgHZtNhUifgV8DHuVAFiu/+3kbdT+fU49m35uXJ6ZQ
sFBw1u1IRlJMXEU3+0wiKry0XfMAxoSv9GU4M/vz4IMEN6YjqvIu0CrUADFhbgcjAE2uopyI/8i+
WxlUQAKJCtYjmtp/twubI6mOKVErlKY6FbOgaWl7U+eEEV72tDN05eCqsiL0xee6wTIKQ9sPH0c9
oYiLNRlmUCX8VzmywI67fhq3Z57GMultLdHg4GfLJXmedOSDq5yImjS4N+7fPPFEMaw0g8K8xoZT
JMzFn2muHpJDC7WYty6BSwkLIfvHvTSsGn3wKEgCGQp7uFJ+Sc1+9AFKWtJK6qwRe/WYp071uODG
MGOflgK7IVtQeyvUPF8iQ+Ixqmh2xnlRf3PG+ftSdbTjSOpT5YFX260hgI+uGR2/9tDmLWV6IMfd
N3cJO1oajMBS89AL53142OQ/UeRtyEvtqGvx7g8dCWKICyZcIgI1mY64VKEq9epGOK+ZM9CALVST
qLHh5bNHk113A3PPMwg+pM+GT39+klfjFtEfn2RJQ8JW+loElotNWg4xzvj0T+pTZb6FplGu0z3h
sHiQo0VSHlK+RVC09xURYwVOO2qT1X7J2JY1odk5vALLwU9T74m8hm+7r6sY1oazu5e5rB27dPYD
P02+QFtxEiFM8AOzTraMEkPCZckszzDZF/1THjwNl5amilseIz6Ra8MRpN98ldNCBoQHL1OekhF3
+dFx3UzfJke8DqdN8zdML6CmRVdMpPrR+wkELT5/YC1qRABDXVNWIVwfQtwq5VzAJ3nY+FOnD8rG
W+7ohI57XRgY1BXOQn31+G5bjvpaYK+0TVB+M+Fnazx4bFsOIc2T7moOtDWK9rDUqukDQq0ZRZy/
wNC6JW2+U+uzKAV7jWkM2h0cuLo4s4f1ikWBWxZzgpLSC5UfargeJdaMUXFs0BXckcP3u54+J13+
SS37w8BkvlGSP7IsJN74oYxFjasRFq8w7PbN10G8RHbSltvZlmKPHEfe+Bgae7zMAk8TafxZBlsr
JlocP+4gqZaAnHrCx8UATWCADyICEf+ys9YvlHKlx2t5s9CjYsLRCpdsdk1WQB1PaThyy3cdT5W2
aeluXEk5tnMr26V54ud1rn7J8+Bk632ZXtJASHxzEgeimbWyuxF2sGJPLkuMV6gzggDkRp+Z6jRJ
KSKzRFY5rIjztUFW895LL4N5owa9gMzBMppLV5il0k32UmNNiW7p6EHx4VtE3zmY+GpsZQ4DP0cn
cF9SrtHS30YX4ILwK7247YGhnSImEhA5F1GxVDhpO+UmoXPO2e9Okp5Qi/+nr0ndvfKIrpGOAk5y
0GZYXUVZ+bGPeN4BNVOwOCyYvo+BDLSwuq/OmIGBsJz7xUPdoxKDiAM1iKN1H9VY6dHwdJNxSvKT
WMMYPj3BKRubcmnRpu0AMPuAA/lBkolz6fLfU0Q5G9ri6riYQidzlf3zAYQzhPlLldFQ3XYRzJqG
zLk+RyEWNqKyZJoSKm9ahY5y1fiskF1IdPXBM3tvrFndHTrxjG0YgzFq6Jel7uplK6u7wqV1OG8S
Wf582mGaRho+A2tMlsC/Mojpha3ODcxFDSZNxx3XXkKnIlNQX/wkk/eWx+EFbJ4szgl5p53kx1Ru
B43siDTmYqsHfPx/+pKv3AWpxkr0bxU2Ja9gS/85UibO+kru0Om1IZzvsNf0rLRpWZp7K5suzp5v
Tj86dHWSCiAz1crxdhsalmFyyDjh/R3Qxd95EUQnZDH62bJ/fK/0dpe1sHQTv9Fe9zF97WlFXbJm
wLXiEHVsNNgt/tnfHLB8V7wbzvXVQ0qEXYKPdNsqhebsf6PO2lPcWsjZJDTaysNTXRWi66Dkh+wg
54UwN/3PoB6cHST571FN+GMzb4mm1QT4yP+XAdADg1vit/yci4PAkYy5ij27CDvmPHcOsFbU4qhm
AM2EbpZ2LpBmrdQBygi7PopPUaLjyhPk6zrKbXbmhXnc9tAMfe3iZfHggLJIfat6QQg5LbfO3swW
UDPy+bog2umIziGX6Jt0ccj4lSijG2khy0Ohtm0EBQ1wACa28ljV6zWUmgkFHg1B2a5Opy5X7lWY
4yBw6Uvh3GJxfa6Lj0xYb8jL0w0fOcGCUx8DmCoFDxkJz437lPLeYvaOvymFll2dbhVwYizVl4r3
CRkrFtvFWAtQ/1pe+cSNID/G/a/KVK8VB2gm5gR4ymYlMBSVYz5im/397Dq7er/6WoHnUy3tR9V3
GSzCBGEmVDtqtHrxUSgcml2BcUFssljF5+oJ39kLs8Xw5iotYCrfExft4aOT8Yg2sU2oTEQaS8p6
Gb+Pj4hntDL5yFoXblVjmMzI2tfbTtoIwiUko/D9oSN0OME+1PgF2alKv2qIsrdZB3n2aN62Kju0
kQVarAyyaAjo+BwIIwenf/JyfuX+GUL1kJ540JDMOYwRudRu7m+6ZdZd+W1sv4VW5r5ejX3E9DqE
3OHeasDUMMMdo2mDl9Tp1gRK+Zm4ukUN8qb/I/tBC0A3xalN2iJvfncylRJcd8w964r1mDHV8cG5
Y/JOv8Fn2A1I8eB6ANlDyLDralBA2qZv1jq9NnsreMBW+HgKfRP7x5w7Tdmc618wgioVbtpfdLqd
07GDFabs4R9ICEjdAVodtHibLwVmJz+H5sIA6QBlN4X4n7XLbKaPYdo3zwdRnzU+U0TNTjIkg+00
qhJd1M4Le32ZFfQU4NHXKT5AlMVCwCTMeN2NSStF7iDg9pNPceIDG435Vk9JO59zhw4cAahhY7cu
vRWLN/PagdkA+mSaJjhm1LNs1tVgZltwTNbPebJFgKVz3ypuzGYNZ/Amr30TbpfSvBACtRGahQAb
psoZSrN7jGyukVdqVzKt4KBIji3vV3rvk6clVJKSO1smrKe1IAHpHQSCSxc876TWTiBBInNDcMgr
kov7RtsA/kjDw5A+Fy3fngisbPWRXt/6QxIlS9pNWpHfHRc/lTyovO1S2HP5Kr+6G7iXDK+7W5fB
hfcXfrDqag728PMRv/p7LnLIA7nFzIYqrP41Ryayn5t6UMzShfpcRDgx4i/1Dx7iV4/IANQ3G26X
jS9eeAcnsDFAsk1P3RA4nMd39YVhVGVtCJWdVh1P3tbUZZaAV3Hpv9TSAiQVOnWJCtWpA2763Cik
VLA0nv1KgEWC3CibIH4HBdRlmDYW2jqdxWbHrMsf9kIef1n8IjWN7hTCcuedPE47cXp5AMuQNhr7
n7j0YjEM/UIV09IUCpL0bzlY6Xx2ebSpV12xwpyBaTVGtArl1aKnb1P2uCOqhvMfoUbvzmDCv/oQ
c/GIK1Qmot3JUVe/dO3LAjjR1P7ZVrp9ajrMhRTDPOSV8Ljn4UaUM2rHC40yh02XsNbgriIWN+1c
TTJfgO7ayQWAj76A3ojMllFPD7Wz2UqhePFfaBjdoPfArxFS+P9vELx0KZ772lIHcyZs1m45w4oa
99MiTSiiBQEs89YVImMPhEEzRAto/wNuQNYKFBIxmrkkPeQZmNzQPu3yqRH3bJDVv5Ue3okwGdzP
MlcyF0lSAWPt/KlSi2uZnYvWNvgiEo/FZJvB/oTrnQ474DMjPFDtQnqGOtSKEN3TmBhq6nY2WPM5
Of0c2QwhiJxRApDsZ2A956E8cohvyDS08FoKhbrNo9zqSQ4OvXxiCBVhkr9oByrUFeYZ9uK+ul+2
iRiW5UpwWR64xT68B/PfBWe28SO86PWQKDs6sKP4hcF/vuEfB3N4WXBnlYO9GCaprSig2/qhDC9D
+m4gp2SezFyPQbuz4KP4ncbf2+v8lr/ctRhc0vXST2KFKp9P7S0fq7s39hBjTMzFNuWuIG+vcJKj
oMi2+LhqFS7V1WZl3paSzQT8cw9q3CAutPr/vJyTg0U+Ac3KXVEDg1SmdUxuntbK5BvvPobosAxS
SagxMUzDKANgGuwhKWUkBJ5Vle2e+DelgLhFWrrpDKIZinLIhLoq1NpJSkZtLxASiHp3FsCqo4V6
pnAImqQjm793mDUsSJ2IwqIIoG+8k1b0KhjkJRd/zUEnDVV+Bbfpcu/k1lvFC3WJ7biIAsOt9iRV
6vvA2IZVYipIFJkw1tbS8vVrRVz2NeRHS+DP0BA1ztHw19cZrbOTRD1r8bnc8hVNP/S9JzlwSUJt
N8Ofn5bk+CGds27BExA2Idki55a+6zaGba1Q/wDGieOZf7jgWtgNBMXgS60pouGnWp67uN7PeOwi
QrtP6FJQ96PIiyXq62/Ar5cmfaPOn1pWTQl962e9kSxuJZsA4DqT70zwI1rJZF0MdKAawZwNUOzK
VmLnzLBpFtdA7jgY09DBquXQzYwzRKZ398KyRKz5R2/AP06GGsLGmSvZusH03bknShJBNH6hcTVi
qe4TpsFeqbGwckNRM0yWfaeJf3UbCIYx3wcfTH2OjngM8tV2Ct0o6SBEUsFDdPn3xh36+acKMhjp
va1ADB77t32pXva2qY7GS42chtKMwrBis+HvLOHgm/wP/3hmUX/mDskd2NIVRwB2miTekYYxFmP9
9VX0P/s+LnyWknq4qWKvZtD1P3JijPQPVbCcZBoAfpvdO5ruPZXJhsNd5iL2dEpd7eFHEEWmEoSB
iM8ars0QJpeyMGfENCR+LhQXnhBdBiJrbhzNMZodGOi8Nusm9CDSw0R7w3YYW+UvbLYYbHR0rbYG
f3x+xnz+2XzAJuJ/XT5Epe5GFje+bjgeVUECA6M2CAU9OBkFkWE2PaP2aypgbOZnRUmXAreNUQDQ
8JyS++ZVP6MaFtC/mq86yRainQPkex83AudkDMnbAM6kEl7TzZiI4YWTcm75xNBzcQJhpuiChES0
c256hokKFuu7RuhL8QCHW/hIR+g/0OLbnB+2hGa+i2TBcrMtldzDk9f7k0TmH1PTXN6hhIm/z3Rd
42gDHea5aH//IzY7+pv1pSVcyP09RDyxHY5KcdIc5u/SAtKd2KI8YLVB+YpxB0+hMOvH7Hi4O5R7
DPA5+8iaFR9U2fvv/dzdaZVvEkZszPxKOlA0t2I3WRI81bxUrUt/UaLom+rkwb1gpWid2rneHWLf
yDdp4T7mjiPajG4jGXsNE5ZwvaZWws9Mz/gAvc4pjO3CcpS6xSbGrnDNJ0S9TeYrKBXL++09r0SP
L+OvS4aGVQnu9rgXcDD6NAvzrAyYGbNkOa+R/frcc0a7RHjzUwwC29GRaM96NFkEbchI55eR9gr/
ncLrashhA6GtDOMw1ck7HZ8ZrpW7yPdViqfGALE5fRWXYknvILNoH7h3beJAwRO2n10rKFf7iGAy
XcuRFquT7dOAMzeYLWfugaM9EzOu7QCEXXhCrdzfhL+XFADADTPUQvE7QlBRsi/He7UuAIZLPqPL
w4Q/qZhM3oM2pdpM2JEBnA1ROMDK/PFS+XP+nxBOFtzJaXO7zNr22rEU9r3cOjD3Xqk8o6trMx9U
tQQN89XBRj96KHF6z6U0E93OvXm3+3FsmlIJMyubKE3jqVjQ9o1ZqOqF66s+AS/+KPffvMrs4w7M
plhdUVhgEtxgmWkNaOmO+8SkHPo1d5KGjGCIcU56/YVLM9X8A4uE5xSF6iOiJi+LMw+MfUgQ8zMN
9jteosFIkIlf8KvZhFnsoj0MSqYP7Uf08NCfWUltC74LBK/lkqLNAdPhpJLiXViYapioW28fvrF2
Z4SPPjJZNAyhBhhHl09aXQNLLwg6S1DfUfHs5KBogHvBIvxrNeh5qzo5dNVuRuU2B/Kr+STPX8hE
7GOUWOrnAhUOYxsmpvmtbykVyyVg9AoLJv8MALn1qBN8oXJcuKpZc8qiJVO+iGN9bRD7xBU2SReu
mz/VbvbVQdiX3ATPFukM93tELLxXe5A5OJ5gqoyyAlihplXORbCFVhbfWw9lk3+oHKbgm5o1aeVI
qP/6M0XPfw00Cm3BcxuwzUcg3TZKtCxgovBvpwe9csp42i6x68tOprRixsr3y0w+bCDE8nvwXJMV
YDbPgYdxxM2MMEorc3oUos8Dr1pEVByQXy6IvI0SQfQY5sUmwvIU8YXTXXb5NNpDJ4V9UTw3MT4q
2N8jYUae/V/Z9quPMcWVt+pI4iJEd8qLJwYr3hC9EYlbSYLY+kmzsug1WSqxrOnL4OtGjb+gWvGz
YTeId5AyrsfCHg0UN3IJVw8iSoiBBj7RDbQMcFLUEdydfVVDWIOXeeY3EsEF2kK9zpzziu9caxMX
FEiQ2Dvv+J7CCJSSvqo6Zbejg+RkCD48rbFDYV67WAQNSf2JI0VL6z9Yq/Xt1Uovov+lVwapwzZI
XbUwnUpoPlijZzHRJJwCn4LP15WqiES+Sv+0rYjixQog+e3QGehhdAkb4/byylKWwkF8WAkPuDJc
L4pVYwNSsQw8o9BIL9LwAZ5NfqhmuJo22tZmZ/knZBjxoMoujZ0JUm/KzC0HVYRvWfmMMGxXG7u3
HJzYkHqK+sJZGWGhWYeiFmQorSF8VzBk4OkcNBBscrAx3lYjY3dur3IU0ZGkhEdZbIEqwKngUjSL
M3xprKawdGaTUsfNOMIxHnePf7eAlyqPapw9KcyIFkd3O3q5oekMz3R/7dUgqEb5UDZTNpTH1u9D
5/yJ9c5O2luiD3FPJ9Ech9APqRvRMIKfgkxNoGYXk1vB7EIUccvxz9Q3uCsDbkvtr2c6yA6Hzfj+
2Xa/UiUd28G/mOuWv0j9H43y2AnC9AEnK0nMQkZsLPOLY/gOCB5b4UXait0dlLvh7iGukkPkCesb
fLfT9gRnEwIxK2SToWwdeASVfDKdI6OYz1jPWvzweAVQgKJMKFRaYzbqz8rM9zyokwvUTAln/2jX
JYgvxp9lI3xRSYmQtQ28N2bQGiNwosW2lr4vFQD0gevHMfbOsJ2IWfag8cD39v4gXeNvOJ9OuvHf
wKcUBnpJ8NgrdL9JMepI15e4l+F6iLbsOzHbEt2IUFIQFgsIoY9gbSJsArUnJ9l2H0hko4EQGoBX
IVhNJZz7yTw4twXKldSmAAMb/eh3oEFOqnHnQUwRDC4VPH+PA+6Hz4R7TrYMn+ZtrZehubQMMF3y
6MHIoFG1cyjGy6xx7zDkDX70Z+ZDjYYYU4k7jEzk5if93AsqMnAzLxP2tMXGuUvLFAD4QXYilETc
8Twvz6K8AD2Ub50BUjNArk0HJcumH1jVcsTit1yqSGxi6G/+U0psWCiFxqqKIFZ23cpV6EhWN4Jw
QF7TiFk2WZzVxSzbE3/0RWnrOEEwU19UKypI2Kt0aOKVVuwVLIz9QlU65hGBOKNqvwF1BAHshA/0
b9aRqGnkV0gcJsaz2dS/D+t09gN2sKE/CzeLZT8mp10sMGKRSFcTtYSKvVpVe9iSRUADHiQeE7ri
eUrBmlLeYYGEkXEbeCFQmc1eAWEb9+WV7eS+5jYHEZ+Q2reSN7cHptySS/CUVoN7IYs1aAkUKat0
vLAlIbq6oeRUyZjHf5ExavYmsOILe2lG1haHnQ+80L3n0Qr4c7m/nOdQvoTUB4T6HBMHJMZSkoNL
hcASbfVPgk6P2VWHqYubYgztqLTH3iQ9VBH1zxQ66oiKsaAoZchNtJVaILvxzvN2fSPJnMEhJDAd
ExjnOuBK9TiNit0D13TJeaqauyuImY4DvrSzm+thlgNCfb+YbprpwR6eAgd6tjvkhx0G3WZSIas8
Vhvd7x3n1kKr22ASvkq2TKMhjL6J0E0TWHY3C94+pbwtoHzEt+ZIa1XMg4OZD+lu8P+yMvy6LMXv
pxI+T+nnFwiTrWaB9V+4z8UVddaHiAVcsBOHtnOAGS+nrW+gpSVSskbsJKachv6kgCWE7c5VQGzn
H5SaMD/w0/dPc3rpR/GiJm3pQc+Wwv4OeoOX4P0RdDNgFKNY+DEFVMD6/28QzmZkW/P0OJcPs3ly
blkxLKA/8zunKHrDS7quug/f5o7jpwrc1AN4XzLzUn/CKWRxqoVaZzo2M0JOa6nXeIbkztpA4ZTp
fnbCMQAMorVVbQMdu3TSfXvhT6DIIQ7WL2gaggNZU1v/hNaXaHATz4WJ8c0f4rEzYT9+yFhIofol
P+/BhU6hCmtge956QDSV2SZDJqKGqF4C182RAsc7+IMPDrPHN/4dJRlpXhv9KK6vLlE5xubGzW3F
l2lN3Y/nchrIB18x6TU2D2rA9ibcOEbgdM0Y07BL2zvEqFbRJO0SfkUsHwCWlsRVUByff8mTYgar
91eiMexmItzJulyFfD74z3HCX9PMiq95pvwuo0SK4a+iVapNikWuJETt6+kCRBY4bSpO5Fh0BKgp
u7i4AWMbosXKBM3iw8Z9BRm0OUXSgWGUoOe/DQM9adZwTLOznHs+YYD20ON2QtBwRFHePczMqZUu
85qRNybbjptJZvOpsXDuuCW4hXjrBLDrSKUBSAw5krtmrqKli/N+T2e31caC20yp8OCPFpAJRpZO
+I7W/vSWUW0iMNTfnGZ2zJuqDmGdAx9j7eSGwxnplCnXTa+jYYiD0Bm3XNueoRIfro5OE0j7BGrp
xMfzu8t0Vj3O12XCykcyzojNfsSjP6aau+9qTgDktf8KF5W1uqaoQaXcmbg9n3iMISxN7L35uM18
SV363K0w3Vr70Nxh2t7GLAvCUe520ZnmcjeZQRHD2gz548AaUHtY9jiFfZ6xJhOH1+Tyfpu5ZTXH
Y2zXkppAvy+cIshN7rMr24ngqo3pGgug2dqbN0zILa8abqgBfhEENkquZ8Wk+LYSD3FQSOxfUQYo
pbRx6ECdLNeYdPVse6r5NVqgh6U6YWPAUv5YnyDpWiE/25nV36oIXH0MYER+gM7t4Ji5oRQaX1q4
hqeo7uqtXZbyo1ADKrbC6Z1JgqfTWHUuJslNrJLpIOuqqToV1i4dNC+w5bwnkHvKHOdFAax5myEu
7rjBwDq8HE0PD77lcVK7doi0x8+fcJX7ClXbPjaGxFNh2PPEBYE9lKQOHg45+LbiDHSzSH6FBoUr
jRiVtx7FafxNVA3LG83U5XalX9tHqszArHHaninIbc67QRR+8bGEtV/DXKbY32F+rDqxC6ErrQs+
j7g2+q+BlQWkbuTmuJaB5ft3Y5MsjOa+Qc6GAwDh3KgPN4gk1WDByqPMdBWT5GsV2KEwd2x1KdiK
2uJa6Zhqa+PMH7VX9LNd0maeuMZ6x6p0yh677ZrEwkG5bHDIl0ieQh1vu4/G4xqcVWAf53DAJqf/
V/sjh03F4Hi/CavXNJeM3IxDTP5cc0tVMY2l3bdZijPuqxexrjLPFt4Fmsw08saj2Z/hmbkeQ1ju
7f/6OsIShyfqERh20eUcPR/6WTwjyck1Bm9FfowWYpQTB540x4MnzeV9THAZlR1gJXjBoDyZLz9O
3yrG/OSIeyleY4wsZrDKN4xVqDV9tgwVks8mBGRNPT7iIMBWdJu4eIpHn5MKYdFv31VyCDGHMYNW
3zoGLQ5/Yc/7vEpIQhCGJ5KphhzmgVeiscIxBUSvTBeSQGfaiXMDyaQ9w4IbllIq55JiMT4GAQII
5FGLj3FrHOefgkN3aX+VKg1YYlgm2cxon61NkF6YXZro80MVTFBo727p8+rmZRV4swZMPrdh7hgK
LZ15whxritBh4Ar4Jz41xQidzaVN3ESOoYh1B4YSgloclpYkRnoaplY6u832ngbJbmitrmTdHPVI
TI/d3WCIYBvYNS4/7ITiiXnCoQin0ggv1nRwsMMIVQ1VZoAC5h9O7a71L4Q3uqocWqBjWk6W5f/C
lP0bnOWJUB53xvKUKA8qFns3PWb6XseybejxvBa6m5gYRS/OT2c1pj9mhrP6LhmKlrpLI8YMhtbz
FqYEpv1Rrclkw9qj5Z49eiNG7ZhC+Pc1PvHdZBH+eRHljYQA7Par7YmnMhZD2OJAPa450Ff0+xaC
s6G0ZWjXMDJJBX3z+05scsFNweN0mA/RPD++kaTw1pwYCaxVO1LJWj9G408OgmfCNIAhKt7w5mOl
mASLk0OBd60eVLI2us5eF8mEBkWc6+DC3Ue99HPqcL4695O/eV5QuNLLdl2aRa8KsRIVXnXrYurp
foydGDi7MAYV23Z03kTuFoxS58NS8E3s9qHQxPxEW1TU/VdGtg9Xws/QyQitSbpWol+XLGeaUrSz
FJ2kSewoGCQUXAV4zXri73LGmxSrWaPAvVfb7KCAuF6BuydxKbMMpYYB05lqNGVbJhA9U42s3f/n
u5JEpxJGqHBgrFWaB+zALYe798k5d80WoCwsvUGe+E/4DIxlRpxRwMh2/E5VNttTVJqmff3YfHji
tIpgNsCgsb8anZCEogprMiLpaehhL0kjWxC9FczYQCG5T1lhrlNASqnEhgvWBvIRI4o+E8bbt0Ab
sUzKLoBVBUS7LXt3Tu5IDPKTjplFJry2XjK+dTaxPkxEwImZbWiqwo0pEbhcy/hIuGkb70qIWHtB
2LZn0lLvzFMxAtw9LMpiPk4JtQZzkvwY8aN0GhdlvHZ0u5U/uvWzGsKdAY6n2T6umI/8BfknbpHq
FUnhwibHk/PKuNVo4tj1YIZpbk65Ur+07x7Z+xRIP+17lMJKyOQsXdOtjB9e99cm6pDg2PjaODHY
H+iIvqeYI5BRaEnPhAl6jxFaDS3qBOF/EdpLPEKCKcun9et49Pc9mgWiTZFOUEK0E7HB9FcHACLF
QU+md6A1SQemVnt2cBqIw1hDhoMYHG4ZtoYM5K10ejnJTJKVijAX5DWk4JohV1yw38zu8zok5VFP
pDt2PrjsbJwD859OHukpaAWgtFDtjvwqJyk6F7uwEFCVnoQi/pKrVK3t3VXJ9guvzJT5po9ToN0C
+3u9dDj1Lzxe9so4GR6MrHoJ1jXcB08b8s8isz4J8xr4rcdKiQ7zub36EamYEAW0zfk25sHGIg6n
q+Vjaa2fdsSq/Tnr4GpgTuggA2+jw5eLjggbX/2Dn9fooTlRXvaTj1Bb6Tw1WBsl7i+IXjCj8FBk
J9roPdtxCOCoKbH1alJGPHgao3kq/53Qn3ivmK00vRkyr6UdtNFXKNt68oo0vsqMWKz5+4lPWV4n
gTnkVf9DgqaPdmTG67qdhtiYdY2dozDDLGnwAJyzowKP3wysZhDcMsGYOKqCNAr+kwG7Bp+tew1P
/IedcTzAOlWIX0Thu48726bgY8x2RIri2YBHQw981f8J4Bg0rcQ80Ur80zMqXU3NiNAi8djSSRtc
+FXvX9v1N9qp5CvE5bB+OTVvBT1ZFwDaxY+mCz6AFISuw3jQMp5vTEM84QCLY/W35VdcGXlD/+BS
JljsZ90cN16UaotGu3KAJQpBBOzlIp3t1XvUllimOHfjHZCvXsEbgcOgfBVdI0jNKyMclfn01I1C
B9tMR16LpvBLOyaQGtgmTVZHHAN6KWJqm9wCXmapVMH7wwrHZepHdVdGqjNf7dpPEhE5SPoYT0S4
1s7mqs4thYYEYSCkebJsgxcpXvQAF4isb4uz9OPRon0kEsyBd77hiNAtgkd2m5qPf/XLlAr5myPI
WSE6LO18Fg4ER9uympVcgsFTxKNJ0vDSZS1hlwWcjSp2Y6SHJEy2onxPCGyfWzmRUvuKO+TSbid5
MEMLbLo+/gWKOh4MebTy7KLs/5E0TbWFGwpAU1oj4xNwmrf55SIfw9IyGSpRjqk5dw4C1AuGYeRR
l1tyAxZzBNfDFQP5sZWNGNOLmUsoq2WW14ZsNrIReknp8whORBoKKLMN52d/6LrzzfIuV+YQlXrA
qOQAca/OZ0RJEFoIg2ym0o4SCS1Nhr+adUo2SBnKg3y5yw51nW/lodxH+k1cAKeZNtj1zeAUVJH2
Uk/UlFWaPVPq4zFb/Ev0kZahuNFgzgsSRxh8PfGngsNZzmp/R8Vynzq3qlvT2oEO63xelqN0QeFQ
3GgaaJ61D3V9F/utxdSE6UO9LOmLqVHkZMi2t64JOfiqgNT/J9S+vT+LN0KV0v1/Os6mFkU3HIRq
2ONgI1Pss4S4GCHl/HiQx6kBSFBGwjj3Nme85fBc0PmwE0E5MMhroSDgG7L3gEVlhF2M7H2ILh6v
udxZVrxVxE4BjSk20Sz9iH1gz477XlF2TW4809GR+Zv1dB0FmSgA4WL9z5WIWhp8/5gnUOqRTNbo
BAbzQUgDrHuUnckW7eFvFGXyX2eRiK+mUURT0/BSmOigZ6V+dnpuFs+G8cauWkr8L+rn/iAnNsmw
YqRl4zgQh8ttfLoS37jzW8PQCcFXEylbMRdH1ESUO1uwZlD2gznFLQ85YITP/7JXZ41o8WykhKC2
oJ5VLaAiIt1VvN5JNS2KcFj9uVVLy8FEqo4lUDS5bPLzCC9CiOGaYWtuznhn7HQvSXuBl37DVmAQ
eG/HHMRF01vRSB/1iHZB6MqidQ4NKTbjFwr9o+mx3xl24B5CWENU15FLhtKRT8aNNSPMDUh7tJhf
hZ5SsoXFDA2SlqAZEIGA4Uik/4h5S2Hwohc7Q6Ev5CMbNK9IFd00+3OaezXjPv0mzpQ9vYGfdQC4
TqOxycvlM6THqDUY6RrdWA9Bi26sqmXPUs2+LdEAT4XNGKfqMGOB4lemdLv2tnfLzyqx3Q6ads8P
wSXwS1o98o8zcnmcqN8CJLkFpvfxjjdY18LDT4EBuFpuClBejiwSxvdGvwIN+Aeyd2b1S5SNr/lk
kiaIw8Kn7bf5yzEuGWEIUTqnhPGyHzKnLNLj4Xl5JjjpPXINtVLfW9QQweRbzF/NVgUUgmKYj7RG
CLUmIEUeMgLKHXjIeA3cLuN6pgY/UDO9oRmJFd1HMWvcgR841OR8z3D22x0HXtvMiUQ8KNkUkLgj
SJKQKVVjSvgSbtuuuTGmoZjfSGefRjy1jKGbyKtCMQQnnQmoSfORGGzet7kDpB4HuJhB6G7aRDEZ
hxE+klqTfqfJjozv/4D8Tr+QVatsI5rCA0xAwhoqMT98O79a73WQwDeHRFFWIk0Uv2uSW/fE5FTp
KYwLNOPxvUxVDkO/f5mGjGUinUjlmZgTty3K2sYkSvShPe7suAB2yK3bufjpymeDu3QDjsCYzLKY
DhtLH7s7SyHbxCLOx8b//+M35w1Od6Ns59Kfb3acIkIS2vruyAO+U/9RV7s1GRPH0DcN40YNnuKs
IFlYkx50bDaQdKov1roSEh9Zmu379ybsnP6rcyaGai0e5H3ZdxjLwfUbajTZvZSP1L20D+mRkIRw
OoHvUykNEYbrIcsmk3qKDaAtYGd989cK9Kp677YxAlpbdBaKXaRMtiU5ao0en1b3jy+kHWq6SEfW
hNkKvkitOiz9FJUhHCT95ZcExFasZ/rm15ppwMABDvb23i7mrHkSHRNRX0THUJqBgNyvdFQ/rr7o
Hqm1vhNpU65VSI5y18VybYNx4nzu34+5ZlER7C/lM4nXVSvkRoWX3yK5nJiFLg8zahU+N1zqxO98
MfPW94iyMPg9tp+9HghKTMGpntTnsJmUMbaCsMntvAI1ReFYKaI1oAcyCSvQBqKkaO/oKTS8DIY9
MIISJCkEUBfLp/NRQD3kYN0BiwUGlgv1Wma3IFYbWqp4YxCEnwpQhbl0GThZWJpCqFu1mJUs4VX2
ojQt7Har+Wb6lfj2kugTQHJHpT0BfHUY38jlVe4mPq4gMx/HWROLtNb3Y4G9IfRZ6Y9i8+j+wN7s
L9pSTfh2kSNIQxUeL3c5CtbTuf7HhY+UPcyTuMg43OHmwEnbR8Tea82S1ceziZCvcayQuvXSNQL7
VhgZDo7MRIuYf4hg2HJkQt10PI7wmk3cTYwf506n4uuoN0ekC0yp/DZ6TIUDzpWysety2WDTCxW9
dSjDvMEx+d4+/hrLraq6T864LRdfXwC7lOPJdcWKuVNSXkR6vw9Xmv4rEG1c1HskwlqbfDnCf36A
nUdl2Shpvk/KdUNLKFSjaj5ghGXFiWNww5IhK3GPVdx6NQxmC2aJv4vEl7RVkN/wYp3ptDKbIDct
3S6TmkOzrHa5fF/oZHlTXvXThyASFGgJICJ067/35MeZk0ntcFNPwXw+l6anMqyoxhqneDw5nmrc
Kx68Q507F6X1DCDv0sWZJtjTxn7s1nTrishIZR0i/mY8sdFchk2kOYxAX9uuKckO2rcJySDoK5mU
HU2pq5HZsN9hGmf1xszSO73mmXZC7HJM0d2UAcqo8c9FI50SzQToWbWRHB+0NqyI+5osUS8vTuQW
RTjIxfgNZkT6CJ8XkexS5+LrlHkrYgGvSLmayZ7hYIsc8rQXOLebIPvlIc3Nu1VlSfssQS4Gx/OH
AwdMTM0bMQTsc+SqLgjknBugOvnPV9L50BbxQF+h1OR0mQwnn0i2IDXFP5gEgzoKzYaxsF1RWp7z
6qTMtJ/d3iKrw2PaYiEvUSGcldyLCx6L2EbtS2f9wkdV/BvMeKiMnfX8y9C11DZ8Wydi41F+qvT2
OM9g0XiFIOqhrbwD/esT8xs9dSZk/CKLBGEzT7W0qHwSa+Qijt3fpeiJxQ40dZs6+Fe2Tx+J22Ih
oJtWvNHEGivJoIT6xrx1dWH1WlqcjZFhU555xzhYXSxR7eWSZI8zstyy0Zompb4DWVa7LD9NvSox
H7L/q9WjapzhxoTv3pzCd/6RnxZ39QvLVlEVo6xDd/OfBg5oi9IzxvHuKtTsPYfRN2IbgyUWJt4Z
6iTXa7AYM5vE5wXGXBnGgRL5QudWRUrY572RC5enjK438vYOZ2hOLARU/ujAssfc7V+OeyWf2hKK
F6CsTqiuTMpyFoHh/E5n4SHJOH1imPRq9URKAByrs3RCo2m895LMX3OpmPMvNqlQ6Z3eUQy0ckxx
4fR32uTRsNiCbJ/zv+PmO+8BYATeKpPBkK1/eAd2Mv6F8UlBxkkr1AiO1tG0zgR4qjazYKHv8x1G
6Tv/jkYOsq/wJB8NGyIEZVIoZ5B+EAVdFiftYXWelKL3nZ/4GwT4VivOCBBA/B9P1fQIwQKgoAM8
KicUCZ0dwQTbDfLb4X/H4ldtK8JYh42tX8rCu6BlKeGCa0LfHcoZXlduplS0a/pXw8G1ogZriwn/
5Z6rC42IjGOE7l03oCkvdBeDDJRYn7/2FsBKk//b9nMpLd3n1sZtx+7UbLnpObjaOUAQjeL8gbLx
W1QX1zx5mKq+NHBTfRkn+SvgLlsJKf/i7SPe2pFmUsgXq/m+OcWfpvGiqIQ8ofbrq6B+bbkKNjsB
IsjBrxfe5y+g/51zhzLkI3QZppdoL7S6na+yKUj2uiqN8y/S1Q8oZSjvVp4QcTPyKyotlhEpuqU7
Lb99hu/Qz7T9lIyTWEBsNJM7uVk2nVmjrIZ53/0FGK3Mi2W9cfU7pea7lGbEKpr5m2tV3t9gzlI6
5EvjmWG6xwalDLWTpvWcoODu8w8eckrMJZfHjYyyMcshChWl9GXQ5v0+jxktnCaa7V1BAb/t9mtV
QdECj2+ZJrt/n8VN6Skxy8NozFfOMZHwWqFfkTODRWv8wACvis2wB2l9mIMs2/2zdAncD43BxZZw
UM+MG1LuLfmNe6CdPXfO/IqSk8oin3joakLgUsf7cjU3YsQThWrhqwIJiHNMS1ziDGsCnQ92IvX3
uod9hhisMvNHPMAECMn++Hu3C1LgFgvXR+V2OE9VWNWVyOvnAgRUfPyeSoWA5xk8CGc6fNOaNPV+
I1aM17zi5q3IrjVyVZmtmPfnaRY1KHb4xcsWoVfutfUqHBAr5Kc9hl+1MDQBGSogfcudTDMqvW7M
7HtSS6HfI44bVki+dwFhb5kfJoNLvbO17QbdI9BwtdnNtmuPcfbFdzYsWj+n9pop82M9YJTH7s3s
RxEbIKKCNTI7hMsILYSD/Bl5OsZ2cRJ1Y8cc7z8BEkJeVslvTaTM2y1NHsqDQ5Bhondb9pkXw2bg
ZmUhPlYnK2zd/QcYMD9y3hTBqSwmG4SJ+5Zr/FIl89YpdW2a9mmyCBl/Fg8M908nyQ3UL5XcsJFk
mP4bysKG5FKg88brWbj0Rp7MfKKswjmq+oIJ7UbW1IQMRTGLdj+ERPZI+TK7Tdj1pciVjbyMJRvm
GhWpJtpWoWzI7f7h57RCojbTw/gl52HDCu3wNliQlUCzSWyWLfuCnEJ3iSKMVakZzYMhixQCwMA2
ToFejxfosLWNR/NlDN3lTojH/Sgw1JWGDIgO8uUuBVReMqEEBWYTQQuk7utlX8QUY7fS/OzT1m2g
PYTsOz6xUcVIrrZSsMSF/uwYl3vKa0fF06LDuU45RZuVl364NoFdGc41ThcoY1Lauo87QP73TOTT
bxx3rlyZZG0pxH+uiYAcSDoIF6jdkrwuVezGGrwKegjwDpzTLbdj/H0NxI4JOdqVG0CCbBA5iX+2
AdF8NasKdg1C53/brIeqRWoUyHIZXg8N8x/d0kszZ9halC/bh3gyPrvQ3nO+XiF6Qm9MQ8dwvCUA
4ufQvmAOgYh7entZx7Xn1DorNz0gD0o81SEOoPYyqvUg6TFIN9ijT6dcDETtF8aBA+JV+VV5YDIO
QbvPx7SIMHWgtcSUzpm5x66lVYZW/Lm/HJR7V1pNn2NZEYQEWRWxcwvP7b9g5U7hGDTX9EEjBM7q
Gl9B4KCbntvKhcoyPZjSVPXcERySxuid8yTTfERG4DifVNgY86cDB5T1UXsXhmybuzFD7noBzubn
oxTXUjP44YkyhePazv+Ns4JUyPSBhVK3MX8+IJQAgCnJSWOIriFnw+fwS9D719AUm7TvrE5488xc
u0fgXUMHacQy6dsVFNvxVQmKlyjIChM8XdQ5Y6EaPdjG4XYrHRrFw2zMRHhdu/X0dEA4R0KOWFVZ
rnEnYAsQkiKGB7oxH0T/WDsze4q3cnxj3vRfAm5PBG9KVvR5R21vjRsqJsHUENVKrTSJN9O3Ozs9
wWGXQGZfZd1sbN36xlLH7hNmfupX2vTnux4q93Kz28d1uoUhzRAYVF6Q8KKmmX8iIrwhMSHegQjO
vVcLd+bwc9HBn9Ksrr9h2zbaYjiPRF7pEpceknKEhhYYy6H0vcM96nCNWi2VsQXij+kL82UoQJmW
gzkUeipyhXlWpy0a3uF4qSLeuL/yjVOTyUBYvkW5y9+UnMqwQZ6+1M6HfQrSJ/M/uGDcR8AwfBD5
SS4opgRr/vMLYQ0Gt8NoqpqGvM7SoOdl4H8V/FOka/vEDARUr6T5q1VmJrn//vIjkS/l31xu7L5q
N+Br5UAP0lSsqDo7/dA9L5hmFgL4g8EySPyc/gGM1bGszjzlOIDGpE80PDFsts6rN0XZN/QOjP3D
UC4fIyhV/EFqxbio6GkKab2i9wZpyA8GX/o8TOzxriaW3wn/z4fMxRJKg0eIEtNU3HIslp1HYaIy
XxAc0kQfP+JTfg8n4CJItQA7opxr7FXV9oTlO8IbIEmVMuLpHAQRAQb4k0jKIzT2zIZIYFSbcU7Y
To+3cYzXpzhF0/b6/zHI04O6RbHXanMkGY3h9QCV1RlRyE2vupMNdXl47r85KK2/p6mi5cXF4Ut4
6iOgBwC4ugCKzFJxQAkktuhAw0X+Nphr3PysWzrQlEF+vxTlSRuVAfzMh2H25Un8UtKQI7IGus8q
TuQ4PfJmiMp66JpG7Uy+rcVvjS+Y7VxHlI76Ljin6HMKdS4FumTJSapqG9RzLeu5CNOVubmoSSx8
fIltUIqI7aLIjrp/XJNtoTAno5BmiWpM1WSIleCb2Syhf7Ru4KfEPRF82cD4y91JjKnzJHWlNbS2
wHGA8MrQm00vAkhdBWy9AAk966kzS/2pPM8B3rl1CzKrtA8j4fS5WupvbxOX4t9jO+RXHS4+Ubvm
mVs1oJtngHsWGLDBgbb1cCo8Px5ofs5CrPxOB3/h5rMF9XkQvIKzsMTqHde7l2Aa80vxD/qZ2Lii
T6+dF5g62CTWKAKPx6m7ZiF+J5ZjdOLL97/X1M0PH6ftrqF0+24C7zzpz96IrihG+xLIl8uouh0F
pgZVolCjD3BYLbbOlw5mf0IebkOEEVkHfAy4ZECiMJF3URqxM3mKUgL/ITf6omgOydK5deksqL7P
cbwxCr4e9lsML+MKYnjNiBqeXwmBh30i2JEMVP0OJBrgzFNnECyAKqeuL5vrdR5laTNn6wz4hiUS
cJTDQMAd79PC0zArVbsjAlJunOBlSvrtS7LDdmeB+xVog6Q14yzrvZNawUhAVLNuEnGB/6Qrj5KZ
w8CmS7XoGFb5z+OvpyP1SeLBgbE3n2nRNRJsXxPUByrAG6WpBrjj47COiEqw5DMy7fo9S40gJeK9
y10iGM4KPKTJd+Pru/xREYKMs3z6Ydxfvjn2cC/4oRFJlZKntdrSFyeVX+Xbk6+CI3O7c8M4J1a5
REV6OZhOge+ShqamN66H8DrVLbToZcUZIOZb9KagLkchsYwi6opopSIfoio7LzBdeHXQl1nkXT8c
MSPzdwaiqyvuIAMin1EcywCkwZLOYjfNGTvEzNZgSu5Xi/A8XOS481K0z7LbTGOIZzgdCGdixJf8
LBmt6YmY0zSg9lOwe0qTifTPGYyS0Wp98yoUUDWejZZGf9BHMaUxcGCtyexBes2vylFW3+vBEdIV
VAJuqu2nWN1/0nLDqNQg73AOq7RuAXMNEXvVam+LcP5N0mG6h9rm0G8DfHNFBbjx1LQ2hiNBRL5F
YHv4OM8OzAKVutCejUPkdDkzhNh9T6jdRytP+SA3Ll+/1/rwF+M0+5q1Mxc/oi9t02hGxH2YepJW
5eQhzLHbr03uPHOx/eMr8FiNtiefT+BsypzDGfuDxuIg6wEig+z5fKGgYvh6OthQxmMAwZyDKbA8
E2t404grIV4y5fJ4O4gJMc9JrUYZwCmatbBaa9vVh7xfwMVa7YoMmPqo+g5o3j92rp4HLKaRfW6F
zx4qsjnmz4LhkuqSrLRYzh39HFymxzEypmoL8i4jwNGBmKmDuKj7Dw8NPvSxIA1rGK5DheotLXMX
kaYO3vGks/ZjZTLQVJsCtEJMLYPd9cyV6KIVcCYc40thDk373S06gIdPi3KND1XTb9rwuYuwbtZB
ThY4OoQYZ4tGKzMzQDNC/xoCEkW4nLq+u4XoWSuaJV6Mbl+chZh5Euewev8TGAgX5jsxuIG9qTT4
Koi6lv539ugjhQjOFE1DYjRjrHot9EkbyMU/2TsSpB/tRjln1mpN/amqcAAe6/o3seJZS5OYRe6D
a3s7nyJyVr6bNxlO2eunI+6LxaE6CqoOC3gZgSUBDUw6h9Tig5WrpD95B5SyBmtffksnbE8J48Do
iPEF8nb6aGgnam8qDrSXHpA+a6ppwI4thlvQ2fSlk9+XHGIL0TxKedRtov1DQeuwEjjJcFFjcWzJ
zykYnz0HTU4p3k54wgS6WezCoSAm/edKCTocnLh+igeYOQlmN/lZiT6A7AuOXbiE68TH3KPMJGyC
uMnanDBpsAIdDAsbGWWGum313p9KSWOrQQDo+scEa1vSqpj+AvfgB2M0Q9wt34G9fedRRsOs8Wvw
GRhbco7zb0C48Cwdzydr/e+Tk+5MrhlueY40uHJHjCFdd7ZcxI6/j27ciupAIB2+tVHmX24xhhqj
BmdfarHDTz+f7l/mGQsT1qthz27fu3FvdvoLdqnKFbb3OyNLbkCzKjFvn7KGJ5SWbbSQbwHjwHDd
+RrO5PZMfReq2TjCM+Uw6wliUlXFyICFUkIf5fMKqmbS1/3Q+N0aB53TOdKU0rjPVOUNl75VWG8l
m8iUGBMxFrxSHNVFfKvJFeuFM0FPk9TY3A5jhbjSCseFM9FZrQJWT1naLSinQhBvxH/Zn5VQWnv+
8CK7/tGJm1DjnSpZg77e9/LvmwOpWTQo6ZgjDp6Oeb6U670Z838m3yCBv/oVx66bYrJX422aBrEw
P2LlyIsV7+I6lCHNt0/PqbH+JhJja8laEB0WMkwoPBeTv30fP6zh8RUEReK00nGgBeMv2G2Y7gb8
mV+sO0PCcU0Bxs7nMIPIUVa2g5UKhwz+vuJywEFX5HDywqD9LDxSInHULsbpl1YSO5M00bEhLrmu
gQtqOJna0FHS7eQWX3cymSYXgfCcoAZucuD4naQoaCX+HfA8NJMmBLcyCyZGxyfNH5Y43P/9z0RE
pyStMX/jqW5L20Y3dIWqjkah9RWJFnU0xzqCe9hJwlxzOimAV9uGYtJNXbnNDVHVim+njMSjR5uQ
bX4MTfO2o9ftaxXu7wcNqvGRYI4sCj9TAJyxwD1Cr7QzH0SO1NWCzEAFvzyQ2SUxLdQ23f8O5z9h
3oAdfpxdCFDmkYl4CT1i6Uc2F9aMu7F7m/264Ld3D/8Ye+tbkPOuqI8uMAO1ySGGYe5VDfwk9GW9
dRZNnW7mfXHhRkU1bc+jzHH6BssNmStqTcO1UHTXTWeJw8cSzlmFYbaEjs8OTEQHyYMOU3ko2dFk
zRvI9SgMecvBDIufPGrlN3MK7RuzxLItHvjTPgAue48cFLFkiYQ0Ny4SVEGHldxiurh1CnwAuxEB
vFlLpN9ixJqMfi5G2YkcJX2tURH9JJBs8zjamiZ7Fbg/sMGx+CnspWXOt+r7KGSP0lOc/crmxrFF
wzoQf+LeSjvshy+wmpjIn4E40lOyzoW3u0j3AGh0dQoTrHeELwxVnwMOJ4APKwjqFlbbSpyzr7bM
mb1G2cICdTd39V13dwSvU6JsBvEgRliWzjZX0c1w2u2Opy4vUSN2Tjvmh/0blWcQCP9lbSWUsvSR
9vdlaz37x6lQWGUMpLzJOEUEegVLJpewkIuqE+L5EEs65Wd9yufwkzv6wleuFo7zZ2Xzn7yw1oUn
lvqLnLjiPRyUvAFT9XpFS3TQqxbLAIF9ydDZBVyLQbMcPELc1ihmK23Hjaf+w2L/MLup3z5NPbQn
8xz9SMoawSp92rM9N30PnQDS9bKt464mrVOtQlXCNEz6GJS6omkhgjlpCF5BytxQQxjDL5vbx4Db
/1pLvqejWz0EFsWZumfVDg1+sBjznoPL6qeue1XSyb1YmfzDB9cVv7gQGBTMonnSUhyivJpMOdp2
WAEbhGzUPt3xhmrNxePTrQ0mWnztIFOJn1gRucFjSQjCubiW87tykPa+9I8oHR0GW4uk/RoRma/t
LF51oEdwQBCDOq8nUnDylNFrTl+4UJUFalpqGwEKUa+G7rSeIXxp8ofya1dzdiggaEQmfCMQfETV
KP/DW2WB5R3PRZ5rdsaO1Va0FwIvRinhchsRv9QrHzbGdrlM6oUdbYUggoSgoobaG+eIqAU9Thlu
GYUdfeYLDkyU2+7EBP6GUm+rvLaA63JkqF8eNgfygna0LU76kXWvyBStCTZr6ZFDVsEOTpClE9ry
uvNERA4YLnEuQgs26b9VnS/Q8q9OuO/jLZXmIOV3A9qpds1SZLdusFW4ywDij1FD4Qrr54R9J+kG
k1NYgJv0Sn+UXCW55erTtNn5D1NnxJfE+I1huxgGV5oEHaHMoZd83T3Ie251K37HT1aJTxGGtMlU
rWnwvDlN50HKAefVbHJHOD74iuQDrRRMW1vUIYNQh8R2kGUgMW5yL7YPWjPoGxpPLAWl4txeS0nz
DhPPCmDBdFDhXmUeflNYlOPTuWJbz8O6LiDstV/eJXiKAJDmdQ0xqoTagm1cFxYjf6BJSLY9sGNM
FhDUNcUUdcrsnInbfcN142wUe/HdE1kv/bLKaKGcuigaPomsMlPRkU3MUNs8ikU1Vp/lWagdDG+H
dGMVzciw3LFidVRh39FO4HKygKF3yqI7/TbMKy805UGI8bkJvPXzvOJ6+6HxQ7v3XCL+vmDJcEdh
crYmXT89wHhNpkxEwfDcaBvyWbztizCvcSYJtvW1YRywbH+/5TZ7mrMrb5+fGOhQ+uiIbklMwY6Z
B94/BGtLhEYR5siXYOXwp1paMJ3Zi146xfW7wK4KkC6VBmRYb8dKFl6SE/Z4ByT5edVdNErViKvd
H9OirOghc77bAgzum6iBv3CAI8ihqvJuA0rFYUT0T3M553xIC889zZmWQL0gBCuS/ukdp1HgWqMn
1uI4xMjgnEO5ovvG1FM+c2zWMIhmLRRN3vEREsHHPuu85ogBt63y6CzexgViD1mb0NJLpZ4gVDNt
X1Aky0JuOfIGdAorNXqzwsjdXPC+FrzAdvsSpdgplfMpY/gcUyqxD73cnDWkBWPI1PdlbmbEr+n8
nmulcu+sjnC1Wljz8MqAtUxP9CMSI3WWEbYBPyqV39Z2LPH3+IkWnefmNwd9+N7GRbxCEHu+Rq/X
hwbxi6TQox9hcZPYK1yBZL/g3u+7CIVCS5LLLZ29goRw81/b13Ft0/nq8fTK+uxETueWaVYRp5rG
Gefk3SKipbUXYvA8s6GJ+vw0gjjdGHzC+ipsGvcbcIhhDD6/JzzeRv9YxAfg2ELcIZ5XShe5f2Je
08J7F7aNMWcgyQG7cp8z35uCQW9YrFz2KbZtVl17xyGjoM3aAS5S+LaSd9kk+EcM6ShfiKQLSq88
phXIkspuswrWlh0R7pJvet5MPnyHT9ClVbnyTXVzWOu3SC8DTZJ/95DVxsnUfYXL/xqQ0XAQqkzD
yWfWPF237UyUssFKIlfrVDmyaGCD62h7GekkfiJNzG0ZZ6XC4RZVGUB6MViNtfBfBpGJpUZsrPEN
dmZ48GkcI7P9vXcYVGAsyULNNiZj9RvCgp0rd1DFzbYY8MXM5Z0OAGSbWhzWm1UnvdjR6Y35mGwU
T/Y+h2tusXLsY/rC/RNgKxNbHAY8nyca5JWgl7/ViUEE1VSbnrTlStpDZE4qaRmsDJdDTi64Axfq
oCWcBxV418FdxFfFl0cYZ3AgllAPYzu5o4wJEfP/EiypWbayk29M347g0KwxbEEhAyXuFzV7paab
ywzWoIHMYyJ+peKN+aKW4JchS9VIu6Z3lk05mHnFuCRe1Cdhm0NXdC1NCzxbIAR45ozAIMhGbeRs
vWlhwakGpDNpBnmsfG9L4SxGb2Z1dR82bb7URgnmTWE3YdNp00nhkSy6qSQ6U1lIHkH7v758gY5q
vqYI6TGMT98KgDgasvhL/pTWV1Dlw1WcnXDYGiODxYzn2valiu8etkR6ym+OLm+Sj4MPK4o7ao7w
em+fXUa3WIMuhs1FJ4RapJhqVWLymqgq1VXo7UtmtV05n894IMgdDq/YzxA50JtQbfAs5iMI+Q1J
ho4U0j4BQvk305Ap2ip3QOqhdVug+s12Fb2liOdHHYacYedZmTRUTNaVH2KxmWtLuYrNSzoKa1kF
dzjo7a4WVOGs/W4d+KvfismIZuLPkevIJhl3PPHqLddnPbUHAhZzicOpYqlHJYwrgbDxhY0Vb+vF
ybO0tABk0SpH7RTEjVwCjmnycqqPo5Ltbu2J7NtU8DPxMInLDeza9lU360vpwM64NyCxTp/zJBlj
FE0StAtM31Cq9ThfmWrZM0hAe5tdj3z2tjxotaYhAMXTffMQLuvljRY6wAYUgDPyh7MjMK17/nck
C0oKD8HdIpROtm3aXU114wETTSQ/ZMP7ABUu0Hnp2EV4j4YYUWVzIoRRAtCDZfTC6y7uVum05bcB
klYk7CA8ryga7Q3rJVx1FV99xAuLWzYYFhQDcQslD0S4x1kzc3Jh/VvHcHqXXiCviBxTcRGk9MXR
/y/MIhBpwzhE5X7tqxsG1y1uMLjOIPFvlTKe59/uSyhII7qUY+npNuA7tle+znlF15TXGQUsQ9Km
QXUau5ynvq4URW9NjzctrvjUz9e/QhUhh8A8PO9r8uO6WpMNpEe1ADk7taLNaGDhx6LrqohXPSKd
ccYttjzH6LB95vCpRWHoCE75Mxm5rZBzVkL0dsMOfEBVxXKUCuoXs2NVY5+gkDR+ugd+e5mKpSlu
P+O6VLvAMtMPp7GjG+6Y2UUv/uh41e02bGqJaz43mleWS7H/8FU6YXiph9wi3AABeECnRY1nsoSB
YZbsLTvGl17YsyGN4VqGEOcHHELURlNUZHYxNe3Pi8wvHIIuhV9S/0qA1wNmeilZKDzw1rNQPdyI
awAvo+7d1B54gSFml/DjLLGk4+nj3EFpXAzCYGg9CohRVs9t2LSyBcRq02GZZ6/Pvd3n29+4B/l2
yNpi1lIqropkIWUKa7rox+53/nhADjSighHdWdPuQ05OjItUdbvYYTmxIZt0nEmn+eGznCG8x2Cy
6eP/if9OpvLx5X9e54XbhRIrMzylqwuTdWEXXvxvMN2KGkna8w8k+W5XCnFOTDT7WNalkQdeTm6b
XccVhhmuh9Y7pNm6OnlfsS6BIgOMsFdjENZ+AavctMGY6+jJaKtaFHe+K5bn18C8GnwZXh1H6v0D
2hxEap2HCAAZt2H2anxZN6rUgdnRMG9abmIEGPajfYXu1Izmmbs0lrolD04vMlqvAeFmbDYQWJGh
eYcv4Ii/KFIveJ2ZgLf0tQeLK77TkX0/aV6uUrnV52cRzSaEIYrUEZSuYJ25C+TXYBiDTIoup0IA
j6B0Uablo7yAuYiligM1WIYNUJ9bn69I1Y0pcQDRlzgV3Ry3PIoWxpEBGmIsWwUqyLnWuKzr78pT
KKa5dZUbUua0R3vPIpbEZmnDIUP+OQCf0IPii0iQTiqfw9ITmnqr+DlrOXyGyZoHH4PtgZnAHXWr
ETvO4ZnxcNla4oAUk3Mp+SYH6nzsO+B+Xw81MBR+NukXAofizbd/4LbjhB6fQjbYg376mfcG4pOV
TbNQ50Y5UN3UAv+7OGtZHXtHf7e1q6Z8vADx5tRPGsd1MFSVOn6oyox5nbBauS+frabz5yoyq43c
2jagwEk4tNtc0pLOIqLCHu0ZhFR8uLO8F0Ye2krswEVdWJ6UR/ywzovDAOEkxGTcHY9FKUx/5L3/
xF5/wsIZJogBraCVsVOPSDyy8/sMl37zuGqoaQrMKDmne3FIq00YreR8djrx+Un+NjoCA9jsPtxF
p57jvWs7x5mFZUhcoe3bJr/K85epPckYTzbCWnkKlv2gAIcgVj6aXj+Rw8QncKheU7BOpvcnu0ve
1ZwgqdotnLoEFJGP+jvnKi+KsRah3fNCdF8xhXDBaRHJR7j2Z6tEi224lz7dvWxyEdcUZCL5r7DX
mVQqq6/uGbckQafhitSwW0ieKMjZaixTimFZ/3K0kKiSz6lo7C56mK1kvfWyv9NVObLsN7cK0Mnx
yieJ1P8kghUPRtA5+nIytRLEBe27HMpHI7IwukJ9Yd3s/DyKG894rU/HycVZVMhyhuXN98zgBaIh
4DEr57NT0xsjrY3DA5sxuyn9XGrqrE49xg/+BInFf2q2mRoxNNLvjr9Ia8iJK/Gk+BXLxKFbBlpW
O9I1D0Taaptxrb1NW59z/UScCXPm9HEPlDuartBV6nYpra6eerV1nWU02Bx6mrVVZOrMLQZPy2by
jfAB9EDtOIDKTyg2sjNTzkn8qwUJX/1z0HQbL1d5ZqrDljqp87c9cDm+5SVAE+U7g0FyvU7/7RMi
ZC9Me8PKmYQLaa+99Re75kKgS7zJzpZ1VHGBmBApPIzVumsXs0TBntqgMSZ5+5xP0chxb1Aye/6z
Wyoq+gXgQ2pxRaFFJ7fAW9gnUCmkx8pqBiWQlDSX+SoJlEIX2uL1zJYFF06kAB7dKICltM8fRdJS
9TwXqBPy0nZAUYGB/Ykk5OVx/1iCnfSHXaMa30cSm7vlLieDnaxSpJg4XFJNoPqPDpbQ0tT0J9NC
uQwcM+VGYca6LsYUwFmnR+Ylp4ZfXxpZm7HP1AvzTeUaChvlCdebahsGhPrXxUY8hTQhqjg87ie4
mgy5H5/NnmtdDZarpJOayOMIbLcQQEzctBI/D4xv+iRBdBOfzRsq+bJ+3mOchRvRCXkiP0y4yyJL
C6G66sRKOrxpjD4wnGDahvoE7sRxOMcLaYNHFKXmNMiE39m25SFuAcybu0Khol2p7cB3dsXqjvkw
pJTbKrtgF2xQHrmdkS6jG/dqWqN1V/KfznSWHTlyEiq5ELVI91TTDYIdG0uAmK1wbBkpErVyVwDA
pM/K4Skj0Q+af4MtMCP4bF9DQpPE+Nnc53iQQjJRYPs2ym7bETGPz2EqQvDvSJzk4g7LR0E3zJlC
rUFjLKFVhCalMKHLNrlbgnSJ1kWuwbLU61omItbQmnOVj+fl8No9nDvoES2CitBiIs8keselzRIc
AHXjXn9B/852vcOS8+Cv6MJXl7jk0SBPvzwHWLOgnCjiLaPU81DDZ9Tezx5OvyefViE0xhMe9rwq
l26ZCKpGwMHkMd2u/citDSmknIhFVDvdIdDvoQ1NIm40CwGrK9sV8RscWU1hD/vzUVzJl8REbsL9
eEb8lZzhkQ4faVU3YUsA2QC60PenY/d2wv8kQ4FURnzACBc/izPysSgCcvsc+qAIJPYosHK4UOJ9
74p7eCuEJ4ggRoMb+Q4vbCW9XXr/T0i25n7TKsdRo4wbWyJ9pLkfDBdVVJixyKeZcxevHZfDhYtU
0cpWd2UvuTWSPQLt5usUTdLm92YW4Y+tR3AhCdnYdlH1nM+DzokOTC5KcDudvKvCN7VPpSwxyl2o
EVKAX26tE7gDQFVW/9sr07bUpL4LOdc6yLUvab9Yyv9l6RqE5eIg84PBc92u4p8NA7bUp/3yZoln
0DIbYbSmlLzdVH752hv8ij7A052ojuyV82rp9cdAurj8CvabroGNWxRfzWxs+VPAnbNx2Gb8s1ur
sPvqVCT9MzkLrA6/J9BR1VxWllIDfpFQRlOeGucTHbUzx7fboSOjhaEPGeK49E6ryDz3v5RVxDqn
QqD2N2w/dm5Wmg7Pe32qYWCgsqi8z04f5s2MF70VhRZcS32aBM/BFLYAyA/YMgNrNZ3N3GCB/xtk
kTBe9qQYaiI8JyPSohgfeW8eT4LtOKzSKXQm+N4kNPus5FLskzrkAcpA2Q+1y7gIR15vbHrNxzKh
2TcOyUIfFNehJJ0F3Hc551Kw7llsMUODoBEPjytkSt0Ac60dXVlw3FQjJve3D7ILwTyGkB7qk+7R
t73uWeUJFkcQb3ZztngjUXrmd8BXb2fK0HUIgB0RaN5sCviYtW+HIx82lwEW/Kf+VL8inatl3t84
CaJpf9mduZ5oTAmYvMqBE6v1J+bELX0k2KwsfZ+mQPPS4o2v5EbDM4oIG0Jim2gb9EtAKd1OwEhI
aLyG78Jzu5O/G+xhsDkdZ1xkX7ej+GTSdFwcLqOKJCxOhLNn6Rz++8xgffaIy12xUiL+tTHxjC4F
PC0wt1/vg0MgJKHJ2CDRCVQljhVz/bft2SHcYdAiw2P7Yl5a/ohxr8fJn7iNod+mvs4yHWAE5C/d
sp7kndyqeYF/nQ69mZ8H80A/93Mxpy0e1tr2LFFhqdVAFCQRpfKAy80qWscE/eP600KVpbL/HeGd
EWtkMfK5Em7Y426Zyo6gQpOjgKRlZTbt0lW9v5OQ3GRizJa0GnJV85QZoiyI5T/OyS7O2PBZFuIo
TJeY7RUtUrgCue2FWAgR7+INYPluSp/HBxIhN/gPeoBCKdBwLMo6uPYJM4oWU6szs6SHxryIOoCn
X/Gt6pgrSIFZ2ZlukvP3X+QBHYm0dukmpIEaciWZGm/7xBXjSnANepZsHMX79d6tjbsKKNp+w4XU
6jJfZocQ2XZKVoK6vPq4JXzV3ho8Kd5bBtuQAUgAbeDMq9CMyY/H/6fI9QCmzZgBkEmXjqHX3BOI
CXPVIoLsWHp8YYobTIrUteeZeVLAXej2pYIyeOqRQWkjhRXqUj2vnUIxIqx77+E+BX+BlggA6nAP
VT7jIS/sISOjjbz1NkZL5A/4fIgjORYRsTQJnYi0h5WZmR0kcQz6fZyHrsrT9VH1Bu5XEYrQ4TxH
cJx73tQgcS2eZkn4Ltq4RB2uECv4NST3iXIDybyy9rIf0kdaogVyPk7coFzXTYql4qg75t6GuMEf
fi8yCzUsDZFo2pOixLJmP5Fg58xFZgGVbQ6nkzX7ZhvZnC1+Hy3p8U9Kbud3qCPb8xINDXBsFj2N
YNtgXkp2ODiybdkYoFxk6MbLu0kYLy3D92POqpKXv9QBZgVQjnJ+nN1u4pEY136x7D9Kgj9XEyC2
f6wsAhIwLdq80vFhY9DZ98mlqygb2dCpFEs9sLrQzM9gLXE/2ZnfiLSC/BQyee0YDhZA9CHtDL9d
l5uTa13IQO0ySuz7OpJxFgxVmNfbNClbCbui6DOx9Z4i5iJooP1vTUJWTIU6L987ZZE5MDU2HL1Q
sIRblVKypMD1BR8JFBLCy/z8ywVPxdXd0wMTOQx1Car5aOz3iCKoZxPKuvuMPthMw7wtTIUPfQEQ
0TaHaJaxFKAqRXgNdlBSzAXvNDU81Din4wOV4IqrKVX0zS3sKxbOf87+figKBfSxDOh6XIrQLM+p
lfB0OovSop426e7MIlPy2qNi5RiUslHVrtjPjezpm+EkAOKJPpKkPbuZ2RDLQZTSC4xbnhuawgVq
Xx8De2BLEkqKCSExqaxqWOfK/xJs2bL8GBIAhlp4UahWdd+qzAzMLPSaySX0O2Aho+2XkoPtrbyd
YEAUlQ2YICEkk9ed7JgwW5JzO4XKva2J+yZZ06yr6CFLtOptxsS3YvxtMJIStnVLqO+oMYupgWYm
Kmk/6xwLAJ/zmpLbrJR3cK9uKFvm6TnwCMwH5eQ6XLtwKTYbjnHSPEXTaBR3vkbJ+Qm0g9RtIfhy
LeVGhItLvzAt3LDbW6Sw8ZUsJ4il9pWcUtr1lRTpOshKFKu+pDLkCrEUyqiUgy3GZuQ4IxmtF4Nn
gmSe/NJ9B5Yd6Z1BkakMBrkt+4Vxt415bycKqe6C3yi6TJDjJ+kvv0aJqx116B+t7jPQgCN+P0Yi
Wtfsm8UWtqL9W0GTSRNFfJ3J7LhncVGtMSRXyQSdeN2bQWNOFVP3g1l5u7SM9A0neoLeIBHJsqmU
YmOKKxqN4/7ir0tWReoOO6Qm4mzg+zuKFS+jRzm8FowiracSaj21payIHpqALF7xtDaV8bJ/Pjom
e2kxY61+A3kY7U5z0uj0DV2gjO9y0l/XvntJlQH/kR5Ykhd+bm1Ff57aAkPuZRKP9nJdLFSt9qH/
TJr6f2lI0/FCAIUraI5m5USBVQyVgfBmhK934mPEH439CKK84GZffyZ9FtYNO1jI70+xBWCxnx9s
deRF2/xdVdlfYSCrEGkRev+1/Nxj+wGi4KUwZZE3+um/F6jNZ6k/0CrGHfOoVt6igjqN90oK6ShV
kpMDCWVPGdxZGFQNZbGea4xxB52cIipWgvBKSMk9Iboriquv4HGMX1qNjleOU1nn5RCsSp953qvH
AiBFRiyXq35lTnsN5Tt6v8492m7ptH27ba6G+bFDEpSTyX10c0mO7xA2R2IIkjWkpQXnlhb/haaF
73j9Mss/RRO6vaQmHUKmkCU3FBnODOWyJ49OyTcZcya0hZeRrd26DB8ORURd64+jj0W8nGKiqA9f
MYu4X+yZnu7obEtYhNhZCzupKMTEavEmX26UoCUAN+pFhITFSYakGS7I34XB0idFs+HnoGjv/Dgj
cdiLJ9mp/fp2Xxdfh+0h6+xs9zT2gJHlYEkBW3lSuUH5Fsom0VHUTWnBgxv3ySxwZzC8IZXvGShv
N66q2T1F/qRNkGbOtaXPhmU2bqiHG+J4MoDX7YQZlxuC9dUbtEe6wZ550vuqQzFIUeRFWcg39J7+
IKzGvyxNDwtNcwMrSVS1Z7KKkzlTCqTJdxRXRGnjZUWo2blqEUuthaLtM3CYIZ1lQ1+v4MpkoX1s
iOTSdrC/GcQJZRpNvBhKvnEL2McZCOLqkE3cr2Zht6dBMYyj/a8oAs2jrQuQz1sP7vzQcINsZFdM
DUft2XrIKbv3CO9f0shpkxhnCYY6Cqzl10gaYZubFOkG5ujCW9DdnpRFjK8E9U4WuABytF/J7edl
84i34AJIXaAbxXjyy4OTopiqP8t2p7riT+7iMSuDLGifdO6m4u6cnp7QtHJKkUX+5z8Y96hoPn8u
BN2bjFRe52RSAjNLo85elFxa7hsfYW8m8Hm2W3ogZxCSNVorbZUX6AGFbkXnyrWiIuHqZxaaawcG
QMomtGKTRWiM9JWKK+oAFS07T1rEuR2xFLYZJXIyiIMaEpkigtFcXSMFnvHeODCk3Tupm1iT1tuy
jftfw8WBHC7hMDiuXVDyAz94GscAxlgd7kUYtt9g+J45C55XcQfw4n1nes8HetkIxrC8bDN8JIRP
jtP8MGCY6EpPZxBP1W8GVaA96weTuBcnlsQoTa7S8dLcYc3Wf53xsWV7FY7AZpAVrhVE1j/I9kAi
JvkJjbaIu8uLwf8W+mbeyLMKc0BYyJYr2hqDz/GxbTNsbk3kJmeOMGWGR5/HrTSs512vbRYVn2ZS
Fua3W9mhojUwF7exTBAGNOZ63gl/omgeA2FTZjNONoULWrSHz7YsiJaqlBAzGEJ5ULdsNsJOCOvk
WXAGvYgKYPT5pEbMhnXqKqP7/XBwmnQeqm+cGe1+YBU5oSDsseIn+dsxLJVAlGMSO8q5WICQZb4S
4NWcxbfBPp7B9ddJ0ePA1h7ed5rWZ3647/SYZevuBKdYd1OqG8g40LVdejVtAx2/Che+3uioQG7d
7Y5GZZyPBWMXP1/BvHoKhsOb2F0crkm40SlVj0cyjdGoLTLtHo02XKTK3yIz8GVCwFQCu+4JovP4
tSxvThCZEeY0mEgIdKFhTOUcI7qjPhGNoSaWzFxju1HTmjJAgclrsR3BD8z4TS67yo4xPoCFwjdR
djO9uEoLtTwgwYz6PUZmSKMc3Gj9PSCLsVPhuzvAe9tbHcqKj5sSQ4KCOVg1BSLGVIUKDqlNo1cB
KK0X+iSugSb+1Y/HjsRrQGXyWj03ONEEVZil7rObr/fjivVStQwzcnYQgAPtIqprVgdYmI5k0TfD
/YtHlRL4fYACtoa+0YrLHRvVeG0rZ1oWII4fS9TBGzrhWvXq0Yvtw3hKv4u+tjjyPrPh4DOEiyGr
WEdWIP2UcDyszaGiZHSxY4uS5bz9PmCTq6LEZ64w+5a/emV+nrrCpuumCT+mPtSzhxhctraOIPNJ
bOXFN5o4NfLPOsHSYPjz+dznlIDGsQfv6P7hrItojq4ECaOzLZD9WIy5avij+CAgrHwrYcbPTxfl
wBpNnLHlaMsseydm46gtcL2UUo6p+7xOZ59NMQ2hgF9ZO0RxNTrU6GdKWkrMFl3Q0fcCUomgpGnU
dGl2xNDdzF4Ipxw7vH/EDRSFBU1SZhWhWhezJ8WFr4tsdE2s+pg+ScaKn7OAFXIM/ddM46f46oyl
EXC/65vSeF9d5BvQPSgiyZMXUOkQHExGyODF5AaA61jrUKIlYOLh2nAnFmUq5oSyUr7Wg5GiOXgc
AXPfDD+e7AKaJrgQqL0zue2HRhKgh2GZ02UThKhDsAVSKRlnqbLgrGy/mCXWUhlhVSD6V8KEJDeJ
PCmKOjJKjgu+/I1sMLw0VqEHUZW8o7K1GtEVbwRQ/rnYLBo5h9KT8fdOXPmIHR/TYIxSPwNZvtjn
EeO+JDY1QniR1T7u8/9884fjHe3hiTABWrEx3UqO2k5uOMkZD1PgWuCvPElv7GbTHsTmpEeDL/pI
Z6yU94CEJ2UbtfOoDS6yYAjUTrCHSqHEtRkN9wOovbUHZm/Nf/yDZlItOoOzx3Nrg8z9ZH8Ji/X/
d55toSg/o2vymweiqWWRgQwBYPt0plbT2BqEicOqKSZbVRTbMV6e1gIRPMJtfRIPrBwTDg0nICGz
p5nXuddeGXGfTSl0dTXh5eGIUwOCf9bt16JxifTSWeWU3CLmpofdRLOH0tiLhcd4Bywbx9f1HoCA
COqcCISVbhGet+cAgTHgkL/3ha0rWoycp8n50diY+K5k7y/rBTChOa1mRgF0yOOtlpEcc6ZWgI8m
V3kCNuzGxJbr9mRxfbKxp/rjJWJYj7/Qrbvt+ppX1PkG1ym6ieGl0U9IqLzNj9PeBkmVfImVqU0s
1TuWhMxqBG3M5QW6OPqJDcfq3eWSHTJ8nG0jjIF57aceCxhpCfnepj19PBYBXZ75vlnCU1x1Yq8C
Vw+baQ1BX9Qk5EiFS7+I+5Q4GSXhgUPb5/8yU0OLUmmfqu+i5TXd1zrqWK3uJLHEPBDegUKvqiz6
zcISrbyP+M2n95dWrNcG2Zzjx0LTINuRaujv+IzaDg7bow2SowawRpO3UAZyQKOpBP5K62bmqRk+
fBvPhOt+dY7ocsIZyMu+zVZrpbvCoHKR6W7CAiyvrbcZ97R9vWRL0wn11QV6i54s7lGvjgS0AUJa
ZG+lIOIg97UXqFoVyUp7i8K03djfT/z8Z8DuG40edFrVCXs9UaN9YcuGSc6335bDaD6q0HpCl+DY
JfCTA9KPYTmuM0PuZpSl3Wd/Yo4s5BaG5SUGDvAjcRFcDYEdo42jU+Z4IVPJV6oOELU0Kjqafqxg
xyNDr0p1FY4+hq7YxPt5F7IAYgtnLz9mLblFGHG/vMiF6PN5c75g+LWsmAK0JhLIwWrSIN1dktPR
xywsvl1zqpDEOLtpT/VaCibE6GajsTF+kEe/Nl1uxQWC5QcXKOsGNvPBVwaM3tB4/O/UBcrHZQ/K
jFKHuoYvuMJF0TLflcMt91qmGROl/j/bTOSOsCPig1B5bbaimHBeR7Hs/ck5yJGDPdyI9l7DcAfj
WkfAs4ZBX760UxWZfnKxuPRsOyYVYondiCkNHLZskHXVNXP61QOusF7HglyFqwx9dNie6e/nbJ7p
WCiFLcN3IA5F8MHKxMsbfx0GQmf0zLhJtXIHCwa/WhuH6EFzSmb9sBbDovAwrbyfrntDgHyQ2VTC
WwuRw3KTNEUxdkuu3C/vk5uz81MjQOZsiQlWfoeJXj5df5eoNAe0IZEYv4fk4PamoMFMANhLZkDY
FdTUcwbHi9qxIsnfxWYFMqce5DGmJNDzOG0EEp6PnUlCTiOh9N6edzVolKZd2mOMvXuJxPcUDvPG
dMuAi4MpKFOZb2TmPAGFppXfYp/N1PSesr1g+cYOkhqidgQpfZ1XAZOcIAoMyn5n7bxERcrN0yoT
H210uAw3iDxippE2FWBkJctaUJy/mGxIbSNPebH0XbFLkvMZqfiIgQsQE83WzYSqoD6ahp0Igw6X
UPcXkEGnYcYDjzubZM1jUQ5VrB5q3yYqkwJnE/7N/5FD1kQrg3C/u9vNcV9RdFWruCrQMFvQWGdh
o4tp9bbSM0d3Mx0pKCBTwQnZGMStbGjltpUh8cTrvuiF72mFYyd4HtR1gZsNz7KX77J6pvEojjr3
/dabMwExrmHTEY40SCAmFfl+Kef2BUvx6VT/stWLXW5iG0Tk2ccixt9FGNT/qPVwAFt23SIrIdPY
uZsx6s29wwJUBcaqMNFxyyeUMuT/xXW70hBIh9NO/VdcrictacVAZ6tvrRANOgOGkO/Ri2Y4vJ6U
hw2qNLJGiOQoI/m6iTRHetA62J1L55FhwaHMurvJ0JORj+7KdJGMgsdd6jpNp36GQCo7jTraPdiw
94waWFm3Puhwcun1qaOZhpOGgBfSGOFiBUGhnIczL9Y2G44kN/ATgdJ/1DSk1L6hVuYzFGGxpp1F
xh071bXOwMTS14ryUR23NCXQBEOBIQF5gFfwRgd7m6uor+IfDDmrSWD0MpFixuYiefNNvQt+2yMT
ytrAHFU/38hidSjF/45WcYaQwu4ihP8ivniNAQe3bVJKfxXzSVJ7ua/hhgv/lkPUbw3rjuMSQz/a
uWAdNig5f3enWaBP0yN+u2vXknnm/3AYWSEdkJqidlm0RWbh3ulyah2/ipRF1m0k7xIYbIVFL9Tv
GKr2L85Wmv302KvWkyVdhy58r+dSlEkm0s8CqpYSvINCm4gMerit/mOu28bGaxOwaP9T8Xiw9MXD
RFAgxDK2wlHt2Q/Tq+sGJHcu4RBAR4qiRfT7BE1Eu3aleXBlXDyhyihdeN87rMe6crQDO30+MsgE
qRIdJDfWo4K0GZ1mt4yvIxscf+6dMxs6xZVmnWCVrUUDNbiHavgq/87jb3fwamfwVoNCkoU7f/yd
qsvcaNUVtEBzC4L+V05Jk5RPjoXmnn531nuT9/iPDbzjp5eDnwocaWTsHzKyQhrdajpPcB5zN7Bh
hjUUnPM5f0u0v9U4MoJ1NS4Fgora7pculah42yaB/WKgJbKzLRxEmX9TZ9olwKPK3JfDNYS0rgej
R96l9eCn0iVrwtAJ/EiIc48SXIyfdV/2bpPMw9U9XR+kA/VRWWLiErOIfpRMgWi7ZuAVjfgaEVv8
+WGM7WnYQ/52SVedJ1hWhUlQE2IpCwNRUuokuZJJDvEJ8fXHSo0T0Y2BBZsjfdV9nM6g4v+S/ewD
s1dsoWp9slz80CCi9LbDgLcn+7I5z+JfEDrNF1gCV05D3c6F6BAVUD09Go4gGHDIRr/NxhZy9mUD
EElepkWe1zEqmS7rixZJc2xJaLGMK4DX8eIEj5s858K0n/tF0IJ/8uVpqyjcH7JwurLSDg+Z6dk8
5/E5smwI6eoRhtfHAWlDJ5IlVXbao7KzFFRzwSapqiK6GCaop7FF+jiFOhBIac4ld3WaKPSCBo3K
wg9izyH4/5/P7S0kKxEcgcIQcT0C65XpsV5m9fUYlZYexFsYIKg0b0ioV7bLicdrD3FRYMohJ0S9
/kcj7SQnMCGgkwxwAprKCDjR6jBh/Uh6x5qXbpMOMn0rwlPyASlo6+5AHoQtgPKrJHDiq6V05H6S
jtTM3urJk6SJAi064aA2ywT/DAyJZCaYhUPSCfYV2QTrJ61B8ETcCDZtMWI1BzeIe4VviXjH2aaZ
VdrfP8/TeQKrw+df2WwSPbffmd7srVhf/EXRazvARCsNar9f/xDvtE8VgVDwKGtARkwZUwgs4CDz
t4PYkTQgQYjVntNlu62paJHAgZHbcFjO/CFGzcZ4zB44307Nd4nMfP3xNDVpWpEMZB8PiIN7C4ZR
b44BMGp/Xyx3dfQDAklINIO/SGok26dgH0AVDg33mHe1Ifd3dmE3IF4a5EkPryBJRG1SPbesajF7
oLD7lm9MFuB5e7vZyntJVjB1jcJcO+i1yxoWrpqlNkGsTtcxyjlvuXNLLw9vqJVnG/95Y09bPueu
iCjxc6LULmpsbtLYli6DrA2R1i+m1AfvaxoMv6ywMiPpMTZpxGG5Zk4V++aMhZ2QDQk3ihbZeTHi
pMy8by4HZEZh78VuxIU/E7bLjAHXH6pxxTUQyvwt0OYZPkEc+TDbcjXXXYffPlPGilIwJ1KEBRKr
oKmhxz3H72/XEbyLfDUMakA++5RpGss06I2oFzYs7w7uXlJpaRO/44g14uNcvjMMdZD7CYOJcdeW
/Vw959xJLs5SvsL3F8Mxga3trEyXnkBjhKhzOT92rK2W8UclrAK+K7ImFZ6/XVfn5pfeTkEQCG6h
YQK8CuQEZme/cH18XydTe9n7+3fOHf0CkqXE+zU9GQkLeUxAt66iPio5wv1pOpqdXBjIp3ed0Ts5
HWrN6cD7h09xYGO2YvWNhD343X+iHMxG9XXfYZ6GUGYUhb3YaW3NgZ+bAZDVa2uqH02jS5WofPDS
hqyeCaiEk92NnaKYDREP8fscJkBlJ/CjPVL1KUTIIZqV2rUSX5xw7o7z9SZRhbeAgKGrr6YrPGGk
MCOvnyFLmxVnqfpqwxL51Um2wabc351jzvHwMyqwvYql28fJQixPrkkjJwCWBlXMFf3hUfqtxwTx
B18D8W6RPmZj4iD7flLM5kDt+5yE55Vt5HSZDB5qDNGDQPER1B4ZjFXB5rUblIzQ4yxhTS0RwVW7
o62ySmfwYPIP6WkqIInJfWWzexr5kpW94sOusTFGhLh17KILkfPcbvLG8yqF0L/SMYV2WzeFDSL5
CZ/hrEVjY8Hfq8hibP3UNMCNh+Qb+A6ocK5hLSAQKNY7kaAC+adFfImNSKAPv0ReLxrmg7lfAPqv
YcviVZPFMW9pl3BkYkMCbaXeJWlQUiOY2qFXm0kL9FhBDWMzh6g5/rGdjQe4R0S6VxGKq9+iyAUZ
yBbImLs3hme+zNirt9+SSwsHOUiHkK4Q2b387A6XTiNI3O/wXUqIrYxfFWy+jw8Sy93jXUNmbrse
wcy4y02H9iRP8ZhuZZBRCTZSLEGZI+CcKP+VHGGBwS/ZE4qGdeSpBunta/yqd2ZghzSC7kSO2aa8
zCI2QIrLP1tFylF1iQEQZlOAYTq1FnlV5ifnoTfHfz5RbPP0txMq/89CmQ4Dnfp1TGjVd3VA3bSa
QCoE8WZXcDwhl8E18pL26Ksgo1hgyOiCfXtoRYW+vs/LiVNKdKzDVu7Lolt7ADtcu/sHKUL5lfUb
I9FzNcZX1iVNAZmqyA9EeQEyFPJ54s5hCcyoukCu3De6Nq0TIrsKWs1mmpn40Eyzc5vPGhzgyEDg
JVX90mgYrV53cnU4G/3GzsTu0W9pdZlYGz/zBZI1VWE7mqlQrT1koLfyqN0Pv3AJEgxafnZHJ/y+
Ixv09t6da3OJi9T9EECTBtwFf06oAA5qMnnqvI4WdCVlD8wqoaALKt4sI20pK1vDG2TUSCmuhqoX
tRT9JQWGPTeak/eMLcEwOK8dr082r+eQOKygll7jrQnVygbArjUg/ayZyUMYyBjlZ63N8arc1VNu
ugHSBcgPCjo4ENUQcfjuKlM1METJ0BA1uF+Kds50aRoGdypojalN2vSGefE42Xq0ZsppQZUHRMNm
uWvYAk6AG7L06r7QFJkAmCKHwW/L49Os2TD6WuDjbPC3VbZoINnSmjSJ37eWYFZpm0HTL/3rz7Cq
ieNr0XsUO+MXKgYEaOQfc//7c9jnZkYMV8oRa4qqLwjdGDRFdFqpzELD2JVJFF8gJGc3ioCVlPUi
0xThWDjExStTH4zfNRDe+2YNruaDCFcxeOsd+MjKxAHZPbpVrMIOxKBYRpW0tOvcTG7Ax6LZpYKu
tnUV0SmOr62uI6xorC91TVtFQro8s+qooPbG0snHqellPciUYMbixLvDsX9+HwDRq+Z55BkeTLVG
Y3wsqnqC/siFIsByVViOVQBH9aPlPbnNxPh29NSi8tnOrbM+N74SF9hdLTxZEv7viWJfr7XV/Pog
5llQ1CQf4Gp4HiO2VCiQkhstdp5h9SeqlA4J5vp/2ZDEgP70YAOTvcDjBeONEcNnESk+u0ohxCtX
EAwfbOL1DbyrxsNptFcjocy17lDIzPcJ983McaguJ/E3+a2J1VKqm0W/UuSX9WiVHOE2w0yZnGMa
zRt6MYqAkWUw/rg6/EZTgZIZq+T/vBD1Wi+ZCg4h/4x+nMDWNSsud35AuhfrMyaNvSlyGbGVNY26
H3XlZW7mZyyNlBkyE9tLjmEJPDeoVZ2Yp9Dw4O5avB1sAEssJGrEQqfkfvs/AOymx90lCS5wBini
HzuRywl+rAMZH1MJhWU47t94nFkKIM0UCRKZ3dwvYo43bqfv/YakM+YXpupClc10Xlq6rX+8qHjs
tUouQgttW81DnWxhFRFN5PryEDpdwHzTppW/3rtY2Us6DwxqvozMxUe2VIZXBFf2McpIKVIW3wL0
Ua/KoRWOumwjE6/ATHT0itQPxCQmyqKoQLjMamcZJgQHTj1btx5whW9Dh/A14+nZsGc0WoyEb5jH
Kyuj4MQYtILaoNw+VulF1fKJfbJo+hzbTEuCzIT2jzHmUMa3xs2PR9fdr58yqTRHZGnP3h2nfHyo
EcSmGpFSYZCJlbdBFZ7a9J8A5shaMK6NQtnAU1slvzovtZEJsGCGvSUSUfkNYc3r7GqmpDaYJOLd
iMNN0J0Mwc5EOp88eKkvjNoNTXrDt9GtnhNoiS5m+8W8w0CFjNqMuWK0RckNZNP8ttw6Gwk02bbt
azW67mUYp9S4OxELoQPU1TLXYycwWmNxNPq83TrJSZYROS527pdBmilyZNlNZUNES9u/lEVmwZtt
KrWZNau1T3tF/Gl/On6km+uI01XPkm7QnZrh9RzlPsDH62pPnAnKQ+TYzCSOxfCOV9piVN2arNSH
OaQWaU186HHk/FVDcQreDiW0vGNlufWPeYfd0stMUixtGaeBVCU4uu/f977VfdXEwClCRP6uunt5
GF1lBKXOzAHdUmBJpDt290dkem75ROX4zELxfG4WP0RESmjP5urWS6cT+zbtFlZIdIexL+ite8Ei
AzMGQ+XOc4h2wqFtEmIw2U5/Q/gK316SMipJVUgvWTI6G+mjwj5kCkJ5Ufpw4tIR2bbYfhD7NdhR
Seu6HEqLUG0CKlj8tXglfT6EllZdHFk9kPpaOEbvKA98YGLoXko/Oi4u2AtzQCxiU6B0EmzppXbV
WE481UDfdwfostELwlOSsTxwmJ2PaY5jY+isEhr7MlJtgSzOhT2ID7mY+Qniz5xbsa/QfOmAQxge
U796PrYX64Glaz82JBg4Ws/p4cT7nLGA+NkoKqsvjYn4beKJqVIGwVpWIdcyQP0HAfzI9g4sy1XF
5gf6CQDfuYXwukkxrUndD/ASmFT9fHLr4MnyZ3x5v6lYpb1WZ96tifb7zipKmWeBloLeVxYdX92B
BayucCV0XnEdllB6ekel7TFUYHiTfpAMDGHYVIct0TLh2pQIFSqF+Xo2B7LXUNrQ8H6RVPgJoZ1p
jZQNl0s24eCI+TpYfPHwo/a1qOpfgBhzzA7gupPjsEnTGBPSQtCu/r+OClHf6hOahp3v2i70r0NH
ncdUYYjlM1qI002ZX1oyJo6/mK0tmtLHUMkdPfg3E4a8OAt6RD46dRju+VbUUy+oQbSambFL0PWP
NbG36ECYvYVwK7QsZMh8mjMaAUZhifyL6xDUd2QiHuZ/tWc9VYO/vTDJPNUhMiQTNhYIO+2BM8w7
8VtiHjjoQ4U01jm9RiFxBP8CaIVdMrOYK+FiZe+cuNT/tOCoEtuFRhwmEJo/dj5lgDZ3usQrMNn8
iZ+pcUr36PNRkqzoFehV5GYqF/eEQVNMD7BMq+oVVEW42Ln62FpZaAdvrhS2j4YwlpIfn3SImgU1
SBU8mq8yru9p4Gt4+YtmkYJSuoWEtbw7XZ41MS1JQaYBQlA45c/pwbHwSo1361v0++MxuDh7Pwpy
/mmnD7QZiqnVKjfFAEqgPwjO/aHHwK5s+eFomg7GYw11wAoUGqRptlI61htQT0H6BOve109tzqYb
kYBqsYjQ47N0iq6lanHcjmNbb6ry5zRJUxBHmPMnLbBXx85u0XpAF4a4JjjImRiBMZSQjaJCFxa0
oTbPYymAwZbHe47PWEdZ1HpX2sZKmM4J3RASHxuO2aoF++glSzVCqcc7ZOOLxC7CQinWce4dL8/m
DwiASRQGUiAajut6sJr27tZpn1h4SuNjc8d45cKN6FmuJ76SoqySam36WQyBVtPh3FS0LNxm7/u1
sdEK460XI0XEt7ReJcAE5DHQ/2hD6ybkG4L2QmGDmrwUgWUtYCTfslwq6JXCrj+KG3txOE0SW2ZA
nxSFUQM85P1F6ytrrrAqzIUBjcV+PMJCJnZB+vY4RRqJ5AxUEYVafJnPkWgMwX3uG3xADWCAwfNQ
YGGm+W2G+ywr/w+LSF+/akgPe5CvyTmTHxwJpjOviXz8ZAJUDwj/opk0CJJFKQArYdeHDw5OTMev
CwPdEkuo/Snkv+F/VhTyrSjNvv1p3quoPHiQYp9JtSz73Aiyz4ym6pt1Ik8kZ3bVCNhmyoU+NA94
JNsacKsfjSJd7FMxgMYG+elxNbIDOIgvEvqit5Wi94HwoyzuwKSYjKr4tzPpCE+5snCvc4HIeprr
RNpVCZ15bDgSqlmVFmx3X7e5qLzwU4fM9mavYRXWNN1hYDtOv6Rb1JkoPJ1LYfTpFPv4JktkVuDQ
OAD+nmlKY1EHuJIp+8qCAzFSxQzBmfN2Bp43ybTK7SSR5DyfjPto6a9XDHd+u0B9y3/4wq8FZT8M
Srd3ifayAXUkb6qYKcpCCf8ub/bSVQQqmNrx+wVIGSi/Wk4AzxjcKVD+c18GmEXEX2nJTHIJ42Se
W/rHeWzyAgVFcv9FgxiveiyxESUPhtd7A3uHpibNmqZdM6LM7egOGzb159TK7U+ai03UThyUgZUo
czlb9smIeVaeuJNUgt0vfgy+g4+rfdNLWvQzJV+5mD5NmJThf7ncvftlQ6PxyJkoeNTA7xXow8jH
kq6PSurao6MVHM2Did81NDH5bUWafZ7FzbQBriIcXZzQ+oPPtky+QP5JHXUK1a5ySDO9uu0/GMtO
DhGLORuYHSHQ0d6kpSsJcsJfXtRQVBZL3fLysOULfvELcPd2eziV7CqhOO/iAN7B9SD9+YKffY6R
M1ONI+eLUbk7KBr96ohmQwqLjsPpPaUzkTuxzRG4rlLvE5XxKZnCp3kl9GYhjhKHD3jIl3EJn/Xa
YB9rsXuLcHS193L89T51Tv+keklPzN3AEi0yk2qzANG+onPkA7IxHm8NU7GBFYOnt26JRc+cC5Hw
OeNEh+7+4sD36IzPYEjSJRKKQs5Gw81CWiTUWXqiMLlpeBwh/6fa1k0HfC+A0n/1hE9NVSGDn9Vu
DImiNgTjE3/5h4miOGCAlxXhLSA513mpu6wVdS4pdpuCwStwbJzFuDIp2oYLTgy2HvQPQJBhZ/hF
KwF6MDv0ZLkluc7RNSHSbn6C/2rBkvEsyh9zXyJT56b7Pm6WtaHQX/oTiwETa/wAOg47Jp7qAi7E
BMVrJadusuFYO18wHra8hFboQ0VsShj1xPdvmRsx1XIvkiQIMmHvLhYmzUpeB9rM0dfmZs1nhVUK
sZQbMn7rgHe8DrVJTi09A9r/1DzNYOpy+sVkUHrv+kin5WXxnns9+yCMDyspwSI4VVbg1YKhDPzR
7/nlvvjYkv9ktZuSUrXQUeoWx883r1CfcvgH/5PupR0pTEOSSeBAZWgU2DSdKGdHGfa/306n+O17
5ogKWV4OoNyicV1kJdRqsMua+O/u18Kb/F2mrgMHBuP0qayiDgrNJS5TEnjvSfyu95r8ZtB4wiRI
9aY2XtwRHhbYdYExiaooDXHDaZb/0jxX68g77EGbsXZZhucXseOLbk3RDn5dbXOOiW3gbNCA5AdR
ew2PL8prMZ9Uhy8zyt7YLkLMO46VoS2u4OPCf9O2DJO3jayBa/FcIcU2nxsOWOWQSDDwXWnBeOZb
CAlI+19klnxWlI2dzcu/VpbAgOn3q2ahGL1JThzN9VhlesuthokqzOcvjpkGH8cudEE/16++qDvI
44jwvQEF1bQzV5GtyyWh5ERO6/sv/Cjvuq5IQdP3PEEvGtslhJ4vB6GLITOwvOXbRma5nZOKl32d
ZCqumHiHxrmL/B0MyzHoa31O7L6UnNpesfkWz1sV3nF3iuA8MyQ2e/LBLWACR9OxmufL79aKTHF0
4+MaEo4e0vomC//D2ijd5YWYqEASS+gyFtHzJ+1JQJl6AQc7Ytm0WoDQ+qy4kq35V/2OPJJ+QLQU
05QLyjDcDufP7kF5Pq6C32E3r3jZPLS6OG1zRp1BjT+TY9lOuR+ACSpHbetGCelygM+ijjG5C52Q
+wDZ5kQH0gNUb7xI45BuvhLL3ilgf7yBqcDy9QIxHjjTj85HVDuGy3Whs8crEuMe8tgVj+XB7+Uy
99nT0t4QnBoN7n28bZ7h70d4Zvu0S6wsWZSSnqS3TjvcYMQQFDjxeZdn9vGuv0j8MTfYlE1zPLVy
3kIrFdjRiImv52G+ACnTVwPmkWlq8TYOnKTH8LZNW4c6MpnWzMbrwVYDJKRVXAnzfHbQmTgw4Cx7
uPQgEVsiQdiyLCciwhNphu0Gbl12RLQJddI2EMwtPV9bVHB3jJlRZsH6ENNpeP/4hENOEkhkW9Lu
uf2zj9FsBsWID6jFDHpqIxlWNFrwaxenKiWCfM+j4aawOglkjpX8DQWo/43E0CKyZqt0rS+aBYt+
zZucMnnW1ls50zCuQax7PmD4tHl8P2xkg7qE8SkOEXuaUkL+/PMK0UZDw50WJIjCoXT2RW12WisY
NWS7g4RETfKTEEUlMMGHBlS7Cfs+P1wHR0JrKrJQ57AYIOSghyFrksZBaqsjmZxjkN5C57Hg3f+M
W1EU8NLciP2t2rv5k9cNUAIg1eoApGVlyWrAgFTwKyDDcXAkQVpDMjl0kFYmozIRH/WFRilKT79Q
o2Wf3DcX+mvjpdS2We67zg4jgkrOeK5tmNtQ3UMWV+5025gvTbYTcG/uaWE+18tU2JIfJESINcGk
e/BQp1egAfFazxdudtN/hmPECJZhT/yQCrJ9TefdtqdLa6hCaXAONOfrCyBghAzI9qNh6HgLyNwf
A32AYmugNNcTONTe5/ct6DuWth0gBhCzAMnJwz+pBLFoHwjPBs8RzhxLHgp18okCl8t2KxblrYME
2eKV8ukOVStKmNJg+nxIW83GH9jCCV9J6wrXFMLkTFTfGrqKt7LI3K8jqYn1e3wHL8fmHPbcaIKK
vheodsOvSAJ8jV5PQK5VOy62gut8amPkhq3TVi4c7BKL6TauBw0Pi4urptDk9PZ0Iydu1JTMsPM/
Se7F91Fd24Z/GakrG9cwoP9aTuoFkNxhnEkt1o30I6BCkoH9zbsGPwXXI0GbvIXdsvzN0N70fRXw
3/FCXCtmwbwxB/9F/ybZi4QZv79c6YMANjz3SLxX38SYgmZ4qkAjDfNYcVr5JSFlf3vijJZ71OkS
preQwZ5BELWSkEIb+u8+RSPS4w9FbrgA326ietWG5acjZOlQDPiL+TyAGXGfFIjrL42P6n/wVZAn
iRqpLMnhNjWGNsOHiznV3xRJ5fyU6Zz2YVp9GjL7CPznU/oIuM73bJhJRatGPYfQQ0KYIs4Yo+wo
hIjA1f1pS+g4V+BrYJW2CWzkW+UsNH6ttE8/EBNETduOyIj56BAdPFxn0qhI1fCzYcfj1vifpyBk
imsqqlATE8wwM8TVAeE/sEN6M9AEVju6EqRNRlGwjWFAKqSbJ0TWO4dD/F1HZcrGQ9/EG/1QT/MH
tNzAVMdJWkmRsQZdttwJslOVxMB+Z3oNNmP5vW7+M8k6PX8FXcNVboIm0r3uc5bzikt7GyKjNF/p
vHZrOJrRFfgQDjB7Lp+7wlE5Ly/DzRwlaFE7QsL1pLrf/x7ftHHbwrNDZdxxA5Sa7RWxpuqFvHGn
PDGRTUyJRhh1DREIUc/UNENIPG01Y8IIlSalwUi7T3kFHMATyNbZ8fGLke8SdMjoUAPuuZQ9owRp
9t+r2a0BdJdhVlpmfUul5OyHHMcwSCy12L2dGZzRU1paF1nwmiZzT4LMQEqmHcUUMpSlNW3IGdyk
J+BYDmDcg8qEorVAUZu+vaOyS5qiD3FIzNkERiMmPfJBKFnlXj8bRcUh0CuQnC4o2mJ2twbFo5F+
QUL6PaYrFmdxeYI1+2unUWcXL0FscLaGtQpcGYS6nKw15LipLiAqLxLopbrz37hXUZ4XgODEjuIL
HXlBfNyBsL1C8m4rT7NsRthl7o8AvRjAAL5n8zgtAxWtMxSzvWE3G1USbJJMGIILJ3S4qjEh343L
XW16VYU9w/EfycWKbFnPB/hxq3lMRLFnqVfzJ+qLakrnBalFFSeysU9CZfbJ8GBOO41NskTiqLym
HFrpPpCEHJJ5XdOF5kWGrRYEepUh66bQBJdL9DY8EYBU9RF5PHLIPgIn/1JVsajPcK2s4B4Ee5WX
cdJ8vWZ+D1QkV1VPcoJylAPJ1EwEyGBOgoZYyb1n6615ER7ER1FCVv9qLj1Kig6m5DtBqvWIZI6k
KUMH2vowOjbZVrKcPZVUWfmLYHDR9PebMhef9mezRpLw7u8cVyKaxwyqAvPaS3fZ7IeZ+RbQ9vUD
hqSmcWbWlf1rJHHzz7ByNOU0zH9A5Fhtedu2Gi0aUrSUXQ8RRyrRrKp9M1a56pWcaIna9X3QxWAn
5VR3wxYHlHGUqa6DEeLwfoanP0y/0okOKSCITeaO5Ss9EKxbLq3dX2JD8QMNfgIi7hfzmYgLzUMC
ZjEcnmmC9VIsslJZmqtJwsNwWzMTvU8Rq3fQVtEGXRJHwYGWT/n+y2tLK39DWZY8FAPT0qJ9PMpQ
1dG5XQZ/Urh6kKGxLs/pQ6nxVb9NZz/67cExR0Y1r92UcoxS5J87qZ3pncBlTZMEEfK/8roMrWn9
cBfbwiLyE3jieodsJzaBFvOATUkDl9a/H6++eYeLGzXRE7lLMYupJxzecwN3td6QcwNSIb39KwbC
snjHr7YzYvONWfN8/zasIW+cqCjvD5jFb/h5uOYC1EZkErTX1QCwf357Z/jtBBHUG4Z7DiHLLi6+
CwcXESa6r2XFC9aCyZ1ES9GiPN7Hkytu6eUR6qtKM3aisR6eeurejR7RPZHCyeNAlxKXPnuWc3iU
mMk19mWiwERALkSE8VxMd1zfCj1qpJlAosu/4ZMlzpeJjOSpCv+6iv+9o0mTNY3VLxnFWCDRxTi9
tYGLg/DrTTxQaFSXvWhSyzSlToCKX8GyM3TSTZv+rzhj2ivAvSVS3Jp6kACClGadB+akQg6eIVl9
ME6jCu5OnztLpZHoMEg0dSzDVOAbNGJRW93bmYjEOdKJoUZnvyFhZl+v4EY273g4xbp4SNL63epK
5Mf6mPJBySh/LiSZ+akS3r6mm7OrjVsScU7M+YsdVZkuX4ZkZt2OYaEmPhgQGsh6WIXgLkqRRGJM
iknZ9NUhKZ9fNe038yteVpok0zEBv/NRPQquIp/nXR4EPbMFS9AaBGhNeJtQi7CrCY/pGs9WeBwp
xWVUh8eyWfaZqIIrY0PRwvwqH0Gg8Qy4Xrk2rYahNQqPK4Wwn37mLTe6aEC+SsiTCCOBfHX46lS/
y2Hsm0n0w/BFVW/Cref6KixVHR4vhOqF9RVQOyxgvQzprvxUdBHsNtUDFXp6a3xsb3UaSuMi/ItE
HqkgmIT6z+Oj6lufUDxSUjsBGvJHq0yGcDtjdp/Xv1mWSqgv/3n5jbGov3jwW3I8wQDJgjTOUfVA
KW04WVIdREfFl3Dj8r4O7181rphqx6UvpFBYRgWJvMhTIB52TwTzeNPWLdiq1lkYaZRViOQTmx8R
PPKPnjnRfAslJsTS0vkHkGT12OzAApTWSTDJs3zhN5zSSVvwXUsI+Oh0PWPjEX86sN98f9O5kR75
5tYRM9F505Sblvyx90X+QFfyXPPUc155+lKJk0n/vzN6atUMnIg3X0ewOdrem50/jP9Gld2oFRqI
wDK1XaRz76Hdb3hEPA230CDzG+Nkc4GZ1g3tl2hvPLzhpO4q01AmD+R7kWXAgw/qFE2bF6+6vzpC
X3Mc2aoGq00vx2PvHQBa55TMkyFQdT4TrdEdQbcWbqPA7bLDz/S1vhO5pW6q3O5uoGUx71ycA1HN
rtWIUp5M+592p0ORdYYyt+FO8F+Q7wNiUDmrOxrJhmsGw/Wfq0W2N/R10MxZRtLSq2LCg73/WWz1
toZxrh2jrALFu4RWvCWR3ejrpt5INTS3FQ+i5+hihEoMOAintLxaSROkZ73nwXa49ta0C/tB7tsQ
yvlJux2VAkwfP/h3hKG8VpN05DbBZuojnzUcyO4Njdodpz2ApcOI//EHdmn5opREo/tbTKQcOa0t
4x4C/oZyFmkArKeRoMTBuw8KfEC9s957F77vQsnrtV9Lg4ORvebeM3XFEwyBAJT2NeQ1Rif/sXpm
SNlPT1sRhaAIfdQsqmCJf5acgwc0A4Lt588o5XsrYJoSi87bUftj7HZ7lGeuTgtWvW1i30R39WaU
GVKmLOc4pT0ZfS1J25dX0yf6U6qY5hB1eacRQaLBGVPfzp9msd4ngrxuMRV+okf0Yy8F+N5ifFH/
wgH6RdArbWKxolR4u0HmP9WJZ8wkkrmiOU4t2gjzxVONyS1H/hJo5IFZwsuroXk1WrB4TypkUnUA
78lmXhv3MKRuG68+2QMjsShwN51RrzkxI8E50QYAC/qKnKpqHAGtWaHfdzior6Fp2Kch5Pq0SRFn
YH0zdU0S4KG7cgym2HvxEfMKHF3JFgkikjd2Qlrt/YEyDcHhUM3lK2G0x7S15Q3HYcE0qWrHxeB5
shotSGGoGpItzbn1bv8O8lp8H0G3F76NeVDgAbxSOTrz0HqYW4L+RwL6bai/0UzW7COhqZsbxdDt
BA5XXlh+q8Qe316EsJsziMbv02aIOzEb5VCgBPQmsYhJ6weRDAVZw1TBYp/FVSWn0kU3MzGNmY6b
WoEs/OgHy0e8ddUHcxtaDLkWmj+xDQmU34kyTXMPTyHM4zXjXyyRHhUeDamfKLdB42Qg0q7a6z0U
IB22W/618TLVzyvn+ib6cRh+oYdjbNhpyTRsRNPz8Ss+mBwmtgMlUCe1Zn8aIDaQcrVvStu5Cb9s
tXxHXvo2h1rzwYVEDtTsn1AliAd19TMSzBE0H+ehqTxpgQN0PhOg+Iwg3WsR9MpcBz6CWf90RVgb
ZnsVvE9xhxMTZER5bkp9TeGS6EdTLSANkKbyzeKcD7GqhKjGOwsPJ/1CyHu8P4N8I9Xr7zXyzgDC
Mg5+gy+bWjpaurZ5lqYWusviv3b/a5UtFHLAzHR8e8KPJWit2Ees/yPCrBzFRCs9eO7sguaVOzhB
ZZR4dEeoSs1gQEjPR8gyo9S55WVbqKTQlQrbbCzShMn3eopjWKGwvwiik2ydi5G8yNEuRaSbVyKR
C3vi7B3sfGNAUphhu7b8tF0M2aKmkQSJbSd9TrIOWantsJtPUAj/99K5Dxpvmb6PQFg9YTM4av54
2Y0ep2CtGyYaaX7PJNZc3pOeS2YiGOxqriA9ojrr7llagBA+9RmfNLLMdUyaFShty6vECy/H5Op5
M+Db1JY6Q8KBmnYtzSYlb1RaiaiYiME6ZaUOVHrioMEgjBkR+GddxAs5dPD6rBP7xdZmoWLQjT/H
CheP4A1xc5QpzJHdNlh9Uvm+66yAv+Zg+NZWjHD2JXniqh0aBI5OM5TcjRz+ZPF0DEtR6eplQ4EG
rkSpLRhji5TtkvLa7rDwzI1zYQtr2cnLM7M1Hten8XlMkS9pG+d2VAx7YGndhsg6aaef1ozwILbV
/+4TO/g0nkWX+z657etyq3+F8UEgd3xS8gRqSGJ6aTEt6WnB1gAN7we209AbwC7hNvDSHetUBdQ/
nrD+IUK2QtvcjWCYnU1xPmAIMVwUTFY67d0XHXEbjm1jH2+3HGjQeCOlUXrRuI2Fe8wdG312o1wF
JJMaTRsbHdl1VoFS926uyX+O1bTTO4wlgI+SAde/LRhlk8AsYoZFff+1Zq3+0aK+8B+dewayMCrY
r+IhK5Umxlm0EblX4UdAzL3GsdRKLO0npc2CU4olKfuqgjhUVLJU3zf1KEGdC6Rs1omAbX4uyISW
ltq+OpOnxrtRqsLltcV/LHcgNbAaLESxwp0E1QOluL3PtMD5PhId0rEwvwu/WcCe3ORg50I2IIPo
H3ScsKnPaONQYKafixVVGpCp25FxEPSXiAYTdESjrp1TfEmohLi/urGSKfrTrlEGr89dNYtYFpvr
OJt2JV69LSNf1vDkStwBekeBhuyvhSHRmEW9oK1LpGusJaBJV8eksb/UzQzq+6d0/0Bszk+pDHxv
IiKL1Z8LzfkMkzAcWtx2wL0yVB5f2t1AgGfubcrTZdL/H86rIlQXP4Y1kYelHNcDAEnGGJjG0cr4
gNNKU/ENRytYDhZarkyGma7KQxBf1VyzRzN/Wl2Pg/TRdnZMo8lz+3q2vivC7hbfTk94mD0w0sEr
OcAK495O5SOvHhiN6GKlPEd3NDpCTTnCmEFcc7QrrWhpHJMsLT7EaO8eVTbedDTDmj4LqqgZr+8E
pYvw5fx12AH4NfZVqOOsSEIVd/46RR1FjRgn8JpwWYMzETL1FCbOJVX4DFK9XMrEXl7zS7jF3Dy9
+LTeyyOhLR977KmhFKx4I/NjyLKaUrhMhIcf0MyCcHDzKuEzSGnIDJzlC5Fpw6YjCT354ZePfaZN
xWBaxypPcKSpXqDNIVrNAr3A+TPkW3NnZ3dF4MxsubjN51Nto2aLc4gNM5Ttl3hsMZ68L6UT+pxI
prgY9n8B5hVxftPD+RRLtasFX0z/bliSYOYBOhaw6ya41u+vZBSHO2zUfbBg1Q2C0J3lyWRwCxmn
cU493MiYCBce8HtHCLuDaF4YOsQivyJKgdcjZpneETw5t4hrbrx6y22lGDbGB9E0W7dhJMqtLRoM
SGliPWjBryxbvN9bfXJs+sd0kYeK1M1GYL301vOFA/vgu1n8nfqfXbj26/FoWfLcBtadRgHAeARu
Pl5QaeMY7zW3f3XPC1SKqchjte18SAfNhNbZT2+9T4mp3IsoWRHALGzpvgh6hwHIBjsK6hDrB7NY
o2b2q9YO9ur4+BOXAScouGu8xNb5ZasfSGew1pa57YwgonCr5yRxdCeqCCCm+IoICAT3Rud5nFIR
wDx+Tp+NRjgg6Kig2degC2zGy3OOextejf/H4DfYqHpGNAmrrybpdUtNgVTg/Ovu/oJaATgXUhAM
AeG+Nv/rzC1Lvksy0znv5MUMi3Qb6bo60c6lKx7zQAnUdCj2N+nkjiiV+Y0PotyvF0EH5ZAXxsEg
E7zCMUBUtIltVL9Sy7qO5OvUl2umrIYbIiLwuqls0dTCVtAwlXNiVsTe2qY+VUC02VC9KQ5Y0s1X
9p6yU74nQwOcyb58wQOP4XTBki9paZIUkpgO14sxiNavSWkg/dVo4DpJupXKApyCVnk+2LG1fmj5
GGmFJYLZPvEzR+bC68FxoYeajn3ZBHIojqxO5MJJzmrkSJnNYEofbA7AbffiMmAiTYCeh46w1qf+
gz9JKblZdCg9CuCCtkoOyadJ4BgsTZ1F+DLLHVL+yG5ynFuef9sOEvMgwaq1nQc5EURVbDIn/1ys
KVL/V0due92fWd+6PeJ9HRb1kcsnrVYujlLdN5XfhVJbV4idS/NZx4NNzyoLfS2moJxei3czHxo3
fPna+T3rPwfVj8ZnbrO/VBD7FoicQ99PnYibVtQoXji/sPMisZikN37G0g9DZECmed07IJIo2tUI
9iC0iI3VK6gtNUi+HVeB183x1Viq+yNfPJMp3juJThvPQyuP3WJxU/KfTWXBa0MmqPXMpgy2Q2X3
KbLdu9gDG6ES/qbXE3GmgtvUoD756q//9DQPrH7Y3cguQKtMBTcO6bLHoYpDLVrbK8y+75Rwefw+
J5SEkkwuHmxvrUwvuqN6uRu9J40iT8El8bObh2JR6rIdgazv071KwGCxWiJ7Tg1Mq5skOHLA0KhM
KxDVfVn/8INlM9dnJ4dFgirApXJtZpmFjVxboWqvElrZAZVuabxqHhsCP/i+z50raY/Bz8o6wV9G
bV02GEoqgdOZBgaH7+YIGqiEeKtnpXk4Yzcw05gI+VplbtfVqEyslIl6IddUC22AtRbAe0q8QGSq
i6A4vSPmUAPWm6SbovKHzSVNmr/FEMxtOlZ5ZHkqPeoii54+VNu310Hcn2597sVsB1Rp8AjpSJVD
wusuWgoLwUErAEaOnGCz2mIO9xNW93mMnHiVP4LKzL7NU6CXXx2t7Ba0XdU4lJV/aplvleLpC3W4
HNGbeypGFd3oThPQkib7hmWG1bxJivery8tgR41dXp7C0ZVl+WsNXR7KNIVBNrNu/xoiPdT97hBC
yyBFeky7kFP3i91enDa9Gvc726/ms9LbQs30irba8bUeTouwjg5z0Xt0nfe9jt1aTqR9wwWnL3W7
yQhsPjkrgVRR9sldK7BYu0af4vgDjJRT/ShPPxRpQ0OszVkvx9Ob0Z+PlGWvoUox8UTR/GJw+laP
3YIpA148g3ccVrthS3Vs6U02Itvozx1+5Q02YwkY9NMo3Jvs8ikhdQXoRYNfEy3tasOauuff7qml
nflIRgdBu91cxkLhuTyhcCUoHEjWrhWruB16+S+IpssEFR3bhCIFfj7CMsNBCIiyNjedV0hsmP4t
xzmXxO0gzIEPrMOH0d3/A212FiYJh+HcpsTr0sSKqdWRnQhCro1FBi4Q9TstAEG4z+tY9/n/xduM
wtVwgTFmaCmyl6OPOVy4sS52yTmuY9+GgCZjPC7AnmufXx2t5vSasDG6cQjKhjrXqBlO5Jic6AGC
he4CFYBnm+sg0pmwuaKp66YzvZpC4J522cfuZyvcJN79vbAvSz5Pqhp3V2S/4hy3pn+7v2dFxhGG
rmmAOMMdJQmh+vijginUSn/SJyXebaanc1VHybNUDsFnxOJAixYdJucz4CTwr3CmiG2D9rEnZn62
R1bNpOjH9sYlIwud3ZEGJ18piudFiTb2u4w0DgU/B1mVxGgstoFwklWjV440JQFt2R+HstzPFLBo
DsWuLvaXi4h5nnEHmAdVi+vkhA7KltMW6Z75yuTLdKBjJ4ZEWojXtDD8K0S2FnL+At30xOkCzS9c
i+6O40FvhdEN5Tdwh4qUrWgnpqWEj5J+TeV8nsS129XYSSK94yrCyJI1h6AwBekjKxhQgB+52hgo
7tJasCNdP7wdxdXwBaOoz2TEtu9cA1QGyU8XMvF7qCNzeBGfCI2t7vVNAb4lKdvtEThhDEZF90yl
sjfDQXpTg3fSMjdqqAduG1Ga0kYCS2oaH/+jjijX/MkKV5bhBb3QaWP1LjPnwi+IxkQBsEcNjVpq
dI8N5wOK+98eI2xiQTlMO5CMj4yJr9Wr/6PyVKyEjQY0H8VVEYUJTx9okrIZmN+UQwGDm0XhiQpY
J4FBSRs0TvZwiDe8wUMNaQtpKoLpT0V0fqhIMP6QW7W27LNYH/3MGYH43HndL5cg8AKMGTOHC3Xq
3ts3w2bbWUxDzFGAbRHOdsbJlKdZJD6Fw5BQUpRwqU87UvY011T6AcgCjUzVSBk2cjgsG0T6nOM4
QWlvKnV8suhBVqVlr0/OOL5SKiJGoAYWTRZ9BATyT/oqr75mCrd2OLJWGSIcwW4q/+5MCo3JQMEl
xL+ZZOeFRcyN2VErZkBUdnVvvSUzBjKlVnNhkoww/gkU+etRjSKg/XNh3UQkJ8WHx27ZVjCcR829
30XE4bphr+p35UhX3SRBTdvxuPd9iwZk0TpfLcCl0o6Z7eDv4DWPWJheDL1yvwFaXuc/wb+Z/rQ+
IrSO166/0cZC9kAjlXSb1IRJmt1w3wHV4NPxM4NXh2MmQmW+ZiEawG/zWqDux6/AyWUkLaImWhT5
375DvHDiCstACpkFtK+vqriIBEXyr+qjii62O5qU/EVsC+1i3pAhhKmGbf5HFNJslhzWaS3HFR7V
NQiGOi0fYd6fmgJcOhm0oA5wTumLqgJTGavMmR0/HJpyty1PCeP1dhXpqb9e5X6mhQ6+CnE/8gR2
0kjcW04YcjxBxOUNZGl1d14/kBPA+9Q4xQMD/4QBK4Z2ikHuKns/ROjbGfokvzF+a0Za5CC9PSYP
ye44moGiEmVPYZEZicmg/Hf5Du79Z78k4qr2vtuTZO0O9NWzH8j5Xdp0lTM5U9ydGF0jhEHUwT6B
33dzO+Q6mSBPKYnCngcAYC9nkpqXAN/g2anOPAQ1zoAoz+CfgNxdthQju42269wNuN9MNUCLYngI
sfaJO8IQyHf1JyE+Pj9+A99n0PreD/j0AAov5tVXAL+xMt/eA62rOKJfhyyW9QhzmM5XbQTaJuHU
um0LMPsyqarXJ9wuzY0ff4+akPKkP0aN0vdwF2CcarEhdD2Ag3Je+tC0VFmRAlnc/jLaSyzsBt93
it54PqrQLfQeE3ymqQogiDpqF7yERbPProk59BptjNrt56TTmgHRqy+5TiJTKCHVUHv9dH/Fk1qN
y1inv9uFbAU19dDlx3FEzhEU8XZXHBnUskaZ7A2BviU/LRyKzMo8vRv+plj+O2MKDrMw0ecKqYiT
eLLaYrUJvX98KexzO/E9iQQAjfFeGXdWbS7HKQimLVPi+lfRdrffnDRztj5RWT2P1AQ0xOPaDXdq
HrGPJOuyWAGQbFOwjRKNWALCX/40+2Ll7QzG2TEQNBXROHolby8exQMHNlIRFJQWoGKFGZFFr/1o
f2X0j+4EFHKtt+vm9kjnZ0NeWd7xxCooBfmCbKgA2R6i4O3NoyHULm5skStnY+sspWmaqvlhY0l7
27wsrTLw6EIwUABoI4xYExZEzlOfs0RJjqO3ry8FewKnXHkXerGIKcmaMWKWE/j9W+Td2PQHe8RS
DK98NKPozdfMq8Da269U6A9RY1ZgZ7DDjp84CalXJ9hoD9Eb2OA0bD1HguunZhjtYsjE6KX5Ppb6
LFzjw+bi/qX3potO/LUo8yylLcMsFCJOh31UILo4Yo/RQeezFInK/t7XDpmam6LBUPFp7qHXVgoA
bVeesq4uLitmN01R/EBqqUWarhFT75cwGUYKQLcMf9HIBKB4AmcIQLXznHSINmRYg4kIVScqab93
AtsYxklwAtKtV+HTrtPqgsLfwCUsoBcZFxifqn6v+aeYHP9f1PnIgDZyImQkOiWY8PrPw7w2/9aY
8VmXORKzUv40qha0SkFOWQXSmkiOfOrd1XeZOZ8AE6e3L5/KBWr+7QSSi3bnSHu5gXnDFfptUrMT
xbkdRzfoIxn/eKRF6Lvw7lGh5IUL+WFxl6lPTxo8eXEEdyP49vzpXM4agW2jzfaSfWRW/bTCFPwl
C1Is6+NwU0vRRuD65SZeJjt5CBNzV252FIsSpyUObOADxzpla7MZ4uWu1Kde3UASvbeLxNTVMdtD
Xud+ciksDW25U2h6brUfFcxkm/KWT8SYU25RsYLsAKxSrmIOkGg+2InkEaKQkN4mbjKyjltddVom
UoWT07fzYfeswMlYuKQfMkZv2HGx3OhJzeh1l55lPl0D8OWVASd0+mJf8ZGmR/hXen3AARsnFhvd
VHW2cetdUyGUVsMmLhazwIBoyx+Rm69L36zCd2mK/Xr66ecOqzZEN/3ynICM60ktUTtf9SRciy+7
Pk27Zx1eOcw5rxgDtYiCj0ls3ZOVkbWZSZEZssP18Msxgwo7pg1cBOV30BYfW2SAw0X1SovQZLR1
cvH5p9cb/5m8QclSTMfzBXiFwe9uYBIHOF8GkJF2Ye5zgs8EURFKHKzpdRbyw3uCgMMDuwV+qmb2
XxhxuPavxOlRSQ/UC7WZo8JJESBWELGAXlyH18GO1Lzc2hzAIkauvMBsxmO2kRtMiS2EptWZ1pJH
lrk1+z9DkkvzeCzFRKPWsGM7/N7KtZcgW85jEfoWe6+I3iGTXLOwbFDWjAXVzRn5mQ6P3HJT63wq
UE3ec7gaVdNE2WTivUeMywR9WluCQ34SRIGl1nkoJEm4RTGsOVR9Xt/Qx3/CKlDED1QZx1B3NAkV
vaCmmHP5s0WrKYXke8mtjZagDcs30NUXuk45oc84oKlMHJ42SnLbWzW5YnGrF0obRt8qM7bnSxrh
dIxXJtbe5kJfPrlW7TbAdzCerVSX9mHNQELDAGzoi4jsdV/gNaqavsyeyoaxV2DIsNf6/A0CQ0xI
MYhmf0Pbv0E4rPQZjDjnKO7zQZnLF6SRCUChBXOzj/p4fL7CK1ZN5LuZQdMTKhY/WqhxdOCgFyba
Cpl3XMSIYuDAWur4nGPtoauxGasZ+MQSM/SlDCALQT4xqFGVQBw7pAG8j21FeQ8FrNmVaNf8qu1K
FIISzC0asB2tyUzhO93JuiB7iCRNgW3PAvJ+rOJI0vORG9V2wr7QmIiIzgM02tbGpw1wJCEmVfrK
2rizyDwjEI8kft4kVJzzBT8KNYJIdiblGbR8ugh8dDGKdUq/1uHEMIcxaOgBIKQil9Be1vKfnjTZ
KzP+qsMOP7rhCyPXV6pVcvCf/7i8oQFjYoEEi12lSPCtHtlS6INGzXifTatq6HTzQetdt3iHjzGH
crPe8/Pr2xFuO9omV5bWF+d74O9GMJ4OYwF2+IJme2WmqdiS3eSVxCreJnlvRKOI49wRO3QZcQqj
jV6wrHffk8buKKKSi2NI1TKU2+n7BsrEsrjpljxsMXUhSb2d6b5xNPoF3fovaG/7J+fp6ONjAx5L
DlLGSzsSVJbN/8d80ePbQdo3tdMZxmDY5aFiBgao40x9/w+F9kgPnkzAzlNhjGltjlcPQrMkt5TZ
dYiMf4HGtj5CZprIArVPix4nMry2bxJn2TWLcUY3oSVevpfpCm0ShZbieG72NTdoMpk/O1iRa9M2
bmq1KeD1TN7zutW6PxubDvRvToG0TQfiPrTVgnKhbHKEQ6HAyIb5hF8B14fIJkmQK9okdxC840AY
NSZPT5eDeoF2/jWAOq59ju+uon5CsiPsrh87XYRzH20fxRX044z7d8zgd4e6pe1hsZyxIWQKNGB7
8jdqtpZ8xyDb7/Vun/1bDpMaLGuyyhWs/uPoqWpq4S7o6A/MNLWPJXF3QIazzYA1EvrlHEbZkd6G
Tx8KhlkvqiqIfBwZvz83hLAsIBoGomTxviYOmog8wAG2RW2KO0canC2Ngkxl6TX4df5cAzAoS0VQ
uMHL6O+wvJtgq/x98k7N08T310iqW3NuSTeKZIWyT31Z2IfhlpU0oH5PipzwuvqZlV64a4uwN9SW
h4EIYidW5IWEheRRc0LLgjyLkfYxvviMzIbdTSAVJIH3VmuwumwK3SIu3nyfmUCgPOlcmHxyvoev
q+0pdXp9kr251dofWeKTY5l+NaJZ1Khv/jdycDYYBbrOduPlSAOygTVlB0UvB4W2FRCSYPJ7Ntl9
cMlAvEnecDHbjGogmdNpwNfIGit8PqZovSjaKROYXm1pzAeOWanXMZffcW9735/XRYJKzHwHcXCy
uSO38Ob39yojnkdW20+79VklboKWa1pqTKEu8xcWirWTjV95cwRVc5v2mQSIx3XIyWABfBsU09sR
6TtsoX0FY8MsRZ5BPoCsQgs1cqkxFipNAqk/pSNIfKpbjcSEpQ5oP763J9fuEppj75PfO5gh3eSo
P/SFB9Zy1JUNCm8uPXZJDrPeThYV9YkuHq5GIy4GMAW1GVhGTPBovrdq42aOt2aIi2Q9QX60dVjN
Q258y0Bkswk4QuAjOVYfdbNu6/gtLESyFA5VSvVdoLEixXUhndr9VuP9H5sCTfscybr5bInzffRx
MFONpulB/kGNZbAiWKS4ToTbtqBeR5Eb+YF3jo7x9TtYUo1Ps1fJc+Wa0iS2AVfd68gP88vFFpZQ
ABzgJhZTjk/GiHPXfumSqhFk3YOgnaqmRRitln84bLU4hTx9MydOe/m8xndGp9Sjvue8kPSH388S
55JHRRiyvWSCbihJ4L/xsNS5AnJVQXuUTuytp67Y4zoN63d8lqjnZHzBjzilVEv+Z7MYFsUj42uf
bHRyZHLU41pNzxXQTK7ECpv2x7wx6VR3YARUUwyvvKQbSFmNybeuedP0InM2J41y2VON4xn7CaNr
WlMfLhZI2rJDM6Yxl8plUlmQcNrDD6KsXFxjNZOZOjrOl96ABccKYCmCrTVGYyMhTSoscbAAPSuL
hmMpZRbGgogtunharlDUPcKVH5Eqrg7R6o0AjeVz8EVGna6lcFjsANI8p9Oh2HfBdS+JfveXQAvn
s8MkGc2yx4KJQ0G5INo/n5onAW4tiPbxzbZ4U0mvtATAK9fC3acAVjG27H/zzA68pVqYc93dnH2o
9XXHTDwCErvM0ZYi0ZamvxPdnYD54/WmOLgspa96Xm4h5hyCmHGZor7gQSjJTh/FzsEsJfKSOrvt
tqw5o5R+mTtX9VJn26Z2Vjo3fb0k15S0pzJyKr8LO9TQmNifhOC2S9jtwuaiJ3eAgv33jvK69MUK
9xe/ULFfPmn5gHtGJn+FKexhxxbBTD9+NUo0HujrHWlYOhU0sTHBye1Wb7XyDwfWSJXBoxiypUKp
5Dd2Fs7ImmeEOnbXGDrUHBkQszfIeOG36vo/HTD3WzDr17RY5FpGN+3YSnYbft2BXVTHXmBFfVmd
4E8aP1HV7jHas7lKqbsKlOqw3vfOTJosH2vmeXaq+a6eOlxnAChAl5khiordI5JG4cBDwKe6rUR6
QFJBpfa1S/+50yz5fuh9Nv/kwSfbGSpHkVp6sQvygUccnr/gl3O48SVLnOtsT7CPvr02FLKiRyOu
ODNeLwtXNGLdUqvpWUel1j+X1mpZ6gMqIcka49vt0VRr5n621CONIsAnsxWseNc7NoYqkw0e3KkG
KIP/Siiu16RQqSiAisBP4FYlr22EPYar6wF4753EWnpfGd7+i9pApw7fFQv/OKaKHr+qKBJTxfHr
W+HobEzUyuiJelnzThnthIouqSUXszi6A48Z83bXVl8OjkJzqz0BZFpYkzRB+V/5sG+Ff0CdzCXW
VhTPsDlyVcAAccTdq8R7xs6N5Vwh0hekPouVKC6s5bVFt10tkIkLMMoSxIK82Dt4qLlCbDBBF9h0
A79vIbv6wYdVyMnv+ilL0tBGQq1ba5AqvE2WQeuWgId4JwUOBBNcCO4lVa5RukOoTuN5/otr9vzA
HINzg13f/zVlCS/Gtu27WxZiGbEchcY4l/S7QfYFN0Fu1PeYdoaR5jA5Hv6w84OscH6f6KQI3obg
m3rwihPdeajOh9bPtKGX1zMkFQvsKHaBWMnS2OIfAjkw5y+eEuaDFB44U7sD82j+oE10Xt0LQuNC
hlqQ60AkN5LuSI3YxPJJ7XOChiiC3WfH1lUwCMoweBzbl7WkRZQnHtZiOdEd8CbiLbXtRGWVChIA
TbD0sBzdtNOmiY+Qwl1yumj+MWOZylWY4gFUPcjxaR3asr+9pWaD0uGyTCSEdEfp6tYM+dfcg8nL
6YYPvgQiVDRCCDS6a/5SSdKQGZk331UVIdLbJJDEZ8L2BR0Pg7HKukd0IhkDdv1iTNy0aPinpuMR
3C1t0cSBu3Dg9L4Vf+GlBq4Q9HuO/00m3fmI+p5AUMmcjL2KsgKQpmnphZ7CKK5xIlC8c/2mh7ZB
kuQya7B9+NWz9KKzPocPr+1afH7U4DT+MMSdS+I3S9HJflyvOaYReUGTKQdsiFteAVGRTfq6fEMQ
nZeJHH1kTObEF6saxO8Lro0bNk5Vkp55+hOpRUnr66cJvbud76U/xWAdxMv6Dnc1rp8vVLivEiiH
KWC1391AXES4VWF0WOzCNMHwHSMY81726x8tPBiunewwvevJqX5FdfJ45fR6jYJ8sjExZ0wiKjtu
R6HtGrQCUsHYoju5syw1FMnGNkZW7dv1vJ39Ow8eoP5+kqna5+UeNLdV2LZNLvakKfGXETfm3UfC
UY+h2WF4iFiw2wmFQw0N0Merd89GBDccRUzt9Fj1Tca3wszB4jdhzOfHoqPq0MLaafe0Ien2hLGF
bgq8vR9bD26ngjS69Pv0z4rQv5JbL5DNRKYPhHtot/fBpuwnrKPMfzMA23bQ3CBDrkLQVipPL1n3
XlQ56E7uIfKE2S1uo6psPFcp/KXVr9Qiljlb6FELiN8mPGBe+L6CGTjsQoOwiHnWgodI2hp0RasX
GnF+PYFg8+YsnNj74QrroYo4L9xWGTRZRX9GOlzCTFZCQGo6HtT0WF0TW5GHLMnM4MQBqACLwNqf
DHVVUlOnHNLYzTK+IDH0R1015aEoQsdrIwONU+NTDaO5tlEm2RX6r9cxHUicRgLfYPipKJK/mP9Z
2ePDcoiLvqHdrJ8X5DF/bBziN0pNEj0dYe6Znt6ZT64Jw6B98qzyJHvDKSkfTpBVlacBM9wOLgZx
AFyUyKZn2FIcZJFqozF5KB9Q8A8DBWyAESAdby35vzp+ziIr5advBuhEtjX4/dqGR5Igb6Y3Zoj8
FNLdg+kHk+4rCDtolSLBR4cYEOTMyLXV67UZgYP17NjlTW4TfbLv+JmVvuwSTMB/uM477Xn/IPGo
2aVu9tsvnwkmqAaNwL8gQVFkoK8b0jSdCcdzgmOyl7jhnydwi8KS8vpqVqQxZHxadgwxcB9X2ca/
fGvTQH+Drug4mDEzJKO+Ky81Z21PphYVO2p5zycY8VRiDicMxdapueWLruS6KzNfKv57ZMspF4FY
PgFWmJYDOuyiGskBzb7D2rKeYI5zDMiwcUWJ/iUDHII0bzDyv0t6+fihcpIWEV7MoTrWk874gSSV
qknxAQFY/E2blKv3/QCPjo8BbAcvzDTBPG1FHS/4P0fMLTth+1CyGNU6WLNGzvy6Hcj672CFE5en
Rj/fHNhk4pyAOa6zDCdCUGFYqffr9Af1OS8YyzxRd+3Pjgw+nIQiQ0jIWklE3Ni3esOp5c6Jyw4B
C5nj2JsWm7ejVpJ1B/KbJiR6oN9fm1f7ijuSNpLkkaz4gAdWusPLZq343/txnNB0D6t7Xg++piil
slUTi3vqnqKrY8qKKBdGY/+GcpnzEKnVaeHr1f467XyK/gkK8CNR+k2UAehsTrH0GvRPRDikUlBp
8gquiGVpVLVMp2+krocIqpQKh2a0sCQAilkoMVgk2B3ERj0nAQemVAwQPA6yPD7/+B96a0frqy8+
IiY7s/l409ztOj5hvX80NUtV2JCez4Dt+2nVIVQ9q/mB9icdiV9qdgkjAMpJitBPt/mYUN6uY/8G
co3/P0r8DpW1VNPDwMQSgaL/zqTQwW+QJAp3SQbtzf/hkgdYN2+tOiTeqs+3x+J8MrinWUBPc1+Q
MC4HL7/xfoz1FACRSgqAmUhiKVl8T58Op/DqXIOvogmaEjfaVL5PZ41yijLFglz5lnEQIBUBPDJj
hgibFXkko4ITp5S47pdcUfXQOVtgPsG2lN2hagzB1eecL3VNNBHdjvl/EdBRxhD56246D9amLL07
ihnVVVk7q1wZ3ZvZka5tOyt9R1gEE/M6cnBrhy+UioPD1fW9TpQWK6hBFjEsHdJ+oAN8uIK800Vy
krLmh1DSzavw4V2/EzQ4OiFDAVr/xIfS4TV3mqVM4AXFK29pZ93yNv2HLhaYmWz+R178IM3amFkg
MGyq5woJtdw8ilwT/EW813NS51LE9GaHvYAPaVfuopMCqFRPbZNxoxKpo3A33jV2VRgqZw7lQRNv
kHnj9LJSobyvvjlZq4YsMVgE+IEhZRfVLVDGJGoqP9qrIvz1lGt29/zx8p8LL0RlNwN0dH0R48K2
sYdIVPCGLV4wDJShEftNm6UZ6mBYqy73KTGdR5c4r+iFEsAIRZX7YOGtaMo/LdDxKWWhgryYJFJ7
a1cQSrDYTUbWDXaQc3WlOuxWjCX/dOEI9g7dXblyE0vLECZCF1sOnJG6QgHUextgAUB6gQI8ueT/
ixtqgT+6dEqwWkCVBVyvwC2dgCEWSfjZZNnJSLGxdYOHb7R/RcqYQp8/9M/bJyB3D/pV+yNNdglQ
hmHMNtPjcQ8YculR5UZFPIFBcKEi4a6+Q72ohV2I6clA2ofeUvJPPATIJNwxa7ZXzBECSK8Nt6bF
LjCECC894HkI1/pFwrUeDv56M4vzGzdi/l3Vc/jpOsBBCAXQTt6P/aiMlMs+mpVjPd7J1Ip9BPaB
0GXy57R0/NJkRlt3juX51MOF647xA+OidxbRQ+m5YkoWr0bRGm1QxuTbw03oFl6W83x24RWivRHI
/ehWMOayCDM+iGkAx/S/Taq33DTtx9Ub+Y+fWAOB85HoJ7Ijopw/WpTi7qnmYBgv4KeRUdI9UD3G
dSag1otsz9DtENuAMrUIUQn7M9ac3kQcbvKLkkKuvtF1synyb/XAFcb1iwIcFwxdwNmNV0BqInqz
SK1YHhLbWQ0OHFQg14phYSEi+nejhrBvoGLpzICU1Od/k2lVGAqNUQyr6KT1LURo0fKtIVFxv1FL
LBOPY2H18iAt78+oHhkLobQmk0Id3nmvdKfV9XWoecO7BDWy8wsadQ46XiTj5ShuGu+Leu3+8QKx
BylmYAVatHvlsfaH3tSV7FRJ+B7qbKDnsAVYsU6UvtheJZ3TJ1pcW9eOrxwv13HqUVVyrztJeICg
LWRHb1fp44A2nU4CbKbs4WTOWhSeRwyx/6ob5B8g4pyLYvum3gb9ucYcHMyAv4N45y9NE8X1GxTM
2DU5Id1QwBCfOsPqvlyEGTis6PMrOaIrNCTC2MxlSM/9tE8F56sOc2JgKoMO7aAQXPN23dmZ2UKq
ytkThT6eQLT9d/TpdqjeMYa1jwXSf4a29iIR28wroBv87BH8Zs93V2VgzxZmspE18yUl5ijlgWly
/GM0jE6yiJZx7xHzyFe0ZET/W7xfT5BJVoMrjt+2q5JvBB6okQcdutYoenMkty//aYf27A8/xwrT
vINBgmu+6I4Oc3FWCTB2AfUS9jTdzJFhYCj74K4bmCvQ2ReBUHwLPOGAyMQCNXFahQDxrZYHQnV7
A1hpEtWqHfoLr2DXfNB/8nxg/sBAeNgAOeKJUHtfxfrjqbCKTYN9rd9/PwxhAyhn1GFYud67DgXj
bYxHw+N32h7CH+P9egQZ+Zf8nvtez8L1uQ9NpCE1s+BxXXYIqL+qk2Jl0unb8F+wKipjqiUdY0Wk
Na5gygiG/5eFs7qWF/GMdYXrZs+ExC5pzQik+0lEEIKZEsQtX9ZKTueCo9AUK/WEU+KN5xypwMua
iRlu+SW0D1kEMlJExVvLETNVODfkzxFtQZy9VtFlaRRDRtslptBY7yC8Gm7SHUhLIniofrKYpVyz
v/KZEc0ZpLaxZ2gy6bKQO8Kx5xl2yAaNLYYrco8aK0QQsGxlGpPrpjcujqZeFFhHGc7i8FSnLXM0
SpAqnr9Dyk+Di5VxKzjQEPXYc7q5rlXLil6yUBFp1FyusoDcAkRMXFspYfbMRH0Ld4EXupDzC4IX
PlsDtPoZDThhm2//46mf/BLn6anwv0iwhM7knFXXIwzJ26s0I/gbD2SfaX+djpZ4+8BncsbKmz0F
bPiXc4n4AQ+Gk7LsXSRkEhA06Xs9c/xh/J3byapW+1icPr1enCFFPpfjBws3/s3RH8cCZuHtxOm9
suT85Uj5s65eJ9K3zEifYvI42Dx4Gh17oqOmHtcOLzCyWXBgePvCY9VOhnkSmZvubzxcf3cdmvMg
L/c92nVKHYQMqL2kSLVBwK56nmGuANtX/jtfx8P+F2DNngY3a2GOdW55GpbnfsrApFt+EGAOUM0I
2w2c7d8aSyd/w4Y2NiMHtKhVY+sDk/KsmC8x5UCCFxa7cFKRZvNPW3fC9Hf6ZXPaRMA1lTbkTcNW
fkveWpsjkGoEMPenpdf6vj2dB/rsyWPSnBC8uCY8+W5tfU/x24+TKOHJVu4SYv+YwYQZhYI4QgPN
VQ/laZJZ90Upi0KcCprFUFKIJio0U89kGac7dNweez4KZSPVHP7KTjTE3kcNMdzaStn7EMR3G1zJ
FaZaqIp2/DFh+xy2VukUJ+63J4BuDzopfK60NngOM7swMhimf1reYblWJ+wNfVqeOhy5uXc4Kaff
fq1J+f/1vQOrcosD0GsCbkdlSS8xvtlFbjIZttWKWPeJWRAQgEDdjsHHmuZ08okH0pwuR4YQ/1GL
+W7AErMjkbPsBhiF5Ct83ec9fRGdQ8KcfeaUhcL2gwUitn+4K6XwD2xoLutoR4iVKrmgfXuiRHXA
rwHtfLpUFu0eZSt5Q+blb2/HtbIIPntsjS71KpnYfHOn0BXfQdNk0Pobb5Mn0C6WA/Y4ZaegFVTA
aJM1/TjD9pO1OvNuTq5eCQGGJHHbCx1fU7WVSaK+BlYUk6l6p8pF4QY3Fscj6+73Swc2KPbOIMia
wBUAKtpQtOcXQR9Lh4Abdu8LeMSaIIRYuPTe9OCcZF2jFxoEiFum5ZPnWLHzP1/qAaVeJdywJ7xw
OWQFaG4epzQnlND+VFA21DIV7A1nItgBXK7vHhdjekQEuR4GHrlh0VDqdZ336dJQ5+u+rJO4D6rZ
9MMtsJDCn6DQMR6ATSUhAJYVQqnwurQMQa4tolPDw2RBygX7a7jlYbazJf0X5WVpsxUYgmvI9ybT
abFhip+qOYlCBB8GxC3KRrbpyISvdac++17XoKgJTOXorNbY/TWcpnONlLgWqy8kZawuylA11fwC
50CoaDDQr4hQslF5eLgJqkE66eOEi1Lv/p9c5lC6K5R3+iouMbv/vfji8Beu4UZ9uD4WyaPpNtiO
9rDCncuxZ0m0NNc8kz8UVYycBkqfXfRYHSyhL0DIP/LG4ZS0SodIcU9YTKnQwsrymMsnVJsI/vVC
kwgDqv/qRW7q88KGbPyenzf37W0Xy9tCW546M5RFbB3H3H4osuJ4JMUSQE2m4YQ1mHgqKjClj8VX
RmFnP/RlHMPFwQx6BKDDMFTCnsqntItYdJiKnb7QKo2MBc+mPsidmZq7VoK9I10Ie2gKqudickqj
gLceVrZrjHKe9HX0g1cWDzH+izKyU4n3KPQ1SGtaH9KSvfF/6Pua9bztwdBmcQgrrPvCw5swLhAc
3/I3715REOcm+KtJ7AxOUUPOyzDP5CGd13rwWkz7MkvN5PmFNRno+b08B+sUkItCzfInY3KRd5pU
BXlcKjzmZKJ8/aNtHUUq8raZswXMU3/LimOTOCyG3OSNt57CSA3dFUzybx253mZ6clMQUMmtdDtj
CuhP37E9/e66H/hRMm75HA43pDVTWAHQFsCDto6L1SQeNqFf+/+LVLnthdBp5srZK2UrlkT2PCej
9Z36RjMngA2Gu+wK/OkAhIbSvDiA+GfV9TpiBnUEmzlHwv2EzQ3U//20gr973qKRVX/1LJ+yGSYx
Gy91xC1dLpTp5Wwa3x8qO7Uj4XY/DMdbPTWuSzSrGxjxb9phJAtP9kmG2fYnAFBEpYuyT9CYnY6G
l70s/qXFRQ4NJFNiNHueR5BcO2g3e0CdIQ6GetjOqH82X689ZzoaW5GJRtzF+Ms85Dcc/aCII56M
MhU6RhRW59fqAF280Ve2EMzGdetsh1AwiG1axpIOlRsCs7gG+EqsFi4bO/nHikm3fwIhX6Qtc4Xc
RB2ZWamWFwLOGbCPhZj3kVS1AgSjEb2Fx/tLqr63qDuyIFsRaX8A/uLT9EB8HxuwhVX/np3gzEXy
Ioa8oTpifk1x+vuHUxqQkc0SUIXBwQOWvErAj5ouPhCjQLQnpnMJMJjhMzChJHjAJRfQICeLXfJJ
3/6saF7KwnjQfrbKQupPHB+wpVtMMRbyvOlLQWrbeL76lWEcxLcK7ScIZRxLHV44nZ/o05ecQSGI
FOjuQi70zQ1feJx/BONrDWH7REXm23RZz/2aKL5AhMvR1/E9bXOqtWi/YjcTV2xmTH0krsY4izz7
hoi83crK4LfaFhF6axw6YT4PvQcmLD1uXOlyrSOsLzpYBxcaH2Qnk2CMwTznYlFJeJ7+v69CKGIF
l6jPjwSP2OLwQ55xPMJ2dlu/j3Gje0RbONms7s2Tx8xLosa0AnUFEu7UByASvq8tkhBN9vqDAS+E
XD1DmNRN7iQ1IEsmVAOF81UuPUS6VAM1sYFvdO2U11R+6XHWCK/29XkvXteUpBqeProXGJ8kDt5Q
o0xiPBYDabINZfEJg0f5LB3pfYkJ6l7I1q0NdbTMF6CSfwAiI4qnv5JaQ6e9wC77Fd2d5faMDXlA
bm/AZQ+A7p70KfC+LMbbGXU7Q/CZ4DqilwtCE71PfMQyxVvEi61xYhpLydUb7mIWYzl2y/nBLxGE
TIzBWcIytYRQ7rXb0Zld5p6rrYiv/SIGr3UILXO0DEnnKEJ7aMQ9DgVWZzW5W6WF08sj4pSJL3Jq
Kpx+n50albDp/CyPyzGItRQZV4MqtjyOzz+hxFJBeQB630owJYn1bWp/F6zOYFXjRqK0gPEVXQys
FyQFAH+3r1UJlc6+jCjfsnDjFRw4HeXLu3moBmlo8SZTPsJcOtwsZzpA1XrV8ZzHjk3UkKuXJKam
xY0D3P41Fn5obXT7AR3Kd90Gy7VU9Z8H2C0LK8FHz6FjNnPcqGpxIuLlyIbBJeBrEtf8+uPVWTnx
7NcdRoH7TI1HOTqV3HeB7n+O/epFUpGRwPC6gQwVTTHpnbSjxz/9VMgRz9zX8Fpe0cey+H13f5Xk
BkO95FeUEtutEV7xQMC3gKltwQBg5NIvGJEsMJLY8Uzm4Wyvs1cn2GTvhqBjTC5tgbbUp9z+g109
zO+6Z1FizfjsVT1bNRYx3T92Pz6OLiGwJFrx3cfAjxj21MDX738A+BTfXPIi6iegp9aane4IstMT
I+7ECI/RLFR53lXhJZZvx5i7Uo9V4YVGoGuEF7CFlMnd5sEfynhLOoRKMl5LqwmtM0a2LCvWbO9Y
JuINT8ofhM2k9xNwRHhb/Wd4NSwlw1SNPDPjOaoKWwSuRjVyrgFWBxLSWf4Dzuwu4tD0Rsw3osaZ
baSMjITNOXxbgR4mbvoQcXXjg8Ut9i27odWkLs8n4Dze+IDSYTSYwx/XwGaJr0iJf4VhYqAOiKdX
XibUns35T5/l/lCG5A9cimxb99Vu1Th1YC3PwB2kO2nZqLSvYzN2oABr1o1eRdNrnl7t7q8qO5iV
YMA/QxP2Bh/WcGa0SO+ad2Yc6MGynKY/3K9b3p/6uQ36wN5OPBiX37pVT1Db7XP6zgQGP1febbUS
+ZnFRViKCJRXDCLfJxwbRaVbTNXqyCFV0RaRJ2pBAVxmkFLyzrDBAbQwSNmpuGhYQ+4kFG/c1XJM
5wwNuCS7m22xx3NxwvAnXQbwpmgWut4qJ5S9WwOmULXduu88FL4sPgprWkjySOcDD8Kx+SaJ80tZ
31qUh/5i8gMsLZdf9cTpT2KsKSkOjXiKZTwDCb3PBJp0RuOGibpDogj9YoI0+LXwXk6sIDYFYmjF
3pQUZNkIGjf+d6YUgTGnPNP9vm25QFN2iRSD3xuZXd+BN7p+42qtbhOIyCz2wWCCg4oREPDYQaen
XCtmIYtFYi9Wf8c3kO+OD4bXZIjYtju5ETU4cefHsHMRIw+CiJwCtfYGcLUudmLuuk6sYn+mTeJN
YRG5I+nH7Yh5Dn+A9Dk50UU8RlskRS6f0X/1gcw5l+1kHifAx6DBpS9HqYda6ACfzRelbFN9JgZg
k+xXQApoZp7NF+R1pR29Z5Qs55/Vs9hSnBgGXeNVbKDuIKxM4hx4iWTpdVWT8DSyr2+JvofzJXBB
PEHbPAgBRbkBhdxPq9N8d6A4R0egHrkxNP2ukYmmH/ZB3AYchIm3W/5xZtM/Uyjsd/ALJQJIXSha
uLD80lVemqYtVIN/Osm+rBmfrQMshG+jjYGNRb/VfTxbFtmGUhkZZj9ZqkCQL7PpU+9QnYZgYHKk
rDacI5WV+0y/h1J1mfv9jdpQuFUSUHfuk5feJyQ8NJdqF4VCHD1WZMgNCNM/cb3xSN5P9vr/Il7a
INXabvw+EoLzSMyaTFsdSEGG5WSDQUd/NTLbvOI7hlTNgUg/ioSIykAr4a4+3k4sUxxmMpvKDexc
bIHEGHVoF5T3vn0aBZ26NY7xgje2dwA0n/eJVGdO6meJ4ZkoP2mfy3XVqQTi8OYbkmLbjmp8yghZ
WuyZgOLkimoG/kHcmvqxO82i3h7TXMrDv4qMHqfjnt+FML/n2AXB6VbHDk/A4NrCUpfyUxeMiy16
HjDkNzQs/L8ZG+mk9i2IyndomgsirbscmpF5NIoEoGPQaeDJH24+qfuDOD6zZfRhNpUpX9CGvg1/
NiUFYZy8IYgkNbj61v7w3qq1GYWx69JUZYma9CPzZOufZ9XC5bWqsABI7yvWGzlhDwWAyUXZU4M9
qoBde14LOS+dbBMDuSkyr+dK98TsJPqvV40Ry3zWUDcyRwMJeybeybIdHcGSsCsJ7WP/e1KIBKTj
oN7Gr/ju5WtZ+0bd5W3iqCNZJ68VFYWuoEru83RqQMGhvQqtVNXvC9F8Jm/CUo2quwoViuAha5o0
DAj0lgOMViMl5gCWZ3m57oML7Jl+2NN+0xgbKjT/npJm6H15F9H+d3cM6qDAbnQnoFOhNHValy1A
EsS+R7VIAj55MCL9wBhyo/aTJVv98epX3t+psSbkWuwnzYd2nCU2u0gai7GqwVmBKNW1lbacjwGP
xAZgIE5WCAw2yXq9WT+Ug+5pUg6ZJLKUObJJWybfl2yYjMZNHgUI2649h5Cxk1fMUbI2H8nbIdkm
j6CXOMktJ097pLJSFkmjRi6lR5YesHfyoI9YFsyApnXG95KmPVhGJhsO25ILyxAVNGoJrGXM0xBp
OHAoUNruHQ+i32wTHCJmvmMptUDQnkeOhwmFcnJ1+7p01u9Rh29AhTrazw2cMbtmJAmkSjhMuEK4
77FsVd+3gO+1jFyzzFMR415a4msNLL0eJFYokNWxExm+MuWKHJEUOx35HyDIjGbmJebA09xhnTez
cewFz74Kj7OeCLeW4UwmEcyCHfZVcr/8hVJFmiWlgMGdETMby68YlcXVzLOiYsyHfdOdiZ6fuvH8
gSHYjBNEoejGs1DEKdCMZQ/GnDUkaI9okN/+egHz5j4I5KRpbhgj/1doMwQjPEOzG+8OeESMKNhA
IR3V2i/pHqIUPV75AwVrJWv4lzIwys35IIzpfHJuVE+YrmRw8hEyMkizpo8Z34FEp1szg71M8nIs
gGBzVPXiNd90OqR20fB8GIdFbjMrgq/t8gh9H1PaeDfoFHy+UXzwHYmkB8Q/ohzhSNXo/In/mI5b
3T121I92lqlYd4wrVgccADvPt5uPB2GQejEvsZDS4+17O6dd25ddRABP2hZtETXrGHhY4vucf25U
UDIjxyj4qbEvACFBBw9kQTPOdh1z4JEi2Iyw6O38hxqgvK/ip34Wc5esaMaKZPd+bBeFCz4rlaLn
Eqbhi450WKtgQQtCu2ieQYCb43Spz5g6fEMP/xWqHhmjStiqtdK3+8SHYM/4RiijmjeqdLrekmhv
gO+BSMitmiCP5x1n1w7j0D5A1R4T3TcjrpPqXaKKL5wZGWxL3VGTe3XjAqbyiaW8mkhNA3vZCgti
NX9K8KyqBU0vIoiwyUDZqZp/JBuc7+qnOtgbFWvccxmsf+USAYfn9kPIEeBTgKWfqNoawHqRZ6Iq
cPoRKXwHacxRVeY9tbSVX86oaZ1j5gZ6K7DnlslDjLESjfYKitGrJDNGLqy086+IUennnEwF1MdA
b3N/rQfwDyusEHUmkBJPpN/h2bjWJz/ZqzIrlTn5NOudwP/0CgFOXVbIDK+l/kAw/gMviMyxTvK8
MzJjP7y1yci/JL0jhrxw7Ys4Jk4r4RyaBnOBclRnioEVIirSP4v4o10O6S954zTXxDQhtT+Okl1Y
a9FmC2avCwcbPCs9OfaQ2gVJyhXO/f22E6LgpdA6elgsKFz2esf2KoRg6c7ust5WoVBmHY+0RYcU
DXkOWBAiPFWOJ1f/HyM4xNvqlfmQptelgw6A86JXrvO3yrzHuuwIXVUB+zf5nzDTAIXPVwB8ET7S
4flTy5KXUNUua4F1NYQhqZneFoFNXMZjydTyC25+E10S8tW924TJVOnF/88AqVLhinfV6LDVx622
s+ajlIdLWaC70cUukZd4eA2JojVTJZF1tKK8j4n8L1CP4VIdiOrcgAjdGelza0jKxTMSh3zl3UYI
PPkgi/IMTqi9piKEvAbD5yIh9hrUIQXHb1BO+0/Q9NsainopH9a93tR8d5JAGqKW0ulv4NHulzas
rqE849xjsjNbyJ0UvYYDXfz9I00wurcv6qgdsDKnapqxUTEjOnlG8mXTJNPl1+0ggkou0YSRftED
A5soRghvLb32Dz25vgCOVxDP+NY8uZwLDshFTyPmaA6nm67lR86RO8ALcNTiPZn9gIEIplWTIjqr
LQKUBGl6l4TDE+Mm258yPGaj2d3PoWY2YO3zoGsROvvN1zOlsJ5a2XdzaGaFgC03k4AM9H/63eHr
JWEDKO28wThqEV7sjrQmjSRsfF7VdSJ5z/osCd+RhG2h7qJeC/zfb+Ag7fhSupr1EhpgmAPQtMhS
lBOwm+Vwgki/cV9qhb7A8hsfw6i3w6kp+3vvB3Kq/xeXOCvs/Rtdd1dOtH0Kou1RhwQSVrgoASuO
g0bRwnFb8r/VWHnvtpEXXyDMb82s1p79qdU9r1U/EVK0JYZxh6IKcEwtpH+x+2sRqgT4yD6/dwYn
lotoTfgVJx/wCX5D1O+6kfIxKKLHKngggkl+CC5Z7t4yRmiSMaXAoM2aXj2xm6XYlXFdejaRqsXK
4LNzx97kfs4IkR1uTadbvt9v4ZP6XDKDxkyBd4cJxlYWxOl2NG1ZwzBV7mGB5bjSsrlBgV3RvItT
CXLvOMb4H+QlZExLnz1PkhNeg+WWA+Gl97n+7f7pI6+HWl1vF5W7KffvNLMvrihurG6OZPwGNgz/
Gj7cvM9dtur9fAImDbRfxY4l//jRW7kGpY8MMJIQSJY2JaiMt3Eyc9fBl/yfeZt7TjFyfdyWyfwl
h7F3hpZWrGKHa3ItSPGHfNzCDMLrz26A2fHZ7scOWBey6AVynD1+W20sd8p3fRiC2ycrqkVa0lMx
+c9nTSjHNtEOWoTkUyxAWhlPAaL1Al1DDJ6xNpYdJwF35u9HR01qE7ALO+Wi/Y6bNz43t3GRzbUy
ydmWuDGOVZ5yJSjstleVWOplAU0mSyyCMAzATMTd3fcxG3MJINATuTA9DkYa/7bHwmqi/WaNuIin
0NiNefj1D7bAhZ05+w+33fjjA6znEap9+huEWU0VF8xyuWUzYDbePzw5oNeva45fwysEfU/W4j5Z
43emX32zkdDreJWcZA4n08RqKt4FyokG6WQwH9/5q4Hpmb+0utOKXroFiTjx6JzTE9CUKw0YOhGd
Hb4iELAyec7g2TBTXOjafDw0VYscK96ylOovhQ4p6GDCbZeT//0W8802aFau7eS750ExDL7sjTIW
0ke822DwOhlTBZ/TmM84xBOD5MdWJ7T1G+ZgSKXtY+DvT/ZKzBDqNsR1Hcy0Unwc+LMDHy9AycK6
tv64hi1nptCVZ9T21Z65nQcdsKGGwdYlOi5hsgELJ6wCdonjZ7NJ5SAr76iX7zmLWL0NoDSyFsEP
+yUjn5mnFDh+f0Kc+iZeGwAgeEh/niFNXwciZJCz892q5nlNppLryFZb2WALpkh+XvVvH46gDcGq
gzN2evHvMKSEQoxKlimFI+Fu3kMVzerwx4NRYjscoyW+RG4HoJM/SFjsfSVI014m11hzpPxmmRy1
JKdoQsz16rXgpmMJPdp1c5Vzs+4K4l2GkV4jJiZ9BlWtU6MK93mfHlCnzHAOYWCuINmCfJGye9jC
GcuTlfw1tv37Ki3VnkSrGMQmrqQTaQLSvieyQmcKPBmKwTsL9WFdjdcKxFj/7ilMK1qLlXnlPNas
PGtdzRDsQ2MCZlVSRV27lT9B6+unJJ/2cecog8s4S8yhSWmhiSJE57aVSIQmIb55JXp9gz7XErjK
F2DlPtUQs6Lpf8646dt/wMfHnalytIk4iSt4uPFZbNMgkxsXb+jOiGjZy9Bq2EsmSMbuyathIdbV
hw9MOZ5aooBerWtbxTQU2jDK1AF4xwFjTLwYNs9mUcfrkHQlg64PlOoEx2pdMFHo2pzwM+g8saSU
z36tuxo3zrSdwOxmy9hIHMmMqgKcXniQm4falBQvihn83DQpHfjgQChs/vgTzSELjTuL3gZoQist
T4EitBzHRLjzRElbcCBbPajCHemLttqCMz1BXW/7th6Bn9sXKcWx21OZChvGA+DCWya8egomP6Yt
4srOxKYyijVB28KlZPXAGh3M3mfDug0jv00qg0kSk4rYO97iT05HD/bIUV+kK9DisxtF62Y5vzll
NlYToi+HfwYzzYgkMvwZegq8Hk+lTFam6Gli7aSB2kJpK1Dl0eCFs2w8KuwvJ7SQURuxFfzR240E
4IfTJofVGq9IFEf30ZbWQKoJ5tco8Zm7X3yrUua76DI31bUOfOA2pbZP0phmOoYYtomwjUYmsFYo
LDQuCc37JwKa3Yi3fQZNTw+8BoYMMBmkjd7u6YHymyTooPU1AMjo/0BGPELKOvhGv2AC18IDeqsU
LKRaGT/7EnduCjuDpmY+/te4GYnxRJjpaRyutcxzujQwi/CF7YTboAvAUB7hnKl0km1gR7IdUeKI
ri6hDi1K9YMl4I31Q2zsdno9J0dxvQ7dGxi/Bxz/RqquOelLDvUzl8VP1GsUFCpGJaqyfrRukajz
tHEPCwuaGZbtiw8MyuOCg+i7Cnt0QJkWrsYlmSsRBYvM5rxMqxH9noagSEmUFmY5bwMkyLnJCCBj
/vXCK7dHkKX3RlzrA16ouqqAtNXXgjyy91I5G8gIfcIEwC9FhKaKP7fLwerxO4948my0cRSZVvEY
3xVpExC6lZeOzfFxCIfA1D3OhqlzHEain76ZfyrINX4mQXHrmTmeIxFfLr3F3QrdTpeXFM+bHaoJ
MrezIBuC+r55GFSIYbLmHfcQ25RT9fkDZ5xB6CorGptjGS4yj1q+GmPqG4Rci29VnR+soiDvaPEd
adgCjXPtEThK04orrqyFls9QmuALgTpSoIai6z7D2iyMAhFd/qz6BQLkX+kzKfIXa18X/GImPa35
fYL2PySICEvwDMG71C42Ettyr9UXHzdwBVthrllHLyM5XN5rytLvV99rYzLhxmPu0voulpFZR29j
E4/ILrDZayxuOlX53uWMiEX9qT7XHvtiBqF6/LW21VCCOrFcckRsaurr1zRtCKpsbcEG6LN8oDtZ
FNkH4g2yvxVG91NjQAoTdzHk1oHFPvlaIyjMWsd2VMochqpRYLnl6HMiHxZKedPMaX4F43AchTs5
8nrcFqrryr3XAkCe/rdVmQrFhV9tFM08aSyh/xjFRuv2y22ozCroFuFXDB1W2b1Cy/6pESxWRtlm
kSc3U6NND5wmN4vEeUuuJI070LlDzosCfOdOjupQM3cNhyxs+Rbf1TUf+myhyyEetZ6U0dtG6Vq2
5Mt6/RV+mTJswKiqcrnMpjZTS05x/pjuLwl3l663Qaw3orPjWHux8pA1a/xuLBg7TowO+/9pfCVt
pWcwtU78sItE2+BoO09VbPLRzZPuecguzjj9usFKg0Wuu/uJFClmA7am0gYHpNAVgPPriW9CX5C4
6bqeAYvR1QkO0bTVaS/ZZTwory53cLsEhUywRvkmlZVQ3S4bp7NypohWtYvweV23m8+bkhYsH2tf
KhKxYsdztZWMl9hHlHOfkj1Lqx9K4iWswA+QwYwJqLni9jpbNhaDbapPULgZed7nTVHV0AQs2GIj
aHPAho+GRP+YaJYUZ/XxfpKWUKZhNP2ujalFBs2YHPEJuYOEFGeTfdZEMCN5y0U0OKzvGBXImTcK
qVuhAzwmfBL81Mv2w7jALSgqlTV1oAoYlTy612L4gSflh91Ch6tWSOd5lOVNL0ds2mBIKzw780j7
6ea4HsG8m/JyeojPauE9e5pnRxsUt5pZ+qPDXcml9bEmVzf2Esy9ggxO6aBtqmSPz6CEUHHtm6/M
jwYTs2/0ScdHgJPjFJhyEWyBwtHRqgTNLJbvWJ3tf8c0t3y3ypKJF3DlspgUIL1LaxUizyY8KNaj
D1sX942tVZrHOYk9iIFgZHbDSyGkfKaHs/5B69dmmiDMMj21kUBZFgeUE9BWTqDuJOtmgMMp5fzO
KJzbbj1PDbcDhYu+HFPFuF5O4/k++IPkQ3OsnfamlukYRu75RufF3Km68rHsXamH9XneF7pd4EfK
XPm4Qbl67l5Vq/4Ui94MVqKIZ7B5j4IduL9k6BN0QQDXJRHhf2QsCr/xqj4RI+qQ1cDGz4uNCH2H
8d1Kmw09VWuHR43aG4MFBuAYFSiruRlr4cWSPB7jC1i8LeVuX7DmaS0FVuGZmihJsIMndVfyQVWT
+6126aIHx6QjjPceektNhJNC1IjjQPpGMhZyn9QetXEV6e1pXzco2M+XCtSEb9GFbpulsxSOvioF
qgszYGZsLhDIxHlNEHS9/lirFJoh5HtGUXiXyiZOQ3wNDQKe2eCydQB84dfptJg/TJE7d/FnwA78
2DNw/M1UyWg9GIiX+Bg+IoIYSMJrMUqHroBB6Tly4SY8oDBIJVgbEMtZtMKdl1d8aClPmQfKpkTI
F7yypEa7ow2aAsA08fvISecfAVj68kLU7igw1Bij9MY7NrBjUC5rT7RPHh29dbn51RJ7p3PFAExq
ugnTcRO9W/PbXwwMA6zvLNRBIUEEHqMTJiPH6oPsleAesveuMQn2npOpQu7D68QifIGUGoVbzvgw
GZQ/9hRU8m5agVFwWXbhkZtekdwKno/guthb/lZPbIE/7x9fWWEPz/YGRagxtSg+tvzNIpz7d0Kb
ZMz25LpXbe9Dx5hQ4T3y1544KPjcYBw0ZcXEGQHhRw4rkZcJZYPDLzu1+aCNadYDYTxF2bvT2I9k
GUK8AYH9bCLUuKLKQcVBiwv+AnnQZmDro7t9IK6OjCbx+UgWOKdrp5A6+Vu5Waxu8yW76QcRkfxR
g+jemxHZc9vJrL9TRG+RoQx+rDp3D8aTY+YP2KuC8XKczcarD96nJamAJbxzwtcN7nVNM2wdSZLS
ChWYXrmsUBM5gV+5X71DVwnooLulRWogIkfLjuEK+Y0EXf7Tb2SagjSVIHmj+yPU1wpbZA2Y4KMR
eHNd6heU47zZJ+sRWiM4vubR5+SaskBd972Oqnh/51k38YX1fRU+WlMMhQzE8fy9+k6I7Tzy+ul3
VmuFLFquvzlgruCiGlBMvtQWZFRkKk3KggPtBZrTEebdNV30KzWzUEnKqnR2eePKXHztSnEjgEUX
9yMIH7jpQWo29HAQU216EjGVx7QhpgLP+tMIZvxvWsWCPN2V9YuwYADtzuKOee4YhQnW+BNps7xX
a1lcZJJ5mHXMXjkXL0ted0Ubz7Ai5YlUp2jav1eDTvoWcKrLyjU3L9tf/rNggFDOMVanpoW4IpLJ
CGj8Vk+7NSwUY6vSRZMiwbqlKoCblGN71e8gX2c0BIf23x+l88Z7wTmeJGlpEDYqOQ4z90Yhx1Zn
tHeUHNWj47d0r6FYJvCD+868LRmwAetX1nNjnhkwRpKGtHg8tWWwVFmw5Hsu0Tcxf477gyC5szJn
zpIbwpc+G18xo8u0BT0dNRIJoiyxEbu0OMsdzM1OdfxJOQaU3am8925czyECghOUJsKgFaR8HRUB
9hX3t6RW1MLmjnMbJo+yJN+aXzrxxA0RBKj95zjlktGNG6miSYh+AAeGyk650CR1Rt1BQ49rO5TK
5etGXyIVPB3251hgJeBmrSDM7Aj+0hcXppAKIVMg++xwSV5Z/SfhCmkTCLtlsAlyjCei6CGPMHYB
xErmlIiHxnDGcJgb40PXJMIX6WQX88+bdl8pNsHw4gvPCw6tHzCodGy6u2X85x+mYkc2Qa/7scXf
aq9k9S76WvhDN5vZQNT66HVqlsOakHS6HZ8HUlRyIC4LrU/VO0hNtItR3vXOfbqW6NDj9XoY1sim
UxVTsxS6vwsYX+kaOkmLjkFpRSgCVsf40PAAtXqzd7b25YimUEEAFLojuuYbQM+fIRiNanG2iguX
wPdo3c6ca2XgI3VTsYL1hS+CchO1hnS0/x3yhULPe53oGC67b0Fc0RhKZevb1nhOXFTc7+vaI8Fr
OSufoD9XLYaXoUy6T4g2P62e9xlCKVevr8pR4EhVSg5vAJgNsxV2JS2Cf1ikwn3eVH+BnhlZsW31
nEbDCdcd53HFwlOPNuceshaB8wxFnnEtngyL4F0gtnvItpKRUE0DjITiWJVsIYXw9hKTxL14gXp6
kLmL7iYt/BO8P2W8gwx/4BYSpCFTxj/yCitpT+qx0llgViTGGHrrBaksX1MR+JC/JXueuKEdJOd5
WgnSyLhL4v00PQlJ4Q51O1wZxSNDRQxcF+RVUCT2VKjssw4vTH7PyYbpxwwJOlnCQc2qINLm/zi8
AW++l2buPD3TaQ1wRiYT8STPPPtg/43dBpXUfP7twqvTEfXqqSb3NptmWbclzNg7q3dzCvpuR23n
th8oSkcYiMc56rE7/uuwXHhjSLZSz0lNJ5EClCdyWQFGtX8GP8tz6lKZuOQzudx9SpTYpOVL+Isd
FnKn5dfVeC1ZreDUjlo5POF41q+w4DJNilpn6ssO+p8X3obN6tsEB/xurusTWZdgx/ex18+ZOBj+
7NS9ZPFMbNmjMzb+lnGPzeofZXNZwqzl0lePhBF7mApFz7fcIEXf7QJ8DvxEFQmG/s5Vt2+Lm6IS
DMZp75VOLdIFcFU9YPdK5oE8TA6eKbolXQV//aHRE6JtZw2zF8OMbCsHi2FKFKPc8U5XJ/xjUYSc
pr91hqfKuK2p68F79k7858DCxLyDtGxMl7iPU/lHHygFq6uTYYimJBHd57+RiXi1C/+OacygjDgK
VpcowYOtNFyn3LTXMCW2YWtIniqZjF2T+hCWyWCl/j82LaFZW10EOrMeQGkc+/lZ83symE5wEcX/
7DKe5MZXQdHUFxEKHYB+3pAxP/bl8vkW4OEQgVbV2UNZ3FM49SkYtRWxvgaBlPvw5KzuAwetNIRt
82xk/YpKR3yLPkotNOdr/hMAg3CHRnS6xR6AG7ABQOsO+ioOB1hbCIa35H/92euPAjGE+g8uSz9T
DF15Xvv2/M4E8kP4vr6Qb+tp1tl+S2dhSzH3z6v+3EO0wqaBpmbUyvqgFDANAt6UIOv27KKN9D1U
Ryifo89tu2Ese6WtOeGFu5sdiWvpNSAEPg+LcRIjlB+Wt6vw7NFp8orgzTEKjguaZ1QB7CXaSQfY
pxPNAsBlNopEQ3uHbLP7dmBWUvSwk3i6X0yXbzOWEIsuzMvU/kDkVFaPqMTR3Rb3UVEbla9Qkz2x
+bjPXq5e3AW9b4vov14lrf7AItdblPCy3mxhVo3SnkQlZEITEbyfGgR44mwDtz3Hhosp1JXNeZ3G
8n7PacgoPye5UQKYGPueD1cXnFIHur0d3iDsHta99TpmyeIC3rKzRwDKXAPLr5SjgA2wZV3TX5iA
0uxzt1sedL4k0bLlNwlaBSibgXGo3t3UlKklVQsEMTBV0woP+eJCSpS3MWlWDnjt2IGt/Jqx3NoQ
f2n3osCjIu9pzd1xiXstQFhbDqufcy6D83VoulMrtLlJU4UaEq6XrBeSfuwUiPiiiaucwtbBTlGn
bgwZ4O8fS9IVodlte5KF5wtYU9vvOMEJywErcCmRJ5Tx0rOgayS4+h4QT+A9eUIj+jq5wupp8t4g
owSnm8zkYFiyOrfW1Iw7LIlPw1vA7mznCk1B1w+BhjGrvWXXTyWXw3NP1C2/JDVvwJmXFTVxYSlE
ARa6VCAcnpskV/7EZeYRNFe2v8biHOpSNvhoRZDhdZQ2HuMNFQkzoPmANb6to3UFJ3vVt8cTqThu
fUSjCtrFmD1QlPgfYPtHDRDI1T50faY/lYb/vSBcNrsSoUiWJrNp9/eJL2MHMyrQdbz+O8nxUBJb
Ih1olGKNdom27gsn8ibuqbHpi0LBCVGDJAF0JvxqiwQBkqws/btOUS66A0HlOTVkt88ZV/yzO6sy
H/dzY+6exeKmdXTj9w7ESjt/FbxeHFwHQ0E86LLnJWDgYDuTiibWf1LCBoaaTh4VS1FGEwnntgKY
v2UVmWpcToFu5tFUuDpqonlqKGCbjhMT206K7XBwFhVVs43o8tPuRzZxeUnjQpYKLP+ig4LpW9GA
BhOgv6NXRx/g2XE5IYVXZkAxLKF7NFnFnuh5gRq9QYEkt/PFYunIm4TPGXsIvReQmVdh8oY9EF0z
lQH4/ya0ECKHHJYeRFoy2dQrVKC7BPkonhskYxzN4tzYPrX6sMRICSs2bDSqSpXQofQON7MmE2ed
V/TbI1W91QfIyXoJk3fSM7ylO2KUyU1QrjbPtzLAMuRGgiiwa8Bb7U1gpz6pNO3eFh1U69vSpjSk
9yG9iPg6XOmc84Z7UwYCRhc4iMxEnqM1rwuLet0cY23U/80LsR5tncRZNnsrupG35cajDQryJtvg
PbAymdcfUx9GQ63nqpLhmWs6W78XRd9euVnELsWtluYqff+QoT7lRvDfZS/1WZx9U9xzUJczvlNH
k+zZExo1CfKd79354d66pxrayHTMJUdBA3KB83XwLhUUnE71LKJPPPtfq2qBSrBNQ8odUvkt3c9J
XNG2Ks4WslzxBUKAmpUR75carNwR/wYq60fxeh9yPsKoOWu/Hup3mvQDo4r4yT5HkISqeerVYu0e
62pDz62WGqijaLp1twmCbE3uSLksc8vVj7jJAyxXqUIZmbzIklfjjAwpeEwkIV4UJm2JVGfilJRj
7y7t60UP5DBk16XXbUNv1ehvjlhll7LK1xH3FIeeEBrZ937eoh010tn/S2i5w0SwFD7BRuamquoZ
2UwrV/ufZ7Vl6OTGj8JBy1YmIxf1XdibennnimqVfqD+U3O+JlXBeeJzw+HQsr7xBoDkVIhOXe5k
wrBWlgLf2Aa9s4Tj6IKeG4Fb2Ee9p13Wb26m+wxGRHBrdVoL66COm2ULaWVzDM9kO6ArAJH1B5Aq
wrFdQGShTzbjaG9FQmnynsG10XLS4q5ojHSmqjwOkGJUVo8QfbIfASjZl8F2v9CDWn8bY178oJ2y
8rYL32NpcgVRNgE6bpjDtUgo8BUxhTHiiaZ3ttQPRk/BzM4VgyPeMb1Hne70Whg2go14q64juKQs
9FbPbhxEi233slZLT7e2tTXyKLr1jIF94+bW6BsKSfZGmS97p0K6lhTvwQgA9Z32LTgsIQdoUmAS
d4KDKgBbBr7+98gu2Q5sslaHOVBnrwvoy/S+d/psaE0bbb5fy1CqRGlfidThoZ83mA4n1wbOkbLO
aPfPmg+KTPHjEWhBDidJTFaS9YA2ASGX4cpGwP/FdIPB2/P3ie+lgtcu0E+mSPPStLu+TZfDfvAk
4DaTEpm6LUZXTlWH8kjvErNuk9pCt7+Ld2/p5FCmpA1EfuQ8G4ZoTrBcMeW7Bgj4UbTCO2ozB9Ag
nbCeOz0QPIPSNaQPrDCHrSgy7eBlNvInfjlldcv3vsg6Nh5XWDolauzo3GXEYVxAuGYI3HbjhhtI
HFY+GVN79VGhUkl27aeQGsQTJwhpdXulTvEfAAFpYSWM66S+3D+disOQa1choSj8iXAvJwfBWNF6
eO2ysDTgJwE9ohn55/sC7r6j/bQMYcfYagjvQsfsgpiMwW92KjVgHB2S4ojMY+jL/H7sIqSIss7o
d57sfpM8+jGhBOkOFdh6jFkC4l+/9cNJyxgLE+QzVxzQLcF5C4xStNWThUrX7aX1MNCf2we2kfjC
9ADXmj3UTJjhPZkhYV0Iq/N6O577KdNkDzAh1+6BShWJyhQ0cSfhIn1gt+gW/R0I+m8S+5P+uuuO
SElIlO2qcLGi2j+PwbO+NFUbzwF7ma6V+SYbm40aNH7eVZIP2bIW4J0UT8IVE+9fn7jc+1CcCHih
jtYPGMzZJmya5Kt4HSHPuqNbEJHIWESVIVQmQKYQje3SAxJkI8wlZJ6sxW02QWMs5TnB2OVv8e/s
6giZJFMHdw8qWBUpXXj45jmcs+u/sZVGJyU6Qi4YOXm5U2Z51ZijenFOxcowUCxkusBKdc2IpJq4
Jhtl1d5GapnFISR2D2qOAfhboXjrKLuxm7ZUUw/I5KoZnM5XSQEHEhQaavrr4dfGDtgmNXoWLPFj
3msBB0UhooCkmXaqlSEs1B0+E1l3ntSCuP70MaFV+5FoG105A+TmzqsGkv/dmWnCVInwlb5GZSqx
RGhzYt6T918lJ3rMPQp/aueg3aaY+jE3vCZk6622eoYp75s74LHb23BqeYT2lJ80BeNjg3O7wZxB
ReAo0Ma00RnUP+QlDUVKIx4Ac+0EZZkW/YpUFiHlumhi28wJFfnuXwPqTAKoK6VFsR0aExGxat39
oBDRKNcErLcIpvWj+wcRNrVmr4OBwL4w35DrHedmr1NieH39TNTRacWAYVf8l81b23gLpN5fO+yc
4n4PHgBnhNiFFKijNLDhfpulkcp4GWvjmJGAs9PGvOwh8KGqfM5V8IxRqnMmV6kaXJgpmrd549zy
Oh6Px3IujGLwSsE1e+vWmlcOF6vnLtU1lddZfMzm6GvxZYJ/ol6XS/wMm2b215n+q0vizYfF0O/P
/ztxaY7W90dz4yu+kvqD5vT385IQfl3DgvylvCok7gUePrjmEWIDjwj42xwZdpfSRpMRMqGtlVeB
r9sVtMjwg7YYNvofzvHeIcUU4hi4bdrBWFqiV2WGVxgDVONKoMYJlEWfGPll3v3N4NqF1Cw+IxUN
4Of7NBovwt7uB89WeD7FId+9X37J6F10Us2wdk36J/5S8GHPuCIbL1y6xLEUUV00BGDBuWvSB0wE
iv47fHs/HNigA1q9ZvzAn9nOiA5cfzcvnNPRP+zWfTj1Kbh49q65qBmfvww5PiVK6EYVQJVNk5lr
v1YobjaqOlBw2RDGH8K/dFvTLQnGvSotvfNlDCsl7Ddj1+XBA7jQSHHb+p27utPJwng1xbxIM9GD
C9vork8Z7GgRngfXAGXGWaEHfdISeZ0SpiLiIixdIxtUmiYiXepvL5mzlcl9QfGTMgb01nDuZ46i
GOu64cWlzkPlfUMIU6Era7Jp7Oi+5ClEUS1cs3FZ2cdM83/JW2A9xWCMYn0ipNNueeWgRrFqD7Pc
7Ad9S6k433kalQKw/nC56UtUgVx4AmkJQFNOfJzG9pXebwY6UhYBKagGTIxUomTFg9KOPL8CymfN
uSiBVaahn0ceJ3cFIYEUdvCf7sHzggtuDa4iPgkRB5mVrbyQgI0UvwVTPC0tpAqo0XNIMOCNd9G8
G2/eYht8XwvCZyXeOYj/RfJVMmt2enQTZiFONqBXrbnI7gGSjUveePWyy+S7a4XLMeDrp2IFmgde
wNvnlfW45MwW3ktRkpCcht96Tm25RI08zV3yD315eJcnYfjVneBYYiajDnjTZxxA2TcMrjJ1avLv
Tswd5tJLobbdX/HB2UT05YLiIzcgS1dnZW03SrchQjxNWdJ0x14W7+pHSO2uri0V6AOAOeK/KYpY
VKFXWJdLs3kUENkiBnb8E6Eu+REwbl8RB/AteGeGlh5/4KMmV24C9oI+uf3c9kp3I/3ZGbZ/yW82
9Sb39yrIUHaru1EhPStnQzNdqAf+6mnpB6w0ESmhbI4l9BvSdflzoBZ5EdCSPOWzptXdx7yENwCN
SOkYLjltMqrKxar7rnJWHQLZMScKYWO1NX20Svw8TglcKIeKw/BOVfGogfjG6AsZ+erJ/bqf+uHo
Khx9SrDsC7pkdy2onKl1Q9SgMUg+BtGESmUUxVXPHkCeBC0xjL2XMz4O2pn7H5dlLT/oaKgB1zC1
G8PLVbtCNtpZ7vdsKXkwf+ldKWbgq2MTrFcSR3bWknbONtv+2RYzqfNoBpxDIYdQykeBu54aRBuR
L95HP8AqZHfOqwmSd3ClRj+2hlVhCZYavpmIv78dy7AVimYo1P+ZCujbYJ9bCuoS95uLwwvV6C4e
aKnFTbPlkUIw57cMiqlxee/SsEN/f3BZdkzg1FzWPlBYSdkuz3y5xwaZwVUuM6Rxw3/zjRTpXS25
UgcZypve9YOaNmeEwQ9Qvq1ZOAI2ZACrIWjQ86zmKIqDCWmBvT/L/TQ5uHbYZyZohD68Vppdfkfv
YeRrCxqy7O7VFNPIBau8q1gnOmbdYWonO4Ts1YLBorLKlR7xNRq5fdJe610mfOewTPhINcUapX6j
eIaYVIOMQ0WfAzTgizG2ONPK75CgaBs6tmTefjZPdsEwxK7DzhQgN5u9O61JwIXcVUBOpn7SzgnS
OBmEW2/cUPCzDg5Wg0O8LEYMjfOQM6E1gWsn3n0CNhvjQhJyRpVaAMwWNjLlfEdVgx2JrIVRh5Fm
YO/wGjpftIb5197tNbMUkc3hZlM+o37QZ0BTIahouHBgRfXyif0b/DpKdBM9lDvP0r5iRxoiKKTo
wJBPUM/oHFjpTKDXU4FpJk9jurmMeNkGXqKmHCuGcnLXt03AL3tAv0BzFQiobd8SWfVZTNL9N64G
tqK4I6tj2L6yHmAynAWE/ZDADpSo6YFVH4sca97k49ZQJz52o0JrsI0jP4HpFwciv1mwUfh6iiAq
zI29j9nf84cde8N6KnsKzDi3DhNUnjSQd95nlEMU/ISWiQkpKOSYaRATU411VNFTDGaW0vILpBek
bT9glACU4Qb+zxClOmNTittEqmoZTUbi3wF9NxEIMPfiydzyJKrmSrFjY9DAxksesB0E1L7uAzT9
ZIM70XtNSGNWO0qn6k1Jzqo1mVbjSuCeXuyJ/iy83g4iU3at4nYBg+s80YOzhAqSY4Whc2eBvxbs
6Be1z2MfW14Vu6Zd33AVOhBIEHJa+q/DMfzhj9toixoMKeODQvmXJK3Csy8QnCMNLkJKB+h41pkb
biOPqY0i56Q4gumKv91vaqu6xsr5B0G2jcwwsSR2THPAewWckSK1Jafhm0+wmc9cKLmwtXNvFeJe
qg2bbZLMj3Z8HKhQqbXD+u450LWcR9aNePVs+/leaL8vHyTOaFGl2HgNXnxjy0mylcpFll7AeWG3
dRm3ENdmXIKUZ40QjvymxyP5oYfA+gA7Ox8hg7knEQiDOZVfHL0krHcF8fOeVY0uTsHjYiM8DzgR
g6kS9csiHdAFJ9tUIRaBVsoKA06zf/IK5TGvjOOjkAKLujo/AZ9sVMmfjyVth0rtEo1zVDrhLq+5
1YJkXj618mYFxGSc232erL9ytZKDWVIY0AYkwAULkKgQEg3HAj+PF5Us+gzlwx1FnEweSEGziFwX
4yl1KCwLBswSLUQDwKYEQBbooAU5Aksy0MxlyBgQRFhA46Dwpk0+PXibsWIlmhDr8plNTnjzP2V2
zNVYuIS0PXXygiXRjwxgO96zB1pT514qh28TUUIDqcaQc9KTNavJMML16UyB29+60IMd3KcGoNoE
JobE4NusT/RFJ45S5he/LiROGc3clY27xKsbNRsHpWEqNgRgCQnI0VgnOm+F534YiBESiDCRj4DY
jokFGittEPs6rGbktr8QTX5AHhyk+ICMrk+5meNI8T3FZqYn381kOrRjXQd6OHY1tI1COaT8HDMi
AtWtpK9ouOxWYB6bZPP1ZVfPVo5pIv1XV6vjzyTLdVSBtxOxJKnLO0kRWAeGel8j0OwXAf2NdSv5
mXtoWR6DDEW0O+3XftnFUsbaFJQqmRBYolZkwBRWz9dBtj2lHSXlZIctJwKguEtL3XoePJ3o6dxw
ecNaUYxQL5VymQ+YQFqeG2h+zTaN+Qd/v59zGG8uSDo3/1cgjvaC+LSFziGbj+svhMOkAXpJD7Vj
5qZVDT7ccoHJoAb9siJXwtilq5q8j1sNGw/SYAYIwv9e7255cWqAx/6BFCkGKTSl2E4fHPJ8UvGZ
4FW5w6NSvhNsIoUgqbxeskPmEErInnwq2wKJU6ml6gWHjbYzr4VEdgLxMl+PTtu3WoiRx/vahKS7
yqQViqOfH6EOSZraH+JYUspZT83HQDQURJMuFj97lEvHfeYGjee9VVao+6Dwmo0wQ1TIPxQIhI7a
JRoTc/SfqCkYWcCzDHacUJAALkVpAOnlMIVaYMJZ7ty8rKBQkQ8/y1HM59h3T917eAbm/H0H8ctn
Zar4f6d+NJzon8KOjttGn6gEqIAfsu0TNcQxL4or9sY0UqdXYrEJJtNd0TbIBjhQ/qmKG2xYZGUz
5gmt93LCPQ1VfviHF09QLC8zuqBiMHEtNwHqPjajtQfjdKJgKUOr5zg3kzwH1STd2vVvG6fp2kNK
6iMr/KFkr29pYiZNIZhNSJK7r+FL/uCFUmV52kaULxyjxSNm2tvcBUK/e7DftXgxVuj4cT+HRV34
EGDhqDjHu3t7EtMsYj2zvMt0F+ftXl8tkGKXWEJ7etS3GziTBhrrvHHWimpKQ0KdFCRJR6xirD6f
oUCPC9Sj3Nro3O6sli+PD9ia3iUjIqVJUUOjDlszUkyRtFZTfUTy7rwoViNLn6ZxgkVE2t0u/H6O
3DW2G1Nm4dqU9U9WCfRzUjFMeQ8YLbusYlz2TfKLhmbop4dRnVgvWpaRRKzt1U5Hrw3xsXKsFmSl
j6n2UR6HY7ILvWCFrUAL5acsDHYWCzLYRM/AvDiif39XBkI6HWH/i2TfgvpQVM0/FDt4XqlwuZrO
CWf3lS3zpTCX/lmm9iUG9BsfImbjPU7f3RI85iWHeF7pG48I5dATY9EDJGquOGlasJKDQPR2ucYi
mIRPcsVNRKIGyDv6RpeBSPQzlkWDMGVO108qcOlHFegCDQODRraY0m6dnqoRHyO8QUuPH//ncUeo
iqNgJuRBEkxWmR6renO8SLPjhNzk/LmQ/faDK1rzMbrs/pyHdcn5vdx5ukkJN/DDMd2cRNSCdF7v
LKxQCWrNMWAbrEi81USwMCjx9VgSqevDZyO9XZ9g8iEdhYjVIbwaJtDu56gCS2blySJ0fFn0PJJH
bm2d3b1Mel4okvSdAlLl03I7+2Oujt3/6j04mL8gysG311TKf+5jmNAFWoABmk4rTy6NXrbMqjr6
TB7qLtBMdB/g5i1SM119glRoywaAnQv1wIzK1Y8MdvB8ejbGTFUZwWepHB7K1seEWrbMcvNRHFSH
5nU4jAltZ03R5KDpr7gm+Ob7zcvGQBG1pe2HFH+oQFlfR0xFrg5VzUxrxs9xq+k/3q2+2D+4pw2/
wIkdEJxsd1045y1EH6Xq18aORImkm25mN+YxfMo7h/gedtByJoFqcgz/5Oc0pIyoMF3eKwakER8O
S5zUWUnnjwj9C3cQ+7pJqe5L3gm8bdgwv2eKQ1KvcMSD/u72py9sZrzsc0o8XkpimobyzKQbXtOW
/Oi12XVfp6CAg+afxZJERu5RofPYPTTP61hIBI/33H675U7STeO14gtAiycvMg2bIrSzszLANPjz
E94Fab8TA/h7Mau/BkmVRRxZk2Afdaougq67YjgSsugtKJxLH3AOBnsVnQsSdun96/zfTLexRTbz
twm5KLhZymvCFz+AC+EYTHID6QV+qNj3IMu6GhY38fh0Zjwtee9uBKMG8vcu+FU0jlAHGN2IFz7x
/1LXiXCStXSfepdF89UcV1lgMaS56G+3OM3qH5UhntO91BnQOeb7kzCpnSSYZ7nIKQxgKr2zmjBS
ysLqyOKJk9gKPSbOm87P7PRQgG/Mg6bg0P8fcjP3jtBmPR3lQJ14cVBK/wBvfuSVCbaDMnss6cKJ
cive27L9dUnxcls2ep7k7MEp6hWuuwZ6lT4EHZHHO9jllVcjRTDzuhymC+eIcJl9s10gLWcc+B9V
Op5dTbMX0aXjhK62q21GC5EEvqVperqNJF/DiUQHrQoQki4W89+GZNomzl/yCbnt3LmGKhepBqr3
A1S8TY2gDjr90cR8X0230F7DUk0/h7fP5gXyTOH6BHmS+LPFnNw6kyFkGjsfo0rXPgOnrbSI/vJo
G7a21OgtTXXh1qHlq/3fvATWPpfRRy8RpV3rINADAc7ymLLCt/MMG2cw7MHxLwxNiXV6R6PAyWsU
kbLlXoKBZbmoGHiuRZKvNv54mjNFGgoTWXt3sc/HthW27M6+W89X6kYzmGuilbcDckcGrybFRzP7
oDE7qN3z4EQpNmkbalddygjaajmQi2lkuBUfgNZKMy3/S53IW2Up7QrndMewvR6Eq/iLF/LJUVfw
l0RTaLCK7AoC1iZheCpftUNfJB07dWxeL6fQDl4TucYcxMuXWmlf8LDyNLqKc47l28j2qSlHFGbq
B5Z0M1zgH66eQplzIlHi6eFEMjk1FUFSW4CPwUSc8wPI+RRtGM/kUhybOd3l+DrW4RqFah7zrn3e
8OODfR8YyfqsjczlFweX5U8eyYlKiKvuE/qdGgmXuqTRG1ovF2fPnwyrzPb8TkfPcNdFNCBKB7aT
hwzGX8PjAtf47r4Ln2kfTwzfrElqeJNk3NHOEpfzfcIXXWTQEMqpI6aGvS7YjbKnZEVrfyJT2KWq
OE9pE+KVpV6ZvnNrn/nPzbVulqZaniabjGD4pumuFqnFwP8e3B1bPpsdhe40K7pC9gxEDvNxF4AC
BFalc4RisTwQ6Qar9hjBcdTd9jKTU5SET/n6KEQp96omhuJn7KkprT+G9aabYV4ha5Yr7xRGa70g
ne3TxNeduas+cX0O+aT/zQOKjnCpMi5O97al7ne4JBu9RMmu+tfGQHKHsyPI/p+bsWFQtRCwNNzk
z2aj5fgaaHya1s72/HUuNfNkTrSirP8vMA/QWoF6YJ8FAOWVpTL1fXONwb9G9veuISUTDZsL6gIM
a6/wPT7iqgbslBiLs/gDnnEjyx6b1aX53jw6whAnzivIUL9Wj25rJd6gqCLUsoBnUl8fDMeNZ5Pg
/ccgiMOeQq8sEUZWXV+47Ow4k3CmN2K7TX1Mo5U5PeQnZZa21+31vm0Mgboccq0SqbH6hW11xb34
kgrZ1l6g361g7EvJle3Y/ka2BWIsF2Dd1sicfJBRnO04Ec5Bk0GGE++0w96VJLSY+TFoRF3XMPCK
M1jC5Y2gGHAT/OuYpMNmsxPwD6k+no7homcxDzG0SJbhj99mGoM8K0+TXG0AKhFHUrpX6lRIxE60
2IeDV2a3XzbrH9jm+RWAs8tgbL0yLgSVIGMm3n4m+ATWL/Qs0ez2RWpoew0RyVCIociG2UpkudoM
r5+9RGtd8vM8OQ/TMhPMqQ2FuF2hgxtMDRmUAgbnfMkEIUVPNXCW3ILOKhBxUkkhZogdtsBkJ7An
CoCcWGUYFOtV+xdq0nObD0iiOgLZZUPVUEfepzyhwWSTDjvJp2YXSzOkI9wdSwjHlZq6j/GXvOZ3
zJ012A2/FEKN5fqMGmTJqhpI/XcUqW+jzJO7HDkrsTKf4QdiJqilzZ3v42Mjefyw3yXnBvX7cyIZ
EB79Oq5HXQRDwKFmOP0fOvJNqHalFKJZTLHMYfcUDfwEcug8W6YK6H6VB/HigigVruCH+tPeKCH2
M0kI/HsBhcfNtmnsUOgruCARI+2PkRS83TzrtETg8ZUi85QxKntq96Ni0CEVWvo56Vn5aEDPa12H
n5VRMygNYzxj+Qr0tcwtsSe6h7KTdJcc9uahHQ0DcjUQGZsNqk/lMWJvRLYMq9o8q8MuZxYY1sdp
1Ytu74vuvwnHkX+KTqFV7X+ryxeXoiBL3hadEZL09nNglyEgREnBourMprsMKM50L+24JEDln3Uc
vWWP3wpOtne+Ol1o6/CA6HtHCxGgoH5TEIaPwqetqverIGOLs9n70Agk8PUB3LvfAEN/lMnbzgu3
w4x0szfd4fRA5Wf8Q8d9QZuFubTVvQ79INNHDXJCg+3S+PXUOT2CEn7bVQn3NmSGWVF2ItSQjtRy
O2n+Oo7JcqfweX8REmdVC8CUDIZDgfAapYglOWNrt439fLcIsBMAytwtynOJ94rT3eySj+TR+dPd
vazasSmtOemto7k/RnEFCm4EOYQw+8bdm1AExTX3BvPbcF3M0dvko+oyLgTlPty+F8ChvrXo07PE
bgAGVgTAzHCVFotRX+hbm2NVqbxMMpffNxw5r6DymXrCYFMEEVY8jkgkRX493yBA8NwaWApwMr+n
2EB7VajW34tjAnL8hUpfqqCtk8ejhkerso00vABbWl8nIbfGlLsUd644ufoYWbOJH4THpBstvxvc
yQcEXpzhY89fSUjA2BoX572rvQoiqNhVQ564UgOMtEKidxChAWtO8/xVhYmdO2tONCNejj529Xpj
afmS1ffvSywQTozgOrFRdYSTgBu1IhdPpHu+uGx8lCzUpoK9XugnDJILzpmAbS5OiraGpuvMRKoT
pIaMysX0RAILOX2aWJ53YY46GIzma6Xn2tP+fgWAUbuRyoHvUshm+zDJsEkrUhRPM6qJBzXLZJvy
WEuKGs2KHk2I5FPgKRlgQGiQiTsVXQ7k9amO05WQA/nO+khh32i1/qKhZ/Aw+Xvy6XpxWx7rJB8u
OP8/aR3wxdZ7QkVFcZy2dvSeKP3pfVqSVgBfU9bz5+STDGF4FOWsM7PDWldZ8oHByXZzwMn7CbB0
hGkC5VG9yUZ2l6ioXovYWcEWXi8hw5XriIpVkZ3SiVZAi8lk15bHgmzKeyKrIGUYES1xXBgBDprK
EX9b7Jj9Hv0VcG1BI0IsqKpJuJDdJ4dGiUAKqcCfzj+au0d33MeX1DkTmTIEwY2s0MrgvK1eQwge
+bwqvwQ6xV6okxxRCglW0rmS4ftN8Srx0mV/efnBM39OQwa7i1ILgZevCpIzf95bvc0lAFLOW0yB
V6y0lNIv39HdczAEi/bapIzcq/FOozE+B/I5jVlnS6ukiSKRVK+XU/6aivqkkNp91nvk5LFXDQly
kLN/7Zb2UV8ZDdUTg4sZbSRjxLegIrDTacWJ9vCbc3JWrSiYdKIC2d7deNVc7K7qI8FliegKH9qH
ccSCQGWQSeh+nJY/JgZk+OVk0rr6jiTSPD0pB+fSJPoJW9OaNVVFPmL/6kXNPOkLaW0fle1/kFxL
VTlShOqrCV65V3JeHxPwQ5F2VGd02aYE9eY6TZ5psV66/gZ0Gnes8p5RlN0Qg8Z6MaOhhIYnJ/fT
JcI4CD0v8mOseBWp4UlHsS95xPlbJBUlQ2L8+3S+EizS8A82ZJrxk6UYZtzCN69U2PXBtGYQt/RC
WN5IMLG1zT5vLTP5EC+HZmzP30dtejOL4I+ERiknhq9+whNZZnnb/9zHwo9s7MENrZCKy226908N
THL6NaefKaIgrRVhvkNgmi/CRn0g5Ina4UAFtdNmtqhZQaX0LsAdvLZ2n7Usc+jTkX0cSkfdEMa6
7Y3GYHsGD+BBZUN4frQHY6EA9guSpE35laI1k7C8Nc5cV8/fhLGH9B9i2BDPh7KIGeKVtiMMD5YU
uv5/0LNCCfwmlR8z+smaepcYCtzjCXKxLtvD9/T61gvYYxRnLKfI3VpnnTcXK/863IlkoD2nqMsh
YR/R9dVHg8Otyf1l2jRBjz0dnz0dWbRd11FGulEtUNoWMVGUPGG3ScOBr5NyJaZoyyJCQF3bM3Ti
9R9yNFxDCa1/qaR8LQRkCqlzQNE/63w4bw6H+2P6h0kZCj6RPPftomTzpRo6rEALBgiKEmyM5FeC
yxQ9ihrdxOF4o9mZofrQMmQtvsxthhcXooW5w4RpZgMoYtjm9xcScOqCXJ0tH+5g7J+5k9toBLCA
y9g4wr23P+uSrVdk2PYR8h/T1NzAKYFss/4rk14mOp2ZCmUgZ9Yppjm7LcaaRRST7GYfAP8IdJwZ
UIxdi4KRFVu7Q5SY8XEWepWZSdJKusEP8hfrbzbQhaJGUI+Swf4MThVlARAs2/Y1ZuF6FYXAEBw1
8NF3V0xrKqCoywisCDeako0vnKpoU4UmJA1UQc5CSgRwqYDUBSjaDDQq5tTbnejyASTGkyVAlnMC
Pk6k/v1W5I1ogvonqTKkbkWi6iQS4qBHygig/s/N7SceGzqJbXgUmyTZsmu8z59YtXga+pzkRXs0
T/7nIjeflCKrawq4xBJRPd1MvthhksNW4z1XIUdyX5C0/jq1ymXKb0h1CkpxyWvHM3hn/ajQnCTT
EyXbEpEjwC7GSeS2sczRxDyQ+VR93l8VA9mwod3vo0qMVpxgESyL/9Zeb5hdO0Oi8iCxvYcaRBjC
6iPtEj2jHPfvrWp+9Vl2Nz57jWoNEOnCK5l/oBJFpPG7uN+mS5PkY9JwMM//VHt0TnAN8KIXx/Kp
bEUWbwegKR5Uj5ufghBkiGm72rC6s0rz9ctEdOtIyaL8CsGXGwHvyNFV5KiGx21tmKqH8YHRe9k4
qtYJ1Ht0nWp1Pq+HfiCtSVSHw59uPOxKLYwnbcyHsYQ0x/Vkvxyiwai89g2bp2HI+ztrd7zjgvoB
t3NY3Y1I87Rz6ODx3PJsmuMo1fks8uDmfR8/JeSxFcrRBMS1v6HQY4V9F+zrLHxXWI0g7+LN0nvH
RLu++MrZmm+8tJOrzMUnFfHgcyiVJQI2YwAGDTIT60dIWGLMKE16YSl3jXdki+wdbOMdkry6GCQ2
DasPI6ksGS3DY/qmIPxzvg2eTFeTMdfr9C8Vv5K3eudibFEdg/95G7pOezQkjslp17+qRcjrwjBI
FweFSEJDrN10H5tAvlLSgebIHbwMrhxQl3bFInDOxm34eilJeZaWHl5cxcq92nyvqz/5k/tsmLjF
HebXW1r4eyp2wtuI0uhaR67ZNJKQT98/IiD3JPTm0LZQXb1xTk1Ku1ObF3Fhbhc+vg+p9WMrLc8Z
BBDeXBOeC6EPaDZyf719LRwVE2IZOaMAbDxW9k/lnPovWvynpAeW5Fh7/bsi5tilaNBbvIO6c79+
AGU/1y9galdegao0Znx1Gx0Bl5EQX+Hgqv+Y9VcO4SWBxT7vsHjv0Ldig56ES4MfU1eipCfoyuFj
1jDm1S+g85t/vF2IcrGjUwtbg7nmZgfk6RY6nXh0VfiTlidDf8OJ+awJDp9HCAT+X9x5Sslu1h9n
+YO144wzjFQi4kjUMELU3lk00U1rANfDv/4PuLJhUGkUFpWP5WoP+U44bS88NrV12T3Fyi6Nw1FG
3xrHpm3QB2RMe5yOd06r3YWbuNg1RIziV/LZwlMZ2poLZMpQlTEXX2HPNlXJm02n1yaoHMKgpyy9
FYD8K7jlS33M77BmqYlj+hqszOTNWwQVRJp9H7n6Z52hLS1mv4hTXsDDf2agOf/gw0OkF8CLI9sC
yMxz+Ph7cGkuFq78yoiZI/q/JsF8Pm5tRfeDvRwcinfhgTQtFWdra1BX0+OYm+8/R5CPhuRdy0/Y
DJE74s6VFBSylIkTvYnMwxXG9qMAr/k3mv25P2KKwXkmY2pGoOkpxcR6QouJKbAzuoFwi/CcoPYB
RCp0ZaPzISOcyj6OPBxJBhdXbIhe8ipb2PedkhCooQxjj58S4mpUMyITyqd598BjJ4NpK4sixzuO
DghwhUSRHAANNnEqkEJxtseQHNQ70E8pnKJC0Cy1zfFK6hBOR1TjM2mM+cE2RocxxwEXhGtFnsMZ
NGiUdmgSukW3TfDEe2KM4A3gqKvVQmDuL/gQ9rMwdZ/zhOZZW/rmR8sJipcOVmXF6bUNwC6SVINn
Hz7Xd77N+6VcwiMGccv7VYTTpXpnivTAmdXoEes6e0aFQbQlHy3MJdRY1arCZiehOMrkZO/kUoiy
0rW6lngqsb/PyDuFi7yDXhQH+AXlq/KBSSbHLNlAiRvSBpPdXI8IEblK60bogYkOH4ehqWfRj8tm
2rhn5iA4w8TYFNuzpYSrcZzcCBfgfedUaZ06N34iSO18oDsjDcZlaXqGFCsWeZkOTUC1cZ1jdrZX
amG7WnMrpdVRQol1YZnR9aQcUYONey2HnVtWYiJtXV3hfQlkvu0PUkOmW2CPi5eir5DiFDgQWql9
5OCSdkKYkra2g8aUbMEl9t+gx3vzY6KRbrO1cAnNNrmKclMMCE6kggXiHLKxo/KyZltcKdLyiMnF
RbYl8W2Z+NggODYgo9fLLKc3uNYR/F1JNbda2oRiHc9s/4f1T0KJS7SvzBD96mC/szeZoCwq3pNu
+lxDTDJHQ5JqXNj+5/I5y5Cl+Cs9QIX3B18K8NP95JaD2El9IF8UiRnJjucwxQuZ3DDPJyF7togo
t9rBKkWQfXj7B1oA9OEGaDtaHR/fwWJL0AC6h3eoc6Oe0//KKqEqmbt1fCmsa7Og+uSRgHlgxPIQ
1FnpbvFmrhHV6xnugQ4Dkzz7wJAXEWQKjzoLm+oD5AJ5rymNDUVq9ueMac0UKjgzF+KLkWapU8Dt
W/mAbwRXdq6rhelUq7ltfcNd7QHBRG6YzO6M8P5a1rxnw9jkFiNOzsKMYauVRoFw7BlVO/DR/lwD
SqYCM+AgSAqFUTh1LeSMy2jQgE9XGE3QVHRFJxu1TOUvZxaryaMxcMnjv3B69Fzj1d2jB/09yYbx
VTy51BLSkmEJ23STSoQhdKFnv5tWo37had42Gs4jLcOVb6XGowhPnW6ykKEO0X2kiwGprkkzu1Vb
jvFxqpD2emLOvwcFU+0RKwMXi8jH4plehVBJ8eSiiElypWAW6W7S/TrCIUQRKLAgs77EImPy+am+
CSCJsyoSmXzAWbCcd5gDhdpP2CgwCeQHUOkc7kqNFBgLSVIe4SbuGkdIapP8bTd3dhwKIjf8OK/b
W/SYDJN+vXrJdYs2tZJ8dhsMrvFlXdJxl8MU7P6qU/sZdVzyL3vIUhKYxM1WMyERuyOfj2HsERGQ
WERWs0kzAuhtxNu1V/HRBWudRkgVGMRWEzJXXrnrXpPg6iTAMYCwU3giWJb/CTCB94Zs7cYtlJpb
BXXVIsaT0JZnWJHJRWffGAz6QdqnuVe8+EkeFmC1pmWtk++/60R/NTGL02eXwevp9qCJpCWqSVgG
SFKbnnmPwsYexj8gGdAvLVkwp7xC3PVUmVidMK0poPBX72DCXKVVnbm2aCQR6rKGKGrBtJLWuxP0
uV/F7hhHrUCuUQtQ7U8ZY+7OnwDryIlhDxdQ+0a3Z4JGa3zMgUT7YbbHnOATJrNPtN616K5dCvbf
t+xLbKULtXO+1vryMpMW2/lMa+/8VHwckxqgkEzhJ/Bb9uTBewtWc6nJydtoUGM5W4HamqqAxEj4
VxLQs5hD0m0xRwqGqnIHtTbx8YdBhO/SnTYg3oGrRCwIirEGhRbA/FERbYdk+gnp13bIAt/yRd/L
aJLYiGXQJaqmNEk4m0kwOZK0YgIydk4zK1eqnlM58695bgjn1OcdYpJzG0SZ+djgG30PrAIinB1M
JqZJuPoRT5lWdLONGSz+BYX6jnCQrkyL8Wn6eplWyQHGBcubfh2KyNZPlfhMOxFk1DVZR//YU+1C
jXDDHb1A5yIH4J5vcN6eDvl8jkNXkGGHU+q/UNv/n7PvINupIlNVz6/zopAmGtG9HIxgz1pqGQfh
B/DVi7WDci3WkpKVJ5RovGtN/QimHp128CGzbQgS95rboEkFTCVzB2kuYl7tuc+rl/yV1qEzIJni
+LGwhq2Em5ug0u6xyjBDL5jmQEcG/1zRObWd5s5gWaYJsnzgOZiaPUr/4Ug+Oi8aH1UHhOSSAz3S
xEjCjzMgneF5YcsQFfa76tQbOXzhbsv4d52/bxiMx7+UjaM1sTa59BnSo/Vut6cuXPSGJOGxTa10
OqcBKUN0yol/vFYYeD2Vff3y1Zg4ZdTLTvCY0ZxdTLmh99SeSP4trH4a0ZQtk63XNG9GyHyukT1q
2JN94nL+QrrgxZ+gY3LHyDzgoXe+6OTICrpS2ZBEF6C/t7Fh24+fd4CMBzkzsa+sZ/HO5f4UDEJp
5qNQ0pCd7bIyh5tz6N0LZpofatvnu0XpVioXRwCLHg7wV49LS1ukh7vgXVmNVN3ZCVJlcg/MU063
aXvUYjqBlkr/M91cCTAGWkTjyOO9dKsPyEHTnMHRO4u6Dw7CBwgyYUb9Nj9PywPC9eTqbk30U2xy
9MRdpByHzHw1a7CJn6ylOgwAD8kYKpq6Kj6aQnyJ0PwCop1k3ibDqnlmAm+dybUcPRxXH5ByOKpd
34O63vJO6Z9ZscQmgE8bIP7ch+77BDW+J4LVXRngFejFFPdcQBpijfPfv25uDwc48uFjOl4foQkG
UDM0zLWGsmq0q/H9fdn8228qc5K5WhQk5SbXZF3bBJQjeyf1x9bg5xqsBJom+aJOcBP47fMTB5+2
IDipAh0qs0RJGSNOot2KvCgmqzjLz8NQNL5YSJ7eDv/OuVGY/Wc9yIiAOkSS7syjPGPn0HLha7w/
gmUvkN9DOY7D9m6SEvAQY1/TJ6ZWS6Z1c7wR5KEX3zL33cd3RX4Ss8eqnPki02sxZryDLcGoan7P
HAvKsdOIZLZg+526L8sKy3LmZJQyLsHT29HWTFqFcrE00p81S/qAGF6QDuyFy5+U+as+R1k/napu
g1rnkZk9+b1iG7/8lJ8hF/SW/itWhOkX8R1M3lIumGgzH2Aw1e1wakfs9Fix+xBqFWMjNNUdFBdI
+nGWlsepZWijoBlpUbMuK2sKDc6L9VPsX6rcpi2eRWsFDa+8FQKHv8E+hC1+c0q0eEtTsajUV+s+
jzz/JDayNsiu35Qj9rz5cekAetbeD4hbjUs0qx2wYTTAOnqCDpaiqBnS3WPUhPjGuZn6pfkb+axk
z7NlWXa2oYujIddmRl70/0DHK3z4DE8oNA8adJ/h2O7jForEJkb0lPuIKoqRrlSIOrgw5WXim1+K
BQzA5EqTqjJtKcNFhCJz/qSNVyycMQWCEveK9oreLdeoixANtPxUA2BSyZuABc78nFDSK4T2d/zR
OdVayL+SGOm+LZLyN2n3XDwLtOlfOzjMBVgsNLD+XJrczIvbH6ec8fFtO+EHpJZLbkWhvPU+hWqi
m8JgYXY3urTnu1YtTEeBQqXrD0jxGj8dcoblq4VTNAqryrmm/uPaly8S87xNqfKKbBuFAD5RoL9u
T93OB3mEj/WlHdwQZ7XCsObQx/eqWRvoIsIge4SPk+GSHOwOMbBtiOvmxOwIJTTvsO4o4h4IF4e/
tCdHRXywyJCaQBT2Qj6Kv00/1mV4ECW7VQizZ9bxFSrZHknsisznytNgQqklshATREHJeZ+tk+zl
xl2Kvy9gcmsO44cTMDRWsV7rNdmYb5jtavm9go7IZoV560sxHgRhVGJc7qX/VOM4yuYVmE5W0Jtc
1WYrGb8SGy0LNkEtB7STaZ7QOo0dsA1vQ3dVSYt/77Onar/uBJv1B2EycbQGWBZDUWvpnVM+E7LC
5U0/r9TetFhzuinAoR2JDcLRYfGdtWNNjup5RGpQslWbW/QPBULIbhwyp5/gH2LphC5I4jzi267y
1m3N06p3Hv3yjODJhWnxgsO/xpFgAmgV4mqS/tNLqokh8izMS+wdkRkT01T1PjMS0kxXpl2H2+nz
RU+SZMMNud7Xp/CFGW4WsIWSJOlyobUG+RCxe0x1Ae2KMhl5Kjzz+euNg1u334PnPQMKMeTuwjeX
yXLU7UEb3My2JYpcurulSmPo73s5MY6wvuHbiDABSXuRLB3OM2thXq/t9dyOxp2NM/2I2foCTLdy
uKNDQF6lhdr+oVLdQat82j8WKexk1YxcLg6vjXvZ0zbV6DKfV4dOyCecKjtr69YVo9+0yaD8ml3n
XKwMu1Vp3hXEbaFtgUVlTnzcLKnsIWyIaWM8BcKKF9dau0/IEfkjP+Uo2Al+8X3Q70pQYsblsj4W
Tk/OyZlqUOvfkxrn7Lkn9XIEQmfsM7jLPZyBUKjkHptWJgqnYIk7hr4fdsmO9NU3ND8QoZ0dZ6yV
s7aXLmUHCk9R4FMbFnMIjSVStKU8SJ35TC1OotBv6NHhsTYoU1QlKAecDQ98/Kmj5A87rCsIfaqf
Rqhg0mnZf9PDvkCSLWs6ejZAEm912nNE4yMYJOHn2YEDtHA9fBaF1zrerWcO2iGJ7rAFXlwCgq62
MiQneZk9Y0r6UvSqY+RUmJ+oZbVkd6A4u61fFSUH+i+KGx0aqvbC6taMf+g0Q8QSEs10C1dDL/+2
fqmgi/iBNyuc1sFTR2nrdVuuzUV8xAAdsezMMW5LQdZgkmW/E/WI25SIqtcMSsMJK/uQutV7gyGx
AmRBni5j5yflQRZ9tCecpF0fPylmAkA/fv3iK8n3+BRB2ZyNuOLGYsikjiER5OhSSHlgQD3Y0uF3
SZjmrwoSEE7WrWc1F7yy4horBCVjGMKhRXuxycmVrCZz59PUonjVbc6HBDYqUgzNm15ve1+37Wxv
yA9yrM2MCLhq/SIT0Sdm3gzoXaZjoDip53JjqV8j6O3zSWoROobndsy4AXv1WWclqMQp7equVB44
HT7mma6v+FcOclOfmQrTuqti1fejpOwiwUSJnV9aGdgdUPSrH1fTgH6Be45joZDmqHKpBIqNqu8i
eLECZVNJsA6nPOBlX1vxPeJqSENqJs5iKSABPqQ147msq9prxKZ66ok5HMU7mpYBGV4Keb2K102r
wehu2hW/p307WVuCA9ytRvDojpax/PoWoJpRLbPJ9EkLO7c6cn0wTq7/36UHAQ6GymRIRYcsgDM7
2jqTiUiPmGT/6Mi0x3hykOKMo2soyGbYeJoKoo6t+4l4HD78pRIuIaa7h1r2Pvl8XNnrkdAmjQ0N
51z7YrK4o3R6jhCHbP6NTL0BgcbII7D0MdIho21lfGkMbX3K6k/2Abw70t+pZ1ZbhrmUQiQaEFuN
pSr//QabSfR4G74jdWTWZUR1EI91KJcaZornxrrN4LhZ+OhH+sH5wUiRP8AeqA420dygSNRVReZc
g8IyCHM4JSLhpyD/F7wyMjKPJyYroETMuT1IexAukFGiaWDXtrVgR2aS/0z2gCZsiERmkXRkgKuV
vvjUN1rugRlP/xmBJjlvt4LRHvB4DZwQOzr2UAuM7OXvoOCO/dyCUp+2bv875NGFufxxTuSdELiQ
QzY+/PDGPZ50wfxQ38wTRWnV1Z1fkBdwvHv+2y727PBhN0rb8RYpUOHT2cg97vSxTM+Hf1dyPQ41
ierzOK5Ax6HbWdPH30Y4+1D4h3Dq68bj5MP5E3Ucyp3tflAU6sW661lHDeuaJbxFaScJ5oXnGPTJ
/EftckrsZdhAfuFSamTycHReNbrCEVbWYoqE5eD1svBlydCDZInsohveFh4NYD7KFqnX7MLUfJ+r
BOGbWhowEXL0c7IaUh/9FwysVmTV/cuUHYkFE0RDFjAU2Vg4V+ynAPiJNLnWMCde+Pt6F4MUiVTL
XhIPmRj7UrUTuXyuIgBGtoLrQfSbgeWneBgLQgm9b9+ufpeKDsSObml5QVRGhOwyd+LLE+oB+Y00
NlLe0HCa1UJv4+5EdWVe+5a/HPYmSi8XD9mXTkJvJUVwAMgtODrwI2My7c3GDQPPYEuu2mZHEFWu
Yb/GZsnmnDFHMP5741cpFV02LOa8VKoWA25PTNIEN+lxFaChgg98gRG9M7X6wYSUpeDZbmjChpOF
W4k7F6b6eAos4NHr0dEuwYPDBO1tKVgk7vP4KmuL6oie8aHddN6W863D/ZnFuD18fFvc5Yr4Th/B
G3klQ418M0BurtsnPDqDhe3xAzxabcWj3ABCRKroRwPdAq2g+P1utmY9ou3uzHBaOzRGMnJ8HgL9
VO5nB5hRJCfa8dxHfaffbqOQwqDmsqdInbAz1+mkTdxcFiEsD6+/byIORnrCvBjCLKYEeNBIyYWA
dZvb9u2DR4TscPDGwAV1V+lupkfEoI+RfBmo55DYNmN1QMP/uw7EwlEPEX933H6frl2PcYldj4OE
wnZFgWiiBUZvwFawBvuYOKz/cHqu74Yw3PxZ+X4ZIDgw8hjA63jgEGnsqFQR7qTnKA2Hnh4mpRyb
kH+/Wlynr1i6UIk1H7tA5FNhRPz1LcDhw+B/ID/gy/Wd5fMF/O3F2b4sxMBfbTgtgPW0cJwIkzg0
+ltYuYYC3RfAbBGBW2YR5RRTc+kmVs60++zOqpB+9w4AaWVWMRtT23QTYxeVcgNCHuDtWtyVOWWh
X9vdofbymsn1/IVxXaWB9kiCJgGgn5HuLxbTqCm/tF/e3AVU4TGs0qWTWO1jg5RiXqHp3EtXnKMJ
UICfx9K5uUJkmwX6zbczujA7Mn1YIB0HB6DmurcTxP3g9z8cCErDVfOQwQG+Oj+6IAf//NALsM69
giIi4IfwZoFWs4t14n70IXu+DU5ds6p5dVJh9RvD7qvHCATCMY1+9TGfE4Fyp2bhYVG265MG59hM
2xJjZzujOmMvkSTSCIElV5KINOK+RJN7cVToAeB8x8nN1WFK0+xf3wLdmOwirxgSy2j+WwDz7Ihf
Nxocp+aedbEfpcGAGyrfncSuOL69gbphyLeU5vAGH0PM4yw+tsJIKWktEP3cXAKfQIykBioh7WpR
lZYzZeaEWWzej14r8FkZfSG2Z/UIXrN8cZHV7T7UcdyJiPv2ZIopm1SnAWYoRR5TDdTnTe6HCpWd
gATmaA7IbKIGEW++2PPSw4LBc+rP0xrIdsVykMSBoBhcHbKwmucU8Jxqzm6Hiw0G/HFs+gxxsLiM
MQdGH1j8E/BX5bztWARwoBp/Lb6Dc8W85Attc+48c25HDDnAvyLhgaCzYbhYrrhAkMl1bJ60gqRt
UXOU3zylX/Yju03D3Aztr8TRVrYJ8YMpY9a3kM6GPwgD6POCS29fZQcRNpTFDAq8UwqGekFj/rwR
RVcE8gBCNZPtzKyw6jR99HIljkX4taesAD1m4inxU344lk+QodSmUyXHYTFEd8mW2Eq2IhgsaAqE
+rYf6sQ/XsZtcAtUbvR/jhtT1AKsCafjmA5r5jepzYH0Ab/c6gJWAsPI88JwLz5VMSk+EiPqCJ6R
RVs/6u4RxlLDyQVQB2nfcQQ0rKPAMt0Pu+Zx1vY1ME/oIpQAoJZbze0ERDgR1avj+cvxgfCqmPLN
bKmmx+bqnGQiYph0oT8Ejgf0QQl2fp+6lTHrYPQpJnv1ywisLv2ANKgcyZHBTPLbkWv2//8qcvoS
tR1prwO5aONBYiyrJ908/xBbCHWz+0KGKFMRIrYtWN+vXi87C6V7IbUexKqvl6tCqyPQRcwze2zT
VmyRXjJ/OD4+T7EGj3jBrcCG46ZT8NfPURWysGY2zBrkkQ+NA3tpkSN61zJA+B8nAfN3QbcdCcok
tQhAjWuNj81xwlTLLsWlyR8cPQ3zF0fETWe6Fhpc0RFzTN562nQGtGUvz9g74ywQpzxfQn6Eghdl
xjKSICilZL7b7jybAlFqDqq02qfs7Z2rqHmlQptgEePpDwOtNg6LQxQ7QkPrpCbn0ZP5RcOCbtU+
LyBnCcNZ/Y9egl83T/x3ZQ909cqpKIP04VEUVJSRHVDI8ICk2QmSxO5Fq4kxLZgSv9UwY6fZ+r0H
w/brNzgdfp9xMJriZlPw/wiYiFPR3h4yvKp3uqAw90Cb3FpOZrBF/4YRErl9rLTZcR4IJ/gIQVuv
lLRcrtRk39mT/qYsKrByqDIC/Zp4B2IiwtDppmL/0RQasLzCe652/+MK3uUEmfTQ0OLTPxAHVovz
BWRD3vuAeZZ0OFHsy+9UY0n8LbtQNWD+KBhSuNXIEF+we52iXPaH9tMt9XcZb8uBvkTwoqjZjxmc
pZOrNvQ0FZaNQSK5e46L2T8uMBCT6lOB/tzNii2l+GhDTZmQnY2AFiYIPw0bA+1hNy6ahezezI+G
tmN18ID6LV1EfBQyQ20r/TkCmPKKLrnjg68El+9duvVWOFgYw7i35/YrWn6M0P3ZhkEc3WCKlLxd
BlsQ4pTe43VYPfxkMKTM7ALUvZLfc99iB8gaBytkC6j4LRvFzeGmGPoWfQuWcey197tU44UVarOa
/ZuhV3NauYDF5D63LCeoittgOQqRs4fmfA2bx2JF4cVds8guE1u9VBr41sNNRYL4SlFTedRTvI7s
JgJuOMCg3JcsJ4i7tegwHDmc/TO5FQ/qpjzSuizVqE73oyURJ0ZRyNqJkVVVm2Qu/F2oXN7tJy82
Tws5YU1S9CuVTQz45uEzikhdDMb4ZyrV17g4om39Ojjsvqluis663vjYeHKjojIDcUQC+m7Lfn8V
KocDu25jP36xMk9J917bzcaZnlOqRqWDASMpEMi52I2zhgI+NuTFUaOv5SyFzSPIeYCfa1nIaa2B
oREQWtaJ88+wjzH73aizdRWphDP0MoevkGn042wJm0SZr60dSqy6Pgfd8RmCrtIv6vUT5ol3ZcMo
DIcdirxRmpGmEn86Itfq8lN45EF4Ld13fZiWMoV22L/c89udRAquRKfnKqWYcyLPee97PnDCjBh+
ntL0oL+JZq6OElYX5S/WOGyUtEvvZOPN6wAN8uCi1F9Cu5TkaXhCw6mnecPs9kT//dlf21pA8KbC
oWuEi800O8a+RbdkslVkgxBvPNpel35SlSFmzBtvNKuPtncRjRaVIFV/wxExCf9da2qcXhE1LG8c
tEv6BGTqYfT7kMUuQrLAzTLpfCKTX9nE4dxGL197Bw8mRCFnFa5bxI/LN7CIeAm8XSRMmFikSzKD
qAKxeMJhijHmsad//52fwyLlKmPLT+MGO0CoLf0KOTnTzwFDnrb2dGpyPMGYCLbQomVbAfPu8G3s
MZKhU0cfVSdXe3hvzqfi1HYLpQOK1iKY7UVgyHqLW7gvNcOzri2UTf0rRhDYzdiUUDCGROwtAuWt
1s8cPja6Aj1hdfgFGvBodrEsziFI9gjM6lII+K7ilApnIOZu3X+lmzykSnS7AdFBsEM6hlNRnBqf
K8MM7wx8/oiZwWB0Df4PsXstDNHb2vLRtaGTrca9y6gmov4+4nS7lYEH/Q2ctlXh8IQb9xH3qKu7
HnPMA7QR7D8uTDtAo5FIY/AuMWL5RYg+rDS59T+sv9asTiWp6Mz3IPIYdmiKxQWLvHEHsI1M6oW/
X+1qA/OB0cXYQlzNQbB4MpEm3rCdh9NVEToAHoUD2PLSj5qoTfhB9bQnfZpg0wIqShWDcjx7FfVT
ur4yXe5d4WKCQvEtTR4tK8KaZf2UhhhuSDFpK5Cn5Q+Q0d6Hx8ZNIRigJOjrDm69//pTNJRATkRh
sNpUWzzKmGNU4n1fKVfnU9EKwZzQ0ASw74HgEGj7CVj5aP2moPuTQ2ukPWrS6P/067TrY8cY2lnF
TmZ/1wqZzju/II6uVWgHkP2wKPLPklgUVpEsPcGNwdbX/r9Vjovr3R8LAkkR6tCPXrFR07xFX+Lu
np0L6uYZVEbJUE6jf1Hjqx82ohOIzlUYfaoW8IyHX/g2pI1VNQBvMvM6Jb8HXLmkoYDUeCWR99OQ
Wd6GmE6Qq+pxdYFM6BzL4ZagcvIqY6JlzHY9M4ZOR1ckOdlIx0dt0sPycEYkPo7sKFZ/ChP0+b6w
hgJ2j3S/P7CrK1VYeGIq1iBhsZqw1xUftKa2nspfYfnQaxwfdilfp2kfLK1voqtKZUwUQl5g0CZZ
AWFnidLrz5sp2MD6cT4WV8SEyq0RkhxuuKsB5C7RumgcprFrF7+5HlcAiie8Ep0ch57XjC6gK9i1
qeLlSLlEdyrh1SCSIfhos0cwBohMEDcv0II2tjrVK/AW01/QQQSqZidjgWKj9Jbyl/CFRUNhjjyi
6v64m699WQmof4YWgjM36HdCRlX+72kXb2x7mrzazD8qkuTXP9o0K+NBmCr6/YTGXjrIvEOYasZN
55jc+jh/Da7GmETJki2xuUABfU9mDLzsRDZ7v+PwQDz8ZzuqAYy4Epv8hbqOe5gL+FwCwvdothcb
23nfsmFmT1yC0YZ6UhMK0JQMbRtcdBJGqBcSSnYTB7yU/RVzNOBT7eWZfrjZI9wFSEb9cgY1KB+3
d3W6yvovrnzN+tsJFLcVlPOs4TE73/9BKbRRQ2+F4eginw0+dOKWeexPZSUxctdbMw3Cb2DyWhoB
x5k7q1jnZZ/DeliWbmZji0tudI8e6RLDEkRs59V6r09olV0d2+W1uk0Zj0nuHpz9FRcPAs9/ZUJq
kkIdTKHb8JD5Yy0lqR23LaGvlc07D/RbtoIxicVgMoER72vC3d/1WvFJco5++Q5zi0mbWOIETXI6
ELBCgn7C7paZ5n5Xw3cHvo/csB4A+hm9vVbRvd4UJIa+u94hzoLNgZmgkFQKBkGtbDF2eOQqmY4h
ukXTB9u7J6Z28FOGTXxM3Vfb/wHj+ZcsBeFnmwViOXgyUGSdMeITm9NowL1FFhDZTvXPt5YybO6J
UgGFpdZJ9OtnuPMUbpATYy1hc+tSlxq13l3NJQBuQXLh3Y+glsAurYZP5+GdYLAbOx9H+Mc8ZSru
5SddelCR/T9OaoU6mE9Tsodxq6bbKjjVP0NbaeQbjWNWnbYv5SSMnV4Lzcjz6MxQwOliwDLeTE9s
twcEF2u0QDq43yJfPSK0r2GhMl7Vgpk5dLSqQqt6lYl3wpxG565mZYkrZWTBplE3WjDoridywa6T
lTjmF7hjP14hucIJXnUcF0mJ7zeszt6Czhi/jB2lakfypvkz66/D7BUIZ0NCg1HWSThGjNfNKI8h
FNkkjKQ8VoI0V5msaRUbez6+QOqd5AtDPng61vvVG2a0dsJ0XPdb8+saOy5zOPoh1IZYsf5aeyLp
jbi586LzHntqdiiIgSerQRHV3DcWU0aAbkLUJ3zO7f6KpvHiiA5B88RDuJRZ2MCloK77NwV1J1Gb
Ojz9MF092M6Jpl+U8r+qA2u7UES9R6mV/4ozmbTKXn0D2tRaD6iCc/4mVwkaIIOrqm2CSt84AhXr
duDyD1oKzuCSiZRrPruGdP5cyw0RX+uH3paW39UAoy/7PGWp54Cthiakoh6R3YsfnK/AnWz7FOKu
Y8A/0brKxN7yTDXA7TINyB9EMvpVnO7u/Ma4RDyaT4abxKYLpzfWZvx+uNLVlf+arIrev2CmGgT2
FKi6qALkr8wJZGaKY1eNXxv+1uwnC8zPxoYv+unjeQtsWmZtcyxlyqfz1s+L8zJWs7q9qUR85nlY
+e9EF6s0kI+QVVPNCr/zdXgX/fac9TC5lHZFJuMLNfZE9FBeyNpCXvQJOV+nmk+/fDLkWcgtdWdz
JaJqtBzFdtrIFldwIeTDYuzqVpSnxLoKRongKrR6NBCHDN2oPoMACG7UpLwsW2bv4gMVLwLH+pBn
qWPQae6Fsn6chaJ8elS7qjK/6FcPqHXRq+bkSMFv086H6EAaaF/0FJFkL4jCi/vggVqOQ/fsrDEs
GVniWRZGyPjr3zNUQdyT9mm/4ZvdnTRwHjaWs0T6dVa337EDdRmatS+dvJtUCV6MJjxIUrSFGeG0
b17sUmwDz1sxGmnQrj2+/IJLi/XKVYjMLumBXJZaYFpGVVMKRNBvVob0FyyM3JGvLojXXLZ0ivkq
IwcbRHbUOtj252hrpY7xASnI1ZjU2EflYZyT9X4t+GyfDnU9R409kdHdWAkEQiHYSk0rEQJrEY2u
DFgD+Gj6PABUSZDRlWu7J3hs8Unaq5NCTvxAgDwsXz7Oo2Lkws+Z1Pnp97pq+6ia5gmvGmZ/R+/f
/+EQflFMT8cQSJO1HvZGQzSmebmTEai2Wnp6vg+h24FeTbq17JqIyXqRkZWhfj7XRid1/9O1HDSc
+YKlJpSR+osnRXxhYqufOL8AcLVaLXT57d2VlEJZ1JlpNpZnuggZwtoTUbnfHQMbGX57BUG8fwGc
SH+PE065oyVytPFCnmWY8RbWVbleeODowJzWQd/LsKO8SFX8B3KI/ieX+PBYda4HV6VOeoUG5IKZ
0ple6dVQ+9+VW0Ce2ZYA4YvJAkZtvQkCAn+xe693spLTuqX7em3OttDfUFxPsYO6uMAkEhIAn/b4
WW2B0qpmXSLRJ44GXyeQXxJtu5RyXjIoX/D2zZlp4ikfojvIH3JlxF8MFenBw0HI3XDBMoelFFoE
KdIDaeOpkx9Tl6xZ+LwSqIIsa0QH72v5MDajXmgQjXb1H1lfDLgxlmDRCG9AV/zuMDk6zcgMyViK
dwMP/rWCgJHPg9IEyBakKSkB7ay+jV4vajKg7QcrFDql5VxvYTTn9Cp7EFhc3pxUS3ETLfJEi87J
5lCxUHLSra/RFwcYxlf7gPQWauz0+fXDgh6BBH+Y0Ay6FQIgWuWjQ/sOZrz2vWGgS9amHs9J9Dv5
SKa2PgtvzhC/Q7pIInFoziHb2BQWU2CfWue3mQ35jH+0qTw1eWOKsQ/kDVKNNy7g3Tpo8HqlOaN+
Tep6ufdLOr4njC5lCFLDUyLrCCgojJJDF4uI0uTerB64BuSURd/U8A/P9zxb+SXKODEkrv5SqDUB
O6q4amAWN8MO8LC3XSQ7YVXkzg7TiK0QMmJN5zRtZ9Z8v2CoXfZskQRaRiJHYbDVHGiEf2AZzniZ
QFQfEVrxIZWsUYPu0oFZAgxOQZA5CyCC+6EvLvylMLRFIX+Hai7eOBrEYB716vc9uFhJ9M8BGBMs
kuQFkeWLU46zYHhcUirKE7xW0dmnnzYmpjJoE5rB6+ApWWtabWHUHtGluuHnClxEEKjkmjrU8Iuh
1RVJUqgFI2hRMMaXxnWnqcBZ8dHFWETM+4WF80vzjDlRHdV8KKvXh4sBomBb7dEZ+ywIalzTZni5
EPGrsS3mRric84zW08+LlVOr/55pVBe0Tsujh7kOdPi30hfOhEzfHZEv6fUM9f1gXDrMKbRn6VHb
rBb3cRhVn//Xnb6PKFcgK1IpDQzXU8zLsWzElQs3d7bv6IHUYHRymTeRPBX9r0O/BXC4SOyjoYhg
OuE56h8SAbYnxQWac21AZoA3t71qNZy9rQc9rbmKEOvYjhHMC6PGBcGq5+a9ZNOhIqIchKIwSNuS
CnrWW4S2LF7sUb8m8ZjE2WUcQroqId9qFyBchr2XVBKQ71OaFkyEPvZRkhyae6oj+m92brRkRDQB
vFeQR2HqCtZW0kOp5JPbJBROHBmVjgEPIoD92HkBX8TYV3TA9dWXhQwlqkwNrkGP0RT0mlisP7Fg
7xpmHa1zfTc/Xc9lfTubboEpYXeXwYhGvL3AbYyM4SBC1ys2jzCasfOTDewlffystyRSBgxXiN9J
zG5epT6xQhKQzT3sKOHgYWZw4jjR6DKz8wr+toc+hF8WkjSnaGgLJa/hqctA1K4WNSzybagUWXqC
K6/vuZ5iqK2vYVP2hh3pnKxGMkNalWuUr+q3NkPZhKHkJ9aQEvu1iJjRtcbZIwsw34taMe+YTnBy
yhqwvaO4CMBr4YXmWlFu5oW7KxY6ydVsCdw/WvvE3kjAO2+2MDf7WtLSC4On6J5saTpxLhjVzHij
aqVYX8aiZrLi6C4M9l4p3BChc8X21FuqW/8tNjxrlwQN+Ywsm0zrzot9GvUPwQf318wicT5ep+Mo
9BdSr2izHn2yAzs9JdE56QyzM20/861QjcEiYYpwg0gv9m8kSHQoveJPpkYyYV0WExZjkx4IPKFe
T7CajAqFw+UMLcc2mYe+ET7bNoJAWTBmaDiFtIsOptEeJDYcL6ZCy8of17L7sWBy8W4gSC6jaSbo
u55ockk9xxlvBhAvqWP544+TALlnkcBUHvWVCgU0QHcnAvE3ImfbbTpPmffuGpIyZQc5ZuBnJAWc
xJVpMyIlUU8gaFnzSq5G6qIzKsBpZqryJM255q9qz8BfpGdsTq4+gUG6H555ihUC6BDt3/PTo6E8
KDqxCEETwifc6WXCzAq6WjvQF1sKGFpCwg3CIxyFGB1MlwFsgSHd7d4z3nEMziXRZg6k2jNux76v
eqRDNbFk/zI+7fKGzWR98XY4MO0Wco32Eb2RIW3mGFEa1pZrhbDAI8X42b4uqAq4qKMemBdXpVH1
4kNYeAnf4Bno1k08KV8flJAY1WcYp17f7iMQPn4wzgdjJ5RhbKMNGZUnv44wItea9XwM3fOU1inl
/DqJsub/YDm/F2mG60wDWjpStqENqcGZanwgtKYNJXgn2JiDaMvIQg3ByHfKit0Y7jhuBx/lfhm8
Go0kkF69xLILLfup9am01YQHBfoxKmFx3lT8sfglWZbZvAgZV+9w4C2tyXT3jWNGVKf2R6JaCwl2
hOXRh4iVoWOSOQefpx49R9FP7P4Oi1K0NP+euLGNhFc1EvOYJy1pOfD5WxpVSV/M8d3ohOMhBOzv
XVF5U50H7/WeoJaPBfLCha/2T1SJYluCUDIPJulJO0Mvj04OmP0AJosO3EbXnjnIZl2B8MqeNQKJ
DwS01YP/3XbeAiurhepYwP/v0x5wrt6QzsOp+eHruOat4eWENor6xn7I3yjIlPpLRcNtLnLaJ0Ze
hiTo/FuWR4PKnQUUAX2aOqZFf+0I7NWYUnjYuJnes9KDmbB4nWCbQ9LskS06ui5MgPRYHemO7/ly
iJTb8Pb7YRI+FawiDOCqsLrkYy1sMaJCZz4A+OPXAhGExc/TFIdG38L75WXdIjhMyHGe/aLX7KqM
XwA3ey5i5idNLNLh6La/8TdGe2/m/r0cH3J03m1+rYVePD024uDprcNzC/hqNchuBuvOvjz5LJjM
0KIFXGAFL5rbaeJKzzeunDoQiVm/0n7aqcHcLiVLsfVR3WZuljk13Qyo6ZgRkJcSJmTS34Frlk7P
u2FrlzfhIRhm2WDjAXkkNsq3vB6RZJNwwnR7JXvduri3diTBIyr/6vMsT4Q+Yp4V0ZKLKDvju5Ty
yKTEZSaBNb/fpYdcT9FSsMHzNfb8vo7Q60Negny7AcpmB16ntEJpG8b24I2BGRW93r9QxJWyYCxt
7DJl72MmQ5QJDlA3RyWIGjwcuH1sM4qF8Ie8yKdB766A2ZxTMlv7HOeHI3XlOTNR6H8P/QtZwINP
vzeCLxbbwgVYBTlVpwJCgehMdyFtLLn8IFwQ4yGpR6OyVzSvUlos/klHVmGe8AM5k3p+o6GJ+t5Q
rRWSuPWImlSt4P2X0E6fv+O+vJPhjt+qqkpWYkSTBrFlAgJsG36wblubiZxWdQhGOMpi1SThT4Mf
GqWVOMeEE4IA/LEgM5dC8Xm/hIAmtXRQJmfdVO5oHkWzNfREo9h5hMUC2YWn5E2dJ3/HdTvSHHoF
+XgELw4CTxdosn0klg7nCpyty3eQXXjSOtr7ySNJFZKcLXVsxP5urOLRRMWddn2/MpKlTGleRR9c
B7QzuKvoclzJkiTWV6Vjva65srbVO7NiVhIsjQjSaJwRMCoKmr4CIMQCjx8YbqijMQb5Lynep8kv
nSiPsDp2NCPr5yFcNY+Ly5S1pnw8nu4K1dbGDfsd+5DCqYqJw6LLAWqVtUrdWHJEodITxGslUiWL
nsqt6T3CHvYj4RZbuehoIpRJuk/0FHWLEUrE/DCAe1JGhV46BMf2XJ0J5BQm6YmoIWbYTGWmONFt
OIIpHCThhhncdl4W3L3wBKY0xUBzPPTviQBpzq44uh2vmkvZEvB2By96y4Mp9ixcOCcWlFPjpCzP
FGRa+x2UVotZeIvPBLHNiZCwTGn44NadqbiMRkp4ohP1YJszPheLM34nqEuJb2xQ0bK0PZxxwvQg
brQfE/RR2YSgUyLPx0cZm50JpoPLZUV3EHwRKAFRPDoMM5fd4Ub0KqkSsPrMoKBIE0q0ODGQWZ7L
VCuYoiNuqJmSpQHy0dMDjmEm3KO18FppekW7LxrwWBICIaTK9D+ASsaDyWvAEmY+eKV9xhz4cJVN
AOfAa6ghClJ1iuzI7fwhJKEYbHbRHiMhynYrLUdzpFOQR79W3rxwSZPb/7A94ciUji1lFfygZXxf
0N6QVC/UvYCIxAXbfOlWWDUcuUtXdJYRSZqNdfwH4Ia/1MZmufvJAioSS0d6eeZf93BG4C9ekiSJ
Zqg9UE7tGsiSj8nkm1ewzzkY3ilcy7N440TYGeaQNeb/GZO70A3ec1YWOJuQBnK6nCF+58G3JuXu
AtVHSupoOjTZY3wqFbsMXLTdTwtx0bC54k814tgifpuGwg6m8QsXZaTfydOjXFjUf4W+2Tva41nJ
og6Se4MInWcm0iphnpjdadgmdYfinKwpzIn0HwqX6Owc5cMW26YbpZGX9xbge/pikVMA/N3hEgEj
n629vs28SwTh9xyhQpm38lWdm4n2slE2DnWjK53YZY65cArItyoV8sbP3atmkscRYnAkFv5lIK/J
A55TgU8lTrFHR1FRRnGXIia5NHSKc5vsiagyOMHRuDHlpYf+4KJ4+xpxfChRSI1lW389seDcgbFX
iSXOHOA4D+VISA4S65GukW23tURA9pCho4Xnc1c6A5rxl4O1PhjrwTYJB0IXcYg2s+1qSUOhOIGm
I2cxa/vt6sMLGYWc1K6+dx+O8qAquOHp915DFD80NK4cAxxtqV6HNe9lF7RwAO0T8T0z08kG0Wuq
be9J0qF7+jZ68AhG5282yoq8+Xze5Pgyy9vmqnInH4GKhKI56+X5gSO5HrKUl0W0hD7UnB7BEtjb
mRlZYAuOjkc/4A/IMXj9yTXFo+O30Nd1as3kmm1Oh4OJVJs+LSHjcTX4wbP7ToL1auwH3O1Ptiln
qDTAWH+XSKjF+kP28F5XzxcNjJnbQgElY3b92pjZAgy9wZwu9VB9wcvagiqa+oryBq1P+fRcFSIK
uQDGNHAH73TraNbF8Pn1OJ8F8Cq02Lydi77onNQ+z+jmMPMuYaZwF1j0vwZp+p5db5LgV2pjgjME
R9Na7zVrbxNWXkTSBwoI4DQ3M15GlGBM+QaqKyvtoFNJnOCg07WGmGT8O3nyErGopGoDJXkWkAzX
+UfGavivNQhXQlGWEzqRaO9O0xvqcIeUUQZuYkwOkb5lBzFcruvD/8885ljOTzVjOq6rvfjWOPui
/t07gTAFJFBEqTCKlGrroZzy61ck/xI1U12tRzT/Ky5NL0XnIGl8LtbA04oboGvbtxQ0ukIgr/jL
ET1T8yAQjO9CVguEcfUTOojdnMgfGqX6++qtu0APTOMYtozwzIt7KVJYb84SAdJ51wbdqoZRWwTI
utpvPs87gdyqFN6GpfjArTrueYdX4eWZrTr01KKNhbYYRRcWLKXc8zHzMhWEOS/1tXHTUjUVp2w7
Wwp2O8VB9QFqPIBWSWTUV3F+tedV9xjI2elPylCOE3YhPXs2fOWnjn9S2seYCNMg8plx9yQzTi2M
ar/LeyMdmYMtxJaYxa/ifpgp6RMsQ/nEJlQsB4tghnNVEfnH1kiIWpCA4hLHSEoaGHEFMDQKrVgg
XhYEEcAT8DwkLsDwKuGQf0CE7eul85aOEcWQh9Y+sJYNf3KK8JowMjX25E24eWZYQv9bdPADR7oW
jQDxpI+NuoCGaX3CMtv1kLXb6xG0lN2MWVq5E6Rwwbc2xD1AI24LOVHkUHhtA4daxssn2SChBoyt
8iwOntjTJmZTA+rjfkylOvMTiFliBESJrn7ubOiFNrL5LaPbS0lgDGgolWNbZDju5W6bGLS3RC8f
XN/3zi8KQTPAWMqeYVhMXYgmydEXGJvubXdge9mzgoChFMGfl/OiW3f4V5Opf6WpM1WScWxjH+9F
oFzlaHvNB9zsdxfeYZDCbWUD6xlp+jBwLC9KdM3V/YPTQTLXLgPNUbrOablc6BuLD4GwOLDkujnL
10MXkl55rjUnTFBmteoiM/OqZqC46SlgpaUMUv/rkkC+NyCGTGw6a6e1LrRhjqnmljF72L35oQBf
r5uEVEwE3+KPdOCjbjAzxxIAsTelb2k+nGrYKlX7WugUHlcBrm9zbzc0xJNLEVegRk2iA5gqI89T
LT5sSXpoMZDx2Ed903lWt9PAcDjlNz3cE+s46Y4IxuM8IJxzd4wj8KlE55gvlNiXNDPSU1Cy6PaV
MbkK0G+sC8LnlmrYa1SPXg8V8twCLFC/miDI92bq7kDtGq56IBFo8tociXz17nX0xzxjtt24ufMs
HwLHjlGtgH9C7xXmWqlHtLh89fvJ3NETo9yp/CHCeRQIEhiRmPY07ERas/Lr0AWIwV7WX38IKmfm
gP/+Pf+zzbR1X5NNqYAZDs1+L/pjWdUhu/NHLLoIvuYDANkRsecEk6WLm1C5mGI9K8wFR2qJTEws
KaOOl8HhsvMRiOpPU+6v9Apm1Dt5jnCzE5RScKQybZMNzBUcjY9hCaUCqQQoR1WGOXBxG+53hVO4
o+uBvDFT0Ghqny5WVMq552t1jMKfzc8NvJ5HkYVYDFbWkpdHI2lGX0O9yPPXJYJGNjkSpPHI7Qa9
6Y87QeDbpAcijbmNeHsQu8HVV/Q5cptuaySvUDfl9Y4BGHTFTsH668P1cPMD5UWgXw2FqtulSRZY
uAGV/eqGUEVo1PON0usFPl+/NCju1LFczxx9RRTy95DkZTwdisP/K/PBt1I3NjH5YOJrnx8v8y/V
aSYeCItTexPRggUuw+FddRXNg29qmEkuftAV2NuCcvfsH0BsjVNA4QcadGKmFzai8bgAAHHxvO1u
xCicV755GFCQbH9zX49hW1/75Lxi6/RmO9HjoNkv2CDczsmPZsPOiHIw3Qu340SCJsImIEXgIfYc
z7ED7tNk7uS9S3MEAyIysu+xyBdX7sw1+wTcAnVShsWIcGzTqyLyTF3S7OBGX4U04UH+oiHQVhYJ
4uTJRqMFkDvykZ9DuHoK/4rOASU54irq8d1vMffVIeNxHxXILfXLFs7rhwgWS0cToEOk1mjA4nEv
qupIw2h8th6tdPVy//rDYHqTLadnruvX9b33F9umGf4D9Sco+60ysQJmVjfpk1sze9JpLeahZieC
Q0hlxy/aFK0zrQm2LQt757IUiLHtojQg/ewLq6QWRkhhd9cPo/rJ47jFptO01YfRbuKX+JBgpRov
XUshmCGvjmzkXOLh4XprO8KHkGvtSVQq4pEYjbA3JpqWKTO6cSNOkxpEBEHE1H/OIwy2hPvFoz9W
gyXegMayAm2j4MD8pFY32fbUtXZm9QNsqiHIIngdCITWjOK+4u1S/dZWnSoV8FR7ua36jKnjooqM
+SiV1QW9NUrhZhnQTVwm5HzzKuRmlXC0cntz3td+7zcQUkOzDSYKKpVsDhCwxqYcuSqijQ5FBEE4
hxPoHSZZrTkZ07FXG0r0a23alj3E6osDSVqV9v+yxzOKTa1DxDdJq2Zv7lnG+Zb/urdJ0/JAIG0D
GqBLMLv7NWy/Fv7mzASAAT3i4acqOPDG9jiwR3OrcqjOarv+HTN2tk1WwhYRSiNUb2929RYtpyyV
H7G9pqC+T1/GXvpr/A54uYnw5e51jTKsdPVJDAR0IjxXxhDVM//pzcU18uYaW5/HnASmejGDWL/M
KI6ehj0g1zp+MO8r1AuM1GDJMC/0f400UCtWhvs1FVBgT18w+Ha/rXLrteH639FcyW67GAiZCmPM
9jiJMosX69NxZZSinO3XVfRCIorAzK91TRZl12+hmJy0I4MyPmyNzvKUcX2y0aPX9pdFzlFSndcG
FmD7QbKIBS9R6uzMICFF6+BMFphZqa3qoj1CnM0WZIzU1iQD3pOH/0jw9g1yFS1bPpG/rcDVu/ln
1+C8SfuT6dkS4piu/adzFwTX6Sq1M5UhkNMmZDHCjOFE+AUHH1Z3uua/4jhnk/S8K76YeCxM65r6
VcdEIrVXQXFlfObt07Kqf8wqJWgghQ+hcIb0MzXb4xpL3bqTorbYKveulJDJkC8hzwGK1jyHg2kO
o7ezMgZLHGy6VXAZZ9Q9DDWa3MtsgN9IqwjVua4QUK7El3bmurMWXv2drdiwbBLjpVN4rkaF7u/G
8K9VQlcoqEnPcLW3hM+SOUpW+qNYyksNdTqQHhqnMgPGTM1Y7wPtfs9fHURYMHX1rr2vx8RXMiC2
e+mVHcehsb8tBzJISSY/pJD9vCyawHq9+wu8fREFSDPcHnz9/ZnPNy4ZVaBDqlIHSw9QByuRpB4d
J2CZx0i87LDu/jXbw4Y7NEEmYL8G3g6aTKwzUyxnBlmc0JLKat+A5qhju/pmXxUWujqzheJ8udZK
vg8diABrbe07eIKqzgVPwdpIdpUozKn3thGAaeuMLtUd+hpnjYhgCZDxrvNTatOaLCPwWMuE4NL0
jSwZGpiiAcKcWN/AO5eJY0LRSTolZnnelsvKAQaFonudqk00OApQs1K+2emx6mM9NcLPh/VkUTuq
PDV4MFOQu9rQIA+devVLz323woXE3+mguB1B3EZNTlicnUOCiophMbjLzUf1Hw97eSHYwa3Yxw1W
XCaiCbA7wJJwKVTtbwnBA9mKTML7JuN6HdbcLMsnCRHMn4c7EGEh2e1n6z/kIjmb1YxaIbmUOiJv
TVtFWXNsli4euFxwoomnRf9rapXfO8tCM40gUJla3cOVaJUgRspRjEpodSjJvU22vFCCeO4H31o4
S3UlEg04knr7qdLnUcIo+ig8DyJZWN4G2aWaGETPJOGluClSIge1l57VyjJ18yN/TtFlxqRkAi67
tJ+IXGQQn1l6LA4tG6GmajeOdIPsqzri/bQdKZmY85IDXW0V+55pCv47pWn5QUxePetr/KeZ8yD0
V1yfWDoMc9fQHHReXdy2mo0WStKHswB7R+b612QnS1bittPs5DLuZqIi36LSWs/KevesqN3akpwR
wW9MTrWOFAcmTR6dK0BoVSTHmirk60Aqt6U15MN1dJvXJF0QJ2NUD8h/cQB0aNa0CKKxnxhfta+t
F9ouLW/2IFwprTvyOeqJtABBQIpx5sOFC//+yBmPRK8R+OQ4UjAha1RoIgQMSL0yhXjsVy1Fkn0C
A659BNzAi923qFsjrtVy0xnJU+3dU4bdIvNo2Tnyvbvf+HjmuA3LGu0Fy/uqOcTVLogZGbVDjmGV
zkmVzSEnjqcqxN4JTf9Mcdaw3qcV1MVAUNzQAd+q0NExpoZRKkZzuV0AccIwtfWxHUZGyzYiaHxT
faD2nCey+EHbOdwxG9QlztBf9fkWDEZM33lVK1ZtjE7NFTSIyz0vjLCSOm3GA72irbuy1uZBrBWB
BUwzS4mqazJ4oKME7jmvpjCcSJuiAo6YD/gO8Ym3uW1So1UR3wRsRj2QJ2KNMUD3rDOxNIwGd6Bc
gDSlPaBnQMf0FdD4fIKlA/chUey1DpV9SufoDoSYz+bQvV9FfG2xvgoFIFw3jDUf/5PMUY5kh/6E
pjaxxmGotruD9kcLlnTJY8yun9eawQBiFxgOJArs1DbbGFkNcA4YnjCpQqp8/jYvayII/WCRpz9v
/cPh/Nf6Rxp3ygRS9Oz4yz6D6q335ueyTiT4cNV2dYraq+ebWcgWhkUyLHuGZaWaY8j+i9GWBk6m
FoMjsEHbKCZ5phWZy+sAdtckoq8ZmCF2LqvggeAw1o+Y+OjoFIowFhBHlQNU+WASZ5XgUodIoZqN
nsg12ilzxwBN/dbmXt1PCC7/o4HyDbaXfo/QtjIIcqW3eT44r1Qs9n8I2aUXE0Xmu0cAFasajBzX
PJt+aEbmwj07VvJyrEqmfZoHQLueqFQcBkRIq/Metqx3e0VJDeB3NX43TVjXZmLTG7wzPW1tgP8M
NMSKee9RzCdb3ql+FCdQssSPv8Ox7ZoVbDHiiu4D0M8cJOV1UaupJ35uvOgpH4VjZNfOBCtLnTQ+
XPWignUoQh/Y62nx9hGObl63ohiAZgyhNKWRu8HReQEWV7vynrja1Spqfpmd0Ro39CcAaDPzxHaz
KhquwTdHjcpD34Fct/ZbpybawO+UIBtOGka33gq13vvFHywtTdjzRTEieRIuGnxLJN5pU6F+NaIJ
dD13PZJ/f1TMwgl3k6aDc7gcFWy2ZdBgsYV+RX01W4tcOsmZZXxDU6AMyX5z8527H5uo+8pR34vj
7jKVOrkMfkdc/7AN9ssoXN3qRZz2qlnsg1r8e3XDGcmbVyVuD8A/L2mzM+36Tmg/obzGlUuGGo9B
XBcDCqdp2Jz+HeIPG6eBOF3VRVUV5IVtkxKC5FB8JxXYI67FyVOVKp3Vks37Ra7L8A1F7LwcLSjD
eAiJxCVJcPrLmfYYccHBm4ixSIRg8whD4eLBldjZpAZaegPlq++oENPr42xvyEG/H4HFFrOKUHw4
IhuPNywa4QQtiD14/Ny/P8SsC5evE3yOjPyZMC2WV5EkSBn9SlMtq2RBdqdaGtM5RXzl1HtyZyqL
LX4Ey56sqzO7tKoo14W61wxFpU7G51GCtpn0ZcFMg434fykKptD9tQATiI2kq09pvLxaHBpr8PNJ
7hfZr/k2FSjo2v1SZc8WLWRKBvFcl4GVuJBSovsMlX3D7Nd7AcTWCWJTSk7KtScU6hmxYNSBl7VI
iKEst75nodMr5KrXqyzIvohuhlCWZffbpBwNtxW+Vi/mi3BF/WTdxnv+uyq+A1cQirWvPZ0GMIyd
07v9fwLs43Hk3SykCu5I0n0nngjZWoqDyAiFc0v4JUAJOOy3OF3VGU0MtmayPbMSqZ7pxLD8maKe
q40r8UxqmJzpBHB0mEKC9A7qMRfSGgp8cJf2NF2VGU6/qaQ+ysZzjATK37SY3mxgYJUatW4tx91x
sBLBqRFfhgXgoCAishdSTtV18eZnWrgIxg+zlN/Tp8wHXHCp2JDZMsZBIjw85rn1mJuhV8kxX70q
fpn7dMlNiCCT//Q3+mVhr/E8RMNfNIE+WbB4Aed0Tv1rX75doSvil3noX5BjeuWhfB6ySFHTnluq
J7rah1jMczud9z/tYGv9hLHsJWus/L4CE9lcUH1MTTK0zpZDM+W8zF+24c8I1ll86AGPY54N2Xcc
3KRltXflRkac9UEk96Yu6g49mMjVUOCzuqWGZffrbZnPMKEJYkhaHvlVT6SpfUGa1I2v0wNU/yJC
KgNIwrDarP1LhfAta2DbEbWHjNo4POYA+d6zCJ7ikJjVfhVkfYFGmoqlz6E5bIDRlYbdjt0mip+V
MCJ/ndEVXv+/XPJm+52kEfJdo9dNImrYBIYUE/xsjqwWhdKbrw9S3XTmBuAaG4lkiFkWDo0jmfyu
TpTDjKEYMGrXdanpwgdwph4oetqfRMNiq9hArdoXPei07elUSkq2f6Bjq/91rhXqvPZJ4JNRGANK
CJnPjiylNIyIVPOp22NaKPYlbC+hzAP9Q8moRp1KtfLNcd+aP25f7uQJwCGr+xqt7+0vJFxHZGEt
i2nSVNZyrl8exq7bA8PqKO9eCWxJH5zmCeuPpMJh2xOhBd4cvklpjCoL1VsmCcxblQlvFUcF3tsf
sU4Vo4VAWrtGupB6ThZ2eXUE3EiPXNVgJWZjeUmlxUgwZyuyYBBytcP6R4i2GvHJfAn2EuiC9llZ
4zgcZlQ/12SrDiviCK7HgOoPoWgCR55mKAmNSCzL1ilQ+gJSgv5c4/4reIgzrrHMd3EvIUmvQSd3
1g3kH0hmFBSRM3hYvPR4Dd3Xiuf/C1o1bu+HLukcYW5A+FvvnaHQGJMg2tqUvq/Ns1gv+s7mIac1
E7k6xxvIIW0FHQqT+OAI7JbO+aELnRtTEj+Pi2H5bhyaGzYqvdPlaMupwd4jfIMFuuaOzDNzLTID
dHNyt20tZGBQSIQ98xFjii+dqTBnK+asXs94LXqtJ0VhgY/y64YoWBXlLIenLxa59MOgMgdOjpYk
9CNdsiPcyzoZmqrr7ZjqQ275pTAMc9ebu/QIN8Fb7KYUeDl+8OFyrfOGSbYTKvSFw1AuTp46EK9p
cjSsGKwcSwaUX9gCVapK+ky0UmrLAAtYAqiTxTNhy9NBhx5BhYypapxvm+9JP62CaMuIyaLa7ODJ
MHv2+UIq4SCI43ZnK3eFzYLml5+h+qbtMDgiLp0CpdDZ+epyqsidtWIHNf0DJgewxLbvJluMbHay
upk8vcUaO2ACtvHe0eXkUpgEZff9L7IYXsVxezGAoBpQ6VI0IuampvtmV640LpscGSndAGbzR8Z6
q5o7z2tyVPDuWu84IK9toxL/h0vP1Te5FxHclIM1jfgr0ZXr1dyprNf3G3gGwJ4vd3kmwobhVNkn
crOeUh/ttHLfgryXU0GE28YENwbfc1gmSTksNb8DRNEBbBp+/7I/YEENzm5Ctsv4ehVt6cZJ0qKv
aWaiO+eej0a5YTFkGABrWoJJE5EiFueoxoORGJlIaaLKpm3T3/B0eUpc6t6CZ7qJl8z6HBDLjvDB
O+c61m0npc/uNu8v0OvBfBbMkkCoPwUGPrtmjyiRvirsCH2eN5dCoWMPabjJkdJ9JFVRrQee05d1
8H3yFlxRRUHf+AlFrzA5qJ05qDpXOe4nO0Z31j+5te6vDudrLo4zyoYPYjKl+94haj1TZBU3qLoJ
9Cj2WVJ0oTj3KjOaK16MfYz8LbOj71DCmKt5idOGEHvVMlpnV3TfUvQGL00wYCslKpKDyuc1Lt3O
j5atioSZIPZi6UKHo3AACAhjdorUb9V1ZwHlWWTZ2YM/8eC8nqH6xAhCwOCPy5PJnW9xct6UbFJb
Ezg5p1hHcmXpgqiQeOjWKZ1woDxw9JL+nV9JR3iwhK2zlUVlfkxzEFATqQqxwKE4cvShKueJDHMr
ZDFniSEsicOv3fvhHXkvX7uoKWgM2ADj2WHou671H3B4CkjAl7hGpfjSmO7me4Pgs/xX6L/88zm9
be1BADSBTtU+bCv8v9xdcm5Y1crtCuCBKp9sq7qO6ORR2HO1wV+PS3+8Nx8CaaAcYA8i1+90ueyh
DtuipWo5QA4AC7RAFwsvqmWURGtsx4kV8s/fjbN3WJdZdWW0Bi24cUSWbEhK8v0qZV1wH+vwFVi1
/v3UiFOBVDz+TEp5+PfUpdbYJsJNcKKRPP7IRSaUMQOum3888jwVpTWnxzX2MxC9eKUg5cVb/Jer
JudyQScxv3Izo6RdIYAK0gHEP5j5t8kRhOTu5kzP1aknhXWmtTFuC2v3yiw6tjR1ZrMaQHuwrtcs
gG/vGtnxhoLLVwh4NqzXNaBUXjaVRwBl/yfZMMinhR4eNe4gyVdmqETSQeN9IvDHMZ28gdqCxDvT
mBgYH+yhxtvJW/g2mBHd3zoH1K2kTptDDczxlNbHYI7hXx1ZVqlecUHedFjtj2H5SJRbHN+zyHSu
Wq5T2SCOVoJvm25h5kqIjMt87/j05tzxykKGVVPkOzek1NMSD+VWVUDNieQv8kvT07KuyWdsb33+
qE5f7kehWVvtrBJGyHeGmAuLxOlTGuATYv2faIPcIFmf8fmzy46yL0fAfKmwWuEyBkjTi/185C8m
PvptEicUedbCqwNfp4v7BEX+nLtlzFyrR890bYWWqPja29NqVoVh5mOD0hxldJxGpYYQDxNKPNvc
by8YbAPYZ0EK/lvf1E8n7vznLTCZn93uDNpt++U7WmnGjAp/3J1lAZDRjGFCfQao2LzGt2LAxeNm
TyGQPyQk+RrInMn16GSCOAr1SHSvdgNadzJkA0Y8/wJYfSr3NRDMd+dfhW2uY4KwTac1L1GiMWSx
SwwjxFZZL2YiBBy+0NM1fF2vqNeY00vqmetUzFNhz/pMgbRRn4nfxfNpcWVkczEgZusPbYkbCRTK
9pJcO9QVlo8AJA+jqQ9KWu+DpKwVtgcPtpe+hxKNXujqOXwVYRNzZKFqnnXZMBdNOQhRlP1Kzbcw
NQSHVKkKHQK98/onztUBjigKvOV6IIftpYKgvrRKtMy3286aHrqbNzDk7XYtIHOB6lnUyycMUdkT
SpymJjtR5iXfGLCQ5hEw3BBBpleTaJoiwXnbveUVMa5pr13SMZHLLFlpt103nHDF3u6t8tB69RA8
BF9RrCBdsTF8BJvlg+yoZ60o0TrZ2OOTFvS21vdS97utcqQ+nWu/Wr5Hiten8VFkh/LB060IeVWt
T8OU4BAIfwZnEEef5XXBwpJ31hLTLj8gZ1ayZAkOWh0UQOZUi4Cg1Dy7g/sXUeuAubu8trbMLp51
qlPD68QGs6WsrUSNL2R5jAktCtYVjlgr2E/vuUWs/nLlnsE232dK2izVqDexa9R2GtaxvxEG5Ggy
H64/WaT4mUtYA5lUZ4pXnyq6lbC5MlkZOHeACffMZZXtYF1rwdlbrUQyxSEmQwvZK2XFkrpuuv1S
KEyQVBx1SfDqWKDlvR0xH0U9jHQ/q/8KTmbV0kLUSShBEX7j4EBuAf/qDh+NP3b+q/OmugtNYhVy
p68ArcHjjtbhX5PDVEYiWiwtJuSIBqO/T7mB7VVYJQpeCQode4/EWbWAXa+Wx8ik35pqt/3afqZF
YOacdMLKZvwQyd4rYmnqafdxjLA/xG7RwLFC8BZ77+e/gsNbwi8PgX5Rqn/u9rkBDoVl6dcCxcvO
Q+SpIExyywuHlK7VArlbAdnHgASHD1F5EZipsycqFzFTP1/nML+pIlEIEuBkBp73uZcXMtI0u1Xw
BV9bF49b/hhep/StmhTvJxTHcEb+WKs0skQqj6ecaIlL8eCRC48zmpLb+AiGrfL83fKEqcKFaxh4
4kqO3xcterm08gIJH0J+fbz6XBsGRsSFEXFjZUOfEb8tmb6d7WiE91P/AYMg9T3KGqX2mJIoiiod
RawXaTLTChxww3G0APYRoVMaTkRZBZAMmMv/igN2EcSYnNMZAQQGIQE5JptHy1zHZMtgQMEPhCgH
R1JWBA46Ai+EpiOCDhQGhQkPCY624aXpT1RL1zBbkQCVpwdUoQit319yXcbm8uO2pYar+H9585VR
nT+ijVioR1MkUb0FGpEah6dl+Of8tW08jAlwCc3OcEAXMS0p4qa1NJOGZ4y8LM9hIQW2Okm5c1om
KyBFezIvShflFNmnXXlU7SdFl/Df7FlkFMBOcVqV5SmGScJwjuasrtUzdJsVq4d9OVI2W2R0Lt6m
1lF4enf8BUftNw6s2LyWbbrgE4+rb5Sd1FTpeebPHhh1zxVBD/pVtmT3hjGhrH/LswOsZZrLyTMF
1REeu1H0DWj5hLJZxjm6ne6h08okM3mzjCHG+2RJ5mUK+iNnu76nKn2ZZ1dP7tJG/fTQ1bjQ8Ygo
oG/aOoOIz9jzgdiMit7AP+EfYFDhetxK4ku9YVC9uPaYXCcWQxkbvgPnyuGy4su1S8+TICDFhUhk
H+93Y+P7udMXvm2mbja82ZmFQitaIoO9UOdpsYh60fRw9u7tgolA5KsL6tNABrkspZW2WOiqyQbt
NJRx4fPo+9gSHQTs42mD2cY3Np9oNdueTjERa9OVcD+/aMphmbX8fKJLoiiamyqVNu/Sk11FJKHv
yVvHcQt9GUJFBaX/e5xg1yc1g/mqxUE6RvU8i3b/XMKMPCu2W1X/dBHuZWE93uvsCdcX6WLzB+nK
/G2lmRGOJ+5Zflb11Rgd+Vu843ICCOrtYIsAKhd9FSW7BpYW6yf1UNnfGb0HPb3GzTJWWQDmHzvB
e7GxbNrMJAwVdLF8qhi7zikol4r+3d8OXz96pEaKMEOnBXBKtLjK58NBOoYPGbJHCn3LxUODUxJY
s5EunXZEj324Uf0cNHinzM1j1MBBhqwrxmBQEDszzFROzUiKNjd4RcdRjVkXGUkfAWiNIyFxr0Cf
73bhfrj+8ad+HIWGoZfjNANOlTcCNKtJvrcUSBUDVlmoVQZcwNsMGduuXVaFpQv/VzsdDIz8zOjw
3ln6eSb6ObXzXBNWq0pk7ty81Gevspqu1wl2YxRJelCkNVHrBDnEJQ3wGHADJ/qc+D+TvlALswq0
kZUkrk30+BRYd4oRoezR8qDL70h2gwPKUR9p8BEJrCFzaOELHqyik59P4zu6L43CEMl+pBcZzZhA
wDkjcUvRfmk2sVX7pBGYtjqy468yE7Jf9114CZ57qgCuqV+It3lMb+5GPbpCO5BbUBxdRepTJPxc
Odr5jfJEuTo5V/D3+MGbO9Y3fmorbmX1RcLOvzTAe0oe476bn88HSRjQDZnuhG4Of8lbCYJxRX6z
q193NQUkHsf0o1z6iiTAKUICEErfIegCisBRYtqvzbMImwUWTEW1v0zStAADvBNuX2tWnQYqnlRc
pqlBNzJJWUg574tyOGe2l6zkq8QfEWLAKeEkFOwpO4aZ04LZrosVFoI+n9QVQiGUafUEJDCulPkz
bRHc0s23CK5vEE+IPFo/kDCr9Gj5DZkK/qB49g5ezUG/BhSVdOQ0l3w8Tj+go1nHqtklVUPqxFzY
2XbNBrg7CDIteUMdpWWDXsx2D9ACRDYtgjq9MZ7ssh/EhL9SC/HE7JkLUh0YMrmEj3daFvqVBGlM
BFbWxqPBj+aLHLuI0i169Y0Eej3XHZ+Y4xFi6U5PAbLuLmaXBjFvoVLtAxJY0MppDRJKsxH2LzoQ
O79Pd//1VYTi0uzd9sFLsBOFaeqpbTcq4B3GThP7NPf1eARZhW03476au/rce/+xp1YTSdBtxLRM
MUpQs1cQlUtbh7LkyFLE6rdg/4bjIgWdDh3nCPaqD8engcD/naOLT2BaJ67AhWC76suArxwgnWzu
MkUa99NmWgks5rHhqEq2xOcpaA44n3HXL3Zl5sleLQfIv4Vv5jdkOJLA2Xgdc6CTeR/SUMex8Z1Z
lCD6aeXboJhGSCxRy6Ibo6t8oM7cP2y3iy5AtyeIZQAIrS6Qm2btrRq9B/BcG+QvdCKnf7ybWKWz
1r1U+C1skMnBR5xurb7e79MUmnDnSciCEjj0+pW2gE0FP5ttSxfKhr6bhgsCbMhgAkMXJDu5Uovl
E9NTVkyRz5FBCBJhMDb26VhL3EFHV9EBTifm6D0AtLS76EqtmzLvpLLTD6HJAt9QatRda/aAYHuC
dYJHEHbDIfTQZWTtaQzTBUvSpvVKOJw/36ma0h/g9l77aGo3c/SFDL4G2S5T6w117F3eSc3neHPb
Ls8s6gQeLT1vc30YC4l9rz72XIkTkIn+2YU+RgUfjf3zCoweum1rCNtMCCR+ns99gQWqZzl/R7Qy
/82vt1Yaw6J/gWusf9KfaXxPMkpDw2IoavN12QtqNKPUoYyQUGrrAC9cQZlQZEnefp34sggDhUJb
Nl9SDL5nLH3S2sqsupdPITZYYbl4qImfGnz8dBrV7pa5SbsqANzBoiFSZNYnhgL1aZcZLJCpmN5O
reStWNcUanXWGViCKn+ksqt3RsqKGJ1dJAwsiz1z+48375at0Dn5p62ziaDAtHpAHJ0B9mE7Nsa0
noyOB0ClLp59re/Bk8JL3tonhAU1aTSjvo+SwRSIo82XZeqPd+iNWGqMjRrNlqA8aIkBfaAn3FE6
emzz0ij6XUtk5u1cgDnpJ/XkzsRoR8ZLZJqXDXNyiGZCYdmSGXnFCp0wcg8NNcDLV1EPVzo0Ez1h
oRZO0CKbrv2YTEUa9EgIZgxaBsbxW/DLpmRZejI14zj4+Q3zdNBiB1SmUjN59ewB1SylmjWO8oj/
7FkGEfrobpl+SVx0WBllaT0jPF3XFjcPvGm1kYQQwfQ9wvnSLV2Jeieh+c2zXJz4kkb+N4qRsQvX
0T2Tl/RvgtUCVh31oLinTinQQJqPzqlgwGg5lsmRtyMqcYcIkA6DwCPoq0AFFXUpPbRSxW4aIAQn
27GyI407DTICnKjXpBXjM2KDV+LZ9B+ZO2j/WHWmz6Mtc+X7NDNNYkk0SSeWuwQ0GszbnQKXMrN/
pONYqLO3PwYMgQMZDfaHaA4K38tTTdpE9cbg1t1/ZgqR2FxineFjo+I6PzI+YdxEvdBoxxWIWbws
5LlWDdDrvp8MOZroGrXP/oVz/pmCyDcFF6kptZUwHeeRfvIqxiXfQqJMuM9a3rqfXHCaTdaQ1NHP
TO3FTR1DdGgQf2hnN/Y/DVDr1SMMceBxiztW+aLd3pp9RbkUqXH8X0TFPHXa1+rC4HpkJ1MVJMl9
F4FZ4lQ5/XDKOXEaipoX6tW835NApSgcodlw/5K/FYaHNl6pIXDXiUbuRzIUQ1MS8Cag9GnrWKJU
I+GjYYvZ6lZsDYALYdzX2GXPrHDXhmlu5v7S7roSzSD8TmK6ClS+Y8TNWfN1A43iru/NTvW77Gbu
A7wsf7HXzyDiYd5CQYVYZERW2bea60qYPqssISToKXqi9DUce9pc1/l6VQDKQDLQwtQYTeKPthQI
AvVlDSXCMuri5Wb1q/vrQlGRIOAQiqwKZZWhDbIAdMduX+j4sRivHgLknD0opibYRQmzakWT4A8k
VSDxmv/JmOapvPDXixJ9g0Aq3JGbQHZnwA0kaZxA3/NsXQBXW3yPS7JAfMK7Lnf7HFvvv1a+NLSF
MzmadN03xEFtmVnv+2u9SWUMupgPQLCuIMzxl/wISj87YXEDjpDqssWUVTDWVTzmKMoa/E6MRPIB
gWcA5gczdJVPXqPs2YmQ+kTyQpEmsANE6wtJQthcCOWVziwUhmod4kWHkY1+bOEE7a2zbAhNeOPq
G+GTQOGN+1UyOU+pIMwD8pUh26JvkUfnJbzk5OZyLe04lTEXkGktQgEY6PbwCsiJdSB+QTYNEaIO
rLFb3BXh281BNCRNOi6SYhRBM9mrgWGBkSGLIIPGZo9Noc3hUTv2je1s3xEXi6rzucXkMgw4Zf8Y
qpDvRnHzsz6jLPLvJ4hQvEII1bBdwzWWIY4xmRRRkd46c/hVhJJjdY7Jo/TpFZ8E3iJwTvHnmUO+
TkUeC58sY6Q3/yVpq9qcUzwNc2XW5IzyACzFaBWnpRdXY1bykJJF6gWe01wx8oMVmoUT15ZxMk92
fHCRZ/vERpKxoqAVIJGKYyDhRhL8/8w4NuI3tEFal6qZYjhHW0dK+yxOKA2sgXzO81+Fhlz6p5Hu
elC63qCbFpFReSZ8n4Fp0EAYuxCkXWN1AcCRIZd1Tn8ghpfPqx+5Y1QO8zK0C2n4d0NpDuooE0wv
dZg9pE9h0aCeFN9cBertnHZEgD+m9mf+jE9onnfklSvJqvS8zOKXhAERTsd63zZUQLbEN6aMXZ0k
oqW2IDQ2+d2D83lt4hZztVmwiYbH5aW54TE+FvGvaDuUNl25BQJoyFeiVmYci9xOsPEDFAbKLxAU
L1kdBRfQFWZVfTd0ysDMjXHDfNDSDwh/0eTbn5xt9gf12/A57UC6OZxpNpgB9OlpJNmzBPK7amJ4
8YXFM+gb1cGL76bjJbrTjndXPr/B1PrRmMU/rrqkCzRcBlbJ/+Lpvhk1fdJe+uC1RDqU2wr3V0K5
GoVOUiZ3bxdcdnD04JECBXDZeT2JRNNZ0UjfFiCDt/qVmnXobl24jUUphCWfgTi7m3rP8H6bWN3c
b8/J89rbb4z4qV070RooyU7ogenD2l7s6DhRndNjJaCgwYg4BJi1cKCsJtTa0W68uziAuB5pfsJj
wbTmo0csIgE5DSN9RyFSvH5R/2nrZgZgRmemi70PfmtfxpVTwWP7TpLIN4fZEZeaOSCkNIUKWFws
JaNyX6N+ZXOFvHG/YczftNx9/MEP6u6eK+rYWD0W41oGQmIo40+yFXOxhD5Rnaq8XFXC0DP0UJS7
qCm1M2BTIZd2FewCmcEQyluww0tow8BQVsQS+2f4inFlnl+nTNxsf1LUa9OJs9oGp/VZsCmK7CiA
uTCooL8fC88z4Utb+PxjrgwMhGJfpoqrx/Q9YPQf9pgprt49cannsXyfEvcAQv4W5x6m3O8R0fv9
pm6iESsS+nuqcdNIfDIFRtNHPvWz81UyUDjZbKNg9BdOEFtxOER+XVLTQNrhKejuLo1268JM4hpF
qzz5Ap7Oq6TVeyk3TkF4S2+ihbCfVW2L9Ouyq08MYG/dIgScgf4hOmc1beQuhHdr9pp0/283ipGh
IryyYdT81moTbYAUCqSGFl9XN0aR8XF8bKJ0j6fnQM00HUwDuNss5voZWHZoU72YtfM3/wpKJX8L
+xdSBZjeMSFcdRkc/TQ3EpWsPzkISWP9pJ/VCS6lMvyhnvq+Po8khVIQil2Y1/CKGjxBuA+8KTHi
+qoBoItHdmPw8p4ND8lhvk1BUTL7YkDb6vv3y+H7HijnjeMpfzcfvRwVK4eZzrC+oOLtSIubS9qC
hpOPg9wBQMdwHKaYugRdqT9d68cn69jSW1h4q+rjLIJp/m4TgWstxiuAA/yG6cURpkk60u5E6Wpq
T3+6vwraPM+4hi3VA3FMseMum6LwU/VpMRazD/lgO/JHh7AlRMbTWUt/xNA21l4e5TfxRdBA2uzL
sSeb54AuY4BrGDh+nsSCRJGTusX1s5/5UeIAjqufdr8gsUt5NdWQ5V2mMhMhB2iRDqzki4iwOz+6
HFjaMUMsZRcUaslglnO50iLlR9GACtVFAg8QtCcsX/15A2Fit1LUHkrdHcLAI2/42HdwytpAeBYg
cyO22V1eY32YMn2+sxgDGEa34/HliUUAQHDgj1G+1UOsr41wuhRy9c3yPtyDF7/OPM2AMdMN9BI4
e8NCjLLwUxJx4lPgeJkgPtXuMg/CxpeguLKAH7fJycV9EZ6GSVdQe5O2IpsqtzPSFpX1ojbvOCYr
Bx0Iz3jtTp7NmD+XwJx57j+7u0ZaBiJOw7X2sZcZgO8FNl5DVe1NtC/qr5FbbBTWcWBti6ZqJ48E
GrCngppkHjZqYHMPsXkfQluKPvX7WHskEgkvGeC8CGh/VG5/u3N3s8q0N5d6GD+/q44oKNgomOxQ
My7/M1TFQ1Suhj1znstrxjMBmXpY3pMCBXbWsZqA3e/95U5Vzle5+aiyXmdMU/gDcT/1PMHVsV3E
rt4bdnX1+zbpBM33cs/tVYP8iGHqzm3hMKRZ7P+d9wafJFXeyRDl6I0I2QMNCSX7K/RYFrxpFcem
rzjBEt+FkGRrHDsydwY5oDdyGp4akU/g87oPk04iVfhchiGeOCa4tODuw0dBeRRrkC1qkq85ZQal
1/GN2hLXl5S4fe5Grq4OiMf1MZmSZEimzwhKlfV1wr2pmP11g3i/hNt2h3JYE5U1dzxVxhYwAzCs
de8SKPRXMgCD/DrcZVPQjHgGWz+3FR2Yrn2ach2I4oRa/09ZeFmJ6Fux4u7S677VcRNPLZwqysvl
4MWeJvwxn5E5qWvs00qG/4bZfjJDP1rmIKmMNoXT3gpIMlaZJiJ+qY/dYTxlJqghD0htCajZym1K
aAjfVz8t9u9yLT1FWHAGY/KSwefdbbN9ITCttR9e+MoOgg+WRTG5puDcR3QCGSb7BG1B0sa2ELPS
ZhK2voS/B7KImxjun9mfOxkzm8nN4LLWiP6QeTgQcX3YFZ0DSWv5isgvY+Nkzfoq2gWeIGRjKqZS
q4CoPQReD2lqHTDlOYJAEz604bL3g5xPK68IzyGGNf1E3F6PbUi5bBCN6gMafYxBK+OufhUjixaC
2bmr/O8uy9i8lwvEEVkAXOmqbs1YHcC8NzrnXUBn0uMEVRfROcr/2w+6U6V7KIbuJP6QGwMoLytG
SU3DnCX07UO0d2f99aPUDRN4cBEyVJ5XHeoUVAiASYwtZlNGtsJZn0+3ITXfC2BrLwqq/ozXj6UF
mEPmzzaIvoyCbiNMx5ELLx++2avNHamPuEiYJ1nelzKqQi6rvHqlYRuQsh3BR+jTxDaE07n4dXjD
5KmOKsMGDvMi8f3CQoWVR8D69U+VgtpELCEFXbhCc7yRn9StXj1MAifNCFcDYdDHFX67H8S9rufm
fBlnNz4kbK7iEeQD2UKHemexD2dI2jtemVD5jaM51p3h1LPPH+xFrXa0C9JSyvBdeigbmQoeYuvC
dWcPSyeKnBE5d9F2RzErKm/r8/rqYU2b0zM6Xqp+UteLlpPQ51FRz/q6ALF8GRMf3I32QVp6ZxjA
I+Cw3LDKOXbKo7a1B29YZYDNL4nr/PL1ftfz5kH9LQCTMhpzkra1TTrzV4FuIxDMx8O6DZ/8/ecW
yFkRmS9bQ8Xm54LYB9Dw7QCatAGZO4bNg0YIgp2c8dX4vRIVrU1isW5no3eZDhabnw8dQV1gs2mv
eijYvpKTNm8OIqEl5t6/uYbdfMn2NHq7vv4Tt8T/y3wEU2f3E3iduiOmofioEAXJGcAEWLzc64iQ
WYmdJqD6n0IKbQ3QDKuD74Nst1ftdB1iwkInIUZiPNa0efurp0u5LcQpfWeeWDCdTRBcJM6Yu64Q
dhVYylUrsy+W0HDYQatxS862JeAdxx7fm2wDNzqmsBMng6ayQOzj6RZCdNtUSv+tawYy4nItvxqM
q7VCduHgyjjyqJtDbEWi5fco4xS4sc3DcUupBwFWpmxvGOzbilwSpYDBvp/4NPHEyMdS02JeG6B5
FzSKg9buP6aNY7Vgte1vKw3VNU4ZJ+d0baiQgF4Tsi+hygMd8A7Cb5z6qchVJQdPQ0LggWIy9WU6
9ID0n64ZtAp+ihrLgOvHyM9YOXkvIthjRskUQb5641v4Bsai0twf/ffaG4Akh8qUioA9OuVqYgy+
DTvTwMmDGGm+UniFS38GykRehJCI3szhI4e2EgopR4IDTafls4LcB9JG2Mz4JzPXbnhqRn3JadwE
58Qq6MMI8JrmBJInSzVndvfrvfelrdJ62JqQT/2jiXThGnkofVIomqf7y497vMwqoIJ7M4Zw56w9
pHjMKSqwv0EJcCfHHeqcXk5OX/OVnOKptmbb/3aQ8QsVIiyWN3bZEkdXGaL/lnO9LmibA+bMCk8C
0cCvochdR3NgGdAVLcxk6M3UToYQEazS0pF5qvdDhYoKOCkes7K00PF0v8T/BaY7LA4FBLOWeX+I
Gv8ySR09d4CRKhm6DXdD8SCPlTgZV2xksZsMgv38gZ1zr8+eWEZxRlfn6gUkmXJD/9o4ecHGSBNx
VA1FOEDP/uavxndhtJp6Bg+bO/JLvHAvaxRmyk4bxL0zqbsO7MuSCRF8yIX68ubH8Fi4N/WYo8VC
3EdQgIYcDVaR0lfetj91EgP/Z57FEgEKY8TrD6kbf+pBGVOnAZ8y8+E6fLxiKwx1Otyu9Py5ICq7
DBWTX7tcA9zfutD3AxNF+a6lxLbEsZkyJqmdUH1PZC3bbBNXy/fhLmW6CTW6KQb2rTnyNm+qvzoN
65y3OS6Nqr5BEnIQ5HLBmwGj8Doh+eKIGLAfJ0mO5WXSeMUlvc0kDIiv6cuWnHkAA5kA6wurgBZ6
ZJ7+TE2rGTu9vznsgjRvUd6kcZkXS3yUrPgCEe3olJx5RUYn8YjJzO6+RMTC+V0b1L9fSLASSo4t
iPl+jbNpWetHu5AjeUPG9u2/hHabdY4Wfpt/kwcBgR7p0Npwg65KNWLFuLLMht6fr1/25+1VnBLW
uf+hTpnMRm2Q2i3YnH5hJF7OJw+xN9gL7VskDhc0RAHGguKo1PHIJzaXRkOCnokrRMr7F76Dx7Rk
aBKEqyhip2kFg8QGvbri+XAy9tgojRVJBld/vg1N5U64noc+VK5ucY+klj0SvHOqLu2/zHx+H1GU
7GmPWO+zVDvGhBl69kkANhrMKIDvcrM0Y7pGtqLWv1Oq82dYLR3R3i4Qp75Y1IVodr9pZPS/lE5l
3EkDQwSSJDAsA8rCl8G4yujNWquVOT9/7R+q4yv+zqmQjhoJ6ekYvFiwvBFRY4OZP68jOT7vToq/
wuoMrwgOgZxgjUW69PdZs2qv62+1g+9o/wWTn6T3xthX4vJSYMEhvu8eYX3z8tI4/kcZZrBmu0Ql
Jn2GRDYY8jyFB7CneC8ZoJuLDUZqDwmIxqK3GqNsGXRhxBvDLjbLQCOZHZUhzyAvEzUInLVR8ImR
i5q/qsPvdrtSyi6z+RMUxcK6K9w4CmI5BWntI97mPJ0acbtlxKYX3kOiOGINt+itpNc280sAtG7o
W4ImE4JHNxzIF9PqF1ezVc6htrcJxAKc/JR3x/lsdjlDjL+KTR7ewdg1FmOFloM0fyINEaP/Fy4C
a0A9dOumyGaVdO7oU5fmtATFeo+g43AyY2ipHmnATxBLaEM8G7Tj7W/nB8PZs5LYwgsqULrRxz1A
EOqpg+3i4X/LjZanLkXuaCU25UeCHhG7jSlYWulJeiV3esTh4lj3f4hom2h5vQBghLhdIdQEx0CM
WS5mHFXNwfuwf15CazRDv9rSJhlvRbha0VinVfjC2+MLssTUHBYjGbfrKRJN9tTUwMwnXx6Hj93B
oOHfQtAiNxQauelv9Dvy7l1WOc6LJJRnRpQdCTUXlntzrvFcP4aKzi0wj2V6vabGma1fCejEOWFf
/mftWZ4ElwKrGpZ9e0r+cyxZoNfrxXB3QY+sqPUQP1ZzeBSDk4xVhZVN3wXO/Zm/Pdof+hG4xWNH
/fDxIuAlLpT2mEqOKOdgh5Re5cYNADEiTYIcH59hs3vqRC6yFcC4+WGIDJOT+gZ9R6KJXcdeSv2C
VVt72ML0Tc2fmBQIMKkZUFzsPu2uCs0bhO7+B0SGixCGb+bAA0yni+KCxflyEkkaaEKrArQfkUDX
2oOSiy3CGsd/YNB642Gc357dXU8feUlIkSA3imoa+M5BHEPyh+M2EiBCHyJxcs8fYIKahHsWIFcu
U80MkDzteT+1VhdGxlf9WbPwYtBA1HU34QEZLv7MRmogY8X/Zlf3BDZg/dVvWc7ndqZtxNLBoPVg
/SF3Beg7XX2FAqbEH97z8WkdkdU+gJnixXoXfwI3MgMQTBhQaaXOWOva2KV+2h+B5qBX2cids3aZ
nRbo37yN61PGcosyfEO+YqEFpxBamhXUtYQNpm6fyQtQP2zaj6MoLc+/afQQOg5bOK/opZO7igSH
A3XXdLteA7KNZjVaR52UpEE/PxwLW+pyi2ObZe+/6aSOVjTiFRlxjEAmQNhxyQXr7u93fQ8A2rvS
S7x5CyvFBSvtb4SIlb/o11fRxoeq89DnZCopTY5KXyOV9Zyn0LH7eoluOwJETMufVTrTAmf0gRgc
crFfGHa5Uw2YbNeuva0RpSYUZG8YIZyqFso8jbprTuMQbr1S6u2CAXOTZb6bxCoWlBUq9w/ZPV1v
aL67b/dtkc/tZfOhZb/gBZnt9mkgbraAE5aP02PjuInBoI9okTIvDwmps61R78HuiX1PgtFfTnre
F8aKky3AyhsvWadqtMxyL0K9tYIZ3aDb0+q71o7BsOMuSvlZZt32NJOaf4oRNex/qR19ygVQmEcQ
ML9hP/edS6v4+x1STc4dcg3NBLr6EoMtSQnAL7Khrf++4wclWr7fx4CMhlld61fPkPvwY8QaR3u2
FjoJDqcXrmfia2NPRwEDURJfP6HnEpuA1QkxI/7aoS/VmdV5rIPfiDGvzikkNMuVS3YBWnyfrp/h
9Y9V9Qsw/uZnyFRWp9rqgScm0sw/bCn4KlY2YMM2iy26ZXeTH9A98aCJ6o2I/T+zjtEXWi6tKq/N
l6QGYVKVSEIVuR0l5cIjxEQywKAQEJ7uf6uVvSVlu8tRBgqtms3A46FDlQI1+gA4Fd4IbPoLFrhV
EWKbVZnj6LEcltzp7sbYURPtaF8xw2gjCC+P/YhLQvMYSbp4xsBDu1oLYCdNzwjuK5J6RDB4yEX/
o/q2rkjLkqY73BINX2ZLjJzNRLTuS6FkMKcz3+MQG8dik19guqvoQjfZd8cGm5rdz/SsGY9lVA6o
/dEBNVjGA7EWBuxUVQ/E7wmgt3la6dMpwVnpI/4V9x2flbPqEOjQoKS2Dnz3LAoiXz/99I4k60M4
Fea6D8sNBMwELvHxI8iNz1gZpeY3VUMmHjILMd5GUQq6Ea49uy6mecB5U3U4e/mXIb906LD7NG2I
gNITaLAgPL+5H/zz8EjhaNPpO4odQNLSCYelmQiGYVHdwp/KTf23NxOGgq+xdJ5wDWEf1ECSeTGG
b4BRAlxcLHOkjnhmjFAikPWXqW3kWbz+Iyl5T/ZejGsyimN09ScnDvL2geetduGv8IskMkI4A6Ea
6aA6kOdJbpjPvkOqwg/wHPF+AB+oV3liSZjbPPyhD0/IKm+KaN9jdUTrXQQ7wY1o5MOB+UwiDOQ6
euXMvxEFL3eMy0eZ+zjf9FaTZ8MEEexS3sUofrB4A5t5Ug4uFxVonPoT24z0KVj4AGq/0iXnxPk0
JvlxCwqxObq7GP903nAbC3/FR1Xz9dBC7Huxoi6qBtTJVZ+SDYmt3MoCeQHPyBEHawROtglUvqUI
04ecY7rE6GSRuAoP3WNcW2BsjQtac6gVUElEAMzHj7hJsotTk4+0qOLIrizUeeQEiiS7p5vQ8kpC
vqA70zAPctcxEUs8oqNfwh6KdmMkPdRDD1hFeYwzXWYDrmcvER9JwiGzLKjG4NIrEl2IPybXRMGu
N75FyLgEVtI8mQo47O/5s89XrBDAO5zlMtGVDaU5XCl2m35/9o7GyBYOa/zOblmfCT5a6SEQ95y1
dJSePA8lF6pIDESTYWg2qI6+W7PSXVjeo4uoK+GTbe4SopTESb796g6K6ZtzpkqXHGHGki/bOJB4
kGxGE/tIqMioBwtbvNpfpB0pwYWSdrzJP7gkdRcey/PPRlH97mjI4z43kbuBMrK1NXWvNCI5WUny
PbbxuzGl8r19OhjXlZ4F/tV7igJEpWnaqMk5WlCONjWJG9fd9m8xG2sIVGCN5VNi9mvANiyqC0NY
kWpklb4b8btghYhSZyV+Ec2kkDH1+xwE+wG2MVHZrXvrP/OngmCh9zRx/KwSBa6KkjUC95+c6/Mk
3P0wjfdWC5jr/M/PFAqvdukVVG/ZLHxt4OLEWAddAEd1b1rckmSk++4bwiZWVUncEHq4RLM3NUSr
GkUyCdnMkWpOwIUEfDadO8c8IP9qc+J97YfWa3SSFFfK9JsfhK3gD0L/hZ135AN4kn9qLkdCgmlH
hE4cAVlNmIe7aked+HT/Oai3bGi1iWcmKcrzI1r9zwYQs36qB+DAXiCQxPAU/1dufNirN0qc/stO
yXkYcnrpMviQddqCc321BB3uZo+Y2QgULMVX04V6WOE9JyPJkVVzzeCl/GOTE7/nknIMPqjYqs6P
ObvBxo1INJ/a5JaM05lR0ZRbAfTgmmErHXz5SkpEK8rJ5Tyf8jvphH6XB+DNo7N6FWVjHlpaJEYU
Dtueu2o4l+L7ajGnEOdcL+vVYAe0XjBnMrLcNX6ug5WNn0ToYlRFJPVI30MVb0n+j465CuSDzKdR
5DwOGSt4/jLZ5QVihnVmfYcyub9sZK8wf/Kw/9cQoeoHZwQHX8a0eE1P1r3heLlRvDwiX/r61J/M
f+R5KbMQH+YQUrD/JgyOk1aBdgyDq7ki2rvKyOd7aq5ta7U3lcxinzEOs7b12gRqTpmD1EUNkvf9
8Q5RqRByF8NswfezVYDJ2T7Id/5f++t3eOPL8g2kbLCNqP91ksvUs/fAGNAoFfjkO3JKo9ZsDBep
1D/SU0MSVq0REcndgAGW3xfesJg5GjIFSZ6rUubrY1IXzaYgclCJkyg4JQ3B/BmiNpu4IMuolIMR
g7rEUVZdMU/poLp9Do7kkHih35DGbzxlCu7H+A6Ws6M8KYhqzGW0xI8KqLLsQxnz5C4345NH/Cfg
b30ktoFe5ksMTq5na/iPPm0hEth54s2aFU1K/fNhfps62o42Sllqrka0GajdoNV0vVKPMSJPNDDh
pZMRBoCSRX9rHodoVjZUWWjQ18biqiWUdIwN6zfPjPacTqIurTtAr3RZBdH6wTKlEwVppbwJ32Ev
Qa95Kize1JUYTAmOdrhW1SCmPMc01R/TWzouVjdnGJqrGEb4D+B8rBGMLia2nOfX7hRTGzwY8X1g
wMDOgnfuO6+vkVZvm6/JJldEvu4yMNVQm88fJdoETFTKVREKQwdzh7o713p04DNRUWsjXp256hlN
LKW4N7nP7p3kyonyJfn9IoLGaqcRVu7+TcXYkAebohJaj/ZGNjTbdNsy1RCFphu35L3jJmATfi5K
aNueBPc1DytI/B/xVThd/63rzq2UeQcguv3XyjTFvC2Uv2RKx2n1ts9Y9xpj2xfEMVSyOCaexev7
vBI1Vu+UFCdBofLiNCpxcrRwme6B0QVqHA4hHoXm99LFljWetmEGSysAg1TRPhbE4mEUHKIbK8pI
U3xs1eKoVMlIj7eyQZLGzRNMeecKsPKWssYeGupsLxSruZ60dBf0vzdKmL2qr0anQySus7oP7QTY
MuE9aMowqOMxZ1aQkXSeHvPcw0jArBYRtLlpFEApi97BVwd25JMT5tzOdSGOAWIGD+djOhvt6iQv
I/o82lheD4fpqccPq3j2mfiU/9mMsf5oZy/m9ZSIMUWRHZtnMydHr9EeSiVqMMAgzGtJDhbMjEgj
jxi2fuuF06oMohBsj9KLzb1AONBvev/GrTiyEqFW7W2gVXJ1UyNRskoMlOUbngRosrzi/oZQBE2k
yDQJssrp42p1evGRA0iu7rsQRZ4s5td5wwYbfhW9wydHj2BviCOK+Y4Bx1aGrrmekn786/Hd6TqS
XZIFCrvp/T5HpEX3QFyWpcA4oFmVWxKzce5tAr0mJUbdYHjMOZqW8sMD3+o/OIbTlhQT9TIFJAO4
cgT9HHpX1oz/PWW67nLyW7MX8Fbz/yjzGPHrApkpn96KgG0H0xVcjtkxPnC39OlfGLKd+qybN7U0
8/IuSK8c4nKEHyWzh+Eqvzn6iyFK0t4XZir3yVGiN8lsvpnIqWLQw7zOfPMJ8Cf2c2RyLT87cp5p
nCbtq/U+6sLBckbTS6dtvT6HRcKDLpk4353fyG87iROd8sTpUsOg3p/phLRGfsMYg9KBxtTlEWY2
Fr1VzCPrSqRCXI26NZjSHEgLYlhDWxu77WAwmI5TJ1qMz51jGrdGePDYQeIKpRXv0jBMqui53T0O
JkLr4cQhrqb3NcW+O+EzNn3tbV05wlbKwdhX8feLS4AbYMQtJRaQc9tucotDUBsFdPXd+Ql3xPWv
+YLn2cETX4JaVFHUUEUZQTmb+Acpybm8ePHk8m2ALaTXvgD1lXBhExb6vC4mGJKgBMFO2KYUdrRy
9m8oUaC/hQd/B7ojTu3gj0o33Upjyrm3WWvPddAaSdmE1ce1cp7IEYVkO5+1hgH37uk0b04PFNMy
bcuwG5n/sEbcXyRG3GLd8PHIT/MfdkqF/csFrupw4o73hWsbb028tHof1IiuyyzrrU+5G8JA4imC
kvlB3/qz+DMl1IGeKRLXNAcKym7SBKWn+wSVsSuLC1GmLvAN79UaWvFg9xJVZLz39OXkSIUtSqum
RNEor62lMT3qmOX0nN+8ZQGlz/mFpTp+lTBVrqY+N7CKy08+86o7lfIZ1upkRbEeV2yL/T4yZnvY
/0cCx46GydJbRgloMyTwvlqdBXNnXabiBYWONa1mbwrtGD7lpMq9R83WthiYuTgLxl60qdhNxNwn
aENI2F8G0fFYLyajwPU6m2J2Z3RK2eWIpc/kis5DFcOhXcnv6ufBaNSseHAKwjZbQdDkyXZvflSP
I7qIH5yKBzmvtPfmsnrRcznGsLG2iDepZfk6TkKPCccN9BS9uAyEixKZl1MFi17hoyL3dM7GCBJl
2Pfujx+MaQJIjUkIRlqf3pfrL1ndAX7mhs/O9vhPBrVPwFqvtiAtJsqlwnse/AXdMrUT0SKSpX7h
qatASYik8N6DWy3ovk8XlotWtF4EIj9ijAqv+1dyNejmdHOvnhWkx7IHnLtK40JU74DaaeDzeNBY
aMDFTgetUOJw4A4jYAHgzwvMVQ2bdxjD5RgPehidi8pCY26ilbRPBOE0dLGaXKGybxdKvRtsFddR
Xp+7U10GzgUdn6mM8y/A9jR8k/hbYh9w8fDpsMpcNas8BlD6XDfHaI6giDKAun71mWd1Ono946BT
59Gl7jinHcjvVyCASiYRzW8ObryAYfvhHYx/KM7lJkCfB5c0zCWPYiZgblpzM6Z1IqKBrhGzEX2J
IwdQGsPUG2joMU6MqjNaesFqqynjY58900GW3ORGXjCrXxRivCWrrQNkeO64KC5q2ImapqGmge0/
3kLPJVmS+wWUL0pfUrNCMdvOJqoV+XYx3iDKpdjUik9YQfkGkC+8nLX5Zp3NL2NEJqonWxWaHDZF
kWPbn4ah5j12rhADlfwKHB/VK4ZfQQbvHzG0EMMcTylMtnTjdEbtUATH2LNG4QtS5II190czSPyg
dSq6Pl3Ca2y2tocOtYpYWHG/jJP57917JQlhu78uQzHNgyHAU8Cr52qi2DL94C1J9V/t321RwHm7
LeN4Ol6dQjjmmmSDqgbBXmDFVAiTLskO3hgb9Wu2uEkBa6D4QiyeS+aMY7IU7J/JSCKx/gm9l7So
GyW4wDtm8G0c+FSbU6QdhtU6ZvR6ddAdIPbLyT6p6I2Q6xCl94BR+iytC5oSdhbuXthyqfrI14Hn
79uYPXWbrKsr2+pvYQULqE6HrF0bfLRyhRSNwmp93tsLSVYxQMVUpy5TM0X/P+akP7LQGMr58bjs
NMl71aKqmctO3TqH8C0XJwAMSX9mqPES9b1GeRzHa/v1/nJOZs3ZG/eG5OZRghK50PZoXlqJSaAC
VsjCjxNFKz2fGh1VOsoy2tSFKdiN0m+FxUMaK3n8g7xuS8tQ3KIo0tR7rg0tzhTAnrys0kWIJD+h
BhsXTlsfhbgqG9c5dCOwK02ud4hI++G49NNxAFUaAAm6z9E7SGus3N3pXHNIANWlScXKlL1/VOD/
C1C3PWJn6NrX+nvuNWrGDkzARk25wyn7B55R/RyuDaf581wd0BiJcoVFcQj5HvUXq4/hdheEAAi5
dYHkxuMe1OihyK+DcLg3+P4I3bHfiKpTYRdZQqTBG5NJfUjX+ztEL2AACxQVxMRrHChLNYRxQHMW
Nb6SMp2kg3/+raQV98J1PUbjYR9mY32mznvOG2HxiRtBb0SzbdhPdGzfRFqupqiPNd594bX0vb9K
kB0ozBfcgUETyQsliY+xWbj/E+xUceiOuEIafgjnQ8G3nBoH5pgcCmZ7mO2XIu0Q8LIQVBw70/mz
dYC1BErQldIxOxzVdkgJ5nI7VZS6ftuxxFUnqDoN4fgSQgICvj2meXZwtw1sdrtFFe6A2Y26OJYA
XKSEHVjGii6ieEPRm1K/0nNEPgXwP1rshaNuYygFopv5BAyiv3H6iIXsm4v24k5YATxt8tLqikX3
M8Q90Ynbd5kSBI8lslpzIhtap43cVxS/bTqZJlMKwK6dXsUNjzjO6qyHywc1OtZKcDWqImUdqt/M
yECXiF3hkuRVfALxPpHyqqp72xMXUhy4tQVU8MEzTmrze5Fb6e4JSCag+EPxjE89/i+Zd2Gg1Cdw
81tEMXyZOkO8LWkbgP3QobnD5L/suN5lNk3bs1xwb5RMmumdGAHEUKo9KcM+X4DIdS5z1LV756pL
kxDJTOZigOrqBb61BhwBJCVt32m1g2FcVBAIUTW0Mm09Jl9AGNaeyL+Z7vsqc7Z9NVjKC4tFswFk
+/NG9K2CiL53GIx5rKf7Jt9gvwfRUgmheCWGu5/EuCra6w6oafOgQ3xLzg2NgtuyX6O3hkPqfpBL
l5KcG32zFkz1sWwxEY71ZGD6kLSOSKcASS1ekuKn1mRaLX4OJ8Nzn5muIAp2EdBLC2cA3ago3bNl
DyHXvOLFSk1EJoZPKVRMjMUOaH517QFBb8fUviUVskzNJp2PGgM/cUaNT5DUjbM5jKoq2oruvUKK
pgY8jlivTt1P795RQRn96DnZrIyKPReKvermxdnGThmmHdRaigYhP9yOyMvevZ7/GlWKessyYN3n
Hqnk1U/bn6y5QSyKux5JUC3q8wGsjkuPSlbclWGQRKQMjPb/NBdhiV837bwOwmscP9PzSX3WJEMJ
OhRqBt/vPDFYSR9AegO1RDjK+UP5SG1oOwvXk40D8Xz2oeSvHnHcjqiERuQg9xKA9F3vkKt+eI6t
TGdukUu9bTTWiyIUbAwdVSC9iWMLwJ4vYMu+QtAYiocAgGS89GZdBwB4+/AbIxpzx+QdmQilLHhy
Br8CFrScxVjz12Ynlw8jpm0OpZRyXSnexLO4s80Di1v6xK4uF4Rx96utxZkDVcmdrt+RkSUYDTol
qGAL37C/oSbmOPOl8IY3vF+GZwKyWNmjPLyMjO5mvdLe5qD1iPdfIg7ytcH9VEorBib5dKH95igB
H4vtUe3W6fWHd135jssaAkkbGXpXIbgfJaTGOUunWeBhHdRcdnrLqFa+zvcpceI9wEB+pACb7pq5
93f3+gemiSpsuufHM0jD+k1O2wwRqo9n3oaMgnKePPKCTpAc2J7EqINvInupMWHDxu/unrtvsiVg
P/vC2QOKbOtsdexYKUXXjWLOPMwptBT3ylrx+97TMDADH4kKNrunu2/QGiBQh3DT53I48SXY1QX1
l8RoSp0getCffAssEKUQQAHTQWplK+KDzR4WVrc6DV8NbKltygQOT9gr6NgDNK4Kjb1gugtk1FfM
iCym7SewQTQvGwI2ThDCeKR+LiZ94WkBa/kQl5to4tZFA8YeCOvqtXL7pHlsTXZtO4zelBhLPH5j
V9Wz8ehTrAydRmxPDtT4/DNm2Fo699XxdSiLLsGxwZsT1RayEgzRKrNzOuL1I1dA5nOKCljhzkNT
IwidQL5vwq67bdtWSBV0aqPRYZ3hlwcD0SHQa30WrvgF0YHuDSHLFGY9/krq9gK4Zz4X0dx8aB/Q
pmi2A32CeeBllGHsKD4sILxtZGU5JY8/f0ltLeGwWHxdXmvcT7kyuSbfhSBFssTLeU94Q38ZkFXl
0o4Q9CmbNOsveF+cNAEe165DcFtVCscU9PCOpAkFzJDBOiudkpANkNwPaHQamLXUuWOLhsWOvcx1
zxuctWGYURw3vChV+8nAT5Ma43vo0anftWBwqCelb+FLVUCyqKy+FbuGlT5WieIjmU6cnkx71uy1
GKqagXon4KsBlJHWsPVdTsB5bVboWd3VFoDGRbsxBJj6jjELBfoVEsVi3IajsAIXma9f2vNZZxIQ
o6YB7aguBXYwNYqY3uPfet+PBv0/popbpSViY/wMzDj8lDfEbRo53uG4Fmxe5dj5qzYviyat8Agl
/rCxZa/j9iC7cy8xNkvjchdmlDXyRp/rSQUqXfs2OxwrUqNB2r7YxnTGaWpHjZwn9xps0gOs6jdE
fthl1UKvKSj5/G7BFRRwDN0NkWE44ZrcW2BhKorWxCfMOSk3N237aWFd2hJ3eV0c3zcNKlq138oL
ITCpA6OtAjDVMxaa/W20lmO/5Ba1SMMba+SsYdKdtrg+cm1p79Nr4OAEsV1+kqYmRk68KinLaKW9
gKqDiCdrV0qLAkh31sgz+jUXlj7PP/+7PeRzPZPMjjwxyYkY+XNSsLIUfAQsCh9BNrfwAx47kf7C
Y6/LFHaVXMSnN5PVhoDZXwec2ER3XQwAl1OnM2GicHwi5wp9dTHwOB4aXVtHTinL16vmchm/rDcA
gdJytkUCOino/tVTUJnsUwjL88C8o8jRnMU9VMB7GHr5RMPK107ADMgduUeKjhvwNTwXGW6jHMJT
rqNK8Kbrm/LD0e2IUX8amFzMP1S8QtVjwnmXgqUUn8FfwExp2Jv1g+o6CqM1FNP36+TTlnhiRoRe
WutR11u3iSTlKM9XMvpKY24NdxlZsFOpZ0LJTEYgXXhnm7Uww9EBPMajL0i0gLg5bioY9Ht4dz2n
LWEaQTde1VGdi9bWrJ59l7WZtbeKZsdUun0+n2peHEZDXuc2Bxa4EtSrQ6cOODUNQ/H23aB7JIoA
rBGX2Ksxj1tEYMSNzv5Ep90zPp5fFmVMjge1AuPQclq1BYK292xWVUiu+QbwNqSXRQ21czKvJyvb
iKq0m0+FlKPyE46H2MMwW218kYbRUhC/k85kc3IFgCjfDoQj83HcOJ+xvB8uQh3HjqNSKAJJCZiH
f1l0oapPPRylXVEFQUrMgB/9YwsNbWepGORx9uJapy1RFhy66Xt82oaaFI06UA36mn/RENpETWZQ
JP6ojt93n2DKUqiQcSc/G9FkoJue0mCGtaaGrmDXFlG3TlC64roO2iSRVENOHs4r0K0j+RgAbXi/
SJGVd+hvLgfeUwFM+cJrgNluaDVy4Rzy7/J5WY4Tyq7hOAsgASodNnt3P7sObsd+jl64cdDFoNuX
O3Vt5KMo2D5jnNGg9k0SC82qnxxGEhcsziJ9TrydGbc9eVvZmm51MHzHRfJ0zlBKSJepIsFdLa8H
3kDTgrPxAOGPoNWVxZZQ74diemHEtD9cJuIWWOq10zNZtzIE7BRNbTgj57jXxMuOyCTJkjZi6Li/
F5RduKy4bFvSg+YzCfYpXvbfU6TrF8UFETwu1bsvQjW5w55tEXlY48r+nTVseGHyponzEY0GjuLm
2d6sN2VVT0YVJDuuYO2sgm3QrrvAQKGIN5unOIK6kZUjqzjeDRbWFmA5q55S3SUCFKzT3anUTqWs
m4G5Mmf7CW7RpyQtmXYUXnMXGYgEj6YozVzGKxgtvXaZdpSJUpg1Bt0wmnhYPsmDwiNeLSlngVr6
el/8hQeQ1Dv2T1+5q0isGTWHkeM7gaGibl19f/emG8gelyBnCcyH3gYWO4xQANDn6/jleAPqOlbp
uUH5z4xKnbIgUcR2sG7cjH52pMTlyPbxMAcQfkLQ/jM1/l/3av46pbtyH5royAu/cBNZIZPupHvO
oXiCVizq9JTV//aht5QwDItinMqNRDwMPJb6Ap4nO15fisG0toZ1bzoGPhZsdvowilrpHPJz4mpG
lh0McZnDXlmA9mNImvCiZ9b37YNyxZc6zbuJxPB7v2muMZnj3Ky3bQwGt6W2jjivs41mY6B1qcQe
+v/cSNsPBJbsBiDd7tAqYYqTvRxfrBkmcrHZlYe91RcVtCS+jM8GE3BODUncJIkZP1aF+Eq1NVST
UmGip1JIMxcqI2MnadHXrGAJYR7e5Lga+j+jApQ5S8ewuq99AeKNjglDIdQ0hdn24w9+UFqT00vE
+/prOpyiTLIGNUOZY4ppztPh9SDCoL+j0PqGTQOtlr2dEnkOl8CcNQuCUoTVjCwTHuFWFGq5EWiP
5ViKXcMm0423479WfF4bhuYqgB/ic+eFyW6lPv+7NL+JJuuqjcIOWtKEaZ6T6qsgcsSO4SbK/8Ma
vIoOtcw5f9Rs97+IXdIA8jC+/StBZpWnBZomWfWCkH3gWwHT8MCT1n0OLN/7lWJ36QVQ6p3eqjdX
mfGRptmb0NhuNFOHWWBupc4KDEG/2lSM7OA7anutv3slgme+cgStiOMJZjExUYW91TJkm2QBVLnY
CW0HwzqOW5oVznC0gDNrx23Tvr1s4/Wp01rClv4ndEat58B1VXvjit2449/yNfm+HVTqCWETapq+
zgfEzkwtCh2F4WwZREAJaNL1Yf8SkmjO3VMyvNIjBmPIlQ12cZnUh2b2mPCPurSx/WWFJm3No4gc
B3svuZd//6yoMs/Wp11IlciADi1SGTxmon7neBxyLBxcSum/xUORP6c+ZO7lN+Pa51evrEm4NAnk
F0RcNB9a/uYCh+twywPPmaOG/ErsN64+vk2ox1GJf8xPUQEaM2yTGdDHcNkrKEhcBVXn9sK87MvH
Sl0YL0x/Yzlc4NO/iJnZoj1tQGlAU2KDQENJouQ68kTURlkRkZOIFi39CZ6IF9nO51XG/zGJevCI
UewhVRT9/T5dVIMi/WpJnJQ3OxsXh/C2M/AqPRLqIO9sqOvWen6R/wEqzKCRk5qmW+huBwIf0H5R
2beRg6UCp5MhCHHNNYQ5xt64xViV13oCB1nt1b99uHR6TncMwzjHD7981a1AfZOzyrzIdWhZzuip
+42tE1cuF5h/zipHojbT8SmjaZr3cQ/in7oFA1rBpA8lYA6uv9LC4mVbmWQy7ChL147gyJzRJtnd
WWBY5MBbjPOzok3mArgBhqm17ILUBYerK+LWi2Jw7SVVcDFJyTFyM06h/Lhk1bxaOaOWGSa8Ckl3
GH1Iq9/Ch+i3xZgQoF6NlY5yxGbXUbT77aWDZb+4ek9InWQClpwBk4kGQrJAuyRkajI+zH+Yu1je
HCTBhrxUVvajkHUaffG9ro/XPq9Wa7MxuVzNNQihyF5rzfXUV8+SdwPZLz8ySukXm5GEOJGKIKTh
1P02A0rY9pX2GCVQ5X/ggB+Ax0J77zJrZme1BqACyRRzmgcqcnSE4oYPU/N6nt9MuaFcJUjNidY1
qUMFcI4EgH68F3IlyyaWkV2EfAd/hdjnyyRU2CwpcyO083gK9vgxyyWkE1AvfbZUDH710sNtTrG3
dFdtF1uGPUQERE0uV97m7MZ+eQxlpQmE1hz9L+Y47i5XZFD8UjeIK+X/0bC8MzuicZX2Mk7JhbdG
7+h24MyTRIyrBeCFsGB8AZtPtuel7ZP1pm6y7XX95qdWPIYc76CJZ5YeafuHaUt28iaul6bmrqq2
2M6VkXsViEZtI1yevpesFBJTs3RuIbis6nnd+Fdd92KBXwJ3LGWgrDF7GcN5SoRIJfkorNTjD4S8
LPa0nsf7fusykTFUuOXmSqgo/ihO7EdgcTyxd9YB0H+yWB2/sC8zJ4yjdXoCDNxq8dpBP7x7VVhk
OUfRK5PjKiUky7QFjp30jqh/GhsOSdY9fi2O3op82g5m7mo4jZVYsEsfgQCpbQWz5LsTVvBAHPgq
pFQ8gSjLErje6q7rDx+4vBC28QbznVFuX4zN4NSwvPXfloRNEVagitNM0KTm7xKn77AoxPHBH17T
r9tlzTazEX90vRCWqkr6FwvEpI9Z12U/hit2KANzty7P++2rfEYaWZDuUS0h65CPz9nr1xh70XHI
qR0LglvD1kDWULhOfA8Xjq3jgDtEAStvqSN0VI5IbLnAGbw8Js1fK7ltQEVGo60pnA4TdlpZOCfW
eRyqT5mE6SdLV/KJBDN+iyTmHoYjiu1qFrFBkEOXaW0SP5G6zu/bkuQNR2DNSbHvhCevhhmn7KFu
pj0zGBdpSP0Pf9VeymbXcpT3QczJzkloOhIrGgQypbVhZ9JtOcBSetZyPxi9rbkAhRnoEIwuHJxo
x6lSliTK1qr9ZZp2uKdP+M9STWGcKIC2yEfrUlHYDX84rPAt7LhZ9s0ceYH7qOGIpaXBSZ5ORZlY
we04d1aBHSayuUw11j0JHH+l9JbQcGDvWbTDlyFkRwWdaI1YtjixZ/fEyZ2yvX0UfbKYP3cI1ufm
32USy6PXvmO+umdxkLcmciERpUb341oGuD1HnBF3Q7RGKunIG/6UClq5Uqix13cbNA/CWW0VRFLw
6pGV7bWq1LfLupqsyK/UElHjFRqL9TaIM2izD6MyC48R2Zy6wlTVqwuTdzbTdc4eeV5cgWvdHxkR
mUm8s65mZ2c8BGrB0J+Ps1fMb338wopbdZrGYGM4Bw+U6MDNSs/TArvw0aUK/bT3Bx8pJQOLo1Uq
9vqaA+V1/64+0ooTap8irBnJRCpgDLoeRstwXS+l2NcRlPol9EWmiD0ZgSQfLsHh0VQwLor7gKHw
5SJhlos3lYwZeTJFBM10AvmwPClN7RSApstdEIGPlMKwP9P7YpdfDhlQd5ykMdvIqP9YPAQkowQ6
lWdPy4bGvppH74zvQzuB5a2HJCi8nmgnxyy1mKbCedwDDqyc6xwiI3y5WiIn+rS/kooAPr8af3Q1
eulkiqz6N43hhVGPlIw+jeCnedCPl9zrRJJ5PqstSVjrXgLv1t4rLnlTNqXlbqMJQx4oM1l/bU/B
xDH+rMDdTk6oBuYXlYvL10Kd+uidk9ZLq4cx+lT3Y0s73Il3xTBnFTVaQZ4iCvxZ43+VtLPFkX1R
4FxfmANGYBsQPO044sCaxFSmcwdnT//3Jb4XidSNePOoaj3GOvcwOiLotHqMBdZjdhZAA+6HUKqq
6AvVDfuVORgIa3YgW1DC1yQqH1gdSvs67F+QfYrquAtoPMm7kHWHNrGEo0+mCVCsWKgeD2/i7yMd
080rVzz8mVdkSDQhHdsuBUSX9jlxWqexWsFEYDyBl1W5gqGNfXE11dugqkg+4mPUIkwT66A/tDWP
nwogkUE+A/owmG8/eCYoNKbXZhNM7qpXcUvpJMMpOzdjpwLM6c7WZVVIhgvrAZaW/UbSb4NPnkvQ
WvuFrIjZukzRY9m7DTWcsQhZmFj5jhCYX9HWp5ZmMR2TLKUxaSmmDc7isiAzvOojnt43gXBhhqf6
nMRy9aqQKYoq0srmBrx0hAZmvpeF4iI+xiuF4HuF04q+6Rl2vEICINEKJ48d1qRub1OGB04W/jpg
WIXmbFqk2qddg7JqoXvmyVSEKtceRThSxT05bCIHgvcsGQonZZ06tNwAj7JWUGsXLIj94/WX8jd7
TXipTqc/srjjbas7z/zBgSGK+ITUbv6N4boN9+MYQ9AK1BkG6J26/BQjZd1Icc5pwyn5RuqDyhOb
BgvioxtcvCUHUFoR9FmpinLyz+Cg9EX+o2wAv8TYm/vgbmBe1hz7h+UKda/NJf4X2ATkeNtRU4xu
/E2eoPG2aIawhr3er607gDOym8MpgSMJZ6fsyFmcPZ2Wvz6JvwwUjOEDe6t2iIA0K2fe9Zq8NY6D
AjLAKGrTODgyyw0pR9naJbQEPUbjGEk5NbighBWomoqilhACPnLkmAZM2jZxroy/N+TjJX1gdszj
1I/2E7JYWuQtX+4NRdn5RwtPyszDsWzRXj995ekegff/RX3vutE7bYVIsXi9f4zsRiQ0RuzM18sy
1tEgjIEb1HcwYxjF9kMrveQfOrlhanzcKs4AhLLXGwKqbmo/6nt4B7kg/Yr+VqbJf+ENEzScGnWs
/3VRjt5lNOmYRjY0t74ZjYrPXFY35KuVEsvdeI0xK8SHfgklnWhNEGvA/ZlSSPuPanMDB4lVTXjo
J0XDkNFtAMLvuaJoCnO4oE0h8jUfh14+CvBph2cqF8sQiQB7h+NQ50JKw9yjHsXJF+PsiaG7sXOl
0bzqhYq8pb7/qATIPEmcTjv+whcUr09081pVdNwKjDt55BmcZlATy/aP7/K1ZaFpeHu8BlkVt2SZ
1DRqq5cpR5eJdPC5o1JRbyNAnGXWE4Itb6JgWB9ndwVS30F1sNIRjNBl6NO3wm5FLCIfx1NgyuO0
SJuH1kQ+DZJYwx2hquzeFElxWIEkJCE3vCAexn4kuztjUWbr21eNynyD0FyvjzElMqiccz7VqqvR
IDb+Da1h72QtfGIB+Hbf4amxofqPeznfBwRU3Z8vAvtAKVSKLloSKd61hcU6XQ7qm3YLJDeYlxKK
Ljco11vW83zh/CaBCeLPjT6sNScRUyqW3rweN7zAkWTU6Rg8Ci/YEvHQZJitJsetHD5Jy91gL7kC
pmz54Elq1S9DsqZTAqF/CaQ9RSqIta5BuGDej+fWEbpOUhMmVly6teDLrcFCV+7CqMZDqoz8zj26
uFhpBnPG9nM7aWxkPHAG3ZbgrWhqftE/rvWwBtMOcmnCjTI7p1+7YVGLJnWAMu3yIyjGX17R7anG
OheZYB0SzaBwV9zDyfxoGFlglk6Ol7FxQVm9iOKfJ+3PnxNDzwtGr7MD6GBufCk8vXEBvwmVt5Ep
gzEY8gnhVoCzBJX8Ea+F986nMbwc3cqG4ruqN0lM99usnZEyiin9/O1cJC/nl3HWMJobjOHGwAUM
rx85XghMj3IbJQZRT1LxELDW3iJHWXRZHnPRSaqDyhqUiNjCUvMMuXcw6dV5vEaQSzOtq0HDa4nq
QNpzYLOhkpFhRD8yBvnEDjTWjv0tcKsXszcKANhsKHLdGv+s5bdndT5V6gxFarx/o6/QIp1MT+RK
xvOtwe0GgsA5qbrwJ4VJXxP+SKpH5DsrFhxj7R1rt6FQ1yyaYjbXyqUqXup/C0eOThqW0bYTHACW
MiLzoLPy608Kg5gs5dB/P5311WcFJ0TsTFeROrgOhEkHhI5uvIx4pgWu6mSgG2lOyy4Z4FTnivrb
uFVfswIf2uFbxLsUf078rPHaYyrbaun4dl/vfP02lx5PWM5MCcdKusTMNeCPZ0ZWnpuLAnT9hyUa
Ajs3ccR+y7TBlFD4TH3Py9bxECcyifV3WX8ve7E9JSkiaPHC45jAyuWneu2x2k+gk4GF/AkDU4ks
EglEtHck4jSsYiLAOfCXUqT8ISkCVk2rV+W2/eUjWmF8eTt9Sevf+oSMZ/4zv5fdES8npQqmKsTq
phl57rJuRNO+YgyaE2Ufk7xsFT8NQAEdLhoTw5ItQ59gcbSM9LuMx0g6shVsNw8Rjg2lWq4Di+70
XMBf7p6HXt6ShBiOIvfXoorpIcFlZb0TEifnMzJJ1QPMzMLN5QSGAbxGXycSMmRH94ygjnkBW3Ef
ZdzylM9ReUV2XR2LEVfIqebGOmGyZD0LsDd2zL+YhCorJRlNhvEwqcnpYHZmKfUyycj9ZQ7ZxPpd
xc24y9s35tEllH1xVFFePAROjpaOg4OyBVT37N69iplJ6LuFr43KHtRl69aQW07iVMEPqIBfzJNA
92/hE0O6mJllprO3JzTalpeuU8pjpPBBkDrhPqm8ax478VCMco2SOd3iZCY6EDp0bVWkIj7sjeIH
/JpcAePRdwNyyAajOUYH1qIpuHoBx58J9yu+6FGagAQZ07xFVCUJVPlthfz7H5pvNKTJPtoAn1Sd
oEe384hOizROiKklAY8l26EpJ0njhxzS4CYeJfMC0QRXA2/PUJUsFSOKnsDQdhKP225yLW3e7cLf
rEIPhe6YqILiwNMbVrPg6ZTzjxmAka93GpnQpWstS3KHUV7E9QVbPqc8sFtIo52p6yXidAV4W6X3
tQzdWDItIDZKIQRevJa63/L820PMHmD1tmQujfqigz6CbaJxZ3x6v+9xbGBduhpSH7GSokSYKLlF
smGsWTBDUAAsAuWqzFepp1ib8rey3VaI3+0OwH7woDxO5tUM8M4aRaNyFRUtYxg3J1GGFDxP/sPB
01p5FBLcLOYiT37Q8pBPpBXYfscKpskc6CiPqPOo1y3di8mhn39o24s78oPArHfLaDHLyBC20gA5
hWlaxgdb0dYwnkiUkENpCYeyvf1YbZjtEvFt6ccxwvxyD2D0OFqYaJsZvSuSgez9uCzengeAu0Fd
7okLz35ZDhmhq5GFrRB1LtRl9I/WqRhp7P5YTY/bUeOwDzK8WorH7CwXE4oFcHkbnE+uP6tqzCf9
H/CtqcqQcZb0KpBE1wh2XJVIkGv4FEF3egBZjyVjnK6CtLXwwwDRTaqnIaa/Cbzg5GVIGdG2EyxI
EhCYBb9ONH22fHKxenpT4O2OLtNNPfrEkF3DppBijDGe/vkKNmCEMCOHd24q3VpkqRRs7bvDiUX5
OOx7Dec68EVxkE7Csnk1bpbH/GvYG0PCcR7VUPzghUGvD5v9uTqUYI4q0QNWAoak277iQOfvxOT7
RGi84m1eWNVMIkDBTmBIYpZx7T74IcBd3JdmNM7CtXY7JvmGIQCYxPb1am+fuHnWo25pu6hsQyJ3
NAuF9chMhfZbbslJQdO0qzJ4S5599z1DrL0aER/KK/D6wEzxlhHhzCIb9o220vSwqX2fegxhPp+G
Y4hlQHwNIAeK3Cgvr3QbJ+gMkcGJw5DkW9K/1fkR+KDcCla690/ffi1cJpo8b8/SJmTCnQrprpai
mqyA4XbMk0KySkdvEwkbAKfqWQsNgzwXzhtoy0AoXEWZxNc/aNAtQoGo/XtLU5wOl7osbnd9eRp7
8pxJeYLSH91TJFi23h7jK3qOQhruOp7jjKuYLAPf639X9VLvKe4tTpmN42WJ+dvgubQYz2NRljKC
1VYd8ZgRWSgKa8ZEBZC1Vjgz6YdVcmwPof0ssRatmvNSMloD9FMHr/VgWy7+505l8A2wndR8RxTb
6vNJT01Uq2KhrBx3EaKeHFGyrJO3ZwwiRkqx7vOYh2RFAKygfnSyA0wP6cBDcn+R4DsbBKBup+WK
8dWhmS8WBS3b9ErnHdaYpc2GrPUY29O1QtXfQVIT0dxklHX9oald6BNehkpbURC3y0NPpbKVw55U
Nxj1UFBnNHkjzbCrSjeSPU88T/6ew62n/dE0IY1enLerjr24phnf6XARyYXA2kfZGYLPmFDdxt1d
ytZ4Xax2VyBvJvnRddL6dULUGIQ4OQjcV5whsbt0bItbfu+yik2VBvGOISrfqQ1VBCKQtTg4rfls
hPM74Xqwg03wuLn1K3xp7wfDa8TP5wjmUDXQ92e8wC0xsG8BQrXnqennSesV6qaFkEM/j2VIHAMU
cOkuv+cNFf5spqv89+mN3W+aRXFy0erqbmNNrqoj6umPtfbOiuGJWm0pr9ObvKMLyiqQAo6OPlWj
WBxwnuxw+yDrtJT5Yv3vuRWP5TlxUxRieaVGgMJDNTL7FCXVzzo4/6f0Vl0j15ZDYHJdFV2IdTTT
WtgvqvDtNjf1okS4fb08jTJMhLMwpFr4HHdYGdjr+kRlO1vRn7d4h84VMOzgIIc5of3n1cexgHlX
DnAmDVHmhrlmB27eet1jn2CyhpbDsmi3BHGV7npuYY3htEvsRYJGzfTz8Z2u3w4gnIQN5coDcVi1
amJK8Qs6W7cP0nlVi+KuScelHKTutoU/GNxDDB0rTy3eJPregKyidVQslv4SQyQ0D5///pScCYW9
lfOP5I4wxtol5EP7gdnLSmfwegHkv1sVjYsz4iK8N4mVU3ut8E/OJgkv1Wakqfsk8FZ6txa+5wf+
7Xbu4K2r4Zso61TGoUQZYdcOjePc0Wx4LX2oi/jH5KxxDnlzo17aa/ZUHavGykjYQLYLcDOjZzhO
BDm8Vg3V8MNMI8LzjUOYEFg6sS7gOjMlJYyD8+/oQhRflyFj05KWxPgSsR+AQTOjf1rnAV2G8FyG
87Y9B03qosYyiU6ysi75mMW1q4WhA66NPr30owKN83+u6JVuK3dZlY9zud/pafIYQxHFEDrcKvef
DKFyMvDQIf8Nkza0LGKYcL3r+OwwQzOwRAzTCQXSJ0+XdogkWPbtZIiTsH4b3FYkxWRdZw1AzMvh
LuL9cPUE5uNRp1Mf16/GcSlasHvHf2pShk5eEbg8Qr6d4GlvMAIja+/oiY3B7nxdYma///evbuoT
eaLakQ9rwy9uigQ5xgdQskXU/Tsic0CQfgUOTEmRiO18ijAOta4M3vFHlDG1+CTRnGr0rYtv6gS2
mUrG10+ZVX8oyjPUfIZU0lNVsW+2aCe6we/DY5WwbAeBKHUJxrv1z5RIihit/SuDZfliyKvRzETM
GirNAbWre0MreMXYIbc1DdRioXmwh15/rTnZ/LFmH5Sjd5v93K2JtqN4WJBlWb6JdTd72oLmKxpF
NImwlApx8GJJz31hGnHF6f830jIJvmIHOwH3LoboWeL/vJc0IgLeqlBEeLrcCmNcl848F/s1mDn0
q48K0X3CQJD1DetpysWPaGlv6FWX6HCdN6r1nJGEMWtWJuOOch86l4UYd/Sndy7df93q/i1SJ460
zxlLGip1Cw2VlUJpVbad/N10pWbFMmDFLdatY0EMzSas/EFY/eQze4lNK0URPZUmWtLlV3MKirBS
JikslcjjZlRCFmYdFOn7aquwu0uXa+aeb+aMzom522FlEN/kqp3khYnyUyK2a4Nc7aKCtWT0z7P9
NKJvebPvCYekNKQLvNSv7kGJUoAFpP72ZZAcPTmU16g9rZcPFPx+kUMf/i7sjud9/7TtNIFhiltO
mIToOLJxkNtKmA1gMePP+whzrXvEpq94anRYDfmT8+ZjrLepHar0G0uyUPmmQHPYJL2kje3u6af3
okqsL33PgByrdQoFQGGd14h6DmxbYTCLO97UFdBclQVNn3NVtJU/OygeYbvcp+WaYnTzqJuIq7Bu
SviYldVoDE/HbBeaYruD801FVyrfkF/QIrOhDHrtbCspZVfxRINt9c5ZSAwUehRUHpZ28PlPYu9U
qeNnxn7G2MTn4WNlLDMIrbidUDcLUz8dXV9i50XjpHjabwn19N/+iEmXFvKg2uS40RTtZXDXtO+A
ln072K4iLwKCzz8hYVVA+nlJh7Yke4863vhpY9ym+9lz7lw5a02JCb2cDcr85gWWwFYUfiLPc7R6
/3bwRkz5thYIpkDmpVJD9X+LSsiC/16Ld/m7fgz0yba8KvJjCoghCsIykexv56BCFN6u4Xj3C7lD
QGBW5DSZOnHcG9ADVGb6kbLK6Syg3udjQb/BnOc/H865vAb6Xi9dauzSVO85OFDoqpkwNqs3/K/d
eOMBWkROIF/RCIfDc16uv9z++/GI7XvbSWrD79HUsTL8/VYImIt/PLnOIrNDUQZW9ZvyMJVLtnJe
1uPb9SUU4QZZHLrEyjLlCf6hpMQOgZFzpMzwbMZShtxPfVW2kYyYpJlP5fQDJfAhCRnYqjwEJ23z
h97NW9amK+kGFw5e8lQhaPVexTL4u4I9muLrhKtNUGr0rMn2iedpo6gAGmwboXqZUEyUQVSzG2kV
F5F4JQCSrR1YZHvwlrx+LkNSU2xsejBUPqRblrtSRwVpTDGSLD85GiwU5hFL8C9PMkpogcOYzRDw
NvRInC/vEhfOff9lqzOQBOSLP8nT2OqQp6WxlaaQEeZtqbDMUSEB8FGP/jFxy+v53inNE0C1ZL2Z
BX1YT2wKMAUhYgH0b7wQwues6cnSDj8jWtvHjtEtQlo8UvVI2J+JsbNMzxdM35J6VVIqiEP7MwDH
M+IHBaA98dieW1Cgim7fZztvZsygxcO90rXXWii/4kDgYAYEQVW4O0ywInQEByn447VjLqR+yWme
pazPFy4GDmIv0rtJ5E9EKak6KuyItyolCo04O/OLYLDTGKmU7icw1ODmh1p/Z4kN+sbJYDmo6CrI
whnDrvsiVNUkwZdZf65JNO+vmiu96hESyVM0Uj58Esy30UHtwRPGcoC9vBPu9KBFrnhAfhKEpCrD
0bT97//ZKVvcaWjPAUyjnCCpJn2ATGPiJdT4WsbvgwLgkqmZfBpFo6L8MPaKwlPnue/ZXhtymh1U
thJRM9ekfGwG9FNrQR4Cc/gQiGT9d59XnIRbol/ELke7nuekBl/EOdKeYTqopT8BckldSTKWV7Qb
7BecDHD1r80FQQ+jFOw+PzExZ+gF1XiYlhp80iHwad+R91o7jXaNt76aYHlx8IoOxASxlMOn/zSc
WyUtITi1df4kRmSbi9Jqq6zJfDwrDmtzzd7YFEy6q1ksPN+12xZGfUrEWMP4Fi5hzI0SYVzM+qM9
7P0iMGXZa7zz2K4OoiwB2HcF+4SMfK/+VpVAWirxWEEZP/LBOaGA1vyKqcnKUHDvAAjMycdMiRtF
qbi3KcXnYT/6bNAbs9+14SmctsL5valuMJXAL2oJP/JAG0mhsEjIX+6NEkNAq1Tj0Uk6lZ8dRM7u
Yx0vUUy6iEHESP7gpJ+OEYMCGuPblCDoCcAfPtzmxZLOGMT2BtpNFOXZlA331x3SEk1yZQjUVr2d
u/8W7iG/26JfLlVmyq7zwqdP5gJnq9+HbjRYXuNfz2c7Nohlc+sDrYL7SD39sddmBstMU1mV3+Sx
omDUC46D+IIWTQfVSQ+B8uWG+pW9XraYzLuKi0k7gC1YXfHFqfjDRz8dWf22+7Xj6XidU7U2ueGG
3jXEztlEqSflzKIiwY9dqJrIjRHStKKedj+VzPPwaoP4m4uw8Q32U+yRH7/i+wet/5TWVaEDn2F2
Hg1I1Y+0RjuQ0uwB53XLZkB+p34s8yWETKyB6HoalreqZGhVA9pICk8hGpQuyj6fcyBu0ovosx2U
yQCYwGAlnTg2kTY1mp3hLNq3m5WsEEKQ6RimYdj7CfSY4FVQzh1KatCqC14pTePUY0TSdc25ZFGn
UGbZJ8jYsdVzvA+bp6Oy+3OZWQSSTnXZSCC0nRQjsfpsAU45RmbnuqKjY6BQGH5LQnHZIEBFr6YD
cL63IC3YDKmPyOntTAewRv31lE31tCFRVGSZWmKj3YYtSCHJ75l2Jf5xpGeopvgKQuCBNshWoZYN
AE2up7r8+/m7P/cHBHIQ7T7hU4ZUABaoVnC02SfErrrBRRwlseSuNkev1fpMZOE7NGiFKhlY4OzJ
bzVjgn/pmGIj1QxS4Gxp2zAvzfOOLvkQ0aAwoudah8QZc2VzbN4TejdKAo8nObdIvsOAES54gMwA
w8u7NVj2ySxwjpkegIa3EmRsFDUq6zhQ16dnVkOY8bnidoga6Sy7gXofwxEcVPWMEI3lbGKCPd7C
6citBrhJmIrxY8O/hpPMFzp+HUT3yi2MefhRw9ws8C5c1vATgly1b3hJ9KO2qFcr+HtSPnsMnDsx
ciX0LhvN+gAInGVPqHcsUkGh4MnzwXOpEX9aaGeJT5bHaSzaUjkaiw5AY4wNgBcCH2THaCAYWRx9
CZvTouMajUeiRMkh5yjSzfVEN5Nzy8PxdCtKik2iE1ylOpaCCTl3XW2vtqo42zzqcDnbNhwpg2/e
dp5B3DBSrjKdaDxh2lRdyg87TaD2JbJqKulvb0jlqsucWvTvKikYK3zmDlTJYIKZHszUcWZeIBgq
PaFxd2raUlwl5FHtNHBBcwZXOAnXah7utXmKBTo7U/IGpK1ksWh4i0dRAPd41xxv9RzmyM/dg6k/
vvQknnl+Hg5UdT4T8nsNvqOb3UMuD1geyYkwqXsJb8Cglx8QMGAJ0TfhgF3xCcmxweVHlaYUmhtX
a0H0Lm8oCXS7hf/DLTozUoRpUsJbk+mV+nyuvA7duQwsANJFysp7JlL+DHe3Pa1PRbPzd/BrxkW0
fWfk2nDKP4VFLKIkG2sJtWuovYAPVhprSdq8Xwt07OkcijUTy86txMdJR75XF1f+d3wFhMyl5Ok+
moqv/CUpHHzthsGHqoq8yc3YXKfSJ65vqc8IAJeBmB1h4i96f5OIE8yq93fAH8/HfBo/4ly+dBMu
xVZSEThGDMl3RuvxItlGa7lpaFkVLfxqAeKMyC48SEWJXTuHb8OLnyzCW3ykrGg9P2JJl6AOciYf
oR1IzjuS92tijWmlq8NHc/0hXGY1AAhiRiZk39xI08daCICIdy6G/FXXYd7bFAh6MbC3DtfbOvBg
z5h0OUlraHs+pDuiBOPADPiTPczRajWZvvZHkCnML6tnBDJuODVqX+dkeew79F9pUmVAQg1JH81l
K0LmTy80LrFcFmhYLASxS38/9sfyld5dE5wDPnHpVuvW5un6w6KIWj6pAKkdWFjz5wmloDpynlBM
D8bsJO8UrpnnmN4YP6fQouXwTmwQaXZnOCrnKUrHSbdyPlHaCi1/X/O4saUoE9oNdlDdRzoPHJjg
zoGIUQzzIbZxjQjzYVusFhUX1xKCoZqaBMDBmydTLDar5klalKkdariq79ahgi8Je3jZoiLB5+s0
qamtKaazX+4dQHMWFstWHewjAYg4lhgDozdMEVmd32VcbjofwHAMocfBgHRqdiV+sDuYYRji4+3p
w31Dvue/XP/3IOPpE9XuLQ3g6BT1RQijgwWI/78JE3D+FrY3XLDEFgcD0pzJbLnuOv1N+f6GnXYP
wB2theexTymMNBPpsiMKkyMHow4bI0kqCPp0qcNvkxOkXVQf8fJExYOr/TABSOoUxKUYPXXnmPNK
TMxMp/oCAJYuP+4XlrjgZoEnhz3VUofCzekFLiU1ElqoiHHxSZosxWg4LoePWBP2VVj0dEh4b2N1
Tsdo2MxFyncJ77pteSRMYzXMIlOS9i3nipfl4RAt/6RZw0sbj/LpALazjRLA+5UP/KByUKovy2mE
PQi/AZnRrcT8L+8r1FhmZ/liYLO1b4SzIG9ML8+rgz2ddEmgq42Jk6YZG3OUMlElbAJLm1Yr2EHq
eGIKjwcp1C5Xpn+JQ1KrjTof55kSCoBAVho64rJmAbn7SpABabtYGuGxfvhvqN7ITnKJgN8nJ4nb
zetvcnShofjN/1eWxFmQbSsw1d73ccdgouICS4t4KgXQt6MMtzWvLhdI1ETp4NtaCAJnCipWtTFT
LUNMEkEwir2QJAY/Gv2km4sIBUuvirqaaFhHAV3az1gDd18fI+GJoe8Rrp4hjXRGbRXsVJ0ZqDwW
J1GzTnIs53LdGpw1Bw23UY1+Moh1lo0f39D/5nZ0AMHFelxvcPZMoEbphJ398puG1HUHermOi2aK
A5OV69hcM4yB3Qd6TLO38f4shYQJYu6WMmeQxzMkQ4A4rloJFFQzxkGr/mIG/J9wvcjbOlV1fTVP
H+xecrrzD+OLbD7fEBuWhA5CDLKMobKP9U5oM+eQfQ3Qy6WEsL5Gs3175x/VjvHosikGjdvWVEFo
n5sNoAMqg4Tm6k6BbCSiRfyFrfJyW998gtv3KTVWS9wv/RBGTAKhXPda406YitgEs0B0PL/SiVP+
vp6kDVCkLgq44yDVRf7eqp0kw+NR6v4tVRLLoOr19MH1Pxm6Z7SZ1aBWzUnUNTJcm8alQVjeq37U
pqrWqqTBt9Sgk+ScnSKATGsw3mNu9KdxAsYil1CX83a9/D/txJYOO1/3yAA4DiZ0d+Jul/+hSAc+
T60NbGR/qDnW5p0FfeD5ZupyyAjzEQ4y46Jw6gqIt5qJTEuagbwc9HppN6bv3RxcPqKVjDrw2/VT
5zRITEhiispeLTh+1S/0Wzc1MtxDDoNQKTO5iufME021T1YOAFHThnAC0klEC5MY37++U7C5wM5h
D2+oz8JxyzUHVkrNgYU3u2dpvG2zBgaFBTo87BBkvwznZXC4yv2KWj5EPTObZMSDqC7f4Zx7p0qN
3cr8yogVdaQqKmmrcm21pHgLjvb4uN/Y7oIhxw1ylD8XbDDbiC7hoiQjSBz/Rx9+9IyL9n44sy54
DB0Po0nExHc5AaiYJylwoUDKPEgCITeCB1wluCwRJ0yFQqRBeTSidwtjeLZ/0Arvj7bEMZ6FX28/
lINAd1auB1OUjcoYSHVYNK1AEpKc72EUgtnJX9cE9fzVfPBlEkOZNQqCzT4a6QDS7nK8JULwEHri
Zfg92z5tvb0pLjROX6hVRJFbX4WSDplAAFkiv7uDPs574fm6FxZJ0pCLIid/XYXn4AH43DKLBwKL
oT0RM1JJBCBpA9QZkSyG2YJtaLPhrjaewMCn+Cfr2PBg67I49MYYHrNPROawgdF9k+vJ/sCqvDvN
UkAjJmfXQWPly3kWBVBGvKTv8XsrRSxsX9hQtUxrDGyPNmLDgndhim0XjLVqxwc4m5VYVBh3rMsI
0vzV/00EWa8co7ZRRGpZ46wKnyQHzZB2vj/9E7fVSi4rGwuZ5v7QqdSKGiYjY78EKQHbwTm465Sz
8JID/F5p1joR7rZK+NSHyjt5XoHm/pkrxXi+K4K9GXybg2hCLMtqiu2Y8zQYqixjxphElWZ1z8JE
m44G4UbgfOmSVY/TbMGUtQqoUHnudspCArCBpl+Ip4KL/U7IzV5vUMo5SNIeM1yWyjpJTWzyB1F3
HpIqze2CYjc3pxI358EytJOdmTgGian7D5ahHIQ+nCcCEd2KFQYeiOX9Ge48UmHKmUB12fC+NMgh
z8BpbjT2q5UtZhkxBE21ZcPkefFxwEx946adM4MEP0ulAHHEuLcx2je4cK/TOBFYjPvhQttimxq2
BfoenNl5xfw8mE7YABxZGFywi/QVgfMoRURoc66U4AsyqbPoMqSD8siD1a47zN8OpJjrRIJUTILy
Tg2i0J4qNkmLUrdmGzsw+6ROGmKf4JCD6UqLtpTyCDZYT3ZjWuN/Sofn2demwacwcRgrDRVy6LEt
fzTKA+u59EB2GbDmt1OD8Nuql473bQNbeUEbyrPQMuM+MfGt8EHKTfwcFRwPIzQ3/8EHQRrTCyDR
bR+TTDAccVEfXiVsF/Cl0OrNSU9pIRtgun5DyyKtJnX4kilsxCODlu6pQ0DFEwsktKfEVV5PBEku
1pNYDFsw9oFaUYayqTZVmKvYxk9H4ub5xrsic6qH1nDa/E8JVzQQl9RNomsHrv9p6GL+3o6CmpZq
sbDpcijv+F7TLCGjmIW96X5r8KWT/BKs4f7i6vPs2ILmRU4wwy4N/Y5N8v9mw+w6faA3SwT7htwj
/To9kqJ1ob7lSej13xBB+gtAcQpjOZmtn3sTF0xyPz3I8buAVj1P2XvT9zxeF5AJix7BVGx1DTZw
ZQpWcc5nVxMxbx7VsmnpneqtAGhExC4wWEQ/aBDnw3HX2xJKz3eoXldMOjPwGCqF9c0b5P/beozp
TrkZjowIDF0e3USu41odKhYjTQ0JQDhmpFvRtUwXZx+yMyGbAyN72uxk1ZS45gUlnad99kUT0O1y
DXKQoSkCFvMMDK9KjdZIsuh7JOdNll/e63PB+ZXMEXDhx6FiKRV2I0K91Rj3bfufEuDnn3VN1LNq
E09cEnUf3gojYxy17Xcfx2Rk7CBT29d6BomAGWxeF7PmJtwlaWTc1xaBv04u/trcD7cGXEeQugya
SZCgevdDb1CKJsQBrB5QH5RS5pdvpxBdwxT9HjSVnhZYHEfgi5U6UudotWcjNUWSpqo7/ABbUsUC
rjz9EeDSZ482RcqGrQLRe/zko2FIcENm84aIXhbp1+S2ahc73B9/Xx5DggOON77vBPMFPoTLGIch
l62/Up0GueaCINdalKmQpAmlOn6+DuiBCFfZcyiQ6mpT+pMRPM++kTPglDNBs3F9FnF1mr4Ij/Tg
SKGQCN297YKiCpk8nV/QEcsG0UBKbuuHH3G/cQpcNEmnhwLYWQY7fKIM1bDLTIYhK0eRjT0UZEKz
qHPZoggpqUw8hQk0fI2kHNhWERdQSE/Mr34jxcSPf9Fo5KtyPnlxpRYkLjIHuZRh79qEIsUt3YOy
fN+ZVm2IdfjHYwQB4fN3gQt1m34wErvry6oV9mWg9fskzynEdl53DraIXEBy/FXt3YrvaVnMOU17
1DDnWCz2ErolYLl+zMM9qMIqaC3+9nm3F8qxeqqnHy0ufafNwaQ9XNxnfXf/7F/XyPQkdsrO1IxE
0XdVqIUukTh2mgrtmZYDSSpx2uwbgDZ+1DYsFbAb6gh3SKGqVIuEm5EIuLM5W5gB9/QYvkdoU5o/
cHgBPfJt21CYPx4v3lI6x64XY3Yf8fVYZj9EeG94DC6KB9cyMYof9XRX4VbOtRM7WzmkxUiD2qzy
4QkfErsOvU2RFPyeQgkverAe6PoJeqJlBSho1X8PRKIsDT3VN/jtMDz3UHrWIKaU3Qa03dYLVIoP
aAvi+a5EVgF2XEObQ9r3nWxPOSOU9XMmNG6fZTrqCPLBWhlvckILXpZ4ATOmNO13I8n3/Cx32qSW
n3TQVbYm2J7oYwqF9N6ZYjpoE+4hdY6kGqOZ+skC2RsAFgGaw1S+8GGOedHO2fM5xuMft8sOv8Uy
TBP/PErX4yvAz1TjzjYv/wCyRmk9qYskVVLwLoFlSOVwCFxIIch8rNkhw2hQ5tRLLAD44iyezx0L
wybS39c8iorDNdu4SFd1MMzDRqvy4q139ZNiIL+PeimAHEB/WZ4ccI8iwQXHwYenhFE0BK7CaHsQ
ZLv9tOqAv8oQRuqljbMN/QS209wdA6TvhqX7BX6012k3SOEut7aXYLFlmDXHSLeLnLzII9JC5gHX
rOGSqS6Ao02LxKlIbd6uP8ixxBTmZ6EgB28j5x2ww74aqoEmbLUADuQbZkswrqp7yiHH59lSgC54
/OQkz4VJ9J0fNdn15JpPtDEx3KPcEGaCegWV+eqj+kGsa1/cIMQGGk5dwhiU0CixKxQeBz0W1U4X
KTmJPJ4kr+eiSMPaCclNQicqnsS7B9NpO5qPEad4hjELcwDAMF2pE/rH5gWisBE8weUEq+bnd+ow
T/FpG3VwaDCUfKiUCvq6+rRsmdl7Uiv68ivCLqKxIaFDJfuCSa/uz4Cpm6v9jmHcUxWV+6uAI9Pc
Bv9YxIp4kkviUoKkWxCMx0JzeOKIIjPh/W9ZHrK3ovu/EYKNrC17lHlKyUIwtJvrBPo4cb+vvCOQ
79vWEILwqlxCSOQiW5pVBepBoIuZD873/ZEvRKPo35YPdpEp+Kyyrq60GO+Oe73BzAlD8VKHd5UF
BUhpHg4JM3LwetpuedtGfkQ88IZ9TXUTx9W6J0DwqfrG4T0ZzYrUPobXFtzgxpFu7OV/dBGK3vO2
xS1EFOSmJFDlzF9Fl8oB1uZzbrZmeFdyUZrUkJXmg8yKhnNEI6/rKjhvgySKCs7z99xp9lD553Zt
i88NkeaDOtzPwJps6borTISENyxgvICEIMkjXCKLoEXO06DRsmwkxLDh4M5eLm868jLaGb82P0oz
fjtS4h2rSJxq96cRtfYS3ebxz1aqnHGI6MO1z2qrC7dBIe3dXVWD6XhNUHPD25JM/fMSX4AndzWG
hzT0Bzy9P+4rjJ+WzBWPco90YDfEA/JsBZc6TlkQ2NM0i5H+9xja0IXjQGXKuvgTi/LKVLzkjmN+
fzRcBnIyi15dMhYTdKiT8TLMrU8lgrfB/cMcsAprt6yI190ymJYcaGyP4tGLx0tdpWFIzhMXcX1p
hJp+jiRAGyt0TX5DdvAkqsmSdcA3fE+jYpjAHp6Q4U0FGJHi8hFsltc2Zm1e2UJHf2sKzy/HR1gm
2l+51Ce+cj4Urc0PffFBnPQXxkgfV39c5LCeTjcQkLKr2QMPV/9OfeFm4Fjl00qfiGz6ZWpq4rSF
z6rhsdh0RFH8iVSijGFvnRTBqNyFUvslN60Dkx7iA+ZRbk5eV1zIqsIIs9tdGLz+L4hWMrRhyQ14
zJBGULkySI/Oz/5VFCXdH9xXiXCTuh2NgR3GrHl4rrt52JD4gx5q+6xTXKXlGQK40vrSmjF5lBo+
Ym1cwapnGP3SSMCusPu77ta/ixR/Zq4jr0FiyZtk5P7yNFi09BBKvBVnllOS+T+uElhUz4ufcOeT
jjhLE5HZHavE5B4SdKt8q9Xb5XpDcTUI0ep6vDtPbcwHp4Yzbq3tKILvBOmMCYfDxKluUDZOY9K+
aYAtShbpGYPouJujLpM0jFf+A3yoNVAKJwNszaucECOeGXelrkziusdbm1V/eFKOg1OtdPg+qK62
eilS5sOEf+yPiNozo+d3UYdKdCcbgK23RB9U7Ip3VBuSzQaC2CzKBqyGfZD0oEjnW4v/7pNROduT
VjzK/Xo83CF3OVUIMtRjC/VDlAw9T5q29Q1qsdUucEyS2wrFp05CDHzX8ShnYzuXaQsY46ME+ydk
4NIzNZsj33UYKnX8rd3ONlOla7uBOoguJnv4CFsX31ia1FM19TOgjmOYHyflljlPLxDHgiGyjuN+
XYuf3QAc5XfTeuIyov51BOokpSldpvgaeOMfpliSSeDv1rSWupB5+GlXbhIyiCGWi6QuxakcEFuk
NblYSa9TplBr49PbnL7q4eSVAo18WAs0f1h8AkLt2zNd99fwrz5r5t5N7YzGVwAGx+OORTQ9XPZZ
FTMDsx0+VNXEM9m7CV0Ke7auyd8QDsPiUl8K6c7tjcjwqkFXXZF/H1j4ko2aMxwwE/aLfYOpN/vH
oXMu+7ckmsJnlsKazT+S6QfA18w7jiq+rPVxqz7DD92KpRlJ1A5jTQgZbikzwZzHXZBD2h/voUvx
pOhnxklLnUb/uVRmK8iJNnbGTwj2qs0MUqBNmE+hyuMoSM6mB+5ctrLhWRpF+HWrkWmVrbDOet96
X/8CXUWSZdoY0YqFR7F3eUcBUdlMMmx1Sws2GYApAw9d3A/qeR1OFu6vJC9mK//qbWMkX30YLM8X
lmwK/JHKFwbsQ1wmRSYKF4+1rAKAQPL9zxLQ/QzcjwFvmPBzGcfpzmkL8v/Qf3DfZYpiikQcO5Mu
TJ/rPbjwrmtzXDnDWWjMzmiu6huWjKSJTmgEwUNhJKmavIBmlDHZO/3ShPnVVLwGGmKXEUB73zBK
cAExvBwzJwmO6tkmXmjRDczBuxZSk9UsfQ9pODDO6nSrw6PiJFsAEJ3YsGC+NXanqeB1bUeo4VNM
l3p50n+NqlloVIO2XAQFM5h/+tr57ZiTYXUxl5E/3UO+zS/3+7FpZ4bT7CrrX9O49vw6ISUpkEiQ
vFGUSW7wouOG3K8M0KQbmY5H7oRDI8Oe86C9BZyS5/9BtheuqH2YTWO6SyhFdecXtox2kcVjDaMH
oLUFg72sVc1OPNhwReR894s4M2E3VLozqRs0oeL61hLsQz9XnAUyl60u16+EbKPTi7ZP7pmbjly3
mNvLPn+iXJb+8I9SgZS5NmEC1PEU06TZ7rNSbdeW37rA17kOq8l/uy832CyZw6veCTpfKmH/EHpP
VuOtG9Pl9lVQTdhA0UQxeN2xL85Op/IpYsUReZ/z69f3gPi8sKzi0/wORmmQiYxnlG8BophapJ+3
DytADoBRfh8Ic6yHuS0cr24olzxnpnRmIeh0dykGGyv3gBINbd519AO/56TKv8Rl+udHJ6ecCkbn
JhKpYvKuNWEeWH+m8cdCemSJrRwSBSkcj39eZRzs2/BpJMJLhCCz2Hr4YJM5KALnmu57DHJ2LSFT
h9CRDpfMBj73OsX1WxGKI0wg6JDOca8lZFGl0u85VpJHoz4nJ6K8GwTIwTC8uGWvY9YPwt39gxM1
6Cr8yBYiD8mdbjDR6PLsvAwrftFKDBG3a7KKpxH7j1xeyzkQ3vMgWQJVM+Zi8q3GjfTq34lJYmSn
gwrB9kJxhoLBCSzkCbcS55IxVl8C/hXn7/gmRgiFPDGeoUepj5NNAP0H3nibJRwPYUdxdkQJHvQy
wZoU8aFlgsB00KJzZ6h3x/idcXa0ZIgqbw7zpNinzhpRDZaNoVIaMwIv4Cb9cSiL0rnr/Psigi+t
4c0Gc4jLoSR3VrktI48mqUULlhxm1rBFWoySK0YtHchR3cabkFVWNdK/ONI2GsJEWfdq3xP12M38
OGqqkESHdNd5DezctLJHMsv73pCt0myq3TgKQEknH7iD1vkMQ471Yt96r9vvLM/AM+vl3k5C/SCJ
01tHVkwo4ifhvcrV6r1hyEcISh5S4KXnwbh2mmnzMD5bE32/A9QFXDEKECjNQFaWoewj7UXFiWgG
SlSR0SuwzQFFrFez3plf8jV1c/FpOu6tVaUFA47ihoEmH9/hhzG7NM1tfg8TCH3cX/RVszroaU46
i38WuwcV/C8G1U1Ag2s59/MPDQWfXeX7LM79xT96EYBa0wsBpeKZWmt+DaPj56/Q2tXpngnJcgr9
NqKp5AWkE8L6QURxQY/oFnGiY5PuiAje7gep/uCoi0hN2md8D3h4lraxm/NHRmlH6t6UBoD7IFGc
fAqyT23Ryb7Na343kfByzGc41EBBzizMjvxLphK9kyaMVvjRTDEVzBoGUoN1vmnBeFac2oyWQnoP
KtXmQOMyJ/EsTwhfV3mgyoIchATCy/w6QXK+YpMbiFUFbkrjoAxJczUenNxqmr+MPuhmYwFoipZ0
bBHu408R1OUVFGVGTmqCJWmqXC4nPWKCQ4NOMjf87LFZy3bTryUAnJzXjFtxN/7T8BjevvhPsDlP
7/12YcU/TD2YDCYPQUOvpXhUFDEA3kaA/GEfyrACQPGMPbFxHfAaUcR0cOzEnJ+prFzBNHXIylmv
AZVW3ntVALR0T71T4L4hxcaJw6s5G3Qnrm5h7nYPcRDGCj+QA2CArTJseHHUYWOZtn3/LrjuMbzz
duYL5Zlk5lZMaU+70Hi+9/IvdFfrJ0RfM82KKVFUCEtc/4W2xQ2B1KYHVB9fibf2Q2mbA9fV5p4s
PMrKs7muDOIz1D9Ncp92O+zfXceBv4UmAXVtAAL/ojadd0JUEEHGdIEir3/dlO3chYlyg42n3vwi
Bh2svQfcWXZ5pTEuFmnQhiJ4yfKUK8gvOkTdQs+BSW6NOhHbH7QhWCV2IRV7b4RsEqN6Tb6gzNZn
8+Ioy75IJ056Hkg8jiD5Geu3BH/vRKR9nmPHN1lo2Va+3Ye5a3A27rYQUiDZX/jXdHvjPItOI/a6
bogfG1824ULeuuFE6u3roojy2I1dU56zBBRgzX+uyMQ7g7/D2LL1KfM8b+JHBfNCKZUaKhYsMYjW
h1sxbwwZquVoaae0X19Jbskmj7XPtx9+2gLt2OIONyrEkxIwt2Jwa1pqOJvgz4c5S2Q0+qg8zQAQ
Y1a+LaF6MnedVlmHbcooq//0m6xGethoBOHY2D4SCVO2Sxxaj9Gu7JiL8muLgExMcBhDdRSd2cM2
ZTOP8yDpFUFDcb1Gj4coRRyTe7yutCQuOPCHtroDH2qDJeYgiKbDzF0N3crpT768kzkSDb9+p6Vc
OMO2z+67JJoj3cRt8HDsIUPzoQ+dJhfYClsOy1iq2TtZnZcUrssmUUnF7RVPxnLPIbAHOO5XUWN5
8Q3iRhuoLcAHx4duG+Jveb+HgZ2HQHunQ4LEdLKK0fx2r7cbGhuYpObfT952Mtp5jdnUysX2+6WF
JJsp78+C4VaEDTE8rer1+M6qj5PiLqn5LkW0LD6XAZQJKfTC4ewv5DliTXrFB1fvvLDtJX0XW7ac
BOCkdcLGTkBCTNMR6/FvCp4PqmxIRNUXDK/BpHxFZV4/vozSlrbzf51SwAn+RMjx4/uN02Q9Z1fR
7/3O3pvsYsRUgW/nUO29vteEnlRhqnYAB1GDfmBE8sL2uiCjL4xBb8MSJe/0b6kg/CIQazXwIOOR
kcKqGEFAET6CKvxbLibOVQtn5PCKYqTiMcuNy7J+LQ+nRu9KUQxewoAhNl9bgK9lN/65NHuUqRLs
XhtE+vDTmMzd13/QYUwcBg881WfylvHjXR2Cn4tzHQ2pLKfr2AY/19GE/U37ZhAfX0C9Ujg4LjzB
MDfLVlhAZL7Z3qcDDdLG7jOo6wwOxkULjAF4SjvnVyOP7sFqMZFFJ8334j0NyCw2D4efJ7S8W5Fx
p/cURi0UGQKr9pAl2TggBySKTlacsSlB/e3EH0W6paCorPZLDsQAkj8j9ixwxcnOIsDMln4owO1f
BLvGg6Upo+N+KtpAL66NO9tOWSAXwiBp8hMbWFin7EBuH5EssacH1psi18FmGsUs2bVU5zMK3sYW
rsPGsFQ3aCnsx1XXYkZvzJbL1avTsvFlgpGRIkWeG4BCuGUlpdwXc0AKxXIjJ4RLiOqtBpk7Hv3R
MnYFZ0P5kLZDDtx6PVViIsKnO27PVnN2VAywFXVReY4HWBfYK0fhRU5CEN1OnJHJavMBiPGd6PiV
vywDssfHtuinF4Mx2XoMxRvWh9isoRNowrZAAJhBFaOKqwA7N5EhzX4HF6EZOGkXRsm7XZlEcr2s
qX4tFSUS/nXWghPhP3lVrJbcL+rAQ8w5xzfI4GcDF2TBcEqXmDQiBAIThxQfi1vWFT+rw0bMIrKt
QPC0ZZ6kUAhsMYhyYAf+xIdhiA7GCgh+8A3B2+WvhJi57CBcIzCt7kEERxc0CrZyQoC1rofa0NEe
ubZDCMA9/zPii3EwDcRZetzuno22JjjiGhxD0CQIM6kTcnsypO3ENV7wT6xZsW8dOvOAQGuQMUA0
MUnkPmB3GaF4TRLeg4H68Dbt6/Neb7ULpGhbNDPgown1qLhaTo+0trFweZEDOl9ZbU81fMTnyJ9a
7mnfw+npCSRcQo0xthauGVLFQmHF3MklMGQdtrxQOkxpKv4dNHqrWMerKazk5qiV0Rwyy+0BAxJ+
278eK3WrsmhwvfqTHfOekN326HlbWIkz3uZmq9o0LZjSveyY15kBFpfSpjxlq5voMO8P1BcY4vbU
s/1tyolTtQ6J6gud5TlbYPwkBDGH+2tzSDGD/BAhDErG6Pyi4rKhnvv7MKT4gB02vbfs5ryc6WZB
Pv/bkAcuCLIx3IFxOi6kHAmBfMSDMUoCcmT5Nk7MH6py2kE3HvigafWgIww0LP0JzsFxzxvhAiwl
Mk4dFcG3yy/BG/grcHOd+xw9sE9KzEsSpZ9DS+fbwAdVU0gi9Rc8gmNw2aQQu/R0YlRONDBYh4Oj
EyMqIpw84JaHiFD/GEe8/wqwngX5Zy/5MpvI6AwZ0+eHb0j25O7Q4zXR3KfIlX12w4GevRaaM0Eb
suAUDbtwTWG58Dep4tD1P5BBgzoadhCMDhvRoTjbacCQjysNdCFjE7+TW+HLTDFEKRpyQEI/sa/f
H2bM0MSBFMdmIZXn/4TyXQS40ooss3CwjLyN3RPG/ToJ7uLQPCDWmi3j9i1MrCJ8EJaH1EPTZGsB
4ZIyYFXWUCVN2w8y2tzyA4TV7FLYjoyGe63Q2bBzsNgXVYaCtOR8PjfTucheve7MjbDmKgfDEsZ8
SYsWeF3mibc6D4w2Rpd1KZ7IKKa1FP8R2FmfA1N+dzr05nbqDRwZb5o20nhtw+ezPBa5Aa6cE3oN
jjSggqgYmVDRiYsMseOXzmROUNUhrXGfYDMCVql2Dq8hTjnd+6kFuJTmVSMX9SG7JFJORrWrOuls
wU68gApqoSSqhwtg3JAGq7xdCoL6t25gPgj6PpbWULzTFhWJ0/I5m/HvgGiCBdbpHLpwVowtPZXy
WDfv6GVPrVJZyWt2zeq/QYzz1zkONIzqrjz1RAraVx/ntQkkcI3NJBHHm8nf5TGWMy81c7PaJOXc
oGcOyvZLFxYm0rBzunkOCCCyas8HU/YXGrPHluMDhSDjmlOqO/y34INXX6QlR+XMAheVI9S2zWK+
W0Q2i2zqbJoFgp4gUHCIOXiXKoRWEHS04O1hZ0/rFICK/QPxgbuBQ1K8XoS4E4KWZEcF/WyxWGIy
HWcOFYpGOlRoEo/Iw8bvxc5EdXGMvMFdPJYxwBrCh1FQJOEHvkQD0LpxKe+TDM1a9nXfmQIaQnJb
cYYVKfSSKqF4sNLbI+s1iMZExSnooaB445QX2sR/1oJHxTgFfwo4RktC3fzwFK1bPq3M6bp1REa5
kdx50PscNqpL+UzXpNJoeaTgVFC48koU0pBq8Ye4B7kVOU0JbGRhohI8cWdaf/9E8ZJc0f4hWHd7
9TKWTY8owxUsNoJYIF6Ybj5RF55iyPGCtDPQbOpENH3W9GOZ58+mkr4m0NWD/QgcNeyHo3WV4Byf
6tuzhO/XjkeMnj0RKqYAZj/UaxjTnITcRctt3sQxe7JqYp5FpJGi/dwtHf0KxbGRJF7wISg+QAz3
1RhvzxIOkMpZjXeb/cyMZzmVzo4UTZdD5UaEZ+IWIGzpZ6+UXatlluKn40E9u1keqsQMy+mkfRrc
8PbMPNhqXp+7ehGdTrbytjVjX13t4IBH+oDdHVciHfW7lzrEMmhcXo/TCQu7LmVMDOiWqvxnq3qX
Q+wpuvDkD3QeviGtEja5LzN7fU0kVmSiJua/S+CiTtPSLFYeW+cI5CBVfnKQJ1MMCSViu3WCiCBL
gpcmAMWT2OjqTKSszi74SfLhkvY36/IR7SwjpR8lqhEzd8dD86X8pgSpxkzq15u/vLwEvq6wcJEZ
TKFYVBT5SsaQMaT40GOBhwZ4AoHGVomG0rByY4s7eEpv2jmw8OoGowCoeECJE10oiHmSKS5R1bPi
L+9kfmjq+QjU67LcE7v9qOSHwpkb2eClR9MKxdTHgl3+ddGhh7WACyOMVUN4J0Lv6xJlEwzanNkn
qXW2BqSnlO5XfldHMJN3Z++pXXyOjBI2j7dHUTBwoVJe7jhnWz9BB+t/61Wnwc/wmxgKo9m+Ybp1
wsKvHRknTrK8nzmM8TOMaKg5PpRH0SyNpHXv0Y7W3nCrxLJ4b9+gJngTBKiXknE1p3KRNZ/R771R
atPXP6xG8KuHxcDtbP1XIDSIZllHQAMdUMWUCKr1WMipH37XlVOXX9QRCIO2QrJhSJd5RgoRYgGz
nNltiVY2lBJraoR1RRwPtuUvcXdSOwumEoJ39JqsWWukz8rnSbPjkJ5voaqdKeeQOCipGaxTNBe2
zc/ejdl40mklvJJMIsrNmkm93zLKFjLNVepv98TO1W1MZosmD2QuDvZ+BZ9DlIFOyr/QrDo6cogl
utU/2FpJxmmgpKbKIdK06pADF4NjRk3mvHWf3bIuAm1ZohAt7+iQZx5E5xZttUqlw9xWP5T/xkib
mAjjxxPa8MlktMR7E+9jl5VfwivqDnyAprr1e0i5lgwh16kRwGqIP8PTRGp/BEWNDdbsJghpP55V
FkE++mKcMny09iSFSu0Fx9E02993cgMq2l0yZnlOwX9Jk+S/IJibnh5p1ctO+8TGTwHDKfWf0ak5
wM6SWmGZMK571MjTQ1vehPvkQ6mt0EI7IgnWyFgtRasb+CcLD5f8WL0o67lsEttxBo1U8Mfe84iR
+XlzbjdutG8FDbkDTlzJdFo04wdLhxoSDhK4sbfryIQ3opBrKTzzZsLjH3HtShwiFlxLRF6DZZD+
Ad1lnTIXdraeyCph6HsI67bbBWXb1d3g9fISXWUaiUoIHTLwKUX+8tBX92oy2tflklADG22Ivnpp
4naCTRtG1BODkDYhE7HBdIOrfzNVQfkXnGJh65lioDPn30QBLwERK3xvd14OCTFNP6fkDinHWoyn
syrE72KLcOBwUjLMBmUM5uKXTGMSzu9pzM6GL/gRn123iurErM2IhZhR8pfMPS18TBwM1LOrgDCT
5y2NwPRZkX47M/3H4ZTYjSo56dEQ2ONshN6Yb1Ul6WgmLfimRlHXqHB2ByLrW6IKpmXAtMOIzP8n
4URjueKOBlZcfHsjH9UVqZQm2z3TkNMQTQ9WLDOTjlW8ANd/bgsBkMd+EtIDyIz759osnZxg1opy
tkoSlfvK6N2stluZ9O3gm1RsOGaSgz2ABxiDvcF26rgNmUIUewX5KjJ7YiT1sDQirSp4CYKlw5Lo
v/8jq9Zc6EGAg+lSl2/pLu3ZhvsjMXe7sAsHZkfVy8c4QtcrXm8h/hKokJVZVn0xWGM+bb8/fYoP
xqCF7/qkG5OLKEpm0/bT0K7pOe6BVsIRfW0FYBQvd1Ro8UJH08o/xqj8AgBMYDV6oak1xuVW3Qxc
l0HfFqrgwo4K6mNfOWOObUQNOdUv6h46btqkTShq1D+ONK8p+8uslwfU/bp1wUTcI7BfPY/lGDBf
nqeRIWL6mmw8BjuOuMVsyy4L1k/FbUrQYySLaJ0FlZFoxislWpz8Kzt1um5jEGk/Rw3nGxlR8+aI
7lpQ5ZIUVJxMoh4w2bulniciSECOm+pKWk2ycpacltrXvqVWXdMPYHhx+kDubhtLMYHsA1c51CnR
s4Y9zJbsQuoaRRCpE5rcSvopuP7ro7rxNXGHxH8MNXuJ+uoX/9BJxaU8Up/EdX+VL96RR3BE6wbU
QE4ABrmIZUHEWBeX9IaQgJXH45jajAIInIAd7vF0rQENoQab9JRu5DnItAKGT8qh2FvBlWKb8HJ/
arqpsSFTYguK0lADxGu54bY3eYrtyNjucsOCdi2aTPqYoYADdr4+M+f+hxi7nQpEJMJGGpdp/erD
dhPk/+f96QB5x1bxaElnuVJV7VFP+dJHIx1Gdjxe+JQPhFiJeGV1Rrcc0IC1mhH6Bgdd+ZIFiea/
/TTGiTAGcgRtFjVChLQX93tVXketZTDj0YWpxaP6bEEk05P7gVhPARQWNOo4ub7rRNVusHRo5bE0
Hj3ccx0L7jt9WSOeB2QcNCJJ1HWuaWzPIHQVyuMZh/u2Uu5LgeYjqm9hbubeP+1xVSFQN9LVftVF
6j4ILOvgqlen0lkLUytvhMJN8Iv8jTBDlQObMd10GVVhHNCGYFFmkLkZUTVnXexGdFsH5O8SxTaG
hp3CruDe8Q63yVifQePcj8m6Q5SM82z41BRbeClFiCz4EvnBVnAaBfxIAWF3f29RllJiX8Mm0c5e
n7fJJMibtFZGGwln5IEvTyWuNly0jQ8Kdv1WZXm3UUjWBItV7jIXy/ggoZqDfg35YojjofILM1wM
Q9b2uUCxeYsyhQnq1ozGoHr7upPEcxacYn/8HTkLQAPnb88EEvm/ibVMGphVJeH/wPc3pfFf1EkC
k/KpGiXvpuhN49Mksc8b7q25KWMRqaoMN8e7Zajc3/YyIQNyfZON6WHb2X9R8SaAWtnSql8pH2FZ
dEWpQ8v0X7YXNTh6k3uBix0UiwO/GgsA9dFDBAfl7m07lkvdfihg/xh8fiKK2jF8f6gbaHRxYACC
Xy5AiMcxmbugRx3gGIxabU2MvN65MK7oZORjdnBA7kb3Ehusqh10BN49rTH00YLIEtfv98iEH4RV
Vv7XpUGsibfOb6/tLuM3y2YZBrBuGI8J5Wrqn08+O+9s7hbL5rNOOVjT3BnW8GCsBr+IKzs6gEE+
2JvfpEL6t/hDkqvdOeD7vlmm4emIeRrjxeZFBHYYMflPavR/9OBy3+RTWyAk/ymhBDhLs8XL9ijN
/7ygHQc8Vz8OcRCKwy5kuFnHdot+Bcx9YNyQBgMBalaggCalRn0UpVBCmTsHYJFXr8BEghxX+//B
RrWOPbAxunetrz4WQlfSdgiOqBeR4QQzymtaptgGJZqIHOUYrtjxLhkJDj+wgUpm1VdTWaHgfrKM
6cpCUNlanJC/pP3GAxqmKWXbDQDNeETJCSQE6gwP3Q6aK87qw25i7sPrWss7BZrfG6Whg5UtRE/y
E45PprQvE2MxEdzmXGhZRTrdehmIyLP8XPu3geHSiFBbs+3W6KBzjkXqaqksPSr5PzPIOnT8FY6w
dkJqPoTjN7snEVxoijHquKm5YnaoKdXcFO2Veaokzwj/oP7AjHBcErHvk6QqMSdKLDkfMnAFG9Nx
T/prEnGhyav3QMixVmHpVYKYuvG1ucq6Lcp9gJ41RgzHnt/OMgiL6UY7wNBP7HHYOi84bk1c7M+T
clk4LwaL/uBQdII/H/Rgrf4uM9ApmdPJ8hcmDv6UQXq6o7it8UaGaL3xbASL0g7eDKtW9wBWRJui
BqM6bDAzOoMN3y0JYlg2A16Rmft1VTCS3ORu9hjWgbz6KbKdfgkOeAKfzv78g1nhNtdU4EE8SCCP
aoO/xKWxrGvpkQ5ELD3ZCm3hq9vqsn+1zRL+lYfBwzasqZFM48yV8WhRMTSGhbmERuj1qsKo4nBh
9/ggrl5fc1S+V/P+ZMzgwmBloVmo6XANv5oORqoWS4Zm+S5vqxq5Wouj8QvSVlFOK88Y9Zi5LPNc
4LUS9OvotNiObWlwHlpOa69/eOsG1LDKR6RC89vrb44wyB768fgU/a5ONheJQWuaYgqF6J5lkMsX
9IgFhrAcZZnpwIAKImB6sIuMDvvEgYB1FqYcB0tuWyGKcDG/XisTlggzP6HaP0nE6QHvGI45wfDI
V7q5pcR/PLtXkShN8cCxmmWmZx3bdb9iYkgr2Gq97i1DYzyWhpx+TBG5ACT9QwXS6qq1y+HkJs1o
WtR9AwuYpil9idiJ4kJkqYkoLbTmZDXFDuPP4H9AyB3XUqpkqzufyOHbregzOtO2lFnGgXb/uNt7
z/9kAdw+/KAXh5K0ophdSkE+nwAHtyRyC+AUzLUQYht6KrRFr4Jk8XvoIQXJh1kVXUsabGlZuBS+
cFDU+UEJYCVXgUooCNrrw4AW3RbYzNBz3ywv9CZI+SW4IhpY3t9j6p1m5MMvqyKZE3zztMDDQTtK
b6q2j1OeCRmC+SIKx4MfAbl5kdyBwOlZreqhjuDBNaX1at5wryOBZSoJXkmhdoFueX8aPMEvh4Bg
IdcS+ixTCFNh0P7TMcp5S4BIU6vY/b2dPe0sf1o2BKj56dKUekvDjOyeRqt0XgfLf9X8VGZvfhz0
KJTpoKOwEYaGLheL0uugLY3ERdZZbLHMTUnxcoTOOU8LjZh6KUJoW2dCZxOy2MV3e/m+VWVG98iV
BBZcnEk1EwJAXGD3vPZcNJbFgVFRjNOIZFW9azZW82vEAGRSvHDchPlTtQsQc9esuTGwjfhJBNNM
F9WiYYSfFb7x5C3E/VeohSfoPt21heqblS0zUcwB4pjudJtA2NK4ex1+27WlCW9mM4QLNoSz/wJq
SAuddw1URepLEmJHYgnBg9C9h4S04Xh6Ivj/jMOLewKp0y7uRIsVLC3mJPPvPisgxiX0rXw0IXoq
FamvKrwZatKsOEa0ypvF5isHwXsw/hG+mj+hzbk7TYAU25At/Bq/t///i0VSM/J/H8xsxL0qHP0Q
Nqp+sm6Fhu0I4a/ejeXz500O6PlGoEgQbTzEosgKSyr8xB/JD4ZKuitMjuIX30eyznVPj8Sthe+J
yUsYIIEJzhqBd49M5QSaObwjaDcakHcuIa/Iq3b9eQpkk/xHsMWdzXocCsi7kZR1lsK8XYqwW0CZ
gFGaOnbCPUtcA4UgUI7JZsctkGUFFbSoHRUWxlcQaMXzj4mvSWZmqKP8O5z69gNH19VnZ1Rwq/gI
VQibkGhhDSRT/X3DtsSOrH6x4azncT+wMImkpOWsCXPi70OrXOIVCbvJo83D29zUhUTD2ea9g8AB
AI9qunyWgsydocP+wwCCoeddK0/nkJ719tvK8dtzvdi8vN1+8kEI8r/Hqd2CX1eRjTfIGiQF0v4e
/eik6h8izM05qeRABgVI6IdPbLwmy+AtTKVAPD+E5piKF02Fha24JZHDBpQjkSKrHlXDAC12Uujl
/vu/Nl3+l1MKsGk/7U5EKP/a770HhMgu9/uWHHoi9sRoPa5WsAkciOu9/GzyarcZD0pfhy6voRxh
YFG+iR1Gn2nnfiUjWJv80uZ517HB6RQIFz+nNPUKmZYAcRjKR5SXUOqEKvUZB+MxjwojtJWSJA8L
cTqAHzwteM2/RJaAukm1hLfMJO1eN+sO6v6qUJBj4PPBafg7J+rY3s3jRnf3mJJ8b9h7Z+NMhtka
PLPk9mIv5R0fHNefCLqJM8oT0Pnkm5CnKTnUVycKaeJd4Ujhss58TIw0V4JDRjWWsSqqKj1OqHRN
XeUEa3ymsAXhb6y58zz3wXP1tUIoEejIxXcDYYjIdXwTQ6pNrBWvd42NEKqeE6UzFGHiVQFS+YL/
RvnsjFnJYnaGmBzl1hGf7i5RfPIAdQZinB+ZEV3NcDsY6ZpHzMt1m2IxTtUGmjwMiyLwy3dj30GX
rrpQ08E+gDKwg7UsR+/pUO9NcAWNbIa1Y7NaqWamKWD2gmphFslE+XR8wB2NsaBBr0hTenffXQSY
bObGpHA82vkgF/wGwMl+I5lAeN83g9qZ68cjf9bBXxx6F3xUqgBQJ6FsikLDn+y4WOTVDt2i2RUU
OeCdTbZ7srbl0JuJ9c8AytOgI4buRk/OlWfmJRjG9FJQhcnvGa6U6rWmX3aWDvHOlL3opLwU0VZJ
BjsP8wYXath2Bx07ZYENnc6w3NFx9F4S0g+6pqaY1pFU3gWUwggVbz/mmqCa0BkB1FtTgHz+GaSa
e4JBvWhuhsVOSd6FUWQh/eRR8mdIRetHZAvNeR6tmg3f1CRLEYxoupfYdblm6aKoFWq3Nekae2mn
XEoOJtglq84bydbMmwRLONqdWu5WmzG8qQl7p1dXsigZkVPx0IF20OAQXTNht+oRbm69CHPXFLH4
CKW4kwv7q/jcd0P422sf8YhGhZfpOa2br1xYak8R4+qs1MZHEeih8azk8EhyD/SKWVFoHrl4IN4G
sK1k2kLlxWrfAGpX2PybG3DRh66BC+w7PF9ysC2ewllXlY53ooZuV1jAHnowKbM86Na4OC2LI5Fy
iVDUVa7wA7f9+7PSpYL1jeYwAU/GiWQ8wHKU1aXN/Jgnq2sglUYUebOeV2QZ19OIjfzag0WgLcu2
kgcuXq2iASoTddWqXo17E0GYcfRyEoakjJIjf/zBIXda6HH28j8hxnwy9IYCoppMDcYesp4qvara
LxL1rbeQEx08x2sViDSy1s9nZNCQgP4M5pY4QFEeaZpe2Vzemy5Es8es3N9CxLYvQtjzyznwDd6n
Ay+u8V9Z2Ih6GWYhexMz3lDlllIlR190t7jwc9sH6KRlut+pJHOspmNQ36YMGGGTDPEkyRSfkg62
BuZ/Afn+6rzb4KB3ElauDxoCFHTmRR+/F0H0cuProujcCFhHb8gcvj2DLjIbO5dE1rzceGCdcaN9
PqKBeqp8oF84C9uz0YEALO1Siw0gV0VSwpyr7Bm23EQyKmIHSGYXTTftfuyZPILfrrLDDMNGIYq8
pGms9P4M5vsM3Qc7XK9EnLSDp6XABuA9yMdoi72j35GwmoRP8U/W7sdbHTe8CM662RV4uK7Pfpnj
D5dfIQ6yXG8OtYb6xP4jwH2xo5dXLAklTLnTy0scxshFlYJ37Inmr8+En+vxEhQHFbzPQ/SFdbKP
kbKd0uI45nsBCWqtZuRHCKMPIttlKoENfZPUDwKTTAZR1zFKdhmZa1fI8flrQ+OrqjBOmaQgdVux
W2psgFANLPCkQBsjDLAmwXPhdljQPxHkf53+g+3GfIJvhISPWqcXa3FJqC0XIDcbIdNdiwRDc7rd
5p83u7PxYYoIEvUZ+zLpidxiaP12qEjtZ3eP+RKD7rgffoJKBGYn+noiK5RV8Q+E3RswyGNQb+Uz
6+OO7t/bo63/Uu7vbJVF4tX6/eSIEADd3wN4yD9YyWOmhPzDukdDrWGsYxw5zvO5wrWRbVxCnEO6
9Bg1XkQqyaCnO8UROW8nKxoYzVjzOnaEfEB8A3RTDsV4+kckGeQle3Y0wov9In7uuVg9mPnRTozL
lq+XTFzCW0llGl71BDsWMS0bfcX+Sy+fmqqtCunlFsr/FVLUDaC/pYsv6PfshfVii81t2png4+fp
OaJG+R4Ox6tYNe/VoosTht9GTtRzIXP/gakr5E2RGAUbMZ2qmDiPVtRH2AF5Gs9567LVBzcD92vz
JouLtkLKfftPhjAzxoTcnvYj/aO4ZiDOCzEkHOeEM5YmKj2pdvkjmWK2DZGYBvbiRjpjouyMKV0x
hLHyypXXZLMSzPGVGGko6izFBf/Un0SAyFuMOu06V8tmI757Aw5fgWg2RVd6LDIoasOlPdC6XXaG
guVnTJarEhNKwZBJ2ir5U8gaTIlqiORncuohkPbZS0Vvgbx1mNsQDAAzZ4fenaKXN5Bvk6ifsxtA
nDKk6TaYxRZzaX8xRSY8W/p6Z3Jdv0erRdksW1TKZnA37dkAfzBYmQ8uPa3EethOhZUWUQocoMni
6HnDrj2CBnyHQwvQMnawauWAFHrMPYlt3nS+cHZp8Sj57WTWP1uOdbVW6pziRCY7lx926ZLvqH39
GxH9rTvt7fYg1Y8H6pvegGD2T5c5VcTvKoQSgeyLvBuB1o+SoUvrnLunwq3HbzGAubJVa7/EsUHb
xhT4elixp7wVowht1yeD4JV3r6nG9tC8N10NPo8xgwuYFfWJdCo+hElO2FUnrX+GGo33KxbZTkQw
39JNatHnqxhinyScCfOTpSIarnYRvmXJGyjsv2oHDvfGrRkonksVoksFaY3sE0/ZNNMn55O+gzMx
3IXsL6eK6pXVNMv+maLhjWAjNesKd4Achd/2EM/EOfxfZyqWSbmS3C1I2vyX1ch9cIlyd7pejNL5
H7d1dCdqx4cfQf9QZwOtVfo1PXUZVW+NK+PC5ztsS0DADeY2fo9KZ2T2+sb+ugpCn1SXKTLF2c4F
t36J1Co0fS9s2hEh3Lehh/ePD/F+1qy1Xj2g1dy+G90cw7jq1u6y9AJrI3q8K6h21KLS19wSPqmz
vlvv86J0k/ZEt3inFASUwrBsno7vjxoKtP8SFPjHaJ42Qt73rYyHvSj4ux5BBx0wW0+gm+hJJkdu
h5u/SIa4klYwu4774bR1KVGlBzWYR6T2cdcMZBoq6Cayd3RBnrH4DjF2FOtlfup6zPKBeCxu4cFa
VpJ3uZ62J3l/P/jwYi61f+ZFLjoMDvf1ylvOZ1SlcU1hvGJFBcbwBSwRgtrni0jd6lRxaUlHzEof
d7T5Ftwt6FLPqmTfN0k80cRGIu3f90upRAfVN6e19OKsdxwJd7NaG+R3lyW2ys30CYaAgX1BRUZr
9lGc0UNCd0X2Zl8fcshKC9RxJDAGCW0Zasw85HZpbhMxrq2wG1JJE7VkXhO31mCLsiGQeLGfL98m
U8tjxFiDylP5Qqpq+MLsuq/4nPYvfsMcU10+MafKOFvsq4sGXxgtE2iXysnXPxJZ/KirV3UGHquO
I5w1Ljqtrrq5gE0z2GyCXwiQ7qlG+Oqk4y46Y/7ojybQGnnz9qsiBrI65xsY3imqB3CAxCbpoyof
96Mo3J6D8rX3+YPfux/up+p/hfrARBisFSf2+86QDs3o/XWzTcj00/QTjNsQYMroAquvaWiZfFWz
bUVssJavl6UyfvEn4O5xnFzbOMaYh2aLeMfQIsBus0b4uzlLATlDszpi4f8jHAqaJRkMRxlDw7Sy
Uv7dEz/BxF57B7xDQ++5X1x+PXqCFeiTSdtVXs57BrWeMKgXGtO18lCG/O4XY2xsaaAZ4ZS113VK
Lzk3KoLVji/TAzcXG7Mazr9pcyZ/c5uuKHMcmNrnPlzX+6mdiOV97LRkiruBQlp2n0o5opFaXi5b
GzH4liOH3layNtkEOOYrZPoDXXcAAWvgjTGAILuLguIC+yH45nSoc/84CddgPjkrxwJ/hsxNaFAI
kvp+FTPT2zmsTdWA+/e7Wy4xNbeVgap527LdFNlyN2onmAApu6tnjQASUKeV93ec5tPsnosHbtUD
pUwyNb++08UkOZ3mPU95ePkwnz1FXr5H4ExcjsyeKTg9AsqrKtEXK5S0YZrouMwh2R2NLS9N8oC8
6E7MuZmCmBDrMi3G5+uW1LxPAFxjIPFMraZ07m4KTXnIiNakwR5GGUxRPR15cl/WUTOtYrzqtmYC
qpZEpvGB/1XAxw0Tqy+Ekd+hL4cutvOFkLiRHhBnyAUZnoOO+4pOY083yudIkI90VdUw0lM3EfIK
n4dDk5D0FJEikse/GTn4tqzIYztTb2uZErpLZAWgorjgXuwrLcDRzK44+P/VrCL8dLpXT23qz4f3
nA4Kjbm9Bkq60SJViiyKSaHjw3D0keUarRXvH3MSZCI8vWf56Zi6d/OLsdJTH1geh1nnUUp5P8p/
XVciEtmOdnzp1/DJ30Go3kFjZkHULa1yMz1nenEZJSZpkc0W95jg2E56iukyl5Y3mUbDLgCOlp95
eeMpFpN9FrPSR45aBqpo5SAdZEL9bn4kKFReXoQzHe/TTHPY/eFqbZX6leMBC57Vw2UMaG+w/cL5
7U9Y0JH2sQO72Y776y9qd/C4mKSKDXAJM+5bwYLxq6bFyt6842+LZJsljvLpdb3r6x9nlqXYN+K+
8wNBy0NSQRqyAd06ZcBJ2f62AU80EXaqYI69xV5f0OFgLuP/j53uMqt6lyCboVBV4Es7G+zbtr+a
C251kPU+Vb49+FnkcIennnyneJ7tdOUFGFpSxBJeWVMBgSjMSprJNuMU/PBLXm+Cnii/IwavrhAS
WxvwsXDOKYjZGPoBJwtyP2QnoK/6zrx9mN93CJbrC9fq7l8oprVfyg9FDWxbYkiJNhPuEiSI9iBe
YU/OuwgaKd5XTXGtWU7KAyRlvbjhjB9Gt2iRIVT1lT35y3KHKgdDx56/21okOyMq5ucPXsqV0vSO
gQmHxoGBoOvN5QnP4NOsHCIWiNTZLN+tE+DIL8E9QQehmUrSTMWQJ00mIFymEqDk4nlxjDbs54OO
KVJKn3bWFT5WN1AfetcCUo8c8mxPrzYAeotRW0MLkrOoPM8AwVkAmb5O9spei2HNIYPe5AHri4Rf
xOqxNZwjychiyX/1geZOIHikoKDOrW/0xL5PMEStULNdBHGrN638A9fKur7u/DqEjZ3z+3qZeC72
a53s0SydO/5arQWoUjMIFVqAv0AMLkwjss6+CTBD+H2tB6LPXRC61O3zMTQazNbQENb8hm082drk
uAaZPek1IK7nxwKCovSTC6WTGrr4xlrdcrVSNkDjmdsL2LMeQuxRSZ70xRCfqdjmqnxt6W2jl47J
uJ1dLaaBAK4kKiOdAq/EwSJjX/2fNbODBuJrR6l4NdyGKZwKjYicVtjKW3muxR4nnhnfm2uQhRdI
KXpkDN68cIWyQR7GrcsCb13IDc8p404+LZjHXv1Wkrr2tr6fs/Rd9S7OHzqq+AZfxJAEbrGz63cS
1jsK3NEcNn2vwibhix7wXTOw2tBOQZ2MjQP6NB84I9zK43ilbGGxqwlMMJ/7zeuVmfmWIb+XtzAr
uLhMcN85x0+ozYHw2ccChFHT2BypOfhTGLPUs9l8dkLIsd5Fgul18IS75S2+DMDUJR0Q/OCDGzDM
wDTRZFI6w4Tp7wkqzNId0GSQ8m/qW2iKfxWd6vd/TrxURdN66SEAo/EB/oyFAacO1M6XIYyUyXpV
TcoBdSQnpPMZfkVaPOz8PtDCbQ+L/aLQz42JImDh334Dsq+vMbdGeMYwMIwUOSmNsF+rx3iIRpEL
dmfehXP2mvQ4Ias02UnaI7IDJrgIULFLEzoVAJBBRRHiHC0zQnsZN1quc3Kx4hmaNA4AeYBFMh/3
CuE/Lws5hKg8al+egI/MLjRUvZoeXp+ypQ/z7VhEPfU9UslNHAiPWnr+fqtCypfk7R1LjdpfB93U
IiZMrlH/+XJ9Uo3Jc40lqaypO3mqFr32LK9F+NyGeb3/k6X5RWlOTLtJU2PnBBAtrLBbv2edxKPM
S0XOidZziY/GFkvPDhOjqkEn3ljv/WmOL7I50Xm5V4fHXBzfJiJVUG6DjpM6WJlhaW+s0vAzELCO
P8p/JU9SR1m8rW2baY6waukp/ggu4SpHuHnvs/Iy1NpNOlgi846VDXTLg1K2enJgaU0eeSYUOVtn
ypBpjVhnNl5/ssTzGCq0N+Z1eXpX0/ezirjJ3+2gNBJ5VZxWZbWibE71vqxs8CdYyFxCZVjDka6g
9YUn7K8mHhQKiCNZLPRiok7fT2zYDBesZsdBq4i9qALlCCgMYiCRedEGjh/YNgMTJsljNb1CPob+
M5KPEBNsGok9x+HfDgEOkKfA4f47L5nioitJKuegk3+OsIatw2uP14wYd+n0idtVz4i3HIjhgyNS
kGWku/WTi4auBICt64hhgS27FsvpaQVG68YJfeIyt6uQ0tg/kxXizDcvKA2VN/PT1jd5AXxDM3Ll
ppBl2V8Lyw79hURXYZpJvJ91Pgf8ug0zsvdoF8Ttj02i9k8oSMKj77dIMWtzCqqidZ5LGT0eA9dX
mnUMcYZmwZztt6Cin3+PgPXuuOz5C/p8IcoyYWmeKOe6uDoixiIKM3BYgecZOjXTIb/e9hYAWyC8
mOZPRX2ha22DDdWQWOhW25i5rGvn4XMO2ZtVxkF7uTOmtIPA9YAEVA+SHp3VCmKP6sIOSNlAUyqa
KC6+MryayAT4sZAvD5iKdT+Rqz2tKjLK8XwVoQnZ3T8MIB/AXh06ZF6kzbNhkB+pfA3QVzDx5Awr
Y7TUFcrSg152xDrC7bK0SPpGwij47qOskP4tLOOAv2GcrQl62m8Obzd9shX1CCH6/doJzBbd2kPm
i1gXRdoxL4YVoM1TDUIZo6JQCiSNamKoHiP/aL/LHMm9sUpbNaKfFGbudBT0ddpH4t/c7jB3b+cc
vCk0JDzIxKj1O75I/E8tzBMiaedKXRrQ9KdVdk4c8EtyicxrxZ5gp/J9RxpSN8tpiDrnU9cDvOKl
EvuIyr0EgmqP++fiNvas9CQHbuAsHCeybAsG0hCy2DuEkFvlne4W/lYr2Le4cxvbuWO0b6hCq5b7
pufMaVLpLTNpPrFJDtCHedo+saXahISTVZ4FOSdc9rT34Gzu5S4XrdW69qZzPUVcfEn2BcyoNors
GKimgUT/96zrEpq2BF5UPSdU4pZftzqn2ii2nmfrVQez9cYMgh0Wqc2RQDalifer4G69NqrElb1R
SZdDmg1qqSgy+Jsh4lkk29Ac0eq/PIjc3HjgT2gVjCb8qYE0zY34MZpmH+T2sVZ86BvVkn6GRdeO
nIMpZxlb4jARSdBcu8HApRsWSCpiQNGO+w/w9s1QrvZiWlsC9XMnR0mXoIkxcnBeCbvrkO2t9c/N
lMBuPmxOSZRdOUJttGs8NOEbGL0ob3I6ty+NnxCIATkAqV/fJS/i+y9Q026seYJ3sOWdi41Kox7R
1XWsJ2I6YV0e0b78UWg6X+ZIm1tjc6i7dyNVVFxEGB5YqwAV+bUGmMjej5GHoz+123Za+HGnTxTw
MaqxTrxc3JnIWM2qpVcPGFDjDsuHfuq2Vcqytupd5b4L6m03Dpc4UhxItYzMS+7b1aol9pAGVlx8
OlVkqiyaOGzM8iITc9NcBZ7SUfVUCZ7mpBNPWtl7MKsmH/A8GBo/aQIr3xs1zz2yjOPWFtawIZUP
RNjx1+sOwugRJN/rv6lv36uqbegARsZ2Q9QY/L0BQp7j95zECbwaJeeNYEuEVFk57yh2mAcARrW3
lz+i4ZhB3dbIqq6bEPCSjy+m48/2JSntdL8D6XUh267itW0TGTprwSi2Ewv7yuEOl4ToSikplPzj
25x6gAhV67tAc7exrpHtMAEGMB+vbwLwz+dp8k11rxz1HAEZ3/1gPuzlY98Q9fd9+gxVqHwAdrTg
GozW4Hv46n/EEzTLOt/mszKaUoqlsdn3dqzc7DMTigEZscSAQGvODTeZ0aeFXOPjsBz641VWkXar
SfRt0acOg3+hmdcuDkPQ2uLaSECU01oJSU1AU0yGx2zmom1o64LwGHPg2gJT0RJ5lgeZ9sgQuaeh
6llgCMYtzszQceLmUEPwXQzxWnCNR1gcSwYrRj+a93YrLSUoq6Ejyn/x9gyhUjp55kVr5RIZzXes
h4gNdqx611OtKDkJ8yzwtOIZrThu0KHaIctBSMpwlEFZjW90MJl5wWtwM8nFDbopPCP8TJv/LNY5
+mUx1EPU5i7ATy8VIRzvAuLuwiOM1dGJA4QKut4xKI2XhCNHVu7/ToyOjoz9dN+6yE4i7UIW+S9M
SPPHgGsDgQ9av16c6KM1q4zm4iGM3P2BmFGAeS5Ofnrm93PGgzfwFquAPZ2gmsGnGW29KH2TC2Aw
Lb2N1MH7tzTAE+ZFLy224dELVNoJN4Na+E3TPJdwF4EoVgM/kEn6iPw+l5GmGCbySM5CSCkg1Vgl
CrOBnZ1r0xlJHyRomIer/s4xGzQ+XAUe5DN/QPT0AoI70Lt0s1qiPDB6lsltCSWsWzw64CmSLW/A
iITOzGwMd5zV/pb3iVHdhOqZ96isLEDinwa3yvxG5mFyukZED0r9Oshe6wb3OQkWAfZO07h/S3rT
AnYmgjnxpay3uYSY+GcLaps1WSqrSE4BL2ol0JFjDtQQ635LQ08qj1gYZa/JXjWvwab/7GR/s6NQ
RTIrecajBif27x0KotXxtcHGsH3vcsjtiX4Bsrk3ghHHdHTTDWEWV9B2Q2im6xelxnBDw2P/sUqH
O45PulUGSoq2LE10jVwbdm6gQlQwliignU0r+y8zFp/UdWm4uZJxuHcTtK1tanFn7ehntlurUBuk
fvxS6qUinJugc+AoKBmU9MU9tVoEscztqVvce947RZNCO0lxPdWAn2a7UlXzSzGQVVJdB/rD1Uxs
TAIcPVzohjlAv+TSNV701qbZgG3GX4ZF8pjEgNMDSH4hFJnsxNoPBhfIwt8z8HJ4UmK6NzYGEd8K
DYzRBG9gg/Hg7QNjllJVwU+kI7TqOoBe/VrqXReUgbt4tJbggh85+tbq4aq150KCI1p+oSq3QFsO
9z7BrmOHGqlTz9yU3e+RjWp8YD8xTkJDCoqP2iylsHTuTrNjsY3C7Wa+YNQa5ofBeC5k+5D7wy+X
7y8mZ6AebYR6IlG0E+3yByqYaVDzeY+P8hAy/LPZJFTYXng2ztJvPuQsiE0Prk3g2Y3wdSpy3yll
ZyExIdSjDm/hUNe0AmzMPxu8xT+u8YiTyscFQWaOb1d7q6XoPR2u3fdhXt9AnysSYxRgkW8UtXdy
ftme1z2AmOyVl0EF2ttFoM6+eCw6Tvo32041ho6JT0qpZ0UoaefxR1ascB4Rkor+F6W2zKlazMxy
tBeew7z/SJ35hkRz96mganNDviXTsw2M9ZLlRlBNSLUbnPE7IEC6HMn4mwSYljwHIeRrQaGrb/Qz
8ZaauqfnixseMIgaMHnqiv/qEbR0NJdnj99iqha66VvIrKZylvqOfGnEsFfWPzENyZ0KEIxQ2xwV
4m/oJ8qO+e8ESeaCXmg9tuetoxdTxpjsP2XUcwq/L4/0wfSBTurWl1ieKnjiycTqWBabr98BymPi
GqZ2xUj/oQOMGMvrPFXHnuMaCiYWMBZv0uslQ5cFj7Mz7PZBt4n4pqGSR6qJMu96vkXzrTubl+p3
MofZnwQPbxBgku/fZXiOpJP5/RIew3JwVyChwzTdLqRjDuJqWbisXE0jlfPcsUhp7KwiVlMaldPY
s6/ROWANsOJCuvE+9nj9AyD4CNWMKc1eRhEa6DahrvAuiw9fiz5CKpNNtTOh9CpnxKZuqvl4drsj
QJvZeIuyUUFuoUkc6+EvgTK2XnLcxk7X3UzbD0fZ87J8lLCcUZuDm+rkUCUdt1HWrsJpvjIac3nc
PnaJIz/SP4wF4neEZPnal1CsVF8CjCgYrjeWsyaSGOgNjHgEtjBlkIzrJfj/wG4UaAs5dLK7Azs5
6GcJKtdZXhwNNR7HHJ283XTIAwxMwP1cQpB8rLkU46sdCiDYv+UkBFZzf5oofiKfvsagw9WMeX9j
iEjWflk0U5UoZ23u5mfz0SP1XPGju+6ywsiLPEdNhpunAE45UtNetg/l5jc2rTqHTBd7sKr1m3RX
RKFUGENIjUGZFqFNAcsdPoQk4cr6NWTlcMc2Pyi3Nb5Ue38DHFev5uGunG6VGzPBx/IcjGE0tK0g
LMqxn5mWxUD2GtiwKgpq6zPG2G66v6l5BqJkU08/b9I8bD903zEsgXkjsj+rLBTxpA2U9hkUa1kD
qhR0HhTarz6KqJiRQnZO0wFbFwGiR1polNsMrIrrqkd+H0ER19mpp/GETU0y0GiX4ZS9ykBP0n+2
f1Bcrc2UGE4DZ1Hw0KHCBAkWurmz4+gR0Y9yNTw8SZ1B3cFhi4sXZXht5Vr6zmqsL51Jg08Km8kX
49qQJ1mmj9znPc24mrqIJ9cK+XiRujkOWq3+c9kpAN1wWNdhDOeB5lkaMM8SS8RwIsQCVTk1EzSL
vpELm+44FWGPwyAufly2USSzJdbg7gByG17SH+bZMA1bpVxKTG+dh9lgQypSF99duuDT6TjDjDyE
CfeQnwXQgeTk8ihR9lcyeJTqzaPwNmaQorjcavc0f1g0dfoREf6NhVDA2sBE8zeHrieTwcGE0hsY
t//kKPTGbfAqk67m/Mfr+0lXVYmNkGgmvIHAKymoy8TgNZS41xfQCXtXp66+/z/4ItUfpb/m1oYS
NL7ncWlMJk7jAP5JhHmPYVVVBoFgELum00sWzDX11Gd9B43PUiY6YsO/xDN46al5OlwfBQZLcPMo
aalk4gwvX2iTYZX33jVVHJYfHVjJ3+fRWC/EIoxoI+zFLHG+lnPBum5JYPqbcj7hxvZfW1gWi/XV
STkGx7SwwkWfKhmuwC7Iu6W+GsmI7LRCPxgAuL5ysP8xYwHfA8cPyOI5gYGX4ybs8RyrFgLBcvdP
R7zLhoDItE5JoXNmyfM4j67e+Qn8zBPfdc5/ph6rxFgDeQltuzm1Ld9xWGQgurMbVRAEGr70n8I+
IiMVhYgDkc14vncHcqqjfEjzERmmLXu7GarY9mRk0WlpqCt8N+MhTYb/6wIvewIBh9hP+xMgOKt5
WOyxnsyXfnbm2ynGpkmFrh3IxoJ1d0WyAHXid7tOaXcl43IeiTPzCa6avTbxGowvnPPeYcDV6iDB
ZNvV+y3i0KwJqoqAxGe6cIS5z/F+nTcoOjrqjrG1DVPVGdiN8MmaDL+Kr3sfCUduZg/S4Ep8PUGL
4+6A6wRG1AqfspZLdd+hKksNzN9yZqpFrhStb7nnRFuzGHvWPMo5EzArHTgvN9G5+MtUkDLZW1io
vfHP9JbQYaqXolUT0XZff/BeO1gA2g4sHBKGYd5DMnPEdHrrBfmEA86psGt5WfVrknF6Igr6bg4C
7tkt2BjljGbSfDskom04QyRIwViuv52NZOWUa3qSW/HlltpQinLAy7EOXEbq+musP0S6k/0MbEA3
iklh2Ie10WxGjvAScvFkgch0Pjy07xLXWOcmXJ6o0gKikPDehd2EqeX/hwMtpvkpso0rtqO/wMCf
HGidwMxB4VbLu8qIbvo+jOe5yszB1KifkzP8FSaw0NbHIm4If1mU4UBTRjVtwsIWaqKwONMCNcL4
wWTbZmcYesr6ja6Kv/HlQE0OhtKbsuBs9dlbl82kYWHSi0wwQCwEDpd6ghVIb+gLsYoDgZiTQyCq
U415BMG7J2GTbQf1Ad+4FjrfvMdQct0Y6ZqWw2brZM7jEJOwH8WpzRcW6wqgjwbWHi6DhBSvw7pI
jMs0wnWu80obeswSYicAdrCG2/wafujUkhiqHkvkfNzpYbtB7rlJ2wTSwMZnhDj0Z3Vmh4v++QwW
nQtkkIYCgXBXr/oSuNAU1ojnpHqNyNTasoUpvsY6qBztmVnEtRidbBB4+bf5l5hn1oZG7q4ut4Eu
Ib/x9ktdEQ4aY+ozBOIUhp2nL7yC8aCCPeXRzhKRXnpc2tY2vWJ1gwZJB+c7MnpXQzsh0Mf1HPCL
mtGtk15GW5kUfKbC158MmyjspP7hEaG51CNYaIfAhv4hQJ2DWSK5xb9J2Mffs5YC2hBQDYUnzjzW
WpIB1L/cmoBFKUUBR27wSJQiPY4y9wlhtdP+PVIyl61c3iraW7p/KOD//QOjH4GO4eWI9MV1IAlj
ifzSqvyHfghidpn9KmEFSgcTRPWxXXJKkbJPs0nrYWWBmuCEJRNZgz3e394tXBBsT0BR3u2bzhId
D5JuzQn0rDK9IEagRcRoK6rLCd3UD/hgrdqFeqCcWj0So3IJDmcvLhxXiLNYomuZ1sjBdVIFtmXz
YK4neoG/kgWsWRcIrolXBZWyQLIFwq4V2PBaSC8prqcP/soxawTFh23iuu4+hJeZpHD1JoxfvWDj
ATDeuH3PzyVZYwPfgyDgv/9d7lI1npbvCYVGuQLxSxoa84I0Vti9ylFYpeur0eQSSu/qvV8M+BJb
jofyfO+NnilhUMuSHx83uZCpztyL3sFvolkDgYzBvrvwVtE+YO/lFbpBhpdNN1uvsJ0Ezh4X0eiV
WkEuUMj7aFrIfwvWmWIULJDfLZg2a0TULbVouxKZ6PTwdjmq8vjtmotg8tjiWqKVdkB+dNH6d3GZ
+xhk2s70GIJgyISLWE9Sq3f/VjJHG3UKJRaIGS7ptbi2f/o5sPbuaGCE4JoeW7f9/xToY0mgHffL
BXkzO82vIGlyfzXYN9zvkRe8PQEUh+3Tgx/qiPaLlO/qV7kE9Y/cOrZVlECd4ovMRYEhMnMDQFxr
UvJotPHP4qYpbo5R20p9CWl26oqZl2bP7ufsCiLAYkVThQ+esVcIBPeqSMqfreCkEwYtQn5z1uE9
Qq+NbM95d7Pa7yCY7PlTHq7y14G+Iwnx0/jXRpzBGO529RdSOxKZXCxGHkR6vSSqB7AjHavv/Z8C
WHiAiWPYzkYQuoffQGOwSctbpVnOHOFwvnU7vRZ6KPlfaUeAXqqtoqS11M10gqS2sQRcLtqRo/b5
98ufZU3pXLvZ1KEqygk/9dBWBzJIvY3nrI4PkUqFcFOpUDD+9qBOGE4V/iH7EhQplvOCPBWQNTbe
cjjQfSShsgmvCqwHTJaJlLI+3Qllv1qj3qkjegn7sT5dADsjHpW6NHemjVdMOVxMsBqorqdOYb+/
Ms4/qX+IJ6a46BqiXNeOnMrHU1cwrzsKcf/OOKqgMwIEYEz6zhVrryqUzFIi/YLhX1OcIQmEozzZ
H3alo1D2BM5g5XrWfk44uv/wwy7Rfkmq44JcNToq6DI7yWlq6/6vjLFFkh8odNchfEb48yFSdmkx
5O/g4GQmQRx+BnTqIDbnoqd9q+xebNbzKVcHLAa380ZfTPync92oteWpTtmrmM1Kllq5aF751KyM
2rgWm6PutUgFvb9lO7m0PVqBqgiGhi3AD3OoHRgPqdLx9+4ExPjDOTfkRsgNASSiPLnBZlt8+bSx
G3MggOORA2REqwtxw+a54gKwB2uYyXRh8rzw7by4dBxW9A6gMbWqSoidsZzP+VgacVEQi12Hg0r2
khUJAp/mh6hslwjC4IPU8m4C5mZqZcuZ4w7R2rLOT8pdMsP60Nioar4uTMJp2jr6pRR2rGiuYEle
QPCtD8bHjiYBpjFLIyZxZUBfHVT3JduLxYVf5k5qrYMNptwiqi8RZ71D7K8kIFPP7kVNJxXyKdCV
RajyknGjR6Yox0fGLjLpaXyszkIFwyP3qdOrTEWdu6P7/IVDdj862TW7mGBEFkonqgR8P6AJ1j6B
A+27CTJpATzZwXft5ke2AcKCpZvzMdvtNNl3RcuAQWS3pjGmQVF6mYBSCQeXlt+l5VSKK9NF9gwk
6rZ469O1ya5BDIqjeF0Cz5XckfwL9+050f5A2w5GWqSgSfQYbJY82TOe145XVKsvD8L/wjLoqP4Q
FwTF/BE0Fc0FiEybDqh25l9RyD8FjuOH3KDjMoxr/3JCHZLgsAVqWiZOQClFfp+r0CPiM9qOc2vn
IFiwp9ZoTuDe3NZ3odZAMcm/9i+XrrjLK90eUqn00Own+PhM7R3wvn1V10KrT3M4LtM82yvrv2qL
Zy9ph6UWtzqer0PrZjlDtAUKfyd1SXbCE96GLfyxODkAn8ZrW49xQ+LBBTisPAuutuA16DFlFTHI
MVVn45Km83S+fOD59nk7zugvj1EJa2aDFliT2nIOFg5ZtGQ5BjEnjYBz0OSvmPi3putio7K3Eo2m
XH7a+27O2NWymKzMVGUb0kH7d48748vTCvoavNpY2T0LCyVBCpzjXVc7AboK4j/sCUJhkYiP4hhZ
WqnBctz+JIqclwoLl83Y8JN95gTXSVrFCnuCZvAxJZEPPOCPCcrReqH8Pbq2lk04i4O7NqlP0gEm
hSC7we+03W8EpXR1A1W1PQf45Dw/t9PQQ7fhdbRwZPNK3EBH7YH1lSu2WNEHmudVis4ZQ3yW+M1e
gR9CGFMs0+rAdma/aGWLtIJMaqgk/KKc2SxmE62EtDDJJ8aCbq5hlx06n3I5om/0sPyRxVUV4h78
FcHoScSOfUeVoh/EYcAQ2s7tGxOw/ZvDYFa8IMCXhS1jMdeF+5i5f1giyqNSNIqaDIr95MhjRjfy
m9G+0wTMogWM2C2PZM7kzSKkU1FgZ4LUJVVA2tB4psMq2iFwKgn07XqufE3bzvAAI3Is7UVFUa6I
QzRy8rGPVSeTW147hNC61RNA4DMPhGQM2tEiTPYHMlZ00JQqqW0lHyRntmQFli0hU7YP1oAlLz0v
0eRhiVAJA3TqsuPAOwZd4jL5j5Zr0AqHauFZtRPNHy0S8YK+rotw3EejQDdeKV+ht97dgCAZ8ySn
hDDPQt1Ix2RUXFBF2hWz4fcXH8MmF5my3zhROOj4JZIHIaO/VxqLYjyM44DsvMfuDavex9djz23I
jGwQfU+CvKhPPXpmuvfLLe9dr6nq43GRwvpclmWq5CEXiM2bJpiIaJDlxbqHezWwosVUfERQnFRA
uKzhuaxOCS14vGA+SCIXFXrJ+1pxjBZQmdFVhroTT9Hzohm/XqHrsxLM5Xyt3cSpYxpBsjNlEzs/
L/JrRMg0+RS604I+qGHwnGnNKmta6Sol5WiqSW8sJTQEwDVPy92FFhLd8naa5wI8QnIEgUZNloXS
OPwi7/3CzL1RvUaweRcHY6uP0UYKBttMAY2EGMca9EME64b/Q0BK9duWgSQHy1VWhQec+7wnzW3/
pU6YrKSDzVtH0L2jn0A7/EsnkgKqtdceenokbNHS2npE22HP7OtX483hXYYGrDKyFDHBCU/n9jhF
ZpLSVUnxKLJtoYQt6EG75mQl2W8lf135mumQHJGmvAsd7zS7qYk0ImTfoJ4E1v0epAih+KkERI77
FTORlilkT49LKlV/OqsbKvrne2NlNXrAy1s0l4KxX9IYEiGVAr4HJM7/E5M1oWF8yJoqaLs630eU
3lSb+2IKCbNzuSS8jVn9u2zuDs3EntnVNtTDhZa3ov60B/QQvkWIcFz1/le/4DbIGC++0rJRp2E+
urNUDPGGcGcFun5FcseAgV68SmsHh1nuhm/LtZlA28wf/324sZXVSQocyl2YqVqU8x6O9eAiBPBP
NPUj8vz5saLqvdRbYtC7FsRdz+jCs6bHrO9vA6YNLM7JLRszX9bn5poe7pTSNkmM6fotnFoCFKAz
WL5bqtIZc6xoz9L+xd8ZR4DUMt1gLCwBv91qbLOZTjpCoxLwWp8kHKaANU7V+AZpZUjSuVfGCU7h
5DiLThZanOU7oIB+4qPabmqIUyNi6uMuQm2DkQ+SiedDR2InG0+Z8QPgoVc4WQKg9XZLnxoVCg8D
ii8Hx/m90SM4TbTBFZIGXIk+pz4bQgJh5ArGzZUeOwYy0YcgBaYoTGbjUHIgqNncVCEsoY558PPI
ohzzQF7h5zhPCB93/OhFdXN0f+hZC0DyvPb8Us/wLzy9VF5PFKdb04oCN9NIXIg9qPB0as0WQaqs
Wl+JQi8T39yFNmJ4/G4Iaa0E7PBzlnGJeg38MPl2CENntB0NpGHYFgMwRIt6BJ+YuslllArbEASH
3/VwvgplFJixdbEJy6INGNG5KhvYAZTjz4CGcHzBAqMFdWY+dtW+DxHoS45SxgEyxlf65zL9DTFA
zj9HExLgVDD0wJ8v82HpkCC8CuSYJMEKoKg1DGePHVzKWJurx4O886ImkW9sjQFMnf1oHQ1i6/zs
K1fibpLBnNTQ93r7KESSyCwS0KRem6/AmJjBAxB71A37BzEjY8so/rKVMCAS1YOhzb8IroIIPSr0
DAcoeVSHj899msYB5fWfsnzK79T7egubJQ015+Vug4Q0Ybxd3e38jT7UfyPJ9/0BZEUH0sAMmzpC
S2nJVxW3Sgeb8OqY2qm6Ipf+MZoCAG9lafTciwN+YW/Sxj7Wsa0G0Ytgv7BSEZc+LGAABn6VxvJO
rdY/MpaArFZ6En8F+j6qksbwT9dp9g27KmQ7c4sP72LIpwQbWy5s1LpYVuqyc+FUuSUV3zzCDIVj
XTbciDBtuXSvxjTCyICrhc9ViSyUTeVk6QoPYxFCHvxD1Jz7LPiPuDcbW900mgodkiu5IoW3JAae
khG84sFDRrDWa2WX04xBQfMSdIRBEVW3RNgz8A+YKZ7v5fiMxhIIrjfz6EvlzFVydup2y4zXNbK0
IdIB90h5Tpgl5PkIPOEzZ400MDvCpk0wf2WpPv76pOdxYz+HXVd+jXFbvV0QJFEr75W+ZYsqGeLe
EhGXjCkcCGwBGgEj+wDBZLuIrSp4aFy8gEmvPEJqYe5iUN8pry3lL98r72gV+grzSx59fPmQu0wW
jNKiVQPQf6/55BqGdjkvXgMhI0kWD3D24gw4f9kwbS1adqj+pKswdN98PJitkPtSCEfOspd+ICe7
uk/U3o/3PW4YpSefS2cE+5YquAJqtgC6qToRu76vtNXBmJUBeLxDHjNm+bw1ixf8xTnF9WKKjh9O
3xRa2T4xWhnglLgJwEMrID7cJU8kqSFRyoKGtxiqKiAEpinmBjy+Rp9uismEjXRsZk7pFxtdB975
TMIcavzK4HcxA28sup118HHF4LWMxDxsrCu74jDL6pJoNfdArtG9AA46+ye350dCdh6eVZ/RXkZD
i9rQ10PoH34JJRESWZiFS80DCvJ8XFMRNAedui7DrjhE1VPQdmo98G9olc1Vh8hhsjO22zoO0/od
tB38PQxiXQOVOdLdQ0Q/84AaDqyuvw195QRN5ygwUfnq4HJmlGxBhr9xkjzno+eqGZ/G1T2PItRA
37HewSJJQ/AogBYa0+YbH4yCmhy4USfgyWIppgEEwWgCZ15uxuTPGdRUVs4xOSfJtH2A+7fqUBVM
CdmS8b5qko7rBwZrZTIM3/FqueIDzVa5mikJQX3htMUlhWy4Ffn1WNVcZ5Ym6AXem/feJ7RfRVOs
+2R+dSq/yQFIBl3XuMiwz6A6YViK9HKFO3QawIixVkUxIhwuKPZSau9r1Pgb7rsntojEUt63kGc8
2j0HfYo1U0WEpPvd/x3Pc5j1YG9ZAgMZzdjIsy/UZ/e4NvQ48C/EvgqccepavZYfTPRbvYAJY5IH
YbqR/i9tHS8SRNK70wLiDwtcZ5gbYv6Vm3YjevmKQ6lRKFSYuSgkrJ6KsJI5kdb5jCi26AdPVPYm
HbQsDD5NSxnvOhm6q+1G75hou1uz778e1OqbnNRaIEv8nK0t4v0+TOyL8z0rrfwzr4jV42J5Dctg
XspTrRjbkgG4qL8aMH2zZOoVMMQzW2ToXEwbqdZr5kj0EioW+fa3S0YJBA22AvcO4jDRv9VVLTvi
HXIHMZWpP5vtLz0+kmUHX2/0r4Wp3UXealF0tZAwkK4og0LDeAQEaLoccy+SqY7AlJzDZmHVp5CZ
owj+AjIneFAuJJ3Boag8hslpt20ZpTpuC7PyJgqDHdiHP35b4qee/umVIeyRHGHoLGAxkw6aT5tE
PhF30I37InILeQRzbYm/6FM9/7NgZhOV6tUAP2Tf8Uh/N+j4wQAH45qqWfGmpciOyY+EwT9VPasO
NPHbazMz4542n+evwrsMl8uRuLVr7QQlyIJ/NSrIiFlyV7oJ60ZnjhLWF4HwmmRUIog4USFjggHq
BlY+WJjG6gjq+XF0aSE+z0X0dMoc5xCtV0iBQYXj7AV4VfQ1wFy53hJQEgNlERIjxzSUG5it/inw
87lC+SpsFr5MiMtqtLSNqR3oMpNwMfFba/32CJVmRKLiTNWpn0fet8z5QVufbSRgsZClGwnPwXhP
w/HGKmTz0vfFcR9fklsF8yarzRMoj5tSXUoI1yJB/5C7xs/sUIwj5FdN1RDvd0ZEGkzkjhUMZtM5
Xr3bhqGAOiO74eGlxnnzcjpM6A56ecHwTLJZWL/6QxxN4IIEm9vacauMyQRPQL1X2LUJvMtvhTor
4EGxHHqjTQliYBbbCjfodRjq9osOGEKSDRd6pxDyxglox23n2+ePRRsqcSzGx/Ra+gSQd2/L5wyd
RFRiQPRzn+vcewZmHiqVRKjNY1vD89g+yVCfEPWLbkDxSFelU/e9AItesswyyVrhUPPfF2j4eUYM
VDh5LiZqJ8O6PBUnKXwsTZWPHNX5IAA0c6AP5gJViDrt7eIAW1c0mTK+u+IPETs8vl0IAnQ8bblZ
iyrfZUNFG+wjIc7aeSFgRrzmTZVPaxjxzVl3cvIRqw827gZmTCGMWdqvJUcrY2K+iedJ/gTY4p41
ncsm0W61vItNXmqipJWYom8MEchCjJaqHWPzW/Aa4fQ1unA8+4XkU5e+EkrRAdwaI5PDxIot6t6q
EC9x9Og8Sn9Mu5DO5qKCJBOE9M97jywGp0J+MAkXQ+Mr2pIHKCFkedY/qmIp03cTQI8tzqFn6dJC
iolP+/IiYV9VrQUr8DinE2w3IvIuBLQt0GFPJ1RQdDPZCHZ8egfYASCnOewMdmDuCYbxV4keAHhm
xRwhprLW1a0kZu5OL0g5Pcba/F+ylrwex6qFUXX7h5typwFc/hSDa0mT2Zz4d6HUM7WZ1tIEDovu
rW89WthEAlD5EWWZh0llPm/SfmgXwnOwLkk4LUG6vOys77OBZwwqpKrBHJ1jGQKNx7Nsb7SAIIfV
qWbFmsDmxR5W5T8bm8L5pXukJToDvLYSWwLNs7yeeu3SJgY91rvUrnXupBognDpiojdwgC4ktLEi
ZcZ1ZHvGWwBSt4mWI+eOkABNzifw6hwpqevvBECrE3WPNqjlcihiKjSl7R3oP1girV1eKxzVypHF
/ZpEUBft5Ej7QODtTr9xgtypepFZv1QGdbOl2Bv3ua7FMe5K+Yu0C6oswUdmZ+3XT+gATBrsi65U
dwwQnHSFPZlctdSy/1hGUAxNNg43NjyO0DWplatYxzhFacpiVTkldrEEDqX2OfoEfQ9Q2S5Idfx1
xKyUalRrjrOcpGs+insopuTX44bWilrSmaPDKTA0MlPs9lgzsOU7s9tuKX5xL9i9Tm6FNIHoruKc
KMleT7jMODi4I7EXKrCDI5i5cROuoxHNOnKbpPXbHlaL9O7ougG0dcL2mMni+F5iXqXppIjqW6Xq
LQIK2GBdA07Auil5x+cVZcbRuCmFhYzJt2LKxECUXCV/blaT/HM2WsT8CzYx0I1GjETEqWSI5nV5
ul7aikznJnVoa62ldQFK7sPGc5HbvFS5CGEyvKLVmVvCNiS9sIjwz3Qsp/OQPrI8WAceIcfmTzeo
JEV+1W8BDI/HKJAnszxptZpGtW/SYN52misy6BIzg8KtHXc8odmSf3vMHvKryPZbKw8hA49VmbIy
zBPG1bl8PEzQE2hF8+zuIFp9Ta7Nyi0b9GaWZ8CoCHRZ1HId8VhXQ0rvStsCu4yZBt055S1fK8Tx
ti1VKkUGsgIIL8ds565fZXJZsEpRUhEUaHtu9KK3elVkKTvAhUsAwoAUNCucI7EfTKq3+LB73JJV
QF9+Ps8kFd2jBM1/dsrUlhhn9CHaUlgfOlj6xy2tYowIrW/Mg/zbrOewWvBkERR0zME+WGuBnFFL
oT+Z7PZBhGtQ+G1H8LzeUGpoVaeiSsw/budsdGq572PO8fw7Qfdfu3UGxXXfhmfsOed/ks/AW8Qy
Ao6rNo3jIjsK1YUeG4mF64tRuKg28kO70ErUh6ATDtNO8Ruj8hSiRgLq7nMwCLfZuQaxPMLEKUO1
FAsCOa+QYM7RSI/9GYUTdMiE+b9kBNVlbZXJmZ7fJsgFg0gYnr8khbVl1L0hwhlROUm0ELqMizTs
Y2XOZb5oP/+OgfAS8sO/vBR4QaQDWvaLZuCojIxcQC7QVOlYohJxEconerc7izmB+mym5kQieDo3
K5xCtWXP4J2V1dewq1wojYxZwa6/qB7fKrWV4ZR8LPut53gw3Y8hyoMSRGGQOZi4GSiKpKgVSPdC
HNyB9rVfMXckR3YWIiPXyNYiIrnmMTJn2aCfUrrHGbpdYFsbcw5+I6uLkmzTFHvKVRnWDrbd69JT
Fou1xSHiDMeNyK1WWv0mmCAulh7ZGDXwZkP69JH9CUiJleDeebSn2EYX0wOOBepcRJnk0kbxiUon
9B9h+gMf0CxqY09ek7ygJQsof5m/fcjE0azBcnKDfFu1e9i2OCu3eTToQ5dYUwsE+hRquInpdJCs
2F5uMJqBXFDZ7MbR5Tv+nJG1IKQUS/Oqp5kChXeN6S9BsgSWziCmU2Rpk8kfpXIE3ZiFTGegtNtO
UPWwTu8X/3cs6YFcpNLptKq9ITIOLhOJRuPTHJ1sOAN/yk26gKKDopkQCY3LuO3HLkkD/sQQuZyt
NHE2GSJxoNJdSVUOYW7YfMkMjU3kCEAMJKgU4V6Cxc/J1/mEDfWR+93IKLBNhFUzbuzhJqZwyK69
aMrOGVm/9/u//x60WZ4l2/fDbr49QKBKnEpaVylZvakpScoivMKEQetMcO5EFYyP0+MOFm+WVLfi
TCo6f86e1tu6EhY2Y69FWdYIZ38egPrf/jfR/2A6/M2vlWqRg7y6p3L34Z9+guI0vhI5ENECtOMZ
MlVzW2RRkdVhgV+Aem2s6VY1Jt4JVpl+TlNoAIGBWSi2N9Y7hwBo1a99p5aeqM/nbflXWe7HE18j
GMaUzcR+k4FvT7w2baNyOAOA91fXtq1nweKnaiM2djVKOqyeSmIDgUYJrXbMIW68ffLMOn5vrC6I
vpdUcVtMT/8Y5opIrDEafuLkceKxJFjv/iAKDc8cfTMZklTX552Q7ry/c5St4hf8RNDBX2wsXplX
Dz2kkIs73eLPC7MCRbnSOwSD5I5k9Wmv//w+n01eryt7qCX6G4/5UpvBGOTWUongGIR9YQIZnwkj
GW5no9h5RRsQVrcXduq/XmEj9a2BmgCiN/PTOgl58ejBFsekRO9vQwO/SUo4iZKC0XvnLoiBSDOG
rIcC8w5A+vwgchp5RrghSILnecmDE+R/tOs3e6jewIq5crLrPKMf7udFM+iGO9NCL4AnQC5yXvpB
1SSa+IbzXaGzKxvKZ5eTJ1aDeJfIDjWNHMop1a+F674MXWpSvWZRxwvgIME6BEgIHWCRoWqMH3ua
7ZjVoCGR/F42RIPOjNV6uZJve4sN/UmGRmo5zyjpKJAk66jFrPXZ5eEV4Szm2sx/fJ4HBWx2OBUO
b1J2q/uQuCbpLhOyXTdHR8LF4Yz7eRPfyaMpEkEIlvJ+KX4B0QSdGDsPl8y1pYB94lDBaN9v5yiP
dhpjTviu1xbFSoenAcSKX3aImxwRw66g9CtN5g4jI3cLN22PgHlHoxumS8EX1nU3tpcAtJxZ1vqg
mtmRaHCKcEBXFvELswMn9ZoipAc8Qmy261i8QXdljUzXvYxWLFfVJH1ZVdyBkhLR5B0SO5vaL9h+
5CkvOaMHwnQTjkx7qDURqoA3OhmYuYrE/UT6PiuTe10tnaDIJ4kPBBGj5s8XaDIBx0++3qo3iHkw
lo5kQaFAhAa6Vz6XiEKYH8D9qxobSBrPPPInFflnG5aWpBhjXsqJfR3tvAUAPviAAEG16tN8PD8s
kIbDkgK7bS+XdztCoYKkK9c8Li8QYzqUUsWVCO+HEGvxdOLgf0/OlpKKJS1nIkskQWNjnb9zqPMe
dlBxLe5QDvAn1qHwDiAV9cuUp7D6dMvFRP1XbjO+KkqjLNqWodlicWnd0+ldWA8X1KlGMgItftZ4
kp1lk/BMQ3fYDfskUeLAC6RFX+uX4F/8qOTq3RWccyq057fumo2g4YsCgBfZFAwHY+3nipTvGtMC
DEnjdBUsbFt0MZgAke+3Nh8mFKWZQzS1cTNuhPr5YSg65GCvqwByRQVJZ0ky7j5c56h1N8d2cCT9
tPmPuZrB1kvU310pifNEpa37XUqBtl0GzHDMa9MOeK9efSdCslQ07LK9Tq8Zjdyu4fonV9MlYB14
mLnx+0LH84QK7nGFnSrard3II9IxBad/pM8x8jnyovjj6fqJj9o1/MrkQmCPPlJk9IxtHmHYHp3j
sD7mxOKUPhM2DYrLUvS7TJpH4lsOAvlK9EAig6uyb91+1P1l7LkTZF2+njOyZOG1m7XbvLMumf+W
gO+VQf0ImhUv21mMPJcC61DIQfaphAa5k9zdLJ350vIdTOWozlZA1+E3tpkvUSDhlboGEK90M94Q
5OQ/rjrnQhmtZFklxzN74wNa0EFcRhcF32RrwbdjCCv9NW1ZWF7A7X5xNzRKWn7avA6xHummN9Bi
8Mg6gRI8wp0KBkYz41vk9lTbcvwoKQrFw6x08qkHQCy7gTY+FY0WoKEp1NFa0sfmVtzMp7BgMZfi
4DsLd/WeDKpbePvjZXdTE/Ezq9O5kCL9bkRkG1dYEj3JZQBBZLhAY6qDGaUt++oJYczjZjLvdLX9
RfjwVqH64wBIaBLadJzNA1IDpuMRmtHUgDbNk2Kljz9Pr1egL4nJdxMFM5Ik8hWR1WEFgmJfTqpu
ctEquFXSWAoPUX3wJzj6LUgAqOYSyZFco5owg028g4nyy1sCEs1nn21lfxUuHZKtKRRF5jTpY+xw
mXxScXKHBoquRiJ7HFth+AhcRs9gvCno4r+nTSp+ldII57vu1wEBnnffbF8daKABwrvoQNjfcRlC
y7+W0CItzRKojC8ojmJkx4onn/p+nt3acFaoPShCek3c3y7UE6opAZLF99b8/EMBVQSclEqbv5rb
gBiOC4BqqHNcZ6fc8DRMqe+u7hOJJD2Pgu9UaGRy/FsDqZT+DiTmmsbxLqNiYbzZQdRT7Z/D+YSE
MWT6fHUg68U4zhKuses89WHrvQqR/08NUsoTgCWMyET5tRhAsuGSBI0pBBituf5K1LBgz/7vdDHK
H7ZdEW3hGlphnplVXWV5VZfA9E72KKHj24BUUdJKTXrrnqoJcBp0fFPvU96s9J9CC1/VIcZ4m/Tu
920OJhv4Gsa8fNtHHYa4ztWV0AZ96RnB7gISYhFL54r5r1cRbWu9h6yYebE1QkIHvsg2GmkJBT+R
PIrn0hby4BjU+5VQtzwTWryv9gamiwGIEQ9t3RU52fM7wbMXhGgLcKsD2tmZe21RVEiA63wjrMws
zaMwfGn6mrc3US6x1Gj+NajV4XOxlkB/x77sB/OFQ4RTxtgvQerH1dWp5Xbcx/pMBVkv/Bhbghfa
K0/PXfVp2AduXrxR1Y43hp9qZctv/WUkcCYo1vU3GAcdzHBanzp5AOKLxtc8B7JUFWzZFC6Yb28v
aJ/2M7J88eeVzqmKBg8azdAlXd9vZ+KuHhXr67dDknYMxqOc+cw4tC67J1xBuNPm+y74/qmbaYPA
rQbHt4ryi1pFaFekv/6z5gQWEY8mgcyTYC4/cG59L4X38DsVfzJCO2MyX4O6/lqJt+RzGC74k459
yHV6Zo41jGz0rixlJfbend5bjYy7UShAwsgDvJPxswC7LbOgNOpN58bQ7zFMBWWQhGeVwq2ouHKU
XB0pB+yi+blBwg0e1gvtlrYVcC612ncV8NHi7BJEeVXSy33kZS9G3ENb28nSfeT5tlWASL+7aQki
/yugcjEwtlhW45vWgaYwUKVeBYGNnz6P6J3OCiXjdkF5221Lh89kmiNIGXhTkHCjMW5jeLL2/R6V
dOBWrpvPUlETFDI269Ql4BN3DIe2BIDqm9hk4/CHWetMXSyWaipu7V2I0TK8XqVsUluaiRVe6An5
CnZxkw5TYfcJ/p7sqJt11RouAfCyIFyaz1oooW2u7O+P+4fWEE8AfMEQgLpprTPBvXK8v28aOXon
ZVfRD6yIC+vBRkht2H/MAfUSa3mtA5tZyqGbZmws8qg5ELaoqnt8iWwiujBLMFv6sIYJ1KfNyLaN
XBgqgjgLaPOOUJBmMsL50lGaxxYbwBSBD5hRuhgOP/Vpaq6xbdMjxP+Zh8577FiCqwFN+6pLqCh9
LrjMFwK2YiTj8zDxfuQ/3W+grGXfAM+/yEuh1dmGrLKxKZF15Y6hm6qMEjS4sJdJoOJS8IWoM0Rw
rrz54TkyKDZ3tK4lBjw4Byl/CpcPOnsWyN98mzBFIC/VEEAkR2HrzDawOsyS2elyoSHzdVjGWKu4
Vd8ZMJTXeALXlnJWbr/BJvhXN6fEPhLA4wDrrNSrxcBgCBHR0Y4r6XEi0kp/W+tcE+bl0kFzkTfJ
k8QDtHUZjgmjL1tHHQbQGi0KK1sEvn1AOTkSFecC/2/g85D02DGUnhVanwF4NrU5KMsI36rgc5rW
LgcniO6BGUqZAnRd0QbL1yLPo2seISGSXYWwiLG8f8dmjzSackRZAYTYn2YA39DDrcglDt4Kg93C
j2ehWaBgsmlPnDG7WZ7XbNjKwlnlcNCSMGjk6qDvKWCeEQVyFC1tWPdKWBH1arCjjvGZ9SMweEn9
1UQXVoiyugizjXbuuqewNb9hS8ZGqXv40n+hfik950R0EbAWaGu4DF6uBmeb/PQfB1isOGsZUoUr
yFfoUp8K4PdHxTEtmrdOmjiF56s0kPDPz/zqnaUKrptIsAvUswSeZ5A7Wf0sz/4WBt65Ifrveef5
RYKKfmvguVodmIO9BYcYED1crxRK56Ipl9UDpT29F3P7Glk1HPGGYo5xWHvS7oeTG2/vqSkY95qt
hLKwa12ema0dyhUo/TYB4W5m/TIYGUx4qrVm1mpBCNGiSkxKZRxyiOQGO+BqmirzYB0/cfS74QWa
TrvuLiZyqiofC781ctBUE46saLYqy7hJdP/Ic+nW5geZbyUFMS0yV73B88OKZ6CTBQQ+OXH/Ydoo
jeGvPMNZ+TE0ttfSKOk/ycl/rtiZkOYRC36APcZd26Eqct+wACxWNmN9Ndere1D5UHk3Kp2aVwZ6
7cBm2S2ys2bGIJEGCXrAToHUmEtO4eSoTUooC4gJzMGeTmjW8N75zVvCda1Jo4T/8j2Ra0Bs/qzc
paqgkfhI3nLwmgD0vk7pwtf4KEizefnocRBbW+xDMhgK/eBZI7NPp8wsU/BMvcYeQAnb/UvNs5N0
01chE4Y7lTAIhO+AW6K3tLaon243Re1i7UzMZnwN85oefPhCUwNlwE75gvWkwIgiTk+OlLhQ0A1m
pU10ez95sds3p3h80c2fXZs3NDuaOEjoAuzGnrCnJwvDqLxCnM0pRO1nU3CaNl8d5BSZdGagc15Y
+vmiGHAr7WzhFInmKJWRvwk0DGhLIn25umKGUMFCTEJFaG7JbFxUtagPtAORwUxkiaW8U/6hs+Xf
94CA3zB2Eo1UAjLJgQD1DzV08kO911jrO92Qiz4gn5ucWD7tHw42CmDYQqPMBJA7nJifDVTnEPzH
JHIa8EyuN1FHVJ0c/93S9KMa9FdN5HUwA2emejkWYUFQ867e8m/e3ai2O2r2ZriuitB04dUPzTfZ
0pAMjifo3Yhrla9xaD2yf+yAQYImhmwmU/5mtrzBtvRelEMSQWdpR8tU/fyXClYmR8+SNfqMIgm0
ar66rlxjStW0cSZU6M9doHjdtZgDL+3to3/rCzraJ95nQARHflrYZM8Nx8v4RxvVj2ajtb5RSE5/
d2eyujRBT8W6MuKSqZd4MUjhkswlRqslnRWRCqNJgssc6FfHm3MJ8scYGMT5o/3XhPlyoNWrWNzY
CngM7ewU3xeuW478BDSb6lhHCKhahtM8sfc1vl5IjYP1eUX4+MyFXcWG++zx7AsqPFSS7y/+8uiZ
/kHW88UUUNho5KAdjG3Vj446jMA2UhAhNxrdcfbi6HQRYiNbyLHBcTwiB6nqYvJzcE1hVJkMgXIS
qULsK1yf63OpFZs+MX1lCRPjuuYqKI5WwbVBQ2XmdGrd1JWl6oc48TlzKQeM7ohb2gwJvum1/5Sm
0o1hzRFaRLFixmeZizE7wH3aoWdnqkWHPU2lcgnGta0YaHkJayfEQ0cU8E7Gvg+MkIg+cc4GHt+w
RTxiFMNPCeZqj+k5u3dNOJfdcWJ0KHSRCXESmLGfA/QhxZSJStAr9qAsVk114s0EBUfKZmSuBa4U
GM72v8KGnYLTfkXzdIlBj6o+tn3mXUx8MOodWI+zuKSWOD+mXFIbmXpgm7d7rNkoPCsE0lrjPj+M
CFJV9hK/+4GoFT2g9okDoLwJT2FBAbcTDqOS8vLgJeLORXyzvUBzd9UU9ncezUVqVI5ug59cqe5j
YTR8Eyzd+jJIleOUj4c/Q8nndARvKlRmMYpE9UV0y0WdNvaNDmsE1y5ePgaamU56cx7qKFrxGqyU
ssMurVpXRwfwT5kkdYVDfkep5Ntw1Vba+Dc9mfYKlNLN2FEE2xxQOlIMVrY1B9c0Uy5vUyTCZSsj
EJvcXtMo2+01BbARX/pad5SNOOXV5KJe4U236cF7yMB1xq2AptaqaABKhYpSvZMQyJaGM8kVko6I
7sdESAzLZTL85SIrIvs8keLQw4k3b/KWT8cJjErRa+0LktQP/oZ9HvhaFuOAozJuQGIuzns956KL
/vgCbVyBOQaO1eug/4hSF6h3ZdQZZ6OvGmZw/Fv6cL3qZiWSO1Y40bUuw5EGDFRZKl7gXCbj+low
WpPfbNZ6YS8v96iougy/EmbQRlceFBTzSB+LCRaVBWKfgbdL9E9hOxDCNpLh/Q9J7WiPqYHgie35
3cMmxEaYPANAUoAuI65bshsL0rm/AEEPVuX951e5JaiehLK/TPGqpAYnIUapditho9C4nZ4zQGVx
5bjY5X7dn/8Bktp3R7hyghrWtc4VZyC0lUMFD0gV3GspLZ3B2hwz1TzKUpEo8PnthDxQtlgOYl7B
+tvX8ddHWodp8F5xBmjHbaDtDe0QIHUtS1zJ3oKyn1bqqoCSYs0/vqQGyBfGHVq4GuZzgGIdIfq1
vElFrHsFhEBcacxKCmQrpkvei2yEH51c6aLuPIuGBGGCXOSU8xm5mp0XAAXya0k45jxQz4agSftw
DqQ4/xVvVEmmDG2L2xbPFb+hILa9zlGD2he+GwyPQvhvXVJBSqk/woLZrB+h8aKdUQ+nHz6vXrhF
b4GVD28QEH7YeK1wakW+x/wVbpPYPNJ8+LHmrMH3yqGeNFWKKAUjWF0fLynCkj2VMyAEqI2ZM7JT
43dgcHo/coQ/mTK+uwXzARetn//eCc4jdb0ubtkAl4W0oGQGyTfW9auxWYry78HTP2DrVrjfZQDH
BrNpOn4FwXzIvjFZzym10KrYGPFY06Ay5nJiCdV5RKK7V5GGyNSBUgl/pI4K6yj+gvRndK1r7utm
erty6L8iUFb6CAxYYRU65MSrYf7tUmb1+5xG1dKK3yQM3xniLXNsbRqfCEvrl0Bb3kgl8PLj+Hh0
kOABpqOhDkVUF8PbBuRRKdPKtjzeCe2rLuWj96X+zpVRubyLRXbiwuCJkFSux8MK5GWmFwdmcsuV
Ii3FWAbwqJtajbcRdAXzyiTVyTA9o7U2IcqjvkQ67WkGdUXmoMKsPiYEhy8KAv1P+gitZLCseMsg
sQXd93h7wtLiTgN4gPnVu3zwpwk30yarVSmz30H852ady27fXd7uSp0J4YsY+NfLFaLuUATBn+wK
YMEhuddoxelgp68jTTDA56wzfa8SIufwuX0kZO8dNzTse4O6JV7m51ae4oV/KghoDxC0MYTYXSM+
DvxtD81UOynnvbJQ30z1nUfnkqqQdaJVewR7C+pbOUyu9oQYGV5NlaU6XeBe+g0NXFpt8tA/5UBB
OpMuxTJmNAX8iN90/adMp9D6M0rBE/rgE/rqmgmlwB5GT3CITiYuOScAAelgxCZ3x/+DzzdQZZZP
UgBOy+pc+gVX6be58a5aMbuhkqjKJV+nLMNwqZhX1vKBYsAjzsRJr3xHDv7iZgCv94bsCER6x7i2
TwBE8NkevcF/qkriTW57mVaFwQDkRAQDcQBCUAniJFRU7HK9jblPV0QGit3xdCGaUCfP/yIsJyhm
aF1H9eY9dENBwfoc1Y2v9CieHkBo8GWxQ235ep039sLRM+oXeQQY/RNy+XGShEDIOUWTJXu+3Ig6
zA9AiLIKmOJ2BPrSOR9OI5cReOKJHHxMvrHiWNcNipAlz2MZ6wU4VrKKkCTM2yCDLnTTC7ti4xe+
kWFa3XcONyvzD9Sdfn2ICYi8/NbjE0h4vn0WX2KkTGdetyYb1vpGyBI77PB9DHmfDWAZi5GK+pNL
PGqCnxpfWK/iOZIbkMhrM3R/KpPrhO9hAql+HMtnY5tIJP8IUqisduXF4GBcUsFyF37lApbkPIks
VsXiAbslfwSn01ybfKPJHOtkvkT3Xe+YdRxl1KnIzXUwpSXJ898X90kUTUZ8vzFeFeVgb/a60DYz
MH8O0zC6zUbn4Zb8FHgBhPsNV5iFLlLGA31BpQLNOj01Ln/KKsqIgfddPdaJFPz4FgCdH0z4PcZn
BYMOL090il8DsZ1jJAFZ7MuutAzU4N5hDcpwuT6SFUbE9ivYaj2qX9F9AbCJnfGVYJ7ZAsEiZpts
1EBuz6x/SMi4jctm4BnO2HWYzUI8BWlJJt5AwFlzng1OmVYgIu7deZHyAQ4kyEqE5Jvcnhl6AYnt
BmkVz33x0sdPHQLo7mjDVNOXS7QJJrkDR8nWzqlYYyeOwhyswoKslTNhQjTWK31l+JczbihoqQid
GDP7mZKhQLa/73BmZ14hojxMzL47jqV2eb8uwFgmRgj8hj6EpaTZjbcvDBAJTjQMGllesf9NM467
iLtqaIc/zbVP5lUhtuWE4lpyeVJSnAHpZ0BzVIUmu+yKfdmjZ6SD0EZX2bBw83exHnn6OABTb90I
zG4XGvFWZV8aXmnjLeAhZxqdZRIBXm+ytHWGi8S7pqr1vSl74zE2S7Khz41req6e2USflQRuIRep
nPd4p9kcpESDbnGYAQAt1/OX5uGeak53Ly0qo8c5mV6AHhHuAy61KUo0ZDn89cIubls8h+0zEjNA
x9Hxyiqo0QY1UlYepidHPiXWyJMLWqSITgRB55XF+c/hi3QLUGiSS/atiXa97Q7A5cVYhGPTOvlN
tnkNVpijVAM4PCr6H58t9PMJuvgYJbZEuQk54zhQ53VELeE5qUFHzgzox8qba0iamHNf9mB7bHjo
Nymxvn3302K7B1g71Q2jZ9gbdqNpoUI0eN/DfMoNYS3HhWKCeKXId35RWhWdBWNgNln6sqbQwtIF
7nsYhSpGG6pilyGWvNUp1TQ1x1Z5S0gblIrlybrbvzja9330XnlJK2NjOr2FoaKakCIK88Ui8e7K
Z2CGFjfYJ0QwJpjhkPAGuMMD7cD+ZQY0FGfvsO8FCJcdtbsfEGTVP8Byi+16cU1MrlIfZtsGXFpd
uztK+a6G3Mx9pr9mzhg3VFx5GaRdgU0flmjCkDJ6eTWrOlZv2XLMKZQ2C+uOxHqCTpjviZp//Np4
9/IdmSehUsMBYdQ5sP+kk1H6VCCFvYEB2zEXJ/w7W8iG9rF08nGqpbXLQ5w0hjOs68ZAYGr3tesh
1FGOzZasxiSONlHr5uGtAD6nOa5Bd2bdQ3vked594HAaTnkwCV7Lt/eF5OjEf5TdxveSHQJ5/nTn
LVt90CIR3BgZJkJm28zT1Lf8Q8lY1wcry8vjO4F2F4VvvY+9KBIZTQjGB4/yLMo9WOP0A3NKASnI
nylLYTQQ/rf8guNWEjshndB3opgeuFE4dVoe/kGxE93GcHgNXRVt5o15pHL+B0jukxFkqElfrlIY
IV4a1jID/4Sjyr3K/zTGnYUdjB/Uwww89jjgXc3UDmNM6PLUyoVf8epNGOvrUF72vNdPnh49ZE20
8TvaJIpTDbJ27NQw0r6OvAPt8v7S3Pkrq1/kuy35QzTV8T2QDOWpVXHGqnB33Otm7qgtBHavU0Rf
fWqG/fl80L0v3Nt4h/SEB/2rDykNcJ1Wnja9H0QEZs1mJ3jvKAvQs080VJhQq+56CnnBLtviUXVg
ST6Mow5hSmPhur9pqI4TSafu0+XkvqoVt5wwbxup/8jYq6BFSW0mS37KdqzMtr+xPtr0cHfDrdoh
E5usgJI/4qcxH2O35XxikjPfAoLzFuDdyZHU7P4WpQrtfT9jvg5/mdYJjoBckkIxBI2EQekRIXkL
NXK2drrdvXZWUgP9qZ/lLjBWA9ZJdagFBJgdxC2DAfUvtfTIMSlZHpNq+ITe2N36pOe2xG4kr2h+
U56GkCP/Yo+ku4QIJIiies05T6BkBhnkAe67uAWlFK9T+BRerJWFFD+RbQNMaRl+tJXQCjMvY0FO
Wzu68tEWMvYakxhQSQMUw72xL4EYZtlbGYCrhkjueh55GUWsHqs1W+TsMeddUe0s+J0VjYjQJ9cZ
tlm/A6NUc2E4i8dcbQDffVXwi3keX7G4ja51PfbR4jtWBsH7sNn+AVhQI+SoxVYhuwUcODc/Djg5
r59lmjvM7UMlmMkKH2+8oLsXWVMigEri1ZaEe8rvG35jQ9sM+8NqVRNiclKwJWjZMXS3IXm3hDXq
z4xInWDI9LLVesW46sO/AL59MUptw7um+hpjNwqn6qMXWA6sxUqMX0oNqWjGKVRvzIzKHuC0Uyh6
HfNXCPV5MwxnOgHrISqLxobyhMk0KSUfeISexuQH4LFOyTiiwKegJ+hQtGGxcbTGw5zXKYNfIVcu
HrEE2ZzzKidksg+gwGCow3lbMlNZmWmti0PkR7b3Cki+ucO25k3Vlo6Q9Lxvp09GtzYQVttzXr1d
eFmxeMILhO7J1PsmUYs74q/wDmZYmfiQ1CZja8OJhWUkTIKyW7WmMerRKNqFxpYT89pEG1xBVXNk
iP34xn/znkfc3tcfEZDsohU7cyd/Z+Bglzh3jEa72PZl/HzMZ9E6IJuGw1yuDTngraVbQ5CI+lBe
9ypA6NfGxTcNMwGaxhSt2JTwRx+08Dgu0nfFbi14jH+o6qGlQHJuQbSnVK/vuzNTznvnnwufsRsU
4zqcSzOED5yRWAJVMvOVifL3InrS9Jfwj7bkoJFBrZ3JfsRbz9Ww4xWGV1NrC5THyTU5RHEuoc/c
DeVp0aQjlm7v6YiRSRIZcTQQcw6TPzdgbFLjE2LYiTudigXkTVchFY4eEg9Jd1Oby4gtb4UpMz5e
7qwTlXHYYvG5T4omZi0qUPxHeXf86xMwdOj4UlNFL28GMLxXTGvyDDeOzYSvcG8XKaftnmbr3gHU
2l4RfO4B6ed2vcrvlMBvKQKZlXxHRZhWXPgKOn3UxskCdT3kVTPfd1jwwxdeeObC/kLw4R/OATl+
R2EFJsqj6PSBs9mAHtEwDQ3uUBr00DuoJ79oQ/39G2NQVvpgDq08KLEb/VriH7yh8WdDfpnyd/rm
YUYy/HHGFvkvNQv7a8al7wSxHwW39Tr50kVn87mra9DTZRq+r3Oiss7a7Ij9eb2+uyDcgY20O1Mu
iPYrYCx2IMQDGzfH945DbR9syz08VNm7L14gqA4F4KDz4FBQz/ebh2H0/XwKLk66mpPgA8LF+T54
agQORB1Kg0KYzY9lhiLMN6wO0PQIra1yeDpKbHx4zA9P3jRs/IWyTOGBOzb8LBR/xydz1Nyj47ee
XSm4paAi1mKxhSbphd8IVLLSjCWcKvQ+dvNG2O1y5tLAUsL1f2jrTkTGRTBhnuLVFEn+KEjmzyNc
qcXIC/6hgokQGgF1J4TKx3wyWXCv2PA4p1u8PI6CrR8cE9mWhJyIYzqHhXVBecWe/aNQ4KOh8Hdn
vHRs8UeN8bmxXDTOF5M3x9lAHQLukLMDon2+qkpquUlmvzRQx4Y1L/3YMiCvzfFdoW2SrQcRz+EC
2l9IPdjoWmZn8XtcGZKi5btwhkaysrTqfBQKP/qcI/ZSDwReDefdNRcJ7XSbV4mlBv++hlDZYqNW
B4JmpbWtXEfvOB5pbeHrpOUdk+GTsVL7ohMUzqu7dwhhQaddBfYh8PnRl78dllLprae0Z6VLn6zm
E4BOxUSTHPgpYsPSTxUBjvMIyFQZPTUPcwNcZWqPSeK8/ibcRfjQQ/vgPNZOAdocyI+dPQ/2F9aE
Di6O9d/XOlmjeF4Dtyg4SwqEJKhNDnOZtn3r9mzplTROzgo4OVBJNTQyFaI40wCWt7th8+DDYipM
45DPZkoPAr7Zsitc9hYUKxJIRiE5wrXBM3NsS52HQ2S2FuhaQVbypx9OgVsmx8iUZuerTlHXOjma
8msO2N0adGUmbMFKr9rWmMFEkF7ErAekraFBRMRqBgrQYJamKblr8MQVvxR+/nq4xWWvXcrDhrBH
N+uhGjq8RsyIRTtA/zdC6RgFqxJpkDCnBjiPW38PR4C2TKfyyrlt+6SgOfbM4xCiP6CUda1gfiMq
89JAY56w/wkNfZQIHBZHxRlRvDTQ2SG0OjaHQKftBowLNg+2QWHka4gMBfzWcDPaaDkZXcnKmzuA
OCM+0IwXPV/O/WHeSis97/zsR1mjnzgQhdmJwUTOyMuHreBjpquOVprG5Sn6az/2aRkm2X0AfVdb
JO7s4TLZfP1noABdW/jNfifOib5WqwOmcwfJglZ5hhCvSx8gJ6cimCTX2LH8IMIg0+VFXbvmFb6R
5xnoCEsgJKIcueI0sA2Q3HXzTdfIw5xkg2EOEytL7NVrSUFuHk+exNYC69kvEUZue2PUcPrtGwo6
yyY4LoaUwdiRRaoQtgV0JIo6o+wVgY7FZMry7aO5oUACpTsD33EoZpqa6MIsxZJrJUfpdXRuiytf
gX0YydRhxRMGEVLalclIjUJHojKWCZ6eJX2/lD3O9KUPSmB1tWZUtPM1u1cqNlf7hViv0YxZ5P6a
MRvX2znmwqS8tn5wmF804GD9AcAVx+wx4bRVBGUJ5o95BYs2jCKOuEHm+f9IC6fFR0lKD0COTGWA
gTBufAWnjyQuDKEsN5SVIGAXQ1kydS9daH35lEPg38jtbYU9H34OfATC8MYCmWKmRwIfjLgWtTa8
TsEIOxYJ7kbYhi/0YIXme6URjIGDUl3FrQS0TmO2lqxc9U+3hD/lelolmIM1b9M+UjHJiq4x6wci
5JpI/XREu4rriBPyaC3pqjzKMR/WrYukyryqqe6NlR9TXpGJ4Zm3RW7NCbZS8+u6DCguEjZufEH+
3ZP8HoFCuA/yLIeetb8Y/9ufoum2EAXspfWypRlSRlR8z9IOCbANOOO4/Zr+jSF8blm4Q7o0La6k
h1KEPsd4XeSm0iyqtJ5VtXcGV+Mmu66Hf7jh7l5/Ra1I20B85l/ksC45fwhoXlipg9r3r6+UoZdY
KPhaLYd1P8Taef4IYmQa3WJ5Ak0LjM5wh/jjPcOs8LkkxRK9mBR/lJJYnq9tXoWJD0Go+pl1ykKS
+bHvimaKkHy7eAf9aNeE9Sji06fWTvNjLw9/jQcl2wx6WJTKcck2+Tza427gtK9FaBtk4AhtXXDu
6oFsIvMgFDn2HuaYWBUrctK5pAseR/oU73ZzrXK3ozbH6QJnlbIH+ACHAwhQC5MZEZToMBkCmNWO
MzfsNIJlvv+4vR3khAac5+HyOqfZVca5n0Odb1CYFu6Q8E/R/wowXGcql7BnsaU3TTm18XJMRu7g
cOBGZnEb0RqYr7Ys39ZblKfiUDEFJ5uMnzv4PHzUGf5Il0/K0q1CTWlyw+Xc8cJT9qrurL+EXkx5
Pf1yzwX0TmvJCBtHX4Ckbfh0gg/dbtrbzyjOFTUAG/YP0Af9w4NKve+FjYPa/lgbd2QLNWaRQkLX
VJEVGWCGb/405JmSAXam7bgk+uaXHKleNpPdomJRztd3YgW9IBaH2NtF0TNqaOwrNYhZzBDWB3jU
E6J1llKlt1cey+cXBctvajhwUUtVNF4817S5mCDMBQWmjCgHAMRNkri7Dyid5FavAWrZijDbG3rN
Kcj20MTJ4Zx3ilcjxWqcu1cfGsWX62gYwRB+dtrJpC+seA7xTVzx+7J+/dAb3sL6Y+eNeekucurf
msERRE5IA6zBV73FHpsAvWoUgBf7gw7X8qNzRO0UhdSAw9YE59TJFZu2eJzrZXx+//f7wxX6ezkN
xbtATx2qOUGYFogOGnJ7TMD+CqICLFeb8m9qpOwEOLqhJofP0Sb7XgdCj3PU1YklvzdXH3zu4EA1
lhMiLzCC6IbDX7JRzyRPom8rdLggdI3EKcY/Liz31WIkDeJAAbbLo5SYza9E14mWnVKY5YqZl+th
RP5jbLdwdeHadzavJpyVGuL64M85A+x6BFLTwMvOcrLZOoRklq/D67jCot+XACyaUxzhWsvAc7uq
C0fiSfWCozXfBJOPxF+kKP4h7/AhUjkMRdYh2JhNsvPXacgAlFhnsf4uHU//e2UByTLZaAV21Qnu
kC1pcnRcYVR+8XZcJ8/o5YjV+LvEQwiFGsHHAC3ETxT3s4sSnDOcwmXKTQgCRm1DDJ57bTVl130G
Lq6JiiqAli3BuBzCC0BsOcjXrtV0YWdzplULNp/W5BvVKpjdfKaqOIy+e6nwbOFuR/NgrHlloDJZ
u8ZsvS7lR/vzmDHrbTiIuGA8BiLqGhp77GCBbJ9MTSf0IZC4B/TsB8UY/1ZEb81tcxZNnGc3asJZ
2y+vl3/LpskQvMj7WGRzUsV9gwCo5M1RLgA0AF7pf+5VnBqTYUoIMJVZ+Yll+YXA7qnVfV3mkeAn
pBRYyF9DMHId/0GhD74JhmUktS8Vjecwme8aFQdIo0Xb8UTIFI6A1156NQI6tQFa5UwwwQ6xNt27
WE2bJuT6Ag4ey/gSDRNNQlRexP+fSFU4EEl+B0HjY3TtlwluzcF6Rs4UgsttjheZXnFYr8GZedow
0ex1mng5OwSOK6gPz34i8w6L4YeRP2FOX0N1/eDHp9VrKEcRcSMEkpFawFzOORGKF8a+8wdv84Jk
HZkgIHX3weZLywG6+9bOuSGaPWluxGIXRh8JXv0DvaCVWyPkqK78covc3uK6O2W2CSwncO3j120o
MOsVzlmOiH5soh4Gp/VdtPD363nl6qmoVUD2bO+ipZ4tsA+sdQPJD3q6A3a1z7HGcfbZeAbuEcfb
x1gDOKoz99rud6poPONAE7e9WZ7MdlfYnK6gfEWNmkpAQOIRLg20b2b8Oxosy60kOQ9ystZe8yB9
m22HBplr/E8DZgQkOo2YYshrSe6CwM+1MoAoEjzAQyPu8R5ufDbxWIUeRvVtJ7043LiDk3UePRNl
N/fHIoakEx6bbevYNH7w87T8JcE8ir+KDJI0XXup3RZl6TxoWgOSiolW8bnhTYS5XItkmoZUXW1c
dOtn5fwm62xPds9t6rwDz5AVg+EfLi4SN3xZnwtR2MY8QIUbYSLcve9ngrldlfcC9LixABFKF42H
qMCp50OIuakkxZ8lryKjZwDFU2KVwbkf1ORX3Z29YpxgODGJ8bBI8sIifQ+Cc6HBQmPE0kP6MoNn
aOFgjJSKdBViq1Kn/AvLh9LAIWYea9UZ0yXqpGtENr/p3wnFMiwIKxmkCXaeueiHH4szbsKTpIxs
YAJXLB2FG0VCWjO02h+0Lt5E7MHw7S7Wb/hr+JaMgKJ5iUbhawB6xP2JBMQeaSaIJIJyG8m1+l+k
R8AZ/Q17X3vPzg79pAfX4FO0+dztuDQzzSLceGP5iv6IouvRCiQdM0K1KBgLmAeYzH0wWTRAcWjp
o9N82gzNKKK6ZJHlHJuVUHSVFfThykoxOz/xcpJbiPF51Tybmki14Cq1SbJb3wEyY9hqqKHe9aeN
0+oJ8Q4Ka6Z0z9DXXd1159sCSSFz61s7F3+PHFewEqGbb3sTX+GSx+4Y8g9fkdSk7t8xYqED87lK
ZBcdy/pdHX6h6+7rWXRMZslaltlenViNNmp9pwhVMHkkSSiwfpaHKZ+FUXrNEu+W822IIiGH4Yl/
dYFhO3v6+0RRu3xDJ0rWOl1SjgvQ1CtREMlRNdfddU9SSGbsbBd0b5RUcan+iKq0NO0BSw4KKPu1
dixa73qQGt8sfBQGj1EruYkwueiwPSPAcwiu0byxjNVCyLamtJ151Rr/Q8T6KD0+VjN7a0zEy1ko
WjLTNt5jb8PZTOEL7045/0XdP3o8+uNoZQkAlwO/tC6hX+QBqSeQNB5T80xRV0X6fe8YDb3aAa+d
csp+LuGhwcQiKZutH26vAQJxz7dQrYSnELmhE+Wnd68vGX69Pr1rUxU3T/Plx2p/bZiHa6pLzNR/
V9tZcXcYxdTaeNLs/Oz5Jjf2ET63YR5e7IQXXcBEdyn9AGa39Ha5N8t74kvJkQV5P9h2QUyMvLbJ
Kf06RSmv4cSMJFnxmPmMVE58DjMl/TMzPL8ObmKzgWz+OiUBLmZx1/YGWg4WBW0a0O4tzgvKss3j
i5bTca5zhwqZbtA2v/7d1b50WBfJHTjenqdt/gFux8j0zGFURGfzknlDVpJguj16HS/iBTIHk3QA
jioV0ibk0jnS9Nzns1AbfTAuzz4LYEXUL38jl9HqO+/NHQiWw+kK+KuuQpE3SIBeC4kZ/edroqSM
u7mSK8xnpL5r/Y3exp8LGVMyVrc/f3L2iAZ9wZnIlMGhoElBAk26CECbQ/LTS8eHQuTV9WDw3bjF
7fo2g0Tg/UUaI3jUZdIqcsyZ24TPBlTfWDKE7tLJHNL2Bri80hPFD6H+B1gK6iz4Y96Ob2S76y8g
08QpQG/5gFd7ktrscmIqLpc1I0ICn2KAsF7GIk2fINYxOjiZkGsA++ijOM9PapFG4rhYpvwc+n//
k469AvmCtlWyAAUSlIdbmBd94CbQGuhIVrdkcZiiHlp1gvVrK489HhLpFyRo5cFjNhEFm6lluH4H
l8PhX6AinfiFtojz6oliBI+HKM+BjzNeOdNUrBIS1S0JIpS958f+ddsGsRoCftlJAfWvDsd56CI2
2wHdAlmtzRTb0Sy10YaYMI2mwD2au5IkF6Rc18T9P6jV+J//wgfNMFQv8bVtcl2p4KAPD5oB8vUu
vGD77X2YlrICyod4ZLBKWDrLPuLOWhaUpQjfmwOtb3zWqz3Wk1eqGGYJlJlvoOnHCCKMyNUXgVIL
G6R/b491/g1cdJ7QHJUcim+Ff6VSLjqlfcfmiTjvMOIfTsUx3Y1UUuIBbj59UP9awcc9YE1smALK
GmCxUagZwsN8A/wN0iFm1RY5xiCsJ9M2Jj5TuyCYc6dKlJXFqVcveqDtIQzGxc/QSQaW0soMgpXJ
nPrkG2AUIshiKF/N1fNHONrh2RqS+mWA/TJrD3dinrPmX/iA8zxr/Xxzxb39Gm1drHpCAMdm2oBF
n+7e8FPZcA01QoBu0FBnaxd2YzD6sgo54i8ikPRHsLhcpFDWC/POAe12f3GgIJKAHaPx9xaNMf8K
SYgFG2GL1tiLpqplloab0Yo3UY4rxqUQ++He4KUeiptW6LH6yCncYv5ZfXIaVvYvyPjx+IPGdTu2
dJMakwSicjWf9lJTEccM3W3NGNUMB5fPNaq600+/EraJLedp8qSisB0x2ditOP9LS+1M+1viJYNA
Dn/2B8oeFLUVKZ2fIlmIpOsPxFwoyWNF65cB68Q/CDIJogfJK5pdiBWuHThi4Ao7QDjPlKPg6fcU
MvdHSo4ZgQ6cLjIPvNqj+Vd1EHyuZiJCXtY8JGmZ9WE4LgPkl8GDhlG0ABo1F6kfRuYSl0DjYcQe
ZcMEoPgxo7W5WxlucZ2B/KlnVwXTZpTR0pgM6WOMr4yQ32UOWhwiNEFpqH3nRDtddVplFyjpp/B/
UJ3TPem8UUqfM1K4l1sLSZ8A9IIdsMSrcYUzBjoBd9V4Lwvqrbffpq1KqXaL6MyOdcd77Pl+P14S
wCTV6DQ1Hz55kc/7OQ9RQgMORqVzsL7rlM156LoE63JkOrH3kEOZu3t4roNTEVTLUqvfvalyFw0G
sX0eNtEhfcqw6yZQ0sqIZumEP/obj3k065OtPdYUMrMK5AMm/Zk2lv0IqbValaKyBohsu0sHeCzu
yYQybvbanPk8o+PTy5MbwVZEjw+/2fMXgBh7WEdldUWtu9lUz4+wyCdAVuIpzKTodifzLXJamBux
tCQddbZf0l5tydlT2MR6D/VapFEpebM7bUsBU2WDCfp/OpPxDNgPk7Dj7Y7CZvC2dQ0/ZBte6o66
g8T83TW0MhEIMf5JNEaJWrpLNy9sn2r2LCysuIVCzQ+XRqEHdDny5kwN36EadRlWLKdHxOBfKP7L
J0o+JnZoJb70lOvq0qJgMXFcxiAS0JoZEZGDEeoVrjiHMhYh9xUH04ofTjpxTnDeN1859u+skwou
0ZAjmr1lwJHPviK+MFM+7sFjQ4vthzYBY4962pedFw9lNbW7pfT1Qz+2OhOjGoiJDUoCGchTaMU9
ZX4KmqNjZjUFZG6r/sKZFv6cFTTHnRqNZSNZGN/MCqIKbJ7ay99dGTWUDopi3sQMAtnWvHNcD+zv
4QhULP1CFc8G07A3jEPvJGr7hAc0/fIyjBBBcQ6+wIOqm8mPRAiVvo9KLF6cnFk9VXA5kItzm37S
r7DC4xsWsLusAHAaxt3ynVZcD2YrrDQm9UWDYF2XkxRO8Ct6YmNipTW5r6M1AM1iv8DSTXWRgMXs
Sl5CofO8v3dnVL3vKd6PNP+tZHlkVVBh2CQLXMxaOOPbaBX259S4HbvyFMg6spdy1AsVKIxqwFXG
pNLdOpb1+fs0eOBvvXTNIA65VRQgpk8fg4ywv1hMzMVc8vc1LHbW+vDVXU+pkGCYwhK925h4sXEE
TcW9xdksEzKRMUTePPCuFBRp/e2g1HjScufdrV1uJt8a1u8Rd2Tpn40VYQCdMIavNpG/Sp+KoCej
fWVwG5qOGiF7socm++qQa6oY2sUcV7sDmVSJyaovsUlAijGBVTh00Xkx0zH/0nxmvTjPusnBp8R2
GWpA5LE5NlI8eANVUK4rE2vdAo9iu++PVOACmzZp+3ittGgeUv22lGL7GdziB4Dg5JWsKk2+8dnA
/eYot3vblkwO//JZ33a+AbMNeaJ8c/XXNKuXYouE+uYcMw/t71eiblTRO3iBwfSOM8TPuKChDjRA
4NjVsJdibV4glxvee4IkTgQyJ8Xj79Qj67r7Vv00u76lqnRRWP951hmhkYE4S1NsV1+tupC6nf4R
qIvHFpUXVCqW7LMc+h1RBnfhRXqiw/rvWIOtV5lCDc8opKQgZ01s7OwXO0JQSFbhZv1ElRMpUYF8
1qqyDNlIffq7b6ee2Jxs7VMXpxoR+qA7eVc/M0O4gCQqpMamWT3jeFmlcd99uJ93firvt9taG9tD
yXRoJp/sHZ2Ud2MF/3F7AcXkKSUiFsg57p+VmfIpKlcRyNowSTsU/drn9iedRIw1O0iQSoDA8zVB
sNp5p+e1XKw8G+7rAIHYOvsACxMntV0YVolZo5PeBW4ZmqJG9tc/SGp3X1dpbMxs09CC9fQOL9Jj
NWASiqP7mi1pk/H/dirJgRDEFngzHwvlIdGz+ZlBwMussP9qHtpWZAMnr66Qg568PLVHNgY/yiy8
8iLt5BJz8n/qbVDxt9UVyXlhjAmofSnTClUq8UbfEzYXy1OX+BI42PbwhOkjrfCSRLYf6GWj6U+5
ulSiYWIYyAmUe36CAinR8ObPc7WmHBVCSPjEhKp8ZBVsQ2yPSvrWiCr2ajodSWVlUbu7TL3/vWlE
c3gjWHHPIRI5gnwOonc42t9N74a20XplLyeiD81KXlK2PAj9j2K1fTjo2zUiS+/bPu5Up6MNwesO
4ETE90uB6PeLNY/ZDTcP6AyPRn9kzTfbChgj8h+ykSNJgOyraNHHJQc6SuStaid9yYIYnPvmX1S1
XLPpC60bHEOkUtmtbZgIDqBkf2x06HLuNsmiswY3Kidz+PQSMVdB3p0GcgA1n3wJYXE9IkvjYi5G
Vor/0M6DXlUbd/0P/g0K+YDBIfLszNsleZzGdPe8O4iMyygfciLJ0MgnZjxaLJGTe/kMw3lFY3f3
GEUWhHmNYw1n4xv8AGbZxviYFCK0B3XQb5+QidiGBJWGPTUR+lkoT98Nz9TQ3xq+lba/I1omceX2
XR/w6UTdFmSBtvb4vXAtYo6tt6PopO1YHLNGwtjm5KF5+fa0nT2zCu5pkzyVhXImki+lrysixSSb
4e2cZStQ5hsCOHH81CWtmNwxTBy8Uzw/x0Ke90o8x6lJvb1jjN65ZohBcFsdFyS4uXy+w7JzaBhw
jYnrYwgYXYeG5KkGaghUTN7218/fAdjTPAUlrC30taAX7JkU5wsETsjNTH6LP0E/53InODqjt/RI
df3ogxJhIOStuw36KLiTn/Q1zsEDeqJ5Ak9GEb+M9ZnjPJC7pgsa2/pWNKhQlOJhmpn64xrOqFJ7
/xCnAEvttdDzmGLT/2GKG8CO6N9v7YbPLkbElsIBRdkZmOSAZzvTNpj9ohP3gq3rBS33ZwhXWfBi
24noPX15s+WtFz+t03eCrE9zJ6x+8IdNG5vXpXMLRjAKmLxbPAwlPVpGzfmBJsf9F1twNwZ7NlSr
XJfbgLdMFCi9ujbyFoEKDSPMV0n9FLvyiWiKpbO7p7Hn7J4+xf4lSDzAMEL8qvs5OPnocGPyE5fx
ZCns7AY4ljZ0QwYvdcc/cO7/jSfH6sM9b6iYEqVx4zxfRGfkMkdn8U3gUKQ8ua9MCpeDhyCGOUL7
UYyvPntQqCxsYvisjRPtO9L1vyMB0E9cyM50kLWJbCfJkPAv41qNSjJmgJnLNeMQOVr5ag0YXc4C
n73zBK76P4af+TsTqvOKxcSS8UQbbghCCgiDHysX5VnPjYTmMSA9GafcYnovAH1Wwqp8CRDn7BAE
4aJIrYwV3kCcc05uhV2LkHeyk9NHauRRArBUwk34P1CgNaU6ixwOM6lNc+qH53VkX6bRD/yjrvpn
zFLuMLd+GLfsa9WDQdY1FPfnzz7cL4dLfH1nPwOzS3skgvJ0NKumDQHFJc6wg7L434M03TlQKCxD
qr+3ncATor3/RY96yGCm8/btLyYyeyR6TmCnjyVMYXp9T3tBHpJ1lPzv8r7mH3898jswOKPFKrE7
ycgPef3bkwgsucXp4MCC8PrQ0ZA59mBgC/RoUpLygAP9fz3ZikKfmU2SiqQHwMeuBRJMu3jyDe4T
OcvXaVYb7BGktKF/uWXQc39rly98gY8VcV66AbEox0a5gATf+rd53paWhfqivp8Oq4Jo2eB6cM6I
jN83S0H4EnYgqlh3sDm3d5DS3c7KU5FFLAol6Wa6VPnmqGMdZ5WL3cH0F1JzVtteVaN0ce8VG8tO
SKS7/Fcu+Z4PDPPEbjMXFe+apd/6Wy1236LE6hBNWmR7I69gGBZoO/ZhVwXoYVLfVhKxJ+2jVGJV
MNcLYtPH5wj+PFiKvyihm4KpT2PceUvkJ2F6wtl3+EmJAIprdu85d4GdleVEKatcNUu7ZEZEQeb4
haeomZMi6MgZJwRXDQ/7wTSc9xATWZF8AoG9JhQqDxs3hud00n2NH+UpsPHRCHD7pgVMvNgEbPFL
StMXKpaqHvA6OmLBbu0mE0rxeRfxwoODpUkwy33h7g3ab/ypLEVpZi+J9ltV89CGImW0ySkIJxDc
xe/0U+inYtJtdYWcSxNd6h8HxQCJJwPlDVbGtatNI9Vn7tJIRtqJgCn9eUMk5QjCxNJEGkoCl1fa
I2nhk4chvpPVx0O06AvVB5bfrXwnrExmb0sJcwTBMnyEzt38UsMsNGIrpsbDksfn2u6s29h+Lz4P
Mihec1lHrLVHzZJl2mNtBHtTCtj2lJ0DWW97/vvk1sGfar9ald0ja15zgfRtjZUU5H5CXJgkc9IC
XwhtOLQfjl9RZgy5ZkBKe9wntr/Vk8IxR7LwbKqH3wIrXPBb75QcabC4vFvR+9dlMkiYuIyATefi
szIzgq6rhyK8BqS/fCBIZjvsbCCD6JuWaOW54UQ+fjw4dBzFKABuluRmxDlx8Ea6Fw8wBsQ71LYs
CTSJbO7m+An4Sat7zy56utNzzwLp/qj99LuyVNFQDlTQHXfmRIFMQ1U5MaFAe5+1+Xja7nNcWXEG
4vOSFUVDRn5iEvaNG0X1fgPXTh/+1pQ1uYvb08IDmhiOMi2rk48VeHLcu0n8YI9b3Fu3XiS3jGxJ
e/nJAb+k8Dwfip7ZQkH3ZuzF6F0ZIr+5H0VqK31I0JWwRNXB9dsVkv17EZL2fiQs2jhXu6sWKlSV
4RmbWsF0Q5y5cI4X45/na/E1FGhEldnA7AFk0Hpzklw2VV8auMx5viVujlzQYJSqcLayXlHtrcgr
e9JDeh6BMohaI1Dkkxzaw4QVH1veNUEohxxhuRL32DsZy49KLVlo2f4DxDsO7ZM1cU8vmsYVQ1SH
8cpcGefdWNjnhRzSqwsa3NmaVjycTtKSHvfsQD6BL/SAtK79D9Sq61u4qXj0TnAY80hULfvIfk/K
Ua+gurh72ohOeQi2P/DRL9JzNXD6+DyyQfzLLuI/+E3dGpKufvafPmGM2Be2q8S/A2+fEgPqReu1
vyo+Lbb7DjRvJincU7m8WyGctqudAYb7u11FoUYEgcDmlxelBXj6UnmY12isZnsLZ+VfBZTulCqN
Ev+QjVUZeqi03DK5lUiOrQRXkuXS9rSTN2so7WsSjkobKnHciAQCXRFf0T1oorCrvmTJ7JAucIkJ
anUFq44R9MrVdqCDpiW2vEfe3BwX36vyTRkyoKIO0obAveZBrZb9E/ZeX4JlX+qmcWcSzdWP2QbH
OcaBnJKuFvdeRN8SAJyD9qdhpSJHuuJWaZHWnLTFLlkKZNxLPS1tzflBdhxufv/y1A5pZAdh0/lG
OYzikXQQUdiZNbWbdf1acjwAzF4N7E1QH64sHsd0fgDaqfh0v8+7JsRgElcxj8727h+3A2kiDH9v
mrDCB1TkimQSNSpxI7wBDEAtMBDu6BBAJa7ahPU06LQXvWYvD8TXYmyL8+MCQfaxw7CorCH3T3Gv
3gTPFWVJzX6CqdzGeO+8JDs2PGrn9Fv2wEYaKS+LiwUp+no+9MJ786eBA3jnCwiyXnVEGupyU64L
3q+W8Db0UlSflbCgTMfGT/FHah5I6RkFYnRdHwy5jaTovW+sSVVT4VMxIKFV7Ey4Ygy3yeEb1+Xx
f8GowSsbszOH57zHtWKqAda9T+N8bnzFgxnx+3NuVF42nRY0kQcvi5z1ppo4NqKoDLKIQSaLVPlI
rWxzsodOmHXFT4/w/DUkIP0YLjPC1qsG+qLWxpM0mhN56S0igVqscgH+xDTUq275HmHnX+Ma+qzT
2ZFYqw9pl8MjNroBRu8CgdEjucRG59wmx4cAv0Js36xo4OcLNH0mmyoqPkdiOiXaXo5+hVrLMeqL
9r2dcVH3AeViirasBxPnq80Gy8SMdz6sba5QeWNJETtmEi/g1Jsj5Bc7DOZR8OBTjqTixZmzg+kw
jb87YyBPXr6CJZPzq+Yd+qRt506gFnYIXmDbprIU5VoNtrHyow0MLTDiuVo+nHZo59GFtmqylZf/
jQZ+WLIdWYJPXytUYXIq8Zdhgxpke7vob1KwNAuVr/tqnHG56yVBn2leH1qIlsMEBNqoTMvytOAg
QttdNQASCbx7q3br1CN9fOLJoHd+9/o9SfJGDz4AqVywV6dcSp/HPKdpVuaqWMCJ04UY9/+gyhri
JHB/hEzTKYgePfUWhAvkhW5q3H6g9v0oiEAcRBqRisSImReMHDU9TXsH6/hD7lHZHYgWwH3Shd2D
gyaCHmuKS5skMMAlMgLI1DE1p3kHxUki7V9XOmiBuGwWnwYcEnhREhq1s/9ejdebNu//soimwpg1
IfNgbkb/NyjASSKkYj+yZo0YtkWj3G3jK2u5DIQOXJRaBwU/hm4jvmYk6yMjGG4O4yUyEQm5jvfR
Tilq8zBVCnm1OAthpgg6cycqVFmvjDgQ9/ymrgjXD46WFK/luYj4pxgs1K/6gIeFW64LbG+tzNBC
I/FGlsqlLZ8ehPh/B+ExaEk+/7U1TknhJFqzSzrsN92k09n8O3r3sV3NNfGBotnz8A1/TrBULt2D
V6fT7RIkiksS4QtPq5p34uTouUEM7F0s1LB/ynXtGSbyiB5oW8yqgOfqPBx2HaVe98kgVFW7loSW
MY/agxRC/UtSmrrI9yWAMAAWkfr8UyG9VYlbcPeAuriBs2UYisCDD55Dklvo/BgzN2YANiRVBM/3
o7sUSWuEJ9PkNPlS9UvUqB0BFuyMuNso9sSLghVJCNFt+sz9JhmSADxmLkt8jw3KOZAT2K61F9ke
VfoFDBFLsIf1EyPnR/hDqdmmK8YbrAda3d56pPc5qp3UhCL/4fG8I20xOpBu02qlMwZwpJCRtNA3
FwwncVkzc8ECbaJtnFdEEMcLSYN4YnOnZ+dAR1/p+35A2K0NwyJG0FDoyxGxSVKpwBhL71BlQZGZ
rRIHCSxrLvtHl0hTm4XWVA+9SZXc4mqLOdFXy9/DbY6cKSN55elfNJQH/lICwvdNaWihhNidNKuW
SQTDRKp1Ym17WlzmQkcfTxmpjrvug5XjXuOyQCK8dkGzHseMNV+3s/UdRbnuKb+BlGnp+fePd2AI
QJm05Jet+3rX8IRby3CQy4c8vjqVQMDGCM7obXRyz83Wmq/UvxZyHwDn/Cpbu/OAa7BYdKSEKyFl
8ZBDGTYAAKOonmDiwdKqIus21rJcol6f691lFpkOzaC9dep3CzhKSEoyYqF3VAKnhNcj26mZMKY9
Odx5EVvqN2WEHr90snrvSl+Txh/1XlG9DsXwRyRbX0NfA5fvhT2IcvK+jYcS+1umvTh7X7zEHIKL
Tb3xyEyjdDan7oOOGpBXMAnseocYZ0/BPkFtgRBBzXB7H9E+AdHqzBkF1WZkNe1ti+0qiJNJMK4M
5wR9CoeAaoj1OiAquePVikBdXS3eHLzT7oLRRnRJiJcmJpriaNRLRR8n144GTGjRhCGwmgsQEewY
orma6Z1L2S8kZVIk/bFFiOLiddwsEAO3AaWD0q3TXQcN6SqDWD/zlCCBhw+io/xLi8tDHNEgJVKy
qfDOunT/jSTMVWyalGoJkAGZA8vtEwnPSWTkKhyo9SxL5qfZAvKn+lY+tx9KvtEUuw2QUk4XVj3b
0oylOJXHNI2WYwDVkTSJ1GWXKFVRVeH32VtANmcA8K0nlk7omOfjBvJ0lLIeZsPc4PbD5KVKzG7M
dSTa5d2GVKQUbKzqMlpHSSYTNhHDNjMf5O98aOVmjTSRHX1rKG8yWr9sEOKsuBtWt/6h9TK3+a3N
LiEZuL5mGSgYW7tv3Cy+sjDC6AloacWgi3we/RIIiCRxztUex248o8WsHuLmkP6wq3/YGarIr08+
OBZnr6vWvh0yb1rHxeRgAITD27UGcVuYVfNin2Uy50UVikTTSoJ/XGpAvX3fbRiBfMCf5UBiJzqV
fhrnSrfQlsjT5HR8Rhp/Ns+zgiSR/ExGxsEt4nSbD2cbCR1QvOEsy6UlSasL23l2uCoAjg+fWttL
3E/bZ4Z4JJ6XWK+J5lWNbEe/Dz/7+MBzxU2JiS1464ecVn2QlrHgDY7ahhtiPiCLI+Hu9FdgNQbe
WAlm9LZ/GEPHEaGMWXngYGibYLAf140xLHS1Xr1lujG3dIT3ZSO36bVM20rCU3WqCFRd/FY65nuT
o3a9xd/q6qnrwdLg/2brN2JKSZw4u+Rjw6ARqHMb2zS8snt0SdE6FzARyCGIpFQ7cK5Vqe/kiFmW
uHkEArqyL0BHbAQjN6Oa0Yaudgo1QuCBwet1OUIQUAIv1S6NL8kSY7VAE0wkQ0gmmMsulm5hNMJE
InFYVx+mvQ981OYOzEMeB+LtsPzWOvHO5w2B+2Iid1TMw0iGUzY3zNqGdw4GL8R2O5XNa8DBXnHw
EqV+aAh/IFrGP6zcA5TWrbUs0V0QuBeyrdKHtKt60umrq7mP4wDBTA05J16kKV5/mT8WS//NlpOw
9GGVg5vbFSqycHzmQ3wuGAAbVjoz6UOkk29giiDhi3NNO70jRGioMUGeG9rlD6n+I73e5RXgTpQd
2LwJPtQyVkWE1DFnm+eMR9dDpvYml69nghfMHNaSYn3Eyte0IqHbQjU5dkIBJLqxiV4cKbf1QAoX
H7vrxQ025QCp+36XVFIf2WWpmVa1Jm4wLYTIMVNm+PZh+27t+CGMo615VZUODzQwQMTqFO7H14Ex
gQEXyk4ggI7PLX9yG/aC9oTXt5rf0qYm/V/YNuZPyEZOrAn3OUv7iyzTPY9oUUlCfODuGmRGICDV
2ubCuJwdZxgitLpnSuG0U2iLSSZKFOJEAM4dDwcXHa+ALyWJrt6GGVF+wgAY9/oWgwfSvCM4l9J3
g3FuvT+zfYsKob3YCdV3TCTFuWhoOJZXyBO3lMhHgE17bDuSsy5nnnZQWZxMM6nl+IZWDoKWBKWD
jJICaOPqrL1S6jgdIDHEQcC7COr+ceFh69spE7vHfptSCe+NDA8KLCGnLqMzRzPO/zNCMcETY37v
ZosCvfCXI2mT3/PIzzWaxNRL08hIcxG/dEbfbISNRPAoL2ChwiIYKMLHfMjD3keBimRXkRGHcbgb
OwrXvElCU+XOrdCG4BGV36HTSvJjIP6UcCTwafKb1SIwDIa3qVpatFWpaOxHm4NhGMSMBj6G3usL
Vq7v25et4DcJqmzm2is9HXdPrX3g6ETIG5gUfkNTu2C+9+4ltwN72+gNMhuWv3TaooQzSKVVjhdv
2Ph0A/DWp+sMKQiYOG4lcz9SBYJIwO/tcN/TuadttL8QqY1n42CmBdkRY4zk2N2KqVNNDWpkdUZ/
msrhOHv07Kv2fOy3pMgvMhVLj9EE37a6b6IiosgVOw2qY6Dh4sVBvhZ13vK7OGRG+aB7+GWa2emi
HPc5wrDbh0c5lUZaa4O9Cj99lGLv+xI/sLweu+62degR4KhFhlBfmkm7Kpthyee4/2vUXFlwcPA7
WpxcXHvPwEsvb2NkCC7c8AKRfjaEwmhIUrRiLvczBs/bHKXK69t1o3MRCrp9llASs/LcuqUIBHKz
nHoCfk5i+MFqNCpMvV0KVdXDJlPqLkI2x5fizyQfdYrq56SC2tiyXkgZzKeWZ/79tTn5POTvsOJ7
qfFgtElBJKsgSyo5NvLQW8HRCP7ldOfLogrzVZCGr4LTb01U7C+RZDgufzvjWzAmea8djEsL6lG/
3W3djgBJJtuESDaOI3Ca3eP1nxoIoVHyjG1aOTcPro6hrha6rbUSXZsKVIkZMcuL4x2rgz/Mk07K
S9/LfRHldb8FJbGGAZz397znGsSsyOeJ2TOynanM3HS27YH+EZbhSSgsEZygFtn451jPWOSK+dZw
gEX1BDD/Xn0IAyFMOXcvKPcswfFrduYbfOZ14oP530CuQGrQElYZNCQFg1NRsaw3ozURZNsuSQ5W
Lejpu6BosY4EGtKiNCPNcWxTebWRuYgcmKN4ibRBGj70djgHc4sG9bvaNgORuc1GW1hQZZzBl4IV
rfVa46A3pprnURvDyKUyThYjkg/F826chzHZRpJDXj5R6Gq8ViWP0iP0xPvDwFO9/29XX3iRjIUa
z1vOKQsn6/6mm60ZUa0Pt6v1IPJnhEmqhqTfbenpluSHSq1EOcEHxHXmnV3ypiJy7hURQPDZkD8l
8UUgSd5uJzMo3H2CKNne88peZBNV/fra4KtouIHHNtBsDlW7Wz+r0HhrQlt/U77oQtnsfFx1MXMh
joMNXEP0v5fePmbQXBe1ZkLKyaABznn5nX36WOFV4C0/Ci5NIyoUxaS+9YaOhbq+S3vaSqNzsvH1
Ozy3U1p9hDO+mfFepPdAcBBprVi4DdGPY56SCv5mcc6ofT6pxkmpPw1hBXHBfiUx1NThEFGRYNMi
8OJ2t1m4FIPr2GY23HqJpOhGbWxN49FOKxWv2PAqXmSEP+q1+KSQ/+VS9A8jmTvXhRsC5Ie86V6w
NXPlzml8gKP5jHuMX8NQ7lgEQekTIovRte83DmaOO+YnQjME6gPYWKvEqc1WAoLMBiydeUnGzCL+
CYlMsFfVeUVorl/Xo3+Ivobdg+1i0kAsQx9YImbD+szxWFz0ufLqBiBvx6WGe2LxCU/6Ug0/fWHo
yPMDXAc7AOewQksBrUIVQWQeemsWcKS+njOqt2ecx9m9CoizBnrmO0AekLBDUO8r31N6PK7j9gJ1
3j9nVWT7HAP5S3H6kKT7UNTKYWeYpN06ySvv6rGVBx7JdEn2soiv1I5PPUGzLGllLiyyXDMixChX
JGW6A15Oa3t0MuSSBokMNcOuWG80lpIVpgQleiZo1tAUr+pMTLyEU2Wv9ZNtKOqh39XX3X1uVgs+
Sme+iY6soxjc51iW5xKLRw7V9HYvepmftpKd3XuqPPwFPIzkHbLuIKUBcXAr3wPf5j9Bw8Vmn8qX
1+GNjl14UllW3bDLXvZuz2W/56ZT7RUunBav4ekGjiKmkA6v4aRgvWt/Es/8s9cS2a0Wnxp1Zp/N
MuGlbXQYazJXn5SusBGnl0UhTs/xe38sOzeQPYGy9Mh+qz96sR+ZTb6eMBw8wVVwstzoNjHhJeIa
rqAbMAWAWRtpwQ6G1ePwzHOJsqfiG3gZKKnidDeFtwocmCWBiuORttUTnefiip+a0zgi+RJRg1dP
iJmNBzXeWPl1SD3gPh2lBNlJqOYQRaDPxU34Yiyc6BcdW4NJ9i0UyOkPU9ptB4BnQz63DXMN9ggF
54JU1uGMYaVd2CJ+umsPafZa5tH86fPmsvBj8bPIYk1GAsvHm4nPyCSH2CH7f6Osxz/QMc/Kzg/0
oF+Rt3TrId20q8sUIO5lz8Proaot1XMRsVOxrseZph2d7ebMaN8ty+GAv9VrKL2YDT2zklkWAI5+
uJ6/f2ywONO89+yqPxEYjJ7pVPN2vmAhdbN9KLWOChuncCQ2t9nfRjmQqr3JBv9ah1ZjyXkSol1A
hZheWeW0uHp/v6yHAUSAYjVevCHVdsyfqG+Ia9LyJOHV0gvHtmUgc3m6mrCL8UAiCbui8zIvuD7u
iWnaz9SNvEr1UmnJbTgNsoPS9VBYlFWlvQ6mCGHJ5vpnT/pvbJppuqecrqMd4g/nknwck5flC9KO
9YL5SJOgIddQTXcdkE5KnrE3tkOJuxiciTE2MG3/knrUs5y9Ar5a+Au3/Yb1oq6smDwjiyfgcv4s
P6yhyYoP53mLJaq5w6XYlV+aCNwNULnRAzI3C5uUPYFDhojZCRaPhNW4ACBIE9G82m2+XIsJDN11
qup8IDlaynka+Q8qqbHj6CQf00PDVwQiVr76HyQVLOKWWLWN+rlpfF6kaZRVNi6D76yloihvMIoM
wpf+w/MHrv838Ieyo6GqL6+gVLsGpuJEGFrlZ+zlvSafsMl0pDFXiQPc/BhOE035lm7zqWhfUHfN
Rw2ul2mo60DK964lyKI+ZTOEyRtqZMoC3j/p5uu0ox2FmplkaJwDsoj4jPTa4qlvnA1naRk6jb6c
o47/ana5ladNMOqu1c2o/fDG6WtoOmZfytYnUzPG8A4nxHzahG7jCAz5QixEKsPRTnZed1YAE/Vi
r0aegOMGQO2nqdAjaIX1neHCCRrkx0/ksOhic5CJkiPxN/8ubwxU0SalwuhP1Hdre5+5l4lOkzC3
ij2P1Gv7jn8PSGPTSg/SsAFFNdWlIahJVfZrUoA3jEoqyAqGV5K/w20FbR7ggHsf5cjwUNNZhuWW
+AEOk8fNa7I21jVQLUsivG6dQCMazUu3WaLiOYVrcNiPqGMxc4+5/n3klmn01KmbyVX/oYjCR1KF
TblSvYuGzd8GsrIHu2y0aVF5eKNG+Ce+oin7Ewq5G5Tg/NVR7Ad8xa6nXoVNg7Ix0mZihVDHJKri
BvZU7D4vX+nBPBmDeedGbqDpgFVG3GVSu5BFxJcN5JA8+VXjmKQlq+nOaKTV3AkY+rKNuGruhug/
lFINriZ7lVAhyoqxr+dFugFAHvklE5iUVUl8/8erpOzJpkr9rltCJRsUFSAZvf4zzHqrKw6L7CTi
G1uCHTYZipwLLiPQ82DnhDYm6dvfeD4hzdFwx9zKkfEDH/cDLoBr1RqYAznZfy0NKh4waA6qzLmn
N0ZKXX+D2+anvBO/hsVqLC3r+B5jtnbIP7iXMth94Jm5YAE30pGaVt+RcikJQIqX9IXSyuiYmTe7
E5sOwg3UD2UMvKsNpXbcG63igYxITX2WoZhTxr+VrNPEdGmHDf30q8s2EOsO114Awm4niUyVZ206
UQkoP4kr0iP7dMkAYhPYjIZyBFYBXBZAryObFA5beceY+k9yM5Vy48F6vAzfPr1Te/A8AwJLW8as
W20VkQ3u9gnC5Kvejzjbk1VUiGRUrygylSn3VOgYkpcWkgEv1YZWcxwn8uViKhgcMCd/BOIuyP64
j++t61KJR7JpoVNTj+gq9+ckyXR279uoVBqE5B8fbWRCBDcUUQ07FBPkMTrquErbojRv6++TY80q
YfxQJ2Q+/KlhBx2lhE91WfsGwZQMYMPKtlvlMgBilaqJBQ+oUvQ4mu+y+SIwRckKMg+K0EVxIiDz
XM9y3hBf05dC63VPMVNhdGukC9v2M2AypMZ1juIY9oKEALIZdWIxTYjrosC1lyvxGPseUppt835X
Ij7tTYXCZj2j1HVBlGTe3ccC8tEy04+WZbftnA6JozeROsrifIpRKPeQ+si2ORC/qozMbtWw47tu
k/OVRsj+/jJABICS51q7L1KiVdZm/+Vq5vkPchXS5jMStOYRcahNrveLMnWqLE5QRM/aTkUVJjuz
1Ni5A2cZ6eCNRXPGu+tvO7Ln1ipyKbCJtRdQui9LIfD2dJwBQC0l1H3bN+2ei7CKUVAT9kNfCa8T
kvqTA8X7XP/I8IXg6ytvIhuLjT8oc0BdInDdwFfdE0gawgf7MFIfe37hFjhSJOpAf+o+RJNc3Zoe
79A66dc6dTaoEVrOmBE7K3tGBFdfhqjwbvZGht2yJ4EvkfGcXS0ypHPzmjAqYO9j79hnT23PWEmM
/EaVrvgcfA0yenAqTjJ9qL6XsrJ4P5j4f2ufYMbZSqjyawAs2xI3GJ5ZqdEDtHZbZW91UP6m+NDR
SNunkRxLnz2lNlliys/iPv96VE5dovljvP5f1LAxJ61tYbQrUL6KkPDB8OcwZF59gG8t5W9el3FS
MTD25Nte/4kvsMOo442+b3G7sFEv3g7UuSwmXiPscVdlt+09Xv5ZqC8dsB2qtNrnDwWKNs5s3+YF
rNetGK5sG+AxKyjrRgQ0RWD/3mPE5oo0lejahQFi+ETsTLM2uG5OTr87OtYpaG7bfqfFiz3ddlQr
O3BrMfrY2LfVAiQR1SPQnTl5qMO0pU6YjnrrdRww07cQLefmISbwhafz1tyzJyiKLryo5hJyTwmn
+wblonNd7PlE8BbCoVv9UwXb+DAf5r/ChhOdiXZWuH+jHjCnpy0p/9Mh+tFFnknjnYIpbTzvYEcl
HSk9ce4CH5aSPHt/gfBY+SyPRe2pXgy+1VF0Dsbeeg4/StqXfzLYMD+ADmfv/FdhhYZ2uDFRUvN7
PmNj/DHQEq/ijWl4jZuSziJukb2fgJWweuxxdXoF8roYyC2z0H5cOD9ANnkkiaSC/Zz1a7/VQnAh
ih+sLosblXPmoyVjXFcCjMHbaUa4KwZmrSrIq7WpwjBhJjNrZiobgS9cf4bPK8jxosfjxJcHr7wu
JHi6p6yT1P5QlvxxZpJA1RilArDhcG+TJ2T93oY8MOZfqACUcdQaZDSzQ9hx99x1Gcg4jD3Nr9IJ
PjQiJ+v2QlR6cwo534KShHhEVtKBO/QJRaHlHBAbAKpX7frLW/othnJf7oYHA326JYc6oNSQrrfs
OXtUDuhixQg3aLk8rMef+uJbLl5+UsANWwDgfPJmjiMdLMgzldm3BhAvHx1B6G2QJdadfMOhINtN
lPQ3A67QUARraMU6CTjs/ycJK+NwHoBbam6nMU398ZrU7493+rr7VnyyfdGWh43msu/JVKELeGp7
wB9xsMaprtj8sB5XrCy9gFBE0LogE6Iwgdto2cgk7JrfhPBvYN/uF9OTaCpd5Cy0Beyll03JwblS
pIjAdyGSUckdyNynZMB4kgjzyOdjMBil3jXWKoFpm9zT72FHsqj/FXFbNmfFfQ5p4T95WNMxNmDb
CFSjzs0ExMD626XhgHrFPjzM6LPmgJgrbKLxMKNbgyVspMFak1SZwPttQBOQBStJI3McQ8Q126c6
l8UfPBr0nQuxg0LUNEZaBCHeI+mU8tFSN8nboLp9P2/Oxlf5+iunSYXw1bpqVc0jDwCaIXYuTzbA
yfqdmFRRXtL0FalwMN2+G4xcu29/B0BQWQPwfuGsp/kDzFhXTv8G3FlbAbZu/FQZCwkLdCc+U68H
dXitYCuhoRnIl3TzEGdrCq6PuDcNFYgkPMySbmx2kO6PLEeshb7mztGy0gPKtKA50yF+9p7ZNKq4
Ydp+VT1mv9vNYYzDyf7shFxGmPT48hD0kBTW38Gfq+r2pq1B2f+Hxa7b8XmngWmlcJ+1AFD0ND/k
/42LtISX33Mokl9f3x9IwfQxpns1+pJh3syCEx8Lib6nklKtg3Ppp5DkaV9fhpE3pt7xssNE06h0
KUmSnvP0hDCX7sg1/YS0Rabz/UmAR1OG4vXOe/zuyFd7Nqwg/AiGSX7cyIIZcTxSCMkXWrrdPp68
DGVgr9ZxH7FbGmWf0WdEcTNNTxpbCcfetvMDOBT2TfONtfaWSjw6T5VZB2j9rZnhBXxnKhGKhKFg
3UCvwrGucoG6MUy9xm0snVMBoyWYr5tQ9BYMLv4qYDKGtpWGxeUSlPXOuCR+wvuvgecYiyP3/McS
tb3EtbL78wOiYBjOciI3FAGE4zfqziAtf1Cra0WoSGtbyzbIBJOJJZx/ux3nQthzsQlGermA66W0
ubdficJrQXQgH9BgapuppxUryIG3TQ64jlC0QmfrvdALwjGv5Dd2Kd6nn4OsezVJKJGA527PvZ51
ccbDbWheVAKO/poR9dm+ZCMSneh2U9BuQQVK9SFyfr7RUhSwKrxna/oA9zXM4Vj5QhWoNC7i0Jcz
2YZ/r9mF+HYMRAf4hhj0sJgQihOPPapvhQWLem/UzwO7yASPMv59A9MR8S+bMPYDjwHNcElsbtqm
32PH2qRNBW2UxgE6afj2zuflrb1UYRINe+/ZSS7PuBxE7BA5ApVNO8IC4Dz5JAKMZiwywghRHr3h
P48wqOJ5BMne9XVXf7eMlQ+V+/FB9QpOHmNZbeTr/hEB3WOqP9U+Pt/Bmcnhq8fUQtlO1Le41IRZ
JCgM97VFeCDWso8NkohlRix1Ooc+xeovrshA265+QESyI7XQw+AUpEbV2UsHtCGKPena9wqd3M08
ZtXG8bnfuOsyQcbIT8+m006/sZ39Hy/q4qnj6tvYHXi+Kp8KbL+ntFS3x38kZyvUYcGA8157A9zk
Vi/zRv4OlHOAbIiGQ4XUIIxBL4VZwTGPZZUs8XBNB9QmKflPqo4jhbf5M777GWnWdN9sJY0bzZoc
3tXQ9/hceOm/w/Am1R4VaTfZ9qPFyojjj05YAn+tD3TqmNp8wBq6HCPK9utWRBq073TvnzBTNJT4
RSHeQj28S5PD9+Cy0UrgsPO/7IrscD/9rn9WooPinypGIenYWK38/rQlnWnLNZZK6QO24z/76M+k
rkxuLpaOOxNhanu5YH0Ep8dQNAxI9zrGL6sxUpDLFztfTL+VbzH1lmuY3epibHmfk3mCAQfr7uh7
0mcBn7SRuuc6BH/pzgBRJdUeQLCJQPtvYWg2USALstR5eifctkslpBIBvlhPEtvpeBvHvS7um7Le
bqkVlprDwW4S/Gkk3gXRmFoqocdL5glCWE2AwCpTfRLuRvlovdGW9FLPNYoH1e/EYX3UMiFmW7fp
lK4VLCjfFp3rBYHVS2UaxASb+PKK8kpE/ZQa3BFdUCvTYD6rrlcAvapP9KN75IvLtoQ8+b4ukgZq
jfUVcqZH+IM4YXmaItv3kgO1TiWbsvyNYLzVCDsu9Nr0Io1//xshnCWTZ/yKJjROBpm13YIj++aT
Jf5egEIChnL7UU35DnCh/1mi5ec/uKA1MRDDMKXRNAlTJwOu7ddzkjlkD+arFt/9AnvlQOOqxFxy
gOTl80Q9wsHaHpCJsO0tqsNzRu4R2klwjFtvxvJL+GiCBGy8AkrlnJZn0dQXVlEaNdK4vHKYh/D0
Thn3Y/78pnEF3vKfNDT+UWHEZ/cO8OpmiX2d8AfWrAkoEW67xfZE5E89G/IVl9DRn3QnhMwu0lcb
oPWm5Tr5GsxgRTWt7x/P1rr9P2qWfRODfCSOBCavhUVCzzRnwjVZNdH1zYgyi6WFy+J+SS318qmH
DPDVhXdxr7f45vKQsPks9Ao0jS0pqba28wADkQZy22JyJVgkv5O8ibT51Cb9Grtz/0SftywzhPf8
R7bhzm9W0ZwaY7fdygtvNywz3ulGf06/YCI4H4vZA6AFDdySIwv7o+k37ykjA6sGkHJcpR3mUNrD
/lmjT55t2yqsu9M2/pw3aMosUv0WIQdtOikM7dPTxHHjaCckB5LVRBCYPiXQSlXoMDalPokzWFMh
XmQIX6huJStR3lU41pUbUgc5KuI8X0mECQsazm8E1UobMdsP7nwIrC9pV3rEXD+B6NKoOPjT61HM
L37VGAgIe1nZiQo2XYEubqMJn1dMBsEldL1Gzrc4kyka8lxKQUxoCa4V5PFX/PI8jXvUugI0aXcZ
6YjM3v706q3y+f2vmkrFmMHmvyMFLzkrFHlxEc1spfwkyzAJlCZ00wcMLDb113SgrKloWVtmUuFP
PR5lLvtYcFPtMlAL0A08nYC//1Bhp+wjnquZQwO+v4C55zoEiirJ/DTVWLu0G5zpSDPZm+o9j5YA
wFCxPdQXgsRhxqrmYOVyOAedkZfn9II47lGEVTOnmz5nz0ukvc0Qd49voF8Vb5IvmIF6Z6/iCsZU
ZNUbQVbVwzEdYmY4A3SaPH0fyMA3lrE/MRVF5w4Gn4r6nVt2OCyN/K1KB13pZwUwO3KecYifGzA0
fISx0iO5+xawsjcmm4+9RKRjfgN0tPxyHiMjlqyywfZBiUjYUrWTxFfUgIHJe2YuWm+S1EsjEBxL
ZQPwLe5TMFTbP2xJLZjPTJh9myiAwvVp/SrVpPTUavZ51qk3Kd44bN/paBtTEslvP0HKIH5LaO2A
BqW9A4ypuurjzV6nD9mQ2muJr9UfjxBqhfWXujJOXKdOC54xQ4UAr+6AaH3Cz23NkJViufB/bNq7
N1zIBxVi5Inh0plvc+C9VdRqJFFtaiyymlPd0pfeEdT77Hey9Zm0JSMQyNCeu3zJ54G5xnopMWBW
nQxIsjIQx2c4fuMIuPAz/mDGqAQXk1H3ZioO9ZoxeL5PZkXdJt5TPOGWk7/PVgAXCwllnfTSPIYt
ov08HOR3CqOfNA0M5dM/tqmG6HnUpUzRo8FVT2v7XMhzbSEG5rSgMy6ZZqXHi2jdwX+9OBgh5Cr5
NRqqQwH1sKTmmnr5KCEiVvVi5AkkMMvCIfeJzzHpY7PZY/u51Vc6uH7ll8JmiHmtRPxWW57ZFKs3
jp8Yj6exrUHZH4VCjvDWtp8rPMqJ601DKfUD+YYm1mC8xiRvieDC3UpDtlIiP447DhZvB3jXEwyk
MUaslONS3NgZcf2LRHAFA/4CGByhSsWmDLRDhAmwS7j4lL1qWMet/EyyG33he7BwXiJgrqzPnKzp
PQXajqhyZqatK5suiuA6zN2GR2lVhnDv4odIxUgLjcBvYg6J1SSwly3CRhRUe7h5S1NHIHw6jcWQ
zOpTVkLzBcaOHv/l4N/FTnmuf9Hmc+IHWk2fC2ZgHMJ7MsvPoOBVA2XPkhVEC3cln3Z3pK90g5ld
1sFxX4OEB4kqtgSc4QnWG5hurFfZZWns+tLURWPx1OkohFaf15Dy5gsInrrlorQ8keAedPLXqv6U
2AQy4dzDNQ5gM1qOklwC7MQRsVq9rA86IZmgKaMMdXHskzRS894IE68mEqJtbR3zOj5B1KY9Ow6c
XnEDncNB/cu4WEQ/P7e2sAy7HGYrmRoedlXwNA7laq9JG0H2oCl/mxpYzkMLcnQRGGrAgADurZT2
9kgWpSbKYv2zHy17zlMKyRfaODjk25Zs8ItlK0OddzEt6vRESSyaM5ElLqogm77MWyRFGe8CJAAk
cEJsHTCuGj9L+rId1gqTrF99qXQ8c6xtZdNjcMkvVneeDCjYYUPWCjBpcClSgQcYe1iYVsGfb1ZY
IvNSjtuhegkQodLtdyLANpr26yybCng9iEXDb2lS6IJdLjRm82PQ3pEFVcYHDo3ONuYMhHPEB89r
Rp/EPoCuny3e9oiIQR8xDeRvxIiHxdFdPE6Q0994lobtlBdSNi+awBZFsJ7AGZugU35xqpwXPphW
ig4/0/P1NwKQWNF0uuad35HdIK8a2j7OljkQUK3igwAwb7qkQ3YSlTHJ7K9hRH1wwRZfFNZcKRMH
u1gkgphBldmT2TOVAiU9h1Ffq0p+3t9B41G93Y8WfOGVPCf7p07P8pAbPtHCV0Pp3WAuH7G9NmJ9
lTm8D6Z4kcLsRaAvWjcBkN7cxFFS/5um/U3q2a+3qIqd7aTuVxDL/8aZAL6kz07WiihK3XbcL3mz
y0c3+YiFpPCvrh2EcBt62wegMnpjRkdHCBTOn4Hl21bsO4QLupnaEyKh/8gxm0O2tGArlgKFf3i0
RUWf/PUx3SX5M8GtRA1/TXz3UtpjZwqw+3HbaCD4woHx/W2W8d09iATnAkN9Na36cKvrmleEFnQD
7EYgFqoSlagraqzIsIeId/ZlUQM/978RRe36kqLIJ16JUm00uUL0CxBZ6VCnEPn4AIWWtvhvLkQh
IYN97j4lrUBD2fO2N0NoYaccKrOm0InjGFa7LTi839lXaKk+ArptSb/pR66jlV2OeWR/adUGNTyT
qaZW/z7ylWh4uMWebDabSG8V7rA/Gyii5Esw2PLz3k3PfrHuF70lLPWfZL5PzkA8uHxjR2LUHA2B
v/FXnhyKwmsK+kXhW1Y7KkgOCW9cQGbQZuEFMJzcxM8Q+sDiNzURFiR9FBVh3FP39IDUQOHclkA8
qyOgGOg+FTypru4mx1hrebw51fgfAbi+RT3jZEoGOP74psOTERGmyYpO7yW20A7S3uyMeqicUFs5
v0tqPtl3X0xKf9BEc4oEs8/EwR+iCKrX1ln2KXHN/xOLVT8d6aMh/WrvGLJ/gCqsAnADI9LuodGp
g2QeXOJXSIwOoW2GjxoP9EKTI21fz4Phg6Tq1qqHo3bnITfFZ7xWtAaF0xX+6O0otvCiRRirxy1Y
po8AV8B038cLQTHCZE28g4nkRfPd6DPjmczz4jH1TkbpU2KWwSwNOD+8d1CG3JbGV62aF8P4XNb1
uGJgjGWSczuoLiv8L7az9izrt1LXJSuaRrOfMfXPUb/Tjmy95Cl+a+MK3DtNxUnpJZafrwy5fap8
wtdRZqiHWlVhXcdtmNkTgQgPcwI/51fJ3JNcKENY7GFXtabM/gEbQNa/CaWWibOs5OUOAILju3TX
WWEoiOU4SBv+WJQP/j+fzs7abLYwEpULjjisHdKf28lLWb+JGph5ggH2DcRD6SbyTB/QHBi6QFf5
PTzWPQkVS3mhF5ZSCa6wv1X20RsnESCJPG4sxj6wesDhioResAwm3ak/SqnPqGf3XuGmGKkmSqix
oby4zL4bEEYl91Ss7tUqIrYlhN4/QV6FjLKAG0p+8QF9eKCH1lngP0pd9cxBZB42FhhmspGfL2Tm
Q8pzJFT56U7HOAfnOJOXbHoVUsx65KJIz8mLbvu2k6aUOm9jCFKyCoGbAX4eKpHn9farEg5SMXXA
MMaGik4y9IrnuGGryT+w9uvOTx1zoyjN/PkUiW+0FXQM5DP38puvoEe2bXfMg8xyG/ga0KQVTp3Z
oXVC7339Xv0JI+FYhSJ7A3Auom4zrVeOcJQqBYkQg4A6nvXlxdMBsSa1N1czw8TuERRUiMxTVD1u
YHme+gFWYdQd5EqYIt+lxGbf/suOCoPqoth0TytKLHl2siJyjajn62pfVoUFKgXO5yfHujpcrC4l
2LJI76HKDvhjrdpi7TjEEfnLBVftCnrYvC+U78vPPTalw8til44xXMzfGf2t8w7BKPCH1hpH7Mmu
kXVfc8VyCdDW/rbrhZxSpzK5tP1Y3lm6XYVp4VchWZ9EgLPH/CB4TwWVHIPKCQ3tp2+PXOVUQZQb
Rnu4EocB4VPxI5eb0tSjXqC8xoRM1ePzmDpbWbFmT7LBar52Wc2a///Xc7d74doZNW/FnfGNGrWv
bcPyA/+F1+/15+o0+CkCo0AHm/qoqV7BKaryMQ5xLL4H8FjXKJytt9kaef4e2lhn0uU8Sy9ZHDxS
srAYHGiqcLu+pFNJ6XYJRgV61+cBJP8/x0vp/rlm+FGofBf/D4UlG4T7dOmeIYjxvk+yKHSorAui
ltyBosSo4uXLd2BS/qD29YR+75gPeDvf71R9zSRFQBAi9Np7LkG3zrE/aBjea+q+NEJnJlnLJAUJ
EqapiGzw/LgFGBTxi94U+V4D8gy0DR/fEOBAZMcuBLb72a5aesP6vHt9XtVGsQmh9UWEHF5EgEux
6OWm9yOKFoQMDOKHwR8U0mcl64hr/HZ0+YhnrFnEF6eMgqxMZzuLItkzmrtvKmeKXRhT8WDcHTyf
f53G3tnG+rITh5vqLFihzJbEUYMEEZgRLkoXjg1ox4CFnc9LjbbaEcJIBqCJaU0DTNVKUqQVdgP7
+OFCgZgU1/qSnHf0SoH71CLzGPHXPNCSrBWln2KQGlHEt8z8egRymuKxkJUOfJR2QNrOdmoy5rE+
Bsrx3R7rzS5fBL07bg+sQVqTxxeW4myoHsXQDSYf8SWOpiZCvjPhnVVKEl6zE+iQwuyUtd3AjYt4
F2dxWcnC2I105ZaSG136ZxjoGdWFauZr0mSolFHvPA3M8V/v6m70tkmK8ViO1rwq0xCEqGmZgtiO
/vk7ykCkux64eLaCS9gUdxNiBRkLJHRov04YgEPezL7Tr7OplRui+wTXlqk2LIDhmElQHGBsgfmS
u6aEVtvvGdXGJdywS44i0fzMVxaNotuANlJOtQlOsGJ6Vh7UWtJgwXVUX3th8vaKpyUj6/dprJ7u
OnMpecK4R5LAl0lPbmewOVyfXdHQAqAme09wSd9uoXKkWSy46Ud2g+iETLy2237Q3IhfZWKDI1+q
FuLj3bW87gbaW7faKfd5MJj+1YKVNUY5xb/aEEqiLU7khWbHTgbZruHG3pZv2LhifaYxkZu69seY
LVOeBEueHBbAAHt9H0c9Yau47oVZNbZoQN1jTg1ButHZ9BpE+w7u0PPADNJfLZAt1ir/zF3HxTTz
rW8ZmsbvFq8ajZRHJXNucy+Rf6AD9VIxLUVp/t5nnScpeQsHUIeF4OHI6X3BjBKMTGcRY0WhrV9I
dV1DxcB67w3Nb2oB4Ouhtlv62UBX3XpItQGp8O0B0/z1uqQ2mPPJnxXnPwf88voiELT/J6gtmokr
TegLQoeXv4OGdfyfFlnbr1YQoGTPIp6ji2dbOjg3EX+DD+BKfXXfWKoAzjsqYHlvCH5Ny0y82d6O
jzHFHngg2vP+eik7dKBce6IRnV/ZqgM3v4hwyFJZ8h55uppfTBgxfsm12sgVGF3f2Q5rcOnXvNtZ
HWkzKtvYdmc/hXmOs02C4r1g933+j279HSiYyhuoNc1ifKNtxXTPm4rCjTQRKUca/H82cKmzbgjz
HVYjlpGHLF09F0+Zb+QaFyzY9Y/EuWzMpupecPE6slWgql0oQRjR1+h/rwtJRdGEfXJyDq76y6z7
Xda2CbQPxPUYCaEjjn7LxLAHctmVA3eRrbGE/AEEtnPxF2KKxRecXwudDLMU8D5mWT5ThPmU2crg
sHVYPmbuMZUsb9i4rcqGlOBSMGl2UuNmp8rjsMphUwElBP/I7eFNX3tG9Kl9gIteSJvvEnefqPUU
lOiwooD66n2+4HF/+uso34HtqnzzTDrItvr3nm7DYKN0YzXWrydUMJAIZAbYWybzeVKvRo5Z320m
9p9Za4WTCPCUDWAowas0qkqKWVdte8aiA7xUjfjHAUghxa58k9nCUDXUAvosU2EIS+iETA8EkzAx
SgLhZHYqrB8npMcZrd9jZzu2p9weyUO0bfS3zaDhdxpV7R6zQpEnmr8SD0zraIHlMrIp4jSkR8dU
cNNAJDu+tlwcOqnQTMgIbHKb8k/gUOhZXhEvWkq1mWWbI8c2mkd0uoRe55QlCEmLsS852IDppaCF
i9y3OlUlWpFwUfcUNTHlE3B5JbZmnXoHoMC2+pspMqWx08Qv+WXsBmmoCWaBeIHYc8p/Q4IUXELu
NzPS6Afzgf9DmOIolLZlNQDEa2nJdiP72zbeLcUa11M+aAQRFDdFNP+5ax9Mj5Eg6KIUbQN0R/ts
oLOY0a77yUgVEYQ1CHSpx9qGPbzK1BhKwREBixzcSjt8latlVqL6m89jOqAq1Db69C9V+IFrsS0J
irm+uAekaAA2wLXLX0t90OlO/nA968BEEhUDORAN78fGniUgoIquNoseg63kUDM6UVBIkWLu5qto
yf3WoI/lSYECbGxaACwzkdXjM2qmJlLX3mJiNODK8t23DhUSwdPxL8rHwUREq1qcLQtvUq7V1ule
BwCG5kECIyiuNJkhEA+unANJhLw/XEy92tTZugK50Ms/79o2HgBGnq8KLBECOeAolFSGElMuxx9d
Hr8N+6vLE3RUkY/w+vHcX65JCRbjFj0xENpuqf6Cu3RufULuQxx5UEYc1t1VqJ22NCyTSVotJgL/
qNkCwPqre5q0b+6/IMw8cBKpEEZtOGhLFxd5UPqdaE8pms1Atct43l2UL4w3CoMV+d7RtxDEIHkJ
WBA5UE9lj8ulZZ+lderFOyYEn/zIVDAVhlH/xYxS/MIHkrlK1AJRNGkaR2LtJDTAkTbmOBRpR8t9
s8oO62IDMfs51vFVUNQHtS6v85zDavoWoXHzhWDE3pVP2GKk6RP0qMZJb4gvp0U4y4aiPLeb9LPx
rObdxcYBnm6jxg9tiYo8gZc9qkgN/Li39GyAU6G+S7zuBtdfEyfvPFIE5aM3dn+hvCbDPs2wFEvD
4fon/Pm/PvMizfCEeiUiFoX5F22Qw+1utmKMRIgN4CufEzoTuQgnI/kwMRs+iIbNxtp6/wogAWAM
FnRR+trSpyB6gz62OLgpb+JJm6XKJtY4EKVeEqst6b0NlwdYSJya57raRFIdtQeYm6Rl4k1NJ4uN
fht6Kmmb2Ss1+vlSpKnuKoYR7fSWxA+7smucoco2SLDEf/j8Sol7snU7A8QNSoLcQeRHigs9Qub/
yWqsg+dlOPdh0C6qUHanLMuTRnfIP3VXNHEo/kFFLPHk8aoZX5GRT4ZjPCZci6mj9f2k3Xsk+4VN
cMvLC3ZaPQBKHuKhV02+tBtsws0IEM/DjnPYh6skroqwh0J5QDhiGoWB/A3WVvrGrde4bHFbQlwr
GJTCGSWOhjW213bqFTRWtQGfLYYne/+VsS3xykLLlxJiYoB6y4OLFUkQ5sZxSA5dNrmYQdXUlgPk
BTjfLBK6ruXAaQifvBWb3dMlvsY/owfnXApSRlhVLe39jpuSr5lnllKYVhZncyJGP2x4iffq1IYy
TrstvuAnsW4rlCLPy8WAH1eBA3RB4/G3IhQpAI+UKgxZVaAmRcc1/YWFClF1v7X8U/GXMfg5BVsb
Z4nXg9vxc5lREDbs3wKwFwEmZyLzrcc1m2HXZtGipMZbBXohel2x2MRvKYta5hQ+ZT1kr49cwxey
xOOOzkAVHQF3dvjJRVsh7yEDtEH6nidsN02ivjftJnDvEBWgGM5zUZkmXjxDqnSWz9fvsARQacQS
Mcina329zWo38sO+d0e1MvEu2h98aYLhX2WpTRBKatpkioQVEXWYTkWRAiB8nf7iXIo8WX8n9ijQ
yxHXnHvVwQ7IpL6TYV3vwOKK9+spE9XizNLhWB6sCZwgqHt8YSoH8FdCmhUbP5iSh6dogf4NQjYM
MIqKH64QA5EefXJ5JbwOG/tu/kZxP7Xq842rzTLwLp5ga+G+UxBzPQwJYHKYDmGCqTu73v33klhg
zNw+oQoL1IOkds5XZDFc6GX6v0htMVXNDVMhrTyJ0L7rgfoPDJ9AmgT5U7arYfy6lQqGN3u2LnQo
qHTBuQ7vad9Q1BuLZIIQsZvyknTgRsEH/20tH2apF4GQ40X01Xv9y2VZGi+eFrCSkpSOXF+LKly3
LAJd6etoGpGSZAbNWpfGLZiA2QJz2D/gxXdwkw45C3PWBgv2Am8Fj2EcjpElXPoMZIy95PoxmWqG
l5ffqpGV4IOK8T+dns/ZvNfEAzU7dqrPFXvGpc6NGIyMWsOfiW80abAMkD6pAa5IbJek2oivPtsq
2hFnJzXv9TO2tEC4XjNbVBGCUhe7FCgUOBVewF7BkRCJDR+Fi+i8TPnrG7P9MrmBppHd1O+vF1pN
etJzcB/8+2h9EiTIbK8EHNKp3rkYVJDNFGi90Ncqh0TwcB0UONtWlXWKSsLmQgJsWr9AGE/x3iZE
rPztiFKCKdr3Lt086yPRB1Vfq+jh9U7I+c9Flg97VJdvjBKKkWxHopmPNu57zAAojPRRRfJQJPy8
0FWolN90+0HH2bm7lcH2FLv/eXr+MwhZGtgUybnUbqW1wwVvb58aIUc4Kpnp/8fjI+JRy3pfx2t9
xyQ1lJrIi9iQb2r99kD5UhY93IwHKPWn/rFMYWt8+UeTlxHmJRk9JBwI19bMlCZJrbrcMaat3Erp
VEntd6qfJkT0K6+dtE+xSmDE8TW3NyKDJtNbDGGkbutOJ8nknTrhbDRDODXy388C9k6Qmv4vBn02
q7+sN4oJNv6PTTF64dIYoXh88CJdeDLFheJZAgWw3XFlfnB61lGVnV3b/K/qFeTLsBhuaQa4DSTv
EGx5gpTxEoMYb+0RWL4TBtZHX6717Hyal80fkiXQhUcpIJMg+QR3GfAVrp/qwKbVaB/tfDR3XwaX
YbuTAc4o/ZdgiXzaGIiyRQgetLqf+EfdL5ZuWT1GA6CT6RLXM2Oxr4jvuVTQlQXWq4ShzsbD2jKY
jsArcgxybatRZNXCmQManHhBZpjqQPrjghbqHS/ve61L8lSBECCRQOPbw0XtbHnQCRLJUdrIALjd
YEGSpENz1pd7sCNdf7BAIIa2B8EAACbtHFqov2QIF7eavPmxj8wZWZzpVuM7dj7/lhMybOK56BaD
T9wIfOJBx5EcmKsPXChZn48F+/COJ/fFJrIbhuh9sCYEt4M/pE3sYy0Y2eDC76jGdXErGffQ6DM3
hV6Xe2xNxqC74gBkfx+w80PwehFWosA83yV/KZC6pa5+iLSw6aeUMaTM2ZwiEIm5oFDR64zgaPYT
7qZ1UH+liUKuh4IOAITejjMUt26bqDccwGmOP8J44wHZuSK2OU5ZuID79WSTkeYas7DghwQzixtL
mO8yzPeTHVjLECiBnjj4gMMDuc9xoJLSghW8fo1EpxE/lOoDqfT4mdVIpcmTfbehafg5pIDs//vl
kltHCsuzACiSp5ROgNeblmyfKu1EAnckHtX4BRshgW3MW44mrLIfRv/yi3e/kp4CJI38MEXpdcmw
xgsarmZIYf+qcm2ZrJzowp/Bz+DirhTo9XIcLGxZegdLHesUcvX/dd3WgNS7BEylJ2HgptiKylO9
34RDXIRjwyXCcQgryZQI7CLr7KItTB/23g0KTrshBgZ/C67/lgGkRhnQCsUlI9SgPQ1dGM4VJwN1
KhKoXpeH1fqf/ELi+qIHu3xRYLt8cjw6ld5kvcWd4z/iF4WrFRrKw4lcsCqY+LaNL2lsEFuPSO0Z
8dPq0j8f5XylCuIr/31Y+rMD8t6ponCL+Fk2vjq3TARigJjh2rCjaNLBtR1Ni+e3W7j4aUVDvvjq
IqB0SniCOWdIW47TIGd5ZSzaV2yYRvsYDmKuj2GMOqeeWbENj+OCh4nHIN34tiswzQqHdLN6XLuK
TDi0gTuIkjAAutWhe52E2POh07wzb8esMR2YbLCfyM5oN1Qox5LQkWLHxqM8lyMIZy+rNDt5OB4+
ZWPL2LLMzW8dBCSirnWOpX6Hz1sZd3Shn5hH3sBlbknyOQg/g9LLiStq+Alp/+PSQueTBbTlJdho
uDbGxTOKmDQpIQCvl2Hmuv//LO/rK6MfQGA0cWou/oDcrQ9DEruJ8jjN9k1WI2wG1kexCHOMX4zg
GFDPCvieqtjzMy0qRMk4P0lug1FkpUpeTG9ZZi8Ml44c8AYyCcJ9nzHmFaXGLWTSxeoP0Ml10LRK
37o0sGP2gHEJAVf8HctHr7ud6uY0ZgqB7puBaHgb8V1eCf8BO5U22cPQOgrmH6w7ZFSgSGpxEl+l
dRXNEQaH3kjXEFGTI25t8hS6CUMQGauPYOmUxfHbM+0MlQUBRu7iqVLr5t4FvyKe+xLUGeEyNvHn
Z0C0logmLmQEPYUouF5Mq84Z9C1OLZlfZBt2LbFBxFzhInH5pySZZ41ptL9Vp4q9sNp9qv6p+sBY
F6OMHL5TRW9WQKKUXiC5rnCm0x/Q6esxN6KM07e/PxW180I0Su+x/1CO5Au9Lple0Rns4yoKFTPk
dSIX/WYUtS0Y4PLPzMIWVqtFLNp1zMjbQGhR1pU5TqLTPFSl0A8blSl1e2y8k/m37xiWZLgZnd9B
yGhrhhOh+6TCrqSbqbyp/IRpfa4Jtri9U6cvpmfQdA+bY6mXyor8Z1TdMgWURwXvAO+vXgd5AehU
fcEq0tW8u1byFhdGkpRllmRofdOKydyAOZPxRWhDqfRueQioZO00fK3udUFuAGLVlOhlo2BgoXgA
AMYMLwZ0AcpDVbXrNMzZyJ9PLcDxdZswbAUDLuG88pB290//nCx7QL7EsJirdtl93uMqycbHPbMv
3Rk2uyIw2M0QxRFpd85ZV13na0Q0Te1GSIZVmFC0Hduxg4VnDZ1yHlZzFO56WTnwU8xbdzc/GXNH
v9ssGNH1+4qJPfr2UCHnR9eKBimvgfLu1z2t+HamO6y/IbFERn8ertlWjaTyk5rafiIbwvv96KBw
tdMtTjRdE0XFlPuAj97f6/TSp+tFKFw4YgesKk8ExRPOu7LlUBWz/s5VWm22l8lf9ZfyqfqHc/m9
Wnx1JZrb/7cRGkP2kYZGI5h6YsHpjOwBIKQ6vgIIrTh8wAHXKodkMTkOGP+09xEHJIjUBMH2vFWK
rqak1/Qyaj3Xyrwdg1tjLmLX+Dsppg6ukei4ics21iLPPTGByHNpcsuNZ0Z52feg05ZqHWcxyAlH
eSyvsWwEHEyUuU9hMvIHn1aoVkzl9nr4HVRec//eThUBMmAs9v6OCnyV1wKP5Vs/APFGK2v5oVC/
tzzaE0oChwaHB/vTnvjeSl9myNOkLj/XhDz3IdipBLYKC3HmY/2D+0yBbqPKXjZXI4S0lsbnwdB7
u+KeCq7ger0Op2Ej5EURk4bUCw9ke2/8FnuLCXTVJXiiX/xxDMwb4PpIH9BTQUtA9IMZnIKvPJuw
rP5ubDuuQrzSwPk83UiojSOpaBzhiZL02/O2s2VXhir1JwmZXCeRWui4UCLC0I5AJQcBMGIwgbTb
OXe59ukHNG0PjLLIFtzbhsXvCu6hzmNhVB6HGVRodNaqsu+4httF1P13ExhyxRfXjxdIGE2ySX7b
xLFiJ0Io7NLB2WJEWKyLt0PGJu7sJ5LH3wEydi2BxWP1zlhTEc8zJ7s9BqopUgqbvS/SJhUIAlcH
LDz/9TU9aGhcwwoV2N7crBKMRCWK7f3GqMDICViYpNsJyaRu4ENH1yNphCh7ZTSNgJh2qal8qoO9
eHl97ZOl8NhGxyceZI4JPfn/Oa64F1mlsusXclXzpxgyBZCKjdCZCKcu61ShEOqL6hLvVQjx6lz2
lHxSEMEnawW0+npv0xWCz9gXrcyfFwkTu6VZkQ7HEYySdMGwdbnk0sOyHhxgPJbC3lpRK8zMLPGt
YOcust3KOV1X7M9Zo7y49pMi6B0xGL7z8wFV3VKEn3w3BZDMQts5IhLCs/lQya4SBEob4Y9J19yj
oH2plw+OYifc1N4bDvbde+PHTh7RuJiLs81Xm6j9BCntoMZCwsh4KAqBhmd/uZmRq6XSfWkMrKF1
U6h6oJqZufsGlOo6O8YC3c+X7B8PLnp3dot+rUqUOWoE4skbcYbjBbFJNfFnHC+PRXt8NADh4rNL
Ccqyl2xASNGk/PT8nRf178MRdzvAq9fWXXWSo17DAFsPQKpqCOrFSuCY+d4KWVp9gHR20vl5Vydf
jNZta+0ZbCElMpf8rAuNPn+gNR36odWK/Oyf5ACfRYzAn+q4rloeU/Iz0zB25xdFOEwuK3iNpmxD
8AjEFKn0JKcDSMIRGM5tuQ1eMz5MTWhXFiRiuclbGTumo0PewX5yxzMRiSLSm6ZpPRNgidynxTwg
Qf2/+7Gijd2PN7abYc89jQ2uHAjKA3ttQe85za4BrRzaQKm4YaONaiSg5Fy4Kc5PInmJrytfu7vH
hoNjsoLG98adjMPgglcmxGo+a4JW4hts9Xbb1vP8ekehgv2iVvLnK6A3uqQQGIEspiUAc/sjB6Sz
1qYIN+qfLtWGt7ueZKaApE60v6GuZypio47RF2tf1maSxeVH/S54M6iT1Y+JUzpZuI0lY+UdMjSo
Q/pLBaaB1W7cJK4p2HzV9Qh1YY69Iq89nH0+cFu80KTKDD1AyHZR6LYB6WW4i39LP3kM2Ns77av+
SXJXXE1Ag7iq+WWvZgCBIhgB65LofhJgZ68p1BKkfMO3KI021JA9b1YGQlDC5mfy/oWfbvzhOiM2
sahbVUdmzFrp/h6eWIhqOO2FC35nZvtEYgIW0V61xuoffZWbVelE6kT10h6YXXeiT7eqiyCLSsT2
PZyI8wVroJgvYOe5WNqrNgxq1vb/0op5AXDoRYPW8LMPcaHbs4b94Wq+ouXOUK1aYNEromAhEKp9
QlaADTQz0wFfiDC3OVAJSyV/t/jjAnAxDDooI1aqF7DGr3gAmaVDhb2v2iZnKTSupbtnXH8+XdX1
z+YPe/8ZJVzesCGXkZG1RFLNtSgYTm57XxcTx2gMAGTb9rsJHyGHNc1mxPGNFPX+7eQVCYWDN+jF
wy+VZOOr7UBg5ma4Q4U5iytXv+PpXs50jHYck07TTTwgb9DkdtVMFigpRVMeq3fKVgQN6lU1rVfp
pKz8PPKfWnP3sDV5zNvSoAoOvxG5PhDPA5NJm/WCMhXLKCInTF+aRUR7ozUAE5CddZOXvOnV9Uyu
EkvYhdKmOQ1gFHZQYWHplcvUvVVmI7Ccd/axkCmvamQP3cCXk1Shvoft7LWtUB3EbcP5FZ6a/1St
QSOjfM2dKLONdyc2vKnCLwht29w+zR/63jnB6aOzK3kgEeZBwcn88Dg5Pd/HYaaV8zQj70L6R7uZ
T/tn2U2GIFOCz1KH8om1ytawMyo3y2r7ZV568wZWu3F+g6mYgL1r6Gz6c4jalL3wcmYPy+4lczt3
zuC6toskOBythmUC2IQoSsRHXjsMfR2qbhKmv9qEvvALN7Qo1DrimxZynfDMjQKKm1jVgsyRnF7t
HaMLqNbmsEU++o8vv7TNrkTX7JYMKAfYP4WBBx3vt9L+wBRV/rhhOJ59PXFV53mS9dkbzlV4yA1R
XxlU8+mYZyTdjK9CAyRGGyYzFC/83kdz8tJlE22QHfigu5+XZw69KdG50eXqtLdX3zcfEMMKBiyy
z9fWcLyQ9FIDcZ+Z1LjazQKyIzloSgCbbVHGGseICr988Si7VDe0SYE+CMR5O388ns/VIOeAz3Gy
U1uqn4Wu1cJ26mIMFGBOlRtUbeOTfSR75IUZloJy+4NLs7EwuTll1+eaOLWrudq+01AU1OUwMVO9
qSWzYEVdIJ/L5jH9q6vRTTRseKbrzrQb5zTipqGW+IM6S1m5B2W4BXOa9FoLQ//VZ8xEPQkmBDOl
CqKVK5W5V3FzWyxgshikvZhW2SL0LoYfEgOFIThL9SkAeNLkCQEJjW6GztVxQ5GazyyqW5yYhE4j
0T4SsOZt3cCzShZVVMDJJw7HlPSwjM6NfCJ917+ibaFVG2y+Z00aA361Y1+fVYwooxtWcZv4tFEk
fwN2Prqu0A1m5EyqpemQcFvnZwClOF/M+f6XMSurUiow1LvxadskBsGS95OTmRNlgCU6Eq9ZKbwe
7TT3hWBEWcIWRdDf0yfFEirNGIcvNHkzYQ7yplorYuzo4thKEyioXjqR3NGAX4wJ3vLAgmtkQEr4
8bxsVaQT8hCRbFTd+LNvWCAh9qJo3bigpdY1yO47alZwyj6rh+SpsOZEpQTvkUyMcJJT3heQVMiy
telhxVq/Dorup+xvDP9lU3Ir0HcEWJNknW+YwR+ACN4V45Z4ScOeMJFzB4AbctDNGrjzTP4FngK5
BLv50a1wK7CNO72k6DxCcX6Hr6kSMspCJK5f4RVUStIWSHnlR154TSd4M3yZ1a7i7SV1QHHI4k8v
r//Swz8JRQcVQgoQxoVE1zwpa6ykUiHciogX45a0CmUHZURAU+m/Qt1DEO7Ismq/7jfsjktrxkS0
MCpI9tJyKUktX2k5zMyluxAZ5DQ7ztvtBsiTmiB4sQ82wi89sl8W6nxeybCNcP0tdHiHyOw/06uJ
imLfVvSLfN1no905DHjrV8+W/veyOW75uTt1mefyCUz1ZTtaUeryGx6633kadwYkRvIom/myDUPd
gcU8u+tRrYZZdX5ooKnIN/AjaM1y0M3g3QASl5SX3tB/87xm0gx763ro1Ela0pbzN8zmbkpJd4EB
oss0vuUifRqEpC4e1l6sEMm9RYAgOokmBM2Uswj4fa3QUiR6Q9ehtTZysufOou6bak6OoDgsvQUe
8tZeenO/lhoIlNA8Wc6Cgc0yuldBLwSQFFMBZRTCN/ZIrrrD+CfLJbyT7GTUceLcV9MFbwUJ8PE0
R2FpxjEJb8QDBmJg1H5oKmotjonefpcxHzVDOkUW1jFE6h/SQSKllcx5E9MILfnefGAita4CW8wi
5yl0pDy9FKCtNHRu1hmqLBAWl2x5HRQI30iDnyXY6gN1mltGPsPcWMkWV4yrKZUXmZUnyyly0VbF
JxOu4hJwIQH0FiJwkSfqMlGmg4FBGBkwrkNxOshuXxSO/TKChF6+0tdOWPamE2R8+ItusNrqcYQ/
ajXXUoGifMPhNjzVkQgMwq2m0HCgB3K0sMMDx270WHJPUaXE2wJgh+rwbDNreZoGuCqGWdLof7FD
bNA7n0qkKj1wvhpzUU6RxwpTDN7UyDVZrsZNnyPWjaJWFGSA2xB5UgL87sUkZuZ1WjJH88XwG4QD
xUtKzvpgYpIjb6sHHiZFNGHCrWcTRy1dtxLUQQTbviDJmpYpinW7sZdn5Kmc3/lKiPXNmPBWCb7Y
zY9mN5BVGbB3DrLhqIv6FEz+NUqEXf+8YTIwtzhLeIo7DuPWDWu/nqFvvRgtG6KmKhzA9lCWZL96
unpVKCxgtHdmGLQfsHjkbho7EITGRj6WRzLDwYXVfugrLALqk5S/lhWqxUtI80tTcigeZ9qhfOdn
BAWwdqmuvtHnwm/NVoMWOag0ha0iTDp4/rVMkGWVwknwslq+IMYmJ0JrhnS3TVV90owTa/dK+zTD
4xo1zdW25jGfQLT2HGab4NE4OZ478sHPKE5M0zUKpqBkzFi+Y/hYmaGwGtnpbkcrcRFn96pzdJ6P
mo2nYQKWPOD4Z/SiGUCkKd7PzG3tSi39ydT9fDVSEhx3/nUS/PkiHRh0bliHpJ17KVK2LIpKNoLK
h2Cy6wTeCAIaAlxVMb1cup8s24QdYn7y7hsM3+EacRdQE+t8/zsv7dhxENQLD0IZ6JpRbE0QjV/Z
QTh6++7/5zWF3Aj1UQE+5yxM/NVy64HZ5wiQNp2TrBd7GLlgpaV2zSchdNyYRXEMF6GbemOpf+zy
W0GB58TkDiuuwrUBXhT9Ns2PW6+D4X/8Ex/MQYdVW4mUW0UOFCGTVlzVyu2ziypHydNoQVU/ChmP
8RPCcrhqhiXHXCH8wkUepZp8ztGg7RZXjza8zBkWmGrZun9ZD1TZivDAtFbzsVgBDww/FHrVUykf
Ek29aI/Z9Url0pochVJKKbju3zar0vwUXWdYbvs4R7hPQhRG+ZXq5bRrH8ek1Kw5jM+4LXkiSfgo
Sa2Obc46sPkZKHFNb3V0FKg5NZ8E69JrGjcLaAS0Oeko89o6eN+RqeZ6QtRN0d7WVf4EqczcpssI
/Mdj/BCc/rlrMa8Aa+QVQk5AkgWHTZWFxpVl2GkudvI+I1ccpMbeQHxLBuuD8Q0V6LsFmFh8afl+
KwTpAgH5z8sGwz90PG5xysMauMxp7SC24fAJfd4DjOXDekkMOXSl5Qljs77ENKf2VSPFynv+04Go
jbLnjWRlIGY5T/rbLqH7WEi6Ua8iaJSp9BaE/VU9wCQ6MdtyyHD1gWudDGDjL+P4kQbiZkLZHI7j
WHX6qElPj6EgXMTMPoGQfyum11YxKobQAkt0/JkhNwU1dX6+I9zNunlWl5ayb5zFKpsWhJCGXHNP
gc/kN9pcmx2TMa/rAaaj4NPowBC35dxjS+Bx0oVnn4VS756JmSP4MHwAWuLHPzGKEDxt5xkTAgjm
wwDruWrWzaLKf6J3/VzPyCVaul5zkT7ye8TuoKcCyc6mwRB25gIucPvG/FgkbfAJz6cWieCOsvqt
2XwjciMOIniN6iwo17HNLnqWiihf3dp+rQKnIKSfpsUpOTLqXVGiGXWhXO9xZh54ijywknZ1Ed1w
82OgQdYlNmtKBEpMhZd2hQq2+90olzLlrDQWCcUOPDACCQKRLYT1G5AlgPBF9XeUNQ7LAZ43ubLh
AKijWd7k+Q4U+IRaXqVn/+zek5euthKuRsdXaxTfwCW5VYUj6niInsmgDLBC0YtegkfFvqam878W
Nx9hxx9qrcMG9kNvlsM/50SqYKFrOdV3fNNKaG6bz0c0rwHLWdn1numutqTdy78KxvalElvYQrJQ
29jleRX3Y2GCwGh7WO8Hh9IJ5yZz/7JeYf7HHGVC4pkWuYE39faCV0SdAeRQ3xVgRvFcKdugCX+K
SnQ+xQU9h4A+5E9YNjpxwo+5ozvelQoWE0PUz39SvLLByMaWWoeg5DTFDTlh3zGYOlhkZPlSUou6
hoaPQN0Rt78/W7GVT4h0QM5lur1U9/JfH54+Ik8XwtyxZQDD4dm/dEqCKx+RlYkF9lnqd4jSJPGf
6ikBeQmuQ/9yUM5NufST+Q5YG+zVk4iH8gEBx00un8J/xaTSj7jQUvcwd359Bk5FextwrSPSIWFb
CutNIQBxRfTk4URbXzKfA5X+kV4ecmq+WKg/F7oX7wjvSpNLQCqd4b/2jEHaAxXbFXGCNSDDchXr
2RRnCwe8TeAhHXptlmxXaeHcFc/Xanc37r4afrahmKKHe1gnhMi+++mA6ZaeSmn7Q8ZTUtZCsfxd
h61F8Z5327VRIyHRMTRm6mKWbZYYf/AZIewqwJc/SpWwdgc+9S7JIospITR+JzHaNbP6NC3NTF0y
BjhF2XG9fwCsYXM7iR/WiTj8PtflZ2CEL5SVwAP+FOPQaSE9cVfvhnYyuNNMOSIfno5BhtKVgvN4
vsMHy5faX4trMElI82UBYVgbAgTWTmFaodRWmkPOUZ71U/9aZ5gvweQJJSme1vxYNsUkzoeKfExm
JLChvcj99Zwt0cRKEZ9PKSr57i9R5/la0GEtS7axoghIdNn7QKvfQqhaujAUFvfBZq5TWQnFGT5c
koLbNuAd3CKRydq9KG1zOr+5nraX4bEGEv4h0FYDF4VxRpocWHvHjyI0msjLXjEloc/nSSJwmXMR
PP0D0ORpmNqF6VUDqyhFzBTNgCyv8iRZfx1zS+6XGvWvFpHb6MyiyQ2KgjYDhSC8NEZPJIk5z9P2
0sONv/UcUOKeoEjUzDEkTog4bF6s9l3qRTaTwV13FrjiiPmzrdo/FPEFgNgMreZ57HtPy7XzAzNb
IOJ7umxgy0INhxoTUu6BamUibuYNvVKWJ61IIlRjbopHNFh+v2RWJmq/S1YV1ng5m5Otnk6zU7JQ
ggFR10h49uOO7o95KPNbnHNE03YGJhP6IcLwo8HbnFICJQHwRpEURFeN8WK1Ckvf8ac+44W+1I4z
xnE5w2cXwE62lSieZuFQmOXFnFP3R0Ya9NPqNnHgGSQu1tA7XKLss9s5q6jK8ImSgmrFcwlIQJy9
KQCx0b5RHXXbCdugF4by3+wa0atvFbIkc9p97yna9tbFtrYhYmVCzgnaRGhDmchu0KTMvBRxepCh
AtI9e4yEfHHQmnOUUJJHlDn6Fk0V3h3N7TRkWO+AwslRPuLHOQihUwr4ASaAJgWejamCtgkuwXu0
pWBEFN18KpLQIIPIIMBxUZWwidZGw+X3BECfwpS/8n9inW3rm34N3JsaKndmDDJ9UbEjsu7/ugkH
91qJP10UhU+n3xfrq3gjIMs7MLPxCO/BA3nyAHlOwiFnBJ7w5g9+LuAw+nvWOWDT/yaNlIYXDnAk
XKmVUx8p8UdsE+UZU7NO5fAThcYSRs7PuUrU/HePUcj/8d6skPJR0xQFSxPJnt2qyTgEPt2d1OB4
uTPz4z5l32Q4F2esMbSE1XenpxTYcfT3qSvoAI0egWUD7TQkysI8zsaNSbAxBFFEn+L1VQ7Aq4Xk
2HQ40/Y/6Ar1vumZ9Xv+P88Zq0dMDYTO607kX9OT5Ct3/VAvsD4lVOTk7KuYxt3om7PJrSlVOX0S
yf4ily8D/UU9tgjUFOd5JXOHpDN471bMkzq8C3kdgXs23l/DlKvRYbqpFiyixgzQ6ZYETxHycxxa
8kQLpTYFo6+Bo4yINL0ujdUBGOQAsdWKUUBwluLOJBjgKZHn6KSaCy8pwDJ2/feWYmJLGRWH5B03
wJD06neCb9ZxsEGyKmwCjMyyyxdMA4sQAy5DOaqM2A4dE+ijyWBZL+AbNdCI6ML6FKBS31t2zxwM
GH043a23AdCRnFxnJ29b5GPh6EyieqDqhuAhcR1B8IPrrEF3YIpiwLhkBcvI38b+nrlZNjC+yi0+
EHBdi9atueuE9EBfYaBa8w7eSoWVlztRC8SYBW1p7FUyHAHqECQWKnQ9M0CdI6BJISCqNh5Xyt1m
hu4FpgstdhSJQOdUZE9IPktmcgQD0/nX6wb0zXF/GCJtaoongSA+SSycvnseCxwccWaC8RPAW/Yz
6Au099yLabdwgo5NybSPeqJw24eS0eOw1NnpNh+CLfzJqz5SRiuZ2CC3epjL60axEZZ8EoGEU6cq
n7EbYJZoA6VMRdnYbyOcDi6AGAxMIEjvmnz4jLCSja3RxqKB8LgEvd3uqikXjwXnitkFo8xybczM
snYem2w1/7O16RciB4jgHly4FcUSfZtt1C99Vk7PoNvBi4hXhunCpH57qxcLqwtEarrpFYLuTEBn
yxy1EwEdIIPGLzrTTf/CRSQvymDavOmoG+vrvuRmWbflQodC01QpFeqR61aigOhI5fdM0pKBl8a4
6NRdGeLb8qBqpUSMa2kNbmwPxToZnpddZK8BgC2wnj8ALiUGTbmKL1+jDCmyRG1clPQK4AsTn4Pz
Dbdyf7S/doRbZFHx17DgeBy+nBXb51bQGAbeBkzrAZrLzCxVCjp2KSf22MmPhJjPQyCWCKrgl1lC
afElbiw76Iz6NNYO2Qqt41vRevF5Vpz52k/r4qpsKAom0v+j/S8CmRvnLYGJpctui5SBHif/kROZ
X9MCt2xw8H6E3Z51L8NJ8D7q80bLQGbaNzXLeK90ghCHSZyfgGReklMoBYAsnscpF+ye/a7Dq6xu
jHdPqzcjZcvZVkHnmNoGEZ1emw7FzRnvSGuPKz8qKv83CZh82rM03imdAyQkF87OPzaVF/HQ7CzB
n4fnhDTAshLpZFRFLHstXz5pt5J+R3+vXtjInk6uixk5guXNzXgw7K0KGYSsR0Iw0c+r+do6C/dC
l6IEfiPwV+lPNYZrhCCi9XiuLdDTIZE+P4Mp7YclXVcYC6z17tW+0i57OdY97FuPq2uUlHuUop/e
I6KseUWlOySOqP9T2eVfZgD0Ly5d3OmEby2+6mjBMnqKCQ9c+uy7np393FlbHVjDqwaCyya7ZqYa
PiD6wPlTW+S0koVoTjKX5WmjrGSnGYmxlk88ZW7u1hvgKQkpDKe2Dsx1Um5dSj3aNf1sAOOH3q/5
cszZlnmM571wt8e8AxxCMY2YUL6xXOuCFimSQCdGe5qUeVCD/J8+KuP6I7mHruBSK+QOokQVHBFS
8PhPVROOwBXQQdCTRZHcxu69Arxtgn8kTg9DYw3hGdfx5WWdEQyY/FoQUjcP8tc0pcBlSGLveZ0Y
z+pcOerGiPxallOzDxeKysMW0m2fQ7F5sNBOXqS5ZYfIBv/VVYZNm47Sr6qUklJOU7ijUa5bNUzK
YzYkUFuz4x1o19H0WVjNCgqUc/t0CSSJ6TmLJYzfzR77j5o/6ip91+GmEKZhmb22kTxdFg5e3tZT
vbBePRiVXsbuBpOSce46oh1xUW3wsCW1h0N1foKXx2Zm+gago9ROVf8ytan6I/Zhgm7NTATa3OGB
A5jFcd/yLaZHSZmSb/QUR5ldTHAoifJ+ykLC66a38r4FFZWegdj02yZdftVF5naoWtXJ/td5VHk7
zKXKAQWusGcni1St0UI6c4yGw1kGuxe21KClkjFFe1RmvkgL18WtLZmDGl9TitrO/ioXtWk/TFfX
pJMi6U8h62Upr/7XeQgKhZqMXPdiMwZbdHlOvvgX+cO0dVfx/0Fs4foPcyWYE1svr2C3Z8c1Pc3X
1Fk5qIT4X9kSko+tbhpiKCPktbWIMZJhKxKy690tm4DukxdI+Rc2ws05ZaI9M6ogIfgcdbxxCyHq
jdiNEN1FePaKftL0rrAbILEj+qyHPZRbSZ5zJaaMtU9CH23fUlhazfHPBIg5mjy2B/wgVMQj0fLe
Nq5cuqSF5ggVAp6dCUWb8SKFQK1UnTvMANahdFD6hxL2VU0d/VuOPRMnHDImoUwp8KQYwctJPGTa
nJivGVzpqcOiENx0dd/0C3RND/11ktqugYT4SOtZkFW5CHF9aQfpre3eTHHADE1A85TPxBOR2Tdq
sHdmFPruLi0nSPFTC7CNdMDZAzRjwpdKtFEy3NXKWN6XemrXSXtS0OX5O7TDKjOk+yoWs/58j3je
uvH6I8JmP4WqbhX4zonknAZUbteEjLa7lh3Zig6fKm9BgasZ8LKsAEknxFXUfvpf8M8BD/8NAuiL
njuI/KGACCrBnmiOvPcf6iaKcDEstedtM8uE4Sj40Gg1MuB++Z7UNNkN8NLZG+Be5I/En7Eu9PEn
XextWCN/HUz94C1KyfFHQvw1TWh3Wcw7ZA253zVIdKbNy9VJ81ZkAit8SxF75f7QpBOh9/MJZE3f
1Ucb7kNbjqVfhEa8H9RatzyuDeo7WyqcjZLJvO6RdMOCpggq3fHxPn2jHwkMh4aq9aOPNtu9buXW
vaB2vLMFLdnlhE59MtG1y4ap3Dlhi55sQSPvp/0aT1aHYQKFH76J3XsKOVBz6b3GZXXPIo8lMeIv
3/rvsc2aOa4R2Btfhu98URr0dTOXlmcsYQUUid7wowFW+fGZ1jdHHNRjCUiLPwVDT7JWiUbhBoJI
RWQyWbcUGukrjugKhNfx1c292qwnkLADc84jw3Ce+t9tpdOgPBYfyC8pJjMSPKu+V6zWxPTtlg7E
ynqC/Twv/g8nZ3kyaUjLX8sGnbUPRMnRiNpkThfTEGwpB/4INSJr5N6TC7al4LOzaq5ExLl1Ih/Y
qn2BSJHGhAm2Xy/el7wQgiiUFya74YggD3ECHgXd4iO8cJpOk3+c43SpvDVR9Ie6kpe+ZaaHSerD
Yy1sCxxL0mOejafxD4AB2k+40ttZEgzS3X0QLPl7AtTx5excqMybWPFzr6NVI0Pjk4oo0/7isbxL
+mSYcU213BRkeIQ1Lx6+YU7x//ymQgt9ArDe2MzhJejoqXuYIuLyqaoKVMyQD9jJ4XCf9o0JUAz/
L9SjvCaNTQ1MOrOEek13GE3WrsLwWi+aXBGixHPd/ybih0lSqnBR3DyAb5EmR2ZBQ5UI8lTzOE4u
lEqd/dAsDlDgqLO5H0hBdK1JZlJGOQ/9W3po6j8pqkY+CvBp6RVx3WVW9mV5O4KRnNinRguQxztN
93JnVjhEPU9kKg4GVUfVAaqUB3a0F+VHuaQxLg6jWie11Q4RB414Yb5TeYib4uBVes4Vs34amyRR
b7ZPjyZMN1pQVvQqD+1hI+H+RC+mmyee+tGtbgav2sW8aaxfRoGDnLwQ+3CnF+gMfRRYIF/dN/ZR
vlJ53etasw0rFKZm+uLJUyO5WxO6kZDIyBCutFkVBcsWFEIRG03s8RQWfAWUzhwIXBhIJUEwAYTR
kGpK7HbZek0Wpw1+uKl3N67u4RPVcAzo9buGcy5M9T+8qhmaEYbH9lbkWqRFBWCVi5frHVzVqRYQ
6iJQwwAjYqil2AwfbYJft5V+2CCYIvwTHHRZabe+UT78w+YIKW0biuDOywfPBvTnWpDanFJX1zvC
5j9DfAK9SMIfJn1dLAfqQNBw66U1/JixKF0n/Jw4kqrVFuxNEoGVhSPM69xSCwN69J0bcolUdFta
298VEqFBdCAyhbVKCXieh3XWWqYRDaQ+TzoqwrlRMjPXKW+aeoWPyeUC9Otgs+hPGKOMlkdKIKaP
muLYxOsUIgwQYF8vzxlW6eFMoJHB622nH1cjzwU9smpCXO4uD6qKfH7tj3INDAaXTHgMFCiUKbJ4
i8hWHBmBhaNd8YA5oJorKqTiHUQdcI7i/ncK7g0gVUiyKN3aDX/c2QP7zo8EP+ZesbJXw3WxORRd
qxSSWXmUkB0y0hK4RcyU9SLoJeA8aMup9HMUO24diP8KiYWzsJ1a3Blu2uJ0HoYWNVrNsbslNM5K
/lHJwkRrCEQ5qveLM9pmCP/FXWTQW5WflyCYZ+4WPTuDHI+NZFVq5qZ6OgMW2ZgvfK6aEt0hQQis
Lnl8vaMSds9CYD0cbq0+jnGBEGT1cmxNsH2sOzudYISE/cLNHkJE0zGUdgOMucipI5TdnIGoR6MS
WGiVpPAjWza30FG/xKnkTOFshWolE/KcP7gDY6XRkb6v0lC1FiW8W6hGACt+sirQRyn+CXcNGPVP
4BnGwzU9YPvzm/LkR4p8ZvyB1qD7LRKYPJ69SsdOepgaeWhY6EO7dvhm1n1QJUdzEk1C8wF+E4Sl
r7cxijzcYEjTvHTJP6pzmwSCq3+TmU3UwcplQoGGmE30F36n+hFmDXFd5YKE5H4O1ERwghk/u2Yk
go7vApHeVJEDoGf+TRf5k7UpJ226cv4QzbzWKFaZSq+CuGCxyA1M0vuCUnEbxdBVYzFKK3FLy7Pc
EMtEPV4vPzqLD+QJEwGd/dpq6XIZGAn8AiCJjrJ47zxfJsL6fBOyoshdkqfykiDYiWuFE/7YRVQj
cIcOWoRk8w5mSq5IuAZRbd9eaWTwAii4+norCcbQtD8U0KRNnpOU4up4adLK+Tahi8pXB8JqdTy7
O2inmuD5gM4G9jjM9kDKmCjYWdacFTIBrrsZlzGswKssw63sckZTZhaQmgV1jsDK4VbSsFNzlFh6
p2Qg1eB2+Ry0Wr7DoLWycYDXwThYQekaDgIVD6BA9rIQklK0hCJ6IG8OF4eHfN7Xcl7gFHlh6Q+0
OV6SJAA6aMYOrsxkiNIlRPBpC+WenNjI9oQaKaw+QEmDxnXHV6O8TiAMjVKXizes+pDhxrB2eCH/
mMm7st9oxHUvObHw1rLeIdYnBl/EFvleag1EyWJxRzN2BPiQK51cPo8b9qAVD/3i90uzWnXIlRwC
QW0hWiNFmY79TzeULL729bo4Mga852P+bpLsqkRUmrurjshK9T28Frxs6lI0leymhGjJrrfMoYsc
yJB3e9+xxIERKaMeOI4uBC4ZK0oBECZssgXhhyjhjB++swLog4yaRvrdmSU22vRRPTmw4NEZp7n+
R7UDIeznmoK6OZeQ31w9d5QHYDMr9JFKJLGLdBcBOvoHAZkgkM4hGaIGTeFnMkN/6xVu2wLM1FOf
UMzMv4Yxf5WN00ht8mRg0oXeViMjI7LHEJGhtP9Y5QI/Ungb3pfZmygvlj5adm4zSZ7j+ubQeoWT
1Nzt2LPO829V5auOszubc03lWT8IZodPmy1ftZFPQqgVkVJ/Us+BGJRJOVXuqQG9Nqci/0W8cYeZ
QrI7hxEUDqu3GDIGukblOHiRtc2YLAlJWrzaIAfqzHVy352HeL0JcA1NPAJo0qa2Z0zzZyaQ6GEx
fLgKcUSJlGRtnwt1wlgPZriTR9pMzvDjWGsvP/Ss8tBxYm6AtZkCBTP6wtJ/ZRMQd2SHyNsEeteH
yXbhb8CL88biRzoBHkopV+ZSU1Bd98Cva62kPDqlGq8caAWxjOYy45fbOzTs4HyDWsq3UXYv3UuT
OYwLzPS1RF1booIyEg6i4PKH0GokPQZQdtYWSJfMhFXLr23sbwawKMizdJQ4UnfYJaO35GOMirZX
g26K30ttv8vfaLoxhLFf+UqshzcLGZn9e0JMVVbSjJJLr1mxISGIGsJum5iFyLZnthAGec63rOaM
/0FnQ/i518YyZMpmXsUZf8YrTMowicyZ4wKEgg+iVxElGNn8wk8wV8MtuPEH319Ov8Xm8GiRfak0
k5TML9ENKXLn3830F7t1RZerHayIsh/HrfT9/e8i8btLrT/quab6n3K6vthiicn8YGmb8wyWVDhx
81Rbsp0JVFu5EeC2btxHXb4GCmZZJfDUSjNZpWRDPmDqPbHszUpU4R8Cc/J//C+h3UybWKsPEbDF
go+XT+Jn3wmPPBQUGfPT7nufhkaxdu8EYCHDX7Y3lZD3SlN/VwQeFXUdoatlt4HbaFAl9fGEZn6P
7AaB4ZwLxiWu06KypVyELniuSmJsdDG+50PFB92A+zsyIXZ3yVIu0iXgdnGpG3jtoQhte3YGLUSh
ebXUJFkA2k6Ksl+2huxwbC5UhxtiNiSP6I5Bkj5k+gt5Vb4ZAKXPqRd0Yw6Uyo4Sc8iZKEpy7pHx
ADHmZb8fhW1I8lfAX5k46FeCUdh3H5vUeZMMMGu6Y69lGR4IN3re911y4pGXJ9T6QJBVB5ODreeW
TVUPkByABpNq2h3HI11eE49VuzW6PZOK9BHzFeAvuulcPfxdv+8TJef3rJt2G4rLJ60+DNlRRpwF
cMLFNvjvAbuEk5b5B1QYyjR8bJG8BdKcLLopiHZFY+Ok3bfP9K7K5h58qVKRkP3Z1ELtEPtgdFbT
AicyEyoxys0m+LiQFsg8aH34GQXYKoNvMKK6Y9A8QtI4vu0C4/omhLVKiH2vLKCQsm3NeK2X6IrD
eUfnnQ7YhBbeAD34tJpeKOJI2VSiTEZ2T37hzkSk5G2aCBCQM+gL3kRJt2t/nd06USpFnTp6gk+0
KeL/4yCw4wxpHHofeFb1/TMMh76XkqkdthcHxbiIlXZS/e6YmJ7cXqhlH8/t5kchePkqXKKRisv4
usqt1G+S3U/CZhKvXRS0fovOMMj3xGJH+N0/DX0XrOrvlhFkmBV3Ydqjqn2oEHZzBIvTMysRzjRA
kcpeELoSzMq1h6qZPPV6rJczt8MMtdyLuJDq30zz4eBUHTForQOPO4kMx5K+hUpDZhGyQKH81tOr
37hjml577Ec7GNseCBLeYT8HhUIjWA3+qnBFhIg/Ay5VLvHKqrFHm3a6YDq5OiXsEpfx2yogMolJ
u0BZ8j54r4RXqiisKTbc5fkgzn2b2ainbyHPU83sGBkFjxYY6E2UbtDASqhaumRLbTNX0qYx6S6b
q5kM3fSP81Jnsb6OoRKtFzLyVwFt7MtSVs+VJkv8F6rpMCQRv2nkzSsGaSXHg1Z5CmAWD7AS5erp
QNYpwSpWL2hPwmxEHR1FZumyitrADAGgAFFaq9B7pMCnoApA6m7Fm7xvceZccGKBOWVpSvsRwav9
aSS9VP3+jkETqBvnAItRr/K6SU5KY0O9P2OL9wKw1/sEmwJ14SzcpJaKwoy3tzEo1wGx8ie7lB1a
qu2Di22Ri45N56SB3DqpNNgCOORxXeLZusMX8xlDszlDWD7ByiggrU9HPhcdBIc4GrQHS8qxDmoI
yYgPEGXqYNjEO1dFWEBqgshSOcXHYXU85BQp1EiHadGXrjMRAW6DhS76V3uOfhZQe+oiw6m/bcUy
GugyDN+dwopSADrJ/FH7Xz44fCx5QxQJ0nks2oN5I7TrCDI4xi2TqQG1BEh4qLtEtwzSGeKUrHI2
uN96t1eVcueZYNM6PGveEMz9fztotHRZz8cUOTQfzJ6LKC6ovEbaFC6C3BUmvAG6rmWoBlcQPXGK
Q9ysbupJsbpOCqiC27NH7ehqwJgBG6Z7mvJqWTOE3oGbq78HiLDwGAjap0cHmc6CvBeHCLN1/J+4
sX/CHjqsIXQzFesOkPSDfEb+c0bKut+5PQfWGuRdhfG2ECEauYSXymfskAWJtvTsXNYyebt0t3/C
lAIMA2cOcz38wwEaCdK5caJ0wFpolDvHyJpaveo+gHdbgVx/k1BvaDxBaR3Mne1+4PU2fc9rjxia
pSi2GXUgGFf27bCSVX2RjC1b+ObFvTb1reVVhaBrfcETAryfbg/l0c0K7x0n1e+uDRS7303LuV3N
yE3inkrnG6DcaWTOG15fCrotd8D4NgZQ9NidLqcD1hT0rD/uSFRGjlkzauqBHv7bIorXBhhA7rQF
drXVNRVqjJWGOFume+ol3Sn4ip2v8+Fx4AA30SInCvTJIOXMw4Fjd7+QT1H2esoCxYkO6sW/ABGr
YTDWhDo/o6TKly/rOqaDxr4w4/NYKS0r601lUWiIDk/jEW82HzxdY3hYWr3lk5Tqtbt0BjTA5949
Z1wV6gPi0lMzrk6rTPWS2CvZpyuJQJ5l3lo7zauEK2tekLPig+7OAasUyG76fbRBX2NQ9HxH9pOd
CHyf9cwg/ZpUnRQ9N3yLLgwM3qV3CjNKYz/RAwP2qWlNHzcfh5zh7qpIC1qsHkf4RYePLomYziCu
8+bB/f5nexYgO9/ImSyIQzgpDXllc0O+2rJvpieuEyNJCs7nbhC5IaOeYAdUDtTTdkNYWCpEs6E9
1fyS0wyJ1Ubvr7niTOVbNTfpK+X+IWun7RFfiZD9MvIoWBK3b+/unfNKLbLcrCCpxcuQra3lLqDe
teC4/NoRG1088WVPCBGfOJ92VVrNsSK4W6wyIZ9R7G0zCf3MQgaZFyk48NF1wmujGxLJmXmnnv+h
9rjRHLYwjcXFCYSRlPn/6pH+ZXcEfWqLQYAPQ5WAZrGBEg4DnuxAbRygJPRqPerGdNSjr8wlpZ7N
YjDt2/l4XS04E1vNi30biFwnyETj2oO/JjqeouKZpVUQCIEYaM6MRdmE5S6WtsCYIcG3CUQcmRnW
WaW7xusvwrZdUfgPCpQprd8LIVdnDxboOe5csMloFFkDuFlzvorUexxEnnMmUwlXAybsvHjXOpFi
4hl+y4d3mx7qO3Al+osMM8/9KojLeThzjnvEJ6HywMbDVDDtcJj9GAOWrfKjZOi9tHO4bZ1ofEmn
e03iPEtYzzGI/uBm994KXgmtxmHEfdj4KAbVSq23hrhJQuiOTHsW0COrdZfgckyjzPG146q5+YVn
oGrK3mlzxQmOHnTyZzdI4C7gMkZUYrOr5KOlC+oePCymNjOtEfLfhs9R9G7GOsS0AV4daxTxDSuN
/qDIPgvoXDhesywK0S4ZkPH2tnj0DhOQNPKdoqhrW5o4iHHPM6GtwyT5tDLrhq9OoHkSK8lNvvcR
/sJSmeGwsCNJU6BB+9n+V2TM2Qmz6jYmSSCbbTp5lvt8vluNcVigHt27P9N7MO6BGRcFuhRdTP7O
UAYKSXUJleOPlBYn08Hg40QAsG4uG3BTXziPlPaKCfyjT8qndxhhET2dVeXi9h/38wvCSbMOkqjc
wP6ATNiJ5WWxDUxYHaVWgny42hCWS627rSFSdq2JpAH8GLoovKHGQ/zkcv8VDyTB07bly9eTEYWZ
PQOuOmwu6MSZte/ewCRiADdFOCYPqVe8yHpB7YKxu/FHU07uEzkgZKqkF5nVHCo5YEkOUM8KIQ96
rRrirQy29TLvO7eIuMhuKqBmcqXRn1oFIzzQf1izeBkPGYhpR5HW6PAu80w20FjS2End91Ns2Wt4
1fuEXmbIDkM2FdjLE0ifjBvfYY+KuXvSxPeptyvXDXIzsWCF6LLQDXu3JAtarsQ8QHUmui77uztH
biKm9H99Ph6xJTBQecN6ypy+XDuqZ6HbZSs+L1SH7IovliT+0kczUR9nJPDnBsY1h4giFkACorpW
noNuD8U3AymEPNAeRMQDLa5GoX9xFQzTDH3JwMActWpdBSl1um0KrPYXBQrdSckk1iZUzyWe3djW
Z5gyHIIjVftAbJPvrVpbV1kbXwvUObQPCTJObvbs67TgjbQECogsVEzUY1FUoqPeFs2O9bswF3UM
AepXcFBsEBUFJJhyeWUtpPTruvGHw04HKkPSsKxo38QV28nznhx+tOa7PK6rixjT6sl6vn1i1p7x
7R9x+XgD2I02dcxWAO4z/KmhPytN1zzxDU9gAjAkv1Aqy1Mo6Ndm4mknsC7/c0/xXU4Kg316JKhx
CYZAkcVAZ2z1p4p/bxd2oAQvit55fkNI6+vdySqej8NZVwt1UB149bC7Vdh6ojPzYEkcfRz1eqUM
vasKPJ6i2ndNhboTCzhMZBEluBganZtu0nCSVVGqC/BGbjaASHQ4K19Y1uHdocNUtS9ODCVn77SH
/5tGSm2BLAjOFoZOPHyNQR0hi0oKpyM2g8Mb5XDHtwPgp9YLK8TUwosL9+54PRNuJJITx+iGX/Li
bP0Lj5iZYVzza3MJnGV0DlaLv9tpar8PjydFJcfgs+1tBxdu1vbhOLbWSyVQnB5g1x6mJQfVAI3x
Wc1goPry1AmrugHwzp17A3657byNSJQIxV+3DO1Fwbz+wnDE7MT9+/qMWhrKFdssFZrBI8YX4ZYn
CQ3IFPHojJq9x49luanDZObW0fTuJaBZUHW101FwUADAOyV4Fsl2VMxaiK20ToR7CkO3Enb2G5SC
6O1VewYT11VnRPnSBfqWWioA0LgM/60ZX9+rAvV0v6ryhHgFDqQnUdekEodKJ+HZt3qQUY0OpU+a
KP9RWcc8RAm1Sjmk2m7CCtLiMWn9uR0Jc5qHOIEVoByUKq0q3MahznSzkluD9NGrUi44/aynie2e
s8JrPWDxxN++IZNpJAHftdw+OZWBYarkgJEb9RiuIGyEEz4uBb+cbqCL6HsxWQ4FnLk7G2NPBw3r
8atiHlaQ9xoqV3QANnWDYJLhetekyuKRXIdiRqnw0QGpHquDxrT2dtQJNZb7XARPwbYHHeBpLDUH
4Jmp230n9G0FEYAWP2ke4XsyNqLO9KD0ktxCL3u+pOUDFUHWV9Eii2Grq9i+m2gIoo/9ecROD2yV
L2rH1P+I2v1VQPhvtcLuqDFgNtD4t6jXWIIG4l0qmbsUdbv8QEa6nl0WxUcHTLdNBiIk7ylISWm0
HgYqf/R7hIBOMLxjV7L+zWJtSNmPJmyqi3MBH6EutjOViEEuk6Z+zXi7Qmfs8DmzIKzpcXPVeG0e
ubGEiw9bLQ+JTx5D7dkLnrbFvaH7SWrsiTURMWjK28turEkmLbvGE/8kmO7/KgjoZ8lcXzgCLDg7
06vIGjH+jSoD9VQiiAix02t6zSrKarVNatcYbfpkKcIckvU32Kt2FEvQrTesxRFtN3iCX/H6KgOo
2UJS2Km+AZ6v7hVQ9Ovb8bCts+D7gJOwiHbLQbIl3cIa4kenPCBoUuR1AlRaKQPJqDJ6bnDZa/mV
RGj4Yc7X/+BvN2Kk8T8D0BeZSto9x4kAWktufxNv4/JDwe4g9rhkmeLYLl7Lv3HcOgrQRPHuF0FY
AMKZ01hA7buNB72ZuJtOEFbr6dFVpTcRLwwpM/aSOHasfdWXA8ZtP1TsMzlTV7UMiJg6gu+6NSpE
YcXqH6v7dkCaUZ4+XTdTLRRkhNhuO14SZ8ZxL8Q3ReQqRXZgKEQqMBlOr+1e+HyvcysFFAiOMVGK
qNmBJ/rU86JrAhSL0ifsGLsATg7CS3V7pm4D9D7O1wWu7XnD6c8E2UmRaJxDwzFuU4DGT/6Jpp6Q
45a401k4HQqOAQFhRxGZ0pwQWTKRCveY50++wwdzkBORUWCqbJW0vVZ4lcjF6TO/kE+Z4pQat7TP
K0OOyZAEWG+10yFlzNkEH9JbDGKvk07h/TpwTVbrSsXfEP1vOHepfNF4v0jRq9hGGY8SBzB0f4t+
C5ZeKLgOo+CfF/X4sKJQJ8iBOmP58bQPe5bYA1co4CzwysVitiIYnu4io9HTQtW+BF4AxT9HPguk
0R2NRRGIb8GZMJE405naS9icHgg2F3f0pOaD5MAeWwfI4IFVAmZ9q2hE2p+o1thbYiBU5q7SqSBJ
fiCX+oZSRswY074ayUET66a0dpmYNwNc2DnHxidQk2EAOt0zHGUt+voHCvRWiLHgcoLy9mpO9eSH
urso2Wqm1aT2G+3ATOJmUfe8LWjbIArqlbTlnfhaaRt/C4VsNFqSd7sNfJS5uxl/qbFPvrlB9p92
s2Fz7usUm55z75JPcLpyEcHuz9o9KacXjaWPFmMq94QIdV2tvTsRe21BlVtI/PguTRSUS8BsXw07
Fo9f9nCGQf9SVdm4zDM2VLzW6Z4trXPfp2/pr9LanSIcgGjlPmzMuQlu7kbSiYOUb65jcHkEGo7K
6XGsQYgykw+N0sa5LxqNjFqBgCq8zDOL5zXwFHAkDmWzXmhmqQ7ZMp/1EPGP89++vbFvAHUWkYGi
T/loCaOnPDQxU42OiJUE0UfMPCRLK1c1/QMPRBBXdtczGadtOw7KKZL9z16HDvanAx/vZGesP6HW
4uzZB9EFc8oGAb0Lo/qlIK1NOJR7APzNkeRDsKDXw5b+IatGuVzHIePCsPFIT4VpdLEQmeArqgJb
ByywBSelSgscwn/ANtx7OUeFgrjAfs4sKkO21+P97ts81uSkek1WzJTCIrJDSlPjxVzBaYxGXIFC
o2ddxaOCJjuL6hIAtif25+QUCyt8pDg30eXPcb0ZqXmMRv7X1l28DhRSc3jNdnV/OjHv5u66d6Yq
TiBU96NZrnGRE0W1oWxWqvp4LVY5WojzDZ7GUGpai7bMWmpepg8XDoWN2jhlwsHji4oH3W3MX8X0
HILrAMbdBB4b6cVY5Z2oJ2seApx6k/7eAW8L2iUMCe3eNlI6WhLw0/6C6CIrfLrFyPSYIRXlHrHl
d/oWaGGq7qQhZxCnkU/uSIxuvKVn8cEmcrbwqLNEDYaJsr96FsdKwRjlh/XowJcyk9qz4XZsOY3I
Tuqb1f1LqiYfEzudcU8XOtCd/e5wcfzgoXjQJIH1lwkdjEF248Vl8fc8Qpdnsrfa/Up4v/bm9BmN
9Er5DAsOqvxpwbS1HWDFoiZQyfzYuItRs79fFRT3XyG26Mqjwjzdjv0oJJP9XoqtH2qa26PspLd3
RmTUTyR8MysbjInDVFEgNq36fLe68T/DHekpV7iDJ5njREK9YiIvRwNh4RbB4qTd47oSx2l+dwyy
+y8T/3inaYZCbofmwXwT9ZZLoWN9IhcyTTudtU8dER91C4n/jC3a6mdDlGN563MhjcfB0kjSNw1+
3QZK6whzFF3e0mU4TesQfHUSJ6sM/QyrZnAcFzzyfuhTe2nQyn3nD0pMIy8GzyreZgTDexrqrK6k
C2Swkz79clSFC2pVMbGFcyBM2eqVbPd8ocMaSXzjgM/Yi7XSP23t0H+BtFpMoWuqvL23ztXvt+SU
4Jyg2OPMMgdGb9gyfzjGuoUIde99pw9wEV+DIRnv6FwkmZhOaWrQ5uOAyx0s0tiCTU9/FEYxAX32
CUYDqwJlSoyJBoGii0IXz/Nwd2rhSEIETghsFWyfeQ3r+TTaEuFFo5eJ1M34Ny3Xrb2nrloRVL7X
8ta9yilLppCiLyf4oXwFVm8sdhrzMWyQmfE5/rkK5gc6L3CC6/p1Vq+0rCwNuw8p3QDPRead62K/
6hn1AUM5h3Ix+8BwAdEgAEaNexZfWYYnXSXO/tPrHycSrXAACETlmvryObtUF3Q2/G99SXZfHbfT
Q6l3oCe+rG9GSFGJK6TlKx0fTPVk8gha/ktZirpYuOA78ygh+yMrpS9NkOxrDNznywbJrxB4T1j5
bhdo91yPDumThYrHfKnOmZSC41SHVfZsUdOpFO6VZc76Nc+O7nhWw/CIe1BQWkDFgYokZWHIvHor
G3KvpXqVF5P1pbGObrqszvgIS1DBrgL3UtGKt2ovwa9GbuQVHOFaKECVhnfO1vxu3Q0nTVqfSJka
GoQIRe2RhIDGfA0IhWH5RxgG34PFxTReF/mGwpPr4huNsAceCQtXpBNi4V657mQdiC+ANKRoInee
fc6XJRxT8VCmf4PlpGIcMEyVC24X0srqdpjaQ5eFu+Nx9SySb0jIyBNHB6nEy3Zc1O7yPMynCmc1
gkj2VZy+5RmHEekOmhKua2AC4OMXD1EW39/w4kgSh/e8toRu+KTMCVuN3E+XCPWuADIh3q5/wiEh
X2rASuKrQjor0V1aht7m7Z0RBqyKw+MfHrqBnD7bh+7QhT/F8/h6ZMUZNZWfQxB2qwZxs6llrftx
uNTj+RFRddlv4Azf2gYQbNARgmrW9TnCN0sfS00EKcgp8osqiaIjHhSUNpVVl913ftT+QJXQS3F4
UW27UvfWKFtwCcoigOPV+b7or17XHW/YJ8YR+LL0PP7s5eoQtEe2i38bEs0X+Oq7N2V+l8+lXu8O
8tGmNABALh83k4NfFRXsd3Po0etJvwBO4MweSKuhCdlERc9/RrI41RsT+OlyFoD2r4Jlm4Y7inxe
I1DaNn5mINukHzEwTMv2hhCaIZ+fpzmmFQzuewnw7POa8OptgHKeqCMGI6qMVvNBLR7YppsSAz/v
k1YAbWZG1uumecxYjPXiUZPCQP4Wgzd0d/Ag6C2w3VT23AES9nNkzIAWIYHQArCsE46Odk+9EPJc
sn6OAYmr8l3RVJimTP7almkdpTzcssNWAea8txeqtdWPDbp/P9GPKiMxrONnLkWekWan2KKNzHke
iAuXrw8ya6i7le0KQGcRv7Q2nvScFDcf3UVswMctKQ4kRF99dQhO6ovWSQ7Fi368mLH3+gjI6R5a
JEv7u24X3ROVYNqkGpYwcti/HPMsS615ioO2llU1HvHQOjx6SaTDFvr82QZv0p/QHcu1bLM98ZUe
Pwy57uyaqSeJEiuaZ9o0Qr+s1Ssa+bVGiPTAZ9Dls6X66MHtVj2fYrgpxCi/8o2jpoiZaDUkguFc
ZF5A/XC1q1g0j/br2PsXmlPDHS36lF1lQWxO1b3O2BAOgf/dsm9rrU1/9CK8CIEsLgzVr1PJFDIK
2RdL9wyjNhIB5T9PubwutWLInPbMYfUR6j2u+hOw2p7ayH7OVe13Q2LGt8Mx+EarRQq2CBwxoqzm
TRfvWAVJD2jJU6ExWTEsY4DoPv8DwCwwHDiH5rnDWEUSzAQl6zdpUhEj9za9ppPo+nz1IfVQqzRb
JdGbn3ftVHWWQ77+gfVZnE/IjVXGqN8VZH2q1c51+KuFQyAfOOeoZrSp3+6LHrdLtYQbjO8fCtFx
ndQfi2KqlqsDL0g+HKczMlmTGh/Wk2znp0aQ95WzaibinPmrNxHz+s5pVx1KDHnezbxQj6KhzWrV
yXiMhnGCxAkpQ+09SvmOx217yOneeR2QUC0kntZVs48NvGPkEz7tPmuoZ3/jvvRW/4jlYec+DTEA
I4BOluEomosVzygPiOPkjLzC5v97DQJgc6mITjAXPGTECoe0zjrnokFJW8MPUHXFvhbra0+BmjV9
O0qZbSPMMYlCl5YMLU2Inb21ll1nHCR/nQBHOP6p0NY2UDq2889X7Izt9jIhrLY/OwY5KMj+9Wsn
ib3JjSYB4eXVAhq+MZRnYJfgG8e+VPZ6aYxqBXNzlXhFCB+VEDmSOO/N1uga/Qjxqg8QQrsba9mE
VpzHMF9a1M6eZvCs8l5ZBzX75yugl3cQiCi+ASaEAV2z/8NbfueYRqhnzcg+tk1dJbCM02RkNBog
pmSS6UFTrveJwto5xFN2RtqBnOjZlKQ5eRw2T8l/pou5ut5xbYFQMpiI1qRJDnsWEHHkSG1lS2Mq
2/e0soZweFAXpX5/SvsOoVutcmMFIyGpvIDfy93LRsPByA/Tf9kVYKG0jdZFhLp7U4jVtvdha7sZ
XPy7YG5cBLVOKW8V9sixlGeJ/+Ksd4TuCFuXUbSCUqk39BgRODohzTWx0ajQPokaxrDl4ZSx9vdB
cVEAPt4vGkDw53+jQDw8Tu6sL2yUrL9xAMLr7teKua4s6hyzwJyjX/tNiTC/xT2R8qMU3X40r3ad
h5XVqrBCkbZMddU4OxpswFsYWvKtb1zz1cT8wKYCDX03XA4TatGwfFXbIfGDwcKLyyfVHbvUZYJ4
nzkSLCb2DUAuZM97kqy82zFPMKxptHc8OkVqsgUJHu17rjd9rkoeNUcEFC72kCzcygnKYQjLwGw6
chlB4JmNhP8+XSTW35Ehk4ZGG0RdyG7hGhLOoOsAEAN0GGfXzWjIPOAD7o2/3K+D8rz0p9VkybyA
ZgAjzPxwInc3D1zzZFz3MvHlaI5IAcUooPwe4scki8S3tjEOEvQ1e15cOOlZvWe7v86e986AeLWi
ge1oO6J6WRQfN8lijbBAaeQ/kTCIdWPrbIDDP0nbXoMA57cZHqK4AZ9XY6xOOvfeP6eJrXnvjABZ
SUYnnN14Rfqlr3D1jU1/p+AE3AXPpIyUfsVPPJF+o7YoMtWAKLAigaDOK+WBXBOSMR8HKOlvNnWh
PyLncULuFWgWYlO7P6ekzr+ifucTK4xzPndRcNe6oqo1X9rb0RqQQ3v+qS/PC362xKMoXlP94IhP
tIZm3MP2Gt0A/RnwWJ8r/X/digf53RJqU3fMzB6/GsI1pN3YvQLdE0UPdXR9LQAszbqaOA35r6Zf
rpxZDLeRRvdySDBfwxumfD67GizW7LpgBW7u1abUj4GkDIe3Ktzp5U3ba6XTA8DYC7v0z632tUnf
8Khzl6JSWQqeLGpPsImsUOOrHiCAvagEsQS+rzSnBl3fBTHPJpOahxBWf7V7DwJeR/rACkPBjZ1b
2jJwHd3T+iMx770Oo3AA8ZBG1azvD5zx8+oZykqzGRL28nul7MNyyOp/VRzrhdDn1KWAQV336f4H
iozfNmKmWf8oPXv6Yic1U1j8APN4uMJrB9FINFpjkqwTRk4aEdkByEbapG3kQd19Z+igglh5Zz7M
Qz6MaQ1Kb5eNIkRCALjWtgfCVtNrtKmI7WJU/1g1157aoslEU104jQWVs480Rfg6fSy5XbqMJKLg
lAOlJVUXV1ogdDzp/QbHBwBYL/gZhbDVDstX5c5p5ZqwrrZsYk7klKOkO/wMAK3imUFrZMVmFPUy
DM8ryYCrBn1RYggJ3Rmtr4n/SAazwZaBWJQaJV1wMCAI4SxiFzD6aJxb6FngiwA6u+AJ0ROzqTAz
cE9MMfE9g8Fbv4XVAbEY1BboOiu2Nzsabjdj+sIMUrP7KWhSNjiT9cqde/dQeLSZ6LWpuw9zQy7q
hEqAvlXazz4XiVw5sySl6YPRYxKxTLD+7xbjvJcByheeCxq8ZWxOzyHOLfObg6ZMB3jvKuJ6m7Rb
XgmleKKp9lLyKnzZVizeSzwY4Rfv237etkyIPErGelEajJUkNJwv7jXwrMEPhrOUPfN3wQfJNQNT
T4VJtOSPkwlAcWQVgJ33tq/N7lcDxnuHuRk2BUtTDj6MNuwDUVK8TftIwz+ysGHXFzJZajud2KPW
obf/75X1BSsCpvuYFFi6ynuuxypuA1QSw6KQMmlu+A24ClSxyNNDsQiLJFNVgmO4csZfnaJoMh2I
63Sc+zs0y93hPqV3LV6fc2amkiXmsdvziYVICGEQ3EF/J3L41QlUeYw9eHlHcg8IXpPlBvTD3aOv
5TIIqlx6Zlf6HOWmiZHfcoRzM1T3/I+9VFuBTO2vCAPSTK7BGM0X81dxYikx+i8FnZA0DBUx2FoJ
nLqQZHuNOQkiP7mu6EOoI6efhk0zgAZgNvaQf5eHIafgZVgvaJgaO/VH2K0bOImtXqaAac9Ynu0A
26WuCtuQIqdaxIgr8Wq2fWSNgAWQHatureHOHjX5s/0CPyQz2XPP8vK4EHwcOzKIIzGiq3vgsnAX
S3wd1I+RXGEcLlJ3L+s3NHmxXzOTSQ1gFvDiUozzWYaxYhVlFV9e/7HUPNscyWfHbQIho+saS+mY
Zh2PU7ASjI+wgNXHf2FouO+8vIX99pBng7uI23jW6Sqv/7ryDiS3HOEME0W9zB/wYGZ63XLp8iqy
h7OEYk9GF/NUMN0aiwRKS7S62Q22smn2UYeUwzyiRXRBZH0gW+kTjblD8KaObJ6BtoUfRxCeO5sX
mKENiz3IUJSQC7QTg0oGtLXytF4R/LwXf+F1ys8zU9gNqYWzwAdW+Jv6Kqq36UZJDAB/k0D1G6M6
u97zOEm2YVCaemEDy9zE7dd5BdHbSQ+N/PM9QwD8oQFG5s2gFS3uYwD0w3f6ojS6nst5iAQUPbF2
V5CvkPCa3ngxQZ3/hYxBmO1tCVIKzFlEA5F0LsqYE7QjKkCML54i+4i1krmgsjpVxG8kw8TOGvvA
6BlOAOnhhZUFQHpZvLg2WoStDj60fMo5537Fh4iJg9uqQ32bETDjdoewXlL8HXYdG0oMyp1SPAny
jffCJn7ad1V7gK3hd4ByHsbfXkawjUVVzqf13slxeUaU3b7mSZcfsooh/JreoS1BMM9fTHoJ3SlB
ZpkKiytJWkIa87vZbVX9rQeb5EZ+NLww42Q8VUUN03lF/YgisQokGe9UTcTSOBvw28K9DeHOKY17
s0g4aXIfupDX78frTmR3WtRUirn1U0wJ1w/BjAnmtOGGQqWL6hHaBO1WcRR0jZ1uSKnD0PJRbXXX
2aKch9/9HYILs4TmwB1Jxm/Q/7cZrsGGL5eB0pCWIRjwyDIWBk5an96fVVtB49qhoBwaHulLKCw1
N+6hxt5JfBuVmDHdOlDAYrOJRsJT9Cvpuu+BcPbP1IEsk2c5FRVWKw6tgbhVV8VEeQd/GbzPlAmu
b4LNg5c+yCjOF/32PYG1aXiURH6aUvY9m0RQtCnzsc0TkBBsUu/DDiGGH5A1o9N+OcPN4CSv3RXB
7Ir/CItZSvGoHBr3TdnOwk1PgVWiVKgL7S34QdBPYAqtk5B/ZwbYFqxXTRrG22FBLVei+Nl222i2
Qbq6PBAxVShcce+h/GZUVBPrdHR6YWnijcSN17yGLFoQfiNo63Jz41PpwhAf56soXDOpbSp/TD+o
M2HHukNoNAmghhDrVCwz5SsnKd1Um9V5WpW8aR9y/aFQ+QrGdDg7NXwvmUa9tG2+69Z/WB62M8kC
i0hl+xThYZpZkSEmnEI/gUOXVwy9o1SVIh8zIr+LHtFR11PyVGOApRenfmHqdLg3FyDp3CQr9eVV
LSeFhFajdDefxiCTJgzhzkyr5QcsVftbWsAjUT5d5iiytEsn+L6W+lzqCAhPPm2flxo1Y2BG7/rR
/ncTduDFf/vfWi251/rdk9E09MvCuOE2u5Dsk2hZMeQp7cVcbj6xj94qdhyn/h7gSGFjE2gN7sTb
+kl4bHJxSH+iBhxvkaIzecv2IbLPhAk92yzdCy+DfNs84ELeMqbGtFkZ1JzVTPvBOiZ7W2HOqQ+o
tXwjmxZCbRaj8Tr1+4BbdxXWVr9UCr53CT/AGLphSQyU+uGn0JPcox1J0wmVgb+WWxS9kwY2g03c
T6S3mkNECFYNHRzzzGh0AYkOLT5fqT+LyRQMRYmyguJx0d7nzozMS+VRulwzSNSaHhTIMCZBcVNf
S5Pc9QbznqFmgOU5Cl8MYHo590WNEjYKmb9D4wRFUle+rKBXHYt5fCvaB4CP5w6BP98rNUhL9UvR
VhddlRdKQDPq74+im+uqsHVUOMTPN8RrRanaiPYvnvRTv5TLGkLgQ+7KC/B7YqEWNY3EAYAa/zP4
JPnOFmYzfUGkSbvl3OaYsuGGyIcoZQtH4x3KQmcyikCg5j+lmrb2NnLI49Er8Z/u95bSfyqu3BS0
kSZfbdSXxWm6QK9bCEI4OAOQlxV7KnbHckl+0jcxOp3epb1EmnjORuflkyOVU4pxCdGDSHBwgYcs
Tu0TLvGxKYaMXD7nA4S9thaDuCpTWQE7mznB0otUvpo/hPfY3bUBjQ4JPT0ILNjA7NsOx8cGIOHy
mCuM7k38LkYG+WVm30cb8xjvIwaJPooXqHApCoRoZfd0nvhy6H1j9jPInQJLUCuDnF9/hiKW+Obs
5kPi+laInaJdSdssj9Qji+M9j5DWPxRVc4EQkVRWNlv5qA/EgM96O21BvkL5ppQgCJvcwbZ9V7vD
oU8KYOPcDXIvjSoMQddLsLs7dwvBspsx7C71brvzSYldaU4TBZy1gp9vFKFicE98sg+A7U8MzQLz
LrGusk4fpk//EQ7QH4W48wIrKnGVYqTDSY4XWFO14v4XbzrUtlu4Ln2qA5/aCErvHI1TlhUQuDoj
88nMGLRFggxsiUyhs39ATZfTbwezu9LQ8OdNXRWNJYSG83QKVbEJFglDbeWGYpfJXT46u6fOj9js
sCBKWNeDTopVIgnB8wuF+sqvrAGVXJED7G/GCRv6q8Q42n5V0KpOKjRyDlf4aJElKQPRfWp8nbwb
BfG0djLwYk4hkFXVS8trdCWM7ztj2ynqMoeWQVyP4lUc9FJoeYNPdVGe8COny4pOUBhYuIsW8a6k
bQ5qhePceJ9OmR7T5zwMn0SLusKLjQKpGxqFiX7uGm2PSlemlT+uzRfl8FZnBr2h0il/0JJtJLlR
28IHp39ZzpvT53ndfnqRyLrY+Esgrkrkw7EFqxqkhMbk/R8ssFprEpYlkTlniP9ihVhPdFdN3lQC
jMImNhn1JRckuYTH0az+lzG8Dkr+e4eBtlm+LvF/eOm4CPey+VUto6W+Y9KVlq8p3gt4NcpixYii
d1cBujjYs98x9OkQO7wkAk7lOuKQvh9uk579mjhyOxxvl+4vMuSTOsFmIeOQLBvolmFVmuADOwRm
DP3k2AtwR9W5k9V32P5D2af9frZ4ctAuR3ZOo/1aSgxE1orvy59lUe1CEJYkS5xruwxedi9hn8lB
yDcJ/HbsckmOZoFWwxeMqGivo2wM4n6GVFWSEuQQ5L43ahW+hMNO9bxGrlD34MAxX5LdA53g1q20
svoONpKy+giz8KT6W+fbj9kkyZyH9wE0vWilUti3LAyo0N7PQLa2F3Uk0M6jzyW4GXVlQRioSJVy
7uEr4iDN7KXDsyDjgE+4Hxt2UoU5pgUKLj4fMMkRRPpps6+AwHtZp9+rtQK5oABuY9mkgeKeXdmp
Sunt4MzNF2svP0wGt/tJyc4prHUTKXiRKltYPMlGCmoeOe7WqL/zazBTw3W2+Wt7LiMdxa+JhlzB
Tf6y7DIAJsORRUNg/ewH9MZ17k1/KG7gpPXONPwW4FBGP+1dZyN1vJTOBMWGr2c1Pf/rcNycaldk
fe84QmuWPHkPK88YQPXqZxASPzae7ZA7kCDbxZOvhzf8yZWd8pjXMbtudWq+IMgvhJ3vP5nWlRaz
HUjyV2KukQ5r9HTRAlfwRPEpNBh7diwVH389pyI2yLPOyG/icp17AT5ZTjWX4yhtuvG078UAdojx
lTxtI8s0gyhtmVtTXor6s02zq71lD9LOsW/tXyNrDw2FwLJu3pBVpo4xAWw33/f3rUismSICa8lj
eSIRzxD9BO6vasJwRKfSQg0aJh1olrPTcAWEKcJRu32uO8VMm2B+8KP8EN3LK3zhUO2UInyDUSMM
O2dbFPN+kxXo00opwW5JT2QujD4FNnvBJyJ+taBWiM7rYpckX5h2UXqJJRxPEaVe6rhxV5ehLbqg
uq3+eYyAwAZAuriQwoERD3KXFoAGtH/YntRGuGM4oj3lR6zbYLAoeFcCvz5K63Tf+xrHnUjCTk1t
A3wrKOn3TW7Qa8z0Qv/kfMFdAZ+wyPAsptVvjjAbr4r3hnGQDBogrfwCMMj07c4wZyILdmHnh90V
dBHXH+v9Gd6hzYySsIkU/KFRi4lRWKfWLEe/ZgyIe+DKkhCkTlFJbGSdOJtzKl9diKossOTlHVAL
1BP+DgizW+k+kSLia41W+qxoVfANYErgwMH6ehXWBMdBXWdDiSTPhWEXvVr8J9EQPaWT/wSW+t2A
jpTzZgv2yUd3qwC++rdFKxzMGTB9AUf2xKDtCFl1Cb4exXSgmJYGCI3cAq0ct6GO+PhROCtbwuRH
UdUXX8VEukdb1AhwaAZI3C1M6RxBXv35uAdyZIWLr5QxdP7oIqa/kWpTj4pp1Tu1aDSiJ7QUnWpF
7ViD5fF/9uDxU9fVG3iQE5Li3X8JPrWkFtSvHoAsimI4FIPfFNXRzKecawqaixxoXVeMEc3miVV8
JkfT9vF7/boQ9KGCm/tz9tPrRUdU5UH23vKbJQhfAepsCto/HtdgQwQwj9ms0HLE6FvJoXL6UtXd
yrz7mBlnC4BYFeaDjd18B7RtJJpH8r/3eqxHV4A8x0BAtAjYQUgsF4B/FlLCS2+sXjcv3mkwya1c
d2cOSjhcuKe+bL1HYjyOVNl3JRjt/fr71q0vS866hshyOAdhQzHXLzUVV+bIootpvX/2V0yL9FDc
zsFLOKMb4iz/dY0WYbz3pa+Jh6C1KLjKc6Z84aCy6cdLSX6Om0oiI7RsDnUNWfg4YtQ0BJ0+Igui
o53EeNrrIDzj+vB5X1gC0s+3XvB6moEh317rDaXRTvBP7xfZsza1NkndGdAb+6uQi8Gwkd4z5nM1
BGTjordJuqfv7VWGtyzMoDGRYhg59yuktfD6EjCKaVrfPf7gy5R6oFbaXy3lYs3RztQqUq6F9DG8
Sed1ytQEs8kapaVVPTzcy+2OjHb23slfTs36/rNDmyvTLqvjDiCNP/ap/oaaOjIL8X9D6TDfipQ1
VULN993mWMbmGr6a11URZoUijhLwYmEtYjZoC2Pk4LWBOu958C36L3ZTtvGvBXYsG+ErxiBK5aJQ
hCvw9ePSkAQCcTyi5XGvBAmZS0gdWLtvIxpxQXTC3K+YQMF8D0XeT6s1wlBpiQW6gn/0cr6zBMrr
3JNMM4zyC6KQKgWejj1Nc6Yqe4ZicDI0DI4E/H+/MIMY9cAAZuckAo+UmdQF1uv2CnqG4nN7pbQR
s87XQrB5lvfI5axhFf36JfA+rMnUIEgmbYPL3r+ldNbdjZQnS2cqHTUVEGnLyQvz1PuO0OwW4rZ6
t5ohPr5eII0MhqeOITXy6fZyOXEHk6vbxzmLStjVbOgZlnpioWqo1KX9phLhA//SdrDwKw4/tLec
qkLUwTlwHnF4GdO9HGYVQgpnSpgsLoq+Q6gSVV3H6rCASp1LXj7zr8gwy6xygcPfHeOnrnOAB2jB
BLCNV3yjC5Jn03dfTpG0gF77ftil5Ln0eBa5NImUAbPkl2AMJ5Rouj82d/Cb98+POSyaIRzVEghk
SnoZ9poee8hRqN8cMmxKu3JF57Ivpw7TR7P2o41CqYvdcguaKnkcUjaLGTeHjvhX3DG8zIkE2lyP
I8Juf20eM2PAJ4iBKTMilAtJamntnjgyulBf0Ft0rNyIbXwcUNa/i9BEAGg7LqFdZVToH3bWaUey
X222LnEmUFHfou+FYpLkOy5dmeTKA8kBMijcqKNgT08qfhk2Gmyc02T0onGG0TLu2DsZ67CXM8xY
FjbKDXAKbhqxoOuR07alOxCYEbJCv+li7+Yf2RKzVJOY9iP40/im8zXr9QZu/Rrtcyqy6PKaKBQf
4YHmE4JyNHa75pJEs8gv6U+8BTPWwUORHFPSMrzQ/lWF8/QAPoDM2vNNCtNJwQ86QLQ0WG11T2nw
mn543t7+yve1oPMCI3wFBt+F8YXGXoLr+b5FiEEK5VNINHB1iXk5Hj46wUGePwxUl3Lcegn83j6L
fgzFVdVsJ2v5Hd/0SfRnmWYIrOG00BE4TuHTp+UdlVOy9wc2YmJass3Vf7hJdbC6/F7YAvC02Bgb
imbk+SVEOfue85qfsoXl314WBDLihJJwsCnzu0OwIQhQOVmTbI0on4HZDp14kQY4+yjGyAyTg8hm
+J7nLf2FdLok5XKESjzmA2HR7nGLCEIjYzJFGLQZOomA66VkznA/QWK0l/vFxpdoaLOww9S1lvma
y7B+45nCzFedh4dJEuliaj2l+GNs+aoBA8hjfwk4n70jOC2oEKGm9O/hXXijOE+tQdJdm02taqbA
sQemGtKMOM0MhpmhWC6I5JCCvwv+FXdhZQ8DyjpVYpaCFspwMkMGxJUXYbZ+hcd7HUMeVvonekIn
KFZ7CxNm1sGo+6kqDlYpHGcwNCvrgO7nZU3apwanYNMMyMJ0hRSvpZpywzpZMJ94dK8k0fo42S/c
MchZy8KgO2zi8zH9fGyAu/+EVNG7ou374L5EibJ5HHJzXhkY43XktWgdIQRD8FL6N7lfjYUxKyo+
Nz6Nf0NXnBs/Ma9+fVLVxyirtTNfEnqW+yLa3oFpSok9qg1FxUF/BaelZw6n1SBY5Pxon9qp0QQJ
/qYWbhPevpe1iANwMbC4eOpEfslkC5Zb29M8tS+F0rj6kHbWb7PQBtiwKXyJgn8Acb7qE09V7TOX
HGFzCM2WFGaSiEsgZmQ3eq4FtFdIM6L95UCdJIvdhq5IYah93w8/X4H3WBc/pr/IvJTWj/PIEU+a
10oNdzsOgRRoagr8p3Vuh99kjm8ABWpzygZcPWoAkwPH/cCFpaQlLiJeo91VP++Q4cvXmS+2HZUe
Pc1K8/aCm+2d/08pjTdHUoYhVya6xcDBHhkqvLqYFru+BWmlIHbHCI4Hvz7lAG5qa8wPfHCIMS9M
FsmdsdRdA3tKyKorglW5zKndQaAeGJlgTAKt1T3ZLPZtQCNLm3RjuKMa5g//iHuo5Ix3s9rLKzTX
8XYKpR/OAxufCXbTvUHJZPK1v7s7FIvePb5PCLUtZgO8nNxqxzC6Zsk1WtRrs7zBKPtUOiRuU/9E
kJ9YjUc0sLgGU53JZfAKQ3mVyb6qu6xR1kh7TJXr9dkuoYcQReMFpA8Ese8qYy2mNnc+cYFDZAzJ
CTCVLYs09MK+tgSRa95O7rZZPNvmOyxpqeqgSSqIWYUpt2+WiXFHCFBfsy4vrnQil8A5/zEDRb+8
xXLqxKy2503Qs2i978gRfg6lHvZNtLZsE0KLLWzKMwrZs7UEgQnOWPLdRokzumjRKlbVeKc4Jl8K
5i1DsZq3YDkd/3ILvvnH61XbPbC01T++RQWE9F0PM9pC2qQPKaBbry+ALvogT3u2hCxPGImz/WZh
2b39WP0guFl6YhAzt93bRUMLgcDXIqpY0irZria9CWoH5bkfL8e5paZXUOxfxjyjqv2tTrsnoitG
2EDKA9LH0v1EupLKsaEEaFK6Qa/bD9TVgVeRs2t5pFJwxJs46pzpYDyT5eaVDZrjWvrDyqhZ8X6R
22V30XA4eXb3L2IwXcHsYnRH8rcy6tELIe04oI+ferQ/H4Z1yzYSm034ZZq4XqGb/ABXNcpsO5T9
biHwIG93V8urrbgkr0Zd4+StQrlt7oFP+80QduZ6dHnDYmtA4ROKw9lWbL/PHzaqHZs+83+PmxY6
SKaYzzvVYnBmW4FOYO9xCva2EhfraYC/kMda1HfLqlKTGVHfsbd1K0KfBvsKYDKCYvjJ+mWjc5qf
/XPbRinyn/UNc4ApnrIoPdJphagfv4zDLZjHwYztzx9nOO1PycEE/bd1qUBAuY/CWOewv3afZUOg
9ugdiPjKkLKVoxlUE2ebOR8gSxe6fEHXs35S63x9TwbPvA5NPgGanUKxJIN6cGCpOiRasoyj9Vsj
4A5XGQWqgXKudReztBGDIGqb8PQ3wnKVD4c+ttwhVqh1rd+AvmfLu2FwrBQXFLIpvoEGGqh6MFNJ
9U9BNzsp8Dvx3At87/L+3XAT/u752/oZtGKuX0XHkKVitGU9yvKKup4aB1A4EDv5crbsxD8pyFLn
7aicl8Ej9fx/mxTrSKlcD0cjO02ZhTNPzfzq49Puf3tCMg0iBvw+diZCeIqRuqhiiOOpRw3Mcjpk
otE38p1VCPD/p1bAxqCu5ftMw707UQJX+EULDGeChuQdaaKDBCBjiV3ftMdget3KrZ65sy9FuXPs
Bh8QVHpqd4h+zrNBwjTZvm3jcLEbKi3Tr4R/k2/IpnoC3wvd9bZqf8Fkh4c4v4xYqK+iBLK2UOTr
M1xC6fJqdE8Nh0/VAQ2YW7psEZ2GYZu24apOUWQJsZzXxmG/8KfaQfxQf+UwbiW21oxv0SFVPpxQ
46KZjQebwdHfX2Fh/7f1qGwixBsMKWki+Abp3+9c7DgoaK07+kZzNgw/l44V5CdnHmQ1F8RYf6hW
8zHr6nS6kwUpEXvp3ZGcNGfK4zjWB+7nVYNegICUdfp+lELBNx/IVDerRlgn6+RyAhUrV2Ove2U+
Z4BkkAE/yB41maZ3y7tNClZLgdfzpXnsqPOHiO9QkPmUrkUiFvk7Uh0R0et0OAcd6MCcYJNlvX7w
f8vhQmHIQExhUNYHL11FxGNGdQXubsy8kN2TOWZdXV00xKiclrZq+TVDHagzePKFGVy8gIV6bhgx
LHLz+XOrTupi3of1oI61w4VfYkTsOY7byNusy4rJYtzo0DTCIEPALSv5pc+6SM2026x46Jd4AAMk
NdvZW4zq6MKmrTxzT4T/xhLFSrw4+WuD1cO7zrRzFqLyjBGnq6Yj2e+PFyLi5f6DtIGAVgsSfkZo
5sNFnWNIvLJI7MzCBXZCpc+Y/gI6TfPf4s5F5Etk2lBRB0Lg6XAGbLWEHpXawNTzjMY6t9PKRdeW
K9f75sO9e5tC6zm6yRbVrc0W8kCajQX44m5RMX6OIa4CpRXYyHRU7OQDqYa4/83NuaXSP6/1JGvP
lpnWHfbHyVb2+YMtDhOcUzaLJPfB+OIfl9gsAvz8KZMtEFO6id2tAmhhsSDbpT9wHF1uQyRsXROG
L4AAs/OtfYYFggqmKZOocwvu3WdkaJJRy9HNMPH0wf/KbhnhSc4/n5MHoGTH9/xZrm6ePRdvMkIp
KmrPp9sab+eIYNsz6lPDccgQJVo3U9TuHUQqs/aefr/UtfJvj7Hdw9IYD/BgxKbzLCh2pkFIqfEy
2H3lXE7TPTuj7Lb40wp+A3f3P/pDCERNzbtH1MpBLPWeC1l4yPtZh5Fgla/IEOAv3bOypPRDqnYS
qDdyGtV4yii5HGT93bUNGlVwoibFQS4D1SHcw/vIHrbCjsiZznH5IGN3xlU+0jXjEYUrSeyx0B7L
NUIsVjChPbTjN0GxpNBTYJAN1Ou5FznfKA53YQdyAotFGl9I6cV/I4MWMsyMSc4sbi0x3n3b3GuI
8kcXR+EqC9qursnwMP5Rx/T+/+zwUOsRW1Dof14foQQmcZ9kLP2XXkyjpuUITzHlWcxfXpZp4iao
ujrJhzY3IjIgRFxg7wR1zSSBrE9CkJJHAtdYyURCHPYm5gvtp9jab/k+1VnXaIaYkQ3NE/I1IAOM
sMZuM2p+A39twfrkpGJxxCqI7e/9k/8/oyLzlNvWueMfsSGlPPYGwJQo93DyvIdJl87yuQRv9lYP
MQ3No9Ix5CA2oX6Dt1dEML5GMY+U8l12SEvJXdxESx2DOj50Hgmm48WuYKIom2i/Ff/KubLu0CmB
zeLRJVGK1dxpvO6iEm/gUglmbwxZxzSaazEaheSItwXtI3v1GS4Bq0EGyv4NMt7VbJNvTWK0e13l
PoRkXHWh+IXqbt8fCdTTg1t1d0Z2ZACCSnWyKqdYczVbbsfnhfYfLJBd87wDHj9TEfaXHoLX2Ecr
aiJlrnu6xDQjrWXOdMTIMhLmN7sfBBaLUsRBSobuD4GL4KSuEXX7+/QfNEwAf8LhcsX/5hDJukuZ
/26wjiKepN0pjmuH6my+ADFFc83yPeTXd7FR17WnEwByBXDXQwe7j6ybvHPufMEOeaaIebstfR4W
Wbnf+u7bMvgnYIolhfJU68y+8yoqygQHqg7KC8179lNe5P6T8azA6PU7onUBA3JzSL/BDKhOOYnl
JHF1Lg4guXmUUhQkpKnZJvy51gwiKhyxhz9vwKc5uw5Ed8XV45UNo4f/w1huHKbs/qqLIzjB0Nhd
FfkSp9jsVfYf6Hbz+xpQwRwTGBwSKyjlccC5whfSUOHGe0BtytTSMeNVFJYwx2Tp1QYcQ78+k+Cv
gnqxy5cB4SEFrwKrew6nuZzGuoCuatbdgIg3Q2kWVtm6/ReanakaR0k7ZFH3Zb5kZOU4GOynALSV
OLsDULf1A8Cc2d5jAePP/xkvxZhqP0cr6t+V+/Oswimr/veCEg+YZPp60yYYRpAkf/aJgOnFlxG0
EJzpad3efxTgGTcPBjVn7ankvEpwn0bTJVw5omrLm1OfD08yBLRlkGvzMxbxTzqxbolJUgRiZyBg
hLgZXikDb1CgxB0GPdbOcpl4WpbycJMrn9hv+Y5xmu2ri32rkpbq/UTEQhvoTm62gCc0y7j17Mc8
ryi0QmibgAtIvmf/ritiIprBtLtw2UAgaWwZiM0tM/5pdni8XBYpj8BWSl7WKRY+a1UFf3jHbqDn
u492d2WVbeFMAXLmkRBVWz+S/pa3d7oabx2yR+JmyMqfCPEF8MS5FYIcd7o0IathQkBu7lZImsbx
NVkPcX7IEfBRVYPg3K+ExUvaiYUTnxbe7HpS9R8PH0vJl6KH1gGO+mQCTNHmkDY3kOUmJc1GUbg6
2qehmDt1QkBueYIPDAryfVrVNcrPILRID64/vkbnzi2/k5ZlgBceOpGe1NcqSonZ8HdO6KPJtTNI
5pkjTDWwVBzHeQNK+wzl6dDoPwWJumxrwoLJSDgdd+dbSHsALXu8bob9JjMYgaahwzPMUgaa4gt4
Eou8nh2ta57HhuVGcq5Ctwo/gCUe+eOlUN3YlLjBwzZQwb6207IXygqLsPFY6awsvYaGTMNcimPz
clvZ+gxi25/hJbVrhSOR2kUbOojhh7C8jtHgOF15XBVWml5EPPim5NaVDiMjpbIYIqEy4jNAk2jM
V+9nuybYbPtwyXHMOcDzJzjtQZ/yod295nQo87jmX84bB8HUd2MzpsfzENJmS7II6d5pIL/jbccP
qDszCstenDtKbqQlbTnF8dwX9aTMquHuvPUO70irErAFE0cjj/ukMgrF2IWnb66nS9YMxg0J8ylE
I8ItRAFNjJJ5clMC8U+IaozxtDEyt2n6BSW04BDeO+yNvs7dFKW78RJhOVyPLHelD4YrwAZ69gPm
GK1na9os+rB5g5z44nBM8A1h5h20J56iZvewe7YVxfTFUSKd75xHywZv/EJI/yH9iMYM4q97XU4i
MyOjGMQ+AuVUkldKAubTHm3jx6I2kzIvB6/jU8Tj8VuJ6iNmkLnvyGcHzRzKX8eXNtTOy3cSgL5z
wZxYGfuFOclZvrkLFyMekRIp46xuc9sjNnwEqtcN8HrbnS3Mdmux/f8q2BBzh0LD0FhdErPAcf3H
63b51eLQuv54qHj9dsmsfSYVVYPG4UcnrOfGFb3pYYkjn515vAb8qhQv2PFUFH1UyRqS4Kf++m/X
PFJexI7V0nM17DhYriwCNcki8gkSxYLmxATR527LvlgS7Gt8fmCLLCvAuqu6KH8Q6MjQo+qVPOR4
JayAgrKJR9piv7YUIMvwvhdF9q/c9aesB865aHmcqcPd/Y6BJSyQdjfAMHV63xEUJ7QavxfL5xOv
Q1ryvWMgSEO8LErWXSXcb8QiHmma35g4xoARTNTIRCuyAq59HciyLpK+lF5I73uazRRDdD2gMvS6
iOEOyJ7uWgW7eGCl7KMtWdfxBmmiNc/fJVcEVJ5+oRQ7zvX53/y7yzqOCQlG0yoA6MmAnRbztjKh
OIroYc38TFtt/Ra0z5fxBKnxgZoqufsGdlwfTjTatguMLkaYgWkrNEQurg1iVjzi8CS32sLo/6mL
8nl5asQFgvFajLUrXiNk75KuohCp9AXgLPbcW7CnErXiQuIlY0m5dXQfJRT8cxMB2iGk9xPhwdnV
5XIUoq7ETfTHWSh67FMVji6ZVqhLwPmuDqD2YJr8SWue+vICkLGQY8gRS4bR7zda2qPbghIsvUjM
oiaAymK6O428YmyzSfNn8/be/k8L02yQO35C0o+m23w0pVD9bOBDMXn0ex3QYS4y8UmdtxE1eLhz
S90PVGpvTjHKw84BM8XmC0pBswpL1kWD5HKkZUM7U1hWHQDdXNu6ZTG5udyn8aYt3t8AfmVTByi3
w6ql3JxArIcLKVrfZpBFgL/FDyzcxaqvFnlulHY39l/6CpkdBno/xsFFn/43hHt2zyRflaecT5x4
WzdIpfZZGCZhLN95gvpYZdOJGghvVS6aaygAOpdF64IP7WtN/QCFjvmOVzGHEo59Tl1+vyRWWJPq
io0KQdKJ7MXYryv3Cvt2QnYdGwy9+4ttjwiZUXUItollAvIq0B8jt+TFRBBjag/gtabX3o849u5X
jgRc1izhTMAfv6hQZbYKRMaQD/LPaYCPsTsDshe5Z3yXnTMa8slbEdYagPQvFyu4/4PjJvJ6km80
IJZl4YQctmuj2yy1isZayXj6L98rbxX0oA2tZYq0fAXcByrknzlcF5Ho9X0mzCQOhX8ioLFOHyw/
UNfqH0wrhl5LUdIQgPKAaUF5FjoV8OK+Yo/rUUIFO95SP5nEWPuomeqjqccLYRRlfNqDNPDdJt2q
oJrjROopxI8yUwINI929iXCgX4ZgW5mpJaxxRwaOf3FY3eWknWP/7jZ296Zw/e8RUNOmC3HMbVWC
7Jjir6p1M7kmGzrrXzSkQ9HTadpP58cFb5P2I5j0aviTce9DHWHu3SqXko6E/afnIVQTywHe3vp0
eSOfqekvucwydtvYz7afOlfQPLzSNQlz5Ltc8M98pfDUt1aCOD3f1w4ae+5qu60cbuYZet3ytmSG
V7tGjUcJzK4jhN8HTfTTTz6IuisgyoZiCUXRpxKVzGLeMQybIAkhSAI6qE3cM046+9X8RPFjqqgX
0PU1SpccyOhkkV0fwZ3AJH/qs4F6499mATVs3oFg7cw1mh9VPOw5XKkAv+dKhE+O9tcVaup+hNLQ
E5v6Z904JrLQ8g3Xkw+Hjb0rvZ19SOu21Iqh5QvzufI17FilcVoT/1Dv0EJ1LZwDWUNc3SHgdU7I
FgnKouphwdMqeWG12BpOEMQuK8nqBacAy+//qVmWH/m1Qe6ipx6jAwwJRm44WNRRreBKxx+Xt6l3
4Jm3a+GiU9aDGUdieNjAesLR675bCvhinHS/00aRzdyHUSUhER/UULBJFD+OvYXnAG/zr+n7sZiA
fN9gRinqGQSOB9EhYYEb0adymwN1AIYgTW2irpnb/KPmy1o3BFDIGxkkl2yXUq5wc2cYXxeKjq/D
pS+EPmzCzPgIZNexHtDnXnFd89e2UxIyYqSLSOSKxloe4ZJPBzy5UrhmxnzheQqKTIS1WHtQfvEa
oWVNOWZP51L3gcv5Ydp3sQyBYPQLWQTARUVrilqV8lb5F8omH6AF/cbIz5gnzTpTl7dOu8pAFPdh
Jlgdxsb3w8qvNxkrsX/dpkObOt7c9mlcmw0aa/TzVbodXBKaT/4Ggies2YMst1XcJXuad6ds//iY
3lsP+k25oRAP7tQsdCcm/LRYNLNUjBFXTf4vgG0WL8WAI/Q4pvQyYR2Ab3C62yDvSGGbyc9oKDg1
dtX5eLhNOEwElZyHeQ4zVmAeFnjSGaRhLTxGG7YUtPI1+cGqv1lpwOt1/Hv0Kie6yDvqYo2Hpu6X
d806U/lFN+cFeliGLUgvGgXkosNHnJr6zEtnXLjHpGJPmTev1lYGKRUYSwV7eGZSVas2k8sL0xWH
l17e79bcAnsoG3my0jAp0hWPYaOkmWXhsvqLewx4OqQ+IS0mtlBhcwej3L3WCLW9dsig/uUvkwLh
HQZn3K8YzMfsW7mv6arRmnF5je9iCbRFm2Kd0pUWv//pLuWPLL63n78Zv/WVg9RQr/NCK0XLfCO8
UYOUC7hYwL081rGBdgvzz+GEA9zjQ48rRwohVjKde/A5Nni5JARNmc2OaWQxFPALaDV2ofTyoK+r
5hQtmEWCQ7uwie8rKOXFpZYwCUrIXjmr6IcVJej/bRg42HV5Dx0wALmvfJRgv3SlEPfm3hcRMKGX
ZeeLYSX5qZxDYcVxYwJqahzSPgkWTh/sl3Ov1RszQHX+h0KZUPYQBUQRyEaf1Mgf0n4GGx0oFcKL
xXvdD5tvEjnoDxOWIlJ4G4MdC2dKsLO6ZlMUtihwpIuzUYYVqx9uAdOQBscfNJZLgVWAIb8KudqR
hGA5jRB7XlROZ+YRRGeXIkmFrwc3hQzEtuMRKYiJiU74L8sWG3SewYiBqBBEKKnqGJPNYrwzQLxt
yjfL7vdPq5BdKrBPRqPUBStpZ5aNRLPPjobe/rSXGfbsxglEAk/OkuiMTjwcs+miMA0Qz4PyYg0D
kay+8T0X8hl8RPYWkbboBPcICjpJB+83QKElpVyYBthfTgKFa4oQxQxYLFV+2TleHCk5MHlZK1zo
SBtWUqMDiNdW8Wujg5JgMNqXOjMOnMjFPSaJWVOgoBlQdfOAlgrl1GUb8ZmLqE4rV6ymIZIjAX1R
zyT1kVnknGiXBIlbfrDtlxLR4Fp51xm3zqsiVCEEByKF4j7JCINUYfnqDSMIqKEmsJbcsjYiTLgK
f8J//CkL2vfwBx0W2s473E+2zvxg7VsWVDLo6wk3GuvEkHLf1RmSxZ2thAhQOH8GEpF1X7n5E2yd
dzfPZs4JixF6/xpafL2sDVchEloD8EBubyuf2lzK5jBYPe/kY8y4QU/ltquVJ2SNION0fvwZXMlG
3ctmD3qdVh5ibOTR7D1EbJRKHGaS8vCBO+/jzQ91PAjSc1z4Qwo7y2s7xaYh/etXhIYY3u2qbJi/
09pyDvM7JSaDZYF56BQrr9hgEpV0lIBbAjA3YyCZPhmRTyLG2F0GGIGOdoQ9yRAbtiiCTnkfLeUU
J2hLTP+Y9Vcmgns/PNX4hG0JznsteDpnz22FbTZ+L+eLxLcjWsNQFpzu4ivqeChhds9czGAPyWvd
aHQPE6Sbm3czpSXj7pkeWFkijeKH6E7l5AgxY5a4FXGszqViptzk2h4etprYVRZZMcdl7khVHGfj
Jbk+sMRoBwSGYxum0p1MxVLaG+j4Che1gTJ6BC5yCpnYscGZJI6boSCUuNIb2tCFA1mn3027B+7t
HGhpwxBkQ8L2J+Z2NcNdEfnD8JLiP+4Do/tULQ/zy2/MToJWTtOh6Ge4Wco1ey1pb/TrOggIQdra
+idIbLZp/Vco1Qrre3C6PVJ9Wv5AzCSf9xagjDU5Doy3stuFgZ8eHmTSf6kItSEMO9tucOCimOrq
MQDM+WX76tpfwMFh9IjkaDiMNK1g6mO5p513LoaP2XiG6z0L0i8DnSyf9NHYoM9zdq82yHbDp26p
DWFZj93Un9CvZfxuGNLT8qyyZvcaWHceZpjuDs7UOqqHQACkyCO+lZuS5inOTuIhHclTJ0MMnl8f
zrBP0j8G7bkn9WM3cwrL9AzN28cYW+tzsPYuqejDP+guPVWVPXNpq+4So5ErHJaD7bgb8kMPS8C/
XNtvO0gIRle7pAV0OZ6WhdxCh6S/FDh9ItbH6ppGGPg22SY6wPNxwQx5GIyK7ufzF2AJ5sBnZw6M
jRKqoDk0qga8XZ/g4KBsczKmqfDYSmDE2ty6DAAmQ6uozuGrc5S6HJzk0nXfOeDvpv2mprlU7NIk
l1znh02ih+sYhR9E7phk9sT+rSR2w/j38Rt4O9vpLTerhgwYvnZ+KhhgBiz/BYW0LhW9VtrFsSfs
s3nxNMZ1LqYe4sID62z2DlBuOo2uXQ9UG0y1mI2wkGnt9JSP2o3/HH88loH4IfTbW4SPeqEamSoD
/rUjIYUjBQGUFHYcIy82Nm9jyPAvvGDzeDukltLsYPJbS9vLm/Te/R8UmA/AqPb4PUDIKlP/Tpv+
vc8TSf/KT4sQ5zpw8AKPNkCS8VaCdM6NE293iikvFR+vyfWUhYlA/RbEzeXOaMmCQ3WutOXp38rk
GdN0ZuoTkpoWLRxoI2KobAQSkpqQDUvxqgjgtnBItue56p4ktU0hMmLVXp4V0n+ryVDNOGliCNZ4
OUqv8/EjEHYcnPsi+e5gvmwcUxghWzWg2m0/N/QJ/915jRsJc1tEWS89SYMrlnJlCJaaF4OIsGkl
mSjJjXQSEbgYp6ZNxbISaIbK+SAAGWWlYAsJzAyvpZEn1klUlmuip2SPJHz+kq/+4IhdoumF5BAc
7lkSAUnB8gGPOkrXGvONifigo15GwGFbfZAuuVy1nK+KATgRDR8cZLMflvOSChYUM8Nw/i+0iTrd
AlDV97tc0wWh4Evy5sPj4pz1crOcChFn528jNthXPyEia9IWXG7j0NMIJOFK9YVhqxi3XImIP70X
9eh9m45vMr9wzUeHS4AkihCutKQdwf/EjcoBiCHcxydk7/ICoafdf3nyDHBlaxpsI+NniguaVIm0
P1Xi3d//QB/+GhlcOsqbnSEnqEQwuTyj0Yoc25TlMneVSg2asde7mt9IsMJ7DyHH+DMGiN0XyND2
Ifa3dyCuR6Uw5UvAfBSkMi97N+4qt5R88UnHoH+6XLDiHL8VpPcKL8NLyseHjn+J//L8WYosUiwv
ezLa2qYh4umpljU3bqcTfusykwILAFqWC5OKUJm4+cp6UreU1t7VuJ69eTX+6u8VltgOqwcbtIGU
Q3BswlJKfCA3J3ysNawXdqL7l6OZicWpgicQR/e/egYtLowgq4znQSmDYYV9WWH7fetP5Bg6QzBG
ETulSU+T3y/fiC2IXAb3H0g1yO8RgM0zrgxc9YD0DK1ZBqP5U7Ko85uSWvZU0FlJirEY1pcHhdPK
Q+EKVK9KtB8BHti85ZqcGEYUWp+BuQ5FNBoIrXemBOXlwjwxhoQ0wTy8vANjJ2huS2eX7/AANXq5
UhGd9hqGiw69T8qWnCSHdFscn3/O1YiF2495fp+Xpg0MVVQWXmIsCMlCNlhLJQ86hrw4UwyJwBkr
J0RpXdCtdyi/T3ng0v/rww5Gsp5a8C7R1j5WfbahlzhVVSRvXrEGLn7CMlr+DEuTE8QmN4Tr2l7p
xsUNd7H7laxG7kNZwYLzLkZ9CrSZ+iclOdeZipsex6i7hnA8T+RkqceClErN5S6dq53BOy4y0Xqf
hE7QrKIaSCevNEpweS3qDGuYFmlybPg2/6s8B8QMPVV82km7dNctkb7HuQ+dCq+FFcSiPDk96AhW
FpAv/k4H75Y7LaUbUV80XwCA3ecgkWND4C0eybBuL5wAOAIAH++yhaIEwZOevxPDfTY2siuNwqQa
STSUTZ8wWtbbvo38k8B7f4TinbW0gieXGK1B2cLFkZivO+qb9E3xsRu1vZ8vrXcp5tB8a4cA8lDK
6aXx56sXbnw3fiPcjBcJxtCXHE4qxIvzkgJJr4GtXJNsryU+tU4R8w4vCA6lml0ESYVN5irh15/k
6nBxjxoHoX3WB9S4UqfqsiWpu+WsDxUoqTzfEeO9ETrZQdrFHsHxrH7TcO7W/uIFtGRSWgAb+tSu
lCuYPGBzLdA/cXYyhKurG7heaFQB44JubpYPctQy7GuYNlXrLVLt7eFeCoKY2spghNj7xCKfBFv4
SyzKntyenk24JmlRtu5GHvnqgFKMkGEoCgAV354kQA0IPx63uOEzJ97qLb/PaRAhA5+gV/rKS6GU
me3+LXlgN0N2tk+AVFG6AHin3VBFnJ5IK6Hsh0684+fYlpEHNy4BU1xSOCRWnRvEP48VWsP/YzbO
Yve+0Op/8+PTtSG/0dfNHh+7GsJYFhzlkLh4kZe8N0IC06kTeuYfXPfvDfsd5Aw4SK2vlpgA2rES
u+SPoXbRkMFnI9IVTy39y4rhWLt/0WiJ2dEqIn7/hWQ692ah+ZV2FtI9dlUOr1zPYixZ0LDK190f
CAul6eJ6yxk0ZtHyx1nHe6OlXgXJ7IjJbnnyP5kgn+df7HlikCMw9k7vOTnDPqw7xG4LukyAyV7z
32BVts62mIGHjZPNvxqWcyqS1Kr9g2qSEsrWqLTaeMFBCUsZ22GokqUQyEtmjKHMz3Yt6ozibg4o
3Df12MVuPJ7pHq2H8JoOBkYp1d5m8JJBwhEm+psFa4mn7CziBp7QkFWPuBAzgxpalJkSrmgOWlHL
oqXXb+hA2jlWiI/UBilSUXfZxq34y7gv5flZEMLMd1yVBX4U2QKjZBh8F1RSks6D2Y1FwgysFC4M
Pu3Qio5JnxPlli97H2LCbR6r94vMchcQAwocWAWJXiKSQNF5HPbV3aeM0qHiFhC6gFSQbMVcRDXm
SttxEDLvvkx7fNlAljhwe43112m8Q/C1mz0SlH5lj2tienOjX1DH83JL3soywdrEvSwJIV00GJLv
ojPNA36sK9oLxQACR6BDMbx9nJcAH6NBB9awnJiz5d5oPBJlruMiKmUCdBxXktMk9vgIepPj1jog
gAtzPbxPUdebzi/cG1flgJdEzgzAUrrwTv4M+x2jYSojsiaSLXX5q0WqNU3MN6wH2SH0o5HLVW5O
eAnwdF8KMIvFSz/OlfmrAFPmZ2tTb3ygkZbDZ30GjovXA2w7d8Xtl2eg2vMP898wqV+oMLL2eQ6T
3H9YTwSPqzAMMihxToDGloGH99ojoiwX6RTfou4ss7cVUGFWd6w3Qp/7VGjRa5+gCVHSvwtkR/3L
K4wiSTXVmNEGbB/EQG/eMpaBFlLjC2ui8Je+1sKinTPOWcE1QzLUT20rmpBC5hdgqtQcEl+pJoRZ
Y9ZzMzzGYotGKGKqIVjughmFlI9K/Cb/xYFtXmSM2M13KQNVoHg0SJOXkW28mISDDBD9/jXt4PF3
BsyYh8Uk5HLRQng8xy7o3yRbOLrCxdGV3lx4zXKQ1AwrlCN7kieSMrY9f+kiZ16JNVJGrc1hE+WK
6wpNxKaeX2d5F6YWanqy90WIhvVjf6VeFqWozliyZYJQ3EPqm7039tNznKrH1iN8TZZ1J/sJ2vcU
CXlq6QRsM1t49l4H8cxxAoTIcS12qg44LPP4vG2AC2vPO2HLev1Zxur8co1YbU4w0VSYtfl1hk2W
/UzjEekfJBLZpx8ch9GVBIkYAU1fFTXDwDCxeilOZ3oHt3/8V3B62IgZ4X7SOhK3VcHt/k8ba09f
90zhO4alAMhvdeXZxjRb3iKWi37k2Hj+38I11mPnawJvnfSc1kHRd4H3lXeIXGC1bKsTxMphO3RE
lPkq2YDQNzQsKOsEmwJCSZgctuRDBrz5BrWJ++hbtdKlYotWFurS9IGyF611E/4N68p9ytYql6pS
SYeiMasLtNbMf3ZrBLR6gyETplhnDmDlgIkKCIuD17kR7MQSYDMMtrV3+TaQC+IUVDQqWkQcnmxn
4Eg4IcRHTfPTV6AEfNjghKQPC31RbP1I1t1VXoAx+2mNCBRZ484yeyfsAg8aAvwZOxU0WHXMnATf
WCGxAeqWawNX4jVW/JxKsQbCWoUzR/RZKpx6ATAgAJF0+Lbm58qU9ifP7bNXpOZpxStJ5J0+A3ip
H9+FSf9G6buLsYfUX3AkZoVjW/mE58pT5qO+gjf8ob62vPRR3A39KfP1O3WbXtw5SYHXxp0dPcRr
mkSkJbCp/8aYkVpN8OsDUIu+slHoo5FMYXbo7AkbsejGtWZa4QuMTkDrVSyLXvM4SXUUGl7vvR0K
IKmwaNh0bagzT1uM8d2qIv0gFRHTuUfluYiC1/PmnlhVaDuJRgLfuQBrKvbLSQfxIGqg9lFhJYtj
bZzcBBTw/jHRwTPtQsBrVCbgO/QjtIpo00UTGW6ENIB8Pv30cGKRf7mf7k3nGhnXS0NSN59dZlsM
VODtuaTPI5Ixi4htmBCi4LM53U2LxccZ3OOi+I9nD9081KkqUJYBficRX6NgxXysUV2WgrPgCONY
WjYK31lKy2ujpfL/wO4bsRKdODo7tJzVkwSwTACLxWXRLUb035TH3R8w8riwdvBSF95dLnCbgM4v
x9F+oj6Xo+WoVU1UzfEJ5Hnz+5NYujx143lYIVQn1XxKE3KatcBd+RomjVCG3WGDI4JqNtCTE/ru
TSkNrw0L+fC10yWJGwL1wEbWTIumPu6vjMn1V3nJ6H6PFGMQGYvz3TA5NuRmJJAi8enqTegEM01d
Ot8t0zKRVGgfyDbXl6fPogsW72GbICnviiyYk/QqSdgiSE6qfEumv88yege9c/2alPCfF7W4BnJg
f3Z3VAV/xEVs7TCU+Ctll9iJTCJ0NBDeNLJa64bB9LWwuJ8EURnhTBzLlAgMXaHr/OoDSa96tvu/
dVIR5Wv4AuiylwK+FHlSHfeMvUc3Yci7dbzJSm1s9vH2RcMQkZwcz10kbzBS2dRw8nugLmgs75Ib
z02/WrnrI3yG373hC+vJ0XzuAL1RxPuKJ8ePPhXFyDne+9/iazaA2Cezrb1GM84C/TGEvnJvuAcL
i+thb8YYHcbiKhdZgIatefVe7tNGVeE04vNvIIgXnBgKnuoRFff5paYa8NeRvgDPTfjjZGPJwvec
QuqppPn4PwqJBvTFWASsipMvkNh6fin38WjteOOs469a1PLx6gIMbxWZCNvNSOFcJtnYJlTMPzVh
I69eh/wgcRhMsFI4Z5v5a1jRhSuMykf+/43JHhlqOHYtjmveIN9dS87s6IDrGw4Bcbyo2EbEmPaS
jowv35LKdi76uiCgr7SV1G849YYjvlndbu7zuouU2W74w62R/Rw/Rct3Jg5BDiLjJZPUmqm7KhXm
VaRaWfIyDqGCTGMqQf19Gyx6FbGvgaCgxth/k68VZXDPtOAqbZWrtLOCgQBA+WCKeF90q7L7VAif
i7vbA7LlozwIEPTbFtOcMdTMq1Dh08SCsQ+WnZDWqHyFg+yQRnbsML2rfoGd0T8tfHLVSOzjIMwR
fWXsVQa1/Fmkb1TrQRzFsTx+4htZFtsTw+rCnmLhuYq9aughqX22oFZGJIEMWS/UnJ4CnJnqNQ2n
zmiarzT3tcCoYA5kd0YjrAWFEP/5pmMzNyyPQxfyMTwNkwVUTPXTFr7gdl9XXTlKVl0BEoQCQSA2
6k6GfUa/jjEaUog/7gr+zR0k10v5Q6xeSoLGK8K0oWn5zM2XmMlY+vLTzxQcWc2N7DIATUfoIgJz
l0b77nYPTbCZ8cMYWTAoer0WQtPCKO5h4Mx86qJCCI2im43eOzcFuY39fp7UMneJ+yfblxyyZBli
lq22PsRGmdGrAqVjG8wJuzGjkPiFm3rgQtzOj5dSu9gAv0g5jkBNWnWD4H74t0BnbPhDDxoVlW7J
+YoOBRQP1jbAMQphYAwzOv3v6uLymuqelKrAS7RdZsyeaFQ42dZDksx9mXVlMItXcg7HbxQiEYYy
WfbUq9UTH+UjXIuNPR1rijMR0yWKEy9gI9sLCc3x98WWSo8pK2jhHEhBuH3sx0HiKoMSiqG0KNy8
4YURNcNCcs5Zb9Ea2sgbW4IfkLoxLcTAm6YkTbnyPu689AgJHkDXg9X5O6B8cz4Y7uZyy5bwRqIM
pKBVvqeMkwMtIoib3VQ1Std8S+gMfvUe2i7Rei2PAFXHwOpNpJX6BdatoIelJDwlxc9ASkdv1V9b
HBEuotqLVKgzz0+TFYSvCYbgryAGqj4ZETWeV6W3j+Bn2EdIi9MyCT60zlD4WDppqWu3Mh+czfJW
hXFBqGlFyUNDk8krnEX17o4gVP6XvVsy4iyw1OY0RSSZ6p0P5pQZidb1NVKgCa/KmFITbDbRookk
6zfJa06KkUkAhnC2PKFcsJXsukXfXRE1pOXKySYvRIJR1JPhFGxKwHY4G1cIPiTcaipKns0EMzaB
oggQ1EdnGk9aUm7EHeF/7haOrHSkoa3lavaro3Hp0mX9u7Wk9a7MNL9OU2+UE89EMZNJ8pzeKnBy
H+wQmxY9JERbXHMm/mp2jsxBkGYO6P7QS5ACvb4t0EH9WXRD306PmEVcOfPcowaSMP/YBinW4KcA
qf++O/OA8sjniLKj8H8uEC9AeddcnittAb8QhQf0wLRxYDoWFl0Zq/bQ06GVjS2sPjObxJgJk2xm
mJmy/GdGJ0O19oYNdl/k3A6qTIq+K2KfCbEgz9oFGPn/vzX35DQixJ1AIsmPu27leXQeu/tiWw4b
o4I6n48cxLm2nw7G11Ngt9mW9dj8OuOHhMyQ9VwE4T5INYXIO0OnB/eHWihpMM8EcHZlaeNo7KIL
ic+fcHGQtAn36w/UQHryrswoNm5RlsPEMHVp6lCLs+F5Kgd8O1zwzKDx2vl7jHvpfqJmB2vH57bc
ZUiF0PBCjWm8mxbsSg8xGXgrsJiTbNMsR8Zi+HZnhHEHnNcH4uzdRArsv7VFwHFsD6edoraS8lH8
3RG/2HdGkUXO9ZRQRU2fhN86ormd4NuRhJLygKUjBO3xVP4L0+7mamJkwUVs23TNZPksEBA1zqQh
F1Pvpa3tLNyXq/zdBcDBfaMJ6YmW8bOUGLCzHNxV8nh72Lq5/qJgCSGveMEKT49rtLmta14IEqsn
79zuXVvlg0rALbg3SkwaYg5b8x4n0gRv/2U8rU9s+QKJcNvVEymBrq491YTJM8KYiUD8sSgYnjRi
PdvCNLycHVY/J2XYTfD/Yj/AcCRQ60TIWwq0030Nz9gu+2BGiadlFYo2teXZD6UKnjPvljCMJDfM
xVSnMN3elFuTLSP8IqshV61NG4vdaduqJ6Ug8xb3nXSUqwgHNGxS2PLWyMthhPLKHUd0dQob0ntY
A+eJXWT+3LO7ScbJojfkXJxfCDR2NMEa9Ya8hQkSeE6wJQPkiz/e63UyjbZjU/lw7TfTDqCRMbRC
hRT3U1WWPlKvmGRUjNm6BwBFeJLoSWVF2JloX+zuH2EV04Hgh4KyQzXOL3f0QTCKQYLufG/HblCg
+K9ql4RSrneHx4cPx7CFjyxbqyo60lSJiAlfRHOXVJnJG7p/BhF82cBJpOeDhoj91QiWHVzpkDea
FZiKokMP9wFpAG07WmrPXOFl0l+ph/m38qPq+WWnQ2SSdw9CzY0jnEa6XiDh4qxuKGpiM08Yqorx
DmrR3YqYKuaFoJCcML7TiWErJG3a09Y7DRJHWw7oshWnoy8uzI6V4EEjlNG4pQGQOC7xDq+5TjVt
rvx2eo6k/DBg8TeqyjH6w5w4KcA83MABaFVG0UYKIF61kn/S7L/nNmsu7zFVea70pcEWwhiYiv0p
euvJWncYgxlBbDrH7d9KG5BNMF4bOg99UGWXd+sqgTg6NzpMZoX3wE4YtMOA3ecy4NdnrhSdumeg
m8TFMWNwE6iuTsb1BgYRxa2Io8qy/g4/SlJSf5kXabmgCaSChvDccZTqEEUaw3q0Ph4F3U/boZyl
aHQscSC/VDFqYbrvhlsVxrR3WLc7GL+T0zSZ1jIiSyB66awGQCO/c00cpdWSmMSMk6E2aoR9MNLW
hOew6NhIsfK+aL93Lg3OUS28gT2S2xCHRixjCRLqIR5ZX9zottImZQ/Ih01+PEMOTreC4pc3D/Yh
nTJYSc9P6jBdjp743F9I6ulRlKukr+rXJl5y0ywKx+HUBpS3NVNCBVIp0DBP3ltVZHF51wABKc2m
2XjD+/RWN2RARXP4WSko7YYddRCbfgp+ow4oG+cWuqv5LhQr9k1LrFQ2lai57H87JgLCB9Xg5RVI
yRx41ju7G60FuUBe9EUokCR6cai/nYj78jHmGIKHgJcJKQDPcHlJdAo4pKbQi0ivaj/4fl05bFxF
SQQ+TXYcWS9xMzBzBOD/pOuKz1aanMCnfCSj+xhPUm++ee/weO7oDmfFBuM0CR0lfYtmcgl9AN0d
YEbaCe01+OxLjiMg5BcjJFhW+6J0UTtgNQ8X6P0zDr7BgLcknRdiuK5PM9UbK+ScR3cmmaXON74L
BRsJXpqJRApv846V4mpubYr8k7WSGtDYL7M42cki9ofZGzIKqmrhvYEzMx7t4HgRJtnlt+Kttyed
RSFhUSyyMTXp5ALkBD0CMK8QwbQ/XWpCJR7SSPIkawFJDl5lbZTiLFsai7/N4NqaSugqXK6rMv6n
Ys4L1IP6VL3SH5s9k6qVdCnzUhveDr1rKm4R/iy8vndia91cS6WBlWGfbo8/eYq5grLSMi85bDKL
up7jKtP0Knt9+DcZ9MItjFdkKSFUY84vWnYPy2+BoLI2qxmI72RrNjMWaj8LXHcpmcyxV4uep6Pc
ssJI6lx7PJH8IPSqRi1EEGRoH73jzTGP+fbW+yZY2FWWNHTXommGQD6loQxOXzef80X67Iq2S87B
UuwV/uezmkL/nx9l+P1j9aAMEiOu1pbs0/Y6PcQ0ERbOLbewUOWu12aLxRjoN9Rn+tjrZBjVVZKn
QwdbzNtMlGMnyTKSlmFy2I3nRlgHQqqWn029U/btrXDI4r9DFAGpFbFJRdBXlm6cTi35vPRAYd/A
vEL5r6w/GOfXxnuJ7bqpkkdUIL/hmUpxSam2fLQ94Dw/t6cTb47unhr6GQ7cTm57GwffBgGgQrna
FR+cWud9w8n7cC/uhiTC9FJpUtzK36ZkSEc9DapcoVik4d6sQQk/CvPluELz80BcUx7wdrZqKDvK
E3YrrHuRb17oN3F46vKojYnxTNbUjKN5K0/9NMGuoqsoLzIDKA4SxD3NrFmetJw+KXhLKl/j/aWR
ShFpm7jBnPC9PwwaO8NPlRfg6mpCzb5huBQOl3w3QDHrPi84mCF1Fk6R0/7yAxvei9lgsu9HVMWc
709ii1gWJpl9J1L0xOPon+zCu0asXLpQVznF6SldZ8WEZzbCFrCHrgwVhBeHBMyryUQUigd9993X
Bk5LpOuUrVm2X79kOB4RtLW4gwpknP4uFy0/1Tg0E5YmpouwlHAnFJjzwaR0RadlMf2IwhpSQ36q
rV0JhZapMpfzkP1XTFtth4l1LszDkPQqrSCGDTYPeVjDbI96TCNmifU6OM013ycp0q+ZEm420hrr
CwpSA9Wc2qf5UA8QzyFtq4Aptz7OK9vegk0J+7dnkimBLdHWdKBkdG1DZRTxzN6G+uT4egRwvytd
ivDuxJVqpfqLtKJum5Bp4ckxctw63t8oIaDEF+wz4+mGtjQyUq5mltLUGeohChEHvArd8PTv3Lez
kBZjsaoVI8owK9FFIgH8KbetBF0cwkDhSHOpZWH+cBLg53EEaY8kOfsOfb1Ynse5N+y2RuG6V9DJ
VWnFWSoexWPcr3YgqvBV8lDhdhWoEe2gYKAxK2In2DZv+mDenPrxjgT4PsZ3egD1+FApXtI9BGCy
6iRNplAYP9QUaH5Cja4+9GfUOj9YaVNQDcMlA1eulPytD7Wf7Ly6bKAIfDk1Ul4uMsi41+EK8F27
eTnyuovgb6CWZj7nF/Y1NQntmZM3SFuII6bKZaJER6oYn9MkdkcFveGxYbwKIWvoY+6qxZ9m5SQy
N8MOaH8sZIQprJHr7DaFA9/XLc9PTNZTiy9vBeUnHtDDokVrZ8YyWteJMUqls0Km+BVfBV2ei1jd
BLNUrO0mMuPjWIuczHxgWgmV2JPFMXzuVNoBjIQBUpOSblQhnAm9okJXeDklBsmsn8VWiAk08294
rdwLz67kVoeuBLgEcnWFvKCGgJI1rklPvRQRDGCCh+Wib+nNLdMnBhHBDfFm+gXtXY1OugKQxPjv
Z+HxannIQrP8/udvJ+pndUgy2gxCGnGX047IqEY+U+IRh5o+AfldimxndXRRIl+KIOSyVylZ83/K
aqvV9ZQbkI+NQf71lLI9LbnaugT1oZiBUNBANQFyi4aKWJQtCw+RaDrWibT3Y5VuUPpLGibZGXfg
hXW5x+fga65LVKNZmAB/DyGyh8awL4pp05SjqRhPGc20jJw0DyQ1RMAATICdqVtSXSHmKC3Qg91s
Nu3cBCdCQKdKLjPjKqxzdn2DB13NgjnY3LfRfoQP979XtbtiezPIjgy9tqx9IFEgSuQvsE1/xlFA
TyTM7w10A8RG1DuggTrOQwFcdD5338HBYK8/CxwO5K4cEyYrTJE32L3PtNj75LUVggj+vPgnTV7R
dvGHf81tWdKMpNG4Jy6lv/XKV4sq3a8Ve7gYlzWlitfhJF3+F/Fd2oVk86q8fcSZIvzfOOZ7SYuA
X/Wy47tdbp+5aZDTkUHXXIcvv6vtJKX0w+KkKV6t59dtdZoVKQst1Kv97h5a/XoAVPUsQrWI/rGa
dCnCsXHYqtzOAz1s+EkCQQIlHRSQuR972FSov8dZf3H0USP6ZIUoz2+Sih7suhffamYHUG63WlSW
yNvUIH/Lbg+dBedRzWDWiZc0Q0+7DQ5oCG2PhlRR1uAkvW+MaY7kAA6mLAW8qyWtZytn+InzaTAQ
e49+HqTuZ8KjGwM55aVCfEPqkNLVZ38PVsT562MvHayBQfCsyQfdVYivIBSAx/mydcPuXUfK9f4G
znaDMgRBQvYGaAQVf0oCcwb5ry2i4wYfiEb6okJuMeeX6Vemmsb7njE9g5eNFB/InbXpDvxwBt4m
jUWrZMnXoPDpd1OSLIVnspOHF0NbwyArkOfFvMsq49KF3rTMu703FRkwfcZVwBJfdy9KsmWh9J03
FSfLzTsTZtJQ7zgCcWoBfxLIxmuDnBvt8LdgK2gKeOcMYqEfAYRkgXmF+zSFAlZ4XSvuAZ5Z9b2h
9FJFXfj30cuXZJrqrcFNWAErQBvQoQZ38HDvIbEpv45foE1elTVJNPrMBZK4DGHTot65g9sijr+F
gdqr2wV5XkIDIjW7o85ZwdFTRWkRsYGaNZ8lQmrKJFIQRidLm7fcI01+kw5AfTzTxpqQDKlkGtTR
De7w+KuJ4zHd7h1oodAiVrzEsrbrQzdkwLH+82Zro7ULIfeT3EHheV0cYj6y7xZPg3WARtolPJqc
7jD+HOA6GsXSVSui9oUXs4AdTRu5XfRXMg57SKBj7XJR5fJ+K7X2biBA473kPwmxwXS17hUeR7UA
ZpHy1eA5QQnRycYk+Tmy2d3IxVysCqx0r+k80wfNtZuG2yCZZOuong24BW+8VwXQn3WW2To24yct
bmBW9u9FYh9HFNKnid35/O9Fm8Tk0c9x6hKiwGot73HQ1lzPZzWSLVLLrd5Z/osCNuSPblqBDxDz
PF6jJk4ilMq1cowM6OttGd+cE/YSNv+rSTu2mSsFCZOtmjXNxzqmCt6TzVEYSrUcNR1hPDSY2imx
7cyusjeFVDpyO28PyIysjXBZC5IN1I2XQaq94LkZ+H51DhTFcFx6Bv9Q9pQb5WIkbwkXmc8Ugr9g
fxrNPlsNRXO0kNNXCB58qBvfALP8k9O+b/QXcxsYY6dmNSD/lmhGFEQs/6gbT1b42y32kPXhuJCq
ZBqypnG09tcH3aha6Ub6RvDUbPBkPL2ZU4/VmsLaTAHv3Pvp4swECPYmBD2Z3eGe56hGy75kogbZ
7nvvptV8eMKpmxUGVLl4hgZGCaCNDFJH6srSvExU7BtLs7qnWgwdi4sSpaWE57rfkf04qXC3weQh
gCkHDsIPmyFPrF+BVmyMG32oSf7d9Uu+iDiaBCFSGu0fcMTvtQuUAwecv8Lh4y5C9IFc+PzTrSUu
pNhlzKGltcBDyiLHc83HNBaL0PM/ksmlBaN5bEF9hj1R8PnKyXuW0tNCOFrVhF23QCAFkJ6UoKqH
Rtos/b84Jizwl2p4+VgNR/rpGgNLQx5ykkfHWPPF0WxI2qkCuo5TnHO9/4D6lBvOH0RkJ7mLLlWo
TIwlbZCwJp2EV3wmdTZq/I7yT/7sQI6uFOj5iR9D9rlpOkEzP3B0bBT+2M7aZxtkG6RzHmVoxPsQ
4ROp9eYIcVW1KCVbGPnAViQySvpZr0JUt/QNjEXwkIUzhUoe6jJNmSybc3JRA/b+aMtHzynmHpQe
L933U0klDHzjwUoWfuq7YO5Z1tGsHqHOOkExP7ESrjoxTzDDv+0HnfNB2HiqSpiKwVgJ1CWg7cy0
VGouXi4wPiMEuoIHnS4IALeJrx9he84fRiL0gL1lDk0bZdBHhS05lkvP8p9C2TiABZlr4X3uy1B5
tuNTiQEuFk/sXDVWId8qkGF7pxZg2lnhuYx9qgInO5rv8iW8diW6kPe0UDzQP2Tf4l2WWSmDdHbY
RTfY46az8VM4sb51biTu0XuUNwJCMAETheWoJoSNioXxzq4q5yIsqSdB3UaebFde6TMFHN1e1GGI
AGDkTai52Nc4UMHir0lpkpXGihB9Qo0ia6Zwf85GQ+uEREynjgF/IDcf3kEjfAA5VF8p1fDbIUR+
PErn3wJ4sa6/f78g83znvx2lTFfN6qBesCEq+EYsv8muxrOFqfI6W+ATsmKU6pEv5k+yni3eF3W9
uUhGB072wEsgBfl/DkoRIFet806Dbd15KnxdOeidwunQgoWMl6HFwvGxNnOOWFzzT/mIkwFYOEY0
tW0psColAySr6U/yjY81XMtKx8jXEa8XzomkwgQFtoUin/LUML3hDj1lM3No5c8BBv9KTVVJ/Bcd
VdSnLDYENB/+xjL/Y8byLdltem1R5+OoeHE7MYOS9aUbY2faE8QD/h8hJV3q9hnwuFIoI/zifGX4
fZDNho//FuHHfq5qyRfO2HEroFwUgw94K1EKPz5taVqklequgUBh9iScm79UhIBixdUxkCJ8TZ6B
jOXVIQ8UgEDR9WabxjaODuO/hhts5t/NXdHyVCWFKg3+O37j2ci5+D5LXfc4liQwzcHWzxE3uaku
yxuVCeyQiZ34hr94yTu4l709RpEd2ByUUl7CP0D0YCG83jHiq5Uc+X88IYpWOvp3FMjMAVhFB4w3
U3RvsWkgSdk5O9RhmJMSbkpF1GL50oj9X4GFnk9dAzJRt8Wba6MvxBSMI/b9++vZzRv0ms4UQaK4
q4xEqnwTaQyUdB1TGg1y8p44EK19c7tZfq856UDhRnxaMzl6e+omuWvKELGtRUftGl7Zv4y90AF1
DUHNjpRC20Qj964XBBVyU67fSD4ucFZck/Jy2ultH/o7/0IJZ7pHCKt0s2x1h9c8Qsh7bIn8Z23o
XWYlgJIj+XLZWU4MmRiwmalUPv0rLUDUTP5ti31MnPk2poM785pYEqXBQCOZWuuKwh4T7mV6XxRg
vmlNTLAy0ITtO3bXd1g1duA9WDAPDzq1ODrAN311idhOYYjfu/o1Xi1u9bpaOlWCogbU9/AH7Gwv
Y+ws+WHVYWd1pOqryhQLapBXsmU/rtdewnKf0oGBp+udJLlQemaacKpjU2TQ+ExH0t+se6In0KQR
jsyUfpt2QPz099eRGxw55jjHptOPfcU1PB+eEdOmYZ8sE8hqCs4ORMn/Sj8pCGBwYGsm0zQS1byU
lTr/lvxe3nETEcaiBHxKEJhDpUrQIePXGyad/HBRSs9mmaCuRijkP/4ewBzrpcMdSLkIER3OO0l0
m7tO1nKqUDaWM1eeQGV8MKnKAvnZ/vNJqKR629W1VIdytleVVjn0hix8DXlW2PFQGH7Eamu9TH9o
G8TmJObcnO71w0tUraN6rVV0eZoBm832b7wKMzwP6HsIP51Y61iief6+9EyphRQGQCGqglLiQj1G
4EPO9OarwY7Pk0xUe077X4MnQ+MUpyhjIghQZ/eaGXwfF0GP4g7+4EfXKNZRmR5eENvFTg2ysthT
HmfxUjOg0uvPBdPZPlzlB4QQvcgYM1l9ylHcKraZl4XXj/SNSI8qZmajffTvPuIb2DEFVv5Vepl7
LTbqw3XtJb4xExu6dJxAgyzQEHAIlBMzBvoPkOy3pl/SdewlXiZavJhmPaQdUx1VoCiaC+AGgx4b
vcy2WxTsr5/Wwc0q9dRukRwYVOy2/xKyRMFW+o5S0MbSDONmN7csOp9zJLzHAOuMElGChsC4YIqa
Obg+VYq69ebWxNoNcNG9qsFp2E7uaHcNtaHH480u0yBaygQIbMqJ+QIgs3kQDxgeJW+Fu2ysUWJI
pN1qfg1G+8ED4tBoS1N3SyxrWDNruvMJ5GyhGh5aEIRnYRMvvN6JfmR4VGVr9gjG/t011TdMtzr6
gvyvgXbB5mSVgUuBEk0mj5gYkXlyJrPCEwuEYjcyQVyjs+XfNz7mZIFqZfdfZiJ0OWBsXGG6nFL+
84beMgJY8iQplYATYeujSUub9P1U++vu6P8L++jfUyLzXRwAN4o4xBbHYNuLisHjmf+zQLg3k3Kw
yiTSmw6fOXQkiwZAAtEXLwmXvuIqc1YFhR2Y3HJec/5e7GZF+FRG+plZ6bf52WY/SwQ+Asg9vvL6
lxiTOdNMcIMpFAkUMroesB+Q+hdmahOg6xl8itBwMWykEweg82YItWZuvQkV6Lo+edjp3LkaDRio
I/Rt7rNKsqJhE7/d8DhFvHQ1OZWz7dOYNJJ8izJif3aLZdYVDFZ1/jdLzQjqJPZsDyeCIJvc6o8H
FnlVhCRnCSnHbsSxgSNvNVL9jVM/SOiI9np2zRsc77AZ0ukAKRtayqfhjhX801OxmatDrtSkiK9I
LBXZ0b0/lwZJAr6smCJ/qimJ0ucDHTg/3p/JR8HCIo6H2RBKJ059HjgxfByuNcacIsgMaOASOODq
YQUOZqtc4DUgIDJClTQsaSAGI82uoAeb8UDuuDPuj5j/iNXqCpu63MAJ463taEfjIL2gsn+LpOQx
rdeTO1lU9S6Zg+R4SgSXFYZ727r5ME0MnrprCeaNfF9SyKZihg92DaBcRuoLR/JMR3I/mb/0mWjs
WGba3TUcwU2OMhijIc5wMLp8hvoPGmawCgf8WyMaF62bo3i5lpJ6hWsc0r9hVBaL1SrOVwQIheRw
xdmyZ8MrRnGzBVNJSei6Ygy31FdeQK9/Jjuw3GSK6ORtxPiF/1/YuynCT1IU7/K1dZeWSYg2PydP
itOOnxRonl1LLXvOLv1cApozmWhP7qziHctAHeKVyq8FPml+JaKUMqQtnTpxccKhg4m0YWtkjHL3
yYrYGJ1VYeCMN5RwYsZjYm1z7eMvio4Y92vNS27i69S01fQBJDxAePcavosX005waknm37++tExi
aDtC3E0oTycx5LnYywJkQJxfn0EjryiwVzXg6UUFD7sTjRpOFn/Tt1LKFd3QfO5WXZYnc4dQE3op
jsXCnAjvmskvPIVvAXXHha7xe5c39Tq9dprQGYd3z6b9wTfdKqc4tL0hmXTDq7S1V2gDI3cb9/j+
yfbeIXxMSGs6PkqkGPkfRNJW/hAcd8Izzs5XbxIsxeWLXPs1JIbmT6MNasShT4lBYNQCJUwvoJ3T
xsZtP8su1/doo7PBL/LwVMnJKREY2TL4GmwbfpV8ze94NrGX+h6iDryXihQQ0NhKoQl/wCtQaf1G
bWpq/LJX72Zu29A+vEpnUlD+P+u+0vmhsILwChjX2WeP8HKXi3AjQNBpR2s6wspAvgAbvG2byb4F
h53ufGtNytn3mGbjM6iSCZhJ044FRXX2430JQulUdIevDO1q+eiBBk6vrPjh/I+4+CAT2C/qWuuv
Um8EOuHmVhBNbv/VTXbYNtVahsE70/IvT0XFkgerPDYCRSbdsZ5YBEr03dfEKdV3Qo3WK2ZqvmlD
C5ZufOlDlLlZARHoQBIkStHztqjSupGBFMo7lvXk+s9Pvp1CR/TuSsU3apwbhWzrRzxbEECJyGli
aRj4mZpEdV4HHNWFUo+tUBZyVSZLphsP6HlKsB1NRuWSNPuaUe3URNRf3Q0jxP8BepyP5tqhGvXy
Czuz3Ezxgh0n8MKpMRYJbG2I/YYEuiHobFCty3YJdzejhwibe10nVESlZDNguauVDCK6r+Hjwfzx
H5PSbfYnuJ8gnv4ylRerJyM/UuK1wJzsoFdl20bzI3Dd+UfrSwlzckcE03vkKPRW6jdjuW9pR7Ns
4MKUDoXX0s68BXN7xW2WyXt3pTRnLbk7POacR95/wwNIOvq8+yzJ+sQuWShRMVu58gLKoFmhiPrk
+4uZMHd9DL7Ym8zzI9ponVX+WpbOWvHJro54hxh+eyk+DvK24Gad9HqBkOEU6Nr910uaIpeIIdvl
kvnzL635NIV/avj+SkpKrTyPdezN4jze940tUDeR04tsccakTuacB5CwnhqTBoNbvvb/htHY8PSl
MLAXhMrCTPSdbXsHy8F/q1iAKLIOYm44+z8aeHxB/8neCyJjVohTue4PTAuP1wvE/tySn46mCknn
L1G1mT6qcLgMPD9zK6pZGuU2SPFwIenH3tXPPSxUfR4eAurQtLxKLFDHo7lxNtWwS2HuFPycNa4s
AScsulbryK2IuDbmj4XR5wihVS4pqJYdnhkXAs11gYOUigJO+gzlj1ensMkLHh6Llb/cszAvSsA6
Rx55qI769d21sz411bK3WvDO4UdtkhqdaFN84/pa7pntMhnFewGqrZXiG1TahxV0qrJJnKPXDr53
wmrFqxoSaVfaPKPeRetTV5r9qv8GoX+9Q1deIPWorO7xSvlNHxW3OADlNQJIYwVAV8vbxl4rzfIS
ll7tHNDu8Kwwi6I6PEvYMjif+XGd3ayJIiZSYbj4pJ/CIwyDz9G1ANp9fRDJFo2RlOYNfH/6OPvO
euLL5k2JV3cVbNMVYdV8JQEGsmdMnMqoCLO0eMNW66huTFviexpdgt1mlyuW1JqnoMOZuWu7XCQ8
avVRT1vKKlNDiltqKZCj4/NLAC8CvzniyPNjGyt7eikk1voBebLO64blRkPZtObrqdA0Wnmwcr2x
0LvANWTHtbdDixmmS3YaN61s3A1uxR0yhSEM1gZIEIKPgaxaKbaW3OIzfSX2Ftk6b1MdiuhxjbZH
tLXXGrC2nKifdljK3SmwjGFWymAFwGungtQCBhQHuG7bQuvD0ec676235kZUcVAfYch5XtMh65YT
TS9fRFmGI5NCLIaNRPDj9yepO4g2TzNaeywH99E65o1EID//4bblz+BkGQFSMvYHh5jkz36BQss1
dPJBp8sLuMQ8Sh5P7LRqbzwH7JmaNkniSXmMhptNye8kE/FrfSZhLGmaYk8TzpWzIoEBbLGx2VHS
OVTyVPPFuY7yhnQREGQ7zftnx74mnufTgLslfGwfyj0lCFq7tzzgOpBqLrQXxM1Xlvz2Y/JXw85t
Z0XUc4LQW+h7tVS5cYO2DO+NCszXwtNB4fUjs5Ddt+TDYoz7nga9tHCp1UrNK96c8mHqB4U0BMHK
xq57tUjvdWqqW437U64n9813Xmxb4ltWhXZ+RYQrl6sfsdDwTHolTFFZRnJqcekMo6+rGzqqWbEB
m2OQ1pkY89UOuaV9QKUifleR4nv9GCJ+T5XkBhaFNGu0efUkcShD4JE/smwiye1eK0iCKIQWojui
Ibl/TxJF6nuhnxAnCAb7NaAUwQw3XX8kLOa8tuQbj+oTjtNRMZB+m5mpVinfJC9uE5bX991gLZOu
aXnth7/uj5IkB+ant1+uCwco+fPK9XP06Vq7FO2u7CLd/cDfJh+G9hPuP8Et/oK8X1m/WNaE88M4
sbAbGb0Wa3J/H88A7/o2aXYbqx6Z5w1+DeIMzb9827hPUAZNfaPtH4vCJISt97gFXm9in8b889iX
K70GWN6XcilChJUCSZkCZ4WM17fqXdxen5qhfRoBdCX1v4ORerwNSdE6BR1uA/wzx/RwqxrScJ+u
JuvKu/P8KrYakB5gcrWM7fuCXMHJBtJKvVWVkPiqYA5ikAIuI6fcMKdsQ+yAZrL6rgiCT8xhaLo6
1OLeBal/haRZ0YwanO29+KiNvQaDSgF9U6o4V4fwddAeu51VNEFPHXX8F1vw5+dinAXuQeoAx9M8
XZmObRunx9NHq45eZgRMK6i04YWjE8Z4F7eRyxfbflrBXQoZ2Orgjm5VRh0J6HXJjeWa3cHirbBq
E4VFWYJ/dZ9PwAsJZvHwpHwhzHS6bI3/q7/zJOacTlXwUxzhfzELrW5KKf0rWcKwyghKDyZcy1zL
0GnwSRjM3cO8+3W8Di3H5gNJV217MhBAQBFphQTh9eO31O/2NYJVny0usPIwNfjZgYDSrCohI7Yn
s1bNOkbu7OJGQ3cWk9OPMXCuB7JUrcoVnZBHBIeKEIhqc9/UZSEMZqqRCgLV3Xk5Me6EnY/KVnCA
r8ttWbu+w1U1JunhLwfIcUKLllbqbp+wdE6xStRMQOSHwHPbg8k6RCKeblcaUXVMg+FGx+v6cnTn
QG38DmKmTqiDE7+m4pZHnN85JcfYidWthTIJTZBhnsUvgLmjKmOJEvcLeq0ygORk8B3wvCz7mMXZ
3aN7JTnX96RUk5yDMUvZRHjrMPena9lVMt42tskYcrQo7otGOiOe1jcMkB5XnFxTy0vDXFRDzS/b
0KKC9Bi9cdMX+wrN1/bIMH8GTZ9eXnDvQDKOwGNog4iM93E+Pf24GxIeoTQPJ73s4ELPEllSBPKF
3PZ2KYfMFto7KfMmCzAl0m0QcgFCmk+kjASYYJpcxZXZ715SL1QxXyV70W6y5rZLhqYpaMhPUgwc
LvhKHQBYFzBX/Xni0Gyy6lg8JIsQW3mJlxrDgT0G9pV+vI431CA54kkyhQBoTli+hgzTHNkGWnY8
oxun31MuLZir2Da607cLEu3wXGAFEXDvMR+UIcdzeYfqoSSPcvUCTmkHjiqSjWrylEdRjW/Pe5lh
vGUBt5kx6TZIK6ZxgJSk8SOwSAe1YvE3JPyqUsRkfLd2YQtnhsWkEGwcKrBzUiPdCE48CNr8CbFC
R4cmwJhd5thog6RmbLF5NAV+hAhBdg5FnuznPAnlC1LZ0nwlZVqqNmaH5KLWGhrRYWLoUuy3Qbw2
axHPlMO3ORLrIbFB2j1FkB3MiAe/IANQDYZHHxnEih0Pfh18hHpLHXQmy+h6DwSc13Z9n2n2Rwy1
K6Brv4dnPmJ3gFE5EliqcCMFK6UQlqr0+PQCCLYUq1+JpGlWzWK0GnI5K1hHn2hxNIWf3Z3nPKJ3
qDYJLOVV9xobBw6z2TRgpIUZX2TqdklKlRWG77d5L5FK27oju7iDqG/yqCpYIu4XE78sSyqu8q5u
uZ4G0j6Dj8jLEb0iQcNNlAvwijFfs4McWygcMDEJ4egG+qKqLoAgP/1+cCtjuQHAIfbKHck5i5mz
urFtzXzl1Y0YUvhF3A2R3FDrZGog1LlnuPk1DLKwVT+T9ua2U3S/KmPDYYI2GA/jMdCXJdYkgL8c
E2FWRJEqcIu/VcnvuH9n+8iz6tFFD9teIfj7cqG/aaLvB9qDaRdM/vHyTu1OKfUhb3gr1oVBNCk9
/0zXDKIuTqMuhKW7xAyyqfKuGCngy3EhWGMr7qrDHmUhzbOASqSbyVT0Rb++3UnVFQuj7znRxyJ2
fOgFAH102saLjFYs51mNBR+l+UmFjDNVlkb6XbqjujL1N69Ylcn0qM7fBsCe0fSM30nPvlCvB27v
wC+swRYASYSzVh4hnL/W0+WVhJtwWjsh0zoBfEGu68vnSry5yR2Y9Mg5033pmnbKU6yKCeKfHHtz
ffGbW52NqOgFERS38Bc3mYEGBuwphM+0OCZ3ciP2CP8uBYdC0ULVmAQzVhvNBmtycwkEegCv5sdc
OMpjYp6aiNj/umfqbs+eWNonIeMguRR/n+fXeC4UHBexqZOe4n2ufElNuQpPv5cpfDcEy6r/eqty
WXuZTHkHS3rlHTzaWu0IrBOzydkT975NYLdjrYhoCeu44dSiUUNap7T1RJDc6Rx9SRCaZrV7x40h
VxAgI1dfE/2eeDozSmRkF+ukntt+xAVLycX520a9FO+UvFezlyCaH9PQDIGh1IxdqGYWvuc7zCmt
lhAlrWO+9USw5Sx1ctEAHgDCyvCxDL2sMGV67dEXbJKqpl3OKe1Mqh8ZqDN73+Su+6yxx/5ACDnj
1khyToVovWdO7UHDd0Iswn5s2uZO9x3EhhMoh6f48yr36xjhsNM2/0R5iNQ3WiPhbe286G/2PsAx
f2GE8cj4y3TTK1uNmGGdsF3W3aKG7ax2ILaSIWk/9gEURT3V4eQTsVLCWfbiE/qrR24WR8Nn0PzX
ud06tFdQ/jgKHbsSQlJELkZ1XjLR/YEL+h1AfCCo9+YI5Wjbxb10JVYC6PptvsH+wEbsxsvqyaEX
ATmSC6ZxREfdkiCI4hP2B3Ru4E4AzTUumvqrN//DnkdVDka5jt9ymWPgp4X+9T/DsSaRJRmxDYnR
CFklp2VYgThAaBQcIbrtPwurr1v5ylFtTys75AnHCxxe16PnHXyju6C7IzTEST9Fki/P86+AVi8i
cXbAQUjBwJJOPC0OI1Jxpx2xkfYGo6BNb/bDCOROcLdfkaGLSv7yyAX8HydULypJf9VB51OmWcBR
xbO4DWdvsiCBsVnuEQg+TjwXUpoEfNWC90dQXE8sbu8geadaN1u0amib2OXgRTW1XjSuAhputakj
dCIALuLZX0eJteUqslw1NoQCrtBW8Kv+1trTOoJzzTwLPiKUtmtgoSuT8cofuC536MkuVFnMmtsV
clG/lJYu4r3HCR7E6M5L6bDHW3M5rcBdL9ntgqbUnQkMUQYLRq2S2Ov7EG8PQSzxFoEL+YJ5HnCW
dyU8rduYgpotBPWK/V+WXygbP313mZnmoHt2hfBrMHomuYYjH+jJgeqXHhfFenvVlbSyFI26eQUM
B4BoF99sIfSMIiUZdk1Tu6v86suW/LU4AqquTe/G1gDAz9AchOM4nKnTpZFXDKByuU+hKgtyShAw
GhUwkAgWAOrHTlsGB4hod+/71tJvbS+D0bsajpr9BgmTnkSsnwIHY/OEuzod0WfRsHSELmaX5qTQ
sxuSsi160OibBQCjYTGBex2NlSbzaVKyvdXKAog7jmehTNc782ZJ3raJUwgnoXBci1i5VUCdp8Y9
4tJs/+g5PqD1HYFz5dYuUZlnpBlmNqv8MvpJhUhsTcvFjUJagfqRFMiseZMHWjc7uOBrR24USTvT
6l1MLLBGQRn4yCHvMrHVSJ57p6KZyxsvoJrHXlzLkxaJEFk/fllNlj7x6QigMoWuOuVS+xEPfJSh
4S+S3ULAnjkWuZc69RqBAvIpDMjMc4snHgu05b2bwhWXyQyewoQAwB2ZN2ZMzeaMHmsZv691AXG1
dt5kCzovQdu+70xxU/+lliUTPOM2gXdaR33GiDUMyhjoZoic/6byn64Fter0sFw3jd9Bz9FkcatJ
A9+fHgzWIF3QBDB0l1wiA6htFFXqHkYE4vem3Mfu9agX6XGDiM5trg81u2HvEsQ3tDlECpy4V/Jx
ADjs3pY2muYLmfaSAyhgxwIEi6VMjrR2xe30iKJkCf1qqSEQP22TjW8+d5Cfz77sfe97H6Un7AA1
J9a1FsVKy8BuMDX0tOGQG/6b4MpRbs1NZSUBtScrHSsthXPmDat+rPiJ1e6L7WShGen8+eosZg5+
L9oQd4q4rWvTYqDPE6PMTn730vmNqo1XVcAHEQpv0IMC5JHl+GYpbgEg1oK6E6n9dieHVZqk3kYK
Jc+50TvOOKjTZwj4//wv2yM3rTbxXYgfEg1kQCzU/iktqmQhYy4POEnnsGRxkVJJrFQE0IFgrD57
eRs/QsJi8nT68LcC0NV1QFOcF62TbFhPigoFhyW5wsP36RagUqTnxiNV2fZ36OmXGymEA4iaizsb
rp+jYiaO6EpDfTdpEkL3OeSOfbuDE1UqcEh8VNWkHZiCuDP6h/KAU7k+Nr6oVehjd9R6dvrkTlVf
Johv5b1fsBTLWi0IjEqiz658F9TEEbB1J0vkC4P32vfawcSnggFvW/XNJ2b928rSORISX8cnAjj/
/vGIKmehhL2wF1aBGmDj7AslVVjESlMZ6y0O7KQuWALoa96T6WyBqZiz6FkoI3dX90B8MVBySFQA
CCy6DOg5stlrO2kfMEMGIzsrM0DpAl0R7YRSulMuy5csbOYWLW+4rgLSL8Mk6pTNnf/IlI5Y5V/D
rcCRmsKtsnQP2apjGBzi1CXnfit0YKY8CIVrHTRoXPSISClpFth4Uk1OUXPZ+xJXsJTVfNGawSv+
qFACx0ZIpPF64bH62nvAxGW8AUw/oogawX4Ym3D/Qg6KDnE+C+cZIlfFU+uyaVyMh9iYSuxgEIqS
mi2YQDiwAXylYf9Hg5ju1fkj5xVpuD4e8gJkwPlmLGh7d4VPlpnCa51AD7pdO7mtusObgoYYdxal
I1bRPzhgVuP562Jv8aE86Cw93p00kd/Q8cJOliDDPUhDxxCWLbaAy2zi/Gx7BpmT9S3nUikS6j2I
SXazQ+AUNvkIF7W+T9wRcMQqz+HD9e7MpKTnjWeZ26KV2FtkFmp73NmVSfOK4xpP+1AQG+B2uXMN
9/QemLSnIM/V7oHULBx8WN8MD1KKbGVTrz7r/TsTrY1xifkwYT0MJhZQQkXlvghVZlQbZZjvNp2V
vMPCArM+y6Gwon1xM6p5VS1l3wDd0u3PsVQjcPv03kBbQ4JkWgsS8ZEPCZSrkIbCVM3leodIJjbi
lsmcpBvFJYRI3SWVo2WTFLnsb5nx13hHsHHf9gFtYIKNYULNnVtMU3SDe6CNGALGPXECeZUbLwt5
0NESVe/Su14g/3XA9bB5EOL+AYKDOhQD7bT5fqllBjcPR7SBGup6ZvV5E1lr2FamfrwJOKTIr+7j
6NA0+qA5z7UKa/YRs20c0ZKbz9DfImeKBgee+apnkPdMnEX8X3N/Ss6aUVKN9z9LjL+dG2VCfABv
P1XkZIHz9wmuS7FELqzJ4QCmlhB+W9V/u3Yh9cE563Je5vVopcMVqPPqljHazTeuZP+mjjQl5/0J
LMSk6+rKLIWY9LVJ5uPnlmFbfum2Hb41CkPN669Q95TAzZskLk1SGOQKWRD0wCDxWNfqvlRT8U7J
cNvnxCzHYKbPUcAL595XWMPQy+f53CRBgdkA8rl6pBPG0jg4bJl40KsW+SA24JNcgfPbySsnBwlD
v8l2IykqI9oo6lrwt4fvLg7tTQIbVTHUKupkkIoPPHVLnlAksKapU2BF478kzknQYZ2eQ/gaNcyg
qhEMsOVxB9VLj8d+c7v7kGPFkeVZCJmdsmlxFFL7oazLT9i+nLpunzJ33AklHz5NOq+XiH1MXC2X
k6wF4A6mFHIHgcnmKClTuCaueOhafGjDfSLarj/0RAlXpSv4Q1myYlCdI0Og7rLe76XejR4DiKoK
yAfmIDnnmvwWhSHW0qfouYWyeamRkm0YjibsqszLDGoEHRTheh7HVQvwieMcYQNX9uLCdqLIWWjj
3XnNeyoGr6gcj6kjVGaO3X/VYVXV5oDJhFEfgTxeNy3AXazdgmNp/yDkRTN8NDPneds1KdQ0KNnb
CrxlBlHMRja1z+OpEO/SceTQTxcI7BuL5YqziVpAlzYPdrICezZVVYOQrAMVvtv8BT3Y9mHUIN5g
vNoHkOvHaVGFZqiPK9uGTGkywYh/HcpAL3pOCUUflpdFPNWRPQzJw6QjxJ6/1hSlRdlBVkM2ce4v
uOmwsjW3ocGA9IFAnr1iO0fFJcuhrkwV0dnQdUXVYXqZbLPfsVI/1sJ2eQ5ve6Nr42TsTqaHJkVb
uh8LsyuP5aWLawsaIK9ahkqklNobTbbuEZXVKNdc5vnbJ5Iw6070lQTOV1E6l8teM6/Tuq2d13HE
QGMsLQrEQC4NvAY28aX20CS0qe0UmVz62Ztnsb8Ki5AMa/5WBvGScF8q/9NJn2AUsDDrKPm5rLo6
0kwEAjjE16Q4e+O9TRv2WqWBA07F/PZTKYpdd9X9fl24n0VSZkSHkbhU/fYo92o9JSgAc4LAjaC8
iWbsP6h2dbeuScI+5jDGgOBqPvtGvC0VHbUNY0AprNMrEuQ36qD0dTytEUitSLoKmPTWQofkEl81
shfDnIHRJWUaKSEu66gNwdpC703jG5Cfg0eWj8NzNw0WuREOIj3C083WsOxpkOXIzDgV2e8cPZOG
M69YXfOZn2tjQgHtIQE4CUUSX+CUtmJ02uPuzPN7D1WPnHBaUZCJJh9wcC/a5qTqADR6wbV5gpIn
gFEA24LFS35M1VdirM/7Iht9Ble1RYRny7g7MaxZzZZly+8TMHdv78RC4z8I8IjxUY/DvTJi6OjA
jWUuwlyy6H/DLydvXmzmgcAYoSEreBDLs30y/5Dc2MCw6D+gPWPvOMreE8LWXoXjPpOA/jJLSB1y
orvcG+OnNIRDRgMxf1dKc5gpVFq+ejvBGibI43g44HDZC5nw94q2297jhjobjXTDsxeQq3NpduUF
oMz/d1BzPRmhUCEMBHPPMIx4KBCE78JXLEYfsOkZDCQOitLpHCVwEgdlZ8TaKNtUtxtq6heWhHSv
lB4ShBKb2gg+ukf0XZSsnjdsdvO1Iqfl0XK7FCp9S68L3QpRoGVXrbO/GpK8L0dRZg5lNzG9d+lr
UK2ONGhiHmKpL12EhG1FFTBD6Vk5bFA6ddhmyYamIBEsxBTgnaPyAny5sEihbvyRWHTJzIECuJ3B
GjtZMoVebbBOmz3dGeKiNWP26KhjfWvQtZc2S3QS6w5dP4FID0orMpvDpRBGfqEu6qYMao+c1jFa
Y1NhA6dDvHE3qh62XL5eSzBr9L+gZR5MoMn/M1mNukbV0PRZn1SsCGWGiOz/GJScXTkmolugmI7w
2J9NIXhprPjxc5n7e9DuNxNkiFGDpRsHhji/9CAdp0XDBFfR6shFjQQWedtZ4hE72mPeSzx+cCct
01hxsZWK0YPTlyjtw2/DszMrSpKFWykXZpMoO9jJExPPYEBA1DJdqytO5lh1L+bviZOpXfXMWnVQ
RU1hcnPgmg4wa2QMjyjdzd+/fs9idbZZE426ufRDe56FCN0yXLy2bafogMYgwhhjW3EGAEcLjcdW
bGo1U8Y7TkRByRoT73q2l+l/MvSGlKVIB0WERS0OK3SjgLPFCh92LQk+3D44/jw5rFXGGJWPLMP+
CeGPj37KsC4MugUPgD460pV5Oh+PrGo3pn4ya93ds0OEcwcPRBeSlGBUXDmOaJfsb6SrjbY5Iymk
cKHQAcziLbXBLrji+xs4qZi/IfRdvzHPY0YzfFziWEdXwngQ4+VLWeZ02FRTeEorMOINrOXMrFR6
QuGTOvNdBB8MZnZHyNqcVK8LBpNPmunT8kb36AIRyUD+lRJoMjL16O0R4hyQDyk+7kxE0XrxhYpU
v2k8I/TYYry7fsFk3JGNoDBevnfQ2pGVBX9XpYThZ6Fc9m/ADHKNmnHhzMC94cIVYda44QSPnkNA
yBU3L700F8IETGjVv0vkqFJ3TwU7/bFHtD6b7cTDZypLVBfLr49vW9WgRXGFz8dCfxtfyQcpksfA
+aNq/2jiodcFjccmOjru8a2Bd1mFs7u6fmV5zE7868Tt/0FbXCKZxjfE/olZJiAt1t7iANeaA0nS
GQjPktOJc2gDmbG4xfpfGOSE8o3WPwwZpIEt8HsaSA12UnIsRMAbQcrZX9X1P1fn2Fk5TwDbfoGC
Y597EuoVl0/68z5UpsnaTHb/LlF6LQVA/EWQ8d9K2GKPEsY83nNmQrL1GeZINtL0I7MhRXSwxEMW
SZpaDLK6kQ/JA7YmVtofIpd5CA1y34t2fojziaach+N8kJf6YWPRxAlCGSHKzKQQUl3gOH9edcaB
xgsSp8R2Xh117+MQhykrHBSb6y+4OubCrV6h8xPHUpB/MCD2XsaC8w2ROry3sg9XDD7+Rn6RWTrL
3S3YIx0haJrefiL8//Ra1gMIx4JcDwC8YUk+bnSOOL6OGMzNwgQovIGnLlTzS78cY0Sb1Pp7TIai
262kfdWFYwvz/XwX59w4h01BCXUcoc7lKi/OIyf7k2btfll4EjonSK3bQislDcg6XEnxTLY8MjeP
v3/Kl+WOST/jEIiHHpFoyjN0xQT/X6vFbtEwwLQsln6l+Q9SFkBAX4VNAHJUnhK9Pqjg9MyoxSot
dcOaMz3Uiykzq2j8YQD1UMS36UYUORhyRT0YBo13dZ/0ArNvph8zx9Q73wHCxGBD7kCIH/1L3wYI
OQr94OSCJR60mp34fdPLcL0ub3/LtdpyVIic134ZwfHWeN15hDuEieShoTdtDbnpOK0SlG1hlHND
/X2dcKvZ1I/2w1WYBpKmRVNPzZ39kCt0AWn8eUb7BtvEDe3MB2r8O9ifbkL1pJ5E3zZl1gnnieBh
1e/FwU7rRPy7iYFNkDwblsjHxoBNc9/hlujIkQ8+Kue0j5T51lWdzCpBgeDM3ZRHHLjIftj3ykKb
x93RrGbuweoDelCtBdMCG37zu5ve64KKqLACGf2EWb2iyjQm+VFeSpIYosvM/2XjrI9+n/khRnF5
JvYB+Brd6tbPORmm9v4Gv2empOevl1iTARPFxkf60hcPI2Sq38K+raGWNTHdyw9VHolqxvGk7OAf
UjiFf/ObCOIa8P3k4ehOWJwkERECA6y9fFebBV8UatfBOnY7wIjnp9Kleam0H66x7vScZNTiJ/sn
AEaLozlj2oMxNXoHK3BsxF/i+PatZYeA7xcjIjHo4ipg7oRPYl4CVmdonpx39MjzXA/LwzGYmue1
eWbq86RPFnY1HbUpyLNLVcdfuBJ8vlZOjTrvmki3Uocn7/Mk2frq/OzGmUokSppfOkqU2SapDPqk
YQ6ddkmR4DSiJKCTJsrjhKyNK7xtK2HUqbJiMu4tRXzVaM0bxmgeYqA8Yc8hOgZLl0rIDDVwBtBr
hTqL8nZUcAkrBiy2HsJ4F2q7n8oZsbepoHjKs9dW4ffg7FNboIHDVkdLOoEMI6KqYZY6MAmTNgob
QddwDAdtzvNLipbyBVHLYOyG1jacOhMXcbN5R2j8YZQ/KjcqeutcTbxZEv5wGzI/2GT4vkkQJBkw
UYbDF+HERybWRubD3yLUP/QgVC+GtyWxttnKMRV+jN8SFirJIxgeUs7MQJ0rRaKwOtEPAVx7YhlS
yj5IrmXGqy6F2dziHGQd60EU+BI1RLKqUymWZhsNVfo4YsvNyGgEL/MVSq/QjJtMiLZDp/skQ4G4
dZcRWohdQ+afvyV2xE+oMgI2TLLFmm1o8+Of/stgoMb/aLSldEKsjfOQ1rbP6O0qMiCCmiZp2nNo
VrTGT/P9CH9F4uWmUMT9ECKZW5G8nurd8MpKrP8+VoRs8KA6I9U7iYURGMmM5PdfNsEtw/X0X6yv
owAhvh+HZazR4QlTSeAA4mIY6iQFa3BtSyJ3AR3R7Z16r1e0pVbOpatX03Pvg6Wt5S2mo+UWZUv0
QwO1XoIF8NP/9vxB8LodIokoffjSK+CP5556rDufn92SJrBkjpyBuaQ2oePxkVliIDKzots2DXrt
2mXzR4wicjhJQeL7kA/UXWIIzAmeUvVToWPnnr1RNLFzQeWeO9eG/8BlEjHVL0DuDruyVZC8jUoi
4Fl28z/314Jn/uthuoeOxCtNRQHdEkFZrSbuviSdyvIITG9sOygQxowDNOK0vrkQGmwtfPz4gdYh
RmLNBp2CQ0pGwkkh5Nplj7nqqDGicvursbE5OWS7esPqtq6nFwHDZ27z2j1S0FJfU+VPvVv7GOcz
dVmyQjtEiu3lXr7XPySqosnxb/PrEj1kYtUwc91g4IYLZzvyHMm4N1Lw+hUF5WTHkS1iIiIw5E0n
UT6L+ToX64E76wvDQU/cDCm0XGO7vHIvsJMwBCGMCu96Uqkkrik2OjKXsw9Hv4Krnk7UYqBIyYJI
21FyAvBMMjG2Ft4kQUgyKOYWJ1FySGlfWwPv7ivymhIFyNPk+2IKZtQ/lV8+XwZW49dgsmu406fT
ew6K1heJasyeL0/wZCzQlR395SL7Dp8/Oj6tqLz5LUhiAA2KKP5fYvBOSmlc0kPz+4p7ypVicnEx
i/5tW/J7fCRhMP+u4USd1VAbQ0Zl2UIZyKQNtAUHwhosrEUGHXzd5DTHieGGbrov6kNAftans01/
d0nQZuSYFRlXJq+SiP8Vn0HYy+yvlqkFc3zQmaTnlUirXodG6xqI4yePbSGvbpnJoypq0SJRHY0W
bJV6+I0yvs+HqBOkAYdRJYXMT5W/sn/5uUrdJWImuRRjabqICGZwbbJOsT37+75kk6xLqQnJSOef
B0J1I/LiMdwj9qgu/WRLV2b4SGmWyNSV13LFFaxsF56NQJ7BQd/TuTwJZSfSVJMHgij9rFjUmJ/6
W4AWuvcBaOV0erVR0G/xJYJmWbYaQAPisrcSY+C1JY1MK9Fr9W/hmwaXNMu25vZf7B2TdcrERUPF
i1KG73xBxNMqsDQnvIZ3PTmjSbD/plhkU28fVAPxxPIKLAbWogd34CnokrueC1SHswr+rfuATKM9
0WtNCzPu5FtvCNzOF9vlK0I7osKOcXV1YCvmwXo1Nb5O16QtMVnLh/L0cExLWDCxcURAZafbdGDK
JdIWhSdilGBCocQ1GVK5v+ie4+FMoXb/24ZOM+XFjJWDtJxuiL81gcrbSEVU6kxQyd3Sziv16Nea
F60pam1zo0MJXJ+I9C5oz7hh9pKtu2QwbNsMadtnxh5HpvlwyRuRoTUK/UY4LUKrj3HHfZ2Wa7eZ
Q3LNgPnimj4HvbRuwL/VfFgdrHwRHzDcVlg1OJRlVVnR1jj10CIbZEzOkuB02cCQo3jTl3DHUo9o
OFvaMeF8uQKIbs3bHYDQ0QyJFIJj+jbw8XpTlkW74xQtqz8jsMa7iog0chIWLe8Qe5cDW5J9Iibz
cXB8/xYs+FDuAqC/CbN/LTvJx9/r+1XrmFxXRg3gaozKeaKNy0tfM24xvpzMcS893yhLmmisk35U
YZYQw+rgnlGacHU+DeodIOoodmWbJvLF6GHCqi6dTsDa8+SWV4nURVNKqIwLtOohKZHbAag6Ph40
4ZNseqb+c0+iliRbboS4n7XQ1/fkd6jpy4URZ32HKVC+nCmHJrqt+7F4mS49DqN6ZSrBP5mS1eou
clmVdbvqNssr6f3yekMgv3/ZLiD6YSwP+N8htoOboLIO4DWsTBvnPmUv92h8qTJbszm76gvQwuCk
fyS8FWrHlD03IJxjY+9B3wYuP3MtP9D6j4Z9+fN+1ug3b56NVekwwcUGMVPQ3Vc09XOIryNWiZDr
81BBJIGlHplExDri5AB5edZLR0Co9csO55dmZlj9skr4W0fOohQcqDiSRA68afJVCNC3EvW6lE7v
xbiuT+Rdm+8WsZqMMAAV0qUUv+kS8jABUs+fehuKwWVa6le5i0Fq7xlFpVL44LXLoV7k5HXEzr3g
wgKDjRUDYISIkz4nYuXpAEPAcIzFdiqn7vNSEnp44yvf/fPXPQFjyHTXJQnntnigftayTPf4wjW+
DoXlvxc3ZJkGOSeTIXdrHYSikKHZRPh9zKvc6pPI90XbwUZAZRO/HnjubjPrrJHjcgivxVmijz7G
qS4ChYfRKT1QKME1BGU24dWhRk3HC+KTwAm5KK4MBmYB4gQgLoO553b6zYPjGpuMvfUle460xXbG
fGCmKUOEXaGFKcRfPgrJMZaRfNdbM8ovx2LUDgQU9TitgtjtPa8kr+PYPtMryh+EM2k+n40n72Ao
a0DL9Anc0AAN+S4nMWY9mMErN6tw0Vta1FIFINkYfOewrbSEr5eeB8PKfyO6ckdnj9TLmcaSJGQ5
doIzUOMd+rVdd5FT5BL5/gUQqzPky1R+M1ITR+NzrpanHtLPl0HZpXWaez37VXWtD14oB/wSdEyX
zuEkmU0SpmvDOeetQ9xKYid3Ph/Y+WjgMBujW5qQWRYPQI419sKsZiOnflRwaagSXpnYM3XTZYV6
hL47jSU7EV3naRHgLb36t5TQKtHQu+Tz9keXC3HECX6/ewW84D3r6wwztuw+0toWoZPJlEdLLxzx
Y67M4ruY/dGTvDczYBX4ZRNBFY5llqUHeuW651SxPf7HFYeHohRvIqdkoJGY+9c+09/tEFJw5a2b
jEQcILBp2be1MrsM1bB1cxhVKGDVmyRsdXixgcZbcDtvjsjWO48uhN/Tn/ulco/nOrg8Disxwy7V
bNsh6OIiVWEA8dvuCjQIFi5ZWTD2CKNv6Jnqrx62inUjTTZJL2FSSiyJHYDQ7nXaLsS10zr0paVD
SOTiCctr+9rEo5umq4mE5hxJYkm3PDbbd20VcFfNeEzJ2euIGpCzOmItXbOih/ITD4bW0RKLuLrP
4/VxMV2AFDgANCht+lZS4PmruK/9FxP9PYG0bHT9B/e6AL35g+t67nhZpv429sthis5PYc3rJlY4
dZxjhDBQPFB6renPwOdT6YKrhzalwRVkK/pZE//2kY5N46an4HP8OraU4X00jO4Tw1TsHnoBuuQk
QxSns1jqyUB7ZCyzicaeJWfscJwn1zV1+H2UiT3ujUo7VY/0lufSKh4hHq8sSiRtuyHC5T1+oruE
CnUoi7/j3r/CURBLEJgzlDb205O7DjFxkcpdmTAuhnboXYMOuTXdU6XgNjz/8PlEY/nCIuKK3Vpb
2a2YDr+pKACXyZ+fZfJuZN0pQElLylt2fjNC1lvj+SXNuhMgmys0SZ/MqnnBg9bmpwMK6R3ZE8hY
ddr+L9AwOIozjU4TB0oiPgxXk39gJzsr1o7IyNQyBiv2zKVngpGyBEKWQO3mvAp78JCKPV9djd6W
Ay1iXmlaUFWtBORVJrOXi8Q9d5ohuWEYtAKKRyH7c+jF92D10Dpft5XMMG9oUooW7P7mqYb1uJHE
9wzJKzaoEhDwRQCjp7PS8EYrxjqU23iefneHzmgbUAOMFlyIAlbqinoIaETfMb6+TCFpaMT3Utea
MqBDetjsB4LZDk/dUBGAuB0OVMdiNLgDGxhMUEPb9uZh1kHEJ+r6URDo9kivoTrBzZRgh/wxyMj4
bZZ3zdlueDEJzrNadAQOalc1SGSN51TuHVYDzQKLl56M3tEarXIoxc97uFgnbH19m/tNRQBz9VHP
bJzS8b6nTSY/1A2LgjBVvkc11j77g5oSQIw2DQ1m4RZDQ1e1810Kr79u6XHb+iSTjwKS/JkCn4ul
IDV9Q7gHUafYEeGKASlCrEE96GfA0nf+8KlVNpX40dcqXd7eCBhfAkJl72YR/q5ZNQKemdy5Db10
KEEJQuSc4mNYUvNXkYtaogT9fVZo/ZMUw4nqi0nYiCy21BbS8MrtaQ3NY8Hwyfjpbp7Uj5zFa/4b
g2U+y6DkUcmm+YvbjxUaniOw0cA2HYMLyNbeO7tZjNlE6TbjMK6gcgrRAQd4M34q44551AQsgJdP
ECYC5knfuKY8+VBLAtRKdRgjpAzXEVy8Lbx/Td2oTO08gQZ/zD/k55WdAom4leeXEmy1SLnm2s/d
ZqfqPW9KUeI5qcl5keNvV/CECbP1l1gCIfzxLQfTcIhMoN1tFZTPpBfbO9WF7Jvl71EHwQJrN+KA
ubF7RNhw2QkaZvk9GJBXODZKb3DRITpaVsl84no1nXvBSaDpC3x2Qq84zau8pQa1hToL0blEoMQ3
2y+qQmQlV65+cX0PXWE0WWfeBzkccE4upnEL8l7vZZqiRsQfgteNopA5j7WFl1kBEb0M3UaI+PMn
2BlCVRQEuBE1XsPN5ey00rrER0ljeHgG1ISx3/x7AnRgTz0tJPohARrzFUYJ1AehUJLtG8MkVoYO
lTDn0Ny8AIxDnDnw2GQGCFW1b2fojj5Q2GVXbet3ApMmXcB49uHfgGSSr+DwylRpub5PjjYpuq+D
eF8bJ6IR8S5hVbH12PhJUKCJTBlCG8+Uv7DZvnHYt1069LYDkVimA45aKQrN/BKKzl1irUa6inBq
5KfUqiD2cyND5oFJXwzSZeMWbRi5PO0Z9QxcRYxFk20tzJMJK2P0ekPML8Yrst1xf0ff0EZu1V5A
gCK80wZ172E/YHAqEnU2ShSbHeWOi2329pTp4iDdPTmkFxUl3zD7h3pxzXL3yJerGIBRSRBOYGkd
4jiVLqR4A7+Ad0Ta+FG6WD6ESjghHv6mIa20R8M00By+gUK77OnZODzAnXdtwkE76R6NjJqzL9KC
eyeQAfme/lQDFJEK2g9D9G4K30VT67zlQwNOLPUBPp7gUKBdf2XxkGlwwZgTJImSBy7aOHa0AHVa
g3TU71X722TgP58Jt4+Tozl1HBu5TakqKB+a9kLxEI+09RWCAAughThd7ju3vnEeOmMLgeEOeAOs
OZPqJdluMX4f05Xl3Ms0THFIVttKKOrhwXf7YXXJNKCKUmDcyX1PjgGgpK7oPbmKBZP8LIg5o75c
N7NQ4Li97sA6xaeMfwkdQMon9uvm1TcdwtnbQNhvtPfHxgBaqvBMdBw6TX1BupGzaJFi2W4G31Th
vtsNekxFimiyDr3icWZ9nT81+1/Je+WY2P0mknegIKWsW4fWZtgYWvuFrX0EMQCOrSKwfyVpaM/8
YPL1IQpFmkQjdiswGAwO8G9RIfJ6aYehLOzOTho76Ao9aevDu3b4wI7q+hveLgFga2iVKP4opS0D
a4oSHI66UfI1tC1FJ4IkapAbsaI88ctIPooU8IocoSSFtGKhMUf3OEzvoE+MrTEL/SaL9rVYWCeY
CAGjQffKAzCuz0WwD95Mj6M8/6QNAalUeg0K0njELiHhItSnwxZ2sIdMVvXyxLz0hGi3r2uOcjTR
h7qYXyMw+mGir8RUg51e0yRzlcNCEeUcweJJuU30FYcaxzuAsTMrVq8a1OD+bQbOmk2amB3LpoBX
5awc1EHSMCPaWdHwzV8iGF+Az9vavsxwjEQ7k8TXfQzhYMMcAT89jKmPd1p/ruH+ZfE7RvBPxQE8
zq19T3KkXiEKpb0dHNeRfzffeNcL+Zk2VJtYOoNEHgispt8v4oghaMCLMCqR1FwZFEY/jlx1qBFb
Ao3bvvWyZ3832JFHd/2eRV6B/K5hGZCBMaD4BGyDJCqZAh4oMtRewjiACZoPmHXe0qIaUwFZeanm
9C8OzWcH4NUFKQUyZ4WNhvUIPN9STisqUBN0njGPeP0Tt1VeXNCRfAyZRMwSrHTq/VPXllhnq7O9
Uo9/XFxFfJJrgNPeNXX4F9jrSeNB1zvpyxWqVQLoXN2Yn0IGCsci7lSqcdZkHMf/MOw3uYHg1XyT
Zno3OZfhGQxbqQdzs966djbZxmWHfKtY8B6isCDpE7pD/sF00yrNbi2Q8ve54Wj46rQ4vt365LSW
UMkdBZCXO0N8NnOfh+J0/7JvXvTdelieIb0A2LincgM5wbNW8VxeUWAsRhhxplivBqrW4jMizvfh
EBhNUnU7SsEtGfgiyNHpVRIbIE47jbyPYr5/sjS7kuuQCmL7u31/SdAJvuBsSp1qri1cke+OfwpF
etu39wnVMUzrT8A4sWOJe744kPSUyFzQX5REfNAVERhmf/RedrQAEd7lHI91INwxyqyOnCRzF6hP
A2SFJP0+aSr30y+DbSoe0MasIMIuvWDDG6LtGsVfnDgrCjqmJBaqrQDGCKue2pyOV/Hqmlr1B18z
FOCmziq9SBiDPPrs2WbPo/hnRvuwUfV8ZmeF33lOZe+YAimKxBMnGNkGHb56L/ZIY4cqGUIDxw9z
zJIUVqbu238/bEmBx830K5HrEX3whJSiw0kj3jGfnYKV7JGCnJIcTPEfeJ5lSKna0ztN2PGBJWUd
euoKtPPvYcaFekg6T7xAKeLmwBMtyPWF09bC5lV0AQ2CTuN1uNOWZdZggXSrSEMMavfLbWa36PIO
gDX2mDx9CeOlevqVZs4QAcNOmKOhRu2obXwqOoXPfFBdPNTq7udBY3rLlvgnJasqGz7XDyzgkcxG
+c1mgn/iwk5oZXyMD6tZ0QP2d1ANa6ZbUeP377vb3GjJUy2iUHL+moLdZSUqYULGWwyM89URqqaz
DDA9cQEparFZxqAV4kOn5g850nVWIEz4D3nORR/N/xnS+4ZWoM7EYlwshnN8PFwYLqAklhL2X8n3
6FXBJfKxh7qTmE+75oao4GhhDg+jmtazMB1b8x9wRH1kBPwPHo9Yqg54SOtNxsTbPBRohBnvCqoz
k911dgUK4lV14PMLeLWiS3QCfg870C2tznUxl3Kj8OfXB+AlA10WjH9JjSZcNX0Zf0td88R8XjMn
zoNRqYr53QuPKz4mmMbU1AvVsKMBUEekBsC4FeXTEV0SskKpzLL2fnYV7E2Pac8wnSSjtGC7Bxoz
V5zTNHqjVw7XaW9BYowsjzaB28SORmOALM2zMscxSaMbwDo0OJN/G8Z2+ahWJJNXHnhMIxIXCQ/z
ubB62P3tjELEaGJ8bnougGQpvpeo9n9IK/jIP3nzcd9pod3Ck4zugOJRJdijI6WrexeQb2c9B5ei
b54Fn/I80B7/CGFysdxNVquwp0AbNSDwYbXsoMZoGZt3p8NEc1Ps4BWcRDItPERZuL4YV1yzJSEk
eR6IEev+BXShxuZbuaYmy5JhG0XXRVoGz4dRi/KONjRr6IP//gyZwASjHt2XZZvWbNFi+2c1JRrB
v8S+fp5IrXTVbojw//IfOYb48/CXrFVYloqz+ZFjSz38A6hHgzAOEE0Jc+G0Yd5ZAzLGlHardOYo
ZAPvdO6KGVaPuiRI9IqU2Xcb+YphxcEADJhqqsivR3tH3azvBuQRYn6nYmzzvcWYrZAnz/u3pPkI
VgoL1p2WNB/txcsO/ui98kvYSqVTg7SCkkrSvR4Vum+ukWEgNV9/pYWprzP06DncxIAOQLqfJp54
T4gDVzUrY4cDrBJnpXYC3oMCQ/eUlJwd3RpH0BVgWPqtdZafl9lME32NEW89vjNCV6jsPHzUWEux
l0n3O6eFljIgw1Rmk6xAiW7WrDBUq3Gp84H1jx9h9QN9M1liNg68qcT/HLhvjL6Wc694VAxdzoFs
XYYehk53IWCNedX2Vs8sj024QRTG2jDwYqcfCZKWgO7nXVhLCmykk2xgkc0SPcGQS2kpxWu5E5On
eYpJ+V+2FqYmNHfQqLl8xC6AgzTvM/nAYq2lD7CA/44M1s9U9XILEIDW/FH3MqM12GmSYoYlW1gh
Khkgr2cU9nr6XvCyQwpGMgLzEJOFah1nYExXrjI01Aru5ldDw6GwEuWrfU0gJ1tDKP2fqZRmoqIE
0b4v9qRwEdjDnROYLhlJicSNvfD3/7yTnIkl8cQoIUIolJX1FtZZ8qW1ibMSEAiQaa5WI6J73I6R
SYgNpr/FEUKIZrl5X8Ca22TrhICr7fm03XMFcjHBoeHwGYXnSTMYW5IT+PTw1pZS5M3NGbP2mU3o
18HziPQlTFI7vLcrNkJBdMiHwUyd8LjrP9Wb9SurU/eB8gq4InjPe1WRCmKXeZVZABBfKmCi9wf2
BpI+KnsmAfbuJF7qej8Dvny8FFEF34pDb65QjWmil857sE0OXgI1Qi6AT7qkJph3IfTju/wSP3aC
Kd8OnAfor12z/kKwk/77WYzJGhawDJW3Mee3+DgkYDvVB0kaLXXtR99U47KHXM3yLg1ptcK70/jt
v8pKjxjPgYeighRSpIlJm+ED3os1Sx1FChaawVguqx/WZVrDP0aouu7U6jvjLMtppypyKXBdujfN
bTi5zsLzEAdylmD6mqb9TWcvuGhTem1C1/eTg9uushJAMu2tSuC8k4ULt/bSHoR/T9HKyQbU5UNt
jOPztcsyMaNHHCL17RuA2PNaqgNqO0lXwH2dsMB0XI6UAk6TeFKb0yns/Bv2ZE2AaKtqJpoTPK5W
/0HRj9371Nm8IsxD3lLDSYvJjPtX1WVkl0Hb6bD82zg6U8EDXaEjyuRZGQMiySo4rY1O9AtNFsG4
oSOQ1/dni3wl8aLlE6sirBn8GGam9p2zXd1x7I+SdSrxoMnUZF6ceLOSBfpeld0wehp79V9TtuBx
BVl6mc6PhSgMoQ/TMEes9iFeOgRdx4k4t55BH3EjGlxPdj+bHFUI3oof4uh0xKQY7bBc3lHihIIu
fxOUnyU+erWt+qZ7WWczTIThu3LIRkBbcz0ZkWA00jK4sO7QtALpavHgbgrMQ+P6t7La6PBrOE/I
1RByQSrXk1rYen6jEo1Q7h1cepP6jDypKYjPpDiK+NhOI9tbsr7NDb0AM3dEe3AFmXHsYbzvzS6L
goVVQC7vokXAXZpdzbhwm0Vwp41ClEyEbmeXTujg5Ybx1nW+Dk9CjtQ5o5xay3XkcWEA30Ht8gnT
bUD5BzG+/NyDfS6prrrpmj+GkRdPYr7snAHXfL9BgxtkUmrBQrUZXfgaSQW0Oq0JYthFaeTRrY/S
rZgKMer2/BpXtxwCHCttz2aVg8EoDhkzKkoekczB/nl8SkmcrXudYsQTP5i78lWY4NBICtOlId85
rSGh8FKUG83V8HCT4rCvQD08yg2PrLN4/+9rHYyOY2K86kOBFVAlsRUeSzZRSDvpw1twMDnmcq4M
tmX+SCypqHn8+4Wv5wEElSyjXVZpOTd38rukHKmX5GDIH7Bm9qP8DXXAVgF4kBtBaMapl0BMMFzi
ujJXwwq5GkAH+A2ywDfbrYgjzHifepVaPvuat9Plv7H3YTwApkyNqbYw4IMaJr5hx6lf/3mPBulz
fQUZ+1LCd51wjwGA9VvLwsZc1T2tGo1Isi9eMXpuFCAx0V2NVopx/T0drcQv7KOG7QFO+Ym0AQlI
xjLynQ1NwEXpgV1iMfCroKtlAoDNtqmSSRs0W/6o0zfGEe5dNkXkxtmGdZCWw02SQ2w47/7j1+V3
pYEVzQ+4A/uwOqlltnnAorf2lEkoniUbRbJ7lAyvmwEzvPD7zoqz3S56rvME7f5gYgTbxMkiNaRU
2htQbLPx02gtN1mvZ5jotCNmW7xc0S+nNKjvlUoRevPa/63pi5bMvPhq9+f86Bg9G3xAUpVIJWM6
Wyi33aQwQQPhnrCM60sWSVfMkfCWmX7Ngd5mLwXgCkyyY8VHQ8lGRfZrRw6F6vudoVJcbWKMUz5J
uoHrvlvOtvsb3V0YbJbngZhW4YlTVJOC2uDL9xgjs/eVreG19WCOc125yJuceLt/RFcS1+jw/lzf
m9BiYGsFxE1pavrYKWZs0yPmxAZ7W5XY50WrPKsjSTnNXos34HpdL+1VA6y9WsqXMtzhiX5cnauX
I9eJNobaE6uBhMaXkwVDImhiSUfkP1Ma/V/ZOVLaUjv1PD2JqktS/RUqLvnKzjl2OVoQ2tJEcppb
9Tvt85Oi8/cRmZmjrSLtJpMm1vfj8288If0OmjoNC073epCjvaXNhQIJtYrR4isErzgONr1l16ej
AS5kIOAKcOZ36FzTCvIDc50M5R1CclsUT5FZ4+2koc5vpcP7YwQOHa95aTzYuSCFDUOtZQgZhySz
l1qUbVrwbYnXa4OAkLkidHTkiZ3LGAAkmyRTD7e/JXX+Ln1GAPQyf47f23SW6PxSgCmcd4f+4oIF
B9x63fSZ69Z4cs+udaAJnaufdZ5q65FV5aZnwR/98XakZ3gc5vAORA8lFXqeiAyVZBaMb4ftJmN9
IBNwZFRJH26V5/dk82tLFD0DQnXH/HPf4LP6h4zgzouY3yk0dk59sOhB4UKK/GAWW3oV2DxSmzZm
gI8rf3uo4KryRGKuHbyzhF4+KFPfC8RgTppkGs28cxCx2nx9GfWtrBt+fEXYvNKkyk1firrYnbS3
sZX8OcYPOdIOesCcAT95Hz3SnSZAgU8H45nP98eQYESCFsHQiG2h+iVRwBHq2lR0JbSBfQWIitHB
HlBEqCEqJAt+mEpuV+0nhENhSO11p/Sa3hrW5ajKDtECQslZxR8BrQWfYSh1UQWP/MyD25q1mbxA
+CWepkp+G2pp6q03laCiV6hyjwClH2JB4HzzrQWG/lDmEPTFRliJEVgKm/ZJ5Tbud3usruew26Ji
QRpkAQShXiJI94H+AvrIkXr/iwNtBw8I1iZyuh23naTM8C4F74cqwIwzKdIMlxoL9wZprUGe6yfD
hPaCiyEwnr6CqdoCZMwvwdD8qM7S5WSx51msbcuZxY3592DJRMmvohNgEOklZgIy/btEJscFf3Oj
MfjhHNFeUka5aMmRbJ0gPfcQaf3551yT2NT9UeQfySZNx8MYoN4rKBJHBSYLekqIAh+KZkEdN3yb
1PM8416JwFCpag4EPO+0MED9SkyW0/eoXkeSD3LNQuVEZpBWZYXEzTKPuBBc0bIyB1kn3daIlL2b
o6niSwP7TDgRnPYyhZLZjKWJv+Y2misZiLKIbDEvn/KJ+4vyVhOFo8nz4NG3Oe22SCtXDm8ErdP5
eGFCw15Ozq3Grl4PVeruGmO4mWxi+iGMG3w+LVDYkBrfw6wWmbx9luJ2ovaA0TikLKG7RtWTW1uf
8wYPM4IFtI2G3t7KV7CRAzrmn+RYD2BTdkRtc9jzcqlzMFzVYDTyfVaxpuY64XWHI+z7RcthdAUt
Dpkh8dLQC7JqkBLJ1u1XnQgojiG3Z7hLam1a/Ci3rh9ODEFHaKqdxiU+QTnXWUkUqCofaNN3i2fo
AouhRNf827esGewjdaKRznwHNk7dEoI/zjJewxWdCfWjPSAQsdgF6bQuNOANnk4cmBPZ0zTK5Ieb
Az/zqAi4qrRZiBFboTKJLx1icQeYzn6LhcxZy3uQ6x8UHkVYrxzplZgyJlEKl61JUy5Yv/sZnzko
PUQYfLduelNENegHz3qU72jj38CE7v79HhMTtLPlJHgqo0NdE64gtCRsl1t1LviJqFkrnuEKNKbk
ktU7oEmGZO6rzp1O5fFpka+xqK95VUbwYuUizN+Apj3xeIOAu8151gHOJk1WK3gBTmSzHIL5D5DD
8jRWsrjlaMppeid/r8X1rswItNhlZU7oLM4+V+86G0aH4sAQPynUFTojguHpIjxAzBhIcWICG6Gs
5sBzjB+8gOaIthI231oikq4FrMv/32od5VlSRJfA9kizH73HLIcm5UH1bYS6K005AbjwMGupRtKP
ypl9ib8kD4W5l/4sz6xqx7Ilpzs1aPCYbccxtWA1Tv5O0lFwC43iZhNw+4lxMsSar+w/WOCRy/ff
ctMAAyJmniOZdBJF/6cW36uEOl8SYR8JLVLeKYj4Af6kF72GNGyyyXkkHM+l1wASGuBLMy/j696S
SxE7ioRL32c4o+f0ic92OoI98hVqDl+07S8jQ0N13QTKqgElyRy+Wk2y2HGlODJArnS2Ht2r0qL+
czxMhSka00tjX9tA9xV0Jsw1hr0WkPd8WyvH2wrLAhav9vqoujM3S/HqYPPrQwNZ0P4bHPIU3Ff+
/urdI9G0iFRPN9oi+CdWz7x8ubG0+4TwqTVhXIQWFXySjF85qgfuTb1lgKrfwB8fQ699C3mXYtiK
H0lSlsXCTOSEUUR4iUBtqd5TjXgJzkhp37VvaILtLEfMez6RjhjKMoa0q9f6e8bhiDwPWJQYrItv
6eLK53JTqmtgj6NKU9BaAjSQAnIBmLRK119/aJwxBAaWz4AED30rv5QEFcXs4h2sHKJnW0kwePpy
Chkx0gwb+p93A4QSwKv0FOGJXRBZjIrYc72u8NYp5n9yHdhscSXMyf3HmdPmu/IuIfFCaktMpXkG
3vNxUCOhPlpCowLsUabPiZWsJXkGS5NXROvS4ZBdIt7hG8S1I8i2QYgfQX8bDY71whzftqXodj3j
zHpuWrYA2NQX7YU/ZvTy9FJ2PoMxTI0MNjsUAqti/KjCQoSv54U4Uw11KO1PM3PfHurm5JfXMqhB
FwB/UmNl8UTY9Gm75r09sPL4yfQGX+ZbmMo/gHMXENfEAH1CJAIDCf6AxwDwKWzTFIUj3K+aIXJf
l6lBEcJARsyQfqHJTbFt8zsBdCnNDfzQp9xEWEW3ZkVcs6vZbYp70ZbeV5hNMCFGUvV3MbsGTodD
ycC6+9nb9tKeaedVmvbWHoPEtfgpm9Zft5LFDFDqn8oTWLSw2Dbjh0BiHOwmR572GiwFEetIaxTx
V7EzQ5bbXY6j1PaJwzA7rX0vq6YREdQ9q8rxkDpfErCBGtfnijtkyJm16X5GmOzc90qT7/Xe6fX+
W7gKbrdbwqfNxD1j2YMymhJDiEua9dKhp2jj8KlN6NZCCVDzY9wHCURwjpFsQ9Bu+VXJDQhjLy22
Bv+/F9h4t2vi/2Im7wvLRIyavIJ3usP42d7fp2vwE/2lgeirMb3e1EGkfHd7ymtvFtvVy6fjVRYK
D7yVyDk/4gLudjxZWz0wsVpEFbEcuqWFK2tYwqb49sKwQ0lyEIKW/me1jccrPm/5qFAtIuRHp1Mp
tM7yRJ0+z4gWYL0zFkeK6xnpg76SPoWyirEs/Z2RLKgIgZYTZBGc8fOTX9f1YxesAMYMQE8LHptu
1E+dUCbNT10rkUFtDG8CxRTPZ95u8khUUAxtPSGQIlDfB2FjXQ82Yd2thwzUs3hUHTMMDPEJpN8c
Xgu+Z+zlYogBtTba9wtFDzpcIXRl9z+AZ65AoMx7AKjwlOnXT4q8GZYD+JloD1XmkC3hTs/Zr2Ab
xi5nxTUmguFloVX7+TuG6bzkP2SPW2SyLPGPhFKNcyR42sn4qWJ9M0v7Da9Vfrct0xNsTwZoKiJs
+NrtN6Mwv6tCHXdz57C9ZNaRtTe4zLASL7w9ynMQMHM4y3WV0lo+v6PKkojYQ7U2JpQrY1L+PESZ
ttHZ9gygBa5QWrPGterh2fnGcfyx2PH9ji6fs4oEr00Mv6lI/P95M97hFbkt+33BwxgivjlkWnO1
ihsUEV7Q8mEof4H/4x5VgIr/HnNhsTIQ5iltyISvh7WDbtpfWAZZVGUPJ0nO2HKiJaQkoyhcZqQx
mRLLNsR4FA7aAshcS8MDM5rb9nnPrq41pgLV9Nxhkc3sJJUUuVGwfABvAOflxnd0yoQPOP+v5eGf
pO/mFyLOM4qifgfQLqSdnVB12TC9cY95m4HmSJdhWMxX7YLG9VxxjBJ6gNcTbIt5/KslX12eVngm
SAjKRfOblv3SvDJNHscP2WgdvApRI8Qpwci5f1zUtexrdInRPAXxvzpjMeYpVg7nfP0vehpRyjh+
/YD+muPKG4YNb/PK45bINEstPLM5iIWkex7iUDCaqfbamOA/oAPGY2UlOxT0U8TMDSGQ8bgs1JMJ
BR3r0j8rwALPl+jp7ow8XEL3ppQYKZ5bf2O+5qHuSqsLCHlOXKpe02Pi2U3r+tw1uKqOygINsXSt
3YxzknbiBEpvBEBUFLP6TD3x49r4RJ1wL++mkDpBmg8o4KAWLn6REl6eHeXNilwv0Uy/6K7PObFp
S2WiwH/G8jR2f4hz6l/tQo2OFN3glDTUsBYTP8ycjsVRkfEsAP1FQAo2Hr8VOi6qLmxntuWpX1O5
w7fkRZEFx+fB4UL0iBB5Kz8GhPGDL3gDO43+APo6Sks5l2rfevizV59uG0gUJKyU8IZO9LpCJOJi
QINTkiHhoBjlE2LiLXJFrxov5bNIbtr379TBBQhqWoeHb8v/OxYxE9H8WZoPyoqAOWOTODVD29py
c9dfJn/quylg+YBXxNM2UzRNzpaKulUP8xBmaoDHLK9YiTgnEBRjPlIOUG3EVSPX2BATjv7bxqGZ
amI7kcYATUDyGJGWdGn/KKCuYpHQAAP2pyVBlJT691b47DqfFXhJekw4QrXfdSzFK8lGXNFFLKqo
nYq7ymn5xjbh15AWc39mJeHH399+XC4NWHSj06eAPW1bFZQIPKuGYCF1qWIo7USqCcQkNfSdoutv
UYjXZTNyJcnpcDZ2oBd6L1ja+/SLbRwOI34sP1GCWDKbrok2NPfXN/uZk9+TxQ1LNizTm7Z/2LHb
C3o7NTNnNksBxAG+mekGhXVIqfN/ztU+ZRWjowU4fgTW0VwjSLPeXcK9OI8BYPnydbndSCMtBzKM
LD85svonP+tREBQmdbHfC5XloUmJiEouPUgXdT4xvnSXtfnVec6hmwpGjwfqzHRr2xxUQmJVMUME
+vKSNG6MXlau14vSBei7ZpHpTUZGcH9gD5GQwGWBCTyIcuu6x3QCvSFJdWDoxni933Q/WMBRTGCl
4tcvXtKjfVMu/aaA5lPFxsy4tmLLu2uUZBVxkEAnZpOzuRJBk3MdDvoVG/OWMsjz2dXuoIBl9RAF
2Bs35oOHronerIlNq9S2dL8s972hWJyicYRnpjazpDIaGUe77OKQsWlKCR3rxaZnFMHt1pUpyZAt
6rvGQ9sFqodpsVb0NK7UNC1Ku+5KJMORIaz8k8tqk8sI4i3xAhJ+EmMgab57sn9PlVGfD0gl2JT1
qKjqzbv4s9U0vhdPdK0UkB0F/umwEcjnanSSnNiiL1q4uHdApIfmsH99rOYvi8vwMaJqsiEmYOUu
ctVgFsXHVcEKdHZ/AkzgYJ/HxUhx8KArGOvBwTJp9xUhJrhmUudYuAw/0CKJ7vkxyNiJfUDT3tV3
L7RN6sqSszrhKLk5pjlK4sjVVFsD10avbNBkAYKMEi0C7GiiHbPvU+aSjl2z7EH9AQIK6YN5cdbU
MRS919QhhvvWK3G9P8yWWXvqgRT/l+Z4cajE6n/utC+o/yOnV+B5xGoVmzvuVF+fcMOoIMpC5G8j
CO5L+pCq5K6sbn5AOemi49yH2hmTfq9/Qv1w4c7a5SjGOxkqIqHeQI1hWBy22V9OO9AkhKqucWtq
+uVFHqB4tPKpXrTRv0hcWr0asfpOuzbce2ibdzbJqdB9nnVvDUVsn/MTGSJ6TkEKnyvofFsEZgvC
MsRP0XT8cw7wOCfggddb5eCV2Q5JjNN8R5MBdzsUTiP9Fc6OF3b2ZEbUam7Y7Xaa6V2zp7h8WiZX
R1CpmFi+koDc5KufelWKz6sa8Q8GuChNvNpH1t+PipCeyUIHppKk/s6vuQWqsOXeGW9TzRyTQmRy
nvFqHGwvjjJTZ/I/oMXJxsDHKofEvUH/QAuQybHmxT2SpjXisGgWRrN8O3qnmwI49v5jR2aTn17c
bg2onLkiiXun/hiQBkLFNwCXQCmPtPLpdHuvOOaQmM4KR3mn4Xeb+Bo3lIZdk+p631Vi7Z15VxeV
EqyUI1pD5o4zckecllG4hKl7uE0PdjddQWI9+glwofG8fXqH6p3ucj3S/9lagCJhPS6ORO/dgv0K
/qKOgQTgSa52ETMFbSUUIC1uM/oglv07sl30NLnU3sZXG6FziI/oLH1dUjrhHVDvWSbZRFiIkHDq
ig+MdivJ/nIRc0olwglP9IWz56ijuar7/AIZrlR8brsJuAPv401HBg7z9Xxmaz6gez15DQvi4ezO
H/gcayX//ecnWwOVhZPrZtd53KAv3M2Y5aTevinWHoiH2NhMGPBP1pV1RU8O1555wnfyT4P/kMY4
kCLcYbLoB2kOMc5byUSYQ8Hkv9UyLMQc6gNBFd/hfE6Rj4cvmvCGrTXnojokdj6zXrc3QCprLxUS
FH27FCD0ba1s6hpnCR4XEf+207l/3zn3JZ5ZnNWvp6FfaoGSg09+c5c3QSk9QQHB3qer22uXk96N
B7HyAmw9dyDPhb4MS8ujQAUwrqZA3d3gcRtyPJnD4+4YkKXMNlFarxSQn865Wgllg7tXwzclPxPB
XVyBd2ydHQ1MATrs2pT5Zbjigmr43oRtGxR+jPUVBwu85GRLFO07SVXJgdOvFzjdnY1DkOAdwumG
gA7D839XQI89CsY7m64EBcfUzLUsmpH8iPvwMqXUhrRmdjd5CZCrG8pU/O4Xm95/BIcBFovHgove
Cn4qImKTG371ONv/dDc7/01DOiuZYDYl2qEezOQoJBmVa/bQCCA3Z3QA2l/EQkmBJ3xHtJUDUWFJ
19tp8MbnUh3xcPEswWHmx80dL3iEekeCsv+iYMaGqBjF4rWefSO9JrF1Xn7N32xCj4zvqqaFdacN
CnKZg1xAouClH9KDsXUz7vkNQLhtLCtfvOC4n6JWOfkSyGZe8l9Puccx3wDRTOcs4KczJaEDctAk
I0tCTExUeKlTTQCElNEQFKUDEfyOSBFENyprT9iEmChbkJtrG5z9VPIn2OaRmKQTqurXjNREWKKs
B+o27ZrH8n0dFjqN4yq8BJLadoi2MEn/8rC9W7InQevfP/pWE1jhN1VXYYZi3dByPKjzS6wqTlWd
nArZaVpf7CtxCOCI5VQmxsFTCAY2K1AUfJdQVBAJpzY82cQOfpPnjBXi+FIXAm3JUcBYt1XQfhEF
7rBmYn+yt5V8Cn8NdQnUeVUbwDLs4IY51TLzHb2aJx9gOc08hbEq2IECRl/O/J8nRDmdGD/qxD3Q
9KTa+imioiVAph6CLKBIoCTG2pZd1sEvArbN0nKX0Jcbgs1rE0f7lK/wIeqLHWOEErSxgv+nUhT0
tjgEm+o8/HDmc0274nj0glh7K9PvAxbsZJuUrZC2vVW+Au+xwiaQwUNIWQHmj7ywU2MTUyOfBu4f
ZBeyiajlQZcYMGSEyYFbr96McL0JjlZh2SeyRLKNQOuFruz/2mcfYD03dVtNjhtjbUaG8hcTWZNb
7kCZJJpsZDa9Ln90nTMQAyg366BfGR8H55R+8nIiu3C/rbY+NaNTeXiccSJq+Ia8o1LtnHTX/jGk
odFAgAQBBg4gE3GBsQa7mcPk0giGKjOxwz0d8SUnxoS3PqMKez6cQ8fQDiwsQ/OXfeEYgYHOABZu
c95H9/NCzzQzZvpEePrNWWIBD7SrXb9bCUluDernPsOthszlzXm5tNu5ZxWnuGxfsX8hDz07cjyK
IqjxHvlV1q3MvnQqwRcpefit+kobu0lRYuxLx9BIpn3lpBRivcEJqQqW5RE/XxK9HLtzS+WbJjLN
80SGua3iWcvs+OupRlZxqhGc3+7rlho8uEKEIbo6/UOjROpVf83pFS2JCf7SaQvSNFtGGkOlfOxP
KUJlgQ8N+w+ZCEzT3OjNndLzEJcCdsTk1abyNi1t2U4kjDqcd1tUao1OVMieC84MVx8WgkZTxd5h
nGKAwcHYOd5cgSoozeNSZr+7lHiPjQ5+Tziht/SRaen8sM8wbAm4LO5tv8XaoGt9aNmKGYU0xooX
4oYBcFIbjReE1nkHt0bqpx8WHj87hsezAem8L3XmtB3IW3ZopGpCKEkEQOwo/qc+XUJfPJxsY4UA
VvsaFMLiOPeSFz0nJnZ6Ual14LgIqjKShxp2B5xLvfPbTNy1ULn2MukY0SW4IRTpm72vlvlo0NiF
Z5JqM8qyB9TfOLIqbg2u/5LVuR9JUQkZsHcROaPWfDPbaiPgBFGtTC6QOqpHs9BgryS72RS/etK1
ZtDbifL2ZEZe6W8hjDF2GTnf4pLFiGPw/iSL+HK6ZAYDICpvSmyDA9nUZrUKP8KjG75pswpX9/FH
Lza/9skKvBo3mErpfLPV4ZwbMTofBAPe+aZ56jXb+pcT08mQCkWuXIJn5xeB46RkxMhMULlUyG+T
551Jvf1ze7fpy+eH7GM2SbBYfV/KD+us1vkesfLs8vsWpaZ3C9gWumx7bAU7jgWHvxOvcF+J2LgP
TjYe6zkPOCO4abRe8Tf1mVbWXYj/A+wcSS19aHRlyFJjMA8XUIcY+pd04/UfPHzrfZTqVr1+Ob6t
iSRB+XJVIvmPG9n2pWeKRcpyWH0XU7mNR72Uz29q4nEGtDDk8RtXg17OTyzzuCc30KiynlnPa+gC
7AX1O1ScIzUICYy9RjX9qJlDO53ltC8dZBADrcaBbcqK7WxIy50E/PmDlWSY0NOtvDwds8omUV8b
z0uxXkZ2KYDeh6bmjXrfw3u4QMYqdIOe+OkHZN1ciUaF47H1S7n0pw1ioW2p5oR00BUdo3ZCfr4C
AcHrGfLerI8jeqyzDgLjsPZWeF1WtUvLVTlpuhI3p7ZoVr2eA4bvYdIwe3qn4Mi/Akxlkf8T1m3/
DXy9TE+XUzpPYpLomVCNe+GtdQqQP0mH5F5nJNKaTckoeocg1pFgEQ6Thl5NwxSvH6uOzqRblk5F
Br1tVx6QUYvxNZXuP10qyHwfypFOOTGlY7R7I6zQ/pBSgo9++bUg7rn4Al0TOCSeXgadtMLvdYKq
dxS1GnSG5diaQ1ySazd+bcdrkLomOUQOL4A5Pks6pnkO4YaR/qL6XqcioZ0rn3d5e4g04ap2xSur
EvF9OXW0txO72fnPoOOb5KDdbEvROeCLk1J+ZxHQpHZYM8pY6l3rqS+AS92aq7aRTJfsKUTmDVNE
OVx7PBhtbcWI7QSrJq71dZn1GfSFdQwt6CE0AqUNa3tydPPyqXl/cWv9KTsW/0YKPzSKVlGo43UR
SQ9PII8znPp4KSe0vbhAW6Zl126dGzK68bXTjazRf88Xs0Si/8RWBu1csuHV1KGYf3VwVCXq6p0Q
mJuGW6ebU7OkZOS7KAXCiA9+u4kPBVbJoiHsJvwZGcPwU69MSkXQZ5dxEcR+Sw5gIyy1O6gtalMG
wn4HmnqWSy//itVGo9G0b/5jYZI0ImUKwn3U3CroHBrQQUZ+lKxX7/mgrgsIy2tj4s1yrdpq1qad
6LnoIqD8l/dD0MLGS4NwQIKk/OyZBFzCzvYXECpEhW5cp2zyULn52822wpmj0RJtBLf8n+AbZj/O
7Ddg/IdiRDElXRKjFy11gkwYrxw8Y4gauJnz+u9Ys7bXvgE7OoJ5Q7xnxp10f458g1l6s389wdZF
6m+laRcQX4uEBtY5SRlQBWLxWZZKd96p1nLmVSIj1atj0L0+F0qCPdCd12+VcvZ66X8fop1vOggQ
5yaAs2YYgqZiPZb1wZ3aa78boBT7uEWJXtlmBDt5UZiY29PDMfurG9Gzk3fmrKoZH4UJ6oscH8NN
KD0qvFw0i06Sbgk/8O8MyHSq3W3zl2meBWPTRQMNVqTkJzVLGyo6Jkhi/qtu4Inrsc4jwvMEcqT4
kGWPVG0SJj0sr3IX33lnSsAY+HCo/x9ZzNizqPNkQOS8tgoL4Khjhly50XEpISaBk16D6+ouJy32
QkWBKOpiA69N/tv+mWLw3mQUpuft69fZs6C+1/fsBf9I/9XtWiKcx3Qixm1vjvDcVxNcwTjEgqyS
d93q+eW8XSGuyvVx0t0/onF1yCeiIBF4+GBKa+qZ/j6SWDiMAXRGlVE2afYrsdKVQkEsfzKqiRjO
mH3wo+zDPxu3OwwA76npcugKD0x7F0pVuRpopUizdcS6c1ZaLYdwYYa3KHCtuk7n7Obz2doAF5u5
62uBhsVqGb+UyB/1D9O3UNv1YoT0rGCY37iBSAz5igRcDObYK94mVPYHcnVhuiFcNqriiMlygc+9
1rB+kc5uOER8fl4fTxUwy7n43kpTuaoVMS8wYUobautlu2UVA2PmnSInVyystr2rKW4rCmEY+1Ib
LV+q1PRvXODb0KLhn+OzYCzh/A84VnVDyKBZdILPxpCeyco21+lepE5qWgjh7Q25Z1POlpMqgxdr
ZxT6Z44TpwwbMuErSmHb3savA0JLbkwcYjdP1cAvEC+FTmdSD0wZO6z/1Ei0M5tyDNwUIwOLP9Vg
48brSjAtplstOaN5G0t3ek1GJNdGadzdb5HKqCzopUEUQblvqcpeoxWtBPdUrUU/o1h41XzwTJWs
1XftbEN+NgRXZIAMpDw/LSrnjJ/6GGAhkpa8VTifRXX8OB0IzHUvZJ7VOJbS2qHIfGrPMxlEtPCn
8XD5T9leNoVLiIcTVE6gvZEb7VJZ2lii0UKkohK/2Twgp0FDW7EK41gUocB8Uofe1zEjt+D4l0IG
Nk/dG/uMf3sy7wiaZOeBD0Xiovaksz2YANeuIEn+/amMYQyZp3B716DzuelHDo+XHIikfoY/PNRE
Y9Pg5RftqctGOUQqVs96r7C/QZW4MmUdmqViI0rBX6UlAUig7JKMkEPGTtHMPu73r3xYlk6bXG25
ABT6E2zQfkYFphRcZhjRAq6uO+oSkwyZfV64s3vEt/YqPlHTXmr9hbwBtKc1Qgz7Zl9r2L734EKG
rW8nnZolF+W7+DvV7uOpuq06lMmc0VT9WtrX3qcPyqxY3LsJ1mHKQpX86eW6jp/nwm02lvusjgyg
71OFqWFI+0odYWlgQ4Oduv+Adn88Jtw9EeljQD4Kzq48Ixv0/d7WQZBbUqP4PkMcQjK9co/PWJqu
77UdbRReGqExwXXXCBkx2krna5Oh7AnHP8ZSONe6fgR14Vnpw4mlPGJo9iro/a/3GrpBbIsnIExi
HTTSKpMlWUFi07fl1QobFjfLP/roqApO0vODOsMhZN3tlptQ/f0klaAUVvdgpEFx90WJhv7mnijA
jbLn4tFeKakU3lVYIGq5qZhXVqKNRGn+5s86p8wsu7IarBZjOAxgPae/FdYzsRjrO0awtG44qHZL
4EHKyPZb/btcNF9v9S39QifefGu6P7ZW2jKRPUtpBdoblMTQjcdirqlufgQoPAYa940M0iOSSBJ5
Q+T2s1V0O/jmGWrES67HfeNUoAq6939mEixo2Gwd6dqjBr+xHKSmw9ZgrnOG0zSgLsoO5KcYYS89
05I2SxKW0jvAjIYpFB9dhDE2jid5Xcdki7H4QeZfXWMInJTjHR6VbepXbU7LlB45UARkyiszdhAU
pCqJjKyTHmtvMdgOl+Iara10dpJ7VZWog0HFnaGFC4lWRIlb7+cKBeZ9C6uMDET+KGCZFSTIj1d+
JlOtZ/p5qlNY7JdjLOku4DDmvP6DYDcHOBAXouPVLCU74/wqBAvpDaRzM4v5kaZK4EM8iXrugDEG
RYbZn1l8HqMhgw3Z+WEKy7GKlOK959iInYPOXNvQ8dPAyzun7ZDxV4ikFHQzkrtF3SdXjedsiMmY
7l5hQ3xeSbtkT2ZVcsGgs/fI8gqPJDaSECyKQl2EmjZG7/vjrzz7ls9CVceqQ7HH4Ef5ApR4DfU6
ClU/KFpQit4+uchB8BlEAXNoV6B8KNtHECPP7aKKE+qEr+FjcnAZjzE5K5f9PSk9O/WbNAlYLKm7
zGJUNNDHPJ57Q5JoQvnsWwckH1bDtOY/FPt6J9JURbyz7TSCvgW7jG/tLGlHMAU+HmCVO0f7Pi5f
zv2gPWK0TpR+tVTYMluNbatwTmEZqzYLug7xPHNr8IFASqiw5SclcqNLCnfNvJDjlbhEEMGedfAH
1AZ9aNed3ttcxfi53CiSd5A7PScy1ICJCl/smaJnhbM5T63FHTPwrg7TE+xbzPBJxbtLJdleYtJo
B83TNKebglQhMygcDmdrH6PGzxl/Vu+q3C3m6zhUGp1+h705fhA517FsW9Xc9IbWJwvZARLp3eb/
snXJ3u+KYZuwQHZd+IfOWJE5EcTPTuJdOODwqyQQ9TqR6rlpyc4jGQrnnV8Fh5C1mpoxJ8joANFc
ho/h6UNsC6bwFz+i65WpdU+fQwNck5QmT6Q95k66ooa+7UwWLYK+1K3lvT/m+BQB8Y67UX2XA9As
Sz6bDmDbHwJNAjrYBg7pt2gyHwfpVRXnVu2qK91mdTcSpZM4dh89g3cgRlQkQK7A5fUSK/HjGE47
I6ISIe0KKnFKvKFOPkiHAtUdN1h7pfcvVCxFT0p2smoGt7pfsUnfy30Se4aN4q+KEckpEyJJ8V4a
CFTFb3M3U9YBMq4sExoLX5IwWrP/SVOdzU7r5+yirnSNIH3+w+OGfNVrXpdFtQLxt1GGk8nHiSq8
VmIR2wg5HVPmKBFWIOD/APVztNvcgVMt8Z7vhSSPrj6WafODSuX7+PGOV4chgop9GEygnjnOkEuG
l+o12MJ5EPpnwQGPbt0F7xd1gURBo0zGIuB7WyTa6cAUUG05w3LdSVyeREeUU5pWkIJOB5rdLUow
WgoBz29fFhSNYQm5CEL9NKNiIHRTwqm2vGmxCfGC/T40cXZSZoBda3Gdqq8ur/hsJxq2zb0WOKkm
t/N0KacXjWGkXPSKVbnfb0Jczh2WSSRVszB/F+K9pu+ug3NVXd3O3qnBLNVoxSyj+2ltla7+sxg2
emKTOGFsTi1uqzm6uxzsHg3Nr+HtFZ4vc1MfeS/M3YXPP/qGwuT+6tGK8fmuphhiAVLrTOES/9H0
PBBf7JNfcOD1bXejGoNL17SRh9laylxKYkss1zvFMhujz9URTekOUNIGFUX/yazy2HaiQcwOHGCA
igLbrXSnpimUJu0jngbayKuf0OHx92quRsKVpqOfPBCEuwqv5OmoqhvtrUzK4TrYqoNTu/JZSeHv
EnUHJkbtxb8VoMRHEGAItZS1475aP+LNpYhUFd7b9n3PDTtakiZ4o9bIlXyZk/2YZ4Z/7iSXo2sC
9vrcwvNjUWEt0/RuhcnyPOFW5AeyT/P0eBZNbVSSteLWSvMJ66flnil9i7CR/JQlmgwvC5WKwN2y
EjC9a2bpUDbO2SWXL1+L3Ej0E6vlEyvbDeFCbLE3ejr5fSOS0+8dUGUKDpgmEUVgLWkWY3Vh2hyo
JHTlC32n7ubK48aTYBs3vpALfWSNx/MMGnG+Idp6d4ychON/b+Nqbm+r6ZopmSOuzFpRSChTsCuP
7x0+V/MP4askbMdjHgQx9PbCeiCgJhfOmUaSriQl0L+fTxGUogiaXosVmc8Wrq2QQVJ2GQv/P++K
3Ff8YFmi/InGrkhcul+OIYFlGZ15mjtnHFdNyEdR2fJHWO6sjwSB1Wp1313zejiseuemqSli/SI6
1M4kslaj6Y4+7ri+zGM/wClm9i9B/csd5LvUO6RO34rOwodOdwV+N/x+elQpDGGpFRS76pkfX+6o
sU0v3DEkFG72oEtIxv4eBwrai5x4YrSkj76J77AYAvomVRW2Zz+MN+xYZgivm+LkSYm43Q+JCIwF
IHWNEGZhUe0Z78uDtQHXNnH2Xj9qOUkTcIkC6ODCxLJ7xMhG/dR3vSssn5cafrKOX8PWjFrB7InP
iRlXD71NpyJoEG1t+b6eUn8wT0sJVIeWe/6gAZk7XVnA3FaWt7AHsAJWI0ruQ9acrlueVFE2L0cR
BJnLkauEUlAj91ECwJvjd1u1PIR9PQye7XJpO5+evHSoe3fF97SmZuPJ3axOpu43vfTtpou07jBE
eX+AhiP2mw2wMdkS+hTtCPcp4pnn/PhhWdqHk2fr7abAO0kD2OasRiKr6siqZ6c8optbQYA1WiUl
rhcHDpBKZJOkiORixoGf9vbU4rMl/EfIHqwaKFqNN9w9tw8+ERF6g6Ybth0g9QUJbDydzHn6NB7j
nN1tvv5vFc5CEipEfA6DUpJrZSyJz2w4iocsZcjOEuNviZtjGQ8FIkGteiCuCOzTYlG/6xvHd/01
L3uZipZKiWAvJfqj/6uqnD9LcZOTW+qssV9W7YO9oiS0AMctcX1YSV8TyTNXC5bbC0nEck4Q5Ejv
4QoJNVrQ2n4HWxFOI6iJ5vDdNkgfh0r7EpVOZQLcZ+BsVLw0Z0WxJZAtjX7JhYbkZd1NlKMpOJit
d+RxNCImVlSetnRI4jqX2z4wapQErpQY0nKgSwDt8o+6l1tN6ORZXBT7RcT8XZswfqvFlir50sJj
5hzj/s9ic8gtrvXHPaX2RkkSQOaxw5sBmifJiBseW30aCa4WqvldXLBCm9EAzFCprQv2ETDNkqic
Dxv2NaxiuRwsJSDDLd6afbgxbApKUTCzYJDROFFYz25i/04GuclhwmRO97EWgF/ghsf0ZJUWfS9p
Ga2zEaC4Vi5ZOFXOiNXtWNOWky10mJ6pKQFcoMB2l/9QzlUCF076KfKC9UOtCQFOSIsB5gXuoWUT
+i8TCDRhMWM0+O0H7+am5MHcx8KhQRq6KMOrvXjpBBXGM4wUntY89IQYTdKrP+hur/3RHPWvuttu
5TwrQp+A1K6zLbnq/mwbLjMl+iWxTjIAAAZY+5c+ZYZ2bPFm4sqQsKoQlu4s7kgMBwKGsI5R/RvQ
kA93t1swisNJXVL6yHW33CEchmwX/3Gcj4Zwjxlv1guxN0aNc6GINttT1lVq1oLlXflPZfJs7r+j
aBDcOu3kNOy/tYhHmEJsrpjuQF2m10anP6Q43Hg+4qf02q33/JdDnySel7YUyWx9JLxu3Wj+CsyV
rPKWubBoWIB0yMvEFFW+j1KZZfA2cKQnC9f5hdIty9wdtwNFonsw0w2T5HPkfGAbLMUbGhFKLI46
y1vT73pcxwgRu0RVsS1psIVWVnb7dXv/fvitIfkh2D02hyzmemDz5FbyLmPlFuFHcrChkDuN9lMz
zm4p6JrUNgPEuSExejlKad/49zxCpq3fhExUJmYHaKMbfWdW+telFJCVzBFFiy9+25K9APiu3xGm
b64TvECIOxm1uL18CKJ6g7E8qf1mAspZaSB05OzFz039ug/36sNEon9zEzePA/A5P75DS7+SaUwW
UQ0ko9IJK07xkpdReC0K5isjteOv+f/ZJ1W72JD3QBvjJn4dFB6eLyy+eKewzALLINyg6lOKIS5/
tfo3VQti3l/gHX8kwcL9YDatNcaHkfa6hFR13RC9896oRAd3hamoWpBa+agPfDj5/ZXRxDm8toZ2
XB/cNINB2DRdj80p4sDo8UYug0VwAjLrA7OZZ7MPaCmvPujTTe6EvVxKDh1rMsBVGGCVcbYkEmrd
p6A/8rbTba+RiVsHu629pxSf/Kr/HCF7iYivkSko1nyCU5lF0+Pz1HfiyO7hzZXRvZSyEhPm4TcL
RmBXYegq9Kjm8+N/Mm3gbJ6bwA7wbQOljRoAfHBToUgwp4iL9GcN85JSOFcP+ECM5Di024zAWi5p
L4szYjA8b/u/fUdwSaXg/VIfrc23PYQyBmlZaW4dsobG7Z2B+UV1oQ/VxZm9kV5hbNUVUNcZXbz5
+DuycHUuG6mwO1YbPwMLuWdhd6bFZoRTxh7QIcr888SAg1od2gYMXhs9FMghEve2/OCCqywsFyUO
vg9Vg+VoysdzeAn53yn8Cqt/7SI0u0Gi2POlyfGrDBReSUrNINW/W1fZtN9TxB/TnEKv/XP8S4Fm
Cx+xsEqxY3HY3BaKq4MUrCWwuvo6EUn2Kl7Bbf6Yi0oYrx6lkkFn1+Tq+Cls5X+SaDF6ICQwPbvT
atR+47ifv4NHmFHQ4tqJndpHdQlt+J5tvnhCx3v0Fh1HSDbR1Vacx2ithf7J/i86ZWFb5mH3gzRb
hL9Llz7Dlxa37sRyuBDDDactwQFBzgk7OSzRs4xv18jPFl2MDMXd+Yd4e0drqZiUoC2Wx5nfoPtQ
GTYIqB22sflKWDWSg3sZAILyeHzfCMHtO5U8j0Fv6RZYsgddMptrGMgRQrBvxbbZjteMh+eG28HZ
VdG81VTR9lEj392LDY62+myDQfxMhPrLCQIcv2SWzl6QDhkMkRJI3s461nObTB7HN4RrXMqrqxN8
GVAwTM6XAsgr4WQoOwIqHQV86ydtQ38e7g/yrp0rZGgl2C5eAmmTp+CClLhbzkiMNnNuv1JsaQv6
X5YqmpSVyAcotwKtZPjAESlqSZW+AJlCihb0+ZtvnLNFviompfU3rrOt7u3bljVocS/V+UMfaA3x
soBbcyYFh7lIOoE6tksHl+g2mWd3SVMC09kUsEnKi7odhKVqj//dO0bjPSCb8fT7hWcPbwo8fcke
ioBXduTNmGP61xcZl6ufTjPB/fFC/TBF0MCmdokBCm9CHPI0QYn5yLZ8VcZ252Du4aI8Y8jQS56f
jd/uiRmoCdKiub2THACi0QcYu1cnQmY5MbS4+nRAm38cxtR8828Lj6p5qtxLW4nm+BvG+9n3Yh78
Ovu5+D8QTyy00K1FddjXvuaFsP+vNysiV6jHatEWkswdkaNA/VswYm/QNjkOhE3053lbYZYnHfZg
Baq5vi9Plc4eUuXHqT44lS/d3XsXrx7dLwqBE3pHMLKz2xME7BKaWgj4g4+i9X53WtKe3n0pS6Ix
GNOv/hTba0urMQr1x2UzKOK7QodWbVAWWpxO6bhOnlrK5VT1/sHzz0wwnbAyAhSe6wJMKEYQmEge
+1gO9joKW7Pl+2c24tWGR5p9Z5xqXgChWAX2gZrsrLdavX3+m6GleUUz/C01UbbiKHiWiI6IgYJs
69iSV6UPtEKYGGAsAun0HLXXQ8AXLRx7tCe/WXRfB75f/ibycGw3oC9zPDOqQB2AY3NoqrHAIR6f
nLlfDpmQiVSrfmXwNRzsSKU/uAVkAoplXrfclGuxsqoBJoG2bpv7E4AdjisNz4Y6j52/LGyKCpMk
lwgIiZ2g2mGLZjNvMQ5Wnk/wsC+zpNi7KcNfjJN2KNjsKWcqHVXYICB4bJ/Y7GrV9TctVNrMSN+N
5WzObelgf2pm/jZoL8SY6PAzYL6eBMkRkH5Cra2X4732qeHIXKTZl0hO5jIUoSzhx1kdGiZCWqCM
d5Lf/P5gWI/tX7zK7t1Tsb76o3ImiC2MeKFwkGkbPOuC3cKoGX3T8U8vwiWkz3WfH2BpqJUi9MBa
8RtDsLqtVLOujq4X8CEiBmmL9c8d63Swc4h0A3lG+vwskkM4h2JjXtpqTDA+y91oJR+d4B6Uq8EF
8BS2aIGfFQPZBl5cqya2gl8vsuQsTPbkYF386AUWL33VOFgXdUZsvppoBZLkSHv6RCzCGf+1erQI
sdlqDxOUJG2i5RrUACwZ1NSCBZjbncLQRLZIqO/a2bgaYpgb6xPP7MuD9tKXOKpTalgUeqSlSEip
HQt87bGQ/aNQLYxUByaDihZ9wVuIgtP5d5rAodnRDxkTyBFMoGDbO2CDzi03YSy+mthJCAL/8+iZ
K9Ii2OzdRpYgrhK+cDt1I60mOb3YBhvJTxpemCdfj4WEm1ClXmvpN1V5iJocuqb/RPLydWfXT30L
4M9hnGBJI7VWB7jUDVubm8N+nvU3lxg+wE3hW/zZB5pYQ+S3q0x169kO0yCjoyabgnNOH1MdwbYZ
IngD+31pxGt/Y5t9qKqqYnlaho7hiHHGdBO9c/fMbk/Hd5yn2lfaL4YVasY93Oei8JW9bqS5lJOg
fjOIc+Xst+RgTc9wVfPAuL7NNosEKQoTsBHovNLdgvKNyy1BNqSTWGHk/CTdjmF2q9kGC6Jvb4NC
2wmO0e7EixOpcbdUnrolyve1fIzCpf62v3k0m+l9xZWXDeepSnrXzs1YapPAeuU/pffLGtGmDFUX
QeapH1GP+hiyynTl4KOekZX32G5b3CSa+Qw5XZlFdftC71xgnjG7VtXngXJrUgzkNWew2vWLLD8K
S1kCzkl7wRegL2uWY5iepLSwhOS24jfH3RTNVa4jWPQS/xvhDDEx5fPzFHkAf4jXaJZX4g09sOil
xfSK22ca0bRTKsalKG1knU5yM0hz+5JUFlvUwnRU60ZC2sDcf26PSPUuVWlgYPlL/grCP4MeF7ye
l5pVwVZFmSm1sALtSmdbVaSK/tZxDuqnKwPX4buAOtPQvOW8Sr9ICw3un9/d57A10kaidBAopod7
XYSFdgz0TKYebkevlGoylzd2NHoUndK11UH0ad+j6jRmIWJ95pllqZrZxgJ8wyrFc8RZvJEuk43p
QEjf5hbLa9Lai5pE+EZ84CstJdD22KILTa2Dj4uFywJd2a/AXQ08FLwp5gudowQNhrq/bfXQxDHe
9/TyGlE/imGfzqDnH0D3AvCmxxI+53bI4kk2j/ZoqDDIOhX3NIqvhHx+QwQvE2dMmfiDYfjdH3Up
MITieCyTLERkh8FCnMaON5LsweJI+N/H8XAl/WacibMq7kC+Gl6tAWMXheMHic8kg2NFssIQUmUe
rvkJ/WY9zgCUQ+PactOmMaR+e+spJOR35M3LPSp48tR8I81JJ2D//uOarYLYULrywqCR/nzFocXe
NczDF0UqstlGpMEejGcDVBmdxHVKWJWy8raWd1pDNOFWEpFfGLVuCVhWuO6czIj0XM4RL7GqzKlt
2J7BlzAgxFxE8FBy44//5YOw3avRtZDHmvjdTBGXHDeJjW/daBi7vw9+l/0oHRAHn+2R2imbOa38
tBVgD88vJtwymGBv7PS2JdYyI5Mo+tCQxSsXaq9AYSGEo6XBbvkGWGYdxGxY+lnwUWB7n5KdGpvQ
gBWzi9bkJqhOGDW7rcwfHUErePktoCjg6y/66Iad/J+uj3VjEG/FJEI2xYwGQyoDA2bySY7Zbj89
Fd/1rXy5W0so3clqHe6t+6pPz42Spb6vpkpvuYZj6tMun0rgs4DBFysqs/BEy19znRBk8QzBipww
m7XiCVHEor9f3+72mEtJRqkLGrNeWMaRPfq3P91CL01R+di127oWbXafDuR0Eydphwcya3L01yER
PjL72rFSX9+iKL9laF5g4pREaplv+klgFzI0b5FstkEykn3FoJXY1SqX63nrcJHj+0VBxIQ+S/t3
sM9hnb7FnKL2M6dmc8PvSToKdmkbuymv0+Tm30RsUG3uf13Nhiir1x765ZlkujDYUsbE9i6tdsm8
B2A3Mb8138aR6vj6tiSImEay60RKZWTnRwBT2Q5Mex75cmjJii1NK0vdDO2c5dRIoW742rne/r4h
UffqVciQ8bSNjRhI4k3xumu7zYRrXQbZ/yR4vzOSynqdMLgW7gAoB27DbbL7X+dTFf9N0PMh09bt
ft3Udnho6Pi8CybIAR7PukGv33NvgiPKjdrDfXTRmVFzX0cArYEWPgTEbrxiSYfqIzQV64d229GS
+WJE7QfXwnqVGIvF+hM1KloaK3DdnFM9+gqBaSaByikmciumHbEMceGERvgkk9aVpYF+P+uajH1o
e5Rz+JNaZxUJVPgUSdQILukyOctfV1OXMt7zZmL0vGABYQGjhsJ0LSHBMhRw6KefZq5AF49xlynC
+vyB2j1pqbK8xzbaRFevtPJBSErhDUhYVlChT6OkwjYvn84FZds0vV+VHp7Ff/XHxGyfb2bsFjRX
ZDzzlwYscxEhVkxaWHtaphXTH9CdO2TtoLQTjVykBmeH5AJd/WoslTidz+Gun+yJZdSGkezcmY/Z
0iYlrSjeUQ7a+YsKvkT+xuFL074KrVPQ6gmGhNyfKN6RudmGeJFn7w8KrH4PL29X0eWhpHiWtDC8
OIh+9IajyHdVuXeza90Hqbnk7fDi4L2deL1cBcDHr8oX8UTmXfwlkrWcW5AHexl3RwyLQJtNEEAU
7X3vNLBStuHMoaJVW24GjjRtfZWcfSHW3H11B4kR72GQVvfXoYphtKVSxM8jSSdLajeWs4luaVxd
N/kuqWF37/aHW+Ccx6o9ha9RrVrHZRZEP6teIZi76d0rqs6bBmIKUe8q48LHBXtP+ackp+OXiBOU
cN7IAyydsW8GFZUZF17fPzruuDi8360MqEAKOGfx2XoyfMcmybuBT6xrZ7dzmK2qoNxKwlJIESoM
mlUvaGOmmoA3pdTz49PPkGEaIO9duQLuKZak1fPInwQOt35bQtT9lfI/kVuk0/nQEPgkOnAsGKQm
6QJ9jtY4C/Eb0OexdLhO2eBwtnjjpBCVeZPnvubDmhQk5i5tNwxt9duHx7LwKP8fdpGx6IVo+CnI
Rzkr0lF81cA1RnHVMtlRLJA3hqFcZp3afTEE1ZAwJaa5lIy295+l3mLP1XI+ssgzg8J2Z1hVZcA5
2fMXkPHeEV4tjz+/SbkbczeF+KC/eHO7bZkxZiVIFgRlDMbzsydVb2b6S4QVO+Vb4Mi5qHD517Gu
hQc/hv08YJjdXUsFpH89N6BP8vuCfsvGoYJqikU4T0pyYfQC/BwcaKxUxZyuJP8QwyHP9F5wCW77
ebm3x0UG4mJ1c+mLGq185/pjmsEj1DcNbGmT7RC0fH9Xm2qqDZkDukf6pBNy3o0o2pbjTNmEIpkk
pKBasp+kRN7a8WITK3htZ1pJHsUF2XpUh6FGWMNxMmFJmC6zZMGTYFPeidZy7191yrfyP4uun/Zt
dJIzgghDxTywpW1T6hlMIJqT2wcbGBmoYTKQsAvDjeIs7TSw9CeaZCUorx9NvOZs6R2x4Vln6Pdf
e7z8gqlxS4J56QBTBcm438y/49k5dQ1q42+HKb0SmRNMKUAiWlfGPdVA261D+4aU9uGbo2yLGa3A
b1YtF9w34iaT0P+qCOu0V9wTOGUJlFyqWkRf4saUF2f3wc0bTPqZn2zvkTnq0pciPO6YXI+zdlsC
obn4q0ya5X9mzx+nhb+plVacOy7qcqgq/tLpvkl72hOmXJ9E8hnSkUfgPjNWV4Qv2BHnOwZ5Dtfc
KH5CGxO8qsFpfzuPLuF58mo8atGRvrNMDa4S9qLB1c6p0biEPwZ8mDRxCqIagBZsIDlQlg19aybM
ZEp9lCCtpubtVfTsEt4ALmJ1/hbt0+rQiRSpRdc/invlqibKSo7mdY/HF4SBOOuGb0Kb0bekxCvz
qoA/uKgYudFDLS0tHp+7EeSX2mwBBudULWD+udiBPwOB8Jd7G1vydoslZ7pwquXrmK35s4jxExDA
/38/smIEDYDD/uogY4cMZd1vZhek62uLv8Tgfk8FITu+cheYw8iAjFKobytNiLHb09CCGYqBno+1
+Jt9sNf6cSRiYnHleXiTDmyxIA5l+Yv+Q019w7tAb6stmftvkvtVlqgdWOpGyRpZUGmwkueGlk9W
a0KkOx4Elygslt5uDDmxDGVHD3sOTQmZHHQIpa1D7VnkgyflKnsaZVHdvMg7xVASkvzxLoB7RaZR
eV4ZdcYM134NC4n+sH1WmPtOk9PGZRsUZ0ENMjngidBz2PGMrgHYFrBEuBdxL0/upKBV6mpamm1F
W6tMZPgvNyWyobGK0xE8PhoFy4V7GKMD8p5DXmTGQag+lkXKU+7p+GWOyTwM/7kofJcv0W+CMdUW
BMmx7WHbnXS66opiW8jNYlTeBnXQZQlJ8cV0whoXvsNQtrijX49aiOOJfK9wlkjJ4sb5irlA1ebd
c18YQOg/dR95+KBz2vn9YE0Qle6n4T8A6OgzeNsA9A5/X6GEjAeAaSYq21EoXBsnNvJAopti8p30
l/AMasGF4eKZqA4zUR/uC1fXl0VqlMdlBYlJyjuSOrCqeTM3OP0BM2L2pqahm4RXkqwxOYomQUj0
gF4jUmKdZ0zSUE8koR9O6hd8sALiN/pAqDTwefjboXLbvomOOv07ZyPOd5KKv1TIiw8X67ao0D4/
ovMhHNSLf12PKmvgtHue7CfwT2PAu3+iKs+JrxKj3iyG/TFMcKJbZL70wY3VU0q9y0tk79zwEYI8
w9S9P0WshRRj36G82M5f40V0eI9yZJpsXTkNpn74BWNME+e+7mth+7obwH+0wvrH/QzDgz/mBtfq
W5ObUFB1ft4jy54MirhH6zLzYzLyYulE86eZXvKolMLkR+YC70sarCFlG7eZVWF1OY0V71pPKgvw
ZGBIj7f+CbfgoE8SYwPy/S5tb8HIDO9OAUvicBej6TrDDilXJuseuljONK06CbHXtrhW2w9sztrW
AN9iyV3FHzRgpkPIjlbmwrB8L5JpzJWRmzDe3EjPzWKAKofurtfrOMd9VIUzJjj50h7xeoL2hsdX
V9ZWOhBt21muJHhXSRrqcmaNpf+hl8C2u1ZcLnaAfNDqUTObjBqkW4cVY1x8FndI1RD6+dHm9FU3
BN+li4TsNVpk8q1VB++2ZmH99QWNJKmJ+h/Oo85JePbzhbJghmw2706W1pgQyZlM5Lqv5iEOax6k
n5BpQSD2LjyJPwWnGFwfjoV/Xn5+ew1Ase/xSfhH+HDZg84znEeZuiiRiFGden8COzbT0oWipsOT
U4wXrNObaBZm1xAj6fHqh7YYnhHHjSrp7TFnaymNTztDvt+6KVTSbwXZaRnurEH96WFIrjB6wHT1
2c3YH0J0sSwY7Wlu/v+MJJYDux/qGoTYyWRhLxrTBeUDu3KAM8UbsUsVKngR7xldzRMEkUVJTa7f
6BrxPzi3741MrkZiuTOQtCZbxgKl3XvZpeUcgcgsw/ghTiG4bq84Kl/hN6z1vV3mBIk3uE9CpfSP
VADKP+63+wax43hEK7Pi59A86lcUIp7oBpz2o+F1/nMkIiTU/x7UUnZkBYxoTuOrVb1jBgAPUhTD
hcYyYIEVHjXdWzday5w84VQDoJOzLp8DgXyL3WHqmywaFU9yx28UrLZ6RKuBAxnsnlTKOP9BMjdM
fkI+dS/hnFxLT5RAGsxqz1hTCcGbgB7MwCueSg1t/HvqsL8sr+8W04FCuLz78Jg2d4dsaa8fMFnv
ZNei6YbsCegkuqSvdLFcF/1TgYmw4aSVgujzco/ia3Tj6uU21Geme7lu0WRkO/+uBIP2juOfVhaD
3zX/eP8TA2W85VDEJtLbrf9KWL15pJhawr7BOY9ucPBJ+pTyqkyVKdRJ7K9PtdecWoUhH1nwtMV3
/910njPlndKHFuzCYYXl845mEkWs5HPmrMd7baAct4Yk9pBs+Js4ep87rTy671y1+HxayIkCxFvc
p5XhsvZLQt3vKZbQ4oIqVf1uAiOiZNs0bj1h8Wz5AsI2LTZ1jRgNHdJUZiyTOLgE0fly31qvbk+e
v96gx+Y5BAk4rxunX4tq6Zx/jX4oopPyG/LzmIAqhxLbFM4PlOQNG7UL/XVPeEJzodEZvwyjEjvD
Sll09v/LCaoUCVIvm/jcOGcgQlZtX6t/EuwHFg6ZESFryySizwzPVgW8eLH48uLj4V1zGhxyMF7d
OrlLw7s0a9sBbbuSXhf2DkhYqEAUG8oP/W7Yw/xZDfbl0IQ/9+Q5Q61WO08vuMo2i/i1eN6/L+GH
sWfXbfSld/t8vAKgo1MqmDTk0tzvESpUzcLGyuV66KLmk/K9uYif4A8IkGaKhjZIoyhQmxJ+hPp3
oOlXqeTM1ha1F71IT3T5OBkNnCC3A+teSw5bAJEWCUjK4QtIUXxmMnhmKFb0Vm6NBL1UK9vy4PMl
YxDnjEwuoDJbO4swCIGdfMfcM3af00cxtf3WrfCv1tSpQsqd9gLd/za/eP0SMj/pJvNTwULO6xdt
39mNoeGXrbmBxWMx8yZcgmVjCli4OQy/ekeTR9j/B2FXpkwnEKZWDmCP+07FaZPBAjYt39sw/N+5
P7ankT4RveiAIbwD/88/E5VhZWsw0FikvShAzky3gC4oHWnnuSfw0d8MhG/bS0uu85Qdpnfo0ATr
bfPqmK12Ssh6aaaz5X8fOoVmyvsXBc0wPxkcWoBsdLdSdzmkkxTU6ChVLA4KNX+AQY0c2vvdBWYf
gX198cTxcuzEmQS/AjhfuE6AkjwwoV8Ve0FmnFH+kZEenS1xjOTdfhoXJKkkmM2byykykdkFHsgT
kd8PTRTJNA42MJHCzzlu4eVB1eSCLEZZGMT6Hpm4CKfF28fOrq8Lfrm/zsw4VPhD0fa4e8pcI6Du
i3rZO6yRSYFsXb87vNLepFvoDurB5IyZkx00vbxE30uaYf1Wpy9YJ8UbnXMVZ0d3vH+rCDI0P/au
FHiu/Vz7APHXPsdDOI8bAIvq0RUYkYCIWr9pmlraSIGxmb0nn87YZCQeCOOEKs/aCOyE4zUgPBR3
go35sdduEBFDezbfOdqbzEqGVHiywON+fZaH6OeE/1Hpx3QrdoDXsRDhVdttqSE6eNRxRtZZjyXa
TkTYIiCzEqqUppGCrSN7fPcEX4DTaOwy5AXDqqlo2qbcGZEnnJ8BPDibx/3gSJQY2UjkMPcqvBKp
1/u4wm9B2KY0jCEhdpzsq2WUr/NFlFoUbpqM03GZXvlJ1Via0e6Nj11YLJAzQN75Qh2osOWznPKT
vB3zBda2xRuTIB28yvtXU8XNWc1kCAAow8Ov1PS6xbcAGw1GpM89k+C2a4Q3V4K0RFUS7ZZk4VdY
qSzTq1UK9/38h1ajgtnL2HBoQwF/kqG1qd17eH/URezbGZY7/UQDDFATrWASGE1JcbJ3K7gzEe7r
sYRYrYsplw4yVyuOUwEnLe4RjiIZaRmwNqXFjAFck3JrkliukpLOPYT9frYx9i2b2KplD9y9t6r0
HLQncStY4OrJKSbYzveO3YN6aLFouQdWVvqJz1Wvj/R1ywpaN42Ogo1CqFdpRG6StSUIVD2rIbF7
UzCzgo6OihYwcwJegTXj6vMtWOKHdvxlcgKg01k4xX6Qe5KJS6DN+Rmv9BEPPjt0XtC9b3Z7YhAd
B3Xqz+jCHKJMC42aSG4SafMS31c9uFyGzgtEGUpeHGQzsXlekF8AdmZfPDX+UT+/Egw0MFlQLS2B
VsfSXA1j4496xH1PkOm4BpG6vKXXzzxab+WXqIzaHxtKGW3RKinjJajxCi+bQ45MrDdIgceSmYIb
THhvf9dir8S/J4RPCTOGVt+R1R05sD/ZMnMldApMZxMFyO0BwKVBHVauUha99olXgipitpfLIlid
v2y0ZQ/9itpPsR76iq5kUqjHofKiLnyY9hxCiA4fdKdtejHaQJedVeO8veYn3rs7tkRU6i2gA39d
S26PgStLRzi/K4Y3JC0Wh0ATDNy8KWJOsnyJAB2VYAlOtnUJn9i46/wyMpbQNvncVsMQg/PaJLRt
xLWKvi9opIN4o5i9qhPjr1hoCZyKjlyqhnE5LA4Czy2ORGSmDtvNXtCHdcY0rgkIpSwIcSKtRDxl
+BJYSvyHa/V2Z9SEohLi2HoddsADKhn+Jz8Ueb9ZYzc+WvdjOZeKAY7H88myGVyX0eUtfWVC74EH
Smwy7h3yJfrJWkIMnsmn432VR/br5DhspRIh98Kt37qBILAoqZ7L1OGXrXPYHU1UHq4Z1QtEJM1y
+iojjGO5oaC9f3lP9bVGsCL9mnMYtC8W4O9dnRDNaEBAWEMYSNjd9xngbwbPGM0K2UvLv74gTCv/
Pmp6hON6TWH2hKrn/bGCpeFMdrEno4KGv9O2AcsWNYaRGOyLRe+znwKw7/hd7EeslXllW4muQVa/
D+KaBQPwbVA/z6m6OUmHeVItogdtC3IZMYCroqWXtVrIRLKAZKgFnkdemx4UoNzzDG3rU0C3LF14
zdEk/Et+YuEk1I8fj/j0yUrGkXjMc/cA4Vrkr6kS9y9LYN9hgB85Y9TCglGDYtJXbpK/Cx6ExML5
epSZhd7khhkY63pLmuc+uNCq2QmYN2HjkyEZc9WugYFreFQTAmJ+oQV/ZEXami8swny759cHszFB
AEbz7M4XMNo1S9j6tOLPdbBfPQZQX1lAZMY8PLmCRgs0BkifLwApgrJqJAN/WRwDtOdMu11exDny
R8mi9ocZYr/ZbZuI8VEe3Qh5eS9vpg24xpKoTzf6M5BXhPtZQBGUHgB/52boYuOmATSWEYQPGmd3
eyUXtqgUONzzD8GCiPoEGYMJHv74GjN/uVF3MEUWCo+9zIU/lODafoocDFu5v3fMZ2JVfJkcnBPn
ReOQdH3FHay6nDj+HfdMN8zcfO7M83bCdgSAKD7zuXABiKVJlyqjv0vCN7pVxqaT1vSLRIWltA5n
X5kJv1BcW1IBZHRMZnq7Dyc0XbxHHn5nDxYo3XSKF1SjS3V//AMed88tAqXqh0unZ8UEYcFIgq00
lkq0h00cJdHhBtfAWmLFUY+M6Y8l+PmX6oxu70SILx18MzpSVuWtsxoH0ETCrIMrm6irmKDgFNBt
d+oPvUfr5ArIRiBAQp7H2wOmViy/BE/mWQIhzEjtMxSw68AYYKb06Jl3IoYUFRodKf8YP8AtfYTN
9q74M+G3Ag7CqtNb6YXXIUYH3GuXx3kHcFuay+qzI/xXXYdNxavwVuKLD61mxkPTKzcN+bcGxaZX
kKKNgMjAn1arNw2JyU2KRSHDmxOFAFhxDuDatFiYezu6Bkqy5l3lqXEs46eR3UK/azNkgy9l9Q/2
r2QYyjiCm+dleMj8Q8wvArLpVTYz2AeCTtlDVmVSZ6qu465oewGZMRhMps1HWssdicwH54nVYUsX
Tm5RxPeauoddp5Qlu8mvjBlmBYLxSLIo6Z0kl0FXSEISMbzu1TVsPdD4MW7m84w7fV+jKPf2SOQM
H0GWd7ny0+HWTVy34Sinrr+4hLX+N0VBkQsOCq2/6Ma4i6OnL8HMI+SHdq4a8bCBPCTOgVibu6vg
zCkaN9yiVMEW3UVfV+QngHylJZOHFoHVE2WWijnsIX+VcQpo+PvMU9N/eHbn7WYan41tmawKY5tW
mHF0Gydj4dLx9/HAui4CflaXe0QBldkQ75y+KqC59O1aJPVUq93cxolNX0XcooEC9QW7X7BbXOSX
P5LxCTcbUkS9xZbfoWixBthHDM27yjllTYBvhtMKAj/3nhyGEo6Q3PNUZxgYKERPnOWyrFsS+PHf
0pqBp0gDGhl1MilHBvLoLOOQq6nzFL0PxIn+K7iDV0rVpkDfVvHGH1NzvM2/o1YOX/2qL+3vTXX2
Tm8IGhJoy3dmW8ai6cJSIqNBv6Ck4LciC6HEb/W3TTl9+sFDwShuS7oacDym++L78UnrmN2cxKXj
Q3oGyV92rHtZw5P8EJCT+jBnHKqJ0MrKnt6EZKU7MRnT/+IHO5I9NLzSC0YJZvqUr6vounLeLy3z
n5TWIqreIa3jG5AFDvyGjPAS9BNzF2V9Yxod6Ajad19WIqyOlsnqYai2i1OFnplJiL6rm3s+ZYyp
pU45kszfzt2I1rt4fJEG6x4jOfWRycGKN8ftclpiNGrDPDFLl4iaFu5skPPM4Rwib9XX5rvDWuqw
SmHgdGbUjaWJc2E5Wyle4UEkX7SjNyHsXuRGuzH+vv/9QQ2V4hmHBcfsUD5IC69vlLA4aKFPDNDF
0wygK6xjq6E4UMyWW/raOh5huT65TsSMU/rqKrfNp1rFsLB4dBA3Eb9xGjOXAfDTs+0zDFi/pCbs
mZtm4zni1im8g7LVmuXILqyulz+dwUnPmD+C8278ASfwfk06J+oflxDxCNTX3nGkpGoR4A4ViTLx
MXosJlFPLH1xXsjPtZk8xfuxPaDQXYd28Ai1/UdFOwHIKvl4ZNImWN5QIwmzctz6JRo9XnnUhauS
zAUC3ptpJe3KH0Kxo9/F8/UOc+UAFJdDsulUroHRrQgZtHaeuNHuqPrmJ0AEd886tCQwa68aGZW/
2kJJRRSkYCtkk1643VoNG1z01tMUSunIaHL3hymR4zcwWGuKCTyAcDPnuEg6h1YXvfXF7ZThnQUB
6H20WQaEi0I8yHPP4x2qfCm3HQ9gAWEBEIkgYjlmQ8wdIT88iEfSsVzcsoGO5FXJuoa3h+MMWtFL
lMBoPJgMxZR6pWH4ZLiNjvDFDj/eLCfrKxiwsnYxYgiyg9KfNfzN9ILeJ9I1RiOHwgKMMuZ6Ngmw
xQlSzR/MzmQmOH6u2Hw4kzGJygxpMChPqhzqJCJ5RUSGHfY876viTwCLhBFNKLLk3cnPmHkWk6Hf
AdB3L22cDDEDPSIrnfgzPATjN/a/cxXqa5g810nBVWotlxeC7lL9zmACnfS6vyVrtC8BjjuRUztc
tJmBOIw0pk7HNc0OttlImWM/iCVKJ4+bq48lMmEHqc/KvZbMpR76/tUG7MIRtvQ/L4TXUnDGq0ZY
7AXNbo4lAlu2wXCIigUYbYdImC7vVLfJZlKx9HYxHDHDflbXdZOA+FS67WFJCRGFpYYwrbhRDz2f
YlF5Pd/z4gHhE78RfBgHT+vPitdqr3FhqXgFcHvwr95QOZhZrMwpGTzm9Fw7GRS9JWrUzF9dsy53
+7fxCH+gKh2uMhOlH4wx39qOlvWp/iFnscqkfrcOnvXPw/vYezeTgeezFYcM3wAoL8/Hm5MWyqaD
glFJ8cPvfOHhoTruz35u8k9FuFoDsl7hLqKwYzGYSjr+JAX43LKtvaDBhWvVmsMczZGkY8fAdABc
S5sHcuasr+t42bm48IYHEnYaW4qYCyfDB5EZYHVNvyp3O21U3iggyW1dp4EOWHPZPxWTRznuS2Es
lNGv2I0Yycn8MPfUfp+XfRfwn/KR3FligiHdvx2++31yngPZWXR1klu7PwxDjLZGWy57RU8auBQE
GMcvZMuAQbPimehCxKW+ii/S75kjtY9yBeFBYxaGdTVwR1qJcAx5Yw9iJlSlIfjc5tXG5/pagET+
SIC3QE8h29PFsomB3HP0fO2BqDaFCm634lGjBeKKmZlylX7kwFck6SebFq0i6AUnQbudI3Ex63NO
Ch66zfymMRSog0b+gk0HYr4Tdfbu7wwkQIetCYCrVqtUqAED7IW43dyb5TMrpGd7A6pknmYuRwAb
fr95J37/lzT79YwW85Cv6hvEQcU6qyFOzgLFPiDy8CHfFxZ1/0oZkRAeJu3oZGGq/RG+Zqj7UDXr
QRAJALTe8p1420lRD+zFMREY2VdqMRA+2H3LUAsl0oqGQcy1njxY5RYLmGJ1eon0AFOUBL4qbdMA
qBaiILqS8D45bwDUzMB7T7lMHa5C2dXq5JDzYyK9xLJOvpC2JBR59EKT++XCGIH68gC6uhWWZtEu
RdZ1kfhJDHbuH+wNKEFiyj+EJlKLT2IuCbcCD+CVo1WDY66odKCCTlM5oC/7wmaFhWW9HyUI6XFE
KuCfcSkBmvHvL08GucGxAkx1eAUFu0FDX7RKW/aPzhzSYU1/um4FQfiTqC68mIJt4RFGP9GZ76tw
iLMSaw9NswQ66R7Dn3u76nk4lD6ykFNnVE50JTVWNlGb+hKOD7gNFkTYYGOpKP9TSVmUY2oUrTCU
2rlE7wTkQFIOK9rFKFfJpRttGavKede4gfjWJp+2I5uqKOfQwKu+ioyZpdiBjjF3ypxxkH3mmw/x
0IqnyN4f7PBLvn7+h7fidamWSpHd9xbWW8tb5mBTXUOHUR1AEIqqBQdY6+jlm5yGDl4mv731jtrb
5mWsMJM1WwHzcVTzjY4PB6WFSbXpGWRhtx1KIIQzF6x47DrtSaLnQsPezOWerzPPpUruFpru9w6y
FADt2pbkkHujkcE3PxBiiEtO5IwRgdC3Oj5oOoMPX45qlPe09YeEFDEHy+QtefP7gxDDhNcpn5FT
OuEoq9AzxR0YLWCdMSavkvHM4a4C1UiVOgRAsrJ3+WueP8DgEFT7I3tvyeQc7C2/GFlJQMQtXi6v
W1kb1WfDyUiXvgV0Bdkx83WLMv+MYJ8BMbHmKSis+VWRMdTfYXk3izwictGKLYisSN1mmr8cfb0N
DXOfPrBtYGUc8HnxeHB5DTsJ8JpwkkgMbVQ3GrqrWpXen7TOABm4lN4pcDtJWi6vN+RS4J/MgwVN
EktHquJRIrrTk1saMeOzuP7CjQ68jDRSEjQjHn78KEfDnCQfQ4Qc2+OhE2gHYjU5nitgsSOOLOio
qYT3FQk9w1e8NppkW3dGO1FENi/pMnCah5AepdyZmjjmS3Wtfmip+RcDavyMwLX+lguDlqZgurIV
F1Sdx/aJKOOhW6+kpMxYVMn3Dw0jpaGVhghP87x9ZOEyurbVvHDbs1xqQDYHP+l0WWZtCauDeUbW
hJ4gJI0f4UQ0FNxArClDYr3EcGbR+DJEegq+q0iG63ENwUK1sM44QArSBKNfotmzW1r+tYtC6ZDo
tsGBatzO0qjEx7q2DY3BKF/sSXyUT1tnJLd6htmOihm2qUmN11doH5vLATXaPtpkvpMsA8PMj/nr
6CEFfktr4EDt+0ABjqx4Ir4emDC56uOQ9Zwqx/vzpHoeiAF50gdxc/cZ9ahaqAVx06wcUk6SRBY2
bAcN76F6ybZS3WK1rNtqd6t6ma9fTgtA1erHNC4NipnlnMvYXOFzgiPWAcrnH0vuDTMVlFALtqzS
Md1j/TlqsEJy4S8BitLQjpS7DQNHTKV2eUBY+9F38Y8uhsp1RDnK+CtaQntu5Y9ymldoM7HUzY27
RJeKo4VWqRDnE99Tzc11RTswIu17cjg8tKMy7FJ0R7BnwsKwmb/72YXN/i94AXULxXtHjz3DWU6r
GMVjUMcRTFyBgtjnyxFHSZGcRb1JDPhDsUjGbo8kH5bznJ0cAmQryHkL9Vj+HH0uBdeGxQU4NslO
YxZbuQN0En2HQv/79qnpN+8DIPyNbePcSJbXpM1Q08uhVLkU5dbzDA8x+jyIjbC01VaM+PVv8ngr
qNMyNOOuyl/80Y1CKini00Rm0lcAZA1EsNZe9FQsSi4QjxEFu5VfRyOAUWBki2T392J+uaPtgTim
w/9JEaAmA/ZS6AdW1eD1+omOBTSr2IaaPkHnZmGWZh0xwp5bbddxpQ2sJoJPkPueKpDhPxnnlhKo
C0WGWvMi6b8//f4p/IuJurLaX3vItYnmIuOedc4IMKX3h63r0ay9p3pe4NqJXBNoy3L5ctHt5F6b
NGFN0BXmYNIn8lKO2aRsJG9JfHCqzYE3ji9sCvtWOx3D9BeWBvCL4vrdNO1kVx3QQZmhkyIYIIky
pn1mkqUbOt/059MXrZDmwPtVoqYpSwRA0JOHG9QMVVyk4VqVn4TtLWOI8iH5tmWtHJ5ecIj4hG2J
/QoJ0uuOX9MbFwPVkabwk0yQC7EZ1KChM8dnvlwooPmrU0YUhel1jzWlpBpIQCagqyLkCdpuZ8rV
dk1SIB97ag+qqMWXnmTOAZlKyRNHjoaH2n92pdHvLZQsyuhc1UhaOvJXeh1/kEIhINusQeL3pKSQ
p9xNFn13Pcc8LNfLTs/G+RtKqzsnfT054C5yDhwrzLH7ZfxcHT8UK6GiuCJDWF9hXsZf0kdj5TII
LYja+118LX5d93Uez2SN7jfuPfwP8tmf9Pg7dI7N8l7a6Wnrpa0kSPPSaqlyosWAs6g4aX9sqRlh
KUqOFEMPMQUahhco+cvLig+JKKye0VFKYNd+8fWJpALLW+wkZhFckO067vEUBxkUxgTXye+WjKv0
o1rz1bS0xQd/aY2oqsMuXeIc5LXh+qBEnlK/54was2U/erPMWoy8NtgANed/kFFaioXKwwBi7NTv
GanHPL0Pc6D19Lrv5x9aKbJ4XXImErBS4tS7bfveFrerZ4JaepUheG7tfhF3afe25Zk4xTo6Gve4
aH1HgEanChWpE7kYXApywgLJA8I0M6TDEvwn+nCY3u9m0/w4P9i/nefOOApmFGEtiO/FjhM6rlny
nvC24DbAIsIFXtY6n7Fqso40hs34SN0KTNHXon2/+r4xzMjLAoI1UxSQ3y7zmqPcWIxJhLZHRLP8
bh0kn7wIfjqnbwmBZ7uoymaRHEgGeUvJu3rYaxyY3KxMFzWqtYBpkdEryYiEWB3SbQgie+6SKZNN
CdU/iVPcXtEobP02eP0ZhvKFGG01vIEN1rSZ8BN+1dBo/Kt6V8dR4Zl38JZlWD+9LznZgyJ1L7kR
dLtZVptb8y0rPVt2YR40GJ3CDPQ8H8Q/2/f88MEmGy929vNba5ZeGzNLOpuLntcadYmUZx7QKw5T
nR9H+tr8UuOMj2qNihgIc11x70AEGqMO0AYxjaaiTOhvRWAtU6/ZTdDXWr0/kbYlHKvz/a/Uwrnr
AdAMMIAKBc2Mqabi0ZVYpqCEuyC3pq8HIWET5y0/xsIt/vbMLJ6WbLeELR7VKicW6XD4ZIAljgHF
3I9qHQbp3lM6AQCL/JfdaifMZm+k3ThnNpgOtCa3UkMlXoHndW0aUN6EmRupGCIDV1Bo+SQPAsHk
D22/Sk4ngreSKAQ1j1OnZaRUoOrJpYnLdfRdzzc9s0iVN93xZ2IZ7zG/D1x9mhA6VhUNzIRnuvJh
USHKnBDiKoobzo9zQxSUWH2AHJTVspAk6OEs4ajybyKqcpDMPmBava7yVEysx37XtKDYcsFUpbOO
pXQ5GULt0TeBlHpDLDe0J0cvHte5xPDbO/63pjpW3i2rNjhMZOP7lJ3pVVuaeckvgMdLuu00NAMT
7PIZgcA8+v1ECjYrqocn3zb5Y9FGx7xNrofmopv9vRbM68g0OLuylhKz0tCYm9RZ+MwvPdaOTJxP
YsPaFwAsImhg4YBz6+iJGftA0X1+JISfAkvwf/q7KSx5x23slbtDbtUfHUzC/w8T/Hj60+JMdffY
bmHFZEybE5ZkXG9NecdF1cznQT0XSHQCAEoNfDP1KDQzEi1vwhv781JyMn+LAv+cSGJ16oUJZvUp
frX9lUIG+WzZUmqKGZ2gqtj0uVvcGJeEYgRRNsq5pB8zVY8G6/OD4V3FunNttkZi1C5pPXzKao92
dPAykZ4+crK90dIeigyTBmWF2CrnAvttjO/bV48LOjJl8YiPZeXdC+ImydKW1m42TggJq3EXuN6c
Uf2WTWDSrHbsshUgZzqeBE3Nttrh8U2Y0vMQJG1+S+nrj2L3ughUkrUPPYf3hl4buAunLI0BImx7
xTkQ0QWrFTyWZ5hsF3whbozQdAaQMwcTwxIEffJoc+eU3OeontlaoqrLXp4FWXi/dANPEpC+90Y4
DG2IXf7LnvWew9vwwK9YKBn0O3jYvPMxOUEhkX6tJrwMC/uuMqyeo0x55gKf6jB0qBlGWB2ntdpB
sgdPoHvRJgd/0/f4ojpQSzM2Ern6FlQmfs6CBQIzDsdjMUQCDbTkSZy2GYOnT0muBBUUSCCUgTBs
1pwyIlUHGCHxJ9OB1YvE1nv/rINWPOSG7Kg+wjqy1F651FaeEJL7z0rq3f7QO1l9V9jokZhKOrdf
1nNQvaddP2st78chn5deyYDRrTExBMrT2jtXwlyQ7UZlqJHGnUnoGXg0lGhXMQxCmyvrjfquu872
JW42NTNsH+Dddb5F/cJoxbWp6DiDymE2XEoEGlh4IbbMuFvirwcc/CtUy8AVVvZdvVcRQWhH6izw
o58W6VlRiTN+jIRJ6CpPzWyo5LgoenSCOFg/5FOOJLx+HCgRTXNlHhwtPW1I05UClls6JSiRPd6j
gmppHOW6GK4cOJL5C+jOLXqbHsmfDMyzdEIGbW2zdF8n1luVNPcG8A0dsUCW2Zj+ZBI5eCADHSaL
CGcw6ZXvzynGAWFtVm6YF/v+sNS1oA/Ec3EFIu2moFocQEMaChg0wpiIBBQRqJdBX+7abw2fgKzT
MTh93Z/shNjgDj8m28gqwTqnbvBTKmDVhLwd4/3MW6W71aprfQ5x31EZFClbvBk58ot9RkWxlcxK
bxvcT9Sx7i1tM6dEO+zBZF75mfHwVkguKNi74EkdfFfb0mw8DWIcmrAosrXGGjO0RM4Fg56GVOjl
/VISCyjyGv1UKJ3ATCICBliP7NkSzMrKPdDJFpg7dLGrxHIzEkHA0sgczrOWbUlijl2n84ThZoiP
/Dz8sR/gOrYTcfN9J77+9VKOfIqO3ZmGmxSGVI+E3pKoMH2K5JA3ewFJiKBdNcEUPUS9zQ9eHvB5
uW/h29PJxifUf8La6u7VjbX1hb1tLYwc8XPTkhodMgbYlvHh7KPvQVYkifOOUiq2f4Iwo5JuqjAw
nGfkxFWSj8xEn8dmNCpTFk1aD5jQjWYHttxY6qcAgO2kG9Ihx2YdX+SgpYkIG4HNPzpF7/JoDtWe
L3njiMFJvi8vjmIuCQGqfRx1fgd55712QSmE7q48I+SdSI/JASEtSh0oh4J73rxKI/dXqfsZOkxB
O/CHFgr4MKG9KlKvH13c0gDV9Tr+r2wub/Xg4doZjjmLPWqp6OKI5XRccyKhYqh9usDzYdL3fKPJ
dCEt73Uv6P9mRzEaiFb3n5DWZ1Fdx+hnVXq3PiHs0FD1Z/f3HezF+4Pcl/is5M4N1fAhyEUmTG/h
TPZF1wBM9SnrIG7csiu/0QL5ZSZV92qtEMJVODyYUYQ7AtevX2fKu914U3A/XKlTEs7E+v6IXvDY
Ii8aU6aWAhrG+Q1fSLOuHuXwhamgWdwldG0biiEZzrY1jPfk4v0aZWZYLg0tG/gioB3gTB0rATRI
eWDx3mhHRQXuY/5IodLUjyeSSAwCA9O4g0xUsRe+cqC0ggy4fIRJgE1rJ4cQkdJWlhcxcokaOZm6
oL9jr0ZDJ3eCT4v5EIZ5IwYGJnaZOumWDsRH5IdztzbxGZlcj01sJwZjdX9LCTxftSwJHOdwPu1K
+6KAe5jqF+X/zDytA0NYgg57q9+b9YtxogtG+fqPmUsnbdA83G9ur6ubQirJJeala5Qg4LTIYKht
DQfJB49URjulrD/D5B1bbTTeGlrGRHsdZTTn3F1H1nz2oEC1qdjwAFkTYh91oR1HIMDYaKHWKw2+
wGmqJDFqEqLAetInVWvY9ze5+XEpoR5aIV9NzoD6XVGIxCFAyQD5tXS+v7FHZfHijyfl/lM5oEVj
OZOjsgVIRrDnFXF81RWrQy0nmdSYJinNs9VbBOX9lWRBuLnn4RVeJpW1LIb3WJz3j655GIte/4Z6
1jUWdqJvBBzf9npAHQ8eCqnw/G8NNyucSyegidPdV9cS34+urHFFlSDC2FGv0tkjbqm3D34M/fbJ
5iKxy5hvatjongrkn7nPtLY1PanCzaLln6hLyW6eR8uWURL1KgATeolOom1IxCZp0f92o5ckHI71
ym9Cgses7mB+RKRJazFWnFYmvnWaJaANA+lH5IpawQVSSD0LYrSj4gS6Bf0A9MoaTADiiZiCCxQd
9156r0lNHkQFNXJ97MlX2ZCEHh+29W17ZOGTdaHV4eUmeeUwMUfxgyhuJI1pKhMcjyBfkB1F8i13
PSZXw6us1D1y8PLw5FXYT5OqQoB9LPp3vsD9bZ+CDKw0MgL94DtoQ1f5xEQLIgsHePfnngOvKD96
QKwMOMAmfz84PahBp9iE7flCfwQtROBaAsqcM0MhSxXj+HZQ8Dc4OtaPdpf/jPQSngK11dKioROH
S41P2hfl+Mx1r48GL8G7pu6ljU5a940DC1ulB5hF10ZwtOZpVwYI5CQpZ1B4V9UDfU4BiU1Qkjqe
2l1D3cZ8ChllyO+lq6gwbxV8Nwu1p0JiQTJ4As4paTFl2e4KUJ5bbz/rCdWWj3raSVGddUwYWbjo
NSaE3cCrE1vriUaz4u+Ggpjdh5Tmkd84neIf3eM17lYORoJ7sjxQNnfwz+xfsJy1NHdUgx82j+CC
laoAOQGZU3PzLIrZJJ6YWYp50mowuttGR8l2x8CStDtr5lhy6ldPpnZDtp9RX9KMUYF5a4Z2Yfb6
lBA39mMI234LtH51OrXTycuYbaRzXY4Yn+XF5niGQnvxZZrSySnA8onsiN+rkSwzYi+FzRKyhsng
gu5vTmbYkItYDdQ8EWJ48WVA/tuC4xnaFY4k2HaX4nkaHqBsU/DmmnIzAOM2aj1ZohOeXmX3YH1P
lJFyJQgxGmQC0RUaiR8s6OovBsrwqROCiocr3YdFq9TvqWfpzGBqHIwB5kP7zLIzeD2Wtp9zmyRF
9Sm6LiMS0G9wqFTG3nOHC7UVsE18FFGvU8mMHiG29vRVNj/w4vRks4LXAkMbmzqZMlLJV8xC1rBf
nGoqQtFCiPUMzDNuwOWG7bcqH4oEO88H/l1PbTWp03MZILTTxirqtMPsSBFRacnbwTuRxJlQM4ig
ecLtaU5djGB/PZiGA6Y6tLVQdO3gXc5F5dtdHB7u8Ij0Gx6XaJs8zh7ip5QJogFfwOiA9N5fLfBH
eRzj/UO3l6uTA4msLXAZgBjpVYEMzWJSWVemz7+BvsFzOzl/C9Dg5slx2hnHeWspeDOicbXElhFa
FRDSp17g5EHSA7D972mrDcsyE7BUU3hDtMH2aN3H/EKqw3QCyDRcYf502evs5EC4/hgUf3E03V/8
diYpTcZwk7rbo1feyg3RF9mU02v4MBExoINLU+Z2CufUSH4cwaJn5Vd2LJnQOtwoxjNXj/P+SzjV
zSubFVd3LBh7pDE29vlht/hNQO1KcvA8xmoV/72WoWiIXUUq3qXwdjj7Uxlzet/p/ZQydiulNu/S
MMb2mnIzWmNVhCVmNdtslIySHghP3+5Z3LImrbSid/6VRBspc8hGyDBFKk5sFxtzScuoTGS9nw3T
0SISmQq/vwO9ytaHocimLmJZI/QuIYOFm3s51TTxnhJXHW20ybpr7vBeitYjZCrlLFtg6+9kw+vP
OMyyMUFoninQ+ay68tlu0nGXWNg5pTivNIdbLY77pRf7s0eB/7ndAtVH38DCoBW+Vu3OWp9fo3NP
EXRfzXiZ4tuoiNpm0TjijpIwM4TVkE03TbjGSAW6c9iEGsyNcNUpFAVzC2d353TntjL+8H5j7xav
9q3PogzKy8HJNcmnc07wQbiiTrfm8AWO6musIq0IWCtXHPmgeKedDoio/f/0QOTTbkY5j+qY8LPy
eoKkdzSBWTQsIyZ5Ahe/cKGOATyWEzu8KBl0EyMB0r/pTS9W0VL35HcvTSHqNo47Bi0BSrXXpoKh
b5q6qCLijeTuKFZ31qGnWTniWkqVMWlbZf2ZIVjYnsNExVGpOmN6wruVg+1GZTegqcWyHwgv+kIx
wYljhu9Piu3k0CGo9O5KHSgo4xtj6geUnnLz/N0j5w8ex8TBnd0Zb+HVEtKLD753Ych9iyvCacBP
biLRR0Sfr80C+2KDSoEYoxBBTHck1NPjGgnHZyDTp0KlWtrqKNN1U4hz24iapxkOYJGlCyWIcHft
rKjWwscRMVWJE0xyv2C4ma0JbeBswL8sfbOUhhewg/CBiA4hhM23WQEmRBqR7SqoMiJSPI6Z6oVL
m/ZkIWoYhSG0oVwoldSQFfh45jBl8MNz/Be3xSs9U8AOn23vWw40XIuwOi/lC+YvKdRaKNMTWO2h
+t30a+YMNsx4wK8ex/3gMpCRjaZNpHejqiPXIQPDY9Gg8efmPztC3G+dISD/S3ZVNkqEVyeXgW8v
/+Br1KReC7yAJwxiazHoT04yBKWZHMtbI6nIISZlvtQ8P9XdjwW8/xYygekZXFFMggIIAz3HgxQM
vrjCbmJiU+u+SZgqIBmmONblGBnSqcjyZ/suVzUZahMOtFs8xG7eoVjfj1dsbws/b2W8b97ACJQ0
i2gao79N5IFKoaA7RCMhTd+B71wd3C/xa3G7WTtU4Eu+eN7rIlcTvU7/NZWzYi4UGU3URr179jA5
7/4a9+XsAjpY5bosjFR1AL5eXAj9jKz0+eYkpaJL75Lfwv1/qPX2mNrp08Lm99OkkIq8jdm9py2x
1q9qPNaHJH3TLqKjuejLM1gqKvX+GZiasp2R5fmdPV1ySlFDtoHioup+nefJNf8mrqgnOvMTJdIt
zTGLqhKBHWWYCKLMfLQ/OxvpasUKwbW7+CWuWxyAB5m81Aaljce4zxszNgKABfdETBQCVGFkaWVs
zyfZVCjq+h4uUgbPaxvqIbjQERMUAbq1ZW1aHd3zsxzmWnc0D3N+m6kVx4gKvY491gI1ph7xEsUZ
qDeq37R9YQIQGl225iXSgqeHVsw0BAZRLmfQaUxmlU7zODNq9O9PrjOyX6fkl3XWPTGBuTLCmOpr
Pv/icGQ+RFzm/3b5XQpnjII7mgtP/5F8AhawW0AO4/UHkakasOWuhNSaSGUMeeoGxAgPQgvlH+fk
180btRE0KhIOrkiP4qpmpeS7ceDhMbD1oY9q/veRsoOf9GITCCeJIpxgQK6yxfh5IhGB4x2X2XJM
kMskWglodoIrmEtj4+db4TKCcBnASxhLXM/rj3UWkrqNi4PLDHE1qStxWAqg4yJhXN4bJ9wOq3Bs
5frMQNUkAKaPJCdOMJ1Ce3Q8dBFDenn5+G1qL6JBtnCs4B5t0bnLGAqYtNa5nai8GyIH4RIcetaU
TDyw2DX0xt8AQTLDh6qpXI4wOZxW0NgfMqVBJtctPUtB45frTTp+ZrRiLGvgUwo59Z7Z6Zcf81o0
zuqQ+FI4UQS3g6my0MSjDiPKhStMqGmDzC7Hc4C4jwy0y5Jh8N15AzUQc6PNBi+pe85M+DF94vJJ
HCZiiJEDX2brH1kVyachBT7XPR2RtyJq889PMxNCbDIYQMmjxeGw42G0hw0lXeJbpKFj2nLs0K2O
iyCQAXrVN2LdWxYCsfI3nM4Fngpp8JGStbJjNhcWnuxtAOtKIkVZc4p4oHsOwJESQZUHwOq9Ne0z
6GdwvYaDtj7pV51S/+LJKRHHlOiOmmWITIstLZCJOp3y4iu1fzu1hvck+wua9XQg/heLcA4Z40SK
SqRju3Cw/Gb8+kywuNCNMD+5v+kFjIG3dMpU11gYMTr3MRoXEUAX6PSHkJ3lBBLcL0OMMAV7W0J8
q4DHc88yrg2viOs1CbIUn+EfzA83DYcFkS2vq9lSEhLIQQIPvBvkD5fJkdtBz4xlXal+0zvTU+OS
7XVRacT4leDaA38iEZy6a9lPZP3kUKWGhSIgqgDxfAR6QRtw3CqpM5+G71wBHawJZqJwlbllppBR
B/q1NXY92d0wKIqVjQXGagR2Piyxwbrp4ML65UYr4w6mjTdZCH1qvGqoUgHsdHqhYt6Ld4zzHE2F
Ta+EU4Cu9x2ts0Mby3EDKvkxE1NReE+MwD2c5++rxYw1+aueqsN3YQDmYuCZyecUmNnq4ahYh4x/
C1BeTqGprYe51xDklkREbJf9Gb/vvBnB4mJZVG50QlyMcChEDsMlhpgF6H5iD4D/Dq3sXRWTAz6T
xZQbWbm1XKf1M/PI5WMHV3hKs6ZFBjgeEaFsR1ARwW8iVGLwZA1FrGfGl+DxCkLfimJarWXkkeuI
V3ZrFnuMO0dGeHtH629J+7n+537dcaaLSH/3g42lAZGoI99TwRO9Nl7gJ8TkHNCnvRp4UvLP2CZ9
yADKK+Up5i6ACin9j6ZXhPTegzwBfWzVAdLu5r93MrwaZaAHETPMq9vwg3f7jf2zgVH3Bs2qOT68
z41ltEpteB6NteeDFyqKVFXdsQ24FhnE5xQscj8z1d94no06yYEHL24j/LTkC3kLqTNeAymu5nHU
Nfbwzs3WvgztaXdiTnrmvJUVSuYmLzv/17fAUcnFCj3ZnGbX1pdJym/NarBgMyqeSeifZpFhpcA3
xCsq0Q+x3pHyLJFeU6Q8YeOY4BJpLssHdnX212oqjw1HtXz+EEwkHqkFEbaWnwjxKMV8NfpTAHf+
XIjQfmHk0duGJP4QSmd3vZdBmfF/cnb2Xgf6J431dIq1AY61P+A9VxG9VKxX6UVEV3j5BUSeoe4t
06klejQPP9N0rSYH2H92G6dlIrNZFPXuAAGHMy3ptffiULdbZC75zDuTx8BsHGryh2H2alsXr1Nv
6YlIPu1DUP7o3R4kzqGEldslb9BNlLF004+rGqHZaAjGr06YVwCnaiF+SeNJE5bXR1Prphl1h2yh
fXsBJyUP59GZCH2QHREDs2jiNHeylhq0lIbof4ROzf/zeGqBSNPYMpTkB4aCT7bjeboew6Z1QUBy
0bRQwIGryFW4/0zLVVB2l8BqBtjf4/b0q5LiN0fLlVlxGjFHNmza34Kf+vY+dB5QkL5qdUBhNCSf
wiga3QlpH+PelFiSy2Pvcs9BJlJN4LDQSDm8SeqGD3s92GyNbzeoS1yn0e0zszQ1ieWAn9nAnSGq
6oy6lSVz+CkQ1zp3FX0Oqtfw9NTKlUwx/fGhKWeXp7auj36ulygwimVaXnHJj/vr6ulAUtpJNtyO
KpjZ2RGI4kqOL5vUc1mmdzHqPHm0GRwoaNyR0CaTUPV9hI7E6nu5X10V2OO+0s9yEHQCzoH9pBqE
hwPibaD79fo4YenLvnAMgzeP2PTnMiZLGGRWAhTYw+KY8/ACMBZHypjbMgQStZUX4nIDJ3oyJ6C/
jsEGVRlJUSEHv5SQT6LdVp8fJK+qMO6cWjwlRKXNvuuwrIM8T/GKyrssujx0HcD/dSkR5b4nEUy/
olaYA4CXBjn+3MJJ24ohx9/GEkyZ5MLqF+OMhkfjGNMXVvmvcw/uKKfsgPzh9MpZvJC+EfsIc+DK
wN5wR1SqhWX/Mgg5F/CcQzw7yp8lWxn22YWGzXzwiSFvGRjCzPv1QXeJv7TClVDEWwCQETC5/jkG
CjyY9hdKpSw8hXyWdMSPQ6q4dCfLwZu/B3eayowDuKBjX+GFdqicge93qz10nGi+cAtnCEbEKcwt
ZB8oJ4wYWzFynMMbaaMnaxgQddY8UChhApjhXs7pLgRW4/iyMi+VmGx1zH96sIfag9ADuf/R2KNp
e+t908RgHGW7XpMligP6aRLGHRTbX7XkWskdyPkovia/MtFpeF6Pm3w6dFcJnTsbPluJvkI2oR8c
1BrrLk0+ZLu93jD0COPm7lcl97u99wOazZt6JUXl9ywrZ/909JERAPRpHVr/VfsLwR4ALGTiDxbF
egEy5nup/nHTLfYCn+CTIhvU5J5KIzs7VY/G2+U0KRBrZaGrLw+wr2M5DFMU2iAaEhiAH6JxUXGY
6PvKCsZpGPjfPptWT9zRmeiSQ6YsSGxpfrAl4pvIoKf1bV3DjFnoZypkFZPJiysS9TYFiIFt+QdM
4999V/omzL9CH1dNgr0uxxkO7agl8WRJs04h/SyPib/WKCyHl6rgNRu7S3HjuwkPnolFV3tIw8ai
q0Qu29AOogBYUTH/iVQ3/kEFJcEfcTmoem8p39PqOAnBwzP3jzGowPxHZuvQkiGjRhoEssL9uJxZ
33BPsVxZ0LZUuU6u2QzF/lSx6S98Td/0UM/7iKyQi3jS4upIefzxpSxwNQ07iHgvfjA2Wa28jXAG
vU/eT5CReFfntUE4aQclxcGHpNa2dPfXkvvfROOqTSiOOLgyb76yM0hU5O5o9i530I+4vN19qmSa
nZESOCudEA4vVSfdYBVJzMXa1wG3IifUImC5rwhhil95xz+SmslHYUr6/m83mxi8WZ8ifHy3KYTJ
P24qDWjnyp+WDY93sYwFsHJWKMEbGJXHMg3YVBVyZjj4rbz63FRAq+GA+0A/LBEuovc8plm3hO1a
df+S+U5MSio2r/SuVxKiJu0fVU9hJtzTv+iLzO7U0r2dyrzZXJAF/BOi+64/e32pSpphg34Mh7ch
AygWViKUJYvO6Wn6nIvL4W2c4RRnCdzP8Q2cQBflvldN9XCCCfg4BCwaTCU+U6AN94Pjl0npIJ+0
MSIgv7zedtfvq2eKWYjxBlXKVBzHBqoO73N1nSXoMze8QsMLtR+spGScpwhfl2AWrKMiDevmQMtF
KAWAIkP06OMnDIiBrNUBSv4C/vT2UZJo5J96Dz5z9S3E1yMht3Mt4jXmu7kY3m+5lkRUzL5IvXeE
66tto+SNCYCkwAS9tOUO3M5JwAlkhp/MWr4TfffD7xVPGm8yfEyWBZHOvNxjEaqGIOtnxPMeyXHM
ClUuZY0oAfyXL1eqeOK3qgZx0clv4aHeJohlp9LoYqHtw+2AgILpO8/4JPtxb3N2cYfP2xQr9moG
lw2ipU8WnndUVPFxV09tBgQz6f7OJdpr7oNPmWJdXXeb9konuza2I2Ai6hQaRzEWn+Fmyh1gEaRm
IeHTSzd3LR8HTpzFxvwEUdY1p08Vv2x5Fis3XpZL2ibxuEEq8EEs720NUaQS/Fx3u3UiYHoZXcIa
vZGb2/8QrIiOl0M8Z2cS+OrpdZ0T1t6GL91Ps1PLcjZUKJqmzvj14tDC4zTjrVaySWdt1Z5OF0m2
0x7Z0etw+MrOBh//9tU9bEI7ExdYvV4Gl+vnVpse4nolTWKPxp36WiF23MhTWbAWVzwwrvHh7NGh
fTyWLvj3LTtV8UOciuoOimum2A/afrpWwEN0q3wwcn4gxGF4LT0X3+TVX/6oK74ZLBQXW2YnCwzc
y4G8+BctHkkC1/Z8GeUb3n9I/Mi9JVIgzUyZvLbOiZ9V0EG5cec/lg3Obqs051fuRKzmhzVY1NXl
hymOhaIix1SDALVRu6/yqeoEzn0fQ9kC7/Kqo2H7ys6txYWuVmwl15K+5obiUgpnIsAB88sF704d
CYgoQzgJTJvAkRJfD097ArtzTHU1dkjyhmyTWNl2zVGFb7Zl14/BocNPIb/RbJzXM3CjRi2yLrPV
m50dpcFjOTxwq+Dee5tHVAEiXDuX2nkxhWHoxcKpLWmGIWqArfmw1K+zFKd4PDq81K7zbFTQREtg
2xb1y5O4+AJKFxELjc7d+4vmRG0RsNwIiehWQVU03t+23leCeO/ZOFKDWzb831XH/a45HNpQHRmE
aRgAqvdZjBfWtPYCRS04vzY2apVFyA0nCAjPDF3XcXV0EehzT1HX3ORwhuGxk0a1brRNAklJDGVo
HcaDZX3Bz56Cklopb8CohxnzxBGUINMK87bm/iOdOfGLx/N6SAt1MoGQ2ywXoakVheLhNNVHFUqv
USxQQopSIIWwooJvyn+5ieQca2jcMZ8HrcRQYNamhahsqeC6dl/9ee1VLuLwil5km6tVQm8Dh8WJ
ngw1mBEyqVANAl/200Qhf1lJvU3Cc1/mJ94mPH9wgucI6xXcQfblDZXerjs0RQHX4WbWHc8hkUlw
o7tn/9gyI+jrLHLJ4H4qQhwsNRbJWnPJDR2IBqURIvIfJBRQcZglkObUKBI/yTSExcAYiAvsZsXx
0IINYdbmqz5TNnFFykTEs3hOwJLWZ3bOzeY0R0A9nrLhNekolOaNWQ/7Rr35tsr27y1+HIZVxSyN
hp1emCdpAy3A5KyEJWFEI5QmpZAA+STqTMZJuQEcD19pvtJ4SjeNMPY3l3ZN4Y6UXcwz15QiHGwZ
/S47OLFjb+8YVayQLYVkjknOwnY6/IeG+EemCrhMOqLv1gjciHRoAuDHD3OMDG6zFHJuXptrx3W9
guc2hdjrjn9uycncm7F8fj9s3P2jGEqk2Ge1yqgmsxr9q6BcmRFC0czf/fjk4e07Wq0xsTUsS3kf
+R6w5jSFmebnI1o5Tzh/vkXR71djCIevjOs28whBsjnk2j3ts4Uwn6yIHln7ES8T7x1EX0ughhx2
M+knRf48GnISBR6SyteGn9Efu02mF8BHdwtAS/Q5VlPzwshaA3zs97CfGqc36gQqQQ6shSz6Th/B
kFtDbw9oUZIe6Plh3p87F1vDehxhmN6hIcgFR/RuPAicZikx2ufjMJCLTteR/4JOkhf/wVHMy4Me
eAhfThk8E2nmE8uYJC+QQbqA/5uxC3Kv9nN8HSB5rqMskrKBG3ru/tQx1a1T8IyEUEkGSo1H1Wvm
S8hWgK+2zlLa6bMv8dNm0By63B+0YrkkEqo9/XzGIzUeS4j+Lr2bCPrWjuI0lmEdijorUsGZroXU
XXHA+GIM4/zF0vQzKwgoTZELbiMoJPJhXQYaODZ52NZqVICZAJTAbj/x4ldq1WT3ZYu24GL9UOze
ex3qK+wH4rNwAjxjNGHVkwecwD7QXB+L5JtZGyx9Aic6Ittt9XRCOWTTMylVtOk4n46/HWDKKMU4
aTUplG0/KsiYFz8fjLczSYy+ZYOIMMHnOdgMfUrYKzKtaIuLAT4ikT4sNrw1JHZljcBM8O0VMWSY
pC9XoHIO1BTe0uWw4hqEL8ASC2JzHKstOcUZ/u+ipttR5b0LxJleQ7Pb17RrG5M9RK6D/WdQWz13
CDdElj7YsJn59Co47sY/yurnhvaL6FdYk9YNX75+litiDYXKt3aI6ViiOUGejY07h46wXRM+3nnZ
PME+dNTY3lw1bOBmCTmYVLPl/PNbW7+Ye1Y3TM0FOAPYFJDjsxFHFQHJrYPTnLTAwx2C9muTHys5
N6EXwrx76SKr5Y0NE0NnS8mt2BX070/kizbtRVtexV9uUh9lWSGObfuB0ixRdl53US6BtKFsZTr0
YFvgKSKXbrMRjBA0Q7WRngRbQHKH5GMqHNeEyoNfR7n1xCiVUGtRBwY3MBh1cu/JffSoGxARYQxt
/+S+Nxl+Q+E2n8M2+zDJMVb0EU3yRUhOgj/15ObIgRb0u7jHDaZkeJNgmuR61MEo5yG7dK2hdZRq
xl6tPrUa8dvrlzToNNhjpJTUhuPzEIMtxnnZ2ZBMo916e8d2w/r3Ky4nX0C3tjO3fFUEbTJEjjpA
dUQt+D4hmEOVu1w0ax6B2LZfFbod3TpK4d2qLVxR+bzKzDtFEge0qQ8YqN4bs54TQ0RQd7RUFzBD
p4knq+7aueoM3hyezIkio+0SpMBwylIjsRxKxIorzdyymN5jtS+A88SyczdEMqFvNu494awZfFjW
SjRyNXcBZLZEW7Ja+Vx9bsA2AwgEJIVhsX0FjbUcdbRqBrmObz6K8ADRLSzvOmGgc0NvIRop60lt
JHJUhlzZtmh/uUPz378qqHAkUsJtidrwK8iKfZjljdNyIkhTy7pJit0QfYA49JGfLM5sd5dZhTLe
0ArxttTCHmXGfPQv2IJBvmvDWZlgtyCzihlgFMYChyeMs+emz7A0kbv2xx1qx8CqIa4Ya5it7lmY
ag+6bM8Gm5vbJl2aOTpdJvtk21H7EJeAVARBQ033u6gf5d3ZPiNEff76QS4TaTpmoRR9vIIC/fiB
GiZ5uQ1ijSKBrzB19XKDNzzB3furVoTxn26LMfgXbkCR2EDwx5MJxczR0flYB0Uu3eHlHu94bTF4
RYpyq2x3QMFtK767p8ZmJQNCt1XXEArxvYJ3pLDinzXQ1VGLsf61jhvu0xIfPR1SDl4M1RPopDPm
TX220LlTIHKfXh/BZ7nzQwRYfMNhFHBf/XxlRxUgbhwGGGwOI8v1S9wT07k39L5Ra/EBmY+DMjuh
MnFd3UlfdmD2smpMrrC9tRsHj70fm9ZZSHvj0cOZRxsz2ZwP72yGDGU8hnNGr94BxlhHEqfzL082
uTxtSX/9k9/jJoXeOAM4cP+tbVm7gUx1jXLZBkPVj+doFNUfRffbtmZQhPsheRTgwNDYrXjKlkfD
wksipyOovb3zXar32XBmiNxiRgTpOcJg9ld5YuFJyh/C4Nm9xALvDejnH5FWsyGfRedd9jRUJh4I
5eSATIp67L+fDUAYsG2LbXthRXKemarcXq0KQQSxyFXuT3F27sV1DGyR/97x9tfsqUEhnAYTVV6H
hdoPSRN7KH3VJdNrq0SD6QnXAoBrA/MDJKG1JhyJlHZfA8MQxwFGAuqanybxwLKog4NlhegBoUQD
MfpelABPrPh7W5km+5FFPaoEfVW3BifVr758VFF7RWBTAi87kBZ9pd6aYB0Nc7QwzzdCDrOqOXN9
Ej1PDYq1g4H0Id0wt8VmVg9TJ+nSeuFITmi2eJJMBNqojQu7OVD2JKLUnq77cD80r0JHlnCocp7P
tsCMnY7EkZctlkuqPgOTh0mXsl0lEUgKSY/ufTqUD3brUcf7n2fbRBE1p/qotlInr9ivdz0MS0dG
gOjUFLNC9LhMmS6NHgndm72M0fb9ews3Hskg8Ol7pAw4DkwiGh7/A3uWSeckCvLfpCMCalMacbis
qj87RCNZ+Yv1w+j1/0sz6gXCf4F9qbeMqr/bmZPjK+MSA162n1PEYTqXFRtL1eHJ83F9yHC+//NA
DlVAOjWvfR+0U2hPn7ljZPZenSlsU+EIKkC+2ihytyWNDb+rdlOtG835lkHobs6Rf6kABLBbbPSw
YxRajJljhCULvOmm0QDXZ3DhSvpgarLHct6wWhjEWhgC9ctjy8jIBUh440xRIgQiAdpq2PuDrEEP
7IVqD7cyQI/fn5fc+o+ICXt1XgzxoYvRyTE3GitYIFu8QaM2X5injjwRsTwSvvY51EpO4O48wWv7
p5Wq8zKQMeqW4Xxq8PpfeannZFMtCqZhvJ3TDwNOLWznJCw7FhhBTzL0SNyJ+UXdvuTpZ4u0ysYN
z8vDt+/zDld+P8C7RUYomYV+CKQjLCg+9YhscnS+sAACLQh1STJHPfe8dRXlZxRD4x3aM4ZImggH
MiLCA9LzKkSWDphOOdptcWi1UGMP0HHhOBUamgkci2kgmGS4s7BIkUKthfVSDXi0sV9kHW64eQzD
Ya6CqAH0ZJXwUH92yyrFj/hfnUhEIhntcS6iyjQ1oRaKrcC8f3mXsmMXYGG2kP2FtobHKC9IZxBo
zzmEWWi3HMfufbCfE3hEiJ+xD2qzcV2hqyuCgO0EiFG07krFQhDZu/qKGiYtvttm2wBGm/ICehTO
Vfigp2vp02vELHswk7WbAi5q/lzxl3AhXTWaQyyPuAyUtxs4PZCxd9B7Px0De9NJxgJDPETDmRHe
1OUJks3L1T0FQ1HnweaSFRT1IliTypwoP7OrFQdcj4HOviEeYxtXAVaMPGtN8mMcRnOX1r3HdVdc
jxWOlkq4OT2Ky9oYXHPhByqklbZugMn5qMhAJoLKRcB8kVA37sJLBtqWqVvhaPshNV0194/2e1DW
BMGFVq5h3h8+N9OwXCekMG7atOL0CHKK81iWIc5L7pC8wkYPiowd28wnkK9zPWGUwtD7llvs19A0
ooHlWQQA3oSwlnc0bq1sqpyarQhgZXHi5Dp3AFxp9ML3XKfQz0N1cVNs6lBJbD8BWzWHB/FWAXwO
JoL2asIR7vFnGRY/gyKyE+qZLU5lhcaEhatsUuanJLCbDny4UT/TwAqX64DdqTazZ4eR7Qd5i3My
OfOJpc3fP5Fj1j7u5F9XJ8pNxoNS00Tcd1SjkoEWkubEQ1uJpavf0V1Ax1N6aqnSfTpIeJqv5GJO
zWKNsyjYDhdxtF/XKZQU0YHMiiTKxcxME4cJtgNrWjBSRSN6sm6iFANtxS2YGOKMyQIQesdYhZCg
bk9MUlhQ/pYmMFH8aqwkdehSf01a3stzOWcet9w2rodmGEDQ9Nt87tG4XzzjvBc43EJPy667X83p
4xkMqC5WaajCTkIzG41QPSTrDUmama8Nsx8nURyQvB/cIrFvRb85tvXfBqLqPTkPMv/arHym7oJU
BJaYqsdEqMqtOBvlZQieMSPsvqoUQuh3LV+cVD6VoM/9T4MziEqAO7Ewn5lNiV4KVJKSuvR5LhZ/
S55jMvEQMXhH5tnoPtjEFsjdmxEJJ6wTASRiqsrLi9Nn7PG1YQM1xZEupb85+qrzFMn2PA7RHtXG
COTM11+g3IwGFvfwyLVkYscE5zHsu7SP6zQcRF32wQcsa9SNroBH3Omg1zgOj/MLd1bZLeaVTmAt
1x4fLZNLlifxZ86BhrsIVVkyI8uf7ygnih06YimBI0nHZbVhgBh6fcus7y6z62TkGzcnsPb1GmDv
A1zO+lg89hgrdfoiRCiaEmxUJnzaSiMAHd6wGsfzNeLX98ZTuzizPBQDKtD0hLpxnfY/x3d+ghUY
j88So7Ku5RDy/vH8z8CkV3DDm4Tg7ApQLEp8gKD0SpmZyoHD5V3K2TVxwMvian4fJcwSq5Raqndl
hPRIvInx9hPoag61kDq7dFUtsO8j87XosEbtLGqXdC9i3JSf5/dH+k1+wvJhMkdj2fYpfNgaoRsR
X/qz1FKGl+TYLdzHBX9ZE90tM0K1bttrDryXP6G1ZMwEloBc1Xnz+pgzYLOzBbtC7CWHE+63Tumo
+JcwCtAE124AHhbJ6tIWZeRjLF+r11TBTRR2c0DwwF44TPBXxcE+rQ19pQHEOQYK8p/evWmtJNFT
C1ICjdfzFXnbPXA2DMaJxgYuTgGw9k75fEGGAlKCx8Y58hhi51MOWXjXtpBM145STbuaAH85EGdY
wmHzaYdlx6PeDd02JWY4D6G7lSPq0mam3scIhUM+D7Z35yjAGghqfJWGVnj8+seDudwkpHSonmsn
TK8tzCUu/u0ggGgJdFOuY/FicFpMkFGvvIy6FJevIINo6PLi0eaW873MDcbHVI/JgJsbujcyprtA
9nQ1QjMAK6s8403bc08o6jCluqITeZyP5QujSMstgNU7tCcBip7qC4l0eJ1zH06NRyZpj6sAMXJn
UCrE65vJ6eqhkI97k5PMwN/u96IuipxU9eLUiz0IK+iOuEYjpGo0WwcBapTpEqNaQ9P1XB73QWiZ
w7IwEdpVYVd0vmWqqxaJjsPO9wkQ3P9eT+N6jFMDjGObbtayU0heF5nxBKvhskVly2loIG+/Cvxl
I/2427qk3hrSBhNZ+31Yhe7UJEObLSBuxnLESPPU54WALv8ivgBuyNEPvtH7hGDcrtBOuX1PReYo
X8oRrks/i9hSfa/4Iuhm0sPobftti3oKZzIVtluHnOPkkT25i69aiYgkuShL4E85AwtfmpAVb0UO
yTIxCGf3DWxeVxAhS3edybvoPG506UiUGfZmtD+i1Cg3vrSZzhP6ydMfmOXpdmolACles0JqPq7j
rbnu52R7jeD6pnAb4BpwAaTaoIY2ADi4epgJNpRuEErbnvs5Bt+t7V3DhdAJIHilKQWn1p3cp6Jh
BOYkqcOfVOQDVugG8naTsZlB1ydGFGez0Aeo/xAOZ1erjFCGSvoSQXCzhSIWIKB2JGjpSsR5TaFT
A++uw1PxfJH7UJwE+3USnIx/NuRmySwlGyobCyk9ttSWVi6FnI5GAjPqrRt355GdKSETiEUMXMZg
wYLqO8yR95BQ5XE8lhpJybz7nFEfqvG2YRkxDu/lWaLSieQaYjj12BsK3v8SIPdqU6Eimjj9ZxR+
XbYKCUjDd13Yyj5IM60l6xmqXzvSp12GHLr34yLmcjVZnnSydOndJODPmY0PhHTayCVK5F+CQgpi
EI8NGAc7iZPKwi4HRWrMVykvnNMxTy1NXLqOGXEeqUOWWZeZoT/gwt5QxP8pgohxQSsy6DZqVJDQ
GkZ90pgRUXgtezTUeii+m1s8tLjB5RcGL8ICP5iyscG6+pEuuAqvRu9TjFXCt9b5i8Ard4ipB2Ny
EkxIbQ5DiyQo9EfmO2gsd/rBZwwz4T6Lito9VpIG/ZnrQUN7gxYmwaQY16MgZT0rR1PUd4J21RHK
WKa/OvRGmkGkd9Y3n9BW66hMCNPL2EJJNhEM8u23OoMf595YSxSP8fU+dF7LkQwC91kVEjp7k6Oe
DfEu/whZYCcbTtguf3jCDyhNlnj49WrJx1EItJ09CHs4qEH301mqUhNGPbGBzUtoWg32e7WXSJ9m
M4/1v9UfEpCAgCzhSlQZia5gkGZGPPZcO2YoqhIDGQE1wBtzY+ABSvFLlxQfy97ws0IkJ2IIHB6E
0BqMqfPGxGF71ZxjEQ55HXX4aTFrmLksZ49W/qflJf1YOuSFndRUCd8ZTF1/vb927jvC9rbf4nbn
AoPWAov04iHofXjs0SHkTI1E51Pw4TN8HBHFKGI5MBAuo29Llf8tx4dgpvObR/JdlW8GaJvUHLzn
j9WZVgrjf2lYoMcttjGJAx+zksfAxZdnyBLrC34A+RM52XRL3713zJLFQqJrW4mMRXz6lKnpWlNI
dHIs4H+d2R//27RRBemur5c1biqZgYQIiNFZJ3ztmOqA+wKhHsNDQwK0EAFe1Rqd5vGyCs092sdt
M4EOFkml8QQQYKDdWNNiGnqxRVU8f2YQ9N08dgrOPgMCrKQ2nY2xrWbichzosw7pw9xBf7Be6yW0
j0w+bFggW3NflkHaHKL4WmYye0Kwfy34tBBph1X5oINH4hAFH5sk+iuL5FCGnwObkuAUWItt8dut
KQB/tq2e//ycqCXL+anPxFemwjikYEmZxG9YUZv7riFHqsaVg61UvFgNX55K9TlCv5FPKUAXaDPT
TVeO511bwoEDUn6qIxiVHRanw892gNIdePo5CQW4/RiRSuFWgexhGpzQoxB3NxThHglWQU3yNgEi
77/K/5hYYpmyQhGgepUaHbuVTqwbjlRtLaPXWovL889PlXjsDUL1iYU5EC8uzABltUsGY7rZUVuq
NulFle/sSC1cHtXvOPPTF2NeNweOuw68Yo/Uo60/6YHHM5CP5blTX592hxqw02qIb+Pd8hOy0ogJ
PyHb6cP7B+6Vkgg7o7jj2yM9OB2eEPj8yZqnEREy3O/A0XXLbGL1Kvtk2Z5OrVbCFZZZ32MphljS
RluRV/5CgXxW2jI8AhijFJqh1MOkgqibW6pK3FC0Hqfm0ka3bzB5Fu6/OIFi9rj3rdET/ffSJ3HZ
EtTRVs0ZESnLQSDh/OjHLNGaNGO1pZU4S1Swd0CalEpQ8mIqk7NmN6xlUPWaDfg6jUIDU74NlJS0
W+hfCGaz3X8q/s1vCDeQezyZQjNp15u6tub2MJY2y2CnrU6qIOVTOMFDdXh7YCl3tVBxcNhpbX4k
3ZEPujuoX8/QQbZni7RAfyiNQSRIaWtrNhYtGe0H5hbRsltFvSjNkQbJOAq6tPR8MJX0Cs1WMgtw
Z6iGrfpI9IkFhUjww/RJlgLO/KWaNqpBD7b9XRpoJaq1ocPGvzDlvVmwXocOfs7sdyLP1w8pc9+6
GdCd57ILn4zIP47biDZ/yM2MLzueYpF8Gz6Fa1H0GlPhLOrx8qbmAFWoGwBTuaEQdSLlb1lJ+hMK
XsjO2/sCOmQKtVLNXtwqbzS+1xrJpJolztV9/nRt62qKzsLXtBDY2ZqJwbt2ax7m1oYkRk/jJ3lD
nhqpqIePNIUDkCASNqNvceinr2YeG+gwBCdO6yujdejP/ag84Gij5gpV+k75qsd/7UtlQwYM5bPV
LFfx+4GKfBLs0Vxp5M17QxV0Qm8cggqeIYZjMQ6R13QUlJq/wf+7Sk4CEOJ936mzQoZp9pStJvJU
IHt35TPwQpshf1fXwW4P84FWboI63J7wEZ46mWfqEiC+2yBd0b9hZJVjgPSFJet7Q8+ATs4LV9fC
/VxGxUrqSQtIx4ppgZ/9jq0K2ouP9a+fQXhS9h5/SuFyJ/RuClGmICoALNRMc7MuhE8Da6l/YuKv
VgNTtuUKNP1oglt+v6iTN6CQQYqOQhaK9EpDajNQrXBMwIXvFNlx9hE3x6x8ss0A8iBVk4CnNHZn
FYPNQAC/98sQj6wAPu4+aKXqauPj7B3fxxye/07BcRMLwVq+N0sqIxofgx8thTYVxPNO9BwFvtXj
yWTR+l+8eu55Vnph+2WyK7yZ1rLoTOl9UbkUsMDHXhM0zhR827qU67PDvfaCH1Dpnz6WdJ9IGEbd
/gZAe6AR5vBqF0sS6uSzkdqZZev15XlFi5erhOh9OPty/M1VKZMV7tK8mAs3vWwmtZJAHAVcRV6a
vJ2l25BRIQD2pDXcz50OwF9/VaNlMHG1y0aI8Ri/s73eXzoQwLl7XWgWHx9yvxuq1G4PavKdQKV7
W6UfrODm2dKWq7AAN7vsCEunQSxjuqFYwe8E3ImNuwlwVJcG1RiCWfbgHkcIRV8hrRP4zoGnfBxj
+T2UHmschusPn5rCnYSy1UJzWRnYMXKLCvOUUMm+4MJjGHoTEUvWHrhvJN1PVpnY+gSdTk6dohIY
hUS0OTxOsvxzqnCsC2wtZA0+ccdu3eRT1f9GBEOUjRybWKVglou12+DTWJCYRRtNlUCxTKw4Laso
XTiZ5Hfv7DlkmBOBvq6jbbMFzzK/H/yF+5fZgrOve5C+XR9A+EwpkwFWJW4qETOF0pMz4GrLS5Q5
YwM7FaBCGbQhPOGcfJIoA8V6mJmUH3AVKAYHXQPnGWZJH5ynkgKVQjVPvTW9gEyLjw8uL4zPqd7m
eXM8uF5cMhcb2CQV4pODizwWoOYjKqZAiBqpuDELwNdVVw3ZnNBmpXkgelHKWTtkKu+2PcWXKTOF
1m5kUKPcilgZX4jSHk6PxUox04E2yxg4GX5HsZObsnEAfjObqoIKWM0qA1HVt6v2Ur2PKWS+r5XC
OI/8K9wuJCZdiVy7V3/ljxBp11uVtNJLp/jaHsN5eVm055j3av6qNNkT7wjuffaY1UMnA9aHmZdo
J6qnj4vJ5m5rNsdiNlra2N27mxFHW5U/U+XqkfNV7CON+GNK59zn53jigb3SAv+/GhauSSsZ8XN8
R+9cg8b52606kbngBjWVdgUys9pDfdjC5UV6/y4sCG7Tt7b60o9b6e0xTcqmqVofGGswsa+0EtJp
3IRwPQlRR126ELMLgru95o113+jewEFPov2v9tRbTXeEOZTYOsljf2cORlWjzo8rxNx5F2CjJ0Da
wH2RLf81Huiis+UVoOMElpnTyUe2lulkCtpepLrBVedcWXFHJen1fQSMJRujbtHzeVYkafDEOVS5
4t/VKBbDYOC1EBPBsLyWbTDt5Kz9fYcyEo5NOfLxpltUhjS07dwD1va7i9zwotrF2PJAQkv/Zbde
TrVXcx4griFaciPms88fk5JYvoHyG0iun1ULNP6zaSdFdQpHPW2JyJAGg7Igrxb1uEH+LSiWRYgW
fDGGO+X8U9L4CajtH2Rv35d6fm78qrHFHa0I3ptwgfcamo7YqB+XzVzhbXAxLJ3csuMG+RQxIoBE
jc5GYtKyOs28Mk5U6GjYTozlB768wsOisNkyxfaA5SAUCL48jccw7dS9kOUlIPGu0a6c9eRkcUWE
GRWiHPJvMXVmqW61LiwB5sJ+97BXTRevgZ8hs8pFjvnEVB02Kfblkbg73rV9/Vetn7yIU1id2K95
HWTmndb6BqJI/CfU+ITweFeGdITSvUas6ikFJk5i7olDm9+48FngtVGozH01lENMzoKdKW1aDJY5
Kpc8rYJIwTsOQOE+DttXKZOGyG+0MdF4txd2KZOyJ5PzaoTHlgU/nHlKi6tHgR4/t/71KbIGIQ2L
Nj6pV1qf9t84e+69n+3HYxwadu4J3rOZ8pvlhJBK7vnP1aO/GpVUi6gSA12NVccI9BRJ/ewGuxUG
XBMTTsatmfI9t6WMdR7Da1kHnFkCp5AKvxlDNz/UZbcOFUVhvGa1WD73ees1c3IaWolLFzgEWXpy
8be8m4bM5ZyEcvttgXRXP0nClLIqmzG9PktXu+N1wK/2p6te0xLDzCGquQFc2R2Iswuhb+sBp8dR
lvIvgZLaaJ9Uu+LBF5MF57771pINRmJzbw8+2pZkYIWggI7UwAnDiIRyEbbhIyz+t4VgU/y9HqDR
XruHXspgH/ojZzRgOFG8Ww9GiUoNefDkF4zX9zsJt8jGn3XhFw3OGlWmbnH4s9Z8YDvllHHBSpjh
I3KAVESgkxdZOzA26Fu/lyMj2AfTTgeSxQrGxZRe1auZwsA+BeGQsqa5IYLrOl8e+uho2IxFbjtb
NiHbO+Po6LnQg67u/LHvOLJLHZq9Zng+bguxZohzz9Z9M72zCOSJwUAUaBO1YOxG5xXzMHSNmT8D
dKINv7QL5flMljF2GQI1avfv664zU1nMhsyISOmOPhzLBkMfR/9WqACo7Kmp5d/VvuTDFIW/Dutl
xZ6g8lWE1YRGvoIUCg1KyLPkyQcTaysg+e952mPYqGgRD84zcrHWc4qZhK+xenmjG6yAbhfkdzE1
ZW3sk5bAtq5aBvYtDV3lezOXgM9w8RZEfwMGmH+eh2t5WeHtk5+V5Z0R4/UbGU1oVkT+rPiYMdbP
D0ANhsnFa2SVWqWn/eX7BpM0m5hdUbclKukbk/lYgXloCkt3maZ045uGqtmGgsgerCz5RYEpzAas
57B6xFdWKRMcel0gjHpV71CAf5yMAxNcQ+qduUvZFn9HVsuKqnmmIaUO6pW4ycHAOdGnF+iKx2O2
c/ACv85MtRJ0GlWGfV06kl3FOZCtZi5z+FFtfoWm12t94XmWxeIUtrx1Km6yG970U2bL1ViwygQ2
OKABsBTuoEl0pwQcTR5iWsF81NPRDMvULjFcl00/HSSiQ99EdHLEtYyHjvxLr4AZeIjW+AKwSXwv
0U2TQheDr542GokkuDV56TyPDfjYH9KSRlVEwuW3uhQblxinWDfijplO2lZjHrjFK87G3I2ulA0u
N9ZAcVqrLP3T+DOBs0jcrTb3AeOFx0i40PVSwa8Ly4bt0vFQd3Oas7ihK1H3g7AJKQQ6AbmrZEP/
4XrZn3XZuKkh5+ZMoqhMKhCWMdSUT1JL8iL6O9OaVHL+zlQt3bpXZdwcSrw+ZRd5J+Qc5TKyJtbd
tu2dvzvzRlOUvVA40tzFwOUDG9yqRwnjm9iSG1pvXP9639glFCNDUatR6VFgnzLWTC5rSCn/WbHN
GEj+fwv4ZYQMkVLZfXutJUDMle39qxtN3phIbP/ERvRlnPThvUkuLF/o9JE6qgeMHuVpJCmRJqYk
KB1EhFqtbmPX7A4TKD3eb4dwscOgprarLB7YG94Xlwr74U1HfdgN8oW48imIHvl93EvnVzHGYZpn
V2STJn9N3JvKGjMOyjWQUb3wEXh43TBpa91/OqIstdXNo5iPH+rTH9BPV8uY/CuwDw/ifzhegbSW
unrOeIjWfR2nmkaGh3NgmnuBxciUxSytDZyNx8xbS9Q1GlWA0f1nFxrdUj0EhfEd2hlxOQUT3O8I
aW/rOHHz0ykwydwfOeTJjk+11StYqKPNIsSLPsQHCaxGateEmbvGIPktyoezcBi+hQs26btHqrD1
TiJ6u8Fy16JEwtXgJbKxssWqwv3xTe7aGAavZns0n98DqZJeC6wP0dDfjO92KKKfmVLgEvWcrxbl
bZjk7D2oEvz4BET8+9gPJdmCSFBUGVLmvf+H/5ONly2tgDPucbDwb93tvb5w9v5MAOHlprLBr4s7
V88u/5WJj+YPOsfqqnm0D8IjoS/+YSw15E03ucb87z8zO0Q0C1a5AUtALrZcopNaKfxWnm0LiSa6
ixHokK67os+FVXpRXsVDKdVElZe43uLz4RM7phZy5ZpKGC/8VhJjf4tNA6bryB2ZpuGcfX8A0SGS
xJrU5I991a7dLdPKlUrs8AMGXAG1DptVzDvQRGp4ed8fnvWEHdBeocJ2/8CmzQHyRBHWRDqdOM4Y
PvNnuWDLtRnJZJz8kfLCXxCAIJEBJihIKB5QNFcBBACqJ6D8YJZtKjTePjwx99hG7oaMi7RIgt50
Lq7ct/uHDld7H/52GXrNfD6+IkOE+ahxZfhUPkvnK3sticmMvWn2W0tQg8SGJRcndtXQAxBlT2iq
oPuCrzOrVSfQdbYutjl6sM2pUZHqL7ahrXyhipBfGsw8mIFzJxVmykeRcdCF1j+QgRIFIMHdMqrs
8hNYq1P7U9Fo2le3J8AXgdTaDfr3QZQ621P5HmGyBlLxOqap/ZchTjLwJMU5LwrCRUbUISuixJme
TVQfoM3Zqw0Qg+cmFy9Lcl8buIkf9VDa70DKxUfQAV4i127V7hu8+47FGB/QLAHelGsRud1TEFRo
nd75FdGr6XsE1yGtkHcrOr6JFYeriy/W0cT7JNBWl1kqsXRJWAyLxR9P5ciKhT+twQoLCvUhnH5L
tuFyzUaSP1nW1QHcJfXJXJHoNMjhAfi49DH0Nug+ctUPkAoK+xKjB1JE56GuYGcIv+GiGD2Bcs3f
UFqirQKJktRNX31FhjMftzxWv/JWWFHu2uJYKmJ6iCj5spgFpgbwKERB9WKCU8YGw5IrfNRjiFkQ
9bYHVly6JfI5kdn/4lxL024AnIMqxj6sAKzM1k8qF8gHO8wGYIkX0ZtwOuafkOe1Lw/rokaOaTVd
0iOkpE9bZlU73e+c4osBZQVJqpEPHE5F0FllZ9FgCVEdLfRcSY0CWDIBO7m1RkkHd5VyaT4oL4X8
cYrimf/JeYCwbVI5WtImp8XVG3jUjjLsLx8pOS4qN0l83CakGSJpd+HeSLgzLWIH9YvVV9udlOXw
eIJymLDOtnY3K8JPVU2AaF+nJCn0KrElLmZotOTVA32hPcTVdev3DR1Dc75q5Ug2mblSVlb/VFun
BXWLqR9SRgJKc7N6Ym3PlJTCdvW++m9vJ7KNadCFHr0KA1zMDuW/BfwZxwG2XMSo1ehIOBxGn3FO
AfuCz0kckkmqvpah+OgKpWP6sBAu4lUudJcwYDlSEe4y6f0G8VHhOOUqMtZSsW0U8GkA9TUigqg3
+DZMoQrJ25uPtdCnxeNtZGyWb424s3Fziq8+KdgDxXrbFh2htH9qEk8bUaQoAz+4gTOpeA5pbe2J
PGQqm1eUS/kvFyKyTdFX9qe/DZWBpCjDqqnDuDPjJnzwHlf4wloTzL7gkH6SvUTkEF84DnpFt8Wk
PXiAV+bB5sbLdWR24o5oFADjbWz6336e/zIoB0jwkTQqKGjd88VdZ8xLtJac/HSVCDzcRJSikF4x
u5IMTpbxX9LnVPqm30HvHvqoQbq8J3JIZZh1AFWpqCrAjhvg+u7R7q1Z1DPi2Kvh+leS/W0V2FVk
9WJhTEECFUIwq6CEwtvM3FUf6pmHaqXFx5y1+k7hjwbA7I4SUhn7Ptp3viPwriyfkR9FvhyjSlJv
R9FFOToxVAz/uGpHY4ioSRl5RtvkJu+4GbGC0R8OABQCmEkC4XreysFN6BNRLoZSdRGyGJfV4sCW
bWs/rOs228XaaXjATWlTz+WELl8fe2KBhwpG2WBoSjyLu615lwidw5D0sYDQACjtRKEsmn3c+E6X
tXOqrrxMhuFd/Je9IBlJIxu6F1L9f2xn64DrrSr1v3WoWALnrrI8Fj+3Gyw6GFPar1WJMgNLcWwK
is/b2bE3TqO3blB9dYIJlCEZsptTDJkmLVFhXzBZwsoaZ4hSNrHRgK24Cr/+QcGqgb62rDu8JZvm
7bO0BQutqGzEF/vK6QxJb/4kM8flz348NadR3Sicw0hdz++VRlMXAoillNYnFItqq+l7T+toeNT1
KwUbgUm2RssifHG4jnrsjnWm6ReacU2+WHnNyrHIzCWHBxkC8n47kmsaAcHE36H0qnPfBX0fH0DV
25YB+vs0zzp9fVGpQEQCevKcVf3aeEQMnY/qgt3r2C90NZfoZpkJjQ6kc6t9BlvJV5G6lPMaOjBo
+Xq9oGnZKeHHkCEvLHTvuF5uRbaJaNFBsfaEa8zvVDEfPnMpP7WX6OJQVfc3RdSithsclhchT4V9
NVCZvQX0qCvKMyPpEaYLfMwCi51I4MXnli9AVLvDLFuu34y93ECribmCVPtRYaR7ExDA5J237J2+
1jAp6EFLand+Ww3+9CkL4sXoT3GbJUHft9OsrRZTb+uTB9VbrgBTrH/EUcw3weOnN74EGGJHR+8Y
zyL0x/isqI+Zus0TBA4zt1h3C6iphbh0d1rFoCZYJRdixBjh+BI0RmD9n3ai9SIzp0Jiv8j5sJnA
NK6xubscqs286l1i7/arPrOrR+FLwk8aYx9h6VoOSwWmhi5hgNasGMRdGqTCyLfUmSC0Sgd3nu24
+tLUcHRatZkFt/SyXh8ixl10XgaYXPz0mVAkj0uibIzSFklA5OhnoqUWXzd7IPuAkwbHcEkBUrYA
Qa8BNhk1wjCw+gQb2x8F1ZY6+vxf1A7757Su7Lu67RDYO7QPFfVn+VjUxk2jbIt/9gkCrCWMn1NP
fxXfV5jHfh8nV80wBzUkxyUW6pbrA0P9wTRYOcKkUsJVs0mq3B2AYIIMYWzd4LptdrSGEwmDbJ6V
etRFSN++Y6AnX8SSldli3Qs7BWOcItUcxx9RwB6bF02uxjdf+yd3vvuLtQ54A1CBaiM91Iz9ck3T
CvOIdyOEo4h4klZ/mX/4/XulSwdrBCaRidEVoPHCKZV/TL5dtTzkbA8V0h16kbPOb7Jfo0hYUSfU
XNoLdCr0JVpfjwS3EVp6KHZ8zmwtKxu/EAd0CuZtZdKlTDv6Wa4iWiAqLN9RzZKNsKOKTRQ0/zzQ
DdFDtglvZphOP9qN54LvXThhrRMyFanv1uyfIgfPaazw9UZtkfIgelwz21bxrlXT5j2IkXWGMlWg
c11XCD2bnjeFh+IsvioKCJ4nsOA9TNHrxrCIntaGyHt51iT5SWi468BnnJFKxvjVa33SBBUnOMSX
ZR/iufUxdvX8rayPqIbUg7Pt0ebrjOoeEzvEG+SqPwgPXLukNqJr0hT6lEWPMzrrtM2mIkGyfEjP
aQ6OE5hRYEPxmPZb9yBiprv1SlpodNTft8ktCNx7tblaRj9hHp89wYzsvX9O0joqAwnOgJsxQKaz
M/4qYqbSxhjWuEDeh7y47jwbw/D+cqMLrRS3OSZJpR3xr16Tfo3eW4nsPwJt072BPtZyxT2kS7GC
k8dyrdn2K/sr3iqrLpqC2rM/CItwIq6qLUJzoeOqNFT/39zkhXrBRn0yCh6C1uJGDtEeo73infT4
vCeg6cqNLwe6PEqHAh25Io7GabLF1XT1QiD7wJ+QHiL/Ieih3Xyjhpd/UqDwfRcizgnn45B9Ye/l
NtA1GdaEt4vXcpcXmDJshBCte9+43RgodPf5mZtT7Jv/ds5vE5eKoa6/aaWEHu02d3+S5mDFgbex
ybUG3YwSIhpjzkfiYscaTRPKCzd8BX+aG//2IJWD4177t7uNl3DxyjK7z1YrZF/cR66Drk/tQcEV
yfCRMz3XaOZU9yTu0A4kx1l0W7O1t5HpuhBUWu26umgiXt9+yiHd60PbMaDSEFqIdt9m8lE3txfa
celtqEpkd3F0dfTvi0W7hJDTXNd3+9fDZGAG0oc2Acg2qHIdqlbv15oRjrzgvX8PvooJ1+o0dB+M
mxwCubeMl1E34uLBtD96T1ejIktTwHxYR1k8dFqDMc1uE7d6S2w1QpHF/+jQN37W+CBauTH7oJo9
9Mh0vENmapYlHMwISLYScv4FGoE4So0Y+x/vns0ltZav96RNmxzbIRNAIFFDzeXRG2fVGAPwuJYs
oYh0bR01qeImKtIwP00Dfexq8jMz9A3qqvGIMsEz88JmcAPWclyIvki24W/48LhqAkLzoHhRYs9f
ANZbYXnRP9nrtoNe13RFogTmZjeW2l2DO45q6nJKf6WMlWablry75BaqhrDohpFpR5iXVMPI0btV
EivgoSPDf4MrncifTKFlhe627MA6Q2hbgFWvQ0Yzv4r+rtDRSUQhGZcyTchV4YWDEW+b8fhftdrW
wPAIenq591ZtBCvSNaPnxdt5X5wELLhCMYG1wUYQEG3g7EolnXwyKryeMdLz0aorWAP1OLoE4XlA
egDxGIejpKncHGxkjGWnuTknV9TIw8/p4egmmMsZtryDrnn0m2HCCaYef/8HvUPEYYiP0a6c0xD0
ijkNU+wplenIPojHpTTSKkoPkcKBX8nNRY4C/hME8a7vvCFc/HHlSxfqs6HFr5dBNja9DSa+k4ui
eVPQzxYDlJ9VVmpOMZ0hrChqNvrgkTOYHvEAL5ePB4UZ7ttgvtv74Jc9DLkhn5H9WivtNFpungiX
P/6ii4LT/FaGoV816nk/rvLDaqGj5ZKUKafB0hDGnH9gR2Si5h5sn3ST2RlKe0IiKoAZSPEJ7SHG
upz2ZF2ip7we8vmiRdnRQiFzbcPH3nGu2aEO6mgoBms0/mQlNrY2Tv9xhr/Zzoxe4TCmB1e8p9Y3
41W/PT0tR2ROl5d051vdlXTx6w2QBIj8fIHh7AiXDuw1KUC4edEXMykd6rTA5+nlbvx2DsbYKpOY
KFVhUHQ96fqzox3gckGyfq8gVejMGJnjyDtLsDjVjwsYqV7KhjQFCZHFkKl7u/tgXoiLFHFSG+jG
ltkStOrHxKm1R4bWWfec1h6eesOhPKEVbSnRu20LLxIcYcbxS4M9ZSiTgxKwOFy4keuNPGPKkxI8
3+O8w0a8DNLLUre123TSttggpL4nwLjuB5KqRGUT40E0vb1Bi8Ax1L8sUEPg5dt5bXuf4SmR3ivo
xWNx+zSZfWKJ6xctSON/hz973MQ/LwQdnWr5gfCmCXRGbCjDtl0L6Hfd7LNNgdyFo1CYtRsC1GKb
9zsve935G8RkVyEGHAXJIPfWYExhQC/p9JKxZxoqn6xKQDxiRApD/MUvdJzvMptP6vC4zK0WIpoA
CuHAt3P6yGfkp6ROf3G/JA4Wx6cfLFa19JiJSuXeQ2vORxKakhpAp21qgNR2cBeujOdNzDVgFHkH
KN7Iip3WvDdBY1R9KWwcezIt0Z1xl0QkLvA/PnLErDx0783sHaiUOFJ7e0jI4KKm542nWs25pFEe
A0liniz86CjH8gFVRBWCSYMWMGl1x/QQeNgngxH7ywsu7F73maKNEu7Bs1SwVw7YKZOy6Lg1GQuQ
R8GtzdBS8y06Fz7JO4LXu6ZkVpPcEV9pi1/gQwORbIpVX9PVlXmc6SawLxiW6lp4jp+dpYGDbZSn
naiOLuNXbAd4ClxqSoWBc11JPW8yXiv+dJXieq5H+R+MZJJ/WJ2++eZT9IUjUl78PtUzm9ZNgKzL
I6b+4pG5fxRRrVF+GeEZYAlqrJ0YE+SVCqjvI+y0Pe/8Z9K576SjahP+ZF9kPcXunAHY/1gyrYpc
+vxv2EoC7nzHOgUfPBTC8q0TLrKaJjdAkKi8ZG0X2qduZC3YuYD8vYyghXgMLILf7Cl3MBWjW4U4
wrdNL9q9nibX0CvsxjAgolEuZQ6ovUe+351U9K5eNRhDEASMx/TyIrCBoGVcDHxJaPx3E+GMnD27
spQM5Xad5c7y6jz0j2ZaHiYs7AZFEgjdlmxUQRWBOK6ISPkWnjfOUr9oz9MvrWROqte3oi3U57AG
KlGhmUISe0bl2vTQdGeIX6qP7ISO6dkC9Cu7Z+4C3v14gG4fJiki/WjuL14p5vQmC0+s7zen884o
YEkIHu5Vqch59qk3D+89huFNrQzqyYqyzaTZshUgmxpQ5NhavIzdo7PzhUWk9vLX+r+IuuSJDI3j
8e0/HvYdgva8/NOkhivfXCb9q/FNfiMEiFUkylpfbAL9eezQf2NpfVhv81DQ5Pw7zAAHJCJXrvH8
/FRLIP+x5ZgXRYcrBDEoAz4WLrHfPSq+yQ4gLvtHLDMe/R0tVQunHdAxX94iZ4QM0Y/rems+74N8
uL4nqIGuO5k0WudLL+FWh0tfV6V8R40jqdj5o15kWC1B+klhQkXmquM7bokjxJng/Yd5/UZQKfq3
znjIqQadv9ryvsVJgRWJ08b/Vyq2ldvUZQ/vLg64n/H2mgXnNV9eIDZER8mDuZ12Jac5suYMkp2l
KwwAnhQE+860rW9BUqJgCI9xuBjQi+52TeSREMZeFSgcqTVyoHN3LK9rzBzD8loSOZ+yAle6F3CT
7G+lVYe2W2ZQgOaSqspu+rEv/x+1Ecqgef2dZpifJ2L+n7nLJVbkpZNvR8rCnhBuZVQ9X5UNCuMP
ZM4gIFUykeqJuRtr1j7qcSOLoALtYesz9PVu2JLYU9WPFIfgBfbcujNI+QP0q1Pqpj20a4f8LNsz
hNp/bfsJDdsZStkghh5SMLlOSHiiDOz80vzBGMVCzfSWqI0AFG6Q0dY+MfDi8LyEotgwYg7g/huI
fgqLPI9DP4CWTFlNwihoEDV9RgEBdc89EtBGLlX0Q+AmzGC5Bsqm9RNBew1irS9qsO5DhPOzG8cs
qK7m2PaYL6/94emUz/c3/OkzFvNdRjkDqcZ7mFv2Qw3fMBCyIwB1U4+CSBoDniW3DtjjRsiRtuiq
4IGon07Q0d/K5Q2WhpBFazprN55wzwUh3nkxiAljr1w3IWp7eaA3VdVYcExjYOT517/GAAn+AYzn
BPHONrorSR84YKaCMTLHmQ0XdpRMpu+yOZVG6EwGQW0ahecplBZrJX1CLPMOuFnW8YbQO+7zz/fc
5G+ApEQxu9prk2KOwFXrkfiNgMW0kmWmosGaXUnRlvFo3HkqYOoSBXdE81aEYU58Ggb/KfJHFoCA
vQlkHkNn2Wro/gvj3LaErhEvinPK1JuE99bvtN2+/PMb9ygzVcMPVtlauV8uIXM34p2Zcvl9dPaA
mLnKYaTrs7DnUohPyfpwSWYyBGfDCKsbZszGjk1q7psXIXlfFMuQzjVO1qDtwshuCMocvUsMwC/l
S5zJ6dwapy4AYfkxEHNnxmpN9gJHOO0cDQCRBW9mPhGszDiuIX9j/o069A6Iw+qb/4JUqLEnvA5M
rgb/ZgEaHiAeYuC8HRKfr/5geSiaslaG9RcKWVung4Jy5sOXqDHpYrzE99ZzOm+j9H9B7JIwtBfg
AXKwnmQi5eUiZ46u0DRbhFKmV2/hoWfqklTURnt6D2gZBsJGl21LKBi2sWTLxvoBKNcJogCLwxcc
MPwZCf1yTqeRN3ZUlHpOqHuiG2v/Kw0EDu2SZM/mXOwIuPzSu9GeeLDge6rmn5jIg3V73R4piEca
LZSWlrh1/YJgoFBP1u0uBJBW5UX8RmpJ0KJs/ae5/ulBB9cvH0awxyq3GKtkt/vnUrDUU14bnf6f
U8oLSr/ywPQEydDj/aKlEA3x++UtMD0dJFOambADL9dE6dNLxsJuNDBTNEz6DNLR+XAqI+WojV/T
gi5WlMHmJQEIKV0TPb4nta/cPCIQ4OXGOQiGW7e85sJMBsq/t3VXoZwylWm0dYp/xtoNnhA08hz+
UZYUOyJ/8oFO8RuQwVbixUFAeUGRl0me4vOxFiABmSFmg6ij4GZWiEMlEbBhsBG5SOPTNwFdiBzI
MOvS2rb7lCvoX77brtzUAt8inujMv6Hzgc+elb6fjlrq5tU+hza5ebIpKtRNd3DY+tbFJZjk6GgE
oAoGFNYjh7C9e9xhkX0VKsUfnM3zP6nqmsldAyC9I7aAJtk25n10vkadGgRiOo53QHmrIguur0Oz
MJ14BDgVzgA2mrw80ciGLfz1m1Mut+4JyuOE3VNPD5nLIU+A8V0g4bGUj/IO3hyxGYLkiBnYzSri
IJGNt30uG5B6OUaVmRPA29tdNyQR3RVYrBDKGpXpUmCW6ZmuxZUFXX5vSaOfYwVfBi/Gd1XqqY4W
LDqF3xjT6gRGhZKlFrCzcC/2gL2EkYZqXXchMbwnnNzAsap+9o9B5MoPq57nFQxfsegOA6m1ksib
5QTtUomNbqZYL9E8yetvsbufy5EAivUxaAsC+ZhhKEP45Hsp2geUgGHeDsiEOpzRj+u/9poq6WZE
0hl6VkvSv+EqGcCFSkYLQ1Tk2uXP9z5h0cW6Rync5FXDPP/E5CRBC7Ykrr1fYnP+C1v+EX8lmf5W
3B/JEOA+NpDZxiSDqXTdVNhVgnjHqnTnjxPKzYupYVExfv+GfUqraks6Y7xNDT6cSu1kYUbOS8NC
v4kBfoSXjQfgJogRGLuxinDv/o5L8BWRwXgrz/HXjGlk2HzhgJ2G7HICkWXLG9swat9rmAOXbTdm
pb/FRagItNei8NrDDvYqVcmIWNbP6og5qHDyWc7EMFnaptmBwPzeQFPeGf2ndLJC9BCfHCTU/ZK4
BajtBuRU/J0SYwHuhbZXaiEdGCYKleyrV2zU5Rt41UOEALEM0d67gqLzhB0I2L8PkwauPdjj6vCh
t5Ofb/dK7Re2b40bYb+w331JBVuRZV1ab9R0aQ3a8P07PmtZfjXiJ57Pzm+IdEhOnBtz0VZqmdh3
xFpzuVrEyjDS8NNkLxC6IiPa/OjPKRZytW1JHoid6O7rzN/WKBmaDECQ8xfoGTqbAZjdK+0X6RFp
1/FzWMxiOJxbzVwpzX9sOu7Beje6cXIs5pJA8AIBzfiWBLc75fwFPm4OBHlVBKUkV3c/OluzuAl7
6cAwN4fVfxyZ3zZA64bXecqBaSh7dDjrohcCO7BN1CS7mTkfVDtjoXwRbgg6FZ3V9Wdh1NSgue0s
BvO7+zVskkjdIP5PBkCTgMVQOeBW1eFy4KgLyi7pRv0TxgYUyk53mnhXgKYT33hcvNL0RC0nbQvN
O17Ck/fuMwWPHOIDfqcA9TbUnLana9Bby0Aov2JNfmbQPY7y1wf9DmVln8xO2vlUou+VHqwXTN6X
fnXFKxCa4wOva9ZzNA0m/Vk5Y4kQVQUx2lMHnpJtvEqJMVg0PYepQPoT8S+B/XSQvyDZeVoZawBZ
mAVtgIpJCHbAEzYj/+VrVpbWqm7vEDWFLjLOaoaUQje6DA8JVHnfLFvpqImX2Fpwh/WYkXxyE/Gs
W2OTH6rUpi29FnUrVMVovrO0Fe6Bd6cws7f8Z2CwnUwuKuQlD8sPmiCI022x7FhNamSvAl3A0oXr
hLZwRXWZYzBFH3mvUHsd6SMppqDO66aiJuYJGSy5FNC3h34j52vCBzHG4HlnrdGYxoQRa4VX0DgK
QVtUH33eV0sfY8qLpxe+APPTL+oudbg4Ijntfr1CYijQI/WSLWzo5P2SvGUbN2BEAqPEiYG284xl
zSJtE1SOZmC9NyuE4mj4o0MaALOe+MdsKBi5w9rXsTfoW6h6xqJY9/UOzcYUjpRBt2+17i0I9Q76
tayq3JmNR77wSPnUdVrRt8/78xEk5o7iIAnZOV/ET1Evruk0HG6zvGNNvjeAcU3yeFtKq1wFzacl
nU+1Wc2bDQCQ84/UUzhdW4mCEsEvQcYrSoJbtewhH7OKqnqd4tvTMRePEsr0T3wQWkW0jA3ehHLj
gomyVSxo0Qzll3ViWKX80uKr0jD4/X30LJnlBH1LHLne/c4ehbmcOKBgw8NnkkicPvH+m82QGO1B
RUZumeHYvwErPrBbY+4jFRN8n6KN0MsDpC4coLOz8QhdDnsb9zbWasSO5+9+7qzPK0MLEe2ZGhrV
9b+nCT8/EdhdBmlZTGJrJojWqsuMaW5e87D+yauEKTX0piQm2e8rBhXk66YoksshZG3+OGWkr7Yx
jeaClkPrRpgRL/zAHgr2FgzGxMgntzV6meDCbl7JjOAnUQGtfkGYZw70wAr+ZAFIaTCnDh6Mam1L
d/CD72RRRjTUxl2UtEATCXEqEbdu8wWwHZy6znTFCqqnQkXV6bV2Ul0UwrC22vWpibvq2565tRwz
w5FYMxWwKjCkihtwJPZNk5YEQF9ksUQkHKPIgENk4XFtqVjEHyttXNV1BlffKlu0yif8kR31lpot
40JW3OxDEZiZJe18VGQ2EgWkVdYEOsNmf/kU1WNk+qCOjn0qbpN1AZI3h+PmGtSghSExMshR7JWA
p7Oyioi0dbKUMAK+SQ3kBYd0UuWBqsjC00vrTFAkSZXFizyq4pMy1MyxXru6Hamh4ZrOsPR1HsUu
k6u1LJ8OBW0lGUWs4LBRQb/mdj96ShZ6g32ZRF59/YTaw1W/9Qj2OPpbCtTKxtpJUKvcBhOcW0or
GsFKu6vH4YW7UDpu9XON3IylN7vlDq4qqNgeu+f0jAGoepuOeheAbUnehH76IX5iT5MbatYHAJtx
A4UhTY1lMHfncFlxiKBdh4QN7ndF+umpIKhwOirKCz7c9lzjaceph6VmZee1MYAuBeqxiVs3Kemi
FFX048qF7Qgz6O7c0wW5uEK1Dpdpe0qDyXcV+imKzz5SFBeMjTOoCLCmA/UquKfHTGGFJhIyo0aT
mb2QJYhK023p5gfl4NoYAWRkwiX88Yk85a1YNi7KMDvaXOi6hbvx5LwCBKQ8ZFqVWDYehGrRoJ3S
hCsgsD4IDxQlWsKyaFnS6j4GMvoUKZWstknW8vUToikJnz8qRTY39rp+2IFOU4etkr4zJYEgsF3N
nUY2DBDdYU4iLqdfOZK05p8yTmGRUIPKwQsnRsqJPol4JZosjkLLZb9HgdZ3eAK2Bxeal22beO9H
0YL73/M9w0BaN7V64lldPBOrvfUM/zlJKv0f8tyoaSzSF4mmYOUcqWpfvc7yA4UGzqKTXvVg91iI
3JUPgEg8/deSujVA2v69t/iCpQgnTfwDp0fuHi/563j3rFU/quhJejGfW5kajeS33UbXDI5gUgs2
qSQETB+uDoewhdVy95H1pZ1vDcXq+FCme18qufRIuTteTfYI+bbHeLBp/PfwWk7a5ox50BI+ieH5
yPZ2nw6w+J0n49ce+tw8r4lgXINZ4nJWMGV3qRF2IZw61gmHa/xIQbPxPyso2LekdsRHDvHixRGf
RqUD0fNcp/sww4n8vt8NVq39RrNbf+we08O2BRtou7kaKncRlaZ5ChcZbqLXgoSUy9F/Bc0uA1Xk
BULsbL0O19bX51Nt0Y1oK/ZvrsHclwB9pzyu9IlmJEHpUDzhQapsjNo9j9d9UYwtsajGB8OID6tz
ruULIUdW7o8sSecHNZhBsC5Js3JFkLxmrlK7lfihINjqaNxe+M7n68KIeD7GSR05VHJyQOuliazI
KAadgR4xj3K9Fsy9awoLMc86FLmC7hpYGogqW+lZVkpE/IrGsvQ1u9cLoNtk2ozjhai5eM7/rkFu
kkj6baP5LO+lfek00gy5Lby367GygaDvLW+I4PwJNcGYeWGld+Rg3MhSqnjfHasdNr8EG6S6n8ug
tBZZ2DHrCEOWfBO+eElJ3J8K6djI9KGX7OgVh+vMfhCpx1TQIpQUozbMvGIdJRTlMe6d4gzA9BQy
MUplpkfhlLhSbijbZFABAHrsRO9340/YeTrf4cshC+CKRCUOFARnG7nBxvzt3j+uf+N02e9XnYl7
z/LX72bKVucDmGYVUOq0XDywpobZCuiJSYcPLRtQ7K/wua7QU4UEjVLjZkOpQiXowqefYV1Xrc9/
P4g5Udzi1hi1WgXH8sxp6D14IhM2ypcAfdxuldxbVHMKs2KaWlpuYJ3hc/9cHXwiJJtE2OGIW6Hu
Zpg11uH2NlLI4VF32yfGjLAtC0l+m9zgqJkboul4XZP/XFoGiwWhKeLCdO8j3mjDd30mknJrzICT
adbZWn1txs1lsiknWvs6v5Bp0fTaGazSxABTdLoSlne2Vl1BVvaSP9XgWJf+nzm5KBilQWtZ3Yur
yKH1nt+x77GEbGWErFnHdm2U/3o9vrtiNPnKfImKDHf2uyyNKtgLkiaTZOqcdrZR7t29BVCG5lfi
cbzapB+c+z8eG3w/YJkMD/kG218NBUMrYa+XJizQLHXCRIG8u927S62faGFjNJcHIDO9fA09OgVQ
dQJjPw1zDoN8FBwl4AeaQipsXdVEvthhx6hsysjTMVaiK9Eqoxj1nAKguwPKtQJ4kMuW91CPjXCA
+XiPMPuF9EP8dXdSE70+JmTC40HUQodZmZmoBbyABY8dWzs1RvkDQ24LO5ibdOl6vC6cIsvfgbeV
3SOAws7U2E20hU+xaIkrSTS6ni1P/Ygx8OUYyJoWsJbjWSfJOU4HgSiLuxOEIGvm3WGYyNhePrnx
5e8izwhRqar5U4IY6DAI766ZOMf6t1LEd3qYyqWMDGjhZG6PPAVFzX4voQr8sLcO172MoEX/xnku
an5GKV5RrlXm7lmNBpJrdu9WSGeYKhRf0JxljwmXPtMh7zSLpFNT+J845H/h4SRi3piftBEkfxJj
KX+7KmKrtBTOnnylY+DmxtVlc44MysNtxdvZzXJb145609E40jXncwgMGt5Rg58gUwtzHNdWFg8F
+/bCoJsayvtyGByjQCN+6Igdjbhz1ONfhcFDTCr1vkCsqXybhAPwImHNlzPFXpG/dAEvAilmbxKh
T9HTZxLaYNJXb4ZopW8Ul9o6Ct68ouxrPcazn3MFTeYulkWeT83mazh6+4rENoFFmwoV70ZCQp7i
lQQO1t+XLg43f7TktI8UssiTgFdStenKksGsA7qQ9RBxKyJtqzmYyNK8ldcAPfGZKGi7JUVfwnr9
Ez+k3s/8SXUGzu9i9DQ4qxKlAZLjRoCvld0B6ba8MWtN7sLJrE6g+y739jfedwKV7eEYSTSF9Tmy
6+dfKsiOKS3rEqeQuWrYv4rbiDZmFZHoFMm/OuT3Hb0BDpGE/7OvhsbtUauis/3lMFdh4w7SMnDL
hQCPtS6wQo5Yev3lOlY0YCZGO96Q89bDfGlUUzHQUrntNIDWkYZQUg1IZbt2QmdykdrrStnOP8Av
gUEq7522leTHUXQsB9f/m0e+Skuq1Mnu1fmmWHRcIKL6RjxjbHVmyEoYdKSyYtgRbKHj+J9q/fim
YwdCVNfiVL+KVmLv2IE8z7utm2YTAspwXT9QKCYS9Zq7GctIfUY1zrNEw0MVvlGc1Vo+da9j7Q3F
w90jFMq1TDVJXU9u6K5iQDyXBwIMBaKS2BLSsB0Rad5zS1y8XthKwkmpDfz/Or/PNnY1F1L3OqC5
kih4w2vNb3WuKSvyqliCB0cubEf+nFoFS+5SdvD3Sjls9dHsynKt49HDMX6PFg6WzY5NUC+82WCq
fXbWTiixbRsgtoTBbQ5mvz+7xrTSIQwKS9V32PfYdVKFW/OJcFKw3TByBsVOe4D73YHLdrf+j68q
1UzzoVi0I+90qRqg/FvK9tZkwFMw9+iLXXxI0r3oJG21vp6Ihn0KfjVs7mRtx0jOppddsA/Kb7QT
oDzeKvc0p9dR6VUOPW5LMeg82EaNDqz/9/633cHlhrVHValkaaLjvS1dm+Mr96UUPPr/LVK64upR
uPqGSqcVFeLY9SFEF5bnTFqT71x1DeRWTYGo8OOxDYdgIR6frO4XDXI6MywY+m5mKtDSuQAZd/Vw
HC6PrEAcoqYH5y/jhpmjW2bZmfUT9V8Ed3Hz/AqYkWkxIJjnqEPBASm8ATeKhyTHSImdYGdJaUSv
BBp84geBF1C1RidzzYiI2tuDQ55K2jPvLFOwQZ8ImgpcSA8Duti1HLeMvGO89dYwuGgXsG9Q3YEB
uKB58KbUJanbg4o735EJ2e0go/YPQ19qe9huo/Mq+zNUuPD10RZ+3XUKqb77Pn2tdQ44CJK+chel
wDEIPDvi9WMOCZKCCPC6huEG36sJPKSpKxDsvgNfvWzRaN0+ke9hqX6cEBu659LopuMYUryxmPGl
lyiN1oROa2wwLS7pnn19Aojx2hzIzUBTpbYdYaBFi0CqzNNKlq6aVWsXGIFuKQveUligAkQr7Zu0
Vba5JzUncGQWTXY1GNI51Po9trzzxvNozh/WpgV7q+mYOCaDq9HtTmfLZGOxTmYTr4hwuEDHpwz1
quzHtYBwUu4k+hbT9lEn3BO5nnFAia02CRob2bKC4OVOX4q68GUNU4PWifTKFcYZN5chXnWA+Q3i
p7UCQNd5Z4+W9F2pnagYWju5TYFm2LQPLDjOvpSg1RawQUC1NwvfflXLg+N+twDIC/ABGC4Ml7jc
6wGjwJi7yhiluULXwjQn5dPQTg1pmTWswUx7WP/zzQXSHOsAx1WlcTBMtW+N0BQtHfIHJFmP3h0B
s2QEpn9EdVwys6XDy/qhw5cb3KQVUCo5OPmrgJXvgTJy/LK0jsMouqAro9m+zMxN/mEDwZh1xbyl
hFqXX2I+ms221u2KHnLDfdjMBgMrcziY20irzlOEYmct3FMhQ3zBPpCg5m1KgMPyySEvd2xOAoSy
uwSn9KNQZdZLogTXKQmlpei45z7TCJcpgo5Baua3+FWsrB/jQRLSomF2rsFotvYUVtG0cFEjfkiz
VKXSI7VSdsvaFsk3zRwdm1OZFitkRgvkFdGuE+kh+/4fkPXSHm0xYw0VBq7dnfupKGfSO/fbLW65
ulczdQL3NGh7X9DiSV3JLcxsCsoz0Q48VWPAWmKHuasIUoPgX7vLItqh3Ite6ti2rsWKMK9YqHQn
CMJSPDQ3ED3Kp79MHd5d7GqR+czj/uQX0jQkj+nWj4sy4wrNnlyNTxtY10adPBuIGOik+0X6T2cn
UC/221jM8zZ1zsvz8Rph4LG7DGDnh+tSLEnt3PE2OeUnDGsGC+6BK5MxcbAD73YA4IrvzI/B6gLt
4+i0Oagan7DkBiC5hKGj5OBjbwTQeP7kpg7bjnnrF3S7+xHOgn5Ar83qWa3S1tBLl1oHyJAxmDju
HHUuCglLQJpXc//a/0V1hblZbDxJpYC+KE7wlqJ4+H+SfsUY2kdfHlATS4QLJ8vqbXQKPdIZlFmq
gWUO54SMPtota1E9hU/HNRCg41hCsJIvgpECFNzJndC40IpOQq+2xQmLR2fFY8sRsf15b2E8vJrz
DFuteeI6uuGQq358ZkEfP01dvZQ27A7T9pa71qkKy6EAvarzXND1KERkhwcUqsATVgj593Rx04d+
gJt7TpphcKvOVXje4uk8rCVsXVQFzsrZS6340I8GzPq2XJEQu5VWIxQJPbZrTyT3V2vJrs4zhkiP
a1IQZB8LYTxCRTCVZzE//zhUKS+aeRU+7N/blNSlKaVx/OEWJuEMPsFW6XTBT1Z3h5Qh9pLHBxxt
d1S5klqe3hnireQZHthQcvKcZxJ5kSzeypc5ftcGD6Rjl7RkE9YFontWMotm/fcLbbq3cdKhkD75
Fk1WP59Z4W1Szu7GJoU4MzR9qNmYoO26JBZqDpDXCNIrtMnHxAOC45bTKFVwvCVZflf5TZq1eCxy
KFPU+cUfNsi6wel3rez1LE9Sm+V7SlHl6F/tePiKl42W4aMyAtKXsm/DAccEjXmu0tYEIBWtYV0Z
OIY8os/haUdwVlTQztUTuMiz1El4en05P5Z/AyzLfj1S29WSs4NYvjEKZxKo9Zn3hs5clBYtDZct
uE3VuhL6u9RARsvv+twmANyyqAIwboX0C7+Ij13TGdmv69/DWNzRJVN4peIYqF7cQkGYQCp9vF0n
F0u0eBOpP/cEtQd5S/gxW1uvT9GjvPdC3j2+K1b7EJ1aeDe60IvLn3gEqF4fTOZjYOUaVjjHbukx
m3W6qqtwlHhlGe4/PJ6ljvrFGtpZlUbnMwff8GhWg90NKs78yaaTcsrcFD0e00MSLV4TMW6jc++7
bYllc/s4/PWhbtyBblcVuGyEDQIvo3KtVJoqno2rN8pCbgmTYF+iKvq+JdXUWbuWSHLGAHVfxMd7
eWIIY+wJ7oY8t4c2/Ut73AYCGGR7Ttbb55/p0ljqho1Qxm8353Q9nvzL56yQYdu/7/ukx1HGjnVw
21evqeGvB5sGrZtNDc2EmYMVWabqIq9VPhasN969ZBNefDXy+f1IN1dfD6zN1y6NuN1pGBVGyHmD
pxn/KZLrYPN7jTzfYjlpnxQe9PX68iM4rNqxjOV4KxyDvS9eZjbeZb6J/1iRZDWXcjanONOg9iHg
K8601Ccdudfjg4pOvmsmBxZseDHhnZh4N0lqzgcddF1q/oiH8YQCr1W4XdjhcLfqH+LVvTkDNB1V
1ys2Hzz9ZLm2xnzVK4zNEQRqycgNeDPXQ9E9aqF8JeyUpQlEpO9T5CZlJZD5Ofqu+wnqP+Y5tqZj
W/b+PCJamZgne6pA42QOmyAes5T0rRC019hvLXopRXsmzeYrEKmlwiUvNCQaSS+ou9EZQt3eFsEB
d6Tarmn6lr0E/cah9MH0sQgUIdxqaaDwfbmDo7QsFj1gBTq+oysxFkLx7z/GgbL5bBdtiRQHoZG8
aHfrOk0FAo0ekEQlEbzZK58VlvvydhoQcQcusgN79oQTc4vYab/LqohB5T+OoxkZYrxbPQjKS1Ho
hKbbadhq/hwxyVnzpzz6bsKg5M7V3TYOeOmM6LaGjgESgGUD1mlWIxQeKR7rmH92dE1kfFWbwYbq
7GwauERDqggADmgkNg1aXYs3M1rtXhn8jeJjIjjNZLpZ1/nMelx/Eo9jDXO1ttcRWwWlOgmC1qxe
8JrnH74Nuy4cc58o2fAlQ6CVOm7cmQgTjZbdmkxRZ/y1JVepI4eH5yZokywrPpFk2HZcqVJzc8zG
XDH8j2VnDuhvVXVTTzQ61Vc8GuAhOQOAnc4fvCYi6a9QjkPBOX2nsrwoaE8R4u7VaW+/GNraFjnB
CLzMP+wGoHGYjQkUV2Z/EsO92LSl1ekoV4aBu95/mbmQsp9Jvthtvy/Z0E1PjxRLdoIw1NGmJKvX
BIUrWhqKk5qECxuy9uCEbxxB0VbAFQJpDlGXGqA4JqaR3yXt39lmAxRGg02qVp0yhCyU7ZgLpFmv
5E0uYhkv4tMB7UD8mARxvP8xNY1kT2nedHtqcNetY2Vt+VhIzLkFGRI5ve2uZj5cmcFA2a1W/76D
Ael72vaWLzMZwjZyj+EXp/+ZiVkspcfv8X3BOplJkOiun2DGnqISK0IQba026PR7bXG+4v4wEhuU
ehmAP/hn7Kv/v8wU11IqWQbxUz75oft9JinkhzuUyw1TaeJWk37OyLdOLWAAsNRsCAyOGWnWMZ0S
UFCCJTdv5gvENChMqXKeJi3qB0THru+EEqoV6/PUZFOmoHQf2B4kXPrFG+PkGeOBY7bDeJODbeTF
8xvbBpEr8vh5R6ZWVnwKWtw8joJJZwr7h7r+xfeoScUjVakIOjFfshzQEET13gNlDdoBNe5A59fP
EobRwsJHvMMzj5RcQY35LFOAQKgpkpbm3bu2mnHLqLO5D99v2B04KoaJDy4tkuYOkyH001hw0LXo
5m4DoVxpkB/xmlhXIr7d+ZLVyrwtwGk4BvXzV3swkMaDM3Gdcw3B0x8eu9agOIS4V5vcrlMzM8ia
Difx+rUi9tN70mwrej2OpfJW2t3/96su5+GYj3eg5WQm7FphIExoQMWuYHgUTQRbZxkRmRjZi3o9
2vtXKeJPirDoAkxGBKwboP1AaSZX4BKWpf5tP9dpi6PouHdl6/4F1kd8Zmoz8TRxwgUuQcfkAU9u
Yn8syoTFdlrFxzZivl0GcBiU/YXAqqYRjZahfOja4KeCZoCxMeHUI9HbJk5oGRdISoFruFEodoqA
Dw37z54PXGQhHW8KKx7PRcqnmIU6KjzCzSHWkZ0N30SdTr6fEpXiai6OzOztltgsUFK+VNiXHSJx
6LLyUA+QpZi2PlfhKOG8ia4fTU/dJRf6VSVlUqMt+0PTIMc3meM7MpWOsVB8mCWdLDSRoT3BoyTI
KdaDZGyGGyX6GDb1d+hgevFz1IB2n9l8qsmjBTI6GVjoX/Bv8XUzocWFuWEjlViYxu332TEsMpZD
ba/uet7Sh19aiNI60sHbkamA1cWdHeIiE6DrFnBXTFvp47POuO+7W1scWKljNZhV9Ws74mR3NNo2
hzRsUx2i1efkSSkYwUlyehu4tDDVuOsuLvgcKyY7HKpU4DQ5K4neSVXWs9Xf9qXFun1sMX2qW2n4
luh2Cod9MoFLEfd3xD8yMI4Q0hIWFYiwyyHVKkZHgR+MgrT2oswZfgRj7j4wH683Wsvh8dFeV72R
MyTAOjSundej6Ue0y2RERCkh9OE6fAvYjuY51mwmmXWPgbWywfgIZ+8EM1RnKCU0QrzOoUV9Azdp
BAYp9P8qEyoAC4vIEDJJTDwRTTTcPF891h365tzlaFTJ8uwbT3DEZdos2y8IoOZxGXbXgaVX73i2
+bd0+SGjldXKBATA6WvLcYi0Fcb/7lChzTKlkmmW8OtoL9iHRlat7UskZMB6VgvRhh4p4QFR762U
XfK95HtlQ/WwcizbxgC4Oc1G3PSxqf81tl8rHdiGl00I7Apccvc+W5SM1CyL/UGqnDTGJ+QPPaoX
8ZSwllYpkxuRRKvuSt8Z0odQJG8qrQ+5GiC7JaWP02oY2h1uEzWgvnCJ9v+cagl8u+4t353Hiknf
YSYCDh9jHou5wyWE1B+4oF1J1RCtR8bXG+1cmk9vFOYl3bg14QGkAMuigk4rPDp2oFHTzf6Y9tcX
b8RVIVJ+491VETgTtTHtNwhux5GvxyYt3ZitHJc/oxfQEbh16FOulMZOfq74V915SpLGbIYbNCwZ
NBh8J9nwWMVfmLzFHRcDqFZg8nvJh/+C5y9LU5bDWGybJPT4yelR0ZoI5l6DtOVPPEyzSuZ7aDXJ
NdN9MpBjYxwj32jQLYAeYyE/RXqhP6l3fldJg1pWWsmF1UVVn7mViHu85ix64pG9Nwdo4WmxmsFW
JRD0JMpIYL2fvixV3r/Cqt1NaUUuxeL3E7Dnqu6HfwonXsBjsLVFKVnk0CPvc2nUi7/oopSYd5jN
oe3n9/W7bkmlKLKCQXMHkdDDVKh0+e5YF5iN8Z0Ts9dWHebqCNbSA+x+tzP66mPLK2Ez5itH0W0I
m13WpF7VBLZfhkDjgVrnjk5uxKsByuxKHTle4HzUm9RmNhurj/XqiS8HbK+CoYyih064b76hEX6X
3CPTL/y+L123hJs+JX3VFDp9XOBuacXMGnmlTEmAxFOqvYpjmHNYFFrXrxB/e56++yrou8sMZxBz
SS4kukbkBLK6fMd9neQv8sea6QJE2GJ8oxyk3hJwJ1o6yI/7iQMSGQX+e7Q21PKeGuPDaeVjWala
zYJiyx4BLDjhKJ9ALrmOv721QtF1lJim9YJ7U7Mj/SEKfSLxDhJkO3s7UfAD495zb9IOHkpv1TgY
f/Q7X+AeZPtYU4B06qXbUyE2tdwFMDtes7GxDynjDLsrrAXk4H9jf0clo36oEmkr6Pq6DonTwBl7
YlrgobiB7wyRrbVYT8x1AdzYP+bZgOhiKKiXHkHOg+W5p8WMJw0hk9yfXaQmq9qrdFg/zpXZXONY
QdsUUVLeWq23gPyzVw7KssMfDxf7A2U/SdxDgs/iLxFdIbwvRUf0Mp8vMJRl4Z8ZMpVqAfKt/XAo
i5iwblFr26n3JedWgiSzj6g79JcwHCoB7pv8Sm3OkK8gcUqyu2oiESs+CSIZHdxVwggZk4olEHwn
1QFFu66cF4Le43z7447nXW9zwpfHx2BV++7YPqJuPqUzIqUyy/NaeACXkqTefavKhMcy8e068Olu
1z5akzpKCO5FoCwO/0gq1+UG/zorCJsCGqq6USyVwbrqKGD+4TqC/8+FG/k4STLVXQ/zKXqiiQnA
0dDgVRG5CoZQemLu/j4mletRSqzLIOeFT7FY7fnHh2FBS+dT6UHiW9E9434e+DH5DwUdgwmhxgo2
o8sTLG/0cGJePmPMnx8tWI+bWe8it3ddUQO14K9ywpL3RkbuCSRRU84INe04TGGE0HByeGN2Yz/1
ulb7fiQtVoEjaVkwcpg/4/aDjIegfMrgnnr7Wrofb7c5o0AUCyOt0uE1JkagOONUYi7Phdiw44U1
iVNJ5M2QnPz2fj802A7vMr2N8bBCY+YLK1fvNIF/9iL/N7+fHTXWMDBHdM7ykG2GUb+OfalAisuG
EPf2IYWHVQYTJ3+c7N/qxbdGy+WtQn3/unXuAXMmbniHrOC6z1yIL25pMc8MN2uNKd/LJ2U4akL6
+sN9jJ9h73524vIj6/VkqyBvYpxHnSq0H7Uqcm1afOzIK6fKmfhZkndr9DDtNlbwj5yl8sgIHzst
dWmIUgsYsv7/CRHu1osD5l1BP1cJzNBvetE2oGcHqsLvOq3oZ4NAB4w5KM7da6vFPnvaH0nal1Ru
9rAOMqePFP6ZjFRbjLdmIyKzsgJ646Wfk+rfVX/ZZrqW383EWrWc4TDjc1fBRKrxvH1e8F3AzZak
5JYyvYfWxO2xAi0pEaBkPJhHudg66pV2uxNlmbaInlm5W+w+w5Zmv+C8r/UNhKC39meSM1RhaWaR
arm/KIuJcxw9wDxwE4gz9Uf/mecfi2xNS/DK7Fq1vkq8O2gwsxJBCDdyCSip0nFDdp3iGfAz+geK
Dck88sdFdNvr3E9xHypTHmcm5JEBo95/+Kg9d4b6Edh8+arXJj4sPvbR2P80q5hKQGVL3b9tlNar
fbxG+LvMJpfDu4RSFqcIpC0//pVkEMD2Sja7IJiRRSRC6zk1fL3W/mLi4N/jzZhGBWmVN04yEcRn
mbjvvWAAXnUCQPWRLGrdw5Qj79ZpRGyYjHdYTGs7panV9TImwuSZI24pJss94ahPo84hsnNqjcxF
Ca56Ge9r3kmo8KXQUskx8Egl+9S3DbCFVOz17LjhXr4KBlSeH+hypnRGOD1LHKxLb36odgrZU14X
zo9qtxikJOJunyk3vtdjQ5W12t+CU0kilKZuioY8UD6yEEMqbvyiCYcBYt+zdY2aFa/k0+cdIVy6
7PBb8ppgH6s7HjYb4eHhyPjhqAH8rS8w1uLhBNHbQvaytBfAiUjVEo/SjDoxRbXsZ0FMXYd+KAxM
L5Jkj55nS9dy6nXUZRhYD81UHMYsIlZj3sliYdUtrYiY9DXP1zqfPw1b8D7+9TKSWux1CwlUTzmc
IK2/DcnSgSliMsvmaAb+vT1xMVByfl5WY9nwePpRfQEyzfOCsyii3KCH27CMiGQZ7yoYAaZabUpV
7TopVJlbvxhAUHtbSIE0pEkC/BbE+Jk8iCZGrLw5EY9i5keWy8vhX9sEOuixKd8hwo0ycc50FrTn
uBeXOo8TQuI/vzOBPvpTh3aVQuto386N9n7EGiBfleRDVMrxrE5RMyU8UiDtz6GOy/0k0IbgQzq8
CcOfBAUSg1Pz6nIc9gqbJq4lSi+QN3FsYVLZw+cmaCjEZUYpaMbiN5nLsiOEds9XV1OgR3N7ecJs
xZj0GRECs6xygVVw8QQ4XQwDvGUil8CS7l8EQk1y7iRccNwAzKKqVG1mcw+6iocaqCY5BCdhJFZ9
WHYSP0B2Py11O8biVrbP2ByVTNlSUerVoTaxnb4FhreCVQBX8/EOzghG1l4tANwpSyo2/f+ZcKqU
inL6EGw+KjBUhtvhQCZn5FeBdRkYDChudynY/zcYOw0z09NKsakhcU143rBUmj2ypm5b6annHl9r
NmdV/9+4Ij0Mkt9yP1cNgJYb/puHQZ8jeJOfEiSzlxnyJQlXAXnu9m21LijEA+ij5Q5DIk6JF01f
WTIMzZmzF5C2ujOL1veO+kkz6RbVSa02IP4HdH3M3Xm645R8l9RsRxQ5Sd7q/vfKvIwfMFD4VMuw
d4Df9YzWC6diiKl19JsRZ1aYuK7QACANm1HWSNZrYBCc0y2Yox2pJuoFSJaI9R4RTrQXVfoUGhVS
zrEuE5PVdUWtt3Y+WYd1Pn4Rl6dEtgziYAYEVTkeDK6OGeOcsfJsjlM7xgeNIQnVIkQF+EbYhraO
JbRSlchscdNRi5/gsO8rqAyPYycUrPdo26/WS8vNf+SydJ2O1XuzRfXybHWUefTFu3nEnp3GygAd
IrhV3FXzPoyjCexg48F1YLXamg0/uCvHDaNLQOj2gOUpGTpuQUpoFEVQykf8/ZoLRsohVKr32rHc
607E/32+k2GmPZN6RhqKgdPNjGe7AemrB0tHtbTjXkjng5vbxLjsnfaZR8pCoWpnXvW0FrNsYmxh
5yiiYWKKHZGO30aLSEDwbDFUStMVU2bVZa+ngSS8c6B6aXDwgIIX8rSkLlTdPavDrvZZNdld79yN
V5fHZ9XEVUuUvum9YIfdRp6aX5gjq9H7kG0/iHQbRoW+XO2fI1XK5HQ5CxrCxaMGuvr/05Vj5PdE
8UjIEZ9ZJ/1Eyk9IJe3nOUZjvpMmg/8rFq3wSSq2vx2D9QA10sOnBG31r8PGKstQ4YAkDXZ9WQQL
pmzQLD2yCtYfYYJ0aoC2PBOQ+0i3LdWZpGdCbmzJvQ8OGzZ3LmLBiozINPWbNqmKCSLsi5otkMj6
cLuy1gj7NielZKlfK5U2jm1pcYPowQ0LPPypmczWWlGP10vm5VC475kIXiHz1nFEE/oiNRFE6XNa
ulWqq82VUTpsnDNnw6M34ZilyFtTvDcrKD8CAM1Pc3AnW6C9mFlE/Ok/LbEq2ePdOo/y3zkir9O4
rTX7PsxKJP4/ZTanjn5Qjt02gsoQpKU2cTp3oPXg/V0J+Ox26Wv7rW+BPYE+TmH4UEpR/a1vgH/a
6o+yh9kLYiyPa+XP08flNGWqDUMt9j3die53WH8F09Y6SqHMF88rcGrJah5yOOFphQXFRYe8Qti4
uC5M/OvcPbxV1DrrKmjAbS0LWYRkYQx3Rbv9jG7RuUbDA4EB6bpddJJXq9FQIN3y2PYTyEK8V2CH
MqQ7CcXVMFWSNXXqTvupi4eu3MMrwggOIasWdnAEMjqCvDn0TVr/G4mMrDOEjXfhWATEbVTy7bhq
qvrF6C73rpkIGr4H/boFwNA5bUT8akuDuQILEOz42B/mQc5Nw6Lubmr01QR9rW51k3UPg4AZWFci
xLg1RrivQxZOWTeVaUKJpZqEYeH6qZiKW/yeqxNgdp2eJ+5lsGHLZAnd7Ly7SRMQFvSj5hftQVix
kl0e43Jc+HpXAuYM4Cm5FJzdC+CqkxrRtwelAOkIzkCjDPu0gwkH6jd7S/SacqbnmmJlZJw8sShm
6oX2kIZojszwO7vRvQDShDKuD+cjHdv4u8Otm+OJpN3Z0vClPWO5xFr5PqdPAX5PkYd2pIRIR+t2
A3qXOomzvSOmTtMdeqV8sLlyBqz1WA4QYPNtgxf1mrxGseiMb4gtJ6JHrNcOXjamUxtLdrsBWhaC
lQYjz+11cieLcNnP4d3PoUul4ChxRGJHJrfNClIG0cztimU8zIa5EHFUSSi/Ic6jA77+EOInFDsp
OUOskOh3XDVsohljcliwH+3PXcPTqsaz/zilQSsV9vtJwGGN49lJ4EQX0dYV9a/lPC/QxKp5xp7N
xSHX1z0g/Is27J9huASRZ4g+kbanSo9CXGYQo43K1q7tXsiJWfY1NooEKJTwbiyabQJyI3KjOLmk
UUxNYZSfRkNFfrElZxauuWlyOd9klt9PShSodMNHK4ynly0nXugVqlimGLtWaWrkFxdLcwEBFfUM
cvb5eTeHoP6IJcXAw20esuVtb0yh6RwclDvaXuY6GHFXcFQzpRLzYTpd5bDKj459H6rekDHb4lTq
EkjdcG8UKYOoVkOG4R5eW6MtuKgAV2rHR9DGshJZ/f/st42YGukRznglFZmFS5EBnimOoiPaVjWa
de3IisD+O2EQGcX5H72j8O+6tJ0kCLjPOsDABs4J1BNZN0+2H6QQmCjQAjlKQg65UjHNkMbNo9s0
0xaE0wHCVUZJPufArP2Gehb1hUmxAlsdx3o3nDhNSlPFg1b5dHlUd+9or/zYyDJTQ5rQ+VUwMU3V
T6uiDWNpEXcG/if2wTGWYxpG1qp99tHto/SdBZwpADp/KMky5QwzJ7XEKR0FXB0sQELHZhFn/ow/
0ppZ+BUXcscsUXE/NQsFbQFvS5x4pZhjV1qh+vRBDBFm4aSZo4HS+gVIkxHy7NrzB/JgDuuwAXFv
wKR1zQvc5i8oFiMgHD6asKRATSvRDJvEpe/nAlVEI/D1xHTzzMixLcG/LvRiOmITa23/IzJ8Xlza
ki7HJ/Uwc6vUdxhC6UpM4R7rKPBycce5QuoqL+lmTVySNUKzfnAxN43lncwxyfiBH9oHZ/1MjGli
cxWzBZZMSd7ER44vCXIaaevthsuDKK+SiNOPfUQugvXZJP8XQMjfimh058MP5W8S6ZQWWyNy9z25
jWbw5Vj1shdj/zl+aMIROyhRbxlWew5PTLKJyKNpfRBc6t9YVDI9OHx+aKb++Nbxw5XbbqKb3lup
GJGruV+gqN5TqyoFEw9a9pi3OpLyvEiBQWoynO31t2+bQ9RUAQAf/HXbiYn1NMji6VJANvaIMM9H
OZG/WMT80WYK3mH+XOc3rtOQ6obGgSDB7vQKNFrl0K4MXln3MNMvKCg4A7SljntaSGB6SjNnA+or
V/ShlYsY+2DTeXX1495LitcI/oEiiOk5/zma/nzafdcmrYa+ZdlDIxmVzZ9tbnU3TOQFaNPznxY9
3YC032xlmHtP428DfFxUKfYT1VJ61YZjcTKg0rbrT/8oPgEDuSQ0wBemlTOucBOYFOfuhNdAAU0u
eazRfaS4wDWrLFU2VOb9a9wK5wc6z5Rg/UrZDWD0bsTh8sfZa+FaNAxJm51Anh3p1qw8IlG5k46h
XX3IZWKKgAbIyXzm3ECIeL4Gt3go0zmNLQHt0RGWQs0kd0/rR3rp+/rXGJVMHlpPZ+8HIZzWD7CN
jdNl/BKKGNhK8ilytx3VhxpqF8bREM5jDgmIDh5uWqLRs2BrAfngBbe6bCEdpcLjdBhoTsQWUOfy
BtM+WQfRjC/NORirsIK5NdaQ4NY9+QdkQiiFg3OS8KhTvCsoWVEw7asI8Q6VvCTrx+H6GdqbLS7L
zRhIQXaEgCPCMzxuPnaMnpWwJwrdfj4Asf+uCy7I4TgHeIYEpBAhaz749CJux0UBs6RbzXN/AOPc
iN2UGMSEA60cJY6xKpXjvS/tgMakDVjlhkXu362X744gngwS9qXpfM0rJ9vqN/r8vewzTmw8mvFn
wyWpNxPZFfGSz6QJkBg339gYgtrcVc2tJqk/ktrG+v0ei9qLP3dHMwD5yQxQdnegSKOWCmGyTG25
pcvtT9WONc+jv9SXcP/bUERK06WsrmCFY/igEWCmIedRfWhOr3xob6JTfpd2M5cQ/V42y91QZMKy
uP09zZKrHcx81hBkzKlQ10UG32jlyleYN1ZDebRvTHebrfCIq3fxxGZ16B7HvVoOkkzzfQ1n77DQ
PLkzCrjvLzxNl0Hlq8kAtbGgu7ikiXqkK1DR7upgchV6mZ5iBi64g/EN2rM7CHJYrwTVgHoBBbvD
zGVNVvmYNCKPJTfURh+bEHtPg48Y5NtMi2X6pTHyIOZL5+kz/nuoA86fLaOykIbB0s2il8mwDilt
aNo9Wyz1znkkwVBPiCYQeutq8gZH9ZY3E7Ljt6MW6MCGFUfZ7Y0tV8EPlW4WpVjwmIrrW6E0vMdZ
Cf9Z3B4FQYITjTqvY17NxCP1Y/e1K1gBRwy4ki/eGjezCVD5s+nS2bA4OZlfEAEWkmTPxxVmaNRi
ugaqguZsblWG5IRXrr0H+A+iTf1GMIsjJpanravhHDlDg5xmo3p22WeXjCCq7wns6eV1GxC2AHOv
zrXXhkQ1QqbPiRQZjq4OGQ0MCH7VE5guwezJcK7ttNf/GkDI4d2fRwYazXmKTukjqqUB8zKPi03+
4zWrta8LeMet716SrX2XdyV1bKeVXeb5BWhG9cFaUg7aPOCFMNr42Ql+Avz0ENWuz15/FdZLulgI
obUKyyY2vDq+wCI+LsbxBwgo+t2C85cL0LTjjlR6MLXitSBHQTsHs2jiH0uVpzONDg7S7w42xryc
inWKayW8dDqvwr5SDsL9Vk3U3Uur+1XJ5UEJM1wdUjOoORwa7rNCofXcwgNE2pME3fY70u+G7QPq
weuZGPt6W2zcc9iANn2NjxyLK64mPYbeXLtJ5Mfl1JLYsie424Xi6LnczLnOZlvt/ldvdcy86HIe
aCswAopbJWDnBho9ul+RV7pPCUk0ocXSFqQ8U8mxUQZQLo5vZJ2oPKn7jILnKEtjqh65tq9BvukY
5UO7Bs5IhDSARzycjajty9v1YVd2GATpnWZ4B7qQcXVlNcgI3WltL5LmTDAP1o3xiz6QdKahnHoX
jLZWfGsGnYKtA2zu/tqlXptTqlNIAXG2Grz+jB9CUQ191gebQbo9jlCYcNPkdmgAGafDuf91GG/p
LayDomrSjGhSxcVm4o8UZQpswNJGGnmVCVMSyVMSApdzVccmBnHWfhfclQyRdjKh0PQfTPv+royE
+HqVV7HSX+RSxClsrzH4S7MdSvKa7cfQZZ3117TDmnZqp2N/Ujx39elc7ri09CSCVcSjby1Ir5je
qnHeM24iAcarL5YLqCIquT8JJL/9ktfaKzDhhHgbm9bZdFI2x2g4rejBTWqTGv9WJawSqEd5xGxG
NCWyT+8eeuWR8tfS9ciAifMp+GSMCYWLdwH2PGaGKH85FhGIbKNAV/+jJ11NbQn4k0NYEVbIg1gC
W4i5+0zxt2mbOgTt6G2cjoBPZ+d1TB+I0gTknsGROU0si04iuute5kG4qew+51CRwi2SvgESqnrC
ipbsmMnHf0Z3weh3A+R6ii7870YEFeaXthijYGbBTDKU039lDsxgzxolNAvyXvCLt2flWhbYYiqL
nShhm9vQZs9xj5F/SyCUP5o70VqAFIX4V0blqntCCXT39EREov7iclvm0Mqd9+bYWyhIkgN+vk9h
5fZ74eMOjlThB01nHYRMYVuxLsQl3yTlXGJFnAcUcuwxY6u/s/bwq0pky2N4/KhveqMmPHicnTyI
FCGSkj327Gu8ad0HdzE4o2SjbF1FUDqUyEdbcaarIjhbaQoFrcHjYDV7+GrJWwwOC94+0M65PF2j
4OuKqU+llHthndg9m7suUWofPGdKzhZb70m98SkIf3qbhN1V9I4Evj4+qDDrk4+IF5dqooKZDOjo
ZsM9oy3RDoJn2hndg91PRq6sTXYwD5S6aglwcyJJfcifT5hFUyx/daivLv30XZ8xTzuu5JoLsyA+
8hf+dDlBob+yh23G2YsC92AgeowLOq/zZ9gZbzHkpp4KEFLxMqbIp5zZv5aDqyk8SdQIGvMxuTPa
yENyLOF4hdYB83sYuFmAFutCdyCon7z0zLhIEabRblbq2HzMoKeQE9PlfqIhEHR1h3/JWsV6zFbA
r5AYJgBgNpYXr/0t9hfrBeyVPozRITaeDO1gj0gqtcKcruI+8htEcm71GGS4xAn5JO+IItBvwdqI
W4d9Oqg3ktqwNuC+bwPEPacT/2JNaT5g9MPI1HQ6hwMsHu7WcGYKin6wPT7fpeEpsaaY0P4+pT4m
+6Zyl1Z+56ReqEuSuJt/JfvD7LQxO8rPnUGsAM4+fc2/KDnqSTxIbIAxiz5zRdn1htWp+qHH2wwA
Ef+aaGYjRXZYQdIwj7ePccMPST2VeWG5zVnZxJ9TECt2XA78NmAVjlQqjGKb9wNyJs03JbOjAszL
KB3MtW4rCyrD5QBpSPMa5g6LvePtOxminfIa+sIiBP9BPIxKXeYlB4Z0IsfDe4GM05uAwts+4rBR
7tLbH8Y38+jiQQsEo1IW0gWfPkaYqC3/a0i/Hj9fPXkk0ReyonYeLx4h1cFmBwhrR0nNXseA+7Gy
J2r6WwUwcoct0btH8O3YOtcF62wM4LSchoaunoFcNkTkdnZVuo8eGrXnyz+kWsThH4Azhxel/GkM
XGp3PB9Ayo4RuoiLBQY2euPLyxr3UEt5U7ClwIVIuVWKvbIclcnBiWCwwI7lsN4vz3Y+Ro/9rYPI
0MS9zPsS5IA7j6MEnxB3XXJlqNRj7nlGXXUmjH595QYsVlR1QrJei+MiHVPxL/EhuVKHvvj6vbW4
w3AWsxniNtm0fuHRS/x9AVU/YFEnGDcvdtM1ClbSruOH0uICTuPbsL31PxPF8crlBZ8EvagkOqV5
YM4+CxUs0Y1lAIQ5uNGAgPZYPUCOz7O+8V4jU/+D2b0t7zwCoFc64G3FHoTw5VXr5MBieYl8arOq
eOC6oDbuSo7uqTfAPRDcK/UA5FMnk8c4JlGxCpVElIMpuySbs3GemL6PHPDG0s5Gd1DrjusSljD1
4j97ha1zFrrJVQjbSLc/rIUTgfR+J1/omnY7zpY/3Q7/OPbyMpjD2Mj4cBY8I9CLNUgwUYMehA3/
N0cAVHo97yGxmWKykXaWV/ruA3k2t1ihXM9l43HwR+7lsPJ1vydDTfZvoAMgmBypyeaJdOUHGlrx
TDtoSPhxGddJIbUNBI8B/hHWoCxemjm7Tt8aes6DJziVtl62lC2GWG4uYATjyZKMvcjik9/y/cC+
h20nSmGjwWPoYATj/wmJS9S0UR7ghvF9w+jbGaaqZOWygyHU9/f5Herv9Tes1eU/Q8Mcmo9/F+va
XCP3H366NwDF0jd9N76mkrhkV1QFLEvE6TpNdz3vSA9V1GkQDiQ81JqPIg0LgD4LT2c2XOu2zT7K
WjRgQ5I780BltRw49MCxQIjRAKSvzydSUmATZ65P725LlZHlhs7KqkVxBX6QtcX6/eMa8Iqyv8he
tgV+oDFMTYzIzOk8kmIPYW66qlWydqhXgjDZBcwWD7B6u4trKh372gXh53W8MhLT5B3uoY6h+7TX
SjHg/lvwtqBAeNZz6dKd/4KmKUYQiwZuCSxdfCSi3AqF+5Ovoc40gc/GRkDLzRJ6Y76sxyjZPMg7
eOzCZyThJP5zPDMOF/WWIau0GgLR/1aFqv9LNWVGJljdXEsM+5l1EKsXug0gchPGcObrMIXxpKDj
cfWvD5SJLasHntUKEAO7f1JbPZfNkBNl3SA3MkvUKUdefPHcUN6t0k4BnHQJXzFXbkbKM8CUnXNX
tXYfu7lxW8RDJv43k01TFJlEQHqCZvUfZzOLJxIIX/tmgkDPbrK6BZ0yhRnDZCQxMLXArAly57ao
v0vitlkViwVI5G75OkqqkkDPcGqDs0nfzaz3He6+idJZVhp7ZnAwjHLWP4WTCR437oSviMDgtV3l
z/jCqYWA8Ho2VTlXWbCJ9XzLeuhFRLu6ds1bUaE4xorKUJ8DreTv7N/2UoqPGJCRQv7WHQCYF41W
RNUDCrAhf8+RfK3lgqDyXHPHfXso/wLYj3u+nh+iExHWr0y48hRKp0QEEB9BKVXTBXkzvURzVMi2
flAc/yTm9aj+jxz+UD1474xY/GgyzKuYWaEodWYiJdEGRnGfF8yvH+dd6BI23nH2YCqUtxEmnPUk
ZeJvFmeB4jDgDftXIbEu2nx29fJSrG1v8z+GyJn/rbjPpBEK0sTh5r4YaPz2rt7CdF1YPhcPNN2X
zAxeD5CpHPki8zGH1I1y7/beZef7ySrbQPT1dcWkqwRydF3lF8k0f+zD9/krbbuHfiS4GcTOozB0
Y1gS5ISozh12phsb9Oe2xC05kXAewz3JZNBjIoPDG9ZnrW/jrswedh3+eoRu/k6V8rrn6ICTVkt2
xJp+ArnpQoXZMFVz17Pb/RgogrsW8Gbvyqw9oXQxake7ldf1pU+OI/z/GYtyc8A/UOC67bCxojaI
Fsn7CVg8Cl/dpfmmNFplq4X5M8JpMggn6RGbbtITy1C1Rl5A/oUI9H51oRAxFFvHG35zjx5+5s/h
bU5H3P2KwXXo0vgahxRUs+6Cd4j0BBYfhaUXJcBKxoLzych3Rnr3vUDdx1OuKLVeD6GMePw3R7l1
VPZZhQiUPDM1sXWwa3JGKEE1EV0aRF55ql4EEKbBd+98AQFe8H1RI6I/1Z+SuqoLVBPvvsiKhxoE
U2s33IEZ9XP7hiARmCsYgiSf8wIg+D885w8WdtCqs64D8dJOKkXUo85tpMn5Ma0CtH4+yeGKiX4a
EDreIQ2M3LzxrKCuJYBWUgl5GYxv1oAWCudsO6h0tj2ik4eHptFXKpmf5NIYcH1Ckqb1jjxGDA+I
pCtQ44qXvh5zZuk+UaNgOB/frRQbefHMJu735P/iqLQTed8Wwbk6pNabRFjN8lhUAk5KIhgt9xGP
5iJf7tJ+jfUwJD/77fR75Y31OazqLDaXVye9cc6U87LQQNeOaVD0L3vhh1LI5/NJDXQz89JQcai8
ZPh4uFvJ6W5IQnMww5Xz/jrbYGlx7sRYlu+w03ps97u0xnoGoDmo+Fmhn9ADmiUsbmS08StLnM+u
nbpyzEnevnKhr8GlV8JS/R9tUroE8Be+8QuPeW1+MEfoTkp0zT9HdvCd2tphdcIbV+K3YqSFtbRd
FDTBlrOYYVUSwBb3ZbQt936TwEhshj6rDPhbKX3oOqZRVZwaxU/hbHDFGZ2bDJEsDPBKwNinehfX
QJsdLwXR7NAw80/axD6MN1JVfUmnmiuRhqNrfLSaHJXImsqmp+UxdT4y3Xbxpx0pe4StS5W1O3Cl
I9LiW94Sgsh6y4aPpWPyAkk1Rqib9zC2bkKrEFvsfqYBV2CbRKCf7M5vFtBpxz5IaZh+uldiTIOp
2+ELHyBctGEnvja+JBRkTowlJP1G2K2pIH368MgoP1xIv4bnBS0QWbi/VpYNDhSl4nu1/+CpBxLn
2vBU4bJSsk6p5NR+i0KtGGsH0/9mSPwUgoy3bIei8dnuF11MuZzMxiZPZN/qGBLqV42sWCcKS57X
KhEex/5QQysjqDJ79tzGh4JFrTFs2D/ex58asqEditPFRSBczV3E7g+89sj2bePQB7JZpz2XW37r
6hT56HO63P4OKel8OzdoSIsHA+ypGoo8NcYAPVijvdF3qPDlW6IIWstw2ZkxevTySZE8gKG4jshU
8kvaNbPL0V0fws1pQtr+i4CIiXtQIF7Uu32ToCm9J21qxEY/HVtkcIhKxHA6btm/1h6wovN8YVL2
jpDNsGAGiUn94aOnvpyU/nJaB2SCbdNY/rUlvGbgZjjLH+yjHaYSM780LzGsF6uMhuPGu47v+vaq
Kx8OM2Pm2tWFLhuwESMd5jbY4S3CLeNTy+QgNQ/6ic0yxYplUXyR8D7jouBaybFkAzz+rYBv/42s
nWtTDDVFwAmCxOl3ssZGAvA8+a0Hvd+qT4n2dLtpTwoFTCqO5bRYP6j2c5dr+sssZUjqezgyNfLT
yxWdbVxATJtKUdJrISFI87qDW81IxY2KfzNowPZUTsc+vQmFKkMpZRwZBH6rRTIqHASiWQ88JNt4
Jf1p2pW5Q5G6rZ7lcxLTY8k2IWr8QKkpHopgc8JbDnnchow2H/2cG7Ys8ark3ri4I0IEjY8USwr9
7n8MRbXYGAoFDzeKCW51LuzHUJKuuod6+ZXV2Czr8bNjvBOuEfQCg1Odq3TSTDCG07iXhjz0uPmi
XTr4erx6UM33QJskA1H2ny6oekkfJS+Aq7UpsP8wpIEGvLsLxHymY/xzYtt3ko8lWIQegqpeBdjq
4TlOMyvd86qD+RKd8Oe43AnfPi6J30NbQxiZR3Ejop/xJsxsz/PCaID5+sFv7yoQ+7X6mSJnf5vB
wOaYuNWOOuB7aorlg7lLue7+VcgPwRVbH1Qe6svR02k57T9lndtfLIYK4b/4TWdLDRK1PIQW+x/0
avHpVq45Sltg0ncuqbfVVSvhkIYecjcZQYjPWfKBgorhojdt3VuR0ssc20qqpPdGCagJWMFGCM7P
tJhxAjumAkinF1aA4JgLDyr3BTDfNcROuFIkZBz08qXa+m6LZu9cMUR1qLTWtUcU8v4aGstrEYDy
ylLGTpseISHF++2IkEDWjJSu67xKW8I24tGREkiusbhzqyPJDb4GIkSlavgxq3lX4mWNvmw3gXdA
qItaqi5LBwJW1ni+8GdOp4BqItzdQxnRxGj40iytFvVIU4Obzkpv+UlfQ+D0bagxsj+1GgtpUyqb
d9Vdw65PQZhLHQTlEd/SKimqf1KEa01wQuIHNNVf5yZmfxz/cwuPjhPr4b0R/ihsmOJ+7NCyyIu4
qaM2+syvw24GHQQMp1MRaXLSowCTcVYG/DJbJmZO52GtWYMBBjDHZINj7s8SbsUaxulPX3u+9ZSw
aHL+9hzs9DHy9ftUIogTdoMHXjFTQRNynnCh5SUkZucfK5iPVW+cddLyat5NNhL8quBrrjQUXbMS
7By4oDKOrUFMeChSz0+0TARaT5HW5W0ahdEgaOtqdJFTuWASlKBAcMow8R7kcYftdIx+wAW2/sy4
pnJ621TbFMEMbmb1zpI7Xdzt49Agj3KfBCBcOS6+mrxwOAn99Z+ZlnUffHdJ+xZqGlTMpXEeJmOk
Mlo09Ttmg2imZaVUTBanOYa9xBI1Ip0vHwxUkvULdplJUG1Goxd7dGNNiZ6xdePZ40XxVpkqiVHo
4dwowGuYfKk20lmkRQyGAbVHV2EKk7794KQ9sh4IYF5Idd/yIK193XfFnTiCbL8+7Z+nUdjRkQg7
zIt8M5ahNJuHNjYAuzu2FdP0GQEWo1wBQsDNM8wW6EylA2iYThAiR322nZqEhNrkdxaoHWKPGECV
YKlIqEdUXMQuusWvHsaoHshx9ctH0gOeEKoCsf8hDRHrJPdBZc7GJWq9GgNsfXxakdLTH2tl+nAo
TEASzGf9zZNZRtPNLWjrbJDHbza5Xut4+cC+PSP/gfraevmnllX7eM8B14hM8SqRPEWOrU4AhTJ4
txlue85NIUWava6kHR53Y++uFe+Jkf9iXG3wBeHgZITsM1ODxjf8pte9cEi6HyGML07jDMfby2iZ
at4KSwgB82ns6zPvaMiVWKFG5srsHd5bRksCqhbZ8tIwidNG3ypL1NkB7xM3xQY3gYLGthC6bXRn
Vdg1dEQEs7H+TyOGOGFlrwpE3mWnLW5YFvv024R7zw1YrwF9e7/8L+x+U0FfcIhEllQ2nxogh/tN
oOuycapUHQu3cd4UWp5MKWaKEA6w8W11eDTcWe01ObsJ+dzcfAvkgjrLSemDZChjCjOBNq/BXE8q
0Odd3zAOn3o5udvwBwPKTJ/GJbO0wJcLXbNAx/AlVkJnhR0LMWcRkU71T39I/M17U563oyErl/Tn
6aMPdqME9Y9fr5uTMEWKCDa7EDOddh9fS1Q+cvMskK4w+nMYBZfDw2Wd744JohRVQu7PA5O92r6D
Wc1UXxxj3Io034pty0psR6I1ul+9NnstWfyZSx4fWlFvsClbZWLennxM1VvsPBOEPoKL/ysy3Tf4
R+YXR4vyb+7uDiNzbh2BSEJtDI2LMsVdJOmq+0zwjQz/bxDg/1Er/MmtRhMJ2nppfBP4RWxi0JgJ
10jj2MSjjzhRmDXM4IWWMwpa87MY1C7z0Bx69QpNpX3FvFewJ2vIFCslgRnaq19GP6TYz9Sk8uNJ
gLTkS0i/3tMjcVfgCyXxEIr1Y9erUim8l7+0pG+1R+0WdVcu+M+rDezIKQcnmGaIe/3BzPXU6LpT
zjbtPPNQYvmC13SL/zH9iET8x0MMO2cAEu7F+TgY8V9YtK8OD0R3nZ2CH/Ub0z4zaWtRVjkoJT36
/2W2GE0ZhDoFutjBfK1ZMkTVPOXnCNkHxgGDwwq9lwV/RXfB0tJZNwoZqRaxgZBIteVJjNvicxT2
mAKuPte/2Pz5+1a2B0pRdRuR6EkZOPLsP0ULdHBqV6EofzLTLCO6KaOL5Kq5WCJXUXX15dhnmkOZ
p5JqVXS5dtbWjYSbpewoDdkfPynVCRKwomYsEbWe7B6MPDJST67y7cYG37Lor3x2sK2Qdu87XnPY
tSE1MFAvzHV7gAurKQHjodBiUQhce3POmJ1Ke3QhJ/ZZOMWARHJRFeYU+8qLQYGklfYQwuxzIFby
LQcl2HDb5Gc/TPVjtDPvDF62MQA1tCxFbNZOSKZUfnqi81bkw0fyXWoBS2G/vdPzqXBjrA0D64vK
oAAD4hvwZ1M3LYyUGJtkztHLkf8P9RjKqFtR3vf1Ri56TIPogl4v7o+CuWxd1Ke3eT0tXAcmduys
ULEBAcse65G3wFCM003Lt4iklo7r/BWunnsJon6RyJnFyWnb/Qk7clipgi09QmW13lSBlI6csoi2
hOp/C0lY7Viv7qAB2RGGVB6DehuERGOm9gBLDddpn2TDXwRJsonQA6AxnFQKn734nkn8S3PDNhdJ
hQxS3IbpQpxyiklxr58pLEKNVwCSzffvKZ0F6bFFy2EumtQKxPVmDuDhSfKuzFIRzEb6vuy0eCtf
/3CalgH1DV5kxcFxaRPsQFfL3AT3GjJmjfP4yHm86pPUhJHsRtxptD1fOqpld21bobKi09P4+buR
eqgbml5LXvufhV/5JWTLAm2eIjqOAnhs8P5yd3ZTOt0gbrVxXLZ+4AmzA8RJqeQsvb6JSdUdkMmG
uvSIq7fXVhSrPrs2Xf1/O5YNxEyswSCdR/g7NJJOTqlZpDqpb5abwr2X7ZWbqQaiupD6R3ub2T8X
+GsOJbAsOkodi2RqR94Q9jOEGRaq15PGl/MO0l4dEZKaR752pZl0JfVIXsbo+iLErh41ljED/15c
yaxZVgx1N8wyWDFnCxAIEis/Z0gLegzeCTx1Q+1WfUNHgWY5p2qSPQr3Hhl28IH7dklygXx+NfWH
Y4V6E/935JE76a4WmleI6bIzSeW4svyfziMR0CUkHBfmCcBXNU7eZS1XTTdAz33dNmMKPiLwEQTx
v1tU0w8R/Dr/d/iZ9sh7LYUDDOW2YcCBcDVya2aMVvzwvz4Zhq3gBwTxQl1YRzODJWexgxsaJHUh
APSbhQaYoypw7+ViiY2GGXpIo/lKwKLU9Wc3WUaS+vXaeer0Gskbdm8c22U9ec32e8sp62FDRZ6/
1UuHG+aT+rNLbSDhW6m8Btitav3G7TuM515mjisPmT8CTR4MEg1dNJRLa+BhNnI55hRRCiNbmjEs
xkiGUwkGkjW+CNxJIcuWc/mRgCEo4Zi8EbnTvPrGy/jco7uw6Au1Iudve28XbHgXFR4YPYlyV6YC
h8evDfxe3XbACJvK2OwxipYYmT0G/VSllws8fs7a7pMX9XRSROf7gTmFAMoI2pRePHuTMznt/wu+
qPMMAnsdafTiZ+6D/3Ic3T9MrkabbYmYytttn/1gcFvFhy0zjTG+c/CYTMFenjbnJaXPwWnwqAxf
LNOKx5kLKfqFBCv/d0d6ueFDIxTW0vdEjDNGJZw4xm8WXX1C8GBkg1XI6JPOAlODxzGnabjKUi96
tgbA9SOSlpBrZq601mP82zi8jk/uS90j8EETTwYRBHthQGRC+D7Tx3Iacjj4vCFI9+SVNT9KtRPS
4Pbo9g1kLV0s4AOx2bN46oooka55R6wDJFNFvtcOO2LTCnYXsrxPEnvkn+qOQW+jMrwIeShxp/ka
exDgAAaaQNr75USD2cb2gLh674A2jdONbbFtNvs+4oT7SrFj9yX1Vlf5S8keI9X6uBXNfl6BejgI
2F+wIeG8AVmtTu3vutJdQLVjJTc+eQvufiap8iaVIOZCLyHcE5SBGHIOv8Aw35Dlp5lVNT3k4k/d
jrIPs7c7kv1TMM6b3E4wvqIHxCD6fxySVKleqPZr5o4yvSFFZdkUCl+uxJgYlADZaLiuYwt3rCyl
pFCtMM76KndtuEGd1n2l38OvmQnZHNZmNdDYyjkEZ17Zo7NxWWvS1gsYZDWvIDp5K18lKQt5w2M9
ee9oLHaNovugUUO83rSPfTNfNRCA7Vw5S2UpeJC4hYYBhEXw6VhtznF9eQjMh9xUp859WqV6NfLZ
l+CxnohpNkt9qUeEMJGqWwY9NGzKPhb/5oGmT0ymkUdayBLCOCcsNU/QxfE4SL7GM7+ChIsPp/Eu
fnZgnWFj8uBBORlQmRm7hPHR/JZZlIHrmdxMRYuQU9mMZgHO/nGqCsc/KeO5MFy7YJnwhKv/M10W
89jUnP89F3gE254OIx3o+hJSnylyLZDgdK2G52iFcSeilVObfw01JyIeGKWqrt6ukQfqzk02kHRd
7OzYujMOZdo6aIxUlB/QF+K8dyYjgAUWQY8kFxkdlUyPqG2lwmjVrHA8KJsXuAhdblz/Gn5fnSkr
k9DP6VRo5iAvY/L5Rfzxf06FMgprBsITacgDVB41AmQAA8FNahLxZ2WLWJiPRyzDzN5F7dTrH//b
faoOOzm4+Zo1k3z6/oSjOG//8L6uz8zlktxRdfrv+LdotT8WbPqnp6XVbJY9rpJBRGXDvsIjOIas
hr+/RcUKiJPsM35bV4lSkkjeA8b3APO3Iv8Gm/QzX46wim9TWP1nbxqHfT4LlTvLNgthtJ5SAa9F
AKJ4gN0Er08ZSFPWk3J81T7jQoCk96nh9jnIGXHWS52paExa1ztrdg6VDLKaiF2SEpr1OpZwhNvv
APJNv4FdaPEuM2oW7hztl77IJy+lYXF0xj39KBJEQeoonKVaGW34Yc/cQ/euk9we6wV6bUJvIqt0
5qmCWN6o3/4pc/1260OHEj4fY2E4hm03Lrxjo2LG4YYos8ndszWuYYC+V24HqYfXdrnM0eT3kuZR
ZdF9bL/fUIkLFawhP3/OUVW+ZUAE8DJ6Anh6Y3aN7R2e9Q9uoi1wMHOsXBsxQRAtJMQtG+juMG4+
+Utyisj1JLFY6QLFlbjt2GmJd/VLfmPWveVTf43tv2a7EVDGKf0XqpH3PxJjrg8ifQnl/lQFwWi+
xJuS5ZJFWPKdw7qjkY/V6HnfM6/uFOV0r1GlKxDI8JbmdZwDHDc4Jk8b14iiT/FQW7T7XL7GkaYu
kaj260kU/K92uD0clnJNgdeFA5YPfP4dFdPdRV7DHYvrm083Ax9gsZvvVUirYAUjtsif1Ow2fWUX
1Ndb/CLXTXaTFpnpt3cNAOxRJt+txfHlqd8mf0kRKWXAoidoGs/Vcr8TRebB4vq1EKKjWHh7Tbyz
cF2YRBkV5GLvokO9MGmq7kcd8Wmq52oht2AShTfvkDonPIBU9pj7sH8fSn1ISqW3Pc7jkRitfkHh
nQuRMPPe6gVetDvnebW4faPTidvEE9vk1LjQeEmwSk+WB9Lm88bY84hb7xNqxVo30MtdWM/noYIH
rtJ2r79LVEHA94qfBgXBSvFznFwApd9lfVSwxxDjLqhVOimyg89eGQKLRS6VxyqYnnKPnpnRvy2D
Kk2+EkFsG5A8/SCdi0l34Tm29S+IwchXMRWxCxPsQW+cJ4KreQVi92Tr9eMMcyqIeSs0RLE/D/21
oxBv1cQnS6kVV5/OOibTEHqv9p3CdFRMNXKp1wH+pR4dnbAf2MyS6n9+grLO/u/1zxqGt2VfsPCp
p76AvnLh1fiwIxM5zYVmmgUrBlRAr32/rTfY7G5KZ4u77w6GxHHpXN65lI3Jhw0G485EYfLPzY6I
Cxe2J9BEHL6AcgbJYY2hItlTQfrYblGUvPVyg8InrI6ndEmpCJKe+yjLhypOsP1RtS/IuJZDgcRA
7d882AJj3KXKg9PO037w2IeWJluOeUTDLdz/2xYwDy1GvIEdWLzqo47KCLRnugwEDJYJctxdwxlO
oVU+4POo1dBd02unl2i1AYY4MucdQC624icO4IRmJb490dgBOJ8CDKYFBouaDmVwW8C1ZgwkLt3o
uXNBp+kOhc8/T8BTxA0syfKBZzH5DJuiM/987H3L2C2ejETWXjRwfCwjpeD/86sy6b22+FNQs+1e
xd8/F3ry0rd5awk4XMnFAgQ2U1RIDKLS8O14EGaAbKvenLK3CrTLh1r8+l7xkotzLv6JQn4lTFU0
DcL2zN/yG4bUP4x9jMqgLRxM7r9oJdxiMI3j3EbnFHm3/sM/vsQ0lyRIhHSBzdVyJ928JJA07DLq
kFzElO2zlF22aTdk9D+IYVHkFW1hqAXzt5rGKkZtJbtrshXqP2nAOtm7++3bMHc70yDoFuCZTwyl
ORm2W/tEurnGgMxIfZghimogET4g/q9bALta0rMzZyhyPE/ADTFKUlcwPRYHLvAFEwmFe5ogQ9B8
cyxoctOY71PkTHTrnXXOueQpu2+7Q8yNYnPqLlZ8lOlR1xfMvQp+UNn3pCjp52sohv9+YZiKTF/X
n+4xOnmQd7D6vkh9FlAIv6uYXbOmUrHJZOlMW6L0DikO0G0llWlq8mojlDstqyPKez6SZAu0jD7Q
TmQLGuTdBlBVgAAhuYcKwlP05u1lTuTwsM41q/YptTjo4dqC6eYBUHQIWdEiAlkDZk6s1ehJISxm
v/qiDX5Ovs1f68eZj1b2tKkKzsZhsmM5Gs/xhgval2CYGLUUqc+y27CyOBpJuY3kD+JIc0SbRg+l
7Ce9EbO546HBRiyQ/rxjX2vv49vY4ZUXOEq2ZsWDYy6ZrEyNfp7xWX52sR06rUT5MAxlebwSsdos
0rUgRF7EZ45NInB4/JZGbAyysA1s74Ymq2/s8l9u2aDyiy4f8yiCe0/P0PRmA/B2qcP34mX/80ZD
yLpu6wTt2xqRgYxO2MUiSyqgHqLl/Bv4fCHbYqiANTsUFGo5ZRzL3ygkHaHSiSgANUZCHp1Dg2ZN
fOtxDWks/TECyAlujOFaMFH/RfhslVzA7m/611+zTtDoxdcY3ZXCy6WJIkZyNh0b5Qe2Hznqbks9
3ox5tJj3db/Ws0uYZ3iDie0oam0IfV3TE9Q9irtLXP0utOcUzJDMBQw3tpt1nwl1ua875o1BKq7f
c0IjMB7cQHvAt9UB9vHjsO8w39IADDARh6TXkbvJloD4VwRk3AB2UsVslcvoZ31R4W7qTwc1vqp6
2QIHzxOPog5ULuRv0R800DfKxX3JE5KPEuAXdKE8MYL5EbUmIu+J+LuzKwJCILTvYWXwARi/53l5
pUjdzkI5ZzzqeF3fZyksFSdACYR8arEEyIbwdzoZe2fp2G//LmubkllK43q0YZhjklT0i1M8d8zD
nPLE7QrTEGZ7LKhU60OV5P8fuNCbkL6m/awLfJyaiNvrLvMf4j8ivo2BNPZnvSDuuGDS1K7PEHt0
o0wO5zPoYZFeT/g8/ingKk1goYbHt2sCTwQTF6pVZKvetQCUXKkR369A/4u2ek9cnLHdyS16Up5Z
zFLCzn8Ke0M1fhdOg/GXc1nmOv6BfEXmlAeF4Nl9rdhFg5zlBvJ3fmpZ/bVKUPv3Wl4MM/jOgAN4
QgJQDNADcdxWH/+2BKkYI9xAmsOaicHUyrz/d0vMRbSroiWo0kqIv8zwY6n4N1KPgPer0lf6hVEy
40KUZvByy+U99uG4iEdmVLXeiOPCv2OUJvrgT7WpA2FhVywvWrU+CWFYCaxsJVQ8EoVfOgxJ06XG
ZjMmLAR575P+Ec5Q0Exx/FGeV/f9UrEpaycrxXWEolGyRmL94ZH+n0P3VG7oVmhSXvlfcGw/tJ53
3kdueha2d1tPu8n+s+dsItQSlDstlTBo7s7kkAOjMT+LieENM+Fo+eqTKJ4VK20jqIRFn6MQb/cT
hmh+y+DPYyZATNguPsWKIe9bjsCiu727/LeG0hC3sm3d1BsFUX4s7kiTKtqyOSMfeXvQZOcXF/X/
H20VmQX04EbPAFsbr9fA2Yzb7RXPEvnJXNhGULAMVlEMKEwCTRArDpyWcTUQCTJnUZTH2RbxMbq0
/BqSmjTWq23lJgpzce9rYDXW1kyzygyicRWaO9Ag/EKN7y7uznZ4dDfXOjAPb/1rEMbvNuyDlxhF
KkDBSBROQBewbDixuZWHK/PQ/aRjXc1+KBjUUZWR/CTvRlIeu1syi5S7l+bIBlRchyUE9a6+5Xfm
8msLrUbgefbVZA+EK0a7l4zv1k/FdE2U/I28L6aftib5nJ67/SJLmJ7grB2BnpnMpOdMGEmmgdoJ
YfzJiTAuIv010bHlw20rbkjI0FF3QYDOsPsd3sobCseTSzg7duBW4fiTu01pqNT9jz5XlBqQ9ZkK
Y7Q+iCC/0NVX6yVlrxn4U9NT18F8TDExdtk/NdA+km0FZBOB4RjfkvHo/GaWVISJQG5nQKAWenhJ
XksC/+QnQokffWdfH/88SEP6hNwimwM9tA38HVqixAru2z3OBKHph314j85AoI9IIFeTHk+s//1s
Y1xocnECHuGl2s4/h88IQrrjspFn/vpDs/AmCvZcuuvnppbF6E+UA0P47sUpUIq/pOGyJxXI7SGt
wzZiHVxIgTlsbg3b+FIumrqPs6m4FfY9KYpgcvciHi4N3KFTQa4/TL70/S3fLpqbAhfKgK0ZldYQ
MOzJ/syMzMYQb/kCXZ5OdqzlulkS/ZGu5ldEzND+kv7sZlMyR8oqXvcKBaOytkNuHmbc/aZe5r3+
5fLrZVQb1CwDXUitbNYC8xpUgMe3anHvGYAHBUQTJFiuVhePl8HwVaggeAv3X1CaSSBGdIjpGz+/
zGiwDClFB5AKaoreKz13iqa6LTbxrRifPw/+Rlm+F/eP4i8ft+4S7txR0rRYQI9QhlW/donI8Kjr
WXln8TQDxQV1yBojeDKBjFZvidWfZkeoSwqFpk1xvg09/cDc2DJjYOXg8QB9wB8UKngu0DV4/vGR
AHccC3nBrbps26ybIYOk780Srm4kiBr4E8wFPz/1dVJpZWZTKrjmeKfMsQoigilZnZ6tvJuiTblU
SXpsKS5+sILKYcisKAJORdDxKZgGYaBvtBy8I2ryxi8CLofF/BVIlsM4qe72rqReChN5VyN9gOLz
dj4GZObuBbMaA1Qc5Z6j32ZU4hJn29jsZl0Pn09Jq3rf8Vhe8rCQyqrvml4OMZxc+eHBCtXRNuI8
ndnNSZes394xgbAktE3hkMxo/iGCbtfq0arsAq1HSTN+9L0WQmVIVkQFPL2HbntFpWj6vdf56qFB
RYBl4NN/9YfPBu2EgZu42QteRX2I3l3XTqXr+pEj+CKTfdLCHt6ZCt8cLkot/255472jZViqx7qr
NwElWhz26qhbpSYZjRec0Tm0fRmG4aMqGQdVMRb3UQZ+ZSdwzQlnFVvZ5FitYP6x9LV8BbTFvLoS
lqgZaZMy13zo1MJiYuLj3UaHwaPCen/LvduKIVLLrPno+WRjyDJWH2tgah63bIiZnaw+V34vZd/T
yPVniRZNLkn5f+gPpHD9lIVQdFPhqHZT/d+VD/+Oc2lPZ/Sss5zsG8hQdOWEvVsJAFGVXJrAkyPv
88kRCmTyOuufbwE8TiYN8TGRVf3vSm5mMVo+HsuV0Q918ZJGpKvsrWMtTRNQydWHlyZrVN0fF7CD
urYFPZh+XbELXLji7J3NF8ChD6V5p0ZtuLzfIzo+dYOxbmmHW36FmSmLo4dA7eYurcSD04EdLydh
+2he6zeYNZGXhoS5Wo4ktpnzjfkOwG4Z+YoRo3JiNd90lMTglGHi1lPL513LXzp2lXloc75egf3P
CyZFnZPLm6b4gp2+q++xAX5MHgjUD68h0Eo/ljp2YbsxSSXUJTZy8RgI8gmn/odH7NiQQ5m3e/W7
acX0oL3tJIn+0JMzny6fC6phbnVSMuQ03No4VvXtuvAL45DpNkR1iu/Bon5AkyzBcTndZsRBUa2B
C9GRjHly996AjH5cjPQKYpDU5c9EcWUmEhXUJ1sV+Pizj/AwYsVpjs9+Ph9wDwD0+QEuFjB5RFX9
EbZ4vaWQgcWUOPyRG9UggdQRocJXAMB4kSYTZMFFG/ynkUNihXNT1Ds6//PocU9IrNCz7GS5SYnx
zCHxE61MEW/ck9PjgYdlqPvPhjJ2UUCtm2MccIZOYBBEz9kqDtak9RarEjJWVRs/eaN9vjSHINvj
0filYaIhYy1VE5AYcUJ7WDJGEcX2Qru6upetO31baZvy9q8VI31uOfWhmyEgKnZ3tYO2kCY0wKb5
pik3L8q26QjWw4ONvkaXPUYPJxVSl0YHAXB5HZIliMU6ny4gD3CNAu9k/VdiYdPzOHdNA6TZ3m38
IevxcOyndDzPHlh9Kt8oWcXhDn0VoL1y4wuMuYQmpugsYuR/qbT5TwVkXYCqE+ZF0uHi6kEtopmb
sbCGb6PSjeaoyU7crvGj55R+mQdjBELYaqi31yRaRY9+z22cNZlQqa/SfRBbpOsUK7KgQQWIX88a
9F9sVpDWtgRVSnCIb0qPeJLNeG/ttHcuCQkZcJapsm1GekA+9TnLb+8fAzMuAyJ1+91j6OV61CLk
PHbNy/tvy9ZSh3mlrAcYjqmOpuIZhkaeQ+D/AHZWoVqwTg5zq3tJ7QIhDNDmfDldlyr+J10lOBWC
RpHoHEXaxsvM9LFMzVJMFLbiF7MhNzsG4LLKSdRg2kyxib2US8KHtSZjtOnc8K/ILVuQKE+/60W4
pdC8fZPL2a2SJ0u6+RAmEmbFQ3yBGPh9i8XRJOJcdJGHr6zWuZ0p3eqO4J2Iw+XskajHSNQiEI5c
v5JvHINxhRVB5c2CKC4deQp8km+Z7LqPvokXQZ2/hu5SvB2wU9IE23MDpkhHWVfZdM4otmD33MEo
oz2ES1LLYdIPXAlTTXq2PhLdV1D9P1PCuhO9KeX/t4z0Su0DV4bEFj0tM/WemBZS85/A1Q4heygr
VwvLgUQ0GCFBju38gKKv9CC/Qzgo5TP5geTNPmoD0BF1f28JEVTSTcNpNxr5omLowRldTiXGGDYp
pwY9iiOnae5h/Mc1z+dGZMaPDBuTgD3/ShQs+XS5MidbytS1HttIXAzmGlF8L5+ve3Nsl0G72PG8
5pblW9bl7/TWLNBAC+rFCOwB5iLxlCMC7XZIFngtcDA4IFN7WimTVbifmEiARsBVNXJj90tkPC+A
G0uqtcdSUSwIF36BrZZIO93XGexJOwygULLldnMZuOomLbS2KYOVnFgZ0NvAoix38dxOKGIY7GKE
zt9TBZOyYOB66GN8ux9fnvv5kncVS2+ODGuoKMwBU60SUiwX/qD2NDbb+utMVjqBwBx93fGd4NMl
QITm3P54H1uS+KoJkhvr5gMq2YkdXKeoif3jZT6S/z4a5jAo/t95JtlmCm0ar9wSCii89jnBQ1+e
IAzpzY1vXqPjG4JAiTw25vjXOtSa4SXr/x9jExsc/9JxLULmqwC7NIPGxdicfmWKJorWhqZnImwp
4cHm6uzxFCoHjDpsRRaV42+THKoFXhrVQHfp9nThh+eEcSnjal9v+A+6cNqtGTDqaAMMpQPPAm+H
f3xPRKm0jCUAmQLHilUnw6rCVFiqgdqkMvaoM4MVMDTdYTEMpS22NPRPVnQD8cHo6SyZTh/O+xYw
y1oG08daBCi9XPf6AUslbMicyfuIxrh7l+EsE4F9zNa0IEMZlU817v2VkEHEl1C9UNJLhTBaOOjK
Y2179YTL/ciQqQPFCtEU8GmJnNgMR8ROZqVfn2tzuv3CWe9Zddtdq2Wta1HsetLK5pyxe1eac0gW
2pOTg636B7SJIuVIvTQiTXlZaUiST+eq0QcxO8LVue96vKgs5TJBo9enVsBqr1t7gSgKJnRLF+pP
CYRPyImBUR3PQmZYeancZ5n+az1iTrep2UrBnNnddTwLhrhdssBaESijznyOxpIZwATNjhJxKhWr
y266rlTZOesxER5/VCJcAKjcWqZDigDSK00UNNhN4wkOw6Qbu0w1ZB/8FAzgjPbrP0CT9j6/DE1g
UH1MS7/jJSViRQqLnawcnrU+0zCVlEH9bw6mxdGL/czrOQA4HcaiR9AcIk8lmEraCz5aBAmlTPiO
Jt8P8crjvv8VOCekXphU/NJa8C9oMGlzCxvzIJRPPUMern8OmGCR7n5xzFOhMIdNGlh09NtF3/8E
hsdTtUS1iYOHdAbvDMduH2dpxtNA9h81qXypFlwD4uGyGizTYIt8F+KwjhZDf+47GvRAasD2vTcP
JJbl9JWl0SJzRM148vSNbw6a7cqAVMCcibOEcObb2T7HBRzbYCVYsBPzBFwURGRXDtGJT5asl8ro
phBhsbL8ROmApyLR0pj1mtznvSWs1XwCMTUh+SsCIaOXW6oqdDJKTZUMigpBRFYhaJ0ZYlemEkz6
v9scSWImXkOeBu359C4+PfJwAXd9yjnW+RNTNKCCmI/3/5DWn77/Qbcw3v17hKJrh20FlwCqTKwU
Mu3kOpodrgd4NSj8Jgw822KH5YQmWVy3cNVuwKzMMD3vDXy3ys+RVEVZdm1aTrcicKrrv45XfDsh
cVh+U8aQOLw53Eul4b1+gYeWlRrpEsCzr/XdJNkKmMNZLUICY0MM01zEr9E7pPnOuc2BDhVrc08E
eMtZG3t44GongIAhj9WS0tF3k2T+nr3ATvaw2kF9Usdwi1tH7AHPmX1gKaGTc/6jUOGTPTOyEc7X
xN+doVlUv+9rrXrLb7NTWdtsIXAhXr3PR2b+2zZIlKNMQPxup5pC5xpCZpFMMae+D8szkbzaycVf
1enqKw2p6bqTN/20Vwm5xKZaecFxoKjnHMxRYpdnSN2T9iLaEeQX4yqqzGrVzXEka3cLCBhVvnob
pUjzxVgSzruhsLypAW9UbVBiGyj6MHPv9TBe3j+FcLxUYBYHC048wg51gx6hRu4Qwef3rDg9uQHD
BwnrGLR6pxxcoj0LI7ZCGWY/OwNEHD/SbW2cbdEwMxSSul5uWrTddVZq03fzS1x7eTE0Zm5PBkvS
N/1TrsLIEm2RX3GlY9SdCwAvQz8BRGHpwcMoZgoC1S5Rs6U+79A//ceCa9CrMHVRYcS75BMi11Ze
zWGTY/l7Dj22loyihPdEyuk/VUhuZ8MYmwj6IW0TE1ygYNaOguDFtf651W/B7TVN1RGHQh2ySKrq
QEhzbpo7AM9ZJzrYaJRkpyFla/LvDDYqIO6VV6rY2904Szl44KayNhidJ+hXLWpRX0Q7eFOJeSPF
Mpe9HVTi9zLDLSjSVjuGUusi76s5KzDJD4iIt1PstW2cwX29PsGA5rmYQ4pJ6UQ9km9hF6MVFDt3
vDpe/qqWFURIAP9GTnUND3bFchwKGS5+uZzq2iUVPwrhQMlrFZPQJuOneRmr6AjO0qIys8LvMGqJ
YR06Cr4LU+EuJqz0gJ6vnsL8Rmp2mjiE2K7aPH6ivm+gECUWOD0DcK64DS/vVkk/3L5l3Mjm/TjY
q1Il9+MIrcGel+1YXMrhWyIPHs7VKzdqFJ4+vCA81XpS7XTQ9eueVDG7rAKBw6/wB8vLYFGuExAI
t+TwD36p3O5B0rfKhMS8GKRYydYYGmcCMF0ZgHXdwz7+f1DWpreYMzyMLzIgLDgzDeAqjJvqR8gB
JeiP/syaqvVjW4DXD1QVy73HinWc8OVmu/f7TOrnBlxjr8OuNbaUr+RtRk8tbCoh5lOHF1z0P4i/
gEG/G0fVIPZuZvNRby1FHg3t3sUiy8KVdTby699C2XcC7LbJkvr36TDIMs29BBeH6AR3EZH4cBCu
+IWeuj9BYr1Ae0EIuqED0bsllejGB/xCtDxn83tqSJEdQ6mLQzuoZhHIs5MLPsPt9Kks8y6uy4LX
rR3G5WRvr6TQcfOyRSfpJ8W/LjLFLZVHSd6bmFzDOqS43VT0LVO6t4xhOJUaIva//K7K4dijWZNF
W/x3Kp12ZIK3a6D5GmZU1C/iPx4V/wyGma/1dettqrjLZkBewKUYVIJOcA3LfOEoCeb6qrAYY6M/
EoUehiDKJQCZ9T4eD3a7l08smUvBLoN30PN7J8Hi5iAorddCwmfY/Vb8NhwXMgmwWWXjVRbtB/TG
H6fNTp2aTezhSmZDFQf7KEPTTz+da/1OJB8fbeMgwQolVvjRatQ6y/jfMl/9RxbYrGi6ClqWLoFm
Jhhoydibhct0TWhpyc+bnRn4V0un6mzdBNPbtF612o+bnIgLOf2RGPgPbyCvOvugyolQwa8B6eIU
qPD9Xyh9CBXx4sXUyaFmevDXEKL6xrrk0ZUUg/OSWo/zf3MNLetTkLg41Z8jPgpnCrBda7au83GO
UIOJcdhca3o+2X28rhqvqPQuWPFRjUkBKWD5oB1aS4Gykss2n4hpSpaZOQBRmKQ4KB7PVOjO0wZW
pt8xMt88tcj8w7VdtLJMtHfXG87S/B1ZgPmvX6ZMySlwT76Rz+OyLfddx19viHeXOY3emM1rYFjW
pxUfV20mgs7OpZbd1D7hzTK6Kv9zKxg8eOQ+/biNG4bvy9gYUSzhnUnS/4Pgb6/HMEzlE59far8L
hwuGi3NeQGlrRi1CM84lnm1pD77M6pJXSqCka9DwZK8yH/kE9+5tJDhExKRDKCa6X9QbeJ9IUbTa
DBNBErO1tNWhYmZnpqExioan54OPyGrANGqsEwRv72zyjvY9v2LVoGHg8m2eb3EtWoyFMYXjHRE/
nShxG0uYvwhNHffap9GDZc+FWc1+SNRgjJbLgpSR4BQRjtBhWtUL0g1bejFjzVxai3qdPmsgT1A5
aMLwooLbOL9n7ex7HFQY7W0muRxkaQef7PvVpMZYG8mk2m6TcxaOrT8ON/5lxShL3HH9qL5Sn3aL
qzQnZ8u7Hw3AomMh6naPSGglsIYvgEwR1l/p0ZZ1lgVdeoLzmkdmDXBjDxeqojUBSxCjO+OmJjO4
tL+X5dJBYi7A3HQFDUrXFWgTUPjMdTFpG+bHtxdH+Lt/AX6rsgsRI0D+BRSfmNpKVLIU8k1v8qLh
GY4b1uDREUIq6um5Xf0OTTHnMRXYsuEBasAcmn/1h8vVpO2SLAphmYzo5+/k4SinVt1PZgUtpWvP
bdENrFWMnlIgTOShWrgbsnDuFszEat123YD+FULJRfhYE8lvhm7kHCC5BKY1Eeg1Dey4m7xaFvj0
L09I/qdGIbfWPOyUJChpGD+EoD+r2blOl4SZgkrz8oqTnAVOvXwtFtTO2igs4cv5J6HOr9CXhqoE
K2OPa+sBGlE3a2TtV0ATR7cnYcxOqIQB/L7iKCERAQg7AVrJW1kLf8d7U48MibiARQ04u+QHzpMB
aMc9ES8PPAMjlgQuhk98ulcxvLqz9zLoT/fYUOVAeXILSv5fTf/qe+AiAfOfD/w8s2MyHpsiBzCh
0xGgHHUMpWdDnBJtCwks/R1ylIlIdCqoOexz1X09Azw2lpf0gv55CcKwcYyyeBnxUUPht0tV0t5T
TN7Xt3tBN8FVoJ7nHrsdP9kJ3n6Jb2cmlyxiBgGPZxq0Hu34Kx3sJf5eZXDf+mjpN/6xB4JurFWC
rdtxW/2UUkG9GqZg3fugZJqGEuJBufM/DJ+Arjse729dKv/Afqi3Y9CKP76jWdnzJD/DuOLgL0P9
sxKmSKQxRYXSUVcATvEN6BgNCmwUlAFqNAtx8p3i2j1on81Nxbj2nm+a3/DGq3Y3gHanjFcNlKqJ
M0BVQsvkFMObqmQDczKZBvIRyDHPqDSyL/OoBAi33plXwW24bkTI7AJROlONPnOIYL8P4vPC0rks
z7ZOJMQloybS2aVIUmwFMv04TLRRSshtdmi4xxVZLsjgSDMX39IeCuCy7Ig1LtRYcnzyXpt5Nrkz
XsOKdtNlyc7oAs0QA5EAG3EKpfZN+L2H7RTeAfuAHxa0lReQgAr4W4jQXpDZOS78LIYmI1x9jgJJ
L2QBPWi4bcDsRlivAvfPqAfiHdfDlS2ilmmpIeuupyvezU/4t8mt0dDPpfX7vtzeGQkGBms4v/21
A0Zr75qq3hNad250ufaa3y0mUgKlvuI3gbqMKsYVcrIba8u4Zo0DqU+qSUsL0Wkjn1gyUvWB4cla
t2FzpE5E4Kq1Mbx9l66NHkBv3vNYnUAinZDOIgkD1diFdWaO7KK+9tEvjc2wIe+J4jWjQKPx0vlC
Gi1HgFULhfr3ocw50XLjHZ7cF0Vl5mwZx5ggpKr2MGsHetsKNMX9yGKQLYaWGyvji6DzRFMoHLIz
PcMijX07f+VxtTH5vu3HQ/QS5rM/rWuIGem5hzV+NaQnSxxY8RxRH7+FI4NP/sYTKpWXc8GcvDUO
5NL5gt4KIrW1lXKvg1ZToNQTNH2faOAK/62Zu0h2PS01v7LzEJzUAGJTdOgcpVSgANiHsk5wW0CL
k6v0eWB4KkROFldkm7fri4HznDn/kG4OdyCsQOp8Ma2E8morAfHIyJOHb10rTaUcCirjv2QeesPQ
erYLnkbILx6ioumq5ThnmU8kBt0RhDWR+xHh2bMFjNAycDPPXKcgyfIngWE2Ec1MR7j+1nfvw+qD
Dpb58ppxVir5jGg11yNxPeD+tozqsDuqoOPD0Ns8FJR5nLWqu1fL8qctdbkD37h3FfZvPzmsPpXu
+vQgaBwkh+6BgZDWN6wQ8S/DGoGHpeSrVcmexYVg3OLNZTlLjWQl3BXaLBhY96HK/J8VTk0txSXJ
U2/uR/l8xRf0UUXOWwuqHE7AUiDd7elXvTMWsfKmbOabqRAhVHbgswfLu84cXF5Z054Mekix8qhL
XxsAPwe7Cifj5tiV4mzYaACtSjjBgg4VkaulVVSAXkDo0TnZ8go27OEhxDK+ElVnAbj1OBaYHFnn
fBnnZxxJGWKLEdnFr+amPLqN1N/c26E6cymDmTU2VNIyFHyEg8oSy3Wf2fgFXRyWCshLiJwkqqUB
YoFNTCZrU7uD9xzrOPawA1kgd2N0G5LFniNlupgpuRuIArnlqvb0NJRlF1ldJf+RtpPqTUm4Fgy4
bvuj59kFEHCm5y3pUeKzR5U020zVer0uMorZaVgi/j18mrCOwlAHQc21T7yhiXSr3/L8JtrL9BlT
1B6dJqEbl4nBkFHbL2Bw82WKCNJm2jwdqaU3ONvy1Y8HHfJOrG72JvcsUKmvzhIJOdkCqEPv8bzE
nCHWEUECWcaIjzcChfX0TRKfrz3qxsGlVbZfRdHJxIf2D4seAkFih1ptXqNSsR/cHYIbUoVxvsBN
QgI6r8/j2t0XNYsgx4ZfEnLilzMOdQRfmRXnm2Rc4mxFebL6DJeINsc45qEtst+WxRtDG4Q1py59
jkvU3F6EeE5XpwwX40DTpAvxP+w9eZch7N3fCshttys4KOWYRzBJRldY4m68ux5W7V1B9rlwixPo
PKSdRJI9qJh5idlC7zMyYS2j9gdUHBGbWtwNpW0HpOFtY9DIRg+wCZFmPKEDFZDJ/g+j3VhNbSjY
umdYRw/WOKk4oSfN1BVJ54DPV5oGf4cF6OgXA7TS84YzJ5impLgpMDnbTZyoRf7wAJafZUpSnyco
3WJXpGIN+luo3FJLX2wXsz9ytTqfOI+aHQIgGG7AZiAd8X098NR8cdP8xsUbPPo4HwpXSWl4+epl
zOEA31cJ6JY4eQJJ2THFpkbMOKc0rHD+WJnyY4sNGrxLSZS3YMhpc75y07wbPQhJjUoYgBsdy026
SyDTVYasLzp6TC6NsWnl/7eQFJElaUJE64ZW1XO8uFdWjLeBhA/Dy0Q5XYNRZsTQ76O/iBZl4LAG
4gSimCTBQ00dMVFFzmcvt9e3C+rGD1zbTW5XEQfFWS05j9QYoY0pyeRnKo+BKAOyFZE/1+1wRobz
jQZdGcbdAmtZlK6Kc2vBrglOy+jTQ4nm3FN08Fuwxr4IpqqvGOzgJ0+V7H8/G5yt8M/+H60Me5/g
ZPaYecSvcCgW866A1M/5IVSwezeONwuKRoEFI8hfzVJhxEErHQ1d9brVYkGKX90ka0z3WRU0WkzU
S/Y181n4WHQ5IFT/S3Rzk4PDaguzQ7gruW2GovLgelMH+5QfWPzbaLirYPMD0MUYOxPFkEHAZhll
cOkP9iC2zqXP8H98ol5eJGy4PC8NY9+WuRR0eoQG0a2qbYpi5pEHB/EwfAauM4iDv+GK5nxGwbKn
TQ+R+O6UJDnmvjWzSW+Dr2qZeW8taG4towI79bt7MMn0g4lITQAolSGWPfPm2VrrFjXAeexSVWta
0f7JmvevoWogoaijajdtR7kXSfgZMv01Vfmc4NoJCW/6QiZSH4if3A/C+DMoNd/oBbeZYkqRPKiu
GrgeDyTfOVLg0CoBq+f/hPsv3Kii//RD9GpUZbuoeGk0z4QEZx9CuuyTbo9okzc0RTfDe752UBoF
FnNpINZZCIC8azaLxyJLuY7VeSgqjQ/U9QP0uqWMDNQjJ/JUq8FFb2KtBxAUbNnXbJOn0d0E+RxB
+Aaca48sUK4Ce7jta8ff8TxHV+6/SkYlKmOUfaciX9SqG1mzhiiMzx4rVP8B4LM2BkdTYfXx4jgS
2ONMj6hOuuwVCRpE8m+oPtA5W9NOKpiRgKZZQMuHQFn47V3L3ExOv/Zd0rkoM0DVCd4D/w+mJq82
5mCLBXQCK2OFo6djmAST9n2x4QI/qiZeFF838cGK4pkB82XxKOy+ZWDnhh2Ar61gqUn4MlI7bA68
bmxhs3cJeALsZYCJm8l4PbL06x48lR8MP06rJbmQHRmijgeNmzi4/p/aIJu1iRJRKIH2HqnSjZ7z
C0rLUk3yIPlqhEAy3gggBtH2Xhx0MbYj1k65rsuPgFxCqezxy/7sTKTp2gNsHo1rsMfXPZadyHxW
izqQgyD4pv2REiwYZHIwTaoLiiYTa7BuIZcK2alYTJrQNV2L8+ckuCFLnyqitZiI/j4hLSHj27y7
96KkjpnHdaV7jdqA+A+rCPufMS9SVcYAqsG8buALogApKkrHFe3fPCLTDmIw/Bpa4Hwk3sRYGlp+
8lzssuzLO/j5BLji5g788+vnVSrzOidxxp1Tf4Qc4M+M/DTH0RuB2SVdyb0sdarhez13PATiNZXc
S0cfL5h4hB+Z95I8sdJ42CHmiCiQnHy3TAEToRS2NUwHeJNxl9PLTXiCu1svabnl0oyLclq8djA4
qUOElL1qvqysZKjPGsXs6Y9n5fLcWSyuWk/iQ2SkY0YZk8Cm0PkiAQ/ToyIkV1yOOdgBUUFEI2Nk
eUTtrrfubigGTkQbbCOFW4oAqvE8bw3dyi3+Xti0X3aCXIKJ4oupFBN+JPkIjofPCDSw6kp1EJ3w
zI+qH+PdKhpI37Z4iJ+aXvbhbAPthtJVGPikZh4jZ/oGNWS4GS1iEdKYOBX8FIoCtPVehn/DOn/3
oc4+dRXj9Oo+ccOWDKPoJ4rrpZWfZ/QwSAPFChtkdUpS5PJAePReix6AinCb0jmH5dMoDDCgxW5q
83JaZfQf3K9Ro0S91hiZ14Ey84icHcy60/vZW+j0LDkfwAaiN2nhjU8e6CjxPH1QmOh0BAFvdK4z
R12ojveayjEOoKsN6xcrcFvpG6Il1JRS+Y2CHdeyPP1yp1XAxEQ9BSa9+pXEIbKTdxjgg4B65haB
6oOtr0wbn290TnrRMmB0GfaEGY+4YLfPJF3EvrNlIgNQa7g0LccWCS4u+fyosSIAZkO/WLkGRYcn
Iv7Z6Js0kmGSlX0OyizOWaCxIOKDwyLafYAfiFHZSHQMj3L/P3CsGV/iNHaCvlOWnZQFbm9UhSw/
d7roJkp+g8incn4e08vyGt9ZE4OQA5XWNHGVWT7cS9oKPrp9CI2w0jOAot2b2T6iZUOWPiOeW27W
otZWAYHZsnDtMVWzBLYLtPsuMJUt1hye1oKi+7ASczXc6l4BD1FFQ8JM0cABpCeITrQhA4mBUj7h
coI+ouRgov31JDkr1sTB5ssIDwruc64AfagVMet/ZgoIY+r01JRtuBa3d7TuwzTjNlO7HDZB8Cjh
YP6hai0X/52Sc6zdRgMxy2TR8Wx+ESIboI5deuYAoqpJgbH4hk2ZkEeAOJ9UwouvYrb14nV2h4/6
frxaT9SX5+OFZCLEUrgY83vrrbXL3UsffyEKLmFOobgpdWofPSj6WmSO8fjLT1JFKXkgVkB1WPY/
mS5QkcLX9rEboOfkmpKvcdksT7hL3VAURrIF+v4k7WlxhDRWp0yUxIh/otv9Xy1u/8Hucs8jd7nI
IePUftZ4IeUQQiHgfm22B+LOtMvbCwPaPjJ/VLmQOSBdOuj0kwe6VvOuK0YlX7PL3n2jdl5H4E9L
Qq/g4HPyOl0NMV1QAfYZaRy67zXa70Mh9b2o6yg9/aZBYEb2fbNP3weqNnc3H/2c5OQs7DN2x578
lhojbKsIuyqloDqqyT5hDfUCHduDsYA4oJ0uBRKjnP9mTwRk/gjxJ3JaKac3wY5zFLfL6Jj5vAVN
3cIxCKbs32M7l+kPwhnLRT4Clq+9jynz1uM+1lAJMNcKWVGBVs+AYGW2QUZbx++cSVLlLrP19Gkj
D4Adz/LyyWW9ZKY1aGojMi9lTOjOyL/JZbhpPS8xRCCM6dNS9HQq3ptXkBXh72htJI2y/QuPxbIG
VtqmGHpIPt413JPf0u6aw9aQmK+qqUAqDrvO5kFAqRJ78a7f3N/nbGyEH3AHonlbB00CGnw8vUmK
3V21RwLpv9QToTE3nr741CxJwWg9BbIMIKAcQ74mFrJ8JVq5OzqhECVqW9DcRgWIWu5KbOcAZ7Wz
ZxkNMPBHAOjyEadOLfgn3ImzfA1a6Nlhy4AiIZ2OtjhpsqtlmZ4EM9kWVkOXlCMTDzdwPrbkjbDF
xO69xpzzLiNAj8YmCEFVEps/MmjUCzVKbkqGPaBkUk+eA/ufBkREsikCzoO4b1RBsX9OdWaeC8vd
nZ1HzpXeh7IDZxMb5SKX0aUvH5iNG16ss7Gp114H22kO631J4QFqC3k16qTlwQgWgnYrOhc0Fo9f
v4tpwNnzoTD+RhYeA2bVd5sXDZ5AmQKn+mwjuzYYeb9y37/WGjLp3UzymySML2MOlogNhuC71Ip6
urcsnuwUUFwHvIe9LDDkfJGRy0qUiMQ4KbCn/re1xswpQBAj1CHccLs5fWbSyzrNde+06GoDIba6
KOlGwHi088PewtGaPAmQFybXXVliVO/GLJR3q8f5etoTor7dRCe/W7YL1kzxEhp7/CNCrLIqj7Cl
c6zIbykxJBg5TtbrrsDJ4OY43IjaHXGRQz0UK+9JkjpoD+fkfb+o2mm6FiCaeCrxXv0b6GAlwE6H
OHY4q46LXgSsyp9cgOkB7uRRpRy/4jgftEch3GWQuI1xHl4/QTuFMue/P7KBi6L58VqysUlbOlpx
q39JDcJD0oIYYRM3mLCqAPsYYabG32QFxITmuAUlLn0W7BMagoYXiytLebd2Vdxh+Qtldlodpp2U
pXvSy3vDs0QQ4q/UnZKl4x+NnUxGNdaWqsDcxtuV763pWktiZi/gLnUmEXzmsg/VTTU3eNryEo8p
wLYWgCiYjC0wdKQw7seuVnZ9ysJKcjQw2gnRoGcQxhTa4P8jjagpWV3M6Qn2/Oj+U3byBlYN1KSS
UGH3UFW88ogICX4s+zHxjzQbWcxG5QTKeJi0gXl5XwCv8ygI/MOtaOundfQvptENBWGq2rkLSEiO
Wp3UJ6LZnOtkE/Tv1rNsO8KuO73BPG04Jjm7SCPiJldDC2s6Fh68G9g4aKah0lqcTeDF+rLC1g8q
zKQt0PNXRVTMrQfMg5k+dxDTwAhkPNbrD1XUREbCnPHMXIJU6YzeaXruze2DAPMf/g4QfK4xi8t3
W9M/aSJjhQtuIBLomw2BXfkUlcGAzsSPrkyXdRCPQ8utjlEgoCS9UodYVKZYTqBEvsKW6iZfBpjR
/8SCS2ZK7DKHxpxZKDFZK9gb8HBhpxEnp+VyhHzJ9cYA+lzpOtx5PdM4p9m/vIXdpY2qtxelchzj
4/qncuNTMVIrg9MLfZJ4fCAta2wgwjF/egfJfZ63YL6/v14lAiQzdRvpmQ9KKlZ+A8wcRBwqBpBl
/33aRb0ara5H99iRFRBC/zUhukT1KsOFmWIMiKhWBJKE3U1ieg9tPe0ma/+BQIGwwqxeQu4Xynno
PxAm6EL8iXXVHsIP7HDrPmP8wlCmkToLyiewT/IOEYXzj7SqjMQ3vnIlkcYNcRYAQXh1odaJksxK
yd7yZ9xiTS8jQ6kAWRAgWuUzbLGmXCUOrdVNUwBSIzfkERXglzckrkLUm4jeq4QdcdrNJTANjXlP
OqgzD1QZQlYZvtgvxZPT7GrJrOrLIHlN9hS/kpVoEP05OC4a/5IbGtNe0uQNZ//Tao4cn+b8dlha
erz++/cvrNHpPU6/wMdNdyedZ+yWMPA1BuQJfLGFhkAjUeXiD/H7Uf6zFGceouhryjSuNw50xxVM
xPXQ3je8lRgopNpQjyws2/AgemzC++BwZKLiVNT4r1ejeFAeCOY8t+k1krapjd88x7lEKBQWEm2E
KYO6pyArN31MbZI/3eH6BUltn8F9pbQ6JrMBIqULiQ+0AJkdZRm9ZnFn01DLJ5QOdr43wUAnp+uI
jyFiUqy7tYa7f6Br/g72Jh6K1oeFC22aJE1q9TB0sfjGOgOg85RDnHoQm8ljMDcPFdM2mJbr6XYA
YYKA0ArsHsriwQTG1Lnqc2tXzRHI9AoqcKTGT7umFeZA5DKqXlLwDRBJyGKyZtd9XTpPX2h/8HId
xSXN+6BR5PHH/sUv1RmbL67HKpnl+hieQDaYJX7YTjuQZUf4+IgjvJjn28rPyIrrzOteERn2B10O
GlHF7bAMkdlgO4iRn7xyJjAGh/8A8OCJXJXDffMbIwDcLsUa+gJ5/Kv9hLjBJQhF0N9EXtiH99LV
bpqY458QxxQpH9aS73zbYYpnMoGnkkvn1wg4/ROqYggYZM0WIgDvSRt7H8auooEJKayKeVxA7Iz+
lQWbkquzY1NUNVz1vu1+SrhRQ0AlKAMBw1OO99duztVBfur9uaWaVsQQXJPUtllHqOtN07yI6q5P
EuAxUJrfzdKPNSbCtmOKMH1zAQN1rf5merv+vQyziHu8AAkCmaakcUXc/nE58QPPTpjkrq9nZ6E2
pvYUZ+Md0yoBMwB3qGn8utmas92T90Ma6WnjL6WJozCVedImx+qD/+dINiOvhdd5Gi0q0BygflFl
n+TKQYkyX54i6rEmkJQjlB79WLiMCY7aIEroWu32E8LwN9ouI+Ok6UYjVe4BpvNwpcY+NK4Ck5B9
Yjl4tglsK7v1pOaQm9coqhZZqry3qUiwtg1JTfmomtWBvFJinilvpBVZS7EZ5sSnmGh6hvs9MvNE
MwQ1Ulb8K/l3mRok1mHxwmvykijfLGQQ5QNQM9ZPgQkbN3G6UGRvSrNKN2PrSi9clhZrSTxNFXSS
X50mb+A1LHE6iYhrpj2ZoZS2o8hyWUP89YkSlEPMBqF/7MkBpLmDqC4vYdsKwVve6O2yPRXpsXxB
6jEY3gF0G3o+E+2Av4q5lN1iET5T+ajQ7vEdPyVPvfX8283iWJljJU/PgIyZbnYbm5rmcp3+exiu
fD/bqBx+v7x23gHhXl74yqdXUACu9PeItyqfWUhIsSnwXYlBRre0b4gLPCvW8r/xVkgRh2c11YS3
xzjiRwakbzC8Tn9knhWrluC7T6FniUUjSB88D5GS6bNX8BKFukpWNGJIO77U0nH7OU1L78MJhIff
u1yuAItespDjaim2czhO7Swi/S2WmCIWeU4S2bdj6gJRo9PV/+7+odDsXMxH2h7eiBg7A+Uv2Iyq
66ruDVP44U0GEHj9g6syadzEOHqZ6OaaZCTXBSNLMaKk1IamEraaJnnGfmpN9ijbyZpD0AMB0Qnz
91UhBbhADu/mdpjDXjMDFYPw4unul5t61NoWJsFAUfdIaBeB0L2chGjpGsG1mQbX18BI0QSd78Is
kbvcFp+YR6KipD1FwKYYjLW0cII1b5iKFPeLF5pThb6VTUTniNzyZbjSaIUhqD11eYb5xMkPWSd0
t11WsPaDe5lsfzdnk2w6nCGaew01bCCQLjo/YTBAQBrsVVgeiJRNLhz1UOdPM/kZi5TY6SgSc7kv
/ZIy1rWdkwtXwucToGtrhH1iXPuXicfE7kchUf/v02bRg2X0l/wdsiJbDFs2BmvLpKk3/aHCUawa
7psfsgmfIjQbLV0EI5q1kZO/PBVnAs1Wxt4AJI6V4R7j/NW38+tmrkJ3M3S59T4MF5SeTLjnjWeO
APL+1O0KJsIMh1tqDLHEG/kWJGb4xwCd79OUTFRx2bJTjSt/knr7ECXFTJshggJJ0rLhzC+ivOuo
7fR8rvdS8wFaW4lBOOHRbb7GSnxxFghUSTmY2jeglWTegG4FV7YyLNwVtoFODFcupbdKTbIeDPBY
fFY/kP4sJMQYdYX+V5bnRXIVV4XspRvMQh0ZTbuOkZzuO0bkn17Nd70zFp1MZ4x081/w8LlOGYSO
VNxxFTP8PF50eQHsHwF6DyGJoaZTQboOCDudHE0KT25PLwnrjVTDknqRWJ5wkHgUtP4bIwrrkVLk
Xd5H+VOvsFGt/QaD52otNL7ipdxxTVBsqE+n6cNZe5Fa8T05pUJb7rR9tyIfWQcoVuO/spMcMjEo
IXN95fF58jNIcfRme3jQR3E7FmVvO+phaLugusPWAKjHlXvQ0JOHzPwDVpWgDHsxPSf3KhG34xXE
SYN8vrDHjvKfYuaCoUOGuYVOt5XS84K6GyTmhVgJTmiwAEwahyV5IGGUsHcBDaWn95QF+2n0Av23
nOh8XKKgCn+eNVPQ9RTVi7p5YqPj0YEIjOKnaBuDl6CrvasJC9T0YWU+UL5NnOtxMQgGvWmcCsNb
Z3fcMHUfnpEGJ4dCP3RvgDMmEMpQWbfEab/w8AiYsu5T2jqwo9kR+U5XYJMFBd+EL4RXtyvl+mNa
2D9Va7aVrPCIjBHgvT2cBN9PZ0HCFQD81iJ4L0RMeOT+OWJRtxWpO8PE8SZn+zM9fISffaC6rww4
USOTw16Bdbm6bJKL/ap8hqzx04XcQaMNUzL2YRyJjxThZl/OcrwlfBXBY4UkcUvyrnZuBXFvlzor
NVAUpITUyyxTvdm6kxwd5Xiw2ZRyKEWqOGMimjHqok7BHzHHAKI8Y7rO/8XOAwCbVR/+DBcfMms3
bYI6tBDqjkEKRviLokxw1Rr2W80/GvFTa9sGufzBaYifNZ7k0H5ihCqyEPKCYDLUtfzq5IR67PGP
TMtuSUbyZkl3eh4nNi6Zt1soJXF7ctkjJXreuA2pCLZzP4lX8bzlYNYEAO//j3qVYu1qe17LX8o/
jJ8fhWYGSex+sTBysPKBLmSZqkLAxEABpj+AdEqOK1JSRhqbFF+VMGZfNrIk4+XeU9wiqe/7y2pe
C+9WrPhN+a5OjxTAVtWVCxDlTTlttxvpsaz1X0sbdSTGlZgR8Z/044+HqRyKeOqgf1VhnthZo1d3
hRID5z4QGjpXblxH+G+KtBA7IxyiK/gFA8rKbUWS0vAQvHuBt5ssRld7Uck/uwyHLpjNEbCUBkZs
AmqA11rOUO1o4EebT45zCfCnQTeXieA/QHMlRpEVrb4aiZdUONkTQe27MDiXbImh5AFsryD9Vsl3
Hru+Adob0KyzX2ZUbl7UECUHBVBcTFHvaNAXnUJYybCZzFY2zP8QuZwh88Cf9ZUxW2Oj3vkeganO
bDJoTs5UKTWih5aaR/Uqidpn+gETwlqaNP18RArIpe5VHcX24aL/ZCeOVyKcbymQs+pJBVJ/pvUW
KTb/M/Wf08Dyqv+asW5vBmK4KMbYVlfgJqhEAk6kPvMZwUb8yjQx3yZ1E2s+hsz64Q2jG2FR19Mh
JyHvmY2TX7vrPO1VWMuYhcItm625e7lXGbX5QkFBuA3wMgWWZsWfNq1fkjy3Mm7txLSg5BO3y/LT
pFC9EcwlJetiRE2SEJh+JOkvGDghKzN452foaeCXzg2o0b3CfaffqzYCfhbAzaYIOTbxch3W2uGc
bOO4SWJZZlkX8F1h4SawMbPJ+e8HXr9mTwXrWqkICPvfar1uNW/xqxMjZxK/s/2b3pBvW/jiaX27
B8PDQuGddJo0CgcuJKWc3txpJbtBOmr82+9V3uDxmfAoxokbzZuyRFVqMdjb60MJfZuUJuPnSsFx
WAF6g8WslZY5uTFsr6NekQno4Ow8EocTGzO/HjVKUjR/uBE/3w7kyj973qpCZTvp6A6agmvvrxF7
mkNpmRUvl4Quw7N5NXyYInTU9kv+QbSyw/V+0KPMG5O/p8D314+vHYFeMYhdUOyMUggDIXcK0OKg
9+Efh+hutuy9d4Fhzjob6aW9asWEFt6QxD9oGWHsvRS9o/Gq6ITl8vtxEWoUgn5fcOw2dRPnGEj7
xOL4XbYZlc9swiVYdlPpvrGN5jcEmXivAB862bIjohIhGytJ9DT8BCcr7X7rFU6AA14T/GUHQWGG
CghSZDft6nSEA8OfWXBo0d4s+of7haOzGFQ2vvwivdJEwgir1W/utxPck835QaAfD8dSSkCD31Pg
MbsTLwdoVdQeQBxdEtgKWdJBCmC9sjo3pSsT2vn4g7QJApGjFA66vgTigPD3R/v6CcWYtkJdj/jf
evyM0d7b24eCeBp2Cvery8hGIy/cCAwBniNzTqT+6/06Tv7kOyqs3EfPkJUM3U9CA+4Sqq3K5/so
nVC62WZHlwloyis5NoFAaa46m6Y6cJEqw+tVkJgRZDtkWUKDEUKUIhk+TMqKyFqswa6bZpFmN2o/
75reD+Wnkv0hRqhanYRwmZgZ2T4JFggg+qxww1RI9i6i3aVtSjoExStR4GODGfJlVlJwG31XzqDJ
eZ4kKbTGafSs+1Hs6h6Iy1BVpJGnOvh1SH83ym/xmM2bpS0w2zQebYGmahQsrbOc9mKgrJMqoRUS
rPyyWlPQhjK4C4FOaIP0opBOoaY+rL3MCCM3CAglV97BNoGi8sQsBtaV+vtKvuG0HGMZAXgMHzfx
p+uR+2W8K5FDMwaLqHC/ZcfIp4cZLG5rcBDyqzokLgQaWS16sxEczgyaIuH2Enn34f7u2j4qC/KE
CJTzEaV4nQ86HLDyvLGgpyOLTsCab2CLNcHv9UWIEofUXgio3WdDhv+qAM+mteRMQFWAlKPkzAJg
UDhVJdGCpHQIEI/4LTaSUq7ZX1z/fr9K8X/6yTaZI0BSvcJCdUs5HxJzNcIjfUqgXIzA91LuoiQN
b9p4ctjyi/FfICmTj5tAdnPiUlFj4jwmO7t5aRBkdt48p7bHOEdyh5QUV+vZ2dYMgHfTkWf0mHdv
Bcc3iWnJOHVfEkabEiq74ffxsLAhJcSiq6Iihk9WblW1NjcNDc4N5/U4XiXxtsasRJ6Jxbpm66Uv
n3VCT9P2SF2P7syQXdzHBKthQyGnWO0gul3gcSt447V+aMrHAxF672yLX2TFtQ0zE9poh3dIRt/A
6xk+1jAkwGL89qN0AJ9SttnFsqksgAPTjgFMADgNHSYzzLTq/pTmWqatubM7gbMN/wNakGsGf0Mu
t6pZweZo30biXX1QmvvNBdcz6It/QmK/yeCnlGp13bu+fXdRocxDVSMCI3L0K1YWr1vsuPF59qT5
CoIziuo1YUZ0hzq9kK7xInAHBBYLMDdcgBfBDdHHgjqyz90JC76UXxC2fRqC5H1lK11zXz1zQf2H
9FUgA3T3wtOME+sNcRf8k6oITxoBJ+WsHGqut2FG7Bap5Qos4aOq3C7zoElqGQnTg/nXlju7PHMY
aMdqFL5vz4fEuJyXC+QFf+T+1YjtkMKfGIsliQS8SIF2wtYuTd1ZS9nL56CgKXesL28Fp6TY+Xuk
fs6unCLacpJC4Vz6c8g4xxJw97mGhVYHJAYm7cP3n5FGMdyXRXqP8cmhM/l19nBa4qmvI3Yr07Na
6hl2TqV626Twq0v2P8O8BNpRaaDc4oH5eL5UiCjSlXti8EJjH3TCSYjmPp2sAPlcHEQMYeTNEw6+
YA0QpyKvNy72d1Q9Wf/e8AsyjCNUdqVGwwsiseF8wby2l5uC1CW1jUz8W5eZ5b/ZNlRGBkQOHbzC
BaEDUQ/0UVztNkytK3vMzv4oSWIL/sM1W90JsdpC8ZSDO4XyIt3amKeceHFS+SHKeW7ggBO0DOLR
iBYPkM//LZN35lV4pWDQNa7Q2TjQZkgYFt0B8P845aTp76dLVR1aqUQvCjBDKumzZu90U3QEeQXu
rshIOWEPiCrE69Mi72Q+viUPWKJvqy9/njJad6WR68CSjY3hzfb0Bivh/XGt5nPjpuw2Lz5DsUiW
nuP+/XU50vPvMJd1246OVirPfhSZ7Tl6w72aPhOdKxtwZpracg7BnD5h0vma8f5wOtPKtrEDiO4l
S+sril/tKbeER+RcspexlmfrJyk8pDwZDqUPvPxtBMRRpWZpgZYUBE6FoEfVpcWo90JmaVWv1F5Z
f0pyBaDMObtNnSYYfx644ssV6EqLRzCb7XpjqVnYCTEzJzW1agbyA/DtxmPwezAioHs16a435TIR
h++Vse8hcnj4Tj1h6CN4ZsD1SgjBILWTDB9GYp50u4AtK9d8PNvltXR3m0bdkbA5VHijHXUWjApK
5yTFYDPRJGEK0I3e+24YFATChsF6s7B5rtqQ3+r8FMjFxIvXn3qbQSYw35lLla/W1qGlxPA7Ryup
gY7ZeBjWyuEUAoo5X4qqqcS9urkfWjqw7gb30Qp2W5TSDSEzBvcbs4W4blgCFBUub47Q6P1Kil+1
oalpGJIaCoF6BB2IVpZGNGAjzqZmb+AVZ+JgqT0T9s9/REBwllJyx9Jyz13bOIrncSyznla94OhL
SzrkeVdJAkbtfUzX4ttNxp+EU9ROXop2wgYWUu2SmULnEGSlhe2auUWD9MzrjeDCRR5mSIs2edCP
HYBW4Vn7nmgV+QbWfwQlsxXedMf4d+o6x7fbY5pNmz/5vqssAbD4rQaD+iQuAFQR+jEotoUJUIZQ
IkpSuX2NeLiOaedWWprO3fUdh7xEjmI3FYlrrGNMaQ0NXcK95hkjn6cTT8mddI8R1h9yuu+6lf4Q
DcACmegVGqqo3hsyhB6M4DpdU1xsEo8yG/Tdmb3ZKlFR/uCMhLeP2aPzQGdcmcdQLV8oEgiRcYL4
ZnsRwL+aFd8beGp+xuPVQJjhOQE9Dz0ndrV51ncTgac9lMazKkUOmGIebg2s/oiPjpjlF9hpesiR
tBAj37bpL17GVQy7dApw1bkUxeHVfCYIMVJ5CUIuTYnXjGsNI4S0dHGVild0w6eN4267WriAjQD0
C9ICMfnJCGxP8Rd2M9P24GeMJSgasyGnjclmczygtaSFCiUEFCBZ38nHvk300+PUtnVqRKabo4lR
jbbklWWpl+g5SZf6ffcpvykssadOlIvSDMZJf/2/Gqy86NVFBQvvT0PnnJVOA5b5an/TYESu9EJ8
cdpUssvL1vFsToZqMQklVCIvGaZmA7RNWuuQE6RkfaGW/6iDBdNpJioeI51os01dXD60Z4/tQ1Og
DxvIXdCj0gRUbQX0Acd1BvMx2jcfn/UCO7Pq/8uPDXz/S6iD1qasrgleiijmMaZpZlgMA7Rtq7bb
ZGMV7LsaAnXfdQgWLKE5xy/iwc0b8F5xrHuC2LqmW+th0OwERlufPss5tw9PuFmucKyieWCspkJc
UP+Xohna+Y6U3zA+0rvM4Hqb3tGpftOvPGdpO9wfJ+Y4EoeS92XgAPDC3S3Xys9z+ePrmXG7PJW6
oPTZ2fjGAbRj6N7zkBPAiq6htUj+RO4cLZwGzRmGxupBKTPJCF2rqLAnmXWBSZo5fGMaF0qwWAkI
aneAv7HOjTKWqClKyZ15+dSezw40Bj7qNawV9e5qDoJnPLNx0szaj44d4PioH16KjZ+owNXyiJQo
inpbA8CaW/DS9KjIb/d4y1bhn5QnOGuUwM+WeHdfMBiqkEtCWAACBs5Qt4/d3/3+TTBp4DxQM1Sv
EkQWZYsLliS1QMypTjeN63CI/xYzgkOMboPx486+/vw6vZzt75UFZg3WOK8E++xW3dTjtdPeLSQE
07XpdoN5muJF0FtGsDISVJvNzIYje/pr+JgPy6n5ydr3v8ubnzk1rff1/nByK83Juszwv7IP/PkE
fEe8xU4UhXw+c5kYXulqS7y7zqf5zVYyLD94UIVaglRTlyPRDM4XTIc0G0W5g6VO3IZUihtTyZqm
n3FxzqUVVepJg1pmFE3vL+bgGxWgPz7x0DXmVA30SwHKqOfDQg0E0tBdD5L+SsfAZQSeLIKfSU2i
3ygBbEIFL2v3SxDc2z+x/jTctCSr9avueiOCE86D00QNQBbzIF4OOIFxxITxckE6rm8tnytQQaR2
pt8iWNHv7as9v3SgHaBIwHwwkUFThIA9oHdqoy+npJZ02xgI1Td7EhzRifeKbAARq7Ovk/VxhRgw
xVo+IchFv18EqcgRjVPa5zHrIRCcxOuv1pj+p6VH4HsOXT/HUiXK2b01jUVD77cfWTtT1PiT4oFN
NP5/uD7wUAODdygGpYGs5FUJylRnKNdOMsfAChEYndMqaUYBjm2MSkxSN1qAP1cOTkv64SLBT1Yb
js3Vm1gTqDJFJ0StMAUfhYRWxVcym1Si7BgSSMiAs30E6q2F7xegraCyEqc74dFLLng42xUHuwCh
u1EgjJzgk+aINqi/uIJId31IP9pPAA9t2Z9TUloQOI+Xg9GQYI3daXG0XRob3R9fF1z0sne0pacH
SZC8c8jhjaSZLutPMAd27wrwuDDLCvLyKXrxBNsCeqeWwfhABabTcXPP/nNU7LCzwQKATo1jHxIr
8JQGCZqOyKcw+takabmJAv1o+4CwAJmBFPcTNAnJXj4tWb748FOHbxkVglEFcV3ZUVbDIO75NUyU
IhftjEwkRiY9644EPMnqhZTK0keTr0dWKM2ZI2zCLdMjp98Gd1c1J3oXkQkRMsodJWBcwl5Yk5nW
dxqvT6WQm+NjW+bhMdAMz+S/VNW+TdVCwNWh93q+S5m6gpYQLuZxF0y1t45f1PeIKJyzxmJZO6xB
IUG3FSONzxi2n9Pv4uh7Iowbxq3z4ekAw61zqAyTL8/t1vbPzT4Mn8LDKSSvrN5yefYbbSbCTDma
Ga2Vn1UPjDHdlUGLhdJZW5/4YGn941Bgi82r8OXdXsfVmBmL8eV1vnwVI8p8ughqMUPX2OkEFQtG
ApAlXIAX7nXifsIBBaRvHBNnzKJ67oB3urj4myH90xMHYzC/48iqE40ebxBDpR3dsSKYF2CKRD8c
Ca6QcDhdLaM2FqE/OWVQHuhJ6KEWqunWyRLATTK9GGC+cR5fmDc6E9CoTLfXHYmDrP4utPhcCc2G
G2XnjOmKFCHGK7KEC6buZpu723WNFcd+/tZitqC5Ig+btsqS8Bhd84un22poIfuh7jZADo9WGMKT
4Lah8uzKEhNiPANDnjpVzXV3MmUY6NJ0vjrRbCdvtY8/Li3tYDAwjvUVRpoMr0jilBPqtIbsvkvv
qCfo4g5PhKZNfDo1MpessK/mpzBb44ckhQaNkg+gq9a7qRFKM0kUl/TnCaGNxNG7y6g57rkmX+Hg
EvZTClmXzk474eI2tmW/N8gcfPG2Y2SBdssfOxyNTjIybjasI5utymwhNZT/BjSWnuzUOR86C4kD
zISqYMiIyNsnlHyzOH1i22xLl0fZVNF1RCQdfiNUdLw58rq14y8X/YuPQnvt60qoKbvh5Hg459Du
iN+96+RMpz90KI4nC/4JovQr03H80IcEbMxyT3RPD7mw57Zr+tOZxJZEuwl66CQelbrfvCiCgSWV
pcZngbNDmy9vpdcr1jSC9CUdjyBr2Ukc9BTHOC+GTTD7V6FbXFU7c1bIJT3Re1zKAlbllgODVnxM
zSNunDHZEsATwcq3d77ByL3WkYD63pS9qZkQocCBn08Jp3zvCtyIqXo4AAS1LHq5CJoLrYLOogY3
ClTIWCYtR3C5rFm/sk+wx30GeTqmxPW6CZRYgUBqdNl1uHDb+rk+uNvh3U1pN1x/n4AlwfeDjfR1
jGp5OG3yZR1qaA/bGRuj8uoOHAuGk55qgdnz6WWKpDA/jydYRjwSfb5wzrftPh02ZXF9dVG/Wj/r
T587ZwXHwzU67B4IPnMkx+OW7WoXyd/+xQFB2JPOT/VmopeL7AOz7G4f/aKXW15H7+Tm4uasH422
s27L3Z1PBTf+/YwkWoj2Kt0VUx47gRUGDGI0hXa/FZnk2KK3rgYsdYsCgbhvxkeCCM+FT4VxwDo7
h9POzKwzp4MV0XcnB9hmNCpG91krgWZtWOZP+EGrRgSmU1NG0nQb6sYIDrHnrzwL2N1ZZHu6qXnu
CX3W633afAuXWglWXAGi1pYWZdKKOPMrsKyHR062cN/GWNAn1+MIujcXGj9LaHEN0JSJQJ+/ibKR
L7/IsvWxA9mvZQ4t3LwPDmy+g/SsNLa9SJUpAL0H2YMG+TvWrxoSNBXK2iO1rs8haelL4BxL2IpX
8z3l92EvL5CNLQ6/eOE/sTe0Z3GUer9jtgsF8/j+IRwVhU5Qy9UMuT0cr9ZRH+az4fDN/9T2f6bk
40thzSLz74Z0AzL3QWW68uTfiSoqnWJiIkdIN5Fi4oc7r01ly8Byo16C2LvNbsawBq8x/e1win8V
sN0k6D07vn31EYUZRnTXLvIeD73UYXe8oGCPS53rBtNgLrXqL/EOameJvEX5fbjI7SvjSpJGdw0L
fA/yzaLt2JvGosIxVufNhRbU3Jnnaj+oiSMdq4p6PdVDJaZrKwf6FYZSUrpheOgGCv3UYei16lc5
9oZJZoLyHyEwajHcGZMEI8RVl6zYVGxO3NEavMfuwQXAY5mFfoo/inDE108lkcxwf+hfqgZutMC+
JN/ZtFRHcTt4mVx0Q+bVyrTzCBwUayEpeut0y/vhdhZ3GfxtXiKCv+A+YZH7e1zEVj+mJS5Tvfgt
hJMLRD62/y8mWW/9QPDr7H9b5lpUbF3D52X9R15lvoAzIMaMRBOsxitRRJJ4krbmX1n5bxydMmoD
/xe1xWJBPjSWySSE/N/d8yoPbnjEhl4vOiEFn8dZ0BTSot7sQ6gzBFJJ5HMwd0Sg372PS7R0yNtT
QQ/bIcxkQbbivjvlsPFoqJo6SGqGMieKOg/tf+ZLA7TS8/kc0k4PiPHLkRZX1Zdy+qM3vWlSmNHL
OVCD97qjxdcuNE/+ewqrvS9VgVxwG4InN4T0enDCJVyPCJNvB0UnGZSpZfwzgH0us4k2p8DMk5sJ
vB/xofz8ZOjZdCtwJIcb//zZjt7eKGrVDL/j6qkkzA9IZtd+kUFQNgu+vpFXluOOJJbe9WI1/9WY
mYTLEx+fGAhaaZ/YTTDUCP3oU3n1J79I0K3ZaTmYWJ0xdpNcMD23tadDqDN7r96ASu4hQ8uYkVwO
eGvgnjp/bQSgZVmIf4WH2WklytDbnKzcqYWU4TdVTUeWDJVRlmAumQQbsKYoPD8JJiL4Qg7ur6bA
1rB62CWdV+z51ht5ayqXPyHWzkP10OWiou/CmAQ00mHYiqwZEfLBDPIfFDfXiv6jfghaZmx0y+T1
9i6KP063h1cwuGTiCU1lg55lGZv6Ofytjija2D3d0f4YMo5TsJ3dbdK5FWhLpkVVnSQQECE0+Oq5
1CdiJzXgwnV0/S3XbkEoS/Kg586EPdg4wnISjGCL73Rq/iFR/DKljIeXvAb9v0WZVwuPR/oYFrzF
FhRmX72J2wHz5yUp6M2roJ+1XbQ+wbjIt+pfziMJBFBUhT2Oohl26Y7OqHwbkwlR1ZuE2eb/9ss0
MMGBQyCaIuJh7b8dmr5Xrs3EVRFjoVE+AOWKQ9hIL52VjpkZWkGMKFq+7qsU/XjR8Woo/D+ru9KK
EGztR666xtKxYZkdmk6oGFqdU3KSvz/3kaYgM/BLCXRvGxKJRfrZcUdsHy6POo82dmY6zaMKlboJ
7xTQh7r9g5dzPqP7GdEd3EOWKdRkGeiXECYBmIfDmWx6MzFmQMTtnT7n0aP8a292IDLGwD3pKiaT
GMfJxwxPtpTzljO47pZMpxmMd9Jjtm3/iRGAEMFUTGlEVYlq3ICALOrLmHdvffyFHDrlPFhUdAqE
srv64wX3WQ2yZpaQ8gGH+sVa8MmZ0dxMss1YDtqoplXfZJU2SkZ1DxqwPUGfKS8UGUgie81IMAD6
lctMtM1eGzRrvCxPzPsRXYTyX0K/CmVO8PkuJMbuOO6s/5Qver5CYBYCLbPi+FPxOUczTutZWWdk
fhKW5IU5POY9e+fq2lTAjdSbpwbS2mZIMQ+mQOI7E0Bf82XaO13BdHpfMkNO38J6sWDLs2BaXzN/
ygbOFgSfmNxNbWFrFb1W4FKamI21RXUJoIpbzKlCI/z8/xotf7Bs5ZtBQ5Q4MEEHWintBxAqEPid
9CAUqMhyHyV2N/tiZWzeb2ZzU9nPojzdcXKnQ9Ru/mppR6d4XyVx5/zCfEWSJmnIypHhPJepkUZv
6Ql0wP0L/4NQtTLnvm1H8QWzmdOmFoA5iUl2CCqh46mTwYwvIoGkgxOMXOsw7gCFSQ1JAZZk/Wif
M1FfoMY1QaIUrHhzO+74/Z3x8fRY8HvDWfWZdGoyslNQg6Ilx9j5VkMIdi1ICClD/PJXKvFnwOc5
3AKyYKnPyk/vsXIcnW1ZVz8MP/y8081x2b+3qngq7p/wj//CqIbhhvhsgTi/6RN1AJOMLqe1bgzB
oCyuTWHmguylq5EUfYOC4QH0ymu7CZmkLYHy8YYsnAdpE5VrbqeKhDWYxmC0R2B9KEvGcDGXyfyl
RjfIuogf/4prbCCyWAV1f/28dc2owkWiDIovZajVTj+DNWEj157xQiDgBXDEhzluo8RE7uhVUhIe
5FKVwO3/0V1sQo+ZvUvMiGzWJfydx2YzJ77CcxI3sYYGAQDHjQ0p2nGhoBTDCmugDOapkXiuGRNE
jKtTIEY+ga4qjY4qwMTBW4tH7YaROTmQjpnLhVIwhLDurkRsI+qPBfBS8/c/xAqkBuCIdjyrb+b2
mzAS/oGehVgM83aYVbmZTomtn9bcLIk3A8QxbBtiVa6ynWZrGtfZ9sjjvG4zuomeE6IBH4JPmgOt
rkFtf6HfkefXPQJHDq364OPyW9zLC0Lpynf8rAdqBE4eVgNF6mUbRo65H7P6UTQIPyG8UnWFJlU2
XpQ4sUaHXaVtHJiSnkkbOSEUQghiLqzf9FFp34H+NLmSz7fAol1UUjxBN/46eHRLPwiolCnjGCyw
m4TJ18agRsnFWmn4ttAIvFVb/36NZRFnjqMb386OrIWYr1Xd3yhh3Ze2ewET4ZeLs0Mn92cWNEaT
UjLEGltT8ZtS81Q4+c4VDVQJfkwkamsaOw4C6HN55CHPAl49cm1KLxE44Q18m1Eg52xM+tLrnnkb
bsdrjxTgUpkrKCJnDmtl0phhsOieibG8XDt79WsY0G3LqMWapZoq7eswJKSDb81N9Kmwzy3Iwnpq
L9V+7abZQhlx4eyNUWapLyTG9o5GfqH4F3aJtI7SK3bZODepaWNlPR8vuS05JdzSrJ8nSgThrBkI
XhGdpqinB/UvRsnJibHxq50RTaoVnHttFp34PfXEiYdBrQ8olDWemADjzrsCM4sxyxf8FAPyNEsQ
PwVG4ABzwZ17vTysyS66TRcDBoNSyNpdWkm7fuxXbps9i06vzinQ49K3d3lv6x5SPV4gL9xGdTbU
/jXu8tyvQaow0bL71YRQf73Af1tCChQCzpDI0k5PTlUrSIDtY9DPsoN70LL/zjhbJ6LYFmrJyc5Q
p1vFpremIBYcKoRkD9XYCwkMFuKeknrzpZbREisq5xcEjh9VgpJG8sAw3SiIhZ5DLzsvtQkd37i3
kdSfhqAzTIxdS40ZVRecLFOpdpQxX1k5qah0MOJb3JFaoOmaZ5wxpJYckGxpoO72CI9vrjCk47mb
Ou6OSmIuRswvzCLiEKcw3GLHfnyTNIyenwpfoPz554rNyBPgjH0eQGKqQHZvWwMO9a2S/bbf/ovH
Ro6Zh8H17f+p6xAunUxcRkipZ4y1V5/jr68KyZ9O4joTtGrFeOjXQ9Ku+iFoB455fStPXZBBMvdt
NADoFpzTZA0R9DzuG2IQAIYbDi2coYx1BUsalSBni8KabqRyg3rueHfw9mVWE6Bh2qHlTik7yV6h
hcP4oJ6p7QawxbAPXsht2xO/IjoW8vkad9RTUOjpbrxX982sX2LKM1WLhbhrhJ+jsWoEqecc6/tz
s52nL6OhhnCGvIUSoMjgKFAz6gOnNDqW/zwPG+STiIu8qNhAeQi/niWZ38FhO/QNCSh39CEVWoVq
U60rOstpxp7Eem6GAb22LxeukmNTwIbzxOPSh90AjdwJQ2ewyFykRPp6KjrIcfDcJ39k3bPXJDch
Xw0i1GYJT45iu+G8AKwAE1oqrMGhWy7molRt8GxfolSyDy8CbpsQWOkm0ZubbigniF1sxzNAHWzo
ZFbCx5JGa4J0ary/Urw3AztbJCbqmCQHqPhADlWSroLH3KobDliLs0+xibtelhh8JNROL7LBGQ1h
ATq0YCIYsOBoQaLmKbYJ1ckthLe9/wP9CIwMVl8E+OnJIAb07HYQKS9hMmVALfDpCTESRxplNMcE
agNRdmw7Y9cgY+2Ticd15dGqrrTpdZ8UsWdkEUnn7RCO35am0AM+Tpqr/qSoRmpCQpbALLvtbalK
nCmd2ByDVrghsF0TdAA2T0X7sla77yM/NkHisyFBAhzrwM4Um0MdR3Ff67oKAq/qvFMTkx/UQfwg
RORGspjnRjXSnpIkvZxbF+MfTWkONgNmdrP+CXYLNRwqQAkJAHUeJoJv3JcFiTRl9L7cQKISfgxg
96peKo0ItKYwbKa3ftH+GHDQfdh9V6kguH/EdL/AcJ5PZysHp3Q+NAifSFH/VABJwZ9EE+FOaQjX
l8HFw5PiVWPEdgCgk/f57mekO2+JmV43ZDO4ma9v5OmDVg4snPXPeexi7dA5RU8VOcnG+u41Juw0
XhWDvg6xBExAFe1FrdzL9PLoC6YIj8dupjhVOdMZDZm2rQaGrI+nBlteAzQNM1yd64+wWmfvCy30
RR8i1iVJDk0tFHHYZiAgGFf/MsrccWdo0jvkoXhHGIGfy2iCA/6IvZygNSOp/6thKDn0wBfdQDfM
1f2DZBrucHIf3IDFHUluJSiLor77ZnJPuco9zrkyCop7XfQ98/hwYg/PwaGsr2pxfwC3RyjTRAJ5
yWw1bN7JluWw9frBBVfpalHlxIY2OcpcImcSGAh4nHuYTJD1jd6HGLMAfWovZgWEsuLaZvAq+q1z
qeovJiP7hMGmLaYgtm9cPjYX6gcC61jlao9ZCE+tEJNIdfz7OFB2YAry4G4PY56S0QW4jxwNsPhB
IghNxK0DrBVkcQ+VpF3g9KfXu8NoViYeCoqzP8JUZjE1AyIBGeA3AAPeL7yDd6DSPw7x3Xu1DSlo
RbZB+C60RO1MSEEaU+/uBvb3BHgHSC4bgO+5IRCkrHwVj/Yg8G9Kl0GnpmffF+JNuWvQc6SOQJQn
6JJfW0zkRHsjn/IejPAP9V9hYsfrmxPoktGQaFhQglg9xcesPmLLAu3BFVGIO1sfkI0iguelEl4T
nK1JVNeIgrxCJhSiJPMWgm8Ir9GHLq7dEWoOpJgPKdZAs6pXtS69KSojPDye+cECrz3L8as5NVkO
pN5tVyD7xKm1ZU07tHkOcI9Pa7emg+QpmpMs1AkdlAJuJvPfBLrNJbdBCOEXmZbkPPkK4VfkWvY3
ttLGo7MKbkpg3N/qgotHSpz0ba27KGI7i0f5a5pILAQvK7zqekd5NDTd0hFDVtyxDHEwJp3oL14B
abXaDZo6StCDCP10fAig7QZs+OrdRWfw+khrPzuhPaNTBY6IuVubdJ0Wx0syouAmdRjBtzJ6MN9c
rFNUgqmHH6WipzxDHaLkYMZnVN573/mTW5lI2Xzw/4iVfYg3HOW+5RQnswj/G1FarmbBokz+r4qs
VUruIuL1bI7TSth9/VN5eUHUhj7Dam3ypkO3RtTfIeXacWyARTBQ4CeFWStOqO+1VZOhzsw/h1f4
LoAnquarGYBVryEHGgGcf297Rl13uQQTtGDHyrR6ymXpHDzT9rXR2uhqSW1KelEQgYGis7lfYyhj
R6Dd9GNeNdcpQAWjK5CY80O2gIKLISqQ3UAOpaI5B2pWY/LzwP0rKiD8xkaG8ctVnhPCBGYFt8jh
RSLYMBFKUWq5ukuMHBgeFEaA5X3697JOhIqsTEEdLqUBIawKf8fCqK4cxN9OUZ2ClrPkhzba1Yza
jIPnUqnwb85ADMW31q92i5t71nNKWZyiWkgC9E2aFnnWRZNKCM+CjVUxB5mkctWr4pThhlfElQc8
Syj9EP4IJY+qWhEy4xDEPfctgxSl5FgOCBZUOI6GKUAYAuGJjqW25RMbZJt2PzvjxOwVy4BlLvNr
pzZQLPqcgc+P0PRjiyWmY8Qk7vS0cvI2ikGq5msjDfY5WGzBHrtg/pztPWO0V0142lHNH5uKEoVc
lekcqIvxOEVKhD0oXk5uAJ3Qytm+deHHOgXDIA/O2ymhTt1DyL4BDWVVeTJrpAwAJJXwpN/nyS7+
K80s9aQy7nhWbQaR6FyKnT/ErrrLT5yFcDHjBVjVard6LqgTN3ilfVSnZ7bM5bFKBRc6i/+IrdeB
6UCcwXYRQBo8LCQOSYkaLr1NWVKa7WwPzbd8CUwvbvPjjf/0WyUveM1cX4XUJ/bVfaNI3GBQu0/q
FsnSdbUWOodTPuvnup7q24sGXDYwcBw1kwiQaotiO2QzCFwlarKsN9yj9UKZBGnr/N60bI40IODK
gDZSwLk8Ggxf1pVNiXfRqsoXH/YNP6vMjRV2MEc/K0M5FYxpvsxPzpJUcVBrCoYk7goZiIhrC3ah
iWj4til1uUjtPJOQOj9OlkgK+LpiW+nGXLsnBaOEcmpKzTZTaIW1Jl7VhD0CNfwfCFdZzzvQRDPz
SAfHXZVmieD7+DDTv5FjKqWmnTerGP2e3Z7oBTseSnTDAZZhilNzxPzuRTYfwYPfpSiAiicgMB2G
WA/WsPNvcCFv4lHpw2T9Vq2E19xFTuaD4P6KTZCpJ4VXUs/Yf0tjD0Np+z8PCTwCbUkqjA975Lnd
s/vUVFsFyCJskAEnFF2z2GbdfsGeGwyB+la6XIHt46mMk2Mkjvnk3UqG6X38BzlJh1f1H0JsnvFe
zg8TtpSqH9BH6bzWvql0+o7GHdCvD4YF98xtH8cz1+l29snKWJX28gEXQLqgBlCJ7z8hdLmV4/wU
bhEN9Y0GXO68UHNbPpMFu9QPe9UkI9+yBmF78taz4SbrXzyKLz644OIH/F22u8tI9ALjLb4FSrue
HSBzAT7EFrJtdg8bhaGtM+dPTUwd4ynmfXhSAqWpeJMUF9o8szatrhlH22AUpFviux4T4JtVHwgo
oAgPBOpb9Rkza4SrHpjQDtCFte7ncCEKqSPbL0KvF9A5TVm6JCKLS80vRbsEDme1WrgnPjp55T0+
4TBjwl7gBxH+X+xxSHZN7H3ZmX/wQnA3PR/OqpW69K447jOOQDvFF8UBGBOdOX8r9qZIj2hO3yxg
PDctCTlbOGrdUvIfxgvWPZtsh8rJ3REzVJWznLBfuXDkpfC3NTqOGZxgjgZjPCR6hmg0MeMcV/0t
Bw0OYCcTxoBfCN6AFEjyLci+ab7jU7/8wGy1xFsfunPDAspO+7at0RzFhXBtojUGg9lLb1KnhO0v
A72e8S3M54h3Vx1tsVbJySNZ5M5tQ8nX83ChDLskZ1mBdD6xdbERNOlRf8HVskitoT0cPPbRYJ7X
/Wdth97zb75z1evBHnnGLPmMuVLzKmBL3I/dQBwA3RsC2ovrmyBmLIyuddh27Ri1nVV+Ca1omCko
mZmuGqiALUVUSs2p9qAQCa0yraP0PY+9rVGsU0X2pTYalt33TaxF6E69AQZx00/YvJ8RKwdGppsB
5AXgIbLGl+4LGw0RlH9xVz4CgWwaaWRjh/DTy3N6HRQIFwbyEaKzXZ2Bmgyw1nhQmJG0rYeBgCfF
4qOle+H4gTgnm81dWkmVOaUd10/qCcmAzLzj3QCVSpP0isB3+boQnxtSMvqzXw8JlvxRhLmldU0D
AZV9VG0rxnnDoqJorak9BgzwzmVCazVrGynb+lVqnk7Z1HwM1iSVJTNKGwR9Ch53/BO/LcRiDr76
AJ45pAEYKVQZgRoK+CknlM0EmrtM1CE+dUWdv1CyJ3AS075a7ekGImmrNob6n/LjAJoY+JkX4AcQ
V/dmU3+06bjfDCg9HnNCxqUN9pZORrPqTsE1fWnvn3EiCWBePUhULneOam4rdWZZ6vU+GyPUgo0f
YAURgCpLjNlu/Q+CRVZv2gWd3Sct4WvZI3EZOzU45t7VJHrhEfAbxXyEw0ss2/9WNLk9bCqxlni3
IB/o+m6P1YspPd0FVQfqiD5bCQvnrvB/Ym5AeKv3UvsGy8kfNFAZDD3goMLvRbRq9pdm/U/NC3Wm
PIoHeetv4KiFEUtXtbY8Qin8n+J3qunxmWXWvYtk8UpllChzoZGYmBLfCafZtJiRn7gafb5pLHqZ
QuyNt+jY4BTyBbspSIqiF1nDTOncb4n0aNZIGUu6+PoYS21AizkXYhzALBDNkZ0Gc+E0Kdhu7KKK
BPdiSSMmuZh/UNTLS2OF310wbIrp+n67MjMRcLwRGCbO2RKnpA8arnK813oZELatKEu0BVltroJF
qlrmuScED+9dK1f7SZORs8bMSK410kO+udroPtxpM08VpI8slnt3QtqFLLWqfqUzPziHq8+yVVxh
Huj76klcY3KbH7kTe5xXjXKS6ZvAzxGgcmM0FEiBFvdFjJVxx334kcfya55XoPSeGIgAOArd/Vnl
O6kqZhkBGgeGxvdvmasuVommO8PAKhfWPrLAn3uFAfbNIqLIbOzsG68/KNEq3LxXGxV9OoAa8UHa
VBUQRB0O/0UT8/OVe6+kPotiGSTobrkipdGaFrTQCtrTrJ7ibUOIIyTt8rBRuseJ6V8OnBvQFvwr
bb8Oo3dvAHkCqdCIXGO9YFPg/UXwBvzcYuQkYUJNbjMrfpUJ0OPNqYhfDfvp1oL+Ryx8kLA1+UMZ
1T1mOe/jUKOV1UD0fga2RUYP/VRw3XpikOTkVYGmxxGfnMcXq/rMaHG197Cy197c028hImnLDNQT
VJrRfEUJh781LYQj3loVIVZtPPJIr1mBR9WFgQUZXUxQGPoy+bieb1Qceh2VfGENyzifIvamnUKO
kkqpAS9SEyc9svWaGziG60+lHF7bdS07N9BOmqzx2Ok4tLSokoYUyrHF7CP9L+fuMTJBZo7Rv7X4
CtgU7hALxNu1rk5NZPliHtPaAUY6h8+y0u9RhnDjQ1GLsIbkCCfbW2vljS0Jwuh3LXhCpmJuyCAK
PEjhsKAHpcMR72MQi4yresuiYYK0lnWaI++xZ9nYcrjj3fIraW1ZfPFdkm7zGHcDVhA2muMbvtLA
T89nASZ9trwVEidVLL+NAT9KSzDTLXhoGMYVbi94pmoHglVzEarBVuhiO0buzrdAzHdzbb8IynNJ
6jeoqkqwcuTARGfMtgUuz8QTeXfXzFR+PKownnfKwVRtdnZ4S44Hl+z1Cc6ca90o8eyRMdYXZAzl
qmI0Y/rg7H4BGr1l2vaPT1C36hJ8w7UeJ/FfNM4N7IhcFfUy4MWvq6Z4i+zoDPR2Im7CS8threRH
tmLldo5L/W0xZZJWUmc24A2Jbx24maKLz62NwBEsiKDtHjOYxJAYxZa1clawugn90L608TCkLB67
mVD4NTGxSWYcM/GzYKLZ0XoV+KijkKht1OvbIMwsSywNpaZqvci4yeIYwwlrnbkb+0uOLFSZuO47
NcnVY1KlN2gdTVKWLUOtNtTYfeuKpV8v8ZWLuK5rfyCblsi9C0dICHwKa6JOHlIYFR9rEGSaxuj7
laWrT0xHmWXgWpUytvUly53omG6csNJB7G0xHv66iZ57n2ZOxEsHyDvJPxhCvz5sx7vbt2lxf8eb
sMFDIEHfm61Y4yg1I7m45Ru9CqaVhm8JvzM9QBy0xJ2rO9cTLJQV6COf6nnSHDIj4zWuCgvYh11J
s4k5HHPDnhOYJSuJqZhUfieXT3uGLIWPjpaVD9kl4NvVk1w0j0kZ9753GV0NnPf7WZ6pVF6cRYy3
oumXJUjdeVZj4mN8qEdIZmQz6JIWd+AXvcgCZU3pKLGhDbHzGC8+h4oPguBtdWD/rABl7noWR1Lu
QuxG29wpvy0v/La/L646UIEErZgStsfcdqAmDVot+28eJUWeFGtZWTHA5APqPwxxXeEW2qgsYOq5
DQpK/2FNDjxZATZClPD+UVwGyRT0xx2BFxsv8y4/vvArCySi4DIf5t+ZVcVcEPSQf6idEnxDb5+L
aA1jnHKqyHtWLAYSnfmO/zPh/26C2ETRwnL4nk8MIx9r0mxt8kGDPeCWDkNFuEOCq2kQd0eOyCtd
XSqSt2nZ5oedELTzAr+HZabxmR178AIrgEnZHSiHsuACaR93a6oboNu0hw5pOq3eF6Q0WYuu5scA
n6d3/JkyYpsckM4vRwx/1iT1eOcmv6sGqh28HtZh99SQnDRNqME30ks9+HzD0GX+2SrjOlMZjPNU
+uURrqUZTGMhvzsC4x3D0Fd+R/t6AObLWGsas/xVg8myuDcFtw5h9ProWGOvKl0KhFccQmSw75jF
XglkcNWCARZcC3bpQ1ymw+1nFOFYC5zBkdNBEAa8SKTR6fMM8/1jKjLWvqqijU+dADsWBjvkNzWE
iDSxb1eKzkS1Jf1oF8WPj3xPpcdlsAhve1iimsJyeOjvZsCdg9bsnrJLKKO3y5oif0HqHWXwrhBV
3povViMSwG0EnLov/TOPt63xiD2A7EIhmsuaPj5CaGliBmDMB4fsnc7XgR8Loq5GZDdYwoFkh9pW
8lm9RM56al8Ta2v1U8f53niUISzYL6Hp2R/TR2VDv/L5b2WAsTZyU7efasUgztBV8vcNYJcbwmgT
mfGAMrMvRqLNEN0JTx3Sxwwi3ezj+cZ71mITJBYeHHQIGCAURhOd1P1zFOJGiiHWeZJvxcvttAy1
oCcNpu8FP593P65HPJ1wkCpqp38n6Meqi8Q1CrlJ7Xu01nrEFD8Lm32F7w/5gtOV3T9BQ53oGNR0
5DeFoHygeqBOPEQ27Hb5MvJkJtkV3hjo0w+RSEOb1OeF5wm2E47aNiv7+8eHKkWws88LowKmHD/N
bHHltNN3McNknD0c+HAXqoZ+ewjhr2krbRolia6RRXmKAnw//OPFwoz5KPZ9yT8P0E3hNAGWCsgW
1pHPpGK2aQoOz6/Cu/Su62sUppmnL2SkwgV1pzL6tKETpV2P1hRgkkEjI/yX6anxp8LSE5Be11Ma
dn6WyZkVvjNXj3ai+6Z2nzkl/57qVw02O/RQdhI1+1xUZsBENb8wgAzoV7qSrEAtwH7ibPN2ePUz
vx/JTg4/vQZIT+2z7Luoiaor7J5ICq9eyiwLW/LNRV4tT1gotzTR/YInOoBdZo5dhYeSuS18flWn
5UUQX7qWz75QP/i8wDLgz22GmMvcj8T4UrnV2urzYgtq6Wm4nyOTFIgUuL36wn4/pTzhERfZLVQF
96lZs2fD2eDnXVUq0F6oIxPe59q8xu+4+PKLxFWAHa4Gv+0Gm36p4M6xzBtTwuuMD1SAKa6k3nXt
o/VC1crr54RUPIsiFVjHhJBTqiOJjc7r8Y9bRCKEh8zSkmoy3ofJ+RoqSUO4yf9dE/teYXb1L60o
RaRi87L8rvlx/HiSuhdRNEzUhF7/xDjUrXtpGliL0gqQtisXufW3gwwyK4tLSpFcKf9IqgDIZIq+
X7HLbWx+f/F/X5ijfRmA6I890PdVPuibEB8n17WQtO9CYHGm6ynVr2EYk2yLKnrRC5mIxkgitp3O
TwP1Z6YT/krWQ7kax+/aGPBEfaEi4WlZnpqyQ9cxgC5b8UXs37KDB7Zlc5C/X3DqS/9z8+EsrgqC
nnYRRO5fcjJIGtPRhKN3tPD5qQSpJmIiA4SrGf/ks1TEavLjvLshqfGJximACrkIENcurMrVdgDR
DJfWpFCOHELX4b6Snn5HOMHtqHBSt+58UGlBhYfCn/jv9ZNo7p8YqKNA9Ut+vCy5WSUKmm+asqpH
7WMdpoLAjDSKa9Tedlm6rdKi6Wn06dT4v7sK+iYQ3Ef3hH53p72gbq1xxCQdjAqQiNF0syWxMHSe
dQTk7uj0VDjKemx/Z1ppkz7SZpeh+WQ5cHga5EW42ZH9Pws8LyXcAPM2QCkLwcOtX544GCdPkHEP
WObskFgsv5tcUJEMqR/nlWYlPj/j8S+U/AzcKzSWDsauivRIdsPe2x8lbaJ2BYF7+z3eXazIRcVn
HHMQejT4juLAnf7Wfx1UmP28aW5EGZVIlK5InQlj00TSmLE7RzeH/6etW1E6d2Dbsgw+LYZac5lA
WSJoAD48g7qcQau0wT3jhWtZo9xrRenD4wIjyb37cc9+BsxD1JN/43knyrKWbATQOVi0uD3bl7XK
UebPPcuIRazpsUVD5ESWFlFwDJ1adlP79nXYvkv2tIeQtjSLdlpvgU1Ts1nnNBm2SqCGrye+WVZJ
vfELdS1EVRjb7avdfQ/yWx44DK1xb6WFtD25EjQzAQIY6B5+j08DoKmTihGe8RGDwjoQmHyh7R5r
ONb0mpV9QBTji2mu8sJ7zJcHRRKb7QC9qXQwIyOmMpNptZ/SMH0si7mWbQ5RDdxnIfK63dAdeLEs
f5aI45maqnH1wx3movcY9WG0XT3RtHslix+Ok7dADRSCz89RY71KAEfzpuph3ogpPpxhErRblROn
CY+qTXUp0YcHWDHaIul1levcqcdDr3np/TbU4avgZHqkQb72ZcYwc1DBKT8iziPMA2fYg6hH3n/A
ki6VvneNCLhZDnahlg3qK1qNA2PzHfbqhUAP1IYgQul11riEy/IK6kXZdWOKDslUOeIvN6h2gW6n
3K+e+5PcmrRAUUn1kPGGGioakfaKUULuxiqCe9bvaPQWiQ1swiYfw/0egTQadq1qolyVB1jSpq1v
0Te3rW7bAiinF3QKz2A1SJeWGeiG5Ubc/epJ28eWmXDxrOesJIoVLRQqgScA3Dz0tjloVg1laycY
cMBpvjq0vvQDBiY3UZQkCKcvPYdEtxZ6gJfcoTggE1oevMNy3jQGVos2WtmP/8D5oL4XimJWL6CH
50JjuIENwzjY/57pGutUwDR8SMASdpr5cLTHJK+OE8LAQpSzxM8lfaS2tpdwyaYf3t65t7l5Ie0d
6lKyvHdPikwTsTlDEz0ym0QQYTKjeverX8pl0etgf934QRmpaO9nqmgZBziuF0bZvEaqwirtdlM7
Y3kzP7iAUO7NoNqKmdqr4IceQBRi5p5mz5tqBVAEBeIvTwdsUUgWVXV5HvnTpony0qqOhZkJGRK8
SY6ivKU2mhGl8K9e3kuusw6D/4fh1UITMiR0ZPbP4EJdaHnrdEk5plk7OS9olMdZVJQyGU0eUDwx
Hg4bVVeMtkQKIVr/VEH+Q7NtNoYI/y+Czq61v8OanNcYU/eNzFiY2dNAt3xaQ6zfb32auWR5GkC6
FH963ul6ShBSHQzZeoNQo8Kb92ayTTOSHu5RjHKKXhdpPHuURpcoB+7vGemR5U8u9ydno/LH72ZL
xewGoMqKzWvlLq2p5ECAgIKxJgY3iqe0JQLg73mI3SMOlA9Y6mlm0mlH0IYYvp73EkBvful+JQ59
xKQanqVqZ8FXfD6CtN7phE6hNkq6CrD99mHEvdywgvVyGqKlhSITBORXxZl72BubleSKznefo5KG
4JvbmLBDFw4qAZhXC5cQlmbDD+eIOLQAP+76+Jpw6Tzo+K29r5NYOS6M7QRDgrUTdd8nnaqU2xCP
KaH3FuyrY2Q3EkFXkhJzUnIZcjA4EN4y/vl6LAFjnfcHxZdO0jXkyctOHz36nknPxw6hC8CyjrUg
8zFUPvLCssZMBZiMNuzEQCDTdXN1YlTywQ2PBoKgU+aCGHiUAmpVqva+9YTO5Ux/ovKdQR61sT/V
xRu8e/y+3Cg/LGbpE8NWv3V243Dsg7j4E2Bq6uca2f8hEcRtsyHNcZlEvYJY+190wA4UIHhP/zRW
pLucKpA5Y2t0k1+oS3fT6vCjbB8wCm3SZwirLsSWvkVN+2qE0/7vvQch5HtEdGaseSINUPpzxHxZ
tTX+pHdeFdudxwvh4LLWR8/pVb//+UYeQAYngNS4ufyGcR/PARJC9u1+u00iS5K6cs/i23cYDUjN
xaJxME0Rt7G5LVt7zBVON/DRz0fqGagWlDqcw48wUHvLJbnyqNwbzDkwh2qyfht4QK7IZgCI+cz3
PwS2TyH7Y8F19/1GgWfp3cCQM49RJ6Rnk19k03zzt0ZZ4u6Qck8ofyFl4FZyZBoBrmBnOLG40jD7
VCXExBaQ5D76F8M1GG92xBylvycrUPkGXEeW4U7pREX3N+nMGsYzTqDOqEf+dhLLJbebYtPARqCj
c3YFwIOU6zFBlp1f0cF/cARu/O//tvJ+5gtzTVOdlDaPaLOBjuHCUWYqDMyGBi7F3BaHiYtImT+T
FnV8LvB6CVHkxl8maBAjyIhSs20a3Nu2/rRcYsCZpWXTXAMsDcFqumRcENSb2SsOHKt6YvcalEdf
efgwSFM7UgRGX49odwBmBCLfoS8JrB0g//43bVdqBQ+HIlvKFi5j4Gg459KiMI9iPSUy0AbUfwwx
riIIfog2wp+lmsdKYO+PpTYqF2uAlHpHkbG6ZT8tss0KFvcZNkZ7vQmZfedQo/jpr0Bmy/P8+7k9
OkY5Ycqnf6O0yrmpngwZaeOvIwgW9kmCW9m6xsBc7P+NTmTRuYvlaxmB3a56A7gmFAjUs5E6oC9F
lKZSl7BWkJ+nUxuKE2ohT2VvSPDW9fWQM6Uo7fYnuJ38Oee9tgKIrByin1V0ZeNS8GIXC83Dz1FD
llc3oFM/B64OcjO45r3UpGPKqnYrZGdr+TuflQX8FWAGOyga1wmVKiEhsYqyB00xO7afoGz6xaXG
MSEgoUnhpdLiiUqRvQSlc4Qehw1cWRQ2pc5jW66udP9YqB8Cvo5UPq4zvGX63ymB39w7AATbLV4l
1akBeFaTfdVB06hgRlP/eH12WkYA2/75qATXl0PsP4JedMdVWRi4Bv0OGL24xujSFMcmgMiETq8e
IX8RcLhHQ62CCr/fBKpCKj3Vxp7IccTv3HdgePs2U7Gy0oYkOB8Jctr0avHKTsvAAOyrsan0H4uq
n7OsaOI1RuYD4HjdPqBUdmAloXkSM3bzJT6EFaX63+CKjUaxBfB68GmcrP8YYu13fJb4uwTbxjNJ
Ob4QohJhgF/5PYzJhTGoqdpwSXs6eHhV9qHRo6PRYx+X+htZ3WbiSdB+8tSLojeZ1yDe6RBdIg65
i6257tAKo8gqtkDVgoeqepqjWVcDFr6i3Gdtf9uWO6e5SCqQOyK02MNgESPBWAiIsSf8w8M75jzN
tSfc9F77f5Brl1gxhby+1eiTfrWWU69N7O55grPB5XlxwvugtBVELW6X5UurVKj2M5l8/V97ZKKK
ReQlOMSUQtkquu62C88zx9x0uFW9nhqUy/a6ecXJRDc1DhfAR7Wc/onGVNqQF7Jq9LHaPCoI4Zsv
9YpdbjjnSMjzggsSKf8S63SdWVlux/i6fbGATSkZm90pXQHPPI+zYVwQ4aYVrU++aU3S1FhgiTdP
SPtX5l0xpZtdtU5iKQ2E6z3ovg1HZgcRfl6qOXAJVWxkw1pobznaUhq5zGPgBPSdKrzoBY8vST6K
Lbf1sWiQ13ixfKA00xGdHiLAeu/7nOTOcSxaL0hteub2jeWBfFcjhL/wzEeG+WLQSexO5VisDgeg
f3aVVYFtBThPTSW9EhGK8MeQI2BSbZnWAgqXvAPvOHn8Hp8TeNilvBmNYiUd4ybK69nsJ/k1ryUP
ld/BQrRbPlbqKw8ec/rp5M15U8qEeEmWjiHNNU8CoWFfW7iFWjBYKVttmGT6tYkp+ZaYLubw0eJA
g2kqryS1usUxo6puL/h2k6sOippapr8QNClFMDkTkbSzIY7jUjpsehxrxmqk1DwDj8fUOESTzIOn
mazzlhWGZnzd+xR34ZOZNq3nSxTqTaO4kJLx7e0SNVY5widwG5wdLvjPs0r5/GsyuGspv+mAuzXn
/Nmr6eadEVwiHzlCradzKVUc9jQR7OZkCEQqatWKHO4fTkr3uWhkkUUEw9UETUSg7ohric/BP6l1
L7Ib6oywbHK8r+IxqX9g1RCxlP3NViW6ai6PFAQExU6THvRdUf1ogqn3ZV7mCb3r6OXh/GrIX2fL
rPVIKDlGWECmSBFbvrdYUgtAxxJcsodkFOxaYZ0+DJKwQiKUnCdBbSlXaHy/NKjX+PvwrKp5fe0O
69HjXKgQqw0JtQ745vJA4BuOMmBSIMOdU4A/ZeEwOcadf0u3WApzXk5aqb7fhRn1MzJGPdG01Pt3
vf7+UotXVdI6619Jl1UpHZizBrbsdMdWpdF5jeAC1eRLVMuhZeayhbgMc6yCDzyVErUFhnNW74JU
59Y/RXtcaeJab+3yCxaqxMQPjP4tDGL5VPX1FUV/PoY+8etNvmgmrzqUbACj5oUt1vF5H+IyvH+Q
fpQsV+SpAqEh6xIkgK7KT3KSm1gS9PQ5yXAd/jxh7i7se3ZG1ocI3o1Ckp6pXwsCD7OKQbiOJt5G
ob0eItWsinItbGxWzw5tnoEywjnj3nmH3kzKuh3LCsJnmEhdevAkgX7MNmlj5ipXnM6dJMI/Dj7P
ORbZbBbBm1vpurSCdtu2kWstCYpBikDtCSW0hd2HN1rxS70CDaTCGxExH4RfJ06g6N5enYrTeWa4
kx/FaLye033DJsQ87wjn0UjyTGBLM1O4lIDY181FcpMK/nrmlT/OYPuXc+Qz7Sreca5oWunBdQCg
bQsHtCeAYWvJuV9L08gRA+xGwn0IHQdgmawRV1U/3AVeJSq+xFZhIeWbTd/eFcEynPK+F+l4+/58
HEVL47oPHgmDJPtqyJJ5knu8gSgKmX7ma3oIMaw3YtShiy8qJ8Rpe0hEyE9FwYsxi5Uw/TAQ2PIX
VeTcGTQkEA8s1a6rfda8DLPLmub+QfOptTFEH7Oh5JAUBKWkqiZR5oX64flC+eKL/StCanK8HDHj
HeZOBO16MWLhALQCYDP8lECj/VcoMTXcMtMyUAiHsr/vfg9IZdbUEwl+Kj1RTyqiOWmx2jnfdx61
hTpHBfFCxkvIehwe+RcRbeiHsQ1odmxA5RIFxhwvJLoPNWS6uiLP84gbfzZw00GupOo7nKdwJk7z
iGUtJKAjrAoL7cJfoZ9oSt2oP1gSrCUFdyAQtg2uRnGICC1RT4a1wtjihJJzRr/FuoTS8W72+l44
lRL0AwMl75qPyx7uyU7rHCQK1auudgNJX7059RI+FwNx+Qc4w41QsePIKSo6yHI4Z3Z/kkEoarr7
hX65dC8xbWbuniO12RoBpztbS3/buKvRr7ngFYjf+nKh2fnhhhWHO9tHJcZTPwE8QEDVWaJqmrmr
VKjwhbcskdM53fk4dF8Ejmdr7wN9KBKPfyinz2gG2+/KUe8qhO7U8HAaHIyQrrtRrvpdsWEh/P5Z
jkfMNLbtSwrlMykonnysUQOXdyKM3pFAo5pK0bp+94RiufvxhLg6hpNHb7bYfpPbaQmFxIksiAWf
8wHEm/jIH95RiqqJwrmAmSMhcROk/Utsnrnq9EtCkUQ8k2CGhxkVxTr+iLlKfyNVltBUTaBX9Uu8
7NxCRazcXgrGL2bTiZulVvoQl/Y1hPidQPn/ERvsRCL8Qoj0xn+8B3z5AAHs90RUC257Y2fgVqAl
t0wZPBIMpa1G8vpNX+wbMRyd0OToMEnEyTWXfRIqjaC+m4gHQsVB9zEuaRpkXKhtXwPdhDIu9GHS
9qDxIvuRpMmhz2M49zqfVk1EZPwos5S2KZLaFiwUwdfreXyUxhzd0zFMQsWGoUC6+LbD6doxtbie
usST9hnb0pZGEXDNJxElxiwflyp8UM4FiqGndfImT+dpDyVGYeOniFuYCHipIgYZWcvYP7Z9uaG3
mXX8uHCotOOdOOVznpWxJp+1HdwksjgHr/7lytAzz3n43TF6CBjJWisbzNvyc5qzmvcQEUWb+D0O
bo6BQ6tDA67LqyV62xFiqLhpifOjw8KgUbISaNHItaSBK17jrK5B0Zm9syN2ofBex6wjFbPKcokH
4kKMx+0bLpUsLH0ZSfW73wjjSiLyohuLpdWXZdPhiXTrg2qstmWfNvrBOzyXN7YucgEuhf7INCvO
fBGXi/piRugAoxM/ifbB6MMdoaVk//Q+SrKScm0nnyprTfoGo1PPE85CLk8mE6BSpC0NpsLiDK8J
uc0cTZVWSHRqBG0EV+uwz4dPIJEnn+J8ds+BhPT3LLWbUlCy1KmvzL7Ij7DwUzRnaZecl0cJg2yo
qOmbICokEIpzJGzHm7miKVdrvO6ln4a0y1ZcQW3dM5Z+okFmo53BySdLJlV4hoCyWGErGvKL7vlv
JI6oRfvYt6I7lCeRQQfe/3aQ4qZZHLjUZY32KnXDgJa20czXjZtnZkZih8hSZMg/wJrxT0DFtxuu
Pj2TgPnCOUOsnW1NDZ5xFpYaElgZphm9N//zw15D/sItosN8c290WP1VFqD75ckPR0w0S/YolI8A
kqRb7FjW2RiONZTzexlUJWvenzONf1WYqgAjbgJ1kUy8KchRUZtgPnHFWyhgDyondza+6OZLcqfA
brNyf1dxrM6zpaGM2/K6wh7R7zTiDw5V4ZzChfdmX9Z0qaySNuT4Ewdr+xFwdsl/PEDRg/707YqH
oTFzLDfQOYld11qHxQmmbgNHCw4DCGfzMAMZZa/lXlHQl+xX517Rn4bqeZnvdwkHBTkzjxKvQBpO
XS8eN5tdlrNCpUiURE9T6pMiR6N758Iy1cFPRJGZ63qFLp0mX4p9jmDQ0HqYuiPdlyUUNUWG7T3U
Ib9spkjkNshSJ5ZmO1FGCr1attf+UuG2DwXgs4jsMFjHqSli7zM958kmSYuZqvgHdYxVu7X/R4uF
/XLbJuyGbEWvuVDktGJmSuXnrbMtOR3P2UQUpVjUb1OejT0tLQzJkteVlBsFxImHoqtn9HUiByGO
xw5u1Uq0UnTG/MwRUBW/j+OiWfhUB+IOcyku5h/+7sdniYDNPkWDHKISpM6u6ARRsoU8PxR9jmvs
Pj0HL7VG8NTi0IYXaBkqjOzaLq6kpZihm8VAZSTxiNxI9dfT9yfBN0GCGxkTOIqd3XTOxUf7mqb+
jsbbVhDZcaiUDJbBgwJwHUBS/vos8j0j5kmgKg2z1b9gFRHX80gZ2Hg4xAdNGYbNiHf+QMikuIva
zEq4BT+KJ8Zr0KZWAOUU13YwXc8TDdqvM40m6+X+iJcP7lDoQz+IrnJTz/V6SmGaY1BWor64cr28
VBxNY1P5QgDg5ThazjnstKwnCD1WecmXhNixXxQ7j6aZu2h+XCVK9bRODu/dhYtrkInVsEIuNtW3
l3GQF4eZZi89Paajg35SjfnvptvG6AkWnaOoa4lcboLBTYwPm7LH0F9tD46EKCC51mqpSXfgNwzu
4SqLofAgFfSJvYqIsMbI9br7isvHf8pebC9U9HMWPKybf3yt2FS/smW504MwRm/HqNChnRcXciU8
15fVnLemI1etIgX7DBo2M22tXdxJSnib/RmLNKhu+TlgDwMtRoe14HCaWS7YY2sl1yHV7/DobRAa
+MDkuv9z87FzqoxpYtVe0A5xaElSjl7y4XomVIn5tq0YZYQifOW1knD/cPs3WYyF7EtWI19N+XY4
QGH1GkhH6WpKs44cSC34GnUFKSqTjtw5Zdz48C+rbsAZxyMNVu0+K8GhrGyi3IuuuF+IK9F6IFtD
jz/w+ZcYS4VCT7QI/Fx+fu5FmgEIO4iTE7FlHBMLWwvEjhW1wbMv9CfLEsFPANRScBhWOu0h8tSf
TgcsWZr4HxFennL5bKch/l869UOrzE+bemG13zavQ02AFSUV7A/8gDFdZEZ36BeShaVUjCG92Egq
8caFy0yh7niUpZPx+LwhH9QmByIYTI0AyTWQnvBa/DiP2fBCgFCgUGRbcCl8wg1BB7/zwL3gCMi1
x5Dqo/D/cBvEyrFX1VXWp1D+gnZ+7+aV1OaNE79LE+s2jmdtMocuJU1Xy9rtH/uDsOpo7ii+KWhV
SZXYxGXjYuimdWetirKztHnLWIVQyhACODrCqEdHzxPYo7L/JuOD3D8hCFFfwEv9D9Li1ie7SXMP
9c4c86VSjCwwfYNkp6sqyiKThM6pStLspqmue74XSy8lrgs3uInh7vtJyMi21ZZF5bZI7E1+bWaT
ZowzPRIaA3EH43KUebyMPUIZenmZNY2r/ghxYF2muPp5dEN1RfMTuiRi+/gWkBH2I+Zt5H9yADCV
VFLIvLXQF6lRBeffOLGHG7rKh2pdILnfjCuoaeVZQbqIW6MbukCE/OpP4jcojOHn0IS93xBZogUJ
HHR3w+lVjHNrdz/S7HUAb9FEabAqJIINmL2ggpw15NAsRKlWu3jRMN/MCeC4qkYlm3EJQgu5lYz5
svClvYGF7zKcQ7k3GQEPZ28q/CivrXVrUpqHgdYeXrmfRfOdVNgP1tbuivtGxhE5Cu4+FIlUsmuj
0oxTlA/yvykMg8OenPS8s+Pt3dm+S2JrLluWaX/XNx2kfQOh2l+lDmIfY0moEhB5xJa99VAAVOY+
JUPrljzDEpWMBVfaR5rJuwpDE5HMsIWD1kiG69Xs1V38JKNBjS8GINa937kt6C3nIuaVfXTA6zHE
g7HpCgGnR5LWW6Y/qJW2Xf/8MglaZBXStb7HR39bMhv8ObDNouOhUq0AnmwvAPSxrmzsAAdZyP4f
hZYGqOWGHz65dORUqK/4fcCbX0eVfVtRHe/6zNQ9+dsghTdtxmRQZjAxITutDm9faxzjHmHvA/6u
FRe5YUkSRz86MXTT/Rn+ZrSpdp3rYHl7hoUomNDt5/x3wdHFwf1qk8livpx3oOMieBDkkGTe1Gop
lpCoTMFrp9TxxNdSyy11FYWZx13u6jC0IrK8mRyHJaaLat9h1lS2Hy2xuWm5eB3dj08n31mkvZUc
IHi51AsIBRxFfutiJ1MxYbOUwV59q6BbYMoj3uHEEiPMbawchJlt4/bTyCVPpa7c79LoUo1AQ7oa
tyTlUBpMDm62PXJMkaEuAq6RfqRulKTLReHwnqYm60Ilba5WuLDONE7s/j+ppgqjk525YYjxb0QK
GBgjCH+pBGVUysShrgaWu9Ph0OLPSaSWSecDGNqgNBTZHfklJH7lHzMDnAcFCPDEBC5it5X7UPkF
oWROaOOeDxgXI/EHSKN9vlLTAQ0BzztdJcZgFbnQLY7QwGLi6wgSmyHrV9fCBxwY+Q0yYzA4xE21
3cw+mjQkbm9zBhAJlgHqKH91qKXOPV1pSqLJ4WBW0gg6+/eokxQlhJktNBmInKWP9BTFlw6IIuXE
i0y/n33oVOukxHLxxTJMZPn0iAUXZzYb98IDX4CjXAbscOutIqas4qvCU/2eKxLJV/fK3XtcdJRR
ddB1PXbQ8rhHdyXBmYDcNgTqauBT5BIeITyH0bhMGB/kiZ73yH+/r847FOX5t4X05ia1mW270KrF
tNo3qzSfvhVt5UIte2udRGMBDnYW0ti3KaGpRnorjGZrEWd9TJnetvmFTTMVNOxeY4JepivKeyst
zX7uNrN5FWU+iAFMIzQS8zV/rTZKUjknCCcPS98fM6jAhpbdf3twMBHe+uaryueX2e7ajCao3HwD
gr/4IcHcqUArbvFu3YSjZf2p1TWsJCxlFk6Um3NbMARZxyqtNXBKeKE8OiIwo9fG0Q9xybQqo9Ox
0reWqNHhmbhF27yy4JKMPZkcupoFrfls/IrRhvd0LSXr1n7QzBnGZ7FAaCkpXklO6+S0WvuIHoRK
J5Lia+mC6jvhATMZ3sePoVSp9pYA7L770l8gxVfgLoSFftBth4/TMGADIupylYvDR7DBHpG9fWw3
FKuz2mIhcdT/hPfu72LeKyUGrmd8GENYRgtdbfUU5++404jaOI2b9SYBEwdrjHAjjQ4Rg7guMrRL
GqdEIPV+j8aHVNbNceyG2gPnV3fF9AzULvXAM1KvwUrH7uJSI+4JqIP9oNHrGTrMAh+i6vsM9NFW
8phHIw3ar/FYAr3F0xBDNdOwb+fpe8iR8syvDjz94cp3QhKSmU4lLCRuwknkxLqxUa/SqOxTFtzb
YE8skrJoRFM9FM/WjJEIVeKwXEUvj8DAWMYRr+VlJbXbWOLQW9fz4fjCzLg2euhsNaF71kdzLzZe
JF+LALR3rUtTs+XOOl/JJE+9WeHCMcM2U8o0kLkv8W9rbajUo6MQ/Gc4lryBBz2T6d8eifx+Q2fd
BdstxyaVg6cqSaB7OWJDxeNafj2lLaJdXni8k6L5KvGPUqnjujOUye+YCQ7S6kfGqcaovrB+Jgke
oovgryvd4IS8cyamI8kbNUT2uBRyu5Vduf9+5qLfkZrVAapWSLWyzPiUnPzUjpx5gnS/ucJYC36W
0XO0FxjZXy2X1Suh6AcXoXQaKGwqktKxNYKalzGY3OGSK1GMmc5UmQkRvz4WxfXeD7DIcYC8kHZQ
qR1QNJ4uJruSRBfNWNgmLh5j6QsBffMLl2ax3SeogkAubjhgZNCtnRHl8YZ2uZRPL39bEzEsovwo
CYzqCGwzZFt1UmfvmbFUdcZeOjx/g0/lLQBDGVN+w9Ci1RivVP3ZP/E0LbJiIfsJLFXS0xUSvitu
uoxn2wQnSy6mT0Jc2ibEYWG99cNK/zl0E8sN8yi86BbLofaMctyKtbzwEF+rr4VJtu+75xj0Y+qc
DWqRoRN4bFMjjoh2gcF5qFVWw1/iGFjDjzNnEw/8BFtx5oiZC6YFnFQECpmntjQ13auqWm+SLMz9
oL2DU9KxZWQocNEL3hu0+4Wk8EyYfgxiMPVxPXajGvnFPSDIYKVt563Q9sKapMHC0lhXaLcaSIgq
mw696F+yUsbKhfkZH8Pj2hl6DrKKqNGLyYO03fZBRStGF6sYUT03hHgV6Bs2Tpg+j3dPPl45mmUE
eie/J40TB7+2FyF/VZvrrTpzyeLnwtTNMlb3S2WyotiVN7o+HZUc9odOpt1LLFzkmhEbHUkOBRCO
+urzovp/VZKU/u24VkbU12BLWK3onK5TT3OpJ+VL9MPxPkoE3WfhHOH6m0gMJjzTiVaTj/4Dhu0j
m99xuxt02bV1xIWqp2sS7hZwFQgDF1Dku7cyoLLmlqFJECwte/7ADDTGOyXz04W7KiZ+Jj/V+si2
I7CIzyyMAKi1H+A13RmrMFtVVDfA9OxuDJZDKDgqIIiSQw26sE9EZtdYSc7nPAX2MIBdFQe56rSa
/Lmg7hx0J4OfqaiKKr8T3ijIeZRe4stUgS+9c6ZRt7AUzIW3ODPR9yAJ9xXzv50zZFLv9cMyTeHh
vyFdcTfhFecgy6UCVNW2xCw7DU7jaaK+x2+UPPajbvQtFBkZKdtaDyo2TcpcWARjz5Qd/xchrh6/
EuXsuitYeURuuW0ummXjBYDZxjQ/Dq93WNixGUMWRxPEx8DJQ5bo3yr2WC0GwBbbc9FAwO3xNDYt
aHaM4RCIe2WE+iKj9UZDgT/RQMftmaS0KXfaR+Xa/O9a7CY/UC8Htwi4pAA1kKEvlJDZ7IlVvnOZ
F7LeoH+sLyEdZu0F7WgFdtwAW5I9rJnbZRiMt6KQezLIkEeNd9Dt++mtcJwVpidGV1wkfQp6sVT3
cc5evHFz1Cap+5HjoBmX2dtW/svGyux4SEld5HEwc4L25w+kSXy/FgpnEHq4rQJD73W1LT5wXcsQ
01Yg1Pl82qZ3EvRsgFZcFlLl7bxc9VrlyhT15HZpUDh2a/07Qk9878jv3s74Mh/52ld7M5nQHNfr
R3JH1YYtGI6KxO2ngKgTUiEzvseNJ6QU3EyjeIiSY5TS90vPVH/yIGvYFAqjhVSCilwYGAtAFWWR
zL284yCbBFchC2hVmE3lwtum/RyqEjrDYJPCUi4xa5LY2b+Eddket7QDGXPtaFb3Wr01BauTF3dj
QM7baoLBbflWuzhiv4f3BcGprMg7VupVtZ2ShuGv3RahObSgQt3/1PYi8tgdpOa88NmkVFExF1o2
a+kWEIq9QpK/kJvRxtAkYG4uBSLV52iIQj9tw9EgAwJBZ4DbUt0MRhu3CD7+CuIOHZ6smFjqNqpV
3e3Pc0Izl+/iHfNRSahVeU+aBaPqXFAHCUk+By0E7A7rxkg33J4v4Wb1nIhGdPQ9y2kyBtTABwib
pL6yRQi533onHPlcXusD3Wqqtn1zJIZl1wJgbqoS/hIzpUDaX+lg/do2aonchpRlebB/ONUq5nn/
oUlv4jqT8n52kS89r3kvJgZEce3r3TB7Oigb5HQOshXn6CVGCn+xkTZ5vOVL0/li57MoykO1KVDA
arFQpDnAjhENfxXKAGbmdMGf/T+PY38HRO6qKESNBjr/V4/r+LV3QDGR4MR8ptNLte/moN2ctdBk
SCKiv0whYR5GIgtl7Wfeva2CjWtVQ1qgvqYu+HwsJo1NL9vClrQCUXZVEZuFIlioQhMhZtuxMnbp
7dbv8m9Y8HfShCy5d4P51i0/1ffUCWJ/OfXnlsMWxf1JXjLkN9wEEshVJRzwUOP7fx5VBRGnDSxa
Rk5ZJTHCvmR9cf1wrs2TspxAxSnLdG/58Y4ALjQ5VKDMYgwxW5gVrADeVNEC144k9HtDs/iEeJNp
IzMiQGqwQfdKYtXUinv0hohp3lFqrjwYvqVKwzkXPXv+TW3GOKS2DpWXerj2ANj34DbTQh64CCi0
dNtW+gy9/0eHEL4Et9xdOoPJxzJAA+WFibMTL0+sbDdpNLcDKZga9zW6TqfasBpFSx/sRukz6szZ
+lHThPYPNNgwuYorhpHt9vJkSGctpLs3EWjxMte+nMPYSdCQ3FarhDQo6fTtE7flIrNxc+JYXWa0
sUxpci2Up7/L232SZjpHmD921CXFxZBBayW4sGEIENJdM/OTy7Ab4hDnJR4azAc5MN5muzDK5dRg
m2Z58y7DvvHg55rq+6ombUP1nsXLKZBsxXwE/Jg1XTVT6QZ4vWICcLPRzUud4tTyH8n/TMq5FICx
bYvwT6VT//7Q1w/pwD56/tssVMxiNVA5F86AEoEOQpwfH1jUQy6TLtnzijN3deGaqzq9PgvERBBa
4e2I/FVlwws5HkHcXOvPT9E3P2jfQxSpyyDN5bOMnO84Jw/FSItN0TI6bznFUJ+K7MCtPlRNXbdr
zzxP+rXpMnTrFCajR3qRarA6YQzV9xpJNQYfAq7wOS2WqAack3z8rynJ/QwRcjbk59wXGg4qXpEU
lA7dnTzgurhxVe0QaqZdA7PreyXsEdKodVzxk2aV2fkPmeXeBBR0bk0LkeG9FxzaLijHfpiLo4R8
Z7yaTzA1pEduQEajACKFEkjHHSmHHRj3ephgqWShsJqusUC9EknuQkeTiBlxprOmecMbdrPDOzYS
vBLnCRsJx6fX+3nrSkeNqGReaZEa/eGn+OQr1sbLEQDEQVCWM/6Wm7OpI0MZ/+bvzBXQ96pKS74A
7wkrkULqKM6xGCqU+asbGNSMoeLTY3P014i1OtIYRjr7BsARK4o8VH/S9kA3EQQe5I9vF16LLcVh
Cet0pYPmE/wbXXwXId5nFesvG1gel0wjPSnAruK8UiLrtWeUStCq/CHcaZ4bs1cB5OmSDC6FnE/c
lCXMfhSpkPNN3WkKU7iPAgd+yc4kN6zS//HLb6cXv7vIx/ffUwiS1xVsnMVZFvvhOTKd+Qov2tHu
LLLziewDMvpR0sISA88ZAlx7vICDMFIE6qqqzmRVqd6nskz2cZsa1g3QME5c6mNYREuzJS1PHRJY
z87KNyVGYO65DDrmMXbaoG2xVGDdT/YJ7IvCOyo2TC7yKerIJAJB9UGfrDSW3IFYgLNZ+hwiqnfG
6xNnI1Yut/YL5kusVwi4Me7euAMsWTRrsaraYYhxXosgKHn636KxUfB59IOBcaJo0WgcL9lKrIkx
Sy6sTX0m8D3Gv0iAAz5hCDB0WNUCf6yOn1SqFJ4gF8oDEMwLqYgBjW64meKbWJ/ABLUl2oemslJE
1T2pEyHMty5iS+pR1BMLj5lO9KA+L/BfpqrNC3cqtBhChy9FrPYLhb/TFdjWPtUq7r1U1bL4+AfI
QcBJ7FFMTwv/6v2pRivBCxqUnFj0PNaGKkSpEmlEL52oMOAFf0nQz+xxJWn/LW0bB8gbX5rIrHFk
crR5Pw1u3hWNT/p4CQ/1cftXNjCYn6/iG/hbCPNLDm6LvEwVRo0/QHBzg4PgKXTtGIIhsVe96GA0
KMEqV2/+gpbiLoIyCtb2LOSzftWIClmXKnX94NPSQPBcRG10+AelrC/angjeeu47yypy9ZHcx1a/
k5X97cniukqS8aZUX3V00mypiXqojOZOqBFgD6VFQ6lEMGb+IQ37ht2GRilb9yThcoMVhLEcZ0qg
VYDRBkIkH3Sq/O9ZeUWo89UzEfVA3bduY0CrnUHvnJRu2bBsQSu5DvUO4qXL25F9NmYjHdiH6Fzu
NIxW2JPPwnb5nhW0fkXh6GHvffmam+WNy84NCLpJj/U0sY45IUTSLpoYZndddYLg8PdOrvjE09Yr
/lVjRH3smsmALwA8x1uXk9KPRJmz6s7gYjbvVOc7MXyMvBU7rOSd/8H09SB5aNE/rhcwtyQMzT8S
r02SrMq9s+ow9Xa1AAurFucEKcuAA0GMtvzwtbt9Luq7ndmdEyTYpKclwunMSSpbXTCoP1u7280w
xKNoHVFpvqdxYAE7fhm7blnorRCULrpbcyPpNGjAAF/RipxTJX+drmLVOx6UGYt5GfdQFtrATonf
nmNmXUs1yTASXu/AJshP2rtDzDKPl/nkkN+MoJKgzT0gYbR2poEFOaiM2NAHwQtYJ2hRPMXm5Hrl
Nt1VsLSxUU4csLKc5/ms43+v/gLj5GvREz/PN/BfCUNbs+aRQD4566fksdaxjELme3cw/HGd3SmY
hSJO+n/Rmm2WC0axY6J7gsvTeH4nKN3VnXe3xZIaiaVW8rBOp3AnoPfhGgEwtihsxS2jTikwQVTx
xsDl48qexHfYYu6PQagN9kEqY8E4ASzGBjF5T9y/qL2m3LJhDzQ3THMbvakRdKvOy90Sq2T0onFu
rlYr9CjGUEzqwrZaOC+sGshaQlL2t9lrRhtDRs2ICf2fx0rN34dKrLaz8YNmazT41R7pSRHIB2h/
9p2IJFHzHb7KjlnhaNthU6VJvmNyK6ceyWiDm8Sqfgf+6X4kEwn+NxzSthR3HGpsTGGtPLvQz98v
F3vLX/Ndbd+OHhBL1ALX3nRZTNcl383mDfL92kJBT3CFnZ9Ie2nKCMjMPEJlrpYPyzzOp0T6HX1y
ExuNt0ExMaBFzGx00L64Bt7uLwYWeR3Y3Ml9atedZqlOOuzkIC8Pw9tDPPolZw3uAGos+VvbDGXL
kk2VBxQvRvLR5G4j8ZFLggmxT4gYrV6V+EOW0sX8WTIIZyoXJ+p/lPpVITFiTeSssE+ZQMHkepqA
HRXE3sq2wQrpkvdm2MXuBRZrfxIAGj8y34ALvCUt+L7pijxuA+fmg16lzSRPDLvq79gFR78rsvnV
DBdL5IKNIY2MOAuQdu4GAGzKSNyUSgWi3hXE/ZXOhyMN1x+TNa7+okHuR0IE6t/kt/P466hYGACb
kQJoKjIevCt8KaVDSkLucQwk/lMWaBw+8mCCm4pmDZpku2HQSfVOPiIQ41UBcZ2PnQfC0LT/S7hd
H2IUtv0jJTMNhdcSP8YPQilyK4w7ZoSPcMYS4Iku0iFpWCZML6o92bMyZlofieFcMOXJcL77XPPW
lG1mD9Kvb9nWrGipxRg0BmsON43LFaRk7F+Fs6NNvqpdDpTr8J6gRFUNZ2vxRUtNjJyAGpxWm/ff
+jan8YlapR+oE90E8NNExoYyTyh2pvs+5EPhm8zvM7n3edNMSjAd4iLpztwdm0FPns57PdTd595b
MX0j1BBJIbOZWIpBYHv5fMkEG0ggPPSut1/3i5b1yV7h1POkaQPaHngjEvSqrpRcPUNImG/NxVLR
oRCx1HEZHrWHgX5JznbbIdmGNABb4ysfPFph9qwl7Ky20fMMtCAQK2Oj6/pzop20IVSQ2aMDNTEy
xNPihVXI4Fot42ja0d2bf0WQGFz66b9UDCVody3SJd9s4rmJRUIHxONXtkEiAxYnU7pCUsUXo5U6
q6BfHe8VeS70rPtXA9CmqLPx/0ql8yiEz8KdGAwcjoGvjZilI+ifMmPch/lUNnNRGuNX4DSX1wpN
HMPcbcpBEExsE4TlKkaCP+5B716EepjchgWdIRd4n/05JWJJGXZHD8bQApACK+0xuXr1L7eP/JBc
a3OPTYmxce+/rGl4brFBqZqfj5mKdka/+RWPbGm9pM0GZ813XAFQLfoJQEnWIN86wCumtQBKi6bQ
IirMnY3QEPtJjiw2x0l4+HsTJXoAXVS96XSh/omHODqPLpFUKNvasVKqtZtQu1RnZW58MaZcUuDB
JD3AR0/G7KY58VINYkhsxqN8urWQPEuBbnTFdwyIQNNa38rIZLuhtb3rKloXNUozTjzZaYHgbwAV
e6+KhHo9LGp7xrk4HAXednzGrP/lIp2onlTdDN+7zOIZyl1PdKoCN1D+CmE+ByoGL78Wf6XMLocZ
fRZZOSWjnJVN0q3DSosVZv3kSbdtKf5LK1YMxaJiQA4068FoDTljbL7x3QiLqntqT+8kJsyFEusp
qLr+FdobPkoRy0KPKmRywO+WjQuNdj9YaasXyrO4R3dhWvyvNsO9DK0vpZdtOVZzh6XKpueXeSOw
PAo8cs0VDtwKbLZeXRkZ8kvE7Dwgl298aGH3MMbDNAgx6mPiqhqoboP4qhaNNM3PJKHxhu1/yZOj
Ne8iiofw/t/DRVCfB1zvYR/sWFmBPkqWlJXAYDGYpjFc6pZo9v5Nj84mXfN/fyBANKmkrg2pqgtt
A80AWz9IwglP74UWysHDgmxK2rFL2J2lYo+sl0vJTqnxvO+GNTSWLZ1t9AApgzzXbUZAxhnAY68k
CUhg3atjTRKmn3/4Yu5A0QShCVfX/V9tyr/ZNlby2rhu6Uay9q4tfFzwXOWvt2YDLtaCOBKJMH3Y
YosAMNm0M77Ahzb4TYySG4NT3pBGgJzH6JOkyDcdPOAkXXKrq+ygiXdyhXylzz+jCg2dNaBgv9tR
gUQWpuKv8LE0gP/08kXoR7Ao7UxSx6/Fy6L8S7e7J9a6+x1RX84qA0VcdjQSPSx4C/enKP7zlX3T
eJATet2qs6T8cjRiFCjYUpw5WnqqVY0yqUG7zDQYP4rL+pbBm9KcVWWHBvtSHdFyAPsBOQkkOdkx
WbPCug+Il0UM+AK/R2L9I7qXZUDN1d9mJhnspVtiPq5ZgIsrifjkF7bZbiKLZYbXECNR/t+clsDI
cXYSgwDqIJFCBMgop4Sxw1KEK6kSMiCjkpfcPumfR2XGlIBSK3RhY+a0EWD8mpoIbhbyQULTtNyg
pwCkTRltQnpRwNBCKCaqDKgDHEogua/8QZzKRkzBYcEOdW9ZH2PCCMMI1aovH7/HrtD01By/63Yj
VHVB2B0aEFixcspoZSBAZINnsWWR0/8i7wipO1PP9p1aKFe5ZIqSmCdxAEP1GVRlRexA8eIOjKUG
WTg9pVQpFqURK+OHtdOkVIivhw1WQhj8kMsD+l+aERC0B91eD5W+3xpJRalAfx2uGXL9JfZcHZCc
rIjFJDa5oZFXsmH013WttlJmtpu3ddC/RPqdqCzkeBE2elNEtUBTxlvcZ62xrHQB3a2m0QNgdpCY
ROj20GjAVb7fc4qX0a34qwpQndNgXTCb/krgqwy48AY3cZ8rk7g0/zh7QqRlOwy3hbBRiL0kHTIM
7cN+FbQRnfKTlmHUNBOUE3gPX1GlKrTSAE6E91VcWRdDd9UwjU4Yv+LF3lQswJaQg0v7uic0chnY
VpYyiJUZYBrlYY0U+GPjIt0BZpBMVs9Vx+6z8x8EJ6qxeC2txn4f1fDYJM0YRGgEoplNfYDWH5Hh
jKGX71g/9LA4wHDjXfeTFeQ3JI/dgY2MXk6tfGXw/+hUy3LypCV74cs7ax9Flr5CSyFFUol1gAYJ
CaRfgkqWeNBTHBB653BvQrsdwMJwfqn67mF+k74qpcPBaFOqVphX6Ro3WAGhrcbFouc5jFy93w4x
ddER+Kzm8eDSC/9l8HhGazSqy2dadUAFvpbgR/haSUsc8lnA7R3EMf8exFc0tK2mWBkbFaGLLsrN
rw+L0U+ERueMhDk7tFw9jdfRM45lbvawxa470xQG7D2GHImvCoN55R8do/LuY2D5zhIr++1x16LQ
EldpKlcU9HRV4f00iooll5rddRrLMbE0OtlTbvsbIUG6xuw+5HttSlCgcaCPI3R8Y1DmR3y9tcYs
5K/e4s+FfvWKRtquI7fkNGIrFmClm4SZeEjANPjaFRX2NHxLrwlR+DXT/uC/gv6mgJP/TNhN7SuL
NlW9CO3nPb6Ag6hgzJwWsQpsOB83NgmK2DYXtiR5CzjWWR0j5s+Qg2tPWhSwNf1TWFBCFcW4PoIQ
gLXniKjDbBMUAv9YG3NP3kzotKg1ZqsNwqreFvtGNN9TJsLbRQPSEgROXMo/bzOZ0T8Yr7eyWWHl
75h973ltFKFHBlRjVOjW7NTDAZsSeXZCofbF1Wn/tBvhhnz9GJkZH0rN419dUpVJ7dHzSpP19zB9
niqnXAU4Lyk+rcWALbGUSKsKO5dDYAetGhCbrnmO2cknBEUBzwOeAI0uY5vABkYY1Ag2KUkNdbyN
CQhYS1Np06t2YAVyYB5OS5TgpNI/NqRZCV4s2EnCRyhXyXm5HR4TcVxW+fvSaN5av6HlFFvkKVfX
+9ZA/gNd+UNWwiMOYJTwd0w0IYdWI29Rvy69oAbAT8qOzBbtvpQ+SJFkX8AUTi4i7kcAJlkto1Fs
UwNCVG8LK5hKrbG5387hTav04Q/dPJUQ/t2yPzchgpSFqXsGXVAdtSB53x8aVYd1AJ8NwsYJQBCo
M8CAuAK3rgJDQmkaf1FDSnYKWCeU15T5Tuettz3xdc3pmTKqHzCBIuJw5y39xUomAmm8+oLRb2HX
Pbg7ULrhE9PXgqYpw90EqaLWmptJJRp9wI6kCZsIVF6r/mmZUhCd2vTGaU1HvmTDlmKId8HmqvaM
aOa8Ejs1LJMam2B9KTLv01bb66Wmgi7NmQOzlxGToyc9SFw4gXxwnsf96EpUG73x2O6dSnePeHa5
DVg2yo0kswkFNyraKXIsbqnEm6WEEoIjgfUT3adge8g7a65BVbvITd6BLTqjoak3/Apov+FSMJce
23IPn3StpPRXTTJsD7ADSl+N4gX/f5KKgGwZC4ddCxxajs3jHZbOHhQBDKjE8P88BzFi4W+7FX0W
UvUvk67yN3x8QsyCdfReoxd2JBsdHPSdXrZsdvdeOSaY4Cehj4zMFVwALleJL3z93vdrIHuQk4uA
8/YdzCUeY7FIVg4pcqjxEEqSJnGy4l0VD5FX0ff4/ClXVhRc1CkU9DLHpQGYl6KQZuJvA1vDiek1
8HUE0/uN2A4ae92D9cEaNpJ75A/R6X7cP8Fq7VPXfLmIezzc+OM/0CNb39eIbIkX5wvwmICrve5/
Jd056fSLAoM6yWZNKjDkbb1hB9LMNSvcIjA4XYZCau0HmLNrlMXjuQfC6/3PQ+qGIwgFDxHpzWIR
B5K0jRec+7ceKZfSLGSYIpQptVa0T7QbZRHGDjY9NAFtzu1TQswBI44ipeDyhe1XWyR+gUHPddR2
bNmnuSCUfydrYDe/sN1Jfld0/ifdj8oa9z2mOWIV3r5c7cDp1kwf3DnJsostROjnAja8shtT96sT
7+jnUcieJp9Bpubu3mhx+Fsh4O6DXb7NJqjaV9AQxkblXs0jLK47Z/y2O/AWweVl2qWFFgcJu/ol
nMhhGBEn5Xp3am9vRvMPGnxOGoKbLRf41amTL76QqyUm81iStIyneENtDr7ndGY9uaqeIHLDvMJt
75bo6L5WSuuY7r5MzUfiQqpP22oXnHQ3JZv/a6xo/WD5Kdn9bbVLW6aAX/744Et1qM4Imb8Y9FsW
3d90zws61luzeJ5QuUvi7ngheK5pgtYwHLhz5zW1myFlgl1G03BkwRbLvW/8OXRvi3jHGu4aJ9px
cjgYpas/5KQ7cypYSE3XwGPwP2bUqaD7eZB6W5fQ8ZgB/isA5qXlWgarpewnwpohxLJO/ZR8KOK9
QGhFni/j/34wuBZsnXTrfxoeziwxSRfBaaa5anXsYbzt46sLt42AWAvHNNH+NrgWGX6EvTo7DQEd
nC6JRUDqpdYqIg1wJZ4Q3oSZZgptvukMv/Sm5aOcefehenozD7cYScYBzqgXIQcnzykiL218nTgM
a8H2It946R6oJOZc4/bkrwdoMLOYI9Ux7aEJAysCTjvMLjSPLuWxYjsVb8oFxd8+qA/PRC9kZmxA
nH3mRjYvTXe7E06/jjjFg6ihrltGYNrOMVbUQDVwNMJrgEhKtSk4qVIiIncHlYAbquY/wyvPoBeB
stzlDAKijWoeRhySoE7f3KXyZv4uWqVzubmjd+KF8jUsgoUctpRYA4jeEXSWxES4oE0xB7IcgZmu
OIxqX1UR2SIkutB8ZazJ7Lu30xGMYLY8EfnzWNog6HxSzzw/LD9NSQb9vA0NTF7Mcw7Yi/X4ibbB
cNRw/5J0YJ0E78MqHc+DpTpNQFSrPOpReHXMX48uVriZZFH2MFuBoQio0yLNDLxEVY81kPDJNqhR
9yxcovyjo478n03U+E+Qd2wbX8FCIMkXOSszErHZoOYOVp1DoxLVbutZjLAIxbvUSUfwBB4z88F8
3E1t0ft2g6HMIaJIesCnMy66H8W93KrGCQL0mRCjL/pPb62sZjFq8MobSIhVsDv3nIGv3NmE2amw
SBW6eToAMDABt8oi2S7BQ0FfHutnynF4BStkdUzZmngoBZC1TexlHRZ/1Wosmwt7hlKHjh8btkut
sgGRgu7F1c7TEMZnwYWJ7weJDMdRDo2RNqoJ0ZJrl5T+NV4oA9SzRXmyP53AorhWROaF5QZoTTVX
XHUwnEzCkLVKWmeaz2b+vD4OaGBHC4Terfc237EPdfIP2XaMSYuobp6lcqbTnvZejW6KFMQ+KJxA
UMjUVUB90SK+cZuoTRibSNgh7WWvL0epdpQgjUDLmW548+wWJO8O8laH9P9SNqqp8qu9UTokNXm7
jiNgM47u2/W0NtdcrPcD6em8egqodjz8p9iYXmmTcoz27qvkiluTW8fKUijHSVUivmWcTf+jtlLG
Uvu0hiv1yDCqIZQmpLyXyyAh+cEI82aK+AwiKzxORCx/02ze2bWUel9cpW9WEHRpG5dCX7SUXEQX
+kyFj1SMsYhi9kWBJp0KUSxCgPPovRkEruPIZIP0cElpNQ/bSRb3WeN5OJxqZzrNdsjkEF6mvTQ1
8XAtImy3Tv65phPW1E7G4niAcjcCBaO+sK/5dYdJdqAaQuEWyxHOL57nnZaMYv8qoGonGElKWi8G
XQR8S40444btiX8wRBNKbPmcEodnJerlGuuc5xhYWTvPNKkBeeLlCoxX+1bpRbOKzE1iHgyE8s3V
nX26va7pqyr1qbysP4B3rkrmFINU4aTlw4E41P743cYhaJWrKzrFh9Eft3lRUW6bjqYgO8eVbW78
7fD4H/zuHw7hd9FAzmZ7B9ILnj86KuN2/6HpXfJkXN/3WdFtNJxv4DVqrhQ92WasO//uSjcU2Uz6
w6qeyhczpLKjVz2uAYv81MYGC7tOhNvx4AAM501pBd0/dIxb7GiaxDT7fU+Tu6RLewS9IbMMa/GD
WwGaxOrj0JOTS3wg5RKFQs5ydDZxHTlVMnGHLSvVhqUGDLS34t76d307r5TErPNaIbnvhEnadkgj
hMtn3XKO7eOqlQVbb7EidetUBM/beBJAN7kt8tn53w8VBAQjs95uw18jwKYW1y1MSUYbT4SP24GA
4QqkL/HSZj63a1EuKdu7Ta+yQi+wZUpxMGRNPXS5xkEDdp3NojyHdOLCxGaofMoL1dBXHSTqwA8V
xZuIPnv/vcwiOheOcDAw6SsriFptgEZKEGBrUwKN+cx0yRuaVFRgQwzoULu+RiJ3PNoaKxLB2vzF
skJMdDIuKqW5xFJK/JMbKKZwK2B8P28A1UTdDKJn3hU0i6qXNMcoB4gsUFTJrBS5f94BbkXWK7aW
Ad5vl/OhRBIGXKNb2xbUBLzayFb0dM2JNXJv4QPgvkeh1u1FmTyhRwAdb0JwWLKR4aLNw80EQESa
KoYntqp++Uv3pEWNaZQuuozKtECmV4mLKCjH8dPFfZJXinCqo2Ons14oGfukpP/VqU5enZjrfWu1
aMVPEdgc3ovt9Y4uRI4s6Coji2PiPFKbVWIDJWfNasfUqsjJJIanroXfDeD72e3uU3ZJhv30n35l
i0JD3huEhrk/6BGDgj6XXxRcRI/RcJu42ixyHBrkzGLKkfV+WlYFVSIEccShrbM7gb6fEiIbL/6Q
OVD8F0jRElRnWeZs14IDMO5XT4tmSkgR+CuMUFt0eHj6PTTqWmbwOH8Y13guqRA6znZ9VQjpVO0X
1SKjApeAyxhrJ+xtkARbI6l++fXBE93aoFD7Yfp7k9rBzhFp4HiHTyb96dzDycgo/JQRYWvUImoy
QneRfBEHxv2Bb2XOt4UdCjSRlNCA4vJwtuwWDvKGuNUZrMHj2QfhCeyMR0XrNjtRrVmFtAp+d451
hmezp/rZUg2USbUET0ViP8YIhhDyUPkarCHkkJ94K8mnr+z/bzmtTX+ss6OdJeMusF2Q3Ys/7a32
tx6+nYc2vRvLIEuJ57JZWSHU1KKX6KXJJk4ibJOyoDRZN0nZO9xSLf9Cj+l39L1dV4XFwXfGQ4VQ
mYLlPke18GLRy0T5IZ1TwfJ3nMx8HzK/NhzbzO6M0UGDF7TrDLa/FFWK8JPj+Tm8g2d0P56AuiTn
fnc/pOJhEYzTpBBDixxygHo4LaiEjuSffmQttu6CJ1QOB5H2zqjgJ8PkTOdTPM1ichSwRQFedsnY
SNgHoJ0AbbAvcu5pX2HWHk5Ssq+yVUSK7bvjXNuYwIuScqxkJ5Gjd8Bxuarrz1nkBZjHSCQ0xSIu
iaSzAsPnmUQrrW3IW4+BwVrkm5Al80OrcFfaxiWh23HJU4uu/TIkOm7w0xM9WTHLxNKrKi9zLr3r
NfCkQSKgG3Ln9drrbzdJkuYiOpZsytEMbiOzJ/AZQKvJ3FEWQ0A5MSBC56UcmZd8ZNuoV01Xb5qo
WKW1UEmto2ZRvcDewaC3IjRZIJ9O/sit50sm/K4FB8KR+ZCJtueXt1qQWBs6AIm91doghfbjxsc9
La+3MQQJ61USJs5vkGy0B3fUBs+KIjWlooZFUMgq+XpwgHpV2gcGcJFetrZyA8EBcjjxMX37Kx/U
jrQLall/MjKyNkkdCh82nz64Cv7HWQKzQVDDE7aqPLcDrHrV2rjMhaTyA0EBUr91rDaGIZ9MZ0ge
oMQNlIs2yeL00LDNO0AUFu9Ilxo4n5sXms7f4Kf7dOeyfNUjcBxqEPdoeKhtl22pMzFSy6vpfRvR
6kf5wAc9yXqcMEKuKlXcxx0Zn1kVeFDWywg5jHve6NoyPlC+mdPIaTcMZKkTj0xCMZOMEy1CmsX4
OBMQJ/IM0sr92LmhWq1I31uS0b3Pd+1Ct0ZGQB/TDpef+WWZrX+Gv1rQuwTi14ndLeQv0SuNlQi8
u38YYuSsHgZ+Q/iIQWJLNDbKb1+8+dpHeDJ6E38U0tOQpymD77BmtSCRtJv0B1nllmh84emfle94
2mBMsH5aobyE5lcTUSLmca+GGgxd/Kd2v2Pe/arB5eH6URE5Gv6Tp+dTdLcxhU0+9OQtoougH4fZ
WvjGU17G8uykU+17FDrzPgyEuR4KMXSqY6zTw+EJLNyFuwe0GwPTkbazMHpSIhDU8lvhui2WF9+f
k7JTg4zoMwRc6XPcmpl3/YNj3NEx8UwJqaLDpoREb9maNLGJXypSfzKfu5Om6If6b9WUeLkJwAug
Ph7Tgg51t5H5MdKQsn/D+7YAWAvEGYsSvwuHjDSuKvuyEaYz2Va4e0gSjG7pYHmnmPdIePNAX9uY
D2Q1BXQy8SFLhwk/SWXp821XsO8D/xbRaBR9LlbpcDVCVdk+S0GLD2qaAPnDOHhOeWIaN9mOh04U
SerONlOzOaT0lCQa/c39Bn9RkDgYU23P8dROYoK0iE5tKZwOjajlurZ6kw9yvWsINzGIZb4eh+C9
Sp6HiY0xD4j2QPA5WkokPrVF2l9dYb6Vjgzbzlb/yR4e+0heRD8Dc//FXM10if01YANFfUTnxDg/
0gyvMNkLLSeUjWvnnjQyDsT5Mvs16iYWdQ10LXQi7xVhz046C/Xk7CzwifUOqE5sSOCFh6+4ETO3
Qb8DcsZCwUacfyzjU8ViY49Nf1+q9DYbIJkLQhcHSYN+H1XOGDK0NMr71SQGaxCxs59Dhwy1Y4DD
lTZx5kl/dL42PFORvZuvPJOSPMjD0fivHuXEy0YbOUVzBkjtnw4W/ieEEqhwKW/SqAqywtKMJ1GY
k9AteQcufRf3e0YzIAbbsSRJ4vBSFyjlhrGmwNYVg/0dBYS9rT2vR3jS7CoK7CZ7n0IhA/b8Rz24
f86E9CVIufbF8gvchPuItdcQC5O3aNcsOE23gjMoihAk12Nu17DB9+xkE0zyjEFEeTldW0vpxnbf
6qHMW+6D/Xb+aBqKBjZ99ryJNpI8q5FTfPcmKWLZsf41m3TCd5qhVAm3K+r89NDlL3BGDg3RWiHw
a11DTSCvNliQxc/Fz2DW+fk3zPKdA0bb70EP0iKW0IJXAuI1TyjMHlM85SJcGD03dJV3rSflurkP
KMY99r//YfzYXguAIGce9Qz9yBPYB00s1AngCgxkVQbbe5HTmmaPA6py4F6z1dxeJSHYZiPcBX4k
puQ9KyEfhhBJ9t1Y2a+DPw1oYbqYuThwkc8A+HIhh/W0HyWjPJLAzvZC7rywSHUFnFdwEoWy6tUs
8s7u7kN1xobHSOpeXEDPakRqlZRitNQoquy724l4bTAEt8iYvIRbTCVL15bcHrJ+42IZstAISxCM
gv8ADmg3zzx5aTyOwtpKALT/GUpFcWTNY0lSZwU1haZqo865SCpLiUWGlJO23R5uLrgibKj5BjGf
Fq4nD0Lb7AtSSmyr/j03UJ3VZOise9WEHkdeXSlr2EV1n8MnG/nH/JSEhezA8XC+qy+AeLNu7A57
WLB7dqpIF7lHOv6kba2j5VMLtSihYJcTiHTERr/6+1fedFdVGm2TkRRyI9wG7anUFT+W0p1mqS/j
KLK+4jSDNOXb9J4oS8Bhv3zA5EmU0EV6s2HoixkDRT50Ff8p5lcnFrUB6LPxv47yKPkphRsBhjh8
/KlwLJKD5gVg0B+ZzB4qFxHHQiLl7jSNonirkO+cJsLc98hD5qSm+6W+WmB7j0nAuujH54btZez6
yNavW1gsFPqVnRYnF9FWC5jqbUztAqIBiu0GMysRH7cTdQYmKwYHGDT7htYawoeGPflzOunzW0B8
onYBDeSPGVZnC8FIaLI5K2sfBo8COFql1MgHrXBMAL3POxFyIN6i/oVFrAwPf5j8pfTLG45lIpl3
2H5MzlBq2RTaa3ca0WMlE85W+KG84f38buj7BtXSQ1J/Ji1fFEGkxGPADV1Qb7s051M69ZbOgfjV
vdKxyFzyHjrUoYFVFtQBsxnYazx4VSH+WR+aWvck7t+lBcYDLgjX9n4ei4EHFbKbuCvrOdlWcerP
8OsfbIcmbSXjryILb/BrJX5zll7xx1EwdvOSY2HStw18CJ5F5apjzHV9O/ssBa4R7iMo6KxNwo3X
MDsZ+c1eneVfTsp0c8EIzJ77M4QF6dIizCAPgwsruK90UMsGoZtS0jpuIzaCytluZt50/tJqyCer
Ux5bse+gCQY62gGD66NjQ3ANHR11YXcb7kKQTfijBPhAHKrZS969odT6djUVQJUM+trhSwhbwQGn
qlfkbcpilEGdiuDoshQe0RMh9VjDxvtlV/7IlVfDxoS43GjFC9shhbOPfZZmgEjldulHr+oNxRBf
A5E4KiLDx5EqnXL8PYn/KjT1GaBqnko9njqzMtIJk4KBmsbG2P9EZzNStoOfEAzM7QJ0kLi66IIY
PVWDMnGmZrq84dpodXGrglSG0iXgewiYlYeNu7wNXvLJg7jcbckXf+bnW1Pi4fj6Zyi7eL7Jfl/9
nsfCEFXHlsll1NFTPin8ZsnjApuoOwXQcgmsmGydRI1jIMXmzq2TliauPk41szFQqvpjXmkgXPat
V+SJApNRR3ZywHIjispNbMWzJqVV+/2EPJ3zNX1KqPZ9yNGqcpfca1JmnRoNnmXs7WQqr+Gc7XJW
QcwoZnolMcVv0PBR3ULECApVZU8LzZ4BhCfo7RcPiASNl7XTxGeSz1jXOx+D88Z348S4/XxdHH0f
ybpoEJRNEQlusz2fAZ8dxUpBIZuwaGdI/d201Nzr2/sg1aSxGO/APPzm6KZunUrlif7W+ox1JF/H
vEiqMwcY8z0eXvW7H0EWt7SF00lrLO/s/v9ZzgQAq66wH39iqfqHEhl6TLCi4jrMn0dmFbDxRRtI
a3mYaN1GSsNBUFAUx5e17n8ruttn8QzVh7jl5xPB/hMVhYV5duyE68hc32DTFAJwj8PLAporNfss
fDk5t/0ENYdrvQqhpqWd9OQ2tRMHYja1IzGsHA3jKuRHhloCGqn6C0Jt7frmeUjLMhu91kiZ/gny
Ftv+H/f0C4r6ULPZyE704uk29w1OnSsxeo5FjyJnAJhIJdNTYDjOotyfmOkpLA38Ij55VEqNhQeR
fz9AzA61uO7mPCfSdVbuWgUSnjlOfCnFaxIZqYsCuAzVcezNsryNiFou7xPy/ln952QhjNFG6ej/
QP17UUdt/fc967WFO1JDDTUh0J8wsRJssKC7xi7LSJDeZHd625KO/2pVtmPO9gEcpzPmcLzsOlZw
NZZNY5EIVK0Njq5Q+aj0N7tfKwbtGW2Y+A+5SOKKTrCgX93FM5h+dwpRHXNSZsVaGyNQ9RbP1ceC
qXwlHk9dxKCFiXCpf8JeV7QRa3Z5Ai4MvRr4elqksVKa+tZAOKQI6C9m79s7VVZ4jHInJXbqWP4p
aCRQkbzLZ7R6vzc8gyAnNPwXumM0ltkKzXS7B703c5y6cyaczymaAOyGNTINMzG5nn3TFACyTNri
AzBZSJ8CvjGu6Eu1UfbSliPHciiiDgLfmkujc5mM7/hlSSQeo/AtTXPlb4RwESTy78GC1e//Lky7
R8ZTWCbLJOhkQgrkYJCS8w1FH5QG/bqCGS7Mz1/JMO/kKI8exYT18y+Evsfk9xMwG7176UIUpKNJ
Uh7bkVI3dxzf6Iz96loejZFzPOzGhsOEKVjJrZmcrnpki21e1MkAl3DFCyv6kiU4mNEXguvesz5A
1OcNQDukvA91NquLVXeI80QZ9ydVayWJD7SG3uSqFGtgliI5Y+uUgKdk+D1eektwdKDblryY+f8v
QWKR6l/Kzc5DkkAfv2elcCk+I4/iIHBl85rxTMlqZ4rmNsqfxJO74SEoEueuoxRegsq9xd5qqC8a
2ZqObbYBBueb/47+HCcsXCZLZRw2uZW84Jq6f7VRUrvKjNT14WGuayArHDX7dsgTXrlRJu6rzpFb
XyyszHyoHZRQ3XBclkGO/zPcBzMQvf7D5SPYJLB7vEYzBkxEREsxIDv1NQppP1UIxSu0Hht3Y6eH
qlmMkobMu9qiXzSrMQ8dsj0/PgYeDbAwXlKQkRhZblPxCfMl9ZqUKdNqltChA/iV6s3vd7DywngF
IcwuzSYQzb1EVheaS1RFemXxiZD/Xfs550AAAHQzd/g+m+dZlCoBl7XB1HDbw+rsBGiI8pA/RZiE
hYdgBcr88EBBowpZyNTvZ7tYfQ5N3Iit70EMAYhw9uI70LbUdmDYtAVdWSO7Skfp4Gh1n3HjyvHP
Czz/0EUzbBh+iYblUbUzMG4byRN1srt1D3ZYmPTch77kploj15aHvlR2RBzdRte9rlvo3xbFQGQC
M760qPs/w+2Frv0M9j4rGxzrLP82DNlsSdTp45IM9JvzCKCAXaiq88LQXOqHyA43/7JM6aGD6S/f
wyJ3lYDfOYbb/wjS8akb5Rcw5Oc+HW9YscbKqibNh4VStqQQEK0NGgOoGiWMCikbnyjCh7pDggYo
FQkIzvN8cd2H43rex7dzltfUIC/Zp1wMzWEVzJ4vaYI+ZqdFcFQ/k35OwhqyXSTdkbZ/3S/m+bIe
KOAK6Ivy3YBA2gwboiQvy5xxh3bJqU6q1DWVSoBwCxvakDD77HE0ydAOuzvHNpFmNtGbg3V7rolT
2m8m3+wZYIRvBtlYgW67JNtBKq+N2zSc6KBzg0C2c8a/DvmzdXSZIRsJdLOr28JxgSunLEFsafPA
hxlVPZUNMqBCjBRrFYjPGDH5xPkARgPAkJUV+R6MGo3OsMuSORXWKOTfO/Jf9i9VbvWG2+PBx83r
WSp5rQEwQRXE0MlIfiOsBS1rf060ecVnoZGG3REYt4YHfDrwacHwiwQh8j5s4hQnaYxtsOVvHNbb
Ukt+RiNntjsJnq97xxeK93DUCoJJzY/7hDir+/bG8fMRdtUBguzasopaGgW4DKA0UGs28vel427Y
Gm9RHzK12i0MBkKOqKU/NMHlKWSuIhVXvKVLXxxJTos8sUbK0pspUsZuL5EgSYhKsTzS9ntkXVkE
CjcrxHtj8EZEahJkbKErmZAHOHaFE8oB2+iJVyGtHG30NTyhbLDqoY9/fhnKGuOKQ3TQdNBRono3
osMIu24Isl2is8Pq+YCOovIz6D6qoYIea356dETAokKGddas56+lEvMn36aWQRnJEwSoLVV5xrJ5
QfTJglNxj676nCuZ8hP8ewlMm8SSUvWnQP01hBumFh7uUFR+/IiF2KH5uDD+nDRP+tDpHeqKrA13
cSQC7q/pnEliG9yDkisoCcHrpBnNHWKbkVV0orIHS3xYNeaenW82Tds15znV5v2tBKlp7e1VjrKY
TCPQU+OK4cpmGyjs1v92tVP0dh0tuSx+bSXoFeHnEzfQvWNYJVFAgjFqdu0u4kpmUJnLsCZKTvSJ
yJekolnzVgH6iCVZah2GGLgCAjnvjM6y7Uiy1ATg3QSECWCCeHy4BmMsxNGjL1w1NCWrOffDkOtl
X86/hYSTG0X22COotB86ijhT4/MajTIsGyN4pCQZX53K/7+WYCMwakWX/WmeJLG2xfEWL0L2/iiP
t1TeBnENXNpNzsDXwdYkxFCl4wy2Rp4RAgKBZfYJLXasLBEeumGhpcctJFAsbJjdlL87fKreWeBr
ZeUwGeGSvshyZC55iw4YBN0AGpG067+LZNlHDmZM5x6KtNfWZHBX8+zGXJTJ7sfWOa/gaxCYBQuy
6oM3+9nRKyUkvHPNwtmJ1Jr5MidSqCwG5kQu9fnBWFswnTisrBGBRoum1sX8XutLpMT4fz1p6N14
4puekM+m09kF3Upws1LG11hoqarpX5Yog4SjIxc9Es84eNDJwXgfmuF7dvmvGlGLXtP5rvz3y1WH
Q9mZmz49hI0xKhdPxdfTF6ehYDB5P900RvNnzPcKHKrb7Yuv0tqa0Trw4i+otNhIGsvaj1kT5BdW
Jsf28EF5Med5QFNhl0nANGicArj1shR9BOFrOmCPpQBLiVb6vpq27ade+JTMOoFxPZssNd6hfbZA
IOzLdgey0GTL7cYm/8S9BhiRGFZV2vF298OrqqCMHSAuKdhJG6mOZA+vL4RshowcxeT8D6XzrG2c
9U/SJGbvcZg2meG5UQ14XcDhPyJ6ehGU09f9uqEAVa7vqzV/vSk2o8U6CIuHBFj3PXZDD0vWn7qO
gUUVURNiwTL/XgI6YhpAHO/2QiggWLxNzZZZGNZiNc98qfgfhK35akMP1JP0paoXYo6GojakDv0d
5AuXX+QfYSUc/mMav9I5Xq9vzLUwBhGNGJaExhIQLNjYTztIf+ZKPHo75jWrH8tna6Fr2QPGUqBG
ogGCXkNd/fpOM69RL2VNZt+K3Bo2VPXBJb2d39LC/sioFkJICJH57Kh/VE63zVnQXEFRbGaOZOuf
Y+DMWvwwxSLr8Lw1cIQc1pXq9lF0HzCuJzra2qgpLm6xpSbSQ/aWJjWBT9P/MLIiILLunes7URjn
wcea/ObAnRqo9mFOH7/AVm5gcCeV8nIFnfMxPR8Bpcb25q7QHbG91iQVwvaRoAN2ygGEjBcFSxDM
dwv9adWoCjZaj8to2Axz9wgfdLqdYvQMcLRapZHpFOFQ1ZQtPRYqV0g/ClBx8OP5HZ9H4sVBoNDf
2b450O9Lmscu8T6qVCIjV7rj+HdlbiM6STxRNcuz42WqVn0Q580eolbt01mmEGaa6C+dqeVduQyd
QewfdHBkokRYHg5aVJWvZO24G6/DTzBWuA9ckHctqJobb8UyXa4hrmLVwaXRYWy5SEXHjXbUa9ID
pYzAgvxtWTlpHzcArV6f3g2AIAvWPVigx3SGKmz1xx1XRxyucxuOGgGN6HtE7fYTdw+IpvTBBAno
st7Xe1CDP2qva+eRxnuWhuFtFVuaxyOl83ef5VoHniRDmUoDcrF3OTjOWGVeFlqTMRjtndD8dYSe
gPWk9BEVLRnovWeb6+inf/63Rca7Fxn20vIixkx9ba4m5zKLXSJM+/yW1tYIowlRD4q84DuUVuXZ
qFI9vV7FcqCg4aKx4JXifLn1gzw4XJle9nhXyamJBIV+ifKcF/9P4lFO7WyJmfoDYNBf0YiFOra/
TaP08OZyeV6iVZW38JpB8vzifY17CIMsuHhJIuupyKqc8L9tHrEZyA6pgMNQnj0mOVWPzogl6bF9
JLNbffgeT2/Glw0n/mbAyHGqwMLTbyfgpJqjIBOCs+OQPBseFX+0qDasneHjvBHLFCqy5nepLFRo
O3pLbQaywKiGReBgJP+c58dUg2/7B5fsz7F5QyZnpE0CywDDsTcvjKMBjNgi/b3mcW0tw6BaHDVG
NTJygN9W6MXfMmq4gu4oc0MpTCcmqj6j7SEzilpQbB5H278jv+xpFN5lJP5G04vsR3stCfbH42AN
PdcMOfkk5Z9VHSRJfa3ehQugCDWpwPBkr8oG4V9O8EXr67ogf0IIzCMYch29BNSu33+huTHLSz+u
9wvdAaEwZiWHldypC8WHSL08O7mS7WK0f50rrBa2g/y8/m4LBuFHjMFyIQ5Re9xfWtCLwK9TBGBE
KDe98+WO6Rhc9IH0z++FjAhBHR7e27lAsjfRvQjuKVB5MapUpp51R3qAnLQyClOkkaB1g1+AAXFc
T4L8gnogiYt5zxxABXfxZ2nEzZjTViDiXBLEMJTKqFgImXvA/fx3rGx7MTwwIMuW2xUp0Rr+FWFo
mQ4HF6L/7KBQkO3bCtgqY6REyINtXo8J/V1+PbqvVVk4J/cwfSpxS7iYxxAbaSmtTFBBJ2VeGI9Z
Fk5zCicLVM+dzb4NGCEl4afxZIxWu50G5vwIqFR7EBdfOlRx0GW8jqDmVt12tCBs8OzLmDGmlLAC
g0atg/HhBUjjeaBu7io4C0iyCkm5L4WNwAsjDz0AbbVjr/EY2HI0GB8LxKF15b+Li5pXyxJA7nn2
wYAm7wmQITXIhXkJQHueVzGkuUs+1Velz/PC2SaBqi9/lMqD1vUC6fYZu1W1TjcXzljGJO6JMGEP
QL78K+rMs1bFh+y0GqJOXnsIYDGAYuQjSxQBNJmEkfRVG5tzD/Am69t/l5a+zniuKt7lhfDZePwB
B1yDuGPcCvWYznDB1wXBZkU4kn4lxxbxmEXryMySGa73pNQrYKLkbggvnNr3mBfRAHWV5i750iXH
tx4m8Ix5E/MqdXeUlu2Amx5v9AV0vFyIymSQcskZNtbJJhdmtOHOk0jv7aH2Fv0ReTo8cCd2T2BL
a40MahIigvE249F44iVxTzUjz7fFDqalSlrme45wUSrr679mtOKHDb1ulR4baoQ2GGplwzDtGhbv
l2xirHSi9vN1c1yovzBllpTt3NgPLuyLOLSfC/x9F1SApGLPzCuZWrvcDad5Od86hR+DQklzi5iL
X2TrgVjvHTN4Rt1l2O9CsgQdVnk0CgJWltsZdnDK5o9LJR6VNrz30o6h+76FAk5NTTUW1K2vzx9i
/0sbMJE3uv9LXQX/bhiIekh2K7rOageOySm77cFoEljuPR6bFy0A22ILaYhyuOwyhm24K/h29muZ
/sDlK0qaQEdFKwxHuxEytbyDaZi77h97r5VvcsHXzbHNerqBkylaidGXWVZ9/CCYWH8tz9RqVOG4
Gcb5bSYCwimQI4TBU6GvB7smUkYe/OLaQwYzOEibCclWXSDNefsIBMchBl5Jr+q5FiBI8rhUDVKB
naugtcA6MnAVvg/eB2zUKoa18bPL6xYWUiapjww8G2fxIcU5E1pBVEb9nxOsSigNoPUox8SuLicO
iQO4dusGr43ZEwvDCTQtLQiN6tZauNcG5E564i4GAj35T1WgbYhB8Rni7U6+MfWztBLiA38pOqBW
XKZ/W7KT09iEuNTRZpuN7IWruSyWZTYyjZ73j7HzU6ET22v6PJ4r++Hp3mKB+gVd3Al5Rbs6oYph
qD4dB10kUIpy7rauT1iQSgSRO60pNhHJIPhIGxHMA/4aavxvZUGiaHhD+5SuHzyMu0bI9eAq7csO
hYpEw7BeAEzn7e/PsjaV1jwe6W3RdDC1FRLOBflUOEixvjo66DqcAth2PK5BPfsdXQcR3Ymr0SiQ
2Xo4a/kWTB7uLliUBWe0WAiAJOwVuet4JcP6yHquPfJnuT+Z/6ahj13cFJZW/KvkQCT2FUb2cRVn
fuM+0q5RdmxRaT+91hut4h7UMvvDSrvAL7YA7V1N/DA4aMpBPeUfFT4g/LQGuzWe1J9ZeCLWC94/
l2WK2FzNyXYbMo4w8qKSTpebgKF3HxH8l5pa1fyOneRLerxAfPXqjJcBrVYP1Ce3SdN7/0a/D5Og
yCLdSmSh0rN8R45tZpz/eW1l0YdHviP1zmD2OkKHGmLMzlERQADGUr1sF9AwImDwQFywGRMJmMNm
eN6ARNTNC3BM409ubZHCA0H1HdU432bZ7gpBUEVufp0rUg9semsdyWzipbdTl2jSWkDTbGezs6SQ
AN3iPh9M6kgA0/tJ+iHI+g/NDpJY0QqEh+zG4JqBVUroOxEzIsJFOO8VrUON8g+PrUzLyE/EI8Iw
aXqVUAl2NSui2Q6cIwPRpcWHfMHzDMVxtjPK1nRdwr9YIgNSilPR+FgHsmDozgll/OADtby6ZbEa
T6CBTjZRZrHy4mGipjJnp9YknXCN+0GEFiQr8ZCo2DLMYDAr/nrrx9NlMlNjupE5ekg/KkJiLnOM
vfXSSHyU8yMmsT6BufwAj9+kGPAVVXdAYBWwFOm7tT3sI+uNjJ9Y+ml/cFsrPNsuWhfEd1099pbv
PxbBu8zfLDR74+kG00MYZtEhBo6jb+Vjnn+iPSDY2J2A4v8hQA0/6mmoneJUIC9q3IvPwVVXPyQB
fAvTI7pGGrIChbc+pEvrF4VouPVrBlEBcVjpAqyiAUOBhCs4h2BqzKtVoWEzsbrDB8jvnORKUVPq
KN8y+GGXGqMxc6P4UtJ9xorRFEhkfitIk8NbRu5M33PZcfWJIh4XR3mW7qRmN8frqzKC/jWnk/rY
SsDEvxUr39cUs5Mx5OFU4iIlZsNqqPMM+NcDum9rEbNfqvWheaL/CCmxI5Tu7rwTOaKsFG2MyWBh
/MMRbvYbZGaLWQOZuUSSNeLSz6PqiLw/MNZaIBzzwS6W5tgZCXkb5IJKO9PwU7J5PcOB47l1bWIQ
HWAVIef7zjKCXjpRvgCuVoinbAS2qj/AsUw1W24A7gG007AtdD3jPzogpaRrI+6yp8vhjOf/TW71
Jguyv/CrAEZAB5TOoL50cMiH3lnXrESned2KUv/KZ4wwATxefZBE1QOF5FFE3hVFVQevdjtBC8bs
HTfMgA8z5x07H+cqDjwP7Ecgk3x/IYDSOfWhO0LeO/Hfe0kwHmzOS80J+GkzzJ17kfZAS+2Wk9Iz
rlzZ8Doo2XryL0WQEoeBwQHNsHd173M2KZOwgYg8DpwoxcnkJRIihU8s3sjDtKX5jJAr6Z4iMCGo
zXCSH8rvfywjpGX1C9zlLIFxnqom7H+puiNe1auaRZb+u/2llOwWvjyArCauQrSSK7HkYX1PKt+p
rw2I4Mt/VoY99KuT2oBh2tyyJMvskPZBwiT1f3FmZX990nFVwj2YwacMu6UraX/DabdrQNuy44SA
R4XdwMzVUkh4CsDOigbmZKKy+MJmay5tp01qxcOUzXO4cGhGccDq/NL+VO7m+Ab3cO9h4a0e3tuN
uw1ZyPSZKWMFICTz92cZulyseyIQafOExvB+LCt98jwjtM6vFBpx/QhhXSnNVtdrbqCz6/dP3xDQ
EWV3qBVa53nfcBF1HexQsOYdqAxHADuqjvrIF5iV8hOL6LrYpeWz0a22snB1/KMzL7Hw6UjCtcjU
zvVYTtHpfPKkO5Z0Hh2lmrxo9IJXRG1qe5bEf1JoBGluezIiAfGX4aYyspzO//PXqFq29QXufRtH
emupOuHtAMVLHvMO9Wkmpk84e5wYXDf5gC5vWgkX82+oqmIo9P08e5cm21KsT29dQ6XNBy69kMwr
dG0Nd3zPFSAwU3lOZLWkykDRdy0kBbgbcdRN8UvaUEOB2FNeWa616XtsZZrzLzlYJ2Bs92nv93mB
XmWTqGnlLhctLfQwKeVquCO5hEi590xGJIYKRZsWy9nLNEAvpud4PO0Hgmkg06LOxIdO2B3FqU1e
HgHbe/Ue/8O01zR7rD2gVbeFooJ+mGBIDRSOCiBoFHDb/h595DMtz3uJKXWeaUffwWnyZSgUUtVk
WFP1SwI7rFR0o6NW9whS4JTU2fN9GR/OzlEsWrdbSWwLCztRTofDxbaizKhQzwRyv0O7JPV0zreg
2S7s7x2lGtn97gmPiXQOmC8yqTgAibUIvC+0W/1MAGFmA6CW+PjcPOyK54PuYi1zbAio34fIql/w
kb0EAo/t71rGKMCg5FpZVYl7EG/xBYhnymVUBGlb/frL/ZukotjtG4S9xHP0SVCLcr50NfDsZG+g
uHg/H6UXiYdMAGdWqF8ULXh1fnoa8A5PROHZo/y+bkA161h54GWYM8X6vHGWVtTAfFSfF/2wzbz+
E13/PsbM+LxG2NN6/FjZ9q43U2I7oZ1Q+QIhlCiOpCuy24V7lwJHKYk223jSHdhUAUarAmIBF/Iw
y9riKIm8KhA7xPEKejuuo3h2mjSfapIl10WF58CXfyQVUYFVgWgOORoi8cgTX+aY5NWnX6LgCfmN
AxwK4oOms+eoRJorhU83D5w+SQrZzwA198KMlg9/4uyJQEEbFuVUTc7R/ZqWf92iSLfXIkAf5ANq
AE8RBKnLhBTQsn//ZBsBRMEdGFBMUKmKI4VZ2c5cVLeuVoJHlS1tORNggwFcNrekzIGFvD+qqNrx
LIxyNFQp/xo6nK7WY98TkeiFoX8vkfTB5j762tbUrDreXc1S4tgwMFqwUy4pa6tjRdgQ5ifQmfrx
PNg2IBWN54QT2sAsBIb8OKYXLzX9STxU45xw8/R5/Kt1a66haBxz+Ws1quKFlN+qPwBsxna6p8Pg
C09esrkLNHZEQK7t3fuCUI+XZTOZ843MRy4gZhISBd/IOjQKVYBTTxTpnexdSUA18GUJvj7IBDiB
WlpdeNFi3gaUdreRHACoxeHu68amKx5rcgDe8ACTGeVxOp0nLVEQD3zujncdJBHMk0cSYAcfKFhz
Q9M810yZ6KBrF5aSYBr/odfBUkCosM+ftyrIJZUr8hKcecBNws22doJPA/ri3fJsWg0tikX7xFU8
RHpqZcM3ytgOwRe1y5M8RwpFw8SvLQNvI9bCl1K0n70/wcIosiq7vf1gw1pmidFrRurudX4AGu0V
uDm99wq54wh8WD/0gnH8qTltAissmSZOiSpUBHJkNIFPMvRuEKg9zXuMsUXafSxvzdImBYHz4fPo
lB5Iwy3/C8neZqKKW4dpdrystUO5yTyFl5RrwjzG+1JNTV0/QFJb4VOzkMO5zKVrGJT6bgbgmE7+
Ix9QNUl/7NiBRIGBVYMb4H25YFJEGDBpTj6FxFPxDBHkYSe0IgmugIEGxhGHr8NCPhckbOsPx2Na
/XAuBvvoD+0dQcrOm7k3hZfydS13s370uaUWhWbF/0bNUiDr0lwocwus1weNwKpg+Yzu04V9sfGG
6gRPk/XzVXFP+8HaxgTQg4OHeD4WApUmbGrNhVyrFQE5eNmsle4SNjS4uyXPUgkj+tzqNn5Tf52X
RckEa++6ZDHmMJpv8Z6r51XYsNcKPiTJbzYzpGZ/Qb8dEBHHZan+n88HM01E5xLHDjDdfw1SurP4
W3z/zb0lm6XQGAL4XqMRaUYcqL0bm5yuAmwT8ApQtTuaErJVqO7XWse9ZZ+oTlXWRiheKOYxySEF
uNRTDjqwgFb0ozY64izIhnr46e7ujQd4tEXVRERQ62zyjAnbqIlj5hlPBqggqdy9KMtjD8KzVCdB
Im0CQ4VUoy24w2tbBFWkuN1iYDSv+m8UKN+EETTmb6Rs7uF+iTS0fTeevvhGZih7K3Uoecl4+HaT
ZFr0v5kglA3uPXzvHEjth3iE9EUCM/h/TqDAg16gn9jrhY7uAFGS9x3RtsZYQB2GaahZzScQs3wT
YTfrF+1BfEBVik4ZzrkSKvYeIrogMPt2otdNDAVpSuji03Kypn2kqnO9DWghr0KuDshtR1J2XhWz
dDHRDxvLDNqLGl5Ew+R+huRhWIEwE818ax2CWYKqk4cyfyga8JH4k54icxof0tjwhE8Os8nY0hHb
QNWlU9m53+zE0RyrbBpNFX4FqYhFzU6UnMxxFeDpFaXkHnVLmHV9D+a9RtqM0mwjc958BENgvBWr
4uUK42LYaGVnnXNZV7JLx7GqFrSZHsYReJQJkDvV90oqC5FfI6ZeffCVXn8gPlR1U1kUwPdMm0tw
AlKeRTQne2TARcEWTZxQQ4vrYB80g4Ua5BomODD+/asxP5fnrTQf/1gqv0+6jAmpNySQV7KhgInQ
3Z1sGVAmVI7A6meQykAaRf4Tg1xmwGVks3Pn1G7WRlHf8wSN7r/2cQ67r2En58QUUtOBlvVYorij
KULqXUqyMDQHPzuMType+AeXVkECZN+1z+kObbZQ2/zA/2sEhnqVXjKACLrUnr6d10aestAyWG00
v9oJ8Ps4MykUAQgRurnJnsMfaKwslALin65fWTKyaSTpzd5UqqaWxVDwOrCCDRoI4LLTUIs/LbRo
USxBcGIBltTP827IM0zUHeMNXlEfG7WxO4JiozLQ1FlDodxqds6vRIcx+ggdWz8j6t8SscSRcd+O
gpf7t3dFkNdl4ATmB+l/FWJ7k1ZtS8fTYZLwX3H0xcevxhRXa7qo8X/iuFnyh0SvlwCBULnk2HRk
4f1BZ8/20wFJO1nAJC2WMkosSnGUPs0pIZzvnNYTYUb4+PSEzEpkn4IDMU3oYMZ2B7SgxsFfQFV8
ph8Qp9AtVDCuzWC67Cj/UsWJsV6psRF0KcKE5Ig6LGn2d8nZwTZskVbXaGtBDbVl2C6MxzZJDSTp
gW4s0GZZAuQ2UlISdTb+Le4mj0aGmcj9+Eu6bb+F9ebvHDwGjWL+zYNVkUonp2BLqoQAfGn6zmR+
yU4xDSDxjLTYVE3F/9oLu4QIhsSkKxicCvKhkpZPmq5M4ilVbGmn7pY5dM/wddzdG/kJIgT9FUJJ
xBdF5CGqyqJP/JNCejyYHYNvaG6/AUGoQ0gMspZXnfi+AYSnRIVQze7JprB+x+NpCWgIm+TumW7P
S7GYLKJC7aQoImSqblCvKjMz29WtaAaU6TnYlwzNYoAlNyZmMEVXql3DlexBcFHqFQrOUlD7e5Ab
xZOzGLx1NhTtyZR2QFtHsul5WXoOm9O033b/lvkzHEotiw/Wbq/pSE5KIiILE5zaxHz0haoh3gi3
q+TbjXp59D9oYeUL+ua1rd9wo79m465si7APKnmCtBpc3yy7cPSHWWjOKA33i089EzVH3sW5uQ1K
3UDcabOLDHs3d0qA5bjX36xU4U7T42/NJEMccwP8frZ/H93e/+4L7knvS9nd23jY2wXSPg0+jCOk
Lc0d/tcpQzUYsPSm0nqQSAa76JvyDmbTwQ+9xZ4dJRLuC5oJKdCQKWAwLR3Tirx26Qm8D2VfvcgA
4PSDKqDDTgQ10DJhX3JTjVnrwl2GtrVp1v670pxvXn7hlXFBsO6cl9z9j8IRDOIIyHX147dSYfF+
8cb/j7aYnF6uDsRep13NLz2GIUrFgE6flMg97AHSluZ5V0TM7lwB4RPpCLXRITQmuKldVu+i4I/C
yujv5/h6BYjEFhaBbbjugRLmRFx2I/gVc8xPRO13I2qjqLlgJnTBy1kTXZ/zPSGYKLeXqQSQka6s
pzbp89Wd/RZTUD7jgZV5g8xB1l9dlXaPhIT8Q0NWTt7pnqbVEFRn5lSPhzk/2u5Dd4w/P4I+QbG3
xnYVikFayetmjSzMyAn9s3J8krfc8ItRatBvrLARfaALvX9BeT44jkZ1bGsxGWPdwxB9pvcoUW0F
N67/g8meAUiK3Oon3zIvKPFkJ07rzjsLXgnUaS2mHZ5aKmIf6zconFqnQ9P2/pffEDX6XSMOjE8C
ugvrlo7WQfPGjzOgteibZf7UUd5dNom30GB80XC3aWpzxz0xVE7L++Wgv15GoKPqaJ+Ml4fdmgQV
4CC7GGoWhi+6pqjIweiFxDa0tlPPQnByY1TGFW38qSM9o7tLcraRz5Fn/I++0yX1pF1O8rXMIjIo
zU5yj7FwFv5jgoFVwpEY1lwGAuOAmHyOHbNbulDa0FShRK/ULV5zlM9nFKtgQneId4ScEWhBs5QV
x/3fqcuCG6khUAuVyjgRclU/7MJv/q23PVo1+FCZ0N94e5LHxNC1Hs2zTpz/c99BP8CfroRpZ+bv
F6ThH8zYlcbQR1IqDjg1yBOXCBWLLxi+oPx861+he4E8Nk14JnmamppZ0D1UxIC0kURUsIEgmezv
19Nwo25l66sPww3Xoen5fwBPtj9TlIaeNGdRKj0LpE5v5//3XIwhAfKlRYicpYQAuvpxx9wkzmKs
P+Yg55IXeiR8abLYxDEDvh4uqdqElmMUVVCd9KVK8/edQ0u8VNx0yagGsyoo5wgipb1g+JwnIlCZ
Y66trTwltV/3kxdXWfqqH6D1aeNcnEHRD3CAYbf1Gh/XxnaoD1k8YtHdQIG8aX7wpfDO45/PDzXf
uBVJyJ7I9DD5C/WI79M7p6cr+sAPqu+oJjI/DA9fH36kLuQTF2swZ7/rz33CY7waX0FvfbzUftdd
zJiyehHaRYwp504snmQ2rOSiCv76Co04H1by6bULBEmKbc8wYn3g/atC2eVUOOIjG46WVZbKYvYW
LEnc/Z+PnJPficpEm/SsAOddhXWEt1n7UYLgcWegeX9MI+qq4qP2vI3WdeHzkZ/I9uyNvko3HZhN
xUVIxn2E7tkVwO/qv9N+LxyJut9g+M0BlrE5gmgjySuF2JjeuzCPwRIjplkdz/qraLE2jRkTLdeC
6l/ONgBNa/lWekVGCMCIj+fr//z3LUllk673biceBKURapAx11fdnOv9RjhFz0CHbhBrH/kBpnmi
UA/xrshwYq2RiVrRhSOLl+KMO8+OhmqqGhpnln5paOjumbaLY/q318R8sR/ooAR2XqIziqDMuz5/
kWVifCXTx+gphUbU4kWjUFX6TtLsesykvNdb34v/092Lc3HQMtaLbzgJF2JjHGVG/LyZJjhkIB4l
ZJLsJS3K6i3GXl7Z4mLMVwVoM8h0NPNdCQckmTM7r6Eb5pOF2eyJ47xxkUlYJmG+DcgfIK9a+kXX
QjWaxZvZZztQUHp8TOgePOvSDg1ckJUocWsFJMIpA6Wz7k73Kj1cRHTDT5FoBMhLGqmtk/iGqSx8
Xwer/4bfn9RSHjZE4LM4Cd1AZPCkxcxAJzgL39uBiKYc3djexHYzh8POvss7RofKQZgTnkZUjOsL
3jbJ8LwLWoZUgZYUlOJ6deHC0xqYjfm/pgcN22UVM199KKrTa2hoSA3dppgPCPMovMUFaSQFdhPP
EyeD/sCZltlxBrZDoYh65hIbOaIu1JTLXcMwfCtSOMCs5PJ2FCMmHcOMspIbawvCrdC1h8Q7kWj1
xJeK19nC3K+319WfGgcTOtG8251NV8uAx26+haYe7uENCl9ITq+bYi39UXO78h8X80fpBF9okNuG
Tj4GB9fGvjDjfjyvLljHCu/X/IHRh2PQJNpzgdAvHwsz3k4P/YhAy520RE6NXrLzroarOhd5mAp0
WVWHSaZV+CPi2jSkmdMOPVqKxUF+KxenWoQb0gXVS4R8TY9uO4LM9/AJW6kMvwU/BaAkIw6xzdtT
mCVRQ1MXyShirQbJW/Q+HAnqs7iR3/mPXKUt8S++YQQ3RDVHUu7qVFS6J3oNoJGghKJ6aYvJj1/m
DYhlXMt9JqTBY6UjSnpk4kxu+q0Cvdg4KEoIJ5SqRpdtYYFp3Bp8x5RwtJj6WR8AnYJ0evtgUJTO
49Jjo1bNQjHaCtSYVTievgNb/b3KnNVa5O1tbTtotIaLQr1j7RvIm5v2AFNnSgJhFrMsp4Wf+29/
GJagMs5sjt/jjnMD5XTC7ro0skToEQkgij2mxgDGSy8IhrO9WwnyybJia0/FncUywphNps9hCQ3Q
c8EjG1f80wnYGWCzT6djG5MFZPhX5hOYq7m+pip/usYvgzwlP/+kz1p8+bvQ1Ra+4WtxZKcAZZUK
7MQurHaLFjPfipgB/9V3K9pBvM1fAgU0j/XLSlWipOEEzbPOGFMV6B9IQKdqEmuf/0unLOWw6zle
q13QcCB9qOiLaF3ZLjeyxzOcj9Ke/ZV8k148aLBMAjUXd/8rQkrXTWKt+iivNeS6sWOU7cp/9RM/
c83xVtyj/Ng3qUeJ2N3/jHpGCRN7p1bz+wo9042otlDDng/XwZ9wtwJ80uAVU6IuOt2sM26HGUKd
zCmSwK/W4ouNUQfUH5zzdjBUkkfdIeQRxJuTxEa7nTGSno6zRDsrgCQ0pix1t5BcbT4e+pxhw7kJ
4M4UWd0q/ojbx02X8HI3wtbMuJB6T7rN/EXh1lGS14puVZbWr3D9T4gUpWuZnX0Yf7WV4CWFZjkL
0971tKR4XMYpzMVcP+4hmGuNM0hqAJ+SD97ZEZ/wK7Fbh3NQFFzM/oE+z9VEYmyhH87q0NZ8pDMt
Uqn2hSLrmKuN1y3xRKYNkADpYZIAZDxplmCkIoieyIvpjsTuAdP0W6EYAAixd18qi0ECTElXhgku
wA1RsGKb116aB33NiT4yqB6gA0iZvOI+bLCtIiap6wErWmo1Pu3e6ToCfNOfzx2n489qEVR8mTgh
31yLjRBa1BFSx2wqvqkaXaeeV8tMYTVMHH003J2DkdUc3BCal9EdFIewTOzOaRyhD9wqlAZbmgoM
8PkUa6C9XFyoXcZLT/EDSzZ2AOMmfJ+lE6OaOP7tDaUTKe8KUSp2hnPs+EFEc8aqBrvb6Qoxtye5
ccq1Xhuy1Zf9HKOwIvaqb736ebeab1N+KzfddRL61eUY30l5XdQDOZ7igeh/wn19iR6KZ1PYsy9M
BC/O3daQLuSvbXkXa7IX1WU8Z/plJdWyfaWR8DsWdjIeWN0LTeUnOwSnXzG0FZ5gMLQonpFOAxd2
zDmBWnGzG7xZAQ6FHJm1ZdZs7Lq3MeW13YhF2ZSMo5YWBXIH05DGrDCG7irNjSKhpKB+hU6vhT7v
cE8NWcFuGutPtl3FxzsizSDkjteh1i83gpEkF6Y1BzZkUsBhnrlLElLlt1Ep0j7KNcxsQ+BTlNVD
7BwEn2W7L4bQqMo4TEpUVu7eEKB3J9cbonGHGuGpoMuc6AB2GROSBBnJvwYvDUK5enTD/hNOO8uo
JbgvWSIjGOvU2/1rHlZuf/KC2hvSSHt/y2BsDwQdYK7eDcuk3B//LKTvmS1ykXpjhxq3ozZnJASb
CfErZlQDm137S0HKNLRxYIJlzAu7x71Zsdl+nmlIPCoG6c/A0Ib6LdmYM2xo/mILJCpTyGvEcDPC
whHvyPbcCzR2B9jTMDn7CYXzqwK/ugw8lsEmS3sxnV4zXIujN4ndVRZiL8dc9fRy0+D8/+X2EYnf
smmZyAXpn1LdJBTdLsLfX8FgUHFAq7O4NrY5yuEDGRPrlw/H/iFJiEURqgoS5CLWU61j8gSfLOtQ
SWlHr9dXlxmd8taBfb2LY2FNcJ3OzLpaUPrqfUd0ruobRQfkhQUDeYWAkhZI455wyOfTm7RC6SJS
Qvomv0knBllXXxT7OUXIrvw5CSfcdYOlqosXQNE/BWHFqOA3AScPYUDbRcMyrru5aWqozaFjlxxE
ip0I4xtZ9FgaUI6Mm0yOow+oqElM2z5zw4TwiTpr1cyQnljwpxWikA2ZOLQkyB9yPT/t5OZYy+oO
Eq9s1UWHLKNm44hfxYp5Zn74d+Hkjt4+EMtcJ5KgSvoNjxe2nQzrsTmFWeUOTIA629mm1A+uWesB
OBnmTvclSKwhQ5YHpX1ZjizSee192jQ/lA1p2roqxFqO9zpo2cmkEO0NnvyhPXj0Hm6Ieym6eU/p
ZS57twwHuBi4BmJFyT9lmgqPr67JetkRMc6ar6kRSuRcPtZQH7joZ0+lD2WPY2TH99A/P43lqO4z
hj4aT+MOHxLpK/hDNKqWzXmer5BZpfHriyZ70h0G3YRR0Fig6e7Oa2js4cZjugbxtuDq+JNWLib0
THtndA5PgcrdkzvjlSz/c0/oTwYUZFMagoDg9LrXDQuutL9CvDAyjyVVaVXGlHXJRA/OY+TFr46Z
VQRl+5o2yI26QsIpCEavzwLziEtK8UWkwY74kfgYioveLW05nV6lVEbH/aiyQGAFIV8/BUKTIAmd
1on0t2zX24a/n4rn3gqKcK5fvmuOTEW5IKwBUJLZ8nJRfuVBUU5O6DtjcT0S96tYeuuRwwLC6FNf
ano+darfHdGJBJYUtPlHE9fFMvU443KKr00rWtkjB+wjINgxvsaLSwi1xZ9E00OTDRKyGhZ5xnOz
TgFrOzyR8V7KqOiqbJcp/17qDC2GLvtV3TKqwfD0AQAUyt9h17Qt/c5nIorXzWWrV8Z2Rk+VLYi4
TM59xb9OIdM6rv9StGSSOY/QWfNJrPPUwAco+lJduo1s2hoWRkkWSOSojdFUGwmk1vY7w/KfDBmv
Hl9pEHJRaPqtXd1T3mh5MxRmcmV1UkBUn7y05V8dfUAjGzoi5WyXsnBPyeaWKb7nH2NNlTJmBFs+
KcIYq8q3/3htvCxPVCv0e2639cwf+yIRigemOt924dYWBmOmbVxP3obeB7A7CnmRjSQGbo27pNEa
OHF3SqgAYwzpt/uQHZXEtZwrOuhceE4fUbW2DlAzCGUtqlwtU1SmDfaTil3laSW2vJF6lX+ZJoob
+TwYfql60fR96dHef/z/IsAL645zOd1ftVXx5rhNqMmuiXkPl9wQLMK5QWmGSZ1h9iIP73dVCm+S
xKEvwjpIIIuyNWLbKKcl7hSi22hPdWq5MBuQyOywSsqHHJbJGQNhoR08GjxHGQ5J8YnDpBXZrhoX
t2YDwtdJd5A8Iiv5KiJP/QS8PYEsSamYgG5djcd28tNEOVtAwEeWfPUG01Ag0NoMfyVzmItQNFPN
YfPvD6gJKsLM6a8NnqqHFXWRSQuHLqO2RX9B3gEIxUsQuR38cyHS9YV8cG5k2fXS7UVKnj2BzObe
X0+GhYpHnWQ6lAmtXaIeWr6q4r7X+Wy1d2991B3+LHafgN8EfVJPdpOx4JTQLrOIL0lYHUQ2zQRX
gcden5Ju+EW3VwWUadFsbcZhYfgVpL0rfDRAymzfxsryrtTogimbmfGNNoJeMSlGel0Np/F5SQa/
tnyrFPbnfvWSefkiqtS9aj3tzaiFJR1H75g3KxbAQZ/AuEc7pBBRWzez8/HJ8ytrrQiS4KMAyCBo
3x6zqmvxoNSddUYzCYczxZun+2vneGR+dp1HGkJTlqlnZrKxnr/qyKyud08Rr7BnNab7e/7yH64m
+Q/aiGbAbukjmzwhBXn0H7hmSlovp0OebFImMrqmnFe2d5LPCioe8H8mERsjYFOGyEwNgHFPDywY
epWEPps2hjd4flsuYeM0rnpwijc300mF9xkH3+iKusRfBvpotFPRbRQzg3EJknTq9CLSC3Pazipy
lewt5QokPWrWHK82YaR0RiVv6EU2qgcXeiJ3s9aSy4NDk/1DWShztkabgDMbiKNKmNG6FfaJcRcv
qntdatbI6PtRImdSsu5x7cV5bmUHbZdB/ruj4HFv9Xgxc/7wqAwzifOV/j2jVW3DGPQiwDausGQe
ebLxk1zLMI/DCrNCBPT0UeFptgWepnQMR2MIgkVTPy9xSzI1sTU/klkUATtr39iwXfie1wXaCjrD
v1B6O4/7SoHVvg37y0dn8D1r/7MLGDrZC0Ka9D03vFAu0mleFpDz9wla5ZwuMRZAgqBEdcrRQcOX
DiYE4tNBwf1RU0ziL4QvngTfaYFg+lAb6I+kGY4Vd/r79rxyJ0oWoV6wVO16hFKzVGvG8YCrQskQ
gdhFkyN78W04UsQ/SXNWp5LvXbwmQeqCVORPKKXh+bu5LkRDUVvgFiSSAo7UmVUq2W7sM8K44+32
/h04rgncPICRK0LB5IzYTGY4zeznoib0JBnw+d05VDgOvQlIQFaJMAMiK2aFFe7hx3K1ebBlWcJU
eUeEhKokaQ7TpipfTBp5SX3P0YcoEtCe7sthc1yW/uNPXfarLecPLXSdM9Lg05mSTkg8EL90YlMZ
mN0PyeRj5as7FQIx5vJQLSyqKcrfF/oQWRjHWoIYFZCsvGRjrBJG++97Qji31EgbojeJYIf3gmZ9
HeeAA62mfGoD5jnZ4ztvfJbz7SK6r3eqi6wmGF7CKqOW4ExKdZBQe7XJBU5Md2c3PYTz4qhjha//
SdBN1DS/xxU7OiZI1AR27bP6ZKAvrTYiCmFo3nkW/8xzqlG5vBL1rgeGToetOkBVmKjoAAtWc6kz
240RB0378uIo6bitUDmfICbxn2sTDFFTBrayIOIKE417OQkIFomoMyV1xRkxlM0tXb29ileTMUvC
7enqhlFdVAnArHw6dlN5qKucG7cXS9OLWU3aljOC8rCHiOG/fCZ8/rAWk41OSam4hcmOv+mdft8S
sCHBzuNbFKxPOUy92YR1uDNd08mTeXxRHd/hlx8BEeqok0W+diWzCnCUvLCJRjDgHIO463FPRcab
PEIiHJ371HV1x4I+KPsh90VqwTslJWz6MAQXTHQ+RbFbo6gGrVUaIANREVgSEVfx08AGn/NNGH0a
XXqaRYfvMhJu99HQuZ/MTMFHLZWQF8l17qEoJo2/WjQW4NcoX5ulsLomEcsIw7Gm6gqFCJxEc7YR
eAGBftSgOzednosKwmyCOQLnKO7MfDUXlA8ghYGR4Vd1xNIkYD68oQ+eZB1ecDoKs73/o8ebjYYR
m7Kgz5qSyN+B4XzKK3VT9/ilLHItXOg1NDCXHF+NOQ9ikcE9kh3ucHZ+t4khAmaIxLru5E/bn668
gOj3ytc/PWT8BHRg66eNIVtW8Hef98U0kaaKZD7eiPU6djEmmyU/DIy30CzSN8r+p/V9Xk67lCRD
IeM6hfajTulbRawmaVnGK4kFFQf3c7FhPsvovo4o80jXRNdDyEjCdj7r87vGySvP59Apwzl/1KPd
S9KecYr0azeNVFnTgX5E80A+gJN4W+P6TNtq7Ew4ZSqU20nu8Qyr1geYL3VrHPbELqKuCT/bH9W5
cN5Ln4QyFXEjhajrErt9I1d5jQvZd+wJllfpI8Xa6cCp+9+4HAUeOJ2zEtvvvRrLQ9bEKkDziQVo
eMTTo8d8GI3PNRbleVqygBKbB/wZzT72h8xT/kqiiwWs0BAZU8SXdSDSMeik3xA/NV4WdWGj58qQ
4ROuAsedgn8IJfyHVDpq7fLMF/k9kQivMg5ZmJ72Tm2lkvFg/4MAJkefF37/da+OeFJx2HErxc9h
PL78bvvOFias4fZWiIDflcZGaB/3SUSXUSHkcVFRLroqmjRyj25IoJFkqZt1+qWMbKE+eMfczphy
ZSfUCCKmnd4H62vsASPzNxVaT4/vFwwsXtfiTOoZ869nPWPBRKSE6JGEwJiJd6mexQOVpUSKmrGE
qmhJB0Bha0A9Kc14QHZY4W30nrh7EnxxHsZPvnVIBa3ORkK8qotW3hroDGvC3t9jG+wrKl04IQIz
ci4My2mso//Ylwm5CwQyYsRJarZ+6lKI7QSfMzh7VnPeHbzbS7c6tdmWlr/trWi9qhBwloTA0Tck
jeOB4499+vo0abQnGJEtX99OJe+2HfZdMcIMj63hET4UYSd/p8yTUEPESIBpoEl8+pf6uw2r5Fs+
MRVZ90RSMe9vQKVMxrZgYXAlBGJfKPcSqgg092a3r2aWZfRduAfaMMnCaw6J0QuGoP/4gSf4fs8f
8kYzzAcw0hvvD8JMDdffd0U28xMPSUy2HjVb0/xOz7NUVhLY6oO1Qez+fRExQgVbJJkmHmWpi/VG
y2ku1ew1TI6JIcU3oceD/k2IqWfzYh8Gjz9pSwmbly4e//5xS/h/VAlPQe4UsCTnkxitA1Z2P8Ze
XNVkRVU1gs0wwsR1eGuzofdOQLreZ2Bh/MqQGr9XqsR8RvQPCodimcakGYjxtPeU1lAK4xEKt0Yg
L74G5an1UNkpbcHuMyBDTx7zUFASCwDFqmgeaaLUI3b4O0izX/bmPrkwctJTaR6fCv0GILKZD/fK
TLgkD+JGis/N8TtgecP4VBTcRGjJ8rUwm8pB1ByR9Uu+SMjUQarj1NWgYBNzd+SGIQrF9dZNCUKT
oKen28GUKYZbBpAR472amJSe50bEFLi3kjxCrZuEhcsJMTO0aC7Nly2G6SIV2BVH/WLy0l6i1UgI
rNbX0XSWYqzFNh++vIuFLA9927g/8z3AFlMsV2sfcXtK6bJ6Oi2n/xMohScsufICdSuKDCcApr45
t/46PEyOURqPpRAZlzUwrnQvTozGjnH6QLbFj+QtMyi5Gr8X7g0r1kU0V5EitH0ajkU9RTffUCuW
Voe6uRbUvBguZPiJvzX8l4hGDp9LoKqQgXk8qJm7EMA9S1cYNa900QH3sDe3kEIcfjU5GX0zJvDk
nPTtPs+Khg5uO1H/OfWsmW6xwzQvrUAS5kkHNeqsbkWiJYlJd//5wEcyG8nt9iJ69v9M3J8eWq9e
NUyMsU5W68gVb/xIvNxVd70+a1rhHWpQD6dGK9dDRKPZHpGpkaW/Xjg7UiG9UMS6HJe9ESTGCFLe
Ih1xBzfOrcdUsdaWvOb7DY442f7Rooctdib+huvcVPpYIlk/4TP/UzKiyzJPNJRdeKW54U8GxlRI
HXD3ddrOx3iPfv+INmk2YO7hRyYtWbMEUg0zLaJRrMTuyoFlYGDu4uy0pGdLOzWQmPoEShcauPID
dQEYSpwcE3fkx8Cf0U83D5GHfxog36IlAeX1f9XjwLvndf5WCuYjCvBBMVXHLSyWqVbzB7Q4mCkx
YFOJHucJktOnqXzYha/h3VlSwujHycPDf1aQSHgKPfFLxIfULG8gb2yMy7Yo3/1hsQGmCuuVia1G
yn5EUScYJonZP8EFjCoV8VBYTfABGntrCLwiBPWv7ZYdszaDTuAjd4NZ0SQblyZeqk30fnWCGTD4
aw1lCN9OWtlCTvS2trGK1WGlVFq4UFENG27M2V1QCywB+Eb2ENi9SSDdLVXv7lfN7IporCXII9yO
LYex4zsTWULXY8LgREwN1mK7gNVA3DZAwvGhdDk03Btx8dQ8vqFkVxsea9xIgx73e9e9tmiCYrin
5mOFRyldXANpTetVpqcKI0WrX0cYHph1cHtuljKNo3o0UmelxiIXsSOhTfibKmOe48HtD686VZJ9
20C9H5duQbqOfaiymSdxgNeE9nRuXbJuYdQLbCmftLKveuY+4G7YO3S/rbP4T/PMBqdomxAc9nRh
EPL3fvDnpGjBZyifLvxuiPSIJ4l6F3kIQMn0eAhFGsXGT7C0zuZ54MYzu5GzLcr3wQAQjQ3aWmCM
2SgwrBpnpacj4q12hSe8AaNN2T+fFZlod4NKjpZH9CgnISGgD7XvRJc2iDYzjPaluhPRJdNhmnFg
r/NHLkwv7KHaqDt7u3L3Vg1PPeINnUhDedqwBDGja8ds4tx7j5oRuJqjXdVKVudHyYd5qF//GRVi
LUZlqRbM63w8m3S7RobCB7zjWb6Y7KFVsOLQ8ZjW4NnaO8BqtiNYymLXONg6TW9ydJMxCU+Ft5NK
CHjWlK4ckgXHb9SSbJ2dn1CffUgJfv9QmjogQhfoyiyDBPRJsemeBgKsqQd1UkVsJw1GhNgrcHwB
TJUWG1+9O0isAQ3rBQxqIUbPuA6zNKZQZkEZqFhwvVwHAFJj0+7Wko9IQxciIjmALxIx05glBpJ+
kEaV715eX6sH6gnaPfGw7ze5oQjRwqLwroghT1ATWdPEVuuYQ5PZ+27pRTlFV+6n+z/PCvedilIE
h13PYjvQ9S3YgOJAKHphb06B3+I71HqU0MCe0CYi3AwN37sOk2GnxtTowyRNubxKZj+xGsOzTNeD
wSEc/j4WIWhHVMyMp/HCychkNKW8df4iU+u8RFbXG6945Usl8O+xsc8DfvrIZb2160SMCL5zPVTj
Ca9u+jV0pctVhz8DHo7tz6AVNr38CF/Xs2LuBRhBMiHRWoVdsA3iau2S+V/SOUrz8BQ4jofKcpR5
o/RVfNTGeHiUHf016JCcsFPlRognYdf0DKwRkLbYMD+evKZof18u7dWhATUKUauqSowkUU3psyjU
6tlyCXa4ot//4MtftOzs3CY6jM51J1M/E6/PmiSq4Ti8u3KO7V2zmV1608TJRIlDiPbRXupsTUtl
LPF4qm2+z8oddFj8zA40IcO6Z6uT1PicpweQxRj9Eogj4MoKMhb0RVTn4fF135A5TLA4wfT3RUUr
FV2upeqbcHW7u9894wtcb8AV+5dm2tZb5vjPZppmcuNww/+BG2F6ZUlORJ2gkNuBJqGP5w37d578
0MATAL9gHOwXGPra0d5wrPmb9QvrRYi3tp5AG4SLYvg/2VNjnefx1zldMhAtcjWwlFZrMc/24/0f
QNxR1laS1mT3XKyQsA91qSsyGmxg48UQDEsIBxMokreb9FqgvLGYfG32hntptmsENe5ODDuwPaCV
dqs+v+jZZNtlTtto2P8Y/SPLVQrupBmJzQFOHMyCFLlKS4fUD2mmNC0GAkSKpixiAgQxhRqOv+zV
oVU0e1fj+FTNIDB7kgPv92u+f4tfdEWv6WWilri4kbB6VtM/3s3ncMMtwJEsfQqKJ3egk+18Mc8I
i4yJvvv2nsIFZNtp2pK6JogCagVSMmauP9V0XOdDRnScZApdAgj9Y+RYcT3MPijVPYLY57ExWqEI
SBBs2QIRo3bNu5pX9GKi4+DeeGRpTQA8qyZHJThlqss5zxeuUinwSMtYdWXSXIrjjnxXmIvkH740
VZboCOvxwb46sjzZgLOJ7ZSQSrY8a5jzUgdxyHza6R2hBQ4vCkei0QQp3tS8KG3Wi43/dBaat1W/
xzLTjE2lYzIQFMK2/Wz7NtqdTFUS7kfkvdqM9IOe6FXLg31npFzwCrwv53DqhCIllMia5muhuw9X
Eg5t91qqLHEs/jvHi70Kp/ueoW5AKFpXlNIF5DYSu55JM0qMzzQauTGHfx7hrmnkMr6rOxhvLOmT
7md4LErRQqk0JoWmIYKaoiBZXqh2JKhciKRb0r98D85e1VohXo+i3UggreWXqCZGyDEXJ/BpcOsF
W31CZGmtI18cVkeAX2XYYdxZ1E6gn38BIh5ts3oHf0XsYt4xL/z/rx9hvXn99ylH3GXUh22UAlzF
El8IweIhm2VlOmU95kbwKoHMkdE0u8EWQbcl2vQL0LQwsx2l3hVP/JrntXB0s+rj9ZpCVwoGa3BW
EBbzbB2SV9Jpg4bQafGZIfdYQadwqzaI3OumBLAM9HanPi13LMlfo9A/+wAabxBiG58omuiJ1jsx
GW4PU3sTdjm2ejrdJuLweI+heZa4ObZv44VR74MiGjt83x/cD6ax3jzI4EsHJ+ZYWA5a3JOoFgle
bG0w6AuBUydrWFLGXY3Fe31d8dFzcDh+Dpt30d+eRjkgBeLngNc/sgByCYGXo1PxopK0yF/3ob4c
tmvdgCu9zmBoVqlDNLIig/ljgCXrfdo261pK5tDiWXEgQs8CMgf9z+NJF6Ej7oNi9f8ZwyH0RJMa
u2Vg6+P7VALS2x8s1Xt0Wnr6xnDNM4EZHIbS2966Fd25E+5veuLYmBoyEUzmHZkzPW0UqIRyo5Dn
2+9aZXkjLD+Rg5UgW7wKtWfLXNTGkQkLQhGOBd3Db3l1knU1p1fns/Z1w8YaYMxpU/KVG2jLZjNG
VPceRAA8/fkvDC/UV+fP6nB6kBtRyc6X1CjcwxHiy7iuIDekxfIUi8KJ3QbzNdiMYCmvdXwIrn+j
143HmFOdoPRRmeKBq6vJ7VTCaLoOQDWDw/QWDGYF+BVzKXBhSt0SX8TGrzURRvWJeocxDNe3T5ql
DLIDuW4Idzg3f0PNVgoSkGLyNEmiVHi1524ltVZecefF/Hz+GFwuFJ+tYjha7o59OG9AXv2Al0Sa
7BeKkVbP0vthPZtIR0iei/VGT9NWrVIA4xP0+mDKGUpqfGpmk6z/Gswoo3szytu4Ip1ltt+AzES3
DnZR0L7nN3qGtMJtq/gJfmCXOEaOZImS9JcN0QMR+LkN1k/3VDCKrDsOQQRqT4pAwRb/JsogBJ4L
5GAwDzZhVRZyqwS3Eg4aT92o869zfkddiuMGG0sbwBdC9dNqtMSWcQYDMkBB8W5Fi5wTzxLcgMY7
YhTB3CdVUJYjoBtJHYKAqYXud9zbGW6ODRqfOaDhiOkmIs3MZtia9slp8j62lQMdb+0SgSbrP1jm
urQZBMJE/hszVlmVclLHdife5FGL3geBi2GACNJR3PqyT12h8RBWU9ZZQmxnekxempUMLNPW+9X9
RR4M61YZr7EQt8A5MD/kiyoeY+WwWm1ZpO8tpWEbJvFPPrf5eEu5MmynRWR3shgnYicIsPIXWFum
IHPDw0Cw79kQ701U1I8ina3TGw42Jp2X5kKeTfh3e4PQfkpEfegXuC7x6eHzNW/FOrSMXG2EiqRg
L+y7jmyMVIXsNCQcShHO/5RG6nn0mSH0KBG+O+FhnQPPr0W7Rl1x4uSAmeVvVtZW7lA5i3b5ajd3
AhKSHuDBfsB2xJfL2sIOag/To0ZgqXCGMSmwdG57mLzLtktIWDwgrshI9hMD486V92yK0RMUOtoc
4o8cawEgkgCIcfJ/2I+Eamx7+lleaB8HwnS9S6Fn79YD4Mk67HrewSmI+nCgGzW7aibZu4wniJOl
ljW8PbaLQNO5XeW5M1mlzCMHW7tD+2xS9YaO/rcCyaR6puBgpwAwJ5u2i9VXDxvPLPeDiJnMEOcq
FTHOY9U5Xlgi4XOkIA0SfMWGg7KVQ+lGzbhjL/76b3nCoKhfz6tK2ywlL3JDyLJClOdXyr9m0Amc
QPEXsp3yFqP4v12hFyz48XXJlNGo9HRSUpX4HrCXjjfd1uWjowWiaoYy3b/BEyiWpYDJi5ixVP8F
OWySC3YRY1KUercc/tDYZKYjX7Ep8sN8JU+GexFrozbMbyUyrL73bC42IR5TXpWlFFHXk0iaw1j0
KAxJVSAC+pWGWseuOx+GXJv5nYniKAIasQzhM7WhTiHiAbN+CRq1Icd9zZS/aoINPy7yjDmyQmQ7
dRhsXe3htISKsMQrm14epcxKvlMj5p+k2+wr2LOwCMrraF9llTyqfWCWkWl4YyQyVS8QiV0NOfuO
kcGOT50ldCUXz21z0WwSiyZngCQsBvgeyhlSasSaoBEDyYag7nNh2OQ46p+3e5iF4xOm30wvyiSH
qNm0hRFTJ4Rcq8bIFNcxuEVNr5aoRqYNuFGg7TMPmdj43yNtDMR3lb0KiNM1+NAH5bz48tL02L7U
XufrtEaT+GgG+zfcwV07z2wKZo9DSURvkUdd2nZhQii/LtNzVRhpl1MEH8bnDvvOAem+ZjeH61tj
gI++/Oxj9BPNaDNaZFO7pqVx2wM+3Sk+V7csdwspcRIuF/yqe3fATpu74XyJDb5QAsiay8t6bc1R
ySXWwC3n4XAwZhC9rePGVQ8ecPk2TVVTSb3g+msIR144KabcJ6aqdjzYP8SH6QM/MK/qdRYpBqVK
eaQ9JBFprekMIrRaUcSZTZ4+aZe915071xcdlmOocb4V8zzArjX+D1tzZwjRa6FAxcZ/MHNfSRBj
ovfk2lGIM51wP7Ra6WAVNhqbNR+K6zbbdD9Rdif52+xRQ+67wa8MXHBT3Io+K957+x78Xt3P7MIB
HibVzLtqFuae7KWQrKR8IR3pPRsambjzb/i6DtUqLhH/WMixS/MBCiMlqecGFZX4w5bN9XKuXget
FYiIwteHntkLN1PfIMoYqQvCIi9YEmOHwALtEXMYXEiLaSCgZ88ez3Ta+8s98dCi5UeLeGlzG8vw
Xn7lFhJT0bgdv7KGK1higonZBYtAkhNaiaPbuXCgcCXgFK4XAWaZKf7v49lkkkYhCjARIEEW0h9M
Lba7V0taqRveN59sQCKesHDQjHHXVHjrnf1Xgn/Sl3nWUMynNrNpFOIEl29y5pLJPsoFTy/cTx9U
uP1yYYTIXZgWTJjH+fFdu5qba4D4HuobLbXhDqrKm4LvsmHc6PetaK/k31x2qQwsyCCKU1PBKf6L
YwTAwPdg688cAJmYwXRIWd3PyaHQi+JUNpTpFbtAooP09qdUCGuXe+YxivfuVkLZZX2CbVl9eKBk
N1tfZSUxzgs3vyS1HH5UI93tqJTQVQEHJtSAzEpDFagHdPkxYVKky6sx7zMOlS/ebzKvJKNfJvL4
0apruQyjFoD7lxDCKPP8VEQ7PRo8kR2xtD7l1ht2X5JEM09LJyoGEiyF9/omcXUBG7d5PhxvBhxR
vlbHeQgiThbPkCKzSoN59kUVK2eDElJBTVi84iadRKW/g5hCMZemXZGSffyUgxMQEQ+Tgc+hLNm8
VO9shJgKewoiBcRNpr8WSrbloQup/1yjZTZ7hDQiYFrlaU/FbNlpM+iQ79vRkRDXaWx1LV7lTWo7
jjz6+yQSzTzb4Bgj0xCJ07/MDS6OFWmQFNC/xxAPFjpTwMbFGEFBFO9MlL74JJt4FbWLHTwrsLe4
JdfRK68tEyGSAu7ELwzY6WU27PAwt3d10WgYuSBoLdKNyJZljD5/SYy437IAlxxl3xAbZ40zlcjr
y36GuuDqJ9CCnQdZPe4MeZ+Wd0tXTuG28sXvN1BfWWnyoER67P+LNud/Rt0KVwe8fsmeAAvCk6JI
eVs5C4B1elyXoWpnLquSSwlpzfCGwB7L2sISYDNVBTm3JD7Z+wO8SviKARkDM22BNXgLKTgIkW3z
33yk9uW8iLMk8nQrr4BMcUzDCFFE3UuVazFpMdpFq6dWymMbuj8rha6CirWKM2Pp5zJ2jIxwkBZw
a1L73vEY1SBKuVroqUugDZXQsjrakadP/ByOVkYeACl9ufS4JXfrX3BvwCTZLpzVS9xEmzydV53V
4PPKBY7kgHZck5BwHel8DIUDN9bWScK9X7kMNra2krsa/dLLcAlmKKqSza8WRZS0xKkehnULy+5j
2clarpk9ewgTVJ+HPyKHg6959PK2/Wjvv9Y16NTQEKGZqBsp8Ml7ogUhN4YTz5uTIas1cmR6B/co
TMSryM1Ojks4Opl4kD5ANZxZNC/eLTcxWHHkOxUaAQ6q3AGYNVd9nAHeZQUXM6elSOgsSm0wPtSt
2U119WfQFuSKBHH7NR8mwcSuIvlUK7KM5eYlG65m3AgZYSREQEAujRzkpN+FvXQ+AGO4U/7izF0d
37uPByrS18hbzVhSfpPgEXQdOG6sTuCmNmovVIP2BMeIBDMLqWojZDtRzV4eH+XxfppXte0tjIn8
8FJVu0/fh7lyzou9jTicrFdrsUDPeS6Tit0XDpZ1uhrFaa7w9HvwNmja69prS8r6/TNorogwekh+
7JtaE9XtqpNFWWszz/wdg1UIEZuPdiF6EQGYOHoD197re2koV+vBlAEpRxQfkb42WEEzGAoYMP2V
J+zRu0QrwBecEIBQ7ZkqzBxHpU+Z+GpR++Qp4YJwIYVFczS792linsUduu8Ia2N25JP5yvW/8opz
jhZ2r6jGrLaRuNQBPR5RusEnpQpg00S8qIoI5cRt0Si3B3vm1aBG4ID7xEp52EzHqXOdMjax1kDS
scVF/hAsf3WVHW6lQuB08V1MJcUGl3OLajMoxVICmQwod1LPduIbFPXezIKWV2Stw8R600/rbDgi
bdafuhs4bqVAk5jN9OAtqEwGSD0hhIZv/N6fNiyFKm/FviqiS8nGHVlr4e7FFtor2D132HLyTzcg
YMHk+Wa8A0ndM19yM5sNxdfF3ev801BINKEkYjdcTJQndmX5S7FwHDYLjkWitx1Pb4rlWupUl1WE
hogpS6O+t+7j1ncD5EePVqyn10NL4wQcjRIAoefKvTNjzsRk18Ws6dc8HxXErpJXz4PYH09D7F7n
LIm+zUiM47kKbh7J0/hlL2m4jVbnR6VGbbt5dRRiyrN+Ao/hhw+X+EKS7mzg26MSNUlldHAzeE/H
vfXSnermEw9KJ6Bz9dlCu25+3MS8OoCKzLrdtp6b59sUppCPcK94kATPfKD+zgJzAflgNnNEoH97
6O95NG7/nFto1O3De/88KcE1hcMMiW0U6jchI7e1zlTqASy3A4uEPnLdWdgBqQAdhTac/rZI5Acv
TjQrZiXeur3RE3iJElKu9zMiKyTPnlD4FEeBEC/xT9nbLYVB0Z1AOEpfhXlyBrgGmACQ0AWeGjbg
73jOIAsJFZTx9cPlwFKZbAbWjVmYjf+WLdY7CPO2DyFOXRNlzaiPeZTJPrbSNIpE8Jb+gpcHEVT+
l55fhcH3tEpA6um6laOM6k2QQ0QQwUgNCmlOH1Uq98Dc3NDzomM1n8txkD+wKIg5Qj+Vgm+Etr05
gm3L9Ob6SRP8JUI3UQWxyWUEHwKt4o5cALAqW76gODCC3auzbIpgBkUgef16WgSlRfm5OQDleBS1
oB3O5nqv3zqTXZ+OoSmHY/T8jyUITr2PiCEd/p1ycuMOEa4prVxuFN8OJSk7q1o6VKxw8EEYUwQG
fG2FBE+XhL8cREttVIWFU1bgbHr7Hpb9t2baibVejBDn2srB5YIb8KCviXqoajvPEA5UXvdqzQLY
4/qEk2sG1pqJ5SABZ86FSEDL1shUXZZySNUxLLy3iF7cLWOIG4+WwiiG5/E9ANpQdy1OCmDbN211
F2/MwxODirNZWRPcNPYg73cK+eV/p/aYa9Doxio92rc1ODW1tBQY0QKoJN6KERwL8qHNz7lEYC4V
x3+EkauRvPyeZtKRDegtsmvl4JPKAN6F0BTF4pTeetOi8m/KbZ9M3r20gdH8FqVyN31UvVuM7ZPs
nP/9knQ8dkAuoU7n13Qxkg4qyPHj2rRU29tyWHUsz2ZjwVM7HwrMel6oa5fZGLbYshbf6+M2JqWe
/8JaVpxID2EC7d2hxy00F5zoUCu61CMiB+WK9SBCUjwxWu9pcbgYqrRdGD7+YHlaklCl1GHcSc+l
mCmDOPSn3DlVjaHi5ZBs27KdW7VETzRJOQAt1J5Fl5HjowOzhdXmnHFm5OYHn4UKkh52LDwYxTyB
r7esAWW16TlCpGCifJ+uRqjIp6efBzK4oJ/Nlp85jjBlH9d8bhS9mgUU3GtjwEsMrxxxqG84byC2
4BV54+uaUcg4wI5QOGh0/mTzvfcpHj4aSGSRELsK4sCeD+T/yUdkSf0jOMbCpwzAnqs/F4YNcAZJ
J8Am/9OhZZ9KjklskjM6ts4gg1e7bydmYTbJ1BgzQjdU9ixJENyvDgjxaPnxkQNttE8XOQlCi4Xs
b8dy3gUvD/QsE74RSyM5viC1O3prn+nu1COBBrfkUxt2lKAWQlBGTL5sfYLHxCkn+wxEbJmgjAkK
rhJ68Hl844ufZASJkV2gyPA/CRVOXyXs5si2vxWrSnoJMw4LHlgQGBGlXSgJqMLIia/3xhZUPOYS
nUHST4wcA0aiSjlVdbcbmrunbsxHKYgXgD5vmZX2ZTVVuE4q/DWVkMSrxX9kRWbUQxitlTIZ5kX4
0jXI9kO2Jb4Ea+nD6haxGG5R4uVmXCdVpZJB5yWpJSG7nzKd5KNy7pzt97tXPqTFRu7uGC5fns3r
RTFvobVdrh1Tx5VjqRtvIkKwo83/JOPngRIdpiPA1ebHiCjv5qy5lmWaylWseKJfwg39F1cv355k
QoLQnUhq86Lx5M2YNAV5/+H4mK1N9qTOE0Atj3inkaCVRLiTW4wGSI3eOoobXkG9+5V8GX0NT/rP
zrBfqWGSjL0RWIDHCnvrf96ktpXeweSDaEc8i0TFzKL404Lbyv9xom/kBvn0YkOgRBcFwzwc+ARf
HbL2IiP6UoZyFKyCXOB8c/plzfJXT1FvMGB9vA451MwT0fNxQ8uQfAwbcnaYm56Ee9J2GjCjrRId
k1HU6UOWGr7HVXgzODp+uybACKdUHKoL/PkJSNUerDEvT9GBJqp8EwY8JWSNvE20/GV5K6XUwj3r
1r2w7XAvJYmRyJC2qfNPaAuQ80zwebBFFQ2gKdtF6skgHeI3zze1/NvflEd1arRNa6ZeaHHaGgOb
tfZYKNTwbi0kdJY2EeJ2Pxu6YH7867Ib9dUEhbGAVjeIiCVdEfw4+FYQP6hJtcZ73sYJllkA+Ov6
7847TKbMGtiBij2rQ8QEFETl1r/ZD1G43eFDp9TGzh7qHtk2Ius/rpIFTMz2I0bFIJNZEQJnTKSZ
ICphFNs4p1Fc+YBbStbqAGjFR+areWKDDkuM7OOf6IvvhhoRSH3fBF58OiaDB3CWaDszh+VwZ4Z1
tAb2rFY7yAZSr5qsl4FJEfhziNFmGUYTBnQs5pfliNLZqxt38IgdDm5j7CcEbauvZBJ67aCgQZIt
gUctBuNGfIh12Jr1yxNKckTVwj2GCviS+wC2Nwq4xnXhNuBXFrCRXP6p6hmxXmrU1uA6liNuuxkk
VFryFQoSSRiwk8ltv53WI2s5I8tmPG8XK/q9kau6eyruwnFgk8zU+K34P13PuI/I1UMgTe7EC3l/
pdZOqflpkLjHlskU1VCTQaK9t6mK8nswSw69OxWrwvmTsET1jT5hJrlbmtuCm+4+xGhdGWjpYooq
ClQ30aic3p1A+AZ7YO7NC659ess+YWzbSyU8iuCDtjOHJtjI58nI2T3vMBH+F+/WOAdONaXsAdsi
roBEKXHASKCyLw+/8KzEbsXJiHcoTuefxQKDvsTqVGNmRHbSiH8F+uHjpCi75fiMM0CzDrXzGclK
CrPeu3usYqn710GQcNtt+MfCnYNiUxK27cEKf2OtDml/Bv9y0igTyCg5mei+sB7NwBcyRu3fVebd
Qp1unqp8U1nkKYm5oWu4KjbdvGh/n34aUPKBzX4z5ODRSgnVNIMr2E1kSCDqn8cVtyxWt4yZnub6
9+xvSqgADz4dAQ2HyAsXEu+fbgDIlhRRQVje1EfctZxYBufuxyggwiI3n62lHBeK34HogfVJ1EF1
UTfoXYSOfdmd5fuqCBTjxjkqogZrCtnHXOFtNEsdTGou8h98NTKFfUaAsMRj20QRm00xg4amAEH1
JyXu305Nyu1BLVKpmMuhNvcocKs/UOg3i/7A5fAsCXFtCzQmqTcsfV5kUNkoE5O/FPy4JyOn9sDL
WUMf5F64wdTpK7ig5Wo+jlYaSgvPBkc1hSsE4SMFo77mR7wd0kPiMzqBO3EJumBUht4zICY6y8wO
F+lRbwHxHpgk/eKpFYU3z1VHxsjYPDCqlsW6jzJxHsPbVuSlMgBm1Mz0EO5DJiNPKPDraMywU9yH
AWQDLiksS42gSvh1WlkJ2tRG01kLYXsM0P2Mxhne1YLCIHmeSVp0mSPhzvhiDNsFLFIS/pa6DeS4
v9c6SfOOc84evoxBMMwAdieUuEGwvc6O4uvKVDGwTVnpxwXh5T7pVfgqu7cWbDHBmvOCotsakMmw
DoONlcFbje1sevH9hVZ+U3ekVIbWihmJlNwr2rHul42NbqRuIueW3QbexcV0ip6scjkThXPiiaNd
LLe7KChXy8q1LMTaeQXgjIROQ0IFerqKxFBQ5D/rcJ1o+IbD2+CnY0eQNZrX5Ak9HdSmlWVjUuQ4
MqSaJqh5mNgmejXFQdyO+kytl4VvTWL021uFIMUGZvLdYmSSuJHg/w3g7EgjfS5JyY1xS3uqRAlr
Bb2eAaBVLZGsUmaBsTR6zjiodP1eVWsRwyJsLBhmTBy47lSxl+PLKga1S7/wFXs2la70bbbn5rlN
Cj+aV1OWFqjQh/JgUvnXUrIaPR6JuW5hw13ifISHbgXKYSxWKIVN+gVhssgFFUX0Q+stgaXNMQ6i
wszHj10s1545uTw6jpbDyijn710mmYOgw5qukSCb2S+xfsuUkPawLl0abYX0vJiLPXUVeonDhOxy
bFMWgrs5P/befv090TEoTHRrfsbwGxMrGiIo2PBzOaF6r5chOaTx72BYboUXcuxuLr3Fp78H5Ew9
VoeiYLV3IuoAN2BEjrMqlQyFqy/77qjiLCjRnuR7moXuYpOLIUv0cEV0O8RVtEL2YC+GkaRYuoQF
qzgNYzHdgrwAMDNIDMt59RuAlyZI9yTqWR6FXjxvyTMuwNa4APrSw+a+SXyH09SOnTrIHmXzvclu
mxccUIfspvVw2JEtPOUR7i6XpE4F6AQwQ2WXEfjQMtES3hRyVtq7hd2miXR0rCSrGj7PvcYACbdq
Cj/KxNvmST06/l0xKzZXA7oYfjCR3MDWQLMG5R2B8ldfgIlMbgd+p/YWWYJtqYSmoqSm5GD7aq/L
nphVnZDj+75Gl26NrU2DlXa+Mh4o0D+WwPiSDNniTWwmger1dP4QAzHgVgdjSd9OWnRR53pcHDKs
XPK6wjHbrGXE2OMyi00k2gcfhSNykwGFmOMJ3rtJVkJv5ieYZSE+oZ0pF1LgoxXccJ6miO6LhL3I
3j7yFmdERdtWydodJp7Q6GSArTHHx0ePRl8M4LvjaYOmKp/5HvdcGLESIVtQugsBB9lvNIUYTA+o
wQJPSrt71pvKzUwkpIyxtoUYCz8YZ96oMiI35ke1BV4YQnX6e6BXic67b2Ykiv/HvhPxR+64hFQ0
Zu0jIy/UbXqWRa919Eow0Xgv/UjqROPXKLN8BSyTr9EMbUKLqE/1+lWzC2KGChPDMX4QdEBR9w7W
W9mcNAR9dKrhjwNhR5D723LuEah0pCcuQrB1dKQ7NAcq/o4J9JdvTTYOf/k8dGXlmHUR4Ja+HVGv
Ywe9W4snDiVMHUpgDlw7vpoJW7mcIpZuHZnKVVdFpCZgjkytUTxYzXc0jgc3ayMiynFn3ViOd3x8
+ZAimD+9urfEW0qjQbVYhx7cj4Lpd/dfHVeBaPY6tr8scQLDfWTl99hqyF2PxBqoZ92OSi8CgDTl
CHhsT8bDDK72tKX40JIHAHQlkcJQ68LHtCrlVP3sQow3AAJtCkSLvhttZWeHPy4ORQUWRAMTcrqH
tElabrX3jxrkmyPAyJj0bJbRtcitaiERLB1OAxZ3Nea3JAvCl4fNkV0Cr6Jw4faYj5JpwERu6wG7
dEO8rhyfzZ/o/yr6Nxlj4xqCmtW8Un42cdLlcE61OTjlCRfUKgj2K48LMqHWzq9IYkE8jLMXhHR/
24SPLX4mKOXFzqUOF4NNXT2liCYdr+ECrxJ7Y5MUcF3q5BsNyWPAGdi47O0Ij7gK3UG4BOqkyGQU
LVF/fPwEdsjIz9VunJ4DNBmjgOOW+0QX8aa82HmLk2EUiLQeJrKlLFa87m2rMv5x4CIx8O7fXAUG
K5cs4HsF6Frj9O6vt1t9jXMQtJ3/T+E7qEEftPqIcPWMtHMfVrpfvud5lUrUIvvEJyuvn/4XosvQ
Rffgom47FLKg0vZTQLLmY0KZsy9xTm7GQ+3Wd+YdhaZCTSlN9VvLp3P32MmsMg9NvaTx1P95JSkR
+fAH0CxoWOY7OvrqO5XMK+zle3Q+G6YFdieLtHDGs6EB13i/KPp7Qm1k0zzpayrir0bacs3KB5jx
XdbTcwgsQxhYwHbUyreQZdPQGGOEqDHW0+da4rKmBIAJtqwJp33EIvjzWl+hKQ9VE+H4MzgwogBP
vpLWxRv6vELCDlBtCn5mO/Pe5h+ievm1z+Odn64xGqwwKIqkUsnx0itv2sf+OKq3uIDGfqNFcHyq
jjeSrUhuUMq9UCaDQ6YS+4x8ydKmLGDuOb4FVfo0YDpEryPosv1pnk3Av5peicu4PoyHyQmxKHLe
lkzPJB/haeye8qdXyZcrmAL0Ni9YyEcWbMgCFLJFWBmga7umH4wS4WySB+2YI3IZzIaNx7Siaane
VCYZbPmGAJEGbBXEZ/BHTFy9/aQ806kymAFxqJTJlG0D9wj/1dQmaEMLVff2PhC51cwCWk1QVTxU
gYCxmb6idkOSGtkp6AzgNdQQ2bJ8S+SBWkA5S2wMvaDgZ/maXxQUey2KMrijurUQ2qpCB16iGLw0
HHpnBhQuNM4dMJK6YY5YkD/X1ZuiKUjm/jL5eQVKlniWhsBEwTm3Y6O101By5K2YQ/AOt5KK1RAI
CSiiOL59e14PXVBUbj5fsLCDn03kTC7vqMQL3cD7aLVCXArgjEAVpHeSUi7rMCP+qSltHKjE0xpq
bAoEiF/Bc1XNd3B+TOhZARhNH8PqmC1kJqAvDgbJZmVt6I7s0221Bvram1hirzU2+rgPmwyKvXTp
doIExtABX0exS6wHaDZI0kgAL+flLUvJdISz5CeujdhGX0ea0JdXxXIpo1JxXiSFPqV/S3nFSeUE
2VwhRhIAE23xhvDadnJXKBRepoY24uRHJu3QS1kExeNW9JGIaZHNeUL59uwrX7GbzivuJqrVix7R
Lp0gSvRmIAbZszlwlEmFOUNcO0A5TXNhO8IhdSMVICdoZfDLryOH94CAjarU4jsfAJZc965cAt8R
TyemDLbQ/ie3zYvLHxnz4iz+U8oLC2JR8JEx30AJBeUdCHdulqqqkdUjL4NnJKxO3gdU7ES9VEzh
rCLz9pE6+XW5Vi6Un0j6HN9bTyNf9V7QXPwX6ofGC4+xJ7Ioy3D6AjuYRRA+dton15xVgdw7tRJm
GIYTAAmZ9b4HHvZV6QHdw/MBYLp7p6+pkBCut4dl6vlheYnh5jDPfTA98W5XQxEb2U5RTHOk5ih6
c8BiemHpKEVgFRLmMK7RrGKRXVuZFRcpDxjs0ZPpfiSQlJTpuEVKAnzUoPSBPUK2DYaVMFTsF3Dq
gij10eiu5Qcr69IQMImRL9QTlG0OjCCCvKFzOL8yCddZrzBlU4GzKhUPIKqyT5w2nn2DizXaJ2AR
ij2jlsdrVJYaokNc1M99EE1ZElUAvrVP6HYHadS97Sw5qpNSpAKwKVC3Uca1NhTErvblAE/K4IrV
KWHhQLB9B0dGvnR5yEUeerWQVSKcn89FUQS0qWcgwLsrNQpZ+P5FVARFUIHfMryDU0MPBWa/L0Rn
SXb5LHJgoEPNkj+FlheNuXhcUw5hegD8wr8gfpVyP2C3LVmW8ze7KUhlt8qq/0zEAz9/Djp3KbRB
aBPbfC7xQKmPv4OpTf0VMPYlDHWbxPpnjbTMG4h8YdMC5VOAGwJ/S6xkNZXAs/4BsWFgRajR/PW4
hEMz/59fU1A6ScJd//rZfiLzQr2rC30xrHZN18N1FhufK7gMpu/BW9koOc9xKpOHAxGNNdk/GbnR
60Jm3hSlVNAIvVWHwFnEpvSYkfE/b05CQfllheXIVXuwQlODO/EddgVJh27t3v220KIVL2/7qFUa
Ly/U7hohtp9FmlB2XreEScFZh0u73x5n121cBkGzN61X06IP0ynNd3osMaiA5fVS7kfSJZSd4VeD
tSunsYvRw+w77YinpP/p0DppHfRXm54iaSiYppktboyuz46dOW1OE8vCR5crauu1ok0/AsUsdXNg
9tVKYCu0yn0dkpO2byj3P8qNVqG0Vn+AQKk+/eaeIkKLyJDwJvzJOCPeUpDO3W8Fz36ccZrJkkAT
v0KbC+fAuaVpmhTSUrA7I0J6OGhM2IyAklh+6oTo4MfJKD/bahVSriK6jaHrcNrLH22mUtJ4yprr
9TXDjHYct4LUWZuin3JAu+6C9ews7W7ZMEoEOcCNg95zBQmrDMIXjZzf6o3gZxNoHlUBEE62AvwE
tQgmQNbE7lXjhboX7oVYVV0FSGsPlETA/1oJUfnjUlzi0J8Ud/CyY7ce+7rGVm6TPy7MlZgs4VIA
mIiNhGqWZ4LIBaYeo9+G8G1cXZcVvoJt9Tx1wolBdhZGD8wsFj1W/wGuYnY+ZU+QpCTZB3BhtSta
f3+hTi7txLW0DVAxvcGEQt+Yu6GoKjLcprVGmX4ZQQxTbr4AKqYy1TaYz3QKumBTZV9pLu2jiBoM
YdV0R0BbIY4yQUtSRBan2J+wGn7xRpfwXt14DMB2BGT8R7bcanO6fmWcgdmoWPS7Y9O9VCO9vq2E
fSnSgDu3XQrE0+fV+XZpjOg0PJOmqkEv6SvkU6Ga0SDEEUwfkoA3BEfR5QBYM8ImlCtYesVLh2fE
6muVTw6YJUW0Wyq8zPTEQLOpBiEi1ufWJcDz9pLjWgh1Zy2UriwkPisP3dxuCDZ/jxhd3zFv4CkF
ZV7agNg0OSYBq/5/GGiiWORMzxMXLPhOY1RW4hnoqB8Vpwhce2nSqArbhjZj66F3zCThKboXlacR
qhbvRq9wuBJ0Tpp4I6qCGj7ZysEy6Q+Mu2wDsvsTfpNzTQA+JTIDYq7kNIsoRDw0sCUT6H4xhMTn
3sP82KUldJOZruVEn2bJgiS1cyJAHTCFeRy5cCXtXj8SeNcZwRXS4p+oXU5Gu+z6CWsY8bfEzLds
pZcGPUKiBgrjC3Hq+ov8d1BAH1eZMVyk1WL1/dJfgdDC5yNFm4Tcu5/ABEOMz9ATIIpfIgxF2uNB
fSeXUbK9gZwp8WBc3fUBM5/j2kFiWNOClTODehRo9ryvnt5DG5+f1NXirstUxX1QrTSc82S9JoMx
Lb/QhcFq9DrC1SjOshT/DTYbJOXChDPR5y5lz9PcqUVIIYpK2CKPNFkIy1CtvF1qkls0JKUDwzBN
qAEyD24e2hDq/G0GCJ8A71xRZ92W7gUIZqyvCvgAjX+scRsuQOQ0+kmyJu4cxqml2DhVCUyzHS0g
cL6NbXXowqu2Ih1VdKBJQ4iUVlPwEgZYvh1ZEaojUzW4Gn+1TCX3JZPQxKVdi2jezZvZHx86pJBR
br9fzpWat/aFCZXQBbpif4MP2AWl2HTyzrUZpVHW0Qr6KTERrvzG9Tp8FisDzV6PBoGuJ1Vof7n+
g4WPHhGkwOJu8046tcH8I2fOYsD4iw4Ed6tmJGw7GPhY1PvCv5wmbL98DPNkSH/lzgvQLL22Go//
usTLKh6u7X+AN+EGgc4Nw4jli8UeVPtvtWLc3/G9sw3nzHAfe9rC6jAsNW/VYdHFZZ1lZEsW+MRu
4JbCTtXCCntFRCP6Tx2tCcOSpao72RVi0nNCT3H9dtunNypFNqfTosbZdt5PNjZ/jw3UjMpJwEgC
9NGPGOvy5R9Tn6Y5NXgt73OYzbijjrmUkSsKKm0GwMbZa21pOd0CX62iua9YtZa8GkRN8R7yCqlW
fDfUqVTbq1iIn+G1RuZl25PNKN6zuBdOMg+7ZjJxEjoqUSaYB9SkbvvUvRCygLT8qABcx3JTMZyo
ygq9sAli7Cbt6oab8Xf1Y63fLy2b1OxKuTrctLApbgof0NHdAiRYZzCdI7UyGYTGcKEZnyGyDWEB
x5QW170jEZRBv/j1rIQipa7UnPxmnIJLB7LX5BWXHEX8svBMS4emOJ4gLNjtaJ7KssYUcH9931Ap
F0oy0aLefI5rCI2cgf6fRI0TQGCPVCKBV/qBGo+FiAFW1FNHUw7aDPAzqpK62WGrjVrme0q4GWiu
H157YmVTyrggOsqGT4Q9e9HrT1h9iYJMKyyfZO4OVxK40h7UmUaBUEGhK+PtQTba/6Ye78TluETq
vL5ozoYryeJ+45/Awy4ebnCUMtvnfM+AqikT8yK7W93TrOCQaj9u1RNoSqcqWJyzCLA2BnV8Gh4z
PeGIn6keQx7Z9yNkj9UW5WsDpDMCVksxy0GdbK2uO5/khpCr9Q2ZWKJQroe72/b5sxHFPfXWJu0c
7GawdqO90qmo7q7zoPRqzumfjgl2JAVSAa362f01JzZ6fyjugVPcBdZ7lumYO8QD099AB+cWNXNT
ZDsGJXQds4XhXlfY6st8JLrUkwF++ewP2ibDSAwfq9bPzi306uRFMm0+8rxSVzM0VmkDaRid0kLt
c16wHkWQImUhxtVBIa+/yKml/YWoSb3PnH2oWEtll4lrm7wFb+KDc6zhqHDH5/3a5FenATz/WuUy
c/PRkFbUY/5DtzbmqzQOBCgreKNJA1uzWBh4gzIqrHhc/Gr3OkK5hO2M/c8MyA/y043QEO4zdfzt
azFKipOYb0kAjENHSvp6ZAw/wwqsu+WVJS70QXpb1ITo7x+bi6PDLs1gLSaMaGR5iSeWosfQ5knz
0n91nc9hwsAd3nveHrtcJoItpJyZVMbVCkK3daUdf9NvI355Yqb64eAmmCb2qveNamFOgq3UuLkl
FefH+NSk5K1arFKJLctQUYnqSKP7YpcnIY2aO0NUP8kkDC2pHv9mXG3aoUqHheOxGvyKtC/Bt5oI
beuhU/ExtVpK03EhUBmGobNEn2MEPGAHy1x3r01KSW+lQoTwBU3/rbsgrs4c3k1iOtZtuTy0UJwa
kuTXGSloGey50f9VixPA9vRcxgKSsTcxzQntWyaZWz46oblERNeGtWpVwOIQEOIOaVh7ECnpsvwY
jxfWqNDHpHJmCIUPQ2MSJFEmBJ5i0+7zL78IDyXKdPsiD80hnwg7f3Xz8oCIPPUo3J7QX4bhBpvV
WZYckWBnNxrXU80xcaLFI8W9Qul4AbcUfzj4yxaFbp9y9wMm4tntV1yhHiIX8Tz2Sn3JvkuiJI65
+erxac84HzCbrdjTgSw9GQTH12FGRZDj+Uy8lyQg0g9CLscMJxDTWrENxWjnEaR7Thsk8eLg5Atn
/VBs5T4t3oKthN9M2Ksys2H9bIJU8nrheo37W0UDMoTdU2JPL2Goes47EKUJuGHiOeYti0y+3NIr
AUCSaFcltNXrXniLZzH0fqFMeBnKWONMZcMihl+FLc6CcSYNNV2n6k8jvruwGhYA946WBbFG18OY
3hr9Erzf1zOh1IE+B8XpGp1gzqC5ijpyiAUb8s4kOa96XrBdTsK767DaEQuP/6ZG8wMmJnjd5TGi
HRm6GiYQ3E9V/IcKsqOZgnEnD4eR7826dn5jNcH59BBuklCs6faJWkQzLk2TS73WMwy2sgbjwzrh
P18024i2g9vFd+A2WRxepQCx/HT8ws2pFEipzeEKRjGm/PQ4saqPwi36l4ZLhPxNeeu9BM/Khd3W
Tg4hNkfjt5iaeRVx/5VJRxs8jJxnyS9/PuUmozM/AJhcuq2R3VA65soY6/pVH7Xa0vOn74HQG/vA
uU44tgEbNzaHc61QS2vhmKbB2+ouOqhEu8kf6aBMBxrNJgkunVnTVvhq20beiKOShKFw/z0YaUWa
0iJgXwkhro8aKDEm0QqJIAgGMrkFRngLFFrullOXPiuMjcz9BA6tzL1AeXOzjUN+0ZnHC7NLXPfM
prxZzNTEomILOQYKqxDQr7WCMgAzyYYNc6LqlEwRp4TemOnxdKBPhw0EJbJvszDqgq5/imvRPPaH
+qu0bJoInslAOz6xloNal8KDuxhds4vXNqylWFkGiRfm1qrgL59jY9dCY28MfH6WV9hAyKZLzI6E
UcYChiuNz6jEfVNHSHGYLUPMPztCBIwJ7+Mn0f4KNursEfSXBVtK+AWfrYCLTYxje3w7q19YNfor
uYPP6rG2BW377+OGwSoQGaD7yIGto62VK9LHKKtgiLuNfnP84u9Sm8vA5QfUX8bQsEs6qxoBCX9v
SFIDqA1Ss1X9j8ORKVRpP0pqnHyu8qIzYeub9ald5dLcXbnGflQmlFotlO+P+IMeBGQAjv4YryPJ
jDBUdZP4+KTiQFtmS2b8oUng0b3a11rxokDJL8AjjAYtVq97xu5aGEhEYH/SN1O4tUU0sk3jdbCk
2adZFixlj4eiHgHBakujiC/KkjoTqvAVKizxMlYybsi2rWd7gv/SqHDSyHyqcadl8BD5PWUtJ6Z3
ioHa9DfTEG30tMu9w4EOPGczav/R3DA4546uXlnb8D2pLznxRjwtsIkrUZQtDV2MD5nOYYiba61g
Zd+wU2e+8Y3ZovORhY6AbOLdmpPm4P/Vk7IIFgmTaXYDz9N7R6H25S4VmHkmuw1+Yk3NJOCI5Tvj
AfWZTK1SKYLsMnMFT5Hd2Oojti1PZaXICh1M8oP1tnD9oyYXqRMbN7WVYuFtDj5SvWR8uMEAgVuW
86MOm4QyeRHbonuK8xe21SyrHvWO4AZpw6sslS6eCnsoz6cpK/lRlCthXxLytJ/CRNnaxxCztiAH
OgJ9k5WLsdA5kpjV1R96DSyEd/JlZ8KjI6Q4siS1xrBCz0ZT6S9vx4xb9cATlNBL3aOJKHfVbdEk
0Mx2rOg3L1CKPwRr0404eXrtGxpYyhE8dTE3fmleRj7kTRPCWZGtDhBtYqHm1avXRIit+9IMwFig
baj1QfAaz+C1LqU1I0O/qFUsXVRtWHT3wU3ypi8F+9RxXv0/7jQ5s/rcMXA31McHpeYiTRVBA8et
IapEkqoj6KUCQhnLu8CLtkhb7IW/ja5LOKc7vOZ2wudtzGd95FO0Jlsh8dmo+yf7wvwbhY2/rlvr
aBq/W8Kvc0lnu4vWKkl7PtWOWvXeTYCNYCXyoinOvrJOaPJedJDDFxaWmkAHIZ0+hWf92cRgOkZq
4wLTlTxZMHuNJp0H56/mEyWWYGMn4m4hukPdKQgs1EqafrzYqID3RmddnkjggyshgblZ2RsxSf7D
wuQ/tJ6cSyJ6qAGBOt23NWH/AGyTcrLOW0JM4lb7c7NYaTC7bmfuxv2iCgSaOG2KLeev/l90jgvA
8yaIZylaU788XyQJcs+sgbnQbtUvYv9vZZmzkzgUTQf9nVnBoTOKvCQmOs571fkG3ZcmIzg9z1iv
GRlJ2zIeWgdPg81iLOJu4Skm14PsxObLmVPQWbZZ5p95fFOfzXKcYPG6hcP5DORM2ZRMbQnnHraQ
q0tAFjATLKO8JRXa89ea40ut8sW6TaGXwCMB1w7WEh31lRlAvOtN7Kq6EDUYnyngmuV8MZczAepN
Od76EW/DDGLJh1koOU5glXjo+lvY8DwqGy3zcFC6sMjpX+gh66hDWcUMflnPx9WXR2VOZ92srH4o
baHHBZMHHPw8JvWjwOlTdPvJ2VIt7/y06Fp3AEo/ZMryxd4eJ5gnOatrM6R/CR34isKaKiIrH1SK
AoPrnwWZcaJPqWKD+wE/XP6OCSTSfLKesA4xxllai9oQqhuUYoBo7VMmfJz0/xuz3libyqEub20D
ifKM3Jp7oNv/lltXlJCeBYOMYEja+ULx3NPuyECBI0fgf5rUHyRnShqTzCuMJlXkN6MDf18OmRYz
y2HDDdrZD4VqnOIHrlhkAZkeMwkoukb3zg5y2yQanouhGuVZbbBUokYeNpdGW18V8TnMj8FdLdHU
Fikmw1h3jBIobVOtNRJ90vKOJEYZoi/wFKCh36b64dhcYVf9cRDhgPBj/dgcVlwMRqqleJAAg0z1
JYpFHTZYwsKEc5+7ZjqtTazCJfz1dbcNAyyDq6azy+JTwiM2dZbq4jgnhViC0dklE61Qn2iavyRt
Bmo3U81zsU8Z2sgLKgUYnoyRuFCMjO5pe2+xAWEYA/3GHmc2+3Hec2jbIuHhk9yP24syEM0uQSQB
VOtHfHDhCV0vpagx2rGGyod5fO6J+QOZwt0aq3fgYmP8P6vabtQu4hffSAy5vlxPTkP4Iapo8tDV
pKsmV/oRuM+AV+64BKLi9RF6VMx/ka3MzVwovNtMcMOp3yK9K/tSb74WYxGLz6uKlW4Jem1ywIFA
7YrJLKXTFEWa/8EFnSSXgb+wRGt0w7UGQ7cp5n6y/AtgOwIbFs1zk5M4SzEVSK8lqCyPHihufRXj
IWZQprQ53xdUCvg6Vozxgz0AtW1LsMp91oQtxhfxDoM38SYDz6GWoZBHVdtNXVjMSp6T/9W12jEL
LggxtGmrsa0SI+LUr1pLxJ+XgXrEadF9HXyBT5xPQ58lu++Ne1hgbULLIcYNP6rwbb19h45ckF7/
amwZWuES3GdooXsfOzI0xHpblvx5uqmyAv19ASL3rUHp7fa0hk4gxxJU6VDPrxZZpcaiOnweSfer
xqjlXvE1vYPEUhM9pjg3lT4msdLw4nZK7k9ycnEOkwnHVVUINj6CfY4l0Iwbl/UmxmUGvaRWU6tA
LF+7QTUQ+eivglXW/Tx+6OjZU2SxrawKu3kw7Hf9SgzGk8eNA5hcCOwnA7okXd8Ij7hd2yqTkt6B
tkiPO4CKUzfNTvPM9jSxwa1nUxKZk0kxOcpby82wJiuE7AFyngi1DE2mqvmT+Ir8+pY0/8ntu+nC
7W/vJ6rhPmGVNGGDG/YGflWvXl0JjxfHkSJ+zRhuCnEhOkn5yy0g8xKnrk9nbLn2oFGn86DVfAh+
da1r5XirCmXwfWt7eIw5oMTxIr4zOK9xO3mUXWwNFB9RFM4rFlFRu80z1nYoaFpu3dBBNkEJ/Mb2
1sE5yQ75gi/sJMeJx2t42e45Y9EU/PKwOY3TXB4+096MVdVcaoqmdOi2REjBHvSxp2pkAHDOmSvR
LQkOJSk7AzI0FGQncFDKiTPhSTALQN1XtKOTK9vXoxF7iY9Tnj2lLhfvV8TEv2ev4QY5jZU4X358
aznmkVNvWktfsJiLuKoHq37kTqNY6PJaXz97fMA+vkt9OaP97HxzHo/b/g5Xt1fgYtHGpqOLdLNU
euvkSuvfkNpO3eJuuxsDr8RGhmU5NzWhEeSQDcc4k3RyEPJnvs39m5VkSsWgKwc6kA9uUSsAN+IP
q2HQGQ2E6gNMd48pO4aNaVRcO58DWTdiH7zHgLQtxXZbinyhz0pRJXk6uddUo+EnMDqfkBBfIW+K
DLa1XRxozifO+RIefiHKLJgLm78t73iGBqXnZwA7QkUGsyXcSfGmyGjhIuANisItM+XVAJkSEx4L
ksM1SqRbxcWa8T+d/t5TcAZW/5s7IilAC5IygDhqtkq6jBIZb3xw07XBuiN6m8ldritn48BrqbYE
5t/fYERQxB5QbYErxks3xMSafdMs3G3+iGALsAW3o/4bL56L6y5Lbp23W7sccFApw/mp1rXgoE+7
DWW3PUD90AFr6+3WrowV20g8Trt1nTGarrGR75RY/quZz3aFHy/udu2jYnNsJbOqFytkLjt78DEI
prahGj3mqVgbBKNHdIeZTMInoWwVYNgr4jd8lmxnz1aTgSyFd6VD1vgAq5/1B9obB4s2m5oa4Lh0
skgqqMVAfwbd5NrNrrLJhsfvNfSkQdnHHBY+88FmiYPLHeqI+G6jz4p5u200Z8bbYidZWgAY6pEp
+orR7Fi4FPvdzDSkBUz//0OidDlpjTcHqpcO7HFzCSgwwbx5nPNv+/EevX7b+WoBK475mRPLrJrZ
4LvvXMDHieXKEd3ujYvjzzfSFL/qwh/azIyet93sWJmcDvalD3K8kLRMV/SAfp3FmofL3EzR2WJs
hHJo8OgsYpWtXfqwJAT8TTaGqXHUUwibdVkgZ8X5+zO7uSx1wdtyz5Ku/MV04QVHIGcqN7x4hP+L
pfrDscllETcUygpmYXtqgTK9ntKHT+yOi/2KspukZdDRH4ClgOdhWyYdAhLdOMjjv5njyPaU9c1U
pTRSZ0bBerT32zX3/pl47UuAbcqDnIsC3aEK25Vq+sqSyLD+opCez5ZLnPKv8T9vKMAt0ZClk2vz
MuQ9OALMpkYuqGChOsGMh764F4ooUXZKMRwE25ObZtRWtkdwE5BAlbykIaXI82OcSSDL0sUzMETn
HH2O5wId6d1O0paSYLflOO0zVpAUkBYuW+AN7wNQEt1PAe7jfm5IVnPsj1loLmT37N3NwLmFAQxu
DfCRxkQUoVCbqTAcBwOfpfcRQKna8NWpRZE18hSOWeyuO7GAHzSn261tM+TgnRG8Fl9iSv8tGwEk
/MOvb3MHLDLWs84T1Ks2Ip6sdLd5VELkEMabixCXBJIUzTpggKztvHJdGRabGtt6Q9VRPPJQxyvP
wosMCtJwzYHxZ+MlFo6NpScTz2IBEgQBf0BgOXdXjZunSpQZmCIS08coycUgJ8SjND89B2d2NAN1
pCxz2ZzYULA5V7ylOS/mJ3eSy9NiOM6jrf/xuOcfEBDMqv2Cfd8XTpP5rRCEwW1U0HNismyGjRRQ
d1WHpTEXZVuxqSbz3rKwzYllVbtDfEcgUptAK/xbyjQ+1tc5PNb7gD0ltDgxu8sO4x/Ws2KTUNnp
5wu4Why3/PXjb5maL15CoC/jUDjYFikB8cFxDxbtuRK0NIiqASyWAuZxYaqmfQOIwNVnJxTXUx4l
G/NmvYs9yzvgMU+S1wVZiR4asncDxx4A5hmogegP3E8JGQxMG8nxYcZkoVKIxc+um7szz25DnXRe
UmhZXiIID6TMJImiGjz08YUrQxS8HNb3aMfFql2HtYhVSFyhgkVCp7HG2XdP7P2bIlceAXbhV4/J
Up6bU1wp7HamJabcz/CJbQhY5cO91GZyqmGD7O6QeaQj8EbIkTyZXBcV39bF/1R608Rko2WuNyJ1
DC69JagbgaUydEfi6gvJp/l2hmNFCH3K0SL7saanO3wr1NCttAbA605p5D4wBZhZN0YQ/xEsiGRa
YnJA6TD8HafNX8xgx2IbWGqetiqXQOPtsiTF+oMV26QNhfWet+XwgXVYcq9zSTqhoZ5RkT51WxLb
FHpOHB4W6RaTrwCtKEtSRi+wvF94Cvv4PuCYYFXCAWia8o5dW6ompWX2H34FPpNSztrC5HgMcKph
D8Csxn769+A3Z2VXWVEJoUuYOYknuw3+CVpiyHMTaxbGg6FE11fuaKge1kRY4BaUXoGWbJnLdRPi
6rV3tlofIeB+LGgHUuPYUlX6t+6aB6Y96S7lZ0dw50vcsY7drTVOB8SRl+tQPHusj1J1TC0gcnrY
3QsC9PNhzC8GRzkD76nLx+TUBO2yfpKP9fpBioznZaL9sOJOWfoJxSNPOz9xk32nK9Yre/XaCnNo
KfWwWF2ONfnzQwi/brKDgz49gm918GGCQFt73fTACB5AnciXdVvvTFE1h9wKJsoqi/VSGzpsgqsX
azlV6HGueyZY3dA57c3QNTaHQAbn2QbomdLyKXeBnGnhEzuHBclVpiIJu71yDpY7rksmXA1mPn8i
zitCHMVQ8HSliPWPa5oswDSTiseDX0QFpIT3cbSyKa52VcrZ5yU+bt+AfPzhQVLSB2wWX1HA4oel
HfQWaE6b5vmKNwMp0gvFGF46G4BFMrGoGLWvZLDHnFQXtoAOzwEq65no24lnB+feOziGWo09gfeD
ht4VaCfWvpKwrxpU6bqvJsgR10z6+Ru6dZDiVDtMMDJKbfDwksNjiNA6V1HiYnjIKXzHuDI6Jfa+
DMrJSX3g8PxrEyJi3CAWi9sNAonKUdKh/oH5/m+JkGxhOKp6AJrZO3t3/04MD8LVZfQrNnkymD3S
qw+MfdyjqQvh5TDUTtPFH3S4TkpmH+p15VIMlmHe5aHeBzhUcsqsHSgpXTGGheIQ9BbCn6ECyQ7b
X1dVbsuEEkhi7RdZ84roB8ivUSULRQ5pdqldpZze7tyap1GSDFawrzlSKSo41deEMNUQvk4OsfMN
zjXxeKg6iafZbEqqAkohzBcTrafFUVSxlyzYNrBHXa/YbYVSolW35VwStn4q4RaRXthLByhkvAct
jhPv9OiayC95Kbm96jura2nzkhHZbH0cIeClZjE7gbqMCZzGSNFVTBpCrdKnHXwTBtcpVsS9CrWH
/KP5KQKcWBmm0Z4NeBzq4xWDxFzZJqYit0RzEi69wQpKZ3enBaJKCJnr+qrueZNVkset/BwpnLLI
5sTVZ7fUup+ThxsWkE4NcmJFioOPeBcy5OfHQCkAQQSwbE0DcmMXL/LENq2SLRpZd/zAzcwUeBws
/javRpGPYwNWCDT/0CZ3Auf+h+ZWYFa9qC1s7G4LyfJ4zpXtY+frABORfZyf1UHnuIURaTfopTH5
0DDrQByezvmxMhjV6JCW7rbUBigbWKvFelc6sG2np35FV6s5kV4JHndYpSWFXn1b09F9sO1nKJvA
+ALMOEAwg8xIUKj6skGuHluNb1EooEm+ga4SFK2r/3DXuWzALQtLxAskbc/5PDsOgoBtZwnIn47G
wdNMoIeb0AtGeZcD8MOKCZfsNuGdCsxoUEf/tNhS3oiNL8RUvr8Pe+wwYSwdd7v1HVkcn81AN9SI
5xrHhqLSzZ2e12GWtK4UyHk7jD25OQbB85dvC1udASnA/RLHJXOPPwS37iUNeuCsB3S+3FXo2jz8
x2/itnhDIgR24IH22r4TonoPrfvfapTNcOvm+aqDXO/ua8GX4zHDQJWKMnNKKGrj+ZQJnG7QrgO9
TS4yFbaBHSQqDJQrStS8OmoxeGfwMVw4JFp36IO87YIY8k/Moa765aya22+uZ14DqY7MZMIWklWs
HVRybqx+CK8kK0trhI6QeIXQt3vkiFFrMMevh9YN/WdR9M5H/amfBziPrGG/1Obx0mLLcKdTmw4b
uvwX1fdO/tPIYsBvIifNy0BqqyuDL/g+jHbyEgovxdDyn2kIthZH5ru9JTx+6IsvZ/184z0GMzTq
djOzImoowPnzgoOHJ5aSWSuKIleWP1V2HSD0RmgyCyzLq1mdPGuoG3vuub5HkTAqQHaIIJiny8Ac
lyYbU2GbYVFpJn4qX1DBZtv0+hDIEk6eIlpWI0f8484OBd9+VYlAqNw46kSV/54kAtInsE6R2F6M
NHdXOK68fRyWnskzlXjaeaR/s/ev/svRyjESl6GW8biM3OELbzbUtya2OaDKVFuotWUsIhprXT7D
gfYObl03HWurHlaHt/hyOk8SOVTg8az166gcHQ1EO4B1hs1EmE3HDHuP58IQ2GtMBczTym/Oa2Zk
Xr+/xEE/2OKZZxy9X33J/DwNFIzeGKZk09Wur6v2SjcQH67LjCNAmlyw23SsK9Jy0GXbXHXbjJBV
LW7m0fNxg6EDzmvd+WWJ2u1C4FknMnW6a+uMTBPvu4ONOm+w/FHvg2lAreeLDC6d6J9XV1EtbdOV
xMxtBJqgx4HL8inCZRqjs4vUtaqkPechC78t5G2ZsK4AsnpdAqlpAgerdYB51+6M89207eej+A0+
Yj2sooTgX1o1sP14wp1yLHGuASWdjab5p4/svb2idSLzO7I0GkycO9TNVvZoNGWU8xTNfhlJqgjC
aLwtxxm/3PCTh2dLVn5qnblN/MYROx+fvXkQUBRjfI/BFype5BZMO3NgBdyQHWp/PMJdG7VrSOQk
Evfmbbp2W1TvItNGCQjT2T4OZcd/JGrz/2ds3OQQJ/5+F7mdVPQTUPQm9FxHLEKmucrfRKQxKEFu
eBKBbPv5KrPO6XZuINBydsSacg1Zn0qV/UKAA/v0GN+kYWlQkklaj47tnnI4bQF4h27AEo5G3Wa+
w+05ttWO1ZuTvWhJFVC3D5g8MPmnNVeLDdrnC6LYwq/BoaG/NyOtNe76iauMiPIYQXMnCZHUoXJj
VcF+zvaEUe4hP64sJ9oVWq5eOP2iEPr5sUgf/unjJVJOOytnUMOXc0BzIBu3w3vWyW39BATzjkX4
A9Eqw4JtSvLlpIoM0DI0dH1VnwCQJC2sUGBxpwpyp3WHQs8GHD+hH3l3mB5ZtY425krPI1v2Y21o
jvFLRQe4SRo5PHXAxhqga/2cB4OmMCdl2f6btCyP+HKSBBkfEziiFXpwrJU7g/02WHiXwCbt/OcR
mqlyLgLbhqP1DGKDvDhx12V25x0r7EpgLrKri+5gM9yjhpWqhLQPsEmTyEzx1IjBVQgwJl3V/5VB
r3eQqVXDR8hZL8Mdtfj/zYVZsrL6Iwyv+E8BnyDJiklX1rZMs+BeZqbduMZPfs80r6OhupZZPDjH
QJSCyuGJOVnT7+dGwOEPF5pr/1UF6/ABYo8u2qbXeAjQL/uo9a6AUnN46ZmaRzKHzd7tjt+eW+nd
tm2/QYVyHByUmnUyzTjD6BEugfuF3/fpYv6AySElT1afRP4g5MAytdYEsXCyJ4xgJ1FC0TJJxqFQ
6agzdaIJwJdYQzyvPCoYUEznYbZHF3iyQZVMlJ5XhvzATzwH24o12AuchLqaUHmSkUZyYsA5L42E
fzrhGWWUprkM8AeRyzfydbLGIaS0b0GeOaasDry1YA6lLplXK4GsmLawy3vizcIyCdcAOdCoJq8k
8IMwqHa98MRc2/Ty5beVQ9Vp56AsdKfjaoBObg9kLq9Y+d0gqW9y9CkJbOwlmm9pUNKDyyIg+VNr
yqblhXIcnq1bjga8TEeV7oJ+X592KgsqCKp5LrdwaJP+ta4LymMXLQhjW56vFSW5cpS/fSfULA6f
f95ufdsESdJC1SpGPmN1kPu1AI5ELSIhK4mIYL6QkjgtZ4FibhbwP9dBMqSDdYPweZt+NGBUqtxO
Hxs30y96kiaknksDMVH/mLslDDYNPfrN/q0+C5DPavQinVhCOg2X/bHCcNd/MFU6fayu0PeSP+qV
QDwnW2O7Qr3kkm8J+ZB87rNQHIxUpCxmpBo5IP49euDmGQrCmqFS4/F5b/eaIKZiaApV3HuQ5ODL
DpGvE1bLral3tUxXSg+2J4GxTxxtcriRZbJBp1EILn8nDtlSw/UPkotowjTkqehiSAfEXt6UvWCV
VfqiWbYiAqHsm2WfZSFT2KgzR11ex+FZmpCc0xRBuOMl+eKoHVB3P+YKs2MrpLW4iupfi+QpGKGY
gEIxM+9GLkwJ0SrPWIsU5ID9sw5qkY/lb7+aJE6iuvWYfuV9YTNiiXBjeXp7eSq3lPUHCq1mpQc9
kTZql1W0DUfVPaj1r8J5rld+N9WzsXH40etTO6k+NzrXCCtqHxkjMwTIBuiEnrVdMHKU5dCqDfRg
F10Cb/1mOjBrCeyozLZhT2k2CyQhgk9FyBHMu+IyXXWI9t1AWFKwah990SS6UpkrC5DJY2q/5fOm
WSwd6OY75Fz1+pYizRGPODRb612h/AOb8joRo4JT4k0Pl949csvLieKUQBxIEQxPHa6OskC6GDbk
aFqBKX+CVtWIlbiEwHiEiaD7PpviCBxwzLE9IyvFe8gcZwgvvatn3cJfvLHF9Ig92ZhFnk+S7aoT
8OyVZeZdunotp5P2IGBmp3dcQ8fItFdPvSOuzh0G++2KDJ9/55WjTIlYFF0cRpeaxqnx7V2vYxxG
j/6kq47ChvWbVqdThM7dkr0dLiFYyNJqoYSg2gzEEfL9IE5Uxvo6SNB3aPu3OWM4crOeME1k5N/D
hKhCKwbgGh8xTLe2cwzPAZ/LYSQYDs65n+EI5qULSLAtBSFvzmWnQ3DGS+W+2tFiJhchD5EwBGuW
6CjyKYJv/tHtW+fCn1TiC9Q61W1qvCIEePeJ9UWBkurEeASmDrcjHrH14bcGQbJfHnli/5EoBkOt
/sJOEf/kHDegdDIt/r6un1lRwVosC9eMGofeu1LD1sEJi78HU6lTErLDM2g+FIJBfDoKm3XtKeX/
CQiBoa7gYxbtCZKfIziWD13MWdfjC7H0wq6inyZhNQy6Xg30jrwCqrVEal7xg5KSrdHB8g5Bxfm2
hH0YWkySkfYPFz77+bhDvZt5cD3jf4vzBUl1ctlNtuZ//kcATPOvif5tBdtmed00EnA06giw7CCh
FB8fTwbf6v5diaMTj9WjxbkIIEw8Y4Sc48vSiZNL9b9RvO60ILip5hfMfFkBL9cbZ5tLj4DP1Mpi
CDkBEFTvcMi55+xPsWGWRPLuGshNfbSHYjHpDtYpXYPRq75oXeAvEtt4bs6R3oItWeMeQSsvVlUf
fCtrQqeCCP+fu4Qv+ffB7aZgsuDCJu7BwyEqObG1v+W1hgwDo0yvSxZbUz0UPsQo9iIB/tBrJy3d
WMHeOP39huMygDGBGZkpQwgyVJ704/Jdd9jKU4iWxFfyFvfvH2POejXFKlrGVM+oTgXqtZuAF5bU
irfPpG/TOGpN4y382lCIkFHMw5rqC9ovBhfqZfUHs/98fZ2PQibcBKaN/TaXG5X0HixnfuIHhLtD
rGHqiAvwZt/u1SoQ8DQKqsJv0wDYGUxu2UUAZjgmLMp7uXXBDtKvDumTtZtCTqYdcRyOj+6JAVjX
bJXQE3odAheueOBPTQxDTWDeksP9QBmSWxla5fBmwywKnzuXRZtokHXyP4y0kZRCAEw6kQ7QZWAR
f0EMnGAuWr44Put3PkqolVNDLp3Yq2OkysYheO79JmXLkQf0s98XI25AUgYes9DkrV8stCVJO5vL
W9Slrff7n75G2Wr+URZsmo5VKQlOHC3fQENprP4m6aXjSpvMDV/ECVrMxNCmL7ObSPC5EH+AuEjR
BzBc97aGQNMaGQy5qrmeR0nujhK8icOe1LzLNFcRibSYLjpwf3IvrC1PJSZF1nqN1JrCAOj8GCOQ
997+O84PKKcHYxlGeht03VhjI1cj60Su5Ycf6wbNskE/HiGqm75O+NOCq3pSSK9ktlvvXvtdUTxd
4wcN0SNJ95HwOabDT+mnI8mVUN9UNRUb2jWcFUvtRShaouPfpMolAlUmJxlGwqWR0Vqmwg5YP4UI
s/D8d+8KwRP4l7Wof4+N/Il1kAMSwgDn4ibhzJ77X7NiYKHYh3sau+UIjpxdAxaRBSB7JjDLK7Gb
7ICgxoAPc5rG+JzMeUCPcBDWBf4Hm+4pPk05GGeHKllveIdLFIdxGGrUv+/Sme1OB4rPq6yUy6UN
UHQlMtOyXApcseIzlQyqv+CnHM/fRq13ZC7sND2j8455ArhH6F1jUksdx/PX9dAlayZQ1T7a2ZHQ
Jp8C0jGLYj55o2y2oq0vQ/YAaaNofvQbp4Sz8ROKpI/dA0xmbvkf6F9LqXxCEqIy+td0tmsMb+YX
FXzOFRLQv0KK0M4GNTm2b+hrqOCe+Y2FQhwWvhCBWyHf7BMiJxPoCtevhLp9uBetrIUNuKwadS1f
lWOnPDHwzVAyZlR7SHMzP8PHB9DXKD/YNLa4jXqLadWPdWISBNB7gPsYdDxmJmFl+ysmOp4kTPqg
dHjkyOWMytH04bjNdcqJvkPPY5s1wGxqYIVz2R+jXsjaZ22fDJKUt8GcMmQTtWniXMKe2BLd1Wdx
p2CqhNJWiy5hN0y9xLT+ZbOOVZ0w8XeppA2LNC0ELFM7t2qZVRE+nwrUfv2/iHTfPDmvTSohMqPW
OBX8/JQlNnaIhVB7G5P1JyWxJQUDvJ8+IyQe/st2A7Dwy+v1nl7zrxw6k9AzU9dv4eKOjNCBxn7P
ggvB+gq1CW5J41eSmGYy4f7rKN1cqYcD5Db70tuhBRsDe7KarQ2v+iitTFkIrzlBnxtYW6SkAqhX
uSI/1s67fuu0qCBEVZR2+0wQ3r9535j/2fIAEhUCY+gWwaAzJUpW7wq+ncYtWehQdLM3F5Rr9g30
6/o5qfWKYpykn8yM+RUNcTmbR61PqfAzolPM52CeUBYyiprQdvaTUok6nuDGLcfX8mczilXL5gy/
YdCCxZDIzbmQp1D+dJBlxtHYl+zXzKhYxH/C9Wu+un+b8ja3BkBBKsFe6zSFQ6UpWJGeoY6dAi/A
qG93tnLNJGqIrDWJEob3ZuEEbGNSf2B3P2sS8kyO7AVguBAxxFlE4n7TuQ8DisCM3CSazyrbZMhd
Rz9ILn1I2GPa8OJ0JV/j7g1g0WQzlbO3eViics4i8azo3R1od2p5w7JWc9Rvo6+izgtY3CecfZgz
BlIKUVgVXCU6hpuCj4YqCaI5DZrSfUHl5TaQpScFuHFm5iWKWimC9nKKlPwPYXDwuZOrob6UvPej
uJ6++WzPc5VuheFUZOO+P4uqUKCQ4UDGjL311+nAT2Z18MB7K/Fch/sIG6PgC30jX38Ov6uuvSDZ
0ESWITyOq3Dici+l3hnfJObqYOGah2Zs+z22yfSApqYVrs/30NLSjina/PnS4f0R+H7I2IE/x8F/
mgjhGEew+ZTUZZMG+/Qzs51LJVloLLaE5y6u2sCt+JKycAiwyuMraioaZ3PqZP/Oe4Zd1sSMvro+
DgbBkuwdk6KsDolhLPKmMXQy2Qh2a8Mjs5X85fhK+dmV590u5oatgF545XVm0ojJKna9i7bM1Yly
WXuUDy4XIlUqhxunv4J5gFvGky54OeTr4rRSz0uLrLDBIj9H0f12Xx0KD8iOcFQ0DnEkew0sToen
53Vx6IyXVdLmq1xkR0YGeh2pYrFODwGGHdTwA87JBwEw79Lqlm34uG2yNvCBOCzYLTJH8LHspWhm
e+JFSvBtgrIJBfmPqR74nl8XLsvlMElHJ8jffBlHV1OOwN5nhCKp2ZA/695AxwKId4n8VEUCDSZD
iuxniOQEd4xePsh7ks1k8AxtRP0CjlSYpAU2vsZ1kgmMjwL6hnSHqy7z9JmDSSLQiQmBThsOt1+C
o5LycxrNqoz15v/RFh8GnuqvDH3Pnzmk4p8KAzNqmfps1VaWuFzpe6/bpcB7R72hGQ/fanOwSqEn
7KrCXjTroBBp9sSibbouiy2nEyOgSTH8YbyptPt2BAbQPJ54voVGsK6zEKKzP5DB4NdM4zVesnnC
fwe8otnnhzH33AHxn690gcIxX6cSqwbbP48TQsEPTI9o3w6PV22ex2JI2C4cbmzigqZSD75BrAPk
njy8VHt1CrlmJwe5tTFVmVFcnt8yUmThtMl95S0sk2aLhzDtkM9OuGKP62BECcG5JiKsWHdNSBFe
dE88en60x20YPRP4rJLnP3UL7EhUEaPtRYjnmBySRLbB6OLGunX/CEniJxqG8lWX9FmEiXDfUYXI
ZctxF7rH15++sywYVw7UBYcEOh1p94RPxHtdY33wsWxkul5epb/LgCMURZ0M2TRvMuiM2YJgyqhE
fiplEZeNuTB/XNlijJY6eLbugH3vQfEKk2yErTv+ejFUJXoVLu3JQurs4M2T46Pj/uXmPOFJ5PHB
GT6dCNheywpnZQ88jjOgqXOEyC3hihxC/NQWiWZu1yvZTg2NWScJX9dPWqzxV7pPUZRp8Shg7auH
V18oTt+dRHIqi4Gi7C1Uso8piixz9F5XM96rGe/c7Bb9PiMoOV7TyjhI2mBOWQEa3lb+S18r0fxz
d+zmwFtejbY6EBZFaCwNXzU4bYfkdKgT45J3hKpK3mVOaJh/f3X7pbGgBHV5tmuhx7IVmWRHhoLs
irOKxsq2I6gU3jx4roi3FKdq01b0DY4JKisvP/owPFtEubUoOVte19XLWqqEdDVm5RuUp50qAcwE
XGiWol5OtezQLAzpHGhTCPEaWsY0eAzPiUbDDh0/2z/IPjoYhP+9ALfuuzEgCVbNt8JwLSTj93Gz
xohTMZ+bQNWNOLJFhaTcmdJ9VFBxI2jWKV7/OytZ3mgEDUPMyUdF9nIFSCPT/8nJAJhV9e4fJyF8
ds9DckyrPxUsDWNlct6nOGaC/IIvS+pBPadHepGGK+uWp04hV1NZuGLrC0CgxJYvhxQZMd4PoKUY
otX5/3xeDHLyPVw+Dy9r3lkr60T32uokklQL3A0JKxHrK9e2pqxIvqodwJj6VxJzBPYsnH+yYLgN
nz7zmo0FLnK0EPugHrO8O2GQz8XXmeffCDzmnKdfdhD9uU3Ia+wza0B5GHT7DipZn53+IoFo2CGH
XSQ1S9HBoAOqg/6ViGJBTg4PILJgVyLgLiMLDblO2ALQBYcxSUQnnb8r89NabSezmuVtmr4EXhNi
1eWIfW0RbmM2VS9bBGj+Rr11biDGAtunb2NMnPmn3pkmBYZYab4gQrMkzjfFiiM1UB45b17q8r7v
PU/Sj4DH74yI9tGF0cZ1Xs/auCToHZ9ZhTbUDAjFqjbOLsQaNNwkf6l0+peu22/Pz7ItUkRr248I
a00miDKnDCoyv3qVrasglk/hzYmoPAa7GH/9TvmPaGDS9eZhhLvJRBPTcqt2OkidUH6QpywkdJhI
Z+0oN07YQhArnkJ7glYddI5NE4A8RC0TNDOtpRBZ7bvdRGI6trjPiylx60pRXPTpXnVD7WK0LAp7
LACzq9Bsatxbtc9hTNjLu9B/XfD9hGrwLI7vkm2sVN7X5ohfHxyk/f9LeQWsZU3zpHeNaB8pmlfB
laZDlguE1nRNh4E0g7bowQ5ApjequXSFo2pN3Md3FW1fo6P8EqIoM4Um6ozcD8E7b6P8rgAzReZD
JM8uicM/gZVTrTWUNExhbd/5Fm1GOioBINYeDi5287ko+4qbpmWIk1pLCVVsfbrxbpiAvJTLcQJG
5BE1Bh68Xj8DCzxywuVlSOwWIz1zkrKW7w+uZmCtVjIjTpeUmSuTh6DRt1TNti6O7V+qjlXcat0S
8lh2vS8V038CRfhCNzn4MHYwVL1u8ouW1DIiIQuFBc/uzewaop1xU5Tow/aLVrHnjgMMxJStQuZB
p0Zb2uEAx1UdvbxEo6eLfWnmbHfNVL88yuOtR+/Mb1zS0R5WXMVLongAybnnE+CzjW4SEdC7GmZx
wjm65hbRr1DIDFXxIompq/S/JW4ZTMYSzdqU466d4iog7g5aWbtTA9J1gGHin9hhcN6IJa8fNnWR
CAPPCKwwQYDuWm6mTPBir9qFTmIPzN2HXHRTmvn2Pzey+oU/kCZv+AL9tUObK60r17PCUBtK3HzI
oU3631ohtPMLX8aT/J7wC1iq7lUQjIh0JQ9aSJhPfcLIRmq7YdHQ7Q3VhFF8wHnfmZ+dw4ZRx0j/
teAyMUvukDi1zTUdthLZlC8vZJhs0Ku6zkg9owrmxXO2xBMc3a67YlbOpkLtpgz8OUKKXu6rIEwE
51mLbNfRoq4hPatWcrASdt7StTPSM/rADkfVp6Uam0gTFO7zJSgYBiSIpJqy3rZSpZrTDyQ5GA4/
wxovoGcGs4whAAx///UdprUKERq0GNg1uX7OSo/kcZgXy7BnAwgo4iw0qsdXO5Lt4Ybm6o0gOXuI
WE2kXQJiSL25+Nzu6iGoCvKAtz/lBCVZGK9Fr+U8I0cwdvLxMBm06/loRsDEXZNzrfwD+ARicOG8
rg8WZZ+TgiyzSmpFVliOm0R8vlPVBYYIYr2J6/W4sQxBA3qROh1PrwmprOyYZD90iMoqwmn5P2Z0
6zMdbAkghAGVYXRc9HX17b16c+h+pom7FUtJ9SQxlsZSR9h9+CSr/lQfj3y9RTDcQ9MJw1vGA/nz
DBA9mdGHyy/b0HORlqdZA1SL0DU3NpLT/ju+faw5XgjNKSeDnBPzx++u7bsZeDEcI8nn2ox28p9n
z1UX7LjvK5y1uK+UMbTL0tsGP6UnOzlWQ3Yx0R6cr1qHT7drCAU8Ab7T5fm+/9QFPeEcxxRfT3xa
+DagOnJrx2gHawevs+MQ1AM5ln4xFPM4EHVkxoh4D8GS1j9Yy4UEYLI/ui0z1A4JNANIT5oWbICU
Q9meSFPrL0WW5jDtKVFof2SII1gKgArn+vrwUlE0QMziRLKnnpylWDmSKesr915DurGDfrvla+Yk
ItDrqvQKlNYFPA8Nmn6Mzk2HsB7YB3p5/vKx1tbfBzLxNxZV2nOts9oRk2oAxLDF3G1j01HZp2UU
kgDnBG2IliG63rb2rmO3aLs+diEWoVZOtyM2feInX1KXxWoX91QPmBWwlAZ2TvqsfXF5WdJVedM+
TU2qhW8y3zv4OM/P4teG6jP+Y0akD5Zf/U6e2qI1eWwB7+j+ydYul0gluZxVVseLIH2MzQUvMJFE
3AHH/q44WdzPR9KxhPfUvlXgoHQJA3swGNVk362FoefNTMXEaeIDPOVBZkTJ83l1EFj3LD9JiKNj
DLTW+dZcu6eStuZzxdWWs71YiorArlVTypyf9rDiv3JT9w082KvkJncO9zKLZzqoWxdDyPT9K0Hc
jHzPICQofyrfyNBu2R3LIvsuuPGNPjOK2jF9KIHqOk66Tg9XxnmI72ffDMdaDw88R1m8RqVhjIoQ
lyE7i2rzYegon6r6fAVaeYW2fmYmVBKMVz1wsSOIb+rcbuM9nGO/+0wZH0WtGUxuuMyKv9xcdjhm
elzdYC+5sgmcYFdGNKtqvbaQ2s35Q+KMyZfOa7XPRItBs+JHd81pkX9i+KCLdhF4IrHpAoQOPa+n
qk8lj62TN5/dPzELNM5x29gYSJ++tkoZiexc/bFauQ9pZ0Fu2VwwFp14gm8OjJeYOt72Zgc4VnG/
Bg/pTkCzF7gXiFc91LBD76xRYFlM9s0sS5JzemsNwVPiu3GcmiYR+3N/i2gkDbc6D6q0Lvbh6tAS
aY2ZT6N31FCf6lAfRoQkOKdVGlkaGxMttgOUbDckD32D4UcmyawWzv2mzsDdDwAgV89JGORjnssP
VOjrmyVTCiUOJAMtFpSjepxJlGtHTnZuOxxRpnGdS0+GvUMXeI2Btq+sGyFnwni/hPMEEGOV4KBi
ZNxHwoc2qsAExwgBsWpO4VXc8JCQ+fFI9e6oOVCKUnfORi4KPuiHohLQuHNrexzPQZAcfXigRKhQ
YICPG8WFdO1/4gQ3fEXl7buHTiwnRKFs9Tsi42gA7HZise08oZ9e3mNGgACohGsXWG5Ku9/q819R
GdZsd9JTjv8TXaKnIopHH82I4CS0qkx6MjH3uyQVVGM9va1/tu7J3feZKDl2Jl999D8g23M/+QOZ
9rIxMQph3xYW5qWqrkSf8nKShWa619+vyjL2p+1pXz93PEvyAEvsIj5+DV5uR09Zl/dRaL+WmI1h
N2jOL96le6PCDzPyMJMgWGV1dmjfK4bJSRh/LJOxQDBRlODnOm0AFm/NeJb+RZ3qc8KlgEdRYr+A
bBtGrVcKkB5a4nz0ZQozG9LnonsQhxfTeTY2kaRhWA69I6374n4jmBre4AWfM3htp+xKNmSt8ez3
glSgPJ3LPbObCKns54b3Q4cz3XF4b1WUwtLKgTwLTj6KK6XjXSoGdDGoqoCm/BKMvRbPZs/ocOcV
E9DGE1obRfBgOEVRfXaVWIszpD+9nWyxFeHBokyHSh7u82hwNyQ6EB1kqONnnabW+5QGgm42n/4s
2SJUYJ3/RbIIhIDzvrkU9C6NkYn1x2oFSpy3HQUro0fejTN//+A2rJ7EEIKHd9WzbT36/iZmHdLy
kszYNodGQTSAX3yqB/+auIzD8hmhMQtrmawd4I1q8fn6BYg119HacXhNhLKhG2+gzivwKoS6eU3B
MwzZFek6pvfrp+jOXmyGhtJ/eYUV6rIRp0ovxBLAJCX6KVWoKCbSWFjtLFFYbM6C0zUocDZhNFBM
LJdbU0PSI30S7zxRa/qvoEfRCENUnm2ACMYKF4z0c5e1mtWP/OaYHWPybvfCfT6MGiz74iZWpoVQ
Lc6kIxVMCuHMa8icAsVeQbqfrh1GiSrLpv/8KxUbUraMyQ4yw1+C+TtzfgDdTnajLhuE8h0it8A8
Y6dtTBZNRYq1yMQijCA5qTAhcR4u7ataM2/vd5CwZmv6VXAvFI1HiMLv7nGJlwbHo+3umxOhkEQr
VqjFsWtJrDtaO3gGc1bAsnL1gMwiph5j6976O7AGZAMk7ty07qBpuahmp/kdF5+APtzQqRE23FY8
CT3hIY3b67zjyOQIJyOxOle2ueOWOygug0DhH3k6Q6UGj1Y+1+dYps+m4dAxVY4Uvn0ZCzu5cfCx
0e99dRJ1cxYMEIKWrY8fHqQWzKo4Xvk4xPw0XMSNw4yzf5yGDmQED97aDDkYri9XNHa6uoYu4pUO
q2/hOlpl86CidJruqX8jDyV0RbCONAi6ZNJ+Bvx8BnMm4DcqMGd2duk2HpnA8mSM4SCiWYLiOyGe
5KIBKebfo+StNCiyA8xcBGvnUJRz4m4/90OQF5/S6hUl3T8RU2Eg0flzbTCvEh4lstNFA+rTP8FW
p0xpVAd4inQ0rnt2YwiweeYwCWE5mky6p8PG4LoIjIeJRuJI4uj0nHdRpWEpzgb4a/1+nGTvlCRj
yAUHlrY86dWAXz0rJ0vlqN+IvG3Yo5DqttnIf3jLLR0xN5mM8JdojZH9DVyrvD6Rsx1T7yhLZ2/U
5/OC7enPFWKYbYgI8k1abHZbcWPyiFN/qNZVamfTUcZkHN8J3uqPj0ac/BE4W3h79TWav4jD7rcq
/Ac7IrFLIdWZHH9FKWbA0VKBtRin+Yb0gszeAcM9MwJ5lThhJ9AO5xt7xSBC1z5/9+si4mIL0pX8
w9dAkjOXwFrxqrLsBi/lcO5LDGZ6KZiJgrhK88n2R88AbgLqMW9kcwntEJjV+z124qPcOoymet07
/9wwPripZAmjPDjG4U2SmbKMyFssoWiK7h4GosEcoGUeiOINDDb3bU23BHy00EFao2gUjex+s0DV
OjpQvOJN/U01eOxCKBv7tTN1mcvvLveRigOHJdK0p9n0ABpriItC7/+L1w8mpVn2yXDxzq3ueOo7
hGFQyu7dVC8zIj9kId1fo4Yz7tMmKKiZojuY5nacv1X9xj6DbihLPwfKg1ePLSQvGXWx6dtmJ0ti
MkAYTaMLJI33IZ0rxM/NTVQq9zqXyNnZLhJ+2lqf2WalaxxooF055125Xr/iZgkbGpTn/O9JXUAX
YphqS6p6Kg2s5a6ncMsb0dD7gTCE4RV2Pd8N9NDIw8e5AnueBvyp6+y8Y1xFvIfmELb1BDm7g7QX
u6kROPMlxx/xg0O8sVyz18StClP6xUc0+VkgAWOiR9CosR5vBWmrPX0Zk720zDLw5hLNqKH6EATl
ZkMzYgPvZRABDj4NIqUSCaXjkMWOazLKSF1ZqP+A77Att/OhpX8tdM6IvBU/hO/88oiDidK+Qbd3
imVSqienT/Y6CWxP4T5Bs4LaEI6tUhfW3PEaOWd/L0OB5oWg6R1KHNc5ukD6MubNJ590EAhOwbNG
aoAVSJAHuD3us/w9q4BobYyyhj+F3DdZBYdJiKwfe5HqR5bn0tht5aX5C5T+GylVUkmFF+awl+rU
eJvPBSTciIYlvcu8gTs+A5/eYuOCViXPObQkWl3DRaxBD/SmFK9LTvQxa77UaUB911ZaGnpwP/Q8
DcK73xQ/k+ENyNlD+Z0Ikw8Xyawo1r6L1lai/vgH9pNCu6uSu4km1wpLksTyZL8pe8Y7SlC0uC7e
i1XtpHzD7fJQfpg28VArkazOUqT9QNkplJ8bAqAx9f7bTbg9D5erT8p8R4KxVJHurZUSULMrkOi0
Pni5tGPKA9RZKhYKNea4pDoH0CyXvDUaVEfRJ8RPuDYmGDNjE4NMoR9lPIbshKnTDNICTaLwyLfX
wMFq91CEnyLdo0UHQvDmM5lgwrUpOis3cMuCJ+sRYxqw5SxPd6jATnlRF68bvwdh8N8fIC6kKG5j
eP4bdAqNTv1BYSPMRYuih62n4yZyAkX1BPdR3adMF2BxwRCxEqFMRxn3mrE9q1C6Htq5VyjJG+zb
i/PwL0X562RFNkHnmq+L9mwjfJcgTbiaOjVQT+MSmAi1c2gst9R+vJZu5Uddw9tvVZUwHxWltOER
sIurisIbMMh+qv7vo2vxR0fHDpI/O2RqFPxQwTgKAH5eRA1L+AZtLbeOuWKAncGnAK8suPiGekg0
vghWw6Pn3mUFarOhJFsULA1ygBea0NTdp15vZFvlg62JtgPQ+eDyE9d7/ikfQEJihXVKnPdepyzH
dtKvfTwmrzoRNVgbqi57sAYSO6DodkC+wkxSNVL2cHHHtnXMCdisTs8G/F3uU6NilcmEcDuXKdBm
wvVrB6hwItgS4VrcfucmD6apDibQ/Y0KjfEV9qSsIcYNtwI5esN+GLNrBBFzEk36x8ftwfQUAzU7
81kpmaHaffNlmmZJp+3fcW5lTOT2CzU4lRKg7VwWF0t9WMCkFHT2dMeNV+xttBKomReS8VTz2SLz
f+4ftuy3uOKJkfzXqvL87TDV+8RtizYvp83VVssn6K9LphkHJ7sHPoqttCzDFj6Blq/m94KE/j7x
L+VVVHKdXJ4DDTEfzQPji57RP6JC4Ju/9R6wiWzPmRTFYYZdxST1lSandxNf2wxiqza4BWiYEqG7
j4KYkon+iWZHDK3izw3y5CJRNDrWgeOY8YphERJ7M/Tg45iKB8FoMl5ta+FvyhTIGQ1ydiUzVAri
11vjSrWXwm5j45IjprC2tcOuihQ/8n3CYjMzVtZj5zzZ7Mb5rXs4yP7zVrQXtvQmSfAZotkJQCUa
F8KhoeLCmVitc8iuF2mcCkJM/ZvNc3F/KbEc4/NpNAUSuoTCNZmNcCPFadpAhsj59AB6Xu/nMErB
oQNs8azkvU/vv4+OgKIhzYMyeFwCp57PWgqocdkRS/OklfKcY0yfzAyK1+WxEffLIX2RaroPq10d
YeVIB7TQhogscY7VR+gt6HXXkd465SJYQYuLb8SR2Z7RMjYakM7IRp8HKIYcAWJaFL21FEa/9tPF
ElUvefy3tTrpd2y1VnzTC390oA14qUFffGwjYmksQeALd4Gy8oNI5w0YenIu8Ta0GnKcEJJdQVeo
CfuGIg0VFYfpCs34gXx1X6CCv80i3dA/0myo8+YqsjgokdqbKBXXi2+EylqsunnYnYK2lVDjolEw
g5fzX/HHHD7SL2Q5M4lLfbk8h7RkCxDHU6citq0CpiCmnjWkDk8yyiU9ubVL603lz/MJ9MDOdTXw
2CAd313zZ8219tOOuaOW+NzSzwC9kJS/KAOumdb2fwZEngD9DBErUv4MRmAbmQg0EonmJNU5wk0H
tCO6Chx/2p0u35y5WO2PIWQveKHbjo+Wgi6Swjz8RqgFYogTiGRO4O3LCieBjveYjQLLPSDx5M9m
3p0XJfCJF9c9F502GmsW+Y1+7wkzKWcPucZ2fF9g8GJMbFShMFFHvPn2aAsIxxU/lJ16p6OVXT6g
rYwO7oskJrrImGAplXWhQCDfEX1oHlvEoM9HCH5AV91fb0eoaQEvpuTabj6v7FbLW7bhfgiMhCuO
bjUeXGblcjNSCVggV9DTCn8tpDRiEjD7nvcfT12+GNleWJqFe6ycnVedSSzCWuaAkghAkRrN58Xk
iO333lTWxeAHfHtivozFegsRg7yzGA8Dk9PmrTz40Sewgf73Vbahd86oQQZfqXwKF/mIFSE6DWrC
YXG4yvsU1LR4xZpBDp3cCLPzjboFlBG8adD22K/3ZvKh4Vl/qgOWYEdmIM+GtM8p1yklZk2I0z9n
rB31VrQ8ZqlOOtxt97xqqYlrrXqkXTuXNA8SlqeZEBSFvz6+88JKgNHxDdS9chMYO/Y9vwzHjkrY
FaAIXbtfVJBj7OJhYYIQvDYdvVWvflclTrVTNvZMp+ZLKjfVDbhuOFhnsaLFGmVtRs/wx7L8XfxA
3DAbVo0vYmMzY70rk0wtQfhXxKQPMz0F2TW2a3lT4aeJep0H82uwHTM3MiSXJ5aeiF6Q9jbErSsG
GrFxZ0niDHAvcaEg+rtwYRB3BaBWWnOwd78NJbeJ4Tisw4gcoIwoPHgiYNXieAoHvoJby4IVMNuP
tNoO+5dfLQ+j2iRz7N8zBwoaVt8k/eYqoPL2O3onMgRwwQ4fukNRw0Q4WzJPVFKkoqy876xMMjJK
mQ7kRZjfcBLC5NScro5sJzHYjpXBpXABoj0AuNpaNQFh5PAXHFijJe/P1mQdbtnQNQ5vS8vEkzg0
UGPBM1A3eOX6pmAyuY6P3qWe97TzzbrLFXIgZxnv2WQoyME+jwVDwaKOxwixQMf2g5DerNOoCo5n
RQCX7R6DIeq/Mh52W6otXBx/7pgUydbAqIJao2vOUsdk6TnM98b5egQjVXqCWi5EMbUUu50FN/de
+T/0vvHaYLpKDJ/jO82Qnc1dUlIhSCIZdo2OCcENZbgUB5TLiqvxfCJLr5avJr0UmBTIehse5MCT
Doqc7aoaIVTm3BReyJGUVIAuX5a3Ztaln0+AZ+9yJ2xUzj9om1uy+4kDrPrsHcd6KdB5tSP/EQGo
9pUtK7v/Vd7AKW3AJ+1WHRQL43ML//9v9GEijk1RlFf2QHryTylUdGAov5hMTRk4eRI1bucvlhrN
skaSUNWP+VMaFXAbaVI0EeVXVheZAsuDtRl2iyaMbl/nGse8nadYx3wDm5smUL1Ctx2mEluOzBqQ
J58drS58Je+6o2GVRKW7gm7UhDfPH43JIp3eSipo+TphGcUx0Rco1Em/V/icTY791BQgkzFBMsXc
Y1v+xClnfl38abvJvhy8ELt34WKAwiemWTZ1wRDT7GMdUdT1MxRLiBBvL9WcKGNtbvtEruo5K+Zs
cuERG6xQV+n1iUNUV32DM1Jw74NLTUXqWh4bBLdLgSbM+RytHoymr42xCHBvBB6ZIbes3mu/K7H0
15mPvT+PmO1Ybzj+C46R8BrfqLJE+E6yYMH8BYvsf2PA1BBoFAycFVAiqPaeYLk9mPBruUoNFTk7
9xZpB6EFjUG36pm4hmq7PGOTLbP9tFlhBWbqUdBxkyvUc59SzyL2pyeASm6EGphoEr/7cn3SNy4V
16gF8XzN85wB1MQt6IYCW4xilj04p84lXhs+HFws/1MjgXXaE5dN6dxq3qr2fvBFr7CuoHMjhejS
AhjOyDBiOGDqR/rjvKvER3lc/aEhblH3cygPzoNuElQwYOCw/Z2ORUHiN5UmsY26jpm/Y2iraMMp
gRdyFhtRaNwJzpqcosg6J6P3g2A44hssWB7lY67nImDkejVXb3sLjWG33zv/Nn+esGg4BXrTI1EK
dCT+ZXFtLPoorr+Nl90KYFp+FNHmHqI//8FWUvABhnugIVt04hTtChK2DWJUo+58w3jxuyZmF6Ca
8025PhXhm179Di+BJhDnsvE9Ugy0XQCzZMLWCY/Q6nyal4cHrTtDejR3WQv+B1mBxzT+YgSeqMxn
zO3jkTVjIE9fRvaSzKA8RQ/97O7S5OwMvlZlwmziu43qsjT+NZ84W0jX+EJCOOv1m8qWqdWcm5fP
he/9DiVZZOiFrv7DYC4aNEI4vK+f9p8HKParmFVLJfEIwyHwVGeKHz+ldAhGXHByHNrwEciehCcR
DaRm/mam+s1Y3KVxuzpfhmZbN36PaGT5ELDxvkAsQcNl0oWGEMsCoWWj5TaWxy4+2AbTejC3qnC8
YsYViBlZach0pKbdVmYmDAVtsSMvL76GYV3StmojYJXXKCkWMI9QrN+Q/UFqucil1rrHQ6KU7+9T
oEgx3pvuSsmvOvKR9MB4MpE3J+oXhVywqYop7EPsBqpIIQL6ljPKKzlhKLCW15sJ3syRycaS3iOb
hyl2pyP5ScTSOkh6gw1Abl1KB8j+gXQ9axBB3UMYNgpSRJjs8z6C/vU9sEaqem8RLJHQje20Zklz
1BD7LC0XwSFXPYUeUknhsgc/dalCRWCebZ1hTgEZ5tBmGkHGvt5YrbknVWn83x76kGpTuyR3VHKc
L5WXyOE50xKN0KIXWSh8aLgOl/7QcMEaXzwTFf+OL6QpKrdgRRxgy3Y/Z9C5Vf1eMtgibNmUbvnc
HUkwyCTcxN6n0334KckczTTSPnbexgyAxRvs8blWoDeXUt4quz6SLqOy3+BCzx/5fyF5unXk05mh
4h7jyCvmxEVICfVuB+yvwEEHEVIVO/SGEpxVR+lVlvwpKTjhqEvlK4hjVtfFCgyYlZRXgQJk8kT5
KTrVpSTq7AbHkGTzvFJOaUh7nZfh+3cSp1b/i+OJd221Ej5FnlwZ1OhwyEzieMEAYTSg/nwz1+4C
dwm4d3xTWOSUUtMB64H+SVI18VLZUi6xcy7ZarEeRdsIUa0D7L2wQNoYsGMEP5xi6mLyaONCIPmG
OT5Rzjiunl/0wzVrdZML43VN08s0pscX+HFy+F769C5WFqh7mrYv9y5JlS7xaiQzk2H2k3Z/r/Ok
3Zz27kDFAmntNSgem16X1byo0etkqfOXZS8LXxklBz57pt2OHMO7fRzURzIAE1XQ4JiKj6Yr3PZa
4vVH95MDJqVz8vN3l6UXu2V6EmQac7rRK+/wahpbT2BLafy+hpQ5vrFVg6xg3k7oKZhCU6EUbwKn
pkXahnl5Kydkl+7Sw7JX4OyBxxusZq9eFw4RI2gQu/AksrR3MrN81AQG47tZPJ/VH3gWB/BRnKRF
aDp7yuzAO6tOtIhgc6bcqWse6VauEILrBJHrTY8aqq+MrN23NKlszsE+/7l3HXLTQgoT2Ot4UgcR
o3B3cnTpb+Wi0J/P0qcEYSzipUIj4IdoKjj4PtJD8ALU6ksmCVOq66ZIYgUPzcMMjhDCYyKfozgd
8GFTHu/ybV9pPj0Iyop51n/E9NiikfUDJY1nAWyFVEeSYRRQE1Gv/YaQ7T2TVDD+39lZtRP1R0tv
s+b4AvFzaaPJyRCFoq0hSZTiJ2GMzY+VxrGnV9+Yl8oywEKdPLTcWPgRVmhxcM4/JZ+Wv8wKfImc
58I8pdJ5hp1cCZsRoflzZXwor4whEa86Jdkd8BiIj/zJw/tkKd8TH994fngwPM6If7n6o44PkeNr
7+XaoiIN1A/WBI124i1otzSrcUy23aaKGrgmkecLyHZEajeuUgunrhoXgTDz+2ulJqlXmkeGz+wE
G0Unc/QPfO7g7NpptRTpSYx9TMERH1+0lOB22R2yhp0PbV+L5SS+cnmIJRqdNiYIahxMxRZC1Rqu
m2VeQM+z+oooojXgWoYIlxLpxwWLpHVkTE6OmisfKofyhrMoJzdGuNjOTFOb+e8OsKcB/tC4906X
OwBtIqtUPQAtw5qHJkZLNdIf2mGH2PQwcKosRkU9Sq0HesdEsoOOUu2/jZhsQ+CsjDTTUcPv/8gY
gvrWlZAz1ZCNmo7JavkNih1MlGFgnfpaiUmYdDXYztjPEo9M8O/yzOrlGwqKHKpCzV31vVL41MJ9
GBb3bU611rMZLTzimTWHbX9zixZtAShb2PSzgN4sFU4W8t/UlACIxwvAKaOuE06DqTWn520og4eU
jKaodn5n48vtJtbXbctY/00dwkE9b++AWZrRWXjkfAyrlVAGj2iHDhRBTj318FVw0IOczgBwzAxU
uXcL3l6mxNSy6DZiTbLStjYiPdyFAzMsL0Y405Rfi2y/b3lusSrixYo4NsV3rLYYU4yQ9Vbf9lcc
wlbTvlJmA64pZ8YPwvAtU7U0wDEv5voMNKWh4t55oKIcxlOCcQvjjrekmq9xenXdHjT8k7LlgNqm
OKHrWhHBz6SleYPX6sbX/1Zo11eZY0dFGYWrcG37y/61XPN+2uw87MQPNLxyhs/QfysTS0h4/UWM
F88SPX5+5ot9Dz2CrJCPJ6laoVH+N6Xgimgbopfp5jVSD62BB1VWsqllpxWmtX9LnrHGwEnbItvd
ZSLaPxCYCWFt7gca+rSiXQUbuxlopDzZDOeylR3E9SLc0yDgx+SKtsCjmpmjO0abKnrctC79+tXz
YUhLhhash26cUrnpvMszbgJq0FYZMIo12umMaL0LGmy3c/r7lNCQ87dOjBbRX0vXz5eniyjbOQn0
ngPsQdGPatzZH1+P5jJXojSBOkCBXYatjO207Bf/aLrpcQmUgj1j8tzzQYjPHk3Gr9ysR3UCiTQk
NLLG+dcmi3yjfGy2DqE5BFoUji1eqxnwdamh7NtGpUp8mSJW1JfHOqkPjcGlYssf1fEwd9Oo5jf3
Wb6CqAWlVvHgj8mMUYAZ3vqCfrdBOHJmZhFjLk9HJ4jbyb0C03k6gGIYkYP0O+1mfKDh8S3nHagx
tL/+tXLc8J83L5KP2bhheRD667+/8UMdwak9B5Jv/Nj8K9Gc8kvyDoSZE+LJ1DeSQFuxRdeY00+D
cwLHw6+2bY3aJO4I8q+tPiOl/gJK/O5zTxLdLGFvdZ0bbK9Y4J1ErOGRha7qZgcTAcNvPNmgT5uI
PQsUHrwrfQzJDOh96uTSyMu0qlmLUJfTviSToqkO8tAulwvnk+fS6jnA4j9oGivvLxqlbOQRBCTg
EwKy4FWH9/xH43lwoERHM/RZ+qTrwPh5W4dSAd9GTf7se1+wSy4wqMEFkgrd2mKURy6LwSzs4xuy
yy4qLoZP6cbjc9oPVXhgdqHYnQKTbnfkD4pobBwuEPa+P82wyhc5mzIfFUslEIr3OkLi0d5eUM4s
1K9bSvcIzESU+mbDGEOMFLWwPoTfzPf3cjS9P4b1nTIH8s1rl3DQ73Y3RHgoTqvO/8NxBzYyyX8b
3zlwv4Z7hcrSVsSNCKZgeNM8gdK86JSSBWQvoBLq9dCUquKdxxXTOi3npOm1vUZhCnhbXjrL42WT
QRBkKMStGqsvqwdpUZp6eDBvGDaG+P4/w3kHp0Vx7N1c37DOtC0hAiucQRejuq+F7m9aB3dPgLuc
bj06ypFzGd21af8lPI81odfRFBhiIQe+FFzY4qgacyACfrK5p+IOeG5SPGcGzVUpTtw9kMfE35T6
8Iru7r7MK/hMv0U8+qpcCqY9Pp6jNgDXYservIFF5XEIFTsPFSWbUvr921Z/CyJbif7m2m4ofWUT
i3PwGApwQnaL9OIkn9WOHrOBYLJxM3NyqlF3/ALUIXtPV7kJs9qADhqOGFDF2iBywyyJAYVMaQqq
pElFH+U38BRFnOV9SWHD8alZYNj/BxznsHg1gqxqsZxucXkFJFXFq79WnO74TA46IsKRdhLLMBIS
thEk3kWOLz6ZU+i1rbJiDMqxC/sgGa5fPggFaA96MC9NVjd/DeWU1Zy3o+abGuem+vnLb9vktoGJ
LTQM1cooKMQH9+gQL7MamzsAsrOtqHIVFJGo4xOwAUdyvVJP0iH/OHSCiK9oBx5tq6IzQic1jg5N
zRZueoQu7fTxadmkHZZmEMuaiHeVJMWlhMzkYSx7vtgcmDyQmu6RyN2zR/0XNNWMREwkxOKKtIL0
skYhkFcGTVUdNnsUznDPXTOBNvP6XaqRmHlvnec6Q1HmscwWq4Py75Ocv+qAko9VN5KbZnx4aGNb
i8ccfTn+2TJHHAkVaDWls99lS9920uCHM2n7tWWtXOvnnttnJTxN1Y4ZohTPSlG9JqSHyTTCB7jP
v7Gpg/Sq+dZnybOTKe8EreshxNVA1J6tWiG4YHe60ORxCnFszuJjf3otx7UwRh80JejUrimdWuL0
WXawoumC3528iRlI+Sn0VsWENuHaATqSXE7fyJzDrZ3WQ6G26qVtfSoGDfb4nHuh3s0twXHJtsN0
Fl+RQKwoWoJ/G32WtpZ7zwXRk6I+1smMdnEdvHI6p/O0y8KclzKfzJZCKiUUiynzJzRvt/s+buHs
ESc6TU7WVaIlnZYVHTyaQg0BKQpUq2ALuaDussZv4fMIag5H6IG/INGPE5BURMuOu/wY+hAycpw4
EgJj24ESNuSOAtQ7NKQM9Uhnxw9tct5HEWKmG/444lCSAiZPsyGaHMLnrQb2tKkw00fYhV+W1bkW
nYa35WBI7TIQAxjoivqlLHDMqDfHy7pUTSkqf3lcU4RsM90j5fjl75ARWXQc9oRnjGZg5z0BtlUc
loleyY10lNvlJN4bw3SeU3SFkSKx/6K9UlZLQ2PMmSNlN1Vl59UIagtqFtt92Mv1deKI+y4AvKA4
8ekKoVm8FR1N6/X/deYKRkWnZZROUPz12NVcKntqqQW8v09hQB2oW4JTf6KGGK1CZCEokA3DSYZH
4Zf10eQxFwsAHCppRXDGBN/ThGJkAbsY4KBpq5qSZRjQH7wp2C0Fe03V3nXSoXrrdVLKqkHs6qDL
FlAbTqPYM2DjWAOnnWPRcurn1bjonPMAUa9mi+lXIek7cVit8V89TMa7XDrZ7P6Tp5BVQdrYWAL3
mC6tgyngjgkjgQ8aqLdQElypkaWb4+WC9cGEbMWQgga2/a4jHgFwc/uZUgLfrmWazFXu5TL7HVeX
K8prz3m8P9GBUwjHPc8t3hypd0Jjm2MXUbrBeX3tRy4AIEu5DFZl0OXoPAWvzYGnOEfYyTdl5Km9
BdLoMmE0x22BAymzZniy88GH+kSdLetBJ1BMBnYG13ZF9Ku2X4thC1PMw3GLjoyTQf1KEAaCnwXg
/ImEcNjiGWRs6F6wk+Lmp1F42ttMM0Ct9uZnal6jBG99ynQpWmAodF+tqwyeAyjeYZkrPL3d01jc
kpwC/qogk8tDwpP52idcQiV8YJEM+a4k5ZbZv352OXiB7KNjJaJz+0vnQE83O6KlBMQxOKNsRx4J
odR8ZNKe7ezuT/duocHbFj3wfpmPmF4dSYqUUxN+R9TbG+Nb8t00GeF6k/IiY16j528bAKMPfidd
jFetHUgg92GP1CJ3GsImHwS7fU/Lpy4IdCUz18JofIizudpee3uC6QLrro/0/DYwHJzKzrSB1Xb1
qicTxHaIqEM3MKTPRfacEeVWai3aJCFQDUmzsvP4jZbTeGDTMhlDEYTrvlQjb3Vud4zMYCO5lD6x
tOhe95XMjfQ3lKP3S2hATxAR5pi2J6DCuemJ/QGfbPPPq6aosfaKe7bbvXm8DY1dyXgGKqRCauDf
8bm9fDnGg73zb6ugxMPfnHEMlU18iC8KoqwvIckUJmQWbgIQhPxvyf6Wgi2a36S6MbA0GU5p4ogC
kOxKYHMskXx+81ZH8/meJ8wsnTuRQCaKLRaRTcJ/6u9Z3ELtQnhvbq9tQq+A9cl6Tcix5CIYzrR4
AewmCXoyEMtxXRkWJ2lqJVIAjkecbF4xT2X13gmURAmY1D9lEdtqW8zJZGXD+pcqvZwEH2Kg7mHJ
2GH/rIUE5RaZHeDsWfqzcRMvAF0rYW7FOvDrwPGmIu4urn1vPAw8Ikg5H1tbx0/vIEUPpgiejcfz
GvUwz8sQwx9yTuAvnldr44exzK6+lftnc/yTnzFBdeRw9XGpKBpM/zy8tFdJyTvvyem/OYCxZgu4
H0/odOySKZjjcS8h38wqZPeABgGIQsE9bDBEWBBSh6e42Rcm+hAcyroulZ2Lri2VBsqoE6FAs/yJ
sjx7aUG4q/LM0dXCO93hyyIMVhqqiM5R9ZE8eXi1mELseB8IRxHjyq/Ac02qRw9pZlSUSmakD0Xx
FcPeqwlNpOXHHsNKYWkAdS0qhCcT3g/JsbxgxJ6dK5mEixQMsqth/fjYGCT3nbuZ1kUBsCzbvEJS
lVQvXFIO+qtTi0hm2Y/38Z+rxZJRtUv+U3mrhjQXosahQImdpXpDgWKjRGkQi2Mc1jvlLDXXpIwS
8CDq5Fxzlr1Dz4FfoPp4QD3C/RRLn7fX+1LxyzCcG+Qv6U44NA4Gyplx9X0avGdhSy5ynUZNKQPo
oKCihH6150Ei4uhrHlLYFEwUr1MA18ZPWoCbTPAdwVFCX+BkuJpvAcAPcm53OcOlgmF2IVbUHmkp
10hXDbVnNqQvzSU7PIjNlC0vG0r9zxXKXzUQFkavKAMZwUHm6gFjlktwe3QvhBnPCRMigb8BiEf4
EQdeR2qDLlsYrOSCOF2Pc4HRb3XI5dgZvStbgMWgvlKvs8exXuDIiso6Mpnb/ETux1USRUrnDZo9
I5dJTgjx1pyac3Fytq5R7vYPRwwzvsJKUXKg2hJVzPuq3Z8Q8jW3lCptsoPqPNpTHqJ1tKxjl/9s
H+QGOXRk8DptDistLFcYc4WXKQ+l2xda+UoMo4h1X+LfDjPffeCrF7S3JaFCT9Nt8j98jN31vHjA
UFVsqnsNINVoUDbgST5G1waa2voIXikGnZog+On2iRireB8t/gH2kkmAl25OjlJh8Ybiqf3Fdg5H
uO020CKxurlDMr9owYVYWRoEqnuy8kZC6TMRd/BNsuhRyXJdqW+sfrvUskj4gCgf532FbLt//Ppd
xVgCXps73nbtxPto9WwakK9o1kXA8oe5o4bUwpIfl8ki3ijqswdGuC4kS+2f0mpCvzXflw3IXf73
qvVQPAw9qtiWu0J6fsg80KcdxkoPuR4yqcvg8O0JoEQOF0yl+3/dbGavwRZ0Xj3Bd6XK7zKmTRAe
++2QZmxQJAI2gNRjVBZJK6R6xX7oU1Dkts7gVTe5o943aKguukR7x+qH3bZUpa7t5wvp+Dh2D8+q
jvWqTbp1kMdxl0JGlOqUZfKCfQ+X5ZWqsU8S+de8p9fZCXGu8JoJA/nCuyU2EuvgYnPpk5YtHk+a
p81+fiZu278s+YaP3uqD0eCGZu7VOVYqSHNxrw7TJBcirafrLrikp+6Tf2RorxjW/lWRhY2n24QQ
3r11GuV38Z/kja0Xm39tuDFtthq29pNo7PKCWV5V90vhytduqjFcKJIqL0wT7CbpcvJmp9/BmCfm
3S9xRniGaxoRI9mOkqkcSH9H9UY76lqJB4Ho4m7tTSn+IZs9NK1SNAV/0HE8xmiwbTRWfmlTY5IZ
qgu7NbDtq41001+XyUYhga9LKqd6xSeo8kD+AeLoazURGP3GwHIt7YHZDGaBaNhGLcPH4XUDjJ2n
unU0DoUtXdrqGOhJEqLd39lXYyA/CSVJNdPi9K2awsej0uEOPkHoUIEDb1uU/Jp3IOCYrfwm8toi
E8KIhliMVFIQryzA2mQE+/6V1J+hbsqRw25JKgd5Oc1AhXyT2mI0zUHhyzLS7nimiPm7qTSrN2m+
7oiis/y4CVM7jwF5lxp7vdzYxrt553H6oQk+Ads+bmbTHm5qi0nrR37NBhSgu9aCvQa7hcitIxhj
OlYTJj+MqWeLCtikxHOEDo4H5N/iVxiCcKi4fNkI1wBX86xbFbFaHAPJ4FB7cmFpOW7N/P3Gy7z1
kmhzbS3OZa80K61TJafrXvyaGUrCzyy4NbhkKRVYbMA1XVA9T93cRNR5ian0E6jQop8+ZAhJcEou
Dm6jkuzIR1a/SvAevQ19terH6b3YbUVFl9BiaNH2abzeOqaqD4/q8MxOX3BYNGhFADwmdbtYwt6g
L9vZ0kxYkWKpyIhidQU7MQiTHqkMpR8XKfQljGUhK5vwG31A+s9ptVKYIzOQWhzy//Wb7VFVax8s
YZJo+C5VtmP8xjNQ971+SyhhYlCIlpIrG5gJcBRuDVPLU+nQd1ChGpTudA5/KwNepr3xK+UftfhC
MeHQZL1jFUGLNYchv4FVeyCI/H2KJr2IxBzRuStQVzNPCQVXZyL7c09+G21EZ5NTa4SSMv3zxz7M
RD+MLigl/F5knKPPJ17Pr9P5nmo3UPAS1MAldXxeLDNND33tru0ZX9QTOHfO9y/NNMFPJmqQ87zx
4ZBZX3klOoy9jI0hyuQknkiBb9IJ6iUTVml6y2ecz04UkrtRzNZFIR7JYI4ZIFlhvOfin780fhmZ
ghk6kpYe8Q5PMj+tgfrEkPNbA74SeS6U+0WpFQUi01bnPzVykQphXUxLoPL2Qw5hKI5CZnC0Yucd
ZNjMomwFJDk29E+u51xqh9sH1AHRUNWReCxP5baloB72e0yc7tzjpt/pwPJO7pq4aV4sELqFpRd4
Tv4ec2RxQxfMOnP2FNkUHLP985FD3FuHYHm4dhUHx9yhj8aOp0CvkR2IU3+PnKVdVWruXBwYnS/H
SUiJxkJm0cLYz0UVX0fFUE3GdrYvtLUMeZjg7TmyV/PznX8tqPw0O9ai78f9/NcXjPDcF4Q8Kp1Y
xq7cGyVQXCtFM78TpuMG+a9JABRwlkFE+ITgjzNt4Fpdji/c5yIHg5TWQgKAGPHy/rrhucc+wuU7
v0msQBPat21UGhmrlRemIRf3p4GsDKnTuxQF1JqEbbFpMwkNY7cYwRn1wneD7q8ZZm2F5QLWWg4a
IBUU0GOfBxA2UhJnfqiaDF/R98LnaBxklcKfL/SaBTQ4sLX+CGK3R6BIF9OX/0EB5NusKcBJxIfi
j+zLCXTcHkWnuMP+XJFmyn5KWUrgLYiD1926cuOFVkkvQNZA/kFfSXi251np7CAhl4hPoQAl4LNb
6NkCLiEC66tdsY2gvrhlaJnoxxyZpmXUImCOrEFjm/u1REcU4mFexeern2F1pIQUcZwBVa1FOV+C
PIEM9hI96U9ZlHpzpbICX/RqKfenDLjhJUIX7no/TFsBZHW+yqzJmzE+chD5BnzoZexNbVCwx/2E
BzGnId3ZfU8GYo6GfBos3bNz/G99NYpt/9K7ty/cYrKXmF6klWIXC1IqUSvInburbbM8mRBFHSc9
5LRaArSMuODTlwNP8+FI/dHaD+tU9jakFBmCMRUjTu7ABQaDn4t3wd3Kwx11pOaRClLLUBvQou8f
Wbg96nCbi1hQQnEOaN4h1EipC1fGdW/ApRE/p0PGWOrU60TmvVZimPt5b0lwxlZY7h32lWRdhZBm
cxTMRbTR9qQKKd94xUOvWYrfXTyXbeAq/XuIE1AYkGC5xLn+vVaUrojUZtbaRGbd+kxjiTlxPTAp
fk+4/kYU3NJwyNWkXUTXwPmXW//x51NsEsKHIO7p7Mmlk5g2cxtPUFoTqtdfeU5M+wBAFzKMWaMO
cvt26GGvUHAOWv40CSVVj129+FB6acsH3oMkSmHuZQLaajpxcyCEZAs0D4pmOlpLArirPBWBcC5R
SspIC6U3Y4wPMCahFr8gcga5/ooYSF7NeGLD7oSJXm8AVODOfARx1vOb3kdkRWgr8X3GxhMjHsEL
ufigikk/k0XuIF1F1fuGsPLHrcZIE1g+jRXTkOe6Ef6Jb1+rrKxWeD/e21Tf1LWe76ps/HGpR8Z4
d1copEBjybeYdPRIuenmlr0m8CzUIYxYcECm9jQr+x/8iXw1JUvFUTsb1V8QyHTedvwGzcCyC0JV
p5dI3mJVZdEdkv5h8Yv0oqiJGPopq+NgldWls6Lq40bi+d493bI1COSTh+P8qx2By6/B4zu1KRiG
emRfo27BWl6hsjQ4I0phEpWUtVoHqCn6SwJhPX4e3sjlDvYeXfogdo8lmfpP5kpUUoVQA/8TC56F
LKJ/OpGXR/G8LJqOpHU4KrZvK7LIMEeJBnOTjRuM32e+OR6Khb3R3X3+Jh7bDxCKCvcF/X2LjtdO
VZqyv+MmCxFhPEr1mqqx437CiJbLFYhPzl9EYJwpLuqcMueNRTJRFN98/1FXAqYF9L3w0V1jcswO
vK8ThqoA7a8NXfK2qcj5fyEk/1muJwY6SLDxnNOTmPobTW1pMW/4rPnBfoNasYXgnl48EYlvY7ju
XDFJdUFRrjQdyj7SxdsOznFGX8W7ASZmoekqi2T0y2bkEcuZCaXAZXiSpiR9K7p96aW0e6CFw4PL
QFEH3I6i/KXs4ARpX9cAyV5kP8u/QG0Lb3m1UbgLe68NREjWJglZvg+GrESgmMYIA7MvsIxuGjTC
gL49Mm4Quwb1woXIBWfNLNbcO9ka4oiKr4UOQei9ciImuefmsekN6EdsPai4DQAohySf/qxRTiQn
DhCXyd9C+46fz3mVP1T5t7EEpRp5kF78D3LWMfSHQFPl97+rvIAeaFkb8hdjtaSjnYV+eCNyrGMJ
pNeDchc1x5ZOya9tG8wdGOEhwf6vjoE+fO5g463IubsUYvsTkdAefQTmeFNl1jRE2QcfoAt6bcel
kbSeyTpK9Gov5GGiWQLjSrCCuDA99FTRXRY/g9xt0pJkpPtrz5y21LfnLR8AvOZhzMA9FhmqhrQX
OA3D6eWIsmCwBr46TuQdJ+p3qbyHruTyh8+U9gepudTVnLQiRnvmQ9iH8cE6aI1k+kScUqODudg/
CaoEfmLMD9MCEmZ0u/mspJaI2Bk/fWpsLZndyxa14VUJiTTEaBvBuZ6r+sddHxPYZ0wmqYtePmof
BihI7IRtYwIzzz9I+R3sWvW7WOD/q5KiDxAAWOwlTehvGTJly8k03BLzYjgCwqgWPh/BBcGkljoW
pCz2meBrOyMflyAQomFimPtPYzsbg3ljoK4oY3KVotlxq0pLb07VMVyO3vU/fuDhcBeMEc+tXdQI
PHzL16cY/wdrGIRItY+YRHjCbnJdSHvyZvwI8pcLlvk85gqqVe0wOba9ijISWRjGKia6ZecRlnwO
farEO+v15vXpJ6jEOCwcMokUypB8RCj9zHUdVWNreP0fzKTBukQi3Cg6uzy6zJSUu3ZN6qxsXgz0
YYSRp5qMYhy9Hg3ZVuBWPI114262j9v3TqKlDlNzMhnpdeBXaMe/sAm9zzOX2Xp95NFw+FTcifFC
oRrqOgd0E3iB+aaRJys6dDgqhlNsmqZ/KWAV+ZE+lmb9gOLPNBu2VOUTx1RLH2DwAXVh+fVFm6gT
PoFq0JAvHiZTRGjVfTspYgIdlFwbc3yZfsKyHAeWCtpwtEgTD+wzIZL/HWus7tDAom5gFMSrbqlg
ZD29eX5HvKqpfbWU3RBtLvQ8gT6x91RsZsZQdKa/2uBozAjV+p/oGxPVB02F9nR7F1x0tNCgqqfM
8C//WJLRc6dYoizuOgPBy6Vbnu4VY+HKPQLC1O4mhW8y7ZwvfF+nMx8PDWpKpnQPZ5mR9/Boa9gb
lN+bp8YSbavoF9sdxdjantWdmu8vgleyS4rY82mky1x9rpGVzHpLb9FTqy2oNBqr7vgtKThfVZA6
nMUw6y/qVpTzrmGvE5HLYje+1bA+6Zp40gJSWjcviEWzQ0XQ5rKfVDw5jW9UeHHMMY5zbP9TE3Xf
XCk9sjk20ZfpMVSGqJicylUYi7rUDqF6fZCcK52tHsCHy4F9OPl2SUWPfaJtXyEmBaQeFOG8RajN
LKmxnRT7ybLyFhD4atkxL+Qnvn7hu8igiq2R8ohMWPR7UWcRg9t5TwBHSJl5oVdeSz60wWPfG+u0
UAIiHWis3/Pi6jqWhiZq6WJaaP6Y68o/k3XW0P+mElQNgKpTdidsek5eIJjPXCdb52/U1NhGecM0
Lbu3r6KFKL98CpSFcH3IZrO24C+ciCxoa24mQWtFdA0WNn0aO9sw/52qprbQPYgc2M8B64JHn74u
B/Gikly6nxhcZ4qostXlOsOwqHu9Wju6lFiM/vzOAc2L85tykYye8om4B0vmtowGirwYaefQ4WJm
xPJ7pGEIxDDs0JI1sAB4JruTNp88RxR1A6xHGw1V7htD0rZ9Y7VRqtN6J7ullwY6Vk33r1XhHw2D
OTAwjGCI0fjxV43IvHcplnnycOKI0IUD2B4AG9/WsjxbWkKx5Eke31EzC4ZInr0KZVC8IsY5vULF
3HzQvr3KWLLwaWXQNrEbHEovxUBZ6do8JCGN2rGOUcCO7jvn4tPRvQy0Sk5LsAONj0tW57yEu6aS
P4kJNJmqtcgOMp/4QRXPBX6jGk8A0SP/BRQ6k7SPCTkHzA6lPlHByqypVTonVCwl6Gx+17ebdIqL
wHbjVTZe02I02Mu3Utp30p7Soz0pIz2TGDCJrcNtwusLwIePPu8EgHA7R/XNiLH/eGQ70DUu+7ga
PEQWbG0jrMIztYtUKBrzqrP5Zg0Rf0dGHAgHlUrHlcq9t6N4QkyMCBNxSefmLT28+IgGBjzaTfNh
J64Sh3ajT955gwez5bDvw/gqa5h7qPjLxczWEiCc9zBZm2jEe96zXMR6zx54A7o0Rv1JlSoFfq0R
h6t3+DCG/MKaIwYDAG7sQR6Fbj0aWgVTVk10nYMTSltnW8ASjgFaRQwAB+r/gXm+Ji8LW8BKHrtv
KfSx40hhyaLq1zqWGVUdjDLkRZNB62Fku759lPHNwKbDjxU6umoHlU5Sn6gNP2Orm+oxzDMcWNQv
STo4q4crk8TdHBgmKX9j8rzxyOdbAaJxhuTjYRQYubv08z9m9pXLr4iLdBlIfuTPaTZUa7dmkT4t
ffmIW6iuY2lZyMGAC6CjvDHMUlbmOK+4bo71n1gh2kvQuDe3sgUiRuAsMN/tXvbxlANpPWavmGnG
b4Ckbd8TALx8v7zQsBkebe6uVkcTc3nsd911tqcRtraSsHtIR18MFeT/2eMUew9/lG8KTRNGP38K
2XdeWPc75fgNVNyViPhpSNkMIvhwnO4f7W2hRVBtp9eSht8DnEsvuKQDXnN62QSoJBYWcckkQx67
a7Q7v7mfeXDLg+COK+cEux4k5zErj5XTtgs5FQ0DTEDq3SntzuX65cZpnRdGDNyDOIJrwoKtTnX4
v16TuLiHftmTrj6OK14eUbMouX8VawjlMR1tXu3gFErBo0RhurtYzw4HpabK9h7cvijUuSZrObxl
WVz1xNfHHBeRiOLXki0cA0aIeo3LQYTGRjE+NsJPVs+UDt9Sgn2J2YKJ592Tm3b1DsNdZBOEbdEr
HWhuTHinDxvICSyxWQz5pNI2dkRW7h71f8Hxv4lRSWHGDghHm8niVk0DqwD+q3GzR5Tfzg59g72f
xun/Q987lSxqgd8iV7uk25/VkZwj7Ag8Q+g4iixd4yUKdarVHbeIyV6vaZwqgDXYpdoteG31uBsb
BDxkRcE1SqJCRSrNbv6Xac1eFmUjxMrQ537GBltNnmVd6PecdW5/tv6m8IG3Ywz7cWXYAYGelofH
6nj0oXyiH1taMp9Nicy7TI+LuC9f4ZglR12dz7PERFHtsMxaXLLirXs2wxHyI+/VD2Qu20koVbt6
goMonuMFlOisZcIPuQHkaWAynYFzlW3w/MWMDwk6YVVQ/0iwOV6FW7QCtFD5qfYATbpO+k4dXLSO
fMdo2lGCrRxlcKlvsJCobkxDJpXrS6EUhLUtYwrKmsdIb6ME1UkxKaAn0U0d9jl76ClIJDcdAABW
lB3kfdsJVrlkXw/Qw1pMbeSqEEhBhXr1Vw3KTULARdcvK6u4XEH84S5Dsc0xTjinYiZZzaeIE7ve
FWODpVx2BL1XruUbE73Cvy2UAOIOz822uuhvXliSXxzqz1jWjIgjbikqIdiF42EQWWtw2ZpMmH6i
jwn9BVPZ4XItB05/tWGip20bBHriZ80+OsxMkiCL6L1A2cx+siFl2gdoKN8v72X8+XL/EIhvyFHT
QTvMHvZjEMFJyIvza9aDNy0SQSwdnYNZQHLJJZnPB/q+H/7zVzaof5MJbMwhWHRtEC+MVb8fziqZ
qFTFhyCJ7iswqbJVymt/rB3pEVr0rDsS0vzZbT7u+qGIjehXGMJMQb8x2PVAK10SqW2D7pt7Futu
5MqhucwP7IIH6i1TgRy5mJW03jwt68t+2ItWjQt5pq+pLL7uk4jjJzpJf8LWuREspkaCNQ50FHL7
p0bsSf6IocoS+Mewhwry3ZHXrK0tplO5e/KbdRr5RplarCAQcSDET2qlsg45wEnX2Hu1qCwWCZKt
eDZNQN0M1bFDGtLqW7Q1/QLEaEhJSu9luZy6/vXkWTPgsVWu7P+Gxo0UEvFwPqCHg2VC/LvoLYyb
mwS2HfHXX1j0nb2E0lPnKbCv6cK77CjBwyMuwwYtqhDhN9InYQ+jWeBX75VhbQ5oHTMdV6aJu2uH
+p0RfJ994IUXhlKXREZjSMRp/HIxdHlSVw2MhtGGKQLEuA79rlP5APguieIlWyYgy9ewMwGX76Tq
/zRXCGZ/VNaJYEP9qnELtTxKkX/4wLCabb5XCHhee6Cl8VviYcLaAxFNy7MHKelDdLk+/+bVN07A
7N/FJmnwLTtkn/JmIJ1egknNeFFyY+cYx/aQ7/MIWqZPLq1Oked2U0Q50Y2c8joRfoVbyWrx1kpC
j+9dTRd3J4fk81DafFgSlZn9zJFy0ZaWBgr68OnGPyIAtKV9hMQjULAAjFwBtlJTQxG1mKqNSL/x
Dn8Dq8lj+c0ThO9m3Jql8cEmY5+rnqf8uxDfRNjc2OKbuMpJjmjN8FQcattLniQ1ZpnMPxZU89Dv
oJRUEuHBwcnWpObj/BpDkd59oV0COtVZyE/D7GWGd2BLIQh7B83kKpw9sfNP5YZyLqoFKgFIZvZW
oQLy/UZo3kcx8FsRWoftuQDwygx4AqCxL+DREsRbX2d9y/2HaSqojYeFtkSsJhvEOYn+Pn+xeWUg
6V1mj1KGqF8W+KQwo2P9z3WSGh90WD07NAPBonhBPL8RAo8KN8XDiyrFA51X3uBVZ8o8o4SskR/z
54tLn6J/TfgaYtLguTwHKtYBc9BGEIznYAq4YdevruVRz1HWfu59JtDEoQqG+S+u10qoWMr+BPjn
Bd9E87qRVJplQbu/luax0XfnrjmXHLnys3otNC0rEzF4C1PQHUPBQG5vygmczMXVfA9x9XIeKg+b
Dje5Lt7k0V7I2RI/tZXMjlq0cdN93VSwcSsQV2cJgpnWYPNOXwZ+NaUs2xYjRjdcvjF3Bi5VHrdf
3m8BKt9hS4G/dPjZFzp4v9fbbJgJmNQ6b8KWDGqdwusJGa3TGoYGvadiuhbe25+PTh03TrlLEuKy
S4Brf5z3qB3v2TtFzB+P2MaaN19mrYAlpk4BEtiCLwnDgJ97jICerGSj/jp2J1A7UlyV7T7pxHOW
3g6tnV3YmPvxDJo286/dKmSa1AzzEskl6+9uEMMH0oBRmoBJS7h73sYajumFLNR8z0B83UCLRNJa
PYf+nKR2QDPwkJQEfOeed5qFmytfzCDuegaBJDQuLPNVnqzJIphQ1oIQUasdTpF+nN7CHFf71xyo
SnWYX9kwOlY9fbc8bFzBEt6jdQ9m3+bGeKT+o7L6THDhdSHEpP2uaCvlNRms9j9aGmDI3o4ICVCa
inrBOXo28MNaOSniLGOE5VoBMgKn1cxj/+Pv26JgLhqmH7fODg3FkDQLnDUBLGEyjIUYhJe1hVrm
EBpS0sScT6zzi2oycxfC0kb1mE1GosI9zDG8hOplhbS5y+l2KsYPBZwWz+mY8OsWEZ4Tiitf9/L3
jIA87w17HcOIkIHJnG64nwOxnfnhn1aDj89WBaHQDN1UTtUrlJiCCqF7IaMz0Mns0a8dES4IZ21F
2nB7KfliRUYQQnG9Y+34HTxCDaeogtzHh90nSaZfmFKjGqnhSEvLV+mDOoFvG5wHbK5UhiUJHZQh
1ZHOZUy7AguyP/XfjAPi4ulxr93m2iElUaa39dgF2Qu+IedT+m5aL9XvnLeMbpF3Qz7SvFt/7Tml
6ouP+Wit36ocxTG5OIyTw23IpCK/LPLsPXd9JJu1I6MonNCFsVXWbRIz/lVGWll2Ib+ib0oyAkhX
MTBHnekY0JBmH09ERZPZzEP5OmVztuKAZQCTaT9zr7m4haLHoeaJa8SMqQ6kc2F4qkYEre79PsRv
ZCH09StLuq28K62LL7ToQsxYlHvvBcptBFhmR4tddTnq7nm4ABXPw9mlYlpkXbKp09eKhzJrP4HV
FtbETCl2EDMr2v6PdmCnOfpUB+BlzD97H8wKbfqw8Fy6tHUDrgpNg9ckWlU0BreBsBdv6cSgDMvE
f255d5peJfEgqlKF5Wl3Y4j/J7owPUX3jbjYSuonZzXTivAWRuYYwufaqE7Nu26pCRUvvkZihDWC
FPhIptjRw2d0PHYLY2a2h3efWwCBPKtQxQPGVRsF5WMxgKgpgV8MgjeHFxxzsF7Xia9JNAzqR1w1
9IX6KPNzB/fPYdlP+3DxmmwLZdhHU+BkwU/m5+mH1ef6bnHVxN/q7r/yJpcPOd8Twi0Y8dqIqSty
oe38boZdgnuqXVDPGFOjAeTEP5vkG7cFkdbMrh09aMmoJIqeUVC5DApsrJY+ViQ8K65XWNCk19jO
FSA6NQBYE1muBiXSGilK0NktOdT8cq0LjypbCJRXAN8kpcxnaba9PBiuc3XCmHt6JwKigdxQbxII
H5K1itr5a4FNHJJMkk//kdyImC8+BgTFU2sOOJh8TIbM9Dm82Zw3UZElgKyaywahfk8KJC49Tg6+
LleLl1aV7bB/B3YXq8czX39SnU2U+93K0Gs1oV8ExYup4HD7eUjL8U4bA0/1o/6ihkjg/iyLIoYh
+huYcoLPvGUUwKfkQ73ZFU8tsu1Lgc40Vthulps0BYtzwup9SwUhAGug7hjzDJVOH8cN0HlWWzZ6
cHKdBlvITk3CuaFEQA00GJra37MLf3x0lGK3aQZuz/Gybww0kTXmvDTFL0ouScwS4ehLKnSxsgA3
A8iHNwa2ZFPfytzBNXWx8AiQk8eC+MXOMa1G1TsEuSsZ4Zg8vpvO+Fflq3jGbjGENMxqoT7QnDQM
l7LFVT++E+qgzdT1yWSEYR/2HUGPFKK8ZvFSwOg9zkQAE35YLk81+5MSlnUIJMRVNc9c71OO153C
SKzNx6eh/PREFusH+we7um4gUvrLD5hzaa1PAQGwFw7Y73qwx11ZAmzMkSa+7kLmaMKxXicAtcRl
7YFdNEkcCopG8/AzlUP9wIisWkTNrRgenut2m5MhpHc3HmLdxpR816DHR5elzz7+gduE2N9mVllg
bx/g0pMZcCqQDX1zq2cQVA7C5PcL+t4t2hjtNFGQWRgQb72feMQFlsMCF/hd7+PIF5wSwroMetyt
fcmU9cpCfdJpMkOrZac4m/EROkCRKJPHaHwKgAARRezfalU3nWrzLpX177uuzEFY1Kkbxy22Pefp
DFoGC/a8RYreWD5v6z3k6YgZHbnn41WeHlMymp5wea7zpoZcdrid4U6FIPUTYOAoI25UM2/EGt2+
BfqmvtIF+gsq5Ts6hbwqBvyPYKjYJ55eaCvF4tAPhOSXNHzC6fuWPvZyKjbpm608rLW5sc0mrfSq
BUSbDwFrpDmvOa4dfMY+iAYUFisRCGdhIi1azkIZFc40SuxPvU/Of991TDliVVdyHZN13WsAOaq4
5DmTTLrYuigLX9MzXdJBS0V/4Hvwa2QHit2V9GjvULFr+MMxTHRwYNSK2tnVvP6ZOLWdBe27+jcX
5WKeJPi/gi+YIdOYbRhw1Am8RdBgb9D622YIii0yiOyliBsgIGpYq571D4G6DE5w39aPosyDHTk/
/GvQr2tUc7bIrkX5SHwWngB7JJy4odEedzY2tDyYBhf4LEz4BOMDy0DfcxWIdqJ3DJ9kTLkRO9le
4XmHF61A3wDJQIdwlTX7KFTo7FCtVqDxnppAn6YYpWwC0FaXW8dMpp4JTCR03uR9OOgQ8EGalhIt
Ca0qxxgiYr/0eQW6ZgYNjXPc60ie2vsbxX/OSzVL+ETjz8L8anmcKxOxVXlxX9hk+7Bz8nUaRW2a
G9422rni1cBfkuU7x+2CZMcexTs7mxkwYtrqngrpKqEBxe/2OM0MdyXO+/EzqHK9+5aIaY+0iZ0F
bjnJ13DFk9+orhKCHLfstBjo8cOvcJ9xPhOmurkT01qO4kASqZtcplj3z/yhuo5kYb3IiKucS5ki
qF1VneN8fhMNE2N6ATwWFDmJDDPGYLuZggYcElqjx5Zy6WvnU2sanhSu5YJkhCSK72ic6pjct9Bw
2Oa5J5eQ0HPixi/7b2uHcbRz1+atGBnR3jwifvN7OXir35SPT/MxrTnPfqo22q0aXmb6jGQ4947Y
lVsnHwo2SVo+P/C0W+F8OulQlbefP4UND5VdElao4lbbGfadfgaqJDan0bgB9/++6X2t+End1Vgj
vKw310aTTxe0pO6H66k3cXgFRVQreK/5MFg8SDv102xrqlUz55a+ssbs1u4lipmm/Obznn/9wjBj
B8Vf+vlBjajBmqYrvQAv+4SvVisuuS6qoE+N6RE9m1OcWxBNCQR0sK+m7Qk5iASaVGJvb80stjOT
tmBRoEIknIMz/kO+IGxbqZzWszeE45QqlPXwNbfz83+dDF9wEFqPVW+vKIqn/7TxXlU3Wj2fcgPj
So5p2I8gYto4Eo9YGjhGVgNGilPuctlEUFI4sOVV3tAjQQpU9xz1qcm4IyZIAlotCplUGsIBpzgt
3ORght6qoUg+l5kdwkjQd8iVm7KX4jvFBF+CxPgrB74q7ksDFDje9+j2fn1vCRj7KTJClLyWLOo8
nizNnP7vdOgmkXQFjt+HnuffTcS/SVzRKp5leQkJKzXiBA+sJEpLsFxLkppgdI47i/I5vG+XskqK
3kEOPWMAai5wZ+K8M4Ygx51Rpr5qaYytn3GD4G4j3xHwTcrdZODMyMWOiznkHI65i95BU9zms+NH
jwzdDGaqNF6pomS/Q+DupdqMPQI3FI/BGaiBdUmTNuGgDuegKiqYmpq4fY2/OMS47BJwsbVuXbo/
Lsxr8u4y5SmsPju/le6kuXB++BkqPv/Erkyz/kdJvnd3iH6CNLKCf9T3FsH94KUVDCMVw5SGmsV6
gErtiGQUCJgGpC534lOTmPfns96TmD0OoNvqkz9BlhJIxOyT7UOVhbDm8r/5S/DATltcLNfQrb9m
jwSXX3w2KInzWOzgfM5GBS0RnDeDuwzOv+AcbDMRLBGhVkj19wSRmyzTyCZRW86fpCADl/y6aDzy
c6A8jWRKM2tqDTEkgCf5Fvn96f7JSLUyPTeTxomUnyDZMmx/bzOo1srMAWTIru6CJX31EPKwdH0M
t/ZUywNYTxqPJva8HMKJcKDFPdjNdyeN2x5PJir7+FBt8tLlzQsUJ032KSGsOZaVFg5E5/HNcMwA
j8qFFiY7NYkzsgiB7AeFaysb6JF1wDZSqvHai9eYpnYS79OFw667ylqM4+jpZj+4sYaTBqMYrUFi
f4Ehi/M5TeeAJmo463y2jN/BBAJmm7l6LSnEWMk/3DgbV4/jIHHhBeBWILlQqeJKjhROxnxZ49WC
OWUSpjTq1e5kRC/cO4dzerWp6pk33Lh/YqOQUFkkV3ibuRhgGK5KY2tUCkARfEJ9WB7oXUiJP0MW
bmQwDlS0b7+a1j8/oIkQ2qnMhIZrMSgkcvmDR51Z499eLKP3wl8o4oPy+6W44e0HfbpEvsa7Xn3Q
2RTI2PYP6xQY8Hfe3tb9Wryr/OrzBDa1Y/5J55irswH8WBure6u8b5e8G0IuAmJNY4GpzMFbl3bC
D+7fMakNGIehZE6vPrDif0Lwdq/OGNDdtsqRVDcsT+dYuOfao+3NfVHsbYcr9IDlsldttzv/jFa5
6VR9ryPKByhqZwQvReWqo/CWa+fcCgDjfA3gyJJqzoL63+GhUk3zr7F4THYOi5KzcJ/OtOPv1IsZ
hSLHa7Uf7t+3JO+XfAuiRTjpWp6I9EsjliBWYUimysQ9Uei7/JzGXMyLS0Ep2RNkcjmRpMAmf0J7
oIzpdGlW0LZnU7YnR4DYEsfxKigFyqpeQjqyOxg7Bbet6/Hs+OrHg86dvAmW8QKTBLKP5GfjHsst
FPnvDkKURZ++WzAjpIFYFaPNA10AnqOB5S42djzgc6bH9fm3a7TVkilw6l7ITc2GwETg7x1tlTQe
UUyMu7ondaMhb1f+5cmiCaDEcPMpCAp6iJ6sK6s6cxHkmzSD6H5J3f+LqzFQow1ymX1zBuW/USl2
m6xYlHCJLhcdY1Nizf5YDZ6KVMIVfvSrLs50+DhaXTArJ+GyWKJUatLOrfMsu+65ivLIIzFGY4w0
/462U1PoAdYrrElbrPz+QEfS1UpzFl4U5Rxx0X++RWfF9S/tXMmcfmCV9tN+LH1zg1uQ43YPGvin
EGcaguMDBjfxT6hsFeMJjVFPaMw0TShynBRIYMCVpJOgKZjP5nW5p4aOS9G6sO0A+xsk0NTuA8c5
+bOfnSS3rUg+YY3LO++++iMNUXESNWk+5VF7Lip/U9p0kBBNVaX56fLc6ruQnLYp+0Da1U5tnE2b
DMXw3YkSamOtb39hB0wtnLUgXYuRR1x8myfLiDRB+meQTU0tzu4zedTpsNkLpaDpEXcggQr1hVCf
GOQkBsssfSEtNyK6ySqG+vacp8UFR/koX/QFlbS+ogC1hFwqsk6usH0TthssQuFCRdB2S1AboF7m
qUMfddocPmZtssRbVhyDjQrfo6b6mYuJ8/aAaAQkKYHk3/GjTxeV4KhYcvIeOZh/9y7Enh2OYlmZ
61zHAs6PMXuVmYGrJVq16fOA9gZY/++SE3t1HHczuOu9todNcg+OlAezATObhTvLjtYTgY60xeSy
zjFzTjpD4Gj3u66FlkaD6EPe/Bb91BHk4QfZwPc+QjudgXenr4l+inJeu7eVDNufbhUsxoxz9M3h
vUKy3K9ngXUFXEige8cwkFmR3dLKVJcOcrA7hriuKnyFk85rMSLr8czt5DbRBPAztJy6rO68axEP
KfqOpZAbSMi+4js99nWupdifL2US3zSccg2qehhqGoPtjQE4Tic1jhsuXvQVPDzLKZX5+gO7EPf5
4XTrKIUdFtdGDychveHVvfuLUijHvM2N8fzD+oD6p+zSAwQbL75ioNNkk86I52r4TkC09hrQzidT
roHD9gJz+JUZwIiHSZLoMirODfBU+ibPgQErXw5AKzK5KI0jDlFs1z6xf2SvFXGVIQqN7moc6IWh
dqMMeb2n6M+esN/Q5qpaTNaH+3iP3on1RbTLThzo9m9NSw5+X9i1b3h3pcJgk3LOt8/l5lizLExF
wK5HHvZuaqkkHeLF8IHdLHHLYfsd2hHt4aeT/4w7fCypXCt3ldOxeUGnUq3LyPnPxkZ8eeWSy9b6
1xQvJj3tysAl3zpEWpbxk6DgZjo8vHqZnWJNfbbGsYHVt6ZE17oe8kYLYGNTdWcqhzPUfj96KCdw
2Mqfod6MvItGxy13pSxd5NwgZ3Ae8D2BuP2bicrb8GGIQsHQ/AhsIYrPA+g+srgEEksQvkqQb9kT
dITAS7i6wAvIP61rBHX3ODKba+9ZqUmwOYcZkhsz9XUhp+Mp20NoZxeAAZyzgAkmdMoPJ00oH65w
j2UGeRj9+8vQ7C3ocYUv3IZti3q53NV3Fj10hUPNQsRQErUMZVQUR79iVtKHOV+WThx3hsYH/sSa
0xyEnbGxOBqIr8AIKWZQj0qfNF9Wk93HQ9t6puwAAaT9WzYPGBX3XnzXMbL8tfE9cZPsbiUbh+Ru
jOFxN48Ns3dBsMvWzs9MKoLRvWFJJax4FAam5mP1+UZ2ASbWlHUus38IyGMMz5EfC9WoQ1BV5hFb
ICbnl01A3NJBK3TO9CnUQGXNpXhpAxizchJBNP88RTJpSgX5Xs+cUX1BIH6bl5jMSSnJYYV+ldxP
3GvCuNdqTNb9RLUT4ZAjN79A9ze+ysupw1mUNHIf9FEHi0NjH5HxsfoI/I/UBEwzSf7H+39W9Fvx
OiWZlxBvkVOHW9uMJHjj8u702kLXguBuKp5xKvCo2iNiOSiWrQRJ43dNrKHUMgKtBWN0gQzlzCy7
sv9QF2YiVlUCZKOUsOQiZa21qvpYjDr4dw9FoAYVXD/Qt9dHPCKYzvp3W38lZmeM8bAmb69wd29C
EN0M+2URywqvQ69lfp8C7McsdOx1urDsm/ui/iN0c0eGmyf+7OOIFYKbimUZP8UN9Bui8CnBZ+zm
U0AwA2bTCaGzVxE0ku+w0iBtM8wnZ9H8G4qCWj88oTD5O1d9mcFfGlWEM6iuUbhKOK8hYJy4xngR
h0pr86PHelp1OpqDbjHPNrfZB0uGx2i0B2fZyZQQcieVVQiUfqLQyekWFdU7ZWOjGyttMLzIPMAi
lWnilyzEJn4sxpZLiJZBY9cyMdn52IQQGOvr9v2woSRqNNkELEUT/lTXTxiouqaxLCQgoQkhwpnv
n66FGCHCLaMGzaZ+BliZytg+5n4FplBdpwqSq16qW1MFXdsRe9NP33/gsqL0a7mOYfztcpiXsk5x
UWUc1IRHvU6ZOJqBWvKwdRJeZCKBevzkc2bti+TIJZIcAIbqPDPqtVGBT+RibGewnrp0mB/p1ADi
OJwThI92Z7VhYaAtqMP7n6eVUb06kPZY91X3j6nBdXS30e1ycUQ6jh9HXhb/GxDr2JuaGEQ37p19
t5ij92OeGgJxF8FcgycYIA60/G+N2XN0JlwrqIQEChQnvNPxqB/Udzdssa40uHea8FtpDQ7MyUFM
RKAM1zCkkACYRkq2+okvaScVSLIHjDauJJNfWYygGyiqDh1wTC5H+UpnKQExC5O5CyzXbBgu4+gh
R1WztU6fqQ3WTH8JJXnu1IpmAmCJ2r9RdNYuHBncTM/m292J4Wi0dD4YJDD8/0j/ohUnrkPJ84Aq
1MS1sTjilgvCiGlbUrHaBkmw6rzc1YSkDb0E6H61jpslUODKNdrdkWBU3Pfyhx0/Mn1uYY/M4Orn
C3FfDB1ewjT83GPGz6N8kx/97l/yGnFVvfDCFhRVBiP+d+7sDAh6Suu++095M7ouE0rUdzVABQEH
5PQ7Y7f0O9Y4TvlQ2Z5Gz6cbF4Nr/3vklmV9pxf4HLAdGcLV8nbazSTi/iUB72C8so/bztdphkYf
DG92NAuQbXFkZxMIk2YnLU0Iyafcm/F87gajwUiUe2w0e+ogs+riZTofi79UFbbCAPGg7vNB92KF
0FuGoDQyq/u7p8aj5W+umWV3nSUssf8tzLhAPEr3oJj1Tbe0IQvXcFlPl7XH1kWibs1xEtBrBkEa
cRGF3BRgk0Ecim4p6oSYFa3+FuZy74+48az/Xo1kjHVa62N+898uMrNI+rtHoP6JKByqqcPPREHs
D+lmMhopUrjuDxhaAIJt29Q+Hsp5eBJ+0aAUZHl2WsDZ/FC6OAUeChT93bkcbny3jpHXodMmW0S8
ezu6B8n343n/BUfq4Pu9ADmA0HwCyRpYHHmZhC7Hlk6OHdgY/HlSwyZYnRGMRPPj0nhxaQwIBcKK
lolW5bVoyBuU3S/nnJTKsMKFLVUC/ky9oeeDrqod8HFw9AE1LureOJO3Nq4UOGsXfCrLF7K13uhk
BOF1Ur0X/9lZaef9APBQLBqCzlofLmO/Dqd0Ux15oeHuhBjZhILkMiYRxyKe3U6B1FUG3g3/+uyj
3EB8YxLe+OKVgKFBGT0ArNuJ0fvMOz+U/NgivL+H2slXHv6m1CiGxcTEiLYabBpgcgMhZE1HiSET
966MokFTmj8QXM5pJIc+NSsgTvulIT3G1Cnva0e3zwDJ8WkhA96A9CRjKgLnb7UJohEWks9mT2sr
MKhSH+Hp7WGqdI3et8oWWBgTVXkcAY9lrF1p0htUdpZhQj3CfkmfL9QzM3lbUa+V0FAUxPOjmXR1
QWFDYAV2JjrKiJ4ZX8tMQB61ZODY8QiVsAE8mlOsujCm0JPuviQbdJTzayBhfIITB/aNsJ91GZDa
08XQFPRXU9Y7rdwWmx2qnplwLPmG8wg9MoLLFbynlWeTKkDLrgQukwBoeDPOVJ/3V8UR+5Gmav/4
9ZbIVHzwKzQfy8EspJAG+xTsqL/jdOf1EwEDejeoqM7monmdJUHpZVRW3OoSkKlGZtMjPVHijG1B
fzeHrct6xjRqqafsmFP7NY7ZY50TLSNq1PPon9oSzGkmOHRkgvyh1+zydSKGaRIRLCjX4Rtm4t6i
4JoLLlHranmd09EGiLiLfH74IjmXAUSSNC6yTyOwG4yEpbCuJCShQX+gQdYxUBArGvRtNll/Wi7j
UH3sf96G58slUIkD20YAtOqUDbrgmGItiIgP13ByJzAn92d//Kry7RIcD6hqVYHx7trxjeg6zw0X
kMPUznNPcrYTXkQtzlAOPfb04hL9S0xPO6HrTXr9VFY5wJuasHJxFMuoVJ5CC+Z+IXarpCeDHpUB
Fj5r8SQEBzFMjTcumPLdLwziQs0Wp594cpatyskU18KX5reeCH8uzdR2WVwQakXWJXYjAQhidavQ
IsbTb5V4V5/abdTus9YhPYGzmIx1u47Fo9mR/KbfqlYraDFSVFJilv6wB/OoHT3DpeLZgklaB5nf
glodkle8RijsavzO0Dyr8bqDQwWOE/cVpW8buHtiFykGC20KM7QoxOG30Eum+Y9DpXes4MDK5oV7
SPznZ3/O7HCpNa8XTKjZOGMYJFdP2gLnW5dDd1IrIWGVKa950X1rwxV6kQm/kINheq10yM1IxgSR
quU2SqylhvKUPTc6F626/ubQt6MY/fVF1G9GQlhxbiWpK360PhH00L3q219RbNMSofr2wrvAqpD0
h3qbJB+z7SRkcVY/qYct4qiwPD7nDa7zGTDnRsgUH+g6zB82TcOOJFOUUdkZwd8NlXejFQFQWMar
WybtG4pC5+fx7WfOt0Q5HAW3q/vaRAKXOJQSL6z+uMdexDKkfpKYWOf+uSK8B5cw74ooT0NhzpTb
s5O1g/cVjE7q2Xhr+1iyVAV86/Yr/clTbc6kZsA8Ju7XN0GV5j/p4cKQHxY3aOSbFMEznMsyw3xc
6gR+b8DTqoI9OUgbGOXJLqEMU/cES81JJUivIvqpEubO5pHjtIlTX34WBQRpmyMXbuctBLfD0alf
VYs6qO+A6RVMwYVgeASAmxGjNsws6Rct9XQpMRjafVFq21LEtxLpa8aN0isPiMe3DW51WuSBjOKl
0pJsnqHWz/SkpekTYeWGbiNO2cPRVfhDVw87QRfsldE2S770WjmFe428xf3KZRxjfBvDd3ifaXDs
AwdUC43jdxnSNKdc8c+e9b3ymtWwRYLob3nMPOJYFewyOjfZcI51QfY+C/Jmb7qKKS74zNBMcwMr
dNq6eLIA6tZKLjJD/0TrN3C5AatH23a27wy3gUUv9RcnJdkzv2IvGQfLcrSwbvh9aNanrj9EUi5i
AqYvNORXbCKynVzrKqtG3qPLrMd4tZNFmmEFB+srDRwggnW9wVLjZOlZ7mikb5Sgkiajtq8QcC97
upQlJijBw2v+IDTYMIjld9kzHjYk6WTbeeMP2l3VapQiIERf+180Cu4Y5wzKZURIszy+C8mgWhVk
Zd19M/R4NBFifZ0vbSM5J4ZPut+7HBsMa1Z3f3ULpgvaeLmkuR5hneIdilj6hs0oAB8XY+ZTR5bX
dtjomgp2Gyd9MqtfJyKJhS2WXmB2/INmQEVmCoKszQOVw8mIH9TPDx5pHCc49kJKk3Vhhk0GoFE2
hnB80YrfvZ7kyUl+Ppi96otwvt5h0/V03TdD0TE7WtjfjQUFO+W+T5i1Ob51a46KaFULMMBqt+jz
5Pot+IP+4S4qmzn445X+bgF0jXbOizitnZRC4pn7XZF3JH4kWEsPh6zXDwNVaiGD+vsjn+tHjkHW
lnT6zoGE2xNiUEueCdjwNvPOuPM9oGtH5XNbhUmL0bpixoTwprnaarMZWonc4todx6GhES65J7HL
TxLya6RtaH5gOF/Anh6eMQkFWK2WCsHxfEVvDzKr+U4QOrQ5irebi/7xaNj8qpe/vlm+S54KZ2qT
IZOUvEgeabH24plf/lE5wzFAaep7WCh92go1FJQdM7WEu+bjWn20JWl4Y5PXBHJBSPVS+wfw4W/o
tORnUqualOLw+4g1hjC8fSDA9+6TwHbMiPWhzcLJGC9Hq5ICpXT54OJFqUNORBrutXHA7r8LvDfY
UE8JV1vadUug5GSk92xPGU1ACOrjO4grcQsPHPc8gLg1WZPwlIpjAlwFJlXqqkKwogYEDtDV3PCg
CZamSKjo6hkTfy/9e5kuZeZy7ARItxllxQodToHHc+1JwgSQ76iBfNDQ2GdGxaR4xw5rUm7Fj/4+
upB5GvzjvLvjQTv8YGrSfpQBTPCUl+4g+BqY8PHdU/q7Z0RNkgUOHGFI1NG5Ctijh4XV8GSsjVqF
Q4bveMRD0T3MItdNLx85Ev3DoCVQYxYpGRm84cummiLhrMgxvId/uoxcFbdm4NzRxl3L3VMOBHhH
JeD/saQ/d3qevbbSf08KGrjChTuYmhT1ew+R448UkY4xFmyuMND9i/w88oOd3PKe5pOwZmOYc8ze
yN4UU/al07ZxLwM6iEfAdAL767YRVRJaqtYBAoL/wb4W+CjV+gJGk3+r3UzOOof8k1PrfqLpaSJL
E/U918jRZp/7/FdxKanEzlLe1pn5qqqTOMOOHki//ocCIbQabkSq7mnrK87vL459TcUh5AQZk23Q
v30IzgDXQp/qT6451XsPitqw18vU+HJDFVgMtmpUqUanSHUwAZDjc7llzNwiqLv6lsH7WHEYpngm
KSzqTXr7IKmU7TEgIV490hEmdjMhAUm7xduGasf0sMI2EJ8KIisrjXN6aELlPHzYXSNuOZlQCoq0
OgxIy+izJrpVNIBfJ0EtKfpiB3DG9DOEfxF10EK1dJz/gfg1eGL9nyH31BJYEUB6ffIWwHmrtnQv
wWwJCm74zJfZYdsREzB+Ky0+rm45dTFPQEUqSJGEo35fa5ed61EVLI/lufGzfkdco3+/cK7m+LJP
9aveMP+bVA8CEKd8n+tIGYteIM+F1MizR/6MPGnqZexy/JKigvgfNNpOqs1ixrA+7c12IytL8Qn6
sHe9HYfgSeDJByZ/dfZ5LnBpQFRAapsZCqVJ5ulMj+Q1lCAZXhlCWH5I0tPyXil288DcScotvvqk
WfaF8Rz6wBIfC23U/tik2MG55wY3pJvAI2mQLqvCBXntsUd3BPliaRl59SAKPAitcvIw8sBQ41La
PEa6JC9qXWSnK/N+aWGyOd+3Ze2XT+tvoBowoEd9+8E3K/ECshpNtT1rOYehHaP3Y1XUkNGdRNaP
I3Z13OI6+kWNgEEkj+foT/yrLmNL94ZdLG2wkV2G5956VKmQzQXToKhlO1Gx+0BPgE7JV7W9u9ep
2tZycU7LXbAgXKpnCPwq6OSsuvFHdNc0eYWJq5J5hvxe80C2MtUjtX4l8C/M1rgdouQP23+XfGEL
e+RphM83BEbzHrFFUyegXe87XK7pBF8St1ByvdyTi/NTNNBgzaA1IUf0ro0CLfJn9oiLRdR9tpSt
ArBNr3c7P9vNuwQyUkFR1ZLzNyh/OK9PRXSNC4YIEmTmwAOrPM23UQ43Cf8fY/Iys1gLfOL0o98q
YrIBLuoBdAe9umbxwUUWSl15PsjyI5O3eD5L7ngT+9aQNfzPKzSRrPanti2o7Uyy/R2uswzwUV7T
vPh1etVcPhc8y/h0iWQCzLuSjzKEDPzmhspBZuR1r7zMcIRI3x/rXXx8U8QcqL9fXGVHoZnMorrr
pzx4yPwvAm2v74oyILhUTjBz5McSG2Ph/dqTHX+gH7aHiM/EvTeuDi5rCYGN53nZXLfGNWbauXn5
8otGj0x85hyaYlIBHSb/ujreyoAGzpdhMZbiRwkVFoWgr461T2IdHMdcpNxEmHppJGmGTji374KZ
nbIvriY9zUhaFvjpgSeKQmbm163qz3kFmscGpleM375nLHQnAx1VUBaHcIb0dWPb7jGXEl+fGaja
ewTbACGddNuP3S8bgD3e8fUY+EPxzfcxXwWMZ9Kmog2S46SvsFassjNNFnoLW07oFoWk8i1Ghpm3
tJYUyDYm7D3X0CySTcKiGYdGOK309sini4B1zppq9ehCu4LPQ9ltwQ9IjX4SnDOKFLC5m/nG8Xjy
T5oaza18hrqxVNZ/TA4rUmJFVp0TKP15goJQWgwzlexOm20YAC+6e9ia/rAWz23Vq2rDclVoY4X1
xVlApUZhYt+xvG/NDGi/yOtJtYKZ/S/sT+N6NUSFO+U35PrixMUyyWJxtcWYaah9/w6FDcwjV6UF
H1jXbfvoMGSqNNRISV3/b4Xzp8A2Ohn/25l+TtL8jaJdqC8VmHoeejGriYV0YpiJ2KGvJ8a1yOim
BTM8GWxCQUzY7CFwpylRoPK0eDvbpf5WWarTEhkwzF9pnn1FJYGINfLIdzqOeE1Ry727YA5ug9pH
rztl4TkE60Qw4W7hKTYyi2J00JoJHMpMf06LLQgQNC8nd3jjvQ4Ijvm1PTXfqY+ijmk/83SSsO2F
UzUz7AC3Eo3FV8zHH3A7GfS+9c5g9gg4dD6fumzZjw5E+mWWwoMlB0rAOFtYTDPcCaEPJzD8Bfc0
SX+TpJ+coira3YjNvHP586B0IY2mrDKyTOE+zE6UZz4lD4/O6dg5nCzIJgpxG2/M3nX8hzjCPMKu
vNKmj66mSuuC0gmUWIPef4AT8xbcBpBre4gp5YzZ+y7kLEyWau7XwJlrrApUjujQdNwE1K0lYKg/
S2YUokJcHnt6iM2heW+5fH+g8C2hHarmDEsPWa08OBAk9AIuwBbeV9m1t6Sl2TQN/oM07Fw535FV
X9b8iKJh/G+REg1c45RpNiRWeZW+mdAY9a0LN2Oxn369vQgEm7sAQa3CMkwgIRWIbMGRDqKhvAg4
oys1uZuc7llHB/EAcKx3OEq77vF23Jy+Y63Ifnh1hZfdKvrqFC5SUAgT3+htNJtkTSgbYGjcu0YF
fUU/uFdtu2VM1snQgcf3ZGcdw/dtgK0t3b2lOkM+21l0kuB7AKfTNVtCqOMZ9TN7DUY4mEWT1rGl
3sg8GxmIT4W6PCghbqVdt2Y/SnbdJqPTdx0WkrEcCb8Fv/v86czxEb8ZylHlzggDPLXprhAMevMt
HcaVCs6B3maT/wYWw+a3JNZu6/VVc3nu2e73jBCndRYjW6xF3bTzq7NulRDYgK9uWqyHy8mMhaak
LqKZZIEwUz9aYcUwjiNeVfZTUT/4cTvrGYHZIHDoTxkw8sS7voXkmp5Q0GQI4593cs/BBSCyQ1jK
FM1EUQhJqSvwL55NYgfoaguhyBCEj8knydHQm6MPBcS+L9sce8mI/cGWiqQOeurIluzQHWZNt941
8ibNwPHg1oVQVORJLwfIZ22lsrgm1gAgiGfWgYbJCH08liSVAFQjHDDjokuOR0ZKI6HM1IyWi/9r
Ba4U0vlEpM3V8QDlsZgoAbatMcKZSANEzGgl8S8ZL5RfT6RPqpMynFezvyNMHYT1hOfSt4xDHNMp
/Xv7KI2McO0Fw07pnzeKXWtu531eyCf7pctBs16ppR6lWjvkJuBZMc8goVibLDfWhAl48d7IdF4A
Zjdvt+mrgXQEIyFKuD/UaTOEyeVf52Bjf9D5njJw1wo188kYRs+6WLvrVNDqk0Bo1zvb3/byVrZ+
2o2wS+gyAKnuyazEE+cM3eLCRxHLOsdIlRzrpvnXxcNQ9cnwwOR9n66q1l6++KvmiaKqJyNwhVcw
t3fElLOuJrdmQF0GBx7QCyjwpOCjQVx9KuhoR3lPHEY/bJT7OvkugiLW1Rghwj6MNEe3EQV+WL7c
FN55biPbghggpKOSjOP/IcV8+HKClkigRtBTwkALf+JZU8yO0teGngTXU2IeoXi/Hhh4qiCRWFN9
XgWp9tvMcRdL8wwAptA4OgFsCScOIIYNkxBHZMCLpmgb+gV8dMjqu5W7RV7hbkTZRLMjvfnLgxyl
1ldwULbG1BiwFS2kMTReY/3ExbEdvoUTKVeOp6heXzMi+WO5097dgXEaT8gnx7tT4TFEj5U1fz70
2BOK54WIuayybNc/4DJmpj20lc1TRp9w9/zeeJkruaZnXFJacTSey9QGL+QSJYTI0qW058VdgU4l
oi9EVrzjswM7Xw+0depoCncKGYefRyV/qItDqqVbKO44C7zUywE8RVXJ8aCkMKu+JlijaKEShPSE
ET5Jx+HZsSQbSxmngO6hKVnxgoklvjTqz+ml6pXWbGX1DqA8TeK9JrVUHqNytuYGcySjSVFapEi+
h+OVry1t46wy2mJPGyMz+MbibzU8Jp3gUoD1Oyx+jofvCL0EYyc7B+14WM3ZxB9AoUag0b+ZNvas
oJD9qJIUMNwUytztvwhAf3NjkHP8/g9Hz2soH2ao9pTeWq0eZLUSut0OoPnxWPewmKmsk75TrqKa
+f3CTCr2ig97PWFAA3WZ1QpVoAD4KYMCdO1nZGbqAgORdE1Lla6OmwXPhSCU/XXNPLs8LpHh4P7D
blcvlY4M3Ph4yayR2BcTA21Ngea8tELjSCcMl8/+YDiaNvduOF9n1OorLAxi0TaURxcbDK+iHLa5
pkih82rZniBuAL20JRgfUBzZPJ/LbkTfO7Pgha9CWlVIpiZYgYf8f81VEuClAhF2ysFKAR6wfXhf
Qgr+ZIhZhPtCDpwAiLkHX+qT9cViruZB4edJ+urGYJBlrkVMyz0FM5APF510/2TLGse0raTqx4UM
K0XzYCDieIgj1fzpN+Qz5mb7FqaHJIemUetFU0DbDqhx74o6R1q8vL/cR0wyJiixY/sKLXOAg9Bu
RTfTUvC+Fa8unqjj4EMVoyN5o/odCicnmo/GZxBct7An6vAidTr3EBYkiOp1kDBRn6KpeOSoIwqB
87Ff10BSBP3zg57pB1qAL4wZ/gBoj6au6RQFT/G7PvhsnYeH6niPnF5cLWsVgRTeZAiqTkZQbOLD
faiZegs05bj8cdxoXpjk2nf6Xruehrvfk25zm7U7aN7chO/QWVkChTAPjFxMQ+rQ3YpNSG9ls4+8
FwnJECdhQdxx2AFQHorsgqdC/v+8t+lveNiAa8pZoo6AFlZztqcYGNOeJwdfklM/+v6roju/7P4y
UCIAfECpt/tKXutUpgTyV35JhKzK76yY3sH+wy6+KxnetZWyByb+2jfaHuyYBB/UWgjBUk0nh8C8
4pT1D57i8VSylynl2Fd65V1tgKxoeyK31mPd8Decs981ib+vkzhHb4f7XtYlEL9RQPrKihi/pSEE
Gs8mSH6FASE/pXdnPWK6IyTrjA+Zv8bzERryvW5dcEzcbLRvv94zFkb2Xh9vGjEBhMCsHL8LPhY3
QYP3GKaOAB0ZCodTFr3WvqoUY+i3Rt8BiNPcElKqkKmELRdmZrSIhKczDXz3Aqh4X94ZR3W/sA2D
9gAu3KLlEuxrJLO5OLYFZKq50E9e3VxCjKaRVOhcCapNCkgpzGoiVpGLtQF95k+aA4MQ28qQRE8M
Tj0fEI62Oe+aVcgPKE33dLLn4bEQeIdrqjfbp+IJUalIjdYNe969SQ8VH6+whBBzNbT540bYqj6+
Dv0kDC3A7o/680+n6OIKE1RLJ+/+RPCN59pQkElDzB+ZyGDRkIZOUoYK2rsJbNEsPSEVXEez1icF
Fs6pdQWAlGnNyfUyNbdPA0XKNHnFFdc5IWHkqpYAu6VKs3FRKHlXDfOkNnJPCdgmo3JzGklEnl0s
ZX1s5e9LSDiVAZDJG0rXz3RUCCMQ/vkHGtuznPu987MZv9F4F21u2eZnAwT1Ump3miZvjHwJIfYs
2z5kXz6BtjR3PeBo7sg4An9xr0FBqtC+alEyAnXKBQ9OOOrt+9TmGGrKOdnOXprYVuEh+f6w92jm
5I51XRfabgPzgPAq+tXPU3qCpWkmMKICuhP5t1f25ywMIznTLaiMlPCyF2BprcIttkKPuMp8P9Ww
XpLxGwh6MBHuj8ByHB9qhmX5McEegR8MdMQRouvzbav9fRLtE9TWLP/YyWVdaINBo2c1nR5eNy/w
TDC+bFuqMasp9G7sg7M2+l6n7XTyId43w63LegUlQmfG5Gm+H0NQPWg2HvbZ0Pup+JrNceHJWJ7P
MFRWmZ0gm4fA87jg4KQYvtWHVkFQTp0hgDMg+E1RF0b2+TOx1Hl9fVPjWEDTid8vxP6ZrXgnpwE+
yLN+rY2q7HydDZ4LAon46cfrMXR1xZCDR6BVlDrqqQf3Ty832q8JLIqJTLMc3VpG2FoC5lrAur3F
DFCe1b0RokO0w/z29ncPOLRSfZ6Unnh/LkUM9Cyx5cF6ZjWKacWq5xuT8bpKFzmdDiMbrcHaYSqz
HIf2OHTr8B1BfG/Ad/xunkOs6K1qCnPIFCdm6C5nGv2qKWMjd0R8RFzC9WWIZkwBK7MGIhWKP6Np
+pgX8OzLR2IkCHRKcAJnxRqsIVr2eSpHYfawSQuDCe3ru5tHO+/Q+Y86xArqmnWzGQmtDzHRprGX
MQSC1Xrujf/Lyx7ObovYN2EOnlQRfH4lAkz4GfjwYb2DQSdHHaedAPxjApJ4W1PHVKnkI/ipz+2k
YjjJf56VMgggkRCj1nTboVgQexojE167u6uhkwZK6hkM5ns3t78KXXMTQeP89NqS15pb/Vln87un
yuW3Hhl2u6eoSJloWa3ocb7MvtwzAocNFTJtqeqQ16g/LE/jKeI92s/W1sp8E8naVeJV/AiJwTjD
kle5T6CTw1WbpIA0mc3sItRrImoUoCK/vcQTHTGDN9MYBDq54ANkCP4mHqDVBMqOTU7WksfpgXoA
HQxM5sn68V+8g8wnfGUicb4it8sJnnx43ywaSSoBviapD3fnCPsn2mHDqAuoUZZ+Mp78lXd2hf25
zjSKeGuTA0yhFFYd7N9R8L3JPCSthAY6fzVSKdizX0MQICI9ZihwK9/SMxQy/aq2zXPpV9EtMjfu
vhbq6Q9Qdt6DgVIJzZfsSFDAR+kvWtrfeXjAvV1izbXFtQsKLh1KgZA57cKFmaukflyn+0PDsZBd
YF8CJKsIEeOWA+PydwJ2wJWV78jvN37QasmQ2Rtw9VPfXbhhN7zi/ppwpkl5YuIa56c0+xIs9Mxn
sxL5JAmwFhob/P+kthHC12YwXz8O0zeQ5uYsYfNFnWk/YLSNcAYzoeJFS0FPSRxtY7I+izan0PRo
6XTbuYeeM7DaD712qYzX5Z4K8f+f3rLZw6d/JGzh6g+dE8E4ET/y652MMHXwCLmGCDbezsXXLSp5
bGFCVPZcMNgQvi55O+zkB/bT6b14jW5JniOA33/KLlg111Bji6zAA8Y76NMQn89AK52OZLWbeFdX
HV38Cw3tuVSfvAPCcZa7sSYmSc3Nb/8BjGlhIFUlzMmsUNNmuPPvYKGXTWKUYAU+cL0GaVNNM0H2
hmvDnuE7Z4/aIlPn8xt1ubjDbmn5esiuKxiw+MYgUcoKW5fYfFc3twY8kZnMjANvyQUbbO+jJ3qI
NiPs++ImUtkK5zW+rE/HBazmOPu1yjCzurOotFaVg/Cg4blrnk9RF4OWxDkuYrshOQe87SKg1eW1
/9V34Ulut6CX/nvHjTd66kV2jnHtT0dkIM9h/QspQo9a4cb98exSp9lD/ztLuo+ZlVS2Ir/n3VUR
NaIg8alznj0HA7fiQ8S6OxsMxV2Hf2cptpz0H1QanVGug7qcXcqfJWi1B/tk5JidmbjORdGwlulh
f0K2nEyxEyRC3tP1jGNvX23I5Dawik6hd2rciQ131bNCvXl5gD0mtAL5pceHJ7Wfy2LlWoRlTXkX
rFPMVvlJkjvFr/L6PvPSPkRaRHxIl+EmlsHlhLqPpMDEJUU5eToDOqb7P8XV0cQXNxa82rW2pHRo
UvJytLAVc2skWFm/73AO4WNAy1lpZgX39FqzPcdDLRceyIvJWEqm2JgDjCdXd0iIpr0OtEkbH2ss
sDEa+u/VLfccnOvrr2XM7oV5qliyJzknsS12yFV0ylC1qZh0RB8FoM28y6NOQEVr0k/4ds1tNTIn
X1Qc4i/5x8NA6dMAOmtzA4m7E/40ZpfZeIxz2pvnOYX3R2uFr2f+8N9DFn3Zw65hi92ESsFLA+vS
bbrmZ7lvw/pt5hWM+xIj/PQBiMB2+/67iS/mj1LEOVpggv/fPuanoIrk+EO61kQzMLMYap/Fz+MT
o/CWxj35PR8Ik8VdPdX465i681PY2Ti3z4x0lexUYzyk6p6Iy8GHSlv0gZjo4wcqEBm9u/LEEOlb
m6iWUfVdvERaffs6L25MChnBF6dFmvte/2pMU9Y04qwMbWB6vCaHPE/CVNVz9Wy3tqLVJjCBa75j
boQg9dbFaDs9Qa7y9CnmWomQb2AKqNKgr4cUwjit+aRjzyxCyFClEHTU9uni4O8A1LqNrJS6Nqbz
Ew6FD8xIai9ncsgBELIUomQ5whoEsKHZxTNS7qge/I5wMjzN7P8BUbVUSMpln1xE4FfwsGirwIVX
K8ilH//hVaKIOSGrLEhllUgVicqlVL434n1Pv/8V96dSTLxw+4rEPzyIXeSoDfSGVcECiErpXaDy
4DN1orxRzNLx0KR4cvqOrFTjTzlNWnXdaVptbwGETIcjHCpQwC/AXdteirGmy8CLbqT1TV+cG3+E
RABVvDdhQdGix7iFltRMhn1wtEQjC5Tj4rhnquhb0Zne1Hk8SzK/0zU0UMELafXs4UP0/5tGod4g
eufL5bsUSG14z0cdwUKGkmFHJH/a9qY0ACcAK4xhHARmeuZ0oC6I3+OGBAUd7AlOWIloyUgXXZFp
DTyBS1q1ptgUPQPZZrtT8WAFpasH5DV/+9R8g7XlxCpRbUCW5OnnyzMtKLz/1PqYKwhEHpZJ7k8p
MTadgRo9L0kmZgmjebYNTirEdi/nO7N0ZevKyRkLUJxKPHHBku/UaWrVXchVpalXd7MXW16GFLVY
8e6BHEoLBCJBW+Xtcfpy5iJMbvgaJM8HLQyARGvKvtRJnOQLnAIC2xiL33HS4NDIY4S7a8sSXq/r
pKajppKa/C0IKDCcHq9GWgju0UXTJN/om9pWfblBKeKf6JwQKpYkEO0epjz0r3HRXmOMhCi98h+Z
AGLpqUSbNjxTQ7uNA8CW/U7coSosjLpWBsW7+q3YZXQa0nSO+mRryAricqLOnZLzVmBFjPADvDpk
+h29vvWZ1NBegfP930cF0ha+v6hxYFJSMkUb9f26gUS5QXadnKmU+am+aAJKeOMy2nIRaknOznQZ
jk3+4ycFEXyuC7mj7DAi6UsBxOrdO+LsqyaGRzsZ9iKSZUSf1LqAn+aiFKkgUySo2nsaZkutnXZJ
esOeqESi/hwnuFQCezEngDLs9+P5hCHvHkxnjD8FDayCVOwOTqwcQUGK5TnDWIE+Ibwj/+AhzL/v
x2zHwmiZ9MOT0hUHsimkufC0LBUX1p7ybeoD9fohlGnXsKrSH/mgU9NUo1oc3XYBMQtv3eESSPD5
8Kashd9AP1+fAxOa52qosQVvo4g2qdG/VmTI30iRBCeQdvk1ybEUWfif6gBaBnAUbFLrixjpXrPJ
WG7AXmX3LV1fxNj/sITgW1MSJodQLJTKv1qWBSjn+NMzCokBglDdC7lKJTgkfx94vYaaOKo9hBbQ
JzEah3VNUo3dc9hR0Nxo9b0XrBuYsts9mENQ2oBP8737CX021AYQGTA547UBfphx/H6yREDAm8S2
fjFSpjfg62+zR+g9LgPLJAIBEkUbXmx31vDs4c4AFwGlqwndj/K+ZOz3QaRBOgiPAPB5KMrokRvR
UU0k5rP4tKTNpdAm+472Yb/3sw9JJbfB6AMDAVy/O3NXe4YYkQZtjJLeu/W/DZj2YtiJt5aREBHX
k/Hq2fLMqW7EW2RCAFTrP8BTtwQe6jd+Kof8M6AHA5zSsq5+u3tR5oSNvRrNmeJnP6E1PBIcMLuD
1SHIbf+z9YAGfzTSBIhpqPXaElwQq6vBOCEH2BxpEtbFAM4bpChsNXQvNIDZuZOKKVn6d8+kaJ0Q
PqACjUHfykgkcBSwok8TQOB/+aC/geXyPD0gGy6A3ZmuavImhKf+e7u4veCcXG5hy+MrwIbu32Bd
Ju8puSeLyFSO9UdNUfSQgYhzSsJrQ0EBRpdfhTikL4XDf2emAGdQVtLETF/IZezHci24XjR0l4Wj
oTa0I/uIy31QQpeb3kiuNRx5Ibdrs11w1yw/qHqlYeH1x8n4md0Ab6j/5FXgUwM9f43N4wDASZh9
v2gJsU1+QT67M/OlljvPwTTbmv4T7RKm3W07DGatG/pnqSlLiQfV19xxiluwxIfCIRC3Hic2Kjgm
8wgvpFl8mo3SIna4GQgeGQqjQwU1xHv0GycAo5r4+x88J+A1uu/lqaD61+oLkl9tfNC6/YhKExf3
oPd+3vxu4f8QWa+UsL/HUc6wtWzEtSsUED1NuAt1ttFhvOFWGMgva+ktjsO75r5tr1YElX+R66Oy
vmjxHdM+PS2itS/oZZzm/mwnVOKxK5dvXwGMWzfS3h5USWarl35cxg4X+sAzWBHo8P5A1IE/clvJ
e5aSvayPK2ftxghR3Yn32Ut7HPzEDaCA+xxs040wyPkurgGo6+XSlnb5U8zQRHu9g0BM/9QliaAT
TVRvN1jNlxwzMDkN2o/2FS4c9dmNtuwfpqwrjm/tTFWTNVBr4wpL0SVBB4efs9F9SpYvRC4JCxa4
FLx5hJJGu/Mu9bE6kEAEcyuMtSQHKyFTFav3GkmtxTJFoHkaBk3GyYbT4/63gq9CX6uyDlhGINKq
MViUcN3pSelw8wPQBFtEFlrEkdM/EtGQg3xZSCc/WiwiYIC+4OUe870jPEmH1gM3e8sNUbxdNh6+
dKp4SfVKV9MrwBxU5sIcwy8/WXqJ81sTAk/31fnc+KPiOIp/KhuCRV1lEklx9FJ9kY1YZccMTD6r
P6gANcqqT6u0dAegznd9lfHF27aNfdMYCHMkhU5AqN7CDXYz3jrZOtAXEghqH6RU0UECm71Zk8B8
r3Fz9ZKTEPn1X1EBGRrv8LT3OGmmfZDxVeKyJKfG1J+dHwa/Vx8vXcP2l6ke7huuclhgGH9gg/Si
3zcOtfCSa/rjLo8QUePPkBDkx3IGjZZb7UDD5g0i9R7jQqksB/LFh+lvC/cjMdcV917ojGhWaQdd
bbsWN5LeaD6P/O84d198bpoIxKjFudaVhO8YuWKu+c8kM+YNBmOCBWV7mBjnBuPUKq2spyol9/wo
XcdnKXSzee1QESQBtYQeub9QGd+7uOtXzkdpcCH2G2crApb5QOby2KK54hQITwIuIZ3Ss+CeUm/D
wZwyf3Xe3XLeuWbScqAmfABR93tEJRtAmIUFJdO2WhKEOTO+vl86aBul834tf81Bf/R44b0YMIKY
R1p0jDzvUxyuOfroio/wfZwtTkEccEPVR4s//YdHEfGJfQQ3zs0XL1o//jPiEPpbuXUtJdqucALT
XtK/f8UMNdftusRbJn+goFMZ1YW6UlhnbbN9lbJ5CxKeafwKzEUTihYwGYIQBNev0f0M+Z1/XLng
1DWftQngECVSk7pmbH+/b1KFyOMEbm9My8RgeZPs1gxZZ9Pg3dOKcbTaTVplU8xkfVPdFP5cxN/t
ZtIp7VZ0PiquoyNhkTS1tOJVT8l3WnbWAFuMeJKrC1Xhbue3fiPQwFwVBDp5DaczRnILZnsD/rCQ
v1I2imjvxhC1yDe04Ucq6FP/QtsoFoqxIcXs5mKXy8Z5dz8KaOvpWLmhcbSTm7JwysxYIWaxxKl0
hpmSYb18iX0sCW0+Cf3ochHmfkA1VXlbCjEKjh3hRFO47//rWNgGC9XPJ2sYBaapMABVm0lfvt47
HEIiB234yyphDwAiY+vA/58gmVFuX/GTHVpG6zC3QoThaO6ZNMNJwf3mAp/4GOUnPgfabUZPWkQv
iH8+3M4zk+yznhwDXPlE+7XtsVZtn1mgIwXWKU9TnsuWYQXdyS8mHGJE8wK2Bi82So3z/9c+qaCo
+JfbdfUeesqPR12iclSw3lWS9mWewVdgh3WxhMFUYNTnfjaHRQkA4T4Ll1+EJevksYaHlFQRL+Vj
+lFeSYIJmflx1auKZI2Pi/Zf0WvUpBONTWtPvC0vQ3LRhGSxVdMxCIAZFnlWj1ybW5HESX4ckJCL
xXmyp/9MX1ZuN4uDs+YLotkZqZZJOEtUOCbwqOjPLRzBzxG7V/IrlPyOCww1OeOyEzU1d2L5IKLb
tOI3+/uem2JAXjFxkSsN5hg65WvvU3VEIHsfBbwId5nkf5oIABFVrcgNmmewwP+J5HTphbRln3GQ
v2gdQ/sPXQgA4K/vj8qmbyvPNohh4iGyZE3nz4aOWm2pRNV1iPfAA+qBe71oWaAYUkTEGkhI+Qpo
rBGU+VI5kNHFXoGkgxZ2OWSwrEDv/OMMJkKdo4oBFQfWepH9V4spl0X7pTPyloI1mvJwMct/4Ua4
smQdSf6yx1BS8xwbBXQNDBQL61n/KmRGmQ3sxPTO8YxN3Mq19X5eM39u2ivlt3SAZX3pK5ZN636W
hGavj81wRFpOfKN6HxaPApjj76zzz3bBMCEtpK9ML611kyRn6+c7b+cpmVLwagzZ1zK2vtaU5rIw
0RPzfTRvHELXZr77sbWWtK4EPYr4V5Rw9SyuSi4JKYal4Q/Q1xwdbI6n+3mO8fZfPV8ADt1yZO3x
US/FiLXQbFOADPgnWu2h8M3mWXoytj2L7fcy7vERI4u/snVnMnzXwL4Ufrd8vIl1dHsYI7TEnujF
FGgxuwMVQSOV/OXUbUhAHvnjw3KKaqKlilHIlGBdF+b/pddF1LxgX0Ue9tkE6C3Fot8NXCa9F/iQ
/obqweZYVhTN86eNySxS61cNnd9Enccibfjm6LLwdiuGSeZPWmlazWnFXPVCsfwVY5JED+5gf02v
2BkQKI4zhJlqvzru322iXnFDdj3bq/GUtyNAIi5jWCmsqCaKI79L4HImq74QzzrSFQYlqVykqlNh
5zuetNmfykKn8aFwE0kdmfFBMRX3AgqSC3klgb9GHO812+RAtaLUeOdWXZXaxfq1vNqd7x2DP+EO
2wrJEC6UEhcl9Rgq0W+W4NpV5xa1nazpOolFqc4fI8Me39dtmgeOPTFwqHUu1FLcnGLdWCaIoYrq
mnV7MmAgVTip7626cJJpI2nbfqhchb4+YXpkhQHAtnI6WpKAmycOZb27JegXckBvsuWZh4gQVJxc
4AdHOF82S19lvV/1/zX+sOguAhRcNuB/H6aFlHmivNJfHhIAwXym3n9HfflP/rZ2t9+8qhknELPV
pAbl+wV4PYLPEMfh3ETW5ZsQZpJvHY+8mLh4+WSp1karWYcdZJoKF//WtMZPUyxJHXzbpHq503vQ
LLkE32HnyhNEmyq4ZrIC3UgjFXpkqOh0kwxi+T4K7jkSr13b4pjpuUfjGAA7rj0TrF8PAMd6LmJY
r2yRaRJze1gKJcYqQwjxZh2ORJh0t1YqTm0JfSN9S5SWSjCjeGrRdmud0DEpa+NEMGB7fplzUfTE
HQrCjLDApP7u4XzAXKKP5o6ctEu3muGykW26Y5VP5mqjSMNMN7t47z7NM76pSxXaLh2s/GYRVxBA
osRYZMxMaDYNHsg+7QHF/DLFx304J4Vym5faXzxbatuyPkAJ4BnntaT1w2RjMFsrFJ5OQf/1cwQa
L8bmu4o5Efmx9NM+2o2T943rp6HKugwfhdjlQ9UKTeZD/McGW4Ac4s1+nvumFAw7IY2aQ9F2Ej+7
oYD/X44anPvA9it1AlnUDdNrQyKrbK8tdxbQz6NjlRIw9GC+DXOHfSw0ynk3rd5fU2cON3CwaYs+
jho2zcBa8jEg7EEvoC+cn2IzXKxcfdhAp99Tl02w/QskFn46OpQ1THuNTxBtY+B07nKd67lMZYML
VX0ubNLMU6QMMRuYcXGs7fJVSOVxBmGb5dIFJMzvWP3gqqiiCPDPSfiV/o7wpcONtF8j41o3QcC8
GYMbCqxUxB71x1dCneMEJoxhqD9d3KXjjObF0O7BeBPXqSY884/OHqgRt33QnWgNRQfn7fFA/d8B
9we2PqjPaRg2XdrTanWwqQlFF0Jy8GZr9Vl/SVQxX9Wn1ikHf14GE5HsS29M8oyfTVa0F2lt3gg5
ohVSqjXF0/Ches3qCIjboDIT7JoPTqt6/R/144wBtupbx3VQdljBqGjwLDKgUg9QgAvIh0GLpjQb
18M0fkB7Z7Pte1MmzTSba6leKTXaIKXjmbINwx13t6qkhegLVKJhhGsolP3ZWm1L3nDnBPmRhsaP
khJ1xrYiI2tMG/wiutdSGqdX9Er87aADQp61iUhskbX3S7iQmFS/oz/viwSx6J88cZUawX3QMSfo
FH4xzX7+HnesE93naOjdoBppmaWHI78MEC7nnmgl7A4hOvW/o6WirsfmNIPb1YlplbI0MfX5vn8t
xIURwCYl4YjtfF9eV3yuXMpbMRrmzbFUyzJRBQCdekJiCe0Q2MlM1yoy0oEPUoPz3CU+94dHyGZ2
xYUAhkIUs9rjg+cnEBlNilVU3/c/iOIor9f7sdKDLvuHAxCs47N0IFjmUudveRVEoDd8eGlKTTRJ
nSb+k+aNRt419sp5BX2Xv3x7JOEQl2V/xBDqffpig6Uto3wUG7QwpY+qI01Jq3g/1TOokHvZkCO8
jfA2Bz+eOaB5tz8FHlp4srFzrBkETPs36PapRDASYoHK9BBi5bf8LQbFUfR4yMpTPM4fXeW+Tiyy
Eo5stk4DXC39XnTPJ+dgkmXjJ+U+LEexIN3OuzBjGMZRpJg8wT5Y+q57I9VeAeevTKdGSBvSoSq8
H+4r1urXKxwukxDRPwCFaGAE43je67A/299RJQQrPj8wrfG36pf+D1XUmQs5LQQcBn4YAmoiXFRb
fzMG3fIL9Pq/ZPWxneG+KaXs4rULI2lJOleqvSvIZYEL/hZL/+OD1OS9gc1Lv8iGoRU7ILztBkii
a1VHXe4DGwA2FDh1AVeUfi4o51Z8cgckm5lHdgtupG7qio5DDHJC+fMx14VKv85vPm2J5ZhINK6+
SayOE3ux2/pSEvhw4EEc062oDHjyldI9dgT2IDQn4UVS2jKBSC7b0PEGVLNnpEqjcjiEGcBLDAm/
7azcOnHV9XW5XJht/+CVbLjk/1XUiW3A/rdWoE1mrgnBYDuYcgwyNEGZC/DXzcnk836trnS3pSei
DhDgu3tIyjjI7F5UrQh3dP/E+6K+WLVktDU8nX3rPUekzQzcjQ4ZcEsz38tKYqIaiWE9ZiOVoWWQ
T8fuYWdahSKrTWMxF6W3OeiSr9g7hjrzpdSwM0L2MCWbj527kKHnf+BG+QjDm7Wbr0MIKHeLuPdF
IP+AW/2Ny87cINegSJ6FWoXQssky5T8Nj/4qKge2ZNyJHMuOWo6kDUzPUS/tYzvw13f+k/2S48fv
HtQWYpSiUJzFcsd5yVbTfuD2BI4NdwmrIbiLAnIK2bUh9erFaevkgcqSM5KZQIMRKiSdOc+tIfxY
vXjXZXip9v0u7aFBMsZeSf3mr3Yq630XkGvGBoBHVtIHAl91XAb92TRQRvKsnxHJY+1tLfi+reTS
CZuOhB6fYz6Id10gKynrws3FohynE6hskIj3qw9SrJ9vM0amNwDYzZgxNFxDLhMqfuuWnOXPqjb5
bn1nKQRdUaw2cEfhqIH0giJ7R+E/FXRvmPVe4nheib/GCJpz0zdcmcUYKng6ybCUcnjbyeD4Utmz
+cVHCBf1nOnzGP/9pDy+cPAffQvSsNmhlvXZrOSeBApqhlo0UNmUhxR4zUU1ulwV3Z89NLWereiz
K8RHnyPeE9zZFi+c/EYDgMhv5xfuANiU6h4YFJBjioQUTIPfnyuEtCyqbWhVh8HObWOB4nqmEJI1
FIchS36rIjomV+zb1INlESQVR0hnksPDvu1gAC2tiYC68JkPXpIOP1zUaWVUODvSpsSsF9w5vBTe
DOstqsJd9n8HkOS3blGIN0aw84Y1Pr95tUws5QqECgn764suXeM5de/yMgS+4vp5r7LM7Wp2xwWY
EuQw+35eYi3g8MPd9DDog1qXX9NMDi+rdRSKOsDJcWazKvnaYi/J1LBlDFZHp4yHgf8Pt/R8Nh/c
cSjCgRbDnqXqtTPzTy0v81UCZrlEQ+c3fuFLCJedxuNERLEaJvQq3sWwe05090R3qwFjz8GpyFDy
OHMaeM+0gbc72l1SnYzATSaly+FOHXOD3Ooz0EcvokURQ3Dy6P6u/bw2IdqA7ssMtEm32Rg82xgA
ymDej+G3JuVfvHeKYiTO3/fLfoRzydYeTTjxxFO6tuFUFc341ws1tVy8GqiDoZg2o9YWWRYVi2/0
DTNIPDY3W2ZPW8ChDgPv9g8FFzmkbDE9LxvXlvI+bIkn+ieK2C1oE0itjOh+xcfY07skMeC7KVds
IzEgo3nYq6yTP4Qlhouf7wbuGM7jrIdrnVEfBjfvJGkXscZG/rRlY+xJIJMhIELwuw1F4j9evtHJ
hIIKfBnf0jYhi0gVvBWGhw9yKVH3lL73mKsgFsT/4OyBpaop5sMyy5n4hsf7nsw6B+r80JeHo6SP
Q8MpeZOuNigyFzWRZvKk5+omrMIdqqDlaVeV6UgSb8APKyFDX7OfvNqi6uT9fPeMM15LDsB5z3c+
IM/BtdybNFMERahAUq7XbgwpHzM6DfCK45jsd/SO/kwHItkh4V0rHlTr0HACt/Hm2dNW/H10fPeo
eNUjLpe2WBVaZtg0Pd2T+sviZgI/db+Id1FMrs+0WlIKOi/vC3DjvjEnm6AHfHTXCaf0NMyqw2rq
pqIzBAa+BDW1Q93WPGbxY9ZqUjfzW3WbAL/OAgOnCzyf0LxfOC4VE5w4zrNGsrJVZawc341x8umR
ZwNMuVf7Y4UG3wNkGQrz9MoEr4WOox9FwAhW5sP5Zy12VEuqIMgX4lrs3MxZuhsvr8X3XI0ZO/5Y
CNvDKQeTzfE55HAFeBiLUMJkJ/Q9cxNo/H7kyqDnsmjjM0IaXo7V/KbbrzekgF7KbNaufrnv769E
eUQxXewF5m/2/5WNIOqfnlD49yomXJz8v+CaHDeFobB/tzI6iwg8jkSklUIuHPgO/ypqgN7ox+0d
Niw7vayMRKSwcDzsXW78Qfl55FJJK3/fR+nzoXYaGj0f0+cIxqwOG6/D/D6Z1mKo6VKs0ibubtZ9
4TFHD86RszFvvhsQ/woKPrxOjqM1xxqFYEy0cNW6HCkV7RzSJmr27zzEv1DPmfuJK2t3IpgCJq5W
/2Yti+Yrlg75AKZC5n6RrHLz6DY5LKoTZQfWsWXrEFYuYCSsXuqtxQcSlucGbwrkMCFhKB9irXki
E/ASNA/FR8EiHlJN2I2ycKqLkU2Ntuoo/mu1gbw1d5wqR6o1h5HjYHveHNo06RKu7bYB9aK/dMPj
40Ixqgmj7upUM5tukEmbhlFBT32ckaGMhWLiI2fNmUTuKQqClftfHy01PpDHnuaJ8ky5aBTSbDkD
TGgehS3zXvrOP/dvgIBjPk5OO5hVjJQUVPzt6hzXwjnxSnUE3KN2cJ+7+fFVFJ37N57EXEtDku5u
yRaxSZawV5crRlmhUWbokS6GIwxLtNPT4aMjDBxz8TlL9/u4s09zNmedExflRYriiHsrI65wAdoE
828UlMt0ombnN4qGGQOXSur2uWOwARAx7P99pfFLvZWW3Xf2ttK8haw8HlB/CK/92a8p+NcNZso4
pupXbG+77YmUbM2emQVhF5MU7X0fbXkOfCtJKVIgyPfBUI1eUW4UMdpva9qookMc8axuxa/OQnaj
Abg0axFv8CiAIs/B94yylZ9GasEEmDDlF0EUqdHPdzfqaQkvHtSp8DEPe+BKprL4lRMOqrUy0mEA
nGI85bpIRrVJeiqqJ011TGg/27DuRKInMQOIo/Oanl2FbFsGBEP6DPcrzGc2W3GC8CHywMGVz0+d
SrY5tceNYNUPBm0gOIDl/ALdDpWNDb32KhiUtLhQEJzLYmGcgH8kAwHnttgRIuEl0t1rCAmmoaqT
oY8uEejCBKz7h8lb5au5Fp1jfklS7fmjsO1HZ2v37/PaGZR4dQtU8EmvBYyuZ/tCDfIssnkXHZvx
UtU4bof9hQBwWOu8uv/q7IK15WNnqfEgvIVMCjYta+10qrQGm5PeseXu/GO7TBmkO1L+sOBYxOUl
42wB+lQEIldgfW4UtDjC5aM8E82ImktDGlshjcrzwIE2j7D+5sFnj+RP9wJRrZAK273+mGbYxkPl
6oHvYckOeE6LgW+0WdiCo8kXZ1tTm4XeFnNvsyLuUQ5dsGM7gw2k06CfgqIPtwc2xl+4N8yyztKi
4NEjcw1TqefgkqFzsOinPd84u7mSj0cWdHrhGDoEe5PJz8asTT3aFSsxLjt8s/y8TpGXZrqBLRfp
hZy7AMG3gl6D8J3Utpxf38ItqIv5Q4eNsx/lah/sYLSBHBLjJ2UlH/IRm61BE1W9AGEGcxnnkfBB
Jz8PLGWHgtGewIbPkc7Y+MVK8BnLLKItFc/GVMXhXF978L52a3zlXq78V9wl9mwMqgPiqqRMMjY8
MZfuxd37VLlyTLvyb63NwJs2yAKapmNlxb2G2DLZFRKAgfjB2Ns8xO8In6NAwSdAcpKloB3gC2+p
577XCKTKOMy++1cBkCjTV68vGKofgp3Ks+Wx89YJvq/qXPMFtcopJxAeu5bNTFT33s/aItHIHcqX
yTq0R5HqEmryCfwSNx8mBGWDQSEgaHgWURs+QxBCnUscdRtleEiGvfA7YZ6br9lx625Ix9eYHoSE
9YJjixDVpoiFGDMwxm47o1JL6Aa9w+L+m8Zj47frBdp2+fBbSpbdZC8hxCz/P3RqfNCTqRQHdqDu
LCGtC1mYDZZ2K40GvnGXfmR8BfUML+MfPurv7uPNPDghx6NAIktuQ106R5zmzYHQwigsozTcNlqr
HTh8A5Amg0VFNnCwoLgQTfx2MXt5qhYY2nqb7ME9gKKOXMVWaFfy9Aue218hLome9agiehwphhyt
++Cb7Iz4nUHmRt8oJ3wr6rYik5dBhVy/QDVDEb3sv5oujZaMU6U3AVz8JFEXmMLdtrbRD0QxbFts
k4sQfy/dnQSIGl0hkQugXGzw3DTnHPu1WliPy1j3b1TcViJnuiSTgjVbqG8CoxI4T8ysPG0N3Q3P
+H1N2/1B+9j1ht3uhDY76FffkZr8YDI4oRV9LhsRPz16Gvu74ZuZeqMrQOPYQaxt5O4Jz1yuYHJC
Ly6teBJYzOIapYYBd+/BJWZJBbwIZyNMqHErT94C3pBjM3y5mTP5fBd/PfPTmYDNBuFNYxCsiBFn
H+0tozReMHvuH6ExyTVtifS3LCs3zZox7fpr1BcrfD5H+U4jIXYp8RQe0CNLVJzEqwjOJWZEoOY9
7eIRLWXSdVxL6o1zU8F6gftKpQiJceKzHykq8GRCcTAmmWFBJJHvS7utoMQ7FEBfk5QMB5t/YqEG
dYECKwpG62Qsl66UgyORzS+ptAvF4rwr8U5V3bb7htQJ3kUrwrlPWyJDujekH1y/X/IP/H5yf5d8
0JPlD4pFeQHhZ9p5ExMoa+ZK5wUlVg/+dQ6HrdfSNOtFradVHShBk+m5gF9146CH+z6k8/iByF7w
fkH+ZVxce7dVGSR1bqGm9yt/zp6sQrK7og4KfOWs6pFqHeq8lDpATAJp3MlAB1eFRiI8+Us7tw1m
PWxKETxIOt3jIlVrm5c1OT0lUsuFYqSyZpGraCcRB2NM1Dtk25UTGrQhMLnFdnSSVp8qMxrPjIRJ
BOIIY+kBMmW5VPa4fJ1trWox3OU36YJQ7rINj0jtyUvJwTa0ef7BaR3R2jxGCYxfRrP5oAwc1NGo
TlQ3AfzKbrc+OM2GsOlsT7zQ4nSW/SlhH27cBYm7v3FIC7JrBfN7Zv4kTlVaCPBF0Yn2FvI17opC
jJP7YyeDEo9VYHelQ+V6voWpgCO/5i5P5mUYyGGdGlHHPy9BZ4GIjudc0kM6Wuqd7cEYu/rPK6aT
GEEbblqIXk/Ad8Se+6Wj1B5UTJ4cU3LqB91DwGHwSI+WfmdEyGWMK9tHD5QzoUWNqMhdWbq5V9E8
LtKwLkA5GqmmUZkC1UPIq7TLsVzMa/YDqLZdQ4kN2fMifnvUWtzcMkM3zxP1LAqVRzD52H9s/g7M
UfOF0THEVemtNt+sa7Zf3yDP33qT+QzCZbt6A7u4GkuJxAluzTtHAAq1xxsrYxKVHJKzuAJsjOYZ
QKb2GVUzIjSgLJ7O6PTfEKh6tJgFAsNRfCwpu4Qfj7mQ+bzuF+bpCHPHvEKMbyoPWq8H3eAMPcpY
jBG32cz21tztag7mviFmJKZAEhFfI1zzYikw6gopZqouqgcUDUcB88BBr6mmKy6jazHl5hSh0wzY
BnOqxfWF4Fjh5NXSKBRMIxLxoeJnOSGMAoILAsDr4xi7urZXB4BNy4P0D+AIp5dAqX8drFWuOwNN
LjFFUexOrXcEuw78LcAVZCNGvkFFYVUd1y4YAdmb4P26QVyow9nqQKtJKuVbQQnD6l6C5ZoLkn0T
MBkAYNArbuOJamK/Q1Mihe0RKE/3a9xUb9f95dkrVfltnyC6CqmIKccHC07Haz9Yln52DL+ofYTv
Kc8CULRTlGStKKncZmuP+hQm/1/Vd5wSOVhQHLshoNeCkaE2XwYO9DNmp4aolNnm+aW+CeopkNSH
B1cTWQqLUfZ8CxHmtbxquy5keVdbNBc/mzoJ27bm0bhUG9PL1cMnHKhNBjeUTPcqIDEFMYu98HW3
DC1JqdrGzDezkiVQ5ctl+ZtVH20/l1pqvtN+MVHmV2TtCwSsjaz8E9Xja1nvIvVHfNh0J0p89MBq
01if2rxmyuXo+YzG68X+4uuLB9OnM5h+ZIqDE44jFeKdCGdsV/ctO9FBh4fvCGo5u5mD0YFqBEb9
eHQ6lL+Gv4YziaxRODN6TkRYlVVM6QsRBJdla82FIP2W9QVp/A9HHBZEt1B35OE7mOBjtN3jPXGX
GciUThr5ybsT4HG0gN7S9UuZsOhYm9A1MqSt0B+TZyKIQjUFPr1oALzBganqyLuS2xl63IO+7dp+
mW99mULuJtL6OvN4Lq715fH60nUGtQSIVqy17LLgwMG1MYRh01sHyKjS1lXobZNAexS45G8j25Iy
Zrl5wf9bej38v/MA1f6/FhngjmaF5GH7JZHGFAzxUFpJzQc6phOy6NBP9Bm3UFdimseJLHtrbgmg
XDj9jWcNyCoQ9OdYXkMDndFDi+DsvuFfOqERklQZ2q/UUImS5cekf+4MpGXnHb3AypPQt+rwm8VG
EPUUr51yoTyRVN3EfWfvbECXNrpe8sjVlY3Mrb9dPHbutoZzrCWKnEvDZKXe8FJa2wvmGyu9TXKQ
WqYaqt1ncjhWELkezGXzm5Z1xLdmPhsATeW8ulntgRWTPNT+ylnMvZcamWLY5SioFTLnDwHFR26s
mDE0vaTRl0l3FyBy9o6lzz0qmT28c3fQLXoDxzI2lqI9h+QYhgmGz1QkwHZ0th9lmtrXsuCJQWz1
gg0Ma8aiIsckaXemkE+A8LiHiji1GmPH+Nz0hEBgJB1hvcWAWCy27AGvnZBn0hFLFXHzzoOZohAo
GR1oHrF2lUkTbqDrJAFiJNpvJ9YJ67Y+4Ky8Et8ZU+cxlFsV333Ge6NWXQzQRXo7QSyFRs7BXHfy
M7M/rMFcsxvPJLfujVLUv1iX17CZOBP6k5xMrcmxNUcml6l6/yzbp0sUxRq+V0acPNm9qDjaVHn6
2djTxmlKB7TCIaYNromh+KKg9iLtvc/sL/IQbcHs38YnBx+rm5ge+H/90qirtQ6+7rrKbaMB3kRE
DQKLXF///Ko6G0uJzQ77Xr8AYFes6dM9KGyS0ojI9WUflqZgD87G9i8ddNYnA/T/C3eiei0fHolj
bcRRLkQi1kXTYvo2yftwwlTdVXTWFSt+bjg8qipdCrkdUz53jwTatM3hKodFULHr+wzdj1vnHVli
488SulIG2FF0RcU+wMprf+omZjklvdudHAV65LcRzN+msDGQrWGVXAgkWrt4Urs6RdM6AJJ8Cdw+
umAOD1TRCNwQDy9zQ6mYpkpgRCV4xEL7E5QkZMclx+PXGVqLWCW133Bbd2qsEmoeNHSSZHuEBy5G
b4Va2a4nZ119HWZINevr70Dko+g1rCQjuFzA2vZccUiAK3t5H7b/mNgnS4pedztVDLycyzDcoE4m
x85eKdJO687jGzWUQXWVQttZcgh3pnxvC3rEV34I7kCKGfRCiYiThRALcB27BJTrvBaYZBeVN+1u
YzoyjR7pBXzermlDnpgX/gc8nzdx7s4cBzu1cysZXqrtkDu/5jAjHVAj848HaCKvE7Pttm+z6lNc
MPj58NwB9eQxEovffQjIu5EaxZZklvXT8ItvikLUL4LTVaFfRe5fxqyLa41NV88Ry+/24id+VTxc
/tEJpSwtWxjAqtEGnLAFt47c59mIU0hM7AC1HobgkB/pL1pcR50qzJU4J/e1qiRyroexFJOBUnrn
SqjWsFBw6hLBH2lcdi79DO2Duw18ffmEsRzFAXrucg/Xegpy0xo8tZuPl22Oyrgbhd3t07z41E0L
QybVGHXs053Wlg9E08HveWYmjk6dy/suL9wakEipg45+gJpEAnnrmhF401DnF6d7km6Ux0GabQsj
0mEnPSYsrOJyGrlSZFqUGgGN/alipV40cOZWZZTDoOUQCRya8Bvse3Zm0JC6OBgqM5ueTOnqNeEQ
4ICsVZhneWuuYN5rKDVs7q0UsbHQ9CyNber94YQ5Zvpbsu1SP+ScjsOvnR8URP3g77z50Gt7J42x
EbrVbaKRoybXqW+Ryp6iBmWGwbdKEjvsyChyKKqfGRlgB+C/e/2X2ZyP7bWyxTUPaKnFhay2GHAY
5WFIAMFqI9xtVgMUJVkM6v7WB/lApVPnrlO0cs8CpHhLcN9Vcc8DuH/eMDQKdKTqkhMFOF38nHBD
bLImX83UjDldcuCAbNGye8NY9WiMoWf19fGA8oOQPPfW3UJ3BtPmTS9dchorljihVciaUIZZg34W
XCfdF4Aju/44Zz4kIivTb7L3qccDTmVX2ZdiqyGv48YQPeezBiYsqzdSGMeGI362Wo/2kSKyvAfG
qkZK2zct5tJSNlNk69QsIb3XbHN6F7GD4jH1+ktDRVASKMpZhe0hkVgAUve0qb3FxAOoOxmHdKCR
/aeb3sRWnzKoYmXrOMQ/MqzcF5uLmeWnL50bYEg1vKcaoFKlb06I9cwPIckeMG2IczZX6GhnRYyv
EJp5/OzqAGCgp7QikrZ31qdW980BLQhwdHl+WTfMJ7z7374sr2ph1nc+N+jrYrDtQZC60mF3AKUk
e1dGA63/sIcWtv3l6R7q9oPGepCHjXD2RsGnFZqHAPc0V86tg9c5AYvQmZHAmzmbB0eKsH0/26na
v/xm3+B2emERsinFmXHPqPIW4Qu0vpdV+Cm5cxA5xTtwGHJh2VvIKlqrIdzgIrzKqwgYvyao2DSV
pQcJ1mqoMMRT3ZZ2IScyEux47q1Zb+4vTC0ZuVXnlnfmAt0I6T86XJi5AK0BCzQp6F2G7tG89mPe
6vJQ/VT53yFMin8CXVzOUgpyznB6K8EqNX5FJmAAHsY4BSytEIKCRermk671mTkCLRWmVKIm4e0G
24waFBmq3IwbW5nTQnyT0B3l1/PMwwwnSf+zL5oPu6Zsx6ZBBkF+jm6jHMC5phQ3AUsVPdGi6EMr
P+5I4cX1G+5HAO7BIJSkDK3arFFX9E7zfo5Sbhsas7jIMQWaOk62UHctBic5znmNNW4YTUPVa0aW
OQEsfbbr+Fh4zAgzhdbcCv5re8Q87ILC02eGG0qc8SqXWS26EzGkTfcwj5FuwO/0RQzBKeeEjbhY
44/O4ikm1iF4QhOfBElKdR8LEwPwgXzh9KNIGXWuUrRptCurwen8+fKQz7aCs4Mm8ehs3kUp/w0E
InFLQ9c9b/NUzet5HUwGDuiviVYcOHVgOaN4INOfdm4AwQFJuzJ65ws0G1tYRj668UaNdGwUiQUL
Ig69p7hrthgsW2V0GAYTKP5x0980OYt0+3Sq0xyqIs/fzv2EUhc7LqvSM9vNMV98K41marfnVKI6
mgwLloRCJlQo8PampVT/KK6ARCUAgKxFL3XVQ2BFUEYWhNpOv59zqf7tc1vI6q5q1Dp8yX6BsrF2
HMi2yxFSJOuxkCnUhnKyQI2j/72n2LCtu2P5D+gL+Yc5he+O6lHJ2HIUhmYH/Jku/XBvb07lORSL
2+fF73a/54FKfeKft3Luajv5uNNmpQZz7hwMbxRH34s032XUwN2DChJf79lZdIBaX7k/IyOpXeI5
xRMYSf1JXW3Pkh3/SkhSQmbUCQJHEvk6bsyaeFH8AS2BLAwxskaLuc2gF+/Fgnv0U33hxyXYxthX
x3rvTbJ/WHLIu74qHLbe4m03rmlEb55xvwwihDB3EHYyB+J6nigMuj5cSQ3HshZOeH9Fwl31O9Ie
p9KD3PN2YAXpnsvuyVy6GTbZtv2p1o26RiH0IPaMKU4RzutZnGCJMWl4Nb+KZ2dssw2hpBOzvDTw
0LtzVo1kKXxRjVhCuHn+6ac+a29GkbUzSixOkq8vKeKYpTIn2JjbbtEgQ6SALaZM99t8VozTpWpy
JktBivOu7AZrhZq23PvCKmiIV7CSxbfUfYBlQkgQvRp9qy0+guzjFDMPuDqZhUmn2qgIz/1BtIal
H2OiOIkT0cn8tbJlBMFrFrT/8m4t/t2E9JTUBr2TwePc12D3BhJmUCXTqKnLLtRnPgJ6XgKnK1P9
lhSHm9IpRsZGFmmuxwXBWeg2z4rwBgqLZXOHKEFmtf/Zh890aJo8/sFzhAwCiT0xiyygjjUN7hPC
ziz49oP4WPwhxxMHJvj3BCjr0sdKqLcl/xgldvijK8KC38//1epug0eP28dZrrpdSm+2cSyH/BSX
fhBpFPyLft9ECCvqtyhEIag27Ehre7XqHSyFkPZXFzXGGJKSbC0rlN64vuHH+zvWipF4ueFgBEEy
F4Py6jGQ6mbkWfSxUauDrSX7XEbK1DYftsIziONrzHPNY69t1Hu9mn9Fzyla6+o2ThPwqI0x/Tte
81SX+kOz6jmaaK2vNNfdyos5Z+rmlq9ijh1Ht2el0OqH9URIkUnIIK2dXQBPq5mFNHQIGLgXgnV5
KOlX4wRh3qJUdkfEhIUjhz3/h7qQdBGqUlg2p9HqFKpQ6KLYmmhgPXGgZbagUmQZhZwKNlD3fGwe
K+769/rp2v1V2ijHHZjd6Y4DiirxN73QdrLKUCYE7nUzxtjUkgb8VZHe7Y+VioU8jjVRIGVB/CMN
ymbgjrK+uRqlWD0QKR602kLF9yhXaDIvRbjSuIKZStz9liUl7PBL0vWQArghNntaHQJV14sdrbzy
6dkOKB9VT79bvmGkkbkC7olXk3nzcd8yi3pwxGsQwZh9H1ya0IenYyrKPJpiyuNhxDJLY+uIcVD4
qMiI3mRCRyqt2LhtGhkSB7XpwzXSFbpPgVlSvSm4h1RCmKl/P+qJ6iJLMnOjaYKetWjyO5raThGv
RAvvmhQfwzd4V8eAVtl9/pLd11ppzN3W6WEe62TBoT8l358xgd9G9UpVWkml/bnwMWoNzcPxv/8D
VHxItWsOsNxliiMXQSNn8+qpgdMB1l4KjxSCG/4jrO4YOCz3BIvv8WpMVcUjhFQKpCeb1NV+UQxe
rHdpCri8Hwm7MHTZjG1M1IORP+A/tETiIQr2ciLHrwU8YoX28wUTcDYql35bK5pnqW8L1PNfryRj
VwTVa2Hb9eng2ab+txQgcEE6uB37nF8ndrjUrbc+ndYE4Pg9ZPn82GT1yHf6E7H0CT5Dbrn9qexp
yUtdQAMcky0waM2iMJjlHcHkCIZp47yXMvTMgEMpSaFQhZmFXdkY1+AEPHs0Ra1AP3cdNQmshBjb
ULa+CzyKxbOIlKuOrm3GnavfvEt3fetOcHZBMWgM3+Le37rowlfAQPZFYLeDgeRyieV0YJsOrImb
Vikj+iwehQyTAoK2Nma5L6fd9tOAzs6qq4AnbvYh/kIvuFQYI3AS1WRp4i4zNqsTCVkzdf09obYf
8yA6TZIse6P0cDXY1DoYIkgZA20iU9w1xRxuRsEYvXegj3czNyimw0EPjwiky84wEATTKpIN+tN2
iVIJam7tbVJDBLgfhL0eWcUgdMs08lSNYzwubHGGkK5HUKb4t0XPI1USoQNZ2+JQ3BJCuVH1buwo
jEtWU3EtgFc6lL5wF46L70wS7MgQe4eJIr/6AoNlvy9KPEISfkzMvuWEiDxPuglw+WHeAjsNvhBp
0P+/0w0QD8W/Pkg6pi0PWRnvm0NdfY979TscnB/+cAT19dtgAHtuA69zvpMcDaXcPLlOMwyToprM
U7pE4Z32TI81QsT8A4nu+SeRArxAbPSN+1bHWO0MSiH8BWadn9jN4fZSeuPTmAS+fpwj0Geqpfdc
koQepAKHQ3hbanW7JjnnKLpAUxMSAlJyyIa5Dbv98HavryxvBoIxoDRG8+EuCSCDEVUsP8hLlNr/
LoF06S+pSYHZyMk6cZvNSa1bgvbr7BgsWLvVdV+PwqMgLLwZaBQEr85SbdrdF1DPjzsq6+uO8t8d
XpyHpN4nvgHaj606orCjQDqjwCElWk2Eph6wTnyugczteC2r56RUpLp3sjnvTmiqDwwlvuIj8Gpb
EjWq3ycaiA45bAQIgvjl4oM5uRgM7sC2P5gj697o9Onc11V9hAcqvs9j9pYQ8xm3MXn3pZQzMrx3
AZAQowDjBIwgPKOQW/MlsSTrLNBYnr9GJgvJwuURLBeXDuIwy+ski1sHXD0PZQtNTa3pF/Ggfwr4
ZWg6ILqTcKugNKueIpzE5W599EdTZgxO5SglWeEOtK5Uf6rKbnyuESNqF7FZRbNwAh/erkBDMb2j
4DizBBZpCbomtbjkk77eiIMV/+fZpRXbHWaT5rylXh4MMU/TdAcl1NdWwoU8hDA3eYbsS83u767L
PF82wuz3un1qJ+eVVx37skek3+FY2H91kJ+KJFOXh8hv0GeAyqBdzTrqE+SLJb/ulGd5rHUmlmZd
ND9P480kJ1ZbeAIMTw2lEoQ53sMkXDLApOLMIj506r6YO/EkLBTUDzZ8F/63BVU+Lyrwpj4jJW0y
B1C+W/L7OPHgQpLMqI1vOU0xdDzpxHP0FLx5I0eO7zYYxBGI34Z1MBT54SRdq0NXrpa9I1OTDzcp
rp6iEyae53c7ulmTHCtj3Qxx3M13bBdGm37b/UpMsJ28tf0qc0CbagBa2uWoK8n6fK4bDmAQbRaH
lW+B30qihFUP/cXdl/PuEJh1AqhhTyvwxngimLvwy17jREiA7434mzo948XbvO9cypmeOA59O14V
c9PjR299U1XP1ikYadRZZ9W7hMflllG4ihNAMZVnET0GD0aWMS3RO+8znLSsmDaAwQb9QWdM2l7j
M6wxwJfl/CuakL6V3IyH9YT/6ZxphL78ltUf2cZEOGBCPngIOjEMQGgIhJRDoxlaw+PaoxUMO7Ux
bCkij3wmCTyU0owwly7jT4mwupbfta0o7yCr48wfh4UN0nnsFUprnCn29QDw6Y/n6pfa4CwVMjGW
gKabfTaUZ1WqvsilPUiWTTwNZz35VybBscewJe4XrRdUYSctMIjg5epCmR6lBXe1Yz6VsJPDNgc+
E1H9EQTIV81UE/KuJZiDGt546FzS8xm+sxoeTJxdrDwyg4AK+w3w4eHcx4ZcQkIC17RKuNr9mNDI
ci59+QH7nfEnoYYFVktJQXHf8urY7306g/o4csbd42EUvGg4uO9BeMNEfe4fhsgd/6gHdIsseDvG
WRQzHBZyN1Ok/P5DUmquAz6/EAuwFmLrWX2go3bGi7P+g/4HEsjkkzp40Pv0pufNy60C4tNB5b05
u4a/6Dwz8pMdkBmXwz2/YMOoqiPcq93Quxw8TAh0BHJxWNO42x7KuILvxDNR3R1XteGPrp6+nJxh
QDoBy6pfmODXRd5YwmfE4EDs5tOvG684E8ZSCS8zwO1j/BnGSXfH47gju6+eoyuXmS+X3Ql/xb+l
M9LuFG/twbpDQMgtCX/FqoAS8V6HVSHYA6sjAT36WpZ7JzS8L+WIQ0VulEh+wTOePRvnemUl/CXk
z29d8mXymHRYbXINckhWPq1yG7sUqBtmrSxHoF5ZGH18GDP5YV+HCUalV6Bfkk0WHMKA7NuJ5zoa
F4GPKuHcWJ0XSDMZdcR6XdvxhQNyLkseuXHDT3T8xy0+KQw99a2jiHXU1q9rHGp2+oeAEdOa5FZD
BTmi4DZsMhd89pyc74S3K5WXbk/h0g7n2Idik0vM/70CpOZKha1ICrUiiRFrBvMNOYP0DMTLWwIo
YUZhgffYhp0iLAqYssaO+XVFTQvrILnc810m+HPtlv1R28bOoa32Ma7oT2i4hSvPbjvKKtKbji1s
SlH0G8cHBdm71XrTHobY/XgB8hiiJqVGNIiAK3Y7n/6rNUImiuUnKL4x5ieuFbBd3rF/XuK22KXi
t+96ypHFzD/O5F1tnQIe1XIGNKS5R0qtsJD3T/WOB4Bq3Nubcu23lLqWtdZk6QiM6vSCmCiHrGs7
v+DrjXPbagxNqSicGUUmsbIuhPKJYFHbMxbGZyRdSY+04odbKTioqgV3Z3RJmxdOEyD9y9EG6XDn
fH1wHO3T0QB0awGHPq4IOb7D6vHwStoh1wqh+Nw2mhPzM23gLeJt6ycLPqTlZadGK0XDMHP9Nfjt
QOLOzheFyxt4aEZ+r0VY0Kh5ERiXr+F1mJd7BvvTuQK0Zhp1SbVpGKzfs+NeGqGcigExMJP5QvI4
AFBIljJ96dJFVMDo3mQEi05mMDjGcCzjOBIxa0wN7tYeMA92/TRJyD+CfefPETfXiKrRMy3kJdZR
Gh0277OYR1YWqTvqWTa/hbxwsZfyVgAMoyH8mOKnG+V1fppB7BOd2CuMdCc/2s4wvw58VA0Y5X7i
XV7srhG+chmsONSXfpHMZi/QJwDWjddNSHFu12zYj1yLnBszC7H0u46Ujy0EOwohOl293U7jAN4L
Lu2l8pU4eYJorBoduwC+LW6Dw+tIrbyc5NwJxdE3sCWuUxqSyRB328i47JIMy2b8QAQExcQVD2ia
QO4t8MvmPi6MqA5zgmAWiIhjtCJ4xb/LafmrgLJ9wtpaec8FRhHytIcs7pYFuNPtVnMy8p84w5t4
YipFpiKZgoKPGcW7dx14jQK3JBgOCYMfYdutKihZImWwqAjB74c9K7Dr8NAemqI31o7JjGS798KW
EOPWkSMV6Kbo+xcNKgHrT3vnPmreYiIvICDgGuzonqiSMoeIl0AUUuRZPURs7uu4rRLt4NMr/UvP
QcH8AV5BrAk/TwvGp5UBURZo4qfPHggwGiQrg36PNhAD9qODfJ0yWEQrAm7/nSnaOLwJsdENgAfE
1gOOC8LHyntKdaQB1rbWdKar+dq4cxeUV39kI15rSkzQyplAWYy1psRwtT1FZ/p7ied7/+91mwkg
mnpRK0v558GPIUOFulMe0VQt37Y9BtdljVmmEIMYjt1oBbYgQJnWwVlrp7rCOweqFW0gFt9JfzL6
36W2SnxxQ6fK00OvsAKAsB7V36eK+ecD3+JDoSIpby/ofhoB20UXZIu97Z1PfNY9qWtoM5j8lCbH
6T29QLYuodP74vXFdlH1iorT19cigsOoQ0fpWBz6GffNogePhnN9fCGWi+/xDYwRfvrPCKUTEoLg
o1otE8t45LZyqsal2t+qb82N1h33qk2serdnfLW2qZ5Oi9lvpE3QVpnSyp/KlPBqFyLcDzzK8745
DgfH4AYd/+fHaRC15ZPMgm/GXiN/SAKqNwjgqWpTSdA+zixYsWMpSRdXF5jAAlbtQjuh2hug+9sr
kEGZOhBHtj/UiQVbnRBV1ady/tzcexJe08c5zaJgBZItWtmXvQf0s3ZgVzZTInwfrU7sMrRnz7on
gGHvLAtb5QbvMV4JUWfuZlCXvir2mSAP2Rdxz49VHylcRgZNj+8Y6QWdH7EMJFgk+denvjNRQmj1
c6Nfwa5k9XbLKVIv/hDcYKysm46NQtLNw5OSn7uf1MeRShLCU8ezXsIKrsTrrRTVdm3voZo2Zy1F
PY96tIawoRpHpE2Skzi2UVJG9hac4MBmsTr/4MCLKNB4ljVNAeD7aP1mc9t72P9SHvEk3PSmpngE
C333gh1yOBi8nD/exMwUOlNqSynETh+0H6IXHKwlsaqyutiTOu8yKiUHrf0spI8OvqBjiq+DAE9D
vwHBr7Qx5/uekUCZWm6xFg6lrGdoVWzEzacW2ZXw0Y6o9zl8XbYibDeDu1C1dhoh8V9Dqe2B1M4w
QyPghf6jqzPzNCq8OlZ3hlI4Khm4VMTEMjXidv9kvR+jq6SDQeSe1tyXAwlQv/Y5Gl9pZY7VqC7L
lf7vjViIYcVY4pWJoHrBKx+6dc+zJKgyXXGrcLzjPtzdRyQjopd535cDcKMJFy1eF4gIseh4q82b
1K9XNZMJFR5txjw6H+XaenKJZBVBrS6LsVT7tYZrCJ5K59o1kyutNxZRdjs5OqRqmrGIcyhKMet9
0OiCAcURPKMsHZEy+PGZ9AKBq2PZpRO20RgfUuuQdyyhCL1UA3nlmTvFeDBlXi3kRCDvZkk6/2fb
fJzpYisTwhd9AuXd7Dy5Qx/cfKoqnsu/1kTNGNdGGZZ7TCkuFK9MQOLn83pMrTw1c9gxbDUM9lAx
i2d0XmmTg3IUqqq70OS/g0ZvQikl53AVq3dyIUXXet/yPY42G2ZC6m/rSjW3AaMfIHdoaA7tGObZ
5WFjJWqBz/7+wn/fN/QJgXN41gQQt1CeJB5ZNaIGgqr9k+4WrSw4JQ9RVcstyjpWkBNYBYPRHOLL
BfrxJphsg8sB8inwyKjMaEhRhOqOwPZYOCdrBlvU8RyEc7yyHJt1dItdVM8npLA8DbjPOstKkcV7
K4kwWagPhKvN0u8+ZY/NBCqTZVyVoQSIhUfSe8ony41tIu52fF87kjdbbhM+HuZlTT/DjNR/sDty
JH9y61vdOEP1etDSxOCUl+PrXhWBs4eXrieoKO5kptT45+SchPCbVXSkVe3Ea4RTkWRI8whdWw/F
Z9hZrbjVKo6B+AVRiQ7DmAEDhYgKTFworOLDN1xVohh7ayj6uAgQnxhF5URS9PjaK/9WPh7Yb6R1
BT1DuRbNAxzJV4qOd9gw3YzmdQben15c0keC/y6c2aiAGRygTVjhSJqydMn6c/di2ajrIqDwdmLe
C1aJpqiC6VwtZn+Vmc9KLk0JqNQaKfEfMJ+NQWLjxU8f2qVRl65nUaQA50xHx9b/VF/KxgntGX8I
HCqMojp9XV5FZwrJOUAM16ZYLpheSpze4ybVlSgYjRDvlYgONefQIMRUOfLwl1kD3t/tMWlrTAiI
RTW0Ot/t843v6uBLQum10SxyESqFxBldB3ROsoRYM6qur4CozfxhWnl66XN6KAxJ29Qol4jgw97z
XGdbjHbIswELw7TTdaZgwOsSzpraDpT7PP00FZG8YRzlSWbV7SyWWqiJpuag1Knb1q8cTSwEg712
GKD5D2hLl9hf+0iPdtzB56gtEWpjIfeKjqw8bSn2uJRnIUFXY5rRS1wuuf5B2DkT+z+pEwdtTFdb
J6fYlbbMTnjyqUzWrvKMUnUMzQ2EgAnt7G6VN/o+hdV7SUhWQTRvSGI2pnESj/g94VOSkgH1Pn75
B+j8/h2rUHjlZI6qXfXoDwBBOocb4YvYSzhPqgLtDa18mWZMlqp3CN1KmQ13aVrXw5Q31rewXl1O
m9y1n8+9eTK6UB/QOuuj5Z0dTy1P0SuOQuvRHzGb83AXwK4EzF9pwzXQOwSkn+pdi5Rdjb8VEvB3
C9Z4zXDzAzGfixRi2hpBdIWbBAgfaLXl9uoE7gizmaEtJ+lCNRBaidIcu6PSNWywo9w6Uj+DjDZd
fZPSTKOQBgzwF832A6SqBnf//2q2ppfUc07HgmH2lvrblAbWsw2IVWhLDbsZfVK3voJXXQSBK0+d
D6oHw6rFCwBbxGrBpmRMd2TEOFZMT+HZk+FDTwBThcfycJEVaXq5sLz/KRFf9hwUKCCcroJoznR0
vU2xOXSgejQHnwNQvkfLnijnn1GRFLXw09vSDWOfLki20LEhzsAwXvQspq8NZITONccTLozEJqDl
1Gb2EnUB07wSqm+EdXMJZ7orAijN6qfF4Yq9lbxZN3DJ5jE5nEvYvySNXP2mYb971aM8io7MZX6X
5VYiZitg7bILQsQSlfdYXeZEf+eUbfTN2hq9KHEzzZ793/LeGwdF3xDgO4TAviWW9JnN28QchdqQ
HQ/5iU+wivHnJOnwLcjDEbqjBz476gGnUykZ4CrEqgiT9OMAuFFxJLk0UkAjnoLnYdGA8GPmzlSy
ZR/MYSrOlBoQQKJyy0N28dQx0WPyecZ4+FN1rzSLeqPSwOvmVylRsfXt9gnK/Ocs8JV7yi8DRo7G
z1bb8be/QslD18Ep26rmgVU27uWnjBhugkrG9EvJB0BnzP2d2fuQnwO50qAOXPCd9lFb8xjq4Cy7
YXYy2wzz3xw248rEMFCvK9dyH6KC4GWdkKiotKCrpHVHUxleZn1zRhIembMHGrP+Vc+6CsRHP+s6
677A9pvnwhR4dLPJcOIAEI0bYK1sxmDl+L2AAj96ggBCi5HuVzIxFMMVacJ89ejSdFpyuXivYk1G
2OKpI/DNVlKIGI/Ku/J2jIQvX3nWkjVioBef/e9RD0gmKB2Zk9npHZVuN7mncRM5vawSrtlczWX4
HfnbUgkG9oCVKs2JSHO0CTqWJVTrUC/KI+hjeXshifHIYBUCgQgjRmW6KD5Q4n28yrWz0D1xmHyu
PP8WPz6LoO9rccZZ7oHAVMXbD9vXB+H8BxJhKTT5u73b5J/FfPOmrwJZt33wTZdB//XDrY4v0Iqa
XPvqEXGmjKYOThn6xcHvobkJkK2hqIcK9opXcSiVAbmzKZNzG5wX4IH4UU1hLigyWJVlozD4s1pf
wJgjslKMrESycou9bMgiblSNxt+cpy3MQhnkbRLOtAKsuTkPCnNWHXJ9ux6m35QJy+h4FNdxmvfr
Zwm2PvBGIywYsmBXFfLmLmEudBROIiGe0BFmCoMsDJDu0EDq5w93qxWWSK5slif2ADu/kSWyjJBc
u6n+qNfN3X3r+txOh7BhqhwXLw+BvTDgSJunnSUswWrTx9Ff/zDPJEONoeiK316xTyYOMkcg4Zpn
c8meZlA5OwVhSjoI5TGZZILkmjRuyLVZMMJXTtQY7BB/dZ2o6opBRw7xUBGWwJGhJgMWBQvCiY4s
WxDrKPtKA+mdjiYHecxL+RjH24x2gwF/HANym/IwcUPiOfPhdJTg+P41Heqak1GhlQS8ZnxJQCfi
ScJdXVjfCzk66kgfI/qlKzoTdHvlC2fxTUHxZqyIeT6LoHbR+oVl8SAKefq//Uxz/QCTnKyU16kD
PFkDfIuC5YKVhp9kpljJwiJkm5FzVk6CN0oRtzX81tLffRR2OmRehjGZ3MhyDno3Ons1Ddx0qDOm
as1LeVi3gBy38bJPm4UeUcTjpO1hw273suPuEOO2dOs0/Z1neVFtXJBdSsGqlgrdVWlKQ43O+rRn
/R/Xqy2Mu5AGlheldffdTJOASJL31qn942b2XkpnSZOBwZUYpJ3WD1TNGy0eQpSTIwoi9bS/XjP5
ivACDhAA/wEQRhcFzUsY5NTxb2LybTDXzd08a1523w+RXeGZR9GKUdDNK9kzg3XJiJClmEcWtwv3
iNGhT203q0sMBwHnHTD6Hqu0R1vGk3PWR8oTJlmGH7ucoQLjp/vaPWXgfZwvx2XU4Ihk1xwk44WF
CTv8kdcRvSpsglUw1Wzqk5QQNlAqvTuyH0k8YlH5ucUhezvBrYAGdCDRHyxfQUUpNg4laD4WB5NU
lbVTY1XekxAYPDM5mxKZw5z4UImkbVCOO9L5JT9daStUHisw8UqXsikDSGDNlZy7RVJ7O/uW0Bni
sePiOq1zcxoU4G6tkPUw+0GXrf3XBwVMv2AcMqlsJMo+CP4dsgn/eZNgSXCXEK0deae02iAdXhYs
vQ73PJGQijBulh5HlSqNTOUh3+n2KTaKY45SN3WXUxmiuCjB0j9q47Q6gC/hshxa34paKCEQ/Q6c
nKF+bWWWHMbwvCsRe9oYLTsZmV/3FzLB2j4ArR8Te8kivqGDqIFPm0blgZwvr4dxD+++KryZsvB7
oaOvVOkzO0QXDLrI5YHcK9veb63OghAof/BihfQiUNIPzpm2do3EYIIAXJKyCud7FktFTmlvuwMn
pt3tXq0R4t+YUCbNLTNg6hPRy1LmW/xdlDw2fGvjXScJoKYkSEfYFORajJq2JCvKcjIqRIDLUsHd
z5aWcN8eoiGi0g/j9VhoQuBqpoKjw9ht0UUuGY8E9Rq7Letc2O5FnnE8W4bgdxTnyzR4Hr7uAw60
Uy2/HZHV3PMekd7IRUBQyBy/0heWoj8FSGI7pnmmmn0DMByeyfZKtye23Lp2WIwY1Lu1c0rcV0kW
JdqYGIbNrhz5Nt9hIteGXME4NFUe4cVSmzoAHoVF0rDeBhe/rMnQll3RyBWe4mLpSu03Nfcv/dFZ
haoS1wq2X/EiPu/gB100qa0Rw1Qf5ykSyxuXJ6n9WMFSrkdfxolqngH12hU5Rg4NMizJgIvEMBxI
Cdwfit1kb4NdYsbCGx05Apvl5uEuzeqQLDhv1v79ue0Dw3y90PHB/0azbKq5aqtyjJggChyVZRbY
Y9hxXuy2LUZYBdliW5oynFqGWjdNi73hh2Uhet+JfCs7KjNngnAeasCF4dt3j+3Ni7VyBXKka0n2
cXsvsIbLBOfveWlWcKqqmKr6qfRHRX+gWTkbQkwk/AcEycRnEXIUUoPRzAER/XItcn3GIR0IsFpO
2yyQ7wjxizuBAaw2wN3UhJBieI9q1pb8RKciBVaRoeSsc3nDe7m9NKaEHt1Nx+xe+PIDbnwCEtmL
+1qEqiNudvd78/+mgsQ34E/Zo3H9gmyQKB1BEvvus6Wwt7RgN0Wd0xs/LqIM0o4dk34x3mcFwSNi
bx93g0lZnJTCBLQZzHU6QnI34ww0t7LgQ0EoUJYj7p7ZgaL3E3uxpzMqFOpiTt0lrPsH6AnpEdWh
3gxIvEazqkU7H/H+p7YnVs3rCJHKe/iwltUkHzMt0Fz9MwbZJh3rJp766IY5mC9ky7geVRJu9jrT
aPqv9l6DIyQ+wgzeoJW7ofExAuJ2ULj5UEj/TthQCzECcvHNtOwGnIvx6OJFgfJbwFEzsLIqWTrq
mv+PqcNT+NzBndX157E1iJhzUGHv+xb21Z8spT+AVJWncJCtC6GBpdPc+/QNbsadvFtT4wqiQE1n
cFBfyygIDrferVWfFzjzmBjwxSFa8jnd+2lhokfqwGx036/UQuPicCq7wbnqiRVR7amvrlnZErJi
s6Oua0qybvB8Yo3KJhW5UvCqeCQWLXmp1nGRFloWs6rG/vrxnv8TTeMu4T/eTYmq7KkXQZQi6CUF
RvjIJ+/kR2aHKXu9fMbj8ozRHKnRl0XeNf4d/2phsyDdOq77uQXMX7nsCIQGeyUNIvHo1NNWZuNi
2qALSbP8Rl5b2Sqr9JWhZiGi/veOI71qe+Gk+1ab2qSUeoXXz433mY1tG3OIeEi5W532g55pZCZp
nRBPAUZLbSfO6bUX+w39nLbOGDhnuxYnsKjZIcHOR+L9ItLYk/fxXEFXJ8yn+Sp02XHO2cztH9vw
CAZp91uQAtZuAQBU6gQaS4/z9XGgFP3AeX+TVU031gLr7E0XOAswEOyd08/zy1SRbunpUVxcWjLO
2mzeY88KfAU65f3igC6t0IgPPh+Zz5b1wwn13j1BxTZCLk/w2HYbC/x3RAO2YOhuuLCJmQyNssWD
u4/2WU1t2O1NUO3TT0qp5HgzW5pg18g7Gfs9TJNGiBf1ZsmRai7uEYh4h37JWomSftmISWGuzJu9
D9VLSYHDzRodriXV7re8lcPB3MEIAPC48XUPn4dG3OGpDLPLb7bCUQV8dfYDyYVmgiub94JdreDj
SMFEPCqbdA37q44HlEtGlL0mxdVDc2+1DAFa/lBPiMANXwi2Cq56JJY3fF5vfTBvjdIWESXIvk38
jpl187PxkvC3sw4BOLPoSuRN7exQk1003L1mb+nXyIDaZrIC1qksWbiebTHdKxJeniIopVz2uPS/
KxERyxEjxbt351QfhMVsb1YydA0BJ4NtzX5eU7kj00mtvi6n3TUymPtxfH6wuKz92XMV+I3pTgOe
ZGoX5VeJytS3ud07l8WbaWqPyOFwNCrCqyslul9Z3OI9K/zrmUYBwobAeLRwKHmjwbzTn+N4TEDP
l+gNuE44FUZ/FsdfGqW9Litl5SrZySCQd4v2FfJgH5LTzwSNmGTw16uMSjLkTVRp0LieTgYZ0exJ
u/BALBhuNJckKQNdC2jyN5n3TFkCAffc72FDafC4js4F6wikBDXLsagG0+z6QciTLa5QycJGFEPD
RKUQTBei9JTbp+2Ryji49kcMgnFTGnv8fDrqAfQBG12E10lNURsbKg4Yr7dL9USyaN4WEIJiBYBz
W3WEwRKopqGbySCeDSN2UH553dcaUQQzMcboDClVblM8pLWKi/1JCkwt5sgNC5xoBIrb0eMO/yiN
jGbzSCNBYxcca4aF/nH2tZxTf8p/Jq8IMHwx7W2hims4EawhJydSzprECdvhZOX7oW6JtslRWaML
298aFMwI21quYLPkTmhvhA8Me9iuBYS1ZG7jYijbtq8NQaiQg04d3pafnK8JKyowKAGoOFIt73VI
apSkcKEl8TmvsF2zIYSKZq/ZrtDaozFsayoxh6VNQltIoRDUwTS6WcEDdkSMrF77J1OzchO/wyxT
w+0STVQz4MkkVAN99jjEeaiSCdSOFOyX+TIyaQ76RnOYp4rt/OgmNZ/RPbn8SQdAXMKpVEDR8EUl
eEqsWCAHUCF22t3PrY6qvq4ICoSYnqdRqOn/0aObuPRglHzpeYFiSFCeXjRKsvcFENnNFAkOcDjS
O1NOGfQ+Ino9SxLxySw9oHV9HykEEDOYx2P4Z30ebQ3Ku5If/+VgplCSzg9nryrSGo/fTGk1erHc
XGXSxDhH+sazZPsoiaCJGgJSrOr62um7FxCPokP3BBFbdF4F6S7dw/MZUH3eRcxFqErnKnhCMcML
wLEiuzjPsm8nZj+YTBHvE7DrGd7frk+D94OpYrfJ5FnELolbopHiPW3yBJnY0oZsBVA4I+DRdYj0
VsMmgJ3Ps7OAcCtZ4cYV7dSg4a4EF5MvBS01zkedzY39+JPXTR4aFlLwVYZJ3I7sVTQ4bRcPk1NK
PNAJ45kZtICwI7nmEpDz1ZKKpx/QrIq4O8bRPV/lUm1H7+dl3k0OgykW14TO+1L2JQYsojWUWtAM
K9zzi3xYxRYc8vpk54MpQHSf3/B3sOcRRpQ8SkxZfqaR3Eiy733cOK4OC6x3Do8o2qjzxeUgp+sH
1Ql2jcocTdGvw5fVlKT3Pc9JHZ8Fj72B7nBInx5SST6PL2kJ3iscvk5mv/VMj/pTUCNV+hccJzf7
xPsBtUIl7KrVNvsh8Wy5SlQQd2vpyHjpf33at+LSzLN0NbSwIRtPJO2tCX4PHDOOHD0jubE0eZW+
F4BAZftNZli1UoaE5ITfMXgrMFGIgGb8v79P18Rp7d+GFZ3Ljav8bNDAQtsdtpRLqS7NJn+ab7z0
ry5cn13eDyybcZL23shfu8YPzedPwPH6PwVBj8lZRCPAovReayxPjf6v4K3rnyp/ew7WvN44fWIb
Pp5WebDWrCcs7WvomCIRAzAFmygifMgnp7UsNKXsMI5mrdvHzT3iUHAi+2p6N/CfHD+DX0I6Q24w
e88OdLzCQQu6eU/5BD8LTXWEzRzl+aIwfBwwlKFY0eR3q80ymInRfDnBbvm9NLxEsVY/CRTdiQKV
9+wArHPTQcLNgsEXvLSBVwANGlbd2t18fAaAHhhayCVzm9/HMfLLa2LhHA0Yv92uwHqFYGfifjcG
U7dLUTOAZpprFvzzyH30OUN2ynql5CULoYgmpVWr0jEpvShoq6wDwzx7/kpMPm2qh5TxsKlpbHzo
SG287nR0UrI4hmWvPhqoK7iKjNV7YQoDgUfZnAw2nk6mRN9quSaCsehehF8jWllZmjPPKfJuXDW+
q2Kpm4Yn+RazbborqpI+7rHz9lemCrZ9KBSAg7ItBIuVwEuSzYTS6YBnIbr/ea9W50Pg/0ANpbVB
y7tqfnb9zEM3iaXji6+MYoIj0zj0Fb3nqRMVAW3U0tb233veBJJPAUQYzk20YOHZIUjhe17N+/Gm
mYjJrv8DXieatRb7ODt5TOKrLWY3hhoOqAWUlzE1MtEkRJtip0OmjH57oYlMiEhy/WtikA3xTQYX
HdfxeMhqrdGV3/U5jTSx4pDy3aHqOuIihA2t0y0jYVZAJqpgKftNmoLqXzrVpj8yn8+5v18UQ/hs
IfGOpXiuZi0xNqTCRegc5UYzioDXROkJLkB69qEDYUVCfcDx4una7cd9z5xpaVNmqcNbnWWjpp8r
BwrfJkn9+d/93uZKwpA04C4XWNtLATzc/4TyPVqvNOz9k9NmdfsAlTQPyQgehByXrdDwZZbuS08y
GngJ8/AVIQfNQy8n+T6COWksmJe/Xic3KMpngSsiF5K43Ylb8ikdydoG6j4u7h5wZJbc7AuTRdYF
E7W8S9QWiaLq8id7T5KJHp7xhkSosjTvH2ibrZxlGKwp5iXwO2Kyaj2oIIH2TQ5Oe+uGrn5iXou+
QL3RQa2Z8QCpH0YuPLylpRCXwOzt3Pslr1VHxOl+8pRRhKbTjnQ29WZU+R7BuT5XCPIxVY938ZE4
HJu//V/yfniXaKs3ny/cXv2efnA7ZdxkJpHftFkZMJI4HjqJBoM6R7qFcByugd9QrFwV5b4q6Wpe
LcRtXqcoH3E2TPNJuQVZIvuyIjF3hm7r2xjQGjIBePxRAsrz5ae3rc3fWKbfhXl6HvoE4+5d+KKa
Do+hreDotwKfD3u1DSxaDxbqEgyJ83Y/EgLsynAojUE6GSrXxBRLFR3yWVtjKH237mEeWE55RJP3
BX9W5kVjYcJGE7SgvfsK0CfBNW9cDZcA0FjGuyGwfsoSVIeL7+5lFhP5NxKdC6pBrN/7F26O23l6
r2FvRB24+IBZU2cN7Zktnr3U4g28ewRa5lYgLKdd+sOauVv1ip0CzP9+J/FTZAeyVW7qfZ0bBDCL
Vtec29ps3hYH548F+2k/PKH0UuPZ6xnNPisAcTFFF2Qip+UJF7qwstapCclcBCLSYnzNvjBTNRQ/
Kshb3L32mNwW+UCmJQi4p8TXRaShkEDVy1BmfJ1fNF/UYv424eT/RpmA8uPgZDJkBObYcahP1Clf
N8lkoZbRQDpiZlDD7oidIIBahb3rc7jYfubT0wEf7ZWofDBk6dZ0yuvYxJN6ksZdG5iL4aBHyABG
cOI7XgWK0LQbY7VcADmrhQx3uZSgNBdhtA1sk6vpDH9flHHAKoaoIOFfoswsjL1IXD2hRb0tPmsO
3SCABaDXzMCyxPpFavKj+axUoQD6a7z1gzup5pcBHPSG3cIgcHTqEiqdFfT1epRKONUGIINrZd2e
WLf6ZV8WfpNIlP+z7Um8fQO+1SU/T42o63b0rBe0hEbPvnsfdU41peSbJzhAul1myPKK0lZM0cLw
jWnjM86Ah2Gy/Pue9BXorxiI06lRAMfTdQdT6dXb8a+PEXJA+i5C1kKIJ3jiDAbFCkp2spqMbt/r
Xon6kdGV5AbI7W019SmPAat9OxlS65W+kZgrx57gK4TTPGVUpnrGtmqOiyNWYQPe3FH9Pz1aBRgQ
bCKYFgjJgqoOPcr+ZBvqfYtY9y36o/rN0jv51I4fhUueeZqRB9FUozDDGfmzwDm85g0kKTVLPStZ
yRFCDfT2YLeHE0cOadBqNvr1l0TTli4sIo7yoSZP6Zdka2hk9w2gCIIP2j7/8/bUpSzvxquJL4zR
yICgDSFpmpZk5MROXpPsaKo0uoJVbPXWx9HlX/1cAtVK0pMAXDN81APYwYIH5jMjjs/UjS4c1wj/
bTA9KzrOOCPqcDOwCETFL5wcp3XCzqG20UXtuNvvWU52gSR+21DIeKlxVgzy0hXgRaIYGOCKhudT
F+mVJNIVE5TsYs9DqN4+m64dcuo8zPSkvUmh9uRwRpr0FNwDGrppw55VHdsvF7o/kTWL3vbgmFuZ
tG2XdCxAKvHCQbnnhR55c/ejRhmfKqZ9DWZNcy5wVIEVI0quQZynHe/H+HLZY9SUKcW8I/XHU7Tj
p6gK7aGg+HynuaVRFoawadrKz9ERzHt0gCJG0CPCScyPpU6+KiwKjqnIbQMG1Aop7y5jJg63i21A
UNq9H/7kc2SDeYr4x81Kszwak/FfRm8iUY8sEn7uf9QvCGDZzKP/JwhrE1cM297nRE5Zk0TFBmrv
LcbxAQcyJb54u8M59MpS597VQRv7jdJnIkTTTSRk1L195Ltc48I9j4qMsOHd0RsrXmhqTUMngMl4
4GhiKzlvJTYLIdsuyXyvHADz6cO9TGuV+Fml9d+kvhhvZN6IecsKbta37q5/pFxQsQcdxLuFHVum
WmKsJn8V63EGocXfZTd9CGsVb4Q4Cl5e5cxRWSxa+/8P2f8HdAOSk/Ye47gHgje2FCIwGCYrC22x
E/vah62maAOfKO/8M9uVg3uZM47a7rRbfIVJrHBi/vhZ0Du2tcwZb4lftjwJYez+NoBy2Jo88WkL
rQq5ncyvA8hGhZsmd4vzakV7Bff9AY+127/Pa+hxmnHo14yQCx8+OpFXMrKBJlKdRjqry9VjFYrg
G99ImvsSxRIrKKabMtB4m/yKBIDpI3cy6dDcxWzDw68ZFPukMoHMW/Gn+s59FGgxn2t7tgwVPfHG
IHgILLheexbvx784WlJaSN4877HR6OElqdquKQRUzenXNPZUqOTnSqJejTJJkVetOFrxTUr6L340
R1BkA819oOd1JmM532BQehndJFB7td5OuAjgzarFoAuZEMrpteDVlPPCP3Zefmb44+HJZ12Tlvtx
b1YDTHkK1xWUwnfMtMjhU6y90/D5nL8eKnBC8cW/YS9oJzOWXisWYUQE+V2ueXAu7qtTDgqHFjo4
VX8cV52kfgQKMzzeGvxcgMMNY2OKXgYNvjPDPCkf/tgmYyVXhKNIZqeA3PukCEmN09rn3l4tykUU
WNzIdHpSdC6fX21uRI3dHkv17qNxxbK6OSo6KadZJyhEKokGXcIVD4Oe4e7+MiDhBNK/iovo9+Tz
J6OMf4dDM0uTVcVnDdxE7vDei42mJspnI+FnWFElEXJmc2R35qLHm4ifi5Jq1njYoV1iyED2Mzd0
XVOwG59d5dMzzmO8qfi8fEEy9BgDcrqGE9zMnUtzjo5LFn7gquWzTxKJ/f1WBpNeZc49x0wlfm2W
iEgvpbCyEneVmWcbRO18Iq6nMitpywd4g/Y+FhepHLDgV8nRFXcYXzUDYMos7YFtnEi1Ooo72qrL
4p19vnNWGjWaftqGyY6Up4EQUCZMcnDPTLZr7vDvFzoki+8htiDcnH37yd8zsdGZw2nBafneBKM7
s5VwwKs8P3PAUWwIMQjgdYc0Dm0JXN8vWxLYld7+pc0Tm2pmVDLlo4aDKGtOsUZV8c6tgCKN3Yqs
PNhwXURSDsjXqeD0mmjeEk/hBwlk55CycuNkKU2cCRwdKfLwTLXKwEpG1fWgRAh0itAEisqG0ZBU
gn/500nKg5CDGsH3TG+eX3Yuvd8ReV2AQk1o2ZmlJgmc0OiCEuVBGt7QSJBzkXNUiWwOqlUynFNq
uL57Hx5MZZt6m2HncfEkKcUE/NIXOAn8Vj9qu/5MbPYPFO+3ggyGBxA8DKJMSVvlHR4POYNwhLNY
ngosvNlriWBmPevuiLbKRZhn4tQhs32xjRfpeBPxxmwb7uHEZMyxTmPi2Gz+oQfPebkDxAogOw+F
QSMvL0WhKawf152RTJUTmNmA7tCguQPq/wHgpNNJY17S7ywMdQao2ir8Lw5mEeurKJT6C2jADoJ6
AWZcyw9AGGyt7EQ2Yy3g3Qx4T5DM0wFsxMkTKrNob9rM0sALsptQIFYjT+NKVnNqNCaLp6Ac34GJ
SILiGBq47MCfsJzhLYBPxuUtF92oW0uYKHzB72O/C+m1KWQvebQxqWb7av2VHEZZc/vuAYBKHIG/
IbaJenLJ/vI32iw9JeU/LhupYsyozJg0dqwOLhW9mrE+qq3WynBtMbnt9U7KthhUljxlMCsxmC33
/q9cJ/5A0876cjPqvXb1PdYSpwnYBrvx0vIqMMONkt46eRqspgUmHFFJPkKKvFj7podrN+8bKJad
LNfDlZj4UYVNzKT9turSrDVMnqn4087uymJ/JHo2KFokOYBy+iMIQD1b3q211D7gotPCeRj9KTN3
jSWJrHeA2P89tVvnuy8FNzPZO8WHe8isFuPL+y0T9EN7tC6gsVAH4cHQa+BkeJ7bZLWs57YlrYIW
YKXHDIy5Oo/ObeHubj+QI3aQaE8tOhyKCXIvXVKmyumwKWYA3F1lpizr5YLZ3HUrBGL1wA0VUTAm
p1zIUm7JAz0n+Rx7K9amOF3WoCLBMyKAGE4MfsbAFbK/vAezD8bO/k5q4WKI6glYcwtfQVLGqFSX
KNHafOVlDvzV9rA8Jc30VtwiGuZSzXyfE/fmHsy8pfO7gg7oOFtDKl+dhVytmAoSioj4xuqEZtVo
0CW6m2aQxv+1LzWZyZPi4XvDuroJTD+qS7K7yK8R0G2YQjN1XWFXPJyH+nW+ITBX6SvzTLkhnGTq
Xg9hc0IrFd/DD55iEbXQsnNZx1OEcba+JG/TWsCz/ljJHt/QbDXeiRemSjqzohP67DOyLM8fKDZD
WgAdXmy8F/PV4JMXanxr3RRKxwJHOQ8038m/EfikKPWXjFqh4zU1hmIlTmV+XK7s2t4k3pOnYUD1
YuNu6fdHEZO9lXVhJNgt/UmDp1ZE/K4D147OvEBM5Hhhs035604FMaJb5oQKufSjpQpnPHsImoDs
ZjCOR7uxCEbh5VA5JLUCAKyivgs9yUq4kkCdRPLGyHh1xgvTefu68ysGaOGMM6zY0C7TAqRnEocf
lCOACnHlHEXuC+3OgItG6wChtBjKxVaQiCgU7fsbCx2mWY36CdYYF8E+wayndb5kZSZ0z33IqO00
5sSZIxh0REPL8odAKz+xbw5Uxucr1hynXljVUUHza0ipUmp8wO8CxKVtcCz0losrVM8RKd2ay3Dl
3vMUtewbF6YT6Lb/yylQMLei+iXIMfKVME6deahCbe7kze5lybHMb7UOoQ+Qk8Ng03iJ7ft8G24Z
LpyWovb7aymQN28wsSF2o3wiQoaHvfoV6vHlqCLZWKatHOwCLuQh1+aOnf0hpWKacjt3rOquYejA
MJdjU2pQd098fUGmArR/yHhAQhCWiyBkVSCyOuGNu0Z0IaGQl4S4rJ2k39iwCkK5h25rUEqiTsD+
Snr7iliOQpdK2+Q0/DWGK7DZos9/KT5CibICnvfihdaO0T9PXLG7E6+gaYi9yheG2HNRmuIPvDnF
+2Kl4HlJiq+i2JbiX6iKLtmXzmp+wGzXhhGZdUonZqwSLS4b8/rY6jXkZn3voFzQb+rO2TYKQVqf
EtSL1x+VY4Czqv6ekWeDYrbhAjEXU2NRLr1pOSQgj49thAK3oX0Fx0E89ROksYjJEOPZ/vmtUbiK
UZMqYE2b6B6QmoyvFQcBsXVjNf9Sa6pDS5d7NaDWTV9Fq4eikgACbetbOHPoD7okrGacDzgSH9iy
1JdLRJnP6ek2tqunH4iZigB6hY2WySv2MJdJ9NLvVZz6khdorOw3/Z0lZKYAe/tDtm3UESnkqgqB
YQxRXqTtL75raHSZa2qtQllarq56AvVZqB/e/NpN3EC/sm6sX5IL04XRVqbY4LtwgnviB9237ff8
yXt7kD8aBRP8c9EKH4FdE4Qg1Yj57Dr17B6dXyg0LL3E8roWdzh2gBGBSH5LyxzXH4GFsXz+zpDc
IAf1T6V3IB3gQZf+Sn2tdI71TeG12QDd4rDCnbQPKcB/rcDZZB9prB382BFKy1pxSKeeH+XrJxSU
kRS7g7OeBx+WBkp8NzyC/dLMmECHPk5cACrVFW2I2CgxkoEynx4VJxo0T54paqQ+dhSFzuKA9s19
OvTp4Nqc9WCcjdLdcOpS3O/1KWPsqWQft5RDCO7nst/x+A/0qTxK8R2/D9m954TTCFcndi/pFCH8
+d3TuDWvhbhPj4hKXVJE/HmCjqPHOpdY/uSwJ1DQxFs4VT6ZZ4abWs7EOOG1uignNAObLIoiX6GW
o8FL/yZuKO6gRT3s/zE3pWmGGX8Gyendulk+PEIFhVafJcl+Q+aY2xwtywgno33l4ipcL8ueldx9
hRfrv/Lr6qv9Uj5HCofIFOmFiLfe5aMGZL75WH+PGSbvRqvfJw7nbQsZAp+xpUQSLvmnyYyx3X4H
y1Iv7S05s5dw7D3gsUqg+fO1DGVxed8u0RsxUjkBhFlyg3hD1/Zo36e3SIBcWJ8zKP1wA5EUSC7K
/ee5DXZuw8FOKii3hd8ZeOlBZRkgDtzaNkzi+NQUxrqCteZnCfmSz7jqEiQ4NHGGbwrJaF9QWoR5
ldqgzycCNFe1HDxlh7CNmRwChn6NKIb0d6ClMbD6VdwvlnuioxcAiYWKDL6LK1G6KAObemLzb51a
PEzerJ9L3VaCZcBZ3+K3dBm2CceCgdr5dUu7Und8v6QlbXIhlFy6VtzDvyripkUW2T9x8CHoOsh8
LCcP0QwCuDVcu/irStxo5JypL/dDkOtOwXzaVSNeWTONE8ViDD8ZCrtn/OO5+lBAkHwjxvEl3m/3
ip8VCbuORnBUnesCJA7vm5D0Soj9MPuq6xwB82HEs+RGgx9N8j18TMuGcnfUoYIRjOcLW0oC/qpN
+WcocndlkXKV0SdfYmKbI+o+t1sp30Xr4c0gBq/RkV57aKNJ7k0awDdZkvnVWfcxYxgHk3fuPWOX
lTsmrhpQlIxcpYM6//h83su4NWPQIrSVBag1ZHkjb3qjuon+lAKInme3U3Tx/9woQRKvF0m2FI1e
/s6X1ezbXJdM9TLYnGxuvAY1M45Auixw8gUBhDBfaofkTHpOag0xmqpRkgpE5bOd5MlRuH5SZ/g9
y9Ab1UIFd504OogatDks/uqHjDA0A7PrqMCCQbJUm0LzGQcQo3f+46mTk63tGBVDC76IoaGYp1kn
+zLvQUYUhe0+W391xZhuRLYlyajqtVR4rxJe1oyfwlNaLVujqVu9mXxvF4nda+T6lFDZ+xg5mvlU
GcOVVtJnORuuwyNOrhJ3s5qCqnTSRFlpLAM7hOVe9x22A+mjgEa8ghxYmQ4HBedXmiMJiDfUVEGg
Nr2zYEM5tQXCQf3DqRO3oE5r1NY69dZeLD/xAstROOwqfNQ1lOepU9bNO8NtwGVzC+lmVwjjB+CU
MB40gMeu5NpuV8hL5CUne29ZcOpf+ij4SQnuxHVwHGTySFPbWtrTmfmqqnDCndN0m7FBn8u0/tjX
mXbPFAHBRFBtgLGMA4L2Ta4wgmFoIg0K1zXXDFubk+7VF38pDoZobatjvS04DoJqPeZah9IGffdC
CpSMEN/BoZcwPc5/Y/1xt9qS4Q2R5yekeGhPdJEBt1PUk+Brhz3Os+r7eT6D6nQ4fLcKDk+NGqA+
CW1ndgytLHgdpFA78RKON2Dwc0UGqI/Y2PDBP4nOqp7c2BJXGDWOTl7Oh6RzYj6hsgf9hRdWbkv8
TB0Xgwk5ZFUu8Py5KPfZkLH4PUylsf8hl6EXzU2Ugw7jU7HdSXCv9LgOiV0TCGas6ZzzVV2Vp/Dc
ElcUSixqlVtOxsTvuxrkDae9LvpEysM0MaL1onre1UUVuS8/yoVnAzYfMDUg/OENMFQI9qvmVO0c
ha/yjGv7iSzBCbSXKF3GC0sO1wS4x6fAU7CPYHJ7ulhH+wzZeGMNtz41wPxScNHkL2U2FC480Ciy
N6KlWyr5srEcN1knHuhvApHBUMvTDcyRbD0RDHBAx+ObN1/NBpw6sz/03ks+bGJ3onL9x6oloLgI
B15w5xlhujY/qbZ/gBJEYL4ok1iiqZo4Do3ySKxzHTSJzh0BNg235CnTbRuRKhINS+raMmCGG0L3
nSoELfKKgY3OTucPtHOHpgZWUkQDdUJeeSumXq1H8+Vyfq3ykj4q499ibeNAp/G/Q2M2vBfyt+85
kqxxZJUahnBDERxvNV9SDj/oihEnTv/oRVpUfnjJa7OwPon+ZmVEUPImt/mvHGkcDuAYbbN41VSY
g23DEKC35FEvPj4M2UBItoNS6s3O50gZcoA3dgT2wzGLO9H51MN+zgFSfq8uA+mmmOdxLvK0qohR
endZrcfEtNrQZ6C9Flqgz2Y9OQ+ab3tqF6ZItv+iEWr2b81x+hdEARS6GGgKNUvZ4IxrPJudpme4
praAgIObXesV0FCRdSEpdkS7aRuENguMo2b+iTmr0SM3mFFXgVMjFHlldYHcwj85KwjrAMc2f2zW
q3JBsYWo4+scnlaY6EU+/LsJsia2X+zu3NPseP3kuNqijnfXTORKJyOHhcJhczCNYMuN4SIwv/0s
gM2KK5glVSR+SPwoFQockhotU1d02KnsYyt7PAIX4Sh+N5L/Gym5f18dH8oHX9aWfy7P1TVhQQ5x
ckVB5HGPzaGwChSLVlsZTK4qIQ+Ki9+cWDTBSHxRCwvLE9VkjH84iR9PWgOGri/KZWwHysqA6OVw
uUJWc8ZWDCtdbZgAr48BowVM3oAtIFCDWv7TsyVv6fCtiwadH19XtyuvwG21ki3azyv1fUjpkG6u
EhFpt1Wtd3ZRxeA1zGn2BhXrvI+VK3zVwny4be+hgcqzt1soDQVolTyeLtoROgx/1WE8WgN8Zk+T
PrEBQEzs3PNnz60YZBnX4JLcIbvE41OuISJqcDS6sk+vTprYbbFoCLBVWJoLTEAkuIrCTp3alSUu
yckR2t8/vczXJEUiz0XFHKRrhobHVytG8L/O0V9WPTHC5aazjsNnh2Ls9B2rgxLYTeuWrntHvdrz
nPA4N4GOzVRgnnsBTiZKc4azMl1x6/8EOdBQAce2p48chsNZRKOB0s/ivTMbu8WdpKGS7ex5PHv7
Ih5yCVZcFGYJhAdxmpYpIBCa+eTAdmzjvssMW4H9xIqtjD1Vrt/1fk7+tJJDWN0P6HLHqa6vYlm7
A4wrwv4H6Db0jFTOkHJ8Kx9VrYSYpg9yYvnhlWZ3644CMnlzPMctIgFjnV15aU3rCIy2p2DaVGpq
w+3AW7ycsnSvhuqk/nvpSzXqDrFr7uV5cBHNCN0U0ZhUTF04RwTXHbtdiaXr1JFfraBWyfGDW/wr
Hc0hIvvJGYgrj7nRRQMtyYlNSnPdL8+SA9PoGcbJ3ksudtIWjerPibjBHikoj5Q2kHCcSRXjhii9
eqPmv3+Nz8qJNhkkbquPMhPT+bimQ3yLps/hn1xcog+TXz+7Els2XzakvSp8P1PUflzElhckHf3Z
s4f/zeKPJXJ+w9xbt14P5ThjpADrFBeZDLKkfWxEWw11qUx1dsOKxBuA0uPpPtSnHelMOeMekzeX
Ht0vOQdcGCCdPW6CBOdd56JWfSkdxXU5tK02lBoPwO/ufsmcXUrLW8Tq44FAwx3HBGRr/oyOVZCL
eHTMJmxRNJVIA9R5i12/ywV+/O8Ft5Gu590uRtS4WzvyIgAOtzqa/KiOd6J8Dit6xhGKXkS3U5Bl
PfXFw1bZ+sl+CmEG48AlnSAtfrmV+Z+kTUCvojWnDNLmAxsHm08AswhDUfUIXRBkBLHfud9L+NgA
UNY5476TcPZQ5K9pbaxQ+psXP5A5IDU7N4n9hPEtu5S4vx/5FHNfVEGcNSEXLl4yv5KKRWDoPA6G
5Hqgn93ZmLTSUFQ4aWmueUwXiPi00rK6df33dxjcaAG0Uu8pw6SFKVRS6dNWxv2kL+X+yeZ7/bp1
PGoaZSyK+8z3dwy+FHEKsz2gjTZzGwAxLxOzEXrL8uQlScnHQOgOMDXog99KvWz4Vzyp3xe0Fddw
KLYc1o/vXy54Nhrfj4Ik/wD9Ry05Fx1QgsOEHkpTlrjjpB2UPGBAF4o4UoIzCdUDKUeTyFhbu2QM
DZfyn3hQLConxqxz09uV7o5hFkxioagDuG7h1VdCQwsdkPMer1ZYsjR+vDzc2I74WS1c71ay9Mbe
WiVNPO6ae5GxhSmUyy4Ig29Cw3H5+ydGCRIqyD4+zOhKd7/HtRm5kvnFYGNdUemxrz5csjehiv4h
l0sCZJ8HoV/B/olEF1jIgvzfdTB3uZsrs90QLUaAUlaZn7/xH38yt1+zv87o6jUlaBwpHNd+HkmC
HS6MmGYWY1j4rR7qXv+wvG6ONEwm3S1pvdOa3pXJBkTK6gwjtPMUMAK8BK61IAXVMCOLyaZAC/NH
t9DQk2q5zqPAN36DC1gEKnx8sjN09SZ/a8RQ6B9QQOTxp99bdvcIbikt76U9QcWsgeEVVj2ig94V
eKf5NNtwTIAa+GCGcUk315XvYOzeyPyROqMxK9DQlFlQYZW8hGcKlfNjaHNsoNWy7cT3KEjHQEhW
mw5K9Bu9MbUBYAb5mc/WAPqnxHXbzrQ9sDL4zLDoJfki7UIFTKzJJQkEemohnzvHAOO8YmxHKUtb
9r0XMIObT0hB2wTGz7DPzNKkkBHhEnnNx81eGdnMmPaEhfGPYB3uFJVuyhdp56GwCJUSTSOUhRgX
tKeA51HgsboKu795HlHnAIJmMmJ4c6Dx82pBf+Yf+xMoE7IrFzL7qu712kkZVhgsB5D8J1XXHnUD
2Jva6mAzc8Zi+UAPbvLxG6PrZZSNnd1hvETy/uwLaKb0E2lB1X0AcgYn/6NMHdZxwj3eAMB7AXMv
Bi4YBK8bHjnHEbaja1TF7ZYFDqqi3GhwQgx5payPetF5spPYLYIlIwVqqhIkiMaj8z8r1vMCvNj/
5mBzRoE01gvc90nt3tlTzlt3Ilw+icYLDi70UI7hdH3RJECpsvxLtd2ovlxsR6KqsGPFCxAZ07DT
Mqjl/Ny/Fi1RbMJMkojOODCTjJ46xmhoU7KNb/TnG8jUXBNfinOsUZk6aH38/qcVXdDo+XmcM/T+
Qrn+x7HZEys7NCbZlcLchhE5DrZt+R6sezPHcuT4vILHDCPbi3T4TKF9RxfSc9YDoDRggigkJRjH
fbjFqFC3nsxR68J49aS4wTd+cyxRgRGbEg7nriqfAcQLWUFA4VTKUVGkU2JiKGvUYymn8IHAF3xo
UMOsVhtlb1hpGmzNd1jn0tVEcQGkvpgYqzRhSZZIlCLfE1/Z5J2o/Sn/wvUfUzB0ulr7TCk7t1aw
b5tAxq2FUZsN9KoUZ9YejbqyR9WL4HqxsrOVIieR85sLBx28UDCuB5XGRlHQ935vCQTfMW/Ye4YD
UyLRvaiDVRba4Ztvzp1eYPOxG4i5Tsm7n4t+tq/410sqG18jQqgCadZJ8Wm7APr3VQUxIaQfbhfv
QbFMUCU3rUfvF1hhxTmhfpqF4sVVa1/dLufRKpddX+ege+CUC4pj/iLt88+fkhuAmQeMVrUu6IeC
9F8ojEUOIQLeu8H/hw68tT3JWgT9scSMPpy+GzrHHXHs0FF85q72RcdIyv8uFy31yJLfYAjf75+s
L0z3k5fxM3kYXMprGX70uX0cHJTX/TVgG9rs2rtriMyT0Uaws6qvMc7w71ufwPWwECAlsDe7/6IJ
ztVb2TWDmtiQbjRzfZZHCzZISAaPetJXXoMubQH80nw6zhtgvbvc4ZlkFTSC19JmDIcXaG8a8vBp
9NfM5RgAqqEMX/oFA6QTWlsFbYk+bJTqwnmuXgFnuvxzPuU+o3G8CSNocZCTRciUHbdnYC0haxAY
prbpiiy8HgmxP5b8sGTpVe/+g6DbApojjGIA8ditECLWK5k1bQNYIZuLyMsYpnA2nA9N5FPwbVv7
Q6LgjWHC9/ZvGPa+FGswKwRmx5I7A+zkbKXQYnhwfHpYzpgBcnMuz8jDOF5b32FloFCCZ5sYiKh4
OmgY9lODprQoj4OpAjydt1KXvmwaBiFczGK8OT04Td5TWj5yi5O8IK0ZEQ9k5ARsDNFsBJn3vZTy
Qltcxb3vCMSkvTX9LiDq6ONCdlTkcY4usYKCjLjPXLqyuLgxDC2vZrYEmI2suWQrA++8KaZGPABj
6wjBxbdxX90Ffedeid6OCuC1QubYrhfXUTaebYNgOBUJ5NEnQbiU6bQbWkGmCynMsvHFNupk9sNk
3h/PHIeNcNUZ2oV62VfUrPb8ddLf/gEU4zyJqILt+9gZuBIx5oDpkjm4yA1OT/lvITFgG++Y2NCi
BPUKiM9IsHEv/vFJMcrsKZu4qKSCTbj5TlRR3JKFb6foXTwvfOQnvSc0RoTOCrpq3pphPrZ1eUBF
egAP7CAjLilL3MmJTaC9GXw/i8TqIAsQeYeQ7VY3V4tHOcgRzaLL1rY9+UoKol/g/seNwl5aI/oL
/2bG172cNbu41oLCSLmA5N0CdxoXuyyOxL4MdAOpZPvIWLmL7UdwWqUK6uj2o0z1PFpf2sX9Ai+H
VSPL+xrOkWo44WbToBSqQYVd9ub47VhaJC6M1TeA/I5cEj9zUvhQkrh6oDhU59F+Ma0ETvw5EXRZ
KbkL045D9pxY8tOmODtVxaKFnPe9dl0OvWcYqxmxlxZtJdN/fiFQt231OkHnK/nogRU9d179EbTn
JkSOMGUISKjZbQ/t9MeMPKV5P+nNL4yqMTSloUMf7hx6DzP0TzSS2OcsnP/Ui2DvCoKVy5O4+xMP
f7CkRRWugqkH0A++PgF8C3/eo3u/u+xYeRs6nBlCnNGpRAQMAlXmsrNA6Esm6ixIR2Vp/z4Sen2U
CsfjoLk8azQFoaXbeE6SxDIGi9ELLysjQ8UxHEMQDqxRgv7eh1mmcWvyUOGVy3Ks9iNAStic+fgT
8vEipp7Ugp0e0xxKqI+14ZjsbIYgfPPzTy5nY6tPFRF39DNAnUVAjiErRzwXbQy77zXPuMIKXAgX
vMBc+khF+cnzGaQckxbG57UE1y6hSNsX7aTmhldfGLu0kvSOYXZYqYfDkIE4WdnAebzNQ/VzP4+j
d3oNIEBP3eHlnwm0u0jLj3Az7K2iQ+PPYAp2XDLMsn9mvw0jQT4q3HYr5HKLtILlsX8HScIVqax3
ZZdqZ1KKPa+vybs3As5amlNjuSyyHIa4biZdbDhS2DWxtrxV+t4iIMG9xonJUO6EIOLR1nuYTrZr
NeCjr3mYs2D+KAZiD+I/aRGWqs1i1V/3/95P9Yg9fze3/ptq0FYNKSS2L8A6P0lMwhfSYk/rXpds
DA30e5wO6fFEYsTdHhXYTwFBE5MUZGjMkiKMnrhmKc2avXqjtMhAomdw1WojVbP/58ZQJ0m61Kl5
cr70HMUNEtHbQuUTvkxK8pEY5oZxrdf66NdsiFccvU78cPytvD3Gd5mC9zItuNexHErhFHzDJgpg
27hpk1fziEjEKV+c14s+bld/9fGxisIzQEVoYblI3n1NgbMqMBfTHydq3+9J35NWeFSAyu/Rln+c
oFwB6XAPLkEut+gks3KY2z8jVcGYiK2YxFq+UIAHE5PUFSDc7C7tabmcDsd/znJ7wE2euXBT3lnL
DJ/+whHr78L+JCVmJ0W8YWZfFGT7MNFhfCBUF7yRLhgB8vMJxwoEYlEIBmKFipLE8wPfRJHHXDTe
EP+KtmKfV1zwFkKcsPTV5pPbngsvXjIAyJePvndiR0ErQj28cerQPj3HTukE2g9S6BHNISZeR+5Z
yHjkqWBIG5n4LBj3vLibW7cadJ4c1/XvWdLR57XTDp8+QQwe0zNaGzrtgGMbCRbG82tNw5PqpLFL
KCeHBCohi3F6fW25xo4U1mjEcXZMEY4YkwGweslDFLI8ZLAx8VyDFROOXZnTcoTd+jWrLS3tqwnJ
402ub+i8fzfzuDP+jYhlm0stWSohEenCSY3AngtERgEBOYwG3O2+oA5NIw2YJQA0Qj+GIHA6NCjP
Cbn3bauBs7WjY7RqWJl3ZqohqHB8n63NOgE26xEwvobdQ5w996Hc4PxUN9Bqj4HjudSk27sB5k6O
7ann+iz26AKqFumw6E7cgaUtmtf3Wga7vEHrS9Ec4f0Oq22iKbbMshlHUu1eUYY1YQczinsIW+Ht
L9NS8qfLU2Y0fFregQNw8JrmRWiF2g9Jn5o/uFqQN+Ovmv1UDykrsknBPZEggZ7F0nsQzT6wYFlf
+a8evJx6kkXihi+qMBf0xoRz3TT+o0XBUNPafblPYBAA6HRFgR28+1iJ631iztgzDM6/9MVluIWM
lymyTNOIuka1rzDRIdE70c/Bzdv8wKy40tPeIa7GiD0g2zt3/Lax7ZI7KvHYclee06NwW0LVr4OU
y1e5q+PkpmSH9L4Xj43scQdWHNnEt4Tc2RPss1hOXKIWb/XbnI5jDNGU5CfFg0dqlj8GnEsaOyn2
5D+X1cAsIKsCc94xtTSBlWqctMql4GMHdZ5rW2nS1apv+CWX0/44odMesK6t/v0IQMealjtOPeO3
HfeHHXkFSq7bxysTllb6GeDi6HOm3ROo4SWGb40JSK4DEzd5OpDjOYmgxSZuDUoZ7dzLDR3Nzn/y
xYLeT8+9cm7ZesNDpA12RYiSnecX0XVyMUhugo8KkmIJKJVNfdL9Mp8E8MhSiUbg1Q2m8XauqKg/
+hPvgc1VPCkeexWQP7kjxmVYLZbKYLSpneAgFRKGAPigQL7YVT1aGLAQqCJwwzjFDetnpCQj18+4
VtAr152wciHJuUAWwKyO8kQHNKQKlC8a6hAecUa/9F7RbMnGd1JS10cScl4hfMqfmrQwElhgMbrk
LvXFfVKp8zUN82z/F8d/s/WEYtB7SI39kh+je3isq1khqNdDn6q7Kgm7zL9I3TQDGUKEHdODsRsp
phtoc2AWZXgjyLu1eDRV+n67M60GzyNp7W9tNFr1AwOyaWDVeDlz6k0GrQAhs/OEDh6A9LQe7mTe
AiPF8JqNwq0T49jo8FQ7VadkII4qpErbFbWUGWoQfy9XNj+DMXEhNNpC0QMDz7BCWXQP/NgVtfQW
TdQsgU6iu4450WvqgmXKhw55Ik05cA4Fe3CVmvtDIfgyKiPra2ZoAO10WJQUxPqD/COcsnc23V7B
8xwKbOlZq3vEUkjwcJxAMTyMcvpCfqA0B9GBMFksYQwPGaoeTEXb5+6N54RqTi2K1IWRU3NrFpiw
Vy7tGPkhHMTZ+9Uizpm1wGRSz3QFH04F9Vhng9frOc5Bh7Q+QoMlIfcNquwkzKSaYYaBrr4E8pET
oeBkFu/QGZ8KEQf+FaNxNcvU5N4h0xtqiqz4pCygMhzftOEGLLHSEWqipUnfa/LJC+XFkIMnvQET
iveo1RFW24T3YyBYwaC1MqY/rLsS9JRdzheCAXuvLLRrbmyNF8gdB5eMNAOLZns2dBCYwYwFcekM
g5GqjKqBYVRgjrLOrwB4fl3ZwxQBmbaHkfZ8TGZKM8YT7pnvqB8692X7/DvJRljfr4YTQ7Gpe5mm
D8m2elskE9zc2uqA/xCwPB7Fol//yq6R4k+2g+TGL0IlIaUrTR29VQ4igs/fNEXvMGtmg7bnhxWf
wgSz7qmd/SHhLLP28yD4+0vp2kPF/MkN/WsjiITqAhtLV34mttIS2Ykz6QPA15DC5sOG2pGkWf5a
OKEhpUztP3wieYLhMAKN/xek4WbKVq1hipQNZjBCW6miwA1/X2X8hQ9lyGHBF3/Z5beaO9SPajc7
S07GjrtbFkxNN61WjzA1gRjI3T3kA1zM5frRmdGUbChqf00J9Z6P6FN9JzMSu5/OK/Duo+9CEkSp
4r9mb7FiwbYJE6H/8xTCDUQpw3G/Ps/XQwu5uqupsr9KYHvDXFWeoF8qErZg8mjOAL3icUeHWzSS
Hb8NZw8ZNmgCbHOu3TtSLcXIO4lWqut2grTJOCLvT75SPPf+SXNo/bwswyNA1Vf5/juE89Z5kkeQ
dPqfH+mWiDMgPzcUBtgI+VYMoOJ6orUKAb7BWBzofwtsNifIytRGPQHuIMCkgQoJ6H6BijSW/J+k
Az9NTzvkzTUr8YcN5wxI5o9v1kzVAgPbNW8aSFm4B5S9gpejHinAKlF5Y+exsp8OEzOuXFaHZTEF
6OgR5vQUgtsnUdoSVGHWLZ9ufM30hE/s/WlVF+7PyHlZKDms+qdx9Ilk6RZzAzsAWy72bUy/x2NU
9uJvgRRyQjZrpRW4vbFk+GfCr3yYze7bhbKJrwSlM5qfkFg2ECCAT6J8etQqVwd0mtuu4djJnxXz
1hPFhJ53IJtD/Ya2HrmiQNyydVbNOAj+tRTWtZH/Rx1BSxn5Zw/0hhZfx3O1RKbQAFXWHHgT/bpV
1PisGIR+cBVeng7bdiSIicmoab7LbhOI+cbPLjFmBhn0WrITqN/VZKywzFb9mEVOVAf0ff95YmnF
7z5kWgW9BK669XvxzxY6MLkmtk8psG2QviS634ifwU1glbCja46XZWQMlrwlavLU58H0GL569k6n
jC6nOJC6slTulmZBZWXDHthN4URUg1OXFebFKbSZzFl0C9KpFh593QJfTxu5mVQ3ugkT2A45Kmat
b2CsSQQSmqqDGkl0wfe4kRMiBlaz5M6T42IgN3aACDX+WZzkDRP0RVvGvxKwflQ3LLhpgVkjdapx
O8d8LCQTDd8b4o1ldB97R9PXcwsTKKbp+i4l876YWUxzhiyo56EavYZ2DMHjNN8gslUjUcSyrQXt
84WbLCzvMIOsUnSu66dCEjr/2U0WygZqUEYM3xmX+OdkAxMyHnPT3NFXs7J+fYlnXaMyAj82xLg6
Z3lphSCoqDAtkswVyyGngqKLQcQMCIde8knsEhZGT7FPHtCCKUaJ5BnP7Mpl1TsctIXrIRQ5wFxA
1c8oMFGxv/Rut9qz5HKHw45Af6OjI/691zHFUu7okOqep0Tq+f7S4ycKaQ/YbCstCU0qUU7Jjck8
Qtj+Za2uhlz45Hn7oHzPVHYxRaPh17JY6x82sfFtiS5QfcezgJJRXXBxzJPGGLGhtd7VUE3gjlGp
KvPVP9U7e0AkWAT1q7GtsxrZ2QQGrLjFTK1OrdkJFNZjdP0uP2Tb0M+rpSUrC/IPBZ6qCmKi2Um6
flDz/y59nIn4ZFegBJdqCJ47uzfs8Qma8IsSz0/8FyqKffL/KJASh6X8Su5JtTsc/iGfD1OWIXfX
6W0zZC94YADlyD3zfdxsvfgK1O8jfFE40URXIAuk+opONtadllf6OrE6weNo9IWVCJYlgxgn5DEN
EP0AY+sOnLqWH5P3ePVcLXIUwGHlRNJvXXOdEsmiZAyJvWGJ1LaeFNjx5mXI2fw+PJSRRxoX9MDg
/s2JqG0auPy4nYXR+QuMX8SiUg0UMFy977Ja3vUZuzFHUT1Lo0+I9cnEsZvvxTYlMslJ2rwJ4Jg4
48xTxujiJ45+laomCHkWK31HyhMm4/1nmGTedGqZ42eTXSpxuKldQBzBKB1vXJoUWevutIkwMPw3
+1iFW+cmL14z/36IUDRoMh9z3soceRS8TCBlPyn2DER7oey2qegsRkopvmRY/6mhkl7SeQL+l3r2
6YWPhzfGqcdBmH6RQnrZ50INqzMtDNj8CEx2n/p0qorbvoI71J8qZg2tZ57J18X2NbMjac0HjMpN
N8j68otS3fzRFyZ85rf9QQEXmAqwRgtDujiRR2Dk39mdOYXBngkm9e8P8WJSRbEd7cM3d17oY5Wz
MPj+lOIzlj4OJzpLiMJJJso8Lu92OKQvjzlSYPvbC2NPkBn2LPdiG14cBmegx1FyMAWyVb9pa4wd
UTL8lJ1mT722TAbCP2wJrp4tA9I2Px3kyxkSjf0irAI9nYgeSgdqlmDO69huQlcDlmA0F6edpCma
9jdp++chXkb/vv4oeXmAx9TfmIDc1+rYtOvX1UBZsZ9fiLKKh9BggWDecMS/iCa0D320gW3NAXne
xDbJRdqfYVoKZFfYVsRf7bYEHi7tEGeV+cbJ35sOOG2jLLuu/38FVcfrOFAlPO5DQkcU8I0MbVtY
tl7UTCYx7ssauoB2pn+Uo7dwK0lledtE3hJDbdOgY/rJR+Jm4LNUrrWRAwl845PfcBdrSA5U1hFA
QPuEpF8XcCRbhQiJtEdgmqgfxlshtPYkARiCiP5c7rxgtcKONusDOfJNHhKU7WGlqJrH0/ATsHhX
DliYDoH8prMctzeOs7ffcReGkSoJ3laPGCFQi4VXlQOIiC9m/fLDlmSB/tDBfEfanRby6979+rkx
/GGB7TB4YymoGdjMTQHZYgeI5cTN2j7OJFR6agEwaHRD9cZT3keLz1ksrlIo4ZGhXZxj6PhlB70E
t4ZJYZiyE1xVNypIIrPXd30GGlh8gzmUWXB3Tq2j3xO4Buwx5h83nI7Bnu+nSMn4jtthGZmSig4W
LgQQrbQBnZmALNgKPUGA0pWmjFlui1qXUvm75Ibt/GnLYBzzAJO2mFReF2ihMeEmLJ/cNkgpWRoB
VL3egO/Oq8T7vUdso78heO1/jIOm6mSOOioVfSh4bKFXo9XLIXxTIhDNeSH99d5y/2V9PXOOrGRz
T5JPzVXlmNoqNS/P/fF1D3fW3TS8z8lPipmMrTwpWL8oB5wZsuEDvig66hGF2A0AiYS50IQ7BD/N
tMzyCsEDIevLAn3yEQQ5kBb4EgIk3KGAxWXDyKOB2VFGdUnGPioe2HN5FVIZK7dO0NzsGFR/TfcQ
pw6uRMxzKWSCjV/aXLXlX9DEAhroiJYaStdjPDlV40IsTlntllHKRsg/0Q0swkHLlH99hMvjmfUA
9VzBk0wJb4FDuwJWbALsr9owK00Fanm79rL9jlt3PnpYq74EOgClAdF96p6tGhEYlck80zuRNZgJ
jj1sQZPFlCp8X0aGs3G6oyIfv0LOuBZVrCg0ckUNjcDi2aXaZXkFsW6V0QaCPZ6Hsd0ILqLDH1Ou
nW9TBs1zeaxf410UovfY91P9RceCXVNzFc/uGQJUGXzwHbXcJIhS+kslDqsktpMbWSunbmq934vv
gd37uyg7e9Yl0XnYx2JnRjMvvLTdMgNT6YTSM4breE0tmFiZPNI8e4nofbBeWa3vwegD5HY+rpZO
cn/hXtr968u4yIg0Ozhh9BSVe0HRdvXBR7x/wMoJM/HpKqhXfoLKsM+7QaEWanpuK73LMMRjJoG6
FNNaSQLNfqyzd7uUZVRCwv9SfIko0yid8SIwuemd/yOCfUXuwtc/5bL6e6bfd6qd8w7nAm8uPO8y
6saolOh30znogiKv6PzRF+iL2OPYafpSfi/SvcLMgWgmSQxv9pQTeogeeWI8B2LY/42qMVPOnWCw
q8jk+/6ovcYp1qAeD3wXGICQkK8yOMX/+xGrBK5ZYnevACd90cl8AeMv+/cDuVrz4cq3+D83LvFt
3vzAHfVfx5KzqkeyPN7G+gpcnGJr6ioC+7M5h/zWwYycVXdeVKxAYT2RjP4FuB/N44LnR458mo1X
lmzWfP5yjVHWe3msKRPAXS5uh+hz87VGBdn7j6jCUBVzpFXRLvOhhsnhtL+7mV2cK1dfnlnk5LM9
7SBLuB+cd5/plH6ym/YEZtFOwt4Qubl6qdau1MDne3uw4L6vWtLXmH5iPCwrvUhzcMVdDBu8GQIo
dBUvHmrUxtjUD+2ehZVDmzoPZAjKkl0p65lqN+4g5GByrvJsEwECbbkz3MIhB6yRd7ON7oQXH5i0
jXwedbCBUn+42klpwdLwjskRtedX+rLxt/6gHHZ0ntE3MmowD70WmT3vRcsmOlP4IksipeTbxsxz
YbafYHKeQOYHSNXzYWUGG/l839fSlUvOHNo0x1lAn0nJ8Dg3gWP+/8qJZCwDgGILg4QtTUj7AUKu
O1WIWrYzszuK7VY8TfsbDnI4SOL5SqUtTnRPr3U6yGXhdxtr8IWViaK+xCacHsHQ3y7ht4N+HnMX
2VBnOLKyCmGoPDA4s3WPayfoIFyE4D/pCewGnGb93WYDJ1CakxvkRzTP13S8hM6Fy0BCxw4IUhyX
VrXBam0ITkNH/X2GgN4asNHKc7VXo538RwNv5C//TsXzI2tokNvDWAWrRaOpJ6lpHbRytvSLzeLo
TrQmlJHvQKwTrUkU8psOUJq7Pw1rvZivMnRWVO8nQJx3FgwPErtbAhb2wKyrcjmjWLdd6/b+6Iim
9bylJU9c99mgWFJUhDvwkgm8MLTwbIKg5VlqRFRihEDomHxvf4Rw4MY1pSk5wzf31HJQQgXqRRS4
wu7pZ1fzwp7giOJ95K2QpvfzIBVYKskUtd5tqmyrXKFTtNzwcGIPknHToCdLzR2rLqfzHiE6EJDp
l245Zg6VdKstP6TvEK5jFZ7iuxUAY7QBgWJcZYOHLoJRVrw6EQabgOOUHExBspjx2Owi0kUMQ657
hGV7uF55VzRkzVpweeRwXizo+P1wdlS35AsMd+j3+58l2U8nxuTk1Jy+5gC0A7Y7LS+k1K9xGIro
Q8GRb3Zr16eKwkloJ1J3dkuDiqwWh2HwL+jJloUUiJbzVRcn2W6yi0H0jE305nu571v8z1UJU8si
b9gDLnQrS9vLZypWYO/FYDubFJl0t1SLoAtPBiAesfcsuZh5qxa+3jtXZK0s9D1YL6qgRR7ia90c
ICaUKktFYbM51Ub87grWz6AglnegHFQOsonvgVz+AzXC7mNBUSDhW0L6Ccp7+zjRkFM3JLyOFuME
e+Tiwi64xcigEWoeP93LHNq2aXdz0wyTK5/c5euecSbHapuLWjSr+QAI2hWAxK75IYPSlk+jyfyW
iL72N1a7hc9B0AjFW+j1H2MiLWaUCLEZATDkz5ga+QYivjV+O7ck9s5vxrPqiaBOTZke/KpmkuEc
QiPV4E0LYu9zLls/G094q7hLoxiff0TkL8wWQIFHsDupQRlq6MFLth7vwXC9k4fikRbkvNPnWpYC
GtxzahKvbbSYhvx0Eq4EW0D8L9/apxJwfdYwX7Fs3LELmfvndww8rNLvMWwhrDHeGtD8kBcll5ks
jMPGZbTigrdRN+wj9631zb2dyRSxCtk/st64CMxucFI9ljXe1VjkPEHk6rBXIgxltfLZTGGXAT8b
/1Nkqw7uWNa3wcNzsdQSrFo2KCTh6D3++2dXonxQM+bJj3t7z1qF/FWgp0t7f1X9CfpiOOou1+/T
MfLB98bfeKQpBEG7SyGYg51dUjJoOFV25e9apb5kX/y2vHQnwjZfP24YHzhG/m0uCCtvgB1hZgP2
1+zctRhEIlxJqz1MxYeJpB5XU8RjgMAzCm4xcHyfpvVRxnj1QJHYBBgFlAxah4Vn+drhwR2ASeIj
HOQyn+du7L8SyU0VvVd1tgULX1Z7qBGou3bbuDyXXeYMz/n9SnqOp8tFvD1C/IC3rFXQUpWHGGH7
dhE7IZQfwS5N+h2Twbf2P3//kpAs2cwzkjmYQVP6f5J1OCowtcHm0XI/eEuEs2R6SGq0Lzta1IO4
JilaAEfaf4kJfipnVuGaK3WkbTzZW2b05ummHJCof3lxExOGP2LThheVl36J0hBADQ74VfpZuJdY
uJWrYmnddpmScRS8PnIcC37Sfj/A6u2i7Km/waSO9L5yNoGY/Of93d4U48bdPUoDROeftbozmC9f
UPNooOQ0i2jHv1/jZulmI9vTKeMxCyn6AWtEJKU/U+FxbYqyG+M2C/j3PjZkPLh1YI0RAAySEutp
NIZhvGSK73qBh+5UnK5MQfDydXpJRlS7wwiI6q+xAVNqVcz4zcJL6k9TZ0QjNl82QVADK8qcTOQ7
HpGiE9+KTo4xIYX7V85+7Okp7mdHGfFw5fD6ndS3c/IA/eeVhv4bL4yAxJV1D9n9JnEUCFuhLsI1
1AMkm8uAKbOCKnW31peXybcvrrWlDdNR7WILycYmCyiTs7/hJ7x5PQMwNd0nTXOr2DWzqTpRa9qV
d1N3eDjk2BsKQYNKSH8cWvMKaOBtGLHzU29OCimnaCY+qRkhLlugsw/lm9Qd1Z7XPYoMNs4txkoX
FT7+eagd/A9t8nFJ/GXONOsEbt4sfh+uVuvRlyyydKy2HGXIPEwFuugtBqSWKtyVIPJ9iYKqwR8b
gSBPwRNpcD6jp1oUO5rRIfBFImVguxzFfBBou6y0sfx/6nCdOdfZpAm0A8p0Tfuub7F8FVWyLRpa
Bk16+qfgFFpeLcNhyxwX3tZDX+uKIMZO3MItBjEwB+hERqOcNOx+y5idemX8H5zmpxMloWTkCjyx
Mlts744VtTr+z5Ml0Xc4JXfQTzZEb+cYl+NLqGVFg3ie3AsqRTIhgQNPtfZVbq19FVwrEgHXbpnV
0/2UQQu0VdWdj07apukmFoRKHWZ+SYk9EctzISZ0GTpP4FEgg5tbQXx9zVLhXvH5AEs00D8jOI7J
FcvJep/d9Q+SeTZvsNCbXX8sk0HOinznzaBnvsKQkrapfy8OHegbt1SeZa+lWyb+0MnGOLhHMzzR
nhU9pgEbwgqCN8ABiz4Ltn+am8T0/rZ8Y8Qo+J7XnzSfks+RjA+hrB8QvEh40iCRzvvw8s5u49Re
FNKgz5Q/Bct+YW9hyk7eFsadgTRfzVCu4HIZwYXwKHL4j2XtBOl5tqnJLnoWCXXYE+I6rCd3TDKH
RAmJIwkhZZauWjbfHkEqakohCPWET5pC0nnU9Ae1h2rYHUAmL1cQUFgQcA422KiAxO2ffYiudg2o
qZ+0m2mSQGPbU6bvOZcmtIrpusRvnNCb8i0ZfbqoLAZ/uNqMidBvWVSgrUanqGiU8l934eYWw6br
lkD/tM0CIqNoCWtCizVRRBlAtMC5ikitbXhV8SPVa5FrlngkPlhIBzTrr/crcpEu63a8Zx4gmNdO
o1kIqIDqgNowiNWuExnXNaeqbp6K00vbdS07/d4CRSZE4qDImyd0qhVcqsfMIMzkcBS+WzKwx6ON
/6ofluGgFW64NJXZVHDFFE4Ef/yXF9T4z+eKqTtbzqGfH9LI2baNKtni4+GkmpHSOvK2cvr6pt79
1YTb//JK4aR0WczeG2Td+fgJ4d1RcOjio3NP+5gMrc+oGxqDFGDYmKwbaIfDVFuqUE9wdcfIwwy7
ndq2WOU6XemcrW6mEhlbAHmD34/QfT09y1heLuB36WoDcl7Nfw8W4gdc7uvUe7v6dMUXNqDy5nXq
MQwAHhdlTeLbO/5pIn5KJoey2/QkdlKM2P2MUNOn5s2hYP5RrdOoWfg4znvd2183gjvSZvj7uyUy
23rZFMp9PBhPABVPJlTnmCeM4krW58o2v1WwcrODrq2uecADt2yNjXUcQyfY5qsz/Mx+7NzfHRld
jTzaRCBk9HYShdwXzr4BUShzJZVq+dstLK4MEdTGfYBrYfK4kx78EGCJ5nZy+NeVFG1oPIYTwBt7
yOyzI0r/rXd52ffUNf9ut9pkf4K6+RWakGMcjslrUouLQFFK7LzXV72C+7CzxSbaKGBYjQuU5u1f
J6mIsyR6fyEqPK8pHMr86/VUdGta1TxQX9OrFS/mLJNsudHU80zWlJ7lQx8rCw13Sk4DBuTgJxGm
p14/GRGizpP0ETypDpqGuJjOTFkR+tae4hqqMLBiExtcKfgDZV/U+uznLCsoRdFT6oeFkbZ9alJL
ct3oe1SqTaxSy9CF12yBx/1Gj05WXWRjheo66PyfR5Qh/G5hnlD1qrGlT9Tkv6R3+jgpWEJM2zU2
KTf3eT1qmJ3UPVeYzvFKimr2JHJkrvn4HNZQhjucGKwIPXmgLZHw3CxH209w6IVgQfn0PlS1hyqN
FTUXROywVcmKo9kXTyE/hszaSUpcoTVp5OIPcPdK0NzU80g3qT/ENo7uqSsse/D1ws0yCs6LHzDA
2UaQRYq6vuQ9cmixF4Pi5FGT240WLl0EHH99QmXZr9fyt0jtwUPuqG0LuOu1UQ9aZO6yzkAKkynd
E7rO/DxCPS60n1xM5PFUw/115SrR5eRR7DlmCX/2ELrzTXHvF9teQKpzLdCMRDhmjzU5jTBg3z+D
6XIZgPat8e5afkY8CLee8kyA/wGH97KoDtZXyx3pO66yz4iarcTIpLmLQ2f3DbOPTVTY01eRaqJD
Vlr5N76GF1b2yxwJMIJ0iIA97QTKzJrOwPcVYpXOLcQDqlnuTuD8G6J64RbknRxPub+oLwnY6VpW
cTqr1Q2zVwdtacs9a1V/V0SQFK9nlQ7vKuQcv240XWF7zQpbpcdwIzluhOZEEQzOk3lJUWU0WC7d
hPnh0B4IFFrgYEKYW2a+e/iHd+vEyh/bzfkO9QbCSuf/BdnLY3DI1cDNkRXpVQBRACArJNQ4haQo
xmtjIUe1uirPhsucTDhCFqlLNaxeez5xVb5uFUCCrWgc5kg2psU7Y3jMG7sxjTvLzJBE+KoB89aS
+270jJWlgboh5khtj3m9iS5CwlI6jKxiUWrYva8g/7V423VJEhb27GnJ2w35f5ZvJ1+EAukOe348
nKqixR4NfIGc/LeO7G3rOcDxFru0u3bxofc/+nTLMK2PWvmwtIlfPXdpNpmEFQX355qWEEG+KXxf
4L6h6OBq+jD0rJgobsnnkF346oH5acChIW6xl8Nu38+fYMgR3P4Wuk62gFHBYLu9tV3MNYGCoH5J
9tusd0QXRQxteGbzVNCAJ2MMI4Egr5NrpZDaD2+HhQhhtbTygwHvPJ3bMv14rVWkZIQaKHS88Cvd
9L9ybPLuY0jrpNo/FI7kg6BB5z3F8atMmsHmeNGTgvnWudRnW0wTJTDSs8bWNp2/Wn7SE+e+nHNl
i6bKX4XZZX5kB1RnijOqM/ARoJ0XpJWiLC5Mesq/4ABBwl3pDb6yWd5gJBj0ICT+8Nntr6wei2xX
efvS9uehSpXFl16w3LH/Iyol6WcB37UptGvt0OOY5yuaHnrPKQN1AgPZUDqUoyH8K4fx9Nt8tbgX
IED8TLW4pq14JVj+/a1MTY517Qn36AmQzGo6ruA0U1wdWoCC6vkPxQaNOLJAfIra3TDfv9O1d3p/
yBG6SLvdABl6ZLAl1rsP0zbXVUZk9FnofE3Geiwi2I9kIFfUb58O8jXjJrwWOlmKjkwL1I9D1V9n
7GggiPQ9xbgzsNpkCKEkxOjLh80PmNJlans5FUeNK9C8tD3vwO2yfgFp4QGM9uvHAAL7y28u9zGs
EgCA9xVKC2hO37GNLgJOEHGtQtM8C3LDjL+sr8w8thTnLAdr+Txp7JPTvGjET9PzhA30c18KtEa9
QMm2siEiTVGgw/uaujuJ4KAEfu/Bj+5iqdOZU5YfeGWttXrs5Cxv7DGx93LX6GB2mRuSzOlATNmq
RcgdFikw6Kuz/Mjg8E1c/NEHbpAGstePyBqO7IG8KK2WC0QWtzog/ySSxNmYr2VTtwjkQzTKNEvQ
Emya7dJI6AB9Qkw6Yp/+B03hwEFK7MvOdA/MxwTKtezN7zlshD4ug+Ri/AF51wKlq2BEwQjnyiuO
/x5CiFrNBEzFKF0+iCM8Se9WIR5zscYGufmiMAQQ21jJoXew1h6JNt45V4gcuoA2u67nUHch0c+H
Y4rKJ6/IkmcLsvKgMuHODPjJ6Wp2AH79eimHtoBuyHVNb/4UpRjC0tcyxPAo3Q5XB8X4qfLOoZTJ
akmD7c6f0j9vqPgCZM4I4KkOKhvryChOq5dz5AbVHA61OIqnPix5tbuqs5Gwh4iXdIXV8mybQq18
NjcIWSGaKhQgIsPEosxyX/qrsFyh7o/odbf+c7LLYiGbe30dgjuVh8xOyZGJ6IsixyCYNeSO/LPN
onGD8G3jFQDFvlRCf4pQBEBY152QLc2+r6Ns6xPxjf3xWQAwe2UFa3SuiDBxEMtpnQGiS2TkqTUE
nWs660ICNLVGraOfiglji37PiybKEDXDfn4ncNSl8LPtpifngKmTTurVBRCRr/O9+bDEovcJPT9d
ukbagO8rse3BSmNEjhGYGNcdxKXBh6IhAyN/ISKVUjfP8nlpv452QnxIKpeXnnNMO21dIyTH3tx3
vukdrOTwu2qgsTd04IQD9mPI9zwtEdcCSiMCqwJ6EtUzFrFRiFCwiOJYIWqHwHS7lXu4sywaOcQm
g21pThF2gvbVl5nSEeF1X7iWfajrvH8I+dlPoJ6lvn3/UJWEY9L9N7sCF76D1+Y/yuuGHhNqdKAc
d5wYMKaCR4u93Lq8j1IEC7wpyifkN+BfVDxAid6km/Wj4n4xTL6CW1K2r8JYyYO0HlqnpPMVxS+y
5xBINhtYxtSkY3FspesAlNgAVsucU36GVJbxIMhGxXbRTXU/wY5WUi3Y6iQQtRqjm2xes8SR8fpD
Myli4Qq5gXmy64Iv3UMOKP+W09d2woFAPl2Q4iAaNccsayvB3YdCmmyZLbV9hq8kaIlqWQQAonjn
wsPfY+WiEp/fVk7AWjTzox8r/vR0MOLiSm+Wwj0KnpvIq5P0fbueS5EDCioZz6B7UiZV5TTUeWEa
lggdnseprNq7eBtgKzfUNW9hn6SvgqztUtNKjIa7zH1jVYAGca+oZJwxhRqaMuSo4YjIgR4g6okA
p7ecVNvoOxOPSlAHhBVzOP700nSnw0tNv9XOH8B6O1QQLyPHSRkGA/kF1V+PO0+WnsRot72VD8Ja
6MTlHPp2PPzZ4wOOl8fulJ3AAvulJHgx1lh8hD0Zf5fhBaGmVqy94eKX5XvkzGgiX14TACIO0qlh
GHpq/wKQRkyphGgdWEuw8dOMjrLlw2XxhCA2egT/kEG/+q90tZ6sIB2O1IljyXzWIyGNfAF2KoS7
B8aNf9dNQvpQ95NN13pB+Y1CHS6MCXtlX+um6lCV69ACHX2lAPBGj/99zrdt8QQ2zGu1E9xM0skj
lhwDqOkxQMVQBsKKDZnUNU35F4XmAjcrknqJzBCj/n5bbdMiTzWYZ89EijvCesZKynWU8YdFlwb2
kLE/DYQp7VJMIPzCPaJr/9CfYkGkOOOv1yr4UBZSpi6/GoC1oErOOMPacCJ+2FyHV0oYgjBxV57L
nMSna4GKydxMFTZteVP0poQyu1UPDnQMyW4c8Dkm2ljFvxo6v8o31zc5u4ipgMvHJJ6ZUzc1LVXb
CgRf1cjgaL7ALqeOJf3eBR+LeEXI81XA4k14sGtccqhoi/ugW1aaKjbpT35bUFjLTlWhrmuDNn5s
+l9MPD/7jcJYxfBT7z5PGznzZtUa/KZyXbR7+XKRdTsYW/ww2l0JiAQNrfKxFI29NJBq8Lbrnv63
JA985+A7Y5Aec6tSlam5D7yiZ41OSTsYIev4OQ9KdWi08XKoQaT0UMUICe/83WynMbvtFpcBylxO
ufnjH73uORcDqbO0Y0eKUcySzGP+QH7nR0kpZa4x1AS2ihjDThUpUUrZFNy4+tI9zV3X8z96rzZG
NEjpDx3w2x8ff/1UBwYqYT6fIH9mu4sgQv7gK0NaEByvBQ4cARSpUUbKwmyCINFOoY7uHaA41nkK
4R55pCdvD8L8Js1aqMOs9kKzQYc1jckXEK6ircvKpbwSaHImxSlsAX6QdPCdfyTMYAVea0PMQqTk
c3OBp2d7/vxNuOvcGS1pMriqdwIdwT/fAB9hmfm4klrulNjpN0xznK+RBEI0PscNX21ztkkz/Wdr
y8omOryrqtdxyQ4qK4HB6oPypnYZl5YQX7J5PADEJeK8p7wVUEo03NXgXaT8Y5d6SHO1HPJfwDQt
/hq+u6mr57Svvf0N0DPQHVsEk8zhBqBpdlWoEK4jpfzzuoAOrxARUFlj665Azs2nilgcKoXI+S3A
CiqDqOsqlkjXwfa5l/dfq+L8k43GFRjJnEIFQVTxTJOa0HujCb39CRBOjR7PtbyjSgWkU70TQUIa
yGoxsn90wErd/WZfjbF3RjFJxpNR9BHCFDZzz0MOblIBHczP0WGy7HHVBTzFoBZDYISDjHFXo3+b
IN+GUGYjzTQMfZJ8vbhpt77YfNbUfKT4QkFE00DymnYdH8ItzqhQfxaup9fzD/VHmp6O9toQzDUf
G2D8dccHagLQjzPLT1Z6YJg6C3Io80kNFVB/HwvwuQYXiIHo2l6iQ0cfbrn4qk2xuRHHIOL1ZhiI
ccQjuThZLkjUfFQrFJqjT2JwqcBQnuk+V9M2Gu5yTYSQO/bqWVqUIU479mi2th1SPYJDIwwf0woC
YI69n1ZP0ogfHSujtdibvK9pbBB1uLJmAOz6dnR1v9kZlRWRZ64wghozoYO28gbUyfjNSrqDKEry
0wGFb1/YhJ419cmopHwbgNmieumK6Emp9xldGi1MCM75Cd3l+3SKvjwQzWa918gxjE5DlZf2dlXq
oEVCK3qSONno3x35iig82I1ryX1cMFJ9ERarCarwwfs3X7/lPZ2HZ9jLr252pApWx2pXzjyxnkLG
0jIO26lBmKXM5JTaPGIZGSq+YQvLE54yCOr3YmiAc5exFF4lBJXV91oHII9ZT27D6BJ7cLRTMfh1
UprLcHZ231xuUTmiwHPZcvHN8fqy0FZ9M7aHoCvV3WjIKHs+J4ApIXHzmDoUGsyX8qVkCfZ/8YST
b1LEsXGw2PQfT+5TLJXv0YT7mnQwidCHqBCk/QJCqyXOEhjdn0gnbWjWNp1dNEHFzCdJYS4qhA38
j+T4uNwKsL0vW4vQF/6Aau54HEF/l/Ix+H7OQVm22NjSW8qkuiT+SqaA7zYDgVmxxXzFingrIYkh
jkW31FJIpsxikY27HS7D0cXn93nu8dNrMIJGISUsk9VjpKIS6/EDAdhwJZXrcZxa84XrYzVjESks
VS9o4BgmrsnQ93qKN1UPMFyRffJnPTqVpsRCQXY42O5SPcJecTGlDsC2gngMuSNtFwQhZc2XC5Sd
5zG3wcdVlMhN79DCaJlpIeciYTvQjC3ktO9TRVQ0fD/yhzb88ATzf/6SBHCI49wfwqakcRiCrupQ
c9VMlnycOzh7tB2qp52jkODTpE2uxJb5ucXn6Oa8OLKi+hTXaBYBBRnSf6TAo2NE+nVEyOjczihm
lCq53x/xvrseHc6q5Qsvk4w/XjRjQqVio0s+II4efp8iT12AXxSxOjQ8Ln/mk+QNYcn45LvfSWaN
TTBWs5NWicu/p/Nz2z/ObojW35ulVmFDb5tdE9X6YO0a5TS7SAi0v94x7wYhTguorBacEMl7Lp8E
tXjxJooNRkot/0PJMESYzN3Atq9fCrqZD2j1DSBe8QDkX5iI04oR0YTNdmEOpILK5awJWg9TgW27
CLlewryf1o11AgFM7uAV5CXue7IlguIMfkVvwUXy9KMqjMvED4OiVlO99cUjUQGwMZLr77Mb3aXn
9pL19I8t4Hg1Udj+U4IboJvrBpqcntFtmAQ8Mtb3OTcAr71Xy800WGy4k8e2gXt7/6pgS4D4nlHz
FXXHdlDQXqOdt/Y/oHPmBSaA8VwYBiq51KKIpNrY4pND2qtMwcSwuCoNeyT1+fKDQCNXV6LMW+mQ
jmUnNAbcadvPxLJCCY9D4pO+6kjTvgZcUx3RBCNUtwx5kqyNXu7DJtTI6EYkAFK1Y9POp8k0COKI
ZhxeYfr2ZNZqJvf0cgo9Mf5FvSbeR596smNZxoU8Q31yQj4lPUpGBFjYwPsxZPHJl/q4Jfs4bT+g
Y6zV8nJ3KvHEWp0VCuOylM6tDPP79WtAm+ZSXS5AZub23ne6ALvAyvdLEXinSfOv++wJgyKEiwi1
tXdsvQoNFZT25D17wCNatbEt4VRPOeujm5907msJxZu/sSvEH5Y5a4tKQv9pS0eqnNbvz5qZ9qAz
edYL1en+03UigCYRA1k54J1lJBX7WSgK7asAvdQEKtJ7F6jckI1efCiJPKszUKoq/u4cPIMa37m9
e0FkiByPG9TvyCylskLVAa9GZA6w1QlAmtTTjzpmnCRtbflOT18FdLR24tdmLPuBOAGDovRl557d
NKjCRSqbpfPEaNFD2Tc83ij6GrsnqXdHmLR262EtdIHhi7x6Z/zymCGRPQtRryMcNvVqibqkKjJa
yTJFNYYTnHViFWw46Gmd0Rc9BijPG3im64WeBBYL5j6+uJ/tn2lJHRRbxktkvuQUQrPbR5WE1UzV
U0vRoncKRJCL1uQpKtLoxmjA/+ZGBOlrVWUz5QtHSZYxT1aaGxXjrEFNkwT+QBa86g/0DCI9U3L9
CKOahj3M4bcILV9YpszZkPti+CSz49G3EWdyCoS5YsKLIgLNtVHUaO9mn4wX0UWbKyKJnDN0N3UE
vzM+1aoMY5KniEcAWRHLYTWwQXAgUHbSDpnIahx6AOfxeuFTGihQEOF8zZJdQ5KlYpZfTxTPfZIo
49hOGr3Jyvvhx69y7DKObIcOGamb2Y73ZAFynizWFSLQR7qZEVz/oC4WN/zd0E+T6QbgywsuroR7
BA6Fk1C8Ik/76tUv2nQ+S5HfCnrPXw7B0klrNmJgwJJMzrC2UbKHf0FbK5lN5KXs5SLxFJN8NIvx
vfUgRDVXFwxEl6pIiNlob85d5FNGYu8PRHpNZsVvEM9FNnqElBVW3w1nJvMAbD+oJKtuq3eocp7b
61e5RgUjCMIzFIF9pud1mIgrAOIcnHjK4Gnb5SNYfpAJbyNjtX/0inSq+ooiK7VCkzn79PbC0Nhw
UTDB1z+SZJ/TePzIWFYY4TZX5UflaSXtjkProT7JeF+sxMJ9I5QDqw0Swl9QMBjtZ2IIecovOsLB
uJ4fh17xwl2bsBU/wL8F7hWmhePhqBP9Y36SLfoYtHjKhIudNdeGj7o6hA0ZRfSV7hrraAnSpH6Q
5clVAxrkPyDn2C7DqDKeMlUWd2dtCvTKhLpaPZ2pPNWd/EhW47b4SDUx+r3Hd56TteLvRkCHEAgU
HBQDrQ9/EQQuEhdscmKS5MNdnKJi/9mKeFDQ0USs5Ne15DnFKRViiXcyQWb9oWFjIL9yuvv9ARbA
jYdln3rNLyYDoTswORjLP0aUyYn3kfP/qbchyipk2ZB9C7xdak6mri5FybhL7PIQvziLN9OkqZ1x
1tadcPozfcpxtkjMyqK7rMI3u2yUigw9wtU2GoY3Auso9BEz0YycC+0qEt/trcpYbs71/JTNB7GC
xO5COgL2l6jMhCG4SS78E30GzHzI4h55alfAVdWajCViWeecuBeQWP44v5XEtvJlYqk0kwx7m8og
tSI1AMyP0phAJLFfYpeZj5AWb/54WY4Hlw22C3iZhM1Oq56wppwonbilmUYpbXq/tc8pnnbNmTfR
Kn/Bn1TZefCOLj4KcvT1TFzfn8UjaObKnLOY3lcIm3U/U8J6N1SyQZA8AaFLtQ/yew1yByaXbdlw
7F/n295Fk6cEQ5r74EMZ0iKJLcZ+DJdH1Z2n1tV57Jp27mNdCDV6Tj6fkK2NXCfkr6y/+HOwK/yC
x1s3xU4qaFUDxdPD1OdnSdjbPN3FjNlFcIIzCUR+YZ/ultInSmA57ipR3jMKllup5Lc5Xhq5RRWO
S3vv55lQ7CO7Ayg6g+/PbsY28qPyJ4BockV1dmvbePARFTHC+YZ0i2m+1dMYjG+brsXYkIuYhwZW
XdHySFV9eDJ3D2F5e2N1Y1uoeOWm6wE1NFTPYirh/9tGcyvexFI2vsSgw/k//yv9nMUNxYExP8mB
CD5ZgDpXP9IIsRuTXAll8YwU2OYUQPgLkyutYXYwK5SPXGILgwrEUkhoiu9KfOKoM4VBxGY1rLK4
Rw2Zp2vaOPE/3fLO23c+8o9+BRn643ITqwDFJqEDSDECBGITzJj3p30c5neI37JjfeHNQ2AZIDcy
vQNDLfY3wgSqqKAkwEhbo2/khIZGGgnIJQXeSdkE3mqDtt5RdP0P4YQrAM1GMFY0A1N7ceZW3R0m
l14g6WlFVpjOFxAr73+PvCDvZky9UkowA2Uq7ySEefb1bwgpy/zPTET24IWmGLkC3DK8Qzw5PD5/
1BorH1EYPmvuHFDl2qEh56pjoADa6dGiHDFfxNUpWHSJgjDEq2Vi1iNMvgPR92dlqpcSYrZiuLYi
JpxHBet7CiLgQtFWFk05irxLX6FZY6ZhIGhVCKaHNNyVuCeeCO6Fgzb7QtMp/WYDK+fug+TYJ4f3
BVn/YwUe8cU6TMwO+B3U3nU3TIl/snC3+qP2T8lWkFW6R0hFgbf3k9QATOCZGH2D4ISzOqAvJXoC
fHF1HFAfXom1LrhdBwHUy5+TzKy2QHZlF1rG2+MjQ/DWkb+fyZyktAhXNxmuMtqrLU9LETMxiTuc
SrGIwrbqAlBzf6KsFomER15eHp44RrylDxshXkp1NiBIh1ykCp29VruQ6/yj+CsIiHpDapmt+mXf
WXr4m4RuG9auMDVyfC8dzVRhq8UtOf3DkXR9v10xbLtps/aVrFiHnPEu7BJ2HzJrOb6vJBt9Ag6x
usUiRy/68ov51XNAXc8f20/9Tksp0I8poKRaF5aSnmn0ptm7oXEvjkurmh9jtrk3cJXGP0f1aUVs
dPeZf1Dp+6htTyc8U2vII0urCFqMEoelMhuVIQZh36/LXk1E2B3pdpyvaBJdjRaU+X4DUST9GkW1
/yv/iZLSIaKS7A/kc68atG9xM8B7TAcZXrq5FHSq3qEtONm+/U6qB0lm2Oe4Ck2T5cw5Bc0VEPEC
k5UESU9MwVLBOLb5c6TWVpgcomi+MloQCHyHWfRUd56nYxMKmx5t+3nVFwxKUgM/sdOwRswa2I6v
PHkRB0aoOQz3XCQ1y6PYI5vrIZVeTUYTfixHM+/DaFNgzOHRV86ug+o6qE0Kcwbko//NZmT8AMj7
YJOxAZ7qCV9rqX42YXO9d1BvfyCQLTZprbEZ2oODVz5kXO3Ftn1iN1JNZEk//m6M70IM7icxgZjA
ZAHMc3r3WU7XW2uohruDrRprMAvvDBsoVQox7W/l1v+jXnlsc5V5Q61wkxZQQMmCYi7uKOBfvFf2
UzjjEElaKbkAMnMvHmxk8gI5myFUSHtlNbKqZiucKf9b5w8NneItz0iA2WCIDOqYQeZtYpXt/+NA
XkfShKxKKsbi+AzyOtoucKmk9zUndF6gIgrru+B/A84n2+AIvkPsh8sI4QfOPbld1tlQsi5t0rtE
Dulbmhq3ww6nqzXM23axUAkdGVfZyMf/3B9OK56blQZRHHs0YBGRNnYiLMFwrB+1dAFhbmepqNqn
/p+GtX0MxlMsGfCyUsfUgHASvw6z3w3XtOWds+S2Wey5Y1qQ/HanmfJEsH7GUbq6DxCkaJezyHOC
xGXvKBT/WjXTkZNL6iuybeX8qv8uLiWwKa/JFOU7BENLJpJ7puSbqmq+K0W6Iy7ZuNuSBQyRKDri
HORdUsxVYYq69Oy7i/zML6m2m2Q09XPv2qbeh/ZZ8tgR6qunjT3jBSXRcZM+5U98jWxYAZVeMJhL
C4FQRsVWwbu+cKusw9Fy9EhM6kBETL8SrrBwYuva6tHrrOatDP//ZkfDLfg0jxKijucYIeM3/T/M
OAe64NVbrB27l2ykbHCMm1VXhR/8H54ERvREA0TaorXiok7K/d8vkMC9Qyc0tNxLTzkYfrNLWiUm
3OVr3fZi+J5h4lDJOacElrBW/oNTNQnP9wv/7zRv7sT+XM7fZyQuLzAR8Ghsy6SZnOv/XdZH9Cce
JPe0LP+TernIvuXK3OaMFooi4+44s+CcNFTz3eFI94UkRJIlQEYPbnyncfhJU3Y6xDSaNCCLqJgf
L+T9kTViIVpILFIbrycC1LOiBJW8zma4U/AEHPI0qedEbzhrVb0lynwbKde/T5xL2h2nJoXp8WdP
/Szv3OLfaYuIpI5o5uyH0sT0rKH0VftQvRWPHgRwUrkrHEZ69t8cUoYyV6G0cV86SK/ioECYus76
mxQvsRZptDE6M2BvPAFcsnRg1Z1AYPzE+wabXVY9FT31nT+tgcVjB3vBDXhCqGdcH3Neqem/u2V4
8d4ZuekjUKKrwBjpaoSzy8CMnlLXFA893mjumAgjjL2RkfGpWXm/RMNPpMzouhSJUWAb/cgpViKe
TI2PhscKXE2Zdz0ey4E0Cu98wUWyzNW6zX/0Qzsj4OEEJJgG/imNNaFRq56J3I8V4+Ff5W2PGT5C
VNNht3cQzHRQZRh2TJHgKixDFzRJQD9RPztqOaudQqzXpxMdPikAMz1fVoLOCxgLbYsreiWetrf+
w0MVCalVcj/91hG0vdCBFxKO4L9jZlzWQprO3kwx/1X0eMQ/l8pUG7j9YLzOVwL9Xr7y6G7ezPMY
qzfqYOQm8e5GXKwycq95kVoECGCH8QPt3gr2rK6O0Jj1sXoDdv+TJsJ6xaE/yBxWMVAk2iQ42jd6
VZhFFv/zEQhlIen0yT/em1vASCDb5uZENYjN4a1lgwUAh/CDjaW2tkOiaDp0Gl8HEPyFW/459y/A
Q3iJyg00cB508E6Giuok3EtN517WnpHrknLeWCD4KpX/WmcCZckWo8vrOqtVnUXsMeU1WnFNULNp
dzGL21nYqx+FNpOt+zla1aJIXma36OzoGrYM8Zf4e/k+e4Ho+/8kO9v5hI1YenFghPoObEaIToWd
ztn+D9iBbIPz4McgS1oE8KITBVVW0z2/BF1MXFVBavnDRC/cRS6nMecIYNu98gZti1R1HEI6t1/j
EnnGI3fRPZLFVLuZfRVccgQcKIJznBNGGFtvJ6bDke57qjqp67gyKOW0Di0K96oMrBU0D7pqfBaK
Dd6As7yij+VrQrG5tOTVPekRmqQmov+IBRDvQkyRO3kdwqynGW7XbxMTPDqOtnPJpFSrJywUQjZK
DcOi89PAqzi7v86XM2PPIFk2gPoFIB4oJIlwZ6lI28/p4TPoWeiPDnqLEDqb/FecfQpWy2ulG0GO
Cv6KJLg4rQhlBgkdVkPYaXwLzJPR4GG7pg1/pqKDLsO/nOYhRhiHLQcFYJAJDEjx/MKyJSvfrloe
HzxjclqQMfelbE1CixsUMEQiA/h6dwbqzZ5A0KvccPmTAqBy8SN8XfZweYc1aQGuuVF1PIgNzqW/
hWVmzploXCZHQ23NMJTBs+ticKJ8RNXjYjiI7BH5zyk11TSR1RHiG1yMFYsmj5U+aSHyfhZwzUxu
JTFubriy51igJRkpI7D9oP92mL5ogW8OAWBa9ZHJ43GCF0VbQuhVYYtoAW4Q192EjWt3cmvuWHaK
C5DiGt7m2fPh5VKvB6u/8Hrx7Wc5VLuZB+Jt0iTylOKjso4PbLNABykAJYZPZ+TxWSKrun4Tc3Q9
uJoc0pofEdgdXFfTpWCz9+lVU8/lgsuOSkHk+sMF8HrKYmJ7Zp8FxScCuv89MU9EMZFIyOOdRYe4
kx2UHdTHjr/vkMRL/Tl2l/jYPeMr62ExinhEjbTUw/AYctlw0nnWRGyWSf4lsbMYVAvnWELiu/Dr
CGn4whIe/lmcpn52sckyiN16LSyqvHFATyhPpUMrgef8OhKj1oumh/3lsOciaZRRM+JQWlthG8+y
TIp/3p4duqxBYC3PD/Gr8oXEHkA1mW0Dns5O8oycf+a2YWROuTKl0XicC3DXFlsS6R86Eb7tl/H+
am0q+rjBl7Zz9j4L9MU0gZaRwTLhn5HGN77CjWoYe/vDxICqSfEUJjYABIkHloLXS7lLyuSV4EsD
/0bgtZB+tVK0y946pnAOCZ+UXWETWrujEHy5FiQsMJSN4ZKIzCLB38VY11B/la+Lyb2vzJipjsOL
NsDkwUhdytcZf1yzGJ4i7r0HphU+DoBfdyjjvzrMtHHCcwhpjvYTNl/zfad1WjBjXDl5LoqHXem6
US2Iqwkt2KbRT4kxMFLhZZkd/TCm16F+j0rskmMGpRkdk/FgJDBYspnCPMeZ13KmRWEWTIdMuJXO
sWEuwlpCI1ZvRix0Wf4Lw4RJMrDx2DvZtdkcywR3ODcS0KMz7nYRnq0bMnKJdb5yyGF40b2v61lf
ZRH9hsJU8mK8o8/qxCOa+FrALBhcXC6w7+9seeSJqtIKuKzebZC7bn7iCPBKEMgmIEizXuqGGPt9
0mFf5hjv0cjsjFt9OTQTJHbwxp6JW1WkmTVVwMFzPLawj3ML0f23J/1/e7VnwmpJDidaR1aYAwdL
HOyvv2UFQsWuGGmvheThcKaKhy6hPowC5Zd/O8DNegc6nQYXlH9b+p5vu0wHDMcFGVmmsrwU9P8W
dlTXhklw3/2w4hlOVB7ThSGPE46H7SpR6628rfOZPbaq9RUgFkGUTKXgW6hC5xaC6KFg9IuEe+iW
SZ4D5pS2mE0+7RjEUSshR8Oh+tH+dCd2H3G251VIFjFTbvXwfJ1mY2xNZ9ej4Rp5B4wVgg/GNHiM
T8PCI/pgKZRtZch3iTOYIbCRvZEA+Q1XLuc92ZhTh3tYld9Ay/HZ4/yAcAWE+1kUY3WotAfFT9RC
Oaks6WhuKlmtTTheFz1t8e6Ly1/HXjmOwEiueWuxF96vsElZrV2VxuLObR/RW5JPdpmo8bQrQTYz
MNWwU8qXXSbjxRvm013FzBU1MjMpTGcQt/T9aVzQ6SuYbR9K/tbyNxwXF49LhYUae4J2TOGxGz2E
WPvhJQeIEJOAI5FdNe7vTDzCkPORCn16k8HSZHPyjZu7r64sqxgTnKt9iqkSXN4+Am6Ye59hpysl
trk3/h8tSW0waJHZwTAHmAfhDh7lFA/iMF4b2UoXDnSxnAwawRpK/9/XcQ3j89q25UjOCBSQNA94
oRD0IVjpDLtt9jklHgJPPa3D4WOGg+f81BZ3LkAAQZT8qAV7eVr1tCjWEFgXty+ci2yKqD7brO/9
z1zgfLV9fEp9S77Z8Sh8OXx/SMKI8tq4DaE9qkgqb4D4FXHayN2G3Aj5g0fXNYIn4f4pAfQ4YRnt
3SO2gRIGIlBACIypVbEnSUPId0c4+tXsVcXVrYtErVdwq6D5T2d1tjrZAwm63l0/HNPn3c4HapxH
GXiQbIQcXSBdXKWmQ2ea5/uPvIJywFEkN3QZ4A29rhB9blwEXYqgU+pODGilLbqyFRk2pvAgpbYZ
7Hex98QWYOv29j5y9QEyYHHGx6UClSse5C9AebB0ImJKRqil2401P9Z6QnK2ZHWcuoztxcBrOhfN
4mMWaZAGOyRwvyoan0yHZ51dqNuZKWnveW17MkvqKp6OKQ5NBbF8/wX1FxahZud3T86RzbOTLWF6
mA42DeLxsybxE8SVbzXk3GgCeNkaqpT3oOGMWBMzDLs7vYlt3+RxoKvnH9ZT9yC6RGyOwgEVXJC1
IEzRaPCQzUtY0tQAgpPJ7+OB/5oUpKXoVQyDeopOxzvCmvVWneWIlBPDxD66whqkx5D8EZpN0RBJ
CiMdWu/UpEhGsGfL/oCqR4d733YCaMEVYU1qMLKFgwQsfzt5ylYu0IQR0PwEUIKoMK7fyzdp7w40
GAK5ahpqaZ+ahbMTLuaX/Eapsr7d/PIzT7Tr9nnaP3mN4gDipOO6XxoTrFzj8isZD7xTqlOj01lV
k3yphO/8+o+rEaBBxozyg1bWH0CJTCDJHTVI5zIuUDWfAGZ7bpfgnCmokzPbN//WEuh2M7/1y4P7
5NAx5YE/8MsAzVhclahMbO62k3i0OyjRVsQ6Lduzt0DlCUyNi+lAwCCNvNvdi3WryHeG8ssp/j42
JrE7jYElj3EfD+wuxgCJRpOocQQ+dczp9jZTMhXO6FIfJGHUc8ziTgSmhr+8NLLtN490hEkpN4V4
WMB9Sc9KfEMnvj1S/R5jZiGRvuUuMwS0U34bY5BuW6/nocyCmMYeS3kZfNDg58h/FxGxnuRI2pPW
tQzEEtcHlMkAamWB/N7bO0mMz8Oa4a9wK+f8Z0MGS0ytSkEtXita3+WMUAuprkdTpGrL8N/ufrcq
x5UN8RLB1i/sMK10CGN2F3e9tLodOj//xjoxUH4AHJEB6BDvux6mdlntak06oQGWyF/MAvAWHpgW
9iJmjjVlf7Dx3DdXSz+gJ7LQSc5KD+5qjuCLCmyy3bJwaS2bb26MnVhltZ/q2dSQlHvJ5SsCrg9Q
3vR8y6dMAYKqqxPcxMY1VTHbWknh8eR/GyufKxNaARULus/LmnQ3fTODcNspYbp7iIkX2m1IhIjq
/nt5aSRWxlUBYviDswRghdD/k2BL/IRBz++QIJISVENhEKD7vbX8WGsoQjnpmpTP80vkuLummCmp
GZFaBcU9B0TFlwPGYU3zHKY+XPWilLvSVnNcrjjtYfQRKVqMMGeFRnor9mG+kDHmtprQ9lkgjtpH
nZR661rW7UKTFpraJzwRDkqkx4TEC3XLMjr1JYOAJdmWT5Jm9x6gfu8z3gY7hgAr6kPoln8H6tTe
ZTrx0/CDy+SYHYIMU6CZwwsx0kBrc+EDkP3oJ2OS2UKwvEzFbUcqfLAgZiEbgNaFapVV4p+dV3i1
m0hPQzRyGc0LJKTb7/VMlJb+p/YtCG9wpcF5flLo5DZow8obTi3oz2tmNboFoTxe+Vn23VZMX2o6
NbXqbi1iHshUbnNW4EcXUvIgG6XVnZZ8uWrearEhSrNdpkknmPcc3djPhgGTEcJtExfJVmaG7tVk
4pqmNTFkr7MfqQg55lfr3bNA5/hI7B2d+gtwmajZkR9wEPsuxm4iG1gCWMFS/DkV0d8IyrDgD3cQ
EN+cNFaRAyUTe9MigULA/z+GKhfeOAPU16O6v1IpNwha3nMcBkm7DjfGzLrb9aZvCczJ+eO8didH
TVWcikTVAjLEKPaWL25drsnz3k/X87Eb0yyBkPy2XXmHyS+5nZt4zKnze4IuiPajiOBIhBQVNjk9
ABjL64DUTLinOK8C9K3RSn1tBaPxkE1vKwN0X/xXQ638B1mA4sn2ezMXGvK2Vp2YokEmwJEB3E/L
s37BdY6GM1oMk9Y8SS03KAlNhU+KnzwFD2UW+HNT9Q0TzlFUtjIOp+rgxxLgU2lMkdqTUutwc0jK
/BRpzNed8wGUNKRRr9h5KQIUmWMN5TxopW+2NwVcOW+pyaK/3/zWyp/LM2iueJM7as9Ao84YeQu3
xksjpY8rma/L54HpsF4/trioGIlrW/nVljZ6IobBaOXYaoYMhEzM78ql/GjDyWJn0LrY0WeAiB2p
CLeu0uXsYBR5EvhNntZI0rHURxeGLJ/n5ylb7jI+4JXYmQe2V3/eTQ7TjTuwLMp6kRijphhUvP4V
Y4vV5xrBe9q9eMA+LtEefEyIkHMLztD4XpjktINZDUwWQ/oeJG3LCc7ginbv5x+Un4zlKjiiJhaL
+y7WYs11jjCgtDXsZqXG2M5d/Q5SasfzNFHkbhXEFozqJckSL0bZOMWuvqSgQYVA4m4haDLl3viY
w2K7kZHKW3ye8MxuCgyeErEKoY2H489ST5zirpkHrSg6zj8y9ZqWfLNJpLE8xorvER1wTa8R7w5i
OXlJFuysdHpadjTGudYLTx007KYwuUyKVbUqWi7WXaPNEqHjm9kpa+e3KVMjnU1a8DYj8CjC5+Ni
TyCwekF7m/viSEAybtT7/YaN0uXVLtwASbQFunAoaiToG2CnP3Hb7H0Mv/I3lM8xmXAn93uWxhOu
cwRNP8cBte16iP7QlyxyfZuOnZA6K4pKsjKd0WJi8W78VlQTPw98ZsK9zfCTEEPpXAruWG+urABv
kF4Xf9sNyAB0IZFjvCjxUqzxwareC7I+P38Vi0YYokXTDPHFF/pPZZe1q/NuL0F9JMDwDcOOqx5J
SS8/1aefZ48v+v+N43pPTwqF/gC3Ixe0S+ZPKgFOTraiEA9wuAItQ+UqiispJpuh8f5XhXigyikV
z76/HMpHpgEAb0ayNvswX4t5UbdC6zNBqvfJb6VWugUKhYg6QjauahqUxh8ZRFczGg3qpqT5ZNt7
1hlHco9FRijcjNYyeBLrQ8+wFERLRxRWMJF1NHdNu9K5wmkWQl91mkybA5hHPUDFY/9On6drr3ME
SgZk8gkzrseWMIji7qZABNK+259A47pj+764Q75Ryd0SJijoRSAgoD+gf+gvLJtoeCZT1v1wb4GQ
2aOw8/LaJW3zX8IyGjgVYkZLjvwieTNOEIAWbKviBYlXeBGTLGOrrvqRA28wOhXaEk4yVFCmIRht
0DPrbOOpW2yqHI4o+PnzdEtHHmVjIgXEjM7KZ/fsDFVoBN4Zf7nXb1+eWCrM1KJssK3E7ACKNzek
ZBi40L3hsgJel/CXwHwSOGWhXNJvsLhe2LE9xh9NTl0+PCdrJL0MZl4qGpqciF4PiZ3fXVfgRzQY
rjcmAf28T8kNl7dl8/91N0F6cwkTrpA4lLUQa+s8Vl1EEniWKw6aCGA0r5sQ934880lMO2gfpW5i
pAQCnZ4ZYR4PPLmLLjMEdU2pGjjeoyPS0KE1jUzpapVqCLph3L4H5B3lMhEIYXtgPR6fg+oNGuM+
bn0axTA6hfHdvM1EX7RxMlH/tDGBOmgBa6/IRbVwx0ndThv2BieMFnPEBCknWDvW+vmzBV2P87UC
GUuttl6ZzYeFdIk3/v/yzUTgsbYM3RCTWqq7+yiA6a9zyUx8P3GqczJHhd9Fq6oxNiOQHebDlI8L
0/SYpIDzrZHpzwQ8YGDTfPs283CTsnv76H62869Q9j/B6FLHn48/cf8wX4FNQ9Uh2rTYuGBh0wxb
MaA0jz+LBA9EJCm1QODHC3GCIkAay42mmTR+p669KaYQtUDIh/sX4oTa3ydETahymg20ujShoU7v
cEL894N9ZxaZCiqhk6E+7AbSnjdeDqPy2QbjIkO/8HFVt293M9+401ITTeHOxg7t/Uy2RGmq669R
4G3yDKIOEAgLw5E8Ke7zX5N/kt+q6j+yCYKPCOD/Ubs1A0pPvqOxn05KC5PLzEoXurzvOmolcrX2
j3tIWyBPAg3k96ZsqB+ads3FyMCTUjtXbocYjYmX2/EssFLY7PLtaCSCWpAWqaQ4JMP+1tkvpyCv
mkVgaBElAGo9pJkeGFM+0pa+ShrmsgqCVPDaNMn6VU/3BcnSiBIzdg6xdknSiD8K9TwmDbwRZ98U
o6tHJV3TJElhxFT2lMIoHZaxrDdXUJ1zXjNvLg7OCLvPZnHl7RIOBuKzQ0z9jR+DlpbSAkSr7L5K
acMsUICItNJKlD713BwPZ/j1G8poo9w5bYTFaAK5yHbT85ayH9Zvuf2MiTsIJlQQDLTXjDDc3/Fe
AO0K4k8cftCk7uFekvwQsraQQnzOiBPckoRRn/AIkAvZH8nPbDzSndYKhxMYV/YXkCR+9HLNWrcF
sQ1NQ+BkAxFxq3PBDC2OJ89MH+MXOF1EOEca2gX0zaCWFzKBGz77bnpsV5/cVoxqMa+ukwuKSkLH
Mff9Ks8mY5KaCCErDAn0UWlmacqxlE/nyUkh389WSH5CWylvxc/Ii7/nZrxhuIJlHh76xRfKL1x/
2WoU9VabZ2J3ZbEowgoomdZIbWueDUbKo72qAnEpRLfCG4znicii4dT530AsJP054oqQLMlXVlN2
7lPhVLxHnFdATzxy96yKuT36+a6aoMBISajQz+byFBN4A2c9KhQBt5aK59rvAKkI8ASW8ym6/37o
UQDzCDsyrOjgBgXc2WQdzpbU6d7sR5hZo/YGsDO4Z8XKaQPceGVhsN1gSw1RJa251f3rdqrZP3PY
FlR9hx0hrKmdEZC8l1WrV6DrkgNMZyLUwhuVUH1QsS7Qow8DHNFLnA7VaSHARWAMPwTjmScCnPer
3bDFaqs+45HZLaQRZKXE1cnDfV04LM55Jxuezh0DU2Tqsw45QOa/t6NiN1PBbbjiwKDkO3GAKCXr
E29+1ZxAoFG4Di0OmaHvg5n7ak/EI4WHTu5ccILGJs5YeQ0QeluE84gjyyaLzHMrftR7g9LjL/vB
lMWgaRzjNW5+heZd/9zUM2bndq2Z43J+ZaC7y2b5fLwDfw8c0Jeg5pCcXwDjNAmRtFCCv9Yl6ftg
LoPx72n14yRXtSMdO7u4wCPZlSjX/8RzeyhR1Da/AZ+1t6YZMekrgJFD+Ii1Oq6qy7aZgsEvzrRT
k5p5eDB+gKI3tZ6v0hLrdac4rRKnrYfu8gGU1m/NsOAanfIqlVsK01YCAJQSJ31FzAKcYcCD0B6/
0HgxfzlE6Cykzxh5Q9v98gMPR/8pXoQpc5O+Pugtt97BMjbxX3mD3Mq4BjjvQxaZ2rfvSe0NXXEV
cjvOa/0xWl/5YZMsCiBJkGGpPcsXE/T3+N/gF2LFj4YnnOuh69hKwrZcMPJH/yZFdMjg5PV/VuNs
s39jDuG7AgzlTAltMMtu5OgEZ54alQ0be+wVSAqHoAat/ry5dUiA1du7jLnReDQD8osHo4KNcrQw
wsTw+VsCMItagWcBKRauH/JY9KLHFT2HkCmC85rbt1hal3QMyZejT6/6ZZTXVnfKHKLJpho4n5s4
gNzeWJFP15y/P6qsD5iFNmmiUwD3/XDBWUWALC+bLTcuPCsOEhhuksTJ2oDTlqJ1ARJWFpCmcwLo
lnA5TGTOcw/wFYS0sMrU/DHduLY1olOeg0n3WU7587OPq/KBb+Wj9Xhxu+tnhc0RHMrF/RZRreBB
m1DRd0icOkmhfcDCiHwECKkaaN40jrtcxy0GP6Sgyku0cNaz3XArmKlPlHCXqC0f7qefxHLalE1S
Xu+2W853tH9VbArOZPJCEdGyEsUcjQdcyF9Y2lzYPTedwp56Iev47FeWxR0IYo1hiGy2KgFC5Jy2
zR7IjyurnvoZiOcs20Vyb3FrR0/nzZZgMPq4u5CKzpYAZW/zBnDuHulBYvyXW2GY3PsZPnw/EUjN
vuFmVmSaK2aii+/YwA2nLMflxvXhA1lXatK2nmKA1/1+kZEgK9Z8qgGUnsCTuoT5v4nE4TWoBpTD
3mDqokd20le+JIloQqZGViGx1I7exN0jk13EXH9r3m9s5RhpHVR4a6fKufjRylBmhmSm8FKljMvW
vPTnXT2VMIBlaYitW/eMx3ubQMuDWjqC6WwBF1ktmuccDs/rpiW2sE9mrN13xdzcObtFfEvyic6a
VnJD9Ns0C8aiyx9xBEaOoMxAGX0TQh02pIN5QqdFhCDIIIwqoLjyl/3sEL/ZMoFk3WekPpF1VFFu
FvHRkgJzFsBLFbfpFcYCgwxhrelrIXzNk7NjhnIXDoRrKVX+yAC4G2E2ONwsWjsDFKBcf9bf1r6A
Xw+OkG9+BdxE5USLb2qCtLmY/R4ySEhm2L+ol2Hfrf8e3sgCf9sbGZKumio7RESZftJLXnOEtytj
soV5UHjH56w0fYLBWaBRV+4oiWXURscSbkVB4XpycjiUNhrXxwUkFbTPPsgem9Bt5bdaDf+23VHM
+fMj+5R8F9IYKrMQalyG3lTlktGs9oD9OkG2O2l43jVMD/cUhP7fb7Ps2Zbd9IRe18BVtXbvYNp9
M7+/5deB+vbmmBa6mgkKUpV1mo8ruRqb4XSCXgvaeStwH+jOLTQPP0mYwYkzGNafSlaN3N65bRLF
6cuTbOqpixCQ4e9bblVVyZ+zPuePAyR8X9Wbppscr+YmQrS5uMMRQzk/klstHZTDCVJvhVoE8vve
6V2x0DeLV5dB1y0w6UNkyc6xDfRDGdRUTTYdCcEZEHaAPqchjuUz50UVG589ZRzVdgHZCC7l9TXm
Gf3O25RxYo2RwByM+p7A0KyExhdxlHP/Tvi6ZKMSabVMty8vDS3CP98FqJE8WQkpydj8FkDRWgvJ
lvAn7WxV7fqV65YLWlIvUCiuQI+C8SXDAKYUnOe1HARVSefD4hlEPz5wrPwW8zdQdTq5iplGYRa9
pwzMPkDBwQHav8FPNToHQ2Hi7WsgEflLtEh9YIB+qGtwArT6MaaAU+UfsEvHHfX7skEHZ0z7AGQv
PrWN74spYdwnsw48GIESjeChv6V/QxlkietA72MGqV7ah+1rIFXNzAjbJBIvAHCKIaWoQ5jrLOUh
zkxutnmILS//KzodQy7ft97UDD0JEVlFKdzgbRwG1lhmiea/sV1TZXExCDV8tNUf6p11w/t9S0Fr
wEl1130LdEejDJDZ/BdWR2+4Gsyq8gI9btkgQwsBrpx/1NITSISqJn0/6Z1YK39Vg6ij2/IPxuyI
QGuP2oPCzFKeP6SQCWKcUCyTL3oEkTNy1ihHd/BW5qnw7/bhCsC8lBCaQ8K1M6VVOZcMHBFOtGaF
JbTsMCtVKObBShrXonXwIcO1FNk/C50Yv5zMN0+kxverYrr/e6Dow1GIo/154DRWLyOzsR8P65+5
nSbAP9KeyRXL/6bSh72sKZr0umX/RefrhOoVvEDrX6Twu1TDknel1yGgwSo18/aW8iP3P/QoS+uy
p6hTvysp/ynnqy/8mZBs+L4R162aEm9Jh0/ZOyqpw/OzOmrFO+aJOy8+k4yD/wV0dfYNPQgWcTAF
sU4VtDqCICWNV6HeoIpczK42/phAIdZ8XvBnJTNp7QU9V5hwkzYYBUUUI0sO4MYw/TeMV7tM03FP
Gyw7lh+DAD4qYPJCLcrnRqxb/omQIU6pwcDOpbM0gJufbYUh3TB+4UiNHfrNlCbl/EKXRKIPrXkS
q85PGsVp7zNBz/hDK5n47pWOHZUT3dAVImto/TNTAUfoqjNrR+WcE553oMcOc6oVMksGZ7biDDR7
oupYxy2WMJe4/9E86sEHPBlJZucjYc1nLC+Ow/dibPmJO0ttWGVvidmGV5V2Y/WxBzDrwGw09zMZ
AWN3Zx6vfWIFhFvt4bN3IlRvsQmTgeHKDXbv5MVbfs8Kh1IpRYlYYEfg6qY99oFW3JSRAsxVPW7K
w8VLdXBDEXrGv2Y0tQApGDsIxSNU82tcIFWP9GtBZ9kTBC2TJ4kE3KJnPu5IZP0/eiEo+X+qsMxy
vcIm73KdDX0VRrLYYbADHYGzwwpyf7N1Gwt2z8ZlAOvmcnc3BQuHeYCPPgFkJPSpRFeshJaY+ehL
jhcF7h68R9bahK5/Z2FkDTA8xQoRlo8VZ56w0xLofpnsxjMYd00Sx8+nQRQyOhTezeliBH+P1prU
h6mizQjs9mSwk44H7DI1YtIzdA33FTC0C10l2Hxs+lGHvhRMBjAoy3b6QCdVuWl9yn/5gYa1zkej
M1K9+P8wCSqQ2pffsEtuCT6SXMTKbIzoMOcjZ9tfg+ENkk8++kJwi2ilKQk37Vt6xgqrruB54WMv
ap4WM5ci9CcILVfVbuTHj+gMhIsY3kWuNxj+vD4pk5w0YGjKw0f+wiHDon8yRcEdpXEwlxgt1iYF
UJkfs7WAjZgq3QpcTOvBJJHgB1sLnegKWv0yBSe6vRWxi4wndJoE1PKpZNkx98BRbyhWimBcASCS
+pgmUEUvqSDiobAgas4RQ0pulnSgVxCS1UifRqhv7cm6ODRLKsvEvurIdGgRGUpXv5QQ6qkGpSqB
HmHJszXrQ6J9aIg8fl00Qw+6PePdqbXcmMbQ/bjtI7WL884oQAX2WrnQJKWsG1SDCk/EGssDstjj
txMmYFvheWzkpJ5pW5K0MHHlVlFrrn9Kx+onwVKkJ0XDE0W9ZYEJXO0iRq1/darnwMxhUqpRHRwW
24bapa7WxQOCagSs0RvoBPx2dhXQo1ghLG7n6gGJyQNn/sSPETyxCkNkWSQqTtmejOq83yvN2145
Okn8wC+oJG6Le/3JucUJMdXqJ4uRZMQWrBiWV4KmCjs+C4NNpH38/m/aYIkIdS8RmGbaNhApJTdC
7NzlcXFg36m1mPxjmW1O0nowHfPPitOAZpZAZ5B9bkRxpbok5WDFNYpc9MS1yD4Rk8qYmfthOeA9
UaPsANeXd8n2U6EUGMQICHo7ZYySfcMqprhdPFSxK/uvQIw4TJ0W9tm5VcMUuS/EzhoHez7a8nj4
rQDmCwwZI0N8L61Qy1HqV6T3U3wkw4bRq3uw9OdZFQkXKGfaT09xJdKxJj9d+S7n2JrLmCuZCEqL
K2oX4o8l04G8WMdL6qIWZ4wADEIZeUcItT40sdXB781m2fGbM55rvRPGn8TUgmB3GDjFmYPFIbAo
Bf4z9LkLTfXdJKYgxdh1iw624+N8VneBr7O3klzMCjbMb3fkjMXQhFVNuNUxbQKu2lFcnXhOIVCJ
XZvV5eR5poycXYhkFQQW87J5QQEaSMBPPjXnrKBeaVbNisuWCDI9DHshoc8wdHMLyLUhxut/Yng2
g27knVyRUbVCrAtewA+CFt6lFMmred60ZOYww9baeAKjIHPsUD5xNqXJ4yb7h+AXfX7XzOi+Fp9w
shLpp6vHoFxEmUbvUue79sOMJMuqTnmZ+F0gLipaDD33O3NDSPpH2so2NoqGyVSln1Wgi/XkueCZ
7emxH0DzlhxIdWDBTa3oqXU2ZdXkDYMcbQDJdjmUCdp3qeYcLyMr7pVSZV8bAfZHqUTAbv0/C28s
IQjXwwmkKYRlwB5EO3Ovqpt1piVVYv1cFQ6i956IzrU2rPIIBARfkc5ajTJqHQPgUrAiAT5UaMtd
KEMwZusbRG+yn3NIbk3sCUpi46L+BxO0opy9PInZDGqMPR7h52lh+SkOY/N2hP/gphtCoRmCeIel
0wR8imu4H1EsNVdhYCv4ddW1+Nna9UHxxYNThHTfX206aCdoXkYxhDMlLFveEvdFWrdpquD1E806
mDwbdfnUlM/8aYUVQMUlvDpayj57W7UO56Vld4GUmsevlQF806d/oQbVo4KGV3uMozHl7/N1cn3H
qE54EqKcDB+0ldNpg2hD9cy6TH6XNMX2Ra+r+OQwpWyqn73jFx9pRAvwUKW3D/GR521EuLoJGV56
6jxQuGpNf301lahYg9rlfKd84y62WXC3J0vW+n00PwBa4Mmvw3LWXvu8Unz3RL++cZtut92sblQ1
0FsGf0WWrUrWJUTtE5siUCZee7lSX5fPk6JBk7+bMrXmiSYfTthUI+FXDJiRX0GcrwBjQEPPHUmF
7+s+0vjFektl32j0yFB+ugAQmKwKDaM3nm2x39zNQ3QNahzYoWkHx8BNcKQxQRiXxNkUqGIqZihD
2gL06a0G3fMWq8S+LqktupJIMmDBNgnLzVe+Q2CxYeacW3w4B6VfiNgH81WPOaj9yWoUDMJ6bYGL
dvrYz8A2B9yDx6uOBxv/bcOvizzpIHF+BTt8L75qfmO5rig7MvpxD/yLGwIiM7M1iSvMR3Z02hg+
ytVUrG+MJwYUOY7/8LgPSsAIfbwaVJHYBWprt0MpURihyLBcNZQZ3p1W9p5pZtgChcZu0eJhnVK8
fMmER15YRs/sIZwzv9NapUYrdsxIqSesQ2gDe1U224eU2BRU4VqTCuGKXoi6OW28ntZvntjxovwp
HHySuGgYLgfBqOjV0V2617mjdN6ryIJ8uNLU5Al7qWfhIwXPnn2EZ2CQqLBCiAFEUgrD7z8R5DvZ
OBPp5cOgWrs2GWqyoZXsONy25IM0LcDm0QtEAFocu4KuvQbKSNlAah2H8EfrJmK0mdfYTDyQF6os
aJTVo9sJ/s2sSKz9fJaSyzB91aXkThIaLVoyaoawx3FQtn0YlYA++7xQsDrdYf4dCj8jbtMheDB6
sv44IRk98pEq2QU+wNmK/5z+CIDUvN4nXPSiJgbQlzwFv5PjnI2mm10fKMRHJT7Cq2havuwTeaFe
Qro373egAGoMQ7V5eyGN0YnV4d0JR79/9BlPeXOTT03VgrYslsTZgjRqL8m482VbCPMvpUBhNLvP
86KY8fkjFN3iVEVatHTJIcV7Q9Tf68FPH4+xCMlhj92Hzh4/NigXfUYQkljYJEJOZ/p4tdTG4GuM
GBvzJKj2vMlyccVajj78cGFCquXNH9RtUY7JSnPy0ex+ffwv2RP68OkAamM09uOuReHjOsuGwmKr
v7Qwzh02UC+td4Giof9k44y/BTwCtc37OfY1AebTYvjKof0nNUIoLQ04e1JNCCG/IUDHdhylAkPH
ZT1niurwxngZM1SHz3crnTWDK0wISAWQmfw2KrqVJk4zrTa8Th9jYNnWepaFjU4/o/2iFs0HnHuT
4ofAOt8kCaZxrO8sCBugoWyq60irwEhQZwDfXm0T4/5HFij9FvcfWMGxZP0dKOKpLHcPGKdj/XRH
09C2V9hY1mkO/DgrRIkBAKtkl/xpxv0rHKwlsSoO7VKMOdRaJlI3SiqszkCWxBGJgK7KPsHctNsx
GKkywHcVscQNMgMjtVMb00X4jLRsWaX9II/SK99Fip5GaYX4acqGLxO4IvnTKVVd+YY8Gr8Jmy8l
3v2zen46w7MhcAVXFwC08HOWV4bzZ3KIOLHU23M/i8WMRbzVJqfdhlE4VzZOUiqOZIb6Gjwfd+xg
We8BBc69bspZ1fnbRdqWtcC8ExOyoknyJCU9oOef35srugdveg8kdVFrv83v8qDV4kUMIn8MvhHo
vqFQmNiMkzZdHj5zLWT8dl/vbddsvkpwUSp77V4ugpR+/WsrvEWfiFdUVfRVTH407Odq3WVNMX1s
wwQY6XSlu39543hBeojI5h7VF+OBguALuJ/gTJNhmkGMunlCeujB54chiVIZhJS2s7JJC6ot0sAV
Ff1DjGMDsXqtJ79IAZYoWQ34ZyaKW9u6wQ6GLMAyffVJfekGv21MYlCDveY73UTwgfPSl4jDi/pI
rRdTjdqvHSEWkJcTjEA+IEO0jQLmqCUSRhAlLuiGntPA891ZN1qLz15vOK2pkdf3cM+Sv8x3tKFC
1KoA5RlEZlqUzCQj0EoQoYfWSkRgk/sRcOUFb2UF/FEhGzf1N4inpta73+jM3V28hw7OYEeZnECL
1pKT9BtfLNVWUUnRNU/zODxNTHwTwC6RaYOJM7KERw2Hkz2nS/fJmdMysrCsEexfgXBf0gNGA9QR
I7V8N0eNr0UA+GUu8grsSxaFbIrB2tf2TzsFElFI0crc3yi35ub+z8SeAPl9ChUO4EuyjQppSPg0
2tc4FFnVYW3nCMz2A2nO7/Bopku59JmhfmUvTxlbtMWGUS8WRmEyqZH9WZfJULItnZOOXqNjDIYF
TzECQbiC323YNGkLd795TQSLINTbOmcP9bglunOcx1ygEpvePtM6Az2659+hWExGQz6UEP5DPprY
LP2MnQnUCODn6I3RIZNXw/kT7j9x7teGxiZrWnb8DcuedslmoTeLorAK4MIn6rVoXy41sN5g5fx4
zWS3BZ/9Zj0zzke+AdavA+GrCWkIQe4hcjC5RWT1tgio7M+zG2Vbut1UwBT+gFJ6/eHSs+/e26Wj
6W/nLSRw3Fv7VFR0eJXRgnsYzJnr0ALipD7MTXo8pK1RmEiFv53O4633nq9+SMhQVQ20I8/97G1i
RXi2j9ILjqsjJmSIcCw2QlSXuNiqTRoi7mEroZzMNCPhqQOsT1wi7UHLGecENAmnFaNahGsXFZ/A
JFdwHwV3Rvf3T6EdUlgs/DkSsq7ZfpV35ipN25IxwGG5Joy6hUZSI0mo/TEh2CRB9Fh5NXpX68qf
gck+IRNyC9yRNsAqN9YY6o0tmKgzd5H270277WFEa4cxsogUmtlWNT6+qVBroWbzqktQTq0d9r62
7n3cGF0qGzifD9vq2IAqVbkGt1rr3neR7REaDvrZF+ilVR5m95xB9cdLEYaWTDCCbg16/1F7Hz6d
PpUT8J6bwPxEKpV+vVI85sV58JywBbIe0enSD93ltXWImnrbCL8MoElDTrpnPbGdJ8bL2FqZrR34
ehcgK+EfOmRbp0ZJeSIlPo17we5KO/RKLA8NpiZCJMJMFYrel2pBE4XRzox4jqcrvVHrTsPqa1N0
mueRW2CJtNjNjKXdMgyGJRLsT3NurMPYdFkvq3FpXKBi1mRZczCsuYU/3g6epcUafH6HubXhGoGy
W0Za771v9Spk9JF0fJLNBWdsgrywADALR9q6NwBCWC0Xd6vQspc5p6WgBXcvPemRxWpY+loVh2OY
6Fce/BaKBma38KuY/Ti/e4AkV7/2UB8HX+C+wLYUx1A8aKdf2cRDCDD2XXB48hGKt9GA5ZUykxLF
KjZwfTTwDRzoTa2n6+JbP52MD1RtlUUEZtPUiM79msx6sT+DGmSeBm60f/CvVGMrD10fSVL85af7
8FDL1eOWyJzeYxiYoLnZqRQ5XYlU5QlhC3tbi5qsn4S9xlqDvEO5JMcAHUPqblOCrUhMI1MmInAI
GOdcbf9EnWTPX6sDLWLvGZY89lFYVOkXYwlDxqNSZhhNeF5XG2V1H06uPvM9RXYTQz5hKoeTEkDz
4X1fOKTI9m90+56aUyHCNxz5OKlnC1QNA9eFZEmTox/EdLwhoqS96fkEHq/bB1sed2cCfwZ0PpRe
uF9wN0r1mu4ShGIKM1HHcxj57ChwpfSQay1hT99HQ/iJ3v//OY9txXzaMVqe5uX8oOYymD7PjRhd
jSOwu/TxaDxjyQLM4TduwUQtZR/IyRVxO+EDbiOS0ExP+XgD7F+GLn78k/I0m3Ay2qfjmOb1tOTU
ScHTF1FItRNp96E6vd8pJejJdhjyM/N9bO2mqbQVFeZV8fU61NaNZ1EGQpmY/oPq3L9lubLhjj/O
8kkv/cjwNl8dE96CokjVPbGUulk+pkKao42vPZ1hulAmW/tiI6ItpF+/EgByykB5mbdPEa9fFUkm
5Ub1rwOV6KnVfysWMMQhYnNQabbUuFinl40f/Dy87RU1bNSQBXfDeJGRSfVo/a0w9gSzMv8FfTEt
aFFIOjuGXldL+2fzmCKRvPEq9Kw4BakUm7r4tGyt8kGdoUpFONLGuFzZwfyyl+UW+uTg9LMrVw0Q
7984JiRI+6Fch+78qr/DdT4NBx3QIoknSbDg1otbY7oTXU95+jVHjwCz2SzLdTcPjFtSjvFU20v5
QGXzzV4XB0K9n8mQifKIuET+D8gzJfe2y5GVo/DBbxG+G0GVi5etM8+d2kehyeeyfkMPCdGgTZu9
fFoHTsMMp08iZXOuDez2UTRXqm8GiFfaiIaG6r8yDP3Yh2MG3MRmiiEqkjslUdgvErS8gA7bAUID
oCcxehwY5NM+J7PkDKD6fsiOc1If64wmHuKiz3pan07PiD/9rLw5ST5s7IefDkosGdN9cLV/Yzg2
J/wTum7JQ3k7ou2LBcQaH+6Uv9bRcPBASFeLaMSrwfxgUaH20ts5OP5SmA5xrhRo+7T5KQ0bak/q
fr6nUwmasMIlg3bVtr6xi4Ii6smvMHuPgvnbUJHnk2KFFk5AD22ObYR91gWRBHDcd3m3GBK6C84z
kMvthjlfg/fUSZdCdZ4ToMI4iwQ/izTQr2ieSaCz6UYJW2WFrxsvjjucqvbwWEsojt7ju8b44C+n
Ni1gbPQh87Q1WzJX8YrrZ58wlbKm78r4ATom9Y5I0lVSMvlXf+g8mWQWRwcnGkZkFAVjQuvgmntl
pHjOwBunNPuyAzTv21SBjR28Yj9Rhp77p0X6ox3RzEX/0s5zQbjlYI2yQDyKB6VHX02ZH3vNXv6b
FdJKBuDimTnqeo9P84zgl5xt8KNTGJj6MRJfg965xnGvodV3ls4rGK4BHBPQIerDONor5rm3tOwI
deKGhHNojkfKuK9FKWnMYM+U6QnnWyWnHBRhpLERu/CCzcfb1i1NKfH0bNIarOCdW2GRvctgy49V
xctWnxpByI+Z9G0VgjJUtn6p2FaAwXvftVnLrx4DY3klOxm8PBWi85tqTv6QpoMY9thfYRVLHI1v
6bK0rKVg9T5Mm2i8RHlW5s3YRawKnSm4evhgHic8dyIxwKrA8+I9bZs6w77By7bQavL8RAlfAmuX
xU/9anona39fA3i8uAmYuJCHnPSM5a8UISEddmcrzi/UEKiVaya0+orPxmPRZ46JvBGhxyfUSY0z
u3xmeb/YttFC9Bg1+5gfBNe61xmblCMhsPGXDRQaux/GdKlag7dzbee+mD0a2+zyCwuRub1A2vEA
LKryVghPp1lCpDpcxazHT/PWEsmqXQRj+8Tenx97OnHntUTFsvUEUX5W6HIXrukfHORYRpRF11vR
yu/X2m8SLGQBLznqFNzQopck8DpWGhAySBBTyD0GLkG3PeMjvYBy6SE0cDaYsqa2W0jSV6W7xN7h
8IIBG/AcReoBrNJORojmKo0wAaXAptXRq++aA2kY61Iw+SjeV/zaZKbxWT7iWUgcggqvA6lBvU/C
1HZ2UVRq4ia5xw0bM470Y6nL6AoMY739+tewgWrkVbb9Thhxc+LygE8v1N3HBRg7kOvpLB2qbpM0
pL1EoYl0s4xbYz3za+sXLzTXVIh0G8wkviAHhjiG12jOAw3HCd8nu+cxu5KhFEg7CTumUztzZcKS
d/QT59hfIhEF1TWY7h7uX/szGnTXCqL/slSUFGaNvM7mGWpX3jC8+WmXvoKYYpWDgtdDmlX0gYvD
zaSHqmLKUYhiyMjzPtfaHODqjAj0GXky4FjaS56qPY8pf9jC0AFaeczSoszsECWazvDWJeZrX4z5
KeFvjI5SQlbnCtZ5TIZ8n4kgkUvHifU4r3iPxFZD91N4UcKg5NnYOUPlAEnthM1XI+Sp2qxK21MV
MHmc64+GErL3QsWaX7HUwc85gxjJ6VEH2JpG46GMDfDm5zSmwmSQ5+cVq7JjpbdIAIijg/8VSLep
dbX9XLEcAX0Nfb1SHgWDGNRIUVLkiL01+te82ops2pDR2foRKnq015A6biZyhovpLYRTwwWK9S57
7cUQtt9p+Q804bxSEq02cXWK+5ieqf3rpI98BW/Xuzdq+w3qjt+yQWv2nOGke5psbfg4ZFV5AdJM
A0VVgaQrbFEzs7rU3SFtxd/yLFPRGyC9Q2UQHV+gxcOxY/JwfxnFYOa6JxbUW3cfCfjlkFIOLfVg
s4fTJO1LewByVmeyb6ctN1QuxGRYOg603ZSRMICi9UrO2KpIE45ZJMs0m1PPy4Xdf4n301u8lKxk
yukhOB3LPC2lg/3OAZ7OFR3uxEXtXqGN5Klde+tKt/0+C4iAgpIKn2vXUl3+8o01PrK3A76FXevV
5f+/e3S3IPiCHmk5qLYY5aaDw8tAg0ZWsvDHCELrbrXOHj9u0NLBEIdRVXGp0BfjBMFjaY3CfNaA
+e3Qdqt7txH14TzYlHVCbuIP/nOZaUWGdcxD2LzxGx++1cDWc4P0B8Wt+aj2e0fpXy6ChiU0MA7G
hPD5afr4WXVBs9kVgcp18xuxd0k+aEIoojXKSNXcJ00BOK+g9rNvSqbuYoDYVQ19cowzpq8QMaXk
qsqUZS6NO9hY87/+d9XeUTHGIbdDCTkbAXZQ+FzVWXyviuUYjsPc8JqfpAuSvsf0wXXDiCxvM8d2
lhh1BlFaqmB1d+15ZLdhdhZA9lGwEZK+7rLM6urZ+fbZVqe2qNJOr0vZ9UZv1JSHC7aN79pR2Kj1
1IWdYpEL30clJ7kqc1iUHSpY4w6egSyMVFibablwfPgJhESernsdVEvrwWSumyMV3NzGxLUSjG/9
Hvy4aTcVoZLvEr4yM3O0XBQWXcSZ4q17pq6d6GYp4rFDdo5umdDc628iY9VCzWoaXGaWsRB75i6t
9PO7XVX3+dQ4wfpKoXL2MsT9L8igMqzzjnYu7RhScls2V/kGgjdsz7o1qdxT0GpFpZrTAtDFNmCU
51UKgTHTVE3dVonyyQuQBAobpfWimMyK7noOIQgfWivqjIWeW9CeWWyWFxWpWBzVW1gltG6sh9HP
hyc0sxPPWe2bCgD0LL31jhBo8namXVgb290WjoWkVlmHAxNPuIPfmrxicGRGVzw4EFYoKPdfyxSb
D8tXRaSs/EyCSCx+TqLYZ4LCsvyLpQhxR+eTGDWYtdLp6wA6oKsyiCCClajthLbrXBHsaJyRdA7G
Z2mDiEzoXrOPb0lnqLP2ufMaa4VNFrDUykQjO3K7s6l39M7xzzj+YGBgmiUoQHPypPt0CLfsMIPe
CzWKYDAnhdEqoDYVY9A5CxwW8pLzCIy7nLqaxMwbPaiOy35bqsxHZSQ84bcDE3BFFChaxtGMO4YD
KAl/SwLEKwn1fzPwMbnybAIWKWRsBkXuobB+Ef61VdUs0eTcRk2VXp7wIpgpBDcFqCGNVDrkdEcI
jj86CkFXV99Yids+rAlMGghd/16Jj1J73SQRXchG6YVKesukiJav7ih3Q750ll3U/InK4LtFPs0b
TA5nGx4BZ4Rv7kQDswE7oXPEoYFxbQZCu2+n7DOipcp2+nDkLHa0I5em3vMc7Fn1l++eZAaU3oO4
kQWbREzYJdFUUDfwdzoQ90oz3D9hNfqUc2SRom1bo+ue/dpYdgHvKdjpqHstM6MOMuCpB3dJGMKA
8AbcGN/eBhlLPUNC9udwD9YBK8cbT1yjSxsyesJCpr928cjDWiUQsr1yWXh30EOpkGRKwzVSU7bs
xHS1xL62lvfMCcscDUu2zFTb5vMnkKxhXu29H1hE/0deqkQ86tw09vkLts8wLojxLqEmntKQyZHo
tjDcIf7UlZw1plH5YMwnu1gyDjJS6TZ6Yj5vVFkUQND02oHJp9iU/691iuUihkym3o73/IqWEywV
7DWQxj3xbxLFtkjkfB/mPJ70XQGVTKYy9YYmaWnmii1rMCgqK9udl2geGOkUKppouEwuauPd0dIV
km9YVD0Q+azxwGUpbPVSZTPyqQJXLN8fNRaZERnY6+5NieS+uX7YBbiFpPnbgW80mGXEFhObzQx/
2yiX7kzNrJONVHZlfJxypmi+oMPlIw1A2Bg/CSW5ptd/hnveFmLG+TSsnx0AU798sfH8PWVEbsWz
uQbFlO6+KUsQE/Sm5Q201llCuEVDB9eRLWwybGp0X81SNE06lJCh9PIyNIu4FEMqieMIDt7HcIb5
GUhcUtdDX014VxTEAPis8KD+1XwiNpcG+JdjSzrLlduchPsjOawwrI7Z2cU6ejYJN/uBensExuiX
IHyfJGHGaN2oByBtVShadXip9AwyaWy0VPfRZalQM4ceOr75CCvaAeoFc6jQqXGNKxZDl+gEszq1
cAeooHkKMBr+0HjmnTHou6I/rS0GOS1EYwohMHmB2ssY5RFH7Q/oszpQUB161GDjStReOLlb/cNN
QdGp5q6NYgJn60zSkWgj1otw8afRPQbJumtzV6xK912ekZPgvK6oIKlxATjmcLYyUzzWVPo2v8Vl
vR7kMLiY6gEEBeS/mp6qqZzS0YYr/gfcB7p2WsuzTFeQi/r6IC1kVvJzREZGst+wdHLgeztuV3uK
vrvIjinTgUQN+7GEPvE/piXf+1ZM7YXbxH1Fs7kOv068AQFLx9DBp6RCmI92FvA6xeDZ27F4ZtuU
WAXCEiRCPFS9Ec5UyF/YqPwIGNjhhgMJXkuQdjzthzYk7nXm/wG1dTloIo3R9eWILEA0jO2+d5mv
55QO/PnnArFgSRavHIuu/xJV0EWmFNWgoupyXUYJb6sQc4Ye7ZSFGGq98B5/BpFblsqgEitG1IU4
IdqS2OhUecXt4cSyrY0Of4IpJN8Q4FsJqfcaHIe9+6YIznJzYDe/mlxtUadWMCfChVLEQJm8NwJH
6PUuRufwn4i6m/9KNQTGUX0c6TSvDI0K2tiDWbsuzqKwsSwPEPc1FYDWB41YvDJYQjGX2cxoxeIW
xnMUfEQJUZfFwX8DaaZP26HYbsBPBTpNnyeQbVw27Vhmmz94V8Rn/XY86gXZv67mgAy6dwtggsci
WHHf+CADtWSVOaCidNa6bRL0iI9fRymlurHVdoXhTaReX+b6z1fxIfPbQsr/ZnWBmGJXizgbgwGa
D22R8ycSqQ653TMXTsFHg2yUKGWrcJMFDmX+wSccmBBe4cY3846I8JaFLaOrTjQ9DimJLt7O3x9W
3X/TTcLF4QQtVGFsWNZE3fWWAINIuH/LLhYKYB0cBGvOW9FnillCeLkFUlTvuxcnj/7LXJd5Q3AC
92JpyxEOoogmgLyPn+DPFMSLHHEHi+jnML3k2CebO8ae0YSdowULM+0L5+0omkirwTNJ+aa6bAA5
HH1Ry89m9pTxUWqn7kWlKy73qSsFvVzrcnGBFJfAm9PtCCpYKNa34B4RO66jz4tz325rPbB0a/dA
xWhB3g9FUs/I1ru4oc/FalJl21hfJ9OuxOdOXYxa02J3L6CTAl36BxPVZWCuQaSpKn3uMQKepRhj
9RIWw0t7dttWi+XK+pe1zgDD+I8vlG9QpMM4Mj3YbBCsWbUJuY5hcT9pVrvuoiR/7yIXRimzEjoi
W73Mk/wamC0t8oYNQkOQHDXG/Ej1ZXZA5EuryDLCKIXwfb7VaM1+P1PfoW0p0i61Ic9zbDFRoQWX
3BZWbcjkzqati9WIVs/1O+3GQDa2ROOiTUgDj5XiRBS/pEQHS4RGOttEyBuOSDSnuNS6ebqcAw/Z
6b8hriZxAg+RCVOXwc+i5loxPNdiJgKC2Dve8x/t5VJAbKDRNSaLjkAR9ql9rsnNiEtTcxoNWwqN
3sBPB8VcNsC1KWHWN08UmPqZX4Idpm3GQrwRMFTa1fk1TpVyOG6qelhfI27oFA59BDEwkX4xs0ue
mkaqsVJw6zMx752Hq+m2bP4ZBLWLaXMvW2drn4y23y/6nXa7zG91XiPctwLqZA99inC0PO46XXlL
wyNllMT3urgl8Rjmh6ouZp87HweDOhWosyo4h1j7xzh2KntmlH1dtAXiXPANa8rOwB7JwFfw1Fmt
w4IGjiwmcZAJJoCCs3Cxw5D7Ip6virJ5oDoP/M3tOLOnGFyks6dAIc2ZRnwgz1IOS1lSTPe5xSeZ
08tQg+y0chI19Z7QeyfWv/FYX7EVNznybwvSY3fbvLkgsIyeIZ/OPdcQpZxhOLuGrUuQPdUdIxg8
GAAp2S99CbHj0KhLKvLpLBrzsJOI+PKPnvNk27JNEa+SYa/2QEhAP1ixMs4iCIxjwYuyzh/ThI6W
F6dl1t4e4fyeWTnCRLQvlg4PhzdmvYsgvwyvX+fg27S6A47eXoVsPU1dqfc9perjpAeVs9Sk8gll
OerQva5mO4w16K2hZbxf9xWoQwBvN0SFdibroGLfNgF1KSZeiMaLPrlFef93NV989KBGoPdNC360
Fmb5aeA0/kY312rlFchO0wdrwax746IA3DvK1n7sohO5JAUVJ0oo7uJ76j/rQm0qshDgib0/F4re
rnkxzpLnUozLeAgiPaj6+EZxI5qT4YUfVy3/jt8SsDSDjfR+LlVBiUAtfYkPaxIwYAnMEjbOx2Xm
iNQMfSKE5VEZkcIvxPtRt5fjtveVDe87UKn/0hfSGGFPdLZH98Xq4w8k2UzGozEHMC7Vzbnp06DQ
Ccz+dBSPvKa/3/DgSSlKZ577r3OvO2xgH/55R+4Dr/9eGt0i7rk7PeLPLjS2tL5BtlD5LCbQmRI2
dXDN7krt1GbJBek3Q3H/+51mt1DFSLHW0AMEE0eY4aVrw+WxgWowShu5M33z5cRs/dYtHYf6iytL
fdcHZwSC6j798tZAqnesHPYACpDH98Pxetsbif7XNIUEIr/t2UQ+FbYQUlblWNYvwQsuDUL2rNlF
X0fCbfrxhBj7d7n34SyDzzQVfPPP2VBVaDmJvRqyywLXO/t1eAWLBWc1eXDKLOuhe90/Z8IhB41y
Jr19M4KtNS9Jzp5fVqxrqAAKickU8yJVyZFxA1K1OG95VvyFUctv0cPZDAO/NtSjTGV9G6+Ag8Od
oYayzZBtvp8D0m6FuxSx/bpyvGpjUfHd54gz2TMp9uv6C55gI5x+lE0Rn7EU6/UsoUNwqyFrETPI
m6W5U39lCzXxkZxCFUQivakeQ3S8UsphiFSQt0hNnHJNe2uCX8VXXryEZxV+XtfyjXdhxZnUcOw4
/yBqKOJWjK5+g2BoSQx/sVOx9Qlnf4UHChLOHLaMuqhTraum8pEYq+5/Pl3VbpoIxLGi7Y0ww+qv
3jBXDS5iw6c76Jjyz9q8zwEl+7Eeu0qh/lmimyJEGAVREf5qR7LOdx1xxs+oZFHJlJU71anZDwAs
p9EyAwZ7gNXbBvDeebJgWlK22nKOEvQxej0pLRsj+q4EqJPyUNAZObaAlXULSAppo3ufEgNRvoVC
dhZA1TMIDmFolkHiQ8fm80oaVzQmNbO5RQCprvwOpWV6DYBwOjrKdNCpxCecZ2qvRFnb8B5nfr9y
SraML5cDCaI8x0b0HlqiUFz/wirvAJ9TruiZ8KxVf7XQx4Jv8pXZYSAPRyzl29E7RNUX1GLnxzws
g/CTAQNI2Z/YeTq//MqVn/O46a4bISNAyPSwtkD6cjqG1zwv5+O6IZfDuL0cRPZeS0ctGBhVzPFF
CSSPmdFyuBTixBIXv7zwmPuMG62A6/7oesjuR4gAeCN4/FCybR54uFITlCFPGobH1MO/Cx/Rq8We
F3A1eGnu5slKXyC7BdsZA5cu/htpthQtbn9NUflIToGn7qgmc+8yQM0S/PcDxufy3N7jGn2IKS5j
BRO8yW0BmMkeaAVibmJAOPOBJwD0HGWWgkMk6ay9AZgxDcoLOzmLxGWJfwcsV2a6EXeV3QpFlJke
2DcaGnVoCwV/Ka5kNTfvDBIwWH5Z9yEcKs30KvkIsZI4LXSKQZDTdz43Xl5pKTEk8aRB0mVpILf6
HSkzLCGx6TOx9W6iNrxJdhnM6i3my97C8jxliHFIaBoPa3j1Dd6z1rM439hhQwk4RVHNR6Qn9I8+
BHzt0OPgW7FMmvUuuww5JOS7gdLcyZd+I2pDB1ZZfsWVPlqE6yLBg4odnvqLv+8gKFXv2a3uApi0
wsCDtJ5JzpDXatS94AcnqCfGViSYz3lc0CUz841un83P+RvV1YKzKw+OR+iEsROIBS2k6a2jM5rz
T5LkrXotbQKBPl3Of/a8MSpsqiE3nsByiJWlDsXh38X/2N8EecS70cKired2ZnobGviaGnEaB+tn
Fu5aVRQxRJoKbyV4fd2dcYpY1C++eymVFzuQ2LRXUZRGpKBRujdFDz5G+kYx18wI7bBtIRdWrHLq
rI+OKHo96xiZ37SrKLIL8GY4N4duMMiIcmPe1dqt7AAFk8+c4nrv1QwrJc2C9qFNryvyJVzrx/07
JeSBx/2wYWzhc1CtLStMVZxqUV+yZvEpVLBfKmZvOGoSqhEi7RrwqLsFwqJ3ntgBM1ON0JNMueE8
YJYIj75O/YtkgVKlffeNTV/JynCvjjcoOEfSRr6wqilPJ2mfaAFMldlepsAbGY7cKCfM650iPLgE
TnYhhM2FnoISFo0O/+fyKpmIVr5jAizHr3dKXtAIaVPr250QOEt0LyL/MZUXVZo/DMDNuAwQq9K/
wggGXQRnQKv0R1Qi8C8nhIl18bKp52wNPzTXZVBSDk1h7RtxQXFGjLFR1hWljZejzpkEyXANoLgw
pL88AfrQRAb3U2iMZKgwW2aczJHE/GUB6sjZnoVxqk6N7fxZWeLp2hQUittzplf3mcK43BYev07J
EYN6zb2atzQYgH8hgxK6eRJwTx5W+CKBtgJQSaskS7VDpe0+vkjDoCFV4sskr3LWtbX3sQEHRg0J
HOxE7M6U7Yta6qL9ydYWHB1kQMpS+7Hz2rjF59aDTN1Ip5+jxJPCjV7b+mBIwWndiK719lJOQSSn
ha7lZp7+lCHYApR/Eil6GmEPCbVaITO/kbTzyhhtqgOaOCUBJKrBs60aOqIDaT++t9ymAWvwAwO3
W4buXNt3AOYkQFi+8WKy9JVQGXfWAmcSQTfY3TYE3P6ZXc1kfsorLzQE7lqa0XV60uSBvQ2ZHe+5
VJLDWjhYiMWKldSihVepg0qv66UAFDfLLWzVZjG7kZIeXdyI2wVU8xuR4VuXtXV+Ky0PgDj/nvAP
7jPRKVSPibGTs/Hbx8bCQqDyXz6Hgwa1LxSBdszRvFW5GMl8OhlFd4OS8zn8QZNZW/VbG5w7nFfy
oyPwwTfTdG3E+pSyKXPBn5u83F4Q4/KBoEHzXSZNU+IlC5lrNi8RjZFPhxxeJs3qgKZUDgafZ9h6
HB4zv0q82Kwuf8BoTLwbrABRbx+irZLUvhzRWrNWWkuTJINWXOp4o9xrdGTmn4+3yoUBHWNrpgxw
zeD8b5AL7EPPgOLddXwXyx+Jvj1z8Hp1JyC9XONEB5d7YCQqonZozqMUEYlxbyZtEdaTuzVERe/P
aA8CG3phKiAkhm2yQYKJuircAZjHiuN/mORaLCwBLFK1ooTmQQ4mf7XyMZs3mNdBZ68UD5A5011w
BRDm8aTtQ106YZ6ueulm1NWxaf+SD6AIe3XWHSooJipikDpzPTF6NS7naXmZizTMCE3/mpdyA2qn
MVY3RKuGBgVw0DOate3JAq0mf8PwIBnja3BpFkWPaP0cnff7LOmhONZdc5NU07aPlcT5FjT3jUcU
Cc1vBBwfN8Fl8SwbZ91ECTNQX7IaVTq1t4YUswsBwzCP/kpSNs8lb60F1t8qTX/yXMKc2REz9gsj
NJVAEDXsVCclvrTP4ILBMxkeNNXc4u9WQUO9xjuVdhUnrLXLVArFiZ6uGEsG/Ytj69FGyxmWJwXI
5vKqaU1lCxKpoUCZWNYvZyBeGpWFVpPBSGEvDYUlcpOZpjwKyqfWGl7otzrjZ0ku+t7QcvoshoJv
qqJHgONoimjnHqx+Xu3O8LXF+1ea8KFm1NguWaNNqEl7DiXQ2yUs2fgJVjf4zLxzgRnB4ZapXZ6H
CK9kVV4LceDLLmQ3X9574JDFYsuAkRNG8rfRtCVCFd2C4OtlDfRACu24As1zyiYdDi+o41MeGDb2
gRQwGe0iigSweiybFPOAIPZZIrBCXPL5KvpaaUzg7PaohJCP89e0nRxG1Ll05rI6MINctvIlxVl4
NzbgeY+Im0du2wuXhO+fab7EFQgUdYQwxqtXYQMxNANvHh/OFEpLRvUBk8YMJCoYVHCPAnklLRbU
dCW5E7XpvIromv6SPTZjIHsM9b+coyVeiYL/BTJ7TvPxW9nIug/Py2ENePa87MIRLnkKBDpqeBdD
DI9pmcMOVGv8E6o3FBiTSSzDriQyhdZjcfEnQMBMFYoiucRAqfQXjzgmsvYxVm8Uv/PIXj59LpzV
gWhy8+2yG0T/j+OISVIZBwcarvEDrdneLDzgFwS080sUXiEjyZS9pPd3TgO8gf4wJSQr4QlyfEHn
6b3JdK6Yop+usi2+cF7laijd0yuRAanXBM9ygspetcrVGlcKmoCQe50N3r/eJgxs/+4D4Te5mUGR
QoNqVs4hqdGVTDU5u3TmTJ51xLH2l9KybnSGHEVX8atpN5huGq4hLAWkOS33WfUzW4yTZlestVdA
rvtzco8N1HUM9KZO+LlxAPYSKD8htLwTuzy2347sPXnjiRhKaZZyJ4lioMvDrMoTVebfvF6WzAQz
oJ1RWJ/vyY3rTEOkgfm21Ri4OfY6Ebz1zezTmYe/tqckFpK3p9HdyMn97pl5Mwy7PoEqkdeSMta2
efQBU50XSkrtm+PO23UlyKoD0mTF06kVPDx99mp2X48W09aI7WYDZIDl2ud9jHe1Q5Dt4eI8juVH
STB2z11VC1z9iXhwEIMvRZSq1w56PfnLgMFh2MrtPk6iiWAhb18WozE0PV6oOw6Fsweu6WstxZ1Z
/CXGzAthyhFySgJgkuuEoOcH5Yk654qC4L3gAl4DY7qegRX2ZiOIaqLzYOdjg0FFcYEWuqCLQsuu
ROZ+Zj11bjcVNine4X+wNT/8lOmuHY6AUKbcpML1e/os/5AeZnBjM1J/qV5rQO4xlleMQqTnJVLk
G7Iw8j+vr6IqvReR+aEBcnR4Pdk9xPRtOroON7vVY8Eg6EvsT5SM6u+4RPuXYUL02dDZ6WBtE9uz
t3BiwdQsTI3WFHhFZhQ4PKV/+mWSihg/V/+1hb0IzO73Pea0jHctsdP4li8d7LzCVUdeOG+6bJbG
gxA47e+xwkix2pJ7T49AoZG08Gh86WGQCQMj9yPl/kTcldwtshXGC1uRhz9xNsspgXOj5FA+wJbE
aKiaNMuEC5r40cqgQH5g2wz7pJ6P3T0z4qDLfC1znE8DF4wIc01cLrPMiNn3ju4h1IC/MSBXvZTD
a9pX6M1r2ov7GrfCt4ae0chJ1j2FxqjwK+ecoZa/YlhqDs2EAeufJv3jwS/A4orsbT0UJENLdA3C
0yz7bc5qgWes4MtWSGqMTyXFAPmfgNACxj9kPKMD6/3EhzVStKCuke+TOi4NbV71iw2r1bWetkoV
kgkjNcTVdhYuDBdB+40Q7RJZ5jYdvOe1+JHy/7DBq993PqPYOOGmz4lnaLJoAwEhgnWm4o2t67l3
uEcaXr4p/gVOxfHZSXMvzRlrcuC8tBeBb/wsYxgvSzejy0NHiB9XY6H0BkoCuJcpz56gyOKJBBxH
K5CwYJr3WxsVvrnsf7on0O7hsG3ofIDuHWN/gGugVwyovBQgXnhbqBuQFy2g6Usaww9b+BOUoSdS
gTYRQsP71Zyk6myvoaJSrsr+KdHz8bx5evvoEc/3xmBlbhQGgVX3Tgkc4zn79kghcYSS0yzjjSsv
Xyz69eNmBBEcS46NkWWrREeVFarNnSwVSaUnGdEEOpQidNoXlKC54iV8gL0unjM9g3L4nhVhwctE
kzkbvXHzISJOrokD/CdYOtpwjxU1rDot9TF9Y8fGq7Mv3VsnSSSczK9DwLpQ4CpnE8ikIbAOAo0e
7e8fkK8tfq1by9dzShV/t6r3WLKFD0fYwb0Ovh2vX2c/Y8KxP8E3HBQt/EMXUsdrvxYgMuDDiW2u
LC5oHYl3K3012evQBLqcuc1Z3DvMl6L4UaEsSztqeNKvibwCh7w4E5DaEoZcs2Y7RgrQgwulS5bM
PbO5TbNKU3bSf7NCTkAz62YzHlUS4uAYuintHCwiC6w2AzUjRoCiciz4fNS8tHGtlrUQR1ahjvjE
apoMTIER/30LWBM2XxZLTWyT/DMxhM8uoIMooyrXBrbqPm+5F26jvFZ77Q2XnXQrIUqmx+4CtSvy
X8uQPxCYexbttDvRgrL0ReNw9r3OYNon11vOj4oYng+ale6QCfWDAH3AGjJDIm+5qWYDO8b1XrdJ
UjtW4VF1Jhorwv7lCY8kO8LIxbT0SRfJk10YjOjFWqXvHtx6x6IQXsy0q9pvY3euKqsxqy3LCyXr
Esabz+cRTD35YZOSivCBEaPVGFzweRe39IE2GrcelO2+72ehi9mTNJpMPrXDOc6b/2aYx13NW9NC
JsbSimg9hbjDszWBO15dqv/qUI+rU7RVZ0eoEJUcs3BMvHqVny9q77c4lm0i8hQ0P+ianZ8h8nnm
zDfmHGlaqGsA/zn8QZSlRu2Xpq87CXuOIPOFRgzHXjN6TAr3I6/DJ/vJMJpaV1kQmbqNdn4YcpMN
w1XGx6KGCNWYxCcjjivTWhjjQ0XmWAXrQirng3lN4vuBHOm6kcCmTkBF1aFjHLII8LNz7KjXFQTx
YcctF2bV37alTsNRoTKPeG/X37fVkTl4NStRosEyJ7qOFJ+XjBWA/nT5s4kCEoKMEmRqwab8uk0x
IjgcrdYq5UX1kvPCCoddVL2Yjg33aeA3q6K/YcMW6b5DeHCRPkBrDf7v1IVwr9nehCrT0GPGVmSU
CqqoR+4nc853Zn7doKESnDM8Wl8DBCq89IwwobJmp+ub1O9dydPCRSCTO+c5xp+7ZH/0wUQbExIt
xn9vm2+/rguDNoro7jHEeak1/Ntkc66eAxXdagcarxELgS5MyfjWFamQ8k2ZJ2eZpxdqMupWpkuJ
DMurSepLuNpChXC3yQyLMfWSbBsFDLAyZCYvhpZwe52093vCcMKtlVNn2H4pem4gQvJseEzFr7Eu
tDBd1LqeZxwSs0x7uJ7Hr0pZAR2JfDCjOLBYgPgcLGRCnTC5n3AB1PDJ8cM3EOl9FO36Evc4Wvfr
5lS9KHYhGxuxdZlCcZ/lJSH9Ih7hOZ5WPECoUW2aGtd8wbKfvdS/jNHQQv/gCZf6734YIr2/dtwM
jPU7sX76BFt4hWi0mMSTz2bFKgZUoZQ/nzmrai25i0sILuMLg9vXK/+UFK6mpATDBxTSUwdjqWOe
bPHN6qb7Op4ybT6U1o+wuSwLVei3VLOYoukjFSRviTLNqxhpjm6C2xxqDm+UqUUG4ymhFfYirfYR
p+o/G/WifbMGIbFmmHeyOj0s7brvehszo/Fwwe9O55zV99DeO1ohNIndsn6bXJXpvF1zfr5ysHm6
IFRJQ9/C08rUcUY+m+VfLBShvGSorndzdxS0C6qI3RM3kjVcOLyLQ4MmN6w03QhLvOQs/YpXlvUa
VA2KLt/QZE36cJUyilaFRj6SGVEZkYVBvMLMXlmcwjhLu+ikdpNeUDxL/19HDdWs/fx5/MMqnbKc
Gyifh3ivilxYWavfwXCXu2V3+ovlEltVt3+MCGHZIuIoTF8iYZvkzMoVmG94pc48buqRonSwtfp+
W5OC+6piZSfNjvSSB/iz9KAtbSDNCjZRml4UcpwTOJLuD6CmGe2WpfKL5Ss8OPy5hyJN2bj6416P
8DW7ZX9j6U+rVW9cpBll1KrqLQ/DJIR4ea4i9RsRpN+6AEkuMuqVo/iti6t4UL4PzY2bqsYtAsw2
qkbFhWj/Ej39eYj8g/tlyZLcTRgwb07izxNaHzejb1PyeiXWSl6k/JVuZaJeuxyzr8I2xwU5BJpO
GNE6iblmJgQYPuqA42/NPfQRWb88/jcIJ2gXrFGl8yoY5gX4zK26ykbodT3tnbgvTvyPh8/3mmKf
xhl7PtTQQvZtLHQ+KqdAg4BiQwUwgpSfxUSMinbvEvECV1vVWcY4GfLUdpRwZIroOF9vwA7zM2iM
/eyy6Yc/J0ZFSSQI4XfREQ67jhrr5lb/U4aY4UFW+aU2JyNBpD+DZqzJ16H50dCQvwmQQkrE0Cvn
XpIqX9pXVfpm4uUtwuXOvItVz0vhJmrhrNRmrIamCiGgDbmT5rR85r0bF9x+ns4xECBcSnmm8U5k
39T43kucfiLh0J1XHg4KQIoAFVkXKYz/X+ifTqvxbaH79ZsmP62PEbtLGmMRGp7GhEfd/VcObNPR
9DsoakQq5F2VfjjdH/d9TmxmnBR4BCZy2waGPFXsMaSsuHl1j7WwSo8DwdZ4bvNnimVhODOs9GJQ
8IYGASrL3pdZgPQfvvbk6/ce8SU+H8CMdQX2IRA8XOqCUfmYQSd+TYz/FnObQ06ZY1P4qUtzR55u
rEni7TIqqpyBCuhdM07VpMjpLBfUo3cKC6kB2s+FCsVnndKjeaRPxNUai5rhqsIKFsv3HQmfpthN
K9ojA5urRuECnBJ5CGKINBScnWOFsSDDnTFBkf5cWlKHumb2+sbFYrwsjWMU32BY+eA397vi9TmP
GUN9a1HQVU/IQvt0jeiJlG+Cttqb5YkHGVwD+TOtqR9hgsKcy6JVuWjnELTfmjrAlZtkK9U6hr9h
DWA7YIdQuKWQSyRq3b/afAV19SvFb6dYbZXV5QCGbK92P9xM25Hqzm5j561EthpjWCy2X8jDUsql
XSdHfPLDxYl55xMIGLqJ5aebkjeM7M37TmbyyK2EfnJStuHMBv+p6AThFb4vvxe61Ck3R2EP1Qtz
TzUKmx+yCFjnu5lZ97jjPX1k8rByzOlwz87ijGdwytUqkqU/vCCy7B39ECLVCcnxmDnU33nwaZuj
68DqIsBt6MACT2iNk9jKWNVEEdoU76Td0ggjfhbmd9L8YA43K7sqw5FPoe4tpN2z/E+dJY7hAppD
rVR4vjlFaxQax63YwOZD1YHQgkdicuIh4IXkyJSvuk2l8bbe/oUzQFB7ZmSuoj7ldC2a29Z8mfEm
E9xav2Su+qr2SctJiWofQJezdy2M4ijkm0zlZ5YopoKnzdaHwpeoIgjRHgRRQmSZxEoHvTJXv1El
eT/NZRONO/P7N2Oae9gamA5a3g1P1RBuA0GK7+ozFFkWtHOVMU+BRm22XfdniM1hHU/getlGSybv
C9ucZmA8XVTHSoqYEE5IPhDE7/pUhBjhJOKn8Usi/jZNjBMkGeB41WIBiHl9CJFjK2zj8EE03EAm
eMt7StCuLlIc7ffKJIGv75+eCTFDjDYR3qlZkeT9EPZ73aqlVp308QXv0WuYapzMD0nL4xyHIyPw
uNTuIibVKX376sC71oGkS7sYzxyFQAowHGga5IDXrIWgyVEXEj2eDqhQ/b2vsfPyzYcqgo3QLOeO
PlKx+LzVq63QFKoBe9dPOFdv6l0ryQ4A27nrJBfZXkJ+LGM+QwNvS9pbVysRASIY6tivfYeKQPse
76og1VGpVMO7CCQFnqSdUAOu1Rj8CrDa9wv3x3AIMSSGmAToI+v0jypcjPA6YR+wkSjf0i4A5Duo
gdu+sxmgsSenZcYbdSpXUr04SowJRCOgWMQYE9MnGrnyvukJGpAJD14ypYw6IsRLZW/hAG0v0Fa3
qI3GqktKqi0T2feKTA5Q3XtcIizlsLhOiV3knDI5eBWvZ4gf8k4V8M52Hob0eGk1jhEV0M05yGUM
CXL/7Ea4CbOMgI4Yo2jzpM7++D1dvBvVU9vPERLnn1WO0J1mjmBcS1BhVdQJIPKV95Jp45FO0SdL
ecfkPwHtO3UMUrqsKO0RQ8ie0Te/rqkg40NbXjFhFkCfX2Szn+hVg1IQM29vtLpfeikNhtIaPbBJ
59LkX6o15bVsA6IhX/Gl4Ir8jn73eaArLG1t1oyjCsZJyanNevLDWCr9IUfLoJ+De7efO7jHoF0V
bzmJDPL9CmCKvxaZS+K44yyt9gArBFXCRJ1ez5ryPSUeNxmmB9ibzn5XucdC2dGyCJcqqvrPT8to
vWFsgu5zRFwEvpn0myUAI2OTYxeIU3+lxuauCdGNUyxAParrZK8tstWMxpxD/HZEPCDSU9Pvz+UA
IwgRbsTYJBSHOynp4+Ed/Q3vzdaKOSMQz9yKIrXADc1aURIsnCCoS7EwcbxzP0XkouGQeR8iGp+i
Jt7t5v9XFNQdXyyjJfRHZ8OikaRM5cvs7vMLBXQU35MJVzDqEWEaeXk7HVUAg8S3qYpAqgpLWts8
Ub9SQE9Mnn3gJd0HKqi3C0tswLuvkWa59jWfeQRV/vX95qmfBLiJYM5JyN+ssB2Q0KEc4Dni3Nlu
e0qs3TZVva2W8oPUSl5jiweU10HcN+nkMvzokotShyttDINCB/Z2WG93olD8vIDXfTBQw4qO6AB9
G1sSS1FkaBO1sb7jFrlf9sq6H2G/XMQageUR+bjXKnWz1JjcqPM8WgKVd3sLVZRc6YDQpbewIp42
gqdO25SmzBi4L9YVdsldFzflLRGcH2PdED1/ZG1sgfPc/lzH1c1mXiMwiYy9IY1tzJFPcG3LyWDo
IWfa0lj+BBdbfO+DW6vY8ifOKvAKQHAZHe/I0V8qxktUVo/B/SY6Q0PmwmUzyU/3oaW1A+785vlW
+mbFaK67Nzai+n7iuXxy6/fyPHEl/DbHVXXGfMgNln8uSz39weWxH/rOLUHp49++Gi54gPX5tL/O
UdTmMoEsvlikSS8lF1sVddBC62JwbCJq1jUzhuIMEvu4jJ8+HI174/rYrZM40URwh04l3hHlQlSz
7sLT2ngA+/lJcbEScVzq2KNAOM7hlTE6EKIv8KTc19+u5d5lzbaVQ3bM4j/Uvo/dY1mEOtNbA97E
/yk8fMu8QiZVdqf9lF8sy00/xf6UfstifSha4b76N5GKsfWMOpnmerpLwnDdiRlPZ5h8duaHf3dZ
humz4YZbGdVEUG66aaGDBnYKc9Tt6WVcXJU9xYGxrVTX0bDUNu7CtVbDx/vTuXPa36fg/Vg61tc7
7WZChnXHb00g5bCTehzFZ4vynRTFGRt4qR6w/k9htRPzKk2Bt8i5RJMUsbqJW3qmv8GdhEUQT/No
KYfQjKQMrFIbcncA7g3JQP2Qki1yh+5stpu7kTuX/78JWBLkotmAoConO9KLxdIUyBfQrb/RhTut
VjsP6uNkING5AM0hFlXhfZjF/TfTXQgMEwilcXKdujKcyxYTqbmROb6bjSGeU3hHlrfHSYR18BXA
c84VgvE3n67VHP6QuAwtkhJ84AGklAC74s+Iwb+olKxRKpkioy5Fu1tctEZU9uQB45gJ94KR+nHU
frxJMurHGr0IyIezC7DamaN4h2wWGcosGODEp06vo9SJ6HEqx4xGeE/mHwL/vstimgxZw6GaxJXW
N9adPFfMMcTNp63KmhHT/g6BAyA4UrtAGBiU44PiVref0kdnaNfbpCZRZYmnPaKD9zcFE3y0bHDy
Q6Br5z13rgZ89EVC9s1Cs/Zdyqv7mV6znX4YVW71mLmW8ZR9vEWVviZclA+hQEomD1UUruA7S0fL
9tyPwiZuPBG9u3YH1WifUCRKbZcEtyw+IExzf+5e0Vx7vznec5aqcqQGK1DuYlk0tKn4f6zmN8dL
khXAqhigC7wkCPomIVG+MaLt/bFjMEedWesfIIPVdYj6ZidKpb7Zo71CtApUcXYq6+CJEpubE7AU
H2KaSjHeS3Yd2pt9xWZq6fg7386Y/SHds7DeUTINRtXgWhtcoysUKXUPkBxb47G1nUURJNBDN7sX
HyKv4W8u+DPjAuzqoGCdpUFuUSaTc2dDbeOdnnvt1Rf84J8IoR9x8a2K2dElDh3/3kNrubnhPfFp
aQ9zAR6fXPRtTxQgWDMFnEXVNN5K6/r/kUopJknqj6HcGqZ8zxY5bKjFDz7OiyQ2Oynmxey25iYh
I3G6rgmw/nSR4GtEBKZ/juKYz2hCbZ+jO+oKnJcBXRUi9sNBylqDe43AP6uaobA5fl/Q3o5H2wNh
zFZS+idVh6HS//5H4HR69rTk7K/IwEdLSaUiXSBQNTkJjhckbtOeZPjMTnw7MFIiUokL46kYQgZB
rvYa0O+hJTG/Y4VZEWCaDGyIcsYKpV/kvMOH+1DNhCHpRyLHm29a/pXV07rVG/6RvR03bmsYB2iL
38duFls2EcXQnxq/dz9fmFMxfc49PljvM9xgwJb7JKTA+FTAxi9JK3wvbxhgLdQlcOLjNc08Ca3j
9zLzeVKPZczAkPqOkecQ0mPk2VJk2TVNy98/YKWA9yCBZBpPxr6b5JeZPsPBgKz2DHAW036yCldR
ILl5D7JQmSFOZkLgee/N2uOCbIzL64sE6d1Jc2x6NCbB+m2VKZug7pWqE3cy2ONcSwbUlg/5SzIP
MJ9gVENINRnezsRVxtOBGvuLHFiPwFMJr+21pCir/0LEA7y46yDRK3JikPTipPAB87a9W6OHF5vP
5VKq3UUUlcNLGUXJpd1/Z2MY1Jcocq4xrLuJKKqe4H13leG054lG6PP5K/gdEtNe+1hlVWhzwBVF
fEe7DIuzUOmht9Y+dY35rYTEkn+/bbHjts/tq2m+TFxILwuZiVqtlyNyunPIxVfjjM4a1BzeRGZa
OjK0p27ECh50syu6haVHtkkX4PwWm6D1iDzKcjUPG3i0GXQ3ly4cVzoPuzcf9aEKUoKEiEL7f8et
itiOrIrgyk+swC3BGZ3HFff3N+qG+A1nJBAxZ2hlvEEwueqGa2WeVVDM5O2BSIvSu51ac+1/gY3n
j496W4t6wt8OqbZTjMGYulvwzCrsKRuW523yWkVpyAPom6wytxdeWlfLpf2AYDJ0FeZIUCyDu4g1
JRSx0wWHJFFFSRArysEH6z9y0GB7UQqCpS2cjivMpfoQbbfMQ1hjCm13jvrvnKsNw9fG3bgoltGR
+9EZoVyRF8FWnoHUbUaQ7EJK8/0qkmz3xfzjAq92ZzlFu6Pe+UzRLUdnOab+BJj4uDWe16UC4c6+
yLcGTUjx1jcrs+wlJNaKqY+z/RmIuCqg8jI0ZjeHtqq+mF/lJEeKvmHLmvue5fwm+ufC42PhspJA
2TwhqcJCy1yAB9ptMtxJaGLHX3zjNdrasIef2Rt900Y883MPPoPAYJ1VVOwS5sSPd/B5oiOjc4Sh
JBghm1lh9zRPtD7Km0ummhSOsxa+tj9uj5xaICXMXeSJnmX8Ro4oBEwMf2ATyY3VWCld+HIucRos
XEDCcZY2LY31gumKwUHoxe4KuJjOcYwEHNZwIfsK7WITjw7FYNEzryK98JYcEa0LPDU37pemGBpi
vJ8Kd5FjMMQbdJANVT6jbHSfji2c5GwSmR27fFFl8AlRMTmvFssDFu6adZRJoiwMrPSffZRGEWq/
iT9jX/pxkjegy4KwcpN5bFDDuaKlzHw03ltg8qNP0sDqWWqJ/J6Z/IZ+G00YV09NXL8ILjd9ZkQC
FRnBcXljGOHjGYSUuUgMCePHip0QCa4eIo/U19cARd1Lin57LCKXZgt7mo3F7HjPHgYDuWxDdHWg
kwoJGm0/+IuBiOvgXivf16Qc7jZ2OyxddveyMzQAf+i4YrVr5pAqRfpHH76ND/g0SbeHXBFBUha1
lceHEkGMkk/S16uv7IcWVvvx7Ik+XE1x/LT/YT5ftm7z6Y0Pevk/JjP2gD0xZiL8hVLrBpip7JKM
FE+FeE5Xs0JLTpMlhW8mvNiH2p82MDWmrjDnaD8fyekYq00+IE3o6IQemBO2b6eJgJxCPKbYrVGB
wuMkWNxebQBuqAh1IKwPdgkeRNKST5G/fERAmM7ZbeHD9Zibrj6ljaa1w8LNQ+l+1MQ0P6FMtJTK
5qSSO8WxB+B61BEdP2mGp8SVdbolmSz8rnSR3B+H5fN4JsdNSo5bF5MLxKdwocGjMQRdY9Fu1cgt
sYqT+MXN3p6Kx5C9pCqlBYEBWejWiKG5/2vcoEQTDin68O9utpVCDtLoKh739/lAIxcL6Qj7nGhU
WrDTlPPB45J9fUkem9uvR/yeEwMp87RI/9wn5F89P7MsZntqgRgPk+7e9+SMa81SSGZhkFfpxRAc
4LXdE8qF3l02dK+Nhxi8FykfzbPM+MerMEjgotTMgeXeE6vfc1k7zdEGp5pqOmUx7tP6rdrWmkfV
GB0btEICFU0NswOOla7qCvX6eoU3wOtjp70CC43IsLbis1VT75FflfYpE6IydQ9a7DTQJGtrqNZG
w23dVgxMLj2pass1vRwot+mBFQXDd2ytUzcjO39QwHyloUX0qgcWsuUc8epAspgWeS9Sxz3GX3vd
IIwp28H92grhUxrd2Um2H8XC7Sbn2lHK01XsfjVnuDq8hQKAmnW65RRuprkLaqo/gsHXYiqAmMKg
v5J9AuFsGYDu88zOdiqFrpyB3lmc8jWpz49y0AgLrJPG3QssIV+LACXhBJBGMCJYkuXdYi73RkJ1
RqSfQCI+Nb2FJ8Iq36CZyJTInRXVZGnKckjA89E0J+iwT9MRzptnDin9DyqseT9bImxqoYEFmmdB
ujX5J0olxsiIIyJsApVrUln9IL1hcvaZtmFJD/SfsbCK1nZCR6vtesyXTBEj9XSUoDtTFqW1ACPx
RV8LuEvr5tHmg73Tw+rxgU4tvDkpDgwc1Uk0Ln5nuAFcVAttNlvSX0D4nJTB5+/wuq3YEqfthgws
25vwvfF/YaoimtgwcKV4oCdhcjrHdh+R3DXsTB65zYJbJhxU2IOJLQk1zqE/y5lL5sXTnGWhYeeq
WQxm8eboRwZHAgrrmeQH30isU3he4OYt3GPSGlcjai1kRp8LxFZ2wT4VbRYV5sI4bDb+tpfV2Kjs
UrRqZVjrmOfyfjx5ZpN4lgUdXZwuz5rQOykejxBmeCfwhzlXcnyp0VhuMyLD8/YXGByXn4D3+gAt
0bfiTRV4BNBN7kRB6x8bvASJfJfXxC41tyjLTIJL28PQ+KG+aQRkBds28qZWwW7kVmBHVN0BkJRs
WFnpGb8pGh9uvBobP/hXXE+rlAcP4HiauA4ridgimaSx3+vH/YgsCrhivYdFkozcnm5Hefqq2s4d
vKXPSh0cORZH8dP+hNWMwTtjKr0WtiLiOR5jFhjnpzkQGwIs/MBWm/5OB2xm3VaUOHEjOEiLD/YG
IxoSOLGcYrc5y9OTISfKaNZnHMK+7bFWBBnhkX+Z5xxowGAhTxgJkC8qkYMmcSsCFPdRdYnvP5E0
Oe+J2tUV5c21fMY8N221zUSHBn0M0Ei+d5znDcRFPIpCpvIhwaARBmOt/KYzE0swzXguB4sllwc0
RG2jPidTrBKCBcazCbORCCT5cCA1eUw6Uuh9z4DR+2ZayGzMA2Ov1pBkwHSJoKB5PT9RaNRgDP+j
RYtxVBuu1GtqIr/Ro2pYJmfvs6BgCOS2eNBsxEJkId7Tcjv7TiAiD/9AQM9q4ViKTa1gHEerOpYl
mHGxcKv+Oe0kniJX/ywA3z9aCp+gZ5J4EejCQ0KqHH6SQlRC7HdFGm1Sg+pY+F4fVW+eKXXYZvOt
+1SJ6KV/LCKnx2qOIgyg9SwjwcP1anYBOs8k7wis5g+zmdFhYuGaCm1vEI9Jp1du3iizXIyR5t5y
6DLEwPqr+XxZcmoL/vziavJLKF9/uSWilgj6YqxM/J0Kb7M5SUz7HubtybV8btVLsCfn4zOHxLwO
Em2vsYzAFBd9hxEY3Pz6wyscfofJgByoqHnvnd06pfEkuQhCIAP0P8E6y2N+j84loRbebmxRad3T
FTZMxmd6B4mEmlG6kbAVagksD5qJNmVjWyOr6zRqs8APyfXJ9Tru3EMSoFreeJKvz2/Fz4jYaZZl
KRhWnyVDtIY0/3MlUEk4xVzlnm1KSnyKE9WkDGRTQp5XBxIr8lDPhn0dfilJ75Obr/oYSLzu1/NC
9yTMURS/78nwOw9kh2RgpOkVFhO46akAbHq9NCHvNZFZBx4Iq2pnetRRQgNAFcfGlLcHYN4HfyQV
LV63LqDmwa2hdrxXtn8ApgT4l4WmteR3+H6M3dh/tOu4j1z7sH0IKwHChE69YcZe7g9FJq2A+a/8
niQ9eiNQCwbndH2JbBmClRXuCf4Zctam25yXRQLn47CO5Ou6xIqnxrDPQ7i0PAQa5UHulUCvBpb5
MvszXayp0pAKZ+AfpW8He6f+xCjmjFhJGEj9ikk91By+LMFZKaX2dWjSmrECVCP7/cXhWaYNJohh
35NZ07yKxqYotv/llixL3QHWYobf/eNXcK7rdSVSwFgczggtq7O1/I/yK7DW20UDXgWTWPe+h0gO
EeF/2WI6ADI3BX7RUPMjMKDZWd3pqtLNUJakohObJB/YGLbb1gCifEa3PB/1Gidsye/X2k3EPW7x
dXIvSSgFXXd2cImXNYP3ZD/Nk9Rv4uq+O7uEs8MUK2OsXFoKZ0P8wVmykBBfuhBYJFs5W6hZdk/J
pbwicyzglQTQQVngDQ2oDrlpOyRX8GQG89XL1RKinPFT2i41pRD30yBesmUtzEI/I4bDDEpAXOWR
fIyKB3qr2kSPJuOVKUpEmZtBInf8wkyZoaR69pea7Ql0ks43j2T6sZB9rgO3a1lx+srsudcEOBX4
qTptFAL3JZQ/tJ9l+7Ei9uiIojMF2Dh6O1JQXkzfIObWzP4eRlToNjm7cBlaw0wy0l1LHj0MCfzM
k2/JiMt74z82rDg9UnCVMrkC1rpSl9jcRbXOFGw/eSQUhKQSyJtC3nRN0OTyghyodVWJI/ppdz9e
Gn2f0TclbuRh/qz9m0Fy7TfMEyGyfuR+UC39k7HQMvEY39I1GPL3tgtgEFjd6sQXK65kQVB3xP9J
b1Be7sQt76yI8c4lMOgH/X3ES+2EPdymb7CQO7UHC+QENPmAILvbOPE+/4N4nyHdih+PQVhnqwMl
6RSq+PAvDSbBOs3LZQN/bT8mbFHHfmIewUrvQo2qef6nDUPxgCueGTB28HYPFglGzDHOes8CrbGX
6YlazVwHbBxpP5TipXxz6ycKDpYAO4TMl9jZogrgcQZL11bkh89fK59uHZ3a1DFEtQ8ptnEG9W8V
1wGRCkRAEeXrCSoQhcQAZHbkgrwzvTPX1X1bVeE2VLYNMsyPopeDZdaT8rWf5WuKXPOck+FvFoMS
I62z/M3DfruqXV2nZ7SnJb7ykljCApYsL9KZSbzUcdnPmXHOKSiGeuQNGezQJE2DvHFZo/7vOT6z
2GUAlc7sJWfNjmimpELnzU1206G5P6O4mHgc91fbISFG2TecrgyUBUEEG3Fqi93Xw5wvVwxh7p8J
v1kUp8VFd/ArOKCRqMKOoZA2YgGCFmZx6d7QTtQI3vsfTV0Q0Uvdxxy3HIM/453RABqv4e+7CuP6
FHMwsp8f15B/on4w4XKWA8bS5Y+vON+n8gum9ISFOc3OAnIdqdh+5+BJjRsETvqGm6BlODYXCw9w
eqeQMiOfbQzvNJ7BUoSvRed9xN0MTFi8uPe5bUTi2/hGaLak4lFUxNj8YgYs2BNKcmU0duUwQ0Yu
2dftwIit7C6d5vD9RaoweJBXIDjdVgYd9cwqtXIePjg0Obb6u0zrg7/nEt463xSlWmBQKe1hdTbB
2+xX5TN2cYyC4TicBqsdSSc4mwtgkTir6JqGM03PGhTOhc+4S/M8RiiSEyFU8VwXFYfz27RHXgp4
F2waqzvjSMCdB16Xl+Zn2Iw+92AEzFLeVcIS43o5out1lIMWbg3F3kKj4hKuBNxprrLu5eEPJ7KM
2x3u3wYf2zdAFwUPH/r5vBMkrmxc6WuUgqH73MP8wvxQnM6tpPWqGhopnROMVaJeecWW+9fRctfb
tA9v7T4uX1D4s+tTgwlyKH7aV+96hLRvmaq1OIEWN4VdMm8wrXRR5SoUkB6D077o6QIZyiWayC4K
7SjPa3f4fSn1XwF1V9xuXEZhpjWSWR3vsyLHuVtd35w7eaqJSWl63XKsDg9beSseiGD5mcIXCMaE
uc5h746akzCOxFyHPmyzUKToL663qdYMhJaW4ZbeJsTW5RzEoEEaJfDzNR5HZnbFPtTlRAOa1yI3
/4tr1Ycd0xq9mIgVTGF3CGJkNyLOPR/bYWovS2dNBnxZ8ZIrMt6WiD40QnOc64Je4eP30Sf7aYQ2
jzPLOl0xSv0HTx95+kC1DyuH3RDCOnV9ujlM6/9e3Ds1Jz3tKo334vhI6OScTVSJiSPFOPAjfGx2
BjEtG8J9tYmpbTYjXyqoaXZZKlvjEF6c6H4jUn69X/MNx7LTwUQ328yKtWSjPZ+g17ukIvu/MJq1
J3Wd0QiVMYEdFpjkRByYEED4H/oWOC1/dnzZDRBRVOsEb5oGI2bH9SPIgXG8g568HUagZMCSGqFc
aaRnfAUez72Vv2z6S03TXPzkx+bVjLvFNaxnPn/MoXfCsb/YrwF+fV9FDml/PqMEyaOlNyYpofui
5fFHAIIQnQfF+HDj0c5nVJpt7IuYnXaIFe9oqpjryU3J3Pt43iDKmph9B+1A8XktjrSxzDTyQpOS
FeC4OHzsaCRIHgfA4IZL/38TszMsG+H6qBy0nDScRaB1B0kyrL0SkL1uClXFA2FpKxQ2acpb6y3b
Fz3DUFGLcJ/tfBs/Owkp9Rls0YWDCMzZpEC7S8YxJo3eWRM5qQZQnUjs01yyEKTu/4Nq/bFL5HS3
cw4fPHnfrkAhdnZjh6J4+f2J0Pxra0ynE+TNR81Lv26lyGHRgnAk2vAMo4tkmSmZaO16d1Y7sr3i
P1FlYC+3ZPMF9AlJaXBxTgCDOM2M6XPmB0V4igm/4/uOcUDTZE9f+TlXtKP2cnQWf4V3iQxHvl+p
PllzMbUsOJkQY7YqY/gsNn3HesHUITIjMF3ebr1pZfVhEHxv0M6yy46AA33+hfiz3HsZHFIrIQb0
vmuXb+NQ3sidusrsxgLcjseK84TZ5yokrekTM1nlUP7+fLNCE9GCbcLSUIgOgOw8dkXPO7PAnzDt
mLm0uPjNAiqr65YPyDhOafVGniDwGz/aid1/jbF6OoRnKIVi6MKPV3dk2XCVlg1Jg0+AYgxY2t+x
TRKylf8xQPGJN/C6eo8abCCozIyQ+fqnlgazfxEzKO8RmUBw5zuI8H9mOq0zLVRJzeqMQYMVaG9A
MlnkHwcnpRYUO46fDbYNZwuWN+8BKHVvwhkgit+zwBnA1HfIhkhUgKUYKIVnLHWK74q9ynbjIrVh
xkyemobadr1BbJ3T76eS2yg6KV2CQDT3P85GIdAr1CosCCRr1pvJdZ2p/VUokSbbW3I5RjNU9H6U
j2/XrafjRnJ+fQMjOEPub+3jhh4UDTNdhFhaio6PHmBIjGZEA4cMQaMwTDGrWKi/miTd5n4I1YGN
FRgxTup5Xy5ulUsDMVXGMPI+nNfPENBsG8I7oH6Tn22P6kTyIc4zACb4/i99jUM+2h9PEVQAyawr
zmrAa8c5aOn7FvARuDovdX6cBkX/aLnVqfbaEsVtnr0jXAXBuH/xLoSXydXXqlLbynYkA7o9EzDB
KbYSuNlaE8m5eunSFJNU+KY403yJ6ahREkLpoexMBqkmDdHWXovNsEXz32HplY1IzJDhoimqC2rn
k/ienAih4euVrjNmRVbxQ6ElXJAG1jf5UWtfn+m+6QXQcnQDEZyu61gPT+A/N2tinJh5d5LfAV+j
kMbPE4oPuo6Q3FstdIMCC/nGM1W5+0hnd+CpsqUGjrh5J5305gF6RTy0jZeO7I2EfNhjIRp+OYWJ
3HYeXSEf4q5y1QUgrWAhOp4pMHDFHjVAJ45q9Dq9HlVzIWlsJDuvhMU2FynyhsXCFB5YtcYUh7os
RJca6GD2BW8j5R3lAw98ifcSybuq2/dm92L7++I6OA74ii5Cuz+QPxKMs94RKVlzqrjjUGj5lAwO
furnTocnoqaRvEFHRBBxNox5+HD/5RdCb1rXcE2nzAjjwnQfSzNZr1ORgnCO1phJue18paS9nlV/
4cA7m//7R7AZgz0kSMstG60fv8nST8zMg/GaWj1vC7qO4iRPjtA3116MIAcVJNkiCUy1dd//02Ub
qrSd25GH+4LKs+pKwxKlQyYLmVOHPkQp0SiWMNrUlZO1CmxenanEJgWM+t/EFaCNTL43xiZCpYBi
aeVniBT01rilJqkusuzfmc+gNUu1cEY0AIAvAQ/WRGS9sdNkO+J17HkpEySfaoCA5JBtQLdlNSGq
3U3wEd+QWdzId7SUin+aUv06eWKdcWFxV09E6AArHM5pmVYUyFsYuYoOczLmZJADq4oa4cqrpAm1
5WmOym03pTfNlTMUkvz5noTOmZfQgf1BxdfgXnXcfKOvX5C7WJUbTFFPg4CWwvxRnXiz03J3Yc97
LNu4ZePcVN2+JREcPNPpBAirTbYQIPZrtO2IRU4Fb+2V54Narsny4/fvY7cKhFVr7cOaZit228GC
o+LH4AMcwkVQbUN7uIL8h5q5T6wzwgO69akAFb0NyaxYe0mNK+4CW/zKJ86ZjMRmXP5o/OjfkoEz
tr7e856b66HD5LMzHIoqGnbgFsOe+rPzy4G+vNirbu0nkbm+1k4FRll1urmZRbfvQsdORrUekdII
0a0bktT78Al81NCfDNPsG4fh5P8xnrbu6Sed5CNZ4Vosyrz9TMjm71pWn9bWGxZDq9e6EpYsKU93
GXqT+k05fphq/ey1CLo/3Lp+sq1KshEZLDq8PftYNDUXKIzBH7/Q1dVctwJ+Y/c2o9omEyqaoYzR
MoRQV5+P0YXgCkumAdTEhP7IY5qcblWHv+WcpxMNYm8u9ekQFo30rlWAW7acWP8rbKiZc1SghYEp
BToT1i9cb3FXs1dR69obf7z+ayaQk2D94vWPMpYyUcABakur5rYMnQ7JDwcW6ST46/CWoOLaI4HJ
I4Tg9zkcGy23gYIh0apair5+oyAcQalFuhuliC5r3DNfd4V7wNbMFD5EW73GgOk52kBXdVBAFhkt
CwrnENAKxz9Y94NL5LLJu1BY43fYDsZqyV0sJwec54g6ecVkeO504rVy3JyiHv9RSkB4BV0mFqjt
nlNfT0eq+Bn07xi87Bsr6YtEzuSELVhEXz4uUqoTaT1mmZ5ILBT6eOcW+NO91ozeUJODoJUF7twK
XVAoJ+ipC4twa/7bUZvr2+uWL49SCscYXC1qSN1r4lX7FAmRmlmWQPPoZKbWSOjX2CbUfpvWsVf9
fI6MBnUn4uaurF3WUP898tsJEGcQMbbU1EXijjJ/cEu+Ge9eVrbXk3ffa/GMfMWMQBW4EzNDDf7E
zVaCuKDeoD6mSd9UCyh9EfLQKoPItCHiH6/CCTYD4kHS1LuimIvlhg1zyLYnNMLxawRwaiPsDDoA
Q0uLiaRgW72BmNVCkJgiY+MkDnxYDplFCppuO5CJ54h3HNgHSxf+3dQEun3pUxIQ94omYd71IjPL
Q1PpdidzsdMBQXWon4jj95SWlS47yaCwEsEJjZlhZYguD+x38Xd7c9sBMDk+fKDFQEwOx/B8kl7y
OLwzeho8uZbAubxJAcoeADml+Zo/QeYba0TILuOCtZZrOyTH42uaI9O7cayCV+/ZFjaOTe3AnT7v
kXDOh2he/pj/SwB3Eoe2iSmUBSachjDYAG8mGMUZkNAUrosYY/ZviI6bUQJwA3LzN43o/X9sKuGe
Ly3xhHEBcgN0rr7rj3sdXcnTpwPNv7TKbP9HPyS8IopGlcGHJnYxQCQNddp5nMFOQbb5e2jVaBi9
MI1b0vfIzUdINSm4efpl6JZjeo+2/5u/E55UY90Au5PeQITGJqlkIAeOWy4WRmJi5EQZS9oPgyUX
7EjzAlKtF9exR6h0APYsPch/zaQIMSE+0TO7TxpsBptNvx7eIRSTkvm76WBUS+5FNEmvG/HjRrkU
hm8fTO0HPQsXFacnYA1ThbV4r6EbPgMv9/oXtMSaVgl9zNDNK3ShZuy5rI+iq2bxSfNb69dFSXGw
LMaMhSGJUt0qYNWemXVoamTX3ut/BhvYxVV3I2uAYwjz/TdqR+b4sb6EWukGwabOw68/AeQp0hjo
lMbEFyLYHjHM5xCeN5Vhn15Gr9vV8wXot9D5f5PAjfEJgISADZnf6DpDKgP/5/QYfoJQ7uIPazvf
q2NDwbeSprdaY7jdksnsUn588vEhLI1YBaTGOnzFCbHlaGl96uZYecCKAODY4MqoUiY3Ui8JaL31
1TCPAURGg/eGlwHeWGHx5tBtoJD/BUS4F6kM7h/vK4y/CfnyDzCf9DiswUFeUTG1QDkR2H3wkB7P
yer9UACmsygVZlqfCkZ/fokSPPJr23w7WooVsI+iiCew1PX3sTViRUi6vUSnw8osQ9c0H2A57gHm
L762+ZXszBujt7ymKgbhCiY5uKTUTnY8S0vt4uq/5eMQNPscJ6J3f8+yC8Xgz2HlL4oIdbZuyCQv
LO8f4Z4rpxuWW5J5I3TXeoCn1Ee+xc6MV/fTLUxUGTPqw+jJ5i1KM0bzEJKI1RLCrxtS3YPJhWwL
bVJp4uPFANPN+9pMpDtlmE9XgBjualMlDIQ2lXam9XhP1PH0U793f0CCtNAcSqnLH3fpTz4VZCMg
HFFmAnG59is0aQ9OTKdmcAdLENCyBrbrz1YTZYvLqxUSUyfzUIf+otK1hyDgJo1f2ncSud3lTHQ8
Ocpy9zUN3EU3ql7fPBvwDxMfp01UCQLLnSWlAuXPHW8+FirZNpQfQTLXo2X8ooW6N7sO0sNSHGbK
Az4sUI1+HfHTFUHRfAP8+UNP933yE6UHLfqNK2KWPF4H3r5eLmdd/8lWxOxB9nQnoMMQ55/UXIY2
vupC2vyUHL4o7dVICUqxXmjlJpXdMbng+gAzCleIpEDfqoVOnF2wz/PRRLuADaHmlqItmhww5hiT
9AJuwTzcChEivpxrODVuHRI4XyK+qQKZEi7YLq1WSS0gqxQoPcmY32yFMbwZavudvE2r/feKWcuk
TFJmQ6zB6jeKNljgBbt4iHXVOeU9Wqa7SasatDM0dHsMbAaTo3/VrMiX9M9tFudeRHQgnIC/tZGO
rmiRqDo1bLNs/pxxfBJN1/JANc9/km8vAlbGn9L00i/bgn4b3NlyQjccq+Jy5kXiTwTwxyO1wnhC
khKBZrfs623syc1VufEDnOJsts2x/vk/zifsBoSyanOMQIFiQG68kSb2zWyXymQ5QDWZ5vW7ps19
Hhoc5d8eWZtiqWOA0ekZ/jdKo9lWqcjaU5ZUEfQVu0aIVWg/hq6Y42krR4QQj2sLR4OkfOhpqCaW
BtuEyGv31EFLlJyb+D+kEd+nQGZpgPkMewwvfBervFopj0yElLCL9Mtk1FZ96kbCrTqURq9T7/7q
lwRtfwTPqN7C9Jy9j0+BgnPTHJEGJhj9Z/Ki8szDKqvxfKrGTrQshz4wFVKrdFPchsLWZX7UZ6bB
iJdmV7UpUanIPDdMBDZBRp41K6HPdUcLZNmybrWtPEqFlYko/oL58Ga63QpkPzSUiXUBHpcNRK7i
UqkW5xJdOCP2ZRvaMHUttnms4wprcoo8GjeSMCWEWbHK17iy/wyZuyBaAukGQbGpNs32+XeLzuSm
ANkMy2Pr4yDjb6MlrXfTdxpajwFtux69Lxqy/cd4ICGquiA6BQ2R2VFpWbLI4ukgbw+nPDh7wqqs
u6a28hR8MPo8hMe3u0w9Cx/G45gn2MH43Lw63AIy+gCjq6dMX8ZJwnPQ5KQZJxu2rrQSkkpRE3XL
DDiNBUJ72snHba5f2U+aeaFT2DAi3woZzHcVTI7D/2va7HJQpV7A+qeSPFsbedKyjvliaGW3r4MC
L4g2Oj3sUxkYyXa6248Cddix/mnNV49wSSHcMkQAop7ZkJX0UzPzMNWBx51rDJzHauBFV7peUbLI
2C6HBa6jAbJ8ZEcGoypHb0OkTl4ri2m61O5S6d9v3LWHv1lXEyye9Rjnt9bcy7zD7Ncvx5l8XpQQ
OF8c1mL+P+bCBNfDfyrcEFq+hBiPdBWDrApsplCGsbZPs6MqdJ0jp5rCTOfFyi9LJpZRPcP4+KBN
lTYenPE8wrM9tJXwmT7IzNStfQSjTL3JgReO46v0m1rWVJg2oDJpAqcK5pBsZn3mTXpWIkz8Xnt9
MSX3wmQ+BUJc2BYmCnxEK5HshTnF5l9PQ1MOSpYM/7pJEflH/rb3Ui2/2eDE+Z9RUzo+EPAYod8x
naPpW4eMINKzOXIKRCdQHE4WRKqCRAURat+RLZyP3r0V4Rb+4xbAStb2/ZMB0MgIhLJdBgxr2SEZ
lftRPEDQ5fVLImeEaLI8tlFLMQbf8ETtwX3lIzrYA6MuQVz5Ndu6jXBd5aae0dXXGx/m36GvXe+k
NwZ/GS+So2trVTI+lz9BJ+cpZoplaUkifvCVyylc+dbXxR69Cf4AFMDbEauSXoXLHwJ7UqZoF7e/
fyKs8Tf3sJEToBvqHoAoCsD5uA0/VH9t37v7QhyIq7L5s9faMU10ihXoY6N6xcbwBDcQh2/xGG16
1yjN+qxL9V0BV+lBG6ltzdFbQ3nDQnzdy6PVpemhHGbNW2Ga/3HLU3bkXYC1FUku4U2b3/zDL5Y4
ZDF+M8JqL+N6H+kRkP+cJUOnstd1Fny8da+biZHgMC56kg4olldhDvNmEkmbTTmkFzL+NDEhlV7a
LUU363raUmSaclqgixeX4LkDXl4FCIOA4gTdRGsHHP4dTEt7foaJ3MGvfWLz/ShNa9IyKPkoRkzb
x6FrsNcjgO3iVztb+jWB+GA418a+WNTygMxT3hTdgUZWDkgUudzasmtn42uP/Hy1dnRAySzHIi6Y
03Fwc2AG6oys6kTBWHO0JnoNKPG+9n6i09ElRfuacvrLmRp8psgjQ11pCV45zVEMX5nUxoHs9sAb
MDy87Cil92kFjmaoWzXYDfxFrc5Reim1yZxZ3ecxJiU76+yiuaAe4MxvLjC5WTzxCXQz7PrEPZUv
INypjwSHpDzuU3Sx736sbn6k2gEIEAmkyiX5ThEqFSRh2+rW81abvoc+Dbcibvhj0aeVTn3MAbI/
kgiCR8AVk2uCxki9NvUhQs34pEutZlC4W2Mzw+OHzWH52PZg3CUHYXeKZf9L0/4WgDPWVMWU3N3c
zQKTG59Fy21aEwSsnhtY29kEtQyFTc3qWqPF/2q0XC8X0HGuwgdj9akfl/9FRO4GI5NDB2kEFeXu
VCe8+o/sV93e9sXgav9rQ7z7A5S5EfJzHmSeIruFsI77cGZeASmwbH9AlZKL5oaCQOHjq4FR3LoP
4qQw4WHkjBSCkZmGrOMd2h0MkN8zLKmsZ5DIlZNe959AGS2xFFTu0gHZzo15AF9JgbBs2yfYWK44
dxKdHMl9R1oSmziSJfkV55uPiaLmaYioXCni+pi4JKsJUR5QbAjLWJ+jNGmdwIXfPqUFDpLS3NY3
ihZzecSrs04iZfg5hYTuDAZmCJHntKFK/K3oiKx04eSs3Da07svH4MN1jxTC6gyAi8XKijnLz0Zc
IM0i+Zg4nPxbnKTpcTq+lIvfrrqKf8DPTf+l1/3YtZu8HfORty+1se6tflPNQlYWRXVdlDNGneYC
zbhMbZpWaOdhHyNXOEYoSn4znRDMi3wIokOcqyayT5rIBbPk8ONGbmOfehDhW7606V9+el6ZH9Ae
357O4ok4vpc8nwxgVZc8D/DW56mnC+V+sq9GSdwABSxjqhQ2sb+zflkRowAG+VOYWuDhsH7tvbWy
Z7hUySh0kvivnzIJmzhUs5Bfw5lMfDP6R4x2ZnKzqHXfcfht77tnyW4Ojw8inXd4k7tsIQ7SD25N
rYWkis2ol6BMbHjPYpLYOWiTOuGQx6K8I8j6dFRWStkK1oC/+6IjIlXpeKLrtdecMSaieqGuVuZ+
DL7tdfsEQpYcRkpyLhXKo06gYRmkAXf4S0jAOQRxStlnwRnxuWyBllH6P+vxUTuC863JrdAfbxNO
RdP4AU2RYSNq9eg9fgUc6/31CHveSkA5P9IzIgMCCqt81t9oCHe+b1gCkSuWqMQEnZ6EY16wh2ph
YB1Qg/UDwsfC9Fs+GS8HwKHefNfBPcA7xZJK44qkee5OzlTCYJYB9pqw6kToaIymME11FDeqxedi
cA+JaC9fXbZBB45a4wPuY/GcmFEN9Z58FeKYAatBDzV/4TOy2CoIrvLPz0ndntPk1NougCKSHik8
tPeh/pfGNVHLCVDc7efKMe4Wigjdwq0sQzCVwYGcGXyEvwm6l9+M75PaJGTL+atf/Q27wK/PElbu
OO2f5Mg5M0+ThdhghvutoBmM1JTcyJCnqjIzlq5UEujfMVoY/5nojekyMHKuV570w052LX+J3r0b
XZRr0eLXFc2WxqpdGUMqkr1HV6e+9HhJ7C8qX6UggHzD8gxbnob8/dH3NGd2qwnVbeaUn3VGQ9A1
5DGIHsIQFGiTqvWjcXnnHHQUiQXJIN+2W8s3B3f4Sl+g7GGRzuXtvcHu4mANc0HyfjB7Jyl3UnhY
2Ctf4YhKBmjSQ5NLPmpvts2czmE5Z6AicvC/PSiBxO3CLXzRotCWkOhTNbYXEiGOJ16YZQLt0/uo
F4u/4uuXq7J8Zo6U0kk7lBkCD/UA/EKQIRc8OYbFASCIEj/skCoFaUVyfnHzLYpvOA1zQBM+RizL
BMdV1n/KGyzlQhOzM5hKqUkdxb679+sD6ZGMjnS/+J3bPCHgCxCeOLfvaTzl7HyV346sPZJn7kpB
eDLsUbKNMCCtKKyyl6mTnzu7UOyo+Tzr4cWBHGGYCyVOqA4oFQ1Cpr0eOqB7qCEA4lZGGw4svGQW
Bv1uOgSorPGxUZt8mIsu9q6DepJhDalhscA/naUlNR14g59zLQcVHcs7yT15n1bEg1Jo1z7A9duK
599Obe5JMWk+VT3hIBy2+XMbDhfMrDhpm2PwKUiLHWlYZlh9eQLmdCAG1an2yWaKcNsn7JCPOsRK
geiceEt/shseGXa5Hk/KdhisOLJtyUR3coUKpCNhjQVw9KghzEKpdzGfuLHe2ZtnuKau6ChdQ1rG
KYen82opybNV7hL2WiOJmTacAGIAjWiT3UAWf4+DcnM0SL1wJJB2VEmXgeth8jF46cgN+bOyguEs
6vix9ZxMDxdEpknd7vrVGpmuLPT0I/jxJWgownaZYALJH+541NINPoAltLUR5a1w6MxvYLIcghI0
zijqLMpsslOUCOYAo5x0FyWEsHcbh3Xts9lrvLt8gCO91nWfOnP/I6dp/Y3TpoWdSEvqOqFRgUeg
liEcSkqXkeGJOyFchC1zU5HaTeAI6ZE9XS6shqz5GRwfswPcEZJ7zxIKEBQJBGsSW2dMxsgEnEqp
/jq3i+3E6kLTOPvMEVsTL8YJMF76Af8dnQP0PUw0T7zi4Gm+x/Z2n7jI/GqXEaRvVutXldHbZYA3
VcFRSXt/XSDfCPqEmFGFP/AFqCGfX49YQrEiTMeAHs7wCC/giU7sWLezrW7XlmH42jZpYuPqFz2N
kdOTdcMf1MvmL3Mz/HRkF5B2ym6Hw7uA770L0czKc21+MVQLLZrcfTpfCqtW5vuoe0YvScFEwJr3
gXAXKxdn4IFCVPO0h+T3mkE+I2iujkHkIkbUmGMirnKdiH6IBBL6t8esYbE3Sb7pM2CuwisUuoil
yjxQAB5e9GRnfjxZXJ5WmPNr19bn6MiGdlTE7fRuOs9vlLMbzaiujBIaU8AkRhXfPccOe8r5ws0w
xN3iUfj+ZLVuEm8HdLXFmGgqS7tNt2EIRqGE9LDsE3Eugg/pVmfQvvNwKnRL+FNPRUCX8T41ON8n
+iA1XN0kMn0qXPT7UNQ1T6udT8N6Oph+BG1bVxI/b7iiP5SbhZs8tEv0RcozmqWrbcjRHlN3utYp
/2H23qpff6qA3IufHir/ZZgNPHPFgd8iO8m6+AQO+DqmRFBJDUdVztDLnoaSy9i48KKBRE4INFK+
y170TXNg3EItrsC+zNXZk4Cwumi7ZBxipAno9MsEMuuNCT+P9UH8z5X9q1gjxaEqf2/nRofNPTuF
xEo6wgvuUj5TWMHwfCHjnRvDmSytk3IJ6125HGmhLGx1dRQfqsWkSj8Cr4EsBGlbYgbjhULdWDxN
ndLjcNiK91QnXqt0jwDkFde8x3SiX89N854VdtYZsEpYeAED6xfpMyx0V/V7Lry+IDFurygqp2zP
NY7MO/E2wr1vSTQ59Op1Wo1UyQYeTir+5Ebt99fY3S/bDsUY/CQiPp/McTzSDX2DUWIDYK/UjYG1
XuKOdXpi3okxKY6DE2y4N2H7unXMw2VlVVTBFxTobT6B4O/GC1euXLUTNuDv9d7BfQYlXYv1V9JI
/h+AZ9CHGpvhKIA35GSFMGcgITsyN4dS/+cBx6V2U6/k0Qq5zEC10GS1HVyeN82/IpWzDLF0/ejs
dTDIAdASWQ9hixbLmRRGRPEhrQBbfiDtmr2yCu6G6jm7P51eqqsg9JzAtXr0FpbUJvaNLI2wHCjh
GhykhKTOCPSAoh24JmFMZal/LlDnrnUdxJz2Jp33IMtO7Ote9UCm8nvDa1CItj8b1mzdSVol3P56
gPxyQ/6ri9Fw7mcqYp7F2yPgD/PD/Dvd2UBrvOw2oyaLiNQzLpJg7Tx2BJDkMJLvPydIIZJB3/Oo
wsennFCZi3wkNbYzh+uHc2HQvEanx3UcFdNheRqFY/A6QP8eAN6Oigv3E8wb69+j4bgMj+XgsUns
xXXRcG0dUKRzyKo9NWY79vCSveebhE9qj5VrC1XQ8ZrHKkwI1n+HPEuaKUuzzg1Ew2tfUZr4qLgq
ucutCPwiWosWqJIAfKaUOjXT4UUJG9NQsesB5cxGcFCrw+4Wckpg7Gi5gpO9qYFHkj0AD/aeiJvD
A59sOoH6zCIK64PzWIZcRG3m31UQDHOfSOH4JTe2HIRX9lGXMjgo2sJHeaL4es50XLq0U1wcyrf4
VlbRhalZAkgwEtXfhZPpi+4U73YrCB27wsacvr4NUffVdoFQZuz+s1CKzwcSSBDiBilQnkGuiWF9
IViGTEVZOCQjZXZwU83+XUzShFBCuKK4PnIYdCP11A6Z/tOHOAWPwqwYZuZUiDJYUu9vhd2BRAod
Y2mGlz2/bcaXjhwDY81mMzgka/ZCxSHz9f2oP8kbwH+sRTjJCHTbwZ1OPblpBcVRYCFsPZ+A94Wf
+lMhY8ThanjEkzLoOcpoRdkDMS8ms4daK1mRIX40qSsIre1XcNPmLFT3DY1fYjDEskD3PwgbWzdS
fgFZq/B59T7RoDeRex50fjePmXJf/29Gb3v99DuR9imeNBmFzj/emZC/c5e0uT3GkgjPyBSPubG1
EbyZTl5tKuphJlfWX7lak6qrsqZesz4ZpEBMSXYRNo+k14DlNPb0u7eLm+VcLTaMtgM0aii/kzJb
ih598Nf4W6p3HfHItLTpSR4m8eY+eZfEolSLl7n+RWEmOV51UDnL2yjybKIHl3wrDGNHGKnfFYlD
X+Im+phzvFTLJU/Yb7JwR75yoKPO5+hx3SQXi/+AaOEGUJOYo0jyDtV4oLO6d4NO7Sqlvzi5AuGy
FGNcBBqcz9P0dtJKvTxgJiB8dKIyACbKvZ7FzttL9bLsjo0hFZSfhaZRF18ES1x+gvBlBx+cBOM7
zrc6QanTEpdFXQfLNLz0fmqGhEYYgVDZI9r45cVHCb8tTnWQhY5l6Kxpp58V3XkBbddCyochoaY1
JfKv+fKHmau1cJzOvvJIfbFyAGXz9PjOxawHHAlpm2scl/o1IhoLYoS4+CuTzkalG+4SKmf3wBW7
VehRGtoof+o0iyOJ+HzxXZkJnagebQCCvRE/KEFBFFuzGo3niv5uekb8I057h55+Dd7GGQ/ZufgA
ws5x+vewAup97DeO1ZBsMM1ilQW7bFRFcRc+gjIW2HzFdqvSANPMkfF947seT2hypqr/4aJAbuNJ
toD5z1bc1Nwv+VHBrhqo+Vjp10yfgTQLiTYAhAHNsYP5QKRTotCP6kb2C30vw5J65NGkjteiVX0+
JHKbgFRlvIJ1kFrrGpnWOnijAWDfZv9/BSR/hEgP//VAtzJCyI0WaP1D1rVmjb8GaVSJ6bgWgtg3
sl0PzETjgWsHG9LCW61o/2qjkEPOqLjf0qazsyDgJOxzM87lui7nnzelZqTLrt8qYk/29RtJ2al2
cbBodMHBOugbg2uck4HXgg/i5z6VErX2ww+Cz1RgsbfILqYZ8x+FabbouSrtD303hQg8bHwKfjaZ
rSYbnqQv24t2PQtZZwXkVO5WKbibCxQAEWu71n5DhIz9PyjIXox/S0uFngya3HM9HC+H+/QgHDQg
WGlomrJzvncTE26GmYbzuSZjeSyMuOhgt4egPDIBhhrr56WfDECwYeTuUTZ1xDWO7ka1N1OBbJEc
j4/dWAlXUItTLQ3R03JubNAEGVOVhmLFBJf2jSuJGiNnj+92sqbURbB20FE/f3RYfa75IvKBr1AA
/PReVMPyyAIcmG9jSXjZRvvUmZTz1sW8oKBngKasRPMTl7rqNKeuVXA7RSHIafxUUQ92nYLIsgFD
U+FW5rGVKo76quxCNhu3DmFygixH2iAT5PDjmttLVx5ie9qluuSQB0Aa8uMk9m0Bl3wkmQO1yK7t
n/K1XvEg69U1LjRPaOtZNy4e6dJ3844NTVnrAVKXwF8FTMSiOMBRrJki8O4EEC3YnF911pf238Ut
ZFTgROoH/kRTBMcmKAv9SedTNMILhnZdVPfpbHw+PGpoMud3FRE6vc0yQqebIjpuYvM5wbknU1+a
NmNtV/Fc07ZioDR6ol/QU+4B6K4rVO6WXwA/feT4XQ2M9FW1L7N5Blbxf18bfjI8lGyNkiHsOwqr
zO/b3GrR2Eval3PiHM1XQlPuBEJZ2MgWGo0Hdl5nlhSu44ZjqPpFNON/vYzyJhuCzjER6uqbQZr6
gcjeG85MkoPHtGqfld1lIs6y08/qranyegOSZ3XbuzYZ63qj6ja0J/qOc0ucF1kUo8dhktUVuxPX
fYFyDYbBNrMjMSjor2bfef9ok6ml/NDCdwmDkQ96DUY7Tm0p1PlsDPfmyyxxsiBx5S1jK8DhYDhW
YYRVM53/ZqgEMfjUEwmo9XMT7uAhqi/rkayQfUH51YjdN51Y2UYCay3l9s3L9++P58flo6eXD8Fa
shvv6Ia8+AtQPtvpkJWOWlkFyWZT3ZjHCDZuQYZfuiI6gGdAyYkgBN1sQjc15JdDqTGIMy2LI105
lVgqryMjjk5V0uSE6tNwlQ0pYXHE3i8sq85kARTwEpT7igtMbuYxzmPQmGa3SkgpfhqpEQaR9mZL
uF6aaro1GEruIQl/p86NPQgn493xMstCmcRz0kGdHqX71kFhA639jhT/KQH/irmhz59iwRGtX3ua
koi707iH7XAAje+Atts/zORr/gaJq+PuH4aMYUmWg7J7ceEcCAs/wiR4n7Bu/tEnOEx7AT3V0iiF
H2IBfDdzn3YZ6RuPTllIQkZq7TrmpsGz1CyVxUyCrhPO/NQzF+R2PcQ2hbuho08/fKi60f7N2KFA
bAE/M2p/sgzphHqItP9blVX5X1iES9MUqvP3Sql94guqLQJHcw5RefpRg81f66hMJjnXPgfoG6nw
ODEDhpqrqvvhxnU1DVzv9HPiRDOMTkpb5avvhkeWe5RHFRskN+X6no6vzqPxGrCRuXnm1GpJmEfV
E+I3NLNq+5S9Y3sqnesQ2137vA6ulhpKd0Zgn4K2O0hQKSlX2e9UdptEz8k9+Y5BDQkIyki9aDhy
XGJMW29u1JuKMzZR87+MDt7Ljr7XRcq2EwlmpAJ1Pty3xnXsky/5xMFWVqkuH7ris7b9FSO5CiFk
PI4qHPUfq+JzWROCigI0Twt11E/YHymhqqMe++5EJr/7YMp0FsLZHvxDiITbQDCKc18g5wDrQ7Ay
pmVZWXmJy7sKlisXdEYRKFuWiJSccIVhliUb1+mldHDS8d+zD+zHxvrJV0l1/rdxT7y1Mm1dzoRD
+tO850mtavQ4GpzWC9ksG5jd+rREYLVESGQD1ReLAubPHtY8xjHIUIjazcfyA8Xih5NDFz/XrkHJ
SUQc4mguIQSChQtFIM++ZoLGpws8epfvgVmhGD9gSrUQrLjs1Rth9v67umUz/RuYlU3qqAIRrbvx
VspAEIYk9jXo1cf/O7B+k974ynNI6o/iSu811qMgZkVFyk95s83ayQha+rWgcfSXvGQU1uX9uFEX
fBeGlfiH69R/VyphM+A7rjMTVm4N0UmYh+yr9GR8N/fJrWAMjxISP2HwaBl4RCOk9y2H2ar7fnzs
WrDBBvXGNOxWqP3XFq4WQNXJdsqb+5/pYQWn+D3lNrNngS7FFj/bcimGZLJPnd1HYEVNmKeSBERu
QeJ4R3XeWTtPBLxXiGpUmjZjZk9WY8fBT2qFMleyMMYnf2wNqn2ayGAfO7n5eAaC0/IiUQZI0XBj
OyGGZoCI9f2U0jgZSM5o0H+L06KRXebswcsKRbJVZWJUnR3gP8YGx5lZagytNGJEFRWBjFlxv3wq
rFFJxCHYzdEA1NfeiWpL+6gUAScG8D2x8rQVZrYBSisfzsQYkGlTknOj5pjrTjCZqGRBMThy28N1
Sfg88tu0qPEPwRDnLgExT/3nYit7QTCIknGLeVsdrno/Dr+5ov7YSs2pxsDBa/o7e5QhFhBmuhYe
Uc59Hz6NSQzKv2c4XkFRAPFfe5GC6PNQDlDDEMzk48yNRymxzS2gUdUpiDJqqSoC9Of7QiQTfy+h
mWBPKL4R1b+XmxnMw329MvdZARDcuJcUDDG47fXki+/IZV4qIzm7kqkvytSYG3RTL8zSyCbH7Ldy
hhthAsb8rHSomIRfCNEoOz9kKX4CYQX4o4qLRZJRm2+UfYB6e1wGBsoK9OH12r6VIET7gfBjNvQo
CTUaKOaqcX6ZnbsJZiHXlLZIAd+Niqb5LvJ2j4jKoKShbgpBKz+ZUeeCRLUHN2XqXJHBJZQ3Qgx/
oRGPN60iPxQSAzplX+WYKvB/brceyn2aY/aT8FoYzi0p6MGVdE0y0aGmqB17BcqhsvpJHQD245n+
LwPNaScvreJEjGs2gOtSn3E9Ldlzw6oxlpKX9fZiMi3deBbvyZ7o1po00EBgcA5GUfxm5Aot3syW
v8pWw5Ri+UOtrWKmpg8fgOG2TCrNKYeWhTfe78+p8fuXYIR3FHzZxUhZ3gIHaTBQktXoCuHPPM/Q
qNk11S9hn05+KfI8gmMGeYb/HBwD/VhRqGyLyyZXbkVhfHGs6yJDAyRfJVUHXe+gk4FijXx7qX8B
kttbQ4p3hNPJ2b9yLZP29N94Wj1juQpdiV6eBFQi0EmsFFifXDzhErncCvhmOIyymyuM/lW8fxFl
ySCgUfF6+1A9wxqChg+aol45SOMDlvS7cGf19xB8P9NTVtO8WLxHieBuyU6Dr7ujMKKdBbeI9aUL
S3uGpSr3TgXfwLQxefEv9P1f/EJ0ZFPh/o+oCsCOa/SvL0heZCodyeQDYfJvSbMpEIhaSQiWl1Pp
zgQ1sOIaP+TV9TMgz4IVtwdWMIMN41IgA4viEpCyGIxs/Jw4P/BFpjYe7dO6+te6qWg+ODIHQkzY
sj603lzpoKAAxdntz3lF9j1x7Vwn2VivsCu4ZpvyA2fhPeOgTsK8LS+7Vlm9g6HhEKfAMRERtHyj
i8BT7+pngUNKzF3h3eI1hq4VFFJQA15W4QOdl7r3lYizEga1G89JZX7oAQa5L1waxhFCm5Q8Jtsx
IgMtRk/SiOjOwv0dEerLFP4xY5fR67IoJB/b+RAIgTTZDFaB/hRB79YU5EqpgM9GERWYY5wCUpmk
lm2dB5yJIa3sy+psiyZUt5KE/S/0GTA3PIFHPr+s8tX+T6VwAPVapRirSfWj5oUkHmpDJU6umtW5
EjHMVsPM5Q17iAeufTLrK+HD28PeTO8sPi9iItTQ0CP5ajQfcDdMbRTTXGpUWZqkxrzoMfqtW972
z+mdbiqKQu3iqLz/c1cMrU8nOqe1U+GZBcrqSx25dgWuLKnQnnrTY+NVJ6rgsEravI2Z6KhfnqIq
Da0pTrSJPp/LKNQuKFY+l1M0InRBBj0Vgoex4uE5aShvsg0YbEnIVcET5e/4PwpGn1zjPG2YGDAX
AuLXsHi6+BkbUtkG48uZoWGsHDJgxcriW2YeIbN5EDZeP7OjDLyl7rMB9vu0bqNbzeSeFAIKER+p
5eUy8S356j0IU+Ni+2YmP3vzHWDaGTxkt/qIgEDs4Q3AlPNg2q+n8/6vzYq+ACf5Oy/LcDTRtOS7
8URmFuwO2HqohnNUZZ0OBlOZ7o2ZWiuILwS8l4R4DzG7v7VBjBl3gcQ7E88N2MwlcorklXxXEgcD
qba1TvtXef4TxWny5Je87pTIsDxNCf9aOg0WMhw979Uwmc7rnUyi+Un7iZfbf63q0TMsq9vO8uVR
vHginipbUtduO/wJ+w/CionkM0gEayizvJANcNPNdiwW/qIX42tCY5DH3m2yR4lLuu57x9+M/xGB
+M2N8zHTlGvJLhOCgOTwN4Hwag1kSomM7TZgSBDwZaMdS1JiZSgBrXPvW+wybDZot7EYMLs+QAE5
gvpu9W5yOJOZCyl4qtwpyI8tU+DvOqFx1pGbr8DwWhG/yzzGgquG15JiH9U38K0ErWEfvsEk64qL
tSi3zxUxKFOEU0C8G57d/WqKqLrNWGvGXz+jeEh06Yh6lsEkrH41eTsn1mPaHl8uwPceLATrBzsW
OVJDJiS+2+RllMTKYglXhTIgcW60fL9KcQW6ROfwqBPBxGXD6XLmcVywYDDEFI+NhqdOmZUJ8p0I
A+okOTC0vVlUAyj1s09REEx4aRP12fQjkI53RP5s3NbSSZ1GYhw8bm0RPFF07i9GJZu9UOKiHz7d
o2JtfaHCdpcIgDO1I3kb0XG1QjXDMxRuiKJLV+sDhbOGYHWzWcNtPGGrBdU2qM7PxnCdVjv3XWtS
ChWoi9qNjFULqoGHFB5sKtZVskHcRCkYNAuJfdJxjl0ZqPV2sz7AP9UGhulQyUO3ganURwXn/HUr
vrNdoctSsEWsFmDEr/CH9CP1CxwqiqNbYY2Vw9J7OM3HYpdipaVnFsidKceutd4St7BmlfhqwfoO
AQSs9KeFuIlr5h7/58eO4M3htvJYyKvUlOG72/ZTnVR7lV921myts2L0IJqNbWY9Y3bBH4GV9mGW
jOK9PxZrBn4NfHWZVV/x35t/+UxmFQnT/5VMNRc2Zn9k34XZHTEVQ8o3L+AUQhby8VqU5bweJOR0
l2Q6YWmtEO+/3QTCuJ567kzyRuDkB2a5F1SfFQ1gocG5y8xGL9LzazbztNYKGNhpOlV0vXBgFiIg
dtqW8f615ycAOsnTojuAgWh/BXjg6W4TLdknLbcYWgthQmcGTGyEKsooOHwnD7ta9JnRz8r9qr/V
NE6WHMDxpKMDr5dgooLkgQdhNjjLkJtd7B9hla+qr+vPwCVIl9CNjq8GnWuFD4UEodlqsEdikJ5+
auSZJ4wIxLvQdYhi0/AklOYdUCqaG/+d8s9iSHB4s3QGJHd7KMNNletx6kzBtKUvhurUDp1wmgBv
Z/yNQQeMuLvzEjCCX1P8znOC1qmKUC3D+iqUxYfg5+bJnbGQuFGWE5AxnnqGqSQ7HCJzhqJaSgR2
esfxTrQuJYIWyCt8kDMdE/h19HHx4CuOUalw4sNb1/9ppTI7/LDQOhQMCAi6j5zrG287G9DSLzZ8
IjL70ffrFzaPhnUiBjaR+4MgwHIx5chLlIYW5yZMSF29QJTpDq7lKCfxp3veSss5mp0XyUfRP99s
vor6NpCVSUCpQVs9cLG9AATFPCo7aJYUF7fXUyysBYV82pPClT55JjK9t6DrAPZPQnh9DJfjEX2W
eexkqOPZZt8ZR+y/jMYgBesPzvswLV9HvUJpmd1qwUe5zL/kNe5i7HYd0k09hUYSLsPXJX30eU/3
xYG1qMA+ypAPrPcGQZr48QADOyRDmRSXGy9c5McgklRiCpc58j2/5t6Rb9kZK5lkZDd4sA5Rgn+3
KMSeG1pFf02UFP9vSQ2Lm0dTZm+aiHU+c3mYNxswKfMn/pyUp3RZ2S/Yad4U6iV33dD7tPC7UUJ0
edoGL/aJmaziWS2uCc2grgVoZa02Lhl9Vf5cr2CtwL3AO6ZMRyNaZkLoW9CqqAeKJl3BKyq4aVJB
MiiqzD9uaHw2q/2TkNBQoTtNHbGP2URvQZGgYvtoI2mVPk7Su5Ccdn8DoOAkHLpA+RWxhQ6zNn9T
ChvK5LZpUm8vIbDu3CaHReq6OqFqHgB2qk4PcL5IUG0EomXMiug58Hkq14th4FSabzhJ7PImQ5+7
X+soEz2CGj3DlUmKRx7RkiIkzaBDehkp+ARYhQVFm8GyrOmk+4V6aUh523gRCP2kBDN5LQ8l4NsP
CPy8z8V/3LqRQ5a8FKCKMFSo6LNAiJaGh9N/TrKQARLLJVwzNK+LX5cn1YlOnQSwWd2pYcNd/Z/m
UFQyWOtjGMQxc66VWndlMP85bNEHbegts8OOOjNgwiXgj6F7OoIa/nffpznsyYj5F6ixhR5MD9g0
BTpcoz8cXMA3heszasL6/D/w4QiKNWeAE19GnSrM1vliPqPtrroIGUufqt7wK00cUxGasKAUxbbJ
Ify/fb+wv9mG5zoubY19GTIZSkWRPBXWAKK9+/3S3zqcaonsSWI1bKzYF+4QNLES2Wgu9WmS5Ypc
/ob9y2vieN6BhPcH0yIwD9Wj1Y5V0UR1egfoWU9rj5WVUgKNbG7f0RtFH/p34ZwdLVM9wuZDFxGZ
tdoSkCeS7T9WeP4MjLo1n5jCvWfV8F8D6C2hpzxkFTSpmEKHYnlHHslE7JXzpNquafIurGxiQHGB
xfc373inCUOS8UOj0PFxDmpnabInTX9K5RSj1fcPCOdtcXNlMlwh6HAUKUoS2hSZD2AgDOF+iqUX
84fpVF9TGuDcvujrN5Lb7JmPuVsz8z2yuF8IrPxgmq0nz3xjy89tr8Jr2gRdbH5nPjlfcdP9xiVa
7RSn//CZqsmYlNnzTZBUvyam9rHRou2fTfYKSgrvLS8ohPbpWOZaUctIVLAWhv5iO0lIIjLmcKMg
K1FWwjyJKDLLGR1wai5wJe6mQpXKR/FerbOaUlsP4bgTBPTma1eJI+nFhQKGlI3SWWtRuHQO27SA
O50I7LVoWVKpSZi7kSDq7X4VDHuNrPzwIIYXXNf4CIs/3AqaxZhEkOvKvNo52+lrPflbyk5j7x0F
2Li3YeprpUQ+v4N08640AAYZJC/OHGFrPuqxdO19mkiCf+LTdIeuFXUMBSEYoMqT3AjneJFCJYkY
b2DRToTWgrr64RNJXCfSFPGEC+1FyRaBSGsWXLa9B60GLfGZrWXdKJn1qkaoHVza9czCS/4quDqm
IDFv5CDgrK9eZUcUKuPe1VBzjxc+oONVKaR6UOFa5hxzY+o0nJD/Gr3P93R7suDyGSs1k/xN35eH
fhPLauZKcNyG9CnI+PCmXG+Z+HnXgduGOgtriVHMlVstvjNIHTmMUD6sgzifLx5aao5fDDXrSx2f
jUi3P5AxcEGLanbB9P1Dt2pYsEGhtecK9L4bHfqB9Qw2prgA/4sed9ukkB+KiNCHtj2rtCBBUb9s
j51bJCZbkQ2pRKomsxI5kak36lg9Hyp4K9n8CAPbcYr+vj6ofQ+1UteGehU2NltN1tQpEKvB3bQp
ziclCYPB6xKzIKL7sF20+ir7bT7vpw+TGQFlGFwE66axk5wS18OQ/nvO03uAWVPlp5b9XQQbS0P4
7zH9jXdmDIbDfMbWs67GgXTzrnK02F9Xpe/aalWKgnGuWGySyKgbNqqE0pjIGT2wPGhQV7FXbQLr
tCdChAV3FJc6En5P8SZUR7FEXlWxhCy67xHk9AOXSG+wJtvkt4qv7jwzbtA5B+Cp2Mv7yWSHLoEq
RnyjYXeivdhxNjQEmbjfcFZ25LiJ+Roe3f2G1SUKsrEiSyHcc5LYhIO7Glydxr4rrPO3KrwUDzZn
woZ07PMDtl4jgZ0/TtLyhYZ8sVnqd9+o9VNd7qJsvLobH/kaXM4WSszaAJaiGWFmtMg4NNnd4vkg
h/eRPbTmbNnW/88pgPgGclvioLlI98PtwxnqePGtlaZay7X23AZe03m3wX3vaQNkQh3OX6Bqzk4D
Pj87zx2ZHxQ94emvNwWl++uYV96e9lvp0gPEWH7lWxhEIkb9xvKEq1Q1z8Rjqo5ZZ+0mS1+YMC7i
9Wtip5vExUvEUDM4TSo9qP5r83rxBJBy3JfWVQAVo5mbmuuJkZ4eq5KoxAymoy3ffwdnXJJ5VHf+
ImXv7cjg1TT3EvvYhJri9S67kJpNgRACf5S4PbOrnQjAzJTrRsIwXCC06gZ6yU/u7jWoS27yPTL5
YzDyoloXic7pE5AU6nhPpRpLXZ/GUsOyloQggsDg0gXNpejw7VOwXEtsm9kI2+0c9Cy5i8Abv/rn
fo0199WArvZq+xhPiVjLOjFjWGM+CIu+j0FlLsyg/anZTG3PlKH2T/enwSHfwZUNT0FTboo9cS4a
f+6cQ/uQQMn63I44mfBMx/H9Ay3c8heSWtClBYw7pn2ES0QOSuSWt02K/JftYTHGOpvfne11TXrd
zjx/lPtKttcwJJveDA1itxn3NbbAIhvgq6u+GKOVglKwRA3cCTP0payED04ZT+Tf5gzDdGYRkpFW
/+4NgEMW24P+Z+BCKcW4yn1+f0hFyRgoe3nE27cMpEFC0nONQD/+84ukKF9jYDJlkMCjTL7ID4vp
0Rg0BXP5jhd+k9ltE6VYHEYEXqF8Iy4houlei4vLNw0pxETe6BnYktoGAz/bI6D5u+gVTo3Zq5i7
zWDs1CKU+AWJIBge5UJGXLUwyvPX3+tTOCfa2T/rrlkUnPN5DNUgdR6SES01dJ/KN+xN8U5++uIS
rXsWO4zrHQK/l+5SYYfcTlCjE+cHSjvEsNdNjNnGGzzmC1CQizdKRizoxtPE0iPOtz5YqqO8Vh71
Go0Q/rYLpQLf1dC/XB/oD922OE2ejWm29N0rm4nwzMjBDvX6pxjBZaGpdOIjlPbK433uTym/P7i4
eer2er845m22Evfo5qvg/+dWJCS8Rm+p5QzFOZfl5FB3LnV++azP0/SQlVhXCu5m/bgKV/KjuEAv
KbjC92ShwkrdEAGPUbtAmtuHQ1lSJDuNEwqK6sxtkDfamursJI5MbpEXep5esNSluh4ob6V1rMBx
cJpwajfWnPXQ1j19+BU2+BOtZ5SFFo9mWnpQvxxexHn1FBtPIsytSqHfxGTOiQNuVDHlG2dPZoK1
w0/bYan780NTQA3dU5yYTJekoYniEv1bBe2yx4a0qEj4DPcx6wf0PAYhAhhnFJ429ncTjWlMTwtV
fXEqSZFcGpNQbaJgv9ozH6Vf9aRRSNzSLMIjhMSyEcaE1d3nyBbej6nO126xxfHXLW48t+p5DEDT
aXj5bU7rkDHLrF/fAyCZiYzWkApK/FQ4rV4ximX1DaPZZOY6V6WKHZb9txGB9StiTyj0R7XzBpMU
tTw8L8AqwQVPY9IqJR6wxFirggY3295JFerukm9eMdrtHIYdPQUgtOnKc3kKL2XwFBYou4G0qyum
WuoFRjqkxen9oDE+wy4KBicLZDURr9r3gpjqVJbK86Y9PDeOPKQscgbYuOuQzHW0LuSru3s3iOYH
mkCGpMp681vQZ6VDkBgzaq5IvtnplwwXIvCTrAjqH38MrXXrsdvqN2M3yHIbMoMsw3Y3kbD0Qw6X
de1fbYXE9uDi9ZLrVcROVyxjXYTWgNbff3rcmx3g55xMQSeoxo0Z+FApXoEpNKxQe+MoRsJ3TTPo
4rFID7yZlxRABibowHYiJVFO4RsxBVmlmAW+g85lpmIJQ4Wq+hUV+TyC2WKSgA4fp2E9xyZzTAIX
UE5Jk2BqVAzgLRVX959JxRxTRG1ROhfZgIeCcEm9MpBUl4uxUBnuHHbum80qmtXeYA87fadDqayP
2HQalT1YziSVbe4plT2nNuqFixnzr/uqpzbRQyqEzT1ARK3VBxO9UOJI4vToOjK0yNvAmi5pzAdz
EA0ab1nQmo7he0ELqvw3JLKUhbFsnjWmdIML/yR5JFk3ApVXVp9lYIviqJ/olkKGOXAoufQY7dWV
UuSjtDJM09kQQ+zD3Ox0mr8g1LO6lsdogwWw6491kU4ER2AZGfna1AzdOGRkwrf99FeLjUcaSnu3
fFG+W0aHCU8P2gbCXpetvJzBgZXIubFqAVkpVUwR1z8MeVb5bmQKgLyz+qpsBpCkTLNUQwHBhloF
9iHuR5ETsVHmHUwoTfNP0KztOZDp3Af67GWy0o3pPy/SrIAovLE543XpSzVnKkwCTOWnV+ys4bjN
pnh/FN9Ve1F6TCm1sj4LurT+DWZCza2Sr+fad4zbC1bG3eUfHQhj0LZtHb6u+z8ig8sY4dyWcnUh
myVrZg8Q1tCp38mXYR5c5qG2ZsI8j1u67HL7cK0Bg7yVffu7q7SufBb6vT5hdTe/Tex+/CCnqIU0
Hl0NDCPxxPsBU4w3ZgjkYqE4wDDxIo2JFYzDybAOSYE4UMVsya1EobTESOzF9+EPyFixGwy17GfE
reaq8xnVE3mB9TRhWUOn9ktaDFrGJQ818II446CRntecS4giNsw4gVAaDatASocwAK1dUddPiAo6
3gMmOXpYfAafKPyWFdMF9891mWbW7s/z4RkV8PJhKdCmSBcXpKPbqYzyZaoMe0RhDryIKlIUXP63
c3AjC60w8Q12LWwgAeGZoEXhfZpB+6OGVOdYU64ThXm8tUBQ3nxQzh3PZQRL/rqIuMoRMngCb0Nk
zqmofv3OrUP9OqzoWqPw7x/D9opyoZHDm0wlBgYvs8+l1ewy9jwzlD7vG0zlaRhjB0daIlJ4I0o3
jsjgcNx711HmhdIgQggQRzkUFycuNErJz3gs6uU9XbXRqX4xJ9+u1HyMuRQxtv07bT+cUPF1UDBA
Ql9sQrXl6+Ep4r90VN+k6XsYeihQUYYGF4GDguKQwvrk2qf/O5woMVl4k6y5ns0MtBaDiyXuQD5B
VnnGtaQJJM5cO6unLiV7dK0PROWTZcDry0DvDNf/TwaGNJ9wa6hls+Z6y1LvF3ry/t8Pk+gy4Rfu
E+L4IIhsA357EQGZ71GMAiLpJ9k/XtFu7y0FVBVfE/LKbEKVy1NIaGv/gn+05V/vcouD6/JB+UAa
Pkj4had8v9h248sEXZtaMPQSvayqw3R9A4gek2DxG+ASLZaiCdy/OWguKpiPIJAPH10KnMEEBoaV
pWVMvoR6mwpk/OxAzR6JVfGkHsk6vHdFy1YKko5vavM6XIssdYP14vVwQVhPN+eZNMX85ImTudnM
gK9JvoRB4K0+3XQYj54/VLWaBzRzHdXsQpQrrZRZoYsc2hlE18HevyD7xPQx8XPxY95aOQjMTJmk
bDDnL583uVp1MbAe3IfYsK+aX23wG4+CQiNCe6fVfmJFNWJJf0golOIEVFhaHPEGG/RcKq9Wgdmr
57DhSNXVhWd7OsfOrAMcPQOSqTVWrpzhECrX6XB7Nf0PYAHzXnBA3Q2o2MtSYo04ZErfWgkIlkdL
gHKEoyrc2jX1awgyB4gawiZzxeipd3L7Ei4Hclmi+JpmRXb+5n0Clou6nlaVq9XV1zTwKFSihBj5
75z38PM6lRmJTVkcOtdb8hP91Rt/vlEDdeF8xsX349iUVLqnL9KtKzomq7201Kti9whsxWusXZj7
lOyK7CcUIqAFLsMW2W98Hao+ZLtuVF1/w8bTh2JTmgWgCI8n3sTXwCQtGqfGDdsEb6vjgzu44X7V
ir42wi15XWWapMw2a27tZI/IP6oT9mrUnlyemp/rpgb5cITILNayFkZvu88VlmH3wfjDiKbnJCD/
2y6NhjhwoZodr6C7QiqJ5MywlPiIJNKi0mp7GMetM+6ezBfaIyq05slSjYEUgDjR4LJtVpldy3jj
e+RnoS1Nw5c88wGb4A59xIme8sGKNOj8c6Hk47vOTJ64FYM2w+5cW8FQgeh9xcNZpdu7lcGOIKNA
QzO7r+NIk4IMQbiyTG0nBkqIxJ92mns8xROHGsgHwSDFjB7a9ZZZpZIed/AyznqWk3ztHciIbDXZ
5acrkMPykuMoCl0cMwXjGha1QwUUXP/3/nH37hXEzjstqzj6Od6BHR7TyCgg/WLet2pdc9GNEO9r
JmQB8dzP6ZbVlnwViaVeT7cOKe2m0HgxnxqMGHE0kNYOuU8Hb8tH+pLwf+1UNsOXxbaOPS3slYS0
A46NshS353l2nLZl5VNqE/3JzTqbDsqMLt58JPWNgFEpOrAJyJrNZ8IE0pN6/jsKo9/Aql+JIJ7m
OaoJW1NuY0oc/lZid8FhvCmwggmAwNoLN+2ggdG9EiOD9UEsJXzHnV2jU4l6W7oqYC3BcBKTTW+C
yqsUzxgxYUJvHPFspmuaNMYu4szt7whINo1Txe0i756n4lCYv1hDnh6IA+F9gAEwDN4OiKEzZzIJ
DclyhgmXJyCXoLmRW6C7zYpMyeZrKB2orl6kD6YhscVyAMeSub7xip/ZVsDl1Q/1xQzt4GvF81c6
BxxHGrV6axUPIPSj6QSznhYuMxqKvF/nmqIYRcDGIyPmkvprj4plvzj4xDuuD7vUbs0HyznHyS0K
x3Dj9EOTEkVV5FDWTz6BikUnvDbzUwQ8aWTuQspg29JxuODeKirr1yyn2qVVNGgr/EH+yFm+tOTf
zr3YkurI0+aUwdE3Lgk0hJ0Ma8dBgQc7CvpEdDCImhaY31SpluR5Runkmy2Zrgwpl0Pg4zcoCNBf
xcKxoGdhx5TfLnC/fLyYKyC+JcnzgZNOsL6QYXNwluw8WgSyvqm2NNeXDC9+CTv8plt4nQ2c5zsK
A5S85kYNe6x8ebVVVcmaDzn/ee1FQykNc2EzlFZGEjXA6iJr8ZCRPdvHUzQ1ruA0XeuCkyOlni1L
iENHJ1JyWnqcsikQYDA8r/1CUqYKijfpyKa41Ng6/ry+X8XFl62dNF0oeMRF912PGnjFBRHGM47x
0avSbdA5vJEflYurdT0fig1/IgMKiPBgb4zQPFNSWUcOG27lh9tLjcccQpKsg9NCgaMHVY6nx8Ca
jjMdXHEmrv0dij1nJ3TvXhblvLi3PJgHcjdGqqI0jusWRH8IONZr7eSmaGue2x3IyiWU2hzZK9ae
jNDa6EZecUMqsNVPCMI2Oyt+y44V5X1xAeLF6OuuXbrIvQnC5czs0YOPwjl9vPp6QmaGY7fwbZ2h
iKdg4Q40OXoaozNXVDEGaMotco2zLmmckFiWJTrNByPZKO8tA12nrGrxyzBgLI1DCjFgjpNSEw4x
yydxIT7cz/Kk1Os7O3YUOfILj/PQn7+qhA1GVimoNYA62gvE4fL1QYY/a+MuDJwi5JKQKQNmGD72
8L7sIqAUcCXv5klazMQQGpNuPrBP97p+cWsHZG7fXpzxRedyXBrgpFg0FHSuaHHmbmPoJJd4BNDm
WH7kEcsFwvGItxdspbG4gJeBRl7wRh8jd32nmK+NcVDIWp+MyCKm+Pp9SuWtfbcij+fqn/ijiw0V
BsAvDgs7Lxei3mROxF+WxXy3daCHTMiNd4rNCPa6c708hjdjiEF/EF2rKNksMQMgEaNqI3DKN8aM
ffLWIXJP/vPgpCU1xS7fLKDPaEp+fHy/fS6ToK6STPQ3TYWbyV3mQ2bBq0u+jU/b9cL8htXkNkbW
yYo2qwf9RrCGJvlp7hdRFg8xOjZ6E97XBq769fw070mKvUVK9US/IZ7oH6fKCI9kjiPDWvL3Ucoy
/TVq39nk6f+wi0Rl+fXfb+4nbvFzgix93xUB10SAx5tQ80Tt0HQJG8WD4yzHCK63GefgwNavROJo
sEEcprG97UbVk6UuxGzWVrVpSw3Kln1zaHvRnwdtdaSgnaRg+Ozp7zn+HwVsqBTK6UM0qpFUauQ0
NyxasdDNKjICJ9wOtyFRB04bq0Q7hHBvcC6R+P+N6AgGK5pBB/pW8Nypm6+XROfSR9gFfeg9HxWp
TY5NvLErwY3z10E1Dss568mxdqsohK4oLoQ9gtCbgPazjb1eq2/bxaDqjnl3zxGGKsJHFjFI6AhR
vLd8IF2niZyMHxwrhH44E1IeNzXqabH82zLLmlIMnwtxwKrBdIHder5A+vkG5vD17Tk7QYAm7AxO
LXdpiacaoLrQQJx0ya2a7rgzdpZxeKxm59ghleM09Ul8/HeCDiYv0uK9HMUgQdqVPF9fUehuuh5N
M8e68aSMYWlId7qYMk6PQfhDw7R5KHvqVf8Erkdv/0tCKMnN4J5qPWUI5/tayLTsf1dl+xV0c5bc
RpFn8KcXw4BUjceAVhZHg3uuhNzYIWqmw1taCaA0BAIyJb1T4BQ6HfLGj1oPQZaPO7OcKUh5lbKW
wdRyXCc0QWypDwLo8cAvyNH4XNGPL+TpHOKwA7uQ7Xicn4l9CWBHXK4FGx/O+WVLtW3KIlHIxZw2
FQplF7dx2pkepgOBbYgZhcLB9sz8Clix8uFXu73+mdWeudlUICvU0+3Gw0qrcYOIEDQhN4sv+1oI
E7cVukwO4vYRXSj0aNd0gCQvOrbUcdT851kAjZio+Ij2pBMdMtzFULX/6I1a8d1GlHj+vRclLWwa
tvfG/KP5Tg+mPZ2Wud3c/VtVdPb+8T/8a2EUyjT/lKJGYCRseG6DC0DIe5mNn8QUNs9VkrNAUqcK
8n9F/5Xs8obN6irgzWL084OpEmW7rFoqnLeFGJcpUstFiaKWT17AHAwtO6bh955j9Rxd8qqoy3ox
wXs2ixFmqfynXtQVg4Rg4fWATe2W3N2i40wG+K2l635th0hKeSE1UoQ0FdydpNWFSAUWrH1E9qvv
7ssIr/EFVP6tZwXiHfyfrxZ2Chd8eBU1iSTPt2MutTu+BcuUmC5R8aROApW8OkupWWlAfzhM2Rk3
9iUxvuvZ2pBiCfPEqyrO0HjarsLDuuiK8x2KBwOE8bWf74ByDGMXjsu0y4rjZZDh5euX6gxCVwZ0
sZqizs+qNkFwtTx1OLUU6sNP8AWgVqY46yumQ9GA/8PS/4vlr5aul3f9qwiZYDlf38xDRpOfNxF5
kExPsPEhv3giPTDtANspkeMjFNgf+UJMauVSZmMzaBel3YXALewCxXYKjuryY63r9xOdSqFOgghd
Vu2NZ4+KfBs2WFVe1TX400xouPUa5mCgn2kn7nv47kJPTIR4BLScZLTCeIpuQ+0u99UN1xW1Xr25
PSeKYCtkIOiU1aGpbQldDeYHCNVZjrQBRwF6f2NFi32/A2pihW3Ny1d95p280I6mo/5xiI+lGOXI
X43KQOeGuL5tIY29FEcKiCfnkYSyKVyyr/jFHxtsDDuo5+A9b7YljDvzniy5ub6sWRBg3g2QvxGA
H4S2sOa5neFLiFgAYYP/Ynd6JdoY8/5HceHYdVbW67blI9R8zs5ko7zLbBaGB7azAhQbGxHS0FHd
RD4EPPGLH3HSxMWxpcQVeb1EUXURY3ljPZ7CT4LhAz5pEp68c0fuWecfT2Dn86Z1KEnMhViCXoo9
gTdhwbYtltH7PAaOr6CzafjvBDw56+tJFQEQq7lz6m4vxl4arjTqrOD7iudZZDwKgHqW2OzlMZdL
DidcVnqkMQTjhzlIhsUVSMeqWUCeBuon+yPPlXRdt4pjAQAYkjo32B5gdv7GzCTJ8us/JLXYj5dQ
yxxiiObiB3+nwXwcmM/zqYcBlNI4PPDgWw9PxUcES3TcfCr1X11Wsbp9t5Tw5doLPy8PgW4EsUGQ
vkoCMXLWxIZgNbEgZLSnmwTBy9ke31t8rram5KP3Qw7K15emp9yO1mx4+yCoI3DXpry4shAea7zW
muLBnqiCo8KQQgD8MB/VBOJvI8unYkBTBiFvlkw6X6lozGdSQ9hy1uvqzL5NiXdkZuqKCyv8Utpi
AtapFIQqS2zCROYknuRqYCvwpgLYJEAcisUzywT8G9sVHka0Ojcg3lM4MXwU+9IvPNIaK8V0SO72
N9p1sh3fVA2ckqAo4qKL1GANs4XXidjxXv9OTpe9d3zQwlkLHl+wXp/FD3k60+a2Qrbc7pScinmQ
tn4tzkz6j3gTgRX3mNoAnGIARfkut/V707RVgIhME2CoqrfCXDOaGi5dFvN93oftMi3FSNRQwZ/Q
3LTwnK+gAowxUQgoeErvyVd211wSvkUWUWl/izzJNCxhfRzFkUaHH1qPqQ0fAhqNlRC+O2uAdHrX
mhyrlAE+iyzjpOMWyi65UIdsa82mwJPwMEiz9jOw8iXCgQTygZ7o4oerXmuju2YubBCuKc2Ta5GH
iXuRaniXRgoFdCJAhnVf2KI+RJKKtFjMy3SBmeSa+JNJCah0YyeTjdMBmgj7fHXHkpA7uj0pshk4
WJPYopaRm4XXBytZOWcVxOkU0QAVh69pbO4h+t/U6veztGvmmsim4j7NHJZqSjrYsLuQnaC/xJFj
EL+aDLF1Z4yg4VD2mVTgssfKaulxKp8EFpVh3sLaF4ijXHTXGuikL2ZzKMb6G5YT8xe/plfgX4Em
/xEiAotJ9po9MVOA7VvZ7kZmgLQG5Yy1zxK7UnGKSidJJxhzpDHkJWv00z399GyPMJOJ1AdOfJiL
x/K/H2/PNi0PLzkRzbAbVFKQGo7IhpgopAdLORokDJ8JfMaPOiJTGe193BMNTlk/D0D3FIvYIVOg
QO3becliCb020AXynvEKiUSTllVhyxMe0jmBtR0NRika3eEc/pP+39O+TMJ+BZddG8o2qEvQKd9W
o5k0rX8K2k3E+7nGs94kPAzG0KoYyGxfK0O/S3QrQXgG5nOAMXyRTsn/AiX4K0yc8nLHiQ1xfUXz
gQHil/N7h8KFeLNa5b8xYz38bTsnVoXkwo42e2cIx5C/Jzq0zFSinkRWZT7/msnRWnrx9e80gppJ
F1a/dK2ff0H5fv5gQuGQELiR8y7FeIDUgPppSBSiL0GO4wO480VnHaCLTyIIVPkRLERM4tVBgUlf
Jiprx6KC75ckzJa0wN1yz8Xqku3ul4nN7jU7Ufcvt1hACpIa7xjPcg4MLnCBSBNKq7YsBUtC0v0I
+ILJ8MwM/AlFfLWHZP9IQ8iuWNf8cdo24IH+HagZU8AvaHjnCPtBjEV79Re0eU7RqrXYkufWXkVN
bs4Ws9IARffVsjWMMhsh0SVgsc5qbduBwzKi+eAQnQH4Ye6Qm6ajSqBj9lxpDnt7O1YcRSVKk8Et
muhrIS6P8jsfYrXKy2Y7DOCohPVi7b39SKbIOAozpRAmFSkz4kE4lWijk5/zWFqnvvKs6RYYsy7A
KLNg07JmHtzCWeKsD7bdscw54TmfUQbc4cgRL/PZJTFSGnIplXxHaHoPFzm0esfmgQZB7VLC/P+H
Na6gECmXXdcNM6aIr8NMpC1gloC/RhV8egP7yi7ODJFGWVpP0t0OvFyuatfe0GC9Zum7UWAwBRDU
BcLT7QjlInSG/V0UdlLrzjz3Qotez2c4n86t5e1DOjKBK0QKLx3a88kMVr9QyQyImqMB4v+AaiAm
XbHUvBfTvq5Vl/tpn+R/08jhmgocaEoPZ3FJCI5FkzXqAXIOB3YZejU416nPR880f0AGt4qeoNf8
Qat4zX1mB5XnjHwe2W350yooAKdqLHKB2EfvUy1tXr6+b7CuxyLdolHt+TMonvsCsizb1ej4uRNR
N8sGw5JDCPDbOZmKv2dZRs5KyQ7rBxWiWYmm/DTnb1Cb9LXNNB2ZUwW3boWDBqPDBql/6oN2ELMe
zDtzVdgJhzPJmTigS/ufNyV070EvOhJtVdU8z8u2NyO+8o6bDBNiPOW6F1ebND44aANtcuvHTbnh
QdZ8ROIEpVEcw9aCmGHCGiD5FRmUWqVLMH/iqZiui4myWLIhlmxTUofgSaGGiFEXdre9PC15lJhz
j5SR0MS2hC93JjmyN0nbpsaOqR8JxoGE0hRxz423BqyUntjif80OoJg1BoRSVk9+PXGYTyj7whc1
24iMltSy73nSMQtDgCNApwQgCrcgNAudci647r4ItRJkR0Mvd9HplC1comU1QOyhPTjMhojD0q+y
wctwo/V4Z1TtO0SbEQjQ1Aa79+CcbeHzL7MkDpVS+iC77R1x/EQJtOe1H5DmVpJ5oI8aFjtpl5E9
gW65FxiE4zCokcX5omqWe4dTVVOBwAdle1kxiPSRNLMIJYfT1J5aeq5o9LrZSQk2qbnimMFPEoS/
ixzbE7l70rLLNRAOGz8IW6ZMJbr0alGiLOPJT7fqdKd5EhBkCu6Spte4qlH7lco02krPYYGFyW5z
EdoNwl23cxe5cqCHdydyodjonkFcDdWDkGnI6slfiJVXMDqR5n5v6ohKPlWE8lGCLWsRGQlicCHH
nCUjfM1kfRRjWNEhVIHRR2PYeVM9thLRsASPl1IlqIyypl0fEY2lDwFADQeZ0366FQLnRfod6Asd
89lQ9pM8j4u7bHnJbRwAAmAxOre0PXD4jtHYxUhgSHZ9NaGTzwythAJQ1Qpg0VE1cKG20B2u+sMp
VRkEOKMRuteCMMJqG09/go5McoNBKGvryKV+TW2O8am6H2SSNN82Uaz990lAUquWqd+dA+QK0ozu
/kXkqg/KtToXA0SwmTTdfGrdknQqBSXuLAj3mJNqkIlYRAHsq5hLoIex4P7cClSJ7a2uEJg/ecBi
CuLu7H6p8qH0ufJ9cHbEbphjrH6jctnufIEtntxwcvJnyGxfjc8POzF6xoPsV24LcHLzq6V1BaWR
5DwUDNAdmA4p8oyl8FS3+kBQ15G4fKSmVQJVMUVRQ/NXdjNY910r9wM0KcTMq6ayY4mv/WoraUAB
4YQQj5BWxsGyXW+cf1DtX6yXCxWWTuyDTcpQSnCUQGRFtUG6foLPVfE9EHpw2FUh8mp4hcjYTdpL
qzv82aN5U8YCUs6uCkdc+ElmY89d+dTLeMBAcMo5sBsX2Xdz8qO2LstOUTZEu6Gre8iTY0iVVwmR
/ScKUuLKacvPMi7UxQ8111zqV1GHejWTJmPCVQA7KR7ZAWsLjFNhyx9tnYXEVQw8clwzlE17XG6T
2lU5tzoBLBog5tUzxMsRV98cLjUDOlUXBOncwEXDhJKsoevo0ZkY5W0ykrKLF5iCKf6vIVuxN8CW
4qbGYfnHt2RnzqmngGkqMNjlEetKbtGshf79ro5EERlOF8I7U1aYHHuskVCG0faAizJQX7mTidGj
aTARaSSHTadHwWE3mW9rdOF2JVvKqYZpTikeYztSuT23V9vprWtvLj9lJPUbGxQ7y+yEdalQKFmE
p8MM+YC7GBaw3rQ4I5qHaKZ7UkCaG/CfTj+4l+9LPePWHM8mGMhCJO6EaBGKcH/TLQR4GEvmA166
tDJHXdXjoPZPL6NeBMlYY4RhH3eYFVx+WTI97kerUREkH763BZG2/AXzcLt8WyOI9RpkUuRHDZ2w
vosCn4Q/mpkqc1z4JwJb8d9fYjSJ5jL7nKQp8CHd18v1pMECLRB2xVc+31NY0yBHriw3IpernCls
PkkB6IxUftm/fcUdaGu+RwP21tN8W+uEZ/7UlELQnmy4gViw/VNfouuH+oOqPMiUBhhW7o5mPBSc
xcj3L2uA9WOM3t/6SPdJ1hCIFvuJ+cFvthJ/UbWYT0YQyEaBeIufxCXaDhGhP04ijygbVgnSK/Zn
4bB+0/cyYkxLG/OVc6s5OXVjIEfjig+moBmpMrKx7Lp4e9bhRr0g//SWhmyiVycc1QQ0tUKzhusz
YBknvkIBskBmwd0+HgJsHkSDc7j3s4bfs/kg4NkR27U6vyxggN6lR9VjQuPY6qFVJSD7AGvwM0Lw
JVtC66rHGKlpCEuhurcaFotLkLHUiSt2V1axCyl9Nd+UVb8DDfbMd4OgTszoo0l3oWG9FqgqQN4J
dMpyUrSxh20zhf0yOaYNT4KslSvtcd/7C1QvyuoqdTcd7/HZXM18r+kOKGJ1gWwbBJXl8eTPsFMU
0tEVtTXBWCfBrnUSTe3J0qGldoMMLsVn+RkenRfd1TY6GpOK5cQffiHlRCB4CKWyfTt2IIC9husO
04RechXtWuS8rdjqNKsms9APqpisv3LwXtrNBbNfXgmK+ceiE+U4rU0PWc0cpUGWFvB1HevQmlcV
8B7Kbr+IMaL5GnU6SeWExJOagYClSa5zca9gB/fMiFyghYMhJap3XekqrS2p1js7cjCDYPgiCblR
SFelxdMSIYfH/V6jomOPNvV6xad7qHwyRUUH0TahC+gwpKlbm72EnnJ/rrrdFNX7Ra62FxNNDcml
XaJDXrZ7Xe4IOr5Y8EGASNK+Qbba5aNdabrpEOf5zjW9e892OaYHdAzjkJ8PU/rfqSMFqWx3KyD+
WKMVziM192i9cxGatxiN5k0OzOVMygmAMKwGlk1Rr8fIh/MtM4LEaUrRSp55X1TXWcAh0XYuNgK8
HMlfCm/mtsxA+EqILOicT24p0t+jbnbInZS9jP8Eek9+PbFDQ6RcJzj+1Ca8yWu0UVelykminlgX
qDf44utpWLONAU3jf1g227sIC1mw0hlIYZan8EsCD4uKuchK/OQdWguka63iNN8xdsTkMgD04stI
El/Btqkm3R/EEKXM+CnHsH0PwsovjCrRjhniAiZk/AMgLpI4P40Dz5/D4oMFJY+F9IOaJsfykRQK
Ajr/tFlJYAZsrZmETBtDvYBgqGXusNn/pfho4CGwX09UbYb+aUM1o0tvbuFw6LjE2kGY6A9p4GKB
nNcHR+CqKqbgDRH0bTup17qM+GR79Iq2K8n8izzgbwAKaAFtyelta4AGsZawfs3V4k9lYEpqdBUA
JHbfBZOst14AJI2oafMRViClG2+RqfGW3OQ4kXdVduE1J2U0sdja4WHoTg7rpSU+t1vpQ37tBT4r
9adIBLC9q0ED61/fFejM7Mdqk2DSZ9rVnIFpb6nmplzrOQUsIeeg9yLSKTUbzXq+RGpn2WzSFyqb
K7qpqRVXRLJZLg9nhTlOOOAHwLicSj8KIktltGxJYAM9S8HcRg+VZQwI+EHuTuuMph21t+HgfUGh
RxRa0H8p8biyA/PJp87uY1zbqCB4krTeMFJH3Hq+yKS1tMlgBL+Mk1000qScPkNMtSBpnOvGGZE9
/XQ0dP14HBYv2Qvk9UmqaaZqODNYgksTgobp4cEyhbcqOuEzbaiy+NqnUz7BhGGJCbxKuBcOycjP
3C4uHhVji7iEIiO7ENAuStmFeURPfu6TvYN2p9Blg5gQWWOMObjwWjLmwrnP9UUUCMXrbHLJlNr3
7o4PDdlSmyIlChSAtyzyV4fC5o45XOgRTiM1iW8UUy5YpQU0ECJ9OJiq6f0v0iiK0fz6yfpb8Zvl
9oQDWGZD0wkndfUO8xMVUhHg+1RUjptPuJOO1h3+Vs4E0Hu60UPX3o7w0sbEL7nOhHwHUbKIuT4Q
C42X3WYZ1qHAEMP+NXDCifmuPjAB4+Weo/2TYDdni/uDlJHD/VIgejj7i09X27xFMVTGujSLH/pZ
IB0fd+oIhkeFN+N2b4pTgrWaJi+RLPCimSNqMrc0cOtVWYWR/vxTDt0udoweMKq6kDnjMjZtejEs
fMuFUfcW+oTqOAQp1i8qtEIRxdUARwEUY9bNLAIL6K1EsKD2cXSnZZkWyn/iaP9mKGZhwk5qaomC
hXcuzE/n5VyXZJBbIH3d8BmUuOylCwYUVpv0U/3bTDZvydHPS0eA3M/KzEJbZXxbniITfm5wnu/Y
SmsOXsDkaKJelaxoW8I7lqHiESoLBBaZdFTAZx0GrbhoedlxbwSI1tr9FyHbSqYl/bpMk7zl6PUO
Ieg1NBwtnciVtZKn5BZ4oLQsiz75OwaC6RocOelpSzFNlez//JpTSjf2gt8TQcRRfjTkwjG/qnc5
OkjMZEVY6OeQ2zZbhvG8rt/JFSKhGizJsqD0n0xLvx5rAEpyAfxhh/1S36b9EethXzs7YG34Cz3k
DwamvTC/ENM4hCAmKc1JKzqsLtZoRQa+vMiknLZhJcTqvFgddbLJHj+ni2gWFQPnNEWXRpu7ngTS
F97y4Y53TEWshmEiArdz4mE5cplT/i3VC94nUhvKyr/MehZKs7kuH/ESWHOW4uYskdRzhIsb6qHL
IGKDsCokDe99mIvBxs7VgHIZSm/fgpzICHHnaNv1gxBpEomL7+55xddLNsB8sErs6rx/ZJBLFU3x
ia7eEJJK7hOC1T6FXkft89x4nfTS6VOQfjxYn26HKBkiP1KOi2+sGOip/BLYmiSj9KnoBdfX/MAg
eSpBw95IQJIyHiJxOnZh8y840yNt0VGiUdXCa4KnqoiOEyQPwqgoDU3ZIhX2xKLOZp4qBTltxL/J
CV5tXR2yx10aW5ZPl/JiV2bdNEAW2flfYHff14IfmKCD2SkgGy//siFLVRwokZSoL9mSeby0qS8/
Ss5CORUgsihQv1v0zVGW4Vd2afd8IXfGfuwSUNd6+nd53+AbeyyPur/zetQd2ya20uBr1oSG54wz
rWnDXqclw3tNl6/BiqDQOfGRMlxifXeZnX1CQG7JR0lblW6pyMjCdofZ2sFdumQLOfOAP1IRYJ6I
0PVPC16D0szWhJy5eCqmJvqSrTIjrxyDlyZzoR+ojfYRzKCdtScxtj7g9FYXxnvhah9m8hacZIU7
a3lAZK7HzEVdRH3tin/kcn2+/8XkX4b9LFhvd9QKq+5qzcFAFF6Qtr9qMIUxWujNZk6G9fkriaq7
IPU7b+khlC9sZbSfJEAmojRxTI+Fdh0IEvZnvKlzqGs1CkljFi6wKVPcA9PL+UWAy1dl14AcncmD
6mnEKXAEB9am97Jxp5tDGTF0yxAyHbjShHaDNRi2tYT5CR3fGlceDIXvhm9aEMj6kNr2v2ljecgj
CVNVc4oJuE4mUH5p9uXroOSVUkl8Gg85u7qS9qUDKeb+CcQLKippUgzdOYFnTj0TpafK2F8+E5Cy
dpGlSfb4aPxSZrGrFHHzO8FfYT5UXRYgbPv5anau6aYeOiDAH1fTDqrzaqdm3ife5avmd56QM4lV
w+n2ITxOvdxHZzOztLWB1RM70ALUCvax26vIbyhROKKFwI0P+Q8TAPfonIv/vSbgZD3xErXSGkei
nnjD9Ibe2Uq/ynU2zUw8e+65diBu9D3yfxs9UjDGF2mVCmb5ggQVJSBlhiQUXTPx/rofoYgDmVoZ
+9ybnVFDkDXhkd1zAAmHXaPbNjyLQD7Phyx8k3qZzo9/Dp0+ZBWhHsU6ZnFuGWv/wkn8CT+umnOS
HLwv5ep4QM+SWVmK9BKxj0mPhlZZem0L9eX/I4bgDwZEvEtd5q2jyAp+wG0d/ldcvHlTmMeh7/gA
PqUPj91j8iSrGFZl1KhWYhkBUwk1BdyWighziWAskT6B5sTslvs9cNnUBqAo6YefWT7dRylKfqEB
eq2vnBHEM/8PZrc/wOguwIxhw2cm8HWsXUUAcwKUgkyL59LMZTcWPteH8NkfnLn157zo4WFkc4H1
cp3S/M/WJ2yMK/trpjGq4DWbg9aVr3NQiMTuCus/yNFcLW76Fgci4Lkp1Ee+gEypDRw4MrNZkrrG
5Y5F/2ygOz8XHGrlAElc0rVpP93173tXZ37aG7IB0S3jIUBsU3mqxjYRn32jbLazis6+acEnvNK5
afP90qg75Xfk+iOR8c/2vpxzSdnb90RKi52lLEPbu9rOL9mT7xZmrtjNhwZVLNP9S13FKJ3P2xXd
JcSEIjDXz0JfmsyJOKWlwh1KLXoNYbwfWYhtk/HngajAB+nMu3mFsluSn7rTo4LtFWlWhwQeSLpT
7pILUesRMskrZ36McBTa/tuP1zNr+SMZ/SPGsmXDSXP5XsgIJEu65bOsChrvbzzVn+syafqKb/KW
qY8FzJBZ6Mp8RdAplsRemXxpbQ1OMeQxk0QxLuwcBc8lrPA/UWhyBhAoQS2RVaNNszfDJ+g1q7lY
OiKTxYhHtNza114RRT2KQSPxiKSlZDCTdsFR46PaZL0yfjW1y4WzrXPRHPYAhjYX9E+nDiMmVB/D
dTJrqRaWPwHl2RZmoaxbj+Hn/S5Q4ei57pmUGfe3NhCi28GLkpWVpfpGaUnVvlHn3fB8FAkf+lHn
n6ogYpUjv+HMrB9s5P3RxXCAA5uKjyujYMtry369r2RsVQZQI3GloFIxD8bvUDf8UQsVc4Ic3q7A
qqc2V07bzuWoRNCV7t0/7GM6AtTts7QriIHbB42a4hDIxwebwyzXT9frUTXs7sIa9Etpf4NQ1YgH
Nk7g9VcoWpmOXCTC9afXhvDrIOkC+9E014reTrLpByryLhNVdqU5GyZEGxt6JLRun4N86eoA9IOJ
cZHMIBpk8PkbYc9m4Md/n3gFVLz06JkbdQELjQUxbDStCgmuP7SopWpZwMiJTuAzoZJ61FSDB958
maDPObhWL2tfgKv/vFcLnKlfiTPRR9NfWOsS0irP01eDewejgey9PoZBj4xj/eitAqjJ2q4JAy1B
gv55Palv3FGKbGROf6RVFW/AWKYpszQmu6Y3irv+4nTyv19+W+TQ9fMzigbejMfgeD7r7nXeVTFM
qtvtmxvL90CMLrgjN4hDJTjamrJPQVbBsb9WcJBs/o1NBVtSwHP7NNUso17r9/ocAAyS3exml7nu
NM1hNn11v06tONU8TEosgKi0b3Q0xKQAENUZQ6fn/ld2ewxR9O+dgaZYoOEOeI0KkT7vHyaLfHN4
Nv0ectDe3qY1OpKz5mqk7gapUvWGzRw8hKc10iwROyoDVKgEMMN5v5KhQjxJpmMdgJtq7w85+uQe
Z89SoARQkKUGBgIOURpR0eS3NgYIBgYgnrES4ApkQkLn3SIwZgRW8AXPHpzeWBeRHUhAG6oxofxe
QIc8VRlsZC9JGbvyKkoPlHXhZAWqV9bkXjKmarJEEoiTkhrMr3Vy+Qz14ykumzH8zd5r271623fB
D0DY/ElpSTaxpF5pJrSenk6F2ZGdHAzNxg5DjNM5ZGp8urQzxUbzJZHoPEbP/rE3cfPXsg3gpX9i
ibc7M+tJ8U+O69JqTs86qfdiIM0uUnvehhg2uOWh2hW+BUmL++4+BSDDYG6UKtMBnFrofJGDvVDh
TwsM29GEaXb+q8PiyjtoLtiUsawVe2r6KtEfAI9TrXKb3poIthE9Kpfa4RMp2GCBeIgRYIenCitK
ANhieMvIu9lakhJdT2ipRcIc12dV/1CspkCksXN+PvGy3mxttT+YFxq0G2YYrw27us292NzFJIdt
i36nR8ECNNGavxObBlRVC24P9pkdivWRxHQQFKXNGZvkNFG2Yz26CmqwgO7AE+rweYAWMPgq/akM
RKJ40D30gbTRLlHN5mECRVwpkgwQIX5eLakyn6w4oza5apQbQH3T3Tg9fjZ574AZjwuTWrrqLdfL
avx9HEdMpJOgcYEqLypLqKe+CyLaMW/FrmmOAYmecPWLJYT1zcs5eNpMc3SFUJEKKa1C8npIl2j5
12D5B7i/cL/J4GycSujRUoWEVavgDcKbvLIdPzrq4qyq6aNcejeGoC3HSOLLZUlF638PEYZ7QELu
vPFf6Tezuee3bn4cP1F36h81gECSS1FDUYR+wyRgyMAYIs7BHA+RWDzj1mdatgr0HnOIfF+fGM7n
UzpQimfdnW7jlJNqI48pheZiTvoni4si1iQaPi8qLPo1qdR6jDGwNAvrkhsfqNFKcJBY8pmE4gB+
GYGhgoGkwPemQCIc0AxjtcBxY7BnTfBnZdOYqwQjMvE/FuZFj+Kl5dom6EB02CunaWQ9GRZeWNXQ
MBPSCHVZAZckLJ/ih3w+u8TPbMNfBBxYj2FRA3qI8NrBZDthY+IJpc9knLe4osITanrMmikW2mPV
rigIdrhkCl8tXmm+2TI4cjlSG3ppjgbdGt+Fdq8w9Do9Q+uj32ff0TiJpa2CIXVqMDa7OPaIhH1Z
t8/bVFzgxJdIecrXBrWXPydBT1iNV8Zl7A0UoR9+aVl3DqfrEKcmMZz+NkX86FhPtY/im5YHUy9Y
05i190LlPYymIQKgsgoJpNEiVOtlkGrSo9ws5MLBQCkQTBNgDodLT1Iw2xEBNJIQaDx8fBLPEnOO
8GfrPbKJYN0WoKluKuzZ0JggSS5Px1y+nVKN/ONu8umIcyy/lH2g6qs2iBclSuqFJUS8dXCp8vnN
z2pd9vTGilwEiLPuivOOIyM/vVI0ceajlKr32kYt6Qlv98xZQTCD4GimOZLVrjY2qdBiSBOL7ASH
fDN6wmT9vpGkQ13rCiZCNpQcpkEP9kfx8Z7BL1AAov6ZIcTQAzcNJZnJKFyF+QBhVPN0hF7c8G2K
IQXmz+44ZEQoMIOyjKi5N64vpORDYvFW6UyP5YJ3lMdtKNYviVhWIbqKiIyKR5L2BrZ/MIpm+p8b
1LgoyGaoUtlo02o0WQwRBGYEmgl+5hjlDjcg9kLzXCnNdI+oK0uBF2ZvKS3hQ93OJHzYfMCWLYyo
f4kZ0V2V3c0A5PJUS9VPjeHySLKb2QQqYzGAKRxfIMPv9CU4KGCeqJgYzYNL9rG11W+8sVRBUhN8
tlYL+LynDvbqyH/OzpkMqSJbMWqAjj5H9cayuilr8w9FCMnrS3eOAd5xqHb+YzJt+gMgcyFHa516
2r1fUAzytcY3puTBhtEuPhJPgYJOS6oLGSH5lB34csnhivukDGySPr0eduKJJeFZzawkKRQRSBRt
stn4H29VjpJt08B0OqqWTIGaxjB9J7VQ0Wr9Y904r/4Sb5oydsa72sQwygdClGfzi7/yLkjilXs4
T1oOqTYd8ol4EL7zzhH2yuFlWmGTD3He4I/bUHXOQTKEx2+83CjWjAgkAS3HNM9Jsv3wM2W/I11w
2ioNA5U+ZVJJig4BwD/CDCfUCFq+jXJHpHvCdbyb3EPeuL0//QBb1dvk37EQknAL7tHdDbvL+/6b
udNiWcPhyhGM/rFKC4oledW5AFdLJKu3usRIw+bhObXyTo5Tuivmo84O0j9GNYmnP1HYNs5Ecfgn
I4MQl6z2nLzhQV4hYoRBzRRXH5z/o1DOQYetC+VN2/RcOBP3V0EDYRXlQadhWYapv/8T4VXLlfUr
U6hnkual7D4rTsw2f2a5N2ASI3csnac1Tyn0LC+t8BxeWBfOAv8m4QjGHEsi5lcWstMLzMdEm5yh
PRbYCNHJuJ71I2GBglU+YdEKFNJ7wfNwKi23smyYnIw5SiY7wD+ZXOQJ5tppo7wyu0q12agjabSe
c+P99iqML222e1WcYXUsg9jMIqh96erPkTgCc7KzJyqnLflj/eVR7GMAGEAs5JvekhUlol4uuBSi
55yeo1sYfdUZ1Ap43IpK3unpDxBuPEsppeHSixASAehm0w8uu70BrZj8si4rXCZEJ/uwqyhFP9y5
FlBXDUp9DTwga4jU9H9Dz01v10itpeskodqD5Vhs2rVx44PzJLpV2oaGPl5ykly4z3nXabRpdRM+
GJfzRfODnUAEXTnP7EiCj40HTGQ9SlGZzh0IpE4fN0DeZGfn7lgwJ0ZFgfa7ZfOop3gktXG7LhKp
/daJbDsbuaTYJ6aUAetlEDWMvwbZ3dIM78F+aw8WlM5p+Fr3gtWJHE+wyYzU/M94lxwSM73vnRdo
/OW8+B28EAwrMplCgVJhHFecQEYcf2xXEMbVbD9fxpmODXVPHT45WUOUoJum1eWxZkEiT/nCzDdN
Kv1igGB9cb/m/5emYcOQVv1rm0lXwEufLREZK/u1Q08aNKvzwamii68SkL5+YS8/ncffUHmfTetv
v/agPzr+EUu+Op3nvANpmEaxBqTtOQhzw1FfazBgtp9l6jVa5PwdpZAPbVcSGDjlzIGQaZOSBz1A
q7ST0X61Gyn35W6volZjxG72FDFSil3S26xyAfUp66sNpNZpKVdrIOdZv7v3+lJuX1xHrLIkVWzF
rwzhxDW/V2U3+VhLIVirkrVl9UpBP8ClMFPqvFuHlxMeCyqJKpKFUhHkkG6ESqd67dMEWCg1RdfN
2hq3Lg5w82Kg38e4UD27ttSZhuOwKbDCCdS+UsfLrxXU+yDpZSws0LjhSp92oMQmTgBsPP0c967f
nuiT6vUpv9JDkNqgh9tQnD7YEEoFa7Br0DiI8mkDpd6K+YfQeZcPm6guK/PKvzi2fFG81oBGKEyZ
PD3M3RNCoWMQo6seih27DQMKhTcJzjO6jhppPMkdQQB3E5i2uSKpB45juE091Jq5nSYYyFiAqLiq
HECaJvIt020VpOJ3ZZZbOL8UXbINZLQ8RtuuJ3vxlO84DbomB/13v6eBi2mIHQEXEZYjBDAYd9yQ
uuLBFf0QFrc2fs2dUcSCHRKHYG+MevJXzrdvrc0nfD7uswC6tv2wgT82PL5TmCKprwtOIHvrvgtE
m3Ok1nz02Yhgz5EQ/TG6+h8SaGeQWIwkXjOkcFDCavBIZKecZv9Oa1QsD57r4T5JxGI6+58ypDEe
BSb3soQ+W9/Zub5OI3XJqgA1zUbOM1z0CVfSsevTE5tMD0jVt1S5PUIcZEofLsqbLQ5L6guZihpD
ity38xVScBX9PB0px0gI6aw2Mn+wIi2rlh2PxZFgMr8PJL90PTGfn4uvcVT4Lq4sMqKnr+62mVoZ
Xp8vehZ4CJ5MlySkqRPkgTYKr2SZShCrg8tEeValghaAPKd79QSB7TTKGDre6E7M2RvDrMBUartJ
4/hmsqdQ9EYWn07ATYrrP1Ow4ej6+F1+D8ogZ2gzX3SCGGTaiJDLAMVp9XvSzJUk19OkYFdicUZ8
e/6TFrHzGzzneZMO9q8032OBpcnvQQ9GP9I1rnbbWH37ZIKcAj8z+sQCU/TTi2PIbLH4qROE2k2T
8U71BwSr70+4RopyCNVcyDQ4LOEVBy79DJAgqK5Zaa2+iXq+IpiP8fJxJuio5ymGXQiYlIqWZiuW
MofeebkuZGHbL2l7hiEHXZJhhn6LPAOmfINHPxZH2AP0xgGFnldx4FfhzuC5ih2WgmdsTKNGTeg+
3sF7YvrXS7AfYFZi+d51pHpCz9hXRoXDhwsJ9QhrsM/wg0/ZTDU01EFh2Pqm6vR93i8l6qmpPBF9
s2uGqGyaMIt1jCf6G9K4dERqrqOgi1y38ow/v8NlB0tVnFvo4HU8Az9L6RzHex+2Xdu4X9Qsj7Xj
T/q/yU/2S0M5pWbPo8uFGXsLoWZPHEfKkqJO77q+gGCtYCkUbRxPoUeaX3/+YRqtCuxbYUhPZ8kP
ZOl3EonqyVAtc3HqqLyMMNRL/dpe1hd46L+wQgACxE6iCSAtOYm1HjUQfo3ICJeYaWVCzRgSO+ir
DPaQzttiztIzMelWpejV8Nxiv7U0+pMcyObLeQzQALKAGoxxWWurCCieg07Rzz/0yxejR70Aqd4u
0iJn6WqPNwBBsMrj2Aa+BR/un4lfwjo7GfQCHM1IaH4J+RmwjHNUrHcvJxAX8LSyTXe5wSe0Q64K
BMv9+wOSnvY3JPn2p7DZ1KjxVI67/tNdcl0N5Xbb9SZDPtXWS/Cio+8iCfAdrLLO8UKdqBBzKFZg
C9lq14k+eb4lSnb0utomNr8RNJ69elLzpdfjXDZNPXGbts4RoZI6wN1nUqtWqPuddvQIamrIm41d
Z71bIK0u143p3ls3XnTaM50Dh59PK0FnQ/x0jvw2j1sCeox+d+0O4YoWDvFZxNkdMdcEBmKdJzAz
n3nLUv0mD5HlQlQSak8UX91TYDwNZ+1vsZ9xBAOtZ8flDXHt2fQNTIZR3Mc2CCb83eCajCBIwG6Z
mny5TbT5szfslJpylppcX9V+93SIqVrM3kEt7q/QtLgvBFNFErxLBJ/DcLqiTpcXjaZRFZkJ3J18
oaUhSmXCZFmr+jJObly0oYvM3oXvajOf73V+BbEefbrkXNBFyI1tVZtBym00VHHw5jfPMGTxbaDO
ebKvzAEKe/AmFZj9uXDH0H1SmsRl0ee25RcP8KS9H49DNB7QgmdUYEEbzpHxi48BALR1InQAB2km
TA/1l4e0lpKQ66NpKAdlfyHw9DyKdZKNeZb9njprPKA8YiMYVTvtMcTuJRXilszQZuVG5hXtNwFQ
gnyQsDQTlZ/lllAT6M80SVB23D2pfzwSd0ex7hRQjAqO2l1XSjU+xwE9TdM1RJvufG7quivB24GY
mrpPHA73bu9/awjkVzD6QO4lMyrQTtZDy2CbhFOguuZySQkAw1TkQxtNdrqXbStMEMHIDpeqmsV1
vw/aWoN2pb8x2drI0w0TkJyVSxCfd7EjWSOC99NAyGjcOKZNieIdHV0yapymDCtL4zZ4l6FoicIb
h3uKzArS5BuX+CrwVhO/ttMk7sUz8+RaxEcxWkLR/udSXWZSCzAn/o1fxAmtGBggw42vU6fxYFZe
gGrJNqHeGJN/YLUIinUnlGwr0Vo+ORLOEQVcKHU0b7nKeUPIgibKT/P4SYxwpfK/kDlAiQ9DSgCP
+84odfCPz/ZbgDT6JSUOZHCmgwoXSkKamykUpjgwdwLl2A9Nf1Hx6k2z9KgfanllVP23lUMulPc6
rsd0OnWhfHHbbjANrND+oIP1Czt9Y6fklU7xRp4d8XIcUSYr1FuPzcla2GJFY1+nqaUscuK1Krc1
f4XR/CI3Ika+HOg+X5cRhraXBCkR60H3zNN/3sQlKnnY/L4a6TAq8YEjNsk8agkRwzboeFB/dRxN
rg/di/jutWzWS4aQJLQmpRAsF/5MS27k3uew+RzXa7EIe7H9iq7KNHGCHDsGFZUD5mUlnH5ool1S
Wctks099JChTHLv3lwzKDyePHNWoktXVylM4oi407qVczrx8XnVtf/IOmEHbBQ9Uyt7QKUBEAxQw
4xfb9k02uGzjwYwiIu4DaddRCLpg4ddAxy6V65kkcCV9/2oro8XPDEvGpe9EhOivUZLdD2L+MyDm
lWgZ8B2goTTKgV8SgrdLI6KpQMla0Qo40Kt8OI5NLpfOeI5WRrrOnbDIlXWi3FeJ4cLgP5U4gc68
5WKOJ54YJivppAF93As+c6I+CV3BWFQRxkhKbls/HjXVTtWyieVjNv5Y9jWc1OqghaHwu26yfDvm
a5QOCh4SaHbTNQlOh3NncnzVvOgDCOt5Q9nGF1G/6PwJM0APOPEAA+HmTBXQEuBLk0GinLAUoW+8
v1DE2DTRn+ni/8HXPE+td8VxawvWwaAVfcKWlSF6RFdsi802bhFKlIo6JXP3M7h3mZRsBSeME+SB
FBVQDqVMw38uylyA2Igui0Ozna4liir7gdekewLoFCST5sG6TKNQhUoSoPvX6srA3ru7aTxLWHpA
4+4XRekDrILoF0y9IDRLQnMcwDVrdTGLfg78U0ez+ZQbGskV8NulMlabl5C8g/mrASEe22EMdh/p
HULH6cBDF9haednzD+qntNauWSMbR9o3i+Xm/ElS1oQzZX1NdIsaHhj/rGEtudbHjA/XbwPBCQDV
V9XqszrqSxk1uZSFbpXZhRUiBJoQZF3RO3fOn18nxniTOg6bsSGi/qMBnZQANLQqKIGeqkE+8wO9
ntncyuQPvfYIHwRj9DQ1C7VP3p8PfhBYC6NxLjHGSszT89LPbwiJJWP+UcM1UcYP/GYdAK3Xr390
4DrNgwlQ8I6Bxia4QExWgWbfIXRYjtqG+FIa8KPJNf342RljXq6Z6v76+d08asBDriiutcG2FXWF
JpE9WuNNL4FxODz9lybbviY9zR67q1XRjRAmhGUn0gDrYvsEn1Gn9231S6keEi9QjUiQFyVe+6JN
uGnV8dezH+CzITau/tP1PwFh1y9Qpo4Ic4OnKwkFfedhXjI36nADjiSVpp9YbpDR9qFBQc716l5K
ZBqpC3+MwD9DbAS9g3IiwI78MVOHSHPukfb4s/hN6Vpmw8nzHqMNkLdRswJMaE6EyJYoIIZklgGf
NMi+B7KqNoe7BV+sn7XWPVDxBoc5svHF7ADHs4n9jb1LGs+pKS6+uhnupSZeK2Ty5QcVntxXwX1d
lzOzuHT2iI6Kx4A9lds0CfqyfLtGPUYGStxGQBttrUoYBRSR3pw+NQIiYTNUVinyWLTXha/9+qSq
xqR5F3W7q+yxVTpQ1BON1iJLeUrVelHpKgcN5Gc+xnBFJ0E1/dDWPZ2IV31FdxrVmKNTojUS4g3u
pYgJK2IHkJSNZ23AJXZUd2872eYxpv3BLyOum9Wpo9jp6WtofnJS6I2vHsU6MdxdOvzmcWAImTpg
Wj3Li/81l9U5bCy/860WyVEHOBvsuqptYqNHT0iAGEJoN+bC2fB/Xsns1IcjX98kpccutK+JVQAC
MHeV+tEVEc9j6BnNZfzSGrTMlKeLcvdY/KJvmpY9J33cIxqeyAr4TsuHZKcSc4vQjTMGflJEFd8s
ZDn5rKamjyqkCd20UIA7EK+mDiR3Yu3mntztcIa9vGeDexOdeZD3ZaLkLuSAv+w0qQRcvXlUrZoe
c8PbECPX+JJMVMAK3dDbyCHVl+b4N9tzj1Z3E3o1+w7FTbIpK5b+FmKlyp3BE+hcddSEMl9AK8hP
XTOSGHz35MT7elPBxo7EMb41q6WJ1e9OpJELgkHPqhGR/UYLjaJ8ybmeFz2JLIdIGVN2QpBFFgfb
f+1DBRi4QNIpRGtCesi5DCNXLSIqoSQbd/H1kZcBw9sWiGLOps8d0lytT8ZZ3aAXBhvuXkjudKUH
JxcLGOSMmRRGZ6yH2o41tRsvQA4Dc3esUnrl/w+wfftetNwFgmEBE4QS9tnzhOx2jsog5Fadg8a+
sX5fENfPeORKWLwi7NBN8rj1qGU+BlOH01gtTQOX1xQ+b2ibmhvos5wdvcTfwmeylmopPNI0t3gf
E0YlVpzWffDSgQdBnPoj/fRW/v5oCBvuoSrzvZ0XoC8nJu07h7HonojzMUrtBPylYBuMfKm81sHR
sLQEBLSKiOwkqvxGkszeMhDVDUgZsKKYTuf2x2l6OouwnkhULRe6eErKZ2e57+QJ/W1qzWkNQ1VR
/wMVG0jXgjSsCsvdSI4+UDcmOIbPrSljAOPsJ+PhJv6GTNRimMIPtth6IOeCGu+SKPAYMwqw3Ky2
oDwCtnKZ9XlYFHCRnaeIqNiMph/YRjQtAbpEAvpRRlm8nf9/3b/vAAJBdc9iwNbtvkn45OU/C116
oSojUYii7rV8z7CR2o5QWs1Z2Ru22QGRJdaL/5VHZzOHx1IQrwHAECXkhwGOOrYV4GYVxX25G1jB
jb+NFKZo0zvLRum62zcLGFWfOqRRNUmlLytygm5Le3gZ8xpJlIsQy88UrjrGT1GRY6VlpFORs28a
QpWYAF04pzRwZIrF9Xex7hEVx9PQELs/XNys5dDTTohD28DXrYXsBI+6HtQZD8vMyLHOdf1psbji
OtM4eQ7IP74bC9pPmfnlyhq+/qcAwuq/a6lV+jq2s0qolWd0hetOEZ7ZwzzR4ljZDW6P6iqpzbTr
YFq+O8+5B3dKy/ukGCEsFh7paMVvr8yXbCPXcXTZPRF4pOhPM2qYZCPNVe+JTFqs76ibI5X0X1To
67WGyHojk7kIgm57myX61DzJnP1tgjQdzI3hUHVvRnq4gy0ftvs1ckHFeWS/xDFNX5ulIifC+HWV
mtuIyZ/KcMkpGGdez93EIFCD38FbF7acUZrjkKf8bi0RdfPyXWhB0+Uc6fKBTU1hB6aKY2UzE8rq
WoJptdwaBwtj7hqa4L6jkuLzO6qhjRBHHPdiEY4Lk5+wq0vEXx0o8kkZS5pqfAgjNP1KcQMufKgo
mDYmkzPM2ipKkl4ADlMTsmQz3S+2lJqTvwbTmHgtbeEAhJhAOiKbIE4OogiIHDh5xhEVCYymXeG4
S9wn1BXlnRO5DFoKmxyNqf4IuPqZq5GVRnb6HzgUic46d97smUwHGWPblncao+xcqkPIw445vqbm
R5pAkxhseyGGNXdNnzmluK9BNBxNflszUzJhZR6FRAPssUUuSwB2sHBUC1XZt9rbFbfdq78ekB0c
1bP8i+NsObnW0FP+hC610zUxoH+/mJX60wubEho/K/pl6kGBR6Ou9BPz1UclMF5QXxi6KCn85++B
HpTDUT70FXCECHRe4sL078rHGwq0aLj0TquJX2GShJCggBbeIxZ1EGgD+O0WAOAQEdO7FDs2h6l/
O0oK03nwIVeZNbuJWKoz046My1vIEZqbQEjUozDAiCY0RWlortbOmBkZbPk5W23mbXGrWtR+11FY
OZ6bm54hLSNPlGJg3zthPJ6dBBwRWAOxt0HbDI7wDreSw5Rk90z30jyGe2rXGFZ1VAIm/kzszOQH
jOwgwtseuttLiyEfUBVqe78EBDZrNtEDQEPX1qOwa6AyWszLzzdWP7ZTN0G2+gHqtmUwJpTe6nL7
lFCwwXtHkkEM1HTzj+tuwEHMDlhNlxL9XsgUw9yGu4mfA/Pr1CW/s3h502J5PvMOsZBU69ng1Uru
wMQkHy2vtUcsPY17PKkTcUsk6Imn9KGaphSAmOgZ8KoEPgB3qLXtlZvDVsCdcklCAKxCSmk4SCKu
1jwHYIs1nFA+wU5kCZ2kKv2cRUgg8IMxstL+W+WUquolOTgU18HBBiI2gxJz6USSWdBX1E/cie3t
3owshnJORIejPlUSsG8a5eq9pmeXFfw29scxEHE0a1Rn2XQN41EbYIwTEOsr/seHuXYfz31vJPou
KHL9r2L5jjKzmiKzMdH8zT64584rAQUFobX0aSL/mdwoyzYxr5QcKtKiMoMaw89A1BdJSOWXjVLI
FODxWbJ070Kq/BC+zxyDhK2HJsTxTF5yyfe180BoLBC8a2ufhrRJ8YVTN0nVTzshj3cqk0Jm/MLC
KJ3ePm8PHWkdXZxQeK0akwZZL5MsNC5A0BULdSgQZc0K5G2e5f9eceISIxb9iWEJ65QAIB/4mUIk
GDhUHnbmkPrwrrH34ysD+zXKbS9QtuonvUPVoeJ1Hnv3e6/kaW1yfP1iPfq7d3ZEYUdHh6RBkMjH
ddhvPIysfgw6zv2QptwwTxxC+VyJri2clzciBPDjuKpfk0LqcKtyNMTJR4ESqKhyJ9d7mIE7dj3x
l5tIz9CZPVkNjqf/zfPU51Xy4fo7YlDIr+t7Q3GqbX4BVxLplsFhx3IKpo65tCr/hDyieJuh4aVA
u/fkuH1llSRnpIx2FuT6Ndp9fM1mG+Ymn+3qal2X09bxZ7gZILA2xMi/nF8vtx/LD2ZKbtUTBxsN
uF9szcYLCKBG2LOb87pjKbBDeYXlGHQZRxTUnpEIq22+9aLcxd3OQtqtaQhpSQvuivL3g+g7K+YT
lq1wybw+D/7iX3pmyZ576Yy7umh8K+pULzhDbNapfzeOjpfqvnBwNGLQTl8dpYpZ8yPK9IJ+/75k
mq/YF8NEN5bSZh92vgwd+dMfThH3Rm64QE7MHXCWMv3ejJnvBpAAe4E4slbQA4HstDcSDjf/IArv
PXcP3qtURGRVGFajSCsPDGm0+VXVB+HKsOo3zVTjERel/Vk2EmF7qFeZBNJNViopoo5y8gJzmX9E
Jpe0+aHtDDqUTfd/vB9rjX7oJsjY4V3Sk4RN2xRrdw5Uw1J+Nz+YKqIqSxDYIqVj50PFm5o5Ay1T
6R+Z32jLFZoRIsR67rLqH5o+P41z/zkC25G9XSKQX4jH3NzgI62n08QE2WXdYEluGXyMcPkGn0xp
bXjd2GgpHl+ETVSaW9L0wwlayJ/1WskrWnC/0Q1TZFu9HK4d7644wuetlQRq+MdLDXwIKfa6gJsl
V+4eyMPqdXo5sGylayqLP7aBRDxO8zrBlh4CHCc+0/7dAO0NjtNoRQ5U6lxDf7TC11p1UxqalAop
LgNSIGbGJdOYu+u4VRV+Q7y8C+emJ+cqSpeGHyqdynbgzC5x2GnnyRztzWQfWqNnH2yJ1khLtQWj
E6gDGnvYG9bvjIdpXjMcOBDPE1rjnir4D/Zm/AMO0f2uRaoQDVnVx1i1qLEe+WJOTE8lpEy0F+aW
P89U5ToZVEvjnmyX+W31oKcD1Bh7BJ2cP7RceG5QTZWouQnbjVRgv+stZdyaCSk88u0BncI2QwCU
XHvIRh8npgsem/N4q50qg5TNJIsoR4YuBzolLcAqedoWh/fKUGEUk9tgh1xA/SWpW0W+XUEy4Hbj
sJ85Gx0poyo91B6eNFRjurvh7JEy8yI6I+cdTSJY6HjNdxZlBekOrVCWKoCZGLh296sx4lt4X7Bo
jsMLaEU5QP+nFqPkewg7HWG9GD8U5DuQABBKjAlwNyvwLfAuqcvS4uiXu95Ny6ilWqZILBQLcQvE
I0BsHzlGNXj/GqqWbMhxZEDlkJDLgTioRVUnNhXEkGlw+OMelx5UYfvFzHLhuqm/cQ19aFAtFAwM
4stmnENyaXkc5Am9WQf63kLJBV7mksvWy8R3ey3Kj+bFir6P9d9HToYZ6A7RRJYxWivcKz5iyU0g
fR1dls7zokTPDzEQQzZwSOWbksCNhMlJgU8Y96HBUhow1gbQTK43IWHzikguqiOf2GIAZiYDetOx
/EalgTf79SCStYukI7yrwSDOfMhjhducmtcn3O+tfsuvXepZcbMwqgsbtRw7aUh7JPHTzrGT4+RE
L3cbHMU8beNCmkEkn2Uv9UJdHI5dy+rur2aEGPez0yUT/4+NzyQumMe0o/Al+J5HBDJPm9/82v+b
NJtywluGoSaKLlFmkcv379Bo2mMcfidZiuxspSky7yY9LimPRl1ntpOa3Pe/uvCMeplrrKd7J/gx
NoQoyofajafyKYJ+C4CzxZz1hnpMZgrwl90yCDEZ/zIlFvlVjSFXJHcyokvZGgRJk+lWq7pwEVLE
JxccTmhfGsJ9tIQ/wM5tfI4HIV3R75wBaYGiLrYWef8nVlq9KXaZhkjRdIDg2qbU6ZzLpllzzf6B
gRTjmvurdwSB8kQeQGqqCE7b3A+YulqaDv1QTbL5B107fYDkEK/9zu1WL3hY4j3XrgHgFy7HhDkt
eilnCTdOb7Fm2a7hkwNhP8j4Xu/qFVKvvrngscftYBTQSGzGIh7Q6tFNHw/0Qdx3NIGrITm/3kk/
/CXZLI4S/bsNWsbgt0OVd2VvXT+wnaWNcIpscP/32aLIsNuKImGDzOtG1Lgl6CvRf2YgSIOkZQ9q
W5Y0W2/GMFhcPzSnS6abDLMEntCJjpON0OKUOW3xCRXzakTnM7YWe/ucgPu27MoE2FV68euw9iPP
fEuXvx1dBtSlPGjUGb+krQyhPaHuwwGk6TLaAS/qzdSMCeptInKxIT0Y4mNVAep1ADpvY7mPc/rN
JdGWABPwLGkmIGbAdJzIV6XbMZxIQyaRlYRg4KGWGPXgnpMAwXkxSzlMzFz67ts3pFqlQbkueS5V
HP0zmIvDqjo+aKhtxYakThGiumEP/pgqLx9jrP/4TIDSKp2Jbqz5Zxl4/zYy+9B1Uf/bwjjkKcVq
D3EZ8/fQy+Gd8qRJuqlZCwLiJOjERPsRwUMaY5MfBohYy7saco+6dd+/vOHNLMoB3aRumWskIfAr
l8ExsgOaORIVdoPDlDTeFiOfTuD+FcdgTjl1Qfdx4pgp8IY1DHbJHDo8Gt3s/Tqk025mPaxop7KE
6HpzCcgSJ7iEioUPSkvczZynnGmNsm+NcByOnAz2WqfMwsm3HpXI+W3vRooxV0cabNfQAFQjIeRM
dipmrw+7k8NNXG5uxIcHi3YNSzy/43l11ou+bLp1Owp8bTvoLevD42XTAJ7Un5aFzYZcowihemzr
K6k0lhwqg4rHx1F4xf3hsrIqW1bRQTqYl4xaQmSsH7zCrSvnpMqivXulIuB0IE0S5GQoqASDsNFY
M4Mgu0By5HHs7HfUeKfSzKvNv4ZxvTCJAhu+NIIlNlndN0kuiWJtmm6182Z2AFYqeSLco519sv4B
+oBj3Q7pHJENd+koSMQwiE2fk/UDMNU4+5+jpKb8QJ15gHIibypD5xOLOkkGBVR+wNvGL2R4Jc2+
CQ6rj/ToSX4JC4EjSRIZTRp/P+TBgGfje5tmxJ1nqV6KXbKgKksKfbvz6AJtqbLf3A3RAAcJeJwT
RWK7ZGOvHrXeP8xeUYDTOhzhH/o8MZ1LTZmMNE3Ulk+BXR1fYRuECSUY3HtqYm5wolZKzt7cVqeT
cAGVUvxZUeteyHz8cHg4EOUMKADxBuiK6tAevirH70TX5KZNkgsGydGSZkmdiukQPWQnTjikMMSp
guLhxrZy1CxxFIIUzQiR6FkJNYD9UAhZO/Hgq1Nr4yzzXy4/m6QvFde1BJVmtzfZpr30A+Ujnexv
aNDLbPbyTwExS3488A7weD4fsQ2EW56g8bPSsoPe0Efn3LglLagIourNjF91+W7CAzMJPjRrnx1d
54KnoDx7YpcGt1cOJD48kIFgGgaxFoNGWDdFZKePknC1qkzFOn47gx729HStHf1oEjobLLk58q05
NzRqAWqAWqczNnkSH537BV46bK0zmRKB7aYqsmcITIZxMkl6CLjxAHuhvVDrR2Q5FckrLXkP03cP
LZNcD0NNGS0QZgnQe6lNYFkVqgYmjxbcQziGq+ihlkjhvE1LnGMBC4Yk0i0cAIhdEqrIlHfO3bJd
8oljvdhBRb/YEXzcsb46HPoSFmhr5BVghW9jeDrM1VoMoPWsyipzmzrH5QQLVIJlQ4co4d9LnRGp
L3VqQijR4vnfjUkm9TicArsQ/mp/rW/IPo9LCTzqsFlxfV3+x8PrWpwIr2C/UYfR7YnGLFOIQ+e5
C6xBZAXZBJvpkU0NciIuQ2c5mGerLI7ZL9cNl6RzCjeUDqoCUM6f+Uyw0q1IzTlVuoBEZy8EUFbQ
ZCJoT8UFm3COkdboefWojPGxk3trfRw5tQH4aeVdealt5/KJnMGsCPT+GXW3Fbk98b3pdwsuNgKQ
72dilvgOYIsUEqMnQ0ALRQ78Aj54ouNMAtsKizgf22NV3iA1EEvWF5/mN1h/VDsX6L4hfWtTmdx8
BD7jtso0IRMZkEaZpTI8ofhLUc6L/k8QKl0/evR/hcSKYyzQowpDETW7pNLoVePn0onAeA1alLZ6
HGQWD9N3hKI9Ji7mNCHEhwqZnhgK9T9MIavUaOIWfRRcJtOgrb0it+9s59P2t9Ghii2CZKntJ3EO
+BoeyQDZC9YVhQonuWYRV+DldYAYQtrQWJcC7807ME2QA3RSEDo6SjbHoZ0wS8xXE5cMGhEl1Ljj
AiIdmG8UoOVRPVc4g24BDh0j49FSFoyorfkK5ZfMoZ24CXOFtEunsutOCr57bTQ6vIqZ/FW/YpLB
bC863XOfkV/XtGCX8Px/epwAdPxCnIjXHTGat7VLoWpNeIaf5MXiNfiS26XY7BhaMPcGyBBu8kog
yyNrHAtl+DZ+Biv9I6lzFcsIMrKBkVb9dUmELkd8htlWqD+fxNv+hR+VioR9C3FzusSYyC10GlHz
fm9/q+cvylrsb+LvFK/XywqHib/RTLmIjCr5FSVFU07H6VkoRBZCnLikvqIAA2IapBB7tVgDH78W
2qRJgPzpnPCgQWs8kGyZLoKwqCPqS9NpZN8j6Gi7z7EsYpXcfrmvcKeFWCiAvjlrR0MlFOR+iYp5
TkDB4giBCq5ckSRLYP68HFQcgZAyh64wGIQaFn7nxg97GBWaJ2Wgy0BFloAxJ78zj/0k4CCsOOU7
AT7ZuUmILEwfnx+qFyIycGJuCumoMyKYoAYm0/ZA5fGoCsq29nIde77eb9CGxz32EOBLPXW/83m7
hchQRCIP81aFwIk5JcvoAPkjj844xlR1i97l07OEPyqF8HoBpS+9FkE6EfuT//3JSU2QlOSvbd+e
hm/0LVIlgNIvrmiBhGxxQrC7oenEYetBERv/IxwxBAXUgnmqRE0TP9DfNcT37L/5aOP8dpEW3DMk
4dQ60L1F+i4c92z4CvEkPQiYQVYSfPDFPknqhqQQUvFRxeVxQxbVDzCbATphsPDKJF9gTDXdjCDU
rTtu8xkEH7B1re4sG5XZIm6QxJfCkUee6S/n6N5YzovOoFe3cDsAr839tbEQC4Otlu/sZjpaEYMD
93pivwSFRo+qvjTdyt2fkBKsm0OPC5ZdcnVQR7UhEj+KxHgjlnc+TBgLZH+7vGE5faa3ERjWstpr
p4RsmB3YzK+8vGllYD77j8nWwgqIIZw94USRYjSzbNE7BajFGZBJJXzJwws5kFFMwBXuj96ixNxW
imKWpaSY+Ce6eJV3R2UlJ4qb/ROIetlhkM6EgSY+lmPSSr5KwNvLY3oRK5OlPnuH1/6zU6/uT3uj
fZyPi0QNF9XzKrBwOYxhrfHSGLEs8swwQ0xJIKyfazUMGpDZxo5p9qHiL/Gk9xCOkw0iNVQ1PYJ1
6LrVrGpgDGgK+bMrUtOe7looWyEYqMv2H68A/262vsSDRma21H1OsvqWt+9t4uUqX0g/IyWjN5Hg
0iCY0GacsZzfQql5tMMXZzOyci8BsG7swjfRsRF0wlOYzKaT+zt1NQdOEgkklS0aiVT6AGwQt+wR
nkSagGhX2t6ZZamyPXYGacS0S+hjulkWQ1OQxxjChTpLoYAyJ4/rvHoNqWMISBXmKQyyiRwrgKU8
M8unTz4jTVkW76wKzshLoTF9uEL4OfL+VO42W6+L6LExS43Qz6y2ARST1BJtcn6EZ4mqzVtIHwoI
+kLBEpi2NGdHEhcP87mc1kqP4VyLmxKt782YRrS7bG04tkmXduzFsr+D0zaj4n8spXhJvJ2Rn761
AzxNsBqjo95CZYUFGnDKfgTfEWqmVI9A7j2i/66Ep9qSuljs3DabWlfcFANxcVg1g52JSMb+CMsT
K4e1doxGawiHUuJmZkmvwaRUCiTwYBsbezJEklnq9UoD32nJbFikDORouueksuD+fr6vyd9mY0at
TIzVNZhBSbX3YGVPCdED4IfKd6lC/D9UnU4Rt82YfjY3DPuXk+yumMKZ7Cp18T6Mf4lGhLuOx0+L
7ZnmNaXS6JYrR1WFZeEpaxb76kKeQTwb6FfgPUj4CSydqDtdevm4kvZZ89/NTPC4l/eBWOk/tX32
ggHigDBGNQ7feGB4hyhGIADvteFbk072tu8PEYf7LN0+71FnOn4RlCG2nZeg4sJGmoR8xGoJ90T1
pPEfd0wD+rljYUEs/9cuZcKQrrsKWvRCmnaot9eYXppxX6i+JBlvAYDxjaW4Xpf2uPRan+SI6zsm
dIQ/IBt01GRvTu/Sf37t76mZOVhkuUQsfBIv0VjrhK92OXGTh5Y/k/KgwxPUOwwScpY+2Kc88ZaE
3tVtaWUm7VHlYY88VQ1aaM766azXUGiM6Y7iP/49E8ytxeED8aHWCQqT9cPI+5hGp/tu2a+F2zjx
QZBWaD9hfqb8j01pujLcAijo6A1LRGcw5+bN1Oqt4E2EiDGhcCu7RcGyTby0WCRjTW3peVSrV8tV
eGVGmXy5Vu0WS5upm+E45Hj0JxkS6+hL3IrPM2lVRB9y1niHeq2xPLVezV9NgrSCV5oQxoVKUnvU
P/VqHG1HDag5JgxM3QJOK8H7nHnB6WOGP6T1ly9HRm/xwSKbzsOB5FFlHv720CXPMAIj4kw/dGP4
2NU6X8t+qNzGY9xwQjUlP2mY1Bf71D6QvAk+4+klnKEX8UKzRFTOv0xZbbUtioLc+bX4GCEcdyMF
OBf32Ayp6cLW2601+oylpFuoONFGqJsckrRtSFcfwYDC/n56pA5yKxAexn/LeYD6uKyz9FHFevMs
2XWbK8zbaOc7ngaMjptFLYY5gAPnuImhi+5h4HYN0vSnEde1Bpy6yY8LldGP52YR/u1hpOIZQiuy
BAgYNLbabWfF1YIoD9TglV/nl9SGGm4Nhw6mgUzykC7pPsTcSIwqjtozuZYAvADPCEU4eAw/bfdv
LPF9veT5O80QVOUi5CmY2a0KkVtJjEPzxZ+rJwqpyUhkhXW627fpP/jjiIDt0zOVeSfAEkNLAPNf
H+OT99GQj7+cFQ9BVk1c3jtlCVcm/4gcln2y+PCOZWtS5Xt5GaJQhal+i+42Ji3Pv+EoPiycUiXu
OFihc2GI2tLh8gQwAmXhhNBqmj6k/UYAl1ryNZB12N9rmq7aaP4V086C0AlJoOuaYRZU0oYHHi7i
cIK6fQWyDSOFF2baPkbVxb6PJnADlSULjrZHHsVQWikZJq1rIcn3su+bo/W1pDC6tApMVupZKSCR
5np8ashP1cCz2tJ9Zq0xf8Cb4Ty3Xy1oLVP2OFJLh/zLFTauyzZtwM2qgk8x1Unvz2xcespiev8s
jgb8rQ7hzg3jnR2poyEutHiH/BEPG2JhqxvS4f+CWeWYiQrGPDRwwNMwRW5mcZuhCFvwVP30e4O5
sHn7Nj5TYqDJCp/lpCsx8y/mS7a8rKSeSEFPOd90c0bIpZXIoPzdgjrugq32J6r421HYsxwiY2Ex
3xjNYYafPcc6KsHq5+Dld75mNXp8/FmGXx0S4Ram8ov6H0P+CfrjureN4gk8CAz6l6xoR5EESs8X
GABXIpgjQox5V1LY0IA3LUKXWxO5HwaU/FQl25Askh0X1yORVudU6s/FTnN76Ex1RqHKKAcNfGAM
8aPWzp/RDrnZOx79BlK6YppzzHr+Pfv9OXSfHhvNHLkmCCQ4T9KV8ZPCSQYPXJ486o8aOnYArdwD
frxkxwks6dUezlKyPGmbJdzOF/HiGvkywom0zq04ZSYtUlqZcsSS/Og7AyH4ChcT9P6w9Ebp155V
sYX+XDZq4SjREN9P9jPsyAS36y861m1aCZGP7+Jj/BXZpFwAieRiSQEzKwqSSsgHMuDyCA8HnB9G
D0mYSn4WKW2oaHf8fj+OmVwWJCky18e1BoJzCnS2IrOrOXBnJ0nLe81Gv9fIdXqmAbX/vTwAWcqx
YY0ijzVitdoHkpobKpaz0NJE4RKIggkVR/S2pjGB+KOaviaTuehr1opToOjWHDCqy3PsOQ5Od+1H
w0xg5PN1sz5Ib/gaep4Fn0dLaec8rjEQHm7ePjDIaCt1tnob47NS+pqK2tFnkl60gHyCEjqm0dtE
1Mth+1BguVLE6MEhupBlSvw0MVR2bRdumqzLF/mqiyzOiM1//E+tDcKEBbQST7lLGAU3Xp/8JB6d
vQVRZW+lCVwp1gK2IqSe709RtQZ2lQfcqeqvR1wwgTVYwZjMTP0II+Koyn0yx8W80VgGRyApZIwT
KrsTT0YK4v2h7nrvLl0PQRVZDEgh7PWvbJTLNp476C3SqNHqImQe5JI/+bWD/ENzJAjwCa8BJRop
+Bl5TGakH9In2H/ZPdWjN54cPEV+m3HAnIkxMOY4j3eBp68xexaMznAE32gwDo29olIMqUzNyUI6
jgbhRz6wGqoiK2OYb8idUXgaGgHol8SlhUmmzmEJ0gG2A7ZhHmoC/5ilJG+LsbaJhE+82QLuVJ5j
5ywUXRs7+l/wZduqlPT0yT0kNyEFRgjHWVDSuE54BxTIp6MHHSOW1FqZbkRcFC0H312TADD22hwR
iAAc1gQqmEFlR0cehnSVPnT/zAEokXqkEhqNS8hKMmRV/E+rNf+VtvQ2K4vbLnZhUR4DgydbYjAM
ZnPZkJxF70RaE8+jOYEidgEYG58wdANs5l0svFxA+IXVVpzPMggxGlYExVh44KBKXBp+b/s5VL2r
JE3Pqk/1vk+A/dupCqrZGw6MQ9U4nwDrfGIgOXRG0ExISNm1DCmdGQ/qF01AbYmzg2pPvt+bkeXX
imdtzOScw4IObA/Nc1m3H4ufJQ3jDYnE5iwd6EMA94O9ZiKJbqTFz1rPiOF5HvqHETkuPcYJQIwk
K8zMmyIzW7mD6V1fh9w/Gop4OvBQHjsHLC+gTxqq2muZYYZEei3OojBakXU/3FV8ROft68+tDQks
o4gQDWDyTgvDRXcRPH9aqo/EXvfHz8rTbWruPQOc81NA2Fl4byYkcdxlPMRJQ2lsWh6RPd+997J6
6sv8ll4F3zPNv/KIgnvAgAzYGDyP5Ws3GOMmEy+FZ/GUU4ODex5tIaE63EFCBrZ65KUlHotAD7ex
Ps8ptR8SMU8CZqHjOTIZNVJdB2wNEsinA6G5vytqTI8DkT2bizWujKdgKOIjQ0fEbuuM7Bsn//yW
GNtNisyZEKTymuvuSNv2piDqtmn1dpT0x9h7VzPl8nbGG1tzQxA4tkIAuWdzG84vfMnCeI8uzNZd
RB0UNjEi51vdenZt8F+ofIZBGBnVzg8SsnSINjmINaL1o6cCxnx0WghLDQSEkr0ND7zZq/qXRW7v
2BY6zC8gFdabOb0Qwx8X3dMz2JxvYd+5B74rmL/aVmi/Max/S32ovTCM0it9OixfDXna5SEJY/Rj
1THLSzaI5rZm3Mm3kza/zVV1qmEFbt6Ki5zJR1YyBYWrT0T1s39yeCsDmx/JjIpUMrnDriNxAlm/
lVzBYWMsXye0rpmDxHHnnrq2zOYtkUCNpMr1Tm4pCFsD8i9ESbNn3wr3/UauK2mcm+enuHWwdmFO
Z+Q63vCJtx0B9+IvCvm/0OZysaf5bpD2Cd2lhdIzmkM74uKFRIBSpHXm/IaW2CQHEbIj0Wz7j/uK
QGmuvXrcFBFcURBzdVep04ShQ7OXBdrgEXKSDw0VBhcJfEfjhJ4ma6WKD01LQ8vXMaMZBwMfr08a
GlmIiAJLJaTx4HX2t7e9p2szVrsh60VubC0R1Yab8jBdDe2Xw08OM0hc3JbbdBcm8gqfrD4XoKLk
0Azb67lb1B1nscZeQuT4wg+L3euRi1I4ozN2OtOBRGucRB1uXvOBQrOFJOlrdSDn0FropdKJDbvF
d4Kl7cObhYC54DnC1tKtY0b+XcsNDhEO9hD0umMa15qQANaPHhAqK5zZ8mb4hSFgdh4Wz2jRpG1d
Vlqb6j5NHzqGQGKbYT60y61ShNZARKPOwWlxfA0nmK0D4ie3zHsG3cqJ0YVFDS6lTSS18zsskTo3
A1EPV8A8eb6HIKSyQroJoK5HUCPclAQd40jxpRcHIkKPb/jc0E/95XmjiLTpk0oT10qQNWN9nr6O
kGTGBAqDEnwylztMyFiap5WvvPSq6ZrCtoj94QI4j6xEeT8HkbaiYj8DkzOL1aFulQigbZrXs9n4
RrXD6bjfJPkD36uMWGpvGp+v/chJBx2LWxLGL0TppYybiFRmSt3Yf9zi2KT0b0cKvZU8+z1Y6YHQ
yGoKKU8KdYrYtilZhoqHeXhbbM3vTdfOFoRDafQkAtK7RkvOsCLP/qWCf3Z992xYhGRaK8N2hpQd
8+GoZzDKAzEOnjOmdSpbtAFue+F1sA5yY4juawl0wP8qDtJP1aXBdVbY/cZ0I/DCTF9yS2DbO0kN
oqn53DaW5+2k7dodyKgNaqP1UwRzihdn28Ep4J1mI/Hf9u8AOo8AY1VHmxlJkwQ38FBlfCnhaGiX
FFZbMwDdAnf5bBjmplzyNG4rUJxzAfaJeISjMCbbHo/4HxeWoKFFpAS0hjjqre6oriYrk0LMocmG
yFxUxipEU1Ww8pwzYQLTcDI07bHC3jqiZatzdRnKQdzxOYDPSVuOo2Y+I8XU7B/e05j+7i0uXD4M
It6vCboQfr1yW9caGlDMTs4G48WJYusqfvbGjHZUn2CUfTg6iCIBrpeg5fBsMBO6WrLstKn8mwur
rGyLfHLLMG+sbuYvuEjr5yuIo/DOT+A+zdppE2tFGqBQRDgVXoqOzEgYbP7YJihhvZYa56dqsQDq
p6wtcSpeT+OoH3U+dITgA52x/VqnY1Rm2UGJPB220lEs6VJsx8b9jn5/F5pmFWakQdZvxbUkugjO
59XXviOBqaVWSBiq6o+gBaYNEFHln/b5hmTOAa1hMQ8Pbs/PB6KmeO2FL4r9fgBlPmEB1+56D127
8ZDGgxYP0c+cQ13tyIn07GNPX9qOrmHBFYU6WzKMx9O8IyihxTdPZJ+Vwd4Z5ZQ+7RXptFpwA0ZR
4m7o4fhiEzEnS1l7NY+rwS/oxXfqBMeW3DX0iYYlAylYxr0zkCmWacEb7YhpePR8gNlI/MGaFHZm
9Mc4VRn03+jhXQzyBYgjg0qVVtDUc6QyYPV/Y7w8pUr81O9bBMWOkELFOmyLVvDJpZ5IctfgT9uZ
vktdNG0YzL0g+RmtsJetQY3wbzsTz9XucLeLKb4bIuIRJPskzwITxMf09tjbAXi5i22hNy4QWIGZ
e38h0RB0ILrhO2D0q7xdoc4OXpJCVXrYcAzF1+erpckWdXFS1EMz+AehgU+np1LbhOyKmHpDYd97
NKf4+Omu9Z4JLU9Y5eLnmfAwplKb2cS9K5q3W611tyiBQ0MTTbECDqjOMVFsiyIEli+6ObPrh8U3
bUu4cioEmGjofOFGI6xV5iammqevEOhNLA40aX1uAJgYX0u4gBCUGxtJxlCd7JfHLUdsvTLSB3Nj
xkR+PWIvCj1zLSf6rN/SP1TEHAtPrftjNjYI8Hmzr4IFJMm3X4kfnWDUExVuwR1PLUGSo0/LPffO
nz0wr1VjX2KS0nr8CPZp+hCVIDXcizNuGt7tWWFfD/rh4IC9B5vpEAJGaf3symhpTowKJIa3Av5a
C9OmQ+T9XTuFLYKHvNriv8Xqqjb1voZZPFs7817Z02nAVNBtjSfRZkNshxvqA4bIevEJc+FORkL8
mLr1MpcYd2HbXc7Mc/Gf0Cc91TZq+BF2axja7p3wcMLz2pVoUi3Olkmi48t+FV2UMwcelBj4EEZn
L3r3rwsFr/GrUybhJz5DR+TaF+dCX2Qm1mBFQ3wNI6rDPYGavHHSlGerJCskVW/R/MISxvj5y0Xm
Dj95DE8Jy3joplMh1f71ff8EGSJ0DyTa1k1whTEkwhpZVBVe/9JwE6KZQ238mBLatFXNJlPZG4F9
7HyRnzqypjffSNd+vz6cnwM69ElOF3qhlS7tIKqgJOIB1b7J4uJcCV/hZJ/jPeOiaWsJDKX9Q9vh
aOG2n8pD3B1f3OSSzrUcZVSpR/DVhyRexGsAYUNaGAzkXLFAFPXYqwFAEiZqklStS9Qslk9hwOOa
v8lKobjiiHGpa/KayqoY8Z3QdYyskP4JuVRDF45yI0cE0zi5tnmFhUy09kCqmOH+FMrQ4HVrNBmi
BUpVOhymB2GqJCRpK/QBBZXzHWkCC8ptNRMGKYGoz9xva2JeCoUZndUq4PRFVSfgawkPC159gC3p
W4qYOTQQScbn5g4nwXSv28wyTJv5b4/QV8MgkMuWcTmOlHwMAEVGgsMb5OU9mqGHsrXtl2pmY8v5
FmyXKEPvR75/iNv1I4IJfrt6eMd/2cTrmXIFkB6BUnOIQ06kFPCZPZAk6Q+oJmIQmbwV7uFgLY/9
7P81eODcTc11mQKJnNdfGwvVvZXuL5AqveT8+PfHWe3OWdF8ZMzXXI5sV8iKYXRk2tVxDY8AhTVb
6W+2BViwrM5fnf0J893WMaJ20wA5dvoHjSKq0fGpzpXsRyhgcVRfmwyaQXGg4TcLfysc2h2zlSnt
iqxU7tMrHlYCaq/4DEyW5kvJ05UfgKUfcSj3E+gXROFlljx18LA9e0R1IvA2WP8WP6MGnVlLFtrV
3Ktd7o4gOTKd6i1NIfjM0ftUdXQ442IQpxusjLNHXPzl6g1jS2VKiS0zuuDg87959pTBzF0wfDkw
zlhgj1ARQwq/8DI2X9suNY98GC8Gxm6oFn44iglqCB+CpanvcDTAo7zBMykTjUugc+NBmcXeM46g
bpI4uPbTSKFhBo1SHR3wdLAl9vehIdYQlw4Vhxzweobnsjq0yl0d0qzTejpQtwIpIkyZc6Wqcv3q
b4sQpTC2Oghk7EWSp0oD+Uw3guYYfHnYemt1x92DVPiEbf0d152eltd5C8IXJsQzuRvSA1zs4wIS
RYtg/iJX1QevkB5C8dHVdgw3p2DhkYIIEL601Zsxe/hivWoxjl/htAKvgx5ayKayopbQXx4HGeli
KIr6svsKe9pVxmV3L5bYITjQruHJRqupgAKaMveZVhbizM33lqs/jPguUPc6P682RUBm5bIAng05
eWneNzL1phkl4UUjORSpdvsG3lcXy0/WFwfSH3a6adL2MNEu9RgR8AmRF8Zbengv70mRqgHVygha
A/9nvnKhrMF9cpU5bdn7hIacQzWgfHK1XDGcMvLog7P3i6dLQYyZE/dHvpthGUamISjQaJj0CJsf
p4XzkN07bxoeBnKraocOIuWrJp3hGXNcBcctHfM2ZlLFzoC1WY7Jj+XR/kYjn4ymnufdfDdW2X3J
B5GQtt0nAh5SICvm72BRhCzC6qO2OqVSUyyYCMf3hGrdx5F2I7nJEcPFTvVzqaBgpzc2+cgjNWXt
3RUFbYrmNvAvQlMV19QbdvaNiy2JzTIXiCmzhhx7FbixMoaKCjkNFSuIzjXxRjqvNQx4OzqSaJ6o
5ViD91KJjjkR2lVAcvLGpHwi2Iy5xuAfgXmGCRZbUEvFEtAqWM0tfcbTA1P0pzuaicMFSeFen0F1
nT/6OqVvLPuzsEpylymUykkVa3zwHEe/1tCQZZtabDqMtbvh3h91xQ0zu1NuwOZZps5BOYjKLZO3
q0LRVlrfzqkaZRtqBqb1tRVsyZKWEZnP3mWQu6bLphjl2DrC0OQdo9sLO3H1lOSPr0sN7VhcqhVj
IXvUSAzp3U3NT0HbH8WKo+kXWykljqKNxfdW8Ii8Eb5FNLni4ea8xSygEqvkKJMIv7Bt9aPwGAA/
GDILmyZwPJ1K+TJ1VrzRuHpn+EoCsr/E/LihChYcjsgXpoHuJQ+gVkasLqNPOZNPypQ56j6iseYh
+PlRzizWzGblz7uiY1Xtc+24XusPwDWzVBzmQsacRjnmN7hbDbgKGpj4LJeJQcNuwI3yqIsypqxe
Q5uc93nN2S+HyZwq4yl5wj7qsmqhCosDy2flE960PxV5yh/1M895qvT44ntt+hsViWUq5l8CZK6H
DI+UtKEc2atDqga+ZLlPK/fioENQMkFHYD/4IVRF1CYAWA2NU7lYR+7f1Edg1Wq1hSzRd/dxmTPm
o5nr8smTfK43rL4AysttUinTsf//EWw75EYTOxdBrCDDRydGZwCVQUukq/KwtP595po8hwcC12VH
LMUJ5mBkEq/CHpgJ+K1TUWb2pkhD4ehfSOtrnF5sxrdbHOuzY4CTHiVnrEmYlOxe04HHssqeQ+jA
3ScHjWvLnsqzquif2rrzRr3OtKHAJbKN1Y4tITqWgihjyvYUzXfYLTrR2P3owIB/5SX5GobTBI0w
9nqlsif4iOpfTr8EjF54eAnK310HboHRhZqv/TLY2WQl4ExBNg1/Yq/Fk9LOSnrqARZEm/5XUY/P
KEvdGaJKjgoxnAR0hCrSRPefwaVrK2PN+HWdrPe+V1ewzk8cDcEWUOI8wuCxRV+bJmBk08w/ZwYC
ZRcBABWBw4WgjvDacvC4A2T3RiJ9UeT4b/0AOozouo7hA/iSbYmHUXO8mTFzHIWfxXoeec4Poh9c
UgEe2yA1zs08e6TIyIAEyGPP3fc56rUX3XxcMWup2CrG0IcAgvKOm0vI8dRHbD+7pKaOVcgqfARS
3VUffDnFY8V8IoKdWXunh3HpBr9cQiSY8jqLWUng0qZHkd0AAXrWCBlM23oi9zC2GN0KCaDrlgXZ
nse9S0zbpfnVj89B45C8+nmz0gHGDtubrU+tQlqZonYaZlayKI+TVPJFNrOFJ3di5w7wxHRjyKJu
+L3kH7UI1ux9hRqg5qvYgZ40X0MNjWgBRaajJvYwhORUErqZtYMzJzqKjXsS5OJkPl1jB8Cjd5h/
p69t6lrbvC/TD+H7zuqKNDoUkiZPRnnTvXzbs7ED4SGwY5dtSJlUMF3JdtsEEAAGc4GGJ4crap3K
2HVt15DWQBpG37CqAlYTEab+bZxd4OdqN42IgsvlnFd32htJfTNxC+mEwwdzLUclh/jksnpjOwkO
UL+Qp4uMQ32Hk6fwJvolKYD6I1HwprMKsQ/gAUYan7nyXLQ+kqBCfVFcpI8ri2DHsjxxg91F2jnH
janI/ZPRECh0UeuyaHTHMBHRyzO+SvWELJabn5LTcLgehMtHq/wxiuSiaiSqRZIGt4g4kI9lmu5/
Slvwem9HGlo1GCtfHYcXINo2bUe3e1wzXg6TeQntV5//8TvLH+ufX+6ZXvNVV4o0xpONOTiEjzam
Pxf/Nrhl1qz3g09tsJUR42/w+/NTr66TpLWyUWdjw/5Jv2XzBjCnxdrxo/MywL7yBAHgHEXXHa4/
RqHMjaVoU1HKFLAZ06YwURXfpVlceb6xdDjUuCGp6iIn8k5sr1WeWVkgozfxK/iIIU5myfJI30Ry
aU8kNUDfrbFl8qYIjIh0uFUAVslMSIJjm2giz+gRp7wVt6FMQuV8jnUloOAnu6ZG2rFBdn5kQPKS
QGW6OKGOPSXb18rNtTwPZ5oSPtfAPf3rPTQtWf1LOncUf9vPkKCQWrdrIFcGscQq+evoMLLy6IHn
8lvJ6cavZwrOYzBtPpiPBVdC2IjQDd5ZJ66Yzq3xMEuZKA1FPA2pm3oMOuJ40xPYUqZ1z0GWIWOG
TfxAoZNZ/MZMYPzGhS3rH7ns4ZVo7Sn7MvdeDS1j/j1EsmDlzBr26g8c8cIswtpQZEJhdgd6Clli
fcZXgZl2+ukrzVBlUBqVPszLVBSAycxqzS3EMJ6CeHMTcFtY7Tj8x80QsPkLxaCyN7YDnlP6ZVwZ
0qirjXwLn76KRHRpdxOmDapNa88IBoFdgUumcbCj9DF3rfy1F+yGJrSeIUwm8m5fqRXivB2XlHrb
XVnwadKcQtVVbzJPsNao81zchUKgZ2grKoJDDBR2roNiFqmnSRMIOow3kSU40singrg1Bqoj61zg
qOiVcRFw1NXl/CzpaawmwSjwkW8Lgg7xDmQdpHnMNoW6vZhd90sGQtyo8vvKD6l6GG1ugqeoUCt8
bU2KnA3VyfSYxfjhJVFj053JcVOZb4ZsO8arMkQ/+Zu9YtZmdKtHtFF1MLmFuQsOMZQ0XrkIQMdB
ulbit6fFL7RurZTqvtVkTRkThoPcRtsLk0PMmLU9lcBjlqVb2KOwq605lYdCn5DxmAn7C1TN/HVS
EoaHJ6latn+/W/0Is5++CptdUAINL4WEITNYPxvOzj8scF0TLdT35FpF/eqeBsIbrmw7KRW8s5Qp
o8k7ezVIIQzmZz9i1qYvA0CJ6yyX4bb79MLPlp3RXsIrnskO4DQbhLgDcL89zlTYShSUtoJRyiZ4
kW76Tb22c6Ky+OcjG1f0NLVA/ZoXK8aRmgPJ2OIURb2OeTvAci8E4iv736aDxfGe6CITXHHKl7su
Kwf4widKuDmVR7mumshkzEMfVBn/PuIch2jbte/5Bg4c+OGUzxHb3+rZgxh3xODR7l3SUAgZj2LJ
1LefCGVnazbLSJc426CeHiwvaWA+x2Yc9Y4GtTcslzxknE+3V5Mrk1yTaGiiQTpSW5Qzipli7fP4
fQPPLYxDmpDLLF4CZyyVcKyZ5i6iFxxOsdQJCX2zmYq/Hw8K2kdfTdU2Vdm7g74sKrNA8eOZKKIf
ZX2s3TNhJ+dWIyuB7rOSS2AbWwx+33n3oS9tPnk/b4DWvfzbqpytOMx8ebyuLMcTVTmjUx4v2BeP
w863+dx0JZdzA+9SMizzmYpF4LdpDSUBv25Ho/5p1iq8SJU7Rj6SK5G7nAcQwCn6/NxArC0npBsP
npCjQiENi2CQSUsr2gGva/Cj7/Yfe0l8k1CJbaS9CW/PBF/m8TZSN7TYhRCNxs+AKd6K6208V+iP
bYGZVIzLw9aKQGAFhShMzV1tyLRuIGCTl/nJXoPx1mkCpUklBca2j+qU+7dXykFWVHWNrbAmMAcT
JTEt/TIbOIk5HazUtteQKMpc72euvi9OeESCvYhrqaXGBrinyrUoTImJPiX4bBNDd0i6583Ju5AA
+aPBoT7qmtAgvC91siswcrlZBBKhN+tc+uR0lfKv1kx/RRaWg/Ld2EwV4E/qG2qGWpJhC3rprfo8
4uEtfAir7AqEyoDP8aG2LIqtqjWkYg+0XxSVW8WkyehT7xjpqp9tBr/ESRi4YdYWxFxAZQ3R50LK
5s+cT97HS7LOSgiYkWlO7uMWPNEjqV4/yvA/8UENoKjV4ZTb5K58p7IElboJtriTx6HXDAk7hLtV
FfVv0H7OIlhEFMcbn6F+ZX6MCONZyMlyq0rjOK6zIkkw47HuHeGWhHnhumN3PiPj5QPldZpt0M0s
UKus+Goeok5ohkqeDcf89ZxWCkR8lLQymF8tsXYv60UVVuHxG7lKyTmheIjSqge1A6GyhL494suL
nowsm/YEiuRcamFDBTmJzPbh15eFUfGDgaBfuaf5mDXcNnhHQ5KYhB645+68tqDPCPtLT7EVb3P5
+7+tE8GSbxxDSME48YdhMLAuHTAy0FHTX0eKuJ1MxnLCDloAQiA3Oy+pbt7v1ZomDa6/uLEJ9m9x
+EG3Cmp/fD0feCR7AiBPcwXSFDivDY32Nxlov9XTeVxb2t6JfbgfriOfl04lApvygg9KHlEWkFl0
F46/81bARJ+wcINqWfwnPxgLEpb+9eeYQJqogRckzXji0hrNlU7GoedpN0xgDA56XtOF/y/wMaGV
BXdhBxpUU7+OrWjwG7VttlWQaTrD688Se8T6F94XN/US/y9w6K9r15/6WrAs7R5Dcyhbil7bVSZK
pZh3OUu1/qKTU4jBeR6puC/ptX2lNU4ehc22FZFqmVE9T3KmrUgiKGXC4hXOfulRJrJZbRmIDDE3
MTEiJgGLk12AserD+t58MbJ9Sz2PnihhgiDNU5oaXmOzcJlb4uYHlyC3cNN7NANi1PU88PmOVjy0
7No4QzzOQ83u4xLdHDqBkKjJ9ntRVwwuTIpDfXp8Lf+O3GJbYS9A3+dxV3FlYEruJ+CYVjZJ2e2H
lQEoGdsk3D9ZwW3/5TjvfuQyeVlLxsda4wcQNleYHHXvjyIoW5TK6LcGNt6DLC67QCgJElG4wOj7
Z1YxNuoO9R/Gu8QXDqzdEZ5YH2ZnwNWbqKeiyDo+JO9Zj4Emqi3AiaUYmsUoWlm3dTiGH0Kjw13Y
2MDTCuXWqJf5YbBfa/FM4AfHd0uVLaV0oTaLqhMUoimnGdKxgASjZ6k1sVU0EFVXPQQ6XospVnOm
S7TdHXDzpONZnYquke3Kw+WILL/yITypyAruR5x6y+lUAy4OT/EWYZjeMC75hosaArHUcrsPJmx1
xdWuVxIzQxO+vOipNkLdnaKa5s+v6SfLgz6UfvQf7o2egzk5SWtUPoOiDPS1yJXdP+AzECNUkWOD
N+hmbHQqr629ryGe9Pb8ov+7euJLO3nXjGSZnwTAmgqfelTxlqTSUB4twNabb8UxjrUcIc96aHPf
wogGEgj0qq1O1MdUiLUCM4T8DZJjnWj/9CMghLuGz4ilaxJafguLmHwwCxYvpuupVPPJIsgchxti
eDUymfG8bUP8OMap/Z69RygqFX11cbIckd10D/3Ti56tDJUSTlJG+OGicnXFwn/0VXaH+Ebh4WKh
hdV/VgzuFfwqZZbwBHUrZ/Um6ZX9/9KtVtSXtHnZNQuu0Oe+MyGhMvEMEVZ0nNrnivm2mNn/uz4P
Hq90LFRMjKN7WmqAZqUy1onPue+63gIJLWSuoQcIo0j4so+k4UY2uTuDpa+b2CDPLGgJHFn6D4u4
6e57qwX+WSi2oGHPqG6uKCUd4I3jRhBKxH0CPkQY716VVApIomKNmtWSVPY2tITsKsJLelbVnE9b
8yX6KzxswJ0GnZRZsvvxHH9CqSYTmEsd5CrhIvaXzgLGYtWFrR6dhn/2IiQ57/lrE1Y3ThiMXyBk
FDaIR89BiG/6dZhXlgdsKG5okwTYCGsPbuYF25gYwJbg3UR2dEYeaWdF7S7IE7yCHAEsrjcP2c1C
LlSJBsVxJXDgI5Ji0Jqy32QKIKVNj44obbpd2Ex5jtojeDNWAxaoFGQarqS4xlgCBCKDc8r2zcH9
TVCiBWF0TPfZI76IqlAHNar8+Ccri52LwvFkNIysfgNwEsbuUkSSiV0R/uS3Kx1V9vUcc/VHAc3K
8dbQn0r75GaGSeQSbCwnA5hhlg7gXcTLMPm6xKMhyEngorIy8g8v1NLcqwRxEgx50SE5eVCwirzy
1ZBspvgEWT+lnyjDlMnSTNmnSufkiaMjVrQJ4+x2pbwS/E48qoZOUKOvp3grO/3MPaZXkGSXH+wK
jzRiyRsLMqxJRuYin0JkQQgvLdeLGmkr67/4GlKPiXwKOWkunILvUtrN18fhGCKNBXLfSuZ/VQGp
veGOul+2FVuFZBujPj2V9VN8COyetZx55/HH5/kb9I1ttbqlMR4riLVDPLJG8eLNr2W83Gy85TM1
6ucJs/hHHZ9u9vj3ked0Mm40nFun/d7QZBesPfyqvu5NG0//yDeVJ57HrQS1kQFZgRopl4sv5yIM
5HG5J9GvrO3Uj96E8iw/n04/H39iudEyEgoSOvh0JUtbb05nOdrbV1xUJqqsWK63HuJ6zy57l1Yr
BJTrn/jJkvuww7HR3PSNvwttc4RV1ZcBbWlP/QUgv3xLBiKOdKEBZ9CgDGHS659RxjA/U6wMtp2/
9pE7TFjnn53jMXOfFWJly/0+JEyu+EMXkSDGuSF3fcn05BLJNdBU8CdV7rju5yk/cEBY0b8YbwyI
I0wK5M4kU1H7IY9kZ1WTknWncLzN1otPy4fV6UznAPBl11kcN9ErT2OvCvlrtc2SjC+2mhyfgL98
SC3F1tT5SMFeEJjomG8I7SBbIbeuY30qAexd96tDNj061QgG3xeHCuvqtbqKk1/9lK4+bHxWhR3f
daffIWMjmQItUnGTwcWQcuas5PIUKg+ILk/BanoDfo4K/FGxU3BvRDjWaQzn3cv4ATjccu/OYLY3
qqu5I0v6I/nxfYCuxFMA1Y2kLvkRMyOEJ9cAAo26949CFZOYFrfV+1PwUYX3V9ZQBEtGcy7ipafi
H4FO3I6COwfWx725nF7YOYWXFxT2CPVQYIk61VHtjoHpvNCV69HJVaXcbnQbybmwXK06a9GhigTQ
WrukqhzSKBOuCZEj/iCUMzh2fm5Ncr9Zl6k1Dtyf7dce5B81wdsbxP65aMqd5YIeO/qCb23/IT2o
4s9feykibSsTwGwcNb0LVfKTBfI0+fN1S/FBrMNIvC8dnoSh5P/3yGItFozDdjpI66Lpyu44LRla
aKkW2sSOHGY6oEPQBib73xkA2PC3u2JC9IroNuO6GhL47JSb5SliVv8+UTSv/G1ORuJv985t/DHQ
5hyAhsH9WS2GUljpLZjgd9q1TiQmU5zFwzz8yR8T7MlZ/5vbKsEKrK1ncmSXaS8x6Z2sj/sVt0/w
Dcf+Sh4X1C1VxyuasmsKCPv6unGaAqsI04AqivXGOo+3kZpe4fREJGbaHF7U7FUpTIzQ46YEWwSZ
X1XjOeYgRxUChXUpmiZferDrkJy5/cn7kcc9s1yWfkwIkbPVN1aYnm4LUHdXA2+GZRGJfub+QFnj
VD4PP32Buc9IDRWASYOKBB4Dj4M5A7y222aZEsiZewjvA5Vi43nOJENRgOg+0EZ8c7HwAnoUSO/A
mrxzw/JER5YyeKKi8edmuDJxR/vcwFFYXezy4TobDp7/gDPYsBDF7ohky8Jq3ohUrL6142ur4uYv
UEFXNKBKUNsADgyPaWTiI0X6p2jS2t4FrGVqE8av/UUBlvQaj+fyfl3YaD7RY4ynexfELQz1s+pY
oIwtx3fHQ6jKtQG8fRuwdSdqWPWD853BqQoJQMyEky9ooDM+kmdJxWW9CG3QQwfzlU0ivgkbDZ1O
1d4+oOgQz95VwAfve4ejiWqeEv4KgPbePTrzgZ8qW6WmPqY1uGQJ4SaoB/sb9cqvtyqCa4mmoZAz
AthBraHkZ7JVSnbMtA6gEl2w2FUz9DWWAxMDx04FzNpBgTXJTZYFoYc11V5ehWp8Sc11GWhz/bHF
bMV41bHWtOU4KRvI9wuVdfeQbm9FZaTsXjjOLN9fBk40i3NL8g4zAezOC9cClLX4VXcewcJjVln1
meJkSm52JKkA2KvOmZeHi1duRBmM7W0LrhZ5LtE1mc5ueueR1yvuRBdb7Tur8ADd3mEgcs4hnpgF
gDJsroEgDjxdonfVslfs6roGQPmU+Q2V9thsetpbIOGQxsbzFYkyia8ChQ7VI76vy+YdxhC3IOc+
f8hO/SATUY2h3pXbZqmd9nB+SK3y2SNyMU1/xV+Q4RMbzecQupymYBtjxqIfJy6yx9C2I9a8t9ec
gRVuWxydg+ET55E7U4CjCkPA9O/mF8tz3fFnd/KQEDPJu5qWpXKPhMDRck1uZMTMUeli0h6Q94tA
HBK0R5ZJS9QzY9QkWa4cudwg/EnK6SwCtuIJ7C4LE9munboiLgJRquNxTovkSvkuWeiTBbYd/lU+
CrAEszlEU23slIeFEjBmCwyQf/SdbYL3M6bWZx1zdMs/MSF26uDWQCwIGtKqC+wYNg45POPjPx0S
44B1AFa/vHWjlMj6zK6bnVK335QyG2eUtZ+D2Y+t0D3uxAQ8JSgxr/ym8HxQGMIeoJORcnWI2dzr
NurqRIj84DdoRbEanWcLA6NgrPFnNAgEgbNxJfB2J2C8dBtrqSydmArDTiz9ue+FNtJ1vN0PkB85
NqLjZhgrui8I91lxRFFrH6h3KPE1iyBhwnESrhjPZ0mnX9cF+gEka0aW34J1uGu7RpcT2hvp8FHf
wHUnmhFbVi6BmlkBZpiB81t1d65OqqAVK1QAUUG44EyJmSG3yPqeMcDuF1TR/Yj5+zorrUljd4Cz
r8EiwFBcRPGdVU7wulFvdbc18/qGZ/rennVfpx4D0VX7yuDdFadoeW6r6WaIQEuntB79Zap80O4c
d/TFHYYl3KItwPyjN+GXQ5HVeXD2fxbQ00t8e83vTUJzdu64KTIPhVdujXBIksXsUihdbzAtn24a
qxsacKeIaBnTwN/ESjBc3RvH/lOoRSGkNeWH26aX8UpH3+nLdINgVrHW6iKmWYlIdWot3exS3bkr
Z4W1Gq2okKSej9k2OJIx9XSe0i7vYhF830qsukKLQgPqVy70Rkj5j4mrZfHRZIQoQz0xOyXhmmIr
i312TD917OupeQRaBJTTpXlJn4yNLQLbeWvVtuP8HtGjV5WRwpdJKLCVQLbd0DNKuQVYhgRrbqeJ
xfZUXAhxX8O3jkGzssZory7TCK6lxSw8LDrosUGDwwwVmkCoaEkaAoSRzZikwSdRIXOgG8PJ5f1A
RJ0Y5V9Yfv4/37CmtZn5r6Uwgu2cqBzqpNLu67hk62C1Us89Xi3XlMvnKtigkRt/3TZJ5HN2PDwp
//+ig+522cNW93Mtrdu6ax8rgkYTLQpOPr0Nq3hTxY0dI3vQ3PW0stOk1ZqFbVLsakcRMbvC8GWU
NvnbO6PogbzxMpw3foVmXOTN7hmvb2gK8/vnIbPmyQAMA95BDlt9+I5385HpyWNmpnoBubnXLg8E
HmS53HtMBq5N+umaVqauFOyMLfhoaPvtHv4FCAT+aJpE5vy5RPHtCJV812npgwFUUbkxetjlFD8R
sJZDzt7o2yMimCzViIyMOnIhumNxzYSlJAZrT+wFpkouq5arsBge6zrL2mKdpBBtFgz5Q9xYVGYZ
GaRhOCsb8USL/qs0F0hcICqx1ySFDX37+i2zgSM/OB4etpdfY/S/q3DNfM0HFwGE5GnCzvcCL/6t
yl2H/v4xzyNs5+0PZFpbeU+YMpNd4x4g56Sdu2xlkWMc3cf/noF0jwBEpY21ZgP+W4PCv8FyvpLr
sj/sm2AjAVfZlMGXTqV8AVcm+rvGQZfpOHUnyEnrms7BroMDG0+lYosuJq9dum+HrwviGNGJmSy9
nfuHsL9LCcVmUMcZpE8E02LfKi0EiY5S0jGNe0iCFPY88AB6D16J9bTJy5LFsOoXtKXntGJhwVWU
/qm2m3KlzYyY3M4F63dECMLxcN2uq+0Im9B3basUfkbBA0UrWo0oZ8zLSXadKwnbXU0LkFtRnmZN
y7m79+iXgXu6xbOpbnzz1N0cHzkwAVwGFNpOrkg66FWxqDxKB0T/1+jIwSkRRQ8does7fHzcWhHZ
5y3K4t46gXILAdo9W4SUXs5Q+320b0dy0eTaulIjKg8NC9wwPpVxvNR5xqKMBpe4xoQkF53Gi7M6
g+Wp1w4PXDagyDz+J42NoYdHKlfZq6FwDgSaUBlFelrAW/SdElUwUhBkVnnDcjq5tejb/YQJeVgU
yFtG5g27czPTNMuOiLDPituTVrqCvO8dGgAD0Z/vcAxyzF9P+u0ZFhfiDjDteZ64bjBfcQC4vRM9
on1uFH6+FMxM8OCx8QP7SJ1e2PSawQvjRyJbTweXLbQk+GB+Z8mzCQ5CqZVBN942IXukaqVYP+Nv
HCJ4zR/5C7AKCO8Y5LYzFoPNCuxfje6LZCXHMgK5/AHcuqqn2fnpqKFz5iNsZHMyfHASGV0W/6i4
sbP/glHxQU2UR7ns2PMddYFcxqOVful3xQctuOGdIglqB18mQodJqiXttn+FnsU+qnicSSzTX/M4
3NxXwdtP5LjRTt/dQgeQ2VkqOf8uvnH9HV7pRqOybHGYdRKoA+kGr33zQIiRy52d55qsqp9vBKAn
HSth6mJm8ZfSI5bqmhBQNZwHS+4DuKyUHBbqgEZoj4mazPzN8ttFPzGKP7h0XgpM2qjoRlikkalF
soiX9/UR+0/XvpSxs0N5ShtjH4QzrEKqkaWj6N+BsKPtFx1BBcYBYmHs3DgbOmPHX7mx/bN10XNl
M/+tyGsLi1viN8dpw7BzfoBTUQav9Hz9AHs18FQSpBZaVvEtRpM+pGwaOvFSZdLSYIgs1ac7zbmH
0LfQLHXZHdYzN5CV7diXxgFxf+tjvkUK9TG0r6BoOdzYIXFapBE7Il7i94S/uh2iYoFhDrRVBTMR
tQwZjm5Xa8MUdRoq/Hk6P/HZXmG9l2MhgH3cSpUjSLlpErPOxj8iUYILQbNmoNpWDPOxCvrVIQto
JM+0kh1A7xwEczI9F5odkAMxdCBuSG3AzgnQC9NSsrkJwcRRZXWYNXpZE7nvVbCP7H9CW7kDGfeP
9GbWSFKzKEW7JMpYFWTOj7TXr/uRhmhQnhcf+SHrmvjynHbMYfVQ+ZlV2tLn/aw6Yf/2ZpGRjYEH
h2FhP5Rgmm1uDDv+0x0jtQRV74Eyj+TAet+jsncQBWCL9FaeSRv8XZK8aMfxoQ44IIPQ5Q3AfKvT
PwoiBf01hIve0iLlbhCdKtZESW2KbEc1s1x7n9x/OiWLYks80iON0dTHqXATqXdgKjNRmaR/Yzw+
c5qcsbeqMiI0MEHBkRj2XCGUVeeswnqmYkI+L0L+2XwU7OdECpgb/EayPKYpiUa8FG5XEghSCa/K
psqXA5W3eLUG1fn4c1aCGOUaLh0mpc1EtclAJc++WEVCcjKWeaT9/YiXwfQfECHR1sDwADIa4Loz
5eJ8NAU6fm2fUzbZmAJFbF081FWS7cwjKQfqAYzbR/aeRyr/dxyqU/7puycGWe/9YcIq8m/U+GpP
5vY6cEijjIV4tC8wZ72yi9AWn/8ePAZ3C2QKzpjvFD+HqYZoZsaFXks7YPclY+vUIjTIZzi+x4AP
Q43qh7ppQ1MP/dd2Y2zFs4v6wvTNdt6Y1QLKdqfwkxI9nNb5wVSk65Mrya66EV+Cb2oSA9fYdSVs
86fO7FTSsA9O76l35P8r6mGjY95wB6r3swAuqxg1kx+WiDY/LB0zx6pWU7OUFFG0OzxCniGYKM5p
sMhP5S75X9sY0VuZl/SlgnOpfe731nqNGW4kcDi93mdJDfMDeiNo02vNgP97TrmP+1UzJyrv6VvQ
pJ04kTEhIqyTUIoWdwidj/VI0UheYK6Zm9ADmOvCSOBTxVh03GYBy4Xw5BqaAzTSBLvZlI40uVKx
isHDTLpjiHTO1qqqpqwAXmbE+04kC0aTkCwxq1xm+j3utw2V4vVYUmTUo1E793+wtdxke2u6aT17
Qgh9ArYxdGZCuYWFuVhD2m34Fpg/gYUPnoML+24N/fjb9dN1vSJXaObrLbAlA5ryUaFVwqgRljS2
D5XmFdZFlpGKdfxplfZ46Q4VOnaKHMgJ/tRaJDKcTXSEQB3kSfYmyqdYdp82wEhWfPqAswX0N5QW
2mDdv5bWCZ+PX4VYIiDndM/kG9X+glNZTOHQJ8OaM/SbuBAgxdrbMylbtN5ljSIglfr+S3in8SAJ
18wv21/kopED9+neUji93LS5CLLJFTIHTD5pWxzLT0AaXDfm0Duk64ircPgWDVpxPEiZExEWvqxw
HAJ5sg0ZSolJusuwtQryCyngdka4c/E17S9FhRHKjvS7luD2/TxUI87DW6b5RmOBbuH5kIcU73nD
NEFBdlxG8jItb+ieA9azO30Hv8kl2r7VOSSq8kgQqkIaYqrE5jq88BT+POCGHgyCPdCIHbNy0D8G
GG+I4giS0OqCY5AOCAylZKBCgCSoD9YAVR/ev/oSYFhbcgmZ8yXvGhJaZvg49YF1vvOGLE1v0Z9O
L0PvxWpy8F1u/vfeyLVNyqTmKrogjOMIIjfTg4TAQ5oIbb5Kq4lpwCBzcxPkVv1Ajfnwcod9eMQY
poJdCuXNbsMp2MlCAXFGIwZW+HDCZToiRgnEopNF8cDlaYwQdQA=
`pragma protect end_protected
