`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfinaGAYB962HBP0i41sZUp9txhpkbUCYzQiJ2+z9BHRMx5Hotgvc22Nw
2jWc74J97lNTGv0S+oePpCKfLuz+HBorVi8a5VGZCBefLOlXkVCpI6erG7YAzaL6itbzpkTfeabW
WZBKRwttRfeXhYmF34BDxsoDdvFhBVeGdFqSK1eqWCluiFn2McQyBA80liXbuSjrUuISKKHlG9YE
3/Jk2uwqptPHVJmZb6pMLWlWh0Zq8aBs4c1d72nJf8JLASBrmQ/hvy/IJ18JrO+tC6cCaylS6Eux
xpzaS9H+gLp1WOEGn6yTYhfhQ7khHVtbMTqnwIJqYOcHL5K7Jx0gRSFD+6y506+vj8gj3TBMCcYd
qsrdprFPPj1pQTWLnNKqEO8FmbmDN91Kb5lAxlgggHMDa0BUNTThHYQU9RBhhuCwhf7tQRDVVF6i
ziUGzN1faEoRAOKWUxBLkglwyotoOaFYRBnq2Mkskv76ciGb2SDiFeElOuylSUfqNPH9BYo9e7he
5H79FOGCf8ZUCjG80RTXB19QG+qggOZqGUcniImEg8hWfn9wYgadO9F/hRrb6j7IewdwJW+MkoNq
B22FTSS5xgRaqYyDFuR4g/gNimFzqSQOviV2SOeSJDwkdN3zba2FOytCnfD905+cCLco/TP4QRSb
QfzO3fTT/9Sv9FJgsvM+NeXFwU8qSIdVekpzKuHl6Qu+WH9k342qmHSe0OBcqKW7rI3BFuja9qvh
ebh1vqGCMR++t+B6UJQxGbFVWHdlwtZXzmGn+bWjuNSxL9Ibq5HhozAw/Cn/3vQINYln0GN6/aCc
206aEfDUHnvp+d8yFspExwugA9248Uyv+U5PZ5dNJiMjg+KSSoNU9HTK6krPJAhr5bRxBiYrwfMy
4z5KQJtufoEFV4R6pWwVQ/8DDSFtmoc/HykYtc6UVXEjy0BM8RZrj1i5AxCifIoSrzvufi2r/wRR
vPqZ/394MLP8x36NOqrVpjA07S5sVt3c6wuLUz/DwXhuFKOqT6zVg+q4hAzL5hCBjrjX3obfutit
ysb4jYjy8dE/wLxrjwzYxorCJQ7ZxBgOCzhBUWWrbx439EXk5vmAuv6KLbXbMcPF6qsL0/s7OmGy
D3zAy3j5JQGc1SzCTun2ur1NdAXAIsmef6i8MySNnbOIeKtKgWgsYdiZZS1EuZf22b1XgB5hjzBQ
Ly68cLqPqOiuJ7VZ5qRIhnoK3eUlqmtgFQqYYgChhoeEA8Hetez1xqCys+lcdOEsUsB1Auacslne
U3CRParFPxQ2pAwXCI6u+Bm13Q/ZtMydkKspJ3Iki49M17nqKHEBGhH12rvz8LQ6B/o4wEX48Do+
SG5linTe5SKvqjHB/AdbcbD9odBboOVk8s34gyLCn59PU5zXdciMd0VagpBFvVncDPoVPHloq+l4
MIosOq8mYKYOCHlkU2EpXlzd4XkF4dz86kUyuofGLRkJEe7WgQ9naFPUDRr4Ahe44tNKyxya1ms/
bqbSnXaxjmj6SJsjDtfWzRkdvMZ0nC09B21bHmQLM8PQvQbpEg8ULb/gBlhN68uiabsF26JMUcQx
+zFGj8Hp1G+cvy8ns78HROg/1ff0Xygr9bQZM9GUfaG70ih3HOsRhxcolo3hAbSKE+LY/C7HW0wj
YTu2pIBwwfqNB7u09D6rQcp1jxHv2IXFuv6rXzf+2swqMLYcfyq1AjK2hMHa/XD2v0cc/pSTaISs
rl1ye0YbWoM6tqJDmUKpj3pqvbCHToeIdiV/ojdoPnHVY4l0SySouVyKpdB9alMybY+m7LDontAf
uf23OaafC0XaM6lQESeV9UZOdavHWGkONxlgPN+MAf/YiQMhww40iSR3qEl0RghBjuEKEkOxEDUE
Zfhu4ikgZGiPRHKs8qawlWHFnuD9u1QI0Nh7wbffKEzqx0KoHZIue/g+cCY227Utk/VWI49DSndp
1czEt2O/SqCrhAqUyxbwqvzNJ9vEVxbm5YPxWGV2veKBt5MwDgu9FRNFoM/ThsZZ/PAR7g6jNPZW
SZxvSKuaavRtC8klqYt6S3+1ZltJvkxg8RZlbWz0M5Toke2T6FAoOrsV+S1DGz7e+Ixn8jCrs/hl
UxSPGfr7TAWzqjV6D9bhyyWBn/Yevka9WippY5FPxk41s77MM+LLIfTKVDMQivSsZX6wWKqloUKz
L2kQj2bGCzGqOmQbxFZD31VW0pKAf9JrrjXGus9XGs9Mysm/OapppyOL2NQHU40s8JsKVyJxhEz8
/vVzHjEM6pWODfkO1fZvr2NQR0SGcMDzhUfzY+76Log8u5ATBGALSmSL5TTMMNP52yLVrqb2Dp4a
Pm0PeKkusWmcRpoSE9NMWLLYAP8kA6SLfblpQvrLc/mSEnPeA4qxs+GErtNkZmmjlxih+EKELHty
t8xlMppTbQT//5lzN8tSSQOD4aVECJrBhRlxqQg12P3EJsbSzzvC6QVs1DSX2YJ2qNK5os7RIOnW
1igLgZDoRiP/PAifwyKgYH31LzNP6c7/C/YayrVGjqlUXBskMuMca0AY/MojJjS4IZKj7mDJOR+l
YCoPSWZ72fTVVww8rlwkTSlTsR4HnVpONwoz+q/u+sLg6+g6cVR8fU8MfhRMM0Kk8tvBhZO036GN
uIVEcsPYLR9/AzN3w6yt7H/qKycVRIdOAmQdpAHa/zGCo3/m2imosoiNpRO6OrbCbBTYbaRyWbi+
6AbONkp9+dMs1mqKWm19UxVOyG6qXECt3cqBsAcJyz9u6zHkEkDF2d9t6AufPoPsZr1Al4ZrQUU/
rYZPigeJtglOE/Ux8H8Xixr8kv5rPbZBJiPl6uL44AyVMw1YCvOs1FMcNYlKk3uvbDiSk3j7Rr+J
V+19ncjwQU2ENaabB/V25ELMLXO1NTOPnwlVkos+zgoDO9rMUzVtzCPLQ6J9nvhkVO7ucLmBveVf
PeV/cK4TowwCOg4aD2kwSxmwNXVpw4LsxlnyYmQgR6pdth7/RyJkLAKzyXPbkBlJOQ4mBBXG0Ido
8YGzhc5WuTdy3Yj4VhEjJXH82RWOrS9vdX7iooQdpIc6pOI+RVYYmvH4eliTagLPDEmPzVpHgse5
dZ7DebgAOgzX7kJdWnEh8q9neq0NBZrGcUikliXceganaN05s4F4kgiXdbY0I6QSRCtneIm8Ue7f
1ru20AOG+gbWS38xtafo8jiG9SVTUAvp0E8Pv7/uzaohWIar1h6VuGbBn2b2dj+xOI0FJeOJymfM
WICdsuAaUwfBdgQjBrIRidFL3H+h5HjymLzWFcrllZrazLY6QJ9tN1WvuJgjC7KlKaG8YFDQ3lIw
SjfyQh9PBcklZXrFDLRW84wMoKB1nyIOwc6kqL1aBMonPp8hYHIuaZSGWY7/Q6UhAtSbomVFkpGy
ikgY+3BW9CNMHS/KwZ8omQtCNJUAHPZieyep2SwnoHxN7qrUVrK1LgXkwvGrlTJ6eT3QHNjptfO2
zPlBtQf/qPUtbNZ9MdwRjfJ57deKs4x0hNmDeNdjoGlgZT+Ns9w6naS//vBrugac6MabJQS1SMpx
fA41ZzwWe27Q4GlqtHQqipGvY6EOOj2/uoJbqayrWILHmo2s2bdu7iJhVkYDqp1bHgQYVxn6+Iou
SOT/8CnspVZvK2X9UTuQ5TXwyffl/Uv+cHdyRUpmJxca0GokZqr7UkKnxGssy2a6YDtHT+DLlarJ
9lqn4dOYdD5eHOyCFOpbrhZhHZr2v7Bp1F8H0qb3PHEA+9Q6u+8iHQkFMk1AzPdHz93k46bSd1xJ
5oValX96uF+06lzLstYJhXUdgnvegP3ng6sxUYW4jeshDwS5MJsOM1/xehpPflSqJa86/jBfrzBj
Ay8eqIxwqv26xZKs2smaZ4uFH9tBE4M6z/F3r+s4t7bz0lR0qQrcDxPU9nBjZ2RkTOy6rxkCJ3OP
xb85JKbWbTpUWi4vyLiYT7RnLbMgV1HvdnU6hYjGET22A/LcRCcWnE7EPIJtZNYnvU4EafPXgh2O
KmwZ656XbK7a9STafHZcJ47dmyx2+qKx0mI1p3jvSLYQqCAVJFVdxqujY6o4MhxMm1NtOWhwrLNQ
YHq0Ub46CtpQXSOncPdWVAdNOanztpG38+sv+pn51F2quvxyp0kUxHdCseKU3VlrhhQlFxxYlpgz
HYrthSztVLjX2CNJkJ8Es3tOQRwKm39nVLaQYmVocEU8xgEj1NMEUAOU0tdIjU3gr+h3oIxZFunA
LeCxvaoDKxCfZwqGSC5oI4lif0lFz4qUZZS/FLcXJ2+D7qbqr6l7ruqIep3iMlmxXjRedmTlsqTh
N8l9pABrR5n5a5YoHFaTzouiSvKChVrpZR61kI0j6bXqboTJAZa3DbZhjPAIq8phDAVpk6Gi2wlG
OjkIwjsgGE5HVqJ9Jtrx1ecbY0nrCjMbfFI068nzPmrRl6P6Gc/OFrBby5IhpzyIsYfrR47l9/Bq
PS7OtOLLw8TEHEtiZZzzqwvu4w1Hd/DJVl0Y9yHuAYLlfLf18bBA0D6umwFz+qbKV8gNqT89QH/w
2djaLGUkNdooSWs0GJQCuzMmfaluTS+l9wE2eomMe06CvWsw+eMEluX/8WQwdSHA4E/a294G3dO5
6sGxxIT2MaZ12qp8gEWAwEOr4MmtAWLEEv+XbOSZhiuhh5AuY9dhYsxevdyT1lIw688ozjvoGd1Q
Gg4Qb33SsXlGlZg/Gx/B1MVQ+tYByo8Et0wbmCFlre+vJSjNYKbbjtchKPyPbtHfkLICVgS921Np
XRGJKkaJnUMmYAGYyb0VRNcyovubF2y6reNKqKn8PjGcU2gew5bEYD8vY5LCatETPY2c54vMr8ip
YrSDRpAcz0Af8LuFY5T4kHUyQpKbrpnVDO+YiZvkB+cjuqhwL4mljCJE9SOVtSZ1WNti+l+unFI5
kQYL4AigcvwBIjGqQJArFjy/4esNdiDa4BdIlNdBkDQoQn+EYst+3tcq80wmpbTsoXbUOyzYTDdr
iOYSb0RTCqyWD69le0S15Y/MeutD9MDgIzgcQM7S1nVlhMx5yRilFRTHW+0WgMnYq7MPhODNQ2xN
CCjwp4QOA67WpCU2bl9zEfHXXx4SX2L3XdR80Lu+ieeoL+pjctqjK+m85UXesQB/QWL0UkNFoNM8
P5uJsoVyQrjxqHSzED/+NgljxZwhWjZXhSspePoAk4ww6laL/41G1b0qMrNjwwayipqAtggBO9Tx
9vH+huh79fnAnaeX4o6LzgJBhCp7fyAb4m5jgP5WOUv5XetnjbpLeHZ2/5htwdZmxX6LCeg+zc0g
V5C1WjK/AKVGL4VKzNq3NqIGfXVaT5IGLAE/km/W1peC3L9BDXXf+Y9pEErOUuloeGRJL4994FGT
uU8Xf0SwOb7GrVRovgXTfSKeauTz2GsHdmWpF4IpHGnoouAroSGIPtaY2kxwMhzaoV2hSbKxBw3r
MsgCOqEtlRzKkSdgn2+20OgVLMQ9ZI70vSaLf5TkJWEtIjYNODgX2sZSlneimVVehMCvl3C4Sq40
FLH8BExwwr64VQDrfvPuPHz+B4BvHPaKy9HpXdUGv1HEqgwzZJmdSCebswiWSZTijHgBHQ4DOuUX
KniMXjgR5Y2oqvtTzzd2dSCqOxuby9WhGVysR6pZXzbS9cKqFvdR7Cx6sY+h+x5Oz7nf0eq/9dtb
V5lpykUxHo8NW+QUdIwEPgfBSwvcwiFAnbHcfcxlhYOWepldUDy5pSIkCZI4E8kHZu8FOCWyRagN
zBq/salrk+lSdGmx20xSxcA9qQmRss1vw97HdW6+SK9sX5qIpVR8f7dwbix3c0ri4i/n4PtWdUFj
PY9y5sVhnRGVKVDdYWPqrpLq4/JaLg3UnU3v/u94xor/cQLEZ6peqrMCXuaDAmRBYqiI4gPohxY8
4kWrBlicgk5WPbS28PUJd9KjDGA5iks/xs1lRmxOoNrWU3lKWZ9BJAEzLnCy+FgRMSjWJGKIIYqp
BG4Qwajh/5IT4yfGyLxZZnF+HBubUcf/Q3j62Uky/gdFxc8McPlstf0Xm1zeo7icPODTWlDwPZGI
Zb9HqiRhCoIS39mLLiyL3kBnUospQySYOjlof6ToDk7dSzdncgMTMRxVxWzYxin1xA2dk03rJcxb
ML16SC6EMDI/f7o4fI07k7iF70zOBySFubNRlt/6gUayjFVxAXanS9vKWh1thXS04v4GkY9cJIGA
+GKRmStMqb/BoSDmkIA6p+SCZB+dynWIDm/vDysyvwiMwZyRHnv7EwwAjxqf5gDinQOD0RkU6kjy
s/lmy6W+vQuGtLEVNmZfH4uYt63rMzkEYjd0KKUr+/u6598FLeoHW3mue+PRxFks23uwKGBbmHNW
+slpw9uMp2MUlXHXbdrq/6DBVWKsq9hZQcKkKijH2WpA6s+eTIIjE+fKaI4mrqCiq6dRtHRiGhqo
hcrsyS5Pj0cZbZeJMCtKlCVw8a8somd67C3RQO2qF44NDuQPpIlQuD1JnHGswZSTSfMyXBKKH6+Y
9aYZpxh3yVl/ILr4pli2Mum7CWz7/U9/JXKPMUejy7gqRmSHbYj4E8L0I0pk3sIOqblxBEHaivKZ
sdtC/KBra1IgZsM9wlcbAm8lTgq7AOjfhaY5SuuPYCK7wA1TdO23D2vCocfwf/WW2IU3i6jPpNDH
qVzUwFLmDB2P/XyY3kNw2jMnQlDMwSFDUWEbynI7K6ZkgbGzkC57xNKMsa1RXzP0GJHkoTDcHEyL
di+Z4xB9Z468r599LlAPs2Xh8Sgssl8thQPcNwpOilDqD1yMfqokLGI0a2vycJKWpc+X4x5PgAPx
TJmPi6isD1RWKZBXE6XZxbZF7KtMCz6KeFDLb8ADgz3FfdIkngOsyIZTALzS2/zuVbWLGQcr9dda
BMsSYcJOMDUJKIgIT/vWuf8oGjJpRQFRxyfpzXyMXm8BsxKbYxYm+au6mIPNWmHxhfMJz+MNYujx
RIQnLSiaGrlIgD/XNUmgAQSsVvazD3nFPhNANmb8ljqZMgrcyqx7MAuDroBFG59UearcNofBXrq5
rhx5wb2Mql3Ldr3fulw2qoS25PUldm/igP8gJ2WlkDRn/nws71yIMuObmaAzUjUpRWiFKipQwkkK
k3mLOp0sD4722VEmGM0zoFdwvUKy6d/e6OwiknPty2eIUouTt49rtNPl1t6uqi9Ik5HjjwiVvqd8
8cxnQh/GZYNNLWg8PJVycArRGpuHnuLVMK5P+FWx1f7FMLYHL5aw0rGu/x3IogsJNxS/mG+fqpzd
0nXseie0j3jd80dPPGCY2Uv/kiQfNBm9Rlt2ZFSz9J0Kx7tonpLc2HVc7QLpaxAsZ5xXc1kcyW5Q
TUTsFezUUA/8qTx/1yuHpbaDj62U8WDqeEMCOI3+fXoa/TD849Gc+OLr/HDjceu9m/V6uXOSbFKv
wgaIy6+y5C8PuW8aAXg589RfSe6+P45hBMq8ZpOG0S/8waQBmKcXjT0Tk81nld/KR+JEve/LIe5O
FOoUzvE=
`pragma protect end_protected
