/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52288)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9TEKvxviUK4sHLatfEzf5YrF3rxe02uY+s9LNGkhIfAD51uzxCRYY1+h
Y0teZiDKCvJxqz+/ihHE4Eva6BR2CTLYBMQXwhoIc6Y8oI0yzVSc23ESgnHPlXc4sbuFdwxVTnsV
ybYQG38U1SgpFNTn8T8AMcmp1EdBUnqNMxbDv7ehiN19Ld5zRanGYgmk2enR+UmUmzTZSvJdCyEz
IaUefIjChqVEHkXcwR4ONScM4wFGlB7+Hb+2TBLDObf/Ks0tejyJPijn/Wg6r77+oiVJA8ZiI4fr
vYphognsw0hGkDgPAokpdqhg8TN9uy+LlVzW03dYav6ViKiwj3PZ6e/zlXdK/zAcXaaNyhUa33U3
FvmktjFeK2JzxwAAv1kL5MPIKcdxHEepEHT4QV9bgcR8OwCOP44L6y/ZRWS/KBd+UDPY+VQnEhBy
YyQgy4k3Rvx/04krNg6rphNMlnCwP//LDbpW9vtbgfHrIhfJCoD7Gqpnd7S4qf+LTNueujM7pTnz
J3SQFlv7WpuB/cn05sq4uNGIIBL2Qw9XYy3Pfv7079lpbBoYAwjJDSMOMqKnVqJMcdIFWJgNTVH2
3RofQyOKHTiboQc7u5tm3X0+0pN/u9Uwq9CIvK8sFFSlJWNaviSF3VrF8g5MGFA0LO57njhoKEie
VE1b9924nn4qrEICVpF7V4chRqjLfX5/w25obOooTNwl0iYpDBv/fXrzUUc52WU8hU/Shf/p66cr
ddYvFiik+WFXpSqdpPcydjzzfZgWpQfsv6p0d3fMxLSkdkoAO6EVAde0jNxwSzUQAKD4F7Yw+Ygr
CapDgPdsk6yWdYNEN8cVL9qMLYijnIZ9fXzcwrFBqK7fuBC+Cw7m9+YLuNVvW+haEIIBt9t4TgWk
eXiA6wV+rR2nSJezjRxA0KIieH0TyVDLdktxHBcfKqdN25oYUFR+KaV5OuG81GABbaS8JcDTaWXq
XDEbAScvyUByl8IAbVhz9WHqzgb3o0omk+ZcglSApvGq7zeusaDFVHnlZF+EqoXaVjiKfLZW4FcQ
7KmymCxeQNIQ48RhWLA5ZvvHTVxzg4T6yDU0DgfueuZdjUM/uexwJfEyWP1XkDNbXZAV6W8V5x5y
kjJEqYWn3Hja2nCkSqAQqc+bx4XMt75JmyQaIGklKEwIkPUVVYQ5C11bxcpKPzyhN/fblK1VkWgG
qd0oab++cGUsMVoubkhW3J62y5ENy4ryvyQ1DU1EMDmb+MQuMj6k67CsztMOeJ2Qfn9ZrZui0T5M
g8Kx2K6cp45qO+fDeavCXpJV1055ZXnyy4nzTL8rrAX8mzbZgIHEm39A7vp+hOSz98HzAoQdiPIY
EO4uEMl0v233zJORohwMiXK+ZApqtIakc4HrGRlRrw2ljI3EbkJnbOufOpwNHS1pYdX11knYLRD3
AWmk9RYj/oO6t1rzuwct58GoVJV3L4aTgJHPFPcY/ZJRR1mwhimsovMBiW9Ni+gGmsvAfwRmgUP0
Y4VcEsc+O2zkFFLJi/6W9mfHEYW1Js69B5AD4AyzJl54yHU6XZyIBI3UcsXfLdqd8tO1JTXzx+6f
GBah9LdlTeyFEhJpsQWeSL4FnYx19Hvb5tF5CTw/uDNnKVd0z4STZikEJ6oxsbl9xTU7uDtIgGTj
WvKG9KwNMZffo2zybeci2Z/39puqcAbRrls7D/0Q4PHz8XrluJYAc9jaIVqYXfNIWD7Dg9I1ariz
D8GoI1WN2XF7Z5915NSnKPmvRNAWfkdGoskMHPyUwNinwlOg+MXhDnk4CLChKR35GqC6WnPqVjSS
Nz/oXaykWO2t/kpuBPzLzZPOnts8e5mKjPacM9Be6ydHPYygy8R7l169meVOuPK+v6dGWPm60cYW
/CnnbhEwVR4S2zOz4SIWhwzb3WEvEagGsakY2wXfwmPP5qAzKmu8Ht+AJ937/eA9EddK/hjMi2C5
JF4ax13edbsOZcnhykkP9wolQgMBphaugFh4fqZ1KGxfUfYfSjHRl7b7ZMMN9QyV3VjAniedb9Cr
xUb60PlzYYTPLuCJgKdtUH/2iYaAIE7rnhYUyMNFAvNkkKzEGK0C2Ue2kcpMDjtK13/uXMFu8ODM
R0vSpcANEx+kJdB5vl9obwMN13mu0SfmqBbKkTeTGKbRy+57imyVCteCWEizQr+CMYJdSfA7vwcE
NR/I7Mo8ks8yidTIHnptFtQ1SidHmnikOlPlKtEpPvo9/y9Ryz8/8Mp9ZR+3ghJMGiiZe5L5cm7b
kNy39HDU+MZ5oVuYQNZcaOEaLhMIxSVi3K14FzIhoSyrzMEuWuP7uegs1d/AOJ7xK0nqWqu+MVpO
RUnlZUr3kKOjnycOlh0qcLeSvS2RWNxhpKAXYMR4vz9BuP9reqeWSMBfM9ub0kcBGh4yXfjbm55I
LVSPrrJ0u3/r+pMTqVkcSW2wwzFkJ7N3V50sqSeUciguGeq+eiDsy1KIL/Ar+P4hAey10DHpBPmG
bl7lIIGwbs4BMJIE/l0Iwmwg3JUeXZWOLPR9CF6WSt/6mbN5CsdmdHUcJ1Hb3Wa+leLngKaK5wZA
ah1iiLzuF9lvl4LCKJNbMIgJgzEUZ5iDmZw52oxGEmBNQbjNLejquWjsll4uq8SHyAgYywqKpzAd
bdiGDHo0je8Q71ApbLAbtUfyGHzWieeGQcSoZpOuQOY/O9UJNR4jA5bvCPnAM6ad9UdqTxWwngvi
8+yUhxvE9LYc0G2yrVEyNBwgjopN/bzl4lk0Tl7mnR3vds1Ai4JbJagNHLB4vCtsD4oCOYkOFvI3
nVzR3ySWKKnmyy0uAWc2/S2jCBnouOnUJWVvCZNmvluMO89HkG4ixbiU2sV9ILp1YOTcOiRszgwC
wAS8Akki6kNferT6ozC6IM6VKplru59UyVOISF+2CFU4sgj/pCAZD+8o1Y+Bs98A97Gl5ovvXJ/M
ZcEMnTW53L850HHl7avO/ES1qMtZaX1Oca8x6HarLcURFLvLnhGPRFT/Bxa1/2ibjfSeoiMp4HwI
/z4BwmWl9gymNf78j3ziDDRe3jIGoHYCvsUuGjfGW+VjEdN0t5+7wgIViXI/pfeLvkD1NAEcDRNk
PAlfQltKBlUU3MukRHaNdnBppExwbw2R2XbJyKlExNAQs1G90aiUW4ZU6h7E6TH8icUdSlNO23H6
ad/oADESV7c/d7O8TWD0jhEiedsMkSL7J2AL9IveoMn976zdRGwU/xUjss0h/keIIP5Ky/uL2TLY
0yJI0Y+ueUXLRfytBqDnkOU/QcJdwV8lViervSsEkSTWzmikY7B1G+e0ftSJN7pVhdxaXFRaEsyD
DXkTzcXsvxD8P/nYiperD4j2pdG6l305AGVbheg+MhBOrqpFfdnaPZ9Vey0531TaWqRZZnfkJ2Dr
uQyNZdZPAERSg4JVbhq1OkWsgXEpdN0nuTzI0lF0wMNQLM2dw5F4oOIZDGwZhyFcXf+bshEW4CTr
fXklRjkyPj2e5BD/RoUGlnQgoW4HrmDiK9igOoygxw0zaVOOyJqs6YAUR38VsATS2MK8DhER3N5N
vf0hxHHkUVJSCz855E1Ef14UutRM1kh3Xcvfx4VrgPd/dlHskqS38Wc5gTqDyVFtPfN3ygfv2Esx
GhdHGntuC3Nr0RIaI27KvnVtFd2yRR/hdjtGagMP8Lrmcz36QL74SSCZrc2Xc6W5kdIDcMAVTxwD
EgnAJKFTVgOemutb3zxQWWaxpCjykVYltvD6WAoky9PCd+iNq4ZIftCGaBSIRfF0lrRN3qTFnzcz
h72PjNOhqsjYFuQWH6x4pW/fwg8gCdQhDxOSJBy8RJRyDkYSG9G3cZn4OxNGZ3dSJIxyV0dCPiZN
ZmcWauUP+hj0Q2leT8m9ESkheJRH9iuCXNA0ANoW9UgUEQedsIdH3xapBeM/cdPisMZsyDkkHo0N
ZZa49gVpv7oGww2uBabaiD9r8ejw5k4u/5AM2nlCuoKd/o+E3gj5xlIQIb1rzwStoXMQ0vJx/yUw
fH7L+S3gYkPAPbhDuoI/9pUjcspUAANF3lPbScS1wcszeaKdLovYq9niGrj+Z0EYINfnDj0ORvgq
4TUwI4r+ei9ZKkPm8r/ADflfQYYlSX+Pr2jfsCpEFfVbtqWu0qbExsLtEy7fhovbezJl/wb7vKgn
i12X+Wc+q2pghcyHquyBAbjrccECs9+tiXsh7Sgf7ecO45EnZNGycutUcUvVyc307yVl9c2xMtBS
BFYDMxvdHLd7S3UtL4eOrcYT2fLe2LKWEwOEvmYYep3lw0DQlEF/wMZNKchffEiLOnozmGrwo/a/
P24976aRf/tQnqmVKaqcGpD6jIlby8SNYkAhQBVsjxsXlrAIMqFMt0j+2OvG08+aehxqknaOaCmq
B2j4Qai/SXiHiB79dOTvmXDS+t8HzDNosM2NTz9oG7qrgKdwzNSj/gT6ZrM0gxpPm0Mz0pKzC7QH
NWG9cQltfDcVhCA47dcP/MbXzT5RUlW63iyQYcCxQZsFQXEBcSIf5zkS02Vbjhs5P7RzLAPejinj
h/4FRYtuqifGJJgXqhxY3im6tuPWpErTqh2dXeubKswkPwgL8VDRbc1lsMevptDFeVmLk9Wc54al
K5GsyU5gifnt7oM+WYTaWesL0hQAcu8VXSu+I6dIWRz7XpyF2a1w+MdR8sz2qNgMqIejOBmx5sg0
wmD9LIQ+vj+129ktIwVxLxh+yz1DHyKtqNtRlEBUh8GcxGWe98Yc8TqaRnzwNl8sVIq+r4pTsU2E
sQiAmjNQFo/MwYPS3vuVteR3ie74r0ywEmw4ukwBXJ+HFdh9k6qoyRFyxwqIomrLXO3p0FAUCKBA
ejiyC1F7ynKpsvzpZeARgtr1qxYb4Ov9wGyWE+dWMF6DLuzqIbFxn3hJ+8MZWJWTuY6/VWTK2/3W
MQFMBNUkD0ycHjEWY8zq+N3rifL0LRhKXZY25Ppmx1+LGGa9Rt5LDwepweOB/nqiaXZ58FXfTLLQ
Bn8w2SyZLg9EYIJNpOAr2fFUB9a0AV3Qc/8kjwsW/rYNINO1Ix1iF8jyPRYUMdNqIrdB1XcPiqfW
zVFkqD/8oQqR6i+zW6jxOF4DfxTbyGxYvT5nqHL6TlRPASlSaolmfiaJ7hVwRKJ0gPXd+bT81XhP
XUy2GD1EBuyh+19JQUvm2FiLC495bRbRsB70zfXtkLrzuk/Zw+skIO5UcXrOLifCL3euPOgk/Xgg
D1GNBZqiDsSMfPLVvlGxSvobW+WTj24H4yZ4mCbstCnf5EURtW2N2eRxM+c3G38fJBzobbP7Gkx+
xdmVxLVR2cvcluC2RQTPWahAASm9BwqQgs7N3SP4or38PXfCWGyohwvpnqrq9d1zqqVlK3E2JZrb
4EdpbQ+ccZL6xv3e4JuKvbs7Ad/tYyP6QJzOQJtAQKK/9rhE82zTWpyd5Pr1zvCi9J0pBtopSFzy
4Mt9Ve/FCw6h4cd4R+MLc068Z0dFtKNvahFiSGSbtuAKZxnCqwnycdbBRRAA+UbohhOJQunEL/FS
B//qDh2XYUVpNt38wJcIi721iE0wDNN8ObEpmPSyyNfzkULi1CwrDpOG3tLraB77vj42YWEGCTY6
iskHqOmJvL4KTD4gmiRppaWayc5kCm1LqD0A47ORRuDN/dvE/n4V6HaNysx8QX57MhZcb40u3Fp0
hpA4DV/8o+qS3rJpkoF+GwDxk6E5tSS6s6BNLPUt4sKHHokic4/RK7iU+WsLaDy8y64ARguzWVUL
3RAri7V3Yy6gqLgAO84EuuCuL6yq5syhQK2paFLyB2AKBaasncHemaIIM95T0PEyyWYE1K93pyAR
cZdoC199G90DrDHnwNWDVhrNyO93Oe1RVL3aVuPdaWVffeE1I2z+KZMJ/n/CuVWuYniX3WkBPGip
dZoHzQzLAJxiPtl9kWaVDjxikrqOnbP066FICE/NHLDYj7Z67zThY84ddtaBAClKBcFjq3KBMd7G
VOvf2DOpf+XdLGtLuPKCM7foRG2RGhHww7SqRP2fjiqrhqUI+TcgZbEabi+WTtvgILrhamxjdK//
h77njV/Rj1tI4nIQubSWzOoKeY4/Hw+5lW9M7X7Lxh/ELFpKGdTuXDGyhw75NWdZK/2q9JHABJUy
T69LhD5Btp+XxQzEyQTbgGEiRLZWUnzrNX7e/DgwI6bKFNXvVFz46fnAWu9FQeRpM/6r5/FIhOPn
0JxG39aYzSgRA8/fbQHzlOT8rLmb1pzLWxcHyse1sQidZChKUG5dPISd495vHrD4ZiZXYySl/tzG
w23tFHPS3+/sMuLQx4uQWdiXlp9xg35vfc/g6+pM6dYdhdDV3sPBz9HpTdwATsk9Dm5imLDDIrLV
Ufe3p6wXtxT9qEOQQo+BaclU3Wc961bbGcD5KUyUafbFX1JFO5xj0TetzuA1HkJDcsKLOl2cpzWe
N7GUjWk8YsOI2ZWPuSKGt1tzsRXDy5QfAVZ0Rlj6oaPDkms6uH0FDFmpNC+wSBQGC8p7iu/rRT8b
idQfYu/+z1/bkM+2d8YJwMxWP2P40orR9tvqZsWBZSetV/dzfs73tlVGLDs6G8J/M6uanze8vGRr
lcPVTL9HRiz5mf3dnZKtl5U4Xihcyp/QHNBUdq0K5f7dQg/reWqUTkQoPKVi/ESRJFpISuT8k+lQ
7o2vnFl/4GByzKKwvP6LbjHO0PdgeXHtr4fpvEKpRTju/gFeyzK4sLNFqbJz9uCrwajUoWkX09y4
Y8KQJlQ7xh7xrMz8sXUm0PRFbGse11Ev5zqu8u5QE6XD/RD3XJAfRacEPO2HvLcqImFjLKhC+8Sf
U6ZwvZkWeG1xCCzmhRgrAHB8AjNYVvQpmR4swIbilUAqH/bZVZTXXeHyWEwX/D1lu2yY8YZa/9MP
mzkZKqkdy5QZGnl1R6zmI4U5F6AVt67FVK2nbKGt1J7zN+ctVT604m5rmcWDSvIsqAvFZE89kSEY
wqIO0bItwzvAY64Tk9ddG18e3QWnzXIyDix/Q6tKCteCPd5fsyqfXKbltavipqneTCvkYOb1sGPn
xy6ENnFfRzeZTCM6pxhLMonqPgIpmnLA4+PxUWz8zPHwtl+SqbLuZLjfdPUWGQrbezEbryYH2bCg
sSzGong/XI7upZD3e+ZGnCEGfhUoNCzS8Fh3cUHtmeuERSh4tAczZiloX+/tF7Z478UXzp5bDbNy
C23lRqrLXqvIm9/eykTCaVLstnohdaaKqq6E1XseIZmUtZi+2t+GEVTExtDmWEkR8bAOM08LViYk
qF1+WxVb1m9z+esx1+YGrng9RLMxLZ/+1O1JFUOjFZnK71M1u/PyYKeKCboePSkq8A1jk1Kut5BD
NWl1PJH/Jow0Xk+rUJUSRFYXk/0I4UzsGM2Oxl8CZ8qbfu4mGEaJxgWM5OtFYdTzzlbb8B6xMph0
bbIa86zRVIebYUbX+zlR9h2Oss4zutFRBMkHThz36mu5gOfGpjb4JOKxbqYKgwItU9UTFUOS0KIi
lM0SQHE2O6ZMfOtK1phIf+PBPVD7L3VCY1UxYuN3fFx5CSJlNm1kJMF0ot8ugaPQtXzcJd5n5G6a
UntRwdpmEwuLd8dWi7oVAxp2Hil8ixC7OTa1fkPa5yP0bJ/d1NeGLSm2SzZVZ3ilErepEdyxx1g4
Tz7jrDmwjogAZShLYc+OvkoV4orXB38hL5+PB977zBmqJDwiVD7ptGcAluVP2GqcgasxCH8JfLDy
5aBqWxU1cvj2Lh+kLNsfmEqffLV1LvOciRoW90+hZgCziB9y0InDmJ3np4YizihoEIVmlWPAqL+r
ZqyUClVRCcU4XNS7t/HQ1yHPkWkljeVPRXFcEjqNnQKaGwOoAhQ5lxKzrbEYxzjA9ApkWb0zWLDG
gX+wrrThx/AVp6hw5cSpMRxO21JHcrbzFceHHJqu9gmhbHyWvHZ9ew5VNEqyamj+8xs9ibjYD8dO
61bSTTr3nueGCyJ8pGttn467qPaR7bD6npxu5rrgaw/mEn6phpdN1DVfbKA22M8L8/917yEvf6Ai
KUDh2q79TsS6mKDBsQyV10pOKJyGzHB1cyJxGYkQodislHtiGHE9ZdV6KU0OlfFQVLjD8COVtG7z
/BQCOsulRjBJ5dRoxV0/94YbXe3f7ezlcfNa9zwmc/yV0SXSyTJI0fBTzoAW+hKEKo5zvuE2+DB+
ElAGVH7llvhhIfg+LZOHq6Iy8KpXdojw2OmKdNjau6UUm0kQW4ptuC6mlSo1Kb24HlS3Zw6Zdy+U
KCNRo/fvw1HAFeoOXcY3elY6evZJaBPi+iBcuGg/76SgJj+QzuWp2/7Szv2pIQ2UWSJGCUIqmodr
AkOSPqsQNZHEPQswg4dS/KN11WiTxBvXMRTDzROUkVOiJlFY47WVYW1pnSP9bMDHuAmDsxqSf4hF
IIwq2LoV/DFItGWriEupACEr82h3/h94WacUlzKYTSUUZmww37RE1jLFGfPJgDjDKgDjHiSogSqS
vRHg9uLXuXmP1k1c0VRT/04yDhLx1PhAxfpzd762iSqFhb5ex8eD2dKPSrnmx3AdOqJKser/aAID
hqMZB01hVySb51SwpzXvgn0kGg0MUpyj/+xXt/wvC1YXMDZwf0Sgh4k5vIByvIYdYedJQYnNy3mY
GcX3gEdkfeuM7B+KUG/2N6ja4e6GfWqXGYtOhXSwayWjYbR7lquvBT0ZRntGJ300DxeIRJh/REqb
Ovd5/38syL4FWE4QNArW/sRpkofEvECFuO/swt7fhsxsWTP/4/p/zvvfTpzV6ZFmyxP/FY5vlj0h
0xsT1nLVvV/xmWeWg9MUBz0j3/tNl2SZ+AJD3v1q/dxuqSkEzDpIDREhV+X4wSyLoeqM8BITDTNn
YdsItJAF6d7aOYn6ZMGXn/OsSuKgKyNGLrcPhOyMXMu6Vkf7zvqkmAc3VH4/CdOWMjI+2aarERCa
BuMhCQywgkgiLp2J92tqw4jiCeteEvf/e+OVr2hb9g/SVgu7UBJAC8sbUzZQU0yuqNSCY9EKMCI8
DK2JPRVBkmBUp3RjU1n5mT0jHofM2m30wvNzWGKo5nF/sKiaRr5NsE3174lU1QEbGWwXhU5I3+lw
zKZ2LuQDTN78b7QuS21Nhl3KPJo9mN5MOuMvVFkN/ous4N6XRTWtr34x/kj4br7vGBsyPNiJ+N1S
8SHFW117GgXxE5+Z5S/PVCjVOTslwz1W1y3JrjBIz4x/fDha20O+ybGHw0PIXkcBn+pVE/CjqH7F
/ST2cQY3tReb8cYy6KI7MsAFEv1D0VOZ6tDPc9dXsu+RXk729W5NCBa0/XR0Ox7oSNu6ZkXwVgae
1m2iteIljSM5afvLBUUwWVMmyntgUBqZCGjne/h0woNJOVbRayZCMfaIsgA8YtkmpkYBZss1p+Lo
zbmpJ3g98T4EFWyv5/GkRveE/FPrKdyVkGbEmUKdi3yD8ZYO2HgpnEtwO0YNh0dtes/wzA+XdZe2
ruYY/zVlMsyIxs3HKK3rLiNixR7PC7Wr3kYyYmnyZ1oBG/A2B4+lT3mSNnxfdxDR9aNJsImJhNem
WwmLtpa0rHOYcebntEqhJBjTz22VqWT1T+9cc0AVvbImbdBnty1jnRiZdWzWGsb+++f0X85sdQC/
xS5QEJgGeSx4wrAOfltvX2fGWXj74/C1YzhuwwUICQ1OmXImC11Kir+HzmgaqmuqvBDNTOzRjud7
6lPcaJYZxx2CnMzdz0+DdnELUDDLOiCtv4YEa1DE+EPItxP1oeVYfOM+DzeLIb6n1xXxb6I/431z
kDyXfRBIfvRpgdXECNTHAOAhTeRnuk8aUY7RdwO4hk79+b9lp7mhwf5XfKcflNHgBh8aB1rJ9W4Y
PlRjGMXYPx+CYk2T13j34ULuDJ6gBZ4khsUghN1onGDgwNkD/tURRaXEihiF+d/pLn2OYBg2Mkwo
Jj27rMB1Dqm8dTvJWtkymS9bP32ONX2YSVbDWRJQUwY+G8094zLzzcAEAbcosauUj5tlBaluuYmU
6zW9+VMboA/sVwpnnXSDSs4JXxjY22J8V1oPdJCj+b3wg4ZztJbnkIpQLg4h6cS9jAHqeyo25zKi
pbRFvXcyyGhy+ayr6utzylkvD7rArcrS8JMEm+2G64q5ELxsEFtQCKy7bWts0xEseycLKl+zPZ/+
xd0+QQ2rvdhKejD1OSgJLBoSPiNMblbpe9oeR9EX60RDm6RKfJueHbFuLfECOjF9vbcKwkCiq7QF
9F2pZvHAwaOfnbRrRb8DpgnFpLfU2qIu5wphQjcUGOeoSjLElwGT4WJTm1EbeFXpk3yOO7iPMUjL
UplwTJ39RbpNXaQLPZdLCCJCzSCdivq4jZ/F3tgY9IzbeP8ho1pANoQ0ktKuEzu9TPzNTOM9ub6X
1DUM06tvFgccb+vOfJtkHN4XGAv+obmkc0u+hS4AqW7fLpVaF+4WkdIMTMW+coSta61ZnkqzVw7J
5aAplMMHEzEZH+uUQ1wFWOq2pht75njq8Q0F8vOA/jfZLu3dHSrQFgG5aIEBUfOvzSys+KnypLsG
MuN/TmEIJM6T4cQfdoMDXAABpi7YoZ5qxvS6WvyBIk3kRg5U5OXujRfIT8ACW/eqZumPjJw3hxG1
ktYZzv+bGg+NGSxl4TrQ2gN+AecK2eahLCICgxpxepnmBaEGzEzHhg7XMKqxrRcuLHG3Jh5a4yC4
RQBBFH7NYg3F27wLSvPoKegHbpKdxRs09jYqgIZYwifUoGB+cH81YXNTat1og+HXZRdChIKTAII/
HbvS9iLvWe0lIcjteXq/O12wJIystBvnIAwLuKrX0hFTL/od7v51x4/so4VeYg4lqMLCw5WQ+sZk
16aL12xjZE3YEtdVLJeap7Ayo1O2lLuS31LgOkgedBc7mvj1iV45u3RnXkw/7108Srwij6QQqokK
VIDdGZjklgAn6eM5vqMZo1XU4anG4Na9mU4mHUZV7BYlrZ7bzdtX6Oo+sv2NNKgpWOkm3YiGBqbS
9M4OLBuHNwy9ngCWdrk8gPHsqD5RhNLDELYBOz3n21JBXFHpVGeYkbXEwQAvLWnUPgRZYy5Jvr/7
Dr5T1lEc9Txxgxb5R8cHQ6+vijPYaRYBzKYiQ7fjlM3utzFw/XySH8sMGUNpBer2Gq9eUrUwYX/Z
UHZ0VqYqu+hutVchUrLnK5Rw4xAfJKOuVUh5uBAq8ELtu14estfBX5uvR5S5/4ZQdFOkQm+58f21
lFYzMwI40nNPb9fgxvlbKZZzPXUueg1jJAyT5VznZkxtf/ZOlGOxBlclO9CYyQEGDn2IOqx3n5Sg
jOs6j2/LVkPwCDbA618BHoQ8MvcAhWuQGGBXwHiwUkgTZfUkhovOFNfIDFajfyu0iXz810j4ik4g
jtW8d3jHGNo6j3XXJXvdxXxBU17f4DGvKS9PKYH1iRAhz5/eUMkqtJrzSIRFLm3wwaADCOQeKkfa
5AvgVlXHEPXCRbOoz6w5TtLMH/e+q6+moop0pyMhpSqN/P1G2bqyUOeX/zVQHyvgZ1FFeJ8wn0oT
bsPjK1AQ7BNXahB9aH6Qel0G3K/0LeQcVV2GqJYezYaIfVI5Ra6Z5BSZQiJINPZnJCunUO8CmmLt
sPGpwtKiKzGD6bjjsMqQ82BGwCD8XDSw7nGOyq4A330877n1hYJpeQwjyE7m+BHChpctjiJkNGw7
ly8EWsMkR45kNIQB3v/b0ODXY8iZ2hx08fYzdbch7J2tAxjVmkxQvRvZU0eJFh3vkv7TRkgCHWdG
Jtwp5OfGGpWY+sFtMRTeugLt3/OllN6tKpu43gVFl56H5Z+DcKIvmrzsamx/7ky4ZjNQUEmlAOtn
3FEd1KU4uOVT8unzisMMCZH9hmHEsvY8ZfPOxc5cL/d8gp4obufBWN89T2x2Px1pVV2nAeQFZ0bM
dV5n/gLF2b6FfJTlmv4IQmjPoWxERMDUgC6pf8T5EsWAYAJOMcoFN50cM69mTUcd7mGrWkQFlRIE
IsbTK6kf+WKfXxAFEa4CZ//iC1o0lG7CKjouj72tTnL1206g7r7F+VylwbfMFsZAAnu2DhXW+Uxi
8ZBjD2Ct2HSQDeQD9reFCAVXCbYnn1/xbT1a7CX3c/u9ksbnu9TGd+fxYGKbaFEm0e6+qMIhTOJI
BiVtK9HLxugdWjEQoh07rbcqtaD9OEAI05gL68UJ3RgVH31cg8Rq8ZhxybUovwyQlBSWaV+80vSq
p+yM/AhN/jwwaiQ1jvnSi3MEO3Ix5Q2cyWfAkwxBpS8prtONY87OPz3U4w9RLu3RsSaF4kIVauT3
J08+R6DdXHerfGpeXQw7dOjDr6LgCHKg46IqyGyHs59dYSqyAAD+Wr/TCGfTp7QM4IE2Q57U9Z1j
X5P9w6swJeBcJ6FD6XbdYiSW911AlrLGQ3Ajjn7B6dhT8lYEwBJu1fSE+zM+Iff1h1USAwaVrPpl
aKjuBTFmErVSorDrI6+d+ZfrIcLAHykUdEaXmyujy8LNCd5lfteq335eQG5U/GSp8CyyWHoU0Y1i
bXlURqQcBbITRfptJcKO0XDZfHBTg9E06czKvYjFNTXs2ocMUmf+w6e2rHBIneOIMduN9eMidRqr
GPDOa9mNnLVjBLkInhlhTy2sACsSEk8mvJpLx3diKnD56dQf3jTCnjoYKskWk1wtV3GAVr+6LnRa
YW36ptk8O7FsCk+fPK9ApMm3ybw0t1izR3OdOL24z+54W9puh8TZiVcku+mt0exFlQfHn/cIz3ZD
j8iGO22G7xsxvQPf6gzushZNwClbnoBSzSOuwqr3SQmjZiDNTKFWVewzTfdicOKCfAs4WXamS9vZ
mGI1SqtAmDjoSgyFzKFOhpRy9Vb6tvyuU/JFVBojRTOfirTvfm85FCX2SWcgqapbipzlzaCiF8pI
2NJsf3mm49PsvSsfUGKEr5ho5i5wbE+jmSleLDpASOSy2/3oLI9bmQEuQHmakOt/MfFe2c3otbR+
sy9p8cYS4spTVddHLvIeJvToaN0xLtkvYavxUZe9vmliy0JnQRtm29KJ9X3s4KdmAd3G7mp/8Osq
NPYv/sIRqg+vo7yE9xaV1A9tTv5dwnB8VeEud+cAbdiSmVxYnY9MXi4NeyC967G0LBo/8d7rNNO/
+U/4EH0UxqnW37MEXefurmV4/CBwhndybokY0OcaKrVOb30Lxfy6qrtAvaevzsNmSdXJvTHGnlSB
MFPQ6Fa+Ys+qgbqmShKJ/CD+Fn7bkHGHEhKDwUnVT64aOEG7Z4n+5DiaWSwHARQZluV+jnIpwzbK
8R3WYW78vkW3yb5IHV1g6y7MomSb/0HyQWorg88+/BcNqgurN0x+6svc6qQbbFYyuZjpmhWewEt2
LS4uZc93CPwPJMdVyhq9wAqnKrGn+NuP03JbY3CSZuJWEFOsy/AivWkpA6bHiw6nsawxPtFmhM8r
yszGatXQBa61EmsFLozk0hiT8YSWcX5uMMeZD147SHuKFlOXmB9q2Jfx3RBzTY6M+h75E4p06b3Z
2nrNhyFwgXcH3Cv7SuvLMyg8SbBvFxH81UlLiM2/Moq9B13XQoSFcg6zQN3mV7+Bi6qC5Lj0+UKd
1WiUUIFWPKE0wWhf8nbzIOUrw7KJih2t95ZP7bmpStPsKbyopwLS2lMJZUyc8AzwKAPxivy1mCBq
3HQc03FBvPoNI+oRQIwYcyIO5PuAR0dUERpDAlKuMIO2ArNoWp/8xdAP+iHWRZHNFxePjokQjMjj
24T7zqafuMoZwiGx1QiUj8j83WP/7t1Mb4WNh2aUUppu+0ialFD0b2r2ffeTnAl0Ksfm9XXlKN2/
PS+5+vGb6XgAzcACYq+lWDaI8qlie0e0tu91lu7PU+jreuAUzjkk45rHYi2Oai4PVeLgHLjb9acK
iVkO5UOfLodPcKlI5rtwC/zP7hOR+ynMNuLoENX8I6He/aWBLn4KNpdL11M4dUOeKbMQgd/C3yOa
rO/kqhVZ695BG2GMzmQJOAsOJry+QD8BGNVMn3snrnzapDYG+cjEaTwVO4iUBfGX3RU2o1iWuY4G
KqpIV/CHsUuHlMxUNUCYVFMmoCXiD731NFzu8QHZC620QOtZ3mBf8aIZQ3DsLYKknmCmjxgW8yQf
wforJDkhlUreDHc2QDmCZ+8anPtjwch4CyHzEQ4qvSEgWJu5tIh2MLQYTwCXUO0MPzMUOw711Flh
hi7CVtwv2/ae0uGvag6XBqUhZFqXxAQNag3WbUwc6e0EykVTymli1N/6eZ6gvnZuCL+yz81fvpuv
jbOs53Gc8uy53yYhfGbqedzsn3S/edq1c2oNf7U4PQkWlEOYA6/wvqzM2PdDBZ8/CcllInPc1LN+
8jEh4ELnWnIzs5LCs6YQsTy6d1LZ5aK0mkQb2tMdyQw6srqY3t+dKt/9nwWC7cfTLKkDgdne5Q0Y
UXH3Q9qOQ3BZO7bosoSSOFKxqQ5jbZwAqbIBxHRVNcWY3SFRwmY0Wl4q8tD6A98iVjzGrEA1mBYC
kzDVMMYAwYHztRPa3nDlylskK7f+lqUs08N5TjrPlZgEim2i2p31z4YCAn+3W0BV3dNGyAGeIAQQ
frmtFHG7N8KA86V06bhNXjiVBCNtRV/vRUNDm/vvl4GhkRfeUFEVYjSbPbS3/yq2az8g1AhCPLG7
pMxlCHOefxMAnXhb1qD0pP+c6tALjfikQGDt3tXYatCtk7BO9FVTVzxORD4MywNiopiXvfM81T8g
ruAU+W7HOdq8AsoWWKT3sd0ul0HvZSL0rHr6jPciy+V+v2v7f7cGmKUB5l/kJLOsFXkj4kfoGx5D
xzij9mgbFQd+y7kypMc+QbSuRTl9beKwaxqFB5kAO6rLFJ1BMQcEGO368+7699ugb4cDTLYrJX6L
P8ENdd8ice4qOLtAutfxE8eibXZ5dYJ4pZNabLfV6uIcOyFitz4Nvgoquf1LvG71QgiKoM+CBDDP
I0MP2TXcbmVQqqzhElMM006xKryGtgl47lxcNa8YgMscEXjzu+l6UH/HuYTqbjNd4exzvj8erYMv
3mMcMMvYm3gPEUm+OAjXNppYekFTtXCW4rtVfoe/fi9qnLLD5WSrSWwVGe6enBa6/yAFLCEmgR3U
AVkbX69as2R3d2/4eLjFF0U067jupSyR+s8r0FWQ83Oem2GNof1HsrVFjlTyGZF45/QXS+/xkYx4
OoKoL7vkDsJzHfYTjxaVir7w4mRqQCBUt6yXkAWxS1Yh+l57CCvxygVLh30T+JD0Iz+Cm4xzVnV6
NETNHhf9nVVu0yCnN30OQQ3mxxSWYh0BEj+gHt200TMOqgKaigAy20WTrV7B+KP5cbcuSpKP65am
Lc/s9SuA9bQ1ky7JbCq2wuc/3opexNdjVhFG7aaofpzX93To2kB/KT4rnroN+1YDe9bWCH/8OHgi
nRKqUUhN2HvpGvwNhRd6wFEoei4a2hFpkRRVioHRI7Sx2KMB/13sq8eE+T10H48TZqVX8v7hkDnV
xGo8lKnKRHf00/HmNarV4NdoDRUQ5mvrfKZvd3YbvmcFiR1IWArE5bLqdU2lyP8bEcOFNfyTGE+f
/tLxfBiXDxeuKptAqJ8ntpMYQylBeciuzI6zfwnZMBjKy6jEJ7Igkbsam8Bh0tWc6qDXu6MqYUix
wT+hbvn8ovx1EvizlkIahx+AQkA7uUhN1xkJ8d1libGCwGsVbethcbUQoPqv+qdazWspW09EAZYZ
C0I6UZ99kBGMCTO8AqjbTM8IKJYLJ+liIElqsrK18HOrhQH6SNba0XwEAGzHbe5IAn0zPQubEawY
WWe2rJJwBKeRzBCyzqJq1pRNeP9NpaBjDTLWZc5cVKj+f2uaWGZ4YbMDOi2itYbD1SrtdwqWTbhV
EXWp5/l4S3rpmxfNnccX2XR9G4IMTuzo4MihVgeWk4S48A+ETveQ72WA64Jb4lbRSPn7aeBuJi1h
MvJbrt2e6bXfzmojoCiYtjB9bFINilny91q5+aE7HuSxwMyaihP5emWfK7+tJAN2IL2idmlr2c2H
BV6bnyc8BaH1NIZjr43rdoh5igzbawi/gZ/m1gnMxgSgb0SIdl+vFH5QJUZ53QFmpOqN/u4t/WN4
Y0U6iUo0m6fZ0k3e4JVWT83h5FCTI9JMAIeavDpVUEeb5e1q4/tC+9aklflT1Zk7EN11nCeaR16L
oHJ5LHwAYx69bweDabeRisQYAdvrpOgukd9p+tTStCuDI4XzEQcHI4WC+pt3iYYC0mREkk4pVaGl
lEYejzuPhP+Et7h5fKos0m181g/Spo0PPawCHosiLVm/Z3tR35NJY9phhlMM8u4vu1CMc7elTf65
Zd+3z/r/bWAm6gj2WPBwC9w9RbSrTiVejOEqvL9rgyaeCC50JvnoofljeTIK2oj2HUOc5ASBRaJi
FWAqnlb2uhyrU+OF1QY16OYoEX1pInoU7818OK2si0uItrEdNH2yaGyLGmvk9cAu93Q+PpQvIEMs
Jm2aLdWtSiJppGmP4z3Se7R5Oy4AsZ5+ceMS2r5Qg/ZML+iFOV32Kud1NIxxV6GhOwtU0MFW9/xy
xvp5DYxiDFLlxg4C4l4xBLawu55C1wn8jcS6bycQq9fBm0nRzCD0QhwwOCWDo7Ql1B7obwnMPSD5
r2BfBux2TPye2GnbrjZ18Od6qd+ap0fMNOpKmhMZozBiIbflT50RkwmY6NUsftyeKHDMV2R+K9gD
aZBRoc5i7OWpbkUGtcJPbfnA9tW8OXNf++PDQzVJKKFIaGT9icKcIlCfLKKfOWp3t/YGbJ+aDcb9
d2HPLiBDfkglvQWIgNb2Lzt2Eszz74Z7B6NCcLj1MQvbjWrEPmg6OyjKQ3Cx8ozC4qv+Umj1RfPq
Xn1DjY+9qnffQYrbsWZFNvR2WiPlAqHzTRZHw874Fh+scrNsbEL+z/M6ZLOQ+edd8ZKuZI9MH+BI
XdPtNE7oy42hK7OiT+DJCm28DYATGcZ7kTSFBo0u0ofTa64GhpRlMbIllp7E6Pz+BlyS4htpREpq
ipgVvllD8rGi7d+smyCP256UQcVFnUGoqjuyWeYJ0hKSGBjRAeO+JapLfqhWrnqnql/fFPyiyIXX
6T+r7szUUrcxtiGPwBBe7wkwgT68zSK69dxq1g/2JjLbz30YzbwhoiM7nXykghZoDpb0IaTd3Owp
/K+AeWNZkSZ5IFagMt5tFea/ELXlwyA5nT0Fw+ZzXqOuFHkPzLo8Mh33v6mWMoEw3hCwsFc3LR3X
fS1BhtOtm42emT2a0Qdc/cLzwowAqhxmj/esTRiKUUuZ4lRg2I9NZ6NPRikCQAZksXlh1+flJrEm
k+p7mM4kwSsz5vcUSF8iQhaW7rs2YYJhdhNJmlU5+0J7wrOTQEUTFGuBSm8Br5A3sCrFE+t1Pmjb
FupgvxaQ0OCiYMk4GwWYsYc4aGwojxkkj+qpd5LD4yqN33gyO44thp0JRIFSADlUBVIeKFCQexU5
HWoQSkQPdp4TIMIpCH6xYxNXYGc+OeCTXw27BPFu5ObluLt7Pa0LIm8+PzSpEtAmuT5kt3KSpPpF
vMU9iWXMR+oPQ+UtBVqz0weFFFAr4w7RsUNYJcw8UrAkpkHZWaqMT9Axgqtr459l3pj+VKjHxsgu
C08rNPidFgFmceyYzXWeUbXUvmzORPs69Fnq1LVmscAeKgvZv1f3rLJ7UnJxARAu9z50n07gcV+3
UYh5sY4mu7ZBdylVu46NAnysOMN63X1EA+lgXpgBPF8k8OBSaWabv0WWB2x0B+cZUvDFtsWP0yE4
42h+O75cImMDln690mRxZZjLXXknlC4iFGqkDO2a3ygHN6vlHRjJX/FWz5pDFKmyICVglF75dJMK
byWAZ0TxigW6+MMxnzx67FpxZV0MukmU2BXZWZLBi5Cqjn6mMfHneyBULDOv0ks8x+xRvGnjiwbd
WDfC2AltDvxGec6OcwPhJ6o70ylgYuDXP0UPsPvJXPOMz1k2QbSrgSCfbW/3wyQkPSKzaZDnNoaP
8fmqjlok2o7TI2EedaUbEragaDhlp0qGHwQMIburSab2VN1ReH7P4QEfRWynm7SYkBgbq+7zROEN
TXksVJNwNDd1Z1wdJdFXvZeDfpRG5QVjub9+Qx0gXtr+eTTlxcre2Ah0KcvRaB/I+XlQtia9xMAC
swDDPcexc0lk04tF3lgjGPVVjZTayrx3wGva8XXYEgC0KpWyqjJ6iXOgCgNDIU+dE0womF6+H7Ni
oC+fEbJLF523K7/Hp7tZkVCutnnnRTPjY4MizA1qeE1KqgnD4e3Osi+/wwLAk0WJxNUhcCd/OhZZ
v87F1UXwtqUBQJBfMSifOZgB1f4UKdLudbK2F+xg6Tth4UIVEXZxwFnEruBTm/A+5DRHzbf9yRHz
XH4sWbDi5xeK60OU6SlwH+5Jazkd7Qmf1BrhzLn1WHHV/3dTy6pVhMAMJyRMufXUqU18hENG/Igy
JNfMftwBB+l7xsdMR0hb/33j2eMQxhVyKJ7pRWDcF9/Gsuy/uEw0+tkRFu8fj2084m3irXZMXhBx
NGFIYRx2voBavS0RKO8mON6QKBXuIbBFA730EHhXlxt4f5I2RbH3gdaEUqZVJ5YAvP0gpbGNfLap
vXPNTS+S9QV7R0Ed0kXeX3eML69Zy5cZm5Wg641726VwnegZxCNSVi9C0Bagu/aeBsMqMMuxk0TM
ADOI+xj5qSoOXYes8PX73kJFomHAv8xZChkzEHDdNLiOhRGKZqonKtVXBb8d9PgoIcbc+48fUsL6
P9ELG9gQYVxwwD7jb+igrnWwrb9xEA36NXtfPibSULYX05ZWdC5uaP/0IG7SODunqE/CFqjoILPz
SDV5/QRWpdtJi4YHYOaIV6lEhB3XF5Dg1FDmxrgnCJvpteM3WneH5yJWKS/aDQIEsG/f6eQAlBjZ
rqqEqcWTs7P+Vk8eejvM42EiRnYxHic6Ii8gV3dU/sS+3eF3x298eM0t0ny1ibeI9W5WwZilF+HR
Vk5/yTWZ3SrR79iTc6Ukcs7t6n2ZN8m6dPGoA1qy9nJOv/96hasJNXcuVUic7xDnoEDekVDmn88F
uqmARcq5ypjrth/ZPsDj7dq3KApKok+Js6jZmP5yK/NqITM4dF6HTajyKrOV335NCfi8VKQOV//j
QQVQhF6AruJ+VenH6y2b+eQwSUEORgEMVD8KSYdxrESM6IsKTatDa/j4Gwbn0g3e6ES7AAQ3Uccf
glsPV1f7xwaeWiLIxfeYzWATHZJSqrGkaTGqrX0USp6eFosNEL1ADNofRoQ3cACqyRRxxNyV3YCU
7PXdyjRCpNLdCu86OwUGLbLl/ZKvsAZ7rC1t+MJIuUBkmkZ1QU8CHClKvPUV8xubanED1pv2VIlQ
tpQ8bYfDuYxp/iVgUpaY02TfiQd+4El8XbZAFNczoVid3vOu03FK5piovkd7pofULz6wXJNy8kRP
JuGYiwxrUSFNGRKh5vE8Hv/OGvWFWcbmo/X+cU+53+aomWM5Kdgd9+fov4HW12ZDM8sJvdZiOMzo
Hkqvt3Xx9JqDoz4SvJ6SkO0QF8/5GMRaj/h804sERr06wU6Xuogl1hB/7a4/aMwjL1ORhlSQl2Cs
wHZuQDwwxF6AO+kIPC21nHzQmIkfutVvPDBt0FySLzAjDdp4VGNekUCHtH6glXZ/eJd1wHWuvTWT
rU28w2FWupBObd5NRGHmeR1acpNnebx/O+Ba7YZwEQ2oWoodM9wxWhXMJNRPQaYbGhx8bQjlqh4g
8p1usGefz6B/1hg5Uq4i6Kxf9OyGVmsbZyKbvkcj4tKF9GjsWLm92zxS83XKKE2zPCls5yB8r4pF
ff5BL49Amq+QUgmkppGgM2Ja4uOoc3nOnCd+JssTVT/VJbOABGnsT1si5wnaMavLNqgTbT35BbIe
EAlrl9M/A3OcS2opsfeqyVqj8d/Vo66ko7lcnQV27t6m214MbXPJ2Eigl850ghG3uILF9/fX84AN
5S9eIN93cXdWW+0ScRHKkiPC3+koWt0FNUe3Qgjk1Aapb+1F3I82xFXReKBtCDMTdcUp1COq1Wju
fDhI6yph1GCFhPiJerpUPUlhq4VlPqkWm8N6KGtg8+PWeZbQ74X9x0zx5U8FkeI40nE5d89cIj3p
l9MTY5P5rA6wjtibem55AveqNIHAYzKItLwZt2Bi0KwXH+smVywhQ8JcwgzeOudj2iBSUF0zn8/Z
uhpT0hdDPaKcseGgmNxa1vwmrih1qWw4icbxlp9XxWhavrsWOVSwAt8AD7YZ0ry5zWsTLpjK36uo
6a683ybp0hiD1asvvZhDIGXU64GddWV7bvqY32kwKvLgd0P34Ls2aYVq43t28DV5sA/1D83QNp0y
umtSAYj6ALhB2MxIZ2sXCEMk65VHroEUKQCavSNlYSU1MQeZgMHGkh5VqecNW8no9W2MIwS6IVs8
awYcV802RiRuXOQrzZkwZFjiUhu3Ful/vNfbQOJqxPAyQvRxLF5BTHAVn/jW4jtzWv/M+2zNXEdn
Ccbz1HT9Da8OM5xtIjTvB/QT4RwQtildqajqSuMxQf0G+ZSXbqkx4JByri2+r0nqvMjqnG4OHWWl
lZG43ZVbCt0ig7ozowxIq54B5YFy5BRZLqyEwFqWqEi/NERLWtib76A7CrpI1c1aI3bUgi0chvkv
fV8XLmzMCnTg1pvf9w8Uf6NrK/gCyo4q1R3qf925bvT9mxdZ9NcL6VSsoyhUbYnGT/XPwd4ZwGvD
FScV+1SXmkKYDNvcJX2stRXPGmbTrBIXmJycCgBwS4ULXh/9YJXa7CANo5cbN1hqrI6zR39kWSS4
P1bymTRrvusynftVX6XM9/3gWMBr3c30zrNpOGQQ7yRkm2e0ZXRm73xbegBB7uSG46C3ilFVfXVf
Vyl1TTxflocbfLO2gKlgl9P9Z2Pu5pbbT3wwgahvIwyUyxHtMpVmdXPqGWG978kbJvqnxgYvv0MI
jEacA1qEJpxoPwWRcjDdttVDioC4A3UuXAZ8Ewejrz/pyrCCxG3b4uzeSrlCDcxHWpw6oCmCg87l
bZANhiOfZs4BpIQ1H5GfuNS1+RghjN82fC3BqIhWSsOqL5dSAYKwt/Osrk4pPMS0+S/bo6qbeXHQ
TTXNo+Ho/HA5YaEkvtlV/gXAAbtoGy0AH+OWqn0snu3tgdE0IshdzIVZ+nnR35VF9RgCxVdovYdA
vkXCceoeA/R8qJFvR/3rcM8PAWEHFnPi5sO27neQcNGtMvNSqEqlD40Iysh0FecEZ38bgK7/lrQx
0wm2JOPG0Y6ZCKTEerd4qqxlMf+X/+535/aSWtujC451UJKo0SOCBb8m4AOxE9o+Uu5qg+1Kku1k
prrVOpA0kW1yo+2PvO69ZogA3soJGShERaoPU0IrWdDWzoBGEKhj1e9BP5oDgKQCwZpHHkbKCI0Q
7oJTBLW5nh//4CWuELnnW5VcPT3zc+niIcgkrzez0QT2Uk7bulx2sukNuEkMkSrcjOgo8DxvYKnR
bK5Dkce5O0JnhRQrfrSKeafmF8L5yXsUAKRF12sthq7RKfTop8IpemK6CWidMiJgpGjVYr67qXAl
UwhFbLd9rwbCvvhYKQjlfpaHEHlM04JF+3iYEPsVIQS6zi7mlellkBrCgkACfvWKw41xhB6s2Sh5
lkgMRxUfO0/FeQf4UpYXif4ftRXUfJLqOKbjfZJQAaRQHCnNbCy9M7KTuZGU33FG9LXW2OfcYXfL
kOfPQVSq0moksfMbP0BxHIxFYTGhmaSulrN/O+vuNhr4RJPs8wa/8NBT4sxau5406u8SCKqESonL
FSCeo7zk2ra22X7mtSH5AIHJ+GmonoVem9sIroWjfGqav/xxxtvUJJ8WCfrksqSnQrGuNIE3Kk17
R5HE2KJ2Vx8aqrTw4+gYay5f+wBfNNCWBVsnxEJTQl3RtrXuTIcAeZRurD8MwT4n76qNtOJ1rUza
uTcvBVkkREQyez5SBk6g/ohV4OMITGiiKASq5v/P7n3eAp2ogVAsUmu0aTASRRXB5/JipXXJPPQw
DiXA/asH3lQIRQADEjKXp39CW/aaQt+8nQIp2lJBizhbn5NZXeXgEBNb6yTUcBbncne+j+++mZB3
P956iredinaJTsoKgHwWdAnhEByFLlPuigZIhbPNbhE/GU7i8ePnF+K9Wn5Wh+sfrq7EgUChOzmF
MHY0LdUSdpvRVYCRqXrRoG0OrEhbJkVV1m4YVqWdcqkLDQuVP+sJoJtIf7ZBshgkFe4K4FhZvzmL
lcFQk+fW++6wdK3ypTMap5sxm+4k2ctswJB+32IFH2TaGCiDRS4JBvG94N5//9fSMBe0HljzU0p1
vefcH2WdxCIZjsID0FphwJnqpOt/+3iAm2F/u0S0+LEIR1l+xiSLMjXhOLtl2vK12wsOm6cLeKMd
piKn8sJgBxmgfdqdUdWD9nb1GEePeOjyWRR4Lzi8jbzHMJ0SIQuOm+/wUZ8p5FClpZi3oBxLQeUD
MJe58poN+37tj126faeGGuV2kO6v89THoC/0f7BbIp7BJfoHxfTLbCcKLI5Lh991SFoyTeMUAw2G
NzA++xsyFJiLvXyXr+x6a6vlnk4hoi3e4We9OakGxUDdbNWJPN6GzXnpBigzFsbeQHrthGZk2xMR
jjrLwhi08cEGi1IH7p3B7r3u4rvOfNZ//OruU862C204yzoIbxXWaBfgDfXF5oj1Yvi50jPTai2k
m8vwXAXQgukTsfqShiTngMKKnrxTQK94yXxSAC0Fp34E3HQgqcqdAA/2MQzTkqN9BMMbtYWOXnm8
Hx71sobc5pzIC0wJPJAo+ej7tfjoyJBLMiOzgWvf+xgladNz1bm3cVOZ50LKamtHDkg4N/GPHFkL
fSSQ5kp2mVR44NWlL2HxyELQMHgo2xnjv68dxyfOMLpRkz10VYbFZXskB0eLxzk7Ibi/LYa0DxSd
57ib0VjJG4C5UhwesyVSfbJ7z5oBHy5KcJhFkJbxOqqFKyZrTNAXD/D47cr63gdvtwUd+V7vBseU
wX2hhBOQ0D0UoEZYT7uUwZL27KZTWtoO+rGHc+Lh0aS1hA12ICvWdu3lhQS0fOKljXfeCBHqd6ov
qEglaVc+1UwMGWU+z/PfOvIxLMKRw5d57l7AFU5qis38I5Guc0KxlYMNkMtupkuh9nv10iLLfSD6
UJGSG61CVA9q634xagHgAculv7qp885gERzLgn/82N0aYhinCRTZUk257IVaY9Sl7qgYGwdVUnTD
hOpiae/Iip5Rv69WkPpDT1AapECrCsTFSLuySLt2L+zT3xQhPqIevxfDn0Tvj3JVPaOLA+Gj7VGf
RQSljeMo2SWrM4N5D7ZifuZn98FS1+vRhfUi5mh5L6aLZryLJL8z0I252YGqs0UMMlz8M/Qumavn
SiSNbqX745cvyS0zu+Yimi0Zh/1osk9nCE4PMHQyWgaMew0HKvBLT3+nXXYUvaHEqcp4oBmOrwIh
i0MQcOvku1FTrKY4GiwIfgNNp5J8MrJwB2pm+JFIiDy2jdpiIg+bz7nI821XGAzbG6L1qeSjord6
9Z1Mc2rXW3xsvgV1UfrDKgnDtkqcPNOXNTwgGEgGm8bEkhNhaI2XEl/d7/ROiS047vDgVO5RA5hf
lsfUp4BGofzpNwlt9n3ibKvKMqiR4NnENLmo6NCddYkrYLqb37FKXnbsf0/YYddQamxDQ9X71Sbs
LZzKoZN0IOL9/CEXdWoIlJnJ5GUnVePweEeIZrLG3970JEJg1OQMdHdxJrdxs57zxPE7P+A2GXNj
8+fQdNwFWYZkhf37KnBNx195zlGZU6ltr5fWnGLnOyF7sQRY3HDE7b03jP23Xnu6kKXV4s0Dieer
/M6LnFiE8knteVLdzElOFl7hxvvf0oKZpJibTjhXa++vKsPkkgcdv1DGFx0z8I9oUEdtFMWEUJlF
eo4NEfbYPjQZSRU6WiE8pvONPuCZ3iLCUkljUit82OPwOiyoJcbjHoMX+DlmnARXF+hQb4SCpNRV
ZnFsYxgxN0LQNZEygkuj/ELIVyvZeCSWAMv29YKEegw+rO+Hc/BqJ0AhCGpCD7nhNGLNCr8KDa9D
2lI756x5GU81Ocul6aBpAlJp2Fzupl20acBzzx+/Vl56genQci9ldE5YyDK6G3ttQzGNTx/b4gqu
d+0sL7JPonh0cXhC1/V4dSVEgyaqr41IK2jG0/3jSFu1XXamXBaF7nXq2xycp4JRhF/rUDjAio1H
Ll7OnFfeXpiCBNPF+FUWYq/xEn5yWW5WI9PB+ORo1P4qC8w7RTkQtCmRGkDFn7nHvjJFjGIDNvsK
rmP3O+w1diXkbhPfUH8Nr1ITa/BMPNeQj4JozmXpmopt7zNZj+6AETo0Z559nmuG33C2t4GAqEJ6
GN3sFraY3Hzmp51jsVkaUTzQAD5Vrt3AuQOOlsTNkNVtCIc0ZTrJ3Dm+UbkbwBi8jIKcqSERKYxy
Qq70RSjzC1r93tKqRKFmlZrHJ+fu/AmrFYzzgL//Ny9xT5Mdt0eCUi3u0zQA86yhd15ykV7VK0rj
tRrN3xGEa17j6N2MUvYjXyBfqalaUestVzN+Qio5hzPvzP4juw2IeQIuYeSdvoCT0N6mk2CXe9hJ
1nGx3lwn/qL9rUhlK5vMKm6nKKFgqtgW6ztGwlZK/FbEK7zLRgcxXdaoiN4V7MdrCxIFeih++z6T
Zy8bPHDygNDULShRfN39ulObIUP7HhMH02kS8RJbFNzSdWwAt7MsHNFrcbQJ7ym0tiS6PjFGAuVN
SjjRljpFNNk6u55PgxVJz9QdX0aqXxUkM0hX0rTZ3pLd2bJ31e/RS51pZeVZ428yt1DxgBKNTH45
5XWUa0UrUxBq9NP/mvKsvG/4JRanAQCecgKAw8b5qWkKu9+wrlqJO0MLYhOeGPPCseIiBTu3eij+
StfYH4vtU6baI+iOHpQMgV/7kos/h5V+UX1fjLk8+8bLABTfxBuhhSSuk1nR7gcboXb82wkvfXRL
ue0ylDoR3OR4xASTQm+WWg/U6k4vr/GGKj98JzqenPjareleRPWixB9gMVNwvVCl+bPnsuHTDVLq
FoFZoOLxxMGmyZ003cil11Ir83BSamD0V7mZFFUOFsb5L8YYJH8sgErgJyeQg5zqNce1xUJgm62Z
LWOpkwvneou0wjhSnzxS7M7usbcUco9fL2kKPKAvp2dj+CKB4IHGPudltIQF+cjJ6lmxetpIxY5O
qL8c2F/Nym4fPejzpBH/lQM3aRT0iv1XL7R50eq6ZtKEz/nvuaVRic5+8qV+Z5ZjPSSjA/2LOx8X
7JxuuMF5RJNvSg6nzWhYtzRQ3oJLb4Sm0MG4B9s53R+hq+kydUti4gWoLvdQT3hSPW5ZSpAVuBEj
lKKcyCT35NGO3ywc0ap+Mf81wCH4GNp8jFbj87O+WoJK2qexF3eazzop9oqJVz6JDUYr0WLazglK
/QI3lEmabbrPpUuppNZM8bTR2uxnVmm9b60pOJd7yV4W58XHCd9kRjy4zw4Vnai3K5r3CpSIC8EV
XvDs25PLmTIWcSlFz2oUvi4KRK/odAoj6egnb5TIVD0irbZ/DKhJQGjMMfP7yGLkf96d1UoQhG4y
FIE/1Shpf1b/4xbf0ZYALlYqxPlzRNDjDU3JP2zPhCK24LFDLfco0oozhJpeK/o0fEB3tKIEbSz+
C3dABr94SdDNYk4u9zIuY5sxGZ/1jQ2FJkOjaVv5eP83g5RScQFspvfQDOdnPSfN9AHp4vc6X/s8
zbXdc00NWMD6DMzlyLsDAOwa33n7dljRIDdyAvIdRTup8QlD5akR2hW6SL8zehWWGrFJUzr2Qaau
OY4lkvvDbHYvWqAPS4xbmXPFbvIYQdXrSr9hNZNmraIvPz8SHPvOZXwxjd9BYmjgoYNOHDpma3g+
PxMd7yBUV4ZQv8uXj3QGH9aUw4maZInUkA3D+usCQJAcRMpxYbarnYmg4FJNk5mBAuhNQg9MNark
tTC0wgbFLD0AKmzYqzKvCm+lPlMT43vJ7ty3OUjXmHll+4n+1QeMnvkNLhKP6hr8cz1pUeC2T0Zm
qa9+BroY3vhV0sbm+Z38URAnAiGoLdu1UhR73GQbnQS4ZIdlxTo0/JJ3yg5fn2WSoapWMsGjRaqc
PF7lM62lyl5XTibIWujdY4JktXda+XC1ulen9dLDJhK8kbMBh5lGTIXFdBZY5DuEpGLsIrN54F7/
ShGWWRAZg0U95IPhpX9W0nj4MdMWwhG/uD/73yGxRi54GavpuIW1h2r0BZAqonRrxjmqrbj6IZHS
mfHYaJQ1H2HoNeH7Xtr9zIsbFy2fKgRZmdJBBp0rbdv5TJlvXRyuzRUDcNG7sI/rzSoiGVuef0xq
SyOh7aw2WNe6KiueEl5WIQaoo5B9TjopFliILczsWqeidDzyXLbSeJYLXeJuDtWgcFOw3oeia0A/
dKDB7CU5Jn8QW0cBuifI3Oa7lnhectwBNWm8elNVwEQlXSIsvE7TMkltbXTJIkigFuIXlQSx0Odr
Rl/hff5DMekVyLQtl82H+BVtbN9FP3+SEzjIGBtRq/4tkrQPF/MAez1vK3zRtICgYETuOkGjJkOW
MZBwVOa9GY6xPfrFVXU+Sc7hgWOTHcglvw8kumrogOUI1T8X1bHVact7WQWjdKxb5RJTDR4XHnk7
YqqXbhOaYSiRgw/n6+aM6a7bC91g3Awb4TAEHKnB+HffXSDS1t4arFdt3v7r5lwoeW3BimPagO5U
MPt7i588kGzUH48Z4dcMjSShXL+qgHPjPPViyPPfgH+TiKkc6YHcZ7aE41znshQwRUjoZDa8ZRsv
sLJXEAG3deFhvGju5w94muZqcieogZkZ3Oqv8MC17DIa6nI4za+zsrmF+mSnAOY6Xd59lX/EBBxa
L4fZsDnRLB5cY/hfgDalKjwvdroPYM6Z9KM2Y67LRwZXrXA9Ei1d/2dH7kCq+C0hlNhhb/KOqz/r
Yd8jWLLMgG3kcp/1nSPdUKSfGa+Avx/VGPV6EMeGHuywB24qkwqOFv7RxdYtmM7jhhL5ArMCWQDE
4S9cw/8OgZShPXd5XlxlNSXvwgHAr7UWW28wh9HFPlKEiZQG1rxA/SSI/kPBfxLYYNnhcwqEhlqY
EL9u5t2w0r149fbWc/S6+dCyUT5B0ivlrb5w/v9sj4AxO0zzYWAxdL5PD4McZPSYO3AfFS1BN4tq
1k2KLKSZRsOomMWOCunnjK35FtGoc0iBx2wavMY7CIiK2kCQxvoGFnxtT5LCu7T62RDEwS7O8WSd
KWgvg4GibCDIRMJnq0BtgjaYi8ffm/D/6Jb/zj8upHDG9UyeDTn5TLt6B5L1KaqbeM1+4ayQHwhM
i5j4x5KLOPKqh7icfBawso9lC5Mx5L2VM/tOeA6eQxpy7m5lAQDgQPyjuCZnPBGMxq8MtjzFmWoD
kuHehB7dquJkPotwo07uc+DSWKW8tnvuo5QUcByS/x4oMx2u1rj2JCgRykRRbT3Mt6lSpPZPccOk
8N3EnRDnhQxrkhYQx8uTyRCpUHVCx8WTLeqOsV/eHfdkBZZ4iVU/abfNQVFJV5KMgH7ofHkmzuSV
KNZvRsdvFC8xcUEk38tsHCfvQgIa8FAh4K5m1TCAg8EdATSSrRlHnIKa/hq7rWVFwr2TePzcy18i
oLmXCm5tMc7acPoP/JfA7wntx4HzIwwSilyLYRIX/mXucra59D1zJVs4mwgh4ZNGN9Rc1CMAW0RS
bmNtnpoHL3BiaIqUd0huhdq+/UlhOlM+NCQGlhJ0JDFogtZYMQlpwN/AHbfAw4ejlU9f5ggTYMZJ
qmgspST8tUqLNlZCYfmZO6sXyhOyZWDKgQPksmEBw2uCajLt/D6YzqGU2LZPQjN2GKT/8a2yEp0q
+oNj2z/gr/1TMJUBSVI2zAX6jTK4IJepdS4n58fHHmA9n9N5hw7BKK51YVNxB5VLQf9wUnVpTDlL
whEJq1tsFfec0w/r9HqrREuAD0kygYank4HwV68ibn8BQ40wkunMltK5cJBg1JFggfFQwOSF2dtG
ityVYq4P6xslRWBtMGCwqp0EfZiicAvzXV4Vs03m6gEN9e83c2fd9VoDX3mzxWm6CxBQeur/UMCl
pIG6L/P4Rs7W/I7ch6YuwZLtqgWXp8+Ug966k7lUMR+83bFnXujdx/CVuDzjG7iIUmKbFARsvOZR
So5Rxf40YP9kkAkepgzLQltGruI2LWG8Tc/C7XChWCMPvFFHPZdsrtdjSE9Hdz+BQ6rGhkWUBL+o
O1cg3cXHdbJHVYKZoz1n+EwTQDfsiZbl4rcS507ennQ7dY+H9SHde3E2aKUpReUo5KJMhKKjdD9S
98pAjS5h/jmTaA1LjtS4Lt14yIi6yAXeu/VokHSV82qJIwBi8jJj9+n+FzhiajCGbF551t2wz+Lw
nP/xp7W7kqEljoy16hEcRCbRUaGaiFhCOYQbHOg+5r17wsBouLrGmyfNHqEQgzVIR0p6C/u+9pXV
W/eeM/b46+0S91X41GjI8VcesCUv+0QJhNFsIXd7KNWm4Jr7YvqxXxac8ucmIXc3NJ4oYiwP9o0I
13EtG1YCsAQkIxhJYu1KgQX585vilZkB0gyp6saFqo0bXh3WPgttJiXd4Ykl4MPIfdOWXISsAW5j
xGw+HdbWTF89/DdC63eEQj8IJS+x1KQKrcpS7d520mjEbBtsYM5QogP7jV27f7Us4vQOOCEsoWfw
Ta7ig0RUCF8tBxqUdzHKTKob04O6VpaHW7x6NPzCWWdAeOKheZy6MTE+PWodTHfNu74SvEkIBhg8
wu0/hRJnSn83Ii7/MhcvRhH1mCx7Kl+IvyNEB1o3PfXSatKe+/hYbZYAdCXX+sp4NozmhxrfJEdh
NqXb7dIrt4gS67SZELtHvuqBlQqYmzdZ9lbLGdqQbESldg7XwhZqPdKJPsM42FOwbDTHWXsM7ufm
59n5UybsKmwOcE0R4zlW7ehctABhPgWyY7ck+xpDvzbT5TosGKac8Y7m+gGmU1Rz3nsStj05e6io
XOyln/bBlQ4ACNqs3AxAMAZJXQbXOSdZ7xsgjnUEA1tH253tb5YbzsBqQwYkH8hSQpZXCeiBvPNl
Q63d4To0UqEgyUWbl+7fIg0XKmFzxvLCoDJ5gKVrxrbpFNF+11pr6wQ6UGNkzNdpRH1WsqNVv/Yk
2lsZBnk03Y+mXk1jtj2NK+EPGENFK8f/lhcxLZMtvGbV35SETdWHWNPNaGToAFybXqOC7BZxJR92
AmVskCfZlp2SIBvkyR1tsJ2gVffnkPfNqK84RJzbNFcqi8YoWOnFmP2OFdE6zyEoumAnbzyFhFcn
mVJfsQESjJHkZMndU0/AhDcUFJeZ/iK9CTRc4VnKbsxJc1tfACsxqEqy6j7KZ/9YfeZKDrI06ZnM
HEA9Z5fjeMbnwN648GtDN/tOticmG+NuRXwiADJl3kPk1o/9R3vBNr6LiHDVxSsoT5uDLdAZt9BZ
aEGyAPqbf85mZJO/Jd2XYDubHqEzhNtmzK1pb7pFdYBj1QpKXhqsxdSynoKqloshaubzl5+ZCvmY
Z//Lpd59C+oJbklvXsGrMnZp+aVRIvGrCnxaPAMd3umYlRv7jgcFhBvFW9PrD0BLXuznl+yyZ4pl
YC7BzBbOPoISPoKuq55I9rPKrYSQl+ylEn+Rm/ucYAGGWKYiAFOQPJUldi3rNkFGeP/W9bbK8X/X
rixx2sj+BCiTgfeaNza5gS941E1FEj2dv7HK3ePU/JjTd/U0qDNDLfh1VzesLaRrRS8BE4iUp5tb
m2zwhdSBOzVkTRB6Ocuv85IieMOXwFx4zl+QalKYoyWV7Wyos01I0DIAXdtth7uhO4+XDi5ckygO
i5CHTgDX3KhYaIBYvT/Wd9v9cLjBTu3nl+zN5+lbPUZzpRuMv7smwoMp++wHPDzuwPYt3jBjmzX1
+zu4FVoQewg4SNgcIoTnM/fzE4Zm/3fRNZ5AyZR0e023uj86XAS1uDLUeMsrBgNtpvMReY8PMaVR
tsVx3JKN3S6fgSj725kn6p7vZquot4VK22PhQp2ldhUUPMrqI/lqWzyTscesS9wqUI8ruG99/mp5
OBvXnE5K4E3aWWi/GEIjEB3nN/FjgcaYzCauscf1jQcncpvtSAoPdxu8SQBb8O8XFQGiqU273ttn
UxppyPQSuDE9J017pCOrpd9EbTNyRhssSJG8jvt751cpF27grECunlUu2KlCTuE+5/vTa6FBZakC
sn4tP+nATHOqBDDCPuGzxzBJel+F+Zs4nyjofZ4hVvaO3ZzDO7vzBYOwSpbfwoNiKdeeAi8FVynX
VcBf29EKrF8n7Y7GiD483ikfZ7kHtMxf0VJG+OgysVQlkPy8zGpdz6u18aHVVIfeZS9sluDJsCc1
/dcYBEeFlWs1udcjXTs1eifZwXQ9DVfHuCmYGnzlM+Ke1UOF+OgZEFymzMWcYeuGTQVQcoyu9SjT
T0SBy5V7Kh59bqxwo124ccH34y3GGJptUm4Kxdt9treHhTmEjWNC1JQxLkvijo8UJkCH4hjq5mDT
TvxdXD7HUGFoPYP/iW2db13n5rZw9z/y4/YqnVgppXQGTv1wPFMnkG5JUMmXwIH+ub8xYfnsK+kh
6opgO+gElRV/RkFwaGzYyXvuNK1NxbqtTYAN30jSDSbFUTbH6yOyy2He9PJ4BiqJjppAjYCnmZcO
MlNwtvLaQWVbJAiwvc453ktqDOL4E7YNYo3vxS0BVrLmNxom5opbyH4fQEhACGjUvpaXd2AQ6uA0
btKwl4tspDMHexYA25RHCCmXtI/86BrNRJueliZQRegnNdedcB1JBIa1Oa0YqTzAayDZWzJ49ADu
J71SgpSTNI/oXHq7bOCnXbODtKUExa7OkmVVh3d1m0Apt/J7gVlsUUOAmogLyYlbFI1TriCrRHtL
ib9b5D6ZN/HtVlyMNQCSer02oBQYi+vFnIvsbN5JSNFLkPxf+aKLwxFpdLDvaTgeLf25pCL0CIMr
j5ZoqFz+ADIVWxFPHnvrWbt2JKAsPDl+bX0AVq//cNyBN96WoUlC/D2xZ6beJ5J/EmQyL7k/C3Bh
2VgPvJr0+wkijY8LMuAc0RDjhwdYoJgWZ9ABJE9AJV2a4EiyzVg5I3vKq+h4HrzvVwWI0I6ZbXIq
4PHN7bR6Gk0/NgpoReNv1dNZm4eHl/YRTBJ9aymNwj9o0FilgPJbxv7lygzG7OB31B/KquLiLOtK
QoqM/Lwxm6shtQDGfdb959vqCsCqsgg9xhemIbR6y9Ywb9rtRmTiixA0W0VuLaY+GzK09s9ZudiR
YB58uGWFh4CxnHWCJ2eRYgRYuqCSMHuG1Agle4QNSvnmkIUOneLtonYK+UIA7HfB1QBmdX8jyk+a
OXUbPDWlmuk5UbgS9UVEymqh3FJG/ibBZ+1T9AIlo8rKGN8G3BTFMB6E07t2w3kKlRZKrFUV0WOv
HohCZKPk29qyNb37TIpQ+SFdj3tzWUU7NgaXm3iluLRxBukH/YOH/KjGtc6vjcPSmD6J6d+DJ9z5
MJqOTt1kFjd1lidwGzCCl4PvBh+ao0btuY4RqNmdSpLH25RAjzCL7x8nH6mxbDLq5SmzE5s+Kye2
JupACpwvkbmtretWbJyeNk/e0Qru5tDl3ZbT+N8WAyukGFmPCQFRLoueVvG+9QDgOu7d/edIEhYq
oNKe/TX+g6l3VF3uf/269rhMY4almVv2qmvd5F6BlmvcXP0B78FqHA1Rd0KlCPINc6jDowLhDaKf
zX05Qh1b4cTe7+f+U0nvgm6YC1ijd5G0st2HUaAmLvBJKXGttBb0WEOxB64+t6ehJKLKvPueOGJ7
iz8hqqKQIemFnDZ7aTs0TWMuN2WmwNoLWtfiIK6l2tTD8dtgv2tmPxt85AwJifOrAk/efmgQ/OTG
2qWTcXJzD/yg5WBLfzkV0gJm/jJjhfVa7vmP8MKpG0069iduYmiSSV3kk79nzpqxz1jfHkVT/N54
I04oCPzmWNF2DnDvY4f9+Ps9/Sg1rP+rUU8nVSO0wu8K49k83YLxU+GKszGoQqYhl6rMPUOKQtUi
MERDqE0F8I373yy0oRX+Ks6gBPN4Bp79h/1MNCeQs70Q5NtPNrZ0OuCzKeMA5pW7or7GwIbeHAzT
mB+YmdRcsHNqZsGTESqY3vRT/utJA4dLqCloR5HVed4qBdaUpiFAfbh+2Ozi9M03sJ9LBWZPiX/E
ZaQsWjLYQrrz2s7rLf+d8bvvOGfK+7PVHhw0Lof0fcyhaTFVFh/6xSTUsUG+akWNoOsHPAMpv3UN
n+5G0+JemTrfcSe8qXgks8WcS3IWJHQDehNqS8r/vlCNNiR7SjhwcrFDlhgD/+T1brykX6IoiBGO
inT7rAZmZj6IGQ/kVa8wXEzE8nnbqPoDmazDnO2CBxGeNNYA4YuatXfWFPq0fgdvFpc1HKd6c9Rj
OJplMZ5eXmIft/ZzMVMiUVLY0MW+0q7CstC33xf7SNYHvMpwW6oNYOqntYj/B9t2e3ZwV4Vj6ocl
pTiAISSYVcpcWF7EEHVMg6iYmzRGuXwtp9rtokDnnTBpFOS6McjJRV+kLLTYSDrCLY0IF9Y5Wvnh
6QLEQDyrwljZqaI7r+ihJxwzKXUG2QC9hB/Tpvb+7wbhQ54qMoCOTl2WHrboXoffFGuOHaGFUT+k
j7+8u+S1ZwRw6J9V4GTLAWTW0+xTAiEHWPiNNFwhQBci/aKHip1cEn03EwQUtWhR6+vc9vaPQi5T
+QfSwiU+ga9dxPwJpW9OwC6bkdwNZjaCUGvE1ww4sgDbJKF608qfwaAGepDE29Pf7ZzX0nkwwPLw
K3OuRPLvfwW2BAejS82DGLp3MtZOfMKMz8QoI50i7qY4XOPaOoRDMEtVLMwpoXRuDo7x3Qf8tWE9
L02Z8ba5JsqphGVCxV1CjznaW1GBVLhpiQkXhcBxxBZCRJsktITtWzducHH4cpCdNPk1oRKWkcmd
sH0arnkiTdiQm9Ml7IJDMo9lWAKp4ciZdXGooyc9AzBr0YuTgsxH7Zb3qfj+rQhBcZ4+fm7QAH15
O8wuTBtqiEFyRVhrLyj38rcuT1Crk0g8QN1O8jra7SW7zFRB1Wm+fjkQk6mm/vhoDk/nteFaUmeb
+TxycUouPuKlEtyaM7sKStbxAhpvkpblSb/64DX5sxR2rugG460kbDhHb5aQz4tOT+269Cg46A3c
kdt6b08LQ2bfBzgVcqpVbkbU8X78H7SUz88ruAev2MlCuvHE2A0Kv1LnH/1oHEkSn//peidKlIgK
yZZvMFhBkq2xI1gbevRloLUm/Cm+6ukhkrfxc1qcSAx5q+bZmVd4Zjcgc1C+Susim5qJU9XxHMZJ
4OpOsGY12uNKJha8qwpKZroRydfGiTFHQLy/IfkHrG8F8uJCjGMz8Wler7vfs/n5ja3UJqyPZCBO
ottf0NTUi35odwY7T9CZwcmHwegdnitivJxH5KgUd3ht2GUs4zODj3ItwoT/Y5EnVjvevMlgTMnr
UowPE2irhpNjv/MWPC74OG2L7oKfV2JwQb2kvqXTZUmY8rm8RHXOSCeB/fuLZ9Z8OMSs8OGpbkKA
20sbBzvAqJcwnTxd2mOmBIx7aQ5RZkmN5DUs7MFw1l/vOTzd4bdYn2vhJUe+HMGhIc2fpMwfyFxM
nG7SYGjHus27dMkwaa6e+XYym3wihNglsTfVN72R80gLrZE18J97IVnGylXhNjJ8yGK/N/YlGLsO
a9KrgT9CarJvHxBw88frMMQhm4qHJLjNF6jC4cEOrS75XdpscPw4GgHLHfHhH4sgEj3p88vvNIJX
pGbmVKSSRzhUZfiAZxaFB63Usdo9u/83HPjWvrDXdw/Bu1Af7M84qDVVGz2s4KhG72xHhSNxHMTf
enkLbCRhKS/Ku1ONVQKVV+jryccd3Vke+YaSIt+xlCAFrT5DZRjw2cEATJgia2wk0paqIZaEtrlj
cagwtCX74MG2cdjlzZ60Wqvg0q4VZks4UxBltzlMOFLP9VE4sUg3S1mht2lLY1z2j9QfI9SqqTad
CXPvtxUGRVq2cG9k58v/TK5TBaNj8wjPNkaWtbsgKOxcr545FC/0KR5+w+JIcAOD6F6C/9fVHHVc
qmV8xvu+yqZJEEmkVh1ClVjsEVfJ4JUq1HorhsoIKrXbKH1+kSDOMnIhCnn8A6bnV60R0occCeXn
GwcSbuNPC6R1HwZtBBfRUm4Z/47zWZEzLBy0tlOg+FiSWotk0bkL1wMINxCMULhjCfBwxtUsno+P
j51ATyDlau++WM19q40a4lTgkzhExVn899bAymunCP0xv/mQWmOMSYZs8xWPgbOel/v2lmoJEMbj
Qa8uYGFGuUdMdtAHzjUCUjgd/4g2U+DYr+pmKKsHjmkj8Sd2mU4k1nihJWNDCdhPH/Je6Mf80IRA
bGp5FglFt3kOm3Ly0yYCMj6w0MrqZ2kQQzH+Y+laGMya+4kukUoIEJ2F/7ygocELLxAh/yo1b3tG
Y3bhp9eNZ8X2QTBcExE+iZKzycvov/57M/2kJd0g0k0t6m614oqmej9fXyf7vhCAz4P9XnfXsHhR
IvZ4VwMK15F3/3nJpkAC8VqWq8NGKvExq98bcipo7HhW88Wz6GsWrp4c+YvGEo8kevIsbVQ+UHQG
eBGWMwybIgcXz8X+yyQJbzs6Wyy8IVXPBJdJot3XkQ/yL+I2wtfWCxQa4tBGYXWU65E+WM5NUF6Q
4eUVOHxKpWVrMbCTVjqu77bp2ys8xhXIaTvhCaDp49FJHJCoPKVbxU44MS0ga7/yvEkU5arGt6kv
ER3lemMfZ/Nd2DgLlhRr0Zeyi/qG4I/j/NCuU9oDWKn9MhovlstEPWDkES74ked1jRvqctneFYkt
00pdma12YOV6WTQKrCgjztk+Mq/IZE1a9ai8r84gnelV5X6W4D2YAfkmB5LTzXWDxHnBpIImd/Gh
SPwPTlr9E85KSd6RfSBSqzXrrdT3Cedr7jqXS5gTB9R/3AbF5gumMrCYijEWbJavRPQoOtuq7PAi
Ujk/Mqy7eyan2FJ1mBSokodQxvWaZInsdv5EDjC96sf21RdOWDTHBiKCGS/6RZLRllK2Af6dJSA3
vqNrrNYJ3nLKx98glJgPQHC3wHCAqGu25csSg2lAHq//4Vp/I21EkXN0zbfbQWsn3XIr8t8zeOjI
XD7KU2P+5wk2v1mdwwwa7RDx7kA55c/Gfp7z9n591N78uNeEYyOk5aBctzukA2bkaAFGYaIBnN1W
KQttZsJzF+easN8EPQ69brzz6nK6Iw6uek8afEBIuK+kacBSjxinQO0RulJVHKJnumicvsqK0eVr
/RMFa04v/yx/G1WObS975irI6vBtwsfd/MLx9tOekuq2qxmUncCdJPyq+1FYRIgBObJrxThJeVWb
YvXFpztU6JC8ecuLcUH3ejk2qM/FsR6wwLcRhQsqn3ETj57SzWNGmc0iRme3ym+LejOttrtMY1z6
4Njdd+ca789ACrSmESLzDB5cBg8qVvjHtqrWAmC97V5ItNCHgi65/GZ6eshdk6jEzA5cKqIVLJk5
Ij+snIl1Zna5+StoJoSA9NOhC0qa+LiZtBr6JWfsguiVUPM/wLuy9xBzMjp+pqekLJ3jRlCLy+4Q
4lO6nE0hM5I/Fpy+AxWex/W0a4NXnJx2wmvsYvYAWgKQf1deEQ4uO+rncrn67kNDXp9/Plq/D/T+
0G7KSzG6YA1BgBXXg9+ExYNJ7jHErAiAR11CqPhmX2p5rXELXOa33Jr3AHygUpYeJRHcgen97K+w
GvUVZ/eaoWQoBO9VOeB8RPugiidWI86xO7iUsGtRPZKy+W31Gwe9eYU/9VwRXwFAg4nfqQg6LpJB
jq70nBKxJny5E0Zmc74ZH7Ey21AwnwDOKP1Ug1H1Q8Sf7A5PXICbmfpGLtLWxWc+hqz4Ig4o6fnh
KulYhizbr4ybCQLcGiakTJ5XzCDv5H51iAwRf4qw2m0ve808j4fboK/47oZL0NgzDB93mg4CFhw6
4+ptKTgx8o2cFEyGmytniELbkEfYk5QU/HUEqhlBd4TOmfi7t4p+BPIoXFnVAFBW72crFsHZ1Wqv
uBiPPGBnzO24DNvvBEBDmLjwcnIy22dV6yqN8Zbukh1xIoQmEkAiHZT+pPrP3Xl8HSYAK7f809pJ
Jie/n81/V0hX9/xj3R96X6vEe4XP2DP62jik6EL3D69wJrIsDRq9P7GfETuUZEycDjsvM0/jFVGd
bOcIVuBi38L6si7YAROesPuMb6vADHuSbow3Tj720TYHMyXJorFbezhnCEf5rLbQa4jb2zbWjr9v
ihUywoVHspjHmPgeqfrWWTsuuzjtmCGZ+GElBpVqXARJ6LGv9vkl+2O/5eDPJ29+lUv1PLJGXVDO
/7YCXTt7erFBbKUyBrtUKbuwY5eFfAW5Eiqk5C46gcYGfy7v7AG6tplfUR+0TkP/HYzARq1ZnyBQ
kOh4VMP7udBi+VJUYYgCiP6lVN9YqZiZ4xkD1OStF6VRI7DKSF9yMnmdSK5L3YljLzXYFDEGB2ZE
nVG0CqtnaclGvW1gQaSaOgdUiy08/amPSijW8+3P7uy+mhAiV6SPIOyTTqnVr96de6tM42LQhhLJ
kPrLlRJltGoRIgBrsbl16UhIlZcbYrmY07cuQAgfFi6gCwcmhB98NqgaiRDE4M4LBYiCqGy04mDV
dQaBB4thmm8T/9IpQMRUB3xH/oeoNAE30zLcz3QeLoggVfI3LaOMWyt1EClEanAA0NyYhJnV1fO3
9Yv3LtAoDEQummJLw7AlTyENVvhiQExV9Lj7HDSB0Ym1nB5+6bUpN2uDmPYBhepU7tWJFx1128HK
ynX+KmeGqhJq5WpvMTVsViddAs8nNlcGC2RnWQX663X/pCwIrEVrxC93CrSLJBRcS3eZ6NwSlzCU
3hAp8tPbxGCp/p/RnbcVexsFTU+xjKZs86Bei0pbmNvkqZTlU2+cmvsm22/Zy5Z9iZ6PRSx3u9Ll
azZNto7TbVv+ApPFBXzXas3O9S+loWZ1q7dxEwsWikkmgbtWTLV88Q12idgWyRhV5427a03zGqyR
yOny6lCmkqBipKgEmujRvAL2mDNUNzShlI/q+u82hgy5azkOL5kUsqFFgqgv8QkhF6wnYfEIDY5i
EiLHwrHBI3JWnH0KvlsJ+cSqZ0VaA7QYzf2H6FxX+pmBliGQGSlX/lYBkk2zrvkWFRfH2/3KgF7O
Jovr8qjoCm5YdnD+No9VDDF+/Dt/+CafKy0LdNBEuaUIz5UUZCRhhEeaE1TnW6e9KoWuXeFyxOh7
blfTUtIxMhQ9jqG6AAtbZpuNjidVrGNPEhlcOOrbwT9bKFgcsXh4EA9i4JDSNMacHZYFeNMQXRRR
NjSn+wjQT68sycbMQvJ0/SrNRui98ZoDbGCvxkffu3tu4e+FzPp3qF9tTmvqOIr8HLrZng74L+1M
qC9EPORXe80aU5JgClF9ex/EhJZNHmtN+aFO6uGUcUfFi0PNN4WpFc400ar2wsf6D4Ngy19SlRyF
C3M8ZPciVvL5m+84uK+rYTMa8cVOU5AWYK2u/9hz6yEsp9WcSrSWeRltmo5IwfV7+PcZ87XehepO
5DXw97lmPl4sB/50ZUzlP8GcY09JjC97Zge5vvstpgUDJ62IKLru3ILXVV45e68uBhu0xX1SmUZG
xH5CeVU7MecO7eIog5KB4UvJy5DSYB86Ut3x18y5mdemuIErbO7qXveZLB9IDoqzPf8Bby2mFgjn
WOyDVvkWhf+8dEzkyXRurRUsVN8yrBJdzHDbkgiaznG2JCtE9jqml/Lz8yQrkgTzOvZwOZOw4RYZ
tQdnEsi0hLbCL+K24qPQkdq/H0DkLuMgx7CLg/oOtVj/oN09e1Ytk0ym9JdPDqCjZhYaurPODuf9
FdrcMa7YzFIhpvEiiQWjVMoHv4c5XDJ+fuU+tkDImuHUj92S0gd2//M9ZY6FZDFr7lTsI55vAWx4
oqZ40sslzUKYKnuA/VbzzPlLUvQdVIUjfqOKnmAL5CDQVxf9dpYgS5ZmVMc7mQ/JsnOdZ8Zo0jc3
uNbsrggif+SBYGHRD1S4aMV9Dwp8cmdKyxPWJm0VfH/ptBTx49K0vF9FAazMhkTox7KPjN6pIr12
GYILlJDf2Lon9PbbqmlO7Pb14YlxmQVYzwRj4NElHSbzIBNz7ag3zx0FDP0rsI06mG513dPm6hhj
On7E8tKIn8tTCPkm6H3F3Z+N42J+B800dLDGzWxzY9SdI2t4bMY8p57ijHQHRQEdUAGT45FIHRd6
twHpLUNGOgRjlqjNTJ0zhQzD1timZaIDlqH3oIIYouBnR2RWbJI84YyULtm8hmVbIega7QhBQcE1
juLjZxWjvUnpD+tH53mq7YOZxM9KOfCLMF3xw7CgFyQ10ZF953Mzu/nuNSX2G3uP4k1NUMAAojmB
0Ks8T1YAn3d7DvKYLf+mbyixF7fLZ9b+LOT2nwrZafHjczzQt0p26XKevlTM/0L0qGxM1QLvdPQs
gRpmnjVC2FwVChc0zUlriejZHUBRpEhsH5w6GQdItNjo4+6LFrf3RKpU3n/HClOf1MkbG2BTHbLn
8D1SOnGsw1n2OhOlQoUGM7jdvHyT6R5QMgxsdLCdkEDzEn8JvF4Q6ONnIFuLpm2SxDjLpZT0V/vy
cQoY2MMULVQTVpN1pPg6cTyYSicyf3/1PCiAq73G4em+XWyqmgYjH/AEPqN6cbOgC4CxXheI0fsx
Qi/O45eObX0BgWS+qjwTHSSrqcnSmLywDXa3Rf3hnn1eUKQvf0varl7hX+HUK90iRD654enOgW94
NCR6cY0E/3UZnPZdEEc0a6FLF2lvYNDFjNpc8LS2NE71nebI+XS2cplZyWNnNGntlkJeEFRuVmoD
yYkImCYQqgrxmHwGoiPCjrvs4Rj21XLyENKlyiNoj5/9sGUEV+BXvq4GCoU0yPgqUmUL4i1pc+DK
y08Fk+aZWkGVN7XXKMYIxzw3xTNvJYIBsQ+Ack9uRRBF9w4gL6tQc/m7qZ/D+WKADyOc22HUDF7H
ioHacf6GFBcuazkG4BvH+dVGjeSBVV+6HRWqQPbZdZBnKhLlJuKbeR6oBtiwdvWL4wymvfOK2JtV
5NMgnc4ZUKNagTLn53ONcVai0Za6xoCPmGSpAdzwY9LIU5dtOsyTjgmRrp/IQHpRybAjY8s19Hyh
b4z8yeg14tJzV47UYvpySS8NOOA8k+NYhLN1R0eSzOro/dZ2l31/i8oF2t7332Ryog6veiG5JtEc
ne/NYPfsF7wpBnT8szg4rTM796asx/kWZc/12wCWeBKUzPC7rci4ajZXoHHrtPO45G6y/tlM3N/O
zjS33h2FyvOjuivA66iN0wTjkTmy889XtnBYdR7ZDm6oA/VnJLQfFrs4kk35TlrGoqThHqpcp1P1
7AwO1PNMCkQKN/oaEyTCJIikyLOEPhjoYL7WPSlAj11ZcbK17JtvAK3T37bDyfeLT7FsyhPm93Z6
iHs2F8eB7RIe8gmWPeKb6fPQRNEwdtE25NC59l7FmDWSTckZ9lG3ASsCk8ne1ssu+FTIuoQapO8T
mEJ3zbOwW22PQ34Zl+y67//rDnGK+n3IpWaqRyV6sTCd1Xmmez5VOtMoczOPsQoUwipHSCha0LvJ
EmNiUWfVuGLCsZfDiB5P4G+Df0x7XiC6/jfV+oD5jc+3wWBCaCqsE9cjbXluagQUWa2x0Ccxtu4s
M/mVWo+eLqJe6k5Bq7oOcOcd82DaTVmr7zom7ytJIfN78TH9iRu3o5HFSwqVou3gihBn+/zJCrwx
zbN+lb/yN/ZeQ3ATBcVHVSnC3jnyAqGK9xeHswx4feOK+Ihp0YImiXmPvFvJ9Tbw5QMVgqkDVYSk
2RWFExAPUG1WwSEQ2GXdZQ862LhXWckOLh6J/EBOcDwE3yeQuabkZ+3SupqE5R/7A4ZyYJoPr2Ds
h3NPYUcq7pkX3pqQJmEtRNy53E9asv22x22ZYnbx98bmbtgENukjNRajFjKZWoqgr7N2+GB8dC/P
yZw0Uonf1Zc4hOCNKkV8WwWRzzTAbNwpcAah52Jh0dqpAIPPa/OOY/vF4V/9v732woxsrFY+IAQN
/c5hhbU8V1ieEb52n5io+qtqGwVx3X4A6U9uskpkjMP2qYy7TtrpqpynswT1lY60WQ1kME6+q6hi
yTcHgQKwumCcBMj1Vhl93gyGjC12587a166aegWCEuNGleSkmwxTXshUeiLMeA9pA4A7FDu1dLyx
lTeGovbBVn44I3zuDyLGtOhWE+VL0PeVxOX6HgiaUx63vxavLPMCys8e9FzzTSqh3+SIfyWiRRE+
YD7nlORLiBHa2DapDjclEXQ8NQwBe9SQxb0iKxyfdE9tVCRNDDsRkprvrdcVzNv0F/rbsvJlpPsa
RInQNaisJ1MLWdN2EpXk2CJygwBnoU2PBDoDv0ydhmCYCulnRjJMjH1NkSaq2jEndHkPZREASC/Z
fsxWRxYIhlcK3IFxIpAl0xTNikkok8kXUJfZuttdi0sxP96ZbZY9V3zTJ+NmXu1fS2NATv/CthPe
HcehbWY1tQ5xB5kBuijd+fKgskgZbT/8Q0tCcyoB4UpMd/V/NNF44cg8OpWVrhaXAV42zTIHOHX5
JIT+Pe6i0EKefRVtsHcKVT7hLibqWDNd3SWJ4fX+7BjVEbGyyr5x+e3kFvOY9N/bue2vzHEeIsl3
DoYMQ8O+a1pb6tgxL95O2HnkXm+wNv0qAC12cOBtAxHhIHh0mhIddMalTkS/QAgXECWZx6SBPOlX
GzsZ728Vl09+KdRV1/8zSqCMw/84/N27ywxFcuR78eFTSIgUMn/bOk+jRY8kUAq/+LHI0q2nzvkK
ua4fg2yn/5tU0rx2USgDkEaVOldiSkVo4MqGXPqf5g0qR3caiG21RO82nWIk5v1PcndwZS1h7BS+
AuDaKg+yuMyi3eSZDPZPtBfg8dJdZItZAKxqC9DqZi/DzkvYV2n61ct339qX6i4AsW+yrx8vT33a
WUT/Pu3NsXwVVZjwp0czq3W1A62v26i5OAkhrezottsdtfh/XDw0/N7ooULkC1yzr8CDdMXuqS+C
BovWGZCEr9QszXOKqOkd7PcN54LLpKu2rB0rP/Xjt/8VSNFmD8La365J0MuwE9egoQnYfoIOjF0O
fIJeAAiszafrTlRLDxeIrfsW5PxRrz5sOtpVMu+k++spDUwCPTy0yOe++s2yRvW4lT4C/dhcm11i
D2qOmMGISdUt2vVIYTEGI36KGTaCwfSLe1d+JfbURSAIOSxiZbHxBSKmKeW3n143kt6Hm0Vye4vK
IEHhQ/U9Y0C29arT9Kk6KgSFJBrcs54v1KJKFG26XUvySMTuY4RoMcjStlL416uQzMVhtAfgnfUO
x184+hh2MSEsWYFyeyuA7ta1Fgg3AhgZP1AoeCpLVUxHHs0qHuDz44iTg+c9TVw2ejX5FAjNHmDy
rQsSizDW4ys8+6a7jcEtYM+c8RuX3Lc6dbwlSPPepKMySG6xM4c3BqI/AutnJC6RTiaqpuDdHItx
EOlyLz/PEa+katn15IwAhdmGA1rwb+bBNSyvqfKEQhvjYnDkAIvCBqA3qUp7jIF7X5lftHRKuACD
nd6bxHDv0PRJQ1eXlH7KoaOSwgy7NsaOxK7Dwi3soEuVsItVbHGduRe66zboraswaPf1+z8NrR84
ppXULHSVisiypKiNl+j5GF82lvEa8mV34+ReJRNV8uIk6wsgut6Mw34Mpox0/5DW4qdVnwU6fFfd
H3d15VFSTLkD4qA3aSWzL1QJCUOWjqnJO9d/UgrdGbgozUlKW0QzHFouwo/sbzZRLtTexZoSbWSX
+4zOOvRHv+dJwn6sYhjy6WFrK+TdUwY35DULLjwWeZ3SCj1I2QTKN7Wupn1h7ntXxRHEuMsoIggw
t7DIR+BdJd9S1vo2eCiyz6GHkQk+qOKIgIRBJWQyRwY21SDmrl1v1s6OCXDxZPnYe9qCZDvKBsHa
J0/4Oe/XwA7iQFolct1QG3vtHiGX40iMjCizFZT2oqFEUGZEQUzJkY1bcPP+ChV1VBEh3llfTA2i
Ncg+Ywj/ZMicQm95WYmy8m/nvYWZIFtnn9dhnoYa5I7TUWk1Rw5ASZIelr72w7QATaJlAdKs9bXJ
/k9cr/AAu/azixu5pj+PYsl0x+mfxg+0bOQSDzLsoHVoHr4NP7u7WAQWrywzLgJrExsBLSd97Qfo
4jF0OMPI6Xxpu7UH4T622Pumsir0FFppt6ojy0phQ2eONSV/g0/6Cwi4InFLOkNWK22l2a91J03O
Earxa2fuXIZZNL5yQaBv+Q/eueP0SlDcPnjdcde4/JQaYjBRWJ3VgXGcuOcHhdajdSE8SPb2ZJLU
mThEH8gnQGJ57amlZUiyD0QHUYaK2CuK9g3NeolrVh+O+nMaKzcI629m4Cexyp9H0gF1uxDgOS1I
oLWxP2qs0IF6sI/KZzMTgQxHEYqq7QxRpwxTHmhZYCMTW9nG9ciQdb0j3429Tu++Wc2r9vpOYkZM
Enp/FlGwgBThp1EVyc0M6zZ0A8NhzCXa4dmLg/gk9g1PSnybynUzZJlm3Im72NWDZNm8JqmPT3jX
nr+8p7SFrDS75KqosFxl30nZJ7SqyJYBCsChifwTKXzAeG/x7XIW/pI0879JlZRURfhc5ZgY3W+m
bckEb6kK8qCOJsguCJ1DbYSGlfFO1E9SwT/vH/UYI56yP7Wb8eeIacajx6CM30kO4HzHGsp6G6DR
UrC7STBYs4LlUpZLPzXMW7OcLZ14jL6/jjhU29CoPH1iqjtrxMDeBteGrT6mBRpNT4eDSDBgT3Fy
wonkdRgEMKewUMpGHtnQQncTIKtJLX712nq7RlKmPq0LhlFtD/3Mgwc/ZkQaGv7UfgPtOijTNIvd
AkU3a9kz7oqGKi8SNOIGsFmWwe24bhZz4KFQ5VEvaolbAaSYPpt9m9zfNPKQVzuypqoUYt6IvN4m
VFc/Pmjms/o81YJE/l6lqvSaZGjA24tCzhx0RZsU46Fzp0UmX+OfBCG2I9PMbyiQFyZCN0ToQQaW
RLu+M0KtfFPbT+s8Jg2vBv7SE7VEMt/FK/bOzG1mP+x3BSoBASW3ka3k4PgT/Inq5t3uzq6Uqyca
XqKzek33PXrdYSWZ44EChOvPuh30Hf6FHyppDZYtGfel78u2A9phPumeCgdyonRDqsr08YKPc2Yr
6x2ufg68TSbv7B09emfibDGp4n5ekyGkfsOi2QfR0fWnaof6uHt2ZpP0bv5DZaF8nJEaB4OiI+Qe
BCx818fOde4HR4Ar07yBVOD0pRUamWiJribcOPKefX3C7M2sZ6QG4Uz9xjZolPJsWtCOyMLBZI8l
wudADqdUHOb8vTxe2arnAANP9B/3XlfZi7njjUfXcZrzcKB2pipDt2wzRk851gN2EXfkgu71vRa8
LE4TRn9/+KRP/J5nCpERnQHW+fn3RrrAaXQprl6aw9lD0XzX0VhxLyx1yMg9edgEf7EYraOrH7dl
Mg/dd1YZircs2HiSNwzOej4eZbvgmJth1WJxhK71veFZxYE+shsWfUsJM4S0JI22KbbXNfRFF1j9
CEn6bIhi2mhsptXsv/aiOEI7pi/BTJKyUG7kzx/BcE8Dmb2jefugj3625XGJB3Y8Bk/Fk7OFLXui
wQV5xL6nv/30mRTZ7EtLawJd7Gzfh0W8d7/E66CdBRBjv7s4dfeZJjuITLUEYJielwiGED+39I94
bXAIykTSs5Y4/id9nK2xOIptoFdGQQlgw8jx8d0HbhezDKUrYd3fn+cTyIq6hjO/zgNujB3qOFNM
FjjpIBt0gvLJqmpzFK6suRfxtbVBMsKUB4frwcU/jorWveciOrmt4P9AiXMpzHQCyuWG7WD4pzRC
DfTjHr3s1tD0xWhoadvYV4weEZqzWA7jNPqHCOX15jBfIsC0Ojr2ggBhwb8dXl9mX0BWIsIDI25q
P2b6t38xb1dd323/NkyTNH1lY9YXk0hpyShz0hJ6eZSuhLAUgMOgpnrP9HOPmBLrXb3OUUtIg/bB
yEgOSPWn02nmXci4PP7lcfGV3RDH4CmoW08/KoTGZjwKhs9nYFac1DeBAbvFMtKBB6WqxuawOh+c
WH3vXG2jqFZzeCl2gmfD90fZEILcw716xJdX9YcU76l2c9c4fIs++EGYBegMiz3Y1h2HOPOv5yC9
iti31G3FE0LldMtfO+I7T+zbaWC1Br4Bzm9IKDdAjweuGnneW8dg1JL0ZbZ3MBEd2uBY23GLz34Y
3SSXbelkzpEUa5zFrcXQIMW2r9E70zgJvpUwHQ4FAvc56ffJAlpQCLSbBSz33bm/RQfkdcbOMJBx
CkBe5DUk72+nHLCy3dMZWkBwl/Rk0SCDT9+RDoAY+H1qqMd3TuqNwQL/jnnr+i2c5tCZ/ZsOh4G4
xnrSwhCw8cO+bX0t+h6xA3crvMYznCHPNqJ82160tZCBTS9kZTqFBSOSNJP/llpI0WrACl1zmRss
3oEPTx7aVsUS6FyAzL7mL1DCFITstGfmk/7UdFtl4lJPfecYjEFVkB/XMfxp+i2AioT/MW60+sN8
gHfdHbJURLm1XOv8TfF+yUWCF5VhIcZhTEZW/YvU8yLgM69dJPd2zsrIGam7XyPI1UdCY9BKXLng
Eu9LlOYMMVHAncvPMs1haCDM5GRWMz3804VRBfJr4Kcjg1c08g+ywROjq8vLZbm25TfTCk6KNNqz
t+p6owgc0tK44d5qH9RSiZQQMlZWfvx/A/jIqxDBwnXYw0QFk7OaaaQpK/fCZQoRtkfXvpN3J+u5
P2AuRzu76UftCbDkKS5d/89HRaJiwm/nShxFhPe4z2WrRndwqG/kK98cWnG8JAlcuIh50T3hMFGl
YoYD8Wsy2Y7FyBBTFzP5qA5QYQ6Lo1KzUc58Vf/a4mPwWwv+gKIPt4s1AeJg8J+uhg8lH18hC7qt
c0kEMxjU0pbxdpDoGxY9gW+PO7JZn1Wx3qgqTLKyNJPf6e7MWg3Cff2cVALG9rvktwFcRyB3ZkSQ
S7L/uE2+JKdM+NR9abkO4acTPnBeC9EytlYiU82HnhO+HNrdBiOBN+UKeJdjhK+4CVwsUeBZvr1K
PIPGPpZHaDNJ7wubRNrEMsj4ohmUOmcIeYs4yx1iYZajau13vBlCjljg6gWHyGbF74AgAKuY6YMs
e5QPoKOieVmi2ugIX8Wh329zj+tpkSCt76wfdyCTtowDkgSHLOH0t0Zkk9MHfkdyK3ktlnnGP1FM
Y1/s0TVwpxRegePSfHZBxdZqM5U8MdcI49ktvIgJj+irtAwu9Fth9q3hpGqbUpc8qlBHcLZYdkkL
+7XGJ23HhvrznEU76ybg/YNec69QsHxZQ5MyWBmhsKuWngyk84vRKAmt0n8v2xBthMXhcGqV++zZ
9XsYS+etpYTLaFcEsTNm9Fq8OXi6P5fKe89AJeLHAvw5I8zCoAoLpVtJ3t8swcE/FdGzUXKc6+Au
KxTjb7nRi5rlhA+aE61Tzm+PUwvKM6gzDM9XArmuDjEaPy6cAAQQRlKfRm2SqozZTMg32HHXduNP
ELgssLodUFyruXaD3F8F07niPxhNZyd4UagbU/nMHhNDqovjkccQIwvOEL41eH4U3PsmH0adnaKz
XAR5Y4Hp+p2RmSahGneQ65bQbdvkGO3+R8tfa80dwNNVxseYTJkkw8RVDU2qNpm88W/BxoK6VX4s
HV6a+NL+4PV4cTtSC69W4nCqqtu/3WLjbKa50z9j3Ji03ca2B9id0Kn08kvtK4cddIDbuZvKz5/1
iFqEgrDT6iQjJehqslhwFoKpp6xXIFZ462jXTZJwQoDixpgLI0Bk8ohANB4VFT4dEsX86IyKgURD
7UCqJGxHA74FZXphwz5Tjd+cMLbC4Gl3ITO+gDx6ypsuwsLZpd2Gunw7dE8b4K160hPY1XxEvVe4
lWZ2GAIdySUdT7WKUsMvt2j5UxXiRUPtwgtLxmed/LfHTGYUC6mzekAsWONqgV+O2Gi3UGIKyvdp
DPEDsggFn9kxOsK4bbdZhC13/3UrZ0YtvCs+FS9oPHyX5MUT5EpqjzWEa6YHLiyhY0Arbkzr2CBa
fvZ/rxaz1a3AKOXTayHGzFftyj7DEQoA8DF1MGuR5SxfYLbQ+fQxdYAXRtLuhlr9PK6LUlPUfjQF
lu3hajKFEg8fmbGMmrr6L2Pdg6JzWFpahC+USfvsNBy2yzH1rIlDPZQZlCgZe0rYDnwwMbey/8I+
Wrs+Vejk4+W7PufpOmswhxSvqV+E3n49i702LpEf6UPG2ycCuaFZpxKaVUs1fBenpq9xlazYxPYA
BYebf3hdi48X30QdBNhXB2T5EvfeflYltdyQ0BWSxWw3GJNJgPKJhClOoej3T8K0cmaX7cGp+qQt
rOeEfPPOqRVCaJJg5MtHVR0+Try9qYzkiLqjuMf73OGuYXBMshLoWhuDif9MiZlQGwSVXDczgBnn
+IUL7WNmriKa89VVNtr/+N+E125Ys2ONhVtSA/Og6/FctjSnNcg7Abbqvp+zT8vEpAxLozLo1hxV
3E4y/sRrSEDB+MnHQUU6OL5jywOO6483H+RfEvmfFTDImpzce9fUXiS+KXqf1PaDCgh+AYvwKp5R
0WNiFd8mCiWmDVPmFeJ6GMqdNTSjtL1SiBs/TaRtBFMv8ze9VFInKpbyTwNEY8WI9Vx9RGQFfcNU
P8ll/2K/Pbvy7KJFuHHmfhZ9GmpzzQVQKm7l4pknjCkgR4BWXwXcXh2dRTLRzultoLNIfkwr4il7
8/uQ3s+edd4n25pcdlrlwkvTqgO/JJTnAPnByPp7gqRiC/xyGtOtjubTFTRiuJT3oEir2QjL5gmY
DFpW58S4FQGfP4SgQwbv+UWNW6gjQWL3pUHjWrB29+KOwvGGQfr5ZQLGYrsUX2tdMMLH5Betp40i
859z0wFdAGGSjaYsIZMnJ5wv46sSMAc4/bVlP+NwdWvvsrFoX6xuYrk1ZFtgkKp3dNRxaCMEBRBx
NUaUeV9t2yZeH+B3Zc7nBTPHQzSUvFvcvki5ZHPqU/LjdIzQYv/i4fF6Fn9SEg1Dj+mV+btsw5ce
7NOMnUoYI4A54GmyTnQ5qwjWrkzV85zpNyHYjODaqA65Ot/J2rXxMjQKIthJ54aHVMPOMaAW/ffQ
RIsAbXpFHqoYIXY0Q2JQRTKPCHkLAXSYAtcaNNNzAUPLpfcYoaqPrWwaJxbQUHHiBxn2QTdxgd5i
1J8h4++HseHWA50K/IFPngthb1195aOFvwOWSsPIEyAUWpi3twYUMrq1aB98YNJgsgVUqAhIGyST
FxLOMnZi9sj0sm2pAigIaM015f0FLcmuXlzMVNpil3LzNIYe0Pw4ANPqM3tAGzhsIv3YD5OFHTtC
8+YZxYJy2Yp0JVOiFcsY22i7SFYD48qzIGrgv2U+M9uCCwVF/5DTjt7H02itDnbUB7X0mEW+NXeG
vCYLa8sn8A+ib4cIKjPvMyo/5TlcvA5VowdG+35wz9AuxHn0mpVEWAw474blFoOqqhdJ1vsnkCla
lILbARUtm0B2QHjf7hsyRh8cW6rAzPi+2FicTmh51RRvs3XPaVpnMGj6BQEVKXnwJcLxlGIIkW90
Lkr7rr4rLTv/Js1DUj/j325TUnDrLCVs5H9GzDjgBY1W1sSPW7FvEJNf3ELWiW9pxB8bJhF++4sq
eAJ20jN6HdmHtytp2MWgeWWdZ3jhZPqAh8K4Sw1hg0cVZ5aTXBWANjK814oMJ1wpcfR8MRwCe4Tu
62xfS3ouDm51jGDwFmXfJYUu6IkiwyX4CX87vKrqkwwONnnq0qThHirlAEgvFnzxlM7w8Wb97zzd
mjSnaeKkWQG3um5k/PQIkXmVP0NrPWCvxgGDoem4EUow/Lq3Kdtndm5OD4EotkcYbNAlT9fG4Ixr
FBjcjycqalLNUtre3PnATVJyXhVm+d7iadgnGkC3rLruyR/8or9EzWX7u3MjIegrEzQC9Wm+vZwO
7/wa9L4M3EJZO/8jU4G8BDXTp5puCu8ii0/wOIEcU20uEPQ2s5t0tEscQRGQ4ZEVWYQJb/DDLyHi
O3U8OHDzgmEZOhZrpj+4KQSi9B2z1HNNxDDczZ4ETpFUuHZy2VEr9g5rFVZxUYbbpPM+zycwc4aY
7vIWiwY9kUipv/yTR8xJPgQMohHYDe6tIw2FevNYeiQB9mcg6sJ7N86fjDqzkULCQ05qCei8A8sX
944HxPpVbfVoWeYbMFKaFWvtmyrXbkfHH15CNTyVO6B1sVTPW1KdxBxiJDSiR2s3yAL9HnzXAFdy
LPR7l/Rxz1sIeH2Z5MVF7CqNysbeKavp2SIa4mQQFp13bnvZJO3CeX02QhSVpBUR6n7HFyuPNMct
eELWS7IgpzGvR6zDt4wf0JjQCnS+5s+wThelwP9u9Fneym9EmllVHMKO6oEpryy2e0EChK99bBWZ
yQskBMP0Mv7jXL4No9yrxplHQvgf8ytVaO6jOdX05tZbfb29lxjv7VRqqlmbTZaTM6/rJzAgRme6
tdMoA37OPdBRudzNwutJu0Jvdl0JFpYaidFp7/mPm0cdAgMruQMkVtUY9gzRSoSSw5jkbaVxeWRj
WoQrO3o7IPvIWpNEHwucPVoJR2kHPG1xWoF3ZzpxXNGBoCh2SG89m81fbOcrXhmvfV//Md6Ql8KR
uc1oVYkrRTQ4DJgmRBgWgOHeo9Mj6yL4i/WK3+GwlEYtlAjc6r0RyrG5/D0vuY72af8PnbX5WUf4
cmPh+XBASSgCRJPTyvmDO2JR8NJXz8dONP2RP+MsGtohir/SgSanw8rDmP8ivlCsJX1CoxjZgvnm
IPkOVaUInv5YIsYftNpGh5zhKdkqerwsZMsZSQnw44xNRJQJZtx14Toh30jc8iui7aLdwURiAMD5
S2pEnGx/QOs0ADp2HmcjwtI8+Dg4QxB9cHu74Kdys/y2UJHkyMu1tGcLWaM7jjxJUNAWCousmt87
xUFiCD0oA7Tjw6MqIana2dkhtwjjQMbmXbEJ9UDWIlhlO6NgM3Py1aM88fHlizeeviJvECRBdwI7
5z8tXdFrP31cJadR100lcHhASkCqXsLM8f3kYQWVfSZYJKAjxodWsn9SUDmbZpYG+da33l3ENnVr
fNo6pW9HzgzBvcEZGKJPEX6rUtezU4tUVrvFh/eXZNxxLpPD7U9AefCZT7Ac41U+90xw5iyn9fvN
EwID6p1TcxxqCICtV/NdXj5lepazeoePWbreMU3jdLQwKG5Ujgfn9ZP1AnkIA/s/GYj9xnGcWRM5
SA/ngxyNfocm/A5SgNQZ0KXYHSLA+38j6LJoK/KkmXbCHwD7cfwHiVbNPuhMj6t3JHXl/4TWFfdd
H/bRmjr4QiBLFBsnoJMWPLdZ6xXUhmnAB9qkdw6J3K8Uvv2uumQaKEUqOV8nKyje3E/okiC0AUn1
pYULcqT7/gAFWSHjpkOIIYcFt1oesopCX/lpxnENkpF14LS9jyXOGH/T8/s+3LOkfson2/xkh+3G
PCgUoxel3gEfQo9TkemCVQ3CW8C+g4jTGrGfTMESlbfc4TJVwqhb7cGBxoUBfonR+Xx9Dr6sF/Zz
A3zZ9CeYjqx7vB1xre0/nsWDfwcbI70algJrM8ZZzXODa29ZKuqhDrzdeo53wk6In+mm3Fj3lEa4
kgGBwpDpMZg3g1im/9puEf9YxlnzBn8i6eg7NJ4hE8h88i4lTYwdYJMDnF39xziihuUZWTUyU12T
mUPgmN9FL2AXhfH/toMWQxL+uAbHIlZrcuiiGJSowOCvfUBMQqb4oSCZbsGN4TYqVXdj+jQ0YsR+
Q2rPnjN7Fs6kiKf+cq392SRSEeBv3nLOOgRGw2KuLRJINzJ0HUbMterqP6nISB6blGj99/LpfHtF
gPRAgBn3h4k0/oVq1znlSwzPzX5wlNxwavq6WFa+JfcGzgWSdGqq/BvPZtjwcE8EPnHWdDIONi0r
v6Gq+D/4ZU7ESKz0ZPEib5+wn8567ccLaRC1rheQLaacaglTWngi13H1CfPbsXE2FXLW24+0vBJI
eb0Jt61u/yVm3Itg+9O7U+9UPx+e6qvdWCc0119ypX3SAUMg9wkD1DgGgsEsMxHSeCSuXv+2pEdq
ibRiWPmMAthrlT3J/WEHtohShXsa1kq1w+/SWf+58TlvO0g+ZkhwTmioxdNEGvxHaj4KkA8FyVOP
ip2ak4tQa1m3fjuuQ1qaNd0+bxr4xHkpOIB9Xv0gpt88CXJfoePib544br2LKmXwtfFKJlMB0f0X
RB9jKqht2aleUU/xQbGkr8PI+EvpLw2r0TPmxrzNNixsMBHZzyWhbxEVE2bLDPO9DwA250SZrnbu
oXlAzendEngtqsD9yxehjwlVnSTT/bhKJnaj0MtzCeAT3kvAv4q5lfNlSaaA703fleIDErolfTNf
gfcs0v2i/1dbWxfyWNIQS9O4UEP5AfJZxwd0meWprfNm/3/1zoagLDcDfJAqK4iBcvcyMgVAmj++
XwNbgGzSAMjgwcudgBbgc7dP3fQlWlUUIu1ol724UuTMrNY6iZ4ap5QGJzUZsMxiMgbKn0arjlm8
ssdwuHCpM6L8tIdRcXdaNZPRA0CVIfn914c/94xk1iAXTlC04owkF75i2Lm+NsQgNqhYxxlfWIfB
zx5upvlle4/bxVhr5kvxLFkQKfaF8CqyOX8fiCsQw3puD1s+dTlk2loY0rfH+ZDcah9xnuJwAqIr
X1R4nut2TCIMxCNtkWIOGRj8W/EhfeC4HmilvVmnpiwwiq6BW4cD7NPjJyqXLrGYlvKLeCJUS7mr
sOsZz34hlRNO4kxOPjPklT8h21HjMQffDrYjkTQQThSfVWP7RbAToszsM6bfWT9/FOPN6DW9hEHT
d0TU6WP1CKrFNwbBQRKaYk28OoViJ2NUkjEnRewDokYkMw80kclFjfC2m/Cmg25Vc9dIYmaTqx8G
UtzI+b3gks6eYJDFS6xZxu1NaqIqcbqyn6wx36FSjBP0iZ2kSigrkePYPzqYJcdJUD9lnyx3Ek8T
nZm6U7Qg4f+Bp7sLkgZxiw7vF8t5Nc5ImsVSGfwIxoJxahmNnVIVCEMgaZJBv5oQ6sFSloVzTfjX
i3kSraZ/xXiKfgKnyHMRSEPN+3omMel54Tu2uczI/APHVHmX3dDMzlEcMcR5DKq6QD0zfDJ4wT22
vindBB5J6yxJOu16FEa6W9aDRyPeWKRXxxISPnjcMVyvU2AqZ5iXf4lKdDMxtP3yw4M3cu5DWzeE
AHnQGuwzfAdRvVNhnTj/EFLpJB7iYeiIZPr92RQZtnFReeC0tDV3WWiPahFOu08JHXZ3XeLIV8rZ
+sUsDNT17DNtB0r7CY7TEOjEC+iCxyFUiopgodk6FxL8DmAB4bXZz90LJkvsZZJYML4F95oDCQGv
GDtaoYpzknqQqo6GfvBnWrx5gQD4MrKoAyitAtNOcFFhdSoOITvKFPXQL8v+OZ/CSIw6kaZ4QkcX
rmdeIuxuMnBY6hl5kSPOLK7yuXKtWBJDDEXFjtk/BrjB6RTsC+XeTVXGBgaQWzm5UUbKO/0yHzA+
Av7/9+43B3uSuA39ZdSnwgQl0suDhWIcc1/ecuwsIo/B8Zjcv8sv+Wa99ALo68T+PtAchzFfUbwE
qrwb6kWbhokAh0f9luGtpA1/wAaFOW3yijHSOq9Bs6CEoDbvlq3u+4kSASIk92jZnzLCwXl0tB6G
zrCW1NyqT4iBEh+MuB4unGx51RW+1NB27VGDEVmIwq8+0ghU4u/ID3pVpUPT3bCOpe26HhDx/Y56
iKtWr8V6qKF/YQYFZjFCWr7sXId3LrIR6iUIxRxIvps5VvtgDjixXpBb3rojPo7Ik865o7nRnRIc
GBzIgqbv1aVN6qqb4Tnndy/otnelfV0jx+a1yWhZieDj7CZk/KiRdQnr6TYOuhZo+J6r+HOBZXrT
MCpeMoGHmfMMxaZkZKK7LDGW5hZkZc2Xi6soq06D8X3C3qAcYgwHgkSuUNjwN8Zoeyx4nBsDRVYf
LgrCMGQmnKxSUzSKT+YC1IBjzyY2udKOFLtFKp24HfDgspr/45gtQpCad9/E5iI/062AO5d/pGxb
9Nq619iaFocnRVzDL0o0EVqSVPD8QmvOjrOmYBNB73fSUioB55ES0nboy6OpN+aG/6WwtCMT+Mjh
HxwLQvkb2OjJrBpUW1AyWl8O18LbHkFUPk7TLf9WteIV/iN/5+sdp7oYo6u5Ckfzm88WIMMVInBM
kUjrVrQRtAlUJlzYwC8wxVwIG7PcN7LsUTpys8NQnp4cCPZbgw9fVLX/yURcjm4yF30hqSwlyfo8
4dwTBPqZ82Hxm2KAhZ8oLNf79oJVWDP84t6SpCtL10oa6VaGHigeF+fJgqIsWBUvrP6FBWUAuEc/
xlfbsVkvw1hO1WnckWPYQziLgEMp0xs4HpAL0IIl15U27g3+7TQf70H0gnhXfmfuHtY7s1VzxY16
V0+w3gWCmCBZhiyTKlDM/i7jIbk68UCaYR+SODIa2d2K6sjJYY5kXxdcvbTZ5ZBnSpr/gGFOwNqO
fepxgJudn4j0rFUbD8hHco87Jqz6XFp0B2hRkaRAazZc7lWrUwm6Bk1z0eWjRmdV4jU9HbB8XGmP
e7MJRFgiqbCIjbx76zKDRdC24ErVv0nnnF2upKi9K5thwdocrC6FWiIEtsAxaObX+Q5bBjQIhStf
4GyH7aI50KSIEYrklO6nDctKX2KrsddxKTNTkITLPVa11/VG8gUPxZlCv+m4k7S9N6PNBEMtEzqn
JDW+eBkMNa1SovQIfvoPmvdewQe5cA3zHy7v/cy5vrXRubZEPvSlRM7BlfytcznP5H8sC0LonL1J
8W9r6J965NaZ0d0twIJbzHQ79Fq/ZRPK2uEL9/A0ZbOyeNwxCmrB/AolYqRjP0K1ED7cUMCFMjx/
FCtKB3gcHA6PKAtLRjKXtfsG7jV01eqP6/bOaoVsCmb7FHqAX5Q5EqMScahSCei833LbQG/svCfl
gir5T9pNgoKPX29nj1YM3gOxfQ/GHa8MTiKF8YBA/f1mJXeKNlkKiCUIsqrx1zyfBiWV6S0+lD4J
oJqT5I34QjQVmE7FR/fA0qtxnk7K9TIydkFirSyHkY0RIleaRMk+Jiqyog0gHx2BQDWvkGlK9hv/
QPI3iTMeNdCbd5JMaCMciCJb9pugB04NQgHY4TVjQLxhTLDfJ4LNchF6JBnElbHtg1x44tzKeKTn
2T6ZaPbLgo8AsXI19fD9vvvanijqaW3GLqAll+vxtXNMkG3LaObYFLgJAT1GO7uxFQoMq85Y5Hiy
p9puOBdNDV5QJaRc6GmAENtMgcdRpM36qHVzNh9lwsp813MUQgfewzJssn6gzrA8IjIvo4PVC6KL
2njtiPkbxKzBpE9Q+kTG8VjHulLCkDAcp7cCjI6I4hB1fa7Vo3q4iWrj77RTg9VIcqY9seagsGlJ
VvtpkEGJtM02wwsOxyfMtvQHp39cVNjYf339imsYT35f8u2wfeu4BTqasw2rLNI7Tp631ucfbbDf
k32iyHr0uwuIL5nUQm8shJzK7DxKLXDT/pbGbRvjkmdanv3CrTLkMUh6BOt75UVGNV4x0Pn+5v+n
YPuFi9SVg68SavmOAbAstMTuLNnePU+5WcCR7nzmjL2Qwgb6Ip0Fn+reXDNmbjXOSJTp0/V8J0Fp
F79MHBQOaAHaDIV6YS9OZpRJ9i1ZeYMDTz/TaypRM0NYgwHtM2bSd2lFnfbKvoF12DzzdGdnwBYC
PYDFHaloAPVHx737g53Mc0nI9znniiGt9eLY9MWJAa/fNH9jVSZlifYJWVbvRfQyLpwATqJFyWLy
Ufu6y///hi1vRBj8DFPd2npxSjOR0F96eTr3OA83HDb9i/GdE8+kkZyeay/nSKAFaUYX6QwNREiu
Lk54QAUqTJ1z/+uap0W1h9Do84d0zQ7McQq/d+9gyw5OF5R/Q6hUdJgKmwvel6nWxIJhbkVODG+b
hUpDrwYwfh63YEnss2nvjJ3plFCR9mTQu00oY+hdbHSStIipmoO2gUtikHE/TTncMbr+ZmnGM1+V
y5Tb+qKmmq/x3eRHM0aeS5p45MQEMNY41MZL/DGjH0mjXLtpwIfkGlFkFWKwP0PvT2sJPAyee7lg
CfiCitCtzON4k21YDv+ppi1oVgKIA4MFcM9H7sbQvdb49FG47kf0Dp1ptfdOAoXSc8UtQMo5EZ9i
ORYROK18e+RKZm9QGWDh33GcIiw9Dle2SZhHnpJ7v6lLwhPCn8tPOx53EVjb3TzOG7Y/4owLKHcs
3OY9b3uygG1SsKRA2rOyucT1zAm46flcqtDRHVQAvlX4zpj34hVcN3xFC2qETl8J+FcO54LwS7CA
ZNqZ8xCIRo/Ywv+ow6hwa6oXUuFan4vuWB80kgsynlq1pQ1F9kZPkoAKb74xNwgE54QTajNZm8IW
CN1KMXCpXMfttk1dEq/zzXWIjIpMv61uz2HDPljaRdD3ov6kCSyga4+h0hXcFDbUbKfbuq1npyiq
0RmOwj7W/sp4/Iyyjk7wF3Yth3Y3aXeRLpvyfmwzvsoSgLQeSwbDTrGGPrPBtuIiXPe1KlKaBMH6
GBqTn6dvy7VUAIiLPqgBE/RWTyLLvvfv4uNxVjyt1TUDQgp9WhJFMjZyhMoCfn3qwEBVk099AUhs
x9fzfWrS0ZGxh03Jx1fRJ3D9KGlcV/nC2EsTkKMpxcRBn/jWH/glfO7kqOHiIiJgvY4fBwqjHCQW
R878nAJwAfVr5cddSaIquB9MQsjyB8hIgWk+tjrbbgKCP08mDMosx06TnAsBFKJpgnUeHYdBLmvx
IM5ZfnR8qWuQP2pVVfPfOFF7zaRO9OLyv+RFLEctckWeJcgvNRnKLkPFtYKu+5ab0FIICRxtF8Gz
5T8lKf33orC9SgQSyba9dxEUPalF20mgKiM0YglWm8Vaozo5u3lsYzxZSsGbgRg+B3gYO2IDoDJU
0CDwhcb9GpluNsQK58D9SEofSeNk2YkB86mMmWbx6Q/UinsvbPh0w2vxfX1+aijD5CyZuGKfUavd
wAJlehcsRwJe3TL0Tws2FX0Y0oFN0RQ69L8TtaKfzVH5J2YKHTk5kJJP/m4XrDdiVDs6BpHN0UgA
3KwdkDLcs7D4asdokym78+4MPVJrsu0ffm4xNq6Z9nVQBcan3hFmxm7v96jXDb1sL1Tra7InWr7h
Z5xDRgpPOaPakRrLItGaf5HZqR96YUiUY+d6+uTM0N3ka8hUHndXiU1eF9KcrKRewXyUrUrD2PTH
w2zClJJeewzfRcwcm9yke2W3OlBclvB6kkFRyud1GOJlxKl3tNXfYcUFkZyG0zkMsmuExL5eBp50
HSDSjxbBmYGqNpDeNK2Xis7MFPLDKnb/QSsq0+CJ37Cc2Gm+AwL2HOU4L7Sm8gwa/oQwjbz/B1+P
eiEudPVj2A+HdAxaEqld6OwHf8oxxUk04duCZOBSf3+LKfvTaGKgyRf0ZwOByOkTWjO+6jotVaWt
9zjv5mfQg01xzFowIXqlb7Eq2hBMTll1S76WeNr9ZH4TWupXNkQ//M51pO+kxhQW+Q04OYn4kepK
VMug5kkxJbRJ9E08dJHMFTLCBn9qQmnkVWDHRmQq/4ATy3oXyGBEhUnLIWTsfeVl1vwSHxGE/9zB
HRqTukw/BpIc5DoUDuRMlQaCeximwS0bAz4VCozYBqSxIGvlUUOmH0W8o768y2eyNqe/6UePGafb
VYRKUjk7koggk2j9hJo2eCt4r3kKnguNhq/UWnwqkPRc0UEbIpZuDE6OihJQLlxhuyOf/RMfw//L
/PECeO4B0yiZ8SDU3t0KWhGo16dsGp5EoblU6JBpnG98eHVJqtv/cnoWf52eW16YwlBIeDfHzvzV
c6K9OO4EmH4scXUzYzS+/CdIap/MPqfQsCTw2TadRUXgRZUaT0RRxN/MrNQYC65XVsz9NQ73pwab
WBbR5NvIFU9C5V1C0TsNwADJnJo/JEFSyqz8YYp0MUqCAzz5w+3LtJiyl993wk89GrC514TXPb86
iznDKMLVzD80ikarxXMrXuE499dWZthetGrqUTYIHfwgDmfdtCoq4DxnMssLX9P8MrpN7zRIig6b
415ZYH71dPlnrN5Z/XJqnKwBL5M+lEOW7nB8bPAorFa1fgL+6ayTssOpZseyIIFzQJCFiWaAh/cU
Urwi6zaMbA0IqpS5t1F1LGqhlXZ4iHmzrC58wO0uczgbEmI3OsUMiXC3/kJamyLOgiIXs5ELGoHT
H0/6nyVtW/H3gakbhzU4w2IvzisqaRg+SvADbAH8CEKrhGYRVS97LK7XaqDnixVv8Q+Ep9d1dm5D
4YZfiF3c3RVMss/wcjYqplEhaHmfWJ2xVyRkMgr/jyTbqPWWRdeCwLtzchuvZYonoeTz1lEhGVM4
+mCxXF2nwInV+2VV3D5+GMsCWU0XJnz+8fouD8oBVP1BXuSGGvKSqAMxeBlBCdwLHmWP4TnHDHqN
0l5xS6hfNj0x/7/42g3oW1WTN/McxeJbfmw4ep4fs0tL8RaLZNRxnz6EBCbzSvIQ6DHmNZGuOqXH
Kx+P+z4itv1AAPowkLB/djvk+N3PuivUnYZiYFWkRPRGRgBI05jzEaSVRneRfdhQuU9TZqJXDtqQ
rViX19mqsu2cReP6edlgudxuzCo5Hpw6KhfhkQarHt8LSqaqujfQpNzN1l53hHlb/8nq4ck8UM50
gHGlvN6iuP6gBIzMl5MyGWjcJF4miolVN+6Q1TxOrN1zwfqRt/jQ4zcsA0BefZrPCGFwBoCwQCFI
vwRRt3n01lETmxgLNSXE/4/0bQ/gVT3f+3hwdhWrPH95FDM1tZzgXA8XEElyw2IvSkM/+vAVeQz6
kIxV3v7eMs+DekZCMubuT2v6AzMkwFwJW2yUFUDEf9oLiFCPURr9LmIHCqerSoVQ7aAQdmZfCa/L
fTJf39d6NnBgB1COHrfYqDptsDHNv8inGETKN/+qa3gjEo7etXx6BorBgOWo+npbQrFKbqiLIsSL
cUAJypCnX9yLDk1tSVihoOxhvUymGxMNzxXHnQJTKIMZnC7emi7+AyKeUkk8xml+BGEw6cgFpalP
tvqPCwUTwPqxRZ+vYkwQZK4m1D+safg1gWKIarvFQGQvqbpKfwuuSnYxzYJMd2gJ7dgRr0ySPN6i
7I2Oyz5zsb8D3/5mlexKROFejyMX24NEnkDmrgqKTzKgejgAn8lXutTmMMmjH9pPhP/DICl33m8T
nsWsrqgIwLdwg1L+G/Kc3dYnDv0PgWGQBfY5arg/ig1lVaFkYyoyWENT2K50TQox6F4IjMw353Qa
FyNsoFrwwUlra5RQGUvLBWVPBr5HVc0IMVOf/R8CvkTvCLSMsiX52ifQEb+tX06J354+VYy61W7N
Q6QS66+HHGP0tMiK4A95d2UDNzZVuYUlHwxFzMbCJ+FUrLiDbu0mPzuW+LQuZagy9DGgrlAwQSjc
GOfjEEi2QRPX+LQ/4A99ORdLVtioD/yhF2fiBwILPppe/9/PEfaDfs5j95cT7wB70pYUOMpezw31
noLVJKjyMLSaDIMEiUi80V0LIaGtFTvSJo2UdPb07z9UAzLuMetdKu3cCXJlabFLfwJCCmvUmlgJ
2xlio7zWP4AfVwMpQLf1CMn5E4yltFEd4QRpfcC0O3zHvHnYSHTbUI3b2CZhEF77sN62DtxdMog0
4focL+Nx0MN27rm3012hU135o3WUsCVCL1ENOR7/offXdjfWRCj2D1VPk5g3xgsltFKmPgZeE28V
fgiLScl5Lgncn9TQqSBFPXFkx/O+uKdCGZFfQO8YurnhLbYWO2QvXruy6EItXf2QFrwHV9Iq1lg2
o37QWFtCTSnfwgX//CXKMNr1iAaTwJBzr4ty8ss15RiZ2Qe47UKUOcR5KiC9v+GmpSye0z/YmPRK
h4EBDD4+BP389lYI9GyeJkf2ValVV/IWskhQeklNiH3Csj9DrxvXc65i6Su1lIt2R0NlFI/eTngH
ThXDoy1xBqsHC1t/saBC2PddifCgx9NZQ5SbF/gLTvXkdzlqJIHwKt1DJN+e+lqHL2VlUlMTbroY
1NF9JylmZKBPfQOHIZz9a/gfitHHkbp2Xkl5Tcnji6K7xP7CaZwIYUETrOJnLtus80TW20A4AR2t
psdUviLV+T/2L8Oap5wSBQ851Mwyp3SftdQC1ZyMo6/7OomTIB3D2f0w9V1FCyWHVWWIXmgQXFa9
aSfyouHwkH0gBDnhk2HonbAbjkGgEN/tJZRflS9qpAZyhTne6VyWHZ28SM4AFKuhbWW81Vg+L829
tEZlloSHMv6Yo6Mcf3/Da4Gfq8JpIejMx7CzeJ4mj0ACYAI9xkb9plTL1D5As7ZM8aD9mWh7Xdhc
cLO3+1dYpd4lFxpE7FKihRTIHg33xSMwTPNP7uTZ4zIEielFjH19fWBtP9WGvcb5uJAgaWjgf+Ww
CF67a1yb5PWS6lGgnGiV7ab2hfVqEgA5aktITcgMdZSvaSxLqg960lb/DCrhN/lekbAJ2nwJIzT3
NeCMZHPM+nvsQ5QN0IwUi+RD1m5/0RuhVbqUvvrZayq41W71s8SU1u2InJlHlB+sKwSuVwD6nYcv
kEPPuiSeB4Lcgsg13/9nOftgE11QQwfhDISRsaTg1x7VrbQBdL3Rk4VK7rQNDp74FmPI8zYeqytH
YUYpSivsiJFoTcCoulmEUejYP5sEszF6vhSbCeL5Os+2KkOaWnVCNEKxJe9Di8m05oYXL98nCcVB
YBlJv4zGROyYF8CGqmKRgpICTHTu7RZAu4Lt5a8xzLBSzdePh8PuJ4ufI7rQrbuk90m21CacFaWl
ev22y/p1rFuXW9qtqJ4VX1DerXQVCR2rMUjOQqFgqYNkVEwshLlrMqTD+JA+RTZcOb762hsHmq95
AF+4l9W4nVD56gyxfHor1+Oj8kORCiksD6I0SyqlfGHhAHl0R38ofnI6YBCwUaTaukjYxyOYX7/m
lUDRpAblAeJRPVqNQ251yUNLXfswhpv8LlXZD3v6oRU7vqYGwu939ro/0wtKkqvnTBp44iy/HwI3
PT4W8aFWF2rDFuKJ4YIGV2g5nuL8fYsyREagppsSvsTkJiRH91fNuFx/OcBKS9nxSIRhgqOEVex3
Bzae+v12rzDm9lTq2sP7UmyLsWVl365CpmPwdz5XdY6VaY9SRCSv7W6A/dQ9xgqLMzJemAmLbh7r
wM6R3vv0/MGejopOwd+TuGUqnW4FSmMpudGjOHflYl2f8GdSCJI+legCQe4ztBeklEEbpNmgaV1f
d+y/wX9G5fkbO1Hcb5JH6LQ3V8fX8drpjmeFvtBwSRxavSxNqsGQpmmTFFBzzhfq8EbeQTV2fUui
uYsg085kuK7fugrLwBgZ7UxwDrNSYVq9S8jNGQDacJFtS3XFGDybEsEwAvZ5XBhMNojh3BYX+tZf
PaOcqE49GKsnTpUoiFsjTRE0DK9EWNgmf0JYjADQ0vipdHfi884if/0HPorq4LGxkfJ6pru8C8K/
rLdWpeub4w/oneM6YRkH9XvlCac0092HK2w6dzm4SF52OoDWqezDRwik5ik3yjZ7Svr8vjPIWrIa
ciRaqbNLNedC1KBJJm+5xa7QNAsJI0fcfRW8/cNI1yV9TbzsODGFWcRL4E6lc7vPu0zG2Qp7bxs8
RP1oLMH+uza9MyoBWhG/BUHbrCCJRDKM1AO+ZakS6qRMJXIPd3UqQ8fEN/FKlKy8lakzcGJ88EQJ
ZBLv34CnSFtKRQQTyvHMsX7eIA1FXGsezq3P8fFMdlWGS/gvxvWxPiUpoJOwV9JzvwFp6mPdMdeU
FsbKlg9PVKd/BSh/D8NE/tv7UneHKtTtJQl9qzksPfbf3Cu6EDwP71hQzp5LGCzUCYb7FnAKAUVa
EbXT29Vo9l2XH3qO5fNoLYzZ7isfkc2rVuV48aQcKu2pKe/xJHpSYo/8oAc12gH1v3rygoo1nbqh
g24/DP1msVDQgmecOniVCNjkmCldZWFGF4xrJhilqiQGSNZ/FA9PfDgpnSbgwW3MmySJhzVHG/+N
j4EwH3b3vUaEKi7Z4wX4e/+MVX1eptft49+InAT3C7worp8U4c/b4mp1vtlZmhEAYuRdeZMQSGQR
DpuSXnBSdiVDr6uGoaFmDgm5dqt11rd8UneAahTjNFQtIQG4Hp8RNXDswpT7UC+bI2ewTsrAyxhX
alQwcAxFBVIlJqexh4cy+XSl4qTQ2z2X3cRH2RGV70oFxKmnFXWmOu89wh+X6unBEhQW7T4jlnw/
ApQRbnOlxczyWOuYpRWf36fMh3waOZEil9cpIeCf1EQjy2v8qSFsljHxt8utV1r2V937gh4iiVXP
eU0D4i4vODsu1s01obPAZftgeOpTe01TQ98LL8EABKQYIvRYDsTa1cVjD/pvpt3UnecXlQEuzDuQ
ejj3sV0vX5bP0TC24y1NF5lJBnb6GbiELM1o6z3BAmIXX3KZR2Wf3eonODiNKESpG0nlrjB8x7a9
gq93dsw1sEp/zSIVm+F+5tos8Fl/+sqLpnOtfreXeOTWsu5Xz2hoPOOo6JqlMxD7EyBi8I/KYTKS
eunNJs5mg2N5jfK2glUiotm7dXYk5+TGyY5Q1qDT9CUqKOFKI7k448qO3yjLw1ffCQm/r5KUQ+50
QvRFu+R2bBXvHQBAXubG7fKuPvNCY7VQoiLvM1qvI9bYQ9k1PP7OPR4FOO3PcS1uEicjLxlvQy4o
GW+hzofW1hJbunPwVZRmDED6w6Z+BufebRvvEfcR4wp9yjCwS1j73ih8UkMCgJb/fFuVuMAFwRjs
115TeaQtWHMkPF61oTXNhZeDxggmAkCB1qHe74VJUt1sAe/sVhFSej5ORBpcvVvzYeZ/lIXT1gH9
dU9Vo3PQH/uI8F4A9FRxwA1lGj8VnagvlSbtoNHJSu+N3UGDLhCSztEGRagD1c55FAnHbeBBasMk
4EZJ+nlg3/XYctASQVpeZKs4C37wxXpgZBFOaBdWkBARxANqPKSIanQ7JeF9bqT6dtoln4g+DLKd
4Tu0uqwmOs2nFKExBlkyxwMvXpBKtZ9l1QAN/fGLKAMbe4koRjl9Jnqi/v87AKRPCj0qBUaKP+Dw
4D7A4zjHX3pLE0CYkZiAN6JhdYDegKvX3/uVnStEbN1PuNmEqWRe/W3WF3b7kyis3uvFpSSevTE7
yAB6QgEwKftPMhoxiA/ic10CS3PyqS7Y9LEkMJfK/znaw5YIXK+8ozSQGW5o9UIeeIUd4fRl/44O
bRFqnyAPT4cay4SbUgQngoaPzJTjjcwmMNkPiYFamdNaOiF9ri75SI/xL/zrs/SYWFpTWNzD8WET
JYytvEQg77uQHuJjXGy7BdrkfiK6v1B64L7ldOcv4s4fH0vhL2PGH1twdk1/tYfMneUyH5o4MgXs
re1JPFt6ebuk8gulloOrCJaN6pZ6ExrLXgRZ+LlZjsKkZRTced4eIgDbhxrx363jK4NBzFD/0pHI
nXqFkVKaPw0O7yKedFnRd/J4mQV+/2ElSENNt5F34BxcsTcpwCprXr4bJhFQH6VZqpfKnGbjYkFF
2mGHSMycKRHrUdihiakkmJNjZ0w1r/K+42GtKkP0mhAYoiaXdsLQX+FXCEwKtYPNUbIZg9oQ5i/y
k/+2sF+hMHFGzIJeVnqj5gn3j7ESEBA4qGSE/TPA7gNBWr5gFIquxOgWrRUplYYZYCdgfOGlk6b7
FpL1Fwvt65vMyV3yw94qE+vKUjSGpRciCyo941qBzzpNkxCOKTCu5ODi+d7//CaPKiguI9Q8R8dd
aSmDTPW3IjUIxftezSulOND9j7i5GGynTM/AaX/gpA0DCzR8Uq/16uavzSxmybwMNZrtCJJeqTw1
SAMQVIk440hlXNmaqSaPmG7F7X/+Q5eOAFDsKrWIaC5K/gx0dYz5UujqdO8dADLw8Hgple9b8R/I
TtjgbbCMeUOcAeY9er9h0EgqaOioDnHr19JGa+ma4HZT2Fc4DCr5gouJrCcaB6m3y0w1XK3Vcvm6
80ORIOE7iYQXCyjkLhgfnmRiWpJ8oZ31ipZqMJTkWYp1S/6HJz3PkQORXpiPiVkpjN9VeW/jlrEH
bwxwVJFwaIi+qRrjcMuT9BrsPej+PBTUu/hkLKT1Vomxktj8MnSGo3c4XNorbv69zEQdZ4YpRLw+
OyDGm8DFazK8hnCVzSb6huCejibQf+BjCe4kIXIIzFb+Mj8gV//tXVJuUnVzd6qRPDCk0jIi2NMV
GRnJ2VAK1jXP/+VzTK/POND2t3zFzNe3azNCK5a0pN6DrbMJY/AKestL8cT7sXtCS0tO8AV5Xy5e
1wkbDK6eaIMnqnmC098o5uUw3vWENWBe3oou8o/TPGGcWZMADaejxySriQz5l4M0CENqCvg5a5HY
x6PA/LlDWugzvJ4l0etn5yG+AJU8bvgCA65qcApTGixrs9oIIk6LAMqptn9QVZE6k32xIGlX4tzP
hopJiAFqcGO0vRhDmP8xmuE10KCegTP6gnovewnCrJDBIJO+G0S1mxyJvx2LefFcw9KKS/d8BgeN
z9hacpmyfc9EC59CAqx0PBJhAhETi7azFKfw17pE3YRm4wx/rRKkNdARLivSBzeni/jxLajWuztz
6WuBANzwaje5tbW1gSQ6pe8y1LZTg0bQZUtiFMUiF9KaWbhLHCmm0l0+MTcIKL+rzk1HLrrUgMAn
c6qah9LNICRI5Xt/+i0ua2p3UP5dRBgbwGTUkh91IpxbuiwjwlWpMn0zq3xtUdCvx88BZ0wsR2Jt
oQA4/UO83+zLMumkrAGvvCUO/YGZjMGC07qvxqXxbAJ57K9y6YbBPlO1+VXrw1146dRXX+rlAXxR
grikQeq14m6GWsLc8zNBS5HRgb7P4yjt6yg19PWG9ogJITbPYhu61k893Vkx6h6vAbm1YsItPucE
c5ZpPhB+lJv3lc60X8gWagqPoW1yxzvbQf8a1rlr5OUcjrv/HeVjLm8spyIHq7BMzlRWTvnngvo2
eXOYU2u377sbdMsVjwv+n0pInNP1n2L/DRs7qvXBpxhCVoPbFfJuwVBkA1k7LqTH1FvjCGil3dI/
WRb1vn3cZ0H59a8XXlkDU4mpSFEdM/rU/begVCe6I1H2KonJvdDLpQtEnF7tFBVqFYu4JACaxKvr
ksFmOunPJG9xwppW+CVZzti+6hcep4px8jYTnTDh22BpNN1rRdd3Sv26GL2q7leJUlTB/faLugmB
wKA4g7fRrFewGlJgZe1DgUA/qcEf9rDQ/J+u1LxK03rBqXyj2bS7EU4972NKUz+G3/9wy0WNDJzq
iMqkHA/vjAnnRnYppCG2Tuxfxt0+pfVR44+sYfWtPoRxVz/tNu1bbLmcb42z3G3C6PygwUIBZGSz
S4nThREmS9KuagHoS07J96+6YGa/TFk2wtWoK5Z9ycOXtbgAGwGiDXYro1KI2WkO1R3lM1I7/bhP
trxS9R9AV+E16TDbDfmtF7cxWPKQWUccrvp0RmZojE1w1W9JzZNHpdc2B9b5N45y4Az2PO7vpOhS
A1b0wweWimCRax7E3FFvfcOBYa8NjbQSna7BK52eMuXjeaKUe/Bf3q4TbKXgeYI2SCyMaj0FvzMH
c+4NNgoc3Gc/uPxdv9u75cBKk8khgBUETndZiosiE8f/kv1PAD01UCeEFm8nxFO5uXgjKk6Cg4le
iqtKUkxpaHYfJxjunc2sZ0TkVUBZr6wGeDC7qwBcO4C0e7OX3zbPFyjX1r9XFQ6ieUecySyZqwn0
xW0MrzO3Xg4AZqq4thrjDWPEzZ+fmzeA2CLDVUGOW1aUdZSbIK7ZqGwvE4AcibYqsGsp54eeFEt7
Xwni7ZuHq3HFxGsXlyzV4oCvchBQOWQe/K3ZSKL/bWVBDEZuYKlH25Ddqe7NTlKm4zKtye2emw8L
trR7aJZuPYUm+rFls7VRYsc9daAI2DubYk3Oe1YSxNoIoYTm7rQdIVUk9XT8J6N88Z1LQquoWWJo
pPPNeAbRqrcYu/d2hy8lq+2/fU2txJURD45wyJf5lWG7nmfWCiIijp4rQU77UrCK2Z/BvHB3QVVx
WI6cfVtNlrHUqsrYFR1A1NPV5Rk0PpL+OVmWxvKWlnNHF7v32nFtStH12YuztsWIWvZ4TgAby6ZX
AG/JRDzKlWncKf+rA4+htHxLx8njjQ0iiQbvTg7klUA7DhjB/3J2yiNtaz/Bmzhlc2fADKGzOSTa
28VA1IZiAix750kZkAdo7wxjl1nTN7LBAqegyckUVnTH8sffEvgPiFMLf/6P01dW6v8OWwSwLCMu
xbO7KSkxAMsis+3qnwq/nO1wQmjTu3x1/DN8Nyzj04+liGMIkXs9FQHZIpJ/lYfPZZdhHTGsh3SO
9Aopg4ee+7yzhyhtarsK6juUW1xbOHaWgRezfiXA2aHFbi4lYGvPw4fbmysk1zsnNkmziDndUB+G
JZoawG/hILrAJrZyIdj7mk/gA3yPlOiZ6R2UQqkh5PtHRiG06+VbaYJY+ciL6+P0T/EZ5bWIcnJg
wDu6u2gSOgX4/zNGczYbpNP7Zjo2K/z3uDOVbAjEr5POYECjzuEuccpz+ajvd3KW/BInRLdz7hQy
Yy093UtOfH6w+KrMzheOGlQ5VnPrKD1WdPZmou+gQBlHRFnjvTqVbAY+jIOdKD/ZdHXRc0Jrbm0n
aIBIZR0NiOZUUHudJQtf11Dpz8fSamo8FuTB0hw3YgpzZGfYfUyW281uH+Zk46vxbg7WanV94Bnu
4eL2TfXVIPADpdBadm5Gj2IHJhJtda/KKuQIF4yUq8iBw3S4JAcbgVqxKNbfpJpEQNb0kMw2Ug6S
cHeuyT7u3XiUD7RRs9snJ+o7fpI7n1Qm6ugxNwLcC3ew4xwcOgxzk/zBFFV0hsPC0A3NwiMQ6BHI
ICo/ER+m2UjCxKEe+UmPn1zTwsFfb9KBhDzFqTRLlf9bu3SyOPo/L+Jj3AQN91YFsgWWZwfK9He3
fhnxaGyIwzvOj4JtGBPhmJ6o1hZqGWoMYwZyysXFB9Vk3/vM7DllQYWmMPcnKQZ81Iq8JcmUFu+j
DvSbp3NZd+eOd8JA11TDtl3Y2Zv5UhdHxfYLshHKrongaQin9EejEU3YBGLKwwgGQxuh0LY5OrRR
ELnlO3dM8OBvtsQkDmx461WcoGbdM9nFmECIAibQVR4yJN9GTUDQ3+oH5CguK5hRA/96a01FATtD
eylfew1+bRhMCl+Ht31JQ0IMgpifPVV/XUmadWY7u+tR06XkZx+JTi2SLZOH1gP86x1tfRnvyF8p
KXUjRmwndJb/JpCX3yj6ZyHNnAElj5xHVOyFxJULLR7Ksfr+4A1uMuY4Syma5LtfaaUiDsXq8TKq
lrVyB9X9J7PIZ2nC/hV20RATLdQwib5GO2lQRXn17LesFfB9jxkpE19bzxZkwPC3Y24z6oIcl2ub
eE2uNJkDqPu4bCeANxnEhPmiZGQ1G5mfp8mrZdRTl/zVGvypl0nQCOID/VO5k9Ran9mAgjJVtRqa
f4n6imp7z7oLN4BrM6tRadhdExTHJ/ToxolCcw0AbMrGNv0a6vgTp8aJnB/7lxtCSFJPBPJ5x8o5
7hXhkXehTTtABnfRhqkyNBq1fQ4icD8tV/hgiI8sMyyftY31FULkwbMbvtglK3qnIVMTvt9Mx0VZ
SG0rEkCtcR+7HJUsZ3lrHihM/BdrwrinDbn7LZDVdy333b0s4pFtIU74SRJbw9emKXO9aooASp4m
ssBGDaTWknSJS8x+/2dyQFCvHaR8T6jMwBuOnOuxJJ+ynSNJlT2MZ6GdSvcNlIUtv3PRvbxVzbfp
lJtvVHettzhjudj5HNY/G+0JAXWi8e5hT+AbRGczpLkRKi3jdSlsGD0akKrW63UKso7OmsoGoPw+
ppyn5seiISSBAodhZWdYA1LgbpKjnoidrhTuNhrfxzsOmRbpT0AfTXMwVHZpb7F3wx08nRGcB/fU
lYYQi3RVlj0e/b4mWS/mw/GKB/FvxjJSRHT65jI+m7yYUfip9r36Cl/pR6S9+VNOFWhCmlPebdK5
UA6TAN0OWPaZDkwi/Y6C2ND8p8w972JxFP1RyvWs58KVY+zCP6Pi9UmvlTF7Z8FGnpFweGD4rbnM
DnlAeuUDWH2xSIpFCPp1eeqjvwCEHNVasAo8CAghtlshX6YSKJ0yMk6AeSBjj2+qqVU9k4JGcrLm
oMxElXEBmUxX3+DFXoZ1DR+p1lBKCQMEx+gARqtYBE8ZvnS58ysfl+XD+y4YfWKww10PvThqzBhN
pGo1mCSsTbAIN2vIDhloe7+sb/yjmgKRzgdA/XgB14yy+igLpN/lPGpRqsqqxex+gYNzY3CTOap3
H+/srZlxU6zYUbQiL2xsMG5XNlaBuUnNGp5dwmj4O65iQaIPWdqijvWyRdRHbGPzDMHVO1F0D9tS
OON3EBQZHTJ3qaSmZI6E7p2ygoFWfRM6atxlbw0Q2yEfSKMb5phJjG+nENWn9UNAeeozN5+skkjV
pyRZywX73UrFPBAZ2P+w10xspO6ya7bd9HDHLxQoLtvzsxVjieUcGnGYJQFMiyYtAyCzbA8db7H4
Uy+OFaQDv4Ai9khx7RXoKJEDLTL25FHwspt2vvFNmCCq+mKk6q+e3SM3u9htgVRFPZIBmYePD9c7
R0QPcSLSv8kZ0bafJ3aG1c1xi+EkE5siuHivSkWUagA4vj4luaszaipBjI9LwWzuDDrf6UVKkMhp
ksLS7JJQaoFu+Mcv/4+02RlpDZ04qvLoJG+sxZgMLPXdsFjAiOTBSM0xnm1k9Silz7jj4yFUBJm0
Ya302Luima3FOZ7/DU5L6Lg+3LWE9WJVVJcDYkytQQL7A51PQN2cYn8BvOip+HFtY93PwcddPhbi
qzRyGXHrb1xzZErTo/2QmID8BCQSD3jY7DhJ4/2ZCfcioVZz8XTqYbdYlqkIFxfqdEZutSgS/OrL
UJVHv1pen/ogD2QQ3VpY3KS0BTXG8W+ivtokHA6l07G77BqWhWo57x2xrn5qI16iC2kRbHxwLxu+
vSzgO9BUnXn6Aqry38tJy5e/Z3w2koE+bU173LbHddbuMCCaRs0AVgLv+GLcC8hR17coY+8pdS4/
V6SojRF/OUOZFjBe/PbPZweWahvPNbOjij6eu4VX7mjFUfCnBQABLhu2V+FDMfkHfDQluNTQ+7pi
s/CV+xx21y7ioOyeGaUZP4rtEoTL3XPDmuBWLrUm3+BaP91j7AYhr89Y+DFB7OK3ea1ULqko/U62
b8obCC7xCIFO71Dd6pSqMu1h7LZYHcvwDvwJ609to64ESbCZMPDjhMvaKONREAZ0zF9OB9xBzTSW
KlgqKh2t4wAXEnkb2HVXBf9ysym4k4dvwxtF8xtiALBzAJRniZQzR8Vc4TuLt/CX+KIUWyvhpRiS
jfxyhvoiYw2s4sPIfpBLekkISjAGiyvkpgZCPM83Fzlf+EDE7IHru8cLMGiFtmSOp4jOk5Ve+Bwi
ZmjHaCsOnrw9Q1m/kh5ev0rTAiglmZdgs+zHdcLS21CZrdgjUvGYet0Vqy72pCZFVmmaSgeNvFNJ
DMNm8jhAijj3VWQEzRV7dsJmcaHDtTlUxMxTY2P2kDbEjs/jfIm8VY9FG2yNU2YRFt18gzIU82dM
yJyxplF3EI1oLjAkFYc6uYTVR3E1wWd5jAlgX/4LLshx+gN8lab+pTaCfMFqCLlJVtGGAb4qyZfX
jznI+ye426Mpcpklmy+4/K38ZytBeDDLm4ngF+L8hgSKssSPbrYteTB3WIYPfL1CgzXapGtN9pv1
nQXhZJ2uaa/w6JS/vEJvtzRcgYBXp5Guu4A4cimOTFFzSgo9bymAkVTpqCaEYpwtyoq24bKoLiT2
8mN4xOUreZdNMMjKR2i/7PXVzPYfnyRHCVqyHBN4JJE7cYsBNEjhWhnfu/cJUjDGLQKeAmJOZuoY
5EFAWufVFj+7BgF2X4yYHtf3cYnwLCoNBSUaqyB9tqP6qyv8jLVDCk7tu96CsRHxAQa39lbA5S6c
4XW6jdjy2YFHJDEAfGRD+Axai1DsH4RY7ubpwFOa8FcUTVXt0vmDSquwhbV3Hbfhw8BdeFUfLUhC
05+5PqGziR/iqIvSa/tqiUkYKRtAGx0y5/zIM/L+rev657wJ6s+dsFrrFmM5cjPlhmqN0Lzyy4SF
TDRRNlVlJYrV2WnDVOxJCZ4eSL1DJQeD9FceBGOYQ/HP2vVFNTtrAYPRRWQpMPCrzBhey/IxfAtx
GWN4znYAOLW5pVpmlr/E4nl46VNY5j+fKYTvFLzIIqjnu2xmF7aA+DkYB8t8UF0UgD5GTSJn/ZHk
MocyZbYD5xIQtlQWKnSozwUy5QJxWd2kP+RG0I6ln1ByI3zhXrNa9sqqSwMfDBYLLnIUnjlB0rTl
WqKJ6asOaN/0ixbPlFaNYcwOJyJf6QwKHYxseWPJ39LzkEoukm3SQC2rfxjOiPrbIJVmUvSrf+mf
kpBCceUYYocBE9jyCSbNlf6qsq0vSy0YkIp6WQ8q7FVQ5Hhnul0iRefZUHgaZoBoD1sUl1A343oX
P81rs6mZseSefV27JCnkdhP5zo3Dr948gbAJ7wMNKSaqOYAXL9lxcT4hz8Bxc3l7Tm4MR5F8biNQ
/C3LxQTyGfZK/IRfRRn/Ci/rjFfrI/nXz/zWQUOx+sFVwD6CaP1ys7/FMzbwW8NoLbNCRsbuYKn1
L7X4uJK6Sr3K2SXEMeRtRKG6CeUoDIqB+UpHGTjLpCmxII/HD7Ze9LMqiF90Wt9ZEQLfVwK9SJVr
QkGKQZNas/7PNIUyDQ78uJq4jsqat5D9ll0AETqlV92xDFvNRKAdw2pvVwRE9x6TQXsexB5zN4hQ
l8eEJFvGke5xkeZqEJ1iL//6urw2sh9mjZWIB1Yel4kPA+q9/DNEp/JABwceOR3YJkZr96zaW1Gw
puJ6kRI768lIuvV7AE6I9eT/wb1U8hC+8dyYDfrR2SX9WJD2aYyyQLPpNfXeXpLc19BEmApV/FIg
IytLT0NjSuwpLVFy7i2Wfv0KoO75HK7n7muaHTps8RdVGgz7XqRYFf4xQSEYwO01VbokWqzc7+VE
uOeOVMoFjECUETSgyR4C0tx1FWyWeThTFfNNYPddKwKS/24sEUoaKG76PJF+Ttwyn2xW9qrk2dw+
GqA9oG+ELTyff/ZFp052Tvyth8/OVb0T9pIlxAjIVEreNGTLC1Nm3GkWe2/OHgpEPtlaYobKnvK0
f8Ur1P0VxqxYK65mXyhhsDb2QISI78cMBoYxOYe+0/e9QUR/uX+pRHjSuuDXBumSfHrQy8jonXIQ
O/w0tzh3DLsNP/EUoLOa3v/B5+AhWD4DWbQ3y+ZkndgL8bEcdWJVVLFC8HAXYvneTJgyQTWTRpf7
yP/e2eZeG5MOhZBrCT6pVMuxtZC/P1yWriSSNV4H6ja/dXf0rMLScn+y+vho7NDU1KZV8Eu2OSnm
q8pYPUX8jvXcR9uWojMDAPWLorzEZQCt+CHgEuSxVC0qy3b2ynEJ7W8kgjvl8mWLm4rT5hu6Rv8X
FaesMpKG9Aoby5UYK8UbNQIC8m+Idy9w46R1Akiyd/nE/l/f+LrOQI0y51ByGcb7VnYNkAOsNS0H
oFdVsAVq32wyDgLm4VckmG8FWA==
`pragma protect end_protected

// 
