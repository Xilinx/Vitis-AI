`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59696)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT++8F4PPQq2cD1pLLMTjPTXpVh5mCVTmh7KwU2ZN0/MJ0FYpIDxT+DoqyjuaD8ThGgWkQP/
OT2OupVrEC0VpMdrnbNJm8/exNqphHU39mDmY6HG9gXbJ6AZ/ZnkaSJixLABYBGQdwnjNSsudfmz
TIPc5ypp0lPjwNkR/iup7djG40UgyIXT0qWDNJrS0GzEpIDFmnsAWWd2Gh0gPC6G0dEc0/ISJdkc
UBVlcIwhTL/aIGYzcu6u0hxmSfLjxzDrLvf9nDytBfh5dnPMUGS4D3OfezsRkbEJ70ArqbgptHiU
3nzjyaW13li0JXaS7wsWks4eWmlQoH/NwNnQQAiwPDQp8drrpbaRBK15UDTL9mEoQky9AwrruTCp
ciLEirNcyt2PN8r0GFg8oTIYazHx2WcuizTxqr4Np4qQs0fSUhVbKe/2dIQCs436d28rBTy2Hc70
1vv/sF6bk3+C+kZ4vl5qNaTAzEXGDGOCvgebwA8roWLd3MeTcFyghXNmVOk2YeZiV1Mha6xyDH9k
mdZTTV1D3rUYlrhrDtZLG8JZCpugt/XfYxC506V7viYEZflqUQyABVuV1eDATUR44nQt6GzrAKQZ
4vd4EmjkVDR2VNDwgu6VuzCT7YxIEEjU/VppsMnfeUcXVwqzIPGjUoebL3aRItFueuDzEF/yqEdW
nvuJdm8MUwFpBPvxTXIdPryuTKfCxoDD5E9lXAgwZ6bR5yel2/d0OdR/Qpjxi9NNwbM33khvUmWw
uv78eIT1p5clZq4EiDE+cT0KH/SjZqYAWevCHRc8QtvAjjlEtO5AaxI9atKSpPranIRgVjcIMtHQ
0EMkcdsVwwGMVIO8KibtKE6A8aMaQh/CLEUESNb2x9RFkEtWdAXtLPhlbo61K8H4snLJ1xJgaUcZ
02nELOcIMuO9SM5bT1Hd6LwgDCT6g7JPQlGwanKvT19fxrWZ2SCRRnzzwve0VUjk2TuWqTMDqY0N
g+kVyFxh8uz01jRSW+5Q+LT53nrKOtU/P1nppuTfFRtqMP+AKZ8FhM8lZ1HbdowpMjeSYQs7xB17
JywkGMDxulE5zuWCKc2Sv2AuTiNuQKdce+CYkXDKRvX6g0WyTEbfqjF+rBqiE9Lxprh4QLRQIrBJ
XxM3FXaUIHyzq7TqSldBGEvm9YmpDZlJbc7zdw7soiaygpxiExFXqukhZgSRmcrRVMn48FrWwucz
iV8tfs1tW+rknPTkGh1x6xCA1ipIM//r3FIj69/ommxU6r7ZTZ2Ji0pn9PDNh95kuudiLIV/4KZd
tVKjmfnh0IMmtVRYspTvVDZvwaj/4OrCvCtTDtwfkIIBIFq9l8LUqeD3XfvPfKq0EPaztwxVYN3m
7L4KCP58Vwqemarpy3ZEjqpwj4lEZLqDixhnAdlR/rJTYhBoKc/M6RgviiS56lW3kkxwOkhO9Web
gUQtS1oxl3asr1JZvZFhu/y06PvoWoNGIy+yAW54+zvf9mlFa/gmwz28kS7zBbxc1B/YYSVINGBT
iOSgZNCrxj9CLlKZHeqwl3g4uGXEpnhJ917kN/X47+hFv/5LbSeJLmApaH4yVdQiCuGeVpUxbFQM
qkx6btsxHIrqBm3nIl6yOIcAERojqVxklvZFF+QDgW0bD+Jii4gQO8Ired6F3GjrZ6DaaeDJAvIe
zXN0PJQTKOJiq2vcLvpz7aM70sgQTNQXd8MJdxSZZMgR1v5DCk4fIT6rHOZdpX5v94KaWzgrwf6E
ghRbPTTDDiB3s16J0SyCY2hsHAtFnfUi4py6UrIf2jQGmwx9krvpNlkFT1DtZxE51wmGTLS5q0N8
0o6vs16zeAWcbYVv+AUK1x1UvmQM/isHBVW17nDxFFGxSO/CyfYLIWQqsldkxQjoIVucPnXjNxtd
Azwcqkfh++8HlwDfNttLnQ3HbKs/Kj56jYU/NKLvN34KXXZRwnPvUPJQj5axKTwC+rN1Lv7h1T6w
CXf68JAvR5UcjS7mCHXHFvJvis4D7COr6zfeT5VKDbKzy3MHwbiymiAchSFT2Ry2mZnySIrQQ2WN
Xh4w7GYmkUWpFbVEbUzmP0ocNqOwcpHW9kJh+qoDp5GDzwk7rXQqQFTaPKSCc6v3QYMZFMbeIGe2
MOE0HkgrzNEzfb+/xMmFslndPMCMVz2LEZ6bntBme2SIl20o9+7I0EX2wgf89nx+KfM+Bp49hlgA
TmXV+0E/GogYb+cM1INrYI5bxABdcThRmZouS2jhv7jaW68YIRfwuRcgBJFZk3SXmkNrW5KBtq+i
Qv4XzPgbA91ucAbVn2czHl2z4Oi93yD9jN2Py4sQXbvOCtfd77VZ6QfX+SpINjo7ZFyBM6jw5JVF
joNW11Y+mbbKDRiW97BrraRFIKpLnO4Y/0PWogobM4scuw7xAh8O+kj0X1LugNDO2B5FEUY64CpX
S14BlOoyjDUOcE9lR3ReRdeKtXNHlym7J5TiTTeb+aDdpZxDnh14Hlx061ioQXrVu1i20wy62/an
9j7xvx6mgPoIlRTQC7FXebHtt2V0WGLOgb6qOeTMhu0Wb/FARDGSVnZms0nZso/sSqRMsm9UfV88
cKXT0iDTTU0CbzDjDmKG6hyI8Fwb0+qPMHxLkdwv2gwnhG7fYMLWPwcaV+FiRFQcjRcy5e2s6S1W
eevj8PQ1aHolLFqCJPgjm8a+JeZwcGWm7dMkvpWSaorp2v7qWh/X9P4dm1KXuz7ivg093/uIqPh8
oY7W8MqSzQbwgIcZDMfh2TPbUn3kATDWCSuYW2ZclzQVT2bknS44cTIn+sJBZUS+1riyDD/qBbu3
9+4KF8dvTZ2oUvhIpAArWjCeLdy+sq7q7IB+cyn4YiwXFd385pf0efexRtP9OLmmweJPwy3lIhlC
ebvD8BksnkPwpjxuFiri225Q3N5g9Y/M4QE2Ixx6qlH9j84aMU8Izt58XuJhFbbBQNP7DS2kguOt
LDkw0eQjl28sKqG8JdIrwIIFi24SH2D3+RoODzQHJPS5aKW1OC6D+MSAfjx4im2uRSbMH1EtBGLO
IFqwa1OKlDLbeTqSDw8WGW4VKmHybAuaihkVz3n3pjTMYxY6TPqCY/emmdaZOxna9pSCRPXRRMFm
e3uUudL8yix+trG3jmhsUpeqNAJbE7hApWSwtYzUa6/nGaTHyqjoCbe/LB08TWgSMEh526oEVRQ9
uMMa3w6r39ZL74FB9xe9xlgfPsj3/6IlTWS9W/1ez6yY+dSL1cVc5IJyOUUgo65ag2MKXhMf4RDU
puv/4Zfxax09vDX4DzKN/AUsMkRbULMJurpCERgVoNhPe7fI0yvUryLjfaP6A/EwT47xB6N7jNti
cdyytIjRJ6V06D70Zxkgkd93W1CJ6xGA4H0RHOiMzIwhlaY0A6CG3E1n8/fM2bepcG5jmn9ll9ht
3xOQVAzb/2cUNwvHC6Pp9Ecz1DV5Q/qIqflPT+G8Z973NMIOynt/4TgxZK/5L92pGSKkj20zjBYq
0unKI+m91mZcHszN8lv2GPD5v4turufkvgcH/MpPt2WoE1WBQBMxaoemHL+0zOTxj92fge31Hfmd
os9r9DJ4S8TN0pTniH30DoR14aGxRIkBM+6t02WEf4roFX2PY9i+Vf+i+kBRFMEh0xVXutj8uSS7
AOM60Mf+icxpt/rOf1e6xFJSMv7o2J6dfWq3ms1XW0eJ6R0ffdRmVTMu0aOse80E7MAE07hqmLlR
sOMB5Is0LA5VyqUwtD4btCVFiSV2e6e/nTYxNWiDxV3L6ryRRS6Vje/8sIxiBtKxjq1ZeSv5h7s/
85zmgutlE4TiV9plmEz6AeZLjTov3NMGObCF2uImPArQOg+j2zJMfNpDFUq7ChqZ+olqKIoVc8to
h/Y73qUbRBPSFCUsHf53+lPktGd4zo1JXk/GrtYZTDH+VhNNRZIWiSDIG6x2mED96Zs51Bdsdi/+
fy1ozIMoeOWmH8zQaWnvO280CdZgyOOQBeO1YnGTC/vrSwv9D4EdlrCN1QSSi5KMC4ha4YuX9RZb
IaPCN4+89W6lin6Oovr9rQgkeIA87EjRybAuuTcLcDYtQW15lWqXjAcTNdXw6hIMsmhyXzbUnKKB
KtZrO3ucKtuk56579RGwHXjXhgRPlaBWCE+zmM3rIUtv4673FpwxA3eo8IuLNJllKZEaztfeW3hL
TlkM1Rdj1QIfqWE4xv0RKWDfxeR+CwoEr0/5T0JDSb+DfrdWjgEXMT71ODk9yFYqRqaprTprbXrY
bgiKGg1/6kuxxIN6/f2ukpqQZZT4DTQrdsI51B2m+nU10F2GamwQe1Obj94Aksa+Du8B2sVrB6hB
WPff9HRt1ZxgOKx7yEDoSs1q4Yo0urYUTe8MysEC7Kb+LQ/vUYNFG0T9i0H1RNyt4Qg8OHe1UDYR
MwU5z8K8E6RYM7jRvqWq1VsFuCddyeIa1RuHCsX+zcucJgTwjPLjGRU0n4wAFU5V4DiXP0DaQz9u
NOSHxRbp73f5SFVwwo300A7J1tyO1i/+Yl8hr1CkhqqYSSFaM9lnNWkUDWpZkBkg7UIwfFGBRMtV
xvzXuC8gP1sBQ2yg3NGAVxIbIbc7nBnFZEMpSveeffj8Mm1G7UF2RrpP/NYhFrxuMM4n1Tyhwhl7
k/PDLj/pQb497ZL2gsg9kU2n+h3BtUp991Zu/5kWPcDRkKByj2eUTY14/LeyM04ZZ/5ETtPACEo2
O9bjVZtSIYDw6gQWXm4yDYDYpw6KaJoLoEDFmrMeEfSOY9PZ/1sNmapd+sD3AwHhGklyvBcA8swh
FEO4FTkzxW8to7X9YofsVJSZ716z+yvwDN60/7PerokofeQRnG/rqcxTnvwguIGgIvfAJz+x3X+b
3by13HASELkwsC8XfAR3Hy7yIaYRR9JrlJ52yy1vSFBPTZgpimhXpIKgJiIIOZf8S6I7GNuYFZS8
ZLcMfLDA3jSXJnhtGnRtXQzfktyI3BVErJkjyp0k0JUbGoxzTAug6ZEbKcaBLotHRkwViBseOvhz
Wgo1KwGlX9vImdNNCoDbhUcN2aj+84HLEXygLcLpJV778EKlpLTLcnhpBA45rFHRDB62M+2Nd4Q/
oi6+Px8YC4Q6cNJQNps3omZfE8Dz1sU3FbTo0ApMSoyFiC2cUPiUHSDKNJ5vzmPcRF2Gpw4RT2E2
siUagKuQKIH87OJdWzI/JCqMgx3dopbdLdWpUxLhtQaOjAs8c+Oe9yx6WD9jjUZYrhaQirIh2s62
IkdBO79mMe6MJvuVVs6rNnY/DVnjzoOOQXe5WqwMWVhUt3/WRZn2G/EH4xD38mNlK1AxNdRsJ6Xa
LvxfzodYJFmb9CBbb56ZH7XF6EO4M3boD1YNsuVVqhEkuaGYz1Bj63rg93a1H/fFFbY9QeIjtzX6
f4namYWxhiL8QlJoKMFqXC4ul7zn/3wuSMhLp/bBWrsmKoysm/CN3uOnpZTUmasKJCLza/nh8eNO
gnOvSr6dkeJ2DDt+TETPrLlFfiitMOEJXTrJ/dwYgUO7HnJ+QAezvA09wrKnBHXR28p/CzoOcbrx
NmQfat4CEpNpTG7IyVEwF17rUvNji7hUgmrwCw8rqMu4tbgDi5ozrvm95lAvwwodiAaiIHqJchYx
axmrE8UATYj78uD4E2PDklE/U0ZKEzUab3RAzCYUDIUAUfmoLb9NvTHhDhyKvjzGmQteomiLobEV
Dc8lXR5OsPCJnK9OmeV21bSKskePoxGOMxyQ8MqfXEHxK8ZHnhdTIfBocjQFCgT/JfikgG9OJ5gm
LBiWp0EEHOvmQbZa/0Oakew204q9+B4nzfOZpd/w/tQr/QmbUWT2+I6ubnIWMZ9FyBLd0xh37XI3
p7mVi8ZFBE+GL+23w9ON04aQ+nUMjP8+p10GqvjyIcsN/tX+vlrhFcmJH1osYD5Ynx/TZh8ehTUx
VK4Ga7dm/ZJsy91oHO5+Sfjt5AsLfrnEDf6rrjKszoVMoxaLx+H17ye3+P9Lan9DmMhQD6XWeOJX
vi1eW9x3jNjyLjXrvn6b3dDn+M1xvK+p1DaOLiXogyFSfVzLKmpJBiO/bumNpFKfKxz0PC6vCarl
nV4M5rBKiVyYwb1JZTfXqDQ2aQaytxBWoeaWznjNxvRjSgFnntjsgKOwz+inoheVkmcDeBpbqyf3
1n9lTQ4ydqpMN/1LBc4TENR+nPw/+pfSDkekOLCeRkgQiz95REozzfcbanBtJXEFOXeRfsyvc3w9
ul8dFuGpeAtYHR5LIcbYQNoxIEPcE7PiJIh6m68/yuTTqK5Hx3OguCKnxppbbNdKegO3nnmuYqA6
ZQWw4SI4zPK7/EgxipCrWMDo5UvFTzVs0nP6nu0zANF3lB3Z73P2M1A8PiW+nv6ecER5gJrvRbcI
3uDSeee5E6Yo/n0dR+5zFN9PvD0AErofjg+4vTeGRGO8Z8XpfbfWSgaLPLY2NA9+PaxtQGoFX6iJ
STwC2ez45eIyNJXFdbyZWVPKq3LJdc3icecCUS+naITzFAKAdLF6aGkcrCJBakzcvBeTv8DoubpN
esuoH+AslNbsvhEHezy2efyCCqixHR21YvYLIvPPpxQfTVnRF95HgC+bxl2I6Qu5ejUvOlANjvLx
3EXxXTeIHiqgt3mEU8JpZjPk5veBjsQg7bJiiKbDQRCIfviNuF7JEhCvIABvcgr9vCjZaB9sbtFP
SGjNCj3jt8eDYdlSpE7v5pRn5OMsAaZNmk91GY3KA110WxFtysHXHLHEve0j5Da4HzYKP9BPtW3g
wmqati+GaGZTBz4r46iNoDOFhBArvPPAlu5sk2CRrzddQFuY7ZIZHZ6pXhHsT+g1DnwLhMczOiVG
7BPLfxU0gINCkFY1GtGtyoMSBRG3q6jknjprnqiRdccTIMBWN4ItJE44gMPrvBE+vGxc/SjtdUTM
xpZs15AYHggApBRM3o0Mwri3i415Tcgwe7xckfuV5lxXyEdoT5AcACnj5yFXV2ZIH3XeoeCLBQ+I
QdV1SzPmOwEIlbVpXwsPYaqPMR9AMJKi1oiZZEufW4/B0mwPyVBQ1TupUDaHnPSk7bjs4+hkRnYQ
ZchS2VXEMoioll+EzXdj/rtEp21i7BJE0zNI3QJXpz1H6rLydkbDshOyK3VspfmMgFQlYe2mI5Ld
1DepI/gGQsJBci5bRXaEwZe9Vlc910BWLgSiXQwmnYQ0ZkfN0dzTP1AC+NPeFqCSld4PFYv9qEDf
zuk183Z6uGorQ2Ut2JW9Ho1161mRKhisVtBYnAOYqI2Obs3npJE+QxgY6NlqtGS/bSdJe8vNgyrT
mcyMA+mvTmagYIQW3azRkeeXDic+s218rOvK9iXaMa7tZ1k79n0Az05l02RXO1urdGVAzlqjc2Wn
HZYsoxe/Qqw4DO+8qhIdinNAE7O0v8wSMZi9LOGj5M1/HP/4pyGRZp6O5ce9UBVIVGkNdEFMp9LO
WFQf6vuJPNwHSCfr7rx8sKTGhl9/cUxznnSHduQBsIdB30UUDtIbsbvp5SaOuK3SfyuNTdYoCdL3
BanGlzV6P6N/dd8UKnQzBBh+p03jfeEcgZ5hUHFeXbLj+wkf3IQQl+62nfeVrmwMh7NkM06Wigmg
KFldQYSb37I6teS2RGYOB5eUsgUQNTZ7F2PIT2hwXCpFTqxzBZ6wZs4gDarSqIUnxRKLEONEfJUr
/eiD30YDi1wNz1NAjypdBOC7xLuNyO+Z9MxReAIxxKYP92++P/Kd3IrnqQvWMCe4j3jEocon2yrs
gFNVbMK1O60hY4kUPew7jP2zRYLBY5fGlbk8Z9Nce0VDU+FXaQuEiVbjXM0LWRvpVgW7W1RDePT6
yTV/RwovCKSRuNInNBlcUm8JGdgi9T5M2+yJvCHI1U2kFfqoY9gr6WC/49zPtBElYRxDIkkoVVdb
kWReSzABlvQkifFE6RskJh8bkhvByWGrnYfTJT6oczG42I74Ydel8F038ruxxle5jdvajqL7J9+U
3oXIkF0ow1c+QU81Wb6bgvy550Fja88gP6vogjeXun2Koy59qnHxZnVZLVtwTWya2f9TyO55x/pb
YIfI8FE2RyuO7lpNZ/jxU0QlblKLJEdjhpqEwqhd2ZUlFJgpqZatmGpGQm2JJIXF6QwuoaB3v8b0
VrYAXO3kfCmqXTk0NYkEK9p6tw5Fjrcx1mhQUKOd7RNsu7jBG7OYH8v0S7MMuGSrnQAeySRJq36O
M6LkwF8ujevAx3KM9CrmV9Hp9pcrIqANXRgsSohzcw8Xv9Wh7FoPmdOB4j9CNDbeF1rmGkJODYfJ
yqbAjVn0QDGiz1ZHOveibrN0MgqUrvVZGu02cGeatF+Fq6GQgtJ0BbEgKdXrY/Qq1e8hmfaeDL6i
QmIpj2fcZIHgL0CgE6UZojXslmJvXloDEwfpkhhgF65r8zcPeEZmMc0DQeC7RbPdXrMQVoQYsj1p
iGgq9j9RBGRfXOdnhyJyM2tpAuNuKuyJNymZuBTiHnBuI1ONxT24SutAbWhw1UhVFGFJ23uzZ6YW
Tyxv9Ui6CfoIMJohlTimQb6OBnZk8Ibg3baVCIvJHcEeMtoHlR1nWeZMByamL7F6W7+oXpSW0wIJ
IzY+qTOSzuv04WKA1dP8tIiVqzHaG9np0BW08NeqjRvDjnQG8tsMm/hi+MjGl9pEm3o8Yap4H7Q8
v9gRoM/6pRuNLU30rp6brVqB1amvhvtsG+Lxo1DWKGF9pGA1rOWrVCZh816P9/c0QgVLx3InEdgs
Ne2OE/FfxUZnGviprIja0d5mpD6ZV0cgB8+Lmxo6fDPz3sNepghjSPFyCepdIeX95VV5qeWRa7wR
1p7W/y4+i3BYkDkFkiGxSR90nZblH7VnEOzoiJbT9g+OEhu+7ovpByZNkbOrMR39NfyPSCZvT+v9
VJs5zaPlvePm4tgrUOT/7gcXoUutgRpAaiuTr2tWBfsS7eJfKDQpupC128L7GgB0r7kIg5nrWFQG
ZxZxdDJolNut+k4mm3002vp6mBES6b48iv3aUXdKVIYMzTeII7NulOqOAqkOhNs86hiCwHVJzxu3
O/9MQxvm/oDsXrf8qY2uPre9naJJ3p7Zq06k6GavZtp3fNUZj2VhAqJOYmcxVEaNKEjYbTsCxNBE
LWSj4CvhNNqiolJQlpz/DDqDUpC567GOJfGYWl8yFDE4GZqreBfsRgd4UzEDU3XviFfnPFUwedjZ
OpUTtdfkK8L1rf60xe4Ah4nFo/+hmGTeGBcAa7yGooHSN/Rr2PR9loD2pANfP/aWbQl6rwO4iWgW
UyVilBoI4khVFv/hcyoFhqtlZn88zj5xJLrXNJYAdRz2K376WKRLv/ufTOnu9hM8pRyXyogTxoB8
v7FAcnyGMjsl5bEqvRD37A4OKCGy62MYPqbblKou0Le+smwhkOmiKKo/zYgCKSP8FcZ86Y5I1hlS
AUCph4ETkzq3A+CinvW5UFJhDOU/7lFgA1OOLrcLXwy68FdrAQEuiyXzIBPsud3QcOnObLmN+OLJ
lozGGZXKAMvNDPLluY8RH0nwtBr9YnbagonKipR+84KRPQlDbuku8yZ8Hh6fkOH1TnPPXKVQjGTj
yUcSmGCpK0UfF7geD4/iQkULCKDV8wtv1ImarDNBVbeALFTzI3eG+S7QUwZm+iXjMi4kHf1sJ/5e
xh3dmsRVKBXpk+PhEw3AsMJUcIktb9orkC4vYI3VdQAm2vhqTRb7Pp+dmHWG8jvxVZeUgOAw9Ugu
VwOceQeyaLupiSPkcNf6A+fF/OZX/ifHaXucfRpFWAM3InFzygThBPGGdp0MMKlW85d0KHzKCyeN
9xA821aXMc5+77fB6XW1JFabBfLyZWh9yxFhXkebV2PKJ3kGqicVu2jMzs/SIo6kAEFylh8MElgz
BcGiJLKcp8N3LHukEdOmmXTDZc+pZp5nrvTh+0+d3gi4ZlITu0RqOiR4+gRSzj6gkZ8FHwSfq08m
pvloDvqp77DA85eNYyD0OdesIq0QuZNop2KXtynaEmyZwXzlbpqq0TkKRXkMwK9p9ToSorwe2TLJ
l0sQsek3kjF++YgWM8jJRUUa2RPXfQ4l/1+Dpi1Y92X8Rl4haowgExHfhXkvZ89bj1fl0Utsu8IP
AwiLWrfayHRVccX72HVF8syVP8NCUnIVlR6xWMKT9Mj5X7csygxIUzOrFeUktvjprXOHiUZxjxsw
z7STyHbV2mRagraoSWl+FL9tQ8He3PwmPpf0z2hcNLRtdPs+XavdoyAcpsBjIMz3PG5T/ULW37hw
y2h2flazM/c1gUdNRGzf9sURWInpMsioO7NXKm8uTnBZ+QHWR/a4pYPaZwhmE3nIOSOa8JK52CtO
3fVGNbgM1HkfoeRFGjdib/aT9vjG+8/lUPF5BfX1U14SPXQhe8hem4eXYpAzbQrs0fYhnGDycqoN
z6qaRnz7UDv5258SlPfayaOBnimkqwgGxr7VOFKHyiX8LgE37G0plM7mZ8OABmEGoOaJIORIwXVd
AU1YKGP1vu1byMXdT6VaukOuJuDIfMPMp9/EubATLQk4R7WHu7UpIVewDfHlnD6HEMGbgGmpTXZN
9xZOKlHAoim8H7qz/SWVMvBMVJqgOZL8k3RWDJ4vXm6POxHo0JIbBxmNF2H8BDVN/efUX/7yN6DX
TrXWvO0EqNE8YoXMED3Y4NEvzLa95QpQgiERf6AXuVQPUjvIQM0CrYYhPN5vd3SZj/H37nTwqS1Y
UV9EpMpa2oEK9e6PNA7R5paTtAKM9JqKfSweZrDV7wKNVutOj+TpxVKDMwKPH5xFn748Xjz7dPaP
vrLJL1KtARSA0xraWDKJN2zxSXyiE+xkKv/PHAN7UG2kmQx3Vt1ki4RmQiAK23OnRG6X89wwvaQD
R6iyuXdU6BqNVBMWCqNq9IkngRUhCyqlKf9Y45vISZDHvxKVXxtbigGUyV9JyDi9/hta9HVMQZEm
+4p5yGeTRQ26gDETioKdjVeX0cAEMjGm5e8xYvQAKq+WoioZN2Qzw1EnIA/UPbgP+kkY9dpai98v
FFKL+BZq2FytfF8EvCX+sZtZbill/1jBfOoiso/DmYhhg2VVUwAs8ZE6DmaR80Vxhk5GJk20SiQ0
VTKO5+bM7JzvvrwagIi7fH4Z61OQtTyvBlXlOSRzE6wFrO0yiZD98JDXFONh+MtszewtsvBrDHJ6
+Xly+J4ribBnBhsoiERXDDdgnDuSPGFKsnSlQipvQiuv9CvKqDZC1ubdUTALPuhdEqfHVAYe/lG3
zwHtE9TN5avOh52yHZPdsxBS/GJEMql/afDvSf+Zr3yMhmExA5F12eX/nFSn9i73DCalmEkYsxAe
Fe/L+cIvDg6lxha/pRtx1hYEbd/DEsePAZcM2jy8S5sKDp3hnLcCNicm2IELSJ433WA/dYc2EMQ5
bAZQjXPN1LbAOFFvHy123xs3aWwdS2ACjpyAaJ7SodXIcDBR1c+wx9sUD7ViyTuOLu/dTgM4XLma
eC33XB5KOAaSNcT5ub5ajo+0L45QaD+d64ZGnogcmXHUnQX7KtmQ5BRVJtuKfC55R17X/EAvpOrj
uEPlQwOqe2LF01PpHwHRa4nZfJxa44eK+njkbJkMJHSNX+Q2PX7DrVwwfXalirhxjieL+/aJSWVE
RHcMzdux28oPvP8/+IPr8ClSuNRnRLIn4ou2YnH4ux1REwqRjgHaQ5AuvobIB1+0yRyAvV+ZuL8V
S8lkX7O40lM3c+jmK2cAYX2+0bUelEMJv8ZAPEftbUIIlo6/YeR+VK2JuAATu+F9MDduCxf+Hf5W
pPV2UBxBWnbWWxUB3i9nm1MbOaOBgmuoRaEo/APcvywSsvxSoun4aBX2Fx5gxvbvgnmulF5TtuiJ
Id/IaMf5efXjBfJBSQgKrMIXFVZ0MPSDEJsK0jozjxx35TlNRn/6Z+G4m27xSGd5pQMv6Tn6b/Am
6H2B3z0biNzixADYQZFgPq4EAmwYBTQ6lQcAADhbstPOqJxV3dZFDjhyZ737r6ZCg41L8uWLvefT
E1pe74G3a92Af8SIcBp9US37CNlDyvYmnYs1wav4XM/m6IBKMIjuS3cuH9FBgQO2szzl3AOjtGni
TP4ymB2ayMG+atQwuPrOUSjwA587nnd3vhdf9KrukJmYPaDZDaogXJ0lG+1yUHh8Q6Yi6qLChoL7
325nYcqp/kt6Ncz9/Mgm7zgkxJ8A2CIY14uNRAma1QOw5f5BdDaQODynRF1YGFFXOe8x4ZyaMmWl
GccvNjD2YCHFNXBoC6Do/dz+sV6UoRH99XlKNLPIrhcti4aGR9WOj+Saghl6dE2ftvdQ/Wu22b1a
EI6ZpK4QaS/4hIySa+R4JGsnrYadOb60s/8DCBnGoAfghwOKoydyrnLclveAiNr4BwaIDAXLhrJP
i/IZczWMiwPbaPBHKL6pdKSW0EScDHk3m2QTUJsuB7LIdENRWrgc4k0qmXFvxXQ08QNxFpeOVyOl
2CLxOgURfc+ku6a6/n9t2lSXs9fUPCQTcJtA06+uOqqW2ZH5mx9eNWhxiBp7jjznHkUSA4tc+IAa
p1vZwbXzJQ+wgobNUCShZZZrinbSUxTIXglL1aLKAKMgxI2d2ebnl5SwalhbeieNlOXf235eZbyY
3wggyjP0cuiPpk2WhRMRd104HvrT8xcqLgmMXTUIrMJoi7pFcAmLLEDRymcAS3Tq6aoq/agvvCzw
zMca/2e4t0Y2tRB/eQrkjd8phjmCd4eIX2FMJrG6G7KMCo5FbQTaQR5CjmKkZAz/BZGn0GI2LjgO
7WRtCJvM0qEmUyJ5tc3JlieJeAerWbdTS5Vrb1crxL5Nv8QNjnCQYu8Cc7/+SeuCt8hgQlnZRYrZ
RYXWO0B02dA40bTB4S6uJb9qLmzFa2bfj1uOzI8RUqJ2YRr4K60XoJEyTOYXJMt7VgTIkJDLr0fI
XfzFSeSHHR4UtbagnpwDjzVyAV3RHt2C8FL74mIC8Y+O50Rt77irB6x2dvhdcnB3IBraebRyssDL
be8d2ZunGilSUKKyDAj4qK71LnVr9in/AGkCYJdKCsSEKbD2edyNMbpCH7WW16tmLfYS1y7NZqst
a82T1l3zolox9aAAfUtk9wkPAM9uR0oDT2JYiEGAura+1fH5PZOzEklTv1P25oT+kMS+3Yap+ncR
a3AoRpWSqwMCPsf+kp4HoiOyzdkMRsHLGVWz1cB7vmFXeVZNLI750ql4zDXgQ5DeQI+fkgWsPqYw
PX5qqXgeiEE5SVnJTwWGUG/NQTW81zhMrPV3+tOYC+KkMUjdWDFMB7n8zlA/tqJws6wqn31358Kk
tvribpCON0KcPcPBc4iL7ugsTlvTQH6z8wSsXY8j0FgIncC8b/pP0515uJphPRIM6L+qCGHmAnaB
WQQ+4rggQ5DUROks1tQUDwszpE7vhQMpqMj4pGBw4If8pyVot2HjZ19i8RBGTc4JEyNje/8VqZST
yDwVL/PUkPPN4Ol6cOzBdReV1d2rrK//HbQ8blmq0raiyoFiERYfTGr/ksCecJiGaQAxIkhdxuwq
TAJVtZ7RjH63r6K9/6ZvxYmq/eAZQjuztTrKPUfgesQIGaBHnqNPWJJkPaD/u77LhU2+PypcqOG5
H93Kd3lWwhFWStC/R6//yabmXSKsGj0JjFBp9bEVtpCDfUE9RsiaY24eD/PXaa82yIZMSOval6+C
1uEjwRDKZ7fyyVgH7GBy0sv8w7od9pN2LruKaZ6RpRKJcGnuxJiCYOwyLi+D/512Uy2BQZyvr6EO
Torri3f1+VDe70WT4bgTyMPZvZCZJRLuJQVtQzOeoQQoqnBLoonZJnKltyHw8nvVQNx9ASDKawYz
zWE/vKUK0AsLoQlcuXGO+z65gOfwfRMq7jmyRtK7Y6Arx7ccp7TbnJFu/Q/tPZ3Pj7gh/d2sweTV
annTACkOvsDcPKRy4oRhy/s0lutbbLEwjd8JHEDs791jtdpF1PaVie8R+6E1sRejHhjluWv0diBc
alrDqcjQ+0ir6vBkAhtsTsUtcyokklDmZKnj23dnuq/QaxK20IgLfpW/mAiNwganZr/CURd5c6Z2
fzxOsI98eyBJVBW1URkN/xsJmVOe2N3LUiPJJU11SSE5/tuTzaDPHuV7ARu3RXL4g21XyRZTimsK
dsyDCSFFgueXQ8If38M12a/vePrTocs5Sg9W0ZYxY3/hZ6aTPZxX0iPI2Fb7S4VthWLHiwI7wDnL
6AMYs+vNsmjHSmaTbOpP9AsOMotn/0v/GGgbrEckX8iKIyFpUBAuaJFk4To6yWH5FttHM+eUH07z
Mj/+UbrEOIcRscrlcY5NaMM+fnblvJsYSp2TBucAT91pLuTk8jBd/7swBC6LSqlV1DhpKCf+Srd7
BmN1Z/tWmxAJTY1llvjOnWNofayKRwHH12nBYtLolM9mHqa3dT2EISJouSCro42rp+WYWc6WOe3j
LtNQ6tXJ2LEEAdj+WCNHMQVFy74ybuX2KL5GP6n4KzkHsUHV5qmiKnZJ/DUevMEitZzLBa7y6rCq
2VH/mPO5Eayecd4eH2eQVd3SoqnLxDgZjmfohCUKcPbNYRzoPRoF+LxaWlpuzZXIOkwSg2FtgKcM
5F2jTw8kkVslWr0JvYmljm0ZeYFEJWf3ffGDVuyd82TsSWegrg+9HL4qIMvHR+HtdmFwOAz+GR2r
3B9eamYJPq4k2IoakJ7aFFVWGlq4neN+himRaY2IckP01AddqDf/tfC9R6EnBlQBTxEqXYjpjKYo
RZ4BsfPUixl0BmUcHx9DpgfcvQLAkAlAUa47Ob/gsuRZ6YxzxrXRkr34QZUT3MzuSxywKRGuBLnV
vJiiI7pyyTR3wLKSGWmjAZbA7i0M0pYNlZqGB8Xa9nhoOeTG/Ot7KZ+Cepf5HxKLpXHOFg1QdUH4
2hBXz5aJ4fBzGZ4DXgS8S/8JX/gHNYshdoYRI6V10Ih1ja+q1Y69i3f42TC69OME2Em7svFatZdW
M7NjgXJTM8jWCE4f1ROyPapNCLC/e0KeF1/AxlUSk1qJueXaQIYOa+IBTQRfV4vNTbdUno2p9Dwq
uwRJg8qENmanjuwF/dyFLrQa7L87lAiJjD5aJoBQslhO0nA9Y8hKnOWzoZhpBU3YRobY/VB90Wb/
HcXHRX1C/6lo0yIvLvCfLuhFQS9ur4aZyd1Mnnp+NeajJFBTwDI7imbBxJkT86rrjyWh4Bvr73/g
Uq7SaNeIlsfYMmlW4EAwXjESoxh5P9uCFa9RDm41rTBaEm3Xr4SZc2kMLP3+vj03rUEqOl+di7ZW
c3YCdEHTXwaFw57U1ni6R6fHOz2mGbULY+zgPc8Lx0JrXA8EczQhvXu+9W0HUkEcte8XVL0lIc24
ww4Dsen3XcWtnYXnsDFJ9b6wGVGYIe5A4InyljeQY3DTLAkq4BYUxuktJYoOgVErCfnJBqW9T1It
dHqIAO++fVD7xPwE0AqFIwqm/lQYbuBZ2iWLEKPGipe5FW+NhiQStsIn9BspLhJLUUrXnbnkCKf4
s4440es3f0ZMSYAIs4BlYduRsxtHEfBSAvzHmRoxL0BdCxvFzRytCIo2dkfcn5sbTNJrnJgR4s3U
xLVXFlwY+vi9uedzlwLaZ8hpE2deGT+pOtEqr6CgBm4z1XCd5W+nQG02IB5Ge0pdQqBm6L02btN2
9AiezISBZMw9/yqJTpQqbV3uG3FjqoVW+ejFT5f+wmbByFMGLWOG8MnqGMj31H4JetSuithfj6dD
v8Y7vGV9A5b438l3V1lPTOAGvMaeq6FB7XuOfeCyZsqhX7Dr4+V+IorQXNATcWF79bvCAuVxt5a9
Kq15ZJ087I1vXUqHs7GlAIVJ8YRj5z5hGdj8cgkaUyn46mFPCK0Zw6Mxl4eu7FzfzZHrdKtuvBXO
53w7uO2UlvMaXEBAZj4OUGmLETQ2xuo/SQaESg7QRYMnEMMPQb9NRPoHT7adDdeKBvWmzIPScKbE
8HL+FsYc2Svu/f6uKrmOR5gzmKRTX5/IVIolgH2sskPYaefK4xsR5vhnVAV4b+wbSTOc8m9RfW28
agvoKM5s5xAimAxsRAwapQM47HmgBECHK9pvLLe1+mz+X8AS+gHpXsMlMEIzpKhc7aAPK5O5efTP
Un//qhhRMAyUAcp8ijzYXTB4gezJXHllgFjHaVjBzwf1hDEBUoRWAJ89cjTvXtuL4A3BCvb4Xbg/
EzOzfV75XZixoYwU2A5ZDCETKk+MCjmojXNZ5f0HqtyDMi8btzL861VvFqYBvw8AMu8KJLYzLjUP
HIkPStjZOT0op1gK/FOY7CidBooobIEmYAwLO1+LejdRmQBrQZoRCXabmyUitGjk9wCMFvmlEigM
euvjkH2p3ZfN2WKY6QsMWNsB3Z0VFaGnSCvn7XJm29076ppf6feLVmkK3EKc2ZBl8z7IUPUWwjzb
Lsb36OaStXS0R7doxjV7kwDL+83RxjRRa0SvBRoRsKoT5msA99YMEnzYB+h+NDaKKi9S+fJJyXye
v1C787igJPGaJHyxPKujh3E/kUvZ33R78zm50iKIW8fGUBKZ4s8yQDNRlOtnv4cCxSDAqRVV80+0
jzBwRgMQdk9boNM6t7q6HTl7YN54m5i5UBWaieuffQh78/JsL3lJCOsNM3XiomeirVcs1yRX1KGX
PDc5fJCWKmcDcCeczzqgQ6rb6P2eug+WnGeGc0pn8E/Zm4VkSAoFwTyUdmW+VjKpw6OprrMiPZ6K
LDgnS9IYZsKi+99Oi2QAtOhlsg0p+a2jhnpItv3j8YDJjf39iqBfwJzR32VrZxLjsLnfS9EOLXWs
ChSbOjgC7uSUyiA8sznhSTXsYeKyKFyg6N7kPK/OSq5843QhaxpiLqK26ppByOv0cmJYKqVSY8L5
mMrWISu4HqY6qFmzZPmEVPuYeljpHCgZvdpwsMFyu8oKu+2p2DAFMymQE1EHA3RfQNZufMZFsE+V
0gcoNN7KJ90R7SV0s+roUbSvP2GjY+B1qfTbAN5rUjDFAhuzkGuw439Bdnjgg31viIa+lNKclh10
Q6SmOb8/90jDfTOZImV2OA333LdOJ+LFQUdAr2ZtJubBg+xcrSL9RB6T1sgGpzby0Krts7Gghvl0
5B2gBvTl3Z/85uhbwAlV920D9DsEIjp7NOE2m/Bs/Syb1J4PADRp/qngV5EmIlgDH3R/0rmAp4Pz
FKPqXQeBg4t3OegsOPwllEVeOYs2dqhIh4AjCArakvxR//kvQUMs1ZMH6H95eY+qbZRFte+IJr/u
QGnLTTHYgTxIjIYTtogaEKr6ZmjJ5Th9kaX2bvSGC6ekR+tjpP+bvW/LTj33VejcCilrDHoHVZBl
MmcyZe9FqBKadF6MKJnw0JmdDBEBhYe1xH+GBxydAG2cf5BLkgksZCoXPikxSJUBQUKruPzq1YKI
UHAMEbdbeWb+J6uHnNhHyR53PLgGwWvVorNcILo4yndKFFIp+ipIr4mdBDOrrMnscyTNPmhpJP8o
Z9956RX9pXnj0IjxcQFFrzosaTkX5NqytAiAWawzXfHM2gJV2okK4sP5JTxbTuIOzhNzMQHx5Db7
iTH/aKASRB0Iee/DhPMf1OcH/+kP5qYgoSSw6Ph1S73+dWZozDVHnoGxijWqQ5u40v5gnBjU17Gp
IC5BiIV0Qi12rcEpa+nORWQXFESlWTQdxkKQasZIRslUpL+bE50ocUsv4QSNBnm4QPZ3cwZ0aftB
fSpqETOBgzk6O/Fh6k2YM4wSjJ/6hVKpag6FR2OazTRrm8uXkbtB1Uy4Pgg5coYHG9vBPL/RFjkP
htGBPxmUUk38u5MT4sJBCHDORVLuGyXUiB2lP8Q3iUlarp5OJ3BAOTseKHAu4FSI4aJbboUH+zKB
Iy85WRdew7JRx74Wofl4q7DQIMwNkePxznLx6FE+v4aFyD22kAVumR0gTlnWhQ6ApeSbFKo3z7py
wfOY3YX8aWNNs9XzRgSFPAlQQ/b7EHalTsdFJ9Yki85vQjVuXBgC17h6tnUy9VldB3F6T3nI4FWW
ZMMQny/FJkwrgZiU9CVGWpiYjEyz3QNr1+S1UeJnFsl2uKRUh5TSxdPyXqSzfC+CRmvcNZgokJMZ
72OWt6OUK7bLKABfc9ZyO1dzY2eEuI2atE62WsU39rbgLwW62WhJ2Oeq6Jq/shn+GT7G9Qj4JXfm
QPTux6mdgGIsyee6NegYe6VkmH3c2dE1zlthXhrZHxtUt/E1Sii2/CXu7P88fQnkhufiHRYav1ud
dDa5BqxZ+NWyxBuuCJ2Rbd9lx8RQVMCp3INBKt2PC69/9ekPJ4xAYJNM4fjvcUeT26fjpHptDB+b
KgBd5DSPmM/okefzuWrNv/gXsycTWb4vviXs+ioUfsUTOwG8TE/76L74Ob5ZpKE71TYVTvfew7OL
SafQTYSm2vWBCeXNLgNI/82g53KRu4eaZ9tlxb3t9qFnX3dzo2cTsUi1V2qmRB+TQ7C/FWwZudQI
1+7lmc3mf4KQK1aKvH9VjqpxU+yvGi2aop9PvJqoMK9IWuupEFEIApoxOQgbeodZxgBPWfMfnQ3s
0bxy+wK3Y3BnN8pLO5ISYXZ+zh3B16DoXSlvUFF+SR66EeUVZFVHAYicCys5LId78xye5neTFHMV
FAczKjWO4kzW+tOc8vwh4FuGL7gpIAJhIjn5kvdMSxdbWhA7FQyb5xj0sXSqYuweVrg1AaMBiq/X
Xoz4jrn+h2wecgyx/jrPdFNi514CAL6Se57g3+a06k/UtlRljzel1amp3KCOsMopmA9z0JmpS/bF
t5o1EmQD4Oocsx3//l1eE73nWXHeDAFkYvcMYAeuG4tQcqJN3tM1V/3BTcjJtm9/NwKGsJuFja+l
IPMuOzfjUjQrYobaww1jZ4sO2og9Y8Lo5wGMSLSWJ+gsELQn9MChRGMm7w8YL59mb/TaOSHVV4xg
5tmwMeSnqlfFDaiMeoGVv9M+ZV1t9SrrTclzaUpHP6CY7/mkI+zxHEQF+Yx5cFmrghx2BovXvCzi
7Q1//+K7nFNK8iOW8OO1Ua+DblBEVlmdB/tSPDOIhGQj4+L18faLIEK8eC+OnWOYA3DVk/wXvmM1
9iQyPyUQJoNhsnlpyEl86rtvDmRg+dZCEV1CUwOw3f1nxJVHwvk35oAw9lVcs0Z5wWX6r+SWycn3
Wjy8JAh0QfOgPWnTOFMWVxa8f2bVUL0NViJPRi63pT8IH8td7qfR0BmHZtEGtEBePhL9JtSQpnZX
2yYnx0cuhMs24MfvYjRI17/4PKl1WBtx8uBYhoL0eezLtmBkhnHlrfA6p7UY5eKHVsxdzStyc2rr
eVnG6NaFVSkzmTphvSAjo3xK71mYKg9LYfo0a9h4ZgJDTaWdKSYgDS8LxNJmZlW2ODwMCC2SkLMf
7/talCe9D5tWChcP3LEbRVZnFYegp7rPB5xqvipejzswSgw2yM6+rbj215RVeXYKtx751Np7cY6s
lPT9u6NxsZlALlLjsZZc5/yOZzP3TT9wTDk4t/AHjJsGsP1NXHm7cpHAgEJm7eskPC+LbxlIQJOx
Q0YjfihY/lcNoRw0LObbsbl9Nm6vSp4eV38eU2aoLCFZgUMKCL9ktR++Qemv6iEZiYAfkobGy/2g
2FjnHXtd/QGq69nrvOhznzsQAgimB3o6HPGS+jFCUbD2iIUn/GVf/fdMuo3g79oXv7K31RjCDE8f
M40cuoLnYp30U8gHeZ1OIv0tDL6BtQTLkrS53Kz4/7TksrJtSbU+WjkBCmAbv+89KvxwePUUP8MB
B4Ry84jKs1m6RDvoCuGk0nayR38+7fMOA/38amWFHZ3C0oPd+c293cmSFfF1N7YNCy47pb1dIM99
xXDCFoqO/8FICvwE0yvEedr7WHOFwvgPuLPSw1o2c2kBa4MNZiJTDYcEokU7VPZ5l86q4YNJLPeg
pral7XGTmx3dTJI9L0qS1mZZkqwrSaZt7dNdLHVx1zzrFhmlbNMT46eLuzziUSMN5dcNbrW8GKOQ
nIGnImLrDVPTLCCnAP62vtqU8vNSt9lRwjR1mxd1NhGbjloI07nURPjOjh8RHcexhmdEptaqa2Po
lrBf6dk30/TrlBgV0sS1a3cbZrGNWD5dnF++V+9paGdgA3HACmwy8ZFRDc9M5z+JCOa+A5T71GCY
g45yQM6LLTzgC4s26WDFcN6rcav2rje5geEk0UVoVxiTega9Al+xZgFMMb4HZuHrUiSk0IYXSN4f
qbkAJh0J1gTEHF2IzJKDZ/YLAT/JFdHBNZZsjTNU755REY6eeq/9/prf8eBBj/rpzqxOpL3RrlC+
7oflqOLQdvQ5HLbNNdFDxb5CuVC0gjMPO6GuhWGCXCacfMAVOfvWPnWQZS9VPmI3CvFRbWiXX0q1
q8I6QeWOxyZMmbfcrH339l42n7OiE30wNslziiEiD2Q5OZ9GqRZw/f+btj7SwrDvfz7xhdTgvbC0
kCVuI3/91GyQ6NvH9BgawPTr3qcRqPnvnpn0hJp5bUiijeNCocGQE1HNHQcusxk0gZb3Z1UiteEy
4c/m3/IJQli7Fh+SwhGDikvQUiYGmhZRNCD0CxWkdMky/bunIMHQ/FELWDUbdNZzoDG6Y8hpxr5i
FrZzHL4grm3k7QPjDJcUXxLUOhZDBobaET52NFTiMeAQnFDzZURuLq/Tu/fiAgTNOKuFsarU/YCb
Kxk5dkCoowPJJXq2xNIBMyUA+uYwt8DobNknk/qx/J7oyCctp/ytyoiWZFAhO/2bS/9nfiBBgIxi
mj6Y+y2ZCx7/M5Za9/0NOeqawIGIwBaxdpGswF/QsTtXuaKbX7N4MZXCG6FWZx3LePvgDlC7wKn8
CnnWvlVykoqGXyawxZxIRILKP6dUPHcg+kU3pEDAfuu9ipWonRopkARM5lMC74rPDm/rvONSGpMh
ULh/yOeU2jXRsPYp9meENvM1c2YEafQqZI9PgztbhmsiKG6y8vqxx0/WGlG3B0k3fEVr/LNY7PtW
5x0DnkO55HqOm49rLUDQxOInQr5CjzUwVzRA/Ln1Zbl2nj3oeqhMBYazZiOg0Bwu56ED/qDjtE1T
rXvpDRjx+6m5DBFhhDOFaaHWDUFmG1uM0B02j8dhFe3aJjMvP9kMl+bosGUneHXHJc29a2tHwth0
DjrTpgttjtLCIxg13/R+bglzDGcpefgvXP0ypCj93e474wJGsGjLHVmrmBcfNr/nJEmdNoHgvcjg
x4T78nujuVJl8dM25RjF4QTqfI9xrrmlQlzKdNuzduXoN/PtrcI2Xos1VJix/n11F8F8iiy/BIRT
PKv0xfQ2FuMfm55mT2CAhRz+tIAXTqZvc0plEfyzoRMXBcqx9ZEC03voh9Ywu+OsUMlTjak7t/oC
oCtAV+kxHDdWt1SKBS3kQA5z9Tr91rLIczFgdAOAD66YQMnpwG+QZbv/H7AMJIhGHsZ0KmC5r3f0
EbEyV9yCnylYCFeYM3uNXeeTVmqgYbH1f3NGhmj9HSSmNgDyvLXmlxJjC5oGpq71h9p9jigp6yM9
a5d33XbBRvig0dQJDRkwXIOam5ENEZ/TVEuSFyxlp5qvzFX2k7mXln6hgjcqKsdgjQpNLnjHGMui
pMYpeZj6YPJjaWuqwI9dGdvTm9ZyzpwB6AsJXpYdMwr9GulvZA4I8aMpxe8wf8PrceDnIYXsjFEI
kr5wA/IfN1dWn0qaDoPjcUzixUQXVHbCZoGpwdEBrnpkQs1VGbR87rIsxU0dEDEfNPvn3/hdf5C2
IwLTP63R/xp/Fqwz8LKP8C8+4c/54lpL0nGfyT5Sa/BRUxslu8pKBRIQY9Iry5DXCAIkEuon9bwm
RW1wawrMgdUGaYOct8iPZxnM7vUedUKQV2NneuaQMjzFrLTdND4Yry25kS/1APOewAUa7AvhiITD
YfCuZJHphzboaZRyZwev51wz0Jc3h7GCHSv5vF0xy5XE7Rfoc3gffq01mpOiMP07QCTjQvr6N0Gx
vVC73sGS1xrVZC34TDCvtVj968eJl4gPZ9FAY0tGlpTs/lZ406cEJBtFHLy+gn8afkllhnyzoeh2
KRnd2ivqdDjwxhf/xyRhJa6jTbOvoK7+kxmEdXGkoaUf/0h0Q2Nzt9CnXolw78jjZBlPOr6qAe6D
SMEdg3IaKTT2h6PZAW74/YNVdYjFaE0Hb5u8S77wRDXxWAR7Dd0F/MaR8Dp2Gc2J7QcOcpVG/uva
+oppDIbLuW12eTI+egdgc2GU5yZHZpHnGzTIULzQoP9odpU2kLpCOPCIHthFKcLBSTZvXDqS/4YM
2xUosubqB77pJDlTfmiODxBXbZLR1wIIF9ktFcN/GQEGKgITlysHmdfril7VGL7cgMS0KMtu5HAL
bc8pfZBzfwD3qIyfZPRT09i1DagK1kve35SKUymMEsGfUknZF3wJKe33o0wn+36TJ87GDUxAHDnM
fvqa58LxF0QDQM8lIH9RHMdRHL6+ZFXeYZBXrRAg+2eKrHDRP6Id3GeamIdv9QGZzfVs7w77MZZs
sUeACSxa9Fhh75DalgdzcpQtCaH/kXGJAhqU4UrQxsDWDGtWkeL+CFkRiLehWOqBKxeqM2LuNs5c
uKFhOzJ64Rw2kXUR717vdl0nKLAS0eCkfsbHhHm5Hacuu4G92oT99cii9EAIX4pbBXXQR+e7Kj9W
kMm0ve4VU+pHfptmaYbvTHFWGobJWZJLd5vJyOjtcYGy66QwJzynRYnW6RLjtFvKSApfL56fSk+I
zQDvRnShtQXDtd1V+nQ8dzVsnabTR3+rgrDjgzR4QdF0+eBAdNcguVo4zFEFjmszYpUW+SCPbKPC
Mz0AWhVg5So2vJqzA/T6GYJcvf+ZZr2+oteV8qH7OsuMZEX4tSX2mKLKRrQbHKYAuNqAXQTbscjq
PhyfjFy8zN14jpCnD+2X2cpBmtpvIwwKYNpo8yOcx6KbWOrLkDRdjMCS0fYIzA9xB69XO2sIw8Nd
j76ETbX6giF/9txMsiYYaqWRcCyXOMaDgBxkvmVufeUAiKwHW9+2DtZuLjQWrHMLbGSUoV3zveqf
GOg9xkVAjl1iUkN/RBP6YZqqZZHilv8SG+WSE7LMmQcCQQw1MhLa/YMvDm4/hSQ5P7F7/HuIZNIe
PPZhy2w8E0E9sop8aYzQVbnsk8Hha3EaPJYfu6iUwGKfq4fO4A6X6Pt0YXxEQH3wFnVWsDLK3+9C
ZC82z1a57TGdCwlnVPdgPYpCDJVlkf6hoSeiuUneigb2ur4RdMWb6FTsEv//XSiAVv+4Kxd7dlr0
KKM+fnIdWXEsY1AHTocY4OYMHDGoP1VwxbLCv2UEq9WDCiK+qn39Y0AieqRpzsZgS1j/En+P6EGg
3Eg1lh+ybLYk5PYD6uK0oSe7Yc+AsujfKcZqF8NPKBt2ud0l3G1AD2P1Mg9aFLw2lKXoO9Iuhjk5
m1KPmM/SEf2aGeQBMHLZsQ/mHf4PqeLf2AJQHsxxs8xy8n8fsNElZDELK/h3Lk4g4RBH1R2ovJDk
8B/m/ux49fP+/ckqeZU4GajOGfwhwv7tSFsUfAZJdHRwl683vBRXtFaVhE8sCjPcJf3bqWdkASU+
ZVnOboNcSAsZBA8Qozcc0lbNVbqpONIJP/9luHtx0wKflqXf16P1RRWxf0xxLpH2/bGe+tkw70Ch
YxQ1C7up5Vgz2tjy9G7+Tcehb6FQCm5WlfsAc9Ldyp3vw/UhAWuZD8W71xX8N7DM9JBUF818V6D6
HQoZ2TTOhvjnidmGrAQNTX6n3X1pronIBdw19xKtgPWtXngN/fpIP9wMNCmrV3a9b8bv7PFk7jfa
JKPP+G9Rxroov67KG0kZQfe1aPp45+HJBx0R+rqp/8ighhtEqpw1YhNYsl9WFFOQJlAeJ9/PRDr4
uil/YaIs/BQ/of97Xw4IpTECi+4/LGuGK7NLw7RWMxW3AjZVOWadP5X+RJevOEZrCzdfOrpeGJle
RL/QMsfRX6kYAscaJTnT7AiTKkZSKVXZTDs/q7Kf4wfrIS5RMkAEE4V3nCUKZdvvytgW5J4+mmmO
4liUjE26pBJpA8nffypjV+/AzYcgzXnEbsyuT1jPHmGzsGp3sPZyH6EfXrZ5tufaQyy3V2D3+4on
aQMYglMVW9X8ydTfCINYUQOfGt52Lg39iU+pTyOyUG4ZDFVyrfmFudeTVbapaUyjkYGG4BG6zkjw
IxW5wYVRxeHhx5J8CBFw6y2hInFkpmrjZzMqV0Z6+Z8EXQHkysDW9BrIWjbq08el23whr9R2YxTw
rDbvBBFPHgVr5IfRwxrbh05JZg5gbe+OCMcSNfByHYfjdcPGBYEdgYRN8iUFborB6mwp0AFWifrz
3gYXoxfX21Qp6Lg/VzDc9L3gO13ZKKJNeyYxuYV30QR+1mK4kjAQDrb+Kx4r0d8GDIj3dDlF8iT0
BYYM/d2/gGbUe62lFhmU2S2uPfXM/8ulRNDnZ4aZ428pV//RFVJ1I3LN5FqyqnFKene+u68w90+2
inhd8XHaq+z3Ob1+79w7Z/YvRwSt+TjehPtFGxaBk9ddTqOQ2Q0x92WrAUd7UDes85sXNyL5lKGw
ZDnDd2oMRGU3eKsOP5Xuu0UWiBCOlXzBDXlow0a0Ug96D3rMbbKPt1PiUBZ8f1VZBQA+weOVGqFQ
x9EZP/rwDHKW+JTuL2in0Izhi26LqxAmKcoleleqn6HaGgv4aqlU1wpcha5s8YTeVAWPLph/bBT9
m+e4JxYfWmISYNLSu1d0pSGu9vB1Tu2+6l7Yr6RS1lY4n62Dn/5UVQZhXwwkgWcUeRBMOMkRt5g7
Vj8KCWnmM91luqCgmJSQPhvBJ5MDKVCQKUgu6/nIsEl7HjEYhYls3i33L7pYM0Orlile0mFofQpu
B80oOBAl4EqEtnSu0ES7368EypovqDGZQK88cWLEMeheopri4s7thavmvl4KIA1Kdd9bTp3OfTCu
xSUipFaAjeJXXtLrMAPhMt9iiq2pNgFqKTixF1rxOTl6n2TAlF5RNZjq6QNNiyz4nzgwVnG9G92I
U42MD/k+A062fVv1Y08PBPaM+eDarHm0jHzXTRreiYqcF5zHrFqgZcri0hOXzyypF+5P5lMmcZzk
XIPNP/lqEkPC5zN5IqjZl3RH/ikRVbVmA1iF9hVtBDIMfDrJDUa5z7xa2Ku/1goBk2qtSm7JHIUy
y9bq4MOipt8XyLUkiEaDCo9hIiTwfx7VNqQUL7wbxkPpMqOhoZeHBYFr0y8/I0R0ZUeG3jEirwp/
s3HgKZZu8TZS1IZ9A/FedQPhcIrjXLkX1P57cLYXNlti2ful4nniSa47DSeYC0uLL+YMZkvQ3+kU
ebkL7gPZ1lGMZBVVIigzazqLyXumc0TnGITZH5GDOQ5AqnQVBI9Xoe4FtRLW8uDNpbRd1cEMzab1
z3dEHzZHnLeIQvM9tl/tRLw5sroxRbDgP/5XrH2N9FVs90KhKnQ7gaWKqZDR/C6MaZ5sg+v6nRk3
CxaTlDkrb+GI9NM8Pq24gUGHCJP8r9LrJi8gLlUnBmbNfr06A7bbO4F4stXgsEgOM7g2AW0EHa/M
a2hYzgfR9r5kQtISfk3vY1I0lV+s6yHOyZt3IroLshIgz2Zhxa3tisEWB9EdXs3SfJHFNrG/k6+h
NsNt6dAhosAQJjwMgI/K1mFQ+OkM7IF2vjaPriisj7pQIeiyZ+j+qBx18c/etaoO34T2GaDQhK09
TZOxpDdRl324NDWjZH5s6t5PIRq/Q1tbfOPd9pSL68HenSOHrVTATIez0UjnZmHwasjyj0bvkwwv
NYLfbuUTWFwZw+JRg2GvrofxE54jvHVh7+KHCNDiDEGxBDfliQrXLJiLToph3X9Z38WmysyCPR2+
bXzckJdhYB5y5VmshXr2pj8YAeIgKmmZ7VR+b0nFGz+5kqOYQqaAf8AS8EDJ1ndfsnvD1PlIXQuc
rLo5Bh46EEg+UDvfgs6H5dGgzatD77oj2QBRIZ/3s/ICBlb1k6/nsWImbcqkav6C7x9KZ/SUXaBm
Xp3NlAmlKI1C4K+XlOIGp3yYxxIf7IpvEaot1YZ8RTHO13tRigcBjTXuvZAPqfljeuFw+uPljpPb
cH48w57SGp7Ppc6VnLmTSgXcnkBLJbnpVhLB7GWc6NyzsdM2TQZPrZoVm9f8LhjiYTC3C3K5LnAw
W/iDbJCw3kRb/TuyBnCAAx07k4q7J8rnGLdqa2aJzvl9LgD6YFdMAnaKeI5NCg2RrkMMhAwSV3N6
FRGV4L42wHnFKWFF0rTJh0Vo+cqzYG7tHt2LsmyEC3CiMszcIpwmp/828EOvO3pNebfCLx3eYy9v
uV+nvQiDO6pjSDExxAPfKaTZ+KK9AOfo1Tbu3CWhXp8FPyPaSBkbOqNUCOuRdENefgakdgBsuQtA
AlpUdo0ddlGOLHr1Yow4LCvOvpzEugVu3C5aac45F+I3vEBA65iaKl/k5XiGK9tO2oGewqRvpe9e
oPPiGBqDEluWqUvjvXPK2ynfilctk+ioyKxyyFEqbe29VxRR8PbwQvVUqWeuQS1SYYMYHV4hVyPR
alo+WYuWNbgtAE2KNwOvTerj6QnWhr6ijmCN1gB9TszIiWWj97vrwu2uumEr1Uhy0j1RpFBUrHe0
hhwgUoUCznZ6Q1VrczuTsJsvDbRY9U09wkBmqqIzOXXu1rtGcAYow6zPQ8fuOsZx9ECSnyQdXqxm
Jwbgq6xYVHnz+lxXoYvmWC/wxu3T6Mm6KPa2FVzZof7A9MiJ3Jfhs0h/em4RdXAoR1EiemHrjhXi
+nzJGuzk+g1V/JSdm9xRZT1uiHXcobZ1FlhpIT0ksFzNwXn7D3Rc628C0wgCqETs1rSRklKK04UK
Amh6UA8flNzNtB87/hFV9LGP1JUF52jHZAas2OJfACHtC6Kd6NXbZq4mUG5+H2pgxQK2IDJobu/+
n/6MY5zgFS7H2+FnTEKAQwvsREgcL8d7yzcnRpF0vtKqgGMqzgbghtKEQ6/wlVCNpPcNWubAJ9Sn
bMlaaGAdPSZ6cIXgDwTeyL7Ra8Dp+YjhJ3z5hDz+dyDLXy0NYn7dNSmjarUWjLIBjKMxt7OGML83
ORlyY2oIZQE1KnKNeJIPlbuyEBRxV7g/WqmGppj56FLHRfp2axmd3XiAsaaWTjwW3V/6M9EXvZZm
MbiN9+dNtZaWEl3d68fNZgvGZGKJUUJEOi3mVY31khLwBEhaz6J3IAYAuBmMoh4XyK+UYZlNhHna
zVaPRlRcTboCzLdxWySCoxGrLtjmbtQTZbLCC2qlRUV7/P2EAQtkGTeP81nYEN1A3QRxB96G/xuG
00hR3cwXDHQCNSyytb1wdBUtEhd87naJwuchUbgAaYulUwsKzr3oldLRNdyTHrvXpZqfIgRTrWSS
bXForNivby9cAVVoza42D5DIWRA0ueul3fEN5GExSGCItDTBsqH8nT9qvxJbhCvcJjxepXD9ToJH
I2vla0oN4b82wND1T9oZovGD5QOqtqe4kCD9ZTcn0gEJQ/8QuzSL+l04SUvXnl4lQL8sUFgorqvT
7fMtjd241IntuhubAlFERc517DsYjwYTwatbMN/ls/acL6h9mK1+2rI3Dzc8O23EahaH4Ffb1mJc
vsO4j/S+UT1+O/8hOlAa7QmMz/+h2Wgvo1sqvfQdgU91PJDNrSnRG08rNz0GxOH1gIsoEGp6UVkx
I5jYzB1bUl/Mw5wuHVMvrBj6lFXq2rFBARorjUZzBnOXlPsWjzMLle3H9ocM4PC0W0JBip/9uetD
GzBlmwLS6GcyKIPKCaIVV+R0iL6c9NL4nYbFUMDORqUgz1rotYQbXw4PDPjwbOBXoW46sNXFGxyF
cH7bGMhtyRASwF5K0uPkPQNf37Fk2irsKMzGxTxAoPiD2DtiS0jzpK7IrTHSTz9QvRV1E3RbXIbj
36ERn6/J5JcNpxcp3oZnpRNwEAfXINEdE4i7A8YEQvoOScKMSIVIxitISqUawnacmVK/1+LDl51f
9zqK7g4aKJMItNupvDquf+r2vPbXkmCwktCAopnuz3oSgqAKkj7o9DdpXxS1/e5X4idxW3qLHEF8
3JRkErZ+Q+jsvwsHHUGFCrSA9nPwhx3eOAXug1ZZIoP2itKtasxFKKi2iL81os45wi1Dxbyx42IZ
5Ks9hMJWnHJzJlZTjWlZQjzMb2GoVqJq4ffz7ljbe7nfr65qEmsbbIbweRlv/kRjn7ZbDUfe8Qg6
lFXqWssy2EQVc22I78h5VG3VJDyiA0b5Y6HWZsICyh4454MosbF8ryHmlm0T9Cm1/YlXYTrg7/Sl
9fHFqEQ57Gpso+Mx2YBL9X7Fyuu8dzsgfC5xWDD2Oo8cYmwK0tB6ao2sMRKq5ZCekipRtZHekRU/
AS2jQB9pnojUIl3x6FbZ3hJI1wUu/AFUlPmhyd3s+ouK1/dwNHa6FPYB5bRkUfGQYlhANPQGG/tk
8uQhMRQhuk9p585tsMWoJhKZOvm0lBM6hDO7ZnP+/TDXeOq/NnOrLpQL4YOWfImuwwgBZJmR4OQQ
BoB6uUafX53FymBHqq2MoQppUwBrxUEC4WRFDJq5Vxsb90PAS3gSjMC93i1mQoMhpe1h9EdHjVHe
n9fQSmgLQ9hqc/C/4+hkVVO7+sx9vNCELTH7ypxuoRPPqvvRKKaMWcjConFShMOTSSlrkzNtDxcT
eXHUYB2PiJlp3iSru2WOLvtu6opdTXpr9sBKdAXosl9QFwaPO/UpxhmQwdF6qKeWPuc8FW+e2erA
RyCqGIJbM8jkIsOklQC0iAblVpipGVDT9jePBHHTppirP/nB0RcltqxnN0lOO+b990X5zUPINFJk
SzC+da1JdYvbJ2D8p11uT6IU5WsCJoN2RlCQXTQRGQNqYbIPUn2lwtxBxWSc2Et1k7LyV4E2jgxr
+TAXq1WXczvjwWTYDW0MErvFBbQaUQKiyKGm6UfpgWd40gIt+SrChSlxLc7iNFF3dF0VI8bPNVLy
Mh1sccqUgCBxRYjvRsBXw6pLpgoYK7L/xAyz26ivkB2inFhAjhyyrhqh9qTcOuImIGgyrpVwekRo
AHO2+4GRwXxtcTYiDdvVs89uMVBKgDG19y7RVcWrB9ClUD/oiM3I86a1f4fg+Gd4JAJfDkrdCk57
BFe9HbH0EKMTLaYCNod7j3XdquY/zooLab2saD93dTQc37XoZe3BIqneETlV+/K7A8FbuFc7Lyrz
UtkBwKo1dLMRr0XT89W+sr7I/wnJWRoGs/FiOfNud46LPk5QM5pfQQXoMCjkp++c4Csu/juJvuz9
Ki8TWHEvNYnc7RatgEKBnCaOK9hFz/ylQW9zTKz9EKOrJ4gfKpCe41oClZuJLUqlQKB94doF7SlP
lJ1QL40cZgcVVH90FZYCoi3VqPe2YIPwWc7ZN88B9C4KjSi8ikQqgNMzXYelqaraV9zd8W/Cwd7x
NL6h5a1CVqtOSMSpiUjJolcAHDj8PwoPv+0x/2pV0aEmejI5Ha6Hco+yegPi5C8gqu2nn7fqGVrq
VB7MKWwGNRd7Sye8ezDgSsoS8FaHCpC+JaSEiT9WMptTg9EFwzPKz0Z/LJ8xYgaryNLpQB0ZV76N
TEKf7+GPwXu4FzvFcqMDFWtGxm7cfw5XJ8ApRYMCftmDnoth1LpNCdrqahamW2ngaKCeVse1BYal
mahk/MNP5TAnJPcXsZ9tZ0WsfPDFuL6t00G21ki4S6Iox6FJkzQ9msJUHEeRq+mDqIjFoc9K/VWl
wLAjkoz4wi8/d3LsUOt137tDGkNXFdP/Aq18D/nTSWa/RUuTG7kUcabnzp3yGGf5YGKZWxSrFdqs
SMKO8yIdr2JuEk2VPsM2EO56faSEjjZVPnDcrTB/hX3GT5CmUGosfzTKn1x0xcK3k5+IwSFSYPLE
1LGUK0LhAG/q97nv0l/M1RUp03SlABZ1vyKGPmrOBnLgwOV4IhuVAIdD35sX5QtFBnDIStDo23DL
/F7HTY7iEGsjn3CTfipM7DeTt6camVzm5VtUZ9hGIKAoyk/BHAJ09c0jgZ7VuFxwLgiFN6liEapm
ZZgYmYgolHBu8WI/GevzuS1jWFOJ9jYaFoVgtqviPLVttcsLfxRh8wNCryjY0GMCFcZ917HCR/wP
tdZIesAejd+NeTnpcxfEKP6F7dehhiwKj7fAR+1zoNyAsuVHvIrfFHiwxZFyvtaYxSrsKOdezXSi
hKas+EpOFDivlndsccUdS8OaHEnMDPZLmb0ZjjFnLRBGXFY813zSzX3BxnA9Erud67uHMHPE0n7I
OWE/3UNeDaRSz3ysR0iOfN75aAa4G8hkaCgw7CCyuJ5CnpJwhTQyYw0Llyq2NZO70PM6Ww5ZN1v/
BkwXpSKE4f/abS/CkOtzsB1FNe+MZOReJ06vfrpyw9nStKdJFrz2J9DyUM6ORJaEp+H6zg0Bf7B2
v4ojUzEWY2uI5Sbb3jqhf3KHPjjs/mTx2YPMciFK8SiyDNuJy8E9/2T/qsKjDOBq58SWyAiY7t/2
OF3IswsiRoBj1pNMM97YhoejYrubvQ3W6Hpu9Ky9vhU0C15jfCPnPVDONUCfzcBTY0S1vTM1T13M
M2Hk4z3GHrGi9vBs7vG8pUjJHai0EDYB7SXJMse0naPfb8qxzW+w8UKwDsVo77Ncrm2YA2/Nw1Nx
4dnnW+E8HBLOyPkE+iVGyuCzSvx1J0sQsc+WU5IsVPFlkHNLtrxJp0aBaRC0G8CQjrJM1/6zp2e7
kcoJvPU+5nQsIyTX0J3E8VdXj0bVr0STt/6Ox7q5EmVvtfLrEBjj7YLPu3Y4LHbhgoc8fZXynKZj
irHbCYaBBOnmGQ2kRff1q9PoMcpOOewgQg/MSjg09t1KF1946nqaA11zJFmuq1X2ZGFX+6k92/d2
x15+4z7rUHI/G2YDxPuRiPdMsMizTKgtPxLu+EChIqsYR9TOdVzOJXMmRc8OyC1F1K7FlkP34Puj
NpzVZEiZDpVQh/GXdjl1kyIw577ihMT31ceZeqzEkog3D6Z/kCzU+a4GW67kSfSciFVnu8Yfk2mn
n/ec1v+TkAL0dcfWSxK4JKS6Xgh7dcaU+AUf1bYpEEazKNHvBV54GhnLZRbKYKAOilu5TB58bKPp
EwXdfUKXG3ROYMy05vgnfUfoivwoQC1zPV9TmJbzQoMfN8N8uOB6Roc39J1QHmxmiury2bWNSZjx
fpFXcxkJ0+mL+95YNa+2qO81AJmv+DqFtsGQeAJvoCGirZtB1fh/kld2ZEcCujL3HVKNJbQXfdBW
xZzlxzeV0KPrPnebcSqdLYPgyFZX4SHUhxkAnGTc7gc7pv0oyzlOQrIpAEwuAtWTa6QSJXsNsw7/
PVAERZI5zmgI/FUW7hRuLV1OKLwybIIf8dzLf6Rx/DnRDUs/sTWFqFPxf4p4DP+JNPbDJY50HMR4
ZVO9fJhNq9aZrRp/p7qL8D2Yuh1KqTZ0qIEBRfmbh6zxP2mBiSSk4LZ/d/E4vUOTa2ph9yh4Domw
X420osTIjL6pVr+5fv8BB1TSdWFgRbzFB5YoA2uyaBagUR1yz6ycZ4ClrtWkhKP1jPaVOGN6oCZg
UM64rI+liLntUP7QICN7koi2WfZ8U7n7YiOwivlgbdyjPe99O34O4EGUvsy0jk8dDhJ5WNad410P
7imaT3pz6DtFHS/5ahaINzbMR5UzUnrMx0GgHO5fdyIKJDcfyeEwinSP3Q+Z1vCIfYv5t4EhI0wo
Uz6ijD5EtbFi5RAS9BHspHfMy2FotlyaZ7olwV7KdUpqFxk13vqVHOE0z0Zq+2NS5vRXiaYj9WlJ
wlS6TQQjpEfyyQgvYKj5q+iW26XEe2LQXB0jcu2vWMTSgAYT1+unjB7zjArLPgtsN1xg1C5IVa03
hC48ChsRa7TO4g6vPCUXAR4Y0u82FiUgi18+tgCmtVda64cxs810fsM4lxKUEGtv5eH85w6h9ufz
9c8AB+hNR3FkzIiMEZkTnJ7c+rrIcMVxCpic8i+vMsBmO6n3YxRz4K2Xb1VmpNkNkb+tE72KJK/W
AoftLv3Aea8LddOEKf2yJqLpm1fYjOzeuWBi2lru43PaKoYxGYYJmAwDNeaH3+1WyufqU8ceyg2y
sG39szktejXqZXr26qWdGm9XEv/C8XhgK75vCj1krYCat50y4nfdpzbCosF2WwdLNPnf+nduBZJJ
NZZ5dv0BYTNWDaonENdnn6ZuifP8HxcvCSb5t1UXeuuoI4k/uPvDxnZVrSqx1LJEuwD/T1zZkhaU
uUQ3v4nsXxWKpktTDvqy2ZdjXQG6QCbUZda89pwHzMFfVtAJ4YzKubWLCcrbBZJVbFGtEDgVoJxL
vR1J2NHG14Ha4nXVllQtMnZDHG2r6eQyjabw8o89sJieQffS0H25/Y3jr7KQY7yXUxQTwj7Ukjb2
I4+CB3w8KzmjWSibzel+GxlbM0tAEwSNnfmqaJWoU1YMo5bkWKnTiW8dF62AjhmdEbx05fITN6ou
e559WqJlet7EYbpZo6fJhE65L5w6IXOVfwv3VLJm+6cRLNmQf4Up+mV7Yb0++F8T/4iO7/xjDs+l
1fuD8vZzM92FO/K2zoTrrqFYKfAx56UX3xDrRG68uCzTSfKx0LlrECfHDHXKI1Fh6qwIWhjPayJ7
/74xL3uoOE3KlRD6dmUSU12N0HImRO3MT6IHxzqXHSrNZCjPghPzvABKGml9z4IAFUt0QHdhiRap
+a+tsNPEyqKefPTi7qSv9nLuN5Pdh62GpnWtbh6DVtFprHpw0F2pKZL949+ClF/0DXKeh5XTyPwI
ed6gWRl3OngUCssp4NOu50u51AbW3AK9Hzl9g7N1CnTr4gownskNeTmELTKWVTKT2eIfLQ6hEvzg
AMZZZx2UgOlRKZBWFrznOM2ptvAXlMZPOYAU1lhpvXAlvJFvFC6JmFieFlDxcVCGwbausR1ft7Jx
1W1UVTqGgmzW5rcycjg5TG6O3vv5t66ZnktO8rhBYZsPjo+BaiZiEWXn4Q6RuJKC6g1rSuKexH9u
FgnLsLBtpg6PBdzE5jED7OwNxU8PlI0rdJD8NnFcYpo/Ave2Se82ASaWSXA5hB9i3v5A4SoIscQB
7k7Fm3+pkp/TwQ4v/R+MXi1DjbQXorSZjtWXhJjm1+I47UKHNyPvsjtqhiN3dHx+LW9HbNhcUyQD
nBra85ezBsDzmuBM48D9v1/ZsybXLoC4dh8CZjKSKtI2CTShKlgekf08JTlTigCeFGzfmC1YfeRH
8ktNCfLG1mIKCS35Cnjv0Sn6prjQsUCB6z+aLuK3TRT3bJXhSE/2z/2lWZu1S6bvLp/lUnlgq3cF
vM37Pqg6ys4OVezSjEHxPu/P+Od6tYe/te5zUJVSgOUqLIfoYpQU5QGcQNgP+Oq09J6v26l6U/vT
H/Zgou7ZpaIrq2NtQOOWtemsSB6fMRZJ0iAKo3CyFoHNOi3hORXpybsQSPRT+2leAMbEisgGczAp
fkgCgJeIMMNWu0UfMyeOETeGlXkGjOOMVV8G0ay9S0d4ekLF00nBeOz4cEASrgBzfdWOOd65TSwC
u9s3gqdy2RaBoatUimhFBR89R2ss3Uhuu3w4MAhgRs0AQ1um+Y2fzFRI4XAiRiW1dbGoUJY9et8g
PJrB8GgFhBnSZBfTpdrlRaTc5Mmekd1fndcILcJscK2hN8tT1TOuUl8n9QOVfacnEHm9DcXRgPqj
f+k6cCwW0AUyABn92lgNQfiFNtRh8UC88iUXaiAzxhfgtrlcrbBITHM7L1kem4pjWowXpJU4Evv8
VMagBwTgNWZAL9DEKNIiim9Z1ZQL+QipdetrBKsISpJvzHGFkV6KIFOfnNWtC4dgU+0bGxz5NfgW
yRqQe78mYMKHJiS9Sjd79fMIj1Sc/qjfSLPPhiK4aOBI9ECsOSTJmIJiviKkM1mfD2WW5mHK2waS
IvIAb9PeIpYyFc6XKVgj50Ezjx3CwdB4fAdEj+sYswLAVusbTzvGwd/ASVIbGly+a9kBi78faGaI
VM/M/kqJ1HYWDn7SpW4WvgsFMGoHp+akHrc7zoISYW5quWBG4QGKPkoUlrla62Oc0S5+JDi4AjXW
mKwyo1NZQmAZ4GnOCGffRJzGFofiuXzIGTKPodAg5uwuYLskDljULO8cDgqc8ZYuCE5tKHpmPFcj
OwRcxHH+byP9N2NF5m6e37o08wiXvDwjfxOq96othg7AC4KqTCM9VkXTV59JINTy4YPW3mMRT7Wa
4lA9tpGDAgE6vvTz4eBquNQni3itux4uvMHzoKG0mV2QrAaA+ttOVbKX+F+5ODwlCZLzvMJMfbPr
Gy0lR/Tz+tX+gsfJRdu4OfbFfCSJc1swXjo4YpQA/zMbUQ1+HMoe1FpFHw6KdRWKk2309LVYgDQA
mBuvIk6amq2+xWpsk6XPAIXkBfsDtcbm6u7JulQHRbPhN0qldJJzxv1a5GJYbKGrLor/0F1CB9Mp
PMxG45Ft5fQ+Knj6sra75zMG7leWEUdCcP+sv1ZZFQ/A39uyk7GVnZ5e4mG5YP7KeOOyMzSnuIcP
ApZ0To17JTO2t9QGjr/n9YQQwmhX7YIfzLKO1gfrcn6M/fL1WK4Fy7HKOQ3jR4I3xPZLQDcDQrDV
vvTTOyaqRz4570VlnSxl5KndrKUjW6GgSf8FnWkIhiP2scmeUojM+f3qpgy+YQlVaH5g9OQyyhoB
D7+Y03QPQnulAnbmizH+vQaIHJbDXw5mYlaj/IbWZuNkwdWpg/NR5NvSPNhNuuxkHGyvkb+WY9VY
D1rAEfRhhQ/k6MRCw7v9BUHWD3iHmGaImr9v/9ZaHu4pGzg0l7sk1p5UNppOmwmSAA2Rwvolug9X
XFJdJtOUtAiWm2AJa78Ers1yeFD/rXgkaWZ7+FQRCpZp+jQVr+N9D6bFBW3SJv7uzM+86ivXVq4F
uzcJYjVSqsSfgz11YUhCAqKZIoW1wfA6weSYG7gM6Iysgd2Gw+DbtsZ2j8NugMzHtWuSNL1m6O9M
MzW1+PGMUYCwdlcY3VaqPLZ9KuOCoTOrC3saGzAJSUYYL21m/xkGWasX+8T1OagrSc2bw3Vnome6
1PNwsh4vTDcGGeQfwopNspOtEHPAPRhnFYNdTqozfns2+gzl1X6GEcJyqU5umKu0FRFTNdsR5x5S
jXGLDVRkLKvF8P6trQ+CmFZSVBqObIH+6OZ6VefsEXVpcqHIt3Y9ITKqqS8xh0eUd3EaZMw0wexf
60iz8fQb+ODa9EUhFLuJdikL4iTy9iCamcl1KJxNFSVDDvHqfzEDyZHlyo5eNo5S1AjwVY0NoT4Y
kRF4NC7YQBoJ/CzGLFmtQIU+fdr2kNXrI8/mpp/piYSJIX8Kvgx29CbTEpZVXipC1n2XXrjdo2wF
0W64zrwWRWS2fDil79L9msqzOwNO8Vp48MI+sL/15JtCB5QO/tedMX+mz+IQ4zhSXvsrd7vB0mXP
5Yuz0fy21RCPmMX6g1bkCX3YXPeFwulLBiwhQ2qBGqqLWwfIwlK8phpRIfdntv8EuNLrjF9dSDbm
LTmVglqX1bTT27hgUoY7W/7tBUrEwyKE6wxaiOaaOpsuEHrfC5drpgGMkz9snPp/uhecWuGwoU+7
r+1KG86MLX7PKw/XpoNl2DBMdvtw2tOtVdy7z6okSRjuddYgwcLsU3jmjZnSkqXNZHX92fx4whrZ
1+MBnaZ8JX8/hAMP6XNVvxKLpwYjA+1PhR3iIEIDdUrKFGUbvWa8ZgVrOAIfovjDTQiYdNkVZU33
6PC3fV+fGeouJBkXZxoz/JTTSnyue1B0kFnmETqUBwg7CSF43HyH9qOTQcHQFww4EUz/3h3DTTW7
m9t9mOTRB5yXRMRIbVXEj0u3M+mdiZBIZPSeEoqmx8uwnX8YpG5EE5tv4XjLYvUXyNbRIedPA2Zx
GIFeRcMDkXBKCGB9Q8PvHBc+fOBiSxf8AFC16o5SZEzG5EwTxXgS3IcYV4bJgPm0NoFViHzGFPzI
ZjSAeYrpdoNLzv0WUdYKeAIgxh6LB0Rqqa1RmdqJYdiWQWZyw5E0rqYcgVWPAQygBySt125rKlBv
l4oGUe6FykmnzL6l2pEAaQFjZYVPBBWT1XNCyUHKIvv9j82fsL2ETbFovyyLnAGM0yFTpdxLs613
vNvb7t6zS04dAic/l9+2Rv61BTMWCfIatjzGRqKoVphrAQlu7DCB2Rkcqmd8OboDOhi+pFSvP97Q
Hl7qBij7UCqiv6lArDA7sS6n09S9/Oq72NhWftp82IHIBXfh12ABtyNU76mca6njWRVJGea4hvSs
etjDF5JT2OgGEVjnwLff4l+zKJgpi4Y5X5X2KdsY4bssR6xc9uR3H1Rftjx2d83RrGiNnyekVYBK
vi6y7fqBCyjohIC7ZMENkUgPSzxOymsG6yJTseCRmJtNOSwguBu43Skl7v+sDz/B/Q9Hfqs3rlgf
Hg2XLb/xCv97imGW8rb0aatVqKSXAsgrtKRv0O443vDwMUaC5wMUhfU8CJvGxIGR2bY8dJ1/x9C8
oP7BjxWCTSY0AR/+48KSjjNn78TLe2Iim03x9VNXqFkOuculGmHul35ALVbCjURM6khs9s8n/TVf
5x00h/lnU2c1Wnr4O7VuyicfAI5mCC7QXwqR3guBwcNnSU7zGuSfgka/qlzP17sdzkfHdKGPIppD
W1HbtgCJCvZXjSnfYfb6LBzRTrSQvg9uKiIOhNy6nu7KmkV5/Gb5MvLgNLEpKRKNM6oDVH88OYdq
5XNpjfFHmm4cSPFMGl0LHJb1Zy1FV9vDaXnZ7gglQKi/EYJs4II8Q81yXKCwKTajnrOcNzVbrFv3
aKK/U68HnpkW1171urHhlIJA04aqhu0Vy8KuYL2SL3epmmOiItTUHwvNt9/WYP7ybgnArDjuf38y
zTnvdOyMx9Ai1Wx1madU+jzmyeVAiyE7QpmYK/HHYOQPBiBfVTvpmznaWxCe0cotsZdy5qDw1mMX
Z2D2e9+fgcbjZ253vGjBCB3k7VGeRDk8pW3KMd3W5y/fnRV6paekOI4EchoYGUd4Z3sTrCJVw4mq
mdbPmj2nNGpaMEXLdBfmpU1GSGip0YSTT8pfP0K+kxk2oL418oHIbod9IStJ/H2jBOmDOUkzy7xu
OAMVDW+aysYyluH4ttlAeWP0zUP17b7tz+T6jhcNsu9VNn5WpsoTMDwZZE+DQ9kwAOYfh2VyReak
ztxCTn/c5yI3NfIbngXb345kNe484mjJoBPlyxyibVXPlVUb2UZWusAl7AR3jc42pc8tQu8vW568
Ft2WUlZtkSm2vghU8vU76JN3QWJf3kQ/5uczAAdX576qiCwOiNpp6ifNeg1U4dg/oiE4M0Pr9mAQ
LYCdv4R4vuXjhi3SFbAcgWKZyUO4xQbpyJrAsn0/WpVP80Dkh6L9rVEnvl7nyJ1or6b97WV2pCnb
Ro9Va3xxDwgVgIl4UUal/y45qID/MuJ5wJ1lXXzdSRTr+QkprDxhR7sG17kO9EVANV3ML1hWvyBs
3kxJeGOSWP7ypkbzKexL2eJL5wItVUoWGLagoUOMV7W2qIWLDPbRKZ5UsEflIK8+vxjcDv2Z/NTa
aoiHqowM5rSwe28v9GWuRIH2y10HSuTeJ1wj8ScBFNFe+epdmGZXklcmu6ijqgvI3U8iPLH2tig7
ANlGnO2c7Odmx/6F0BP2cB0a2NjYTX113/NmWdoAMseEHEpqunBhDa2F2WyvleuMbIqfgPiufpWV
b+EGSh2x/0fCV3KdgmbfQtl4eX9miqtjlZmqfGYf4F+VrvgR33Kw5/BoBe9EZp/VkjUrrnDZ0f2d
Wq89jVgnia73JwyPtzx9yxslPLN4KK3JYAqUn6yCKDm34OGiYxU4yImai92p96MrdfIPR0S47mPi
RHmmIc71l5GSEHHzkuP4oomx/lvFToT9/UxYNL6HP5t73LyAVNmIEvWqwBl7QU8TKkZ543LG3Nq0
NRnHVcjTz9E7hXdy38fKq5UQAmDUA2n/ucJNHXjzgYh944iw+XNddl07JfAi4PvK3RmjqtpgNL3W
0YqSLjh70QcAPxaDYxVdD1yBnYONFOjXbIYvMf82A0HrEDI9FdWx+AaOb/Z3eLgOfMV7c37hQNC+
c/V/g96sgSHmtPPvMws78yGwvcVSWIY5sJyRis+V3qbEOCWhm5gEyR/iraGF1OzUQnJnSRZ1z9pV
44yj0oyQtIDnMhiqGzPi7nWl8Pv2s1yeJSsUqlI6gVvjQcLpK/xk7II2EVNf1CVZ7RGSUqf2b5B6
Vrxg6k8RyWoeuPguuiPxaEBRplc177UTobiBEmv2z9RgjFQY8QYMwAv/C/5qkK1mttuS7sECWrz1
TBXY4I3bP7J030u0Fb+zG8WviI5rNyyLvex/fJEmb1JosrZJi/VpCxGKrVtJS1luY21Bp2/HYBQe
ap/4dPRfv9+h//wBEbkVaPZAeipjBP0RiqRYqDgSx2wP5A3Zm2QLT+F2S10ZQ3JvmltkFqMSiKY7
Eula7GJhjybdZ9KlByWdrln4KooozfMNJemU3YTWbzVWAIPNt97uX7epcqwMk/yarrn12AxgMVH4
ygFs6tDcjVJXQicb+qGiEcQTx9VGn6Y6ZMFV9TVXvNumGsOgP92QZKkkzO/fD1T/3CFYZygz10Gy
4QvPHqrHoLnW+ONORSWe4G8o+Ovlma/4ZW6D7JFs9pVkmMXXCdUq05AZx0rZRyXtXxnzBBSGJMM2
LFiAF0ngU7QOYy0oScalZr68qaSDH7PJWVgi3q1yuvjtLi/ZNePFA4CPQqyemDLqnhw4RJAJ52cn
Z3GcTV6MUEPwqdyAqYpADAhzk/xTIAlVmYb8h2jSTJ1e1NDlJlY5pzbNaIBBWY3tr71kjWfHTvTC
tUqiXDHC/ezJuQlVpBBNJB+1lBqiWgTPmehmIv+R6szmGZ6WhD7KwkJYcLY7RCU0XbJnVoKjKWPq
iqT1+JSmP31IG4qMcEtUxSExLvgg1NlYGFqtDMvcfOA9sVz5+3IGNODktil91MJwDj9MkpcZegWm
YFFkyDfLlJ3bHmnOa6seUqkVyUmKBXqQTT+i0EyBn65DEvMWVBaai+NX0Q8/s1buAKmranByr4ec
8DNvTvmvR5LosqnBBSTZ+1PlXW7TF2+Bh3JAB8vi5f3D4B17TBVDFX+XIrRfG/5M3F6z2JxcEEDu
R4poF5aa6Rn+k1Pk2nBXVoqOsZ5zwzQ+Mww72oakILKWurwYkP9DPuvmx6COt3ETlPshHCJDEw/H
JTgbot0dhTvYlL+/8s4pwRePFsp051MQIxbeoScN9dcGQez44P7jBLjeGVUSTBmKidB8CJOrd5vN
vfnFGtJPu15OJacpj7Yl1ntFW3VQQj+TNeb/JtP8HqdITxBaG7OVyTruhsBfrwl1tfXZmqYouQyx
aVaU1f9mQCK57eHxuuTZxBrNELW5ykbH40B+lu5XhqTlTlgFiUQZQ5HBFptam9OWADLMI7Bv4iC9
NDgA2+/dByVYOKro+9wHQnVUvJLGP9+OxgZ7+aP031wRaN3eN0JSPO06+P0j7Yinvsd/0z/P/LdG
y+0MN00RKkkIBciguMPDmtl/ctuhwzBTMltW3QcRgMBLE18CBp7b0xcaHkGNywHXy9hs1ttDnW2F
hJqqJ0wBmFPI+JDH7jsX5DWQ/5KGpCe9cQsPXtwfMv59IPIXV7AbdF/yUwkwXxOx8VP19LinXa74
9z7XxgFvnBfLZ8GOXxpOM8bpeGEHyb/0tgJO/JxuJ9QAOVAe3ARTQA8vsOVk9Bh/7zumdrNbWi5W
rDDVN82s2KK9Pym6qxk42VicHnXqhBLQTgQmE6MZXz6Kzpx2SquNBEaVHlOkmvkLjrjaWmecF8vg
BYlIt0jFJZJPichPMTRUuPM8uzKzHgdPkr7Ao10m9riRwpv5TXm22rQV4QIBxKwv6siu7vaDKEmX
aNEpIm/oDnzoKOVCtskn4BnCzi2Mn2EJdW5MJxxZMdPnmZKwME0RruOJ+PfhhLgRBQfV7hmzRM1b
p7AfzF4p5OfXo6ujY+5g/QhKg5wQgIdxKF1zM8dTtjdwhArDwIbtZ90WP66LRMvbKBcvvHgZ/GFM
9RNNCJ/izKArLE/20b9XFpRduns+K3g7C+9Cj7bRV7xKnj4jqNkc6BXD5wUnNcInD5I8UuebAH45
2u9oss/Pfny575jeKUSHmShrjML+G3ZQ4mPJgzTCtwpfCImDwXFB2Rmt1EPq1mxV3/I4i9mJz5xH
EEuB0GZrAb5hfLzC+9B7BavhadRZGeWBpYuIHQ/PM2S4oKJt/aTUoV+HfaYjb/njs2Gjz84xD9oj
mRgDRA5EE1+i68WvONUgPyrJxBwx53eCv6U0lgw2B8uAZg5M4qGtO4wyLXFaSdf9Vk7I5REKcI2h
YJGqIhE8/zJKdF0f4Fv41BkuSCkgo4SVvT21TkH29FKywaCdmyiTnpAE7HtTKahbm11iuRPRYI9N
Ls9QZAB05JNXlNonsUVyDqZm/JUtWrw1SIH8TRl/p3mzvOO4rMMZTb8IqAadHBSuQTSBAH9nBMxq
4Uwt+ik5wtBFYInXdaoQoSCGrxqJyhDLIaCLmnaSAIdO1RGIHm+ycQ0iGlW4iQwMVBekxaArMl3Z
TdkNeqxB/qhqbzMD1c2ELfKQWTBRYHTRmSaFxgMaMYuPGuC6m48z9LnRUCGxDsF4r3dI6pDNvuyS
Q4Zftl4CajH2N2ie/dJhyjcbj7KXtyMYmxW1ywRJKy6cU4EtWVnxCWdPgOd1cSZGcucXrEudAe34
WRRKmO1AyMo+I8UuEMm0umsOFli+P7hA1QTUGpDcGmR7LwgURZ9OQRXbAZP3ESg3WcHM/3Dv//iO
SftJF3kBQCmyNQVSnjCLmstCi/Tv+Fnf0SEWDYAxWg22tE5gMPvJ74fpdkmYgauZysTa8BMdDKzi
ZOPbyGVq5gEKETJuHvp3E47pAn60yEapTMB3WfTywSVaJAYKo+gXd73g5WXpWnrNzOcKecgQDrWE
5F8P9Fjp5Tmp26usdroHPThrr8loLLsrDs1SUXr9Q4+jKC2TKdLf01Zhak9GWj3QQY3tBmHng1Yj
nPll+1aL4A/QgTyY8Km8kVVFQuI7Xt6zXZ9j0lXmnqejt98rGz4rA/h+8QG4qHLHR6hG8060O74x
jpU7ExqEGHu8Ftv5Dwqx/p4ZOS0iAaZA3XbtTJD5fPF+VVH7/0/4EptRkH5lJABm7yYIcw4lbew3
m1AwSZ/tjDdFMtstQCRbzHosxP5Fnz0UXjZig5SAk2V+7G0q9ZeHmk73HLb36FWAB3TF7bWd33+F
acpbSlXckBQnvLZQ2gleL7oBPh+sZ4Vk6bcw7L6nr9S9xGjaWd0CizxnOfuia7qNdl0xq2Ts9UJp
YXNfZNdzgqMSS4g8tBSHKd5fZwKw7mTdVtqh1l+cGFuAdrLcLb4EdYzdduHNpsqKoweIv9LHOepy
dafeXU657Q1ImDoGCsffcjURQQncIolm2i3c8Di4c30viXIP8dMb5r/cE+lF0AOp+u/acsVytRh7
6ibQXhKsKQVUX9WILXtk8y7b3DNeOL35itoYYf3BUESyU0VZMjSs+yOvOPHVJX1TEroqCeOsDjuk
YnFoR9EyO+tPCZsmcGzWENoQZK4mFmm6dAc8P4HpNvc/4SFb8vXZkv3zd0xQgzDWoI1IsyjGsF68
Q+6mP6oWnpP5W08p16sD52SQS3v6KdllfkQlSK0PIu/jlWzxSe5rE/8pDtvSvgz4JdR2PL1Jbzi7
pKVaQUkRGVI/NKRLqyBiOfs5Hm4DtIjKT5eHsXhmFKD1TBOckFo/MjdnpKW8zULc5IP+uQWKwBib
pymwMs3P7PBVXIQwnoEBOlNgCeCR1zWiLKkBZvydYAVdD1MNAtIAIyDbtX6AbHpDZgBIaD/EJ+Tu
6gqK9byki64zt1Pp2KL1c0Zfhr5fBU8jJpnwbOC0rgwUWG4fqwB2ClVR9gHlG4jhmvHu8lId20IB
vXV7j8q48cYIQanXT+lx29+j/p2JCXJ15tfuN5cyWdOYZjMiG78jzkVZtG3fCfeR9C1tcaPY8+W+
DHQB8KiUd1F9TMs0AuM3CVuRRpBagY7zrWF0GM4p/VDhjNJT1nSt3827bLze1cBt0X3U1nJk8RgU
3sbonjm8P4yZVEybQtW+72EIIx9bsNWFt23bj6e5YnOZ0PhGUOefp5fmtithXx+kWtmi1qb3opmA
D8L1zHAo6YC9HEHBEMekxDf88CtR4X+A19syI2WpDvXXqm+sGWX7wBqAOIxY3RH+HXRrB7FvRhfE
qWDQ/ZFUWdcjpos0RTIyeIezKFiqZZ2pa86zEW97Wpbp9xs9j8w811hDl/ACB1cfBZWRM8G1VgjV
5B9MBlwUE32efyueJm7ZT9ZfW+nOD0f/u0q2ZbNj7uGBWoxR4L84BIKDyxb/5QphBIPGvvlQgfcL
2TWJHZriGNVn+d720/Xfr+x9Pd0qqRDJN5xyuArUfe5Iz25zbTKm7R1g9qoTe+cqtKR/veJudf+1
K+sqee59L5dZQW6XCs9t4jVir1tBwgEllgHQAVHOHJQjM8qY77dLdHYzHJqeiYQ35hYfH8H/Xj3c
0SIqPIa5HIGrRFTdINkxhjLNNtEolTpvorGStBArsRUsF2N/2i+cHmSl55zs5CyYDrXJQU8AYRM1
QubqoSJIx06EQMIVTpv7OLk4zgMjNYpj76X/xOLUf/vuGCwy5+zDOW0KLnQE5ieJCN4vdCiiiDcb
XadK8niKX9bvzprhBlUkLojfu55EsPsXRiRGTA40cxL3qz9nnK440LgaIe6eiSZlH8CDnRg14ELI
YD30sJy8SxWLi5VOQH2e2SzC9Xp5cc3SKmzZSNiLSAgPPW11Lbd/vQmMg04OtIXKgWU1sAh7AuZx
YI4rY5nHdKMmTxacuyiGbW+uiNxCK0HhKP/MLvpGoiVQ/1FYE+ikmVsFtX1hWOurdMmUhgRYlz+1
ZxTU7s/X1Jl9HiZefAAX6dv8aQzPJvYL910U8U+8IJe+UbDqDnmoMZFuUX8Km6XI5SNC/XLuZ565
hX0+h3BO8gKLeEQ+mafzU8J1jDPc6uFC+Y6u+veIlQcYDnx4ImxadHluCmc0wVszdreaN0SaiE4x
9Oi9y74PWO68jf7jXkP18b52GtSARTdAKy6FK1RMlATHPH7/KDkiXl0VeTvIcRjzjaH0kMHi1rD7
XXeWguQ+qkV+HC7cOORHee/RligiAegas3xBlHmMZbjUdcVniR6nxst907sbMvd0g5WlUBqwC77C
0iffzihbn8uLiQRZ1+BR0cWpppgLfOjFFjKWdx0bcGbzuilz4uQTjqVJxHYUxuT5LKLRqcC3NSM+
PhOS+QeNY7YrgJYTRCBSPON7+oGZ7AoXp9WxKXQ+7+XQ7Do0k0kqWJr5aPHU8kKMg/fhnDNqW/GA
YOIR081WeAriDWoYTq89j0bigaoRBhPFcvRuRL++qc08Oa2RTU4OlyACxw8IIfBLMgpKISVFTzX+
PVtX0M75L8G1MsFgCAFNJuVRW756ddnLecp4h31eOYbpJGisVeF5wUYRZiUzz9sDnq/wOk+KGqoj
Gm5VHRQk2DN1XSqTAY4QK4Uw0Ms85f8z7dcXYDD5f5C53eIMZRw8CymUjVOXxP2f6L3M/1AXhMqB
8jBEHD7YrVvnUhMWiah2UCvJpwF/poYFi3P3t5t90RFRU9SsI4ngkxdQULjsDBEYGmlPL5CGWJSZ
Rr1YQ3M4oWHzHsbYrB9Kt3SPrvTmZQwAntgrEa27sTw0aXUy7hLO0xQX6MevnWZhNc8ji43CrZ1U
q12E6DJjU28ndl/1XOmT/TjsYqKErwAiB5if6rzU7SDV+JaUsDsp7fvI7MfBSxipcUWxB5URmZ3g
wIn/1Tq3SulmsL6ecWKkC/lWlpq5U0XUg825K83vtSVnE6/kvYj0Zfql4exq8+Yb3NCaAUy90rGp
hZYQg5lRH8RIYMXL7slXAEO0q9UCQpyk2Fi/eV6Cu2ntTuNuJE+lNsvgvk+B+LXPGzLz5LHhEaqd
ouZBZAJEh3Insel9DvwNucqnQw9WqKE0m5Hqj/Ze2bdU3eR1BHfD/A754sQV+kVevdAlN54JRc47
c6Vcfalgn3rKqomnS24gyDNP/leIHCljpp+5KRRhp0K0H25Ybkm0NUfjN0du16bG49lNxx9IyXal
TdQwE59R9TzZCk0Dv1LqV9tWybkaNdufYD58CKYUzFyvu2hUJdidokaTOVvZRm3mcumD/sWsS2KV
HdRGjp0+85vRyxU45CGIY9C9xOYqT3Uo97ly6UNI/QJkN7bUtvgj5Ks3ee910p21Gq/e6JtmQusr
VWNPaq0H2elAiYAPKwRXlonJbMsUo3TM3KPuBnsTyz+dSF7RAewcdjRnL2ITeJ84PMTqkGxNWs2Y
oz+oBHxFD67AnZuAO/o34uPWkw+B+UC/SHs8PR6+wtLwh3ARnfHOlQPyCkd1AxXDlpAr+NmZlXVm
9N0V+PogrKjf0BfQ2OCC5kqd7pUK7/xkRR5hsARUEzm+4ICW0LWW4707eRjctjwLPtkc4Unty8dw
oXo03jSSowgcmQAXSxAcjgO4f0PZIB8Vyf2h5eOUD6MfG3wKPDklQEN80sGJ/g5D43zGNxazVPCW
XrEGKBJaUaIF+FuL6Nd/b9CuQhilgq8lxb93I1cyss9Af8EPgms3SuZEWB007G252aDJfxXc+xc8
BoBT7zTOtfcvlO2pL62TUmtzwS60NpyoPR9Zd9flirSkjVXwiIIyiij/2l7gC8DW9FwEvaD+O/9w
TCfyfbRFrwbu7c5vmkE2uTFoMsM3FxzLsPxfiG1ef9dnxMys6Ik+0uz4FpdIFKyJlwrqxm+PtZgW
vs23gAafRYTqSQiL5CzORMtFGDYn3KndduswgKalklJ24zhmUmAar9ndMOJgl4xUnkSaA20k/DEC
+SsaahY985gps8YKMp3Ut8K+YGLSNAjM/ckZn7WhdtPmaDqa3ghzYLOE3j5E2+3im2zaO3QEzGUy
shJnNahzwVx+oqGVx9JVRbnowTdkfSV59ha6jp6TXfgmYx529bI+8MTtmshuQO3aeqqmvz76C/DZ
86hfDBt8oVLrOai3kk8F18vki6W+jVcldPJD06w49h1D9its2ZjKYQ8ltcYynSOA6dC6Mt/nbUXL
piXKHB60qe/6dvyXeOHin0YT2GwXcL6CdV2m3GDXhi7cDNh5jJPRjvxC3CMpgyC35i9NN0hE2WG3
gu7FNaYPsJn+GLVncHeFx+zYwJSd1JJGWBM+J/BJ5fXzqkvWYevtlcqmANrVIle/WJSGN3oSXzrx
i3b86r+DzVvjN0K7NviO2vnqu0unUpS8G0eUDISkfKcfVrDaE1MG2M5B0iaOB8brwRwNNE02P+ye
AtHsgr2bS5Z+niX5UjoC5XQV2Ty+M/1179sOUrz6f3A3yaE6Zl25NCxf6OQWqVpdfuUqz3zR3CeO
W98h2qrA0/C9Rum216qqFrJTTvrybtVxhqJd6Zs39QtfEPCopxrB6+R5ZMAoTA7eGKo95EV9kpoH
TLRq0Po8BHFplzYcHAjIxxe6L1bf/wh0CUnIOYrlivq+fI5YQugoPXvf4QsDdPfOu2Ll1Yuf15tO
KKaTtTxiuJNLLEu2D3F+p2uKkhlzrodsjiJHit4oIPaJg0zZsNyCcswmtKy2T/FJfuWbFqqm4HdY
e5Ys5k6bjcVx5kEg0n3JzgrrgA4Jlyg9a63aVThQxxwu+wi0YnR3K3ICbU7JiWjPUaA08jBpU9as
zw7Xvp01RaeIMflYVrrqpEYbf0ve1A5ugOTOGx5pJfd2rUoMEpLW/Q28oOPIAaLaNQxv/ZN23izM
oToGJqsXDhgeFbZBWMAoHb5zLgyUiJybX/1+khksL2JvWA9/hwX2X6QwGPWrP0aFoG1cpolvY2d0
hI+18mdhbpTpfTa0QWA+m5KcYKd2h8NUdzC0/BieTkSSW1DpgaqCGONUaz/xWGJNvCPZA2CrUSTV
bhs2rymR1LFmyqeJV9EdTqCCk5Jnr9tfyaarhiP7T/NzQVISTASpzXMjAm1uT3MnJWsSk4QySeoE
NRSByoH34QgbhmUk1JvDBqBRBIqy8OtqjnX7dg49Oqy/H26UHXJlIECOXWDwpveAxfBsM2JsrfO3
2laROksVJgc6c/xF7hA6xvfMu9mneTBCh71nhCaOcm/IRvcrs35ICXohu7AXb7gZvw+FV9ObK0Qk
5DnhXPVWSHt282I6zDRN2eoTufkLRLb8Wxs1u1Q0KX3lxNfRYEulCMgJbRoaA97oOBHVb23ur+Rd
Q0rkOIxCt/4gVz0NonOaZ1WbmHkZEdw6DPVxRCjVTqoXkxPDL7E8uA1f2IopxxG2wNGuDOUqg0w0
LMbll0G6404fdRMEF2h1U9NY/Uxx84Y3G2z527pBqyBRww2QWI/BSJmthoV8f7e/Rm7pefJtKx7U
GTcmemc9SoOpwgrDoQBoPFRzjpDiqoxe15V53AIYwrVLBUNwI6F60ftlto8Gd1xs4XRZZo+slxjt
k5oicKNKir+ROHTDFwRyoOf71OU7fPLHbZ8n5V9XGxQZBW9Rq3CW0pVy5lqo6LZkueH2XWi0WOnq
FlbUadyOGElmOrlO7vsSBuk50SYk0ndBkUl80you6hc8e5Zi1t3tR3jufbXf5RDDCbgzu72lDWzK
MpXZAaGMYfA/S+jI/217rhkIM84jiiSK9aAFuuFsZBy+DX4IHSDbh6MRD2u/1Y6bLfU82WPCGzEL
6GA7hm/RGkT38FXll1+UntYea3A2nvUk761f0s7KF3UH9hY/8WR4zeUasKN3rBm5/gHRQzpNNzVi
ApZJVXP52ZpwI1qMP6T8+2si3SrgChz5UGkY7sQ0hU5vH5isehu0aD/+CC+8bL9e4f1+YwQXEprx
jGvbxPGjpB2LwS88Y1T97H3R7ok+YG0OAbTV1oYEZvxAGbFkVLDZShiETkCfD1NPsXeNB7mcviR4
W1lBJFJ20wS2E4mWQ97oB9gh3SdzjtX0obDJ8u09Z79bX2K3tMf5r2AM2heKoKQK0lDt+gjMvY7l
sJwn+D7aluoPEeIaP4220AnWT2NzQ9jhaVEKEKmR+yQK5Vo/485Qo12sa6hw/EwJmDbwtVdsflA6
mXSaCx7VYWQyZj1zhR3B+vZg991K69fhVSQEQla6xUUxlP7eng+tM7CY/hPk6nXGblIfMcfW3Yee
BijZFqMaXb6hlDtmzDkxo4AOTPb02uj1WQLRXivfUwEKTj0HfQUMS+EPJCSoiSONG0+GhF2H9SSP
MpJswGi1xdo5KgTd4foRx3BZRZXxvxBL+BjUuGCxu/Ax1MMc3LELLMPv6kTElgojkNnCPAXz4PG0
kxcoi534yNfDxDAdMcd9QUMhZS8aKx7lVOqOm33czZI8MpWMXxCXIIDLvx3AoNsxVQA/EjVN6nEv
s0GBcukWAuTzhRUN57q54tBf0C+8dWo7EnWNgw30XHvB13IYZJy3koz8uI2K03glIKESUc0dcCNk
fbC2tsqFrAqHpXulTQ7rCOgHcvFzS60K9ysKbMzpOGDdH0bNvWhw4xCCaBl2sJn40iD7snuQOGYL
tbwQdrnx0Tr2L7qkESGAY/azDYugv2h8njaMW0pVhHGeDr+yoCcBSW4C0vQf035hEPYktks/AQaV
zL81sEuPv02h/MSzeQAhsmwbqazcHsYfu0T6GSudP43TOEMQpbsoFMrwRMmK8CJxDNa/sQTOHFrK
cpYJhtK5m3rDhMjIqvuEx7DB54C4oaHGY84vrEBrfrajSk1gM7NE3nMhM4+A1fBHMTePRvhwX/Dr
8zjp8cjZbHo7vCnQRZSX7LQhIYWo/KVZMmjLmfycRJMsueeTr8ADc9DpEeOVkwb3+O1VLiNvYpE7
D67tc26HJib8ScqIbJroekhI0UcHsOf1ycezkGUEH+HwpEW+EZ7ePVjYV4bjZ0OwoEkd05HllkLy
X0+vb3tnzMHxEPvvZ2pVHlaxroer4sjCkOWbs3bVyBxeca+KHKtDKVZsAkHc92UA2b55OqpWxrPV
k0gsyAjFxLXf/UN1wrbCiEFoSrHzYFArBPy8UNR0B7wlIir+m+HSdO4TneOQYaJ9IU1KOerNSEoV
iLhrgKvjOyS+xvseZ5kgqQWoGirFFjFOAtgenFRYgStlkkUfLxunGfxJTjzJ5VenvDwz7lnTg1aN
lsqZdOUxIlNxL7d2SEjlaRUHFGjRQeB0fzjv9uw5YRi5H2mafrWySi52aN+WEAZTQw/688Ka1Bvw
vOXy9tWRlMboXfRbX0hSPTAPe7IBoFLt7fxvWA7IfshrmcoeTvu/NLlQmSsSyIw8EdWoKeUcTgdO
VRVTt7vyYCXewVD0mbWoeajuP43wyHkMD8/2g9+sRjQbTVPBM7dg9cRL/DExQgZ3Bdo7ecv0MetV
YypNtWqShfF1PzZ2++VqZUfldtq4XlNfG4xTlTW7Ec1+rd3QBRwwwwc42ofccUIIBNDOBu3vtXCf
cwIYqnbwk44MTIRb2TKrEMvN6ZbOtrNCnr1ACAkz+iCgyhRgF01Pmm+vc483m10WdA4jPTSLrjyU
gWTparqW/7xAq64Kg+qZs6RFole2Raq75jNWSImteGAyQbrST8Jee2Rx4axUEiHuzkAYE3ppdwLS
oQY3mncq2yHAV4BWD/8cSCwb9T/8KTqPg5hq0T2Ee6nTQk7g6IzMqge0UahnsOR1O6+mjZCknScn
Uu+EW/DYJEEhrRLlA/THB712DCFQVcfnhzgaunh+FASEG48cRYb6aYmL8Ri6n4KksMh2wQsWcv4L
aF8stVMV6ccDUeecMVt9N4y8b3rAmElY+QD8F7cG+osbXts/fiQlWi3uRrRnv29F0w7IG7Tfj44Y
VkpIQWGWrSmWOzwSKpipqv6gJa01DPypCEj4fq71eOhETFCnsDzWN8kJ6n0vRd6WlO7gVtKcQb24
SR9J/J9SwIo8mFz5UTFLpnxGgEwuezGX334W2PyWdufNjgwL04mf1s60nwqDK463lTCBaZBYFw+R
996w1RM2imV1J3MMH7jxj56hmTzcxR5Gin2jg4zj02+G0lrEDOR4+rA2R26bvzmpISOW5ZEXHgjc
o5IJC/CX3lwJGkSUhCSZqhfSWTYhqpvJJ8E10ujsXSaGP817ztJ7p2ng/WrZy05Ed22QdVRQMfal
vkxCVPFBCvuYC+lsd4dxJPHvVYzUGeZ8P9VvQnSFYc2T/OHFgKTcZChdmO8EjvJI/p6urMvjpJez
WqtxbKsZSuHDwwpQHt/IapC9Xar37ZCUvksUdQSArOcrS785Xn/9b//Y+RiFhr79m5sRfzu8JocX
RceGJfvLXM4RHMUj/FsyrKddcO6+HDf8k2yB4n3wsHXcz+ECHkBObun2ZWxveXJAekYatkUO7H6b
6mQZhHeJwp8ceXykxLsaSyRNXW3iT67mUgw8UmTXUZNDOi1YivmdgzeMr3ZFzmzm5UX3eay26mo6
MBtNaPXw5D+WjYKLlMZBlsKgo+PjwPSDY26B2D43HIvfNWMmUT8Uj2RTwDIRyRwwEXOI2NqHAcMp
zKdCAPt2oZNM6DTnSRMJlLck/xe9Y/DxT0KjjPYMz4Uqfisk0/2nUKBqee2hIZ31kiRDhuN6BPJ9
xrdUWkUrpXMYL76r9D/RWiyf1NxbkkyJT0Bd0xe7tRf11PB/KmZF70RyhtdrX264nZKrFlwKeVyV
FVc41kxziDQH//7eVFI7A+JL09oW/Fj1qNxmJRElzJT0Gph3wIlqenPnazK4kb7NOgaC0s8RILG+
jW290zFsHfXeUiU2eWwI0FOWgZTiu00DhZ3LKsRAdoGK0zzVSau1dJAEJRD9rWB+zNHIHJModMlK
gNqFGOS2rBRvYrwqsO0tkJf+G6yrHP358I5hMDiGgTtmL4BRuHGyb5i+cDwuxbAeii48xqSR3bHB
Nl7qYyZU6LMAUvpHnApOMS35JI0nZg+IFHEhFEhlqzRGEzTh35vkhwUkpoeBXYZ8DnqCuPXAkIOV
Z4BVEyhDGsrpSa9O8zCYhvL5xSgX8spu1gtFkuI+f1pS0ftEjLqfRPE8luoXgKwbEUcANHEKB5j/
aQUE1BBCCnbRnQizAMqU3R4okRosg4RRNdCtVyW0GHFik0wU7M+jQ7r/5ZPIWnoyVg6eE3VXchOw
LejEQHxnipIYBAAEf0/sA8mIPDqfSR/NZgkD6TyNupoyHabO1wNz9dc5irQHoRu20mmUcUXFSGf7
ATuETkMcxYfcV5/S0N0HBn3P3vZiNumcr8y1zRUkZRgSovXQ+eDxtVKftq2JrMay8eHOiDNfrYud
+lPyBlzjz1A+ugqJdY65V+vd3+ykvTyK8hojikDK3iAQsg72wcz6mXtwOtYgSipMYPnD3F7T5/ww
JhqPiG9dmgzF4CFNRDcHDPvrkpwf6EApWPmGE2MZ/8PrwvH1GXE4YUGrp5+nt6hl2fDPWBQ5bKIT
7rzAAwutDCD94EHiYDrqw5jp9do6iFMHXkprat57M9aC69+7EHBvhzIwiRXnpdyrpEUosLGKruU4
vWoLZ3dj7LTHFkwrgPujPuNtsAHIeNvPbQ74keztnNO6cfX2LuBbILFxaEgdXCp1i0Sic5C9qTUe
hyDM68OTxZiVj8JkjLtlmMJ1jSeOb2nuSOGFYjcJYmzKaIwAzL+UbwGi49+iLsSzFbteQ/EJP06L
gSioTreA1hVWFseEheJXGcw4ZN0doXpFmk0Md2hPdZ9rRBysqPdZqNHtagpumkHqsT+j7yQnEWMQ
yajBB5uJkv0CgROCrLGc7UnhWyZMRPI46LgmP3e/CGQoE3MIqlRCCLri4tvjIt3JwY+6hb8AwIgX
wAbx8C6C4ocNCmS8Cca5iF9AGLvFny4QTcGGYbfOMM9/NEzcg5wugP6XyTOcMW/CI4f031N8j6C2
1O+aOjvM3hLxMbJ006bVSz3J1U5NsrSGBYyBojiDAfaEEQX8YSec9Tdx4wg8MTOWYqhPesVP8ReT
jG73bDiaE0dYRijLwiZUmMd8Hr8vyka9i0B8Y1mxpzxh/dxcOrcQRYfNmIVARZpmfpYq7/d0ISfl
oRRQYqN8CrJk11kwUQIL2rNQ1SHMhix9zUnyqDVS2/ar7zJggYIpYSfCReC+2+LLck7Ut2bIdjQ2
aI5cZCn5xBRsRTInQ8wdtqOAK0TSxHF66JrwCb3dCdRGJppx7xw29IgDluKgPo4xlyZ37VDWPcxQ
LVowYjP4/DKkUlj/uobzVtFXXK74sLAm0DLZlDYTUbzF1pCItyoOyNbimrJBDWIcpKyZd7Iw0/o3
/iU9c2e/ZCrrk9iErJ0SDODCJqn/hoVIest+iwi9O6a4aXbVtPbadWahQqfHOFMsXl7Y9mw74yj9
vb14ildlLArwMv9K8qqvW2Y3axkpO1AFDYwLU9PTNnREC8XBPQz8msX/F0haiuiYWtu7d1fiyrAA
XDkzVH5S/TvRnEjn0WtFVlR95MSuDBz9mRVtvuSeSlpl1urDP4FYJtdF00UXh23JxKwpgoO/FbHk
e83wvVSldElmNUMJO/Sihl/09kH0sC+siQdrpTsxAAAismmV2jYGQVFhe/f3L8/clUhR+iMh7eql
1DR9hmO9jhwq/o0p5T0nuER//wEE8la0vaW1rXnfiFU3bpr7sR/H1/3wBJggtBrCs1FKs0Yrt8dH
+laeq0+Gv5zcgV+hl0oenK/aVk1hyWMN0etUJEQ1wEJsus4muizR3+F8zZKIb1iNsIsyeEYgjrgq
t2jCODiQQOVTvm3Q5/zXc9EcGvbjAyAlcgevYYfShuPBCcoYI/rIRNLF9+9otTvEk2Bbp2ZDioUv
7yIqS0+BTHuNhN7SFXOsI6TChv8WOFw+uiqrceYOwwK892ebNdNqBcT71OfVt/X7Yy13gqe7P3BT
sKohDMX/mqnutJJ+Qdw4MFSvewmeoqjhnG/YadwDgLNeyoQGn7FcGNbEG2Xw585mXTpFzSBEA63T
u699OmR6i0QJSoja3R85/LxyrQWXySN5QzrL0ePRctpQTc6T+mvXTeghxYe2g+o5A8+YvsOukaf+
7DrHlbFDIYwchpcoOauF4wc01BHd8dw8DsVQyVJh/pd/LcJsVjPbHeN8Fm4WZe74Qf37Erusz7mg
cFRXIFEpvjqU3PMiwyAtu2SjdH6JdO3nyO1EOOxDt3iQjrEuCL+FGSAUw24cQu9aO2SvEOVp6W12
hFJMaQv3l7mIc3mYnRzmUCoXAuWx/t8Zqeh/w5Ig8ErD1I44tlCXaQOtomuMCtO5FAUTy5JRwN+J
BPp17tQHHJg7Xgrrsf1cRmxBxwPFU4NxZHPHaxiuAxsxQ9Sji9TP6TJGV6PB+Oo2KzCNIXiyMZAp
uF33CM/jAcBK5V7VmMzu48zI7ztZsWZOOv6OFEl9Vj/RpGGyGDBk0qhd8HIltFBSm+JDrKbg56Wj
o98lsqZhGQXWoHWWg5CNVmyXmtFcBun+Je2zO+XyWh+Xthp/Nng9Xpuro9lcO0KdxO19WJep4nKk
txVNu+YU/Z93SzUKh/uaZ1fVeQAmYRlS72w4oSUqnKIbaETO7zIOCHd32ruBvFM6alGgZhMIq7a0
+InNoti8QbD5BVZWGsUWBJ0b6RseLHT6ocCSoWQ2ntv66k6YvDO0mgXHeK6GcT8fe5whlFIdEv87
qhhn2K8k2bPjUoSNmZwLqUtQoMWKU2tLpgVOBQPFHSq/I4M1b+oMcoKA34iryPhrABU9QpO60Eir
udxVoJCMtJI/MeKghh0MpJ/lfIJv9rpk9KXl1GcozlHX9f4+2osK8oYM4dgXu0lsyUe58BnFjouK
VGf6PageN0/1S2zjc5pz/TLMxytvWJ8MgSkezkpp1EXPhaKZF0tSQ3HRLGwQJFlqv+mqogwG3A7x
x06+Orfv1I0mYR5qpDP4vw0ExRQeI34veE/RHiCZu1S3y+QBY5cTXbFwEUpc9Yztk9RFGMjfdQ4l
7AB6rsJ4HGAbZwYpR1syHQPvyA1TCT387zXmHGE24FpNIr97b+LbfJZ7PBTckQdFHWH1PKEdOOOq
orDLJfWKusBGVVuKvLJ/0CKNJ1+Pr7jmZ1fEAmWfvjyUC4VPpxLiNe53uE6wARY+PskJ/M4VyGT4
Y63/Nl49cv01YOyQDSJPB+zDuIuNK7q3/AAp8rhzF7b1VV54maUbbjcp8mb32cj3dNmjlj6OuMQK
djeHm0BYj1dPX49vupI+09hGoxe01DhORGzYszEscngV+zhPiZiXBxCx7+MThJhI8YRJttmH260V
ZIsGdBvvydUxBXst3SQCb1Y7iGS5JnWntfVtNFbuV5avfcebWEYmM3qhOHxfRqVsqjFKW4hnTloP
Ck+3ziYYGLhAQErs91kzuvonl1rKpixKtB5lzCRlkVqTtBsQnTbLheDHSp5MqGGXTYGg0Hj5G2fA
n7POppYyrIPpOl3GfO5DLGa9XStBmU8lszDxJgpiB68zQpzdlmOvfVj5QMAShh8Yk+ImFuYfFPm1
k0nEwlv1pHT9Myw38KD2s7cjx6jlE3dqk+S0EW8msU0CCSae2OnvmUu1NuDBIbKdlyKA3wdeG89E
wC3HkPtVRqOGNGEA8R5V6Sh9CiQ9HZb+ODQ6oqJhP0exQ4vp6q2JZpmjZ7ywQz8sa0tt+jTtCiow
t7MgO4eTw3Byh4uTKPqDNIe7XZXCWPer+jfKhdXYpwtSoY2c8YiekkLZw9yl3Et34gZJb2cnKSJ2
tE/SpW60tZHnUGDNOFPGSZfMN3K8J9z9CMNMX48KV/1uYpfIr7O5hwDaGsxaVUVvv980yIifionB
gqVHzWwlyK3EtQDa/h0m06KMdd0ilKt4qjDuvvBdcmPvCEJDlS/0PEQ/FUhLzWJMW5bLpXkCrxHU
LJf9DEB3B2G3hhZbTvDHIwbK5RZLcYfCwk7BztscYw5KbzZH2/V3r9NA7XviDeyHApW5qjO5ruge
ebtAaiqkGpRjqYcaSzuur7D8m/wRmWiWDqoUP7DuVTYGFaa/1OAM6jLdUgS3JFTMeQyoTdwpkWmt
73B0+qRJ3er9GAURib4ycIXExsryupHY09k2TTIBFjQyjcFNNAX1OnvjHNuGlIiKlRMMK8tCqT8e
/+yhvxX5bIH/MDL/29J/dHmYmxR8Hx1pmqcUPSm25Rez/3PxAiy8J9o9YAJSAH9OoRzSM7gjrxnF
NepnvSY9e1DbKuRltHk7msA9yS+tLqK5URW+BTCIjvz7zZrmM+bCCepNdmnIlnTkMUDEjhY31lkT
I2J0T7cgYl1OoVm03Y71pZ7GT0/KjFIWQrLdzrEnCbvnRRkCgFfngI+hZgZWnIponYgmDlB89WGW
7zv0RfEtsXEn5InlPPN/JpX8g+fQ3uhiVPZjb3ZJd6SzszaozR4UfqU38OYiPtUq6QObbvVfikU/
Z6kBtcGCgDZsdIW5yZLSoNBfpPOeTWZUPatjEOYONsl/h2jCeK0t1WDlqNXydZAc43NlEM58RJqn
8A9dM/++nWVcSs40ONh2rMljRN/NYvYjnhcTuw0uBrKRl7LRpV0T9vmYzmFXCBFOMtWrCcfXR00h
EH0BcJQ3K9ifr9oKxY4qIeV5NQNB1rkH52J3F2yzFq3ju2GawG4LCT2pweAqPTs77EF1zWGzJzij
Fv3P353+543F1njkRu0459gAdOp6H7mOU4mvFKvtbnjYkjUdMDR5i16/sxhSjn0V3W4kR/YJj5Gq
ZUY7Hyjy9eyZ8HqYrYOCpRRv86+gLvLH27Y789OFFafWnTvXFJbHahuw8D9uYuWC/cGJf2Zw1kdt
TjWT+4bibPy2Qki8mz9iArlPwJoD8A73UdmLyNvVQWN0LaWo0oS7m0W5IGwEoY4te9TeuqZc4JQS
Pt3DeIYU1r0eo+FzDNDUsJZSkElee/gNSbZPOaKmGSxj2t+5duXjQCvls02MndW1cbTSLMMuNKRc
rKeBnuOeTceGZAtSzUVpVFbMLDk0S7xOYcBnLzzjKNqYcUyCnM9xyMePzdZfCzmcT/OPlS6m7htW
p982d/tCBcsG/T+5oGufRJH8jrAK7dZAUCLJ5FOJveKrzMD2z/BaERE8C/eID7w7ZMkqWWpdSuQR
l9Z7RxJUQMbMLiYCZqRPQCK5d3GXwfxEbcSzvOjzynjTijepR5Un/lOhzeZ+hdSt2yzooQE5vFwP
SrEdWhvbwqs1v4MtCLcZU39/OfG1jmU6ChU/hU6PxOWmsXFrgn27wAo8svWEQFYX7r5OxioL4KHb
NTdtOX/d2+Im7ldsYi0Pakq3hAmc6s+vFTolnAPWnFMgm/FQZs7Ss47KFChT8SMls51IjFMe1Eqw
VrUnNA62KpVHruvh+qrjVdUKfi5g11Zr11G1VcT3TTHFPyITMjE6BFpwQkRLrjeIJipKB44qXxa5
m4kAk5yxDaO9menOKIQ1bkS5Pf8OAgdRoQZX+UL6qoavkeIrae1SgtPmQIEp7hVk8n4BpsA693YT
NysknH3vFr01k5mHhVD1OD6awc75883A9w2SO+kE9FRAfmA4lkxSQvzHYELYHWz/dAVtGg2YLV3h
GAp846Dx6+tsn0RXG+sti2RnMJuRW4KnEuUPPCBY3BjueZrxEBDwEYpSPq+TncQ2qKOvLZJwIF1D
jpRC45kCCXu0cOBLE8Y/zSUSjK1ktXwQrWzzyeN9/ZBw096oj9mxOnSBW2ic0Tfwe1BSCXHC9+tf
sOpkdElc4FWKzqrWw8GYCYLcgMQ6zlLTIRWym/Vt7qxBRIe+PLa8R3dcVc+JG2atqy1UqNJZTheQ
ykSJXs++XX+0EcK+jwCaAG7IYC4m7cbEN8mkqPR8DBOzXCFO+t4+B1JSPShiTs+ZZMOI7zSMH+3l
sdoAWY+q9eqbAc1fNOvlCiz3KP9zZTCqN6y8IHD2ledAkSg7F0NL6d7KYsae7ysPl3B4+MelAaVF
nuh2wyFL5tjWug0aRzKWFsknGTTDNhFDCGmOQfA6p1AdII9wFSEXola1tPfscxqZWJ3qTdOXwUJ3
yEMpNKrDPkCa/k+WDAx9gXt5+qIM2Lnf9VrdLvtakcV2TAnf7vOXedaJcpTSZ+7k2kl2qUlIa7fQ
qUFblRrxUr/MuOjtfirmaI1Z+HzKUNLd9sEM5/oxkM5BBdkIus8LE0FAZ91ToeOt/PPlaL3oWz38
jIalNSrws35QfZJ6GgfJaRC2r30W/NkekKNxJYs+w2sLnL/CaILdkMsKn4Bkvshp0UuvRUrcKYed
2gR+FFysmx32IeQAHEMLWpUrnHxha6V+h3yezA+uKgZX+U49IlYUKNOmW/XP5AN6L5IAeAsUqPxZ
F2fAfgJUiktYSXchy5I48mWujNuIJk4YarrcaakctzEN3bfsg0/fwo374X1RFmQ3JoC1zNi+wDBj
uS5jS8YP6ggZCL3eoMCoWWsUTbBoqFUM9W34QrHdaCmqwLiwnw+2sZzvB9DUA/cuvGFBTMFmcoya
p36xhv0+Gtu4U16LHF8KNM2wWJv6H9UoPfnu6KuB1wLtcqIW3s7nOpMJ6kF5O3+ndFU/KDspzvtJ
548LWy1w9rGLSaMuAuGuclwEcLbv7/rT+GoZmrHbzwXUh3I4DcoMzVeCcZ7E3Rr4x1LfdcaRMvBk
E1WXdNkkC2CwNkSrVhnrt6VJjGq63MeKW186nQ6qvkCvCa4PCs3gRPW+1Y1w3tTsfII+ISSh7iIt
iH6MD3pVLAGKttgwbfMibxHq4i+pCCfH+mjfThddTSN+u6aBVFrvGIAr4tYazc/wIHrivVltOlWM
zUwdmyz3UgUb/yDjR4SF5dKsh+34SS7D7rmGWgPTMQoXQQDttx/E0KjUX/5Qq2TIBZSVLIcb4i03
RSTEJoAeaZGn/FrzBhM91G5QlNa5/inYdnvb2V76KHchH7h7QcQ2R+ElCFW9AFgWWuwfeWb7iw2/
oc01WzNtmSjrxYnh1hgMZrYJjfCxhxKWhbMA7UPWPqu9m3ulGsm0uSsngKrAUUmn0sOoyQm5P9NK
UlbdMkFqRCvFHvntM7xUCEW90JpteLumYHiPDyLmblVlO5+9figvcQaf4BWorfOQyZa8+WLkj6LW
tcKkqHATRYif/TZK3hfa1Of2sohclMpdCG/vM4BQkbDREz6+3rB/gWq62zkhzavbgWtzOCRYbG0x
6uPFjaOB6vmsOX+oCeerBV/mkskr1g+qO2OEHcIbKQekx7bLuAf8r8rIHM0E1xSyLH9JnHVVpRWo
+fGnr9Xjce4c3uOSN/wQJvrrKE51MqdKSjpHjthJpFw/apyMjzt2wjn8PX6cokfxqa840U3QdZ6d
FteqPUCsLUHFjGXVKkAG8bLGUn/ag1ZT1WuR/OpRsmiG0kF04bjy/IgGr8kqFaD05SbWpq5ktg0V
u93B9z6IY+i3h6cf2eGDzx7iqxiG4UKRakqXtDqxSnJ18A5yEuCRb8CFrXvbq3Jc1CsalqOFIvBa
jtjggogxQwOkkcA4O2N1cB5GeNWojdH81yZMbKIwDIrE9Bg8m0zBWdt0RkcoMf0dlB4cc5+uMjRn
xlbrX90KvHotWwCbWnBNLhmRpluZ7bFT8mv83vbWlPpcsYrP4tCbEOTZf6yyuTmdDP3jfIYzrAXu
V97/0QVjRVBAiJc67moJYJhTOMbS20GvNIChaKHI/MxhNOb7CGkOn8fz30uggp1wXuChOi4MccJH
4/wITn9iBLzI7PNKVYu7WhbnZFqHoRzNiAbnANJNpGeQfyikQeSpZ31EngwsGdnv87ZVczmTPhtK
JnsKFDq0+Nhjhpi58Jqx1OwKxe0zKIv3SMf5N68kdd210//SFZp18LuWPMbxXyN37oDgS/+/ECFX
NuinJ5d4IB4qXC8GR7Mrh3dSDDOZLlAaFx8zhkKbv6DDIC/ftfDMWN8tWRGYxW7CFFm28PNFXdeb
g7NNPPNxBrUxDPdUoetcnVzyk1Fj6T3AsCPmpczH6kOWliufNYUWopcfqhyHqAa9MwRToRPVCkrm
REVrO00gEaLYGhGxOVqKGViMJ518BFejwSIAWmRzzavKUB6+nh/kxpL0+J5uBlug+mUwm31F6WY3
8WAgBA5QmydXs84RfhybBom8T9zZpKCb+t7sqJQPXnxchV1LcrQsVQQELg25TuqDRjF2gSVpqHdx
PFQAfOt8mbuBXnfUkQhqG/WfTvvuylFqYStJHOxiWn56pIQTHI9CHDfH1K+OT4fmbgFEQb7fufQS
TOz0q2nMdqXqksE2vouuPZ7vAYM7F0DEtmTESV+rzt4so5vB7Ol6ozZ8sRMqAomrku1l7NWD8WdD
4tCAuZGViLlMCcz/kp4HrBvOzjZNZY2fRBJmkLAVNsLGA+dPzQ5Gz3w+83EAa/tBVZyopMLxhA1v
t5rhftTDmjf8hFMMtbrELPXfM0XJqnSSzAX8RRyPF1zsxII1y+jCoZsVtUSgrEOiuFa+71+88hzS
d4ttRW2GzJ2M0u8P2pHKWOt7t8y9zLoBwK84ROkQRCXG4gBeyfs9I8puy9vzk+QQdeQ37nUKBzp9
IbNjyEbM44Hnjjn92XAJp0IHARcIBFi7hUt/iW1BVZVJp4X7D3JINQvCuAi7gHdOmh3WymAMPIwk
nn6V69yBFIK6bjtxDkZ6c6VQI9xrlKtSDxnL6vKGLguC/kDZ80uA7koMfjXSk0f+2m0WvwMsRLYY
l3ieU3wBDAtVoNovYzapBAfX3JhcQb4D2FqBU54huHRi/XfrvDnkQw6kTn9eiBY+IS9ES/5UaIk2
Bk3U+hJeJxjHGC+SJ+ylWxr4i1UzKYtXQfYgkCwqgJtkNgEu8iZLLD+waRIGATiXHnGPqkqNrXT7
+KCfeKzwvhaIbIyvX7bDDrmSUrsObjzrnfB+L97yJr788br0qeiETgW+Ap6egLnwXQtXzWhtDDJL
lsuO/3om6qLI0pJIEJbU7CJL6TuNPqBdic7Atq7Cs3tbYbKw7lOr2Gi2OtGZUEvK0e9isS6alW6M
523VrL2OKPxC5w9fYAhhw4pdn2VkJZ3Al0mPlJEyo5kG6pHwE7rXgdYNrEWh+mNpV3Cyp/wiavDS
8qvT9VFtQlRbQlbFh/ej/RpLivnRkuyBsccUbZ8SG/WVUMwaCARZZwXoXPm6EfJGrX14Ok2jXqrZ
7BCpwYG6mc45RVSQBYlw2VNZlHHcAF7I2Fu8qwyo6sXsYrvKXqwXiDQWk9uuK8LzLboGnTdeqZMy
apInXE61Z72JcCytsP+c6Q0jajEM3+uwBE+UyKazLfqVidARrR8c4r0fKz9FporH4hahs54AFlPf
7+ptim37Eod8i4FXne0hTTo+cUW0USGyj1lNaZVnQMSUmlnxzC6ztGM5/2wxtVsf+64niFY+/q/B
DO1gx/DEttAxv+rl3osuDZKvHh66o1hDHfL2KMdoVq1moPnYsJG3rz4lkFYeaph8tUKx/vAHSxwO
zt6U0tBAO8egVv1+2eEOhCfekA9B7HdqW86qDK8BOM532ladHmHS8+QWrtFZ2q8nTUGZf7jG9oOp
qjVFmWhfOXSDjOgCP3wYcSauCEpNvWkxdH1VhS+3bsxovJk3JplwAMr7ezsN9e2v6SL8R74+oljb
hAyj3inW2a9sQQ161xibBOytbaqp2AsSL6DAiFpO1/faAa8wR1oh7sn2YqwN6b63QNbpgeD2mV1I
uRFDeOwC3z6m3DyR6vU72mjf01AaHojPdd8gmDrkpJYvmKgcYC+zegbzYftHEigMc4Iu6cfzK4eo
S2awlPsH7NusWvituEDk3eoJ42csIEEqt+hE1LnpaSPWcKMnIy9FqCDvquxyi0RPZGkxyTtEpRln
EugIFGnx408vEm7qKmXjZH8m5pl4qH5jTbcSnCCiuAqdTyuu1pBFwD2ixl78mxXfPSVwk0YWYtwG
Q2gOfI41XvPvKMx1XXfTdJoFXR3/rCwC8TDnk1Ge9rSzdlgxdbgAYRcqyrGLeu+a+Hb78NjSFpop
ZsSzBy5SxzxuSA5IOn1WF+PZ9DlgrMWO0QnB4/4du6GrT7T1Q+TPXsPXyn+XSxbQauWquPiAVXbg
Vfa16EXHVT3eJoIDc3yGP0okgt/km1sdIDlMe47cgFhVmur3IG9g4sLlyedy/f5rOV0GW+v7eO95
2jCRwfEBBtvhvZS+jPhTuU6CvV8OGtghEU+7yzKoCVgaaGrl6CXZ3vFWU9adrcrHaJ3yuiGRcUWW
KchjDSXsdMNZJnwhZR2Lifi3qgJxL12rr+tpvylrC2GdnGaNav/2AkZV3ggiKrqb5FkYulbKvX98
3TBklJRRfMebrRRACDVZwnAW3SFugVbsnqx4PhweHQ6VrSZaCMADNjWBApaHv8TsuTSb9JmJABOq
zTwV5U10Jr6tXUdc3QYoJ4ku7K9B+pPu+o4MtUmHm1CgFm3YqHTusn3A4q+3sIJ13syDAwmLh5iC
ADCz7Jfp8kMI0N4ZL5v5Pui3C1l3KW1RTGmn2ziLmcA6+kX6enRa9+SBU35DzxxwF5YsXqxobWkT
CaFt3Pzg3s/iqCwwT8kutIXzTtv7j2/HJIrc6on60Mjcqu4a+zUJD89V2u4w9O9erraxXSfD19qR
0WlgpR43qeKee1wkWSMZem9miT0WeqgO66CCcZlwR1tE6kf/KAqRZaD11zz1HG6B6B/rsGmRmWYI
tGIui358JXtK5IhdgNxuU1YLtBQMlbZ7WQTE9kKBB2OtciAHrw7T6uuhpFoKdojFeloDhS+JIqFj
5oDKls0ugiAwhHEKOEZ39r2wfeDmQsDiHeQS7q44dZR9V8b7P4E10eBUFJkM/dHU+n924LRQAtRZ
BqXKRYScSbvsYGZrl4PRshPBLCP7s1eXzys0NWoBUIjx4DjWNGKYaIIZbQf0YKJXhw9+TF4YZZmL
1dETvcSvt5Dnwecq1aed4IUWUeLMenyNjPDfcfNz6psw9rLaVX6pPF4HAzu8KJ3X+NeFP+C+NgAM
uqYI/R/MiMok3mMOYem57oO8bBOY+OkRRNzT9vXT/NsDfIqpLbWAPoYU6rdvVIq9Ud/RHFkz1j4I
Hd+hL4fKdzNYdH0xCgcpKDKC2wAI6nnL/jMG96vNjO3I2NxpBQJM2FhYnhT0h42Dec6M/TTLjtx1
we4CYssyQf2AyjKE/uS9RbT2aYG4WY9BV7RVExIAslYbfzgDNGdTGalImFiguQUoZF+yiAd7aeUC
qV+WjLk3G3GE/nc6GufLjbJ/8Yd8xPe2H4LwvHS+78kgpBIORAF8Sohz0fuFKbr3l5L868CWpwnt
XZ7LtulD+QNPHG2nr4D8jZ5SwDUkTy/FSg2mlqsqQzlUEoVR0oRv6bcfcEwzmtyYqI6fCOXIygzQ
PAiS2B68jcQT+p78xtomHy3zU3CUBpwZIS0M+JKJdCp3fVQmeuJdQ/8fFQc/Riw9sOSEelrn8aiA
Re1KsmGcnYZdDU867XP4Tz8gmY2aFTxS/E29TdFppxe75qK41vR+vBX+9525diw7I/Q/Flh9G/bc
cihwOKTjZzN4Vu/cmc8gfrNpm92pvVfDXAbNYGSrk1IChrJMQ3cOS96Uvz9fhnpEIrJBlDLNLRzb
pBldHWmXdzkejpxRkhH5vwUIXRPBDkOvTqqq8Y9uEZuK8RoQ2eLkD8gKXFffpEb1HF0RV+W0UdX7
DYkufYGxjOB1pRZdWSC/kuw1Vq24iqrKFfKeQSIcjVAAhWXs5KOtTTlLoTj9i4l/qVxmP1FsugRG
tDL21rVQAZTni0R3crjZLRmaETmKMpFw7UxzyCGlgWPGZoPcmj6huNMOcbkgrkYtVNduYoVTHNaL
Bt6O+rslyL57kVSD+GV6uRtlZLvAvzr8OurdVumIUUHoWBPy/uURxPYWPGW9qXCcEU9xoaMhpBar
Afnly6oxHqbBqkSRUfsm7m07qi2ZMyPoG7kPZZUFuVhZ+LPksnxTWxNAUv2amcxD7cJDZ/8FNBs2
S9G8w5k8IwhoUmXN1o7dT7R4ewI2M6ehvujO0yuNAnE6aXU6WdXuG8dlNcOV6FdzCtNLC3OVQEwj
hJYnHTC27hD8mJVfh+16T7N2e1PqprRFF0iqFdCzQTe4CzSwcCXGf+Tv9SDp5cYUOGwjil3k6MZM
uVM1zGQS7ZiqYTAV3XcIucJV+NfyCGZhQbQ8gBM7NjiHgKUJFK1uy1IyAS+/HgZx0O6bjIV9qBCh
Qi7wCDYrVhHruhbVzY4LEvesLgrIiB7p/LdNyMGDXnr//spW3iVtWaAH9D/PCZONDBVnXRiP30Qq
+oj/YFZsB9afca+rjOZX+3LsRPUl4k4SpL8XQXF4Hm13ankPF9P7Ev/QrALtUBxSwhmueksXYZeI
/vP1I/VNkRr4H9N7QrKrZhuCAnSI9XSQXqJqWW0sqhHEFJNF65c6uMumbL6rKqbXYsY7RRCrS+4f
+h+cT1ErAWeHCkYYFX8AqzOihgfUyz+G6Dbg2ia6oljoBCbteGJins2s6QnzC18CI8Pc99v6wxJS
1Ue6bWJPXEY6a56uBTqnQKPuPAKANAbIhgjkaPcSxtpHsiPZJX8IFRlaZ2CTbBZnEebWvJfFgab1
RMjbvRvtu6i5Z9oHKf+XekCilGRTt8B97v0CIT0HJio8z90gXXrbhd+4FsIHKiH/d4Vqc65T7btw
hqqN3k1ssJKjPLQcewcjh3Ev6v/bSUpOKJypjINi08WgHwm0sdsZ/WryKHzPmvA8M1pDB72GaBsF
oXIrW9/6HIHhOQjdb9DFynFeF4swkgKiohVDeORiKENnK7u7oSkCMtrneoDmhRa2Gl6ZRJiHSNjk
0lbyAJ+dRTzpf3dPV0QZQn5iVhCUeALyVCKCOnAX47lLuTfFfXaH1uNHarVWOYjDXCGKk9gjvd5H
Fl8W0t+JXubub7pleMyuToGd6sVjoqCgfCprBS62e7hyKckPGPFqX5/RFZnKCBSiVibv7wphzeyQ
sQUrdNtUiUECUP7GNilwsgfSM9o3bkOTDzJzPOt6Y9O1DFMaaYAtOjitOpymcON/oExoogUW5P5a
eLWEpqr4aQNcNgrsAK772Ue1rl68hvAVAomIiDGfFWjJIBCQCFtrXsvVR/NFFat1I/TlL0Oxv8y4
l1ik4A+c6i1lKIuhCkBw9OVXbLDTPCLc9fQ/uMWyofqXlwaIPchR1qQW8JsEtdvcVO4E6j8kQl0i
HyQH+8ae7of/c4Y1ps90biWRI3lz/ZCIyoCwHdCEYXmGWhonsmVu04R3k140zNuxoByteEu+hszA
e7OSYm5EpZP5meXDqtO5JqtK6dZAY39za5kQ0SrqJ0hb6Mvv5clxvAf/Dapp7q6HTcUIOhldsipZ
FmYArw/rHIn4YXNsCrL2HdCzGf2/BwQ4tgfpR8rDyg3P9MKhF3bhG+y9ugUbF45YlRFVWMFyFu77
S/CXWgJLOKFzhqbZ4Hmf0NZyIkzQiWRcXHxhAtDmhubPiZXelGLgdznC1BwuJn0xM3P9qE55cqFp
4TGweis5ajokt2vHV0paimlThqwol542jGKVEFxzij8hS3iYnvWUJoPQgfe0WNbBYmeEeaok/B1q
L+UAcQbYLPqcccFJcaIj/y640CD2MTBiXicPab82u+L5/cQm25+/iJzIQPENlq6auW/7Dr+PFs9u
EOjNTVnl3XNMi/KPlDB2f0OdRzaUTo6PNEOZoUe5qASLqf0enXt/ESJ2xiVGkIz/nC1s1mXjdTCt
QH9wIuPh+sY6l7Qc1rMCgo2PI+Kt+QoNsU54Y0rI3CgJPVybs5H3vvHCsEVqQDVcsdsOS88aQ+Rj
Wal15LsncJNiDhEArD6YHuKfFo4KWhiAjR+s+zPVsrEciIzAYGxD+EVa5qkaOjzVHVs9AnhThR0j
z7CjXk1Wx0V2Ar/yvEplu5tphIcsn7IFe6CdCz5Rd9OVLbmd7B7Z33JH++RiMsBhlKG+eHw9KkoE
DfBv3QPsoNsicK1p6sqQnP18UjT1xROFVjiIyLAYKONMRyFXHLp6D8+Sh1E6nz6kS+B+MK1/uJ/M
awzRdv8/crSc+sHn1t7JUZzOf7WkJddgHrGv8ov/5RJGu41sDeGQeep5Vy1AVypq90iWnloiShZd
V57GSrbvWnY9MyYdvBnoQBTy3fkpvmzQ6/xfXtsmUdZ3RY14yETHA4eSFiPzFMMNvJnlae2tGWma
eYfkBhWwqVe7ojDptW1uzeSUHkRnkAK+qUxBzcjF8ZQax6Yz+WxsNL8hemvMFAk1wrSs0M0kU+9/
9G9bu03FsyakGHG7DFOErnUF2Q/yJRJduCbpLumpylS05fBtn7iw31Mk7/ZaSP5H89o7vCvPvxzB
eUwJu4OJwBu1FuLGidFXAB+MyLokCCiq//ULygfhxD7zRB0C0BFIKjPVZIAtYuRSYEhXy8fSR8Zp
xV0p8I8ofnw0+wzH6GjYXpGuu911JbbA6T+Bji0nTwfhxbTeAY2i97tqDfVwaAPTesiRVgZaoEW8
4CPxplSU/LcMGIKaFm0QG7jl4OiCBaeagNJwZg7g0Cxp+Wk0V2bIYZLqyRnDYnNoicYlskFWelaO
dM8hYX+1ELt4aUErZ2+epbgTjTjf4/zcWDL7/79qwMceniHFgwmTNti46+p5Wy5rCv7gZRiwZZv5
TyiaUsFXypR8DDgnVGv2RqzjUb+QhCGIYnMU0BLX3pfW4X1uRQas9r6BfUu+1S7P1ZpI0ssYx71v
nA+fTU1c94gB8NwDnEcnEw956pMxmoFDnTh3n5Qcn2XtW9/N86HvRXLWWhzP8axVRykf+oJpQ94S
KNpA4zpOogzSg1inyvnXs7qyg7KFFGXeG2aQCXCJ+mxSFPn3B0Yj3M0+v3lj124yodKdEcF/9z0n
svNTXkMewgbsFcVI49wQ/3d5zqvqzj9POno4XHCRQtQA0ScpD4pBDuOdr9VpSZSleBcnNW7/75NY
GWu0r8roID1EPGn8q6UeSvzwzO5l4lBU3LfvRMChIa7Ih0ByYCfMPUi+ZldL9yocQqOmWPJm+yP5
wSNh+xZOK1drh+I1G69NIZqQ0XMjmiiI9Qc2Xq68aGHiBTaUZhnJt6ynr8eZboJxDmNZYfQVCTLJ
4/OngRJ7nZXxQ7XUtphM+3bS0ebLnOwYKkNmCCuXgMUh1zUAMKaco3xznz76zvFcd9AS/XZzQxZL
AuEq0bdF2QBn2/zU/daf8VTsH1cArA2zLj7FFIDVLo2p2F6x5vI3iBEn4yyhYbPdbUl2AYlfXnXQ
SqXD2n9jFVPxGZnFQqttX8DmyDGnt4DEuHJKnNJkExZK18fxUZtS751osq1xvDF7nZoI05wOmHF4
EF8EeTwunpS2pO8ri0TYvDl1qv9up/co/7zN2PdeVnJthR/QFnuuxFzshLXojWZejAubN7qt7Lid
nOufGd8lWE8RHJzY8Hu4BpcJJ3GvUbCNiGCgRE2LLwFJfKDRYGigTTHcyxQqmMZq0kq3J/cegNFh
ifvIUvfi/F7pia+Ug3O5+BMH6NUXVjaZdaIEqT7TZB/aoOQ0m8WvuJ2pRote+zhx9W4bNt4t9uV0
YjUdiWL/qlnANM9/ts0UX25OwMh217ByiZcNwcoaFt5HZXhK60ykUDmeRWyPOxjj4uEAU3qTN15n
4Ji14besQHYA4zMv1I7lEveKfBJ4GqwvgmY2wG/yPY7CLO6qAiKmUlQM06Xj98C0r+cpN1Z/FH8e
YWqwHMZnH0GKV+eJhnoZ9/rBkhvRzCw2iv5JHW4W+pj6EaIh9YVNcF15TdLcY1WrAnvQh7bKOxms
e7jqgwTShaSwir8S5LpO+WeWtEunrXmUvxAkFX9AWMUUeKKPAFkKkFBzfaCHmEnzZlOrD7bVYhp+
qESXpy3mNZNAfrA/oN8lTxNk2PNmJ/oUsm7FNwLzjKEXV1RR3MIsL36I4ib2zYXkk6y8ZVGDCFFo
YN96jjQToe050Eow/VUa9N3gxOZvw22oQ0t7Q8Oeibm7janjLzcL/DltO5kPAqPgd39Ia94wZvsr
rIbHlBGRVr5rwV7CHtT07MxPNSFo79gfE6bt6e5tqXzTWvigJ6lCEjYlnD6G9XGxQjg2SdY+nCbA
FUxHOf86TYE9z4B1RV5+LCZLgb324RVZf2HPqHqM0B2Q1vbbWWfcH8XqcIXatTs0VDKBXCJ7AXZx
6TJJ6qwxth0+P1DyRPYN8sVuiGplf1T6Qiqyrz6aS4k7AdxQmnF3XEKvGSqHgKyAfbqqJnkQdxEJ
GXZDXCxfkv8ecdP9LmPhnU4qrwILfpRct5sY2mnzUWtRVpm4MBERKxovevdMTKI6j1V29wY7Nu0Z
0Q+/REwzHHThRZkHcieUuuTbyaeY7O6bOG281ra2tbDYTdjXnGJvMFAQ+1eW/i7zsH42hIAU7OGv
QN3pv/+GIfw5Hvw7eOK+HWspIyvC7um83e2J5YYiz663kzqe41vx+aumSMzevfxKs8QNb6oNtVua
PmX5IbU110rjU/i1qaSigo18xRNnrE3vCSonB5JFNkrHvkBPesx8ssEpRSDho14Ib8S8T2Mjk/UF
KVv7S+z/rzgR7WTh3aHxM8QPPUIabEv7feeoMCENJgmJdbiHNEhF767rvj5iMNWMgeM18tlzlxlI
g5ToSagzwSPxB9rnk4LRlXxlXGGrVMxHNkqMWexpBgiLWsI5gaeAZppXUaAc0zmp7rp4qCAQl76/
AwckCRunp04FF3k/iSGz8sZOD+cZdrwnUB2hKZEMzsGF1MCNz4SeMCbwf7NHzLx2XLVxqx1L2lnt
4+YovvMdlrFU7neyv/O3+4vhuoAYWk9+S/U5D3d6+0/VkFDerQy5nCUfZGyCC67j825sm4K8h6+T
CXlseP7n9na6Y6VXuS5RwWiIB6AJtbqzkORx9Set6kpFmKtJwG68y5Y0xbghhxTb5b3F7jA8D0Sv
MtMRQCyOSc8NVGanzwQDt7yf0+wQxsFNcbDTEursTWFRnCFjHPs5k2O7Do4TeCoSbg7TpP7m0omD
X+Tcwvle4od337XdOHJimn29/b/g5u/gWrxY/5ENfNdipARI1SbOKAQWoUnlwOakXtSBGoRTC2xs
W7bdhwmTcmLPYcaVyaRin5G8YrhV9WZWC+tuQWAsWdVlmZ3NJw3UJ+/HbpXwRJJr729QRknVwJNR
7dWMoBucS5RK+9prIIg/nO/BF9iG9rj1+cWbLKFHjPNs9+AK3W707v48rQJBhUAuC8xi9W9C1E+u
+vnqEnQ8p143kzgiEXB36p3WbZS2yLSqTArjx51+JftTnTmXYhFpQSSE1yIbCag2+SMZqQ7pvkYC
PjDGkj2BGLkVOGO8RCzT3zDARRCodbifvfKNEKki0nPCFVeBkhgdFiyhYsN5oDnKXLS76T5y0Tx9
Z2s56S8vOqZ1RpuwLjR6eShUHNSiCrUONJGZePrCAoegkY+dqtGoC1Bf8WlBJn2H0sE0KyCEX0UL
KXFePlOofvk/IvqYsCt2VdVo2+iXFP8CGeBaquZ7jraizCwR2THhB2rTLMxduvZFV2VNEbmnyIL6
Uu/mBAbJqdqqBtpp9M3QmZmtZ5kvjbfr1fflv8YomItITT0bgtLtfLLEE3RVWF++Gd2eJEN0Odex
UwNawnyB5UqSLVZhih9QY/Nv0eEtux3gqpp9LJq5RRAaUZgai8JYSqOc9uQ/N4aqPED1BPo5PSjt
dLm2fxm0UxLrLeneOGbecPHtimo+vRUe4lXD2jrSH+/IC5JbUZ8BToPpRItSwAz+/evvNWPnNcLG
xM7uTzBGJun5snOPuzRHuge7s9wVzmqMEBB4mvERTKF4qOEsJNAHUoIgQyjZX2Q0li+p+FfnCK84
DJWsWImxhAKnLAGp3Nx4fLNU2Jk7tL6K1QM9or1BbekGe5GzlqZuoTI2j52kAcRDB+5r0n0UOl/I
nEJkMaRfKdrpW4+CHQRgmqiHN8+PUfsB6tA8PcbjowHnySF8Ny5cyoxCLVq0LD9GBQ2RvrhkAeSY
Sz5tU8yDbhXIJvVw8swg3lVt1Em6ZAUmrwHp0kJ9W1bUsHfBKcORHYvDTmYoKqljIMZITqxlvbtQ
l8ZRvTKGjeOgNeQUgeU9BWRuV+q9l5DmkrjUnGLDkbx7fiNN/0AL4GNNvp5dVwQcQ/1itkRhMaJ8
QgaP/fCiwo8wx+/gHsb2sngwNNs+oUyxgzok+M8QuoI3QA+Kzfjaw2NcbaxYrkuYrfaiwtgfa+vB
9Udi7rSAyRBhT3zjVIHngwOYP/+94Ud4hsRdKidiMZOPfsUg6rSuqeBVTZTKCKz2oIA1L7i1Re0Z
6KbVnz7qRCFwD+pvdg9Uk3fgNVMsgt+pnr34Q5jBzlJFQsMIdoIbhI71q5fqjVRg+u5Ck0PWeUEW
GgDrAMI6d31z627AQexAsDvzWQb3vo5Lag7E/iNIGnN1/IEP1QCSfICoqZMw33QttpCH9CcYTwU7
6YPJufehDkTPd/5Slzhau/7QYPmRwW4ujUHADaCyQplBzXqB2PeB0d4dQw8O7YhoaJQRpEtd1Y56
VpkFC1uS74unZ5F27aMBYK1tE0iu2XZ+esze6lKOoL+6H/11OFAmp0muO3XtLZaokKERB9rii/uw
ywZBVOyNMlfG4YyU32bT7lOzCpQq5HYaYUXk1fIa15falvPJdur2cYvtWCgibY8e2gpMAYw3IU8b
y2B63ju1LIK9TbLD/0P/SC+2Fcog2r/44BhHuqB6t6YEtNg3qW0gww1pq54r6Y3HpIhXaijoIqNx
mVfLElWfvuM//n2yusGm5Xy3CefZMLKCt8kHTFPNtGs+35FEinGO8ZwEV44fjGCvA6RB0qCWUQfB
RtVDx36IPfhtP5v6k96pRSezjonaPRJnFZCntLf665CjN4gpwoKd24AgS+KxME3XXoN6/rUp/9nm
lFH941HDT0tS8pPzs+Q7IYH14xliRf9yEj1hbR13LLKBXXc6fPquKp+BxU4V7ZfULHkGsQBj4XEl
ytpvS3UwQPml8QTXSVFwTIPK0xJS6wiZjm9Z0u8bV8KlGiTh4BhqXDPQF8XRyF/YosmxwLGj6prP
H7+78FYPFYjigfhKUsO6grVq+PvSUjjaCZV7scuCzYqI3t3HLELLPg2YFZt08XoA/xr68hjMxZtp
5k0H1dDrJB44YQrv/d83yoP9aX73bJmvKuMInutnXqzS3QGVdS2UL9lmHdyUDTJ/I++isuSLGsKA
AlePZXmQiwi/+ObrbwzXcRoXcHqHZv51NqYjC8NuQOGWXmENOQurYtLP/6kNGGztIOxFQr/Nt0eG
dlaLl/HyFVU5UM2paZn9X6k0ETYcGohzy8qUPRBujASnj8Z8M7GDrL8TIEQBRV6kWaNtWtu3jybV
EEH7iTXEQiAgy+4kyNa4PDMT+PzR7zQrHnqsXOfcwPuvLGOJaBh5E+Z1wXv3AzLZbl4Se0gSMcsr
LUnGCeimnfjgwvrxxON4bjwKCwN/MY96aPojHrdZU7B7Imx6++TGwYfaU1byVMlkzbl/2c7KrGGC
Pywx6OkUTwBQPy8JGR24zl86JCUXGN/SHb6oyDraoehIKyE6DkwunbQedWp1p8X7+8yJAgrIV8Cc
ti9htBZ/v9ho+ZpOWFmRz25Xg9L2WuMbW+tc15CTwyk+rsqPn/oEgPybr4Ng8CM7wvasGBcQZnIQ
X+l2YqaQXiJVndI/dzB3cqUE0+St7MwbHwBs8uuPOVm9ywYPGNZa9DFJf1zFA1l2Cq1cZy9cEgA6
WgqFUBt9cHth5RKy7BqtbWoMNsBXjP9HqNfJp9T+KsAErgs3ORtsTy2GgrkCiie2ktd4S1QAyoP9
/YhdBmbQ5ea0xk3Xt6ghfMXCIOFxA+2E7rKsGFUSQqQvJaGAPvhK81tvFM2uTqz9reOMQH+wo2Y8
kPpdWBfGVb4l0cx/T/FVAdLxZw4X3G5SGBjqm9Js4MF7bsjhjlFKGhLPPxOP3jxrnQhqmIISeRmg
1cmtHm8X2sbPd1l20jFSLNSFgXohgOVJc5OiTBfTs078fKF5uX0RqnHDDbo5d5nMyrP9bWijwj+0
99Hy+/9xks+293SUlLVJDA7JttnNbjl8jHqK0j+45xbBzRAJwy9VpjXd+0ixunyMS/D3af43R9G+
8DB9pg3sMyPBJPRCv12Q+uTOycN8IHIbM8gODws0pCpEdMc+8TY1VwYbqXzlJSrd24hxUh7wK1e5
oX9bU0zBC8QWGIreFgi2lgfT6mt46bOctjTCAiiJ8cAswxTmw2niRaKIKUrsRG14fDGjy9VuXZRT
E6Ae6AjvkZDIz50sV4qDXV5sTG6SmUn/1IOKu+j/0SLhh6ofCtv2Gt1DXGKswXzZtzoiEvyaDV+Y
sfLvo1Bjl+VFgk75QTf0qfYGxnK0IvYlgMwu7fHL6KeyPv3dDOzJMi+sGPYqTQn1ZO004WwlWu2U
mfTR3+rCyuqKEPOaDXBCCNeYkXWJzP2XlsBrum8jUFQvjlmJhGFJ6unFED8JWfeKUB24Y0yuPk2N
Jb5YWnUdKaDU6U/pwxlUzQVfRhNveMtkL5/Iuzm3Biit4LyG+5faaDIWY+wB+ynWEiPzS0dZCbqW
QZv8SZq3xexvfU+8k1Bj1A+CSO+2hSF7z6NYY/C2ok1y0w4LtrPS+9kG6V5ProkupZUS8hcGuJ1r
nfCA6sos3Px2zzhOIajWOK6ZAVjkyjIq1Q2st9T1ag/FucoRjuxOeLAwWOciS9oBl1XblSgF69gN
GNvy6MoZ1bocCREp385qQe3bJbQRYuLQ2ybLetOTq1ewm4UngGS0SPwqkOWaXxhUU2K4UUqy/5RN
ZeUdxiUUJUNb/DdwbyjBb6OUUiD4IAcrQAB1xWJQCrsBiy/8G5gLQ8vuyOnMw0unpjHrNMtfE6O1
ZaR39ZXeDZiZU9Df0fdbja11kgNuyOyKsr4n1+czZDX6qdVtRFqZp4wcgG6tKM3xQaDO+4AOdAp/
m1BEmB4VqgFqi5q8wJXhZjRfjcjDuSNdBak2u8BEQWc946zACVsg7OxnIQm8RQ93fXDhjG+iRLhJ
yHRArrGFPjbtBB6AGt+jRLZm2AhdV9omo7Rm2WQBm+13OlbbzmIybK0Fb9vV+p9oCSVDlA5WoPRC
VCzD61CDxAtnQoeMDVmVlpe/TDnZlFrU3d9n8+/4nOnPdp501IZFfKVVAMaqA7SjIV10n1GWZFfG
0h9pcYgu/Vtg67kG/RR3YocklN1cnSY80m5gZM/D8GzkIN4DT+zeI3n/G+PP5uSnd+waY4znoujq
UqsASfuRg4ROLFAlOF+GQ5XG8wXRZqrO6DCWORczedvJ1QmGqMUoeCcu8PRh5aW1IorFureWIDB/
PDoGnWwSPlKo4Oooi25gLdsxxQVIDpcrwXgUtxa5Cyc0Ri8CnHqjhXZRV73ACRd9P5h2quqsERZZ
TvgL9MAEH5qxyhAKs52TnLWUyisepuoUz5WslvwO0aGyhFR+BAGQynh4hy9W2+mRE/HwsoNa2EcE
rHqjhxcZ74wQiGsxSY9fr2bilQQAPnE/v7J2PpiTXrUtdSoOdvKY8vLCPAMz9LxgAuh42XD7K2ut
fyFDmqNqIQBMulEelF5JUR9CpVtzZ2CisPVPUGuuPjt72kSeLMXA3OkqS09jGLsNv8nEWJrMe9nA
WsQ4i+bR5WhI8duhz8L5ZrrxdnZbo8dytFgz/80ulogMu1O+M/Rb1eXQ0czUlZ+5fwkvsxFcvfgV
o2BNYrcnThiWcbnlEcrWp/jVLhDPXlTn1Pgtqz3gocqkq2ScMjoW8W3Fcbmr1olhKeMPHi2Ue415
H+rRbUKFajNAbJHkhStwLnTts14+q0li0V4H19AHX54yrIPTifvc8CEpmtGO1EHtgkNhM3ltf46i
gP0LedDBkngklc5wr5BSEXH1sqknKq1SA50BYyR7QgAp1MgkmZatzbZLECwzVdvoIkKVIOvR6IMC
oTRhJUzoQe8aFuTvaq+x2qqfuCZj/U+ekaboENv94o7HW5wdMYq58MbLY5lXTeC8f725zunWl80+
Zlp3HLMAnbLZO4LHO7alCssewYk0PEpkG/07MItue5COl66Zlvs97ueOwkPi1jJjgdaObXKN4D5O
MJLOIaHcHL0iGEz2vNTXO8Kf3ZpaeW74m6p+ISEvydjQCuvB5IxU/rO7bvTBOQSEYP1c1o0IzI0d
s+Hd9D57HzmWL3UOzrpKQrkf17zMbIkHD3xvREVbMTh7C8YXkbEjPzzivRcBYJO1kORR8+IO2eBs
JvRc6Yt40RgIpJr95gp8yuW/TiLuQxUYkGVrsqRF2Ls2sYc0pM0ujbb9zWlpQn2EcmUVJHTPqnnd
PO+70hUyzDF9LtjJYJH44wZxVfaEUc1qai64J6ihFY36z5Wsn0hj/fV7i/3EOT1YV5rn0U+RZtp3
H7rLZ0fZHRznTmpFrJhCYQX0oY5n/6ez8aMFNfvzvuz6Gp7GtyTwmMXNLxQ/xz9Z0FiyliZ173Q1
kRZ/xAePwfwZrUakL8WkHn2pMJ/dP9yRR6jU7WhlhQBc87P6psEDoGHamk0hjVCGJDmPRpajkakp
KVD+OW2H+FNa1M+Lm2OaRO5J2tyG0l2vspgzJiEFHE1vVDBEiZCcKcMhIHEJ6KUcL9BpSJBJ5OYl
6M4pPvW63a5vPybefrGZ4rZgfyoD0AoExyXjCzIBt2AS+Wo63zwHHMFY40rVpPfNl/9GQX6DhtaH
QS7SIyqchqtCxFtX2QQcvOquIaqhJBHqL9cXUnLfcTI7Vco/jhp+p+ayvJQp/oraqm5hDYUTzWTd
/aXN8P4VScEuZb56NJwP5ySbmKfpF4mXCs1Q5h/hZ8yKVrT7K7AcL8iYjvkUvvtvGOIsD3CZmUBr
X70JJ2F1WozmSQSWfiLSxeynsu/o7dMs4LfumSCxmyoNXvJDYbrFGiBFDoDQp0f66g2gztIZ4oK1
/wb6t47TmxdEqbCX4eJ5maNoFaW4nRoe8AW2P3UluL2361ejISj0mgExeAIWmKRI+QCR4kzLyUYf
EgVwh4aq2RYe27pwC/WddKDQPyq0O2K2WxVBhqHxWOAshz2pfI2+Lodrrz0j+Ev7A5KTpWjzcwpw
tkf9iHtECdiwQzUFe5wVKKSXoGlCODePUFEzsVxFB+VD03MnBu51arm4J7wdiUoPrler484ZT5JL
LGMsgyEPZY/eX59TRbCOmojKnByX2PJ352jR8Y1QienCxI+z92BWRoD+GeKGYiYbtFdwkN1pu21g
OcK0Mme8yoDkEyYk0Knwsx34fS56Bdx8G59mupVuewePXnj4fdEeOUsE12buqYiWzTg2bRfBrC78
rS/+IMXw24DJx7j3JAiFEFSm4IJfqthq4fowkkA5Kd4tubVo0b5cJObE4LrCvFyqnpb+YjmWYc9c
juJAA73DGGU3o+RGDtBo0z2PaN2TUP4aXzkrpNTv6nsgbCk1Sfu6n5nN+kvYyDf7JH3mCFRTjlsO
5L/k4Opa1Cw1WxkgrQ3oGb6vH/IeupLbvBO+eMvQXryUdPqFVW765LSfP8tfhQZEt77IWP/ynjxQ
J8tm26GgRyS9MmEcj/kvp5VjmWis31fdwzWoljL0ZoRXDjr6ca0vMeVoT8wgHnMT/PpdebC4gN3k
dA52i0Vj/KcMF2yVM649BZyakQBhd86l/pkBVfjeg65xMxfrtn16KoGGrWn1gMhrXsBW4ltfk0W8
tzUWpH5fmvU4Zf/G723pxn+3G38TEQu66Spz4PZzzQZg9u2Nnd0uPUl9VvHy0HWA0gOOQwF4tRuA
M4djJphLFg0uz4un9Am6M2ixNVvhystJH9zAZ8wAZ4oSAuQqVeFdOwSLjdaX3w/VMQGUQH3zLFag
NLSTfK7Zin78wgAnnS31QoTc5nQYjTtrpzygBKevEWSvfD2Lwe7kSqWUa/lvoAjKRv4pzyyjQciy
0a4kGnrEyjWc8p6eUFy+Y+d7pEPwvXvZMqg1SzVJftZu3xRuDyedIEbokj6rGZq6UX9kmRHib3CK
2dG0yB8Et/1eqbMN8kcWIEfSTMWuTZ8MB+koVi/285LyI81eq/cUnmvbupfzC+D0wpxZ1mVsJnYd
Gv3KG5wU+/mrKhQp4pKfE2GwuC05dZ8qXj2ZpdnKXsj2B3/8GSYhnb5W6hZgTtqycqrMNT2Bj2Wd
Ef1jdZWr7Nw7HdIc40sc+hQcEaqIH3a5R0vQ4dy3jf6T8cm8KNK3CLjUnBFWcONF5oU346RUcOh+
JDtMKC+DLc04gLT0QkEB5dCnvsBVwyQr0GpqoPzHq9+y7Vt8OoMTz+rFNRxBPhQ+ckCv47dQK8M6
x3JlEMyg+PhKrimVYDLqZvbXqBa6dn9uwtW9yjeV21ywuPS/pmm+5T2fnF0YVVXq4lXQYO6aGMUs
zeTah/5VCAsQsyx+oemTDPdSAvYdeDZmWgvVFWGAnx79TL2pOGp3vMUOgmZn5nadVPkV3glTkMA3
BCS2y6KHc83OqRmI/JSvC4dFdqTwtM3BvxdZBpg0k2mR3BNyY6XWEjfr3tETvh3CNEfM1m6DTRnN
HXQqK5RnQqUryD8Emb0Ta1YZnt5qyQlI1gSpi7ZVQUWKGF1zgaYiEsatrunchAc9Rpj/GAEDgHYf
NOMTIZIt27q2AH8RrKMDVk3cRf2uu7VH0BG/XhHQFIXuFn6hoyf9OSqONiiJ7VhN+IEf5c3lMrvY
M5hlUkfxOl+wf9I1dOv5eiiytPHIlsHo88ZFwW+VtzNf27COW8MgnQga463ZNd4sVnVBIgwOXLR7
WUMK9YM6NiA5ZmU/xiH+hsU0TgGXmVWD4yyktBqScnQXLQ/xQhO2XGUv+v/JpYS/8wVSuplAA3s4
3qMitvrH3j23pd9txCW7PzetcqYn6WyOHoSLs7F0o7C3qVOZxg5Nqe0mDOz9d7YvCrH9Q6idxWcc
zp1z0wqrHlVGBS7BuaK43ii8qP3NNSZlDzJ9xeufn2c7TS9eu1fklQkXk1vasnPbL/0CnQaSYR/b
f3FFiXXi0xVW4I42guTyOZ+SHU9Cti8pQp/vzo2eheN7j07a7um+d9u3OTYYIIuIAW9p6K0Em+zk
mAPAwEH1YwVt7KQeeWFnhVYi2ZBEuk1act7nOGgOMm7I2rxLp0EKLDtCR6yWXz8oYj0sogp3hh4g
0tyHIDKXSIBotkuRc2R6Kv62JjFyVnUo9LZxw0beIt49gdqeNwyUtsoQtXa7DCIjtzbLZDRYzhDQ
MUzDTPpYSuaTe4PxZVn5AKdHBOcANNz+FYKNt141IPLG9/BtkcMb1oSTYGa80J4fTdnyQJbgYsTy
/iZDAtFPnDUc+5RUfi/SXOEdQdc9lpiL0k8+Qoj0ZdVbGaOpCjh1qBpaGryivbYgOz/msB+QCNQc
xlAvS1I8AHs0c6bgN0mU1EAn9Z0lszrIhG4fm++DJtQ/rjCq2UNQ1s+3mXnoRgyyO2GKcUaTmAnR
FPUhhI1THv154/mBpxRX4fwt8UPDsJ3XZnt4FHkk41sXV4/ppzulSJd0Nr+ZLOeYUIuho+serxJ6
xFO/WYC8eYJ6LnUGBQqqfb1MxqCQvolWpdY7HcEr5wG/nspCSAIowZCGCQZvt62xjOOun6jyl4w3
AVUiXSgcZ/btbDGgUFoorZtqYt/wUYBmel1C87dB9+xm12O7Vf3cPnKvrnBzkMIuMIEZmiDCzvyF
2pCucD+U+gq0+ZrAmN8K2wJoRtr253H7AWPomJZ/XFvdfyExgYrMxncugbTVl5joNKMXov1hCbL3
4e6KXAclcLAKvPKln+fq4dESsAr5d3i0XI5wk3bNBfK1NHoDag95Xy1jSCMwNapLsLAuYG/1FQYX
R0BobXvYJEhSpLDjRcTgZ/o/lQ8Tv4252e+7bLBPyuTvxGTn3YCvyobP+RQc110dYKQ8MHTHZOqD
PKfe4++26wVIlXGppZ6/GCKfZV4sj5Y/RtK+jFAWay86/WMG7h/4vioW4WorckGap0UHBTLIi/Xj
NzuNkjXIBWFg3V0GnUFlygTlu1xDVqiesOSkGhCLYZjttUhCw35+OF00CTk9cryXYQ1jaIyJMcgH
+dE99W+jgZCU1pKSGUsuIYVApg7DTjZhkxBggxCthCljq6hC/G6TR/y+IdkX+Qvpdu1WRKUMAAxN
WJhBSa5AR3Sbb0blBrEvtj0aXDN2ok5O5p+UiuIL1/s70ZekTjv1SsWULw8PgXYVSctQUko9wKtx
WUCc0Exin5tE5wycwar6Ae87OKWYeNjUOZQiKxhA+IcXsbe21qhHlvLGX/+1X5DOTi0Mk8f0Lu1p
AJch/gumv4uucsbbDaSTav1LZgT0fuoveipX3/nmT1IJhbKu+yJSRHbcG6V5xkCdyWg1RFHvMsAC
cQtm0I8EDSKFuK0hD0oe+DkEh8sQ7nItB7C9UQRrlSVjrH9+pguLozf8fOykoOqPz5tYSCH3WAxn
eEuPI/BQymt3mvYGJgOimB9QAVv/ebA1lAvj1r3RM/j0+zJsZfW3sP/zImsor1WafwtHMqwLmSD7
eeFV6WYdot/3K61DkTlnhM5EHxRAwP5s4rn0Pxxp1dPG1sJUhXczUCeatS9YkMkFWDHaWjivPn7i
I8PiN7EBx9pDVuIMyOR2V6rEwwMfaXbNUV66bqft+wec3e7P5ZPpfozXmD6cNTw5+gljrjbqUQDV
KQfFp4vpc6mEUiDJ1GW+IGhYCS1DnjkaqVASDb6gbPpcTqETiflTi+HbLoTEnP4jZok8oJo14w6i
bpjoTBukexwjUuHqQlmm3UgaCUFvq+KJVNiObiW8ORDdIHnpQfc55403f0cr6YiT7asBULFMp9lw
OiBga9BmkH/gP1GEug3N39RVBpMCSQpfkegpSF+o4dy9iK6ss6s0XJNbJHtSt/9AFQknv0eJlOrk
AocmFuMKyQcn/sQr0N9tjGpADireKVh25s8rWBjW+/zdSuR3HtNO0b8JgPbO4w0drTuAIBlnBLZd
S8nW54AoJHMqkYZ0GV0ps/xdYPYK5BLH/HewHr5c4a7wauqdN0c2JGXngZWTCOo0EJNbfOOWogaP
jtOooziVnBcqaCJpFRapbONJmieSza+DtU+LAesbASP+Z1zTbCkX+9Me2cJtn5NtoplnrJLucKXe
8bA+RF5WFQkrsj4z9Kmo/1zWxmgJTKOMw3lFvmmmWOWlrYul4mx4mrjdGgrG6DVC71O6YbTIAR5x
BUtsHo8S0Js71hnrYSwAoILMYrr5XZT+HySFEs75EzrDwZADYaNfSL9y4V5ESZTl0RDOnm7Qfwsa
3XnOKzsFAT7dfexTDRP9iHohdK6ep3SXSFo85gSEgtYJn5OZAtT3HLNzu/ruaqDHdZu6YTu4KSRE
qZy4erMaRpBPIvRFMVcKsOm+11vCU5YEY4VkqcqhFwOAo+TMr8ZPVNzf6GvaaDNO1eewwKkwlJiK
Vn8FmafbumiYoJwuqk+ogyFEoT7MvbMhEH919EBH8zDs6gixcqwE4ZWa17Wk74YbN2nOjJc0OBCF
U4gS8tYaw0wm6fVPkSA05CHnivc7EOqxhlck4jUhu15EAi5lubsaJABcMpS6Fth3JpLjnlrtfmpW
YLHtnKOBAaM/RJgE3w5V0aTOgQuinzebRVOvzk8wA7WF1kFdHMmPTYxxiWoATEgHXbWlfRgloRf0
Wkco5c1+2aHJt/93OF1klCr39QtVCqtqnNzisjbQ3sF6blbiaazmtx7aYxDRl269Je1gvlsAdhUg
V1lpEMhJVHGVZTVjnDYsGA+CXhUkGh/+A26jhvXF1Se7RrH5seCQVWIo84n0gi0fQty0tOMlJ+he
sdZAaMoo1IEyxX+CBTRPEhUjvpHf44c6np+uNq2Z473cDNX1I837a96KumjJo4Cfwd0KhsQn/rup
26VKlT7XiXJuQMZ1XkgMuZ2CyufVXBKDi21UuHGgPPDjr6uqGZ18K2/O+VFRN7XzdyzYEQO3ceV3
k5vQ/5Au5UOTqQjS81Y6RdLkOxvuH9V/fKXOJVD5go8Aj8lApn9qbWMZajkp1uDJjurkLQNzzejJ
1+nPLMvDc/JQRAe7PxwbhsKx9CfNa+lV0WypfWV5e0/19tP4hnnMMWc72CoJ/rqXT9RDXmKYxvoc
q6ATU/r5nxiw+rRuO1FrcuLRwoomwuhRP9hfuTUzxYvRbfW/MEbh6MDRCnhgfJoL0JvMtPesAep+
Jr2jX7vlckqb7v0zxEReLGH8KAygsqZVn3AZO1FKJC30GeFieSZ7cU3Dg3PApCt6gxGmLTRDiJN6
9ATi8epYsx65+4ZYjKEJgfwww5rs6vpca4f4TqPQLG11+UmmeJpHOCi4IMu4AQt8aCvZ8R+nC+wo
OVRcO6b2CL5qcUWnz32ZnmkHsY7KogXOdv+UVPgdDXmCfNlFjLs+PwAA+KbR/g9Whg6Je+5ewEJx
GE4LeUs5j0SjDieSKWzpmlQR1IgEHnhqKwl6PkhJ1EBE0nbxXlIITyM8600U3kEvwtdMoGQje/NG
1PANiMcFMU0WCDHNJcOeAtV7MSAFp+tlKYuk+9r0huIMltMiZQcxJjqacZv/MZDBTuDkEQ/cLdS+
93QuAfc0cQViYGMBSxa/S+tutY3L7QYTOwsCnkJrPZZ92vHZnshDDBHJi2frFtV9uDtpEhXZOoWF
P0/lKKU0MIfZsEyH79VPzNYAx6OgZIBpOgqIfpBo0LQCOtxfi5epaZDL1ENK7wBHFFlNMzym1Ywd
B10d4+Fcl6ZK1Rkox7cHFuGYEwk9/pAbow9nMirfjY+UZeEgC+lgg5IeBuhJAqOHkYqpInOOIKWa
3gHeHN6Pbp1D4lVzjXMngqd4M1b2YTpaSv42jjCoD+red+YtNQU1ijCLc5jwvAyufDA+tsU1/hr3
s2z3kwjiInSDyx8ic8hKeWygabiLbdWkfLuJ0Mz4ENFedEqFI7t1TyxI+6lDBSsvRQKU5l+9NlgD
NkxdFNxv9ogc0COV7VaM9gxRPAq28KaWil84AvFFDt4BY55b1j3XbedLbxfUilx9uREIKj+loZEw
iL4YNew2AzPFUgueaCri+gJpzNO8/5h1QEFyrsLJpjG4Ri0Q8ktmt2EjDgzm9Psa0woh0DgaCOS6
gRFWb/OuxVuPaqQM7zU28yIM87d7HlC3SR52FozMIh5R7OMLbb5aWfztq9bvpfTiC3R6s5FxOrPI
R9j6/sqCaWdMJut/fuebRpy7Cdg5FS+Jk9MC/IHBi8Fs5v9DfdYlm7D3ZlOWOrUkMjVWcoHWwKEx
bmIL0WIOXCXVbzaYm7OmRp/Vob3ZVFllLT9kIXK9hIeyckenlGhw3zEfJTq47Tf2zHtCYm2rBjcJ
kgFCY+dO28uBCCqfWB/IZcJu8rSEao3Fl9jZs1rUDbxhPxUj/VsielPr1kMb9dPa/M95IlNOrVUu
YhEQFzcOSfKhZb7H9C3lgtA=
`pragma protect end_protected
