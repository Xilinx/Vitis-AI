`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cpmLTnckjJLm/GJhnEEySb5724
XCmSymMTLlXyajuUkv+nefl4yXy9x2yAhXfBlAkKJiYo+BnqQEh1UNkLqYAA87d8AoAB9ihUb8s1
IgM+IoyPR9o3uY+NiwUbJmA8+WWguyhwiuI5cBoSnntNWESoTGk94tPn9TbimmCK7vJ2fB8ppcY0
dzN/XzQx6rnja2k1n9Vpi5cSISAq+208kK6K/eOIeE3s7kpYpnZ1FcABWMhBsWlFy9vQNq77DLCH
vQTzMzjR/wZj9RgsgR/pU3rvXtLtkUDA/6PI75l7BHrpLlMLOGYsw3Ktut7NFvI+x5JYjOeOGqV5
smH45YmdH0hwITy8hhhfGqqpqrcOkgCpZZHdVao6VBq0JodHgH3TFuTTtNcGEJqjghDhfKi8nSJ+
DxV8rwcd6nt2TRHcGDjN3Zka3xp341UWVdbb/8IqG81tO/O5Mh8W7tr93Srf5UcWIQoUd7PC1jGq
kzeCcYrLrzP0GE6GGb6zwAPxblmbJxgGkn94olzg8jjVpoD8EbKZVZd3iX9lrKFUMnbiiFggWJag
EXfGV8b4TYwWVdU2vJ+pM/ur2cup+yPJaOwCXJ+kL4Oq1vCbYOtA8qBM1dHqaFEh3rmLikKLQIaD
kWZgLr2a39uIWlU4OOdcTa02pgBCaC74fGK7YwfJ/vI4asGigLzcfNzvxLlMiJRNOOk+tFtYLZIT
4/ESdPsTzaF6Rx30e/cI4zSBjYuCokkE/o1p/P2PH3k6jbSYWMB59dWoVoxvpgMfzopAP74d8YrI
1Zwtbl4d9qNDXgvzv+g6gf/xHw2zor8//Y2/fxBd2wSotcLnLvIkfXsDcpjUyFZG7AKo60VXLRTa
ydjNe2mpv7TZAnwWAwAwZbtdJraDfgEOyL6QwGbtrG4Mefab7r+1GXr1HV/dpgm/lSIu+mkIM0Uk
HuNGXwrymHqZIAFqNsziBtNQrIBAs8ZeX2ZfYdytR7xdZlYmGkmfUz/FMLrUEl/Ht/r79RDLef0h
Kko0e+4vftuj0i2uyTlQNptp/I36nVWPwFWE8ZPPSSVqX0A0xLaO+wlNsAp1jkNqsh38pMgFT5YH
Ev4egx9b/XaWWqE6jua816/eKpUuNWTvBMSWIX0qjjbQL33q9VaaaYqPjVYrPgSiH/sU1sZ2KNFB
8A3RBX/WjjAwh6eURLAThkdwQxP1OJavSrM3qq1Bz7Vs4k9vNMBy229HgbMTCIplK7rLBvrMhTfo
36EmbF9PDWjifGH/MePlmerfQzXA/RV3FurjBzQ/gEkFKjpeezOzP/Nz+5yxzymo4nAswyZiHIww
8YvZ0SPQlSgmDIFwYHFMuvUGhe+emfBcoCKZqJ93nVZNJdmhjfa8DrD+mqb5tj63QUi4mElBtRWf
ujnCY02nVyH8Ri+ofHNDLoTMNJXySN5cbiJdQIfBtVYbtNL/kSEpQ12EwPZ7gpidwgXgDJ7Mfkvu
Svw3uaKNPzilSuSaDI29OzmvBv0ShFucmEwnSZE+FAveE5Klh2JghV+264C6ocTK19r7h62pAWt5
PmspLP2S73EieCgd84RsFSF1jVKAZSXGPgononltS/uvX1OKhW62raQcYsFXa8ufksxsy3vwRCq5
Fr/eOUTcIpdwlTtE7AepwKsk0eDxh5ETb8aa7dejfFKSxRnPRl10txKfkbZKAwYZysUdOAVLzd0b
jjYm5bwIouCwK29I/1LCLKcOv1zgB4NVtshAJW/Qhbe48joB5BQnhQM1PQ8VNbm65cjSDTNZHYEJ
bohASbTAiVaDJV6Fuki53WxTusxfQh7/necS3ZEH0fJl9YuEtlxGJLF/6HbnwL0xId/hW5zluH1i
e+bcOe31dVIb68q4dGCFCNk92zzUc7sMsDRxPr8mAmQV/+jYjW0uJe/t1Wps715Rv6tY8bCOfylI
f3BYDwYx88B9TAlvMyPiSkuzzT/qe8sXL3Jv5cCPaWdjpzqLaPWg5NPB96XYeNczu8Ov2Tposi/b
yxqGqEg9Sbi1DLku+38Xk3maOjGD18v3qVdeqUZBEGLVwYUnN2SFtyiCx35kka04GvrJywkV8KY4
wLnzaBsFy63B2poK/dnDS0vhwM1/4YvTzOqNUgV/f5A5mGoCSpUMpb2t1FJd36ku97ZygSatOELj
4ZiZrM53LT42uqjxaQW4vkEvTy2thZMQYD6dmHuVADLlMcssxxFhGurdeYO/pdBj6fgRIbCI4MvU
ZnB2+KbchFEXh0ovd8A1XjCpZgVIvSh3j6lDQIJ34SnwRx2Q8/KlICBmgklk87qDn/yWrHiof9sV
aBj/IuHcINeg/L7ISoViwVzXmZGIR+DD+klXmqcIG3J9D6li4InrCibgf6xYtRM4S3SzBBtu8fgx
sF5SjFgeppgxTS9OJh4o+An4tpapm/4lNxJp7O2Skr9KPiUiKX4kSkf+ASYynSQXFnMe8iAE+0p+
ARPihIKyjERy3gMiqeZ86vUvaBwTrdmPFStZNvwYX1gz5x3v0hPut2Xj2TLbzwdqLBQB+wVYlXIv
20U3/g95PkzwK1EuXwSimdDABBrYp3mrZ4iCmT7eIRubstBnjPPGfDFQsf0MYiy2s1OkD0U8eQbL
LURPbnHW6JEVe1D/CK41cOi0xVBGmYsHto2cYZUyXp6NS77kyXEbQ1N/0cUVqsHZyIfjMpHbcTAv
ZbSgTINxwe60a/Ktu8hYUNKxLgouLru1pmQbrO99E1RkfC7uMs6HCRhZU2SAxgMfvydfD2RRbMml
s+ySQHCCHp9Ohth0RVfaoIh3erUZikE2sXiwUDgosNkIR5bolD3xo+nixr20Izr4LGFt5jS8finK
vK6zE430oay13TNdwUhrzlIxWpBMthMes/Wa56CXZR+EHvR4mXAU4zOZHWbjaqnqhtgRQoLrhZSQ
+cbXXjezinedW+dh/iBhDadjRvK0CJVBmOSgJ+TYZGaGUQSjzntxlWvI+hEh70q5zufovaLlgWSC
QY20CZfgM/ojZf4F+5ptwinyR4FBjLAfhiTbu8VrnqGAC0zkvu5QWuWTqKAGdtFykgvQCkqY98h0
POkZh3+/Y6qxgfMcIYgvRcwWntI/7D38TF14FCnIFNh02jxMDdF5Ksuaz6aLDDEznX8cBKmbZ16C
brNh9tZqAhTIIZ5mNdIvovrvxE/8ob+DGZlGg1otNwAvQZ3AApHhTAo3o4/faFbAFUPAyEx/yURz
ZncUqWqfsBj+jOjYTapCKVCGLE7SZzhXZ7zL43EJtFORj2wR9LjxrngzVywARdx2I2K2iewcqxjd
iuYU3FpVBLpv9fwMcG4KIeadpPuPv3R5Ue7BRpwfULDYltk7z+b5qiX1kvxqHkWl0VpI/masJtbY
Im2CYXtArm3Xxbn0Ioy5ZhFpVPl6DeGn5PWfYNdqynULBH+3dBSy5BGraLt9rhwjSM/eZ7kw5mKB
o6AvXSs8TRg7nXD2re8IHMXvMrkmEzOJW7rA1TlebmUGR2fT3IgKWXxlKERFUFzm7MHE6/kZh1va
5J3uIFef3kUKU1/I0GiS93ocCAK/z5Bajw5umCTQJcOrdTC+c+oZ6Vr37B2R1wTS7zgFN1XG+9jl
/tYhIT3/nFrF2a9sOMlMZ3arWkRFNCLymTd5Sd02GbjsGsHgsYmr02oDmtDgJDqFs1vYBJRBBtkD
bdBl29ryPRrSHo7tT3ELGvgqrxtqWa7GhMGbqW+1AhDY8auzzv+dNOLqgmAUsmgtlMqa63rY5Eqh
JfnNcqbkC5rxY5Kl8t3VXDOLWaKTqf5DyZBa6+r01uEgjSb9vUfddzCYUQstt5dW1WhjQlqn7mYi
QpXaqDsQ1/ECrZXZOx5es2BZ5Gcl9Zjcc8nhNK3Xv4sW3/yP9dd0S3pY0Bx+ggW/kA7FRY+g43vd
rnEL0TJ+n5c6ItRAvTpS9P7jxXIlD7wyyfPMNA5Moa1yaj/CmRsHUO8+xr8yTCA/IRZwdh8/pHK1
xdwGYNzB4Hq8uVY8iEOGINX1+mzeW7RSDDf/aIc0sy+OehSUbW7JmuouqtNIqAFG50IZPPgFZlBC
eg9wSk1JvKiojE9nEpDOoLB+miKOY+2XNbej8waTVJdkYUtg6rKPe+Zs+FGx9hwdepzTFJzASWLN
cMSpytQqjRitpgMfOviR9sO9vtPBfV55uDbJINnccQXb8vnjA8OfF3AfXuMRWZ8Iua/4veFKVcv/
0UFwwZtx7Y5aSRM98aLzMB2Qqb2xgiAuh7DWUWmErju/0XYfjcFiFpi3Di/DNt2uH3vMzUt7NNKD
bNl0cko+N6ft/rjqcMiw77qpPMp/2z6iUDQddJP9WexJh7QN/fGE4DHjDOOAu2B71xpyleZWsq1Q
MRa4hjQhqej1DH8EUvzSYlO0g5JXmFL/WB4QCt90cHQFeIttiJXcMP+I/PgCYNnVkTAAvVdDw/wn
SN7oPQwf9eamIK/lXdOA18WPj2J695p/FWrufRxXkMdp8AV9IbRKDRzauCkns+er6n4F8P3fcMb3
+BDyGLk69rAs7m5mtqvhRT2DI4qHOlHmoOFa7Zyhqrl05vB2oDcULyM3YmfSZRUMVV6yRBi9b9Q5
E4RY8yQ/ailmmSA5vbaaNARPKoQYE1F6OmvKWO7WU6nA5atzdVZM9DnzpWsUdmFPiPyTgrPKcaq7
1RCgixIYokha5flQeHChAlfP+lN4SM4zCyukRHQrwlYewIYezOPBSDrGTNtYioLpegYgL3daTJtP
damduyib9x1YiT9y9pWl/FTU5W6IHUSMnrXyNi+DhFGIsOWYrWbnYMVWUyvRLHAor8mMVF6+7iUT
ke3vihwaxLO/BuJ37JQIS3jNUx0fePTWCP9gY9CM5XBL3VJIaPx1CN/UcMaQLyAEk5lFe4IZ8YhX
AqTPKLSXqxQ80MWDc5KYNZXM8/76K1YMO7OEG4TwbGvmJLvL2VrH4MMOkRKW9ElETOMarnuWarg4
5zjn5yI2jiRKEtUz0f/SOZ4dMovIFKbT8TOoI35q1Rsol3yuVa7DKReCA3MqRokt/ngcmFyKQbZ7
0w2zllLKpVKjUAJuyLiUjb9SKhiNk8KQObJRKr18HZrDX8IGf/kWrfPbgmkJHkbE+gbsqNCWaOsD
7TVyGom5cCbQS0bB37HDrPzrAvnnzWJhTgVdZ0RDYVBHqOK5qk6IPmYP/eZgC9KEOPa2ofc6MTC+
NELJYD+Lhl4oJmL8wsG+8xdXHBDY/qKfs4v7tWOckwbwxK8qCVX/5IElt3Rp+vrsF6aLEDdfzD/B
xWiJU+84F/a7HfqCo3cOCclUCP8d6s7OA3JUh/kxCGEy9eSJazK0nakJWVQOoo4ki3J4835G7tOn
YNORTml/FWBEKUL76ASfUfr6kAb1ZJOvHvM6w0rtJHYVqTBJSHq7nUCnXjoAtzpp+FsEiN9roVui
SxTaVtdM5je4WwTZ0b/C2al1qYay7OsroE0b7wHANwoYaPRSHSm2/zZX2A02xG8aldNQdC/wiB+3
hyopjcaRqg5D1dmHxFJTswI5NyAD7MmZHLfk59uPwbYjd8tjx7RRokeANqKlVsaSuI8OrmGvAjLX
o999kl2fJfhQDrXiMV6BM8vM7XzizV34hkiKUCe64TwzdYuPjLxxZv0cj2ObysAP7npHCIbTqB/S
KVwWg8arWdf/EWw6YIWbHW/Ijkwyy0CDtU/HhssSv9pR3o0ER/DI1zBuhgCgmGUMV80bhhza4j+t
YheSWKQY3cWbF97jKltI5ZA7mVVMiX9xR1cwtJMs2iWbQLvM9Fh3kQP7YARswR1kgGc3nJuRC8B5
XfIJ9sEw8vdOYmbvYkHfBvTU7e1rB0+eBw54CUJNaW1bv8ThdzNUZqmlSK32jFRE07Zlnqx224jw
j3e+Wt37516FRR/vfmTNtoxjLvjxn3O6vVTS/6o7PPotzSQ5vHOJ4xHQOHySR5cWouAcDvLcJPSy
0gYm12p/ZgyaVHB4IzW5Y1kRyIeAwyd8IcD/DLcUFG+4bzpHBvgSj34vRypE6X+XoPq6iMujjQly
5v+73rD9boRAQq/SgV0OUs0SiR2M8qvCT8W7zp2VYZLi5UjMTlguRbHYocCb77n1zaWW6v3JUK66
IzvcQm07KBekuinOK0y1C30vKdh6BHeJeK9S2eKX+RhDrhgpashg5KLhGiHorqd76VtHdEALn9sr
FUCiJowz25jtuwK94QMfpFQo+4ZShOfj0zhuKo5k4e7GfPDxliscwpGSrWIUm0LhP1Zq7mwD9oWG
asgfpPQh9Avwh8fD7Bp/6OEWw7SWpL3zlVa5mOcb9NlV0mLgPIsbKJ7lpPeyJ14LM941Go5cGsex
cNsKgliwuO/ugtqbWHlDs0zRWI15iDQRQUkf/SnIEjMvt/Dp2v9sbm4x3sk39U/yZFMkEBinf0xP
unLPcn13JtL68d341ohiU8UWQpzSn37b5NEq/1JIW+74uCXora+dXaUtANyj9RgjUljxWirK7L37
bJ7CmDopYJaVCTJ+x4vPaGRG1Ki80zx6se10mnS/V/WppfvnPP/hoWaXBNoqgjj1zUHEbBFfMEAZ
pjNbDm41DEH60rn0geyTLUk1HXKRTEodFIsQUrX6C52sNTpCJPihT7cYdF9F/NYJq0j9YUqVRwNb
7cB0HVWb2MxXtaL7EMN0kQn56PAF8vKhtjGuhDr2V4P56vxgmGuAEQT6UMBRxF9VEBLY2rBVVcv5
G0qpxtp4RxsA10ZMEDSOzaeAztCyM1AD0DrnC7kbwirIqsVgv2VFOxTP9qQCWAba0uKfLHC9DUOK
h59n4OfJSHc8HWHB5+w3I3mXKVzirp1+bdu4sGP8ouoHnU3/j3lx7mp/GjjL+LUUs4FqlJDsT3rW
dhpWrh8SJ/paqwGyCKtR7TxGgDMmqkqe5vFgZ/3GyGas/Q2d7sICgXLZJVjK6dQUMqtbxHTctsUW
GZx4sJBfrkZOgkzQEPLvmeQJG056uSHB/fWCv4J3pCVvRfyPE8f70fbgz6buOEQvQRqAFxTdNHy2
vJ8EIbJiG0XIe2YoMCoz2+h5xr/RnhLzk50ahCKjQ69Dg9xWY+jveJ31j7VapILvaWkTle4ZlFLB
A5R/xeUNy5U5/fGwunF4n9mRrVQqtwH6cD4TPtkPzCC5AC3ClFNPh+RBKW3dT/rk+etoSyaPgMv0
u7w87iNM0b9hhFZUEBhPEaVYuHmzmoisj/kE9FcrKysQTpb3/zi8HJwsKRslVNJ44rVczUn/qSmW
hcdQSaw8jcV4Q8y0Tomr28rtNu3CKXvKyUeNx6StLRJUezz7mZmZX11xsYrrnyzHoyTz/3cJ4fCv
beJt3kwcDB+M2akjwa4Ecvq3wRzrQvNpkJr/96eM0QmKrnsZtWHVbfcgRjans1izbCHNA1+jRH2b
1wQ57Mn1chaKauUAFABskuTHHPFRDNsOU9VHxXu6wRFNmAOvTZwY9k1kW1r8W9BNH8DPsrszka9s
iBEji0O6wZrYylgLg/9lq14Mozy/NnuDG4ymTq+6NpOqY/LeekGQPODxy6RCl8NvAbi5c3XbnHL0
MVRPmOVwnfib1KcwrhcycoBGvjknrYymSWrVgxAG6tRRDUHfpz3LSwFxl3Scnqa6nNgOvt//djWA
N4D2YfIqcXIt88vDA6IubLPcZyxBP5t99fXd4Dje6T4Fu2saVfqjnCnJnnhTIA3IesoyL7CMu3l1
EAe1GMvcjAbhEzw/Kx9bsHZ+cExih7lEM/QxJKKKDDQ//zqyiHmC+H7lEvPNvm2lm/GHh7uND3VP
LLi+RWkXkhHVl/8yxybTQfZYS2FjzrVqX+kX53BRpSiqknwdJXc7BUGlTfNIl3GBDBsRSC9oskYF
nXqwfsODD6Z+PC7CVWGCn19pvN0YC34A5qklt+5buO4gbaixxU8YYoQ3PDLz3pHFRj9U6FBw63p3
3iWGy14VMYZYRRAw/mbPGXTsYfYn4yESwjXJsClRKbJgwSzo2oB6/AJfqeiPuyhJAgyM/LITaSDe
oKh7Cf4XGO37OIUY5FBBYnbO3E9DB/Us7Tp3CxOmFt24Su/L8uxEer3CB//tFrJ6LNwH3WXGXCps
qo5Vj4ohufOji4Vx33q3URA9kgEE3d0jlIgCnm05Md8HndNw8UIihZ/yDX6F/uWsiNmOiR5ZiqGH
45u1CDzASQhdPv62FK46pIf4Kzm4yyWgHuh+7E/Xu0ImG5xJXdultqCcAzd3Z2KjAbNqKQXgexmZ
dyASQk6wP7Sm16KrLnpmh9uHDOYO49oSyqTgNV2ByddQLjbT5HWOkfDq0enH9phXBib+CyA3iu9R
PH8zLqbAbLyyEuMJ6yOVD+/hBiroGMeeomrf2egkJKuWMm6cMyfAudcVCxA3xDY9yzBTrOFnxnzv
d/88srZLAQ7bZusWkFOtlvDeCctlsmsvc4aZ6lg9DTIwJkw8H1w3lxsh1rDnxiGO9o0lsdisAFg4
a8MlKFP4FI6PcI1JC9rN6o2DPWpfA4USLy08D+70ukf6VbgkI4igo5LtKAs/FAwy5/SNR2Kj2SK9
fzojyho7B85gXwLjaaNvfiE4Uv9EvaEp4v/gnUnSLp2oGqBGpXFi5R+Iqf3TqOO62rkwXA3WrTV2
50Yds0HPW9g4D9sLYJqkKyg+M2C4wtA9fC+lOd41VcdfI9MuSwdPBdfx4jkDGqSMd9we9xFIIWim
MvDyaFzphIWxtW9HBspwRF72+Kqla/Ea8Mq6U5dn3bIF43eg2dSroNlULgvcan34Xjhg/ZC+XiTI
SuLs1Tu/ujGL00gQQv7YeXpp19UyYcDYEbMdsf4VW9jTCG0kvu5WFngj25bx2idKJwarLzeQtGS8
6h2K/GWyacyOYdyBp4FHF4iIN+SjlvW4+MUIHljkLKJC/bdNyZob6J6ulKnWMv+Z++uTAA/gTlnc
FYMpKWrm/2e5ljA4V39PEO2hUAoVIm82YqLHelxhFdfzMBsCTOBc5ByR9tXfWTIEerSmIFtGf8wS
yzxvYyT3rGSpS5nE8HWJMwfMJeflFwx9vQlsg7hg4J+/1BP0ysft82F5I+vLbUt397afTK0Q0+ly
s88JNqHkR6tXrM736jpTfGH+/3tIc9AdB+w/aoi3uvpR61t3zdvSn9K5TqAZI5PpyNoCWlShJ7oT
S8LriFeo9kYWpJpUTz9kPLi7wp90M6DYgl0rNGpLND4jT5XW9pRvPf4UlxvfPApocrP9DRCFjbem
YcGyPBHP4IgQ6+/Vm/0WXpI1tJjFihHC0xDm0hrryX3JAd5qX/NXgDRztTzNW6aoPjcx8H48qSSM
XBv3PH4rHblHs2MOvywuFpB8opVMZQ3qz1PYgpKb1896u/jMyph6h3AhSBXzR8qzY3/7pSDfgD8O
vkb7U7fiCf6Ln0j6QI+Cu+xYhy5CnEtkygPqcBzSXz76kvGswEAT6SlifC0KV3C9GB4D6wIZzO0v
ppSD3i6ZXAGyrbLzv7/e9CfLDBawyPcpwqKP3RCCfEBWALZlleb6sU2uGaEzLBgvg9wMeNpe7pZV
0ON0Pq5V1UJK07CMHoHEhXNcYwDs+G/1t5ZW1UC5DUAj1ZhMCN2u9MYDMW9JejTrGNQ7pKkpNQqW
ALvEXIcuM3LLk0EXX7kiF+q64TLOEVJnoetlkW9JqdIb2l4kaLCpTgPnHf9UygmsQFNKv/bSYk/C
DhVdujtcP5Ubvc16o7J7Tkqv2tUd/9NLW6LqXmqDgE+JRJ6lXBiURo6jnZDd/GKwku0S2NmAkBZd
e/wEEjocX5YRwwiocc7ZJXrdxbxDjmIZRgstTyEqtb6SUPNU4gc4nI9axIpcDCOp8dgUJ0lylMUs
aQiNm2Bq4HdT8vV9SXqCBHNbBEI4zKtZ4dQSbcNYV4A7ErfMKpwlmNGja0bNm2Ft+hv24P0gz4W7
jUEs3Y5wl1QA+Mj7z8NbmUL+z9FnSJLHtrzF/HnITNgtR+MNnPa6M8qwLvEJR+gq+RxA8/4/Yy70
NX4MCybVJcuhkvKFr/8VJ34HnVtRysHETO/iVEtz5NsI6sS3ShTtjfzbwaJoSJKrma2tW1JF+Ahy
4URYP9ey5uMT88Bf+9FPJuXuLWT/2ivFH45MIWXoMkJ9lKXa5zC/VWXfHkU7wGQ0nhhHtb2RrOY+
R7xUKWvaTIaHECSPkMSeF87ImS5DwtLActBWXAGww4+qJRi5jExfuP+jybViSaF/FFFYL3+CD5Kt
cOcfe20WJDQUdRAFFDHZJMnk6Z6COn0GDPCbdVCyopYAb6a8HhzHqghYAGaIYxHQPGAdayZdg1V+
Q2M9Q4b76bfyyioRKCW5fii2+pjr+NdXi0U/edTmTXsc1OP1q7zwYLxMM6ZPhzXSr7JWt9+KxUqR
wkiYy4pbFRsCcPjcNVTRu6bGbBeyai+gXkIXJpLA0KcnWotTKvohLAiI5EmuQg+Gvu4T8HMwgdq/
7PsgIN5/4PA0+n20lGb9/ZWY0hZoSCFdcJ29A6sxZLuEn6Wob3QKbKdNBZVUXPXakrUtZMK8jKu0
0pXX3GgKVc1NhFL8qPKV82f8Rvslbkad7SwGpwMsDe9YaoXH0MT09csdlClOCGZ0j6P77Cep4vNN
3ANQtpC8HmDq1zYK0s5YtEGvRyVn3HYZ/e8dAc35W0Au8bmhZoXEEOBCGCe0K2VT5UrbiEaL6iSM
utjSgFxrQfH9om+lyEMI006lZEM293xq46yKS8ge9WzZle3mml4UfhU4dJG+k34M7gyJqfecKQmo
uFnmRHdQBXh1DVokn47N5w+R+3Igi6kge0AK7jVDGkDlPEex4ddnh6yFC2/Dfb6JLac5B94KGjHZ
722dZX9xN6ol3T+92ws3+qLduL55FCY9V8leFLfPp1AT1vVmzx8O2masa7ES1E7GTtupJ3rYwIvJ
ANLuoyNG6gSwv16O52DATHLnV/7HBgY3jVfCgLpry1f4h6XRgjM3TAHFOqG4se52gRZk9iBNgODh
t+siRsvsLCV/QlSaDNXjOyiQoDXqUmVJYjJmEhlfpfiLIgkurR8mGN8MBcIOAaoERHubwfbyGXew
9cfMiXDgOqF6Y5pQyQTHIUg8RyHYSoUYzYytTT8cQ3uNs3RaAjy7la7taBmL4ci36Kza5ssvnu3u
h5QEzEDc+XQGocjdImCFw3+FbLFj4blzhgOEm5Gxw7DfiW8jMI/jE7DlArppYhnL+6VqmTY7C9t1
0NZxXT9EgKOrTiv24mSK0etlwGwgoZZvLnlH5RHzkA7zG5mUK6HMpKzLfOGFD3iQkIJfZFaYS2pt
2kU01E5CfBVAftCST1Flx2TG6Y2EO6ZiRFu5wBQF3ym7pEjwElYqHFi0pX+6m20LNY+8E3mnpf2I
/NrG19mvlOxpKKYudm6vwn6SDxCh8u/VghaOMz96JyDHvIeyob/3aGF6K6vzQzj4Sy85wEeW3C8A
LvHLtm8NgUQefXtKe1t/Dgmnq7qJ26YRQjlhGtCKis7xgaupMsU5cZzqEGdV5/2VxLTBpY0mjuOc
aEfAFbgN/6zK4lKXrXKy7RprtgML+dxr6X7AZozsQLcokohOINAeKmXnw6RE0zt54Dt1nMFinroN
lPpn9YErcbvtXOLQ9/GION/pfjl3zHMSylqlCx6CY6XHJ/cEA2pNef+wGBTNpEM3xYR1Os9H7m7s
m+evi7S2AivmbU0MWbZGEnL2BEmItrYGNjCAzNK5G1ffzijzxDSzykRMZu+eXnANg8sZk/snfA6H
yhcmvtommVhxEVJjfVhASeEiwwNleeNmTNhQnRoZZLxpD6WYnZrpFKlFIbJ17oVWw3O6M9fjVWy+
ez8+8UuPyjuXqYd5U//LvCnzpMtZ7HTyk8Bp4rhWJ8qxdGxoqKZmeZnHOQxcSpwXK4UMIbyZN/7X
7ty0ifSz9SZcEuFommSd92DIooia+U/P245it3zLsf/JB+8DkZZcPgS6YzHuXHKptiByl7YulsHL
ziuI9hhPphH2FDTndv4mArfHxWDjrA5lKt175QpVlWIanFREwTVc/IKRb180xFehtDPBv+0fyjnN
XjItM/AMPdbBuGAr41KlZ6jrOiQkjR0xxQGXUTKuvG46LObB64aeVvS/Hff/8xXDVJn6XhCWxiJ1
KsdTmyoG9vFHrfifJiXwoKKhWuj8BARmp8S+9m6oEaX9sw7AfF3/NyZQv0C3NSwz5QSr0kAtW26E
Hj4RiWjzwe/6z/bg26YPQChHPQZ66xNYkziFUDQ2ZMWTgusyMvOoC60CeStLHu5cGvgrbUN8r/iw
Ze45tkBLI6pgPMxaqzRAR2sgK6AeUgi4PUKGJQqnWA/IWHYQox34wW9GzRzEPws3lpK3baRmwJcv
+6YYrWMtgoOKd8Q29dxcTRi41Ckk06HE0CWlHs+mX+B6yfwUzHFUtL8wUOHmOfiEGD8K5x7W4g/z
yJAtYQw8n4781E1f+ODQuTAeOmSCZiXc9mk6CBanLkbpwqa2nZLL/FzU7NYOfWDunKBfbduEO3bl
UnHbNDDBG+CsKmBfTXLte1mt4Ewve6Ir3Q7Z/WYGf1mzmDMFj2GiSROezWdFuhjaLSYkZm1J0hs+
1/kwXsqj0HP6f8sc6nR9DDfP1mKsJ3oi1298NKSRTUyby0aIpBDDNnmeBlKWR9+NewrvRVvncGKk
VADPaeHu+PghvT8lzp609Cxmr3TLWcfZTF4O/T3srHCTmpZla2pIsFc6TrPuF3q7FHk2JN7zL3d9
SMB/rxwbxkFg/ZPDitAyVJbv0zy9jJJxZXvOzOX1MUFkl5+HOsQj2M1GIjqezaN3RAvwisg7tvqL
r3qRld7nmGdpTAyIn9tbXKudlkM5NjHRjYg7BkTJMound6EgMQL6a1DO5qLugULEzNesCmsw2qyg
9rIzkdvvPZ+Fv42lRrtmLD5iMumoE1vBzINLouYRwN2uKzhEea8CBZ4XG//ZerP9VkHfCR+zxMEJ
LBHIKPO8KuKqeiDSff+4MmHv34Ixe7lrl45tfkMKcrIb8LZzYGgLNUV7DUyMUXsOlpAuwFMyaF1i
7cxL5de232KQgLTcq62G8x8X3hdoBFtW8/OJpRCcP1TB53fnoKf07MXfy+9QVKsFio6Eu1zQ14ys
8F8qfyRRSpNRNvmUbz+TD8OlIVH0HEtJiCYAb8bTg7LUvx8BWMOx8t/aIkIj6nCj8Q75cYzz+zkd
/ZYSLnu1C8IQqDLKyy+ePmxawedF9iOUXa7RufQAYNr1mm4b/gXyKncKeFjKIJOJdORGwT7JoBe2
49qTGCfhm62BiJz9NWTRIMyn/RHbhG2sDb2WFx1ZvXQXlHmGBL7QpRBN3b5sp8hRdktXa7FWgqFm
OQjWr7oEbYk/AOXxxxlg4vuCn0cJSW7+q55L2A3F2eW2uPo1/Fnx3AOchN4EKkV9OWv6NZ3QUcf7
2994hnhU6PkLFZ6JwJxieICeGhRW5qHKkHVuGLF3tdfaSVn8JD/Txq7vRrcA993uXXyL5gQ87Eyn
W0JSh/kYJmbwY2jC2Os45NB/QSotc0I/zH5R5EbroEajJ2OBftTg57h3NRreqUdfZQpYPXfbOL2g
nrr6tEyeSoahEfXlU0/IhNyhsmIYQd4arLmmKhiJJheiiw+MzBw82o06PyTtBHBflN8gnnZcpdef
OzSJ5GERvZK/fTutuIcay/OTpGccgw8goKWjHumSpFNOhpsF51X7wbBGvxA/w0KjDeKCMCOwzRsK
Aealltuyk49mS77hPfUZq1xJGwX0P06Kyn9VjXoeAgLNbHz1CMyUE02o72vSxCNP79yVpanWcF4w
hE4xy22J+cThfZTvxJ3Xx5yETbR6ZBtJo7QWJUz7V71S1F4IJxR4+Tij7Yp+KhOkc90GYBf/Ofe6
Zb8XgAsUYUbLF6CyewqqUo7tB4D+vjgLqHgJmtRjv4QeByxSOxeRWPmX7CImJy7VyALYE3ZBgtSN
+D89znuv4xgGGd9Aotx6vwzsuiGgpfOgk9P+WAfC43uNpLlGjBDFr+h5mY7vtS2gv3v1nkwf1XPJ
Uq1h/l3oGwVh8iOt9iThe+a6G/680DLlx1UFsaLrhTKfFp6r7Ixy/gPsDLSUeWMsKMQusuXnB3yR
pldKt0Ttr3BY/4/5YSB3NWdgf0OJ/7E7ZX6OEMaWJIVoXzDRC4mXqRIE9/+ijQMztlGmKQD0WMv/
E0++1dOTc1rlxxqJbd2/SG+6YMlZlADBn3cT/aI/q0Pp1Jrpa/ZLlIwKAE9jSRSpVH7iQnKm+7Na
UxIEX1o9IIuGEHw5HtwJBSysnubShS931bFJuSSNSpNO+jJGK/Ud17Z8vBDN0fCUdBs9VTNnhrn3
FIlu3cx5mO8mrSy7wyogmsY0UeS2003eeCfgxT6NF69D8xhM261XIidpcFg6g/SEAJfnbU5x8xbz
6tAbxWMOXwYaa2sQpKfhALA5kALGA/lz2B8gziMpw8aDpSARrKrNsglL9KDcqRDD+3KooOg8SWOJ
5Tazg3WMWHvpORsmRu3rdVAAZqd4MjJKjVhjbyK2+qF+HNmVSDZmFHX95zD3Dx5e3wDO4sGqQzmu
gcetp7oO9hggyXj/AoctYuuFgag1qj1DjyzHN2+8W7ni9WjVpj0R5dbcGD18uUug+EuYwb+1yahj
MDQV8TkHQZSsNbLAGpmJPLiPFxrqcTs5RfQJULDAOizyGo2iPrFh97WOqVTCKoOFBcwc4Tj+yVY9
Fld1nGHzRRQhGJlmPDd5NgoJz3QtMaTnS7G0fM818s7degZVqWlj2LykuSEoPhGfMDYRiODaULMs
4xaOeF4ztmEz2+lz1YOU+6D0sD1f5Qw9cllzz1MeXkBUgYwD21HBT0+yV/eP7CmncxHEwgxOOvBj
WA7hnNBjRaCuuiWKWi1DJbU6K+2H+zHX+Sgs5dUm/KY9y+H2nYOGndhhU5ORmhQGC9Ut8IfNlJ6X
7FyJky7vDc+8DFpiPyzf+v5+vhVjOuy9y/ShtIqE2PjauMxF5kJ94R2eaQhsuk18b4LNkVTp46ci
B/Bi4ytAzUX/E/n47nJU2Hct8Trj7mt33xCi94JPETX2SDjNEkL/n1NPG1HiSoL/Mv/jh7e7G/82
OLpxjyU6PiYba5hyI1Tn0K5FJvWtVWwEoKB8MX25Ryb+Vef0KbwNK5Bb5H0v7u4mzWDJ0wzAkd3N
1rzb96AsYTCm+Y6GWIqd6/WuwD+VAQT270d4DWyhhP4P8tKzHHWqN4s8oadlNxU0kzAA2eVzxhe8
ZCjVX0F/ZLARHyh4JLF4vODVQPPCb5le3Q73NOWtHO+FDyCXpuP6uwORl+PcdnYbZ04JUiv64Pyn
n2TBzc6n6PjDWz+i8yxvT1Zlb6USWU9xywPC/Z07BMxVC8llkHemlVhaSugZr61EBM1X7+Jw+6pX
MzEwT93N/sKimZKxDzOyzwsP+Avumaz+52qIqoudkHtkLQ/iN6t9412uT4aiFi6PTBjY4LwGi9tm
mewOCCEMYExm1oKveZUX5i8m/qHzB3Dosj1pglq1ss2hO9zF8P+ISe3wnXS9i7+ht+OLWIIQMy+U
3qPXH2MXaX7xYPyWH0L2HF9/GDC9cZt5lXOmC/EYuuA9eAGAo8WU9iLADD7MbHCwHas1Je9Q3ZNm
Fr+i8yVBbi7ChC0HBsT8UuczOJef1TD0RNoxsOBDZJ2wNwY7a3pHu2UrUqGq3PHMQ1IHMQxaC/35
ewDshleo5UmvNHkdoa+feD/pxcIjmCUqpOMzwHdTfuZLXhI2txJyqpTYsKmq1pQSotIv0Hp+jqpW
KelpUwEUbWw0x4kB8jikolplmiDvtPQ6ZZvLVGSXjPZhaVSxFcxd3r5omGJ05SsbmFyTlOCsztHr
RWUlmNYGSqgzWGTFUrYYU/Ty6VognAgLCQUZKt17SlRkIrPE/7+YCuGwQXRidzlTU5bGiLVzxy5H
W+kOEeOqeb3BRgNCzA2IFCE//wcnLSd0MQd9PZx8Y4czLpiAdESzWPCf26C6j1SmiWK0tfsoIm45
wkU2GFs+cxL1042yBEPy34QxgL11EwfntkG+L+MnDzEMhQgCcR09hKwEypQPQ0rv+0zJ1568KBjJ
EzUsoVUEyf4HYJIaeexTMwr5cw8NgIkvjWe1n1/dYBZ5OogRKkwJxv5I1PNMn1luJ5yZJeBceDU1
747AYbfB+KmMJM+ZIS2AUjBq1VCA4q/W8RiL7UkE8T8VALW9xZrMOCM8T1MWnVp8xjlk7dpnAeCp
qe9jPEidsx8+AlyPZF79GUI45b8JqzmK4wh8CHd4a1VSXJW41WxCREpXil3N/2T4A9i+owIMVKVk
UZq+qu3wLZ9NY51Qt/aTKEhKWd2Rgj3Fmag49gCUJIyPBZHjynUCO97SdFfYSg0ykPb4PfWS6sCo
XqUmaQ6jXL2XRMH5DB/cJdIHMa22LosZRwF0ML1JuEYew+7ko0UxFKygmbK/0WsKIDNKaky1+Pm1
juPJGwvfkACXoF/WqrvGggpTPF3gD432P6LJKXhNnHcF62OK2X0YlrVb4OnMRBDwhhdC0rDZZ54H
M0lM5LyyXhWp5po87rkn3ugwkqOaRrAuqSUEIeoL+wME+Fm9WwAolwd3eSVIOWsL5+ULKmCBQ3ja
HYC9EB9sUTxsAFSbs2JPulItKE5/o4UbEPnsjuGk+xGbBd2ExcgjCG541d2PGb6Ru3xUQChmxxWK
xmiwc3+ivk6TysTrHiTHddAAd4Y5vMHnArk+pUNKYCV1HN7JtpXCwzZJbPqI8AB1pCwnQ6WVCeYo
NQDwf1mH0Vgn1MI5mPuNQvVdDeuFOrCP2ss46PLJemsWC222G3qiVc2GqxkrsapQduJrCkqLJ840
mL3nJagwUEdtroJbYurByw7Di7A/t2zStnvf9Df7B0M0WSDzdzFHDkgyvFvJtNrt+g7lDIgPDWNB
2iN/GjYKllQig58PrBy9dpaFhPfBmUDmnH8YyLvOg8LCqgGjTze5/HhEubUcPIWVNY0TzRydwvWl
pbEzDBJY7V8EJeHxkAr+TP9TLLulscWRST6aiRnp2FjLOIUQ+MKbdmqz1m/NTN1wk3bOX1vrsXxH
/rd8a/2dYVAsgaF5TODFVBM1jTFLHKbRE82RBKo5Iv3MxIPpbOnmHny279tU9nvhW7Rqi3jSWE63
J4hy+H98RoY9O+VuxH/QGyi/uvCGVilPlYTwhO7IT4feIVHqwWOrZ6LxUKOeihzaq1uQ4cs4eZzl
SO0gUuJHm9Iq8gbfy+IbcAKMsNCyhFAc31gBl3lacYw//17W8JxgAL9ngZD1YYSluMUyZEkKlbik
K+AZ6lYcYnQzpy5g286uqOKY+FGxX9iQOX3bwzJUwgCREFvuJkl1vKjr58xWpxXnVSn8WgruqDx/
mWQj6QLJOKxFgH2PRHdqyQXWtDaDLJFHUelpW9ZSWaJbtttwA804K08j2GB56bxprulnIdJdRhaf
mmWEBBCYMnRlu+jmDzK0ISzc0s/7UmU4i4rgq8mMCJ1xDNC0ZQvqo51knVKLlMOiuI5iBeTX2noC
y2AJYoQ/GcYr5eMs385VQuJRRguJ69i1bW3IYVeS5lqLUCptTHL5IA8VLj6RHSAFv0SoR/kcLmA4
YlhbP5pKOGtHvPqEA4XC2cRDDoAOC78eaNySUhiIfeOJSOfsa9YQZfGkN5fueVUuwIzYgEDxc9ct
Lb7dxpZByGbFXxshyIA/5L5LaRCB+9JyTU7h/utvR90k4U4VKRXTtpre4SaZ0kqpY0gb7YAcZ31I
v3xAUMEDYJV57HyxDWW8KsU87dGCOFAImT4CaQTvo8GIEfCVliH01xUMd6iNhPNpmDJz8o905/Qq
xx3hAS4tNr7tEy5C//emfB8jvMGGMhHhHUbnH1WlvMCF12+EaUsHTzlAwIVBPlsvBkCTCs4nKWSr
jAlX+7z5b3DYuKkW/qrqLwcG6fS8GAO6JEWEbXHnyCg0MxzAIZXg5ahXZ+lPEom268CEGobpygIg
Mf3Z/jVSBqomWw35/uvp2qLff7meDolV9JPdUga3hCGo80uDzVtDXO0yYLMz0nP1O47bAWUibSNK
IfYok01mi5PCjiHlM8pUB9lRw6fbiAK96U9RbLNe7atRI2HsFuSBsVAqJxY3bF4x7hbJW/yZPuiW
0pRHTQDOvHTD6u4DyK38qIoXd9SaE/JrkwjZ3iaDXmbNFfvjB9vA6aJNZslrDmbiQl090ZZ5qnVP
Kqpd26WMfnP9QvLy7JOvyuoOo26/09l8z7nkXP8E96OiCe7bawAkhvD7YAChTcIxfNFhGeCyFWhJ
bMZtqNUxvBxNp5AslKZfXywEXKH7q7mhoezC+I7z3YwGcpD6f2zPi3EFFVpIb0JNfUb5loSmwa6G
8TNHngX55/kt/ByWhGMo7tD55/xSXeRs5p818dYv5+f87Pb19SdaggRNoeB3m+h5ffP0uA8A4g+b
mx2G5rJ9iZipOoMwskZMKYwN0AbsOX1UerNlcybNT7I7K8R3ExkneE5J886S4mVWuafV4GM5Ay7j
0AZwGGfFukbwqPII3sAmL3tEf3FBAvHDgLAUAo4FWI5kEI8xZl1hMsbCpYJ/jDi7BlsQTyQxDbFG
vpV5M9lBokqGIQx7Jum0n0id/pmjf8GwH017RMmbhFJNicwXORQkJHY8g9Rj3QIEBUpEeQ+zsvjd
Hp+69snWsFludt18BKCsJ9ekNbJVTQ6pzRPmZCBYGG5dRg8AhhW2H4fLxs10zziCsdRS9equ9Svo
A9Zk2KGN88Lpt9WslyKK3JcPo9GPGHw/Swjf8pswvIQHzekpgR2WrlitBY6DVG034Bnssk+4KxKr
7LhkUxMwx/oeCb9/ftSYGVf90NLqLF8BZg/kmCWvq4pBpiwdsiEsWWfpll6jEuaxf7L0r5IqSyTZ
bGOKPdGJKwLqnAldVs2MaUMBPBTj0tzMXTOUsTxXE+kzt3uVagVaxQP1Uhwxv8FnQbCllme2pr6m
ZbsBhPYVApTvuhxavA1M1Fd+vrLPlxZhhqz6RIzREqoXPbm3FOfoVngyVRWWhV0n8IefXd3czTx0
rnhVecvh5jHzpgcTeAoVVcb0+jrZ9Jg9tlOJPOj71c3GxWoRUPaGIRzLmdfKkolEKcQTBx/jIStl
J34rVrYy+w0OIP4+TBMt+hsxj0/Mf//mqyj/0TyP0ahUGlsbpHgAXj0sQ4IkgoetL8c9SdOeWfUl
7haIsHr5x8sqIRHBntSU6aX4eYnOhrVF1NWSEcqyMV+v5ipGNKypinQJgVgZfvaoMOMAjrCO/ycj
KMt60kEEw4KGnuGE2lqPG/LdvgdLfWyCFiGsQ661RRs3uuUlyLfSzufrDQXxwuBDSImZFfMkIJKP
Fba+iN+31+XZ6yaDJpQaLaZ2Zb08BRbGO1Nvmbh+0P6RI9cVE3TMtWZZlWOwf17qk7gpjlxaC0K9
hLXG4z7nLwqAZ8cY3KeLRTd4t3/ZN/rH79xAt46iYGeTlFSyCR+3j6llSg8IeshpvbltN91blWjh
xi0Lc+Zw9EjCqAbyUywn6slaVYunOWEv0QHWuwNYmsCqW9gqCXESSpsIq5bsZ4w0yrOxYODxBF2b
KNaCJdgKV3QSqQT1LxqdgCmxrU3LTRVpYn1qP9M2ILBZviMczO5RdZhmgUfwYAhxcQfz1w/3j5ny
SP9cyFUcB3CQFZcGzfl3Hgf0sDuAbMGJLMYQf97g8ppQBolG/Tifq9pzpQL4HMAYxLcoTVq4YIMz
DanyJNn4KYfhALHjz3vYUJOaF4NTLSXWGNc/ocvxnTZylVE7rMvPkpQcL3Ax+gV8olKua9Av8BoU
PBiS8Z0o0NzzefDH5WbwtRqtILeDoqJp6j6xuWx9MfA4Blj0wGX9vmwNpqoxAyIRbeRo5kaFiDJW
JEWoCDtBK2bEjS1G/4yJmhOa9CCNRifRxFkIScOKzCQ/iA/88+Sos/JzYEl6xEGwhYB6tCORieKb
NtWp/vr2sz7mOmcl6dyxR30skEniu5r+qxwlKu1hL0hkWjG3gpJVEqphBNNkr5eOGqnbb3baBg+z
CxyB9bj1C19jjFcjVFOyrMVAsxA+Gt3Hi1T7HsMndx1pSBN7cOALEl5xueEPrS3HHKIWAeYOCqla
79qk6Rb/54Fs8LsyGEu1zvAMGoAZicJcsTNrYmz1S/TWmzqoHkcC7vKj5oElgPamKecVysHScV2j
KutHUhQ/5Z9VpOZVWcj/OgiRZw+WVhLWO+wq+Dae8HtysmPOc83eQotluxh92mFZqvOBN5Kjnm60
NkgpqlITwzg2Liqeat5tjbuPIKj7SREr22TC6k95bYorD384A1KmbDP1EmkEAAYfAxIV6JDiI/+v
UYLI++fuuhvP6a7cBT1DagNrZRz1+Iui+uRms/p52cReWbWN9I9XAi7BWfjg2G8QkBr9GFmfHDk+
knSR1i1NRKOL/3PI4YCqgJkfMyHU41PHs3UW+x19hin5mjtSYocCi9dlULjdeOp6IX7mIybktQoC
sLkKpITWXHQ2dLjlc+nmXuGBXMAZLqreGhq6JlHSU/doxvvh/Zbyq5NYTUKAsseZ0AaZA51PQoX4
Yy88sPeQkC+OfO0DD7MEDVQlMrRmjhWDlQ4/jLl8vd+H6wSeiTYRNYwtisDiHNtPeRd5g4qjX8ES
uDBW+gCf5m+4y6CdRWB+14zxRO8cvr8wYE84MmHkCsWoVguhSwMgw4mqK15PKnB6XyWzCm96Q4bV
cdLsMmOrMGzSdNf5TEmDfIQR9dxezjwTZbfiejHgIbbYN8NxFTR/s/4xj8dl2QJ3v4I+2L8K9W3V
6iSmaFpfCTJ2kBuOo94VCruJML72KnYmXl21qqSDGl01iHH1xf1p6ROItt7P6G4689dUOpL0SN7j
E4c813WWCZeEOXw/UnH+Vt8PEGNZNEmPc36czAQ1G3mGJvLswHRA8oT9sBVt8Z0HucjGJjAhhrMK
lP3uf8IO3haYSm16WIbaM8b8hIYWAAfcRoRSj2mRajjRKin4izU929eEIMbmqi6MWr8r12w7iGfe
AQDhclagxO7lAvKwwA2xm1yVIZgkaTe01ou6xKUZx7lrnUpusbbxZUsuuTfa2ryYcxMeoNULsXU0
8ZryaRo/G1ReqKicDoEFJHb/hKb0iNNvVNVKnZwefW3nCbTkjqOC+asz/WtQrg97/3iGdAf8gEm9
ds+tBVBTECaSRxf24J771PBxXNsXaBP03f5pcaHueSw61gh3L4pw78bG87elY3cp+5rgWbVbT1LW
KIM/xcmfGM/s8xmuqX5wdqxAjo6zTCqgB0iWqgjBl4W24zHEvRm9QUtz+szda5NKwPTBDJNJ4HNV
j2wwS+5dVmU5NPJeS39gIB1d5mhDz2tMio6K+OKxJRJJqQp+Vwiyf0W6YM2JF9JVXq54RIB/72Ku
vuvDtN+mk8qeyO04gXNbxU3mjwkgpIZg6woHs/sJW3s5lQwrgKreRnFzdR1Pgji4N7L6o1fxCe4B
t/iWf8jPFvS7ezFkUJa42hCr2Xl7Bb+NpojoVf7dSdFLhClppL32bX2P0ujVrBjynEH7lcZSb0mb
4nfe8Hx5Zg/zfBgNMVTwM9BI++teOZmJxIVHqPNalDnzMgnPNQFPTyOEBCHARly4uVou1fnH+SMA
RqkkSXMDvdUBLygVIM9EN+XQd9NUETo/gzkKmzE7tUAhP9ObPHCcbEeOozxTLjnO0/dJCyr0ivNS
b26RKbe0sn1N5C2IJsXC+I6CE+NrT+bdlTzpjxk+4CTNxztOh+zKWzb2dsmBCubyfUaZtDD6i1BH
IBmSV7Bqrv5NJrZXCem4S8jAnV4Xqx1dM/ULPPmzQ3uH4WpA+2ML7ryHz6iup23Se+PvdDRtO7s6
9UA1jz8gCCLeDdXvTLJe3DYAA1X1wRXH4n2JRXcZreX/E+KOFfLOwXESvu3lRxXlTY5VsLplkuy+
i3Al3/pgssL2DO8E79iXq5UPhBW5Ipd359oXELZwJX2O27hBMyu23blQjNg1unR/EIw9kZ5VIgEK
LepiqygJRugBzp5k4laA6MAVza9djMcTRehISuRJtA+VcKQQHhkAq7KHTt4fGciIf2gvcoUUP5Ra
8xym+uMX6sphjaVYOg+2G6Wakr2lEQynzlDu6+9q765eX9/H/Vnh04JgR4Ri2rGjRVOqRTBRQuNP
IM4qV+ut3DMRhFD8dxoLWSwSzcwq8aIS2Ym+uO3RkLtVxHy/cLdusOW+n6yeNT40EZ/+iI/nQ2CF
Nz57tkReNSdTlNui/7DU2KDFBXE4VH1Ke8j0Zoq7YXIsHt1tIrvbw015tShLr3UiJYYqP/kMC9eh
1ev84WPOkDucp+Wni3/iaasB+icpwTbyZdjzD9H/MMpNMUW8wwuI39GFo9uI8oETBvyzbsx7PQ+j
S0Xnylw8huLwZFvRLD/Mlg0vwvGrhwslMOeyDB/KVMcaXJ1CSCu8igBYw+c3QJ8nN7pKb0zjJKfp
3B6hZX+qf3RmVUnRf4BxlW8p+X+/AOyYusXnsHAtsdbcExUrhdIju2baZQGYSKTQsvLZofRWh7mC
iLIPkz0czdIzhifKPmpkO5iQys6ejuHt/6zIwaKONrt24m40OBpJpRcjfszGu2hvIcKNlrIvqFd6
QeqAUM+COsQ3+pm84oAtFzX1fqgbQIG8wGNsECy1p5ZafV/jpqNvjMx3wAdY2JE8AX/wlvvefDp9
9lvJ1AZwpxkoZyiFPyIVfSbXIohBrO9vDot3N29sDbrIKdKeGwArkJKa99fp47pFixan3Lzmh/5I
6PNOoa+weN68USTo3EGYB1IHaF/jJcrhYjm4N7BUmqfrh2JaqIEtDlpUAIBHgSNlnGxzp0A9Bql/
F0T+olrSciPA+gHHU6Lhz/Vp1XGmljGR0lxAG0+Io87dY9L9zshlFYJgaF9VIAR7u6YyhKOlxtdz
NVlF2+0ieCmB/YvSl9R9vmAqZd/LEJJWBE/iIU3uVl2GPHLPIIBmyGJkTX/XVTM08FAlFpeW9DR1
cfaFbz8rkLm64rafFcWZpU51wmRjIDdYv0xxYcWjq9+yzOkfl0Yc25e6bUGn287kFEdZj904/6cP
Ll1GXXtpR25QteOyHP50S0XZKReHhK0aFHqidGDiojr8+VdU1u5vTi7UoBwDBUmYwzPkrZYjfXaH
xve6EjTHJ29ZYqYr5VN6bJ5U7Ebpa+hwQhIxIaKTVzBNjuVRwWLKgsbizo4/zVlXVBJ0CjUcO8OH
vFxWFMgRNBxqJ69iRBB8a7lrgczg2QOP/sAtGNQsxGMWRz1mcDl0N/fFaLmKd6fVWnC6R+sOYuWI
oHbJcebIH+VNBxbMUyx4mQCwYa/kTaatui/sVJJlzD+f9cUeDUVwA6F0aa2+g1ufnGwKGyDhPC8V
7J0ZMYPl2UaRy0onfCeS0eOcWib1yBk/G5UPrdkcPWLr54Z9qQYqK++W4vP/To5IH2Vyhy12ntEc
6KaLXKS5TwNXLKq5fi74C+fGrx/xKrbl9GMpkZkommSflNsBXlKCXjwrNPi3OzD4etTlEb1Sotyi
m1C+u34QhT53AMVI7Zv6gNwUIVFr4sO6gmIc++zNcM0JzkkKw8JTMNDd+JfZyAthTW2e6TMn7DD7
bRDdBpHmpFLT2Fxg6CIOYNfagiXj9N1XFoSS1MzpNo0AvwsR0GVM48BwgqjJ+dsWMNLjJq0jcRdK
hvJlPnkEpzj+LSil40uZ7AM+uofV8wV8REj2oLmg5apEfQ5DeQdL2jtcPdlhTb3RUphprqiSe9rR
Oqyqh+OuOqTSejSAa+GGpiFklTYGO+f88KpR8QnmDOQSrfDZDtXUI0q6tCWIDKSAIEtQ8WdW8/Zo
RWuZG7jleo/do5sO8lOMS5QsBZLO8aSKxiWyLGkyO1Gy+heFdV0efSq8GCnkl4XYvfUALbVTa97G
03VGOrKxQQCI1KWMLoovs2PjyVc9MA3yx0j2lB+MXYkv9MNsQxd8lY06tMD3KDn/iN9i3bPZ9Cl0
2XobbnQCXOxyId1aZBkSO5oxEWxL8u5gyYyJuHJ7bx6NO5GlIlyPYSh/ivyQNAaQpIqpIXKglqHI
vzs+pcf/0JZHMcwIIUNjHayh6FBbM47h4iOoiiGKHdrU//kNeiShWhKLS7KnERFWp/VIz7+geiD6
fl6vaLpJKH/A4YMuMBUlvOx+2zC7a18eWkiYI4TRyKtFENOqH8YDMnbBOUec7lD/C6Ql2bFoOzj4
Ss6vrtFHwNYn6vDn+S5aTTYzZ1mzMSIC/UabwhqQQMC5Qd45D6dqsPIo/RTC3r9r0dfpxhmiYfS4
f/OJ1k4dB8ZJ2oJ3zaCeSR29ShoHauHcOUo58v8TSSwMQkE9B07i3Tpk6CK/iGVDXtWkvsfC7IbW
/SV7aya8l7zpFYFWSHlG1TiHdV5UddmwFUJHb/7LRC0iyX68YbkylALsbJxwW8B/vLWWdmaj+cEC
tyGKxTOx3K+HILaGXkIKhKAjijcQLRc0dyMkRhJvL4dDs8FV3muZH4UB98y1+xFdayHkXtamkhNA
Yb2lkQ3EWxKiguPAEnx1dTmWPknxODBrImf8MZrGtJl5bRQ2S1/iALfWK7p9PgbFldYQCG46VbUS
LMN6wyBrNIHxnX/mZOLcfPGLnfntyR0lM0uP4LiE1Zr4JwhzRpHcewFOsog2QMsKJJy4NfPwPBvT
LpshK8eFAhm2THImUXPuZhd2J5g4lAqtOcpW2bXuc0xZ23cEASRvvTQbG/T6GNeTURccr5FKPWkJ
NMGZglQTkW3ib9gGCXN98aSjj8bZ9AVEVgNsGcX+CFyNV41mLABrSZ2NBhM7fv+xTyHlE+nI0H+Q
kKGiS6eS4p9IIz/ssMeYsQNrAtQWlZ1vj09ApYVDO/zDvWrqcrsBb7IilYGOgmhUl/OTA08FFOxT
7QrpD9MG9+xkO7mQaBa/1sbX28g5mXB1RoSSahfOOpwtoaEDGoW6R6WRVuDCX8r3TcoLWae0Vh/r
gvHnWr8GZBFoQEeqBIWUa730DVl3B2YQIj1e3RNxRlBlnFyres5RMFMpFEpErbLF1P+czO9Ql3fs
GuWpsYPipw5bEVk5mdqUlHjj1Lk5MN9ELU2K9r/z50E/HoE98drvwihJ1RyEWlmBJOcvnGxGjkn+
PIji5iY+OeYZ4n1bJycfk4LVOkhdxjZDC/X12crXUhuXvgHGSVvI8fnRxepB+p/4S8W3hi2Uqf0j
BuBb+507MO94Dts5r9P9yx3+NXACWpAFVrxauimUxokYolUKgo2okQ7Osi2wSV28wvmu4vtlyP/q
w1WgZCkX84vB7YiuaIvaKPBivOgY1wBoCwIOL6xET3P8KLj1946RsK9NRCZUvJKGLlhmEcKe3JVF
hnVUpP4veeiFnS+RmxaPQsZK2/xsCBGAA/MoP6GTpD+icXOQrotAY/vQuqA3KWHqMeR150F/fe3Y
NZ0KhDk5/L9Xt3N4ypkTAxdktWLZ/bJDN1aiVZClpa1C3GJFkB3CFyhyg/WOqMItVNU18fuQNMYT
PvU/5XDPizfWLQzjCh3fKP+VDrI7KsPifrFHUV78ogk2exK34WVgLkJPvEuFs7IsLiqBNBN153Zj
ZEFO0xKiihnMsHkQHV2iYvyqgwnXoHu9cv/7SDcJ6SGqOBwxBE5TVT8luqVhT9/8om/yws7wgT3m
pY+YvnhwYF8VjNuUl2HdLIG2L+/qBKtCTlSwFkAXQjm8A7VdMtJubJzUaoO5jmidzCdsBq1q277z
QNZ44xOuKk0ny5T1rnjMTTn7zOeoJuSEL271DmteFNJRiQ8Ery+8lssr+shEmjnOPq8zDCQLz3df
aKOvFTRbnhMKSxwy+EHjY3PQnKCw6qFLeM1/yuFnnxpUdjqGqoBlm2mmxI9f5G3xkw5Aii3pD4ff
sQ4+uG2iH8a/Noh9eUuFY4sXIzvZ+FpgIeQptqEhXEyyeHXqqTcvrEK3zl2Uv3ly5qxWEbuoMDB/
/dAB2TQsySFlGXjMKhgbokBNYzJpM9GYWKVwgPBxjhwPiVf16qSd8T/5N8zpQhU+BUYbFQC0LVBl
xuY1Gs39na0ybbJ4Qc7MHtmYbGaOVVukfKxVHqlljhyworlqftubFTTyxafFdVLE6Hh7DxWzPpPb
QCS2qybhK2/yuqabJBlGWNTuUAqJxZ00kUG7B4OPTynT2B8N/iUJgmPi6pS8zBzWP6ALQ+D9dQi+
qWCz+/3jjtdGEzVLD7jTaOMTQUKP3xS/g61Oud8hUuXMI4Khxby4YTjQIn4nfKhDOKZgTWsO9YjF
hcnAcpHcGxJTJBPOmnt0jBaJa5Ke+NkgqyrYfpNx9MC2A49KbOOZS0soYQ9MPHFGYvRWSSHMZWNd
MCtN7lT5Lv9D3G6zzSTzFrgQk2/BgfYdNqdGJYEhM9Vn12UkhtJjcmroGAtVN45XXb7XYx5tlyT8
9X9h7l7H1U12WGWtszOqa/KWXEMsulA08/V50bwEEPYfK55y7ApeGHQMt43AJqoMAfPsRsOkU9cL
zyiC5zHYN/3XjZg0NfWq11G56CDqJ1jDH2aYSW9gCEva0ODPXxLe1G/TDKTCno+XzZdj0dlWNi9B
vP1bIxKliPjxb+3CNz8ucm8OnrbUYYmNrV+cIQy9HL2eMJpy+NkAJbNjO8hQ81BUKgJ2HqWBsAWG
Ro7WuCMUHi2PyGOCIfYSvPxlKzkGxgK2ALAI3PYx/BPRnyDW7hfhvHoSTYl9U71WymcCXmbmWvOV
io/zteJrg5gzVcKbfzjM1iD/d/4LikifAeWL6pCGg6cByHliv+iwYxtD2RqMr4LrDkl7eMT4UegW
fCKtSSBPxvXUFPpuBCcbwd8ostfk8COobXIGyQddL/1jfs6FRqR1M5+OveCzIell0tSQ0DnU020u
AqcmYE2DaeJVV+6A9rsHQdB05G0iP7ceVFX33nd29ICK2iooSHk4RiOXzQpIap6Y2KipL7K4NYPb
5jnW7K0v+dMRLOnS3aLU3ajO4jp6UWljzJOjKiQEl96B2Q63jv90rhOLJe7F3Ejxq2uranb0Jm+A
Fk2d4AT/kuWhctPJIH4s+/63HjR9VP2AQgGgucLAHsOrOjlRV304Aveo/zmoulQMGGSchVKueNqk
4zTNu6M/uHGhmRB5WgvEAUuWdYMC+/m4qoaRAGXdgA01yrP2jeV1WpUdPh0QyyE+ZNjRCd3BVAiQ
wyIG5wn7YyBwmy4m+SdtHU2C4G94TvqWkeDwm8LTxM7M57V2HyQGkMJtVHBRcnEhbB7LjdHZKRis
ozxZOU6YcT5B3S8jqvimJ9p3+JWnaBXFwvS1g8VpjWSV5crkc5nkSSDMCjZJV3B81m2pmij7mWlh
rAOFLPr5ZuuoS45J+ypupqj45gLLNfOHMk3SB+BlASmF48UtR7xg2sldXr4itufUvQpDvZu3u3u/
hlIxoaHFp9lKstGldkXmurY3wKiFUc0NbKjFzOTq0vaA+rqIFbL0jvZXKAfB4UhQfzljdHB8z58Z
NNFHtUS+CE1oiZrOZwZen6vReYJ6Btx9eNjYNJoe8XgD4vX77nMhiJibHHacazDHYynxELQ6btNE
HnjZhweRbTCjw5whOdh9jRQ8PVING2iD/3udhdatFqPa09gORNta4Q+5HJIMpIIyYOkWDYo/GG1B
/uLonBFAdtQ40KA+7rRuJRhjJG3d62gvyfD5UQyfQO5iRsBkzxbtWNT64vl+74Zwbe0tZQL7iwOI
QkxmT8Fd1AYSjcAo6w8OpopIJOh4tXKfJGFCQZCPoJI6ClerIDrExXnRhcQCbLrxTnmCZseJhoAu
di6Cfg08vdsiUFJJUrwmvPeWxr3B3wRbMbD0KrvG1liJjw0dqJB16bA21JPVAxHXI9hvQ+ktUE3v
yR3w1Q2uJ9bhyVFctnCWbSgqRCmlIiMou3Ozk/oLDr/x3SEPMbdmNk+3AukoBmKja51h+ztFm/YO
2YSpom5UJYKGjQ1WhDo898YrxYJD0pC0sCm81DAgK8vIUS6UHotP6ggqcBEh5T8+LarSmk+Q+9/v
J5Ct9QlTzfqkkqX3yAz3UI3+GwPBoTdjLPo/MypQHHSdiQ2grM9xnW38/QsY7rS1WsDdPrm/+LBa
xD+cjTm46gufYfkuib02n6Uhs/SZKSjd7fRgR/aBVO9cl6+j7giLkPh2xXDqNnECJ2ejbki1eIJO
UGpBNjeYXgiOs9kZICQtw9exYVFyHoSwksYJazHJK5JjN+EYICe2V2dbVe3eyAj+C7uS/t+o9EIY
izXK1Qk187bJAADrOczpiTRU+Ogg6UNbrx9ySi+R2qL4oJyCKtEEDCsITSLaMedG7YKs0iWQXOOh
184cJxVFE7LD+oAp2/46yeUoXPbRTYdx8kjKmJ70KmaYL3LnCl/P083SLhIV3WQrU8J6sPEWklPv
iDwOWEWrTFvhjH5JiXHDUhmB9z6dqm3ayVEoTj7Ci024GWwV8p9PKap7SyYotdMaHP47G1jPlOMx
M31H3zkYNgH7sF2G87M7K+keyFW0NSx5THghmYkvgDGdb16ZW0huXrm4ywADGVZFt8+iDfXFPnbq
AILdOWdERzQCPMmgCZS26KYzAjW7gzy+tlf3eAop99z2e7kjeSWbZyEXAfufhgPfCWC/mdd+tgna
ZYPWtxSKM1jizzHrf7SpQs8gDqphlVfn4Cyvgzgdb9MUmOEw9JrehzU/9nZL1cl18xcMfl3whBr5
vxVgfKyooqJZ/PLrmMR8pIMOPoi5F5ARuSECry3X/o3HQmKvAD5jLTbz8gSGn2mo8nwVMgzPnAX7
vLCudCDsjqjAF1TEnSlgNSyIN5rduta/MCukuT9FnKsEr7V9amgP1mkGRnz39U8MutVck6VhEweb
z3iuNllENG87ABTgAZyk8j/l/g4cJh+rkbav6V7NoqhMb89HHADJdUFeJiYOBoxWBLQrZCS2Rwqx
ycwKTUVOo/R1FLJPI9yckiK7n7qvvjsnftEw77qPSDBpPeLgE6r81EgfquQWwHBiR1L6CSL4k3hV
REzzcESorcD6UqgM2DryeH9JW5/iqJQSOE/oqVbTeL1Z22WF6JPPIGDGjkgx89iWppyTLj0ZtVLx
S4f119Y5sDAStwhGqePH6GLFNFtDUE+gxgzTw7ShCm/l9UPQN8qmZtopUuTTWac0G/G9zHsLp6eW
dviOHcE6bTC2OEs4yViDoCFkoWrM5GAZuN7We8LT3kD1TsiQXQ+5TMIEKVxKcovmXz5bQuQs8YAk
fMRI1+hw3kMwvfW5kgVlBYP8w+Zm6NDcCqsNZDIoww6puhBGJs6iw0BYa7CV0xFg0uVfRdKdy3qF
xWEsRN7oUX4TYgnlA8I1ZTapYG5KA16dUSVp7Xzu0ZpRqhaPzlCFT4zfB819oIFwF0nm/ViNPvX1
wqWC2P5r8dZC0cy2GyD3afOEFROfCgv4WuFj8zOhXueyPZXsqTYL42bLiJE+aiblhNMEx8ndsZQJ
Hng63NuVQw0sxogXr8CR6o4S0HW+srEbN4/kGRd/453tATj3aXibOwE0VDdrN46Wujhi0beSeDhI
Z94t+T88USP1YzcdNmgaI/tO49lu9K7c0vSuSYZNlNO2QTlDWMkgjDwTu+l41kLD5oUTK58eJNWL
TGG6VJNyo36nmwGvzjNMuyea72Cgelw9G9nO08u2c/7Aepv6jVsgc8nQZsXtqTVrBFrNLYAAhJsL
ZAfV9+3LAAWClN+qp7p4+lGdl//ZWgF5lb4KHhXgnWabY0at6DP1dKTqupgknhrhP07GswLWzBrm
TESyw3lJw7oRr521hZwzFXgYmt6GNhr0ULRQpJ5z+puHGQw7UQB4KjcLYx0U8kKk7OXxig7ukPxo
IYebp+/A2SZISasaVLDS/6wgjV+5RG8d5vzHGicT3ZlkLm9n59Dbufw6z7WSzYAfpxs/XUzXj4ng
OwXo3Yr9WSUIKrFwN4WtFRzD2CnSR9lO4W4lvzSWVzfYyOfB/japqDZ3pAk88oWW3HDjjvYSMce0
ksylbrcxqw9zzDnHoovwbEQT9+4wmmsuKwZHPgtlGmkVjId+9GjwlnXX3gQ9UaTNwN8alyy0FFyw
rYck2xWjsPwIXOclg3aARAgRmlaakqEtg5KAjUlYVirbSyhKI9tNB6SlVN4hFjBcHJhD31n0L9Nu
FkOALntaQK/0Lu9x8dAa5M0cVSG+v7p2cimaQzvcF8Kb45613U3VmksWLSS4w7o3D81e6QqLW/Bs
tiZJceKN4n9qORDh3PWykGpKG05RR73l9tA8FSidfRA+9ipfr5AHXe0xJlVCjSgok+u+VaPqGV0k
HjKvGnHIYTblzkFotHBK98Ozgb1K9s8aEx5ekrkxcNYktX3OPMuXMtLcPaDVrCObYnwj0mS/ZeUW
oj/EIBIntwYi7b91EN2bgKcLiZXn6mQRURDUwc6DPmuSoeRBk+z0lB6r4cwucPt9w2nlx5PtN8Vk
sEGl0bvlm4YWFMblRSv3EEBjKsAdQsQAXcQFn7KV/Ll+BPIrXnBK2o1dd5ysk7IAfbdOz6H+8Ds2
ikXcKWqzMngcyegBGiDHDbaMFeXb18fgIEnkASqAyKt/xLGNXV06wGhrFFW1BZB3G13CLXkNn0O8
JYz4tasTTvWWxDwDJ5sTF+gCDyIF9OQyNGseSVP2IlJTe17ifE5tkowKFKC3mJxUV81gECUmqf6S
YpVt+w3E+usTydLRoyeei/TGVOJ++ap2NABYSKB35c4RZY0bu8vTX/qRA9o0NCFHlegsFfja+7TQ
+AUKhcP8gt0RkdcSfHC3XHf+okFRyS8mY7SRBRJYQIvMjL+hFPd3FJh4GyzfjRESgaIlBIrhjr7R
8eqIWOZU/SmCJMzUwGwK2CLoG/dmfa7LMtfNXAzxag3yg/TS0ETRh2HGzVtuCdEtvftf//vbjy6b
Kle58oFqRY7QRk1IrcaJRzG4Mhb+/7+9wHEf7ghMH2ohodzMF5GLQLbiISGCchEB+dNvM7hZyu7V
ZGo3JzMFkUHKT7LQWcDHCK/HaU1Ied+Pj2q9L7pxE/wkG24Ost0d40HAfKYrnIcZ6fLB/+cNyDaG
g4XALTryrjh4CLEJjFilcLks7M5jcS/SPpf/LxrdBvTJcSbp3FnXdWyPqdhD3NjlJGIxc8BXkJtN
GlATefRo1tz8i9Nwj/gt74pqpn49L0Uh2Ho3ROjajJN4zaJVIpDoxsEDLm9qyPrCZP60ZM84Saam
vkgrRCjawmliVTORWgNck7ha6f30oscY7dd5a3V7X5XVxI++5FCgR3R8NG9/x+Bk8iV5NfojoPiR
FC31VTMEMIUiVYuzsufHK7KKRRFmdmlsHfReqB+uZNxXXtvbcuAa0OyQFylFMpacP2KgT3cmesLd
0CryrCXJJ3SttulJozFbblIAiBG1MsBmgQFD4tD8AmQzvvAUdd9fNVaFInCZkc1zjmC9IVwO5xtC
KgjvCUua/+tWcsg/CHnaFU2NwaM/OPdH44e0K+NCslXsUPuLe+GMGFHPHsVJBTd6nUm6NQ5wqjcE
bSFqVY2sJWl+wve1Zu7lmH58n7swRyFrJJLznmdWfWRJTdM/wpdUy5IQl5s1zwn3w48K3/0ry85h
/VGkq3cTiGNQUJkdb0PsZ2Tnzz71YDrIYYGx1Z2yb70HxMHecON+VJ4N2Q4nV+79aZD8gTdN8MWa
o7iRkgsn3Ck+7HKnwdkUFij0EFupAvYJBIZwKAJRb68l8nHaUkaN0IzxCqPhTeC7IOhGHLaX7C3B
jlR2cFEoD+CQtYuTT4NBSnw9dkr8P/9zLn9shVUL7jWRM/LTQ7MuvSItaficUTNeWUyk7cFvwGKy
gMjRDzfAPNZaWx3Ycp3tayovqqt/hJ7c/nC0bgxbS89IR1MSqH4iFy6FNCfHQE462Wnt6yDZhlWZ
1EngoMo/okNhLy++j3LwtSDGB1xdl5QeXqU4kkUycLTymRtApc+slGkbk+iPrzT73J04j+ILF6CX
qcUuY5Sjak+0zOQR/HkJkwNrLaIZptMUpD5+NzUTmQKKcHcJxZ9L/ie9wuELqRBamy1SroMVsgTZ
IK1+Im2DqImn7yLapB89mDQkhjBVYzd4m9iGKP78M1CVjnIguO4Cdd4Xl/FgR6k7HdTyP2Q8wLAO
2uP8Uq9N2prTX94x3sJPD3JZRJ4+neGXSREUUyjUbXQULb0Ombox+M2O7ifAxrJjf2yGkc6ci5ZQ
MT0GiBpU1G0hLwXCrXQbjvy+JY3tY7giSwU1WF/dwCY6mY5gSZgbp37OU9bA0esIGn4WEvNldysv
kirh7F9IjyldoSzcSF46s6MTMvh+jJfL6Q17vaXNCez4GNTaGB/T8AXDFtHhcPuM4f18NKQU9/cQ
JTPUOKv59xy6QRGjNNhVj3YnoXOQb4f7+IzGJpb/WhHHJ6KbINu220Lj42x9pHdrIOwSIsVVSUET
1kvkKJG0XBGVSq0ludXDjPpT4zkksaVGJtKjJpMn4p02AioUcJ6n7E8EAo4e0SMiYjr906I78H1z
xUJ1tuCvdGfvb7PpaYrPNYed+fgulRAGe15IsbV2UfWuTS/r+t+IPhFydijATQPIoBqMk406UN8x
/MuyxR0wcxcv7pTQK8DEWHIbdgK8P5iCTJtwutFfHdLQULdWBG9v+jQy9ru11xo99i6LWh00qtHX
xnJOyrhiT4aUgGCWGRAkFJVdWhwxgDjZ6k72teWP6VNcweshYGPRnZWb2SnQ0pjqmLtMS0eMaXqg
iHiMUODu0yijIeSFwf3FgEaPymyT2xjNUNVTvetezPQWaRFmzkXypV9R59Pmu/zo5OwDQpQIIQMR
wogenhLnXVbLyddAfrtX7eviKlWTwZBbjpwMjz5nSBHziW+T1wYdX84ROgstxSD9G3QQnMHgxi3c
wIcQPS/V5SezJaM25T6SPsr6mrc6HdAZbsxeP5PwKpAYlX0eiXnefF4a4OzqiUMkf+kG8EKdH1r3
fTYL6skwGZMSqCSH45E5niMb28lVV/TRO/G8zSi5Mq2T6LGup1rSSa6CSy+zZaVTtA0XmK3H7G6N
/ZONxdSo76AfxVgIH0r8kE1dOBzK9vQEZ4L6If70/uW0/0YEJ7NFI93mKOQN+DDa1uMuJbvjOV5W
RLmHtMmBw4SDZ8U6SCQ1NL10jiDKmdm5dBWyBzzUnuayVDHuTwbxvw9HQFktyF+2EoytTYCoRP02
rt5Ui1lf2eobqmOgVjjvKR4xljsATlOLGyNwKx1NHnC8K2UYlvt7zd000XOCkRlUQjTr2xn9QB2u
sHfrJpoyIyrQxI+unayZmaDcfJn4iMq4R83cjpi0P1Co0X35uHejRLvJLTWaeeoIzdJeq97EEqpY
+v+DUuRtP+ZdEUDNXplt7mP5oUIXy0PGAwllhmEn34ra7JW3Vyz9qThDecPm8MCUF/a8Hyl91hml
NXwdKaVrI2811XWN0kOXl3dOeuozRlOtoXBLYzSxnvMbgS7zSFskjfs0u2FWCt0dkA0/0fFaFLBF
NtZikj0D8m8xMHPZOP7RD0nXxN5aPlnnRKDHvkDItV9W3AcrnSbgs6YDWHn4r5xuIifB7RWfuAQn
wZNI6AcVJDP3z9j/ugpbFWG3Oj5+tkkha+Q9+dnq6xGNOm8eEWqr6XZrbcWTenyICe05RkKbzqTV
6AJBegM/QMtIk/ZzCmOPrD4Pof6R7OSKTDh3+iANW7m2A/8SLVHock4WMzgYAhOwoWSvI2rlm0Pd
7jT7hkX65TqQoLr9N3dlMyhVqvTVm8zzKleGB1BMowUuCQMglrZIBQvQlM6HMtBqd3Cswu81mcY6
rgRsiqJL1gTb/LSBSYaDQRDaYcTw9SAmgezUfYt9hpu+kWIFDbl02GJtqUBz6Y1D17mlj0ztsHd5
QLf9HCFoISaNWxPhsE+3YWy05Hp3qjdp4VzYC7mwp6YLRNgmuKwTlAtVBHhaa/1nSzLtO2l5d8MT
Vx/fI1P/pheMUJCSQpqrB5i2Zuqdj2WjGTeQJSxH1ZLFQoDOkHNMn80Qt+ZwS8sAt9PuRKacxjZB
4DwOC83cr0PfZADkIfC5Gs4zsMPR2L7lg4/v+unVixcCejP1+y9s+17eWKSPDEzOrwh6lTI1Pepr
YSThax91lfhcaBXadnZ3o9shsJljS8zrpvEWYTyquAfruGGGFTeo90c14G8vpCslOC0eqUK+HkjZ
BKPZhl/UMlwpJBivq+e3m8zAbNLKlYBglDH8SAhGyjlKcVYLOeDzFmc4aodxB1TLX1OW2lnGqCQj
iCe0bsqUBVG7RNAtQueIOgT9vY21E/5XS4idFz+MMS7pjJf33MG2Si+73o+/N30QctA/odzNbmwa
uGNEXUojsG9rtqvltDUeP6DPOLDhAiLOyVAnwCxWt3RMjuQILHWY10BbjcK4GqxsT00tJvPQebtd
YNDKn0nNFTFxJxInfgcusClqs9fnsu1MjKuJf8VCWabATC1dVoYkZvvZxvtCgKt9sTrENedGtGGE
7/Yb1UaOuB9nVnwJw6/PHBfywLDw7txerfzS3ajHNhUp2Sj5DMtWP4Xgdy08Wt4SPb7VRKzKK22Y
+aSoUPzZSBCMzBX3tklVeN2p1TpV6cZoYgXNPlgOMi8Mu6ej+nsdCSz2ngw8awpwDBnnyk1Yw+X2
v9Vxslg8DmLLsI5FGNgVeK3ZnVRQtEj4Uu9XqfBv0Fk7Eie7MgwW6nhMo5BRVT3UX7i+SQ/dciwP
hLULfLYypuwRIQfvmn96b2dLefexgFFmebsOpN5SoH8ipKmEpE3EEbVDGsaBMzB14O+ZP+4CA5K8
enDTC5bjlf9Laqn/ramAN+F/LJt/MEm+h5IN8718QDNTfa+n34axkz1Kx59JLnjLMVYZvNY0H285
Ea/kd0vmSOh7tJRYzqnT3ThPuVOlbumGLRswE6lWwVmagTlwU2U5ReQiVofsmXXGuTgjYBMUYcIr
xsl2w+OlFDZtwrRlSbi8xK9Qd8lB1c+CUDOqIkA5lWb9fUKNtzBzwIMAvyqkDkhVYSshGqkzsGU8
8UhkBIWbfa1pOQ7r5X4IBx8D4nueR+/D4jrVwG9ZHTZMcAnXY/LAcP/bsgce0Fy55bYzS1He+xzx
/QHh0kdIp2K7ORkPKCjngI6ovfxKnRiconQWcVJvHOnIJ1/pFuZHcEWZtJNW+AzfxQeKQcylU/Xm
HtZMPV8KFJ/DeYtAmIybf65L5Shj5dlmgHgS8FursMKd2gTt9R5yE19JKOUrWRpwt4HwqjTxoJp9
uBD3SB+7cdF8arObiB2hQoqKkl7EiWA/qIttlctJQBjYTt18+7YI4gss/u0TVl/6O5gWq610KCR1
/B8fmt98KwDtbCLypKTHv5ZnGelvufUKHBqR7WqgpE8bU3Upurq0j5FYqsoXIge1VG0QmXzhPxn6
7GGtHi2pmtKONNLhaPWCUggGi5xWUWBCqvjJ5ig7Ea37LM9CY+U/VaumA9iHD5NGzq9jQkID5kBH
t6hXKCoWIfpfQn0DLR3QVitU5Ya6aiz7S1AeIoz+dvA9zEEejwQYWfdtDQcIBBt0TVQiKhVV1Yad
PTuztmoRBY32IvyQ0PStKV45cMy+4EP6xXhai+rHAN9D2dwrJQEvY+5N9AVtIkYSwpBhuorL2kZs
vBkFfx445zWE57fsVP64Nb9ap37sQfxViBaKmwFq2NGjAj779X7WAXotbAEcNeUz7/cvmnuJ3JvF
PfDJKnTjN/3/by5ks2nRWStEnp3ucCjCLsGr3AZAce76nk0OW5H/Eqz5MN6qSGK3Cog3GdJvWIsW
3bAdL2iUbfTRT379wMqX2kMwCUFvDy3e2r+qusol0MmghyAZ+kpE25DcRPbLH546eZV6G+NW9aLC
9wvHAB+bZnZLhII9nVbz+nyCIaHDK3Yue4VUJTan6SyLmJS7pgJjMEYvZ75ENuzEv2sakDXPZnOE
q+s0j1FJNlCt6gHmZB+qgsslxjaFk9xPv3Ld3fT08yZ8dr4de/SLOk5W5+fpl6Jci6zhGADZt8+N
HREkaVleSUEdH+MXTbg9BTncpLLD49HzlIfUNwEEIg9fV7FRIrysekv1IsQ/GaZKMeoAfcbzlxVU
DztajBBlrDxjIYGLGMuD4nbPmzveqy7Hk7+6enwYt7xSVdZ7DLTn/Unj4LSBSJ+KQ1bN9b2NklhG
HqygZPPi+k8C5KwiOVrL/zI64i7HHHMvVSgt3u7WmVDV/t6c1+jKq4VOaonQBpgV21sssA2qj6rw
BLEubkD1lHWb78xt1UlDVVfSTKJ9UoRw9rXk3C7boYrbp1KSg/w/KTDlXYQZcl42xj5Ax3KMJoeR
KMSQrlH1SXcckf6o/lWBlDs1/dVCp7VcN6WuwNXiflpT6KZQNxWG56co6tQRz5ZUg/AC0+LBolmM
pfdHrWfprZEJgzXxSizPejcAgIJeaviYW1Onrpko8j+LZ1sMdu1Aqgp7bApxLI2DlKfhU3jWaFrg
t9fmf5iUl/fXtlAG1LUnFREZfDwo8DZMHTEiQYz57pO4JL9LARoeDA1PX2OTG0q0/+/G2+LYUYnp
fkvJoVdliRpTk06jr+Tb+smdjfURgdCV2MmegS6XSW6qIEFlr69bBH1yy9sL5bfzsYIhQ8sviafC
OD4fy3Bjk7tqtOb32ia+To8h2o+WIPV7OkbTcPEV2pSzENOP+vMl184aaDdqwstNLnWAhnQbiK6l
pSWWJ032jwK7J+8BW8Xzz1l2sm3vyMFiIuSv6bhYqGyo+FesIRi3tCgFMtQQElZCBd2OpnC2sK4P
ks660SoVqGa/2T5w8R7o2R4v08OugDxRGRP27fzGKXrekPANOidWdCDvcrqm9KQOUKkVJIgZVf1e
yc0hUicPQkZ23NhM2sfqvzfY9ddiSiuIxrw2ucAqwWk88vTubj+t93Trd1ONBL8zzpHQFhywOS7K
8nzFVArEI+ELmTQryzLG+KOKMqYVEKxKhk8wCtN2KrSDApto4hdaOgDTp2+JCOgMoTnjt+2op2X2
KvxY8lM3r2xAWb44JE1n9u+xKSIPTGuGjvrpsQCi8K86Ow9GGDQD/3ym6gfKt/2MjWX383nJQ3Oz
8QXKE8z96melJ466knYaj0+Mh+ze60uB3CReknw3fsqc+l3dT/ruZjDN6pWjIZAEy+Ws1seQKGm8
Q27/kKpwheiXdJpZbfBD2CLfAwi9YA2w+O9VgcXYobTRp633LQm/z4P6Zp3C/qEwZ8L6eNnQ958D
tnd1Z40q/oD6lcdSGfJjJfX5TekL/KspfuSOdN9WiXOfL2sAGUzM53WTHvIdjkQj/hBnRYRwVMhP
Y7FUYeNoBPazzu4xeIk6EsxUuxDowANOoyjf6fbWcz5lNnZDkmZTq+V8PhZRHuvq4Z79MqWc7AGj
f1iywx0uVqrYrCK0msxs3jMha8bMWyqIi5YFH9NWFhVZt576ROjpliz/SPVAjAVTPuCdnjT+cgca
G7VTqz90uwsPqDYTWKAuLQmMN0jSLLu72+/QSqmKRAJP89igf1FUZG2NXEiZXT+6zEvs7sV37kn4
/Ca4WH0Hh6vIcUf1niKaBRjMi3CiQRVzmKxugyVURv0NJi2932CJQxO3B9wEYhWR78xpbL/E9h7q
xxJXhGGXLMnFTP4mienCFNTPs1yCj08Zub5zLFjTfo6Ii6UD5R/8pFXfQ7CGYojARj9pHc572bQK
1UpD9gaq8xtxWp+0PAmLb6IkLwQEPE27kW5w7HmzOagr3Chz028wT/ITfTpK/5gJq/3whukcqWCc
xV6bokjVAK9LDUbueFZCa+vdefV5yP9c+fbeP71M2t/w0N4NleR/T3w1isJnjQmfYq9z5C0kn6N0
01Jcy2fBJjsIcwavu7jBrnUDSG93JyNFxULv4YyBrs9t0LsvWNHX0DsmUHr0JjwpOgCXxBpEV2eQ
kypA282PxHkMpZruV0fQ8UOmtf5NDRX+tANw2ARhS/dD5nI5ZILkCVAGxPCJIj3/Col8X3DgGdAS
KBu9+stgPa6z23hJKSYGByIq5ScCheMKgxKoBMBc94Rq2nrs2w7y7cc2ucj4M2oiSHKMa/zNOnwn
TFlmOcvy33TZCxQXnR5xrs2eYgbYojTno8EPGESoTnYsKv3CPHLrkZ0GiskTBmyU6QY0cyw0X4p2
borT+vxClqOT9d/igmamh883tB+KK2KwghPTqKN9CidrFTS1ev/8YmiN73QiUbAYIjhpcllmpCrS
F0cudqiTo+sUAiykPeYqg4Cr8vLUj6key2aEeIuK9oxYVRrWrBZTJjb8a6NORzw/6fnT4ctu3/Zz
kJK40oiLzqy5wleRNW2+DpFwVZIBGbNcMIhuWFxwaoET5cRReM02DYEC+8B0abD6T0pPRD7/iNbf
Ms41Q1ZQAhxHUVQcwTBkGY/L5xW57hWcOE+hTr3ADFLytAGGSse72Ql/52MV7LXfTfn/dH5IGE7Q
T2WeA+xSfSBbd/y0Om9hUdQJFK3+UzzkMyc4aO79oCn21qot7XPYdOJqEV6TOgW+Dxf7wmooqyOu
W975fU933KuzkeBBPgO/1xV+XcEIv0S8LcHQrkF/tMru+l5NlOaa5DIpN/cHml+kVTb1D2KTd1n6
pJoaBgfYC/x3AaDkU3z5VQ2nj7DMyU3oR/bUTHqQXKqZtQ/Nqr6CPNqwYJ7y4GUE4TxJDnq13GgL
QKYN3PCrSJ62JHokvk6p5YyzQrF0hPY2j5pIsFLkCMgp2SBjYt5Vjd4R3C0bMo3nDawnhNdwZDLT
jsRCEZTB2NUJF10X9BIGs9ZABSgziLbmt+6uV4iBzNQHlgu0va9jdGdtbVmPFByLGA8FLSpBwQRd
foHdLHde1QYYHidcws8+bwu1/DrTVoPUxH0EYJN4wD4U+lyTz1tyZKSEh4IQXFjY7yg/hUGzCN04
4KnkDM01QTcXaT+YglMy305Xr8pQRhJPwU+6KDtqDkgCho4KZdtMtEwJ5ZJIvYn127qgCeEb3kaN
qkyvlvK5pES1SjLEaR/pWMXGzKznqcBWrDcigOMarO4mKEEZWbNecPSVYuhk0+58gb/VLvj6u/sd
0Bslozpoqx4UpRbhOJHf5IUHujpeU2KFABqrLAyug8aIXv+gmWO3AIuBhR+X74dA0DDRm42p2+/W
HYMVRm+jDmrzrnUzCYLNGaqC4DaDwMFpsIw5FY48C/hf8wc+MzCSydVrILGViwZGI5EsXb3QTrlI
9wUreZsZzScKfDb0wlkSQeB4aoiMbz3KS9Z8BPMz/3LaFvv73tT1hwqlaJ6kA7jqIqpISTGAnDVP
YoJX/uz9mweGeMNuEG9po7/Zuwj4TnTsIw5n/tJTaa4bi3y9cLFpMacT7M4G0v8CzMxekWahHdzi
IErT35OepAWXbCy3f5sDVafKaaRmQlb4/UuZQcVOzNaQtnZC1iAQY+1jcITuLSKRYMHkAKez+JBl
WuoexfvX/JhpJzW6gM/2siIe2PixZRdz4hOI0VFv7fGCmxG608lZAlLfG7ZRv2UmRYtqUodup+bj
tr2/JpBsP9Jnz0fhfwoczKUu8JYqbvaBjPFZWh9FQq41Takk+GL4bkL8FPzLFEmWczkgPI1fFHn7
9h0haTjczcGPdGTQGjML1Us7H7PZcARg1nkqVEUyd4IurLRAObUlmJf6NqGYhtviHBgbr7LGgPpi
Aob4UeJZCRgS3XpuA4I+gQT4Ej37sEkURfgGwJ/p+2Bm6/ZDwrsUm+kjAqqKnnk+axxlpCxBHqs6
pNflNhlbspcQ3vSvbNhjUVmx7XgNHEiKR+ezwoopmtXyYrrO3fI5DaBYrDiO5GShzeJ9pD8OCwSu
BplPWZ149SRdIltcpVAzQjzo8aE9aejD23rCQ8sB5H9KYzuIwvifNXAm+jl6P6Gd/zLZQ+NlKyCO
g9pqy43uBeD9n/WVsx/dv3mlLLNqSzLffdM+hO7BwRFbXyxb/w41aaAZlCjJd2OPG1n86dNF36qH
7cqwitRlH8UdQ+UhyAbhA0tkpd0nqjC3UVgDcrj1rKAXmW0+442JZSs7tFBDjGbx6HMZwcuppF5P
gbUWi/CuJNeQiK/lVTYKda0nwXJXn/YYLSymXjWJE/A4tksASFYmiVEB0+ZwPXjRpMfoocJLeYjU
6hTDeus8a9QGZ26r5Ox+4CJKDO3o7rCPtmBLff/k4vqex1lxN81JWC0GLq0tZ4/SlbTAcvaF6Gt8
xSoTeeKPKDpWAzEyNgXImBl8JGncyf2kQSGzPKLl+v6EHGPo8yyAlQ6nGDVx+/JKlG+PeUtCBBwC
E6h9yl9jGqS+Magk5EkfLRZ6i77NZNYmO4vY5K/qKkXaeMuQkAXND9CxlLwvo2KBrAZTSPmSy9ie
Cm090idv06SEkKCSsDGXCP20pGWKHjlvpy3S7YUIXUw8g87YXm5+sVZEHAxaFon7EvxS/pw5poXV
1bcGhii1qLvr5MxIxFyumXQYosMvagd91SxX3H06hbgLmYLHir7dYiup3RZ2+MYz4JUXBSP0T2RL
m+UoLYuslBOJKoj+9tcMCItsIczsEjyI7TmzPu+6qINV+nWlku8GDyqDrdoII9gjlZ+JU0Ks7L8L
pbJ9SAu3cy72raqERwZmXvlFYMP+aYF2y2eLDiKEso7ahX5l2Go1kn2mld3MJZmlIqMUxUIiJgL6
HcO5f0mgB5CYwNsJWDkE2tpt8DrBpocmT/m3I6kB10m7TyLSm2Jf+1XTvbL1RIN3ZNMKrYvtjT0Y
70FadVFu6QoqXe7sQusvjRXYpk6fOucBA1Di1YGveqF9hdFGha4m24xDjNXGx4mOfCvManHYHTYr
Q+7Vq9zMV7m2T9s/0AtFQaYZFAiTa3Up3JNUrtOourFluXTbMcuQCObOtk5KXL9UOzn1e9geGrpv
Swed40De63llVjYsuIR1KlNS9xhPjW3cCtzaKNg51dmgB6J1ow5tTLUWV68Ks6oSrIhZSJ9putQl
/RhIlHyz7Q9eyfhXySjXAlGfss7Do6NlVLUYv7RrbPAOEZMFPIc7V5jyunYhnzS91Tc7lok5hCAf
bQMcKkLI2bX+xPwfDTnTGs25pDg1clsFC5r7N5fKd9LLYFQ2APZVpwmP4fvhc4TKkJ42/jL2QuCz
FOw3iTbStKPiXqTcIZNqjdt2P7R3Rck/ipavZfMoC/JJPW+T+4RrOpoBNWYdF0RkG9eUeWL7joUV
Vb4TmGKN5KQDaMySJW2XlyqwlYYIi5B4DBPKqopoeYZatnGEy2QK15LzQLt7MLf7Hkzs7dO3F2u4
4ylwAmxIxnkcatdgkx+zrjfGg2eFCSQD1NKCQ4bpQ7f2OKQfqlWgj1uto7etbOa47hmD/TuQSu7C
nI7ayghr5rY4fp1iLl/xW/iraht4hUZMvR1rwJCKTWdu7R/BW9oEZcYQGvErnXFdSHC3W6iWXJr2
fVDHeJoq4cwgL7wiyekkvQhq1JBsSSmf9gowgO0PWmJLEVDT24ehw/m4xmxrvS4NYW3Ni4RoSSAj
4yeWoi/vVqWsPMSj+w+BZfXLPnbDaC2+eOr98YHHC7lzss/Xu6CjkkKrNQ70xKgaRJGxPGJ8tbDM
QWXHQuirJq27jYSD8Mv0XDsAdoCi+XaoYjAL//0+mc3BHFdNG5rTJ4mtf2Bslg/EcLp8pISFlBx+
58ShfmS2R9EiqGlIBRprtZEObLdzqBE7GYrldnPFmrQaPUr70gTphWmkwic4ZCB51dSc6+6Zyuty
aY3dxDpA/WLZS021A3yeD3K44NRYuK7Uijt6jhwabvhL1/E2pe+daOZ9dbgKpePJDJV+ZqiUtS/8
1nD3vit3529gJ8ZTtesxXcVoswKkyy2kShk5Bs4ALR6MCF6G+QJkrU6aC9f/DNTCTURw16T1pJbW
BX6IKzZqv0Pa3j3TMuqCgYrHTdu0PQox/FoH/ZKcjGL4smSS0vfDIIT4oxcV3/dIG+F4O012YorL
+2LFo7Cdk39qiLksh+NmPLNuVmnxiiDjvbS07L3mTSRodiSSQipNP6T6nculzvUBMQxHnmmS8X3b
XkS+9dKeV3TDch03r+VeUqHreyWP6w9XAaAzTTX4+Zh3244eRrq8tr3USwnxfugFUeUlaIm069/a
qDffDIofm+zFlct5lzyMz7EUd5AK4gqSg0I4AhXabRu3xspJjS8VGyHox4pIiLgbqBkiZeVYHEao
Pe6D7F3ZdsMlZXO6GZ4OUNyv3zFbh+gzInWnpxa1MBgZfWqyBKFIiGcqx55E59NcYMh+2LFs5W8e
ZR+nivJa6A0puZWPXDQitxMlQDerLSCwy77/oAdwy8sSqN+avnrPyPY0AvxlsRjA6NrD3rOf7iUy
QaA+JA2/MIfHv4ARBtqw8JCwEJzP39PQOomd67ObloCfcwxx4GfVyK63b4jR0CQ9qDkYjBomQbMO
DJYJjxKDWCbsZQE+O2PUdlFL2T004kfRlZ0BL9jZGtOpgEN9pgX043bHnnqAQlOB6mmwwEq2nrL7
bxAjiK11InukNQCT2ulZw6SVCVKNfVBTs5PSgRFbGFG4Ti0oe+oVBsyBQgTy9/82WbhhMERjQbLs
YfJ+XUC5jsygwndhG0mwQVKFstgh+67YI3XQOkOCqNFgy+ELCxp/gbg7ej/DaeZArV2yvDVoFACh
jRk1udQqxFN4B48/P+Y+G/jHNU4Lea6DZZJmMhngoTwhzs6kLcwm0HO4DJh29EaK0APrFask8hBm
q7FFe4id2eLI9tUFhJlDMIPKIbLYMF66UpWkfrF3G8CvjGQE4c7txgNug0XCvDbgAgriAwjxM4Cm
0KvPT5NyAUG8LZ7OQAIA+MgXI2iEBAbYPnk7UDfO1PDpn7CGzZ0H0pRvE0DCIIor9RG5F6jce3Ie
irRqszsOSPkJQB+J3G1/ffauYso+9qEFS7mqP0rPai8H9MDq8N+IySirBH1ZiF23Fom70Cbd93fA
ZhWZwG1+iiaEGS6Y4FnxrWvXuMDD7H7OMWasfq99uhW7XgBDys4WLmBqoEeXnhghi7xlrxMIDu/m
nwkrmt3od/xURHQhXY+IhCi8FADFC7IH84J0Xj7MLDQYH9roHurHfBTl6i5K3OYjc+kEYFNCc2xK
JFJgOEqsN+8J7on/XjKh4tYjg9ek0wJqaZDGGef71UfbP7Xu/tqgL4/elTzpaHYd3krGhSTpOOpy
24tsGDiTgyOsAlS0gEju1FF3Ch6nAU2ivk8Qw1QA3+Bp9hADHh5VdGEGqHqB9EsJidXAcujh6+x0
IieDv2sN0mi7DJcoKc6P9b77NFrEi1eXA2G2U3WelVH3l2yd/kcjLiphKObp/4l307mSSVeWAaJs
1/y6ch+pM1Fm0lyKNfp3vJErj2YDjQcTAflqMAP3IRrrIuKhCL9TBJNGcJhLQGLS3WHQF/6cmi7/
OcKcndxt0YBP99HefId0WPZkJ0TczrcNAjW5sGrulJhaIcbqz4AyjsNgswiLG12BRzrQJpKj3nJY
JmBqYbZni28qp0OC/NnjBdKPa8HdVyKUpx0r2oQUCEkWClnRS65EG4NtXjYo1mmbK87aKlIVTt5s
XU1Vof2uK8SRfuq5zMO3JF9tQs2KWnDm8VjZGyoXIcOf2wvNiSPVmyaLtBNxyNs87OvqcfjRBpYd
7TFbpYYDXyEnrW53kyAehBatBHlSbX9HYtV2mdwZsu6Quxr4K77O4XsPuEwo74Rojjk6kVByi53Y
jQza2DxqsARrq23XpE0RWGl0cs7bEpR2GErz/p5MpuMQPpddwScJkV64BQOHeK1/vtKLxS03zRNq
bGVO1AOjPUFUlxIf3x38DxFyNUmlh8dbK/EJkDdQ3GP8dEiyH4TRGo6QuewXUe/mEBPa41RQj87q
HrrDkP04AgPO1cvDoZIm2ELHy0p7E1HhXdXD9tznqzBId5mU0UXikBN8AMOacWeGlxuv7YAG6hHh
VGdCcV8YNiryL6p7Yo1nmudbV4ncq/+4QluyZHfq4wCijit27JQ6GaFG6HxGCVLuHHRPOb4x9Qfh
gGtlv8w23C0czonRG2+lvuxM95LpmcTuZdxDt2ffyO1LhsBt5rFjLR4CI9B4im+0QXcNfOJcNsv7
nv2uZYL5jM2pIL0+WARg5kHLsdRHIq85DcHQDDbR0sUAnpDPpp5QJhgnRRJXaotJHtHle+jfe170
/NH5K479rcQmA5dmS/4/y8tWkmt6L0DpHOnjoqdRQlhGE11b6kwQYKGC+Wrer22IN+Iei1ixnrUs
EN9/fjWYmglRBq9kaT9n83VW0ooXChg6ofRRXEaWd8ci67TxpvvfDaZTipTGsWNVrjxf6AZMs61l
zHZLZia8q9qkXqHfVspmYCmlgN0CVJ5+iFy/JqZ9dzxeluE0Jn4cogjZtnshQwYvpD4rgP3Ti6h7
2lpzHBU+eL+wOhvTWLLyiUo4JepZy23+Vg4wdbIb5bHCUx+nAUDj0QN5vHqZ8xKaUrwOZdGMtxlV
ttN8ncjBgZD7e0wKwASBkUUOPs0KjJEgWOxTnS/Z9YaKkeahZD6YGwq1ux1Lz23Nt57sl1x5tQtV
i780964fRPe6/9KAHaPGPezr6/UYUIRFY8FAf7CykfsvW95Xofx9T0uULADtuS/tbkj8WS0Drwz7
5xGXHZWrO7vi3HLGa2/mFNK8frvKZxJNfSREu1NEHTG+rZtNwUh6TQ1gC/ehYFrwB4DsMecNi60W
pwn+JgoP6kwXHk2G9N6uKsAlxsqOOkd+rtEmUgbkoeDb0funPowTD0jB8dAZi92fQM8aEiiZtndT
eNLgC98qdUgqXqHJlxZpts3AuUqePGhzaRHApYkTsEV7SK3cHw/SHYooc6zUNeoI1R2lkPzdEEon
dAivIG9K3S81k+QqHRNo4Cxr9YPdZwtCLqPA5fmO2P07LwBGZTVfWeFhM75Pq1S429SBWlTRGEdv
x10xyta+XKYzd8qap2e0ipu+J3BQwa2+iTGm5GckMSr8EmE6h+7LRQUFAeXK4psnCIqajP7JxDID
ePyo+Gq5G80w2H7uv/pTQOBe5RBrc0mihqyX4lfb7VsU4wCSQquHRMvazBCHZugsw8Bvm8L4dmfo
wFxFL+eGh9YnoGn9K0u4X9Ah7i92tVf564jleOyjUD4+lA59e2unKwWWUaEGGTwkLH1X9L3Y4eqv
MfDGjtOjQP99Aydom30H7ZRcRyjew6YIFKRXLqln7rYZz1BVL0kB0YcFPW4wvlr6eF2p6qwyMZZq
qcIK9vyaCYvzaClkYBEmWjBK99vM6ACD4HGCohHIC7oTrbcspGLv566L5zzf8QA3fZ5QE4EMe0Iw
3feNtLWooxHyidQYD+HXBdJTlQcXBtI7z9o+60bLAdvyNlrxavoOBEtreDHQqII8HgHb3vEMGn03
Kx2lcxYF4QtrwqUEftvAah2WIpTL4S/dQ/miuR1t4JzNuD53h6I3wgI56IH7LjX5s3/1zS36rNPy
8n76BC2gpToNw4HT1VQ3nCil3oZFls4R69XalQiw0R+2dkNNIBmVTgdD9MAl3B2huHBUC4bEfAZ0
7u4dPrGDdeA91BvCWi3U2If1D39d7oHAAr0hJ6ETkX8sNGgzJPNXBI75N7KBlAEgee/QomH5XRyu
1JTVyHtfE12Rg1DVv51+erUJXFrt4ayIKJIDb0OLIQiKFFq1rv4tL5PfkUUHUvDoEgOqpA9WJYtE
wkx3CZRd0735Hx0b93PMw/AKShIn4y5PAHWHdriJZAcJuGmAPp7osasjQmWBzxriTLL5XOgOLZn9
va+1331TVODq15oTmAVeU1gi4sRkNrNyKCx4+LP7fPBSfxYC4G3CRbhiFZynIK3BIK0qRbZsGcnI
t8ZeOqmnR9pCEctVQppVCHlSKww2uFZTncIEd7SHBKkkd8uTLRtFaN/L6fM8JGCSmc67y3Ndbgro
J6r6dV/4gTL2fO6iNgY/4/9aVgqeNVjNeKAGC+QJzeWw/xyAOQ/kPCTTlo+ZgfO77knBXAC8vwtA
nWabDta/JwOPg6nunPa4LnBsUU7wMmpRtA3tG+MpITgm+qgqODB2neYwrZSjaComumf1KyvdHqDO
mpwXKIQYb6otZTAB7fyY4Mxl6j4qBWPgNK6OLIODp6OMpJAw1Ad2dqsBumnnQ2fdFTuSEhTpE4we
x6jkqaIIsxgWNjgs0WrEiWwnfo8gAEj51ixEE0i7CCnQrv+ye2+IzCy9VW7o/X+q2yq8bRLN9WUN
ubOIFV60Q3O61fD9aeckyxR/UFY9w2goCOl8Mph/WDq/nw/IomMdccCcTRK+y6ANMSwcZy2y+NGN
vxSBV+OU3WfKSEFqz/UN0Ah619W8WeVg/Dt5ErdEMQVTJhL4YrVny8MUPWsuOhC01Lu9+KXzXBCF
63xtTTl6K5iJO1aCzal42eH1hvR1cOPn34Inj3hWcOi3WQsMNjuXjng9VoLas02cdmgmf4o3OmPq
kDnbtP4ojtwzD5U0sKkCmjzzO9KFOndFh8C6z34CUmmRBgdumDbuSfA9SEwEXo20SEIX6BQDjTDG
6inZn+iQEpJsyFbGL4rC/6PuEyodd7Jnti6cfiWaYGHA950bKgPA7Yh2NJijYeRIwRradFqx6y8F
8Fxx50ztYV3bC2h33bv4OxGwtNnMMsiSjt8Yr6xy1iPtPp7I3WCIbb2KwJnFbQy8Er67FOFmhc+N
QVJwEFpr3GfzFlpflYW1Fp4m/u+0PuGlCR0IOWfCfk5FVMikjmcC5oYxeKTpNnnQR2ngp/LLL7wO
QI8OIi9dqaXyYXvaRy1MaWAlirraKLu5NdWZJUGCLTXDT17y3QJx7NMSn8iiNNOUGZKxfQar2HkN
bnkvs11vTokc84584k1nxW2Sxazg8pKwcreE5zCZl6U8pomgJ52DtvKPfqPSJZUuJwZHrs4LTqAL
C3UDcaSt+AHm1laGvsXJZaxI+uiNlobjYkvUaELxA8RrHuqyiho0pc2jKWLP/Xfhr5kfpDY1cIgm
EFh7bR/k7bR7E0dCaaV1BXdPxkttzJ5keWA9ap3okmMxc5G/DTDj7R/il8dT3uLyD3wN087QSRcg
bh4nmCzfa7msBswBcvVXwzletqtpFp4JNumW6sl2utPORJIG9X3R8AlWOTRh5EH9n/eCyXQ6HmqE
GiCGkz/QId6j7jOeCley8bmJVWaSmTkY91NrSEDMw+D6Qs/67CgtUfAVPH0fA9s6QUGnFOIAOz1f
7XHQFWUrxPdnIyxmTsjvu1wjaTsnrwygbDnwuIVRq3JA60BrhycbZKZjm4j/NGwg3JWKH+krn2Sn
xn06JvR6UnZAon9kDO0immqt0XJzlwMoSS67xOOzCOGW4pFsYStp01gbjDFBPs+H17mVDu3hFQG+
uDWkgj8/7KIfSQKwQ2MWxyhG0FjaQmwf2E42RDlU885UUNXbfsrW30AhQUB3NUYm/jKalRcMEtcU
oKJHpiQMnCti66cSkmrplM7IWXq1y/8jOrtRId84xmJ2dqbsLJ1FH1XeSnjNtqlXK9QDBfbDvuxt
vIVMCjywfHpxP1qXgYFNI+680U8A9zBLAwGnsk+JQOLlKaP0nAyRWnis9P/B2UNNmtfiyDZ4nbPt
FDb7OaEaCsoIWFs+edJjjDfLzT5BpFnJu+AkQ6Wipblc/nwmK4xJPsvPkfnKvKXx+nJXaIEUHLnB
BVRpqkKkfQBgEZnwHvKlPvWbmqGMg6ET6DFEKK80XwLhTVVTuVv9MKwv4nr8DoqODUE3mVPuGvU+
rpSSxPmCiaoO3Odl/nScWHLVgDALXFy2ObXv1C77PYIwzxCzboLnZ+RnhAb1qGOXE4jg/M0ke0ae
fZjBVKLB1uBUBBV3XRUg3SnJIICzFOkX2QLY1ugjfFz+2Dhyz5iF+nMurJ36BgnHwplmChDRvzuS
VwqI8A4DwlPCGeiBt3xuoLbacBUL9+9DUTTn5BU1hk+KkyKWrBDn+O3NXRA8uPD2+YtLTrM/ugzc
6O/K++h+F6sGsWwbHb4JEjKZppYkJ2WQqHkV3PvckKpp/EWbDnKxtOxTCSXGMsihyoC8UQA7OOFH
4T9H+SX5LMLMHIz2/L1qH0j0R70I1MzbP48/98aOXt9hsLWgzjBMFB6Ijm9ZrAQZ676HFO6cP80x
R6De1wTcmqE8YeyfDBuzkZjQGGlEk3tvUBN6iMuLm3e7QI59P+NZRz19L5DvcnN54aU1enwFW5Uh
Vc+qOu9t1SP6+lAf/01z1hQTxIg9GnkMfHcQA+Excyu+ZjCUcXjD/TFCL8YPqRt+emqGCWW6Ea7n
sECNNCtfuWfvs7dURciP3g/nNVEtKOtzOltbfYK14X7B6ZD20MXovssjDFCni5nDf8wRlWmSqPMr
kW2KzpmypubGOsew7JjdZ7IkDFbG4WCT3WIXdHa24OiTdcpOqoy7galczNc/nU6+r+RnVPALEcYH
7mIb1KFwsduQzPzDU5EYep1ZlAOptlVdtb5jh1xHTsRcoq7Mynp8z7Z02owZc8cNRf7o5LtLocam
tnCCY1CAuK2fEgw/PDmYCbPR2d9iNCoiPPq82XL+DpV3O9AM9faW+TTmCa8HwKPuUAepsi3ixbey
sD/nG7v2HBRgFVsE37kY+rP9K7fVW1zCeK7Mw3hTta9v28iaRADgp5eeIKcaazFtA7FwTe0yHOeL
dt3ONCyNRIzBSAnqVfEf3hp27Akge5/zcZ8Of/1hOjDvzBpIX6OlV/9lS5vEO/RTXiPnkb66hLRl
X93b2LCjpnlQ7FNZ+zMgAywpoKDftpYCjpdRsksHSGpozGVq1z8f4MQ8tb2qcHLuMTwQzU7hfXgO
VUS40CaJgnmZZ+Bctr3wXQkjcy5JEXpg9G0q4AgmzZPU4BJLBVWtsLVNjBvPY5eUwvVevNILcwrZ
sbjNiDAie7E5ov3aCQ+Clz3MTyuNeO80WQtipq7sc8/E0JZnVKtDL/FTcWVFYtCYxsGhEs08ow8t
EsA+Si0WPDyPjkFDpiIFEiaWeB6S90TVp7BYSXnqtYjpZsnP9OGKG93w1MvK9D13a8So9Km7IoV+
vyoQRJE6fIIivsZNBJJB+lfK8XuR7XCGc2C9EjR+a1YmFebPcpE3yFpiSposSkIX6wkCGSULUXuS
pjOOzDm3yxBZY5wq61bYWG4tdo/JU1Akp4d9U0uJ+YblC6o9saR1rXzhsStRDojKnPMHo+CI4kcb
H/fBS+TtEzp/rt+SaUomI2kVGGKwuCf0NbjYfEl6AqUtgox3fJUcdCclRzBZaGL9bVDK+Wz1EJKX
zAteZ3zJv54IfmsYPOGo54tFWyKN8Hs0wtmg2+1oTBpHAAZsIFVBUPSR3zeSe8iFuYOjSvuHJ+No
bXsCSsY3b090okhbYpaMbfeoNAPoZTq2YTWJKPYBIIEkuHiO0bmOqZ0kwSUm5pMZayj7z+XP153V
JzkRWYirHFEGVcE/vB/gPA8lIMJ6UBV4LHN+epSHut24KquEuhIdyyQjEUJVtyuVJD+y4i6k+ygF
M6+XkwHAxMZmvC1grsyF6w8RCa5GQqUcLWNLuFZWR6yQ2vUBaIYKtPZBO0aXjH5OtuAiMCYE/U6N
gBtjvPHlDAFu6U4vE+8bdYrbq+TgBHIAQI4rj9kVtCnF4b3b6mWE3qRYEGFAJKNWh1AjcP2hyZQk
3vFet9rCvOGLc1fq0r5bJPVT0mph9+TYqEC/kKtS7P62nJo3qpzVZQCHjQbpZDi8E+jFzj+EsuFy
l+ZNcL4JVdAtCKpZcu2CRz9WWpOUzpwXEC89BVS49XBDMA718ormNuO2Eh3BqF0ejCYDDsqgAiRb
hTkLffDKBoHgXBmJ7Mytz5HKC21zqQOiKODobgOV65859e7gU19ZctSuRmoSP9UXs5f/qeajOWiW
rxkw5hGUVdN+tIr9Btnq2Ms5rgQ9YsDXZ/1hY7X670DlxBxN8/LGIZ0X6bIaDp2MuDaCqyKUhFyc
9EjISKb1c6vJpjETbbjYaFGogiH5zO4eM/0nC6+ZCRNsBD3nPucqsinAA1v9PyGgLZX1j77BlRvA
QthHk5pJIyry4qLM4pFQKZ/RO0Me7DAeve2VXptGmuMouog55UoYeCNzVtUXfnKETOYnwdLBxobB
KgFUsjgz5nr103pFPs152Q0EV/FxwAVWjNIjTQD4jdNAl2PvEDhiIjmIEiY0F5FJV1/6JZslrZWi
NSeK/uJztRkgwnYHaeQ7OEhc4tfSOx6bCoF8Utun9tT8BfDcyGQ6MCaWf9B/Nr7n+5FFKNdtJJKQ
JNRycCWGdmG82Y3YgNf+2VZ2qGDfH+NPqlAjm3vLKx+Gg2drpjdb0QUfK5S0h7ym4DqUU+bSoAot
wvraNwa9qm3Bwm9PfTTDcqQcG9vqz79EFEhuwppdUGQjLk7dTrZX988IdbRMcHyhb+q1zq94xfX7
7aoasfKlJrIsO2jbsu8vM6AciYRx2C/GFVLrKcocK9r7JpMNIz7SzQLfFy1roU/mVKQGj+NG0cOl
UDfpk3ZbU9v5ZsOjbTzJKPvannlzDbxLNxAH+9dY31cCJpUcuXtI1H06tg0OOpa1nLYPxlDmv2S0
CH3y+JgbyqlD+YlGG6zkOlERpQ5uZrvT+kJYYenJz8j/7+9FUA73hIh2IinPvzTsXPOH7muknP8b
DAcMWq9hzAX10DBFxkPK3iO2EoY4l8Fcv2f+1cbHmUmxtwK2VuEfri+7NmnQeoqNkWSzmsVLfznw
HP/RjoLmFESP4VIWGzGw9zFxIdJqa0RarHSWQF/DMJR/9591xp/az0LygSsCdS0+0LzCeuSkKVkC
VqjpKCTaT7J8i5wyDpaJB6M8qs78lrfzfYVrD8jRfkZgOAYN7KbqMmWC2b7uU+9btKdSK1W25IeL
8qVFlRMymz8wLL0EU6nrfwTRQu1TpPKCJr4dy35haiFiciL1MwU1PHm+JLyR/PPr5MXfrdY4ghmE
2mLsGSQ9CmsPG4xEb9gggp6CyDT1Zl26BRwkG83MExnco5JFZQjmUN1ed73XqlulUJqRBnLse6AO
HUiY42tADjrp6DJAE9rZmcn1OJ7uxUyYGz6MWJ/j1eJXjGchVh4eZrPSbW6baeR4/CipFx5X4Dm6
NmO/ztqOT5GQYofJ90ckPVmwrdgK92kogC6zgR+xILqd3xpHswCC7ndmUeRmwJIJm7iqUgDC8b6W
mJf1RuaUhGLTq9jpChRdvujjx53Ya3tTtbsUSN3DNrvxyb3sE0KturtC7wLFPoCYRuJzHvbjrUQo
BhmfJJ4Mk75ru0mLm6J9pqI4bubGiqGJcUF9SFsvZwn282eiO5blJJ0UOKQLpFpxIxcctfaM2tjI
B7YU/wQXH0rLx/dNr1Xwbo+5mmwpYx7u/G5NcvUKnkMNFo8vLnw44NVCrFTZkpmN8kHixVvuKKfQ
3dCRFRd7xWBRacjy9Tbr8MOzVefpbEQkyrdcQ7psR3pxET5Q0c96zd/rT2/W0AbsIfZ6wm4ZsYHp
mglhDOnDZjqArHVFLBCV3ngIRTAN3GXNZTZMOqwx1dnxQZx7qvVMaBP/AKuJcyL/NQUgF/DATw2J
lxxp61FFq9z/njspyxV5kvEdGTOLsQPtkzoYyODCaXaDwbUB5FF4GwX3V7jV8Fovt2FKc9v09b+2
cPVp+qnHfPjX+/lG1NquvI2qafBT1ME2mOlgn3sLWks7dWzstB1SRv/JSdZSKzszudV4XTepjQF9
x1kWi36Cq6v6B9eRIzKPa7s6BFE6G9oHVRKDnjC7/69ZRsk7SbanmhP3WoHqKPHyGtLOFs6SHYm1
wH5KRBsjFkyyRE+LduCThXSAFucg7YKbwtNLreo/fwSqysBDl6geB8f2S2p0ayIZolrDdS7PPWXi
kiyHPPOC8KeSuwTPzItil3hDT4aIaktmOUiWCkMltWoAaiRIsq0LmO4bqvLE1Hvm3Dy/UDywjcPU
F4g7rTBlpL89lfuL854JxUiDSUPpaY70AtRlRkhrjo4HPem5J6+qfqsgcQHVgaInXnEdOaoNWu7u
s2Zw4Yt6VadtiClUvnrNx8Rz0I+VqM+ErF6aQAxgRfCXgUR5/gVsDIvnMPIuDsGqIjT69VKWzc7N
PQX2uhVEjy2y9urN1aiG+aTQohhSAKCn98mmHpxfratSBt/IkfQI+M3m5QiJorDYWBiWRO/vwONR
3WHR/f73ef3i6CbaA9iPN8qjTyoqMqp/fRj87B8dMTi71CZWLiXkZSlE217uxk4pAv7gX7Fn3IEo
5tcJcXRUsNgeE4eTCylocWTqW5FCDxkzF7sJzH4KDokqtxWXdMoKQGxdjPxAnlbqVljcx7ZdG1dk
FlcqAEfa9H9Q9vfZrWJGWSEil5Fqe0D7lwHsC06cnjuXmgT66o41fzHp5EcmEyS+Gi4dWNn6hBUz
V+Gz4RWThfm7WkvUkKvifuxXP/pvwryeUDwQHIfjM6BNew+nMZ+Hlu4yM6ZEcX58ELDjJkKm7Xpk
pjXpx6Jk+IA5byNBsTi7pG+VRdenvAoA9Y6AUwoVngW4j5lg/iIJyJ9ueoTocUq5YUbai6puKoSL
wLiSrFbRFT/hRApfJPfsrW7jUXiK9IsfYEbiEKNP51j/R7+tsPUaEvW5ckrIEN0gZxW8HoIzZJlt
HKMj8KnoXq+fD1UuvzMIfD7yvGyVfH+D7pqZABVHaxLRqCcX7icskRousxXOOHfcSsuYPc1r9MQa
7Nrfm2oQWEOiqZsB1LbppQ6tbxpoien3+zQ1Bm5VwSb8pLT5icdNO/ZKjSLxCvhWlbpmyFi0d0hI
EE6J5FPbgFwRSJaEm+corRWDod1dPTJWPE2KhpWDdNG0YjyRgkdlHbdmDh2TcNEhEzLdrmJlyJI8
QzdKndyNadQIr800ZMXQrxhUGtiMlWPKjKuR+YQo3cpGp5Hv7fTKgeZXEDfi/a+4lNxdkyIkSJdN
5YhHrpUzXyy1tV0OvRMcFTbuPFUrZ7RzNY7pxgni8/Cyf/qUgWu6CSzMVMScOFElsoYcT7kGdIZf
YnWVI3AvF5VZK9YjmAb7U7XIJ5phOZS6ocS445VBjvxWo/gccFBBpBU8cqrh03QcAvPoJsCqSNbi
bekl0EZ50pFf5QBJ3mqSjweizsVzB92Q9u5p2HaUy9bQJ8YbAxbAdXvkbNjV+Idx4+0tCmABYXD7
ueqZcIQN/2SiSbgV+7WLFGWvPoIOYuDDNP7Fz70CCuksavYbaOk121ICjPiMpiPVO7z5i+ylOdRx
8l8OJiwzZHwnxuSfQBUbUHnh8DuPtK8bE36XS9tTnrPaqWzqVP5qR16xHBUVrAGuhXlfggkV0whR
y/rev2QfWpfdF2uELlc/wivPlElFgDnSCc7fvIODtVA8MuK3Jd513HmiR1oM3oULxtq/tXOzdKRa
O5aRVMgs/E7kjXiSMxgp/4DvqDtKfasLkmkwA39Tr6ezNG/YJuasXO7rNR2kkc7n7P4la7UrsWoc
HlyNu4Cm6y+MmPxvcWBMEKjDHuLnjzGC8Ta1g6kAlT/SknV+I42hE37PgqmQIhPnQBcjOY3F/Tpd
yAfg9kOL0gfgzusXrJSDbgcsZ2Acz1R6wAGL29KuPGnGkj09HiDr908wDBbIzlUTktLBGk/rEylA
psAo0fCPzbnOodreWTAGiEcxErNh5wEBgeyM9Xop5RckCaYh59tGDn/H4dgF14G0WzUzYS0aPk6Q
v4jBQPinBMFca4PaGbTgHNG69O1fkiwMOi4ufxhYsBIt+9wYQKqhq20MPF2SaW3G1Q4MwRyFnXLf
bQsl3WqVhd2db6hprQUlSPLAcyLUlP0rXj0TyU9Qr8ihm/aA1K1JN/yhiqUp9YqXNUlHc4fytxY2
VYyVKIYNAwdtd6+sJaLPeCa734HyTmtPWmaNgxm/VB+Z0bHq8DccdkuW5VjaAHtClP/GKlp5gnnl
PQW2R6T+VLmNFcJW0wfVBsBOvlNuG0O0EGZ2lrQcqmlBa8+seGcGHOgMSn2jSBGb2NBDNQD1/1G9
YNXeIGA5jZdUbfvQmrzL1axHQPu7pnhySAxJUGV5dHFluRnVAYMWFJdvi82fI7/qP2lQ7ggmI5+u
WQx16wm4e7NfzqGanTPLlmQxqJQ5jcJFWlo9WhBLiB7FrLvD8ZzgMYokxvEzRW2XzNY8H95OU61W
yr/bwoSzM6YaTNLofvB97wh7h/wb/kAPyK3ZbPDa0tYyxdZbBLl7V935V3BAAEXjIfp4XsNKuuz8
W2DzK53hA0+SeD+ulZ5llPWt+AB90deaDdj8EYnGugoYAI0p+atF/Wn68NBiwBBPQ86bJcTZa5Lt
JzeZElATd+nTB6jQIMFoNbRc7MHR9SmiqaA2RYdlQHr4/QBVxWTwwwyIhQSM9a9osL3o64BAXCAi
/R38CnG4etDLrY4LA4ONxPCm1laS+UWXmy3r+3m4QZnQuntH+zS6ehvrWqgEzWKGEC+wDY58+Gxk
3qj8froVAN3WR0Irh1B9vEvNCPk0UMAV0b8y89lUrverZltqFMZYTykdPUP7V5Re5mMDsuuWT6lK
VS3vQeQX8VgrZF5lEE2UaFQUIOcmP5jK/BdrsJX/S8sA1ocxq9l5oik3XGn1WZUANv92EvOWCWU9
ja72h1a1yenI/kkVP5KD7F/4aq0f1ib6nrzTCHJ/OfyddZqC513D4jhsGyPSrvPeSB9wBEXi0PuH
tlv/t7WFgUYs3AxY9EViB+H0TrJtQDZn6xbaMj1MVJjg2jjzoxo1JQpDHcFuf1B3DIUPizRwuVgM
qcBe/4vCtl8mliOBf3I/nRckPAOQwi1ZVNuJZ909HalPR0EO1sDkYY6ETHW1VwzVhdhbkdlno/AL
fxucyhLbS37UcDSXhQlyn97XHohkVK+IXrMxSheoa+X/KbLoPkTvJ5dp1RzuDBJQ4bpJ2nKlXhDD
DCrJOekXCMo66eYLN+j7n2YTDjAjRdVhMGgJb5u2TqrpB1Ms49cjQlzTcKP6vPV0iXUKTrtGCWpc
c20LPSrhLzIjS4mzFvHgbMOnbOQcI71BYnB+GPz9p7Numyuqa4LESzQDKM7buq9oD13yGV679kOW
F44QR92lAHhGDFXIpfGnq5xHsivOVCh+pFkvwUpJzgR8p+yaLpm6v9fzdvJ2VItQTIcopxnhRUfZ
gvnqD3FTdJvnAJP4w2/ClNyhDO6uD/ktO7qpFYK7PDoolLntxMSvjaygIkjjSOq5LegHGTNC1zOv
juR1xzZbhN5NnseBOzXiR+ADEFHqKUSrEjqPrQwqkZhrfn3Q2qAZXtj9i9gNy/w+o6ZWV9aUpzIS
74qchbhq9WoeLEzp4Yy+VTeuPWu/zey31DmIXlfq240jEbDZtDpVl+QsJvJVo0nAlKDkxhIdUYGm
6D1tkkg1a2Yuo51RgJDu0NXrLAzPRcQZquFBMtgTfJbU3Q7ODXgek/2e2jKyRx4ef9WXCjFy1hOE
4QXHd34HNWc8zn6dLfL3rl844IOiKfnAB7yC2AAdlr9EloXA/ZxxgsqfWbGrFj34L57A1nY2Zrnz
CXg82ksteLuHph/Mz9299xoxtyucIkYmMcv35W5zlRov7+yG1KbtoX9bXwMGw1KWY9nqGjcbCBNA
CGKIO+TI9wOtyjqXjIzK8RE7Eu1XiOq8uQ/NXzxLmQl3QAugzqmk2Fp2RYyHYFiJaSHdJXclgEuu
F8rLhvILxokTA50wEPGVGIbkNWfSGn0UzmR/gntyk/7ZD5c05GEBlN8Q0V7Ye34fMmAE/gKj00zO
LUD+YlH8Rx7R5XG6qhtmKUk3FWxST/GDItSsvJLOTaSgcdvPfSt+1164WnXuVtPU1ILqnB7zjm1N
8XwG+9ArpGq34r5MPlofXLN3vMJkfwttn2q7LqeFp7DVBQb99PFQi79e2Jxj7dqqV7gv3JGgluuL
DyPLoC+WuBIyLVnEhXglLIdKQXsGQAxhGTCH12eAOzOhCKC7Fy/WsHtZY6QbWpgcfNWC7ZQ9e75o
kkyp/gmtOgpwiS+xeWmdPEPxoFYsHQut9pua8RCIX7onbhxq1fvszqVDZpvLq51ftd8tt87EPyK2
hQSkJktmsibaUgBPjOC6jYb5rzwSiPUhvm0BUrG5EnC1BXwEMQS+hjEqRuUOKX5wEV33jLC5qjNe
nqlW5djOiRw5bgTWYA2xbSP1ztsq/9wRdRMGJYVbxFuYgi2wpst2iTKNyOJBSmDrF/v7lVCFq6qE
CcnbPv5PSPMqJlTANTJfNz2o/WW3I6MqLNL8kyvcz3BAfAAZElJQfhzBIOVK/yF3XtDEebKKy313
QoyAR8V7wcpce1oykbF7q/uMAr6f8221jsopcfX/QmVfwwGpKRB3SAECcb6EUHknfyWc9ISIh6Qg
AbixOhbsYiR0wSmG2/BW1KA3KviKMuZTTsNf0EXxN1gNrwcRrOxQlJr7cNG7xpspZuI3b3WfqKXi
rRNJ4m8vlFy3T/C/qBx2wu+aC/A6H1fNGkM52x4eK+z2a06nDTYFBpj2Eu/jjusu3A90ZD/1jvOC
Rm1PwBVNGhqhhz5AocLlTAIE4naRFJ9K9AaI58EKC1tg2Lth8S84ovVF+gLAVFTjJU8GnbUy4Izr
OAXb8QotJIrHs9rCEK32qr1ILLiu4eRdhn8iPGqkaxLQaq0r+iwhavH2OJd4AACr9WCn1Lji6cqA
1vqwuZITx8QU0obcdRNZdskmCUgC+q6Ylh/B+R1GGrKrug2Xqr8apLKR1c9uWDGCvLOkmEOObTBl
7jtL3t2XzidZGYZprAKlXgDZGalpmp+fue5hZZnI+91BroHQUeNVEDhGDxjDs6FP9rvlkj+/oiqS
rGQDXV72er7oubnnY6hUjl6CpVejrCD+Pvl2U8ILR3dSM4qb6UwuxoxXQrnxZ1AGwlCpAVaWViJJ
sRohHsECf5kn8N4PEAWrN9eDlnu47RvjteFtMGnB39yMU7bjF7zZXIFY+pHLsvWLvxMQG3Rgbj0G
yNWjKkZw6OVsPLxLCPNBL+WPN8SQYVjuVtxj2ze/NTAb2WL7C8iFsWbh+Tve2yIiqf/vDDZOWk4F
9g6+IzHbp0JWx/s3i1GjtkcpcSDFspQmPilMc3rAHfO8LqS5ktel22/uN76udpF254F+cgqfGeVO
/LDU1DdFSRxp804eZu21BU7Lb1yNsvyt5MIB2zjYM1p5c3VkG5ePDUzJfStIivFj015tp+fE1ZaV
pyClGXg085s7J9+tTzeXDOilYnCWYmU/Vk+Z8I5AQ7ip8PSk0pV2ybaOhrlGCjJjbu4aLCbsh8lc
JNvZpSx12aYvJpZjLP2KotEFoq8v5H95upRgGf2m5PRk7zkaWIPkXxCHm/Mj90Nn3ztVvVTTV3D2
fbbeGNhkgewS5hvfQMIqDd9RS7jml0E6oTGaIP4A4/+/A8/o2IJDDD5Eb5orY6aDTadIguFHK+SE
a8eiPQQ5AfqGG2qLQWkhJbTzjlpj+cvP4PcG2K8pza3wRnR5cDKFV/FzzFeLQiGpyiTxa9XiWqo/
aTeZ1TMK/I7QVWyoD3O+O5jRVyyzlUh/J6u+ByN8MpmSaLUkjzBKjgLTUY6t+iWRNJwocNaNOQsX
T2rWKCMdrMUbsIgvhLV8qNz9IJItHYfS5NGNvX96Hk6M3N+2fe16STHZkQSRRZURANwKFDw2ZjsW
dWRo/+TZMZvtzrB1Cci13INhINF7LmyxCXSfOstGOQaW4C53LvrP5UxBPGfRfil8i7yQf4kzq/Zf
X8NWc4xTpxffW6lRJoMTqoD4dhUN4Ceiabu9Xuv4ZEZLh/c+2LPYeuF9FW11m23iVq7W8oUKJvbW
s7TuXP7s0rdTNglSANtuDAh3HcX5+2/72UBBLH+hmPU/1nhVmkDUBXVF281m1u0bFotuJH7znsrr
zhNRMZgPkXeIwpLfD/TIxuIw/GdFzUTlVbXRkru4D52FadUVvYutJFCiaprdN1Mlj0LXhGIDtoi2
nktInLQVpOmGX33Fc54hjCooaukNCz1UY+KFutVyl7AYDy0bKId3+W2ev8yYoQabMhsUoIA3E+wR
sHZeXTFCAXuApWd3VPqAqss2Pt/6h/nnw/kOYR6U5zwUxguYzmnmZHfe6Q1UOKjYTzC6mMi963iQ
9EvvJeULRIsOe9mDx66h3UccH/lF9ehqiCHePWdQbxW7jTzljy6YENHDTxOnPT3vJDns5+1S9Oiz
CZkf4Whkb7EkhVeEarxHd+kaq2CR9bIY5z9tPLCDWcFjUofPiaZjPmSKoIphn51gig4NG8VzQbic
YK0VBcrycxhGzUExnCNdT2YEkC83jaykAe0BCQRN8ipbE7weadjXcBeK7NLG0xnfG+3d9X8EZP5u
PwNQVkuuVcYZGWYWGb9oCzkFTnaPts0m5Xr5bR6C3/3Nntfs9/afP9DCSJmHmob3mHAghngJppK8
fOheh1vi/WmxkrhJhIjL+yg08r1E4bbsb6dXmCnmsI7RjpMoEiL3W7sSHXjeCmYLtLKhb4Lo6cW/
bJPY9alHWBd1niWTpLQvlAxCbmIDMiWGb5bxjxjAZ2OqlPzQsFp2puOIx3nwCsUYPMSm8ObPs2vb
MzidBFPzh6/BZtDrfdUgtxdGyudmRJvc1ji8Wexb9t2rSFa6X80lvBXkjLv8a1IHySDU6G81UYKQ
HjWDXCgNJjFXjQf5mPga+P+WgTFtTWhsJHsHXbsl1xXzteOiIHpGGInzEiJB8xUGGkb+IuPyuvZG
p09/B8uwMq4Kmu7nQqZtZ8C1Gvc7ewujo0AS2TLPbTPGHxK6E3TMnuMm7Lod6sxAfM8HymhAHWg0
4WJa43J5TCCDCU8RUlMj+QThS1IiyEEqX3lICnWZZ/baa21m/xYjeIGU9xHgxH5YCn3LbJraTKKn
omk5ieDBfacgvHKOJHwBy12rH/3D8GFQ1dRqGxrs0klyy5U7dHMkkD8GtT0sx0pN1ynvJzp8dwDD
nUbCFeLcTKMw0dzVsjCM11CmBOJLHm8n7lYX+0u7a/Nn1xcboF7SULEN6YZeeccxo2Krm2EePkAB
1QS5eMys3D8yA5WM+eeEKGJnHYmqn9kAZM2pOy54wdiaP0NPHqG2tlje6AsGnlok92Dg7p384gWj
VdqRcWFhX3aBW1T3aGsrIgWc5EOPpTgbbTIOjVBzj0cBN49w8xL+Gi1BOWKW78S+u2iBdauHQeWm
ZRU+kfEhTA+QoZ/RsdAZzlQy7tzeFgUZsa+vhKBMgeUflLz6vb0GDNs8KPCsMu30qdKNLvJXCljA
W/DuSnMKVRcN4mwZCKE9UXXkurtXAs98DdQKwI4zkfN4jOGUJgSjC/Aia1tg6ozoxBxMRMNKHGza
Sf+j0Ab2x16cY9lEdyWnkxurxAMrEwtt9cia8uA8+f4dpqyKAjEw3dcu4FZGJOgSmRUPy4r+RPhi
nsB+sZvCwDuuPyTUpk/lOxxCm6DJGDd+S9YM+QRndmZQ1fXiY7Dpb70MCv1xBdVDNVcypcwHTzvi
o7QKoCeZ98bTzkIqgZVCJoFkeHeNmImXQc5oe+Gj3Fx8H1ft1aJ/KxSW3A5ozrEWqYNx8veDIoI+
k9Bw03vMvo8GuRgJ0L8FY5vthq9D7WU23c2BLL6K6oxJIqSCZ35pZL1tQgrikTQaHLxp+jVb0w1S
QUFYqn1kMXFEXPNeEguzGVQRUTTOsf/1hoNHgOpdwTVOwQNuwuyTle31c/8M+VZgLzgcpkMw63Gw
4jX9qSgj02aqaBq8c8Q4w9ssyYwgmscwb2y7XB6OudVHWA52a8uDEZXos4y0AfRS7Rb1viSN3vKU
hltgV2RH6xoetTDNHNpFX3+8EE1xDJYNIivuzjPx8ZOavt/n5nkiPhJDqC9gyy8lqVlJ46kIWcDN
bCaCikncep2uJ3SjWk+wXRCj4Xmi+rJoM0rjPd9LEHmQyvRdJ7DIMuqk9X/2l+f6R9/AZTVrm0sj
EREs2YZWRCcg1pqNbGnNAZsPUbMW1rZnghR0RbNNJ8VlRTNsfjQXUNsX7vuc/R0RMIN2UAcet+1R
l7mQDddX/mMiSbLDZev5YnMlZ5LkbzJB+PL9Svx+tolynbgfR8zpHo6JSQ00X03406RktewBvWor
QH5IQKPYFRt4zGkPtwwW7oKU4ez9lLK36I2JLghfxP+TRt+mfO3uxqNHwc1/PXlPAjf/wIGI+gTF
OX1dMa84nPfiF/bRXRNlNkXYIassnzjQBlgGughntt+iUgXYIhW6Ct2T/SvtTElVEeZS6D3Svx6d
cZj6CdCPhJz1dVGPs2uI+UC5s8TDQxbKQYXvGgyxmL34fk5xx7PEQMMECkhNQftNj4Gffh4nctty
EoJUrG8cJg/QhVC4cTRNxR/59TUb8lZE/xQOOLomFxBNpPYTt0jwLU3svQJ9SSyAK8sXM3bOzOOx
Bdcd9E+QoMtjY36eIivSF7Tvj+LsvSSsfe8DB6+xeZoAVonIvnJNzrffc5lcNwLormNyEdWp1iPo
2njnZE9j74wLnn63bc3P70gy1GmdDGWqRMO5FTcocpaddFaOQhZg2nApvw1INwdnL9JaA92rYD0G
moxDNjdgbaiv3sSPL9o7MlMlzomg28+HRRQkpWO1FsWlQR2wH9lXsAvtPFnZOkc/LIv+YN1duzt5
Gi9BujKatvaoN1d7NTZq1Dwy1JoDDtFPdeRWHEKWMYFP0fE4wVcgqZYWTQnmS7PAkXGBBy6+0iYM
b8emnOE813n9UKQW/q/aGIIAFg1D95yiUYHFpO4093HDxa9sbPhp2Rza1nOCPVOMLSgf6O0H8wLh
g/SFz+RC4ZNFRKSWssJ6JaOEeY1W0rSZtgO0J7S4E8XhI7iFprjWhna5u0HXP534J8lSp+6mwqp6
Rg/dGo2HH6EjMrptgIS84YWtMY9tI2B4wTeEw50hOdOTwyjysgMgBRzqXzDTNFuRPvZF8UU0HaYX
LNAGy6OyVBOmYU1QQspGBXwNOzgS002+vHrM6sTlyaosXtB+i1KfQCkl3zRymlwLtxbtnx04t+Ck
fGQq+XXl9ys+ejy3Vz5KcBthPfOLjLm86ueDkgZeWqKkckEL9/jxmYIzolftJwz1HYnuOGWINIDy
yezQHUHCjDKMQEwwS+NALSIrCPACt7WFh6PiJghaoKXjTKEOg+J3hNyQO3cSFUt/aU1B9IvRQ+Km
gxx5wxGMcXu9Pr7tGt2pN5Lh56ms72NESNF9bfWIJecWBok48TtF/dfCrML7b/wUp2YbxQ99x2jh
VUfPMA+7mfVscPaLQtV1PZHCwvLIixUWYCfe71myUvF3r0VcSAzQpT/Rl8UCfM6DlHDUNRjwV7Dd
pKZ+ilwRF0JQW6fOFiP2CKZi+tfgmyPIVUpx2A6DvG9gF1pyUE3rCVsEGfGTp7dNK2MORMGflbnr
zUk/Avgmzx2rkZ6nBfWeo1Oo0SKRiSYiCguESGzupOgotDQs/soHhtYatID6cNeAy0LiYqQH9dQN
mleMghNhUQXJHmF6ooP4h12FL8yYQWQENjs3WHtnFULlLG7GeY3DO5uOB6+ZIVJctsOUknqP2nQq
LwP0J1mZc30d6z9rSG4BrKfb6nJFORjoNaG8iUL/E+XN+m85K/egtENShfLCNNSFXN76TiU0Vg6H
Y4aqAT2VmRvzdm1JVpPaq+QQFhAA0iSMbO8WqgYgyCvYizY6vvSU6Hq1Xo2oF19giRChMS3QSUGx
k7IM/BHYHnaR9pVqgRtQypxjr6hXna63BPG7i3XPr8HjBKg7gye/bsdLyS9onsiDOddl/ZPGh0jY
YrtcMj+56fNpVTmVhCF1Mw/He7bUdjydeErx80q4K4Aiyy13w95b2s194BcVeMDf4+rzzVBKgloO
RhDeLqRY/kL6VSJ+5JdWhgdVcD313TWu8UkmuSjNObLrGyfFyZa+URewyg4A+cfWOBR4P7SuUEl/
6l9HOVMOE+eM7XXEhle0KulVUVVaAoKnvUja+Pb0vqFMuds+xCRIECya4ztPbbc9SFnwHLu96MAI
zDPd+DqlKOz7DCcmzKRnltbWeWm/fLYLvYx4MAKxKxPDrM1IhZ8QEkDwltlYlHGlUnKYSf0YHd4/
JOP758GQujzDT8/QHyDN/DMbrvMHUBHwXW6SRSUfbcEYt64zBqiA8N/ox2mvjFZra/f+J4oMVtJu
UBIJHkF08Qzz7B2ZiMzIUvaIZSn7s7zFbpS/O/Uxqe+2/Vz21aO1oIAnBsv7zitSn/VO/mNDmK89
CuyzfNV/EYyGHRaHLAhWcSGk13Mn2Kp1kGCAvolF59bWvqOxGF91ckldB0Xnl4TlHQL9BKwsmnwq
5g8xbRRcOya5uPdt9WpUmMwY9+nwNtDI8ztIsY2N1FTAFt4KwsiLTqalaYyvIxj9KsBvf+CoaDnt
IRCFG1C3RtAwr98GFw1I50C8DdZlph7XtYU7G3MreTuJIO2Ah+4vNQjlUB+62GDO+WA0dmWkk77t
pJ2B8KHWklloIwfv4yNzZR0AgQLkLpB7KTQTieFzFoRnRSgl2GtJMJgfRUAcXnXEvuSKbl13rCYP
LT7XDBiZF5hhVqBY34fEQeVmnvEkeHQxYeJz325wEnF9Z3wXwAK+3GdGdW8T5mIDrM4MuS8jWtkK
rv7/5Er35asL5f9YAWUOlHCcH4dKDMRH58CZCqBc95pLEiYCdrDfbQFDtFiFivOdgv7jJYKgG5V4
z3K+T0QacpU1s+GSCXiVZCHXWQ64wu/+M+2EDrDvH16vty4c1p8aHD4Ly9PdEhH62UGMWda0nxUz
SSDfjbZnFpT/RPXZ8MrbWE4GfqgD3kERS+GrFTKUVHhpoQmM/7O7xH8uve9J4bN7mPFzj9dysVtZ
iYE6dSkSqdzLwrR3erxbwV9wvNv0iEB+hBj97MsVWsmvt0ZWeKr9PVtDcPLvXwtcSuxeD6n0yP0D
m9i1Dw4VeeyeXvZWmb5chq/19G7fVteJQ+XhftqbSGxFd4f0JYevabLju5BFOLAtr3Pg86d9kw8/
mjF355P7P8PrQi3nREfonFMRdLsgxZiaksxE7yTG6S0Q9j9q0Xu1C/7Cym4mnVwQgKOLnlA4k5sK
iN2Onkq9j75n7OLBgNjd1XKP2+eJO0JpdkAKdUEj4CSJ4yu2qQ3q2bO5S0bv4sG2vGEj6KVGoWO5
s/eWp+DUFGpRDOMIRzdUGa3BFGXLuGfkDeFgWWlnjnvzSQw0eGvKGbxCMdAZLkb1OgcaLpqyB01Y
kvv46WcxL8/0cUGfAx7AkPI7RXvady9eVDr4HZ1yIGcdBVnyler8Ci4Oa4kyAIV7c4oo0AS7XW5z
iZcnkwIN53eGRZjs1VOv5AEYT9eVObIkihJguaqUibAuV2EEfnsmcUaIryOvK9WVpWXppD7nA4ge
slo+QZtJhr/FLrLFcWf0I1LsbQWaOjdMDJihNv+oNBcAYmpZUZlwRjYX6HSCju4VUhk7EKXVUHf3
UidYmP4Vha0YyIC3AX93MPos2GZNIYCYfrdb5eJGL8cDILhX1ckArHSB5gBRgOzZskeyY4yZVAg+
cRXSXNj+b2a8bVooIs+7UyEseMhNIHOzI8gRGKaXaukIkvUUEePqCRZRwCFuwVpFmpC5gxWnjmxT
yB6EwkpyItFXd7Ixebl65bK7M9YOqz2DHyc963tbrc15oU03j9GrVu5takkPy8qLdArYtDrvnzbR
q+k0nEATIMIijYIpbU6SXoH7lnNnjOdOYM9E05es+Q4tvYhIhm4DE8RkgBhaNGFEXikgVBZ1GM+a
0z0poLw7Z8uySGFaFx/jSiY84hi0XJQelR2c/FNOu3YUg/u8nMfqS+n2n3dRmAM0wtt+93GSB/Iv
2dj0nzbxn9pPghkzUMbgqxnupjnh/b5whwQ5P5t7pPDEGcpT7gH3gTcix3/QNbzR0pv8j5EkFiwT
JNvTMyNLWtlQ5/blCoPp7w8cLLbBpX0KDThPnl3/dcJO2EEDPQTlGdi1QlAVTDscdhYSwl8dnDp9
hRJy2JyQYRuB9izJgWYCXptj1AwME1xk5JDzQ1H4aND0GPmVdwa8vvXPXa8F2055OnXkws4CSA7v
LJagPt1PRABcbgjh8P/mg1TW7wUlO7npdkUa5UW7GgXuYS4PDu2n4LWSxRQ/flG+bN/fLDS6BDSK
EYE3bKpJkpx8mbIiLzWhETEgNlJnOQ5w1GsVjr5rj4H0so2sI1dcpPg9NafFplKkDX48V1Wstom1
edLcM0q4dPsWRTXsRapzi/AbulOuI6MKl+e5y3lI1nO15PT7ptZaQbPj9acm+zcvoojraNohiEOD
ZGWklrBGwZ1bUw7Uh76H1/kSmiy61+paDLtYb/Ty6YwvKTUVt/ZDB7GE/f0YoWrk5/jjz9n4R6dm
mF0Q5sGnXsWv/aamkXvztRZhkFW54IvNAqq2Ixzltqz5jQzdzkktciZZoyaYf9NNYEBiJ49SA/8E
eLPF8T7Xh4LIyjhoA08FqApsIeohSmzMnovjyAVuFq2lFUWyO+hR/V7R4L4DxS946bkbbe8kn4I1
C1oZr0Nebli23rwNMHJpAgb0ZNyry1ygyrQVY6BYUirkdMnHTSduhmxU1iulXAlOnVqc7vryskJB
Fuyj6w+jQrTXLsGYfkt+HDt0c7XRZ1XQ+HmLdXhEcrPuH5PI1kTsl/1t4P/bJyPpZiVTxGjQ2rmn
t9Nut92u8G+1lN0QHPgMr7IWb/6vi7XSYE9qRUUdZdrkNQupHiSZYVAZXCqOGfQ/DT//k77jnVN4
BJs3ydVgE1vdNhEsGtIUKTq7k59j1+k3+9Q2Yy8xUMVKS31EbTDqZnxftEpeaxDv1UDb19NIQogg
VT7qIKixfm4LnCpjeQAdbNtVFclXxDsBZaPhQ2dUTglHqQKGOX1yljD0mqUAb09RDbvcjI+OsoBu
BvR57yngP5vNFdKrE+p5Wsz4TaLNR67ah6K7+fe8IBcGeiYlNSd0E9RQNZIB5jsrnDrm/DvbjZrS
8NU3R3nV3m4Kxg6TD+/c/aXNSS18Ye81rYJKL07iq1/wP8T4KO9YGRvtEsTpwaPo8ReRaZ936ZGr
LKBPy5Mn+Ovufx3OlGUqv+ihBJ/hIMQwwhzyS+hgZ6JTyfg3FCznrkK+sH5Pz96Fm+JxeM1E1mM9
KmESsyhNBWTFPsuBu4txLApOTPKvwnCdcsOkiw9IrjqKT7DL3gonD/J2AD5lwDbo7QB86ULokjiZ
bXtUA09flxcnGdfaxOMdRKBViHPTowduOQ+8R8oUDYqKDG3SjPVuQrWOPrM3uZoIdfDfN5a2CVQk
/q0jgwoHMaGDC/nemufVdAEuxW5WeEvlLwkBPJSOEsqDwsfCps+WofT01e8lDodhhYBOvUYr5J08
6EiTxOAfuwispeKOV+C77Hxj/z2+d7ly3ZYVMsoMa3YL2R8/Va/m8EwTZqYqmmuOUBVJuFHgYve8
UCGi9wieH5QRv/tUfzXbq97yL0rM90ndVUqz77EPalq0t8d7NR7U7B34JAtg2L8/Ci5r0n2Y+EsY
1MfYmAyC5voG304CcQ8RgbAe5Ofai30qNSctohwF0oHyBFOYaOxkeWzCzCLEsjBB5Ns1P61Bmb37
1PvbYOQKegW7JToptT0eVXFlhSc2lady1aK4S3Jjayk+KGInzX97rJzXD8/y5HfJ6/WdQLGBU394
tem735tPzoWCuSoqLdrpyNjZTOWBQqJrrFiCBv0aGnDG9LXM4JRJp8n7MD3uJgsE2STdmH2Ifl0K
ekzv101w0S87NpruXRzUP6LmsygTeav66RuQw/AaWvE/zmMu/sV1jVQKoeVkwBIZLuwGfvTkyQtH
hjoRjv9GneoIF5iWm/ZNcGzctIk7rD+JuxSlCRJ11QUBiIXG5oT2sEVh8uCpS7N/Sa3ngSdviSI9
5yCOP/mhMde6sgyg/DEzdduXsk7SdrW3YAoQW+yy7ca7+MFiUpZchC6iDvGs3W/971tZDkj4NaEe
nd2E6T1+q3POk4zV5M409rE5B9XzDSmab1nrSaOuSXAIRlm3tc6Ksi9VNOBWsy1BwLVWk561798/
T2EI8wHYgAuS0+HuRuK9Dg14ylkK/SufIt0ar/KiESiJAv/dcw/LI1dIMe4uqpKxan35+rXZx8uK
ifv6/1YuXLt4IvRaTf9FlIZiuT1RDorpm3AhK/UYAD0B62UPp1eZU61CirbsNPL0zsg22rcIdSa7
fcac55c2HNDokLo96ikZ9KNNkrLbwUeEMis/f245DIXs+NpiKDjjpPkgtxMOv7aiBXhw7nO3LRxE
k7Xc70tpwcbeiUfIDK90jKdnFwX/B+5Ds997fRcHPXf9XFOanAQk60nrbEzHQnFUHVaEispHeANy
x/0/Yi/avlqDoYcejxVZYyQFoTx+Yx/vXLtCAQrkoIuKBYANQ2eqDhSAtIRkYWkvxHMyzkuyV3fW
QDWWSN8G0CCPFKHt5mowGBsr171aE7iZdnrviD260kKXCpXNV95cetNTCSBus6aRkrF3E1teTKxg
X/H0X6zD5Cm3YgI25XF4hvK8SbsH9S3u1udSJx4w98sX4bNza7AMOGvloMwrGUxDOHQ4l31naOaB
vMPmlAprmHyyd2pdRJy9gjaal0nJsTMLKU4ikp8/t1E6q36RrDPD/9elHj8fiCvke2avlHsljByT
90eYuxIkptsORMUfoUaW/Xt+6Y3vCYnb1CObLPv97EsPVuoiAmYYxwyw42HhQV9tJPHzmmv3DvA3
3vcjVAkLVnS0Hl1il5lOQ9U1VHIetQYhdY87Gmus6RSMbOCqoVCNcnx4O1CxufzoCdXWYh+96Axs
kXieqJWPtmuee7pEeuf+hxm6rWEl/QYMBRTIfmAnpF0iuFDMq6r5L52U7fIS1koboXCliRw/gxYB
dx1iuV7nDBj4fFe97/CSppUAGjV+I12mQQz8ckb16WuMFzmdPHnpMKfjFXdkOy/QYqnqnVnIxS81
yyAM60NMMUkocJpEXckifnIVIki9M4ankoy0dIU4iPdb63oUISeMnwxf9nzlpBO74l3UGknZsxYz
bRmJXZH9RI8h6ahHHSEkgjktpioNGXHH7n957z75+ARSTPhXXKPptq7F68z9XB6+SoQ9Cg8CzDeA
jcB9DKLY0bFK1y4r5KtLM1JSUYL6TKnzWexoXx7zCjzjd58lVnM496buG4gIu8fK32qU+5HJJCmX
NbIdQAzm8CxzBXW7UtGM61doB3nNAefHBawmt6MtRPtNpgDEC5tRUwNOj6PLywF+ZvAGywhXyQ+r
79bwYchG02A1UIVOJrvJP8nhx9l2LFXTFSgJ70OLDJbBU/fb3qnwDE89x/vQUpcIwxtVTo4yKmHy
JkJajJTwDAnQkKzRNIwynhu+GnVK1rxSqSzICGPDBzwsQ95enq0V6nwUmy6Xwl/ffw4LS5h/uOLF
vGnSFEeKEnLZ+UnXfXuMrCcsfCaWAIooul85EOq1mHXHtksW49Z6blOTdcF2/hfJljhjsh4mUIKD
NURQENUEwUhuFXDQu7ZT3AJUJB88gWC6OvNTasTjCiuPc9pgTKO/1rwA+RzFh+DSWU3WqrmQKRY0
ABGR7/TdQEjfSXr9F8cVIy0V2m0YuBlw8078zsaUJe8Dn7KohsPirOMzoyp3xg3JnWFIFW/wrmKd
jmmyLl6LPP8RE1itFqKCM/cvVETGZYAuAUa/fwcimzrTfkLV/vriA3b4bsT5FlQJahWJa8PVWldL
uZo4FkrVjNjJrNOGlz4tmnRrEVDNDHeh7TiqpU/R+zdfZZh2jwnCdJ5dpIluX2Ammf/bM6ctGq5c
umMFypORuheI/569PxGPX9sfF4RLdBKsgDEpCU9sIQUB+24SZKT0TBdbBzgHKKfoOiYvYpGCzaMD
aHjnFtsxO6as0R4Es/L1/STscCdEbhYSmTa6W7O3gs6hVREH5feYTh4c2yDfBj2ISGiOiu6yskHY
PNzPx0pVLYsQC84r+tuEz4ZHhc2iHJTb1BV8kcLXo/E4kv+J7k27YmqRU1rx6A0qDM4d3mFd2eij
M3VqmJvDmsD2J1/1abT3ibPjZK3n5kjTG4ATAeiD67qY+xIGX3/lNUNSKmUW+qVzg4yqJRZ8Xmb+
TfZ8NkN32ppQLme81SHweFH5y+SRBRwbfTV3ip5ey8HkLzvSJniyjAVbs18BNUmH54Tor8X+imzK
zGhACpyuTN+tYb8Ru+cgRjYEboybdDv7U+YqpXqD58gvEAu80wd0xeqJkZSA4QUZkj1Wd6iGmsOR
TOmzj7OpS64g76R31wlB9xOKI1YOWCnQu255BmyaOuc0Y3+FB0XeafG4NNtqExKy5fTJyGd9Q/Q1
0Qqu2AUGdPn9N7uLv/IBcxji85Ln89FV4/ajdZXwoM27x+KS1zR9N74nCKgg1hdMGFonrVa4DZnr
sYCLnuLedQ8x+dEY6I/mK3GvX6z0HP4qJ7tufNu+iEVrtHHVO20TDFNw7SHnFooqX61mjDpG9KMa
vm/dWnkLDsldzXFzI4fxI8bEkg0Ctl1DP0j4QBmMaHeqL7zUiF4CpLHGro0CZCqEfBT9bVJrsqVb
t/mUT2H+9NGqdhX++P+Sk8i8/jrKTYYn/3IEagtlcTbCW/0F+iVYh7XmxLnjqgfqCvy3oeCc/olH
X7X79T3hANH5+qSxhKVEFhwBlCIAfdOZnS2J7aq/N48YvJrz9oyzYgNMzLmuTARI1/nCqCEdamQr
KseorIxeN9bjqjLG3Rk+RLbnsFNB38TOLKz+yigQ7NhcQw3hu79Px3SEuuMGrrVsrFx5lZFRKDRd
Z8Ed0E3LzcPPjfJiKeTK5fYe/c4/nBo/AvSZSguqbPK+/9OedSWMamjiejsHx9ax7lAnQBdAQ4yh
aNug9Zn7AeUIKgLb8OGPRbvdeh8zQb4olYgem6gLQIqZ84ZETwtsQOFApjM0WqVM26Hf/cRVscbX
NU5XTR3Arm7TKQYB2o3eXBeli/DrHPivBoNMxDbNJ2g56fMVnGgzWLIYMdi9G9GQjmbCNVvpBtYH
AZ1VLYfFC69UBs/S7AU0TlZQA0nS/kNq3oFjwjQPD2opyw7ioVNqitDHGqJoCzAHZFc32TQS3CrN
uNxoV95cdYUiV6Vq20hoYnoFzem9itbRe2I4W5C+oXSxMq1Od5pukUnpeKQSFKFirgW0PM+6BB4N
pV1bhoGQL8TPGWyTgVQPwRoZ70d7vn+7FqyZcSY2nGHoCDRaKwcvj2/h6fltJ9MTD2mioplRwGXf
WtvZz5Pb0eU1f989hWW0SOB8nq9RD/uvrw+AthyFBUiAa93nwJe6LpUt0wdnp9ZxYls6R/PaPyEb
MVBj8V/NtG7zi3S8ENCL8fOn61gdhi7RIlq4QJXQWi8qtWFRkRJAM28D7EaoXKHuxphB6KgpCt63
vPO4priauuON2Sl8tdk9k5G1/xxuyQznGszyxYSoZMn1USGH4rJVDdjGwiTHvff+ZeGES3bwS6dY
S577ZsRlwGsRWLfKcgGawv+OqzWTIXKjDnt1Jw0zgqYgiiHTDNLWMJjgBQIj5GwgxUaC86zX9pJJ
7asoXRPFNnPZcNOGLmvffEhPuxEddEyp3wr7ABuI1KID7RcHUOnECPOQvHV5CpoPlQeimjVOeiqb
8V/GBKgmFV448525TIzznDH9PT6EMmK12YV+kW6DUAMi73iQVAy8yQWYxAAiAiYVl5tT2WuKr14E
ghLndgwwXaUYxHoec++G3F9h03cTFxnFySxYBOqyzgJbehkHZuXAkEGuc/kPMEG5h7Z5njj5atFS
an5+hTV8cOjCgsMWVcPfwQ9eJfPrk5XUCLB/mdztiQFsVATFQKPH/0223OUpxALMCpZUuBqZyaOb
O/ikcfXKZzmJDrExnYkvcxx0iF5xfPzJJuFawkILSKdvsxXhU27Odx3zsmZCQKaTfhYlyvWWjVJQ
5hhbFnEb63SDHkfCSPNBy6Nc8jH1/UjjMfD+aMb1Wy/MGik/Qr3EHYKfVVf0BISUA0y3a29NWLXk
o02aftM9lni68mMZMoUix2e8oLnZg32PryNZidg82l4D3OgznZPSxWXg6yIPnDvpA2LOWCKg0WfL
DU5Ths+U/+h5Nwre7nxDwsVgwgIYjaD6rUol/gXRar3MxkcjHZ2iLz4doVt1v1oytoycNxOdTlW9
2PTuEqYe4WxldGBoL2jO3KSGnb5Ce2Hr6JhMCAIEz4zvLF/C/BgBVidIxQDAmpNM815Uq6/C2Scq
vOSxFkovdVfmAb1/2xuWUpys6nKkR6/DXX0BEP+LYhKCouDk4eK+BaGK7mInYdsAnckpPt8DneXc
4WT1f3Pm073fZL5VQQ392RniI8yPR/HqrhUrbGYp4mrnq0fAob6vMSiHByh2+T8sGgUxRhkRx4rT
H3dthC5gdMR0xaAoSdrbrmU19uxGq4hIbpGcX5pzPdejCzpb5NGCeLxQlocsKp70eh7bUrdFwsm0
9RMzhJswHGOM8fBzcUiIkvm7odBXFVI4FRq4XxBCS41RoCzqGzjiuU3hZjJ+a9z5dbdfpzI7s+/a
dRRRtUYjCkAlaFo9NwDj9viE19UjUilZ+W1LEJU0nAbdgW0aqWvuxmzFVhxY57L9nZ7TJH+9ayPO
W2KfiNhUVfcI5RhoBFZIHix5HrS2aglmiSyOs0afFxhh65EXvieYX0DOHt9DCh3MvXhnBHvEVaXE
yAP2TfkG2S+bRBurBdc6TfHDHTqE7NnEd8q1eUYvnfkqLW8ilNIm+ZVWcEAaawo3iYNIE5GgNXZ3
NOjU1Er+Ni0TSm6hS37Wk6WXZNyC6SkVwO8A60z6spIYLsssW2ahWdRMUPF8z2C4v3lKTEGWG5gd
Y3ENPR7Rzl8jeB7K8YmJLfhisgjIt8P/uDEp1ShJV4tR66akJ87+VoEc5WKxAqwz8UhjfClNu1Dc
UEASZ6xPn5aqfmnfP1Q3RSZApKf9DHoLYSjHlLzDNOcWRpx63nDbQrp9CXZn6Sv8jo3Ey+NjqEjx
Op+nxD7GTFBCRWtAQgsPURucsWKuI0SGKbr8q8vNY6mXj4OMcI2SEcTnna1Tyxp1AWe/6mg0UtiY
AHUq0XBVDrGyUrA1JcRUe40v2+3Db6RYKvmdPNok2PdrL2QDuQ+ghO+duhZ9VT8nGun0oNhQhFng
/vo2wPECNYB4Y6B5kYKZED1VsPxcEJ9JODRiFRNEk0PiELJMo+lgRCq7bNN3Kku8BHDkONyOlnIZ
6cO0dOeDqStOzYcrMMZNAZTUICEHXd2kADqhAclAOU/Mmn0Fafi2JUMC/oeOUTR6IWUWzgFLjXYd
coEb5DS9AME+5DqKg++82/ptbRE8TaImDFyyDBKLHWD3UIzX/6f1oOsR3Qr4wvu+9+LqEOikkeK9
ZABJd0hpeDtC0yQlmRjfvXZZfEHhsxIjvHJKOhosvwcmWeuS/H5yzpirEmRd9+xdAaOoyEDSqSEM
mm1OtNNwsEnRPHmQ75t+GvJDh6uu1bdwNcGvteajVhYZD97gDCA3JtUCfxaxi+DQ7ai/haMofXMB
5eNe9HL5iqX9/SCarYLKIyaSFCyVfHYMrWYFGTfCyrIqypUiUA4WsfPqLNuxqQuTXpBVwGoCWqW4
wChbtdCpM1KPsIck9JdOlZxPJL+tRUsTBgdfE2nHZm8AzleGX6PvAXb1xvyPx7vtSRP0BPRW5Nt4
WkVarBKw8LKAXoOffzv1iV+0AZx2e96leGtyIPktc95M5uJTWdYZqIOxwj6lcHNOT4VExLd6JDLx
DijXDJoVoiNuiAeeQzvCUTxiHqt1Jff91Rr2HAFhR9O3IEPWcumgans7zdaxAewUdjoG3IsyRtoI
p3M+Ph6QKsmAfRT8gLP+7F41IUwFa5b3mP/MhKxxG/vZ/op3CgMpv8xBMBXJsIB2JCWqO6CXr9i6
XkwK6a0I38vBbNWyqSYlqpTI0RoapRzNZg8Q7cpC17mHSTeqllnqyIIasrRcDTCsWb3+ipYcfdSu
SeGIWZL8FWj0UyKhRB/sEi0S1nep8eaeu+wHjAXiHh8qHMfUU3UH+DRa4uLzQJF5QuU8GAD1zjXD
EnVLxyHr/dE+wAwVnaLxViRyKyvjfEKSDyB10mPeiY81eoDFWio15i1LWNqx7TyKa17l9JLGtXYy
nO76vFkcOLkQvlNNqZm8B5Miwhdh7XdJucOOofUe0YbNVz/u8EuRxtiImrKjJioa0LrEw2994+A+
DtkUdp5ryu0lYF8qD/L+mrCQkyyzsRoOKT7+rO3Ij7DtpJBvoD0oYPUcfTwECk6pMXmbBWhIrpJS
9bpxebbYzzqkAmNBZgOUObnCxeCunj3tvU6eyNt3nGsY+9WL9ZlvMX+78OYM46MwPbwthPY4BFPd
Y1Lt8JCTLvXT7tqvdyw5rHal5Q2yJ+mZRCeXe7mke78dAwBkCFbQrPdE6GEVPkpDNTHIbf2WJdxt
a3lLvoiQNWbav2zOU5C2PizaJWzdog7drjVaSFD49OYN2un/e10bNW7RJ1gKKjtQwGjINQBpufOj
YC3YiMNtkybNdCd8GurTzEaG5JeNECSdHevSKAWAtGCKrb1eVYT1zg+aSNQV66psNTV5bhc/2Y1O
lEnlRSgqPIoIClUIVyJsqDzsG/EVS9PsHtI6Dppu/NCAXFkk67jWtA8mgQSsNDzMerzU50zEpbV2
BDaXFn0e4SloWqg0iOzfNX3jzPlIXF1JouZX3vJst8Xr3ZYhMslRjoIVfBCGXu2YBZrpkDcPLm49
5vw5NP3UDOqmKSCgARYbIMnM50HFYvXiadR+WEyxVulYW90XusEbKMBVnaKZfPVsLe/8A4SmfCCn
V/7qYbZO7NzgQ37TbWsRSZ10AeotwlpcU8GcCWRQtgbIyguv8MtH3MYZpzCtO+oi27Ig5OpnqrDi
ZV3FoCsWpS8PJi86qguoUPjJYwOkEw5SVdgTqdfC981gEs6W04Ri4rSoag+bV9D+XfBtKfchcqij
BftZ25X10YqWRWWEibtTkUry9Oxb5br/V3azGyKxYopSW6/r7C7n1DENoCS6kfRLNjWev581TrRj
n1kYzgj305OsSFvXXOhW3StD0kBrn+7yHP24gc5uFw6cserMaR6HkO2YIZ+c6KRTRKhnH3755/Gr
dOtUbs5IeNLzxc60bHNUAHy6QvtDNxUVRcYomiKhG/ebbSA9jIXZ1BErOyD3jbAfEshtq8joq2wu
kE/7euu51Eoc5My5y4cE0YxiWQEWEkl39Jhidf4RDURDyRD82G5/gu1Tqcp8NERn1EV4EXYKRjUO
Fq3vm8klXjpsvPiDSiKteGx9H/3Q3yVFbqDPNtLFtyKE2gaqO453lWoZw7mt6M85YCT1iMLpV+Sk
WkyIh1+O81tav1jm8m9v5Zd8gRUHhulGhxFHIkHhvrMSYZIFUyBP9PG9VBwNc6oNfxk4xOrOE+Lg
htYujdpu6sh8aQ4SibSghdmIHkTj0/sRCbx51+bScvAOylP4nC/0z9OdcdSFQGam/qzZqB2N1gYS
qjafA7fVri0vWqRaSqQNtN68GWUAbu0o+bk9km6lg7d6PcvWzNuaGdq3G0pD+gzRVtv33Q4kMXRl
4gSYB1/s0R9GbDlTMTWpM8bghrdTH4pFdKv6qrXl+2Imcf0zJpW+kS+NecfA6NGhAK0bAtnaTALV
c0yL0gJcUBAR511E8IwKlC2A+Pk4Sl/thkzMBq02Fok4li34owovJBRJGhZgjdzsHHw5BURXtl/5
Vh93O91Qe/GfgB18RwE/jTLtdDrpoT+VpPUKf2SS7G6mVuG0BWg5RbBOkOdgDJL7TmQgVWAJtzuk
yKCn94p+r4bg2ug6f6Ql4QIDQak5VGbxdojt6bpDpsm8ceRf24U1Cee5SbkG/qhtS5C3kmGCDzZ+
MTeq6qwWbNif5DzPo/sE5K2EHszuwYJ3oBH+5HFnqtz0REpfg0Nj52LuQJvnRULWSRWtmxECMOPk
6pWcujHQ+9AclWvtqzMqJp3MGB8vIEp1DMvAeTTNfSMzamukY6/S0qOE8emaOuR50slJHykWfk1/
kMoJDBPlC1dhLGdKb/n0C4qh8tRLuGICHZ36OvjBzC0bHyZXDtgxjzf7bBrjI1CCnC5DAapN+EN6
7SAx7z55corC82jbJWZNKvlEdy7osnUOIylRM/rXWF6fLWzTDH0FK4r8Tdgw8AReOnvfeZ8NBBtc
pRbyKTMWR6BbIzG8gjJ/zBHUtGWiiA846fFniSYvjYRlWM6Y1N8M2AAhbiL0MjIey0SyxLHD//f8
+jQWn9kU3p/9/n8jFAK9b/yrky6g2XXRddXh1JnWwl5i5JxwQ4kuALPj+XHDauolqBT69NGq+aH+
ozOrfOpMyS9pUsn6qm4/SRc48pb7mPtGfdqG2P6gDzDCRCYJr2RAUnLCr2Mi
`pragma protect end_protected
