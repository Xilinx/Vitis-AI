/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1082384)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B6+vDDKPy4X737G3crGW8iE4VVVoNbUIaMHFfjg2UT+gnHncg4x9Cc9Xp
vwP+6WPGeRcSnTaxpKmOrA8bgMCKRFDzk+3CQBQ62CzudgJ00ynp6eSLMebkmwa+7Kp2/GCsKRT/
RDgEiCdbm8BsFcBs/w4FUbCH+r7CfGsxelwYHjR7sxCbuQ+uvmFRzEpv+2xM9VZ8qBzs/rra9L8L
2lNzrgxayznWp6O1BNVJQ+faiPHI6JZj9BJbU6vILvAjlnIz9708kZ1LJNjicI8It4lEk5H9uZzq
J82s9xVossu0ZMlfCyS4G4HVBk9OHZcJKQsbWtMKXDc1yjfgLXiXcZfHf0KxmPuhZSkvhbE0sTn3
k596S+S5wncswEEOZvODnMIa/PS2sL2MknHcI/gPkXJi62vqqkg9+v0WubRgrhDG5gAh3BUuHlu6
e8CwkP6KYNW5NytttneekDPJ/mu5cSUwSoATyJLOlTJbnuPbCfDTXIhl1+ot3M1ibOY7EZ3v7Oqq
yFXm3WLrr9J7Z30/WLkZJIoxFzzQCTurNznxtV9knTsvyRi0rYBRtKaFAI1e+HomCIakzTAgBbiM
lsO/KMzVGc7KjZvMl/R0Bq79wJFAuuqNY01UQV/b9b7nxt/nFwN0UIdHzQsljie+ZUM3xDCdW1s5
U5nfR62gafJ7LcK71eStpwDQVdW68/tRSnRjmTI01vuQ0QpMwFZoooMgdIXfrbzmAroM/TjPis3h
mNY0RkA14aCqrPeF2nufV07cv0++KEaGLzMyy/4PXk9QjzU6VwA1FrE149hrMrUmTgiUmEEHaYDj
du8l0wdfo2HEEt+EJkvrYXNQxZmhByZ7ATT1qJ9E1Mb7FTcWV6T11YYkrng+gwJ3ekS3Qgpsy2Ko
7HlcDc/wY93ykQOFGxuauVLFCkvQ7ZTp1ZCSh+O+/gxmNTxPyERXIC8jXRmry0ZnRLjS+fenJzfw
aDqM8mECoOYnVV2Qm5IDOMmYrfI+7H2U6yX3HwCTaR5c72DPGo8A/Bpeth7nFduLjjWEIWsXDruE
ZnLNEnkefBSTTXaFhxrz+gS51VjX0vr7ALSjUrhelaqfsTvlU5caSlw0KEw8J13ABtqsNVE8nYjd
dooWT07432g00iknS2YKqGw3zzOr9v939IGqYCCy6b3PBXz4Z9p1mDVI6VLNwoajwghD5C6N8kl7
ZJsORTVwN08UFb8A6jmSwr2774fbpRh2Oo5Wb2cAPq/Ngum4cVCkJhS1IPewjGjZGqNqsQdXVufy
ddxcoSRUUv0+mPfm8xKH9v0YDkeSPOiec/bdwHxW/Wefzn5P4cFihpz6n2DidcECR8a56OgTNIy6
X6mUYZoVl1gyjq89F7wn12xq/vYtEfSn+EZtKS+hIwmL5RifMQ710EGUvZ9C/H3TeqEPAIOWbEzC
h1B+73MgbWbhh2V59/rOzaHf+uVcxGRRwxtYKmqPc3cOLQlhukXdRFdlU2lLwT8licEavvgYS3Vc
7njFbYx04W6hXIE6wkzwjUWJY37kzgV99M40+5j6mP7M+D3PtQCSS5HyiORJyhsqBQx9d6V3lPOO
N/fh85dBOg/eDegmpb4ZMf6HFXzPYPpJ3VPtXfKaQlIL6g7rHyFgjeB2HgV7uNwvEOTdwYxn5eMd
ng6P5llGQAPoonUn4YvpVKqm/NYoE+2TFPxlPAyR9IWgwWmJqp2/EzUqwjIffFYI6ZHkH430rf9f
TclWRd2uUCBqN/VfGKGMdkaTnZmVxNWHgcUxyhA8+kLsN3n1MXCdo70Qi+n8ITzGwAM353PQc3vY
g46y0VWqS8o6yROC+3McUAM+JGjvyTEUfJLYBkzAcz+3dZ+I4+AT4+X6BIn4M7HcSTOiKXjQQQDX
f+IOr58vvbHmyz2tjXKyA8gQWEmR14S/aB3d4/jk6PurUu0sf+T1e5aEetNcV2dCUf2FmppTrZ/x
L2IttOllsS0k+k4Q/cbQO1SRAfQZeC5+xuPFuESfbA/mXsJgL8ctLruHiujEAYRLnJ69kKTVZtni
f+kiABrxpaMMoTbOHgW+4KrePzh4uGYmnWVIY6gZUKfkmnSghjltNtsjJ1f74ovhpLeCCsgranUy
6cuRZ0UJhl4GDfcx0RDBTb3KgGijMGEdTJofchClrIohEqw/YguNkYrOcz6fLVUKiQgxDlDIc7KH
/eKYzdnVk+IPMOBFJPaGTPbAN/mk4kMGb3v2FKoaBgyWFn7JX2cc7VQZ6nrrZxGunKutYE959qNN
IZIGZp2RHaI+3Bn2nV2Ff+gW+iIhQDMyQtIcMB0St9qEYt6GufKdoKGUY+D4bHBlhyFN8LKNmRsA
vmmi42nlOHg1hYc04sDIgHYrfXpwPfznR40JnLUpa1q7iDnP5EQ5aLtt7tSJ3ZrCljJyQr88op3r
cSF8WIQKM9taYPMcNcqCojHoxXS7SOZ7o3+93I8duNVvwWl6eYmeXC7K5dsGuF6YOdNZQdlX3QrX
QteYSbj5vDeFIgO9esxXfAjL8El6PLwNEjDE4sNT8nN8XMCMBd/EaakeamSKjrbl5t2wfhdvKGLC
XPv2fKcoQhE/a1OsmuCAExdJ8eG0j9bsETmbn9iRwpGzK+jmxYpnxbn0XMtJNwZ8Ox2EWFS6ijqG
HlQwz+UJFd+7lNM8gk8Bn+ZdsCH/6D7qayR3pIrSEf+RoSkkmJKTVIUzH0XJz8WT6xq8mskBVvRw
I6LM/CXfrqLy7rMonjiuPwQETHu24aVMlgA8c1nnIV0InIm3e5yPrtOBxNp4Gd/bn1biEHiiKKFQ
SDbpZ5tBdbDFyvR51macf0fyWnJM+1u+ZLQ2XZHhgaH1EoAEZkjYxYcL5qP7lKsVvvXBViLJxqBT
yoWp6XHIUI3hC7dUIFKHivJy2iTZGI/+JiWgNHWIptPe5Ew/BXpIm2pOoChXsbctpKs7vbTPQGJH
N5lp8hBISWm1lGVZKEw6ja3H3X4RYMs2e/KZky0qBclVlg/iOxDuuKGBhVv6fDfGpF2SwZQxeXQf
MqrtfLDpe+3U4v9y9wLIJiWsluSEuESrbAIbHWpXecCMC5sw2eP9hE+W1ytQGg5lqd+lVaTYgiEj
zELrTdylqD0KXGvPvJId0rYMra45zNAg3ik+UTnene3royjMygfAh8FkdI1TKkzZvz1tJByh5/e3
mUI0IXQmsuXXtC1m4OW6+4IFKyepfRvy36M3UdWBuLphY28r2dsUcd3UCWAs6yYJL4MK/mjMzCOa
pqS/3x2lVsAKCactUU4DcUzsk0cPHnz8B5hOW1K7YffirfkxemA+9HSmKnwiVzYOTgjL6v2UIUKW
KrqmqcV3q44nnB4bVcLL2T4FLser8HAK1ex42jAOtR0ajCUGXM6DYCjVy7Bc+XfWxzdDf44pNGIi
texsUwDoE4+KW9GHweqCRjmyUoG6c7JwJCpw+N9UrB7PuKoL/D7oPCogl7GSPOyl1D3D64a8MG17
VRL9s6HVpn1wWwPrKPf6Di1Twde3dk2N6s4JrqQmu+gdowyIBrw1f7n0OSYvPLyqdhTpvTMtMte/
WA2w+3Nq2PtBdjM/BovO1bBy2X3SFKhUQiiUEocpGlC5oNTDIBT+nncwrixRdZ0KxvTGhLPuexyq
g44jEyd1n3tqzxIUx3oNkbMPs61PCTJkJAb+B1RupSUcJf37ha3nEIuV4SGs70Qo1HE5Mv2Bl0Op
Q3/6ER9pakSg0fdx3gTBobGvCHd3cYgNpjIn03n51f+QozXPKlQ/64LMfsGK11yvsd3N0cxXVuuM
fbFh4vVCdmp3UlXatI3AEkv/b1IGrVIByYy7BMUlXuHOBfQ/U9qKxYCuYGTFmxSsj+BDEpn2SadF
tR1QXNRvGoY1qzqTCxZY2YYz1hT7mgS13qw0CP+fdg0hFM5CclsqnzfceQqBEFP1B/iGhKcuwiNJ
sMej5K8neE0f0TalP7lRNR75/lTiuj9KJgCg25y6BHkF+Un7rYLU3z728O1usiZ4z3YWVBLqmmm3
sUKIP/wlFi6u6ws8diFuArBt38lnW1FjMEv6kiqOsZTUZ8GFz9kTnzRoXFR6XRUV63YNYPvHqFPV
6blBPPg0UW23RplWKhmYelnDl2Hg4ACIIZ9ERkI3q9N7AJgy+AUbXtVSkpPwaTExa9LMMs5ZSZDc
QgCRJiJhJUlnmUmt8jyI4iifwdBeojF+fu9dvPOTHG13ehHzlX9gGG5JqcH9Ld3+vfmkeiyD+fe3
n8+TL8nk0k02g4DXjhrjh8mTUnxCHg07/FVnxzoKrYH9ynT7WIUxDi1QCcxHrqIjOo3xucDvWMny
2JfVZPyzD2qnjtFmmwRvG3i/o0eTpPS7YmcSLVB1uXKU6M623ApB4ZnTEtL4muz1KDnvY9sJiZQC
AiBzjxNV/CZSXePtmYS1F0wXnEzHoEG7WfHJoEFQGPB42h1bWirNIeovgR0m39o2d28hWyIv+GO3
ezptHUZ77JrpH0PoqggiHZZvNiQMVzEGmUy5mTHD3ytgagKGQvNySoNEm51eVkVPINuY/4Up0Bnw
QuOOop6gnEpIMTGdaHbnVikLN+P2TNn7+0ztb5aQACkZmoU3S0gbyQwT6u1t0MZUlGbdDAOG44a3
iwiGkM3q2h5Vg0VbPgNVoaTzNtOnhWKsM0YPjsosqznZI+HtmF7VYzGU4pA1rGii3N72f/u7B1A0
DzytFJV3bCLp9hXRWYR2tUNo53bQkdclPPm2bDdsKRtIon5nK79c+GzYcmo4vXBym0RENrKMnWo4
D9iN7eK4cQCI7HvSGNXt9D3WFxeM8/Kb6LMX2tjOgX+NroDqCKnI5pXVPSOF3pnuY6PonrQVGqIS
dXg3iw5FMWPOMtIpdPD0T5yUcOTnxfSGzSij5kRzwdzvilF3PtX9cbf4ih3o5r0/BYbi65LlzXnU
HkzGHj1/lVbv6veVOH713+O1eVz2ZOqCOPz8XQEqHW1OZFSC7+QMydfCvKyV4DuY/yD0F0A9PDA8
pYsmP2KPH3aaJGFe6CxNYDHLsazC2042N0sFac3B/2RMxwwaHWzmXlr23EZxnSikVCaK7JFFI0RD
Vmtv6amUL9/jTRbLH8TsFRuJS8IeOj9nvFiAQTvZJwpEKfE4sV4KQOA3wwhzac/GhgkzNF7v46Oc
PRmrHb8HcOYxJIjxin2M2zuuTz109qkUSyQbuM+hVlVXvbGeJRNT5ZROCLsf71WMrPeF3l8kWQqq
WWGtBTLHp9Fg4ONBUC8MQH1BAvCSADcxN4dssMyBuoNCFnldLIV7Tn3nbRKPVRYbRp4so/yuvaYs
JDyHeoaHx2kpWO8lE6HVHdDa490IE+1013U5Hu5I08M5FNGirYXaRBxTYfJ1CYYJb9vNELxwVQ90
BHIZCxV+BA6bd7QVSAfUbKDWxKiOgvk/GZEI6I/VNIlcg6y7b+eJ0ZyMfFPr2aM2g3HnzyZKkv2r
vu6KmyrBO4mEPHm0//6119bpgjq1bH7DKSZX7sSLbNpPpoTrcPikitI9B6JundS4Bwq6he4fkb4Q
oNOouhqoL8P77dFSn06Jcy8tgT3rue84Y1cdFiXrRXnc+2WvTxOVfIYX8l5n1nM20MGCpt7lVfjx
1ITJvXO3PYOLuhg2zzeWWGPgbtmN1fQJIHdi4drgQCMKLt/CFm4PSCZ0EEknAXoY5h4/k6In18CN
bLkdXCxy8J5mOJz17jNmS7r4Mx8bzGE7Vt39y17Bmox81MyYkOYNdBj5eCwXqT8Vh4vgv6rxc2DU
Ilxy/bwytYv2DDzBnfo8XOHFX4CTEUpqHer46KG/vA/VE7WBRHVBSQWiwfOvUXOGttL3iZY4VnGY
aVIdn6tuNbjIfAPZqaRFxOGY1Ccp8p7JtPSclJdaq3L037gr3uhJw5Ppp66d9hphetQZos4M+Qj2
k4YhtCqYlCy9KXMJeyL+HS7pxH+jlghuFg64Vp2+7Eb2siaJ9yJ4xvlhDG83XDzGUbMA9dXFl/zu
ajYiTlwf03jWtwecVhSIvpULC6DvyBGZlQIcLH3w7I+LsdjgCQxPzJ/8D+XqLHtVYzaywGrKED/w
QrFGi0FyLamqll6zJA3Pbmh//VwxigCUIvNWBQesyr3cP4+9tlCpCnQvM6l/1J7ygbeFMCNHjwL8
22OcsvsNgwF7su+ZvDHE5Way6uTMniQJEsY9OIplVL/zrRSH2/EALAdP7HrGCQfXBeB2LDBYPakI
myYPWTJuFLi3Z+vD/WQXRWfVaamuE20Pk44bw0XS9AWiDCakvNXRfQRcstalpJGqSVd+jCU4k4vM
oBiWMekI1pLL1tVfTt+ZY6YVQMHVryag7dvErIG2qWN+gbYl/yf8E+Eq5kEmqin/QovaQnCjOCmi
AZVdd9z8CMnM9l7cFI3rAr4cjHqZM7i/mw5Kvti56RGFd0DEUpPULDDuDRg1E3r4OLp58ZnhLH4w
YHqlbvwrCw4WDVdjG1WBidL2k/Sdh/eIrDXIdAdQTMaiZciyJKcEAUYTCpjZgmormTwqG//eavnx
U3OMj9qm7BSuASOOmAdh5QfjyL+yHjGKdijNXvYKNZ2qklVDVNKotltoRbJgIcZrhBKaWB+RX+1w
d4uSBxwe+rAHZ4cg6Aqh+T20wo5bO2E188fMkgtMkYROUypHZPVeps3covyW4/bTS6xoD0INfyQg
44+cSNgOjgdtYD830fIyMsI2jUBNg6aYDnuTEFrynyCDOLgzLorAlrBJmZbsCba0zU65BehDnG+l
/pOvKO3vgOj25Dh8gCZmPTjyCRNtHrgkXW8LzV49mbo4sGg7K51+yaKHPQHxU/CXH/V+rolmQgQw
Uref2GoRS3k8j1gvNbLfpwPX9DMsK0DhF+MSxgF0VZzsq0t2YVN7IfVch3+NBSB+1ZKRrC8abj3s
IjWRR/EoP9QeaNzVJ6cSL+1drOHpC/4YfWGTd8/bkws8DsIZIX9LnnSZ1YKyxrUdSJ+aromfA/UN
pVPCRvQF9ZGdO7+145bAdBAto3h5MhYq1Kouvii7qD9MFQ80m3/GQWJ4BF6m3lQoiM73MMn7obHG
+sKBb/2QdrgWpBISfPRgtKO6R44qSNAy46O0KygvA4XpO2Y0VU80LDQ37MXD+GQHmwq9FB2WKpew
F+QSuPFgYrck2N8omQRTLnJbpICHOcedn5wMq2o0uCAlTYI4WFM7OesiFOIllkkPTGjTbH/XAckM
rQzLzlXjjk7XD6gIMOFqrLfOEfLWFhbn3j9QC90ghGAfjw6AEag4RwU9hGD6wc6xMOuD+m0ybl/i
IoWq4r/RI29VTOZQ6CCsZtc8Oyonzfw2z5vkQaO/NWW36Es6hqrtUGyaXQeQapeMwMc9UBm7Z2mU
UvX1eY5i8MkYfc4vLWglguzsccdh9LU3+s5WIiebGhaNvpp9k2aF42kV7q+KqGoQLvVhEx+6qYOa
/GBMYHqtowKu7H/w1gNyXi7Tulvzwaib8c+Rf1+fegeBBiM1kw2cQarCTlrC+ezpp+DsXyKsvkXI
nMgdzIvyTV9QguT2d7miK1V85qSxKuIloGnmUEa57vNlwBL+L4sKsokrTpjnEMkNzkychYOnQEFi
GT6yK7IN7f4W/FArIZBROpoqxiP4L4x0RUVpTSpV8ZGyX7BB+wptfic5lBHJxDs9vwlEsR3fSQGQ
B3NW7AX2g4H7da5MooZi1r4bJsI9hjzGCxkGCuOOQdFq2/JQGCsG8G77b/MA7C2DEVWfRyCcfZ+l
82nWV2P+vd88zApq9vee7J/o0oQVmQMAZP/hM7f3m7hbmdMsfz3J8Youp4T87hNuJPV1bvJ1Z45O
LRvEHV4MX7Prfukf1wqvdD5pORDN4n0B/r5psUpeehPwxckN2cjx6nmD+NDFRPkoGLYSZdNNck9a
CeOFSt3Nz39Wj5hadsWIU8AGVMN5b5xcx7uris2orZT/Pvgypq5D9phsy7qjqDRw+MJgOfpbCAdf
Ag5ztI9wy1Tg1K3VZRR+1nVs/tEmEGwp2udBae/vx3nf5pJD7RLT+IvDaFc+ieGXtI2EQ7KO5jnl
UCWN2bOCxPKLjGB+CU2VRMuwR0yVtzo77KRP79Br16s0X0Su5UAQevPEsX5nhuuB4eZhneSmHiYt
ZRVyn0PernifzC4PcAJb41EbKhS1QUkaKtcRrlyS5nbSGoGAFqHgY9xAUIcSqKDL3fLnSxs9QAkq
4Wl9QR15QIVQdPJUcVqaWQ4JER2xxmE4Lxp4p4nuVQfaM9bquZ5VJumPJQaW69JdJpQZiqvpqGBN
BO/cxNw21vwJv4Iv9yfwKdoYdCb94hvPcOOpn4H4RcrATIZO4MsbSkwivQnVsHMTQxoEUokJMQO2
xSU/LhaA9JFjp1C8p6iM5J+A4U/HIWAzGxBP+Pj5n/UPIHL/mG5tnPT1wghrwoVKdBJ37+SvNAoB
hElL6zqtq3gdKFa00ZN/3rmKMFxJyzUUGnBgLkpELuZuSuQb7vvs+Zxo18jpNU7ATRBcEs2qZYx9
i3TyA4x/ASGFdWd678j4fjKaZyCKChVfLDxfaHwu9g9IzEZiwIKcA3U2gCpDPO0/bW7NHnF+6yH+
6DWwXeQzS2zensuKWs4KZDv8JHbY8787GWHqj51//JsUh1TZcg7fAkJi+jp149MjEgQSyLkk6gCD
Q3Xhusv2XLCrJ8O2RWRIi3gd7a6cxs1OxzQm0qHEICgZqjy2dBlmclW9a6vfYRpVNCYnjgssQN7/
N6eTcZgVHneScb/fnlXOnKjTXoUWUeVbnNDnSYjyRD3gzJoKj4okIWyOgkGkiRIqhGq3vwUzf98C
pTP/nFBPRJEDTGb2AyuC97RuXUPkft4fbR0ZUaCu9+TwkH6qGpESABb/cfFtHRvoPKk3GaHEhn3v
c4iqoxLyYpd3u4QB/CYXk72B2hqvFBCQOG3lISHXNGefjBXDydkPz8XRG+7Jq0R81m2FSeT4hrnv
eEx7J3/pBwsnxAMCw+JSKzSQ7a8Qc5CwNomSnQWvD2JI8iiMJNkJAZvPZYUhmaBHoVmX3pgGE7vq
QITaGpgF3fGhWBw+KWs3X4SRVW5MJ0zOnYr37MUdxrheUz/mKRNaOHTHIu2gE2mooCZzIAX1xCnx
c5AN62mvhq7n0IXy4dQXAFtJ2+/K4SSU7Ej//n8IO8egkasRXtmv2lOPV38qMIVRPGS9KlR/z+Ak
dqyM7nm7dfyCLY1NAbrecv/AzYUlb514bMsxTKa2Rl4wLYIw8p3h9uxK+zyZnTfOK2B+JLyskWJJ
1i78G10d2K3ZSbSp4lHRAQaJEWCyfL6Hdyv1jtax4fwyNcHOq5YG1ei8YVgyUNj+Zy73erOknHUF
WXnayhzVP8H986yaikS1eD9vpZm3uintLhZ87zmqk+q3YtKgKR1u45oLviR1pUH02IQw+rb5HX55
zVeMp4vSovnsPLtbA+p/RlnFgBcpNONF/KgcVP9/dIEJwNdScACYvaswtsg6aM7nchZoYeKp2FOF
WBJJtyh6AjE0TB9wfnMBWyK1gWfAseSeOSoc9ViqengH9HZbq+TfKfmDCZNpsSs7TMI4lV8s/74B
4hzOoHY2Merod29zLg10JTbgINvcvx/ptWiO0avsnAkFdCBL3U1RKKpuRHSL8smDheDQgukwzC0M
g8N4mG2Nc96lQFeVb2AiBdX+UX4Rf7Ti/fQ4btBuM3JEIA4N8H6EtrZLW50c08WdJvdyd/Gy2OVz
MPM1sDceeZP3gcBu2Cu+bqliflFLMumWkgyb04fm2tMCwC9l49cyOoLWRz42pDBp0OXX7QPc7NTN
mkcEke3q0kP3fwRDyN+9HeNM/2bHb53033XfDB6UtU6QH5qK1scUjT/4lKjNY9OgmeznWt8TKDWa
M/dpg5SyELA8ed9XUhDQuksfFLc+vrY6vlUqhRwJFGAitkOP/1U6lcLYSq17jHoFbjiuAOvZ6aX9
heNJquc0M4WK7q2ud6Z/hR/+idIidjK30SlkW9S5tm1SlidpVp6RF/2cnBWbJH3QeytBSFbe3YOo
xnbjzHVZbjAcFebce1WBpga8q5GekKxY+0c9CLApecDFTVqPjlBrBR1tx7HYGdxCHnnYD90fSI+U
lMguE8Vm0pSfUTzPjuPyo4z5ipXZzTJP+giZ7ScQ89kjPLd4mwf4a445MDyHS2k28QwqOaMK0+dJ
LTDJq3ASVhv37BkNC79OM9ht/ib7URabrDPj8DgZP+ccWK/4rlZrgvyMrbypKiRMFyusOV2xsWji
3UqRg++2Fg63VEGcj5pIoFMcx4I1EpJstc36ZRsFzhkBv2atj9lXoSCZajQp0Z+aFQ03weHdoGFF
PmwsPfiVSam0uyn25NgzIx47LJ0y9Kt6ZKep7rUR6Syh+c+qLueFOboek1uVfUiF32B7EQ8VYA/Q
EnV8mItCsD7RgznMZJJEHmThg57pMdFMsj9yldy/K64rk3GWal9s9fEAlf8gNBPAJHZpuIT+nju9
eoFkIo+zAyLIOw4I70s2FmhIXbMNeacDe3o7qJuuIocY3mEHxzIvpQrx/ag2NBJ8fD1oZ19aSv1N
SIh6EFkrCXVSDP6pHzNMc4r0CX2t6Su+vq5MUcPGtcr+MniFT6XGw+dik8UOIIq59s3/wDnSjWSJ
LzpvS5H273RNCgE/oWSrV+iRUKhlhBxT6T5fblHWDHs1f7vbEcQp8kmgooW8/XZNju7N5YcOgp5l
fk8sTpgcpz7SBJhO0W13IPdcwpDhWX1k9XQddwhEFhGmCE2eKly2EKzrqnQFvz972LoPk8sU4RI4
ItzFL3/6Vu56K51+5PiH89THgGHytTrMUMxwQcAzePjr3V1/FOffzCTNftU48TyDMpncLzBmkeYl
muM+HGj84JAFq+hn/ipHRUY7xz/McazCDSPPXhNY2oAdsSE7vZIE1tcgO79LfadAe5wucz/+ow7u
4gH606JqhddCmtK38INuRi/GMUnJ09j/9YbnHu8hC8w0F/5VFr+iWuZi7vizvohoEjuoRY0R4j/x
7/Dbr9fC79uN4LHpIFcSXKK+VsHiq6Nr9YZl5IQZYOC9WMLQc11L4OG5tqvDTnJVgE836T6G5cGY
PcYYG1EgwAAwEBxn0pLX9Pi7XdlTypP4DD6lwR8t1Yor3+AzQG/HyOgq9wK5XYcnzscCy6K2vc4/
f70KnQW3ByjyxDrEsI6bVth16WIuRpODk/pNeBcbll8NzghsRR93cW+OBxpPg3L7cANyUmpe7vOq
wvTPUKbErxvOINxmRB1HRAicw16IKN+3iCYLMdTrxeJZrCUyXdIezy0188t70ekspAvdsqqwritI
Lwk2S4/GFKL/hrhAKU0wepoFS3ydtEtVA1aaEDBnOqgr03duNAYITBHQx9FzEq6Q/sj/EmfL/I2Z
03RPcTagAx8xOLWm/yZhUVRqtgsKt49JZHtE9VUCcjgzRPXeeGnxaSMgN4lqmWezHE0jo5TdeIsP
sEYnbldSDs9caW4/BdyUR51D2QZv9nJY61VOKmhtv/ep6PQxaj787UuWRezdCexONd5HB+yUrd9B
GWA7ggK9mSe4mp1H+AL0Sbmy1Z3FF4TSJqfRN2F9S50Q/16CRam4jJ+mxERUGRj2RiJdWY88iRQa
xptgkNw48vUUxtC9CfBn9XM8xM8BObsTc3t3YORkUD/Zc7lHuv9AZoDJkcaRiNk0Zfgshb2TkjgD
IGWvCd4wAWj80kK3cPxsIVS60bMXw7rsmIcDxbrLi9hB+3na+ofm+nsjtZNy2RWvA+QLBeefE+er
1hTN+rKb0RcVWCBviEP6eCOUXLuWlviFiHHTrfMg5N0BqotpjzgfJhtE2dVKxlv+uZKWGLBwwEvO
/OKe45R+bG7okmuIeRw13ZCRYTxw9wwJ2lJy61S2ZVh2BXlbkznDnIlxCvP5W64jd+EPePEgc38O
GMXotgKw6HUnNoJqK4iOFMZ8JUkpvRhhSr5EKQhwBSbCP86hYro9MIixCoiyGFneaQOfpecW4D3B
fi4pmqKCP7dy44opt5gfkeoJ1wOMdMRRMY5hQygTMxbqM6SQ1qLg85uPyurllgLkCei26Qu4f868
29fs4pynL+pxZnZJefASJ5AhqgNRh6rsMmFvRn4nFJGCW9dnWi4jmeTJ/b6Y9N+MrsuSzVOkCV/C
0zpXseg6y8uB17egkR25rvi1RaQ3Mn/ZgAwjF6bBoYMMj49uWBDYn4gLdTjgLq4HyIf8cojoDymN
PW/+b4ulYmNKmYM+z7SjoULNatmD/v0J/8ZIZ4a4JFNQaVZtpDJKaXrQaszpt1tg1L3xJpXsqGqQ
eF4FhtxmSN89wKL8FmOoutIUiwgz+NCdy3AfvtHBNbPBFztzYatA06f+n3mpI2Q5n+AUA68gU2vk
97m83p+a/YTVaWrshlKn1NoAKp3nu8JQ83yOchuR1pvnHrzYcH9dN2bt7yYrid8hJVGbpZ5dWSCH
1qjwFrIEG6wmBAJg11ErENyxTlzeG5Vd15lCxGPemQp9t9KCgJaMYdUR2sml5I5uulvs4TY9wwCj
gCcaqwfUcyxPO6tda1xueVleJcwIEri8cQiRgXuU2oKIH8U06OrKFdeH2SbKgTZ9muNS+RCFJEjR
WWha2G965EbPy0mQZ7flSEokg/MbSQ0wHoyngtePTcvrtNeOIq7kFv0XRBD94Tqvz0coG0G0xVXz
iiRTcRevwE/+ME6C8fzxWbXWCSVJa1q1hhQf4LWxb1mB469WNfwZUBXOPGTWptCk5z9+wJDMITzp
+w28yUUkvhNZWhDgLDwqIlzLCnf+x1Abh4LJlNzezAR0USev8/U/PFqJobFxC9FYQpd+otvjgie2
2z4zRxY2fi//JNkBW7I4j62hTwEtEh27pK9qBrt9m0MZWZSFFj+GPEpnEHhEe6LJSbDGXsRPs6O5
UYAgNL/ztipx+YGFNROMZav2Jp6mC1ZKRyol/algwT4cEGXGgc55Tqbhbu+jprCp+Q0gPnlScp2s
s9G97PNONXdWhHoqwP2UzObSRjhJxmFnskSq0047YqSYSoDMC4BghQSVQ/ZRsg6Y+LCQNeWgz5HM
hnAYzuAt16Gp6OQZB7BcOFpgiN+LtDVxofIwubokH6A3OQOhwwoPyd/j1Oij/lOm/HmUikCu4Pmb
x0iJRKg+DRrDYGW2tqCcUXynnFhehCI4yWjKX9FzXTMYLga061SejNE4ZIHiCceQi7VWWiicYNPv
WFk7jMI48u68lYnJet7GaeMHPxs+xWaY4RrUgN3v86i+sIL7P+oK0Ejkaz1dHNbhYyCbbNCBT3hA
BDOMNHAuQZNBqJ5U5wKX/YBE8ddC3Hfx8gHrQsf06j73Z7W7H320KGWoTflvuaOzInDd2/4Ne+3k
F3DvOkWH37xO6PXjmsOONt5loWtwpbBnsepQgRBO88o2yOCfBYyab66zmHlP8BtKDMwCmHtkaCcP
AI/OiAQam7UhOXOUYWZ/nsFYJjCXtpzieVaQ4/7RZsrJSlwTIzFcStMOJMZ3eQj6xPod6ha6QCdK
q1k3paSvTEBk4XtJ3KgmiS0tzUsyihbBVLQr+wenT3n6PK39iv5dzbfSzOylGUKSbKJ6+CMqZk+C
DqjnIbuLO0sVgS5gU/Xu616JTCJlqit1X0r2tkpFkkeyh7wPyR+CMiHYeaGQAhAjVraT4lR6+d0x
enL9QCFW1i+85S6KSNRZ//Zr1TQqy+K6I1JpB696d4xNoJe6dTNSNFbNGPDj9FKRagX3AhZUsRzh
xBNnTA1rzDLhk0KfOkrxoVT7Fk/vCSerJY3VexnEE7QuwerLZYxVkUrKggXd84dTMjOmIW1n7Kw/
k909to2q/xFMjOMwLdtUKClToQFxPOWDGfNHQZEjwgtbRaYIwVik5sJNwLl1v+rFkUl81afNJRZm
UNgfyl52ew1qbG7PIBECGTlOGUWmrixXRhgJH1LjA6ZF9939t3JtpO1PgYLnItSXZ344Bv//hXWD
GQ4Cgd8OuDYbc6PAIhE2OrljVramMIDlLNCWk+tKd6kyhZiXvluebKu3faogDDF51Qk+vX1pQ7Yo
HYyN7HIMvGoB5JhqrtSoY+s8Mg2MmcWXWZGyIr9h2dPp1EY6xxNGrDTLHuAjzy0esZylWhJ29xBl
xtaOpyHfVPMabjIo3t+nJ9zB/TAT6zi0QEkR4733xbZBYEuLt/uCTdz4ErWdrovOk//1YjBENuTK
PZleI2VK56xJ/PaLuur0zVs8yYPi0JOhz4pB+kmY2belWx2kbw3F4DIPyab4E+Kg3ziwVXAmANfO
69f7qDZds3HL6l1eWepnxTAQxUaSP5Z3KKrAxIiACj5lSQVGnXYzSEkU/xN6c1cIshQYEJ3rs3y5
yvWJu2aBe3uDeWtQMLLLYgfIaEbwhsTIN1CNSEKCDhjji8pnL8t3DZtmm8OuT/t9kvicUv8ixSvt
bC4tFXdEmwahZ2P6/p10W1Ebao6kNd1eICLxmYyaIXFqF7cPKIeh2SUs63UgkzIDMqy0Z5/shdDk
B7rzJTZ5SvLXpeAVsL6guoRnyweTgivWj7uS8C3ALYVOZAbiLjnsJv/4OcQABtZ8F5k2DAQ9FV5c
voL/yBGFPu6xEin8GvuAw2k0HU+opiJjOsDteaL2kpkb7V3/u4AIYGAly68JzO5gqNB0UbUIEWgI
BxWFQfw0LDGp12l25//ero+xq2B7RrDescx9LY4LMbmR9UMepKHloWVTG6S4KGkeyxADp0EsXe+m
S+kg4igSxFwoKCqpah8cfs8VcHDR5danOz33RsZLWMPWESz47GprC8b3eZt/DMp5sYYXXLtcnOpj
X1R+Bquq14hTYjBi4RYe0G49kNykm7qQX6/fHc21IJhRi0jvq6+LhKuupFrnIi4laBc0PVN2M0EU
5C26l+028pZMhxZDqucNmcGxzJM0gmgq9JOxTjiHFEaydCZZRnTIwd7hVWmyY4Vjo8Nemq5USkh5
bqwTZh1qLpJ/N+8yfFi3XasPVY3aEKVbP42LQw47Prv9ZQKT09zYd4Ownfdud+hNGShDFmWn999Z
Bw6lQ1Yrz5vgwh8UEnV5dV1hwKZdbfLfyncaQ0+0afROsWwng9ywy/k4SEJ/gRLtovBCVNggkcbn
VEmY8PNcc8F6g3wdskMbvu7k0+yVmOrFYjip/mF8fcQZDdrRiugquO1U+16YLhrECvg0V/GGWWMr
clXdZelmPz6o0yBBuVkC86m+IqnkItydzQ8bUg9pBwd8olodhi2giaCYwkB0JB+jUhPrn2GEPFlN
C7WMw7bj1Dth5iSiiNUfEo4vPev0M3Hs2LcS5EGC15iHgRSxaKEqaBHRvyRhkfAUd4OcWTZc7MKr
edaUUWWkZ9YUPRKSCZBCdnTrI2H102k0dmfS8md1lYx6yzY7eeqcHPDOR+FLVoUpxHoiLv/h0yTw
IVG2ro31hskv3ey14sqLbDUcLouuyuO0JgHkDaANYuwqh3jeigg9e/UqocN4GNwGkr7hxXsQJbP7
HFYKQjT803dGpHbQ+yGKMhWplhscr0hFPn3i614jvJrUqI9+E1UwZBrfCDCF5KuYYRGYUs8TZPBF
jNFTzDrUkzLPHl5ubFAl0ntqCh+9kL+Ocm2rK0DPzzKbNHvGw7dDGbbInG+Qrh943t5CL8aL48IS
rYQ1phTihSHok/ivs7/ug8sqW1StXAKngZAjcnJ74VK2j9BRatAT+oRUAWTDXZ6Q6+uq0tzLOGTM
D2iMf1i2lwTPleb7DUm45Lg9r+Zbb7nCzyRHMK/C3yRePZVugbfj2+Go5JYus3myxv7aQzWYt9kc
TOfbHfXbqDCDUzOkoh7priYFjy0jRcSVSGc5oKeGcdRM9ostYueIVHXn6zIvy61BwOCZNXqppwDL
2ktGVRGXMbAsX22ohVnUu68TW/Q6L364UUqcMZNL6ZH2Opo/FuzgOJjaeNiIkk7gQ1kLo5Y5LNBg
KDn0DuJ7C0d6NqkAufA6/XDUQDn/gCERijtlvR4TCo+Pq3MYR0qqyqgd4nj70fD+S8rMzYyUrmwU
0T8LxrRKf0x01gVshTyjjhfvzG4w8Qx5oXYacgWneJfFhvCdwtmflr2FK6yFGu4ndPaTCfxWmL8i
Bn8XIaZlCJDLrRJhb8xWH7Ba7Aui6vFP40E3ZJGjhCCGpjo/IRlk30+539uaxWYBt/2RKcsoba6O
ZJuRiKDwuBEJJuyjq5AKaLknIDGlaFMUGSx1ockJXPOhXTvtOi7O56xwZBCyU/PrbsyHvrnE915P
0qx00q0V1cda3KjydjqMgI2te27+5DCWd3wRBpsjS2+XkDG/B6r5Ihq76poaWuPhy5DEmyivqAvl
568LFTF2M7KIAZ2w+viu/fGDo8npZmecGmvGuvJOVmMTvZksOryLQE2A0n4/PVSMNOKeyk2NGCj5
1EplvxvKrWIQbLF+v+tkETdqWd6yDNu9DlEtKbYBtPWeq2QclPOMwVMwgcaeIMEUcfpRFCAPi8+Q
BqBB67hHsdobyKjto2R5iF23d9YgtR56O5yqYFYlnYanw0GwEM0msWReNPhbE28rSm2+sjJFw5e/
WM5RDGSXUZVYadQHLoUTGVaL86LNfkYbyL0NBLthuZAhWpnyUksR4ILTXcoWzmY7eNoQG/Zuhead
G0/XWv88+j2wEkQjV8tsQvGPWvbiGLUOvdyUQsL8KF4cY0teGhy763fUIu5u3ZhrM/slhMmpZhX2
wpnoDu89uB/h4q1tp77Mo0d4gVy6BLHZOjHh3JjxR/UIWPq3nuh2HO3a405PZ5kXM39pv+sxZt7Z
9IJwZL+OKG5YZh5LeICLYUZjQetY5yUsUA/ehPmgMwzoes0EsRolef56wk5XCfOJFUi1wHDZTKw+
LYjFTFNGOjvYAa8Z6kB4kNeMhF7ted3BkPgHvveZOialNt8tVCkQBvaKMNrEyf1xkN9EZ+6SHG4h
/lgFu6uFHHkwykcU4LRPhp234oSPPjFIbTtNKNR4PwPrqKhybSJjkAztWwgqvP7dhMNuSbvpue9H
TbM0IbIDMC7xFJ+pdd139fLn8h0GIwekteq0GtZXS45a86BjxaGisSYgelbnWwrFEu/E5c4+HlX7
ZDviZdgXJnNH0rz3ugGRmt7S0zCnX2N13UrXT7ZMxDGOtV8hqNMDJhGZzeYux2ppPkvKimu9Tem0
v3Xwrd7ZzLwhOOmEtB0tooh1WBxfpW0VjFkKibiwYdPQThDHqf/PXQKbuXfA6r4zibgQu18FjBKJ
lcwGP5QEXsMyzE+b9aZDpsvreilDt/Bvd2stWz1b2D/bzg0nC5Qp376n5tFMndU8eU37yhzo2SP5
NNKMJ3Y4qidqcnegk/PoxkNrC8tzRUX551Ij/DaLRSlzE7o1pbFDTYyveTWrWt+vWMnZeQw9AYuN
vHFiIvvPCUM8Qe/h9tOoVuphfeJlofXBS/T/tzXksAzTSe/Lndz1H3dSanO8iKbdy0qaPxuhVJQ1
zVJbG9i3DBPR3vkThgHodxKC1wjRq9hvlasWxu2BHDaDPZz75UGeNn3Oz3kDGT4iD5b2pH26x8cn
7f0QHWZ82+SFFSYU1PWW8Gqq3dcUJ0Ur4bAB2ECAiVQv3tOPqEu6JhVXikXfZHkbxcJ2kdtvGeai
Jm6pgjQiYgTay1evLqqOMMsbyqv48+2U86XrWs5SzHXHp+BEmk7+V1dC8q8CAxePRIwDCmBsjO1o
Iquz18deHreR7pMZg/VPGPlyScAYShlxnPHp0bu4460HTIJ8Bd3y0Ccq7xd7xhD8WpF5lg7bONxx
9E9yfa7KHjWnS6W36sqqzEe1fnmFeBoggbi820lIrhFBbbzRxG5BjqleAzTU5LwmEEVo2OE1yzGF
n8p9qf5vmiribZxu3ezpamEFYfVh4fQgsC76zPCbFMWAssdTqnyE8GYgCIewlB+Jk0y9HhzAk3lV
HiNYHDg86D2zPJEahtGjfft4Pco3ZcgSvZywm6/k14D9ef7ieKq/erkT+q2+/lWdDbH9VD+J+sQ7
rIa+fcsXmxNv6+i/szXkTSj84I3sn4droZ7ysaeXU7IRV6e46qcq8+fD9ztD8CUCtL0t35nbvPAo
24yGlWE/FcYwqJu84NZTHnfI0iAt/MQqWzfjgJubU6rlfs57/9gYUTQNH3x87j6UnxzirF3j/uGp
h3oXIn9YfOGl/oEH86gteFkPg0HbSmJnYn9IlnwuX+4bS0EYuHGiCNIiReQAC2HnOLDbcwK8TorK
g8ecnNSwu8oSdvyTrpGBetkrcXqqmHOpQA89VLy+PwQfbd6TnP+OHV+n3N+saHhCkqccXWrZpX1z
vFKSLy+Cf4qB4t3pUJw/AcSDwr42GCe+L/nd0mBPrfFbA8nu97y1ngcDSbngU1M0AMiqbQt6/x3e
Mc/1wNv4PCKj1lxMG3fxAvzxM0YUDO1B9NrJcRTaJfZi7cywl1pld0zTQjr9wpel5lIBbsdqhr1A
PFjhXtQ8g3rwmtrLspJnSsMI6JUnkp1zhj3X3MoVEK5CrJfwpCRxIsj+vHiRhpapYMrTI2nvylrQ
75SCnTftIiUrdRr7pDI+le7V04Sxl0XVng/RLGC6zV4z8GypfSkhcA6yd4R2c33gx6xAvqkAgGIj
ttNe2SJ5p6VNCQRqEmRoq1f5iLOhTGmEZCD8YINIvKHWXnUmdb0rYCN0mZg3W3NYV9KSPRtI9Mw2
nzCbrXoa62dNW8arAqCDu/NtdghE9so772Jt5/iczaMv8CdIDa0t9IJpQEQsb6Kvcz5Q8sHr6/nZ
FC139/U7czehSWp41kkV5u3u4AldxDV+XidwFg5dvw2AkM2iAhub/n/MKw8gMthENHDUwy5JLiLr
lqla6oHkM1FNtnuCZUX8dBM2Fi7QLcc+AYXOM2CxX7FLUntroCwKt7WPTjetzZuIHATK9ga54p/K
lPQE4PKAkJ6hva2JABBBhmULNeq4goYps39/vOwDyiL0qI8cPb/D2jnAfkrz0n+GRdaynaiIb/zN
E2pz7jMpMVeTjsrk0kH/jTvEweNegqyS55Zo6khmsXhPcrzJoep/Y1X0Df1lRKeM8UZP5id/He95
aUkDV89ilfMpG6PBcHCvmy8rnwK+i2zUB7nj3cqO6wkfyNEI1Kg7oCEUGozmZnMThjh/qSoL1q1v
DKcuKmCEvMYofsrgtByx14I9y+RQENBMXHXS9eL3ycUMhbLEajbwvb0UQqbMKd/5pDhiIU0GVdbF
XQIMeAkiPFXRbg9i1yPc6oPzJ/UXgJ5LfEKTUGX0PWuQKp84MnW0g4KoqH6+yB+lCIE3MesfLug7
S7IadKONsJCmmat3VdwZq99tOa4UwmAisG/9Fu/0YZvxmrkuwbQBGqDMkWe+QUJaItby4r6njbiD
/L5eRUHhHnOSM+iM+fpH2QMgyTV/D9ZzNe1yRPMRGqhOFASqw6OZd6PQVfCMgeQOX/konHqSkHqQ
GcTwYfTw2OFNUAeYrhhPvCBIlINNaMzWgp1GLEdYLPfMfb+Lfa4Ao1Q3ZPsoeluoxS6EseulE9FI
na3yFXQM43JReku7CRP6bHjQRpw3yCj6TALaoEGOnKp20+Ti1XTcyYUuMm8uxM+6JgMM702kXIeR
Q9Kj9woFjQcsBSX5xloapTEwq0XmzrJVUbYm5wuYveIsuv052Q+Wf4G2BRr2Tu9RtrKTV8hJuGXt
F/gopRSIYRFiZ9L8G3i8zi0dMdPVld6G2jSXNtqI/8E58rQf7xGsO62OBb0Ooio42FdcKYAwy6CN
g04WtZxEp6czT+BIIjwkGe9A+SKbFwCP4R+XH2j7AEM5zwtqttGEPdwEXmbKf/hD0tOdeEb1ZaFJ
384wxHOZrcmmkLBy+LWc/+ErZHsq5GDSUyGt6uJHOrVKzazUkLPiNY8RACXpmbgi7mGKHmd+GhAO
qFiASv4quBnsODA/+GUcarAc02WTnJaHZCQAEpwSoIxAoShIYYaYqg39sRmvDOGwPlppkNJliWwL
wXXRtcx5ToabLdKlbEQ9Y+PLrXWFs43vb2mTiMxz6DqIIylmhXaSTmAWWdGP4qjD9QdvyhjYKKw4
iXbjbvrWgy6q6SUR9RddCZct+DnZq6M4IVuCITiSUY5FdCMvJXRc9KXB+4oMPHnGnnSngLfpFvgy
9uBhaKr53q4Zyh0TbtbnPTwKpvGtku87rNgb9Foa65jlBpo1/pcxmsFHXv+njXnrw9QQ6EtGd8NL
mQtkx8WFKFybP/WK36xFVat7K2K91SYJR07GQRs0Ik7wj9Mx4bdsgPhSWDLAvQS3zcNiZlVVmxNB
bQYjn1DuiJ898rZEU9wjogpNEJw7LPyHyKAZ+a6IJWS3qO7n6ycXselSr6CFOafJduzmpoKP3W6B
UQXlezT7+J9qGN5huzrxNGJelLfJtD5LHu2qcw7pXwD0PQXrM01+KuVVNFz70IUMzRJs4SQES0nt
IH344EkFV03vKJb7PXxPuCLQsLV5HTK3e1a8/NLHnkw7elE10i6MkAk3saBXBn9ZFcDrnVM0wCZf
RXYE9p4SB3FNybGOimnrLq+qcYATdRR7yTsFWPFs1Aq3mX9x1naElXFvPWlPC86CZqn9ZV4wpged
5v60pT9K8TbpsCccPiBtJ8zBhRvTus2/Gz4/NI8pTl9IhjiIoh4ecngayy+bJKzLCgfMT3R1iaD1
H6gi2B8ltlqUJhpCjqaDE+9sNToAGeKIzePyl6ZVrlqEXBxMsQkcWNUcbXBys9YVtrwcCHKzAl89
QPA/gl/piM3fu3vWYd2UadjCDSFMRLEjPUum+MldL03IpnLwm9+4WXBewJf22qA1JgEzNWVNlfHj
WdNozrBTTmwGquQLef70QgRY1VzQ6yTuPlBW/ztQuZ4tqyfY4Ti35gBaLkJlWhRiZRygVUIR+GCO
HV9wilT6iIIXzYu26NvCwp+JnB/0BeS3veYvB0BFZulc0pytnG+8ZNcovbXnZNLxIuflyZqsxi77
t0JQtRDy4giObsgTPUB/sJn/bz9IT5j+KDTmpQHdibVi0VGqQmZ7/DLF/d4t75kLDfH+jDo8gulA
ldF2C/OdiSfqQcqr4ED8PW1hsUUx8cLEarP3BxdwwdXx7TejZ9tz6vHBQcFq/lp0BiFHffXL0e88
sWjmo69rZK4oSzNGhPwN5e6VmVKiDvwUHjhfEoxsjiWNWo9mLTLyOFYrUL1/J6R4qK1VTw7aNXOa
INFYKXhRzCnEMdyjTnYFh3BdS2P/nIyWGhNLYJ6QlrSeoAInr0E8GDl64gmCPIs2pjQL7xEHj8hP
Ae+Gi0kF6VswDQcgX9GLv7QC5DfAF2/VprDGAW4caFystkz5y7jsZqIYH7IetlyY2OJjCQ5FF01r
xd6oyDuLxIDlfxMQdzum91cx6k1cm1n7aWA1D5V8Blea/fACEdhdy4OXhoCW41TaOzi6ql38NyIC
bnwV9GUQdP5SwJwe6kHHAKBoizDs5Jfp0GB5ZBA2DhZLD/ypKhnZ9TFTPprHNvr3p+d3o1MB1UEQ
DPXOxxBXR7I4AlFRySOmzMMZGREpDQXiatX4Awxq07V+s+iBfExx9t+EXZHBSFqxbD04bfH8UCVM
+8g9AhMUwTHaVevVJajxoRsl+SbqiM0qmGQb+hnnmxK1JerVn6mKwFAdi4eIMNmSGqM1VdDX/zfm
2h+63FKu+VzR4s9PU/5Mu777zfX2voIHoBbkDhsaLz1WvZcblgoCjl5Nr+ngylLziteg7C7qO3iX
7LjSxEVZNDVqdieADtqY/cmWyjhrcrNXz5xQdMTkSGK0cnTsumz1i96D65sG6WEFLP147L+wTR/G
x59XmagAyHqnlEHKa0q5EU58dqZl4HywVheiy/slNZASVLxa36DMPAlZN8c5XfIEca3gcPHDUeFO
inTLPiQ6m9Rnofpptt8CC+oYxp4SzBlhzg9ifSJhixUOCXgr9wyUCUvb+7BIq581VP9w6mwuxHGg
rgn15JzjHpKWFLlazA5xq4R5MyiGlMizSaqRBrA86ES7vSCjhQrvgT2ug51WvgHOGvSzEfB71ToG
HidVkYCVIzA9f5ubkKJXtJtB1h4mpqq9OG/mPlDj2MWNTSCiRSkboH3+y6T3FQxb+dASWS8+FXN5
NBLy10/g6976USBPQ7OzXCWcAJhSWtLMvMOvD4kj2N79IajFrZDPze9VyBEsSu/e33DzcE5JiB14
k8yGxMCE5D09PNV2IIhGAwB7ToMQGGM5jfNBWqABVWW/ezHEziZ01FI7AKuJjpYYvkyAZOSiHHHl
nh0zeGhdlaXNK102VRXRPtfnEcV+1yAy1RMeVnq+o5QRhdlU8zkwoD1WHyzKu0BxnFMfm58jeJgY
FIKDOM6GLtSvMGS4YISzoV4JDG/E0pyyqFqIuKTPbgLF8e1M7d/pFSV/mZx787LgKmaqo3fZqfib
uh2dX4yKqWfSIRzw74nhjlQYKNEfleYFevyagJj0r1G6RgP0NXDx58rDi5zwSjbzEVo1M6mRczCV
lyQheDqCiahxEL15TfPK4wTLahWbSb/OSJKSDS3YfA+Arotr5pK1uSH2lUaBivvqNrsNAyGV+6+K
bnRNKJvyvep29AkW4CifntoCLFyOZ6Rpj+s1bkJ5tTQO1k6GoQLvL/jD44qnG0Sk0tOPOTYdFqmg
S2ZnW3NTpU0Fd/yyABK958i4HhaL0RxJjs/R04wSfMU2siNxmOCm6vhrKkH+zoQhvMoGkjoNxRK0
1yBlZ+Xdk/z9o2QUWI3K3bL2fBOTS5bT89zKjBtUNiDaDTffHGRx5X6P9V8Zv4IiVmXQGMz2/nt4
ll9htJ7mw0EpPXDN1gfd0r2EzhiHUL9b7utRDtU8lK5pme6LgK83/sJW3BZlSRFymKgbYdA+xciN
NXtQ6/duXRlJey5fESuQlXo3XuvT8MHRlv+Bahkx7SHviKXU/oUDDEWsh0Lmy261YQcN+mdM7Xyz
giOU+HhDRH8BHGCbths8eRpJtjpihHHuOHuVBab/NKDaoB6HO0c45fGgj5FcHM+8ct5KZmebcz3H
PS4mxLdMRec3Mv12wAwDhei6BF0NUrQaDweoTemP3ZbUObJe7YYxQ8he8b0MNvPYpZnq4dGK5WEr
CuyWIzigtGnqnduDGoGpcdUoXZ1AZofEb0pbsR26nL+Mw4ehz9EsFRfaGs32ZXnEJ60oj7UIoVOM
oG5akEp6dv5EU2g5dO2sQJ8d2D1hXKxsjdHunjADUbU2nKY960FT8SxKXD5T8nHsVwcURoRHNtRl
G8HkqKBtA1NVslRu+SNtBnuNO6Vrg1NuqsrGaGR3hxCWkA8D/q2lgB2IERsjsFAbUnPF2btqVEmY
QDoFOzMjHWC9ep0+0i4fpS56MyeGh2Re2MUyFrU0STP/g2l3iRB6eNxzE87DfGN4VVn/t+bCbh+/
2OB1clAj3Vm98qj3dJ+H3tpkvrD6dDt3RRvGgj1d//z0zvUZK1CdS6Jjz+O98odWha3ksj5+7Jah
KCktMN2VDbZk0BfkPHlMWBf/nz3jV9Rck+0dl3za+1lHnHkuluY+K+rNmBnlgpJggrSsKG7Mx/bQ
S3XJLC0pCHJQqFhiod9DG/k6RY9yfpwQhKSWm1rgRFXGoSsbqCusU+5bY8jq7gzzz9UQAS1ymOXU
7oKPto4SHCHDnsQy8qDwjiBtf8/K6G1QHg0po2UeGL0F3yX5ZE6jaYuKO84PghQFIulq+yArW5qT
DxSLuFeL6ccukeB29M9UxcftnkV42Fo86eNU/FQWh1m43dhER8tacaoPiNxEywPF7JOXgHtya3sM
H2JqoAWzI7Dptt+h+gKbwbZXmNoJ8kUuSutBCCre7LnDDxcAzDnwpYRuwOr7ZuVuTTYIiP3eJIt+
UpPw+gAZJOzgHBf2+LmGCs0WcSNXqQiGN7L3MeDp07SJzDU7N9qvi9ZUyWN3A64njogGVUGX8HTS
Recb5gDcCzlRu/VLvLk9kE5XfARP2pzj1xd7rA5P5XRiAo2q5+hE0EjEuyT/Zp5P+tcCBeM1HzLZ
1Zm6R53YgOgy9hO72DI2gOITIS+lYcsehF/80/z9nu40TVlrXAQd0Ad8UekhLNDz1W+/1KrJfQ45
hBBPvqqzAGzWv+KUt6jMYUmn/ZyRV5bbdx7akmWwPzkWjxwYhpjL3hDio14lts3053+fp4nnIPkq
nOgIF71whAZvoN8FNKApyzkV6EU81tmc0yGrnFxlTK1hnKJTHO795yeD2bIHAw37ccnfmYjAkfQt
7drsQkmjErEL4L7V2Uco92YcMx6LX5DUd1P2YMBBSCncLxS8XX5vPo9fUKLgVsKoebi+kajBqhva
TgNS9iAKWAR5WNQLxNG4Mm/thfYv5myVm6zENuPNfAtzBF/sP1vsTBcl1VNYVFNZQY5ztMk0Ld3f
7uY6U+qYHVcFJuTnZGtAvGRrv5jcqMbt/mvWchcEfCD81j5PQRlXG7PpgCboUHNHOi+F39+TTVUm
ST0XAhDDIbccNyYtHMKK/CJgIgRf/8GTt2YAAcC0OcJswzYghNDzZ7Vc54inVn7oBMIQ+OMO1UJH
Vjsh8I4JWIaY1oos8v6KuVFnZmm9hYZYq2PiW1py8P58kfhx/cbEO8K/ws1tg1RXc5PaEbDyz22I
Hjmn+fMF4K/GvIm9RapKpsbYt3YiKO/xFuqK00stc5TzK54PF5kkpLysCujyiHza83lVux9ztesH
UBrPuBATouQTYABzEO8Y/QaVCD4L2cT6qPO/dcaXHrXjLvjXic11oOSBC3IujZG5qoMIyZwKKlMy
QjDcHsgGhj5UhmfEDBjPN5WlvQeD2x9wW4v7d4Y/BNAmnTPw/sRVYYmXYCKTsedZtUpORtwsBzeF
mGkC61WSgV67I0A6TQTjOFr6e1618chx7uUbdYkjCMpGEjQ9ixKtn0HEP90L661C/16ijU0Ojbs2
gD9SoAOoCJD5CDVUwoiSmsB4XFALT3ohpdoDGNIPynYuHnAm/NMvdVf/YpqppAG3jdBpcIxgEqqW
iPG9UEya2uIoWkibtlX2bdF3DC8Hwknw1ouZfhHCZbXFyDJ3r+FNzVIgxKGAcnRvm80rv16E+ti2
IRAf5hrIiUvTZ194FpPIsbSRhhBjyNhr+/y4nLQeqE8bCgXLSp5cDKOC2Yrlizho/JClhMvN3P0J
pTyD8xpK9pmNT8Rq7wauWPDxqaaiEo7eXpcjvquJZZTqJvbQsYE9woVLjkCSEb3bXGLp4xGm+P+b
qHPq7PmRxqWzN+r1CF9Erk34GC0CMv5wPj6inv+oOSsT5EDhFBrPFZ/Jwb8BSh3rrZO2f4x5n1Uj
pvwf17eghFVrjx45MTA2HuY/QDGvLsRI2NltSTAwbpWeLscLWE4o2VBYoR18nS8fFUTRPpySS3KZ
NwajMX7QqbkEvs1PIV5s5f/GEDbHDsULzMKON5SIsY0krA0armtN+GOyMhaqs7XLQh1AeOEQVhgP
I4v1SH6nvY7U0ChibcZJeR7P9t3u+el0RsSQduJAojCa2oB2o3AKUDnm872gV+79VerryPg6kh+W
Sk39d4b8Nx79tUB6htSBLzyXPzhV3HuPOL6OP9s2Po1Hc9Zd2z1Su+LOCymHFldVW8DAimqHni9Z
p4uT7xsSm4ui5faPBp8+stoCFeHmTt0kryuAXfFEHXHasi3rgl+StVjEzfJ2NR56NUqXUjRhbrVO
uZ4g7WOih0RLg3IX+jCP3PzV9H21dyu7LlbyBl7q+P0zPmBN5SLAuvdAluTxHCKg/Pduja0pHlFV
Xn5RIvpQTOTwLpZlPGKBrkbgmfSb5Vuvt104YRPV8S+/OmaaZbMusJ0OD8ZHNOx6wKxWaNGwAmb7
fLhE3ycI82UC38PRIenBSXhqbwc2+YcEuEfznt3Tv+3PBLQ4h0cv2wkeeSa9ILpCbbUKv+kqwZxU
+lKQ9fw8RdVxNsG0SbEAVOj6flTyi1iWc4DB+UEChnQn+kQPxPqXKH8TNpnv6otKP4oS255topQA
x0LRf4wvg52Z/7L2jtcFmrIWiIaLklG+ss11j+B5vWh51+6uDW0F3jeQ70o2GIAxlpWAiI/HUkQg
Ro5E38kOFFbzY3DzeNRH88sB6BAAa/nkIcdx5Mh8TSYVgucg8xqeL5LJPfzR8gpon/eUgZHAAiAm
/zb40fsV/kpVttoByUdXE+aT2Kz0ny07V19sXMlr1CUSy7JRsUMUp7dCQA8ZfaS1LT6w+CdpvBHZ
KHVabWC1KLi2f3nFBRbHh3YKOULr2S+G2SYDx97ObyBvtNEX+uy8+jrAdSz6z4DboI31fe7Gr2xL
p+2gxJvDZ7t3ftAVFV5yVgaukfqovuBwfGRlieD/tQz40emCG3P85q1lFK+eRC5RcGt1/6YiKysm
vnfKQKpZYJ23T1Vi4rFBK5s4lNv+AF6z8xUYcV5aSepJ1Thbezxn8FcQZolG+7CmtxJq2nSZHxjY
XF0sb4NMVK0B/Lnp0YUeLZkSnFiX2fwsQBnlc5tS5c/1QzeAks9P1/Jh7zh6uneKv9T8TPuXDo02
OHB4KL+41jFE61uF9Gql6dWy1PkS+mtMn26kfKPc6Ba9jRj9UtD6x86Ejw+/AoK6eL7+Y1eTU4/X
eD7x5ALXlIeoS/zSmn5VQB3UN0ks18PGrKzzjazowvbb1KCyWbXGAOl80PTQ0RNPECvavuRnUAPW
TF1YsC1TZSFMV+X4KUHWqQORImmn1i5u9vPXl4EV0BSndF0vCyes0+TgUXoJqVt26Q9khen7IHR0
trWSDQXBnwGdCVL36EmP8h+dVmEIgyo8vyz3sLFkgnMdWjncvf5mxXfNWvAYKy0IMyFA/Jhnhh/a
jLMXrpofi56tkAXXjDItlTZuVuSIgdqY7nR13/OpXCqpeLp0YuW9VZ852E01kRzIXm5Rc9pOLsXN
f2/BC1/6BBLxcwnHvze4swNPvv5Wpjw5Nz8Gs1i7siwkI6G/eEQ2bWtvrRe/olikQOdyII1OCoJK
C9XiJzbwD+9YfjiWWbU08ibf5iF6Slr/SwPK7dS//fkzoFzkHk5tZ15HgfuFCqEQFtlTOBVT5+mx
K4tEzislf4DjAFt7jZuB0k8wyYiZStlfMeOr/60ATXkLYDb7A7FOFU3+gfuYr8ewkSuOaIbx4gRa
oeEUvxLfyCkiFBTp2pT1a0mD0a4CE2FzmIioPaqAi6tw1NZeRCfEvE8Xtw2e/Li7Ym70rkPaH4gp
HxxQMrCVeRgWPqHWdEdv8FU9ZVlGcJIdifAwF2uji8JDq3yCYvqmOJTDWNU97WingqdSfcjDyWmC
bWfpIQREYUSHy1qSUDDsyoGgih8eMLNlc6+VY0NIpecJ35VIWf+N8HuG1KOnsJl5FIFu/Zi9Fpqk
fQOL/9S7aAR/+wYQEXFhhuybtbkT/zbgpQ730uVCqZr+BA0a5wZgQsPRkmgkV/5lGqtfFTRNCYPb
1/NDtunIRmXJLw40AAdseUbFqVmuE3D60lUqMqAo8DSHGGCFKCodaz8qyIsxrBqQOCUxKlaSr/3B
s3kbti79om4GZOtUIM+nJAtBYHXr47pPWxZEl50uoGGnpG6B30GBDK2yIqfXarczUey6NTZVRJp1
QAKsLWDJ1A+v22zhHBW4mgVGaialiNvedXSmjdIvKavEN2ynHtmlwH2V5uqSq75gqQ5YVCvLd6e4
6fFi2wiLbMjW6fnMJVrz3bRqhjpu5B9XHrC7u46tk2RUTsM6O4t1sftFhUF0TFo8ZeqGLLfJ6vPR
/90rSStz+cyefn8n1c9tP+FVIQS7lKKxZGOSEV7F6bx8+e+xMoL5jHxN4lTPSBbN6zFlxgyVVbsP
cYpA0hiJrVIWHk1BJFSeayePITjxpItTR1CPsJg3iSA0z7qyGBTrapUN8sLhsYDut4/gAO5Olugx
TWOnrtypgLoc7w7X1PxZI0Vco21y6piImcfNT05DPKu92oT+CiVNcPxiE4SuoJAW761CvlYKOPi3
a+4Q4UnSkBRZPcFtv1Kz/VMp3vR/o1KeZ/ATbQXUPJ3KHKxKUNOe5hrAllWHp71WNzQlQZiRiQV/
VNta17jYrIp+PCUuAXiENhnlGd43XQt8QRcUfLXDCAojKv9LXk7YNk2zKqrCP/jAtTt0PfpH6mnj
afQZwVO8FZYRV3u9/3iG6PBuepwhEwvqXY3JUsnsjxbSKWjg023hiS1lsEPavegFuEB2X+D3bjoq
bzTlfUq6TTska4CDWJHOCZCiriEn4mt4+f6sZ+ZfvRTlluT576/cvbIC+YUHqZW0GbJbejPgzJ4S
zImAA6q9JtViyTYCoKPelqEH+kwgEBgfiFeH7ijzr+l1woIjwqL3iAs38VVcKi1+EeXIuYuKR/vU
Kb9sJwpdGab00Y1Md+VZIK690/jmxzhuPFWsx61+bKVgQuipUKcjFrbajs3vvKdozyvWnNQHbG0P
EpQG5GFKWhbBRXAN3i/v4YadIVAJAF8mK7mruMR6fGv2WE1EAn4cNHEJTYdiofs1r/AU+hR+ZzaI
MxIR3M+VLTSuAfCrZ5Y36l7oUGotk7OT1mqvmzPKGHLk7l2yAcM8RjRcBKy46tjTRFf1DA94Ji63
5riFPQDlJ+Y8HwzYBLQ/guc7RJKXKrywPYBDVVWsFhxT3c1x/FhMpLtqiwsG/E27/1xcBcyJfjVt
IDjsuYJbbEGU1lYVq8UNLyymTT5JZbWycuZNPHx4qVbH/ZWJDNsG05n2SOrMHmrYdZ22QG2j3DJ2
wkMxkVkmeXvMr0j/pqSZIUH8gmFle1eyHqK2Ve5+cdUuw6Ur56u0jP/GoX6HA16wMJHKSd23XHjH
47c6Y1K3X5IOrPPi2nLRkMnVDlgdT4G35sxLAe/zoZb/IHP4TtThXV7NXCSw0pXNvvy97lOm8DfC
qXaQIad2lZM5TvOWbpAafj3I3eGlgX+rM4/bflF4D144ldW3nW22nJTBSlyTe0LsnZGDO879w++q
PENdf3PFEYwRj+ECLhDQD7hLIs1nmHs3uBd83PyK2IzcnkQ0j0zxrjK8cuSEwNp79TKV6SZtOmtv
oIUBAYsgJ+hni3BxVn8KIDxokPx5ROyUWH+IdUK3XJE0XdUZZE7ad4CBPqhogLDdB1YZ3ry4zArz
AObYj5+/3owBbXQgah9fcJulJZrZYoY7AHYCeLjwSuOT9jKhjI2RqcShX4C2krsEoX42ZbbBpqwQ
vSYvrsVaK+hUvQY0f14jhYUpTj0aZSyfQRvfHzQCd+vBK2No4CSQEuUvSwtKF09dn8ZFfbXdNvLY
Ev8Pi3okH4Xfk4xrAQyUXEwpOCLPQLptdsHhKn2j0frpTZvDxHJPstmsI0n6CUsZpLu3txfYPZht
gGGd7+Pinh7ezH1YLrAMBdDBugJeEnc+B0CZ4v5SknBjrcNki1Eu4fopjJKLAfQrsDtUrPkrKUgV
6YcEd04uh9/BVkX3fZeoYYaWOCRkc+ZNHj4IpPm2nBfvY6W7VjZunfOn4iHKtJr185u9qJ2br29I
7odbDhDfesGKB/97iOhNpkOrohR48QlY7gT+IF6W5YjD1453EO11nf7pilzgUfmHu2TlCPbqjjei
zxe3g6N3RRq+MfChnNWPGoBJvcLmnVa2cgN4EUBITGreVl1njDx7kEBa+afK6nbAJMIWzwwF623x
yQP1GOcZOc0tHlUTMnVR6cWaNZcAioQPY5E9laTDfx6u7p5XeCK2rqzz/qad43s65GqMCjRbvoU+
IHY+RZ9me5D9GpEkW/r0WzVhWPd/yYhNVcd01MUg5IiYwwXqB+qTmRs5PldJL/NMD5MErl7+ozZX
hT4q4+ZQ7HwgyxY5JxXixjsSTyr3wKIn2Fm0iCzT8NsvMe6wayWR3PAkxmKTjWI5esHw4K3JGPh1
cWQ3wNFPPR8mv55xI72taTTkCXFjAoDTs7ipOXzopN//vkU5ldehb8ZY9NfYhCtXKveyTsVpH6iF
B93/tfjM+krNIXUjYUrnP9Dq1I625hEDRSO1Y1fHqtnsgkCvNEsUsngVf3yYnMC1EpPfYchQ18Ee
QmUFSL82KxwIhqkrqHzo0k1HEkNak8z8asyetW1J/KrXUWyNKADtcqZSP7iGDNlQB59tqZ89mWGz
9O4HhCEtsb6oJnvI566qTGoC5sSvK1rq/GfwakM4xwmuoqa3nifW44+ZpasbgtMEVxqzqK06d0zg
Jy+J99QJ3g9i2OUK0FZtiMZEKWw/EdjsYaOwhxIOLltjWQjxa6nTBlWBhmY82GbUxizaJKUbTFSL
nX+qdPL+IypT8tik4gWA0cw63kfr87puud03pUGUZBSD+3ZkL31H4C73PxOytxoejCQzee3icBAA
TvxiddsOWVG6rLMAP0l7tLIkZkUMAj67UG9J4JsIiWVh0j/HX7ojAl+BnFXu7UgsWJSgYtVs/Xc7
HI3MIaRzc/OK90BOTwjj6+IBeqLareLW5aZrYpdjDH29frlH+AEff7uj+8kL4nNK6QNiDJaFuBBN
ucv2ib3Y0rGmhJNovAwsNynBoSnveQXllYuieg6FBuVdADsOJsTN1cJs67BNNnsp61Gt3Kml6hCG
vbCm5R+hSG5FnYZkJZgorik+R8OAZedtqq6z3G1tQq2wtIfpEFDccBV6LJ+nsToMdijzeSDtwYts
BYIQUcj3m2XIrRpkh+iuXgxZZVB+rvIiQ2jmdw7Q0kVbq18fSTu6iB/rGNv04WbvE206CzSEKFLO
asRhZk34lig0Me9drGC9desC493k9+xV6C/Pofs9RCSUBogHbBV+44qKv2JfD1pVeSl9ekXjOlRZ
p5Q1SRBLxAE2X2Wm9xBfJ5Mfb2DsKwvmKo1oTomzRsS/6zKk2dLV11/07bvA30f0qzurlywk+Om2
AxzPSQDMWddjuQjxRPN4V1gl29Ht20nxEhztP+ZB4/JWmt7YYx/BxfZwHfJRukUn+lotuFdDw+Nh
7+Xm0ozKc5tMBNJguOA2wEMhOJFAcqIIo0W+Lfx/rF7NnYq4KQkCFOrLkYLzjt4LUgXnbJ8LIUpD
1QaPP9i7Ht8yxlTJ30S4mCzQ4bpLB0JOgnKNx6UwMy5KnIfNwP90a/GKs3sO/3eEGD8/E9WuIeqP
pFfM7zXLxbmONjq4iWcwUUcLIMksBmEpBiTfukMMBT7Ouir9Y+idrXnOt9vJH8OKnoc4D7sMCOw3
auCvDhxv+VCR9MuevblagwHIiZJ0wl9++N4sYm3PLquZVHq/E07VJ2inHyIIpi+vq6LZCkY1eWyJ
jUAggpoHO+lienxW8PEOHmCenv4iAegkGt3oHHSXxEhGMjYf8ne3JNbdmViVMGNw80G7l3dLuJd4
2vWWaDG44lFpPukpcUQar23oiSmbYwAlQOjKzZ8AcNaI26ypjrbkTEKl/CT8C7b1lv6lhuyFykDV
Ep97QetB8zxq6a5aLCR1RzF5Gijq64cC7KZqMZl3hH9mL5aqnuFpzSZllVjc037RRnjMDqEoxo0E
O8Mc1h95D6+Tplu/9NB9GufcdnEB4fGuUSOnSi2gTdCvk30roweORQDeLlehXYs6Cf3dWEWimVGl
NNGRgteGdFPmF3KE714W8cpECXBWtHc9j/Ns1zcmzyU6VGc+9+5c0LFUp7k900lR3kB7/SWsivgl
XHf+3QA3gq7MWLZHvPTwX0gJWyPkPuiUEr4KOvHCwUFf5ZrVi01YtEEY8/TaFSgdAQKul5bxg5Mz
rTsuEjJzGsC8iQ2bJ12n7iYm8oXdGWaCmRyT3yQ2H6cKscmLH+ydZZ/8V3TIC2U3FWOg+on/cT1B
X43jKhI669j5H2clHfd5VPLcUAJ16gLbeeYAI5t0H/FmHzwwoTPwqo6QSTUD0pfuIub2cPeBqK79
Z3xqP0UjYDhIhCocLbVpHmF8nL5fvpW2YBfs14nhdNdKGabgLDJ6Kj+xjtuqou4zBNYDdfBSk7UK
Qa8bgRaU/LUbORZGPOM22Bz0GUVxYLpeUoCAuukS0ThoZWgHVMl+NfPteiLus7KZMs8DGqrw+ehk
HviLOIuYXT450WkDpheseYE9NOD+JNBpigdDdi3+pDqbb6yXW5DWng0CcNdOzDt/7UlpKrBRHKDc
nZnKPFzO9aJWX5eAFCu7AsQefSFPLZewdiHZc8ZZM4TC0WXuVMoymaS17Uvvj0xm/I48/RT5qYMQ
eAEHssKdSeTumJRxnU8FmfNFqO2oCKC+IOEnrhBKHGdOtJkujypoSipWP8k81j2Hk/SqlQa2SjdI
k9ArmqfeTDXAbuxsu1c4wBIHR4edOfnvtNnialdcsvkGK6DAg9B6D7ujd+rSF5G4XH63ylTzUnI6
kTbKGv5wB5G8GG0CdCiIXfDSUgqjWlDxeiuPZG/xzwQwRd55nK9++jPM/65t5o3zZtvu5I09HneJ
ABx+ytMDkJP5MQcLpoj1NdpKYnJ68lDGvg1h7G+UXQDJ3k6YmThvWhmk0YmngTlLfRC1vcJ/EItV
OeaCSDlwRrQ2qQBi9PMk1WiGfOBailFi03ltc/BSqaz+uqorfDJJt7NfmQyWm3DA0fdh7wgWBM9r
eKZm9uhxft6IDY7nu9mL7ltGTgmb1OiRroKZynFBU9YvKudwU6WAWYbnfYKYpvNLQvvJGupQRq5Z
00uAK8izWQdPf0rIw3xesoCnAwgrYRhD42y5J9kTXhPPS1c2cc4J/aW43rDV01fdabbwMvVgEwB0
Cxl7w/kM9z75kcny2RfgHDilyTkYVUuRn14XPisN/CQpusrH5omqlSwfYt6Sb6cQg+C698GwWyCJ
j9oou67/8r9uFuC+uKsUwGhodGFYjGNYMPjMJ7FGMWqdzCYZdPkgtcdQFMyJkMwh9sMifLPFbMfk
IKfQGrmauU3jJ22qtqmxjQCKDq+yeDcyFr0wPDLn4lbhLajXKe1mkEQFLolh9BQ+H0/OQ+wTigJv
nHf2J3B+677LlRfyJMS+vnuOpFXq6zf/cCtr1ydX3p3raWuw80+jdYiV/J6DGXFVY8sFT95uEd6C
EdFQESWgsdZPOkgF3XzpV8NzKCuImbao7cKqNB/3iMYkyX8IqR68fOFmBjiFf2wobNnEYtmbj4r5
T9+OjJKD+pyMl028/NcR4WuY+UwfH/z1jwPS0cMWaqxKmP7pltvID4EP7HdFodk8EmKyYCzBIZbe
Spj7WXCp3EK789iYj0Du9+US/XaaghBtjbUDK81Hp6TmiKFxi/D8oBPVzbISYrWZGox548FDR0FT
96teYHwf0TQ5wAlrRy7+zC7aQcZv/GzbDHgo7K3nNbIStFJQBOCGny3JIzDDrxkOvZvrxreS3/qA
q1gehONvJsUTbOXUe7fRudVxFXeI+OrDl0jOhAYiGAtswnHqFzOlGccnUWWELgXEg5KPiUafItC+
Aen9VXG9J9sbr90sDwU/IflJicRCSV/rBDWrrqeQ8QYPp3T5VS8XLmNrOdma118rDr9ZFC2kAWdg
g/MpBED1wM46Xe3vDrzQeVFpZjr3ApMJnSknch5//X2f+EFUkbG4cyVas7yznuhVq6gSAYTXwtY0
uMvfcA4qd/zMHnCTcDr6qzvLW6RoS/HY6cb1DCR8gDUhnKmn4R3bm6pskA3WvgUib2qE+7e0Q5PC
Jxck2sM9hkXTJPPDYlmapk4B9zOK9IvVzn2q01uxEIxCZtTvy4eF5jhlbCeaYVI146+j2Fsh+jyL
yYOnnJtYLdpapC2DNxh9BqV8x0lMXOpxq5kj7t91CXnKlMmZNubBwEwgwQkyEJq+c4qky0ZVdor/
GQ9InSEuHLHzaUN+4sdDlRDkea1nL9wsLNCLpvYw/FPvjket2rvZteoroJbDI2GQ5ntX5HneD+Pa
CJjtjKX8/fTks5D95gOOIWd39Fhv3g5GbjEDavbGVuoFueWU/UaJyCKjf2t8nEzVtoLp8gofsiYe
+pYTe5dao4B0nBgtkeAEDts0Of83Ch5IZQ7md+SiAMt0IgPo6ePHwP2Bnb8p1V2KY9RkKtVH7++Q
pdZjnNgFrxiw/5M2xwS+sDy+oLnVQG9UQO1d5LfoihrcQqyn6/H5fG4aqbs2AkQq3jjKUQrN8FQn
9nniFanqJMhYW7UzwMja02qTWaWEZ+eoJnmPRGRA7A4eADIc6o8vemvitEAA0YLRsRHHmQIRcqwx
fc/R6XobOzH3RyZ1b4BKxdDbZwwW93cCHuVa/jCe2OOWMGvgsor9MtP1OLpyn+K1To3LCL9Rwi3V
O/eEA0MQIajQJhU/G1fKW99qq2Q87sHtAkwqXBwQgr2qjx3ShYvsiGznFZuHYWSEwTvtKH8kLVeU
5OLZfzMsR0hjjqIP01eZCWq1whmP3BVrxkaIt1fzMaSKUhpodjUrSMZW2DwjySXZomJ7e7+YcmIY
+TSp3LR8OtbnvZbHt2HhJDxNlvNBOO5jV9cSZybz8Cis7v1EXu+nz9IXbmbe4bRBVa6cOLSXbuGU
NPYj1L/EQ57MwQF3yVJ9nFHrbA9mjELxOUDKDOynmuugs0Qwqsa3IdmsgSsiW4qVVVz1LDITMf5s
V/gH9cUouTGq6bcAitopfhRXv+goQyw/61MY/CTl2mjgsJFDT43tqLrDaWKriTVyCmWbh04PAbuh
zfZc7Yz0H4VCqF/eZffq/fVAhsgR9AFcuPdhnVCjptuUogkrx/OoCFXkzcP/BWDKDdbQD7sSCOPn
Myi43jG59laN8OJWFWnwnxpLPuK33sDc6m20++TxMAjrQdcbKGIwPe/P6PtA9fpE0ES8lJgIwqFK
IQhznGF1JkgDnmiK2kxD2aHhalb+hvbpfsqTGmd24JPlH2+3q++d2YkaMEFzwP0D1mCBQzqQ0Bqh
HmcaWjmQxkktvF3jJPonR6egP2Rbv31AFcr85k8KB2Df7ZN32W5DBgSNMdfmjxXByGeDWoobh4FN
HSTo/AGH57N2UhUshNtVEl92Bg7nQwhBXpCSt96QAzDo9nDZxwZ6mjbsoIqnO0FZt5i4UqKXqgVy
Phtr6mpSnC0T7Wj74wm1pKubq9+FHSwcPlFtzFcEdTnpkYs8ZiNXkqSh2mGFLhtIwiyoSow0EqYO
qTOVZ1OTx/Im1hyb457k7UcozuKwguPsVKpwCWvCdxUdiYqlDH8KhseAM/WJFKP3xO3ihLWd75hh
FGhFIKvpIfZTLIrvbFWAxvSwMz6L32C+oMPGY33WUxWZnmWfPny0VRSH8EukRC3UGKa1O2a3a751
KpqhvvuIdCzaHHCjUrsM/zZd9VW0u7LsuWDHhDFeubYbH+ImC0GBXpNSE6AEHX0UjQKJcR1WaprC
1v1vm3ZMq4nd5AegMItD0rXJ3y2MFzuNemUq5ZC4/TfhuSNypy50BKzr5cdJvhOX7zOaTZedNHyH
FZo5aVrigoXrfFBtZGcEJ3yyd2BEtaWeEauMIT4g8eF8V5IcttUAhcD5/GDwRv5ISQDXqo4PUZLP
PFotYsmBz1QtVakzP205Ik9HmrksJ+ZS5d1RM8fd9qrH5BoCUsrZgGUEs/QNfILxUNXgyTBrV+bq
gAVrBWThtDBfbOas7aNqQnWUSOamZC/nf/v6e5U+j8emlwC4dk30OHKQzxPPadC1yEc7C0IDhvyc
VYVvy9xUm4RXs5X657qFq5omBubssDZqPK76QGlkoANWPAC+/UdkQrjP0ZYv+PKmM5fzwNzIYfe5
R+giz64ULFK0EX7FHOwXx+Au7PWckIK+hhzQAGEZbKL/wTMu3ha3yl33GEBQ6JcmIEbt0VIDjnUL
gBiYgUtOquC9bfn8uRTRyqF8pY1gjrORO73gXVMKOqQ0fdKWD2rYrlHmadOg1FghMz8cNZjOO2gl
TRhq+zcAmYRkc4lmNdsEe7uV6ekj57CwpHk9mX2GYTcAWzVpJniyeYl6NfY9hhmRE/IM/ONSW6yA
q8Nv3/ambE3joCgvT2utdBmpWGGRmPlmx9NNvzCBTrj4v/Hny+llgTsjrRr4GfS/PkYrDLc3JdZg
15ZWx5N7jbLWsVLTclVq5CKx0ehnSBcEgynbyPX2yFZbZWdK59jN0XRdyRbp+2zeqq58u/TOC/4n
COKf6q0MJZ6aJPYk/iD781iZH3a7uVdpIxsvIwNFFrcvH4WfQ+Hy+sj0wuOlFM2EMNMu0BTzIldF
NiPZ/GYeyJSH1dZjqIk+AIfJyFtJ/Yus5I9m9RrFFY0mWXSRrfoGaLl3IIC6hHVM1JuERPTpufK3
PbMwu08kqbbhuhzBM0d4vXCyQ2zV4Aiy87szzonc1sB45HOIQHfo/ceZNi/DCGbuZJ/2Mg4Ka6cf
b+4Onpxtdytgp6yAt6QDU2sCDv6YV6ro7yb1wWiVimg/dCTBu5iT3EZGRUt6gssOCv2JkZVsHDq4
iey32AmZP2SfFzsDVTlu86tB6TwTKvJK71u5W0g0DjHAmA9oNwLTBTWcKhNPhx8ub6yB+3S6EOb+
tupgPdzM7IqfLy9YqCsLZYXBA5v6SHM49HCsD0YAPV2Tii+6ZAYP3c129ew+4DHBFHik/YvNRzAO
OiXnanCrV/nJyj2N9ACXPWmdtfX8tVFCSIpy6+lE73WmafgvBKyiOGUny4h2xtv9OE3ZJoJfOIzS
Z9H/Hs8RavNFlRVaXAEFYoh531bay/OOqKjsPTUtH7Yw5VO9HlLp5BeuOgfRh+Nw70MH8x3qZ9ar
DewTpNdYgq0FjE3FBgPj35+DqOouvqohotf99xO8y2gf8Mschosk16xTQE3ejW0KR13B0PIJ1kCX
hqV8tiMrnWGrOxiWCucKasJX8DLV8f3I6hxnyQ9TOsxPN/k9VomTUfpngahTL/gJC1AyZRazK5q+
w78kv25l2kZUlmHsisfkda3k5WIRwH9IPv5tefpY2Dc1iJR/1uxnUzOBwYIBC8hlqjNNoxpbFE+B
M5Dm7taoFwtuunxFp3+lkx0RvALZtvlU7E+M5nDraYDXNMytAE9AkxcKh0Y79QiUp/Y2947YDmbE
nGgN/BNoSo5FxLdkDs2LpAZsuK/4YkL+45coIdGq1FHk2BthhIAd3B5mMg8lVyA+1E+xLqPeGFsN
qKp8aRJ3ZV2UgyCmS8Gg4ZGAXmEC5HREgqZDN4lg5AM2jz4ACp7uG68wUiykQYcpBELVFbOBQZxN
CY8vS1HoXhM5IThp/tBPsNtdw4ru0ptlVU6HjzLczosXccqmbNZapszaMn1n3/BWfare9YPUaRf3
Ywm9cZzZzS6kxZ6N4t+dcPHycLdZcC7UXg0uVU87yRB4r+BvEDx6n8SOUD3SQz0AWXOZRX2iSWyF
kkKzUkGF31f+lFICG10kToxlgnI5vkXE05/HM/NqOSzYf/mcgOjvi21rh55vDMU7YbXPL4XlEoFH
Umm+cOXFeVDIZ5v0apXEfJ+hV7uMh4bQPuYbdIqdAtn33s+8HLxGR/YwxZOTvqiasA2Gs/2vR5by
RCE/eLyvFncQ8WsQtbgpeBzoqr4EzV+mnFRVafiNWbZk235HeQh4UxlZHWeRt9YRnhNXNPWPY9k/
fGhnAGHzNi0EX0dQMbvW7JuY1aGesfZCiGFvcXuJ996GCSuvl6q+1o39TXyPX+hcwbloOqi57yei
MrBlg6VbTZ02X2xP7rcL+Xf+Wk4uLlgg1VY5QvhC9BRJYFmhC+TRwZ1IpyCVztkZm/3L6jAt3+en
q1zuGzqRoDr6BCgFEwS/mA6ouqCIOK1+1S7kJPit5k312klqaP6wJF1J6mCZjYTQJ8GQRA06cOEA
RehLFcgKL/V2156WVrCQTYd3akralyseUoKdWz6RCt43lfrfeP4odf1sPprEPM3m9nMWU7ZW4KMU
mR8YjPQ6/rfSrTh8p7bQkmAZkvfusMrCcWOLrBohcNj8XcZR5kR36j+5j1eD0M+O5IYQHvFlcavI
OwzDP11eDSABkIKKeEBGqeAXtOdhkjKkGts0sGCny3+G2Sy7ksO/KGC0Rq1JtvjG0hqPJyvnKgIp
Z8JfIePLvyH4bMLIm8ffNXkr6qMlJdG1NTD9xNRbiHnfw3706KpbL4LmRMHUTrLCs+X34UB+ztVz
Bz2jx5ij99AaPNe8/4DTYoUcj7YjPydEDiC6J0j4+E2unBEwxMseJQjoDqE+DOVxUKNaTsMH/TNc
LGiSsK/GJ7VcyVqXATF5zb5S7nCwk1I7EMQplC+K/EwLDKneqHV9t/CS5QCY6KTIpNJ8WkHIDRYM
Yvo0JsMmlmDUe/MYoyFg379mWF/0MwSgayw49/7PjSneZaskvI5gNsw3PZD2ToiCl6MmFqAF9hwp
jXS5+odAbdfGcMuJ0KB293aBYuzvkSJk+2MOIcvu3DHklt7VuIxZYgHXqPb1unpucF+sA87ZxTUc
jFOz4dvMUFj/ogJWuQfYsqR0axHUkgV2IFbaoGJdMfp4DhCbWNLbZGQeFOrLO2oviq3aw4TSnIWa
/E98wRJPXRj8YJU5+8Dtr5phty3NmuVxyInJcifSGZcr3OTzth1xXg5GNUEPjfF0y1OD6PZWuH7u
bJj+6ViOLO8Locr2i9hwrmAYWTcqtDvYcGL1VKoGSSD6eNKdPVeewltRlsTfvh66h71krTZU/ffH
EadwdXUEAt8ifDGCgro3tuHzQnwI07waAO0OQrRwlgnXaIL3ykR7/Bq8SDBm/cW1g0sRnQpYE/Ds
liRsqenFHBC2PyR8qnI5E+BFMtWZGksI/wwGhmMLgKzzJGOpanwsa430DOPJ5W0bzeNrbkqYu6f1
Bt7mYYFO5CcAERZMeu2Gk69u8vUUhO5X+Hl0p994PCanPyEU7y2DqPr2CAJH6x7EcvBlLDkj4XaM
g5GwJfKKN5S5Cty/9d4kAmAR/rALBegulYqqfjgNsbXRyLFbMiDyzjcXYKGxD8qtBM2ewQC6+stB
I/eeCRkGV9vDMJhbshMroC03NDDJTvXhbhoc/nBpYu4qipKr1rf5Yy3OYsaHAERRAKmkaBsJeFjf
QTyyKdL5sBGj+AB8wPI6VgQWni18IcqgMGlxbHsFjCucyzSYMmFRunRR9BO9G77Q2V64ZwvP/yWH
dg3JkpQUgN7acIAMvxiU94DFyVCuoY4DbrUd8PWoqvo0CVuXyoJ/ZCoIqZU4UWL6Jng0ejFLJdw1
VbSfMkOc0U4fpbAVskgxFx8mk+BDI887Ozk/Yn0HGD3r06NlJ0vZI3GeQ7fXkHcokp86hGtSC8+F
kX9OYSGeyk2qIFXe/WawTKiyakNZ7tW92k26FOED3m2sVSvS/CG6zSLGpS6zsutmqnvaCUAMS9Oa
i3PvBUoEvegNWJdSHSaJ37PQRtk2UwRwCEbiFK2BzNqaPRxHJ1i8nUrz218xkwMRY7J9RTSgIb5W
Lk99iNsi7K+8VqR7L7slhCdbhHOX3NvPMmrpJT3POwbt1BBLOiSSCt1MB9rPgn7NwTUDtQe19IcL
QxfRj7wSbXDxHBAtwyzHrdM+nb10fZU9XH8bqXP8cRJduwJ5QrFBbffGrwA8zAe9R+lFlrwozTsq
ilzh+ad9CsU/lQH3W1GwbIoYvz3QKk57cbiTg5cOkuFEbYHeGvphlkL6CO4DlUkzg+Sp1xWki9Hb
A7diuE+72C3gz4hNXdesV+XdsdPU9DfKpKKs5lgkv4b9ZDf711PZl5BVLX5s8mjt8iQIIFBtT9r3
w8FJgGy2OL3zM1ZE0wPwatx4tyeRPe9n6QkZTvdWBsN1YCC4dZdLjjF7GXE1hq3N2gs0UnbIRYVl
bJc6aX4qjg1JmfMAnPBae9Qd/Pg3wf2PjLuPeC94a3eN90IfIyfKJSUDCZR08a56mcYgBXdg8M3n
XaJi+BMHptRDjXdX6vlOiwCG8aPFlAHsCpTNdvC5LaksQVoVDk55FKLl/FddA6euTkGZKUmzyxUR
sk1nNuuJe8Uc6Ug/Yr3ER5aU4+rtcSLdo5s6f6Qjq51EnMd5KZUaQVMLT57anXNJD9Xxyt3Phxn1
BM4WwtChKRBleGJJmV3OFbfhEf8XREO7pdKzlnC+hbFopSBK5n58JURh9+Sx9BSxU5lgYvM3ggja
fYlY3YZNq1rt01xZ/27L8Ibw2RDEQY7n5YlgY1k2PUH58xQlF9FE2DBLs8fWIzf7xldb/O2Lbgyl
ifA55HLJ2aogek6Ahk8xvO2KOERbyUnODPU3vLWAwjp+kFdltv58Y6kgZqYeN6naeMGxWyFAtamM
y3FSz/OlRJPDFZDR8kOEUilSyEpDRG2xoUeheEAlr1VbkhRAN2uzgc5XziWMy/XIyy4YPV8ketRN
9893H22x9kua3dpjw7ucAK28lHAbK6cp4dEct2MfFb0JHPGhe4J3qpcd1dgr9YioYPUV0JKDWs12
VR+jqwujgF+RWkiN0ZIZDVh+8CvwVkY0o2fzDGlDCGlrgY0WSxyVFjZPyjpfTz8Aqpc+0WCKtzfT
fFaHy8meB8MXYO3KVVQCcgB4AUbkofERI3QsSMOLxlijUFzN9P7w1g4yUXy2dlbvsCck3IAMMowY
fbV2jShfqxfKM+Ht67akToKGSIrZ1U5Bug3ZSZXeVWTWA679nR55g1DNfEC/yMTzoLwrqd58BVn+
1P/pCkNZ1Ql1Gc/M/ZOcOeI3cOuAt5gacI7V5T1DvAU9RVXj7tPf7htjy0YNRqdBII1NS56YIKld
6CJWItR0XCamgkXDoRwJOz7tNP7YkRA4BGzqVFWz2stdC3Z1w8AfnJsCUQw5mO3c7wP62IXqvXza
jP9TAMSOHuedMGXyKs7nYqV+/3PTTllek4YmPMGkzJdoQaQkSG/eQlIV34MOAoCmpbLKiOo8uRVT
0+BKjiI1V0ffuAK4u8iogZ1oO9iWKJyCn3M8OXE1vftdGeWHYg1ZGp/DBVU6exQHF6yGzrxLkrri
Xz0zEukB4bn2fl0zE1ryThBq04e7mKT38etnrSTow4hfD/0lKa97mBGei9wU3reeYbGrWpJUfK7e
VcPszcBTRh0vZl+/eTzxnCTVGiC2aedIp7QzqAKV1M1ZALCaJ/bezupc4ec+y3/jy3+IgLueZtVS
8G5qn5I28dDOPXWvFLbgKv52lHFj8dBU302LDPeWej0w+v4vnPPPiUGl0Zosq3cU1QtJfPkv/fXg
7NjxfRqmTAVu7ONHB0J8JNjVNGIv5C7MKn2lI1Kh1gpmnYiFO8kQNrdMC7g/1bJUXivMOHVFfpzT
pBQsy6taXO8RAP0PNzCsjT+zkc8gHJSjZ6g+X8obii07rkqdEFwRi/n/QlrbnCVoSatmyfrJRABQ
7PCz5LXR18bUKPYxu9h+JXfoLnn91Y6QuRE9BP+tJAxNONAFsoRIwPeoqrTnEVH1rGK1dTyhWBOm
argnqb7T2AMsC2SooAURjbnaN22dinI4JniHt7UOOHH8Xa0IcgCo52bLJnvILk1o4jmWOGQBkicJ
PJwn8C3sba5Aa+YisoogoxgTQP5qyHtKVP3Q6AbwmOyRXxVCwCQvEGXmO5yaLUU0h2Py0Lyl8yr1
qFrGR6ps8X8nzLNIK81LLQaN19LrD6E4Pemut3L5qk4CZ0bWtYBsKsQsthhE4LeltNDwjaGLQ6FU
Lg/oaj+J91RyoEZB4WWm7gfb0Zv4pZ/7RssA47fzEo7xcYRmhIpLJpfXdXbX37NMOTlo1HqqGBoa
13DkzBP7drNUWLFV2s3qjv3ZFEF/3eTYdGVa7qhDQG6AAF9GZR2oNqB9OHDNxCW15GZNebyLH3xg
iBuGi2sg4BIu4t1HNl1Lk9WoAavZom8zduPrjdezMdUeEQABZIiZub/Jy4rIAtQgbLLO+d+3ziJh
pnL6N/YfjrLX8faxRJiAREuey2A3gXtyTfzVW+5G47UZHT7jU6UmHzg3xdD8NqRZDkxXo3uGft/m
dWx7GrrAlsDK9Z6m3urO9Y3ZALCxFUddkp9Qf0duMdmGL7cakAdNqT8809xKbmWB3EY7KaaCatyu
gLNMl8xvAuIXpTBkra/CxHsMy5OlnfGhan06u5Cvb2MvDw4Sww1qjf09sBzIHBo9FB/LeUBYE30t
XPwcL8ysuAolfaQQUxZ1scz9o+lTspreisl6i02WnMPxc0/zIM30BX3B6F4mjWAseTSzIQO9lxWi
GgjUakZ+B9Yk17wGJGGK9mWe9gmoSfU21ljxA3ZuJbooGW7b0UDyuskjZsItXvr0B5iziytq4xdA
BXh4Jnvg9b+glTVtcZiq66tR3P8cfM3Bz32Ma7n72QOYC0BxUeYAxtd1ZFHjb9eIDUPGyMXmEgGf
L36acspVg8RmRiKV9r1Rf469vn8RyQB7dFH/iCjWEJEc18UhNrD+8HcUNXO8maqxKBzzxqRH5fnm
zLHE9vX8z0ZPUZ5js4GXz+PBVL+rLvZ2oN4TIGMsgkTL7uBn+/3XIEYJC76obhLtbk9+Mt7KL2Ir
EI6skom0hNSyVYYMtQR4mwAudeJh/fd/4Tp/e70HxevfZYXUl/BpOFDTCnKUxrkaCdSEggdT3lk+
LKADfA5/okm1DRYe9hzQcy2cea5/wpnkUlLdb8J7vqvrNi1d5XadoGFjFMlxz9DZr+G8sh+rCwcR
sRqtSBMdBhhc8bbwq4atieDHRWGgvcIHZME07sxLvjJymQNGsqeiC0pX1TQtDE7vctTgg4qoxJP/
tiKtVfUCqmcpAjzxvpsPcSDKC9WkVzvvaPRLe3fq0js9B1AR8P0DSuSQ7T3GbcDtmvAb+4oIxC3v
86iA8xv0ipnAk7p2TDOVJ363Ngv/+yexp9U9OrzyVsi3CC+PG+acNgWYmlNsGd4VUg7FsT5y4K2G
IMSgIN9XjHb5BNxgi153TEiyjj6ELGpsf+GMRTkKrw8+WdCB95R/k2qWAUZjIs5EsFYKDbnqbSS7
ibL85viWgt4mpBfECBPX2rNHAgr2z3JshWJJe/VhNVkxTpQ23YmL0nn1rNmmh9YIQwEeg3hCLncv
NAuavKRvurLN31I511PBcTWVnt5U9HMy4KEnQMdt5MP4xvCyh/ADchBwszShPhK7kNSeC3DVh7OP
62WVZZ5fuj95YcmeoMiu3rWsTQOra93etaWhLcpgBQda58Xw/CcunZm+s44yGBPKdofKAO+KkI4y
PjMt8HznfC7Y+xJ0p7PjrjDk8Gc3OLDyIjrDCOuYKi0v3HjDSWSjWxJ7l1AAkDlLDMUX9suQwuWU
r5pxmExi2H/KulFH/dqwjFxkPynGf6Dz49UPwJtyKUPliPV+2XM12tMkFRc4MsApRWHFyWSJJR6i
J9mL/1D8Knm4xElZXPIE3BKrlWwux0JZZxTA3KSG1KvVjccva9hmZnd+qfmB7VIeYVvDxR/BPlqE
aOvmTwu9iDUNRctmEdC42sNaDHkph5Ye0lBq5TUfZPSo4MHwBOc18fg/3eUjbnP9Pry6pR599Wir
iYFTkrMMLcL47nJoFferT3Zfov/xuBdZXdFiwIWJNTflbasU4YXe57sgmDi98TMyzIy6UBjWtySg
5ug3xl1prdNsSw9LY8I+0K78tvpbhqRrUmLeVWLnxej2bXAPW0/IsSo2+GzYiDcPvOMKdbrOZPwh
ia+kKlvt2YkP9XfNrpifdb0CK6A7ud8kyJgfbb0Jb4EwHGd96hAA2FFFL9pxnxy6k3eFz32eZpA3
MBVBNUcI13hdGFGafv+OD4AMfqe42dvS9m/Z2W8Bw8uK7PatQ6Jhcq3zSzVPWTR2BLUPimXIhJyo
aOs18fED00sec272ytJU8HAdJyeNtfjs29QYTZLM1v47qJRR9bvvJ10vKGyAWNJo0BewxqJstX2V
HrFj3TzSJYhoAA+TWbwllm3a6PK8NCPjDauADJf/TDMBEW77RHhu90VOO0AZWnFIiXlH3Jz4+f7x
m2eidFP2Y0194jT/iWZeomII/Umyja5LA/aTXIiffTyLmjosf61P2FbrurB2yFr3kjlbSDnWbvu+
CXTzJj6OUY+hTrPZHz4f34OkTYHSbUoNraWXMCpwGVrgkZnvqiWw6wELaAzpsmfTlVouZ67+A6L7
+ASQt0DF39hGR+Cl1fON0l6guudi0fT/5HzXnLTYudPIv9nKGnwdhun1UsXn+MroLAjArVNAeydE
EAS8QlKhMlgDLiQLCuVwNvYPKmBL6yci1+zIxmk9N1HGUjgOBXtVIVxjzPhdALx9eywkVs0nlgSI
ADMbu0FCuYaWQHiZTZ+YSYKL1wyVXfDo3UcrS/16MYcZuSZzcXlJTdLSmnyGzVl5fd5OquJLG0gl
FWjZsY6ob3zqQMk31qWMVM7WGCkfBQNZenWuX8yvwjcW4xs+JSlTxSaEmHuwvbEFKT6QVGicTMk9
Alr2GcPQaInDOFHJh1xqF+46GkNKV2LTo6TBrjjK3O2wnCyYEZWE+44mjqgMmcbktXPM4YpZJ8t+
jCiu2gdzzlsOSKZ1BboL0elQLUl4qgFP8WTShwRmBJL533Yx+DEXfJIaC7O/Qeu+66s1xmyUDaLZ
UwQbD6w9PRoy6MFEVku+WFU+JqGigyJZyFp8XN9ERU5q0PwVkZIiHW/5ZHHOEzKdYp5CYE5gEQWQ
OAb30VLN9mhscuaP0LIxJiyBzvhEC0GdoyvPTyWOpS+QAi+P3SIAZwz2rT8/TgTIg5ZBmIQq33q6
aX4ZiqPXNXdalpo6QpGDaasGl2RmKhmAyNhv7gDyoyz3CG/pt4vCrQV6MUxP1Y5/evJtYdIVfR31
XGPQPvKOWUysdQgU/YqVQOMiRPXeX9O5jSy7ZFtpAY6xalzQ4zkiRPYwp0LU0KhkuycnluSuII/a
JEdd4iX3HrP0FyYvTxKNbCpRs9oVJ5EVu3Qft2oOqOyFH6b3zOg2dHp8o7Ribkie1saTg6WzaQGN
Vpt22x/zKL6OanNH1nXnfIlI9uaHXyC3Jaf4vYhTWmt20pe+rvgLgrwKqDxuOwQyeqRTtWc3HXeF
pJdP7W3Dt1htaVm0fS3Gg4RQBUqoIFZ6vLf8ZRUulqtbo26N4LkmF/Bmo6Z5/74EU0BVMhDJ2UIr
j5JZsdUDoEJQNfDmxpp1qhbMGp7eXZa68Ueo//AtVk2NUv0cYJI7V5joNzSF+ObA+EfNtwwqxsZ1
u5FlCm6jV0e8uwzw6gcNffdqXIARyLDnPNaQZOfr9BlU3MxUXue7NrBdzzrzmbvZvsmy2/9cSHBn
FIciygt45An74FLzxnOLHvtAZfEBsABHR8Lj91ZrA7ZdDP5Mhg71UNuKDHIfspM71L4Jwfj5SBgA
CKYvVrQaBHKL7rUU4B8Va/eUnBSpTz4UeY020y0Ony+MUtm0UgjlwE9PcfI9cu8n14ePDruYZTQi
1KGP600jozlwwdBDNhk+KApohLtq8qzt8iJXoSfgkkw3tedKZYct9b0CVbmb8F7wcOGFG+lzSM2/
Kr/VrFZbGzFY5Su6QhrwRjJ3hAfump6QlyRAqCuon5FMxZnNtiJ8tyrW4JuuybdfbtYUsoltztDs
cOmV5Qsbl3QD4xUbJsKHi4HiCjCcvvdyqz0WXqfVUzEt9coGN8Nu44RK8PPBPKoY/gxV1Rj5+POv
nJeBRn9JNmkPY2rhSyomlvK8HRSSvNADPlU0MW19WWzA6jcqVFSivgm8YDH95pt1+4Lo8/ioJeR8
9absFdRSIloF4GijhjxAQBUBUqqKxn5jRu5qYFVVNQZc5MUEFzt2VNZdlyrFjhyeRHWsuAKZdMo2
DObmwPMb7Lj9cbFeELebRJCSoepCP4ave7MWWx4w/1RQLDE+u0zbq4GmpIBE0ZKY3H0NNdjKhC5k
JHWPl+lERX0jbNmuZGhu59CcBxOrc7dMAZh9MSAjfieh3rStnD1zfuX8hf0vWr29pSLrmy6C99s6
FTflf3R7Uu/vM0b1HCJBt6tmRV92EX7Q7B/iggWuD+HgYNVmDEl1qRhAfihk/iZNZtpQlMFyOAvC
DvXq9S/A5dJMySOFybTSngtzAskYZRwiFI913LcJkP/bcexYJxBAKpg74LRYFo3HTJNbuzZ/9+z2
ZUhzxRDk2g4RWpgJpxZ/ad3dhWP609naM/Zutiszs4zizWeXJDn4wzhh5peL6gIB71RGr+wmalsg
jafg8Wd6+9p84ZwV+Fl89Imz8ekKZXDQbdcn2+fQNnOUJVrDGkFImC3Ansx4kCt2sWiAGM68U2It
ZWRXId0uGLSR/1Ju+8ggXphebgbESrn0AAsV4FyJK6T+AiTReVJCjnOxE48Oz723v+vUwHIzBnHN
0FTdPiGlSEb7eNtbp52Ak1vFydiT0JJQVt8DILpE0Zg45YTrhnfynBF010ScElZb0jN39Ug8Pce6
9WPBNGFjCk2LXXwyC3RUkSWI0t8A5jyV/QBz4xmoaHdOfYyjjswn/B4SCcOmNWyr8JJH6vValTcG
k0BNimO+xQB5GoT+nNeamtxDQFZ0Zi/XCz1EZ0geNYGdXZgnCCjrViB7qRGAv5cm0AqnrG+AaCdV
bHjldBhPNn13fLPedwoKceb9xEomstQQUXxeztKFwHUa4OIHd2xPTetIddbzvf8sztviRZzrtntf
WaCykYvfeHe9WVWIWVX1mWSZfhNCnZCNbUU2THaLJKU86t1yGNtUNc9JEuaAsVdQ0+uUpkWh+UxP
nVQKZWEGjIbo1xmzF4lroA1Sc2RWl5jOn//fzfd+BDyeyVCVyCaw5qDggToAfVxk61JKeMdnTrqh
HGmNrtZdcE3qh+QiJDyNNbbc/TD+0XRd80QGhcuZPt/cAu/0vxmmvHU2Nuaxg8QHFPlP+GowSPw3
2ZKwyy7Ei+CBRW5TqyA2LcoIQrJg0xMyCAFcwyWo9/K5OU4Mem8u0lv7VlrThpbocXfYpnIe6A0Z
kpueXIoQfW9gkeShqb8f88l74Lo2yBD0jvAw6CltuozVtLXu+qOsM4SLWjOwNfh0Knz4YR78Z4mt
+n/3rDClKy1xLGYLJ+dBu8F4o1QSzgEUnOehLV6apFOFldun2zqRzCQOyi3cdgmaWFKzKy5F/iDC
O2PV6j/P1pNkk2f1VXem8oxSembS49QQprkhJCtmDN7qOU+E0jVbEDSCE16HW9pZ4nx+7Oqs1RRd
UWxMrfKr/cqsI/UMcWkQ1SLzgUmfrH6BPqgjlcSRKgIsvdVmxNdxWKzQkk+O+XjkCfP1G8jrXToo
pTFcmtxdqcAeaqMf1SgqMYsgjj3DCwguyJJJJpvRKEBApIHGyCYQTGvgOmgyrZ/KhERzSYqPSaLS
Fy4jXTEscZxyVMnNHjcKiI7aQqnmXiK/jH3+Tlh3CVF6TgGmLl3yNwSnRRuXwCdKqCpdnzWr1jza
SSBQrTfxtNxjU/dxnMFyGy0nv1gqHV/h+tF1BtlwRUH6lPcJ/mTNbD2LYto4xZkRgm4sYjFxT5Ln
xFc0n/h7GNFDvGcCs4GHP7f5NhZnNwpsBmAsG1CA2Utcau30uNm0woUmCbMtQlPcS60guEEbWyVr
AV47q05UkS9E79Bz2ACxBZJ8atg4G0CfGGrh4ga6EOMjuAf3cn5a9JiDZHhsZjoupCo8kVVgDxz5
05uDxJclf3k5+n3SB0WQwe54p44XizJQi6JNSU78xegB3kXjrKwc4t95p7pV5h3VeiekrIkNiQQm
siqb8zdjvwyo28nd/SLE1TKA2NIDkXDf4y+JoGau9GJMDbpRvS4vI6gcSFO47i0tcLjw6iC9OVbh
Q0ltY1rW0YxE/pT7fhUFYDTP7m2c62P4DX1RiMnMJSb/dfoU+52ntC0Zwmi6d/wmKFbf7hzXdx85
baY/6NQunRQbihsZ07f9aQmydG2lptrMxUVFqjLAnqXwd//uBbUz0w0sYwoOE7rgUAbWTAjnjerj
icz52aMOgKHHSMC7iFreZGFHn6qX9qfPSg3BBo3aDkZKU8WU3bHb/2p62GnThqcOF54OF3fIoD0U
6V0EUE+1NLf9Cc3PCJNwn0BbhvryCH+2vVXDrK2bCC79TslPR4aP2suiHJWEcbLt+QTpNDVtICVg
tP+twEGk7dipu4YLrnFNxFwJ1IZCp4FEGF95hozOOih/2h/cyKDuLrx+tH37NolItkl2PAG+aYnt
WY5EqY1JCkHZiJSCb+0Bx8iz8hEQXKn+HOn2SBBtXHb1QXILwWSgOlqWN4gDbn6FCs6VVq5uE+Pw
CjEQyAdFgZgI8ckuArvrR/4EuI+5hTcv+aCEQy6TBSlKPU6mPBUFy3lplN5HC8cBu/2fbGqNidp3
bYbhdFxuWLU9IGrOzLzofn6GBBHeoi8W+K4OBkbXbJLogdEb2VBuQDgZXEh18UH0YfyGYg3yZ+dN
DvVY16RKSdgbWvqAhHSg8BdAPF0nwUPWPcNQPpx6ecdq+GwrcCddhBHj9turXZyQtFHRvKxpfbYX
2PqNDTQgwmLrlM+T4VA2ChUUvXufHLXjkqo2lg0JwkDZGiA0mzpG57jSQdIFxbDZQT5Pi6vWXNx0
XvSMij28Tp2tYMiRinFNAkVcDr615cQWYgCGHh0p2NNXultd9yPhpvN5ntN923K5r8CUyrajFd7g
8u4Y496zLwJ058XobMmz3HmMWdW52R5T0vS0rWI1dr/sZLbT9tvgoHrAMcTYqOyw3ulzKlYJlEAb
BhGBP99x1WajrI4eiU/ec4I3L8tWiRq+nV0u5T8DzWHGUIsGAus3mtz6BkpybekuFgFohaq4ytn3
4aJdsCmvfxOi7BQibkvkIy1fo90epo21Md9QwciuL9jiePBGA7Uz2UrPCIJw7kVXigq+irUMjYxw
1BuGfSnW9QONJE1e0Ck5bZ8t18Q39TUg6DEuiZFfDE2/TdOmWZrIjQxiHK70RcknaevkzFnBO9oO
KAlRic+nXA6nwarJ64JCwojYznX8kbRKNCnXEhb0oAoXOYyj10aMhXOrX4iqHvetIbdeZ/KyM/ui
OrapYkII6KkdVBTypFV2j+JcRVmLolED0w+G/lZKwBUbIoyykSHjgCoY3pkihvCB4KdqhG/bPxlO
U88TOLrIuo44fcDoDdayBazow5q/xGrGeBdJt7+naz8y/PVeqUDxPQ5/YjqBsqRw0OWAAEaxEP4O
iQsNTIxwGO7MlL5Ctu+LbwmbjjLPjP12fu+iCci2/xnQUBDthR4+ZYhKV8kKKZXCIM2d2A8zoBK4
2fHF8gNuvxoGuT+r7BtxhEhgL3UM2uEvDM4CLBPvoKUdziTycMxWN9xBiOS+6HnRX3JfSfwMLT4M
CLWyt4KGhz0mVEzzDyhjWCjS365hfYirNwu3FCplA28HPxUwi7cfUYn6VBhl9mD86bd5unokE716
JH0KEnEmyDYQ7bQnX+ESSEhYQYeb9ZqwMbngScBD1jND35RlfjgM71hyvsmv2vXjldETBPzoGglJ
6GeI6t2YNrhJPnRLNs5Goa5aWgYMALg7GjYz0xwo9rHATZj0Jrlcw3Y4SHv1P37AfrhKg1jRXzN6
bioSau5q9gz1JFyCrJOkJCH139XVdQkp8hpZAUkjFYnDOSOjLqFyLB2f9/K577JBj1U2DLNGUldv
ppaV1eeS73W828OS5xg2+X6HIgUYjBYSPLZHqu06oWpcmLfwGNkdhTrZ06A06UqFbEIBly3FPIVN
EVvqW/iXXwoeox9sSQWTvte4vcN4qdN1g9A2nd64IbaK4Z1tQoBtz/sNp2pDBmALaQ3MtOGO6+4A
OQ8VVfg3O9KAppjfF9giP7IQwZ07ze0TtrzchV7XeA7V5MIuSoMOjuykEVLdBQrw+MYx8wWCGKRV
CxQdpT8JghHcsxO18vuZKeMJt058tgpz6JpTWEsHvtczKURarNddMicCDMWtqcPvC4vlpfa0gnZv
DxcqloV9q7rQJBbWUltRSi7DyTnQIWqnam4j7mct4WMMJg9I1gSMujy0PAX9kgCCwg0qKgAxHjtc
MuE3pCq4ScdnD4Xp3Mda8KAQ9VkbzMKBxCyfSzFJIeMQdjFfmokjFlHQm3mwFqj8ezc6aORQo0gA
NJjKX0RnQZGGbyJ1ZIbzlza1Iqll1Cz+OXOi0/PYphAkXlkMYDeOHAxWG22qmuPODp8usLwJfT7k
9t8GL0oQ8BVUsFtobDknHARJAK/KbZ9OcxMVwj0rzucuiGab2iJR2BmmqG9yYzQC9bFKKzRPXpxz
Z4RpD6SS+VJ8K2mnihLWiIFmq4h4arBeao7OjLZ3yeNefyS7vUHWwSNeX6ud3pX4T6//WoLssWWY
2g639BStHkZ4hNyFpn8+UOmNi09hIWcWUsJnoCEPcmTP8oe4JX/8p55WajL4UQwcjq2WXRZpN5jN
qL4WiIr/0JbcFuzco9KlLzlvh2NxtniQmzni9gALbcnJ3Pwc6kYMxl15t97GeXimiCwxP1j3oMJV
WYCR8sR52AFUylQUrrbk9hMVHJB8JZepJGEqUdjArtokGhfiqSHujPcOsN/wvlCfYPwR8QmEWyGM
/UrMXJJ9bSUSVjsNDuIMkcCqBCombdnDPoREDavbxT0cPOAyPSX5FuUX9BypEVlPOX23rN5jw/Zz
xHtm387qNIYklOT8n/J7jRvXivFDOsce2ALLqEl52IXTxoTJbc/M5kXcclk9WgavAQbLKcGeMlyD
m/7n0pAZQNOzl/54F9teVTGzW9S1DPhuE7RroKC6xOVlJYOGX/IPWERoqzyX5NmGE5FkAQAm88wB
mZwVEFlvCowPDSHDTelZM7s1v4LTZ7wncW5gYjK8ZMDiJFuJABNTF5T0cMqMJRq6fsyOFeLW/2kr
ijK8tZCU0WhZxX2RmFLSvYo3ZkHyfDhO8ZzAldOa2Wrr/bHczhVer2b5/xns/P/BuvgQ14t7gMdm
vPrXY6yXhE0Yv8yRabv7bpDjbqLTRDn0Hne5yVzeU10wxBRu57WfUrnbvmB49bP8NpXK6UpMTNqE
QBIwCsuZECiNC9xKrkjHlKpFuKi0PNnvHiNQ0xYtxe32pErzm/cnb4FYLo8LZMY7Us/gTstDdZA4
6QcBBozpzhac0quP/67BB9B2B6yfazGaqPeseazDOOgY59ps+6iLFuYRA0B0OmDmZWhGJdcjHfLp
sFk2dESCGSIeZ2EOQNDvpzTN+fyUFrz6e883XWfi5JPemHEyFEGTF6DMzh8CGupJPYBCK7ckDuPN
yU5SYyn4yS8wXPN4d8omnDt3ndc+0p30u4RarTwOcdJ1k6CtOicy6zEV6VbjN7y4LMekEqi4Ptp0
YvJFssCvQZejK62nEcMZ1TyQwNZmgBoqN8tOdFA4dQpWmCX4C7Urd2xJIhf188a92MIGO6T/ofc7
r/lwY1ljOm/WDsnTRn1w5UpaXI3hqkeqpKNiKBJ+8kxkq/vdHXaP30Dhr/d0BngkuOzKmn5e80On
Iy/QGipn3wMZL0tlMpXm67w9OOHVK5jZS+YNEmwoxKFHRi7uUSAS9WgM+aVyLGhWfzzcIdPzYAlv
U/GxXscFy+HjxoURNKSBDYVxUHb6KGmnkkfxck8YQiaR5DCgOmsxXxgrB1me2Mym6wVw8q2LXxn/
ODecpB5NNJxBdHL4RwgFS1ARcGyeVJ1iOLXrx/OCB8442PCia4Zf8JIUzxqrapO3dMpLvgemfotN
jzNSjQzgGDZTxMMrTVt2QiFC0kkvsv5CtEjkpSXpkAPex9QF4zmuheQMxrr2unCUm6TyzFoK2/mM
fNw4l1lHGF8QIR6nF2XDkCBn0OdjVrFrk2FSPBDo2zwCwO0dQsd1fK97fjF8k9cAs3G3LdSZZcnB
qiEdiZufY8p3vFNJPcHoszAItd7jp9/Ri13ZrrtO74gmCbs66mb2X+WVMlNfmUa8cYphs1+vt71u
HIQxtpYS7ToXZhYunIgPBv6DW6L3xfkmIz1FH3AImi3/VysVwXDmB3pXw+6HTJmN43jBL7ru/r53
YE+LDV7tb2xlLkzCZDodc73WV58dH5wIkAkoqHNBc5Lft/vVrIg1BT3+aeQO929whfpRztCqF1Ik
H/K/yfb58eeheI75bgYQwrWnDYvdIIFWd12jME25FYcyCkPLhK/V348SwEGrzZnDug7FuyLECHVK
uQ+MD39fRAIYUozexB7DOTlQy5ilQ486pIIP6N56DjN01xWSd+5Xuxh8YqgBtwgXV6SqNML0+DCb
1niIVQQPxQQPLyA6/rJ4fqXAY7MMTnwPf8ixCw9CGzc4ZglSTftQufqTKIqJ4PaCVLYgTVGDAkYW
Vmv6BWi4Zm0pyu9fZhNoobPyVZNax9fg6DTo3Jbh/PGA0PejLhZS/MukKjx7Cr9lFZGL8XeRDcmH
yNshm3uByFhls/zFZC0Q4NrlcUxkdw21kbQMJIRNlrE999P/zSQN53sUVBG0L/vufboQzqzzDwfr
pLiXU8ow3l3JwjHqR0rdJD67S6On3tMApJcMNG9K+JKjYUdKgYa6Om4k8jwMCdpRf4AhKolGRZtM
pXMUXecNSF5ij0IjdM1NncZNVz+h7bwXp7pAfkJyqk2dAoMkV9dWa3bUN6HfiA6UViW++f9O9N8V
iUHccBiwvrR7rRHaTqB1Mg0oiMrl8JQX/aRwvJPyRmpfNv4N04aoVa5wHAwIeNK78sw6P7WFphWF
fU0o4e7Hhj+kVzP0dVdVuiY3qTrkXT11uU0BTXVOiQIDrKuIe/gDEFFI1UAmnTiUQFyLx2vnID2O
tbKt91/eYhNPhKhOm7IdL8Rz6TCNiHyFx0S5TKEIuaNLm+Joxrl9aOlliElMwwhTcDK8ShEui5kk
bVRKAY0GuYQ9SBssQT7FTQjyJMmLy/imZaeuLhwnSrcNRkcxTWpA4UUzMViZtAvArJBo3gPtu09X
U46MTWO+rI8JuoYC7+ussucaUU8ot8HKGKtN/cJ45w3fgGVvyXdGvyFDm0MbXPuXbtfMgGrbbMnr
2a/EeaOLlgSVqYAcE+N9WpUcgR620xLMisHPn6nqCEne/uhGk4GBtUUo2s9z673neVSQill/u4ly
pF1bOdJuEApRrGEl+XBNb+3dGb4gYrhTwGEBZpu0MdE3URUjTIT99BI+sak75GbhcfA5FhBv/M7g
19njivRs4X3r3asYZBBGyYbzf5elCv9rpyBep7SEQATR7IwIsP4fmY5imDwzjaO2cLvwTBnna2QS
o4aPKGH59sziehI10MO0ArF1KIPN8JGpPUKJ5dVXieWZcxz6Ifct7/EwsQtcsDQGHhMLlBpkzg+o
UvO+41ydjsIcSgSediJoysiU+JN/XPjfJ0VK6pyHzuEed6d4AuXa8Prq5ZbXccwcvDF50YdJpe4p
Vk4tgbAaIFeM0IV8/zzsXX7Zy0efz2I8MZoEjUTMaNCihq/0OVuebJtclyy0+XfgpNby1c0OM1jj
MqJQSdxfYbWVKQYJLy/w9Ldi4+379yPxgiBxnZRFHVs1/03vQrd58SZk/EcHc3uZAHjHpor6VNJN
8YnZhgpxIu01GwGV034nBTZCOlLmMRC7S4x+1Du1X3ARXhBJnQKd7LTqZOzs+LWI57R96rdC6exq
Gw8/E8IupC/VthHcI70ExI69/d9tO2Ch7cEoAQGPy3kgh/BcwQB00w3eaKdRcSaf1yLgGK1BgH01
+3VSfRYPlrgISRk+I05kjlCoXzcK+7V1kh3VV4GWAHup8xGiQNJq9j14JgzJQjLtVqN54ULcIyC2
sMY/pE9w0ACv/4F+3VnRPOCz2crT6sIVj1YJRWe6t649UJ3Kha30e6aT2aCctJkopeC84JfW6TWB
hDBXqKl5aEh16mudyX2UUUc+viucJAnkMQrGeQE+FhKDI+bbnwMR8jxEFQ7ebUh3ap0uSY+NA7Ui
6E6znFjMUIsDf+GKd7t7/1EkOYEi04jfSgib2g8dC/J8+/10+37zj2enEs4RCZDGQRhYpxDMMbde
VimOk9j6T4mkTP8kPhoJN7aE/2Jnt5p55MYkD2YC2OP+v7wP598AOLHutojQoNJUqaAABO+pO6qE
hZh+tuit5uayqSDTOfl9BJ6ufOvBo5++sQ4Msl/OAcaDWd/+GdXMzqqglrSMt5fOKyRnZeBk9tAQ
5Q0SqaqeNlXm3sjgzGM7LRIWHOGPr8IEWvGdGv0+7Ze27obZ0UkSmUd6XBjeaMcYdIicpSMOuWj2
9lwQ2iD4RF5FCOEAbHqLYIPkmucLGGEpj9O03BmzXo6h6gI/WhxEcfHacp2SybFADLSWEsven/1r
GIe2j/G3L8KtR/TAnCoAK4P1CDpC51R+8LAlewXyxZZiC1g6l4QTpdgB8MvN2TPb9XkAJidZ2fPo
zxBao0W7gz9ut2CJaeCQbge7YeUj9LXdCedkzCVmS0MuJF7Jir0MBMamPfPjU31Df0EsEgyT8mVP
hlEEF7VQVjjW0Ux95n3c/dVnx3Zuw32+OuxsyDn0xKYBr2Undn1W42vWZcnMtmafzYu5A2Uh2O4y
GO6XQsiXI7mgHE6s8pTCD82V+Q0qsvrMSokO5Ai/olSzk+dH4GTrIMvkqtPkMhH30JHFZM6nrFxf
jhC2KuZBemY9FF9H8M3sJm+7GBhJxRBrpY8JrdsV6OL/GOIZ9EdEeHDMbOdcgZ4v2YU989TWyXO3
Ct5c8//wygXocHvwuVbHcdQdrqOMyMsvVsmUoCIUqNrfiKuIeIfALr70M2VgW61xdyttKVZA7pGM
boIoe90xnOKrppEUzdyJwT6Ju1fLgubFfuozjdUo1+G4/K4nrXPxw3JCEQOOkCfvA3jID4B0//qc
1GkMrCIbtqok3hfd3FyU6yP1+VOahkygJwBGKQyw1t9ArGylOeH+My9lj039gBubmNrL9v3Q6ZBC
byo3btgyVh+ErNGLvzBUUJ+u7/WRm6t+uqqV1ZFAVn9eDw3W/gexlu6s8s0piZHcnTgCU5mqN3fo
HRODpd8MOW9VHI8vPDyUOXadQlchxB+x/e/DSN57e00FbmMhmdViHLF/B1WHywpCq3QVsdNaHXrh
U3sy/HUgivKDiuNxPACYiwKrPqDWGhEodftGhCYr/J5omoeJZWl6dV6lTukp7jfmU8Q4nlJTZqWY
9UebxGn1wvpAzFUUXozX2OMHqN+cpkrZ1JwETTYQNBWmjoFQ+7sC/J+L13NlHS/ru9oIt0LGpsi+
hJgXcoy1wc5tqF9k+NVnIXCmkANLM4bXJDoYFvLXVubPfj14+OxYD2gOR7kmtW1hSugswiRYhYV3
R4zYjeZHU/RRXNNI8455kSqVmxWNDMsvD7sLC8giwo8s2hcxfWJxrYgXVY0wSSzw5Jt+r1N8t2ZH
i5uphAoK+CZRUC8Le/mH87QIIRGKQw/NoN5qZXCCIWID0BuVsMxJ4qZyH13Ki5j7xE7M5f2Of6ZG
XVvD4AbOdj/hkOcRZr0r+hWsElfzW3cmTDkXs21emS0qt2yukjrAMMSGRQ7tjD7q2z491KwUjqC8
SbcpsRCrYXNSdnvzlH+leGBYbn6kAKzKEen6tNzAe/hvsMUTfHiA5McrbSL6sED7dLgpg6glKqfr
pja2OKm+9fz5OjyJXUP4S/LJQsUpO/YIs2dJFM1iLgan9VMlMKXaSP/6wAuGcPrV0OZBiek1CX8Z
eiNQQgKNudoKIGdqCphRaT//4iVPvq6LTXzmugJUjVUb7P+DxuES5fStIXqi8h58oMWHhJOsbAwo
ihGXDcALAZcqOht2tozYs5dPjPfrB0AF09Z7oE3ZBRvp9RdWQZnXXzWdXweHjXltSpAvjmthLTYM
WDshyTG/Q1RFO1E/5LZNu0S0qwYDV/4wMEH9Ojt4q13RhEE86QnxJ93t05zd8V1+L9UyvycRi3Sm
E2yd3DJbjyTBPdNASgWyET9MOM3Re8/z4ouNgVTpSfIMJlAtKgunCIdJnXKmzHHrR/7fvU2qq6zq
DoTyvW32MisDDzek73b7ABDQdWs3EdhpbjDrvpZR/uMiP4/MoKRVLSYByW0mPvViop84bXOq4/3w
y09o529YMqEdjs/O2kZiWaUApcq3rL1t9x69YULy5oftrYA4i9/VLGDEpG2oqkxgBx3IXEtclznI
rflY6CzWclP9PRP8NM4sK8G95gxMaiLIcrtPicm6nLwF7sDUWesDosmcgJ7e7q1hT9HSbO916NlC
UdrTSjv4NhZl7RNxUn+DPg41o4Jd4KvK+KjN3rkv6qwYhT13E/XzMs4BuO/XnfngVvvPpIf+T0xd
9AvDpGbirMsIOkyPmCQw+LbCZI5hqyEH1eaadwQaqo8W6XZ8+lL2e+hnx0LYHiAUfhTWR5v7hrL0
hx5eLQbdBjomh2A05n+9Lm5fNk1aZcFomRMVMIsIjLbTkfucOSVvGpoCYmCy9heMmXEaIxnxOAeP
ltI0S2eimhxij9Gte3Ys6JVqxQhjHZoI1W4/W7kIyPFBB5zb2KB0bS15uP+RSjWwa0kLy5Izc9mh
ec7IOm23xDBUFHCUPjqPqToTxP04g9QrvrXI4TP0HVa9vgIZ2mIxY+31rQTvAt0BRFPR7A4ec087
ooMcDnNH//J9xbrDqewp67DZUbCiZE+uJnj3HabCgbHzQdS2xD5X/RG0Ysv8ICaS2fXLOGaOepbv
U8YegL79+9Q60A9Z727sQ7VlJybE4tv+zTUthXLvkG6NfBvEn+b23zOZ4u/mhaYf1Z+QS6czMJvy
V2LAUhvyTQsCPDPSy4jCwPCi/6MOl/L6AuayJ0WOJU9kgead6J7URfC1W2T0dZotdYH482MW5Yb/
IeXYmAkVtmJ3cWo7T7TwLG4q748z9q4LVmA/nPs4H0C+CoYs06rq42o665ewMOuQhjy3obBD9zLu
et//AhPoCErdMijt20XdV5OtjVOnBu6hNhasN482bO6itPXwLndMOaUe0FiUeQgInsO332T8VYl+
Q062wygzl4dFBMCZs9h2DB1w1p56rNfFzA5ZnfS+mt0Y1/uIGHLHPkhKS3uS/bl0YFJ7a714/+0K
E9KFTC2OMvTQVR7/hfRu4dfyslusOI7jxcZyRQQ8iXFEK/ZNV98qDfvWaM9ineSwQG9ltyueWuA6
GqHOYNr4Oz6RIBWwB4SWYP3xZX6mtrAW4AU7u5uAKwqSru6tYX9aQ11LBNUNfVJI9sn20vifNBQp
f1awa3SN7IzEPeRRzd4FRzo6kyQZ2lCd0CG6c+upm5z19Qa0JD0e3ACyyVI3Azm+dKcvB1W/umP2
8EJSTaFdvO51A5cy04uRDzuHlivFybaSabLBCFEiKrKagJ/UPvT5K0/bWkO+xwLkF9yNTCnlMPcY
JSMyLmERhHHGG9LhpqOzeKmrdNxd8fFlkoUQzfp+HAAm1UIYplR4VxgPqu6wEbnWpWOGmGyl2eJe
kh5uzwfhUol7ikk+yWUfS8CluhLXJ3TDQGfyo766PqijHICTNvVPQcvpASBXnIe3PKscYrXEDwNF
N5cv7MmzDo8RvdGm68ThNSUZ4MNta6EsdcqgeFdrWTVEKMtuXyYMoetlKSydYm0W8J0eTT6HuBsB
NtlFWlzTtvR/yXYrxqyuGEj6ages+611+b4LedzZiQZD2Z6p4I434pJJW4v2vb38RIWHTZxOynyw
IHmpCDnidJCDYAFsKjMGFBhWWfvR157cImfVryWLQf/r6NXKRBaax8RPlLOzqS3PBxXR6awTU1Sq
5dqkEWKBVSkJcUCsa7UFgESOH4uMj/IxYO10DPdEmWtSIS2L7Rzbzu95jlpF97uZAEg4BPru09aY
sRY7RMmwXe/eYAkbOMqe3MNZdnBgRMWccOugTxFAebVgLWZjseSaA5O3/TPljpzVEONCunCkcKib
xihc4e1hDSRcH2VWDDB2QcGkC9HCxMFdigJ5BUk6vmuBuDyRUasvlfjXpxnywOnwifJRWUb1JKGJ
Sul1xIQN+Dj2iGSuj8Sx4UjbQH0Yl5TchnHHe77A16yAVqZwcsrsu9W1WsEgRFJx0syxg8WPGaBU
9IKHQvpf45PqSrUSqZZek2qvODZvKrVacksAMz+AXHjRFVVnoweof2Z6662Xmaq9dcm+zvAW9rPA
RXSQzzxNG9upmwBP2efBiV9byavAFzf+wgxBeKpebtZp/iqBHwLWzgXiXxG7LO/VlQV9yN+pSTGM
+KPDAYE4f7ZlLIzMim6pgg9sqgXUK5/DZ1cwzi5UwV1erWYlVsR8G65hD7Lgj0t9OvA2+auEsZXv
PamYmhJUllD/SoHL3UN/cUe1xcJyR39NAFFFBIZUUCreLvIrxSI7Jz+N5L4bVminvJANDxkDSlCR
3d/B/0pnshNTg3lDJH8hU3nXHOc3e/kvM3yVWdnUkRV/63HZAxoB8/KDYduY4heQ1bfsXKKNcPYw
ZDAaJRqM7Kck9eSapLVgbPDZtEJpluJ2Znr/tDYTQraTQaX+EprcLfrcnT6UOqw6p5h46otry1yE
uqofmAwJazVHGuIEOIVp6LMpAYq8Wb8ovwcpVXcmWOCGS6ynwcWknaLcN9yBpLmj9+iQITYKIEX9
8+FvweWHYs6oI91NRI1JLZ5cYkE0d2ZkF4OwtKOiV1Fzkn5ZvoeX3S+XQi/XDp3clNE9BIqXVcLI
EmVFpo6Oynpmvx/N1P3jK+ZG7r9812h20v14nClHc9DNhTOHAsQkIr0R6dGve29tPNFIaVVyF2iZ
J3JOSFHPUFCbRapEys9sbFk6tCOb0CpZcSNdcclBTg/LZ3Tn3zdfhm4av4qfxhfmRzABNWDq9mzw
dInybcgqM0OvyDHSxeRfZL6InbaTM8Gi5zQBvb7DWrF6enegNdtMOSFX9DO4S9oaj1ivBYjknQ2h
RpLzi4fBoV/inxQOPaAqc8Pl3WYQSy07jXScR+nimZdletvV42yefEkWBusRsLx4bc8Ni3EAc20l
9yQ9TxV1cH8/6MZ1p+cPOMtbaIDsN1Sleg9QMEsFzHrjhaSlxAj8BaGqUBWYOJM/vkr230ODPayg
L/fYkyphmujPkNlX1YhCkp3o/HXenMSO70kGbxoAK15YstIT2t5RQX2hp0JCxnMPVYN9QVD6g272
k0p/Y4T9qopaTdRl61UQIvWWTb7c9FELjBI3cVGarZKOgx34vGP6rJZgnax5emQhxCuXwe4oL55D
sJt/8U7hUqk+bjsBhAgJtBKOZ92cs6wy++Xn2eG+1UAE7ELzC+wFP5Q8W83W7ZrujgrMc614WC0n
+HLSZeTm2UxvmqvIi6fQ3JzDQTJEq+LQC0G82zr2Q9p1Qksl1xTByqrd0A+Tb+hJJIUsOCq1IGzp
vAkKzaIt/6lumsb7G7EMvICJCa8zcOoao48NOpC/t7i5ZbNOSQnR0QjaVqnfKWdWtfAI5XZzVW7C
CXghDJtWqdueWx+7L0/rZWNsiSRJb8plui1Lj0HKiYldyYHKcsR6e5qi3elUBGo5gq7PqoOhV+B/
4V+2XYIZ2OaOlXl5NFaiWr7qMwoSphRooe0czggdYx9Td9d7SlzvrFGRBKwW90zi0xO4czgS/py0
vLgXfEmRSKaMKia5crV/J5ExniL/CVAkIEWjAaZYbZIlx9Pe3/SJkMLjQjpNCTv7XTwpzXyONOvW
+4Z/iI+q5PdjFKO5e7UiQC9x+ug9e2+KYnfT7xwr9iZSOyJLg85YdDBdZJhc4OGwF5kR1MrPwBUe
RA7xAL2byPAS+YyIbzPHrpRaDEGpaJfdqW5Jh7TW1q7SAFZLx2xXLQD3iLyMzT1McQGvAhjwPZy1
dAcAuVJBxdkpYdctJIHqEgRPlWYTH+uwUFyEfbxjnxs2XmzaZzEHLozsfLFTqXdTGZm3rqVPspMI
7t2tBZlRST2UO3GINWq5fTaJnsh77P9UUoqct3fmYEAaheINWBnFt8Y/oGKnAFr/2DCHSThl/J28
aqEOCdiGPhqQ069JVHNXKufF4N8molGGFYoNwdxTQsIt0Z/55qm2eiEIh7aP1nUOtLehRKkVWBwM
f9V+CvocxLqHDBfCCzuSf3D/H0mPIKeGxr82aoBDLeZGIcPijlqpj9w/ZdPMy2rlXnEZpEX4hZ61
NVhw1KHK/9BsNAhvU2THWS9YQczmAtCvG//AWvhWlKMufzMeoypBy0tt87BUnhgYgAmMCbyuS507
h6bxxqnrguplbNR6/4pfBrc9RV6tNCFCxEepE3Aiitoop5bzDSy68BDsFsW07RGcZZZc8RL7Kcyl
ZXpYT1YChg9qBWIT0BfzNucQYhy3H2uuWRlOTPBQh7d2GUXjilT1iipZWm2WnoWzXc8yfsCC+Hv5
4rxqWhUG3oP9D8YDAFUoxhGNEDkTeATE8HIw7cdIL5C1oZyDddwW7DLp1m+jvtQU+LADz4hGXmOm
JB6KrFVQH7Uo+Fz5F9X5savWYFdnPkI8fneLgEMVYad6a2a8vfDNfzToBwYVwFfsEubwh6emzKUj
YNTTTkhuofsrXWq2Odt2XhkShRhT9GaBJ+x7UOl3/xxIPF770nbkBpXOO1uMKwi5v2RMZ3HdtqP/
DkspbpsdOE842KGYb9v9dNZ5i25ggKkLwb8WNnejc5yzc510+VisNHCQABxE84LXxmBxGVG0dgjt
1kZPWrIze7VESMt3gjEZ+nPrBPTRhGVs4OGVPPB+rwgGaB53zinbT9ohQEGTc25ldGFuFj0P39Wz
MF1KwPQuJyIM90AaFZ1cWcSY+ubvQRAt9cYJGTPmFYGiwfhMVxQQ9Dqpul9SvX7NE4Kd7ZqVp/ju
YTfPHG5n0I9xkh4R1caA0x0y9k0VIaMxoYtNnQRLJZ9J8zf/eVS2mxD95l3KQcHwDKDNZHQ9X1oH
XlyfhfXYkPai3pZfE1R0TJmc8DuFvSV8oDZ9o3PfKvEhNC/DLMiqR0mKhoZimTudZEXxCjY1dssN
UxccWoTHP05wcvpMt0b4vk/Zns+ICo1ubyZlOeTMZgeU2dTuJ87SIhA74ngKLQjYys7otyMjuiVZ
he/K0sRABHuQYntAQhCXLLlqo8juD7BvD510eaa/EvkhgdjD2lR6IIW6VVJZ1diRYBWYu78wCv7Z
2oYIhpkCbWwuJSgH4zsB+cB3AqRtgjDwyPau5G9phcHS2T1aZsBhgjAipiFVApyrBoITb8zU7lgs
VV9NL++vahm5yKL44wsu4b5WoqyFKfCfICKjXCtpJW5pLBUr0o4pIzEXYQkRevA4YBCEwP1qXuKg
e7C2EJH1fR8hZrluxUJE5FMOL/9yzP+YlREembqSpeL8cgzIqFUIusX1DXZGgdsfj3K9Lr3ALei4
4MWTMLKN6NA/b2S1taVOH982Jq75gMqJvAVsD6JoSq3/rIQUw+6qA71wt6oUKd+M8g9wa5Vv6TdM
gEaRX+3E9EaPAwwa/WQ5poKTjMQOFRg1O0NsCKjWAKB71nEpJO4Jj6JYVFLdXgbZw/Pq/HyZM5ib
+VUiKxIfJFbjfgXN6wIw46BfA8nv/RVTOWp3zJJkux4Hi0NKm6Cm7Gv/S3v1Z2XiztZPU8AkBXmg
FCk0wV94D39jPr8KqPG7FOJ7KNhNOMv15ECU2LSGiT6WWQN+WZIwdHwlZAE9tEhbRBTH436uA53m
JVoGD1GSQN5niVGNUP6U9W78f28Td/jk3951bXZbHgpjqdBVNeXDOHu8XLcGFF4v4YGb2RRskW9X
1RN9Npoxqu5HQUu8IWuLScZ67cXvxYmOyYZU7VdhHAVJsqf7ndb8FeiSVCHLJmvuI+l9A7RyNl5L
grEYNOALjAcKu/uSnOlgduIziwcZtmO/6QtcoNveorYLh0pW4874CxxAJycsO09BwZCB/AJtKmjD
Hg5Nbag8hFOxvbQIFcNr5GKMGk1y2+CTmFgCJ9wGTu2dHMwDBh77F0MvldC+a3wZV9V/GBgeYEk7
r4wFbSp2ildI/8Y6gw/5+7fede6AdIl/TrX/HJ37q9vkWjTJIXwON3vjNsEdVu1RhGQj1SWwYwpX
m8mb5FEEDBA08Lt9VN3BES0GE2Ot1H0MsedEAAcJWfpYvStLgGGN73q/Ee4qvBeZp1A6CJStO0HV
4BNiP6t3iVp1kjYIRu6MBH833oYe6R6lFVO1tXAsmyTp6SEk340wqhpTVigz6rXMFYJyTjIYOq5S
3yf3kolrcM84IiAJp9Z9taOKxvPk9sRGqxM/AOPF/CuPRipd/dXtJe9V069wbI0kdmfNt2TQrUXq
XWpYQqAIJfMTC0273M+YCBkaDFerEa7vLfL1yBvT1e+0K3CWZKJv9qWNsFxD7uPs8VdVUDPfVlew
0EmahBhcJsromm1ir7dlel/X5xHJp/z2qPIeZrHVCHoXRGAO1c4BCpODEqHXe4S3qgEBJYur/XtI
gL8gjyRpGSTBvKhibTYLKNyKs2Z2egz0VndfqHsJ0DND+zTFKSYI/jTRM0mPk/2g4HdpNLAZ1ozI
q86xZu9BKSj53qKqlLWVvkgORafur9i7HG5vcbI7S+2yUzUfbbqWv2teAUCpBKkzY9jWwTzMtsNa
etl3G82CrypjmyqEaYlcn37Uasmxy+ghFNN/h3IV46sjKEdwGFatWXClboJezgihlqYQklVZuYYH
+R18J8tiYc1KLOVSvlpDfmtAMI+wceiKCiOKZk0tBbrw9LC38Mm561GIzxBXtLGJUV2Dqidn1d7E
v3t5s2/q+Uz8EdBCThF2V8jousy0tEZ22N0GqZ26Cbq0oBtPIB4f9nf+yj2dnuGMOxIPlutMR3n5
PzI+mdsa1/Ptrr/gDecuM0eUKBV6fQ2vD/EAY831lUfoKAEnq2vvIfjXKRJp8wWYNNoOncC3Y284
BcFn6mfuXtKCN5P+HsnJkEYRSWZbY//AKaTuUBv3pYqKAxldRgF9ze3+fmgkX4xvfEd+vZVydziP
0RPVW6bV+dlWFoDRW2J15cJ1Qbk9g+YzoMxcL5E7ufFytC5IvENIHwt8TQvgv8A9ptQZ75YmVJQF
PE8aoJXaKDde63pX85cRQNqHZgSCr4xqowB5DOMAdNOaR6CiEBY3haBZVX/fMaU9IyJbc+rUQnhA
OXg7qg2KpaOA29gtln5+jTQQHOzapaNzHe6mEw68As8LfUkPdsHAJN652w+M8Lmi3x2MbXY8OYb+
6bmEOMHDbfnSjhJN/t5VO15xgiK1e9J/zQgTh/Q29Nvb3APT9VyzrM75XUzrI+4ZJlL9392IL32o
pBxu+w5QH6qa7qUOLkazrebbl0TSrp5T4HGoD3seyf3XdwgcEox++qqI0rXsOVQrgr9JIHIG2M22
lC0cJJygVq6EgO4Nj4m4rtiVi9jQCijPKPt1VT34k7FKkGWV679UfNduTFbAeAA8439ZsDqHbwTI
pGi5/7uEUIiPc9PtqB2gymdapBMnD0w1GbeVfogDzdXxckr74UE5Vpfrr03rTv9+EKEyn6OgLA+P
4ULwtU4cX8fSU5wROvUu5MySqLTjhl0mYPEkP1eYeRgV464AdMh8KmZ7Xe3ge2UXfFEETIOn2SmP
/98WwblRx8uEXp+2cfV7MDibZRf0bBaGwdlriUaxNjwfX2nZUPiK4jMenk4Tw43MyDdI6OvIYB5r
9MS4fhsUNaKpIH+M3/xIp+jnmtY0vR84wniZ1JdQuebDcc78iv0EJGBxgXodvWSUEo0AxOr37yJS
/SK2Grz1SSU0wgoI3cqgEcBoLNt6kcKtpuiy11KZsuX7hYKC/J538b1lmmW3LlBEl+lkTVErp50w
kxIzSADTITWCeL19eVFkQCn/cf5Yfi30+thmpIx6VYArDhRfL6Rj56ZyuIj9WJQAbi4zwTMRM51y
0ad3Wmu5VG3QBzfzVhfHcpRd8IGkPuX6D2CkkI4k/YAEYYVhDukF1jYWceHA6a089tQaK+vaEeYI
vtNcCr4z8P+sKqScnlivjSRh93sfIEzRwnXg68T7rkhQONHgqzWzageY/WnjqYwTmRrnA0XXJJ2Q
Tqnqs3jkI2dO2b2SEE5Tdh4iSPkztGKd4QHiVI/sI13Y8UsbFgOwEVAtHz/RBRAVspi5Tk4c3Evu
RT88ylC21Zajzh2Clb9q1Lj5zyV7CpgF7XAuRnrv7kAgWVc595AFdXvvh/uLvGrYTzNvZB6D7+B8
5SRoW0g1nbUPV/tUoRoDP8QZTX3v0uxVx3kCuLHvK5VGpoCpVJVtQRz5+topXgA/tN2RcGEKwSeZ
RUExig3PohA/PTCWyoR1AScxmhlUllLrme9lxd6PibYmZCt4qy3Ht9t3qizJ1dlOkpAhWTdwJ4s+
LWkONKcMaz3geen2vnk3lBDuSH/zNUzrBl9c6BxSMtQEbtplavtM6Iqa+gyGa5NEmipoy5SKjK8w
PoRy0tH3lsMBlTT0E4WhSyxpfCopd9KaRMVJOQJWeVCH2CBihZHgTneMVDcEanAhILYETkH49q3b
fxpqSr8YGC1tXPNsnZ9QjOB37uHSJBGBS+c9HuRF1fm1laSircQNw1nX4a1ONMaX/wQAU+zv7tlR
/XjonMFfdiftptlPfU6+blIj/ewbHpcD0XLBa9TEycg7Abs/tV6DfaU1hDSuEigSbdHIACPVTwcT
wk2K1Pue5KzVznMVzGaHr28+qU8CNdok+GahhTMSHcqm5eK6wqcLGuuoxmj3R06tYTmm2lwGqOLp
GeFKLZaxCLu5hkJIt2STYqhMsDYfnC7Kx7VtElNaNqK7OcIkkoZg0ZJyjJl6u0+zexlTda1IlcBO
GtL9zaZ3obgDm+q9OO+Np15FhonkhTnqoqxQVrUoNJrl73IuvL8XU7NJDct6Ay1e4qiqCSBokILB
AyUEtAnkf86cBKFL8+Bog4COTzJVugHrGC61PeJ4tBchlizVk0vzLcaANz00PGMQ/BVlSwCF2exD
+HnviecxKdEmngbqNy0MBvfYSym4bjd7kCDFSmFRb1LgdrGOv11G8+1QfuCx3mqB/5sMm/+8jJTa
f8dYs5Wrvk+VQjADf/yGPnQqrzgUYwHlX8H3Bi5nAorMCjhaGrEIEyrrMwV0bs9Jk/8EDG0jqOtB
BYEbOoGPuIDa4yHsVP2NvbDkW3SX1nCxWR2CDMlPaYWVfR/nkhwGsEtW/owkUU+kacR9Eu/IvJqH
uFWXpx3BKJwRx5AQmU0Kls7DcmtikhKNLWmI2VXWzMSpCNAl1i8T7SI/McUl4Vro7aYguAMMPpdI
vVHAFruwXFX/eaKMOWPAOqSZeFCHO923Ou2NoZvbhP3kS68P1UphdnEhNqq1UVYbxDD1eym23Ykx
ABFAasWOcco/xM0eqtmnvxBY87imD0U/N7l13/ZIZEd3WPsGpyqo6oIS3RAV5w5FVXGbRichC31R
4q/7z7d3BVfLJVOwj9e6rOBf4uG2n7BNBPX3rdN8FsoIdz+UenB1Ks0GfKtPA2DU2TWXLq9+iCx9
OhGAkSTW1TmiuJz9awrDG/+anRZV+oXNfAvqOU6X/PpHuUf0/1hVGi8NpmGmiSPxsB5p6RPne9i5
ziOmhg8hpgqbD75aQmoUpRKFrpEN4DMB6ZP+LKkjGQuAy2M0C+Uz21QZANsjrpwAw7HUOCwjLxU5
J5l5/JjlLHn8h42DOE142UB7zPbIPMLYJqOfndGoxYTn5I0g8cWKp+tIZPFGn8OScqzc96WeTDDi
XVlSoJjytPWvhtnJVjKpsglj/XqAUHWCuEBX+A/nEw2DtSGbqxfCyi7P9byCKS/Z/nG3bn/fgn2Y
Ry4j7oqbIFSCvHcQLEsb3h/FsrekoCFZ9Io+xcJ8WLBSb8UrV5zY1YVBvGBDiy/CXtrxk2uUN3eT
hZGt6DIG47TjgjHJRzf1SZZ/Gd2acYhcicgAlkIgLQJi3bmPyADy/j0vSmLouJJCzG128nKmy2S+
YLQYK6y6lPIplbRelcxzuB9ZSSwabVU56/5+fJgnnjvcHYnA9v3T6K2aFxVOVLspjYz5ne0RQmZz
3OjnNic2HsUbx+FDMjA9LWEAzG1KAz8uYt1axpK//Sz6y5GM0eymxzRYUCuUqv/D+qf0LjfOcDPE
vxopYF+qIApe2d2oiDHYRb3Qvscz74lU6bbYuMkAalPtrbuPiO8Cn7xr+Wq1L1jfgNPNxqxPGUjj
YUxwYmnkbxJbl80O4v+3m01jHezuvL8v8/Fd5rbEChVJnj44nMD1yppWO/+axFrfBovHfGDD7STH
qjQ4Um4cng/jamn/cyUtJrqOuLpCu6l4Nsa78ZiIoBwcOynkDqf9ULoRIeKOWqCDlzyisivKOXTJ
uN/qZ6/LK3fIJrLHiyCEFIgG/cjCMH6a0JHnrYjCuyR/BoZEg4IBx2m3pmFJ5bPi3B0F+eGYeLxy
yMS/yIAdQUbx+v4LfHufOJoxOqAogZGrWJKoYvPqk8+T4peGvbUDOvWgLvezdwxH+Di8z/g8KMYg
zCMJB2ioDe/5loUgedKtNUBsURgK6XbpnniaAr4Jh+j/MCattnj5+r3iTvP8fpFaKhpolKN2oYMH
VAjfo/Bs6WHMsWOOF8f0DIQPveMvt8z25hjJl71eoLFiALnd+0YYyb9dyki5GYx9xwbVy6J8BzMg
msE6tqFpc+V+p0v//9Ug1oScD9baocnG/urQ8/gGKOMgEqvrbsRpc6cVzS23DvA4KjBtDtsu+QxC
MTsUDkM7CIR5BtXFnpsFKGMMWRQwUlZ+wT2W/MsyfSp2rkwuzC4lZuL2mzdjLzInXEJRDqR5sX2T
KxT/acqLVBIgUy+xqjahU7nqnBRww+0v3rTbEA6acs+Eaz+iCzmNCQ/RH6B6u3ym9i3FQsIgR+wR
gjJKbcjfVu+czQu8MnuQWDKhhb2EX0UDVtErQfD9MQSi6utd+cWnsWr1ysQmXI00937KPzPdlDKn
TMULF6C8YMCVK6IHb8ZuyG6DS6mG2mYeT1Sm4Yp1/U1dsdvXslR29Zxkh1sXuQN2HcYcKhR2nSHB
cE1i7F+mZ/bNSKE+HJPnp8DzW+5FIea+HbhPC9qoc8pCRune6ppphlen4IN/r/gRAjMIT7Y7Ttt/
sHJfVy7YXvtaTJg4wndcAAwTULN4ozM51DD84VvEuiNpQhz9X6wusUH/khPvorHr9SmWsiKIEcdv
1r1EVj8up2D6i3TOjeoVMaYSEVFYOVebneE77bhss5muT5MPo9yvyK5+QPF1gx78ouQxscrrGGXv
lI8MOpOAH16imkD47DO9nRXkcUkEU4y4w8hMLN6Y79JuRB2uB33zPLJhpjDbZoI6KXGwxu5OLo/F
IfaGg0gXBfXqifYxFMDcdI7qCoXjDfQ8pY7dzzhVvil6BfaskrqF98u2j43bAIv8DODMWOVhRrX7
7nBWTp04i52yk5T5iuwJq+VhyhCQ5UzFlZRDpW9lJUqtb1A/10R+A0umhTTAdO3/miADX0QO+mgj
E+gqg1NQTVASQH0RIvRdvlYxFd+LZHa7Miv+VKcY9jq45SBM5c33vfYcvSlq3avSEy1XwBCUqFDt
wToybsbWu8gVVRUcPxJDhMq1jFNAtYTuFG9cAN/9I2uR5hefNfrvY62ipmLd3/PhGiqeZ1cfTFbK
FvJWEAzGqp1+Cs1zvFQG53SI0wCIXFaSiJrw86n5q8lJx0qOms9yQ7iFvpmiCA7SX3xufCsnj/L/
4N6job38Dttz27XlKxlu3jRDAmo5JC4D4BpRD4Oke48fu9rcj+8HxC5M9GR1ZU4cfQw8QeTdmV98
ydQUGBo/NMwiejtcE0+O02mtk+UjSKD5HlDgFremP1OZ75X5nY6xBDIIAsZspBVc3+hwhaT3yz1n
3S5k9rG/0azsHUN7WEMP0T2xSZETLKLupdTL4/9EhB2WmBIrbxf92IBwwb8XOSW6jVuUhYQQ0hdp
8DC9jrcFYhYt+GNPDfxq0RIGFPUs/ZEiFGVEVjtqKQs6VlMijgvsB4R9XjmI8r82Qk23wxmLddAB
fHKQX92kue1V9kNwdaeJvpAqp+xerBhPK7XcQqB3RPXcRppRIIOaFFtc1Fu69Uig71aSc9zkBPMZ
S531etWp8I//oE+2/eCFuCIVpQoKVS1k4LhxZAoLhvuRXlBcCUbau33X2ADOptgnTCcr/Iahg0L+
1IBwHMck22+YYkWLlkllwrmIfWMrXtdkLE6CnePB1Lh3Uq6HU3C/bCHhx2+TzoEOK7BbEqlkbCli
Xz7i8NBKfgVZ5B9QE+m3WRDBTD4i7luitUlHZV4OCqp57wjWlSxeJ1aIAqjqo/Mk6XiXUyUgUupO
cVF8nKSZNREF5Qcb9AmfG6ZPOMk+Kn5twDUkfVA7JJxW27CMcGbdL82EYXnE+aMfKH7Kc6jwubqb
OXwJfJUbrWuHVQwJgzAB87W9G/byfPeiQMlPSG0JpGi4j4fqvGBMqr6XD3tsMbDHn9U/oKTCN4Rv
ToHGlhFPPXGRIF09dW6XOnWQBeLN81XdI0hAuRGrav/uQdpAifVHh1pfH86x9sEIqUxs6IzE7Y3A
JX7EM3av8Ptyk51dd8djcH++eOWYkchttAL4oaHWR5jYU3naXsrWICjI7gR7yXU8rZ4AhVCWBCt7
zy5ehCYSkZtOUJZQ/Z0NShKMbw7q5B9/wv7iRGh/wc4NKjiDA+I040HxIRmuZA8C6nWD8Bb3J3L2
oD6KbOqZi3fYII0/p5rj+K3fweC0H/u0c/UqNm4grVaJpYFOjyDd9MxoB0akt7a8UYsI2i9vBtKQ
KxRV+wceG1e3P15Fa9B+sRyQOVQ8C0khPZMHh7c8ckCGket6nayM0AkDBo23Iu8tBymCwpN0IYMI
6B+ie+ZmxG+cc03OskEd8zaDM+8IhzZmYypzSF3MNF4jO7ZZMOGp8dQbW6XswTIFFdPq3TRsyfuw
LwEPykV7hS4xWzbzybS1ynT4W396VY4O5Q71UBCOQ8CV3KxCkvNm+BYxSLCzK9E5HQYWAbqh8WW0
cRMf6RyNGm0oSBKAD4blD0Ej3oBU8VkOzkiqQ8PuMs7fyB/hmee5A8UWkaC6Gdnnla002654veVo
E8EkuB4v8pDo97yZAJdaB0bwNZCOeF6rvlaaZC13DdYSiqvP86eZGamgronw/HOUNoVTpXq2y213
uJyctchy9TZ4aQ4Nlcs/lP8kbdmNy/wSPY/OoFHBnJzn6oJ9r5zmLmMgL4As+0fKWAWhUnAppT/J
OjDXjvHVZyi1Zjw+8xoZmFGAHPr64pv7gxeQtcA2KvEcGfh2RsrsrYed7xGVzBekYRT0z72hiHmR
LpY9FvRfkk2AYJOoiOKA3MiIFeMO87/VxkvTNBkJmfJaVfTnfARr1Dq+PNNLJzmeTGYBmscfuYZ8
S65GjqrLMHroEQ9CWoi3kL9JmlRVcROdRZmCZAAvPmb6iRDlplazwidzb+UD+EtUTrhVdzGzJUJk
g8FhpywJrwpWKI4rKTYzk/MfitveNLETkORauR78ift+Vqc7WABj+4/k9gnKxPXnzet6qWtO333S
bbydbrR07qJ8X3aZaM3YVoqghxI73d8zkFESgQCIS4rkmRHf/9urKO1pk8+blaGCUVYkaCm174Xf
jgGGJiUbvmu34vWnx8oZE2ObFV57oZ+mY6RyJZhB2c33yaFkzB9SsGit0Z3ROPQGQXWJN8jywpPM
CrmPKAY44FgKekly1l3/GtGL9qwEwVGLhR5hGLXswj7+jwuXb8ETT+YhSp5OXi/tzXXxatUIWeDy
xd1PC2iTLh+ARy6iO0oIUlukMTh/A2S4iEf0rgDGHZYuVG9noEYSZSaJI9SAJsMUjheFKjIG6QWS
N1hBhyYG5HDGxmoZTd+FSm+WahTTwOh2y30SmOQbVY1a28RW5gPsB/KlDgsXwY9ynpIw90D5X9Br
9NmeQ8w8rRN+cHzs/z8bPX0rFRyBvAtt2iQO9SF2it1Cwr7rEzlqBvPATjb5uXcv6KZY34sbn7fW
RdC1M+kxamn/uvdw3kE2wLhQo/bv+uMCOFNwLoZwfFYR0BVbYyt4hnhodQfwxhU/ahuyWLDpF+SL
WkmXWkOk6XZ2etQt4/79bVRWwcBX+vZnSr1glvHhMsdlDTFp4j9Q5FlTDal5WznsvHYn57Guo8iH
gL4gfH4WEQOlk1/9TEAaAsvb0qIOxgF1azqx59v9svUjQvHoQekziqcUMlnHxlF+UrNX0w3ZIVEB
/NCrqtI3z9R1X8pk65mArVdDOTsoWvri1Qun82PQCt5YVrkNT5Q8f92Fq+xSGp4lyoLn4upK3aLj
iIPtTclAvyZ3EDyAfvCj/FPA/rqVwlUoKolrYO0slBySHW+qTEDCd+Upb7as7/HoMFjVeZ4qTmM0
Jw4X02fQb0A7C1IVcM4d1nNcAEGYVpPpGwZofvwP9Kdr0aRi4/RAQT9LSbr8nyW2zJGMQIUb+ffP
kHaqAuVshYB+eqUHbgmj3EwasWS6SfJeyRPelNWYUQ1az3gkYZ+QHy6hJfgYtztYJIYmw8BAhV4M
+Sz2u2yPDU4tK50fmoA2hllW10+qNFmbgfmvKnPy63mm++VtUc4QEZ3B6GHg7x7PQ1e8DwoM262T
ABLDRVPt4AE7pffQ4J7rzJUK5eVmhYXDzChmZ8glaiT4FuZeh3bfeFPHi3eGlevZHo77QSiUAfpp
vvUP70zpRzYnWijGDCLjwPkTo688cdS1mNhZYUvkR4enqzKBRetnJHNeNG8BO6Wwk+VKFNq6/7c4
TNYcC5KFZvH/cs6FuM+6hTD2efCNGa6SqibF67DlvoBHdkIiL/I87yG8hrTtCHgSVOY4CCzCFDkA
5xtkuWLRkamJFJXqHcpLPSNTRpbzRW/JY6jF+VcJLtjxddi8an0dXODaF3OmpKUbm5KO5ZT9Bw2O
PU0mRECz2Pol+hTbd/ziIWCQvYBBAtwa0ZotF7iZjs2pzn8M7tYplrpbTr8fqAahTWNSpmqx1hMp
5fvKl8GTAk7zePrQadQlUT/u5dRtFtAkFs4IhTT39uQMjb7njgQEUUcMm15gO55PnnXstvvuBdG1
POjml8C6mJXRPuytrUbwAz5OsJnyimRmy6jdtjXtwkLwWgZti9ZlzwzqassQ4sxBIjcac7jjklqL
fFhkjtLGCTOcJES6+YBaUrjvLjoCzCLFj4qNKsfgpI4YgaTh2Pf3p5e0/WVFk0uz7CrwoJyCm3UK
5RYOYQIp8aDX4f8wvhgYwiWoChPJVcXyftmeOxMF7azrATHCYoxdtxsJaG0KclhmN+hBc1Q8tyBZ
tE2BmApstkfEfbZBO1KD8YUMd5AAld3blnVXPSFkpiRn/yhY37JsRHgGe627yeSWymc4HMzI6m8b
wFqxt3LOYBym3GeTpOTn8U3UejQYfRqYWIx5dG7hMB8/pnyVQxIWzSyhZjhZvxW39h2YNGimhDzM
d8RhoUvoqjWMxi/CcUTsTyyDGbbKccn3KzN6tkrAe0EI8lPQkbqwFqVGb6azNdz6EBhRFEnd+Njc
1u+XVba7neWO9EGtFWGghdIKxkpHBFIfmVD1B98yYI8sapC/qwzKlrGJpDBsBuJjwAKHTe1CulGB
r1VO9OhiSD3I/W9P5SAKspZjocvMk7QD2+0omwj0Z9QW88HLTlZTQmZGDqCLZOnahklYtQxUBFlu
iCa3U6A9Y9WyMYMiXD+olYpxSpkBryBpR7PPrFs4ggOLsgfNxawOAYK12TEQDc1SJdD40Swlvt0S
zkXIcTeSa8zvFUQXz5Sovt6d3douKvVgSkWyegRsVgosYfjV3h2jaLALCS+kG7godi1MxWhyebNx
gzJKNJO9fIxhCzjNdU+4Z6ftxEe6InCrw87zT4PpVnVIsD8yQ4WPgUjoHzXRu1XMgP0JueslxRdH
+6sm69UvgNiGY2alul4IB5UTnwdSoIQo0lRWH59In4vczB6/35IzD5I2hWOcbVZkEdsxR5TiFM/C
UL/pdCCLWb2PWLXt5gB+APAeMsYEN3WkKd4NNkKxzZZR49A8D6/uUwyLeAw9tWrkyP34KFnR6sX+
mXgjalsweo/YXEU8e7SdcebP4A2Mk+vl/62jjXap+iZCIzxAnk9KCiQhm4/g0rogrzRJSNYqgWVL
yWbE2yhRMVuo+8HbrHb+DTWZHXOp+NAAcMDpIULkk98imeLshWj/mr6OMlmvGLXKnecbrWDmnMqJ
iY9W4PBNdrHi2p7i4hc2thB1WrTHI0StmC07UxcjJP0JSzV0yB7v5DqzT135JQcR0ZVGLIkD7j2A
MGuZ9zb9TcTzuxEfHTl7ErR3xklBoq5Uk+CN5ulIE9gEQiOlKLsKOjAbu2cAV9D+cK9ixNNJrCk/
CUH72KFS1RGfja/wS6u+wJ3HIXMYgpkgn9KmXK5lQkh92kiAhGv9DjAXBniCuem4cE7DQ9q598FJ
oyWIIDC7RLeBLshdlYAETlmuC37WEZiyp4I35+8HVLtZ9KlCYDKaGj51z+MLIPnt+71QcUssdzWJ
fTRnHQRBL7eUW7AwbLbv7zllopnaBHqVfY56fIQtsdFdg7/dEixIUxIfzQSth/hg41JH0xR9pJrn
sN+mwJ/ts5NRipKEAlzeSSNMSIrhhZrYhGIdWfOhZ9iGS+f6E55tUVc+01zUd8FeAgCv2FBKe2hE
lgLGD1pJ+L4YQwzwHh4kaK1nP80mW8dxb7xer1yxYZAm5n02ggRphTrwtbcEm8dgwcL6SB9otsnX
k3uMKle6adE4Yby6EyT330pysnsW47sapmcTRaaC2G7PdaXNk3n2oukfIlSmPVPu0JWmOFOv8Og5
b1pG8SmzI2WHuF4wf5wraxBrPkgfWArSpNKGBFH1NdOrnlxKNjaR7kU15OjWg/eBRZuhYhU3HZsV
ifQYdiWHxvPYv52DZd9e003vE0qUrCA2xyy+OD4EFGdbhLJdGIf9iT7HRGXhWwi71woUn6Vja8Q7
BUbRK9MpMqhtnfr3TZVhzwU8g2LyyAw+rH8+NNfiqOIUgYbq2p8D/NPk3xCS8RaIYMi+mDPXb1wO
4bE7ccQ5WQS0LPSQPzXRN0iAlsm+jxNI9+3jCAZiiLduPTpKB5lgGiuERgO6mawiE+JtM98BVMTb
ylqh/TJ6+9xtiMZ+OZwgzTiJRoWpm+K2iyAFpXRnVqQQMy1nrvA3tBd4A+N6YOeVmFWDgwWhEr1Z
Q6KIibbKGfqQpzfTwI/Tw+v8+4DcGwGEbVzQnPcZiSnvdiUcArJBMzAKwddd9EeuYjYPm1XB29A3
jWGTr3SawhKTpijKl3EX9QlJgdlpwvJdGnmJ4/ByISNkTZpZEQaXqG9VjYfYvwT6UAxskWdY8hVw
hp+iWdng5Xs2pzUBIgv3DJ+DsV8My9lS52emIlIobs8RrYPlq3HhCPCMljECgi6yDUMrDt+5L/Fq
39pW2OEPO4ac+yieaElYeqBqc+XtjFM1Zd6+Y3fl2SyTb8RwVKjS6gU8XpI/pwuk6ZMrfcyZYLiG
OCvVDs+T9K0PbmUTBcGat9mx8pJNMeXK/ql1tKrVvX10y9PxgE8QoiI7PmNI9CAmcdrrTszJaX30
p1kdpGY1imeUpROpLFyolM4JbwcrS+xo0iw+quT5Pgsyc+KPsu+BZADDdj6xWxHrlzcVXapBDCKk
060Q7kL7+NrLqYbr4w6PIMnHOiiJdI7zS1OzPYoMhCgQMkCf3cZ2ZMqAahH2fqF3+Em//8DrFtaQ
Dd/wisu7gLGK6pPZJEhE/sn2N04Xf+6LYUQ5aPXniRaD2KrxHQfjxuEK+DgS2fNeKkph61Gi9s65
EnXK55wbQQ48gBwl/xS0mamdznXdYYJtafFpit8rRTpxV3vKJN3VmTVGoqoKcl8nQ91q87oWEC8r
7hJ6xfRO6fEcUR9jvnIbPh+xrn+Hmf/tubJe9p50TzCTayZ1SQtDvxvfSr0h9iQ8nLdMpWgAjroo
SUzkcS5qa/uolRn759+J+4naJ44BcZ7tuBW4P/DAlKGlD7CxasXytcQs11gGi2dYUyLD2AJXN199
0jKO6rb6yFIyZmDc15nGIFwxnkO5CkLYbkg+gmHgEXOqtIqQwGanRsnG7lPCTLmAKukYurPjlHwB
zioYglvoGCMk8RdgBwJwD00V1TxyCNcAgQv354OM4gTXp7J0PVW1Ns+EiDbQ6f66kv8IhRdEjra+
npoGPHfNo3ArqE0y7yXEP9YlL830nr4T/70/qjjbj8mRLw9rPYm/J4GMOEA1V4Fs4gjsdTEeKDZT
IVW8w2e6eSONoC1o8Smnhd4edF7eihLg4d8dTTJNOSeTCyUautRj1ObiVMWSv+4nz5SVYljPco0H
D8LntDwJgaF9vK1bS1DS7VkS+Z56fLS3Cdbf6dXGBgHXJ/g/zOMTz1DE++HXHpojBbvog5r9Y7ix
Y/2vhlQxeDO7qqIkQcERrVHCPtZU4cOcsJ5G+GDtvXcVj7d8DxjCXppjHXio+BEyDIO0pq/Yztzn
LkuiFS+44RdSUQZPoMr9vDum2DJuwS58vjlJojnCEeP0NpTIGmRjRvdX41vq2b1WUp1fxD8UgvZa
KGTSInnB1P/kBZ79xAtBvBZglv21jFvMAaRFCoosR0nESkB6PXI9xgac+dZkT/CNBP6HZzmA4J0u
34Ik8GvoSgA+rTbrA3+oXEblpZ+pLl4F56Mb/hgyTKhYKO0xfWkvRRvub4+/Urks8OWdG59xYvBo
AaOIH/tE+IPVQ8AXXEzio2VSZzE8lr8stNq+B21UBh41B+xCvAhjbWAZZIDSXmwznP1JTNs6Qi9v
9Fg2xMYoY5W9VVm52Lr+CAK0OGnnyBo8PaFXNm51eFaSJP7klUdjwNHVtY/V3NcL0Q5Zpfwhev4m
8Iew+l1jhucVU7A0EXH/TW5fJ0nKcwB0bovvnF4e0ReuWizeSnyJHKYgws4iQQWRa4W//j8Bm2sn
CnHSXkEzkVDdk/OQyz/31oCFC+MKTaO5Jr9u86YPy9S5mAly0vUNUHOGRFWRzdVQd49Gizf6ZA8s
rPkIf0EcVK0VFgr5YainIldN02CbaZjKgRK/v9pvWQB0QbSJ+x7s/o2vqm5xx23wJ8I9HF6gVcrr
qLZr23xSsxRTtjmTO0mZ9x6kK92CYkVWd3VEHJAJ9t4MgIteqiAw9XRzH2oa9/XeFQqPSz8qTxaP
Qw8xub6atyA8W54ZGaxlTjQ0IYt+h28F6oQ19y0QwQAgpFzkOnutVxhfUKNmGnh9ehD9ydscdMsk
JqO+LtvAzxFzO35/cYu9SWKUszQslE5oBZ9ucbEJ1QrT3qvtQRWrCg/k2MJB0neU/9h1Xsn12VY1
3k/givIo7QdT6QBlro7J93mdYD2k3+bLasRsZYQHU6oLnlt8lQ3/eLSYiaugxQZFAdhUVqjmI2dX
53OQqryj/HRNI5u20ZVhyQrPiv7YqDH0YKXOFf4KNpySGvovaFjYlVn0mPyy3/4n8L4QWPhDbgRP
bd9s3kUyf2IaYulWNHK/O7yoB3x/aV4y4+Zk2meuQuCXFEcEFp/9E8eYlJKI47PICOlXJvQU/54f
rrVZ+t3h1cqm7DtOprcV1bT8qJuR9FyMjzREBYML28r90i8kxjDp1Kmthxj5fkg6uSrxpVr47zN0
vLhOY79sZ88CLrpI0AophVVW31E2r8JXhAeE80t980MkcIxtkcAsa7Bv2sux2+7YVUnW6pHy/M4U
ZumX7Ar1qUjfwMklZaOezDWXQMbp6tCBOu48nXUWc1UHSGlySSYC2O+rrGxaG9KLvmfHLMyhhJZX
zoiz4IlLV0XYKUNKXzkRrwGfJR7h0kGjBFC9I48R2vHyWddr/g9lZhPvbx7zyONFbekSnjjLWuaT
ogyP5CluFkrdnfbcGYAYpbLInJYyu0B0Vv3GzbRbK9zS4I/VHoYJT3j7xjmeT+E6gUDW9EKBByZU
rSWtMoCvZOfnlvqGMRoy4Vw7peKelDdhuGNfKXnGmYDIMDy5wisGN6tC8LOO2L+zaVm5GLxafoPy
hoPitXXY5F+wobRaslJiHu7zlShRpN9sxq9CAFzxL6InOZtpNcKt/++vHZ+PwAhaP1p/n6wfWO+0
45BRZdYOfF//mIlVB8nQmFPVhrGrvhQ/EankyWP7U30SpJVQD8BJyC7oYFhRu75FOEIrhEhVG7TX
lECsA7YPXj3vZ3MZr2KmewwxPW65iB1UpDTLIIegXaFeZIvOCG9z2ueFZaok03sk7eDwHXv52P/5
g8/CNbmML8xnfh60ooWPe2kDn3XkPGTCkqScR5vPAxRYcul9Ew17xxBLexCcai2/y/026pyeu0So
F1hKHqJJj+L5Yicvloq2lZEytMUjNuklMjuuDfhRfzENgOgYF65XWPQIr++QWFbt5/OoNA1GWKJ5
rnFZPVv63Ww2H9ys30cBnQOs+sutYPiIV9BwIHcXjr+97xX+PWFwTGeF68O5mja5KlXPKKy/eODW
VUN+iyAUJyryW3HXHvSazb1sF/o30MFDIXhJgtNDRybnpRYig03TBJVsnEDezWcBQv0j1HiHN3Rt
G4+urMIH2mf2kiSDt1UVPyZ5ACxye1AATKn8JkA/c+ggLBDIFuIYxfumRIRPhY+qPFIvFwNIEKDM
cT3BiLXfPCxxAIbbq5qtVhIEsgP+576JWM6nqvvaMNAtqS5z6mXbp73hFbqQuhCUW6GxLN9jsky9
ZD+K71PX9mQu/YeW8mGljIbCVHmORdypm30xOxaOb2PuGdZqRHED4x6PXydNZ/UVrBW8UjgvGWgz
+DG2NfQBhFHH9IXiRmXROosNnT78QOzAjP8ozXNRC0Y1SQSBuevHwi+fZcH/6FylK2FloiqKOncn
nwak0ps/pperPMyPXth12AvAkpaOQHY4bpFuyHOYwnmlvRgDcMKJplvxxpO7Fch03mjD8BhDAr4q
G4rV/fgQPBLLCVJxQob+GidHPIvg3MTukuNkE1BzQxrh8EbpkDCwqQAZjq4bEHI834AIQj1kH2e7
kYJS97ZN7D7q0xu/UomB99wPSC38Hh8hYh9eRIj4TfCFZLyfyVWz+owzv0xJ+UR0Ti360vJCWOyj
W89ltIhZsSdkKT3C1/rNWYuOB+NwCr5ULgx8jULoqzpblGZ32HutVdEnC0kBcMQFFP21mzs8Nqwl
2K2kb8vyNyymy4jAqB4Jzbzur9bSXyIGwLgsuVKV0DdqTgTd5aItEPWe5a7glu80qRj1VGswJGio
blIBq3NeMhl1GOt97nK5IKwBZS9hKsaMExOitCX877SyK/McrqyxB5wUahsBi1kDpD0tmInNQ2I6
LzBhynrDsrrlG1c+8yfNKBEeE9B0U3Z/2Kc0EigoxJl8HYBcbdjRuSqGXB7aoBFLCoeytL9DWGnA
CiheF1lFqSD6balw4/XL4J0MUYdL/DwniYT969YOqoqlw0KvEhaAfYxSB9U7ThZIbXzIP0ko3scS
WP/6lWRQ0iCPgvjH7hwKfZfH7FsuNr7fgIa/B6LgrrbhRDlf7+BVbLAXoWhZ8w5BdYzU3oMn+mX1
qxWdC1mrTBiv4UpS3AviyT8tOjjkp3IxQA4OROio9T5oa/m8/4lu7suyBYYieN34WzR5L1YzrnT6
+06+2CsLK5sLDhpE+FtClWI46PcuWaOzkwAydBHsz1e8hE4BcRXYm2zmV1yghWDIi62YkoyunCA0
/t1Bjk/+upjL9yDdtTxQUGhkQTbZ6L69hEmuRRHoudk55ajcMPOHZvjFZ9Ds9tptBqv2upvdikWI
w9RjFruNE7NqPl0T8PSmuBNEibAAOnhQ37muqOFzxiGzZrsmdyTtZey0mFFmzheOg/wRPQ53+LR1
n2MLb5dALTXNGYp+/ON2M/uokPUijSOjwL7gO8vv3G+FkPy1EQGCMxKOUBrpCeEfXi+fKSASTq72
WLPqHw2CCmYn1b42JbcqzoBXJLCFFn6VCeSQ93pA9gmTGShKDox+JyPdbDDV1nvyyGl6rVRwhP2Y
ICY/j6IlC8TkA0Gx7eulKx9bLfiNCn1wxnuQ5/8bNgLB16AVIsc+vaVzINXOQqaXaHy3CNJNR9hb
eaKBSQGcCnQeyHy0+4FuVkeOtaabjcAr+wxKl3TJUcKTASFhHk7WcuxY6nIsLTAgNLr1/wGp0d/7
2tp/fTY7rb5Ur+UKlqeTRZ1bVhkyTOHEQz1xoj8SZmoa9QskbpdI08T2zxUo7l4ZgHjT8JtU9fPo
+1T7KOE3CXwUdxGc+wP48a3fvecXfzOQZ9tFOB2/bIXGdbJYyMvc66ZADPamusCZHjWwzSkW90nP
5kERlB7hf7SD6xLpTOwjBd6r1rF6Fq0BYpAVtJgVebuiNfnFV0+xZ/Xz7DvMj6U1hja9nbBCSWnj
rRPVD55GuAN3HdB5lSQ59d6KBG2bIlZs+0vyNngyAkO4yy5ZKC44v6sqkMkHH7z7PxAh6ksUdfov
xmq5/CP/w7V4lBS0pW/Wz4DBqF7K15RK2rzgcar2CZtpuIVGe8h3GAnDVQd4gQAS5KrYmxALcA21
iHvV7FdwB6KZD4j1x+4w9PBQmkhDJHpwlcNR0++xiKctR8Ld5XNXbQh+TagBO7kBC7AD/U6mq8B/
7mjzIxD0k8xRVmyrqP25am3eWi5z2vHwoUV3nemKLUDlrP23J1YOPtWyOq04pHT8pBAmauMFyLMR
kO8y9goGBRt8v2+Opyo5ZaZO3WtJatbi4OhOXGoTQ+u6OJlCU6JpLUsoR+d4vKw2X0CMLpKxHGXz
vpMdwSwFOOQjJx77kltqkOD2ElnPtMiMCJeM9+Uz+lOCPzlBR8SkQYqiYNCqmqhP1rRImYOp2BbM
6jBvt24FBMN+BKxbmxDORVMcYFudBZ8UrLb9CXN6dRTG7NB0TwSstyEJRASsoi4n7O5Ujcf0+Qix
FKRa9Jp6lPAO3DxMUhLnl0PfpiAficN/5h45B70yxWKEzexZf4+Up7TVKkiC56/H6+LfLwMf6fnI
EMnGLwdS9+cNMuhR49TqXc5kHSpq1y3a+LVlzKVlaRjRRqQp9H/xzsZaq0XVK5yhRUVq3qHGjXa/
rg0Te46E5meCDOCUQVkUy/L80D4/7hGjczQPkslMJY55CdpnCvdQ2CR9z2AXx4F4bCbI/hCkn3Cl
1zOQYmO1rvjPU1jqQLsOlr+qdZW8kacAQQ49kesC4yJ9/bPUVIFTKnP/5zyUb/SVIx9+/T8AxY+X
fDuK3z8C0LgWXYbR39jUEC0tDrA901TEmE+N0+IjMKkIV7v5rSb5Lmzay41dcXbEHm91PF2jT+t3
ty8b0KQ8tEzTSM4vbAi936Bl8F9xe/yudsvdglLf1jD6PnynYXlQ1IrEPlbijIZVjlaEc7bylpCN
/1A1OgmMpWeQ0fz8ytFPaQbS5jdX1WCA8FYrqoRZmnv+1izNDOHeksJuxJQiQHUvSCH5UfGTGI+A
GYJaSzj38Bkprt5aIQrpOW1yKw/ACRZFM2hHLk/wRwgLuYoK9xVbtLpK9miaTyuZNxZHyj9NebRc
eBMV094YgMHzTjgJjXUaYubBh0Z4F8WVn6r5gRlwHuxB09Clnlz/BbA8G23ug3ZuZL50g1TiIUWB
ughyRObVVV0Eg+D7vvU/mcXGMuS6N7stadPrrcxydmclokd/LvBwTbuz2hVIKPktCow6BbIa4c7t
iLPXUeHbokCEN+9t84e2M4K18BdLqeJX2wccml9Z9/SrtKnbdMgLqm8uKfq7FMnqG9szNDLmM81q
tJ1h+wK7n1LOkrFBQoEioIi2+z5VCUQEW7//WldEvmBmuPY+uwoBhVRbjyvnQBuPWnuEq3QholbJ
+tmNGTr6HqYbNs2qc4e1V2rVNTFgMEgLG3IC1/s8ad17wPC7/3ySdVDsY2sJkoxixBwg8T8ALgqn
mz/5qhFNTMS5EjLLLKDO5iVm21L0p1ksOG4qy6Jm3jBUBFxT/+CmK/MloiEefrsnqPsVVxyqcrgw
AlTpyJiI7w8+qDjxw2qHp7XVuHvVWLxG/+0H+0/mWljbDUbdT6Qj0n/l57huuha3CINrCViaWvsP
osLBeKdU0yqzQrgwXHYETNdoyAftItK+uJzSUfcEG2LhX5ItMhMPbnKZiCdHpapNsb9U91cfQi9d
pfLJRc06ztji8MnBRIIuiuOaTsBIxH4J5oWE/XZqszIcWwxJyOdfeEPmF4QX8MA6EszqM3ha204z
+CvrzIJieMU80ChhR3kQzV9KjzW1fLMFZ5jY8kQcJd9y10d+GKF3WPaue9uv+oCYOGZ18II6go7L
irjo/Bqvf7S2VSUpP7+9VUxRQYNurnk2dW6io3W50uyGLIbwAm4LJPO2F3rx3iQiww4NNjxT4e7/
g5EACtkTi+fqN7NChNPZcNHCwfhCtMHLbKEc5t83eEWjlK1P25DhtXbndUWpixXRHjVDyDYmFYLV
VvXtfPOQBD976kD6qAH+63+KOhZiYuG0sMnJhuSehsmLwE/Jq34GZ/F0No3KNUhjBPJC3liY7/2Q
kKq1L2dR7pnsA+TLMhmS2Tb1NXrL+KNMdkLD+SGDuY2wn0uV0tPgDGnSklBAEofQYMAZHRNtqPIj
1OXXgFtSBiBtSosD/Vhj4hd2UDyE4sXZevYJMxAj3QwkJ0ur6vzWE39E93aDhoBjVM4zGpPlL3Xu
ZOfHWs7x3Uov0l6M/vWQL1LY2adTXeJZaXZIapzTewxU+DXrNsX2JZIMIoJ6DxrblqgJjb4dmPN/
W/dFyJ8PyE88UiRREl2TTjvUDhy7stBfL05x4Iifxc7qmXZvrPnpZaV/S5Jfh4pBZ7qVynMTDv72
JBowGSNkcmS/2vNav6O6jdu9oD/8dNgECWbTIaUvL9Jo8USaMG/IMppVTNG9esCz++TdQ0dZ/mvT
5R/MUPbjrzTRU2FHB1q18Yp2ip4xQF9kN4PPWaNcruQsEhNdNkPyBetmg62yeyDsE3oW5ch+vbfr
aPMPGOO+wc5ivkrNFGJAzS1Mii5TvhZ1kl1ESojedOpZgRXJxhGZG23/rvYq/ETDX5bLTfPDb0Nj
4bYMCXNw2LXhcuzcydmWzuq3UH5vxepOfXnz6FspH7Gqi+322J0mJT6iHYqZzTAhyo20UOLNncBj
I1KlffMEVLTfbwSKwl3jycS6GOtqCCUO+OyGaN+135bTI6oGUKwTdiG8eyXul8OvwdVh8iDSh7Fl
QW3e+mOK7dlujzT6QcogXJwlQST2/U71l4H+8cj+9cf3HT4FN72KmrJ1TKbud6HIAWqJNzWvZwB/
VwdxM6tcgQ1tbiYVUO3gdb9YDWI5EpMN/6Z3sdxdv8ORWY7WQZ/zk1IUmvTQL6CB6hE60iVNl5FU
oMt3V5ip1bN96Uamu5oOofHIAswuEgLrqJKQMbULHgn/EwpD/wV4mc7Tfo7CPlXwOkL5SbTxHYW7
cUo/u4TnhbBwcUmKrg+MsbQgN7gRC0dI+8yna8E8GQ8SxJHdVP55w21YimI9+r0ipJTc6SAFmzMc
dTMXmY6x0pac8rub0y4SYX2vZTZZ7F0NIQ/YoTxs9K55i7VZ8nSnnWP0s1Ueh85kUF0199CcEz77
JGrn5j68BWHhuBUfHaBF910wdyuP/Ejk8BcmtOy3GOfz71nJBy3iRWjLkB9TpWsy6c35PKqlJkz2
trfEjFsSJP+GIAkkTb6CDLwp8AY0Ef7vMX5Xsw6OfJ8EaybHXogNQV/HYPvauHPMVcZCUcfL9kWe
UHPZayQZgX9C5FS0FtTX5yBJwJ1BRIo58CuBKKKB3+NyYQOj9xZrFLicmoF0nA7ZiV9KQGMKjD6b
8E38fr+8HndJf2WfOnk6bRexcZOCVRUT/iqPqoGaH2lkXxZhrbBKCYJ8bcQaSd1a3iguDsr+Czph
yGY5DaCl1QgqLiLDfcrtclW7F8AEsr0Hpw2NeJyOSVq7Rgq+5UftU9Ti3HKSo5N6tvyvtolBZolQ
k+V0RD/4wEel9m065TH5KhYwjUxpQ5qHuBFecXDeqe0BStlrCWWEStNTsc6yz/bOvfr5MLMSVVRH
xnHmv6CTK466tKHaDtfNwRSOHl4/IAiv5ySStY5OCZomCdRhOyP0+NhL0xe31wlejx+xIiJHLTlx
0v3R9q3O1S9PqToBm+32QOkSJETzOQmjmohHfXhjdSrF+Hj+oN2hSFhms+h3tSXU9kbhpRpo7R0r
+7TMEZaf4XO1iS04fnVP0FFZ33zyttE4Wy9MAeTQOp3hfHqj19MrSqYZaUB7TDYS1W2pgeYFR9Ix
dkU9mIbgooxY2BZFCSOuV98tn2RviK5fkS0+OGT5zVQf6BmAzJvSUyL8RgeKacnfDn7Jif71lycz
Kd96z5PrqTII/u6jZoE0Nd3mZI49dZ6VhoZJsZmowBcnLUr5jBO/SprJpT6j/kR4tglV9p2Ih3DC
yZoNsKnsk4dxvURc8dLVj88/8BYcM5d8G456RIT3M0fUQMkPPh1HmO3q1CQxUj3oQEQP+MiqLOIX
DE2fuBoIiZXCtvA2ICelFJAlm4cc+s5o0B3caYmKgkXxMoy97skC9UtJTAAqWcIbowHQDEs/ma4x
2k652XlBPx1YLXtYiHcCNMCdlcbPjXTYWJcSth4QO4wqO8BRMqcRaHrMtG8DYAYOvHGNL/EB1Nbz
iRxSXbZ6GIUkKrkuTtdFLcW85g0WvE/jv5oUNnJROjXyWefaYWH5nHhKqXy+OhMDj8wAIs2b4zGc
ZTIq7iJ5cGqW/GC/o+1bzJASqApzEr+JFzVWIT54/uysXDwHKkd2Jm8tuXe2Y1f2cZM8+oCbn5XT
t/CFoBrg9KyQR7cjpOuVIEJRSjasiofH3UgGUlSn0UWx7yF0H+zuTEHBi8gfR8tMBYVBNmGZ0Z+D
oBZIKtAA+CJlpOm0jrRHowx0JH1jHUYJR8BT94VpRCiVZ/rxYnO4ZkeCkaVQ2FOOGfgqWRrRTmEY
SRrUlWKcsvbKVvJn3wo4DzBGC31sXKY0Wsl33zBgDF6HXs60EdeSbRa27fPBn4rMh3PmaHO5S8BE
s+J2PmANBaJ7QDnK146yxCrwHeps6VdpnWrj0OFW/fnwNyMgbgifb2Qc5tZ8c5y4MWrm9Loyficm
itLKuBO1wQQOa1QrnWp/SjHgAx7ZZ8FEhTY+Q31zoFUvUUWSUV4ksdjZ7pbv/whtOhm11RVPWFl5
cyH4/IJMMMOP6JiYEHrCWbfpiY8UNbOpz5Kspw4BAnHOzHkPtmfhisSD3CfiKLVbV9BTOalDa5cU
n9ZQi0+z8w0S5YNSyaNRH6N7Mr/92N7TQEd6iMvk6YgAX5Z54XjBY0mrUXkOZTRUakcksy8b8iSg
LfdbtKJdKZwrQksXZriZ4MrFXJR0r69nyoGbfsnE6VBNzXHGW2NPBomM+QSe0cuCHFhcrjug+NXi
bJh4AHSN3vP1J/rI7FjSFeYPSsJ6KWi2vVqw2azHTE0K8iuXubFKydWKsYKSkfzAweXI6pF+V9f4
dmZHLIhlTthH1l+nGuE4jcH89NaWrMicRWYQC/wZYJOB66le8BXzgTm3WzGE2edco5UKNGWiwooT
96Lh1Zif+dPiqgwoCf1+bBjsC6oIgFvAl7JV791gKLKtMjojL/bNLaFCXeOjdmdx91vndA4I/8BT
jqDwQOGYIq0X5LVCrdEFpw7rDCoA0f4aTk1xNRnQBo+w8lw5pGOL454l2B31DOrFMLvxuL0lZuId
ERiSHNsA3d67Ahv8zPvcMncuJJ4AxuJ3heXCe44FtdSfn2nTyEkM/UVm8xCQ4bH6wsKAbu8kWvgc
ncDV+0HpFpRcRt2m4J0P8/CUcmlG4vXSd0+TC+STiZ9a69jKMtZqroFLeIBI7PDIiMaMdbwMuTCB
TMeEb7VXBfhOZgwlrKhTOtRb1sdbP1dUFidtIYYzWPFRYshxDEGELzCfILt8rZF5iVSVSbvOH17Y
VkAmJjQPZAHW1Re96pp/b3cWQKf+mCufCxdJNvZc9DBolzPO6c7lM8rxQ/mXvEh4dddpPDxBN1YA
7hb5CnPUv0VNush7dNfPCRTKE2p2L50Pj44yVS1TgnbJTkC0vKH105zWqZnR8E1gmMr41v0nUsB7
bnkAYuutMFGS98rixxwhGV7Bb97xjTE9o0f+vs/faxvs5kGFHhG4YPzVOhZvciGEARuaO6mBO2Rp
hlDnbnst3dY15Otax8s05EumeupIA6ZezA1q8oDCBc7qLpedFOjGtFBaVyJbD1b2IR34ifE0gCn9
gGaDQh4vZRrjo+xm2WcwrqvkHusmsO5YLj1h6Rm9Oi8hOaQR1bDMWwvRbmuZYq7iEGi1PPb2szIX
VXA7YD4JZrmv4O6+TS3cisxVfSt6WoLftTEqLOMYwQpnP1WszQQFWxCw6RTw9ZGrnpZlAX05td2O
NGuXHz/QrkNd+Xoq3D+Yk4TRSczvgnKsF6fccOJEN0jlU9O8VfM4U0Ne87Ls8sjme4xs3qNN7KEg
roAK20QfqQsjnjTNV4XcwmOh1Zns2Tb82kkgLtiwI01cJ3UfmeBWFlPp0gX2CARgEwy7Yzh5UUpS
U1J/s8JDL5JqkJW+NXvUzyl6OGwncaCXFjUyrIpc4iP/3mH08x4GgsQM14JXfAPNFtd96AKAOWdu
nH12WfI63lgxjjjxzzJmeNeaS/AwfI2rqVTcgE272GO9RosQoiuX/j0PyQv9TYTvdLvGiSHh+MPI
dZcCQwRDil0hDie7TOCuuqfCN3fDd8tfjEeaiIzq3BRHabd5b8R8k08i62ERGonFdPMAb+GycXMw
lLcKId26SDM8ZS39St6Sq/Eg6Fs9Wldrr4601G9DXQKb8MhYI8Lkoo5V0+pFRqPGjiuIK4rcg/LN
poyqPR1dqI3K7GNgpQkmrruWIiJMUHijhvqWRbSiXsC3nkoGjOW3DZ2WB3o7Nwln2eQS0IxqxFmw
EvQA5FZjgQqZoRmQsSKYOlD/Sa/49trdrE4W419mo/LiUxLt0xdx8DkP6ChcPJBrLfdiCAc/plUx
Wf0mz3CvNHT4bD8pzIALdfdHtbYrFMxSJY77wd8V0HnDTDfMLKq2OkDl2siySbQ//39AYGPS22Y7
hXN409TvUI3MuJDyVUd2vH9zHTDzK+bm8Ag38qqpaKmVCkFDleUDqRQJBC/WHvHc8DwrP0UX14ai
6AHiCnz3Z5qpUk5B1OO4ZD7SwRaolZljTqVU+VtWYGesaVUnqpQ3PV5AgTrzpQr0sbjoAT25vNb2
KrndqqhXt5eAPBWdHkkhq/lcFsdeyBBc5E5vKBqyWFb5CIdpGlVbUmGflUitUWrCwyrtDzAq522/
1bJD9H6zy5IDs524ewRQFHybN7B4u/yYUz2J4TlAiX4k7Gt597bIpCE8Eyh/liHPPuxL/HWS9V3z
FNqqF3YrQgrXXckR561YwDw/ACa4bEStTXWag6JsQNPbOFiBBb2S0Qa52hjIMei/yP6pFWf5H6hm
zuAfDXW69jckElKIFqi+VkOrbMMWhwtUILv0P08G2zd2EIHEG4ZdYt45TVCFYUCPMNGhj1eWR3Eo
vjPc6imS279bbgB2mduVJiBOuiFv6xZiCsFaQOz76PBCJczkAubZgmkjPjs1IMx+WdXnEiCD8DSs
SnxjXyVyB7QIjwAJV+tloMxAaK+dBKKRt6RoZRmtGatn/VbRc2F4TnzJCL/5fr/icxy7q/JxdkoI
/oy6Mgb7QtJoRjSmJWSAJlRay4qzK8Hzjdu3NITWD+UXCJszJETxD3/SoyAuEcIAU5Fg263Khmro
6zIGcPbXxXfi+21t6BRHOElSje07utNaRornMkMu2OH3lHSzDkJ81aEImDUhcNb3jTcLk0G379eZ
tm09ary5Rc8YyQqVcuCupwpKrHBQHZag2czD9GIdx3WaEx2G1EwgN3Krk0JzWmn2aZ4DZYdNc0wG
yE0JkEUI9qD8/yIwpqjOJPvBJTaKp7Wgqc8D7paRZSHtDzqb8t/8eUBsYElTix5c3TqKaPyvXQwS
o59XMHBfTAXk4LPjRDMTx8Rv/xdaFUsjdYzfIJDGdZrHAkIfxoRfPDmaeh1NYgAJLBoXu9GvLQ7J
5dfQnG9HSFHzYbeenAlmPY+qnRI1rjZZtLk7yOHZjGpEa+UKCg5Dqx7J5zw4SkgrU5g/Rn9Bl3oM
sWKzYA9l6ARmnW/muLDvT3feXEmnFTPTjPLHosZg91CQZfiSsO6j7pAbyFqESX80ERNR4djqOGLD
Ui13LlKwKXkeibOInpE/ii1Ntf14+ZtLblQ/U4V2jsYGmqnlfYJT/sbCeGmkV/lHxC7juXO7L4Qz
hzNSyr3LPUE993K/NRSt8qPNciI4LnXoSFBz745mgBYdh+5uvc6Ag7gHhOW4+/Kd0EMFQsSQ/RHV
QymcCyvbvql1L+AwC3ufOTH/wYct3un2cna9e+mQ2Zt7i62BFQBZ2DZvPZSuxh86wc5WxKT2d5T4
FpiyEDanQQyTZxjinXbeUe9LmwbxxGIEfTMGvVLe34JQlaMgpJ5xeg1I0XQA+dbQYxqCLYK2g85g
oXgUjZnGZf3ha7B8mnWRUszUO/JCx/VH72zT0u4rdAnDb51Z7NCZjZqb6aT96pPLQJcfEJJH8RPy
gCdEAvw2pynbgIXyDipzwzEk0SevOJuWLdn2LY2EMysHQNuv9FEXSBfNbAzsTAWRhHJMf0+DlJJP
ZhrpM+ZK4EWsfTQAtKgFrdA/XJ3g4pNF2DO8CWJGReoYDke/bUXJz/SrunzT5qy58fxRYrYcANex
Ututf62iwwFaCXhKWib8+87YSNhUKZvRUrmRswFx2v3tChVKaz9M0rWaq3sLtOKnnJcvEyftuopw
O4lRyPowD2rOdQRi+PWgAjVIvkMvuI9mGmsiJOlHNobVzgqly89kDFBZU246++KdWU4rA7OpreWQ
wxWtOI3DdSryvZWPh8O1+WI0/sP5ALh754pDNTNSQ20vCWPzRNs14UbK4Zm+je8Tug3E0oojX1E+
0SWqlHLROvlKAoy1xqWGKWRUQbfopIsPF7uivYLdJ0LYeIxZiv3a9Ge25REXCtlEjF/XfxQ6FLtD
QtRu56mqGnq2h0H6ZyrB53Eqg71Pe2kx+WpDa205l7d7fPKY+V5jPWZDrkPP1ALOJtjSFZfWusNU
sv4TZ/P37IXW3cjeeclSYrhFWxCF6eW7ylZYvrADV5SQ5gbNV/8HwS4C9D+PBD9M9BKMlifvZ/6k
d/VBaTyzesdXqfQ6lKolXbF6nAcJrV0hw48vQwWKZljh0bmGWDrXi124zc/xaUJM8m1uPvTMsbrQ
XKJa7U9Qulda8CyNJWIYYorQOhN1+EaM6ob7SRO9UQ+B4AdRmc83ko71S8un8U12S+InCm6D/jSm
LBfpTK10udNYQUhHcz2m+OZZwZqfhtWBHRfXJbdyLkaLc1ZSdPkpaKQSGL6OgP63a3yoCeuWC6vn
t5aNDaFr88/9ZjEPeOQZGSWpKyrE3YWpC1UKPzR5a2baAV+qweljZ7V5KXxcLffW/0Xr/h+nFf4p
dytk9s1lAIOSP+xmb3YZNTqw+o1DsgDfFSTkpdSm0VegcHDa5JR6LCBBb8N394hs5+0JrUVrLIQm
HmEz0XzgeZvmF0KXwRFo5K0BWaORfqZAGXeHKrqViqs1C/gurRZbfnYNzJ7Djbe1KWC1Vxm+x7mQ
Jdx70N+m/2BZGeU8d4Y0Ii37zyNTlpDVdm5/zZm8+a1Rr8Dlt2KjOi+7LsV8rWnMnXnTxAU6ZzWs
OVJz7zcFOytG6G8Mpt8pzZgBQfsaKhtonzcV2nPEWRK1RJNToJCg3x3X+lrvcq+BMsRVFSsLqomD
1euUwnykC0RrCMOy+CZBtchzROTgWL28fJnVvDt6PTZbgUupwXaAJPImkCig7y50ag4Sz/tKpnk0
fz3foBSbrLYIE2ufD/CF+PRUpv1YfJb2o0QagsWFlxSpStjpfqyRFTZ7M4iH+YWBsljfaBoLj7x8
XD4lhx46Yx9lKjGtpvGQzrgkXCx2yKtdUviEIo37RoWNIkCbCq6+QtSMGXukmZt0+RGUQqtHtJtc
xBvL661Q01itm7C3H1pylBWjCwi6Fk2T5u8xTMzrvhMlZGBbcD1mLpC01dhkLzQgrVLTkYpXkv1z
0eJKl8HCVCbYoAaDOvvrlozTO/bsRwSNqaE+ICkNOVKiAJx0q1WZny1kiRJUUvoGFv5ZgkcKwy8G
TlUb+Qo2OsMMO89qaBibRqpOQquY7VF2LgxbZ3tBKlFg9aGE/h/49lenzMamPlHIzIasAWEU7FNl
+fpgww1s1dMbAIqgeBVNS4k07CD0Xb9KUzG4SkPxwu0/lK5KrPP4Jp9UfFnccuqG3l01BTvDoUZO
YFeBcaplZF90RmlP1S4aoo+8mzlCH0yabe38SHBfRBxSY4MW/Dd6nVvQOAVI68wd23BBJsOpCS6b
162GpkUB5wT5SEwxcywVQV0sNNUy0DtN902ntHG6tjAwzotvESt5hi4vPPpltd+Bj1Z2PJeFKkAm
afkWHY33eSUXVDhMp+SPgd55Jiq2mKtEaXjX3354A3SmJUD9/FuhGWPa3wHmkRu0kXVLbNmBwE1C
R/XbBZLrXLMaRlmiYjd4rOVZMcTNCtsbdGEuQWX0HVtqKwJX1zJl9Yn8X3Z6XyBNZde1Fh56TzdM
VKKrAewyzsHsoasxP75UFfvgHYLRdu2OpEnqMAK36tBesFsYncXYxfCHvjuqSKtX7/AWrZi5sthu
8Wer/xz9PBOH4w8OFmWxQaPHJC4ZxZUKBASaswluBjl+wL292VC5Z7cEVutFve4n7qnRP5BkgOx0
MKm6QvqieH23ZProIojOjHrVJ1qFPbVdzeTixWreID/IVWAoU/XDzl9N2JeMMoKO2lxCVkEzceJ/
MxW8zG6O8rJB+Ho3g8Dj0Ha+Y2zMmlcVCl+oBE9gRk+HTFlnqKwiYiKGgnNXyXtjyOvlX7WoHamn
BRE/KeOCmk9KxT3+x0ySrOZZErk8TQNH9JwvJEJNNx4mVaRffiChQ0VpUVqeZ+7lcuaysUHnsDDW
XDkK9r5ajQoq38eVyspSPLQ4aCOd7bbAmf2jRhBxL01C6l+mbhS0pEb+HLD+bdTANIdt3bK8lfkt
TeqT1++46w6p4Fn8dkDL+suFQER5VPy0ldnKt8Uvk64o+spIVvB4oTMIr33VcbaRiYDBJ6S2Hdwu
n/gl/WB1Q6DA5E6dFkxeRmXKvwoVjkdvJxYL258K5C2FP0oyX+jNcNMwk/3KkSPJReVVsz0UmBAe
oATs+rbCdD1x5k3Hzf2zwAIZFiTYbN/PvpJLaeda6azzvHmDBOPnILDU+ByuH8ttRAldMEF5sgQA
OBa7JU5SCl1LMpPNfWTMEHvJwMTNkFMObzjfW6+viH04/mlV/3u8/8BnINvn+Y3sRKupApInxRri
ivkifkQgXfDlEmhGKH2we5qXcWghZ/Y+UhljmCMWnDHD/tpnvqgWbylMw6uKj4LcFJO8ltbTaCJS
eqjQBQ6Ox3LVSaeAX/TqtICJ83gCyoxre54tPf33qiV42tTW87XdYYcC1wz9OtlTghcfeAfMsg1u
oh3a08QYBHuL+6qwWrqtGn+PfmtDFYn84DV6libJWDzxWQVhEf6glAJ2KQEBviQHycaI6OS6auN8
BLKPPAfb02juBQRa7Sp9ZN+/LkUBM38UAt6V1RlJqe2ttHYvJ4gmgMttbksFiuYHVIElNJZtZVxJ
wiGrMVRJyjt+yTUQMyAqi1lTbtUZIWQ8lH38fcxexCOu9pv0dxeWslFIqKJVOURoIeTuck8jW+QP
x2Ej6wQYvqmCjMskEXgeiQipIycEM6gQ3r8K/kVJ+pHiR/d2ajjaHrysdfRjenrNNhgqknPeYmIE
QUSf8xztfTDqxecntXO+qRtymVmpEtT1Wyu9V/44xH+d0TlmkjIyzpzWWsKNWL5cAeGWBXKeHEtn
V65f0XXMv8mtQjUbAGTlaO3ZBDJMR10t5X++7Hac4H4nZ6nWNBa/697NOOSkbDLcIuGwTiLjU/xw
aWdLQLf0OTK78dydklUtiI5fkg008HjlDoYbEAX4ELw+fj3SmKVRbVdGm1id6kwG934M/cArjf0G
2fe4IUAQcJCZfH9wV0R0PBV8NfIn5u5mDtWaPCuEHoqSABiFHorEvZ65BdTtNDjw0Nb6mAeAhv9v
+Ib6oZ0v7hTmKoAkXBmffmWGzcAbcicsdtzzLtWjVCpEidiuKCZkw+rSHddu8ggH3V7Dg/ttVGZA
IEW78KozGiKNhTuY5lIda/YvBahLarR2hpsG2RQIectL5eCIyarv4aXTj2ZvmZ4XBQU6nKSK1kto
g+B8G6DUpDipo3nTCypnQXiN9uVmgg6NsCrQq98uRKG4bZIutP3a4CsrEKDkiJVytyKwurQc0WaX
ZqEVTtgsDpT4q9+QFL8iDL+jzhjnQo3iiPiZoAbxuJ4ACtXLrfB4ZIsuJ1zF4IEsMBLUGxdIl6HW
xaWupDA0SR5hP4FD5whL19hVvdjad2TKoLh9VfVVeiWiRFtBEACamPASqOvykWd+6rxvc35DMa14
xXZx4A7RnzQrKQJfdqAv6tFi0jtZ8fQdnH9XVzY0EayIP3XDHqeQx8AHOL/N2T4FJmsuV+z4YASU
mftdyoZV7qlvZ1rDvRFTAK0lYHTbhoAVJhbemM2VEKNROPWfn1o/vUvBsZ+pBmWcg3lrSWk5bvec
Bn+YARFcKWiHukGr1ClW8j8DKL+A17oA9BUU22FlJgrfJmajAiMeX9uThMJmAczxwQMADkNn/9Ke
gWXe6hWYKkx4jkkDiwdDwfX/xTlHa0o/IouAE0uv4vaV5IM+j6Kw9c8At4QVGdriw23b2U1r5m5k
NOZfcv+v27wdnrkA2AXU4jD4xFilsFbMtI7V4z0H8QT2FoURbBr/AWI/PbQFpyVwGE9bGdOmTf4Z
PJwH0L6XhO4czS03pZa2sP4MWM8QoVg7RuZCalPpMLhkmmuhI7SQU6iKmkZbcBxBg0XotlthHWPd
eenScetQ9eWATXlyfA9lUgpm/YEtUbcwbOtisE5miYnUc4yIyTZBSN55uPLWCKdfL6MZSX5ibYok
8r8q0lgfzgMVaN/lwQqcY+2BsS2YMDZ4jjUlaqGlx6ROfFI9brkHcq8fndaB8rnCGI6pdRDpK6VG
zSvhygsKcQGBvC7OpLhfNuHZXyC95PDChXLSwhWdfWn3d6/ZtP3bfOFYipRCg5q3MzeOSXLuSOZA
cHeHtSxdWy6fATzH2cXd6TTMbV2tAG+INcbAwTscc/AQ1eoAtgUoaOTABM6D0VfNg9nwKVQT/5BU
Do7AJcM7IHFEbpo2cfKpuyoKBTeri0fXwuRVn65+Gzzf1d8qruzw2vCVGdwffWZAGw1n/23VkXTS
C2DyzQK2MZyTtzcw2N+9a/OrXWQkxe4f/yFSodU/389q+oZbhSNsk5N/r2aW4V+z4qYtreqR7Asf
/oT3qlVmHd9v3DTmVeZA2sCGF8rFRgWDVGLMRgZq+BvA4ePO0lh05OpH/+GQ+IfxxNbIAft1amjr
048pi4Nkliou6mw8ysUg85f6WboPcgbGos3QRjrpQMSk6IMF7ov2B657k9yJtkr9D4yZAH/1AC73
dy8kS2a8BSSosqcTo6DFTo6cc3B3n3qojEq79E+uoqnLYL4gjeB4iU0wzr6XEFzyopVA+k9/MoOL
qIfFY0NZTeuPmAwhLlOuzV+79RVZp7aMmgNp/It9VnFY6CkwUoD8vKyOrAWMJAA243Ll95YUoc+s
UP6tbhrRjsf1rEr3gcNYOKxATlD+XbHUILqvctCiWqpE8DDNXBE0W7Wo3kxSzCl6h+j/0sUyK+pt
PnKkRgNKuWNtgk5IELx5lMZkFDNMrcrJAT0bd0ik4RreaFu08rpP/uJ1BFIJjyqq/qxyIrAj8Omx
VnbP0wIRYpHCAnQ+HNyuzSiCnEf5PxgDgfKM5YMZtmPuAf5JhbSLgil9FefZLOml3xQicZ5WkKEq
tCp/Y72mxaGww+ppULrDbsVZzL9ZOZUwdPcjRc7Tm5f2C+WXdCIrzN10dwE7Q3BeECpooC1qit1q
qCIIiWX6j09SP3PNjpsr1nvxKgbvr/TPjpiSSrKNNGale9hQmCyiOZt/K6y6hKnXk6l7BZ4wyc1v
FdcCkz/qwVfueZuRSaU2HRrPgfLQPL3CbfQGVOY5qpsKBm5rnnP5zhSo3afkI+0Qz4/cIGzINLhd
I+6652Kp2hSbXtQt8jExXzUiRxZ+YJ/lQbLZO4BWaXkZpRHHvw5/YcrcmPxUZFfy7kzOtEckVZfR
Ta/kTzk1jzNUWbya4wWAIO+zlvIejM/eJZ6yH1Sil51Zjsk4q/0YHoNn8cvsUicl+eCzsa/yY+Ba
A3PjvOjw4iCI0eGuEKOlp2NvcKMJTre8OX1QPlY9nE/Avhk7rgWOnP4vcYYtAmx5wV0i3xXd9gXH
mHWQrQTV8ZDPXgEyu85BtoyIid4j9yTw1F91FopcAG60VRBlQ+6rhPBehHX3j75KWClYHqjxtfzq
4krsWNU8dEgfSoPCAyhIzmiwflfBWC3rR4gi0rRTgld876k424Gl83o+J/yxXPJno2JIQhilEQdK
RMZv5v8tO04UzFgB6Gi8SUs8INpm9oAlDlRSiWsQJUNtIe9WB2Uhqda7lWCJU1MTfTy5FSysTB77
QiKZRzs6oEWNsftxsQj+UXD3Lgrc035ELE//oQ3Ozp0ybhtvowbth1onVccnreGbQ2TjuMIlWmhJ
4MaAMEI8rH9JvZaMiBySBDn3cDsPDCTYUMcBAa9L4NI/E0V06de4mq8Le0arlmY6tZjv345dsKFX
nF1E3GMvWQFenjz1jdq/F4E/BrKrOGqhhzpZnMTGAus9I95ZEUX3SlOt4CnxohdxZH3gtRdmF8Ku
hcmu1TnDPYCqDmHlkxI8YKCWCYiKfbgpDWnDWK1wQcFXOSd9Q37I9NvFovmVAJRANB/0oviuaKZQ
XDf15uwz8gAHikOHH8Vevxt/GZgicpLOyW3jkn3B6+wo1Fm7Bjsw58B46OETP1LKG1mANGfMBbaZ
n4wFoeuYxMY2XrG+gPjXND48dlPnl597uC4+ecfAMzL5Ycqq+bGALNocNd+qUdmdChGtZEJ4z/ek
XOwcttm6dV2autuDv8mLv74mMOILeAcoK7csucrdv1vpTQv0FwlMXstB0AU/oP09fBNiEvUMBRiu
lA0h8p9xJOc3LW8So+avnoUemp0k1sz3hY13bHIrQ7YEzdjCvUB7/xlr6Zg1nQ8D8K5aZ7Se7bo6
kHl3OFP58kgzq7jsTwigIyoFVSdm134INtfJTAq99cT/p7yBOaPXEe8m8oX+723jn6os5CTCfbXB
D690dLFPigeM+cx9klqzOms8FroQHKox1pwrzRJrSe02RCiajYe+WKsb05BFLrEgvQ2fOyKGscdt
4UrB5fEg7vKwPPXcVcq+h6kkHeq9NNSuLSqCIb1MutS1jrwlduXsY4ug+O1bEkWQgJyl5ym3iWY7
cJ2n1ANxORrS47tc3KvqNGPa8Yulz+qXN7FLgC7Zz+my78NlxXnAAlXx8cMSUjXg9LgJ+8NmCM38
Zzz88ylZuj/HsiM5F45OvcWPzHv+/TIgjIhS8cbHOh4LmYTQqRVZn8hx4q2Sx6HML4i7ZarpQpqK
+5QoQ5hfIEhCUjP/g1oLO2VATyh7ydKy+08ZK8KNXfw1Ysot4DENBi6ldrpmqyzry0e/+qxnPNXi
Oowbd0q1uw8wy+b4EPa9e1tu94lmXAi2vNiiwn+ObcX5hhcTNB73Z5kyX1lsDofWz+/P4bQKSE2L
dVZhHvvf40+JsXHtI4nY+3wQWq0aP/vAlsbx4SyUA85MkBsBgevglxB2tj7OvIXGODoSWsIe8Wr5
sXU9Iv5qmvaCcN3NHVrRUXoOgHDcme9sPLU188sGNpAeWwA2ELufJG6Sdy2PB1b1A1CmpplqvVia
wL5VGmdwmtwj8SjITo5b9q19VucZFSwBphkZwMfiGd5etdHqCb32ZP5nc5oOJdZtyUvkeR+b+s1o
b+P/436jSTmtlbev6/S7dx1+mHevb+XMjH6iYL4GiFSoeBE5o2hsHHcS8qzega9yjqYdB5HlOjqq
08ri3t9eBdXCVIyeVLkP73QJaFQ86tq5lir5FxBBMzWxyc62UwfkTShI4NphlXPJg7JeQNR6peYD
KT8GsVu9/sOwGhIIkUhrGWretkXydiJW4XwMY+vnSb5cVrMKYQk3vrvj+dHR3JRZW/nXuQueZjpq
GTgRxU4prL1HF7EeFTPCDoWojdkPQCCnAWkKU/svGYv0sf6l7w3b5Q0MMpJjrw8Tl4Mt76gMxA6u
qa7TJjXeWAdpWtL+zmgWsib+guIUME2UCcByq+fAHhlFplzYM2OfRgsGCw5r/y6DW+DZdqBRxXQI
O/X9CoDwtJkvvAPWmPpcglTy6CCpZ6xcGgn9i1Z8QWcdCcer0HaS9ADfd9wOGO2NmelO7JvKuCq1
ptPCa5TJV5gU9yBM+NYBilpNkTXpa3cXTIabTaxmGR5UJ6EWfUMlUk5dsW/3qhbFH1+nPVTQ3GBk
20txqWEpky9BTl3v+tGUuUQMRq5zEba6ogWEJT/4VdBCkw5nfgy/rLmznfoLjj+x7NfB2FKsWaV+
TNkPKZ7xUysmw55QWAUOdJRdN4rbtZx38lNZKUZnTEuV3mX+BOIfpb1kTUj00eJUJxhdVS/+e/uY
F0EnfdjdrlL09NUftX9N6M7z7GUtTdihkPWEzhM+HRsOraXlNFsL1uFaTxUnPwwBSZ7z5dd1SgsR
RGLyiw8UrnPrSDOGvmR2tlSFQNd+SJbzczkloA/KDuaBG0VdTlmWh+zLz1xkoGf06ObvpyYL6B8R
ucUyGK8Z92N7DuhsL/a4SNk0aoSPSxZfon+rxspXDuMIF64xai9Hm28iVtsy9Q1XDtlM4JqqfFLF
M6smTV+vn/xRUzAep1Kw2W1GKjdJ47UBIvUCkh9q8pldDINzt03TUDvjzTkjx+zF0XqqPUHZThRR
zV/XdTppDKabBdlx3WplEqtRE1f/yp0+qlMkq5CrusTbZ7nBjUsXYVdCvsUtfUFLWTBiclYEk3Vm
eXn8vxZguX3+RHSgg1BrTMss2hhABtgy55J4O4oIQa7atoNxQG1hPV77sNAV84u6i15hH/5+sL6j
I67JvNDtMLKL5tIUAOkIHfbG2epvs+P4rBhUbkuVJ51FRrKCBxWoXubU/cvvPYSKrbooHV32ydpU
+lX0N1nFYupgDeqj1d/XFJncP4mZMzF5h46bmjhVVraAPfg/ISycUE5DSx3kT1o2BIoZkjSWhNy+
H5ZQfzD4WyNbLgL1a+GHf8DCZCJwNUU3fm9Kri8e+USYeKmEBNwiB0NCcEd2+POPrQV1QrmzvTrB
rjfnHTTPugT8sCvhn69nPe9TEI/XUMbs4iMhbB8pN8tXHO94n5gQKXdL/3M9pQyZtyKPo8m4poDm
RDO5t5ncHSOlHyTc3gasQGGefAVxyWfADwXMfC/U7s4j124EdSFQFvgDhc2j6/XYqoWxmwAdLcv6
JrbASae45HuyIFvQZf+y7qfh6z2OWFQk/lPEljreXQ7Lbo0Uol+hXOt4ZuAX9zyyHzr8JIA6vCFl
nmezVAss6I5WlJe3AS9/BQYzaG0+9EG8n3LOnON7KaWFEO/OSmwqXps8x4vxpCfP4mFglbTXiRAW
O+OnBWwqkwnF2SMayTyrGPz6qqXfnCQQFyThM1snoJYh/wnxIV4lXPmQP3XjjVJp/OD/UdhSlmC9
aNatMjta2yNqYaullRsR9Sj3DFuSmFMVHlAg0ZdMXnX4evHDZsrZgOJ+gXKqjsNSasP0ux/PIdac
AXkXGF7NoZrrhdiucjPZrfUpHFS1Th0N5O2+R5AHxVxIGWwUiStg3fN2Jmx6+uhBFT9MyaYRoP7L
OfwqGAxX4IYv8HZ3XUQL4xojWjBj5nAksMbizWRdSd6CaDzsNc9gZA40SLULOOm4TqrTmm1EncUq
qmoY+nr9YxtC1bDKlxhQuua3Gqh7zTmwg1SuuLWc4sVxCIkIAYJ2CsQLCfZtPZko20VkOb+As0Xs
xcSA6qN4huBBAKJOeXmoP5iPqGo9PCfYKpGrtlpEGZQOVNJy7QFpZAD5IUEqW+6eGb78EzT90b1O
q72onrOojdDmJuh2Dg5Nm1Eld2iKLNxGGKAYAy36yOMOl1+cn3SKpxCj8IUDqqbzgafVkhE8raoa
XIV2Rv+lpjQq85P/CWjQ+9ik/FyoZQz4dLBjmXAp1Mg4BWgyrxBxb6pXcJ8khe4pBH0w55W76AB/
dVmmAPGpM5c8jVO/ajrRJTHG0CA4cHpgQxNXQOmvInxgVqv3mDZD4tqr9jtDC1aIf/Lsw15sP+FT
X47CfR+u7jO10h7Ts+kh7oH/4dgQQwPoSpx7Tb2kAQcdX+Lf/l7EampPQkf5sF+77odh6+YkA/Tz
7HCpTO13oALvj68RYljDME+D9LGW8zB7UwpD1Sy23/S1xBtCMdnXtczVAN/9BURYzcmscjPx2qOv
iyFLaciu+/F8jGn8WB7+cgXARe2LrIgaPHgs6TPvsNZOcd2tE28lGYHoN6cFMoSz3mGp8cGrE/SJ
2PpVcLHVHXtMxmhm/iUCRxN1GhLCW0z+W+F+ria5escSFyUxD6ViOsfrZDYSc8V1TtpNy8CHxory
g2SeL509REY+sBE9iOnfQ8jc+onUY2Mzo1cHvJDYTZGx9tYZ1L9q5SWgsb0PUEe4ey0bk3Fd/xjJ
vRk4cQT7sB8WIDf9vpwBWgCGL6eATIbSDLgtYmfp8FHcRg9GFIYjXigZ1kNwIgqRKZ4X6cndTfKE
YYjN0M9WjhL03VjV1eGvufitcHsnuCe57RkKBvz4Xq0N67h8WjNcVsuFDFZyaoXmFo5i00pN/yay
B7afWdubxQKr/L6Y2tRco3y8jpHw2GjECLXZdg/tAItvNyruiR+KM9jcZe/KLrfBFUOy4vd+0XP2
gQ73nt6Su1x0TEvQ8tNvgwcH6AHHTfLBRUQsigfRTuFP2V1Lb5A6mgZYwbdG2Cff6Qv7RrgIlFQZ
YMGoVhRNbYkkQ/tOYlV5Lt4CQbaJSc5C6VNTUynGlxV2BemsI20Ki/UBkzWsYRHTV3VjkJHw9GyB
UqhSbMz74ISvL3bE38JnotCYCz+vUvyXTHcyWd8Ykiumz3Uti66oAy6ovs2JK8XC0H8+jr7KvzaB
K6TNprxAroM756dCNhKDI6lwYkoS5hFAw+DzUWXpY6ZC/SnS3GAq82u8JsKM68ajaZwn+rXSVEzh
6+q2s+/OicFqXSsKenb77amsXjHT3ZEciGX079oDVAfNbipFFhsG832InnAP1fiGzmNfOfDFCxew
rPrukgdPx8SHx9upfmZa2exUxIrhaAtHAq3dzjMmnPUPrsp7t5yDgySyT22mqgz54UY9aWQas2XD
oIfpy+bLETrnIJLkRnKlTf8Gs6x3BsV3psZN3C1fA0Qq7kSw/Itj0FoaeGsrKobA/gbY9th7kqKi
uU3VBM2YkBAH4Tb8dkYwwMYkZg0LffpNjGI9z5Vxl2HqHrDhdeHAEdxA7bX5GciLuMURAaQKVZwR
fZiUwBKUyO5jZsnIyO8TZOHcEr5MhclWfdiPJNAaaJnehanDrP/Jzbi85jlvYyX/lsfz4CBLcUzy
5j1xQHp0pfv1U1dR4WMUexaoMEIwz2z8P0hjv0rg2BXrlGECI7yD6RA3QKgS4MMUQLouFdEx0YU+
KTIL4UlzmZ2xmj6na+5Zk4gKHrF+3O0RMweksVo1VP9xI43/IQPDvKmd5uyXVdRg+j41dYqpAUl3
odCLmsZyxx8iG92S8AgjRzHuMPTq5dlu1r86OFzpzfPmeBSNgtlrlxfHw+8+EWeWqCi02ZGa6jfN
CZluDU8BJjHdCV2udzW6Itwq8Aa/jqax50uTGifLXs07WFazwzkpJTtlvT8Jlpw3VZvY+0cGqBJB
qPImHOgGS/E+g/XkAe/J7JsnFddN7i7ds3Ea6YkWe2ei7AJgSiFMwLby+S+zA1/OFcCj0GcOBx5/
vCZXgXbZmWCrcnBeOuXuxhsGL7+fZR8WZ5T+pyhifUuBnmijTCY2vZdiD9LMr/Qz2CntL+cN/rSo
2Re8ARAjHgpCxpdAIQhpXnlzS3/HE6+rngTbVl1mySVWa3e4EGLmu1AU2hYIUNmaYfA56bl8LH7Y
KxO4nnfA3fAIKuXMHXNClYUzhZjpiykO+350VzStjAijNb8gFQh71D9cSzbzC1qn4bYDQyx06TGO
R59CJ2vmYZ3NtcG5AHmSuQeLGB2mREvOeNMhCiD2ws2B5vxTM8hgdDKFuFmLLbdcu0Z6D1gNKqxW
CUxF2xYSG/fop3HlG4U4qDqPalo4jchdEoWpAzZrarVsrMAex8DpNuYut0Jg1tt6KKGvCsaCxAJ1
YdScElsLmuUuE7G7FB7Zp4phZV6ySoW6sHUZarJ0bRQwcQhgge143elEHQFm2hG5bDhFrNV2uzO6
aSzUKIt/XiAxlG9p4BRFxKIKqQV7w0cEdQyYWYHrRJ2t4eHEJPY33YB5JLc1m6aEUD3vpLEIgZfq
7CwK4Ze5Ab7yxnxw+nj8GRyD6xfLOKQQpaHhxTvNxemW2wAKvOko1aGO/B3ewaSyv9wqvOVgImEo
B0AQ/BQ4z/nsLR1ZV+AvueA3kH0xpq9diFI/xJFZCHemYQJPeoQfPLpzfSRKfwzYqde4VWLn6yiI
A2S/0Q/9khW363nC5LJ8VCvs1F3mOv9Xldi0AjFtZKdGpKW/KQteOhbi/rk6JYCNBZaRG7yesNAK
kUyvAsk6fg/Q/x/f2nKV46KFbktYTdIg8fFH23/H9GGXOyBYJtEFBFhcDzzaNAJENSyihulNYrsC
4PGMU50DRJujWpc+pK5lJY/xw2sJWBli7m8WthhiM9/FeFYxthDZqA+DTyU5XtvhOGdR+rkbklv+
9+Ji7CqZHaA8bb9oU7A2O9nHQ26hFLpZPa2vQi4EQVl6eXgNqZhd1oQUdC4yzZywK9zWhsQmPTSh
oSKgdAJR3mwAfj+jj8LgjauFL3MYavhgv6lk0PwBf3RjmSRsS5pU1SxLTJ1ING/o62wN+/SDDDMl
5iTd+kPlb3XdiRNuTcwK48ftEZidAesJYRd8qiCv+vNVEYD+PY1TzTFhQ/MdEdA3wbDs/L+uSdex
QIpSodirdWdGwS8UyLjOxMnxsT+Lws4fbANtNI6Hh7gxjiY6NyhEKYM4Z6s7XdCa7m+4MHD3tuR0
L8oNGoJet3SF8dvsAy8Kbs7w2Td1BD3/sluaktR2tLe1nd779GtKGsPLRPmYjMPKlOVBG9gBobVm
VL4Hb8XsX6Z0LfczbWFvJjbfjpD0IqadNaEWNxlCWPQViIS5+aUFNzRjwAWGPCB7w6SVuNGzrdQR
wjmmk7Xz2mxzplQD/Yyroj3APjPrM0oagTfm61Jn8t2p4aRZmoBBxSJfslnPmD1mKMPK8Pa2ejY4
xjTbCZoP2Fr+t+/7PiX+/eJHlebLIEJtD+MiA+EmXoh0Rb5c3R/rNFLJWVdWWqtdT2EEBrpU5AI0
+lukUPNVSgsjtwKC/SvSMmxvfe89ooBVFNudO6P+xyouS60jm04HOdGj9BVK6bQOMHMelxRfnOsi
PsSu9jIbaw5SKsP2cHAuDBcFA3kliMGlJ+gdXS0oIZD0atSEX/dZgIn8LID5fzY9jkRNt3iQ1Fg1
Ujoj95B+0wtNScKnjx+b5X/TcckwMnrGvdKBRMPk5r1FUP0m1Xgqsq450uCJNxWBeJhH4+u88vzd
sYPCtPcZFt3ojZd+mbsecCWHwAn5iSYWDtuMGYtM3jZbhLAxU6uPI7Htc/EsEdkLaXVtL1mjl8wE
NcmYK+CJ6531DBJnwKCmqjEPA+ievS4DxjXn4e0yDLVqx35AbfAxgDXds6cAW5iIQh2xdQOpiTFM
0IdxsRHvgVJAdumphb115ucqWD33G2uH27xL/LJp7JtRD4QB7amq5Nkk3g7/hRh0dZMBxAdS8Xpq
iMpYfXZQDUHlpzVK5nCdOZ6AKrF2oQlBCL7JGEAGpimGgAn5PvRWYGfvvyE7gIK9ow2yjkpTXLhk
3cmz8KC0bdSlqSxP6EDyMEU4ePUsIPG5qAnnJVXSErvhAn9y/FfC5CYz8ttrQ9U21X+Kwq/GMjB8
kEBgVROaARQP81Fmkvd3CAYCjMr4GOZgm+ey2jvvpQAm9uSMKDhuMZ0PHP12F5zRF+dWov7/gf3K
ynwqFO9ksTvXb7fcWfOpv2wuGUf0v035X/ASmjCY6B16nG/lbFihXVXZcHdqjpPxYHl4bs8kB9Gr
0ZhXdLG6Auk1C1DDCLnu/U1OSYBWk8Otv8QxMlLdBONsA0IBGER69RoI4PUBOacnGDqwJEZoFP1y
zrS4GXdTb3ju+Sr2eVhD49i3xZo6w3Oe78R5a3wOXpgw9ykVkIahJwwl25i0WceZvitYEYGWETn8
9b26eHowVopf1oPKISg2OX+q0V3mrJ30SSGwhBPpyk6M2KvVd7oVwGXoGvX9oU5gonQ4Q539GJhi
yRhQdOS17kHCeKSlIcmSSHzzOML8Svx0wiUbLSTRogDckYWiVPtAQCQJp7y1kf5asM1SIDVRWJXK
rEjagTyZaWhKJ46MvX4AISmb7bTHFEpm6BZMfjZHvtPYl4Fb1Wl4XtjeSmIrGlzFT1zaJ2XoSLkW
s9IMpbcVgFdNeKFIcwHAK2KmY+HLYzOpoH02UjgOzeH4uHBXE491pPUw6Pw4IUtCkJyr9ZuGBPLi
KnErwV5QjSl5k6Y/k0hDbz/A/M5OkwBtLfZLrJNzl9OP9dz7PBBoN/IfNHxU0dUu2XEv8/ne5NRE
X9/oYP/dG0C3qhi3kjDkIq2+QDt+Ut0if9h6ArpNeRql99bkgjJf3Hfh/68kRiBjMEQ72E7k67y3
Lg+lhhCwhKcOekYRWl/km37rNtlWylVcwtiQlS28YX3KWSTwai7dizV/KsyysW7HwERORdUH384M
/8+c8LrV3jcuMso36ms8tCt8+E3K7WsJaM0DbfI83HAgoiOKsJAm9VMI1xCW6XwjN9vBKiKbcYRK
JoZIF4CA2I2fsqlAjv9ToAlSjehK2GQUX78PEHj4/lh03CdegfEfSS5pXDOcbNV/HKTeTJong2sx
DoslbYJIs/QqcZJ2jkV3Ifp0oMHBtLPH4LZhD7GQw2JDM9+zieETQ6w9orXV7xLH2ATRHeqsucXS
fdsH2BYJbk+bYkS/yI1wDjM+CBtHcyf569atOGOXFLI4n5oMd5Rm1iV9jwk5TIDrYZ6zNsiE2Hzg
0atkkOPRDm8wKaFORgm41YQ0vS+DYviRG5WGYUBZ67sqfZGoJMnmgAsQ8TKdEIw/VZFw4W5PFyy9
rKVCMwRIz8/pmXRqPBeAsCohc2jLTK1u+MXr2eQCd/shrim4U8inPs6o0rCN5d4aw50xbFRSYC/W
EWXJS4QmYaWYSvudDCOMji7B3rSIpyVQpYNdizG3y9Q9njEHe6L3rJGiZHo4VvJMbSq+QeONS/xN
2UNGCEHywteotApCbFtSx4RFvpyI9NafQR/G+h8FX0Zn26L0fz6kXyUFwB0Lz2XOwvv+FExHgjUj
CloM7m1rpyDYmx6yMYCcaIMVAt6U9SGs5arzMfhSDQ1uVkRwu0QozI/AjFt4fT8nAU3wS6LuhVrI
McOw3fH53CeV3xVbpUBuSfXwqLAzgfU0xsUWeMI2Eark2FpoLfQ75IFeRijbiOG/1ORfEWSy8iLC
VQQuMFDPNvRUGcoIsJkI2ciqaByudnx1QFqZq+eBc/jSqMqJuagEfCMkS0BM9zqJ89v6QJpPsJhJ
ubeJ47Mfv6/4YTwVQmhLx56dZeY/CxZFPWKxGfc3ARrm2osBqv9PvsybRUdLpMYq3BtPn/it2dUd
4RKwYKbD1jpcMS+RB45NhblqS1AzLPucRmbwl2/ly/oQTFB+Slth2MczIz/rNMZtY0djEelWwsuj
894H0ZPwWygAsTzbf0Qw0yyBNCZDKPvePQ9kjJL15P5SLs8KDeD64azCnsE3sIIr72wM8JOYxBxF
4nYn1CVFUE2iI1nF5RAN4xDfecK+/eKLFKpturpHL3kMQDwu+m8tyUXqZ5co7Gve4kKZOLn8jPCJ
aRcRuFzKyCSg7TGCiJEXhcg1yhPc+rodFv3Q6vG9kkM7GndfEzeaRyoXrzN0IiQ8CakkOHjQVJSF
3IIdfy6j3vXJmrpE1ZHe2Qt/ZWZ2i5qu04ARnS2I142yP2OQ0m39Fy9hqA0V6kLqV8b7JYfA8/kq
dH18Ixjfaz60J205BSeomIwrrDIwxEM5lpJPr6FFz8rlgnBPXB19wbbi5G4bBVbDKHVJSVGvkYse
yFI89cVjjNZzHAaW3lNdmtmOJ9NHSmccLjLMNOU8r3whh1mw5e6W3FjtB1/+yoh48SGfRBcERrCI
dOUKpUt/J/EMQYBFDnYJZKrK2XIitl7z2uUDTYOuagaoAl8qj7Ok+ZLsvWOh/CmBjk/3SyEqAILx
kyIs7hcy7RO8to/l32Yg/2iJkGlD69DHehRIv/BLlrd3c3lriCEsUma93KkQZdJQlTyX15gSN4TF
gGJaaBr88J3hFYdGKi6eKmVo+pGqgA8uzJyNiI+FdyDWNUQidp1jpDE4l3sJREy2IXx+Wvw/4Qmy
2ieObf7eLdQMbSRWj3cLN5N9tleJzlmwLkOHMMw1/Bn159r7R9kiv+vElz1rYBr62vJ45JXs6MhA
EAWYzifRpIO1hGwPW+tOBOKknIz7jVnN906wNQheavk/l3ifQkIPgrqfMrQ5YVx+8hMQolC8RSZ8
2+d0hq4VIFic1IheWGUL1J/7Cg9vid4QqnhlNoKsmcPbQqZ5h1MTke2Yn59sHyP4seHkL5EXBQCY
BDpVQeQmNFKwnVxMPsDl0GmOM7P9FpLJMKdn6j6uqvVgDnDTX1yovxzEl/M4UalNflsI8A0Cp6Qx
OYoWTqAI+nIGg+xWUNGjl2FazKjMECzs3FzhrI+bxlz2j1nfqBw/YRVBCivshcorB3yp2URgNBS0
+DydT8NXzxB5ZTeHGPbXS+ZEyuhvwS1e79ZRry5kAwG6RPUM38AN47+zIiB/ejTBJ4s+z8utb0Xi
XmILICYa+X9bGhDFwVKIutA03J4aQb9hcV63efJAa+G4/D/AXjeHcCKfi1IMVleAwbODznXcPsgn
dZJtF6ghtUp54AMtXbMNdgbys6i56EI6p+Cx+1MWwaYKrzQrJsp0HtEvZ2cglt36wIsBGHOs4+/o
mzxDB/dIU2U7J5BZEbQeq8hLDg2J0WEtWMlBAxvFVtUeo+FffCHS3V3bGt/jqIBB1Vff3+MhQAL1
Hxg0WOu92HpiAxHVz0/12jkj84foLcQCG369y1bVkk86Sh6HYi5wE8bl9MbmiDJYQpixjvbk/kTv
EQRssDyPByDaF+VHWFFQ9zY4sUsxkcU9lzxGL5cD1iF0iRoEmPLkUycMPia+kuzx/weMaopv6QWr
KobuIrLNZDdl8ytNtzf2n+Co8i0NatgG2VtfMi6OlgA2F7Qao8mZ3TIroZmCtN2SxwY9Q6eU9HBT
2+QsNemn1Tx//U1LPDEmb6Qi4rul2xJ0WoLwKKFfen1HyXsapmocPYSKG1qJIMD5qdw/1cX13/RO
4tEUjPnAy6PjreylLbuVB5YSq40MOaFlyH40H7DRxZBVw3mNtZgud33IhHljR3f3KxdieLoBNFHm
wtLyJa2JnqJKHfJxGrQz6OH6GNNfGoBG0zpjUAUteNZ5saSKjGyxjt7Yv6IK511drut4FgwSH/8j
gcnJEK3EX9l8QfDJSo3aTE6GJQ18XEXjiI0UtEXz9zxmIu5mJFF7+if8BrLWHZ/3/yCGtAn1lqYa
Jzu1hqqfFJ2SqVGQK8r1LbzkZUkfByxsoD5f0MR0DEeKx504v9wjMrflHj0qI3iCD6kM+jQm964h
igZnNTR5OXcSjXDiZyiltY0V0go41sxQgmCK/bZrMHj6h2vAF3S0yBlIw4VXM7KVT57s/K6avAdx
mOGPP5V0Vcu1JcyQ6+i7spwYwIW49CJvU1Amy7q2CWaSgm5mAaa9I0Nvh4p/xjSHP1DfCS1boRLl
Jayw8MdWc2cW+LlCmc7mPVw1X8kUXTblsT2PmX5+9fsDs9mpPX86hyPVLWhvZJMYsNOEwmkBtbhj
IztEIjPMgW1qaqL1PzWK4w0LSeZOXI+MiTjD6b2EXYIFHHWgNOc+9lEigEXKIFA2ge/h9fIjlMP3
8DauWl15z2uFFa/SkyH8aqZc2hIDtzHlnxrxr+lG8++Tvttbffr3vBDM+CbtlQNYApPAPLrcSpC6
CHqOvRsb4gYDlr2Sc5OGPAS439m6T/Z1HcwXmYnOHirSud5DVvNGKlQBOnfFfXqxBMvpGvOl+yhV
hVdfcVPKQnAUwv0LsKhU629z4UrzPNiJHO7yD26hnyV8ANZMgeKjVBb9e++MOLUxDxTciL9Qps5P
hDEsL82h1vCr/43fVle9JInwvlzjYW8B+R+eugYGK5BtnIJlFlFTMsC4Qibflf4V9rBM7zL3RUqV
XKzTG4iG10O8vr8AQpNzyei9IfEA50iudx6g/XJQ2FoqzTxQg3CPd3z+3UyxolvSWq3dnY+L8XSV
kSFBbSswn5INhvTmOn8dSVYZvb3RUq/jTTjPLtTZieS+t3xM3gMS+UplkJulstLc7sMpAjfzVhoW
mZaO7obrBEhIIgym+kXDsaupfCbuBSkSY+1/REPzeuAFnpiwjyHSrvE3WZnYQ9MwlFiuvpDHfEwN
yVjWkKzwKt98d69oZ9KeU81CyepQFgw8gju2Ur4DRBmEI7tarZSwbjpVKEizgi3CjXl2y1/a1q5r
YYrnCS3IPiWjGaYm6HdWykDTpGKgrxB9VzNxXXr1M7cMgzkoVuttsO9MReGHaufkt4OLAjBi63b1
l5590SRRmEBN753iCVRKx/BqyOakJT1P8HZnQoQVUljOTRrdjJQDF3avE2VdnYhl6aMxLt/a5v7c
kLSd3I1tW3FMf3erySRVrS2l8Ry0CnXFApYFYk0gqweLTYKwXTXzWfPJRY75N3L1GCmfJDkqYyEc
Y4bAjN8dcUsGFXcHXnaP7XkBsZIn4a8Qdrd7IXiMy4JJ2A07h2oh5hvLZqPxdkioz3t/Ydp4x4Dp
Lx9PwymRGCU4JR6M0xXCEPJwFTIEYRqe64TKjhdLxvyFlY4lNeWhxu6bi7UJhQYeKHbwzi3gh6vS
iSHbvslJxoVSp0oYhceT5B5u5GVZDVZMMrHuwJ+82DtQuhJqX9LzWUcC7RjD8fKUsAJpzAJRl1xD
NIH6wPnN4QFNSeoDQWAzYM6yQfK3S0G5fg4LqgmwWFu5KEL78rxYzn8mjH4R/sK/YVaccC9naYtK
szbDWLqW7XD+uxNiaJ/t0S7xs1YQ7wUZcHR4eVL6+S9zCtF/YBygOTsNIBVQW6ZaTOks4EGGi+w9
hKo8PWCUqm+GmZFjh9IjOE8DQBRZyz6dQYZupa0ye9WgXTpVW0mxZzK1+4oDRZemQnKdxQzeY3zN
dEmr9KPpkGfUdGGFBzUVPWCIZunjiS8vBXFRd4CHPWUn2iAJYyd0Z1g0ura6JKtofyLqXSZ99PqE
YF5mvvNn5cLdzHvBw8qjKf5NnvImlvaqWSZscHQbTt2ZgcOagF8G5Pv/M9X8+GlA+OsuR9ZILQUV
okXnHutvEIRAlUGkC114AMsfj2AKpWKlfST5Wu8lhvWGrh5S5Im8uf7a+QEEAdudB58qm86KAx+p
EHgII2oy/qdktiWiezHVPbiD+UKg0KirfZKVyoBVon2WYeaouffZb0WzwXZKKGmSAQV+MB2nu6/q
Pj4zF/5A1/RCLkgaWG13/6VQ+g5ntNwjpYlob4bZx2lSKNhHCfBF+wA1cSR8f4LjaAnYONiB55k5
oUrYrSLXTBcGWNnsU/dgV4fvyuPQy/9qa9nvZlcVgbix8uBAFV/eLbLBTukNzXNGLit3Ul8EmVVB
EpSNRAi2LWCCDGBkfKRUWfosbJUW5wiAgWgoFrcMu16gcKO3ufCg10L0jh4ijTXZ4M8s9EXYroEz
yOsb2H0gsrSmUEBX4ePuXybFaaqG8+5+gQJEuhAr0aOI5uDkLsilawtEHpioKvrFDJTs6SfmP3ST
bdPPAnI67SBArIDtaTzzYyL5PJLfxq2NdZaNs8cVvnisDbyTYvbsjtTenz4fjxJFcYtZYgc6byI3
CEL1y1DU3nKfngPYgFiYDzKTduDgN1kWG9dZAKJW+gc49Kw+YYrOvRQ8JNHwk3npweNfvDj6e7FH
bEoYQ2ve1e2S4Uc9yvP7QeKFm1PYhA6/8By/GPsfcZP4NrQUECXhdavjrpSRKRTaAJWnsPLatN8l
7pzWoraoP/5E4aDSJ4v6JgHEiLU71yivePu06X6y1W26zv3SbqbK/oGKuEv/i24HVt8iVPG53Ifg
XWOo6HAHSrfDtTvAiWLSc95Gvaj0p63U4dSafYJdCi7SxkprXdQfrWam/nSqBjpdBUDF4soIxwfi
VRVfDT60O31Fg693beU8EoMbwr1HV/56lQ17ru4UotK+4wkWSUEkwXCMWHvGPEftQe+OD2EET9ml
rvF9VmhraolVsXEo7wfhLsm4c2H5uJ8RnKAuloIi7FLgVPK69EO/D0XuEtNmf6NmqChbIDFBbLL7
wpucR/xkF3tz0WwoiOosHOwrHJUaLutOa+WuKHOvojvZzM3XVpcvVJwQOth8ohp7ITe2a8vbYIeT
NwAyv+QIzVpfDKWG9DcetuaRariZmIi6WZffWnevnO2NWxNOgQw9zGVNO4YMQ6pi98Xc/ae4L+Jv
Ah43NZvubXFrifdZTjS2punEbKozVKC6qQx1iI7pyRycRBQfKxIRw6sdUwX/eIGc4fwk4Ao2Oydj
FMZfU6gSc/RQUbZ848q2vkPiV0I2npF3rY+vJsoFwZXZyG0YYL/y0pBb/PVk2x0Pbs52yzozmrX4
aeO3tMtIbUGgAVTLgizRatKFml3d9nSadgp4yCZVZnD2ept67VRDlZ8YxUQxV2uX3iyv852Usz0J
jShCSBSf4vMQFG2xA3kQFyOD4ruFzQnBjNc4Dn/mY9UPij/1DZbzeE7vGtT+WqtclYm0kqp1TBKO
Up1Z6kGWmPzT8EuDXwhounLx77THHOxB+eC4nhrx0BsZD7MJdMKhIKxsQ0Oxs4Ahjgco3Mju43YW
hwODzfaeplVleaTX/yVh70f4jVchv18WBZOPhhlBAs3s3YOjg4ctpggTrNYGMA7J1bB1sj+mEf6o
30k2eASvEKPYLPoNzUuVvPxaXXndMPN1xrCujPr8CSxTf2J45pkYEiQuonO3sDEltu2VnmwR21g9
3ThtvxyLp1YXEu8cNpmzfbILe8ZphvYLvEI8R1P0FPmTETXX/6+f1AuPLcQxEyioysQx/tzN3Zwz
+vxDRdyvHaX7RKf5suEdTscqrDxaPpnXqwqZzwXdLqgnR4LItfraYfU2yJLi1W6VVpm3GrNIHG14
5VinWbyqjVhwAW8V9WzlW8Zi4MvLpnHE78R3SLjoFoeDzl12itOhifYoBZBDhrfiRDFZV1gP1Exp
LuNmM4544zoMKJWDCfTvPTxC9TYmiLlQGJgdXxxNXH8TEsTXuYgjwX50TS7Q/saCHYSCe7LYf//I
9tUEckHd7CL4NGk76a7YKCIPJeN2wxWrFgbHOrfA3jb1bfr+4qbR1psNwC0sIZiQlXba1ELJO6Fb
o1uzFEsAe+XW8U6k4aACmJEqLpMDMVo+KShtdWI53n7/Hb/FLYE2OujSyotvQfCGcSEnUrg96wWk
7brD5wEsxiUhVC5LR1J+YQ+E+GrWcj2ap0/J4AmyLO9v6o/oMxKODVOynXhuutL70AUGsaJGmWic
xXfxWWOSdOaIUMNJo1NtzMXwcWzFhdQsfzMCCUITDvL+yQzX0UcdHbYqO20gBM+pP+Cy1PN9t2yu
wONZbmeL9eApVfcNvauSq6fVzVOhONa6hyf8/2ywbe1ANe57QZ1yE+ALCNGDQQtsw4U4UxK37qNC
BJ/Kv1Fj2QWdwT3br0PZW+2bKraDUTzv1L8b1rm2JeKzJTpRNOCwF5EU+zs5XN4W4DKgBqpR8aS/
J9lNzxoK4MMf+rYiQtOS/pi3QBC27lpLUNOUwyG/pd8xs8LUSvH5hMNi6ze39cpRkx1joUILrxLR
cwBcYWUKCMpmbqGgDhEtLHee5hTgwEaTks6oj46eLzf+a76MMmMfLJYwLyu7hC+849/j7BljxCWA
Byb6bZ5qDFQs1F+a7FnUN32+3fiqmNiT+IEAF7mqZpywY8+w24uwYvTLZv+gVo8ZBVbgWcM/QAKp
bEwERucKh4I8oLlSCEwgHuAt36ePgI+pGflZUlYg7jjCJncS44uevBa723N7ekt1QQVEuUTT9S0e
5semJs2MHR+YwYm5h11FoDl1mLlhx4hquasSUY7JpBebjRXdb2CcWwMKGJoBvzGCmWUhbq/R8i3O
bb1xPb0UQ6QjsEqqgKB9iz/j3geYx8FzRzm1uAd5W5j03+1G4J5cDVsH9yaQt29sswgwhMeNFnrs
b+1KS4oWKtJhnaxpjqFcBAkHH/ALP8x6CzKxlbqDBDXMG5pNatfLHso9JQjr7NICo/LTa+aewWTI
HXspbKbqNxnvL2SzUxhXx8iHJYV4M83nWZCpz9Mfx5rGZSWw5O5XATNu59W7Rjiefo2HKxO1BiZU
1ryH0khdbODhZ4vVfQL3TMDmGbPDhd82nc91/hZySdKgY42k5owlx+ymy6eDZVtD1kK4WR/QHHqe
5aQw98+Po3c2A48dXqixuUTQz8PkuII7KSd2pi7KFBHWdmZruA1tx5gR7qucmtnKmJtCam4xWWfL
jq/dNCSUMwskueLp7CcFNk7v6uefJ8zaisNRKT0jJCEJ8jjUWt7vgAWo16xgYEmWQwZo0BIS4hUO
AvVdYH+3lSR+Iy7tPUIVl5eo40kX+W9PnYIUrYHlbBVZSFWGQGIJKK5uyByYnxTfa0KANJNZ9Q/7
2UFA7WIgiq6zRGliSXQBJ+bbcHwu55QRPolrivQ/cLtSnwILE3X2qYjZXEcrALHOigRxwZtc2JuN
m2E56lM82qvReIu4vmsBCO/Iqcr5yj9cDL0HFA4jovOMGQY6fTAq/GS/rxQzAgHdk4/CbmPTQzzV
D+aE+TSZsioTOlGLQLo82X23FP82GkdyggUSOA9e9m9ehBkwEQ9iFVRka+Alzfwm1GpYV4hi/lA+
7xEO7bJjB9j5dIFTBP0pfSk1NdbNb1/3637qoVCYH/Lo8JiGt9bKwCd7p8tEgaFzueFqT6v6H3Dm
MtWQQLgr7k92A+gD446bdy/xNXy7iBXvXck/SHhkumgpRZrbGlraGcjUsoWsaAXMkj/huEqzgdTx
Yb8l512L4VSrShrAfRSu/9i/GYylGafjwmZz+71rQS1Xc1kvsaXy5uQL+zkXDZ849KxUJCaPlE5A
XuW/TFsgKkaxDY666ErzLG88s1G3LJDYhvletRhSkLUbRanmlWO24jq9o0ORmpKU2rglECeSVudf
/wYNMnp3kfHvJwyNxAJWk7KpagSa4pravAwyUwy4usz8B0elqaeTcSKu1MTThjqKl3hvRURKc0FF
KHGlaNJfl/6BSqOS7lJT95l/PAU1qt+H/LnrzcFA+hYGZk/vzQl6GAZ16Ppay+IuJ7FmQ/VjMYFO
m1cA71e7N4as0jxiB+r4O5qFEkBuOkx/TkRLYNj/ohSCuGBWE4BaxC/HRLAtqNXuJy+RcpRR8/RJ
E2zRcvvoR/b6GIN6S0PUdmeW1wRYvuThgngIBJxlxW/JqyyPVX85/5IRolVrt0xx6sK/XVqlDRm0
ur34b16pkQFkrb6aCdO3X1KJJ1S6cliwnGkjc+2PeN0HX4tEvEE1a0auPxm9nOZxrh3DPEfynkn3
dyrjw56mYNQjmLuRfwMDCFFDcjNV/+DXXGLsxoQWk9xRK3XBAEf4tWzusIhqlO3YpPsxYGL5Dw7a
L32FVFGDwMQ2bFRgQuZXCJnqhgb93rc75vCN4aUjHQJHCPrwWnQe++k61iNhoNUbNNbmx6+6Cwlj
/qOWGTU/rZlFE9p5zrYXgcXvWcyipgsDyO0WW5wnCbUjDuumrhjj2yxpTETdXxSzzym4xjMQLxM4
cmOAxwX2rBqfdkBSpOHOWevCwzsiInyaBAVyVeTVeeDOIflnk0Ydtn3NfxuemPXfCZ8HMsUsMIas
eDP6XNPm4sKntskrLbxbqgJ9w/B1c2cgclbYg2xfnr8oFxE6MZ55MmIPCRuqfJEjiwD8HNCZyxxv
VGoSKwqgi9p6yqdl6Lyb8SskvrAqD0kZ6G2UGfLrLGP+2J6QTdLtbAZdPFEBBLl91O+rPggNjiuf
hezUK+tbmtjsUH51eytG6VeXAJq3Ha87pNdvCAPgwjm/NZv/8yLLHLpHb9NPjdxPx6c1TV7lnr+c
NI7g8ftGP6NgXiP0YIOQIUhOpVKvfvBC14WhLCnWJ/HCLefPlHVRisGEYHQNsaQ9kQrPl2JQfzFp
3XCH3fsZgbAdoc+NOSmU5OBIEMP2slZiJvKHCn5elk6spMw/QvEzetFcQZVo30NG+12Jru672t9l
9bkX6klm28Bb+UQHWJKa4M+NHuEVEJdfbeaKhW4+YhM7S0BHlK+XvTjK7l1uouDVaOG74bleuE9K
5TAlj80RQaTZFDiv0F1hbrKAdvOdDVLDi36w84WMzQ7r0Em/+dakxe72fLRcd8h8WIwwMNLtgj2E
BKtuzhr1uoHPtw5fbC9LeNJGNRsRA5nWnINeCrn6sN7U5E/brUswWBQ+0PWI8VRCzGeNj3wdA0Kj
4gBf/032YOK5zuePdalUN6zNraF0g9E4J9lFa7dyyLifp6C2wwLUmwqJ/lLF9nw5gx8COMWD8F+g
73YBvfruo9pILZcD4qD3Wov3vGFjd34ob6zKLRO0PU+4+4FgVp1Jcs3z1xV3vURumsiB7/Fe3TPc
G1aYWO6W14AIYpoPdycwV6aMuVwEbeB75ET7bhNKoKl7vhj9I+HHavraBVFx4QhkZlQL9+4YhtuW
Z7xcJMK61aXXmXkxKPgd3xEaZvh4Daku5lG8d34yS8l9+gspILMmsurweXeZDGNs9RJCmltc7Mol
W43aKOurj6DTywbxVcfYRI2cDCvzVzcUHH0XtYRQXYwuz23lwxgZBi2ENfQZM6uInRqpLwBOMecv
vzMEVlXFgBGyJO5feVRzePFZXqMd0HtR/qgQmwfxiTDIOQEfzFMv9hTx48FpkPqPnUtwaBCgf8j9
Ucn0gOC7J2tm8l+0fwQgyOGqmxFe09ZkNXUklsr5rWLrcEZsj8SfExzWoLLwj1bJvUyVc8k8l3cz
7laSvFnwBIUngNzOaCK/SSKtcdMIRXO3ObPDh6fXZUVx2Yx3z/OrJs7AO3Kn3Dx4tXY/gjFlUXWu
CmWC+oRZkRjBQ2ounoW5Dnok+pLzeMTRfmVqrziTsn4KNb5ZCpi4Djzlcp2kO763T2ye5bAdl9Gk
42u9XD/PLc2U7aWV00j6yu1QsC1brKt6/Vu8qS+peFgKQYRvPUz7poNtA+T0e5NYfaJEo0S8vsBt
Sq9ulnngIWL1SbVMsXiN6J3Avor4EddX583tFPMDRgTDJDhr8U31owBHUzXduDLE+TEj8ocL21xy
2Do5LuHX4PkDBMB+p2E53ewAwknhfjo3VHsJzLv+g0xwcqGNpau/pkgQ8zbfliH+ARDBOBXDsxBa
iTqPw8tFWN2lrNDCrAmsFTZxay7QwlQE5615bn0KMzW1dGskfQs22Nh0dBen6USHfbBIxhe+RDAr
nkh9OxrrOtftZqpOADZqfG3as6QDG24ztfxLsyTbX6JdBSvwYGDA7vvc6Haa4IcOo8I71K880zTH
u9B7qbl3wOqk52mMrn8M5NNm7vuqCeFK2VhmH2sbvo7piNafbYLXBYRo25kADexkNU/9/DxOEPfY
GaUJZZKmxw+YaeK3vvT1Ky4Q5CZgIX6ULXvcoqAEgCjy0qE+aS/u5s1W0oPlqD2CbmG3tqMmsNq9
aIXQOoDtazZWUgPTxD0/bOc6i34E0HfJoQaA9HX53C86gM0zx7rYarn7xjjqyK/NHj9vmV9EvrxN
E/ULw2lvbJW+PY0ahmtwYhMmWYgJXUATPn6+S3C+/QflGXmmtr6rmcWdlxBa/K1zEDQZRIGhx9Fu
4DjkBjifoiYRGI91ttACHh+cOWucmsZtlEX90wvQS59kkbEvPxgOo7lV/UfSSc+2pmLyFFw7MocZ
dyDJ5kKPlw9TNcSYQiMgj+A0MZmKC3tIPyEqrNtv4V0bebygimiMuk1VRoapPnm2Nkx6uBeMlKZu
poOZN7oq/0SMAEFTAHWtK6vtpIQu9/NVZSHZ/ZWFxSVCqApGtHu59mtPYlwm9Aj4ZR90S3DxUoC/
hZ0ip0zV++yTFhCYUyoctHn4a6qerU++CcT0O2wryECrF0uoLzKqEjChbbU5u38+3K61eE4mEgzN
V7AmzmbSUxM2eOGamyd0YnQYmunPguQzwMcnO2i2e2Ale3AMpdojjrfG7sV/kQMpvUM/q/Q4/a++
E17o4Gh71y2bccMkKIynPwIQW0VpNfdjowWUxujmOIXZHonMXEdmf1diNak6+SsaKS4WXgcExbCd
QeOlg37XPv7CjgLlhf436K91V2iYa9QTE2n7y7YFNiH6A+1iPd7qF5qq/m6vW5cu23s6OUNW5xSk
OWyzcpwceMedSVsJEDSgJ4mr73zaW72H+DXgO1STFAJvT/a1ZIUyDsvTMR0Zg/2nCieZhsUzri9P
sZiQHQCL1XIeuBuCLfQWsI4RqwRaClmCyMqsxej0nkxSAI12A0vuaz4uGtizjZXwyIPonjgXuHPr
BuJ/hF90EyeNeDYF8IQnj97uzD5U31BL8gEH2Tl2MaBBS5ZHazQqGPmUbyqFklbkhs6k+sXxZAQY
OehVqgjzD3svLy21wJ1GjeW+rD2BeM7DtyWG1cHrHS6dtKzqWiN+G+EMg4FG/CIDH9TN8dWotpov
NI0aG5/m5H9AUDG/y+ebCIgISJPn/m/ijy+CHXjaKC/g35oyAne43ug8fDnZjDjXcq3ZXIf4vaQ2
S5gwvUGDKlUbTNf6VJyiFeSIeDHjGT5ppehOKMh3wfhMKEJPxCv4eRfZ2cFDzU6DrW+7xZThsEWn
XIsjzA/0iZnux9e1yp/dUYKbcX8lrTPQRZ99EIhAR03pnC1gI3SAqmp90XqrM3PdfhtCk2FrpxNQ
h+itw5YDEEsBjEYlTMjM9zcCYiua4UGaS003yj1BA1RdVl6s4apijOKhvjsKz30jDWnAOha6yXOX
tKYaqHuDYk/0VLMYInnV6XgH4muDlKjrgY0iQj7niDFlaJHDKOLrOcl+W6O2FHJhtWRpSZqQWFYU
b91Xj9JR4FHw2DG20mliU7qFk4aMbiFRjvUwllqLoCwmONP6ydyWcmahhxoUKc3ioX5NU/3dKXge
uaI/wIOV6MEdo4ybO8g9hx0ALsRaddVbwrDFV897spMpzssLfHY7dmdDq4mq/XvLl+efuPgRbH2R
T26t9xV2Ao+TA/xbLKM4HZMxfe9L4MlERG8TynK/RR5LZZqSIVljzu1zZTsRIq9Y1og5r/9fS0CY
pQacKOGMc49QpeCpZ/I6i35ubcf1dwIMbAvB6obIwmQhylIgtjPKtK3u6I2StyIG9ol1qyKbqatu
QNGO9988xuayKzHObcNPCDIsEdrxHNfq3bqnzXCITxZPGOovQHbXOVpWmYrhTI0lcmyYu+KVhIKE
S5pBPwy30YK5qkHWLxfbbyHGAgGP0jIyUv8wWMwLNbaGEg8NUC52zsszAdTnBOcUc7L22GfRQqJA
EIpRPR3QUZEcUcYqepDfvr6Vj/QaSJ70RiH5RA3Sx7HrBI5Oz9J2p+f7OjKxZO95SL4TaJ9yWXnC
4hXh/aVr/516sT9JP5hNkKFeUZXLSxnR4TDukqnqmH4RM3DQ0jLjbkr7Dh9e9a/4JgyD6312Ufnr
teNVZsb/PWrPBLHf8KOx6tmUv0roe8V6MyYPuFGY7wydhAWxz1nsnglJaSw8hcws16UXF7RoLP6i
tgG8Gqv88EqBXu/NMZj4L+Mfyt76chBl18461Dao+UJGLA+wpIwZnc0t0ipeuqXitv+NcEg8qVgb
5swg5RduA+cE9jcvAX2WBMFdbGdb/8QChrntOvjEtxnowzzQ/mKT+ND04lGKQR6o65w4FOMccegK
hnxHFHQFhR0CGQB/drD80SxEMudkhcQ9/Tn/VaaSwAFCYRySNAtv7FkKhyhZrBXmZDrQCJoWzsNv
ktI/Rayjkjh5w5e0u44Qv4lSfRJPI6rrux4maLE9B6rNvNte1o7r42e366l8eZ8c/gtj82StpBQI
1VPtroyChBVgA1/3/Bt7iyJknDWZAtgHxI1ejwyeK3KoDdiG/fBKbE1afSZJdlltQewWstnJr7vY
rcJ6XAxirEJJnqXmntv/DjWVGhdkTupgWGq4nzyhOpMoKycdyHW1JLyxqo4PGevFS2OZHMyVPpXy
fDGSlKQ76uBRHWtJno1HpXriV8C+yLpzFuVpE1g3+RExGj6CvQ74Jjdb/nGkyfncGP5XmQ1NcA6Z
NMIqy48CjlJw2S7tjl+hhA4YGV2wgyjAn/EW3EXLQLOnbMlD1Nfsh8t5I8NGC6Bi3O/kNqqhn2y0
+rpnkSW1r9/oYHZEGQjz6GzMAeIuk6YFG0qFbp4uLj3k5mVsI9fA9fBB8WSgCSxU0Elp7WqUAtjD
bqCLb3svbV067cDEy5HMBjilzmNlIJ58qNqP+B1W5ZERxZSrfq2MBrn1DT4J/o52FsBQ0w4NCdjN
LBI18mUyegsSgV2aw+HrkwVKWr8aG8AxjnefiDFv47h/nTyLnHVNy6Pa82pnQTEXljIj7O4xw6Oz
qCO39B5zQGXULSDZaFV27jb5raOUHNsbhuJiZ0EohDvjJvEiKcbgjAzhBZ5P7LdMuHl1+dnLXxCC
1TkWJVeu7Z5JFOqQRW3xzwNKmIX1E29KF5sCUewYU96oOLaAwZzqoUzvt3ZjAWIOaHgAeE/eolPU
cpFF9kZEn4OQBUsk0vcz2wcg2zOpEpaFrLACTWIbjLpzUIZohTdkHpQm3O8sNVGIKr0si7OvkjEc
ebVfChP/qowfTHszA3CqLDcCj2z68wfMFXKUhYyDht6ybD1mQSYDczq0lIdTMvINgjK53tuuKTcp
OjnohQ5qbVCWftam08cwEgqUDgWpRgDeU+UuzaylWrrp+41W0t7ufz06TmQ45F9f9x9EjA+mFWLv
fUqW0cbU0HKEGo5pzNAd+K/1wZN0uJ65PW1JrimT2BOR/VPCUr3Py0USwvXv6bBOKbn8Q36UlcjI
nbSm7yPt1z0iIdI0u0o7C+VE5hFQToERsogRr2PvZrT3/SNIZf4q5XxgE9AtoMP97GyKXLYmINdx
sXhCw2JnTBrd8nPpd6vBGJp+GTN2upCHsufHvWWJbjwAj0kWuuh9c2V4s3XBCEdsaXV+SQnc5Vx2
BVb2r0+qYh7F47y9cjq81sQwAun8Pw0Hgl4JAeilpbPQpGTlrfKVXtge07gVEXIgFzdA1cYvK8lP
0Lp7qyRc8blGMol36HQskD3BjWGZ5C7WH8WHjvzRcNAN4RZospdDv+71u/g/QuMq5YlP+Qhb8QgZ
2YSyJpe0mAdz5X/tKUmnWOC0y14jQRXwUWvnB67gCeXCHCm3SmVW5tRHuRCgpY3wfDd65iPwio83
sEkcLBR9POJhMRE/K8um64d6ln67EXFtbm6x6xxTp5fFvVrPzj3olpr+U9ACDk3rbMHlv+QXW0V9
sig22LqEYx98bJbJfsqMa1BIZFF8upd/KCbJ/zgBtKzCF7CtHTBKPuy8qJt8cYlXR3+QYob78z95
JvifQEd5GyxHwvavsKlbbvjv990nLmZVWgGf8ct0ajhN8fqIkoMbY9NbQZSRuKV0vpkJ79oiF38A
mwP81uu5xwOXYZWYtVCBeWtE2cg350gW8ec8ne1OJ9kAq8We+maLKNlQokHynwqgJCsTCI9i/H69
+D4nTCW/ysxDFujgZjf/U1ek1q9gywVMSw7opi7sOtVdONmdFoxtWGK66qrhOtLQkHfxngIY0mZe
uwB6CXd7xVEBQUyXZjOtS5tcdud0ozWEFb+M1c6JdVjn6F6iYUo+lYaq8YCipTXSyxG5rli9+PhE
ZSfAONZO0/jb4QWAz7UbZJIsUoq8sHWEBGFMQRiCaQ9NqF7JKYegW8Xlc1sRFKkKhvwhKvSLr36A
MiXt7yQX6m2MpQCN+n/fjeL/j2d+pkdVFZ6IB3OqfA8W0pOKn34zFbnC19kaVi0Ea1BIXY3R6OrP
pPIpT7uJ3/Poa1iLssJUDC12Saxs/ozust1GEVprKjU4oCLED3uuHAJpF/gFPRFZr8VxcUmsB3CB
6vnPiCvD736MOifwJKbOTKbBqcxpkFWOWTf993Jk4EWfupPXTHt1eRQlwafe+OJRpzZAM/mZp1lB
ldLW/MR71J7OGVgDgxprse4MiDBbDFsnaZ2bb9EAqTiSEuH64cQbhTtD0DFaq6yF9+n/tjcNl+Ov
dgR0V6/Ks8ydw5j1GABaIdl9gFGqk+ymFGFEHHDzedSw15WTXOmYnNGVjctKio1CC9H2sSpzMQxp
PtP7csPz5LaWxWJGL2jsTHEWBPFy8sqbm+PqocVccOUwfwE8HWLWJcppkHsKaxCAa8EVAquiukcN
OTxV3I6XVLmIb4N+roKJzQ0ltQxAT6sqQy3JRucihi+E689LZd4ZSEh5+ECo9cvbG2hc4ENENmIJ
+/M2Ykiw2PjPRN04r7/gQmzgcvXa/3uuiXru0VZUInvlnMtVYGIhkN9sgQUTtLqdQs0BYyRQiV38
IZQSuaMuwTArFTF5DgarUIwEGze9aDopiBrpfsg77jGi7yU5hTB+ji3eijV3VKIarPAyZAERa855
ITsSOtnuma+X1dIgjIGvp5+FFNcHpvHrrRcdTJmH90AX14GiCXDPZsUaMpFNKEDDKnozYKwD8VvU
gSmcQIOm60hBrZgV9JCmtXU2DEP3xAbuLfq9boMQYHy3KNo0WILA0YxD5Vz4ADiglSjy1VHwljvN
J9few2c2TcJTsqTu/TNCUC7tjW+rGnaBquH4Y+6kNN0CVBjNEaDSwtKRIHcwzgyIG2Wx1VukqJuv
F9BeE8eCafbSj654Pmjd2qZhco9SNXSNmvgEf4IBrgvyoVLjJv/EGkdzCv9k9IBpUSAyEPxJ2m9i
Her04I0+vXzm3+COinSbHuG3L0V4J3sRs3keBEyq+O0cPe+A83aT/1Vi7w8uQSQwrIl5xuz6O4Zp
LChP+PXei4CNmNuKi4OJk5odaOcaOhhVHywt7hWvMPDkq/sz1J3DXmzHJz+MInXftESEE7CCCwm7
MqfF552VVF8jdnJjrAzED436oY5MzxckK6bM1Vt8aepwFjxLSlRu12hfRMlD3JJ8dsMmB7LxDtOU
vNQzhIDXFZlQb24DSiYVRKHuuFOUpsq+lRI9g3lTHYPYZ7X2q5XU4qLX82BK6gd4FEHmOMGO5A2j
vKItJO8sCnw9T9EcD/IoopX74VzKaP+wsuHFkzpB4mRSVRXltALWHvvlbDGelI9klQAv6ZQZwg7H
pBTNyvNtoUM/klIPH5CSavvO4FPY5vCFnfh8alccAyFU8okPkQGK+WMswAeRPR2G4ai75KwlbCQg
RjT8GUFLtWkuU3mz6kcrimdCA0IxvQT1fCQqoP00W+NVQoE9bkUBN9c717EqGB5tsU3Jpe2KSxcK
Wif23mbgueuxAKZ0EiFZLWDoQPsHrjoXcj0JU+r0/suz1xnxpJDZhTRy6yRqQ0nVn0a0Mzscgcq1
yzv/lyiAFQ0RI/U0OnUjcglwmtqaX2gaWo2vRvRcmgXNMRcJcOPKp/8BuV/yZVu/7I4IhxBTx54E
FaTkisTprM/1n6neLs0fz0xT7OqfqohcbzuJH6AuMsMSQPj1y0yJUC5H9PLqe3AYiuipYebzPQii
X9arYe7A6coOYPbd2365WDKmE6FZAB51t7PWIvS0x+Kg0UrZK47l79FLlqG9Ij/WMXkeyMh7pn5g
K6rtZezigkatXKaZo8yXy2xE8k2AvFMpg/HdXP1TDKKe1edD2vl/gWHlaBTzZZ+XpoZtF9u9i3Nu
XwFPKXK0AE3HTQ1/WB0eOcYZa07H+4OvJ/0JDzpwoy4Fkbi9Q0oEXx2TCJgvZAN+8OpUhhCVClT/
yHBMuztdLw32NaiIMKxeeFxYoFkR5kpJwrpsavrROyPMd+JEvy6nzrKBaez1n6kobLwRhL8zUjdx
rkOVqo1wSTkHOXapAqFHfG3BIs8+eX9txSMOpdlrzHY3wfX/+zacnEM9k4C3zRtEBuU9rOVB/L2n
bKh0p3s366Nezz6YGBO/rHNcaYu9a6/ceWMHaWL6CjheJxF6h40LMIeFdYEHslBIXEQLyBVSDxYM
3T9WoGLYK+N94OyFcMHysbBmKkHPeYdkA2xcKYY8InXvfV3L6cXY9L1e8/wDUIqZ6cJrB1mnf4en
m4CBbqzutCpafIN4gYUfPt2UKkJeJtAQ7afoTk0VwcCjsW4YaFO+deOdiVCafWfukvGBfH0z0oSk
JEIz6bz2RQlRaWyLb/4aQB2jhJZMTp3oSLmyohh6RUYDdJQzE0WRhLtgyLKJgNe06mugd+XYdp+G
WxjFqYKjnhuWc5uEIsiAf+a6kgxsw/pQPZCpYvJRzBonKO2NgMjSOLbt1cD99heQoggdBJso+Nf+
XSUguf0c1Y6cm2iGk8woi6NQWPunXSknaj7yO5W8Nu+ojsxpChircX4W666nR7/bcedVPnfo/G0R
k9xPHO0hYctFJs8fLIGm80Q7kFOv49G/vpAWfhvH7IUr030eWuBwn3WRULdcfYyQ/Urgw5EmPkBp
QhQtTPr1RAnhOhcFknzuPjDrhBKpR/tWYmgPOqSVDOvtPTv8spFGK+EnCdSlUnjFpk3CDGwOvJMj
eKB/knHg6b+80Du/gz05cdQLvRdkgjecN6ZsNhZUygbJKKZ//Y20liEUUWYHqGTHrYdk4B8hXz1D
AMINYEU1qQ3jBotke00p2ox9AKpNOURFqkH1toeYxi5wXEMX3VhEBCZUvhPJSCTZot0tvruXaFcp
ZuAmd/GBAtLHbuI2oyhf5CXUjKmwZ6f2ZUf1wC33SYdmaqTj3hfoHERf3Gq/FYe0nTNaDGUMESHo
EoVcgcjxFagOw2K/Yz3B/EKJW/bPjkwfDcqJwb1AQ1kOce8sj1e/RrA2LyUiv/yb+jdABZxeTnEp
RscHUD6wBHcdVkF4Oy0bdIZ9WahLLi9RjPin0NhXzIq4yJoprR6rMKGc5C2g7Xl/OfBFjw8nKvIw
liJyp56E2RnDkadAumo7P8WKOj5NgncRHtlw38dK3fhXrg7dUY/lOJ0AnH/dXD1O0eVImUGI6WqD
M06IZTfGkWBnTyS1gdYo9izmXqiKmDkva1F/h2fitFhV1mSVAoBKDIMA4p7RwLg5pYqLpi6WJtqo
p4dXnjjCl+mXNsz4jEQQs9+1+I491f/fXQOQdVAFbDKcAAmlEimzp4q5d0L5TSVMhBbzimnSt9Mb
yhgzwVV04pMge5/WAIgZxt7xgOddhmlj2lkgmDW/cWw0g4JZ9JdBTZHZO2eLxT47pLyNt3hejPqH
oLVgWLX6gNa7r5dZZBuREVIev0x5P8WsQmzxrJvUWT189ESYCCBu4Q+b5DHqmqTdQQXLLQaYsrNa
QpGI0iTRWAHJKG1D+Npv1V9hPE2bxIieOszwq/+LxjkeGZO0SW7gqRjMbwslI+Zstec+Ocl/jydM
3SQ1v61XVcwoJVujg2lmGm9m5Xd7lIrVI3a2nxvbo91Eei1PqncyN1ZAAvecCRDJCVeKcTiZw/qI
8EVMbHl6Gu0A8vzxoGpp1BmomADBd2laqIdaOKwCMnYzD8uIhmfrpiJYZC5OZhkWayIYGh5G5cS6
FZV9E9R/bwMtOqCDJo9+eMi9TICSO2G1Ff8Hb22mMfX56QiaJ0/Yi0Z/is5MT0NZeEUjPzR4z8/x
9vIdwJGML4ec+3kvXjnXHzgaFcONc5WZt+bquukBJ8Y0iXpQm2djjWw/BQ8DvQ2d644id5rmwkLB
zEbgyGeiLhLaijIFX4MSf21JyEykYCmc4xPXjl3Ih9ZWwd3ZI59fBmfXvV4BZHn0OxliQE4vtJcy
X61cqC6TrhetDQ+TO1EF/f+uGECSfQj309ePbvbBkX2yrXmYntr5ZIEPh0kN4LAzr149OM26TAjA
1E+UHId3cZNbKHIHPnKHF3OKTAEBNleOqNI43Q/ni/rvRVEifmq3TMxtHyWfutHvq3fqL1qNHWhv
S//gkgmBaU07f8gs7QJuiWi+r0Evz6n9GSkKN9/11xkMx0j9q2HJWNNft+jloL0ADuKes4GW0y7I
yy14sYzxyKfv8YAbA6JqSQgx0MwqR3RixDykDt3RIV09MRTYk9gyDzT8GXM+/P60H4LUVAOFACjh
WbkZamONO5ZvckRA21zwCChu911rsv9qRfeXEDu4aBCJrcp3kXDWT0H2gXaKA4N4G92yOKoiAnJL
ytQK2sXhehF8zZmSZqlxfsoGWA+JfNKOysVRt4QviFlseuhTy0XLlMHWXZix65ZFgvAoUEPmMzZG
pW9UwAB7PIVzF0ZB89O/CaThC8cU7ixB2UldWzcxwPvdrJ2yOCpAqnuw50HFWOsQ+8safoVmvefb
qXlWgUx/nEHR1aDJ4rD8cRIzXzWlVS/3urRrLWzi38AxpwardpohfBudESpk366oHTfjumzgQbYx
MoohHRxTqD+TaHS8DuysbeAMe3RY2bYv7ghgTtgCuDaZG2u5EmPTolko27u7TsVzeBim6vumEiz1
xWjP+hIylydJ6bUmioDek28PhQ7JaqWCu9W+ZFUxptRLZhsjnm4+zJ00zCMFcvxBJM4XFoU98qoW
oFYMyfi3VJ6x/WkgRbfpnN4HqDrowT8QUYlIjTVoxZRZ8Tm8XdurYODeQGkf2OHYNEa3HspchFvd
bo7Rk+17YeiKL4Fi5a2JKXef965uxNifmN1aI6npuWOcroW0w6BLU1OhwsiieLSdev1bad41jyH8
rLnarkGHhTXqNwqv359H0oksq5FGSIlKgHujZWyjlMfwoT3Cip+E3WC4k2v9KBBqoTzr29mZHjpr
lyuKjp4HsBJGd4E/dnUa2YWRCnlf6gPEUSvKsksCvBA089wNkRr7Be5LO+mZRzwWa/WQ03jQjk6y
q8Nsj9xWQYjskYwEQF2AJ8mPADSkqmqOIEGrMRE3kttFIU20+lROed7DrFe2rg9kbEgHjtPhiP4l
CYBGCbPNzdBWNKJCIJ2jyVQnRHKBH9BqbdcxCHkpCiNWnvgiW6GbNmLQTUINxklwV97HQvXJt8h2
5bjtP/OBIs0KrsUny8WydFHa3Bf8nl9hXIrDqYQbBooiczvj/ESxk6YWXbiPyR/XbmUGUinAUh47
4N+LMseS6a/7vrvXG7GNtycMcP/LL5a4qO/jV+8Fz7ccE3B53fuUDZ5nxZrJXLODQsbUjA755uyX
GfMFMZMo0sLShSbYP5HIM60M2vbxEFZMsKpnhnqJGygLgVvzBXnp7dICqa363iA5Pj/TPSOHgIk8
ytk3gpF9/1rLUYlxDypLCpW00Pby+uzxAhsZBt9LLJRy3vAme6HQv5efOd2RmpPIlgn/tDEjw4l5
7f06u4dX3iQnNrA8cGlq+OcRFHIGqSG1L8FA14ioMQd/2QUYFUYWiU+ZyI2p4dq34hovTGwobCB4
L3A1UobYicbA+cJKIZb5Ii31ouJepVuOH5DyuYg0lHMkfN/+MkRRGasE7hrCttwnpT3bMxWNmw+3
PqLFiD09DltCXLTOO4DJ5Ny30gMUKitKu3lOSGcI2KTLGkBR0HGehaCIdkbIQRSdNQHavLzuU9QB
GxNPS2rsbJVGshwrCXzdOmhjSpO5VQ6O1r75yGxljJVwYkKpdpUKqX7Gg6U0VlFXKYNcyE3FguG6
/ichLf3Vl/eHZilr6MeF1Ss8xyor36VNNd74qlPsmdNCxLVV7PTyYEp9T6QGVjUjeH+Vtk6mGQc+
r6gCsUQVrDOGh1a07vyc3ewifpZdL94+RKaR1/L2Q8b7acaSTVWKbS1d+Ax7zXmiAEgxoIUWiFPc
igUcggCnCHcPRg7NkkiDJ9OD4WUrWbQkweTMGi12NtFV93ve8SFCxSQYaiNCSP+39T04CL7atUOb
k4cN79nur96Bk92VCCzX6oNtlmdho5hviAnn9zHQuBfYBHsfAkbz2g6p3rnV4kqwSsW3iRLNqobZ
4zhMOGPGNY3oNrkfJaaSEdcngBGBIC6GbGt+jXuRDaRWe0w4TnuCWlL86vzvd7pvtF0KLFlzWLwq
5uEf2O6nIwCQowqBRUg5G/AoT8A1LfYNQZdScNB3MPujJLgFDik/wRc2ptwZwDVoIE3aSeXIiBdP
LSExUPjwAc5YFOGemQ8oQltOvPnhAP3zfPLujBOnQkD0rvlRByyvRWUV04JgjqiYSqjDh831LYd1
bbRLV7uuz5kjLrwvL0qzvF73UPtgXx/aF6sJkMjVqVZTNv7ymRK0VIp06+ht44OpeXjc9BrTGACT
IwKRKbq8/2k2C120ATIAmK5443lcSCwQBvsXWaAYvEi8H1Xm7ks0f8ltrafH7mLVvWD+S2tQNtcM
QZ+EXMVM221P0FQXOvgsiaoqV841XHeWxqZ0LLps/DUQoSuTR6uNFlztsMKXzDtzhlRSPd6KN5Lx
ckcO9ebO9PO8wy4fskCCJtPRgBKyyZ6C7hAHEVY/pZkR77kTzt7vFHrrQx/TAl0KDLx+UdSCHuKa
7fVMD0EUnnewSVTgtVpbcFeWhM21Eo/meRJeNjpCjU1zr7hVHEBbLXcmR0SehNMb+xmRlpxvenGT
XtITeM0prY1E0dIuX6rWq6VTBiuMijlX13IZB9VEMGupfbiGje8pIf7Amn2q3T4oVBE6BoT8San/
X6R5kYihstZuB18y99LnQKQyO+aQLOefAZiqwVltJw705UH4ILRbJ0ZZmKvS+/bT6tRk0lL67p11
zi48ubnIQC0q5PM/IOy1LtZgIervQg47DpTeXTy6KMyCpof9Dnq2H+ZhqHALvjqk9psmrzjDZ2kT
v6kPb0hQC9JiYHUu5jIalIreERDnY0zKPOcQY9ARnxgZIsK0b5KoXRDJ09lN+8WX1ZCLIfiQ37qe
5IQd45ECSSyZzdc2YF585e+TTGQyueMCdgxhvGlnzMkzAzFnCF4drxAQiLTb0awVL9+SEn7dT8Fv
ULjospMGC3RNa7CRpQ9y8Iv4Xy4dX5MgP9KzitH7fLxWp1ZjiogaL/ol2FwPKpGfF2PADSxr/DsL
Wvv6vrXEAPldTJeKT6RLI6NcK7KovHIjnjO6sZpzpLP3QFhniCMIjFUoL8DOWf3+BKc71skmYO6V
I5XmeRsj6h+ano964PdctIZnAwx04VS5aeTA0i0kYhRZ10Ifx4kpNJr7ncUK3jVLRrnyHPPnZu/7
6PwTY3OwDQab2aSnFAHBdNH3p0YVRDNPBT4YQAu+TX2MqFoOdLM2wtMz3BHKib9P9AxvcdNJKXk+
FhW0HfM8KmdIalEIzB5mvGrT2dmj0VyivQJyjRjPQOWCaLvH9AskxietGTdYZc4NLW9ldpaCc2WK
Mdol9/c17r78vgklieYgpSs3m9Y1Sk9N3I6nqeHZGrZ41NDiVKnCJejvXeQb7wwwdsAtCWLbi5S4
GY8RISsDFTOwJ8n+L/AElWAME5iR7qlWG91j9Fkhl07V1fRJ6nGS86YmrSsNaDEXEphd4xrnDcOF
iWCzevTZJtQYSMNydMYQa1nOgcwZc+FysfrNB/FljsYomV3QM5HDPlOFiSQ7jpF4rQI5x98VC0tG
PhaWLV1xIm6ci6SIB3nXDwyH7Gk6IiGIAOXQxsFxFiytIyQm4feaWxso0AUA988n73d5xqUK4/pG
ERaL4bSERXoq1CtGHNS9WRKznPmXCYcV0gl979MrWRl67MaHdBc9/BqFyC4IcqQryE7ZIPQPq+zQ
4Eh+Vj4xYuK0t4Et6oNxAi/JoAOyVhuuCWMa/I8VIWPYrv4bbbQ7THWMu5/Mt+l97k6wvII0DnH+
hI40hmf1Dql8C+majfsUbLMSaXpvkqJrciPm1XB7qN3Cud6sLTLH+wwkWdVORPzmhzFNDs79eGar
GVafBgNCPSkJt9GtRaTZBO+j/mse56DiE+Elh7J79qghT/ISygaad+3QfYQUJuUZx4GcF5UipdK/
ZmjiJmZqe7xOiEEkIlsoULbh5+g/f6Zm59N0sbVU12m5CF0FlwhQvMo5CS1MJFaZAelpuyWJjcOE
L0um9iwBx1cskU3hGpUYa/OAtv5+GypQKzvavO0hhDrFl/se18Q88VhIGSUa+bQ1k1OxdUx71lcL
zLwA6gkBeUxIkraMDetWIuv4jf7obDN4eGxZ6gCGB+kjfC4xJbun0QN4sWG1K9w/cPBEs9tO6Lze
U3LiMSbRYbBKrl5HK4oFTKx4t2An6DdQ/Us0s39UvWVWH/X/u7dUGHz9qT1qDoS+WB8wuNDXrdBY
TUyzcq8AvN5kbEQrGj587RRRYBerLNDCQDiESxr+8oIvhVCPRyKeBcjcwi8yaT8V2LFNboI1AiLz
SWsld9UZ/DU3QXSAMMOchOmLqgtWepc7gqPRg6EZ4aNIIg+tt0fNxpqANIX+aHHD3QaRgRco8yFl
LbEueIJZl2Mpt1jhijfoi0qc2Gq2dPsafvYDltoJs4WYE2ZW7ptsxjfK3n52grA0KTpl+XKLuzoo
YQXS33S38oQ9dXshd55Z00FzVmaDXcRxXIZUBXAR9eFE+onAP7zSBxSY4dL1Iom2cgGkfMuogOp7
q9X5Tw5bKXzQUQFcMdslBTiMWOOrK20d4an7Y5azhg9uEt6naFOi7xPwM18/b6dnrdSwXlwV+srS
zo43CV6mAYmjk6hA8DCq1PWY4unddfdWUSsVio18ZlrGlFtskEqVjRo4GZlURiTz+M8zhHPYzak3
t/WVLCu2jOcBBfws0WS2gD4UQ9njkUjMNgtx43Fm7yUnDqo/JVjCP2fc3VfiSjFn3dPqlx4wf1ha
b4en4pvXlegkhbvyuU5yP+CTsGrZPYZepRkXmbqWNNB20+KpSEUvYkxwqgxoQBGV78xSruMPj4Ba
Tm6ZSzfn6RNrpjaoNCHwox1iFdqyUC8Ly3CgIYW++mueg7VjajRIIO3LGkOzbvqzCPJqpWj087so
0J6v/fplEiA6QjakRAD0U7+9ZzFtj42BVVXWLy9gJhzhlFVrDdYLwVKPpHe3PMjZj6PVd5gPyd3f
YwWMeoq4g2y0hEpvJc6DRDeFp/4915nbeVPhVkAVxGi9yyBV785G6M9ND1zTx2waggF6rGRheX++
ktd37iZ/Lf2xqHlL/A/mBkv8p9Q3WK+XAevQ/Gw0wXx0KNLj6WFad/daTocYvGW7aQZAmo54x53g
2A9mRIeZWTqVDFtWlvVE3mS3QOEWCZYKdebgSlozcNLhnVFf0vTVEef/32sZhu9szCiPX4Ht5t6X
xWEZ9/1BcuFerWEn9GIGCR3W/ywWTqxvkfJoPex6Pr1ChrHTGej2Zoqf3kwf7GOfwlCYmIedRmuQ
yZX6c7o+QPFQpvllblhGpE1OLO9hHj694+BHS0mxiaW13N67b0TiJOVJCQRwZaj6ZkWzeNK8dzUL
z+mtNhZIWUicAXHgSWhIvY3SHWNNbSf5NeMw/r4PRVUAYxkmr8ND32dky3NQirTJdhCLOyx1s4IZ
R1Y3AzwfP1XRU/7MQXF4RNQN2I1YOS+5BYFuHlQceu79lnCRFT1Kte5I59cmzaQDlV8XcwJMPMQC
tZ2kdi+itI2qeoFxL30WuSXD+jjtLBj06kDnhZ0UbjYcbWZLVzfGJF3YAakI/0Z6jTrsKk/XWqRm
XoVKSYkMkE/hmm8Cc0j+yUYJcn6W8OPAme4sQKCd4fmvq6/QMf9XAuEbM1FyUci1LaLthhvKjm1r
49bS6bKx973VqNgEjm7AZI0vAsxh93+TUqKJund9Ey4F7A7nXmhdtOLSpwB/NjE7mCntEatmB32d
0zHQ4kIqxjnVF5P+otrBBNUfTOxpZqaBZj1AqC0jc8LjHjxGJGBjZLdLyYJvqLNku7e8RhW35irt
Zy8GBEixrlv6wPa68ZyjaK+lRD1kJdnSJhqeNCxmxEqcBb0ppLx5zDZMjUg7wT9gixXCp/N8+v7B
HGa9e/C8HlgIkh4JImNINyr+L5YqGjtS5rXWxH4KYJgIWtk7HtPcVwnDT2q75ZdfTDPuEVbnTH+i
50VJGMioJgV3HTVhUw00Fup8oGuXNfEdrIbeL/v6SbIKHrSjihv88SbJgSc0ciGc6saQllLYLsss
jb2IFCNBacXgkhe6zOZCOMbmxxE8ugtZHJgaQJbb5gkY6ToSTwNJM1+MP57CBFZMksssylRvhfHP
go2bwuf/focTkVFkkKd9M+bSvzA6LXNEfnSS66tt+/zyi6+TdFeR+dj0n1ISAq+OkmWbZ4H1F1Fa
RnQCI0YnyZVb0DXRBkQauQYSJLf+pooPHqhU9nXgM3HrgDUkB9V0ZM3XWH4h++3UHkK6NB7N48jL
28/iSU+zwdN8xWQnw9f6CGo1iUZM49OD4PoBk3DpDuTYGBdOLUJXGZibp/cMLvMMwRwIrkSE0kTi
rTzpCoIswlf8UIin98lFLwy5EPYg05B7kNDOPe9L+JEkzuFSfxevQZj6kWTKVrk9rVuTCObwnOHi
mJ6wt5xRAs46BufXPGC6jz0wVdZ2LtkCcdkhUuvmyj8uLTzI7SJMkEc+KdZphUjjTDXrLx3x/Xtv
x7FjCfkZejuuwSUcmoaER9CjoCQqePI62BH1foikdJe46p2/3b9pjBUFMExZALLf0wz3luTk7meG
nIft5try/joa0lwA+aSfJv58aevK3aw+hgZ3i5fMPsyhgtLoEpqKVLHdTd1nYGcLq87lWMFJz6Q7
A9CVWSktwzyU3fKFb9KtEwzgCY074dh9WjTEfIhQamhwcR9XyKTQ5AsmhCHSmpIIG2kVXwAejQBe
LVLw4RwTqcCGZGei253qC4Rqg3dal65rktXh7bbkziVPuUZ/KTbZGc7AvxwTyM5kqsK/vwwyvDyb
38RVPQRwmDybWzmCUB/lRhDFzfxZM46THHLR0jQK99VHxRAMYw4xN7TAo/oGW0DJ+doWmcM/dype
KQroB1Qt2hZDYWtlzcdG1iOVwfD9Ko8dNxUBA3ZrN4aT/tO1aWoBL+nqC0qpGK0+jmrrQJbpgBOP
lrfBt4xDioJAByU9qvv5NR/UBvw6Y5kiv9AJevQcMRLW2bILqgra+uEGKgvZVp065RawffXQ1glO
5ELFIX/8Br3R9Jr16eGK+5Ys8gTVvG4AsuckGgBZit9bCRBy+NLgcn2edB0f0f3sZSdRW4KHWZju
6Av7uqMorjEb/19PdschnxYf0Fp6KG4W67f3vdP8tcON5w+Ug7y5G0TGHUxSVyHeGJBiYIMy95dd
3LlGARlFhUtnR4vmb6fsSqbGEh+r0Sar3BIkt7jwHUuNNCoJoq5hpeHD9I6t5uHPmwZp45vuEIwi
KAiZjRMLHwjkvSOEEerkx+EA9ySU296nz/sXn91TSjTnlLlaqo3iLMsjrVkgcXsApL2LH++KXkDx
OnlLkXXfe4XW7fXwKJrc3uFVz7qSaXtpu1+ieKm1Kqd6LbEJeRpjb1ZOSSt20WjxPishKGRQ3p3Y
v4jZVGY9Hq0huj5H2OXSesz1+aStTyFvwflqJENlj01713Sia4M6bWU/+LGfwnqUx5TagkDmgDXR
xL1WNCD5imhOdEWc60Rer3tW37IAZgCkl4AfKUgs7Eve9/ucOm9sLabXgMiylTSDuGiOjev9+/rC
aMMPbzxZVGZ4wsdUk+G7QOqF/6tYzovVooflJV2qjs1Oq1v0eSCEbaZeJx/Hy8Gfn0uzUGe1qGlA
3qsjjX6NOrrMT/k1CzXx8pxGBa0IiCffK0s7Y9yn0ayJbOpAOPwCJ+C85vSMH8C6vbl1Z58TpLa2
ULPALrJn83XML5+2vybZxpzttkosXxTq/RRrtylhagOOU+5ToaOG3MLV8aljnTE8eoyrr3O7c8o0
zRLB+fj4O6mTWDAWtZH/Ov5jXQy9AG6GoBbBeLpt7fASv0/99H+u43l1jIjimFl3kI4xSsAfDAMO
PeJy5UK7yq2Dbrnx9xExR08omKyZVOMXPfK2/UJZOryv2Q3fBjtlOiaEmfql2Y4k9erEtM6UFV4q
rzf8UosIl/cDGEKrW1jHF4QKpMbEOjZMJ2QEMP0qMMni9ZufpLcs4SJ+vu/u088Vxv5MWCU8a8Oi
KuvuBuBVbE7y1H1Qs6kCGuTreL6Eq1dgHZpJph4dK+BtufHjlAtLCpAfJU4zFDq7DgcIi4U4WYV6
D6LEamnJGrDDUEYHhCY+96xipDSvT2aQLQLVQu132PWcfwR5wB3dVPXULucfHZcGZQ3ezpMSUzH5
w//3Op3ET/OTvS3dFOTArHyHuLkSn0+LT9+2+cHin9HZxz7b42+t17NROIdu/aG0qbzqWH32Xdey
kctNBopiERYf19u2cadVwt/dki1t0UYi+ZWtMhaqF7ZTs690BzoUeSEQG7O7cX9uQ+7D44RLzjeH
2/RAt/pH++57b4EjjFPl7VcJAnowCSEqjszU/zCmAhCgC0CMVIiuMVFTBmMtlfkFPtgt6sEu6KV0
ksL6Y1NZah/8JXpCBmMkWFFSW5mBNnWcuuJXqF1Z5cOY+UNXAVYHkIDI80xjMAeAOO0f8zUVIQ22
NkX+t7qwFf0mURp1d8dQjIgCJ5CGtCI8EBBjmJ3JtnSLyiTZYYCgj8tVgD/Sa6QYbFYlztFQ/CDu
KB7RW3TYlxyolFyvw/HaJpRHHn29yo/Y5Ea6c6dmzcdSKm+UQoWnuJz5TZxOyLUjVqt5hweGuTrb
1baps1fY89WnErtgDK2/vcm3Q+3PlwYDOdUwH12lb7KsO0INmAY4Few7azXLyk25TCzwXyfLiic/
8VyX0KKT/bSWZ4d1WeE3vmcvR41f4GC9Gx430iK4Ln64XZR4jRh9Nu6UbrmJD4T6M6v3QoUhP5zC
WOOg3Uqv2c+hIX9qBYyC6WLnVYz+6AnH2dqFnqRVsCCyllZGLlwLdwjNokDeeF1upix1eH9r+6P+
oeLRmpGegvd9zA96GaxKUnugMD+MNFHpcMHzc45iMpKD6vy5AJbqrztZpRqNfO8mxX+ekALvbimW
fG4V6GYaWRpnsiov66sDgmfi9mKZnbPBsLyY9grqN5ZYK8DPNYggGqV5pKBv+gqaREM2okBP2I6h
GABFHAwYfA8gaL72b6x01Rg8hRZSi2TaXwcqJjWqPL8hhjHLgRU7Apj7Vu05NVTSlsrBivWevloj
XK8hRlvCh/vZdQ0tvfd+AOfRs0xR0IoetIf8NGMZqPdYNFlBDCuTegUyULi1OWfXOfBBF12gRUrp
Lm63qlCRfJeiKMv8OaIstHqwT+yHmJI9ce9CICu4xOR0F7+k52vrc5ulnjgos+Rl4gY876pNtAHc
lEI/cO+LKB4Yfjxt1Y6Kve++TLqMt1k3pRwLOZqglZSuhwU4mIGUw6pcLldQnclCx1z6awctzJob
b8lvt3mCIlV94kyLK6VKRKstIL0BhNsL1GL7eDpsma9mOH367rvc4H1ghYSz26puxHgIFeaUw4sX
8EFBIRBmMsBYsy0CLhqFjAdaRPoFLQPh2HIJLzmXLWYQBfLsWXyPEFs293AX2ElGq2kFn7B5KagZ
c+HFK7iN49PHaUcx7YIfQBa1wmciagTEnJNipQ+g9lvP4FdZdtbJqY3ZSWYVTpulfIsWqQcqMq70
m+AJabqOXLJRk2xfrUwp9irODmIgbf0MbYWCNarV8N7SH/OHNp20UWGYu14jiBvLgizjcpW2Pdek
tzQtZkH2RTCYZv6eUFLqB3Mnr57GghvkpamPoPVPYCNC2W4UxPjnUwInmc2/HNMK9S+yUWSLAehr
GYpvRVf6FyfC1Qhp8RVA/v79isHKz/cnY5XMzVhvUfzjGRC1sL/159jUFyNlJ5zoDoWH76BMQPNh
6sPGnYE/uqy2HkSovsbx0uTlYkg6hUOYup2xP57hOP+cFKoG6vhZrIQz+au5J+ewQHMvMOovP8uF
W93cYWL9Ab5YW2NTDuzbsYAgTtOjBpPGSvm+7rmgWOS5FwFyZudQPrZ9B6xkmudl4q3x1AugZBrX
BKTqBxoN9bjqrj3/zpcZ0dHGSIQfapEMLNfM5xQsx3x49TrK/U6p7OCmDfigNkuC3PtCnxghyBox
/5qAd0Zp/TBH/5s6YLYghaMpdeFzuIWr8Ml+DDIhdBfnEMVtcQnTWcmFbcF7gwFVt3nZ/xsvA4BF
nLUVSfIB8MidDdzuVYu5DtaFGXn0B/SDP7EFWTi/9OoV7Qo47WtVtAPBExJ0wjpKFKcrOpQxV7kI
NFMFx+VQmX0QDlVxNdJZdn3Wqy4YXljxZpzjTwzxDGqD5QKjUTnBG56n6jyj78fWG/Xnee6PL5bg
tE4AUAPvU5fu6Ez6uTR+JPzez8cWhBeQpbHY2KUM9qql5wFI7J77VIST8buXTgluIrABB9KYMyup
4rY5wJosx4ST3pI4u2YCynLWiEAQBFmO64KC/TGbZdqpTplkMnFXrlsiTgH5PgbDE+n/2C/LKipv
RvmCfnWvIIIWsA+EIaf/CD7solOS4D+iEImBRBnYiA0fqtBXzMLTa/AYfZNj4zfyOW6MrjjGjJyF
uUKCrXqQNjPOWuPHMcGB2SVZPmBtpeSaGk/ueXm+xuknliYLrOrpe3IQqMLO++u71CQGu0EXWlUL
n8MWUlKPU2WYh2Vjd2V7am8cXEKmzq2k1rpSHaKGlC9iw2GjTM9aBb6tv19c6KHy1BOL5qTkrCqv
d4TQlRfzhmMY/+F/Se8cvZkW7Yjwx8sgYuzj/Rw+nOtFG76gIRfvvx0/ujFat8stvBNK/WtcXjHN
M9EWEyfeEpDYtQVLGgAvb8pXPEEkYOXhTPATBOZ0ZdrMsN+7/2f7DH57K8leBOGBM936Pmykc7WJ
7VNho/5tSGNYtlK+956xDuEmMHEAyNOZg1L1kRTKXRvMz5kvrqD95XJFWWp/LLQoBZ0kbjJGVoBp
aLie3Gcj0u5wse5o+29NXvU3bmnleLmQ982kePQYyUpuQXIOVuSW6XcyMyAaBMCxgjaDcIWNPpEk
bjY9qMxdfZJox7hl+PBCNQiJnZ+i15wTAomfTPB2VmMG3SB9iS240c8q0PXq5iemdz3Ol2DK/yR6
YqK1kSRpdcKtYIvciPvgHyXAvksOFC3AHhzzzcd687JyM+O3+nqkrmoipLWeBJhka5ctAx5aWTQc
i4X+Ikb1QahYQiAdwMwQpv6Xgi+4gHf3pLGubeshh2xqGHzlFdGhERWSOeW4sDRn3EwGdlI2AXBt
PZv+jBHv/AeY7Win2bSlQaUbmVQ4jUmpnpACkNBhYpkr9UfHHFRt4mSxEnMlf5eQu/jQyLiUMsHl
sjcnHLPR6L/I9bRPqcE1dUDTgf9Kf0yeiW0VOrOBtrIlLA0RI1UhF088VpFJsRK3+hi5jXj5nz9+
+1MBrRu4BDYx54BExI3s0HZpk0X/a/ztSOe8HX3LBofZINRWmqzNmuGNz4fGsZgFzsFynjru0x6S
AiVDZl7XYU4Vw/taCVYASGmm3sUotwPApRvD/pDoosYRYbQWWK0W05cKcfCU1edF/RloGz56SVBR
boFRlWlFjw4QhksMo2zmiwng04kFHNqoReoVN2zFp3x/tTwhdENac1cysySZa2vbFje5az7ptkoB
BplZH+hjj0+j5z0RbTTScBI3OjdiW3Pmetz4q7vaJ7teaTDhH24xGQSk3ojeggaYRmpn37iFTloY
pAzeX1mYXT4464vYlP2LFoZz41zR3449vU44AjYFqIb3VMUdLD5S5vgTB7a0S62gxmAkgZuiz+g2
6XMjBNy3zdGtQCayJwfn11kYTta9oKH6q0HT1ohe6ur6DPfaAFCkdAI/RamB8DhC9006UqB9ErYO
kuTNHI13OZU0qymRAlYfQCRiimPdSByMQL7/rQDuWXL25V+YSJylTV6KTh+wgI6mhqDeS1KZ/mF9
jVL5rME8PvR+BtJfz+ClE9b3NbnjftZV0dRlr+6Z5Gp/q136mvYQ6zVbCiXUneq9y/Kg4GB3mTbE
acDbL5OsSISuxDCTeRtQDPFuxP4aCnPyjqenfMJHHO5wGW2lYzIFteIVsOKNHWzfJARo9aNcUHMu
1FbFdqtozd10/XQXV1Jh+c45YQUS7FFj8vOlHTWjPFKkOlHpBYH9206t14kmVJw5siKnVwNF6tFk
vbFhVUfEWKOvFlNtDZhfcMe3um+XLHICS3sG1wdSIL7iRsxykeTBN85zBb6AgRteYDiNLsvYe3B7
luzQAcX2aNabAtTBgnXpVIsbh/lYCkH/LQXIhHvIN+iFdrHRICsTVar9t8nXAle3gtOYjZz7X5KT
45Gb3BgTg1MfDrVGDMPsoB6s/bko5AA8zW1gY9BSCSBoqa9rv1H70scoOXx/fLNKecLwoFUtqe5u
VrRn8Sq+UUNdeDXqQ9vNGTM/270nSlZxutWpESFjXqj6QhNhmL/uhnkHblmbMHogJ0PfeaA2p8Zg
eWlMxLI69wBQEdpaNGw3ZyJRJek8kfIwiCEdYbre7JVxa0fCU/MO6aE8oGT/JcxCsqbWsdQA5KT3
+pposkH/Gvb4gnt3PJ9vcIVxMfqg/xSOIa/Qz2Zk5MzHXsXi2Gg/znRqeR84zvxMCVBBcfsjL92v
LK1BPWfmggMNZM8nQEuSQ9xQ2qw2TNMrojSm3054g/GHnH0mRvyLqG0Tbg2rmbTBQLt4Mg6ooh2X
ZfEWmZRND6Q/ROgGbff+mWwwFYLfr4JrLsOxFDyuzmU1N60S3k1kOqQKqgdUjyVGneAm+3K+2OHR
pJWYRKMy8PzRatpEk8MuPEuHRiXqP/MQfk+k++XLQtjxG7X3pHV5gzVrBLAL3Np4pSNmzeMhEtpB
gnwyz8JNq91VxHu49tTjn+4kB7598woeBRwUhkTa5D4CAn/BL5y2URkC2ZuAlfwL4FEaJXrk9Ati
8D32pWMePyx6sz/pSo/w2X97CRRR3f1jtIzsB0qMtJN88dL0ElD8CX/VaGrOthmNUKkx5zrF8yZl
osRD6b3PtqOD8ul8I1VIjyxF5dOiU8WIuOlCn0Ozk6aDaIx9rI87fMVvRTAvF2JbUSdCHXThJf6D
BQUzyjU5CIweLUz+tMaZU0/vgGSWcfRJweduGu8U70zQHA9xA5207TDUtWsqOInLqlxuJJjqUkU1
fvAhLo8FEaerJqEdUnojiqP/Qwfsurcx47RvlNZt36x++feUYsKynsqwVd47Hd5M53SGAcoIX+V5
wlnMwJNUaGdJ8y9RK6VdEauuKJz2WrvjkU3fZjL655pUQbtUrM494lgRCxdIxImCkTiMh4+OR+mB
8rNbcuD6g/iTRs/0o+VMZr6CHytqPDIo72oadSXx0UaO2AaVt3Yq4/2OC5WCYwpXI547gaj5X275
Kxuw/I8Uk5REsJkdrgPWAsSgOpjB8OsLuKiyFmi2ofbb5nqEErZwBaA7Phg8X9YgFqu22FfnJMr7
+IZDgZ1+HL5yr4/+7GeoXTCiBqXS/86LzQqoFREoApCyMteO9FlqbqMT2l/i4d7BAwP8oPBUMwjz
gZ+JBahmW/DEc5kZaRpZgrYo+CW1q7fGI3na1cCShJYFfOoR2fWWv7d+QZyJDdmWJCDqqLFwoHvx
UYPgPY4lzhKU+o6q5OMtNZK8xOIJSkLCyBqON7PMf6HUKF2s443eWHFL+LT/+SToTjqNgeiuLfFK
Elpqnku5d1MMhT1JGylEBvDSwgtmF6uJRDP37BEvjmvpVJZxEtvj1AHZ95fVrBVQxIB4md4+4+rs
U/QOIPBN1qol+wogctRkC5NH9XAxujKjVPN0nE5sGrFXYDAnLP4pKVOK8E23rNyVMlejlyhll1p9
CXKN0+uvh1sXDb1n8UDAYLlGGLrsMaJYaXvagdR+xEfOs5cqll0x7qQL5ZObzQFH8ixl2Hm1CdNg
UJnjjpqnF7ExOCWZoD32ztI9ph1Z2QbPJYR7m7BIRY6q9OEgQytCrC1TI5MccdmLzTk/Hho8ObCQ
hl3nXYXYcUgtacwqGondZLBQ1QAEE0e5UZjFYUTBkP+mpWLyxURcpNCCkKiVHiBBjhKkofIz2HVF
4v0+SlKWsuSr/IeayDS2DN2SJH9YyLNLRs9e+bVzQdEabuc/YW9QtasbKFQKatO2I/s/ram3SnYg
VjWGpJSa/g+ayhviEppEivtsiq7pXh+CVIFtjXdIIbufbTSzlAnEDtE8CrCRV3z71BRE5LEXr2N2
vB3D2msmdfkMQi8NRvBMpTWEhNiMw9Ug1pJjpj/uC42Fc9Lzj+uAisusueRrYj2hTRXEc++ye26a
zH+b6YTV0S+G9y3rHrnBgQ1sS/mh/XDuSePjKfZkk8jjIYbVwhZw5EdlxLxcI+IZCwZrU5HBdc05
NiuybruZjXNbnfE/pqymVJ8If4sifA6J8/gzBcaD9aTiMxajjafRKJAbMAJXUDcKs41uDwdlT7nq
K+jj3D9r+BmXOOlWNrYRp7KAKC9UMkmi04IoIWzhZqdhfo2Ee5qhfMfvawFpwnDWYfcnHCtbdKj+
ESMFNf//eOLaN3XROou65YVDGXf9PEXBYuaPv3SeNV/1gv61t3EKaLEjU0SaP8UpgQBJsrOcRPf4
Q8ad2SlF/oKI1oxe1RAJ6Hy+eD9hCTZOLO1bLMdU7BxRNvZ99uIFJGFMDZnYQrT1apUmJr5X6xs1
oTLfX7bhKnDgPaVpW1E4ZfzAGk4z7IexOOC2Rwu9HO0n7iEUdmhdiamQ64s8pN/qNNXMvjoR0Z9w
YdXuCCa9zXBou49lQA0lj7qOkgEHlkbbYSPIZgVSGs0SRuWHu4N/l12WGzQGEdjn85cWQXShVlwZ
526x/qrhuavw4z8Jd2SyK7Pqy1FzcJkVQyoo+dvGsRVWLygdaAUBL3KPQYl08DSCf7K0yq5JUW4v
qJlVp1iYe2lUIptiPsIGajo+VtXrW2cCBZsEJ/wOKPXoYvQJTIAB2LZmwcA0+rfExVYke91ozywT
MfM+YbIbClG6HMTs0pTrsvpIycv4Ps5sSEzOahl+6VWNRWD8l1+V/WuUc7TY96JFMJOfm60El2UJ
LshB7uC648qzTJY63wVhe5JupTzEezB+jVlS76XTC1Ytezy8R+Lc9jm7YxgE3SQX9sNinDhxwqsX
VcbpngPQFolFuCfYZQgL+UGErN5H7Sn+6rDmqhZwXb4qOSu1+6eeKBx/8/9eGeDbhfPLYvkIZblu
S09Oi6u879h1FU7EPRzihQlUCs6t7FOTVgCTJUpCqbkHhuxxJ+sAW+ocmCj/pViE6qv8T08ZGWgL
06ZRsc+kaC76mmEAZcwAH2LTKaTfaTQox11bG7qcJ5mK+dZJAlhsDLRxhslMLVyidGZvBT+cxrh3
4InbjYOc+8rtEADpT/xDv26HjTbTROaW7832VyuLCn0pJ5piAGZctxqqfQe2m+rMyTzZ/caTBL9S
mICfbe3EU3FsbYHSRctSB04TMHv8MVC3FWxCrcgtZ3QhQQsmluRA3ItR7w8+NHjFjfDtw8K8kFu4
mcar645MPg3pxsBQpJyuN2ZmZmOKouDFmO93RD4V4ISBRYKj6yoXj27GbLRJZzSl4FlP7aJLgQuv
lTlluQh2LUV4Li6Jo/OULuGOt/4HqhcQXLHlK7NgiN2u9B0zIREZYkLnlxVm5iTXcwCVLnA24rga
nTpviezHb4lXlO2RqL5pTcfI5wM6/AjVuQlTekwZ5veer7tOzmjshHfumBTs/AWPk8znU1iEzNJW
k4FptKLHfY3aO6bRrmvYY72REk+DVy1Sabdjwo7eAH9AAgdqajoQC8Og8qUp05elzvhubqnm14O4
WUHoq6Cr0dp0NzfcX/4w2pBhkybi26anU5vwMHCD9paeGDuLHyzNHxJzwjEvObejGlE5LpdysPoC
Rq9qbzrFcdLvvGB1PuP7p0+CqzfJ1GvvDEgSuQyca3/inftY2mDhmP8a3pLetrU5JNBQuIvBqbVC
PqiLA+uZyWZSHuswdlt8TDLrNEye3H0TeDkBdMBHHNUWsWvpd2ZWiZ5hr0ka1/e2G85ZomJIaKn0
YZ6imTraQ+8obali1pnF3ZZAAci1cFH+6RlBAoQCIkTDjfIw1R6uBo8Slw3zmK/hNJJO7sMAEHtn
A+zoaRM/7gATLL8uTKVoeaM9FkP/+SC7tXgF197oDhzu61/BT8t7yZybcmM7dbWOaZ1ca2o5caDD
IedGQD2o7T7HkoBpLXmabxC9pzFef3nmba77ZGfM0oyNbgBfqXkb5dol6Ah46S8YA+4EZ8aFABvj
N851q0ZapsVMoCLgXh+VW2+gU+vHhzplYtD1oVp9zeTaiTOP5yRX6so7k5Lc1XO0sqjdxvdNTqm1
o90gAt+i5dMRPDtK3sNt2DJzCKrsNEFdfU0FY1K1m0ScLhsi+nUU/lFVf5q6nUuaYwK3fEo37whh
nR1Ar0BSa4S2JQnl9p6ROh2K13x4RRo6q6wysuI09O6urtagOm51fMBvYiRNxho5yoKUCuTJdqCN
FXaECr7Qw3lzh1AB9ruX/2M0rpdKeUS5+8sVK5ysRo8TvuDK+vzhKIEm8Zp4sWIPE8pVHckJa3Eh
TmXDxMdaxaO1iwexeOHr7nwtDi19oyeElfcKnlJTHxlbt3mMyAWEtYod6VDEiXqH5bK0KjcSk8Xp
OeFzo0CqIYsBztoqJyFHLfQlxOtL+RkoWBIqAvOfbn/h6zqs0Y1VjGr7tR3w63+CYtkazVmaG88M
ZGb7T6eRu/dQ8xoFhec/YEIg3KYxPUazKpTONreRzvgxGe12BnSj9QqeBoXw0BXcD7gH5gq8LyFn
4c/9Do45F1fN+B/i4qqzogl/RE4acTFQcSyY5Xsm7+fCHFUXw8xfwuX6XCuWHrdjJ9FG3NjauA+e
L4G62C6Pl+3M5a+iI0ipv2Z8GNGtmDDJlhywHHkvScTDZkVHhmDOD7tPnRcEmLwPD8+rH5id1t5i
N6Z0LLWDbEkjueCZ0RHkrAOu86s3dKZmC7B8izKO5sf5UBj7uNU85oUAlxLQrThSnig2wzF8hc31
uZfWinj3t1aVE7p1hxT89PQ4oEvd6BlAG+6DJSegeErjoQ6DiLIsz/YH+nWW3VvlQdKgZh4l9qVg
wd7SocGaREeVx5ZdUcVCeKlcBdd5v4EGxoJGT3qUTLADIjro927tMF2qR+T8rbIb5gavUzjjFLWL
aXbp8GjPiKYbFfWq/08xWupcAqjxJjbxMW5pPmsd/dEcMqhJNyfqWaNDpqdUOeCfnRqSYmFgOcYv
uof1do67QfLqJahvH76evU89jTTw6HtmCAfwNAdDD+GUwZA9Obuas8YF3H06l5EBttiAhASJSrRt
KZVjohQGYMg4cKO60B3rDuD0hSuwvJhzM+xTcrcs4xy7VPO/2op5y7CeBVuUetYL59Ln0jxb2+9G
5Ds7pztUQ7CG+4/IdlxT7scrMzVbVKQQbPXTNSa6/KCSMHMRjWT9FLW/uWL2wGxp3DeakxzDK9PX
kOwBCKwRbbKGd5c367kkGoM9ldpT3xJ14F+4nen0oVOneGQf4VWYid1KiMZAkm//iGbRuwqKCyaX
1n2xQZIhyKQ8CPdZ4iOU9W184RkRznLIK2F8k8Gic0pubAEGyDH4OfnssiV89TTKCb0lmADQxeAb
lRV8H3xtsKuTkLGqt3Ya9Es9kFs9V3L6uUXlE8zkkSvp1f2nJrvX3f3DhAwqd9lXy9eac/zpfZuO
q4izKkUsWBUu8Xe6uwaPHlyT78Z/rD/eK4oSv3lcSHSXqkWmdWPzZAR9qun3GtTIA18c8I4Ayesg
1IGxrGXe6POG0yP1Twfjz0wpilNlbBVqdIbBPI2kSqqXm4RdmFpQGltbXqnLAhizmEjGotBz27Xo
LutCVsk3AVX471oFciC9lzhP/znjtdtgo9NHjjmkjuSIFG16BrEAtzf43udI7zq0fo74GPytJPzE
sdcSO9oq10e0alChyh3miYh/mb2p2uj037KYZ1GyFA0UHGY4rWajbOs3TBK1nIdo7uL5P+duql1R
Ze73t/6ECWLN+S6ghlZ2sFe/jdEmRlPUUby2YEdI6ooeCkrk9vAqRHsKjoDzk1M4SB7phwJG+mzn
elR30ZHIGxxoiB5YFpHVjeZeAsB0vMzxqfd10VuVgRHQSxJS9vndg+tJeHIS1XuEPv5O6j7SAriV
floiwllJY3EHngvygQjgR7ws7iC8kHs8PzEhlIFliNmFvwYpHjMv3f41NCkIeLBlA+yaI20hZ/wP
rajpbpwFkpMlRRg7CvUsfWN5jDP8vFdSvI6+a3kJ/c7ek27c58VhPAgbhXZdpGv7+sKMAf+uTvQr
D4QgDaiSjddqK4XdJuRQpSwLuQfOC9mGt0hvZhFZP1Syz5UlQ/D1gbMepxx7rzsGPm222lvU2sca
EBcnBxEiupmyZr7YhIC0Uj4cLrGlzlCHfogt80/BkpVO906WkaN7NsKZzQc2/oB8t2qGQDoDwGLw
w0+vLTjNP5Ne1JeQ0WttF0sSihNiKKyC9R+R0hgSRLGzeqCdjsafmskdIdW1lUlcX//4qcL+Ckp6
6debPn+V+IsNfFFQ6W1NdUQULpYBgkt+29XIXQNdsBLXyqVqKnsri3q7T8DhJkaBkHnf1o9TVpyC
mcnzzQYI2azN6u1f/3HUYpFk0BF/bHRHOBykT7V0k5OD5zO0Z/A4QWq7K2b9kjpMnY0s4VoSiMIx
yDOvI59Uig0G43idCnw+h4kkTE3yM/I9ZjNCc9vTihmqsK0XRueeJV/2JS7ePLJE6t1pUmBPu9p1
yqUZj0Wkjt3w0Ba6A1fZPn4WkGYAl8+JkACr/8E6bGQK03iGL5cwGF6yJcm3XJgf7LQluUE/eFDz
zUjVPu/ecT5qAqsJlydQIq349VmvRIMpEqF39GyEbpVuDXAJQVoG0K7oWbO7dI/AqYSXOP59RIBC
mcqhVFm0foCNzXznKzrZSREQVMfj4eoWJD5EkNiOgFxgOZyEmCjGhXiV2XXSqPLRuiEeyfDW5+Ug
GsWQPz5HnOEz/+FQoD1sqW/1sP1rfds7ZVdMtLXbc9jHwI+Y76w76YMZ0NWOIc8LZjMLilw69Z1r
zsI+gSkFOy1ri4GPj6yyDs34R+PSrqMH1PVNlCsXYqSeI/Irr6CNg9qbtVsJS57l+ovIMhOV6gMc
knlxQay8TvFrdIpDvv8MvXYPe5tZWVcQfGQiMlrtteuekhRAXKDqFoTJ5VkJcxcVF4CXNVciJQZy
mwqvp3mC+V3uX7A9aiyYI2qGMNl1hFYqirdqClIXHLd/eyzn5NbU7CTRLV73oZcGU0rEznwcdm4W
VSASP2MCFMhrR07Tda1HRN0gSW384q94L0rfuSOEDKaKWgzqx7rAz7M+wGHrjeEhuhj4qEySDR/s
8eoQ461xBMRA4ei6HGzXZ5jX0dlu4G76xD0H3pUXuxDay7s2qtwRQ2YSY3LgTAkqym8GdWo5AmrV
uLYJ6KtkV0R0eoR/PVkKl2jQtZKlJi2TEkwIOu9F/FMMZ8GxA3Foxug5tFD2OpCBgNrxWOVZTTiL
cpFfc+8a9dMI+xpZnbZA9xMUcWfKdFnr4n7qnVOrlV70AhYPTilkZ56wyUSliWZZVFl4mJZPpFv7
+PKcvRUk/dHhL5bfUzMU+QV+/fvhkmEqUBQds5PxN3S5N8LZxA6ZHWrCJRacaq1XPs4mym5F68S2
/dfSifXDzqTvKjiqO0UcznmbqpE6srs78U+0LqWAR5MnLMfk7w6krYvhDZ/FDmR8SZYxPTBqty9H
O2CgoHStY7tAUu60DDzNNT552j0Hf5uN+P+mfXzSAMcrtDEQsqn4hglWqXgI6FTg1YcRxgHTRldp
fLr8AurQarCj8i0L6MmpF3ZsXJIBAJwaBO0VMgTbnFzksZp8nluxugfMyo644Ps1beLqmT9cFQeW
KkJVTTIzzp9hmHTZS/G3/j2TMMi0DRSz2JypgQfFie6RfsHkoT0POYDBygVp36LRJ+8uA6cpLHPm
7oVKSZD2N1kkC9a5jn2WXNuJMTcCziQzmM1yqcGlF7DKpjqn1KaXHl84LA9CuytRI21lAF26505L
mgImBs+WJUxaQ4ai1ga063UFIi9z0ipEqJ5I3XYPeoEMlwd/sxOA8U8gn/fmjxD33oygFGwN3BwS
SdusU6YLhyV76NRHdhyZLdQujAMVw8dXtAGn2MTE6dMwuUnw5QdwQWd5oo04avQZfCCVJdgZH4uh
fKy6U0UTtGAJ+vnjp9j4ArLgSLxhWvTOvJ0TQiu5JLmdkJkEv2XSmT4ppbt+s8KSHoh/jdFWqSNC
8C6UX2O1R1LJvznoZgm3XQ88mTqZ1Rlubl3OeO+y1oVXIXxLMQhfQvTg5266YVhoyoQkEZvV7P5i
0eA+nW2O2X1PczV02opbwX4parl6Q0qASewDTAvnonCvFZU0UYjH8cwQ64PJHTl+MrO8pWopflhJ
jkZKRDa7XtmD8bHyiVXAgVvjlM+PHm8T98pEhmd/RpBCRmuaNCwj3opPb3Pu1RchMBFWe7iV94KE
Uw9RlyD+SJ2T4h2UGwDSY7caZ+f+FxhPHSLBOFFYmRK024KP/KjgP2yIzxxNG5cgKPklrJfa4Zpr
K2Wcdqf2fkillD61Ezb9RVzToiJBCAQqWVN2S1z1HA4u1qfOPdQCjKgiOMvd6p1YHg51tw5ayn7y
Wnqn+EQkyU91O39IGMlXthGq8u8iR2DaG9ov21Ekf0lnEYA/OiTP7sjSTySa8oEk9KUTWUGha4G0
jJ8VZ9maLgQ6MOLDJxGi9yVYU8ETy1BTT22d/UsjJ1reSUjl8GM4CpOf0amkxbfGOhJzA6hbyrxf
vTVPWzELjjpEGbMqu5+lHcREq7PIZNTLGdWWe3TLRgkkMrxPFzQnV1i78wqWVRBNJCiFReZrI9WB
OYMNnrB0c0SNYn1aj6f+WSAwGy/OH0gHsWfj2PShUwPBSCBYP/UsKN5oqih2CpktnUsLUgNSIUsb
uuWhKfJn7BdBikDJYEDZQDobZyQ/Aarvefnp+K88P38MbZns8TBEsrsWjg+nTHtcgArm84ShjvmB
GNyjQS8/tdLtembq1zVQTvEZItyf1t1MKe89mocOrhQUMGIqu3WdjeB3vUOF7zeSXFKhJeT0+HIi
l0/d26ziqVw9sRHLwuj+Lbj9mE/+BMxPWFpyP2iN2rDFjdI6e6LoAK97u2HfqgPlOpNgfgvN6gG7
d3Fc8PcL1cgVeQ6UfAA8KW9Rw7MNkA0ovERSByFenKhnYOYGcyFYySkAZOfbRyEbyfWyEUJ98sHB
1LJjqzML8ZiVYqQoxvc9l84nUusn5+3fzmaPgrNXgalArrBJXbNjXWUcjJHEvzJWj2m/v4B5AeW4
vh7YLvzpPB4qlrMWeJiHMhHz02AdUYbV1gS7/VMN9h/Mad2q0TwJxI8EHnIEnR/Sbmmz75f2Voz8
Kd0DKZW4NP5w4ayU1y9g/8glMb86ALYQ14/1zvA5xbOSAqyRkUhn6PG8Ney877O42QQuI8oH4K1P
uZo7dG9hntQVpjjoPQ4PxZLHEUAnvJyk3yvRayQT0StWYTRhVrCyd57MZU9n0q1U6IkfNeYxwJs7
o6s0nWPXBel54t2FjKNDYhwsSRsDrUYCS0jzRtH4PztwGjqriELyDzCHJ8KlOlzqSeaYIhpVsVqq
rMZwQtqrsWwFdfcTByfE945hR9g5/YHBiM06YQoT2BACgMPheajE+jeN2Z84qJV4JjdaVcDMgSz3
c72C4KqWPlVVrjtrwrD+FmI1bkd8TKC223c4V3E6x7aDSp4skHifeB61XyOn9sjVS24KiUKlHTPb
I4fsalXFhy7GeujCpVTY/31bIA9isl8BLCPMrlirFBlvzBWIIqcOLJW0pj/snaesAMTirS9d6fpX
QGnb0PxNH+5lzzwXwfZIy5/EAV3wluU35erGoWzEZZ1CPGRs2X/zflaB2CBOnK36wcL2x91dhrfr
5vuwMzhITrcBiT01sIfSnMwLrR4G8Jh0UF2AWWyoamhYwpty+gdIP3x0S/DkoGMvOlbSyq/X/Bqm
VVcDjikG3j2MefGxUZwKd803bdb5bf4ac3dix48uPaE00B4Lzdc+5k6pJBIEAnF5vqxDgaZX4h/e
bPeVj35cGLs4GESKBe9cHYRJLHAksQuLxD5NVxDPXbGlz2+f//U6+J74jPnDwZ0dZ97GPDHs8lFu
4dBrqmb3SQsC3Dq6jcqq4QrgNhRMCU1tBfxGBHESyAyUDIX3oSndXR9LZZkXXo4iQYWQATPfX7Hm
qfQUW3y1jIRO4VklHpY9UVv1+jLrkjKxHBxtRCxoZ7uTxzHRQKAMkEC/1ItHkTrfmTYbaAKzjYE+
2Pvu253DEBSex5dJ30KSwbTQNaJYFjmsxwQ02myUTJr3Un6PDRH05XHRAYhj4L6IC86If3/S2W5x
FoHSjF4vfQsNMahZe0gS6gWdCoRTiSB7DEYzcVFEU7UAqDGm0pdjWgV7+GS1AI6pU0+mvvYdSTyT
yDnNzNfUVNMiv0za6TlSHLW0ATKwzUFB9Z95uCoo/wQE4uQGVakg1g5stpMwIxZKiSCVg+Eo3kqZ
rWxIpUzbjL+MYZcPS4gZxVnBdcJ2uh6LxsKtdx9fNH7gwwojjMN1yD0XHj0gye2dQRJ41v7LyWGe
TmDQlG5G6H+wIWo8vKbwQvrpWL3o8azRmWCrNlzmEGT+GFtWoXMS1FoxVfbmUJlkeA0yEWzLiNra
av/q3RFgZqziOXUEsSRCx7tEEBoqL8/7lxFVjfTJQDafHWSMBAIAdR09xwBziqS8zjKHogPgSc8k
3ebLBCjOFkGj9f5q/udmEvcNf+pEEx2K5QEl05xupjkTOSoBPWBVC5+MSL28mhT7ubYREvFTyfL8
e5poSLZ3WuPpmvJeHJG9wD+6idTyXiIAdyJGhuB4poFphizZTSt/Ek96b7s96bxOcABvuTSSpoml
JhRM3wPA1a5gmciLSAiumJ7Nyda9OOq2M+NTPZxfDRluHIe60uWSRjkkT943cqbYbvcA1Ku6Irre
v1OKiCrRzwSyuv/NeuNXxwZx8rYtKjFJFQoGR+7w9y6xU9DZ87EknebqXIZg/1oeU/GBlS1mMHnJ
Wdm8BrovFW7+vMOB+F3LJFC89Nq8onRixj48FBtIcfwRi98Xg/M4qz/r6j6sO39Vd05nXpQ+VOGX
6FtPfqobSciFu71OpxNAzbBQxaVI6vDN0JXXIRmODQQChFa8RsJB8ddrGcTWvGeKJPdfdRF+WHIJ
0i+MBQAhEwcupw1N+CCBxIS5H4ExBd1+eMMzwvjpfnzathH4nTxKekKbyVEaINiCgjxL2Xc3bi1l
41s/hf444JT3F0JS1PJqmUA2cEwih2sC0aHuNzzm7AQY8np7dWDUJu0rRNQSFin4t8oHo822+eun
UycwodrDzKYLlnvWb5ObrK8T3+DlJ4GKu9U0MsLEy5nTGvZ3yQDhAl0aVCoYcqZ1dvFGjhzIpU/V
pXxs6wr6ZdizoGZMOZVShpfu+ICnuwcvwZwFcXJET0ehRxgrf3XkNkgOLv0OaZSsj9/0tT7bbow2
1Q1NxGDgkd6RZjG5DSwAUOe5rCYzc1ElR6g/Y7nF8YidNcyEhh8YIxj194wY9n+vZ9Q4lkkzwdHl
+SxOPQQRthzTdimQVrPw3pBSUa30y2ZFVF72vIUCY/yaoCj/cpuqXXZbvV1SP3/gwnKayuWvHbvW
CL+l7nUZdl/eFjno9JzfHF13jLX+qrZ03ldsZJ2vDTBpoF3U9flBHxhfz/NZL/ycEg7xAzlZjaCA
udLzn56mAcjPfA0CYEF+Pe7HZN41PaEMMzqRf8Hw1HFUnte/dX/cWlbmI9XQu1lbCNSXAXcgV/mh
OsNtM3YGfSmbYm9sFMmm/72P0EpYwd6E/5kZ+AhDGRfN9Pa8VsSWtnIi9bOF0YCNxxwy0gLzskP5
X/2/T722+ObrfH3OdxpfxzxV/5ivoba3jUuiHaRDcJW7iZzNORiZmB20NZlqX4SKjnnzJsZbYN/q
QXBwCgB2Mi7pOAi4fmvh3C0R4PweVJ6d7nUQViLL7+UAOeQrNBUeL/4hBDamL+pgKMzA9LGlWJbP
z3xUbuCJKpZOIFw4mniYcJXMuqkNjG+Rxz5yRgx021a8b7B/q4zNJnj/CkfxA4Pbjugd8sQcl8Yx
+QMW6Px3AZN3M8JhEluUaNOlSnHfYbdoA6e/tQRDl6pPeU4MIUqO9uriK90vEoRqkJJGiv4WFf4c
vsenyFHAkXb3QWE5mYSaONmIGAx2wU2e9UCc7BP63ZcmynhH+97vbhIe0HNmdw/pyAaFjQrDNOUU
NzB69mjWQ+AA8WnteW8fLIInO9fEi/oWaa52je6s9bXetQ11l64m+fSpEn0Gd3/5RmQn3KuHHta6
Pd/4HiQ4uh5jOJoarIoE8c1bjIm1huwvh8NBqnRZTfCT/XUp0tSjVfuSvLu3ld6LmWSGFz2Jkuum
tzHhFLqGfN6lnI9GAKBuUqLz6Jqxz9ECwPqNLDFCPE3BjwM1QedKtGFuaCb12Alo2ikKSMSJf5+V
Qly4JHOlTjjg7vx8s/+5ZAPBhltYn+kafFcDYf41ISqNw2zF5pas2w/8SJuLEG5yC7jrh5PEKUS3
3yEXgcT1YnK1+ZCrS+hyoQYiNt1k8ER/3olhUZZ2jaAKyhjRseDjNCOsO/t6eqOjJN//BsSJj+nD
ZK2Z3h7K1TrLyGCBKPxhpgxKSHNgwxaKhkRSytfwocTETmnivWTlDaJKzB40Zu8BMvXZiSEPMnyJ
U4K939k0yQF6s1muwGx/lfW0wZmKN1z7wFkOZwhC3hrc0OjtuCLpVRVnUPeRG4pYfcnzmCq4rGg0
pNSea2bEpvrTiWiNtGuZmn4s8GErGN7Uev5DoA9en071q7uC3NGhu/Y1IYMrUD5Q96C/Il6D/2Fo
K7I2R6/038sG54GLoFUifPgRZlO++AfTYDk4PFlicASZqmRzmw5tY8T3gwicPo7yiD+ktAkWOQQd
+LjZIoNyJ58+smp5QqtGAgcSxd6fjWiZwk0Tuj7K0+P8zdhT++VXkVsH1l2zxem7V/dckuxiB3An
TZXjEnvfpFuCSYz1mXWR5AyxvC3afE5weXb1aKXS/p+tKpUb51hIiHWRa8Zm9L2IZU4ZbhIAN/ec
oj492ZOMYzc66agVwqsfAAYSOLNWlyKkRa9HyySbuQfmorDY2Bp1CsMkXCBJVAicKTRPLn8YcjjY
fx7s0fEgU5ogFK7ww+2DpQMiRZgfZgQuukMYc5YBtkghW5C7hiSgICQCq6NoYFjuWCrs2l9Hv1i8
Eh0YyZ/5ULYwnv8wJ0cIi7SRmpGNNSTBFw6nW49vLZBEtHgjYTwfV2JonwZbOmQlJ5zOrwZlp1Bh
W+jRoNmhKHB1vtVYOEJkxYpC5CSxstyBFCK13KYLg/4WdnUh7K2GsCHn4cREHQcAbCa2PIy9N7OU
Dp+wfW8QKEJe+He+0o6o1paPvzZn+379YkXLqsAUmYLU5uh8rOwphigrQGIeUWX+R9Nza9RFiFoK
dBxjC7hlsfy5qE9HUELYHBQxrbG7Wp9oNL5mQNpHRPoLnrzmb3JT0JkSgD1zt86gYboI70BDLYh1
0hZ/P+/FxwWkYotG1aBn8zB+jPhKGoHEWS8Z7U9tWgcFYysUX0WbmaIygbVMepZxNny4R0RLTCxJ
nTmt16dlc1ebm9gzu4AxT5Ln55mPO/SzY4Ym/8BhLFPOHM039KqQUk8z/Q+QN7qB7hkx69G/jRdM
/s1t7EW71d9SF1pCDfQ6fiEX/J/69nn7YBsqVAhrTV2qbWfE9lBKeLYAtYlNzFBJXr4n+dj296di
GJX+qP/R30Qsyp8xZXnAYnmy1IJh8hzR2M1c1wUANZfWVoB7bBfOCJDMPyq8QHz2HaTZ7ktDA9xy
tYr9VpYZmsb5LmqLOCaFtTReL5Evw8SvMZvGLcCn1Zguzmg/f+B+VDMjz1eT/3SE1Veob9MrBTO0
sKcUMK/qgQaizqU7gU7+1mQ1b7/auV3y3Sf3WGz53Cr9Wr6T/99gXsl/33R1phuC4haudDCyfcUh
7HBORXmKUMidXJ2CEqvaktuiauzhY3F0drkhVZbS6/2SCGCNczKcitWup+khd5h56M79egZ1y4PV
1UIIbtadJ1Fs89tPz2mNdbha3MNcfzOmY6ZCpur3q5bAd+v71jepuN89DvYwaCzcrgsuKwvN/YmC
rs04mvGF8ICqiFZtGCzCqyNyG35/H3zCLsAHFCvaxmFyBmglQX3CSPlSKguWtj0SL7EtnIGsNF/2
5bpnTZAP9rcjIQxJNtuIhv0MHeRdUZNDI/PeB+3W/CUym//V/Ww3aMSMpVrWEOY5d/XG3pSFyF4T
3qSOPm+9C/iz2e6RwI98W4R/iPSRHjUlv3BSqHA47+4/mTVLIOAlE5urn6vTEHuV1GxX4eck74f1
ZlTrzFidF8/3x1/MJ7wYAuZt9a30Vagr6xj+O8Anp3fJD15eYZUEZqoPSm6ZGio5xvtzLFb/Vdi3
HFKnz2Tbf9TRoDRBcovZyrwHwwG9KtBnhhbS+y8M8t2XCq05oImNw4pR3HRuB7jiBnlxOChMsMgY
HqXMYCDflCx/iQZ6Y15JwckQwH9o8rIYYurkaLHysUrLPR2LOY8cSdYjuMd4YdbsRHIY46A7hp5h
JDx1t5Vwo4pNNwkULJcTr8Dl7a65maz+vnMXSc7ZMu7evX6LeUlhKXpb3Y7/kv1PiYBFsapflY3S
KaooCzEaHrBbMOZFoPjVFy2U09xm5dEP2PGGKbm8HyfuCDA47/2MmJskqfNcX0CeAKqJEtadxCbi
KINmcFo5Iu/Hv+0YJa4ddcAEYkiYEWqxP+XB9TZMrh7VHQvjt2978TG0QXIK36s3LW6v7PNr+iki
zKvQhCxMepSGIhukLYt7o+Xn7nked4ey7p2YYDtcB9mqtPduZM4kj3KRh61iR8HInt5IsnwDk4Nl
0IBlSh1yOzHATy9DVKB7xV02sxy76r0aQC1VQOmS++ldfvVJiJCvb1aWIxEtTU231s8V+pY0jJ0w
b/sOdEL79oaNV9wK03hsr4M9o/WdZdnTysl3xll/LnP3c5rKavRVhhC/scHO8foOWWEjRdj4t34p
3DTyVJwtzaRmM2zXafs1dnluFSDL2YE0+AMCHO4Srw7F41DuDf4qxoFzff14B74kZm5Q3as6ikBe
xAO3xRILzZSrgXU6ALaTdVaQLtiaOia+B+QasUWafN4+h11UHslW1o8ApQEJwi5CRe7u1w5vimwi
PeTN9per1/rmIwPxjSA4wNLkcPoREzokKgiIuoyVKcAE78sMKM1HmnihIrKfGXF2L/HxWPTU0hNG
FkzdmkCCl1sccQpHOgDEnHoShMTAjvhqszMnvQLWMI5y17YW44op3Vtj4pXkLdrxtilC4PXHg6ik
BmUSzeNrOvnR8hrNjVn00zB5uoYvUzmu9F9LoTQcwBRL2l0Q35DIqiuKSiCcSJy367h/vrGe1kCO
mvCobUFP5cYP5o32u9a7MmJinaEH5Cr6JTeK9w6zI20J+QZ+XKyMu59B1ELUYfSCLLlTVvwNVUZz
gBEQpWUJEPnnqWTVi9IxNU2cQz/+4bDTbj7w+QSo9Kk0C8Sk6ae9COOBYUYLExqxlcqPpw+pnHNY
8+cPH2x03f6X2PLkIFa9hwYjMjej1cI6Mc3tyyH/WY24L2xQMXB6ewbcF6CsF+OAZc22aZi8sAuD
/IORkhowJExkJV22MpLsHbL8emvbegBCEQm74e0X0BuGDJfaAxSKgfIl+7oajkz0xTcjDUeQ2P5t
upvy9XG0a+52Af+fWAAfVtK+ZaA16nTXtdckLHLsKKOthC00gIAOoQKyqMk4lwPSCBfSl4loOE4Z
A2uFfoYNmh+hoHfxGwbpyKfq//NU6pOC8rrz6X2XR6ozWAwJlInBej7Hkzjyp/pRdXPnTltQHFaU
5OJFoCjeiRsBGLaHCAUyej5G8DaSUcIFLtkZ1i5wL5iUR+fqP0/bwT+S+tImssnTMryDl0Rx+eh5
kdg4UcfCrKoqjGMH1I1z4mCQXvriKViODWCIV0OxOLih6Q50tsaoQdNZgpegXSGnhu6MFyYUlxu7
tx0fsO1mLGzSavZHD4KlU675Kb/fpw+Kv8iao7MgJeG+VpGp3W/7UyYmWX6u2uW+cKf6iMZVX+BC
ovhAsMd8rYziIzLIXLusakG+lfRwJPVu61uZq2BKWkJIVe0n03FlKXNpRSj19DIxN6q0hQKiWmkL
9q1NUY6ZkbxI8D1FpBml8D6fP5Vum+iZRo9frgk9hDJPJoM0L0f3lhwGhrBvKbU+U7sU+W7AO8Gu
vbvmk3lK4eos254EqgmuyQyTTqgJ+AvLZYaWAdYQKxwmP8Qqdarlj9e2YqG0NnCj40wq+Fe4S06t
9m3Mlx7DDkv71ABdIwctmXyg5nnqIP/DVd3Mg0ShHB96QJWQjELQX6C1fQ0mEomV8R9/eLkw3EiN
jXvFFL4mEkiBFGAjec6kYWSHvcIiH/hrH0B/zukfr4Z8vnsrfG3/SCji5x/lmZX8Imd3ll/Jasnr
OxSuGkDZrsTyHetZTd3xMQjlm/Xkz0FrXzaWMBqWTBDAy6gtx5WNd6Yy3HtpqfsuhTuP1rgiSPCU
C7/lPmTCumL1dFVNoCfqOO9PUyiP072xWmPNqB/dz5lytzB9PF/gmD4G+YJgmo35ucJcL6GAF/zT
ykledOXZQXUdvJ8VrYD2DrwmCCl36VzE7DUjRikG7wvsTM1pRD7+XJGxagYyNDFpL9bIhDS8vY4Q
vESqQeZql3VHE4e7oE3F0f95bDyPxOH0ZV2/yVvpaV4j7TzGMoURrBZLDO8Qvvpxy8M0TSRpILbj
h3l+mQ4SgsfZnxNySMDVJ+bOo3QfUq5nfDcphLYJXKnXoqTCOrO3lPc2UIg1ECxS9LvE8ge56bMg
Ni1Taz65OI27/wP9gvvyH8/rcSiwSW2nn39cAvPS0wNW3+O6IfOonIiFNxYELQ8eW68CvlfNYPWg
m1xqdSgw1VVoG/2MWCmi33mYaMsgid+Idrk4HNYacTkJjNiF9xxMhI5NCAK7gY2qMqHG4cs3pT2z
IXSoHzLPt596+eL30s279oxMMQJMMVXJyCMgkWb6PIitYuw8A5w9R8ap+8TNio6CyAfO7khViq4w
kBiMT5BEbgufHcUduELpLbtwV/CaeN7avMNGRtXinVT04SY92WyJyxQ9CG6VG+FRxLY7siWdGoR4
EZ760wwonNMHW31CXCVR6fwE7QFcFtvkz2By5QbqajWLdi+5iaTnuazClWEwF6FsBqjjKp5RjRT9
8dz9L9RUzXKEgm+obc/g0aoWhNAC4WAzFA9fLnWNQ7HLzbAwYzM5fptZIXqzumP7sIQCBlne3D6d
7KaRBFO51axrfZ0jXZnBgkvhiMBKlhI8bqICb4q+PkWaEPwL0EjLXvwSccSdvptfjeAIorF81XVC
3dWWOJRipJuXA71t0Pveh1waiaEuZbA+sKLRhs7q55nHDNYKlvDJg4qyTi8362CgYzWDOcVilhnT
briRd+0xqDVwsV/IUyIK+/PhT6csHdTruvcU0AyYg0NQpa2wf7Wyuo6HBMF7G1gdoFysX71ZToAs
XjG99Z5jqxLeiesWic2NZ7/iu7atBLcqlZePRla0oYi2Iit5kuAu8tlzNBzn3ygIDZ608F96RyFH
FymcThB0S4HiqSk30d6ECiFCOa+6enOkYVOKWcayMoF/QoCg6xkmynCJlAytKY18SyBWRb1a5opr
/E7Ukl82saR6+xzeUoDPm7Dj16pGK9NCCEPl8qJlgz6jRCq3nwpA2VJBuP1cjbSSG1f7SnWCKp4i
KyTZTw/VuUM8rDhTvItJi3dkf/NrWqLkxGnH9rXxZDBpE0gBsHIIbbkL4ATRCd/rKhs/JEju1nvz
RUsV81uS1ueZhxq2qLD1S28FZv1i+UjbAln9hkbBD+VGxI2f3Lr2i5OZxfjcH0twB/Xp9CAkdo4M
D6XriqKFvjXiikFXZWvva2gWlmC7+syEE28Si8Zk2FWlleFzh9Uq/4a9u+hFWWWHGed0aeedUoIm
A1F2wj0Zs9QAC7gL7iR7ylzBlWI7ZzSodF/bxjQWxucJjOqGX80dTqBeFoBu7jv4DA/LLuVfi7fJ
5FloMP0hitP2wyNiBJLUqQbYi9rDASLN7KBq6OZt0kZSueaMaZSjZryoa3B85MhRn5ciSlTKIlyx
46Yl1NijYrOyIli66zm6Fbxz9b+LoEBetwhgRkvVTBfeDIAd21QIXxCpSMCW54IQGDILLW83WEBg
bcQNn3SDMjOmsuKoNN/6qAGFyOIPZeexxEAode7Asp4eMDyxhSOrpO5St7RNynArHBcCCMqLdLxb
z7lGnIizNrU3lNr25CB4Lx3vm4giZIDpf4PCnbskbChoIX6LWoh8sAoF1NjhI5SeXo+cqBI2r+EH
218CJmhB99FLMJ4T0GSK/NuS9KUobLurp6bwFjpLat0kHp+VHxIy59Ufc0gUOFAgbbkTI/+neb6N
PTHEpx0V1NTV5lcn+ws2M5RuGhCSjn5/9yCYMP142YGfyyf9if+r1kEesgdnxf5mds6ZN0pJlYuO
bILI6H1YItWl2u2hzWQ3I0iNL6q2FneNXQ+mLwkwHxDsa3iTW1OhjlhCMXiml4FGq4UxiWTvyemW
w3f/Ow/AxiQOq117ufdgQRFbBhDVa35S/4pfENYqFMJJt1vY8oiXln9SOHrJh6L9Eq+FvPrvoxaD
nLfiNIIVNXwzRO839+BuNc5XCrBFloS09ByRrJ3wSdd0BQph52OuNZEgoMR8xK5fB1HCGvI0nuRr
RzvcD7uTBnkXcueuQPDuNTweXkfykMdbzOR3zm1pePN4kRqs4Yy5hZw8CeN4VTNEuDxy3QXKnaCL
Z8+r3DmRCYNdrj2wtTANUZEeuCs7FpfTBAtguveggJcZexY5lLS6zdBfYO5uJ+MXo1ENMFM/DwuV
BBOWhYPEWfTRIUViijtMQdfzJ9W5N28GYwJgscSrW2er3r5TzOiD/bDFpSrKE9nNxnswwRdNhv1B
UMAy+v4R7FHilOEodIvqtkP1HaufPWf2N8ehQPLd9mYZMidAFJxiGPJWUvNRTlXFHkobvqZD0sx2
snPJ3nWQk7Bp7/yuApMzD3idd0MwT27zoMgFONsNn+3hRJwwOBoi623uHmD0ly4c4XEp4ILqLdqh
jK775QHCiGuhQ5p58hVJvGEZE2Ie02gBQA7EPBtjoulB3ky/zRz0Jhn9EgZGouRX1MU9XlyVjhkR
lzDmZ+YUeIUPzMIp+EX1+gPpmabLENSpaPnVmuPorPyXyWbgJ5o7J4aUn9jYmGiU8YGpfI5djCmK
zDcLEzr7Mw5enePXLR0ylL2WV+e8MkISStTAmpwmq8jPT0LFo+9vd+TNr957OZz2+nEM8+Ea6ShR
dZZDWyJqoLkgHFpC8qKUvF3pWXFw3aExL8yZQubHBxBlgt2pHu6Im1++jx0IyKz5hbz0E5aLDdvU
rTZwiEGI9UB4dVmCXO74c1SoDRKTrOpGcEG6qSX5HQvOk1fn+3u6kjq1mt4nz9i2Jwb2JEheoqyn
ctdOuOBFP9+BkfP9zE6deSHbdX3xI/J6jHnTpY3kXRHzAajn+iKJDdwp+rrlsmGqSjeGnSRzR3Bu
DN96vOwOixtwJx0IzREcfV9rcKZNgMVIw0M36T/CbUqArqc+ehkspFWxX2EYKWVkBjfPMR5BY4hG
ZbDARknvB186dcFtGRgAxtKsMU9Z/jFUCsTTlI4qIwKbfekDByzaRtAqzaXqcmEat4Vru299rOWD
bowASM6M1r+LAQ+GL6zBuoWz7xDws5t95hzaBJp6iZneqwYPxC4yjbQa9Vgy9fh6kpMryiQU5Myu
HZm1OWVBlYAj+vtKZOBjq1+0rlQc82fYAK6kyEP5phW/MbIYQNZO/jwe8D+QbORTW4MzO3lWF3DO
qQiEmk5VmbWBQzCAJ+aX7BZkojMolbYZimRDr/zU5lcagzL/pG8coRRGoJ19HUpQUKiMYGLafXfu
O6BzNZv+aGC3hU72WQqMBdiuTE109HS+tWDo4XcrloxqOh7npe/SyLmMw2UhLUvcQ80SzZuN4OAG
hpITbthjH0O4ZJoiFP1P+BK/jlhTZUVM4b1vVMFPlOEcbnggqA6PASbRuJqGRk0Q7eurfa1fXdx8
EhTHjBiykAvVRxf7/BpsFNuiYtZBxHkuHQ/Ooc6SzGQcUdIM30GxV4B7Sm7CyTw+D+C0W6RUk946
jnjqty7z3bxOA2sS4JkbebN2dYlKLBGKmDKSkSV5pynbPy4axie97JtzRGx2k/dB4lI1Zdi+ugQ1
Rix2/4W9h5bE0DETjSMOF2+BW3Cu1N9jpCgMUMmm7NdZ6C5xBDt820ONVAxbD0e2G9y7V4r4TUY0
t3A9yesMBlDcJvu2CMEhnV2bbVXVsMZczxDE3YIIEae5Js3kFDRjOcv67oLb6jkOnp73wydkh1uq
dQPVA8O8999W7y98LsNHDCDi9uNzBax05cK5afzwEcHNoZf/u43+zgg4pE1X7pfBn8eSCmPI4Fc0
VWjQ/G23Cm1L18oL9/xGgODCikbdvC8qEQvJSQCEfkusHO9D2th2Vweu1SJFE7y94gws0xd/Tz3Q
eaoxb28cCEk5Np1LK9leOSF8OxuDvAekJ77oZEQ8r0HjMkVRuatQdPVlJfjUHXnB+/3760glI9al
zXhdTMdZWPZO+e6pvoG3mhaxyNGyXTUJxtG2QjCOrprsYzeRSuzTW2ZXnvZuVD6cL+gI+hBEgfIB
TXH2co+Ode4oElOffeR2NknRRz5iGug9Yyhx5yy0O7Bv1qhkd+eOLdrgsDrc7iOLIbRkYBxTmVIV
BiJcJ3AVnoMsyw0qjSH3pqzdvKXCleFqvKtBaR8YqfqP0jlliUg0rL4NP54DyzqxJ+KmzL1xf73c
w9/iZvCPkyhx0/QB4fd1Ddl20iuF8MvL8/hVJ/PIZwnVrLO5UtWZt/qhc1ohVXPavQzjq0fDRNN5
DFuU7Hy3EHwmk9BFQtK9WH7A0lF4bURPX+xjqgk0TbkC64nrHE0i07Kkr5l2zhiohqFI2vIvkeOv
nG2t2O78+c/0b2sOFkKj6unfGsgaClbtYTNRbP20rAujnwIIsy0a1qQpPbEb9IMjQ3oMUeFkh6TH
9KBgTFGcB0NvOj57jV9VMQMgJQK4FLmc0jllaROSzSdDJwx9RmosgmJ1h2xHpETfOfMy+p+wOuH9
ehovp+wVfvtmZ73dmdfy6wj3eZ4EGVSw9cOYTrAtiJBdgqFEVRxdpgZoKiKBtvThKGc/2TAn5Lbm
ivZVM4cTzECMDTsrVHpf+GAq2tUfGfJXHWXojszh+g4p/sgrr156YvdjlXZYunAyiAAkO7es+RsY
uX6I7G/F6tN8esYHiRvFbsLMHd4IRFkzecg178jvSb8swPgWn8S+8nOPQHlovN2vDIwCt9sIRnqE
J6g/d5hrHx2htdkpzFl2YM7jiABS2SQ9h/uWFaqm6QtfOkhyK2MqjZk1Z6eIzUtLkAlmC8BhJwqe
hHDjwEQifCMvMIxFnpDSoKxeRR+nvrt9XdxRxlrygaU3jesXzNw4XbdlJtRFtKr1yJ3PXucFYbTx
ofjrt7/ZNP3EEOAlT+avXJt6H1PfZYy9/ZEN/nbDLJ3Cz/jZaNzT3MTnGpfJa9ZovzEpbFvm2XWl
YM4omLcrhEhfDCps3aCRcSqR0P+8KDaboNtoKNsFFQAl5U0+cvUd+/jG/NMOvDzUW9bW9E1QMx6d
SEI82K2Wi4lLQjy5n70QDkzzbGGM1eMcbNzmdjZBxqbWp8+nPoZG+Efg5MNwS7T3useepiVP4yZe
hNeDLKHmgWFQEJ56UNSSqqj+m80G7EwcrEQt7LDuL9iWpEs9ZhM0LQb9rus6kEhpgcmJ491NEM+F
tIMAOLEklgIBXHRMQU2YQIpAwFFmZ6p8G51oDLadGpR0P2o1s3/xcCdM2v6I12Zg3HOVvVDjqvhY
HSJOlZ6zFDNN2+lX7y8zqgG2k3Rl/98flePu5NFYSSnrx5y/qWMeW3+1Mau2fG+5fJEzO6NIoRjS
BpIvp4kTgmRvnUxeQgCRZu/grPFbtiJrjITHXh660jz8q0r41yDbVT+Rc0s6qmMGgUOBnCtr8OtF
nUjlPZXQktdhpoBQHMxD5qgOff+XoNoImFpjm9bRiqBasRjSQ0CPU/BVhoybL1RihvlLBdvrlyXe
PMlV6U7L42Xpkw9p3DEqMkS2i23wY+CvpzPgWAVG8ewKcsBCQvisQVYIXaxMYG8/S2EATWhtzZGE
IgsqmYtlp6FuQ0FmHGH9zBRzN2Wc2Z4qWno1GQuf8DZmdlgVz4yURxJqD6tSiaocqtpGYSyTVoez
88W8nPs++w31xFoJl7G7hHhkfXlK/GEVW2Yje2bKzhZA1G2sZt22oZ9E7SH4wHYI/A10vI0oYpYi
5AR78YUXLZ/9lHSMvzTHyMYIgDllF2L0An2tT/12VqmHYV66UeK88++ldAjXoVB+R7FLHt3NvnW7
kyg+5Tuj477RYhUb+577SsvihhScZAlA+Xz++Su5leTUO+DLArhrAv5vsCWvcS1z/OJ90YdcaY3u
ijsKk0RlYwScYwVsWfBhRUnZkouokMTrKOiyKiu1GPx8l2fh9U2IoTokE843A5/dzSDvRlg73INT
8sIST5pgyMD7UAQD86wvvbohWKtPlZcuC2us6bPrkm6o6NShronBPnQsRoSnha03L3dREEORx777
VUG7BD5g6N4i0QrVN9ga4DKiuT+bAX3VVBWDh83BC28XqSqFlFyofzz1P/+CATQngdbPAu9+QJhS
E1hAVTSA9Qpai3WdXED1jVXCkmwO5TOSIZkpYI/D1KQndU8q7N60J3tXMpfqgJUW567/8CGmm15y
lHzldipdrP8/VGZS1sfmm4NScNmHiI+ad2mvEnqZ8pz3eoqrwhT6jWqdQaNujGARd5vYflWhqR5u
ytkwCPOvNoUZk2FeWhIkH3UgJM2DGba3Fa8z8EB48Ydxv4XMJ8fc7SqapYpD+zUVe7NiV1K5Q75V
FTL3dvYMXM3CDOMlH5a+zMxDwoHbWlivwoipIR79e45CgWVu3Z3cxmMtxMOu92rHe1Zk+WZt9MEt
C0v7eCwecQ1OfF7hBVCKOUVYwQfDGQUa00f45RxiKZnjwQmUHWeYkIVjtPAb8wYgQ5eKnu9v/mm4
h0iUJgce3QvtEc+H4kVlGTvRAkOzroHnmaNMoKogXz+4sE62+HCgWgv1+sSTTQFx9e9xKgs4lraz
6UDG7v0KqhQ8mU7wC6Xn6gAmU92J++pOlxq5C5dh2/bmjr/mNoV8YBxqRN1+aFDazce92V7D/6H0
jDTRfLWOcH6bW0x+98Ii6jZXQavTGn81bCQXi2KyZVviTRuIlQoXNNJWLXOBiDvtJnNTSqky6a42
phMP79cmoC6JPCyUftQ7c+pHI95WxMq8OWLtrG8TsxdCicn42YiMtGG++NEgYIZo4+v+J39bsDCY
QkTl5ZaBo3H0kfZQ8og/GM8JOLv7739oAuPi29GbwiQ7CuVhXs5t3lLERki9TFdPS9cTG9+Gjq/W
ZTm3aM1NElWbBBUmgH274Ni2afs3xARIPa5V3skFdr69TcxUuIR4SsG0aTA70RuQW/4Su5uM+fNS
dVOkhc6BqSpoohGp0nHF0ouZL3zsTt4l6xZeWQu+BGPMrnK98GvzLIrwBykpSNo2gKdfHdpZYPsj
cQ1dGTaLp7nbuXv3UfdSB8LqZSa/B0J8/LC0MzOda/PRme2qvqVOIeKI4LaEVeVXPk6wY2+yvfGB
sggYLGv/p1vIOw3jLLuqXFKQpxiVNe97FgvSg1sy0mudt9RkD36hesycwW2FG0xEy2E6rRevUEzs
Aja4K5cSMN1VmwF9QCy+rMBZHELWkRgK5PhxZ1T231TkZfz55ArlOCdYMn8731ArD9udMC5Pnpeq
Ht8f3Q8eYx0n9R/FI75kGGTk0OOIKba9hjILqGzAyzls4n0oCWxQ7qGC2ke8MpIjxGgkr/AZpj0C
/KZD4IQ8Acg/R8RyZW3jx9wo6FNos127pWjVtv+k+9u/Is5kUL4ZKWwja37hxzVoehTZL+INKwaL
6UL94nPdL4kskzuiEgs9QDg0GZRo58rCzVDuvSPcfjRQIo3fFPrnz5FLzO6nqsrL3KSMiH+b9q63
LEjInk2J42kw5TPt5thLWR/TrTQ6l3IokLAmC6WXbQEceIPMEY2V7V8Q1PQrloTnR0VLBw4DqAfE
2hM2NPvBhxeN0SJb79qAotioQVnqhETlo7z7Eg1QyIwNvnYm3UdS3HzV7PIQ2vVZFZBi4tEM4tv9
SWoT3VdkX1WrCVVUZywpYXC4GcO2sXzgmVJiQzByj2rHepZ2iCMpp6u5KJpAgrFoqj/r2w2CEWTR
Jzc+PVfvGbK4VWQcewDBlDX6npWLSVW65KWKpkcfQiaFjz/zKm8G308dP8HLuNr3oE/W4O2fXS7U
H/tTwh3y4J1HBqtjyRDIyZHBEJOvUWWD75VeAROkYdv1Bq5suancxlpFZbdAakMAVgxyPwh3056a
2CI5jmMVTy8x0xxA9jPeXgWpGZOF19ts7hCMV3BDiOVR/tqnUzvPtAnW6LNWgwWUbfEvYQjW9x6J
56vyU21Iup19N4CczmkDpMmQ2qrRnEGl2Vzr2cwwug576SJFl2vuMeCni1Q4DWLgZ6eS9fZL/Jq6
n8XGVyhVcKO69+jQDwbcdoPkZKDw1wEhOEhMCZlDCrB0r2UAF/6EbdyPBbvgWS2m41ANrDS5Pdh3
/xANACNHDswe+sILEk84eeVvgQHcZLPMBoWVEy/E9Y0PU0MVLF3+8U2l2WzFYD6eshqFZUU7q+B+
FT/UU4HthA1QTJpLy0tp3Vc+BDNgeeOflTe6j3sg60Fs15E9G4brVcqmyhOJIdix3PuFJw83H8iW
j5L/l/ZExsn9FFdWVVIe/vFW3/F2M42kWhlTslpMKWqovqNJfgkGdtr0mp+EEeILiVz1nBq54TSi
eRhWrU1r0rvY3BTzBt1SqWF4ld7kWGuw4bxoCyfx+XNfE0DUH0B1gvkQtRc/VFD3QAC837uJZc19
TBLyWSwDyYEuww/WZ7C6DtCYHE26h7WQFqbf6e1f7M50dWrS4OApbpJC8cTH6J2wb5Ma+V2/EFj5
hl1jszWwfCgean7a1tG4C9ofl05rpubYLKigOqHkkFGUBusch0bceHDq7lv1tfJCg+xz9l8jTm0b
rPUHciYo0v5WpZgnHMtCutWvSs1BPPvTmahYP3lwzsDCnCtuJnOha4BPAqKDhU2U8q0fnLwkggjv
3qpTsCoFs5DNHeIuOgQPLFfQ6Tmh0HWvn7auExHPNeZOLzr3D0f1dRYGTEeQHyDFfDskLIz5nnbe
t6tszRGeE1LgP6zvMF+6v1aAk2HSP2Y9yN9HUHvHxLtnhfYgMNj57TRgYhwLgSYa+FmbKIDa6g4M
Pz0vxXWqSseXJkVGVjewZ+BaWYO103JCyGdoH0gM0M1RnscIMPvKlxmhuiZ+I4tPiyRQwW07iRMn
GqIaYc3IJj7lVWR7FzjWrcmimnpAICszUlC8oyl7Chpn+D6/Pcn3ScPJHxvZkL5IUWKpVvEa2kYT
ZS8haKv1pXJZY4EgFd81ZpT7MTs3hj1TsYITk8o+Qt196nDPeQXwuyZY3jTVYcG8owS4XtWygqI4
PzwerXMamS2qNx0PXY4R4kwgLRuNQrnBH1hEwA2UqheamuJc2KJhi3OtUdIqdps4SyAT1agOTiEp
nhXp2Pk5LmrvK6+9sQJyHHpTxqGRrvP5ExEVDDJskbJ6v0/nPpmnWtZpn7JM1z9JmfZQOfBCQRKL
Fai0M6g0dXIP7rZNnBtv3ymYD+R1d/qG6qwnVVL0o6Jurk4r7cIRUey0llY761JNYplxFtVoBRuT
S3TknGkq16B8vIAkghVldkQ38H7RDMgy3d3pFjq+lcczHYQCyUf70wYHmm+cwtHDLIYn677hVvxJ
Gm5Fz1s65dUU/r1SXs3kLuQxfOPWfniFbN8X/HLQR4AQklBLSsvYc0Hmd2pJ0xeSMIWkFRM0WWN5
Gwn09pCrotOMJcx/CXwHpIcSLvgPMzx54BhkYYyFGCEm3nLPXZAgLCYgmVTXN7jLUdE2r1t6LsPq
4utsd/zbUwNmgIb/7kSGjd0FI9AvgexCpCkodAkv4oN5bP2PjDZP4CYM9eRlJF1bAmJ0sCeiG9sv
09bcyX5c6Enw5KHbkcFBwm+VoQz3vuDxe63XPTlylQFMXVl9VxyYMJSvz/sR+d1aSrSDIBPFM4E3
5y2REAYjWufWiP2E+t4QVHWqiwOPOZRm/l1+i2AX0t4kRXMHY9yHMD+hA872XxZKjYbcsecT7Ott
SK2DISVsc1Uc6yT4AWM8BAR/IzEwEt5ux8VH0myEfWT6RTx/iYUOTGerFL/EcDAAoU6VEJXU3Qdx
MKCGNxrvS7Y+P8cCd7L7R/wTrbVE/LYimLbnzwnLuFxJLNRsoNYzdxNA7H8spCfm6tFGtwzT5kh2
Hxtv+KHLReg83+vMb/UZhCRU+qaM8h7FeJ8eAOuwglsIioEJ/RNAth6KUWLCgW3lKG3+mhEb6vcU
Uqic+tnY+uYf8ov0E/CX1s0iz5F2kPmqsWlXhWdpzDeJ0OQdsg/qSXtR4bBbQCYJsbwrPYYj9ovF
D/H55mrcgnLX4KVzrECFyOMPs+dxdJD99cGs8UN/+vftGvMdfhiKe2bIPUlF9Y+KOo9jflhreznE
SnSkgUDVdvJvxXt2OVSFIfff7xtfaSoP1RnF4D0jlmY+x2CE39EnoAtA9tXVYT8lO2WAnApqI5Pg
DkQ2vhnKB5Qj0diUYdyUu5Wkk9ZquY6VyBmKRwWyqAX58JZZyVoEUOaFqvTSKC9Acbt3CqInTpy5
e0bmmOkdS27Qo5QOgJzMd+5LGZN6batEReDgQM1TkDK7qJFKgjD1k89LRoljQoSY3hnHFar3Zk4A
A3E3lwwodWliCuv5MN1gx1UINItsgmpyuQy6KxG3ICQBmPUs1RA3FfKbG4jy7GQR1802lEvnp1se
hHMAb/POU5yao2Zu03AWhLqLn8GmumBnai1N8ksPImeeqQabPOHtsf28Rbt+nztVxqtoEg3HoWgd
DSgk/GpxbjS4Zn+N/jQAPodaUK5L938oZmz9w/f03wzb/S1P3vny00F0/9KtcIrBrtRsQeS47G8b
joSBsBCIjgCwg1kvoQ0idmgieGx76qV7jPQKxImspmoF4t2Xhay6SokMUcgJ/U6PqALClOx5sad3
cEKbJZKZp82wamqrPjT92+QYD73kE0DNj8Ei1CO8RmcC5bl40AWoBnNST7wAMyuX5YFgsuIeblxF
PkDdtlw9oT5j7xSrIneL9e4JlZXlLlzG9c9u2JjXEqXJfb1YHfPed64lv0NKsS9ZxSRnPGtjCzZn
/wFx4VGW12WbYdaroCeq5TXeuxj8k6trFxF+Cw18kGalP4AdpmEeCWbYJffwasyxQFRjlaQkldk0
dTAzDW09asvXZYGrKD5xdZrYKbVPNjKFhsoR9NQJxoRznSQlCoZAbsaHcIGW2JMqRYwQQaFRq7Z3
xhrJQoeVuUY91U03TiduUrJ1vaADFlRBsG2erkerVtgiYGK2yi+yDWh3C5p5HekPV0czV1pq1zCV
ZDMIplAdcwU16az81tMPf+J002F0RstbJ5z7Pzt85vZZ0PPt1oo/zkqzrsoPnNWFR0R+hVXjlobK
i8w367y2DVi4XIf/WgJVYlU5ZjfD5Kk1uftpX/BMHisA3g9pCxrXkYz2k3501GoNU2NGh/e7QR1d
Ps5+575DX+twtX9QcIHPwh9UQkgCpCe5F1svs/YqH7N+OV5TZYh2b16pxKTxO1rh1L+iq+LhyaR8
T0M7I2fYtgBXl7ria7JQvNWSI+gvcTcoGYgGU1FWGCigzr/yX+tLrIsIoLhRKpYl6Xz+3bGlj8Tl
hcrsrADGeHGIlwUaUnSjEppQoY4PpDR7Xol0hXHtNfrA9AAcoZgRDUBf7X4a3b1YSnX6eih756rV
Q1oMDzzjxQZh+ShRQ6RFrij+i4vrEFetB25ev2bwu9miZLlqi7rxaMEhjamR545rr+f+lC+hjwV5
T/X3VFfAgH4q6izwTSZ8SE2EnjaLcOnaBRvTt9xeC0o6My+yU5Uw/j/jvZYEp/O0TQWTFWTj/oSe
Ct05n7Jb7yiJG0XlkW1MbGLKY2VHpAqHpBs9v5zEN/daCejh9EoQ+8zRp2sJwZkZg4l5EFMMkJJp
sqwwUMqTWs+2jFVduDzrlIEcbIC3YZLAoJGI6NYJx0hHHk9TK8LfgQFdtYoLeWABar7DrVY644vB
lZIQhx2Q59y0CnjsrrS8pgTckrYg8uQgSCuEB3v9d5zdMpEmW1+0r1ASsL5PGil6N2ktZ/7TRufy
FGiwddfIJf3BLxx6LVmBGwkVLd4UwCrMojFvCiJeq8iS+qfquE6GL3EZg7Oz+Y+sNOoGUx7+fNVG
8NT4tDbjBbUSho2kiDWkBQ3zg4VOFAqQrfH8LKPgxLM17m19sU2NT1ZiVmVa4suMKc5iN/CLdJQQ
5wEW3bvpCKqO/o06oRtN8P8fzHvIULDwMMxSKRaw7MpNYtPjj1B/rDBX1AdC7unGkZnR+L3vyV/g
7aFfNkvgEEckDUui9ikkS3A3VthcvAOfkIPafCLRa1ROo/zuB1TYgYzIRFobIhjbnzBTWxXyXlnW
PHkB6fGikOVe/nMi7T/USL0+/J2z7dhueclh8DZdZALF6KJ8ymzpHoOyF3JvKqdRnHhenOS4kkNo
Dpt72FkiyhPAZLJcUzUwzn1g7PBsQqKRrQdnhoebAqGgHIiN3CrVaWaSlDAH3GuLSmPOFlLaP0T2
fh71rQWTLO1rBOV56YoEIvWVayE/pOcMt/5Emfd9i9Jzt6mfNQlLEJXhhmgz4YcP7U7oFbWRuOGO
u6e6ltntwX9B7r3Cj8xtvZ4CvHyErtu6OSZwUW1BN8vNs2T12nm9ul20aXA6wWfA8XY+bqYhqpa1
WurNvT4hhDNmDl/Qcbx0jzLhWmgvMHJLBO0bR0iaP8E6cpggavol211s7A1G8Hzp9hQ3kfo7ATTM
2ZuT6Q+lRkk/ClKIX5MpqI1O0/jQfzgRs22f4tZU04DoEgoAvgRLdZPZ3uwgPBWEq5qC8jMnIjpq
scElutuhOJDInyJZ+Q/SwQhRSEiuarCNusN3ixGGJK5KXhUAdW4BpRbRPFjx9+Y+CzG3vBGnaHRi
nM6nyX+UCLiQzaNQnmIYtsxh3dzAWUXU6r6BrhLmn0gA12cAAeoQ9W5d35+HQAfDFRxslqpGJIAv
ATeHN6zkGsPVvE6h9Sk87V0ZHHwwAP7mHBrl8AFw3pbzE8qTLuIJjngyyIIUDD91nB40NWFB66F7
TP0HDjunUZIxvLq13gqLaivfQFiteSfx8C2BMAPWroQlHO4zmWGS80HXdLi94dhVH+urw2xfdYma
xsN1FFIMMLpOqlpq/JtIyCORC2u1viEi56QjiZCJYzZqsCr8BU0+PY52QmysUTXGt+EYUP9xjRpe
CQQ2nXgGqwm0ogn3mD6ygoKdy830XtzBrNAtVGa+dypE/Weu2xSP1o6IMJGtAebOUpoVKzWs8wZo
8GBIq4Qsh7h6EiuuBNlnrYfTP3ylAJk4j/z/QBPe5zc7xJPktTWgId+i0NTAJNcGp3PgqT8YDJoa
qmOSYbhgEyY0BKM27XfVOo0mjxEARxU1oVYlXeGb2SC3QGMRi2K/L0NG1SElTy4oHmTdhWSC1M+a
4DZ2C5mp1BGrHxLzPHy2r2G3oyT0arN0OJMzU01ghyXYdQ+Pyk/0Of/tighcM5FLG64mTIYiJ/S1
j2vSLsYw/MplTeCT7mCob7hsnUR5kkq6rGZDViswz2CPwlylLz/cb0orOPqCp8lLUS8J2Ubmtmls
8fNH21Tzh0zakk4Olo5corP1nD2/d2BDOapY6AEA993vI8sRTbF/zutacESrdXQTYg8XrHl++OMR
pTOeiQ0rRikV1uMkNqCjlixm6Zm4mmBQHzK5kZmiUHEut8e4LJFC589txbRUDcA4tGY5r98XEzha
xxL5sg11WsI1tPNYjk6z2NsV4bKWJFvcjyTYYEkwn4Rkaon3S7mGz2V6Vi14J8cK7flN/fl4GAD2
jqIN+WqwCNTyJJcks+S8GaZsAVDIQpX9ZJ8crbZw9QH3TeywPXU4Oge+1dt5HGuqABsndXgXVYnN
bTPYJFWQ7iEm5vRfJrIwZtImCVg17K84DoV6NgBo7CguFYLe7NGJMquehJXSE5L//d3whbMvTA2h
91yKSat01ULw+D+VRrtOurLxAQyojZMNB/UnJ63xGdmtMPVxq/4DlL5m+QqThq7yqhDjYwAqajdy
ceqx6qTv0n3LdL0QXyHg6az5SJKPVONQiv29IGveAT4nN6eMHg3ljjnmSkVH1hiwPb0ZGIuBnbX7
1VowIdnGVveVuZXrSGmXy4W8GRCx57ENf04oWvqzSlKZ/cym48alJKfiKld1B92egAKkpRK+UvgK
ymEHNrxmdkO6vohubpVTW9tO0X05RqN2cRc3l1Qun+2WVIAdRiFzCYL6KrZWeHpVtl0OFfjr0hsK
eQJMFowBX4+AG7J6QFomtcARUoYqvuawHgNbj7jsB4n8ieb+XY24fZFJxTFmvK5q5ahOGIsQwsmS
/QPyo5xaQCGdJkuDz/dCkUOHxbwQJDxEQApmVQQHOjKBo0r/pR5YELVENQscPmKWn2CDFsd1lObj
7qN+LjEaFFLfEqPQEMIETHCS7+BdWcETJJOsNh1Oza4xWAb5yFHht/x2OJ8Fp7uKnS5hqWjjV8fs
LvYrZPW4ImI9737VV8DlCxK7swk9jV14f/ypTuaL4VGrtmyZV81xpp83CRjIGcrqxohJLEfUiZPV
LTWKixl8hGsXoi4PvR7xpWAbwY94xKZxqO/iW3PEo/WGpXKfd/bBzYPrSXSEbNZMR99gi8PIDZem
DIEApLi6AzaZGYS/84JOtSzZgoPqkKKWZ1ajUI5XsqHuE88adkpYl2yOiyuKZklOFyz/kvCxM7Za
LTLsrJTvuCuUjeMAp0H1cfTNCL4vVj00/AgcBNKSW0Y6QOuPih78E5WSsymNJPHjN1O5VyJx8/gi
b/mewZiUFjaCkJnh3Jx9W8NN4BbsYCN2WlbWHKsxECQI9GJvL8PxerLXGa+9PiMNLlDcfy54g0Ew
SCoItyHkLP9t7XqBhBWxE09rYo1iUonbRVRXptDruzKDQpe0cfydaxSYP404RkCLHFgZ+SSJnaO3
Com/SpF6zUbb9NzbOZecqRdwNQ4ZQlF5Bk5QPjP23WBVAj9SghjlZ0/eSzC5F6D0nIpDnTuJdzUO
wC9viSOv2zj342t2gbYMCus8FktsGyIsj5uH+9q8QErp73MkLfP0DSYgcBJb7wT/j8a/qH6FXHgI
mzUpeyIw+SGcOTgBxh+GUp9PsWNnujgMmhlGSLq3EtgzaeIh6BLOyhmYQE1KjYHd7RGGhdGcWzNv
/hDdRMBfD9Y2fbXrUAyXONI0PG4DrQd2und3v0iazeG3FO/DoQZBQSRZ9l+917ffMBl3yjXd/fs/
dzhPw75NP67UrBi4/beks7vEEIeCtBGFxKJOF7ry0v8uyTwS8MTfOJT68bPJxUVWtHMJFNMLFDuk
+zTC743FGdgmICFwwNESLf0EpZKvMRqgaUDWsfpLW8JPgP5TmCzPHdT1+eEE3QIvYzBnK3wFoNCr
+azJiinhyE8YLJty2FYbtVy1MDPkK7sDX1KInOWj0+Zut0wi9EampgOAc5S8e70IUGbOWFGF5ZbA
KNlhVk35UwLkkdnT3r6lfM09B0hK2v0FnzX8YAhRKE7ZZHvekXWIV3noCMuut1pdkqM44P3crVMR
VAwur/qhAOm9vWmXuxgpP/xy/9ub1ycuFtf+jRwNUXif4VutL1vW3/+O/GzPa643FabIvne6lEJ9
JQvNmU12AUuUf9JedRywmaG9QnoyC3vpcm7Y2X05xjMduT+MSx3Lf7Un44qbWHrin3rYkPwklUUU
tbC3el7WKtepsuZoc4wkQwogyHwKBYDGMSvk7uE2lMuC5zU5Tt4M8B5Q37Crd1eRAAkRiHuAE8i2
7EEympk/k6D0fhLIcf4PfdkiV+FjGfeLUekqmBPTSMfiCnctNhFfQXqsNw+lq4x2+4bkY+ucSnub
5OThNIc7EVUvEC5geO9jMYwh324fXlQ2VtrzHejxU7vSnnSslSlGpB66qMD8CcD98c4coUnl0fB7
73RlvgwE88fjkSdTQL62GJhaUBJOMMFo04+Kpqhc99LqA7xxD5YXqnGhYVU+8fL0KQG3qrHsIg4U
X4KM3MEyzBFPmfMZtNaJTpxJdYvDK+thCt8/K61Gy1MkVmdiMDnr7CiqOhBHoAAzWzIQGLkMZsfZ
Ov6NAYbzShxozl7wsnZten4Zy7v65K9KSt///2NL+YlpT17njar/AvMPw90HxMmKRsBMG9r87OnI
zLfITCp0BMsrvh8hGJzyftQcg8+qK2cfWmttvnGd1ARPJQt/0F7rjYEf7hun5WZHnn5awbSOW0hu
fg1q1NT22rg/1T6L9HkDNcGXz3vjLbAvSGAN406ylzaJHEpWhNKEwjdQJiH/rfNmXHCfIWV+fQwG
tta8ck9deHWsWQrZUfmKsavK5E9fYJb0wmNnFMzSdLoB2Y3DFG72ksYrF9ACZXfkDEti6Yt5zRPQ
3kDIzyAw6Pp0Q7JymFAnbWy2EmAo41j9BlYbVUq6bDtTJc+6RBIxhiufCK6yBk+7BmKZkxrpxZ8M
qjUvIZsdPvVHoa+cxbo9Iw+9g+jUWgHKO9DG2zRmCKJhmd8hAQb3Bf5hSWrGMs5jkq+A5Jdvj1i0
0H1HJZsKFVMW1iKvRWIxAP+hD1zB5X1e5tu2gvCIl0mczQjqrFT+zg3OuRgp1W8pawJp4WrvYDrY
jMRCXAc/EddaoLu9lBSDt9hlwCkW2VJwlWOIi9Yox3FFqkBFtpiuwVCufBjGcyJ4Y7nY1lh2RQ4B
RfosiKTyFZ7M5y9pnqz0yjRwFLe1fdH2zPg39EICZT5Og+jchHgIO6WVCPcZr2Zj7ERTMHWE6BBt
QYMXe5liwrq2eCCSNCIZSznGwanxs3RdTIMuKr4tRoPUiLM92AHm531X+X54sAKYO907NEQMNp3U
CcPsIvKQ1YIfWKgiCKrwxSIMFnwH6OWdsUfdzbzlVIWbwKOmesdMWTteJF5hxcktTp/k66+/AnYO
sICrsW5OmKa9K2fPIJ2Nvou/lv40t4jBdQSUCJioc4xSyONjj9flvB64F4CP8Ktw36FhAHtfdA+0
KIP3r52dACaBd33WsG8J8/Ue15ltJuXzISo5W9VeQfQffiyWplkOKb7HDyvCpQf8NMhEQIq6yRKL
U19t2mtwoj4CWeh562qygVv81fjDmUt6LsjC5GCzByPJAdTOltcNl//43DEEzBF7zXfbsjsgb07t
Vh0C4t2o1KG28zXGa3r7Qegjij18m+zWM9LFmVL8E3LXvmz1EHrZAOfKkyp3Ud7xhmfCY5z685Qz
yngHN6QIi84+OWysmFyb1kMnqCigKK+LlksLU91ZfLhniQrnNosnxQOjOE1BvUpkN89yHLdKxhSk
DE9Dv2Pgcv8CcXRDthCv6+/gVJEPAIqFl7TlXB5Oh9zZteWDl0KnadlO7XUGVJWMmCk1wOuWe8Pa
cHZ9UwHJvJ/76lXVYEcxQbvgfDAleUyRc3HOvtVV+qXQdLCgaUkwm0LwTbaOjo+Dv7+xlVKQ2LAM
gouJtG6OKZrdT6eFEtV8X48VbaLIsT6hUuncZHggOhXQeraZpNj+fhcIXI8GmdTNqx3OwEAHs4Kx
K794ekfhYFoNu5A65p7ORNSrbdhxENn6i6pOxV9V8ko/sQMHnoI18KCtu1eQnxWKGTmc+rM45shS
qpx4R2uRdkQ6Pv9H6zgL8GTiqx7pjwLd8jGFZjRdk+eiOZraGXqF1EDiTbH20EBPQNnHf5tCIvyc
IA83kUnitD25NcjkMLyQZyi0kYYkWHkExLAlV2zyGVPjFRlkkhVNfYGbpFqmsYm+UwP7C1A8l1cv
Xj1ylOJF9Dcw0oQJJHbr71RBXKrznB6jXNKkEFNN0wiZFT98gyWNYF94vkhvWAvJvoNqQaSNURJR
A+u7YzFp4w5hPWXvl7v0x3d4E19BDEtHm4gKCYmcRmkHJOIEnQrxIYEY5ibfIAU7oKO13KmZVX0k
uMylrHjPU87oKj1uhHB3Zgb3KQZPXwvrOYPTZ8Xmov+h4qu8HxdvRbNgGHEEmOjTaXOGvHymCuuU
5Q7r9jKPOSmxPiuuyPbWKt4re8WqxN/UbKJ8SE7qvNiBo9OOMAugWcUTGlE43D21ApvaAhReNcuK
HtDj5CZpngyrURuPa04TQJPPuuYW7gwLcShImNokS0HsZcY4AopLCaePWf3wt3lrIHM1uwggUKz2
82KhHlAGDCndFJDzJLItnVV3H659KsT0Lk+fyiX/rZ4ItmboNFEgKj2aVpOpqOdojaNmoVd4AnhM
kQk6MsXf2m4GHbbf3f2LcKqW1pQsVEq+okNK4FDRlJqvIMIVfM6h2SkTN7wmdD0tgsFWpN256Ckg
40yXsFjklfHi4NMT/vO0aD+OeRaC/c4d+aw0coM6/wUr3M20xIRv94JRawYfLyRfSXMnKd9SX7kD
6jUNhpPaXwsyWALPJtFQPNYk1VCWd++yYcrV6VB0LbZurIxTigotxwhTY4FsQtTL7qDG3LIjTR/g
nkvD7H3JChcd5HsMD0eMAQZYNvMT4awk4lTa/AHDZ/eSXjm4n7JfyMCnIsmmMvNbmmKK05vYpkaa
GcQ2XzGCGgu9GiVY6RMy7HmV8ypiRqnbhJNDYUapEcgCvMxmojq02AzRUitU3siAPSJaR1uE911v
vRbLsxusXa3YFo24Tfv+yq8vPQlt570eHynZ6Fqo9OfYMBcBhE5kEHTQiwu3mg30sQZI8nC4nXju
NnHs/3TIlhgOyx3WliBsuuSnf1cs9MLtigO64oPZVn7DjEXWAfrOcnAjVhmyJz1oIZEW5IJVpWh5
e/DVc3OO/411t8ATqQ2zgQ6vbUqmm9Toe/BU9pC6xM9EzLxmEnbmMWYZQrUK++tsbpnon6gCJEO7
z8QFIHREKeTk7OoErSx+0Dar272p+mS7wY68DAKP/lRrk7CQ6/gzSBuRzRNGgnkTaLN1TmWnLlyM
+gRE/CSPLhlsR6UlLjl8WEqe4ynLJHa/KLSnTWUtdibq20yRZ1ejUK7K4Hznt4VJX6XgBI566pyN
YhQJdbWjXMPEpz8+w8zbXUNQ+NNL4UFc/nXnop6U9Q7zTtZBDIVFeaL8tjyE1ksqIEddhUxm3nsb
mH88Z8syetdw+vLQO7Q5wYIy0vVIfME6MqRzBo32IampKU9DCfQu7neoCZQ8jhgtFd5m5DX40Qxw
MlGOosOw4TWAFuLIkBDgFBlqRGzldjZkLIQ+bQLM6oPtuu3Z192m2TZI6IGqqpFdNRSeOgzcJep+
UZav/zT9vZkjfA90Jm2iMHi8UMVWWxvMGFG9+ePgfMXWdkqnpq8WoogGse9ZfHLF0JpFJU8Ev+uo
fjuVFjWn5iBs2Xx525pdwXjTQqc160LOmBFuN0u0cpbK+7O6B9vZM0IoNRpyIVvIG5fiPo5/vZS3
xXU/i+CR0rZVnMif9m5svCELMEWK5EQ1zHFNN12MCqPlUfefmJ0wzvl/UX/hsUjufh502XmzDFZQ
wzcnOboZqkNZTTJuoGlKLDgC5w6iGOP19moxMUhvEfMv9P1NjkhvD5eZyhihbsQFYK7upMrXf/Om
P95fMr7dt/gkiK346vLStfm/U+ivxq9yM1nAsiP6wbpAyqwKFEvBcuDDBeZTBpxGW9gKG32fZTOw
PloZ+A7MlHaKw0ayNhsDHb8VtTekxQ1mLQLx9ni78y2Ca4ZCYrbslr9EQvWvZvtBPJ4t0KKbxXak
haO8RsPEbBHq79TD6SMGZQn9H2mqS4lJhq7b3jgiOyplfvWbuV8aRgHIu1U94hrmtpCmtN7L8Sin
JDKtbKyW6mbhpBPcqpRkvZplogd4lBhsddERsZFDRfmBOYVeatzPtNegexKclkJ0ao7X554wfP97
knGjCRkFeK76jLtLwOcLY/+7MoCpNMLFdwVbZ6/zPT9tFLRoH3dfoxCVxE6+Pd502AOMYdoE+NUq
801Uxsj4266QkTbpWT0yt+GNvva4G63T/Bs6hCVF+0bJp7SPRjYY+gzfei/rbX/g95KBjsOUM4v6
RP/GDYJQc1CQ3bjkAiKYV4lCeZWtHGip2ZDtG7kKaUNVoBeQnSTtz7hPEVJunCHgGnxaBm1/Gjxx
W/RorFvYgDSu9+x+Wm1L+mQ70DsSHE98Ff3LA45Nf5yb+1EGM7F7czQODxcmHp9nNo1Fj/Euf8uO
Wj/OITRwPq91h+/nYpSX+Nxsy1S7yUS4bQI4OCYEbVs+MPXXQwzk2w57LL4L125ki5I/yc/FYLm4
AfDvQWLWg5+nXXHdFHd6BTfYZXsfjKbIiEwF2Aq7G4/R0dM6ZyW8U4Lkn+hiCYk7kQLXZGrxhbLv
wpMt7ro1JCP6MhTKSDLiT6eHpYKNGJircon7B1nz+EuQdJ6uXSaxufw7kFaBXTNELfSMh4PIwOpL
mHoPitK6AwNWRRvuw6SPo/I+RqIiqZ8bDaWRS3gRcd21IRdlMnSuM73ZpSPsthgg8c9xkal3GumU
EPSJCHPNdUgh/GZmel0X8Z2WHen6bNgzFCO03cwUmxf1g0PQAVsS84tZhpTyJDL5xrFXnOs3HSdQ
dpxxLkNU6ehp4d+BfVzphpwtkSfi1lxLcLV8PAkiMw4Y70QcIJOwNfWwiRzGGrEjfo941FUmHCs7
EStmbY8q28C9f/Z05Y7+/6s3CsUIHvdFPy86sXqcXB1Ox2f0u2c3cUS53SJi+7oSHSNuSPaHxPMo
B2LY8FCkwTz/FolU+CIRvWqGAz53mY3oUveu9MvHIYkXxm+v/axjkW55b6eQLar1GQFa2RBcS67y
mtDhg5ksaFVntr7I+7ICm4JEo0EEB+Nz2/r+iTYa18h+HbrmwOrmip0GTOpJbKA7DgAr95bzhph2
NvihKY9GcOyNqvr1QCE1jIcQoOKGwRQ1TSi8ABtSVGh/WmcNs39r8bUltPTkzL7HaiMI3InNmZpv
lppME9fh2ezP98sGrmAkIcapP8FiwV+NHdca6DKedGw4fprPGOtD7zGn4UlXULx1TruVm1grpLTd
Y1eyake7c99/K4st593iEBmTdobC/CZoX8DwVhKcakkipNkGnccCSmQFcP/g48IgPMW+2Aeec0a0
LDtvFQoP3wbukZ/0IaQoGzDNrlsuR++9AoHtQW8BOIb9CU9+9yd8Fu1ouJuxRPtl+Y2g+T5Pk2FE
/aJ97lQnOfuytybrFnfuy9AWb34wl99r/RiIWdQHoZZAeUMYjqiMcBin3tQkGvZK5HTcbmyP0Hjj
mbEi5vEZ1LhbaYKIYzGM0r+CqlMeNf9DzAJdxJIc89R5yro4QuIybvVvinAEvZiCDC4wkttphhdv
ahrWqoBi/UjDQYjeyn2zBZd+fNRg9FgVSUksmSW9sebdpCkISh6FfvnHQbY9j+XzxOy2ttpyv+nH
2m6FoYf/wFRWaD27ytgEvah/OFGdVM9FR45w5iuFmWIcDneG8dGeW58iW31HZAgMKblbz+dmOPdv
Gy7sa3ExSFOrwrOG0PN9/hnNYFlJvkpa1rR79nUCV/BiMebWCH14AN6NHldTuoTRYzjJbjfwyF+r
S1iwaTuw9VxYffQuApL9TNsqYhZWxls6tU0lJxvBaqkGMfiM2zuav1a5zqGZUmCzlQhJiT8Fls48
pBogRgqc8vvVcOBfxsjLw3m2nm86tvivLM+T3zeqJm1dvYjUIg7GSNQAXqgW3uhskVeFSlPwGdcm
w19i28enyDju3rfHhEnk3P5ZdI+afCD00Akzs+WDiiRi+ujSFMiV89LEGPFZx2AQe7DIMbqWqCuj
YJjL79GHQ0uhFVbyplLI180B28/kPU7bD6+Y+4tKyp56WoVbLtEeZAOI7O9tXJAv1K2zITf2Jq2P
EXB43PpEdhLFMuFPwdWSf5bZZwuZAD9SED6yYx1mdJFO4gKsbe4byEmvBogRz5hHOgZhYgQIpN60
XeKdqzeKrzDgtpLMxYpmsgeO9/uy7Q5/A8Nt/xxtnDIlHRQavOs2CN7xRMJnEcQ9O7vrgctW2Bvq
SKe1L+QJsjepTgS5lKMhRVR7+EbKn21zXsQEAFGDHCQQsvpmNRlFBVtPDx/arHMAbWixdxi+sqFU
s0I8dHQ4DrVA4UV/rGALbcLCZ8ijiKuQSdMox1yXL+Vu1r5UtpI5AUpMwRuybWNaJtDsWI+nHi3U
GvzLwQyOpCmIVit9IaJT9jiQ24VJmA3n6lssZq71zy6+sATP5W0kFNI6LNhtoSdY34bg/3QgdKhS
dObnn88IOR4EqIwRzokxlBbWVXjlyrVnlyv2fruDXrtMBd3BKhvngBCuXmopNyWM8Am2FiSZo0rd
N2blKJ0LJJB7QtzfwzRCgcPolxdX5/BdinKkloYh5bpOUY638NT61Rvq70Lsh3Kg14vCeNvHq5od
ND9+pc/fP+nkzidXS/CEfTXOgu065oX76BQSLO7NTTRUHZpGW1iA2PIE8p0SApOnsSPG7Xhi1K6u
rtoZjwNtatAwS6wqVidfY1P5YP55gBHCT2YevVqzZf1xTvmUcYzyAfbhcLY1XcSr4LOmFG5XSTBl
4nIst8KHbJ3jsuRhl+CXRsurMyuXPHO5c0EOvi/k68xwkioDeYsf93Qph2bvwfO0+jX6YMcfGQ2P
0LISTkhggXhCo+sT0yPlPwMPsLpOWE7dJbjFVB6CrA7MHc4EXxM5elwb60qTxw4tGLwBd4SIGIFo
oFvmP411dLPPa41il680+xxKxWzPglOV98k6LmWJMvyPiA5N/HpXWGOas4Ke6y4sFuB+YN05evRb
9HQhnbboHyluYV9hcY1yRub06YbnI0+goenxyvHRKTqHPMz7PoRC6QW+C/z/jUP+to4KoTnRH0fn
qBcavK5yVp0FdfjLqz6fprFHrK+p0PfUQ9HEmjtfUnOhQiFMH6/+a4JLMu3ryJs/Y6Lna2xnXb3l
bor/yqnweCy9+DWlKvKrWRN9rBPoR25aF7MrtNIHEAJV+2IW9a/TbHOY8TrwnQJFj9RNa8waJaMY
JXiMwqiWeG1eY/Q0JaKlN7DMjmveksD9H0+XaUZkDuoSZvFj09aOrX5ZPa6l1q9JDAPaqiSdYi5m
5hYM4Pj1+j+ZE5sRzh8WOYsM39bi+35YZL6SFIYR8bh8+yN1G3f84O9wY4wlN/O/humgA4S0PHwA
C0b8c3d1qgVCoTxYwB9fYOAvmb0H6QTBwhKvnkdTu73dqOdjih5X8awHHR4oKt9Athp7W/63A8Lt
Y8OSMCttrpWZlfmd6B+b96YHXRy+6O+NJcVBTBgt/4uyx9xP/rkIAG1+c2FPrjEyJkOPSVeJ/Cbn
jB0pyYdOAlM9xzTHMdbuXJcZRsfKnGkiwjwa6tQM0LIRGd1Ox5sTYHuSrd+n5d6IprRnvbmvwuy+
sfjjXkl1/6bZB+ioapx5bj/J3pN/xXwnRR375yHNMPLVdMO983jrH7fh2NE7h91j4GYlRzr9hCUo
SVqsf7kVjEG9nhzbtFw2kKqfhGk4+728Nn3Mn+lxrWNMyESsyiLLOsO2Uuhvfnk8cZ77zc4ch3FO
7rcNkMBl7Rw33Xp+qxMwK1nupJUqzi86tDGDcnz4cLH7NZoBmWyA8kvwU3oDZ84Ai6zxgHY1DQHr
u8wlk64ZFz4AiUYUkoga/3NUg/6dAp11bQL/CzoWfakaM1FITwRKgVcNGd6LFUojSWni9k/XW+uW
eFe24x61Bsm9XiCDpOy2W0Cs+anKDLv1Yd1boNGgC3KSGMLjWT2Ew0kpLiB4nP9PIDMv4wZ6i3J7
jEhMBHe/hShzEVkGI3L4HvLdsPtx05FToeK0I5fUqr8bjLNyuFgqVeBfxJNW9V0jH0pCKWAJZwVL
kPRVPe8VG9tuHS6HBPgiAwv2BAC+dJyiaIAsokqGFM9HnPpQUduQMlSTQXkDvAj1n/N/izA4JbYk
W41qHpsU6bjOQaT2SuW/0AGlWPVLc1Z7DTRFIq2o5YX9EMf46V2Sreb5N+k3flI/sR/wvamsO1BD
kEln4zOa1RxxrH04Rfk6eoKimqH7Y6gX9uM+4ge0rw9ZWMlKmtZ8hJcXHvfD/9cLFfHlAhX1DPEH
VZbKMLalo8JqedNB384VM/7XDWijSGyubfXiEUGIn/ATPchWXb7ojapLLEtsmgD+Z9K0idgi0ga/
PiRdv30ah6og2g8+maXaLFm3k4SATQRGceAGNFVhXQ+/qrkcSya8S24DhHG0es4wiY+WV6g7ons5
rAuQfGxyOi+YV3Xq9chjVFyzQJKxRwFKRaez7DvmgnH5baoAOtpehpssXXjtTfnNoG1So4KPFjlr
6iegJZbw4lmJRCJdBzXEXuPKlYYWwbKWCQ4Be3JLjxJj/Bd7531azy34NyF0rmw9Hu/+nfA+pLbE
HywBVV8EKb8NmU68oOSY7nzOAdHqBgWAW+s4A7jBGenqTU0hzIT2/QNP8iMkE8scNUn1t9W7/Bwz
KG1z5c9Zp8c/ULdP3ctGqlF7j8mKzsIUgHo5wh5VgxWl40DWBcQwocQWKGq5iZgWXS+bBpHiCTaK
mtZvY7tLKFzvF84ITBrpidTAtdW4bsmAtCA2L2i2eSxDjWtgVU3Kp9W7RnFy8Fzia5U2oytDMi4Z
BwfBRx0tuOOFAaV+B40yyYBXpfoZ3rYLY5xZUyghv7swEF4T09aovyPddlz+LB9j4krpO1WYPyky
4zQHuYHGVtnNbExBMgnLQ3jLy+6lEu3VCcxU+rd6b/rQdBYTBcJu7+UhzzlFGZ/tlTfM5mTok3qf
1P5HKs5ItJVYkJv7lT2jTYEFTXWSsS2AYGid5/fitr3kihllBbW4TRUo3EhsONTRBu4+mvowkpXf
4bxcl9u2qQTA5l/pkajLY/GR/GkqHrHK96ra2MRwQcCMg/JQAimtKBRSWTMzdTtFzuBcwhTA/443
2Ug9ayNlDaN2aQHVqhR5f3Xh7xomxqSgt20yKFBXYeYqfn4k0nughPPJ+OmPR4PA2ni3/l5+ei/a
vkoczhza2PRCx6ImdieNPZ55vStWgeGhLiYEkxOgCnSHqv7Ypp/kfFq4Xn7XXvhXm3rKhNUVL2I6
/oBfpWTYhZcbSmz6O8BuZreUfF7L8157BJHoLYm30gWbPy1tYbjUtIy1Roo3Wq/Uf3oIrPsMx9NR
Q7VJC8G7u9yU4FJRVU25xll4Ffg78eYXw8lTGheImf4A5ygf2vmsjy36rB4qYBjWM4WXVpOGn5Fx
e8wVuYADqXyz8nCT6ZkUxCLmwq0sr4KEnjbTiHCVHaxNb8lvpkN4Gsngr0LUcnE9weUx7rVKhO5D
GPIc5jGI4q3ZI/MFmwDZKzLzSwVHdpWhHlx1Dm8cSAcJi43eXt3zm23rTsJdh8DwLGlEBClVQicc
YmWcAtwwMlouRTB4kqWPGV9ce5vXdu47M0dUdaZxaw6UKqPH2p2YJZsSzzNUgiRyNyGq8gGZDsRM
7So9uVoauELlcCtP93csIoiE5+t64uFDuoYLGoo6lsOQFAbB5X2ZH0Tm9oNqb5yknDNvxvmiaqNd
sobd6gI1H6l9NT4U++rSU0oFlrcOC6fg69l0M46PDmQ645ScpLfKwVba7BXfP6d3wxry5RIcQtTJ
4PkMysm7npSgnLUndEwjHBEIKZq8AnQdYsA1TOTyMIsTzYMdRIV+xjwWg7eP7rxcR/tibWk9mp4d
PS0PVodmWZc7QgeH+ErnntiioViS4WGFtERc5xl17U9dK8e3oWUeYIVdTwjEB7CZTpkuljGjidSH
Q0dXOl2ArUb8BzyIosb6lkaVu5Cwqi47UXrB43Hhd3RN7EZTGTqiSXEMolCo/uOBuryaVbtjLJyi
na82SUay+gmvdRiW7xmD6cYt8QgqcPQxEQAE9oNwjijxW1ff7e23o0IBokKXy7CgBR6dYGAOyQAO
YT3XNOwD700YIT/qpZayNjZuIjC80oEph9XqbQg6zMDW3Xm3fv0iWtrD4CTPCphvIkFX97uCwaNq
ntnNBhSfTcoeJ4MPXLfzwgUt4ZLteohl64DWJsowFilCDd0z7UNY7OdikQg2xB9GCLyCdk6l1Zp2
NtogmeH9Yvt+29yQSCOd+7CpJR/H+7b26FM29+eNx0NqnqsTVdwd0+0sbPyWe34vQrF0rklpnOq0
Wa3rn4DwNMwY0qXQw3q22ZfgJCg8laxThlHyV516a93SKs+rco5ChU1uYB7WGk5mAfOoCRVG8bUU
225a3Iw+pR5Ym2W49bfz0PpkJ4DVTJlnZACzrVKgUENqlttdwFLOgiXS3nVHzsjQgI4YDwSxmwwH
N+wSPF3NDjqyD7Y0EddvMhmAam0TFLR1aLzFfj9yqF2Mivef3/8C8XlMRztVi2WwizcQibVZHKvL
mvofBmsPW7FTcM52VernW1KOFGn01bDrwEke5a/POmiEjSCPylwL4uf+Wr74I2YBp0I7xrATt37e
64PBEOyiLShbLJejb7Fz87E5aLbe7CTGsvSRZw/mzFVzBDIn84190rVgPRPIA/Q9Xq0ykB2KG0iW
gJL+/l+pzuq6NI7yw39Tw4R2xNkETVYZ6xipECfKjPLLCQ4x2J95jWeYxtSxL3Mbq0apefWa7Nek
4xsVdBId2w9jaVDWOjZx2VcOpvwnwlzNgVd1ClzNtulMxSwaHT6BuEtxkaph39nqfvhhMfKHO/jG
hUPiq5jioJLZxRgqIw5luOw++nF4sJWH1laMAAcIA26T3hGMm40hWWcJng1AvZiiqaQ5eCZ4j5z5
WKxoDBmx5Q3N6MdwnfIHFLJsdDg8qnPl+ptBMvSqeHG6igUyCAye6uspBe+ePRfCQ1tELYBQxkR0
6ROZEO5B+TwUaEiV+ciF3ge8GR5VN4MHar37AtvDpmlI5uYoFE4VW4u6DvByyeLMKPUqVH8vbVHT
3yIHLQJLoDddIhCbQVCx/7i+Xx5YWR87xHINMu/koHhsLpeQsSvjGkDFDeQEuT68E+t91/xxhHhA
3sjeSzHOUdUIRp+SdK7GXzgf/7o67f9W70kKwOfKJIhiJ5yo2ENeQgM1wxR04K9KDsgyGsh0uoQf
NFTU6aiuk4QOvEOGknb3bbpA05W82RlMpHjj9aB+2opbU0EoHLiJnIA1holH71WvCyLJeONQnOow
hezCSs04Kim02n90CkVydLRXF7jSX7hkt17yDpPXzS1arq/xl2zcpoYCenooVPd8u1eBZ/5qVwQy
T8bRw2fnyB44+AaGjezNlRoizd0E0KzUl7asNl5LTkRKQ4nVS/49W8g5m2VrqZrKTpy0LUIxXdTf
3DIt79Gy7vDQvNKx7UnCENcA6vVjJm+W5wCrLU+oWQLTDrA+FfkbfrpRKxc+3aTskvloFYFNMl8X
hqiET++RQ5iohPPg5cioPtwfxHzFHxE3n0kK8NpMoOy2dAUdEnkoy+LKxdHkijizXlPHj5/ysU1O
0bb6VZWxneLXK9DRKBpUBoBdX+S6kZ2baMDidt9nWcpxoiODr1SldHsAU/lZlPdQ9juXUVfSq6wx
+rPkpBs+koqWZQbb7p0Qv9r0c/8oLGMe/3XnQqKCisyiBaPkUj22P7JNGskDloaYfULpDAz1MDKa
luPBPq/6pQXHvYVeMEnDiKIVDNb1ytmOp8ACE4MeuAuitcxeKxGZgIsPpbAn84JRP7U8AW0m8kSz
DPyNhuquShgrhOegf6exjPGDerBA3akAnjZ5ZEwv9QE9kE4IWRDROWHTMsfJsn3pWZcO1KKjeM51
iY23zC+jeWqTHbjnZhJmG4KHB8jN53Uj7Lxd2S1jymp84M8oN89kfeFy8Y8kjowk/cdbiejypia1
BZ5ST6NWYKqdSZOEhkfTMPQkRvgDdzbsTLWgVzMorNkb9SOTgYMp4ymXaH8lpQYnhAEPJUCho00S
FjHvfwWMGnqkUt86vyT729oPIPujCenyQ1HEsO17wCrWOOdQ9AKJIChIK3YkTqw6WLVHYDvtlU82
Ta/Vuh0GoyumOCzLFfz7IpOV9Fx2PcAqlZgTBwedI+N9g1aE2uWAW9Z42Hxcyc5BUQwdOpo8K6DO
NcPsDJfH+mpLXMxIbJR1tgbJG3/aI2af45xxisX996FHaEdyWczDkzPt1jlFyFv00Xpzt6tipy0E
Im7sBuQInK+une+cltPVgdHuGOq+LkloissQt0oyZH0wVa6aCMsubhR6UKq5HUOniU3nrLYQWlW4
INmG9AdFWiUVhxHRLruk780tk+tLa7sSamho3eckK7dnW/BKi3B2/O0CH+E5mbTkhrdc5EwBjefd
SDQHeqilEwdFVFNzsyGO3FHkKkkN0Da0Mco5HryHZaSKOlYwLzvonyRWF6zVDKN6fRD6uY9j9QO4
37W60x/xunlsSPJzi4YK5J4KEnI9FZfOBaYjv3Rg6psGXj0WQCQZpYcpJJNb7aRl9CjJTB/bgY97
XD04MWiA3lQKDj8O2vYMS/VDNWyNUZtAEcuNwvsz8hi7UtcTKSmeDddoXtEarzmG2RBNYLh+sjP8
i7xRv9xtUqwtVEHeUtO/QvaRxPsNLKVGeFSOPY1ABMzdqiXR4CTQX4dVIJzxhW4FiSxSOeJUm1t5
+PkwjikhBc8oHQyPoEYe6VoBokLbX/aS988cPF0N4Hb8G17Iu8I5jOBB9cnCeAFCrMyAWTpXDtXh
dh8Er2qtLo63nHkVj5Dy1C8cSBgqw9YTmPG6JVoxw+zqTIcn0paREW/PHrnTu/BdgNudDdp3DDhx
y02oR7MZVjWvLMuwPjlthW/BnY1NTDxZxE31f9t8J3Wlcj3x/8Pal140xXdso4UvPGCp4R8iIaLI
aXdEThW6jZF4SuawxCsb+TVjBI9BhQ4109SXk67I8gOEKDgSu/zspfb9RtSVlo9J02qE04VH7jQ3
biNc8ff5NjDqTGN6z8GomP7qZHcLGuEZfcRZVe0xeP4P42E1kbLdZby29aswgy5i2E7TwNG7UBcN
wvL7zsElPGOJY2rKsZhF51v8ZbSmyuNhkbLSzsr2nD9QXEcR5XYXdjOPRlUyIbVZOe9qPAAYP7UM
CC5DrK6SPcP78WUksrEZDSboej4dKOMAf5/5QJXzqoFySZYAdua9udIdEcpeR77Y+XzxhWoF/xyW
FNqe8t0fP2aOSdUkTfsslx1ktJtIQGV4KFitjDj2dNEzhWWRdu6j8Zts976iP1+8MJPS8CZYIhsI
ogjBPUgSj0VZUPO2DqRTDNO7PyuaPaZT27XhXCXkvKPj/4T/tyvO5XlTfW+uSPX+zJH1WijGi2TF
eP6jUvCm0/p0n+P7nWENzxlRFs3awC3sFCWXiRwKH2z+Pku4sxshFFQsqr5sElrFOtvWuVw2B1i2
y+FuNAhXhzP4oV9v1WJtLQ8uv/FyIWRI572mZvWd2K5UoYLceYWaf9OM9PnWMrnlhcJJ2iXydaZC
KUQfP29IpMdRgrrxnpn8AbbmARX9vmCVspNAv3j6fSOYJdrMeaw2Hh9WCNhbGSHeig8P/eVesibI
CzGN9f3+Rs8ZKOR9CFH37zzpc8aojXbQsOwbKs6AHkLqQxfvcFKcUuEHYBvtAbpoJiYFMBIEPN5k
6jhbGo8+z5Bw3Xo7aT7u2D49bxqZa79Kvt8ofWClR5xehSZcfCsu65TANfJP6WW0iERBvMEywY+x
YQXBH+SL6VUBqbck3pyJnco0r1TmJF4GlIdSmcIOrjcLMk4xBeYvh2WOlwwUl7KnHGGCGe401f3A
9BuopKxPEf76TshssJxmq7KxilxZhM5wqfjT4UgiktIGMpFCUhfjofSpTi+UErjqAYI11+XiT/NY
PQDaxTqJmLj13DDpcYnMCUey8F5YMRggDBja78FISxgLA/7cMFMqU9harNc0dMw/asoy5DnMMJXA
MHd31blivzAkFGb68SFnqrZyVpBLrg6mz44gW7I3c6BP+4iS/kWDvEYBXremddXG61TC7nxb/p8M
cAYob0aGbax6x+CfUWmRePP4BlvCpQMNjDuUkPhEcPMy1jNVvSMioJTxhOsGC0Ve0AhI+0AMwFOa
MOEdxcyB9oHbV/Nx33ZHIJEbqXiyYPPxZDzFyfj3KsEkjT6VetTXaV3XUCXbRhqpqA85llLJtt+l
YY0X/XAJTk7bLwNnA9XuCai2NP31OBT13rm958FLqgwOuvkQkGpPUKZNR/VvOCJ+o+//0HUirZ9E
f/jTH8mO4xtScRLzDkaDFDTDfJrGSAXzbfh74BY8b4sLbItd2Otqhv+qU0+ksj6sqjfbphlrp1TV
sgd8gbFipdrYbFnOLlr0Q/YGK+pzyBdmJGIf/+c1c+DoqnDDqcr4fiu/ce288wJfK2jreGdurgA8
oklzahRN1HlB3OzTSyntImoo9ggkSWrlH3qVbSeYlfxV0b/jeayLGww0VDy9XQMwqX7sh0n0PTR5
g2N/XoMZPpzdpUW3acmo7mFJVa02kXxVLXjfHQfwSAVVMoIrLrihFXSyQXlSK+c9A9wits82Vh8O
vLwcY3xS6UJKAEYlmYgvGvYG9fVIPcpsIghL4D2559hdvvTE6HnIlqcLeIi6Kk2K1gAWOTgBa3oI
eNkberNc/5H6784xGRKFW7K9PsP2RXK59YAcXS+VvI3zOpZr/ijbKZ7cM766h7X2uj3pto7EMcd1
cm/mmrCvLmo2AfCTms0y42oIA1LeemyWfc0llUNaCv09DzuvgxHiI+XCAzAS2hacVeyyiFO5Euk+
V8SWHy73VpZTtuTA5uSO44yA6OMl0zXNzD+ahWNMhSnnHBoQbi/ElR0mR/wZanU2vSZDBv15GGz9
qYp+HpnEN5b2V486qerh00qWpRhoxFhAhddG68979d+FSPgYmNsnyLZUDXp8IAjiUNALd/K2r8uY
mL+ki7nBWXBeiSvjMoXcVEHeMVGi/Q0WU916WNltRYM7apP5gIRQsAt/9WpUKcMrsxGVHKFN7eY5
kEhyPA3fhXeVIpC7/FX3LJLGzHQwM2aLw+vAyKtkVeXyxEIGm1X7Aum7n75GKELUL9hks7QWXuvp
Ug7Rdzxof3fo7TdbLL6kWWYnOM5+xw38/eqtpjOrmDnwJiFWYg7fJQ3wY37Mh0o5gTFvEHDHwb2A
rTqR/6V2uitWCS6s8gUNPPGqmuBpcOFdVtSNjAOPQuDTq5i5UEpZqGwNqVqAJyiJCLxZuCJ841HE
kKI9FByKC2dNA6SrxzAtpysI2bmjZKGdOWrYZHt8Mo9dm80IOBxDeCkUOtV9VhuC8l7fLms62T8C
gl4/wisk3fck2Lers2eFNjThw2GsBXYaGnaDfulDzQ07mpk2AWurkc1OZlPYoVYDaoiFWwylZyGS
FomPPKz7E0GahANRFlb9wZQfwOp+D6NwP/J9ZuJYAS5NhuxawdxyUFgSQu0+Q2kmzjkJj1ULzGp7
cGSHT4qj3dX+OL8ErhXd7EtKaykrKPgNYeDQO5epDWATt7wnc/Kz6ZlRze0JWVw5CKStQBLMQk4w
WCVNMVO3C93iCvO1g+42maqPDLf/da6jGtOT+Edy9sb8NuaiKVn0dbuBD3mE30Ns0YrY5O+tLNqg
nHPQgX9Dfr8jINnhnMiu9g5tFL8oeV4v/ELz/73el/Q/nA3rvoJCOwfS1gvdhyjNJDQbzebuQSMh
4o/XQDDEUgtr89KTBTWjrDRnQoS/KjJQWtN17ZtzEASmrE7R5j+mZu6BWwRZm/wFWaiyE3QFCI2C
ygTrMErt5WBb2pKVCeNZ6/iElCP+v1Knt5uR4yG3yxaugcQbYbRC+L4ZsJXtfu0pUa6vTxX16gWR
FwownRbbjpHJ8PsADb+OhU7Co/8FX43z/XMxK1NtPgfj6oV66Ik5Ap4LBkrZF8tjTJ2UGeN/xqaz
rZ5l6pKrIuxOL8+mXdt+RstbYWpldoKBvnXlAjR7a1gAY0hqme3RFijqYCdyjxDvJZmED6qgXsEx
KD7i+x1LstjvhTiQhCrA/wovyWwXy60zO5jVgzcE1L9bYqvhST01VNZV8r2Y/LmwX6K8b0IQXCAS
xn+M5Ad17NCzcjI/b4QLev9+Fg2mpnN7EmWxRMwxAygJOG2+qZfhEXIsdK1coIZ3mXtI7dh5EzoT
FxkheiIDHo7kJ9CMxDoIN9R9S4qIaMDfAdL43rGQy0pJx6thxFNhUdbDS3RUM0xDl4m/mv2buaxr
EvMSjrMJKCBvuZXGrYQ04a71rnI+zrSkrZrsKZz+hH2lplZfusu5LdC8MGYIZufCMZvuqOrHKltO
k6Y5t0AM6bG0GW3OR5K/hD2jUAxv44WcFwDl0EdqFKAG6xQyrnx/8S6QVaZQuXt3RUoRpFLACaP9
G4cuYTAwxtii8xRE/qq5049qDec5s4WpC1l5NWnWOlkE3pIeQCHZIjIlZLoR/ROR/C4BRvVfOEN0
1wPRx2ZcqeG6w3+Jy3Wfy0UVg+LX+uhkTTxnL1oV5iAQGOJo0LwDAX4Ire2qN+qj1KkXGpAzEFAJ
uaZsYmS86g0owvkOtJ9sYryGO1N22HLVn8V3udNvRlhVVyMpojgq0caG3MkrHo3jKN+k/Qmzz031
Q7i1tpTuYsiDNjCWbs6t96hgNz9vWOX8OYQLK5DuCd260qLOdvpmpmiwPpf8p6nkA63vLiCFPlKa
pCt60IYVKRWLvwg2VakzUqIO4Gy0izLTywKVSORGNCUvvMvDbta5yWkdbEYZLhsSx8OqjyulN5cl
t9KzZhI6P0Q9HuM2tUF+i5CT0LEdAevORi5QLiglBDrNReYh9cJhzslTnSxCBW/ayrrW8vrAIcv8
c5zc659iHq0kZ0nX50pcEoRJSxma0//IZ2Dy9Uzs1imJYjY9nadvLZXoBUpdd2h0zJu3+U+BtGeM
uzRkCpu1IBAGE2UxsM+BPR7ThBOImVDPu+3iNlmNxR/cup5pcc2UNmN7vMe8kADuThb+3DQizUvi
xCqDNcEbQkfAS3N0y+C6jFqIAcVmoZ9gVpmG1e8N+CdDgIx8iOt3zkyw6QVeXsxVMzwboeSjMXdG
cYOTrlo27w0/XwoXKdlKKNEUw8sXcR6yyxH5l1uybARQtsVR+jF7nlcp8Sdvtkb+BE67nQCWFrUK
hayoITNm7oAkyoVriDgMKfagjtpPWH/MbL1HJFi5laEhEDuM1qnz+tHWa8b8qi6nf2vU54DhT4mq
LkY+VdRzJEqTs+6qm4BLkk79AUaYes9Jlk7xXc2g5eFiBOXWsHqwajiB8CKlN1EShRzO7LKKrW5a
RbuTsPeRkmcn4jNCpVzWjwTen8V2V3hAxcRdyXQVnvZZ5YQIm49o5/AkzIQD/m06aG+OCODoDfT6
MjycFVxmTBAndYoWdNfu0fjoP3LkwXc5fzjIbYR+FAJWsP4pywMLCbIk9J0NqXY08lra7zcthWz9
Wq5ympcPFfJOhSPcxtGDZo7GinBUVSUpmqOS8S0T5qs1BtAQzT8h/bCX1D5mIRaRUP0EMhYyRMWe
doyfa8VEdaoLi2jRm0IZhWMRlqipHnG/ypa5mijuVi2fwpYMMdT9WleJ/YcHimA7ShEhizMlVx44
uM66m4rDavGeIbp6ozJJ5Go9TkOrftQzvaHQvF1Jw4qAyHMW4tRbML+ICaK5+cvfupuoMj7e7orF
NWKaF58oTxTnGv08QwpcVIphE1BjQrK2OlgipybPElKCcgSncGffHDCdxxOyagdily4TLtXmX1O0
0EkacG7ReNYkmH1DqoaI8TnC+Usk0yjWDa4J8/ccJYpgu9YeYgaDkvG8WyEAZzZr97A2i0mKYr1A
XLbTpo57Q3dxleLFKwILdNJZJlkGm/cEQEiw84AHSga8xgNQ9Ie0R9vrs6Km2hrspKjipkF3nPNC
7IbfOLyVnvkP38UqNhRHS+zYAVKVpS0/JQY6I0qyAnkGcI5n8h3c6y5WhkSnkyHGO8Hm3WOnFc7m
MOBydtitPpUg4xfJLDXKvez78gAvX/nWjN0c6171fVeZwwK53RzXATwwRzZSQZ5I3KQTFjk2E0nz
GZQALdC6XaMSgux9g0yMN72AhKNQfB0V7t746zs4hdGYmJ+SR4HV+AXT8GPqqpTVXCbGMPfiEvAP
0hEt3qH0rlh/ffKsbMiOwXzCbNlGTSYqBzyKZG/oAWpP5cGEoGr6qQw9Fe1tnc9XND8w5xbyVT3P
b2gN92a5h1vQoCj5Lzo2hyI5KwUb6umXg7L05EyThFaJSc+hr7b2znRqJVXHh0gO9asjGBopLwWx
/yx2sqiEZmNpXpFxyJC+oWYOsylDhBWoROjEnsbGMu2BPUxSwFDNc0dZYJ5wN9sZX4YFwRA6OtuN
t+bjSxuuh1hzCLSUgX8imC5ulCTyPaVWQVhrvGjIzfxe8N1VVjHgoL9RMtyt7WFaSXsNTOjI5xbk
GJZTt7oOCn+RU7sMqJ8/blu4H3srmT90M7lcC2XV9wYsOiLsbtT+4hQoR8OzcENx040dATC2uGqJ
3dYtKVyfxx3RSZTjDal3e+MB2MEIJM42BSZ+HPGKZ62wPMEouN8/Ic5ScExVRqIsxprQNMsGbFtn
r2HuV+yJiZrTmygVyT1qH2ikQ3Cf5yuBgZ2mBXkyDXmO+T6w/eZm0W2NgS5BKolu7ZIugesvlXki
bpezbns0HaEJvioN9ls5ZPdWPKFwJwJcyCwetdhtveaYPTdqy7tixqXReNMq86VYKKa4vk42TY4W
rojHSs5zGbr501RMYQqRo0vhENWxp5cVbrJPV+kXw0f8DdbKhR+PhtbdEjPEbMpsgdiDAA5OOEpf
V/50Qy4ovTbXsxR0TSSTNvIYrmeVq7kz/yJFK3vJDkxBTm3ZrLyxiEjvjFQedUbktgSNXG/2q35Z
9xUA9FVeISVtc5pZXXhLHJjLpG6K/lyjSoPNbJIvwan6FpowCVcYHzXhn99KirK6g2jDRITtfMlY
Ai7wrWXe9k0hXsLBKRwbfsc5LVxLhLsaKlHYsnvYOCPa4MSruDmehO++4DKyoaEPx1rS1B6ylS5t
QmOSbGERFlOGK2OaVWZpi/aV9fDVmkfhLr9qA0WMyYKyuFEaPBw4/JMzJSMhwBKDwfIlVuhkvdj3
mPhZHPUsn94584lCXBpm8wRWvAnE5ULqpJZE+eO6SUvN6tq4p6hhtLOz3wAx6qwde6uF1JSDmKJ1
PxoL7GRK0IElyyaX1Gs+5iQbKdWrNMW7G1ussibIrCi49gU/UzO/u9SlS25/nNO6KEHqr2eqhGx5
/mH7K+N3f/aGEcogA+mFHqXDUXxSJ6qtV7r+yAAKhKJoVXtcyKOOQDotf+sY+8R/d9qOxBgcP1ae
2tmwO5n4Iy1GYJM4/Ad0sfjqybNrZOB6dsLpOwenqlxbkZGX0O4rlDJpZZF53Hl0fe7Vl6+LWNUG
GviiJm5MGtXprQRjTRFwGHHaXciiZ5yA9xZ+3paYTCFoAVC/sAlqPImLZMQF1u6Frr3XAhgHYFI/
SEpfTUnv/wCUKli3OHOwRj0w++HifASHBINzR4qONd+Hxk1I5KhdNu58ceaqGDQmeXiLzkcFmLy0
O5dZQX1vQBggHt9KxcAFmJ/JgPSEGPKrevNQ7GDflWpT3Mw5l9qfMhVx23JYP38RHx5iU+2hJPgc
YE2zUDJBtl/Hy2jZ2WCf30G1iwF+eYOBZLb5m7Gy46oLbB6+iUn3vQqCHf5Lc00DtTpFs3bc6iPI
cE6FkNrcFgcrqQVaVYN4uRJ/igSfU839pLOFLymPTq8r5U2dkvmsSt+SLwGxQznr25Sf+uNa0Qr1
YSjZagQ2OXS7D+Q+7Hy25+hoYQviGUG8noUMVuSQmRWO8hzlMV+dsKd42OsX5qXGsg6BXWxdvMfT
lUILp45lLgp1XozW6X7y+ERe+mFZ/USfKlkO6ma8seQXQr0MrpJyfdmJgnlCKfVoVAQiXSh7+sCy
FMn+n3CiP7RY1FvOKgJ4vsV5FcwGKvePyw40c6l/eFAUjwXkFPNWzJLD1mF3Oo/5c4wqrUia5wPh
FcprGb+4cbOxOTAkoQ1sMUeKHFUJj7xC4QX8BGb+Gr/2OHJr9Y3/9hCcKAw5A9Rz3Igeaqm9Pt/t
7zrvcY0jWE0iDohzZE8fv9CW7L3U/yrSKY4h2szwOFUA+9ES5nV7kKGm+hTPkRtDYwu9Lj+VJfos
6HJK0KPI9qmn6xbXDkEap3Sgvnjtm5KgDT7A1bCwonwqXx44sIg86qAmBJzavZLe7yfDGn+5L+el
oQo1jU0tayM/6fB06oFIBZkAQ/CS78YL3XHzNIz070ojrRP6BK9pObqnCzVPSTOxcHfEpu2MUkTm
1h3l9AzqhYvUeQFIOr3/D1qj7mN82VFjU3AtRaAqJrlttGBu46cmrDBBNW63D56DcMEg0ai9cmxM
wUp0E8TS3xkxFyibYerXtdIm4TVKZDpZw2HCPSOG55a4dUwqp7zqYDul1ZmAjgYUs5Ye59lEgUhD
1VwHxRxCsGO5Y9UuYG02PKamNLYIKWajhcngpNTXXVDnUdY69OcQfPoePRW1DB9EUePjN55VgTP+
kY+GcFxeA8dN3z16LfKPCfXpwEjZ+H25ZNbvNi4AnbxsmEPvVu675gHAPCnuXVcerhznFdU0nkx3
tH+Ujvns7gtcNeZWp7tEXBoulP9psdpexoVf+ShAVKTgScKGgh6lsWGYs8AfqJ5sPExz2flhHSbf
WA7AGM5kPaL6tzT2M8pnzNlRowp2IqtPqrLKjWjfeDmyXJ8eD0p06Bs+kWsn+Cm5nOWYPdVHoRNH
OCdELzSxWil6IajuTHWqZgkVH1HsIWLlAvvhyFSDdVhjfj+ohuYiWU6vSbauMiRpT7WFtx/sCtHv
9xgzJuIUpvneYT7Gb+YXT6ImJNP8XcSxgO+VKgrNflgZdChpSB2EjcAAhMm7MJVpf7cgyCHxos23
SRKKzMv9QSR4HXrRermZA8iCjC/+EKDyEKPTOQ2m1oSddC4pn0W0Fr4VUFcOGjyGFFz+1+dj8fQ7
f4A9CZoodzIHgoX395jns8C0GOXL97z+a3fFOl/JlDa53EDd9R6pFDGI/O5GnSRykEVKbPBS2Kf7
sLkDgHoHVnEns+Pd4Hx7cRC1xAUwrJaxiX1SjDV1faNOG7i6kz3C7ZvKD67iECSV9GK3UeP58RrI
wpr3gWKvGVAwJh/CiuYVq5HvHuPjpXRrf5jvkM8PqcvHmmPk/2CnYM3zYXJM/LzqtYxF8JILqI7j
MwTXQpuluoACEq9gy+M1Elka3l/mT+4PaRKKeDtmdTu7ZAvkzeJ3gArw097hqWNQWI5DB2hGVpk+
/eHZSnvASRUfHYB9RqlU8HaXFJ/tCKYL4fAtAzvt4M1MkbKSRpYRlWeXJCReBtn5Sp/DSdeqBZ7X
po72R/kAbm6x0V19ZEXhn6bmjjWbn/Lo7vuhE/o0/OOf6bAy0M69LGcmY6khNiaeHuERwf1yH3T/
tOhn68DIEEyN49l4UlpwKL9o2s0ml5gpB3kf0ldN+pErF2pb3GHSXbG/SNpSPdYVMks2b3XnempA
fOKipMSaHC+cmuAxAshH5nyoIIlAMgSu9CAtPmC7Kc0sJ0ITuniZFpbAKROyQ19EmLmmjpjk4evH
DYkhYq7nClQ6/JuuTvWatQyq0EZrdxOyYBJ1o1K7s5wC7+nqno3trdLkWBeWY1jrZsffXWILe8Ir
8sIBk/up3n9Y4IOthpVA6QOnD/dI7ppSSzIw/HfQzYvkzDefaZkji80+vpzF+gCM8XoiiDlP7Tfr
cXM9cbkTUzRqtGmU57bgzTxWH8YVKnNANsqXi37vis4ce1r3kfJfCtNE2WQguNppxlKs0Gg6Rc2H
S7VpG1XrxICSWa8Xtn7/WoVnLDz7UJK1hvQzwYHD9zjyiTNcwjjPDJ9IdrbCGdH//0ZSUyAJNK4L
ep+zihgDe8h9nOlDl+1h5U5Y0rhchA7u2959JW0BgSLo1uT8/VNoXsOmw+NS9RmaL+UC7frN/3t3
r9tJ+kmcpR9eOnFHGwik5N4UXbzCZ8wsHu5L2vAwvnhaNf6lZ4JRwHwbt2zE8t7LVWuHSrBDwL4b
sk2+HS1J7GHTpUhAO2VSKwGZRdRd9OjDsYNBobXviwypseoTnu+9Q7lPW2Xnj8rARrRxfx6j8YCO
q/SzZFcGvKldCXmxNUUWDcjXbzIF00FMoygStF6idGoj5S4C+ECGOyNh5Uzo2RKANhrS8FeimGS7
bk2NjaX/rv71lu/12efqLJSuHsKesgS9YkHC5vL4efhOPzi2zVqp9xEYDkTmkgaX4X3u8Nxc9CN6
RCG2kEZKXQQAQ6GrvgKDGfNKH6SkscByqQ63SfqwZe9GCOTe34oQZS1V7Ez/rzjMmyoWQJnpQ7lG
Ojt1NVC9P2XyESGHYbsYQ6WECuFqaSP1BvR3UrEQElapESUabozzcWi+MDYCuEzmfkTL8cqYFlcu
3U73A3Dyg80eXqy1hrr79U34NTYeIaviv4WA54SSAPtZFZFNHpUexYMWobnNbKTLcXlzr2+zAxf8
5I1QYctZWws6y4ETsvLJj6LTwL/wKvzWyJ6pitBnleAVBLiz0U7d2wrPGMb1PCfmGe/iPKKxReGP
dO3rYlZYy9OHaeNfgLvzVZQWYH3unBv7JoCcaxYhISxrHIGoy836TptH2KEjzCd5jX3+hZHbS4zQ
YEDDnD0MDBb/WLrzF9UZe0rIehqlO6ZZe+7sUI78UdMDEAqwOf0tQjeXud2o72etg6vnOELvASx4
fvL+g2vINMH9QRQYP4LCM8yzbEJsmzXkoqhQg6DQhwt1PnwM2cGSwsZc9kIXPjqimfhZx357S7AI
ufidu9zQAAl2wniy2hQQbaVbIyRJ0GHGRbDCp9cRdej8KFG8bGAf2Z/u8LI5Ny0/fVM5CACWa0FM
QVTUxsrOpajuCX0t8cuFkPPWWcqXla0bafSGikMzGRpLovPGX9VnXB+/TBrLf7oSR9fjPvFMk4A4
+IyDYjJohiZJTs0Ezedxk0rR4SS1NZQFnxCm1v8/IfCdKeoRbqrDpNCZpWf0FF6I+O1g7Vymn+hD
S6uPBgXbmCAoZvbjAX2MMPqz2XVfWbcc+IgOnOtFleIp+4niP/fFRujiS06hDfxF5aWUC+koDdvj
MXuoIx/anNgRlRgBxatQQCNefTnWhv3UGIIjyYbrfCNxzrt9aea1RftRPEueb46PdqgEtZwpWKUu
F4pBPNTgsbT+5ACvdygasIRHLRp25pK1Ox1hMic6Yi5ig/Cgo091UA0zxwgNgtB3OVMTC7nS6Eb1
P19v+JlKrZVEbL7BzWWwJHgfV3Pi02b0XlaZklYzaw/pbhkIh8fueFNnpEOklAaFpsCLc3chruqr
iQGNBPq+i7C6tQP55SLV2MzJXL1RTj1dvkxM/TxcpjV7oILfFy+G0vbiNeZ/+9QGYrUbjm9CksVW
1OkN/gts/zrnvJP/4PdWb0glgG33WmcnVRjZKvFIzxnHbfhqGwgHhMfKz+OvHMv/C1pPaImUV0xY
+gLpCQiGYL2+MZw4Vxz70C8LtfMGQbz+/RTsI358GFS9yGA5GBG9l/RfArfgag8DEiH6Xu+NcVXU
pkFy6xMpuaLNQ4umsIlH/Fx5/gF26+Z5CnZQ2klMHlU82fTxwVhkTUkWU5pUd2nFySP9/k+LIp/v
7y3ZsJRRv3Giyxwy6Bd55x4a9gcEZBg4rsCRA98V6QYWkwD07KYiFK90+dG5S1GyyQEQuQ1K19yE
uD7IdPspXWbyn2/NQRzZ0SODOqMu8B5J+opf7cM0Cor3ApVYh1KqbVe835stg8P8qlken4Mcpn4H
Kj3Eq3fclrf2h5O+C64vh38b8Edi3rrMlz86nz75O5xJYYo1bwFSS1NVApxH+8bGdhPeCwDGeX8N
I9DA4MrVMb9VCOCQnm6pJAoD9BacyRO3Oqcs7a/erPauJqSRV8K09JJYVblZns1cV1qb9Tb9ThdH
asrz+1R7rOYOfrg1YiURtp5JlbDNZu4MdVxG7envweW6LSCiKJW2SS5ZFaQemFmlLsR0WyipDLpP
091i6X2Lsnhizh11BVM49CyA2MSyVADB3tX9Beik02iKOP4y+AevEz/I9qCe4+Ji///A2sJSA00/
OgaU8KI0L8rTK0ae0aPAQaMZ21BluzvIwXV4H9kEcNb5WJ5kPA8n4RVpmEVhDlgIw4p5y94JG37f
7Eop0nFQ4CfuDpqnYJFqs8yRgud4/ufZR7Yi6mmRu72GfQkGgiaaGnVvPrKMA0k5LMDkV8KsQbYa
SYWhgFOgN0+XmzP8Tckf0EUXBx4x0T76puRrwhk09dqhEpU63YYpJwCRn4geOy/IoFBGVssnW6dY
AtxebYaa8iJlZjAP8W9lju0xYq5ObT9NNe5lObHGfVxMiZOfwVHhIfeeYl/4IApH5UmmTVU8Zcm5
OdsHnQoRcSLtSiRi/tdg0jAjsSNPIn+d8GVAVj2EqR10TYA60wxVQEcDQTcjje2OLbb3XHttSt4s
mCoGWeU6tRE3kwsPBmFkQjIifvC6SawpTktLOjt9PPAXqKwdd9oymeATc6vgdybHK7++i1yF+wo2
07EQpR7lf/H/yD2NNXcDey0MmsCob7/3uvJOLGmLU+d6oGXHZCGjIKFUyCS0C+5A1k6lvL6DaQZt
4InaoIgaTOiJahg+qo1xQ695pGt0L355Lmaxpnn6G7gFPPk6OtpkMbH0RsqP+F2wFYHj8ylQSwhR
yot21LWpYjbXA100qNBE10F8DrhVG3FeEgvQivfZR7cNxJCScZYt7AZSUMCcQj4lZzHp1+9O3sit
qdid6vp4WTSd/aYXp5v3YD47lZexe7fvl8EG4ONd/YfPemmaqx8JsFshpmWJbnlb0ReZmYt80oft
QsuluycQ8o7k2j2IfpsvqgoIqAgRJd2BmdXhOYJTiXJ4N81wBOEdIyPNuazJcIQBY6537ShHx42q
EZEjhDlTzkf6CoMQlHRIyiZczE4UV7HJXaNxr2G8Z9PvZiygabPGv4/1BPAbSPL3OQWaZQ5wSr4S
gE6qV84Zlgi9ojCbiJKswTMJbbib0Cwps2BIjSfcUFZAT5hGtl+4VhdaDoaEyp13wRkwHZY3rY7t
z2dkShc9ElI8R4tLS3gATYfwSVDKqiPXlpBjf3bw7N3Rfmv2TRILOhkQpE1pzUICZdGXhgKbMMYy
XLQ357c8YDZKk+P05Sv/KCBDOdmXK14Uy1ZNcLRxiQKKZ/XdFxNwiXuR1v6o1bW9a2rwLWrIWsdw
OFi31a/lWZCPJZc/Vq+J/WaODRFBw+/cWQpSB3YnGoJXLJPdyYZCNFCC3v38F1Iic2Gedf1/dytH
ebTfiIBGLmFEszZg8J87NXb5H7PSuaO4Ykwu1lzVOlljX6cogtpWYo3VetL3GzXT1DHO6liBQV2n
XtLELNTotpKkv3O3pPAUOu0uUzGgh6VH1I6VlP4IIh9xjbsRXz+npSqGq1iDC8brm4bElkJWsPlT
Za3Z7I7eMTLplZwN2SXDG9yjuNSlnVD1ALrwvIfYRnubVpjj+FD2qfld0a2gh8kGUktW4OdHXZTB
OdvaIC6YIpetg/PQC1DfSpF+gxZY4+l9HdJcO9dXTltAlTuxZiBobWamoQsJP7tobdjnVLb/toKe
3Nxcdn6wvVtuCpcchFnC9OjppQfq1UwUOqq5WgWzqQ6JpKLjuiOODp0cM5wZHasI7M7aHsV/Qdfb
Zp14vtSVz/o5q6o+0MrmmrgbVM+1vPVPuXQcG2x3WyE5dCxoztqHXE0jp00rb2TWJUzyn1tqsR5K
GSLt4AvLMDrlqcXutOz84BUmU7RJKM/kXC223hwt7gUUqpo9hgC436Qhd7kDs/suzizpkGN2QVSM
i33GmQUUPch/GPCjDwuiU4sqCq9MHH8WjHXH5Z/Z7bpPjxjWknK7QBryaa4ILNy/xTG21xyx+i/b
32pigh48cHzvDs3UqEU4DOe4k+MEAAbgw1jZKlInqM4v2Ws5tc78T4Xed8jZpYRWPNO4A3TnjX8w
iRuCC1Y8cHj5H5HFEl7yr+fyNqbiNYfwsSu/tgx5hMGefgG5wxp1vkkH3TM53WeQgiDthlPQme29
3J4sfoJ6OrzrL4UPu/kw13okJVJe5WKaXjQnVTtCJF5H1qaTS3Qot1ojIiFYhFO2KAj26q8gPG/R
QWYpGbcnwIzMulFTtR8FJRVrbZF1rQXLUhDUOiq/+SduxKNbJuI7IGvR/06ynMX+EQi8e+hC38GI
KLPYkzZcRauPeCHXFgVr7ITtk51OZztgZIFJuHZeMM+8A3a4KjxAMrw9P1tfcdTr6z0801zqaW3j
vD+tOwoxlxNvU0rljcIVvN93GHo5vn3Afafx0g4DlRwnJZcYzs6wuDMmWLn5lbMKbONQZ1mhDzeI
8y0siCQAyY1Dk50H9DgOsiFGPC90/J8yihkiT5c4yhNy1k8k3AJ6bjMmz5kEGzEfhkqeT2cnTrKd
3Ag7YSVvV1xjWRz9qmMeUYVd9hQ5h89tp3oqpqyTD8XZC2Yv+rl80PdDt9mN1ZCmpnxYTCDBb+6Z
92/WMlqOfqx+vqQv5pv5GOYTEJDTyVUrHv8URp+wximcVjUEAly5hwOKZamIRac5QC+1LMEOjXCS
ZiCopJ82panCCpPr8LNnmnkCHxar4DrvoTyLKBnfW5dDGM/z+t1m9E4jgQplPrkNOYT/Xu8Ib3Qm
s1WpNHIUDyyuY5XHGi4LkWbD4rMjOrdbW/uH8TD1dRnPJe6Nidp8OyZBAu1YOtj5B2lvAXgJS6iN
3EGCgjlB4HO7t8U6v3w0eKcZFuEP/5vmx0RRUSQtJBvABpmxiwRf9G2wVcOokLJIlkOAxpQKa+T2
ZYNlSh1VAQiOxJaNk3OSllidx8vmVK5gLgdX6bt82oCb/IC/DCMAtQpp/7f8V77UScG1rUtYvD6A
0qaRvMkuOcHhTlHFro4llv7+Eqpi5KmrYILDNzMD0hmLRLsWpfs0GAHWT/X73jHNOYBmj/G/LyzP
/YKMVE31FFffIeihUVX9mpJWqxMWkG788f88RkgmHmV0cqLHyZrHKyTAqyMOFT9dW2F5dXfsTKs4
eBXBSHwHMcuSCmkOfhmXtcAV2Na40xcZ87siPh9dB+lIOzFH75LObFz5WPoECK57v3SmyDZM6z8z
CUcZg5rBlUtOi7OVO50uRbmLolk5QhcgaF2XRZaTidO/1mvYKxXa/eftnAQXExrrfgho6aTpdBcL
+18zn1vNZ/CxuZCF6MgCGnqdjmf8OLy3eJg+kXAObSQNV3W42Uc+3xrUNOdn/x3wTce2ZfPwAyS2
/P4Hn8TfCdnSgQg0iV/bHbHashd8zWokSvBAt/9RIJHmHNxjBsymdusriyLtH7NzePMN9I7NLquI
EBs0/nPf2JseaBjx2cZr9q5aN/WwzCVDrxpbuOfpSOC/bpOUApAKJ1tzWxv1qegxu4GamR48U1RB
te5nFAjsKxEdgs2ilaDSYD33YaW2xYPHBzL3pQoETs1B1mkRZ7fQ09uTPbp/4FrI6USs6VefQvyr
B6A/+WQrzBhfS67lW0R4lzjjv2juazvsKrwcNLEcoQS7m4cuLxgI10lc7CMMx8AHWSpcOh8BK91e
WQ7J0XXsZTAXrlqOeeyKK06rC4bMX/uo/82IKJqEZ3iHNhvu4AC212iDPxekxhABXcKWIFobPIyJ
ee82I6c5ulObK04q03QksFrr1LknsaJrFf5X4cAnQBIe4v7Vd0vavGJPPExihBkm7xJrSHo2d05V
sYEMYddIB2bpsKgDTc8y0zckgJJfJDvV3QjtzxFRn/KPFgPiJ9+JzgyTZXQwhRjYY0Rr7RSrPc6J
MK3wUcvXK464wiWWFSHtQPEn6ShboUnr7tV5H1WWZ0G4pOnfGL8Yj5xVafUMo6sTeqiIMLECanNV
RiLByDWCWGNAo62obhmyGuEXNELtO8pWI8Ix1HuhFrsny9Mp5jHXzCM/Mkep9KEjdI/4TpHjgi8G
QTRdPnbN9pda1a1J1Rnh+6UCaC6pMPjRqd58ynPP/NZZT8nXD5ewbrGfocWXH5oo95C0rmf9VUPr
22mcqjeS5B2Ob3WY9Y7VLUKzPlBdq/LHGITUI9BRaAp8FFtsQ592eYkOFJ0VPi1Jloel8diuss1d
i2MGeLlWS6klFPwJCUX2+aWfijmAvKwv8x0kIhCQTrhjVL7pQN1DGKnhF75ExfjgMdbgLDTMFVIx
CBnAuxUec7Oo85TaEXRWb+j67axmLWAeUaFifjzDIuNdd+wxAAQWOyQh20Wuh8Tpf2CUn9TAXEuX
IXFGA9QeLoxdZTLvYyMYAiu7eLlVj5IvU3H7Q95G265RgH2hWheGC1WEWkUyGADkUi5YSuaOfJCZ
TNHCY1ujAYf7sMU54xIlb83CPCiq7sT8ikpqGBnAaY1USb8DyzTeCJFfLwM0GlDtaTvddC8V59b1
6kis+7Q0iWmjnuxrZfVFbJ998nKisuC1z+ImyFNWdRkBgaaXKJx5ALOW5WrE03q6tXq+jov5MKhp
PfIg47gcrnOjRUnr+8lFW4KbOTFMz8CINvurx6Niqe+pTmzWk8SmIQoBOykWJ3mH85uTWcwUqAf3
TyNRAIYsZogpeAsoyMn7xN0fNtD7bKQRaZZIXLYZtG4HeDx/SkQuW6+Nx38aCevoPmSlArlKcOUS
rGt1JD/uiFQUibwc1qZoDrLiGbFhVdFb8isVWCJdI6+VEhvQBt28eJfvEhf8qCYIAQa7Saj4w42s
SCai3vBVgnp6f5NltivmN/883Ro7w/14AwDNfSyNO7dfZkb7ly0DXkmY0VIpT0u0ogPf9+Nz3txN
NEuOdDPxBwfH5PyHii5Is7CqOX4vbTr+ml3UHjyNGdRIzsARu549guNDtMo/RIIklAxFZ8zL1bdu
IqoSS2BOyY3+NtqvqaShlea0VvT8LNxJPkXI/aI4+8lVnJ5dAFzSXW/ohSC60gsbi6fZlbVcOiEt
820eXbs6TJLV9IirkmJ0LHBGHzgMOFoa+FlHhv47GEOkTEFPWhjOu49Lqr5AbtSMfjiYPL5voJ+U
qa8d1jKeAS+Fgal0ag9QZL9OgQp9+yavR3qkgJMYad1TXfhvQItBHtCAlmTZLagBDK9d7e24i8RR
o2uMCvLXaW+ZmrQcG+BIsrz8snJQPA3ofT+VCOuKuDg/RuZJdZDyofxEGYsov50RQvhNvkPvC4e3
kP2G3HB5FSFGhgS9jt+zLKavl5g4qmuEjyWdG2KDtC3SlPZk8d+wXx3lGK1Wwt/vevbXCK6upikW
JtyBbZSBK4Mm2y/Fg7puEUKHEFPTsJJ28RuGUT0wuo/ISy7C+UHK7uxOUx9Hqc4Qysz/FBueFqdf
wLWwRR1Le3U72f5SdDDFpviVOF2mmiD6nzBX1Bn2RHwRy7GuP2jbCe+3arxCJUPM0NJ3DO8XhmHB
mbG4DDGH9ecWLpieNcUY44D+z/z5T209Xg/sBQcRJgjXUEvHOa8x8Q7bnJOwQ8GPegBDHLwuUVOW
6Q6G/lIEnqapIzk3U5IRh24wtnmxSu5LDFFEuSdby5hA2a1P0CEkDLc67AbzolOZPQSslnfXjvlP
JPSCceDHsfuEKO4nR+ykBSoM7yC96sry/wu4Z9iApcY2mm2NxvbUxnxL1MLtux/NFaGIXLPisD2d
7ii+uSBf7ojoiA+WHw9VrSmNZDJZyPXNz+lP5CDG9f6T9pEEh7tcD5ZLwrvn5IURHDOMFd3/WUGl
A+/swYP2aUwy3Jkue/NAUuTbmJiJ0YrBGATHBM1AvN8TXIpR6RNOijB3DExeIVywlZCzhUF4GGFV
pGvuXNO1OZttGR4TD29vU/sFM7kjCPxzjSzxJvta/QbBXqEbExJ67wZf1IsUjLE9iDHOw02m2PPV
4spg0ONYKtuHC2Y7Cxl2OchA8Q9lKIa3ohOopsY52o4sBw3apc66XzE6vawyDzEBzKHrE4WstYdM
YYqAScA2c3Lw01lJ4L6Fx6JD/NvJ1UGCyZj0Q6go6ddk8SCFVmogcAEzwRfiHft0YHMjyPheOap6
YS2aufC+6zWwA6Lm8M9tU1EzRBt6bEWsNLvnicDwLrvCuNZycLWYOPxXfMFwkRruf+/YwDigzF+W
bV9YkcxF/+RmPJ8P754rCNVMV0Fp9NFzvztAkLFDfWceTIY7rNZBExxHMFv/95UvwiTRmB5Q2eNJ
8ngddiGTMCO6FOdl9AmRGnTjKi7JsM9O/uWwGXRB94xRdZgZT18VlZjzaUyIoxRuABhSTzfTvwU1
a26Q5NUX4/RFCHeL43+RiCEO9xU3YRxluKHoA33S/G1FRxDMfpg4l+Z404GT2QD+yTAnW4G4tLB7
4O9dMItdg+csbiDugoD7SUd2L6WDAuolQs5cj4/WIWjZ02OjFWopSufTVd/1i5saplCjbTFISiFL
ACohZtXYDD23jATqqnNQOXYEMtAwc/o9Ng1h1/+ADYTE8C4RHXvxhFNrDRgkSZaV9vp8q5S9s5f8
wpXKrpG7E0+r2n9VqCbgpMa0R/XAkhVwAd8OruhBk7DzjIQGbb6U7pM9saDhYlwoMIKWkC2LItxB
ysomXp/m1gRO3IDvjkzULkca9oL6CmYqbM2McjSUY385ezhMUBI5zzvGnsOPjqfTS8n/zlbyDYWD
5CjBLTusL4m7snkcvFf8ZeLQkQIytLB68Rb/NFDsWA52md4uTerJK7N2F4s3eTAon8kvhzIP/77a
Qc2WvCZgbyDV6PKWlLoSE7WajQOHyMY9Obw7fFZxQ6ohWEA1zIRKEgFhlNr6EzRvteJ4ctAcxsX7
Adqt8zfY526YuJoZwwFpdVO3y/17JpoP8d1QWU6skdkwJIXOIjBPDrUI5FeyYp99/565B8/mEkhp
0zmT6w2ip6m9l7xxb/RKGdxm1ImWeZTzmoMvBZpb+iWTl1/sxgWtDPiWYyxHOLNcMrK0E+vbeE71
8zaOriWzr80X8eOe0L2kPcr3qPfqVBS/RIaPw0h+N/FuK+vYH33xa+NQbZjU+jqYDhCpgKf0+wL2
Gbhd5F+HbnWkwy+a2SM05KV9pKPJ7GNLxyuMBEBTs+O2dxQVkmDATYf48pAtpPai3F46EBFzZS3I
Bq9fSemM1C9+30SU+lATKIDbsNWSumS0M0xoLSy/UYzWIe+aHVosti85rymJYMrHUixYS0rdFGE3
Dwbq1MGhK7bQBiU9rTlAYLvsrIGxrBWwGM144NDOiqAFqx/4gf+NWKVgYMbW8PEqVzr2uGuehGR+
F0sWNuGeECUdBF32GVlzXVdAxQdshjD0j7BX6gdm8y+crVRhfdlN+WjzlC8O5vKnu5h87s+28Jp5
GtX5IRbH6pcPqM9Rw+6pO+II2aP7CVYhD9CpHf0wqzZA1pBLH3dJ8e/3e+j8elYD7T+2f5UfhB5f
sxCIw19KU5wv32xVePWHeQyCpbqLm2NzAgQ/EEwsZogCV4y40U4okCdEH5nSvB581lrKWQWcCYEi
evFZUnz9iaOJ6nzq7EdKqO1jXTIXssChRFMm+cucgb4X1VvRv4iWPLJ0qPexTfuW4xATWI1e24hq
AxcJtHtbWWeiUs1OzT70/FSyj7qpIn0ye5TZkFValgcLnsHjF86wY+SqRMasNl4XYB7AGfpUIYX6
4VkmHfKsssJAvP7Iq3xJbpxpTY/Dygus5HH4tZI2u+N57c50xkEKmjB55JDNltJTSk+RiTraMZiI
RLaBkSKSzzGLkiZfZL/HC9mQodYwrDNGQuTA4Oxew6CYR56WAbDGX/kaJn6pxvGwIcYazKxSbiBe
VTP8SOAGT9OORdqGZZhlI61BsGN+fPVcWAdZSl/JXBGTF82eoDOwfPaNZeRhhUwACD+mOwVwe/0G
EPjYVx08V+UwBAZ8nV/tW58GP2sFAv8OAbCbz//q7vw0sQ+2EEn+rYvKDQDFY8VvhyV7e10j0Aae
1ceVjuf3qWYDAXvYd7/fCMgtMNvO9I9F7ec565L6RPle1JyiY7q90is8ZHw9mUJZX/IAEK+mQj7/
NnpEFiPvbGl23pkRb6WljMk/eMlHVlsXqNBudrashpNcG87bBepb12ldJHzmGhrbDGdAuPOx7O2u
sVvZF+O6+iq6bEU2VOowSkPsoM6Se3Tltv4JEBhVGlZOXyTBn8/jpM/PnIrs6TMlKFzsK3clP5uS
puoresAd9g0wzpl+J+HUxQ0rKehy+WELfyEe98doJMBc/mIRLZTgYVJUNbAVpOCVluG5OFpzFUMs
i8fVFPjoG0zBzyGF88ObqQCmBITDHr5er+vVKIl782akPFy1fL52Hek9uo1pnlYlNrOUwaXiDo2N
kMI2Qb6cMLyYcW3wsk+NiQ67bHZKurp9jAhskWY28BFoQ0XwYDB3M/qdJcV2V7TqHneBUxMIH215
rmWbqbtBpX69LygtQTh7B/Axe9vi7cM94EsELrJEZU7qLUwK9Tao6MO81PujLLUn0XxYXKXXbNcD
uFCuTA3COsg7xYKeE5fUAXw9GJjS3AkYTeEbIkQv+QPUHiMDbuEiiVxh/tEwNKPmRvkMRhPFFm4q
WAsGKrwzW+usPAQ9b6u3J8wfspklvgZzUwE5GpVFVoKutnW5yGyZ5th4/d0MZG/wKUHFuuw8KD2J
FxjO0CLpVT7BQ/vpejL7aEIlFTehaYV76w/nPnsE2Q4GWr9EkK1jt6x5OihxdTVPQxf/JVWcZxsC
PuBpUpu+nXQUh+AJL9A/3otsmZO65tOzejR/X0uz07qODoOoA3n+JIyTAyJjK3Dk8tu4z98/iKy/
RLrhaeY/Rs82+T64nsB2HVMOiTGxwK5Sj22YQoqmWN1ZgYzPc5cXMbPQbpWoR1GNTka9Xgpo0H1W
2eBxmJLtUOWXDTWGYG1FMVomCU+9oqD9PEowO3FjKcXjRq4WYViJ9RmdQjj0SMk7lFGlT6P7fjLT
YYlBj9K6zBKa8y6MbcsFRI1rrIIcI6Jr5fIUrlS6ieyvQomkVprWlrz7C3cAWqml7zpF+O+7B876
uS6cqlQEPs8nEnxU4kTWoWaUUZxLEkcJjOivHrPygde4bfWy2/AMWmY1aFUKLmsSv1Cl7PKUNDQf
j5Bdsi9vRvnHp1WOKKDKfd5ShWLNARdhZFH6DUfbNsFEkgAb80I4TfJqsjN90jiiQCThfiP0Iyvy
gMDehFjJPl3VK/U9IMpuOUVQUKLyqRSd5nt1X0/4CLZbny1Wo8/thp3eom8p3jLmPb8/+aaigPf3
9ALlItbgUjD8a74qyRtZMFi8QcvbO+fRM+adAXsMQ6QpnanB+5F60f6yFO4Dgw22DJdZlRacGIqT
LQBW0nHs/3R1ukL5/KcdRZ9TTc+eRO+N8j9rynz3DDLEBL4/K42YXML+Lr8qbxSO4Xa+UAUOE18f
I5AUuu9nFUlO7dAadBZn//If+ANqaUncuIXEXHdC5DezvDHha/YjGhE5Fs09OcixE69HwN/IpcNJ
HGB/CiBwkKa6qSAKy2aUCRcUwo+4nbFBvQchhdH7JJzgmzt7GQv+WH1TRdBoVTxrMTrDKuBHj3N/
8u1dOq5yKHYoElAQA9ErhgbOio7VmRoe7u/3kKhJ6+1+rBq1b1Vsohg5MlX7oC6zMvXgOyALFcAV
reTYZC+2YpFh+96mV32s+SaZcvAMh2SSXmZoFHM9qv3AXyYGXkOtQKfvkl1p/eUPxUY4WXsxnMWA
hmBJuXl7XskITkPRcoHLs2pBq4fPeZuQ0t1Q2bEEYf4qm2t8Rcfe06Zgxoyzi4zuVCF4GBXEYPyw
NGiVWADmVqmXn7gmemaX4LXkHZoH61BfM1cX1+8ObGRvhSFl3nFmU5w3QilktWVd4ALlX1FmwGsK
C/M0LzWtNNtdxmEtiqB2nXPAna/NJflpHzuNeoq0xRQbr9u+2PvCZTo31lGb4jJb2vN3qHvmMNQF
y42Jp63PJDaV/gSES98WDsX/s/YImg+ykDr2NzKdMu7jWvfZusDmNuDWbUEN/ddAiSrbD9NOdljS
DVs+HYdlVnoN2bBSpg6aw7CKkVigH3n2ZVPPQgJrzSYzcQKcf6pjlTiZtN35/nNcuQojwIkvqPoH
O76DxlBStWU5xLbtUrOVZxd4AeCJbnu6918JjqjDzKkSAUao9OWjPEgtsMnIg3EI1y8/qukkpEmM
bhRPAvV4RifPEhRp1Prrsjvwq8WA9L7f5r9qI/IeIsOJI5QxkpQ07qHOxWBD6MSn7Pnbi5/1b9tE
JWaxj38x5xJS34N6AZhJQrT1EsQdGwy2k9F4ejYXWM7ykXlihTSguvepVKZarOmwEJayh6rZVO63
iF/sp+prihcVuola0PpErxIjL5caQyBjBj5ccG/pku1fDEIfdKYcCyxrq+1t6Dqx4TsChEUw+HDq
wJQFqg+UULX61SqhvNuqNin3tQ0GUmWpJelSLfBRbCotDe10mGseoH0Hzi06fhIWgLZB6px7lTch
VpmDc8yUrVmnsyR0f51FNtBvqkfGkSq84FEkuByam18AZjZ8pzSqWdds+uCWfUcfffChRNP9wR9o
iumBUDNtRlkyIuJCRECJQtzvbccv+eRF2FzNK947xIHu+k03Xu4mtzUtpndZhkNNLA4PBcNx2Qg5
teh5wTz67hjlAbJ8gIJoG35CWoGZDIIlQAGGLYMwA2/e6T0g7vtuAoU5WP1tfjDYfdzo11zFWHsE
maqqZt8tWsZ9rRIRHQIfTrAuh2Zr/pmDtIjNbie8sV/hU2FoOoaOCDluhTODiO+0hee/SkDwDWQ6
yc9yZ2w09/SWrd+QN+dNiKG/kGwEIeBAIyOxPlWD3JZJBFNRsanj/TK6BvhD6R7Hd2kuG0Pg4gsH
kAa30JngVg6KR5XDXD23qQm6/3Mh6h++MKsz8J6NGwbLFIxaB5Zfk/ZbEB0xmUX67QhuyFPjMZ8h
+10dj1Q2Rpt1JBYUqK6yLWiswyQ3MHiB/3e6WUrrOuNCIt/lHXcwY9tvbuDFQtGt0s73y1V024Av
K6hhHbBSYflrXqx/q1G1B9OEBeUfcfpI2FGcIouMTq9NZU5oY1HeHvlv8DRShS/2mPd9dXvX0Eue
zfHVB8qxWqnFc4wjK9nAZVCd2EAcxzSaYiGfMSoNZ79H3oCAJVzxnuBAx6pSSs7KYBUjIZO5XRxV
MNmu5uLm8VmmmmM/fx3EnAz+sw37feKNF0hugY+20CHoQ99VJJL7FAFuhRR+IdeP2ijD9JGcadK2
Yw4jstVdt0NUtIkBMbYJ/eCqcmRvVdtkuLt/1NRabB9tWDRj3vxq76yBGacx/wER33Zvm8Q/K4dM
3qVODWJD5lhvp/cf9IJ6fztRCfiTd3LHgURrEUVopgm1zeGlpISobugm2mrG7zRs8yV4fqIrM0aZ
eini7YgcEC8n5p9Sx4O9jAgIo3uQeF29oGEI9BTHdjhYXTvi6Pkzrnxh1TUg1N7L7JoZ8Go7PfH9
yhGh1Owg2EERXiLYcCs0FWXHR1n6alnoFVDI9whYSooaoa9gtBFKSU2wDby8CoEmf7B8lfXQM0FC
MM9J+IH5x2LnnFcpfVjoChZ9t+NlXEe5LbabxOKWRAwBC6GO+peJjLE8ZJGsXyBaHDe3XpmjPqvc
5CLKLweU2ygJ0y6KuZfTv7nA9646IJz3qJBcII5MgaGYicsnizdLj0Cj/Srf8JwleIBlPEwy+JO7
gFrJKEGp9Jb5BolvHuyOX6FCxwKdS7pwxEhHJ3AnLTvGq7qFgLWoFLYRW5olGeQPI21fcWMkWdMN
KIQCijYuc11WgUF1FUgqgrqZyBxXkwawmeOtqgaFuuP5RUjuaWL8Q+d6DObstVfzH4nD6MpxYKlt
77Wbk8OWOyclN9+l2ivPVkw4CbNf4+8MjkZrZfKl4xXd+dofkwDw40cMjd8GqV9nDeO8C45ruzh3
olR6RNIdIQYbkZ6ODXv3MsGdJzOCPwRqkcVKziH254PzXhDWdlX8Hz0G0ROzELE4zeAYORaVyaFU
XGTYQAYSRRBUNk9PlaoN9gMB9iuycLFCE8jAm69o+bysLhayQSQbiZfAyYKXtrYS/sTN+7mL9tu0
Md7Ncxo/pSzynXST11PcEOU08WQnzRKe71wvJ79gzYvm9PrxAmc1HEgv9myZYG7MeNDWRsX0qUKI
bx2YqTRrDUQrqFMYEewWTBkUziCt4qsKiYWhyvK9PYr2R+2tDAM34FbJIiwGSQpERUo1A6S9bBWt
2zYTeK5v9cpqw/e8HMBMnoXjGEd2osw5Q4Xl+H1RbH8Mqj/VGDqksBqbzEJLdfkGfmEVx0bDVtEl
A/XLiN1DsdTwM3LV9XueVT5LTPu9RVinURyrVv8BIGqmQGrDhzuTUk8c7ft2NQw5WkvG3EibJ/DN
PNHxjEgSWxeD2saqp+53jf6Rtz7+k8VTmE2uWCNmhKzTrbmJyHfteAZ/MPMXYC77l9cQrnQQsZR/
K4TrHwxWC2lFxn2yk0WHG9CmfcHpJCcgeBkR5KyvnnLri0Cp+sqcB0QB3N+tur0XCmA9yb3vQZR1
l+YwCu5MUVEDj1Z57b2g5PldTyKtLCWy4abBPIHpIIVjTj1lGkF7tKAg/mCzpFzqdYWrSFAsaNui
5RaxhaJ46cG0swXKdxHGe1InK97isA2WwS4Eaqn8aPvE79mGH6VVemtpxQGYADnTx+1ZWHycIp+C
4htPrk4x0ZC9xxuS01tfwYn7wd/kWvnCPHIfbTCHHl/i6xmnHenlkbS1hblU7GT4nZ/8XQsSR6m0
+x+Ne+wqHThIRBje1PjCj0VSwNb9S3TNS4PecrWT+IPqHnROI4B4dVm3JqDi+7W7yPTICXkGvu1C
BBhwwQmFp1OSY9d63AoEh29IDdvLh65B7B1appiV9s0+9kETwuyixZOfMcxRgmyqugSB4EpwzIhU
F4f22cZG0deKMF6zV/JJgnw9XhczkFnI1VOfk5ra1iFyhYMfSbGvx4M8OgQR/SL7EUsitZfFGHph
c5zf9FoMtFfs0suJoNnqL7znoqvCfmHxAaCuM161FbQo23mbhNWwj69IBT54nXXXp3Dq9gOU3pGY
g6OlAlsBGnSwNWML4/qybKgkJMqGsoCyL49wHek/H/n6vmhz4A9Qyvv6xV84s9Q07ouKDhfJlz5I
pOh7XHybT/nBx6z5Bcb61vuJHHCx28J7ojeKrjW8I6czMxr/qDTgiGpifG3wQcesSu1IPlu7xzDI
teA5RG9BCei5Xl72Cucre+ZJ6JzCsAIy3KVHsIqIP8x21Q+OEDfpNyjrnlysUYC7SU+EfuGUIeTB
DczkDK1YuzkudNYqGN0RDdMWuZ75gY/4r9U+qEUbeUnLz+zZCjCteFHpGthXj5fcPLM7rrCujvFV
28pmbdD3mEKTBS46BbZPtChmxT8zglv7F9bnrr+7pA4HegBhn9v86mfK5mkRJbfJVOuLWXbemMfB
lnjzMsP/gf2OiMg14OFugsT/9Hw26ViymOo9qwnoYC4gYTTGNZ5OyXXv4YbZbrasEM/TO2YGVQC2
Mo3Yd26PbCxek2piADrpRF1gMYH/ZB567gbUx1TNKE1kcswoeUYYYo6NoNFYh5RWxvsgsdvfForB
y7PiEO5xa5w3u2htNF2YwoLN+WsviRi7JhP3FBqFwhy6rxXC7E35u6gbpqnPccvT2WsBAQKnP5ul
wWAvVvXhGDgg8oPpTweShwe54ACss0+OLdoT4w9tyhU7f4au0vexEwdZJsUoN8+WZbv1yzIu/P01
Qklhswl0/727+VJ8R2+39up7grjljwrNNz+YYTxQmlL4G/7UXqsyQOPeZAq7ubYlGD9UcE67OeVE
E0gxlsExIt01S8B31KP9nzLIsryvdyK5+3YEVo83frpoEf49bIz46dIsfHKFNZ7K/wUP4kj3CB3r
d6tFjq3sSKHKsiMOLONCK/L7n1NZxeVYV+oHKj2KguqYh/Ux0mGh//yxxkQLksKXI1/OnrwBIp/l
OW3l/gGhsAHoUXmHv7H9u9reDQFRfAnjRBG1hcVHUBOEobNMjG/U5H18vMaclmR2lMUpLKvej1rY
LsvPDrNyPoZ345A2ujWIUQAC3+ZaV/tvz3demN1j/LHPaK/Nr5OK5brpS7nzzVcs8C0JHPbfeRJM
LMYpxKsrMhCO+nkWZYGWiucGS4p6QQMeVAP0idHsm+BW6+nplVLQvUPqqDY8qsnTPlALV2nHUn3D
gb3vKGBx18I6y7JFeRLuLClEOX7CYlMQVJvMWTofxha/DyJNt/vTJ+ZqgXiFofwo/zBpkTV2RoNB
6yADYIvJ2zgxmMiej5u5CpnT+JIBvRB2aqDK599ZxTeb+zO6lBSzBhym6ZwlHcbshpXcHqXtvGml
sP32E4gsskvS9aerZ78g1meqy9qp/lPahirSp6tMi0RDLvvPWCpMx088VvsttU/jpw1cWlRk+T3A
TV9VYLlvfROY6ZeP7JjCRS0ZJC9ygodmPlIj5PjbCLDxQC1rd5nX0My71i1k4M4UoRd73zR//RqZ
eqA3VgB95yUW3qq3mTloQSDV8Xvijvw9E97JSBn2m9YsxBuuuczqb/YfLiifQdjEGeGY4f2w0GbX
5HKXr4yabj8pKLsFDRoikIF4wScPmbhNcVcLu5nx0ndCoziJruAjmdGdzXm5crorVnXZRXXnYgFO
2jBLDiS+p6ucEnd30KXNFO/tXLa3opUFuL7GC0frZ90A5fnlBK7vwyB002alS2xsKL50KncZSUlZ
BZUXXvrlZyQ3NDQRflXi3QC05O+F0VRZlAF7OKJB8RsHpVOpxGRKttsNx3CX0GIk9xn4VIVbLSJJ
SjAJJEo4Ry7kYxJtuxmpMpYSkGZI34xSwZyubzigkXEX2VZDsiaLdf0EKi21J1stD+DBPdnQBrR6
wxaSvjaPuGiW2UKpuO+k+UGKMtYsugsDglmWvse5/J+EDrSYvVfzhVMGG0Evdqk4sEPlpmUwU06y
T0P15TE2r7k2T2Rb0Hy/vrxOTUjMte4OtrHpAwpuOltlBYKwxcdcKVEOAqA/3X8I63UF41yfxCvF
ozsp4C+er4YlZ9wn7feGIrWZ1jvzjK6kVsTGqfz/yFq1w2ChPmChe38drIt0/a6mPVDAuJtcpYB1
fM6den7Fx7T4z1ECwOYtf3q/tlZcLEICDFAuApgn0MdPbCkcUWXrS+aFs763F5PauLJPb4f2NOhf
pyWLiSruw6g2OUpIkdQ1h5x7BEjSWIISAHg/i0O6utqzHVpjSq/yXKHThXI955JPuuvJn1n9EmNH
3kFjIdC+Aq64f4aWAzJVcqBE6PFK38cqhe6Q2UQFrdHgqgmkITpIIeeDi2j/raYTkJebyy1WDLbN
a573m6vmFqxCytslRD9XCgy6AenW+yEc/jL+Hvm6+XeM4X+b7JL72DFQZqm8+NZImA4tcexzC0XO
+IJ7sid4tqabYETXB/h9kvESLcnacp0nmqlVlvvy2WmD5N6MugD6E06IbV8BcTHOd994i+i+hY4z
NPS7LWxQ4ctoaHn/zipjQkb9ADDQGuRrw0jMFV4GglUvgsjpNTjyg7Rjhkzbfpb9knvDJ/isWKnB
cbWZ8DQ2g6O+kgv87BESr2qXzdcWgin8UOsNHbriiWTMkL0JVsfQw81TBxi9b1xzam3LPDKH/BPG
S0T5K9ajgTsFHSJC7115V4GbsNZyeVu0zjKxyp3tHZoQAq9oJeY4Ipdayhv4mQUg/1l+rg7zaOlM
MWUXRr2uY8AAk2tnPaPUTs3yiNv+iXrPmEh4ORxje+lErXMXtfgcWlvoIknTUVp6eu4gXXdap5bO
HjwY273GlH5srrPooY4w8qU/5jNP3Y9QmELYVXMNBJNxujxZCwuAvWz4kkIC8eZCU6nk+QDk7Ok0
swhyVV4YVLNA3hc3SFmH51IUnKIboHmQdiHW0QaCQao1vEmzg3LcxICMKHEpf4vVp1jm4rqSX11N
zHpSrcSOOQVXTB4VoBofNOV0J/rhebleG6dAIAkETITTZJH1Tkpmutx0rRvH5yf8MOZfRDvIe3ln
qR5fW5NbM0yfYmhriSdxn8oP4ENta5fvzmj1ylhBHQqjzc1zpR0RXlHA1b7Vqv5blhTa8z87YugP
svFYth8jSG4PBxAkZn2onKPftcpxUkk+Bbu1pe5bsZQYwopHDG20F3VIL9Te4wu2Ba139n0UR9B+
2l+h2k5gQQfGnZ1kXPhygc+eQF7cLwL8ASlU+dQDvoVuzTGUrWsAu+1OCZq9gm4iee8RBxvWrh/f
6pu2w5J6gYSaL55E3iuhcFXtfDkswLJ1zyGR8GROX9J0R1Bl4YBkHpRqbFw+nVNi6hCZ6NxAGFmd
TlOCa9By45SHoBPU3geZEe0oRB76PYfnCpJWUgyk9IkNFxboA4Crha1KTaZhROoeCl6xuQIdsuGm
Wv7yV0+C3Wajk2rsMGjdzAPuYGH4bvY14G8XIjdbBHYd9O+Ja6HdtiQfvtBxKb3SsUza4G9U4RNY
IQgpK61h0M6hsy1cLCjMBG2cGOErzg0qoaVpxtKEzaIL2Mz/3zGh1KV9Jxl2jlNcVTCMgWmzJBZc
7mqFu+wWAV2FzW0FY498QroTtJaRlZTDpfYd6ecJvcVpbySInx/QocMDoI7MKelf+ryq4py7YCH3
ZAJxM4FE8LuEN9KNwwpqesXvPRiH4sGLVEHugs2Of2ryws5dFgGtqyM0LQVH4lV19ur7fC7pp/82
AgE4N9X8DcpJyoTgez2R4HtwLTGkuG46pPSWXgQ3DmtKJyolyFM5MqV5jfFLu4M7uaZ/JepvrwZ4
16MeuFPwWHfYOjhNbV1At+W+UmAcAbW3M4L2KJKPqil0fPvK7J2C8ja2IFwivYMWNsYvmo+LJ1I2
bbO8lWstfJ8fdSG44+Y5YYPNnG8i1Cofoa0jHzw62uQ9S5d7EM/h2GkItDEFwmCzp8V/wBiDMLBy
eKMm//SqWJ55ZYRamW93/huPz64w88F+oGsZizSXd9Pi+PlaNaz1wWCU480rcTIzlmGrVlMYgDiA
8MT23Ty680BMJZugJgu3DJUbiuHNoRPPtUZFUOKRwKfo5zIoJAGy1Zz0EPc97xp0QBQ07yEV7EDN
Nm3yugsOfpsjCv0is7hOXBtyt9omN8bdgnmCIiLBopenryg8lNdcBmx6SYkWlWuUmhXtfMg4Je91
Wuqd+XCA6O/7E6QmX43AN58Jlq030/oxj6VbyLtTKyNqapy7bS3xnMyOHPhHfpHYim20RfJStjZl
sQzOgpC7pPjsbf3Qs6TFPwvpXzH9F5btWO9mBSh9rEoSyFk5MHW96bE1LdXdYMGnyTWKb/rEicKB
TR9U3AUqzNVmn0VF5hU2MrwF7WGJ89V7u59IM6zzJxe/6rlH2GCslLWQI3JsGktdy/rHJkSltKXv
BtJwu/V+l5LzAhdLJgBeoD4hZaQJu809ysx38oy0wWWzUB+ekG5UD6SUN29h40/ScYwgiN49Cdp1
0pYZmsFyuz4SHqrap0afQ7l6JawJu8JAS/+aErovsgNojJcjvJiJG/YXUcX3dA6GQ3G9aUgT9Kui
10PJAYVCB/us9amvaVGObLdZWXexDunuc3n+6Z9DSQjubLvJi+OByaPWdF9wB+f8hvFVlJdcdusf
V5YP83+KALiSytjfxBJtsEAwmtSe4NWp6XIqQGd8phRn9rxR+vPXOaPFAiV8fjkWvelve7qP9GtR
G3CBjy7gKWIkXuwBYVKZoMeqnNlUgdBpmD6TtTz82Angd/sk4rvynkgwUedc17JfLYCApyHwp6MU
5SvmfD6HNSNElfsG/uSB64kCMWrHJvPCkAyAgu977Hq/pjEbrewp8pIHxldWT5GkoYYOZfGbQlGs
kXHurZn30Y5J1FrcEIwFGYlllhhCg4idmDBgVjkfeEtv/bVMGGom6BIkQYdmPZenT2fwHgN4s5Hv
xXvLqIOQhpfd6iGfxFchF73m9TD8YAtssrfFQE6+JbLWwx4koQmkQMlWJg8o0ZbQ5egywFov7z4N
FyiauYvcD5XQjQhPdaVGqy8R3jHggd80tcl/NjyHvhKoyEuDUubUJ30W6EHe74mmAm0iTRWbMb1U
bUhIf5ajhpXx8pVb3eFH+bxKXZ7BkEyDSdYw/0AJkEOUa0Ev81+Gpz30NsKRCDodWx3bX0Ss3Mav
lBr92IzWqLK0fvjhV3VpRyFX6mAEkttk7SK+uU6afKoS3axUDk2mBWPHoJgqbz840dWC4iUPTOhw
drziRGB9Y5z67Adh8aG5ynOmU+rMU8HVLdkfk8+mTL2dFLB0UMr2BIOSKiQYWHHsw9YC1Lrm/6X6
stZyDB7p1dHWCSa0PnuDSFb/nXBrvn+tjCFKTWMrKjit5TFH/B9U6t1hCz9YlcEURkBcNmXkALq7
r9kzUXqPv0lEvd4N2/zn8XNsy9nrzhArqrUCRctcw4HBYSjnekk5dswiJs8IM3wVihA8hdonv+8d
b44Q/6cCZUVm6h6K3qnaeqxz4BLWzTItLeaWXlcgr2tnVgwIlA7lTz3afUcXop+CF/Ro0+GPCcXz
In2RIbX9/Ss1N07UgAxDO+Tzi5i9ucyb8NuAPIperk8EUpVhoUDeVHWqqF7mnZmXDkfLlyYs5bzG
h4UGNQ5+qkfEnbGwUs+e6lLV+COHZZmZNF2vL7/O2kBgGuAkUgt+kN5WVFirL+L9P84FJRoq3l4y
0hrJLSPykhF8ATVAL6WKw3hyR5VAqXGJT5OVYVDcHKfzPgGIJs2e+XlurXj70FOL4K7bg4EYEEMI
a2vnsUYffWolVnD9RKnNc3h9xuJxUcabuONm/uQh8rbSlKgOdJhrcQXsB9PS+mMtVsK53X8rwhxu
AZRC2DowJkVA/nJyulS2gFImHwPB5fRYJBsjVKJniTPvoPNEQ5lcZDHZanimN4gdd8FNTNUfw37u
KL+1S+2EUqiMudiL/cmXa7y8wF3zy98tZ3f2dh7nSFm9XnXKIK+hmFNWLiXVrqUlJuoBDjbWHdz8
TbDV4BiMKLkGavt5HSRhbgGPoEbZ03sFsu23jUHWGcfSGW10mPGG5gogv4AUO6WzkdPGfErOaFO+
gStOcKeiDR8dthuTxLpkBY073X16P8WTnP19kF0JPgaubVJ0+XNyYxOIZKZq270GBR2OFde311v0
jQ72RBRbuFILboas1DYp+kgR2vmovtuFHCwi6Dg7z3LlHojC0RtCDHqud0tM1FirovNAMoFKvEbU
tF6xPlZCGxB+cfRsaLMuqABdJZxYcBceON7b16Ew/yD5YepaElEFOb0IADCUgXEvp4tr2Vaernkx
C8Uldg9eoycU3hivIjz/jx7pr0gYzjGeq3f/HvAeqek+2NvJMzKR9vJWfSvKiYArgIuekBMzZ8Eb
oAHXHK5pEtvPyp8YXeLjQMhuu5wC74sq5qiUIOGV1otSxhTqHSgy3abbpGEPH9FMzvw9nMQpA7NI
pUFfHHJDjTr5AF3sWLpILLE4SNT8lefHuTJK1AUIXUd3IzsA3+R+hcFcfZ43muJi08xiaTkUFsTf
//6hCPig2U5E4qGOzQ6P+t5XCz52wa6TWlFbHc8hb2HuMN77bVmogL5uFfBpq14emMm9efYDe6Qf
iKJtYsiQaY0IFP48oLFjXygo6Q7DzyONojtN+Two3U+CgARaROQy7ZgUTmCb/iMh4Ul9ojsgIWoh
U/TUWCa0UVsPxwvFBlUl47PCgqe5lhAK82b42frVs/X/D7BUsDxBK4/I8ssai1ey5GC3UZKYIT9M
f+V0hctp56/d4+HrxPE6jwHDkkjOBaufDbjlk1AI2QUx8fkDAtDOt7RjrsriDNk8EyUfrFmKraa0
Uq2cGJxh4Gr3tnmXleZ0DGqyDJ/6gLTPlYrb0fM4Uc4wazCvCfR0bK4NlvYgVkyFGZ1VM+/aMH85
HDkMSUIrGZ32zmGJVguyJKxq75xrhC1Qvyb28okyV6o+D8NJrepq2h8dsnRCDImuZraVtU/l0Tyq
/aaNYFVKZngNUheHkLnmKoKVKgKYdhmS5E/UzaIpmK7TCtQ/lVi9QU49uM/p0w6P3aJUf1q7oefy
d3bDTBaGAXfkm01NDZnRrkkAYcG08IsoZF75DxCkvoLvbdTmYLmfV0EXWW9iDgeDq8I4sFN+csqy
Ps+hm4uRiNHU9Zuh87mBdl/9QAi50omzlILldk8ZXSC/LlCApetMY1JmxZhknbCnrECXCV5Na9kp
hUDTNE5uG3oJ8Dk7nntbAPI3xNo7vectX+dJXahNPccf70g8M6tXLraBopUn4ett1Y6fD6tuL8j3
WnIAHVYRkYCHOobo5ZNc2HzuJDRy4ntnjQAkf/jEVe2WCTcWSBAkfK4/xybXmpNGjrxVUf/U+zAo
/QJQ/kcfKGoGt9kKv1xo9EzLqn/+MhM/UM/aMlF4KatqN40VsVf7a2upNQxdk05390MzzXPPPTda
hIbS4f6u/inU0coYPecyQW5Li2E7AvZ4jdLHHI8Yj3zIt5d3ngKwZzdVzkRXbR3n74QgNdsiocV/
domeNVA+x0HrJJgxDKBt49DaTM9YC1LcmY0q8FK/RRR3h8/DJSthWfbZKXEpVOX+EZa+ztrtRY5n
av2gUHMfRL7FNnTh4XIoulpmzh1bJre6ruwrOxkkSnjyD8O6b9/BYc0xTflHz+ptivFRsOMh8HIR
bj9ubbZgKWAVx/JBLcmPwjr7z3eIwvUZ3LPbQEesl7pj+K3sbvMDtWY8WZvJuXLRgqDaTpg06EtF
9dxHib/wUr/kIp/HuV5WkTBHqyi/FFfICSxO7mBg7Bh2ljd2YcLQeUPcvPWZ6uWLxvZ2uEaidMqp
sAo2TOkHrEMdCKLssdOHfdH7Q8nSnQUOUhKtkpd41jZxKF4IRqEdAm1RdJtJq1K2W6Co7h4egxUb
R7QXcFXsHLZOWhLAF2UplbEa+q9cZxppH1oWn6GRkKNOta9/VyI+t5Pbk/fX/fJuO7ypt4ehHQGp
goLJlNxl7KzIGyi2uvCJS92Ik2WgcIZak9qoAU8TI26tKXXVfNXVPWe3IsPFqrVdiiV4O9oayW18
89VacXGtC+K9VHBM7C0+TxcFDLz1xqVpsZgapEYKCk6C+u1wunLxiabTmKo0mJGc2WombxHnutzf
ZF9JZtIURZA8VeFtVbLt2cUhYgdY3pK8it9jrruuzdx2NbHo2E9cNWe1+fMPYtaM7ws/3M7oOk0u
7RKE+231jSEvb/7FtHXtfqWcHnBBhc6MvOSb1czZ4sRwbLa3i6hs+oY9+kHuHvSDZCCR5O0B8ryK
jykscFcj/e/Fdi3ma2liryB0cY7XnBtTjLrWePPksAsGN2acteaXc3koPq8dFTVQH6/EuDcCggGC
7RuYTavPxz3zsjiFutPvyTa9s/OlpJxng3vRUbh8HhnyrWVOWLt2uVvcQ2LCd+ttUVMhuUaZq55n
jmUw3tMABem1eIfMyDXU/IMBMO6LEcRuGb59Cx4J9Y2wPiUMBu7juGJJttjVlQDaGd5LA/1XwQmu
t99wsx02xhKbJWOG7EHX3sKYGYXIvQPyQbD6FDuFm91fyRPFaDCiA3i0IMFxVmTMI4qSyhuv/rbi
ORg467pZWiTS0i32SoGvVpj+vUkderUNaxC5+eVTyx6Kr1e4Xtwj3vQBPXqnWej+grX6b5MVR0en
Y5KNUaRduPEBHR5hUfODEOQxN1pTHmiXjgreyJPXO7ZcVC1GrZ+Lr87jwv0vVUWSzvNDBQU2sB69
J5YMmfx3AIHbAjozT9rLS6u/w8fBA5OZS7oDG8Dorb0IUZ0us4dDE9mXAnWh7PogG+XcI9er62Y3
rWZ1M/5bAq+mMTrzocHfhQ4h+iObkfFPI2YG40QObSVQr6ChtZJhM/phL1LBLLOf1dWMK4rbrbdJ
BBLMvT+hUbVflYDHQGr1/kOdqgkx9ix/bUdX602YXFEpW5H9uALleEV71gymYdN5or9rSmV9gfdg
3suajiLCortH2EPZTjHbJbHKdBOw374GQpTFTducD1HgJx/aJjfJNdoKRHL8WGn0KK1O5OnrgHWg
6Prfxea028lEXSMDSG1/VrJEHr1enF9Z5LeSQj9lPsm6+jNUMfz7h+EfeJetaDgFMFQlryUmy4UP
k5jK1+iyFXVYyuSHbsPvrJVJqr2qpOKvU+PX4UODxTAuB7N6Fv6rfqQI2pBojeboCAuslsi6BLyv
ALMXXlwLvdOZU/xEPzzvKX8s9wiCbjKE4MozAU507YaFQ3pRrbIlXN7WwV8WISmYyLNfeY/oQiDp
ZB5pEey/sE30fLKWBhrOHF3f+Hy2HRI6TgSRcKFgkRWVK4SDgPyhjTCL1V0d5Ci9KRCpBo//ZIoh
sCMmVcWLWMGLEg2yGV6NZRdUhMC1IUGSK+pVvIWTuMd4m+u6nedf5Xz6OqbUKk2Af1jc3mSsiVVs
Ex0SAX7QKiiNVjkUlImLNJ/cWbUmDMFfzhtEoBl41jgM2Aa7mY/e7lbOW+x+sk8jUBRjyMq58EMW
sHgNbhdT6NI7TO07SSOdWw0t9EHPUyCdT/IoD6/ZolMGLM26JN7TYFrj5g/AEsEre72ZA61g7+88
/XNVegSQ7sd3AUwXYsfJgzLrmdcshuTiEeJzHME/oiFqVX0gOJLHdgk74XI/vTb7AprZW9m99HxD
+nCTI1vgjfhX1PzNL2UlPSBLqC4zBREwFzyGYq+/fiXIl+lXEdQOGPKu3qzpWpFMARZ6ZBVbsDhF
Dxlf6Mw+wmiMCmRZ3KED1UO5/bPSrc1Wiv87+hYsp+Q0cxm+8LY3i13gEdrgDbbnizINz9pmFOOh
vl2oth3818bNo+cGm6936P4pH3kA/jpC2GhpIw/YIwORedrW39w5sTWsiwaNTZ3W/rBAVq1Z/a5+
qWIT3siL7cqaVkN/beTCJT6Hw+7zYEx+6ybBWdnRRfYQ+HKyf2Y0kXUvO0ZOGd1zIUHaru4n3ezo
XTxVxV0stK3+pu/cOmbDTxjHIzbQo6lMF0bNtsad3hKAoLNNFqghVXwUjE92bNsOj81HnU9nKiG2
K8R5YgQ0foM2nuqfi8KRXvNOjwHhQrGkQwlZeRfxsbAJOB/q3RnxoPcgbVGfwpZGdnIFNP5G3Yp/
kMbBn1hSLJ8fOSiI9sJr68bojigesCIK6zZrcXT44KhdqcXQ9dGM+xM6/ZUeiuYZw20jVq0V2mRd
4c48AFAM58jdSYSYA1z3rqn1CUc+eoXRgi8WZlQeKE0ibg4iU68IkTpY9UgrbrA7VK7JFFH/jAlt
Y0jtt+QI92vQ0pzKOgbn6kYWhqNFjYOhyOuEQRuc/lMu5mGUWVW8AStODiCjOnZ6kvzpfETgq4n7
YIWlu2agioAJt4jpneC6IRi7w59xsqG79C+wtdij1HYrjRafoc5DlhGJjE8OEIY1sL2IGQw17BM9
Jjg2ZVzW2UJc5njqLGS+RWaNfFiSEYgVSHzL5u54AsI9eLQ/i+hVIgBD5nHX19Qzu1G1eMafh4qc
YcMTRT452OqbRMifYFNYWyxij/1fVJBF/y+RLeUCZhzGqqmd88aZiErN+ZvSWm9cymHuX0h1Xwpu
qGtDFuzX9TFxfcsmxZ/HVC8TBafsEb6IiqNeH/yDaWObMncDmqo0CK0Mn8wPJzDsTJVxEQLrdijL
5Gj5fZxJoszOH/zn2qvd/KYotgNLiX6YDFId49bho0Ssp1J2jxt8/kUV4aW8ij9TXcvA7bcNf4A3
g4t/Rm8JqzTe6JOWPC0fFnY7wHFcIOexa5v+Iosa2mvxg5F2sCh1re0E8iE++XymKzinsuOzEwHP
jpi1nHTDLDBT0tpC6lM253GXWREVfEVliB1tl0obuW/Wr6hI8hrmr5J1gs0RjH2ERLoyBqJP+VU4
VBxPacbgd4NNooJF7f/xxazcUdL621JDKlvYXicbtnkP31y1QXDziD5gjg2S56oIozEIdJ6RJag1
49NucModlV5K1lrVQj0xjnzNgGis4P9ywfbt7hDVdd8POCwGj9GwUw6vsYZs5sB3+4z2ulQMb77i
fcC7SAfTLWXAmew/ul8g364/U5fJRrE3MIkFX8kJz5RtVb3Od54ppC65VnfRDY/moYVQeB3WHfBV
9I6TAFegbA+B83O270qSHx313arZ7FB+Xl/skhJq6lmxuKtZOH/l46AzE/rSIACtOpB1/FBpqQz6
Jlv66DrzrFyGI12c9cvRMmX6FuJIxb5p5LbACi+vIanomiNC7SKvM/g1xEa9RcprDZNzz5qPPQqB
J8bwB0z+XfzRIHhA1HS6SfksheGJI5EcjOOJWWP+TpjrZA5KLMmU0bQmOJiukyfXPINGnF7oG3a7
5kkcF6VDLF+xfMD/gfkugUQgAGhwR57pCrFGpJ9GirAttPfTbwRYlUvZClEfeHhwoXS/vmSQYwy/
wUro//rBalVb+CcbednYRXVhJdjKb7+gYIHwl/TY9sIdpQUTddqHeZgMpSVaPbuEOUYNKoa1eKyK
EOgUxkQESsXHWaBxMxo1G8WVjrDJ6csYLbYlGUnGeRRgqDTcW2s7Z6+YibD2pLiZHlGsBte9tZnq
7g4nFe6QqSKv89GlrbK8Ip9CJZ08tr/9kkZNMI1MI/IAEyOMOwgp5C0WJRR6OIGLQVK75JXJTeSZ
LsbiOVRD6MghXjJaorStMrImzMKrpXYprCe+XGM/AKmkEOqZstBvcrlWqIiqxGRxsSNcS0/GbaKg
m0ojtbrqv1ppn3a3LX9Yrpq/xmayjrTk+WxGoFcTrM0ATxe2Eg6IAyJwTqQmUALLQP8ELF7MB+AV
5e5TZdDGuU11OwXJKG+dz0FXGrzwmbiUSiKWaeg7GRDjMEPOk3SaEMJR3NB7V7cgL5X+sF84bMSp
lbpxfwKxTwKY7C9QXXHYni/Lm8O9RcHcR1WPugpHfgCTdwMWPXZU0NXfzdkfsuXRVw4QuP7xND5Z
d2AnwqTLA7qZ4qZRZOQCIrpOEIOTaKXSmAdkEpoGHSXGY/gwxjNpqvWN8aBhpgTIGCqWXwNHHTRk
LlERs2qWDrVJxfcG2SwYiIXJNL5PBNu1dmnu/OIb5fwXgAIaCD4Aa6+fVfxZx3su8R4IsSvsKxIJ
hK8Mz4ufxU6yvMDMHwgYYah/+6i0MfYPGlFhSxUMQVRw7GNF+lvUi2IHsFW8Z1nNh2vPKNFXNHUW
dc0nU8z8VQWf4JQvmUFkWVVbB5/VQRH1m9q4kbRbJRebQSoK0TCpIm65mJX+FmXmgTLoezJtcEyj
UfhPvxyPcPTLVRlA47KPJBax7YU6fAL+bGMHpWwtUFgO9KYIubn/1HeE7Zgfbmiws63ZWAwZqW2u
eJDhDzfgC/4/4gxb3aPNX5gdXd8x2xRc5nDsM4P/KydLIMu37NsTcikYGlC/ogRfwkm+MlERaR2/
AGRtwR9soJhFq3L7JJ4GyHLlXAayZsBKM+xaOOslSVOAJ67EPFTw9oSmvGGP32cB/opiJI55TgvC
vpPtfekbt8kh2ZwKdnboaRzXsNwIava1ThjEIT6Uhu7EJvW9hIBWSxN+uVBEagGV+ZhLJJwqrcTu
/3bEWbNXaDsMzokj0xzd9QTrKNQoavfFud8HWpp9rm2DVyyrYz2XSVvorwrmDlZQ3c7WhAL76R7F
rB1uVRicBB7AvXfXag4BgyUYROIy3UxxmcKET4u2Ez4RosJXfpSXJMwJck8UkJpmjNTSYfDChqUa
aqcb5A/U17tI95w4+kVS9vXSMbk/MnbgdD+30Y/ZfMOpCdK0Z4NlKSadavUMwQNNDDsYVgwQuLE+
sFiH1EIX8zks90opJttSsE7ZsP7CfAxpZUbsIjgxyzInbPiNrX4VRqV8PnMGBQdsu8rhb9AEyfLy
OqZCUjiPGnyBaHaw6apnLYIZo1jsNM0bGI+HOJM2aGV0YOEgmUkUmTP8/T14TAHWDeDO0prby2GI
owgxa7tXq9Weg3f6CUFmEH6Wc3lvEyYPpQkfsVtS1wIomG25E2+ClluHW2pLvHmpMM0+h7iBK3ML
WNFgPst2iLGoJGgPNQZCQ0eSF0ewmiTvFWPgbbhuXs5zdwj+7QAvErpLHceMzyMVp8P4Iooi7v9Y
hlWnKaGkqhkMGB4Y7u83zf61DYOcWE1Ii6WD1Vd63/McE9aKrjie3noEMVdFCwwL7pMgUCMdmHhw
us6/B1Qka7zXKSpXtmZJK6d7eEAL+GuuZHSLqwHWu6SHmDnG3H2WwbrtK/pOSXc/5R9K2Xfo9ZTz
Lbl/OKrBir+2HPXgSGT1rm+vDSI0aXhV4TAdx7+xfhOjV384xPm2X8ffaYLVJPL6Ux1E3oAZwBh4
/8GUOv/yxurKR5kt0Wtfm5YMGpyvJEVa57dPYpintWbeywPxiWEfy6V3JqAKONvxUkqJsFVmtgyJ
MQ+grAZxkgBT9PUqCOPaFP4gg6KSQMINk+LmrlENp3q1H7H98rlZFZXYdf0lCDex+VaJTHNGvHw4
ETdeqibQlLXmOqYi0mRSk7R8XDcCa+Ov9HwYjZ5Tbe00SibljkItKNejotso+OfJHDLw3cdoKV5k
XZvHwNLV7gCOTV3M4N+IL2ox3VDI0u/o2sYiL1dpl4hWKjGx7us5iqB8rVyXjK6khA/T+A7jsQiI
htKbjQvN59s9TwNwj7CgB3CGLADHglzou1Jw6RtQhCk98SC6sjSIVHZWGIzr2sHP8l0xBPDbhhLD
PUGrgWTX1Ngc/qfj4eBuQwhBjF3Dw9PwnKYNy8AJHKjiX4ggPesQXdGfDrEXH/HV74Y7KOnyclMI
+8f4UV169uJ6D8LXVGWZBPN7zZ7yxkTopgysTPUZ6OwmYh+B8uj2j7jXPpVPZQ/+jvFEffk8pGfw
y8+pLKZlMwMZb7JmVf0TaOxPsxXZ6ufLSYSw8WA1nLGifdS7k+WBao7JCKKA+Lo+AOKtob9JZQTO
ig6zXsuKoG/h5ySj4iTaQLa8C4ey9FLWZ87G6Vij21PCsMMVpcLrBJ/L1+jexgjgeLIRcT5OBqHd
fKEfz34R+BVvJN1p/1FZiH5L2hmr1iNoFdNYFqxTHJRh/b7qVDFEc7lqUvpasgHZAH8geuQKK9aH
92jbwSJCGCGZNMIlJk5g/t7N9KYUgQdboh6NwbFbLdOYz+bZectQurdPvP0AG+j2f4kAEIdQCGnN
OUuN0rfGTTpPrHU2FiY73cJ2UtjOPcSOYAyOYyG3MX1NQ5mAI9cIjhb9CJlxKHWLXnUvHnvLCvlT
1YLYFftxjDjjYl5H/ZXKr/79AFPG5dQZbN5iglrs3IEAVJXrDrBsEvNDNBiImG+aa9OC3+ot+ljN
A0Tiu6ia1SYzjjv9jospe8owiky0ei6wSYLzC71GIAJv0A/WyCUTIZGyaM6ncNy8fg4Q9Y5P9OWp
j6STCpx3fklgwlYL5MQImgguxZod6mx6CFwA1To3O2X1x75Yah98TOP+MrcLJ2h7em16UHDa2jQ7
/YDaKvChmKddGrMuYJJdCSpWZMYb4DXvsuJErKuGuanUeiz0jxC0b6U2U5ihnFbTP9rqm0Y7R9mK
OdhWJsAXQn3i2y9/wMCSNfQ61enHEhZjx6mXT0HZdaoBkXntfKrp5yr7FG2YFYfenG3JVVUmhL85
uFHBNtkSPzMntporOpGGTk0iahbmI6RzTRpWVijBNa2jOblLxdkwFg+J+9XrHz7o8pNRRL1BED71
NZY55OZ7WGG2UVymH29ZYq45HZV1t4eoy+vNW79maFtotU77CEZf2S3FfBWO65dbxLNvyjF6cK57
dkf4NG65zaDvzp/jZ1ODHLuDaQNp7M5Gi0XIGsza3UkJIROeAf8UkupWrKyDGMIgSz3g7r/NeFa0
9MJ6M4Eb8l8Q8d2+7EehcnYkylcPkKvJpURZTYBsEQW6rrA375fzbzUqUDnHyRJ8FIBknhmRZk2H
9JJmTXjMMMfMEuye0DAWSyOqIkIx7uEgpM/r99e9Uo38sL6w3IWjZGdMc5pH44SiIUgMKFeae0zE
BEmaAXiFmXfRvDJnSgecuq9lbciC03pzChEi3OMK4YG9usOHPszEll1hcSIjaeX1JFsMC8zTUApO
OygkhX3hL78Vu01vxsy5uVC9v6h0hTR6jjdMbOPESwQniK55sE23Tp9bApWUX4Yeiny1h9d3vRo1
q33gRTUspqB1Lzv5G2gMTs+MKeqwgRpBSDAm954sFPAacIAq9TPA2wBWc2hi+4EckfvXlOUV5DyJ
Pw8osFhw/8aGTM3gTRGka0gNt0G7Jb2lWrDBdc69IQUqX0lCy7lv84mEnj/cz178yyjTPpcoKlD3
a22gvflEXX1tzfhIhkb8TL4YkbbKdemKTaIGLz8C24YzXagY7GRU6upcz9+W3ZEM29H7IMjONgMW
1srxKqIzf5Xk/rApBuTHf2Av4yZTtrrcT64ZoOaZ5JLdbUNkr0/qOFXOE517jgvSeOYi2AwJfzAd
9De8NsWflXEnWM7LphQX/2ysvv+6R0ltLYuCwjCCvQyNaXwXqV6obIHGqvdTc8yIzKAI1vNd7Vn6
Enm9T/s3ZHZQCD/CRRvMSPa+GGvMw8vK+DS0xLBWMKLjVNdAAaLec7RW8siGnPd+OoOKGqOAnWx8
hllxVWrGWO1k/mmcKeTzUgabMdtqBnmqNnOPzGuyCKMD5Ljg58kKL+R9/Kwrq5PNICGaoW1AG1TX
RkTDUL8GFWyxqtCIYLi+gEvGQsMwtrd5bWj+lCWQnZJel4urXmBgpnZscHWJBwt8CIulRBFWTvvF
gjwhWBMKhlghLI6d2mOV62vITsRtH69D4J8snsiAW5i6vDHj65Sk4VVE8+6rcsRU70AZd7pgXyMg
hynwxZM+3w1UyW1JStKkSfxTvMiwk/3g5BPcN1BW9R9GyCOCO6DMwLpwtRbkyf982hWZ9zasvMba
p/rG9ZQrRIZmVt1g60fwqaj8mKjB/CTsmr/u6ReMMAytp4YnAM+uOFb2bWsdG/IyrPh8emx1gOqn
HaTfx1qovyz8knAJON9+lWBVQu1qYywToBedK3/QEZuGzh2xQlOwIAubU4NGT7f/XKPmp2On5QYq
PfK0lPiNUvCrYF6w1OCm+i71Xmp3iNJR5LekFwuPenLAFbshYNnCiet5LfgTIL9/pfTEj4kHiFQ+
vsXTMM5DbwnBuGgWhTaRzRDgDzYMFUSTYo2XsIPFkjqgTjsEBnzMi0ZHti7PstX8/eQS4/oCPyhp
IoPn6fMgQDQOCwqe82u55TfuGoUcSRCW0jervC6g8EgehbWoRJY7h3JkwQxD5s6lrOa9OMyECAZU
P1qooDHaFl9fMAaijLaSsPxJ6DScOOkcSaM61jwAwu5kPQJPvnQpXqma50/qMlVATFc/kQUwFYTo
kFQE9jLkzvs+MdxZrxZp5UZxtj5ubjFCgj2k61PioZO/cVvUa1drIiuxOn0NGK+EzVBqmRXw7T47
XTcELeayJPO3zL19Vtws05cZcxmwAIjJjYnwab3SlQsBY1CO+tH/wSmbuYo1uF1dlIU10vxqEIWz
7UJHX6UQsRmdtjNXvYT/WXl9pKo556IeDAoHR4sKGh4W5UaQtfBitaA1kyGUBmBv1QoHPjga6BM7
PYQL7QBqlQF3zPPX/X9J4VSHOii7yvblAPOwcfyn7OHCZcjKTsQgp8RFq056CkiRamiRWL/5OW6e
NJedwkj9ZzDPwf+KG6R/0k5j4qfvhfyeL2SfLGmVmw0ntwyhpzTUZz+SrmOXTDM4THCuDCD148sk
f6VfBgcx8Z9bb1hEbUECVxUQMIJNMivQ5DXVaAMkPtjmnKuCEwPtXc5lLBDvvFabW8QFn57yT4em
762qEF9u9l8JaFVJTe7Li313XQk1qWKDK5xgniT0K9OdfAqfMSDBeGZExZChk19Kc4V3AqHhecBW
VrBnjDISyjbnMTl3Tsp6jvwtZ6zltbjCh7NIPrZ1KuyMLtfc6/lJDQ4Esq/Hylji3S7Izmeexk8R
AcOzVkyOwQItqKkHzzjlN2hNjdwINflcs1XlfiozQOYnn7cL999fMI2VErDSbGqw7/wkjGUh3YYE
4VQFE0F692+9PO2k4R4rUR9n/Dt9rmfaj50UttdwTH1whMsTnvy8xv3MqpU4oPR9PvIe04mb21B1
8Umzmi4AZCcH6ZBLNbNLoE0FoHrA0w7XzS0iSSk3l4JlQwToFWsa+Fxp2vg5h5zwrl6PibUalgq7
qWTqHj1/LxnZKrkFYAJxKKdZ4y1vLZbA0DYAm1VX83D18CYFxGGxuIEgO/wwN36OWDP4kxqi4gYP
87WdP6uL4qxHwxL3vcB84VOmcNn4hJ1uCzkOz87XQHQJZOG8Pon6GZpV5OZ6oI/rWVZqW9IuiDDm
Om+ynjqdyYeDFmzEGnGrnMPFLI3SBRD4IVPIEYR1ZR++1xA+x8cOB3yopudiQwUMzm+dqP1jpDcj
mr6vpYjpP+9Vgys/0h3uRDwc/RY8MJ0pH8boGOKnpVPiIEsew0uGKDs25lXwhuWyxvm7KtoOpc+J
xFZCAlgqjy8aa+9I/19AKYJVvv7aoFHyhS8VJmPCHIyGCkHNG1e4K3K7Z52V9ra9TPOrLyPfig/4
eDdxdQ/hKXjcqSCmfKCmX3fOvK0BKivGyqNplHVix/QvIK12N9whpOyP3ImmE2y2x6cpSQVbz3ly
RHmIP4aONy8zKIH7Yc3ns4eW0mF+pz5B1aLPoSkYx2OJbxizmKmEOrKSJuLBfMq95KS4NEQ4T29b
PlgtNlQHZ9MBFHRmBhQmOIYLlVbJCOF2qHxkoFlvbyKDIOxoQqGU3Zlk6Jy72UCoDlxpH4U/pqml
bGup+PhlCDdQeftTySKRN9S8dP48dKDZenc7enncMHhQmPj9vEn2CvdfMDsEZNwFAArOclzYmmSS
ZuUpG7s3vgcn9VTFGRDbOqx974DCJ2IFVOhfId2nIqZGnpOHeHeOz115de6R4jOn3kDXmqIv+5kE
3ymJX7yPbBsYoTtAAPO9bkJiBCwLtZ3DetVR5F0l+ec8YYkqwA7fjsAI2bHe6V/k1NWhflMqoVQs
tTrdaQ9r+/sDpk1ONwIB2pVKldZYAdxFKiIwXNLABRKweklFg6dL+U/IyeX9qy0ciTRNvqPqTqgI
XZSfy59TBroD3RagMDbI/HCcUbbDRmpHxb5YfXkys+Q2dATjB5mMjaNTj+R+AEWGIS8Z3NNB7z4Q
BpIvEt+IMhWE0Xf8o2Hzu7I96iDelVN4R89JDtp+7XDFc3VB/29+rZH1Il7P567lwjy6V8SU1C9n
ZXuUkj3SxtCRfh3WIoF+pIMxzaEhVrcrdbWEiNUejHtCaF2/FWEj3Fk/9yHxSbNF1fFKFcaL3h3i
EabyRT0ZXYuSuTqctMsfdUzqiaXHd/DN7PPw8LIQBvQ/XEamK69zU+oXT3qte5kbRPB6YUgFRJek
QRCpDroFglXS5efQicVqbyFQvEvvKvEyk7KqDde/f2XQGNSSvVRtvgvUw7xsk1/b4OikId/GtWFM
LgcUhnK0/V4y+JUycaPt6ZuWgHH+A0PRbad0SoP2YNEjdxWHKOUCwz3IXzx9gHV+SzHOf2ErOV1M
QzFetkEl7kukNPZlMHVrlrlHMxMviHBvwmgrwgJgT14hXio6oYor5YC05s8CT9gH+ywuYImUIGGv
he4q++NOeAShv85orx2OWPZ7C5vTlqLiW9nxFasnpC1tjfoVjAkudXLTXaBcA03ns3teipyqxgmp
q9UWsHem7Jg+xtAHMsvHW3Dz7uELgH0nK1twBQV92g5EblfwhU6OvkKY6y4NFhytNqKawWvOScDi
e6COe9gfinncfeaiqCVBm0r5i1Mk97g7RE9THyxtk8N+Ij/zIQsPoAElvGQNahsnDtuf0EVVNXWZ
OPAVKWBWXaKoSLri0j5/iK6hOhrF8y0/rdyGX7rBPM82jts6OwVVq8YR7XGJS6EnQddzeGMWj8SE
WXqaXgc2uFnAp9gYOb864sVCxixhMAzLVYGNSFj+6osRCFbfVoeDQpLinkQqfWEwAq+8s6ioCev0
j2Ywpi1LC0Jpqb0f/THJNbU9VWlO5RIcNnd3oKOr/8Fo/iTc25CL1785CMQ0zKXhjRsIU5palEv6
ZBxKLsa9/1SQGYxEJPP450K1l13qUIspq6f3DMBMnkTluEXPitrQtP13rj9pvLOScEvqwAIiIjte
ssTtvuWBjoevyKe/NNFddG6vjtA4dNMeKBZYl1sCsvwKVNfUZJGaSBBjC7U0sDhsc1FNENfLp7i8
uzLtP+swpyyIu8kXHAagx5suCFrJmH82jxP2/Ze+UvvJluzzkDyWmNDwTzEcxfTRcNP7IMhPLNrm
PH36pUJECoaPldYyk0XwT+ArnnwOs/QTYWLbihbQeS3Fd/R47O8n9kGQnKCfKgZwjtCyTWtwJpHu
fg1/0+ifdsGdJbELO7YoLeVG0vl+ZpjJqhV+QFw5btPzFJaft7vNqzsYjJPNbAeMhnY1hzjMVLAr
fzU6JqiWEXY+E2NYEriW+nNXM/2TeGFOlsMxnJa5UOSTHDwZXOz3/031o11cZE/8ZKv76kdNUxax
Pqy72MAFrDIiiKy+tusO9v4NXTWFJFu95/R5PuLep3QJBsT5QathMrDZ43PPVEgPkcrOwStBWuEJ
7RruUAbEYwVPWIn9QXpYeMRB/FX9ULDsMsiTcw7R4VxXJXWleyxrH45iZaRKXRRu/fmUzvfiMY8X
co+YSW2Ui1obdD6enEeYbTxTJVkAYYrZAXyerakhR/r3q/n2hVYOztFJu8bAlj5sgMZJmLLQvN10
6FtJtr01no7SbIRCjjhopYpPCOvs3YWZjYNr1W0En82ECE24uR0M20Wl8T0ykXjfqoAN1+PD6Bph
l1QWGudtW5WXQUh08962G3PxDtxSjmB6nuDYhER6sl4e9ZnqOI5mWekJ9W2A1rx5wmEyksY97617
ib90Pej2yLR2Xcj/BOJAQVMSqadY3ivVzJWpqYuIPeAg2B8o3SP9jdsSSC10PyQMO+UfXmzAi9xA
QfG23hwZdOCuOIDAXOLUBrsbIo34b3h3XUtMp6gdC5snaMDTENFLyaVdsN61E9iaNFp+tujgXc7c
lqvMC1VTc0s/XdB18cDGdwwRiOd/58IV36LzZhFYO7Vr39H1tnCxiwZSQT+/VV8kxf5ZMfz9fE0W
LxJTU2c74IbY7PFPtny3C5LLBST9nVzXonRv615KENjpGF3WwEH8xsUpLiv8oNWuwKOdf3gp6GCk
sIyKYUUE2hPYnaiQ3eMja0UBXjtc2W0Iui+Z4UpKhzubhig5nggP7BpOR1WWgzmQ3AOPRIUVQAKk
EQRJGTwAGQcibv9YBaj1rf/hHnC9f0qNz9VZMnrLBPnDZZCzyTpVeMfRPQvFE0rIsZtqbKjVwa09
I9Gl7WgHMMNBZEP9C8Asg555oOxdVMHszFgTCcfG7SgijleYR6Zdodfn4KWAPBpu8sa7WBlpHGda
5Lol5UNxocuXLmMPG0UWhjEwW1K/IhgRdP5a3D8eoKDCiw+YxG0nMLuvjsq22XYSW+uH96WMnE+B
nDaZ55jkzGsKx4RU7dWyZO1wIFmokWXujqmyvaLD5myoIJ63jjQGkF/Afp5pc77bgvUma/oVMzss
g4fJrYZUK0yo1SERuBWuwVb9/nDy4llSoaqBG3yiASW25LAEV1FtURUKzZDVQii29RaglgXLl2iI
E5BeE7J7uk5o5Qob9D/hFnYEEz8XeIA6oIjZ1kUV3NGL1O0JVUdnhmUHX20DwSqO3nCUW/Mm0hcN
0Xf2/Z+cneZnn8vA9MaDgTEOwGN5sosJxLDV8qOuXehl5DgIcdPO1mJot+ikzJLiGYL7QQXLwC8Q
QBxipza76j8OvmhG0C+CWvKeUIqcg1vtTkZ9hzFrKrKhOwSfLGcRneh3h6zAyzvslTMGnNJt6jUL
QOoEBGgdKTBr9d2HrJOynvtUI3HBLHUHq9G97MFbusThRXPTEMVKEmBvSw18m05Lh3RQ0TTsizij
FzQIoAFkAh1bSgEmmhRkIu9yEp8+iuVUlCYnVWVgEJpIehobhiPU5WmfC9KTrnECgMkgM+7XoJnj
AcH0/ItkQs0PfLxWexm0YQNn2dXv+K9FQBVIGvTziRMXsJGa3GKjYk4yWU8KlbKwz62Z7eHuiKOH
5k8ilSgZGamoVq/hSOSowtqLHx00gYOB+DY5No62CRygn1xLpb1M/sMfxhbSnSyW0yxyaTucceAq
GBYt2uLplyr9/YMBmeCkDvzJQ2tpToZC2xgElAyrdCL20bA0JtkdogygKpsh7d01QqC2TRapinJ/
1NMbn5u5sMOM1jiJt7Aji69RNUvVVbNi8jB+f5yZeg1GHUmM9dToWOsYBlAgve/zdtTPqlQF54ZQ
I08v++X1j3vnZtzcukjwLj0g8xO+FeolKQBBbsX+/mawGoQWuYaVB14G0Nn3QFsRD5VlmNPGUAjJ
aIQBqFoZ5nbBzQ1p+/Rc4LfmafO+Gkd5huckuAnrw3z1dD1GUJ3pif7qZZ8DHnVxRlVa9B+693c+
W+5PLVZdvOxLeyNBeiRYw2pv2dMQzH8MVPPVAzGiMN59pkKuoj3h2MGRr7cij5msc9yTu3ZRNPYO
RHqRC1JIBq9cuyoqpi203bz+FoX3WeFaqioDtRazLwGQLuwJrQzT1ZIVfVrHDJ9WOKtsIotOMQWh
F1V0MvyN8+NXMZMqStOmn9Y2my4btxUkJBk/4dY9L4vBge03Xus/Ue5QGGpCLfOcN1Vs4+oLxhmJ
vpR6wTmUv7dp1ThRcpeLYftHF/LHCugLLN0tJa09peVFgxXTJs5Fs3VScAO/aGuzXVhFAdbrzuhj
lR2k0jiahnIw+SGGTh7q0UDnWluDGJ2yL9ze/4bQJyDsQJJnYaj1hy3dh0jnWwUvHbYLNZaa1osx
Pu2k1GPx4ke1R8/Kah1JKHdSCcCWglmWOQ4ICR1tIbLRvnAIH8KfGYE+QQo6fWZ9Q3hTttPWzLRs
8LAlYSsKOidSNb4KrlMbaTzOXuielMKZbRmbIzkSM/m/WnJLF/snGEQGh8aJiZDR4OCP5zWvpqzI
/PipaNAaNeUUowRFBkwDSq0i+hQpr95jOw+RkmOOlcXOOsQXilzmEW/dpXAwsxTM21taT+bXb423
dLc8oonBGt1Tl4bWIi27unrcdHQ5Hnn8ENRpy3Bc+iQ/YW7A5GXtiDns19KNNFISErSpISZ0R2Yq
D5ARLDZkq8oxcGih1a7++6wpVqv23XLTVKKjcIkU6H85fg0MgWznz5P8DjyUMXWufYAD5klgSsXI
P9e7sFdEp1di0LL9Xpd6WVEsUFc4qRyo5EwqzFgozOPhAtxy+eMuetumBEP9eFq9D5Eco7pTfbcq
WUF3MiONobEM5br38ud2VavC2Zn8kxvzJO2JzQpPZZXIL5jjU7LN6oLIlJ4VZakTs6aZ8cHSQEsZ
QVzgypfqlRQ8A556iwoFkEYmEkSc1l6YKJkwkqFqH0t/CWwsF1VkLCNA4YmHgIEZsimmDd43j/Pf
TFei08Fa691GatBSj7kBLJ/i3sCOYsTSET9MjEZMr7okJOw7OgQkWjxwZqHSRLeH+i4LTLSe74G1
SZfJzZW7+BqxF1QLCTvzjcR/ke8yzXWX/1gIBXAMXxgQ1M0lu3wr9+zrIbwcc4FG7QP/bA6e+eIV
kBlHvxGaJyVNmPLdksFY7byybAlkI+ga04dSpISasMfqVDjjJQ5njXAZVamcZqIna/LdUSSJ7HJQ
CBEksZABJgT9A+SA3FcR1LUv90mBsWRAurls9KHAo4hpBpyh/orOgL7eIEcjzbwTqYrT2/JuzRY+
lrqfped3Gh9VtK7vNkQLahL2eLDQCpPBzsVntI89ieDnghfRYJfgM2qCm60qI+3xtyfFO+6uWr4x
K/fTQ5QY8uHZ8YSY4tYj21LdsJdPteoKd3VmUslidoyTlRFx/GiNIIhqqVZsDIr/TqEM0O8DB6Uc
WnTb8cb+3tL/uXdq+8Y43KQqcy9GQJA9wQ8XPJlk9ASvKt2+7A0sdquR+4hp+1oh1OTkeSiBzzCV
TIAGR94P/1r2G+EWzhfWS0q8bdVwsQx8w2e4xf2SLsIdTPvL9M3b3K/+8Q0aI4oxcg55neomoE2P
0GJ04AKWMHUjG5cUcylDqXSxdSGkVPbT/p/7QU9KcYFjIPysLJw/AVau4QpjJHYycqqkI1Aj77fG
tyvexqcPbhwX+Um5DWrdYV9HijHPrFWgQNcmZfB/yiv/UrvYvTqe4EAK06aXdOFSrycd/kbokTB8
OFeF1U7urI/smlCxuUkb+h1dbo2VGBGJqbxeSbWvr+rzLE3OEKtQDPH5s4urYot06tdBSY9HbJ3x
O4FTf2fYMpezPU6wrWgdSjrC/sJEvpLlXVFE/DvVaWNHZDMBbVixHnkDUUpcCCxqciEsXr8ws9Lm
lMb+H+XoYg+vSMgzYl5K3fHDWQdXelestqYq9t7c3UmjC/ntqq1pxGBcScCaosaFlv/Ui394d7ug
BLGNCDulwLH+vhrKNSkDEVIWspVGLNRqCiowRQ1ETqqwtjblpCr0gZhN7/frp/HvXTYAQdMjD1Oz
RB58mZYKg53s29Q8Fjp0pPmCRDn1zx8Whx9pTUmauiziGo6YLUcvH4SGythQ2wAANFr7AtqGymzY
JqFj9ncyPTI5ZRH8Qt4Qs/lrhL82aPD6L5M805r/q10GVYnxwQQbmZ5iGf4eGWwlqSQBrBsOM690
UX0yge2K4KZSUSG5OpxVet1FSxqt0go2AtSUDz7kKwjz0vFxYxmqIjS7mhe/rdC2UZ5arSPgVrDg
iO5pnvUtuqWAYgIf4GTd1aPgn3sNy7X9RkELnk0phtciLRrA0Ov9H3dJZOUDPIhhvc1/g4HGIoKH
p10ndybHL4XrV6kYfoeyTcTQJ9YOdw4Tqf0U5WkmU0gGJKm+X225w34BNlbm0iGgMTnK5lJOBchH
XPCC6Av+yZFx5G6OoDKMJBpntcsJU8IJ9vGD84ytRR0mnPRZPONWXNFHBPEZ3vGWQFp201XHpqoM
k7xpARKgmSwo/YG7mk5Y0TGgtZ5v0GUbQw057uWblBm0cTKlvGroM2cNKnkX23MEy+4d+Zxs3QHB
j/j25XwMq/B77Xx3n63DbexaqadBPqjIJJ7gRqwEUks1D0WRcMsaK9UzKUuFIrGnG2RfFcIgQn4r
TcP+8kmSB2RuoCdAz7exwTbR/vBD8fJ2bqn8F4HXO+Cv5d9jcbcw8hl9LDaYw+mrHTBlckTF+k8c
HGRM7uUqx+/ItfRT5NzTO+Hnfvp+zI9+vo+OGUxEsZjLFjBbNim4fHTloCjz7moXoh2wM5d8SnNE
PGrIxrasveWWCJVbJsh9OkCr2kB2gUq7ERyFL7b9nFHT74fTUVd26tPo3m6gRqnUOhGCCd8FeYJ/
ZI8qRFOMkS0RO1E/ZhjuiKH/2iba9V7mUqfAZRTGCtO59iEjcUzF5SmQHY4sP9tz77y2LXihnOLu
Gf2nRuxT2Mnc6/rTTufqNmmxF12oUME6mDk0olG7IM+f6dJPVJ7Om1L6HDjO8wkvaZwC5S1XLA4o
FzyIc2hFkGHpasMqxcJNWai8/ORzD9n3NLhh4mfQyfzF0HOfgXXPDnHl658u4/pl8acpdzt0PbPg
gzB4o/pggwDLwFEQ9WGe0myJqTYECBMhBWwUKAuH952rd/A+9VchG7DYblonHQ7nnMFwM8d9vHJT
qASpTpXuGKzU+yaderbn/ArLISZBP3uu/15Nkc6POZwXxYh1LRyTmOvFLbjM05+gUJvvQS6DFoWQ
ErqxPNev7zo4A2wx7o24c4R8o/UpeZ1XHa+0Lw8qwtMfJCuuafSnKbp1f3cCUBL4o5wWQ9zSyFEe
FYKrqjAkjaWOEu0HQU3dFoZzt0LgK5AihPVfQk5B7rdHRaWpheWCVc7LXVAsaoBTeVVhSZfsJx91
57AIqjAiksie2TuzmMj1hrmSsR76lpoPaCVxT4wq13NSo/XRiREjjtlO1A/MA+8353b+nkMoKzVE
sxEvYPJc/dmdVNH8F4d8jf8z0cGmV8QsFNFAf70SRtE5Wl4yHZ+2xQXMVAutJK7sf2xLaARAlIkJ
Zy7Iqd7DWkdpZoebrmPJJmYq72+UaEfUygHWu2I78byjsu1X3nITQqdAhywoN0qHGSf8kTTGl70Z
F4o8cwLMxECuzgM0ggdbSuqGeF0sBEOngIkzd4HMSJgSiSASo04nf2qyvfPEbaBStTqWN8wSJKWs
qaA54D9PKgTh/ALdpYdfYfDhxsQlUveTK1Aa1jM1IGgoTE3XatQ+xTo88uwEnby5LzDls5UaGSrV
T7eo5hh4xscSyK0mz/dzdC5GmjW++JyH7651A7THYwRfTI5XsfPXZWM/dM1nmLiqtHLR+BSWpB5j
bV4VFJf99P26Dd9r+bjCnchMApDOjO/OibrjGk8lZgxjSIv7OjecSXZq1/mfSZSrmhSXTfMcL8Qs
49kHyJpGAtbx9xUe5V9ypkQSdyv8d+2DWImBBev2CRDgXod/q75JB5SoNwyv9DqPUf7kyeZRKwqZ
gYMz82RLxQ4U5Vu+/OEgehOIInq5t6u7T9QfwDNxHOi8rapNvayx+MPjDu/sUQzlbaL61nUE32vO
8QM0sHxbc8mfeMlPEwqIXSUNasbBEr9W1SXmNXTsGjAMgSEV4jHyA5wBK3p51xnQhgqwvBHVDaQy
7EFOnz80zlHiRJ0kNpP7EEKa6nwJrpdU3OVOY7ucwqC4SHjPnBcRLRlfackRGrUyMAGRqfTacNzR
yaD5aL50lbNfpGMxqSqwcKVYrPQUIzPkT2aaBkjovHbsruzIkvMCBe0OXdxlWjc4dpqkt2W4MT/K
obNw6nfeOKdh/NMLKSbTlGEfTfdF4tyaOyIeEpcnSGZmlatHWYHK/mX553dZCZc5nKkmLmTq7qEE
7dyoSNcbKzGlDiEtJMy1fuelSdLfNgB+EwQmnnPurJlOH2QgVfasqaPFpuLx2XyAMI/bBsxCrYKm
oIv1l9vwz5g3E4y1jJT6NtsGgAhyoqDJh5D4G02XJJdqv7GRrZVpnXfpk+NZCH38L0bxPnXaLAOl
R7UrvMT+Z20FvDCqEILlCAdrDCgUVeNjK6/0/A3My6p0v1Wmm+K7CrfOijX/2ry1nCE42wHMqFk4
wLuP5KF60yvWo9/P/iYw6U9AFFMxg/xefxf3IxeXIivvV8Ormh02rD8GqUZa8oxbR+4ohhUIKG6E
6JofbXtTnP5fb/F+8dj7dDdf0b0cdfRZ7+ntbmKYU+luZ2VuNMRRrRbqcO0TLHRktJsJMn/Tepv5
YW0nKzvSChYthwrvMfAQ4ptm8hYGPVE0GlzDe3Kca0+loq/wGe9qSGS9xmlrqgKOFtJJXPTYRmph
J3jWa0ooidl+5v8xtsFZh6X95Y8eAr3ICq4TfGdzf4qQdUiGWJPakmEYrlxOakFJ7ntUYmrLhbpI
6l8FuKRhMUOAuozpJYrrKOd/a68hXvwmRTXLYZTa299UFFslZcUUe/I0Nd5N4npmDtipC0Si2wep
Zh0AezMNp6jHk/HA0gGzXoJL9qqIJ7JVX4oNv9I/Es/ZclXDOgXjkRrwj6OFRRpcxaSRn9wtR9n1
NpmaCLrDKxT8P7h1FXqb6i9CRVAd9/D+yvBG4bE6W87gB7jswmKzsWJXGHqNP21ajyAQHgJyfvYV
1uXQNPX1MjL6fgB5YvTQ2ZPgfO5lcALWdah6Wdtpv/FWXgpPTzxaTjAQtfsWgK8GgnWz/lW+AzBj
uMmUE9ELtpp7L5FhnPnnnpzRfQS4h01qtr75ZSWGgBqkUyydZz3ta7RStCWySO963ftXVu4B8sjE
DnUQMu2nmXdKv5/4qX3x5nsBFwulyQTKTvmqBuL/BRNL9FsV8AoGYG7oin99tjlM+ZZ6/3Vyswpb
GHRuNg5+8XZUTygn3RdeQrmJCY+/dAQcWGSRnhnDH2y/+71qdLTsx1Lpd+FV5jJqVE5tqbOviEpu
lhXBP1sogJBN4UtDOxTfPBJOtKOl+Zk5A+F+GbsMMBkzOhe5ldMBoMPtHxydlHOJPxaElr9nxSk9
6cAf5IVZRYq5dPmIxtD2mbp1yvdBaRoPCcaLx+GbS9ZpfWSmiaBj7nQ+Lo4PUJ3mD3Gwx7Cs6Cub
v45DDFcTpWYAXlm2CnmlbJlC1DmvudTLq2gafgMCD/AjWNVu/KZoas+Ozd7UyQV6BBwUEv7KuKMa
TQJg8aVxCDsM9g9+DYo78wgr0u+G/+hWIUAN0MlPdH3wrfQIzfK78zKBCA6v1MiVw6Hzcq08nNOP
x3YQPsAiraOtyoHM+ziIZGmeASIcQMveXT2XlmwJzFA2kipZR+ZWHCgHhX4vtN9QiRrLZ4pRgsXa
gD462T/ekktCOA8A/kZSTtfL5NCwvKFq1AFBpJUbTCyBq40irhCsD4Rv7GsC6dDgYTQczVZKCV2f
BrvntlCs1opsFf4UNwyyYklq1SY+xYKT2MeWh4HuzMYD/YMKxnuAlsdN1d6Tn4GFpvzWSf23AsEC
dmfS9sicozJdqEAHFSaUPvDIPJT5jHp7sG5zgCdb+BP1c8s7dDC8fAZi5JZFYMrOAtJB5fMAVzSr
dgGFAMVHhp9xGqGgNoZbAGc5+ynn836CVeiojfujEI85eXSFmyau/F4Exp7/Mba1LGAbIaPzJ7KW
Ucr4uPsfk6glNJq+/sjrMDkx/2nv6Wz2J0R0/vgKxpt99J9AjzLymvWcoMrwq+8GIxGqQE2K0N8U
YewcmvbVfJnOfJ1N+sNTCjuyMguHPNw77zWutWyXi3CTU/B1WDlTW9RL5FUcuqLsSRm00us6jxCq
dELRbgnFJt/m9euR1eIcXXyRcHLm0fY/kRhQSIndAsCOxZPezVoy95Rxx9NWrlaJrhGf64G2YhLF
RHq4l9bvg3QoLyqgHzOUKOc0U1AGaJhUr5AbZVmpqF336OHP7WGqaPmS+HPqFQn046r0L1G17heT
f8A+Sb20Jv0x9hmt+kANJfNZt/Wf407NgOqy2JyMWU6lVCWOPYBuT3uhvdgbFww+/GFoIveIaHQO
ehaLAnHwaO2JBC4puxLzZobPU7In91fNLR0Ts/It6rGNcEcCW/ufwq0cb6eNBhjc/iuqnGIjv89M
6R2M6lAu3ztF+8eZT2EWwRv5OzJBZ1mTmabFsQOpHW7orehyoa8IN+/kD4h0/Q52LSVCOuI5wkn5
TSIZwbR5UXs8cFRCiaEEoub/PPhtsI6YmzmbgfPMw9Grs2FNoF1toFUME4JV04rY8HAAVkPdt60s
Sm4t1VjdCVil722G3fycmhvou1B05dr/AJe9nzmFSqeWiGz6/yzK0YJTUHoh3p8IZmziO6j441pj
6QrzXMtljx0uptpkbT+4CdddA/uSvU8g25LDhx2gvbOeQ216v9ksXv3nl204Nmj4YX03Ck8indyP
xyC8Frk6iZrd8an8N6/pPYYfzh9FUQad26D7GYzCTYe+O2BT1YvWQkj886nIsDuX5kZFia24BFjX
qnCGA3fSDUkRNgDZxBai+hyCaYeHjO9OMGpGff+2DCgGMaLTYYHLkueH+cm2rYpWXpVpG3aDdnTW
CDwXUE75dLaWuVsAxqKloukQwtKfRMuYl3A4BBWZlnW7QpSwzsU5h0Kk8piPPZs5HDFMdbQYUrIM
jgppBLFIvohNIQ1dv0MDEjXhqIUHGT1dQKs1Olll23+SFj6RYG3szpSb7/YZrOxkj9WbE4HCRGSc
zPVv0rgDDdhZB7G/3847HpUOeOcFLj44Yz/+IpfSK0b567sHis37jMiNCl2x/QiI2XFqb4yhnEJk
3tkV71WK24nMTlM8rtnHVpy+X3mwAKzrZjnXEvtZx79KtZ9DHzk9kqxX94gWxivDeWTa6e7IOMR4
jC2YdtnbORXE38Y3BrmBJyeQUBNmaBq2RDitEa+lu2bothNseuo7vZ2mT9EiKRri52iTuuSexQLL
E/1DYj8+yTirOP/q87lko5oCdwLionIFy02lIRdqjcbVw/nXjQYkn5mILXL7/DXcyFyn5VlDDki+
a2BkxDcklNuZrt4l1cVddVU5mvehHkF615PnsTCH6FvOB23DDRorhldbWiaWUASTJBcGuF1Aa7aU
0d3px5O2Ex1zTssZRPzU+4uUfYAxngtMBwIOgaBlinY4ePNmvjkyYQoaKG2DyFOgMqWBRgyGeWis
Q4rj5DNmqWYgzuidYBWl0dTTeSRkHLmA8yes9QwbWMtTzfGe5cFzx9rl+EqUVQDrZVukcDNtiZn6
SjI0p4FDqPkKx9OITwD5GJbU/B/BuWbP6EfBs8NNZ9ymdrKwFm3H2VvUOQ2VNyDhzMM2M9dtbA3S
7b2/gL7Z03qmpR1FOtB9zEjX/mV2ySij060gpUu9fu5vbrsOnY7g/qivSpvfVyWH7nZ2UE/0Bsw4
vk9sLZ/2W6g123uuE3vH3CXMcDM/nJA/mgNCftGquz7SzzBTinLWe/rbl8Q3Ol6qRRWtrCHBFjY8
wPvgSqdegEiec/YwhOnevjeb+dPHhAHc3zr+Z4VgFKOEsYyo6UuZ5DtHUY4TKzWwMJpR/oSVaM/a
Ax2RTLYP4/9938Z3qC0nqyi1zsRLiXXO9b3H6zWxb4nTVcsoJTrWFpjCJbpCM0V+a8mIWqRygNPe
Xi4cHpAujsPRg5zSQ91CemI15LC1RskVIrbGoW8f1GuqtSY9fw6L2Gr1nGkSdwFNYaHui5NC1LQN
WiSoT7L2s/euk2H07RX+8Qv8xhCfIwbOhHyMZG+sWipcavFosf9i3PFNG8K5DwE4oD70OlI8qtbk
PD08SBcO9N4Qp8a2a/mfO3o+Oue+NwQl+lrtjDglxBvkGMddvqzU+QTXETMVJNUJ+BG81YeA3+lN
UesQ7in2dBVTpK+AlgWe1m7+gkJmLARaPkWjykHmtmAWjLF3VUQz0jpaqgaPjbQLtfKOxDJD/8sm
Hj1va8mBqzxy1OVQkRimoUKNawwYV1px6Xt8klchifh2jFirrgCvmq19Sm+CCenZIDWMUaFpXrS2
GtFLQB5jauAYQQKD7o0MGbZptDrBVRiV9zo0XdGyiGHzVE4752r0Ew7hvDN1M4UfdLr4u4wdr5l9
bwccHUoRQV1rdoIoccK42uoqMIAQNp/t+q24lE9usdFMZFoaaHMNty60bE7duneWUbQDKIJKiFJL
j5+vs1UzXV3zWhbArUOah874khJ4/yV+0goRJ7xzHJSfRmIxyXTrE+Hvu3Dks/PVXZ3bujLJ42WZ
Y0kZASR+zjk+iWnCee+VwEQ88dLc80MXD94a6GTsUupAX03Uq86i22COSiX2dHsQqoMtKEAbEdLA
eMrdxv+vd2mwc5TX4xy2d95vNuEsOKUBROEWJj2dxCLuS6+RlkdwTTd3POw8w4a6Po0WwlKodPhj
27I8rJni5FkeFmUByOEee+Z7PTaEVYaDDUXDuGWE7EZ39GXOP0mEhyW6BvJOhmpA/BfVtdO3klSJ
8D3PsNfD3zZMTQNhbja/BwhABIzUceRGnQrccja62auVh5WOyT7aTae0PxeQEE2v3j0P1wXqwe3l
xGyEBgJmyTC47tw8YeOlNHtT2qsV1v1z8nQb/YcEaC++lxxVxythqIfmgMf3A1YpPjJqOI810AfX
sKTUTIgdOUHWzMHJtZIrdM9dJI9tm7pDofymz34oJFXlSJoNUsxcMX8gX/Syq0MnWFw+YKSocDb7
SrwMscQIw6CKPoiOIKGPNM+FDeb9/e6g0TJAXnEl8jajtR4TSSKgchmVDvodI/o3W0RIWH3AmQGq
EDPj0giZbvQvgSyk2kltqJKsKRtY+O0YVDgzdT6sT3vhYg8hK0+86Rt/CCDigSLqwDuogiM57+W3
Qmn3hDoa5MJq3BZDIYHN6P4kWefZh8PqMPiI0XJx5MzwoUnOpQY01JJUfzveFmhSTNuM80Zglnlo
z9OtgKEPwECYqwKZu/2sIcYWhssc1YpFppX5njReX8g/nZrsPXwpwprSQqb/JoReW1J/9924iLgr
rpsAgXo2Oc85l9lwsjEv14u4OgYbgGXc56Nr28LwUMxqiHqMpy6Cgak99woqFlSDxkMbkCvss4uB
FZAjOSra9RFTJsvzzMy3XQjEu7ugyiRq45E4Mfpv1V0UBMSvKapxW68JXG9VGeHvsR7emqhcb/N+
RRWpz7thrvjBY/7/lrFA5toMbvMQO2C+EoqdoBDqo3muKnhP7jrjPyc4P/UewXW3pPr0TkgKq03K
cz1Vkfc+75C5aArvpSFTDbWCG/niSJQ+yjRMA6cw0IoPyxaDUaiKSRgr1Tc3BPki584bZgLW2G1E
MSc/fw/5qDHp3mJ1QFyKtHRKq9lwQ23oANErCfPkVSlXFVTqPFMKcLVIy2sDTUWWbyoDEmTrhK3+
54WUwqgNTgJ9UBr1kL/2htP60lDm3Gh7U7T8tmkM6LogP0Zjzvz3h2R0/YJYrxDydLtmHc6BDOSu
h/0Vq7fzbPemhbxUfdmOvMJusPy1EbuOfnmXgGWKXdNC/DRobSlu9K39JNdCj3fcGWSB9GGSbKz9
W8dWJ4XXfq6vnWQPhl/a3A6SmWXKa5twxWeZJR5/sAHpPyqfcG/zhXl8tDM7Dq/NdR1qzFQUyffj
F8KIvZhauBH0ExHNPu+vT3uUU/ivg0c4jTtEleZRbeJ199V+qyCzq2/wA/q4ilChuFcMWIPMfEgW
6SkZY1xCc6JE8dH5DUnHvFVa+3GxzDq26Kft8IL4EYbISk7W19n1vUVWm5GEh4FDfyw64e6M96us
yniC94qwhBowjCBwpG1c90lukjRAZj8+HKTqM7OfGAvztLE6qLHzxTyOCW7QMq48gZTEfjycPWET
100/tVoUXmVHbCz9NdCMMs94EEhPXKWHSeSYxkYpEYYFUu5hjizimzwD8iEvx36AfU8zPKR7zv+1
bWai3VeG7fsz2dhomKpUt0DLRO3+uSAHo6k4cF1O9VMZaB9iv3zD9unD+NxiiVuaPTPghR4QHuKr
D4uWx8+XF5V0ByKRk/OpkwFTwTcO2dF78hpm/5+eVB8O+E5KOidJJAlCuOubnZlkYnOC9nkMjCGI
vbzVl3Rj4E8707qIIrcck2eIv9acyZ1BgqWRtoeUrayEZUs6lxAbGb/UcPg00njyyqvn0fKNZSTd
GX3Nop5MGchpiOok8YW2vYzwo/s7PfFPO0Ce1S/B+Zbo1XCkUYGDTipw3Zr4Cc5PKb7pYVjSDEiY
9z0Qm+Tigvql0fEXLUDVpRG7zPhBaTGlgKj95LPqKOrWCngjl8Oy6+ancALxoMXtyeyt/BxYYxMa
6dE0NC+AAhA72chpJ9Wz5AzgW3N9lLnaxr2tSMLd5Zuu59AOGFQ6+Zj5oofPC7R34+G046q/GU2A
XFXcWTE0Cj/Vf3Ujff5piCdFF+ortCeVsJYeGhvR7K1v2Ut1rKavb72oQrk95MzAWbK+NbrzCNth
z22yw3b5u0wEOmjZHVSY9HGVvcQnyYoSVz2yiyxkdd2ktG3s8pHYj0qXf3OCRA9VwDHiTo2YyQIf
vpOtmBFtj0wZLu0a3fZ5xQIE9LkN3XGL1tG6wW4UPvjWCuGQYZl2yj8f/wKixxV4Dvs0152Dlo4V
3NXyP17XFfNp5HeF0UeT0YKDbjOShBAmWMwfI1N6d8eggOcG1JBBtlRcTUqkvOxrX1JPJuvOkcHr
uBeb+I5y3xgFSpbVBqkCqEvi15YhB0x1o7ttU6zZ6QT5DQrf3KwX2pSYsQVEZyWsEoZKTME9BNN3
Wworb9iT54cSbdLBnLKiyYA3h4ScLtSHOcyFydcKSnucAJrsAl7Wy3+OGPrRnjN6tmZ8+a1jz+Wo
rRBs1v4loiNsABepM1VThrpTI0HaKqKz5Q86YsdklieGn8jsyT7VUih3oeT5odKKCatCcc/zdrWm
ollmLdRO4K+LoI0wbtKql51LvpvPQP52i56dPwgOwiMecdqOVXNjJQpIsQuYf+WJAWYuyVxC3oCa
+X6HsdyLq9DDF2AQNmuyPavorpInw6YUdv+koqybBAVtQacc376Bm3LeVAH3enc1LBH6wosKF9FB
2DsGtFZ8cxusu3CQYk6XhaVXc97yngXiQvkGe3BrSWWUddiMb6RXfOiFxe8NzcBQwnxyfweAgdid
LvdSTT24eXhDwvo96DW7RfOIOl0yH3fjWWKLHqWT7V06Q3Il0lwdrm9/1vdQBmyKvNGLYTBlsbCN
OqcUBe9isX0M1t82ZiVokKd3eOdB2hFEbzj9Tickp/Ovxr0pg1e7cNkmJGQ6mnvNoG1Cryxpsr2l
cCwZ9g13JncjiONvxkCH52PaYPGl3p6aWuUpwB1ft0RV9zOSxfWYIHk+1g5u4rAkb4DiZ1t2F//l
U9VcN1IfKZ30wueBYs2O3SqkaWBEvWdrk6lqlr/wd9NnBWZ2JwXpKARjq3/ub/ADwLFzNOz7j5an
xEmBMTrxF5xtoy14lVpqQEC3cG+3sT+LDQxnoVIQWkU71q28OR00w4Wr1Gn4SsSNDLLC0Gy/yHtB
VEWApC13AShNHb7z8PpFFy8xZpMquW9+nsCVNQRdbEOBV7AXLsW0uOJc12CzoAKhIC0a4l0OSAGm
mhvEu7PQhk4yU5rtWNtJLkya86pVf8zIR1g/GIyuLLrOmn+RLM5UK7KaKIqbT2s8YGqhoLHLynGv
pyqssbT2N0pO3JUPWLpBarj9Mph4Tku23YYMWyYJFFTdR1p0BzoEeEVWMWQMn9dDX39CHYYoRXJi
/Ad6Q58EEZeQxqdI4VELB7XJgNcD3lBOZODoHUYHs8Xt/5sVSWDM+udPnzi05jopcoRhUAFzFygZ
gADshuLIstP23lRziueSJHlDFie30+9ePeAGNAGaCXTwPW868yPxj0WwcoL2QeF1eLVWpvBhjSIO
ILFmx35HAPFDPxQ2sVEBo/xUUann36XPS6bEL8/3/TpMEc3Oc5zIEFFg5mUE+A2UrUgIBsvi/Fa4
92zr2ud/FV/HMXvP9AfY5BDVEJ1wo66nlICAezT3A1MsR9i+pNaMTkp589nMdg4SllFqS4BhGbQg
L4vzWThFUBrmVvdLvChXHSKBAEZ1t5SuiQnNWJKRqvxCsMQZAmqGfWmTnGpa8KCax7Cjy3OS97X+
ozIZjC/ozr7KXacUwpstXY0Z4OH71p/SHRoX+gDqziup4DVx1CWHAzOnW+yVBvUuNOV8SrP5oFkW
HiPV47gENivMZzt9RNZxUS4iPnDzw9rI2az+bSNxu+8OS1Q/xCZUAIn/ptys3cLSnOHScmdF20VK
+Jq7lbMn3c9XsruI9CQRUOan/4v0AKsWEW2pjLROoMmK9wrjrC6MBtdQfiBhqjFT7xtUeVa+Fqr+
fPD8Y077UmjVetv63MaVAXxz3op3Sy3PK9l5KFu0iQF+yUXmAQyPMLxeJo3s/6+houtJuCI+M6iV
49w2NSZFVvAQMDVv8sI1HZWorp6IS6eKXPDGaK21rLQP78OLlLiZgUeuwfqnKj8o5+En1VB/vk+b
jzU4bW0O2Yn8zYjB5qx28ROpUnW+RhLbvQKaZIqUNJkCKcNPXwDDEucgfwvbVGEftbHosOc0hQje
5XoFDZctkLyE6LFnIr3jtfAdCkorLz3FQl7IX9+Bx1uLctx3qk/NU1V1GFANlF3rdc+8MCBfDfo5
WqGh1rt7eSkaZb9GypXyLA5duIZQICYxrDzymUf/M6p4kcdgKbF/K8y+YIojtUNHFtiog0T0jgAZ
T+q04lMH4lj9CFxah5Qhur+UNbIRp0H7ZZ97Pb3mFiGX73yIwodXzr7Izn9E0jCvU2/LNUXjuAww
/cN84ZJey2/BUdTFAe6B/uk3Wpu77faVmL98360RK9pZ847fey7pQsdfMmQKxIVaI67Ep8eRntDC
31Lao8QQ+OPdaMwqXIYwNEmMNQpXMxK8NoQU/w/sljMdpG12J6OB4m4tvaZ6z4jC7dkC3ChfsAor
sGJvq8/YhzzjYhCa4yZdXWQkFSVJ7IRLzpaL9WDiu6aAAU0nGr7i5Czc+azvs7xm5ImMAJUHsvFd
Xjg7qb1j8cxn53H9CvCcVSpCnbJk7SGXoq6/r2zM6uDrUY8fWt9aX9iSat5Hcy8LE36DeB4d+JVg
+qzdoZNYTs4gYF/JJzRIW+3X/VHMWueFMjTjlSaTPPpoQHV5b09I1eLcyOTLB9LGME0mQ7S6wKkG
bHF19AuPL7z5XklVrt7wNjOoRjD1g78VwT4nAq0RcfN49SSAilqbgyWvXhoagNNTzYJWvR7NOatA
pFjrFqpeTuPT7WswBFCAEcl6Qykhll9r5PafMKXGmC+HnnsbgFvj/QJ3AMEPV1QiR8oMpm2vaPrc
xQNn92UuG6V2m/zo10WWvnp9UJ14OgM5N65B6q8cgRyM/J0wqIEOwN1D2tg3P7lbUwckrVZsoD5j
1GKN3Ddz6pGU6OgFysbLNkdHT3ppMvWPzwdijgzlnTUFZp5QGMq48WwI4vK6irGJ9s0g2gphCBLA
4VofpiSYJL7Aq5AayjdPq60YnGl6PF6zM/9m5NOEX3Kqzk0XxzS5eMVb5CHaZP4/f1HhFzBr9CX3
JpmIlwlWf8yFD8TTcPmNXz+9TavYF6gh+2cKDIom+jZTIm7krWi1j1M6rGYKt0S8htUKSto6zxKW
V402eZBUbK0gOsJKHlRrGivEvvDSDBL/IyDigQ37ZTbYnis//OtpAcRQIaD1rBnuJw97lvdhJ0fC
A5wp+iIKNHH/GvpvNDzQWAdPkBrJNVEsTsnnCZPJcFwbiDDxshuaZMxilZXjoY+D+h7vog8EFYYQ
S6JRRbhl4Hi5jrnt8ePm/879TCg69PIZpC28OMcMVfkijc8sTh4k7UeNXb02dGksalqVNy4foRod
EQWxGDjPQMoted0wmGcb/qhrN3yLM1tWytF5moeRTv+kAP/eR16Ru/CAC3E8Hz7f7eBjxX00R64z
LBM/rzJni5DS48hCx1u47jEna86YxwttvijrGZ/OKNPWDbZqHhQptxUxywp0Ku+0kMBsHSEh+ZTg
rfXnrkdYMWv1nG1lY/OiuGC7+DNpllaI7YaDD9vHePT/bZzNl1ktudbQOHy3hDmLfqsVfkjwFUIc
L/JDA5sZyQI6dPSeAEyh2pCQ8l5atj+lSitnVbtctOWPnWzc0SpIN8Vt0LNf3W83KEV48lMKR3lk
mLykTT5fPsJGqwQT4LmVO+NA8UamTM8iFFdhbLp4ot95JEzwAUOIFgRwALjYTN35Tyd6Ln4giQP+
oRVcjxxS33ifey2Ab+6fqLy9bM4TNg0XLF0+jisaNbX4yYF4466IHQTyrxS43/2/ZoJ2U87OwofS
L0HhQKXl94ZftULj4fCUbuiPzIJHNs4wYihVzjYz9eutqBiawjcUs8GmMMYX8nlPvNqpH08p1xdY
w7rJJtpbhG+zRSWiYYfrWmB157iwuCmi0NlRcg3ktmyxMasOGPd+h6yP+htAKZ415mWU2JS/wIzs
zUJ+P4W6ICq4NTTtN6s7sijEQTdwIOdbumfVRDtLt701htIutER37lMG5eTsWZgFbsH4lhJLfMA7
wUSgkkW5rsab5+KnT0MYJT/3Ve/AWZIZlCZu0RzWHNX8+jjpdRz6zYHraHYpYGD+LHbGRG/GBiLk
g+my44375sbFOdYg/WIu4txp3TY+p/1R/G8/xtRxqueQDdS87jGI/hDnFTrZ+2ONXKgT6zFddSBM
xhIsLfskNWbCfS6uvcTiVzXcHmGRI83J31NTpEuPEVbFCuqCKhlbrNBkXBLtXNtaH5MQF4pt2X0O
/ozuX6DEB0+KGMkF/005WJvGma9Cjewx+3e7pjNNB+tW3AFuU4q1Uyz/Msc5phG5cCFSJjlxgreM
YLwWu2ZdW4zFZCQd7rxTTH7eAekE3P+oEtjyK71joTUYv8US3lF3oRRyMukIbPcxG4sIgjsyIv0o
Owz4woKrtviK4Ow2RxNRSheYcyHOFSLYJmJAkXbjdVp7b3QCKsn8/A6WQiYOOjzHJyQEEr6pQkce
AEN7YyxqqqCiUODUNEwDv/0jfu5LjCv64oOq2o7j10Dj5+lYH6LlLxtgUvTtBBJtYAeWnrb/eWAx
HKu/dvgpNPSO37Rxz6dnMERgkN1Ofw0VQmunz2hnz7tNfa8NvFA0vTjxnoaAdjG15YBpsP29jJ17
Yk9cBB7F3oR0cEc5SJRY3+C9JSRLM0feaLG1U1hGZ613oWmYtFiVTuWFYWq9+o0tZAxKV5wYQ0kZ
VjynXQQMrh+qks0rz+JxwFvF1DqtpXZylAhhyMr8TzvrYXQTdVYm0KQDa6E1HxVnFxSNiXPZ3tEC
rhEl6pLUndcxtfsLUuvdE99zfmW4BTWeEinUDO/7Ez758dx4CQ2eg0rNJNTgCLWGT1bzpaf/D2LB
ao1LSWSdLapFBf3ToI/fTr6hgC0oY1CMeUJWc65KQwel9GaYyvo8w6eWNgWI9aHdJGGteZV4v2Oe
K5oxlkplGdUKIpxeSD8eb6Gal69Fjghhm60dMfM7y5HBL58y5C1Ojf4CUtjpvGZ6N8U9n+F/AEpC
X8ng45cUw/Qjnqndzs+OPsyvo0Ihq2+hgR78I/Ms1f2A8zV7aFFX7HgIdLlZSZwf+ThJXACdH1vf
Q5oSKWJ098fcM32diEj+2c19z9yn112RcBmUbEI6Ze73D/m34rcgYgCH+rW7aCw8DPNoWhxrTg9s
iKhVgELYagXeLVmLwWoTy1QowKiX6gAD9mEj5j41sQIVFdBr3kWvQChSmskYutETLhk5zEfNPhWU
40cGMEb66j0khTx/ed8uy7dSPo4EvFYosoKV+1yC0r1RkZOTVgr9MUPXLyEamcgocvJSsCcXjR8U
LZzgjPXbhlRxvSIfTjhmsX19kDQG+QrwAV5lQ62V8NhOXxw9qlds9/qMWJRbv1WNEw069Lxc+4xi
FA5xSaIvGsn2Tw56zS5ant7XZ7tNNuab7c/v68ipfcSlTLn+IifEo/9YDp/3ZIArnyICsXdgmSeO
KubyfomzGePdFvdEKKLg1nAgmVJBmlLhZbCXXLp2nlblscnx9Wngn8z6er5m2SeJB6aGUtYWI56G
844eBmNXTNOkeBiKEp82VewdsaxQKgI5I7IdJhwuEaRF/paUdtD8geyYT2y3CFAlGTN+ZF1O1sb3
KGj9Udl06ZAzCW6TmznuAEr2PvmkkvX8VIR8iAIexUca70wIdaEwczhgy75UBXmQ7pnJuAmMT7lQ
7ROUpKrzbQYTpPKmaBB29Kd2kwtbX8PSqnKsxa/EYNshaYLd+cRdjjdHKwPZqI7JOkQ0g0UKZizt
oFK6b3bKq7QJ9WGb+psvfo4Y8S0eM2GhmaIMK6qMYQYCmLEZ912XCvRX1XiWjrHvgqCCz+VDVapf
ZtrySNCG68ulazfJ/g5c4ksaRyQIy8sazVce2J9/2DahBdRsHfwzgXlwLMCGYENIRDhl8pTQ3z54
vRZGJYwlfBMyA0neIIgCXheYG0aLJm2I5VzPIUO4SYJTN0AXPqR1G7nAoUnkR0CZvXNlRs08Fheq
9AsZSauVDkXEXLyjUEHwdtRP+jCLpjbDHiPFXdN6TLY18oapzmvn7mbFvaJ8OhyGXeAY4BFY6kW1
dHJq4/SrOYGvVaZtxDCIInaagc61umpD3/JqyBzJ02adQZiHpOr4pKbWZvUqLq7ulYWyBcZYgYNC
PiPldbLOQqiho86hz8OIiEpib27IwHq2ejpQnOFcuzYp1ty+zZ6hjLFNqqMN8wyF4pVQb21k4wOm
x/Ila0mE5mmd8kaVY4A0VtguF8+uFgNA7jz8UNc+dKEuQQL9Zr+I8hyPq0KrcdXmSz3+OVUaQaEf
7qnb5Gd7U72RWdLRFcltlsx7AFIOfJ07WRaDPoBYpRggYNpzpYdMowws+Xx/6PDISvA5iBE8s/Rr
MbPTHZajqkm9fe9ZnTfb2cPs1VPLs85w96z++vGgyEu8VzzRawh9a2hAr164zrcNQnoWnuCK7yOo
Omr05hBhwq2xPWGID+YhG7lLPmY1ZBEVKQn/pQLnzY8eQe3bgll8EkF5Vw3hrAs2et1lVlEgc5aa
/rml1Cy7SQ96eYs/S//dvfXQe/bYQVmIaVU6DYumfJ4wb9vbg1ERprXi+NgjFjK4lckPhZn3Wta8
5QY7NTfagm7d+1RIauHJFhLP/zgLGhSjmfpkjmd3PM2h+wMYCENpmTqnz1EIKmvVBUKVYtS1car1
XQzQhXrgze3bq5chY6poPQwUJj99waM7d3yui1Gkgl7U1QCfSQgJ5SJ5BtLhmdUqetsMs/z9y4ww
IKh6QSQrM/P8jv3HYzo4Gh3CgI1mg83IZOrYTFwmc4LYx4ewdMTznHI3gEC7QYRQtunaK8+KM4Zx
pFuLIVMm9u6J6VDyTmrxRG3gpdARqV2fsq1K9b5rM4AFWGeXpwMYbjb2qE3cu9Rp0TYR1QTpxmJS
NZ8+jw8itzp7YWYlPZYqpzzig7cAdz8WTrLH5IQhF+g6NyZ6dV0gedva+e0cLHb6SZw1qlPV3CQQ
aun6oAo7ZdPofQ3b9xwALYXbT10SqJWIwIhn4cMsZk3Zm7kYiZQosERY+NweEdPSkmsx3x3BF6h5
WnAbXwOyCVlhMPHQuGgTHWUGQmIqO6k6hIo/0SLnuZ1T5HbgufueoBpvsEZzsG9ujQ0QVMJ0VJX1
2gCrWdXzUpzLuEHGKTScuWLcu3pg07LLU0SnU0JQZymbYALV7wamp935uXPyZvDZMSF9izcljCN7
8Oq9U1LDhTtnvKqvr4qZ3BizWMkj5C+j17snnFQ6bi5cZsQmaEDVd5/96YomQSqtTHs6zvfyu3WJ
t9zWxtYWl3fwaEV/7Fg/Y6Dgi7mH/0Cza6bVEgWVsNKv5Q2xO94KKrpBwNTHjCageUo9ubdjd7a6
GYViwy3D9ZpuT9jz+jq4AXRyQcvQv00yGr8yXZmdDpHEKKa3HgepTjdfOdsiG1wY7qAfxxTL2tWa
GvUVkjSF5pFyuKlXWT0bbtNlyewxo9daVPxgx3MQNv46+ORN57fZknAOZOPhSxEQMv6IFdZkT/tZ
4bNYQ4XGByq/oRrzheQTFPrzWW1aoHE7DPGQUS88LJqps7vAJc37yP29LgyEkm/615C/pNEGkXqW
vrFrNMZW7CxAUW7lh2Dpd97eJkBpzYPlLBo6P6UVbFmNAabzug6IypEfuzUN4mymXZIsVlkaLlol
0u4SCAQs4CnQiFRsyaxvx+kKbOckOiuVId3sKF1hIMTgHvXr6xIHzMgigpMs8kgi7xar5VW7KM83
iWTkFW4Ua7gs/rP/XyqegXNC5BQLhxqKjMD8RPUb0FJhwKPejcQPnHVd3+ZGSt6cJK6oXWABnS1E
RXgQjYPZV/MFOIwRnjLXTxJhDGu3Lr8L54HKSoimCGRbZYv7o8tfsZXXwJUHAvXwKrynHcLRi/ef
pQuy5QnwZ5siC3IQQfBOSNexaB2N6tcWKEnDcvhY9RQB13ljk1SooJcluUVxUZ9B7xmTFkHSZkQ7
4SIfaPRgpiGESi9OWiL15K1y6pk/Z1FneKJ6q9e4EhFx3AJWic84dAZ/zg9Uk/riqN9AA3wYzq//
0cw/aReAdl4VsG+POJ6usJPcqWQP5XssSjjJ9U59weFwOIjHXJNCvnJ1zKxec+gekzq9qFYS3+MW
8tm4yWbC/uHrbGRejo7j8bmqAdfh0pyVXtbDbkE8FD7DBtZuMm1pNQIv82R8/wZZtAm51wgfOCsT
NmBiBNfY4YrzD4N8DIg7ynzCIt8sxzWFrRPxznppEHUMz5eG1LUCA5tbHteug/LYRJbX5xqNq63K
pGIYSTe27+Jkh7IPMQ1HcRgU7MG4Kl2YW7MXIFLWJODQsuOLUG4Fs7SqaWWC4yP19Ba43YWhdUsq
wk2262hc/GF5Ckoo9F9pP2h3rRnnzgyOxHgjzC2i2BwibpMeiMLF3jiEIeMWVDT2OHBVk93s6GjV
8E1gKsCOExj39SIRX3wYNnErqBvDSRlH67ywaI6m4gaG+AMtyPHDu7WUNEBE/uTeNzJpHyHfm/Ur
kirYT0t8jW19OCDnTIeY3N35+91JTAdYeNMgOIWPR7X5R3co43+nXaSB6khhuaWs8k+d+yLYGp7N
36BiIDslm3Xq5X0Nis20dDyNVJfMveTVyreP1F7XZwDR0zZGJl0U/lfBLQb6+HEJY+K6YwTb+4R6
WKp0bDT4nkw4ev3dIX7Ea3MYLQFCHFGL7H51RaMYWGtw9iswEbDfG8340hIP3gvK5Mw2knhHqaKT
x13zY3vBH15o71EWtJSKXljSus7DkroPl7fSbSlFgN1WFs1uTJwxojCXlJfFWU/pEt/1/8EXJBjb
LfbX73HeqgiocPuYCfqKhonyKc1zq9H2nfn/Xl+r9aItZxflmjwqGN3skILgQ5ScD6eiLPb4+Ole
YJ6JMrhqe39dD7t7g2bzS/LRxvPvxZEeheBtBzwlpxAgccHofyu50BnMputyGx+uXwNlxD9UU/AX
HCbv3YfVfVclH39Jh4U54MbZD8w55gYCIC7VVenQ8I9+L98JbNMqe+84Z6UBq1QtHLGNMlD4rdzR
Qt8/KWhQvYTwVoAMJtdXDU638dJrm3XmppKstkO1zzBxo+uwgODz9vp3OJ8bkIoPb2MxyBf8vgUy
eh4XU53pEOyYZLy+mu+P9hTJAHlu+SjX+jXGzPx1b48yjg8VWMcza0kPQ/ElOnaKxOClvYWDnyNT
LajPVhNaJ5lQtkJZdBAB5OaEzaBaZ61OB9h0p6CxtkiQ1lEupxf5kcg5gBtxIQ0NOCZ2gxvUXNKJ
Y/h69FzPR7sDD//15qn/+XO/2VI8rMJpr2AD2K51sggm8Giax0QXCbDO4chMRyV3OAYwN4RLBkd6
OEmHVaEvL1Kuz0IkpNhZu+X/pRRZd5B+GjeDDqIhNXvXSJ2MZTK2eG+b27LMhQyIMyx3EHJO+17n
JuilmANnX28T9krHjr96NXpJhyf/yrHUic4/JYyj4j/YIzAGk+WJr8ElpogOy9zZA6YMqu00+KSO
kYyJY/Jp3xr7SBre1xoFdKZ3Fy5R7gG6ap60PfHJMt4u/4i5Kd5jHFsXrQOKpOHJky3QIR8m98uo
HQtD5gw44WmDIUlyKx7QHExbHozriBViUBvuWx08Cc2a+BKsEkRKyG2WOeW1L+xZXALKMMal5Kq2
OX5ttOHh7/wtpBeD4JdSIOayeJ9lsFoGscZT+tj7s8Okb3q9qIwkVvUNw8RVqB1R0VSnLtE09gss
laX4UVlHk75gPIjLw9BUWYe8rsbzVaOgdWUR3GiBzDBdl5yglidZFNa3BduKU0uGs7WJ+LNGzP+E
aTX9QAXKkwAqB0c54RQYASvXLMCIlnuRVaG7ejyK6iItcR8EYWbaIDj9JCf/59U5HQs6/08sQK67
VBxPFGvDzzaiWGZtGPirpeqAwPB3MCGaS1lNrbJf1GAjRCAjmSL0VWSDLDDUyQjZP1j33djuq6tE
Inw/Jbii8yWoY2+xGi2l+N4lzxxm4CkO+ZagTGJ2sZLbDbYseYiWx16zq9tamDySAdjIqYaHkLh5
ceWzNxuVmLvX5+uvrt7WhPAfG0Vj7xvu0oNq/TTgsd7BTwipx6M2UwuwI4uNZMNgOrnUXC07JgAE
u2uc75oBQjO5ztv0bbZzJ/NDlrRGPtj0VTX0RsrSHAq/MzbTshOT35B0nDCFihXSHZdcaJGAoQz0
V0RaA0WCzOhNOREsFQcRjm/daogs8cVnqBc1zPa0ozpbSWqeTXG7HNjcAGWQYAhnsaHxTSFhBU0F
frpk+24leGHu3Vh8T/gsVJ6NhUkIOV42Ym/perupRej27p5mYkWOAZQkWex8Vxqe9XsXt9HssdBN
2nCQjHsHbyx+2ZNE2CR8ti6r+1/LE+hzxlKv+InZpei+5Chlr/ECN+qLdy0ft0E66NgFxX2yHZBV
Zyo63mE+r6uxh0tLdV6pt5TjcOIQqvTMFIvN4zJWDsGjgtzjj9zRQq0hISX/w9Z23xpq265qD2ub
shO6rk0qYywIsk3bVJX0Q1Jgx/E8KP4me0wF8eTmaOSFyadGDjK3HXDCwvJ1ydgQ+NxyOs6JH3kz
5wcYEpxsWzoPgJNe/IonloZlaiaglRqEH00CkKsXV8O9F3YGBxwC8dqyTXs5LhuyTGCfUzV8Gbf0
H2jG042CGo3PBIE+q4zw8n2siilbltGOesBAm5bHP5SHtrlNFiR4U6+jdDNeuNtkTLBUkGeJORai
4hepbjuGBuCr1aaVSivTtA/jIcuGCvCFYGDJTREezhwXtGRrYjkWRzCsBe60Cr/e6du9kEMGlQUw
lVzHOrCtlPnn20UgNGqSoQDl/0+DSvuAjh532x2yAQ5G+tPXwmg1hTKxP2thbcHU9AIIXDTFbzf8
GillkFBfDbewvHC4oARDewa5zzVe5KPQqDfVtBz+hn3hx+k4lrw8E30Oiu+z3PZp6bf26wClnjg6
U/QZBYk3wwDd3NHR1jJxN8AWvQlQUookf/rPYf7jK4NrqyJ+ceBfVF9jdudhHG5KN4p6Tqdj9i7O
bxYC/07TyoeXZluTbdZDdI779mWRWg9Nk/ljqdEDD9lgXiRZRFpVey2Z7bveWz6rJkJ1OvY0WQQU
6GLy2ErjSpiEx2JR7NpkYnkFcF6Wm6z11M7yGeJjBqey+D1cc6gF4M5og+21csh5A0VwH/lBLnj1
5DcbdpzNb9t+c0WcYpMdZZuujVkCDKBV+9O9bpt12qTnSUNDnZJ+dTRKc8byY+u9XSeUNRWoXyRf
lJNMhL5fbOZJ8oq4cmbWUN9sd62cQzJC0/SgQbIQeLBRLHlu6XFKDadfldHJtCewhH5Xy3ubicKF
q0Pn2XH8CMN8V1tfp7mqlVhWH+oR4N898d16owW/je/991bIMoJz9oZ/pHyjTR0+N8d5ULVQjPGr
k4eQSzd/rPaLR72cCN2eY8uTLhYNBU0Elmm2XNu4bqLqxXHnj5XvqgPXrwGk/8QUnwdRtkE34XgO
wSAh+Xb1Z5Gujlk3N6eH5rfUAc9OYZI8lydqt3l/ldb485aDq072yMEjnF9dcuc4c0l8w9MLJG6y
2XYOw1mvtCHIHF59kdDAX8+Yty4VnuhJiNvrPWtNVlKHhyq+8Csw0bjT3oOl7cuZ82yatz5I6YD6
k2FGsUtJO8HImyO2ce8DgI9Hu2BCG5WaYRe8ChQrpJMAggCZoFUEE9YJwHOQJ1F21w1xDq7bFl/o
SVHB/KqIgafITEErgQn6fKwKAS/d5c+/8FskgME1YhLpFVWqD2cNVa+jaXOUq0Oh/2LnFvFamCA8
xpMBRgGgDwjiz9yQMcRtCDOL0obowEXP6Gb37hnRfeCT38aVzXZUFQH6cXHBK10F0MZUX4nQfnYJ
p4Aveqf18jn/C1ItNp17mSkCDu3vOnxo16W1UzMDHV+dZrGcxtbvT1QcCTfbNm44eDAKt8cZc1Ci
aAjbLs9TNhVioDSciuwzmR+teVe7CKhh7HgDQpjXpot0WwUAw4TeQlJyXrU8IUyP7/nC+ptIfS+5
jI0d+TUQ3YElgjL8a3amGrehBFNri8gyDSeh/4Z3qJpAjZL31JQOE599GEb8jwFK1nkc8sjJzCS9
13/FDSe47R63fXglW6rLBq4vLvQtkJbVjC2YB2wfqyxZ1hVlI8IlSP59g6criW5o1GKQZntJRWtN
p/uk6s4cxlOrYPmdKfKN/K0jpqpFr4TPwRtra1E+F1wii/EwI8rJQkTTDZOWDR5NIat+F0RBtY5D
VAoNeiq0Si4NX2Mhd1Exj95FmutST4AGX86ZhMSBRAf0dQcsp8H/U69Swok892hsbMWjZ3rxnKoL
phoDGiCZMvQklHWnqNJPGlkIr3LhMn7eFabAEPok10U5TFnzZesRewgk0ifwTGsTHjzlddfNyACT
eojsAHkZPepeW1qY0m2Bgf0zWfG8V/vSS8TfHdauGvXxwa3Ym5dgj7a+noa1lcl/RbCC1SzN3c4R
Pjdfk7Jl6xMEsgNE0qELtAeHUkzk89G/dN8mMnYLAoDN5BiETH+uSuZqUPc1g4o9yV2TQ4Plv+xI
cEY+PEgVmDW+FMxNsf3BRLj3LrpSOgC11dbaie3oOQodJk51BhgKxYnCAMU6cSQn8gvIvTGXBN2i
eaNJbqloBU2FaPV3V/qvZ8+ibk174jacu/dG+n1M7JSP56VbApvn/CekJs4y/aJfAuf+HYtcffdt
WbhohI802H5OSqMF2ge2b8/j2F7RYCa9vGqdgLpb6DVvtnPVC+nDdDphMYvAnnqjHo6OHA5eArKb
Tg24DzwuaWdLah4jRguFeJRbWWL9Twdm9cDYgWGM5bpKj1bt7z5HQ/Sy9ua9O2C/QosyIriPT89b
dh79gXWZbLo9d8/biG8zk7gBJtJeFkmg2E2k8H+VGCeISXVOYcPrpjthqeO59IoAWajYkDAAGKxd
GGb/3q84/cX1txDOarSioi3RJqRcbrYMUEc8DykGw9m/NXv7KChADdJiEATX9GOHqJF/2lEjQj0N
aqXVcuAdyx4Yks8T8pXnHlh2O75Jg5EwtPsmnNDt7Jroo/Z+L3zBdVaqhiF2bxsmjzy9J+zQnNyd
Wfdxr03KRJzkcWDTSUjAEYPzPpIWvamQhbUNRyGfVgis4AaRxl7vSvcha640DK4RVya8Z3hPQ+tQ
d8uXZmuwmsFeptKRkI0AqJ0XcI6c+rf+HPKEfy02iavRBlyiwv4S/GDykccfgNdeLXDHw3M8fhoq
KIhiDdyNg3AAknZT+vc4c3sVfJi5NrdWAV2NjCTM21cKKg9Mwt2DPwrjePHzPrPXJ7cPh81jJ99Z
AYI3kuogDItsONIpUicSiJL2NatWBVC2DSDrIakfnYB63pbjXxfASj+tmxp0BHeMzF6LCZe4ZCFh
bGrimbnRBbJRyS/BByarB7HoArsQwmsJJcLmDV24lsPauMP9+6fkm+VSif4ph4xk6HO8IVM7fpgN
BRlDY6tbEjAmgkccA0nEB8ND68GhYrNz8ckU2NvfAhNsa1m3r1lcqYhpu7jyrpFSUdIL1JvcFlkb
wGHKWgpAHY/WNP5HFfW1ENrR75XjqlB3m6+PgLk+lSxPJoWg8syAvu7YxAHaFgM4THfBT5u8EqPz
IvlDZLNlznu/83vGDtMyVCONSBGwY1PafAWiS/g1Npd2/s+OCmdGtei5UBqZdjyZiItztxNAfcej
py+J8Ge2ji0JFCQEKkzIH4vDFznWbRzUfF5DL4YHBKZ/hG/AryvxCRYYGgt5kdnp7U0vIlV3Ac2y
6rFHYVcsQ3CN6OvR/lKfouhLh4woZAQJJPgDONAKtog3OO1hXD94icgYUp3WVeZOm6/ucWL83fod
yjHDITcMTkgPbUKocGkn1FIQvnVpTZmjBQAOq+kUdcuDQPBgWiYuR1WQOfJlVTweqRqdd3l2Wdci
ohZqITNUwR1bCPeiSdDmJmOZKEYfQ7YzGnckgFZqzC84KNT7/S59s+cagg29YUfE67E9OE5l5Wth
YKqDeWO9YMm20+hNvytvnzYVblOiscQwRxos9KSt36iALPudd+lD5/vDG5kbqH57/DqjxQuiZbS+
m1IM3Eth7LTcWFbY33Xxoe0FIhdQDzO4o1V0m6umIxYjIb+ACaGfvl4QWtODArtuefp08aBa7ZxX
0QElYuPHd89Vxwp954l5gWqcQCQYcERAFJh96zoifW4dPlAyMLh/49UAqFOjWtjtZbUGLjWR9vVp
A9UZqhDR21Kk2c2Aerkq1jhha7KQaJl5WuYnkIr/tX9wFtzifPKy3j6cXHwJkPcbuxDaFr8fLBK0
s5Z5dProaVIkcI9tWL8G2DAkIhwF7tDrCpI1YjcbCqO8+h95effbxrrJqQOiXR2DDP1SwRIljOPs
hq3lCcjiYLb1FlSsoBHl8hMSczO0oD+6xlWfA8RJLxVBO5aax6FXupUL5TcCZrbhdK6mDFbpc7LO
W0BhVpNw2Xewc6kqzvzEBa7H+Qlr7OqXc6L4eDUCjqZrG9JSq9+eMgFUpsMPa2HTjartMYKzpMFW
NQYSQpLfi6AHR47SKN4a5VHB0GfpIpDR1UApgRjH5MsRGQbJcQ9jjJqxJD+pfvi65HcnKysKgb63
Ov5lPsn4FApTn4Jqf7aQxeyZiD9naaHKy/zjeWQsG3aSi9lRyuw/STHtwobnnSj6up4RCXp8QmYy
tzt31WmO4UITdKMUQ5DDY1/pPFT+sRkE+tvAlVtIP3VCu5N3AEDkM7mgj5mhBpmok6frgFoz1axl
Pd6RuSm/0dPrXsXbstxFltAQs0JENAhm9EbGmHJpEq170dkxDlygUhEMOI1NPvxEwOS6xCoWnJIL
x3G1T5CX82hW3Wj0i/y0nZdPJWDgrHxSLYRzTUJQITxYkFaFG40C0/eKiGyXVBk0dpCW6MMoyY7p
1rS32t9HbxfLOie/zi46W+aVzhbxNaJaMkDJWzi4GKx8s8HXRshegxw73A/9J7VEpTBgf1hALgL8
1Y1FSHrjgHKLaeoBN1aoIjBGNsec6tgJNGAs1UtYMBFmtp1SL3NKkh4BA2XJiCpbJa3963Bhl69E
lwcNvgXt97jSjJ4auCZ/dfvPawFWNmNI+o1a/3RWKI7Eeg2/ijQIvlqCuAhDjE7FoGRTJj82NAcP
d4AKTgk/GDYUiHkgNEC3kug7S6QRihIObH2MRtLORAPEPx6yylVeYY8VzuMZkUjE+Vw+4otU9pjN
/c/0cke5Nz8vzZi3XSse4j4gfSndzcGoa+VZbEL83qoiTErAy1HwNaSVI6b5jUqvEddNiXrdoKj0
kv354Sf/SGmzx+pVw/d5BSrwI4NzppENb3hRLGEGuqB2fnDm0XvAAoqkv47NtZnUXJhvE4rdjfTK
Zfl6xWIZ4datWSugnQzyU+RPZy3ktyczYxqs/noYDsBEY7ywnBJyhKbiBjeSKQiUPAeVi9tDHua9
5XzjrHSBh92OSdRnh1Ip073VbBBzralHtDkvwJVLy1Z1EY3iqFwinng0o7at58XPUXSJkQeYzxKX
0m5Gsi9g7RPuqHBJpEBdnl449cBZyEG6jOE9mNc0/T7HcPTpqMxbDzP/yRarS/0xbKS5KguRfvM7
J05AIMo2a/wBUgMp+t77BRsdO+39G6DFRZZ57xdjqAcnMuzZc55ngwDwVUZphb1Nrh5wSjMV8Xwh
5u+dJjSoqTL+hQByO6io7q5mSt53ty3l/BFsPnjJ/Df83E5+DqI7CoWQK3B30C5gcJUyEpEzM5er
CGLxGrpwD7CLdFVo5a3LZypnbCflejoaFa1BRA2PMpQbepqhCLpxhi9p4ZmNNOYA2WNnKQHKndI0
uZTobyaXX9RNnxi8oQvjHNWKAmdFz6o7FiCvD2+aCqQ8JELWeyTnw2yND1Iokt+g1ZRQ1bXoQF1m
mTZ62Y1cyDfCFNrbxM22jfLlhRAmQCcadQu+dMJIZucKXksFT5U3RbrQgJxdnRLqObFhzuV8zbDX
542h2PgxnJEE4PFFP3IYI1kWdAi9Gu+f1kuJI0PAuwPBnttPciKIuBgaACVJ9o8cqRvCq6ikur3d
d9t13/4/2z1HB+ZkxJtXMjXToIWXVi4Q87QCO122OpI4TuwS/S5w9Tx5q6d/wMNX/oyZAUtVd6O8
zQGY6Rmb/3iQ9NBCNEWxsB3c2X/tdNaYMz+9U/pyqUJxvi3X1ATDMbY3Nfut1ljHZDUMrZxuUuQT
+Q3dQJGOV5hm0GRS3n6ZzCWzm9ziXSffZ/ryOHW98AuCK3tkD33ZlPP6xIjPzmWVQPrnQ8ZDVIcb
zXcIr95MYts2aXdRN/EJyaMCdeI1cz6WqUT42ZjRQ/cAV4G/wvegcYcI7myhnVXgpXgT0JD1wp5g
VFQan/cj76EclE5xTYqRwinQL0viaJkNEvo5vFa9o9ZuaLcXzXKB7lSgwFT7iwnMveXTld3IwXgp
hKPl84FCX9SmoHWdRuAigj4gXkNkJZQ4FUEt0oh9yjtM64y7y6RiMhJEBFZ3xrbcaQbLAvwWx5en
Z9VjfKBFddRqDjAAV7tzA+0YoYUzl1iXKPDPR0ZA0ofdNXLIJwZlyZYZWzHhv4OUuHKBSPMb21G/
s2z5V6TjP5vVoQB9zk4IKpNjWDGpGCzSsIap5tsVaLgACK+7P0CJO9hyvMzfMXseUf3gbxvwpa9/
EHen4RIRcWhI8LOAh28mkSXyla4TT1/mo4zSty1qozvDcGY4Ma+eJBmLMW3bUTRDHZ+Vxe1sZwjU
4u9TIRcLZVI0VMeXY/eolwYNcNSCIT8BE4E1Acu8vlM9WaQyN4UiHIsc3XIUElHMWRjADguKp9lz
i3KT4gqi6SexNNnj0S46QIr1hcGpQuAyXLjcYvUHvPOG3zLP5hug9CkkDHlrURFb1SJJIKKfw5nP
8IDuW9Stvow9fw08Szr2DmOszGq204bp+/ZeQkOOfnN6KG6eotYZjLiGekPiVCbVwCjV/ir0ou8i
yveENQ8QAxanenltO64LfWeDxoq2AsgONcrIErbSOqpUWsYf2ApzP3f1LBfcEJfbcV+kB/FTEj4K
2cfuA0VvJq6dI8zO9hBX0JWVkMitPTbmKhE5Zqo+Uykv9WL17/sswih0Mq+sFQgwqcYciCV/9lga
gj3S7cvaY2Mjm+3D9yd86/g5Tu8/ja14RS697eeEo972f1uyvdT64EWaYtz5Ee3CS/uALB5ZFywQ
eM1zSWusptcyZpiaud+LCgeJ24+QcLyADZyJCZKxQrpqe46S5AL4YypHtIf5SsrbAw6lJ+ll0nIe
FhLUe0cr5zA45/QGkZgY6sn+8QhrXoTiTRiC1F++zr3mll2B3pPjA6NwbcY48drq4g9qy/JWHF9a
cmOLxQq1YL6ICeWfdsVeEQLB4bAhhuGNqXrqI+NimdVQO9HF7QpdE6l4dzLBUpPTv1Z9y8hRWQ2C
PYP3UFIVYJRSh08OCd8kEhA6ZcFNmLSzJkHdxQ0hV0F+Zjyu4OJt7dwE68MQsmwPYtEsAUGmUGMe
AcjSseWzoUrivRd7dmyw86K00jiZxuDGZlJFM9AWKYuGK+YO4U5tXa7ckwPasx89Yfvs/z0dQ+c/
0QNObl0tEyHfsQCOmPYb8dxPMhufrb/C4yAHqzaDcVyOt/48N6gQCirZ01Z2WnvqzZM6eanUGv2Q
xOPeVBRSDtYlFaJ+dt5fGtHJjiqgeYmar7OlhfejO+KYYmf5aIRT2l/rQuWQrvMmJd05j2ZYcTJm
qjSXc9LKR55FRDJ8FDiz2/cdcHbmYDU3ySqmZYyjI5eJWbhhZMeng9cVOzCSjJ3rPNbG2QOk8c7E
EK6IuBxx6UWY79KiKmTkYbBW6iZCV9KnbhrpnH7n5xPBGfbB4A6YALphXD1Mq6BrKjvJ91W3+kHY
RLDP/v+14VjwbmYQpNYpItEeZXeEnvdxw0zaPY+N282gBP5qnaOkEIxKlGaqHZrZeKXmNZsKZS06
MfbKCGuD9SoBP5RBVAryA9Txaq274yO2Nzy4pe9SEPBvBAgXvJIZjRWMuBcyYMd8BmBzCzRxf/YM
8Yotcz9p2PGW1E37AdHyBudF6ZHeaDDyW7XC3KKkJma/ybH8NTWo1IGBXcA6yFYC4zm4H62uWGvp
1UJXjiiM3FrMbuSUCOfASGweZlDK+sElgyUsjw9PALv9Hm1B68y3iCd7iE2LIgUHMvqQjtXJVGgz
iKpi7T6ywxcdUMFcsaCd9BHJfWMJ7XC0CDjvfxDt8jrDRGSQfzH46sO/mWf+hTl8h56c6bD3ilYV
Shs+BxHMpqPHxdZwI22aivicuSmJ8y63amv6nNlsQ9oQx5IZRBpuio3q6d9j3EtkRMddm03f+1WJ
lubLV4B9s9fyrNDtKFx9E7meWxPzFRUlXKuVvRNt9dLPA0Jvjw9WoXMlxbn1btMxlxxi+Wj8V5Nt
6qurasZcOHzHRgUa05Rw8D4pF7x2HrZwwiFfcOM/ATHmNsCRbgjmcyG/aMwXdNcDDMs8wmj+fohd
P+JdNZdIrBJWdZPqnYuB6Z9YhtF3dGPlOOA1v7ay7NxZL8TAFVw6wcojpt35FCeD8FALdyHdVEYV
wQhJ0y/0WJrUjNJBxNN7zRHpIojprqcpdJ0BLB771i410hmr2Wop+aP4GXn2pAe1VV7y4TBjnxke
NrK50CpdYRqJeZWLN2Aqcze0i/WHB5eQ8eHoxXkzkXbzeZrfElk1VIqxPzDtGea6pfkmj33F6uzV
C6P+EKgyTTDxBh35ookmqhYOC3OzwWhUyKN5iomifcnYQNn6nPhZQ/BhRQzAVjeh8pRh3Fr/SJ1M
Z+4vtGQR5kehQrOEykYyMFEpW8qvZ6lLK4ChOuxRfhEoKU7oP3UEZlUvAaZEGWOCT3w8JGOA4CjJ
W+76cTEGRBzwe1f6P3LjNhPR9/82UPyPXvQHd991AVoRklXznILbfORXHnD5EzA3bD1mLn7Ny/1v
IFBHsUW1aOVaFASoU6ET8yfaCNAsKSL+ccevY1u9fk3Pl3kTv9ZlnmRS32xXG97QvsmdtfukxinW
ykKaZCXVTIeLltBHC4rqV21Fj+5Hzd2x2udSM18R1W2goo3MwxXYpoj6kkJI3WbAukrspnC2UAvs
kXn9LcR5wxLLeKPkHIx/jO1qT9DpxS61B+ikSXhVgMDawEAZK5HaFrleXfz485dxs8ByiWWkxzWa
+vlFp31TK0UYxXVZlCnt63FYllOf0lqxl8v3pzz69+UuTFmirtUxcRzbtjSBxUTAeLEcYACzYxSm
++KXsGk1ALdnm4J/I4yeuJFymAwkFt872yLrGnr28aTHR32Uen5KIGkpfFIWHPElVk9SthDw6JkR
Ccc2lTTKMX859zPwozwfiS7Eyf8nxGye5VvQA1JEoybloCxIaNjI4uvbd/TaB6f6e4KLW7E2J6HK
1aYi1ua/5oUmU/Z0bio/3DuLM67uYk5zYrXWcb8TVsrgpr1kUEClD/BBsUO2QS5DPxmYxZu0Dfy7
D2fj0aLRBuoUJ3h84qUxkqD1SxAK++yre6r38EVDfHMAR4RlqWiGMxkB1Jll4bJDusebp0WDdAyG
KgomZIjSys9lLMPEdvckaPzv5B3g5X4iz2FYY/OxgBbu6cF6kUn+8YwF4MO29/9r1Yse+QgXUSca
Q6dpPZYhwdQ5DPJYeaEBqOaLyNYjcUevVWBSKJF5b/IiWTo7dxGSPdDg53GQuFnoGAiRHzVNqGVk
qAZ/0Td1TOK4Eh/Io7xZwHsRrMAJ4W9w8woWG2oOHzF3vs9g3au74UX18pVJ/ai+E2dcglITERfp
RiUTFYTS5e+2ZkLppFuafir2FFH+sxMtmj/4Ee3ks6wIT8MuGovhDppZI0o/Kx5D8e6rGDDY/4Ml
N/jkM31d/fF6/aPXLgr7PHAhoe625+DY4kebzAH4C5EWsyvP2aDm3zDUOohnd/7XNdtxsjeyH0i+
ZdCcr9ceMbvOkJ4Del50j6y9pyUmQRZHSz6/iVdglgXzcYvP/j/3L1mDJ7+a8z+LgcqvTd6Qst2O
uQs8zDNIs0OlFwMby9pC69KQ9UZFqJInyUPrw8DuDc7DfzMqLUfVuE9hk10eFItLpY6h7vKbAkb8
FkGRx02kPNNQd7FZfp49fIcu3bMgUj9psiQyDZhmeOcfM0cU/RfB4ByQA09fcRp/6EFMd7xa55Rx
lQQ2JvqeNDB3Pkd3TXUoJv8qdt2ok+O3fJHR01Q5K74PyZBfTvQd+wu/uasiUziA1hBrzbHWJ2Rs
D7JkNrMn6oQ0BWb2PBX68Zb6jjya2w+WWoVGNoKe6hxkqSZOGKQa4QEFU2FwHcT1mtXNd1qVM5dO
9uOpS68lt4n7rtv+RqUzAIIjYKh/e/HWSiBlJNTHA0Iio7KzCW4wKOT/Yci41Ulc0ysC9QJC4FLN
fwshWrTUFi9hKzqzzDh/QtDqMJDBlRTfjWs569CO3Iurh4Y8DdwvtBW5KWfm9J3OuOQG684Fuedj
0sKGW2Wi+Wq0oZTMiF4Eat+NTeEZ23IEcUA7P5pTP/FARBjeB3XuMYFTr0C/CWM+aLMZu4v2l2cf
JDLPW7ntSepgO2Np9jgS1L02KmB/FJQAVPH/7FKD+MatXSycBnQcRaONtvhYNGy62Cd3nhDrx4Gy
tj1/kdVd97PL+SwHVZ/5Vt1xViWi8DfmcaZI+wkBe7jsaoUZB12h0mamPQmynJOc0Egfu/QChNIE
7rl2hfLQqoS/k1GtElwpBcsgpj7oaz95W02HqGNbm4KVL5vMycROob2wkFJ9pIT29xtQ8bnaxBBj
msIgQ44qebPVvj4uwWwy6LUlhTdbvXW54iUPIfH2+KhcwT9RPwuVo65IvDysmwx96EdDK3T/xxLB
2ojc4F17IMDTgDL9KGh2dazsmqhO/2Tqzp6KBmz9g5+BOdHCRmjH2AAyfLG4nGKZY6P4U+Bwy3BY
TPA6ADJELsWIhsu+6fqiVdchGx+xza3w6+aaoCCUNbrkBJE7rz2IBfrg2NybZMdGRV/XjR0urrU4
Ly8+fKDDsFw7IAnETL5C2vCMAc4atZhG/nUXEX/5MImyc1EHxqHeZJLyUI6rdpMNv5Ed0CEr25H2
Dlab6sxPIQqGWpKKKZ4PKpJwk2s8aWzirchrCr/HMYMW+JyeAm6xpGB1+28KT/0aSrh4TVzA6IHG
+IH6F7MNb7x+lADRIwWAqnr2GEtC1VTLzlYQ7xCgFyrr72PumqwzlE0xAelug4LXGBnSybNV5Fzs
7k8ajDk/im0iNM1pFb23M1f6Jaf9WTs7jhYh1y2jrjO6K6R4PnwjqVXVX7wmDB8FhYufBP/XEQeM
gHjjBZ2JMFhfGFwJxLO0xL3Er+K/ZptscTvgMUWQyNQCokf6sm+vCzVHTK86VBaiIQvemFumlXx/
Dk5RUbYVZK7Oj+7bagHzNjT7nUS5AS31wTdbGs1TfBX3gkNoaFZ6TfrYCwei4VdeZ7ffPbg02Sg8
sZhxMySMO3Isi2l3bkCy1tuqNmnQMboC1y5EX8PyqDBnpbCbZb2JMvikSa0YKlo6V031+ldZbtu8
kLlsNHuuD9v2z6MfmKi5L0wvOGx+x614IyYWQuj+xME1R4DEkW1dm4HjWzo1b6kGe2EYXa4cUFDd
DcmJFWWTaCpHq8vhg4rr+cIKEj8Ahvbbgp7CVD/9S6WxiTkeIalvXm3qal0iQ0hcqcCSzXwRsfLf
OHKL52i0xGLUqOvdSzdhvBxxpeC5J3DwsCuN3d6R8wS3wGNTBXsYM6bHejVywEzMG4KIxPR7sfeu
Zz8pNPSOcuTkZwhZe4BBnguRhLF1/FVongLfOt+vdECvShJOx+yS0Dtc1Bb/B/W2DZxE++w/X087
JPu/xIXq/U1QDqJrI1MKgznFZosQUw8BvrNapXjwOQsn4LTja1E0jvPmZCMGzPWQDUJqt+YpJxwk
12a0OFHvok63Ev9YqwD47NH6lPYDGDCV54ydJ7OqMaBPWuuYpAveYKZEBOJnTSj+jpJTtGvNOTRc
8npDHA3d19pyy9gDgfQsokD5En3CMmsM1Sk7QPnggWDvh2EOuNPuqHSLx+oMMySKfja4o17LVy9P
MmtGHg44OOUW5XLm47V7XcPrDX3HX9vz4ZFP+BfbIQ6cDr4FzPnDDgpy/w0W6BDUafl88FGIn24q
82BYi9SB6JoCAkyvIFkGA7g8PbkMSOliwav+dvHLFXcWRBYTIaE2Il4HAKCuST1fFgZEShwsBf59
BYFNIr4V4FlFfc/oYfEG6rIu2E2XXyXij8qvyKbF5Tcy2VK7mGrCdR0FZMXXpBEHwhieHdeamXpC
28WZ9RXZsXEz72N8iR/37T/MdPnC1XbmWloKdJ/xx0JQ3OA3s6DX+lYkdMVPkT7pAY3fOLbKt9Ve
pwy6eE0oRMNf3dP9sspugbvlFn5/kxn8QqAbRF5hUwHidJ9W34Mhn0vnTS/+aW1q6nbyBqoTuSmE
gr/8Dk6Hy5b5IopTTWlM5EHhitU5Cp59yMsRhD75ux4DjnySk0R7TXbaUQ2gR6sikVf/KOmI9fzQ
n32D4BsH8G/T5NEv/BSyxS2j1QcnZYoyWWcKCoKSHGsvJghus4A6OAareuIOljuUokyBxYg6VNrk
7sYxYdbGTKwTTIqcHg5cjZKJPW7CcJlSRs2lLXAB/odxM+XJwwUO86YUhQdDUmIcWSrTgkGzklmn
YISwKlu653+4YrHvK4hcEGj6jaSoOkVsNNdGjbQyoez8Vv6PyLzHIM6x7ixce5BWPo4U3oo/m450
C45KHGk97LwoUYm8ShzgrRMwehamFucyMPCfR08gNpoNoZ5OZHlIQ6ZnIkgVSuVeFnumAVoRVK9y
pgVk3H0IZqNmTqfwtQhqVlGykhcNoMYnhZtXgGGWiE/7tQcenRPfoZL5F1cbxNt/Q4LnlKo6sNFw
sYPZSDfZvHxYgIrftysERZZt32F5CBvpXEeFdHyJHlH2UhYt1KEcPlKxNZq8LjQA8WqZG1flaWNW
WovMPU+xk1eY0qRVuJweOM00J79kmTyeVLLdK3Se7v9SvxoL7fkJGgdsu48bcJ7nxSQuSY1l5ZR4
TPfjFHIzCXNuahRWESgM0nLJDpO/RTXuhNJTuR5IIXRBEKWTHigVjsHHupObnp/OwuwPnUJhUAvL
n6cb6A542Okyn9STEU1+6VkujD7SAH9jeKdidt+QGizCut1bMciCgJ9T3uiCtYl2u+C8T0zYF0HO
2TqKvLL4/pakV5Ms+BZN7HzlT+zXcgHUTbDSWIicnP1NmkZ/EUr64VqMBSgQ2PwwnMtiXlaBfXqb
nyN6oFshQh45vBy/DewlVpKCxxtJIFqmNNg7OwjcSBt7eJD91yeD/SNNGNKYvv/cm3jIYcvxy6zU
c+Qt5fJrbyl9hHpAKilHClSLEEMH4PQjImOX/RxS2ZdIoDwyd+t1EEjOBTyp7aILiz7ooEU335xH
xYY7q7I38ysIcovfFaor4VxlroMeYO6gmO/uJj1XcqaGBLySJCBMjE9mmE4SymQdXTc84KwOenHW
sE7ngnPG6xQu+emFoXLghhZQSkvJR0fGvB+sI61/H6/lgG1xm4lII/OyvJslVdCQ+8GvEqHnSSeH
ptIiTbgS4J60dFzkjC8cA2PY3Tv3wcGmPYcLASnAoY5lg7bpIOjrGTRyxPW7fG8kNQ+sJIMSSVop
D7tqPz8TEJinfZlVSuQuFycuwidgeReFCCuT3NEgelMXJepBRC7h9O+elEVFJIYCBvC8qOCSEQoT
sum3PuhOgLxZyZXti/UeBFJrHrihZGV5IBwcvnuW1025qlpDWAF51DTMpA/mbDCTyYg780nUvgXU
+L2JpdLmVAXK5YtOX2uvAnfclY1K8gGOJtE0+y/d0NpWS4K03sr4lu4Atd++AOHtUFQ06zM7fBnA
bkcUqbQz1P8QqQaQj1xdlXSzPfD21bOgdOPfGoC444WPx57dHoRXXx5FkcIgKAsU1rwC6VmdGnT3
czhSMYZzscMFGz8FgyKw9I7n/zEfJ21srk7PT5J/wU/RVRb+/pnoYPors3qv9pe7tH3KVqrwTLbN
lbIiylKMb1DDHI1ZTtGHYo7daa6VaHImnVG3mVCrC2hijxlvTmD+DjxaZlatQFnX9+z35OHjmEuK
oWTpw3zteTSxBUfydbCFS/kRZWDM+OlBxL6YOUt4XdUrKNs97QLJe1pBsYXZz6LQqEhAGioMBXYM
85wqukOlabDbUJUaGXrkRcCmymRtGvN1daEn5j9WP/zT9B4vOwvzx2CRNhqPV2mvmTRGvA3/ZHDU
pMKbjWlOyWfRBiIeJe0EvvF6VMtTjZNmfWdmQf2xkgLWXM4RQwE2kbKweEr47g4gjIe8oZl8T/+A
EGSgsVG9O3NhQS1UGyrvIZkKnbdSu8VaZRDxEIL3QpKZDGb55ITmXVNVOJTS9xJhvMc2HruU+rSt
CYs0skuGIMsIToX/k8GFJ58nLy8q/ETSNKK+3u88uyycyxUPThL7Qj3FGVOrh0i9afQxjZBCis1p
iB7Vz6yNl0Q2hrgM5JtNoYf84Me2GAm4P97Kwxs+eXDcVL4bhmvcIFai2ZVnw8nv7ltr/JRCAL44
UFQS2gyXJQ/upF7VhOwndEDlycE/5CzWeNSyqeU9tL7IAN4OYTGNlXSfyjELtNGveAgId5o1KUgI
RmtpcvBndxYLtL19wwggn9yKbJ7PH5ql0Pmm77kSH8nGP9AqThETJHkH+9qtDlnQrMDbSLTWvtb2
1C5EqHzQdrClN1K/963V97Xu+NC6ydH03UjVLaSTIlafaxn2p9C+uuIaY6Ts7BjR+HBmIXxwRGRb
v9MnnZ14jlE7Ow8z7Nvzwe7OGediNCmSOcrIDzBholV1fCYh+ahBtfp9DRTNQ9/MTUKFdgdeeBqa
5mXsEB62r6wFl9H7F46CAFFnfn2DoU3U/UaAA7QcgmX+1GKFMNJDbh8HdCvQmb8kSRrTZj9YwAXp
FHFY1m6quz4r23qH8ZGXXrApXeZ8w20aPPx9WWU/EQRrLPhhz7XBuu5pK1bhb4Jn6jxy8+UsrVec
bBMgG1/1eZoH7KJyIoJx2BFjAzO0ekv2uP9Ixjcjx2Wu4i43xKFSI3UTNSEQj8hhtpo5Z0TN/dQs
20vJIWfKxeI5Ksy/WUyN0KOJDIg0W2eC6cLskNib2DRFDO52S6MfbN794qGs45oCa/T2pqpxOb0L
zBUtGZlFef2m9939H5cSZAHSXWcuTZ7/vqpHoSJJkAljalYxOER/I90NgVaKIVDIw5P7crPy2L87
4qFhsE+BEUgDwEZuX/+SkoeikiRfE9NYYYT5723a8B6h8qVug+UxWiphK/1VGecKyq1YBOXcwee4
KaBj3MNKDjMzHHKVzjfNrdco8oE0LnQMYbWYMEl0aWUTD/tRk3yib966crKYdGLpjsWDvjUHyXq2
JW84pFV3nC/bfL6c+yMzeFXOKBA8vIjD2cGB4AiZPlVxCkBXQZs18ya2KtRO368PTPRS2H00y9FN
RIxGL76mnSlhPV4LRmuzTqt52MYwH1tEx2dig3z4AGDFqWYBS6OC0VOEdY5Mj9/JYbMF1gGZLRiL
Zu13ioIno1q53MK1+0fHsuGUQyxJJoXEBT/k1GR/EDOnAua1Z6woTJnujj+jbehAZM+FuO5Ur9bL
GWTC64pC8fkj+Ji8tWyW7Dj9pCAjMNqw822kiBVb9jkL8e55C1aJxyPISUBK7l5bB7SEIDkv+68m
h2Hm/2XwP30exp4ZY22fWgoMnLiJt3ugPE2bj6KMhWp43XXVp+ye+OuLELo7AOc25EOaYf/3hTdE
JV0g1IFKtNmBEttMzUdbXLBsRo+OPPwDRBCR+6/azih/AnaALl5ITx3G5aIZqWBAJzOBfairAYxH
ujGG2r+ha5a1Sg5w+HJdcgQIqJsLXp0wbnfw04SKDcbNai4I9P5tnKXaWa20ot795V9uYy/ig7vc
dGgvL8sxvbfGbn/bIrfjj5Int0sAuxMYSnWqNy9D7nEH4vT0+lUdIco/VFw5ya2bSQ40aGtdqQ0j
s5hxfU7coIMcNRTYg39XcICD9SDPTthy3UCSTEKMt9ck1pxdatOQCn2M4AeFsLJ3pyrU92wfEqxr
kemjbZKjZ7kZsz6c+mF0/UfZYLtALreC15CICLE78Rkvphexer9x1IOT7B8RQW4wCsnyBv/MZm4b
XfmDG0s5RhUGySx21csy3iSKbObizBAxJHGkYeoCfEUKAryz/1a4XZ4j53uZcksUr/l/xw8eKckO
+gMfIUQavl2GACUyRA8I8anZmu9oK+pIRefHUJB5P6IDaWyVPU6g/ssRyQObfEpOvV4ss7bcOosQ
QsBe8krrQFQ9YgfGraFEMdXVH6NUviV5tx3GwqQiv4LHnoPtgJmzz9c9UXxyYrbiwxVehkAiu5LF
gDB4VdihzmJjDo8gC2snGX4PmsgG2EevLDub5/afgPfmZOhGGWLxXSffXeNwCVTdrbLp1bfHTqbB
MsSdEi572pXsvp3udrsgw5+P1QWYmat0Yt9SRpw3y4oR5ILgwX54nL4IgaLQRYO59Wfom9ibRGKV
sJWL/bCxtqKb87P3LOojxntXKg+9GHEQgZgr4ENGasaNaW1Xlze2j5SVXFC0Hc5knf0s1sLsMP/W
ZMbJYIsQtpzL2ziRI0aLfTjHneI6Yl42tVt6R2/czAxrOJykP5czRK0C515oFHEHt96D/k3BeLje
QQ2QglDAuXRzh85n5IGgXGBuZpZYtpmj9cx8qteQvkzCMRIo9mTwtLBS3hzyRurYMTKNq9BDCEnZ
SGpeGiZdk4MHG+Vn1HzJgXXz42gVrGf+nNv7RdO722n3BMpI9OaXxI0srRCOQbOqF56j0O9OUvas
rtRdaGnQ2Vao+1l3MX8nS8EwSc59WVkfQsL0lh9ZIvMtV4j9ZF47VY6P5aiDn74s8AxxyCvqNZJW
5wh3yQauVRfpvD0kCnODb3RXTPXykFxXdjeArz9E2SfqHF4jS+mTK4ZFX69/5916xefaWVRHA+Pd
dMi6ljA5c2g5miVUgt9of7dWqJW9EyGCpJ5iMn7hf8O7nOMRzn4xz2c4/LoF5RcGCEWmGmSar0mg
lXdcLxMdaQ4tTnFB3g4Q7t4BBdxuCOYHmjxC187aJ6HdByY07NxGwbjO0b8a7Avyt3Hjo69I586D
CtDuoj2W2AZUFbtjrXJMHB966DeZbGCZ5LrJmPwke2bv09CXUF/XI8l9Tg8DrzTgKEG1OQLnBUAo
BWlBC9GfJlYOyXERPW4U/HaxAWSEd07kL4ojL5c0PC5AsnvMiwHUNomCNfFm1UJefJ4NrMTZ87UI
L6I2H6c6yXfDtvGU+tDXkbexa2xXTM6phhH3dIe+pHdv285pinJKK5xUkST2qyjh6ZyzYcL30kM1
gxxXgw2KwvQw+zUseNJgIjIb9xYkwZNjQngSmi1TjwWYZawb6CfwH6o2HXgkRnYUcy/GsJlvuuu6
RWoBBIFKZpMNSuAZ8IrfXPx7Ih+TS1b3fQHgX53WlhawCoNn/mVAn2SHjzYOn4lguwtsiSuHY7vK
tJvL/CQC8N1RkQnw3/VPgj6jfN2kSf1rmctuOaHtsY45cpmL0d+ZGVfh/DDa/s5nzIMPwWtPISmP
w8TKc6gC4LKO14ndGxcImtW17hnx9XGC+6hR4DoLooJROk/yiCeBUKLvsCJLRid2P5J2Mi92NLub
Pc+tUVo8aVSu6uPRLlWl0XK8jIaGegOaSdvq8qDsdjvs3Gv/fAKLMIouSvmmOdPYKIeI3r5mW5m9
imTOmFhHigRtxjjMA5To9XgcY5Sw6brKIs4ThDxa/YoECKI4OrCp23bn/lvU+LsU5nFOU6Gv3n57
NqTq+whUCiPe69XquJXYm/j5GJJAXHQEsA9+wyODm2xaJ10T5nu2gVgtpfvyvqFLQCbH8Mbr2/8j
FoVdbNVFIk2MznDV1vjrG2U70HO74tzzCD14kDQkHqvVoEveE7r9GyXAod9wq6KenEEc0dmpPMh0
NFgvNlZtLKjWd+pOXYZsTN/9QKx/EPnXhNhu9D8VXZRDhJ3Kq4qokwQHdHGl07FXg8LfWJ5mE5L5
/DrInmP09wQlrBHMZFBXPVNb6pM1TZOB19Dr1RzymgSUpZ2+lhyP/JYL21zS46o8WcVsvqHpr4OH
ZD2k2nZsSvbMLv2d6ltaNe0VMES6HE/ulQ0Ro09ZhGMZOgUFjK4+dOWBKKEK7UhwSvGamJAtJM5u
CBfmbmlG5SQOGh8PK/kFVWcoA2/DdlInui8h/qhKDFrUMESB5Ps3QPaCLnNMKSofQFdDZccy5qwa
TawIB5Fnf0A4XcgV2hGdbkwnqA86Na1XvhWywv41Rln3KJmm+iv+MdEOedTKE+kfGnikoH8hInW1
1qz64DkVfM0A/kiWcOucPX+zK9lxM/PyX/3dfxSvA8H1y1DirxF2yeNda2VdAnnrmsSULT5owKQy
O3JCt5jpxXhebA+vUhm2bxKsYvoKF1Y+nUWaKiQyjyH2a1G+UtDc3E+HJZD1XCheLb+43ju+PvcG
IC8Pb4GJu7MbyMy34DJQmUxowTDu2Zu97A5pTOvDzGc8lyNYA8pTfO9kFGia6SdCDM0gk8Mq/Sy7
OWJayCW6Kd6dCZTQCf/r47TuWvGN0WuaJmo9XhnkA5EnapCNGgjqKTceXiuuGowi8d5SGKtH/MJr
UUb9ZyvflY7FyhN9/vAVTv0RnJ0n9jXhrBJHZsjfxlCPT/Vy7h4fylUyhDSs4PJjTrCI/G4jPYYR
iu1E64OK7AlmH4IVXYm9dK84/NJZJCozlHgLRjgr0XTaFHzx/4RziVq61Omjja4gSeXF3FPj/Sho
aTf9tS6fs2UVP4a4SpOzrOUGHHNvSZyPrQFs1RSLrfTzR2FaN0qsGE9Wl/iCrFfO5jMndXV2dJFw
/rQswHAeB6YaOgyjqZY2TKzw+WUC0NF4VqDkuNDsFBPMdqRkl4OrlRzKX+X8zD6mZOoJ/4PkUzBO
cW1CtESOe+IISRJVXrUMsXRnrjjApeXfjJTRd7ZRtAKcjknvxxV2s1CWpJXN/+q5WoxVzWEWKaZm
bsXTLNxxAnIpo0zHH9R1Yq1kjd2QLx8sy85HeL/x6yBIECFSJjjPcq7jHLh+5TUVCuwU8Lw4WsZP
VzgeNBuDEKDEcT9J1uLB+g0dRdSxlBnV5Jzg/DFM2jrMazvnfXCtwchq7l4q8ObaiAoGlyNpe4ns
rp8ZL28ufT0ITC+eK6YOz3IcUCotoEzjC6sDu78L+r+0xQpk/XP5YQJnSaZtzvXSnlNSaf3WWkit
xMTm6Pj8bWtrqIT0MitaR+6kWTdANkOSylw+hDYgoBhoK0rNOORNjUJTESvW/kKbXcb8TSeSdQeK
jqnqY4HAeNFmFs3evSupB7ulnrt94KK4GYLbo2XwY8spn5/hbf5mpFr6+7COsaOE8nEI/BpBqp85
0l0Tgqc+Xk5B2vfhAFJyQv2T04C1d6mu67Yb8ba44Uhq4bCn7a+GYlL+HU8wy6OFcsWGUby4Ybcj
4saRdnCYSnYK+3mMid9Jk8HJTbYrvFkptMCTCHxH9YvIiimbGa/6AbTvFlaJpUUkp/aqUdfSQjfE
WN/T1n13hLw4ZOEWaGnqZZM2AugLei53cDT7ZHncAHchAGL1lPy1/FjaFUtUpGtfEzMTAY9XZ/rD
Y0wNA+/r4p/5G4/XwdCcPXZ6CH21qi+RBAbDT7r66ieZ4C0aQP8QdTej6b8czL59K7buUIiaCSWd
JfX6N/GPwhztrwTxA7rQksTcQ45jFCjpSwg8lstqzruUI/Ko8E2pncntCABEcrtXjVXsDPrQTlK1
7XerFJg8buDity5jThLZ/14FipFDX04qe7w9WJ/dRD5D2dYb3rDITl/w5ugCPoN9velrTxh94HJt
IrGbfPX+ofoyhSOKW84y+y7R45+LtI8bWKCjy4BXRbpgy3vaL55I5IT/HKY3W9gcZ0/c9CMGH3dl
Sz3rItYj37hZseyubXcswPUeSbw4KYQcM2lQPJvA7Rg0zcEOdLCTRZiKG3tWvZIBTKN3m04XPAKw
GPj9uudsUhcq2jyFPmLuktgH+vvuAXQ39n3wfaYUCsjENam9qVoMIf6nCjvU0EqFPhpJ7bOmSAM4
h9TccdAQT0LbP8hcBCUG4Ffj8pInHn0bU5YYseavpLAkpEyxu12bHJFzUXEZEC1NGdDax1zEp5PG
TzrZC9b5pcHteq4/Y3E1EzTZkzzAVrt0S3+UYUE8oQStGxyaAm7847ULW0rC68hmiGWqLMUKFoav
NrESsF9QC6ziw/+YLq9pzkNUP/3URneMHWBHs00yrHHuusT6FSWQQoeDZrkKYH9/AW2qeLPvAZQz
87XcCUSJ7X2OJyEbnfj7oLGenjoXFLAa1okWEe/oAikHiWWS2kIYcd7vykV2rMgzWOiDIV1fnABr
A3Rb8Wd3i7k5pvB0F81vNMmMpm1H/qie8ZXaaXGBOflXehDBog5ePO9h/rf69zTm3s1lqC6GIIuO
s/aoO44VNM+GVmBDVyqc/I0hk5Y2zSbStIlFVhppe7FAG4y25/BCndM856GOhmr4wu2lK0DLqd+U
IwxEChstdqGN3ythapsW2b9Hfeh+Ne/8Nm9NBjweze2QPzPMHgq5HrCeiXfWlyM6BytKPNewfcM1
NKt0PQ0hLd/SZsHVYhoKVojj9LmdBcDVKVgQLaG5lsAsckzQo39BWJOKJ8CvOQOndNd4fZubJwhN
xJ24YaLAnblUAMYoX+GxhWQ+jMsflu7+fHBHSjvHpVtHrZXzDK7EhBC4lPLO/QY9DXUZ+vPswjX7
0mbW2NE/p7p3gZebVXxVn/UN+6jF1weK8SH6IKQOj/aC4AKkTqyhRpSnK7lw2gLj1DA0QjQlruaN
0EEFnWFk43laLiRBGZ2dps31ffuJXFVtG0+hGyEvbz/54cu6gmj3xFUmKlBs9SQtMdCj8WEMZygy
ph2eZbkJF0I1bG2YdkKXBpbghaionfngEZ1Hwu7vOX1mUOj9MZcY+7blNQcFDoqF21BQrVYhbEVI
GVJHWTufaLfWhGhXDlz3G1YotWh4Z9GoH6vn16Y4ilf3Lpn6UrdX850hU8hup1xSFJUUg6U5O1nl
pzOZ77XzXOQ4HpaW/fR8cI5wBORBSITAt+MDEWZtOxqeHOx1xqRPs6tyHybfjOyUaoJ64N/6H/Sw
UFLP+bdQebqQJ8maJ98xHSgp+ucJqiayKNlvnaqAqx7E2E6tFzDRLDa3Pf+VHEevzuCtJihhKNpJ
Si2p/h/uO03mBd6yeajTqA14U6ZEzKMNGpgv9jUAz7lmUpga3Zzn1t/9jnSPpgNXqUnBCzP2zHHy
ZCTlS+vxyztSLsxhdo81vafB0uY4FGWY5od03Xx+z94QPscXZaXedMv7YbCm5j5jP1aULi/ZaLUJ
jO0r0Fq4mJOjPgZtfOPGpyXIfbESvJuoSLhuYFO5wPJrDgDZbE0KILXKpdLgSWfE0vryHT4BvU/4
sNP/pYcBCR7MNWZIxogPHNgJIVKZd27XS1qsN8NOpjFRrb10qNbT74hxTXUqXc3Snu0yh+aXtCId
LK4g79fiF16TqXelRYN7S2hUxoeHa2oTRyaYWHsEL9cMFrNQeXBAbj39nxcJ1recPz8/OHz23Za2
rSV749gMyDLgvMTY7CyZ28NjbX14ka6rOSsCBQjTIQLjR3IWZfFHRFH5THGzRTb8704fKbSrzMQC
yvXK6LCHbplwflSy+iVMOK6KseQfXtgy2bMPR0Hsf2YG3MKojf8m7V3KOQ4YNWu0eZreLrSMnbPO
LK1SA8WbJfhvi5kP3ueI/gT+4xSSoo3vwNb6XLzjmSFYApiXF871ZNKv+wfPJ9rfhpEC540gOBBD
MC4gfELgW7DLGCpzJ35Yu++Gkg9/6vHyc+edKlYJSkAO1YPbNt3gi78xncFANozh5DUiGNTpbydC
HOMtGqEUEF6AaOjCMIad/6BiO/0cReNnvIwWNrL0quWsGA2sil4NnjgXEH9bgVpkOZhNxsHLvl1M
EB6fQHcn39QU+rUBKBD7j63cxolPhNxxib36M4cA/FrP1oWg9TFiXrym9Q1It8JP/VsMwC1I7Jee
YAeR6KDYIppSRO999jP++Q1LBxod3CikrWyexRW/0TaIq/7uMexgcS975ntQv8kFtqETxZUd856U
WLoyL7zOoX3qwV8ZNbgCmF0dFkUQdbcFP6iTQdVlS4mGgp6QhljRxDCmABF+WdEb1BM6dP0pZWiI
JLhh4eAMHUTF237qiN4ZfOLwQif3cO8JYpu/GY7C3n3XX20uiWZ74ZV1MNAo0iiw5b8Tg+8Q+K2Y
MpoJHIpge2NoexsQB1d6JnNO9SDvpB9skMFTw5VJuqe8lLXp4SsfmBn5aAZT6HtNrILE8EcbJQ+d
frE6Q3kBl5awre3Pq3euPwKGq4vRS5aB1hGHqYIUOA7Au/yalOJkPnXlsM3oaehpCHELb1GAoxqU
9ktu1Z3Y9IoXOAWIpJD1Prb9B5fc4kwYhPVBrIggnVe8Hee/zFNiC2mox+99ToR4Xau3bB2t6JHA
stpntlC3FKxuE304/fQdWwnmJmlw+POrU1vpVFbFsha49i5TdAhhWMOYjkF+5UCtjhuctkxdwf1/
voQRLHLoAftqiJaYtc6zPKTCz+4eOFu0iDnodOIbouHnFLG+w958xAn4A7Ba0YFzGCQG9eYBidQL
RqfpGAdO8nPjuePFsbI6ZbaOpxv2T2ecFO8BqRs73+S22r9t65xPIcNq00QHvqcBtePK4psiQgSn
IFv/cs6m0Ez2UG4hH+J92cujKp8cw1raExcnEmUzUR4NOFR9UQmzXvKVs3NOT4EHlaLeDzqwlawR
1Lj+lkNDM5t0Y4+i9bbiyEVuKdgMX9zgkTk3KXgGAQ7mUNMDdFs1K6Q2WwibA+9gAnBxDe9JBiUm
xwufrAwA8UsbNsSyv8tqoXcbjNriDirFN4n32+343NCREHThTAalv8vQtig8jHTGrQnGvO8XeHGK
LqhBRNKQ5/SUn/Mp0bFtTlJVeijzYpWl9uNE/251XTEX+/xKQg6tIruftHtaRYM25EBIH9csKrIh
T90dQ+ZKsgeWs3uuyVRi7quzRsO8bgE+XBroPCDJFwqV9PmOeQoWoQmZU7807j9VJQes8u4FgTR+
o7Wt/qkA5zY5F1G8lDtxbd07nSQQA9sx05yQg3Zu7ynQmmcTuMAs2nqMA5OWfT4d7MQHGfzWcjiJ
yqD0aB5qVKNFhcLeoALIKyQqyQGTfczaftV33xpeMM20cFbc7VJCA+u7M7pn8vxml6VCoqueoHK0
au1pjVLrNlC3Nn5Xya4TBIQuFSl3hVF8q2/iSzsI0+qa7AjRhMNaAxWmIBfmyZvNZ3mp4rbdqbGm
nxNtB+ob7i6QWRRBPq466VB3bHGRTxbzC5BqNQHC7yIpxNKSEfBCHg3PQQHm0hwdxKTGTozDxAUJ
8Z0qg5AISmt3IAAnfPBStvk1xTPiTPaJk0I3ASCfTnwLSHvU6PDwons1a73Y6rWUa3toaZs9/enR
nGzskvFB67BebndJAP3DD4cPVs1C5f/4ikVR1LJAkxpYz0xqIOFCO7hDIpuRo5xat0tpQOtRb3H7
Ya06ioX+rZdWXL4JRXlOPskrdhTEZFTb1BObUCSdqrqcmn69WFnqc639mK0zQUOujT6JMKeupAC3
KkvqMhgqFDzwA6A0TdDPemmwPomX1Ap0+sgJYqCIbJwBFEaFtbcmXviWXMd7g4Iz73XETapLGBKt
qLsdbM6hHyNJXG9sZzzg7afS3rjYStP1Ai9gU2Zoy6S/ih7R7t4rZpKc4xcQ7Ht85Ui+mrImhNLu
0v2vzIX7nzQgJt9o46CFT2H9AAzWzllrWkbXmFkj9tTSOhd+OPILSBT8MmfDp5Nu981Co/78JSZj
pWyjy29+ob4ZeNl2WR/NjLW0G/547liZKDqKoF98HNUNRcVyF1dLHCrnwQpU1mc6hjzrP5y6HZg7
0a0cwrfFxBFyoQ0Q/apPmVh/oY5eIVWqG8+mCbsonnikRsBtu9ZWdIp7ayYkb8thmgrVfztv4FgU
jCMLskpD2MiXIQ+bAfMbON5L4q7KBp8bF6y/Lswxx+4PZNE9cQnjyPkWW4iC9AtamLYWtN/4qWnt
KsK/wskcpffRPiBlltiGnqXrSqHnW22HzB55JiAmt0VB3Nt0NrI4WKhUYwz77ShvkasX+IVDs/D+
n2HvZLHORlZzdCQIZvYoKh1xPBjNcGhdJY+ZvXqrgw/94KkRMcwzLWiv92ginOhFoardRkgeJcZ+
JK5g39w4o3MSyDcfR8BwB7izS+CQ0usf7JjElIZylF7XSrd9nzcWLK/kNnXqz02z5TGO3UygeDXU
epB1TUEDOMzMybHS8zHhS0TxFYF2APOi21K+pceq0jt16kBOX4y1i+IK1Lra6XUbzOa7Ki9q2Evy
c/3C8YJKNBkbw5RES+z8Lv2muOERydnA8G5fUSWLcOtILEsbHcO+tNOrC2xVSg4B9vJkWGwLZ1xm
K+VIau0idECL2G5GQORDLWiv510jDlUp/2sVF0PBkFVA24utMNRT4n+37SFdaigQKOo6NOoU2Z36
RXIUcILo7RejCdwbTYRIgQuAAwHcDWHurWnsUIcXL1oyUJB+EU6mMu4a0U/tlxpGvp2cvrZeP+Lq
mq9JLDF5etrQ7CVkRivajXmWO9s785SC7IoAFSAT3jMf5nVtCSP2htLNie5esin3r9KnOtlNMyOO
2O/S3ufFpTPE7hS6nNuRTGyelMC0Fq8oIvoSZBE0ICHriiDIXGR3KZo+6Yhr5qZ9qJLCS0tnP/4y
8SWoDqIYvGB85D7UT5zd9hmxQjnFOe0Uiu4SrXtUwAIf1uAXZFSEzEt1RILpZx9iJ9vs1E32KMek
HlwYO6kyPr73X7aCIkd27/Qoyy3WyqV+wOYewuSmYebh6CNCKoetegW3zaQclfFivWJe01UZD8Lp
3MGTMQGSUYI2U4VVR8QoLvk27ZyiaOdHWJdlm3sxQfL/1xxOTdDwAnEwEAlGD05fkTy1Vw1t2B4K
pdCKvqsJHdOH52NTSSefEGVztrU7RJ9Al3lsfNqb2qQVUCxE+3RlC41pD+pabc+SzX1UOAsG27hH
xaDzhwzp+oklHo/9cTRSPhrkMY0inRQdxiWX9C8c7HKJhRnbG6qOuzX9ptoaZQs3ITbvOHPXL0f8
K6rUw3mNUok+9y6c1c+oQCpTB5EjT5N6uk/jcIGDLbrKLviSfhtU5Bw26lr7vXCXd6AvWzAvPLLz
MrUVPyXfjhQ887K3wBY2cvGhkVMhXSAmPET97WLYlj9Kyer9Y9a2+zxfnJIuo40JVZZSat7FsG+v
XXnvvRRJnqoC6ECdHuvzf/I3c7wX5bajKuK/ZJAjKcXyhIH95Lwf/SeHUQHQf9r9lCP5V90xuddF
Mupk5nlxkyNrQYJl8QKbARwJ7V7a/OJOHlkBi6orXrXHJUBx0sCc2Jfe1jo65tdn0ulJlxr5jRQM
igp3OWZEzdwebJ8vZ00+CWE+W/7UP/46Vc1tzlIh66MOkKqyBcWarjs7BTzP1PtXSsLTpvnYFrJT
ilqJz0P4Iu2nnp3kKGEPTUVCdlXa+5oeShlffFWpt2noxwBDMnM/AubbKJlj4dLlVzzJBJhIjTbP
FBl6k95NbzhMsQETVq/j+avbWtVvdRY/2Ee7pxeIyrWMNJcPSndN57m3AoQ7zcEZpyxjTnnQlL0O
3Ef4kv4OLsx9budTGDRPnDMy4tWzZB/rf3vXJGjeWZq3ZF3p+8UGhkVS8AAqwIIoNwqGyCPNNVUb
0N1b96K2QcvrL8Voe+PXHFYTa9GQnOW3XhnfV/Aju68ui8zertnJNglJbR5LWco/++TXwOSot2he
J7aOGQDAi310O7EgNgkOUBuy3NQpTcmICAFwngpEi8sgLuYUmKBCFeI+yHR6sFAzg5bIL3yAkjur
ozI4TZDvcYYYhdli945BXA/Rk4KGrmA5PEmpvCbUv/tDlnwJ9tqYrzudSTcLOX56Gm6Na2sXSnRi
HH22wwyWe1oVMt89vtNB7SLOwYuYMLTudl/O4B88wAeQWOv4B0rHZLzQA7mU4NYc94acYxSMH7zL
357OTYyus6FeoOIGw6uqL5yX4izAXjGpBSC8QWOMjjdi0nhQQxDzgL9bLgzr1x7V8FxV6nx/3p9b
8nD6dUJIkMs+PxUafK1naNLF0PH9mGmK5GXISe7byrmPEZ18mVepgTO0M+RCpO+BNZYvjdyoTZwd
rm+NLlTiVdspuPi20xuaQiWfmDacK3B+l4xQwCzeYyG2F+ME7vvWR+vzT9mBHt/adxo2o5h67hdP
BbviTdz42+BEnHsXbzpmw1uODg9QI1ODAP9geEpGKsmEGs1kZLYzFHbNloGxzPT9iMgmaOI1H5ZY
+Q6rzGS4RM4cgi+N8eP+Bg3KoaGtdAVjmt4Mp4zb5ntZW75oqu5dzJRiW6uO00GCYW3FmzNAalHU
3X5OldNoY8tR/MQUCV9XvAfoOmNXPKhcetTsdh1hofB6WWDJHZqWJF2WagLIfE5uO2MR8LMQOgU8
Esn018XpXYkx2VSv3W8c9wmDRo4yk0SFpi3XvUMb1mFWCq4qa15q3LgHRauVOOuGkD44rfw9Guy9
OAHHp2TTUEMksXBQqHQIJW5wVEUKWG6EYfUslN8y5h5rmH3AF7qN68cYmd+mXIkoDlG3JRcMtYQ8
P/6OLgSL4d0FDuZQ1CnrLzwY4O1DHuU4BkevS3j8F3k8UxAEANr1o7pFlA2B11ENY1sRNCExJiCN
JzCHmtKM6S4RIV01XuN6kk1lTjCGtjSCT6YEIHDK1xoSGCYB9LgK7bR5V0F81cP9gwn2mbaxENBh
g1wnQZQJt7DZFZEVFzTkhTrkL5cvscnjrXhHeY4KKhyr2pgeduD6bGyZOOzwLnYdL8FlDRykZIUz
BkfrbEqWwiTIiNlJurYP2wjBIJDEexsnDfApwcTcYHoaUnzRwgrfe6hOOTTilgmmNSCNcgHN8HI8
jR3f5Gp6K9/lMz8ewjrxaR3eCCXMeIMp+seAbIbu3MhebO5eefEZhzEGObslIKhmcjTu4NdDYxNb
7IXAO62QedMi53jGzuPO3JJbxXtX2hTSPjVoo/1fkb+b/2pfxbmHE64SvV/l7g9sDusDPxKpLDeV
/us6FLgXmXpvRirWAD2TtLv0CyOTigt/rG0EFix7iDahSf/7FQRrMsGbfcP89s17dAzdfVJEgrJF
W0Xq26o1HaHvU/loRwICpYioJGskeLyhBH6BmS8qqKSk0EzkBSOKXfPn/9WzBn0ef1llla4eWmA1
bm2X+xVMa+w8dHo5jzwdwSTM6xOBvjpneNAOJDMOXUChnEUZ+G6g71mphDYzIWfyOleBu/KVn11A
3fn/BI23kA9RMZk/PuCzRRphGHNnfkUcBztWiNIwZk1PjRX/XAXFrd/QWpxGkUGNjLlTKPpVUwfr
SneNgUURhzKKoxiwK8+3wuNaGV8WSh6ysnsDUrrjNIMRtWE65i1VSFwsRbSFV5KTKUb4apV9ruIf
Ei8Kp6gShtgkmu0MUUG9L12MemzkLz3VuHeHZlAvqy9VFdksVn8PqbByj1kp484qEyowihlrC8uP
a/n2UgaFtrGYuvGLHzHK7e0axmT8//JivqKLfdpno5pzpVnZxb/SXj3DbTsAAdCkh4cveoEa6d5E
cX32SvBezJ847AHLdk6ZIuknaVa4R7VaejKr98V5Kf6f6OhLKvSsUlaLj3OWsttUFkwrmjNzXeYi
GkRjSr/78Tv/W+6+8O2ZnP8/RaHMnryR4tzxYC3eFZyiXm0oJKNnmPIC7GguSMGseiXaFlxb4vqh
u5BubiTD2oJPH4tfj7Bpvpw9QcWgRQfMKeCgjxFbTWJbN6TU//GJU13v8/OODv0D2uFu/1QYeZKl
UTnP6jJRHmRRikWKdNbBYrL4PXZxfFokyrHpvcAligR2iqJquGKjDnsqlkzpcnM8XZK6bGo4/cvc
5iSCGGy5I1vJesj3F315lOVgHc08Utv8hLgPKkY3Ec929mAckRVjIpdg1hoL1oFCxmp7TCt/Vfvv
4xHsRy84HQ7aa7ocrMJLp/W/Go0/g0fRJhDBbXmhtdd1qpGVrBX4fUsS8hQltVheZDTYUAY8Vxa4
HkaB156+HIr8DeDEcQLOjUf4nyRyTlI7Hi8wqTZYEzHmEgiLHiyCJir3rjGRs++1e3WO9hcsHVW4
ikgVRqeZSl0erdSCjWcNhlxygZFjg+RuVsFlbZ993feT4Z80Gw+xchR5x7e4KSwzgbttw7C+lvvq
tByKn81xICXt4XRvyXUwMxsBAcTbzBUAJnh015yja6O7Pf3BFdaZ/ockmNBr9uvxDBHwkqohJdbD
+VKTeMg1gz+/ICzchd86fL7eEaqGfO+AVlt3kUfK26fyKSMfvIgdHMr+ATN4ekLZ3CUeCaR62CvN
j51MjnUVxRfEtCCVgjWhMeTiDcInHfH0ZitDAuPf2hDXCKVrfr33kP78evtDTxpFVWkNvB/3Pi23
qeuI1H8Nc5mSiHWrlORd0YOOvruEyVHx0COqbr9L3mv7AG9/r1ijgM7EhFq82mOmlA4GDz0Y5XgE
0ulfu3mfxRBLOPKE6MnZ7z/p76o/ea/wXgWq7HjVH71jU926Z+/1/iwSRUyCVmFcNzPYpX88y/Va
cN274yJcUpECWmESDKnnXziDC80EVw7WkRkecRyF0hrgg4dpyQDNTAQs5CeJLtv7cb8wkxGh4y/x
6hxbGXYxwqp0yo2efhzLgPboRBAQrKeB1xsouJIvXjmuHwSulMmM2IUrL5taIHvBCRcjebIgTNa3
FCUSszyDB7DnbtRlzZXsxekU7PHVL3xlMyQuH5TF8TLQFdixfWLBbrZw+xDoVDsMpNCxrAerZws8
awmbFi9N+O+zrHjO+SgcKuSxSaGiXYjJelo88hyE0g+CzZXSRLXRsYQOLkgaFWLPJvA0JQM4PlPg
prwCSxClL8XP0esCkpxZnjAiuLMud1RCeQ6d8xQ7mgSlbFubRy/e9/RSzr37mk9UOZ98G5RwpKc9
IGExnoehMTO7Jm2xaqPBwPJra9Kxb0ImUr1Hve+ynC/WSujFYz+18b43SMDI74wj8AHliKwDhT32
RnWdP51jHh8Yy058TGJU4+egkw5qmBB5K1MvfTGYZVKwVhqy9PSRfkrOblAKYA241bvIrn/SFhCZ
zxoLvLJhk4QtJ09xrLToJGKFKPkB2gMqNj0BtFLUIhCY99+F+gWXUA6a63pIcMJcuI8sXRyG5HqJ
FuoTXFdmfBAQMwOU9SIK6+JU/zyeG9RwV6PdK8xNTnbEBPM1Yt2wKxwlvjZ40CwcWdE0eYbjySAO
lzJK5w+YGa1Fso0RXuI55fWII45KaRNBA5VcRvyoHIN6DurilDr2bpOppJ/15MfVSZqwHrOJAOLt
LaUoeD/YeRSMMPh7nUhLMaes6j2UuaW8AMHQrctqyX5rXSjIHJDwL8/Owbqebrz5Q4D759OM0cy0
ijSYyZ3mJ0yDMRRhzp7J50fx0u7E/zQMzHebvCGbNCUDPNmXhLMgqlqefjV7JVa3IHSOAfGiF64n
w5X4gi2hmR9SeBDiOPO6sqR0aWvIJj3NyDzdmYJGHqp/g2cXA9+BF0T7G0B4bFaVhXd5qCvJ+FME
r37jPAiMIuExS45Z76MjQ7PLEBFjsR3/Rd0xXMVAzF+vzrveSHeAFr2JllNqByXXFZRpU67rDyHO
KV0E8BogVDtQeemmOzrwbjlvlqIh5P8htB7PloC3i5RGVBVf1kSsToqMCXmWCEMGn3KGRU43mWVe
YrMoZFYRjjH2FHj/1JJK043mJlvKsf7pUUGMmCa4CthDaHaDXExIEfwfEOGPe+iAkSWlDUOASS7g
dRZWtctutZsj6c8/L+aI97hOhAL6qU6KxfE+tDVzdYI4KQgegiy+mLBZGAvbfvYBDIUgBuBw62oW
1SuPo8LX8TLnTmjevRCyHRJuTswRHIcW54xr/K88KhDJEhzKkXA5PyorLlqliQHHTaXxcB8fST/M
bdnedtyn9zDlsq59bHV6AiL5NY9LiOzvRF1bOdZkqMQkSOplrSqfmQ3ykM2FdSjbRuWGves8ZIkV
Mku2E140j7bymotHe9sMH3iJbtE1ttYXsNWEzebNOhJimLED1QbjApo3DAedQwXujo2BOkyXGtDM
TXK/w5aUSAHUhc2F3KufN5qaZTC3LsG9sbxQbQAc6D3+iOtx+n8pvrm6Wk8o6pu5lImnf6FVR16R
/+fiKgjgOam4YcTFZc+DZU1loOzWgEet9OKS/TxpL+9trs8Ar0wj/Uo9ObbkQPLbEi2+RCWxESqE
an99VbroWPDkaOpMdLpCSGlEqA6jwt6IfH5TvoE9rBIQmFOC/98TNfyUAUahtv3/+gThUguU27RI
CHiK7sjHHxBoEnav0lnaAniS743oZX9MyP43s9sxnozP8ukEDtmzaNgejdQve+FXxGfzujHt8G/i
/7bo/Prqftq0Ioj2oE27dUxPS1Rov07ZhT/OVjb9Kl8pj6Dw2xpPqJ9kjy63cVys8U1fbzG8Z9WN
ojB3VU3FyTOYAV7ZJ667wOSJGbccr4bPc+d5feQanJBpkQCGTSKu8meZXJWZS4iNJ958qeTNEujH
Bjq3UjkJEXuNycQB1QGmAUuZnt9Y+4/NY6szfuTsH0VxbLF9pJxWpvrKwDvgsE9PDG6ah7vpQaem
TiQAobN5HoRhMEIdd6uf7D/F21I/+w0tKZrilVu4ASBxhN6o+l8MCzVO37jPEm7fRsOTtmKkHuIT
DjspSNQJYVckxYPPTmoOA6r3hEsaGoBv2t2xrzpeZ+R6tXjz6X70W15IbWe5BuSvhhHCkv0FPYUM
Q8LlT7cIGoGPrNZ1vLEg8JNlvk+Ab7TzxiDDCSB0i0+HFv9QsujNWf91Uh4ehrWZ3tI7sLplioBx
x0CcxxJ9RTxQzngYHR9oDFCowJPcCvLkyD6sS202OHy4AWDHo2721yEXXLRC19HT7ti3t6MnCzNT
+Dmkw9uJPAexGAC8bdov2bPMB40NLL6oSpzPLulzqz3o7wgap8+TFCdDDmb5Cnt34nVJGznZHFaT
dnmMtKbGFMwLxrw+ynLKUAK12w0t3YBZx3+hOdOGbWLkoNvzQONuFXoYyVeyQig0s2qbq6Q1wz/+
lyIdcwbm/JbH7vHExwZzm35xS9qdgTFXNhNcOwsx4UYfH6p5MvvPiV+AGnYgevhq3MIyBYOqLS7D
kh8RCT4W1Ppf/128YqsTeriV3KcuDrOFg1nNKOqk8G2CmpD7dEeC4S9+uFB8EU7SLq0oWXKZQL9P
ftDFqJEsdtRr/MQxW+IHN7RZX8Fg+ygqUGKzo12ADlzevUcIKTSo8EtMM/6MCbhgFa2h4bF5a71b
g9GWurN7dT/8xCSgz1NfQkVq4hmfJ2ykSRkFC7ru/QADLc6646nLlzF7VgwCfBXiDg8SzCkxblmq
NJULOkJwNhWrqKnREuvlnCVIm2i0z4mMgX8lHsOLqkSHUZQxeOZTfBkZGeZ4KxQu865P/wXoL4j4
DRU86jEbAXxtTekljIRMSb2IhTHVaIHW8uYvbdkGUjTdhI59PHataJ0GgLcPbs21af6XR3D2T8PB
sj3qUVTnayqByLF7xgAD+2namYaB3cqLke2Mu24anveT9TB7oMU87902sDKJ/TYkEwuV05eWlR/L
aaNZWBGsgC5LwwefQMvF5fuONvCdifcehDhnGAmGBnJ8nxAtuna5QBeg8zwcps+26AcdZlMuMRgN
Cm8aDq5Re4hbpsEyLfglTp4fV4GXTdnkDeEqz5N0n6oqErVl7JlJApCX2w/KeoviXytulHdcFynd
JzsnKuHyAFfDBwDJvwSIQ2BKMg3JQEbpVvWLUiSAFoW8JYMAn/IZmReYQD6SLn3TWJ5P8nQ8L72h
PHseG59VUyZz6RfKL7gfqJEYAsJAPceHXcOXB7OY1E4Tge90KZax1cCl9JH48Zt8oA+HRiFST+xd
Ry5cyFdVRvnEsnDtDN1HTHo6biQzPUE7JJmSIkUZUpK2EdY87hIMUbz3/W+ytDOk9sQ1xDF2D4K5
PrBugTRWF6Ox/FSjET+FDFAyfq8so6voPHVzeuSb4yhchVwnUUqNBWkZym9f822zbbUkUFrrxeFI
tliSs5kn2V/nHgNZmV8bAU7O7wK3mdpEkDHtA2fX+Go1ERufZPCTy6af3SAp5B04UcgfTK45Y8Mn
m4wGl0fNk2ePExJl5lMEsww5gnBtSkMIa1SA3fLe5HXLOoTKi9ppqaVpB2yh9VffQwymsaq2BRZE
tFuk9jLTnTJTvrN64CegbPpC6u44SCDxD/Tu0jlt8+MHZBZHSPR9Jn1oLKlOtfE+NTe0z0aWPc8Z
8j9P9GF8J+DdhAO9t523c8GVj3h6GABPbetEqkQE6hBqI6C9uUMyBNtBPeZPV+Ng6I+GUTxmeZza
J74SyL/scle1ExkjCmpPtc5lVQ8XSVnEFZ1NdAVjerrDjNfcEfUowiY64zrwzPJ6TXd2QwkRLACj
pp8Gpy2Hgj+aD0ixfGrtSWWC35jexyUKWlywf885hlmN1qahEhU0StXfLAhwS7cjjEx/kFnlcO0n
bed2Le2zsHOfyZQmOvFWanfO7wCc0twYRDCpH771NEueTnQLlgVZYZXgs+bZjfHDH7YibWc1CCxA
hsev1oUFYpdAfkFJd1oD0lC0xvkKQBTqWuhqZzxduUZfloPhB+JpD3eUqV2o0lJpOmj2pekDO26M
XdDDcaxLkZ161LwyqTIEEb7KFWpRveb58nIgpHLf4juZNep66cTJuI3YSkblDc+0EkigWpTel82b
1a6nlP68dWJHcDMXoRwFEnA0qNs+7h24YT03/EaowQLV3ASvudJBO/kDR6p4h4Vmur3INXq1qXdp
vR/nOYijAhLaEQ28lACLJDfvotZr7rQq0/OXqeE+SaElUmV8aU0S2Bjxh0mMjdhurIbJpyeRQNFg
Iy2SW1ilQDlFsMaEKaKx2ydLESoJF5OlaGnvCcWWzCzblMZqkf4dnnvn3Xy0XjREC6unChJj1T+f
y6yyJaZZ39jnEnv3lFE1SQnYbm9QA5sM9SqClo/1sBX+zSP0yQPg/J5KsywCHfSnD+C4BHDmvmwL
WbTlFXx8N8WfVESBq3xne9edFsRCkxyZMD7huSY9T4LLzhaxaOlykp9Ce6ZFnQS772t4zy+TTaoe
kSdLjtlstO0+Df/eCzu8nhlb3NScMzK+9AIgYwEeV+wDOcCGJG31KtsSHO0L88AJzl/Xbp8xw37K
lIoN7nUwzxfnUO68xtR5H73Y5DGrJTSa6WVSUhiKby8/2BiC3suvRZ7RrkS2A/x+R/t4wBYF0iJb
92D46/THv5a0yfsKfDv+xA5Ce+nmCzi+YBE041YQch96ginROJSL1O7y9JdwUvtNpmJMFV8CL4yf
rlJ5G+RByEzxrvSQ/PZFGhBFVNYx+Q62iR8u0krRoNJZB4rpRPd7PsqeLFI390xfdIO82r0Y/XZB
9hyrd9IIELDxHYzYmJjZ9SEeEVyw4J9+03aEWuPeEO964Ds5UznixWBI6QN6fa0PpIJ8Oa5FL9G1
Z0CCBLGrk3sePqS9eZ/AIz2axiS5+InOokxwruxG2M5yZWHe6MFiF8y7MKTLZKxVUdzX10yvIzS5
N9tzCfCNBpbXKuv8lLLnc6Qz8eCkK2A4BD3HSfhZHZEz7P1fzYvk8C1tadb71MOA6PTbv69Kbk8b
3H0fdg23PTDwbYT2/G2HGfACxqxXfPJ3Xe8vMT4g8W4cC9i8VeyOFYOb/7gx7oqMdrFE30grC9vV
owQl/THwTSFnH9/uipAD9OC03QRVvkHTr+Cafa7rqoopzZoxhhJ7X8zKZWrBY5HE7Dq3CVnYQOx5
8wyLIQ0GXgNgjrY3Z+1LGbVfOsaygECNTAjTDySCPRhEx5BxOrd29ujijHf60F/p9B26p29uaAUO
QABrzPzxy7VONXCSxbd3bPp3rsR9Emkgl70TFjPSpNHhwZQDuPFddcC+Jy+kQiwGisVfOC1hKVpo
rzEvH9+FuA2Vocyio0fTN5WhY6n93hXpB5kew83ppnedYcOR69QL3T0XQ6P9FpIr7/H5HSDUcOP3
gXdbtDoBenqnsm5s09Q1yRBt8/gEK2BYfKPqlUqx8zLCJgaeY2b0KUafiTuvHtLi4qNVB7pK4R+/
jMOQVTScEc837u+OiEEz7bhbW65IwTWd7pCF88UmUudxgoiXDJ2+H4AAHUqrvrG2iWSRyOqOsj6m
XXippGHWJ1dDYiWmDjf+S+k3wXMuAUQQrMGgHNass6yabEQ2l9CgDopMrpqZfwz7X9X6UX0FN2wn
/hQ7y4voJAotMn9xPs8x19YKEEpfqn3xqpo3pZCMrMZNcxS5h6B0dEMgTjCi84BaQFOXvZm7E4y6
GfHTKEYineR2g1ZZ7GwW80cQXOWqzDula2XvNft8fgZu059AyKfGsTzTpFWKwLn6xDsZw0egrdbU
UF/CBn0gPF4Uf1tUy9UnK1S7gonWBrRfow+zgclZhR4q7xRf1WgpkGZpXkyA3OEmWIXL6ks3ECOO
fJqEV8DdjAURzSW2ff//2YbqHQzqxGVPRgKEK4OfnLLSeql7gwFc1QpbxjjZLwgAWrn2OJd3e4LG
F53eYjHJiOFkUZd4mIAVFWWrf3Zucjk8rW0uSIrJwlN4y1iptZGbMZy46KexqV4kl5OzoCB0jcfh
5jA17yJUKH5O4PlVx5UX2InVtKhxbZ2gfxsz4/xEAEq4ois0XSIjm2cgfCR0TzRlCCe9EFlRip/j
raA8fwjeHK73ueEc63Q2CAxMi8ft5P9m2n5467xUymKNyy0w4cUdNuKr+OaA5NvqceoevN5hbjzW
7UZNjmIJrsI3ALCN0OL6j223bWLESoEyQEGD4JAttD5TWl3i1NjU6Guhbyfy/0OqYYnl9ZwBA4KX
JrSBlS7RkLXT7hAcH/jN/Kfac0lJRjCKF01B/t3v5wClGtc9e/eRe0aYzcRjrs7VTctvufb8P/LH
1rjtOEYMEkAHyEe/uWGXelU/Xyxtr+o7tMK+0Wj6aOec2J4CGUmql0d/avAHqZpm9mYX3kn/qXhm
cDoK465nc8OhjjL/8DUzyzNufmVnfBlMcnYsY9f42AnOz1KuDlpETCG5EZv+G1Edd7wMunCSavpL
QEmJyVuJLgmUnIWpVd9achfg5JkLH0YwAjTyALM0Z9gUq5T5DJWr6unXgweXKkMoDhxo5bpmxF52
Zg/Pwx8YMvuDMCBPVZPeLsdjmboInOFWKFpk7TCvZNNqFdsKALDF/Hnr27x6EM480j6UY4yigD16
N+VB6eEb9Nv3gdaTfF6I1a4QeCj3Gr9znRnrYm67FWspsxFv5aVwz8sYftGMxVmZxed9XVi6KAfZ
AErRDZhDqgFDAolFvHnfXE4VyiyWNmi5tKoRd3lYHGd7HRYui2jKO8M0/Lmn6ZC+IPmiRBt2obh2
yCHpnC4RSxcKKeFMDezjx3xxD++JR1UiMqKJ+0KX2xJlcRAfWwDBDPhU3aEAE8Hf2Fg+X97kKxye
AVW1t5Ezf7rafJ0qIYftXhjqF+I+27LDny1PZRSdlR3xRpLzDedKOXQRLldP0mOOH2WiRoEwIIng
ooV4tnzNyd8pVfNqWObJybAuXw8rvf/hEXD011jrPiZrWtxBi5Fov823SMENYTB8WLDisKZUoUw0
A1WXooUfqUUWFKCxP2gBuq5y3f1qc/YadoLDIaSeM+//prnzpCym0FkRcnTsqDybz1TBTxejXfWR
WAWKjLVVZxujdyM7mTAWgg2jA561WxbA8hNZvw1wWiYzMR0APtzCg3CNQxLq7D3aXrh+1T4eEocj
72nQh2uFqIcLFbwpjC5M4jqPBzC5EcNoWGICmRzh2rc128plv/ThKQx99zzgqued85DtMHPnqb4Q
XEJ/DAKqd4fuV3qYfww/PSXdOFXspO5+Jwubu6sPHBY58JBtOrc2U5e4JB6JnIkrrA23U30GYKlT
XK3qDRPVqVj8wQ4AgT55mGaaXZZCJjq7I/CXQhHjn9dKKowL23WU4cpsF6SdWkBDLPrgKkCSfaT0
nfT8GFyh0j2d9nl8CieaoA5JNVNqgovDkDg743dIYeQfikurhMuNuYzuuF9ijtG5JMuVdkKYc4/O
oAQArhfG5a6h+bMXx7DU0JNmTkeh0elMThJahJdX7gvzTH7vRxw+xv/a8eWvBjdOfLs4BdFULWec
UTOCUqLTp2P+cMqOIe4mK2BV6+qq6/4EhDj0HRhLiJEGnaLQuxfr3ZhurBzqWUaClWoo0UIoSngv
Q96OaPNVGy30JPaYsbgz0pJHmvkWExzKZEplx1LQ8cpKulGQR8EQwNOzMwHBH+ajlQSlc3Cyimbl
xY43ER4GKMMhxSDQ2yE1adbDkmeebxhHHwFMbyMtFziqhbztIP1I2ajiwhW4NBp8R8NawIk7LU5H
xu5JC0MNVo+ge+hcb2E5UQtdrpzdun1P4hQwPkbTqVtJF/9Q/NozD8DLmBBk0CDnul1jY7wsfse1
XwiNsIcmFr7PDdhF7sJZ1s/k5jUcLtWIDAFuQc+nlgFH5qfqJ/pKTF05FTQenLwJbFeWlOuG60sN
FSTKNQ77wZ9EZgIMQuIBSWPmfIMr3bube4feymVxSsO3Je0kSAX66Ah0kMou4DnpG7WP+R7UJfxv
SVMRhjnulM0eCZKtWeM8unZ4LW07QEwhqbspElfvrWLHiHZLRGmMFCAoTmEOHiOEj+F6Bmmdndcg
zW6At6I3isyrGl8OmkfKR8LORLjKvkCW//Ow6+tiY9dwdfc0eO3lcebyqp3G8IHAxfigoOdrhxof
7fCKd+baDJK7efiBbCVvhm2Zs132SsLhpQuhwzzyDHLPHq7cfmX8Xq3XYblmgG1uNrE5+JiZFqDO
k27GLu7OrPJ/dGMIAiJ9YRCyivlwOmp4ioNAvUiM6kf2h/gDBDsUDkUshJz1f/sYsDulbrdHO7d6
zP58Wr7qe9krqArUap/hTcEV51NRLlKF734XEa8kYP4FMgzK1axCfjT313u8xcZgCsz86jNqq9uT
VOoeYWUO/2M8RQaHPoVUi0lh4b1TDTWyqz6YjIHn7S1g7d8XLY8vce/YeveQpiwwS8EXlInyMDsg
zXrtTrumtVAY1ccQCFSJIdSXEHGPraf6wkEYHopYfYup3viO7jjdsUp3X93/Nmvz5sJNzkrchyvr
hEOTmt9/kbfrG6e0hcyrUvzhJtqLgOH46KTkvtuNcXYuGBLmI6AI6xi4//F/6EJ0EPFw7T/84Ty2
1BRiP5KCJHGs7l+/24BrxOOWIZ7QvhaW0BWnqZaRsjcUJaI54cTQd7AYnb7CHkJ8e8UFTp/XFaeq
pk4CcP59tQ4c/s2w55RuZ3Sq10L5ZuhuK1+JF2/aTRGDrT3158qfOFZ8e7GOW4EIf6VE7QwAlTS+
pEUk/SJ4VkyB8XTogDhuNVn7gUGy9EA1vjypVhXeFUKojw1HPkPj2BgmlpHkDVx1V6xTt15Zn2QB
RQkL6JwMxGPy4o6YS5Uk3XNZ6keLCD0h6zRzH8SS+Wq6NzyMTjIpRA9t1QFQ4BXSbRxBNSsllPYS
1lFsXZR6Sb9/PoNkFrg5IMeAXH4y8tJlji6ey18GaJUZAAE4/U1VRuORALbBf1m0zWoc8qALVmRK
4LCIEwRaZEAdWfoaw6pXN8AJW0Oo8onNOW6j2PSRpRrsWKGwlqQDQyMQc5l2/9E+rc01Txn5ja9B
UFbgvRZ1S//hU5LCOxgQlSTKUn5LYAqSvGEdxSWjrAqsbx2h3EiyH7c2AvDUM7LGrA/47bOiv3zR
nCJJdAnzUrk2rsrJ81gjQEkKZyY9q2swVDRu69OdfrCDBl8DQ9cjwjDbogwV3SjmHFnOhIztUZgH
AJhZarGvJAjvsYr20Va5jxsORS9/L/1mFZj26tcUMVbPMf+l3Qo106ML+lpLyYfw24n4UmmLCMUe
lVD3pIx08vB3LadiInPNtCdu8a2AGsvzwxKJ3tSTqki+M0soEpF2fObY5bxNZLCrfPAPRJpqIgfa
pNVwL1293pRmiy7CGeSZtKtfNJWwKmSJCrrIaexSjjtARLs+6bb1IAWnfI/lz/bi+0QBuP/wjEmT
qCAvl8sIJWQKkEnJJa6/87i5sm+yq832R1TCunEzX0wV5WRDDGInzBlwWCgvUOUMHLkNxiLqNsYp
dXtE1xElE7wG3F30fAcDrJoOH3hW9+CkZygjJaa4FPhooqKXyNFsDQabIzhEtT4yUdHD7x2h0Y+n
MCz7K5wWxdInA7RJo30BW9PetA9Ed5mdAQvLXzHZuNnK3dGv+oqQHN703+vbq3gW6WJxGOkGRs1O
DwMkMKDmSt0HjGp7msH7+J1ZtlqhojOIItpeAHn/WHHzj3sVChThjgySQnfdyMz0l6tk5P1l5WaP
d7DzmuNssbNL8xNNvTOMGnMfyvI8qhPTrshgrmGA1FJkAfPVNWjZzWvKMNGr/nR/UTivVhdPTEDk
vG/Tk3g9rUGQ++wWlzVwStGOjahUcu5bAjCnJTl0Probb9QLpvauqyrRO/elnkvltPYaIZJIktbE
+o3DHLb6bvWZKPShnpnUPMyBx8voBg2pSq5BYHEssm17dMF7oAKQzJTxKebTuqy2Nn4sJDp2CFuU
Py4+nyx2p4sRB5Fv6ZORxPRI2BnMe7Pn4g2pJOzXdvHouiVklMCEmpEzbrfSaK1J1EOYrVeVA5a/
B1aciKL4sDtO65PRdORGDl4D00QS2ZpYx8gsTS7U4ChIX2sRWi0coiEJpFKq/Y9XeG3F0j+nedaT
R8uc30Otcy/J9DcRkcQv609Azy2wfvWPjRlfQ3WmCqWO77Y/iMLOxLNY0Yprdqz4xAj95W8owzKC
3EUdm5yUopmBGVq9sgStZyIbC3+Tcy0drO52kjg6KTqjGhq/y3mnLRkqGY32Nd6xI2B/g2MClCY5
6eUxV7qvSQ3UToIzKd9dekDL39Z/mJCSfptbqRy14OGDkxmX/Nsg3XH+yq6vFolqCjvyTQoD+77x
ZGe0EgBiDHgxfTJZsfWryY2FgZ3hvyOLpA3J27WULbwU8OxlMtlE8az3zkLv7q/yzDSLfKyohOLq
Mng0ZYCihxKBaoZTB4Pz2GP70zoJzJB7euK3BQOeqg8RfSPY17f3WQOgL3YIWkMtzqshE0KIlqf+
I960xWRdEYtvKit7rzNFWxqrhU+HnyceXOkkiUtUPRaBvrE0GpHirvcLBy7KfL3s+YYhUSR2M3lS
9gJrpkjoEnyIIh3XfNVtpTCB/j7ebTAzeQrH2eMTT0WjkZu+0Fp1YlpBz+5MNo0QXR59mNrDl2kN
rZIB3DW2zkOfai7DAjOmpIWZNNROalLRV9aB1mBN8JfcRPXZHND7K9PicFEo+o1MuC9DseieWpab
lCxsapqR9PTCQPSsSTjK+8/Su2n0qLAsT/5p1P+ICATA63M+BYQJ6EV/CkaI1eZqunq0zOB0I0OI
hxCWljf6ZpbjlPJQGO51UOgnYmuZPKo4NpAZDUAeIkiBhQaRxVo/LE4jC0axYCnPN7HBXamggj53
TRrKpHOj8dC3I6NYZXhW7h/IssqcrPWdIE0PK7q6Pypw+IFdHn1ynps2LPUwoxptjo+rEuucL70d
4EnxayJ3tZDIBDyqC6WN3Zwh+m8Haagsu7SUhA/FRBr2KoXXp/e1zPYDW7F9j0Lii6LJ8yM77QnS
rq0lfyAWdP1DYBIioBSWsqxVMWkqWAmljMGuBXeb2G4u2XYJqtqEYR8Dq4yQJX4OBHuk/AESsd2m
dKXioF+2YoA6IA7mpiIUVMzZUDSdkFJn7Kg3SoHn2CKIii+s/dt5zOUrdDP+mbdcsIKYFeQpV0cI
ZpFQcBylL9AL75jyVAc9ZX2jIEcefhsf71W1xn9glUTk2no2gWHOtbUyuXw2+krwu9HEVaReHGi+
ozJWERpE9NvUKXas0ZIGgVyhxvLC0XJFk0GwGK6TRuq+9JjJsMqcmwQKASX70hSrHySxYIgj2GoI
cU5YS8geTtRw4gXMJZKe1kznOFOn0gSL5TNjZqolLenZN8vMdDchxsa09hufpIJlEx3HOW4d31bK
WpP3sOoLXOdgYiH3u0VSyGqrpN0LEeKqWXuMBkaPgWA79vOMclHPTzjvurssQBjs+wGJfCk9sKFu
pdEwlEfb0N+46jcypW7CqgJFpIAvl7bjf9G/13IlSKodOTWQ7gGZFgLZ2wMlucC3dcAzIIS+b26w
rdmZV8y4dYQ3Vl3DzT2UCpFddzIw4yuxNh/CAjior0aRw+azRAgD3eO2EC6y8ZdK9qv2smpgONiE
SiEca6dcAKtR9n11iQj4vEvg3J/pfRlLWoKGHuNcLFpQMttoBs/gPnMTP3BTNgdWFz+OmDHnDgrM
Ym47CzRrZBGHV74cfcruss95nmgwL725Hwo9dKxZbRjvUx5PsJG83Fy1WqB2DRwF5O4S/llew5dI
pxr2IgYLfBgLA1sYEUyRb2nXP7MlhZVTtohoIuGuK0JajPkL/mPyrO0T+R9IlQ0Ng1WW7HmX756A
Af2BCSqb/M7iTgCohppQ+CoDdMzudfTr0sSLhqIIfifRGX9KKK/6HIQP0n/7P5EMZG4+rh6A0cQk
DMeJFc5RK/bdg+6/S8+jGGYhSL12QDOtBgAuxXwSKO06liH9XezXaHA6SiGEMiaOKmiw5LGxvzx/
Wt39XnDtfKBgdq+nOj1FFFMHMQzDgwjdgrWm7Px+eSMQaFz1bksdXRlXKyXFzjPXsewn05FrWlCJ
lBKua0YSZGFhJrvnhQITQt8Qp+ohgbEhQ13aDHNd4snAtPuqFl81LkGRcJ4AiauHpzIM8CMTTwfW
kQ3hgCjBUOluh68V/o23KuEU/5RWfeX7A7b/TX6eg5jkJ+HDk4DOcq/Qhc342fFK9cGq3RtBEYPv
r5t9U+qUhikh2WdGtgwtNSc1JYPKvqUCcdcb2ZdPimYfKt5AY12COpsjAS0irJkqQ+Z2ZBRjdu9i
BY641kvFbkLRJjWotjTsv4x6gYj4BGOgeNkfDqucF/f5YuDIUxPFF8z/cpxnmJfGMGca6FIx8IKh
mxn67e1iROH9tYLtBA/A+XqZqZ9jYjZsk9fY6SUWYkTAuFTCelPhBLqQRspjALsddhYCr8Ay4IKv
Px0W05nXevsuCmxalzvuF3OAZjdaukbY9yqmtpyOtGioiOdvsocbmyJC//6HXohPSsYRsCSyZSLq
Jceg2g3W8qa79RExuHQfHJA2c9IhhIptbkXzxbevVf3DDPcFB2lj87A+koGHKpB3vp8PvNI3ZTfu
KGMGZbT929uYCJTX0n9gPxgHb7J5/C4I73YH8Je9HxbSFyB1c9m6ipfKsU36VfnJNQrk5jYTLkrC
3N3SzNz8zgQOv2LVinBFoKVw85PTOw8EUMswIhH0qTeqcIifX1gZ+KVlRbWXj+zC0950DAVc1CI+
ei50Ord2VJ+cH0Qory6yn+r5ptnEj2H9aqTZHHaV3gOSfJMOhRHG0RRb0g2erQoYUuFOdNjOEPP6
+T+t2BGke0wzd757Ox3SorntNtqWWGTI5SII/P/tSlDGKK78/vKCQL5mkAEziZr9OYwVELYT/GzY
E5qMUMew9sLJL1DWC9atqffoXFl1PFLbbyKtfDxnwPkqE140b6wz7soA0B9qmGhbIdYFkS0WWJn/
XtXgm3fR3k6OCm2MGnq0IYyfJl9GAYM3hq5LnFhJJ9YfE8Mpze7cNufwC+k7urYNAtig8enwchpp
dcxKHe/G7hWWi6fhE23QPq9EudbSWVU4Ntoka9eTzrJQhNQ53Vu5VSMn+beMGwZ6sFghVoB9M5AQ
8I/JixnmITREiJbI69qhidMOMCPHtmhelePXgQQ4hPnHDj28BhhgFc/SoNxUakKgly+OLD4YKewn
oR02/w0jJf/fkEDYXmQGo0iA3cPaKm1JtjeUssysbNxW2j5UDJIw65J3/JMgUtDmKl3BrsvnTaJC
chxgp89rMqDAniPdDLW7MZq+7WetMHLYPedWcVmU6lkwj0yuLk3g3X9fhSQFHjeMI5ecyxDKYPnZ
LrZdAea6lNABSl7t1UkTHQQuZKyBBEXX6L1+5HKjvH916R/4WNrzPuJhFw/yVGuCmZ9GijWgdlXe
szmJ7dOx2VgdPik/SXCBC1dy1kXJ9SG6OdzuJ1nLP0APjsvtrciDZwuN3yjJUC3GGVNa8S5/9m4f
uXin0j4eXZ6aByWYiw8+cLusrvmq4iuUy/t6QI1Q7fLbu+dhGi6SpWKpfMJ/EHQY/nJJEjDLLAnX
IOkYY4R4+Q95CMaY2rpQyelm+6MRqj2BYGrJUUc3Te08jnYBA8pZgCFSiBwJkmVjw+0gEN0weVpt
sqaMXVCC5KQjZtzeH/1HXJc7R4ont4AqVF4dazMSykHw3UjOt/EPtiLThTl4OAwUNC2hdlghnYmQ
Toqj8XX2hVCE3PsP8qfycAj1xrZtZgdaztRrJj+0VGd2CniowbiTHicsamrfBIOAdI6+oOPcpCxU
RQqSH+ZxTZeDKsTFx4AgZJLJUeJ5OJHOvEqtqB4F7I4UiHAJ/NWf+UJ6foQ1P8WZJyfSvC1zNAKm
wHeChetcnmT8LWRO3Hqqm6I4koKFZSW0xjU6PmVaGF45KkSsbMUeJHduk8DIimFIWdU5kAhrgH6o
Nl9wAgYT0r5joqNEFagd3L3X8zcmsKxglrKCttQkyTKT9/TzHBQ9dwd9B8i9bTW6vwXn5Zbh6Qig
DLFcysCVUA/ny/qp/u9VniJbuV7ZGvD+KxZyrBTkDDcUzF9TXRp7NA3ykca47pny536mWLzNOy/Z
OE5Yx0AEMw0pdQTyKDk8yZZmma252Ql6Gw4rnAm0/wnpEHBhCXHi07VfMfkHjtZ6ju2nXeO2jMmM
cZ609SpLI1aZwLkwx4GYXTWU/lyvL3YGGqcGCoFGEVYw4M8QSBTf5XiokyPInzHLWTTB+wYGuJYG
ppzBTVP9zEg3uiYRCwFpxl8obMeTVuHdIlvG5+1WxTFabONXrbX2xG5QhiAGLNdcUOvrkhIH65rp
87VyRawPrSB7+piAvF9Gaogy1PYNJ/bzt9McAczRb9ikmn24mOuKxPnL1cu6h8q7gUt9ay96f5/h
Uxepk5i7LBLy5/6H3/E6u6S8NOd16t+i4Gtsu123Bj6DV0VECC/5NdadXF1IJ4LIvwAmtJ5S29xn
D+BnW35Oa80e8gyq05lwKuUfFeBeHKXW6XtyPhFzJUP43SyfU79ZQD7vmSzLVlpA/AUxnLNGZ016
FKw0j8w0h+Xo4U0OV0I9T/kdhzOwhrtTt/jaN9cqUy3MiSqpRHaAKeF+Vwxxz3b/TT0g9f/K/liu
GDuQW1vrEl987swRtHepbqIY3kg/QqlW9IQZIrXCv9jvMZYWVdth6xORHzLInb97h/pMoPkzJcf9
eAGyjadXpu06//lGC3+7/bH7y0XZuafh/IBIurEpxwafnH+WDKMDKFRjNJq24aS9rZaw5vLnkN6t
RP63ZKhS5zg2bRT1Aisg64JT5pjQu1ICewyut2eq34gvLOJE8J8RaZkS/drv7ANAjrR/w5ehIgkc
yuHa3rmbxZzNeoQj2fM95wW6q29kPoqEe9oYapEZxrxFNB22WP19C442+y5Fhdu63Z+QnWWstAvr
yPBULU/1jiLahrC6eG7CsLX8+/y9oyAbO2RabhLzHFhfDkzGel904i9epxSOm99w+g9NgsOR6x4j
7+X8ZtifAmtf57BsRIs4vcJ/8iROOUBpzgxlCPH+sYK0tnPe9uAodYpAK+HbpnusGm1GocPDHd6P
YRCad4FKtBV/rZf3J6w5km2jq4M6pxrOCKr7yVplXBelMpvqXcdz5nYW1Nup4pvtlZl/rm69zbfr
7mKAGKBs46wHsxPRZOAYrpFzAZitwAHbpKj/Y0hU5nEVmimkYe/rXpm23GQocWuSUzLIQuTqJndc
pmj+dd7uWWcwebyK4AQEakf74OE1IIGjD6vRcI2prrruS7nYhCfbCZdkJ3VmBO98w9qOn2ww1dHK
24y95zBvkoisctN9cXAmGe/OhAGRGs5k6yaaDSJtRxihFZDlYHm1p6YT82nxATm6njgZ0McxJ4Iw
ojsk6S/iK4WfcSoahjGjeAPpvsvrpdO43NRbxJYezH4dJySd3Q/PgEVtDjgmIW5ZzNmP5zYV5vsW
NhNusw+walQFH16edB5ecanCDb4V0x4kNJOSjYc8Os9cw5IOET3g9aOZ3JLW5/+oAJtxBl6Njpy4
YvUEct8HZpfNCan+/zLcuoT8TtGeAOoH5F3urdOWW9FD5Ho92osXOhMc5CIS6ttb9nA0pq9hK4vF
nuyOt66lsNfOJJACN2C0jACQNzbIthrr09QlsWYCvSdjHaE6IWbggv1/ktAnhIs0uRN2Pr9VDKZu
HQV/hcHfkj+szF1e8Kjd0FdEJ07fawB3xrXGAiHHYz9X5pYdrdbxw+cV/DW88USKJFzBJr8FII24
HzYQ2FGeoNF3wiKq6WDui+fDaS80JlZmU52/JTQRnPAPXzUBP8W0+gsizpyPRlJ3NpT1gmG7mYlb
mNw3pJSxpMA14whTMHs4I+Q7/1jqmQzUWJXLqcRSoeno6NhS3VGS+IeFCGDrVO4uUJQ3uWQUmZMa
SRBg3IUdgsyq5MWV35HM19/gWC+UV0bNYjlEwJ9910H4JIvJqC8MkogT4dZ7jJpaRy1nsjXeYywd
FER4A5eXGrE7Q/CWP3UZAfKAUJmceq9x5KrgRlNIWQu4vWAZOOP+k3y6mAOLeJhWAckKU1Oqapl/
62nEd6x8z9exRqpWGHcMQ08m/xjsExhXhr/wZZ+DmfJyuq8gMLz8yYm8n3EC6orKVuSN8GZPc6T8
auwQWb0OnLKb5NyA36lVuKnHMaq7z2+RX/oUmI0YKxDHsodyHF8P6WTdbwsjc4wmrSeK/02d7fqT
PsuYgST5s9X9bQg/liRyFxr5kxRf4GLSbBD8lwW2gxFarMgGz4QEcTrcWSYyruw7VfHkeGcT+rYn
b4KGQg5EkF4B74uKrhbazLC+Xv1dvJH2HAKrLDe6tnQM6GfJLwup5UTsXfp+fe6+OFsKNnByo19h
qGC9rigKlTJlKvTvLPXnBYx50YgFwb8/lLHL5aq5QqGLpYGk9ND8Wdp73jCPhq2o1nWUZbLCDUL8
mBT97g8to7QBYnhM7rMHV1Z0C0GJnTrveWhlH+T6Ifsa8MR+NvC4xhP0I9242aeiSnFgbsXTjEbi
twhYuWHPYID7zPnexHj4lXEbr1Gi7pn6I5fabrUNlKXTnSgXGhiuWhUyDWkSbWCrS2Lslww1CzWZ
tbtDd9oJLcwMxAwQIPSXWame9uokH8jEYfnARSWuXDEUx15kG43b2O4WkDkxn0nDuycEkm7UBeb2
51XsOtL25GQSwUPNdnaZ3bfE7J6c0dUr0j/6TNYE9qoDKyUUrkTEre+aJpUAgDJg33+daunKQRTz
aqCtswhfe80SVP5yIiFVKSngeRHa1kl9hdnc1egfXAPCfOTJWKFZxnIRhUJdVXB/5jJQekSMnZyk
w7npKdmBCA9vJ65RYQZF39APGb3wJ22kDfq7Lt1swHVVhMKcW/Qbos85F8CTnlcM7tp3YYH4gfrj
2EPF7FIdLxYZUL4bnmfLXSD0bhuZaqchS4rCKab2IN/4SyZFiLaGe249pe4l4pLJd+Ke5fNIpNex
X9yJu4uUpurLmqLy51sbnW1k05MWku/SEX3wN/mB/5Ip/VQ6gUCxCKdVlt7+bGPdHgLIh4jJX2Ah
v/HwMEKfrAHCjdfZKdfA7i8wiwgT0yMKxrml/+XUkXlSDVgEK2nv4FUsbOmU/bN3yIFd7QOJwjUt
A43Js6rRCUgY8nAP11Y8Ixl+jXjkWsi9R3uLZ7GlYdXRoXPg5uBdVeGdpC4rqlcqZFGAWwP2PvPO
i4AaWzlnFPmudZKtY8yWN5xEaWQBw7gx29uE/mx69jlykLRd9GFCISmV/lVMnO2VihFT1oTowGWJ
6jfe157IvTp/8+tv+Ch7K8d9n89C/wjcicWsrmuDsTVhRzcPvgCgUjWSbd75SENWX+OcgdaQbPGe
FcSSTHeUVZnR8U8qB0inKllZwAQ+vDTZqb3Jv/N9IL+Abl6OQEgI/gv+LewGSwXKmSFqkjp8Bnof
C/01fVZIhG/KTLL65It9xDyU3I84hSHvWv5i1yBkk+josQCizfAC8x51uweJ3V9rO9Z6JEsGQ0VK
jY6mmqHlF3ZMW05fQqrxkrzgL7U8sk5/9u5d02Bnr83zdbiaJgeqRz8TUYDbO7X67Y9JGuxBzs3T
LWwfoU9goIg+06AIlieBC7dJG92FQHfTTnla448AKm57KzrPhMP+N4o7cWslGyGwzlM4AP1Gob0a
zlBkvECmzNY6OQ5mO/7uk7+QSebLLGhIFtaYIk34WHRdMCpjRb616bFm4HSDDCXA1dFLoBt2jNjd
eJFhFIbh3//oQ0I8MfapyZIXm9phAvJUE+9oXtjaVdqm+tqvRtbb7DA8zJXPnZpG/05wdLEaeZkt
4mNhRMeI7xIVOaOd3SI2pDf43n8XZl/jD9p3G+PfOUMSwV7AjIJ6yKs6D5WkPpxRjuwtg3lISqB/
ByGBcCCvwqE/kxlafEkcEsM+ZGNsKEbT0ClIbOX0NEPO4rLg5jomgtVpQ7neJu+x/qAsKZ637fW5
JrVZvES3/6C+HndVz5R+CpdxkHKf5AWetHLij0TfL1Zzk2wiR2SDIykD2etdvhoyxbEEDlFHr0c5
LrFl/jVjDoOkBL+tsUBKd8bem3Re9+MTzx0+mu2Xk37nlvrFYwuXNQmQ4yFXzoMybOjZBKXlrW+F
uPVmZdxn1fC/vXgxH/QtAhBfKfN/1NyDjydTcmAZnrmqx3M2mvhUkv2KU046y2gTGFSe679r+6A3
4/ZBPyvNqxvrqginFiM4M3uz8wuEdy+l0alyUMRD1zH7nuBDVjqoMO4SQ+bHtXcrfjWoP26kkibO
2cBguxbyToAqX6egz8QMfqlrCOpyeCTSUsvOOjx83UKNPGpxb6QY/gRh0IjWQkXXwhGDlRy7+Q26
Cs171o17ETSvvl+52B20F19RLix8jEBLhVsqIUjDH5jwJgrET/PekbXRrVv+LQxQasPQS5qFv9Nt
flSOjs/mqq22QCv9Pts9IqhE3ANabS611h0FtmZLF31K4np5jjP82nlRJZoZb66EGu7UibjEpXZd
++ee+9ayPzGmLivryCMPm7uSOczsv93cU9KpJm+TwbvVrERTE84lqo+IlNTxMLwfFNBPQGFfxW5L
zN1T6szE/DHLsvZc9v3l+VWimwETMwlZBhi9bgBjm11HOS/mOHN8kQgaJwhLzLm0SONP/wmisiPp
hBnNh/vQciKmVhZOFsb7LyRucSVLuYH35zcm9tPNomlFLI7x9wrIigWU1sFeDhsPfSDCQH1p5V42
X4VBvIdp1KfMunTlRDovRnxWw5wqm3NIWq+TTuPL0oqBGdOeTQDAPvtA7LGGv1B/mrxwGO02e4RW
i16YGGap/u0ZpfdGnQ9jBmy9VuvVCZDhN29d8OwmbFsBc/y+55mKh1G7ClFCz7kKvHNXsVNloE5S
JgggtupdPQJUQ5+SKuBvT6aqcilxf+CIyqg0HBbt3W2P42FhGXV7nwDGBzkHru/0KPEsIIkQ85b1
/L579tSWDE9yuzoxxmHuDAWaogD1E7nPp2MhwXKvI0j8WDi6u4PBsGq3D4wbopvI4hYw2wa8Lmc3
UCOkUjJDbFRUvHPelVWTYlTwP/bXEQjQ0EG2+nAgoxrDkHCDO2etcaXh/86GRf6BGewWmrdpq+Xz
NdCyBn589fdjzZHi+UH71zxDQpjX0/pbkZm7ZkuYUjcaYmSCtScTk648cdBVHRYZjuhYUoX5KVRy
hit29LDBNMcQXVqgv5RRl6lN5jzOQSdfXHV1RzR0CzIl9Aln3L9fi/kpQ/heW63iHiBMz4rmcgto
Aqy/4oB6Q7rrxflrBbXhN6+z7iy+t292JnMTffLCelOuxfE+g+fKLCUSUHc/BlxyaKcf037FJ2PY
7Ko6ZSQCDqT9pS/pvwYuCNRp0i7qjrw/jciwelKTgbfMR/ga3ZzJkFKMTwtrjbnXzRYLhDwfO0HE
oLl0AFF7RF979JFolaR2YO40wcZtmJySBSULQuMKTyVpXT9g8uMpQjh+5N0MAI+Pb2XfedZak5pt
4p5OpGdkGQACBhLqaHU6nR0p/ToJMHow6tc05fjNnHc5MimUYm5M7t874gDkBGNjA3PGr3RXkdQg
LTnrNR/F+A6SzzOgdmRIc/IyPGkIT+ZVfVkbuOZTvCiW0wUhNGkLbal/a5CbRtWlvkrT9HV6Q09F
lNWCq5BuS2+sPLdx/RbwRXXP+BbpNx+oC3LDDB3FZKiDoUx8YLVZXiOrOqGMM7gHul4xQbmYxI0h
tlb23wes2ICsauCyla8RFdS7Rjbugu+BTCcMppqtwFsZHLJ/zKc2pOeHiq833ybMKT/eBeeMKMJe
XvdKWhVoVK8LUAGMC7ejFoJOF90oWF8K9VNRw05X01bW9LyBZb+TbpVucuuSA+q42iOv5oQNO7pX
cUC/oYods9XC4ov0K2CK5B6zYyk3OqrV9n3R6XOR5pcf/7vUonYTzeu1aj1z2nB0VKzkm8gvt8ma
utLJLCagKaXX10X/LI/sxDFaIx2cEhaSPKUiOAV4FkvYvebEvP9sa+TR73IhL4waNL093dPqHNJo
gmKKIxm2EKa/Vku34An3unua4Z2g+9i/+BJ0U+9zshQDfhbvNn4ze6O0sNTeQQOJ4o1KD7EgeORo
/EHYmCRQAvYHnJBIJsIlaYzNzV98FlImmkV9a+rNIIlpilelX4KHJgFCzdgJFiNTn9KltM4z0U5i
ydPu0U3vAy7dxEjvS6raUePsqpp48ALP/r4pxFdxOGceUVGjq6rmYQYtAoKWPhydDI0AAuDyby6Y
zvNisY0eSR5pPxpgaz5d0BtNnO76SgaAEM3bGASuXcakqar2Z8ETCtuJmoMWObbcT7A+wJGYPh9V
4HvCj4yDwhqt0CPwQyMBvyyXEdfPTjfhJkKo0xc+NafUiflKLeRKgdc++AaA6ZlQs2z8pdxY7NoN
1r3tTQ/R+YVQ6FmGzyJNAUfNrv8JBAhze1FBS5AQq7AbhDWXzX7l87LwfXvCur81LT4xFIwv63J7
3PDfI8m61Zo5GV+ZqJqgzKa6UMkGA23SIY3eblLl6jKm6EehWmU5YX65+elZJBw3Rz64C7EM0dEZ
/36F22zDEem8D3joCQnpon8R4ZEIx1X6iGmKdoCxnktFBTLq2BaR9iNylzNKTUAl5lnhSnYg2kLo
WHXIKLqksR+m5l9rXZkeM/P5kNTUvgv43XH/VkUETVNweJoHF98vErceAxDW+9Wk4j4HL67Zhtgb
KQxHHIaeKArj7mmtVLyyNymlcWCYyntZX+az3J5B40ztLq5rpiWZIw2MW1BBU8MStQYgHVabxSpa
WKfiyyW4fGLJ5NSKaHkZu+gRhIOa+7GQA8EG0sMpmIgoKQRNd/Lx4ekF2/8l6j9d4M9hNdIRdDJl
6+uITd79EaeEpf1fFAUFyMpo4eeSbqgP6n4n+LNtk8sprpzg3vk0zGtdQ0etd0BZCWxmsDiiIUKG
wyxn8Erde6qof7SwM+fJkRca7SmounXApKlEMPd+o1J0ZN1Iz06ML8lNx8c/EuyYmBlVU1digc1M
WJ//sA96jBZr3F7kRnjzGtPjmIbvy95kFMQhHwtp1ytDp1lVRlqO5C0RY57WP8SPJ7Dsmf1tyevz
p5KMyPimpXw7hTl6R3tqPZWB2R9kScHrx2ZJ1haZxGhSRykacjV0EvjvjLcF0SAq0X5V1fhu6cvn
MyZ2Nibv2WhVytUXNaQP72DzJqEaS57SOb+38+li04tiwxQS5WZCiGAW55el+KgCsq/N5qrt2Vif
Dkiv980LyQQXy0t6be2JeA8tfOw86rMYPTxesGZ2CJgOEZgb6WBtgUcSP99OyYE+jEXG3245or61
mDNXpShJO8HlZdiUywiGaODrPCCMm8Sn1bvwKzbgMdRgYRh77MvZ/07/gkmSUa5Rnahb8L+HEARX
fmPrdip83KSGLA+N5SJW6efEdR20/Y5Tis9bGAzJkdLnhYdrih50YHBoIaYDeK/yx7sPp0Db4cgh
013ARUAmt+9HEytAP/WacE77YRZV5lx78zaX6H/18JNoq9kUlbHdawkviRNj4o7RBzcAqnS/ATjV
RNU7SJ9SqZlSBQMTZhWkWwXK3m09gfvgxW3Xb2i9OmeyyZR+SGJBy3bhyAm0R7nTCE5pTD5LnLUa
2V4V9/BO8ySzWUeE/FMliqoGZJofD2vItsboCUaOn++GpXWH4cmqA/htVvY+/aT5fuvsWHoTtfFs
DA7JtoFxOitW9iYJqHUhZP3SiZ0ahC4Wwv43QazTy7t0I02C3j08hIGcTzzTdC1AMYHeGAhwwfTm
1iMaNJCV4rT5Kz8nmgEtI/4OsClgnoc9Ncbkv9kNXf24UO7P1wHKOvPRisTGsv8puWe71fb4dYbA
w6n92lRTLbHF1OU9Zjhsh9wXyxDTfR6DUZPqANg8N0TXQAgQosOEPJi5aQIUCJIYrBKwJAt/T/4O
MOF5oIdNF+szxuyDYvlaH/ltbkCteRZXo2rDS8yn+EthENkVCGrsPoiSSCXTqoDRSxXMBFLQVVQq
uQ2yOx4DnBQ53YXYDnB9iTQDa+tMwn+8ywvFTmNtc067WpeAZGHu4zyRYGQYV78Ebcajlfmceooc
MQ2Av2gbN1mfJeeIkCZDbUVcUPwtMALOl9FDGk/pmHk1BE7YrEuaoO0V1lijov2PYNhVQBFJjWMq
FBhFE4e4D+UZGJ7LDRXP6Alfgk562zwQ9iXJr0PQ5O7k9HLKRpef8MCBUk0/Uht7Hx3f1Fv7J75e
TGLuiZFhAeNXFuvj5erBePAQ9iSthEFEWrMjf5T7sp/YZK5F/FDhhE5WRy2S06CSGD6R9JEeC5WD
0LFEcU7qjgGdKI7VtWNpV7ruN02tD50i3WiFub7C9HwLwin32q03pzbMgIg3Z2H9J8ny1qCRd3YI
9CzCSDE3/lHL5Ge4URP7y8Gb8i4JL0AYxLH/0bVFf3ov4XX+G6JVxUYeVyZbSz894Pu8S85zorDo
62etAD+ynXKsY/k/wS47Ku9kq3btHCyI5StKA4U4FasUNGQKyT/j9vsTMNdh/IAeC00cEwj3sqZV
xom2aEcXNTrMz2XXQSFH5eFnrCr2myLLZVQQOXHSPVJG4kSJl2d50IwA09q8XyAzIMe06Dp+9N3s
lqBP7GJjQaO6K9uMiOSxo5cv/VsDFsxavAlaVPd4LQLcg43lv0//6uXJMcecGgokacv7+ul548y2
zKKG5EgLvFOFwNFmOvCk49X0AEbiTEbakkKTb2hc9jE2pxqpFgERxreXxLAjCNX4uwixJVeO3YmG
446uOrpqvkgo1JY2NIYRhkn9RBasbtWdef6ujqabzM4gOB8aAq81sDvwWFghwpzhl33HPa2ZFrJR
HJVXyvWw3NUefz2zS8NmXifmnFuhgNUfPV4RDk+2IVThhznVfYMVqc1/JBRvgVscbBOg5uz2rXV3
mk5RoQhm3zxQSrRxpybOHdsIdbZ83TalQ8YQkF+ohsKDQtRMVQtsKQlv6JdAhd382cAGMh4ZNGqm
mBldRCuZkUJ54P1iWcBmQ5px0UMm86C0UXXZBG9K7jDSVT6wyFj3iOIJ6kkVNGoxaCCgr1BwlJbf
8Bhkpm+GYWG7+aW2MOG8ST5eaclzyYN78ODE6XKI1F1ExNMC876g4TKo/Y7GKlpheyPKUMQtk2pf
ZVMHJsTEJahvYXYBC8mGS8xmVeg/JsXatQYS5p+vzuN8SnlFaPS9tyESUwP/H8Uax8zuQ2Iz3tL/
H/0HFdTOZVxA82Orhtz9SOJhg8of1KIKAJUsT8xeqEvLCZsjKmapzwAfirSLT2v4hre9cBvpZovI
Wd/RxDASoj+FohegMDzPA9d7YbrbHxwQMLN5FxGMfyRpqXPooQNflkdYt6mAwa1wa8/QVncTQKtA
kAWk77hegIqnkfO5o5fHQk2Jci7YHuXPSWrJpDxfgdddkOK1i6X+2sW32l3jOVV9DYv2Wd0cPcRE
Ec/45LLsdj54ySNBe0rQDYfEJBGKegDStK0sbryVZWZ//1RdIVO3yYNrLMk0wdXz7Y0DOvZMLrcr
8Th/PLBhemTQGYXIRVQLTfeMZSG3LsdAuw6sNgwqbE69OYWdNsydQkx0lx9hT7hyVMdRKpRb5gc9
T6NWrgQPzLCMGP5rorkW2hgJ9LjasmfVjZOq39mkIfZxeRDObwdxBNGjwgZB2/W5FmGucAUrdm37
QYyRqeDpusw2x2iK8KGbsXoa9iO6++bLSonVoN9OcVclJYk2sbvgeH1Dqw3O7Tt6hgvKFTHhwg2/
4sQYnZ+nlQaegBHtMsicN8Y2rBWcZl9BiCTpQoCtj8jt3uFnF/M+Lj7DhJ4O48hI4gKBoF3XjNsn
Vgf0YSNW1C1Z86QWHKxyKFTUy2/VX8gXgQAF4ebPa+PQvfklSg+IueEut+oz5pum57d5ZKycsvOZ
sZhBnKoy1JOFdRTQtXzT8zuVBsyU7zDhungn1Gkv1Eu4k5IEyK5v/8sEcJOGuSskFGeIoqXXEPBs
Dr1nZEOCEixWO0Xjqz2bnh6RoVnRixjSxF+6jPBq0+UWyXAB1J8zGEJf+CZ1odaEuJNQzVKfRkzH
shjgA/1NNlnRlV6pOnoXncmf7cenwsbnfgIvH8xCqiA14AhfGx4Gu0tFCHJsy++X55GWDUVXwin/
G0sTBzMrlG+Hddb/8iaE5fWWDl7cw1Ml202d7ik701BAU4OUzuZaGTtumpsj4pbqnCfUk15HhKjr
0wvagjn7QUuX8XxyvbZK15M4LxfQ8H6DKE5FIGm2KOm07BYAi6sRwTRdA0syRPNnTbJmwcUxnVRZ
hQ2RSOQNrEgNZPAOj+78hnN0bslFymY+gD56gOkrWwJpftnlVnqLK+Vu5Sj5ysD3Pbfvdm4xtRkv
fV5sx2hQRYDEg7RPRI2MgZH1ZgQ6SyiPHH2kwycOGK7HL93uOwyGlYh1icGmPAPidMYp9/XW0Ajn
l4H0MTl93vGQ3OgFJ6M/iDiCm1QBxuhfsqXpdVChjC9KgRNS7oqYI4VVq+eZxZN8Gz3pbv38JRwo
pPKaJV9Zl/wDhhkbcN4+v6OttsxXePbR7O/antj4cdrSvpmlGseXWG7g2lObepFsydgCFgGBvQ3r
SCUjp3s2ru/DWCeB7ZBKZIHdD2Ly002X2FMCTomryUbThbgUDIp54l5hFGBCC22TCHzLq3fJyS3k
fDKLnu15B4D9/GsGkHnQ384RzfTc9FN4Rr3PjT3RVC2F2ndyjeG8CRJGAXnEijhV1rdiKqwsxype
yNJIUe3YD7Z5Il0pBuetbHEi18pHkPpZcyZdaTZtA+uW6jaxYGkMrdDoc6kv7NmCph6rwhsf7cCb
cuwscG4tRJ6bL5l+6hFhLhJtn4xi2RhPBQdSM7vBfUDi398CFECOkx0KN7tuUcgNSvwuFniW4rTV
8lbTUbP29yZZW66g6q2b8YTnXfa0D1PC6M1OHR41jcSjrvzcFKaVBCY/MzoWZ0i4eXO63w9ABj06
BARwYQsdeaBjBZJXnpnzpJuTehUIJBO903fq5aYTIvvZQp8lje6PFd13QC3SeWIwEkHGqese8uY/
lECcqypyE1al5TixWXRy0H7RYq9jTEXOCpZLBXMRTexFy3/Yyna39FDvRevq0ZHZcwN6zm/wqJFR
1/Tdt00L9vLF0/cijhf0ng/QgNngEJB3MIS/Se6vYZR7PEcPw5/Mmu4nKM0hfqx8zzcWAfS/tF06
+KQwUN9QE42UA9wbMdBseB3EHV+pch8NOuNIv+VXPXxd4cC1/DLsP1fIuzLCG9TbtWNFeHWFxLf9
i9ads7LOMV2cmB91QdqJPdtxu3+GmTu+KITrVmmDbim8D12WrGwLBr46NTj283hojz6piIo0yZri
khtcuOeoOq1U476BBBFPRSGoA1ACFTnmiDjBw0+K2zLxgyqpKw7wVWjPtdOQsBCqb9saeNNvlRvD
Y5H5wk5ImDJKYCbtHETFCMlAQdaOCi7ceYaTQnkvQLztDFye1QPPHaOUQ7JwW8C5CU4r63guXlwT
Cm47WH5tFbKkuwXP1MIvWLi3BPrNwZI2SglXRCCG9jM5z9aprmUUfECEjvGshBqSIFE1SflUrvvn
LgjcECxTfggc+jKbSoMRcMZgtRmckCv+vvd4kOMI6KpmgvzTa11y69cm8ZyrSSKt2xQZa1myM3eJ
j9AG6Pt6twpFCkXeKbRzYpntA69Q2jvfK6M0C5j5PEqL/3yzUZ/wNyWJEtCD0MePutj5mz0pLZ/M
b6vZqjCNRl2/DQnJdCm0iQfVmi6DRYLgi7p4u5XOV4qB6j9wV2HERXvkSMEktMPCTxm+RyJd8Hpe
IUqbeu0OBRAe+K4xpquJjYj7pSMNoWBOMTNDjHSwJXjLiTtH5uuNyMiYzWdtMaiOLMN/8GxdFVG9
a4YqJdlydQCXryvCE4E2B7TPpZ0wCjwpSHB7+6hC2AGLL+MBujixFvHvQPa6N6RsbHF7YEqh5F9v
4M+61D3mntO+NWe1MH8ovLF7bluVduR1K1I/CpXKwjYaSR12BnifWX1JNITypWzR2f/2ALVYxn7X
F+Jb8M3RuCb8gP/WFwcXOiesEbiuZw4YYcN3a59P2uuS+YkQjyiJXq0zTQKOwIYLq105mnJ/zzXP
EtYl54lrLamEVqa0YOIyPF3E79IgfX+RYfmHtUU1JOpYsfy2sxgn//u9WEVOaojgLPTxKqit13QF
kr+WJj82b0Wv6mfyHFOpejinRhNFJ0vLYGbQ46C8y9SggfDjr17D9OJeauuwiVewd4gtY4Rzgrf9
jAQOkGMz4jayrl4Rx2OWP/Cr+1L8El/neEra1uajiArulV/lnQnHK5wr/W8Huwgjt05S2us0s5dn
Kj4KPpnN+08C3/wednpKnTYau+fnab7+1TK9qribEsaVdkoBhfh3bUadb3UO9432pUv5M60pCPRI
O5Rpjsfn4iiXW9LSm0gY1LJPwIkA6rcfutLZJUdy32p+Kpb4HCoIfl/wlkm6X3IuAcx86oG15kL5
J0oSAOSxN3QEJJQ0zW/BC4E2qrTC8SgZXUSwxX4BHcrLqvyAZPa4rzYB4owKmEXA/NPCGOXdaxze
SV0iiG3slorHUK1KXVjBPgUBnPc/mZgnqFPogfFQFBlvukWUw3IH626oQFYLp/gX2vWabJ/xM447
Lhie4yOX5ADDc3Zl02xIqY9oEkIPiVE6iJKaybOe087benLMe+ey5sGYe2krW0EqxEj7i865HH+x
m2t20N4AtPTqlKmuFScag54b7FAabDV6GrR0CVApBNDSToMsEu0+TDMp7sJghWIKAwKDsDXT6M6i
86KRDNA2jBZnIDWvUgaJVf4Gr1Kw6rW0E6oEQawgf4KLz7QGdfkob5bSaFcFlQfzmFBu/olK0vUQ
b2PekOHD1UmJsgKt6R43tjhfkJ+jcKrMEL2zL+M4efC3RnZQL4ad3GLmrE2UVpo9GB+c7LfUd6yC
CHldsQGEs9LOGmTddVJy5XCmOBxyOyUv51GFw2Ee0v3o7sfdrkNKiMNbYzvgKACJLjFqZnMRocTg
/2e1k4P+M9BJJLQ/SINUQgpxdUNMIwQxDg77kckhLdU+KIzyUU+2Jz0ahA++uehKqqCx/1BAktwC
kNgDhBzDKtlhB5A/PRH5kWdrDRCIPdtiEU1z1bg82u9R05+SNuBcbRWOFZYJWyiHFhi7f5zv8hMn
dZirpMfkbQFOqYUWpXE9kPRrcpQ5CAmj3w/yVpmr9zsg77FIMmmyp+Xk91Z5emDtVSmb3Eu3Q9Yr
MLtS2yxRec9CgQEXtwpYT07kahLS76Q1iHSK8kl+yv3ZFqJhjwzzOXtODNU9PtejMIyOTYHsFY/N
aEj1txjHS0OyU8j3KEHBZenBDc9y1BXxTk9WGpve4d+hptNOYsJ9H5zw5WjYJJGFxEOpbEVZnflO
D2A1MbKaF+IpciVJ5zfdGSLraNtsOoel1sglhAyViHKH6oJf2jxK56hBZABqes2ydSALQAyHCOMz
sRAVVIRyNp6gfVH4H9D7lDKbSEPkob1u83etmbk61Mlj3lZzbTXf1M2T87EVYdgC4WADNWO/A5P+
PbmcmXR0IN5wctuLvaP8C2fn4jnKgH/VSOpSFiNP1qBowgd+J9WlunMLboXYnt5BYNlzMwNrU7IF
FFWF54jILNbUisHYsDgXqY001yVKfJe+DPDe74Bp9Aje/zdnhed7a/q+1QiIqUCr03M6U8R97V0T
7ddPPLpJuhN6F8ZSLDjS761fOs671ThJ4Ttg+2biy3BQGXz5kCqtfv26XXnnG/jDdMjmyUN7HYOi
j1kpLT4ey2hJNEBGTuS/WKihqaYnOoYs9ArM/WKmEbi6I4AZkCqjFnQKOE+w10kqbYneN5dkzPbs
ZJ5RPA0Di1FnXsoG4zdfiXEasAxTpVDe7OACYLY0JMXRmS5yDLIu1cnY8ue4MChT6TCkF4j+dmtN
O6YGTcO3ld10+bYJcWvA0BcVQ5AssszVzJFX9ouy2XwMa6mwSx+sq6AVMoy+0CIzZN8AOh1MJfwU
t8iuaoKtrNFUR01QJ6dGgGBXgx28GM2bQmxXuNKwbM+PewG50T0N/0uSBv0kkhJXc99eX8RehuYx
sX4reY4FJ/kAwvQ/IZwbEbqUkm2jFDaQ6u7igOB8JBX3TGZwiMT86acBp7vOLleh0yjFHDhu9RnN
yCitc5VzLdnfPUNGA/3Da9U6BAb4KsbncHdGeumH97YyuS/vINf9TmTcktlmJGuVHhVYGF5/qssl
fUWuR5ss0Aa+RtApha0xMsY1XLYmdgAyhord2u5oZ3unYRD5fT+2w4AEJgZV30JU8w31q86Dybc7
U2NivmDX5CCmfdGICH9WNbXbH5vu3mYJZZUhqxZArhrs2YPyrKhiJ5fllj8fpXfDEOTG+uKlHbFN
hiPeTzehyE3RRzD/k1HkqOwBQR3vGCrXfgnidNcI8UXO4ZHe4l93Dtfd+PJEPJmL4pifMlUaxlX0
9sfbQLIsHlZ/lYyXzVVDSlhLe6eDoXfsWY8A+/UwONV0YligSSnahxNVd9lr8lD3lpAnUkcoXSgO
k6o3UWjK2Z+iOKkYWhGAkzSlPu5KEPPAhHtcVUX+Zfxg+vVmf9ThvvKNmcDAiPbIfTqDYl7ZwU0e
+AmTiZJllFRw0paa9HlGjhpctjirJPA0LMDGPVhD1GvpnLA6OZ3DMOa4IC9A5hjyIPS/xsORyV19
XGtJThpP43jTSs4CToT2hjgnrYl7VtW6zjcO5U5JAnUKfWozd2o5VehvpXtnOm0+XBmv46e0NfsW
sd1dxsMxU8x4pswxUgcvUzZJQpybYJ07IjC5BGuYG08hsw4hffck5HNoUhb3T3Js4AehHFzrj4LC
6v78wpT26HF6L9180L9B84xy5/Nn2fYlqlEF6B5T9ARr47uD1VfjdhXAUyT09zpmlQYxwpVKVSTl
Ie2Np6C6ALAisQkwITh4FyF79vSCZ76KteCHlbqGc6U4WyIb9ZRAeU/QQY+YK2EPx8h0hDKGwx/e
IinT1h7uu4BuD21hwqS02FRcyTvJU9Ma/Hs1BfX21tfEOUl9ELSxIy6xTyAxNkFBwgaZT8y9Qe/Y
yUH1IdOJd9qa7IowKeqtYwcTOeWaVQkCC/lxpCHUekRAlpLMh70VE4cFbQXVz28a75G9m9n40iXh
+r5NyoZPUADba8Dz/RHD3q/Y9oDQABReFlHZ7u/+idTCxcPPIq5zeXR140vOs6Q9A33zWNroKmGO
CNfEJ1q2kEaOJnzUArchLLTgLjBtUWxPVuKsb1aSz2JTKWh1vIiQJJICkD+VgcH9Fq7VKOn6WQy1
pVXQEvVz94meA2R7bpCQhyQfM3hlAmL0fuE0xZAtuwGL2C+9eeQWf6TZCi+btpS/7gdX/9VAFLXP
8iAHuBg4S5f2jErhuSZOJOeYAW5+4ohEMdeuexKHRSoBQLNrCgbEX5igGvqVdtCtgFho+MagzRuS
LpURczwfSIf+kXkRfePqnQvZOhZAyki7/dLN4HdWd3+4ifwA4DNK8q0nxBaQx0N3FLkDidsoDXpv
3PrNAXwJGdMOxUpNAqRL10AtS8Y2HlQ0tA1n3FqQqoyARwghUE1dqkDW9GrcHBHgGkiwcVK/wu6O
OYnmLNdd6nh1O4oAowiBhywD33jp6dGlBi1L0iinOeDwrr5CCj2WY3Z6931wxdr9M8dFGYl/6Afd
f519pca0a54IgIE08XBsjtZL7wJ7ipB/mT/vndcjucEkYa9SyOfNKix002gYzuD7BJwD2HUKzOQ7
WhRrhseVFR1CFJYFWqqRdYq2OQQxfyY5IHQku0hv2Kp82eZH3Hl4/SscHXa4XJE8vUeakbGwCBES
QYjAvTNOv1jqV5Hc/vw5aQ2hFjO8525Z6f2Ety77/39orhNJxcC8j1tciG26FuTGPhtxZcQXM7B7
Ed4+/Zkwam/G3Rh336TGZsUj2Ym9688E8YSC7c1TIMs63ej3hHbEjlnvJ7qW0nSS2m4G/8SRvBSu
JjlCvXqZKnILiPS4MLCU0GOh4O0QgAZ/br7mWb+cUrWDedfbiLCAPlrSuy2m6ZsR60lzMLTEUJlm
oI4/k8HiGv01f7UOiCaKv4/8pp6BrsUPJ4Y1dghe+9pMsRLvkX2O8zPPQMw4sEv8uLOHio6o8teh
/7MbYs3AYQ7fzXrvY6sHRm7b825zyjtG9Ps5Jm5LZRG/sx7UDVhHbpUtcAi/KbxD+vMbrszyDfYf
51Djf7tY/6pGIoib5vw8lii1VGQrrOIYQY4E3rfG5TvZhAQfmbl0BhX+KsaUuikM+ZXok9Q0OIAy
A0BquAH+FQCfM30ni3lNLiNZaGxqEVxfrwEokQf50TlQSVhfXyOKAyj+6s4kpt9c/N6tZg9MO/mE
w9UcB4zFG6Xbrl3ocx27+ONrYPTvgKZa0NWM6uEp6ni+Gik+HM6QS0GXOTKrLYNJujCdK6mkoHZi
f3AdsJd8Q/iv3AywtQW8x+OQWFlRbJhhpWZiHjnXBkvZ+F8oXE4orCLCrbQDgejhpRcVwU2jV4eY
7+idWV/AKxUK++rJ/bRXxdkiiNFWSM9bMfQ/OW0OxaGr9XGVh45a3Q48XrQ4a2ApuQEIpqV1y1tk
V+XMhU4+esPSj5nDmhU6+dFZkvPAeEONaEJO4bvam+p7Fo2nziLBWIRc2r0RsdwjFo5/Ik08qFpH
n87F7iM3so54QSP74lO71rHsAgWeo/OQGRO6S+P+3YmZQT8/LFIzz3xt50Q28fmLSKZyGoea3Lxk
iyTQBCBS1oe0jMHNxTbCtaj49nb+ZjUTYBvIS+0ugYt/WHb9AO1Jm74EeiGUYfM8WU/AEd4PPCpo
KJ3vxSiPgFD6NN85PbuKJcrdzLhfb24s1Vy4YzhmYaJj3etMiAChtPx95bMgSoTIOAuo2qxDcA+Z
kEY3aefVb3cZhM5w8ni/ru2ZBSWQQwwnflmucpR+rncRBoXajNawHFcxNeMW+GcPk2V4gbHSeDQs
m/BsS0fMkUyA9Yp6Vj6KhwynTYAMPzO+wMsbt8H2+PkrN26yhwrqXyddl7Z+5b/WNH0gEYEbTULn
56V985wyHI7xT3SlwZoQ/whgEC6svkYo8jesVbTt3l61R79+KD2SLNHBpE7LgsNhEXzaJ36PsO1S
UQ/CCYQvM8auGQKss4biCfP06NCfHrH0qDKM7CrvwVAh60Y2kiR5+o2zFg2aaJBzfbt+se/hq8VI
hz8JzWLkrKLhGAM6LSqSeW86Z0woLwe8HN1DWi6uygGRZmkfr4uBtI1D2eEtdxSPuV3IuyF74Z2j
Y3uAPaH2FEBf0EsZQHXRnQKBh6h4AXf2N+dQSkp5BZp+HDO18GkiEjv1UYHF6QZmhH1O9TmZjQ4A
+WiTvRFqVzwE4qD1DfmL/xZLSmpSW/OWiV9U96kfXPwiLqnliAEeARi6JqzdR4bxm99MRnBR6YqF
F5wf9o4Js5DvbneKYj86bNV5ucG67cop9lQRjaCyg+sUREclUsNKxh1j8DEBpPPEAZbOKGNogzkq
2tL3wWBRUDL9cigDtNb4o60yQ+h2VPPPQIxD9PS/STM9WDOAlSEW5oOkBL2m4HEcQyTgfSSbjdIF
kXrx2GykMUCBwvowVjZfcgInfhXU0N/YZknOAom+v4bmdan17pUd3Gc91O0yAOCRWgup4ZDIA4Sh
GSwP1e2RPvsXJ1hA8FOFlgdlYFdbJ5/hAhhpGSKM3rHJUstfuAj/Xc12INeeUH/Tahwj2LqOKOm0
daEhV0zSXG38u77DT5tGbP6AwvnclKGV1B7DuSWRQyulh0ZxZ4C+qTVvG0wfDs7L1XpbtlKCQ36Y
NJS8CRbXfJpObhz7RHRT0XfhxFXGGiaShDPO9qrv74L4COZfMixbTA+69vVDdFPO21eqWCsUEh6I
AZPkRjh1N9cDoSdfgRzDN+1M9OMS1aO0ir0h+ogQdjFwFS1ll+XCzJg/G0zoBWGpJUJavOvQMfac
+mDJEz9EbT/8U3UM8LVxmub1JWvOaMYMx1R9/b7WKg1yBkUeyH9jX3w6txOkRNNKNfLRUeGCxPvN
2wGKSMzGSZF3huF1qikX4Oar/5Ecvz4+fsJiChsYgweeViDyHk4H7HJ9NjOk5l/GSASzEyudjJNx
TVDGIhF2oU6z/YDgnWLR6jY399h9Sco4rMsnS89I+JtNFC9AuZPfCrdkgkOy8o1jAbWW3XE6oc5x
ddXsJArgr9lGnngSIZlIHkfZng5x5rjLXs9/Lyp0JtBIiU9XiAScvTPfuFmufrQ4tpvmTZG432j1
LXUHvOtNvYuPSeUTa9LNhd5UXkSvbBBrWplp6wivOmrumSUuVbcSN6k/zqRjWj4uKRDL3mflXbTa
pJIxs86wLk++CDOR+p3KK4GCLumTKn/EHCG8gyaw0H47wRGPVtacVImmDFfK4G4IwJ4qQ8gLqF5j
QQMOvDAULLqP6Judk02lRmnYSrTJd+da4Zi5+XbusdVSFg7tC3t81gVt1gwcnRfI5eIsIOgYuJun
goDBfhlxyrEMH5QT7TnxiSq6STq4KCR+tErP4yoX1Xbt/CiZd/Yzen5vtYBlz24MwDEHeM7g3wkM
w/gVUgUgpo1frvk/uDomEGDVYNKxotwkvisAQyMm9GuKaDXypMQRYa7qaapQy4KzHWp4CagyMI++
cEm7HYCk89M/Dmw4rMa5SoV9HTgqvhU50CAgAmzXeXPPAtmcPctMBzm05qPcaRJtGUXtA5XDTnlX
Y9QJAZS9KTlZJ/pNDbQHD4UBPaee/ubWogYRL71o2RJ7MhuE5mrGTu4vWt2lXDWVDOoQbKzFXaQc
W0FySrwXQ9mOmTyBeT4GRXC0NoVrVyzZO8JOUhLtBtg2vkzPHBUZlPYEonE0tzkPg4aagH1sFjd5
3eKHwgbRu2Kk1FUlYY1q9xbOEf4pYVMvflStdzve/LFABLU3vxuVZ1KgKdMxKas6Ysh9Xj611r/R
W2pFjoANM/6omaFUDII1L6tcaPxXQgN01MbizFBgUE6NMPVuRl+pUZjij9szTbjEg9fL5qOncDQO
TUnip5/10PMXfDjtoPpMMLg8DS9yYUVnmHUDF56rIcgMKU7dgVXzELylotnMxZrX4Y6YLZvcY86G
5s+4XtV7vWC/p0TuoUmAC507fqvrusrVIOPCPtC3Fj+TI4mquko6r2PiyNDcn4ECLkb2fqUk2qxo
MSranY1BiIL8Rd61laJ0DOFBK0IA+q59qcfvHZTmlApUqOluS6oxx8GnYnddMZB6kLrWF5KNupMF
uGc8JJWcKzHy9WNh9JpeP5cL2Y4bqM8u+QBzaCMxtwkebaxkz6z4LJA4dTZVQO7sikj+W/gINU9b
gdPEmxRIm+TVORXvGIrxuUBntbtQxyezuFDpIFxGsRHQoOYgEVNT2U5ywRWJBeUVmSG1rfiZ1kGT
7GGQK6qmydEYW1Km7cqaRHfTzZRmEHuO2242l9G7hZ9LKJgNLGRsklDJSR2ZfZJlze2FZp9CCMdp
Tcmg+xl0/4tMwpsszIzOlpdT5r8NNbg9VcETQISNodTpb6owgnK14DcEa3qlT98drVExFl6SJUvt
Xqt4ug+Qff15iWMu7FfOk+SGmQ6V1Gn+4n01LTJte4kzFtd5KpHEr7zlJSFQr2A55afPucZR2emz
Fwvs544aOxNF/23b0Qjtf0S7rrw7AI4vhemK44A4WhyUjKT4J8lAGl2kFgqKDteaD596f7j1Ef6k
75g9jDf/RnVpfmLDDgqvBRXhvQXetKiZjVH1dwk3l3mIUCAUeYpOmcmW1KCStDiLUxKtz1S0zWPd
MnBnp4zGA3VP8vRad/7cQdQbu3j6nI/gRmg1tWC4ckTz/ekGbP7TFiPfX4lcxinfzBfz+XNdh58T
WMcuCJoLa24m8OA4ljyKNAWU6CT2VntHgNioBRUrX+zWDl8LVvU9QkHNiYKDpKVgUrJyBuXtfeuD
zeVa5Vo0LctbEAgYjdgjU1LF56vHUyqIqLArdCBtokAAcW+SeVEOMqTFmX4bcDAmZZvJJW7C6n/4
yMAMitsyeKs6ZF3ZYbRRq5FcxhtzqPVyPSIDxuSRGH60jpWgUoSt1H1MNr1MxDFqlRsWgDRU+pYO
UhGPtQ42GCeINknrbwopGuCUw+o6bf8igHQGlKqhBOTlJhrwG8SXkFl6+Fj4SDI0M1oEAVxfB1bj
sA7PH+4GrVaCUfAf5IPNgC4kTuJQnaM8nNev28DGwGpioAy+/k71NiJuS7CLJobAxdE02bINqDn2
Ai4CwKaqiXLEQs5yWcH+XYxrzPmbCN4W5H0d6ovSd209lsAomx4+AIPfSY/kfkQAHDZpxsoBicDY
1NSt3YKsuK2YPxhpt29WpAZiGhIW9vewnwJd4o86bT0bwTYefZkRvoASJhgKvSKaTVwZEpY6FH7Z
RQbjsle5OG5ntg3836HxgPBQgNKr0m7MwO3foOSxTEaw7dx33onsTSB2fm7bynCQdkLTF43pvBsh
cUh6u8EwHK9KEZwQzL2q+qhzUJs27UCWpxWDTLTzNrW0VQle1OYPZTKIuf7moeGsumcmzcWSWzav
hgNaTxlyNfhZkFo/d5YNFLAvlRJj+H8+upeNO/hrWPAZEx+jxKoIh6UBJU2F2FzcEeDphMPe6vt5
2pDMtJzu2aMM0VUw7aLiAFxtnd/lqiBFL2Cuos9AcvPtuUK+NdWsYdcT9+uOYgUa3HTs2Aij4k5f
HkAx23v19qa/MtZLBGy8bW6yOugmuvM5Orskzz4q6qJRZt3vVY5zvoVvX9NTDV61ip/KK6l6Sqma
b50xUp0loRLefh9PDi5o3wf6kiGFabWONwlW+5C1TWzDfke0260SNm2SOocmqSRY7WBfToYNpWAN
B4L8vwU7IbawAgd8mnTn4XIju5rlf80Zk4HSdV/VrsxlwHslK+Nvc/xgF8otlGOkBGakUPZNNEpa
2J18+5S//OVytAuB7D9YwejiWjcv/QdbGO+CiplCvPMMuau9wCiBOUmlZnpXYxxBT+6cM+1v5sox
BKpA3f3Fn60Ur2obJqPF4eOL9E2J/6YDI1kDgz42IQV05DkmsqjQESgAkdRLnXDBIrDVwQySTfb8
xdbAwwxTc/kdl8YR1ss4Js/3WodRXdybEmTvSzahzM8KdkZfRDGxV3EWxIWL/+UTllCU4Cor/B4n
hsXU+13l2pXMzW2mIa781rVeWVZIJF86l1614lvjgIKkg3nRVilHHkOA5oFCAZ/2IFgUz4mowuOL
n9nxYhDz337sQZiC5W87FWihm4e4vUd9n/I/SvQ6DAiJik+g5bLyyTOFtFkxnKnfjJQ3YgHWt80O
uZ1OkXq+4BUJrnoXc1w+gDWE9oQ0AIWpFyzw+yDWitdwoJo33cwpGscujrpRrtwozv2yNLiUZFt5
m9EkwXL1eMeZolftlS4a3jlbW7hPYOPmaTxRNpvxXRlRN/xO3Zj/kePPnobaIapTZhqQTTpB8hRu
jZVlgxWLi9epT32/c2GEMzzerZnJCHiql+bab9LFPK43xmEoJxm3vUsrKROGY/xZxpwAyLpk/4Nv
1Js3JFdN4aOxtvSeOOXhYgTc5n65RrdTTb6AqEg0sGKgpHoTut4c8BUPKEjzHJ9KUvKm4sK+Krkh
wwhUS/ghHhDsbrkQF87HvRl5CkVnEA+fY564KO3YPcUbdUF0NzAfmmIjBfGoWBQWMrC8md6Ux55k
1teN5BZP1DHtETDi3Yvy7AIKROo4vAvyTtE/fNdldmG6M7256MxwRFjhFm5GUKCKSPDjKxgQSDgd
/9noZTTd3cvd+uLU5vkws1zghDWEQqD8EYIR8iLvThc19pVGgClvLQQ1fHMzwZdi84H3m1Q3CMt1
8Alr7INQ15JiT/OfKo+TWFjVyXQoWoBrMUoA+NCk14p0/YaGfmJpG0qL3xsNyuot5UM2Rsw6np9p
7W9XfxRiUAaN16VjMtwu/JsxJa7wVQjeNKRIH7leTZodJpwJGQWMOiLGU8CVKWZWlB3ou4+C0yse
xTTA5cZS42Ik66I7ttTLwjeKAZXESo5oeEGM2nYFwBOPY+kK60MgH9VmDUc9e4W77vaGNcPcARcn
t4K8Y+kiNzAAdUKaRRxfnNeQHdWpsLcFP4bXoEeqKTOzlTufqXv/sGSO30Va6PrZZ7vGoWqqTlqy
txY8jzRP0z2BfLr8BpB/vIwVIG6XuVWOaezyAnJFvyEBAu0MUsvTIgNLzXbnL1fsLWvojZJRDJPo
TUB+7imya661ntCl0E0qAtQmQxtfZ/L28zWAgONrbrDwiUp+CUgDHoaO0QaG11EOy7jkv8Hp0Hus
/QFKG9Doo2wocg54mCK3CovnJlQY8YET8wNEw+krIlwV1Ef7drShL7rQZkVsTFYAt4gxYt9S5REY
+d5JaIsbURRG5RFD2j3YF5Um6trGr3UT/DkVLmkKJlKU3IlXO8YYUR53t7L+3nrUQyEmcq54EH1d
Ki94j/2V2HetdRR7MEF0rRbGumE3MmQUEqFW7Y3bNu275aLhB7wWlXQ8yXYK0ioJMnsrQ/jSeLUg
0it4T++lD85dyRX5mZ6vrAx0f/Y2IPWvf0futqE8OmQUdA1IP8PPV5D5m58UpUjJSupHQThwwBDB
hsPw20Z+cL69OyTuj9DMfJdkmztIBdQ7ptJKStgnAwEZSU15J+lnYTa0GLRgk2kq/A2t6k+QphN6
4oEDWd8flyHAyPKHyfdds99nO33k9CSX55Q+xzVG1TPyjE7PGBXZxnxYzFy93Oe4tNbP+x9reLbh
WbSTimikypw6aEGZPCwOEx+M/KeZfQsS5/d3yqZgt2VJShRA5SKgzsw9Xd7T4mInx1jQ+zOoZXj2
3JE+aqoLPXbTKLgzGU6YeZjF+jbeWr6N/h5Y3m1iXQSPBLDyqnw2nQFuk6RxPM2sr/EvC9Fmm/oh
0FSTTx5anzsXkgtULkpGUXFRr+y71JocnL8ehkLpuYs+k+v4/fkldohsSYQDNA+OjOxNHZePXsvO
Ez38mwh3A4IN7IKLBTwLpRp8I7LdMq3txiawOTQlrjFSK5KlfjtImJZ6NFlBIV5ZqgJTrnzcVowC
ftIHcEDqaZIBYbb2t9/X5udOqYgM79Li8Fj1kA2R7D2DUK3gXuD+EkNxyDsgiKNsuvwFwTCBAc4E
9Vx2SUqVtXNO5kYsCX3+tgfULdp7Soz9NeoyU3HB8IyJJ2hcaLbnFAtvuGfwsh++bndkUsmJaSN6
E+QcWdhoDQTEAl8yNJ+jNKCyoVYPzKpw4CZZewZKKKoakb1R9JTIs0kbuIBgp2mMtgRfdwnsa5wk
Xy/tWDomIRP3nGQeQ6ywWbz6psSQn7nywYm5PwITn37MOX3VJ2cVPsRZpt5QNWlhWoWEKU6dxcqq
eBA9Y1AaubISjU/Jkmqo1ZGdOCMaWNlWfqGBhCyoAffl0Kj7ej/WDIO4hktgC+ErQdG2oHQBt2zP
gfePx6r0MRpBL/k9MJEOaT8BhirPAkVMThBmmrqYwAdKmK2YNMxvjWAnny2FoedpDGcqYLykTxia
aWmPNCmntu/vaagFZrpjLMwsOSwpKMTg5OtieP4RUDebvjPVea9+LdtUi41izyD+/XyYrfBRjtjx
RC2YxD3irxJdC2f6Vz9tG8wjdeREK4V5Scg2i9oeuFOsOpz0Q2W6bTWRt1s7Ib1RAjb2wbsk9jNx
1ul9Hw+dkOxMwiZPOppjVel6ozm7cIvWvrUkITVjuqMiaZSN0sZPtMaP/AuiMhrCJLRsGGzqmiaa
c13cUjEozf37CuF+HwAHEgNEuBRf17jsf87v7MoV4Az1N7AXEyk12KVq6ht301vLWORmMlp+byxz
PxJCl3vH1B4NoxkJ+TXBCr6HkDWc0E7S5CfseSn9i1uKCH93QslEx6FlQOujGWJL94U0N1uJ3ZXY
MYP0Hjw3Gw844mpc7nrq3Xxj0oZwIDnevoBtT1eu1lc0hzC6IrhnkrvWuVv56j/JKznLKvMeGOWw
glvVVgfEvIEP9PbK6VU5wonK4vt1obCl5bHwcUXXDiAMCTOcVYWY6cCPXCZ/pVqk//D7wWoPIUdZ
EUNLHm/5urSPKMYwjoeQTw1pSNVg4B6r71vhk/isRWJQs6LS2NJTrWdfUdQMoSGrq4EYMGmlkFIK
FtNmcJVmwn/OizMxXPBpEah+Bd9RTLLrVkMqND/Mu65I6mKmrvTFDx/MZoON307v5wcMT1EwXO7t
yT1Z+2LSe76xFBeUDqo4/JewzXpjX8BjuHtVl1XYHO1mavsKj9Fw9gRaOl9Btj9eqXEYWNs5ci5i
BoT/OH0w/GFc8wpR6dM81pGMkgzhDqX2/SE0VKuvZVoXZTD+UpLcfN/MZiL9UsboHR6y2C7Ca+sF
KwXwiTw3fy9E5R8SRiI9MMNfUNixA5jeDQlD6QCceONeK1vMxUVHQhrzJ7HOU3k+iJ/c92I28OHS
MMnk1xlw1vWaK9m++zxpNzZrTt9uWhb9vJ4NW+ok+uH+o1oGJCg8qP6vFxQcXbqDlQzXxXdCjENU
9vEfOWOc9dHUAcHNfcXwW3nZ8RSy6ILJdhKeNAXEV1ZzwW/vGa9EApM+DiY46IBR+GZwJ0I4AEOf
NBqPL7zOea1gq4am79524ZmpBlaG0ne2JFf9jXMCzRtOHUwbdktwj0tFrRBrWxk4+90Iur2VUUYk
zd8/atRr8Up2RttSF6lliCKqEYDhlgfVNrIdH/F9VegHcFJjaWHcbrwp1jROD5cYe3wZxPmD+ET7
WRGiY9TYP82dZQ1hV63jbV0VXk6p5RCLAlWcW8jbZJKj6erQNDh9P/c+EGKQLb7C4Lxmslm73ic1
zdD0yf4KoLfPnlrsBQ9L+hkdpvNvZco9cxbui/ROMPQ2D8uI6UqcodunqgMGF+zkK3Sl0FMOeCyR
nDzRBggQCsWFT4QgZ0HywZDSWyVA3nu9pWQoxyKc7ed7gkzpJxGRhMb1R5RpXd9GoTEQ04HKCzS4
gymhAQI7KRIAljsO1Uf0W7+22Gd4cJX1w8fQ83XW2i2k0PlyiSxMC1eLTMU1PwLKIC7gp5Vkjdvi
RPnoewWH7O4UFK/qELMos+Kx8Ox7fD93rl6WBgkM1kxEAd31nBHe1hzNTztdTARv4U6PkCSw6H32
QV9BbRug+p3S5X+DOe6ON63y0ZJ8JYrwOyRuETEr7cNqdh7bl5Yh7Zl1LK7FPmvppEQd01YLYUWn
bTWkkcJt9VkTddvCS3FQCB9V6kByWPDPYrs1ZdxZQ6MAof6c+HzLl7LTJPDV6sZELV1wRG/MTvgg
v1Olme/W4hhvb4CIrlikmzE1wvlR72BRSYaaG85zSg2QO+cGSGQnwlGYIwUFNQpIYWjRHxUUPNM9
vhGkuvWquIM/HXLj4hHXv/fuskyueYXWtpO0awH9COc7aO0x1RDUqo+hIwthz5dlwgR41sC1/Ebi
2THeED0ibhyjhTm869TnF3QSbLGM6yV4F5ZnXDKsDO3c+5ocoJ7VWsYsctgzPGxo6QvUuQlzU6v+
vSnISrp+21ivAGPtpRybRqSoDcvAexgOQ8p7J0CEVzgyN7ot2nZuX4DpRiChg5qXeQlXm3mgah+M
OTA0rObN9v0vYfJZMOneywU2BHLeJuwwfiaAG9iVvmGCU145P9jzD9jwsi1Ocpf317KUGvDOVw7H
+IHVI42p/6avWNxptczPmtVpIy5w+I4qi9m5jAqY9bdkYDM7e+DOQeL8+E34/BbAIKirjNaS25NE
i3bevow1qs8TtVAxemQyiI05Swq3rdoLujdG23FkipafuWt/fjq1qvr5I0DWygaLcvIsQDmoRdyz
NVlWokJk5k4px3US39hmQxM5H5DWUDi9F2Ybae25EB/Er8ojMtMChnGWO7qS6NVq1Cd29nf3DFRJ
qnqoKpMyE2eDJhxJ+BRVYWV0J1EgOMt6j/t6Wa8WigKLdRHW6Sk9an5yk23puH8bM3b35Yjqhfgy
1+icO4tWVJh7WJiWrVwd5rQnzQ4jgV7/2ap0LicUWDkcNQcF/ZX9jjKoyQnKtgaVhkSnUTKUKuiS
HPNMCb8/PcRkVOWaYeSM9H0II2XTwyP6bNXHbcuUP/64702JkZZIth0NLy0qs/oR8VGPgIi0DZS0
D5S6kunn8OHXSoZ68pQSGekHcCxmHFucBbweL3RxGKjOpG9bvgLuYj7DiFhoMa8AafSo0WBDps46
jDExW0Mz00mwdTnhlYrNkjnMZo09dn+thQ7oRo+HL/ksYlhfzg7OjqRgcxpjmyLExCtcNde8/Jk6
gBAF/6hWHdVcHhw7ZLD6v2v8zsTc/JsM8H1KlIydjrphPMxnIYtcv7YJ+QpFQMkIM6uZXxCMChas
hxFHSHOWNy0x+yslzAQZxZ17jhm4NgTHr0ldmJq8+cahNTMMUd5Q6rl0HpA3dJP5tdkZ3ImWYIEV
DCc6whdQmbZh/QQxaytRY0XEiIpBOAV3RDr1aIAVagUJJt8xq3Cq96MgLnrS8r/RGMBsE7Sdzlvx
qe1I06tIpIoC1+raItCZkJCo+wNX0dlOwiv6hc1Zm6zdm3Kb2+CPQ2R3b8OcDigXTsvVLKuR9+Wl
8mUE+50KbmFbPmEwkZn6PZM6LfZTaj9hWEJ1JSpsjyPI5RNb3o6tybr8lflZXA9LWIY3E7Y/H+kZ
CgM5UPz+REX/q15lqt4qvYWmfbNK6s+agxDg4XeyoJlJeDrKV/cQlhXBwtcdG6xoCziixszK7CBE
5lUJPuOpdDAjeAA3aPlKwKH0fMh2OGOm531jfZ2c6d2IKge7LcnM+yh5HJ3ZxadNyNJJw82U1FXj
Ae/hH9YMtIl+BVk3NwHJ1UYSVW5ehKdnCPJbi1LNIJyJoAnZLSdJDGE7Eg4Ie7EI+W7dyyk66lqc
ZS2vK16JBksiz9+YPsEQ35cdOdre3QYtT0Xy4+4UwhFPinhwoqoFIstzStVhd5wL4Ftk+H2F01cu
dXOhwQo7Mfj/JLuE5nJmd924PhkNrfPV2Wd4+1Bs0VJ6DCjx2BW3Adv3Kugw2XX1LzI+7MeAkgQl
evTXnyAUaP6mR5vd8yFbeJ/2df/VC9ma0a2kh05vK446rvI0g6NlmGPor+UcHz67yWGJoyidOD70
sXgGuxJNFMX8MuBMzfV6mWBRtTBehk+zML2YRAFHAiXiXoumz6S3G/pL4xj07DyG+f5T6g8nzDk4
Nu2gLu9eX3P73Y7onNCMyrNSqsI/PyeeSvjSViuY5PRKVDIQrcRjF+YqgIGb7+GvfYhR1864P+pY
OlewlU19/UxiSLATV5u7FV0GFcseNbKHj6+psZ7dyW74qFE0pPtgeLE3M2Eo8c5HBNhgt05ialn8
E+bSdobYGimf9FfeYfd0qsEUIzyblo93jtOzk6PKV9QhG/fwXp8eqWdljAuouswlQBVmk2cnSwH6
jigDJMWHtHLnJtYqwgW7OPe+wwiEzFLwQQ7+a4FE8eir3e4Y6Ue2hPXvIo5B7JihlVZo0KkTAm6R
RXSwkh7z63npPA7AQ9cC3NtJ74uBKRCoSW4f/dfawa0LqwmW84EHiX2QJ4Qqww8yY6zKAifii+mf
Ag/C1NCUrWmipw6a4eIZlZOjZnTuf6rciH3p4G7uHmIlnR5C01ingVMdLsZOC0QfqXg+CLvP2aUU
2OM6jF9s0+PNPDcytIKX+0Ik6S1b/jV12VC5oEdJEr+ebTVD6p7ID8qlTWnfOM09QlSTMmP7SSQA
epT6IXwpeZovQzOCOnswOd0vWNVjbl5zEFmQFr75bPqirTHgwcvSa73qoXtLk8a9+uLA3lun3Ase
mKASaS6XNr4tL+Yc5PAiVKUAdK9nUqGKac4BeItRU6e7aIrHt28JUywlucfISx1eDEsKPqLlO5GI
i5XYlAdjJtGQCZERS3Jji6vRZrFZgJykAt3XB52A8qLvxwEE2aQ9ow8C1r00eJ4pW6PWGVUjz19X
MjFsZDu3h+ddAI5GNVifMaCWnHIX/UC9K3Cx5PQ+ZWgHmlJoEwPGs0bkmYnWjH61I32Pf/yUcVhn
AA/po1m86MfzACBRnt3xg8kox4s4YOkU/iBZAbXg5bgmXGe+WeyfXuo5Eu63dLNfIZWBAg8Zog0M
wtZ4IgMl1disNSPIAh7QFbDWzolHizoTXwS8EINhyLz9Nar/0A8xoMwMuSIaR+WdvyfMzBL0WzG5
zn8qzCU2OXgRv6KNzhNGs710N+/88uM2wj0j1xmvv/UT9kgIadI8zwaCwxJRIorC/A1rXZqmgRWb
vxbq568u/NNs+Js38CypvPANnK9s2rveb+A1YwX/d4rHLsn6LBDRGbQOS89XziliG36jNF/8O7Cw
XSvDBJACWv0nRAFZAbDiMSHzjt/x3sc063/+xdSTaFn6KYHevTypezUfgD6forpSRKuYF420ETdS
nYvCzWu9+IxuEYn1+BXLemaRgffg+FW9AK1VYnfAYz6b9JSL1FoysE9+ZMST2GZXyNrg69a2q4nu
xCuUQjAS+z4o8LENnm9i0e59/Fgl2dKBQq719ebf1ixI37sZGe8H5HR/kvfHKukE+fnKbHnaT9tt
KIAdgQjjDdXwbsbqP2O4Tt7lnPZQRfJk7A0+7pBpCIzEHqk8AQGlsLusH1mkhNxhThNiuVlripml
EATf+ycPYZcXkkzS45zD0Yh71jeCLG3hFNdEGOu/yPqMtTDSBKW4JlzRqoKMAFjTz1kO5A5TH+gh
NRGHb+s8cPpTRl0iyZw3UDOPDjvFMrzV3A4thapTz3Pw16DuouNml6sZVVr59HacrCjzqfdvUlrP
9pR+mv5EwklLqzFhOXEUncuGk1PMpZ+LLuma77kX07AJcrLTf4aSR8KmwD+h5CgQZl6onKYd9fJq
tS+htpMHHA+CXgr/SInGEsXyz9hHXmup1aqjHW0xBUWIfTuMjwrHX7fnY6bQLyUBq8wz636Se5W5
wWSScvzTS0MuabmxhcbULKfU4s4dOfhE/T9t5NdJvD37WfRaWB2g5uvFWdRwKYWlIL5lyowP0Q9D
Wsi+Ef5P9iBS3HbCkgVk8o7BOX4z5zEd09bAakdMAtCAQouBWxBDAVD42VLSVLU53lYbwJrAtjRu
7r8e+82izr7K9Db7W3WiXCT58o6LYwF+cX49bdilAdnsoqDjE6xI/PXop40Lzhz1gwwJtg+5kSpa
oimPf4mCVlyAGu2y0Km950hC2XR3PZStGxNzoNT0WnO70Jq1sMBm6ao/FedSb1kfBGjV58Jur6ni
sKIv39VuvwyCoT1yZXknSVpdRyTkX98+nxhpJ2dVlfBCVKqpSK94CJc+JdGlGQl7BWUJ3YBmPULy
/wZwSM1dSihKVzL8bsnLcMWTonXrX4u+oGqa99knxO6RFpRbmBC89lm5Q6FX7XVitMLrXtAx7aYf
leG3QvkxbsiT/GYpi9NNLFw9pFCTEn4on+qPJVqCl5GCdrVx6tHZzqZeRyK2GylFe1trHbruVtWF
FMpD2VlJa+ZCkPVuTyvO1v28qTrmcqfBlIaeP4CT7BRE6OCPFN6xkP5vQ9et45Z5GFDOb1Gd0OeW
sI8QJ6PTbzXP42vXFbya2Qdnm8b3xTUf/YwtnhxYkRCb2oQmVZpL/qSFOHN6j2G51JxeItEwvB3L
bEx7ydJXyEUY1GL+nlQbErseeR5EfuLXXiT6xwHm9EUS3pbxNEf1+y8hHflDMjVMt546qrqKb2tY
F2nI2SDPsCuMIc4Ddu6HYsVlSXkVfeeW8ghhywb0FjHyV0LP53xytI4PY6Ug/HntTIvlhEgE1Bad
lTDqnBrO4/TKOvZrqA9vRhVTyJ2Dl7cyEGKkQ+lZHAbph2ZkYP6puPrhvuteo/oPbfWVG1NAUZt5
9pESk66BaccyLc51IGafipbpuwTjXb/n8G2euyaSDy1g3ohgDMvr/gtdiMb4I9rGRA71xS0eyWXC
pkI0ir2CKPBE7xHLSASGvdTPN9ZjglGIf2ikPcbqR8ykoRrus5LXTOOG8noLlJ9N7LeLV5fktiwp
4a/GqR8PpkJ2TonX++37BIEGBGeQ62X/vm8Gwpn7i37GucTBK1JwySvEb2WAU6LmvXJ34Hy1hMcf
Xh/fCoPwf+QkZC++RpyDQ3ujG/AMeNEjK8wttUllts09UGTHCNt6Csan40f0BbdhaJbZINlmB+DE
EiMHT0UldRmo8pAaXoZAV1etlGYBUnq4jHDAmoIvLAU7W77VYrDiSFpAt80sdPZlMd1ESfrOai9i
5cvyg5ZcV/9mNXqyYKeaep8BXOEOP60AbbSS0cbh5TzPkzL61MiEpeHnl6dLdFNcVOzctNpGXpa3
F3fBCCSD5pAu/yFAo8D5AvLJOnf2569zhRPkyWm8m65ghOxS9VMwEFJsJszpzZyZ2uGcPTeJPySP
7coKoUTQ84PkYfxVbwuQrukMPBe8FBdh+zr5EpHxQZNtSOPxPkG7Nafm7PohHHe2tHL+tMc3yqqt
l21S/qPyH50mAzQDX9u0AQmcE1KY3mdY56jV7lWu8skqX8QxerF8/2t8RfQHX2xivimt1+hIbdMM
kAs6GRBYkcxieVewVJowaoJYin4Ama8wIxIsoPyPJY1Xo1GauP4rtW6zuY7+5R5YyEfCpYftbex2
mn2ioJyZBZ4Qj2A03gUZDXB3/ULJQ8l7wK4/Hs2w16p/IpRyBL/P8whEiPpGOKB997R/T/M0Hz2Y
rCh/UVTniFNJCkE/KpLitdhbJYNikK3ay6Q+BeCnJmFf7m7KCa1oOumG730zzFWP/z2SVmbLsHTX
AZLUQ8ZXvx8+jgN4dC3j+MaC+vwSNBJhsDSa0HckFcq686LdcXhsev3mdLdsRZSDZ55Ywcxk144G
WXPLkpcSiize3T+HXFaw5qqRAXBblzv43tERzO8hh9huEF2bq0mWzL9l6fbwr9IRUUNxqyx2Q16c
0wE7RWCs2/d7eoKe2mBnwdOqsc8z34VC6UPwdTRFy5V0JoOJ+tP4CceQ4eyh5DRNjGlX0zqVq+f4
ZyZgu41bbebrBqk/4N5KywcYnTd2smm14sAxCdO1dGNNh2npXVbXhzQjI+a0l+JEoQxrh4RbLUZV
fAFqnCHMZAFvP+49tkhZD+VdcqqGUlgzsM9P6Xl00yYX/ivvj7DM9gExrAAAh1TLRdbeUoFZNazB
80kBVmjHbks0sN2blMJd9zyIn1i0oCsLQuIg5qriVThWorn7Rz45lOyWcZM6YevFs2Lr5I42QTki
CO0r0m8z3p1n+sjRClorIh2yZrFVwYEUxci5mqljpbIOGvKIbHd5fbxrbt6gGKma/v0MxT+WSFNc
B7Sy2nyB9xusf271+i41dW1BIrgyqSSii8mBQExtDR3L73bx3GBEjt/qaVeTgcWylewsiQKxN0qa
+DS7PnQWgChjv7pCb2YAO4lWs645HtuX0+Uimb3reMMWQ9gOWPf8C/E9mApEBDtcsNw80La5ZzkV
Jt8yeeztMkv1Q425G0AX+rOrfdrXblO8JPQF6yeRNUk6aiWMdPZKzWA4P6txZAhthxAHmG0C/m3W
KiVa0LJXgHZv9neTq819+OlRotc15paULz9Mqep9CkKz1713KHtKg+mxlxTyuEMw8sWhWrdsnM9B
bQJ1XEuqROv+5lfy6wbDK5XGF19RW6HeLqE48YVD6PvO+WqiGiTTOt0HICuR7Z14+HWRoZeTkr/e
MbDsycZFh5D5z2LAahybjzVDzhZyY+rG86Pmpz+96DOr6a4aCsTMqtc+hC7H9XNBNqe8x/A+y7Fw
OqtxbzsNMwslJMIni8EeiaOZMcDJM/zEm2yV6KejIuybrhMuJTL0NWHnJroWT4kazP8AJDTdwoxQ
SZ+oRyCtP0FRkk9Hwj/TI4LYYX4Vri9cWnp/BE1sAC97fW1322bziJ7LXmGqcO9nGxwdpAaUZ1RG
aKz93t9wBz86ymYwMAwoXx4uRE/0F/P7PqqrxC95wBYLqOSE3ObEA64BG/iqQeJL910NNoFbPvcu
Qc0zvmaz1XyZ87hJ3gPpJMus+taVLgDNe4KaJ6lKtlyUn9mlSJaPYTFe3WHxfmd95zu7FEDJKxgQ
xfyaBbOD+NCg+AM0fHcOrDog/tj0QCfaRBwm9aogrr6ehwDOwDHa2pxB33RJ9uvifD6NNZmuqrVL
0H5VrRWfPhsSCB+ekKjpz9wQJv7NVkeKfTgbCR4npg9keNNVeqeMgHGcBljXNqfVSA6bXdvyzc//
C7kVONh4aTNtddmemGAOs4uCAeCiB9z4qpQZlXyb1no04so2a3PELUFU+JeVQuIY2wDqb3h2r+ma
AztRHP04oMWw2O5jd/c5kuZtyUPBPGR4o9I+voyuvqoDyG1yI9HhwF3RU1jKKAFEFw2Af3/2pLRx
WFAIfeot1/9fk93cK2RmU5qBkhrO0rJ5LWTcw1FPAJLPEY3ppHipRQPef0CYjX5QNw0QbeMYqZmb
OgOK+xvlQdnNVcFKXiT1qD+mFSNxWfInvSjH4NYdnNnuwrg7XhZ+pn1KEkuB/JMF7A74D4ME25HK
QVfUmnaSuHHas/3PvbanYf2HY4WsH569OP/vkmme/2iOjRhr18UzK3m9hLQ3I5+XbRNfaKICYKAm
KNqqkpxqij3AOVxeETw6K9TnZDgN7tfjezIwexg07PwpcuJY6thJ78DkU7ldAO4bvC0aEICRJroM
Ow9bcSdgz6pcINp+b1BGaI2CCLippGTv9xXPcl+B7RFrkbkUOKHjl9GJqNxAkOYG/LI1ZrpSbvfc
pWuUBXDEBNwBYY0LlVHEilqifhyope096dZY10E5UAv2CtuvnPxbd6pPav2rfNoEeUjvipTCVdDO
oaHGTYEb+au90+UF88+Y7aoBDTlSumYHANy0H7O8KVnnZ+8Zt4ixE2lK+uYr1ui++vmIMBbXwWvr
p2he3D53C3/TeVcfmku4Om307dU9DJLSmn5vAWfhL3QilqGWp31oTDA1Myx/EsXcwzYVfiFrbXMY
w1PLpvqCiLCZt6hWBbJ6UhRJByvv7RSx1wHymXnQsiJkrdquST2dQ+JYD7QqnBcHe2LCRfVTAw5w
YMMLzV0bTSDgtu3PisWeViRQyo4xJZLTduh32pvkGnGaHBPyskWQtayefrFCyoYCkqhjUboTHT1x
Bj0jntwH8AEwW3PLIihGlFO8AB0NpNl0/abL+iNA7T1YmkNjqrOKPhKvhpM/FN0kXgMQn68MNun9
dClh6cHmM+MrvvCIYZwnQVWeE3xmjUPfQf0RZyi3BUG76Fr0uD3aY9Zqzy6R3giG3VfXwMsUDZtl
mcUEcsnEGD+yq/Am+9zAj0PBHbaqc7tIljzEkUWFuN8Bmw82na6epFe85M5vU+CpMsOFlzOeX46q
6uGpLb6NAruyfHPZAI4BAv4b2aX+y2F+EkQpL8EvSW/9ebewOB4cXkp3aFJLZmBYM9YzIfczrpo1
gpRx7PoVxKLZieBcqR0iK5eTNPL300CCSiRqIwWMxwJZbA3lMi7b7BHnNF05TpTv6u3g7QxrD82V
0SJUWmA41MocWEPYLQBFpNN2JkkX+nZdCvo0Auw1f6zegg8k5Q8XOYHEhDk++CL3J9siUjPMsIRz
/gbPZFao/yS5Wv4izW3Sx9S5rStPOXbYldDzI20kqj6SR/1jbe2pPO0TwkRXqFeqJdbRRzJWe0XM
iSnaUjD19A8piai35LdjCvTiEjbfj94N7FGJfS9cyGgekckplRq2QNHnBG4y2H32pBkjHIKLg6z7
SzyAulAB0hMDNyT4hm/sa8IQm6D5vpwR58mDhVAVgsSRxo4t8MXR3k6A53kyta+PnDs5pE1NJUGm
4iq37+8UgXEpCEwYg5oj4Ac/veumWxdqb+UWgv4TaQsmxKu3uiTC+okBKtCkTeuAKJnZfdX2B4Dw
zknoswgPk1ShazAMXWtWsMYSbynPaeZsOIATI6I/uKp3D3rLwaxgbXuWR/v8HrimiEExErzfWKM0
gfvQ6C55aeCh2TX0I0eWaEugiF/LU2MYAtTBz7c6GHOW6Nd+xqKrB0DgE0V5U7i+ViltUvM6KaVy
e4F/WCT/uzkqbH6ARcH0sITI9yUezZHL3aNDg+RcSL6eOzbob/BZiGG2FNT9XEzNrvOYmG26swbE
yPSD14Ur4tSb5Xyotlhe/OVGaWjUBp6O8H4Tw98DNnJ+OjQ4gccWDUeQy/eXoPcm9zl4I0Ub66O2
ik2pQOGNIRhpz7HIdeqpk4V82eEjTQvwy/8HeAy6RSAa4RdS9WZEnX+ev05ubj3e6S53hLPG/J7Y
wkrQ0Cxroj4je74nlo6dZgJxgALyfeMOJWDXfA7jpmPplgNtiBdFf22r6aVkIej8yfsmELMcmy5D
2ibtmK5sOgUOZE6pt8tDiMFECwuTrmJf6fC8YJGKlCp1e23YsOF2hC+0eYZCxLTkuWgtGtEiiBsu
i598RHCVK4KmrucNWlyKSwO+g1W2pschFQGgv0o7rToBtPLUeEqEeS6xZcEDGDOalH4tA0fD4ivS
Sgyfq+AZ1XZL8Gf64eF6jRUwxc76jejvFxq7hN56EuyB5WCqmXPPiursTpWJpJe13UFv9g+zP0QR
pl7Wt7JIg/tz6AADighvwUd8AO0JAflDWE3lzQMiLDkGXHOdRIKkA8LhmIvs9YRYS4seKEz8rJYa
kN7wWpAnekcqBdChwDKKXcJhzmmbglae8li4BJqqPVmE8so4VyhXnCZ3yzjyIcLlBjARjVuCSVWp
hzOUIPfbYNXOkCuLd79a9ZZGF4Yi/4IbjEZV9UAXcccr86dqz2kL+E29t82HSYZcmtr4aeN4laAT
lQxDbVf6dixL3zCNZqjEL7KwxzeKvqbqDrrgp0pq4aka6+JS+kTz4Ba0itBGqmxEdIE/D01AzYI/
2wHjcQ0iuEvy91SW1AAkh7fthQ7LnMaedgDAt0Dghs1Lsc0hN4QbAtteSJAsZ7qynTHQOXLb4ikC
idgpA22GYuoV6xzFyrSN5iAqGcqW6an7r8NR75CKJRse3fwyfl7DN2t/Bu+7NSWXFZpeDqdM52dC
jIZulVibP7fsLHUAA+SQxtJ2UR2yrR2Ur9L6aIilGbYXp2SON4nhiwK3D7TozfRZaVfX7aDPFKMQ
2EMGUjsmCldXhCWAxs+ZDQr/9gMI8qM+ATUQzkdTzT+FtVrzST5LkjTvTUe5/eDf0+ZnMXcBg7nR
cBeciNIN3NQYNW65xSJh/XEn+XDEmBmWMDW5yEKFnyWZiKo2T/BN9v+6SstNAUUiTDQV6ElPR1yv
EDUw3In6j/Jjn/aybdKF8/89nWBo9YsF+rxdXALC6SH8f4QlFfh0wTIXx/YW9PRGT6+d+5g80H2X
qRRN5FvlmYK2aejEbCkbgPIsGwBxeEh2Z+QEuIcyL3jWKyLE4b7y7ciOnS6PRMx0MTTnTpID9cPY
uD0JfLx1m12J8yJLvg1qrtcfovCK47jpu/a6fEtIpm2SF21QnGnllYyJZJWngERKqYESOjhENHd1
tr2bnfpLwKIHSJ7FZ+5wRZDMGgT1/dd/pIj+y2INjNNf0YOeSCPvAMUikvzkbZzXa4dy+0LK6s71
GBCqqn0BO36z7qYVmTo8b+MzvDNSEAde6n6Wih9jamjGCqDxreD8Lw6+12wFv+PSsYTfVLMXjTyO
0wwSAZgz+/c0tOhH7rHtRQBi02e76p7a82KHwlux6IIbPlmsXOcMawwCLhOkIhebgPL17edCEzjM
j4DzY+YmoW+hdKVjObUEkaOMXSe8LYLiIoTy0siKxOIFcr3fCK7FAlEBsj5kpYrdgQwgS3zj6RzP
osCdcnO87PV2UW6wk387LxURmeRJ+32HyVsj8iEmYV7GHISq/PmfJpIIeuhPcjmk9gDY6lx2THmK
61zcTLOJcR+WLznKgzYlzZbkDLS90kWwDlLGCSc0GvkkhaVJalPTo2F52Kc9vB8GO7ydZCjS5617
me71fetk6h/lTy+ig+mzotMNHPVjFlVVAGgh4l7PHYoOVsRg/UraMx6MrzcZgfmnspOCTvXCYG4N
RmVooqrNpYoKseQNYp9fWFloDnRuomMDHqaRRkc18YL/jD9ATx+745xfSdznRctbTkd09tKjlGBq
aIyKO8fOosHr5gvpp52UJ8O3UtjqDB6VT1mlwEoJ2fCuWHSz5ncBfU1cW/jOrsWoEXkutTAj4v2g
hlx561i/wNgGt8OXGnYMtYpUlSI7O1UCJJq/5Uxs1bkj/cqAn16W3uwpGyWvQ/1XZbj0URgeU4zH
EE2IYJTM0G6+wcBZPu6QcLwoIZbP9Mn/lMg39Trfrb+UwSfnX9DFXetHOsPYrF40xlNq89UYL2gT
j2uwmWq/1FKpzAZozjf8TwMz44DybCTCl7CZ9DKbo0rfpKvukIjLpA2hIpgAgW9urC7gX+js3oV0
ADgRrYhbF3pWGq3DtHPO4VhN/di0OEltId0VLSILm255Hjm2PvDbozzMI29R1jKTyrowQnC/VvPg
SRuOjlmrAkmWyBAG1Ob2+y2cqr6odgPTkHT/aIxa/LcHnUaTIEycEKKwDuVWLAP3XMrcTFPVSy80
mtLRjahNpmVrqm0UEjYiHERDpXRckgbm8Fub3LuGmF64sFTsJ1ByeBfjfvZoizWombNZdwjHMWtg
haIa8Khxb96DyIReoKpZ7unt0dleRMGCkU83ObR3NlKWDvKq9OFTwSrqQV1XqTm+aN7exW7n8wEl
AzSLNcghPqOKZO0wC5QaQljnFTyVOSm/UAKWhjWC+z40nKQVAYzKuY8/x71LGzSc+PfajeWS+MgG
MNV/34Z8WNvsZKHVkaAhoM34RzrxwjD9j+AaggRjLCqLaAsvtvdQiryhzaqd47u0RnNJ8bDeOdJh
KgRMlT5zZ07xiwx+L5u7SJZeumAVOmjFFpXKQsD58fkXAbQhienAEybAyncNdHlGTYtdb7OV5Qm3
VtvcsmlHK7qECClcfyQPdPQZSjpKqM1+irK85PGcunuuJq8iIEvdfiY6hMS8G/b+zKnuMkiXHqmk
C6pboQJyDMqnECw6fBxcn9G8zw9Ut9/MILQpTxwJQD/Df1Aohb7K51yhFxa/BXRgcjqUJSQrb8Jd
UiGLFd27gjIVG2cZVLRosllU8ZpS4e8Np8Bls31+fO5GRhz6fpg28hwdpkMcQ3K4zj3Qzu1MtRU4
wcZ30MDzOtkz/woofqjQF6uG3eDpToe2nQhaRR0n795h4LNdSDBjcubWuK+kSPdhq77w3s/yxWPU
TBdxnEsEhL7gyK6SUNqV2V0wyP9fYBA1lG0hTXS/4H7qYt6q1bYkSB+F8iyGmByuQKBAgxW4P5nq
OFssMvyBpf44VnLLsCMbjefpzWg1YZEDyvOAOFhiAXoLRcqutaHmMUT3QJBgoWMrsDUSIfI0YPbs
VEEsvVEHQv7AqcihPN9qKDsR3F82Rrxg3hggW66dHn4WcjJlZTUID6fg4DTpqIDygcIdc+mKQfrX
PgKV57LVF988JxFpFPBG5qm3M/ZO6mpfd43/wzgjtnjvPzSRtlgCY9BjkEETO29DT36qg6FPgg9K
8aYa5xMh+6iKSbmXLk//OlFBFnjuFY/VNMy0Tc8xMgF/GkrY9sKxqTb+DnGdJOAUdMKR/yX+PZGO
uE8/uYvLo+nY5Ep9Y6jyZdLTFbzZBYBqZkJ/Qe61UU1N3oF9rWtcBfoDLpifKxS0K0WPw0NggIin
aFRQZh61hrs3mfaHXkQ1KUQXqiwWdZCKekZwMH+fvjH7zt5n8F5B++bPhN/WF5DGmNKNL5i/7YU2
M/uguRrxxhlQXnga/sb+T/1we3WpZ96bVixyrBNyMLgUWErwxADgjcll7L8McWM9cyp75LqKzyhy
2sRBjkY8n1TAWYHVnJPkCBuGv83DENGBU6c210LMBzdpuSkb+vMRz0cvOzOh1SGt7OcZovoBW8mc
ugQVUY1qaZ4Q9+8tgcTNkUS+3mia+UTe/vPMpebtWKAtGVIfFu+6Am+i7tYxIzl4COgnHibMkeje
PCx/IT7WTb4Y2I49F8jDjyliQiUw7BGhHnPRML7/kkAxrYy/15LpN5itQfIKVgi3iDNri4a3wY8g
0P1lSp7tkVwN8Naz8456PCB/w+w5BZOtRdqqVloW5PfPWddjSKbmqU7rT4QiF+vWODvy75weMBEt
ckw35X4O7TIbRyxnuk0gKhqO/DWuPfK0+9mTa2qMlSIOUr3GnV32jXba9JYrdjJJTObWKoR9wlKo
U7S6Dj5dubzWwssYJ+uBOHCUlJWN0o6h/zkNwcQLgXfEnt7Nz2id6bbRZIj1TewEsB5FAvG3sp9A
oPIDLUeg6eoZPVmQJN9V19MR0a3sF8wFVa+ivXG5hwom3dhCAlkIPwNpXXKXnsiiMUsjvmPGis9N
Beeb9vE77Kqt+w+Dz9xynX9yhOiP3vrFm+U7jwLx9330oEBep3lbxK5sGrcXyKDk1NXnpgrJli59
0mBWrgI1TTgm3sNfKwmtatGaUBUDH6/pTFOhOsYv5oqDJN8j9z2VQxRKYhOEQ8HoSYx99q/aSiFC
MevJXpKVFF4a549exHwgaqZBTc2tMzdFf2181x5OZvd3YkcqEMgAvriI87ONDusjval2OhfpKZtt
FdhRDvFDFe1W5X4gs6JYwTYt7gJG5ZGM+ChjU35ltzLrHeSPo9fv4ad9qFXilFZDXMAFk6bM/AL6
iux3zIbEPm1EDzsIclNA7xVb1pVO0C2x/J8vv6Vp+QhN5/Ciyp5KszOcLDoZDMZJHFhdcPF9rMuK
zmxoGBUrJeScLIyRRbiVRCbXb2g/T+MA9tLoaHPM6Tqw8OzRDDMd/y6IsbAQGy9cMkwEAAlXSScB
Utq0aYDGgtXjhgXFPkbWvojkY/IwOX0n7wXjH3DK1rjImUlAK7hJSBgkGgt/gsxLmyGgIawaJvQi
/78Txn68DACn51aiSeFz9Hki/qP97JoY0pxcAz8o00zXq/jfaJ33FBEqTGj87Hx6USODpNnD9GgC
L5/WwCgY7WAgkxC6qMzSVpgtpBsySgPsuUsw3kngttwc+mDkTpn1vtgWRcbTkTzlUZCyauXwyD46
mcQkTOv81YDNvSlq290R8M+9yMqSiHXA4x7hHHHmBu0cr/timxgP+lqBzGnEhXL/zOnltN/k9thH
Zw5CE48J2Pv7HiAEngcPJ5z9beX1Xx46UKZMzvPRKYeb7fAuDLQrQGVYeviVJ2QwSfBIK9SMdMNw
2FTz45jRABKWjiD17Ft+l3FW577jJj/8Tad6oKhCLmidaYEs34Rr15L4mNbOsSqxPqtAw8rbFkWv
G1URj1Ko+6IBHn6W9ywqjEVfuWfuzWnvAx8PH1is33RYNkGj6Nna59pPixMpWr8/bfYxJNhdEjGn
nkA4RkErr/rIqeEmnlbBrd70Emtw9XyQVF6IBp9v0QmHfLx3sqCeiaiZnjAMkOjASGmg93aAd+Wh
c4rirJWpMgO/5vCtXAexJZHozDZ8iSezCPl4ALAUUvOBMlV7STSvo5R8te7KZuaCCMpIczwWKzuP
FzI+y5kuBDkn4hmbGD6756bFXBprF2RJE3v41v5i90tlQFL+Am8ITUSLkHubwD1V2D3u793Ms6su
Wav7kMYZCxUtY+wTtI39UcO1hxSOBUhFEHpiCP1GMNrWDYx6nVbMdQPOG2dB8CXKvICumvCbpjux
aQwMgBIFsl1zF6e8z7r2mpyv3OyZH3MMnpEfCkcK+1T3c/0fc31pxXFOzXTbDQQQhiM0vrFf+PpE
NVcI/1c6DlA0Xh36jCpPNuySaL5a44PrxBCX+YUdaDGXo0GqfL68onELt5YoerMUg3Z+3qAdH3cd
awqssd6Dbv48btW20BRt8DSK1DI0bdgXe0SBnOYseDAn0kPX0/ER8Mn96fRzNBjSDYbsTm6bGhtd
yY+qaHuz9PaBT1dgIahDrIcLHShafY7s6btsDeqa3B4lOJdvIlBIwjDLSRtJfHJe8/av9Qtr3BfF
blnIgGmnPAtRRdYzye46ugUgrVur5NeGrd08gxlPFDohWK+8jEDq3SLKv88oJaPyW3H1IIgw1hwE
7meZMlHBcF8oAk0XTQp2l2CQF+UN+ZxiCupLV5i/cMaFS+UR4XoqWpYZlreKMlqOUpT+r+GroxG4
2LLaGny49y6SFSthMmU1NhiizCn+eZRfXkyFbJBw7EA4tIXa/m6PTr048lkAcl5opJ7xKEzLsgQQ
UV+6SlKzs02lryA32bF8x3jJFwn3V5drCpfNiE0qKDSuSsmz1hXM4SPqVmLOvCrFXgvuTaxRmo+i
S5OYHvpG7SK+G9CyUlIMpIbG1vBrO0+IMj3ug9T+RhLZpWFDMbCa7ePNGEGLJTflE3Fqg8NmpkIo
lYgnakhyVlWn5Qi3WVnBZrG00G4a78LsU4JgcaYPNF1yz4ykqHnXs9MEzzR2pIeAORpy81AiS1ZE
/3D74RsWg7zSU6geROnbCo2EH+/lifuhYkw9aBO4LQbDpfnWHzUA9AHgJzJ0zcqBSa4jGWY7/Jk5
nwY8wiEUFpcCNU2YCTKnicVOi2oM+kDeY5tqEovQOk+mLriA6XOJADnpHq7Zyf+H8TLTfqnu3OXK
mH2GTc59RNLDato8HtjM5IheJTIv97Phuv2MI1NN2B2xXiyuZGlLbXWwi+xfd1oUFmxMv2ejB3b1
rmW46HGmwhJqceMNnPZtDyuVVihkCBC9VFlPzEXeot+SE6sGBPU7qkCvCSXIxzq5R8MSdEc7DhRF
pR+y2An8gZfLSXMsqnF/VisTH2O3XlKsy1vaJSvoLSlJKD5Je/9xWfMUoQqt2d5idlRu2qAOT2yB
j0WtAbqRoOMaoUlUP6AuSz1yi1J44keFevfSO2qzH3ZjlugPMnpmzDAKuDxp1RRbxdqZCZ+LXB5t
pbxqrNObpEv/xLZbP4AxLLZm3zeEqsYI8sd7HA/MszKheXRl4W9RQ61w9wQ25CDEiz7IJlO7Mann
jVIdkft5QcPKGeW7JC/WYOySmwRvJ9Kk5BbCGcJiZ6vfv042gYOxIGNsDYrssHBXtckiz7r4hM5l
goJ+2HohgqzTsiT21a6IkMB5V9J3gfq8DVWe+YuvTQ15eB8153+v4NXfvaZRIDrW4Z+g+ZA2rN0h
gWn4zqLPQmWILcK6HfIH9r2FxrfCoGPJTmVIfkWwdRAVctmEbbTYNvZfYViz1k0ofWBITTDBmh4l
H7zwFMQgCp1yoBj5LtTaEL7WlfNpY/yghJLVz9ndcGdnqUzlbTPVbeezAEIEXhyIXmAWijiTfLlc
n3nbkC9rUP2EEqnLm1aCV8goE8a0epRpelen3xAA1zyhh7x024zceHcu1Pb0kyzcBQAs72z0qd21
iSLzoYm26eBFKm9ymMvat4y5/6vjouFbepJYttHAmmtdDfnmK1FbcwdMMJeFST2jfAXPfh9azWWs
3U8O4A+qST/vEENKq3BKahLTUKxAV98UFlkmJ1XNOXAOkJE39USQYMpXCdN/tCDmQ2XEFtGrk4VF
ET/191TNCx5/js84dYCl32/lhLAmDG0Cv92A8gXu4bKHR3ZUiw3Ob5twpAtowF7H2WcXM7v77C7Q
PcX3fqwFF5d+Y7zJj9dDZkQ+gp200Ja+9sFADi9P8hydGEsZpHNWCawcq+ZIHo90+0evS9KmBfhk
hxI40phWRkuFS+L8saGIuUi3lZiYJhJ7OYvEsOG2N89VuwQfUmfoJZuhTj+XurIkwaOCrmpf3ba9
AN9IHq3DX5Kcg3rnMh2GNvUGigA0rjpKtqIdmsg2DOiy86WXPuGaZEItgO0+sS6ZfaxV4AJpy3lZ
1k/0CX2FPWgaZ5snPQKwRk2qF42hB9Pg9N8+Utl7JFFrBVv8r/CqykrCXCxU+NauNx1Yc1BzVlvT
MzUrLRRhQZB7A3uEOmNGKr4zNb5KKXVem4n5hKFCUBtLHdWPN/sRp4XnTe7UrtH1WomKhHzcWVaS
B30NrlOe7XWokv2MvpkGGBq0hdXbWxA9ovjVHUHkIMkcwhkkNbb28dDXZ4UnQZvtOZc5k6qCU/Bd
qwnI0v30SUGnBUQcbyBkvTzq0rftBfg1eVw1qe5WXjwpBVR1kwkWUpGzw9iB6eZGLOiyRvE3bcXo
0D8yqZXSR1DXE80WvZq8Cd+pDug06XvLL1hyNWz1rq+QgKlU2+dYplmXRX7mkPTu8LRMGEQOmwSS
APMzCxOnDbQkURj4ShK/SJt98UUdVtDBYmBplhjD8NLIAyBIhcQdplAm1aStl2eH9LtZ5qe5muQL
L7sBwVufWAhBV/g7EJPvLifGXfqWiszK1Mxt2Ar3FcqQBWMERJcBpp000nusRcpmaY/HznntNF/K
Gk+jC6q5E7o03hoimZlRcsg7RRGDYH01KfsGOBmVl3iMZSUQ3fn2ntNviBITHVkzkbHFpoCHsUS9
58za7F8W3Vl3yOMN7QV2ZuUugQgY1ouJjBvOhHtowk77aLs1poCVZJjwtQdmCxLV1WOS4BaEjpzx
Ke176y5XUhyKhVVzCSAq34oUnWhS6NBL2tFaoEtoBSHKoV/eHvDlFs846fxgHRvr8DtAzYmePxa+
d9Q7l22baMsxB+pv1pOZEXYFAJEbc3QLBSMvRtzaPVrN7PoxU910sH/JzdBFg0tJw+RFCKPMSjv3
T5YsBm9tLgDaeAN2lvIeJIycMRRF5ZLuZBsExikk4drVFhDxoQiy5gR7jlp5YFjYT+QzU5iysnyB
PY8iEgETFuWAENq66gqsPskQJdkz5sZ+s7bEBQ5gO4eBJjAvpOewcf+kJsmtxc8oVmbedpzV3NXi
m64KLGKm8g+y6pihNX7raoUPPThv+7hZuDO20d5Z7itoAiHY5zIwneMd+UI28FGnt2CCwrgKP9iU
MFfgSJW4+OaCfrTxxFff9XJf54elHWAUzlEcuQ2E+PSLFWlNJEQH0dvH38NCA6X0NnB3w2MADm2U
kHk9gdgdnpKJXMhvcjd0ece57s9b11AWiLZZJbQOyHg5ykoYdvuSzAuaCs/UEr/zTL5WHlwZWkIb
RojdTViEXeysT2JwJcWLgE7Q+/h5eummibMy61a/ixkNzTl1XtGA7ZBuy6vkv7fznzFk+2DjUzPf
QSg6KZIJAHG8BnStIqoAFiCClztzG7BjX07CawtNtfe+eXoS06TrowBHTgT2rcK0CVvrryE0p9gy
/h5HF75xXUVEublNQX1exxgoeG12sD4qDhQQP5PEMjHfsVgtwu/ff+n2pOYnPaWyJOPW8dohUkRy
JrNKVWka6+7UEUIzCNTzTyUcJSfv2MSYDjZ3SHa14hhDVQfuOVTjOdWKipF73fXZBpV1tkDa163I
9ZsVaytvTXCUrTYAP5u8cRN3DpvCWTrRNQ6j7wv989gKWe97DHterSoxOCIoZuNs+1SdLlLPUJPU
TP0qj6wpV1CB4moc/0Ah7CAdJPnxoy13f/OtdogsVqdjji90+uD29Cf2BRyrP5xMPB1g21ERj1zI
MYsJhB8S141qvMT+Cm15mdWZ1IAIvuwJHzCZ2AjNHfsumjP4gdsaFOm7IGsVFwVnR3LwEiapL5DE
H6rWU4gNCsIdZu7d7yebWNt2AzLPSBIqzNhoHkGZ1PWIabFP4huVnBe7a68dy7lMkhlyW6sro9at
yG6q5KwJqfAukbcnThyjViJlaqS8NQa9BQCA855jNrdr8ZMigF6DlPTlpmVIlsu5guLHmjD/JvPk
dh7OtSpVQjYd1B3mmFcug/CUvXaZ5idT1SXjQv8wZdR/u8j0Px+6ptmLRNyqlwM0SmDLHHvfl4wT
YuDSLFDIK49IRA36pyDusGnnn+p9CH00skj7kgJLS2iBMEJufqXvNWUyurn5CZInyAUm1wDKnZyh
FtyxKW/aIN2NBfS9/6kNjBwgZXNXHjAa1qPB2Xen5s85CmcUtI/IG5bzRlb9IDwa9D+mQpEHVevc
9TFqF00CS+AwhWYsaL2hVDrff1S/WvoZSv+1mcG39+JdUrVqet6IQQnzG/gO2ZU1FrSI6R64SeOR
fX/szbAJbNOJbn8BbST2acj6UHmFzV/hxZm8ngcOjIGPkGoNYGlYKQdcPT0NtcooQlOy9QrCbaPF
sy9fxUls3QolP3qjAa5vTBcswNewU79zwFuB7zSDTs6Yz6lH04d9ASh3wNl9eQPJ1qQAJLGT4leC
KuQ00eoIOFSNPRKDMTmndyQsZFJ/0ESywrnmXeZybf2Pm2qD444WP1bZ5N6KnUelcaqUo1rQIvnT
kSMBJoFpKNZAkcSq5Sb2NHAzcs+0I4ZNp/YTBbGApO0Mnpu3PuN3lCBIljMEQFR+grcI800gik66
cg48mWmr20CN3I4ldpOAcfXDtYLFWCTWkCrl96RmqvtGADJY8NAd7Yvbbc4JHSI/MLX1zHwCYOsp
3h2Z8XWE7wNLw7HiSx0JaKvpdPCRbSEC33ZctYYML7K2bI7Pqq/UcaEVjIEH6ULKT6z/OSXwYy0p
KcdNbLMrzLSHA8bO0fQKPJZjoWVcjAcV6np4/C9/93rbSgm6XBnikCjkvDeJoVGnvmmF5d5hKOZn
N8c6irafORTD0mnOi0W9IRR5Jj7m2gp+tK52sjdHvI4jUZwm5soMLbbtLTtrC1SJDnMHbIfVQjVS
UeUNvdWssqf+o14xL3vdjJMfzyXb6SJ0r17XQSWa7Kjyid9ves397swnCaYIsstGAWgQYPKUz7oV
47CzDRqXX1iq8nf8WVHxNolUhUM+IlW1Tta3//AVcEMhfVHPyhfZ1Hge8ptBziX8YNIYIXJza60t
sIXBWenYsbWpW2eZ5R/XdalmDv5rq9yiUNKjoyMFWLVfnEirnktdBUC8igWYTdYKQjLaB3/Z4btw
nH9rRH6Z+6WLS80ouFKTGgm8HVeeywPhkVPAnVQMZykoIhQYSCLJ+jfuF2AUlgEfTrKd3XEmnJgm
bAmtXHfwcoOLID6vQqiDhYrBK1TnAbESHWX3c/lLtmBZPcqn8BV1Rqexc2DDO9wM1Zd0boZcOhae
DtUw0WNRpuG+nvb5y8MLfgVY0gyn67LGbIAZMmEHEKOqnfhBAWVYULQSsTDWDbA0WS1Ymzdtdwg0
mFvGlaiNhCf40OO2YTyv+xuz79mUHNY4/00DuKh8fLWetfEpFFIrrMUtFrR4h5uGsphwZ+sEsCp7
NXf2+gMvTqyegOoM6EnzKnCfHOJnUw649DWTJuj4Dk2ZbDJIg+crhd4BIe7ls4b9aCc5M9CaevTm
3S9QIYjSnGMuROn/WyKHdQn8T0P7NEKmhP5nbyb7l9XLh4JXiuFP/UELzq6yr1P5ac8Zu99ShNZ3
w9t64LI+XwcOSPV7/FrHk5rJJRuI+vF9xjtCYuCrtrVisZn/rN5b6znssCm3sF9UeCkm4HY1EWIi
7IfOfdoUFBGG6JxvayGVmRBFHP1DNk9XeVsg9zKICh7O2i/YNO9GvMhm82snvDBN6NFq/XJp+qlX
o/Wa3D29vgou4eGaWA9cOu2UQ3f2dpJgNUaAZQasFItlbxUoAJALOpJGDBSt6QweO/OA2gnkTE49
MBHwlh5XdF7qPAcPWNJWYpnYLfket3I+l5YZ2igaKLvbWRiZl475LAMm154vlxKojul5T4BABP/s
2hDSC1N1bUDmkBJUQ8dAht/s8tL4pOGnW+Nynh1Sy7XmoFxdCo6y2hdQ5BMQOFSibMS3WxKdDfSC
dqH0b3benfTUHHbJuy97FSnVwfqERV7Zg+IQXWcfewspWpTEjZt7LVwN7tm+Ol2H2pBmHvtvjZ52
791esdTSrKfPUY6LDGNuRjeBZqmNE4WXx2DYBq+wkGAhX/cQSVCEjuVRIsr1Shz/0QAiKmUjRNem
FVEsIQWAfp5Tl4DH7DwKDMSghdBUm6TsatcnWoE1D8E3PiynU808JV/JwWgL27tIY3UomUeRI/dG
/F422Lv/Q5y25hhskXiLfBbCk4DpW9+DPtB486gkflDq/TocdTCHY1cNHyKsOumc0O1s3jJS+2jh
87ijfL2Uw2f8IjPD/pHVNS32sVt0nyXT/KL2f6LQbUzP0NvO/Fuoe9qsYGy/E8P+QC9Gn0G+j6//
VevRvk/ce/wguvwBIikZ5R5GcqsOPYOhQzsge+wuiyNgGWMHdITMvEG2E/JXp+nTbhCVKQ9rKEIF
IVBS7semyW2dUYfNa+ta3721gZlTMACJWbYgA4n8ZiNanKkUolI4cISnDbRTDEdel5AvTo7/V5mv
LI3MsayeQuoua54aVefFa0Aq7Ko9wSYZReoLFHtUr9a10lA4QV0UTj7Vha8bgepOqHZ/K+gK4FPW
QOlPJmdr/XWuJmtpIOjq0MeGEi3R707Tu9eqz3+Pl/OCKo6H6GPtwTAm2af9nG++5/z1mUMfUgQP
onktFH456vWsCD53XGG97A608GjqLA534qC4MKXopq/5WVdpuGRdQtFg/fJ/BBdjJvR+3lExh08X
gtJ5kRyPeTpk9O0zMZdDaBr+AB1lWqq5pl2gCPx2KZYZuLnLyfx9zxNz5rTyZy+X4KrRmJvs6+ny
whr+EQr0iT4Qm1lbICAPypE2fsfXqBl2dPo4KwT8HaueT+UsJTWwxH1Npqz/wi7v1jUBYsm8heK/
nXbOAvdGeAQjYMDgpz5cuRZwzaL9FjvFRmHWv7TSF9JHwM6eBdmLZHBxGBdyn2K+9yXf+xYOAQl4
cJBYIQE5m2EBITEmxCdvTJpljlO3z1vMTid385d1FFP3gNvzw+PepHfSTAHBEBrPFijHkMwvSVog
wlEF4Lx+N57evrNCf/iOH0Uh1E0Hq5ZRZ0osM+zsxVoLsSqKHi6REJWV015tVSNPXJ+UIUkEFxAq
AFiNAcQDFdB3IIVfBBSmEk547wzABZ+a26BBZ6EBa5j72Vrt/rHSqnuDDFDNu9oRrQuaU2MOyCo/
j/oZ+Lh7Te9YS4+SKo1ClAzLa9d6iupO8ruNZ6Tf+t9QSTyN5kq+2cKXtBANb5lP8GrxqofroNMs
9gBbAS2o1frr7BFG0iQyBNhGnMSC8/CvT6ne96GYtNHIKLEUyAs/VrvofFn5gLgCkOJGCwuAk+qD
GiXucGZSQiYEtzge0teTRqq2O2WhFoisx87ZYZExjGFA06gJ3EsdbFzAsxRhweQ9kYAtlhDmZEwk
frzMoevDPsQ7M4/WuxfqtF7bNcr+4GaPxYeBnhAgK8ePuB7Gh+PGg10dE2Z5QWFpZZJ8MFAyYIHm
4MU2ne77ws2WE6RUTw1QZqhOeSBFEG+C/+fWlDkin6iKvspEviAuBUDiMEDWHBKClOpdNhpwhDsJ
U/tx4Vgfz+Ii4WW0f0Dr+EO93cPUkbHgEwHZpS9/odzBJM4f1WzaVp9Cg0VMvkhhwgvW9ilo6/Xq
Ik9Han3ax9GEKHUJLzUo7QyqHtGXZDXX+f/HtFQZ5pJftCORJqfzLMAXUbZQrFtR5R3zmUXVnFEP
N2lOsLylH3ZDKfyqMqzbtsYeBuVc250feQ4mMDE1diX48qq3wcu2MnQmCw6c83DR8GC78Fx4PF6i
c4G2xyOqSWfBg/EbUX8BKcrMW2ekUg+0pW/qe13WV7zOglgDSqTIPX/8jFPk+Cat6fe9tvQrHj2H
Em5j3VwOqQVgSuGhrY+Z0MP8rLtP1e+fOG3LoiF044FSqoYqjZ/uPl0pKVTYun3dtkO3u3Ama0FP
Np6zSkyp2pTH1/NVLzCL7ellnr0xMp91bMSmVPo78T/OYfQUbdK0gaaa5qgZmUD+bVfyu0vJfEke
f25hcEELvDAJz0P05lzdOWkVFLBr7KGpIS12tLL8sKVPqCav4VxVYv/wIXYKOUh5/4fJy9Ukd6B0
5TVhVK7eCQhT75+iMZggbV11nDLI7PPw8xkcLg5OFjiOc9QMP/lZRHB+C3osbsn5WKpZTwcwYK/1
F5kxEPSnIsatCThPIBzKvZvYH8sT3DUCLmLGxT28IuC7Nc3gM36ojBa/ztDkPABdJonAe45en4Pw
Sy+R+z38s1VEDge1O6xT+67SObwhDFlPYzdDdO1DcTa0EAfODuMjR3iXKTF6SOuH2WsmPX9X4tM3
pHG8/S/ASptkVVZaxYDTI2GuQW5O3m7nMSSYqBJyBRXRUjlKvvA6W/UHGG+Jp8k40DJWJiNzTYsd
70AsP24svm28qY3/RPA4MSo5k7WNdqrODy5SE/hyY4WJ/nkYq3F/gItz3qQCr3V4QD3vhjcS6IMo
7cqECfTtptEZ5OqEUNdM+lM01PGwwHe/ACowHFND9CpYrhQLVq2grws5cg2rf/atAhrPqBn5wdk2
WyQEtzEmAg6LNLQ0QurZtnGpiLqDz9MEhDsZF7KR2h5m+R6+aEHz6hQyAPrt9TvBvpFzlYqWPBcE
578dbsBKMpn/g77eVoOZ1n8BfWA6/X8acG5CwZ8+5j9phshIPxtDRAwVWgHKdw10VcTNIlAyRli0
hz+h1uVcQHECtYaGaPwPyNFI2qbiQi6mwsPNqWZj/FPrNyWxL2X5pFzxjEnwbptWjVD1sYWjwK26
rtTsAfTnaMgg5I68mnGXINV7+2ACldBNyJlRn9N/DrOh3x+FFD0WUeorfDEYO3XV/IGqPQ/Kf0SW
HN6K2EGDc4FwbDl5pvn8frT5IiSRk5IXMXFm/a7B8qU8qvPuZH05vf6NKUlD3/Flg4p+65BhgESl
v0Tx6BM/jfdlhEo6lV499IGdkxnIh7N5ZFHrR0LhUWloVhavhpQMYlsjuP+LTWmJy2cPQIEOklAd
89FkVrNdpT2TGCGQrjqHXLrlxG0dl1gR7K9IOAMUjClC0QM7QFy063EcJbGlDz5hUnnVnHFU8cqk
lOV5+Jkw+ocyOSgnMehQfctagSbSdYctZxH7Zc0Mt5HzMu8XTE/a/kK/WdQWLrQ73CCOUWqyHctS
kbpFLouGcV+/UDf5Bo7F2Fvu49iSMC7gJW0QLLfjj300mOJnmPuNYd+yx5IjLkAQCDr1tUowqbrx
MOW4Keh2aNwXtaaM+iAgmKQXLlonrIs188XIurrFKg+DuCuKYsUHB1x2urh6jroHIaf8V/TqYsAZ
f7X2DY4io66xBUDwpCu88b4wsrG/80Hw/QezyDm7GOz63UCORGEXPcy60YZxu4A5kMA84lWJRUV3
rRUKCtzN1fZOdPHphRj6V4895OTb8gF0Uy/VA3BILvnQePuGzmcu5/wKHnVwRPPEIOBhBn6STW4A
GSHGxw4h7V7I8dw9KOsfzFpyQKAJPvPOqvBYMM84caUTdOz+BEO2ErR9mrCCtRPP0BhknclsDdGb
h3I8Ob65IkqFwePx+MeLk6AEDxH8V0pUuU3zq4dWS5dKDNu/E4TC7NFTUaL0N1akp/xhCpaDgKw7
rJhhKWeAPeMGJ5gUC9o73LqjInNwL4lPJ4GvyA9ZkvFc/ttPavdM4JNAFKK1dyzY0iuESfUqg1W/
z/pZbN/sDcYSVGtGnQKpanyH2wTVXbnJpu2KkUCiq7h4vtT7iRZzG71bEJZagTVr4c56XsBTZwH3
ZpB7uwsHIkPBT/Rbhm7+Z/FJOmDPDVMhZyxh7oyZa360hgUi8UZVuf6nvimYB9PXj4QSPLFAcrzO
Q1/yxKgYUOzQbfRXKaI8S0lR91Lw1TGkFWjF8p9HlZjpQ8ZcIuGVZ4k0xYdULMj3LO6wKMVrSt/p
ZZHZ6IspoG1yqECaboObw675NIbQmQdRSaGDGxtvHDzV2vjSsY0Q5dD8RHvCdU6ih2RW3FzXcYjj
qQJNnjtJaRDlj2ZEIsD/0mu10ejx0WVWdToL2kIfUQkqjTswYCqZUr2pdUyQV0cq5chNuLDmvhFg
HaeYabMqgsFlvxKyzqZSUllPKOwV73UX9mdqUNirwVliVyUKXpOW6Et1Rn5ulyw9FFqn5VmFk0gF
8dviN6mZHHsdEALfWHh0hu4BfwIkf4jBg80E6yFg6ktKVd+IGP5Lkc80Ju3Ho0t2jeaNADtdlB8a
A6sGhcrV/NZDJHmBRHDDWU/2BLbvqb0xEgN9poOB5sPzjlcQ4UfNEIFGvU3/mA116edPuwTDsJYf
KpWLTbKik2E506BOVNjTlu66J53Dw0JOUL4FyB2syLtSkqGBlCaSe1+DVyh+0QPc1d7OkbiIi+sD
Ftg3bqI5wD54No/IxzlixpEGiRjfZHvkJ/tcGWnhuEWor7LvHjBw27m6kotYFDPvOXvX7MLrlC+C
vGD0WXoiFcGbpPy3INXEssfRns+S9ih0riwC8QxXL3aEz4mxEciQmnPO+a0E/M+2MRxR11R61bJC
mYL5P7WJfryeqwJ7B4rKM3jeWiKx1zrN19hkGYx547CR9x07JxW6y/AV5eFnrNrnNNLkvQzu5fkG
bpZiyw5lxTGc7RUdFeiBGsDp6M7Df3s4HfRNYArLWJpZACT0Dn2NjIHDLwZQoX8XWQTM/MYIwJsv
xDJBQd09ud10VYXPKkNB8+C+d4YKeK2zTufmZILyB9fPphGdsNcC/wkUwJRvDB7YFtMjV77utSVy
vhJbq/8RI6u0SwM9kZ/IUfEKT+D4Z2gK0Ir7FtfhY/UKHk9ixU3V2jBY2ByFQKcwPGab0eJSCf5F
9ld8HXmZOSA28MT/vgpG+zyiaEqPf2nrpe9w6iaF/FA/9IaFixCLLMSAefnxBH8T2EXHK263xLIs
XE3ipau0vrrn5hXvhpgFWLmuWRuzykLRdHNmEpT1/19g4lPg/MTlGMq8P65BgrzBTVyMvLubKF7m
dyhteQ/4a61x56i7B3F0RCUK/IlWcsrUCZ7VwLCpiC4oO0Vz1dzie8oyVl7l+rA1UctBUPlQuiUm
bDlpo10eZloy9NKB0qmtKdnY7UYTinnBmFfLo3LEl7OCfR9VizJticEeTyeEAAcCVsNUfun8CWTj
JaqqOj1bKubnjDrfrmOLxoyrw+OBK4fIZvIqR9XpliKDDgLn1FyF+GrOW1jr/DQDTt9KAi1fWz3V
S7FFLIsWJFlPX97GP0vKXYsNpA/9Zd++cX6IV8FYMu50ydecBc7SSgzRDLuwRNPB6D/AMW4of+su
CYhPnRwmmLBbSSSSgHaOfF02Zj2+E0UK+S61nkCJRQskJeKVZnaEOdrkw2kj/6yOwyNxW7T7o0er
R+rsJ4nJdCvkCapDQowqMJw6N0y9hdws3NnuQ3swuDJnyq0rAC7p7v1crvdyTfYqb7s8Y/RaK0xr
0Or+VfalrCFMu+Kkx5d22Q2EQFdy7Mfg/6b1VbDNTCDsb8dYPT6xpt2lExWFpYo0L5wAh8N1CYUS
aAqj8uYXqlAxTcmdAhk+sfFfEEmNb2663YUH0kOJOunv57TVDsOm+/2HgEBzzgF75uiaolgtvme9
Y9ugLj58nxg7aUjW6x9tofg0ADnPE0hGHQ0D6BI6gjBM8n0wfzpyC6LBGOgrq2BKNFq4LnMx0Xje
EKxfrG8T/m8os/HkCP8aDvrIeWrWb+/1gsmR62KB2L9HMo+NQOXLHaDmflEmT6/WnEKEh802QkBw
TGR9vjj8CpHEADR17/XmAq/mNoFyjJK2Ft+Lq7StTuxK/H2PV4rwjZ1uvB6DwR/4hAy3b65WUDxx
C5fTSPY/jQ6LXfAVntroNWMUGnoMTyOre0/R+YaKLljKzZFie00GNrJqNADdhLe2UxaqollBeFmh
LKtUEI4INdvagns8RDloyJgwO1SrH7g6WkOQg7lYwAyO1ngqTaBxYj/7oHTDzliDKBtcw/QU0GE1
flXtbMyOB82m6cR24NcbMhVvCukbwacRQn+2eaj3KXiFUFkA7dpSGziChhSTEsYFUVXpZ2/yqjZh
T0X3umDUteGhzqFASJEUVVsfX/TDjBF/M0pSxsBEeT7BJm4lY0Mmmx3ITa1Uj8trrZTeUphqYcnH
5c9E+v15pUIvVuG42CqO40xr0LLDx2oX0g5ILMNRCuYg3gZ0XVP6AFZWG2UIles+dMmXLnSiPNf/
O4dq9hFSDGEUhlXhsS05kfepLhyTorf6HUPE1XTfc6pMLIf94Jnd7xVugxvKyUdWK1A+3AA4Eqkl
1Scg34/AzPZEfniQ3y+XUaYDQhiKSDPcRqGpxcxE9KzxRkDv7q72lcK04g49VydXgSgf/OPImyRl
qey31pbSpOBtJYpH4qQ0OxuZCeglcEsCyVvsjKW8DnKYoFIwFDHZQG8hQGb8iKST7VFT067X54FG
coajaIn9kuaxhwK05q23ZxfZ48Lw5ZcVgX2i8omfpbhlSTq2yy5mH1oQ8DV2U6kN5rnpm3mr7/JJ
wULlAHIXFNTfiPhE5DcHaRqsaPf34zyuUJEg8EyNFce++AXEBH/EWBXARRPYfL8xwLslyauZGNYy
6DhfHogBhYVFfqp7kQbsrOcd71injue9KLqMo7S/PBs0opclntzABpkes9VmHUpoWpHsKALq4Cyw
P0Rrf+M9O6q0uv1ZnazfmDJGNFuoigZdZ0U3TKietVZj/2damJ8kpUwhLVGJiBg1MeIoh3lbKCxw
cSw5ULj3xR6UE5G2JdW73UELY5LWvto0pLV+3XAHmXo7IUy+dZ7Wz/D+6j71cUqM2f4sPu0neoQj
lk6vYWENJytgHjJr7CleEIU2qnGAtlNKN26hUIqy4dfWQ3Tkj6aQZU4gb2PG4M1gaWzU7ycfR01o
4mzxHrUJAlThobsVynBI7+BRg8e7WkM5zeYXyQidTDTiz4qGmfV6ePyspC4scRSxLyFLsHYGVqWb
3A8PYfXuw2pjpxFhT2kiAs545/DMYQfWTdBrgYTh/s2Bfeztw8V5ntGJ/xAJQdEff1bAwSoEb+IA
qvBGOd+FFGNxDO1l3UPy4u1nC5Xt5ijPhmaKsUWGmkUDWOa5ajcz2tV5R+K93/4Hkqhh3PtLWAnX
zjnRdyY/o9qDykYCIQEkJNXal0KiV1/vhOWcjfn56dVXbiyGvM1xrg365Nj0ideBe8tMIR0TfrvA
r8g8dPYMdbUcaLUWoOEJtAPPSMP/DcaP04EauTqu/E73+ARRoD3Zea0q3hyqgqycPeChDAUdFOLt
/fUXzUWe33PhxJSupRW9seoslBNzuL7AmX+fWyU+tv0gJANL8Encct5Mp/savypx2pTJMms3n51o
xn46B35jebz4CqLVOrMu9ZHTNt8i+qj96cJhZfstLeyq2n7M8v5agw1wOvSxAYT98qmwBF/22DuN
ryqkpy5Yi5SV6JKBGfOrqEvDYplZBjXp305xN+LZzapuNnoSR2ZA2An7y0rk+H/8hL+GWVfNXlHK
NMQhmu1M4R7XkiZ/oM52Q5nY4hPZFSDXqymC6yj+/iPx/uObaJ7J7wzOfyl4XULILKRSpGwrxfFB
wk+vrJ1c5uC7yuxcLkQJxDzjbYuqwFWcyUiyudSqQkMIB/4z/ZIuvdryoZPMXDLmMxuT8UFAQ+A+
kkvI1uQ/VidDTzTAO2mn6wRfFl86ZluXPqp6VaHVkm84dAniTJ/601IBg1ZNG9j0InE2R0AGWqnN
nEEHMQaLmQM1XRjuysDR/IOcXt32qHct6l6oQjOfcV2yqP7XCgmlwO9Ey4pqRGSWbh1EeXg13DQ+
zHU+XEy22v0ceDOGxx/UxhQv2LvDDQHYWaih70FEGLKzCpuQVrGdPHn67TySwd58Gs9Z91to3KLx
9ygYTwcFNk232oDj4Q7JmvAw0fJMnTk2lx6Sr5uOTFZwp4gamPlahZYJjKH2nrIU4uk19Uxz4Piu
akUZNyzopoIwCEEKpqQ2H+zNvBmbz/U3dLtwB/nzKCqyID9sj1Zb0vgPwh+xufLJq+xpoTnyxPhF
g105hizpW+DPkcfG8ub/+S6Yp3NqL5IFRFbA5QWqSDSuneG8JZr/2VNJ/7IQOlntaLOwDsmnNP/T
V42WjxgC/xji04poxNGMtAZe/XxNfoOCSGsiS07zDU+n2XF4A1xDeWIRkTmGJklB9GQ425IcL2nf
3GTU7jN4IdSQx6jf7SM4jNhqbZ6BQ6mOIy9Xr+hwJpz8sbaTrWfITfADZBUka8Jf5WsAnn/rQGFq
4D+JeAGbw4leHNba2VWymZ90uW9elFz7vhKdskUO3SWSu9CURJE254mP+qy7cg4YuY667suDvMPV
0TIMWD6NQFMmcaH09QLy6/qmCFRj9sLuMusRoAN7EtjIgfL/R1EaiR5eOcN8pzm3ujh9n73SpGLE
Koq6vOjh9YWVSRXNczXqPVj/ET+Mg4h6iSVpMArKeDOLUx0uhv+Q2uERLtDqpmGkug6bvmruW8h1
YOOrBQdlzCY5nUed89luv+mXIc01Lh1iJ2XI1/Dr4UJl3U3cPsqPQITIbRcPLLbbRDEQ+NjTfhD7
1eQxRDS1KtUCpbfa1WMPyubyFMLw9biOVfOrNklC/Ma0xmHzSopwu/KB2W7uIieJYQTY5Nvut23i
jcd9d9libPXFrGCibOx+JEstME9yF3ocCLPq9KWPOKxOHY4f8/NH8pRvPkBxv+yRlF5//4ptTswl
GWjTAkeBjGunc/Oo8hc5k9lTuJNNOreI+i7fvGqme0v28Pvt31WSjpWG1QPhJFmrH9fDShcW19oK
Bjgj8hvYUvwPGKc1rADHWAeU8fLeGRcmlcNNwPwiRMKXX0HhM+vBLfXZMGWRES27HzFjDP9Mc8Kl
dEBxy8sgpHyrb9KRaPNWGLJ+tcBc5RLPHgO70sIY4eN2uTX3LbL1JoCJAxC6UnDmOX8115mUmg1z
IHQHBrJs2qTZoXT9Gt2BSlv/VX9kpgf0TOaXRfie6ijyA4nmkCibK8tbuno7IcBRIHCXZQwITuaP
z0NZLrtyQoMuvJEg7Ds5sDcp7HXxco6AoCQWqO8izn3MHR9SoY6J7CBfwfq5p65zyDf4cnFnlHrq
VhbA2gLURFG7oj4PDzsOflbJ9XgEx+wDMLhCtFjyPQh8zsDZq3LkfwLu+KwvQeW4IEEOSBxgvLnd
XKdz2Dm3hYWRH3ciG8tIFvGC83A3pH+h6WoP+qa/YnjyGbkKZ6G+8Zl9tn5IS5gJbdXw77S6czEm
bfyKcZRVeh3QysYjsJXeTd5By1hOELb1GX2ZRaVD6ttNM90GFwazk/V8z1/hfhoQy8oHW2gOsL0k
ovkEfboX8JmjEtK4BTG9/mrJ+xsSnSLRruC+O3XQR0clRsPJYaSqbZMgtpnethueLKePpkmbb/dG
uSUIZfYqbWrzwoNZhx2GD99b8ANRC245qTiFYt/6hf9mhL2h9AYkpvDvEi7hwbLqbm6Y39ATFloI
O3ZkkYTsnnakaGKA0fr4xdVoGxaC/xirhmKmfFLoi2+pun+QPaLdJ2ILj/pf5DCaJgyHbE/lvVNm
RTjhXHZUhxJXXHJOlnOBlpM2avnuYrwqhwfSBksJ1KyWuZ5/uzm1faCk77WVGi6ffLqBx/GyqEnJ
CDB41z/vzYWGr23Jb7NXO/f71E2SKuN760TbLevI3Jo4GVYTBCJbOn5zGsZ8IyfYWlrhrliK1hA7
H6IGlk+vUvitul6y2mcajR1iDhu7SrGVD0dOG3PK8/ypQai4YmtgIeNQsnub2/sRJDjA8KSrW36n
jY/12ZZP5fvbtOPY8uPWK7b1DIf8gpwAmEvv041tn/Ii0eB7oO7l2/QF/n+LgJNnuHubtQMoviN5
U4PwcLC3WyORrFgcqVwFl4qgwW9RInH0tP10+f+7QdpSazH6LCdVMcuCJZS44sga4YTKSYYVjsli
u46S7VN46ISM1zhxsqxQrUknKErPqBUlSmSpbr9EJ6Df8/Klj8RMiUCiVxUXgxyHYgabGnr0y5/9
93VE9b377XCXuGTYDw8HiogAiaI9sOrtV2ed305ORtc80KaU5mEHrOgOR5Q69Jc/5YzT58Fuqeyl
3R6/tVOyJEmOtd3EKypp+MJPYcbvmMdiXR64Y8twp+YR4S86VO53psxkJ838NQvWeqhECsckpzZN
wSyWU/kHOXJ1eQq96LRGj/igcGV5YJfgi6PeqeZdZ2clv+ang9x8gEo5UvX/xx2LFiipEwBcWL4r
g4YeyI+ZTW29Kf/owIjk7Jp4xDm4uR66uc04brZQ1xsJzuIEUXj7opEbiiHilIpxReG27oCe0sMr
0odQiaI+dbfC7T6I3YncBCMJFg6grWxI9jlcvpixh9NJ/WD1pplZ4raExdvZfgx/XIdsm26jnngX
1mLZHTI3MZw8FA01KlQLmmHHCJpLuKkPBmqwu0+Qy1v8irCKcHiZ9grk0vTEBrk0w/9x0f1NJ2zL
ZnE2pfyyR+JvhT7itqfmBVICfQAirowFMoNIvp5rOXHlgL3OjFxGz2krdpWSHfhf+aqWyrPRcgw6
K7Qa8jj+ZRHP4UYVl8RBWY5l2GPiMlri99Mk9+rPE3K/ggpyDOn39RcDWtYKbEboNT/HVGDuwBFx
I59k8DUKuvk6fFpCsxBpM8dd6JVR1XN4Sk4Vww6ZY+7D9uTk9BOYCVG4tfAVJHrsEyk+I3RkiI1o
U+20XBXgnMG5h8j+MXSFgLSpazTd9+gJzmnAXr2Zhl/U4B0uxizbmYx0mANlyB9qffF23jZWM2FO
4rC4lj74zNyq2OhYgKa0kAR47SopXa+U/jvi0GU0wiSlNDrtmAsvcJWtzip2FFx7npFdRUQh0qS7
JwP+ghM5sIduUcSP1Ar47cVgtmt/jEhY2ifN0Fyw+Hr8vrY3yX4jb1rq9lhZQBJid98CM9axDRfN
6lpNg51PU8f/w5HIP3jLDj/SqqYwJr4buE1PYRk/sKe2UB5F2RMQLvR/qHn5g1zoi+b6Xstdn4sy
pUIDyQIVeEHZdamWwiam/8xm+anAanfkB/Ba0wiXc4tvuDEYOIg+QyDnauuhjk7YEngaAFwYAZMU
9HoItdAY2RLeGNKAd76tTy0mb4KeIVKXv2b32u81WkcttWYP1HHqE6ptDXTN4bfVdhuDMPXL9VU3
fMmOsq2VZVpXP5uKInFNrrktvmpcIcO6fxi1QVbu5BumgrZEYseNipoYikYd7xtMYmUhuIEE84MQ
vOXCojq4MUUdnke6KzBIs+fJ3c1d+FRKQ0+zLZy2ZN3XMZ4kMh7K5J+ij2LdTKuKHrCEAcYtm540
3JhFDCWDWr67D+sEXiZhTjHWBgtIJeQzQ6VqTP8Satev0i/XHAQlMSikGotLpkvWxY6+gjPnqCRY
nh9XpWKjO+mCZir9hwXZ0QQ+pRN3K/YqpYILYdTCCbwJAfWq9NjeSei1emwhasjQSiLM+Cc6bNCA
oygHuxkS2sfTO/02C8uZgEtXDHs4uv2TZE47L8uamzLjZZE+bCCUF599FNB4dhTFlEwjVkNnGfk4
5CLxbtA8Zg/Z95iEE26PBgNAt1gZAAx7T1x2eZDZ7rY/CM/6w6mXzzQuPw7HMamboyO3IhED7juc
3O6kV/0uDvq/sBIC7Kqp68lI5QLiAVOijXpvr6n5McrinAYuFovD7GCCV5LfXocHmd75PXogS3qG
/v5WEouiT2YmeCmvmNxh5ngGQOdE+Kgo8lbIw6eV4ne99vUgzkCUSiDSRt6+LpymEcjCjSK/jhLh
fliaeP6qRpBK5Gtu5gFxI7ye1Z/Yt+ywL/QhBT/fzWKDuUXUPM2KcFgFcjLsCqWyNhqR+ErHhZRM
18eVqfvmz7PnpHKriv0Wc7bEzA3ZuIQURMAOYUo9G1RcG8tpAZnHANr4gDsYitYBLRso7u3WtOx8
xOwecIakU40DlgyXShNqNFqsG3CRqqjN+zKsfh08rAOJ015N4Ihi6kXAM2BiGyJH9H4Jx9pj5fFQ
7sFUZlinsXjBstcqIFZEF4SI+T/dys5pclvtUBv4DVLClesa0RyonJ/4znD2rQerx1vCTIN+8/Ky
zkmE2ZbgyrZdSOkqU7S2sCW4xJBuUXw8RhISRghW8x66uw91LWHE/bfCdJ9622oDB4fxDuMLBSam
9szyJZ09NDmSSL+Q+ErMW3Or2ZNxn/4T2MKpM+92CBMtzcf1CjtSlEplvcDpkfgFxmjvx/Zog4U/
cGZkveZZPNzigzg00xtYHrP8COrb05IhbbF3oG2+uh1hzTDJNAPlkKLLN00+R++0vzK1WAEY53+I
gCaBgbIHJZ3kxkfwaGjDTkJrwMCoeWhBi+1C9491naGfbXpB7Jeb121M5f9B5QBWrwubHNIrNnsn
W3iI0cH2lZhbgSx0HUghQQzrfW/jMCxEIrAd4eA2M/3x8lw6iTrjO4YP+AK4XFbLu0gbtqJStGi9
/lWNpxv/BR8vVenD6WlT7nBp4ImbhLM5+E840z4qgBkWACKzuN2iC9MzWixuOS9zDH/huZ/cdt3u
+fVob29RWTHiyO/Bc2qoNGDOVndOUyIpfh0F1NNgLybcpLuPwl/74+Zw4jKGEPv4jVD+HCleReYD
jiKve2DQCSXL2frB18apAB7JBL0H7T/EkC32lLAodZoGqnrnwg7VJwDMIZXyNRlhzmkaINgqCzdD
Hldgc0Yri1qzIZcp593G5dxxG+NbtFPsfibQ+GwO2LIJFRx/KuaPZDmb7ntWbnJpMvaRRA79PCOA
PzMRWy5CLeN9dA2r1l6l0M7ykFjscLNgggIOlzWfkUJBapA87n4gh+wjF/POS097O0ImTBfugmg3
jVPVTO7OEN8SK8jGyPedjAAMKrddzXpbzcBT7MVKLXCA2tsX2n6IR0tmQJcauQQNc/cyraKqAThu
6RcqtGxaBuZ1hfyrBg0W8FRRn5tSpjMmKLnLTZvSx1XM22iqn8zQ8gUIfA9TsSq1nADwpsEHtw1E
g7zGbm4IG+D1lxx+LEsvqEWa+0CAzj3BV23H2mgUqXX89pYywB3JyMsdIJZZQMUFnSTL7Hc918h1
ooM3WJsOTecTMQu8tMiGgZbHZfl0EbKlB0175njzZNrwwvHF06gONJADpQI6KARU2FvCuOU8d5TT
X3L0mCyFuT0EI5qvE211coQwE0J+21XTIuOgnAhri6yadRqlIvT4vdrj+ZQQbH4aWRLdiTjBZH8n
PPF4MqMqrtriMvMZ19ljERHshyGx6TyrSmqcuYoLRI4ZlArmd4HSVBVZ4NUGNemvikyo3HuEzxma
YkkUcFCpGsGRsdEgpqmIM1hSsN1Yjelr2PG4rK2/AOH5jdxAp5YwvK3kFUHZLu3o9ZxsCbOMNrLs
HwExXF/VmmqU0LMjWDiWpTtXRNq/TRO0AfDmEzc1vej31yBYDtOOjh5qUI2e1JH+3fccvKyQ14f2
VbfqTU8TOJslk4UAITV846A9Wncb8ft3Nq7fc/tqYD8tIA6zmDS3grEnS2jh9Bn/WBRhUNmmSdmx
tnCrl6ofFnsDGcwnQqGTMN7DHKq0evZtdri2+yatJQUWbzBBLyEB6Ucy54X/QnUnk8++uqaZmlMz
0ixOybbeiIurweO+qg8I7YrjpvJxBuL3RGpO7ybcUFCKF1CGpUpddqRAu9GUs9Fn5B8XRIji8IB0
dIhRp0yuQYge/A+zByYCSRX0W8nragGr6YkEYZDflR120CpJ4Pi1OFrkHVlNLzNhQuvdmaUn8nry
WYXs+8lhYd14TBS0+aQ8pON4I74VjiWFUd7inhuhNUv79scaS1+2eC04lVxiRMAlhxJy5Oj02bSs
dvfONhhwO1Q6oENA/OppYnxh19SEZMGpKsyU+JoOxZO46mhdf2cziT8V6dL6n72B3dnONAUQhIu2
VehCMguwAhV0gZGPlDF46U1KXPs1cJon7JDLxJFyBR5NLh/2Fz/Kax2ihNglUnpongzUhnxPuA7y
V7QoebjhDd3SUeaImxjwJ+PouPhlcEfvsXA0yTilY5ZqA4GAjlm4OtU3sPeswmNzGFTo5Hqs5nuA
0FA+MuqMLvnkBrmCnAP39x8by6R0AJD6ikp2jlqNPJwUFrFJWGn7r03vwt+gTn+E/gqDdCoNu5Te
ZfKiLLziSOPJE5ZsuWPFE/hjtw7diu9VDgaOo8p7DECt48ahuIs6X6XITA9b4KPS/wpOCqf6CiKx
h5dCXV9F0Emj+Jf4prVdAIhmSIKcGdSAOapQPXIz7C3rpj1NTf7gY9bTnZCGfbY7YRRM5Qp3ASPJ
DJEx6kGguqTOdxHnjoJdxX/PgPww4ysvMxx359tKzHSnpzdbQCOdzNbbkuTZn51V0OQBXummX464
Bwb7jug3FBNY4DQxozxvrGYITZ3+H42pj+/1QWs94JhsjJlWVSbBaH2hJUWUpsE0RzaWCAxsyn+5
zLosWJa960a7DFbw95l5ZzFJPXxGslQV1mwhpDKK6iIfa9kbuRgwfgW9H4SMj/udHFR4G6yM7MQO
h+PINDE0mWGPeDvXl1bBWRRw0NIZOHio71acgMHlh0AtFvOsP32DOdHtkc4vkc1A9vxhIwUVDX9y
y0/16ulQ9p5ASdrieqjltv84ZQwgX7iIa1MHIRVkRriflouBAm97LlhM6gSVlPm2Jhc6sLi1zXMe
13+a//vlxXeYa2wtOCLx6la6MHczbMnv98MwvmpicW2WofgwjymWMz7S3t3hyjII5U/zy3X50XTL
XKcJk+8qknX6KBOFNPyG7IBKqtZmfihdl8Sgv9hpcO6JxGHkYdCyhTg+nAiAtnbBHKA/pMKlMCpB
Lx3TlWA0ehMEFb5sMkMqhiIk4KCJS8ujZdZK+OZaVagadFVoxLNJtMwkjahr7i+VwRMMnw/IeB0u
NBcO6ra/hqWA6QF+iGnEDm4vT3MJhn4b+zAl0rciRrGe2wykr70EWa7HH8PFMiE83KU1SytxIf0R
jUpoX8SvvyhsSGRyFnCbOkO/Qt0sPEbMTmM7l1TFJZgtfga8+ldiKVItn5b84y3OWXgtuJQKaqRK
fEia3HKFpACAzMS6QWWHcs4nuLUTSAT9ysnfxlZ2woParc0ICrhdF+I8dUugnMaQZ2LL4FZjgld3
2nFZm/kOVJLbkSLl/KxPbTo/474gLTo3/W6OKs1R25ldSqdoP7DS095mReidwozPytIpQpV2YCRJ
0g2pFaVtdXtnliyefQN5h5YGIpDNVSLROD80Bd9x0oW6yiLPcIJiUSFeoat0fxNsT6FtyG34+xVC
PjlGYOW3q1I6y30ajgQzlD3CTsivxRC8zDgEij9ycOvJkM/0qzNQ603mLL2Dd8phPkWXuTXi+Qvv
Hh9Zv3A1c8uKjPfGS2hpEVV2fRLzZkIn9/k+fumoEPm4YkMOejWDQwkcXEaZS3OHX4T7o5v3Z4Jz
JfmVN9NVj4m2el//MROnIOyq9AAYv0tqCg6rWTc3xul4kEYM0UdGvwJWjrAN9bXSri6aDmiSZQii
Ivl1yA/rFiLNkj0BfmDMZJetoSzHEA8UDJbHEGrNI5Lm/mOP2hm7mfBxvhjuhCIsbCweoR5+gGlZ
V2cS+ViwmDmYE3gw/s3JA/k3ZqqSAe2lPkwEiqVsrsHJN+OdkNDuQbd9aZCD29TbZVqfWWaf+k8I
Noj0DTK2D6PSKctR6LdNcTx5ukqwdN8De42tYXR9nN4V2w+gmbz3yY7zoj9MWa0AcIFgMu4up5jz
gEeOmOa6ubR097JF4rX7z8MB0KM7PlvBjdDO45nqmXmEqnF4IfRcIK8LplE36WP2iDWoIcCChDFJ
RcqqW9cozUz+cDvQmnIPgifeVhD051pnCq/aUbxYM2XkPeS0EiBaT4lQ6Brw28Y3BnLwNpW8KEXM
wFJ7jcSfh9/ZWpbFvkBKCpl6jqaUWDFJM+JFAig3gPOGsw6UbtO6O0z6+w4/UP0FPfFvk9ccKpjH
Wq+sDbw+3V0R1UVQFfucNJz8/I3pYsHYGsBUyZ/Vm6QUw6tf7wzJmKrkylGs7gYWfQkoLyIpYbjA
x39mThGq/W0Tr6pUdwkQQn4G8S8iLry4YBJ+pbS1R+9MCu0tilx1Hr/ykrwSemCFz39+8uIKv7k4
Vb3HHRfS/wZHdS1DPcrfjJjEKcDrChvBldiuiEPdrZFSweYiNxWUApFhMqgE60E81jJ1oeyF9fV5
DQfO4mIyftdFQMUs2G/tKt0Zh8hB2BTE64CsM/AW/aX99LmgiUgO8RqhSX5kIy1KXs1okogHFn7y
Vd0OOrmU/q2JeUvx4U/hnSfkmupqlzKm/c41DLPtZG2HPxdbiBTKRNzHVSmhh5Rti7jMEOF6e8BL
zH0OmaGgBcJBAqJXx9PVolIGsbzG9IzXDU+VJaXAIIq3xO0nn/eAfBwUG7U6eEVtjVOq2g6NyKzg
tXKQ0OYA8Bdswvo+1g3M/oou1qcxyAmShR+zVqTf8PgvhFaJylNDE3CV0Wf5Tjq2xIfPfKQwtPP7
169YuvGEROJHb02yEMpqeYDXjTKYHqguBCjsO0JpLrMWA0VdGlr5Mq0pgH+n2rYogncDJDjg5s7a
2lCNADD/oddCmsrmjd/7rq6fyHlR4anVRI8Jd6j21Or63g5aTVmMNb0E8pOuhbv9gvAsm3W5ey+Q
gUt9T3d+Ii6LsqrSdXnhh7RuhWeUAbXQc3SOdt1Hg17c/UDqVzwEgZen+8yp6/cdHsXWptUTkK1T
cxA/Ij0g2yt+fzmHedHt5p8WNVwI/rBcRPCGVs52oJpqx9glnK9XX4HmS7B23nWuh/5ahS0dSwng
72vPRspr+r8y1h/tKeAs+CrpTScmatQLK/bgGEKHgJpJ9SmZJIFX0sA8eY0JHlPnKZmC4/5WaBvL
kRDDa/zh8nkuofpltXciUX5Ef056IT6/U3XKwfL/liiO9MS/CRjTGyDrlq2l0v/A+L1CL+yLH87y
t41ALe07pOgm1dfXkf+h+YeQJcpkLG7KFwFRRQgsfDQ2B4TfRch3yp+AOQojZLwnbn5q7CS5yIGo
/EIB9NG1RfXxTGSI0iNE5fQg3kVmMsB0kpFbbUqUqTTngc8DTCEkG9qswTK48GK6UfDGWtwLjTYQ
bnEpF3R7IU8BS5S6mnZXcx7lnyy31xrrzhB18bWUYS85JXB7PJ3p/e//pXR64wFu5lLnHLHfUZbq
RzarDAjXSbHzr/jQnVyvxTcdl4bYAkLj0VLkW2MFkBoo93ysAAQi7Ql/h7VpPNxT2phGNi4VUrDT
ngC62i0mFddaBKXvz6sRqw1GlipHs1YNXBPcPivMJ7xI6T/yGxzLDU2KxbxvxN0qxz5BKnEIVCCZ
SS0Dh0uK1nbAX/ysNbvlmQZ8RMGTfCbIfrKq3Yl8PC7vfL8rOUf0wKwGWDmTctW0a07AhsLchQwt
MvwhvQSHmj3bfvTR+sNITNfVVxvESxV2/8mRvab2CwcrbbyaNN6ZpRiM9As8gvtkI2rAtGgi5Vz1
x97YCXaYbbMmSHxGlaG77cTQjiuhZ5uDdnHMJ6yKmiEEFX9WHwzvC+nmFXmv9knbpk0jQgYs2ilR
L0vsMM58lniIfVo/xNY8lZ1/CIyMkyREmr0rL1Roi+mGCe7CvWMWeuc5CUdbKw3h3PpJPrv0HY/X
s/x2t09cet9cgAONJ7PuPfNYpz9a/jr9vsOQpqsol9GrWIq/6BTzyi3ZlIxPtEUwgLaEfmcaoLsx
SByE1BRITRSTygFxGiHItwjF/AI2atj3QbZt/lb3yfO5792mIPyqdGlW5OEa7G7k9gz0+ClRUJ5W
5ngOKzp1nn7bZe4E4eugkVo648x0cFwhn5jmwVHxqHfyleabBsBTifJto5oPrsVkhO3RmvZB8gEp
XkLSCoXFvX4F7whpFz0QtjqoVBrY7Vvh8inWi5614URPA2T9A+Fg1GhqyUaBvbWkz6TQICNI8wly
sgCns3KQCKoOnKP+GLZyNFImQl00pRNO9OWfxGq14ylGzC7GB4B5b4CilO9N0yQxgkk1SuQQ9p19
9Id8h3LbcTI/2GE1aL3wnwvrHc3zfSZolRBsCY5MZuQOdR81hGKhZRjNQZXKM5nTqB8/IpmgiJ1O
2Pzilf6dtRhLGT6dRU5CBZ3SlIjFgT3JuIhxs29/yw2X445IwncFHG1Yc23RIcUonoUpoW5gdtd3
MW/09g1pMF2VqnYxn512xnnSuhlijCVYGsAyxUSH2hmianWuud0J4t/G6eh2w4bJvXXry2XKcHm+
BgJ/kVbH0kd/iOunlpT3qMWAnyalCgoI63TsZ4MGmfDmfhKqe1LlvY9EkF/4Zqomk5gYjhBnAJGX
bVPoeIven5MIIAd5sZ3uE8GXYyHgkYHyphncNFbyRCyUqRpEvrsGx5ewYsQrcBKkw1yvoKa0Uj1C
6NZyagQjNrrNeT4CGuoV/n8jRmMDGWVI3wSl96afQ+9jc2m1nVkfHh9jYtI605dlswHJHuaKBzzg
LA1n/SJZHqwWwXp5x9nIvz9cNSduLKk8Gnz9Di1Wn7puNLLgS7g5XGNNPPrC+Ph2zJmSoM90JJlH
9UpFFekUNhGnmcZ1acg5hihqXYki7VDTd42F/MM2Aw2etsPPRmVZtKEGY47JWj7VDTnRVu/x0onM
pKyZ0tJfX96CQoU6crYLCK46tuXTjv3OSwSREuFtnaaItbvEs8O0GnNaZXvOVhhtDS3mWmUbL90g
3nIiV0Pjm4dA6EjlKsqiFfqcQ0xt+gzCzuFwA1ir2eMgO5vyD1AY1ElEp60pzn2cSO08PzDTCIX0
Kp+Mjg7QFTKSp9afKphaX+zg08XQ8DCjyW5CHPvPm2WyScfDWdW9TheMIMkN9DVFoO448wG8pknP
OyXrB3iBdUtx/RIIAS5YMj8RminNRMTq4v5xRaCxqRzMZdFsB9gm6qXBSWKuUnqRogK9fweN6xLA
SY07f3l5qqBSG1TrFQ7rezH3UrQoG8MhDD7FqtbahMOeoRJWFSnYtdQI7oTetN/nXZ2c90/d6W8k
7G+B6o3jCa9jonTjWXTRUa7k8Z4RTD51LIi0r0QgfZy4KRu5FIakOQYqYQNZduzEYyOcSaTNJRjb
Rf1VPj3ZAZqXGjP5vBWGVq6MzmD56bYIqTI3wsWZrVPCIIRe9Bx16eKufowBbzH95T668PfBx0CK
ABXwOfzNUJfPCiuyt+4y9Z4i2IQBVoTFOGCP9n/pvi8RedzoqKYbVYDB4faA2BsEMXsry0vClFoy
HNSH3BE8Yq3AWiLu5DzyuCLPjmYbxUGgrWuhnnwJs9j2Fv4GLRHMM+meCMmijeOky6n5BztmdK6/
NsDT1udk2/EWDSgPxtuf1cym2CoxN23h5DnncqGGmbnSXTPJURXwhB0BvnazcZ/1BqJO0IKfFjxh
CgcEzZIzcDPgQ2OaPhWddC+qYS2PAm0db2LW5T6qb2IxXC5Op/dcasOmEOcUL9nCL0UGE7YhqqKE
/CFgF0I+LuSEv3rmV1rgDwsiej0uXTnWbmdxRkPYPsk5zxqc4hMN0f+H2xR7vWqDguwoZ6yyntoS
5SkNQT9kKtkJNdjnjqXlIATec3Aep4zdzS3dDYxAtLJ0U/ETEh0w4VbsfPC9JFqxz2ub6cwpYkCl
UelbmtsXSqHN0fLLxiFTqEB4WYU1qIACrPK2QjFla3KoTRvbJoEazKHPYgiv6o6bCm+yqXp3JT3y
YaFXSRu9xJBjzLE5aMpL86DjBgTG/95+ymesdT6jEQaOIAUX9+a1TkbaC3bzlzMI1VAWRkWEFWeD
fwZ897QCnP2Ajdp2j0XORIPGjSsTFRVOXKwUo3xZqZE5i5JRMbzrg/tvDgASesIrJNdBcTtt0VZa
jhU1pQqBtwt6tbXB5vzd4uoqzQ+2aB9JK6YmoZvnv8RAQaW/9ILgwBgEaBm+dSSX6bN1Q5Rt+bBb
8PXK9tfyK8u3CVOmaxjmPda8ipRiZc1ezDznEcKtiZc4psZV+a1MQSnCv2Bjr2Iyosnn4K3HWr0H
HZ4txzB4pPINGaHXnnzy7upG6K9N5Q3+LhjTgQMNBYpeWVV7BqKY9poWVo384k+V5Rrxw3Y5+a+q
0wBkL+aRHw+DrKk9wY46ivHUJDeynMAYfBo0AqQhpsMEhGt0oEQ5RY2JYZ61YM0+ot4VurR6j/Tk
elPBDpCO4Tw+HoGLm+gj3v9CABMgLXPUKQTitXmTk2NO5Rv537INc7/0DpNcbQBSeSzT2lkKjIjp
UlPO+Wvqnpa4eWFCnMMIz9MXLlgrdq1+2ANaS0bkmrcmPh9dPS7B1VRT3VRyvvHaH8NbXudHFWI7
emonSqp/xeYV5SdT3hyD9BMLrRxj9Wwb6ZsOan+CWbVYckesS2nuouXnnhRiuR1ntrGwuvh4x9dr
mAoWfG5RZNPfTRRORH5HBF67bBAniSn3/oE1PZLXuGH3oagd7UAIzScR5pkQYPsSJ4GszafRIvM7
cnHqBgY9z8IzCWyTOVf6/5xXSVFzwXv8U99SkkmCNju6ei4AChi5I1n5bBprP28N52bdZTaX3zc7
vdCbKdZHwc460gBT7QoSyWv547+uAjvl6uyQzJG/Br53oDXDB4JFNgz/hVGXYNyrvJ+fwxmGB/EX
jRQlgbree34s6m2j0qTxlBnOf5okCmEK3fa0Pj2BcWjbRGYQ2ceLh6Lv9YvEL/btsqjsYFaN7jtR
QpqSZkRhrZwlxO3itL953roE2kAom6n1DTRsvCvbacVbUQg6ySdPteonAnytoHGtS2+ITkr3F0nQ
AfnY9IrvhKYVJ4iQPDlMwBR/QOXOsW+kywNEcndRiC9EC/vbbyKIIY+KRNJMotV1sYxJoXPbsr4p
XuXxIp7YdXtuc1tK7mLwZw5g51u6hM4yPY5hfSDaAE56g2exaJBEKFbz3Cjc1qC7bUtt9pgXVS5R
3MzmPwALu8Hq9GAuqeYlg4iL9E26PBMq4PG7fJgOA7JXBsWuGz4gZrd4Jtm2JsgHgXd33yu62UJV
0xLTiw/XD+05sICKWs2QZJQgn+swg8EhMh7rCBWa5hs7suHeteHGCcDKi+RU/Xl/cTDnNwucvjTK
2P+Z6G3QaEzU4G2acAQyLzjSiFb5wxZscktKRhQ1DJhporODouzLGbV6FcD56q1Ljjl7KsPWcTW9
H+SirpFybO/yp7xi5BO9sm3e1jKOSNu6m8a9vVOWRCNsDxrYK1aAEJz1TLVN90mqxzbCsSWxhYV3
ftu6y5pb6e3D3QXr+S0g2gDT0AwEh1skl1H8JZbpTiqTll3lnuQmu12RuuF9Xompv7H9RunPN+J6
ExjCDU0IwRjdZTy8XR0cPaWX+IPMtZ5PBTGGLjmaV9RtP/M/FRwPOXik0hWSH4G+Ta4mZyw573vn
3gDgdD0uSpS3TqLKEKCf4ysWBB3bxF13EgCpmNNRg221lbwjl862N2Srp8rudWN+fq7OPpUaeKrW
tnRYXEsxvrL8AfFr2SC65QLUKS9/97m0qgLBDv+suw9s34EiJiIT4KMafIUvYQM4/rM1DwKZECry
mPDxiLdWBslrymL6WeEv9DB67cQUdCbZAr8aQRUDxPHhsoVunBAYtV+5BrgSM5He42030f7SIDmC
OsCv3EOg4kF4EX0kcO8plEkOjeSJ0UPVDyVVmS0RUzE3huyQdflHV7L64+RiGeUsvdZVMIhTDu79
vEtz3asC+2yU1Niq39mM5oJsbUw79BPjjpSTMDReC/GsWEhCx3mUQBu938+NXe/4vbt/ItOSYPL4
N5sNCvBb9HGUAq5HOPMwqhNqrt3xmyFcvydWWoO33qOnTCJTzDkwb5BW3uzurAnOMz+cLenB+ueR
lTNDEekILgxRxmPL/VmtNKVf2NZsOMO6/OUbqb9ZG1AGQSUDtg/6tTErb7GidFTV9ExXnu37KYrp
e65wuI64T9R87xUP3JMoJdTng62OYhOYNuDgCavQhkOeSKHn5QyltZsadOwRtYcobwh16oKKS0ox
Cx6N9Cu2YoFkNxSwJNuabjlwkBQKVbaI0xP8az5RX00s7wVVb0UY9fwRoSBloX4ddHZpweoFOM10
XtxVgW6tjTqdYCg72yVQK2K3RH+TRnuztU+3llhXbDWV+19SkZb1Qk98h+mMpWGwRc37ySmC/bdO
tkyIjCMsrgY/tpI3oJg4y0NlQ8heegMGNQpTbvUEDXCIoFIHbX7pxrEP6TX3TP9nwE3VLQGUH9CY
om+izqOlEt8qurlUXO9Ig+61GJyXJg6d/ylZiaH7sKMMgY0U8ybS3kcwiUBHTVFLeP+MXOQc3MYB
2m5bni0LvcUi/lPdlzzHd1xS36hRL4PjFCv93MLLSQmuU49dDEeB7X3VisW081rfDYURvAONhFnm
VAAOxGWNq3kn7WHaeJL7dSZiTaDUfMc3bsk24aR9Ua/BmYVF8estafK9WzJ0L/qYKxxeCkZd6ole
N54zWSC/STYbiHK/AJ+7v8cWDuG/EWr18+4Zcyeq+/PIquOYKqXQfIebugTp+JoEG2qiolEnNg+1
q0tmql4OH8rLpFv2YNKJwVOhhy7Uy1qsD2XxYTPRoA7D8OKVDhE8CjbtV7yDwn5x40saV2eN/Zr2
UJMW3F7hV2dwbel+77erv3X3Izqve/6uFFeQNZUd5zeSJGxIbqheYK8siu5Oz/9T5IgxQo13daRT
4RKnOded7Kcn4CLpLCZtEPcxQSnUcUDHFIIeMYZM5zTczbsnKznqlS7quPzfxGlZhnWVY7W3BC8A
4hlGMelXX0S2K9GJvxO2F+2yf1wMIqZn1NjP1qCiHBLBT/LSKv3IKpNj8KXCfzla8up24RttuJYT
E712hCAF82prKOvKiRY9BGRFivxzmQOjZU8X4JYmyiSxw47D70rhww+MP7EHeYRHAU2SSXR8DHLR
kQecdNfiGEt/Es7Uarpe02Qiu1qV4//VCD71h6rorsZJTM0wMmFMXched4pt0wSxxOKuAuAbaRiC
ayVdn0PKns0lxkP0S3/92iN9Rh7Y0Ppi59qPyF+Bf8hPnO7Zkn2Q7u+QrJkwjryITF2sDhExkQu1
M85+0Nt1FOCrkMqADb01OZbXWKLeiMSF2Teo/gtOtDZiKS0VaWzoUxW/gmkugrZWTbP7YtPzF/bQ
C1zf5tC3kgzxNYXaps1Fc+qj9CymakUvOKB8+FU0mzUvS+3GHeQm+2VMaQu1UhdspUBYjSeODPLg
jiHwub39Ru/G+QJr5pqJxl7CieqXCarxvCrG1IIx87z/qWcYAAOHvuINRbh8JU+t6Q5HK9abCkld
y6Doc04uj+E7BpomB7obvCBMcsaOEZoAHE399TEg+jbhqGpg4qsyLAFbK++N/xq7BeDaS+Zq+NLJ
tHX9Rwmm/y6FisC9BbgTS1bF+m/U1K1CV6ZwRbbmkPm9u17Aa29F2Q4nncjtslgAFi1+cJyrB8l8
XAbdHSK6PMWnWSJbGnLhes8xIfzoZXziBNMZzcbSpnuZCIdkJGDy+qDyE1DWWn6Imt7TCNs4GA2Y
cj8Dy99Y3CRklltnu2MyRjl1W4Z3uTIMZvkAwn7Cjbhe8dVcavoDgFQCqaSwK8DA2BhDWX6vjEFF
Xo4Eg6OfT5h6h0ZxM6vjE9Al5BzNIiGzCZ6cCUQNGTpd5Vxtt/bYJ1mo0f1ElNtyxPt+Qa6cb2FD
akV/MyKxwSYT2N/CybDmCsG7aOYkSBgITcWkQUVFktcb58QJqH6URY5nAnvFrnaBJJGTeQJO/Da3
c/cJx4I13CZDsastgeOdXC5GtLU93tfjY+NCTf5cuSxEmo1cOBxOyCa7ItiozSSepi8iw9JKhQAO
SfG1yVGirLEBShOPbWhhPmi5z3FRJdxL4H3PlVJxUmbmsV/DkrYMETqs7srvq2C14pXUcQYOr6kL
W6yx65BiV/dEz9gISdRN8j+4wNSFCIDeMC6NMpfsE20salM2sk83zVQ5bPkvnVmYFdR3k+MFKNe3
Jz+2EJIqYL9B49c6AWCVQYryHJ5d1sxHLeBGhY75VxlsldA/X/P/ii2+BV8EWrk+gd8SRi9Y/twT
zDtYyNVjd9ypqoQ7kuwNI9vjqudjAuMk00Xc6z7JEleNp33Kino+RrMX1RVH+814Inps0w9f8efz
pQuxZLLMIrwBhJ1YwD8763TmbNTwid6fIu/B1EB9EI7sTTF0V7B3NcCtz0nkIm+T1p+It38wWBlD
c1rV3xl7MJ5pqZQAQsaXsr72QYcvzto6Ci0ExY7obJ5OKaC3NaUAAJmNweHkGRVDz7QZBY7jmSsB
6NDxeUMVfSosyFOwuNi8JUKVuKsl9UgieTX06RM5iQXS7Wi2zHS7siEcnXySf9xv02foahbDO0g7
1ki3wbbHs3TTE7DuTchsOfaTAtwyYKSx4SbznzLK1uOVFUOhGoMB9CxWNpkhRZqjMjr6oxQZcH4U
9ZHVhRx86h4/5ZmuU+tEdkPCpybJ2fEqm++Nu1t/gagOnawT2L2ItbxmaoQZofGH4/aslHnjzukX
7LxaUa2f6j6IBeeG8rtNK8ShhozCd1PkCKoHGVtnvX60K8pjYh+N0mmIfNs1p/XTTy9eg+2x1q1j
koHLVQG3FWS+1Yawr5vtV7YZDSjWuqeFkBV5MZmD0RZJcU4WK1hf6BdtlQChCaLex9T3QKFtsKtX
y+BVrSCpBMs3Mq52VvRUnoPnicfDUZ+OI1l+03bBx3I/BCM77c1bd0TLAOkLlmD7lZ0PT+LHGpI8
SPWdCIPjxIPjXx+beCMtK7ss7NaGjA5woYqMMA65XmH8kEub++uEuR/BhsHxQ7yQhhGL33GXdQ2w
nKnPGp3CuKILAtkNBrZgKcHzYbmZSxLTUDZnbUP/rZJIgSi/oBiXhJ4fCZUhExy5+vnY/tPkGUoM
i+oAP/F3dEZmsTms3YXeAqndaEUMBo0GTZ+rL+ig1EuJhyuMkUI5iwcgCyUH6TrGiDhjvzrBXl6d
1lwXAhQOHVzCOhjN05fmD2W24DE1fI6DKciX6lQDdoh2yjfgBc63BVGb/HeHXBj+DPvSXHOp1mAD
Ga2r1M0+gVhWbD1/YX9+lcGPEM8Jg9EkFToY+TD8zm9Mfo/mn8tWtoLUoEb1lK5vpZOpSFCGvn6S
u/QH1mvdyf5J+Qz1XfINAjHbk1yFHbtOOtGO9rxFBMaQGBHmg66MhrTWtzLlwyd00TgaWarsBra1
ztQbhhwkk182roOLDVbT9yk6UkC9oPH2+jRi/vGzbu3ZlZXiWWQGbU/AX/DhVK9IS9BL4GElN1az
lelcu4Ju8LeH/5OyTN8CmoXfnnKZHyiRLeFFoGjntjFdDDNy+P+Q3U36OmrG/P++OTMgyvovE53P
LF3i2AG8th/FRu9J+r0e1y4aJWhORW7DqfJxQKEpTQHxkMfW64NlFsg4LaWzg3P1oZokFN7rZZNq
S3WU/uL5Cu6/isl6ndhm3Rur+DjJ1AxJbe9i53zOZNnRwBI22fqWSpQ+D2YrUi/Fd8zuIzSEsTcV
FVrs/tZ276/ggZJYdQ04umOa4Vk2A7+pswSaia5mGZt/8+bTB9BlPz4Q124DHhEnlYrTPHWC5st+
dSlKsAwOCAvvBoD6uSdwuCxezjTzJnfY8ftW07t4EoLmrbtLMy32RrtmcTDuw5b94h5TR9KPbn+D
A+QK49Mtxr8+ilFybGR4NhTM6zPh+Eq1e6OZFD8LxwzZwI3xX5pk2ECWJGq81PEw6AoLqIjwet5N
uhoInUO74VRzk23UjTLSUSTgaR4Qrr8xKdJEba7JECRpsnty1G90HTeCdh7+6OgZh9M5ohc92KFp
Y8G0vBp/f0ZBU8EPAVXOUwwIpl16faIX05rLBRKLqfx/IrqaP7B36vlvHlhVVUhoq7hWwHhJcFWz
emfutKZX8AuDWzP6fdqcrv0Zr/xQbyi2vaasCnFwKCG4kbEQfZeW8EeU5+mSGThpkO3V4ww1wAjt
sCVDYQMkrdgemb/ao0C7o0krLVSrAh4L3jggvCuzQMxRzZy+1jaSQGjdogIq1EUinD8XA40yXOqO
5/njOD/pXxtjieMVQkMtXfmvC3Jqke8prd46UqhKViTFwCUr7cVtkEmde5TZB3ZxT3c6OwA43zL0
WuZqobB2BHt+Ib2rSJ4tsrogQLy2LYdNlWgF1MpJ+9nPAeJF3ne8JIz5aV9fPZweLn7DRAAG8SZj
hM34WwHs78iVAjMB1hcYGD3bTu/K7uLoKFZ9ep3eErGrJSetCOjq/561P/2TltEq5zFE8iJg7spF
0NKj/UuOc2QJrhJy/GGCb2Jvj4siBixrySesJRslshk1Me7Tk2nd1rjIFmOfE4bdWNSPEZlWIwlN
hXVB9nYuMrolbv7+D4Y1yAfCsQzpYWyZOHMgPVa2o9lXHK+b2pXRn8a779QHV5qcStWFpp8P4cDK
woFDQKFLjRWha7yH3TZzisKGE8ojT5BA1r0PBoFk4fbezSg7yqG/VvxHg4FTAoycETGYB1/OdhD/
Zm8rVbz0Ok0Cd3jkVnaTRewv9ZokB4X2GtdmUuWMPurd+Kqkako9J3A7nnL0NcpaaGfzPyqNwaTG
gCvX3mJT6pFjxLWY7FqYLtIVX24Ibgzhtcuc+s+QEFprcJSPTfWY2oVw1QeDceFNkEjXmTKQrRvC
y9VM4agDhNJRb933Q/Q0xayCfSzhd+w92fLRZQhncJegngwkiV9VZN5OFmWR7RShxYMbn1f+cJPP
wKoL9VzpnuSpbDKORnsaPEt2xMFU8s+/B0bDqtB9dN05/f2YvG5X/P6YG+Xcpj3XI/9vXDXfffV0
SwESkKB+FPFK6M9K6WgMk+vGkBhSn86p3dkPL0GzAXajlSWWKtMt2xld5eeoEBWVu5oFpj0veAcO
IS43aOC0AGBoeP8wamaYqWw6FO++G9ASe1TQ3OU0u0va3QxiH3yBTUsKBPow31M2YpvBotvAXhLa
LBO6/7Pz7B1GUuI4rgkSdf2eJ4ualCfvrUe+V7D+nZ9svUEbNXZuumkLGiOG7EjSbkNaN0Cq8lTI
CcFt+Hif4aEDlaz7DE945dkC7UtJe/GcS/nBbNKNffC35B91Wq3SSNEUJK7dzqRYaBdN2eIKS+o1
0IkRZdYOUsBLeHHlZGL8Yfs/N0OHF2eKka+Bom4wLOWi5bb90fSft5sXt+/IxCVVUEpLr4fq7TJ5
hVTdthSwO5wEKJz9ab555luq2vdkXtm+zR1xpvryOP0jxySBQnN97QEWq+ToXuS50vB2zuO5pUJn
50B5m+Ls5CVtu0g3kNMeF4rSIkRUT0Eb+rlXpDdHJ7G65Bi+kEPikU/9hWj2+jc2Zu9MkMxnovzF
iSCdGgUtehxnreYHMHCBsLyKgSvx/SrVw8r6o8DxYPZ5+rVVKzNpmfCpmZZEhKR0DN5wWqMa/Hu2
0ixPzVi7xL/38nSBOoNI/mGgJyAzfJ/3x4dPc5MXrPUrTTpd6p3yBp8iW7PFULTbrh/NxYzOiCDD
qbVvDi099kwf004ZCrw63AQVhyYeA7UqwTBv8PfAWBbFVDyGcaQBH26PV5bpdXuXmXSFygs7YctF
6QiY5oOtsiBa0WJeB3NgFPPurKlwHeul5NXtyQKFNOzdTiie+Xrcb2E8SkAt83mFrrS25PiWaLUe
mJzEbU0EOVj1WFbYhn/QVNEL2sJac6YK/2LbrESWnZ+jspQMwaAZJbFYkUXLrzws9NN/gK4oHX6Y
m1FbxFNzdQhT9pLFIp1aRJTfQ3oseQQxFgpqJtl4VE1XQJm6r0nExfj9cZ33rkZgiPSFxEaOKKAq
rlwB/kK+U0zvVDizXfNWUUXnemQ5NYGhCvs7IW9OVkRWGI/GO8RZYoWrGO+giJYK/owTcxp1rT1S
MwAKKJ/RKQCHFQCXBwHIh6zywSPHQK/C6IkDP5qAAHSMJHiTFEk1RvmKTmgBN8iW1FT9/2ypEdHO
mVkjGtEaYa8Xz/vxS/+ZWqOmZzqafXsONevImR4Ll0Hn0Nwf1ElFLUI0+X4+v37k4IwSKKWxBOGi
xvttxWMq69mBcGPzmMZjy6BOLeMmerIs67X1y4itSCIGTZotZbSsCaFhex1SZ+s3pCtGvW9aDxiB
1Go0cbqAUC1XkchFfs/3elQIuqeL1wpVcWxIAktqCuBbqI29ifXk7TnGyVMsvwhCtIo0Ah1eGL4A
RR/HdrINQvLbzCghNQXNPtbWiMctHG2EiDe5UTDsr5b+dxJQ7PeoZK+oymI5/7ZP+MzVZhmrN9Hw
gwsywTFWjoGTHxFjPj5bBfXrcjnZmcTrb0oz2zwIRjrGc15FWZLMUcFNqDG2FoO+1kY6chjP3Vdx
S0XqCecExwYCmuhyGj6nYm7lFIQ1bkMv2NnpDfy51nTodTpEQ71Xr3nQTYux6aAgw235PFkQapWU
04tlOuXBnf74YhJRUieQmDSIAbLYHMYuLFXLTE/zRpNqfcRHUzMA2waKVr9PUrwmLmH7gThXSIMF
e6VGACJMtKG1bB0VtfEjsQipimgm3PA0o1V16ffgMUTFaMVVTanARWDPYF1a6xtttjTyAncXpJg4
qiur+xk0BCJ7KbaZeovqPP7nwucqFUXOtzIA6sILpUTPUaApGziZuNAKmS80BOxPFKLzr+527R7o
7vhBIUiu+SJNjuzN8XrSmxzif5KQgny5n9j3bbwYuexUWHm6Vg5w/cLn5PzPa3MW3e7KlSW1PFFO
xjZMuAhmOfIy9e/moeH/wTj3ZvJJivXRPy7OUeN2c0bgltL8N4x6Y5bKKzyy5f+BLy95nz38vZzv
GXBNCEq43VqtAxANAv3eS7EG5c9JLz0QyGdE4G/xplWEPHe28/EzKJPrApxJRKrsfWKe8xqXtPlb
SQIDOKNQlARFhyzCaRDH3r/fVFi5zLsMg2aKz4A/j1bfLtwKU3AqjCBPrCh5Mr4kE/8I52gk885A
p+B4eAld5Fe1XzYsEioF0tVlEvvvyk/DJuHkJ0cNVxydcoNpLPqEdZMMWAhbd2uyHIdZB3FijScO
eo46oQ6Ps7dfedSQGsY8WZb0B+m6SWWhk033u6KfEVyCPSrE56kurq4RQ9FmdG4GgrF+1Fr6Hvv7
dEvJYdFZfk8KBhcX3ANv/vNA+ctoWmuEu+LB3hy+z9H0qNILSLqd/msf5eh5XejpneId6cuNzuri
w9gzU4L1Fm1Ru+YFMl58Zndzs7sRIrvIzjEASwVlgV24LfQwUGZ8a8ODvg8FScQpdLTmroLUUrEL
4cs90mcHYreGFQPDhGQnG0OHf6yTRdRn731QDRexlX9F4AGw1AXCC8zfNINDwR2p3B/1CGgaqdCn
TqXXSdt5Vp72wLdV8uNlB0mnSLkmf8wfYImY4Fpg3hc83ox/hXbLS9vALfCPu4Jqw3nazabj+rLx
a/djze+rnbzKu/JGXD7igFJXifweKKCQcizc5D6oY06YFIuBHJolX/5lKLA/vh+yiXU7M4IIS1OW
ymmyF5tLtGZGc296L/D8vhGMVvfx1B1JCoq4tYYC+dTG4fqSq1JSb6ySjzVSIhvPn86lr9Y5MpsZ
a5dysAVIP/QnNbg2iB9S8yOByUBABnupcv97Vc1GFAUREhBymnWNWzuNilFCvPBXNhmYXfTSdFHA
Qq+OVWCXNBViA1ocaknc5jsK9x+3qw8BMHSUvABDKSyRipPvGzjqVXQzmyCcuO2LWo+luLuVCwzB
MByFuN/Nc6W/+xSWn/z0yAYDgDcxkgCYdwK+gykAXlcv3xyvyUtdzUmJ1dzJCgk3oeS5eTfAStNW
+ojMq7DKABtojoZKpp6Ude/BeK4UAtuOIUMcmCwMwICPUQz1K9PKwAGshbe/qkwX9Ib+0Xz0Cf8D
6r/URUpkeyTVwduo3yRk3UcV06v7gka9JWCWAb1gabyoHxvR5oodINoVVikUu+uxWxR0/GPTeriX
AWgjU2Ha3pQE64vUN8qNcpW7PWTETXSJxyur+931ofAYJ95ww5z+FTNi1jy6gtSk0qCK0VlgDcCg
QYXmQC0Edo9Z/N+3r4NwANKAj+Uw+VZaVbEnPu2gec8c+uQDJu3g83DVIE4T1UmPPxvd+JvF3pZI
ZOoktONEICUkP+Z2lrbzhOwU2Oe0VtZzzfKIvLx4E9C9uM8UfNFSI+tPnTVZBH/3hBPScs8QjADk
I3FqEvWZ8pQT0jBGwFIpMO0sxbPAJCfqLiX12a2zePuvAof2wBVfVDAxlWYCw7afny+GPJmyFJHV
9uoHOt5Mq0aSc7OLLQeo+emu2jZEwOWmWsdJd0k4rIG20ye77YWRnzIGiNcwOCi80xL0L2xQ7h8r
3v8nyhmKUtJ6zHL69zmdgfwhy/D/ARvxsn8xhnU6Zp738TXLEJZJNPN/EBsSTvId88cqzwNrFYPf
rEhOnEz8sHj5BOFQItj/NL/QS3/tywbMCuGLnEn33kQncY5JM3cPveoWPMKF16grVOVIq5y7Fi2Z
8hWkDCVthZVtrYg8iHkNbdAoyWwrs+PcgFXsBRXWz5iTKAJFhN/opPhHFbOJrzQKcDocgyWnnitG
XJLxulTCE2mFZbgzDH9EMUHcbaTPPCNGJ5XQ3o0mFiBDUEZQxEk9r1Ajucxnqv/MjM002S8Xqf/Y
N7ghLfduW+snUcYdF2CW/6g1ChTRZ8FwOQ3i2R6sIVhrecJDnnCzP5ig5KV/UQQOWkCVV0prk9v/
84Opp9Ynb3BtJJg0BP3hUUUsTUgRzboNxXdPA+KmJdeP2fHl3P3Yuditf3v7JDxGzGQ3rcHrKvC9
M6fCXgzn57xHG3JsQOzJNDW+m6hgeV2PHkQ3bZCer24j/9fH6s040EKnQAFwvPJ78elwplLU8XIW
Y6dszehrAYrZ5AJE2MY91sRfH29U5N5e0zpN3f47D+ypiSICYJMYINr0DSZSgO5+2ILcGd9w7RyO
ENFDBsH3h2+idt66lVSywnVytwh7ChWHY5uRr267rpvgF1gfxNYcjFe7Ehv/o9g7dlvzaO8Ib4Zh
NyxSkrg1XJKYtJTWsbA6GMpKhgFb/NJO8iJJDiOGCKAFhpg/AGoIHA4Aq/tyNR9StQSlWQVK6K+e
ne2L+SAOPAcMAQQousuwMsEslJ0MT8sxMROn0KAFIpL0vCbtzLTOw+AV3TX7NaTqW3C84Pb4uEhF
Dmh79FgT+Yh1u4SSlOlr0TcjRieqw9RSmMruqyzk/QZYySCC1LiRGN3SLNbw5KPZXgCij+aH1VS6
XxMOaupfmSEncbhJ4rAf/K4K3Oe0xnBZ1lXj2k3IYh06rGLG+DkeGe3BJwRKttGxS+WnlTxK6UxK
ehWDXdiaKvw/X9OzwATL3n1cigeXzoN7hWoqJbtYiK/uWTQ/UxglJXWt265Sv0F03v0wfLeP5I1y
zE8yIUM5XfxdKBMgJm+ZFr0/rFd1e+K2bskB3GAHuYLBb6yz0s9pcrBwWkIrur/ll0NhJCTzUirO
pgdGjQZxXQ9j4yNOok+zkNXGboBj358MF2i2IRCWhaxfVHiumXyq+rZHLCmaBVVpa7n2H4Sr/mIW
Orr1pj+IdfWE1CO2W2T9nNLNj/A6zXSDeBXm9mSTFPmDHxNZvH3D1R9zreBrLksbOf2UaRMHyKoa
BH09evtyV0/5aTjieWvuz90vBtGOwj5RlE2v46L47MecxbXgZOoST5JKnASQcTK0Wl6DAjfovctG
ru2I28t8kDfxpY+UUz9tqtq3W5+SX4Sn7ZJb8f5N6rQ0ZMcEMFu6hHfCWR2q1lLhmSQvawknVuD9
qgiy15e87RBcNqqU9uCNcSfg+h5/FGbwOSry4GxUah1zeFeJHDCVSYlTuchmSRB4+kStfcarNsqT
h/FRmpkg+SAtIEpTHoippaGk8FM2z+cTwXNmnh4NanJ1mv9itWESxWeETsQVOQVkuVWMCOSDdxkM
dhJbye2wI9fozZL0xnAShKH78bOxTHnL+c5nbpFP/0RSb4Qgv1eTHbaG/GzzqV89baLXMw7qGXuk
udrY29r2I7xN6nKCK0u4QXs+E6QPfk45fByhy+p48W+Vrl1Xfk+JYDfNNjRZDhk3fpzYDRW62GL9
lr4/TvTqrrmstspKGDLCT4YkVWx3VdvfSOBPqioMoXmjvlBU8uE9NAUB3Ke6ACA2s2/xy6gpuXzw
+ITJ/RdWcCavGtqWHhzZhYwxpfiMxe+ozv/VvKO2SV5xufpvfvdDXAFf4hkAx5nYzQiIB86TGNjl
DBhC4UxIMJmtFrglgPyAZsJefeZ2/rEI7dJ/vVGk6xVsZdLSxHl4h8IFjUZSnJHHfu1doFt8A1qi
tXBTcFjyJLXltESiIwbCmI6wiQYJaXQK8ZxmLEOtTepNwsGKklqDs+E2C0WD36yHkheiCV7gO6XR
Qq+TQjPpbEDHy1GwZLiikveeeCorUKB2vGm0b/MXrYXHE5NP7J5AcAcgK7OeUqm8lCyG3BigFcy8
RQfiR6tFx12ipNUtSFBg9JZBI/MmOkAI0lyZMjN+vYnoPnQ3NY5dkAiMQY0+Vovnfq3UfYb26tfz
NlXwmzjG/Y7QTHkvP4LTgm15acC0mPCiEzZqcybpUcxcTfvtr9qLutgCK0mhXi+0AcFb9mySmP7h
3+ZRmaorsGht2kFcs2YcKhocVs8LB9bEI2VUS4pN5RlMiRxLCEB66j2mqYLpNVByoYPS9NM+8bSw
7csg99ksKYg5AzcKdxfJ2vlKPmevNfNGLlRc8C5BzeKHNjfjeQ/2/9LFH9dIxJ5Pu88sS8bOACqc
uKGOeIVjeNccHeYHiAzhR1tVANxzEuG/SFXcTUT780QOmosKUJfX3KSDLQJ/zR7LtM01LptxZ9He
3PggGtF7iqlFI/YFT7pnUWCq/Hm18WNIqtBsy+ygnYxs0CV9T0XCRX59q31SRWo37oH/CsefX0U/
46IJUyZn+ah4pD7BYI0wFvL57qcs9k97hzBptH2NP+LSqQgmUzfcHJg16QZqIwOTUlJbKBPYjOf8
QFQHdmPd3debXoVpPbzfcx1OeVvMKUff/YTAFt1ID5ZRBPdGiJb8qV9TMgSBAwd0NjpyUuTWfDPd
zWf0wCsIvKIinexy0VAg9cZZE0TjMzTOxjxE1hrnvTS7fAMyMTbqcTF44TuoRcG8h1I9S7BsUThi
A4/xwibRQvDbP2xysNjlnIxWyfnXjJ8YtCEE12M2NqvtROFdbOWNAw1tQm8yx+Nc3fKOqHFVknFU
Zj8xN+yJKGA7K1YUNV/TtAr4i3N8W1CpYit9H/oTvCK+1UT5ZYj3jL6lIjvBbhgaJ72sLc0i493E
A0Nxs63G57ASLEy3Qavrqv2TkznjfHE2alkWebE0y3wDdrJqBJ69z/7dMnCn+TC/mI6eor9E/sQ8
rH4Crhw448qf+Hm6frPC4imu7qep5CeMrcshYmXLwvXU/dN8aZYxatlmZN8QIFiPvrA4eCEeuGYF
7YB8Al0TeW2+oZI6RQhC8O+ONK0CBQyJLbJLzhmTCLyt1g+ZjUrotbPp4Q5O3O1Dx59bObgf9VW9
ZWmmiZ+cRuuLRwCff5U4VDFe/PhiD04QDkqAnzJLlCbTHhdUAUW4tLWIRItY/W0vFoK/bE217OrP
A5g5jVE8GU14LC44dwL3qQREWFjI5AttTXLsl8fuRumTD2kNHBr5SF5juFMJ1Rf5KlJ49YdEaT37
BhYkACKUJyD1Kn5SvJiqHC4+jpwET3gVGYdwvCz/MxtRfGaYP0+yT6sXMPlRiVzc3H4WirZZr/YJ
AkavWfL7I4kfVE+FLZ0uSojPqFeQ2d2lFr0kB1QqMGgzmd4s+Bcbga6s9KC/RNi3i1V8vr+sA7kp
sXLYIdvg4FJzwuJXWJ10wTSEbGF88b6GCc6CIAkw+F+K+erGidiTDDvGoMTxOl4boMefwaPCOZbK
aOClfSiYbLdzbo3HV0GPZyWG3+uHeY2Z3d3fJLiESpbhBRSrIXCNfNnHZ3FVIA6p+zkBYRdEIXEN
H4E6CY3C8hh83ntS8n9vDH6mc8MxmekdbfSsAUbIzxmA6f19o99TJD9C2Yeu5qFJcngf2o5TfNpk
RPS9bO1u7BAXO3rELiSwcD3opjOtAbl1fmiOr9ieojxUtiUUDjBhFUS9xzrRsuwQNYWw0jQBkVWO
NnIml8sbVRI6QepYGCazAXzK3vlFqemmk77LUfUTtnJqSllKCqIJdh1pWKKCKXDptWcDepGV2Pk8
QWL5ZV3D8oFWrONUyqgnxyQrL275pc4m6GhHgLSjXTwzaB/Y0qU+VdK697N0IRjjwDb3ZfsQlOK+
ACGwnT3y3FVnvekXnBBGmMVG4zsQtcLykR8T0IvR56stZ6FKwNLp3kOKFh7F4q42lc9Ohst+QNgO
C1E4pa8jvUPlP6qlX0ZKJktFzyMpHMMwhNJ7HhQve5yfHuXLHL29ysY7q+AmFy+FEu+BehZpJzKD
gSQGJPdlDy8W7J77FxHdXShRgGCVFi9FxN6rx8VMnMj3bvFPNw07a6kK+ZU/C6+Oj77t/OGEOj5W
adsMPiwy4P09PXMByQOZ+aqiVZnKRudXcQSNxWVomG3gxik/EdXmHIhdHhzqloXudjHzSQoeTBAw
/0EJ+7n1lYh5p3i23TRzTD840d0hbudZ0FZMuShuWVXwwaEaXMQpVF01RYIqqrTTN9cdpK7zV2+J
Xzv+TvuIZabR7rjaKoj8LkbzU9dJzLBe1pV+1qw81zbp+7i6jOPEPd9IDRK4HUiSGvYAq2u8eg5l
YEmAJMiIzwBQ139Y4CYjPCwn/1ooQg8e0xJv8XX71DW8pk3O/CsVQLq6VIRxtXtgGPYWjbz9ysPw
u4ZEZHLSY8wmw1iltqRemWvBDgnHEHLwGjlqzZJK80PrsQ8V5vQYorzKATiHSv0/aMEE/GHYg0XD
tt8zFbO3TvPpFifZmu9poJr4cmEOEPieOqqfWVbppHuo9BLz37Vml7IJdpt9zCs8UT+vOzPLuc6Z
gPs4cT/eEsCCRdwt9Wq7bFzdXYTRsb970B1Yba38bTshFAiN8n+EIoAZEzQe2bsuBOCRXkVZDKnM
IGtScTIsmZHcXu3HGuQ0WMd6+ySSCcornRGRjwWnnMoOGncuUG87HOBQNKTwjyfOIWYYskZiMqhZ
NCcgLjV978GlUO534v8KHF6fABrJB0Np/LImerMkMug/tCVFVTGBfFFuvNHRSPIpVxobhY6TQNig
AWDT8qiADbqDLLZBjN9yTQfR/yLFto72imYT6WPleLEPEjFL54Tfje5+H+oYtW4AULME3CJZodRC
CeIDcQ2EAJjqmDq4XpYEHD6Yjb51zWraJHcXzDJJE8F7LqTvHelpD8oANlVi25HvvdD9qTffRlxo
bHcZHV7C71HMGJ7Hci4AWh0RvlyfHt1L5gnhpcuU91Bpap91pfHAPn9mbUGLdc5/yfcmJvDD7UmW
32XSdmVU/I8mM6ugcsrucS5YPlp6aYWsmkPwMsTlEhLyo8eAzP00t4Nhm1tYmQwDn9GXFrTGtBp/
pd1MaG8LAm+JyMizAsgZgXBmfmnoINurONlE83jbrB3kNhEkySDIDaVpHc9+6ngAbvoLaVrufJ/V
qhYoggQYmnY+CHzhTlm6xZ/tzQ0qeJCu0UcxAU7TEY41r5HmjRIUKGxbygPdsVc/6SaQIo+8ug1p
ljc36Brr8iC8Uf7v3ntapSDDm68BZznIvRRB+hRtASXKteczkh+r3RwzYEUfEkowrnGH+h1vN2ia
e4223rjRWDGlNUIoaNZdYyR0MZ9svaSZZT4XPsidUeiTVhbq/mPBz/z/cNnhC1vbYFQkhOUP/zvP
6X2ai8pNYRODkdPgx6chpQzVA0iIflwaTDOI+JV1a2Y78mn5FgDrlx8n7o0kBNdxZD7FZwkML6AO
fi38ttFP/NexE1CK9Emj6i8iI5TNSOQktjayS5JSP5oITFJvkHSkZFAwakNSf/IdtxedOfFhqwYK
dnRx1lssIgHOlv55/wrYqoCEnq4UBicPJ+n9kqfLwbcsVlLHj0sH7yL0h58aJxCOaXc23+XA6a/l
5LKkASWB6Q0SKHCAIH6AtWPKSuQDE9LiwFyWVXT+GjncrcnQsK2gZUAqY0H5tHyw8TFVKGZB+b+y
/Et3g5ival/GLQe8JM/HmiXK1iLVBRcHaFGcaBUzSRLTftBDiumDx7vohjyQc1tBW0s26GaRgAWc
7vFjOoeHevECIq5CNDZyzUdhfSgpV8JvnOAXi8Kfrxgy+Gstqca99aKOKNWgXwr8aOz4GzkdE+1k
4mkzmE8X97ohudmcwMf5xB74XE9XwCWDFrN2tyGF84gGzT6T3XErK7nKHNiQ1CkFz3PKqZm7T1/3
uN9aRjleOhxd//FLd54gZxTRttQjlhZKBcw3xL6+mg9DeJarVWtmT6n+oy3aPGyMjwKZTIEztuce
Ki0smNL4ldbQeO+Mu45JXiCk2F7xQsfNP6vNAlP5xKbVJCfg4Qot9qnyfZr/rRu2f2srMRqflKUd
8PSC7aoQSQJFg5CatkVdnOD5IhCz98/sd0yD66TlWxQkmhM7L5pahnZHKOO12We20JFGVOPoogEV
8ZpJNh7EHu9PQ1Mp8yDqkMoVPBQ8HfXgMsKlCgKn7sNhhv6GkFeW2oGe5LMuCVBsg5BzdfuW0x4T
JMgCHIxy719tPbRoHcw82hDLfQ6YbsvLWrTLWtpE/num3l+W0hGDRvcfyWfjQJtmH6Hs/tqIECXC
Tf28emlMekH27vzhC34nH0qxwv1DPDR2xYq8mv1YeOY92rFQYV6eE832Qw3yD4qEli1w0u3DQ22K
sSIHYAXy63MKwH27kSFJfzEXn5bEMpKIuqbirngnoTU9KYWAfZ+Qx5cjuKbk1791P5CJa4hh56Vy
4WOGuNS+OMiDOA4X29R/9lu0eNu2JA82TZBqL8AGPxik1AqAixygCaR8hqYhQzHwrzK4Ba6v5rsh
JvOo/wjAq6WROmNwX4AnFcZvjp1JfeClw4dSApmeBiDwzDwULim2afou0hPeqx8q1LdznTsjMDHS
ZucgagduDVdRHYrQnXc32JVUa7z2n+o/1Zvi/NYramIR82pu2WMH7xYo1enNO+z/MEwOEfofacP0
o1ZqzA6Yy5XOi7lDjNWUtMtw/oXghWi+ulimaKEJXQZjmVNXotpqch4rVHxjB1OPvlg7J3kZJ9bD
JHXwgmA2CVcl3U7i9oUgdrsDNlhuIqTGbRjJVi/szsl83BliZ3K1i9tH3z+muRCf0Mdo5paEXTXd
Qk5JAM15CJiGjPjmj68wk7AQpsmx0/iXFnTTbKPtgHv7U1215P7tiTuzgCcrpM7Eth58kiolbGfq
5QpME05toFeXFPdbsv7PriD03H1Dnz9HoTJ8WjfuznWL7SV9EA0PrhRCnav90ktp9tC2T6C3Kika
f/zxVBq0Oh4eDrwL9XIN+a0qTCzv9B2WP0lP7vL4KImkGNm7HDvY9w1qoCvoC21Wk04TBLcpF/b5
vzhNBBeoHCQ8p6JW42j06iE2604nFWCrc9ZAduvMmqu3OsGrGNcAVyp6qSBbON/lE4GE8i9SuGY2
AMCgZV2JAO4gcgKgM9bVgRI23CMeILn6tlqUhLRX5Pm2bvvV3jxukOdArf9uBUWyx5+WO9VD+B/x
r6Znt7/SqwVww270kHN6z8G2jGXEWrOPOg3PdqMXoElcYGHYOEA+QY61x0m6fn+q9JYiDA/d4I2e
17hMl/0TMFmpMSxGunw+cxY1BEQhBRwuZF+H0LL9iyChy+JzRVFWnBoWkyHi9NGBLYBWLlyqLwQC
WnOj/YZiWhrzcMg5L9YV2KmSAgV1SBZmQUYrQeLNL2l9Fj4glF4H6g+Pw48hHx6/4PBgEu7+Lm4G
gtSi2DD/XFvmsQGtGwCNu5B9OinMv7VEp3fWOZ1k1ottAjgozqgnHgr7t0L3DFxZHFQvLb49yocs
xFSkla/RL67fhoJ7HRojNOUV0GTLIK4vE8di/ri1AtKNE1L4dJqL+mD5ZgZNEzNNPvUhtCRAO61V
OTkedFgqMSJa+vDVKXG4aFUvppgDSsJDMcwxRfzgcZ3gfKzRLSPRHHycHBuEPdtqQ/5XbdQOsFZF
T+RsQLT7+o5bE60cw99MCDGQI8oumpTWQ2YgLNzmN28PznuYPs1Qt4hcjiAaS4eZjM8ydt1Lm/Gy
fsSA3SQpLqETaOl59qpyGDeQ0SVm9xpNXiqaBUq5F7aDVmfVN55hFgrAzFsXp0GIWEt5GBT0N79d
+dK2T3KyjWRJEY5pVWvDaQ6SMZqYuLoRJfhss2zTMZ2k5FERo1XlXAur+ZMZm1NdbBcaNsYXXwLN
PANWIiRWfxQZm8nMX9S0HTpLuPMSCqTUHZqTtN3LmuGYjxnFKgxDIH4zbD47LhGjQzCkU5qtqqYj
Hazn+38FzCuN/8t4ZfrfdHwMmo8n7EOiQ5r1neihu6GSnYkRtNrWHexEM+1hjuYcDCoYjj3Mz+qk
Hou2f3Dq5LO0DJO83kqtAfpc2LyFSGWXPqM1u4XbeddPpu8q1jN+IsmJIBpRQLGOkgeY9Foeg9jX
Jdz9yNzDe1ATLy+uEzoNyx4h0lBymGinC3AaVSRPjlKvpjbovhJdk8+Ng22xqLNkii9IBuHgzqNm
tdaOYyr0SdFeeBCCGZNuD65LLfLEO4qT3C854czJWI4ujJR0T13G+9Fu6yHX8pyZ3Jfzou0N79Hy
9PwUvV0Ohd8OH5jhgADSFi2cZbImLQyo44pzBg6Zn4pF41Dq5WhsH7zLWm8J/oVwONo6kGJwi1Wc
MCZsSZAQIozY5rIvkz24gixH8GPjx947upri2kbOo4Z6H3GDUcO51ffS1G/UWOVHCTxHrFqst0Wv
T6QOPAoX70eSG92edgVi1E9AJs7Si2x8C5SL4sA1f/89Ryh1Nv5FTmSmeAwYd1mDyK7v1jyv+MF9
/4654YcHwSzTFIZR+NBoxHEHQ6S7MRTdZzQ2OYOgLLQNTzchwb1xqb3aapHsF2PcIaUWld2RfaVr
YVStrvNqdZ1C1Q64fxqzWKQThOF8VH/6wGHc1EoMVVYJwGxfUdb7FzcN9rKcgcj+f/hQbOaOidHz
B9kWZjM6j5jrTJZSpONQCi+/mqrFPa2Q4PZmmrD6oqqgV+uJiw9AfXBYaySV9JTeuHes7sky6fkS
h+AewddJ0kD8WQGF3beXuzVuFzKCEbIrXGo8zZOl9yrclWfv1MZQbuguEVudDHpsHWG1kGyimTE3
0gNLQS8teDDXRZEz5H7pwN7TgkJ+hZywy9sFJoQ3CW8WD1LnR1k7jZvbWyMsBTr1HF6WpmQLdl38
mZ8H1ydNic0pkJvM5FWf3lGGt6KoCq54uZ61Ls0rwqE2znGvm4fErl6xCoqNmjREpN2BdO8iWlvp
FMnhSsb2NHrsy/b+ZiGLay06824BvEtnfhM6dMDeHgiGMAMjgEvziF84LBRTBUP7nmEkwQXPDcec
Zj4JhwcmsKceyQt+6QteMiBcC9YM+ygIgyXZWkafZ5o8oTqmN84mi75wVEesx4REdPdanHesgc8g
Idl3xXFNEYdJb43XTp9TPsirMXKDDjVLhycNcq8/uvCnRd3k77CRKie0cabz9u0tpPotU+22GAUA
d9UWY2em+/NNky8ycRwpaS3H5mv6bIj/oS3ZtgROjizFHVbZMAIHpFXpJ6sUJdnifKkYOv00ygj8
eOFGtCZkePDTnOP2eB7EObMjEumrl/gPkXRdAvnVDTdqYQjHAeWTiy7Lp8FMs/wYWU8p0YVmOCU/
ZNCrzojkh7Y+MiH1cHfqAlJQq/jlFojkVoof2gTZYeW709g44kn9hNI9gdGIlD3+pNKsz0dCBQ20
vjYDVKc8meSsmkyQTF28i3X4vmprqcceDrfCGdlc5YqHlZTF0AU24tQE55d6K7CEC53w2bEwQRMT
46ufJJQos2PuVUOSgGYd19X2j0TNHwF72I5IthBRAn35QjVJfA7U3qhV1z3EGlGPA+A8KVFcgfhN
SQ6BHefp8xSFWq0TwJX5FlX1yjR/S0s8zqDVXbEAdLvBEFpGiDly8Qxqc8J5ZGqpAEhqweXcFsHi
X36iO+Thk7CV4rm3upMwzwM76IftFGDRUI0Jw/xr+52gQqpGSfs/KmuAYTE7MUvfIdn+TU1Ozu1h
6jsR/u2qhdVOp7d/DQPmJSYs347BY6ZbrijsuldiaeGIfsTBvjiM2nMwVJjtx7EHpX5vbZlsgiWN
oR83w3qaqoIGMmLylyxQIGwRvuIKmEt9ajJMFbCw/XJgWTZ8D+hDjEgR56v5DiJHKjotrZKoGZ35
61cVP4wdoIPs0AFc2HwqgBdSy/WhJJBqqWNWDR1bHs6BShgbNi+nyVPzSeiz2dOQyVtOM7K5dMNb
9jIZJ9IUcGclgNB1Zzk1T4wzylYGQk/A0q0s3L/I6VA+XutwXtjL8aSa/DS72RlCzAvcp7K9sk5/
bR12qsvYY3GjcNY6afXUbzAO4e/New9XHiF7OVCh0oCkdVQaOTxozhg5Z4MfGTDgDLztGgj897DJ
7T7xrP3B58PMpsUvjcVQk41NS8LEKcgIVWpQkH5ThbjkUJQjdyHhmphgPXFZ6pQrvZtOL2HYEXCx
+Io+xdTjDy1kLasjtPgUnlvNBmx4V8MDoZYxvcl9hZXTuUpSvLao05vdLVSRPyKvObnw2PnfZST1
eGKCZhk8BR+gId96SlAH9XoPwffyrnGdGkKf9+mNtSMNkp4SN666naNUzOsxZp+b7SKTBGIRkZRM
bPCVNMh4udK2JbkkNOlGxCcqrdV9S5g8l1J/K7NbVcSRsNHNXLQPdexK6GSTj8rJeQZyC30MijB9
rQuVHGrPuFMruSdyOPSNNr8Gbx9j/qNQnw1zQlo0JGGKSXkUpD6S86XdtAylIqDumfaLhZI9S8QA
BSVRTPkxVzgTGRwLd74d5DGtqzdP7X36YHTovsTFHh+99haZMq00iaxqaPjMjEiYYsQrJiSk6PEM
s8UKYgDVdf1wqwJClAiHUyIRpsItUWK3zkiaBwa0YnaRVEqjvN9IPXY4vpCTh1u4myvYPrNqmLov
QI20BL5VAeM4Exlxi6SJYYOaUlD85naOxYeggtmtP5umzA0e4i3ErdbJsAfpD1ir5Z1uULUmTb1t
5cs3Xxk3BI+e00cd4OIU2oxWsp/lHLPWd6rd7JHcng13b9iszLXXzSUJfYGfpjWE/z1e8Mmusl4J
mlMOMeDDEPaOFFCEzmJddMQsxxLI482rVJBcKIQIjiYqWTCAjZsUVJkvnqK/U+ZIO32DlSawvrQi
bUdwh+vEErcFcK7dP45SAnTmj/F+iJOijPDl5PgOlTwjzHc4LD/jtsq5q/vO70rrLWbjiKt/QCNB
7LIoSRQ9kxbsR7ozaQKtZ5lISwi8mvJKim2np74a/af5dsWCXh6m1qlixplTBQYSIQ4oNAPmnVbK
IHUi7DJJZZn6r6ZBrelZzrJJqrTuD6YaQh8mdFmyHfEbj4hkmG4uiv/ClAmjZtNamUCKzXu1lGJ1
LotFhQ+2u2n9GboPXf9h6BgSyab8eFdzBoj8/tC1S7c0rkUZv1fympfxSd29RBn4sB3vtK54KwKt
WqJGczi5kGB6RJUlR4bspm4AyOiUBFHompgmZX3UvknJHpIdyVaaDPgrLC+cE1QKr1LLYK7qZxHC
3c5a6l+z8chRkWsQiS7/GD7EwbXS6t9Tj5mSTAJTC5Dl+3tsPFr0sx1sBLR2W3gEZ3/wZBBKruGv
9s4lLXH+99w5pDBFxyd80YHLue1JGA4CokQR/S/dN6o22fcy7GxJBXIYkpxP/kevqrJc/D19gDsK
MmGtMJ7XZ0NqrNrC/k0KKSHLsf9cS6Rn+TVkPx3IBhWSAllKfFMKWHyz3FSv186125zo5J7QuaaX
e+oFMU6fCa5j2dEaRcjy2VJ94pgCfn95hr2PnC1N8PVDNtwwiCs9fVYTNJDrDULPUJh4pq9pkurk
g+3qkV9vWJII2xQ0uoT3TLc+8FRso+sz4tSEW7oPfm0NY3kYII9DF35YAwfAF2PKUmMI2Y3Zw0AW
dNoan7CIpxXHbbqEKuBI1luRiJtuT6BmyWWEcZS6bTwy+AP3zIKtu8/Y7odBB+tTqH735qq1tjNS
HNRp+IuqH8zQsLOePzeARBEzofpXrFgB01qu6dYUdA2jc7UWLsYatV45jv9hszT9btJyyBdf56oF
piINrFf1JGh8eG6CzftmskPslg/GIZyJbAXKz06MkgIvzj3O6CrOZnwFtGA0/Jv2g5o/v1BfuY9t
mVbNB0dW1/AUEJHVjn6iDlnZq3FEfNxnTccj0D27Bz9aVxMP1vlu0LeAuOTmSxZB9jO8fr4l85Ex
6t1xYXDso+pe7eBWK3yDCygYHslT8NeC+MPsqqd0VBEqSlYS0B4SSf/3roVjtIrkOXq6FtKfW2DR
aTjZCTXgoh+DS0sCt5YTOgGVAftU/V4lXDbFc9du8czeaIpj0FXclkocLU+wnGi37rN3lZdXoxBb
W70O7ibyEQW63/qa1khVxkJAwC8WGowvO1UmKCXV03XUWDIrQO5xBB0AdL+eDxO3lK1CqIqbnT11
5X8aqkB644X1UEoKfQKcYmnENbFBPrYASnPEpC50qdaBefXe/WhScuy3MOT9o9vJdYupajgRREGH
cxalVQeArj20oPKz8LhqGZ58aNmwyLhNjCbsPpOKW22aG+bZvs1nUPgPrScBXwrOULRAmQPSLeyC
k2e5HLpIvXt3i+emiCOPhYuUMqdCHdUTTscBMRrf5Je+T0tjwv3Xd/TPGn/RyyFbTGCKOxah9yzY
ruesnAMzMPnL7Xoa6PG1wtbPETlLqe6zOoL3QMfln8gZ45bP4s4OmVq4hZi/iK8bmTqSniO0ne5b
1mPCg36MI0p974tZP6VYqavjmTeDNO31tO/IAJwq5KSCMK46duoL84k+SrYTIzfkitYWFUk8JkLo
ic4PFedNMo301Yrt0Xnp8QkrB6vpdnt5pq1/rZWlOqJv9myLj2CQfY0mWqwKBUpG/v21PRule9wt
YNfEo6DaL07OguhYwBBljkPmvyrHoXiYrs7TMgBlM5ZfLr+9Jq6beh1/YPfSFAPkeIRH6pSWyCCb
+WqvTWFdgzNK3Q3v6tuH+kGMYav98V8Gm2C4IwLkpsUC6qqYX5/DTvqJdV2089sQyqUuUWp5ljsE
6Wg3/h/H9hvxc/NmWLs+a3uVQNMuWlKPLt3ZD0TxCm/UiOpRfaySp4evX8dT71dVHBVtVUItCUzm
nVAL0q6XJee5XPAS0km6sgZsyF0ABmPUWKvuIcr5fBJRFf5wsBU93MQwB71dJJ3kAblf3+QpVkU5
4AE8QGtol6rxz0brXPf73+2xLmx2bzATlICCtxRiEehs5kHm8uuuAma5N34hh6Q0wbU/YClK8i59
plrOOxm3XHsh1z01fXNUqR3hJL8J6o3c8LywTYUrsV/FR1E9tm/ujPfrh2TLiiFIaGIB4XGIB+9B
2Y1OqhSu+BumpFy7gZ+/mAbAPq8ctnHxs9WuEwTosh00+A0dvHUwck++XFQ+FZbgodnz49t/obJI
tVsy9EQJkidte6nDBFpa4iAAxXuuPXLGocXjpG4t10aWkJ/BhZ4A5wzD/NYF/gm/dku7yNombhvE
u0TI9f1TlMCoBtVbntGQUpc1Gn5dGpfn2Ff/5bI9WqjdbP0tsRr/fL7jDMFMXxlpQWPrHqjmWn5q
G6PQc1MJSFHX9qKJE/jCaxhj1N/G16JJeNalM0kwxk8qDUebNXPNEIv+8O6UZuxEJpqC5UgFO+4E
z583G6EP/RTXqGehPOxgzGxz5Lz8inNnXjNE8vPKen3TvqQL5n4uRKbfZ29hynIDxJBfUaqicOSd
cX5gJsWN/31Pa7nm+GNRrHPJseyFJ0WNYoH4pFgZHfTlaohOCklFSl98YbG05RK3WyPmu08+3m0P
XzArTLPSm4EwndGDtcdBaG4Px7aEAhTyiwXY21gZEBkPTTS7ravOZr1k4AcTk3NQrmRh+uh4LNpy
nGZLx0mvc/C9CHtMBmdJ5STW/12VIdJLUqxbgQ8SfZ+vqLwfRoBwQvOUHkpmW0nbDaHZawH6LPEa
JC4tuL4jUBO38IU0hdqpwMz33WlA9mOLIbu94UbUyl4fQMWwhbdzCKo10011/iqVdoEPWD7TPjaR
RLdYmXp+w7bHkUlsKOS1oMlCODAkjSOYjFC9xz0M+PDEe2sDSg4zhOjo6Nf68Ummb+DfATut2zYy
BFJ1QdGAWQsI7mGaL6pTEGkG4DG1sOvngi9M2UjQh1QhaFuO3l9/xIYHAkOT+RcDAdSKM0MKftRG
JUUVQG5Tmc18HQN5iK/9kqZ50OVBxwJ7HWB1aY+p7T/lZ+0AWQNmqHutSpMMY0FGIblMCvlzovd6
Hxmmc7wdsZLGuJcPM8U7DURG93eiMhFT+Eh8CQVcb+jLumGiPPUhG/yhLcQ0f7x4f7DujSVTXeNQ
ZHzrYBawfy/KTtSmB6JBpT3schfm0w1TVzTCf/O/5axQ+C9cRahFdLZ/ylPL6YkLIIONITiruauJ
pjHYxhTpeyx8NuVdn/WpmhoQI8eB+vHmCze48g49suZviV5SuZTcX/xqlZj2mKfeCLfr1Vr4ogGk
zIVyzW4IIbNqYSH3uRckHXvenzA8BKoMt6e/gQPijkH55cNGh2bR7Hril6OHFlT83840SEDDQpPk
OQcmVFDcJkud26fo+txOgA/HUjxxCRbb31tisD3Z6SacqqGro4nscI1qbyFnsnhw2vAEQKiHjhdb
cvu/940I78vKlRQbUuOUGAIQvwBsfxsBr03flj5TFz5HCsNJDzw98bf8dLMJted7aeHDNeoLfW5F
8F4YXgbJsJSIH5qgJoh+T8TNKBraAhT2jTyEyAuyaHtPNv9MU3Ikp3dbwpifUhLLQdOkk+uvJcs4
CCn6PCUNobuXTk2W66mxw45wyAkMuAwWjjbKtZ1PH5TxuhCOrJnSiK4rl3qY1WsC5m857rgJ52Kj
EUULtR5V3z2Zrj2Vruy1EfPKvNSrUVKiN7oLrPB1H8vS28+13yiRvm/1VhBrupq1RZepvz23+eIM
b/Wyj5l+o+0V8f0/8B/mbU3sqF0fZpOc/Yq/ujVRE0a6jGkLOHJnBfVZsh3Q+I3nkyJ6CuNH4lnp
wMM4NpcNVOuSjLIgbnlmxNzWAqf5tbbKppxf5DzIG3gs74MsK7fkpTazpztlG5aVK3n0cTu6Kh3/
IWzqygk32lYJpXR72oxei4GFoDt2VEtcJNXp1Z3DlFIPYXCS0oEnKrZVYdBGJ3Y7/vv6PC9pXpmX
4Ol+OFM63vyErifkUax/iIDBMzAki3f1EFwDMQo445qHyRQB6+Huwyui1dRrE7Mnx9z9CZ8fSbhn
ii6I9HEf1vZys47De/3EGnEE7E1w1KxRSmHNisTKUkXp5KKRQSAK6Z7Riuax45oYKYuuatSOyQjZ
UmGrfM/0rJZS8c9ie20jPYidpzd8hkE8VCawMtpZ/CKOpmKLWFD9iEkVsO+OMZBoCq3B1Wu9tokp
UYIE22gVaZh0sGwm0HXxS2LtVk1JKGXnNwgNp3EOH3Na0RKDk6wtulIwb7VEIeG1gBWUS8izwD1K
EWL0oTLkkM5JvaN/3Y4NOU1AqYeN8+ZdjAOLWEuQN1if/P1l46djdMtW5mpgBBIwbqpNwWvCowui
Rx8Cg4dDkNvKh4i8qX34DuIBRZ85XdqcGpWWiYKXPrXO/xpYCgDtebwZTb4f/kMrIYxd/vXJcAaL
dcZBKotT4S5/su86MLLdINHwbHs/0MASvMz9E+oMUz0jwihi7lN0uZcOqTEnp6jMbBE/YEnmuBA7
As/flq2+A5Y5ejMbyxesMKdyepE7JMTW8SX11OxqTSzjhyso4COTXfhGXoU4so1wHyXX1kRVRwRF
PwbIIrqGLJkpA+9x05tgmDROqwV8XlCiRywbKBzjgs3TWidTbnsiESZdybJf3w9cXxRklCGcuhct
kbolz6N5SiFi374j4OMES2Tr0e+4qAWl5q0qCqmaIRQg0kxav4+bKvnfvJlxz8aQxBl+m2XmaBCr
8I0cxi9prj6eehZSXDn6tqIwCoj/u4XgvRIOHXFwre5ZeLZyRVmvL4Kela0LSETA9SiedhOB68Vs
1DAzy4pm4b8VMVyl9rsM/ORbKN3pWv+YVIhu48H8sJfRWWCxs8fIHmn85PUH1gcbLoFdSr/D4oTh
O0gL3ckWja2CZwqQwzFnn1a79B1lW3Kj1exdwFYPI2QLBGBFcj/m3WXG7P+aqzHsbbPuqiCN2hkJ
ZDOyfTmOMZtDdMQAkZ8m6Y2yi5y4zCoBtdTCQmWjUX82qB3s0bcq0NCnBkvcDAa9lHmR+Xml0wv7
QAK/zjW612Wg4Rsv3uPR4xF378u2BehbXvNxNib+c3c0Bq3pezNlSt1mDMnPagyJHfesT8YWaDDK
x+CoHFp2qc+ifyKialhQeO/fLPVE0GywGA7LHeeSHPOLpFcL27SxmqmLODvlt7slXMYsdk4GDLDa
FM8hs3Lv5AtEJNxuE5N0r8xu9/HAo8p1NioIpGgHgcJKFFyUeGi3HqxWm7eSGRXO4IMKJRzuH4Oo
6hCqN8by7FLAQbaQ5lPDChu1AuPG04pqUMfXwmqW7kaPnGxdarLGX0vRftFly3jzxkED80OLY7fX
3R2/RYhLM+J1lIACb8PP3/J7iknPBQYze9dWvaRshZ8xD+YbzWM9wZop5rftV8DY1UvFJkZXMhZP
I1Z42XGV5rYR2KKKrUfxN2QecesES0XzZfDxwHsReY0EZZFmCbpTfsl/bf/GiCS0i9g8HtEzlkEa
YEdcGTQYRHafZT04SvbuhJ1EC2iPOJQD6Q8U3LhXL9fUiMuzVZw3Ym6t+bMeewEkeH7W4R17Evh5
K1jKXDOO98z0BZOr1GBDUFQdD5q+Qm7GIyp0qVoNegywO5f9JejrOHFj6Vvw9/D5tCmQcXurBXU4
tB6SBvQ2SciL1UBTfk7dIJ8Yja1N7x8R8AFllqBDSMTXFGDmWXIi4d+/qTQtQM36Hbdw68ibPZBT
vuPHHY7OO52jLhy/tqzY2sLdU5PpDis9UhtxZTMDsf7t+oyVtjVDhaFUcgfE8DMApwiJWP9YBE2p
qRlmrdmfWL10hdxJEYvVPuCEKYEntMf3LiT/7D9q5nInl4i2/0mHfg7OkD1jFswehWobHNmc2+O+
1b9NgB7di7SxgLeJqM1fah6HRxIk36+AEin00kUIqrySZ40Vuf/eUZVHYtpXIqDtONWAtsbMNTq9
tEA2Hm7hSdhzttmorENjTgMvhh6md+kG9nxuonrjzvTZOVZYUmRvgbw2nd0lsbxEruXaUFJiSv/T
VzT4VCNLBBxcj52FXnf/fjDVp0AQFJxcRdFAvfKCheNouu+ISpbrUIhxedwko/+7KzkAaWoKQ+Ax
vOc5VYyGNHcY2LerGlTdEYca/mmXJBYQIGHAGgIWOmKspbOF8XhIeHMj8teJ6EbFBIMsd6JkZrTX
QJ1iQADUksBpJLqEhi4SvAzbFGSTvSqidJFYPpC6fL4R5H1KVW4EAlp0jpTTzkD7/Bd0Lc1CN9JE
GHtrNcgP9+4m1Zr8U7WlUaS7WxAthMHjKUGNyo+rH58itd5wLo9ewF7lbZf2a36cpxH2RYV/RuU/
ySkmaaL99vPZe92j8s4bYYum+kzob+4dGsSstrxJ+NA3c64yys8zBd54iSHPCg79JKfiyQ6HcuNn
NdlXw7/awuAkQJrlJD3+PMWZG6o8nToDtu8NwdSiIzF48Afo3mfUYgalcdAVb5+lPL3VQeLPODfv
cDxHw0klnOY7ujet9ZvxvGEutgTlaKVVQQPRuwHwFCy8RYLigwP33VzN9SvbJ3HFfQx0a1ryucX0
3cTT2JHPdWYdU+s9QImsnadsYxJVbfy7tA9++v4SgGzxwEP7/yEuTjVG5q405wQV1TvYjRBMoDMh
OTbwrXf/orqxIo2VeOTdiOPzoc4HXRj8za5kxdCij1/5xZaBJj09hF7tZyo3yPpBGfIx/PJBIAmf
+JkvSqo4qY1M7rzb1PHWcYOt1iqwYSevZIbaTuyvyyXwBQu4s5dkcCcaekvjqcmTbqpsYqZ1iywr
T+hLfp4bf7wtntZNC9eq7S1+hsFJAJQOoRzuT4tLwcKFfaMgpcs49tcs5FIHPASNhZpJWbRLvO4V
sp8MCYddGzhNPduZ1N+nMliYs+3S2mQN45LOIAWRpXlQVdgb9lfMpY915sTDAC6GhYO4igIz3hGb
BxCB3ZCzR9qSqbdzDgVMXXdo/mHwPmsVFj9HqalvBDPpJ6HD99gqxeKIqogPJNZZHJHURnotb+56
1ZULS4XmlJNEbMGNmtlrvNEis4b+8VO3ivSwFoibyPxanhh7e87cbFGi4rMnn4k94uo5V3f6JjOo
ix0ewm0fvt2TATIWMr6VEsDGJfHHwO1D4nelVR2ItRYf9qeMxNQL7TAFS/Che/Vk3qLEaSYyuyJU
sN2V+HhIOSrkUtazPitWzkXZJWRz+JgL+P/TGnc1Qcyf4vruGl/HgmHNFjcxpqdBRvR8BEv9b5WC
umlAACqKpAKj9wYbf02hxDBa2lPgYiAo4oY5Q7hOm8GytrJSKYBur6hoyCOz94Sh44f16ZlDL9fB
d24CcCc+gHASX+CuzD41GLUs1MjRts9RjdToDjAzLjJbuwEwNkPZ3GDqOopwAFKh4e6hrtkwACpn
nmaq3CH2CwJPHgVD9CBvvkiGGdiLlZbqFc8lb8fGA4iykDJrTigzMWvz3YO/SB09ViLG7d7CxXDt
HiWsSjXmqqzb5X9Zh1x4hYRlG/NfuYlU821X07NCNdlLPMk7PRf0SK0GiTmVr2ssgbTfE/pQXdEH
Jo8k5WKlI9jHNC2GDdU6GdzApcLchCOp5FnSwz6bH1D2at/HXkG3NJLtIqyY2K1HaE/vy7Nx/NCE
5XnwggShlgO+PKfzZL2UjQiuh8jr2DChdBEM+0cJ/HDpu9mR3s6kXAmLtbLodZaWqHRk0KNsj++P
g+ddc1wS+r0MEfiFSdWZUKpy/42iCpTIhnX209b46yguPdg06IJaIk/X4Yfj9TLyb1OQVAoRjWiJ
JlwrM337lDmFc7Ya52+al4pn62dmdENGd4d2T8KVzm97/TCUapiQxWXmd6ZEpEc0xAnVZ52Qyu/r
KrFMyt2xHF8C0qm4xZLY7CVzwd3DSHdjTlNU+IAySQhmfqZ97FWAN3FCOUp60dHSb4EK7/xdyMRp
1Y4m1HK1+Yegh9JCXTaE4g++8UgE/FScJla4ABilHhewRF1Qn+nQV7sgUOnfK+XVKUFyKExaxfPS
N+3RaXxHhJmBBemLjiTTqQOufVyZaMJ16/gA22XQlgA5rKzvqQwHVmusWdRqagS71JvR+pYZZnrf
l3R9aH/mp3UnYcEmbjnE4Gip8tfQKA20C9hxcfYumwp1Lx47hPVRGIGGmfNjMKzIpMNeOuUBrftI
/a7iagUAmnht5zDVpd+pRVvbxM3cftWU+nnwAPUWMRB6JiytYKtp1ccHqTsp9iwrLZyZnEak+hVz
vNde8jIeqkWuSqeY4GLPtt4u7rgijhQFIrHFgTbr9Q2se4rIlEJfQ8+F50S0/8gSSubPV5LT61lI
4fmhSdBlaLxWyo6Xp6A8U3KvGlKKimOQqzoiC6F6UZn6U4YgABeB07SP4+dtD0mToh3amPwCIG+/
Vl/c/WpJ7AHP5lSs9gMJKSu2BnA1Grmk+44M7TeM9rGIq8jABB8XpE/0zaoL17yYkhwqbCNFiNFv
IiJ0id7UQ3NZ++yRI3X0zdI93YOGpoLr6y5zo6YEEzy+UPm/nUKRrT5iMUHNW3+TvvkX+43CXljr
5vtaCaGd949kIRiNeTbwgxNZWnv3AE6G8yh2CNrpPJ5jk/PInpZehjtcM86bkM4+LkMWjR/WUyKc
pZDBtRfKsclItuUqHKTn7f7d0oeMzFb9vmTCynMZseZSsRcLk0BInVO79Wtp/PapRIQ1La0qOHTg
j9N6xnp2TBvLZgOZOtlHUwv8hPbuW1rGXpjB8MKurSv6r/XJ0mEbl++qjykQDgz/1t9pxgYnIra1
wgTs+bMttCc26MZpLM15NK1SpwXYqmA7JT4V2t/eEn5EBmjNrKQ+wzk0vSbM/392LKQRx/PPSgCM
fzB09NVjvoM4LUKx6xMk1jQW4vNfVO6tJxOzTYKoLAI9XLIN6Eh7ZnzUhjna5TBlw0xQRd3AHrFf
ZykBI38lb41Fd821FNwusFiQl7d0Kzh+VkicRtbhZ8gwQKZO0ZvsyZzfO/t185IU/mSQsfctzT1U
5WUR4i88h5LcsGWHHWBiPVs+DhB0gXhDmBMkjXVKmsyxtF3xx7aBKVdlIg4dEBCEMktQRFq6cAAq
wmI2tkpCtj8FagL1ZQDAChtfrc3yUYHJJ9IYFgQ0o8cYLxIKoGUgIz9eRIMb1Bx+VkQd3yQuXvyy
vzLf7e9bC5dUJD/b2ZZfsI/GCZkOLYIy1kh8cAHIh2kJ+9/HH0iv5juhjbUql4PaR0lIUbmmRNrS
BwoGO5cmb070BIcUPiPRoRonUDfrNgSgY1fsU8tqSf1eZeTpCse4mh6B9FaC/8KwdSVTnFh+8fMg
Zo7DIzrsExJt+ePihtDqq7WVpu2vBoi3H1qtY/qJNiMYpcPBWco3U3dUbuGlwFXjEHPUgMlHem16
/JXphOTQdatn1Msy9BHccGKxg1ncVPIUdnxEwhNA28+DonuApcSuUh4W1a46y2z4vjM31dbEzNWq
zBhkZ4lz1OF/fEApPrOYI1vpOsjCMT/1j6dCeDNxg+0eGdImu8i+mwg7C9g/gPGlrz9uAzh2omyp
vlGUB+Kd4UlhlqTq6SvJELZD+zn6M7/FaCD/GU4utdoC3s7IzEwyzybEs+mJ31gVwPtjpGWsSMEp
vBdVa/IVP10rKJgT6oR90U6lJ7A5UF4Kc6LZY1TgBqm2Zr7WkhO6AGhWkQNv02D14IajD6I1o2xB
aMoWfqyVdfIgAjG7IVHKvFUmBF7UieaxBVY1E4ZcTWVLpK5BIoyM2lo//WcR+CJdduwALrwgSNUX
6eQOg7eYPQOn6b6qDQOjOa3vWwC+KKS9ei9A+WSmW0u33XYyLTVXPZ6EW0W2a7suYdnGHP/1o6lq
4wgUDwJz+Rv29Y41FzbOuSWsfK6r3LxIj8e9erz4cxab0uHZh/WAUYdF8yWBSsuOJOVasuvPW5mf
egfNaHoS3gn0IyYyoeb+Rj3y9Jf/LzHoCArrO86lkdwqNHAzSpTRT08QBC0mlyvzP725mp3mMxuJ
92LDBR8TyuqlRy+/HcTdsXuwVHb4CZvlNmqGxGvBOMBaSohNvXZA8Nv4WVakT/qW/X94iqtR5M9M
K9GFLBRYC6ahJJO+DcRjGgineP/FnxxgpEa+DKP7pnb7Wh6lrDWGMtaE+lwXVsgiJBlangaRfnnH
S33MNPFJlrurRmS/hhO3ossaXwJrSp9aYVFl4fiUktLWNmPop7IKsMm3OHiUWRkNdZA7QxJhj+E6
beFyqjsdWHJ5SRbHVTxWSzYlBG/3zTkIc8l0x+bSZ43WSM9lMFeG2YoTi8kX09mkAeq7vdUFf9u8
puDg1ZgusipBJ2GkWlh3qKRmEdwOyfIdYrXgrV2mnYyFgaITY3+QolSMhI6AU/UMV3o7/OGfFX6F
7KHP8slvdLblrNbB3L1L9xh1tePQtJWGiXSlr7FqIQaQZRlHpWSdlrUfIPieIVPGB7ZobAcpNJFr
zAC30F0NrxYEfFwb98R9XUBqUkI81gDN+JzIh+/QkieT8fnk3P5UnRYXNBA7OaKI/9eUU4IPVVgZ
0lOG5jL5OtaCO3x3icDU/W1VkSjC5fLyu36xKIhISet//hrghQgclTtUZnb5hvQx4d/75p+rNV+q
rks+wHDsTDBXozPgfBitz8yfmpOjsAZsbi/Jffb0xd71jCx7DTDtb3au1boTUNt9itqwzqy5farB
WSpP+TkyJ3/w5BXKWUYxBOdtAR9KUbLxgn4btj6L2/XFtA5smQQmyW592+CpiQvcg+gZt5/bJH4E
+ljigpikWsGYuH7u/VyJTWcVtBBTfTzeesDcTKtgzIQck0LnoL2Z9z+Z8lvpM3JkKG4lWcsrzmJ0
eHFff0Kz9ThByi+e0EYBxBeY+KMVoFflc3j66L9daMcWEJWgv6D/hekc3K2L4lvIvOnCL+HrU4ky
saFG+Y9ACqka7xLHyDVD6hHoI5fKVkIGY5ZjWSFBsgXqsyJscWwJ2iJFWgI169Imnj93WVCCmCoS
p6XOOw1IUqrjUToxG0ydAa559VEqEItTFYR9vJgJxAjIEu8HT54rIHnGOAddBaD5PDSw6/8NSdxJ
/y0yKIgZMjwJn/le9vak5wJJLfi21ydqVk56/KAIGZe3HYy/oGQcPr7IKsZGSO/1LZdNUOCX1rPm
VXvolBBUsPKYVFowgMFT7SrYKRj0/zWvPkSZmLRPtSgCSFUJfJHfRLzcdAvprg6mwjdgmVJtaXoe
tmVfVfLn4sVJvCjOe0kqnrGExCL/lOqCwRBU2qH1v54pa06CW8ORIq2iLMtgCTrYBLKBKjq05VWh
kKZoYgNtCLvBI6c9avZ7UMYcwP8bVsXd6ncung4jE87ANJxNnzI8oJ6vSGiZxs80OZYMxeDB7FkR
g0FlarfV/iLcbI8CBObC0LLnMKN5MmB5YF7K7oGupkdWh9fvb4ZCK3RWsf50YWlz9iSmt8GHg+i1
1Lw0hwO4lPqg8WDED9EjE6qMLYRbumbuc2ZcYAfyELzLnr4NqkKeEDoR/6M4xfCgubNH//oll5RQ
9rxWpM1VNHgrSZMLy0uAK2cuAVHEiQABiMs19Ffpa9cSBa8u9lHQJ2jCAYKO5lCp4KhV1qpqeZoC
T+MZ/aNHhMmcP0I/wZ2DbpV/MRH2Z2eM7PloX+W8PjoZApColPbcQYiCZvR/ti2F/VM7/vA7U2ue
xNGYdl5l5eIp54amIhxMc5CNpUJJoP5HHRsy7p+tQxdJkyOBPcmuhtBje5xI2QyDnHfzS0w5K8sW
EWVfKJuIMuOpjX4F5gMp4fz0dx5Ay7yCxiq9+mQ9EwRjAMmng/00ac8GhVgQMgSYK2tW+1vmq6iC
vM/lmikyIhlopngmwlIbe5mx2PN3pJDrf8N/gD/ZXHI8FAh3MBgLBAZ/zWmrT2nD2F4+RJQPCCkS
VR4BfPWr1E3WhVAv7Npl/nK8/vvYH55u+ah1RrZjcDVKLrV2zzhoFk9YC7OG4QSRYT4qjU6myrTU
93xfTO++9B7WJjLwptY9N1jYd4A68GDOAn/zjnlpzFMZTReateJWubJnjSzxHR4T3gnIkYualHpx
zr+UKIjiafmSaHDjgH5n6gwR5jpZlhdUT9M9JC2A79O4V3RnHx71vRMhylQ2KCWdC7/iCC4XQCd9
m3X+0EhktXZNz6toKnQkLYKv6uZcL7cpWPABsrcLdIR2H1Ur6mWlSzKtaqAOPpybF/QoI6RjL/gT
R+eisAObDDuwmumuZt+CMubj2A2mvfGcN2u771IkZL3YF5F76iCNh3Jd5vKxfVNkXAOqjAiakAu3
XyVej9JU156dQSLyx7UDccadVI+Z4BuwLNi2UNFMfGrLRY9oTwKVEHjgNPl+n0YrMYOcweDSA1HJ
s8nkoWOs8lTgAMdcC+Ajm7wWhn1GW1yDPjTWuKo1lllrVlgdhdWSGtmCZbVZ3jMvR/jQzqLPIRT1
zYFOPpUWQVqRmvAa6Cfp8hA2trZaxdIhfySk4wqSWy/EjATCSUXVmXqM2Tj5WsjRg8fUPxh+c02s
hSKdiNYse2Dgaz3GxYA476CH990TGpnzvsqX39fX0Tu0qSJl15JUCffC6kKE9BO0Lkretg/AMIQM
QvMYg6jxVKR9Pv9GAoCC6aHFu2Go9TQwUs2GAhgLNUnkxCFMFyC60gUHgFtgBzKrlkuQJJk7wjzp
E74IJpEKx75pbOxwVtxbhR36CkfT3d7obdvjr5eL5UmxSMpwafBYoaFJYucBLhthtIMmPlo/8Wm3
PIq15mu+T+Qanib1blmtxfpfsxHjuDncGwQLlI6m1G5hX5s3H4nDsnmGewPEfodGVRdIGpuNCE4l
9u3OtMCiV5WH7rrwMMw2Q1aJlOpU6zZQAOa0AZu+gzEigwtxuE26+sGfPdyuGfrWBVxf3a+OoZwe
tJ59iIOgULNF/F3Y4t906cfu8fCSxzMNZNCm/XUBn64Cv/uBakfSssNoRqjo4cppBSC+wLHPh1Z3
ZswD5zoWAoDacP4YXfcQkAaHICLRFUn2AuRty/x/Bgr8fZx+7xtwIAsK8OjDthUi67f/RS0KzZe5
qA1a54VzyIrMH9GJclVYVGxwfYxAutX7wYhYHYne3oqhjralPrLLrdmMf0KG/EOc4wokOwmoOmY6
RbjvPAhPCx5A3/B/dabpIOlTOHW6lF6ZEH/Qy9zRXS2/q6eFDnfR+pAu8wEnjtYtgox33E9YUa7q
ai73/x/nAEayxnizAziEZfTsyHaAePQt3hklHrU8ww//mE/odUre7o8Zet4wo1C4NuG+ORkdrlwK
ItAy+bhEbCb6BP29W1sg+EMyuH+p1ICWfxRLYt6gSNihYsTDB9G01f3TGhOrC5pMveMnF+jXS/5F
YTKUFjS/gRNTHmh6x8GDPFSfgKzMsQlmSRwfS4E3KtGtV7fi/BHSBg+1rIxomMjz5SVHhQPqywNh
vjXxmTaUYUagkt4C/bM9kjjc4CxvY/m63D+0RtblvMjsjsFEemHTGlnH8I8/9eHIVwYHYQujHYbv
WkN9O+EDlybfCfogLqUPOytrF80cb5XXq8aGdTZF3qgdkG87laASByyccTt9Dhsi9MTtmlvPN1IW
VswGqCIA5mULbGv6W3y6zFmGO5HeTj8bdNMJ4uQqGjfNwkMZvCbbaEKZCUnB0cWe7EzaR4hf097g
RPOM17tb+wyDFJeoR7/WVgjeBv5wdzcfyeLv9PV++HX5hMhudzUAz/B7kRffqY6hPdafjy47IV1f
L5njVeexp6k6pHkfHQfdIbKC2vYocVfS73z0sUevZli6Z0TAm6UTxKUDWel7pfzu3pXwry4g0tcp
EQHW7c44NIvK7XBUaeUfDbXeW0S/d/NRlfFkqgiLvHSPfHC+a/1IjNSW5qRVEhiYshh9J6H8Z0wx
AhiYaowJZOVcy2TS6ji0GuskVloqBojoKVvwNlrUJV0qhuaAFlWhvu/LzihqBvt1lp7v9J5U2jML
j+nhl9ZC5Sm/uY8qSYY3hs900RlN4Qwa4Joa4MQXGoUuj4tkdRQWoPLXOP8QtieOjxux3OF3Nel9
/H/HTDcGeBw6leA41lbdmaMW1jv7Cc9lybCO8j7E+jROrZgRSMlvLIlMLAVJiGvy8wFkrt/HSDAB
QjVPDSP07shDP18XKFSShb5ztVrYXNBnQsac4xhWXUAldSj1HPO6xIMjPR7eBtj7fI1EcvzokgIg
W6b5aqkb/HegMcVITerP5lNriES98wl2sTchsKnFiA5S3IXhkWVbaFupe/6Ygy15INe37P1yibuA
Q/sybxWJv1wUX8DhbP91JVpW9KHV9XcjcDk5EHVe95/vgBMSyaxYd5KAMUkNoxS8YjUQfPSA879T
i9WsuGbItvlPlHO+zYfqrdpnp9Tw/bHBicmaIxgcXQ+aNzvskj6eOhD/8+ZeYE9Wd5O4q1K5u9gw
YAAGljE0tlsnJcOeOOli5lCdrpyFFg58fRdECimjoK8RHStalgBgE//E4mlxKOwyiW62Hr23OO+6
vnGc6167oL+mKIlfQdYcyA2amixsJwYLuvdk4uh9yMfRiXfhug879jQj2zSivUwZU/eo8awIcIFq
3k/dzNDJD5DzQLnLIMRTl8qO61c2JgdxQWgp6/LxtPNcNt8UOtLavDEqJH7rinI/I5RUoTqLFAep
KCfAm9X5fKB3u9Vrv6VP7DZf83243jY7FyJU23VCCRL1e81nEnYRepem/3VmuMXCwRsPVxkG8G/2
+TZ1HaqzNEDL7jdmdld8etKeq7zTzLTjANPAXZ/QdwaiIZYJYsSEyEv6d+isieXIBfYTVCEiVRu1
m97eIr+7Z6qcYUZirsizYNSMzkQVr+Dfjcy/iTlcZSCkvYUxsyYcYfh31QtZ+iVEqN5i6RgJlzSo
p/EdwWYj7P3zFrNUd99cxKGqM0a+TCfWl3zDDZju60IDC4phGJEfSR54Xj2FJu/s30v55I3dy2Rw
V0H5oeCj9DokccQWoabGCLqOOteQIFSHioldHyhT3rtS1vIXw7ZIaLynizMO7ns9ctimTisKV+ua
eVzPCijpCRSq+ZcDuxUSnrnbKVC0bfCeLAipkdc//Wx75rF9ti14llZDDPpKEmW4z2hCwYca+K13
AFOItVS5IEjRFubMOHHsVLXtU3HJ4m6zZHjkFfuYy7TLm9DyAzm8VMhLmAbd/yRlIWkD9tT3cWk5
g8oGV2DKR3GAdWsuRwQFbPWktsJfZHV9A/vb5pJbHRaVneVoIvLWtEyD4LuJshMYenkYLdu2rqAI
KsGKcAVIi8oE1qQjlAJZ1Zn7Kd+avAtfdqoRvuUFVEcYy59dtCyt1in3i9r0roS+RCi8Nk8ikSp4
PCuNoM1UHTjD4gKtPpLk/LNY1eafmAxjUREa5bhVAIDJjae0cfWD9JYq1pHX/Px2KZcqZhX/4C8i
jnHxYPjI1BPmKKlN5MWuKpkoWg6SlAr1TYmB2l4ydr3m12E8TjQX0TZAQ8ZCff9C8UcylJ5qgEju
RBL5UONMhfjuE8W8MyzPiqjHX19n4SUJO8vwBkVgF3TGm1GKdaUsVUyAFUF9BJIZl0Go5WXbE+62
VnhRR4fBx3illDKorgvJdGely6rnFy9WpuMC63fCQojaal2HckW/hMNGy3AZ3mLj40fMFuOC2tKF
SWLOAKJJvNe3mUz6AwjMxjWr872SGTWv35PL8hXPC+P3KK+JSbr7b9h6u84MGya7Cwej+PZqfCMB
qyxhqexUVeLa/2hJFtyFkAuAZMQj29tyklLC8NZB8ZJtzCxBNA/8WWffKg0RGLywgS4GrMwmKtcM
bioQwz3Xbaf2sVFSHfE5pcEd6oy+WvXV35zT8wwqoib81gPEV1es2leDUVfb9RhqXz9KBo6ZRUQb
OpcsOqThV35DkpDzvajcypJWTEOrVFp/EhAceq7RakW/kNumOj+aVjDJQKxphI4/J+j0uqTux7hJ
cV3W+hzCINWZxmZcTNlV3wrKZH5ZJNBGG7ZxM0qC4qTEMkSX/xmjzLP2nsLEOWkXpZSaKCxOvLCo
G4PN5+W0BIOG37ti1aRqGyymF893vPFc8ciTdMIAYAj1xkVTU5A71F4eImLjf9MR1sb3RsMdfAVd
lXVcgmd48baBkf2jl8XC9jPaPzN1q5JxlwniMWSNbG5QqCkyzmQJX0CX+zljMEYnJvgcIcPkoJUY
m4dKQgpXHE0VhAUWE2kAZcFSYu0C121m43+RiJq9VhC9SVF33qbcc26LI04KKJ3oHa6FrGcOjir6
FSlVDg8b9dmsnmZ76wfaiojrOq/NsEhcVKF5cFrMIeXSTHOhgvnPKVP/0DxZCqvV7NyLzb3cEdMR
HK+KgqaaUgMCqqMASRIbJD9kmudprnKChQ723vCJQkoqo8QL/tcU0TxJrqxmsT1iQe8LZ1aQjoOa
nVuynA9XrGtUzIF8b1s1nuHbetTbz3GvjmspLoS9yfxRKo4aGNHAN4m/7xKG7inMu34BH6/V8GhV
qK24kmlUKs9gmpHhjJJE4aqLkbj4ufggCIx+kmlsCZeLV9LhKcUoqvYJE3qdtgx8UJDfWxIfBQHm
R2nOr3jDpMFXZdJsHqxsbbwl8svcXe36TGGyh0aT0sv/2Z+BaeWWPuXx1baTd7at3UkaAo6au5kF
KXt/3Zx6xPgxW+bRm8v0REuro8wjAVL5DSlNC3MGJlwFP+2OCxZ+DRANHwrNjeXyGkI59UF5qCt6
zFWIDbU/U9Id5uMbXrNEPmJOmO/l8HNTIjFLR/a+bDXaup9CmiuKH8CW+lVCsvq8ZUqJOIQLDs2y
qiuWChtiRBzu6Y4NArlWTDBdh9QvRQ9zG3w/3y5IhfdpFzds/AZDJ7pfOBP1ii6Pv/aqp7JhRraC
LRoYnF2Q+ZSd0MLyv3jO3PnvnBURHLoVqBSmPhmh7xgSXnnMugh0b0Gs7kW4nR5i1CH0JDaLJz+K
YtogNWUYAEqLObvi0SnDAtsGxtBQCZcarAENOLWhOuBLwEEE0MbmqDkZr3Ol4Ew/0T+Wdq4z8dLN
G+vLqRv2uXK9mD2T0bbCyFlKDlrPfCmqi9EDQszjhUsjjeQ6SL9AcNfg2/oxP98TJx16XJ7Cq39j
fk8cjyJ/UgQx7e0c4PSqbogaCuwK9uhaRVKxTa+Yi5pJL4RP8/C59iA/5ANa6AATrVZpOyHG8V0a
FaYhBU41kpDF00ulOXlhhpKF5+RR69mi3Dmdytv0K3DLj4jLCinlM4dYspSXwIqF4rIVbbRE+imF
FwaFpPAqifinCgzkTpF/FEGLwJr6ob26gJuo6TOGRlz//wS410h86TRmT6EFhLPD4bgkziR5XHa4
bHm1bStFFuF9jmYHNXwHZqjKvSLFG5+l6F4HBOdhhksyPgMDneGtgVB4sxodNef6sx+WffojpnwN
/Oz+UkDCnWHinzcCoiZ2BADYsGywy5rfuw6Hui6gZIqV3IhSFQw5mH12PlgNsVX28q+acdlgkM3o
FNprhaD30rD4CYNuHzd1i2cyJqMlsxG2FmNOohrzttDUqvGxUIig7/zUqaUklfm3+ch+zOjqRcfn
R9/ByFmuaiMsM4iduzJOTJg8U/mx7SsWsKUiI0+Z4mp/O6I8+V9wCDw0cb24biYVIuRYJNld4jrE
okBppjL3tPDv+trDrn8svu/1vSDFXjW41EUm/aKr8A/TxiSV6DLjqBQ4zWYhk+cZQDV+mOH7WrYg
GgYFpt7mqY/VGLJehO7IWdMQhQj/AEqs8rBJ2Gy/FsKsK+2w7nt8xzzX/WfNSxxXpwgs3fqAWXpr
+N/f/tpzvIO7pMDOK6nUI952HnebeZ8CE7y6yaGH4eFJsLpHIjBzYq8Gi2n3Ozc0Btd2ZXnCBI52
gQ3GRRo7yuISqzORredGByJQkiWmjRq/WN7xkk6U2yPdZP2nJrLzicyk115id4uhZfoDuBO3EbtD
5FGLQfvoBgvi/5BGkjbwo/jAbezYHYaN7rnxImVh2IRObUr4ADtkgSWnItSVXjhEeVuFRUSqMp+H
zN3RL/8rhQJXPOcmB0pj/p6NHVNQKnROotKLtxp2bXJWmpKKlNzXgD4J0Mw3TuUwFJG+Xc7FYHtX
Kvq3b9MT0AclzYH3IDJTzRQJw7DB7JYEaie+57ylT9bm0X4KkG10iIr/46LhWWY4DetkY5lqLC7U
XYznhqLZrvFWl7tsXvuKCmFb0P9nZgNzisRSHqwqvO6ywMgrpbkGdXtkFQD+Zz26jMzLARuqAQDT
CtNuRFyxC188Gpo6/McsHFcepGI3PoGKtvnWqJ4NEcKgIZoza2pm/hOwPaYQpvU4NTEB87MZDfX3
LY+F4YOjsJiv8sUwz1mkKtoLq8K3u4PSTYm3U8XvFlbH7kwMvm2LjnMJcISKu5Kzl02KxiZ3yzRt
WQwdnVVaUHiLGZjnP/vofpJ4MELdi9R1GFFGPcM87noiPD5cPuHpo9nrFBS52RA3sYK7lM/a1rUF
+EbacYZSWZhGSqYdtsVt8NiltL2yeZHbf76wAXxUYf7/7ZwRraGvCTE22CsXSAlWGH3VSnxznsbH
/iOCZo7RN2swhgnDUdmVSmVwdqTXTTFU8hrsgRW6PzA8zHNb3r+62tV8YndXKWwHL84vHx5bhLEl
0pAEVU+nABeFG8g27dWGfnJCiCHB/i+GuPzvKnhheDbvrie2G7dZJx+f4uhDkwHZas/Xr2wDHrbf
o9AOw1M5QzXoALz18en98F0CHzAQ8dblUdm16SAhcv6eNLZ4Uqzq8dccRlXB7U4tIs22FihGhwMU
nBT1yPeYk+u6geC7YJFsdPfM21Seg+abc/i/B7lCWI43W11lylhXJWZY2ksxWgqcgFvZfFDd1N+r
mk1b+5rB0aSgtt8jRgN8ZQlXVHu4DlY4Apwa35uqKudIETW6tM4dU8UM8Y81S0uEEzX4EdJYK+JW
3E6MEV3C2hHfCsX95HsTobhp2SPvbxPtFCaXcuhi5bYf3z61nAbblqn98Knx4ysFivUQpWFW1ASS
rrmQsRocz5m9BMk74m9lrKUW2T5nyiWDco96teu4HS2sQuWkLBYz3+XlqWEejfXZOJGNW3iybjaL
geMpwjuHHenAaEbODVgDRKCV047rvWcNjToij9lLFweTNxBKeEPh8E9SnWiR23yDDRrHNtQ0gRda
T3oFDGpsgrQI87Ynw5b4kFdTCVPWe5ZaYEY53IeF2DtBdNOL3VgciNx0C3x0tTMFhrxuCU3Mn+MD
fxhAv0qGvV6U9ORwJKHK9NFLae+lP309xZL73F92Gf+FajAI878ZPmJ+4NHtONmsklsVU+afbLnC
v67//Cxs79tj4m7n536Kmb3PYBjmdUGxxM31/uhRwAXMVbQJpt1Vi1YRlE47q+YiluMHdfgwdtne
ZZYnfnB7Onc3zvvqVeioRGyF+LyFFsiBMHYrKvaL3NjpeiuuwT6LGgCl/4GpCOfgnN2S6tygKkFx
2P7BADZ6mUzDi/G4txZBiLfo9AqfXTiSdFbMGqKD7q3LsRAY0Hzdp6qunB1V9YzL9JoerwXTl5xx
R5R11OjhF/TvEmLrOF3VpCZNDKHrS3vwXHm/iuAxWMaIFIZkXWwAf239eNWH9SBOiSNVfUCPgVPf
jQyYVwsrtPD4YdOOkWYeBC7A1JC0Cc6tm9eBDNBD3lIcOYVDABj1YRXwP/uPWtpOLpyHYfYVXGlc
utumruTM7vIvKz3MNFs/VtAtmDOEhL5RLBdbBepvX7OmhvhonC4oQ23TJqqokTaFfMHjxj+1G1M5
6qIXAwHRtpaP9Zm0j5FXb1qYqigu7+xuZH1loou9vsv17Z0yB4nTOcEtb/DzaROwLD3VDhItFdK7
KaBV3APSfQq1h7DpowE9ouwBoGIEm0T68QQtme2pC8aKUyzk0dXOfoJGk9Zo7B5WXjgE3YFbyfxP
KzBxzug9n36OzyQ4SCEg2GCYEoY8OsgNEYucyBn8/2rGvxc5Lgg3gNiW5qH0vDwysdKgVixsCUNz
i1Ih0S4Th1IewgXhXJz7vQAAZ1LaZWwscvbqxUHpq9WDEz9oCz6qOpRG735ZxaplDanXGe52KwsH
LttWSb7SBK1pr4+bsxbKaKp7eud9s4zyqXUdmhRPw+GMrFXNQDLFGVO4M0L8gUo6q4CPv+cuYTog
7qt82/PVEnLFh/3Ir4KTJkTChC2CgBLKC3IqgA+IO4X8UAfS2f316jBn4ixpJwm3WgmYh1Op8+43
qRr81h78dFb3z/9zercEh/Omi5Ykesi0UcV0A1MvkvVosfU4LEv0CfjIz29pKSIuvHWAs49qSeP2
uV7/hA2GUREKRqz7giN/5JDRXj728ZypQ7eTlmbosLaLz/Bh2qf6dlSxvdIiD3I9Ev5IEFn1f1Rb
7xOWaQg1Z6W4SRZVA2jKZ8422gHYRR7rPDIHZVDCKERDu9XmaV+h/nLQwo54Vb1f/tWgtAccYvHl
jmzwEFtemBWPlzHrWBRYl+1RxmKFapTR9pb7O8TQWbUNysp7kyTnNG5+ZsHgVXCDHsi0seam77cc
tPBW4c0XcD0Iaoc8aukW4yBmS23E1H8anGMfhMWjSH2/l71K5Fj+mDLyqeeyY0g6srANjUgFVq7d
Rp6G8IGan0s3eRyekqNAwfQ2wPR5xIX6CDUihtVvjcx1DKjPjhRyGMZDufFOj5jp4uFNKntg3YsQ
zpDQe0gXxZ7sbnmd1njI1pGYEcBMqUej24r8thkn2u1PJL1WguUHVD7k0cUtbiLyelSnHBsKFkCI
Dnr2gpX1JffdwbgP+bqvrvc/RKzR2D5aLlMKh9GWyCT4G+hWOLKbRJVNyOffa5aJ8503pcsULTau
G2+5IySC16gtlq+YT4LSedt+ts3FJmBs3cagW74Atc+bCt3MVTA8SloBwm7P5dc0JfmZOr8vZmKZ
s4GWSAtJQfS7IYo0mBNKzf/UBfZbhRvBcs3WA4uBmLhHyC2M/zqL3rq57mGDuRMLeIhghLeqoqhD
cYKVh2x9bzSQDeui4xzJaITt3HpmrzlynKdzrEAHbV5SO8i5N2XLFvYTk9qu07SsDfCuMkcClm2q
b1MFaDxpfP8afCaeAbOCE/MDSXuWy9y+/oui4t9Z0A6wzC0zP54IDzsCbdLhl8/w6xkDBvwUXwIn
ldO3hS9AZRofkilZEJvWQZNBmYCwdP2Jrl5S37FU/bXg0kut7JF65sm2fDFscMBxfzruFbsotO4C
wfpcJgOgr749nCwFLXXKlsNeLZkwLQ8R2Jy0lhgvikLqDLSP1v6zELl6JVJSNa3V1P+zuELXSHuo
3pvsynHqJDiWpRMCgd7zzfXaq0cCq55/A1udPi4wLpaeUNfGuc3ZTdCFxKrFTK4/jkYepSHAVicH
4uGuPydvcV44PYHxJbHAK2ASt7WtHrK8iIXvxWIagj9gXQdqe5shuRYzWdtC5hLiF1zwZ+4X7kDj
Z37gZ2S776h1UMx/PrOa5kZ3EXD0LFMXnApp1GxfBDSGAFIyvPy4Y+JEfRLobMoXFhXEoZFBvHTR
6tv5WnpNYcvVhfGra8M7WsaTmIyGDCwnP4J7acSGlj09MX4jZBJBXsoNVrpucfxq5p/xXAwBYLW4
E/hPXaZL72ALadKDpPMibkcJDtpvNPIHsOkH2Y7fs5dlD3lamW+YeKVCJMcUSew2LYuizuOla6pe
G1+3ftzITjFIG8DJIPL3mow1itjBKlwQFxJoRdDE2e3IXWcyNFNkuLsX5eNeCBQHHReBZLVIwH1U
tIrwqNrhe8AqCOiP6XOmNoMcVFyfxfDeK4mgGS7oNjdeaf82TV1DN30opMJS7eKaR7vyLS6EGSS8
gs2HdqbS0sa+abYX5b5OSrebEUg3aZoAXuQeVTTTuGU40eYPpuddGfkqw7Idjev/7+J1Uxlu+jQ8
5EWiQ5mBU2nhJ7jiW2muU/eSjaZK/2WAqr7BZKD6yd2aYNhAppyKWsiT+G+l1R+5sgMXoDyFBrCf
Kj2z4U4t6Xn6Of3vj/51eiYuuTYyzvQD7oH5Nc2liBvE6zz8RH1ewobxfZ+oMqrOTHZukmoKzzfe
YWDLBk+a1NhKJuEVDKVmKJE2O2KA2XptA/KcrZSBN16vju7oH9VPKVvsDm9tU3rx0WWwdKr/5Uxd
m2tH7Tse9X9Gd3oY7rp8zeXA31Ufc/QHWZwVUQ/JG/pdmowpPk9XiZTlRQxEdY0DK/ttSyeuA0BL
7KwrQoi8vJyUHKpeNH9SNaAvpmxUzKtLUoJlObfcbRmF2tlyjyaSy8ikPJwqxL2biBAMFBUl9YPW
bGPf7C8SgShkbrjRmLSgzU8BRDkAoP3L7GnrSybE1RmLt7o56YX/d6Spf81b+/c2GhPs4mI/j2/2
O4e5O0AWUxZrCvyuTAz+LoKZgEr0LSK2psbvcfAqtYWuEy6D5lEwevP4xUDxOxpCo2cvwMWSWgAd
Ce1V/99TFYCNE5o8zyYSlDoOvwv399sOG6z/BDk0EMAsQbRUAo5+8tgioH2cFF8xfrAhbuCQxkAw
EknDmpbLv6gbuoHirD7t/rMIBuvNjpCze1ZQQfRGhang0xOgsyb4zJ6M91ESg9E3kBDBPmVPiT6U
d7XZ/MO2WlspxlNLSglqeR5xujviACpoAQf1EijmVKp6D0F8T64YbOq2MXejyJtnSL0trQDTdrdh
6MjqvE2Zlj8G0cGpxVcdwfBgoPyhsz6vDK/virYuaHMO2l/sXf527ssmek/d8bDmNlyDrbGBY2zS
qZuqZYsx+BhTPG3hmJpqn2Ni+Iu+MlAg1nAUupvX5qQFqo6qtKL8CuOyNFjSUEBx9ympP8ozwrff
9pfxPNfFJPlOqlfK3bJpHPDm7zoR4bn/ikd4u+3bGZ/NqFcJpNUHHMBI1tpHmbV35XqnUjVR0fJj
R8etetotDplVOY1ff/BjnikRh6Stqjiru1O5ouHTc4UAQ3KLWZYun96IK8+tMKQ2B0mNK1KOct7/
fUjibuqHOu0Lu05ygACNHj77ksauz3I0P1KDpTRF2dKAJxXaPYqGqNauIYe9xuOg1Si5BIiCKVw+
Z9oyh5nqgPrB6CmQPsZttNS6GmypoMWIZJ5g8Q600lb1uRng2VTic6+k8ArF9QSUhHdWPurJU6yD
FtZdCnImOKYM4PmPDrTuE91ejPuGxghjUiOU73ylymyLyxSiBHVzaEK/zueqfb6B4JlXQTv7i1tp
3yVeMtjESAvP74WskiUDA8VtqQw0RfKs9RcqZa4A8ldSZl0WQW0+QSHPSi6UGqy9Ad9Bd/yBpXGY
qIxtdLkDf4/iPhrvwbRySWf/DGap0n5/GR4qNnf04ZATlmxcSYeRboNeC91Dy4nr7ge6+YgghlBZ
E5tU7CFSNYnxaVNycA+muBi9b0nzIpqZacQn/LCEGHkH2+1N1oJGDLaPrdLZf+tgfaU8WdfpKNMd
jMGarGGUjz4vpBaiEy9H55i5LYLuMM4Iryxxdxy84op+mtHoj/bSfO+y1fDIGtFNLy/LFlHj9h/C
uHBpMqyLv6nE995PSTdPO3n1UbI7f/EpHLrJoXnuUtrtfkP/Rt3uRVtj/UP+JceIaE9BD7XY7oaY
snFwf55Qddtb76bOCFzMaFF6Z6S9q1u8Pq+ZLzxhEolvubGPt5q2J3tyXewfaC3Vx04M28OWH9Wi
eGukQ42Vh8LysmDw2oTmPh0LSwd6j4Y0g63PeGB/t0K4oiHCxnzzwoI9aoJjXBE6cvrw3lmmpbRe
wIAuh8OFQCfhdAaC/qEXyTPr89NAXNxuUik6LtyYmUfTZOIh4CG+m2UQKvaSLeM3N5U0i5FI++BK
5xR23l0irf0UgzDPLfYSO4MgVZosMJljMOipi/NDIN1PlhPTINqHS39QWanpLPcSgl2uEwasXkX6
yKHenNJdkmZ3XD9k3bCjWZFCavAH2JpcuhXfAfcVOrhOQs2Y0Hf9MkZhYbXjkOXxYO9RjIDuFoMH
UuJkRpaLWiN6nN3CeBEuqK3qns3LZDNKRYESJiOHwTI5ANHMtQc866Ydd5R0NpryzYVAp/nmcYXs
Q67cXyusHawlZ8tgrVkr8OIVdNamwAvG8D/qnRbgk6At8C+RGQCCNF59bH+J3rVLD5BmVMWIJhzW
S9+ANjasgitkxpclpeA5vI5hzh1BhipVcXPxWhuzVCiytuys09FgB25AHfviKheVtVohXRa6cvCK
0GXKOMzU2jQkw4GZtU3gnMPi795Uhk0XYNJGzfoQHq8ERqTIhJUIeNThKLD/Ca1pCBclAg5DbLir
qZW01fb0m9I7hdtVi5zpZ5ztM2Sj4HkLmo8UyrF/K41eeJJMAP9bYNEwtwZQoxkKpPXSf0o+Wnvy
d86o0/rPVJI4L7D8G2EUlUWu0G0A2GbvBxn2yRDQgH+OMNLyNF0iSpgh9GKMQy5ouxGzH1YWT1xx
ui6U6ooD/X3UK/qxMSs1NqKM8U67vTDGAmw3ynjK7IFUYfcxNFGK2mQmMcqqkulGq8/c9FzC6+wj
P1l/LBK7MK3g+mGcs58WAftHGuyR0kf29toFycg8bT7BCgeop5OTQjEcIIFOpAnhocv5oulxfik0
P0gwaNoBDjZtthyc6a2kufvcvHmpVGbwVr6MLBTXsLhdqq6aIJTZNJps0HqUbqIhZ1TJ+tIGpPid
CkaiRlek/uLup2Mn5S1ETXd42mq+KbZBiA9Pe0+N1YCkBDSX6buBD/VExiLjS1WYt4vfLxlWMGkG
OOeFLe28OF2e81X5psT/mbfXbYf1FQboJOP8GFx3/ytZfl94yLFttta4DfYpo38W45zqN5aUVkG6
C8ViU4VQUGTgcn0w8BnduKSlS2eLVtXeVfv8Jl4upjMr44yubESiaqeSXy4yOMB+v2f0hbvClp5u
DEscFCoVszcWeqlFwGs/+plsmbXOtwm1gKVAeY4kQfntE32g8fnzjvWWWPLD6n9JrKH2/Rze6gI1
Od3jlaEZcYGvsYN+AVjb/h2kDAsJ43HtS6/c2Wccz5//dFTObVEvNf/gx6rOtnWQY2ofEh+NUEMi
qLC6XQssr0OFo/HWL2X7WfMnNcLh2C0jWBs5eAcSVrq2cs1G3v1C/E95gOnf3C9xx4sU9fyLmMyM
0wsSUlQ/3DU5fMkefYokKL+DQTmUxKqDQIya2h4lJasytilIVMMhD+LPMfzaqoD/EzN5jLhe0Ysv
xMNWMFOxbtP/fRawFeQ0uHO0ATOQ1SZvSgwOJjbJDNCrVb6XUdBCZFQpGbuf/OBsWPl2HRC3aVNM
uT6DqLWVT+cIOMQX1el+iIA3XZ2qMydWIEh7aRzEjD/Fr8kexzgCzZLKaJrWsbZi+EZDTiBcKB5P
TyoGRtXFTlUpmw7Y4CuajqaPdMigG+C198Xd/ns4EERurL+TTm52EwIjvHM+KPzyxqmgopk5hQu6
NdKu1iu6fubJitGGIL4eANIe/b6CWW+NUYa/sPcThf7Fw2v0V0vm7OmBWScxyNjXI9FUHCdI2Cf4
xJa28lZFb1PazoTU9V3EmgZcxMty6weduF1aFiaVYm/cCrcsdK0ZrWgj/jP2R9SpSV2co0mGz3Un
VewGccxlm7JDNYObOukn9rLhNNW93jodAtoO1K9iRtHLcmH80nnlFWNhaAya0gJp6tE/baBiR77a
85EBm6eS+FYLzjUplDUWvThUYqCUdwt9zDQ3+9O7fD4IijGe0QlRUUUynxY1zDywvnZMyzlpFWc2
f0gr9noo3PUv7UtCXHipjbdqAN4JSSoSijfGt3HkVi6ZVAvVTac3pKWBbwzUBA0MwciEkDO8UK+9
pKFw6jl6j+gIH7VCT/ufwXkzuwbfKNCg7EMP0eDYXfjypJeZ7zYZu6UBS8dnMIZE64eyx4tX/9KC
VNjZB/bKdFbVHwaeFpbvw3scZ4WMuUl3r6/jAOBv9RznmwR662xJ4rMARvLlhyb27OeZPY7fUe0z
a3M/MCXa34VZQZeK9U97G3QTzpF0jM6neeY7NiACapkjtFN5UN+vb5l+sckF3kpw903lhYS29ot+
KtineU9/IcDeI4emgEORBYUBw4Lw1EVecV3C3X1J5zhh6vXazTWdUgamBNnenemNkm4a4vQAi2YE
AqN+LvtJHGEmwMp+qu6bFScbTDgKs6WhyMNmaBctfCtNSCLbAZKraP3v6Gzi6hY5PBlMFl2AAhAm
JT2bKFCJubmEr3LgjbP+0g1qgwNpX1l7dPIiZx3SIgMXny6N4ZeNwM/syn0MzIdLSXgWbAtoLzJP
2BEb9U+SJsHugiQJL3c6PcXlIwtmXJ69dRsv9jfbdEDqUD5l06q3jX5hHLfSTXa4IC6pHl6YhDWr
vI/q8ksFA/KXSwd4qsX5bCBvl1++KyFxc5jtP0DadXJHR+wCKrXZlO34UvSSZLThvoxQPhPss+SE
dCxM/9JwUdiMWVGuVml5+WkE8ham96wWgrspzwplYY7w7uW4hbV5x9HwPRbnLornrFIvRCbajbYl
p7wQVNVgMIwY0oLVWDGYmEq4w9JnjHYV+esli7MqFMEmWNvnRe1Se5r/IvEkIaBHvuPbzSIwQuEh
B3/c34dbIvyJkNLjvZoba67Bt4r+g+QBl/cefsNi+2MZ5WF66O9yQNOeYnBgRl91exmoXR20wlWt
fl46Oz3egqXcUWZZtd/sLyseGEbBBtJeHdXtppjC8+MNSiTNtqoIBzafGQyPNsi5Qk5bhBocfXl1
UFw+LdYwIuIooT7SyROCSa0lH6d+O97Vt7IoPhDPbp7p7VwoAnqGQVAbAWIpK1NVYrSXVX8xWqCu
aO9lv1ZZen0AN8BDfbzQNKz3namFmsOo1ckM6rVCoX6N/1aXPuQb6H/UG7nPlBImS/KbSdxdu9Gj
7UfbikSlhBWoJeQDmXFstFjD2A1NtoS3g9fcqqbCfyE2+a03D6Wtg5wEIPuVMWauhrt41i4FRVke
2n6nkH/zYQcVdL56fINo01P6S4YePNEXIL0iXfyagwogeeKs9y1VHBowaOHnrOdv+TfoQ/guCUJn
SbnlfzMzSnW/OvQangV+Mi6W0QuSx1+2DM4Z9E/s08T0i+Ce8D1j1+4dy5ffexTwEXpNppYqK23H
3EfGukBLSC0H5ctlWve6AW4p681r50uKwUtZRg+womnrbi0V3qrlJTtvybpiawf5Lcf6mt9jxKcG
/v5fyCjdvWkhL8UEi1o+rbKBEgd0rDYNWSfKxz6uDVzxQIXasgXZBU8UDvhoiz3R0ePrCHGSWpGW
P+ihgCcgekew6+qNLmN1zyk10hXpGVt2Ck/gcVRXI1smllbQbWB1I6xsEGPI5RjHuXmMluCHCrJI
nX83vB8FoYEwrE8EKodUOiQPTqRo8wcQBF8cmNn+SHMFKKBrbLJYcthemdId2s4aZQ0SDemtysI8
qlca2eCW1LuWf4txrWIMZhio5iO8QlVKANMMMPrjkwUjMAUy4Sv7ScgNmZAnwsdspbp0mHkml8nK
G7tgNNfa+HdNRh7Z4oSwLNctqW4PJxNcNErnlCpO9pV1iAjwYO1KwF3DOekaw95tOTaPlj+0r7ah
C2AdKhpaXL4FpaB5sVlJ74jDVOH2Pgfl2yUHAsWyvbHcgnX95iM7Q4qtNsrjVnbgYjVGZCUN6Lq/
lYof+w7mGl4TUFK6WLvBfTcciSim5oWX79pZfyFNxhYXLlLCCZUTb2b2c4oMSiyLdfxF1seMCaKt
KtSfBAlW2zoutf4gZ/0KIT/okuu4C7bEVn+CxmP87C3a7CU17QfO2D6jcBJOpHGoBogtAsbVmvlR
9YKFm52Y8120RbbPZZWk/qO1JP8LJ+CNt+E/6IEPNKUohqUPr43OskuwPNDmEBC2oP0Cu7tRWqCx
yAHX7p+YXMyUH0HaSNSY1tttVX53f60ajKobjSegTmGzhwBJa8/FQhMZ2Pm8DuCkNxeBWi2N190p
eipT+dQlgyALwaQ3JudqR2kolN6eL+snn3ND3UZBSb4TEVrdr6S57n9yXoa9LzchsCgz+E7Ipxfc
rQg7+KCcs5A13TOM60zh+8ANMPfbBO9PyQQF74cQ39Mhg/q4oIrqh1p2ULwRhqjsPJbdWmmsKUSp
S78DCUIF+OmRqsCiilD0xVNrR9IYUwUNH3WKM+RHXh09h//+qb45VXoTz0NPnWEP+1LHivBRL+FC
O4kaALSswdL+XnbAnhH73GDv152hbJZQSCXPLslv4wF7HjYudJppZzsJva62E1RccZuklAf/HYN9
+fQCLvD2zQZNK2MB5KVXZwgoGlEfbQLVAr3FJH/8sBpy63Jr6FaFh2L043mBRdh7mQxhe8ASJ/6p
UmUeKqI87HWKDvJHHPgdzTM+2m42bW62XLTHINLxafG6CTCXkXRs+ZIKa7Yo9FFpEhSy0y2C/ica
QA5ICg3vV2KeRc43D4bLIXNERw2OVxx2mwKinSIzwIdlCYchbvkTNaxEFxZdkGaN8kpjGx6GmGyc
S6gGz6dVTll1mz6ME0MCwUvIsObfHA7jR7L2ORLL3gOJooF/G1IX49Vd4OoIATm0Xd72fmpmXx2S
ls0cEKyJ7TJjE+DD1ZL2cZgGft4rm9Kz+SYKFtYwFxAxZaRvZfEKAKfxQDcCEo6+SFKkh/PomlxA
x1uufknpDYuF1qtx+jy1VOuyR+9w4H9n4bE4tTjrMKVp0IuGJXJ4yzLiSRZJrTd3UGoSQerkoQ6O
9ITQu2zXmCFdTv5adbw632hvtjYgb8r+FGKwV+S+JoBykymeAL7QLal/Xr0akVeJe3IJC7nBE/db
Z1TvcgToM66lMHpGq88rz/ujPueCedDo/hCD7C5kZXzVVY0ZZQqMVymexUpbRgMz7ZPyHtwurvx0
9FKHeJeji5nXdHlLKC2aGAx1fd4duCiBbKOpfQcM5S9REk7AkuBN/xjddJUOd6MwK0UQTR4nzkuL
k/qKBCjC55mzSYoKmnQw1M0VV9lofpOOip+xkikCJtffW4IeRszpqOIeevbglKt3OU8Qy/g0xuu1
mfWKKZGao5apJu48CRMcsW0zvjTa5kH3Zd0Tx6TpnpxmMzD1D8rF3Tq7+JO1sok8Yk2hE/hEd9MP
mcHcbi9U3oFk/VNkY7BQdYwKvUfM4zHgBG81LinF7H6zsQp7amnR23+bv+z3XkpcB9KmEoxkgd0E
pLl/qoQceMdKtBIaFEm9TcLnMIUNjGpzzXF1cIsDa+FdQsfRbqWgMStCxVVhiY4oVd6kbuIM1OLr
fbfgq4jjC1Ws5ZqGPxvpj4qWuQQKD+zYOJHq0UWkq/AHTUroWbdyy94ZDDuuoSv2L6+arnD5yqYu
6VmOsVSdwBSW+f6VpmTG9EjACGqAcjoE3FMW/ZnjgL81GIHtpxvpVlrVIeggVwwWJD0GGd0c7KKL
1si17r9fbgMme1MvSpr7+RFi6DlobQeFtc/8lmyqC7PWf8sw/UzXawQvzrDszJm+JHaq58Pbct6u
ETUzkmq9aRaFaUoWe3/jDGdZriKRUCWyZ+TJgxUb7yk0sN5HoORTNNfvlMjVLaFQ2LYjDOzPOEFN
Jkvt4+1XP2Jfsiqmf7VtddNw/4gADyQ4c6u4yUg6DmnLFR9yeThtSTKBrLV4lgyYF2PVFY52/J7J
LEm1EL25/rf+b7EPkkgOMSk80bnhDxSuBJCDcY53br7orDsiwqxOkYY5NJrHqHvSC6tVOO8YntMH
P0FNI3QZRQLuWqu8sNqs3C9f7fPtqfhcAD1cY05SIYpGqd9z3DrtjX+GMQjiz2INjuclyYJm/oGC
JS2rs0xlJAV0NINZMhRkf76hHdPeRSbinXgQAGl0IEzqEs78TfQcYKjly0X5eCoY+QgnYQCQUqtt
CGYRekZcumlnU1uP4S+FTMgPJqFPJobYvKKJSznZpyqj60w9jMW0giclxdsZQk402PZeaXHXFq+U
ZUoRgUXbKmmmZpix/zLbt1x58gS0n0lfFLOUl2tjelox0aMGUQ4NqaFOF9SXqmGdZ/E6R4XD6iWs
KUQ6BLJXtrzAlSiS/LNCV78AHcMJ8xzQyIm7xNm0+aEzAtLWkZjh2cAhiVUmTXdvuOjHgqZuZOSc
aepgcGCXy3gF84pvMg0E1RAHRT4MPMrFGXDHqM/r6wh6Ki7OTcmr6jhc3OTK3AhSSxfFgEFnb+yk
zdQ2eSVT7GDCXCE5OpR2aYV2TlhLKAIC1gCxqolTxCMkB6idyKnrmbc7ar7uz2c8Q5At0LOaEpXi
MqyBPQN9lehirRhYWAjLc5EimrDnm2JGdZI6Drdeqo01FXUjmDiPWZxhl6atHJ+KcuWBBOB3EmEr
3CPHroCvvB355PBm90PDPwOBGotwDACETnxJLzg+Meqoaz41ogQZfMiuv3TTc5nHSTicSjofKBBS
qbcnv46CMbBv21LSI3GWHY8VC1COr+Ym7bzogW/IrDIKM+v538brDwSVJSZISNkqIVwWtNM2qoSg
zv64f2M2i1iEnL5E+AZ7E8BkHA6FPHPIf4TRmjJfEPBmMmzn0FUkyNxc+P4SX9RCpq8DIiQXm4Rc
kFueFoxJlJDgSbPS2VeB/7Z1n56pPj/vP0KNIeuEQjPzHVo+K1OWPjRuXiAjz/4h3sA7X6tKTlY3
oyy9SKMjx40CA+c91egB37K1ll9cAf9GQlKZ7DNthzHh1J7Ad9HZi5tj0y7x0YR2yz40L3ue1d5V
Tn9K9KMzpEf1EK6wrPOAOmw9cydnFmswS98Xl15vzBOVJIuQvRZopFxn12unbBhUSZa9YLHjYHD2
b7YL7Bom3+8dqIEYylIVwG7w6g62CrbEkNKilG4fn/KVV0JMCzdSzlhFyn2IBU2goeGXLUWUC6I8
4O2/u5Oovmi3TiOwL3+2jOfwVoNxmSQSF9N2gVShGEAEMKCxhrXOpfexdHO4FwINvbDKXfQM4pAN
AGV9xJJfqklgiahW87oT7rzV9af+cWOLlRpHvoRAsUaOci1nO2QXZbarLI0DmzS0486vd+3mtcbE
/PMiGqjr4qVxG3Xm/rEHHC1fbt/rDUYUMHjB2AY83Eso6yWTpuO4ZlEbQW4rvc+y3H2/Y5dIEa0Q
1Q8l79KtUe2bb2F4Ybf41+d1kuFh5W3aEyqXyGbmKbM4IcRPMojFXRTEzbNGms3XtX0AN/wVKMWD
1NkjmF0SbSS2etgpXRGRVXOxfUCF+pKFCRE8FHWDC4t0ge75zN67ynNJvpKSPr+AVIiXm0gnh00r
pX55H7xIWzJhVMK8t98lzJLY4ottHUt1fcn5CdD9AAplPUXhzwMXQTKnZxgTEPdHrzLEfIQl1g3I
iTkjr7KM3K8CeTnhojQzRrqqOBP/oUgs+4mzR9EHx8EtO8g6BSIvxGGnItkLldd8wMZWVlmOveka
QG7VKd6LrvhUcEubLUSJEwTfzgvHmQSTT7Vm+MM8cpvEqXQTRnQDWiix+dsaInr2A1LP8n8KcrNu
LdJKFtR88oNKHXF3v1VcRzMi57IG+TAR5dtxGmZ72lx/OyLpifr87ZvdX9cvABEBtSIQc1sMi+zk
Utxr2JhHjXEYQ3fFJVMoRq99tAEcNOlaLAJgO+FFfnP39dccQJ9lf9b6Zq8DCJT1iIh3XJTrfd82
LyIu/XaFCTZz8mXARMlzbRQJLU397UE8UztjXQVBYYL6KI23C6ZZH9e4jVid+feKQgcqPNrjeMsr
C94R9O5vYhPeLRcT/w1ZExiXn4hIHWrp4+8knX3LJZ228C+zOM9w2lSs2jwrqgoe44qzcPsEUH/q
t3Ix7rLnIC3WfKOPe2REw+o/wWk1lZ4oHjRkAg4oZDN3PqhQjyi5mwv4s9bHVXS492z7KxMhLBeA
En5rzcXoUYf0FI2IgEZuJT7v7WhcFGWpdO960KzgnHnm2BS5LYOTCx3R27zZLhMlgNKf90pQK9LR
bxjtd90Zy0OWL4BQN3spHMVxE/KvsKNBqAL10aAxP69QMyprdyUWVIhU5B0W9SxanhuEsgMr02sP
sw2xJKUqJIA9uhfDA62Tjr4Iv5F0tS02azIc8vhIVQESNmZXnh8E+pNiIZlrpkM8UiSJyZ2x8M+o
rrlHGrgdiT4OFkdaZjRB7BLFQrD3nb+wBityWUZiifLLFnjtL1rzvt3u5CXtmQivlBbdIyBLM4K2
1jUgsV3NJMoj2I6uFo4FOQjAbtcPrN1+0ErkOl/HW8JkiCKUBSzAe0HvuJpLTJrj2SP0BCONgIwD
F9I+9qsYi/VXxjBCkPY6I7dAQisJ+pingnyq1C9yQKRAFjkDwGM7xk3naSsgj2/fTjz+7bFWxAcy
kB9D01pY4lSGNuylbGi627Afp/fMeqaiFWihePTdCNbbvpKrE4pbOOjrg8j0zE/MVBzAKIfcDSoA
SLB6oFrRhdY2HfsIxmu8gSYV1HzfPCg2WkkYJKDsabndwhFiAna6pNSzI7JE/1USYqBBexA51/IQ
u5T+vspauRWeaiO+MnCg7RLuL30b9y7Vtkp3snn6DS6ILmd0NHBWnT2AUmx9LFRUZFcLeDl4dRjJ
JUtrv6qxmYWqKrI1y914h1dzvL8fkkBv1cfln1xuCiIIea8f/3udlWxz46bhxQlYrePDWDNmFSrF
TfADixkHRYMer8XmD+7xcNJdmKRWP9If6HnSux3Zi8rsGx4fVBd5Ijwh6XJnaWZmGA01so3mswwU
aVpk4tA0p8Lc0Pyajw3r4VxsRwY7LPQULzN0nUDEZXTEnR1VCSiSpmnt3EML2ciNJ3zqLsRKwzLO
Gf+kxnzMyuVOMBbPJE3qtDmhDjjoirwaqh0FWLGBOvh2JYzP1n2rPAr28TnaWKRKfIt+SqhDc9dM
+b+IN2BLIefsmrxtXPbdx6wiluDyE29OYoQlAP3vg4bTmOWNb0jn8w/SYIFsnpi96mpqoy1tmxI6
mJkTSEJRA0L7y9PgrSUIRPkOP10MkgclV7LV0MEgmnDvUXJQuTg4riwzl7BOKlSRUlzPL0zrCQiT
wx3oATsVjTbr9lvgZpWx6QW8RYnW1Jq5XFOgGXBxFh2CBcz/aOmOFffzgg5igAyDz2RDmrKw5BTb
HJVfVH1J/Ts/V2h9M8IdqHGQuu9l/6QZ26GBeYONPM1DFBlWq70+EVfpKZXhewpuNzaMDRKvTHKg
VKimn7/1e8MgVjkQObHlonRd0MS0LZPec16hEc6+oBrTCfEFDU7kcdiCEG+z1xTZ0qcpQZV3vXLE
Y3ul17eYbkvho21THaUjhxwuMJiFG6Du4hpeKxHvziAlfzpGQSL8v8sOD84AOaZFwc71eWsPGT+o
qb0ISqv4esRKNWQkfiEmXxFfjVVtc5Nm+3VsM0qmq8Gn78TKFPtUCV7Er9e3UwNumqwlMMEdbmXY
KoWlZMU5pQSUHUM2YZNhENHezge5Sdsn4NZmqd79lHHjS67W5n0UIyBZpvnmv/P1TOEBCfYRSw/0
fmSzbjTL8MyJ4ocdCbtrnLnoUijpemdVkylbKGpG7rj6YHxjzFPyI+z1SrRv7xorOvi2vRNy8CrN
UFTR7al14mObZ0lJfHURzOCS6Zc6ojte+FwRPZolFdIa9miSwmQdAXhuEOPPSZoqhD+MZMIuDVvo
Tjzl8JafLheB8EG5IemJZv4PerXMtIhscFJzxIaroKwFGldDyu1N84OjqajE6OeNx4SqyU5CohHh
B8yRgTICaDK1qM4L4jKDCxFCicoM0zXArCZ1jl87Bpt7IR142L00aaUj2imyWJc8Uu8T3vRxh0cH
OEUaaF2nfH7j+gZc+4H+Mlzg31yI+aF4OWPZuTziE+zLyEa/8hOVNfc0OTUmsuSFZTpu7ESZbfZx
k2Km1bk2jdgDoePNCv/k+/RgUodY8yyYO56IUQKR+Qx/3JInnF6jitPiMNLuwU4AD7BvgsC7AUWS
Kuy/WCeUSroAdxxzeYjbLSoq2cb5FuM6dxHhaETzJi7VQWzn/JguQvENmiQaL/GMP9+Dhioavz3+
VubnOvNiLHKlzJ1WdzWUKdP8SemMJjLexhBDSdlcyfRVYbbp17FIRJzVCppISLFvU1yUQJcnG51Y
loWAFz2r0XBmfbt0tcaijtPmecRLRCin4hy5J4Jq0qbafp5v/YqNdrgCvj4dxNYuJs+ZrC6E280j
JZ4SWW/k4JtaUO3O0+VQZf54CbZrgOQ2sl2AtBESzxuChSHdVD5oU0ISj8hFwOvEko7g8mgWHJTZ
mHTwltHgaC6Ck4lHkIBQZXWhJaTvLT53ulNvTKDTNGVRh4sEF0RLj9TYiQM9qrb1kwkzhU0IBNUe
fagRM/2WZOznyHh2VfUuHfYt04t9RRiMaaj9mPM6qLfaxuMxG0MshB2fwdtKKtQUHgTQMu7BuX+v
xEhVwZZSvnK4oU5i2Phq9bu7HDKpYrZd/oqyoMkUN4t/avGr8yWSp6lMPriD98q16Ch9rYM7mlHe
3nYgv/6e4I0lgyU7tiNQCEW9XxFN5HqzKtByCHK2AcZzCUYQMMW65LwhH4SOX9JbWeWNPW63pOzS
232I6dG3T6lMWGB9nAiSPLr+XFP3NEZB1rfUfU6WxOoqLWhjN0dbzZEqTkysHwJSwm1FuP//VDGh
CkTWnI8dbt5CwNmc31BqLocvw2QsWMpjkPzjhocOgebOdOUq5H7lu0Cf1Zw4olJqV1GxR2n5O62T
41nhn86a1Wlb2txD0y/Pgss1+RsttFjxEABP9FEfDlHFEZbg2gJgVEPUcye4Rw6UH48IZve7NPZU
V8ycGIeYw7nyHEdPTxeC7tDhj+Y20fc55AU5R4QRbORaRq75Mik4wdXDPXBUayX9NQi10jFhNro2
YgBZWN9BHx3wLzo1sdBiA+8FJVwx5MlREwECpYag+bXwAAbg8yzJOpZSLYATRNfqTHdtsJvEKPs9
RBd2ziWaI6WyBYGG2tqVkfRkH6Dx37hV877VI6VrZaLqmNGU8qv6yI9RpVxmVwpwGSFRB6CkPb62
lhvQfDURGtrfZssHborXpgn9wwuwwMvxXslcmLbgwVozo1VLyEcZohnMLA7NOBaAM+2t9CJ4fL9Z
wMvWTCsIw909CrW9LZrlfXwjdp6YlV5Yajv13Qa2UEmwAiuUZ0KyntmEIXJm6cDgciC8LcmrZQdb
xXxtIXvrP5g8cpv56dt35/lJnMkUg/0d30Qo3fHp4ab41qOonYsSnAauUxe0v+BEb0ifatjprK/m
26WiA67sKwPEPa62eqskbrlXgQUvsbOyeTOEJefYiP02LJIXzPUJZe6vmNvz0D0rMJpjNVZMvk5q
B2zB/QpMNWIGDKJT4iy1pytECQ1ld+ksjire6LKb5781N0PrT7w9jxZ2uwRrZdFX34wlhxaAqBhf
rJUBdHMyclCp2L2w5xVt8gtWCNnbgNDsa4bYiVAMmGmDZufj844JNRgEjofrFbDkkQ/DfWOPePl7
71EJ+W9BmW0C9U740DBVQtotwOU+NiahXt6ygys4q+oQSE34Viq5grBmzh+5ziwEItski3a03nPW
hCeOiFGE208oQYiDbwnCawmC9lzNWm3X/OmfxZmFIUs2sHE7SIcbY36UiuWTWmHQgrgIsGXbA8Bp
k4SjNrdcrFZSWBIIrtMgjHES6rOlqDG7VAz0COHvWTmeRxJlSyJzgLZTpFZoKsAYOjDzg9Gbh1c9
3oh/DvmJjot8Qx4wiN9cQtutyvw/hYbYgrtrpyxUBwIn6qJcuykf7OLoaPq1oaP+EBREWYcrEETU
dOhujs+OeVHLO6NN0aDEK9NHKmZKEwakGuBw8tZ2FkRkcxe0vhKsbstZgDflvdmq9X4pNdqRd8aR
VOLna8mpdgdpBDq4cyMuEMHDRfMgc3v/T/rKFgaCFm0ZlEL13crZGf5YfPsNWJCxY9oLpOj54/Pr
NkiDSdGV9940tOFGNLZ5wHO4eJqkVW8sEU+D1dEX4QXyZjB7kqa2dWt2/0HfP8bgd5PKB9mYYJXc
ucFdJSzbmbjEcyXxF306sLcsgA6SaysiUFa6crSW+QkYIGeF+CC/Fhn4ysPW8rLJf1kegH4nrOJl
R4QFgTqE1k486RWEfLXZyW0lVzr/NHTXiIgPmkXc0nJC/3BUxBQ+M9jgPFkAiCME63hM0CMVRA01
MCQgY/DgnGGs2uJg9llpz75VTS/TKf6dnpEq/URjo5SUnzMFtEVQKbmdmUaacabijjqTj+VLUPyo
IRp1yQ9dxFnUE/2f6+Iu9nxnnbF33V7aM4OiqzrOwXCCEEoTXiWRX/W8q8raks6DHo7bx+GvkV4w
XgMHtxBadcgsWvlminwkL1RwWHm/FEezFOCe9WbP7Pgx7hT3mCaKSg6XeF3qOTVidWUsc+gnIwnq
RkcFO62HdVtRoCN8+6az3YZZwK4DRZS7bzWseTjkDMsrSd4bANuGv0scEBXMBMKBHTM7TYbEF4ai
Nd7rIueltZH8157u54YvTaL7lQSjCO3G2QZ4X/2muAkU38D4WF3Tgh2Cz8cIhZSjuPANHDBoeH3N
ynorprQ+HUp/X5wouriAYdKPECyZWNSQFY0YzzPuEKr/T6WoQGXokLdsN5IkoZm60Mci30uGxMDy
Yxqubel5eW5y/X8m+KKx65OSwdO32OesmqU/rNVQTmspPvV9qvW0JERRseThgRiHFEMNe9RghHVk
wG7MJqKbp5TDFJMfYCxuYd7cJ4cyrlzBWLfT1/EslOc32A4N4T/b70G0rr27L7JBRC0avqFaH/BO
0CZai9YjYsPtKrnPFdR0egXuk0ybFuXnwJuLWod89EF9d5mcmKi9O2OSoKDVTDEIb/BzmplDZAEE
oSGDOgkct4Kd9hjSS3RzZr/WZIFYw5AvCoRRB4tBTLqTHJikotTc1SviDVrN+Mdlg45T5uZ6qjh4
dSd0n36IhglD8TmSqpuWpEzGox1qg0kU7OjvD1KAaMKYmZlGlY09h5IevMXrNDESKsqZx1SPWNi/
NrEuLgajAVnb+407NofATCLXL92KlCcDWL7D01E42FVNbcWAvkH+nMfh/9+Si9QPCeHLi98YB4gA
NbX2VjPDqVsc4yjlLnH4BMj12jyg2qjQGpD7CIQ7HhqdRqyycTjYIRdtvtbNOwqdvrXFrlUl2E9P
M1qVqbioLz3d04TP//d/4Y1ucd3w185Pkamie9eiEqgRvl1bRhl410QyvIq6l8p1vTHh/eLKa3n3
jpNJHcMRQQXK00+q9wUkTAYxDejasCNy2mCxYgItJg4Y2QAlIqSYOxrd/lXWxosZ03uv/GDCjqOR
FqQCwFFDQpF5Nw4gWHBiJEzYvvBdtBFokV6ue5zGtHxdWGzzxlPlQEzQbFxV7iFQyTmCcztLsZh4
MDr7xcPbaIN4Qb232qdmY0lrg3ZiB+UZlivT46DrjxG00T/+bUT9BCSYOUeSoPruwgvZuIXSeyD4
HlCFzVMfkbhCextJ0PwrZxnEwX9YNLM5GdGCyw/W8yuYIN6GwsuKCqxc8iJmWp4Zr3jce3Chuohx
ayBtvypUxUiOekpPBhRKvYqIVMk3gMjx0KWJ08ZSGJKUsGMOEagOXr/PumubKxVqN5RHxRh2qfdc
EdkNSliLBIy0hha+THuV2tDAmgT6NDabWIjLDpeJUCUV/Wdzx7KSUf9zyGW9kF4lN+WvzChUGrcG
/fNDxasYcUm16rVzR1B6M0YumpicAn2JixWjiP6WOp2zk8gpnSCAC11DR8Osfo+NTK/pyLC6cohX
tnNyS17mlMrTkDxlSUb9hht8jIOizclTAAixMk7J03c7AZ0Q1UIiSV0530yr2UXG4VK81EJNvGmp
th83/7nXZg9bjZ1aMKD5+sZKLRzzKPK3oz7uvKniUes3BqBTC0Ps9wBnyYXc3/5fQt0t/NmODD1r
RafPqES1TwdBGE3zkMXmEFlHlNP1Qq4T9wpVIEtqlNot/oMvaGZAZQZLqZw+fHjhVaeQ0dx9gmS5
R8Oyh7AhDCXNU9o4iUkeHkSaH7sRRQKhnONw02E5Y2WyUn/cg1Qg72aTcLXdknL7ju8CMc5EIBVJ
zYuv/t4br2Uo82bOZ+o9YDAOhm4qt12nWmlTbfKBPvMsJ+9uaReixUK5ZPQoU/ct7oukIyGTc43k
Gzk5lRinjoW/OQffJINRNuBODHl51JhcMAxYauZ5QuKgDEaA4lw1hJLvyqqvF8G7ZSf4fyynqIdj
TMvbfqA83rSx0I2qSSEE+NLNjpp/vh6GyXnbDNvjsBUcS/6KTZjLrCZeeKNLNqPqDfzd2o8xAIWf
weCXWNV4eLg5ZMdP57IF/fqX1xLOKwwsh4Fj3aemDjCJj9d5qsxxDKeadzKLYGxM6ptT5VZ3z1mF
rEDt1r/o9ZP8exB7muIeOsv/F1usDuBbw+YeRNgUuFC7EV3lKAIFyxSMW5KFpJBtndsVw7Vn0F3k
WRyCnp3WJ2FafFJ562xn/pz3mv6feKRGoad561mK+vDZFRtmkVgQMmWfJKXCNCZWpL5QSjDlbDTQ
/ECq309K4zVl4ZipV2zEtptOvrt/d2ytukfzOwW6PtUQikae8yRaZ/ryBc1XQSgq1Slrl8z2sz6W
DliJg0S9FOPAvh6U2TNkzkvzb2L4+Q3hZOmEH1od8JXDalCuU3QW+niq8tbFg6MbchGYkL5OwBtI
HK9own2/8HXT4R0gOQ2i28d3Gy0TdnbHuYSb/0FNxz4pb1kap22cN8DMIlQZI3lPfsQCSGGxYXIa
vbezxWJPaWriJCixtYDynuZG6XLUIwnFnGLStssFMa/x8ElYUWjWJNg+rZ6qFWklDX/y3CEUuvxb
aB4SxyTLz9CyxkzqPe2sJvLSooPq1j3ZGJ9dD4OmY2h7YEZGlbqt6nT3WjO+uLWorzUYXt/kzMev
bWyyrlrcJhe9dCW6nyH0DY+FGtV3vFhS8D5K2DQojilEpSWZ25BzcNg2DcVKZbbOxnK5ih0T8AJl
YsHJAz5wvB7E4uPLFmaNdMgnZNNSRZ6k10VxEZsAh0X9ldOcULBzJMdXpLbJQvVVEST0sgnmjVCC
TQMozmmJL4D2pa7TdxoGK4rZ4FZXbE04rENzucnLvSV1x7OpeANiqKDAl2gsHVX+RNb+HrAkCdxc
z+CsM0096QXiJIO96AfeDlDn3EOzmmpPj14rFJCMwTqh/gkM+NEQmi9dDWasi3hAMf0z+GHIwmxM
DzXwJjd2mQ5jx+WsLnc75xhXZ/ogPi7wk+0WaV6hDIB7wOQsXMrMLhEZoe/8J5jW4wj+ky75YKDV
NQo+TxmxDbhluNBliG+g+D1VDwxHTuEXi9iZI4YR1pL0Ew/s8T7VG4ZWDosFZ/PF0Zb36zASjYWC
isnNWe5CZdtDqk4RAf7XSqlWRNr2z8bStwPzsgo94HecNsRHHtjBmxQNTLTVuvNS2K2HX4tGY4aX
1UmGyeRa4G9z93t4sZIHpr1PL83r40IeSUTQTYcuUYp/SZ92MjXQRfO6xbzC8JP4B+k3d+mKVikU
g9oxSMV6s6jD7vmB604DYfi/nxfvdgOZ5klSvQiqkHyYCgf0OI94hmwmdm2XF8yA8OwtHpaRS34k
hh+put3EkJIT9vSAnU2mLYxBRyfKDGjCor2tZ/8Is984bZ7f7KMRfhaXlVU2Jr8Ie60svZhMRxv1
9MQyQEDidamH+wNZ42sEd6I6uqXklVcdJQVI06vMlktrXU9VbIK74tkOJ983DyMUN1mmB7evs/U/
vCLruLaXqHfWPHZDc1vyKaiNidfol2H68hf9AJyKYGvUR5iMwyOQfMyI9NpEnnywhVur31VW4Ad1
lIn5raFPlne9tW6IqDtfSvDp/d74jTmQfXQGVIcqiJVvpgAJboqssQVqNpw+WGO8ltmiAq7a7OFD
mu20XsVWk+0epGsn62gzWWaHNe0AR5wucm3GojWSUQbBMz/ZKaT2nV4B645VffZR0Z225vyi2Riy
JohKNtnA0FzbLM/zFxUDujTWJKY8Kr4unoPqFIs39VcDgGi06WUFkokVYD/6/Kclw0YgJxsuuV7/
m9OldLJyWatYvSqNEyw3z88YR2q/7HJPi7vfStd4TpVR+wIAoGC8r4rnk9DCy1/dHIWq3zijYQr9
1kFQhdDPcqZMd3XFsLpIFtiFeA1mz7NsdWmKojNKDAMXUrhKLSSiL3D+WafnvuPUFq+ksKLEdwVp
HAibMm2jzvhI1NN+K+BjvVUjdQ5mTJdbnvK3J+UOUVKDIHVzcc7IZIAVVr6b3Qa34YVRAOXuV3dW
91k6xXmWNoeDI4mFL+xYAbUQRfwM6n5kTqw/Mb3/LCK4IEaa7FyhtDgn5+2jgZZoiWagWG8yRHSN
WsmwEb9AzIleC6jO1PwImFnhKYTpPB/nxxGxCa1WmGgE4BwWKYg2vLf24zy1x/cCMtsaHMFFuvjg
s+wF+6jaFKouIQbC9K9UJ5+TGBWagUc2SxRqQ+SBhgz7AYhNzlZ80H4almvcOOMkNrdMXGBHpgxF
My6nMFpPUvN9yr6FPm1KkufDrkLHrdLlLxQekWH08JJ5H3q1eXmBCuX47ZaadkW/rcwOwqJKWG1m
05ZS+1+KLClQfADxjIThieONnD46aao1ZzxVx/+4/8YVHNrk1KNTjo1m5wKWpCNv5QaazMfGCrdd
0al4lz76j6rU7TD4cSqWz9Mc0JZ0xuYNYnn5ui2L7KgWtmnglZ9mm1N48tcotaBtO9DazYqJV7Se
XaDd6wnNDDzFeJuajHIDNSIgvzGype+aJjk/tCgjMMvkcYWZ0mo7vaB2iFarc3HWqwTrDzsKKsgO
lzUJxCQP+W6W5tduc3nDkwMXFzAkvr04jKYn4SKOMI+zEfaqs1H0sAa2HZLqkYxqFbCVrawg5mFL
LiTBzWB8QAMPWboJtj2mfPinbfz67gNaUb0Uzt8YfcaSGcyTyipv7CBZGkPwlTGHCu43aMGIyqWj
lIueYLFEc9l5b9H/8y/R6Le3Rha5BANbv96RHHs0K6/Zt0qQnIhsQ+B2QEipN0Pzg7DoJLpbN6rb
na403O5PrpdIFWLhP0hxBrUE8yxO3whBk1fF9lRnsLQO7tN05nv9bF+FgUF+DfjpzuASaGbKSGz4
komYct/y1QWdSa82DAkiJ/D7jH2At4RYiYXBCLwBEWk/VuKXtYFZ6NG6g5l37wvJePiemzj1ZpM5
4/jQwvFQmqTsCe+/khGIt4s1zyatzSasNsSjZh8hVzWQMoseZM0G2+JGbbV7oMDvmVvB8avpuDq4
O2VRGs95dbXwFxoOCi/Xs+ptIdF59sWaYdJ8ETPXhaSwewPl38okTGO46YVjdennCQcxd26E7RsA
t+WZ6NhehbA8zNNnsV8eUnc+CCX9ivmY8MoG7mabOdla5lu+YZZyR15r70X540sjlU9GUnb+RbTO
bATatBBqsXvTtb+EyG+bYayUTAlkHZUDvYjtPYQJn+p/z42GTrg4GiNpoIthVLZMNqRPdQN/R+/N
Guk0AwybAYmTZ7/Ptg5O+KR6SUhs5ZS6oNncJ3M7kdRx1w038Jkx7OOwA+1bDchKdIpLTGzFK7qu
K6kwDU0hCEFYJx/jSqlv0xpuyTg4PZ+RIcX4ymjp82R8Z3mCE5F4ZBNAmg8ZcEccMf1WbaLqpG2F
TEhGc+DlsI58xbiV2YZmtjvSW6K+jQcsaQmA0qP6+xbsizCdJOqrng+UTPR99b21t1TBFQZyVpNL
zxq0LS9qDcrZuzJ6hLPIXoyX3iOCh27BHr6m4wxXmT04frz+4+JWVLJgbMBbPX/AEKDL9WIKa3eC
9q6pR1KYYeea95gggS482OVinIaONnyRJumzG/SOcWRLTsHVcdluJb3w4BqLDy0rB5/XRY+xtPds
pe5O9+drNZ5YlDrssyZsmzmWd31M7ZltEFTFcRWaVmyq1BcUToqAzhYh6z5NjNH0AlAJIyKNCFVj
Dn1BqMvtE9ZqaBp5KkHbjz5XFZVhF9oMNTxSmOh42J3/DVavWqVL1vSIIIAHGC6EaftnitSAiaXl
OCl93fh/c4cOEdSlWD58SX1cEsGzUT84b2E2Q0adt6bTDzd1h9SQtJNVk3lNq5QKORWif5yByKK6
f6J2HC9NE1OOvu1DEfHIjJ9xyqq7kr6ZWUIo1/EW7rFZTkUkeLvRlitf73oZBCVNexvLw3g7Pxg0
9IJVtsNp3OMT6VAlTsONOT5PVEpcqM9CiNvRDcVb7mfw30irlfbSse35N7y9f7xH44vtbaD+V5PK
ePAfQ4Nc582dmojMYPihflRKtPYTkwl0ezA90cSiqPLSsg+gjyLLhzBYzHVLXS++TmOPZ+u4c/iB
/prFJBBt3Umbm4I6Yqwj0LtJCl/IUAuNgP9SwDu9jvP8UJUQSqQkGPEB3KPVpvRntf1t2cmEqRrY
xY7AMH+qQG5megOsdHMAOEdFeNpyMiLdKKNqeE3dziw+8vWqzP6vpa0szSxvHdSXbJRM8raEjZfo
RQjQXImCqLAYfVh0XjUDnTaKxFE2VB0380RmrNcSrO+O7dYYbAXgKG0JMTzt9MJ3sXJtiA55pj1r
V1JqR+Yb65zzaQbnjeng+vMcWUidYBvb366b/h/wHDFAVMUz6dh7pMrEkNyb66E1YCvHHbCTOnFS
gPAdkWa+AyZql3YZcWbBOxDNbSIGMG6VHBPyb7zuFUQKfxyDc/+zdUp3eBib960mFcvPkJyq4vqs
s0OKWANygPeRj6hsHQO+9YtlkRQ7+u6ckW1cXc2WFr8cHKvsf7WX17VClZcI1DRwD8mzcsNGksM3
GMX1/aYJmPb3OiiLOe3oD56ffAFa43M+PrC40pOFWsNk5rsqhpyoYTvTUEXaD0lvIoYpW/fMc/ct
1VvpYf9CNKdtpR2UFDrXm9Qphu/dmemVjTYgE3tAO+3YqM+xJI8Ltq/RZWzISa31C4n6FhxBHRzT
5dwTFLp5Rb3Cd31yhSI4u65GnKK0T03yMMWrqD6yx8WVaOYi9bM9+QCfHP6RTMRUjxmAY3wNqdXa
QZkPIUUyjjJtfvS7F9k+eOxiloKLDp3+bfvB0bWEdYPOzgX0rjd3WRWEzz/kYk0e8M4izQm+DpL1
/MJLEAL0VEpv2h2ItATmQUhadJbTxyLA/1GkuF09duO4Dr0zNDDiHjVcIwo0co/IU6WlDs8/J17r
kCylwstQh++qGqZwvQlMPIU2jISZ2+ifEIeVKbRr7i+KXQ9k81PQhXt1tPrV9RIphIe32YMOHUwn
uv7+Z04Ki/bZ2K6EFjiA5XUEBH8LAXfwwrVECQtPmE8e4e889wTT5dPr3oe3qgCSB3KZ5rmJHnuD
Ve89NfHat8dJuzff6lFRTPfWTJyFj/8AmY7VViAcEJfryYT+k5FN4eyGocoLJMq6gRa8qP1CabWe
odaZrfSUb6yJcXfbKvOduiP1Pz1RpGYV704dPMdom6VfPOW8d0RLOX3lN6Dgl0jR4ijXbz46N0Kr
xWe3actOcas7DiyGgqbU14Fffnta40i8ZvAB/9vdJvxDjxqmUmoVGyMbridn4LOpc6bsEbs0dnME
ZjLaRryp35+kPggJicaxtI3boHcpxd0MoA8b9hsuLkNfxMfeE/KsyDZDZQQAD9kYJr+sKTEyGe/p
noC0agyrS6kf3YZXBF7O95Susa4pe2aqVTyJrDoBc76eGycJHQwAnbMjYv/k02k+5JkRyAUKlhF6
FpiutWnxx/Qh4hPZwhnchZalLmX/TITrwJvCieFoqgkv+0/MJolniWd8CHlTHPTIlZnvQ6jVSuHj
GEYD3tI8ZXNkfs2U4MAoukdfGLB/V5UMuYNo69FxtmqsjgX5A4slRmMO1dL3ieq0Ny1pe+apPztF
5wiLHuEQDXEtYoL8cd4OdcCj3INh2G8fXxiDkkVnCMElJ+jMMpxv3BAAhlmdRDJJ96DDIoWgvLas
HpoMvh/OxirsEYFLlfLWvuhfsvyZ7FNdSjMiyHky5ObQLlvx8Zc9dU1Utar4RozZEPDRSohWj4h1
FdkLj15HX8C2yhUaQ7rsJG0mCvcyNe5tIjOCthWGQ3fJF74Y1yCag5AZiSKXv8f58V6LRwZswBg0
qaOHqeuZu1Rfj1RIWyd6+/oCw9rtLEh/ObjrG0bpiIXFuac+V6bhUN1QDou0D6RHZTxr/tIC7tNI
E+Cd6AETIc2KDpUk3Xjew8eLjnw2H94LXe0l+hDTZEnMkG9BbdDj+xCc/bLVlCOh6Nzf8Gt6ecYq
8kyreHeqhiEAbc0P/f3J+mOhJL+nbA2rMcd5EsQ9xz7dUTTUtWquyQU/EGAeynHEGvy/nD8Z15T8
IHWxvm351U3oBcx53nMOFyx3vLCALKNFL68jGcnN1Qpq3rWGOPyj+7OxXiyMhFjfUl5gPdxPULCh
tOFDqeH9nEsPUwVlW92hgJgPtM/muQIzp/loazwNLsVj9M2b6YfZR16to+V58DCzo38SkhHUk1d9
Fd+6KnuaUSO9KNReCD/pH/OSZly0ngWBnoFMHbOZ19SbLixBm1Gl1GsvwxEPWxBltb84h/bBz46J
x+fj08jCrD7P6f/IhFg6WVFhS94jogR60wQsErZjJ4zgBSIk1bKzWSkvEAHIIno2n05lVN1RUccc
34AQgzRX0Q9JgrKURaGNskQa6XvipcbSSuEBAonC7BvS15B6EeN85/3anyYrI4BI64tGGJu0TfGr
kBqpnhIXEBb8TzQ53GBNsUxj3rmHx2GtmQ0SIpABLrj7Yw99gA2yNqHaqxcdv2ywBm7VExwae0O6
084lk6yOuzuz3hNdDK77Xiuupxq5M/fzqu4FYhkjtUINIPFF+701lpD7rrsQ6EEp38KDR6gK3efP
f7fqMnvrg7NfJuL0LpsphY2TVZj3xL9myK9RNUAxG78irWYZAyATUxWF2inDAeLlXMG8zvLfkVkH
a8Rhf9Le7+/B/XTFjoULxr14sxB3GtNyv5onBJIbHU6wrY80PdhoSB6ya/reqJsBaZ+AA00I5LL4
SphCTkGhPaxuXi8jFm0re1g+apelBL1WmByqC5rXXBUyLzSuZzNfZfeuAihYM01yHeINbIYw0Z2I
X+FbfO08QTbOWHiSAcvIPuNYJJeLZaMt3YVXY14Q1l8+hL23qVfXkhTR2Cvx7e0qx+wM5QI9H6M4
zTP5akOVhnj/pLLJSk5QyGRJSSX8o3rNvyCzOQBOKbLL/y8apAS8bCB7sBcBkZ7q1Q9bT+PaqSKv
fuAC4B+ToSvfdmAhSrcgWfPxx1Q4oEi163de2sheYfpai+m0AcOXcr8QVSWsgWkgBTbpaWARqf6b
N397m40Yv5k8fbPMRxgw+DqwwKKIR37IyDDE6v9nqIpY1brRALcQfODfgEA/MinD4gfgU9LRbr0D
tzwE/l3qp110roRrpR0ElFgV/C5DYCHjLH7bM6HLzw/9IGf6dr4Q3tP1b2ifNwKT33jeuk0l1YOH
aII6udpEYkY30/uDaRQkc4KqB17Bv4Q6lh+5xmi5SCcEmxj3rlPljxQ+O7yY9GGvlCpKXG9cmsZV
SW5YVFVUlQDrCBxs+AeB9f4Cw6KAn6xq+xF4mqZ5JcpKDiZUwI2QWSs3qp+R6WKZXaz9BIj7R7m5
Qnm907RR9ozSc2igiUYZBAK/jTb0wLnys/ukufMNeOX6SFZ2txeJOq9j+4Bat9vudrE8QSWJn230
9DJ1km+1Py4onBsaG+xb0O6S7FOAVaUIWgSsMfOawzk5IQ3Mv44bl7ZMgG8T/BfYhX5eLSQ0h5ob
qVUG0VnFWPS+h3YsFjVxx2GhMJPyjQnZkORCLryppuN34qCq6aNMZR0SNPqzXdjArGrOIvsCG3ui
Va21i5slxrU6AH0jpAR8m3bMJpInaMFFswJxRls63CIFsCgqDjUd9Jtd3r24G0aA21d9IwRl5reM
/amqv3oSlyu/hpBXtKgfsQNBzFzL3mMDyPp3xucMd5leuytlZ3CZSfjnWnqVr+mUBRu9jko+4E3v
oYWmazwG1w3741CdXt4PxZ1Io+n0PLZnjD/4Woq8eclDhkCc0x/Kzn7dR9y7WAwgCp5g1Y0NC3bB
pfdIWvSbcWlqThQHNyJIdZ+/XQmmgKRMA9JYy/guvpmXt7N2qS3jIl8XSY3+mEiz3gxdM2ioNHTo
cu2jMzv2sDEUE5y7w+H51vDY+TaoOTgGdReoDEEWV4veDP+ouQOQfkwKTjKspePH0DRt8TgyJCSJ
Z0epA7pSWx5eKqp72oUV2nrmyVYl3erwiu7yGjXXTQmDLo5r0EMMGVRg9IWI8TzAd6eg5OKLPVd8
lSUesYPmao4lhkZ9foGqtBFmjC0rMQKROc7nKGkG6swjkpJ6z5AEgR1wdmYqXyb4t+vhTZ28Ng3I
Uus+pxQymtRvEfqT6OrkOgQmFot42rwB8UH5ouUVvSYasQF/WCAZwEMOqmMJeanBCl5gluKk8i+L
qiGzzAllGGkcZ6JK4fUUlc+fr59OWO2L9efdauiNdiAOEf3xa4hQr9LtZfsLOer9yDntOOQX1Um7
Jwe6Rfni8BOZvaxKY3lAAIUx/TBP13HQ62rOc6vVoKYrAkrzil8CCBBvB4b0wCXqvxk7nKIk5HOD
x+RkFty1x757KPaeN1nh88OjTUV2JqGNlGl7QfgN0df0at5Y3xewfR8Hy0tub5PmED0oisAcvpAn
ae5dXuxbJGH4+DIYXOqkGDaHpKFASwGMt+RIUlY9jppnvmEMvKaQXxjHzDi+ZcBtD6iwyajcQgbF
vj+Hn4F6pXMQlRS48oGZiiRPoeK5PF5jE4jMY54THRbsEV4p0Av7NhcS5ladk9RZap4dBVoLRYdX
wCKVyeP3uJ7nl8bbfMnJnGzlbL050tGVye3S80ernVoNF+lOnl40TM3mWwD4UhIf89J4wtgbYoAF
1WeichkTh4tplXWC5T9vJpw00bs2jgIZRV5bD/6GhQRuSMHEaZgmCndgJhzkCjSp6ummWmAyZt41
6VEAtbFMoMBrVxE5QANOX1LDUsly33RlO8rze9VY3L+aaW7vud6Vj48FfqJNWsZ1G+XhybCPP4r2
4h84JwU77+suNYuc5m7uMb+Sr083mq83eawlx0X0sAeIH7dXs9U339meuOP+LT1q65G5hasmPm1K
YLwGxkDTJYTOCJYaRN6Fh/CCNpaNuS9oHnM3C3LsosnGpigVpAW21mprt93PhnksMXSR6WVp6/J4
hYzHT01oaZzI9XFNTjCfXyDrLa5QY9n0SKiMNAu6v/5ydVQVk0TCSkPxvWrp8TgV7PxOw8v9CiHr
xRY+9cmdkq6ZWBjtZRbbS/GRyMtFte2yMraZHOipI/nLZKIK9zToBhLo2uVNiM1RaDdGV/juBrtq
aupZGiHuRnwpAO9FXhwDr3aIMYIxeBPahTow6Y/GJGqltpfTupzrMJgj3WTedM7kCOPqqzBe1ofK
GDoHNc7nCdXmODEnctwRjEnqDkBJ5Gah5uabZiWB8H5TwlrxrA4zHJeb1VPPgOutJUL3/v6IonLW
zvZt5gogz483ZL7E67uQY5Sh+I/+EG3nWiqyYbBznNaKdz2FZsRH9TdWy/9EMTwZMVc4hcv2ZL+2
l1lYudg9p4PUMNVXMll5BBt4/AFBvdP71EofqWoqFpzBThQpfH3cCSelbKgBTmGjP8OjJ6ChNHsY
GOtPjcmmYVh3Y95qoLK2DaHsdYXsXAAjfEzaerTf0NhLirHeDL2mRDL1rOA8P55G+fKL0t0jo5cA
VTlV6/c+EMyauKvay7lLsKyTSYttN94zQ2aIX4zJO+SISPAIU6Pf0TOL7FB/doEYNs4pJ5Btj7pt
aQxdwJzqA7C/h34rozazMg9k5r9JvnCgrMHoGOlN72Pc/EG1Jd+3vcZEZDH3owNg0sO2GUs2oR6n
ggxyZeLhBSzNwllTPyVZDELXeMzaBJnqjzeAr4Mw8E/HdyuJRCt3C0ywKyzvOnCAaXkJ3axMCuew
Ut1jbPx1DuG1cd+k0nHrVDNMLWo9uz0oWzJKlDKCT6CLLW7HfjHatiOI0PXVUjjhHsZgWtvwt6y7
Lwz0WV1NRt0nMYbVSj8CZhcUCkBZKhr2gIVBHNMOI2rQ3GgED3NUHnmP0igExCHHzCjGaBMfb85w
UZDiYQmUZiW+xJ0lBr4T+9RN2sitbPJrD7/AgurA1xS1zZBhbA1+CkHHGLVba8l67qdjNdqEWiyP
+75PKFrkV1oJKCHT8SIxttB63bfNAkR4COFhg7viyE5Sf5XVOU5plRaQsktwmkuPpplipU0qXcH6
7cyJPsNJSGJiQIp+rn4j+tWjPAsH9yAVJ2EvAuFQIGv4ZU6KSMczBkUe4u7DZFl7O06ls9YPt/LM
KS9ASdug/hoRqxwYqJWyLPBrvYp5b921oq79BP5koQrLwQ2uGDVqx/DibPiJ0RGij2rM3UL9VAgV
CEeQ7Av9UfRAUqBVIAnS5flsEQ0aHLhzVYU5vuNYnPVUCvhyYuNc+bjfwsxj8p6c67zeTEBCWQeS
dAUdFnvbM3Qb1YaioR+IqSDKVdnIs/jsmiVTB4oKcABfti+fZgXb4aHGf6AASRtvBH0HbHM2RwHN
K54LEiFC5lkG/6AltRG0PcCgoJhwEEG5DWmXzwMokLvkEBGoqDCyuGQWrOUe0O45Xkl1gpszfcd2
Vx098tX8Ma1vkkuFx1t5FagUnN7V+ikDRUo17w83dKP37EAUNOmXZKmsgIiLLkhBZq7709rhWAl5
BODpfJxXx5jzEOHqj46lLJvMS+fGfjuym00OivE/juVD8PYmBqkshxGrL0mlhnoqggEv7R+GkQRH
BGSeH7jQ7LdGL1aW+8JGVbZUZJTouKwNqlvw2HDjwRABDtwFlsQf2KFqMS0878rT3kHCGNFrmgHC
9GWyU9Rncf7miUur3Ao2zcSdxGUfxoQQpIEMnm4JT8Cuf6msP/xOIuXWdlpHR813OsYvGzKzKrz3
VyHNpKHsAG7xZcWOljjJ4Qe59DIT67nbPS0aW9/uVPsD2mNyTuyau48vpDpKUo+HJDiV6dBRms2J
Y3/9s+PfiyfL/f2f+wzIgn3MbKBXRbUVv+pVwT1EodjdAdP3HwkYOPPLPPISNRTaIsOmX84JtiLo
P8CEabhxTU+U/EtNRjAMGfkaTInh3YHCskoCohdUxD9aGJs/pH7lVvsPdNxSLHVrk902kU+1/XvN
qcG9gGCPdIZN49VIt71RBEpk//B2q2pwZDrTZ0wtsCTjTtCoY6LI3P2qEj7uFiqfJs1D1FX93FlW
eIy6UH1gXpENDGFEQd7WoGC2NQRKm4bIY6/xQUpvUOPQRgtYrPD/nrJ9HG1TGIhjSPeAUuZdFKV6
VMB6mob8ZhcxNCZMi9hSteBhD47mxKhSlhtrHEmTdgX9DSvdbPuN9JKotaeA6hfs8TFdPe8dXV13
hmfNCWjHGPTwIZDMsEPAc5a/JmdqvZAc1L0B+w06eG9h2HOmvZ40+mKd/Hi1O5ofLDJkgVE3FGLB
d/1ZBoQx+Mn3yVDQH/hjojh88yHrsDsiVQdAquR1w5qC/hH0YDT8WIsI8EfJwRPi2daH4QXvUymq
xcq+MAFkoPL3ysBsgJwAPmVSuvxTf5hHaVKEdm9+FalLfs/R2M46Uxx59HYBHFtS7f4+uE14x6wm
EsBmWbN8AwiPqVbJBC93ST/VeX15fyN63mTirTbm2jgdsg1S8iMHYpBYNQzMQIz1X3tQGMTFNl0u
fQma/M/5rdASRBmQSufZg50csIDaZvgV/b8UsUSnHn8YxxLDVAC3Rc3rSnsvFiIWCbyCVRzRo7Nf
EEKV0RQvl6F4cVAuN9PRJgrlQqtbZf7fY4KOU3yV6viKKhvdvgUrfzhtqLGREPLiRKgMOgzhrYRz
tKlwgr5hoh9dV0G1VfBQ4bmpjG6rH+srjqS9jI3+FpFVguC58ldY+Vs+xpiAJm+NjRSLEQ1rsWzU
ee+3hYmPLKH9vAjoym5IwnNX2O1jZKGZU+X9nFDk6pyfyTG2oGi1Lu8NaCXAUl2sSv4cQQzq5c3k
qYYc3yuRRdkonAaUK7MeYq0jjZGTansYh0Vpa4FzU6n9am5nVEh/SB3nJtB0OglHmTrttqgj27Fk
hsve2ST9AcUnA/YDkdB/I4DJEDLuWHVxI042/1sy7yXnC+MpoILF8Qi59maQfWx+QG6L3IMI3lzX
bOCh4/ab+uOX8wcvLv+EjZt+3emxMaPh15Wn+uqepFulElC+f97lUhkcYbOBXXeU75hr9NWPAH+1
EXfSW07bW30Xxlo3GeCGIG0bZ3jb7dkynsK4w6Eju3gu3+T6P8HE1ZcVtSLcwzsaoS5kWKR+yRfQ
9ePrnfn3yrVip6/UvcFxfAEYgFmVviY0dsAvMbNxINN1yy0l4NcIIlRtEqktcyWi8u/grEJFilHl
QzaACj1xRVZxFnHp4f6/Zivv6IYh7+pBBGIVI62NTsBINaWi0CyGBlUYGO87T13HJRdK2pCo62Zb
SNjejyEtjiOJrsjFzhaaccV9sEnQTkYti3rAHbgJ2ovV5RcxjhNzXY3Ok1wUspWF6N+8DpzWnOFx
VXl2zxDtpsdDxOLS5aQmNKa5DU8cki41y7H6LcuSUQjFZI2srOPcTD1haSHkGjRjfUuhKis/7696
EBG2F6xctm7iyTHZNlcu9sedaDA5LQH0/HKX/uK9HZQA3jndc9jp/f1w6/TX1fiB4Blf2VUYq+1x
PYt/jNyiR2fCYAIq/KcwUnbPGiDCthDHrgsOxLS6+u8G2Mg8M3Z3KNWcurwcEOOeOM9aKsmM/kw6
U++1gJRjJ3Vw2EjhRcUbD8dHVPxtOUTQDdXwMEz6nKOLX3VNxB6XY3UgXzfR7LOtfRAQL3zzbSbP
unK3DdIAfOnvbJ2F6lKsT9oJHjuX//kVn8+/9pnqM1NnRItD3UGo2oKVIMa7sxBhQY8g9wVK1b5V
U3pN1TIIxIQdeQ/stDMbOR5l09IXXjAYcpqs798r7qH0XVYjV351ccz0bpLrp4AXHHlquNo3xmTN
HRO+ro2Um86SDKyND0uifwAG6H38SzwiiV/HY0ZWMV9Fvolp2RjOwuIab6zk7hMWj1cFrUuoxV+/
Qgr6N4uxvHv0/h+0cZopqW83/ZwPBQZkz5nJLkk4pI01HX7C2/92L3WbHo4w19jsN+VtjyyXXLJ5
eDw0MU0+czUH674pfHKJ5fwIJ6T0cWQIp5ZYtLeHYL7Mz/SQ6mt2o+cs6xBn155ilX7BclrGjq8E
CooHwXtgTfSjm0xNkgwfpcNGuaPxVE0Jdcjfkah9iutaifGl9FCAfbAky9r1yr0lt6rSNptjB61+
pdqhDg5xcQqNMNeciQXDb4A1qf5e5RRNtj88WwUEVdUzu6VUpHT4JMfZ8Ds0JE7vEqonRqRFIEvC
rxptP0HHMjT3bzVxwb4LAXTgcMR+uDSMebZh9OelM1ObRKnfUcB9gAL2K0yjG43wKjPmCxq/vJJ9
edZmlpZLBLHcUxwtL+1AlQ8HCUhQd6N8Ib+Ych7PfLB9B4edYgPD4BovDIVPMXJia4EdpucqcULS
hUQPHfbhzKHvAtSYlde/FaojLrvXVvSfU8xqcoSnOlCUUwXVbGDAgHsGmN7iCfws7B69H/9GcvKD
PaT6E+OizqYfxEbXZXWJ9Tjf3K6JmI0STtoZNBLmhxW2Fxma7JX63f13QevEMb1sFehBXCi2E3UN
YLxEaMWZonqwDHzs8Qyoh3x9jdLSBL+DwOuorOODmDD/NA+o6U2xmNHLw+qjfO9rV2DRZRl9ckJi
h2ijcn2E2cuH8X6k1jsCoW2KZoXunbWEwDKcWfogzM+T9J3G1EdlXLsL02tS2I8QvgttMdIfWxfa
Q35+jNTX6f3a2eFwvJv3lN1vIVjjMFa+RSQoJZmlgnP5F7fej2COxmkj7VaDXybEzIvSdatqXtE8
KIUVFBjkMn0O6ltzm8YGTsYmXPMBsEfmsT4bBWKzh3iUBbZRwFNcptxwfP06hZ7C83S+ajCBQTdz
EcolE7oCVhGOkwV3NLzSU1IoGacKeQNzm2N0kPfoNHG8AcG6vq97Lz60jkwXuGn3hrw1UTnYyoBu
fwuVcwvC3IQmq2su7Hj4aJWUAH17rA9Nne/tt6vbd5XQMh5ZUSewDEQaaVL0pcAhGfYBZ2Wsg2n9
Ycw/5VDxSu6MZM6SaNfCDsf5Hj1Gd2dbSV8F8xj8vccsR4OldXBfD5bGnGlcTN5OMI/ADkCDnzfp
AdXu2scXHnNbagVn6gE0y4iJAaDnXeo+WKyMNfU7YB2FT2hLmHhb7Vcpjz5XVf/xogjqS+pt2m3I
JYvXEgJfsuH6mK7cjfQaIEHcnQEOsj2lDznaCILlPNELnQgHvx1ttLDnoQ9Mf/Pfxe8lOBenEsyH
a+IdFu79t0w/pvJTADzLBI5fqDyf5OH6zd5FpxML0h6Afh2SDbNf7Qmi8o2i8mKMISwTSzk+ukih
Pizvqcqj0+zJ7s70ww1Rdv5NBM7zc/0jLJ1Rh8mFjzyZI2LqVgQHNR572HZElmDbb9YR+D94w1j9
XDK/1yuT2nsiX45kQAu532zxwSaJc2/B7i16E9+vANczbdQkWvg5eSxXqppUWYSBmVUDky9nwwmU
OCvHSof9zVaV6YVnWc+h4ocyKP2gWwJeAXtsC/ZBvMPGXGF1viDOW2D1XIaTXYofTw8oI8HrsnNl
jaTHjORG1q9H1s4hXRAGpdZ4Pvx3+Gt6kyynPFKM3eGb2ZQvJf8OqmDlZhfCr5Gx7ndAR4KcXI5N
tNJl+0SHlfkZvfUNrpGy5s+XrbvFNiPaf0ZVjbpK/+xpwdNrjJQKy4+DSB57tg84ac0rjbyxltZ1
CdwsfESOo9v5QBWWs+yvjw12kuVO2QoQx2vwxeYz+45j25OiJvnU118fW8PaT3m54klT38Oz5gW2
Jn8T1u6XUwoIrm1rusgewOKYk3SoMuuUca1sHHD92kAsbPFPkHJjXdzUbhxeEC1MTvmqTEvnUnT3
bxgqZsyK1YJpUSXEuPVCXUc5JjyyZSyRPqCLWQK2t5YUSXM1tmItGJE3rIT8Bq7HURlC06XmfyDe
4rKmVs5OJA9IA/vq97c9fNbFMHQH/aVs3z4f/1NKQ9XVVjHR5Lz/y6U7Whws95LSc/u2HQIX92gX
B2R0Y54gpYhGg6QOFlPy5E6RBZTGMdPXUHi7jc6UVNwoEdgeU0inQ8wHsEOjuPi1U5PwsUEellyL
Y3BJGYBOUGhA5D+U1Yf0/KYf1h4t21/FyNIUHo3LJ9oLgpSZ3PTj4ANGxR9VdoS3Mvi46sXM2zTv
fEa0W5qLf7MResVYZ0plOlhSesq+ID6G7urLTktqsHtboG4P/J9kV3Fk+Fg8SpsQ8DU0BLUGNHkt
zdxyLPsy+BaSuXeURQ5fONTyCbvs6Rk8+go9qogderKY7wsfc/T07NkRO/zgt4BWKZkyvaxCQTS9
2k5+dAcU3p45hKUres1FzlH+zF7gcBzjgAhR7APQotGZ6kx/dvUAGKmcLwoM47rJrbIQOEXyQC9A
Em2lE9B7U4ebyaXJTmfJuanzszLBIti2p1P8Pjc9QfuR24lGSAeZ7KvFDKXddLVsfrmDezw2sxaL
UhLZZ/38UjUZjf0Z2gnCfY/Bf8eFJm+cSaLb+9rdbBi5n7humEnK3u4kEOqVK8UGfYteUWwwYmQx
CWoxFqVkkc/wbb1KoAK8TX5wfe/ZKi1xV27VD4WtKPYdC3d0YUF2U/yPr9iPjRggWLw9RlLQpWFm
3vGVSGZ+XpO2ht+iYzuyZKWNWNLcYw2sXKxX3lmkYswbbyiKNaVYtukywU2+yXih1IVsuIFrWzti
+ZpzkHDfcXRgJrbiEOS305QWIhNO7DrCr8K4Xcmg7oEsPpA/ZWHi9VVS4zExY5icFJjAMp5twWNp
D0LvQt1KEkLS2hxEg9evBr1OLVvPmG8qQSAKbJazdpW6ddCsIY3nDkIswbJGAwGlKdxCyeKkdm/f
1ipNLWS46H79XUpjIjo4R2gcSZH/C4dDm2MoS4fCahSkAZIgRGRPtcjBoSFk7Hl8qFI4S+6G8NNG
Xuho5onrO2PGisqWzCOeMwdf4mPNy9gv1ravbwcEvSgJT3+IszzrmdkEJ8bmpNZk6WG2tF+lIcED
Ei/QHHnswWhMG3uuKc5b7o60/WAMUARg0IbR++x/xj32PALCve9CteqB45S8pd11QxseuB3WtlbP
VC29dQbI402qu4xGJH3+qnPAp9N839JG0rM0KybNzHky+PsqRJkK0FZ0WXAbux7UUDlnSm7/go5n
RJQtIboTmpFACMrqgssFGQ+F3oAr+QjZ6ZIgRUJBxsOA44VWXpU7VFClx64kDm42qzLo6H7hWSf8
BNpUGQgUEt1drJtaU+Bv2Qmsg12K9TO4OmNFuK+m4LTWce2CP28N29ORQnvZ7oCz66Aw+72MKXlI
VV8zc7g/W5yCs7L3mifQZ923/TVK7IbTVQgIi1U9OpG5ucAAOuJEBidv3WqgX/JveaLJm2T3kYm7
EI0/7vCSrp2wBPtcZSyGtIZ1OzWqXiaL47MGo7l6Kd/crhvPoYYhtw8dJKg1K+mo0OvDxjw/hZEq
4LPwBQj69yzNSZKeAIdN5fE9zicHe8USTRpWtHb6zQOdnnXoNLTPgrqBlCrDQFzX+VvQFYrDfHs6
a8VurRoVf+PH9ZjN1S6JllpNeS212zNIIffyFWKYSagNabLmzzFkTtENMnBdtCq3u+jwDU84FO20
9C6DsX6fLR6sJz0w/n9eM3n1MOfb24ezVTuhKxjDxnoffYQKuNEj0OnjWY9YHdbRifGxXLdlGhhi
qkYOUVR51wlCwuuv/CfjJHeD24RbwKssIh32OrLIKeK7Zv2TIw+zuOj3grfOfjPIaJa6pGdyG1H/
SsQxUaUysm4uX1NfviX/+Z0HQ2eHpOQ8VRAO8Pkr1Nk2pQP4Rj2+wT562G+QdQ6nqPRhQlSFUlbM
rMOIt0Co/+R0YevZAKkV8cRDINdG/H9imuO9Aq352EwPg1duJFRWtbLljx2wtiXPEO4doT6IBHXD
mncpik93ay2wc3nUHuuKQk4rBktmNnrqlSBIjkGVF5ZcbTKPMO9kIcJN4zx/ekJlQJ1OEoA5Skfs
lUSXIIio5I75SyP9noPc0ycdBub/E/9w0uG0AEHVC/k57hgDuFciqYzvamiDrOD9Kv8xdkVbXsSc
JplpoQGnMIZKjU/CCq6Lodr/7j3+YUp2oQOjlhsalH4TwsEO3nwu0DRbhsQxbIsK1Wm5Nho9nJe1
MUCK3lmgrkJSMETsIzeQyj0w88+iGBV41R89i3YtRNhNdxSoZGzMJTo0+nVN8nkcWR705cqZhhUU
+DsogssD0UeGMW6MAs6H1WePfE/f/ePenx9qFUdU/7t17ZzbVPfsdr3Amm4Cggojj6EkznmemTVB
4Hffemqr7GrDP/pIi3mbSRzGwTdl+YNF2OFA6jmZTYI2cudkM9OeV26mnvTPD9s8/0F5zS5KVJ2K
Cvv8ZFU18Ls0xxjS3FhQEyLr4ticP6gcM3IvT3eX1M1kcXtjuJmrvKvhn+dzx0/ln9kM80zq/55N
9D8V1+Jezio+1Fa7LvHVLpQavk5Y9Wsh9hbLpfU9iQNd50gtlb8MyycvBUcXm4OLyEXX3lbM+Y7E
HsqEmsarG+vaZ1QwjVmwU6LAiiVAjRyGG6dZtjsLZcWxaZxQ4RZO+2i2FHi8HzJpDPi7ycBxARkh
adk5YeantuYjaGc7TLzLiA3m2Z7WuTdkpgsF2jz5UdRwdkYERJDnjLIHD8rZ+kc6F22uhrupzbwX
yiqX9Evqx9gOQuzY2JoUBrlS6tlB76ah422vfvPXo4vVnR7WlUyygIX1s1ITIHI7TQl3iOpsmWsC
FJeiS9BFhJ+LAuY78rRsiUii3VBICZ9nTX2t/h8rH5Pcp7ZQ1WPFjiNHN7EgZGfTHftG+y5Z7BDn
uE7ERtpXhYZdqV7t1zmGPRHohUQ6V7dxZBDAQsyAJR5Ze3BnNMKNsNeDswu4094dIP94kPxmdgS7
MOmXxvvJ+/WFKST8zdoWVIylmO6CMD1cVTCXCubsX39RkNH1zNSGTMXo4B7sM+Y1p1gqgVHNk9rL
nAH4MFaauMO90qHz3zyqTz2IVPWUOFSqIMmWs8v9ugtMQ1v8oLvfbaH4T+SDNm+pHbzqESILS7fN
PrwYOVLFCy4OZQL3J1Hbb5ARdsfw1QRP2HoaLqtntUvVcZgC4/Si1gDnegcQsSOte6Lc3DbzmY8w
ctlifPRo1+Ncjl+WE1ak6WOvcmV+IPxvkv+vX+7UaJ8DUWpfJ74+79dd7HjK2gt5iri3tQr5mQ01
bKf558rjUhdlyO1VUD2DStGzyeywGNyZ8IwhK61MWewreFK7yX3wnkBHH58AUQU7/UNlEXtYy4Gr
J+VnZ5XwaVXAWj2DFOMZiFqe8Jz25F9Wy1YwQ1sxQzRZSNJoUABHRh8OA7L5XpWlTrCRGkZJNFkU
mai73PDUKDVK5rGAFsVEfHyH34KPBI2p4hICed7KRPkpec4gFwJu501Mcu9T8bL3kkXT8nmZJaNj
SrAljPFPSvw95ED7Wi4rOJFkr7+T+0xN8MhAs0KSIypn3gQcztk7hrHBA1KiDauOoHq/Tof2Aobs
jJA3UxOp0U9kVEkIARYmpZT4nAwmGrdYOpWWtOt+KQX+MecRSuOJ5cNFGZ0CmaCVSfJIDp3hOU4T
17MLY0Y0g8Np3fkit3SZsEt9mPzfHBGLRt63Fg1hpmcHfwlsq2VuzKwoYOJVZ6IwV8ZFv5/FEgi3
8TdjE7uzR9iZGBDyqw9gyk2zG5By5/YmgDQjmbGnVptWmxAIsLmz29zB7beBjCVghoyoDyZk5EzF
9FKmjDonlMYmJ/LX70+E2lkJ3xXTdPFs42RoAvJxuyIAFrZ+JFaui6+RfwJSiGnDZA2ao6mHBoYa
uYQTrTwQ8FAGrv/2b4DymlMg7XDCOD9O1ejxPBd4I1RpRMiaBZNFDX5yxZevhkQVoS+mqUNHad9o
Uc9LcDNZdEebe+9T51w8yD1lzpHe2/NCcKe3SOxEhthdHZb58fXiL1IZHvkpEyI82zqETIi2Nh0l
aOvRmU4VA5zo8BoLbagtWHmqUOytV+GjQ9SvSrHLWG3Wvd3sGdgoLOnrat+AtThxLfsZQ7EVNXOe
bqCPcMAsM/L/hTi3mTM7yYDiAgbjuueV5zPWXO2YgiiAxkC1pXWh6QMNp3AY+J8uI7R3vU/TWn8T
NjQ7jbzNBGXE5UrWdQ9UbfCAJNI8i800JRNVhiVLXZbmalZBeI8mObBpmFS+AgXVkZGAvm5GsPws
z8S2pT6ZoUB8qCBQAO32YlDhZaK+Z7uZX5frJrDeWiI5Pemt0OjFRLUKcTSbdizWzo44+a5WX1e1
fyf4Euqq7DEjWpH1jaEyQkqDT18JBv/2dIKaIK1bVjjX61dS1hdxTcC142FIU0th06ZnqMWFWIBe
+Z3D+EfHIbpsPAP0hF6nTmpMpy0E59L5mxm6zd9zZsnt/rKoLPWAOs+PF7qJAPwYakG5AVcj2hjA
G+7iox4ZXxz2yo75OFHDcRH5+eXKDaMqtqpgdw38P6a/30PldcnYmMV0SIr/2GGmRJcusfegr4ZJ
GWqXDV7k8jdHsFO1EtL+wAqYkt092zfBv0aBzdwFoZsDGTL1uvf6mbExPnnhCXWFSkZ9Q1bApl75
YbHQFGcfdigcqj53EiHzR/p2amwIPECmmwCYFrZuXvFyQBdiPpKOzljdIUmomFUskU3RouAU1vZM
ODqwtkMFvxXDX/twcwBal4UtIKgxQ25f+v5cG4WpF+IDdH1p6e/qUwSk7Wnz9S03h5bN6g0ccGRM
B7OpVZDQvIgUsLyAg25oqOeFv3YZBIb8L7vEOVfvGkYWscZEGpz9Zg940ZPowWCNK2088OyCR/bz
5SFAxgf+N6KeFVwxSA/C0ThjrR91+8w3IoI9vk+nf7Rw9sN6YOwjJp+K6CR1qmxcwY/63ZL6Obsl
esege67wh0R5Pn9/1pR93/IV2g1xNyrTFSm+CQPVp75l9pR1X5UjrUKXXCppFpzQ/wGjT+5orNSq
LfYvstWefDodDDoWkI/6Y9wjJJElsvB9ke5fqkZgtyucF8Zf72CPrf/4KxjSXkqMOFtQo2+O6jOK
gFv67iOlx6AKou+Xsd2gyxaoxSbGfemgNE43H5eUq/LdcHdqeMK3oG+0+G5Y+RmgAJ2RZ8TMvTl5
DnVk4INOZZgtI6j/OF7sgJzzYH7Vc9JxqNR39eyINcQm8dyd8IZnCK4MPVPD6igcYsF9UTHbg4vn
9Edy9JQD7M2kecvhV9WbPqeN7GnNdtLip1HO+IBxP4QpSkjnbSo6D/KoKU3c6Rr/QRmzKGn03uA6
n6o4Jwrk+QcGFKkTfOIrGlS3TpDEyyKkZvwkxvPxA4cGEsZEAtSsRR1DCyGUoliYqXb9EQ0yeFZR
8gvaU8NzcWNFZbYVZN4POd0P7U7Ez6jeC3zsLawgbnpHkvBAAb8n3V9NQx/aiuKHAsgajmFTJDWE
PwM00ydnkBUKB6d2glD8EAtfOHWEU31+KZwSqNLYwhjoppe8tEaulf89uQy6slXW473H62wvNytQ
+/Wm+HqN1l3LvQpKA2nPB4KFDggBpEIn3suP9SHYsHYzFaGOUeAQ06IHHLVDrHIF/tNRI404KBli
SSbuFiDrlUR6Zkt6qMrZUSuAfCCTlHVEHy27iQ7eBsJ3eovFiAg0ipJ3mujgLu/BzTFU8tdeMTkp
4Fg0knEuVHBOALqEJMa03vaH/UamO2oLr37HBzJsiwsMDuwUIgzmd2QUJ0wlIIB0sPULj6aL2Zxy
ApESSjlFQflUbkmR/dj4MEXghf6TWMl5pAlJ/JStA6P4t7x+nM8VSK4Y8PxrWHKvw03D7/98cE6w
qLtJmqBQ4uAfH88a30dvCp6fFFdcAvNqI8C3UiyXGO4mn+DsO0dFDlRLKZAaSlnM5RZDs7QWYSQe
qsu9BdU0GjTP9cFQmZRCHsnClpPMz04zxiGgEAtoFmZvSKPk8Kb+CyDzswXQc2upZuj1d+G4QAuy
EEEZ6hJO75/nen0HHRg0chzv3gWqJ2ztmzGuN97ROjkT6HrYn3XHbG+hpHKCLW2wdPoTUEYYPGEn
v9eE+3004HjfkjdzAkFZ8xwkTqXQUbaE8TNS4IdkG45oSSOvvTxw3ksYoiNTTansvcf9v51OMlv0
mM0aQUerhMYCX/KIBM9+4js+ELzpxc5WD0uuWkigKToqS6DK8lrUP3J5NZm9jJWhQR6dB7bO7586
ZVwH3a5sGEdUARcQkusX4maGCUUFbBm8jOpN+gyqwrQ2JOCW16pDsXsWcOETwXZ1b9G9WM+Di5d7
YBGcQSZCaFnSphaEqAeJj8q3evGoXJAWclXGCGnbpMTeFFXTW6d/YCI0h8XnTfH5GcnFGOB3/wls
PqBmO8SlxNU3bRGUwUUa7eF6gLXnjuPK1faxGQSW+R2GJWkh6ONR/m4IV5+2QOGPItxrXqIiseVn
MB0/9u9cGWS57U0Ug0KQPbc3a/f9rUTiOa/butu0vh371jX7s0uYYjOcz1iR0L2M6sEcYf6rHK10
ke+MCxwIRNJKQdEynBd+TRrkb7msNBiy0chUDCOvrd6Qt28x/ZwoSKOVMCvo4G2ORGyxNZMyIF6E
Hjn2izuNSDorOj+ASjaWrqRc0doFrlmIMKkUCgIoQPe5UIPPnQgTC0D8mYATlIWpHkJkdEfqzlWW
6sIuhaBeUY7esvy6Sjalf8dh8NPrn1CUZytIOwQugSW4cgdHv78QfTU5fPQz+uQcPHA03JN7gZG/
Xu9gGaNd4nPTYC6Pop94Ga+zQHiOZ19yVc0QeMMUTu+UyKhlENOJw8wqPSvruBfEa+TdFlu1BM6O
f49+MAnw4r1QdKv+z0Yc5n+c5pfiRP9xj8OORxbecoIAOSkWOTN0aQ3k0M5xf0no0IaY995BZfmv
IWD3TscaGr0MFLYIcXAPBlnI0lN56adkpTjtTZvKZsMmFh2G+1Lcvb5hFFdy9uOS3X7bsyy6NDmA
UA16viGAO55TaX4iUjSz2EaBz/9UOTzYpWye1092v5RlXHMcQduo/mKRSDg61D07lt/q99y2U4Qr
SPM0xlvNQq9W1wVrFsPCxZq988zvrGFrNPltbT5uqa6rNf8CeAXtb3KU5QLRGeGb7SSKrcaLx1I6
v8ERXZqnaiJMhR3nNY7b96t/84isPYLOvOviVyCPah8tvknNl7WMCWaggC7HpZH8nBnHyI1pY4gJ
cfT3tGPmE9UYzn9TXmqO48iyDiJtNJ96Q3zaKI8awnGvOlZgtp4UFxj7DY5cYFBsvJv1Hc3/7k46
sINPCyLpWqwAVW5bc7JJpwTipijZNuPsKtGmKRS6CXc4GT6P+jc/Um8XlopbFarIOPV0uPCsYft3
QapzMrkX0CqmO6mCJoCzbgYUTNqVrjLxqSHHGG5e+VxIOvwzHALvf3oeapaYu0LsQt9X5GA7YtDQ
oIRQaRZT76ATUCTmVJ1WrDas5aiClVm+h+uEzjRp1RnwmOhvLEpzjiiVNai62NRKSvJ2fFfstpWP
Ji64Fm2NfiET6iEwqp76NLskjJJoRbvYjwqvHeC1bNG+06jeonGKWogOBFE2PEHe21KGwtq2IDYN
+ogG3cHcqS6c6ZaDh+HsAadYvZgKapz6GG3vnZ/cGyH2pDbwqr46x9CkNTE/d6ZR4krh2n69a20w
aBKTPFbtAhmYs30Vf9ETkXEcjRHlzPmBtbKsNSqk9ID/z9dgQLZQ4g3h8/+maUfdxgfinrxpZZqF
vqpx+xfj3johdjUqdOQH43iZgG1AlrBUCra1I9wI5lXx3lSnFUMWJKcow5aZie4VmEtJ2nrjwNig
PjMjqKScA7uPVTFFIsRqdRNzAjbk3we1N6/H9lWi5LXJtuXdzZy0qfzaIKGQiujN7c3HS1/gxFVq
wEH2y4DHNT/Se2/D7h5yk0BFLBZYPr2TcaSZ6iFsaAmacRIvijBZMz5Taa4ByhPwVpa2PZ5UQL+T
Gx+vCerl1Kk7GHHm/+kyDUBsbb8rQX5IzOCDTyMITnaLIKA7Cr8eOmRvyBPPvu33UQ1DFpnsqwsW
B2QUm3COZHrsm46pK2kSoDr52hXmclCPNiwIwUxrlJkl4IB+SwJDPKi7RF7tBcxZTpa15DXhiNNa
I+D9CWNg8cRvmN3Et/b6W7EMbvfTuCO6mMy7fHNtGsRQKAX8wf8X8AD/mffZZvY3mtu1LPl1wLkg
8p1RDYxA4jOW7pRjgQFqsnrhUn4v2WK9ZbjGdb2+ZmdumlIX5527ioavhXSEyJSGA2oLA6bOpN7q
dcYQ2htfwljN6YRDdpBkgZ3BlTe3cwlBUf4Yg+8QubLSnHyhoKiPPpd+dirwU/ZVQMSJpeuaW+vE
QNjEGWbgxVtkxmIsrp11eig0Lj2VQgooz6C9c19rCVysg0U2b1C2t8y/0Sq3+ufPgyiTpt4siWSF
jCrl7xubfB71nYRhvcHYMLLse5d6UTtrTN5qMpH8nC0Y6+BU65AbmWS1duaCbWh39biExvFug30Z
jjIQ2NiinSMG5fFJpoDDBM++1ThL7sMiAS/rFKvrwVeiDVFCuq/cOHbAthEKjDFqSYYCLUdHuIat
aceHfE0TM3b5Hag50Jq016qBmDq8F9m3B3DuFJiHYrI6ixyORH5ZEaJj/w7SzDCarRfpSX6KDRpR
yQttJHhJfu/SSoB1OnwG7LAMW4Wc4HnroYQZAEJTVOf6zLKeaoIOYUQOenTEs95XONhlyYQm/TLb
88ob+AuvkFWD1lij1uKHa95hH1NvTnfmyN7557Od9AytfxRAOAmXveAFF85RESAgG7RcgI2Qj0CZ
kxXywYlN5lMkuXT8xZzaA5v/9Ooeop9Ld89xHLb0M/ZcA26V9deZ3eSFMSZ/2muRySUleysL07GU
74HLm2KFqUIr6tHcG6BENJHGHa0U8J27V65X55kQQNcp+TVYGfMoAutWd3KVVVH6+dYeHkCdHSu/
ins2cYcWrU65QrO2/Xj1XwwByFeyGKDR+uHcY186kUmjNnkmr2UvCQXF6tz7zFNSclo+8FEWLM3H
DwaHeXAy7DDBhbLWpGFbOmZX4Ds2C3gckT+yb7PFgcCab+SvFmn8gIgfIf32W+k23gAsAp6nC42y
8/xEsJ8QjqIOzPY6EP/CwWwwt0KMLIy9TbS0lxHh3AzMzNAm8+j2Kv5HmV6aLI+PgsNMh8Kdo84o
yjIZ5rIxX9ebdi5kqEYPWbcmZx9164Ui5z/KUacXPmPxEZJlxFm03oEmtrsGiYhLHmGhbcbsgws3
54eeiqOwJf5t1TkdeAeb7uTXlj588iRCLXcgLCLQJe4v0RMwjKravEkNeg5GYdvm1iZH5Zv5F6xs
adNe4w64hZfNFzMR1RCOSwrf5J6Tyrf5+ypaz3vVvYVPojH4Rfb8zBK9zZTJsLlmqWhwVn592vtk
v5E1lPhz8h4ppxhJtCDZgR0vjapEAKcv8aApy5RDdkAX8X+2gaFIsVxDGWr3Co/sQ4ZHdAybrkKj
vHtiPqJe5tmzMRKUXd1FtbmH+aiaZ7Ef+sBpq1WdrTJ762Jpg5tLA8SIGQEYlKLtZqzpdV+VgWBH
lXFIpEfUQ8bXlSHgKhKgaqGxtO8VdILVUPk/HCdFtJ1WAAxCUXhyCubDyP6Q6zzuBxo3J0nmQ15b
oT8pqPoqlwZ2kUtLxDJGc8sGw1tZ+1YMeP4w4eNdMO4Kh1A8sCaMMOl85UVYgu6peWblMJ9f8cyU
4m4aCVYkpHnjpCWEU5fXdkHwr3Z4GoZV+phBbwV3g7VnysABiVMYLIjpXTzjzX1uWnfGe2UJDN35
VfCR5NS5Y+nkgUYWqWHIvY7NNjm/BGj4TI7F+FeHkEgZWAvRmROCvd3jWNJ2TijZqeJR6WRuT+Pl
CuYVoUIX6dRQvzLilnA+EojtsLbohBTuLWwuWIOHW2fxViFDzqjTl+xtqVyh5Najf4z37w/7nt5K
86B6iT46w+GAE2WGZ7D1Bt+f6atGsNXgf/JfT79P+8agy5geETUOOb367GjSIk4ijVmvN5oP2POm
ZjlJBYRJcxdVaFsz3g6bv5PAt0+1JJWT/+s0fM2vNVLKn3fITW2HRov6TmrnrZYM7B8lE7WKeNRC
9qPP0hd2Bb/n6KM6ez71EN31Wz/cQuTlmsRU0aTDjv4UX1LR+CO/zXm7G8L6857m7yPNmN6xbDmt
2Iy0DEb+rUZB/ymwDKbGzTRw3kJQTd7tq8oxw6y+H3cJ5aMeu7tAjWHI8R6P1u2fJNUeCFiRpNib
s05yhk1Ml6nUAKDmWwzzCsDj1+GUfKEpy088lGAIdcyTNlf10AW2Qyr1nEKzoYLlH5s0bZKqUwMO
prng8u1BNTmEfiiL4HgHM8f+iTJ6Qf43uGybOyf5cdTNgJeogPP4+sH5NRVIcE5d8QqruOsuV7Ud
v3iYP2UWtJC6pVz8KXe3g/zn/E9cTa40Fgnxdq2g0KRUI+ubR+fTZcdJYMA0LxPQTV/qqD+Bzm5K
crVgB0VtoChpYQQXmBHmg4MeUKRqMQ+FMf+QZwlixgdNAagZr9jApRMbA5uwSFT7bqMYRX3a/y3L
AdxtiznCsvtPgPUA0iD0+w9sJ6YvYuvgWFaqGtMaGfYG4rGaa6H7bg+YkG8lGw94asKfthsn5yGR
epA+B6OgxYV5QRpevP/c7wYy+XTJiQmrWfQcXkh8/NuIuY7wscBr898qT7CI1OI6+WSybxWqNWm3
SN6wds89bp8CD706l3igjTzeEM8Gyl7WCLtUlCBTGkRR5x4WcP5c6dbzwocYDQz6mrMlBL14t93f
IRoCs/LzicRMNE9KEuc0sWgop0zy0c2bpuAocJ1FLmLdMByvNPoRKrLNQ2CSbQORYWDZMJZ4Dp+n
hkBbrRpizH6NZIP7qS4LKt+uJq2PeA1E/axp4wrrj1qlxNTIH3uB2+POGivqk6uVVQ45luW7zAfL
Fx0gFMf5z5uoy1eTvOQT+qAg/k0/aVadt+CGAEfhN4lBw1dEDKlT9l7/toZtQSLlSq5jZk4vzi4q
dOKIARAy8dflXMkdI0ZjXsDkZ/mwdmdsALtLIpQfzXEpiseuZ3ffu7QzwFLBZYktvFdCmRWNIokH
JA7cIXSCdOIN1HkPrYU/gHpGlJ0CiBPL34bpSCl2WRTCnGzqZ7pKk2JYB3ASQ8uUZ3UKdZ+y1e3s
rYom5Xzd0mjsLninwHG1rMLtrbZLg6LzzzCQTe8ov/Fj6is4kMO4Bsu4oAUjY8TnOQUV87hU7lhX
Hj3SNBZVDdw2IUVR+Jwo/IkrgN2QQcEDfbgQ1xKLgYORI4sOrq8/xDSEW+mOynxyq944/yabZcVT
wztqVr5f7AzkoGeeiGZ4KvZQn3VqMTcM/T79rcLC6eRoaD5uptd7iPwU3dit5lXzXVgCCdliyE79
/64u22HPoLg7INbrkDKp6oDqYVCSX6rAmT5W23/p964yKhIuK+aPjf1jqMWafNgjamPP5lg73uCu
4ylWTw8En0Eki5V/jawcZTpDNnSW7VjmJPHqyHmrKqJM5nG8QBg9ct57eID6SHG6naX9INwVVwqn
h8rV9/5y3sJr2jqTE/mzCakAPvOb668U9VPTJtQwNmsG/fdLcuBxpnuGVUx7WlMyHX3p1uESo9AS
T2DAt5Q4Q1ZtZgwlMpu8LQgMYa7cWE+NjaIhs/kDf+7iXf9tQVIm9dWBFSTIj7eKgfxvJh3SxL08
tbAt7o4vcbaJkAvl3eiGU2lwkXtGHyEfME6SQ6WZQTGWnniIIJxsI8E92SLRBfNMwxnPkHuB/efn
/dYxIo8ZYPVBASoKG8Cswn/bKQRoDNwKnoVjKCZ6foGJeoSyYPtbsoDUH8Xs1j6gaDo45rlT+Xle
PGK6p1G2c/ymJQOwFzIOwgmEsPzS+CuOL4qdZObC8Bgrllk6u0hpXpHmQub2TMqriey//8gg5yjS
RqyzA7kJMqiIBxJgqwHJHRUw6Ed6b/oRxy5SKAPPUYwfeLZy8Ud2R78Haqvty32qtJ1fy+ZN8aP4
NvO44tdE/g4BA3KKKwF18Sxl1TaVrFGxuz/3i01S2cDKSZJH2rkJURnMzcVRvEx8s84E32nc6fha
jj+Bxb7Sv4TjNIs1kkeywEKh+HhbOuK99iKuugK7HgSmG04ihvWhK3VBVdgCbzcrIktoAeQVosdQ
61OSNTfOjWaw7AO3SUUvkbPRMRDHaSTwVAdHTpedUkyDm7yj2qqaNCV4sn12SSCmfSsTANS6DBTL
cX6sCNS/w0qNiFI9lBKZdr3wuMF64CFsHgRpF+xPzzqK7GDnRLp6CnEuY+yHJtIlEG0utEQ6oPcg
UNlwSdS1lTl42igr6rkDb7KMMVYTb/XhJXKk+pfid53x8bXH4jOaeuS0WQM380n4hcsV/gE2PNSm
3dYkVML+FP0ybZDX7b4PbYvH1xzT0HXcM7lzAtpSEXS4TNjNj5zW29fuTXnJXQMfQz89smSns8Lk
7vRbYRS9nyrcWglAbrxrsv60zt/82QCKTJmI/Q1/rxUL9db6P9hlE0ev2zaQLKUm4NLEwHPSvYLG
IluozBB751K8PTZw0FN1PBTUC8x2SMvkGdbLtkI4KFP4lhZw8GmtzrG7GHd8UfweLiiJZM6/flLv
gEGbLi8juhFXEOctra3xSMDEBxkxFUn28B6VMXgsZDUwqLpLdxEiuYnqAdXmQi98wqDwbfKgMxuC
7UcwuBM93pai+f5ZzIITPUxJItxYqK4oVzl7wb4fHQB/U6lpnspxzNT0iqgeWT17e01O+tg/RNZB
TuhFi98omv0xE3Dberz7iVuNnXqI/vAoz306fZeZInr6JFvs3lSBqvgC1hjFTpKOtFJtT6Ya8EVT
0x/Wl39LUROpToHVzQmCrzW3ulNRKCRnqSuj8R5SwboCY0HvK34Zq8ig/BcoMJqsafJi/D3nFFAD
BmccEKbOA6pvE6cgc4l7Gzzq7lLacJ0NzGVIt3Wt1Y8T/uEod/WBXjmpf5r9hSQDORc4oFvBn8iT
RfEobpNPP/+lj7BLevyqx1O6BFK4HI28TKt3T2QdEn8Skqx4jipLgcnJfZOZrzRapvQ4Xs9HAKAy
/tsG7eqba+bLWE+q6O6sWxwSytJBoMgApugEf51ch6S2U/UKYBgLgJjbJPce+t1tUxb4htWrzt5M
jqyxVbI+loch4ooiksV2qJU4hCvGqRfeovtWJ/7t2tI3e5qZzxiVh2eyKUaDw/rLolAuBAFYRr6d
y2kuEUi2Y29Xohzq6J2OVMpWS2W5meM7/2renbA6WO3LeJHKFeDgYXI2o/+EubVZ2R5YnZKMKeCn
DoGb+MgOlNZN6gYDPwZCwQwThYmXZxLVwNgzYz1t4sKwYVRUcODxqYfDpBci9hmNIqwQV4TQRPM9
VPax1T/ja6ZvjF3G7sGPttKkWuYmovQRRwCzd6uJ1mRo5EPQkQeUF4Vbbk6Y6PcV8lHwUjLfSIy0
9ZPAAZJngpFldwj6ArDPUuYYp7TSUaTwrm5gZyBEu4vqFnJN+R53Cr4Y93fpVXib3HOyjjtVNU3m
Daj/gsGixwjVNei5u2iFhl0CPpRqejCgEq7v7PYI+X1GajNd3d2KDjdUrEHgrNJEKWWxAbVyY2NG
x8+tP9csXoMyYQzZseuvfxRkVl2EMN1iizAGhzGNts70t9fzfZC2DPucAi4TwCgC0Ww1+u/Llzvm
78vjkc3fhHoBlNkQtgXsY+mk28H62kRmqhBd3m7xuWv7h4ESbuopI9p20EK+P1zABYlP1fDrUM5I
uK5ppCpF8XwwLKo2rcBHIxUclSBjaOwIDIJPIudG7tSEfx9kSYWDWJG/9CXCq5KuOKTCD1aAYIDo
NI/UEOqDrqwYLzQHzWow7wCilGwpYgEtKJJ4VqEaeqfJ0AnplT6ZeTOq8xrv+J0oKQIRuE4eJ7Ts
QLUduy6adRf2pbDDPXZVdbL9ZIDYsTyJSWeHmurotCrrGb+K0rfuxNmmX0+NN8iE1B6pWLTnknNA
8ZOos5RHP368fM103sc09jaQa/Frle+AG80m7PHV+eNU7C//+Mdb1K1u3BDHAaQVmMMzyfZTuJOA
hdPc1uobbiqpO+p7chJCW17LVHO9K88e0USW0AjxcQMHhndTt+cdKJEz419TKXMConv19kfVDYtg
YJzCjPrhoFkwl8ppOMi133/I6SBVgFcrgclPA60f/0EpxVdrRDGNUzB29njsc+NaqmO+XhkPC71D
21v8Di3WlHbfB5XSXeba9XD1hK+CLmS6SWNGGH2NXB1azxpZ61IHd5JmyzIWwtrkiGemDRfUKw7u
X35MK9/ZgZowjZ6IrCJ2KVwJzmIF01KINv/1To6mftQJlmgMHQOHhhCxSshbm3pIhAp7Da2b05/s
+c/q9mSXZDgzY7t5hRhdn1gBfZgoAEzMbvr9QNNGR27tc2MYCxGNfO+ueZn2ArFzrkUY5xlj0v+U
N784aYUGCFrV5Bfo39hnnBPyhwJxGmxX1xVnfQOzqyADhQn8EQYCQzsyBIb3mnsbLRmhQuokaJkP
9UOlX33rqN5pNrVvIeK0fTll5VAOk0sEvZWyQNFgU4wRGvudnNok5aOg9EHcIS2H9ngCRLm8gUB9
rYB+KcMbIm7u27NQJJuPOgdISMz5Il0UaGew7Gv3GX1MYOtGrp/SywMTpgO5PNw9Jl8aPBAEoHbZ
nFPeG51PX/0lYlbJgYd1mgMDofsKZOJDN2j+LgfbDVCoOe1JcnSgCmp8OTRHDFddVfW/c0F9ATmu
yIuFca880yVWZk7okS33UfJ0A/bxvvys1wcdRzP2khaL+vidoB/PDwpQSSUxpILC1ns+fGjnkzk2
7X7Rk5+RMxNdrl1bO5sxhI8s204YRoEvkyjHt1aT5XIGg/rdUP7vZHUXOibn/DJ1ygzqEe0tRu60
89nJ7zI/1ExoHUdM8TaaNLA6ETePN/LsCqyKaQSw++ytCsshOlqyJpgMIDzX3tB7eFgcjsTIYy7Z
keTjF48N0dgx6Qv0JObQ6xtihZsCmaE4CdUTqL6cn0QU5KtFBlL07EGyRr0ammt8jUM6XRejtwdk
abzAqPSEsG8zT0TP1QdJ3q7Bhe9thNniMrgF3//4QQPJRDXlJlnhhk4BAldu2peOoeDv7N4iVoKg
modlZqjgT3ZteZEALxJ+W2kgQ5iz598l2JFzF50zBddf4r00Kt2kPa4uktobGZO9X5j7eqt7JBYa
GNjYWctZ0nVjf8cZPFlZYnL9Ea+PCu3VO7d9M6i+Q/SiGkD+man+Lk5a16EzDDRHQ4NcdrdAsoxz
NoT7fPwOVGLN7WTvSJdAGQUh4IeL7y1/S1A6ReyizFe75ci+ux0kN0+rjHdYun6R8cMzieDgw/Bo
MX2LgqFh6ZEXrBJOo7nj3OkAkrJ0FAwYeCZkG+2aRuJPkaMRnxSaTJGKJEkg3ic0Wl/djCdBTiGo
8DEaWDJu9gGFHCTmK9xLxBAb1L1jEYnhSxA92gkxJZ7b90tYMOItn+qTyrPrhp6IJ9jC6y53wL2E
EcN4afEFo5K4b5Pvuw5feJ9vKq8Hr71nzmOdy5qagYe0Uaio/nCXUY5CQX8osxQ2oVD2bCI2XnL9
qDllqpAGySMz4L3tTUnnTx/518XkqHJO+kVPFOzEJso5pgpzt7nfEUa/RviSBHYgfyZYphg61kHp
bzfG55sgXLqR2M+aQMCPpLYm/tNLUIyu4D5C7OzjRLZ75OzKzf/wDIMVEAIsVgMBoXhSu1hvtifp
ize0ijm9nDsyIu1F8/bcyjVOvn92BgdX3DxsYqeCh6LdyDiiEMIB+L0bzqtd0P7BnQ2KVfY6ZRP5
tBzw630RNk/hJuPbnOMuzxNS8yIGZxzUAN8WkfmkkQ8Hm9hzzZqxpDLsCGPCk6LkE9T96Qmb7gIB
4kglyEC+p2QE3sWYQQFA1ZXR/U0HBrM86alaZ5Vsp8a/Bj1KrYkVwQfwN4HqyjXiZ0cxIDK/zq0x
pMRkbLEFO/yKCCDqtPsFAwlBGaxSs48odzg41dyxkSPuUBkUjg643NS2eIoFhu77JFhEc2qhSPks
uL/1aHxjPBeGY6VOvqu5n8h+vHwH/SxCJVrXnRd20F/JnhA6r7qPxSwKmenbsikqzgQ3KmvSiu3C
sSTqNlwUJTcIttEO5akNlA6OyhV95uUEQ5o/DneWbRpJj0qzSMzEY7uoHgkbFk4t6B95atqEAmSj
cS5HmE82VuBxpVzPK0r2qmpjUYaZZjGotha0/Qv76Of0RVqfJPMrEZmQHZ/eB3mk5vyWBiF+klLs
ZNIXal5dFX3D6hHQAvT9PttYLe8Oq6gYDPNj6ifAp+82SzE+Tli/HmpVXz/RR8DLtatIT7kkhWMQ
+Cl2cFvsEDOxZVs9Y+yHD0AXWT6RoIXYACPAfMkN8w0JmVarKq6q4xTwEpMfiqBWX7gUg3k25dA2
KWf69tNBOjKXnnPXOilq3oz/9yYuDmdGQSd2mqxqRh4RzutmFG0bJtq+5AzXDWhX4oyynXcCK204
n+Naas2LcUQ1IgtNW9Ob4+/u+XdEE7EJ9EdmYDQgLsWBnsX/e7Ug/y2FTxpE6idPjPCAfGQgtiTA
IPITtwKQdWWm77tBVeLC0j2DJe1BEdwkm2DmyDM5utVULrR0mGOgt5FMBn+Y9lh6V55LENUv5/I/
FJTgvX15VxmU7m88Fqy+pOcaA1HNsosOjAJk1pmDvJsiwBkYTOYFp7zcR4l6KV7WL0KGZQ25l1fH
/1iDTtcOfh0FA1j8IvVVtoicUEHDpBK2szK4QkgiWXZFmPQYer6ciUR1Anpp1hprj/r7IIfwaYse
bDcUWgd28bShHLSrh9c1N9E8s7n9uOhNXzQv9Hhy5sJLs7eYhrDDtC9j/pfA2b+dXkadSVcUB3Su
7q2QwDXEd/FZXD1h1o9AAJoO0m5GTE7LzB7cz8cjiuF66qAyCU47F/gv6wH2BCfyiVwdwWRtvy50
qf5GNpnslsTaOgnfcZ4oQh0JuQubTuw5At8dOn9+lZqWKVlzlSjkCW07yf4YA6+XWwOsUDkZIghm
9l+cvLNIfMy6td2uK8LawNinSDVvrjNLIwj+bgFkVbKeCtkb0cxQDBjY8SvTGdUDPhf4QfS2aMfb
TuJr/89QYrnaUC+WRVjrLwpaNGLBrRmtvq0p69a/V80DG9W0Sm2ehOg5l40ycM45QPv70mYz2cpk
38nvK4dKr4IhX2BlN/Ovcu124Iqev9K6CQppRIVfypOFGt5VLY+spJM1BvbQKHOjBTYF66426URn
K6nrkLVV1F1c3UA97U/zRDxc+tBJU8YQRoppq/IU+EAxAvGNJARCRD81zoLBaYBRRSLOLiIBdPPu
xzmCfCiSeZ/yxVlQlDJAri28s6R5GFKDMlPxh1jL1KFEaCtC/rWFZD+BYYVFI513wH9Qq9IiXsbC
R/MZtFaSvGyx5DTj7Sz4fBP7DOo+4ZdrtR6RzsTbqvUxrUetvGnyWNjuAS00Bh3jAhjxBxJZE9M6
ymR4TyAhFSUmF81eAkOksAr5IkHUU5pO8+OOUv+Uh/8tJBs4FglEInhn/EieNT4ggqLz9zuJzQq3
JV7Wd4eT6s1JlxTmSok8XYQQ5d0D/kr57cqLUAdw09PwxAE7bVsg8DO+fquWKAQMDKJaOI7dBiHp
e2lFuu8jN8rvBVhAwChj4DvA+ktZz6niwEIY7ClQsVic6z4HyKct8BjMGNk8dK3zNFxY8y4DEJOM
JdESnDw+S3v7o0OijOwXgclPWkIsgAaEl0TnYQ9r+mmiWasuzGqv6bwXFvfe84D3QHN4RLXOjzJ4
A31c9rvmF+8ntpmYzVDxRAz1qOe7y09wmGYqP1vS8ZRPynKpej3tb1ieidhWHhK8IdcHGvuSbxG6
1mTwdRy+YRcnJs9/HmYhuiFfPARFBGnlFpEKwGWe8rQy6sDATg51dXyBWjPYuMR2B/kGbI3PQm4h
q9xMtYK4ThVuPD4mWoLNBE2l828ckNmtr6WKk3D6L1c3qMPVU2ztuiZkjvWyQ4O0w7BAjEqf6drn
W1G84kxRZ0o7wbLIF827DqhBz4YK2zDoTGAw3Rx6542kluToTHDMP4g5iF/yKouNM0Ej1ZgumOOA
2mShu/c7COQyg+hAu+kOmMHiMxTWN7FONHPFiMhh8Z2IVGJgBxIgDEX7v7vTha+qQdu5tKg87sdp
mL3X0XEwpgIPA96UcuQLdOYehTI2v9hyH+lERQXs/n7XtV+IH/LwL3aLAzriNHlIpGGjy25+aglf
iDEUPXWMwOf+IzGBsJQsKs0hSFJgRTdx8RpQ7PWPF7a/Y2OJ1uiiycmW/rKdybkw/Go2QRyng5vL
CIYN8TWauw61K+bbSH5S8uNey7ypOejKwZoCFVhFJg4GqMLm629e7mRLc/XQ8gPoVZi+SRAVdrSH
5E9t//Gv2Y+xGCdhk2me05arBeP/0DH0SrXIlDK1nww2424vtG2lthBV3yh4QUUYizo9OkAb4cSR
7Sd0lLGvFTYIVAC4FM/Ikl3dRldPY9H5hOzoYhSZIWsr6jM9h54C5FPOTJnEE106y+X8L+47D353
yBhzE8FsX0yQl/dx7aSD2HPCupdN9G4vfNWITZ57f5ViAC7lL/G5PZjkWtiZJm9vSEXXUxMpdPax
oYk7O0VPpWtll/z8Ld3d0a8n6bem4fqyzjcpxs5wicBbQAi8/+tXHokZkjtTH/XGIrapv63HLw20
ZLk3zrsPEEDoAxxZ+QPYCDD2Kt5ymS6563Y/u/8IuZo9BbdTktyqjXiK31fD7jB2LfbTk5w8VixX
m5a64nNbV3ekYDPXp+ik7Mus/xNsvto3X9dYCmW3TPwnisxQ0nnYhzjiZRXgnD4x1x485yAEQt5I
vhkr8oMnVadQ/BQrAYcxZQLw/7yxWgNr5GqbX6AGEbs9XKRHh3UoDtEhbkPEXvzU62dsE70CoMIi
RUCy553SlLu8ZwZvedqcgHI5evmfVac7lLYfCfjiFtR+V8gL/ypdlbOSuFL9UADKXSXOQPYKVU0p
gXdm2jbAOmXQLUXMMqPuthNjRcJU8JqE7P1citDRkDAmGeLV4HgC0fVcv2kMqrhkdPZ38FNTF+XB
waQVrCzapKO9uoQBTmJ/Gkp4Pnx1xaap6kGVBrXrHBuv3vEo0HlNRwFoCsTms9FxmNXVKJunizVR
nxo1yVBo4TnjBkYZOpLdYQqugOlUK/R5jfxpy7tVLBApnWNRvjMt4ZfD1gX3WjQjNw6YfvFnnvlQ
N1wnLj6jl3WM5gDsXLTMvcCo8bwOe+z8slKB2tiMPwLXs1RbGJwJIlMqbmWyrrOH9HTJWAGTdwMC
o3XghLxzMk3ZLnUbZEc3X1xYM7+plPL0ppIYsemUjL649BAC6JMglrPH/l14H807bv1boygpQ+Mg
nX7eNTeY1fdGbWW+Bc+jBpDLOnYMJulKVlj49vBS52NvIUfs2TFBg/OEmcklFPI7Zw9Kcu4AkdjA
817UqlGYSLKZVnkmfjXMgCSiI/xGa9UgOzGjW2H5o/CpDCwzGJamRrA7fEzMEj2o54j7bvOvNgmT
O2aYeQZ9BKrRaDy88xkTR3tXT+h08G+cLj3vOBwX4ri+7XOLXUuJKYrnap1AihHAJdoMdN2NQXBI
zO0vsz4+bsl+aWBb3ryWZGQ98+ErY/FJuUK4FAvjIniUaKPiR2ERdQrZg0nanciFK1/KLL9pZWvN
WPz7z6LHX+v0qZB8VF9PoQOLP81aU0dXCwxGbUL2wSXMMKaIQlM/MlXDBJNdfP4ULTR4fEKioevM
7osdQSJ6WmvxrxPad5AzxZgkLcaxUSWiZgP0nV1eNRQkKbaeam0wk0u4kB2Hi/YeXyonBcq3eb/b
gKz/WY24EZ3c7as90dbNMugAHGyv+sKTu7jSBGtdJ7RQiR5oGbqRgIOUS64LlQ4pWdCa/oh6rGHi
YJDzCJQHhmFOrSaogO3n1WtoDyxIahKI9YK/PZnjQk1FG0veBrN+IynC4DlDwTkgZ7gbudJqEZNK
Q/ChLPsYSYEtCNfpJXcWspelLh0IXNwcrWITc74Jp1E5ANRRSU2mCKe7JtDwmeM6FlSLMXoyj3L6
Z/npH7m+TC3L0Shm7D2PSf6TAXWNdPnAwp63dLOXdhrLOSZ2I3thvsvIFY+5fFY088jiA3bNem5m
wSvg3iuw4nOp9Gg5XLyA0xI1uMnqkJYwA/un5DSTvnu2rZLXL0TpAFgw2fj5TBWWRmQJU0js9PTX
PG8ZUGwlroOfs667RaqqqB06IE1rzmzCvcwTcAfYqOa5mwCiY2tVu9hz8pk5sEQrBSJrifr7a52b
j1SayDaDcNef+ArFkGjcE8Mm1yftojbnxpsXuSmR7wq2fFN0jaMGXBGPcg+U2EGRjja56Ax3jKrj
fYdA+X3KjADnM3X5Qx8zbLrsOLKOtNFoBh8eJhw3dbLIri7e5jOuB4HxwpOtPzEZyV7NGSGDKB+w
/t8KvENJFs9Wf+I3nJ6dAGEgR6v2rpEUmtvts13HzSiiAZslBh1fuj1NDpsme+rU/yv0pwHd2If7
3n50RaFKkTVv58AggJ/1H9jjWQqrPrD0N4zdDHocHHQeknjXZBtl9RTtEQ1TlZinzNyAKJtMWuUc
0xrLcTGMgmCLNiR8DVghqGMjvHUaI4nJtPXuDW/R4Q8pVwUK95Qwh8r1jRCeEmE/Cr83n8YPBVI8
SRVQi212Io2M8rQRSvhSBR6eOvJ10rqsTcPNiMGiBWcb1empd8FfKhHNnEE9CU88wH9OiO2Ll/IL
AmX2Z4WtksQeDndU3xvSRf0lmu1BfGA7AJmmeX44tHSv5GrBzK9E/i1Qu8JMEVw8L92TuJqM8W8Q
vR1OK/iUJdyJA/sDcdUHX6OjazgOeQDGaNKMYwvQaLIIG3z6RJVEMxO1VIV7FtOIaPSmjMc8ptmv
Z/ETTHfjQhjjaHZr0KQ0LH4Yk0eIKcKc8hNEyEvNybEiO7pZK6HK07jcfSeTg2ma4q3D6Zl+R4kN
nIKcOdTtNK+lFfrY97BhYQADemuvsXgLvH4UMzRBgUW7COUMEEv8c+0+Anj4ab0hJB4gJgUE+96C
Dyok2gfWwDLsLNu008SrGxrT3Xcii0RGiBqUfpP2djdDF/k/fYIbF/Y7gomSmq++Uhidtkkkssmb
NcUxB76+pTtI4Vs+YWl9yQs7OM9Q16O/SPDFFdlyM1tiR/L7nj0yNXeaW34rlKqGnMHkCW9vtKDY
Qtx80zyJgaVhY79SucnrrRR0quHhN1mMUYIxQfpuFNlDSDdLeyoqJNh8lkKfBHGu8KbA49Z3zxmH
NBhhJMy2vOfYkWQHMPhmj15LrUE7iLWKnpB00BUZ2xt8newdO8xj3+RSAaKMxRALbSbh4hNC4Tl5
yA+mkkYT1AEY8WoHXX7bqoWhWG8RdfnZAW9zifkVJODjTbuy+TAf+gk8xF4OOKtQjn29eWysNIUM
m66XwaLLNVWka7N81FIfe00CoA5c+JZaSl5qnxO3PvNU1R4VI598lRTA6ug05E+Ntn/9RDWip+8c
CnnDNlSow/E4Hdbsg6LyPfqgcaCYpXkFWmvkhQr3q3VxGWgMRRZh5SsDhKkVaQHGBihCsVK+tZE5
wB8ZIMzy1xFN2ML4IZ5OV3IoJ5MwqHK4acjEAshtK4qBmnDcFubLvWL+TVk6l0t5z9EU4CzhPV82
9qoyif6IUF4TwL2RQPmwFc+1xMEiqTIKf672SDolvV/Djb7sIK35dbV53cZUTyxkyrb/JZBkt9PR
2VzvxYdM8oFwy2UlMa2J1BqaruQp6Zsg9os8bq2oTzwfAyQXSe60962S0zOSKf5DsVd4kdPMP6WO
Wf3LmIAA5vDdlP+ConKuq8xK92MnWKpg5g3jwIoN3ZTZD0UHBrP8NgSZP434NtzrbCF2DG3OE9WH
Hq5M1A4wOS+G1WdeXZxgxEih0uO4J3XtILfkD0H6ZDpMNs1PqoOkUKn2jcF/WnFMJqDBB1PP4Iwl
G7kKwAfQ+N0HDowG4xH4RUfUcxds4k3/HvmUWUCIO4MBaeNxFLn8urcRg4fuwggb+CfIdyk1k/dM
YYxYxD9tw6s7TCSZCXwRDIzZAuEJpCXwIDWWwohg3JNOhH7tN+6LbbaCx476GltVhGoLodbGyNIv
s6MSAMpn9z706ui4rjyk9oh//OGStxkndkqiZE+1/Vw9Sd4obIHb1ohYwxtBwVXasdAe4D4rwDWg
W8P4v7aXicYnneFE/4lgHZdeDfDzYLwVxYVEce/s5C6yz0VTGGoazPxRCgsWoQlbx9XHRl0p0OoU
jmhlt7haTp8vrcWMMbrNkcFSRTDBw9H3831Bn0r27bKRek4XJ9yRNM/791nNCIYHmv5lTDzD0tCU
e+oaoQQ46h4QWG2npoQ7gUh1oRKa7nXIL0CVZSfyfYPRL5cVBtQyKBjzRicMRmZ1KaRC0Yw3vc6/
cI5kCtRZOXb372aaA11I1Odp2he29TUCwDSHAMw+tqvWRA3KRXY0nHOZhMvom+kNjMl+0tLgJbCk
wgWnAxZgMXPC/k+3/L8y696u2UCcD/h2869WYd5GVPO9cwGnnBNjOB+1E2nAVasd4qKRP0Ow1Tyj
F5V+ocLWhbSksX2JyIvTHlWn0ysoFnzrrQ4eJsK7ANk1TdXwwVHKla0C9WDfZlGL5bP8uq6ejMiy
Fyzo6R1tl80nqkojLLB+A56i3P74k1ln632n+tAM6suSjSa7gjmpZUO1rOb1Ec5UKD7xEZibK+cQ
nzu/z2rcNZ9UaSUuvpHZ002rH1dPeIhZ37d6UQUqjCHhcTih+WLJTZN3x/ZOH1Z37EpaB+hA2GXI
CQI5pqq69M+Mirfwtvnq6FwNspE+jhaygiLKj65IVEsiLHL+rjd/QDmzuXqFIlMxwGSDV5KZIxEK
nW8sSinwycfMJz/kripOO6vKwwbyi876HKZdEZEDzPQHe1UkSS0JQhZGDAprZgF0YCtgojuv6rv8
8eSaVDHcKl5QrFoGU2PmdeL/hG3IU2UjKmli9KWjK2awb1kQ1W1yLEVUIQNE3Y5DLIyw3292H7di
KCyYkOh4jZkuUACFV5Wxp/0Ck5U6GDBmWZZnuHCPcojiiGgXl5KO/W1iEPMzl2bmv2qv8cmZmv4Y
kvBRCnqBDZxKPQxDcl9N48EJvxNLFrc5PFd0Vq9OAFLitI/rpo3ql/Vn1UN66Qg1U8k33izsddx9
Qvg1A+QSFuZ2J0OJ/TdOzwwJvRs389Kf7ZmzjdXAhNW9dv5e0Tb6SfQE2n+7prPyiEkWbkMZg1IJ
y8shDwfDRzdejgWGSUQ9/nTZPOb9s8htK0su3Qsb5s83+wyoMzHTvo29/F/oQJ2SbK4aHPPXSmuo
gXN7yhmImA+VtoVC1WuKGSGIbQubE1xVgqJkuqhWv8xmp+FIcykPH2o5ttM/UVD27y7SY9RO2o90
IGb5HkkeT8l4d8y3aJkl3Ffwq8vQgAPabVqS9+B4gOuZ/PcEwbAoHmDYelwceR8GdFJj3A9V1xdZ
/V5gRjFjQhXrRT57BSCZwSaFVuJIDAqc3YhtGlYOh1I4dpdngjyRVCgQn0zN/A8L3jOSXvq1CjV3
bbq5Q6HGOtwbe1P7eB27t1FOhj2bYitJpTxPXm6/o2COvtCawpjqtpAt37ofZrHdVmnSQ3j/Frf/
0OVWBqs4y6KiFcdj4e36OpFuZETqOVh2FmGJ9CveEZgdeq7huRBEEheiDyL5efOaTCT31uhvivcY
yLT5Tq4HsrNwxo8tuNxAPqxm0qFt3Za9Qb4/ecd9bNzSIlfU25m1nDRAodxP0K3J4CqRZ60M5Mgi
ryHkwgq0gtnMsXxBwLH99MkhSfL2M4AcbcGXcp4ioWRJhmdxeXigSLlsOt/jQsiWUQzXbIry/YsZ
BDXmIQOBTJA4bdbNZVnFHNeJlTef3dPRprPux3DgbpB8PPGK6x+8a2WRlCMAPpbmMlNPvegkop5V
A/0gOgIRyUji0AZ2XSrWWVumMed3gY3DM4KUavtJ7psUUPVNFL5btSRjmY/zD4LBZK4UfYkDdWh7
rYkxsMove47uZph+0xu0xL/LgIPb2LuKN723XRFdzdpsvwt6XFIyx/zQkNDPdYG2BMWCZZFM4Sn+
WiIwuQPlP9YP6qOrLkL8y1d1PS4vs1qtpDNPF0xpeMJdSnyv8FB4fOe7bn/ZLxHQr46iT5SCAVpH
eVvs1c6S8twtdNpkLhxWM9bp0jHVzz9ORnFy/EMUl4WC2mHXbaTnkAXgF8O0cEwRYbzlnqlQbbg5
J8pocC/xCxau2Tka//n+EUYg2F0kw1u75NYpYP4eWdnmPBMIQ+A/e77c7kZZNwzat3B61DhAtZ8c
0m/4TcaeB4NUfkd5pHiPvAPyabwwMX8rkTAmX7q9GQkOwxsSkR8W3BhDBSjpbl/3Hw6xysmPTIQh
HX8CA6wppKQtObVzmr14dqb66nSARItn9aJ3qZ14mzxGJmp/HeEm4l8qHJVhuB4vFIOsZd68tuEu
K20a5viUm2fm3pu6WtuE0lvVkrLY/P+GF8r3NPepQVn4wpmrzjJM1HwsZJUVsDI9hEEGDehEMNzi
91VLDgRLRF/ZPRgXb+vnXILy26Cvf9o0SJ9EAJnsujD5L/ebEKqVKWWR74MQBIgqPTRuDS2/SmOH
hdA6f+Y+IgfWUzIBubcab+tPDVIIQe2/ej6P+zeIdRkn6rAQka3njUTKn//yg4fG5+ofwadzliYW
Ch64ON0iknAr4tlcu9aBkYe4xpEcu2k4BjpmvYMaQzoLfHA5Sj60XHYtpjFrEzlRFbhbMGezFM0g
Y2ohZRTrrG5ZdmtKV7MPQQSSYlw4jfonF/nJULfOr9lFCGqI+gbx0Sxic2t+QFfkPe2Ey9Wnrp8g
ykQEm/YNhqhJMU3YxED3yqiozPC2Ad0q4Sy+pmrC337WUIK3kJF2x6BHOOHcgcqBasOztsfqt3wp
DBU3bwy+8lsGPh36uhiQ9KhlCxEQpvFwW3KBN0m9K8TYrLxE+PfVI5bkwYGRojSiV7IP+aIhMR+A
Qxg8AqygRW5/cCwS7ZogNTe0HH6ma0yJnKuhkouvC+FmfJ4xZA9bm0hRzKSFqbnk9gbHdDeaT1eH
tQ8BLwJsJLwbyS7/490OLp58WXj7psKA3flZYLmLy/SwG1KOWcwMsG/B0SYA81qlhoAXOXDnIQhp
b4+d1CHjqtM2SLjHpdcGrw2BH5WovRPyKWEkGmsG2o5ZIxMQCD/W0g/+IYsIfpOsBtwT5spHbdIF
n5wAejJWTyrcY6yrIV3x8iRcmHjKAH9RbbOfBrw9QNVvG2PK8lfgvQlieqHH5Lf+tR6KLcGOdr6Z
LH0JaU4EP1VDoLY8TWT/jiWSDoMVlWBDnyLtAVAyYtxb/hBeW7Ae76EmyLb+aZ6fBz4mWq95HPzj
3AKcsBdTY0WP65NKbHO11NeKYvdIyobUetVp7BkK5B2HqvpgsHPqMdj62V3g3dm8LH7GS3HFkLxJ
rEYj6gQDxuWZShJb4enMNCE+8LM4+b5+TJ7mb5nurw8Pg/kfS/3eCdb9zwhsllhIrQ4YR4IOW2PV
p0oQgurKpkJIWJZ3s6jZgUBZqPkVFJRL/1BH1oiYHeZxFYrFQt+avMRu4PuYK368oF3QfdrZR4iI
PeSEHtOE0u8tAjGlr/JqOnZLnPhimMwMUnCpgkQkin8jJ229ChvLzFR+OYrKM8C53YjMp2GNILfw
V0KZiD7N881M8vMVhR6gfR7AYOpEpWh4mar+huMl3cIhF3TdBcruqcfH1jJReMWPa1DYyMl0Xw1Y
0xDDXyMzpWdltgXfHXAJCjRi+SlelWvoIAaD84lZ7z8fhVy6/3AYJVGRqLbNDXGQj8SA3zQdYhxq
HvrKnP6M9iPlHFNsg2WJNRwposWuQWi2pD3JkV7EmC1Yp3cDOedkinm7tmxs3z1cYzf+wZEBvoc6
hXQt1QnMnjce+Cq6UUMeJKia/TqH6dlvfmM/Il4Ai6FotS4ur6o8Hxs7fj18zFmGb1z7mzqNCy+D
tnvxlcQPmgaO4Kp4xChBif0adkcKEJq3CjYwj9a1yI84x5qpKuTt+rXO7o0TWdcmggHeSt1GTp5W
zb5hDVl/vkVoTrVPuWIctmIw/KxqOznmKnmasoHwE9D+NONeiVkp+gPbTk9Kum2OH2kjJJlihLF7
1OvOeLjDu9AlBaUhjkTZKqH+vxSUdVCewtBzwqccbC1ESrLojaO4jlmyOZvkuLAFvB507b7JbfN+
rK7l+jlR8mpDptewp+rySoMy63AvJhTiDyaZIa2hMW9fwDoyLwdLT2e1wAqyU/jWUGmGV3vS2WZZ
uldtstmvqvJ7xnbfXmYkCFtSJknyyFiGJ5xcZwZlwTYaPlGMnlf+Kvc6QQy9e433WsDcbKsHc4Yu
VcY9z4q55rhqPqJMZZ2EeUG+vmmhp57UgcS452hrEvXJgNN2ROLMI96jLVJWHAAJpg5CmOx7K0To
UT1OZRBtG86m8wgRs0a7jkiYAxhYpIlpSEfQOCi+N4lawqtVVUSOjohvMmzUyupEjWNvEC4v7Dit
Eaq3hQwHjV3nf9pVdqMr0pfdLZQK0Kc3NNJdv+7Cz0g71JF1yMKv14BTIvbVPZnqz3XLVvukz1wm
FCxQNEZj/VesP86PRjrLikUOc1pcePeGlvrlUBpsK2RCDHnjdHkPgYjR38/i1lUVBACXJN7AAOgI
5r+I/RMXHOvFiva8yFPvNraAbzENbQmzH0W1i7Ahrpqk7C/ko+8RIzoAhHhm9GPZE7Y6uZ66j8tT
r3+gAJECcLnsgh4wCA/XHc2xxSWXcVWyN2YPYAC42Pr7jB+ax8TDsk14baSMBr7qp8oUWc1/q3Va
y1k+c4HSDbq2iAl9YG2E8Lmcdrmt3eiS3dW8OdDSFrxUOMDsgd2VcR6b1frGyAxi1Yb+ErOj4pBr
pckVPBKM20dDtC66Ssq2a5AWSwNzIoHxF0/RWfiwYZ0ekz75Q5jAVzu3DLIhN1b4hWw1yOzaBUqV
KGtVAPMl+dBd9fuw+p17hqG7M6VyOk3sksEvdCm0dNwRG2uTelcYFYP4a3kSNvmrYpFycKGtVkej
zXod8eAifZNyUshbFdYwWB8mYxFHAweA/zcZEZf2p6NbsOiqVMYNc5mqK5Uhztq7DO/9+S8LJ1L9
r9fS7aiJD4G8MwsYoACc63khuxpduWLvIZRBcaRUk2UDE54NZ7bzoHDbGs5T+JMXeVlOGntRJcc/
8fAoGCfMTeDHLjWoEvJO8hETP7CX+2v1JwYIs1GMcEolMMYS7ai0m4lkjI9QpTD1QoNXBqsISwpe
r1sZInHIUy4SjHIYFTeKBX9ONwYhNBtBnw9jB2awlqsdZZf852Q/kCG06+ujQdGrL0vNzhhBZX4I
SDUGSiUOGxjVqFWH7VPpOUXrCYxq+4dgjxe5qTYaGbCbXvnZcXP8sYs1py+8vFNrXwB7AhvU5Kge
HGapTdoTHT+CBYAyCmQ98WhuPkcSRqAavgqcpTf6pxo6Xxuir5iaMIzcIVhnKin7RSUac3/enlPD
l2tFTYEbrR1C1Y/4LfnKxAajXWnzWa8nWk4WTxzmfEzQk5EZAj+xV+iE43pu5KmXoQ5cxudN7hjD
oYZo43McQitX655Wh7shcWcX7da5L4yLkZQUCfD7gy/h9VP38cto7FVg8pTUL5cbOKkjuHMa/A6L
he7DDZbQ2QxxYj+uP0lwqCWLF2Htlj6PK4irgq1ak8lcmaPG+7hjIWxT9aEZ31jFx8KYHYFeOQFr
3tOQ7UmNUW/KZRTlaS1LEGD0EnY5ToyMvE5YD6c8SQhwt9CGv8aWPLmwWRcpqYyEVIRCGG2utkMI
pLkSA7udZ3+YWVFLdohBPmhn1XvbAnDYQ3yd9Jddn9jxqbMIRa0oXv5KEcJPhtiL0LgAQQ2cnLH3
XQfozUcIQzxLmABfAdRkBaPw/3kQR3jsrVhduNq97uZf4TtpJJkiUvsgzkv66s0R0I/HsNxDULnm
Tn9az09NK5tuuuCK2NcU2DAv+MU77OLFO21M+RpYwKC0nc41zUYRbhlKV0ANCoIB+38Xs+EL1zRt
gWYUGrvjK8B80UIGJ3Wl07zlBbh13ChXm0k5fl5cAn7QEZJfopP/8XXFOrOj3FdU8d0goCdIQU4g
ZLwRAMiTThJeursfNz3S5IUCQDPdLOePHNO/wIqAiEBSv6ajAnDe0XEZYU/Mss+05mgTmZ4UiwXB
0M5s6Vhxmd+1Pt/d/9UT/PNpwP+tDJznHMdTJxMU3IS3TuM8kBY/KtEgTbROi0t8C/4Uk6tYCQpL
mZx4mY5b+2xAMvDsC2GkXSQT9tViIyNWH6ouGpUR77VUq6pFbmNbkMk/+piAlEAnI6rxMxMDA+AI
FC9c5ySsOk5G6Sr5fngxSAwJqD38Jx4S9wv+CheHXmFhzSCUXQ4tEDkWfPf9/i9nUrUfeb8Dk9Cw
6nEoJJPQY04s3HE5RsCAt1eIwiSSGEJnKPc82S7wsZdRNpW9NH7I7HTLFAy/3uYaA4hSpGjbyWr6
Wd167tq5CvwfJh/2BXKFz1O/hH2CKSZ6Xo3euyBLxM31p8f3z+PPIBu1aTEv/Y37zZz8Hx3PwakE
sZtJLHtWNLov4GE5RUMJUNjUnTTBYr611epW8KJH4QMxE0iBwYGCV3srvrUF7L6nLUbFAR0/3Y6a
r44txT+KyUAFLzWNhlnN6Hj+0VMj7HYBzdPLTExXXx0+RyJv9qczVPSZv9cNJ0dGwcdzpuc/hz0o
NN/NL+qlJ0nsBhHZuTLU33gfX97IgpqSYxRP1izWnuMPtfdseWMmNEu2I3zrRfRdaab5po1o4o/r
7F0Tjn7DFEwxTtWV8srTFpYif9VsCrL+C0zYOGYqeRjiA9mwsQIWSQ9rbOY5zo8QxXHTcvN4/e9l
lyQVy1KZNYkY02Sv8VQPrzhfCnK0bgIA+97qvSZ2GNrm6CkmKiKTFlx7eL5oCplC7ztV2DQ4bKc9
zI+E0yQYxwD4LC29k91VVH+GtK5GhtY1+xKZaxJARtdOamSjUBAua+BY9z30UcsqVwccSN7Q1MUE
BSmLzQ/L3Bz2QRHJ91lhuuSWof/iVEe7P8eU9oq7d3T7ItOmLnV6a1LqTcLQoHQv9SuREkZ1lWok
/g+xwnDWPIYlMF40UuVAt1v4CkzsGHKO7fJAhKwuRC6CiZt0k+V1zAsT/QtpAhqmXYZi+g5Phsho
wIBghpnQR1MvXcxN0aWJs0RthpHH5CmqidSDxSD0+n/hBSt+xPV6dk003G/gBS4AJADo0mScKO2w
GWzt6T0YmJAiphbIOxdr+KjyCnxEKsmDu871ZiNRUinox0/o2Z7eAEC9D65CivlVD8Kg4LeaPqZo
iD1EA5pOquNTYXEnCQ0krW6/uiR8k3d8rQnp3zreQG45RGgWh6FB2XTFbZQZvPXn6ts+O9eDPrbm
T30l436CGUCXX1lGDnMdnFwmNT7GstG1J8WlX24g4NpNcSSHqoO7ZeLcVzOegiA2nlizyB78lOOv
mnjIWBGAsSOPpp+rZkBi5Mb1C3kYNQmGw6ClaRz31sYCz46CgmThzvWPpApfhPnSWhtfUe1q9vRn
rY3O/ZpegeWQaXzD5cGFXiKEijgryhOLSfo0ANzYx+Gqg4s+PO8FgukYbSlDPHe3d4mDWqgpxEgW
t3xBaMecti4ENNf+m/1Q7HD7D6ZCvMQbPEhZjbk1/ejxvp2elH11Ry3DKqwAWWilCQl5644LPsmA
dSyy09w/pCLb0UDr+yXLQe7kf/C2phrqWcWNsyP4pVVP9JaCBXIS42GIwi93xlpBgruUQYhQMkps
rPrCVL0csWsXmeTgzTe8Vjxn6i8k9K3SoWBube1frVHGG7zoqUbooK+kPyKzlzj3JNbXua/7a+VW
OxpU62/sWw0VixBrTLsmsqmCUB9HKVar9K1wZdtDh9AsJNAhFAyLieArz7XaFsifKYl/cQJ84rL6
isVEk1USF0e7j91l/xgmCIuxejReK2tJDitFpC4NoljxAca5I1QMy3aceJvWYlt+0r0mcy44jzQU
63MG37GlF6u01LJ2zi0zmnXi88fJ9TJd7PDTUxIZFwvS3B24hEwsXFrd956XcBatY7I2g52RN5Dd
a46WIEqEKqKqVJ2aAb1zhOo818ccULoc307EK+0JzqSag6LWzpfeP337qzKec0Ae7vWb+sUk2YCE
pSr3YiM9b+H5mqrH0UK9ep0+CLurigiptkisa+l7rLGkF+NNO5r0QblsEyXndl7IqfOnYdWAm9X7
V+xDumqcKmG4+3Grt7p8rFzbwpq/Bh6YD15pbvKZVbAfH1ATZh+dr2NMui+M1Fguov+zkAJrrtPf
EJIpLQemGos6ebYU7V/g4iTe7Znk7a06Kqd613db0qpVzH4V6zjMbYk16Qj3k28ZCSoQabWncdRj
urLzhIoJPoPlajTqagMQzH8v0ZTKoxcve2AiIQSdOr75UehnPj1YtDB+OyuhEIwf6mOfArd0+auz
vVZVr2stjCeL/iWPbFvaBx9HyLHMwzGyHi2RYbVq3Bb9BqaKWw2qoFJrTSH989BqynOaAbjbsWvv
MYPL3TwjjWOB3bVfgS3YTlM02ENXAgpkfw0njhNvExn4trub/RMtr+K8Ip2X4eXgcNNn5FVK9pXj
u/+6ItJc8UeHsGCc8kAePc0xGkoWMbJM6PVqXAxE8nhBp82rFZTPDOd9e6AnObxKRgPoY0NL01hB
/+MOKZ6IOmhH9Xm0rx4qvTRFny6E21Ah2L/hZi87vUB0fbIHY1NB9zkB78m2Y2ZN8OWSddMD2pHP
iFrAtpBKNY+gxPEPmkulhVBH0BDscZFcq/Jh4730ZWwVHYpcuXiRROiLLn9MIPpWWAtIicwohhlt
qz7b6QeApK1ZKXmtcFCcyjJGI+7AWKrq+joMbWfUzw6IP0Qokn+v4B4XR82AELT3K740hJVmlURu
seEtUyWYLdCcCA7gtlxyIiJhAxlAIVnpmReRLv4fjgH2RgaGlT0hLxhLNL9PIQYPgGoDe5FA8UJI
eN+0vdxJ9KxXyYeXXWlr2hxqqx/X4LCSilBPtmhDW9Eytnz9rNABo4xh6X7QJRSSSyR6157S5IaV
6h2Gymp3T8h1hAPRGz6Br8P4l5ahDdeKOhiBpzI/Cgfd5yKHg9X3tCVMgEuSzClkiJj0PNYzPR5L
IOT8A5ydJgE276euhsEKou0DHKmuHO/KF3j17R9qK8gkODZbKiBHBzBym/nTbb27tqbU7oHEr/u4
sc8Q0nFuwVvQAA9WYZxf9oWYOhgPBojbcbrG66RrFEVyAMY3/WVeACXo7nGdpgeV00nxRnjrk6Ob
7PRvz7WGzEwV7FOY8uTJYKu9hOttmQK/iROmC8PRz1BEt1oeqBdipqxZXB3gEUB+/TpadnfGtytj
4dVwX4n2c5zhnaF6Bl2bySh/gWFQV9ZPYbay6KeMlHkWf8xKn6V6lRGH/9vBxokGVvMigrC1hxlg
8sm7u6bbvSKZvGQk2OHjjp1AtdCzOe6+WL+ROUmJJVnDJghMyI9boD1gT+HRaRZC/aFr3VCcGemb
+2u7EO4BMFCwSi8w2XJx+liuOgSLzbg8bU3e+FOpORqu9xEPPZFknF2e071iML/i8am3dLjG82GG
stEzvZiuohKFpy2BUcyC18h/bMNzMWQZpAtjNUf4M1vWp6h6kkioJkyDTwirC199VVA265mOs33p
bTj0CPGeo+2vHk27DIm/MfIrF27fr1oFD0kaMjglxoT2go8CtTLphU2hOKC/kMm+2ct05km4dLr4
uRMM5ZolhYc7p05/0bwOitvrE2lf1ABNaRTbospj1nco4gOz9MBBBTFbZlcMkyoWxyaKiRlXNhLT
iYexD2dkoos7aAyGM4GxN1CCCrsMRvBdhIZvFtXxWSAxlxeRSPv94OUwaljzKes8JtKCP5RwFD2S
NqZtNGU6fZmZlh+AIzeS6B3vrbiJqVJELnijdboA8VE8T6ELsnBv8Njssxb3vQoCfXVEhn5aG7Cn
EGOeXVxQB+Cers79joW+2R1lFCwD6mtNZs+OWKAzL42/4iySxLI2gqqFCFHn5Ic9z6ouIlvKazi5
v6mq7E27a7BlvG7R37d5+iUw0NDYCdxjXkuU721Sjykz4SgOiDVMB46jHjJA4lPHmeeEvsJ5YF+b
LxkjynWyExt9i1q61bhB99GVBrWrr5bs/OzP/G9DUOCRIfrAePw2W3dmvYBoAv4EslHduUTmU/JU
wyh0f4WBSYjMeqo7/7aa99gHo40hB1KFBr04ESMItwF7pjJvP+sCrU32WymSe18CSw1zNtNQJyIE
XqWDzJXxkfJGOsTKlsCsCA0T/0BS8FYy6b+GeWWARxTA4+2UgNFXdM9cFHwM9gnhnvXzcDhz7sKG
3oe7Zh9WnupBBBvTCNrHxp73HKw9N/P9SFsQfFXtN6jtnRhAj+DJien0ba9xpyn2BjOihTXQ/oCD
wx+eOcsbHVzVtG1H+X+ab5h1PFPQblU9F/FZSeppdYsb5QL0jyVm+//wF8uMxQaVNCTWsa0EO0Qx
a9tZekKnDaFUgm0w7G4A9n3ISgljZ3eIO1GEYGr4VkJ/jU7OAGfdjSEY+sHvSvZPUn3bXsXpBqLA
um+BT4rodk/AFAwHeCCW65wp80V+c2+IFAGRJaV44G/JR80nKThwnmrLszJUAeThEkZ3j+PMV840
8n6X6a1mT5+gjX1imFtvRCrOtkJjZ1gzbcSMDYCnSNp3lG5ddpk2h7p/rxZvYAHVtcrtCnTYb/yy
2PJozdjCG5Xk89REUZga5Z2o4OkRsR5IcHx3KTBRXlVD+cgMN7sx33qcCEilBvssj69PxH6yqMR7
im/oyUIkwaZPJkjpQEguHBoSrLmQOs08emR5JjdbrGHUn26i36CCZXYDg7C6F+l62iC+tNC/EEpu
DijywK/5LF/w2i9EJjVGjShotqofdkPB4/nNyM84VP/2JRO6lnvBX8RWrJAtE2CP0wKil6JP9DLa
jlb57ceOPCmptVGvLakw2HfHh2cmWnoQVz/eaXd1UZN54KDef4CcTeZUBMNzRlu9amtw3xmewA+L
9C1k17XtR16yc4n/Z5KLdMVFHbg2T0a0as8jQ2WWbCylSypdyA37Dnzmp5Kz4fFvpxQKNjOdKrWz
9GVKU6Ou45A35n7PUUN+FnhbduwyUNsG7kOQNNg8+ssG3sEZUsJgEGd2DYTPpicwtwciT6dW0AZR
y9pNd/LKR/BrKLxxd4dQQwS7CMKNa/xOJXVW+gXwFPIfQrg2c5R1CCaJP162BI3R2IwVygmT7icV
VbixHlMpkIv/wII69p6BY8J1i7Nhld2SiLSFutgv7bkO2QtPkgJv837PNpdIdTt96Av/t+GFQsH1
do1xP/oBhU8ruIKRc9hMWDPhCQy/ginRXQAoNc8obOsyyVncaIy7Qs/cdXxV3n2ptbjvtEsmQ6Nm
Gpvpu/vHMr1p1xAvrx44ex86ntSblSg/2pqJ44xC1PWq6O57XNF/sDYTNdGqozOo4VEzoBI+lVjo
+tpEl0OR/3lXsNyRrpYTwO3YKOWMZQmB+p5OtibvxouozY59svnMbOivvZ66OtYyrn2EekcAyBPl
tUVQciNreNNX48SoesgUGKJjqd8Q/srW+bXQlW0Ca2epwZLpm0z2dYYrye0geqkrJNfPe6YCp/57
dspeTUf4uYYXhEIt3Qgrefru1kf/lsdiHfwglQ4gd7hrPsjLF3ULcXUKpvgpzCYQNcGZS0AzceE0
FvWea6ttV1rYit21Cj0FnK8JVUujE7a9hc13/oN+G2F0y9IlxChKlB3gimvvt3x4GYUXx2uwSPOO
pgScAyLXovyvaTVGFai/kWJW804K3SiW3DAL0pb2/yeA+au4yDDrEHo9HG+awDsJm0FpSUOTRtgN
Dp10jikFuHOS8GMmowEQrqmuadT3xUasrPxbuKCrM6JGpVvhZhzsA3I22Pv08thudc5bkpbL67r3
Rvins3lf71es5wgR1YJZSXLi26WXnjYWd2rWTSUqZsrNPLMFNhR5WoACPTUoVcpCR8MMXUjeHfA0
an3nPFdUHHAdIRJEFG+ft7ihdODtDEYFaoS+g9urypJ3ZsCaPm70Y6WhDmT7eKYvlZjUJwhTq2ek
V4KCpAAVsCy3m4cKbZ6VvjeUfdjFZEnxvu7xQQD0/6L5ueA1SF97u81pw4liwQZCiAm0sA+YhJtB
wXuAP80+E/i/a2TOHjiMjdyXC0+WBmv3GU9qOFFkct8gyiC+NjfmWl/M9ydKpKpGAvCn8wOPVchp
xuicMhWj/A5imOalsdlmBqOUOA+BocVm0drEB47MrOGmhSTFlioqaELWOcecrxbI6gsX+unmH7rq
OdIBAiZcj9f7lvv54Y/TtNdq1kylAKiMVbyqOEDA0/FrjUDYm1egJO/1Oz0wIMYepPICgMPbh5S9
Ygu+vZquKVt7rc0t27WT/uEMDT085rs6DmQ8V7Nrzb45PFfWZvhkokXwuMd4RrZMQzaVto3xbPId
vHZzFcdYMCuNAnYE2sVeVouKDh8vdE6Bf2mfShJ3J2tebVjgjZ0jO/fp4rp1NUcxgMd5TGnOq5zz
dwjA08G+TieR01V47OQgv4BMP7aWMGEahoz1kb+HlVU23X5rCeLqSRZHfAF6SGKn/93MerPsk5kL
2lIXu907bMscxcKEQAgt34Sk40hqtoHp0I6PYgb9Hh8dTVvLaBmSQ8yQlJ1wyxZlq9jyRaKLovl4
Vg5cs9OUZGEiSBI+TRr54oVsCK56YZU8mxgWnfa7i5qlwerOoxx5o+RmyOXn2xfjTRInwxiu1VaF
M+/fQQmhchHsluo8vgn+oP6Uiw+S5fNa+xt+drBsWRZ1nKEn+r2GCYD+toUCPZSTMwwnrcjISX3A
ol6vtdopeAWI+yrb+gqZX0fQsp6CSdDsIC1NB/QxZyKlOYJDax6G/YXvEnd1J3y3tTcFnpMKg4z4
DqL/Zk6VxryWRDEnar58AqToUAlkaVAhfWGSteKWc3bQd8S94bXoEYBTt5uV6Fz2P1ClFyLwNUgt
IDRJ+j6UB0RnDDZ5dFJhYyLGhRNk1ztKhombOzzpu+Zkx5HsjNNkAYgNCN9JCKvNlDvzRt5/cEsc
TVbq6lvfEYCCtUPTtqAFNxgbH2VxbmSQLwkrGKO5hofpTRn/PMEF8UOdWYsH5gFVvvapsJap/Xi7
4dj0cRk5GsUjyPsuBYaFByi9L8S+PAImtRlv+WAWmM/4leN9WCWutkpg88UWfsKK9HyTR8LFZAol
F+BmDPsHuL39OIAa1K3/1rtX1sf9vYjazVjwEuNoNdIu2HBtkRqeFfMUC5/+iO4ql87LhxBlxVcH
MDuLdtHD1agZ7MYaW1vvEfPsXYhDueesGt+TBFnV+d6iMD8LVa3nI2RHwApMSkvxPoQEG99rr2u+
TJTLhV6F90Yx8L7V0tTZ4VhvRVpx/zgxCpGaE5dkTzoe3lMYl+Rp0EJEADrQkbN3ECyb4Bp5xlb6
cLnF3so5f9r6jjbu7ZJH4OsUsomxDnZZWKByjkChb85gs7MXGUrBsBtQFJS2MetSulc3a87hLiFJ
SdNW0vZqC07rp8/r/2o5PO0Pl4/ClVh4JCqwJwQYP988a5xYhsaaF6+yfYS/iWG6Kh0dUSY0TCq8
20FjGl2i0djMTFaJW7R4aEDxU6IAoCDi7hw8EdYmZ/jCgmPTB/voVaVUt5tOpMiVJGCxqLTq6/3w
X1IOHT8I6SpbD8FgqrGl2GeFIcvKgz4EC7INfK9jVffctPi+vWVsiDli5YC6hFOA1arnhbagXHf1
Q3b5oblRdnCYuzwc5nuQoj3cJ9okiIgLR3RzlTRbxxXwqe4tjqQB4tN6kiIyJcl0A3OlRGv/9Yqz
nYn7UakLxldr/pxSvR0nGx6YdBidzYpy9+hENinwxrN9Wqi5OBJeZ9dY0oiCUDsUFUaNQil29LNN
y8LG8BeAWL4uZELf1m2F0LyDGXiVMFXClyge38KyfmB9y6nlSCjmkz2qN+unXjhyU0hKFQQH7pRq
A49LBVLiXaE0kRDqcW4ZIDiwPvPSnf7AT+k8j39bSr8m5EfvkTNwc1aeb1hI23aCEoVia8yQ7BnT
fENAjEUfcYv79NRyoWgSoMimTwVWThMdtr6toUbpWBpO8sOlkvMx4JPW/Pmt9r6TMtb+qn8NlEN3
LyICrYVa6HpI7jYwoXik6zTos7DKNJiBdnQwJP5vVAAwCFBkypxxcJbqsi9VuKl/Ti8mlS589MJU
OLXaqMI6KvYAl3j8/7yuM4PVhHxaTyxDgO4VSQgn5CeKi2657NgLy2HNPSRlqkaAy76p4EmZxbR4
1LQHLel6OP8ZI6/x2bSh4g4WsN4uH6F2TKj034uudPpBzGzMuYJZjbCjhhVmI3xhWeItNKBzPgiX
L4yNt1g+kCFScBctA6lQT18Scqi5hqY0/6uA4+2gJoYt0KfLzknd7as6JNrBEYTjHpfapfkvGCBa
sviHFY4IcKqKfHW0gJFlLHaHreEWLgQkGThtkXjklhtDr/C2nW650fBNzCXRmelk6pAP2qxD3dJI
4H777c3IXvjhHolxMcdHUdhVtpC7f0aaVQEHYP+rQ56o01BzzWHUnb9uqI3+5/F6wemXtYk//bS7
emiOSPKrBiMphchTMcsqFcOcOk7ZZXF3yO5wpP6ht+NdT89C+93d3cFJn2doisrZG44MEHPNfun1
+6NDpYQlAsXApwHvwdeWY/nXkTPQO2VqzLeDVN4YXHblCah4m9F3KV41g727NNNfHzU4LukgEjbu
fPPER4T3MeX78iAEn3Yur8lVJL/7A9v2eFbHPJ+X7EYjAt7fci6vWHeewdaR3ItWVcbUr8p4596a
eRSlQ8dRHYluFRwHkPc9AkdGfYZ4Feao6DpF7TsJ2/tZtSzFIxr/jXitDBZdw1WEOLfDP1WlktsW
kvyTiwBK9KkJ0hNyp1TgB2jwZs94YNQ4nXAmckmgNtt9LKuN7ciTbxXN1G72UFUO2TQsR2ZnCiTw
vggUAwQ7rnezQxV24K7vjRpL7ItFaR5Vx1+FS4f+KtDs7zcTN0dhCmDMxBaXhL+1qG2HbwrYX+ZJ
Z3XTKLXP/zTo4ypu1ed0vGVhtYslm8B6hmPX2esXdDFaCuhjrI3uBzBdtaYvn94LCI0IZiQVd6S0
LIv/7uqnbT7xIQ3b1m2w9il99dY8ikDJJmfqVCEL8lncq14SIzVC3C+WebY8S+IC0vlA1F1JrO5l
lrxlru7alBTklUCBlq9l9B5QkPrfKhfBFIRfVsJgcQTTLGBMxhWlt40MWUBtadL+blrP86WFp0Mu
S68Fqn81yYO/9NEIJ64AFq+zSUnZgNhuTAzTXxY6WNnBVe6hODAEs3bGvn77C9tS8gG/J3WRVffA
0TCQ62WnHKOmVLlG32u2Su/eSUajr3f1J0E46t3TLDZrHVPbppGvRRe9ooTwEoYhPXS6yFxvKfSE
ogRnNdh23C0mMzN45ziYpaUMucKzTFg/zcJDOS6aXeCnwFo4D/mvnOdRDpO/UfPSioEDcLtBo8il
cHTDR2qwJQEM1Xi2PTpoypVVESxDpbWdgaiy660LSfhDtnFwKZ99xTxPo9WOL6zlj69cMYzANNWE
2I0v0LjfSq+bdlVVZVJ9dRj79VgusRsGHqHhcknxe/GO9U6s+ax82nlFH82wtIax+ND7mgY5oicr
8PhRnlfzkOkFsxQQMo2Sj2nmykPdt/r+IGXHKBE+gBjSaO5OuRBgAmZXyZfC+s2h/ZOKGnnuADUc
t+F7TW0j/+L2w00chM1YfPW5XkonTKS2NpH1YOMjhDa/5YjjFKGy4X9D+y5SzZnUww5rPVBMSSfE
mE+i9scfQ1Is4GwFrF70nK5vpAdjXUQ8xmmab4uAzycnzPIPXJrLTMH3yy9OOXxXxJeNo6VeyGGJ
0c5C+FawYDt23/nRhHUa+wrzMjVGNtjY7REPbFo2+oY5xY1tSfzESJEGV/zJvd/c4ClSfhm7kzEn
j2f+zitPbBV3KZO87LCcrgqHsIEqC0e4rU4vtpUUWsv4bshHNUylRzgib45Pk6gcHvG0tHD/SwEv
e1v/95Tcm9Uhlno68SeOjftME4+povJytI8Lc6O2wOEku5OKEvrAVBsctGtgyiGqbco5asKnLq5w
OUPzEjPhvVLuIC9PuKosnEJFnMuAa14zpXvJzV3Zfv3DTSpO5GeW9mb0gqv7CeyjXo9wCzX/yEZN
UtuzEzA8N0GNEBVgd6uli6bX/JrkgCd2TLbvehcqPa8jYiHypEf9buG1MsIB0YIh0TK9DmaCrPiF
NquzioOOTNXtYY8+1q9c7Mp4HUSgHv4Yx5ci+YAk5mR26Jr/dUue/CzlILQxjFcy1V66SfVtgn3f
LvUXCbUUEAJZ7AjKJeyRcAK5YBP1f0osls/B9XcBTidFj9VP865g7J/LVnX2wrS36rhtncq6vBAV
u0Yw9evhhghpZk0RLde2xKrQBPpg2/8i/yEK3hJiYG4PaIhz43GDwOJmFDtiwSVhlQnVIs/Cf8hx
zPS1yFc1lu+vJMWC993HbhPpWO8p1ARxDsi6UG26rQMVdfgbDEG3rqt+LeLFS0cVaILIrcRtxXuk
QQ6ayW3oiH1DFa8v1SWbIBun6jl1uei/1687W0iSMPSpCMBPOqO91eOwenZKqtPqhmPewowEQfup
mX+tBPBFZaUtwvTsPOJ4El5j+MphxDCMNciNJotMddHmdlhY9DycOopz2TU/9qoMd7gSUkOLmpvn
RP1PVsBYClkfJGknvVOTVPO8fvj4yBmlF7TOpCga2g30cDbNgXUTlcsu9T/o941p9zcvv+HCh/lm
7KsNW66e7VMDmpZSz8RHgQzYnPS1qCqsGYeTd53UlDNY/4ZxVaHjiM2wJhI0mkifP2i3DmZvwblZ
5ndkkEiMA5nhQKOfkUETvZnI6rkwC+x0Yy3nQxcDhWO81bZCgwrnA3od9KJw/dou/bGvTDNJyWl9
7pENYMUWbwn6SzaW2qLpNHtwANmOjJrLqdUs1Hd9RbZxSlIfS0503Vp3o1hvK5sbql4INd0Yd/uT
xVlzTIibLTFg0ijz+ZQTQVv6UCW97x+uvxs0Z7ENYsaFf8JRqgYLBtvNeP57cgldRKxEyPXxt1Dd
HSgxoTFcKw4lSkkeDjDfy6P7Ea0polmd1Xnoqf/Nykiw7NzM6CLqnjuM7kK3Tz4m+dskqVmA609h
WviGLmTv0R5ZEWK1+AtSfEl7N2rG4KSpJfChBovHWjWNig2p5OJuCeFpT4FeHB7YKfjMj/4cx6Cl
FHQy2A9lM6I/zgegFSqOSI/Dw/cN4mufZH0xbB6EAML/B7fPyX3A0npHwLCQ+XaOTtcK+rAMcVbC
XvGytBad47q5Rqr1nMAM88/k7KmRTiWHbqiifoK9RUxYEBLd9wrdFAWRxATa+7JlsEQ5pyVKhqGc
kjE40JG3woZe/e16fbP10WCtBzW3G4a3EvpP9fmyTFgwUu6CBy8H6vP6rqRjsk3G9OVneOav7H1f
1ej1HTFG64X5LSwq58ttD5RONH5vhhRkF09CeIUDOsBvsy/oKUeRLUCFAoaJeer3YAaz+MjR54aT
eA1WEcTG4zCMeIvTkIvYv23mzSfc3T8BtyVN+hGtE8gPBh6Dm2Dl2FWGBx9x0JriTXspVIGhMcGb
fURk5QYwwhozzSdQQUNnlAjfVk25kuQt/DqwFXXKnh+ZGOBpWof44TmpdyEKnwIzV9QjJcKutVLq
B1Vxh6eY7rfrdAVD6AAq8UCCOw7Oxg5AZtiEa9cqD3iLB+jjXfo8l1FuhqTJIDymXv9ine/E7E6d
VIrNUdPDuKMBBJJZreUOkH1gdAH8wgcASmvdNKdU/zdvh17zg2q/FxVylwLe4KgmBH92RJDClmsM
MXvnLMuFoS6FTst03a9iwnUhf0N43gbO6ocZMogr/3ce15NXNARxbS0Flu+CpYrmmAnWslAIz2t2
/bnZK09Wc3XQDxnMKGoxwBeM9lmtKYDYBgOKo1D3xIXJOfsmnGXa4zQWIw9mVskTqE51ghkej1Ft
ZupJzCC3O6kOh2rMzRmgYNMRaLtPdb9y25Qndfqr4M9ofEe2TuM4Bem74f05uJkJXOmia0fD/4G+
4tHFj8CdppotrAeEVVaaihsZo31erm9nQfovQgtowWg6io9idtck0MPSAcD/yri6nJum0Gcc2Go5
0OXDRB1i7oTMRu8AWyt11XY1kQUWZrF2sokmWyUHvjcSY5tXjEhPattnIx+pKbV182SEk4uNtcTZ
TwvmlhcIGBe/zhLeTmJQdp56qLU3/urhLIhr/NUgOLeJDaL/W5VrqNoAkik0DcfQzRK+qNyvKwJP
TzUt4XiSIG9F9TycLmDIa3Rz9G4WdhN8BoHqf9XM46bUZ3sx9Or1mnNcD2n8tOBD9O7dcb9+6VjZ
ZuFdiEnlEmJkZOnBPRJakaXEkMPp1lmGlWNq9wcgxXoysK+Xm9lIJ5rM1Q2OmeoftfPaUBuNHC9s
WLai4iE/6Z+0GrcuVxIfDd6EHkushUoYTFqlmgsUiOgEwJj8iwa0Ngkvk8LW/j6drqEQibyOzwGc
EykcSdYoHE5f2Ex5OJ+UtNot/hWc+ZVy1PcV2M0GyIMKEV4KsZjV22DQ983iZar4fGoP3Gc8sDON
IVxqusrwDQBY/wKTK0D/mCdQS5rG4dl+Ejd0t2yigQgHV+95fNpkH0kOWMK4huCgayAdt8OFPzqr
QdIlo7aQyiaq5if7BGVye8xtZ7oy4kWsJRPWXXgBO7ZYIP6TBug5F7YyuQASpOOGzMIuttwk+VlI
IAUAoNTQL9F4iMxQbKOUgW6+iJUd6g+I66Xr9WZLC6UYpt6fz/OkFAEt66P4WbHQMxIrjPYnHKgB
jLcg6pAOAJ3eeZyKgf6ZNyhR2nXf+FIbFWuBvoLc9M961VJzZ3VuMs6sobCBFPsbC0yjsgXBeM/9
DwO7Fq9pohg1WfQZJ/LB472wMFqNlSh0RuP6OaS+apDKJczR0IMZ6CICbvph0IZQo4Gyzs3OQL8X
bfFe+T3BUKX+jtVR7tsAJGX6/nJ30aPLvNiZb+ai1WNf04II58qkM+2J9r4nfBubxYOJFmFYN7Ff
DFusMN/69Ou9R4DVcfrHCbiYpMDUw81/yqrMPFwTVbsCyU9HBYXcojbVyr2N6Gob+/dxrOLDXVHP
+R/O1LKp8BnucblQKufZks6zwksXo1Xt7ggDETDmGPeIKzN10Ql3uZtX1r65pZi9KTnVpj8ivJWR
R6dhWVISWcYHPqLGGmXPYza8ebQo+reBDp3pZIbRDirSUsMk3MWPa3wEWBJ5yOGwHh8oBgbSDmqB
6Xo4gO/YFFgItQyCJwnWruuJlDIjHs6q6T9YFIet/Sm7T4mH34G5SGyUOyLRal9eRbO6w1F+jQWv
/0HdX3cOTyReJ9UY7ASUHs7Id5dIxRRTkcAKa4wPHr5Qh0ftkwjcA3GTbrWF+iSi3yaYx0aNIiMo
rKaFzXZFnb66YFFHP82y28lkrskWlUXWeHtAsCD2PSU4K+mBP00YyPBxAmmiER83KdVe5xfyEEMx
dejU6DJpN10fnrvUjAsM6NRP8so+51WCFsGY+BSyIXdnp/t2mfNXfrWaa7EGC4uQT1jqXdb/kWnS
7+ykOTy3LaSVjqXlyjkqne+wmu+tvuJNehMknS8DvNOUR0RHmNREldWaOEI9cS200ecrdUMFWJQu
OLMW3+2+Iveq1WdiOWqnp1DlkweYwC1kmE2gqj3dQYsSVi7IIUA0hZ5VE14/Uvld4QO6qdBeJDJH
zpJ1YoM34fNGzupLC2Y9h5wwUWQCXvhmZmcIkkpDTrC+ivhbNXduU5b/+1Vmpj7PJpYRv9HXTIFz
63G0bsjXJ8dop6WWkCc1YTejprA7rDD+v0mAcSpHfUmfRsvj+c3vdH4LteKLJBlLT2LZMOsbktFF
NXgxMmG9pRbS1oc1biMQVg+vsC1rz8jScHajOBMhp6mu7kFlXD6paG8SqAAjSgqN2TaP/z8RGUiD
8s89bKttc4vPSEt5wNqehrmTvv/IhLLYPMoY3RqPSxxmy/1QMhHUt3hirmIfhlDfSq5oHQX2X3p7
jKBvND3BMU150CIpFOEWtdXQXKsebIOfIjTHWdDRYPbCRt3w7h8ia/5Ix8XsEFKBivQc59VUJukK
WqhnERP509zjTwS4o5gWrdV7JS0aK6hu0PvtcSAv7/yvzsntNVBlphrkYeKQTU2S7xuXfxed2QCW
wl+DyKoYWgrHfGIf5gmcO/VG4OLr/0DnS6siSUkm8gllAkY2Dxx6Wr3caBAqMdP4JQ/3aewAMWFG
bRIs9+iAZCmfTuijKX2jM1D06U3aJwZMk0nI/6UV39UMLELD8kExjzTH5Ps7ttgETlsgO657yBPu
bw+oOXkxX+04Ssbjb/PspzP6hhsLxwePNP1zSDew7Xk4PX6b0vLZggBlGSUgoe6WcrVUHiToOQbS
higL8wo377Z8MnomRVUc9CthqvYlMskjDCZBrREAIeGqv5TzmmyQoObVe12hcg0aMBJUBUtCPxAt
MRc1BeIKLhbFCYtuumY47FNJbBOmorPIhvPKp52Gd5sVSymr3kFOYYN1mwjFpqwVzHEOVwlchZCB
QkLT41alGRhCAmzFCeQzt4BK/9QwFG31g8Hys1c0YO8BW0L4bgvwLOkIbTJ9rTaLYc1va7Mvdz4D
mNTrSPfBX8wReI2KofOm1DOXaa6lZ9vC32ovlOd2cDzzB191X45VFimIIladGjPAaOL69p3pGM5V
tvU+tPme6M3jKbygqOxtB5cNwYrdnEelOdXlB211vcyY8aZWw5Fmc6JPjSyF6IiSzgFPZ6m9dQmI
S5Y13tB+BwOnRqDrNssdXSdv7AXpieL37w/4pN5eAVYR3+yv5PczVQOAtWOSkbSlufV/lRrcR92X
+JP1f9Gv4GPfmqah+kIcjGKhX3HRuTfL92cyo1eYUjHxbL/+OQR23B6JBcaRpD98QjlylF7IJa0z
umd3RMOurADRabyyzNF/nWVUNVyQ+FAJmmeelAUTAUUzUxuUvBntzIZ1BILHfIxbjnxC4NVHzp9Y
gpwR6Ewfml0/rxu4JC038qJ5rec9A2GTXcq0mK/GCzrSAJloFiL7eHU5+u9uwAMf9c4hxCdyI+HB
euDr1JS+9fmSPnDBkoCQNTxwRXZ3Onoj1jyyZQEVMjkWMsSkT9k6SAgQ+qbcdcVQrpXMvjL7AYLA
HzdDT4r+/x+ytoXu6p2GbWowtTXCr+H7KiIvnGYe6FNBTz1qY74OKO9yez8xsQ/N+eyQRzM7QxVv
PKsR1brsj2BQmyT4BtigR/Xv+R2mtvj+sEx3F0RtqsR84q4+AMwl6+6QAG1HCAtYRZaFwLnL4WI5
+Q1qbFAGRB+0ZHGoVtWKRDSj3DTmY3+wvbz/mu+bMyTlB6R1aaOh0qcCkpd6CNO/D0Xc1pDOiBGr
FIhIkD9ROKxu0CkuEiBe8dba7LMoBKOhn4LaUyFp37WeC02ATpkn0YcWM/V69G+6PCtcB3Iv8JT0
MwqRI9Kc5Y9GhOspiTSYIGkgk59jWNW6vPVx1c1pwoGTKARgl5PtEJ33B3O98Jo/lh9iA7ETYJR2
9dV5/fUOU0pUJ7tAI3K95QgrnnOsHrP6DU3r3DOZ44rvxVdnDmnK+7fCAiIV1P2NdEqHaGYHw/MP
jroO24VD1Gy5pkQaQWJLS3TUWP9Tu96t5liqHumgqXFCNcJaip6SukLL0l+1rusISTJN9Y9L3frK
ZqH8tyFWcT7A8hftf7YvMaffYrGDv2sUJXjDBXFy0g1ODOjEe6CdsSxwceAouLBhcYZKBIBVef4x
mKc/AggI8XqTxSVJA9CEkCwHI1nK4SIVgcY2+LqF+mhW+ZUm5IKcX2G14P/mAvYhpmeoAnMuhS7a
EsC0PjhzIWDpHLhg5EUPM4XQlUQwYycuS8mBh11/tGlok6D+csdKAy1M68IMLh9inDaq/ZknItEz
EBA0JzR5OwH2FVytRsNsqK7HCRamLhvLh7ZB2YalfI7FeS7gK2Hnq8N04PDQtw7+bqgerynhkNex
hSNtnIlPNk+H9OsMECxuUFlpzuNjLgMkTTzYPmltyJLv1JMRzK0c1gYLnKD9lNI0OUQB6/IbWpcR
wxcPrpHjlBW+Yk9AbZI9YPvVj5YK8Th7jTFRKlY7Lg7CtjbTxu19hPf4tAFR51Oz8gfXxnRVdpKF
9o00llaoWQ3KR5cFQetcCYGYjTRD1J+D1MLkGewNs6igDqAwnKzmQWa0cdWIyvHwSdn+PtG9JxH/
ihp/j4ZlZjBtYffUy3HEwV7d/2dfAhJpbnHCYzJdE5KFnqxxPBbgnIdLgMezZTZmtBxm6xAQQ/gz
SXNq6DM4B6GsjTPB7LCkV2Fe8bQEnLw2Wdy6iSmh0+Yp4n1RXvkDZBbRGm5q4Am5ui8s4xSczYf7
eqzIpMP0cDtgSaJz59E0A3W8RhVFTGhIrQk/hcTFxyhkLe2QC+vT0VOjgEY/gnmUdi+4/Afa5pcT
DwNQXuEH7S0gQ7zIT1+pdviiQgcIIK5b/L8SkJLB22xvfEvOnZwatdzjvBmdKO6j9EIupTATGCXS
eq+EkZp0Cn6yxv3MreTNaI+OR8+KhHzVetROeqMYjEB9MKoP8tPnnxlQAFnDh+Mtt+k+ki+x0TV+
8fv4YL0KLDhrC4rPXUTqJje2QifFxMJihRQCaj+G+4xwNcu1Rob4FoXJLYk/NrP/9E163XJQDDbs
vWoLZ66olhSElRflIBQ+wKvuWi0x4Gqv4+s87h0HJKHqZdIA82YUJy5VYUr9Fuhr//nMQUvz1IOX
aqNq50h/rVF90sc5SNBf85GpUbWlPxrkLC9cpB4YTVhnAN+B83RDnHFHs4HeWuRgMStN0wnWj8sz
QhAfevSl0xNJOMJv2nR0zwxz+VE4Abk8gMra0UIsSHhxgK6p3tvPsGJlGKZZtQ9ydY2EyTFqS+8I
4TIyxadLTJOIwJ43gsVOKkc84wzKoY0bBh4TF7h9PqNssZ+tnvR0unRiRRFj3KxlIBgfcih9VJHf
k8stM+t0Gh9HV4ASTx9sGkwosBd9t9GQVlrr0Ki1utepMO8G0M2GzFClz3p0GC1sa7ZlhbUxehp/
gaBElEYCHbd5TTQVMBAupqNNEcIfSm7W4KLvQo1me8uERbr4R9PTP5R+3n3yAE2dnvI0gD/hVyOc
uPTOp0+3qP10K2maLHh8d/3AiahNBsuYj9Y3T5IFMNL629oy4aHwJ9NahXgGh5y/xied8viZK+uv
WdTQcacFmzlbofxUK8FaCABTlYhH/SiMGGKG2cA6BuOFfGxyXyCYx3VkIp+V2am1Kb4rYC4A69Jn
Ogf/AE9KUo5eTcXT8VTGwY54pDj7ZauGtwKiw7ikFVRBP4i1kvKY5p/gTBfKpfq3JG+rm7Jpdtjp
4WUz3jA8R3l2AQZo6MKrEQ15XDJ6YkUOegSqE7vZVA4XYxaijElSsOon8wV9flgqiVeygycj5ld/
sOSSDGvfNzvh9o9nw1mqEahagt9Z3l870SxKewfQ5iICtJdaoaSBlymhg1WcwRqScAAGyg+AZTxA
Tqd0rgPVzG9RTblEdlSTzvu5G+cLq8depMYz3Yow8ELwG/Z+Y9aKPzRyHFYVLNfDTxMPsWSgoQfu
dKzCmFm09kgh0w5mrigJg63PAmQ9Ru4f68xqq6r+h/Y68NGTeYcTJyf8Wuq+xR27nWsrfrZrRIIJ
fE7nC43pHjRsXSvCc9irjezFKJUQzsNooeCmuUjcYGl/jFKrereZybSNTQZp0MywETaw6Ud3K0hy
UZH3FtGvm7m8VKZgPZQsYopls3lJGiMOvvx7y/h43Av0Wu2dPa1u+a6f9OCFDKndz+USiTloDxYV
CPzdgGEnmMwCQS+bLTezP/GdvC3LPWuL30yxV98pYqhs33tY7RCF0TfVhiLycK6mYGS10fHFZEh3
XLa8aRAgk2bNSx0koYSw3KNfPyXASIp50YQSYDxn5s9Elh0+h3FgHVb/w5pFuEyzrQ/5EcAV3Aq+
lPSFQp1v2v3AUgX+AOzSeQ8OnGsixRTFcNlC4pRt6qCe7e91H595XEO2w49ny7/HQcd8HhKNE9nn
/WlWFU1appOxOeLwJtGXTKLJgDyl4ngXrnsJ8ZEYhlcNS4VsWlJ7pxvgElf3YHRsjA7KuLeBvxV0
Yv7T01umH9UOgMxHDYiI72NWBtbDyw9jtd6COaiuAbu8yubxS6lCCVAoCcSBfQi9QEEMiKY+d8MK
9bK11+yJspAbSOFijHA2mDtLR8Wam+Grd6+7xc021C+8FWw2CQXjyrCb3wGrXN5g0A8lCXzW5w9Z
zDyTVAiLgnUm/eFjChodyQEtUYyFB1z0MZDkoqNxyAk7+tcOczbBP8GvAHgToQig3IDVjf3grgZ+
TU1EUBktZkJ6WLL9whzZaLGb/VHSfuTygj2UkzTMM6Oclk2L8183yn+gZRJuLkMsd+TXrylnOCGp
ePTffrkOEhRiLaZhWpO3n0g8iVSOX3aVSYyJwLjnxVplStV6yhEJTaV0knnJ0ElwFov+WfHkPyI9
shTanLpKrk0k2bNt7RhB7u+nhwMgtrNf4iqv6whIhU42R3aaJ/vi8c4UomgYRA91rj4qYx14/LDr
JuS3coajb+PX8K6BWm30AYdJZTAU0ebUEkhYNRUZvHenv+zWoiosits6youBiMFaxSSYeJ8ngRl6
RNYGMn9DTtbWoQ7BaSasMREls8ArHJ8oP9vkiBZI2WXVKHNC5o5kKUTvJM59oplWtq++r02YjHjG
vY8tbCnmhEaxycIc8EOlRVUnQsaSETps9YUHbV0TtzB4xc58H/AUiH7deAYFJZOqsmOoGTT2Hp+f
z+sZmRbQzm9eOL8twNSWZbYs2Etd8St/PJL3PbmEiWauP3z/mJUahDlralKwDtl02yflPbTrHZBm
nKZZP4Oz+d4GR9VGITj6DmFDpEYaix5VRIMUHtFnl/m0r6G/i4r6XLQ4RlAnaAQDD5xnaRRCOtJu
SN7a3KzADe4PS7Uqu/C8T55EkisD4vy/3dHI9ZhUo4S6ly5lHVVlZNXhcDmQgU98+XwYcJHz+Vfj
yzzZr9sTYMBAMig4BIacy7/0xQU1209JV++J7sAJ2CmXEj1tML/FWPqQmZ42xPihz+U7++wsqG4V
pG4tciJ/G7wrnulwqXEvUIcboqJxeKnbeHx8s81aCoeGl1pWI06+6QjobZTvObPEFN0iIszF49tp
G4EKCwLYSy73WHoXDtoo7tUTz0Fto+wNEX6TCxxnQ1mPjcWxyJNw6pvL7qBRCvtL9oFbh4PLnJ59
W6/lTEvGdaQuTTV89tcwPtgrTv0SgNLmYkZ7zqnqeU6B6UMLbqpe62/PQMvxmb6aIahmUQIXE61m
pfCHv6sPgHUk+PoJmQ7QppgA0zXafRKKQXs51LBR8Wc8H+d9ysi2XlXIWtjSJbBUPLyDqP9tf5lp
kFxCLLFsITM7365C5mwMlKRtMyGtHIZChY9IVmDLiyumetv8sh6p8JKecBHcd70RNwMwc6w8JJWf
CZ8s4RkO42x9Q5Q4+ldU4w1er89YFswwvT+kojLt75Zlya1Q1g5dTZvkXv9CCPdARqNTO3Hmatb8
lMdVMax/FkRIxObpVFgDibxBfYsKyYzBvJVx+xB21HmG7brqxPrMucAJdp8ZXe/vJ4xd9AZVwMBs
vx6xjYotlwocvVsS1OVM7mnwxih/T9FXIDa9FYKzWK6BozLQ9316Den4sUUip9kX7hUsl3dUzH8V
ZFXz4T1ejDRfCbgzXvvViaZtHAhgJXTvCQ4yZP9Mqxtj8okI3tZtviQeL+rgtQoMGtSpWx8ru9h5
sisDvKpLkVKHDsUByWTkc8tEMVxtWQOzQlJsloR4s5kqDBq8DUIuW4Eoel64Sph9Yays7enXW+3t
S2NHcd5QMiYKyaim3+y3SIt3XCJpaoEP6qXxwRPKmXVk5WEWH2v+YotyTlfEgmzmIQ90AIIVJygC
Mp3rvM3Sv/7rfBxeQQlmwJOTfzQz2qOlyLs0BFfyEVs1Bi8TO+EA1vo9j4dpMQ2Tb03OWu8OI2m0
wGkTI4BUbdycpCv6XonQlJlXy1qTxV+rST4HsjV4sakKqgokwx3AvAF+jxLtGjjzQsibC53DF4VO
X33tMeOWAXXs3rOkdcxVdhp31cI4we18o/9gkK2re1vPgiek6yun/QLb6k8/DgGHUGDnSXyFA8MU
5ZBuj5BkwhCMhKgW/vFG/59HeoSFP1oHPPGzuPdHAqOuzRxjUpo2A9WX+Bsl7/Xv3DyZa1l4qfp+
erWg8tS8iC5xrhaHab/bUf929b3cVpLtap1ns6ots5CWBnKennIPG34GDTrPaXXdCcs1ZLrWy9EX
Rv1ohemf8FJH8+aO2nhDVZ/c7EQSuk82wSJJMRnCrOmAWEAA1BUBOp0D3aFaUGINkjLog8ispnLC
fH02yKB/I5362VHRHMWiY0p1yfFk706ysoB+oqR4+/g10eZCMs7it007HL05I4RmP/nkjVVmrLwI
eY1CzcWM9dz9Y3skYUMHqbdZjkmQOvXFiQo4o8GNGp/1kxaNx6T5tTsyWpXIvsjPBe6N4YFDAsD7
xJRghIb8J8W3aeWzEkIS2E6fk0qJSmtMHmmFRP9dOrCSmlRhedS/xivFbT28xyoZZchC2k+nn/oL
U66hwXGO3kbYEDDb9819Pf1/JXsSwFq6jf1lxkE3YKRcb95r+woZLQA7nOnyp7dE3u2dOD8P/s+F
YjDMiPBGHceZhGj2JxlP1i/FqVCqHw/belngC602FeKcNk4LP5xw1CTFQLmV9WRUbrwcytlQsBTY
hFmF3cifKk55xigOXURXMkf3L9fTmEVyOSPUxpECJKtSZIuITlpg3ZAjAWIBkx7bTJITbP/smyF4
XfD9keLjGMSPGK1Yv5QrPC4zFIkWXOcUvIESnlWP+T8yLY4L0r5yhk7xgJrOvSDp9D9Ky9UtjZTk
sHdocKe8RQxMciekHRDToRw/uAIIjYo6zR2YvL4+hH3Rpw9Bpc79V+I99VsiN5VVUWkjOGLXUFVa
9E9I+Ygl+P7RFu2dRY5ZyJUoNP7VZKFODbziZqV0vrl8OoPJt5EOhgHG7K7TwZ7CllLxgiMSuY46
y90oXMKjS8rfuH3ZpWzAT2ekIEujd4RTZjO2cdAF4PxRq97MfiVpMrAMM9wmw3cwqy/uV5ZYxSfR
kxtw8ERmFz0+5kgnln3sLsP2MLiXhiFgHRS+Kn9x/vn46hdsOe1fEV/jlCRxUNQ7QubfpoN+qcd4
souWxtNhDp1QKwVaWLVZqULy9qMAckdezSGdf+OQTCkPsQ6K8DV86o4GSz76KkbngyrlHjIXF6ie
n576Z9iWOizqWI9ExI7QXnRyZGymo7st79zX3CJbYOcWcO8nwbTgzYx76hbI4wC5UBc1ILzULkFH
4uM2wj9LYlzHMkMNVMrWh1bKWYpRJ/arCb1d4U2rWFSzw+ETdGhFdFco2DkFK/3W2hIqVHKjdhpW
pSm7nk28Stmof5IIuhmAu64IZUCIPBM2vLEmw320uvnL6zWTqErVnrq3ttjPv2EymXKU9DIqFcB4
3UNcuuU7HmOY3/UwG+Htg+CZodeQX7OncC3pcmZWkyq4b5dEzhLK622RhgVo5cAymjW/pNPate02
tkMIy0uW0ar9yCxv7LxFUqVFX0T3JlElU7kJXS3LM7H01ihkn/2odyOkuMSCSjP/8YllEGsTpZzw
AwOTIPqD2P2cfoinuUWwjbJYJy9xT2jo/MQs9UGIoWjK0BlIeCvdtXFNQbzdRbixtRbeAAJCt/tc
xRR0dyHirRi+Ngx2jGDzxIu1YXwjFaPWu6FgSZKLIIvhQdSgu/jqOyaOhwQoPs7Ew0/09OZ/6H0Q
XdLg/ZCrn3cMm4s5Fy9dUIna1GCg+a0CBrJp+aerViy3QQzrAPLl78T+9otE2EA5KHgomhyn40Y6
ggsjLeee2h+pstHeyvdvBmQhiv4kudsilPwsdfZn29Hk2Mj4Ac7ZENO8FKNwznBZ8b88qNuEVw07
+mctr3kYpTFthgmyeMMXINioyXp4JNPQHhZRML6sWjXhTfAiU/Zp+EZ/Eli0Iy5oEyPDE9D4ndSw
Pr5R8H1s57NxjnOTeumnzr/kgOJf9hjna34SclYxF/etZSk2s9D34aILVyUliN7Dmz3AIkM9OdOy
AAW/Qm1ctNUPl9OnqoNNl8Azhbh34L7A0BK4vEC5E6/UGqp96JbMzCEXVqIG4KD1mWi07Qj6G1wP
mgFk68vPPOH05GyEj+P9hDOIgGj2OZzR/Gxkycjl1gJTarv1MwjI922ifpvRVveH443UwPAa095g
rRa+rg6d1vIuUdZo7yupdTFuqHX0/EtnjKTqkqe7Kxxm3bxvWa9xZQtB3kZ4XuGToY2HMk80aTDR
omakbVUb27myiMPtsmQUem1d7kuUXmJDcXeE7O1wAKRK7VdueppkMFIZt5w1M44DeVdIbxX8X5vU
wNOPJUHk04ttVnAncRO3dB+oYyJmFlydh/7e1yS07ro4sxTLj/UjL83i0OZsrBHoWO6o0hzETkAN
nRQiWqN2LoKi4ROGKUhi3HHw8Gj8zwr8J/6FUVBXykNaP3vEs7yEuY0Ta1HAODTjLKd0EwaISBNg
hbMP4kTgU2OREnMcTN6pQoOcK9winl0hNAIEGTcGMRQiE32r/XkGaHd17wLaYJr6Yo7khp/X5BcF
iER9DWPOclLklHpEDfmvmVHWNxxsd/lKO2e8YbHfFgVtGBaac/dJMhid0oVAKCe/TMB1xvwQ22ZA
PM0plgJXlhhRRhLGS1YOdbSVEJYpM61qOdgll2poaSx53ybovFIZu5P5U6H9P924AyNFiUIJlJ8N
GYyAvRNjzMLAmhNcMylc/Yjd9CkNXWFjFLnhOGXeq456nOTDq0qtxypUYgGgNvDn0JlMEaDkU8xL
86X2EAQT80d8ORwLMEyiEYiMy2erP5+8Bcwt9d0xVnoVj4HjjX4Zck4aOBjLmNaskZb8iYn0d2xW
SZ++jFroIYswsn0sTW0/Yo7MgvTauYm0i7IyMVHhDEBB57ewUMTbDHrKG9s3zamLLXclwiW5ZTAP
a2zfCEupmATMARjONuNpiM51ztGLvdU6Dx+qhiKxSoh+Tutf9DMNKN5JZqjDs0+WMk2tkETxJq8t
wnjgMMvU9DjVeghZfry0qD0zUjIK5Ra8beQsdel3MdMHKobIVXPZq3ZWidQUzPVxHD5hvfaEZEdJ
C+94zcukKNQsQjPPFsomwxLclbmKOSZXy/WzbjV4gRDm5UjSrHZIC3XG/EGk5ezAfbBIzrg6ku7U
UBB/VlhS8KtazwO/6vk4hZxJzXz45us7AGLBpXyRE4dZ38uNAkmwUvVvNw0WK0WgHquT03ZqsmUL
xqgEuhbrqWpsSnLvGOkorD/NujYttLKqgy2Q3Fkm9ds2+evmQe8AebIJeNOcWviglz2OuanD07mN
5hvL0yRUziTl/hw54xWAvYuXP+jYHrtjQLunK9rR27X0NPsIzclztnS7RtlPKzIiBVtUN+8nB2xt
9jMUJAhk0kEB0isIUBdVR6yD3OOwkswscsWqxtwUvQZ4V3bHCuZThUf8fFObQyBnHFIISP8Ttkkp
cZwRKPQadsqRQWYd9UBtZYZZNhCEP1h9Uirbw1hoDkLlPJjH2JBA2j8BpVq2dG1Srfzms1Twn9ip
vUeacve2X6b6CTvW8K5LHr4khvT/Qn2KqX848QAEmzrjLpSvSIYcwrFF3f9n8pecN6vHBiKHQqL9
wxphRB4Yh+SI1XY3Sk0B+8cfmdzII8/VUSsDLsG7Hhu35DZgApPB/YNXLsAu78DwF1SlUKeh/q+Q
AFwFmrb88u1CeX9CM+wdshfbMYXCWXLWeS9renhiS46ghG/aS4As74P26cvarW0M9Kqygc3mRy7f
31rZoM6vf+N2tdcFczNmtvWB6rlzME1QYQXNLh02IbNvjtAuGmL43+llglaxCLMmk8w0eq6E9my1
L22w+/pIfgzQKVDBFWP0l4KkIYt+6o11G8gdX+sm9xciH7LmlMG3MAGX1hj0eZUjTNntafov/JrE
z1wlyk2QV1UOnUxuLU9FhIQCiNWxQ8rhRrKasQ1g2in45PJZZH53BXotZNW901b4vDz/RH8rbNPY
FhYeQf8gAy63l+k00qmmeo5NNE/vlTbl3nBhqrAoRWnEFn7huTgbvqJPtc9JD0FnRqEimLgq53cy
WVgS2SBiZXNCc2ZImzovKNhdFvui8BY6ChsfIvAmWmd6qPUBIr3gnRTUBST3pTj5kCdMNx4ukmKD
++GFCJqM5PTKyp4LHb24JYnovvwN+XdAOyW8x3xexXOXcnawRhsNon0/yPiHPOnLCPwzwBUZMnvf
rlSirW4M93qe0d6dShEHKGQGsXsRe8wUeHucM0b80cQLzmzwiELNcNs4mqapQkvlWnjkXq1csC9Y
brjIQTrieRACF5GdeCMNVOku2l1wN2vwVwtVgJu96GmjTDbV2C8Sbf+HanmH/R6cJBJAyfr67dH1
Th0N7B8gLko8vEQUvgBD2QDN3xzFoMqORtT5jibqSIMk+pbce+RmGljVXXT/2gapYIMVEyG3jca3
cIJdq+y9uped4WW5qJWHrxElToKh2sRx4AsUOJykKN1S7icw1zyAlGv1/ECC1EdJ6V1ZlUw5bx1J
8LKlXzUecFVCstJUwq883RxPAWRge4/UCPAxBPfLn+FYEsoujPV5I0I+NB41/efe9amwX7RiCsDb
BUHoAgWjc0EtnIblVMX43Ng+/saoFXgTLufahcduC/ji7yVCb1otXeQG1huGDs69jfsYLu8piD+o
i0rYBmY+9jReYrfuQPwsYqLseuBO+SpnMS22QCZrOnwhmQ2vREnLp2ujxr5ZSvdVim0sQpid8VJ5
QXjcbooGZVwQXgaZ1zwKRDkGNcqAljimyzEW52g+6+Q+xMLzIkFCTx6Z7d1qVEvhjY02WgtK6bY8
C9Eagz/eiu1P0jWSP4cqPSLbqK0J+3AXnZu4nTEq69R+1FGgS94FX6iBnbsyCMnYdhdaAn0i+Ee0
MppOpMoBfVOnvyHWKU+/XPdIskhuEANYEyI8wKen7eyTd5oHghW3j7yGbrV3PnDiy9PhP+KaOHM8
+JDvl9gIIu4HkPzvpc4PBg8r/wWNHryft+90q3xJ98xEOV6AWijz4W3iYzUSRWhPQfNpo4B1gAG3
HoE6UzBPNUpcMvhiV6Q+570zG6ZEbeFU81Wzc//59EkaAt2pogSjBD0G6ijc6H4XYOgJUM7nEkuC
KV/j1GAV+Ws2i5mq1pF1dXZu8LX/A8258YgRoAaO9F+pxo91xXqdPvHwyl/hYnH7eIzqG+uuTIeb
WiUWcnYViDS834Uq7TAd+/TuUhVCmttT/iWdzYmcRD1hBUJ/AH4Ep4y9EEUljZ+ezqd9TIs5ULzk
nXgKm9B9N6s/2Q8LEN1poYWpYSS7SW3tRbZbVIRUvJ8wSBrJuGF5Yw+PVD2NFYi8rCFnb0XdcW0b
L/hpKtWl37nsZ5/gsGDd6X/iM7aej04EkgqwFTSkBjBiHdFCrhNwWY2w7x6GEkIu9eKtAMYxxOjU
e6Wk/Lz3+oIbThPf1QSmaftRZXwzIxMPuGoFFE3WP+IxfE4EjxrnPj3GBdzoWbJXRC6IrpUBE/xL
J22aELr5zBhImaJDQ4iZ6e+J+Ca/MjKca6xBvBcSFfc8qPmLNkj/IzN7D/5bjFxVBbh7l+DAVT42
ZziVxMT6TkZf5fNGuxrDZfVmNeIiw7troGdJEl8tb9NjcW9unCLZgQ1jAuFzTeOGFqyAT43iiRPV
7CpdW9I+pe5fSJ+VXjHdxiBmLruJX771oyTpiH0+9pMhzH1PKBva9hsdS3OJhIGExFKpVg2vxKsx
zJWKTr5Voj2y37B3v3proEQT7WCAvWXRI63hDpHwJT/ZQWidSwG9LWrrDbrDnPy6dFwGmCgJodvj
+GF9TKoIj7hQmUieEeiFF9sssAN+6MolHRLrR8+tUmnJNEgVJO7bkF6gs1Wh5Zbbbp9SOL0cU4dx
vMMCfQetOyBTzBjMDaoDAXdiE/uvkTabeABKjtsBwROYr0j+xN3s6ShuEbVO9mqO/sPx06k/5pSx
/Pt7BPhHeaZb5xzsveyzLN84ZeoRrsk1DSi9tDllZvySrNyNusOptlvBzadbAUYNtbBLzHGmUmoW
3r28YxaNAI7PBI4IjrOJMuZO0VhnBncDtD9NmrkghV31zVChkS3zNj1nv6219gspSIgVoJfNJ6aI
goirRdUOcq45Uscfhhdo1gAzn3VlKi3Z1t2qPjUeIUWx1LhbIeHf6yZ8TUYzf7nU5NQojrGe80/z
jlkPGcaxBcpdO29ZDlB3VoFK0J1aN67gzX6QXc/Fr3fT8zfzc07DFJkFQg28pR0bY/jHwNnwc2mA
h1yp2yd4AWhh4ObHyuYKwe5NAyoDnzpB6+FnKq0JcmTO0oGLqmeiUlRbP/57ampRMbJy9Rz55GvJ
+YOMvS/CsTIyFuFhgGIzgdJaMXGp4z9574Z4+ntAume0P38KmRt5AlqeAowVSysDVr8/GO89S2L3
XIoVPgtoSx2jWFeLBgEq54yDPluoLJWMH01mEELlCkJDlwO6hVyM7eyCkTAKAVqdJ9F1a7PFFCCE
B8engL7iQc990tgWnbcRMyobnjAADBI+rtjt0b5vl98N3ajzKkV0MHcQvl33L2bKpptT1oB9PBxI
cWFGJb9msKVuWpt009Gs7oQkmZzj1z7o2/8RyUvsYSsjElxgY7+AwTxkP20A0nlUYyYdErj3Owv6
uuYnCi7X5VDFxcaKExC2eGjzCKe1l4D5mRGM6m2QBcFsA3h6IB3U1nm/8cmm25MfqYG93+IjLJxB
EsErAhzEQNLyXoLhBVkJFqHVdGvAnqRbPlqsEFKPnhIFlPGz/UVBo+5Cvci1tp3r8KHDWchSAD5S
+8RChp+EzLvWhIs/GXAO7PxRFuCbzZYpzLxEZV35YXXOiRG7gbzCNCdyX2mlw+pUsu4SCE3VnDrY
ER77Z11fhQB6dsU2zOLBIdF+g9XVF+Eq6b74t8yggz5QDCYnu/VMjAGkrWc4HnXZ0+RkzidP613i
gKWH46+cntOMJiybxhqwNyWLMh1/5uduD0gsa1/J5RMgTOd2u0qxoiAzOVYXNz4hH6WLCrL9KKmH
kuLADbW3ilD4GxhcgCQPNYOBU/KRfyYBVBGpkpvdRykPYEiyC9II02r7QIUNdNJ2sn70HsxPohDY
kwynwzQWZxDRFJtA8Hofiy7eTdF7XY2sDBJ90wzPDJ2rpHI9JmlVOH9eSPckgC3j3fim6/0AT3x9
vlnb0YNU3YbeB1X07TnVhlWL+JOdrLz4oYuKTu8z4CuLtGwYQ2w4FXewA3wQ3HKxisiSbOyU8oQ7
2zmoD4XDt/5KJi9Zz3Z9SUfKOB2OhZQTr6wwSO0Zpf9+wFVm6fgWA/viZDI+Zl2FzIvPYaW78GM6
htBF9v0D5vxLwf/PHMaSMFwmma9HBBZyXIV1upTBMvR9E/pVmT9aQAN/pbCydsWF0hY3lmewAG67
LW2XP2CvIVmHfEMKh2vjbhj7kgNc7fyFy8beDgJflecnt2K1EkgkPGSWdw+0RKuDoBkuE8yMtnSw
+GPxs1USqekxB4Q88++lcktGkGkkTWvGzecnyhlSGc9gM7LSzlpPHwUYFMuYwH0dBid4dWUrbbeg
xRyTszNRHyHtJ05NSGvRwy/QtEUKZHcSCFm9Fdu0sdBom8V/W8pk2pizIMPZiqgAAQ6Yrlp3FRoo
d1TxJf9fO+zqm2b3uce6X3Fkdt1DkXk84NtHp7NxKqBKCLsv+LLWRbABAzWq3LS1hgWpmUKn9uhz
7nYxciwsIHIQXK6zLYEKK2CGLIKritvGvGjwxahwYSGKg06qWdIUpGSRxaZmBDzLYJoZl5NcdOqZ
vBOLvgujxDxP6uUiV21XdiL6AW7ZRcYjXDOaj/cfxzsi4XdMOzciShpQFDi1y9C8737ZizwiNwQ7
h7xj9jZ/f9c4/jwneVCU0tM/zP3bwDt7AH6t0r4BWuDSiMVPTmwXSkDYkJF2964HqNOZsa8heR5q
6I+1IUVUVPJQqOTghwYK5UEAigbLf4Vwz4lHHUOb0/iV0Zv8dTcTqKflpOyuy3HJSZEq5EV1JIk8
G7HzQ2+X94zSY2LA3v/xZ2F4SVkTmbvkdwTu3GvktryTEpD/HSbGYN4XNBwiXv0Mm3dwIwvajtKG
udc2roLSm4KBcZcBxUI8ckW2xscgxdh8ho5SvM/cLEPABM3QtltDRytcy9//cZ+MGlosiaNIqbfJ
OxP7o66hY6d1PdVuEMS46/e2LvqKG0RMFuhyqDtiJjk1SqqFWD/JlHShXN3BatrvfhsMM1vSJY3L
XUxoMtWXZa0rVTs2scFTiiLdqS8oxfrDFd9fCQnO+yckvw5ur0gXzPaZynPZmyEwnpsqVHh+rZZp
46hkZF6s3fCwckphYlMvcpz0dh2F0d9dgr0BZRwIbxW1fNPTuG56V8om9HsiCITTIiJKkhtGGCUf
0qs/If1Xc5i4WeC/yAjnXmbf+fonWJyx7ZwkQnuttpMPhAHf50y+0zaZQ1EJNg6CKFX/1DlnPRRN
QWIowd9BRjLGDhXE7J84TddX6jAsPc8NoV5psD9I6CDboVh2RGhbodscdTWtq0YFy4CkpdrTZ1xy
aJIN86QxIEShcYBljp26xJfjkUBj4ZEX4y7N8pmsz1M03aRBmzoQaYTBgb2HZhB/S1woL7hrw+Pb
kjpNohoBeYY2ZznZEt1lBSSy5rE3kkKlVcQXcP0PhHgeBYt10JmqjXohyUBYfzqd62vxgSIXz3eK
n3HU2z2DZFAHrXnqh44PV8YODDW8DaAVFdM1HAympGldRO0ibUeqhU5s86xTr/uDe/8mX9yFavvj
MGftiQFTE47vWLs3JslUV1e/D/EgQkTRccMTCgemkvj5U2RIcoaXqYSyfmGW9kfvLTqsAAaLXBVF
lI7Zvf6+shpYKqT87F6OehVzTLn4UHJXosWju6JUhNBO7XbWWyMmeuk3DC3qNcAUBV2yY3yszxsK
/OLCJWuMbb5QG8ofDBkemBv6Cwh6X73LbnBHI/QXzLXgI3RPNr8JdQ2fa24ZhC83DqrMU9An6rrv
EEo8v8xuCVztLztsoDrho3hdSjKbylkGxKivdrSQye/MthObETk7VNu9O0Fzff8j8XFoH/V4gkLf
MKJBBTfMC3ko9RwlGOzTioG3bZbGb/OOdTUzoZaq9GN2uPJ/5l8xTTkaY4KKSdN1I+3jJyU+Tlbb
Wl1KsuQ+OkO/u2sptfARdhpM2iNd2hQHS1boOneVjSTSjrXTqJf92NKjfUnhAvykcYWDtsKhKFIe
ZysUHV44NFpyCbXFR7worsnFS6/8Z+fVWbUBXmej3GM7kFflArxE0rJhQR1zOINNifqu93XGd8w9
udHqMQlJtzVEyvOJnRRJrt2taIpIf6aeq47BykehITBebf7QLdugVVu7/iZk6wtlcqGOj7dXJM3E
iJQCvZO5F8YH5MV/11D6sxzooZrIGjJnmmW3U+DyYiJhNzb08mpgu5KxGuGafqhcUELVSweeFnd/
LQFQg5ysn6qsEY57CXdQFNGFr9jUR73KYjnU7tdyjktIMDgyWXpxadX+H3wIFLZkvGlq8mVMFspk
A9RZEYRBxzXpJ4y/jU+m5P2z130iEXtlYbk47uYDMl3dFxaev8dSQH/3/lSHa2VgYBsXgO37kxhX
AQJuBG2bW+b1hlstkNcTIgBa+i8Soocdv1D+Rc/qig52HjQ9J1khGE/f6j+Q0OpWugJApgQmf/os
0pcORxK19+WS79qO1KBL4lWb62nnqYYs7kSMAawIogYe9iWMa98ZgcLAswY5xMLLUVv5uSTBcJJ5
FAp+wQUrzFWxxlUpZ1m8KKkUxKX50CQuAl9o1LwQiTMVNh2RVly/DdMwu+A2GPOZDCeN/sxT/pJb
qxvA/vCwj7bVKjDKsQmbn8T9XO1zoXGk/w9MaPTzgerkl70heX+1fuZ1qDLqc0YG3KvunDOrgJfB
xdrnZqrNvhFKvJNXNwphVUuSaIokK5MMSqEDNMLUlGexxMdXy+4hiU2WvHfJbzhXDbHCBdfC7OcV
Y68cs3BiXrntGNRXPcg+tBemMYDn2FCz1lvsEmK5GHsrrtukS2JYKQKevAmlgry+jJ+BYew9+ThG
h7q+3qI1mIe0yLpGgNqv+wkJ6kTH5yv6DMar7aoXguHPOskyC6k0l0adwia8QWAjXdUJo0J6jag4
Qvvl5xnMBXt9301mlK9WegtB9ncjj2NNmP2r0d5ivSWNoRHwJBf+FTKtip5GMLrTdGytu+0DDD5z
3zmts+9hlLegb3i37J4/u1p4c4QA5B0eG8RVrIL48afw3TUA+wUPdoB7I936r6vuoSJVCDrjzP2U
kvVr5eWza4cwJH1uk0skwShddLjBbWF+xYNTqXqIWBex2xH1J8aXn/Nru/m3ZH8n0SqStbyH1a1h
AyTA2jp6poZ2BN869hSur1FyYXJCUQhy/armSSNJYW+Grf11WggBziR1oxi7dBeB7Et7f6taj8Xn
bOnmvkvbykGexP5CZWjk70GJ73YXqxaM2OcGfsL6bFJ2hW2ENrGTl4YLwzL4WYMvi431wFkvGMAZ
1uENWuAVgVHu/O3MJRvhc7Km138EiZu8Kr+lWFIF9MkhTO3JmZ3x97IxG/psUYhUEz1pbBt5iqN9
CD+V37yCALBbfsSWqonEm+R/c662tk5M1HCA6EXe2AyI4znZCtmPEA25FRFhpWxjfyiqrF6JEPNj
zHKG/L2ld4rjRBMYODe7aoQGlRJX0h0L4iz35xihtkmXyGkYUQgLSZ2BLQfqLLMZsK0claAd4iHD
7SYp/7+DRMCcA4hx0E6QyJYcl/XjJ+rGJ6tHlntabrK2/J/VdZx6TM9gIHgZ/TSxabC99YKNwesx
65iYVmY48o0yvtbH/Flto5gdeUx8Ok8FO4Lef1/6UmqlNNoSt+QwS9ADidjG1tWsgk3WIEpDho+x
H4F7KB5HO+cCawIOV7QTdRZkidP3DlYkfQYpEYjiV0V8ei3pbB2AlIkxm8XZZM4RN33q9XcjCVwF
DZWOB8sYykUuvvFe8a1k7bjezfxz7JZyXAuTV8BmxlhEU6xkq1qfirTOnDkTDv6ja1vhnJwwGgT1
khoT+iDqdT+NZiVKcps+jV9TRrzNztJEVcv2a9HJfI+eqWLLnZZXLyfRtJ4FdUUls23XFXhLui2R
tM+/syr65joeBuIIdgcwsKfH4mJWK9smAP0MpMHhbwzJrW60UQHdt1WTHmncWNZlgKiiJaWoKlsp
NsmsI5wc/r2dJnm44NESvnQ+icerRZOs3j+2PsZGnGGXss0Px1rIwfzgZtMueqepJ1ETSvO328ft
YaLhrnQgNp+kPF9ZhTPUAzz/Ek2iJ7tMcc5pDRf2FASpJJvN6e61SEVgxxQwQbKlBHczW3NmoOg/
t+oF05LaKtFuAAMEwbhO0omqx2GpAyb7B5bjGrK0CzD/s2d6OwenDni6KcWbip7Xk3hpKFJw4kpc
Zjw3sR8GAEslF3LH3iZ2DuUEyaldUa/zdpmOTA3rZHs3SRxauIdiAhJsONp7A1UYKXoya7mgj5/H
tkJ3cutCdaBUdEb3a2IkmrmRFRxWkxF9PXXAjiqR0Aws4vuTU/Bdkz9njp7zt6Ws2HgFgkYaUNuJ
Sp6I7pddyj1Cp0cNBiX+xa6hEeowvSZacpAgn9Q+F+TAbrx6pqMJivHOJpJheFSdneDp7T6Ojaup
LXz3E8QxyrxGvkYBaxqMXK4+7xgnlI2rGjnH3H6Rh1UIl9ai1UrfVnzwMmy/7QENZeNXU/RfBRwf
A6BtH0DzjkyMxE15L8chGfpp6VhqqBZCltvIPg93x+QeC/1LeZMi5ZSaxlky85RwWrco46s5EEI3
eXc3+woC2czPr07Ge57xdNoovSupp/3iFd1i1uZ7E7RTsEFM5LoIia11XwHHlcjkPHsixkQN2NoJ
Ggbn3rg/3xi5ntvxlvaFBRPGwoeO63j4nfBLvq/gm6z+oflyMAkx0I7z3cACbYs1wQJDUfmTeGOZ
GDAb5vULPQGxgj0SiZEynoxOJMiiraq95a7ypkfH5NlBc36aJEYpt9wl1PY6qm/LBnkt9EBrNGUd
VShmGUIgcoZX/MUPU+cQPBHt2ybgAIgcvxYGaayEk+UW9B3AkO2ZFOyMp9vyfXrQBtcCFVs/owfV
q9FD9O1gYzt0v3frU+Qe4pOlg9IhN78X57iOSb2pFHHJwsstoXHTB706r+FNWPs4Hf5+6vNf0li0
T5oTSngJ/KwrbO6EfqL0rf/z3GVGbPb9dc4R63kMlz1RZ1Gn2MuKIZm9D7ybH8fgkCIqnykz/bXy
SaYt83052s38/HgP6m8u4AZlikguUufRIw4BQLaLrYscdb6bf/+3d6l4CmYmpFIVo+i8+DeIcJ5Z
m6RvI6wCggOPRtpETnNkXFZJFHows9PWZ0EBjATeDkQYKfA49bW/dSBlzRH5LDA33cdO4CPRD63D
S272ZNoSZPeUwgBJB2P8juVE9USkhbzJ340B0gEyMVLV+5Z6NgdT9Pe/jL/rxGEQTkNsMxLu50Fs
/DmA6kTYYaxt+tDfQId0Z8L34oB5T5rXl3AY/0JgbwdzId2Xie9O6Noc0bWXuMKF25J2qxO9yxPX
h0uojs9zckhgI59NlrNlVciU+Z17o9DZR283f+BOEsPcLvymmsluyFSaCVzA4Ar1zzPAHF4BD2/Z
PqZu1CghIadY6zjFPS3lWkF4Dc1MmXyOILg28H/MSmJEDjItoqwvNaX6z3sYlgHrNEkqEapyBAAj
BmhK8UiN49vU4P5UCDbnjzxt3fMSGcfPEI98vAP8ccCoHfKkZNGI4Om07STcbie9/xtqlhA5xvT2
ZbmyklxPFGaXe3GUsxZAg/DK6+8aNXq+cGXZ3PcmJAx2hWy+p2w5TbXf023AaZ3lmKA4wSXuQPJZ
h3ZS+ZU24+bkpmyyF9IGRajBJvahFS+yCI63V+WZOMDHE8dn/jllY4FU6cjhCJUZpPSB1MQ9R278
4mVIYEaCuV404lSP6JSid+/C7yEXW34FEphzbnx/xIGSvy0wo31INh4VA/j64tH8J2EFz/xJ4V8Z
UQXDzYCJKKrQny2dfcI+157sWLKvCRWI4p9XGodGWC2fOxmBpN92EwL+Y6PwH06EoQEC3cj29qVm
hPZrY2W2VMObNTXeYCfiHxAAR9UMjlV+H/wYPmjtUE53KDOqT1qvjOJIu/w221H9X7y4lYF3S4wT
WmmmaVYFhZ+eGZiawNCyRtMAkuI7hwpZdbLAKqOiheBb53tlv2OvIy+JzVTHskHYLhM9VjpASQgG
z0xWtLBLs4HFsWkUKID6sLWu2g7pMxTgX1vcVj0koUZRJuqiq+z1fBgumgNZ380MVpC3zlAvAO+l
aitulnUaxwjvdqXibNX61AN5+Gceqx4fD/xrR4hYFD7+flKw4uYUr3GNF7laeuLLUpYoD5Sp9nYB
M3gHkqmkMQmN2PJ4SibzSfUd2PQ2czLMnabI+npJNj4xlf8UINjtdrWSC41ZXSJcytIC5FVMuq6R
Fo6y7ZtZl/WFTCeEZeLDxva/uw4rCh1rwVpXXoqThIbexx7fLcm9yRw/MerDdXHxIYXOJoaq/Vo8
QcAFRbFs6VweMVMD4yJW5unobhWo02Rsd5I1xDgUVguH1OYipCFg4PSOP21Y/LcaT2IqZRp9C9Lq
Vqzp3uLx31ZpWNSt6ktiC15eV/4lmuW6aeFYCqlEaB+iH7gLMkx+Im2GfVNVmRwdrnsVlyoILChk
iyqfQiOQpiAeV1Je2ugILCLMLu3o/Yb6EvepXPbfnHaoj+2pMElTGgbWJrBIrbypQC/k2PeAPE22
F1WTBDyrH5oQ+vIoOK0Eod3rrxa3HRZnDo4KWw5CkF/FjuYy99iC49k0TJQ114GzbIxcf790pdEl
iYpXMIWFtCzFAhCWEkvsIebwCyL9gT93g5xJ1VqOZm8cGPi8Lz6zLWG4tKtEATJOaCMD9g4SB4ta
/lfhOe1YdNrNy3uTwQtYvb9n52M80bx6JtX8XAAtTaWzo48hxNj6kzyeESB6RtelE7cwBqbgDBjW
xxT4DcupPwtoGG3rL2B3qLjt9bDc2kinDCmBiOnf1TOjMxrbIkcDua4DMskkTUCT8tJvqKysqQiI
QWCPe7i2PVqhlALduH+jpMSqoExRRPTJ7V5+eqQRtrKZD843tjhWRjlGUCcD60uXHopqWFwwpN6c
6Y112VCzy5LSNS4LTJXku+9ZzMl5fk0G8UPi3qA0WFc5hy0XwIw33GYakIDiBoLPG67t53pYZIdP
0rbB9+F4DXMhknYe/7o1/PAJwjOeNxhtAfuvrOeM1lli1ZqkhEEqo5t60OORz6hhHbgJ+zwgTl6y
ex3VI+mIbBbO+MHf3m3jzmdgzA+6ikrATiZsvNS0wZRgaaGfZHK4Lib1hGPfNboWtfpYR/nQwBou
SL9WNMvv8bPnEolU4kWiGHOf4QVDaYoNHPqmpMVMjcp74fwjOylbCdPlxTzDbXsQl9C3kLMcgH/M
0nPYAsYoZP0SAauIqkPsGp9wcrvhWLeWzDqH9e9R1xFK+MMifoJpvYTu0rxYr7EL9CCChR9SiJOr
oQ+k0PlRRVNL9CmNXfz4ndqDFgCKdMYS0IDNgPXPkH9snzLBMMzxLSZ+/goekx1xIz2pKKMkqRe6
ew4tO+IJhy0h7JWFSU7kqii7fZ5Nj75I/YJ10/E0cFWwWFvusEqzptMDdA+fT0GM142BMfOrqKv2
IDtk9Vj28fSbFf4QyV+LalU8tWoMhDzrp9Fz3sUjYOLJ8Km0vqpapm57ikO5C43ZkORUM2Jha0Al
Ff1VsMgMpzp4YKj1F6z3Dnyn+Ov5chgbncj+okxngs9wZvPA5qTH91VFmCF+6+c5GD9K4PU4Xx5r
2SPlxhlAQNmJ5L6EIgGP9Imb2URSRgA3H5v6Z2Xlrfpv6tm1DTt8mr34+nYmbaNh0TDA9mpY/hrZ
YnMlR5NAVjwjljdmgniftWUzvnjN4Ad+F1FsZHiI94mMP3McOoncUrZKrXVMfI1uzukgi9ItOriO
QxZuW2gAS740M0YCGBJkF8ALzlCIVTzEpekx3b0BPmTJ3dLxw5B6k2O5u72updMMHG8Pfwz7jxmm
Dl3vVKiOwLM+AxWP7QFDFxo+LZ+4fGi9W9NU+9oF2T9rYQf8MSq17bac+VMXeI+Gnc3NBBG4L2TL
Z56QQuXvhY2CVCGTgWf08d8TAx0w9j84qOHfDoZIRm9zNx9amessp6zgP/KM3+clClTQ4v7MtRtK
TJuaWX9a56Dnsb+v/fZ+dyV3IXiu0/SMZF9Ga72xJ7nnbQHp8+OI1ETQwLAMSj61hJu/dkrRCYdO
rE/gSOBGwyJvyWtEfgYIwBwaG4o0xFGSAnPh+AVHzsf8Osdi1DgJ3W4lMwpkSUE2oZWOKNSEWd5f
B7ZiJT+dsaOmpUq4HwbcCeDiYo/8/dkOhyEtr6OWx5rYZOig0IH+XO5CD1+81c6RJs/eaU3g1QCv
YgF0I3TGvMJCKJP5g7jqvtZJyOmOQ29KYkTdD/bN/RKBnMh0b5eFrwuY/skxn1GV43MssvvXqeEC
UqvYzDtIeppAPXyeC038rA4sQ/jJJOH9UTgeqZGQB958HUpmSVmD7vONZT4fBubYrsRGFMSx2E3M
fd69kjvdY0Lfv4zNNW3ePBV3Nn5e3mPtG2pHtXtZkQtF0QIBB1UyP1gtlqjzEL386BMlA8/s56IX
3iVf8OBr4Qwt8X8XoNRiSBLt2jVCEgD5GI5SBwhztXVcJtC/b3vgwBxqjN6C4sfpAZ3Ffyx7Fcft
X6Xl2Ays/GUi+4/+ZL4fs3QktV78akBB4blBgo7sf5pSn9COhRwjMAJ914wc/6TJGt2w1AhLEl28
BAI3A7lgLjWPBAebw5IpVbsNlfcvy4QKmEiy8r5KHJjF/PPGxcsCO9UedbIYFj8DS3GiWa0MKQsE
YxTxYlGHVKDJTrgK+Pk+gx6c0UMiWU9Nai/DSL+um8AJwml6Rua1rP4OtV7ceEwWJl0xOD+j0Ce0
4KJhzKciho8pLJV1qPBRHseb8SDHYP0YEP0eM1SH5dxkWKwk7PKv7Hv35qyyqnqywvcTN4K6e9dI
3Hv8x3yerpNMHgAdAnQGlfSu2/dWI5qglFG4yRmWLJkisHtb9yHDb3x+J/tkmWaw/o9nQHH0lY6R
03x4nZ0nqDzX99hP6SthH0Y8tyzN0iOTLIgU4xAECGsove0eZB+VcoQJTnnF5MsR+47vumQDmTvQ
BgcGy1VhRg/qyDS05jh0tdh3fpHeJhkCngfK2cK1Oxv9uKGEpq8e9wfs17wFgF00sjzJCgtuPEqG
kDBwBqnlcscqdf4H+7xl++G3fIxpPJ8I2Qw/UxpTzcfl1KNv/9of0Fja01iFXXxePGaNPn1MgAOj
jTRAUqCZGKg3bpp2+j2nZD+2DUmRqGG0Z9d2suI75rQdkDRfqqv0IORxvM/MXZSJ2WBmDPuuf3JB
8/diUyTb+f4GI7+fNI06rN0H9MNArUUWyRgOJSEqDvydl3EDKVlOTM4POKD+KXmaYta6Q4blGx34
EdL3/nuaL45ilBlLYWexCeHgNq9essVkEqYKgfp2UP5k4ykJt4f80vJK+J+AZLr6M2NrSQRS/HCG
hhqqpnHi+w0MH/vxZgZFylhFShfK3ylkvtNqctv2dpm7K0b5Z8JpiGfeAlzCKD6PwCJcS/1tmfaq
zIgRz7kCX1tRtEvND8zd0qHIq1Rm8sbKiEQ/TmQ54xcmC2InCI7Rz6kA54dk6BSFGRjJ1/L0NCV5
bEYSLwXg7Hndhzr4xCCq7ek6P1MqKYfCC8U1Stqv+HSW4pkTa8X1l41PkcbjfP/Q1DKmdu73iyB2
vtWLRnm9o4R0lSZ9ZQa2Nl/FopDsfn80PJNoT6Suf20QD2A+sCNx1Rh/phHoG40znK1+i/15URB1
b2ECuuwtdyzuE118iq5m+MQYUHD6Hgg7RcQau8fV6TA6QqKj7UbjtQ648eJkaJeAt9aTff1hiPCm
7oJPLtdM8l8VZoT1do4AtOqhogpQ9GRAn8ca87ECB5+m0QHwrATzsG9jMtlq3lcD11SWBO0RL+nx
bm6RBj5U66RbF+wxRpUZvYXoZvOupT5SOpsUChzm8xMj5tilvyktPrzlze8vzw+iZm+B3kJWuvWF
zHBRdfc3wg9edLqzLf7Ik9ExodRTH8CNJMbDvqZNHTiS12SPhiiGfHUb2Qq8mLaWGil0GT+K48BN
mlpzQ+nrx6AXMZ7YCvtEQVzGYijhQhMdHWTbgj1T0XajW+noIsjWCOCAX6zOZTv/TrlDTlg9v8Ze
IwbPRqDjn3OdE76y5ag5JO1hJVEzBOqqpSv51Riu0HruEZCEI88c4HnFOyz4gPeAx30iywyJ/ooC
RgI6pfJl3CrKLnf7V70fodUHc+2mCGfxaLrQOhyfDS+fGel5oWhCToYVz5hykIq8jHXw3Q3oYfmm
i6V2fmV8m2jUnMnkc9LMtEvx2w1+4697GcPZyLrkFyS+MYB6i8SdQBbeRzfN0TdgxxW1sNnIYIzt
lQRFFZLm4iPNezXS1eV8UJouGetHIGb6OMiAdM8wCgY0jSAIUEq8aAj9fBLTfF6ebMCW0XXqRU8c
FkuiXr2M+Sw+2FNIosykHr8vUyeDrjN9rd37tltWFXILQO6ro26OIf8ZgTUFmE9Ep52/faDtXi5d
RrpzweOSYUPImFFPkkHeFEMNiya08/O6nvsilcu67ymtiR6pBDZyLSkfeFDThQaJfLm/OwKpxeWg
KLxX/umz0twykYkLeVM5VRLD1w8Kghius592apP0kTXhw99lhcPzOKALX2lN6QBd0+USlHrRJKT6
T/flr54NHdFdsupwB80WzSM0v1YDCekfFSSUmFNE2aURuUNt1u6mQIz9Fmc9sXSXs3AmYqx0xKQ6
l/z9ohcQ1JImxOIJbNbx1hFMpVEorrg30qpou3uD/sXTz+3MOx4/rarkbx5VDr5QG6pCyU27jssj
JdN4Ply2QKhWA133TiW4b6iTCKguGoXzkcGWrQbbA5jtLWfc6n72sufH9LQEfdkgY1TuZA1GGdyQ
5Mn3adzy3yPWaMJUehm5uVPRI/eG/VzJoxbKcZuWNLe6w1cyndi5s2kt4PWXb6AVWne/cfdGNdlV
zwjD/cXnxEPG6w8QJ+hvmd8+MpRuIjKzZ9ShCKUWy3AmA5mPMFiBNS70x8TyyRN8QayLwh0CRQK9
Kg2OsmrmjEqaO12YYMfF+IgdATK2zEew6NetL05gbNM1uDW2ml48wboXmIfRIYtQlNPccRKfOzUF
JS7NzthIn5CtpryGZbmPAGKT3JultvILNDTH6Yqfi1PwlYhYStmmU+2AORm6lJEQFYDxPdy5J/kf
SZRIUf2GaWuRLRh+QQo7fz0cWMRxsVMtuQ9NhYtjGbv/FhF2OGm4EQC/62S4eM6Y3EFwC48MfY4Z
dikokNJWE77oXRgGtWxjHK136cja/QYEoVdSGR+y/GpIl6NU7oWkzEDgnuc+0hOgnhGdT3jP84jj
XoyB72GEfYrJi03nxgxhkB8XCWuRFoF0SmOgWVFGZheQ04+FPFUthe4s4zt4R3isNkw27TTVN5At
1ZXsiYuQ43IQmwqR+KPZyuk8QP1hdGv4yuqANfx3Kvzxqk+bvno2e5l0KLmfHMRkez2gDVGk+1Pk
CzH6gNfeWH44Atog3kjp0C0f6kc9ZNBe/+yOi+eXSJKT1KsrobMViMcGwpLhWjBFGW/YtHvjccSq
FVV0OrA+KaaXTmqCs48q3kCW8/SbmAlSXr74mu4XFDt5a7iW+ACnUsaFCW4mZVeybCUP4tL+p8Dm
58UpJl2C6RgHRTF1jdQPH8knC3tVhazPAa3EO7yoTNBAYFjb3bYdheKt223LwywEUqFIM2UwJdaQ
F2Ob+qOade/4lYRNIggkpiw/C+AVGj7UNNur05c18KN3sIuNPZgmgMIGJ1NsPXdrm6es14gkUArj
uuH/LWn+zJ5dKDFRZkelSZo/8raR9hA072odoaA/flSZDElj1dQZnkBHelDPT372UNXRg30Bdr9p
3J7Zh3G8kQOFM0jduvjU+1dh48HfQV3+AVsrdituPKMbyzrL9+EYlVAQjjXziWukVIbi1rNzW8km
695xoA6qTXOXDbEM6pJDdiiLxfZSAm54XAW4QcrBjAlPgNCXkA9a+bl1SnpvxVgIgXnBSImKAXW1
CteJCI0c/uWMt51sjijYg0AIIuiKNCTmQvgy+qFwQMRk462aXunlSOf/hQA4tSjqXasgX37uKzOp
B6dHFmfpKA3n6gwIX1FiwzPtK0VBS1+jd6p2zx8FoEZ9nwLaX6GzHe86y8soewpbkq9HD8V/uOWl
7N2wO0CXx6lcFeTIobvj0dLZklFvmf3Hz0aLEA/SxAgUxBB9kESnPemzQHm6aGvdia8qzaNhb53y
fD83H8tG0PZoZWkTSNkm3baxWg4OJHpdRqVqjOw4dWyf9+cWL/NauoMiyb/b9WgKlUIeqPpYgP4Q
naifCXZdADTNaHcVE9h2SaUxweRzPR+ThhNAw6ROXYCmnqrL/jIN1EPLLmJoIGAx2TYxHHncRioS
TgaeEXNzxQHJezWXULAZfYCOQSccbP3eV0CvRsKo5/lsHF8ULBm54jI/uYes8m2cztqnlHxmUXso
Xq6jIaTjqnh/pKxQ9XnChXnh+1/6Gom22t8EidUFBvPayeKVARAFqCHuzlrzYAvP9dywI4WvavIs
PAcqTjEdjzxxjfgFaAXDWjZgsnuzVHWa68NNUkjsRIjYSjFKYHqKulhFgT04HI4zacHmVACCls5G
xbnqmdnysKXpIqG8ysJtapdTZbFmP+e3pWa6ETamvwrUX6Xg2OxQLKfAgw4nbmZVP8mlwv6gPfd1
voHseyADW6TJB8V5bLATt67WaeSkZWm4FxosqQjXst2AyxscKRG4MUutmxj4W6Xw3+i+bfG4RZq8
vR+vwmu946+91FiSIpCtcWgT1vqCIatjPlAwCOsLOL5SmVMDZvAqghtTjGTPqNKJOJylkiqgRSG5
/V8gRJV2XwlwLRkULuEjmlvrfE7aU+3xC5+3i0Jpp//e3+jfa0i65HCuF2ZB8wMc/tXJKeyxKVOb
Zo8pyy5NpGGodYNuPhsptGf7D/hVaWu/waiXi5ZTgdahXA9GN0hXHk/HXDnt1luQ+RfvbT2ttRC+
t+dJP2ESAxEo7X7D1Wq4w3xBG16m1LPtwutBY1f2cxU+sLi+t0fQYBZGGHM0PS+ojngt5KDvPopx
wUDZD/G89QbW0xuBGt2xvpPtydsfy/9rMKIa2/FBpwsjJJzohwa1IpC81DKwsHLamowU4+93Lcts
FRADr1Q5CMPen8h9ckZGEdNhf5Shv/ps9oLJtSvhPiGG6uA27tqAg32KbenjlzftwoZLgJMo+5c9
SSMEUQu7YRrwNAPCCixKPzktfZbuOZFeRX82RkYXVhA3ewDe5PgHlp63y8C/exYBqvYcw9I6uUdd
/n8aZLQtX+ctXVaF9fetAaze2cU4+0qHevacKPDyeznGT7DmfyDRTGtSrM6qQeF0HP9GY4f90erS
RK1YgePnB1tFUcOVAivecbYvyhFIR1Pd40tqG/FAP+eRU584l3STtPzxNMjXdb6pXampNEHfuwKv
aejtXynnkRhDH9HMBD1hPGHUBF0Ebn7tGx92PBew0cfUUtLVriUEJ0ywwqkpMVSP8UCINVWZRS2h
uXWpoOBXYBbdmq4gNXDxwXQD7tv99l346IRJINI4S+Re+ugjkN8Zs4iLZp/jB//JjqAl6mGny9yS
ZZwMM9VZueFYxUw4wbqonNUDzXkq5YtEwMi2QAOble3Yd04Z7E3fZlT/Rx+eAd2/fq6RdozirUUC
Ned9+8ySYFvflNR3QV9HaCEr53xRWrF4wVogG2/xpxU2rFP4lS1da8Ywmy1DMx0IDrliXISb1aoB
JuKW1TDguTXHPsQwHl0qHP1qKHRPffz30TLqrXvNCFFFTCCZQ2CTFeg/M2kb0Oos3pmMZB06qlvo
3+R1HPkC/Hz3bZHz7FYDVpmecJT4H4rZ3OPcJrSC0q9LfH0DlFXUEUQovyZ1VyXOSz6stpb/Vmtw
KotI/b+hkyNsD/j3zMbe99Yp5iQRMFXn2Mq6/iEc1klpSKZqZj5NQv2PHb6B/hft8yjrHl/xQ/yf
YqVx+EtMiw76GLYxyrOcX45Ftlj31etFYan/d6fzt5VviymzWlsd1gLP+PCCH06jXH3RcMteLX5/
C7dT5e/LfAOrveQxO8/Ms45nOF2vdBoPFfjDofnRA2iEBPP0/syKn5NUXhb+nElfkbctpyTMYrTq
TkWOzScsXzE55/Y9Ab+6E/fNXuaXq+yZmAXY4ZvnN/heIME0SQ4vraYsHwSwQ2vpvAVA+riw9U0t
5McJWY3+EJzfLC+KOLJXiatGeZj7vz7WWDbOlqlaTtqXDVLgb+q1HEjULXJoCfEsMqjcxr7BNLz2
EjbJcQGkw5hV1yxC+2pBQbxVbsuLCOh/Hc1GHcCmx/C1lHPEW4wZqiqBPZNTcdDGfEq4t3mO9Q2N
fjm/ztgrb3mCACIKO/SaEtkPV4Iw0wPGsyxRKb2yX1hxkw7UDqlf4TcTBqWIF1nKnzAF5f69TK1c
sNS9+3n9N7ke60OXdABHLUeCxmH2aJafg81TjkWLY+0wuRmPM87VA2jXXJcfbjsduniyu2awrzVD
OMOtz7Y9PXUqtQuLh+d0w02cqz4xEZsa7o2jSWwrshUVpGsvKCW0xO63fbMxLQzot/VfEc69gsGo
R63u90md63NqwWmtelbmcrIWhkUiE+74TsIShstGRxNX6Mt21yab32NXcEiaj2w5tkUaCcKKuwWG
wvuX8UghSUmgQ91lUChzNyiAd3PXzaE26XpT4B1Nu4z9lmqI1mhgPAcok7vtDZhNNe9tNKrUvEHm
6DgFGd+NGPFk3M5lYZFAzufCazMLEwvsFJ+A+xkdgX4/n37AMRGLZmXfglhN0cxY9JC7PIzSqVTs
7f7mkOB/peQrHy9EwEdttew4M2a7QewYk2DA1Br7KKFMuJ7MChauh6NBvDi3+A8jsrwLQThDqdQu
gPvoEX8wYnJqnUHU/XN+xQBsuxE7Qeep/2p0nc2Nss77ZHZTuP0g9+28YV9pnKkg881VTWbb8Foe
PTvUcfBlQqx1BRAydifGQetfHdIKlJ6z7JHtFyVEr5I2n04ZWbJA/l2IZtTvtwNDuCCrRaMBtnEI
inquIkIP2Lc+31hRiXjWNTzv64zW6Wf+kjrKCkShRDXjszBayrfdToKXcANPtXJR93SQhJMMYVYv
Veb6oKths2pxEqFhZR1nKSjmf5waYo1Xwo49FTzuwMOdgRiVEq6Xr5iTk4KRpUiWr543iOYpgzTo
iJd3jQQoQ/I6LNJBpTJ63+CwCfgrJGGqUCXNT28CRDtFSPGGxJlL9T3WXEd7ZrbHdGXKZtXrm4Ch
3Nrzz5PXyNGeP7mKLp+8VJLuLXq0o/jTGWtDCdMbCTHeyFA4ZeXcpJ1Cc9F8R8Qz0plLI+ZJLnv8
B8g+g6z4K38vsE5+3c1vC/ZuVwMzci0fE2nKcbQm4IJ3KZewmByMwYZCxdsRgPNNMx3lNR+JLtV/
x8qc6AY/t2joH6eftN+WRWuGe3caQb2S1H8KsNm60qXFIIF0nAYkAW+VsJPeL9EIMgKC591o4O2r
cjRiRoA3jGc7DPl86jTAU/XP4L8JP8UEe5bsT3/TYo88+lYh0mZ42KUPgUWZSPcuZDnzUQiTYGah
0r9ATXuoGreQ6lRGClTBJi0d9sX6d4D5s8kr7cQJ4evXMnub0gOYw1rwZ2QGxTJxnejdnAluaI3V
hYQYccwUQ9KhZFSYS+zGrlSY9yTl2KdIGFprzZNQ5+HDPWwYwjabbt1A/ZxSi3JTtMgzAVGm3JDu
CaHMXhhnnOhpQ8NdVqZwAyQCY0xXs6bFEa33ZdPvwUHRMEchVanFNJdjmBBmoAQW3xgxWlEO5DiA
glnkRHS92CrMYOnDmjI2ZD+OVbWkpjKyyTIMfcwP28Xl1YlZPgau+8bgIJILnOMXwc5Rh+S8pVil
v2C8isGtT4MgfKB14eXyo+pNSdPiS+BV46dqg+iDcOo3NxLxZSAGIuT11znSDLI6UPK5GZonp7e0
HQDhFmhBBtKTkHorfpFSG8W4Aqn7+Wx6w/bqKg9nXK/3plcw8vc6Z9fgBbpfil57BtsvLCTbpLd5
QO7fnqS8boTy8nY5Rk/Gm9h/sk81XjoH6eQMWS8cutiUOgoIXpBzPhy6IhgMnKyuZoISHZG0J+rk
xpT/jUmSW92CKn7cAzJNp9rxTtEeO53+O0U5DTImj09xt7YylAN54Isu8PtbJN276RzJpHis3zrP
n5AxAfqxlqj54WC1SfParNdlZducipZOr740wQa7WT+Hnv560Ju+x9GjtkP9ErvimCSINDUUuCh+
srx2pMYMzcH7cAe+AlfyjzQptl9EkqS6BfjF5vXzZCYmVfn8pIii6q+dTSM7AwtkcKZb9v5PDiNn
QEOpDETRDbUndFHv8zJ8VQoLAaxj+miiKHJ/tzngGVzx+HDflomzFxahinIK+3pWJ7WrQ7pzL3cO
yFRUFDmaqQ1dQfTrP6u/iWCW0VrH/DmgUv3Ty8DWFnfPxYbDxhgn5iY1T4ZTvEADRdx5rR+0Phr7
v80ouLQeJN3nR2ETt9+cV0wnPZ61twOELPz6B7LaIO4xrnA5d9NIB5DFwCpRsJbKpTM9ogzCNyqv
QRWwXp1QhYXl4ApyYUxrSr+ZB8G7gzgs+pcdT4sjsE8TeGRSzFZfH0maSoD57hGuz46D265YWYWy
UdCxi4mG5K+H577u1DuKzjPcVrD0fSpw2alDKXRuxLLxn3hH6TZ56rLnREG6g6gOPEyR9kCRKHhC
S9/IaGTGDao2l/QZp/8ZNmJOtORRuj3oNPE3deOdrnMN3pr1/i29ZK2zlYR6jgFrb3EjNlGUa7zh
0D51VlB3pHM3mmoa+4K+Pue5wJdJ7qgUlM+Fw+/Ao3oT9URkdGj+HZQXovPkMd9NxlDK6+8XTlLH
oWUvWAYhCmnEU0z0Z/9VXet8rci6+GXbpI2z6lRqHqGW4igKmxQTEy8DjPQwvUicdd+LzS5J11sr
Y6a70UaGs4c53TPM8qM6qAgWwuxgFNmyzPDjaoOArzPT4l9slydOsyL1Spp+Lr+HjPdLGuK07i5B
rSER0AaEVxsyPDZwKH9ZjPa12wPqlLAVUm1ThoWogKPehFQohlg/in2RdWEPI4YfaMiqNy9AY7Lk
3JYYhnz1CFR0/coVPo2neMKWzfHEq7z5ITaxtVE6Zf7227HgpSfS9aCaogDwQ8Czl7nCr3fWl6cj
Z1te87NANVf/SqX5Z3WNiuGfeB2lzsOzYjPUCwnCsnsdrpxwzsRggC0jb/g6843nppFvtLfJZzks
tbS8K9I6rSWSHEh9I3KJw+4uqMHI14odpPETcpE81KBGAtOzb/fAxec69axRLaW3lsGRzW1z0koQ
FAhQ9LnWiXxepTweqRPbx20rylNB6+J7GK4TTe7qqWmN0YXHJKRwqs00mhLri+zNyT95CjdYpkO1
0MsvuxUCDJxPTT/Jg2AhPN9jRR6qA7CT3tAweR+Z20X1RwGNpiDLycb1x43fjNF0/8QwFr2mFYoP
FRy4VrXVVNebhpoNgh5mpPb58c/nteJDyacGlm6hdLxJDFG3Ly3QkJYj+3U17oWY4N8gvCgsVX5Z
JZ4rErxvSYXTlx/so2alCQLrqlsISMUHCxfTmKKko2uucTYRJ71HD3AU7gsqQ1b1m9SRhSZQ3oLq
MLk+uXiz0ofTJa5Qv4G1nxYNoyRChk+iSE2o/7WN6RhfpwUYuGrLzCBEGwy2ew1MR7Tp1bXzpZIl
KvAxwmoOr9+MLFBGJFdtd/HsSkLrhuGyLA+Y7jnpATD2E96VVWvP1fB39fmlndrQvAkUEdXpzRCY
7T+WpB6dbLUcjkVnKeA70DbxB7nTbce43hYzPcet1d6bEgWHDUFhoXF4XMta4UGrqZXCGi9EHfAN
ExSfLCSmDKS6aSBQBhXhUu4SOCTv9rryn7egJoPMvnsuBX3WQlefVatWIfeuWjxcqCGPMN7iVXrh
GBizx+OJOSLO+y0Lk178kzEQBh+lKnyO4tDOzaYUBr9ppD7N7SwRCCmtp8+faU/jNKKILFN/ZHJv
ZiiLuF3eqLQZku+utDRlnJ1orkfvXapoFhH3rzuaMF+KwqSYxW3UuRxumVozwkJM7PqG81nhi2Bu
zIGmfPQoTCs7PFQKAzc3vr6+gGIW0u+eSaZNuk6TAG0wIt/gcI3l9Y8rxOsJtlKOA8f628k2Otas
SU8WldsepimaUR1hwPascnJKv/yVtAbbSkrxp1DsVzOd6AG4gKGQWhK81BclAi+JKGAwLHCpFMS+
cyE+E6DC561gSqhSMa7CEH8m16ZS80mMJK0YP1b4XU28j7T98OhoQS2q6mz2V4Vtg4E52JrXwZKD
wklg6M4wDnvsxsPua3LpVZ+ZndSJrlLfWujYld4D63OzY19C503CxJ4fTJh8gFmj01tWpIMhoU6r
62Aqes07uySJr6rj218Bd5fHEcQzXWdy6hqblU7tTHVb1NBmPcyBUBUDpdjaT8rNs4jzQLGTyc9b
7JKWwHSM0v8cQeHTYeR/sAKUOUnSpH30z3H+WWNoHimMZDp6HltQFizLcNqpjbm2/MUU072UOjk9
/iIYoSPrzTXgisNwKBqK5iVrpUYwijMRkqVldp2UKD1wdDSJ2BoY66IaVrq5+UfmVSQ8xLrXyyHl
ANsE9Rb6ZSjFJPk16u5LlUTWGKweHAu3lCa8PG0km0exnGDE8CL9ZsBGlQo6BFK4C/h2l6KO9BxH
a+mr0ph2JvuKs5k1QuUHOd2QoSAZLP3YyjTlHp9lMeZ32mrf9dnCzv8KNXlarTTQkglQ8tE4h6Hf
3ZMAPcFTN+Y1kykZbaIKBko6/BmH6+rAwDvCUREscvDMudFDmsiPe+kotXgAwfiFWuJ7jyX8uexB
w9QrFyI13LWUyevJezeAe2lv+/auv5kjqezgJypPX7Z6o/8pclqR+uATxb0XPAbgzm97JBw3kSeD
i4Y7Um5HTEVypXWK60MTEeDNEzWwTmnKTeklztz4tr5kStIG1G9wClSARo02DQE5qS6LfD5K2Wnq
0A+ukcIdHber+TEdS3R/w7C4N79KZFHwaee7DwDMWOqjbt3PK4g6oq1MBSMc8XRRXHJrNUTOpRqf
XfmOfSBsww5c+Iux+x8v5vZMgcnkMvpEWv8+8vktVSLywOyWSCVAfJOC8MMqO3NlMx/nP4IfFe4h
s2LiZ5qcykYa9ZQMV4cfrrWYhZhk06kq7TzjTk6O8QwjEXGXQISPBuV5YQAz0z3IhbOgrNvOmCkZ
eN69V8jVsYX/0jUY04yGassE7ihMGV0U4SvHVbmqpOpo80WT98o/Ufry6AZXJ+MKSLDCD3xZ4pIy
H2r1FRaRCbNwOBRFiFonesVCvv7j1c5WMFHzp2k57ExSWQhExUAxQgJM7VU3X/rxAl4q53y7qJXi
gBoXkgsw/HIwgBH0xFlPGAXGOUIxMcpj5u8tC1qlYqqNpmtHNfpXPrr/S5NtTdpYqTLZxaz45Pes
iIJhLDtg1fEk267yvfmFFCa+6VTsUtPamcbY6kR+YjdqasVqWlsYYUuOMd9xxMtDU8VNls2FtmMI
M7DYgtfZ9OQa+kfw7tOgSPxCE8ELRoqvC2YvO789VIWB+ce8o4/+RTV+hF+vcTwLdcYAf7MNmjhf
EZA3PutUNOg+2FJjqQ2Vov1Iecw7h4Xh2mlzZ7Rqkf4oWN/1yEVzZajgs5JEXs39RvUbczehPchq
w+7Um6YAv15m/gcO1ZotAGunkA8aqh8lv3Rud6JDEw/QFCfp2Vr0GAXEj8epz/iemI6qckoA9A96
h68u/dADAT46zz9HU4Q9K6w6aUAdnDtF/vYQUJ/M+jsUcWjYIiCAKy0Nw0oi6rlwhJqsj0p6vbBY
NTYMpCMfHOd1hGVNdH8MJXM5ABLnggH6wnRyfSLISxCDqRsH6Bf0jJZ8mUlRBtBb4g4mJCfEGXR7
HupAEulS8CmF7DlZXdtFm94v5V1Dn5jVq3G0LvUB/WVGRi6OXEBHOu3sceX7Wbluu3E/WgBUJ5eA
NckC63FtIM+YOTrETwotk9g60u4uHIq7yMNmhihA7IQCfi8i/7Z29Be2Xjbk/mgBwasYjIVegtb6
BQw5SBC/plLS6TIORJ+3i4dtCKA9yEZm8FtxUglAZSRoMrIz1Z/6NdqTcX/IxPEKFlQKK72KqACz
Hxbc7stgyoFkzfo6LVct+uV1qM0QPQwgfjw+IB4WkO9XGC6HyWshIMzIbQ6kjLoTj9/oOSxXtv93
kq5SEOtSZaO23fEDLYTsMEiaMXq5lz3uN9hiVs9NmXb9npCZ36rfr/7ylqubHGzIyXJp9tw/Xs8W
zcJdoOO5wu7NH5koCAw81DOFSQB7nHAZ3DO6+gXt7l3/ORgYJ8ZWw5loj2u5yT+20iKoUW+PjZBi
JUsRKmEDYYedHrAYG7o26Ta7pFYifDP8mPg6tfBR2r5XPkpvuuu/wZq6vnrkQRVWfMAkVYLtj+Kh
Kze+ZnoK6yAQ6Ftfl4f7WlfbBCF9i/T4gdLVFr27d6PNQTBKiHQ68hCsdhg0ABXPzugFzbbK7pB4
37BqKTeC2FTyyMD4KZyX1pF7LY+nGu79VYOfoMmaNUufsVRRN28I8ujv2prMqpdjMvFPRWP5gpRb
I+xnhFR8MHlrjP3gP/1uIn1Hvt7mFMiA3i1jOYlOP0IaO6l57ofzkWAWBupItsO2ZPan4Bnu7ZT7
Ugs1mg4HpwdzE/723RLj80/efwjzQfhBDxaUFn+Imb0AFJRbfKrArpmwBS3fM8X//1RKtVh7vqlY
1sfxpdQyewQil7TVTocgqv8wMLjr9cot1zo8xaAiC/DPK5weFGusfCAwbUkCdmJ6UPNWk2RpNOVd
IP4jeM1FyPgY56sBA2H890zFZOAdvPy5EOCj61G7cMINLu1SYD4eahXeMvjwN2Rx5Od7vuFqkqxe
nRiMn47BOltbQynA1mjTSusKoykvUaJDOIyC0Jz1dUN34yaISYx6vv0Xwx2oTcTNrPu8MRbf/T5H
xwzwWCrAMHwJ+RzU1fw+NNv3xWIs6YjCmFaibWLCPHiKiFdC6baLTQfXxwwILyOmwmL0YUjTBnKm
cUdqrVUUbModuqN3XA7uiOGBjJnPanD3rnfjRKVxO69iOAyii29cIbi9jyteEXTex+nePSqvIbtD
2YgIDLnYKVifAAh74hKYl1Z1CmY31YHxyv5DXyPeOaZQ0A4cIcsLRucAsoZaqYUNyTR3LfpufTEW
axddVKkAhahkuqW1Sj9KvUnxBG0Q2apby8zwPXAbW5fWuEDnaYAPyifV0i8fb7PY7h996cKGZret
6NN7Xk+nbrWITOTiMy0BWiDRJr7S5xoZQ2+b42eU4hhLntH3tA0Yv00mXuDSuXoruDCzW96Y+w2n
Dl45wXDy1+3eaXl3Xqr3z5PJO9/buRhE8PZFayRi2sXQ65ecu22JasY+gvJU9ckZ65fs2L2TK5ee
dBhuZY5Efzbw/7Gy0NzNHhfnt4T9xZzKEsMSr+fCYoD/yar+qktNQx997yjyqD5cB3/MnYleigM4
esNpY03bztFUfVHH5vDNYpbLXSSzikj3XnIHRjX4U9X/TNocT80dho1YiwgNqX1QAynakfopJEKb
fy6Atkvcz8ESgVeWPMY1O0+JvmdkMZK34WuAkdGWVYlvUB7FwOmUugzAKzb7ysoS3RbXmK42y1H7
DZncexv4T60z8MYVApMVkgdAotTvKAV5fh2uoIAs2slot46gHxhP0A2D5QFam9bq/xK17Y4hEDwS
PSkHNu603EcQMKw69lYYLZivztOsmoXP3gRcA5O59AylHZNQ3y3gIE8fCXp2Bmen3f+ohZOJfWBa
2pQAjV3q94E/2H627GGpssHqBBJf+AwOqt9r8BXN8/9UU/ZDcEMCgARaM0Jl7gdNJZlHdRytQep6
eC/lclUZhjErTut7kEAjb/qoSArJ7vIDp2chTNyGE1EQdlWZC44rblFWB9GtKiz2juOEjq7MqBFN
oAdFRTU81P9TZCneX1z/RoVSB1om4aM+o2dN1T3sqg+ugYDzyGy16QTM7fCjJov9T2c2GnrXMu+V
4CXtyADBGgt9dES43z9T3ND86rpJ4cpRAbe0wWL1mnvWlBdbJvrRA+fMTJ2sDuwRRUxLddrb9+dr
C6meW6/yTLhXMVYOZv5Pfnwz3NCtpR3qKkG3Qdr+yfIGigeAbYxuReY17dsgqo/vQgI0A+2ZmGjZ
lw93KI/lujjTkMkXVJpVXAvb4LMX546EDX/swYRZraB0z7w0j26HWnJ6EcVTeXAF2VpWSmxHmkL4
fAmopV7Rg4PWwt+CEkF2NgmDAnAYDOr3vW0kBiHG2pBBBiL9VU6r+wvlJVQaTW2wq2QGoSgZU1K8
UQe69EUpHdfbdcRFFqO7ec32uIxF5GXBWHyV2X+SSBhFRYgCRnzsnKiSQdSimdNVOyrAtJLe5Qv5
fqzIz9nt9jt8v9SxJilG3L1NdnfbRlKMMEga29CV5gBhcHKEg/R7P8dnY3OiZacfRpvtw7LpttTH
6N6fW1N8S9b7IPsSTZD+K843Y2QBVzZn16pICUc7GhTyOFVJOrJFpedQrKwnyJ2WttGP3I2mWWRM
qnOOECHmpFjY0r48qvbQ23GQ/UPGapqEY11t5Ssic+lqIH4T+x3SzgJEtPZUHs5JU+k8e0AgyVtV
xu+msPM1zpULyVJE0CNQZe5N2ICyDIxtkrGJMk8WQIs0b7MF9EdaXchxtRvBrNB+2ErwLm2cdPUJ
CGUJpCM6Q2Jca5vQqaC2kK9Qwbr8AUnLscz3qxdK1Hd2LxFzxQSA11M5IuLWV+N6vAXQYG3y9ShO
sAjinput2cE4Iiw4T6jd6UFbCIKiD9xZal9x7q1W1Tq4vmur4Rt58vjkIJSEZfJdLnzA4cNHRJKH
kefAjSl+Y07BAeSJKD3lefrCCzjsByZ6VRKcedd6GDwfxJKy1VarsLFp+vYfIUEr/9RIXv5setfi
lDLsX9m6buFC8e/41jUFB64C9G2Bsw4biHTu8li9jcEHgVYjHZvqrVfRijBd5h/4yZ8Yq6d0qbq/
Idp1PHcDp6tnYJVOwZQ5Xvj34dhG8azvTLqKhRZFBMdnBev+GMO3UjIMNsIr6o4U+x1p47JRjGah
a8NFI+/1Eljez8tuGOgVPDA1fkCqFqJTfDs+jQT98rr6akWkRNpH5z5JUlBg/7fPdRrgObpYogE1
8nRd0/SLnz2/SYN5jUhEfCA4P+hbiWY1cemHSqwgXcASWYMfwsoYeainA0TsoHcNN1rmNyLIqbS7
dZY0OQFmOvJHMeYJ4F53hdPdsEEjnExXXhjBpXBwpPwt4emUFnx/uwyrYbP6QCf7a1keGi0SDFx2
SW57pOgGWBgFmOTMhAoOkw5bZoqcyDlz8uB3G8j/7jNPx42RbFtaoFbORpTg8KjLWoj5cd93bQXi
nCBA0vVIE3sFK9BMYG9HVH7TgQVR++l4j+rIvm4sH4IWROTmzR10RxYT/9HhOA67sp+y+qOsZESJ
l59SMoNH+TSUxVbdQyDCxXvjLwQURT8NOhUPa1fDbW/apbIDklajLsdK96sNyKaMcUYqQ7f87vYI
ji0+EsPfLbpRTichi02Ly/wsoXFRRnAXBIoPc2qU+40XR0XfuzlBa4J3P+tvT8a5rDI9Ysp2vRFQ
yvyyLTroU6uvF4OUC/08jnM8Pr0EGoNOd1hiV3TCsEqLgZnhiyNRRFfjYiE1l5aYmpH3pK1seAMO
fCp2lBWj8qbv+mzOMnIofWYp2SfH+yWGPSieLLOc4cQ1Ii7sWerlq41faE3Yna0bh65tRv7JafNP
OC7nmBmGZjlFfhzsmbXUD3JEakpkZJjicW2dKwxBPF9cf6BMGBDXfrv4+qL/NiQPZi2y1H64TfXF
BBEThayNuYkXAd1bBwXv8guNyIiL1JFtaopa6EyBDy8kPK965sIwdds+Pqj2/RTVUfG+3GP58kdm
JO9XGBLMEWksX5aCifxMFUoSezuMHg5qP1gEg/yd/m5hif5xACaXPiRWHoC89tTBVpWCcF6I2M83
YleXxsUJduIbZ7KQqb7zmmes60sY+DGeBi73Ko6pZA+Q4yToVWh86Uu1hnpVXU7TEnOKJKfJU6v9
/tgEkI1/dz8MVAtao2DlDhWYEFG2tS81KxTV7EJqu1nuwm/Z8JH9AJojR07FPmwYDmMZurt0WBUY
gXKmA63g7mSTLSTqwYWNzM3a/inB3zMRqbmPdqhQuzUTUeFZoS8I0fZDC/XSEGvZOKL6PUHpE7n9
HcCXoL4VRNf1Iwzx83IwI2AAGXWjuA4rboid09Fs5fQfFs4lKQQPLSvOBNMqmw2/WjRq4oRZOOk5
uMuNbEKmCsQzhqru6POkHb0jMmce7AjelhMvPuG1TdqvKn+6LvRfgUtfLo6CaF9O38GzTh0Y36YX
sRvyw0iyNmKFWLXVMpDgpEVvKK3Jy3J744YvaUZy+TMNawqBDTg+xvI0dtV50pg60wORoRSpEani
g33Z78Jij119U7pSXyjwhWaNlDNOILjcE96AKfpqx50j0Ip0OVWxPTsoezz97mxqGFbx57p/Kgcc
0EHUFkDQDMSgtFAodo0rjmFcLRhIMVVvQyrKTfoXSS8Tt6Fzl0MlURkAk4QtEguh55pKLN0CAzNT
INGeuwsAZK2WN5KvUnv02+Cfwi26DoBXrlo3ybVXUW5Vu2dqM1REd/tL2x54MOiG90KTGXfwEMJK
vT2JIo/DzCgsVeoeacx3SoYwAyPWK/sJbTZMJHegToSG7rXcNVdHDVLKqQy8p2NsxS3aVgk6uAC/
M8DltvJos9lWgxcImEOlvjSrsJD7T5j8+LsCFZNAj1saP+F2vckz1vgtzGjAIQxGqV70CkBsckXs
D2yowsvPYjdJlb7F6ftRA5vkWd0XnWdjSSkjJdYgCnhJMr1gLMKGs5fZVr0rCRBMpFOC0E+IMxyo
W55GEMjsS+yIxQfPG38NVtfj5DjLChxNQt7PWozTUQHfxU06zg6f+3qODyt3yqw+ZSLjg96XacRz
45cKhf70zK6w3zwO2DEMqWQZ7YVTyK28AVcEudVUFwU+hWw62plGjSdlRjyl3PDy9XyLcHDHHnvk
WOUbBdzjXAdSKco+5HWSZgz5Zp4RGCP1x3i69HkDxIkVoaLE8IIccQoZbXvWPE5wW9JGfDNBBf7J
6s7SFMx0dwPOKULukjFP5xTh/PgtaVFZlimKIyW6ZxvTHQsvEztPEi55HyxS/Jmnsan8X8N0zRGA
PtwCyV9Rad+M1F2y37g6OOTH4AqGXUTJVjEQ1CRAenGlKMcD2/3y8zawiAXcigAqGTbIfQqoTB9V
jRsEzNoW3rmZ/dr/MrgTk9lrxKZR1XyTL7qj0y8eiZF+CZugnWOwkyRFBswzPcnefMgfwEDto6Xr
zEKa9gkaEM5CYDrwLMmdx8JVJKN92D6PA4Qn1a1Cjehr6yfqq2k5b2G2/Lr0wjwwDVB94vfyAfZ8
/WzI3ClMeAHcXu7Z132ePVDBXT4iQi3WqgoJf09wefuN2q0PfbXqsMDJRlMeSXp/IMkSTiLGlz7a
z1M8ptvECuGhNm+rT0X5f1eQtkc4P4JYDARmnbpgPVA1mS3P+UIcalDuXkWD8eWE7YQXKZZ1Q1tb
zdwZiDJ2r0Xe2Wd4TbgEnUN7QbgzRy7zrNcGjpD6xBUBri1CS6evyqaXZGhwhoHrUjp2SRnmZvci
hA7bIPdYR9LaMXKYZ2VBJEgzAhYv87a4ciY0Vy/yxwmA/rY9ZCuUnngDRQ3kiH7NDAKezbAaQIFs
US04wu/qCUS/mS498j89DFiXhTTCmnfzg03AoueTTQBuoYoAdz4BBowgz7SJLv2ghT5UeUnEhddm
aYj/YKU9v0dp43G1wOrfiBXJMHgdndK8F7NfRgBY//79yXqEM1UCq7k0rHGlvPAnq1DJiYcbXJC8
u3UGrEq0wVK7101DzgkY5UofwKcorYAdBDEGD/jj7oRN4pRZveWR3rWyrjVuF5ke2+Zh42sYyD6H
b+9XO+G5n3Z5PhZDP+zLPrP9ix3gflUMpOimgdJ3b5FhW7J8g0wptTEXnbRs201t8tuybp0KZwX3
AQENb5kkJVIf9dVXCBCdFPKBvMPyhSUkgsZQTtCZdh636VnrJ3ozHghq71CAH0POBE3UJPQKiBEO
IaR02AJoFhE25kIuDLSDDRqtlODYtIsFFY9ZKr/LEp9c7KpFTbTFqzQXRiwWSrNobQAC3C2DO+zc
MjOU4CBOL+7YMBEpgmtC9ZePq6JRPTNMUOtMfNZ1ouRPBxWdAngTrd3eeWIc1igAYez+qOclg9a5
8DtxKqzXuM6VHfWCLBQU3Tg7hOFsljvwf03Hjt1SyXIf/N1Ea0Fg1JLeOYDNLq+jWoeqFCsWh1aK
qRx9a7ezUIsYayQrrhc50QyqE8EObQ+QFpNkey+Qj90eAu35ccaMvmdzO3yGkO7RPiuY/M6MLJu7
iwgy2fKiOJ+eTIx5PByOgp8EVg9/3k6j/mmSeUZPMIYOrIi8VJpKgi/+2tL3f8DRdsOJdjFsuHOq
iiQxUMT1rdw6r5gAWemNM/bZtM1Loerm/g+iSFUhKoVOsg2To2zf9VQR4CGScVtO3I5eT/R/ys6o
9feAheNbufTjIDVvND1+MNWWfIJEQ/C3SGuAOrTNfCdaRDwVsUHh9DWA8G3uEgslU6H5ZjlYrQxz
GAGWBlBcnrpQsAZNYBdj0V4Wpn9gRWP5qV7yJDA77lMuiFyRKWaNAEG62JAV7J4Kj9PcJErjTJaX
UPkdITH8DIz1QA9pIkJaao1v1bVDfft7JJH0fhj3jORprz5J8kn5R6+A+tasP3YSVi6D4ZZ1IRZq
l2DSd+7vosgUr3xJd1rgTDiAij/yxOqBuB8Oqw0M5cmxn31DOSk+uqF4lR5e0zsSeyU6uMn4TWyr
RJnFA3Ryxbeym+MMUjZlk7SrUwD4j2XYtoRpQiuSdfsrk1Q3FvjncU7CTjnlzuJrRl2+69BSCruM
PsRg+3MFqeT0JEryg1n8qbQdMq910685HYpQ78Ve6lzer35dobv7lKuTPbsTtbNRPpmM3rwNVLUY
8q4g6+JrjzqGkpVxSESDDOuRYVM3xnBO0kwnV/sR24R0R0lOo0nqXfXlj8J3dKPYFzsIT5T91vCO
q0COVD5vkkS+FUNwF22sLdFoU5GEHh9lfOno7jXuSCfSgeBRZuwJGpTEsSC8IlwI5P9NRWxYj7km
aHzdvuHxv17f7DPDTZJPTZJa5BZfLdAWaaSFRaPE05iuvsvG64YfHllGFBey3gsHAHWPFhoufkHs
4Q6D749MlWW+4srJS8do7oNdk5U83c3IZcLRMuskwixl7ODLxigMPx4n312BaAk7UICnWTy53e/x
aEMaf1rwBgI4iwBsunlbSs99mvg4L3bXt63KBvCu/n7aOIh44jw7MhrqXW9VZbjh2dr/D3gO2kbL
Vpo1jNbr0de/yy6alqFYSyRRW6mp/6tLYCxberiwXjZFgntbcAoNh8HM6INNr1ilGzChbph6s6T7
zPtD0qMQczQZWMiDRAw8QRJ8KB3c3oNmy03xcTuWU/7SGmz93JG1npOxEwR/AyXPgi9rxb12yn7v
XKlM7Nc5GyWFtDxV3yL2+jBCjbD+OjeGlKTSeuXT43hcu+Y+hEtUQT1PucY61nXlbK5eYSNpLGyG
rtJrHsSgO/b2vScDU/kUslih7Iuyrr7FDvqzuNyhagurb9mABKmgkAvVbuCgrevs0qlwnIUkvMGY
ykydcwn12kfELrVtVCk8GVoF6Q8ujYXCOuiEc7sLolkWgDF1E3NbeeHUToucnAh6jM68x9HlYf90
g4qRbC1jZQTKydiKL+3SG2c0SiiyM81tn5mdVhT2/zcXq2HQAvOmPIRAI23MH/cQMkBLTxk/Neky
9lH0SGY3LHQpfJJzenbch1O3EFLqwDQAZrcVzMgmkC/6+LTmehqmZFAJ0XGWpgVPsQOSSY5lfx8e
MaerVsZFevK/qvya0GDcUH+kuF/c/KjT8FjKP8ZfMyibd6/M0T1h651BSJlYZMRKysQ/S+Pr5Slp
9z3f3XsUvnRgTBjEIxaRgIsEi6sagCV3fwj+t1hzm8wJJqFY8ErmqPOLSVmk/wpihzXlA+/WuRmS
LVxTpFCsaYjzzSVLK6gajOnC+pfzXGJRRb6fiG0duOIOXSn5ctQHVx5Ol5D+0MCdSAidg9ra68tP
A5Vs3/E5n0ltq5Dw4hC8Jg6J0k3cKfReWNpQIVv6Upce3iEVTTCwVGcg5Nrp2X3v1B+LT3fRvBOL
w+trRroew/EnwxZgPT82tZIkve71wGSIxPq0Dx7o0rZVFFM77A22gWOXVFNbAai9cq0qOtecDbqk
jZLNSNAfXi1Sksc87jT7F+Puf5chwUKrGEJaPm90ox0dXDzuqktJqFJpRXUqqL8+R2+jU29KVqqc
OFQz9X4aKrmps/k8gWdInXnj1j7ypevokD6jYWxqrd8Z9f0gH94cXbxutqpfN+kzw0JyXkrsChBt
GAsJmeFw+jSlRJd+ft23iR07MIhNzM5wj77uyDDMsysU6OCI7ksfZp9bVHf/BsYUEO4mg2O8Xrth
ReWacIhoySV9MjaNVa594DdzMBkxHUrNHSDMguTolSTukLmjH5R8rUIclynd/JiBLMqn2XZY5ZPQ
UdRK5hme1Tsg5QpE4Jnbjd4Ztbu6A9rRE5whqp8bMgBHcbeo1R9eMP5Q/Z5AxPKezwu/984/Vc79
7qaxRqwT6dqYp4h62/f5rSfdD+Y+aYFO/gYlHMS0IKuWdtiX632WmTU/bBIw1HqvWCeG28+/U6ji
aPJxgOa0TRuevnQqKwoZ6y/Woeven9H4ukIpuenyrVQqmQsK2T8ADyvgdbRHaYjs6RANJRG7LSKM
5I5zuE6IWQs/wOyiIL3KBculgbHBb6ZZuIB/VBnNCFo8a8n47BVM90OTc/ogiflphac0z2DCQ8ml
8FJ3jAfZF4vhvHXTASXg1kGhQ4f4KC79iz3o+JL6AOtMp6Vlm33tKeTGtcDUrKRasgxApYofOjXn
JX+471eYKVnfXcwoM06Z4v6iIU4W+1mWl5QwFtCwQJNFiqSXQ/EeLhbTHVj8DTbNqwcjOrJO+eR3
wwOHs3FhHb4joEJO/3fqDDOjmu4NX19JCeWdh6K7evInwKgJRwL4L7fznrsVQ041NAy3WtXw9TzP
gz/+6KZ73iI8Ay2dxBGzMWQEbjYCGt1pCpAgAA4KH/zv62C8CVxVcxqaLNsH9Ndtmp6iLxfzqk2E
Ei7QVKdL324lKMhj9r1qn1BGp3m7JwnfXzLaUXxDaIY7Ddn5dIJgwqOFMJ3gEs5R422ToEGhycgA
kM4NARDBsfNF8WBpChk9HH/bTa1hgCIhYYiuWMEOD9NzvUsVvlU307Oo4T7Pf4s/jeqWd/Flxil1
XSbCYayfwANJPoSdWeqL1lGJsxSsiQpS2iT9XenHwIoSPaRu0vhQnjAsM6kQoeDIpX6cIY5gfTNZ
frlvqTCmocE56VI7uq0RzVIt0UNv7Xq84bKrt93PvgqjlhCI47l8NrIhNs8g7voxYdBujqkJpt9F
QCpTwful457AlIoAk2P1M8TakFt+aGSx0TuIqwOQZkp7LGuGImLqlCFz4/+XkUmlbvCQwzSk8JnJ
yllEM6DJ8sTMNwJcnBRDBZmQjXyHIPuWpxd4hrK5MPH2ChjeUzwhvfdHxITXurZAv5RCsmQ7JfXq
iEhYyHaXXzc0eTUTc4gthWZbKWQbc4+xxYj5EKJaglpcp6birOyBwTPS4pnm6Xj7J+ZP5SW8476G
faQFV5py2KcYyiCKT9zEuo2CBF6fcFuJcXKzFzp3VIR5WTpa+1xr6zCZxwVrCAgHgosahiuPMloJ
z1YbqAlGC3zeKbGkrbQcJKIRT0Q/6lpD4LtBsSta9sqoKDzj9MMTqEeHJzhuvqJ5QUhw29iu00FX
1iW+cZeXiDA3bma9hbBIp4nSPRYMz5o2iwr9wgRrfVgZvmt2a6zAtTS/NsgOJE7zv8QJ65SFWsCi
GyNT89DkVgktotLrsIWoIDIn3DxneyxJ54hufpu07zEZ6K3x4n0tmFUBW2Y1dacLUQduwuZERMdF
VoI8IEidAIDfyc27+uD8E61G/8XuyXucNNxhJbCgfcG9ZE2lUxaLRKcdY+TFZn+Cyw2k/ona8Lz2
fGaqNqdNfo7sKH47fWaIMfBjUChGOb16G+CDVuLJ6rPxKnwEX2GjD4+H+jHoJzrEFoDA0/ezKGDw
v4bXdpLS1B8BiK5hacuZngs9ThTZ2cyXcZj5JmjfBEVTpHBEbce/A64+fHcIMUB6LB1TlJcEo8gq
ZlWAoIbATFBdR+LRdL24n/7fs/z3sWU2+P0LO9M3rHQ03d8oKkRgbgVKTzVS8m0XBKPIN3e/u0xu
yo4MCm7pCzKrG6KEMaczOTQK9XMK09kXKHU/POBcnlnlQCKBAPkn965Wlw3H8ZLxDpxoGmiCFVjF
DIakidBT9LCGvXvmYCO6lPFeT3jFBc18tF1YSPRbmP4FDItZmzTpC/uT6na7KHE7C+ro+WV9Wugp
EPMlY8eFUurwRTIk2Fk2eWrxdhmhim2IOTHewtRhsagjp+irXNzi8/YMbMFinl5y0+WHdZ7kJo20
34XAiOpjWmmbEiottMTpwPbYIq5TKOri90iJ8eZsvDByHE96le6ewqeuwhjHJ+9jzlmPg0A94Ofg
1Jsb91wroEYVwLS3g/nDHpJwlLWc8AWb/8da50/2eOCHbcFWaHQrLwuIXwbZwGu+hJGRhWiKBa+O
7GGU0OgbbIHlelc2LweXhzFbTOOBuJ8dkpnKAK8C0nkGe2ENmNJZS0FbICB+CF2pMxzaG9lnArho
cINQDiLpfRa+GQKNdEEl//WUtiS2U/SjOz4LT+bNNB01splxor6gOTyIZrx+/aWaH7SNhqg3Q1Lr
jO/QVnfQWAxkYl14G08sDKzmlz/CFicjWO7TeFgTx0uT7c6fkz0pOPh0zJYqF3btYL00OqOnGEGy
NgOlCZZtdUPyfFU6oQJ19H2CRN6mScdeqsaoCQt9igTjtpxclvN5RqHmozQEpZK0IoFaeZTernIV
J2DmwuCzGRKerF6Yml4961UvrX2teyUMmVQJz5dzVsgl6PNs1R8e7tVqlxapxzA1YLXk7+1dHcxf
picKwIHeq66qV7c+xqHh+2qUm/H3NWujUe5r51P/QBwkHINbJmgaQrRo9vc6FCyO0EbSGWDf72Y/
SYGdivLuW9fpkEFCxjozpKnn0qdP1EllWk8yM7hW4UoF4D6kfLwWR5CEgV2/gShy7kmaUXVTlsgP
xUANaDu86xu41y/qMU3/3JoxSI3lJ2sCpX4Vi1aceD8derZu67eZodIZ53z5cAXGyojK3bG1rHKn
UvzlZsvkIeBw6cWNiMrwngiNNjrZeU6/smiXilbWV408g8J8XrNcrm4ZPJPZ3lIZzIJC12FcMgVv
f5EWh547maSNy8lzd6wLvIc+9Bzz8xcvpTYzfvh5A7qbgTnSl571W5OUjcDejh1E4K3GwgidGEOb
MVunsVRgZsHnKtwwPdycHSIWpthwAI+yu0esrMXgVTAEhjzwmh6gyqWIu9/sAYWVNOnstoIhxQsO
1IdYyfCj2qRBxOEGKK3OvEwBoHgELgIONQHusOqjsonqqjc/K0r3rMvKlKdvBVwxuESOmuR1Kg8f
fQUqkAAyq3ii7iwTAUmSK3BUufjsWUr8iWrn1WruM9VLQaVneHJee4lYIrJ/P8CS76L1cZNWUijl
QIHynKG05pP1iKE0dnIHrJHtBHYpum2VsCkSo4ww6caGckOQ9YRa6DPe5k5NpOOoRTekKVc0bCsV
6caEyB4pLTQWxkzmry2Zz9KR6MzRAYT7LUYKjagHJS/ULtaSImvd1CnRzEnmkbl40lbIAoIGN70X
axVhw9wUUuFf4/skUiLXX7OcCg9ZiElRzJ90to+S0KvHmiD0uNwIgPVbAmGcvLac5WSc88zbGTkS
0m3a82pLtFazzvQoFgdwXglEvKCDfUmU4+kOAd/2T0svx7RMmLuEcxlCcnJolvxBmPBAo595Vr3M
58N76NXNUN8m9Y5fOBspVfcxNriMG5rmr0fF6U202yi2qbObwHEcf0Tu1EfSrTfZff+xLZ3kwZL+
JYCq2ggLSKZ0y7l65lDmw4hlUW9sh+GTo0AHn8gpv8nTBHO9wt2MlYo4obHimMOVNagNj6Rw+/gn
bnDi2z/qnfxB+BidEZNGSZF7YP2B/8BOR7oY6JKD3owntHloTJFNwLw+NmMklnnJk8avMrqtJ9Wz
n7tafHyMrqoKw/ZcXDGtszuJt+tJLJJE49SrWz4FqYqsDmdX9YJdaq6bdCvPF2HHUMjlwu2mWksD
2TFk20vOA/DYcZaJIHo2idNQgEtIpNeqd7vmWv6CouxiZwshDQMaR2A+1ASbx+ggIvmW+9iU0gyr
QTdeOZun1Yg5+kH7OfL80geQuBQJ2k4FRmnx4Hcy7thC+b5eO1g4hPNYEW1wpWg3FTKAbvpIt1C+
JmhYQtk495nYvEwjJOTnjDHgc7By19wS33f4w57hGXUPsIAQKBUHpvXMzj9u7mdkU7NXr0EZubE8
HFAxrhPprF+H0n1HITyg0nbvruC8QqALyde/g6wtVOAI2gBKyAdnSMDVap2lXUZDoY9Rgz3deGNe
t8FunhXajoLGmUuLsMMjTgDd/YZBZxkHZ+trwqYENVVVzGxP7KNR+DX/qAGzddyDDxrAS4KFYm1L
TEQR5/5GejhIpj1ju74f6+3v/Upa/TgDbJN1+xl1yM76SrgyAnozBnMNjOUAu+ERRX58WV3S/XoB
NDJplTQUKUflmJtJJlDed6ZpNJ+YGnFN+QvdBqvPDw2ywvYv+mjueklOyVUcuf8TU1JZTWr/XXyg
7Br4GYixFMf2n0b7T9oAqZC5jwagLPen4Jy+vXK8K7T/WEV1/l5xFsNHKriK7x8twAfuH83byFUi
knUkpdgc0JZg6MH+bE5Uz8WuHRcD5AqlhXgq6fyTBMYCuTxrlEMxhYa5aPVLptk4asd2CX6DaYu+
8CXQfkVudv75CdgH7l0iEtg9GenjfdprW9Vttvj5k9UV2e2i+LAdRPESh6xG4SD6K1g30Hh17FMP
rOiVBtvpFpbAwt6gnOl3aUDb4bMmADDDadzSt2MPQDQKY/VbGOz5hfEojlaXTrDOv0YglHo4qUkT
9OTIOqEmFYxT97WmwR2XstmdPMF9VC4jWq2IygkWO4hIK0HjuQpE01KOGGaa6LiWpqFWJk+LtbpG
UI74vDDjrX5sHghJl+FwA/ubMTKqNy9HVXbx/WFtDPHM5Dnq7av3eW1YXGG6cJK2pLELzmgdJkgr
OcPJ1JAqqvtxW8OHM1tYPitOhVWIrUnMFq2Ocq3uqhTdngUrRPtwGhNPtU/Gzg3w/kDz3KTYqS1Z
G7jWNYm7sEy9OQVA85LZDQqPgCfmFKwJ2sgGEWl1aciV0OI5pU1NVvzwvPpU7qutsvsYxrEiBAw+
mYmm7wBCDOT8ZPuEGU93LPMSz3U8oL56tPSWg8criqG9Jk7Yu1kEG9tGW9F6I//FNYSb3o/TFlK6
O85DmE5l7640ItpPYAkc+opBfD5c5EGUOTpDsHutwDzu9N5KpsWc3Tx4aPCwlYepsUohJPKyNyUO
FUHu9/JU665Zb/UEpTGYdXQN6WPA0eyBn4qwpZODK8KRA+kBBB7nCnXQBDQZ6dAVUmJC9CNSR+Ko
loX9rTWWxORYny6S/Xqupc11C6XrfF2KvD1hVAn12Pt1gYk9EwbanxkxmHiTegIiuodAFkiwObrb
fgmvD15S9mRZuUh6aFfWxMjMenBHVXICh8SPJpFlGs616wmI0EyKReY0z9bWFM7+hV+wGE4yRA8J
e7kKXSeDozuIkQwAI3q2Qr9w37tHcili9jsCm/NnPd9bXta+p5eslgoV8fpGabGelEr5UbhXBobn
La18c4DdChcKV8FixJvOhQB5hh44RUGvXFtOHFTEQUsljwatFJVDQwC6ib4QRVXHoTjGfWLVmJJG
ZCLNqb5QePJZy3bSxq2n7BVDJ856GVMgFxtsjaT87ydgkVdcY8SGwXrBf6jzXJarVVddJd60O8ZV
/44o/r98SQKCbHxZk+dyMACNQelig9YvHOfprXPqcMsIMbGlKZYyCw/6sVp7oVH79CBWOHCKfOfN
601oNdhMtbUnZMpt9yLTaiwZHb15XkpEfrdc3BR2jTYGxP5DPo+i24lNR2C5dLy4qbia8uw1kcE5
9Hc+b1+lofTMtlCGSIV5FDODHLdqXwYNEopUlJVkW/FvrKdzQ3ElOq8zsjbD8j3J4JNfigKR5JKe
dmwUCGFN1Xewl/HI4q/Pu0+t2YA45CXpkLIPIBjx29Ax+4T/ZVBIim2viN3oUG5p+BLBgqMGYu3N
YEM2QjVojFvja+K59ZwEg7/6tvGn1bYBND0kb4M4WsCs9O0rhW5YwcAWj6GhcHa2cJuvSiDGYR5K
F5JDBzfnSgsnx3kdaOipa8LVyDixqzbWzciNyYNHRiZM+Rqo9Rg9YD4e0UcfissZyLEA3UYiBahv
shMzdVrErltroeef4pOzbuIoI5hmlC3yvPb8SNNs+pMadn13LiJFUgvsK2JWEIVvEBWvpdoiOJiY
iaHYytlz0g9l67C02lXnC3SMVbhX/WWzFAhrJHbPTrkLemtZmVshlFAYjHAFBl6raWN4rpukEdCx
TDKATKkvqUSwbTwVA9oX4lTO9tPoTY3lBr1PEKfo+LhsGKD55cbWjZBu+B4++ACU9QzCH6d4use/
WP3iJruKuC8SxHAOWIACQcWwMN9sgxTcIH/Qz6yXb6KofYRAwoYqQFrjBJibv3G22H2muhI64sLC
5KZwVxI6C8QzRqtlQvNiWy3R/2cDbTbRhoNl+zBUhgNYhBlauxpLUEHg1sT1GcyeBAImSaljYJKR
W8d3QiF2YJe+5VfwkVCm/G7/cBmoM6dbvq4GqVAt+vvL/gqnfsDZRKqa86p0pzCIju9eiNjXKoCj
sTdb5yWCIyAeCb43POEEDOV5tvhqdHokOLOPAgbSRVe0Wyn+D8xkOfjvnGe90CzhKDwY3pOLdenH
xqwrD8G+bDeRM4YCCXyds6Dvl5m4Q7a3lfimJqCU+u2JZkV73oqLdUikmZ/ORWvukfG3MYPYchfM
RXWxIt45taBl4j97NKF55WAnQsHAVpol0LSff59Xh47kgo3jQdn9OBJuaH9TYlmEy2GWQ5QFxjFa
pWHOEj5EpSj0PRXxFQJ11XttPyhgcPUUW2/wDROePeTsAWpIYepnZQOWZIDWB7rJuSDbHQ0DD8WI
qF1qmB6QPuNhYBNZFzZv1acwMkVt3qNmlHAUfjstoK3c3d6C+ML/MHq6K4FUEiMhXXZSbPifRcI8
ZfT3WCsEyt0mPTyLLOQHG9h6PIGhfiLTI4qOmLbSFCLo535jGYmUfvKIsdGRpJUzF3UBSmeD+8bJ
VhWmlZCZYCW2jqCRDQrDKDCPnoSz/PQMLayKgzC/0h9fAatZgXWbv6MuCoucSUuLN2F0PG+CfK2k
OxQQjKbwGv6LVGnbPj9r90zu/9UT9CQXl7GSYKpJbBjuzS95H5Ydhx9WWYO3ucirPdv+Y3XO/0kE
zqZ5+VYzKP8SMGW+Y63uFwAohTCI+SctSNWepWqSIED7dlDZhNp22oZkz43ooSMuxTVkb45yFdNL
r4eV80od/95YAn0SshWfjrOMI0bxASfrH5yctw9cgrOo2UsSCMbujJXaLwz3e/hrRNGZCPffAgER
GtTVGGTDbd2w6JJJog94/CvAfgJg/wngPq1xPcngkr6Z4DstrHp+wyJcblCV3pTn5fSoGbBl+Zqj
7b7EXsgE2BG9M3OnHUkM4V41e/RYOsEMVB5pY7quZa9t+kmBGcKRnLn3Tz83ybY6yxTu7NhZNCNA
6h9U7HRwj4GyDEZgVCLS+kMpv7BVUBK14tmMuKbsXrY8e0oOuiFiaS3u5aNjn0/10Q5d3nQj39GM
PIQARTTyw+iGTXTRzNf/cxX3aum7TxxD1UBJsi7qKnX9bagB4aNAorKNh77dfsUK/3UK1TWxpraJ
Lf80/AhrpVsY9K/YpJYdrU/W0An/6jVQOT15BNdP2LDmkWCOmf2yGPa0324NbexA6hzcWPlNzPFM
mbyfKRsuJTIgS9eagMA5ZCVM635vx4FE8wa8njdaD+IiHsKjFKOcF9GoAlq9FTq+jOBMSkuTujYS
f1PCb4a1B0QQGuPQid45fgAKx+clmZ7goZZekYQT/glvevF32wuJq2TAmj70NRMTHj2VhHT4w5jM
eHEhDmAWxbHmouzH1Vb+FqubCUcio7cxLWk7KUc8oAXHZNw/F788RVRLKyyWU79TWLcUyNP2iX8T
G1zhoHNRPtNnHDEJfrsOlct/LLo2jSZzK/kwVDIBiUk9/T08vRtYgABFBaDf7pR9TBpmbEqLNur4
ZSKsVIpUQbsGXz8xxDyCNqERO3niTJUgn1Les44eyTBvUt2X+EwPdtzm3bjNiSEGxlduU/O0S7Zg
ulVwKvbfyl+HbrUqeoDiZnCme5zRfFEQFnkPrZ4Pxt0Og1WrefG6kvA8KIug6o7/6noU2Q7Xrk/a
tr6q+Q9/j4gF/BVqMQpULNOlb1RkDjwsWn1XR/ACyoDRVHxMO1Uyu6URtfCBJiKNa0ohX+WzC22G
QJFhM+HdGm6lA7CstAYEwKBGj47/tw+7goYi23Ob6lnhvND4VZd6IuXJwiMJkePrtPiCfEo7Y0gY
VozuRkiNlEwpY2lZ+oWgoYWSEYeMiqq8noWqVGwSzz31rN57RG8cniHpSWv6lgKLhpbk8cBU1QBy
ddFUEgX5CgCkCYTVCbFOc4nwvXj7Siabgqop0C7cjZ2BhSgRFnr3DZTl0qkekc/5Mr3jBlClzXgd
IwluTq8eP/pOkDewWKhZIMu6VQEypPZRc3fwTbIZP/OCTU9qynmRi3W+Er9VcbiJb5WFk78JoG2H
zajn/JseR1cPBRZHIhcHz0mESUufrvXP6EbfoaLzTnzuQIx1JDq9jSRmSuI3VabLjQQLxrlQf0vr
Rhn0hHPtwG2e4NxdaXrbYrCNlmLyw2pe0ql3evIca7Ec+COBsXiDGMb8LK6qU/BnsH0vIksrxwf9
yD7BVuNOv7s3IQ4hqpnaZjy9yJL9ovC+v8O+EZcnvIMT8l75eQLIYqOffix9CsM8zMMfQMvg3Jsl
eNNt4LnUcVqN4NUKgrSmBuo3ec+CrfI7FcMIFm+W08e/K0xc8l1oIcR6u5wnlChLUOHQ73mN1c2q
ZHdQELsxgDYLB4hd1yU0dSrl5I/SuSg7nzRVtOWZMLQRAjRfkOy0tQOJ0jDX8EpmmX/AaD7FVxSg
ZQxCDbu0YMn4JFcQNsiJ8SxCQXUcX2zbwZltbPzEwJtsd1yCt03CebMOOkKmX3tzGgpvXJqddZEM
3ZvS/so8HSRlg0YgZYraaxBWY5sJwp7aTLNnaPftX92mmWb2fxpNPq+NL0H2Qif90r8FGI6Mzcjn
VIfji5QJ2NtuKNu5VBhX2VD2Ul8DjVc6c5Lf8JyFDE93HfTOqjz5BNFczvMvOQRpwCkC62CmCd8t
fntOovldmbYKoWsNEwVg15j0Ij0fHUGZy0GMpyvjn6BgML8vXIbldH18o72Y0FAh1i1VGmCD6O8o
NdIPyRAieJE8FrpFk4At7wBk0dnzms5M5bderQgPa7pjRF6aMzgxuEY00EI6HbiHvF9BJ0u29LwE
9wB6NI8ZPYJEwj2vUR9LRC5vPUkVhtE9AHzcT6yggQLTUU/C9fzz00SAtenyQHSvy+PM57B28l29
+LbeRUdZxjSFz6BEsBoWibdgX5JcbPW0kNkDCioRZTUZ4YizYTKDF67AQqrdsva68+s0G0X6eo+G
NHjm3sv0m2jtqyHHXKRFqCE+QKlCb7TmjQ7W9e6w6v/O/WIivuArB9CCOwQDfw7SgfjXuabd2ohl
0P9dlJrGkp26vYzJx/14/UuKHr0NP9Cuewl1r+eRzeNcckK/ts3ZGuXRj44s6/es9Bnjk35n8nlw
+2ucY1O6tf1KoB+eX8lvgS+2TD7etnH78tx2r3+T4wyA+X1zz/eE5MoWHBoQzBhrhRfzum9ecCJi
2KoNGTf9QRClanYMqAkNal3se363tCX9CoMrNMYIMEBGzNqr6URRBjmjRoPMg9rGqD/ExOahjWOj
fRrhv6xXUMl4B1eb/tUZgci1Oe8tY3nx5BmWBkXMlvX5rCmy6ENwVAJROomGyj4fySvk2pLV9pwP
G1Q/H1LVxSDm1v79AZo/pCYi1BOapwBiP7m7tWmcMBX4RvOI3lQGF6e0rv9H8ZjIPVtKxLnc6YOA
s7a0d9S27fyUyopcpnG7zSXyLA0DNGhs/1PHdVa7Fe/ucwToLDAdhd9+nwDNyi02dpFBkz4YbhG5
EQFJW0SpNC3P+EB7l5OtvaXgPukjSR1GXZ8rN2T55bG9Lg914mue1vHMi1M0Zpg84jxj0R7Aw1eR
G+aAe4ZTC+Kaak9XwGKGDiUCFRNp35w2aYI8GICIqDNmSWTwf0OtJN2d2hjqUHf/kNN/FkHw8mDN
+1y/Q1xFc9XI3GK1NylIRNA21AAYDZdHBrmeYk/lnrnmCXPH79icMQ0vh48hSluzx5JVsak6W6yx
PtzXrEnWa2zx/l/iSz+7QSXRNJ32y/vHK84nOIWgC0Xso1rPw/u76wWidELj0JEsNgJ1oO5yrbNy
kFodLb/Jm/donopxK37OUuGp9XcSI+wEs0exZ4HA6gwPt208EBW6ag6sYOIW8N8th5HXM2hOsWVc
HBgG2gPCsDcLxt0pmo31k6iM3RcwzIShT9k5Yrh3YNUFQSkU/fwzOTUfY9ogqzRQGxuM6rpCpRdz
qLivQbZs2SiqkYo+Am6p/7fV7E6rY2mleEJLjDqvaQINomCQzP/mRSUw2lcvJ+sKseXVmmJnEm6a
mZdEaZljlmAuSnrd7qvveWFUss1JPh8bNNQhXyN1d5Go5ZbIxv17qBIR54yznPuVcXOClIGPMZnd
dN+WfNbYSwgX5QzvjariwFxpeQR8i+ZIgdQDiXfzwwCr8uZpDl43LkxSQRnXgbjObqlQWIQUhKgM
uzq2cMyEjEvkEdu2Lz8kea3+Bu3WNBRS+yMdJMCughvr0nqdKEK/xUeLHW+Y/axFZpNwuhvs1kjG
d3WwMIG5x+LiCe8j4ZdI1TYBYr7gk/mzT8iJo1eVJYRqTHBCuuJY1pIlpljXdpXNJ+I3n+v1RFfd
3f16yQ8ov68swT8bp1/0JYT3KkxTGW8Xwb4PyMDlW+auyoQ2EZIw0Ym1zORtsssQs2vU1S8pIWqn
7pckGQHgRVUB+4UvmZUYPFnAylqABpv7+U92cohQN9Gdf0EqtLbgMdBJpCsswveciBHGBBZiDqot
oU+y+tMI/AMz7BgzgVfKGNYmHHG3YkCkeiwy60rexOhcWlEHzhFK1jyaAn7bFtyuQ4ALUDfw1+DJ
kYguYzOHhpJud9vd2JfSMOCTR0OoPht0lKUpZGETvQo3BZ/n9Njew8uovblxE7AHXdldpUdHaNZN
9mfpPJZGvd8Tm+g+7EBD/vam3H4JCKMX6m1JWzhgKpXWutY4NCKea0yxxYlOZJx6DZuac4uFCKqc
gBM6uHkF3UuTeOg45/bMDbYuCFSIvN2Z/Z0JuXCf+CkrADt+19gyKdqDCbQr5L9scoUrwu+ZEhrX
3F/ZDzKv3IVvrUhfPNCXp42C9qjiLyGqLNeMBSztsZ2FEJdVGxQ8Zy/ayDhd3JZL6t1ijCHlCQUu
7Jd/UiofZaYKZnFOfu0oQl2lsxCEVZ9yifFpPPqLhmBeHkLFyQWT0xWiqIGXijPNM3j8ikaSCwE8
wQJzbLuycqrn/VfsqVVX4LUBNCiP9LKMnkTsqkt4l/K3wDavVgXKoRp4xDl0qx2TzUfHM+LtbuXo
ErQ25ABETt1QrskKgEWUANRwSuBlqNrzIqxg+jmA3hz2FCFccPI50c9dYMjMMPmPZNqsqRyJEzIK
+G53oAcZLOsGJpHEyNBhRl8JLf+g0PjKpqMrSEpBm8pbGJPmHiqiMtLnBtyQaI0OmkygcvkI56/f
ItujD9v45JK6ajm3N2oBoSgyFzdtJpiaxGFcN9tBnunyraIuSQTH47sNZVmg/L9fWop8v0savZcm
1qnzLRet3DY9BkpV11fF+YIvFnY5WA2Wlt99SOz+3jAzkd6j9KqGg5jXfzMJ4TAzPmgJLAaLduug
N9/IQeQtmR2LUK3pE/Dl32l1kFp4KLuxTkPq0ZWvesz8eyTLJCwHTCrY3BPlHkLpwMuoczMNdRXA
+LMrZc2IsVgG+GkJRjMybvLziKEHk0Snm99y2N29a7VyUCYEM62nj+/VVtLl+KreTULmmY9OVSSE
YSaQnWLoj96lRKTI76kjYhqQuJ/0JnAkY+mCn2THqoNepSVVQvJNydy1mSbbWmiV9FKWV3b/GdGg
X7eNnxwhonjnC6TQ4rv2rfdhGa8/NXSCqAA3rPxYnI97dalMHT+P/57yt9yVQg9EOlPOOFIizU/C
QIRDTSP8FDDpdpPBr9Qm9rpZ8q898/CaQiTbpx3KvBt1wNfUJXf2FRMJbteLX5Hbie7WR89qLG0W
/HvDkH/Jf0jWDtPLHuHMLoeMd6a0S9u2j4Rg82Y3+oFaKgpl4NG95fLt9LfVCWi5ReEO7Zvs3N8j
U8JMujZciyyDnQmNGwd7qEqk4DHfiNTM8/dR1ITT/G5YtE3HC3vPZK3BU2UlUW0azVtiq8py/fOv
zjf722uwk/+16OwMfma1j3XmPEzY738pBZAnINr82OBXZ7QifpQi7WiEp6Qrpfruzt5eOSGujaRs
jnQ6uHMR+99n6v6DslR3OZAysc2RlZnuV3Q3pSJqRVpqqcOQWzncccqZ+wbKA4wmQXmumIwYZC52
4DVMGxAsDhBBO/tpRrK+9X8pghxwybckCadDrs3RORyfYKJ0yLaF9MDJ16iRHuHcARM9Cl6LJVka
r+vmF2rgSPVD3WhaEPtQmIoNJ5zO8VNNfwO1v+NWMCHmD5tS5O799ZcrF8HLB29doCmc27B7d15g
Tur89m1bUfWWN9p4uvDNZ43nlOGSYnFyRDMsJ1UHExlPtnzKmL6c1w6NXyapT+NjS8lr4LzoVovl
lQNxKGl7I8YJslnmWc0xfsZFO3PjJGmbsAl1OUnwnKYpetwG+jGjPBm1CyOwmHcUE4gNYRE0K43v
zkmnzHAGSBkBL0hvxw75sME1ioqPzR7+h39U7g15iU1bppOF4rAve270Wl5WMu5Y7PQDQHwlL0dD
Sm77w5JzMyGd0PzXGMm5IY+YqADaK3TnNUQGTRJFPSuTKsyvt0N3acv8zipyLNh45scQKWm19123
3/EPUotW3q0vXERJ3HicaE/CRr0Q2+z+dmDqEl2dK8gCHNC8ad/PuuX+rFNf1V7eQe/9LAVFu/uq
M7Otc3EJ2PWmtPr+TsqvXmLhqEPlmQQupXdLLAdclCQit8pNAzEAt6WBHV7F7ceGAgSoGEc3L8ag
FKySlPJ05jAKSSS2KJ4ZVXQE76qCcIfGjP7CsZmKT0ew0U5vPPG//eER+719eUBxBA0S/i38YEpA
2E8h8zVOKKn4WxHzsEgMU+hVLr87ZZngvozLOsvEZOKZB/jMYhOK+6zt0o1Xp14Dghc678QUzNYW
1VUqys1+zU3inZR56A+ujytRKku74K9c23E0kzCNePMo8YeqjKjhtDUH8mOkinxxvV0/2ghrgPTg
mKfPJjGiGDYLfB34dBGHOEX74R0f825WWg/Fnsq0MsBXweW44AqSxQikvgblcKEOn2zbSkPecmQ8
UGN+F5kHBxWKVHVYhvpM71b/MbndDZagwdp+g/cVXwBCEPitQ+mPAt3QisubK8+U6a7ob0S8GjiB
h2SFMBBE8V7jMy5DuVHqMP+5hxabhRpYzfrZVbl1f/0eqy2JW99AQ37kFPEUDz+F4XKqV1TdBpvH
H38l6x2nbbxsnDGxZw2jJnMpwxAA8Q2mGOgp2tdcpxS/VilyeDmI0GR7CRtsAu65qP0rMXeWFNlA
A+klYk9LxSpkJmx91Wjqz8SRJIzw74U8GvyV3QQ7LpqGiLz4TW9EWIrVuW+P31DLcZxLKJ0dC3df
XQ/Y6n5yS399BEhd9Ae2POlEFHZS7E+GDrqNstfo2080fgFbKNiBH2+c2YULUH64dv/G5AAS/ujM
zuFhKhMzzxdqfh/MfM8zmwvI4rCZvhGqpcd8i0tPB64XKCj9z788WVa/vSc2Vp6UxYmHsU9DDNHR
JV6yBXeNjd59D5oVAP+jYXCgVeaBL3j4EypZ5IDcAfswU0/lZrxt9peW6ffia/1V8eDo2etB9wki
njoMmwuAR8h9l9EEKwCuJAblBgJRkkMnp3GbQQ9D/XZ7Re4nsdxi3YfvvGjN3qMwf6xd9UdILRXL
YsqeCa/Tx/sJ/foHiJzcUyse6ISRmyIYBvsRrPpASBdY7oSrlJDsClU1YdOzwrddsXHx0OE6W8q+
5hJ/5Z1ka+a6RuLQNF6B5sbml/fkRWo9y2AIIwpZoIlBpQkRM/UpIqhMfS2Q7ToKD4XjfDelhOW0
UZQAIkpppmLOL63Sm3pr8+imLZAnJ/5RzUH1fQhxH3luPTp+ciKhKqZxpPFyiXtzec2grmANXc1f
68itk52s5UlwG9kdk8L3QE2xmE4PCEXYNkaC92Bx/sLGIAQSiYyMgZ9U3/6RyM+Pa0XcN/i7kCKC
vt6OgbhHFjg/XH+XrMy8zhFF1/ilxddnPup56DWTc67RGFgiqf/9aHDiw/azDpGpbVI9PZz9EEl/
gwuCE/JG9owPm9gGRoc0PeSUjgIEQwxX4TNlrDjc3HsUKimYbCKvBh65bWtq7uN7diZxnYnSillD
N7/sT1og0i6gpe1I7zJwode0H2CxwWKr9o1xMDoAHadXzwBam0B8gExNIkIq95DbE8MdfDf57Xg3
FRb0rpbjbtsp1eOeiPXWpFxTbseJBooWHaATGKIpodiWxdAU3qls7CsEzSv6IRo9u55gtPA14HJI
7VXkuxLQGQhsEHlXvaGwCWjqXEO4ZhFASyznNYOIHyG+Hdkn3Hz3kxMryDW7af6CLFoPrenU/muf
mrJdQOnbd096aOK7K1mPJFDGO7kKVe9kdTODmwOSl/Nx6nD0F0P/tk2uI6XLLy/KkdvigBJ+tmOS
NRyi03DOguVrgWwtK0Qz7TzWWpCFYfnIDRwl3ypPy+b63+WjoyEZHZ7ZVkA/9WvhKbj0Hbq2PThc
A7uwCS0O4vQgRw7+5+HpbmA/LpY9RHMhQFcMMAsrsOdVo1SSddvodQff8xf0HSCBX0BqhYHRRlAA
9a5GOrwyoedMptBpAMOw4w/pzMBoxFDDpEjf8r0EZXR4ica9z2zD0caZXtFq0thtE1ZXVchiyCyv
j9lqaq1rdd9GEM6Ch1NxQ2oJpfSuLvzLL/Ev4Ml55XipJawAOe8adeAH//KJ9JXkm0Zj0Omk/KXP
2ViQP54hYQ/e+CmX2/jgVo5bS9RKDKChTihiIM2jqCZi/jqSFhstnNwTqh7eldWcNgRtVQVxFsPf
PO9hfUHV+GUQuL2jae5kONztnrnb9hp9ANu0xahit6p6aaP9lMFNZDBDornoRlLEc1m1FHPXvR5l
853n9iMD4sMQfvaYK8cRbg5Kc28TVX9B3fDv71JTdd7ywCkGkCsUrte4nLb6A1KGVi/iuGk5882n
colui3qAFzb3/rL+P58xJjsDFCsK1ZnsR47uC7/Tw12GNUmVkyBacCgujMEMKil7h4HsoOppwdPz
vUzfs16p6iieJh5xb6JNYsQ7Gn9Y9L3Eo5NImTNQxWfHIaWEpA+5FG9jW/P5r8VyKOJE5wDbzDyI
urepMpBrcTh4yDjiD0SlaaGKKhmbnF29Pc5khO6Bu328CfJPXBM52OcI1EJawnxg0Tvyrw95WnxI
IbpGeIrDdwk8SBWvAaypnB24KIABkoMsq59gYA9HA/+3DuzrppyzHP3IpJTWebm3mObNBEcLIq36
NEhQ5Z+KkcIDFPfgt0fizB5hv6JTSYNMZoB4hMYzsKk8cu5+v36IuadYO3+j2LEBXVefFij6o4Lg
4zA6MRdDcCWpj9ltonAeQB1ArjW8B7Cv0z4XnP6t/I2ZB2kmKTDnQc93tybiebvBf+Hfu/QUHsHB
GYn7FbieFBhRPps2hdiwvviWLIlIOwyev7KZ4jlzxwcsvL7ihXBh91HXha9XPeQv8jgWnUp8GOrf
ux9BQ2lBcjSnYuHY2VHOIsYF3M+bkyK7tjaWPYwahMlBv1Pmwn+oQQMcrWtfL603CGtbcAn/8VRc
GZBmA9BU6R1BFTL7d23Chx8eqWnuisG/s88lq6po5J46+1B0K/yx5hp6qtAYTSLISA4y5Nl3Hiv1
ApS5kFpIarYcmco7R/1pCpgBrwWa+j+QumU/Eehty71KP0+M9HynYG8Il76qe+mBRo1gvgh/DnkD
t9/Iuf/AoOQq9qDtevCgvRmmCbTMimv1QneVuZRkyfRAGJ6Nfc4ZLbNpWJYuPQ9tC5wnnmGNpJEF
GZRb6b/2Xqd+HwK5rYntbd+bI+bO/29C7spy0wEk0pH3zp8Okhg8K06onwekSxwaqc6WpUR0bq5X
hQi5hqzVx2XmzYQOg0KuoebgOUMERpSzBihFG/lONkpBfmxWeYaRfn5BLvdfhGmPsqLy1jzZnFBQ
h6v6oCrUsRmWWXls7wF2CdMS4PbNoPqcXj6Yn7GE/D0LvP35AM4V69cfBbLpdYrg1/SJNx1oAQj5
W807X7nXFXGYPCexNHWiLN10DScXaSQTQ3hXCUwLhlq6dmt3QRMhoSxThJKz8D8xZJHrSuRg/85j
SOA71Z/6DIwKAyB4Rz9Q9eFxxnbTWInFgGAF07nLkQ5XA9z+sxTB8syo/7YKXbpnuva0co/pdJvJ
ztPdtFsg0Mj73FAf4m6pCNg4WBk00Nlm3+bV4fAQaKGVz3ZOX11oqPmELK9IWvizcLfa/1jdHUfq
E/bbLgJ/yPoZDihuU+2sY5Xflm9oDbeGRjEUpa1wTc8sfC0aFKmFxs7GjcUL+LbhJnM9tSno+9tF
iVbRagUeHqRY/1zFherrblhw75/HCSXKjIe7eWT07mdItVJRDD73JQOReFtzyaAdCaDrhxWKc6Ye
1oDoTUt/+3yc8bTu8eRZnApJ5V7oYHoUuzfRq0jAlDwbwsdHcwA6fREx1uvdx6BiF1OFQjXF7UkE
D1yr9UrAtjQ4+4UwhlpAlhihpP7Z7IWWvKw6e3cmtsaoKnu8CPumklWiYW/K+t78LDeFY9Aw8YEe
YqBa9hWrbNejF8s8k4aG5x2cu87dNbhcjqgfrtCKy5XfG3xlwhpH+Wo7qrFgTF8wTpsKzzOHFfij
HMog8gMUB5IvPbO+LWfKBQbfsUh2LypJUM4sBK+esWd10heCreieMRs1t51eosYAugSUFb6EqbN4
AnTFz2ssJvID1tOjkztgdmV6HBQ2ixLdgSkRw2LTjCsYRdwmHGypa51ZW37VffqRUbBrf1jD3SBl
huS6hIp1Z1qQYWv4tIa1jWjdwqJ5OCc2o2WObwb2HMkAdCHCxkcVDXOxdkDKpDqu3E9JEWDDrIWO
M/y7ZAXhzEwrJmIP2Alp7MAlpsHIVwtmfPqLKq+Ho/dk2mMtXprgVcjOkyIUpc3sxlnEPk3Yl6o5
whU1zRz7u4NlTcMa63l+9eNlfBDuXWWsjrQMe8eDU0MzAZWGuFk6ydTW3zXCUbjgaHLfq02DAiWL
0bEq+lIAtR9JAsr1Kyz4ZBvZJh3WBQmCVW23KxcuMRGitFCCt//RdsLWyvflKcKgbos9yka96oYq
tmchE1LLNeFNPXceOAZfYDwrukmKC8OwNyFiuRNQyl24SF+BfrQlAkwGCEio40CrxThttUdMj2Tf
YbPWrIQUPrXHQHHbfp5kypzgV69XFtgNIgKdTNMRo70aSXWXXsApinBTx4ZQvL1kiVE1YqFK86QZ
oMHw/bBLCBkoS/YtWVF3jPHtEytXXUhzmqoGuYQBEyCS2XpHiOCw9X4n66QMmMdpAhBhl7xURfUA
VJmxMVmDqGJG5ZO2qeqlgfe+Zj1zm49/7RjN//dNdrc9AXVeWM9mCskqYgCOcO2cw9ylE4q7ZXar
5X4Gd4N832kKpON+eTXf5hFtLSMjaNompYD5Td9Yuz0l6cJ2oZTB+nLOa7Fm4bmcHX7KqFQkISl9
95ccbM1vqPxixOg2DFmp2MwwVGu0ae1ZaO5pojAKrplSNUz9j1raVVzKFFPexYTqeWJ/tO/jsaLq
b9nzRJ2chq01CDj0ioQB8fLK7mttxuIZJ89dPI11Gl/YG4DVjvzw8+wftPXMB9hXta/aRRCivvK3
5vUYmAOuXtAqAgMntP30kWikTvLGgNET7UypZzbnGtRc8/FQpcanEYX6b7jRs1adpxg0w4DvcEC0
weR7J3xTa2NDOBt5di8LltEO+b2RPaIK+svHZN+4HT1TsZ37tPjr95CKQL+3oxLWOBtdyOcG3dX9
WnPdhOKG6fzDxa50g4NSu5yXP3FVBSibRZfFcoUTtsDw7/8qWdKbcI/IBRDzc4JbIzWTsVEV9mfA
LYhzTILOZoFhzH4Yhhjp6sIEQAfQoH/bunuMkQnlq8VGe/hjzus4/J1ztFzZH98TxZgUuHFxxt+V
1tdzqqNvhHx1GIg1mPmumSCXd1OEKWQmBsu560i+/C/w3xT6v8eSEL+wGNUIuFhwOR3lJ7fVnKp7
BL84zwUiBLNIv2vVOJtNrDhSDB0FGO27JY0ixvHYkqKHHS0LgCl14adyGwey5xqIkeg0iblTHH4E
FpnHDvP15CSsfRLFaa4UF93YjNqhry+ZKamsa4dcEC7d6oDdosw0y/q4NZPz4RNbzViKcBp5nyBM
yOBFqDgAuusvJyZQ1vTGkp7JFcExiVYC7T/5H+sAyeNDzJQWViueGg3Ia6Reny8otJGipBVOSkW1
7GRPX+nn9L8cIsLQ/kp5PsY7aVRyKIHGtvHv45Mb+Et+njf9Nc9/fb61mxhFlp2vadzVUlOF4pgr
E0q+YmWWhpU6eVdYTdV6NlDZ0GWOJ+Qy1HhjcPdd/k2391+oP0Qf2aLh9fxcaZgZXLvLC3ojfsfg
tZF0IUUgL9sw+L25EQMk6xZQq0S0ZcGwakQ58LIGdDQ6X4Yx2APH97tttG1VE74+4aGI4PMoQlap
uRdT5Xsl0/NMLgo2ayPMfFSgvnAxai4u+lpUMC9zbfTTf1OpCyH/touyEeKNfnWhmj/NFo7nV4t5
SssBZuqDDHSQuRE3s6UoGsgN8GeWRdpWjSPgFMtMuBMegjkXxwY3DDoxVm1wMP4CHpRPdsogHlZB
sH6PPM/N8IAMwRCDE2jFti7yRT25elhgGfcLw5nkOaM3SZ/Nd7sTzBd13O7l65d19t4ayKmbtPVJ
cfVhuiGz9NG9pYN3VPMB+034X8LMyjyVb73jsNjQuyld+UdFQjZ3NAJSQ1MVi3MQKt0BGYYTwKlB
WNa35cOUNJ5Rj/pi6x7brQIS+Ik25+eW0pN5Bz0hMKRYR4n8U0zhrbGaXGdpCHTqqWGDvI3O7s2o
xNyPdTz9VJoPs3ZGSCNpghGJJM8Q9oTe1hVeWF5E4O5xwSOfq8FbvZKC/0Fruczh92c6p0jk0+PF
wI7A9RmSiaxWu4WpNm2F5zrJ/Wxe6ignWB/o390r5UKVOpDDWYC0/HRZ8YTAsHk5CWLs/RCOZs+R
LoTBwt51Bked6u3eVhan2SRqw4gadkm3s1uShVL0Oo9HWGsSwid32hJ/n+GKSYfVqxuEFMN25d62
WQB2mBB6oEmpfzEQGR09bmGjz4nIHe40sfwaTUcoG8GHsdbT1ovihRx5uzy+aZS71MB/gguNtNiV
q2oRbs8hCRGM713Sb5MtT01hjI5OP/Zl+vnWPaurJbo7IXinY21DqRS8TZzC3Ga7XBPGMZcCYW9H
cfjkmIDI5GGZ42gF3uC1S8hNyvrYMQWrqvhgw81QmEAG41VimTfV+ehe9rOJYJFaDX8qPIuYI1Ng
v6d3tNdUQxFQGnrp+HWu24TNc9z79ihdNHgBBMb1VPHeQOZtoXUDSaDaYa+bo6d5AZTX0XV7CB2W
FkyOAyQYPUnnt9UFfs3YNgw1FhPRXCYnUZcvKBajQZxaq8P5fuxZJ0NmmjPFA6snKcWAfMwPbS6a
qcTAGQohpFE2pwnaNucggN7qLjNrjV+xCR57mk/gZ97ykhqIKXFHhUvYpt0h95NWpWh6PaQt5Nlj
J3MH7i4h8ymKQN0AlqodSwq/05omfg2X9GgxvzOjJZkfA1ImQ0g0kyvL6SA0Nzk3c8vxHRCzWOsC
Wm6bWKtU670+Q5cAUdKn33YkW/G1vT7XsLbMIlhNEmuck4zJscPHZopxgqyd4K1UnVAV9y0ztb5R
4uPFrgNH27JGLHcRfyWNnM5njPAvlkhHIvFwxN1xyTYddoDN5vaNVGdqu/jUPH3LkKIhw8TeNSLO
2+uepyC4MaXfDX0UIx1lf6McDh4XrHZrVeRi090bvb8eFyokDId9/hFe7b3S8G2xGyU5svRJ8rjk
D49ksyLZzNQejdyYZyPVv1bKGBMe9GIYQRqGIVMNfL3n1wFFCnuNVCuHuji4IWJiJOc0NwGdvvPO
/h9atYKwcT3fpqbe+JthimeYJl9MHvJtl7Ivex89e5iDckZkR4V9nJ43eouEd5BINO/RLE/+v57v
ez4FAXriYrOPr6w6W1suzHmGXmCjoLeErjId/nIHA8tFHyscgC+RlbzcpgOHWjsL5Yeny7DSd8OD
D9u/PaJiSf5z2kpCINJjOcrc/bunkrgm5GsHchcTTCmzLJHMyIc4txKnTbTR1DJ9Zf6izBNWaJu0
Fi/SAPSAfRxb6Fi4fbHAIRxOJcfESp7jco5mvLGpWzwa/wcyv65cTS69zhsFKS35SL0iagPUwTeM
8QCa//MT9UVffMa0JR+cjnl6CMAc3FzvDyO+GnOfOIlqWacmYZ1/w1r8YQ3HnIG/5tJnnzrtcJmi
ERuhfFyrJslNWi5tNeluaqLjfi7yeeM6P10kTaOMSpI7gIeIuvT6g5RdvlO5wq9cwi12pznVY9fE
cqshBx63pJvOABAlLo68M+8wIc2l3muJbjq/OrKFbva6vFYGRmlUEWWcYpShibDz8Jayreo1Yp5P
t1pcwoOaId3fjxH/z7bt7RKBIc/+uN9SZcIhzrLBS1sc/PHf/ibz6pshWbkbw3XBk34MrERkTzh0
OUQXaWMrdEPxTv0jZDYtCNSqTpIW3+N93N0u6zb5oTViaBnAQKEKyZ1Qd+p3kAXIXSl0nAAQ/rXl
h+W5j4/7pe/6T1emML8gElRXZCDn9FIJytlideaMTomURla7LhOzmZrBWy5Zsm5wgVVEuOCgE/az
enlSN8/ryaU2SSgDH1MgTFlFtAUrk5D7s4r4mVhMr9MQdvqKkUEfjjPRCEocAbtGDIJYyIApWI7J
Ur48XVPKQDSNBTaKLX6IH//EJwHo0V38fzkgajavFMNbmODMbM/klN4KvQyZq5in/NmJqhKcsYbM
jlWfmD9vszgKBQqHJSNuAbGryQR1f63Lb9yDeeYCPvN+CAHgeomNxxsp9+SGjd2NesyS/yDUdnWi
8ZlllYVm15ikGlplmzOfz0QCdUYSNWgSAkFra7u9qF8wuOQqPSN8cv/9hi9kiApiMom2vquiLOOV
zbrXN6RVkEGUK8UkWje/0gcWOqVqOAAy2T5DEisAwFtzx84cNwwAJRm9vjCkcmHClTL6OKykWfP7
NXgaDzBWbly+HZhaGZgNnM9TxU775MMnHe46SssuNHceY1/7gaM0bkH/LuXeERvI7n4SSW8j9hsk
RHq+l6y1XwahFy50FbKY3EuTg6HmNhna6DBQzxIYHEEWgIwvFLMGo8NeLVC6+yejMK6GyY1MR5oM
XWka/yBPOLTHv4vBNeQBef55BqiZN9TGvTpDiJd4iP54qoRX/tpKW0KOQotxHA5tbwWOZkUxFAiE
IgqOIGAwxRdxlx4uTl2pYGev3Aa8CPMzu5GdXlOiJbJbzl/ctLtxbRAbB986G+PRt8BNo+CHmpHK
3EdUCNl1d1nNJNIjWLQWLk2KngqeEbZm/OzNxU93ikJQ4cH8b3MYLfUrY/HO1kCMa/wWRfp1wwFM
0durFbRjuFEPwYkL4HAWlPDy6Cz9J+ThdlAkTcICjl5MrVr4Chral+kN6wXpW2+GjYo407HHh+q1
QIYqx+pwAYJxwyf960ItxPQRtFaR5T/Y393xha/Wrf73t0FLW7vAh7mst10IsM83G9mJ9h2OA/HH
xLv2WFf5tHnlN730aYGAAUTK2qHUAvNlMH7sFrhVZJy8rh006zhrDgJMPxYD8seys7JbGaMZNTE1
OLq+19Mdf9KQv/B3ZfmbBRWYA5EdnJv9RGPH8J0Wx7v1LFCH4YbiVdhze9LR6SgfLaGyLDgV+MfW
dsaTKhumqjG7I6UBdMMMC/9APl6oQuFtwJ5J4+X2v+pyCSBXKiismTEJln07Wq3EnNBGO+P/JE4I
riU8r/sRqzCj6gCeMrZyJTZsBzQKYIXMyyop7z9FMe4gPwCbPCiCKcZhSxZDMZcs0ww+ogwmiksx
9KPYL1qrlQ8NNoxnSPFlMujhcJxs33T4Dxhc/xkyXNkQpNvDLWeFYfg0WuXNF5N/vtL/h2qEb3+I
2d7Xzp05z2gLdQF5yryYNHYNbX8Xjf82QiyUqOGlUrG67D3AjItkeCnx/qeuxLCQPsBRj97Do4HL
60b/0sN499RKE1KaG8C4FhnpOBEWfRZvGtRuQzL7KvXsMgfqwhn3PzB+GpsfUuyKJeEqiiiu8+V+
/PDE6I0Ezf2nt9a/6tR/xnFqC2mEJpq+Wo3cZx+xW/0ZfNFWuUEvPTriuoSAtmGnfSo8BM1H6PTu
c5h6u1Ec82JoXr0txlFYDtHN88eBwkBAHRoZ773sHxVwBrM+aJAaWBZyHm3Ln/cGVBgjmZ4z4D2j
EiLAvISceR/bU8mKzSK0TH9QwrS7kz4rRrdwx63+KgWV0MtMaB9YvLfWmMIG7Dxn2BKmOrDWlzTr
EaizmbSOekmV6Nw15nnb51EoKXwhJWdKiuRKNeZAZu59TKRXZF4noZEb4dH/pglwca1Ye0jHWuOv
73vi3PMUBohpnELH0s5ofPHNBgEW9Ltn/8IyEsSUw5vDhaza+0lU4db3Yz1R2GmpqC9YT0FQiqpp
JcWjjknl6HXCZYqaBpKtolWVLx4OCRIT8wD2phabNCVYdkvMNQlrpPKlvugx1Tky8fjDWiKvks31
e73fCicl8YN3eLMy5wcz1PMhL1oxV3UmIuU6G383LHnQw2Qz7sm4/T7rw1OMHq3j6FC/3YeEkygr
anAQGGmANqXUdsIG1Z0MABcLiqWAgBdeis8fmuIMr/rSMnJidFHMH7nYocqAMDx1j4ol8RTuHCM+
qINlHfRjDrjdPaaT28fIFJ41MYrvJkY4dAlgKVRZ+4yboSVwh55pvahDlznXluIfRe8cbMcA9TuX
J5RdFlb+KTA7h9S8FqSvR1knjCT09cuGhRSUjDK+LOocD8k5kGkJhnEtuwNYzKd8BMsWJp6IzYU2
qhyTlTqb2TQKK+4OHxeSTaRDY/eGnX7VxhpsymV/Hfi5v7X79BOVhamQpQ7OBX9nKD5XrWZnCy5v
cWxKKmdmMy4LHZ0WIUgHbYIt8p8Ijq/rFhTkfMOvJ8OiFioaWPMo6QuNQLHrd4Y6u7JOyY8n00Z+
Mhz5Hc5xIQk3FGu5Jw6YgftjRwSiZ0fbiCZdxM3JkI3pbj0bUvN6FYGIEExE1yY74WUW6NXL6kCI
GJ2DTMBMxROBOrnbZPUceag88ZqPgItEbUIQ7YnzsZLMdTtuHewrUctrJe9Om41+Anuo1T3a2a7/
qu7mxtYV2o3CgoTe1DlJ/SjRnSOVi+tedXex8sExwhYgjVQLsZT73omF+K7UYYsid9XkHEJpYCRH
oHEtnIvsGjjpZumZZXUEZ9Y8yPn5ZPLW6yTcpKan4pxgRutq6XhJRi9tNEX47HGKAGQh2uKMr2Z9
ORSZPx2xOJNrHXnJTZZ9tawjnl85b1fFHLuyQ+T+5zKlC3s9UQGrRSUu8OyoNpVLaIKUGW816Uwq
3pc179NxEEv1oXiqHVoKSWUSn7pO3vXRMH17W6/rVXZKxaPoWu5+HAH+YFMYFax9MjFlix7oRXbV
E/rVtb9w79u3+tIVJO/M56ohGathlGX4AeeZspDM4gMOdZzh5CFCL0VgfkOAJjb7Xo08MZgE/zTF
UT+0jBBCBblOhlXwKaqDa3aWs7Bfzzxc8SRl1qr+V2JxLlePyJq8KJAau/JMh8LBcMJ6xR91Twlp
9wfr32yFFKmMGp60I9BwoWa1kFLv1ISJw1ALs03DclycZX0WRs7aMWuNmRvTMChG+vrqIOmRi72o
znfPUnh+Eg0bgKi8SIzzyghOWwxqd9s+7Ks1m8TceIt21j5CzWh8P18lc3kQROrEEq3EYKgZ/LDw
N/F5VtG+481jdKPfnJAIltjxaTk3VzomIVsj1tXGOvm38vSDlpk/Ju11lNBlTlQX11ZOBHdGREtq
WetW51nslw1GD8K2xOghEB2bBPOqQNkj9WJy6UeDaLyeyV70l6bwUT2N1MSK5fHRiNxsK9tjgjJ0
8s56Vn+WExc+fFMA8zSY/wls/l1yEEtShQF2CqBF6/x+gC3soZEFczXU2gQ77y/qmvTwWJjvKyfr
bReIe41N5W5KXMnFXxD60znl1s2ASIUpuCvTwuuxi+xAH259qeSUDTh88YTeqF3dnayppXVdqMVZ
T4aWJk07o45QMhbyY7TjZoG0xvSkygUyHlyhTUSSJsZ9afzsA7dRwwjw5yJmW2MksxpXHzm1vAga
b/sUaJpJ4mMJuzv1MpDFZCmlaKkQbCXNB5wouCLGaHP/Mqbt6rqAgu5mDJTsauQHh/vU663rMBgS
lTdkZ2MELiaFQ0aXcrVtynik2IFOMOAvRptp1ciS8UL90+zU3aUSujB6C8E23exK+BWHrkKT8345
QodncJV2E03Hq8YJ9yuUgD1c5uKR0kE1m95BEXFgGqaIWT1IQu1/YagBI3jXOo+9ePj8CRjynX6X
yf48mIuA4af4zwvGDrg+37FCmvRCNFnVcv+b/oFEcc8H0Jv+xVq3jXQZL30wIrYUvFRVevEYz3AA
FFtd4/dPwcukGq7hL2qrA9kfxDCVpDwPD4lq+0wrjI+Wnqp7SxfrCma63HHUSeSBJe0H1z+h1zrn
OPo16qgVLQ4A3yN/YVlgwKudDujCz4mBCT+dIeMb2AfMTnbbaTMQg3qA7zxFyvln3n3yXERp4QWg
b2dm1kECSmdkex2uvQN9fpTe2MLfRrNNvK69f/3y2xZ+o/FfHgyGj2y6oAuYC6LqxIzPobBkInZb
ErRJjrTF+w57Ob5Y0szwJqHKvUmYZryooV7vp47oii9t0CMMRkDBvkrXQjmDLYKsOYmPbMcQDT6u
2b/TfU887+8W6FhmNvarhfgxNMd8fkM5yaKDvgbk4Z5XFTyHzgO850sh+C8Fla3EfU9dS+PTVWGp
0sz5YuCim/aVOwNmc35srrN842M6wZ4/Ypy6wBjRNjRlflWqoYZHALsdTYct+xMmh1v05fvdlANU
IlVjFYGxiVYBSlt5mLMkKfW1s6dKIYTAYTU0ar+EfQiYT66Jmq++H5KIUbX+/qrEn6Cy/O58oJxG
TWDLyUJz9YjbUZVDpYbu4EU1viD7LPorc+vwVjYlmLb4mtPm9cmwZ7XDxwABmsu3lezW5dZd7p2w
H8yZjdnZ/KP0HvAI5IKwA0MnQfQopHHNb8hUhZVEA5de1VkTrCMxevHnpJ7kB3ND8LYxQRaib10G
HI4f0rzAlPhcCCaGpNI/Elt005NOQEbatGaWQXFeb6lGA3O5d9upp/6ggKkpFdkx3fmSfMBAHF70
tRlJCvJywt5qvGcEKW7hBCfzPFz2YHqZE5Av87UMm1f7NFnJbAFnETaWrx6scxq6irgQWrRHUoKA
XeNRyp2kNRx8w+l1wiHXAnIWmhKDa7nWUcllFwgzFLUeaQFWSGD6vFOj6AmnK1y8gdpUotX0+p1M
2m4bvvwQJgjR4eOcFopJQk1ULyLYn9no433pfRwr+mxniguJOKA/QJ46AUnS/+0oONKvg4TC4ZS/
qxqL+cpzsC7Zklap+GV4XpFCJ+XkYu5N9dpfmoGXDYRX6batj91EX1od/kqcXC2XG1EIlI0uG5xV
PU82niVCwCLxklfVK8Yv8lIU5qDX8CaFuX0iMEYOOGOwKXS0FpxoAKTqq3m9+tHZiFJY5TT7dIO0
15TWSU5bqD8jKf8tWxoqyK9WiYDevKNtWqr3+h2O3GiZqYMCCFIT75MqvPHznlDdly7wYsoPpPe8
cJFsbYfWnqxK6WLjWD72T7bTZRLZVMsJNV/4zkIWEMwXBpiyuKvLdBe0j8trvQW4ZjCoFyssKTCS
IxjqCpJAPdBsl2IavK/ABPHeuUrckTC2wqZxHjS0F3dZZ63huFAeA+2eNQWtZRagukgiSggRxYn7
mVhpFBEFYkGuKsG+wRJRdtZcyK1MydABj1ejErjZ/YeDAzhJNK6p738W0YFnvO39Pqp8g4ombfDB
zENRQMOgalycoNLO5BfYyLu7DgS2+SPE0JCyKXCvjWDHk1O+tvl5E9UT1+mBoLXyNxHkd361Hvyf
TrhEqVmM0eXw/FgI6GdU2fBe2OJwtNAtU8BK4rP6tT5cTkjna8vV/V6OL0KN21eV5L+lEUMr2008
sasmR5gT6HVfq7ImIOrC6DHYNvCxzJSlZEw4u7+XFM599D2qPHEQLfAk1v4yzCLsQ0e35JJCkFgY
pgDJrIfNWqwP37CsvBwsMHgEz5PrRyLhos+7vRZob6au2VpeHIOSHI6b0TE24Tsr96Ouukj+WMOH
qEdviMhto04+yYYZMeGUzRR+sCbjbQt7aL8YuwQJBrRNKTVfDaVjTc1YnazPuiZ91m71PFEGrbQp
YDkZGtdKUCVX7J7bxPJNNAiRstvRloPEvuiUr2kcNUo3lY4Ennnv4X9oboTOz/wUeSBSvRLbpNU2
PyKmNkk5ybJPPtpJTiCX1R85iglgMRoN9lghle0JHAK15R6bOFZOTSzNPMVjlhrX1YAv/6DxECT9
u6Uh65PfO81g2JMJBSW+VgLHxjFyOBjcSE92akvZrbTgjNOKzjqGzQ6ISRBGR3L4P/I4OvcySsxL
0zusJ15/32MMeWuEZ6Sc+8tERyIG30ZYKl7SsLGnhORHY0tJNMiXlVgYWwQx7vhnNqjYIhHUbJFD
LkzJclqSSPFYHlM4llY4vK8H3J96DLPLFAi8XU04Y0bRB0GnG9edhW7DwjDRkAjBlg/TkT3JgmdE
V3c2shItNENSvWPShIenn8+34bKs8gHYp3Z0PDVDDXA0cvYb5/lt4rwho8VsbQRITWWWv+7hdpuU
G4JZOTtOpLjBmB1RfHH0ZmXDs0aDJsuN85O26CP16rwwzYyrZCbIochPkKjaCYvp0LR6usv8v3/K
nUdBceIoUgRV6QFUvJJgADH8dvLf/uOYiaa59hmAY3Tfe73G831OSLcLgZG2iuvBdr/t9oDV/hQY
CHHXTOVwz1hU6f+n076j0/f7bHmqF/mJSxGBp0bkyoYR3gsBZqlkU13OkCvZ8ZFjRY5lRT/A7WwX
YCNrpAKwym3nhDvaA16TnFwkHjEH8fBoIFfnwPTz1iHZ1O5hZESa5CBKX12bDecL12mZT6M8jRtS
K/aANHyYU9YjjB8wQIVqLAmbNVoaZw1CnesvXb9g1hb/yftT2zsVQPy2862b1TMeT6hRBNQc+rdb
Gl617OHYwIMHQPdn1ytSJBsSBaTMdkoMCq8/mo7RhRde7unBOoBxIqAKk++aL2428UGiEuIMKjzw
EEQ2YTvkwfJdk9cSbo6PV94Vmlf2ecbIzHeQCM3mSuA+tU6YloteyzgFZQgHhUIUXYXsPsdgS54a
VJNTIfMlUSWPLZrTraXy1kWZi5pwTFgfWYcS10RCgegVITizUrdsNAM7IlHH29d2SglnCekQIozu
xFwSK5S6+ZplBGXudHdyH+maWg5sjkLy2kKmEWX5fZQiX5Po62mo+TMqZNGQhTuWbcfTlIElwQyk
KRWNxwJL3njtq+YSr1H8vCHt5fZBEArEimD9QT3hrUtYzTozF5BL5kip9av9qncRNbXX8F3cQMeF
mrXhndGucUGNSw5saAeJHuUNC1ilbfszZOw35Uv7jAls5zb9ZkDCxZBuDb3f9/nu9a/IRoYDSxlS
05H8Usba2SuLcEKjdrwikuJ7VMJ6oVSnbddtWMukS/tG/fecArkep1eFuf48y5NKbKrsPDeIwmLw
ktM2ka0zxYEfpUXljNOCbrO/12QjoMhf1IrAfYQ3KHmKPgBwO9DPKlVY+v+ECRuUeqNtx3CAZck4
cJ6GWDx3T9jBK4/5yszVhzUNqhZDy9tA77ckOrvk8LzHRryHyBCdKrvWpFaJ6jxHqaoq3cz2hTSb
T7arx8PqW+3Al4cJda+zc2d0qzgcv0u/rdxoPLHoq0f6WWEwIhQF/JUjSnQborzJ6j+jgQ3W5bmG
NHC4icnSw7277J5dzxLEc65STszWvOeZfT4FjCk1VeYFpv+JMysSvBYfB55DFQWqlP3febWxFmPU
T6jHZIVK1Fr9rjh3zMeLenEHJes9QL7Wwy/y8rSRdMw64i+Tcnx9DxBPVrGqt8zuNC2uXmsEQ4G3
hAGXXJEJFmwji3hzDy+czxYX2KPGta4YT+B/Xgvbb0l75E2OSbQKyg3LjMiQz6fu9k+4LwK/0QB0
F0/meDsJgjcYzsmxT2gkG0UYsNfhVH2opcz+lJS4eAFKTlQeEW8c/zE8BpQhhTmRAnkF8Qz5NKvN
Qw3KPADlyTFRyRl4E44NzezANzl3YnOXCoGLHdJcpGhsicf/4FZiOAeFCfKZMuG4vPd9f5RrNi3x
wskNXerMZbg3Pwk/PGnuBM60t4X1pxnrU1dPNkijWlUaYrsi0kIyLCmolKMG4KbtrZ7MDUFCZFqX
Q7/q7Ja1EgsCyY/kYZFPL8zfJ51j9xcq5tQ45TbdIz6UD5Xey82thOs2KQSTByyxpDAWHJFgaXUZ
Z0TrcwWweiYRmFcd/007/InsjL9Mzf8zmLabw6vIR/rpxSPhgt8qu+2Z520mexGAH9s5EdEWfwLT
6vaIWp66JzKeX1piriDAluGMjnoHciaJ5Pn4DokL50k/hkKC/bOd5wzq+vDttQb+iTXUcp0CNHXl
uqys0mwJAuyIIsn2znpeMtOy13SY1NmycyPVrrLpuV0Vc+T/Sm7bh+2v54AWuwFWqLubPletQjB7
P4qcqkxMmTjSqELbwohvg6rxHcWOI5DgFSc22pSI309WGyv11yOZRJt4818F1CSM3kc1HvDYTorE
xCpdJC/yAJbAFq0IqREMsLpaZ6iR6OUdqFMim4Td9G/LEQ9Q7lnHvywYC1mTfUevtL1UuqcsAkNt
Uzk0tRG8uhCQdQoy9SXvkxYBIfjjpzJ5kH7v3cXGkl4tecm4NmQD6PNRczPSeRwoeBVVAlfDHB+9
Kbj3I0/rzc8kUs+L6qM0NpwoH/daxBM2qEkZphC7An7fZheWsdX1AXth80cA1vs4lp09VjtbVnOE
qC5AssarDv8Zbia2ezRT8KPrFSQoSkEHPDAQ4av31nDzke/9zabpTbmPvgnEeFuK5P1/y+nA6QEb
5n/SSOoTRQE6xqUWfvyQCb88QcMRc3BtwCrB/KDqpUq3xiEO5N0QKXr7QsyEBuoG0MP2VqOYq2JY
dNIbFk3AodKofD5MsbADg/vNSeAd7Y93QIew8d22bum1nAtp9q6yywApPwZt5Ftq+mlywrfFWb0P
rKPOEOxxfC54346bqE/Lec/acTbM17c92kI/c7j3hhjijfSsz7jJPdnEOyhmZG9k8KH958/Ab+te
erweFY+g2anHBd/+rLkTQgh04fsuuQGl0ItghZY+b75veNrvSLD5YrXuxoShyzL0qJaWSgZPy6wA
AlJ+6wVYwicLV7QrxS2VswgvLk7vkUa0ARvkBvlmwU7cb7ctwRM2yvhTOpk95rA+biVOO2jzfuA1
Cf21eTfRWhmC0NHeI8ow3bzgZXMI92zr2ET6RnhZ4BBDgopCKQYUiCxbvSpb2bMRuldK9dcNhRLa
fdhK5WjE1nv9n/hEOHUIRYIWabWoBf8snjtXl8PzPpdL1Ieb2LKad6Oy5pd2+kdsyaCql/mXs8Ij
JxqfpuxV8GoVKQr795szog2QYfoYC2IV7Zbven/y630gNBB+BuQvCpMApjH1l7A3Jp16XI+BRLX2
GrS2WBDAsEGAMEW0WnIptN3DINiXlrEuSQpZQnGEyAlpbAI9xpjcezpFIYbH8iATjF1PHqaWoWGm
sgW25YVFsRDUxESMCmcP7t/mnfRODRR99/5nPdGg8M/EEgritsvdtmguwV3z1HvjkVv9ry/F9dAK
NS6/9IiUtUJzPZcH9YEZVRJ1Lv3fY0oLSPKDwILIVUZhVcXVQU9iJRVc/QyCzuG6sozOYBBjTLoG
Pt0UPluNVihIrk7wHsW4y/aTNlMwAIyJWEnNcFyftMyX+/7IyEof3zzYb72/KMtiMm/lAxOG9xAh
aEAvQTJGuC4UIOVS/Lj6TaZCcOriquWLLQV4KRWF2bx4MGWVbu60pzoG+7EDbIZ/MRGafH9vZBks
PMP8rFhd0VFEP4XHyJPYIdPaXYTuiKyit7J+04yN6WMpQYnVkFbvwQDD4AhnfjXcEy6ZNbU48v/K
J3pM+zZmydAbkDu4Xec1geeaDON4mkEjtyAH5FpjsIiI8rs999L9rF082B/hx+IfybutXnA9DEzh
eG2AmeqGZ3+PXnAZ0F6sDfh1ntl/RE04wp+v6awFHS5fa1AnSxb3IxQYbwInq4r8gGmZth79yMQM
qgBrB9nWqCGwVQiL7V++HU2LVIfvzxcMh73rlLaiR/FDQe46QWB5ywduOptWv3cnGFMQ2uV8T4MH
VPIv7TJDpc4pKRFioKmBjLEFXr00xMIoYhwPloPTda5sESUoILYRtboQIDyitm8a10sucnoUvkDi
L4MkYdVbG6CGgw/8DvWdf3xNEVuZW/h4JNbD/+DyUt9T2SAG72L+iom2iOfdTUNSuPXv4Y3DlVOs
aBHIlVFm+hQtabf27PrnreS7BfzHLldOwei1YuLxA5K7y3iO++mskd0tTw574bRLpIBL+j0ppzw5
X53+Be5JH3oMGkdVoN1jUOfzbCP+wrdOR0zvMNlo1W1wmQkQOAHAi3/tIgP7WrM+jLVRPhdQf/BO
9auZmivcSE4OlyttA+RihJtn5QkHJv+g8h9WBNQFK1lAgDbb/lAhcjunMslRD1yXaRVB4FZBeDEt
dkHnVjXI3/3HPYZY4KHrmGcAVLVcm3C0m1GQlnjDoDAoHepjv+GEtb4E9efCTkQtH807p9f/tLFI
aMo52SYUYMh3+NFMeNyPmFi7LaVV4GMdaC2c2RIjmnaE64i65Clz5+B5gu2U96lnZTXODN02pHEX
kMFv1gyNdY7OZRjGx8iOyZf8IzpkTrkUxuWUh/Z3EDpZzIqyxeB/TnNIbFrWSWHiQD//zwp6u+H4
yHRhmJgHet2KiZ1pDiD9Kgarq25Yd0eNOZORrvELm8vdYpH4wa50olsZke754sp59B1NKBFsdJ4X
auruDA/W553wGTaEfLflM87j07bH5LkFl4rusn7GlR2lzV/4DR8BXjM1rLdDRB9EDWIJVE2r+OhG
19VHconjeADt4BgphsFpco2IpAg2dNjYwPOCLdpG5hrOFNRnHhJRud9vx0R8p2KSA8ZwymuXgAxd
/mThL5T1E5t0sAI6/O8B055yljo3Hgiy58aNPxr2QyPj4p75rrVHvlWwn7O6M+T0/AKFsT3XMo7u
27cFOPh+uNIznGhGfunUD7EPVFHZYDDaSt+h3/cQ+E9nHik4atFrS+qhba6UhuGfLo5HqDwxs8aj
tXmteUMvBpY77eSnEwse76B+xTDP56e9zU4zLIwbFOnpiMPjxgrNNP/OajAqBIvj/k+0T6S5SK/8
78Kn+zmW1MzoMi2rETqOA3XsQ0cafnDEuZm51LlB1+I7vkKMpczUUMRCQe79JYgASaoHjabBXror
BmxF9hiFSsmZLFJJMEC4KvH9SJym6SKuORyyLS3Ayz9QdpTX3A1wLty1VhjcssqrrsSCnbzgGB56
2Ob56SgW9wD4++8YN/isQNeQ8ZU+2/3Noy07CJvy2uU9CsOZqAhoLEYrA5V6INRjjOP06IXCDCOA
0gzmnww6CKS748F0tC09XkUDVmwxJZqowEaq5G9tQcclOIgQlykjB4nB8f4JEtebuWUx4ndNjIay
i6J6GNceH3kcfRJZW7Xxud9WwwtVPmlKyndD08cautS3wJegmFlundZtdZgF12aiQWXn93nZGg/t
smADF2fWIzz5hVoc1jaP6BAoJ6hxwTtNSBcpOIFNTVBn/VpXOlKs1Hh9+3XsbqMXJCre2crpI8NP
S5bnSgbhTx7Gyl1jU+D3rtfV/qw8er0r1YaoxxftTU6QbcexAW5Xn/eDsXIW51t9r4t2WLc2kCJG
EInM571TmxANiKJ9yMMDtofw88ZKFAUqAo4pZE1/JFrERHTQH3JQP9pnGuuvv8H9r+lYpW78ZsAw
eAPkB9Bw3ircjD33PqHmqm4LAjisvRNt2VEEC+SdYSyflS5Zi7FqzABcCs6/5KwwaGDzytqsoW59
BGlU7sUwJV32da9xbLIgHt4O1sGO3wWPt89cler/VFcIr4RfMPnhNB1MjnE2QuiQCtFqcvtkYZYD
SukLM+s344x9iX+RItmkFzy4PBH8mYddx5KKjI/+sJIt2LzFV7VRiOH28RZlYEBBaXHXEzx7CZdG
XXgPL5vkekRPNS53oP81AMZNxlpsG4fpRxxLLCDxJqtOsGHOcZGfcodLPr5+BeEgxhEM30hRSVsH
IHETCoOWUUAfBRwkZ6UHwauky+V7Ft1TsbPzVEh5dHQrZjb2GWIfOKqoOTNf3xgSXiHvgKIRa3UM
egzFAyPQrI5K+SIswdzDWdyHx9sQcoNRixdTsLP0gR5DKZ1sn1Xg9T1ZkN2mATBWC99b9ZF7HlN/
/00s2CDYiB4Wx2eR5ciNgkkdRBHYqw9plDLiFbHVte0CN+xYoz8NiLKEhE6WW7rCNiaBhg3JDSec
oQHQtSSABvjGLmbKc4c+moD745RxZ2bhDNIcgKQTQgLye16SiC6LZ3mLz9En+VNXtGmJExv+5Uir
vpugJmF0Zyd4l17jjPaNoKwRCx3KCOXuL3SIUts8+0KXNaHhiiPs5nZMDx/0LSrHQpJldPY54uXe
dzmVVfCeZZgizJphX0aqvImIX0PK4EiP6Qg3r01dKJ1zwHocdre2o9Ths/rXWnRyXgYMdBa8TIfu
F+oRXdH5CwXWWQqp8L/IBLDETBb4FEuIY9lQKfuNhAPF2Z9nwSRr8wTHV6zeaE6oB3u9Jds6BaVY
yAjBxjnuleBhk4tCLEf6NWGc4hctICB4wv43fWTAwGfnCXsIC38DR1Fvq9TeOneY2KWCiiMikIJD
YugU0qOTDtn5ryEjAZQGGM81uJ8pxZ6EXXd/7kpL02ufVoxIQdDDQHsiNundnL/3iW8uc3cIoWbV
6mk9/nODxFGMM43KArwwOYPqXG+fF0Qe4w+ZglIaCD/6LM+VBqdkLBCJpHkop9nRyXTejANFwupC
fAbCCDtWfkKxGMU7Q1+m42ov2CIBl8wVPa06nsiVMA0WGT+9DOy9bygzMVXsYaKefAuH4DFaXiha
0S6YFUQpNRd/c7CZLxn24B8t8tgAD+Mg1GY7rFiSHjYn2skEZ6fc/QObibs53w/t2P8g6sSjz/Od
bpvqlbKsH82Bmek4uAf+yvnD6OAgp6/9yd8Ii0PQKx7yUAR14dAAz8U/1bQ1kvqgEZ7XwEdKejmp
HPNtk53vPNrnnkBTmAT4SBswg+2isWH6g+V4SHw63T7sNBzbGLKKeXszte5qPOB03tZG8JWIpte1
iCoGQT85bd2jByKF30oSruOLpwE7pLUlDHlKaxVMnymlKesxu746x/DWWSYATlk+T/ctmB/4+NZc
3bKlDvApcIJGfXGXdopFxM6L9Dsb9A2A1aze9ZcEpjsF0ZlSEUj01uouagBoCVL4ua8cxOpnPIZC
zf+7+8YFS67loWrHrJ3VdondJx57jrYyooeC+vGJ35XdLJ1TV1YJMU6wI6hJ3KU+0qHSlpA8aS7F
DjNH5iMplq/92Csngk47ho3nLh6pyGY+wfnEHyrWBHBzTNRFjD2bGNAHBFI7FL3EaWFIqDqrHp5S
HEpB0jmgd4vvxmB+3kptYz6/IiDAWviryJaBkaxLeut7+Sr8VM70Q1WvnN4Mqtgx1qX9xXHM5zYn
aDYVp3vLYOz07WOsNn3sdQxPI6x04qai9XfWPnL8NDtxg1fbdznh+12iBid+07yF4Owrm544TptJ
pey97dwXLBw9i2U3yxrnGt0xOZeRum7Ddm6RYhco2fqsEg+XmtlRtT7xJwqSivkw/MqReIF0YP+2
ICJ/cz4NFE4MxRq1ktH2JeNZo/MiDCqCMF2SRSrHAD+WIjSWY+rJVkrvksW64AARQxk0Cj9aT6Os
TN99EAtaL1k5ZNUe2xwku3+2H1NYD/0aTIyHJI100Ys5ng9Kw2+n0RdlUpYS9fU6wD/0y1B7LWu0
UZ4yANolTTy8s/gz+9JPMshIsnBJl01t88HDoglFreqdt+2X4+JEmqgng53OY8COj0n6yTMn5pje
T3UduPmuh/9nlldDr5nIK8bnIkTUQ0OqYp1bPi7eiTNdvHg+s52TeuwCYUL7Wa0ntzXC8A3A05Zk
jLUH7RaYAJgQQnzPM4zyDX4C6k8ysn23/zSOxQmJx4SJ3fOPejoSGO49Bx2m0Zc0gEyF3Ppl8pN2
J4Vzh4l1touVC8hDC2I7zaVOY0AWWCNa9Nn0zsZdnFieX5DS5SuOgY2RND1mzgYBWoCd459SYb6n
RM+gW/6+HLNhx5mLnyE4vTwsEaU3sKjmbep7a9XPPtjNw6A94/8vq4OpyIeHiU5hrCuLpEqnkSKM
c0uoh2VpBL465MOj+k9q/0Ha3Yu4/itWXFQhKN8xauWLkBz1CUXVdHZuy1LwocJHViTEv7ee4xp6
63AV9WdE2Qbc8kGkVfFcNlWZP+PJol6NDBNo3AblHEeVxUtzKMLQplRCHSMxF+pkgkIvrlHtDodf
lzr/X5hqAkAmY0qVVXjaLBBDBTKy1ND5a+ugMe1EehuFZsARNNXWi4KFRE2gjWeXC2rgrLtWMxOE
gJ+9MxNCenaiee4msGWk/cyNJmoVpcrHdj0nd5spnW9Yif8ClwZTkxCp2su6Dg70MBWfHEJrwnWb
ROo5SSwlVm7I1CDILXeTma13Ml/4f390GpGNGOzQxbm+mwieAgkg2VPR1EL0H66f1L9pmS8aiMVX
G29sAaBq3glbmeswh6assxfLbJ+uI7sr+KQABIhuv5W8bTcJvuXsSVVSngRx5SoslsF/VKd89zgQ
4BMCJUg66823WrSX6TdAHUyMpJNHglV/YTsda42nVMiFv4fa+LukBNLyOPdDZJ10bkmANzr8NqB6
//ZnTU3Jmw6MYsGdzqzGqFtsl+cmar96Bc7/lr8wljkaLGE4EGfJ5GDTgRfYMeYPbjl9VPoo2Dcm
kj4xAsOY1cbf2r1PcGx64iZub7y88gEUCfEf332CvpwvhWLDhaN+8/BkY2bW1QfpTLvqYiQkbowd
98vDQ4GcaYuRAQ9ljQuibWRGJ8eNYJ9GkAMb5vEKu+zcl+HgpQ7gEn8qQzd5a6U9zGRacc4lsJGs
hmSBBtE+YCjHZyB+BfGddoS5ITPL5ul9xAEqPCx8eHQ8sDs3FsKG7MdtMcCgkmNwd3Grz4sMscvu
M6Wc16AgYWmjxvlsDwjtSe5xAjvs02jqDm0AcrH3fRuJtGiocFaZP1ONZSVM8ZqxMuwyeraVEbYF
w9Df90fUWfJ7UcKDB2jYc42ZVrQoU7QkLqepavi8JT3SiAIOCozdGSIP3Y0PW/yIwPQrqTyZeScb
LHfKpYmjm7GNv8hz3X5Jdlh9u20cWkR1aw0nBzI9yG05Q0zzeguQQ5kh81svagZfvpioT8SDwayO
QmtKa7XVYs/n0WJIZstu0Nzjbi+1uNxtF/FBY9cPAxDY1lAaTU8zCg5FdTJFnRW1fhU3vLk+RWuU
slWN5yCcbvjWqStr1Mnd074bgNxYwOXvPQmhl6b0zbfkLj292gjAEv3D+eCJ7aPzHNNJ5ohmMHR2
rBBL8AGpzipGyiC1fBWTsvchLju047CGe50Iw/UIkswdFV0+otkXhM+LS9rD8z2OcuPT7RtNFvcm
5g6w91uaVLs3Xw4NCyWua8tt9I2Q+PluDLqp90f0saKUPHBdRdQh6HFb9NOQKlR+CKxDGLNno34Z
H3TpXrHv5S2KVBkZPW7ERBD7lKVfv0D79sxG5OZxHm3t2/R0R1UMLZKx1LSjZpL7zGozVUIsQk+W
ju6kw/ldZ5PEM5NONQnO6D2BVQpcYqh7idTZ8GDNbEYI/LnuUP8Jo5eIFaeaD8teCbiDfaUCjzdd
JRw3O1c6aVbXNQM3olgrPJS3aW+NRLvCkZESz+eI8gf+1FC38bsJQLPO5UDxiadhgl8pqwbFJSFr
w7BdL1QC2wY/yLdppY1h3cpUmMlntOgh7/P5IQtf13vAKkifT8Cf4L6K2TxqeniVTp9HLIrbXkjn
HYTfrPeGKCz7RGSK/nH0kYDbf1KK8JlJhMHCPRUP1jRQRFUP0clCMLurofoTWDcZoJ3xBQLOC2XI
6Z1kWwEfWfw8enXVR89Grs7MDZewjSKFvPs+nrC3z9u6rJ3APmpV5rHbjrg71Dz3P8fABLY2vIll
e77Kq37FQNu648YUc41mHO/F8yhrXNY+CgALCDJhRWOHHSs46N8rgyOuqtoiBSELPrasaPqJJGRH
LmUoGPh3fj3YcTsKsqVXewOPj1eHDKnA2+OjqTDAaY0dOeLGlJ1Wj+Oa3tiH8SFoclJnm6tuaqPm
gZ60Bhxmnab8ACIjzuTYQCinfYpVysuG2iyCyyP7wyUdfDeSJvKo2uLVhQKObujAX6po24zVYZJm
9uiwz51IYsfFJT4k3P7A1yPbgq9xuLSlOohnz2SxmCFmysV4zx0dTfy7xurKxf3HUVVSdx45qCp8
iaQSjasTy/aif5Z45dEGODvvQepvmMwjmy0wcMZoWPUyq+UFzAF3HBisCC4MCQqv4P596xQB3sO7
b/LkPFTNQRHyd6CJdvI2aBRQX143saQtBmGs9dsLB6ziA2TVv34iPu6rF7Kb4Y7LmIxD+fhtGqmh
oKZqxmF2xVTSEe3IIdUCSSMabEPmj3R0kNaGzlGZkOTbqTkcj+hiwRD2BfXJ7Wgy0SbtiTjwBoW8
mYF3CgdSznOkB2SB+ixe8VK5Ab3rnbjTpb021O49w9UtZXZNdnKOKlgg82u29ik9nQgmXXTtAi4x
ZAaDLHw6s4WDD3xj+yPDI3c0s9WQhUC+SypUWF7UWubi4U5Q/tWYFEgKb7Xa2gpYMR+eDE246gon
aK+rzpekmLAJhoE8nuMImQif12dGtqyl2/zT7j6MRT0gJOGKNcUaHDwLOj0gADoUsX+PFOTnnIKg
lY/MLsEsl/guMknbII6/h8HC509JaIEq3E889NDaN+Nui0WIQghVoXvwTfpN2tQ4jdbCPxDV4fZO
fTfyaPAJAGz3XCNBPDk1DOyy6IX7fI1ab6asGF3ITRxtVP6+TbGKy1hO67xPzIeq+a3BumZA/nTM
RucZxzybGq/o4XHJA63rfnokdnZDvAfbXdPamtvlOm9iAfSMgPCoQSeGl2/PVBlPnvP0RBNL4oEt
ACngoPHlJMxBfl6xOwfFUa35b8Aekf12mmeREbTWy5J3O9G+sbrTurZpvafTIJVMU8owrpdSqAsn
Tavc4+fStCSCLPl5Li8nk/ZVPzHNY/mTANxne925TNvzNBPdz/XFq+cxzth7stecR3K/tGByjOzY
OlexlR7ZXVBxGAfF8aKwzWC+UxNUxbMJ9Y6bCZkBOhy41oa/GwBGXYSzA/aESXNOKrhyiks7tdCX
r2pN0lZ4ZVIoJotx0TtSZSkri+6lX1T9IHM2Ik6rhJeTtVFduYVJilgJlC0Q0+U2RKBStrEf9ESo
w9SQGWgNQsIk/j/tGABfc8oKNOLnXa6K5wI0wOkry0SBI6gu0Q7w3Z9FZCQFLLxz5I+WM1pZGr+1
qj5jeuepfCzkVEpnzWq1/mRjNEdU2abX4YO/hfyCcuP1eSI35YgIAQK07XMGDOfV9Gqa8CKYofFh
/XHinfkTMaWEyg/gJzbqRfLxGSvemH+xDjPlNk0riXnzz85R93X2xNPKbGXy6K35a8kNEYDwSo7Q
rq/mR3A8maXcG3XLn7JgCN1YxlKQMic5IeksHa6BrRE3Dd9zuxUdjmQFvFo8UTEIBj4jZCRZB8M1
W7Yh93vmIxypPXqVU3qz8IDoa8MErp3uB1JXt0lyasJ5PXSE/4ukVFoyJZ+wjhjkM39NaSFWyiRc
NN32nJzNm42+BE/5P/EbISLcyimplpjRrmkPG3ewuUvdRhvbHf5CCbQwAZ3bzhRKMLQQ+mwYfpYk
ENLW01pq5GlHUit85WzLqkjzPb2gY1FExYMhGHDsspT7yGSIKgG6HRT7INFVgckfXlumrwNyPks8
xuYA8M3/nY2/26Sk4j1xJZ3p5QbjODjxlKc4kNHz4LX7dAnLdcU63P1L3A24VBWM0N+zkzsjBQWR
74/2iWU6saRax0X1TJxO520tRFvWx/vbA9YyFcTiEOqTs2DBZji2VZ4JrqR5fYg3rSkfVpNrzJWJ
23v1Un15ZRAolqg1MVqZLmr3Byh0RQX4QkcLTdlDxsp+vXKv3LWkjpxc9/QgycM8nyIclP2rM1OO
3468wGM46QUrHyZx+ZkjvWI6wMofK3/loGP1pIME1e4nEmyuNM5J9v9zkrK/xTsqjHjUqkhaqgyn
Uq8/gfryUZrFQscSbwYUgb2mL4X7/mdu3yiH8T+JofE1IRVhrXfFtO1OjedIwnGmuCyGbJg2CWhx
FJ24hKnmPgnGbiWe1MSC9zjb0MsNDDLlTG+KSBwPF2ad+FtEFzayiTRSsq77CsD4LW37I6BFimer
AvNtiMup77js+0JgDr2yQO+SpHshY0YVMri2ij7jV+LHKYGc+OHoMeRlro/SnCQYkmydRXAqvwK0
FQ8vTZQ3S6LbYjZy99FWYmuUP7SRQ7+gvbk2ipr7Q/PTT3gK+qF59WDpu2JvkjK5EqP2JlMV5Jjm
R4ktQ5a6moqJzizS7kx2qgIF3o6YvpUJ54Tzz7yMKtDwrhAGbY3m7Wk1q51tNV/mcnNPcC/8F+nu
kSxWbutS402uOksT7CD87dD8RUhZF4I2bXYuWjoUfltb7gXUfM91og4Hx/zC0bjocZ2zEAPRGXCj
vZcge0k01R8RZTpZT6Aa3DLDJhw5k5vdODQFZUPD/bBv/bU1cz7gXFJGPP+60aYr0RhuFPjmytTv
9i1B8HEqNxTEbAy2p0pTgY2kADFCSPBjeYwZ0zbTBwYvsrdbDy+c/9d28uCpzBjtle7ofQtwa8Dl
gxrxZWyz7UlTeh4hBIUyzeMVIQN0B+ViftDApn4jcuFBrBKlg6ZlvCSkMrqK7pqmImtsqUEI6Edl
DYaq6R5Q2fd/vZrq7y1D+JjvzUUXtRVtYrpPpyY/PYidOAY8g8VbgJTauBtd+gCjd8XntLVnyiC3
OT6Nz8fwcd1HgrtfRcW+ZtdXilasXl8oCNk+yTkLrvh+EAH09GaorGmEGcTh+iWUlYDSUfSKcD01
I/vcf82gpFVA/3RUUCBg4hyONl8d20PQmW+GBMc4f/5bPUM7gZkgnL4NW0NVIgv2hyLAAUs/E7NO
I9rBXyLAF3H/scyrWeU3MBFqwCu3zX399Pwi9o8iciSdwE2QHKcF71MoyNcDVVnSD1Ivd/Yi8Yi8
tDOajVBsAPERdryoQpjHEC9n5PUjYMjShaWZB6b0SXN9/C8x2YpAZHk1GYIRiJcXXKITTZBXrHAH
chmRkVRjbH8zvlQmE494/JWRl+AVHrzDqpF/eriULOaZ2W/MlbsZtwsLrEjWmS67DQ4DquZ22CyM
iD73dtl2Tk4pvks7kyJU18OjuMRJJC7YcJDghamCWb2K4cS4nml6xInI1ta6AiLZ4lVbpWzGiFkZ
tIdsHLGHrSzZYe5ix1ZgVU8u19YnhFpo9D6QKqESuBuIpWwYP6Zb3wFqZY85ojtMvCpYaDELUEj8
Eza/wp+KbxIthNXQlw/ywOOYx0PTTFNey1yG6MmAfHeP2fBThLo16laUYyaNYnbMB1JC3+Kg20jz
WN5mKAAxO+WecLvSUbiL+0B1Q+Jdv+2L3KXqCVQyTxo2I+4dbSNwToh2AnLkQAKFCZCyrwMhDlTG
PhYChMdzvmSX1QWOkBZOKcSKS4xPgwotNiju5uAjIx2pNVDr6KG2IrYWiowLIJwhTDyzo1GmQTsv
k3/LjWHlwfmh+LJEzhmAbediEliBkmVc0b6EqLzsXyGO0lIII/UNX7Nx8PHcuCJFBrXlMhbiDSCw
oPH3rH4cQgVULflu70KrYxWhpKkhOzd9CQTfMqO7Vu5CLKmjdnmWbGR4A5GDQkuEbKnLaVLvDJSY
QP5/V1BbpR6NCYbPsSHmqOjbf60guVWYH1BS9MmZXkkYi1lxXslATlfTxrr8+slRXpxhGQ6JRx8Y
B09TKYWE/O9c9N9hrBLNoxs+5/Gpo7yHhjY7rZrQRvVrk9KtdGyNy16UZ59NFHNbIkjAw3m+tz5m
xJpO3X3dKKOdqqi9aPMzeuN9m07qLKkCtm7Vq64JfupXSAngO8CJCwIjPZtADD6lWDW9FTspWy9x
dlwpTuBzp9foMDQ69beS7cmoS9IlOyAL1ueGzDTqSPG1QShi8PMZQhr0jlVWzM6p373rUmCTMd5D
zATK4+1GkxEZPV9xuxrBLSg1hf0pUi5CRHq8KLxeOkCWmWcRVCTjDZkhXOpZvcs0wANBiUrpGL4m
pd2Oqta5MHZvwhgpGkmXarWzbwPjdkp1SupCkW5D6N0zWR5oYYjn5dnQKvyJr7YAdMGp7/DYS2NZ
nysFqW43VWrRPopmbt6VeiN2hhUN4W1shIy/KizSk7uGLdkS/rVzzCR4i1a4gPzblmEPKX6whtcP
fufpYOupeyIAOY1sHWVZ81KXtYo4FB7QUKDCRXEFwY3JE+4juqLGDJpQaRqjPOY1dCGb2B1Kaogj
fevO0TS5ERccT5tCH7aOMAUyQ/ltyCvkD3ggaEAzI7214GvQchmA5YR93unPPU79ZOFAHjPp0jMr
slB+GPg/q7iyZcOpuepULpweNWQBc6wMbFTDFXPQputuVKmrd5NuErH1bbJIlqpD7ifDgl0iqlbr
q29yw92j3IJ4K23mnwEWUpGB2iJ35FcC8KawqNBIZ5pMhvqQPOeWPTUKgw/S+LoqO98ymp1bpYCZ
mRupN2SuuHIGt+q4zU2HDPWVXRUvBXGOo3qaxBKdIRi7H86zfja5/mAfwmgaephLeR3DBLjoYGyO
6wJ2aw7e6ek7Kh6xJ9xMYn3jjQv47zGSNI/QSe6eCBYRxVk6Z4M4nteceCl6gej0LFwuCxPFnVdz
7LBr7d9txIxkOjReO3wPSkzTKsCuOuqfvvU7Wg1IFsOlMJm9JloeYDemU/aiF7fsellKlj2/M2p8
7UUxWar0ly65QsvjeHBtRgMzxCkag4thTwXTg+k+j34dZQa1FeH32Vsfh8cRmBNxgd9/6htQqh5v
IafNbueJgZttyRkpO/GIdufFXV/Oy1HlQc/s0iedmpwOIT9tnoTu4hJZEC5FkmooTPjdGuk0AsPC
5xbf7uCQWPTFBzJVhk9PupjsggdRFzYqN3bsv+RH4us0GyB40dD2YXyUVecF6eh0TAIunYDAqjAm
8x8ycFu+lHrCEQSWJq/47Wzxzn26cBBsRT7dhgXbfNlMKyWVijxsuxb35L+WOu0+0Lo35VqJTUm2
NkUnypDrp8Z7MzuWSpe/28NHWbuRKdLDZOOMN+CMYgbsg2L1kUk7QUuHzy2zAZjk6rM7G6VDsXY1
AotDuvIUYFZwynzpgRX6ZasqDUGELQo0C3sf2hJ4A9/J3o8gv9odOJgAM2BXKoK0Eb9maT+cKkQ9
mbjVB+ezptdbA9WqepZyzZT9eTmOt03I/1m+UAHfy3ictLpRUNAsxzr99u+CrBByrj7ASNYrNsdX
K+HsL9pNLGIEEymC907+a31FsdGFjgOaFZQPxikWz/x8ERabcksYkdV7XT9v6olZKqyqQfIMFAxd
7gDy4wqVe/+X/bd0uGLpNZjoAu7u3dTWjny1ucjmnLTCD1kcnVdyZfooQM//2tNQaxzmFNLJUij4
75UXBjG+3ZM4jZpz25HUz6ZpGKbjTXGv0w/c70jcvnIkp0FD8FuVzezpGp3GY8U6qWih8mFJWKWQ
wOGraRE9mHcwYzgJ/q7uQoPIQ0dajY5/0hQ3widT1HEs91NLY/lkfv25vmVKs8M8gkZp+iYvad4d
zEc4f9SrGzovrTDEUl5QWLcbwX1Dg43hnIz7QJ+YsYgJrFu/X+pkb6X6MrZ0BKhpSxpx70UEtN9E
Mg43BXaJ2aKcOExFMhEkUrybIXgLEvdhgal9wj5WGt/mQR6xTt5/GWQnNzOb/De35L9Dg+AFK/Ji
kjFrqYo7lYiAjW/lK5P7aFAnz3F9/NZ8lFT+5xYEHE4gY0jZjvZymM93NrxuuWBGDVojVD/pqofO
Kqyl8E9sgCdTWbcihfX/Oy2OyPcR1XQ9asgslcrR7iWaLReXRIrq/coN2SMoNGxiDs8i6hwW1TOf
IS+Avua+1eg+JsFdQk5KmqCUlLVNj3KeKnyosTEVoAIw65XZXm/7xp8QSjrekdiiFOYjYRIlLQw3
wVuZpAp8nPCoc0fSL4fmPN3mX5Cqh7WxdfdO6lDR69MLxD7NNsPIjl4PA50zHUefWnw5/u3ECEvJ
SW8LR9ZDnO9whQt7HRpM0EWGAo+MM1wRxtLg8IG41chHbeX/PkDEnqVbFKMHGNthFVF5n8qDdZmp
3qq6um06kbUyU1MzbxlEZDV7AkPIrd3Kuz75gYri1ULKhe/OkXaMSZr2A7wZ7YZYLp/IxV6eZ7Ni
OZdaAgJJoecKwWCQEGyOrtFnV7xkVgK/5VSfA3AvAkuwe/0mSk+edeJxCTvgm5kObv/qdjfS37Cn
lh8WDa8RS9y5oYZn9GLa9yJ7vcNKCsVK9sdxXd5Scmt37KtA/31P5kyQKUG+OSrQi1CXiWowuDYQ
1qQvi0bAE/RMA6xiQEweBvJpFvxT9ISt03j3zu3IjHw0gUZeKO6yHLJKiEmLnmnNJw3d3OPLcdHv
dduN0wK+twkFCojqx5y0vuvijxpYykjUsgWtfrHoMpo6pEYYm3lKh9mb8CNjsOMWLwtyf0QtwD9l
MBHHM4XjCbdGtcRookFrnh6Hk3szjvIKFLv6bvM0hkyYaCRarBeluaB0x6U/lCcB9v4fcFmB95Dv
Iq7vvn5DiTlwWxu5B2hJyND0tbpPSogDXQVDWA095lM+BsBHhEJbXxRRgn6aVG0+0F82pI+U2gVl
V8KjEXE4G16KBnfY2wD3+8e+AWlMlDXMsV7D1Kmoio9LwfCqKM4eHdbhuH00Jv5zRhpZG4ZNukSb
IsdP8WKSs21eXhb9bE2dKR4qiYAFN6TfAaoJ7Ns9rOwp5KGaKCivcEutE5om5efxeDcIGITvFDye
vKKziOEu/ELsJXQy7fk59a6ISMh3ITuzeFmGp2LUqyoFFjcN+3cc/d1QZBLsb9cGCsG0APOt17dt
hKFMmy6L5vZNmPvBsNhqFd+akukQxaBSItWxg6Mxb+Wcd/MdfNCdfYe3oabG4gE0LRYt45JrEl7/
Rq7y2ARKmDHOwxCffjcDoYDb2c3yU9vH/0U0Gx96I54C9VFw3nQLmSkUmAxMHfPG7nZZw+yxcyDU
lldDY9shIIsuZ86B157oFRtOGyyjeLhlc2Il4IApB8skXk1IYZfoAVLATX3FS0KWphH0HuCAtcos
E/escL2ctYqEL4odAvS6J+rwxyStdqOwRt8aU4wqPL+BiYFwGkG4XjSfQZYkXW4oEm6dFYsB3GJR
iNnCLok726G1hZ+hQxKBRRDYFf+JXal4NsF+TYj1uTN5hV8vf/S/KAy4iHi/1GvEsxpLCPn00IpI
jS1wMCkTCs27zakD9q4GUYW8x42HKVes0KkubLMypzSlZgFLOvg+6rVi3TYRwoln5rDdGp4/nSbb
2srTin8SJEbQUhFJqxhxXDWvvJPg6jDJatJf7gUNYQKveDJ7qe71KuA34sd9fOtZGL2IuQHh8h9Q
AM5+sXc4bdwywaXoeqtWniJjrqibh/LNQgE5+SWG1pMgu2Bcn9R+sTZRixXf8dasdud0qHez6phl
54BJPEoElYJ7dJZZhHnNeUXIR3IrgF25/LRH+L+8+ohadJ3EN0onljMEx8NkanddNx+0jNNMpC4Z
nBLLeNyzykoKnNiJIsDcM9GPFSKwZRtZy+0sN1bMosUHSJZEh5jVOrVE5efbcUKKafYfwey0YMN/
5JcmW+B5JHOPweBKIbqJzXLNPDkceJNN1yy0P5eXXtkfeFLv9VSFsQrMwBjhuijfZWa1Q9vyHLv/
pl4ekfU6p7x3flYnYiD2Be4swf9LO46WGXKkxgKVYQ4OXdTv8Lv17rbJ2D2Ejp+p39Ab79G7VZlN
7G1yNgzBWim2csw/Li4GTULD6/NZLBXmQlxF3g9sgize7gFHrGLqPE9/1KXZwLxuI3XHkjt2UAop
SzkdGRBmDTkNJvWIz+ZU78rZbgISGX1MRcnq5Su4o5XL28aWcrihfEYIXFe/NOynAE/FxkiUtDma
T8Ds+MHhyjVH9jYRUgXrhkOq/sgpaABj9a09CMPYCUCfdHQNxK72wcvVZ9gUMqfXckEz0KQJXJdg
87rtaynTnnhanj+WnICfIDW0WEZsnkClSi7TY7Sr9WAzhOXskwILg9FATjZWepDQ1oglGsNSEiba
6dPQpq06esH0tdPj5z/5rm9Te/9rU2Czl3aRrLDEDFT5z5NAgl99VZyKOlRlvNWQsYKtjA00Y/E4
JZITwE1rrixe5qad3PL3uzmQrFwK+ny09jv3RgUBP6MYXGOSYBbO33Y0GOp14Zx0jzj3MNkK830R
AaHKu2TnV36zFEbL54MOvbJZPwzd21NPUX6HijXgCKB/cwLGg5mTimwJiQjeakSELAjiOkc7kAJ4
RFbeWVI4QnIlFymvaFdszHpXT+pNvBm30wHvmtmTSWC9qYuWPSfjX/tGa5uXlUJC69+AF2jugZJl
EEqV8R5rYrLljsnrJN+Q8BA99ALiE9dSOBWQUXR4D7biBZr8dlln60iyPqrTQVvoPcltrzZoKIW8
GYUwD9MNUa7HMYyNmkkyiDBl/24AShPoPVRr8/17sMrCGcE2GSJLL6dkjaeVvgtZloD6Lvh54rrR
CmkkjM4DmMxWdr7/sXQiC/Md08FTXSE/aDYIWkInKywP1x2z1aGqxK4nmKL6Put7BvyCi+RmsQ4K
vynuGdJUXs+epOMcZDP3kT5M7UJo4Gl9ZkSsR4vfEyVWgUoP2gSaizIhSyPqDv1EfXWBC8NDmSvr
u5+cCIzmokz1pn72oZvN1raw20gkCcD4oVrJE8LLLGN3co9jI/T7QdV1hSJHOlPGWFff7dPpDaOC
5k1MbE3tFG3tB2zCOyF0yBx/pYdku+iRol6IOG/jBXNyif7U+1flJgt//1oiWZG875XZCWnNyCE9
Zkj1//owoDJlmAW+hVCAPD/iBtoPIdrh6H20hE+McQf9orPqRAqTQYHUB7qEsmHKmrrGCRliCsAm
HPDi0aC35BmmR5xCv+oRr1tPXMqDjIKMKzdiKzfe3uvbLrbIWbGwWwADqnmspJ8aPTUBahzbU39Z
xlvAgvi+7n0Tb/aX3AKRs3sB97RxoMPUZCz79+rc0dsw1BRZpywYe+dkB0cwIT03wnNHinYgQnku
beAishBpS2Skdi6uh03dlVV8WE/MmRiD0nz8qqYnbttNjHw1ugK7QFlp1tNlUbfi20yTPZ6dYX04
Nq37kovsw01w/Q4t28huhr+DOmQzBxqSLFRsLvaHtU8WFKGwkrmx2WsfIAZUBYnnsINwsDhZ3ly5
oiHAPag7yM4AcaoDvXAZlZEYdCLDnUWjzp8wdsS7cmGtzI7ogk4nVGEYC69OLRBYEchl1I3s1yYL
A8bhwSaAbyxoR0/eF55/Gp5bDPh45ioFJ0rtoA6iFoMff/wmjWi2yhZ7xNcG9LlFoFikTbvyGKUw
nNmiVyj+6LeVgZWHpt8si12YEFKwe9SamwtoAtN8ckrm5UfyCSe4HM41UHcVeuTOvrlM6vxX2Oht
U2fhJyOOiwZQgIKFMokV+QOvavqFlQaDRdJwNLWPHi8GxpvWEeRqEe39ePRilG3IuO4RPHoAOjka
HMCzNV/PlCnvo0fvVwoZhYU+Nx8NqlB3eP2N5H06xdXokyhAvW+FWcdVD9YnGVUkyw0wrDQyFBZA
Pupx/3WdgDWMv86f1L/x+W9oYyRTCBrsXhamlV1Ip7e0Rah8GkR1ZdTMM4t+SWkbHdBSHbON3TwZ
OBxUEU0l9WbtYBHxKOK8Kgrh9AjUB5KmLgalgSVCam7K+XUkht7GV+tOXxDn/2ITNpSmuK6nOAWO
1/Pa+NoaT0rCy3vTWX0LIrjZBt/0eLVQ+NPBJb1v4ZI4B/Kg5VdBLn3yru10LJHU5XPho3wz7U5O
ueinCPCFN+Dmead21H78kq12I5Ix0n+j/Ui47RGfZO3w1kErs8aBNzL/f8Kh29BdM8KpaUvBWUiv
+0nN5hylmDZ50UKlZ2OKhw93Znr8cbQ8lJnwBXwveDScofqDF4X9YU5wHokAamOKEBvmO/tqon8N
6/9pC8mbY7oetTwPj4871rVYBo42obiMhmUWFR0G65B8NWcrLi25xPUJ9Us+O3cpeLJ1XMFYjVkd
1c9tRAk04o4xHCXSzomcefb83jIsozqoLgoFU6vxmEWwGE5EtmHpVFIeLIRvixeYowWkjAL4PFHz
Uu3pZBikUSRQyx1XkyBVExeG04mhGsf/wseWuooICLw+4C90FmxDMjqkJ5vJcmWFaHKSUO4E5on4
ym8nB81EOnifgADsQgVcWEP+FVnT+erLZ/DTV8dOs3m3mrj3wDTlyO+E/hVN3xuCYO+noC9TCNT2
HGddJuZW256RI1ggr3B+r2QL2mhFrX+COnhwmCYUjY5mCG6HerUR3kQUNVjLKaOk2cNBVDwKXw91
7sVaVBc0uOW4ogsTyGrb4k660JcTzAhecqijz8Ftz3eXpTvi4rQf7HDKcao0aYC1VLaFHoVFGlJb
/4sl5KfrfYKPn2oL7Qc1lcUpRrJrXQhzs+Nul9pp+bJsDyArkEGLD0bctyZ6q+F3JCvCFkgLp8ek
T5JgF4rYbDY73WyuQifs2IJhTf+Xu+bL162FbBfXiQCUxLFpwUUkzpU5IdhN0bbWer/Gfg4Fi+mu
PlhBbAOSLd0+8IFpVuQH1r/ex1zX80JaLNghnN9cVxWRi/S2Z1y/qoOAmk9RxgQWt7JdDfTplssn
tAoB7kURbSZfgpZjNlTP8Z3FCv/ZfJtAz9dtaCpCGNQgH/NMnxk+Zexq+KoZs8e3N38/BmLFMjjg
B+A+z6jyWd4CNd102QWfBmDR7M6unVfvd9eomgj36VhdBTnMw4T8rWT2nbjEvH3qFRywoop0tVGI
g6Nh/3Twb2SGp7ge9lvUiXm/HSqwndPx2m1qh+LQP/RAcGRExaKfhkpEYFCakmVGmz+3bKeK6ilJ
MMfBKkaz7BS1COm3BctRA2P5sgRJiKsz7mF1m3L75vwaPHC/w/ONj6VIdx3BU+vnwvtkhExGgTd9
ZTjYdn2dwWEZ4p6YQ2oTZ93wHnhmMPvnjS9cZD/9QSfV0VSBxEaCKg8RgDzq6FlCxMMkwUsglcVU
+oNp1mWl+Mktecahnl9vzaHTzu8qfzD9AnuhoPlWTpwhsgOZPl9NwvqioS78eOsZolbomknCZSNe
ZWq4Hq6WOd9hKbe6lGO+yV9wqbSynNPjPv9AGW7aGBT4XneZ+CqiAvZPn4y+xsp6/SAfKJyVQ8rH
Twf24F3SuwfwYGdnFcXtqcAqts3xpqDEV0J/upGU/LH8wSiTK5MrcdsINgnLXZasHU8MYVcoWzXD
hsZsk/NX52y29qHJbK+oisvmZpWX905+NwqsrgbklX+7+ccjs/IvKNOpkMuUMnyYVskZlY4qJ5xw
bPs3XsRiMVqK3vHsXBtn1AHqedyFe9b6KB9Sch37hQ3gOTwsnGeuykbZYILSgnxlpeIYAORg5CTM
/dHbcuAFE32FsjeNMldYwKz4OFjZcLWTgEbnDVlavdpBOdC33iRAmENbEEBFQD5czZi6Tgo37pPI
Or7IoYvql51I129Gj1JRy6vEBBPtlvXO1cVxwyut2bRVo6LcYo7ahHrNgZxL7HAkSAH5+lYjeUai
JL4omBD1UzfpHFESJTRICXBSVlEIT2zZtDmHao0fgmsNbKw/ZdyfL+akmJdlkv+WU4dsL09H6Y97
GAzPjDo//WsCfFAJyrzlIw+ErOdwAZhm0jQnBNtCGoPNWPGdr9V8jsf7HAcvGOtt4DhyHZwLGjq+
TXXMKhBYI4Kb1yH66LK9jP8dnrDljx2njCgdf7Cf8erwF9OheFnTRYtpyrqtQrRmRjmSZ7pXAwkm
VJKRtusa2aF124sFc6zJvkjUlU5oPQP1m09Qj/GV82u77sxuoZTt/msshXfLWsD60DW+kcbiEMTf
w70vnGAe4Eh9WS5iflCHokOSvSFalDKdjdpMgzpc45g6r1M83A+8hms1ZhH5u3t/umfK3vqp2UNI
DgW5jxB0+3u9/HT6hDLTPBAT6nkEUF483dv+hSU0OfuYYh0qBLLElH9CSRzWm08K8s1Thp/6hoyu
Uee8oXruVh3nimpGsdF6e4CpTGsU166Uo8R/gme5knVHI6C8pQ/WEa9TjArAVs3AQnhdh6weZ8ja
AFzH7b2Nfzfg24xhGlS+kowK/AI2A0UuoprKxGAcnxoZhN3ancxy7LUnfcV2pOfpyOTwFHkgzpPP
HElTN6gf/88KBJ4lkC2CW1L7zC/3r96J2YFdpdNxBqodW1peJStN2ADcQr3VuIdVIBaGR4SLYNhs
4B4xdqDz4G6Aeo9mqCmpCXM3vyn34n11C/qZE7Fr9DrS67JSV24+XinoOjC8xeXr+vI8ZAnbcMIY
tXtAcV5L26z3hWUjiir6J+OGsuOa1vhWGmIHBDJTLMHsVVhKxGGpy1gvmDD5AHsTeuCL4PLwn4oC
nTZ8OiPBFcdXlNbbvDdQSU2Ev7YIp98heNC0A3ABTGw3YISS+VX8Gz/M/I9vIOm2r93tP/HpEu8x
oKpIZxHYnBQK//DaaxfLa8rBN3PmQvjMhmyRTAtPnVFYV6BEaJuQviL2PaOtiSR5RUEBdhpmYRSW
gvSw2904Fqr/rLgNE+oao8+aav1ehQ0p659V5hE+4Xh/LFqvnitvQUGL7hn8AGHoRbpqQdG34AEq
zswKG4PTQkAPYgRahfEPzGLOXyck5js5dvC8wYoff3HxFGHKXawx99X+EsSucmbpFhnXmWg3SppL
BPhRUp2Tp2BQgvq4JyMpKeexNcaNJKKwF5ONHnv6pivdg7jBVCx+wzF1v38G49wDCeL0dkwcPm4i
G+aRsc9lsmg4c8icZfoAMS+x7sla9eVBqHCchwDiKQTRyYHoqNpHfAUcD03IMPGElsXunhvgzx6h
6RtpWCUpUSJ5H9pia3oLP+UhahEq2w11n41Rff0NUl2m6lw+BzjacowUNN3wBmrfPsrMskrAoy3p
/bOhe78sUDAghXfcCuwby27eIeznU0q5QRFeMUr8PFSbaDpTRW3GDDeR+hRikDPks1ZgAgIf/cYn
jRX+qWLgHLWc275+TYCGO2ZwFON0V4leURVlZaVxuZ46RqFVkr/B3hbpVBksaqFmMd84CgP8Cq8Q
B6hRp14FOx5djC5/zev5Qt+RCeWKWPejSmQ5/dmwdlPIm6DMOs/SR3IDWHBR3z4CAOVbk9MsAGYJ
bH5Z8Wo7pJVgDSXo/YRf8h/LkAkA4JPaXmwl+KQRjC6hgdQwFTZ+ZsnIMLa7xbguT5J3r8+6MdTA
G3yIaY6IWTdQYuZaNu5+fuSwRkLmxsx+ZPwx7vtxsXHQvi2FR3c9HtGuxRiCkK04Z1+lxgxexu/F
4n49bsNb38kcCyaaTymHU5bcUxhkGWgZrRTNNoOkg+nd36wcXJcyszkHyMKXWwDqJYgd54GOm31b
3cRVMocMmpK6q4rmX0BL8BwCaUEZilKadtwFJFB/soEn++NYNSr1D9hU2lcreAlquLIVg5e5BNOx
M8ytQTCaiZc3r4o0uQrsKISIPTZN7yuj32MdmoLycI8Yvc2CUoDnOzc1XgAEisPyF0pn87JYjQ3S
uLKMziXCjdjTifDRkAbMF3TyJRpeDUggmShCosnQRZeJrlLvZrkIDShUSd6U+doir7kXF6yh2eyw
Rv7TVuIwYTdjIFE8QQn5AuYQwP4w3ech/Fanf4f5QZLqm+WvwGdD2dl1bdPIvQGwZv3J6YNhTMAU
aziORCvS4cYlz+yMbWWixYt9hc1/COEYCfnSvC53OCr5QGmPncI6kslruaC82C7PjUNGM3DBFJdq
abJ4yutwaPr2r8EJWPOJD5lsq6LFnISAo0uLSmqXbgxBpbrAPlYhdmKcc8hM6aE8G6VPVOWArVxT
8RZabmTXAwlyrNa5w9PA+haJi3uqpVxxcaeEheJ8nH9MyHVophp1nmCF9wCOarT+dBoJ8zO4KiAc
sGUz73XCdB0EG5vkagJa27RumErvNzeq4fIqRprKl/I8zR/xo8HDAxDhnD7YNLvLMEE1vhCyzl14
4lltp0KDP4/7zaR4W+7YdSfSWrgBYgiK+K868EcBP52eGqSu5WQkDErIbZaTg1vGBEgtC2JgWyKx
lsgSSN+ULUnn5zE4YZp9OIuijdGElWik6DO3U+oq+BdibEOabEvqO3ZIao3LLIqfPJFUib/JUVoW
3H3MpHRARzuTBYhRRBVPu8pt+k2thSgzegskkn/qas3dgo4Lj5gp+U6A3IhWw4mfCP7bj85B0hZs
5wIJ82s1MBCK4DaWExk0Fjq4pK1LtmdFDUCFjpXhCu+ns4nxC8FY09tQbU+lrXgSVeFLV74AEqYG
4J17QtUtmPMF9kN3eQB/VTlMNKZvIklMtNr1koPnpTcBhwXpy+PEkAkDCqwRSxp2Ss5XUtZmBeIj
hOUpvFVu6/H9LeAcv5wl51jBL0k+jozEaR7s8mq/Q9f89uoSG5bscG7g9U+obDY8/axG4ZSA8TMW
wPFkYZ7iir3ls9vl4uB/mHhdD89mNpOGQmEBAgkKBQfY3Wpr8b6eGEQI9RxcEeVEJUQg4h9crJ81
bPSh04kqIok1WrmqrE7jT844/sdOawzP++6bk4wvKteMOeWGhr/jInbEK+ADHuDEjhj+JQnPELyF
m1o8lhdaBs0Wx7O44ABGRBOH17xkpozrx442Kq4JbHsUfFx4gWqYCm+/3I24u8b0pVWNanZJav5a
K4/HrEreyyb7obZX7fJp1vIiQto5ESQGQu3hwm/urxfzYhOdLfUiTVdW8RVXNXRftTnqv4aVvbh0
qsst8GoX2mLjVUUiElGOM2atRrKPMuRIU7EGVXlFQFEwdZ9cc/CMmFb6+yygTsGkHPgUeyu7r3LR
jO4DOQF66fgkEkP9VnYxIUP8Pcy4vG8+RCZyojuRQkShPmyzpAHHzYX5MBo2m4B19aI2+trUyO+A
fiPDGkm2wTJto3aVrg0A/bw5aeUKa/zRrDOHbBAgH6sLXjMUyjwqxzSpbyUMT3elNou9M87Kjn57
PrtYKKJz1K4qK0XQVwnMQa8Spava+3Rv2yXW1eKW0WFJMOwxxRMpt2zUVVfCw9llzOircfCgpT+p
XtTCZc5snv2HROUyFbd+TGEUj8FBsgwbyDUCimAFYR+Uc42ISoxHdKuc4R/AZX+tuUJIImv4yY98
bxPcD4R6D2ogfqNwj6rxVgey1WkdubXxKPkgy8FT7JEm9HRli4loiFlDuqFM+FPl+/neh3poluVP
VNmop28BO8l2MIZlGsuM1rz2Mcr3ZeoWD7oN1D43uFBW6LSjCJxDVaMsTjxek22VC4GOqTlIxjHy
os1gNne7OGK6al5eo7dhXq564gset3U5Jp9JSu++VIy7b0yeGcFtbLF3pd9c3PHisOVkrA6qJjUh
1KTncWAM0oB8Wo2g5x/7eaxp+JPJz5qzpptBqt14VKWzJSGEewxr8EmacT4lkV1NWbtEiVmvzBs5
IguAukqrKGoGnEUe5nccXxMMA0TSToikh1uaJznz/9HR3Xm6kTHODO4VmKS24G9iaLQH1kWhDlIK
pkdWJ02R6iGKNwph8XYF6sys9ynWicr5YClXaqGOAvs6sPupmi/M1/M9mxyw95kdWbfJcIePGzUC
6yEAZw4p0LSpbos7R+rVFFbIlBbPXJAMuzY9EpHiTJM/GEvdeUrmt9gB85s5OHGrHWHzlliSi8Ch
enSZqxYMmxSN0wsL/yX3tcmGeTU7/p79BtCLS8IPZjQvtk7O8agi/TemUdUQJYCBSlnik3EFs079
NZI4qwj7B8hqM6Pqg8eEqBI8e+aPd9Sdi5lOHC+MzleyFzBVRSu9zKCjoKsamFIVCidbEwT9Xeov
71OdrnhyY7y0kUwi0pGMDmv6NVfiR/1WtbGl3u76e4xPtiVc3Dwd0eNT8l7rbW0b5M3JYyACSF9d
X2VYRTAeHFrW9U9izYDy3oqnnCNS5GPBdUD5ywv3OmV5JWs5mMjWk/4qCrScAUpfSZt87B8LNsV/
CK8Skw+OfUKWRvDKdpZETDqJ+RG0U2TMW0M7ODR3iHQlJQbf+0R3q8aN8AzqjHEvGL7Mqgn2dsq5
UA5ajBE/FrNvkm27ERTB/5IaNjnNmJxsxX7lRDt1jeefH8W8j+vsfNw4SXPNqSGXQnhqgTVJMgmR
/o2cQqapG/aTygltJbROWjAhymivStk3fUi/AgsyxkI4uZjNfBxk0MiZ3YPg7x3wboqLS/PqMaZc
8SF884NRGW9O1cqPGyt8r8MkoNMPh84EUc/VIFEXAV7FUMSc8LNodnVHVGJhNngsB4Lh7z93onhO
gjvSGkQpWYH/DQ2k3WGN0ZMdtdB6h3RnG7C+3gqLNvhMnrs9VTzOXv/wWIQymuIxQyTjUwGRbhc+
2/C44rS6+3WwemdZuCfvGs6Ee8nAQYseyXJZwHy3eEo+PDlZgeQsq+VhAZniZ3FgBZj/fBAAuKTq
wtBQn2QgJL8LJeVTpXBM9RvxsQ0K7H9V3HZaGARzBAG40urggK1IkGJjn/DyxFnGniKEXX9POlSl
+wh50rkTD2VG6Wrzq/86wS0eEhu2nQEzOu+miQBNkB/mTEJZdgcO5OhdqMAekiMy4M8PfTH9Rl4c
v2UeDTZqnImroD1No9fpwMw4jvSgDlTTs0jeuiU5Yw2Ngizh2V5HY5/q9FZyS69dTV3X2+Oyl8bt
LaKMn39qSw5vbwZOcE25/Zx17e03feoQzHWzZzjJV5xv6i1HStBByy/vfjWT+lLb9PpHC+1qRCvV
/r1zJvsdbOU6WnlMPqICADWAghgBBVWBK4VbJtfhHrr2o01URdU/B8ETpUhjVPd8qTKRtFX/+bt6
Z7vz4AJUJ9dB3sVKSawMlHcH3LRTywd3h4tYkeESHhRUcqetjR/WqKiPBjsBUbnofyzOzAgiFwqx
oLtU8H+rF7P12UD2FIaxNLHuFx0U+Eove4lgJxJKDXCflnVTir2ZDQG80J/HHr9nCpxE6+cYXUZf
X+H0Qpog7PtwDfIB/gMbjJfRFxdDmueK9tJPkfZeyRVaiqtha7IlZuGLhsBDjWzc8817Twvr5Oa8
TNaVbM5Da0fUKociZDlAvL2ktawm3ULwxz/FmnYF3UR2vmw0ZsZVyBTxr+YCsgv2d9Cr+lX4y2DX
KskFy22Uy6HEIjabE5zlUrZHUkbe6gY3emelHBcfFzRKcYJYD15ULhYayd9Oh9rLHhO8FvSvmU4z
IQqzhvcr0GeD4JQdpAFjxFhs8IB9DyroorCOtcsJlaUntj9E8MINlCbsnEXSWf+yOhTaQ8Qzea3r
2HIa0VmZANuc6/+T15nCQN9wtGplyKJXn5Rrj0n4cu1azgMRTYV31tYANkD0rk1K3VavIv/vLF8B
xFs+tVNoki0cT63Y7BO7Ex/5tvxU2FPAVkiI0J2ZouEteRn/4Ncc5BMJjc0jSlfRPT1Zt1xfx8tf
rvISowm16vzSh7RnPZ+I/6yJXH/ncHLJWXNE4QkQ2GAE+d+VbmtbDkB6Ev4ma5oS8IBhVyBN28p6
pL6uvoMMMoElAgmyMpaMMyqfJ2u9Du1zwt83jfe9MfgwEQsY6OFcxWyPDt0DFdIvBtEOLNXKFeIw
Ae/N7qqjidVC0DDjxpHOaP+1FHoPJLLoH1jg1SR9+URq5XeMhsft1gIAKb9tbHr+p/rf2ZoxeQ5n
KAYTBmlq6j+MiLIZVb69UWPiutSBPxgQEs8m1ZooZORNnCzzTvV59IB28ptEUNNHCt1fVCCs/2W/
5G9tgrhj9hUrsDcZnJ7UxAfPkSzBWbPUkQRrDGjQ2ngj+1u7Ry2h9O2il6yz4qf5JQBVdSZsdAJT
/CF4LkfwMM9bXeTwkJ5qyz9yiT+D0FFzvUcTMTwAZ51aDZyj+N+zdb1bZYVsbAtPMXN6eQZusx3z
JlZ/ATXA5gpvMy2pbwMnJq4kLQxOMaeG8NvE4IMYrqmnDI1ixW8pwePxtAdEfKS9pBsstUnT4ygE
mBLaLUSefLYuEuK/eu0CNfwB5ctYsiWg4F9vzGXxDv/J895XFtwmWK+sCHgIfYq6QLl149q0yYit
YRaxKQ47kG65j0Vpro6wkCZxQduHN+CV0AQNJYYFrdR9MU3uETJuUirCCE7gKvJWYDh2L7Kw4tUS
U/U/3JzJZiu96Q5f9oWe1oo/7Az7hBhlBQBrvvBuM/hhxEJyJWQLM8lp138ne8rzN+Fwot1Zz0Qm
WnEacXiO1a14hTeM7EhYFez3jSzoulv6aGplpYiS+qsEmfxN5Wp4/IvYGUZ/QHEEw4yVWBTJpmUh
GBMH7RlGRwzycLRcY8SiWhZr9Ni6QNsRxBXMVIquqEXMML727STmt16NEMZnP6tyG12A4aniwrwQ
/zk2UG7zbzy+dnUo+OTSWHN+678aVkvIrxR2ENdZSOfxTHmyfxb+tqdqyTWbB14Mq/Ucu9SRk35i
VNmLI3pVAFCs9Hicn++iwclOKw2jVCGiAF4u9MW9p9cyfP9KK2xkxL9GlKJKo1yLTaiRBIX1XWxh
iWfGI7C1TyLwcMiorWXnzpFbBHZPcPTWEoBzsoQm9BlRRNaWLpNRPFrCxnNoX+7Y681uHaXqvs6T
uJ6KmD0Dh0ONr0xyqdyMXS4xQ/V+93WwWTGGqWxHUDeDs58ci72MI2K1w5g7TvjzC704pzMGZVBD
CS38st6+fbgdFQAhkD+M90l8ry5lcC2B07sNe8yZWPKpafPD1QyZI8tDmHdOWuZKD7wkOiRkRGYy
s6u3dzCI4IxDrYx84r/I34sVznm7qwEl3KUbAyAtDT5V4Yfi2TfHOdE5/az+yp5FSCHCYbz6AyvA
6yiX0KwGxXvBvErGsUBRp12bMSPuQpbSQB5Eu29cq86RB574yoz2yAx/B6vRiA89A+dw4LLwJ+ZO
CGvC6qyPuJL10h/50M4Q5O+zv466yRVEqsPoBxmoYXKapyzFjiRHYMotHWM36eFHM0O/nguzyikP
hnKT5LlO5BST8HpnlUSqhQhrJHYst282ZHXrz8PAhPqFcW1X0l1lM6nNVOQ/jZ3glZNEWyn82cOk
aj6Tx9rXieKhW8LGWmGv4Ai3VzQ9I7i4FKgfPHcNoY6OvwUzxmKwDU4+xUYA/5KiQJhDrwN23bFs
NNgLCWA3UzHkEPc1CfhqkhKkShrC8ZvQlXHFh5+1K8LuFENkfJ/hl/HkzcWqp+IuqY+IwfNr4ypE
HUdSZ7a5jJMPZOyE7fSG+aHKvDQ7jWgrTvMy+9eY5WQgp874L5Yd444lQgGXWRVQFZs2jkEXQkXT
/3NrgP4ngSQrDNpb8XFzmHPfA4BTzrZG4W7VfxcAdmnaigQJp1URx+LqiJTyCLKEQg8RRAGctf37
tmZzrog35VCnPb7jibiwFbklCAXPmDuQ9BiUjcTUIB8rTQg6Fl3QGm2IWRyzRQHHgLlrpuLWD6Eh
DINPWD+BZhcBZL0rUWYTy4Jm7abUczJjINVLAMjqMbkYM2rK1jiUS4dc0IxGOTr4WMgi3ttYenLc
8JbBB9jRHxmO4OTwwSuELmke3HwrbII3Xn7ty8G0wuIpfq3ScWP9VOybZ843B13ui/eMgkhRaBcv
0SVMlfzPvkiNrwMfTzWzDexLPSYv6mjGxE/nj47SubsUsW7gvQNhJZXb7TmJBFgAAsrAA2BsdKLK
n5+ebdO8aBkLiZIbR2H7V9BowRAt+WL/gY/I1lZu10kgDDis5vga+3H6Kxe2pFvO3gMxj7HRV02o
oY3fQ6dImAHR6sgno3N6dOhXVKPIGh8stxxoJerOleUh3klF1ez/qu6oPdeuCbxyVqcF7ESaUqVD
ZyOK4K4deHFkhpGG8Yv0AEvV26WtTEorQt4kNwnhuoStbrI575I2FDVIkFWl57mUI9gELvEHsLan
qSGMNalfnVLuxXOON+gZq9S/C7Jyw2Ri7NI5WQdrVSw12sU7+plvtz5vyftbaih0PrxMi5Zxcmr9
PyCGMrzGSBoZzUTsKMoKJXcWlc4Xbd3gDpXvxRVpwMigt8Ocnx7YbQillfQwUSNruOZRW7OA+OsJ
PslYZhuAQdE2Y6s2MUf/bUILzvmeSokfr8QRAlBetDoSkxR5/BWdp0YiMtFbQchDAGuv8yhotc8Q
lvaWO0yE2L+eDJ9fyWxCmAOEbr3JvC7AbAHCGCr4nV7sfKhkJ+G+QIUaM6ekby1hc++DHNNAArlm
bDWG7P9+f8+qEkwCHBGBVVA7/XWk/073Y8RNikwykjURysn5G3aoAJXCDiGSgz0uaYb0Ha7Kd/xw
lbQBRQVUUJAJcO7d5EYO2lbEWreOD/KLrgb3Sdrw2gieR2EzYbfk7zGK8d9De+NeJKe7Tqx2IXdu
Ti/igCZRiH4hKx4GrBGAkWnEOPqOvMLtfDBw3WnNguEBYjP/heusQprNC/ENzFgz34lhMeVsK+BL
sn6JNZzcmTELYmJHko9CeQbskCKr1lOTYR7Qct7NMfllvO+w6wcEXOyV7+SqDe1LF7xLdB/avjvI
VGOfEuAtYh2jBvqjb1PEiRMu3JpmXwQvYNpLs7WpkMQ+f+O1bb50KThtLrHT/ep0XbEzSkevgCb7
PRwJIY4tV9qNHXV5WsnZAX8RwboSK3IGrDVSlB0lq+PilVcZpPkuxX66I283+915dTW3VPjw2QLX
2aVe3uz1W9MhiDbTxb7uzlnN6t/UOxtqbEcvx0JqihunvDmYb0PuJXdv7H2cx79LzbXD8sZIu0QG
mK9ssITBP1xu0lFRVG+T1zevoX4cm/4JZLVy77F3KtDQNYBhxMjsHdneJUNE/PlnxCzBialVl4BA
kaH9BHGhqLGinllAGtZDareXuOGphqu5P5JSwnEBNPsfrBzVv0fOcu0O4yJFk0NUP5VbfIHnsO+L
tGzMOVQAZgS2o7I62vbRGMD7hUZuBhE/9CGspd2RnAH2wbgLVUNIfF0GUIkUTdKmFbDtEHCkzS4U
/VZ58aUpF4/joLjmWrz+eCR+rlouz+7yoBapE+FXvnluO7MRB29ihD/uKbeYognVkVO8568AgVhm
A2G4/ohjUm04guDlEU37FfnjXYIM0Y0ipy5BmQSjluL6hZRh7YPLHpAlwoaqqCdON68ac2Zj7Yvm
FstzJHmrn9b0salUSUv7aTUCD9KMdj5UhpK2Cm6cwkM+DmA9yljc11nhHL+0wuvRJYuYmb5CbP7K
skEL38yu7t7RPF2pmyya4/eAurXhKBytI8fiOf1RZMoMrhf0RavFfzs+orwjUOGaU/w0mjLzV4ss
Um8lC9xaVxlE0GRkS2e2e4GpLlDkamJyQk8LyahuVbAXH5x6HpOAk1pe113ewH7qFe2ic9Q/pBbw
SLUaROQAuuJXaWi5mIaRcdao9pm++xHos47f72B4Rg3k71mJBhderg8kY2f5UsuYp2sWy+isBr7F
7UIJyciTk8IyTb1BDExZdQu4vizv18oBCyE9TVcHE9LDbBoj3CsAkKu4VS070RpyJIQYxl5MYscV
D1E+WSw2exJSy1DIjUxRn0AQCsg9h1chkc1u1D6KXCYfKiPNKHbbyCjeegXawsSUskstguA3fgko
urAAzOY47I4c8IgiK9jPc3yhFrWax70fU47Oc+aGMhsotfBYSMi2LFQqhXCYgEwLB8jwJct7iiqU
jWrS0XbVZbe9KRmdRMa+W+n8hfCjX/N54QpuMRsdjqFuLqjp7QESRMCOuohbSPaT6j1dNiOwu3iw
8d5vgIYdk5TXfCXQxOV3buPKstvE8ikDQNbOsiUeUMVzxu72acxtWei/06KAeBH1vZNgXAQK4gEu
DTRTH+4Ap1mLTkSbRfx/ZBLQOsgWwjazg79XcODJ5bONz0xyhzQ2KNHnn37vQu7iO0fyOsVbHBun
PQwjsowtticiKbMd1kVBGr1qfSg1iP7x2xGYWNrNf7E4b8uhG+NL87n1VTX9fJ0vgGuGar8LyyDl
ptIwrmznN4XVyxlqmtAfzBDiszPaFttdaQecwE019GySsdUseh4W6l+mC5wWd6tNttc67HkDNPf5
sy2jebmVZGEnL8/CPiwXwfLgwkAI7KHAB/GOO+TL1sQJfAqutN58tPYkug8lrXEXgom8zWl5HW+9
5MhLzNwRJyYjFtfOabkFrQNwAOTlhKj9gnUMjCIutEaVoU0mQE1qQSuHeCzn8z/eeW5qmDAH9reX
Kz/1NVjlYa1DbjWrSem38kl4EEn7aYcKIntvuffAhWDfsuVlkGA92Ufs3LN03yWlHYuvTSqwtC4e
chQJq1VjigsZRpUbEF3jVGWtgjRxHdqzPDAxkwOD4uAf10IxQiSfBDwByGr87pUE05bRfPHmGz0c
LguWkcXTREUXTFoWvqMU4SgRu2tNexub0hDYocpvGTc3uzIUzcADXUkcGbXNoxvV57ipPR2keySc
RC2E/JATh5sgtuEanPUAmO9TIhK4C60POhSlhAiDVMVAafqqkh4KCrEmhi3kK92Vbmy8hUQmxYEY
tKD2OS7zbDyP3EmILIX3krvtQ1tq5cZepzbIianeyF6AK1mblNiVTSh8uT/QQL6kcOHGFnS86z1Q
uax53PQLaPblBNoOg0ba9scjBMKIoP79tilyr2KTTHYOQJNIh+I9fwL5k2Nt94n4L0nHa0mDPELM
o8W4XVjbk+5bOJVzRIAReuA06/XUkmZHo4orpTXfyllo+HmzPPU+tXRHttgxvJpa0LM79zaM4qnA
YQJZLeHc/HFvvxWliSG+pBuu6Wm0sQAvcwvqMJitKZVu1fm+yuMO08smFEPFZxvcPaqMXYl4pwfD
za4To7JYJI02Ao759NCakWEmrx8DdIC9cuGHmSnVZsc6zctO8msdEU+paeAX3+ehJCp9MZibc6pA
fs4rIbRLbjc0+Hq5yTDEFJ9vx6uRP4YcJpYr1/n2Mw+bjcArCB8azONBtm7O4OFDT7avVMu6om33
lJmqmWaUXiitT3ILBA6Vpmq0B++oBBtUxRDAgNN6CXYGtiliUk1UfKvB2H9WG+qlCNuiSUoEIk/g
mpiT8cGuAF3IwaolIPfGkYRd427Zr7gSm5aCsy2jJ6slB04+Sz1XLUaSSVKB59Yndh/pZHHjTDmF
sElXSQNJuV7C+m8RjGNoB/tcTAjdTQYLp0AG5jFSrP8v+UodiFWZUjdHhajcoKgzht8yhbG2XaIP
tRE5Y2JEA9ykhKoMN+jnzN4HMAobJDNm/gMNl16ZqB2nvPw+KBQIhgwN7/493IDAQpEnqmZq8AAK
cCManVHV4vI3U/JyCZVVi4FiY64UFejUuYZejARRB4vPtNbXSB5jDLBBofToylXLykFIsmqLO/ey
ZubmFmR4yfYzbSgDC4ReWl5zlQIjr6v6L/1jGL+ZOB88P9k+njsmRk0N4xhzRSsM/VG/yrK/kioR
DG+QQAWkeMnmjif51Zaxf9HCrRy0BPA545+fqQ6q3B6q0cu37ZJsS0IxlinbQBoA2zyjLQzhv2ZQ
HSAKi28PbhXVrMN2eM5e+ScvIaIbEI/Hb1SXkMK9/eWpIRvHkKGDavV175fY/2Ccf7hOu9H4qbBw
5g02qSB+21B+2iTzbEpkHwhWbAqCML2YhyJ2KNBZttr/7EZeXDPtYOO5Afec2ajp9Vsh2gdUgWnA
QGeVwuEvay6kVDYDdYrgPdUm+E0Gr4T7fYL/OILLzxIgIk+kDGY/Njbjl1TQgZBN0vchz60j971L
PoWSaFP4mIc+qSZ/6Wyhgs0lmNyu0IPsyjgQwnNCn86z7avWTd6mkuqhoHQOTvFqh6J1v3QNbd/o
ZiYYSr1gG3F0rTLNbfhHaz55+SirxcccSYnB2QwtCu9CtJF8wazk4X9/jcC61c07smU9lXevELg5
g9rSjlgojfgsthuZ7ibqojSium+z7Pg1nDuOyWQSnV1kQCmZBVEg53EMjlTFp0KaOoHgWP9jBEyq
pFwHACp69+p5dJ4qjkGnMOiVnOaB/1nQ1c+QeoShOoLbmj+8u8JpTk/hPrFTjPISMGWEeflDRRvJ
y3Ew3MBMCCO5E1X6QXoHe7SLKbCktXOyi+uIlddXnci8Z4pseGJOKpf8fe7WayPo+u92CYXT13Ut
gTNZaKhy2xrIFi7dymXkc0G/uOazN/GqF7OTJ1trh3pBWa/FNEyMP+e2WMBTIgSni9j9Rk46c+ON
UEX3CasW9W5j+1mIKnKld5CBONwxCiMjWP2Uok4Xt8U/0oTRL1/gQgISVaeaj97viiwtCIN2X2PA
TwWmDL7Q0N+xjtapLZEUTr56IAKnW5LlArxqqw4kip00ccvMYTpH2GVEqKHHVSJSNeXZBYKe+emf
YbN9H424yc+6UEg+czqKj0S85VMro2vEFiW8YD5yKX4llu28RAsKLoYbt5hGY6bRBw8B/nqJZaLD
XzUmgDsM/nQBath6jnMVDKtEe4NgQoJtwljaiX9VZ5qe5bnw6Tlrp9ysByJZp/TOr7jGIq+t/+U6
uq5T3MSmkTtgxfBhmFk5uEA2kbpBjlOq3qj3YOFI2f49cEvRe5eyjnbyFAQZfBVUWWBd5uAdvfJS
BohTazzVU/XttZfCgrjNv4F1aXfbM2O6KjjR/uO4SbLb8C2Al3rB2fAH0paABcxcDL3rb6hN3nz9
ZsSsi0LRshn18EgSGD3a71UvCZCyHYBd804b7JGrQElOCvm0Ash7B+TiYqMJ+kmmbGRYVIRZ/Wzw
d2xzGOwZeE90zdsS3GkXUyNUn9/D7HZ+xzi9RK7mM0Xljqum29VHmaJxms0DsLOd4YQgW4EF+RX4
gyjjRkug6PpNbeMy4CgiBl3igI+W72LLfyIfkV0bfm6Wf/G6h1Va+p8BYlNZLA44ES0EZ2Hsfdvn
sTMzPCHxddudG2MeHqCITFy2kP79VlPUh/zgDMRxGlDaPVDQ/ER2F/69jSjAj3hfMmKxtI4rVg28
OIHvpsM5UiY/lzhynV9VJeiWgMPWBBrTRYps9Gh94eH+ZQ1fUi2tOtjV5O3INEMexHJmd0QFYrQx
eTx4OBlqH7fG++rF9DCxcxudetl1+CG45wQ00HWSyMXSCEBNWkJJEN+FTdmdUUY6bJ6ywG/wYCBJ
LzWvHja3WtqFxp9lUetv5KqNjxPSpJOfTTMA0RgfwcuvrYPlOcbzzxWFDixgrQMOQgx6RMa9GOVT
PLliP2EJ4nZxQP5iV0xAQfNwqa3JVIPi0DymVqI0wQD7qKlZXA4G1hEOMhWT8LKkSWL72aLxfjgI
2MlnIeoDff2AfC+a6tNrP7hs6GIW0KGA7aSQk+4ooX9sf1JIqiTks0OYP3x/iFIQeMBZTa5HCTzS
J7fKGw6AkB76QrjYFMpHMsOMC+AUOzkMwtGrW+V+jfcfWgo8sAAT+0RJ4aVlSRlj+NSC48FKIEtW
XcLCIakTcVJZSkfijmlx9NtQJapFDTbm1/nN7zl3KZFlwvOcYzZk7DpsTdbd1jEsjHl2KbdlLld/
2FWmHNIPb38Q+p7fZR4SZE8zqviTKeHVE4JGqNTTBFuHnur2b+alKLbBOXUVrCh9ll9wPPfX3Gqr
JNORzMnF/EN8zJ6QxjeQ86d79nf+xFFW0OGxUjqyZLRGXp+zoEsCtkUiBUAbqWfETyB8NQx5/Q5B
tJiaF2PYdrGY1uYZIxO/N+AgFZfwszlsFv/mb/6UyUVpBPGMqfw5WeIFjxak9AURkHzMOlfUeA+R
bVKUCRVQ3r/223C1vbIz95A+hIoHRlpdwdYZmqJdPG7ejFCdgOd0VPlm6mkfEOpDZlAxFfb49Noy
PtFwJAk59u57PsjGp3rvFw80ARzWhV12SgnNewJPL7NcA6wwVjVGCyKiZr1xbgF67jMtwZ/5Vl/k
d76iNi31TiN94FCxoVH06EEs1wKj6K8ctCDmmFLqHuy6rLcRnpo0xa6KGK3BGR/vGX5g1dMxwDWl
sSWeOnj7YiBILJ2vHMGZiaZmnsGAnpBXi56VmeevB+wFkz2cgLf/atc5TUtIIxmUUnesGGsZCQWC
syQNl1T2b+s4LfvkJzqlqBIo+aQcubZ65P0ULpLVp5EPpc5RAXz7UZCxB40psY00Q25HqtGstJQF
5P6LLbVjWh8fjA2krEy+hB3uRmW77XqspmA5z9Dv0vkcKUiOl9TcsP64pBPxYIPAsMjVWryxLrcD
jBm54rVxQgurvJv6YZ4p8BtQwYA/HmHgtqOJpgdfhPVFcO5AbK/98QkPJrFkwfbxL35aLWRe2+f3
+IARCtF+J31RpIiiUfHG0fZIbrjcqEdl8eq4NHXw0Y4CsFxWLCs37iF3NC6RIOOJPghqEe72m3xO
yiJzuBR+Bft1YgOiQIje6/KUg9TrIY7kCzKPIozZZaxjWuRgZQvohbh/GzM8QatU2bUHMvqVpdUy
i3B/OynqLGSt4F48/cZ49rLd8sBqvmZ8jMx+zUtMmKKz8mrySeVN6MgWwIa43sxf6ytupzKmzAW3
K1k2kGEagovbYOdq8jK1Prx7Q3betEDOHOhhMPveWFjCKSI8CNuGw+MNaXK7lrRGjrp4ta6dHdzD
bqh5kxK2EnhTziIxUQvD6d8SSZo+9G0EAEvP6SL7FQkKkSmjKqi0Sb1pzusTOHXUNjKA1GtHNZYz
3lyql71IrivFGRZHTFF4FedHT6AocobZ9zwnTMZBYiALei2r37Hdww9lKtvGOOzmxZYLPkWBTrAV
Qo6UzIYIwLVsDyZff442E/vMqOUQwzO9yZ6/Rd6xLqtdrLP/JOV3vCnVF48GAkwDwvKLFkB3g5tf
81TqGX1I1sK90qN+QtFCC/gFoyNQ1c8Z/2Ctz1FGA1MQIB2PjCJGtxwNm79wughIsN20SlxhxYzP
8l7+CDl/nXYpvCz0Nax6JDElJ3RszhZGB9IGq7GoVBHqDHvaWv3kJdr0n2iSfQJIkaD2Im8+Guzo
h3jWvG3G5yqSdqIh2azbAfu+B8JytL2XNSSkLuNfeybtvx9p5kXfM1kE34WlWggQ8GyWnrZ4Tlm0
O+eHZQpdSDRGaxjy4HwDlHVZzEBMl6hIwPJeK/8rtqO8Xj0aYfVJiQ5NpAM+DzhaygbWmor1bcN0
otTA8Xs1NhkPpS3KabjTPMnyhwqorOuQ8iN4HnqXVA9k8Ms6thhFbETcmT9Vyl5k46o5OdD/8R26
uYhcRH/Lq6lwr8ZS/LTQqPKgZU10CmqoBlM/IDKI4VORti+3cNDluAm1TXRzbad+VyGfnQSI9k+x
w9YxhprUZ9E0zz5QH1EcH3iH0LPx9CrCcfNLhes6ye+9gfqehDImEfi2+pOvaeEIu1S0ga6uJ6YG
04fTNd2nL/pVpsSYjbuqUv9GropRxryWxJ3DtynWm/deBEHE5WKCG1MS/19gbTzearYpI5Kg7yyP
NUOjD3qtf4sMDKzjbdHzIHmiB9o8ifk9Q86PRhA7tXYxHr6L5F8KktptQ0WhNUq6pE0EMTSjZ5tv
Tq8S3x3gcYe3oQSueuBRm3nEgjcTvcfrLJiIC9PvX1uYDJGN3NL86libIsx4mEarKQCsfoQm5siK
9FHCVzD2jKlDn0gLrvH14uFaZV8Kc67xL3pFL+q4VqDgiQNkb3k5TnPADvnuSHpPHFix6iXUr//L
SINSjhxGw0F7s97mKDOBNCkzHIBtVGC4jJShv7fUUwqCpf0sdoPpP6oQUaPrp86JUzOhAD3v27XG
eUcThG1TC7jsm/6Ad2ppb2cL6NHkkvVoMrcblqZSqMNtz+42Plwgok3YxLLB+INfYOqHTch0d7uz
Lvypf9+cx5QGzL4p2bUQfUKywiQuFc+9IrjJQk94SIJ4+C4DmnxEVaLrRfNnEiUhMXIIOrL6ukbf
2oTEjYslEZvSZPvl44YZtanip/8k+ZCEjStSbu5dSzhRA0IT04BiQJofSpYH7pykANmKf9StMB4C
OhNZAbEtruBscvVh0b2mUVRfL97dsP9BR2MM9x5X674DL3isyhNcjR2rMo1kUud8AFAuOmFFOeFz
78oN8qIea3bzJi6h48euSqEtVLgXbPHmxIzNG3boDn7uvyqxT7dXX0nQTW2ldkrnYf2GgTLQJMw5
j+WhWsXOFJ7PidhB6kebTzICrNRXOe4ZQ0zBgJtN+WsOAuXrvdR3cU/6HnnRW9es6EWwbIOXso0s
rtOXA1euSKY5cIX4Vo5+0K7d0JcumDpZ/V13c4+ZrX1YU0Q1q7uh4cbHhlhzq3UXC0DwstrfHIcf
o1DtUPEcg97xUx1IhFd1w+dmyEhH170fLLoA3MUD6t641pz3C4XE/K3mM3d3ydxSmd+PHQv+qkHj
DJ8LdqCSbY023/Rm9yqRn4JVbEoWU28lfoO6pvaMlO1aIjAT2t3+cuGDekPXUtqtUyBx5XLek+SM
RfqI6cgVp1wUMfDEvkifR0EHNNpzQu2VfJeSSbjUS4oCX3T6kFEHypFyVqHXxI3MFAOTAPEC4DKo
vnymx6QDDRDdOKpnSVNwZdq/uXVmUI9Qo9F7EuRA472DVvG5AaEKnrehlw0r7Zgmlg5yLKoI5gJk
3DAv8IAB5q6VMiye9nhB56ufk4rckhbe/50rIowpuwA+9/lDoui1t7IjPlpHYCIGvsixj67LmsCd
8dgwh6+l1BxD6z7XJEENA2XsGWgUotNSfXdNBp5u5/lDIl8apsFs0LR7Yu5Ngb4Hk/tfCLdcvco8
VIQUm8+mhYCXjXcqlZhu00Wg0bnxLa8HKy4NlE8G8OVi2c7MMvPlhwN3i4w5iVkFj4sh3skm8o0f
fqIMDAidM2yYXExPI4tecqmPx+hBd0opB3AGDQM6Wf7NxdU6GQsmRQqekw6jBjzrFqTFm/CnemxT
zxF/0I+sRW4w+Eko6wiEOiOnUdZ9KIs7TR5dintwPLBGg9TDi0m8ESSPSEmfytfbJlqd6/opKBBE
+UkLZzfNYvToqGuhwNTlT3cA05iYzcvb8H2DBOJLOhC4t3sXkK6H4FAy+i2ipvJADMHIS7Uo9ObH
sDLvUkkDHa5Ttwzfc0KhnBsphxfRpj45AXU0gKFXUgyjs7z8B4MEIzrido9hzbGS3sIl6eoGjRpS
kFtU9t+KxsD2Wu2ffGj3bwBHtXB3EebTWndsnMpF9kMIQCkXO78ivQfFxRrJnRRPJk8L5GqegLAm
oF5F/k9EViDi0Y/+WkYfaq/0KQ4yGOO5ZhI66XkQl9G42QwSSKwYyr1ot0r+7aqA/vaSir80z/+/
bO+GE0HpuRJk+VaQ2ptKxgP4egW3c/YCG3rlSv9CKB4uHK/dJXUDQ8FRX1hYtXhVM76ZzUW1sMXe
KrsMGFbvMdmEZxahEVBjDnhH9LkTeTGGWk8VknAM/R1S75/qBLkqeU16MIja59rBgIIf6RwOqFma
hFmiy4v97wlSTCVyP5r8Ne8/sH6yh8p+atdL3LFeHMm7rIUvIaOmS29Jn7bXya2zrYGQaoVJkQ3p
T/APvfdGuWyi5azIG/xrA2lCAeAeCl9rBzXQLukEt1ThntHuzGSqZR+SKbsUoLLXh2vVjMfsI4Nf
K4HtjOC8GH+EGj879VxTbg3cHUr7wYfGeOYtc0Bw1Dw3dmaeEz56fnBJkQwxuOWd+M9uw3FCDgPK
75swpWWrbdNaPl7s6tUoN6N0U/G/H+JoqN9VvMGOf/pRJCey1hzmxtgiKRe9OCox2pM3mUsPKaaR
E24hc5k0SkGaGM/BKXs0SPHpy6HuEkNsl3PUieqTA/d2S0mICJP1dYvwE0Tv+M0LNLMru9CqXAfh
APXa98o96QdCL7bfCzvA2itpKp/NxP/jW4mBlsYrXk7PC7kcl0yCFao5AGj0R75/AgLGIkx+yLJn
QL8FZUATxBCEJizFZQkG1PPeFAEde1BzYHtQs4zKrwwAHp5Xky+Wji4sI86mQbG9GhvFI2Ae/eRv
55sRbzGYzZD4zsbbQon2Xa2WTT6A8VjSc3Et6QXH0GZIc5T17+0mrELY7KpPwGLgkntFZyFZ8g5O
4VTbp3jKcLmnF6WKW7ywP0H6YV6yQP+TE7z4Lml6TjqXqC/F4ljy98xbyRo5drP5i4SW7pr1dnai
BycB+vbkpGBpAK6mQ+Yt/UU6KkTcDywWT5G2DoujHmH2cN+Uif0TJ1WaqgV9aHqcLVB0OC8K8gmi
Ep37PhpcHUqEwZvael6k6CREkhVHaHYfBwJ6cscYLxONQ0OjsRumre9TU+bgb+xvF6nEkkyUv530
jjKawzNci5ojOrDZfM1BJBZAmQC2P/GK8NVI67CSNI6rE9zff/ft6Fyod76yE4goAMRC+V5wXkXG
RoMkusdI0wNNeXjU891M5tdJ24T+GSfURxzfg07xU7MwAd90rGfCad7rc4VL/o8KckrcC1XLBzEH
YeaJuFFu19CzSdS/8fetZIBPTFzNNdSXekSS9v4PvinXMGjr6zZSoTX03fDcsv+Xf25sXuA01UKa
S9j03x1apRNR4Y8eG6JPjmjC6d8uo9BsgpA4j3NWO3qT5w0xMh03HQhuuJ2nmxDwVnabGXHyGlmt
2Gjp56v7/obXDJCuOkl+F3Kyl1NgxfgwIPT5N40p2+qGehT8WJtOnQi8YrgphE1Z4e22HTFt+suu
6Hcn38q4znuWLSH2bjl66fV0syhJOFpczJRa2Q/ysYlT67zGMOuLTrYESCtgkdLZhZ28MXYcYoZy
+Ng+LFdXtm6h2uKbAXWbs6MwE3PoAgoF8mGoDwi4ikgKchW3urCDBk7+1TRA5A2HHKaulcTlFJV5
z49/HTWp0Z0YTgvMjC0EPTer4q/hcYiuweTwkPV4qaKNlb4RNJe2ymOk8N0mJagTge3z3jY82nUC
c0g2UWbereE8ON589+cPNW+S3GjGDFqG8xYMAlPi5R/Mnrbg0XqoHk3wXqX/OYYaDzF1kLqPquuf
rcGvKhLmZlAjmOZ2MsW7oMMLRZ2Butig6+qocVyT4dIor83kxIIEO2B68JvRVi/USrizCq5B3KS5
ZzjFr4jhYa63r8iog4JKTt9RK4/2GKCxU8YUevrxUd/v+5Tx3FWuvkPvZxUI724q6BhuhC1i+y4o
CbKwBhZpIP4DrjXJdZhZyzqrPXjI/WFLxMR6DiYqFPQ5JQS4MSTmg44iJN+lASTTczzcdm3Sumo0
uR3OnnY7uZ7oK62mg6DFD8dE8BXhhrFr1x2Zr34a/VAytBJrgz7NLZm+2rwbO2W+VM25+eSPjfj5
n1Ld9MPYWy3vSYtrKN0zBBCcsavKHLJtHCvTgpZSUrhO0hAZm+CKqF/Mq6FSX2cu7D5sNJntNiC7
UFBlxff48UT8al1XNf4xTr7euBSSDuzxDSN94SYIyNp23fReGsBwuQZfw3sY3DbPkHKeYoCvH95w
o0Ixj/lj0duzJk2oBwOOM1Q4Usyn+HbQ3DpY08E4k6jId9LRRjXeJaHOMSAEFQl3bKvXkXDSaVbJ
3o2tRCmmRuFMrd/H3CeNEaQvebBj8a/PZapcGT/sm/p3NV+6EBuGqrf67CgccnpkcroWpdu6PeC2
K0jzTeSde3YRnMppp9MIEztdKAGC/yrOHInYmZN7s57TSEWVbEt51wVJYsus1jOnrHSOBZldqLY3
c5aVjJAMFJ188TeSlaLXeURdei+PPw6049hnOtbVUX1k4XvBKqm1MOCiE9HAHUqvl30kEzcikEXd
qAeJpvTt/cafqftEdw1K683JnLfY5Xv3wjDJ+ZWoBftqPKsIPE9fBI/aG3wLMZ7lBZIpq6Wm7uv0
zaXuj8zklu2Tj3ymLXMh0gkdvFmubQOFbdEDv4bI8Ra3F2BMHlyt8RwTwgGj++ylJ3/sbCx8KNfF
IKc8RHOpsquae1zdLF81rpZYoQiPTdG/xNZpGqGj+2jBPiZchQDMoDtSCDgTTStGC570mpCEvGrV
mSYkbVhqjNEaFwHxDXZuqGAbvAkJCVVDPiJIvDcGwkIHL7SAuKZ1jOz8SfCpr4HOiJen4Fslrl7V
TZ4s8nRBcnrY5V/hyMhoKKky9zUyVaw6QlHrcDbU5trhcXGWs9SVt4MsunOBUy68ZSW389zraBEs
pbVUfrpDBlXrwKoj3e8YkTBC4oBrDIMe4h5N7AmjUncLFRJYvnoGEHNsYxdEONEjjz8/5fjyZRDu
1WoegT/af7b7VvjdNNqjgNc7yGqPUp530LAq5NbDXlPjwUkhuzh+qrZDCNgCfY3xB+ag8zbS2eU2
+FC3lj3e7E7w4Zk3APRnGNoWkZwmzjvCin7n6yCgG0v7AMgS7CsnNHX+SGy2Ls1ClYHBgTVOG9hh
iqxn8FswGC35UYS20PcFZJ81gdR+UMoosV3K07/+T2VDbVfy3ti9iVdWsNssdQW7wSsJ+Somu9uj
UtizrIHOuuXLXC8mqcVF5G6YZQHt15k0E3vX/Za9hkbln0idgE279iIPJgy2gAQ3OsXUiKym+Yve
O3iyo/ZfTxFbhqs/WMk7E02mEAhRyTf29vtSVCYLVGGwO3oqT+k+zR0fvJRD3O+pHDUNW6Rbcrzp
8gTL9t+c1eBpKSZGbmeC6KOj2kviv+EP5jlboZHcEzyP9rg4bccRF3Q47O1cZTv9MqlXPMDQXwpF
aIsvNqmeaIxo80TNb27249H4pZZpXxOmdSxHu9sEldAiyt8NMnnYqMYh8qUk1nX/AgN8XaVBQ7Mb
os7eiTlR0d6cfqXKIxyZBZONP8vI2vWMw8W/Zf5NBh7sfpKyW5f8owRJZ2fehRfILjJ2M+S73xM/
txUk+EVhlg4ihiJtT/NFBohaPLvzGMx2oaMimXbtZMRA4E97LBlRG6O8Mbt2JdQGGoFJHN4eZI5B
bx5NG71UTF7tT4IZy9d0s+NgFP0Oo76My+17uZVJQKZqcOXhVTJhNtMhKPlsDoTJoFktHAr5Juld
lAf5vmxb5kAJjMJ4Z2QRnil7AG/XmsL4mapfdJ0r+YZn9KG7pOW8bzXFVtkS4GVByL7pH2MCkdO+
fHEkSB78F/Gx0HrnXwT+G11Y4LZ5+OX2lVuB0illnC0L1MUIpOE5Wd28ers21PMvn3txlkgUY3aM
gPdaYI2gsg7RHLeuE6D0DbxElbAEfHQgSF3yO095K2PBlBMnejAODMS8w1XTnkiqR/SH1YLJ/37F
A1BVCqIL2YIwydAMrAtEBGHTQOANcqP0ZJDUa/3ye9VQ4Gw4h4qRA0SnNCGCMth9mjGfvDw2dcsM
yXaGSf6VEksvXO3vzG1KTZujmX5Y6kEIjpLDpnLO2UrRYRiXFTORlhzBxw0YtXgpt9Y7eFuwRG1f
LmCsTIEQv+/pMYxhiV/dd9T9/uT/hlqCCap7PWLd3sL+eZ6YNNYItYxkMUG3A6RBG6nJ0SxxlBU9
kv3NAH34m7fdqYFBwYIM+jgQ+IRDUj9/IAdFIkwHN1LKNXoX/kIA9B8sNC1tlSkBq3ZXH7PBWbNa
16yISuze+6LFtjFx+R1TjjWEF0/u586vVcyYgG4vrEAKcP8v2qF5ThycfFFRt4Ir9JXz/hR9RXd/
Y5CZUahg1aXpfmb04dO1FT4XUp6e5Za7hcH4z2zU8PYle0CGT8GouM2/1cknSvqt13tVAW8BQ0Rh
sAEEZxuz8pc62GplXXPSZJWQGbfJDeZtm6tsJee1gVs2jiiqKqyNPjVRjV/PXBlD2vfH77iaar+C
oR0dmh9vVy/BlZQ84iCLMEgc7MqPfsppejspjqV/ZSU/FNX+kceK0Uap6S+pcFGuubhUUxU9rZ9E
0TGe6CJQngxPc4UPpKAQdD/Ro6iM+IjT6F9OcOmz8+jERlwGDaInldFhYOsiXOj4MXssbEXwnpcl
ZyCEHdPvVAS188YLHkJfCTnJbwHknZF+peUHouOJBcC+2Rs0+lm1lATUzPZypGF3yBsth6dW3rVJ
ZbKGNmnM/wpyVbG8k3XGxF6iEZTqUvUbanccrVV+a27RR2tJbhBBrzeC+9CsGA+dPgg4XcQ4R9xD
pNvM5WchgW0p5PKmS3Yg8UxcatXc1I+6Tw9E/cJ385cuqEc0PNtnXbmMJFqQrg5RzOaQ0qt+wGqe
HCR6jFy9TlHnkmnA/kLU1TelIq0vltidRpEd2ZlsUNjg6Ei3HvaYcDOjpqGk929YmbdjkfYXy7y4
m0B8aj+uooPEt8UYbG4pNo8t9oOECXtOOKQ6bE0X/fpKcd8xGINhTzv0iyfl09uRY9KJXPJYzwB0
XX9DY4LpQHHyuXdi0UzqKqTaDD5LUl8jGg+boHQDmy+RkHRltWwxaReig31uS4SjE0cL1fXmIvXi
y0vEqi74kF8bcqQJyPM53UO+7MeZk6dO5/DrbDfooiuhxd46L72OjQS2ZVGVLqMSOpyXteC87Col
qxWrLNViIVvzIB6fvU0heN4zn/sI5d0HWD6BUetnb77n1awMRDXLABbuoytgoalLExSk7Bu23Zge
ho+obiCh6OSSy9myqe3+B5jq+ac7VbTDbimChvLEbRX01c4bbpBDB2oTOY35iL8yMN3YmdfJHJ8L
FHURYiuZAUBJKkfHwi3h9XVknuS4KAGFsOHGkDO8T+emFDk+sncSmB6Hu2qh2pOw4GGHSrg3+87T
ADVAhWulTKFYQfAgJNei44wqFGGt5qkE7SVRfpAUZdtgChNy/yw6dqnjM7SukA5bLHop0pMqeE1x
LdBsdniDxYMo/efpumh9IriH9sua0NsK/kR5Z621Zu98PaxWNWuC3titytZ3D4ZoCwWW1JZXXq2G
YUdtW12JKcIJflQtu340HBqQAqgTyMqFKxBwjulsRXqMl9HCHkLd6FbW9kWgrcvN1tcUbodZncCn
yF0BXR5FE3iYSX+2VtjOAGu8WyDyX4YVRG2j3BKVeLmma6IFm47/Enljh0lzqkN3/sK/x6c/NsCj
joSNclVdIIEMiPkp/wqfZ1mtBz7Bc2GgK+c3KVsnK6u2aG+cAE52/ndxjj9A58y3ayjrgKKA5CGD
FKn0oFdXdt1iRX/QOboNv1jJ4lxTQuQ8ujMTg4M54sDvYoI5wFwJl9DwB1OjM9H/JitUBeqwdKgw
AaF6tWpyi50tCWGJSH3nsMCCw7ytVSzpPajr7PIc8E0y9avjl+voIOlao/BWrKuILOFaxD7lhbAw
FTaN3l7vmosDKahE/oP4yyNeYEghEJtRkX8HYwC/q0FCBhhqqzxlJuWHGCqmMXyjA0blThYhyG5o
ZFPFFrgl3d4PSY6TG3pZvBh+GCxFrLAMkI6svL7IHKosjUQrv5IUJPvjkbN0G2W03rR1P7zxOQx5
+1XenGz2Qjbw332bPQraoWz7GvO1C7dvnccF6ghmmAOn5UXf+EdQoPLVcEmIr9AAr01kjxZR87jz
vqjgRlZ0fgiAHGgS3eku53uJvpswwc+S2cSxHnjkfjmIJ9l3Gg11B7WK8/9/vjltBFsQCB9dwtHJ
sJuw5KPv13lsPvyfex751NGXngm+4dHAtC3i7jlqMc5ggVrdFh8oZO3J0VM/m9d/75w+PgxmHOkB
bv2jNEG7V7Cdg/mim5AINqRvSfhrKiqOFkWAFOesM7Zv6Rky6xGWQHAYc2VJCV9nniRo3EmAaQCg
MOTkr0AH4go92Plxq08U6x+TCZs7ViDk41pW5kWDimNjINtXj+SwNNnjIWA03hDZ3QqwI62ljL6Q
8jzPzmiVX4WTA4DNQf8WYom+7wTCiieeFbV9KSXYUYdth5mTII740mdQvOSa8g4uugCfz/++ROzg
N/m0KvdPy5xRsBNTkW+l085B4g0drkenl0qC6kKGGoufbg1cSSa74yC8ub1oc6Au7MkDRobKdyts
bB6dzWYNhg1XAI0MyJ7K7GuplgqSneL1PfVRNbca/F457DCoHu/fXh33OlgMlI8huPot5pnR+1/i
8vHoVkqSA2cWZplND4d80RcoPpv2AIasrp0+Mglta4kLI+MLnxIRq4vhca3Khfs0HhRBusRL7rkA
GFkeywXff9Zgw5t4e2E2OqVQr9J5WgodiHXOyXOXYyTOHA+yktKdCP987mFFEcGYoIhrXQXOVYtO
7EqtkUzgnTvkn9981EZOnyHtUAPWf15lLPWdS5tcCfoqG06RpH/4sephUL2RK9OqwYvCiH16aO+V
uLYeZoRBSKa4fey/7Nx5jlMoVvq8kB3wMJXLVZJD8XHCbZxTDO5ma2clktLI70lEfa+OIRtQwNOA
xrlbTVVv563pWD/eA5k//orzOQPgyp3Em8lVsf34lgIl5904qx5RabMOT8QEfkoHxVvDRl3+w8T3
U3GHCJpI9Aa58YBCCXocne08GmoAx49oZNXbRZ76j7uc3/FJILhnoxLTlFebzahhf8x2C3UKEi7N
5tVtuyil2eIGVi0rudE+ENVva6M/CJiJ9frkGPgM645N+uzPgGWJiqoJwGcR4p1+cPBd3Ig707ai
Pg4bZoOZvTu5eCOBOBQXzJZmXjgKMwGvxQdJUzrsCnd/JGR69BWYkBOOIxxHPGTaMgg4vNOGkK0B
uTikBSWycHgT1dPdXBBmekTb8iS9Rt4scJygqqIUwVfGzHnQc5Lt5J7if/RKVat61EHQEdar0bwu
96WzCRc8sXTM6IZz5iYjg3FUabwkBxeogXrSkCKleK5gyhgj/uJMwOj9ov+ntsR5r+bqU0ZQuj4F
mrwTPXtOxYxt0+lYuJ+R2c0OVQFy9EJCybEPROU1GFojm29ql/YSwn02WEf7j1BJxglg3SGp9Cvd
y7ZjGDZoykqPdvahOj8grKbiufDY5duHgxjRRXIAMmEGUAxU+HQVjWdZbvPBGXxMEXJUZKv/HSGv
/obUKnFUXvNVGYHaMTVljqkiVmdJlh39XWRSe1Ns7RCwTxf/CAFNkYtD0zRsJKb70ZRCpib+A76n
glZJgXmeACiS8iSvsGL5nbdXJnYRfVcpp2sSGIQriCCe01BMdvrFg5Wc236IT5M1bkpgH+AQpfEJ
/lAcCJvGzgw2u6eLPUlTZAt2e57/8L71ZYXzK4L+10OWCsBG4RbJAMQtIEszmcoVoxg6H5SZqN79
3Hjk3K7CmMlGJ6qVK5fZHHcpWbj/D4H9MwhC7AFmQo7p9EOjYKBKfBQViOCU6D6yti0V2vzSq/va
d3jITeGLSY88vaynHZ/BRvAq8wfDZeMtqAJysAJLht09XJ/zL2ou5O/CV5cCjg8J1At7d9yPfO/5
JhYMXXYGsjUrJABf9olWu88TBL5Qlpyl3+Ub083thaqghxWO8MGQfG8yWxGRviwU5jzySit4iVew
2aspq2Qcy0DJCbI88JI6WVDIj73+b0jSUHxWGwA7aLP21LN6ouxF8yvUfEW7MgNSrB6fqsP9uRaP
SXgk/jQLyYbnb+sTTMXugvP2ak94MyAwllfkxPM7DsOUASYoTGDFj3eHNZTLGDVqMkq4hdbEDfra
1MFwNgmcUe/IVOxNbBG10KUxWK1DY0GvlR9mA4MUmD+f/m/WiE/+1umQJVQVxXXjM+hX46cUzRoK
Beg9PO3Dps7VYon0oBx+rdAFriuT0Mezybn25YFk0mz5Ok2N6xrL70V/EUS+caaJwrDdCYrtpIlN
w0WJ+gnPnNStNd9trwdwvE5qhC9bP2+N/TG7d+f9fdz6K+YUjC6m3yPtX9LxF9A415hBO2wSyHTc
m6b4njN5kMk3r4/kxy8aF7/SS+BDLZKgT0WQW4gQFbn0jMngiDvaQc1cIsj3yao+tqH3AbWhG62u
6rz9tJv9UjtQqw8lhOCnWJp4Yj8tl+xR6NouQzBoIue2J8zR4N7WIsoLKynt5nXgoMU2fLLuJNSd
gMMM2uRCtPbgyNpf/c+7p9DLJ8AEDQ7luprw9sGA9/45zpnUY8GkMGPF74MP2i2tXjAr7XeI7QDO
v1Y3v6U8UaH1ZOJNstVg6Jbf3SLfWJiLKjIP9FgZlatU1tNtdcz3foxWhFSD1VSPCBR60vszg7T7
IILhOIZqHn8H+T3skRbK4BYiUP+MRYNvEsriY7w//uCyrZQafqQovPoYgVKM3NXj8TKHqtjH/L21
4nxIZ+6xdwERdMRz43JYOc9y9xLP8Oe018/WXhsvljf2EnTNVK8GCVn9tMTF1X/Wzk2YPppfIFgq
plvlH+/DWvRPq8FNcn5pyD5dymS23uplMOvREnZ2UeQngUeK8zWmtqoEqZX8LwFpXaT3+lT1W/+c
c700x4A1A+cbIGgWBTh+UQoSoL3MAswc0aexKwKBiw9+b03uQH4QDa2GqeF+zzAxh/O6XOdHn0YP
f4iQ4gQx4SrJ+XpjoPT+jkVRDBidVeT2LzKY8NShX2/C/YV5I+y9ksS+SQMbweA7LDyJQW+k2ePm
Nl2bzmW1DIjFnfKuukdXlp1bj9CDb3+1mpQE+VqStTX7rF/WxIlkN3BrYZp4YU2Cq4VlfNzrjTjq
OhJoB8QH+x90T6yByvDWOD7PFjf8sl9q0xto9118xiHiyvEzs6p5BWUyhxA7IUMe6nd2aVMVcgQg
/o61FFWKxLwq/2ueWPGTFQ56bh3m6wuMTpi/2dmxYik67tcBCFdWdO/ya0walOemVZeuLFaB+Ojw
txpK/zBELANq4w/5+zbOD/wW2TwilJNo4/wxR2xrOV94jyQa3zaU4BveoVGOPuFov/2xt0o2Y7jR
kqUsY8XhNvFkDrd1RXRhZEqyS2GuIKj9G/Jqan261w9ZhsJe6HQAu9EcoIBXLnLEeirfMl1UbhXK
SBA/l0I8unS3W0hUlSTOJM/EfN7dqU64LzekwcQSFYH//qPxERMuK5f/Xuhkdj/zLbRHUNioF7J2
0XWUJ/IITlK1ZHpt7ijd9Gfd3pVkckDgFske6KGOaLvZoi+WiN7gpso7rXI3TUNIQxirD/COCzIj
9e6aCh99Gq8Tzkzk1Ly0ePCb4G01CLixgZIw/sIxVCrugEhgIZtDDe/GqmNF1WCRZ7az7JErtSH8
r8JZELyYagC6jzB9a3WQz93AI4gEMZ/aHn3rKOPCXHXwx8ONBwhlWl94yng5p4NbKyhduJsZNQIk
HuJg6aGlqx6cCij+cVeoIWgWnQgj5/TTp/PtSpD5Q8ack8pfom2IJ5J0ltXLsjLjq5hr9pYLDNl6
3FpR40N75M8HruN66J+PfJljskjusNK4kzfHUHK1/j5M/+bXimYf4DJo0TA3H/Bix8zNuywxGUev
YIlYY3pcEmnJuEnz7hsspLP4bORLzyEKDpyjPSR9QeGndmLodLywltwaSE68BILjTjVZSqniR867
oZJ2XKWfIu8AZTJ9+sDxLFgl11T2qwyX1+IIVQRzKLHW40T9R0YrSFpjQieR/Rx0VazbdkS6eSKq
4W/n/ofE8X0JhYfg4dKJVxB3tXtxykA6Y9Fm0p8Q5v+AdEcB/9u/NdA3sSmDL1GZ/GCkm1qv6yER
ylEjhr/AGK4zXC//qF3qDX5ebzwWvS4SCWTNFZr/j9F1qi7PDXDCYl7bqcCPR649OEPp/87k+Bbm
lHRnAcSAQEYoJJpuLKVLO+RV7LAr0DsPnrR0ew4oKf7xAsd5p/tqTb5H2aiVW2BRDfhtD/zUFLBA
TrG+3vlcbNt+OdUlcbZd/TXeSQv8GLkrJ7+VznalSnKyUD14QPcRPACRemLkQvfvnhUG9D4DIVth
qTKgDYTjcfhR5AzzuZuq0t8Hx8w/Y8jNiVb2ZCMiglPSbxUmm+NB4VsX0aDWlAHCY4ncuGFHv3RU
vogaGr6mb0pvVGYlkIuAscVj7S/unUrItSr5I+6KqCXcw7KIY0vcynzemgYw8G+FMbzV75GI8jpB
j7ukuqv+m/5QkXgnSUuL04gqYf3cOkM1y5O8cT69GulFKETmmjZJ62F6Cprp3sazqNszdA1zjAUP
3gi5mtH/vEc/OEPzKotLQct+59ZSl+irr9gRV4DCGQ/LfCfYEhL89hZtAxFapOFLeusmMRZ4cEsy
ypi/UcIfvadglVB+uLFLTzqX/bfr9GwyY/qR0NLVzlO+ZeSoQZwMrc/LEtwH0c78Jdqh0ZVqZ4zI
Bl1TXuQFsiMizR2DjQlxtH/eZkgm1PJo087XI+mpx25QKtP3yt5s5f01bspD6CQiil1H9ANreDHy
VVzDqpUtZKZPYZZ1ZxQpHdiknortsGOh+ngoVp3jkHZdWLVVNOK3CQ4/W1WGyutc93uNviZ2A8tJ
ZkMKKnJKqDWV0xjE66UAxuD5jg2TuYMdU6iheMDN/zW/HLpizdvMORUgR6+AL0xRI+Z76+Ac+MFt
8K0OTyhIkjOMDnZlqvYsU/ii81bKqHWrX8w9C+PkNQmqcgIhiAQTOhoeEhuHjzemTrLmGP4UFD+D
7Isc8scSuC3Q8plNg4suxT1sWJog3PBlrWv+SSo3xbC9I6pi1RenXa8+a17Xmgcx2qv4fkJR/yvh
3dxEz4UOAEHEMNPReXrurfWUNyiCOax+wFL74LUhjA7++KY2KIv2QP/nGHNTxFGnLqOZX4TpHMNd
7XTnhE88prbAItfuni/aa7JxhEtG7Jxr9CDrBLpG2vXVTl6i7h9dA0Nch+SfxitRC8nDfz5tUvhB
TBYYOkM2YQa7YLFmnaDwB2kUjZqDwvlwwEtREbfFP6ygIpwyqMlt147TnDjWzJiOry+fEKZCEaLL
mNOsn5qbiMZw6Th57Zygc0xNVcV3x5XE0P9HN26ImiADV/8iGVAFaM7/NnM2fyk27l5sywPgIc5c
BEIwohJhDB2eqYTL3uhgBZLWeHThZDoNeWxDXcaWAUxxKDO80sZie9J8h+Vbv2OYtfjVghCkoSg0
kNxbVRZBa0FQa18j+bvcPqiv9cQRjvOhRUdSEE7bqP2Z/T0wlnjBKIzhYMl+MkQ/x+4mlFaDA6s/
Vu6QtQ2tOeBc4R3cSYt9OY95YyJL+XRWMETb+xSG6JkXFMfs/7PdF4JueC5dFCavxQA9jHfpe6RX
JgL9lMaR0h9b2IXUMqK42zh18fx66RA1GUCj8nWaH3GXobx7puz5Brm4xXVcEIE8fn0/aaU73kj3
I7bsrrP/bm0xF51OZhlHJmuvLtjdjijO5pFwNYByVWVU5LK1r8XTcLLuILx24TUh8QNjIciVREdl
9Mu1bb+W/HagfsQ2LKpMM4I6nse5Fmb7KeW/QbAtXX1FMsWeguHT9DKskXiVRx9fvGLHn0qcvjkW
b9F/pFy3Ok79VS62H2OCLdvyzTTCS0nvprG7EdiuRyRnwRBPg8DPUu4x1/l2KmspR9WoR/Iz/v54
f148n4FLLKVP/tlWqBtiCMZESeIzyM6s3GYuHUbp/c81a2myoyLIebH/SHU6xCBQd84Eau6ENItV
4CNwRx1/jqs3STg8uUciThddg2TZkqcA2OZkYvM9+lwdEGlKTuzuna6rKyU60OLwYgKYfdWq58sl
IFRCblyEDOJZIY24Ldh6rC6Z1Yo559d8YOev7dkNA7Zpz/CxmiUlf1h3BDF7LoN3iiA6ysTK897e
kUxXFFwBIVimbHsIs7l7OJq3xV4t/BsuQ/MTnlBdZ2h5Zv+KXUGMLm3HZmZ0HvcQkMUVn1Dv0xvs
K1RPke0Ymw9nfMs1lCq2jFrRZ5Fkdh8Ci257DXQfU7SJ/lUxZi8HEsuMn932OTK35hFYwppPZY5Z
f70BdKAFLfQs6SjU2ECafX7Bdyi6tKuJsZlMMKV35zYsxmVXFQMnQaupwcbEf+kwqDvi314wpKqp
gdZZYcEev8VyZWlDysdvC6J8iKwAcqygTVi1jauvnjXJSp/RxS7yDcoEAam8TwPamp1+FCMyRAzB
oOMXUZVgCgvVBAAwhmYOyKvw/SUrsQnZJUqrO6aVLesCnUXL6Df8Ag3Lz9vP+lTbIKCGoadARtp7
o5U3tMTYvHmcH9MuBgTTm6TvtyuzBbOUMZgQ0BWct44LaN94DO4KcxLwguRXZrMPA+dnjNXs1w71
S21/OFsSiVHD9qu82iCYaYoz4kX73xV2FNCJVi//Z72JrzndKCgV9OFYuCrtQFAR1SxwiFK8scu9
McLomzuYiSg5jXNB6p7plRYA5QdX1C67USZB6SUFJ1C0vBXwvdEQJKt40dtIvS87JMi9JNxxUS6r
tMguxPnR+4+m/ZyDSkFieikVvwqzzzy29pSEu7fbHhi5GxxBMP1d7vATgAGUab6Q8L3dPTSGjN3+
uvgLFU1Lf/qP6aPzVYdZHfRWvwlVlKy42kR40S2lwa3BlAuaP8m8DDN7DkGoeCKuRybQpJ1+84ou
0vyml5vEjqrJXc0BOTyuvGbL0Wfmcdg7CCXYqUcIQxCx6cPbEixW76NEA5cU5eQt8ACO+wDmTI+N
QbeOoJGsBFmK5An/hNf/7+lU7oV+iv0g5jfs/WqwA/FyKl5pIBPc+kPds6LoRzHEuTwVfc38ARuK
PY+lowy5QnkSGToCxd/j0m4pmpnGBJ8XAhVJuIVsYxhzCDrleS8x2Nxe96a5gLeS5waP4zWSPqLC
pDhN93LwGABK3DUeYYZ8gX6Inba6YtJWP6bK4tLHc/nB22JWsUph4xi9itmVnZvwYGZpabdF7qLn
DTqxAqWsceGjmKYtLOgZlBLogUKvxRjwVChdfJIxNyRHXdDgA0XC/04XkezqAZugxHXUl7qKhfEO
/7M/vI//k0VQOKEwSzlfRKALdc14gGqAg3UEcINw7Qjpj6NDgOxGRZmiQ8LKQ4hbi1dS5e9crcgT
4ZQXk1TgcFELZBvss0EM+qzpg0O8SeX/WC/rV9Sa6+LeW6HB/p4is0neJPW+QqLZu5HDtKK7tthw
+IKrq63/srg5JERT4NY4UpEjlmKayLswsL2WchTr14fPiDbEfNqdS1yi6YoKh/7CRK78QuWYInQt
j7wUcl7vzV+j802e9w5i4kbpCrlJ6Okl1slemC2zcBioPXGfvQofVC6XKR31mdcgfJrkmDOPMqzD
1zlwh/C7p4HVvrRmPjXOpwORsar6WQ9XVwtEXO6mHxO7e/+sY13j1rAhhmYyvDpyFHmrH/czaYdN
DSmNiY1dvLZ4+zaFuQBnVlOlIpF+OyLwU+vmmuXlUqdaKUOA1Ms9PjAK5KAtrstvV8pvvLAAEw9x
os4LtXX6qU+ev043PNv4faFibfGT/3PLMaAq8iCdizm/vmh+Axurqen8VPac9bvRPlhQoT1a/y+0
wTFmNMqcvGKL7GqmR41sCX1xfZWxmylipPbajhBmydDCIvNtq1yQrg9MGmNxBdCLQv+hZYXQnJO7
EyljpVscizqPex6K/9ineQizSVn5iNfW2u7ptd92TwTp4thS/nirPI4LYFDaRdGg96Ac7V5OoI+w
euEdGSxibAiJ4gi4rq3XPj4cQh09m2CdWov6IDzPfSIglPb29JatTGbBJ43zispCgkQmRli4vQ4k
x2dQMEiqvOKfKFOS1e+xuZ17Jrh1JR2Wmays6RfyZTfyFjSX/KlvnWJ2gri8q32rxYPoBZ4lIDD4
w0Yw6Jo2p4JinsZpLXHDrAlnRQDKkbxmfrW0xubRi+KVjJbhu+TuR65Ntzp6ypKE7nG78dw5QJlr
4+XK2FKcO5PKgv+DwSO7FwIdzxPvdw+zKRqmBQ+kppRsFVNQbjZqydg+SLc18hP+xaD+KWjzt9UK
XEDVc5BrgTbaNGUKZtJSuchG1SxJysrsS3h7f/uT4aIeKjZEehDpB5w3wUFOz9byOnY3IA54nfUc
llmenkvNr+GDk3ye5olJEDIekcsc3OnnP+WoHE23PFbca474oHyZT0l9Tm9BKFOoTULwVXNBQYi8
Id7qqda0pecIuD9v1ZSizZXgO6xqsEeb0h0qzzC8DPcyrcHUWep2eESndHNC6mLNQwEyg7Eu66UF
M8I28pb/axudlUovbnXXOG7DbpWwtVUtL+OXqVoLzH1bdyo3ATrGLvZOH3vSG0JOVYSHrQL1F9Nm
Sxz6yrhaRzEvsQQGCSXM9trQze3AFvpTa9/8R34eDwmCoeFmFRBnqMCzyq6uti9PrrF2lVnjXcU/
kjzqfVBltl7lmw2PAwZqF/5QIicrVYlq9iRTKgwtIFqG9C7ObLSdRlSJqconb4KRdRqkXJ/nLeQp
QJ0unoyVG40rhubicKjBS9/5Jk6mTwApNRmF4xwEMogJcqn5cu1SfpBV7v9bpzY4Qr1ROqPKdls9
odqQosSFaxEvOR+Ab5ckOt7iZOTxt24fEHgzueW+cO13HYFUH+ohZEytzlMk1ElwqVDCh+JDuo0e
l5YA1Nb00SxB4CUKQAvLuEusCTnpvyojoXx8BH9Wsw5Ct9s5H3Rsw9iUOlnq/yidPWbjr5N8xzVr
AnAgpWw9s9BzKQOPB3k01+vci1QKobybIYM2fJdooS8e6j8t1pnxSb6tCHrYCxtZ+9WQgpd2DPIe
GSVgEH+gkeO1cWY1+B+lbibQot6RLCgBTs2eJf9ZUwsxMj/9RTxvRVRsyxpI0r7t+EArbvdmMYrP
NtEWAY9jIxOj+7gku4oo696nkxilF8qRBrcihaSCArOPmeWuN1g49UAETiAzaWNi7fIOIAvhHpvi
H1nboBtWgOrF99hL02UnAXeYL3aM4DPxmOUMLcupuQF69NhttCAiRm+40KhUybiOZYUpnDONNazb
pXCIHjoIWvfdu6oZXgjpDIInf4Rc5Six1IY7GXWRgXOOfkvd3tddn9zq+AhskUKqh/Gfpim3VAzh
+Yr7kB6XMNwZsiplYYz6yb5k8e9RINeOtIeRHaDnODgtRzVdHLgMlRhvtk359dwKJ2XeoexRt/I1
Lgv/6JP5SIF+Lq1kWLipI/NodwXP5vlT+coL/GU1b23rCpdpasoy+p2Xv/3FL81AT2s4imbN+797
/uFX/3vE3Bkh6sUTIZsl++Jnsg80D32bS8ujHUGo4yb+2gz+wqgJMVTKl36CIC2MPK9ourDagu9H
Et4J5G/FNj6tcWPXgpc/ATKfGDl35tIv6o1wz2LcPUFsyZFTsGac5Pu8/BkXdWxe0sutYKhwUy8R
zv8cBThwi8cdWInI4SvnGh6xt+Iscenq085zb1mhcABA4JpWYmfJOoA8wm9/86Fd+8lvH5kwctrW
a0iolqGFJqeckVWpg3iRXkAg3o82JOUN54AxDoWao9UcbVAiE+IPnTiwnMf/SKpP0qlJy8TuwYYi
HFjCM4ivsCzkoqL42LWx5zxHHWirS/d3E3dwbZLFSBZuLdoVSoftxcsKXK/ftXRAYIOUsE3jrogs
O7Gq193yr003uof5CmoLFTziIiwvNjf+tiEmk6jEut7QRw16x8YsOybyq/cvCtlKpqSj3d7oPe2L
W+1ziVTltmpUcZOt1ivosAaGPdX8e7fmD7D8/Yu0w337Eeu/Uv9QyZuSfvFbOzjAj7jI8xbqMIf9
ZVFulEaiVgoIWJ51wb6qOguczqu4EpMiDrf+pGOZmZAos8TG3FIGLVdd4C3rqQ5lliTyhbW5OdIA
Sjl1yp1yYgZi2sYzWpEhmFHRUb5pv7OK/lrkPEPJx7rdTPLQwNmdGWWEeVDV0MGNcBg9sYphdzUu
8TVCwKsHj3n7fNI1LeMyj/kmNXf0gC5eSzwoFxpStiASYaTVERYQeDLS7V0E21amPMZOyRyGSiub
MMe8SaJyZjdnWOfLcMr7jMSZxO676vi/nQ2bAo/XdV2E8CUa+XN1NrU+rPcp96ojKgeIOgMBE+5+
sNrL/N8SMNbD/qeXnhbbDEEQLhW0UZ8PuDNNipHS9We+sYDYXSFPGXG5RUBs/SLLhAjj3eExbXGL
tVhE9YJFs3M7qN0cgr1p8pApnJSFy+puSLrwSHctu8ijxbMj5UBDDSN1+T3LcOgr76VXu2OMjUvV
LKBnvGit5rF4jA5wpsSRVZ94ucC3frIz99g2bqsD0+kA072SLDZdql1bzNyDGbmBQ7XNjVhZVcV5
cUBYpR9itTQqeCohu4X/P+9gheYeVLRqgl0EZ9x3UYGioosQzINkYNqqhVEb4a+++tVhUMV/3EYe
IgzHDyi0zGziFFaezzubMcJNKJCrvN9E5ggjKSzkhyB/pz+uyP6ce5CfadkvAME5u4AN2fx9jKPT
qCiBrTfJekNE6UraKhyoJzaF1gV+2Mt9gMSECdKc9kZMaD0ohGDU5zb2wKThL4dU6YEoJ9H1b6aC
8XJ5E9g1MhvBh5c6fncreXMf4u3O6RI4ZOrqN/kLWuCUdvZXGgYYzMatPGjj90oyOQy7ndfb2LPd
SLFc7PqHZbxiQRsnGNLxowstu6BJ9Laxxie+loCLnvcHiMW44DhEowzVHxDdwYCLi5Ac5/v5z/DR
AYc+qkd7Jr9sPnHzHG2Mhdms/c5tD6hLXWSpx6qxP1PPeHfBKpDEdOWn11Ho0Xirmzs0wOqe3dRz
+0OQdB+nynTuzhnyNJ0AYzNBVukP1f7pFdi/IOf4EHpBtg9nycGuM1jpPJytm8SncdaVQHIO/HiV
FyPXcuutp/qG8BQ4JyTWfRZdJyiAd8o/wQMzOsLmrV805nw89h/nMlBotlt8x1PrIt1acOCWNQlD
QwRB2p2X7GB2xxtdQ9e1nr+RcwylICkKrWMMWYAzXNWFyppl1a14b7pW10JRcFrtdTsEZz+3ne7Y
1gdHKajtvtnhlw+E68hvlcEQ6/jqLJJTUZhkscGAiuNUPrvCpXRLcjZIsCOfmkBVLt+/viSi+tuY
bGVLOkoa4g3nc1pSjmdR7InEngj8KxOv2aF2IlS8bqGJL27Z/2xVwCcypxqxksdnWcUGLsuK1Qu/
+/v+c9zAR3bjKjuGzZw4S6wiVhRHbr5OEuGRlfSA1DQ/VD/0kHxeNLUo4C2afBXQ4j8JnWQFv/ol
/Rsu9Cqhv8/f8E60XFhEW8+ZZTRuidIftQSd9EFY3M7gtGBV5b4BTT+5vr1XBV6X0w0At+GdmOZj
Wd9mB7A6k5r4zCNAIaIBR/Rg9KTEPWlnoXXhTvkIGqsHMT6dYHcCpYmkV6NwhOPnTbXyVOMk/JDv
fOr9XF1iTPFM7hkKA7W563IlARKq/g0db72iICsrlq2aVoKoG5KaLk8iZ/KtGYeqfCYaVBR+L5Vz
FgdfanwW5Iqy9f3A0Y71hq2QagfRDZnBn2HP+7sSszKK4RQYMrb0FQKn39JKksVn6mHKpg0Thsfc
qep69T283ix8pLDS/ktQDqg8L+Uotx4V+zx8bcyZfSUo9ZiH0Wy2En79vErj9+nCkaXCBxVxtsWy
33+FQSbiMjobLqeyKZHKSJXcjdILlGJQ2WHwOgPm52d4aWKxpr0mHGo5cR3OnZPZagdDsZ8kqct1
tA+OHpsBNhX0AZv2OkKhgk61jPvW38JSb5aavrn9uZmPSrRcVZUYL0Z/GXco6Tmcx4gqgr1neWi9
po9pAnexD8Dgon8FRRQzdP9SE+3i4FmBvkQLqYi0T1UgfzHwcL46b1yhafz40IvdxMCrZ5s9Zh2X
fyZe9lP11iftxaYqnyaF7AoaFd0yWpSkYIbgDAmx79KImlAZbq4rWQJrSaFx53xv+c1cA/w/9Bh0
6fCFEtiNbITOY46OnIlPC5PaSYRYt+GUo+yiODg0eYqVUWG88yHptnjFrnViJa1ceRfbYm26naTe
aY5UUEYdyAHRmKiEObHk2WEXOEf/RYbmVRnvWqSUuOavnInW5PvS685Zoc35AtzVrpYwH4FtxbfR
E8aT1oQtJ6w0IjXEuVpn9MN9bw+iHw1TnaILPJkyjWc6bCgJjAqr7aHl08sYPUUfqXC/HHo/4itT
o8z9Opj5YE3Z/4knjdMvyR9JJio/GOiFN3zok96JSCFTrs/Yob7C6ckxyjruwivLGVs/hippo38R
ZHE7owkBfMNNivtKpxPO2aLMIpsOF0OF/dII6BsUDZYdHz57Sgw1ITMklwI8SaP+544Pyq5W2Tdq
uUtstS6s10rXhhlgBdyDlaOUqhun7BkeIn7bxOvl8TDCcPZACYX1fkoMI+Zvk6rZNvHG5JXGQ0/m
mIfpRLZrNvUROU0z8oCA4jSj3FTMKFWI9oMiIATFkQlGFvPH7jo8t3O12g7GMIXKvbq5A6mm0Yas
SWlYhJc0XhJjQRKPG7ZrPs5Zc8wQPOAyLYLgNcs/UXyqPH2zxVtlMLccpPVgRhWzTzF08Q+bp2vh
wbc1JAPRf+HCYVCPtEA2RgTjKZk45UIXISEUaLVFQtEBypigh7jKkyeOQBCro5PD8t4HWiVmPErD
rivIOGwS+PaAyQIJNSnmhRDS1tuBfb7dAMIF3KbTsbQSqbr/mTr3VQWOIR9BFwDA0Cpt152hOQc5
n0qmyv3/kaIhWbNMnC/8eouNnCxPbP/gZKTVc6ZUha7t7tyGmK+j2B1q42MD0Ejcro2W4/KW7eud
giBTgGpj+R/cVsm4baixNjtItog9RVetz2XwuA/0FI0pNNyXQWm4GDVIJiy/42zUaDAoisrWQPs+
SrQzMf7WbLVowX2uE2WTgzy/BVnbc9XU+BIrJIseW+uBbnMH8saRrKlAAv8VM/OlsE3F/tdOjN5u
qOIlK8nis/5jidaJAoUhWSL+dQHsLDy4BzDJ+94s5+cw31we4IUVvNZpir45XERoJIrVEocQ9eq8
wxfNIPM4KqfqRhsL3gRnc4D1dZeLoy4WkOZJ1CoLHhA5XqETLUQHBbZqK3I7gKF4u0LE5YK5PJDw
hWEQE1slRriodhEN6ec0YvWC5IUQXtodMZVFDXQLvZS9fyJeVMVTNY3zvaF97fcduGnP/yE497JH
qJMHF5YpvZsLZytuiOzlgmzU2IkZ4g8QK8xLp6klNbsV6as1/jkkDEqGznilookXZ9b02hT/HLVf
uwcQGC+sIPdkU9Z7/ivTou53Qo8gF+gODDpqGsAc4nevOrchmvT3hj0SIkoIk5JRnlRm+tQvEiM+
t/pxd2mf+c9O4P/wAzG1E1EMwGDvwaIgeMJoIY+xmHNU+SoP3ktRVH02XoeX65naqoMKknFPa05D
7247EZm62i6UW5Gs/anMQyhMj0IbxL7lQgCqzjaGINtaq+2CkrAI0/uVXfIVkcH1zb/Mpmixe0nB
rWbaCOHCAPeS3TZw8fv2ak97aQOlcF5CA1cfIqtWL9+H31Y54/bxIaHHxKvXBOiLMueRFExHjvSj
WFMS4wIm0bEwmjWGSPgEFWisYG2v297/LJFraxLHji5SbJ9oDiksmGCKEtqsn2qGD7MlKMOa5Qpo
Zc+JvfUeQHhmiYfE7F8/q7rf0FEj3cnhHgN86/zPvh0zCjxTr54G1egGi3JouOKoPXYsri28iDfn
eB+Z/eTgl4TEABmWJiHfj23x20oNVPOMUhCNI+D92zdkWfHYQZjuFzPBLbfjUYQjACEVGo6EmYJ9
qh8KsOmifQgYJJQiboUb+GsByIp3sack/Sk/MOetiHnvLxQLVAxtjIl3Q2RDd2/2017Patw0zr3F
QJSdUy5rMQoPfc1vBzyHVQrIL3SSNo65hFBbYeHLu1q0T5WLNRzq1IHlFnQmCvf5etEkeG4AWTcw
TBYf9lLJWU3O2Jw0jnXIHf7OFzlY9rnJ845VFVJIjifRD7pvwNuyIvIz1Z5FfOL1xI/k4p+SPRRX
KvVr1pZrmlUn0y1JwkTEEVEVtV5KIcYm6Htl1PoTw85+GfX7SHbFluTTdPRG/8YVKdb6g+A470Rz
f9jXdNicq34w2PzZBu7l9Ti3Bb+4bOR6u8rCY4wGRecQTxKbhbr0ckVpzQdaxmPTC4CGNPWQUYVg
a5X475CmnqCHELlDphy/B/JQkU0HYwM/NvJyqhpwzOoyzghnmxc/m0TxylIBWUmGmUqthnV//cdJ
EkR6Ob30XBDnXxpFqznYE57zFB2i2JELT2RS1El/XGLBsoxFp4QYrL7c9QiYc9t2HaJgb4vGLuXh
T+t3PrNZ6SaonMXlzqjiY/9szrA8Tg7D1M5crnJsn7MhLkHLCfz7bdYKfzPjqX/E/+eVh6CO+ma5
2iwXdm4AHyyA8vf4zbM/7Tq3JUBcynaJA71RSfgYsZfsSwaTxPTmjMxejKlsg4+lkHEwjmxrtZEy
JNONKi7wdpp4Fkcliv74h6d2MtX94hpYcm+pChuRGlvaajILdL4HiSLGw3Ixd43pTJC7C8GN0Q1q
zUJfKiOGr7qreS0xX5OBBnCcVDvpGxwy00wv0DaBQ7Bw+dVsuEAKfIEJr6wWekSpOh5O9tTxkjKo
UWXuDYha6fz032exmkXcksohgKTCGltdwFJTZl/qXyHn57ysbm78HzHOH2qLWsZVjhjRJuN5gm4j
R5gAQP9Ee8bV+h3Xg9ul3ePb9R/c6sxUwTbbuKEy97M2th1+vAH0CZKRlf+zIDG+b25EZscOmbUV
i1Efi6naQ0ypvJ4X8BsgcmYtUhx4Z3qrwpvbvEF3aQlmR3vJXp1PSi5yUtcnBmPiiP+fv3ceLZCR
XBfh6dvfC15MZyqtwkNSiwocIPC3voKpl5IwYcXwNYHvSN48fYzUrR9RZXwdYkIrWl06DcRYWhgI
iLNhyWmWH6uGcCbjAwxuQUMTXRClJC/hVs+o/Al+v4oe2oH/q4wiNKNzjRFsE3bXwhr5sAB2dO3m
QwD6u0Rd4vpUyVzESO47lQlDoNQ9l6EAcur89L1bO9eIMhEZy096dCp9Mwv8hge3tkFryBbKmbeI
m65LJ8TYXJFky5hyfOrDd5KHAbK0Dup49iScR3Z4p3dbXIZgZ2m/DxxVxaHnYBlowLXz/Izbo4yd
MlJdVanjU1VLtlWCjH90JeLFMBOu/ckS/MqTaPnBVCSRPtAYfFow3H9Fd0LBv3mn17OG5FbvKReZ
QtXwoKWtjexidVKfMWrLNfqnQbSQUr5o6tupQo6dTtK+/xy4Fy+u0pxZ/nTjKNUPIPR1Chw31Nk0
7qIcyN4coQsj+5y7dGGngTrdHA+nkIzXcRY1VI7Lpoe7N+PxCZ9DeFQDjzMmR9PBFE0VvQPRq7PQ
ebEf6+gtkO1Xu89bhlqexqILqhiIWr+AQcUO0duN3WG/d+TCviRqAOGUryWN5J8N3cFzx/OaunmJ
fE6KGXc1/w4TymVjrPdlguGGWcMylOgl2Q9XZgOO7ye5dhwsFQB1/XvSTXme+NcIVC1YJkQqjlhS
1YamIvglVqmnxX4khiF0suCIWhByY+mRWtqz0IJBa9HbONTyNWmQasG5rfsajgKaQApJvRSYWL+2
BQKceYn5PTeLxbRc7vhawWggw+cKBprLzxGrNYKUsbp51Q8poQY7bazo30nvXzm2zgFLq+RHN1wG
dyPts4B9FCnEUhpf0M0OiIbw5Y8EkHu7B8CnlBlndm4dVdqHcosOVespHFobs/6MZScq/FRD/31v
EThi+46hR2gYdzb62zw+aWPNXazuAUiAEdM6yL0/Q62Pv4PMiVv7DvvDP7iZvtamCU4xJjARp/2T
kxkvggKHpHY4v30x9D2x/SK91bhTbjqRit8CYaeofkOwsaFhxjqyNovPuiKqqTS+AZsmHmXF5gmh
MJ5bbohxlWgcgpY6FkPwL0E8+N1fApdlsLgOJJ4uPYqpk1PbNOJA19cUxhpftUJ85Qd1FuX0uYAu
mEonQnNYqCO9Bmd3EDrs3kzKe7W12ZExJUSGvRKNFcvmLoMKsVlm1V3n2P3uND38OIxiLfOCg+5E
gvzjtLeOr+3l1swLNENwbCmUI4GNiOoqOZzFznxlgfdTtYWrFY8k2wBrU1knAZiudprIkDf5NHTv
qHWE/A6WGDuT+4i5T9LtPz3d+hlsN9FTAnyBxYBZ2yr71NywwaQHCF5AK1H4Dk3suVcTnBZK5Mmx
lem3Z82g04qhRDmwNB2lvGO0Mm6ZktP4RohOJ/TwoHeIEjk5uB3Nv0DqYbyuNxDwKNIplYa2f1MJ
P9wdi2PRf79gOePMM6wLTYfOQ678LN+p2PP2kvra2/OiOkFuK7FisiHejSq7nOj7F395Rlzn4HgQ
Huja3Enlbtpfxri9szx9VDw9urYisslq/ov/avf/VQj4On3rNtUKi3IeJz7Ht8r/bHsSQ73t79Zq
qSfZEiv+olL9OTqpMlAeU914Ckl8424ClQsTtVn3eJ8OWjYVqJH75YUwLao/+KP0XipNXXBppbM6
QoJKaXuderBgA4xVixP8dBn9xAaSvov2aUF4PKNy1XKnGFI8JJgOhkP78MLGC/fSgjA+atodzswf
55lcfwVV/R2SU6yMYHW/vmxjEhHZlToEu9dCtlVUBIQgQy8f5T2pveiN0OHLSd+vynx4KOaQHx0Y
gl5KLtMD4JJQ24EImG+e1SLdHeknj4nxM1WzGfKAfGnzTSz811OK0SOrmRsWnsIhqjc/vGaSPuuu
vaGFeekVPB8ix1gkz5FVRMDbrRXVlm17tx4Lz5gkyvY46d/I4LNWph92cCONQv/AkaA/bMAnUloT
X1wLknL8fDcVk7tn7E2T0CncI5p7mOFeH11cyDzEwocybXryNVZj5NKFlss7V3ScjFcMc7XetcCV
5i1vITM4X5oFQK0t2R/eEtK2NatZCAiLCGxVQ1Ish57bcilXwWwmXzi27KYtm4r+BlgrHLfMNa3K
/N3RE4zQxUKDSs8HKEH5AATgAw7bwNgJlCmIcccuAZrEsENabxxGS23TjmEJopASqf4+EhnFRd1E
PR1zSecIq3UwxYp+mu21epX8Qc9Q+0RYi2RfWqNuKQQ5nQ0Pe+fCBkrUYjrgLfq1oRF2ENOaO9VT
UkBZu5qwaU6eZBgA+RKmYYw4aYDfYKXQM0SURSAzSORoHjg5W5q1NDHL8lg90cBxr+Kaxo1+FM1T
OkhPy1pv0CiN3/CYtuXFiOhosBZnL3WR/d7BPPLa8v47XberxGI3oYDmQboad55KSDEXBAXZsAyG
gJirJF+QHstCMI7A+m5HJGICg6D12RMse2bsxt1XMXZwjvMOLnxgvzAFKtw9VLYW8juQ0b8RsNAN
RIykEM2uCqqJ2szSGkfI2zzRsljI13AZcE0yJQwYdpJbKgPnZLxqRdoe2zhIbbishirYwYABCmoO
4u659+SWhDGy5yjsvLEpfnZ8lnXrY1m0Sz453Au+WJWoQU2qh/kMHXcN6ZPqkwh96dOwGj2q7Zy6
O0ZjdRX/AkgDOlxRoY/58unC8RiksZ1+w4Kt+7L6HTykE6++Yowg/uBbddJu0inGefZA44+Q0WR5
cNAUHTsPlOh0Hs9jhqF5aHkYBIFFWuMClatzpZL8vEyzDFJf1zi4JsPlqyd0BeiMKOHTmr9CeCyt
vvGvdEuUhl6kDt8eq/8qRW/Xe6nJKvT6r3FyRgeQZmJUaI3ud5EVnSFeMVyQS5wfNg4ZtqbSQL66
DpX1fYaOCVAElM1UGputCV5H4Gp53UQoqHks5lbYB2gkm6eDoQyaE9MuJB7dNhtBqL3SM9liVDS2
ZQCQ3KvThQSC66701xuGDXNj/A5EeFhQLmYiomj/uejXsKeD7GTmCPatj1i7UTt+r0Y+mHKzlPtg
YBS43+l2goEzZA5dkmdoETtA17/GTVm0vAJZk7sXfMu2RAKQXdgSqw+onG2xl9iEPi6NAEuH+rHQ
oamd/Ne2h1J5AVIlR8OCyZ4RI1OecIExq3L9lXwzwhkwYzBh2SfqZVvXFuKKdDBiUXriK+8k8MSV
CISNAouYtGdbDUQDb/qdwV4GrqpBL4REcpD8DxV7gMciKWE5/n6lHb60wlNvG7Inp87xDZmt00ON
lx4tY7gqLiYK/3QT6FLsa1Uj2VV9L66PCQQogipERQW8lMTUi+jmOO/JPpPavTkwcbXj/dJFHH9G
Lx2stSdzcMHFCgzCP2kkHe73t/oAc+Oq2aPu0uuLnEWQJnkCi7KQKEdfNEgKynt5jhFRUiRT3tFm
DlIspzQFu8qVJfcN5vRJ0P1m+xBIT9LrLQ8su53U5o1rVDG5Q4FJz8M4J4c6gTYsFi2boXIDfxjt
WUVtK4k7vD+E/VOTTCSLcQJscyO5bXic4iCvYiYc1YFpZUgZjuR+rgs5UJO5Ev7HnBNyZCsZlYKy
You5nMZ4FOtzhewXrspxe2gQAbEcfquZiB8BYgBav7aXLzLm6oLMdYjiO5b8Rw6BWtFbpcu76TdQ
XQf7DgOhyEASfW/IWC43u2vq2U0nW8mPXRK6LJhIB63Y29E0y0BBrE/PEH4VahovLckv4ggOKYlO
PXWeGxreTERDdOQoaI+6fK5dqKd5TgqyyVpG+rvIInRyk0g0Wttw02orYZvT1pU2H5uhtjUjzIZz
2xASifklekGaVb1WCY60TMtHeD8w0vwH8YvHjVC2J+cF7HRYEmmblzTa98MOFO4iH1vI7wBVVN+I
TMrInVl4UX7anfR9I0oS5oUrAAIUrNhBTji+ARoKt5KvU9WBY4fQJjHbQpBrmxUoUdhEtdVzLX/b
avAqGQOLJ9TwpHnumQ0gamOM237+2impuPFB8jw24rPBYqWLvV3D4XTqZ7aG8NLyYHn23244zIKo
T839rrlDD/Vh49ShqJfnUTBvPFPEDtvkA+nRZfbEZawRBeJlvrqyIUr5uD7bEKy0tF8vv3xcdwN4
tB//Nmw2noAg61Iud0cfgY8UOs3dBs8puBmu/gAARNDgfpxaQ3AC4MqvdJEbFb9V1C2z54hok8H2
z+Rb6dBffKly46f0Uwrw1lWDDPXo/oLWl0sivW89LRzDtqb/5KjO/WIDGOSgGMA2TCLrnNQNIzgY
sZTWWrXjcN+WbV1NdBDCnQgqXS85L6okswm+Ac+P1bKiSZbvIgv5w//8GmmAjM+XaTEtmHortPTW
yr0PeoRhs12dctlBWfrhrFpI5H4nJwe7kcXECpiqPtDAGzXYer91B8XRB/qG5tnDZuPWRK/A0b7W
hbj/BjIRH/+zLW1oI6Oo3qY985zEaILJjsjLgJ9n+babKoFJod1k+AWQXs86N2txABuoZ1LxihXl
VCFn0kiBlEnVAbGLWK8I9ebDS48wybGDP1pBYSW8ZXBNVie92duv+4Zc0g6bUE+ueuvUz2RgtCfI
4HqvJ07ANm1SRUEq/AZU5fxpsN1c9Y6HuCYJ1HSNl7b7YfrCDViAnhdxM1UkBGOepmn7Rtc6lo1M
73i0Ci/nESWef3KiDGYxsw7CbJBtQ75SUXjiVE7VrwZpv6bG1KcdkOlG8MM20pz69Rs1NNP7Yd73
aLiTgPF1742/G34vXCqGwWsvD4RDgz27s80BG+qLUpW4Le8EPeuIDGONesDRkA4mdIlCWd22ntUB
G2bm51rjMXKPqfLjoZoX8acH9/qRscvL/amihD5P/bGq2eBsmEix1mc2RfybfkLwfmNl82V8VuSc
0n21DyUBqSmpP9nHk7CWmCYbNgqWj2KB+6MlGogpSPXai5x6IP5SSlJo4Uk2iWEfzpbPmR3N6jL3
0qokdVpLBgcqvF51N1mrjwRxxN39TxYLhLAIOjEW9+uiezv4/HHk2BQUxhGrRhWOGyWNT3FBNp/f
KGH46bD1RkPFQtf11eff97nPDVnkpAvumD9iZIqixXlUsIQGRpfLntjkI97QPo8949Gt4wbGNuJO
/wTkSFO6/QZXCptvt0IQGgtJkMUGBmYv9LsO7Cl5vlnUMJSr0J2U0XWHs0p+cR+IEh9gkcZvokD8
//0ZfgJTFeAS2MQyHKHShd+75x3qcm9TajrgLGcUkWoptbJG5lCFp/e09doK8Oi06bVEiH2t8Mhl
LSGLJaO1NybJ9OhCHb/Dz466IRWLu4dPgone3izJ6mkPQoUHlqxnKsmyTto2ltP1CD62YkbiepyI
Z3JszIfS+q/XJtRa6pO/ZEPNxR3sU0vlv1dvP/NhXAJ5m0qL0BIUcayji9KR6z8P+bM6yuVLs/AB
EzjVqNOI0fMkCEU9dpvbfhUiA8ZyVlJiHWfgN/CO88hbDamL/gwO+sU3hwP+7bSaI4nZo3Ex2bEj
C1zXHh6a2ERVA30cZ04WauSTexEdBOI4tArpQJ29Uk93z7FZeNJMemBKes/BmKj3+TgnzHC2Tdi1
pMr6AmW/MF7V2dnnn19gHxAcDwF36crX0m+hDAEJu2tqqz5ysXJU3YMpK0GQLNkoG6Q6hG7WizqF
d258D5411+QnY9mdS+BxPLfTkJkwNK6TDI0kFMYOkKGRWrz6Ymv3SLRfvtFf8726wJpHzGwNL742
Yq1KJawk1B84JOwAcH8hAcXJn0ixHZQjsjRGWS8+CsB/qvbfjqlts2pP6i43iv5J8APIwe6UyuxW
njSN6lJSuRVH+AZGQOU1hRO4nvsWbWh6Omd4az85Ww3Hdtp0M2uquZCxt9gR+eqrO3B/SMhB27hM
qrtSyP11UCN5D8xbWuvZNoZBLWokgRUjWdZ258d4x/xpr/2Cj+JBIiVWg1so+y/z7Vs2c2DYMPEc
CRTIqd7m32uaPG8CTfVvyRP2KBjoQB/6LoJNevNQIQOXWNu70pm3OrBPyqS/XuZWJ/KIuUl24VdQ
AbAUWUuudkIy7iQV6rKK2OP6wGzo6fsv4tieMZY7T0E1J11hL8nyA4TzXrq6lv4iU+IZ2y7I1xKM
qcjf+Bn0Q3Si9LTbvsr21SE/QrT8rCjYKnEQ2xpd4ycRqjgZxbrbPM4d3G6XIbtkTRuS7zzUql8F
xrB8V/Fcum6GM4ZqnvfyYtMk2b33KKc3+9e4ACTtXtdvp0PosYvNYT+CPgcRSsIbxvXqg0jwzmol
Ne3ztk16/FUoApnTjH7+/3p/Ux1ve8IEROi8yE+IsccDxnQP9YibTvuMU4YnXIp72v25G2m51AQD
Uw32/0+2qF93K2hlJK2cmI59mW9B4vi0Zm2f/Rdt2WGIiRGNmbbx1OnNBbO+zT9Bi9jrZMFW1gQ6
RNNgnLrWWrwsQ7mxzClAp8QXjXcSex8ZVq2V3SECw1Vx6WCG1HAWjpMZ7isDXxtHPQZBNwhTtd2s
gC2+IUj18yi+2puExOa9ZzheowWARS/xka3P+dwBNktSJ51/E8K0b4DiOsXYvJrcMJCw8Btn8SYk
qacV8JT8xb6pT3FNVAA9D3DQUs1YPqShf4he9FBinjsAS1LCfkYQWiy7JuLj2RI6KlnjTiMbd7AF
Q/99tf/UbWRyJFT6niah/Mwg7/yy6DzWwyVuF9BM1lwGAk0xgr3fU9N2AvPsn1ukr4Ul+nF+1mix
8eWHuwPsuwsZJiFhhUP1/BKYEkAAEiB+rRWvC5fXvPjemx0E0XHexzeoxpaQwTlY81tx24FqLxon
xHExNWdgN7F6aLDw1hV9C4ytaWkNU4AwxHj2FnxvRogSiqNSdmS181JeIJoo1GTRphzDmaHgMbnO
bPovwVG585mfOKELjbiC+WOgzFuilEOjWtVlqz5xVTSqWISrrWy9P+xD6N5f0gmZwnTwqqukBdRa
XY/I9JYCH8kbbamehJyTbLkVRXOya08m4pK95j2ypzvimECfgw/wkA6Kksax4Munf7/57vkkHykk
pNrrVcX5WlBwKXL4pqkM1FSy7sZiB+lrl0UZGoIL+P5k1fIcYWMJFOvbXOlQkUShmMLspH6OARSt
OthqMFSlDfsFNvPPdgJ7GgUEcLXLHL4X5JaTGsa96MBRdF35wOV5gPP1VVvTDpfWp4dYGfp1ZgLG
Amj4MoLi/kFqHvBohA/7nKtK8PgCwyoN2H6agjYhCT8lnbG9s0epUGP6qW19EmDy7TCEZU8DIDMs
9ITzAWzP/uDOq/taF2srXXaYramVfN7Jmd17x+vlErz8DjrQ8GjH5dAqM0fiVV+yRwzKa/3oAjcm
m0H4jVMdseiphwFgGvkRcUA+6IS3/oGbZtHR5P2JQib+ZxlpuaNVXgwgpXC8BpblTrj8mbgqHQWa
5xfxzvSBuRdm1QPLOpe7SGoS/8hm6jH8SIMGChwJ7uyJNXyCAyjw07tBaArJbq18VDGMSD0Z7sFG
/klJMNJcojCU7OAPImP+Bz6vhAbLcfBk47a8y878MR7StVBw4//DhpaFWSGSKjtImD62TNA3bjmc
XjeikH9j3Uo3vNQU/1/C2MVvQ8KIe7B16qzIWqZt8urDmzVeT1oryAAQ+7MAE+zWXAkxvuJFJiUk
hEE5wGf0ZPg6vyJ80J88RscJGiP1FFRhfZMpvRhnCZ35Ymybt0pKAPhjRllSvLm3YrTTk8QSfa5b
IPdV2KiUtoio68VZZ/Up+0i4LumosjRMtY3HEzekieQ8VpWz6qiU0Tgy7RSk2aHH+ydCRJCCE/P9
aBMgNGL1lr9kQH0qANXsKb3Q4sgfEuLgy9n0XkbdM9WOM23CYsebHB7BHoz9cE39t/tjOoAplyAg
G4TAmRNu6YAA8jVn4EQJl+3XAU9up+7nHsu6u9xaTWsUoCqRO3dH0cCokk5RBgdMINFInN4j3hLo
1/DgXJ9o5oCPIzLYClBR35xfPFLeGiaQlkSL6FOSoiJR/BUpA/vwFrrpGr2ZG4mjBrEul8jtgt9j
CoxPf++ux2u33kh7lUkS5vmc7s0xc6pyQdovph7MGpf+ZvEW4EbHN0sK/om0JKDo/INy3qcbKx8h
fFj9gU5kfIKwehcGY0prEYPdYbJkVW6SOHvxKYe0o299f2p0wZE/LgM1uco67ksU8e8dEsle9oBN
7DCQ3+FHwXW83bb2TYI1snZ2vwnD3Qz7ERUIAnIvQcpp8Qt4n3v1p8da44r3GApM/GQc8IonFNyS
yfGG74qCqaqntX+X57aXE457vAdbfDm5y8T1cGZTUEkbcAVJFaTuY5C0THR5k94VvWRSUL3Yw6Ua
5sq6ttViOL9Lkkq6BqoE3pXpjWlZHWYa7e1AVJdZIWlz7KOw2516xkIr3QXQpAzJy3Rn2qOWOMm5
mJGOt0iX4tlf+A3ogH+jQOsQk+TpNTaxfzawX/QOL4d4FSRiXkRq/hYzxz9kr+B8h8NnwjEaLLxG
ZcvVQpR+7BIwx69WMpoJSrRPc9YJWcF/NpalLBVQUCOcjw4vMUy/mAyfzgjMzKUe0/UpyFOYFHZE
HHmR5UgsJoe3fYy1+6ex6dxYhXJNheR1dMCa/OUs7CV3+oTIlvp20tvxysj6efdfVl317ZXLJVqG
GzNM2GQDIxVj5fJov1xprI8VwQFneFmn/quS77pv+HIHBXsQQwAqAagoJgAaBTnnPj7J7dSLt+w5
RPX8F2KZXPOG6L49NaUMHv5Ut09g/jYReWN9R9ayXyDhsrTgOLQzBYiCMQmt6e+XVm1XKlTxMLac
KlqLGhY2ktwb4eNbYb8sudYmuLqlo4RwuSQed2K56acx7SvtTUlhEJVZvpGPUxpCpknQY13yQhhB
x/FR5uKq7Yt0clt1vNmW4m40HJpzsMJthF0Ohk9H6KjUu15NNWuY2E++KXY2XyB3MQA5fAv7lfNV
eyYkPvEOHVkIEcTlB/Z4hhfjJKxWa0S9Uj1a5kRC3X0xklsBiWC2/7kUmHYcP7pkgXMMDycUVQvB
AP+YeI/TX2vo2Ay3SiJYueUoWPOf5Nl8zKQ2XaxTEsYexIyvidrWBSx6rx5Sn7A9YErm0hdgjCRV
L5LT5w/l2V4jm2cxJZhyXsc1zrXvF9RrOHuUgPkAiD/KtCK19IQVcKP+4XOce9tfYE4kynjVjjSl
gotodOKc+yAZY2RL2cdQhTKGw9r+N2Fuq7Szb670qbelPufCkzwFrvepoPypErSqWvL8LRVrZvh1
op8wXzXBCLeOskXVha3ZqaZmMt4poRZ1a04w6lbH653pF6P7ZOErkPKXSWGs/PhSMY7vV4gTG0Rv
o9BdahZPyr7VJA1GFu2V2mpFmRUUHMS9JNaH1t9X5kTCb9fAcU1IiQgyGUOoGWNdkcs11xfc9aek
Et3neG72LHneeVtGVxq7Mh+IDobI2/gC4LmSYQJ94lTwHtlgCi2oGLBCIQo+ApHUqpfCkq39ntZc
sphP5cuHxCaz/ffVGsMUqvN9UVWMFMmGGhb5jS3mg2mtpoxjjQw09JV6wPCPPSL/ROkvD7VhJdCx
P7f+JjLnGCA7APJLU5JgE0xITvjC3Rj+rsUDCOH/dmUpTsSIbxr/F/t9G0nnRMtP9JU2+57NWcr3
GIjpRDJnn1r8PuC9iIALF1tySzbkulknNOkq0WFK5cjzu0xhhzFcb+KcVXJT3BSaMlEO3D3/pZAA
A07aJMAbQ5imAX8jHcAWSxDj+AG7jizhBCj7qUnKj4Yb2L9TjrEIuclBOjhmTAKNVJyBpsHJUTRc
mrEaFKHzilgLOTYpB5T4PFQ6/JFdrB/j2LyZhRo4UI7VarzyU1WY/4nS8+RNvG4NiP/oD2nYBEfe
Nhfwyyfoc8vd0cpt4DquECOUuVSRz1GCa/d56sL6/0UkXN9JnJZW6j6sEYzDIOFnBhq0Ls8oOmSH
IGCOzQNm73ogIWC2sfp6y16761gL+/nZTitG1D5Kywax1dbxbShtTaFVTLDnxbG/BOi/BEsd6tBY
ZxiFpWZRRIdtqFFiBlMIt2YL/0skGLnlGyusSkNNEs8niUW1ohQq+ZUilnAOn04xnR5v82de4UMM
nnphEdxr47BC4Z9lmTpgLEgUkD+d4hgJ5NOoz0CwOccY8va7HOfn592zRKXqBFgUW1OuBQtIuMMv
SZoTPeQGIf0PW9k+1K8csGkLST+wrUb4DPCl0SdL251PbmKW0p8lnQ+vq8BafsD2IjDO/MJwaXeL
KgPHZ8IWoOUvALgD0yxqkWFQyosp99K50wtZHcwwe77FWAhj1krwjDdlZOGfEzOMaEarD8M5zfYv
wQKjVF0s+zwn0CKDPP3pLuqaZbYiAsPw2hT/qCSWi0juKYkdTsxrHo2Z31qmmKk7sH6E7VJ8r9Uk
l6AwbAOMB9Ua+MSjCF98t0EnXBNB7egy++cOkhYZVEjuyaM/ayGIxfXne++sSVD+vlkIW6AeE+zA
ByCciMLqNKjOCzZ4jRp6DxYR9Ky0OoxJhBVgDuptw1KbkecFgT1DNoWZD0Zu/JIkaga+JqFTF/fS
aVR5R2RsoPPHRHWZMwy2neE8FR/j9ffOEzXU7yTbPBVhFxqgdXkmznJEG2IG8QMTn/evEttTIamZ
9XpnGmo14mr3vacAyb/+EDYvKNAUbQXer2TNXyo/B3HvPTbuDwxd4jHINihkkQMq1NiQCYb5RYEZ
gI81Y31pECXUtXJ2eOHBuPfns+G2RDGCNHVlfijGzMtUr8TFjkaSyFBlrgbt15WPu9avs6wv/951
ooehflJwM3WS6hjX312TRrRZ6p5g7SVTSpvYlWwnJi/xdQoVbCTCMrv1FHPWrRxlYk3G4MznEPxT
UwPhPh0qyu502TUaBuZ05mN8tJzdGjMAo5O+vusSHBtyxXYPMhm8y3PrVfmC7lvo/89Jo5yy/2bs
gcKIOamjb20pRGq4q/qDbPizCfYxJi7X5DevGFqWIdjXlKURtkLxnUgLzuEgOD+I6DLRs/D1h9iU
JG3uBTyBIpB7DiZ2TqJUzzVfK9vJP9N672ZkiHuhUgjUQONFlHSB/fpdwoFbyn/dDdcKqpf3RzYR
9qrzDGTRH0uCEOK3pPl+DNDucmZEhq/PvoAYlneCcMp/dbXbs8ouqjulgi9aCtMA0RvRC4rj7emT
VBW8ohT/haCEo0k50wpQVTFM+W0vC5MgGKtdzSO3nn7ptSK0+He9/6Uejq+QgkJmvIso+pvehOIA
LX0dFqlRzUY0u+XVBZ41e7+X5gV7cmP6IZzp941kdNed8VhJeybReoPJDYqLTMDda4copJ8I4omK
bYoroIzN1+5kCJ63CyDmKHwc2nnwKMpFg2pzXSbFjg0C51I9hcMx03+0HFuThQ/Hh/D76Mj0QUQN
TpeSluh9jzq2526NHdf2PcFEjTjNuY3iPhaNM9E10zoYIbj5QcWkIoIOORXz7mCA11fCSgjriuOx
z4F0CF1ls6kf3YZ3m8EwwbbUHfDW9QJpIgG3zX957AYAqgLK6CvGQfjz1Ldv0CkMw3tZFO2QKDxN
nh5GNb11ORM1hRpquu1EhdtntoF3hMyCgOJls8I332j2Ev5E8fpKKxlU1JsrsR7z/qlYXEHId5ck
WthTRmLun8kQqk3ypP7sNrWS1rtH/hqiPf+PG8qhcAgHjbEhivAHhasoA5MHf2s55kA2RAYXGTO3
ZmPV09tgwaxCbQlruStk7a5mUucCgitHsViuKRcTztJ1B8MyoSTsOVgruXfIOIHNl3aRvpMVw/R+
hOdkGOdxeYqi9jgHbl/2d3liXNkePi0CIekpjO49O3jLw8uA69IuDZGM3INfpNdKktw0gI4rjaaN
YYUCalrb6qgF0SdfWVJQZfhvPW+nBHOlw0X1TpyrI2QtEngblSxizksTKlGpo0JjAeuk3Dqn+EDQ
DAp2Xf21gOBoe3kSw4AC7yiREmvCOEXYUUMK8RWew+VQ2dREjGcMPLRf15Ihl+xw0uV5oj3lOJvx
ja8ZG2fC2nwix15xUl1Tq1gc3xIVIJ7UQFRmUJ59B4pslnRSiIOoM0ay3eHcO8oCTrRe+YttwSbq
Ndac734SDNNo61kCDvlPpB1AlIGlOay2Ffy2G6VUkHXPy6rzgMGmz7mgq37hIGEKasPbhl1Gwr6+
fjItJ0QxKBG/6PIP6tSSkdzA+33pg4rOtQ0wVK8qx6BxpAzpjmynOdzwS/WBLQSZy4cHh7qVGpO9
RjZHbhD753zA/Kmud4I1h80Wncj7LeZCq5g0GCuWL9ZyCimSdWeprCNNuZUYDXz1JUIRYuetf68n
q6fZK1HWaK7nSk2iEYYbhPQjQmUS2ARh0zu+EYutH2BSl58mF/paGWc/WulgnDx03i5b3bKdMarh
A+DkyTbL0uiHrmFbYdXsMUtMlgzndY4EmxkoJi92sJuYKD4IB9sEUABNIiFFBRE1/j8/rdj1scnH
USmg0T0Ac5ge06iVe+KUegyk+6B7XX3IgQA32b8x2fq06EfaJ5GnlAyA5UsB3bLpcGhW64PV/dVN
33K6YChgiC4n18mZ3gCB1RPnXFtOL+jbcjV/x7BykgiBT7rC+SNJfd/u+sWwmtNNbYQlQyEHtUXl
f+BG4xdczFS7wUSSq31a7CGj9iQQjSRPyjz7beEUy9p2O0ZJxiL//o4dEXVG6PNWgKKa3BGNFRUq
Xc59WimMdJ9VjAO27PalEseKkmo0l5gEyFqUXRXOyIJffJJkLDyXlFXiENQxDjp4oj/1qy75/1Bw
jr/1PqvcjC8+cHEudmz+LXk/s9j4keh/5qQLy07RaI0IQwGrDw7RczndE7vbQ2PRvWY8VNxi6aas
IaPU2xrdPuSaJt8BFEa3Higkn9HJm7asqMcBCpziBcFwADRIf7ZzuuAoG79+k8SAIWjAGfDJ99MH
s3ZLeB1g1wEjeQREPcbHeY5Wo0h/fT+IbL/QfLree649SiMqBLRdlJ6S0KZaIHRWqSE3NJtr3Fba
vtWzoO17B/cN4NWFOpqhFoMJ3sQqulm/6tutjSiyi31/xutilQN4W4nUMs2+1sYA0n45EnjhSeyq
NoWxZ+F2IKM2BXF0gpaRLI9K/SMe6WhZyVF0D679+h89GdtW0TCy4eGrfKRKgfUe0q7rX+ueBK8H
RcuZyoCMLww6Ev8my9F4lOPeWpYZ/JGomfa8qP4pG+SyzEupOS0VtMaRZOoWTPiGA62CEBG5RXUl
3RE8Na+XKmcX/TNMrbEm/2uu/ecCzjTtquwO01HR6h7w0H81Q0pqdVqxJetYHkLvfd7l591NCSrg
Hfp6Q9TwxKhHzClK8x2a8p7rr0KEaDUUKdSryBbLIm1vN1WyG1dE2fL+R8XRiR4x3J3QQduqo5Rx
mQAqY6fTckOrE/AywSpNUPhltOxYT8cI6KvZJmI/+Wppe+Ioj76u/apqceMLukeE7qC2xQVcyM/s
xpBYThCU+dz5qGT+6/1pPYYrOuwisvIRnZxSXEiUitiMZEgmVMOwaK2rXw95SrK8iv0TsKs5C5Yz
ZWHMJdMte1TrS/61TJvBo0YzzPIrpfPU3aJ0thlCFcBB3EVCymALziP4YbcB6XWUGynV/YUQ8rF5
fOolloSwxRydRisViVQxJpWB9F04bMbeTJSKkg2nf54TlyVNU43HcjFUS6wrW0A+mfKX4inl95IJ
N92VpUUD2HnZWTpWNvb1nBMCX0uQ9vCYTDNANk5Y4gpDThzTqVqKVcphfIol5FJ9h6o7W1JJqUdt
QYkLPjNsBPh5TJXaSzuQs/AlNticXFGm0PHBpaiaZMLzIGmwscT+As0gB1AYTh8hlzq0WpZzdpzX
YmPVOSq1MhvqL4lAEJfi0t7DI7wbNV42Ymj6skiGSXNv1Sd8FEW9FXkQOpTWhBGSLt9upylC1W73
TVZZbXArrGUet9dlKoFM9c5Yp6H9MUBLGOKZOn4ipvb56UM0cCVD8LauviohXFBOPrjwhdVQP1f2
k/kQiSRsAdH4/jV5+QDW9rTsqaRH0l0ix8PzcyUz9BagBPcdotXK3mO4lE+ddUqYcV2CNZhgLMDz
qY3GcSVc1IzD/qPG18Tklnr2l/bXlszhfYSCMMC41a6oS0VVuHEfn0hP/dtQPinNt/ItsBE92MtT
aRM58+Z5RwBSgrYqIy81Uq4LSyLTRf7VXHoXagFvA5QtySnbDtje5DuwNRg3El1F2eBRZcfT3453
Q9yxFUvs7ZOrnyvv2coNRAh0Tjy5FOLUo7u++sOO3hT7sj1tbyV1eSWqZbT4UR9IeUlV5T8118EO
qbL+FilcnELOOSwORfHNXZ6FCdOxBnuRhH+DAdu3t5qQ/fsMkz3eDbMS9x47+Dn4kX7vPhudMjdj
8yncB4o6YvrytHhD/CgcO1m+tMLP9NwplpXBdWE47q5Bgx2bESIGlRAyo+Kxr5Zar7Aa8bTNrhmC
gBcaF2xHHi4vLpyWC4aa+IkJN7m/Wqxn3sL3NRsM9kh/Nf2ArvKGSMZMA8VNmtyCw79GD2zvygwi
brfF5tcJFkIxNzP055Fq/MDqOQLo3AxgMk/mv8emYT7jjBVPkZoWwKTI9nJDs6Hbj26e3iqpdfav
BULBgEIGfhIit5o/4BGkG9ujF2SWyfG/P56AA/bZyVLpfP0i0ee89YWXCj/vbwPkFJMqQhRED1VX
X+fCI3JrYAiUBTzoDbKGi0/kEYsd++9CmG6Wo1JymDbPdbwR+r9MkaWnoihC7Ki4/vcju/7Dx4Su
+OfhRHKl4sHZXaOfhgEU9HVCUC84KPRLI1WiK6RTKh+Uy1QfXG26mvN5xUeuiOVNrglLzXY0axn2
O5JvmJrqJ6vJb8X0sNULf34h6fsndgcXGTH3kOSY4j6nouYKJF5L62aEoarZER+ydDB6xJTXTfyC
Um7hcr2GbSRVawKKoDzFKGblEsEOfa6N/bnkbHAiYsR6pGrv/qIXuf/PRRHamJyp2JaaWFUnw8gF
0cEEE5UYLmHEFfhuz82om9hcw4cjeo7HuTSarc1DWnDEXq3SMuOvxyV+q/QzMtUeqntx2SGtMzgM
oDmEaGxIWZ0/ZotKMA0NaGiZoQxsMBmWkZr2CI1yyRxGbLcY+21OWXcWq3+OmT61kthbNBhTXCoK
PiFijG3metSubq4pAcHCq+YViY6dR2rZTln2xS0+cIMAVMrAINAEk7XAMKUm+IExqkc6QGDZMU+5
fSpwy4oW5PoNPjA0vK0Nz44X0eru2s362wcfyphM14cg3RQLJqkLwi2y6+NfX7yBxEJtjkM63xoJ
NqvnyN/LIliIyBVTnk8oZPGl57EMpRFSuuJ7uIfniobA39QHfJ3TPkPFxyIP+Kynjui+EyjM7uBF
yKbOU0TVE6+pDx5UFdHvZ9y3i36DHWyyaMia7iPfEEunDqGxpsev5q1Uu63maa8P5DZMT6J7sv/f
1a9MOQE1ee7ZXUkbqyvkzrMtXrwnw9K7jZSsSAWAL0T3tqQLa5LpQDGXwqKUWBuMBRLvWh9iX4Hx
tZPrAPp0YQIw/dnvTcqPQIfWVmz8d598Z/d7icHbdVzBA6h9GaFrms1il91UK96I3+GMbjuEq9j/
u7Q2yDSW6xVwcyX0sTzpAdHKo7r8E1yVMZlTDA8qiUyENQkA1hQjmlPrSOeUsDlygtgsyqt3AQuO
U4AiYwkLOQENCSbPbSmZAnMFAnMoa5MDDlGT0/iicdvvsEP/9VGPncXZKohTaBm08ysYUYpiC0rs
cusgc40/qY5yyc7RJnL1R4wCbihjha3+vJJ1MCw7ZtrC7hYwo/zpIBX/HnD7Fg9OmDuJqYpZkSP3
DJ+8x+zPpjHt+Wnhiw9uUhVYe0rJPwMZf8Y0chhNcsJm5HgfPGRRGiPN6nPnKb9LbjUAoAbN/TbL
ijw8eCxnyaJ9fnfgS0209zTD4YKRGd14jzFM0dALMjfhVBHL1LtQIixbQgy3SVMrhAr13lM4oW2u
hH9YeLL3k4l/g//lILVTpr5ro9W6AM9GOc3GJcWgndOrmizjK/jJp1cNREVaMIQpUCUNkbSDlNds
Z7SFWMoBzgwAfxkMBoUMiNgVom3J6eDKJMegH1tBOQotUrw1fXI2IZjpQ2eXwpGBSw/w9WKBdmEn
1GUbnq6k1Nu86w4m+Fe/xyVXhjYA6NvxjP3UZS9e9U3YtM1lub8YgF3SsDW4x3BH+VO67Z7pqI5D
5OKGCWD9PqREvSD0x0cyfKvOiGLMQTwNEa1tHh67fbt67tW8NjPZ0vbTSOHqC4WN2wkQIJ5ASFTc
JwPGpkxfDPuLd+sJo1/Fxzn0kxElpWNYgWyQ0mVYuAKVdBKBnhknEJub85avcUcYKtkGsf9MRXmt
bpg/n2ilUq5AXh+IBydaWul0hXZkA0kbThA5YRtP/SmbpsT7tLAIJBWWfh0JfyA+YjW1SJsdMUZb
3mbWQyVhPdM2jQs8yGYU+rQjZ9jvtdi92gxe1Y1eHYX4hQq32dXfBfRhvfTZPd/zmVSRqG0A42cZ
cAYg/+vt0tzuHS6wgwJM+eSxMbUA1c3OT/uHY6fwrXMbZP+hLE0td3RMwgaLSzqljWn0wwuCOijw
jsqtzQI+2RWJA592DDU6eiVQuTGiu4SKtl6rxW6lUI8Nb1CexAfADdEFW5rsZ6uxDM+DchznNCGZ
yD1PrarVB07wsad7+EVN/8xR/CTSs+oOSFJOGkVS4vLQ+euHNrubvtKWME7kngu+lcY47YGWYIRN
RARYS0O02bmSXVi4tfUqBoGgBuGO1gaz9gaa8yZYRas8l5B5vrDlGAF0hUPqCRlPNSS1Enqguj3F
0cG+qfW7+ASQtJed1g2ug5oD4mOrFcfeV3dOARfYbHD2aoZDnXLYr4S3uD00lmIVMiaAWATtcoV7
mKm5PEioO4alNOJ5FmroLybLJc+4otrJaOfz/eNBKNysWRzbJs6gl2QDP094/NO1kbY2WbSTX1sE
ChspTlC2RzLsjKNrjdVrKVFgO6Tf1PbOR0DQMNRdDewWUxMGJevGOmpc1f6R1Vyv8JOsq3j55AXq
2IJ35HntA6bLbHQeAvUOmIQOH21DRoYrM5fTEZVEzLiRP9Z8mWwW9WtmM9EeRejSmjlqJFqnilxP
TH+fZE0PGlFpfM1m7B5DFryNnlfuJXwnqr0Z3Y6qN8RCaaurnwwnpEVj358yHpbTmeaXqCW2I3TT
NdkQ8IMBGggvFJA6i/LBGGutDrMjUOWCp2VcnPB/pl0U7MFqYH9xRV84OgXx1UIDCsFDnAEGTQbV
sjIZ9PyID1OYyvE4aj4/IjXeWfsJDPlSixHc/FvqkbJVn6FscDnTZfzlYVbqX8IZr2FTjgepDMbC
tsk2x1BMNVLuGrI4Ukt7mM7xXNcy0l4WnLOzMZsUBpWCdyj5gggf8paIHf+riJjlc7fIt1HSrPJH
VuW6SjNkEH0fI+7Q3yx7o09StQzm7vQRy9QX18uUAYgpDz0uKn4inBUuTwyjEObj/yTLs7KpFZGk
otd+wjqruHip+OTvpPEuSpZ8WGpax+hvo+qzsm/qvuziv7WZOdnNiH3wnbbhYS1oIv4wkaYxqF/t
/4e/L7XtHeIJ/WNh9NUeySiWyDehLniFn+uVLJYlv8PAifJtM041uPQ2BT/WuozU66Vrl9g/6tUS
c2oB3kLEjitEQ13Y5QgnszSOo3jJGv2t3sUfNJDtwzfEmAUSmRxsRGid2HqBmbp10u8fpPMQMoZw
kP1TLZjNi1zBUy5ydVEPVKr9sNIMP8MXTnifbWIC0vhjstVpCnQ+S5CKqWfZ+NgG0YXHOCSitewz
h4Crn+og97nzGoqjecaK7QN3JVLIqFUU6rf7tcx9NpNerT8FwOvvOafGK/Lrz/NMxKb0L65qfwbT
MzjNwB4cYoNL6gFRRATJVrKZYGJJQyJ7PJC4HzfUOqwXytUG8bqVPj+8rH8cZUPeGWxzHBpS1Hjs
2IqsE/wlKc5MEf1R6V8+A7vXmZ8HMCqblFtZpUw59wP1W1u8u9468JSbD+X0Bj7CPBOIpxUX6Ykg
vrcsM6yW5K6nGJhy+M6B0iIB97zkMGTN9VY2vOBZpboLam1U08CJeRxF6tXxSnodsebkRVotceIv
FRuhEERJXTOc8CEO+nx36jq+olyjaXlFqj+Do1rea6ce4WqD3kokXIX9i5W1fPRgZl5r1BHWfnJI
HZF8Haek3vlv44T7e0V6e5uWus9oCsojqOKov/IcUHx3b8rflGPnw78xDo1rMbH9xCs/AjjOl6AX
ARtv+BXhyeUANckOnGSSETovE0fYCER74N/ZOOBCQz0v1P94+UPTQI+yf7oc0mFBXG3ELe+isErw
eOLfMW1twfVbOcjfeP97IJJ0CXpyuz1LnzAhi1PaCAJ8pOLgYIbHQMYxdj8Rab633G26OHgbRYae
oAc7EJIBsF7TVB+lb9p+W/bsWJgVw6gBOYo95x5Dku0PKtH61JuGJTxt1IhJiqrl607G3cbU+gYT
802nWaRYbpKsiLfEw5hdHhx3F1yy9BDc9JqrjwNm0NCdj+Tc4AWt78uIKUNE1Y7trC2zjzWLamv8
yYnM1Qdf/PxkVC4xCfxGLxXvXIr0c8xL7Tmrmityk+prBZUq0XveP732ZW9hskvlXEo+zw+p90N/
SbrmujL3xd89cKwBEj3JnG1g54YZFqykkgx457TVH6ay7hnFu/DeewzYJus5U05FbLRNacaE6zmK
WxlnzCs8+E6R5VcU/4kLGsa+Vje+m1hFbxgf4TWKoSfwD5XjeITc4M4uJMSeSqE1pfsc4fOus2S0
1n3HeWl17CABYDeGd3EsF+7loycHWrsqbpuJY0r8rFqKyH8iv3Gze7ndPfiGLdp4UWEVNJuXn1z/
x2sPlbd1oexRQ9+vx/5cnekqtE9CWbZ7QdRt0fBixEAVbN9E2uiQnYCrkwsicDmT3F6nsKd+lCr6
mMYnXPR/BObZByS4PGgEU3eIR2tgdZ+skjM2/QaRfxevCr8JN49+8OUaPNZCex7rM713jmxpQcaZ
hqkCz7IFNA6lhMgnCl6sGZ85KglYFHuXuQumPQ2FwHG+wxKc6p2Yh4mSDkP/8G6phQje1O+lsjyA
0znhpUv5OoRNfMbu34RHxNM+6cp1EP4SlOmVUqdPQACzBpwdaQokjBZqHWqFzpfseHtoOCUor7GE
dtpVj7CnwrCTbr03Xqfd6vqNNRCXnGvaZtnslK3JrkArs4B80ZsR4lMA5sbj0U1NKXBGnbl92ADH
B/NCZl3Jsi0+znK1JiOxH8lRNe6lwk2/ep0KkTzWz5+fmvF8vUetXqnB34ruTYuV0L5i3305j92s
YLuLMnS+TfwLSIkpf97q4Jv6Q20tXlJ2nIM+QlcH79OTvSfBkRnnzFFWO+YpaM+dcA+fuTjbmllS
DuP+MVctFxbYlPiNCFDXwoVPYgQxqrIAn6RR69E03dFfeddoGbcnVDnvaiKbQm8Q00J/1qHghcqz
og98JrOacowAIm9i32+CtYUQxROe06rVH+BVyMH0/TLsta3sYEHBMM+CIjMZDc7kXB2kxGLoNvhZ
GZ1rkxy1/rfzhErDULhPfBhzJ71VI5now/QIyHfj9mXRYb7zh5sgur6iIwmQNk+ktaGXl0+Ridr1
r4O9h1hh4lbie4oKpV4d9eVvTApW1sSTH5t5TeJ44uRgBNwU/+COjkuT97Aw99zEi5UITG50DZqN
ah7VhSA8PZTUdqiei9G0waKw5quIrYL2FraLa4LYiGRF32LPa8vNjpRMxdMPwWZLtGde0f7wK+bO
2AbyqpVFiC3qu1tPGXGm/M+87E38799n6w1GPPd6WqVvmagWAEpB2I6QwNM5RwhgSrlxtT2PW/JA
AsE+o2kpp25KbHyyaorsweP0MKXleQ40qdvhzr8QhgiZLkBb3ZkgYfF1YA5AGDpcCO7ibp21h8qR
AeCJ0QE6NCW2HL0Hk6xH4WlroqJlTLFvApo+JpRsi7RbO3eHQ77niUnsH9HYfVLltYJzsdnCun65
vvZTerFC1mKHGDpAPtExXClhRv8oS3c8ahXiu+nEBG7bRFV70Y/vvr/XPpj1NpVSXom6fP36Kkwe
jUuJXbOxu+CEDg92QI9q13SNjT3B35KIyAFJVZY6EJUOdLuGUyTnwmtlOprCONu16uV1neKqAUxp
V6x1EtblJx+kClJ2PkVAx1YUUcYnCKp74FejsDdReiTe5i2i8zD1jLSzWratLv/kd6c9K186Dczq
UzHjvubtd3ZbMzIOs2J+VYH3dxFfDRzE/5COwkkzkeL7sUtvGgo3pMOamS/vRVDDBvALmNGT8yGX
v069VhadtMJ7SnMajDJkQJse5fC6T2im6qwdECWg6lLlmcxkWla1xiqmfWs2TVyzdj4FJsHu9k6E
Byfhbzn2wnv4gVZSZfMSrIFMw7tqZS83mN12HZcWl5ZzKzqKq8xuv7XitjG/D9hA/3CUQ+fS/fYx
X3it3OjqVeG+nxT2f7wk8lGrTmKiMGSAcCuAwieuBUqPdrU8goyMmNfwBop/GEnAm57gYB7u7eqh
Ni5JcwTZ5XCInC4wwmfGjizntiNLykB533RBKgdmd5WKq53h5MJjctJ+RrP6p26fScnE1yo5YcP4
JfAUOLosdSMXYX/sv2HQj5tmKrnibOwkr+9fW90g2B052D1Qovr8c4IRkOQ6Zrf8kxj5Y4P/imFL
C63eJqEDy+TmZh8dK9X1vgyuim5hrsbwxyaHtx6IzaQOryauzxtY84wL1p223X+33FDxM2usbEkC
a4Gnxz4HuNNkblJhDRApum9SVufVXcBcV2HmU3MFWHUNSl6orKYwgHi8uUiUPb3uFue7x/fIBgaT
60RtupU9INJg/8dHjEWyz+t3Cf5IaBO0b7I7+J+qs2ldXe+yRlj99GffV2pf/0VGiGDlb8LljGdZ
XmWQuXJ+/MVX0qnEbqaHNF/OLUpbXQM8+lhbggWxj6FoXNMOjyW0w/ktu7hBErTQ/hV2uSOOvIkl
Z8sfRPE7SogAft9784PzuoTsKLKJ66fom0WrMyuT6/0r6B7tV/Wmjw5yJ+tyyXThBswjHwE6m7x3
Wqw8KDvat7Q73ryso2QDcB2ulYEsMP5nSNIHqcQiQ5ZBemol2iY0gCi3M850txDRf+VlBA08mdey
mpcIsPnLQKaQHNcuz8XzX7P4S0R4HYWo4lJMgPtl2y6Qn4MJpFBqg1h6H/CLSlq/YApxEFPnh837
WVMsSjkTbX4LZgbMJtdYi1iEOsRCqJADPcBUn/eHQE9HhbvwK2CCxAg+UA/5G25ahqmqccv9rBnT
jU+DAsjB5Kfh1lgeON1G+Ld6Wk1H2XutdPUMu+X0CZa/c29vSvPTNWuGT5LU1tZs4Qdxei0aJVUL
LjgDEDZACH965yt//GnWoE99fPChfR+Fdm4wQR8QVgpMDukZZ1wkSkY77Fz4Sz6BXhmwFBdzo023
ijr0itD0uVzaWL3zxZqD2jtRjD+fgmeq4y+tQ5sCdcnDEabsXh+WZduNUJ9h7yi6E4MUQzH7TkCW
iUHLjcEyc7gv9qLfzOMcuy0fLziZFRdQS/v8k/vQfLOLWVLWj1NHKTsji5Ze5yZI9CFJc6KLbxUC
dy1pfznSizWioJeONAE9B4rJv1zxB0mh3EdMofgTulDOL542qs+pFmqDIIKMpKWM3az5LAYK+kci
YF0lXtXDE1W/NK457bAwN0a8kujQvd01mL4d8g5NPhIcrNOeAOIsbf3MfPsZRUkFx/lr6WDtBHv1
z9704zZgEYJUi8xLHEsuPMgGgPS5IK8M2WWz+SYBzdjF5cH3L2iJzy0+ThTXm7Ke2c8Soyp9STPx
ZGIx1jAKOcUY8IfuLlVmhwFTNOReEtmxr0eO3FJNOw1rQWAjDRruGVpQ1EcNXIFuFEBLk3fulXMs
ysY8bekoi0Mx/6Gnig9FK47eUyrooc0LrFVeqUfSkIKuS540GGWYzDcel74KVQMoYtOLEoGk5zmF
IMFAPk2sCH3RXWl6y/KNYsdBwCRW2RPOxsYSn4oii6Hexe+hINeYHxQGR35b9wy2uFL/zrBs3Ttn
eX8rbZkdctHJBwIsgQ8IhelvEqWeN1V3/m5R4dirietq3/bgl+qVgsIoyKOCav9TH+FZtMpGuqXn
hhfaO/C1FN4KAZCe9FAHU3ONv61VVAMza+HZV227WXYNcR34MHxbEhvDQgdH+eRLpEdGwNY5WBWC
2Vg30KqS6M6O9GxyfSBIrHcj4QRNqqsCtnNrc3R6KHvJaBOvB2sYtDYG5JRK+C18P5GWOHf/MMO/
CAWAOUMQLa48fbe9NXa0upOA99YHLLWztcBIL4rQt8gHga9W1HPBxSTpit7hNlsRkmOI2affKGvF
uaB/RY/tv3yF6NQNOWiV0wXwBDacyMzduVcEw6G0/2V7RfUetcj5h+qVS5c8qowiPqsEB0JOYktC
BgF6I+ZBQhT6MldVSQdj842FURoGXHjaexYQfNGj3fYBrbyFe+igtgVDGcZ2677j1re4+tfddZG0
dOOZ20/JhmplfJP32I7/axnwMGQNwgcYGmCLAf13PzAqvUdYPxu04lG8F7+3U/BUTTWmztoQYIND
Fck0VwD6jCzOoPkL6J9G7JaJiIP5MZNpfh225kVGp4jCaMGXt6pSdqokhUnmBgj54BdZRmOSIto5
fpMM1ORoRxwdnIQXYZx22wqxiyoWt3thniwYjSGor0YKSVARTPc3DBYv66lrULM0jC4DynEfwYAq
t+bg3KTFzgt0B0vXmeFLd0N0mUOftGS0H2EqU05kVwYl5/yvbZYGXAcQM/MunboFHKt2ykAwPMzE
eNzQbLQFaCvzhhjfswSDfMsOwOBs8Hjbi8J1RQ6gVvJbGAXxneWp76aNM6V525XDc8qmCLAthF99
qsly+gB8CdIWfr5epY+oKaj6shqxMFqkrRenl9E/83JRuf+R676v11KNMbXM8UpN408pfHaySEL9
nQlUXht2au+HcfJz9SrrUPNyEfKlSZRxY06In0tPLC+l/+t71ZOOHcC6C8mc5ewWwLwFroVxEDlE
1mLQdQjRty3Mz++hNszSDLbvxXE6lwjO8qdqWUe4GxNg0kNWKoNMSns8OojARyHKfLKSste6A5Af
kkvcsX1TannQajsFF4hFeLk8hOeMYGYgP71yFJ2CutSCgyC9IQFa6zqVGcGvTQT5VZZ7C9oxsMew
mUQ/62ETnFBbCJ5z1/GOCXjxLet9uBLUaPi+cv/xNqvoklIT70aTNwDgNdn9fBpifcr9uo68/baP
nK4exrOh+tKuY43Y5aWCNFEk2KzMKI19aTrkHRUbn54kjUsD4u5L5tJhBrRfD+11URSKyvHd9jdv
Vxji+lUvHt/Dpr1ppyrH2H9QU8g+HVjCd7fM5DpDONPyW4RMIgUtHbbUQqpA5GkcZwcHO/B5UiUP
jWkAWL+QCEJAzHKQbXj0uiq9sJZBzVM6A6VtsQ1nVoNCjx8NtCAsMneF0CwpUTxEoel9efZUumhB
B8znnbLztGk4qBpps2peAThnXrtLeK46T3+Roe0NfahByjWXFrMug7OAfGiDte10ozI1B1PCyi9Q
dsOpAqxi7TeWpE15uMAA9GAMFhOvbJtp+/Punj2a2oC3U25GWPqUsWt3Dqbp6PBQUX6Yxr+LSlIq
3Tf5RG/wnPSzMIlvtXlT5htLIG6NCvHHWhou3cJArkA2g/fs31vrA2w72rPeYpaynywGM8i8Dhbq
5rL0N8HN1M3VUsEVR7+KJPKEaIHKJwnN93kkGzRhUNhHQaVNkN1JaXBQ1qdfCC67rpfh5S+IPqxL
BMkepReVp8LE/XlmC407ysY2Pw6Sb9TLV4c6VHxLT0JgCiSyAM2N3o4g1iZ2dRNzOsSpHgQqCnCf
ZTb/oZVNsXf3SOJJ0kxXzMotnEA8WijXziGUZ3tsCOqLL2u1SrwatxO+JmjP/r+Pi87iuftod+Hh
xcOf89JHCAT9BVzy3tppqpBb5W0lvXSgI7Ilhjctj9i1+LraUfiw3664fDn5QypMTJSnTWdAiTiN
Ecxjc+C/Pc9LXTOSOx3996O+iewvyPOXQq6TcFGTBMgisORZyBqTyyVisA3+vhGJvm//l0fLyZWm
mLJIvSOHyWAvmYGyy4sB71Wev1deUStRm4VMR1qQqTXY5Bto+KileQPuE4uQk3UZHpwxyxLwor52
S5+qbERYce1/gVRkbZ1wGgjjTZ9WQRntGjtlZHttMINFlGBJ7/jPONe1nrDYIYnClNdVreNAYfCJ
PCEcVsqPuDjhsnUisRiB0XVZMFvyrKwfA/YFrYkewU7t8Q59Af9zjCYUwIgtAmziQtKzFEESq8C1
NIfsXBLMNGB79holAqRD+o250Iqez3UASEUt3x7VkG9CpPri/iLpdIrpytsBVf0w76Yess5H7QuL
7dG/s7BccWKRd3WPtC1wiWVDMSANjMQfR4vHEwFErTvZFC9SM3oZVbwQlOVXHXm93fdFFZxd0EnV
wPeKMZgab+nUtEGDH2NvQ5xLpzb+br/e5RVkDFywAnSCS95Gx9OcTbBVlM9gv61iCYE8H6mwMscx
YL1gX0FpA6U/LJggKlX97gfWDgFPIlPHwVR37sPzdgdjp1DXaAFYLDlojaind4p/AiGKbSykhd1p
7mjQh7GveecB3DJBBwhooe+nvrmCqFaKzPmWN+D2CesqLUcp7UWIFeAsZ18Nq46UO+ZaTXoDnBWv
Te7EfiJS2xCiABhmNt3p5WyQyiiT8lBOboFMfNvVNP1/0MxSW8hJb4nYZcv2U+NJQpYih9p0GDOi
PsXW5EnFzv3nAPLIIzmiE2X9osnM57vp7hk9e+MRwPiF0ZyTGHkK0/26s3+atezFrV8FHIeRUm8l
O6oBAD1QUsANQjGaN4Ne2FRPuMOST6E6PVrEiZQNQpp9GbpN+mWhWzs1NVmx8Lmd4NxQW3e2sh34
haIfC7mi+vNWu2ww38osZihtXtnDrVAwXNVMwb3iVDhxyXv99tulyNoOxTLtg40cX9HtEoOK8z2k
IDD7tim9GRPpo0PyjyGIoKi+dFZl41b0jEF4THtfJyaQvyjXp5tJgmCwYSKGtt/4SPpPkE8FVqLS
Ca+CMOYGM7qF07NIrbtKH85NQcoMc0bXOWQ8ZYCLTeypY3KajOhPM+eXjIu2gAxuJKjqvmg5Cxkv
1GbtOKCiIi42O7ObtZpMKgknV8J/1dWdwEMG3iudUDQWGTGnvIMEjjAw6wDZ0v7MU89DHpkUQn+t
zv/1+lDtlKU60jnGo2GFBlaODJ0joDLe2VgY7AvMJTGp4T1MY0OrdM3XQuxumbcmgG52SKuyaemd
k3etlAU+M4lkZ4G5fyD7Zgb3QDVGL7boiG1VcfNPE/wjMAsvdRKScBkOV6YUuEhfikOKcOI2psie
oFdBYsY1NT5w0dTBsnU1ewrlsugrpzsQVBrGaNx9kee/0khVV9jfneJ89J4x8hYhB5QQAanBw7XV
ffnBivZQRoE8zDS4lo6NCMq6PmbeLN47WnC601llsMLsuzc8gSVEE7vWSV6Lub9gO4bRm/30jhIx
y4kJ7XT1oc99NiImfmxTOV6PfkVRmthd1gJOwnpil/NOCORvrR3tjkOlumasd5rR7E95Pf+aznsZ
LxqS3oIKfXaSIM3r64iG0YquL7VH9H161UeZbBYG2V0e5++jsCBZUAedsS1TVmQDGY8+BzIoscN4
U2KRB+fOqLZrSQYHhZ29IHY+01aUHjjr7Mxigxi/yVMk+uSRvYJfCkMGgvC1/fPFc2TYv7gyoWiw
Iho/3IzYmsOdkxj1T/Cl3wVXikAhkkE+CNKmr8X9VbASJxHORUwVzEshpkk6I4NK/yKwt517W7gw
qsBJtOB76hMxjRBCCntCI/388Mr7i0r7ypzl1pbpA8nI8hSKmtILIXdFfKaTJWbJE2ZhKd1kuLdm
HTa06HrxGKrF6HAS48F1b0xFVgQTZ5ekrQQEhL38OxOYLA7J5/Y7yX1SToqfHY/tXoxarnn2ir+e
NhH9MvoZrnxSEqHBIWIG28eq8jD6JRRL+Gbtw1NMreirQpfKAebbZiLdEqZ7hDFETL00XvD3fYaL
CLl3AH6Hjk9tSEf2YUGeVWyOSyNEiZix4jI4hw1Uwr70EZpHPcYwzvaxz9Wl+MU1Nd0sDEeIbi6N
P30Eooam16U9B93WbOety3qyXlLT0jVYuEJaolyYWsyTEm7mE3M3nR4QZMXdl9pGlUcIF7TgVbuY
wjnCJYfVujNZyUd3g4VEMOagJTRU6DN9+0ftAaVrEX8j2d3cw6yQYcPMlGLhCwPXmVesxcMpea1v
HPWgRh04eCYm7cakepOJAWMBExS/b4Nku5yOCHnSKHfd7qNKexEsdU3qZPPypIt4AU1DBJdAZv2b
5Xo5ZTUTM/IcQg7RjUWWoRv/aBnbCU/kocBcJ8Ttv1EDlzyDviAKWr01OAK1YllDuNugUpNgLXn9
BRP6HMlbfM+fIOsIE4q3MOnxge6wj3KPBy9Zjx8bEPxJwPQ1ovS72XekJGe845iryS9S02eV7CiA
zCtAXc36UhZGfAqTWwn+C33QEgqOG3Ow7L8AMVZ888OC65NYcw/lMmImxyIfkCyV3Qz+O+FOh9wM
Kzq8C9UOmmjokAW2MMHeoauu6YcCTj2JUyFzUM1m/paxUPm2GJX9FgVsuRD2juZeK81oOQ4N8K7g
+B6Q0P666WO8iDH4VNspKJfJjA1wJi9px0dIy62KofMFi1ZhOPUdkjxt9IKfJilgbhO34TvqGs63
g3UifzkqrWqKhccZacGLtWKJMt4WRN0KvbfNgluu/M/vmJzDNY4KlN3Eb6BpH4bq99ivhYtNaTvp
WrjZX8qFFuTBS0b6D0KUsYVrSB/IvopAAjACsr02PtZC3PENLnVVCdbaXR0Ox6PKDygb2u+C6r8d
hArD8JYO5X9mZxs7qeQ8G883OwRXfnOROjjUyCWXMDePSvSpNLcHzRiPsJVqd9Xe+jKIola/39rt
VFfyg+75oHVWf6bGZtcR/AySKjCSeHWDiKm06+MtX/xd7V/zWiJNRj1NxREmvZKkXBmI8nm845bq
ZsO2tE1b7It8+JeCIDu+hMZ3bn6DJ2VZs5tZTsvuCUSfQ1MbUlzh8e6vAKYawzDWdrt6fXefW8Kq
RHuaDwo5GzwTGlNbjkhJCoj+RoPv6xnt0omh1ckdfHTAAm0bKzy46+aHY8ov5TYonF95NAR1Ufbs
oluQXWbmwrs8LtERS3LpDmRZ3+m0jPmrmeZDzkZ/tal6PcZDQN/TBpeRg0l13bIBOAcmFjnxzWxW
zdYKGdRMSz2SRa0xhbHO8XkXnEjbw2pvcvv7TDpGwSH8uXQNMflKiU4Oxw0F16Kdh5KEJUiSoalP
P45afets6SGTF6pidLIMlEh4q+Xf1VMBBdn7StO6l9nCrhM1rVFXawX5XuCKLA5VZobYvHxaHRfT
siMLWEwnIbsZF6W4OkYqQWdb5b+d3V61Q4fvFaTCyMYb5gGD7ufA3zkxoWJ6HRbfJMbvT4HZv2Q7
a4lFDk9GufOoz6UJ+/v4BhhwtaEh0xL6I8KTr/hWABLt1m0m9J2J6SnoVkTrknkWFxIZQmkuwYj8
K8VEiJH1ZNnjoEjioL+zNJNvU1nfIySc4POQO+ZUHGbHAhQKA4QS8h6TySa41CiftUs8xRUwzqYt
uHeeU+BHdAMh6alBAn1IZMLM8WcMWTzQ9sdqlldmrNQ1gnoouxgB06APn0TU0GaOlJvPBKw39aOK
uNg1bnR6sFnoa4kvW8vyk5KCtr93SFCYTXM+P3hf8j5z6G74imczls8Sk2jwfqNsI8tk4PozF1Cx
Nhcs5YEBeZFNDT1EjcH9epIGRyWYU194TAkZ9Tp7wn6KUO79thvIt9v/E2NDeRIlB7CJYdxAWEu8
NPxPzz6N4mrXpkS47gKov1+tvJAJoP/izidSl8E8zPTKQ+83v/XPBwpzPRHdGzYvkHMSRqHTqBxX
2vAk2YR8luhz+GnGuv4d5t0pNnqzBF6Ye/vjG4sVH97DFImRxJro37WFyp5T3eyYCnHGqHZPtbGn
2vZ8J5yC6vrV53dnIqRHLGU9hvkKnXxhwwKLRfWAQK7Ug7Im0AypjmY6wTSMGNin6j6LNtO8vxqp
ClS/hguvekpY8oGx7if6yckdSeKZ/uq3MVXOhtl6d4e7E18aqLuGNpYcE6iCXk3VSW8xc1kuDqZ9
KN4dl6JeowEbCqW/bjTuW361XQfUuVKtR/+vC7WRhcopn3svrOqZFsB9u1PON4yC2UDjfYGfPD84
ZwXDznzuqjf5VyOqpFZ76UaW6Cep3O2rycaWCM/5e3WxytzDNUVL3Xldvvk6UgekCIseZKN84c6j
VZOeU9BmafDmnSRM4bLNqeApZV39MPp82F6697aaAM/Jdt+/YV0RN9fNqUKtcPXF96h9EfXikeWH
1fK0fTfPNzVW02958/zAT7AYH0mUl0nac9vRdaUnR7g/57ESIO3dHjhPntRT47rbzbV2Xu2cSmkZ
Q6FxoxI4/hV6ym8aYd0o95DgXP6zlpojiyE2T7oF4lGHAuEmf3OfLvrvr3JHvn4NBE3x+ttqa9L7
IoQXjirxQoGZ+zlOvEzwXyqa/leIme16PT35aGSV8pgHUZJePduG0WDyGfrO14ZhucBP1Rsnaao1
+n2wMj58nIGuakyVs7qT8d/vCMMVhzqKehRxo90yLRdvNCSz99J0EvyW/iK7r04vWYbQR2Zg4iFI
E0sDWYWCGhRdV4wbrbn/L7Rp/0DFDNf3NpuNQbdDaqEEaBskYq3SV4HHTu2KQe4t+igAttZ+903B
yeyj36+lylBxCZMpwQqnLj0E/yHo2+uPRccwpf1Xt4dAdj2+w+Bv2p8OzPJdFLr8PKItqAcPDw/4
8xP8baMlMFNG+znBYnM7CGbmiLPtQZXdr12B8kfmkIB47kZ3gO8+kauZewjUfdUatKzP37ITvXkS
qMueUvvq5L+M8wNdFSIOc2neUJeqqOrSWNRbPpgQCyuj6koV8nBxWA2Fax15U3WPkXC0Hkl2gPFy
fGhEY4hLTwhUVd1xm/cMVUGvGDKAvcMAS4HgqLrp0tQqcjm3QuPyaZ7jwX2APfUHrJjH1355p58Z
OWZttEeyypAFXqv0nSxKc7JiFhSGf56wfS9D0eQU8vjGIRRfm+zYQrHPhAQAHnLKFJuRuzG8xTcy
LMId/nVrRQrtBiNo/FFMsjkV0yQH9gpBPsRBNmO7kZku173QHtpw4FYqcPak8AV1n+zg781zM4ni
mNBgaaxA5JaAd69NBlS/qwYu9DS0IGw7vxhSOM7wMIv0Yn0XsN4y3mCEj0/tmqwTUiPEo0A6xwS/
qaz5o4058s26X9PM9ihLvepbUIv2VTCxSZMZ4DE0bVNvJSBn1Adusw73lGWGd5SR3dC5+9FEL7+7
UECZeIXz8E2YJkzdDEaTRkWuwGX2MLxkyfCrVQOjtBG7PT1iLaWcAa16YQqpdEqk5YQGi6ntY/+m
gulG/5wZsypw86a5L2dvglgnBhntxHe4ndXS3GB51d+oXmqN33gZYhg2U1ShYQ17mTdi9puYnVyD
WylK2PY5qq7oMLj1hSnBy58aj5J9ms9ARIWXb6iJljYysvspewuEWMxwdqFvQR23Jdx5k7plDP3O
iO54v97h+7LbO2w8D8th1ZxgXTiguUXX5eQjcIxzjp9S7rxNYBm5S1ov3OwUhLv1oG6oFHd4/b8t
uNLZE2qn4NNsWWITdamWLLcFByioGAMppogezTxRHG92OJih78oiLHCzOLmDEi8j+YfPSmIS+jfI
YJQsQ26lMTnByM44VuxHfXvQuDZVoY+8BjZL76u/RvqyEOYp9j4hzDtvnIJLHK6ZcnpPcizNrunM
59gHz0O/bjyozw5qjKLlqhoDrcuFQeD9BiF8yJD6wb2ckw/moEQIEK9a/tX5JQr6kMpbLOZDtKSu
KA1nQresYJyV4BgHWkrNBx/AYmkTZS+qLO4SMxCsZ/PrSgYxvc1fzZKHXRAvnPDEXZMYTZNVGHoF
YIkEF2m3jitmxFee2VecROlrxj5Obf/7DnnHu3tJvdCfF07egImBhxjfNx2aylQwOIsxfpXFbaWx
cTBvtv+WfacPlY4K2/wqfssG3ZwUwJ1G/Nd6hRviIYJGhhkBdtBZ+kZvovrUdyz0z/XZvC40P68F
Egu+xQ7Vyufg88Zb1L+RR1uFCWyqAO3fqK4SlVZ+iIdUox5eS6x3nH9oLnoICo8lQHhG6aR/mxON
fqwjJeGtj6QrCWVdUC7loynuyRzs/3XIo2TtuGJyZLgf2g2VRC18Ltv2edL2acDK4pSETY7blNo0
U2aZLAbJbhnLjEsQlxi2UDb//+htR97s+E4uldP+tOUtNW9MC+Pn7qxskmRSHr4g32HVzMpNl8bH
1BPYkfjdIqFlflG4PsC2zgiU5PzKlS20iw5ddllFqeJwxaa8RpsNoZdQruA8WTYTVKKhJ1vVOh2D
HeE2O/btE7P1Kiw5NiecnON7RSmVMrG9mPok+zmKAvouAXmhhu+9GEESsz/VTZ5ZT/jouoF/SF+Z
FXKocH4Q8MXOueh4Fk1Xt3ERzlJRstxvzj75KO88aXbFkpv8gY42x4LXbKmwxLvsJyPcPzzuwcbk
mnYVHzYi0beW1DcrZMgNH8TvfTSDfZYm8es9V4FEAVhmYefm2V/VByvw5d4E+OLMpV16YkDAb/0T
xT1sQ4kglQz6Vq1nZ4nGc6MrBqTUPia1skQmdF/NOiWtv37n6nSrAbTV648KnyFZuKRwvkYsi+yz
cy0tD+yJFd6lwMdQtI2qEkoaJdUPJyaZ8770Su0GeqjgfRCO1i9sW3MtAL6llODIlm+LlP5k+3nb
Nw4Fjw8PJzVWqYDg6MHRwgGM4/RqUn02j2+7UOoJ7E9hUDeVd1wvAIzfvACn3vHyRy5Tvy/NdGS6
vaL4S33pyQ2yB/52+7o3+ei0jMHzN2VDhhbIH4p6mZc/v0Bdxewc2/ezKje/IzOrWcKBi1ySLsyA
4+MX2d2EVXa6VPKDLzKQSGbTCHjd4CDRoXD8VQpO+lnMOPHLto9FGxjumbFk2zd6RIiIb5/KKUBy
P+Uv5xAtfppHMAmgbEU672WZKGQ4VhT7SqR4/LhPIKb3jiKoxG8RN5+TPS3iEfccnowDeV5/3Pyp
/rKbybSnXXJpNr2ooExhMck2IFV4jGkK3oBBYVKVMFw2wkbLFg4y8o2tHSoqv64j87X72ZJs+ESM
0ShGUWYpVq/8wf8N5Uk5gVkqVR+aNx5Pg4+5EnSo+49MOgL5CvBLVeCKXetpjs6DXLiI72qO7xtj
dnTBR37v7r0Of9Z3BDCLdaeKqHGlV6DcGJsws5UQP/kNhEQrWn4N/WmMuPrGFzjc4W+pQLnFg5Cb
JONNFtUp4cBhJVpRLHd47HMEOv5rdb6PeHktk2/my2i189uO/IQf0G3MxyNImHMxBGplJkL5ZoVH
iPxASeVcPglvYcl5VLkwqG2FbbaKU4Rh/s5C6q9fuz5DNTkvyiVMUHWNl90rf/TMJ73WzX4Dp+v+
T6qNRQuVvvsbmnFd8sjLidj8DWx8x9Ygp0MgxSoxfqBb1h1fK5LTIPtH7CgUz55iuUlVJGIDzNqm
M91E9/UUIRabk97wpufQgvbe0iv0EmVmflh8fN+BsBCbw5loj57GzuPQnv/FG4Vo6ZmDYHvpMghE
caAh83f4fhsCNGEM4x6rKs+k4xIU7GMQjByNjHVsTtFRShnU2tXcdcQf3K+oej8F/nhf0wi33i0i
Q0vVGG2Cf0eebmNdc7STY0/afBkN8SDTS/Rmu48jkpBnukNlr2QmbpUyGH17HJkx0m8F86GE7oM+
g1h3SmTYvIwwGg3jEiiyDQD15sS6xUKCHvCnNPHiOogAA5zMux+AXPo6SJhL1DRIOy0BBMjA4AxA
RVLM6oqCvFthjEuIbfU60j4DwS21EYuX+rkawn8sw2VhSKWS78oMHdmYhU8yPDQ/5t7VTCz+avWj
wZ5K08jZQVfnQqMQcNxK0sTIEufJKt4M0THX/dIDJ2iKLiNt3wPiut7hFfVik5kEnUIryyKbUjyA
tNbikXt/4JDDMWyAr0RVqvmQJOWXDpIgDsYsn80qZ+/Gov3+3ZnYvfQBu7l0Z4n4SeruJdTsnpBS
NYiVZpmSigPdMfySZggCS3iUhuEzNzYpAmbawcrr01Ngho6uhTanr4ehrWeQbom8cs3I5Gory769
ke/zWxT5dhXk/lYha4dY6OJzF9N2veulqq7e3B/sc0RtTkG1HN+6f5FpppQJThlMVjaxwzb1NGt5
3lBZXnGh2bQH3pugHdrEkKra3jpadNxm8iB8lHdSXJAAWyWxVXygjBhULCam/P+2E5loHCRAVwMr
88uVTNgtcamcwuQPJ1tQd9tnCzjkku+1FGBJtCJTBqINWrrOY4miLc+fqa8BTAQ7a2g9sI985OFa
tKXtadDha9rDivnXaKziFsTQr0/g0ad9oj8HcRwBDmEgbd2lkfxIpxj0ucTNMH6BcySPeOJnm+qe
MSvXRlZg8lnRRVj73G6erwMCzBf3wz++uw+cgH8WGlnzYZHD8dQP7YXc2O5e5/ZOYdnH2EzLI47L
44rQZk3e2XyyddNh9hnVm3Jagj8UjmpYOFEVyk8AQ0kfaSBFM1Z/2UifCJvWLVNqDSjEBUzrBEFZ
YkOARc7KIfIr5ht1vzIOiO1XfURbKZeLxv5/JPvqI3E0sRBgQXKzTs9ogzigxm4BTijsTYIjrRTG
gpN/Q55VdXrCW8IDL0eJ2NCfNsCvDyZzVjMI7bmfy8YnP/Ht80pRRr81ul1A1QlzUzvITsVvNjkl
ucTz7l3lTr0suk+4UTnU7Yxwuo8AMje2cZl/8lItCTiw3rCAsXGNV6fDsEHVy7dgcTSASSo9HJc9
bW5GnHwxoNdxIRKiDYL+NaRXOouTtd/HITLhDP/58tM6Tcqj9DRbKYit7b47IAGixZkpokPs/ZFT
hIBUwaJtsN7CbhBHXibU/DQkQd302j89HGhlb9IU0BBKeAo0+sV2njti1sU+pqIFdfdgKGigTk6x
cIHxpAKBVqyYZwPwu3XqGR5QjbxtwVgT27DyjJAM1RrpJlVrNc8ppcRvDkPE+BA9OQHXWXVy7qOI
lHZ+cteL3zSKK0Hc+h7X+JuIiM3C9PauSjlJMEM2fenvSM3NVJBO0i6bgG8MMe/tpBUZEBmBFoxQ
m+1Nm023T0E5EPZkr2bJ0WmuOES1C/pMUxAN/NbFyKlVooWRE+nT8eTUN/soj880VmaMRwIuKXka
ItbNry10u+S81m05gncqycDSHivu8upjrbZEX1uSpqiFwWqMSuooqhhYN+VEdHT8oXMqPzcBly+K
DsEeoXYz4rUf4jA+dZjR1cvKv7l1fmhKyRy5WK67Yp6/2NZOJ5qmunSPDeXD5Jojfgzpz5Ty7i8v
cgjAahzC7pCXIWHkNbOJN4t+4+KmF980BTx3h0Uidgi3nP8eTbVIlhPtIuaHf3srsth4SEfoHaHC
Ryu26BHCboJY5Ud58lvNCQC6/fopuNSMNsxFJiz/3OEDVsiQ9BUFNIYGNBUZT98xRghAErWWOl+U
3qJw17+SYg7wKa+XSCiCaBW93BuIhfaRUoqYyv2ez0XXuIu5sHeHgmdvVsC25AKKaBqyJSwZrJHw
fZKI86UiRAl5Vi2RI1dU3s3fR23ji1+n4dohRy4pb+c73TMywsY4zIJaHenPO3n0wtm2vBk8qL8a
7twO1L5o50Y45UjznnPlFcqJ7ejvfhKriUs6J0shLabcgRPUtNXEh9YvQUrznAALowQr0SC2QdoF
V5kHb6gS37J3eA7zuLZCODjJzYnM+AeJyEjK71HRqFTsmUVA+3uUgtrjTl6oZoy8cFdz8MqAlomm
Ozi4LiX7F5ZtGCeDAqQsBIpRfXi5wFQFH1rp9Wo9NPRG+5aFojJ/M2v0m3XaBEklNzZr3PHKXSQA
QlPu0me/31MM1O7iXNe7MUtcpe+IXjaZygL2vdVcLeyl0VslKVrP35/eQdH6vIaXQcNd1aExMVz9
aPTk8+YKpghK/XOp53llf2rtToqd/E5GhtSn7lMqbEpy83zgO5DvZ/Rzq89RwGIWKsqC26hNWHWX
uNaLkrxbWiIwIwrmQUaCkn8ejtGFO8+D38rm1JDWOzyKGO8etnl45NzaFuv3vh9LGp539w0C+Xil
dpbiEwMKpXgyUWpoZd5m3czBeCF7IoCkI4v/r1HfX11IgncAm7J1/+lqnetQZYj5EhhJp9gGuuyu
nosrmlNlBueBSSW3tc6Y+nl97q4tYHhDvlPOsE/PZk2LJfxIc1XO5BqAfypjmVmwqUFjNNSdNUOP
XsCNgjr0YZQ5ctOYVwWEZK/JjtDZsLhV3s1oQdeK6tfrZfe/cQ2m+UblnTwjdmAKiVu9p8pV4aAO
bnBd3t2uL97zq97xg20DwDEL0aGmHubIzqTq4ccSq72YHB/GOG5M+7PWbXZWpKH7TTkfliMgRSkN
AxLqXFIMu7WtLPVaFf2fCr4bXrtmYeFWQ5gnWOvgZVGP5iqUII/N0tZB/v4xquJ1UHGh7203bOU9
MfyPqgI8UXhyPPPfGGQLJW6o86rfABo3QMvtaCYZ578bozbnteDLHBXaI17FW0o1UKNVaCw+RCjf
Xe8Q3NiOCw2Fpcg17J9qVKm2lIrJ4O3IlB0pjBl+5YH4qc5peRH/95vAvdlmExtEdXmIcT+fFwdG
esCmj1adwG+CcZjlBYBTLNaqoZ+Tn8Hm23MP+yE4RtvxGz7kDICh+xHkpMtkuFgRuWNW6NxQYtlu
lUIj9ojiy7R013HrdboZTvImpkyBSr5YOloAyUyqv2ERDmfvFzsu3tSYHSe9uyI7kvlELfggw/SN
cUSjLb+sRXQZ+W3/puhjkhWZqEEUERchj+qRa+c2Zw3bFBQkLYth9IwHoPWZSeKOC7IYBCaKUlTe
2JF8OfgeqbLNytk5db5hyKWMLXSWxX8oqGsgck1AoZbbwEv+Fwhh0rMcVIRyEwPtif8jGYqnLABZ
GhKB7g3PvOHpIWPy49xWsD4tnojO0gmkSw1LZPRR8pEM32w+o1D8nh7kR2BiQIPkl1Dbk2M7s0gn
uwuXzJlfGFLDgAEBGjFhjOz1WMhXtMqlNLdzGPTobXFn7XdhPZq5yZwzbcGz6OG+ryv2P6x/4ny+
2YyjHs7P1dTwudmMO9/sXeBxvY9finkL+WbRR7HN3YsUzcD/N7IWS/pLPT/WWdeIOkwRoWOyKd7A
iUgbBb4sRJdtx4y74AeB04Hwt3dgcjmXN3hml1fZgAOKjH07TPbctQfswM/dkjbiiKha9x7xwhPg
3TNhJUlg3IPwdWS/1/UghmmNg89CnaEzVzxT8zrDIKaOJg61Tb+Bk2JvqDa8Bity9tBmTCNyUlla
dLoSxsk3dMxfOD/1G6K0kcDOoUkBtfDWNjj6zRmQrxeFKQ4vp0tIHna6hIwJB6fzBPLqt0lcFeb9
p4swerlaW9uGNQZOc0J/MOSjfCr2LTGHUxXhOcznC4c7s6MvboqBjnb/fojbL4wXr7o0fxXYUGxG
S4IL2/x7BZA1yGYyr9PMbwbex6Kn5B9CEqMEaT6LLZxsa7mYWy+a3vzTwawe0TDZJqK+xtclS4+i
vFDfSQBZihwfshNrTpIgSIF33eY260T6XKwe1BqAmfcLxxUHrdbrAR9e1znrAfUFrQm5AH+xL23D
vc4KiA8R43bZo6d/G+a3sGu+BlHy7+w+RUJkCl0YwtNKjwWvLX4UI4mHG7PQg6sITsjEWtWBwTbX
eC4pjfGfMbbBEBSdN4C31YSu19Gqs4W2obchtJUqRLOjA4wkgFaiCf4dxD+Uqm54PGTgg5ur136C
CeOVI8wbvX1PGZZwxprIifbcyeaYZ/WZf/qTb7fl+ca62Awd9qv492nTgJQUw519DHaYZAxKMK8y
iWVaNmX6lWvFlCoiJHWaxsUjh7FBhf7nRBOtCaJ44m2QsKalYqlS8VKuqzNq0poE1PToIiW1TGVa
2Oasl+bYvUBWShh//kHKnIVLpvljG1/1rFoeoaf7GmdNPzM4XKdmWKYFAQ+9sRZfdj3IZ11jw2q/
Jnyyve/IlPeNnUwbPhvHuKa3gzyJ73ySoN+ietl45RlbeFxxzhvh2bnnLr6eRwBhhNJq/ZU1uV0c
kz9p+FGX4Ma8J4ZbSe5JLQJZQaJjth1rBQp0KWHCTTcHQY63uswyopUIsIdFBhTPJ/zJk+EqRuWA
Mz81Ce+IwsODsEZGApCgwdDCQuFfBKacE+iCDccg0aC3y1wZxvUH9y4QPdSr0hCZlwVsB+vGm4AX
Q7sldF7zBZixTXYqZlnn0H2g8nCp1r0V9hgtmWAoaj5k1Jt6mA/UKnnP082N13vUWpmmsnDs1Xqn
Mfc2NqsZGBlQHG2vvDrWUA02LsLbLh5lLitpoYBIASdCynXNZu1ip+NzLHbXbqStkVl0GIv+mz+B
kb9htRLRdmsNfFtunihKe93C8OMDiIkHXB29fwHwOAv0YzxWi+K/DRedGTk8TBshOW1VQ1bv4yPv
wyBjjAhg5AFKpXavY4Tob/rgnh04XvaQkG8yMv5w28NotslL3m1W8Df7pJSLZsDsYlC6JDJaapyP
JJLxxp35NUhnTN3Q2S3SvJh75bBZg+7nSMtzjRoVfykax9kdXZ7pEsTijuQUw6ADS/bXUUp6KXOB
IXjjxCiZbw57rmqXbfklMAfbmv6Ej2HYZ3Ps1pkD9uG96YLZ2QB3fzH0fTc/tSZ8P+zKKSZekrR6
u25pdekHyrYOcsp5qdYGZQ3708lZcMqpDpuRTPe2YGbka/xUDrOh9VxaAqMk0V4cv4skreMLMdj1
ZlF3viWLbwYYnUxlBVqkm3Q7CigYAsfGs3kVl8gyz1ftXQS0FD655pXBRkpBLPMQf9D4z9En8Mzp
qGNg2AEAWoEV8kqaZCeJ+ROz2ILViy3oTTV0/5Z7rSIiuBaptoJrynR5UohqlrZBRgcxT8AMSlwY
G14osas6Ii6SA/cjUG1sXPKUD6Xb9oqorBIZCLsdyPrEwghYjs1YOHXBVPm6P2srHNW+hyzhhZHu
I0Do7f4WCWC+wnwaTlm54PFGeiUMcUBtyQbuYFs3ZBvRbuWgCWo1Rie0UFMqKU4vYHXbMkr4qzc1
nW7Hg7+1lbSFY1C625mw1ARRrcqJ0Q+06S27zQnBLxQi1oflK2n+p0sgjc9EWZh1zsnIX81Psbz2
jS/WwAtLrcH94ITuUlFxmZr0Yu5or1icMdKInmcaqIJd5y6TYCClO/Wa7GjZXWqkyaN4qS5RmuxA
yMJmXqgd36K3tSTqWzJmF4vuV56jqDMm2lyeIWfBqfdKX75FRweEtyg1b8fHaU/Ad9FmlJWHx5Yl
KRdZ4iwMrfJKBzunPx6sBTOpLu1i1IxgLgC0dx7+S9iYb/felXuclNo5BdeXx4FAt+4AlJW8jDg7
Kk0SscEvq1CtCyHUEzd0wateCrHaEJwWFLHRwkyqhMcNb9I4Kh88X0v1KFwP9fCAv81YOWzQ7OJR
FJxB9akGjUmuEostpyEhGR8VQqAyA/cjV4+5aZIEKHLQBaLotEtU66WjvJkbG+l2tOzmpgG/spk0
alSQhiIHaINQt60fDvKVM9IoWTS2CzAey4p9ZJBJKLD1EC09U4/ZCQMIeMrgSUhTyg/2ytTx5Tuo
cT/91G7VWABU6q+M1gRfbKRc2Uo3reuQZzIiXUdUihKxzeC13mVHjWMVQ02r5e5tKplX2mmwDhFQ
igH07tWNCf2rKkKmB+BRHdwq3ktQqb/0rgqYmU0eM8UO1ZzHVz05PwRSKq95T3ZQFCvrczoac1P1
2lJ0BnGvioo7yCbn9Q7NNJtFqJSn7qRggqcQ6aNHp0KTciMfg+LIIFfvfMku4pRiJc0W/e+S7DNU
58i42SdIR+KbhxdUQ0FszPv6z/pmrdlskQSgAIB3dNY0Vq2ag5IkeIQeq5s1J2sdEc7L+dUo799/
/Y+AcdJJw1L1XPE3OqIRuerOw+xWIuIly7CTI1+1BX//1toaQDHkbvm7dRP2ZkC1ZEzf4Ij9rM+4
BuowYf5V/urSqSD4IWt0KnmW3mn14lAyqwRk29ZVGRpbOUf1M+K55ujJtqSVxHutWSAKTwgeN8hv
S2J0ez4ExoIZLdWmGvhFpp2FeBB7+tjXFM1zNBLjVcRnT2RU5tqlNjJl9+70a4pTiO94FifCnNzj
+R+q37V9P92NnzebSGBeeNMU/jT5kSobBH/4dG9N4eMyk1GuviEq2BBIER+b+nGIs/50OKvI3O3d
Tyqc8EothqyW/I8R0mzW3Np5Xpv6BATqp/7E0WbNVy9Pfxf8NyiX5med3k5DA2hssXq1N+KijDy1
QSP2io51jCKw4CyMpHrsPESECmPvZYZFzBr/1qonFE7YgUuFA1SB+uNu+z5SGhb1RrX+cDhhimPH
ri/BviIAN1J5CQQRIH5bRrb2EwD0uXurmFj0u+oDk+YVhGwcQxDLu9J+ttmQkJSWyuimketaQLlc
m/LJEz85LYEoQrQn7jOYJIbEXNfmpb2F1XgQDjse1ijuPclh+YGEcNiGfFZaBKzZBMcEIcMD1Cht
HBg5Or2wvrwWSgD2K8bkAR00k8zAdDHD7Wb+xigTaQXqs6cfydiaJTZ9SbXzU4iqcHtFVGF/Cy99
9SgBANdjMyrCFeD0WcdVTlSgTqGtVxEG1B+HOHGj6xH/3h7jB2vDBX41zN3a7M9jNr+E3cNCBmT0
xwuKM8PlKj+uT3jK5zm4PZCPv8hO0WnB/rwqJvglwqNzHGOKJg5wdKJPnVtxHKE5SJHhL5LN0O/3
eqyQGdCIVTtMO24ffker11moYOREaIvyqRoSRqT6SeQcO+/TX65OqexXw4xWEL2McocRbu/NWsat
LhQOZHuL+i8ScQBPXo/ECrf47TAE9XLAYG9Aat/8PqCpkT4NxVF8U9Srnuc5V/M7AGbVQZufITfE
+vRRYaFQj+danD1Y9OyzEm3F8FbDHSvk3VI1c164Azg1aYYQhYcIKGGJEilx7w+FtJdojVuxY8Tv
7gN+viXq6SiribkSYodb38vDBN9nShCYdl22TuJUymLnM9KX8IwLQaCqVLgwpQRBiRdJwH0wPDny
6sjyfx31x5p9roX9R9RpZTy5q183tGeKwxPA1mMKhBGJ1prA3TqXebuaHntc3Csb6VBNaezifD8d
MJuB4Jj8qQd6zee8oIqZNmYesP6fPPg6/4YKn3q7iz/CU6MhmfH+nOdMXZdMDqkXdGoAX5NVn05l
qodbUiE78DD0gjNfqJ4V05fG6WSRCilUi7hRuoi2DojQ97LatG+rYiwuXo2WTpHru8RhNoOH1yKQ
Rk3ZAiNHgz8H14bGmBuCykjM3G0Ng26NOa64NECZI8gACnNyXVftN22ZMVpFRfVx8y4aNt6jjtGF
VNelhyE58PDKUpKWcR3O5OL6VJPugaXk0UPFYo713XMW5PZJclIu4fq/bZaqDV3tRNvhpQKUI3AB
HmzP/0ydPeVDVU2dvs/zCj60vEqXbtkLQqiIIB2RLBHq6KYZ2UFnKlN1QrOriK2yoG+R/y8ND2VO
EQbgxxupfX966yXx4sryOCF6TehZawsK2LIYLHiwJOMYJCKJiR1eO/Wk58qA86l65RYwGGZrs2GG
D6W/3ATvLLXUoBuTm8qfPjjkT0bC7wtJik/yRqA9Y1R9zVm+cIVyOHEClZYpBJzBv5hlWGir7REv
TKysclxLWEthdBKo6TfF25kdrCV3mM+VGBlDOf+Q5fWRjAhJfAeZxk2KE4asYDe84VI7pMTSj1x2
n3vjivdaMDfnzMAEz1mKfOE3pkJk3TdL/0Oe6H6XWQ209wCOcDTVMWQXPpsvAZYBXNefadKn0PcN
OBbWLCMD4XMAcwYmm6F/Co+BvEPrbFTYNiykbevRVqeDS0bMV9eJMFK3wRhrjsvd4ZtGQJSQbEyM
BnYU5qAbGhM0RcXT113d5oetA7eMyZEMLu47gbZCSunrPdR/pyx2tSZdUxmot3U7Mmq06V0lkPG9
WYYOSiLPBbuHysu+AMWmN6mSRG6DKw/CzzGHCIzWvDIMRdqOTUpDizrn+Rp/0rdCXqR6I+3kSnLR
F1P4gObNwFnoGNQNqyYum3ikMNrbpSqBhN6qRn5DRZfuEJUEqmHFjnm3aF+00uVy8qOH2oH8gNdX
17vBCGuX0xA6+gRxzyy3VudT8X7AMlSf2FBFFS1BpTV6n3G7pbjMe1iErDKEkmUtaPZvC1OUGOwF
6UxKisgMYDVioNoBkq/1QtnuhHkbHZSvkVf0PKK6iYLKAYxPZ39eOjADUHI0iF/k7lSJkDzY/X6I
iqsMNHtTAe8l4c8WTuvG00bWaP0VFf24+HWu2keLZj+shrVBwQLLpEDn4QcLh2ZtESL+pv+jjW20
nc3MCHry/B8VFbs4c/IUa7TQLyen60ZfvsefYCVVuH3QapjnKu+KsPmpMFVLYb4l0CiZ0bCG57ll
nzMNVJGswQz5Bnxs1PdGYFLrHWg2OmAgiH3UfAW2VOfvpre8A+7kmV9u/9hrJtDGW0cg+AM2YE+L
Q/gt1hIXJwS3D65Z536WJYz0p7LwqGNtRV+ASMMG8CaKjKsKtMwQz9xPoRPk9Mvvvqi+oOk4J7NZ
aUWU+iX8stU/feiALewqnA8lauLZENLeJW0QwZRTqu31tIdEY7WVQ4ofZ8nxi6/WvbkgcylSPXq4
nd87MrqBp78Dl/f9Zj6rgNoqZDqp+RsvYVv0sUA8c2AkQBaIUvHIkarfNHfNmthmCMrKktyVhxtz
eRpmYNT0jGnJlbJAt+N1roQLu6GWrCPpujBH0GmeeqksR4111YTyJS6gB3vXAkczp0iDmH82C34b
SH+iuc5Rdvrn33W62Jlp+OYJUZ05e0ZtT9h3bYSwmPH9LCKaUYUKliFcsXiRlj1BqxprT+DWqBel
rB4ExEpq766ru1mo1Zr8iTHXOcopDQ+ZzhV/w072Z1sRCdMnaMptxJ7cQQdUG49UhXn+1c3Ayq7t
OOGDwNTb/4nQQqw0zj1iJ8237ANwqT4sdxe3x0fCN4oOU8ZNsgzvDQDHAlJ4b6LPkbfmVYO3XkjB
SRLP2rgk6I6KKL2EwCyNuTKuBnWQuFwbsGV0Rc0rx7NU3zKThI87lhPavP/4CiX5Mu+sIh6YqKYl
0W2ovnTDkVwTQiU9Qi5Ts3Wg4YAbql/LGNU5aibtEznuKW6KiWbFzu9J3BE9RkijZb1Qs/YGc0gt
D32frhaOm4iTZlB5aVLp5TVDUXbiuTCDjNDMW/XYB8ig+KlbIblgrOOjo2FjggSE7Ja1TxA2SSqV
abUqnOyE+Rfw8BgDwKojz9hcu0bDL4D5/Q8YzVAV3AgoGyB+n1gEzCGBJnBeVYWNB+6IHrhPQAaV
kfDVqBKK0enpoZkBDlhNRsqscXS6upSdW768Jmxt7D5mw6MmnvjLh6Ke9yFPFAszh+2WWs2jcXWd
mh0GnUSTsQsQ/4c/JzkNQAUnLfE5B31mqkD2cqKAO0FVa9dhKIedNfqAlXfosvQ2GoK8sY569Whp
WkLwSx9J8UqcXHHPvhN6iECAMbRBtcvUr81AtJuvA2OO3iguNyOArzjufM2hJD3Vqvzt9olpWt/P
4mV/opjHjmJRQDpUV+RtFnOuz43RcvVzs9z+JI0R0MNto6z0Ns8hQBYaU5bfmLTRQ75wOgamejcj
hukR+bbZZriYVCzMLcYoJbDYjfs3KTkPoBZpri7rmmT5wyOGCuPA2fhl3WTjQyw8vffICvs94BEl
ZtFRA9Ue0lOj5xIFwRl/fnGdKMaOdsw1G3wZ1rWlLTG/CazlwtP68i9OcGhLvQB6h4mTl1PfzAqM
C4aa55qAkG8XdGU38ziQZ63llN96lbuVm6R5zeHAtOupv4kdBHAuMFT0fldl5yHiLuRruAQ+E7JC
9lEIUJbR+OYqLaq8jkONn2v04i9doxskUAsDP6/dW8xIPJ09SnCkd/Bighd0+cL2li1GgwLiCL1X
yToK1ehchDjIGpLxYHjtSJFFqy1D5uf9daTZz/YKLMWE2U5PdKwG0lC659jaoaiu8lRTaNR57+4Q
1EspLVa0JbWDjnnGxu1FS49N1jvQ1beIgEoI8EXKgrJ/nT+Lea3tauhZWpTvAhd+UUEfvdwhGmBJ
lOEiEDydSCkoti6FkT05wK2Cp90iC8/sTLraIsYAcjvgla8QeROOvETAvf7gNP+ZvDQqjlhUhKfZ
NyodGr39jimKmz1PFfu+0XOoaAqdqg2ahJQpiTJveRoz4SG52wwQvIzexYnRh41bD+zAKEFTX/uU
a6XPi9sFd//hakWFKh5+cFccqP4kTabrjOlGEmge46D84ILIV0GNYZbFbdbCnfxtJu9gL9Jp+SFp
n9xliBWHIZZHSnAr3oD7mZmbRysf//Y6JNs6m8OHVLZ4uZBkcA+lUqaNRgpnMJRjrmsiReZuJlm2
59AzXBwMtIa5ui/cPAwLJMDXQ/FXqN0bo/9hT6Txc1PrcUowmk0+ih5S5PsWBk6wx9wWF1DJcBQa
lYOibLYqa3YASXT25xWXXSAB82eS84SUjTwGf1FVHFbRAx4g+6jyC/OrBIzZk38hZlFywe01nU3h
4co7OqxdvQAufE3Kxg78gb2sAQlUPVXCR24XHbNwH7nbkeuStj6fkl6zunogx7HC4MeGnr29wkXn
t8Q+S6fF0abV9DO1akbNvFLbrLuYUdLCq/suM0KopIqAnulNwQp5+vCEWZlUuv0Zoq+nebv8EGD2
Sye0s+exg56pMKnnplBTUaWJS+aKsAC2LDtF/DAuUSJvgAj+rSnjf5crmmP3LyT1poMxbxAiw887
7tTNA4rzWUNT4JG2j0jQFNbOxlnzqhCb7Yq+5lLd2lPfJxYdhR/wcaYmvJTZDd4eoJYKc+y9O0cJ
E/BRWstfSvmRcBHcl0FW/Kf4A+jw7vmlPwWol2/zKSfa3G0y7M++AR75ApeVfm5wmwKfox+/8kHa
LTkTo3dgdZFpqbxrh1Ly7KA6Pe0hNtO3/8ZzovDY7tHip8zjsBDPCc1vwgUuMv9LhIP0COFGu1IB
H/gbv1qjLNHOCsz7t1Op/yT2YIRMSiTb0pqd+xrqWQ+7ju6b+jjovJU8CTA1TViku/8CX6V6hk0C
ArmXMPz0Nh/uQts3ROotm9a7sBjgMQPE/pHvEPA7hffe16rVLhADOqKuakoXuQH1/zE/Blzy/WIt
ZDz1Fp3ZFix2XetCJlTVdeI/vCbl+6fmuL2jQwKCzEUBCcaDVH0vU9/pILDGy/OcBA2vrmsnhYi1
aVrld1PCllH9EX4VYe6GgMw72NCETRqYlA7W0QL9O9Ybt1mnTek1Zfst2GOWoegnyWuaIhFZ6zqe
ancC2MU7KY9oqXklG/lhr20MluM7Kc81Ma/SB9sDnIWMaJpmOLi5unhZCqCK6dl4/aYN1ORDRzDU
+2b335T+WwspjijGeYTCJxReIbLB0OXKO+ADiIsd4VvracUenU36tE3zy/flCONjAB/mpv0IbKRN
lE5XFXwrzNoOaVOrDN9vjehv3QwuLbhP1vv6UU2ekVP0DN+WlcZYLbdvZ0oFPax7kpoXc9qValIm
n5ZW3rpyPC1TQzKi1KUS6fO0jiu5zRWz1a0cooIMzuy6afBobCeKo150RqRmodJMbiwwV9GE/ckO
GHK2E7U5oJ1rgc7pCqrTxOH7fMj1KhluM6xrwOecf/BmmsI6Kc1R9OqLNV60EiwueEI7IDKkUDab
x3dXn4r2NB0Y82gea0cmumCUP7J1ubquboK/2c4vXxjSaugkm5+av2XC8X/0rT9+6QuhSo3dbeUt
KNkfEdVW0TidJFWqwtY7C8EsEQ17OlMOl3qG06BWiYPlgvZZBji/aeLqVH6wefwruSRnXSSioGhm
8i0KwjMH48p/LZByZ3SXknCTMGhwSjdt+Rhm6Qlmkryxmse2+cQ+3J2sWdknLhBVMuFI1y51HGj6
VUvm2VV90fa7p1F224ywQ3Uo7XCpnrnBW0G03PFm6n7qTy920Y1mpQuY1/FCgLPWOyzxF+rxIhzh
k0PDSwBTL8j/VoR5wMTb8oJCODaYQ838V50sE0y3kXz7O3p3cAoZUr2tK9RE/tSPJWekzjXn1s/s
rZlqL7AJM2NiIJvlYp1NDuYPRzChOVG7cmwRq+nZl2YJgen6Xngrmn0qXl69aq/CI0zeKdTuN9lo
FWD228KfV8Ra2M87I7Zb6FeR5rlOiY3tHkJDMkr7yfPhLfrAzeNVeA/EM/h5pS/q62BOyUxTT6n0
LEHsrALWo2mFlNpUhHtrIuElgOLFRWumSBosEqnHS1hEMs8+zsMmc076PeM5fG3KOGV1Xk2V3eAD
Wj6narwN6+nAh0spPq6PiWCo3rkzVB8DXE18zadtc5WPlySkH1AvdFzzbQl1A1DNy/yuDsRBCeae
YVxN8tSLuhCnBI/XLYYv4BmvP4Q6s/acBxIAhUA8Mlz9G2RkBmFmNChBQj3h0m2oO0c/8aPAMFle
3XJQUJ5/3K6Z/+EJ4l6DhUASjST8lquBGr07632GbMPpzGjTztXQlJdg7n+fN6KlpDXAIJpAEjVl
3OXQOOZtpopluugyL859swSKFF0kXTSy2M0LE3sDVOaQtQLetMYhQhaO2+lrFVz/9sdeZARMTMj+
1AL9eoT1XktV+SeeruwzzpNmTI6sW+Lv1WpSdkfXbyWSw7dhlKIlt/Su1cGLtLgKP13oF8a9r3tQ
NVA0/DXKBzxHg+yEDmKVY9s8Gi2I9fLSqPSsBQOHnqvmuVhn/pzPkSvgIvGI4/QMqb63aadY14n+
gvbw+pd8nxVhu50jxuvy5w6enc7V1PJ+tjdLW1AhJNyhXlPAudisRtsoJQGG1ixbP2kymwW/2Dwo
mZQnTH9ajIV1zX9rYiWX5ADdClhF50cWK+tlkvloy6RRm2oYc9OUiW8YFSzogf1AM6gX+nLvsdo9
a8vdLOk85BweftjS6BA+zVFFU+nZev+09LRIkDnyt6V6St9zqld0jhaL/1bjEMX9/22s7sT8MkRx
EHBTyNgzO5h7S8OSa6B+aYV8UaHORp+gFzQVqbCkPSW7HkW9O/6KDWcqORSa3SblsPEjvfog2nAN
uJwsygJ0QfiakEnKe5Ag8xgfLkcEj+j1lVcMoNgtzRsl8ui1jZ1+/qMAFiaJ+WOBd5YrNqkahI+T
8zVVC4qiCNBcoomhjfyhJvePh/q0xRbZbFb6ok+5sX6SAOJpVOU7tNOiX4iJFHHR4qLP01Nad5/h
etcshEWF5zFNCh14fzrw+qCesl5E3EHA5WYd+I1KaIBk2OqXAetGT0KUFvRjaMHUFSNKtaS3HkNl
C1PwwBBZTw5gRipDopupVRTSILSutFt06GdcMEAEMV4JBOzrYRsq3fbgd7L9s7QjyTdOFUlfpeRP
SyxSHIXbO85Rb8MScbi6NEc96qiNe1KKRmBv7aySJzlbAxODDvslE0FQ5hP3dZp6cgmRcqKTkXkh
OGpzBAOg+s5LbOL2TMMrs3r4hNy8o2N1NcQ+FCwZn+7QWleXH+lFWeD4sLPV3K/zGR/qWFY8XOVr
jQi1uuqrCIb7Oxqe8ky7I/iGhRJqVtxH/VTtm+Y5eiXNSn/HQori1/nYInkHKJ29esBD9TGoVzK8
ky0XPpph1CPK3Xh68RBHWTze4MRTQ7GcwsUg9SR1lmD1OceiVjoNVunV+iYX4RocN1tsGOvtrI8u
+6FfCsDG+4Q1tK8iXkGvEbNPW1kRGmfl2kkxI6QxVL4LXTm6uVrFMgadI4LrjJBGclvq1fTiKnGD
4Ocas4/BP4amrM5ZgxPSf7Pfevs4djfsd4YbjSbt9WR8Q5XFbJIKJvu2LFTEqSDfplsqXwSQwbZw
XLbUA2ngLKTBsTfk49FdtzyV08RU5zfkqZy94RGmIK2+xH+Z813qrGuFMJ/rJo3Ce5+Q4onaSoJK
FiHVSNISkz4dYbqI/dsvklAgmEk672ymCBTecXvPw7PpoVrKL20sadop3WnVGl7vUVm+nOwkp4Bw
qdsojgqqcQTQLS9zeseq+hLDOU2VGw1Q32QGmtnwspamx1B4QU6AhyA4lGmSI09f1vjkbM8rZjzW
eycQXAJYmJi8AepNDUWTCXsGCCF3id5ViSVCrBxcGjHUKmWs9eTTuKPBwErxBl/UWfljobnB6h09
HZlolRBZNnJzxLonOHkL7XUxQYk4CiSkC8lysyPbJv2rmFGqbMrv26cGkUZbF1FqdwjTjkwrIogh
H4D3g7gN+i86i3zfuHm9wgyT2XPD82lLaEn4XMGloYfX3PFD0hBnsUJ4cJ+fEUruAQwmG+lGCO1H
GwVPP9Po9CPZOmDRDvrb2QHq7ZtuLc22xjrXkV4Fm3q8AADLntdBQ8mWBJDzmHHYmQ0T+Tl6JSej
LOm9Kfd43JwjziVfefhC8eSLNo86/Udd5lRm6mTx8x64vrf4WxNfD22dXDxPBVlWA39qOUFXQ6MK
/Pmcpj8R4eALDvlyFq9chPEWU0iTqSgGjp5/dTB6+mr7r7Q7bRtzNPIb6aKyv8SvNwewRzSa9aeX
zyEpK8GHx3VDl7p5klgImQKkFcToTEg1TzSk9aoApsUrnDEVx2+KrH6eLQ13W63p5Lbhpl6mTU5r
QznxHckmMRBKe3LngFktpPtaAX0KfISYifk3ePdhqdQbfG/wAJrJOco3KVcsMPrGBfKQ0GFSZYzF
pUOz0z4bGXJdcySiDEGafAbu+VN32dp92kQy5r/gEgJhQS59jTUok4PeaywDdBw4x+D9Idh7SIqI
Ry+xbl4iFNY0SLTV/yZInI5My5/ZPJ4+a04edKjLOvldbxMqh4SuXWDcsLJlaU5SmcHMuKKke2ud
0rPBkOv18f3/vW1A+aO9yd+XH1QBnvXFakx+Io5wNF/NqNnvS0uMh8yP6CUFh8KPT2CKFlyFURzn
Y6o5yOF123Ql4ZSZTnaSxWjaIPljAoRiDEZn5bZgMRHb/bp5IIcukxLMgFjqiKsj7A4p7GZylQvz
UfFsd5nOMA1vQtYCjBO+8B84I+YZV8dv7L3uqco9UZ1iaD8leL6yWB6uEiyDMnN0aaltbqGYQBff
g3hImo3CaKSdZyBVIN9yXQFG1EBBbgvrGe3aDkE0UFGn4KaSlmdgE/vEimAU9dLQC6AMNnUMiExz
pYPJPx/ZjxYWXPPBCqHlBcoagXqEGcM4HVuBiRX6eD7U+zlOfEb0Z72ZNcp/kRDOKZl6IR6mLs9G
cnTrpalgWMDEGtzLIH2VYdPMlTrECsbo4v4tKfZc2cG31Z8YUuh2m4UwcnlO3LbtUPltYtY2C3vp
OA3Ut7kGlDjMCR/amioq8dD2u8hZ1cFq8Lg4sYApj+iMIrgwxnY83xnew25xyMpIyFr+62Vvj+aV
o4WfDgrqZiq/WHkEJIlCOjT8QNIDohtDwz66oRqzBPgNLd05Mcls1bNIFgu+IlfCP5HCkk/vxlO8
oWfSsza0SsCtwgtfuiciUA/mwFlKhEMmNFCqvSZ+8LvW6NnSxkaeeqHwI+qu99Zr+x8JATAItQIk
lGnq4dYZprGbVp5qaiFVaRmPVpScdmZckSiBshT1zLFCVqidx61rWeuZ7RLb/tLClXTXmq/BqY0y
iHWUX0pNPUcOv6Aa8NBfcauHeT1JhVkUo0eDiPUlcD6TYvHVruNaHFY1nCxHF0ipBJqgsILK0CW+
2ZcRo5qwxpQN1rqKFW8wX76Km+hLsqvHkLkDNfZ9/mfDGCzz4gbgz5N+yXKSZLb/xG4dews9R6b1
sR7QXt0MGSNZfOuWOOiw1KRSp4Qn+D4nqKIUbH+/2LGxaosjLunfH9XeEFwzf9gH5SV4q3zxOlMm
xuTN/U2B8t4/j99S8OpC06snbkwcOEj8J6MTGkcsX819gWXJ3W3pITCL5LaC8cvgTHM7nbZ1vY7E
JJuVUWSKc7y6PN0P1thMl8EVMHcrEaHEjc0CQ7dkXISWrsz1Q8NpHnVTqirhAngAI04dG5Q3h/hK
ium8q2Quvk11otoFff58UbRK9n6vQr8TqETsB2tWZ5pIWuWBSQ3hCYyk337NPjYkpRrxM7wFBiiL
+yJb3o0zHBUreTGXknkTmndc3JCd+l8Wu3+Eu4XxHXCbTrCTV4KbpfXPEJpaHxRzOsVzQgXuzUWm
ziKeH/76hiI7zYHCzmd2XP8uAc8sN1vHxV6tCZCYLviwrPdysHwxSBpO5mUeSvsRVrSAHuEfH24F
ZlrFsiJ8yWDTOwgcb9mfF939Dk9fm0u7ZRioHHz/xNBj2JXZyWNZExFK5CbUcOMaxBDoW0B7HCDi
eEMeTZ7dJMfpRP7yqOgkqUmnDSSQGfI9LGUo1IY+ik8Ama/Jivf98Db6cd7jILmc+8w2WofwW13d
DhdwHXKmkLwzPTZPyib7Id+DEbhF+tB4Zm6Fu/Wy12MSTIZ8QsKUm2ajK3kpAi7/Y1GW2dCa40vy
zVeCl6DoJhBnMiWOdXuz6JsgWQVQVbEvwwLr3Hy45otqlACezh1gILvTkHyyYLjBgBjd8cX55aDS
aaF612aBZ9wHo7s0VXvYz8g7huFaEM3GVHeGXI9cDTzU6R6/ClS5a62ntNE2eb5xeQmbmFR8f5A7
LtDmsoObqD+MNdoubeMFukwKmnwt91Y0Ejed2tV4V4Fl2Hh5jJ04CuaXFmPx6zLybZSjpG8UuXEg
KBnygx07CeRrTcESoJLLAffvql8siYlFVbttxnRaHZNowxvM9K8lEEXTfnKctKmi0tn94QtrEd8Q
aKlBvBxWqFEp565B/1hyUDhh6i0AVes2Dl8EA3FQbPSCYmfLmt1kJQn7tzhYkIahmY3LlP+kG4zX
AZGzeSIgsf1MKP5GoMCZQ8SWUgLAQJmN+HC2Odw48Zh5Dk5pFb+BIz+pW4V9E5DYaF5daUtNWAOA
ZmcK/G4ghht+j3+iwWlZvWxtubqFoJU2HHc0yrQHDN0BIK6TMV6i3DXhzR6j3u1yBlMTdwzF7rIB
G5cBK9Oc7aAUuWZlACCjGIZ0FL5j0bYZTQSX1q5lxjHIbDUQerw+kUmktMhsch9CPE6DgbMAsT3X
suEVkcliXBzr41Gl6BfU1qEXhZ9cxMcT2x8yk8kWu78jrzezfgXcszv2PVoCzw5Aq29FIrENB3uf
SypIe0de+dMSjsxaG20sN6Jmxu+X3Mam1OyW3U/vm7VyMQhANkk1qDAPyZOpWgrW0l7N1C4JXRQW
poF3OSjjEAEPGilbOWtEdH8KeM/KYwPnYgwWPwy226+Ut4Y2wlnE2RbJeWJdcWj46WI/bc4MhpuO
cN6dYe0gAIbvqLn/fEvqCAqiAiyFAs++A0v0BlEeWbaoF6dWqKSdDOv50ffnSXawYtU2gti3vO8u
EiXFSWpaJe+mkNTtUtYddUs8v9ro2CnsYCQD9c9siZf2+DWdV9M2EAd8Qs75zOcNJwwF+sFV+qL9
u9kR7tPlKgDRfxUcjS63kQtochZ4bq9YSjTilhnaKrWBhlsFqPYArpc2DTf8vHGEauV7ImGwaTJY
gLJXi5gX7pd1YFK3sogwXwT5tWSo7i8mcpZ/08r34nOf6KB+PfU680CLWPsOXCz4X8em21ckrhyX
QdJqSbTNDrrBRyGdSLJUZfUg7V4CUlmQwJOHQZhu3LpqzI+jhgRaDmgO6H4ZYbMYn79eP9LBGDHy
mtR1euKgkq8EVqN+yM+s6PcdmHPFUoNcppZhsAXj3YMaSmBwNVL5W5Z5ajwEoqFA5QBoH1ypNl4N
a6eONjZM4QzXE+YKQB4Q9a2IPIZMS7cCfN4JLljvIYfyk38LI1yuveVphsC5fnT7etzdwVAkBss2
asea1/3OZ5hhzhnQUu9/f1ZHqQfWvkkzEGgvqqk7PPhhOKDggooraKSPYeCNUfZhWKweTeLyQBZb
PvBKFRe9oePo4n/73Jv8MQFUihDJ3v/M+BGhxqHWzjSF1uyRYk5uaExQFxs87o5AUeXd2we9XcLo
WzUMLOy6LbYSN+SWLk96v1kUcieM0SFHa9ASW0luxaJoooQZMpVBWo62y2zKumVjT7TVfW1+ZQXC
YGkrLcISGn2hUmKf1cZ3ENmLxepxzORQxeiJAl6WnBcyANwj27eq6Uu12mVXUG9z3PTkC+2Vggau
gJSb6zcK7DDgA9awW9SiV39nYwZQiaJ4X7xBgQZ99klH/r+l7YYJYPoeD9Cy1FDD7fajO1aKO0gV
gGr5NmxX3BDalAupxEE1mcMt667zHeqkKA0CtwVRDwZwsnOd52dIU+sJymkp4/5Y9wrNJ56tCwHU
eiNUd0r/pQvwKcxJnGZZTXqLO28/PEg7akAlE9pWBo3VEr8/hf7jDukq3WtEQY1RJ9uDL8VweuRr
ItKc8XpNNkk0iD0Zhw8Oibb7LY1pfe4xbm0m0ooXxMu14BKyOQryli8PbTWt7h08e9XWB8nw4zcO
nYypMi01koKYw4ar6VtvXOytN5eE6q9LGTDBhPQYMrHlMc1akCp+JbI9SCkjDTgCdx2uS2Y1Ecrn
KiPg6KnSTzTPEcN7qGiwRlE/Ms29ozBqQJAUyzJpPIh4AL8L5+pEQyKTfpQ7uvsj9Zz1QJu6izPy
gcSd+NNZTfQjVz/s8hyVaye+OUo7Hum4+Y+umyDy4XE2goRmUJUQ7vpy4XFVhwQMQ5RfPwWPG+0h
oLKQEN+AJxH7BoeWBl+q2NCx+NWsal6XfovJh7Cf/qzbnI6mlYrrqLgfz0aRzPvFNN8Yx070I1Se
Tl3Y0HGhGfH3DJRo2pBAMkY+VjlFcXnOfo681uQo193NysgUpdiwBs+NEiYsOMJ/aSaQmwR6vpcF
7Ql5BUc7IBsBt4EObWz6rlGE8VDKmyZLTEcRrStTSMKDZdCnnCQcq1m3iuDTeW3Rt0dHKl4Rc8dE
SffOAP7xSM0Spw1GoW44o5vzQzMP32JrNePJpSzvGRDjObmediMGMWqjA2wV38dzPlp6aTa0Eu7n
Isdoo88VRpoIa632LnPnd3ewhTyUBZNdUlDQB2+154+Apg8gH/ZXyT1Ds05+JOvi9Xj7WkMErUfx
3cDs+JpbbYteAJ4yM7bzR4imQQvK7+xTdturK2hQ+Rd0AYewOnjziIN1cBfSQ0FGdMJvfcCsu8Z5
G3WouGq7GFTKrlkSlV6Zx++raAucwK7Dai6wiJC/GgZ3PbwlkBpV6bla5aCiyuFk+yA2a0b4EIZd
7J9zJVXBvSsjkXN1jmvpgq31BVl0aapdzXyQCI8XQEdOLzKodVkt8XaCiWWsPUKEWnifRh58GNY5
AIVVfn7QQFiyNV7VKQ2U9UdNN6gsESvW6vADFNYLZMJfT7XSmIULIwQzchdU5H94m447ZZ9dXOhA
+QGpsavH0CueqLkntL6VO9zgqQiGrijDe6OtU3a5HH+/t5l+KoGA3zzGjk/HPL9Fz9OMmYzBx7Vz
Oty61f4cnvowHb37Ai0GBWPGcne1D4iVykE0/Z0M34Unl8vvHRbUBBG/4jJx637rrY7bCEhc089G
5J2s7exGAaqvXNYVVpi6ykrJv2Ii4tM3eLVbLfBrm9ODdIDgyjDGkcOZVfMaPA2hRd1C1RbfqcLg
3tMdoMbPj6kt/FGXwaGfeDgIQCAwV5wVgesZa2xyjVIBHdHG0Y22TmZ0MusjeJs85k62xcF7V8Bi
iBap52h2WMyyYcYxZzXNWjCkERj9pMSsj2HkXcdy6P1g2pYCrjl30zeyAjdkWQ9Lhw4HZ8YjRUYH
bp83EXuisWPz1L7mscHhc/u3UYfBZqLknzgOztv5eqzC7iA6DVYFQJ5xAApVHq1E+ShQOYGxJO41
lwzyJmLFBDHZEhn42viondxgJt2H0QSYw+VDJwKqZ3uGLYMvJ1Ya5KENhbMOO72P/ED6O4qt+78m
ybbOLDHszdtBTuFoCD+wW6hoF9U9imDNdDidlCQkef4XrHd8DeBot2nnRILpt7cnESTP+lbnVQNG
bW+f52QpaofsleAPV/aqa4F42PeAeFgZWiYhTap1N6rxyzYiP+TcLoE5mm/L71gJ/uDWBaVvw5/h
YelsT/MD75JNSGAVQb087ePx2UXIyWclJcCtNca/3N5cUN2JSS7UBVGnwMVbpqJ1MLj9/NPSy7K7
9XwLCHLh3ynqEdArMqhGSYs07ctZwvi2L3IAqLB5G01MKOVwVM6yC7uAgJqm7kGZoIwmvqjIgpq/
6rVzKSCySVe9r8Au1a5FOQYCLXKeGSgdsVCRfd5VXvTD0wBjiK9AGff8VL/9gmm0Ql2JWJU90gbx
WpUu6Ii3mZGKPxrongpnibYLnVJhj1jPkbh0DP2vQJKcc9WuCq9s88XeXr5+npgseNmM29SYG+CC
z7kN0+ZOsiFMB8WFQVl6ljmqk/+OxKY9/IJfZksDSmgoY4jwxHP0xOV/TWNSN4ExPW7mvez8fgRh
XYPRqYPb+2gXF4AntPB/RCXaD4wo6sXwgp2pi7FOMVQhQpbXwdnMY0xe7OsTRZ4mYty/5JA53T96
HXG0QJoRxH5708kBSeMULILoKisAJHyC11B0qbejwP3rY/6urab5iaDW4SxxUs51d+iYbNVxFOXR
kPGSgxoSk5UmQSXE1AURBncEqck+R2L3nR8GqQ0akmlDZ+1IpeJrw3hDr3n8D4Ee4NwjgeiktQk+
hSFik6dK9Tyux2d8uk2+4tvPmjDqk6fJSrVWxR8ImFixmgCTumZBCxWy1kybOrHwR0D7f+hc0DuC
xwocmeUBW8WY+p/WCAjkuHUW73JZAwzcxdQJ8K5+R2GwoIhO8BupcUGIKjLQ1QNbW7/gbpL6txHc
guQRB+DZtLYYy7P2O0wICE0S3bQWCUisZjtPydxxnZZGEPUVrUy6p7w9+w2lIPr6Z2MPZRsmYJpo
WdeZvD1Id9ogoWSHrpiqswhBKcE5sSlJKWM1ey0/hjArF7z4G63tMGvJyjPeX5oaN0Apz1attZrp
nu9NVRgD+9fqrF+F88mMfxV3Dbq6KIIWTqHm33P41/qAFH/XC3AtK7CKps+Lad7wcXuCoF1hY86u
ZMcqfprLaFEHOVnHQ+Wx+bVMNKfRhjFgj4L6LSluB5XHMyZcKX3Hj3peoNKX8kDlLNryU846xgDJ
kxkss1hR6QxE6GURGZJl4gKpUM1SJw+wccPJz//gKeyX+NZroABDGwZv27iwetTRxYgYANfqKWxh
XoPHAoN+XOx/4BP/Q3HnX4YB7KzoqHT+MqPDuYQWRbeQ4gZCQvodTtnawHvliFmnyMsBpitGeSQY
Cxw9yQIrx5Zd5ymDRnOTc4ECRg4pSRpQWM66UgC+gbZBQTFM1BflRIcFv9BESxMbMYE8E9f8F/dk
5Umpp5sei4FdmGNL7GNccwfwcbFDI3TrsH9WFLFzunzrVlNW+jBsYYaj8rJiASmX4hGtjxxFnM55
lxeQgYBXo7Mr196+Yrf615NJ1Fk8rYyeM/yMEwNqH1ZM96hRyjU5LkUMyg5wJ4xep+DJ5ZLuSlms
vKA4NUlcj+fBrEa+1Ond3+iaVrRRsRFBMA+XDPPjKUWmV0dy4Y+jV9hwUk0d4d6bKHN0nhrP3J11
p+bOYtx3qlIiZReiIRJD7cJ94nfPu8kmxnY/Zbb6ensxmVj2mJkB0o1tdg4MCIbP+wKR/umuBWcl
Ix45tGr7i7aj0LGsExDpsCcJbWrV9dD09GuT0Zbr5DAuTMqGSkqUf1GxWqnkyXshcSll/bzL1hFF
BbRLbBr6tHGc0GYaCvG3nU1b2iU/srRhnNcXLwrkJvc1gmNLpYTHB0WJOdpqXS2iXkaLu9CWqavT
vlSg0zeb7OnexaKkL9ULqCAHYXb6HwYi8y+i0VySwLI8mfjDlMVobMYSDIJyTojp6Yo9qXLzap5t
lTCTy0APC+PkiBiRW4onGN2PAjLpLNvdTBd5psw7JAwnzu+uqMxUcOCR0taoyifFSqWyKBTBCckH
IxzZQSyVX1FIf+qFYaJPcu4sau6W01jmdAk5NdpGpx/oKnNZSGarVZfIzKOckiVTUR3vatm3bt0w
ogGo3D+NsHroD1cPt9G1woIIvMGYo+FYMay+a29VzvSmP0MJhCKz/cwky0D+CpCB6w0Em8js6wHE
1g/ovdQ8lOgiHrzzw0dDLQuqckAvPst2gbt1DcB2bUrIhKiMg3Z1o5L473sBWeg/CZyCPOBhj+P1
gLNEdJaXttNQADVIW8TowZ9Oz+qBqe4V0AqQgBij1gZnRuEgpqbyZBzm+aIMoTMczmnDLsClITDv
jh9zLwsumrxaB6RO8scQ6UfcQ5csB3EIedlqhLwkENBIxi2FoLil/YvIVVlfX3oGUmCUlYY4849M
IVb8lgMSHgtHF+DZZjjOA8M3/gaLEvu7arNevMkJrSjQmawslcaQBFiTS3Ap4+Px7hndgmp3TMwJ
8D65GAiFVIzlWI7mWqVyUi6/x+zU3VwoI0O3/8godd5K3uXJcWBroUxyWUqmm817nQCHbnzuy4q6
cqhwus8H4vy27qQhQ2NwjCGd7jcvBtadjCT5oZ1zT4QqzrQicqKgSqEaJGhUpWmqMk0WofI9+urR
HyjKK30I4PB59lWgJ1DzDnPkquEd2nwCN5rm634T5nnDttyhN4yMNtQvaDjKM7HR6IGYYli5JBKL
Sz0nZjLn2QJSyK6SxG+yHcdIv0kQLyyFT1ayL2nfbz7Kvydi76QmC/rZdZ1/Zcp4RJdX4ETgo0co
fBbELCfJfljsE6dRbqiRlOLG5Q3lrxu+szl2YSsGecm/oXOqzdRzcrnK3kLnW6bFqJikzc+khpnZ
pxKdT6CPyjvSMKKA4IaSO4O0JsY8+Fd668/+gSCZq0l4QdSZ2ZMADxcNjnhWrQNLGk0uEP9ylikN
hpPLe02+RxSfHs9DlRXBBbvj6mKqv/J0ePYiwjjYqavrxfFCnEPKEfKK5noRXphobM4aqLm8B0wI
sqoPNvHyy8+ar/D/uraeaa+9VA3fbe3ngCW5U7dtmEvKOQGfdTf1b8CRKWP62oIjPrFyNmZZQint
DKUzyHRYqjaX+qzxJlhgiV48ej3ed0B3fWOQMn03b4iApmRPP8ex/4US6fy/31u7vOzK2FRZ2vyX
/nodpOwaVY1w1gKnWaBmTK+U6z+mtfpftXX7e4GRL8hYRaYp1yQ3NCYv/LaEuUbDaKKlCLsHfxb6
7ZDwl/cn/M6vm8oX/SPLxyDL4aL17Mhu1mtzSGiQiJ6tIYBJVKP+X4iempfoc27IYzd5I96W2smJ
yORDqO7SeGck3+Y5zs5CIV1S9rh6KSJKWiSi4RrlnrmBMtIPkpSLQditRMk1s+fuqUmQaBL8DCPl
zpxfM/MG9RyoUfHOS1xz3KT7D3DPKgJ8bD45c7wTO1ee5daN0aoGa1+9hTr6NnxpOmSF8W7P9SuO
6afvsu0Q1uyMdvRQfosA9zOgRdgL88Ze71SfS9zuEgbhiYiPi8+dN8Dn5JMd4ZIR5iYwAAadwDXR
Jrk0fwZND07mwhMHDzHZTokg47kH4XRJmv4TqdSBpPSY5LCfPthCMGLPhW82uKsFgoPCAJw/wjJD
oif1V3HnbhAGc+vdiCWq1lbbjXzRBOPyTMtAxoY6MZamDA5z0f+NqwGGEbgoSOHCOD1F0ginEUB0
bBZSz7hl3XGXVp+50em5nolT32fxwPi9ClPTHceOfWLKIbSf6HxU5OPmZTAOn4scnOp0nva/0ZLB
VcPrrZyqSUTjTG/iLw52yODLXThsV7Pmdrk/o+8S4YAs6ZF1l+xnpyK0lybeMQK5DMz9uDkU7u7a
GeRrVj6y/Qrmrp0JA+pXvzRKu26kXjicPZnWFRSXyVvpuAt83YxTge9qNhNW7g4icdyM1JSopS7Q
6ukPWVUu9sEpgvLbpHu0ZSxOJZydF/4ilBn/JrxJp8BVHV17ZMo4Fj2Nv/UT0lfaKtf+XMvYsRYP
pmVmy9JwIAIAK2ocb5O1ZbYma43fKvDekz2X1hkrXzlkXAarw8bOwPmlQvrJQ03yy2fsZxKSMNrj
boPpvXv2+40IFC3culysNeLnpaT3UWvfsQOjM+SEezYoPDsHbHx4JIcCQbsu60GOv1LZGCuJbKaN
OICgJZdt0HMSACTnD0NcdHJu73Y+TgdRZKxvfZBnT19NJFbWXFrVPWu7t8kowvWjXD9MarutkjF+
dzywtJrFlzHnbthtvdjhy1rsbxRUYyOuTtWA4NNYQld8uqB/82cFVugzLrkIGPf9Nhm3o868OFhJ
ht5xU62KDWKvkmW0O0VywhHjCrhPp4Q4865l73x+En11FShIL/1G4HEQx4TPj6IkzZfB4/S+N07j
PhNWQu4ivIJrockZS8F1lyPGMEYz/ANpcxaQojgI/byTJ575uhlmNhwMerc+drXiCGoYR6CRY4PN
8a6GMNvFMTlxHRi4s64IAYyqu5dDMduykgw7FTaDnkKWVwIDRAOlBU4iwGNF6T+pZXRw9ezW+V91
8D1Wop+viwqlflswMrNlmO/W7RijMjua/mlJiL28Tp2a9f4FczLBr1fGU/yWOmzwJfZUFsQwZ/cZ
dJoMbODjHtnk0gOrk8sHagWJ86zNlerWRIoWHOs/0YY2pPKSqkprT/YRYx1zGiUL7o36S1ZlOj+b
QXXGqHpOfHeAVlP2sWkdHEdCoLW/QQ4bHDIM4b3fl9sJTaDjHy2CPNYHIUfvcp9oEK3+BYssnXPX
p+VHHChJ2ZxYzVJ60YJ3SgTtHH2NKCDKnW/C0olETJKULZpx4rBa6EtmItvbPyKc0V4/zlTF74Dj
qb5MgSaVK+NHpIs4OcSfl1M2EL3QvnMkmydLngdzWxavkxVb5HbEaDMfA6EOV97ElAprP4e5JrGP
0atGg+oZkfkBPJG3m4BbHXAj4Up7d8HZOesdG+dAcgYR0PV4yRAstH4LgBRxL9WP9dm3TXq2dvJp
5Lc6ZTEKC8puv7z1UmxaYbykOmbbxUpfguJyKx9rkzOvXucN7UmUs6Z1r9cT4AxgIit00BWRqQYI
1vbV9+pFlQexkSzBLKcncym0nVc4K1KPYXCDAQxI5RqaUTCTpvTuAAqvgfN5nMUJtN/1lXsLEcFW
LLEIvkXRWRqkqADCQLRg2cFRCV8j+0ZjD7yGiCRTx/1qPTXCrMTjwOIhJXz6mbRD4XKW8B569IAT
DMfL6J5l76cWRDGOTVxiIIeIA+9D+G7rWnLSRwN8R5RpZeoWUrWoTC01Rq2cdFwCCTvoMW4KYRpe
92C+ATWzUMDrwHaJHovn2C3IrJ80xHSKpxA6pcqmmJxayrsW2VrVMQP8ZwJ2sa+ktgwaLQ/i/UfS
CBcBmQCrueu/tz0gRA7Uau8jA1LC61g4c4eE2bYmfrrKP+QXe0k48g0/tm7SxXDuKquvXUwtcaRb
1X3ru58nPjuW0NQoFKlloejL1tntlh9/7lxty6E248bRjr5ESrRhLvkYfLZt0DUtDrBPzDg2/2hF
xZhc///SEbJAOwwBBK44gkx0T6fvVHVe0psA91ODBBjqrmY9yxkEn1rucVOHfzFXMwSLi9nDW3Ni
IK2P9hMbJuTbcVXIj80kymG5P0NmGiI9ZILpWDKmRt+RXy56ww59y00pP3ChoxRgTJ45Tua6m0jV
5RwVtknqrEHCjTayWl36XfJLqd2uYgXxLJq/IU3NZBtyA6xxT7vZGtbCJdHnQfcq2AjJAgp29Uh8
z2I1hsa0lnJjr/nrGB/39uamo0Z0l+MIkDGtfCZat6VNBj61NzntoCbF1wjANjqRyvLaFuAHRS+A
YXkNByaAYVvBj1Zj2CvO5aRgC4TLDptcqFKaivt5GNxGgtetqmd+MowbybUefy1k0e+hGm2vcUh/
aXuD3dtsl37YHps5YLE/ZO+ldNSq/HsLVc6lGPC4UT7FlxjMSgozNFeP/jcFDCgPy/2vEcxdHX8Y
/V4eOtGxo46WKt+/87MyIraEbT62cJ4SvsCW76M6KFFokciezhWVQEI2oJX9jcrQ8MF2zkK2MecK
m5BWaANI8xUWgrgCbCjUAvB06lMvlNhueVfnEhzAB5kX9TQ6UrGDGkYVSW2ZIKnqnrIB4cmIjUpa
oPqtZdnieYqQxikt2vk1lCMYsSIhFbYhwUrHBr4R+DmPvoCi8dg2acoevDyAxn5SzbNPF7vx7oA4
L9xXEpeUCBvymyVzdQ+g97d2EqcaFfvQo/5+v/3v9w03tdbg+txBEJ12cqI+JftJtVcuf4fYy4lY
7z0/hFdEcklmfSx3OLJImf0dElZMBkp7x3lF9YFJ2BpgoLoSVtnFLk7kZIc5nl0juZyX3+DHAeF9
zpz49NBB+HhftYF6Ca513PKX2Jg56QiDyzK/fuwzEeUaiiFpDimif4h4WhQ4+J8ag0riZ3QuHTbH
hqKXNT7MafMXButoG+zj4FnBWYBngg1tmJLoyxkQ3Ko9GrmDfxBxyScT5WaBryf/rL2sbJRjdW4o
RXNJtQ6QokeMdkCxWTR9HwVtOeOm0yJkUhMnkICORwiGVyqTQsxET/P2+vN/uxeFpNTjTsmlVm6k
qDhpcR758nClQo9Ki+iuulQVxT8L7w8KBhc2YB21TwfpEnJTqma2Btvj4XdNAx+Li0J8w24jY6qR
gbki1hYwQfMfq+bkBUQ/bmYUPXk7koZNvSxpI7caJy6ZJIleDQO7UkrEdg1Je8fhlIvjdEf60lEt
WFHi4ePsA8jd0dIouTQsEXqw7DEIxZV5aGb+luCxMZLJjUXdXy1AeYHvEf9JWgEciPL+8sNcwz0y
wh5DKIgzJL2+VcA1YNhG1Lglsm43MTK9dgIXnoHAoleJ1crPtHzhTOYJh6m2PXC5/MyJtGwuISwK
4WWYqofC6SGv5O9KravD7jvDQ85bYUWbruBr25GvqR8W9XHx4yoEamVkvNmRd55Fyu70kHZrVoLe
KvvgL8vW4rnNv4gqLtENMEhB6R84tQXUyCHMH9sJpSGMdh3Fkrt1G63iRBVbBYybAWnae6QJRsKL
MArjAHVuArouckTeHF5Xx5ahpWHgjr10LnEWu97TaYbpJqdWK11zAemu9XgIA3mQ2DyZvKbs10tJ
UD0VyQ0ns2ErhK7dgo913MXC7zgjMCvQF9DnHcv4rnzBH/hwFX4vGolnQzPfdS6oq/B6AgwvFWQ0
BEPzdL5i67L7ScbCbEY8QcRKxMPCd9GEKY1mKQVbaTki1zZlDNR3a6upJneOIWifZ1HtQ7iOUryD
gFJfuijhTGylT9WoFsmPZjaxfXz7JUbC8bqXIinBGqZze39K7FBzOb63Wea6O262Q5akVFTT+CHx
idIERUKaMmcdQVrimtxbdJEV3ZNEcoBbH8ovC60F9IIOv2KDf6KSFHQ+eg6CJVb0wO4GvbsOPgIi
F8Ljn6khObCHAU8N9/p3bR/96oLlPuo2mcgT+mnAxkGtbYjBAUZX0ajmzt6xw2z7lnjec5j20eEb
ZIS9nq0eHOs6btY835pGvts+tk6u5DkUwRF19UjALJelYznz+C7sxzyQfk2ZrZ2SpEiwy/NVjzfJ
/wOlJjPDPr2vNlJ2Xb1uAD/+dwznPJAf4UOcexdoyPeJktV+haJlywLqu4tSotXOwIIkkEMp4jVM
OuvNeYYtYZHLgWAy+8i/sxtQJEAfLvGthSMPOtLfUcsG5AVr/9sQU8ea0iuJTpgxkECzFsKEitRW
8nyAdkhCG/7YW6n5DkWdRpwWUuBjdgdhUV1FvrSD18HEcY0bs6i79qWLtMTtsRAPjqBmpze7E8/R
V5nappA37KrELEi4PpkRHa0vTq9q6IRlYmZeBazktMYEmsUl3SNXR9ft1Ylyo6eXHtL+qbNzfz75
eHq7l+pjtlQUSPNHbwFUWimWWNNH9+hQOua3/cICSH8r+tQdxLftjXU/7aQjb06Omhc9hZ54srbJ
/b+hpzLJkGgIGpZhb2yAAYGrD3aELGPfdOyF0JFUWCDbzpg8WwO34MqeBxH8DL1AJ6FW5VkAjqSx
YIvaOSQ8QIF/VuQsbtOq9WZY2S/tDXx1CWYeS2Dt3JjgH8Pb3fTArT9bM2mG44mtPl3YaeSQhJmn
PpeL6AHVRCFN9qFCwsNUoA7AYR42PKHkRXkfyzFmTALkKCNfSxwY1LzuDOAA+8d1cWWEPSma0id/
g/gShnrIyxjfZISQpAwktFNdA0TxVjrTkoCUNiBrqciLoDfUCtyfCe67ebOwMTq2SGe4BphJDUB2
89zx9JIxmrB5vtr2hapaac8DhHrG+JzcZo3DxhGfvObTynYIXNU6XR8WamECAA7LfQOrscJh5ALB
gUtre9Xfk0lE9tMGhR95H3B9cBTb5svLokVryzS3JVXoe7VaYWPKsZbKOZbjnZkCpJlmXGyRUVDg
NpedUn9PYvPDccrbCExhiC20lDPL8rcn5p9RdYw/ftcMfQIoi81QFrvs9WNpRh5mQoIDl0hDVmvO
BCrhzwSlM5Dn4nDaCeNCeYiHTF8uivgC6kSwftIGTiAyzy8yAS//r7PhmEhX7x4XqzSEVikMw1/8
xRFX9QSmKi0N1xCRModGEBDHMhAaCR0lj3JZ6vrn2ec3DyejT3Lp6hTU9XDHsjh3mv1MJ5qvLLQn
RK4Xkiy2Jc+CMta98J2gRVryiB8FfftnIz3r97H26NQF6alnzpXap+ZlelOZdO4Oe6Dp0O4L0tf3
Mrt1OVG0pE/ZzBvB35sfs3TWkm64Uuk/weujPr84aRfzv+ovZcdKI/PJEydmwUENlCWSM90hL8Bo
xX+Vc0xfG3PPAhwK424cLGiIAH/JGuv9bdKJuVoE05zTW9BKqzIPTTrjmXsp373K9g4UuY1TfWrt
pma43CmPi5/vyWh/fiM7gdBphzpY64CBse5lml6q/LIE/PsrkbpH1KITej4hyD9//o6JGOUdI4+l
i1/qND1jfbrKAuZyf+miXweu6FPC95sbo90QZ4GalvEyDGzVqGs32+0wb6w6hw+a1fWnU1ukEPw0
mpFdWkJKxBKvBCh4loBeX7TiIkxWYHaQeUV33y95M+ISo8OXbmPn/l8fG9kiPqUKw0gaxr/RYo1l
fruoOzpYpqEsoqfJu/lWWiMOYZ9jiHDa/xJPGEKi8CCT6uizHqUgxiJ0Fu4+BwgLnEeTHY1rBKkx
vSc+zvgdTdlQHwatyeQllgXXQovdDCG1NIAYIOJYZotkpFCdMk4RFHVArJ5HL8XOiaqplq3kExEy
0ulF1+F5D/6IHHpXCG9BQciVECJPs2KPagqQXlGiP9nEz1s6M1aHOR4NZ3FZO8pBC/Ewa6yC5Dy+
f/wpHTL5Q+ZwjiXs9lk1TG7eEy87xDVP613jw4efy+c6eB2n7o9tadWO+5fU+JgFXinNbeHu200g
Iq5ajQK2GkZxWJXVq+eQlztTMTWQbf7eTT3uUKbYb60uBkgwuwi5W7rfHmMT0tLYYFZaZTLNJCPy
8T8fwFhLKClAl7RsO9RRDF/4QTV6+pEoxAx+bwkqiiCKk6xoFtWQ4ppw9v8lZ7rkhum1wC1C2bcF
TR7c/OVnG+a/OL8gX5r4EzQJM0CuBkcd8Rlzl6a/cNYkZl/0xXk+oyKyHgbOJ3/xeK69el3gYGxt
jgEwxfE99qOauMlloHPHnZecoFJVqoX2TS9nXT34zRD1BvgGtOOWyo+gOdL/P8B6YlRM5sPq/1EK
6MZIlnH53j5fIR99PWrArcEcrfBdA34bnz5lJIt7SVZvhvc/+h4bUOKBPoxsdjCHOLKb/q+R2btT
ZNLNXj7MB5TbKSe7uRV7jzsxUF0PWJQr7IsXX/JKg2dMsKAKIc/WYZUHMtKnZL1CCAGxgR1SLRul
oaBROyZPANWwiNY77cM1w7SbcZfXCbpt1/K889Z6P60zQVPkYKeWXrzj2QNmYXOu+SnW0kJ65yS0
3B0BRwx206Q42w5SnQ06WPkEHRkO594Z6vmCxcVC+pETQeaI5WaHjgtDEzznAtE33zgTwbLl728V
Y6BORJ/3QVSvyNGiLxs2AgXlelFZONB3XXa1BXnW5jwDRjPWo1k/1A9tlXpC12kUSkTv7wZ2tv7c
XMeN+tH4DrbH+W8phrClUvwklfZbqjAZ1aaO/AFwb1uPLp/rx82lRiDcb7FVaEZUEgLKvQyrkY4B
yr5XFKLnycW8QJh8C/zgRQjHYLOcWUkTEsCOpyykCMkDLUJEE2nK7v0N+jhc4jj7aqaMmLgCTMPD
W3PgyC1fSOi83QSReFDtEVuKrdbTbe+8Z5G4yi6xvex6NrrA+qxJDQlPNPQ+xqsSxdQowTcg/hoy
Fq2ZErXpbD9zP792wGHUmArGzS9KarjrRL5DMwV8fNADzWP6yBxvZOVQElFY9h16+MqbTJE2YK/b
QaYb3tCMlBY9sTkY8mgZpatupZfRYBYYWyoD8kLaqSRb2GN4ezkZm3s7A2G+ZooyyZ2AD83VkscC
8ZURGvc3rR+4KiEoArVm9Exhkob9UyQoldpQaHcwaUHc9D5GJmkAVtiKNV+Ntu/NzNMcZxr83QTE
huxb3XkNuA0aox5ceaozVm/g+9kYwTKzXoOlourHjwi4uhrEiGdImYuxWZ15t4svPCO3aXvd55VZ
K0ZoXpaWlTyrvYph0+m1SPlqsJkUpKi4jiEVUN4GyOa/KYbSSLOOkPhQANbUEM1jjObLxQ9w+Uki
/jWofH3SV30AEIWyPVRZLNP5+ItLnNxTG2a0SfDGNf/Hm81RIQftEYHr8bgDqn3LrTJ5jjOJpnEo
+FALf1feSwmkKP3ADudDD7Ky/bB+4ghYMOPTkk5f7yu7km5VHgrzwl2PZ4Kv2rIa5K9Otm1cFOYO
05n4cPTNVlB1HoTr7LtL9UUKLhnJ6f/xDlHSDPXFw4mRAMlAZlrISYmWISZZbgl3vuTCinfRwTa3
owsgvSpbVQ1+NXgKsmDB1hKylIv4MwwI1CvyxP02tqlCURZfx4jbb2bJHGdJG8ZT850BcmOqRQl3
J4utElxXd/7CmgZqRRDwYcCZ/g7nng+1UoAo5+O+qPBxucukifBwHctkmTAh1f999ED/MNw9ckwD
1ZHMfgoA5y7MBZ0DDt3Ri0crZq+EVSbonXCr6PGtaHHuWKZRvnIphs2EsJdGViQCTxXEr366QMOS
cz8wkEMKFiDJTw+POreutMcDD+iNB6E44idI956Bs4S5MoRvsbzeju1NmG3o0dxsSBBW88dXOKOI
i/U8oSxzx/xK33wQ8LdDfMG/5qxo/JODIp2jbs9VvsKbH7VzVi+7Uqi+HKiS0MB3f7qM6ZTuyXCl
PCgsTEpoFuxNKrnleRX6S2QJTXbIIOtb7re8Xhdsm5Z1FxiqRnMhU78Kt4kzzpJwC6IYmOZzWWqV
FFhRicmytzqA2alNTt6xbnklxOxV8cPMVCdibbhpHI6TGufhzp2aWmY2OEbRUelYdni9qaMbnM3m
YTJUabUEwMFCZm1g2Iimwc/gITinYU7Xk1/fCNUj0UZwXnDwQlu+TrQjoKoEXN/Ro8XBmduHj1aA
DMEJdsAltuNf88A1qyIfOQsK9r6MDDV5FKJXM2qFZoRcSZhFMGO7xroQSiVVgG9HB99BD0ODjMJO
h108aqvhie61SAbkIc2Y9DbzVeL89ThFe7/g7grsfOn1VTYzvAGP0richTG2K3li32LQXEFlcx0r
JLnmc+5ZmMMCmTpNQGcft3Cs6fLEVQiz0dPTGavXk+nsAx0QYbkEHn0t47xAuzfUdqfI/5GHIaek
lujZ9TOWdJU6pzKGtGFb2JOk37RF3tNLV4nnfWKumkfSC3sOJgXGwmZ8lWl167u+AJccv8EIj336
T0TNAmvKgvmUYt1moK0kSN+HpKTNBLSqFDWUZeZNy7z1T5bunUfeGhxeh9JJsnZLoz718NJWtb0T
idRe644WTVmXZldVOLZL20agsWqx0iy01dyLyXucgyXiXsERIX5dGskaaYnIfTHP5UgBFOqLmkLA
jlyWiWvi4IZej4TH4MAJL5+SXHRgwNDle5yZQh7YPGEtVhJM6AtYR4HyGvoB6UzCtZQV1Ie1olEL
9mdDyVNrBIuaw9L9rACUFhfs+LEvEA93sWAhmfCJyLK9FcbiULUHZJgKguUKNCqKVM1SsgGoyLpB
4sOWZLGDHCEbzVSe80kpNbOUDzDdi9/PbYqqvs0TPZmzsg61wgHqOl9J/RqasEhkiDKb8XZp2c0Q
RHJvmlsQ8TO6S5yMFKcb94iLezGLYJUOys4O0hMj62EgFBut5ZarjoHj14Oc8JLP/Hj/H6kmWCws
28aGoziAe0L6YqY3+GGaEGZVZ/dOobZhETAv/9UFbkvImeRpriZT17hBVTn5my6GlcmAZDbTfHFS
pV3wfbNhpeKWDTKXOI0ct2spZgta+sf1wxPhM6Y+cxVEQQ4/1MbFEb2rfJ6H1nsSfEM6Amh70GV7
OHo4wEHSpSbxMQnhTnDpitzyKTHjNsveRb5UwIsQsmq+QBh1/dhjhs/tl3mAsumqtqvCnBhroDRL
hD1jjH1RQJd6PTnoXXibUR/syLIXEhKRPe/9f8lqt4N7zPpFHWCZYeHweFIUG58viX7JD2xd3b6z
al7u3ifZAlcScLd3/gL36Jwk8VYarXMA4Xyem0dt+wwTJLHJUhOCXaeszWMW01BjQw03YHxgpppo
9DGjx+H6myRpFVLoz3W0lW6XS2ZlGBZfMyjMnp/CWv8SI3dL41oIr1yIflyuFeAWLtXmMX4hjjDY
1kOiUjeYB7wT6NT/PDCZDegglp6Fbmvke5vdCxhCKkSO33JksmVZOrSEwC2qU/QlVfDEn021dhN2
SoUENFSWCF36h1sxORsc4iZVINyrM/Elimn3evLWYp6HUuIOfHtuhw+VjmhvU/9sliP+lJzc1Txg
tkWDxgF2gTRrkw5c+KlGx/mW6/SHaXYRRRM2kb6Iz9729/VqxIOZzXYhq/llMI83RQt5IVkYfYiH
T76WtcfXEhY6UCmW63WO+zGKXzhQIZGIZSvXN/Rp75Deox0El+wW+bwn6CJKhlSTI7dUNxX3Knk1
YcV5SvZwckwPdv54sPbN9UfLk4J45iDHFj6Za3E1bmb3UqHduxKslN6kGowA6b/c5KQ7JHQRoZ+Z
/b3ubW302AZurBpTFJH8WvcAfDUuZvJ/grWrEq0wnGXIb4B32RUVnA5f3kPGRa2DzlVgCbMfu9kf
L6FojDoghbEC9ZB/2WJKMNOgJmr2qEHVgFh8d7VzwKeSLBeB4g32feoGWjuBsWbAUqU7Sp2sgyrW
ezC0FCKpb3GvqdoI9IUrbvE1JldBTFV8p6NXdHeVzL43+W+eRaEiBWPDROukSME6XbKEUjiD6a8Z
ZcGKWO/MLr+UdLw/nfAQqPrULlWgyeq4gvyhGF3pm+mdORgUebXF03TaSzLgS3J3ZH5zXJTseabG
RbdLEULdGvqwhN9efBqo/LtOudunHyqM2Q/G4Pz4XMePDQmoXO2g99PMn7kSS/B2x6Lb0PGPyuUj
xe7vd6s54rk6QDB5SN6qLZeFA7OGtFZUr61oOkI0WceM0n7C9oLwFmRKfwUAzsPjcva0jlcc3Mj6
oVRFE/jRJXjcnkZe2ZD+e2L8Ax5GWmvPAsMLtrEnXeeP3pe02YsS8GrxvXRxS/nFq4hInBC+kHky
tzQpSvVOQB5x2wIwryNB26zoufQcHOGvrSafaSxrv1s6HzUU+hxrBMCFlHvsT4i0MZX4oM+4KGdz
TH+bCs/I4Imbt8VMMhQmUPq4FmbdmexBboK/S2pPQC3kWOOTdJI5uqLYie5qv8MdA9dTK2LuPVEr
qLXLm85iXtJsXUAGXTF35qL5rUuIAfEIKIW9WEGHgmH20zYBMNAjESnaOKdL4gewTNgoGO8cGqTL
dCNlj2oElg68w20uqB6qBewhFK5mN2WTXZeJyPWr6mEoyBV/mNYWMeXxGgmoESQBtRiRfcxLaxHI
CMMUbk/QuRg4s1/FVoAa2avpi8ym7y6e9GWIQREgmdxBP9uBVBfeeoC3D7TEfTt2d496uvBFMQES
rGu8WmhucjhpFmNUelqS0GQTgWByzX/PoR8by6qYH3zmew3qIwx8Lzx8HDEiXPoHWD/5zsBWjLMI
QIturd6ifKCJiRPNI1SZgZauPFE9qVMaGNsv1RKxhVV8tlXa9/PtwPTTAAaaoyTq3Ls0K21SGrcL
wRloxGG6dljGSkFM7CR7KcDkFh/KtjMCZphtzXtHhSID2OGCSTXSLTAvrIAzVyGbWIFsSPO4ShTw
uXyaT3yh5ZninlS0BDFPD9bTOTcT4rM2LmFSWK+/X8jwk9o7mAWHKmkKEdocqXEkJ1CqRa6NFm7/
GmbEBOwR9aNUs179doypZ8ojmj1ReaEZTeM7acH5C7eOhC+fLIS6jfiPMs5bb2h8qnzMhF00immi
6M41QBi06iod0/yVTXNnF8jqqgbYzBxN4A30EJywzCinjhRErD3ad+9Pj+I3KR+xN57Ln9c5eSut
S9aJZQMW5K87LRll4SYy0pnjBNLZDKf61WPUvjSEb8LkUJ9J5kewe+T2i4zX8yrt41RUJTD90W3i
8AkaWsXcmhSq8EDKFfXXzuo3OE32DTh50h+WTEBU6rmCTQsKxtbFSLnBBSXgsmwWiSbq2v5MSt+4
Akv//QdWSxkROTakftl/HiAQaZMTxmdq+Y29Xo5R21dtQMDhNLCiRMghBxnkNwNdtCHR9XWw/8iW
ewEfqo2M+xHsKsMqFQdVpYVWQoskkjbF9gdLbLYrwz0kt7bdR2JK3QFn4mIo0xa7ohpbJpNQ6dG9
YsC8VwK9YTirNIdI2jbEGW9ByCdCDwIxGWrWjzhIdQDg+ZgZhUN2a1X4QOjCj6gF42qej0Of0UNO
KA6Vk0ZvV8MbK/3Lad66GkTTissux7oW3G19c2+RXcyaXif9i6Zd9yrWf/aFSPfQ9OF6grfH1edq
DFm8bXrcL+NkoO6GNhlGWWE/kp2tKy66apoE52izrEVqXZhZJn1/6ouOZrnyv54KYgQAxYpGokqw
UDv80bukdBoYKmvbkipEGoHbVAcwhQhyXgNR5EtEt2iqEmoAkAyncXK6GlVmcE6dqPsvJz3Usx9T
gwk4D6prxy08toO9CM4YMQr5DeutYyxdYW72HWwS2i2j6CZAjYOlXXlKyhQ0I74TIYgcgrL1cpZ1
ng6AYNPC1zSmqWXZW4zn1mY51W7kGYpK1IvVKjs/NX1Rf4hqyR1QYklXHuSxDoQd2U9jB/97dWS8
CP1WfZv+F4bCg01UBfstRptRpXH8IsX2k5fOe9IBSrqi5EKFM94bcPld36tBDcrS/rJPT+21q19q
skOIBem8xdLMMdqTH2Ymm+3mEpHyV2PhNZ1j4AOlUy79P+CDHhoYckqdBJibod7/sjbC9k9b7BT/
sXcGXuKB0pa3S+PZIG39TcJXF4LCaJicC/4Me5C3P6BFEzWLbv8lk20e4/zdVd4UKWkZirKwsgqW
Z6Xq8v3hXS8TirNQYfGEudJJ/mNwGHzt78s8Fy7IEWqGdJTQNxTMkFcM+7NcjDyxiN7aRUSUyfc/
H3E5HnhwMvoWJHNfqdARDSwmG8m8aJ5D5cJTBC5KLBszYJbcPWguh00cBW0KEjq03BRnTJfRsPoQ
QzUBBuAWzyMu3GLXXLB4BiDQOVp/y4NoWgJVWsjE11hCflv7JAb9rMo3WANs6lMbEZPvC1EXKbLz
BhI6SLgDHHXUpbc501XoZxrMwDH/nkXqD4O6iZ+BCwC0VXGhvPiB2gprr3o8F2Nnqot9efFRESF8
Nxqn/DzjNmMapIDQ/ohu/LbyDno5tyTva52PiC5bJwd/HYgm+hjmzG6BLnRZ12wQogOEXjoXpgfv
bkMQNUJNYBowbLKQyAfVU+r6Yv3+s2h0t75EX4Si7ey2/Sb9eg+R+ZsPd6ApXKYaVRWbsaokfGxa
LRKs+B6svc8fEkOawNZYZ1/AqBT3BjxHLq2SDEn69NR1S8ql3fxzPU1jiZb+0d6hEYKmFEb0Zxoa
2mBWWCxGm/a3CXzX/mGaeHABXr3FihMN19gxiJDJlNGlShNVkin/s6iiV/Pxaq/+05kFOWbTG5Ym
dXb5QZCrYzVCEY1iCJcARH64RBZRdQ0vG7zTrcRN7EivrcJicuDlQ6q5ExgN7hWcrdQvqcJE/4VI
YwqJxC73kwY6EIF/eiSkSsK1cSclFnLBIryXVTfijLSa8WOPkjUPvMeNu51dvqyvwVYaFfZSvVWH
bKg6Ddv/kRY2uuLj6DrlojcnUT9hGfdtVna38i1b66n5UxXhalZSxbAbtd3x/n6aKKNJ1snGPzNF
JoQLuBgMHon4tPS3T3yHIU9sYypDKUyGOeuGUrxmTeV0LBxpnrnv+WfLXdttS3YDOvJ5lDgq3J1u
gXd4yRhfP3pwGXSk2f0rKvmgL2kY2swagfqOv8B50ctiaB8XWDUYGcMW2M8oN5/qMwtpaTS+v3da
Hck6PdTxrl9btkbSToyBfgkZddqjobS7QQdMibMpH2cnOGUHIJ6rB9xccLa9toAgCoN/3p1JhRXm
ZyPYMea8Q+ew28l2FLg5xUPpGr1tdUzPgwEeAherplBReLDFzFnyBKfIJF/59b9B4qjGpWBM5K4u
AlBlPfrvo3+6J0lDsdz1ZBRAvkMkqInI8oRKRkvuM0Fmj2aFpAwlViCEyqfchCm/wXQkTCFEZ37k
t5xN6iYvrs4okvDKllyqWOL9kNX+EIKDuwX3nLWihOizqE6kEvHqKKAi9+rolr+VpbREX88Bpffw
GHpa1bvHPF64u9MesJaF0JpeNtG5lpT7nqMYQj9OIc2Qc3Gdmb25p4Gw004aXH+/w113GxS19PW7
xk5JQgVDlvz4LFt2dtqgMaPFAT3n9PzHBC188Uml/CrDxj6LzlQa5VkyNe0k8GzOS6+gvwqRG1pd
6Q1hcMVPpVsbPpxC/8itJKS8dA9sR4cx2N5zG+fBjJJOFe5vB8WvZlaKFrEfMuwg9XiZffaTt/sf
iGQD36gV8eRA7NXzkddpttDA0ODdULsW32ucGADG5ip3IrA47NI0dpd4iEiNKrkGzRtuBjE/PMep
PKXvDfmDjnOVajPhF8zcz9IbAEJ1jBv85SGEKkBntujSVktQZui1Zscba0ivoZAUsXPlMX2VX6a8
ca5JPtklE4KLmp3cyXcge93eZrKyWU7qBjwcUPKCsiIsA50UcmT/ogS0qtKEsKEGFnRxkeWtZPwj
w7i/vPU/2AElrQiqrrlIwPckRUrg3PBYGd2ySgnLH5l0nIhjkRD1E2TSD0j2K1tvplXDRkA6UcUQ
5uoe7WRX1uittHbV4q48giDvEQxwA2QBDOllQKOQJHnqf8QixnHZhbx43oUXFzAbMEE6ANyFKqnc
pl7oOor5VGlA1RDRzoGhlvZ+Zy4Ne1ASEQ45UvQ4ZbtxgJYZ7zNQujvRKt+z8frHaLvo10mOGynS
wGO+EXho5y1Nzk2DbUzeUuhNph1+zKAfRgPbfK+3llScf/tS4aOQDTUjKisU9DsQ2EeO2PidIbNj
eMO2p7h9KqL9hTECPGIct4YpXCDiq4X5DzVWnu1HL2wciMA+7poMxyHLn9ihJAXMUp1TbRZKIHyk
1AUEwul2lk32GnpxxtxnnnFngPHEv3vgBqgy4Sa8ST9L3b5vkMhlikda35I/TQvuJ2XuUN2YiRfa
CzwIadzL/X4RggwrGCumFLcLwTuyA2/C4h0ZLX+c710wIpgVmOUwLzFBPA5XDPLgkmYrBb1xX6xW
hrPjkr2OTJCVziTklvLGfIaoRUGPJPLL+pD6JegzuhuQVRz82EpXHWv4FQSs6AGkFiH8GSXlh6OH
SWmgogjqdaZo1dFO+eN1OoI3KxmhbgLaSyqsooGehCx74euVn0dEzCigyHox12uFvGM3L+fCYA5x
0qtGsOKEGsTZEV2S9ByDryDbj8uvNcPFoMmmFr8GlE3mkrxbIr3Q+9kNNDQFwlmDJ9gBwhb0UTav
3OUr6ka/C5AXr+3bBXW6ogFDCryvJ689iInNHo1D4JwJVwBJpqj8ZGbdfpk/rXSaElnX6rBjUt3d
3o41j68rlcmoNNvaFj1xJhaRCjZcftljvL16f0CwKCki9th2jFOHC+oyvDWiDoJY7CjdxY5nefc7
9MnF1s6QFgzZot3pmzwpZl9EzOw0iTw9oWlS1Xm5Mw/3KokazeG2xF3MU6UdFkjGW6OscAgjIxE8
MdpjGzM/aZcx7j6bhNIQC78hEAMCsX5Hzcz/x5xlr0Ou7asXoS9xz2wxiDouvP+OmAS1La9rmcbS
yJApXSQPbW5vpCxPfXsmqpd3uxVWoJ947Una0Jko7HhyGP1NCC7JNHZzD/z6VUyw2zXf3WFRjdVT
CtKVF+jOZoX7zEldQMJ7Oyp57z6bASBHcWzyxsOWzslQ9rgu9QGr1E1bSRoI6Ym3vlh4wZnE76MQ
nzk+KqVDB5Nk7pK/6AYANAEWLoicYtojIZlIlhRGM+6ZY0ir47OrPpoREIkuMv/KePEoovKbyjWe
52BIzJCgcMygfYqvQtB1fsWUvz76kpvsOSpZqR5ak9PxQtQIpFhG7nqCJGqnA962SV2ff4Ya97NK
O4vJ65BDWJIdLUYDCPha4oOacc9v+4VA8z2/zyI4kElWxt68IwW4JwkrHs6N1w0fSgUoxL5dyqjY
ZOtYBcqkeuAB95v7uJm68cccF40qooXUP7aHcy11QJ6qXibtkIgSq5iCBrFlMushM7AV3q4L1nRw
nkX67r2FoBTzsN5R4P6AK0yYzL9OE0lXtnAyiV8kP7uKn4PHsSlTRZmgi8a7B0u0y4RRgF7nmtMZ
hFCoSoqtOpKlJApA9rOpMGdU3y3f6Bh1Fg7csy+ger4hT+D9vb3+3RM5VQM9XxU7KNqy2fCEnQVE
QkVNtby+5YhJNA0Kj5Pwl4FhMViAvlGc65qiO2UyjoLSsx6Mu8qQ01kgoowOh0zXFBlKVbCMQ5LG
BYdc2uacR6ZvD0kOX8OOJr9W+u1PkOgCmlcgtaZs1wsVcH9SHC39PCSUhufk5LDdBeuqdliTqsGD
UNSPYJ1Klt1eJc81z3a9ikCf4enR2EOeXNBoJTWUKiVG3CufcvrOI4KYo+0PFVnGur8Uvhq1Y75u
A5te8lwq5akCDyfQI7SiTgzk7t1Oae9LtooviH8ua+87B4BxF7MTJpF/h8o7z7jeXJY2w6eLpTbi
HcLpZywnWNEJpmmhe5qLQczkXUbIS6uQiJF21lS9f1KTY9jgMKBXoANmVBBsqB87K/NqE3v/rm5o
GFXXTJxLORcDD3vOGHqVDA8zwoLBsSJSH1EabCj2Z7+G3PO8+FHbdYy9wGnx1nLaIb57WI8i4Lcr
l06SupG2g5Ry1HMq/kAG1m6g7OQ34rLih70Cob8WYmjoPF5W/kBit+pLqRqycMhl1v6+KRmBrkyg
PgGSKvJEdUhuG8M1mo0GziZ+6n40ur7vBimE2hXtjHhYCrtW8a7wbvL08jMmQe86jXbAVIAlPA9J
svBd6ATSwDSGHjGoZx+b7Uq7M23RAzKueuFyaVVWOf0QHc4cx5tICb0rbrwSngcQWlWTVbeoTqYC
2QiUj7tdbtQPXfLE0E35TJS5/e7n8U36r0NvChhAA4RO6aJoeNKZFq3vREKCsvQfLhE0gxuD+Jvi
V7aeMKNlgp3SHYueICQnYnar7I4DlIdibYrmDIjIgKNCLoZF+IzWnM1tkM6SrbvdHNPtbtVBhtt7
5FdKa27f3T5dlEh1u6ZHzphxz2ouABEw5CMU6eFnZb3XuRr5yhVU8r4nFvqqa1aQ/FadPBPtIP10
i7Qgh3EXFgQu+eDFAu0qwMS0QQ9vjHVc4sy+DeOagndd7XHkPfbjHKb5O45aQdd9xAM4qbuSv/NW
ZWD14EuzAGa2eTbdbIxV7txwia6GmfUs7KITNxrBC2QT6NN4sLCxHRyLtXvH7nJapzYVoxOiD+Sx
lT1hB1S9fxu7qqtyHHV9ak1kRmeCMKXMHPTstqaBoPabLeKgakNkUEeAUcT/TLlj1JGb1ji4DEgR
QoOEpL2rEpCReA6bZV6yi4frXu3EXlK4JqlJNW4tLleFqe1yD1Mmtt4eAUssUCIPKtHUYlvnYtup
UpSewnfdHjy2EJnZ7PKMYzeaakpvSE74ajsjz0nlfy+X37AvMqDtEzqOY/UzSu+ZO2XT0XHjhb28
oV1dzWnR/DajoOK25nMKpiMAcVcqDpSeVSZPyc9DFKxFiiDlarWqrKYj4foJO3SPhshEZEZUBlRz
G/SW2JAahOF9nR0XVTBB4O+RPItyunZFkCjHHrYeuuUKDqPWWxwirYqudSkdplFn12ej+5op4fUn
Kfu9TZnu9MCoawwRg0bpcpHVZLNYxrhPb8y/80+E31BZEusfRirKnvfzSMQBixe53c+npGJM0Cm9
qCO3g1XDLGfwGCc1k8GxPK2NC8aO3/lOcm4jBG57AR7r5KuDjjddNWwEAMymMG4mp53JLcJMPkOI
edsl3y7BPyc0twbFs6/XyMxzpOwchE7b/fG4oVPKqXL/MVh/qkWqRyAZ6ZcAL+Xm8iDG0svqtNw9
NqBlc5HQ8bS9vkaTOBt6HDA0EDMoEGaIf0f9Q/cAnsOgDLgksR3585KRFyTTzNcOGNghbbRRSQri
lDiMl4FXZSNDwZYdW21LpXe4KMfaCadrmTiTLX/hHZnZVTY09Gbyw+vS530xDd2udF8/Jiv2h7b8
5A4AkWPdyQmkJKlwrK2X/QabqQ+Es3VwCPzYOxJJ9wn25Cu7hAsQbxIBPQ85kJfd1Fk8hghbKHPT
TPc7PvZ0G0vzGM0xxWDpQJE4b79+nugezICN8vdMdXA05nTOEfyG5SwbME9fy918xDd7R73RLhgO
vukzFw5g9FGMvRJuhPF6vBkTiV8GOVPdm6crF6007LbfGprEWd2nGfOXT/aF9O6x62VLmYDFh0QQ
0EK1AitvyDo/B2bNiJmU25WAeoY3Pl4Tk4sR1Zje/W6n4aAo20UmZ/T9wtlEZLtPK1mSggk9D93G
RuBr+Rw7Mx3rw9H5EUEQTMk0D/jF+FivK666WXgqEndCbPRESLi8OKHMsKuRZLyEdyah+k0D9Jx6
of0cfSGgy4pT3V0ZYcDNOSHpiOHmlgpEG3dp+GbCyEvTtobwJuhmAB5Cz5POQEERLO7G7rwR+/Ex
2EoHx7aLsiTuo6rFiKkXVYn4dyzUQWMRJJw6p22B3Bitn+rjLoX6I09vngFYrLnwNQUOSGlak2uS
a+0BIhHkJvIpK5Hh+/bqN8F6bNpSNL+y41X4FQvqpM9dktZqDLmEY9LLVHP++WZzLwtTwAVCR9Lk
BljGDCrGrjI+zZqa13XG0JyVioya+TNEwI3V7qU0LqDfzHJpC/cYk5TviBYSrLRiwiLgGMKEUtgd
QBLeaKxY4qCqC+Zk8YI9SZ2rxfoFgLwR2M1Wn27kPD9nJ2hLzOP0Uj1NQr5h4oHxXN4mJZdi2t39
+HLDDwQBOIaxfB6hu5VCtEnH/zr+3dSOuWXvIfM5tlt6Vg0c0O1lvuEAW9/6diu6XpsHuEUscbSq
hlD6mbXa/JYjlsaWOjFYbZHrkDLkUxAfhzM/+aX19S/nqzY9RpwqqSRp606bMBAoZWAlFwqXztsM
5EywjTo/D66GBpVUtJ7v/lZP87iG2BtYis/21t6/nlgv3Ea9kUFZzM0J1Bkb95IREJp6EV5tI9WE
JDYVZsr+IR4knM9RSKZYeKC8SZwO1eBs0GxVuQIJ1OFAeq23WLdTVnoBxRHA2Cq50GqMw1p2zLEg
krRg/DZ0HwHra6Q+Lx3NXGaE85EusgxLC9WjrKbwilOunrX5wkDWrYp79eLqxVV00xUS15KMbbMK
2lOJh6q+p/LBxBbZ0KGzsOQOMPWiimiwHOuBLTpdHEBWw2GpBYWKN0Mon5vNDCOhFf2RVJ+nvdV0
AYZ7ObkPyd9F/GRYcQ1GLbaI42yN14dYy9mhFD8sV50BCVGx/u7r5WTMQpUMExD01ODQQbgHc07C
0N9oHCCtIMJQ8A/PRjuZftr/nUF/xvYu72pI9JkOvTOAs9rftYe77MQswLarGkWGtpdE5e0paTPR
K5VnPEfy/OlmoEy9PX0YSkWvPohvrILpcIYCKZyBvHzV1UKdSapAl8iaKxcPEX4EsrhT1DW/P394
s1E6XM/Jux2x/VVWfkFkdQHTNzbvJo4u7I1qCFqzhBE+mzd4PTPkWoPxCkKX2YBiC+rOEPMt8+TY
Su5CzzB9evgd2pLq04qFaB2HUhWNHc3S5L+jjT4KXLmBDVFmAmQEmsYMMEgECt8DaQR69nStVJwb
UGzjX6o2kAQxOk8IoFnFb7TfhVb49IVy5mScXDcw92ol32oD0bPJ9OyrmEmjzJW9bshTM0vQCTo0
A7YOs7ZgVbxsXrX3Jq8+tHkFCvIOB263XML1cqHaQkPrNEsOaM/UWYvZlqviZrZjdbJ1hQHJ86yR
rlIcLwmssgGobc30bi3AANoAuVqFHdLqN/piPdDxoEOa0uzGMABTW/7hXovNC279k5kpx7cgNY1M
7qFnXJGlZyVzpG9PiUX/ZKjTG1xHsrTr65d0LJOFt/6EzV1HlqW4lIemaqIbm8i+qbM247ykFpJ7
Su+4EzLCAZztRPIDPPzHz6crSx/vm9djy0/myieQHPDwoUGOymF+8AfBkV3LW5ltxu05NE8Tz8kh
R5CJoF5I7nlnLvNh8zVBRiKD3S1kydbh3BGXFdm0j75Yto9dYFoV1X8s5p4EXVtw6R23RZJlpcF/
b1oOfSQsNhrgqKUTO3YXaXDXgvYwKtKo/EWlUuZVTg7GXLh/FtibZSOveK8f4qHJsQLhPXro/cam
XePDI53xjm0MdBWO3uQXln8Abqv9FW8/IKRlIhIkCkywQ0iHulMDxqQojZXZMuL4IWyb6AwW5M3f
sRycp0ZUkfvy9QQwjWhO2jBWKZJBn7KmlOGlDzKSEHv2dVeT64IiZclNybarYVjIcgMRv6xMLYxn
ENIOBxcgaMz0jRNVUIC13UOSYLqpW5R/1YhMu+LnZmrNtALdCR4ZcvG1+jmibrWUijMYglqo9Qka
4vb/V/feJ+Uefcvoq/7AUEdbCDUocjdCG5BiXseWrJJeF/mI762gxufQ+8+xM/dJNZkQwb4GKZtQ
RLkSu6TBUOTjxyXHOOZsdK58757Ci0SPVMnF3ypt41lvcFtt4+Y7s3CdvhaUsEN3fE6YR0mX79d7
V0x/do2C7Z0v5YdFa3/xhKsE93wI05hni9qMqZ81CHfpifYnMajUR+7iIhjk0/NbKCrpCw6SsH3q
jMiEf04CSzt2xe6HAI3SP1U9rKcHsTgGH+2gWP4Jc5IqZ/SIFkjj+1UxohEfLMtSSYV/gF9uDRzP
aI10Qin4rmretcWGGqlAZDYf3QdShtgH3mWuCXLCioSdIHzPrQzJTQKJtm9HLb3qu/sh9thfJvDQ
1VV/5RRZD6LQko+S0adgp2CNvx0Gbutw1oegHp5IZU7tFMujvMgQGUNI7PpSnO2lamcoKfao1W/i
A98dtCHJrEdL0wc7cCY0zs2H9mt1ctuZCNiNyOHoWnAphVDXFuyLGOb3An/4ZdIb5t2XEsQfbz0p
yMK+4qIq5Wk1okWNwNL5PrYm7csLqlDMLPj6sSaRdWpKvtuN2poALAX8+cSDQdaAgU2EXQhsMXzn
vgeOkzGgZksQTz/MYNiI4RKB3MOsC/VAc4Gk0lRiwvVgrwRwUvXxJ69qqM9SIvvdsxGi36PZR9s0
Dy578BwU/kCWakb3l0ecUau52nRUDIxLDtq20NRhByZYQ3+Q8yNHlXSlF0Mpm2Yo2MjckgI9Rwp0
JtiBz2f39CK3TCvmvCAx5yz4MJ72q0IIaKAijQnXAO4Zj7dy5XSafXzEACfcPIgWfJwGSs880Rim
m3YvtacSKP2ngtnoUfbi6cR66+yd02kfOrVL8MpWIj+PjSvlOclHpzawjUYou78Z2tvydBitKT/a
KoHNsXBwwQhIKpJYYi35rs39qGbEZ6ZtlMKlXo4KJeOAS//haNzEjToYXvlEc882B3NQDVWZ0AOH
Dm5s3S7RZtT0m290aUzDh/AcNiLmweElurOKOPYr4v7laBqL4QKc7xenaicAuDb/RIzfHQvJEa6Z
GgiwraTllP2xVtRQfecmTPOuOQYwpbdd5iP4XOzHDtYEtRVXPUSLbt967hAOC+Nn7J6yfdoyulkU
zUUTUnlyWIA9xNLJUOVlWlmlIjVIvY23/7J/SIwxlx+4AfwnzyX5U6kSPlRZLjqh8CLHtPjRJHmv
pt8DjFqr+wcH0mc1OJ2iGZ8ZcBQjAEtecUst8iZcE9KS4UvUd8KkQSb6bACS/wF37AbOLcgZL417
jNUtN4Y3gxsz60BLG1A3OlFeUWqYyrXYi3bULUQwCl9LHL0pB5a5+HgmbjLmabnH25v3dCjZgnI6
paO3Ox4S5PZ8a9rRuWFDBEnHRyXyIOJqVBvDkzSYnosydlHPILyFji1GAdOBeTBbeMFGVSXk2fWY
hZ8+vRn8+7jpzKZspsMwWQ9c5/573JAcu9nVoszfdOGfhvpjqYDWw/3rIiZzZA2t2jbC1r1QFo9A
tBIUpL34yYDEISTZ680PTFiuBvwZCjJmM2M6uTQ7I81OkeHSQCaADyx1A9CvuAl5h/zkuZ2OtbRb
AZLdS+3AiOw/7YjZ7rDA3ZGT0VL5ggMwEYffEsfFHqzks0at2jyZrjkFq3GPliec6lni/Y6TsvTs
3DxfBi4cF1iiK8UzjmCoL3tPYiW9R0TD+uYK14XJAumQewvKca2Qo59/xR3GrzJLrNpvA51v6aQZ
gwHHaykJitCG4WquunyI3HQKtX7bvbyy0AGapKlguEBMDCc3ERHY0zA3kNBP/rR1b6T415GSZTkm
UM6auuSY4ZD6MWpbCLUylH8uGok3PnT6IivW5jKthXmzdslxdP8vMuzIxBK2rt9T71uz4S87nNXJ
iYIkPFU10wpQ2dMrC89Bwj7RE3l5HrTNfoucXS3H+k3zbaJx9cVzojje2EKq4p/5Gt7+ctXapusS
IcHv1LYXokh5iQ+AN9zn2gNbcE+3gQYIWXRDmHrAdBcPVmvUOyX/p8NIJ1CZKR80M/tJH3qAEcfw
ydiRCSJYPAu4a8AWKU1G+oGm4kclzwpFqMR0cOiZtdvMxoOutB1DaXe1C905U5PXXVxv+PoF2tzg
Lfe80+goYsVUgnWbaAx32i4nCBjJ7ZGSPWNp2oxyL8Fs4ISZJVmrDiZB8kEU3GIqu9BHMDyRW8XE
/80lXz+SY7VupyZv/WWs5fSpnKghMsqzW50vAFt+ebUgAHhkdsu7th2GLdYbBiYOp0rVSazoXdwV
OT5wwY0IAczrbMAf/HlvL0i6n25H9JVfO83V7/HPTGlLPIm5nscr9dyC/GjfKPt/k/mG+M/jIwu5
HjzGrBmSJF5jYN1uKpUI0YsIC4H5pm+1UU4VoEyS3T/Rw7wTUYOeWtnHqKLY8BZEPZ+cgl5yBcqm
A37x1GHZsItgg7Fi/etGz/Nz4XXdqBSEppS/GQIdOE9OzR9N+szDbZwUsgxGFLNQlu18pKFlyROY
LQlQSXM47djX9gFTvdaQi+ZS1p6jYF2Nzm2YcoH3jNnw0jd1mKqhnS5VlTw7frFEhKq0LjUOu8Dn
w9Lg/JvEKWesDr93gpD99uPI79x/n6oed+Avvw7cddhRXditJnrn0cvaksq45fG3+H3jrEt8nbg8
EivF8Vlaj5YwRwyQ6AchrSOrWwDGeupkdH67RT7iM3XpOC9fRj+Z0dEZOKD5BsAzNQlxnH42pMtY
OANcPvE65US0eRLPAvXoXAwhsVsNgMu0SH6/lixlZVMTT8BDEe475J0DfONVRaZkGFWrqK1LNyaP
BYF7r/NxhI29LaXelEIUuzqiM6RMiHwlINL5Vlfpmsuhrrv2axxZpNs+wO0Fu4lSo73u/hlphZpy
yHn7XfKXeNAqi6qdaWYzNWCln+akzu5pQjXu9bYq4MSS3bPtJKTmC6rVa1Kzka1HjlJ8WkdvF4C1
ZwI2iQX/4zrSsmWhXOWRCcRBcg+mx9ANYMw5vKisJ/jjsyREVhsIZ10qOfndg/BQpJU8YawyXefe
y7TtXsec0RW/Z64GRky4+C1k+XgpRZTzaotIPTfQ6W8vehixxAGCgqtNdS5bFhGHLkRF9bza4vY8
LurAKk8+eTM6DCzH+VLXJdUM1+2Y7VWpxJYysPGyO2hNlqEd7P6FROjPYAxmq6dBkRDT1XJLxqn+
ZHW56yX6Bce5pPiMPQIt0bKoo846uA1VEHSOk5dTv2+hJTyGb2HEwA724kNZIglO3tMsajppUyMB
ud0vl7UYZEm7v+xsEUB9PSsO1l+0ea6GHryXR3NEn/ywZ4lH7xBJJH+xKpl9Fo8GdCiIVn3iMud/
3We30FQ2sIncjLG+J76/eQFGyDSzSDdiaCi2USFa/SKR2bSmRvJtqkSI2Bx8JSKHUQx6NvFyy+WS
90nnA1UFRJ1CPf1gvU9MCvqk2Je/p/gAPXz3H0v69AZ6Qce9sxCZvBcFN84bekNLFnhCVRpwuDcJ
9E+dsUIodBWx/UM35AYqk+ri4PHdxwEg2/yuYXb7QezGD+oHd/3pJEeBvM1MOftaGeIbFeJhDZ7c
ydOn0Zji5xAM2CTZewDIKdcywNA3x7FJn5fyao3c7r8oJIQOgB3Xf59kzh5P6eT655MWYp9rI6bj
Rm4LgxhGgxCSjnYV4ghAQ6w2ZJtsn9G0NxwEUEJJG5yznW89IT37qt1q3eehd9s4ixCB0CV7nWPC
dCvmO4dcaqVQywJP+fUP3VmzpHwjr8G6PqsJZ08NZdjaKoYPvFhpnjTd4QUFSXUrG9/9CqKQeKwS
ogXOlRzaJ62D/7rK1TWY4OxN600PIqXrJo7Ln/b8jEPTIicO/DyL226R1hiKdUjh18D+QYRorgIS
DOyEAz39rsttnWaCmASoSBHb7szHivui0Pifejx0TiJlyBb/F6ZUqjzcql7MElQ8NLcADRVftGzy
j9ACFjSuWI8wgdR90VaRCCXENIdR/nAsEVhcN52+Rsxr77OdA/1fbAt5cQb0vIl/VeVjcqwVNSKc
oy5JsB3iBliEw1MW/jNuT8sby0r75dcukNgb32NU635vvfka/IAMxIC3pEv5ZDe36IQ11WcjAMAe
lkXmMdDuRS/+KBhZUUgryVHNsEJsYddGM+FjuYTu/EIBaeEFZ3Jh+abQpeJsEVFBxHmiZQuVA+rO
1sWKeu4di+oAYgbAnt5IUD/TguMY7+HD+D/L6QvaPQexHBxnrXm/fmEGUOYS0uKrSfY/7HqnzPTc
yAaXi4HFmu6ozNjYQWMIVPKKepuPWrU5EtnaPi5Pt2XFMLcYzaBWZAML5jI9pPr/QHytlzvxZarg
TqxVnbENOeT/GRF3hN/p/+I6UjxTQNCaJBqLh042FiXz3CM8A0TcvBCnR7JIXfpGjU787iwBUuom
FjPfNqiiIL9BN0B+ZyYted+bXtdVGQS/AhRsPtJanjviCsHXTtHtiC1SEm4VxF5eifStdftkmAc7
vKIFIhdyr6POkqZ6X9uz/CExNJt6MMq0oKjN65HHAfFQ5B3d17oeQpc1zphOlfUvo1Il5NHB2N83
F/cg4qhWnPeTw6zSIE4fUvUr33Hs4cMXA1ebB6hpIgR/jfydMkK+nwlEqtiU8jhM79Nn1sbNyWCh
QTzs8AngMkHpPlT6OAHR4XFjcqBaZk7PuzupL+AayP6v9SW/K77+riQdYM0Y77d3uHudNtVIKAG9
slgv+VCsuRG9y2L8/3egMubTAwHJWv5qrlrjDWiSmHNvxWU/PZ27I9x9pRfU1Q3Ld+XY8575Y0y6
D1FeCJ2FBM98TmI4eeRE3Q8x5akPvKjMnD5DFBEMStjd0elPXOAFS/1ywvdBphyN3HmumzkbnpkY
aH6GnGYt62djgq+3Jnnx3x/4bh25DK5VFrUD0tB59kyxnhbB/TOV+d0JgFcF64pt9i2dB9JEgWWx
jgJsg66mn4s04gB/fpHz2F+QI8O9YQarzdprAiAlVlLy6PEeKaw9v742z5USJtSuDKlyGPa8GvbU
ZVEz660VxiU02SW8OCvhm7sHtBRGl1ihW0wO3VlVxctje1p8VPaAuFJrlaMr2H2VSvfdOpsfVT5s
MQ3nbUgt9gNdHDSn88XQJS0pyi5225Y0YPvMpXo4OeFp6dipO4TppGUQh/FYYfnxqhPnk4XeC3BP
IK0wZ1UwoCJQMHfnPBW2HHrBJ+iDU9K+CqvTkFf6JrMdoshLJg6SajXlTyFlpoB6i4bZQdFasjW6
VmAo04CAebjvHpglLJbTP61/TBPYpqqyV4fOvQvrNF5WFwuZ38oHppi6D8NRdMB6sJN4c26dQGLl
LummRCbnTHa/DWTAQv+3rrWMl1q+dC3sT12AmbTu3dztTiBwMJfkp0eAoTMsUHJzoMvIQeRQBGD6
/5vhOBtkuXtu+R8zyT7s9q2XkLNY7D/tXA122fnsZGGVV5nidYcA/sYlF3iqfecmBZgpfhIgoiB0
g8x4QGc80HKoV8CC/CdXecPR4eUb5U0yHJSWih7quwQeOoCk1Ipj214FOclDR0eQD8Uye5vr/EHD
XA78T8HS+RrENfRwAlMMKU79disfJRQ48x8nV7yanVKdYaNvRs81jcT9H43By9wqG2WryO8/pyDw
V71rHJYWxjdGG2LLPSVzvPF+QrVlAGEcfuYrfOrDEY3fXBaO6LhWTy1DeJVzmpetlKKNuN4lB0AQ
r5U/ZESGgZBf9fIsuSpMsaA69W9/c0bpfwnsvK36IqNR//oVzFoceFI+YgS8d8t0rcsKwy1OOEwr
bO6Q2+fSjxtKIlSyCRivo82IOJAsJRoFX/Ulfv8GeuyWPpeX1sWrucXRslt/3dmoDWchHtY9lkq8
SLOkj9+1O2DSwOUNgSXwrMANWadEsC9J6WW6rrzYRIqjY2tdhMb5BRAaRnurKM4E6dSgLrvd5xt6
wW9b3yCiAin3+Xpc85eQlYGbOEbqF740KZvsUCnrkN/osb9K2vhrGB8JkUlbU2fJ+2gNE46/YNAw
QMENQt9MWEP5K9iH8koGIpQFzatgfqD/gxYVNcpZFaaUCyrRrQQ1ykXdQNrWdjWJIo180iL+p01s
FJX0J9tyLk7ZzNS/1oa4uwlHKiZJz7L0oUaH/qamthmbf8PTlIdMtvfkNkQE3HRK9rUPC3YZf8id
+op1n4jr5tfuBT4E6tWmqL9uBJ6i8IokQBVXiTGJp2Zbf3JdopNRYi/1ZmSMU1TNTQqqARtF8tcg
XjyTOn2ii5OINghqKSjKmhU1j9d3HHueLBZGb0a/AMt/Jo+Ibv4UsANQHC8qv80tA97byLxOhMMR
L3intcdJJ09JrQb0gKNvEx7xYoTruOFcccST3TTJ6xzQsP9QjJHtuhn2NbuoS1v9xNm9kJN221TS
79QI4VgpwymZxGa4F+++b0cBOuKi8YBBLu5sgVxFLqwjGmSQ4fWSD3u2P/B8SqedHNIsBpIkWnxx
ZRIIC0q88wCa8rBBht+ibYRTEemFg1AkHX4zwy3J65ISnhaN2ELUisx8CmKhEmfTpX8LeI/hlhHS
6XRAcG5O0ZRsQ57EbqVrgCc3ftUVJU+YQTMlXRVhGVKzj1bS4CoEYJgHmGmcLqDruJNVkyBjFPbo
OnTvyWGEPMF67rJiLQfG0NdqXcHCJMWtezfd+ThExRlajFOVHftFNYrGDD14GlsamznSHoAL7fOW
/XlP1fU2Iu0iboclN/dMc6C/VAkmHlsyA2wEVtXBmKjRZO7+YCulFcvgd2KveAugf/UGCJM+vsJc
T1y1r+raAWZlsgnULeahTqH43nShoZapcclWR4CwPpK+OHtKqhQm8dr0FVpdC61MMt4dY8JH+dIi
1lXTHRuwOGstmLFjhIcwWSgdW96PAsOYbqhX2i2V/6U4shMdWUEsgXLZtRpAKiO0cwUrkL51LOom
mgPao274PUvpjOixuhGqbhOXodsijwRNN81nY02nqjW+oG6I0JwlNyFfigPFXxXyPS1pixUD6L1e
PM/NjsQMq/3WWOlVEwE/jI6MBM2jVRePtwzxA7KtBRDGGjbBL8REInxQReNF1j7m0M/etviXkrBb
KKVRQJveqDFA3f9IELJB+3njeSvEWYgnMFRQmKhkXhbHDzWH1x7ywbNq8gJjILjl2j48Rdg0LKyX
Mpt/sE8oHvJPVD5IoaCYm1ilHfzIUoxgBM/Kq6OHrAGt7tP7Gkm7sG+9NGxCEnVwLJYynVQhZpfj
cw6CN61Pe1VZA2Z2Ql+gYvP/O8cyTrg6o4XStEy1MeN3woot+30gw6UAxRBRjVMMumEMHrFC8nkE
gxJ/Yu9JC3hgQtE5CWfC9qUyPKCCHF92yge9aAdLyf3MzbNydHz95NAD9DdlkKaQDNTkpDrqmv7D
eShBBY9E6y7cE3hM0r7th+ikUHTgEBfSyH7/fBOwJty/Ubkb+KmuSTTYi6Uvc1frEfWrgKrRsvf0
fuPi7+3KG4ZxlT4AgYMmA9BXDGmhStEVddjNESZhlD0wVgk4LQaVpagd7GCCZ4uliW4gCE9/pEhU
jE+M8SmG4jxIIw1o8fTot/8KBkKdL6jgt0Uv/JYpt8fFnoGShQeU6Y5ArWzbzFZbLn2KaKrEs0xd
4pdhVouLiwcp0Nqup9/7D5eFmEnVFfCHe4wikR3oehXO5/ZAMaaYmAtLMjNEOqvabFlb5gVxJ8j3
rpeLieuJ3QsKiHZD3ej/hjSK/74cTemj2AYHVIEnDT1oDvdZZ7rvrH6m2a9ZJ4VdakkviaodTobs
1Mgy7sFyB8/dwYZlQ1CAo8UaDfEDMwdTcvmlT6S6Xhm93JQZL3jZAN951nuipckrtUGVycZeFG3e
vDC0KNzMBQT+rdbfLjg6l5ULaW0jz2RD1N1X2tBoeMnNu18JjNXT+jMg4KlGXC7XG9lbQJRjgUQd
qnLVF5qq8DvCS8TDj7VFH87nWO/SHN6p/x3o028pvt3JjaleQojlkdjO42Fv6uH2i2hzHC896VAR
zrotrIBf+Wbt3NkfPxyfmt9cJuWJG1e1s8aC/My6F72ONfjH8SPsJFXd/jQTGEhIXGGAc37kxJ/V
goew2rPwKr3nBewZyMbncLDKI2EscHNBjUUz1himp3rR6Hj03pn1RzlHPQG7f8bs5USmco9LHZc1
aGIy364zIiOFyE76+Et5HvfyIW4exuQVUXoNhGMSBzwWADZNjxQaar8PXlo71izSNVE2p5+PoZ9z
kBcab4IH64zE+PoRRAYScuZKeuhb6vVZgvOXe9ent8IvQZuboToalICaXfFZ3Bp4AEQ9Pw1In2Zk
gEWwA0lgfgWKUlOMTNBJPP22V3ShxZy8Vjxd7dkOPmiaNi7qjvXi2dnqyxsh7epSYjGcB8uh4GL4
gwIbR28P1FfzWRkupCA561EccUBsybCoS+bhoNnwNknSUgV5Mk5dkLaNDIOcQAY/HwDS8CGwvV7B
2RzSjbRmJtO4t7YCR7dSBh0pH4mKn2SRdXmxsgUBP4GVcoaO+8yTkSktsU+DjiNmRoy1yEjqT/5k
es1teTpgbzIFWLZv2s1QUlIiBoISDLA6A1eQlDtiIdsagdaN2nkAoLEguYiJLX+MOhJH/Z3i2sP6
4C7DrTMnwzOdN1AVQCC0s9AIpcaQqDq5Pzesqj28Gvs9AbPGuGJGt8zGprSg0QPVBOfShCo2LV+j
xeqG3YVYnhQWmdpC47aVJh6uCgyXORvcJ6qIo9SrJkLEzAKUlGiKOSOfwe/WEcAsATvYU9aAGCMy
qFPP8Keo4gdBtOibmdoO4Pv6Pm8+WXG9tJ9KE8GqCu4kX0BnEIpV06XX5ZNEvuw4DiDglQP3ommp
TpeCOvhtGsJUl+JZYTenADYCvo+dLwJqx3T3/jNkMcbR/91EmpRJ05C/4erNPFSlGBI3RohHNdj0
MNLL3pQBB8s2/Qc3AH2RaMUgIozmTF5eXLpTdGjGr9lJRqIshsMfVglhDuxsJLanBaoVPHr9W1sB
8dfbuj2Z5y4I6JFpCq9g0CWbnU3mMoNBvsdp5mmhkOv6OLq5aJQ/AztZHrWqXNarHIlKSqciaTBM
pKPO4FgHM1McgbaC3AeN5gI8MHTHi4TmXStrodcIqEnovW3/B/QOTNKiIKAFGfDEr9vWuWvl8pCT
sRICZ9MTfZRUBvgEaTp70Cm+b6b7opoEWXs10vpShe5aqtlsmovz7uN0RbqokkT+GrW4T0NYxd5r
dmUnu/YN7th+IjO53JbyKkYG5cjZilSUtT/RypUV678KCMEH41kxxayjhfgbHz71OHq2aIWsDSzw
ux1PgRTrxwqtW2YrUvsjm1j99PI53Pnqmpi3F5jYCBwUYkatrA5B5CoptG0++aHK9r61hBW6sStP
kjRg0G/yTlgn1CvR/RE67c3ONqscxxP5NsMgAxEuovK5uDGmVjbJaJgvLLtgY9qU0waGFkIF5xNA
UEjyeL9lBWFZ7z9pFYNEAquf1BldbMFLk2LlY/DcjuoVM+G9t176nfJxjmnYm6zsIM3NKqHNR8BQ
5bB9/FWPvdiqESh1+xPxj3PD1ZTHV3GYeIaZVvEMGt0zcES0K6RXO1+IdmIN9MFyVwJXjTFs3bev
Zd2ZTIHoIdtUKbpP6wNJMb3AzqTs00HMneIMF9xFRi5G1Wx6jRsOACDXZkSdYNWRuKx7+O9wLMXr
QZpVMZkA/bbbKayDOX0f10LTKn2a3J1scfSSKaSVJ7gys6+WgbDu1LWX2mH1oGMjT4o2CJaQvZ/C
6lIIJjlRkXxw6A4zN3ZrozrFoDjz97Wguh7s6jGhGcAm0lKujEJURoD1zjeeur2Kvay7mNUbow3r
lYBqcX3I86sfEKX1Z8ssLzzt1UExH1AY/856PrcG2zwPFd/h2z2DtGeXycA1oOekwnyBtWaC36sU
z5JHno9SndgHIXO44kiSMA3UcT24F19ibftU0Rb3tUaWP4WFyhjvMIF18CRdjm20Zl7I3f/f3vtO
BTH/Z68058Gucc7nvSgQEe5hVfw4eXAnJ6f6BN4NC7oYh3gdQGxFfbWqjG+98R1hBJMlZ2+4Dy6j
Df3bQE4D7BeJrZrkkChwAFPu6B4TmB6r+kYi+URmZpS23AoUb8h9GsoZ4V0AA7Dhkpn5+vYqCONQ
zHjZlAOVQnNzeAc1SDZtsYdFuuawNVJNCF0oiHLgV8eKXAxzq2Dqdcnu8kGu//nOAt6NudK0H6Bf
VdLlZKB0M8KgN2DbcQygqjvqOCUdyZgHrvxk7+YROoruFIakMNaInm/9KMb+g2oJ01vvTRCmQRxT
0bhoMYWkQMxAEMmtP7GHnLQH517qqn2M6bDCeMz6dHwfOe8maFZ/LjqH28Js+mEMgM3SrEwFefUv
2fILfMAOpv3ggKC3zM3lbW1UmLWl84Z8fxWFIWdOSusNJaoYaz9D1bpsBiyqyoy9wL7cRJk5a+zl
AydzNwrIi7uDCeN1xzhxsk41XIe9G5OaP9CNoPCY5c9O8DhSAKJXx2Dzchlh3v83GIJ0sHw4SSFY
8oTX32XqIBmpEzMFsQERMrv/jgof6iR/R/AVrHbhj6Zi1Wx6Szv0xEOf1ctF6mdENwory5ZeMoVA
XAjMGsyIwUvUddijbdYAhcem4SHwNfohLsLmjDHp9lO1BMuea4BcAr7CsY6dTAV5ZUsQhUH52Cyc
yDuB6e9W0fo5iKiqJVDOqYF78HZdp6UfpBeefP/NOOY5EPJApTK8kTLAx4DaZSVkTQhB6jJVVpXf
yU7MdqQxT/+6UV3OyuU4n3DOVWH945PkW+oo7vC1l2/jambHE/WjXwAD799GYYd8kmJXoLOugOzX
2l25Kk+Eg4O2SnU5actixC7XW5quBes9kzFUeuV/NJSKJxtzqdPX16mmEfTLgm0884iGVE7Qg9uj
Ay+szgiZ+ifSdikykdsX8LvHjjGDySYsTktk6qC+3TgtJebXRjcDvWETI5R/K85BfMKvJ5IBqZac
IkQh71/KCrXnMOu1+i3uj3NFi4Muw/WrgHCYvIbt+j7AVMYKdU7oEBdGpg1E6MbnvWTBLBc5l+lz
4SSw/p6T06XPxPJQ3dpNC1QN4Dbc0cjGRjcFPWxspL7+b7tIQjkEhvnpm1SHMBDyJ3nZRK8x5wKR
i5BCdjyUnLWGxSzpJuAhz5g8/6FAj1tMGDtNQGZv3yic4dllzUqcvmeqyY5SdCluOaiXW5V+HwKb
Z6Q79Lbv9/YG24+zZDH2rOj/FejpGblvw+iqyzAcyxJj5Da8z5YY8czhR9yGPPsdIGdIz86k/6eU
EUb9ei6LqVlTVks8nlHTuyd5Pv+rurIB1cJmSrh/MR2KdKZtmkw0nc5pXWE++LKzqsVbyF2Lrtwm
cXFui3wGoOp4ZuZvwz+UlNTi/moQpzOjLyftAz3WaDJ64aa1ekfp0ImJ9aTbJCEnuCJsPv5kzGj6
lhxEQfVyvBuTQhYBOeH6pI34hFwDMB8DLJh+i9ONSDl01BrZySQqqsEj5dX9qEcBsgcNOAgadQ6u
Wd3lTWUbNdS1RSBtrCW8/OkSqnptuJwSyCZuxPViJQB2TftMhC6Ti4kfYkRmX+gGsnCeLsuata4n
zA/5hVw8V64wmYLRI5Xb5/gYlDSWTMN+YrMZXDA8qaByO4Nf1jfbEME2ClQho6s44X6jJHOBNP43
DMJRH+cnR4/ljNdXQ8asuiiS9SzqAwWlPfwf2OKGzLvxBFioPNSUpiipzbCNR/wxJKlZtq9zWoxS
b5Q0inmPbGNFKU9ZqE4vqXiS2MC+yR/evFTHF/hv0kixMszI2sTuS2QaEMPgxhCJ5AMrGX2P6y2N
eiN9gbrEc/8B5INg63qYdZ5hSedDIes2a21wZ1YaXOHCracBK0nD61V2P40cioWv0BoRgnsgVVy3
cOtWPGHIoS8dDDLnJCi3w9SRYIGVrZqSCcfBYvxVVvhJA7Tvfre/1gZJ3jLGef7AadUNScJc5zW9
NDcyLZI9voDtvmG+dBXMFEAfudX+oCA5bcoIQJla2LpIq6w1kS++8syEB/z48Jy0A1Gsj/qTxXuV
lH8k98WRPdT29a6AMuwgXU35zUemSjcHe4suzU7NLmUsr6TH+P2xqeKa2K23Luj1UMWYY8lho1/O
uYC3QOf7U5op9QzgnTeBP/ze45GWb8OKnNKP8EFEA5cRHe9YTq1XgH8tGG1qz+iElz5v8du4szEi
HvXrHH/VLjVTOnBbebZpM+haPwiEBWYpHnDGK1R/M3OPJ7QSeX1BvlFrA1zW27Uu02gmZJzCnMql
1/LH3xdQkFcyDJvXsVqhWpWMePds2tew7qJ81AOVoHMQRFlkGH2uaNGXl5Ii4Pu1eH+QwZGF9tcT
xy4s06LMkzcuUzNtfHZ3rfKUohFr/0kV/9KMiM6YSMh78oLGmZgAzkd0rS42GJSHUGmbsAqE2rqo
OyckXWyjpiQ8Yy/cRI3ywgm2SEVnCwMa4beUEuocR8WjGqgcpi8q+ZHRVQCtno4UuFj0wXi6l+Yv
VvNn0nVS7AuMXx1J5Qc+zSrHw+RQSt0Eeba2qVX72l8n7VLyYFVRFoYrAgeXoDPp0envA9HNwNLv
HqDGtGteZIxNOlcgWBqa2Rg5gisdS0EQSynoFjAHT+T+Dxe9gE2jbSavsg6DsY75I0riBj+TwoQR
B+Tj8NLuVudvUiKvlMjTyEVFhPu3twUsz0lnPM7zOqcQAvl78EiDBBwu0K0QJrtRlA0ELeNI7tc6
KHA4Txdaju0BWNHB2YTV0MRNBFzEX3u8zPazXFiTWLHBxKJEuCOpgyhh/AEeYnyFF0lutfQq1LJC
GNJ3IOYjNpBvZkUypG0kXKSVU4Bul0MdZG1Ad68cEukYjsaIMTcGBBWU7Z2YDNLKxFuk3oDpqz6f
a75AafD2p0VmQeUZnw3GpwkGQxhL1zKZfTlrACcyrgrfk0QCEz6N/2d+Le1kYuUBysJwVYm7JcHf
vrj/wrXffv8fbl1rH/EA4e6dlKRVQWd+4k7KJeDNNwGd12y6lOMvBb9VwQ3ehhvo756ZKMom/uhV
5sWdEP3PKn72A27PsANB+ukxFQ5fasX2klh5fpvtgRjzSAZw3B/OSVnkHAMuonRTHW3OY5o5ZJ77
e/uu1tj9npIhnmV9P8lUBS3k18sx/yQcThcZE9f7x9g3kujiwHWrDYohiCecwHAf999UrFQG9KNn
y1rJBS2XV1PZI7CmF57J/3RP+lrWaDCmSeulRNCi7Y42PF/B5M2PyAMWfjccM0u9jSyv75vMNeJz
eNK/ZaOxuLjLK7C3z56DOKXVYnJUj8SPRlKaKvCJ3NCvrvBWfaGprhzdv1fNhW6AteGcxW+6iXqB
UKz7WI0bFyLETE5OwzdRX51uNS+7T13Bsgldye8ZUT20M16Ai0aHF1jfL37RckQmhzdu0vRLnCN+
k+IiA/nDy1WNuoIpIzS6QiJC4bx4C1j5HWRDTm5hf5+QmH/+lbGb8NY83nK6zTYdwX3Q3ANIBs73
cYdG3AkWyNK9qioh1dDUdjhKeLGQ5Q9RxY//UjIum3P7Fq+EpKtxa/Ir+fF4/V8YD7RI3Mycaze6
7C9hVW89nZcu4tu52d76pMYhzBwj/yuQGoeo02K2QktkBleGrzCzXAZ+MLOQd+55AEWTupyTEbam
R3mpZiNNE3cV10n4UT2x7ZQWl3Hjd+7mu/zlXcLx0b0VaI1ayGdm/Othv7D9XKv+FMd1GvG+nzoa
YxLNalH9k8vUOKI1JwWFYqJWL1ZZBt4LbZIu+qhFnQRyb2mVZqtIfxYHf1ElHosMs2X9h5OOM0jJ
xvPzAz5pCRFFoTQr2vQvdwawq/68HUuwtUlhD8L2DxEHmh1VsqpdV3ueBP0oiqvIlwy+Oe5dyR9E
aJ6aeCPTijCN+bOhhcApyGCefjDoKlKQlqz0E24hUvBiqEvc6LScbs4I6fPnYOzUQuZ5hPKovmoY
B73PLDo5iIum4xSRRqATCA+6wRzlVpUL+AaNCz6MYbifG5WgGWK1Nuv16tWrOuA7++2i+liiDNID
qlcetTupWaaOGL+GZbG98X8MV862OMe/BXzn8e9pPkupzQ24agesTbnzlHhv+SyDotfdKd0SsI/x
5oBc6tDdqQAEPuzWadrnDXPc7eTyC7E1u/XN4TaiqFT+sVpaISgqCkLhXJdrxZOMhHc56imOASqx
AjMu1tzNkKehZ//tw68XWhs7A2NLDEuKUh0HYsW3YaoGXVfOgPVWOr+4s6M9E4faI0592nEXmvjY
42yvmz7U3GVzq8iOI2KmZgpnN6bONNpJndNCCdtDJNv2D9hwNTHOHZ+6YSVoYEkVqPqUlExCVpgC
jiB2Ha6DCcE0pkenWwtx6JxRK/wZsIljd2FwrVscozYdo6UJTjL3Jtp8EJA5Sb+Stn83Cr78jmt9
F41CY64T+Bb2r0KdmDKpUdBFHgVzlz12i67KGgZ9LSo0zAHPm1pZ0w10tdb/yaBLnaNsGQ4XSlrV
njdiIc2lVdWkfe+tP2TFC3Z6OLT0AZHPge/SFiexRNI1ii6UhDThhF8zi5SeMD88r1B9px1527V5
4NzCHVfS95JOApgx1JKT3uhAqbGtyH4lY8u0/nlC1buJQOVx2Oh3FPpM9i2Gn2aMrtxfeB3NwJIs
rlWLsRfv/pNa6jEn4OL+mn1irTPU/JdCiHy9P9j072EpoujW2m3yfz/quylrQlOfLTQE6S/y6gqy
Lfk3ZvwdFAn36AI2xNnaDKA4HRn1n7NbaIXSAE0uHvkUcZKNFL9PG22PpK+XcrlwGBcZmVZ8cM63
2qQKF3WEjSFfPmVY+68meeuDgsaR4TKEQrYljd9AW/QYYHrneiBXKTycEJ1m1BweM9Vmelr++JAk
HYQyV3f7dCmUuyWGotHJU9IdkYn5vZ5FOL5hBTIVJPN3UuG+l4+Zt1/uQ6ee3r0AMl9IkELV2GnY
0qtDMyZq+jAWMDfrGRf3iYHMx9Uv7BKwq6k+mXxfE0crs7eaaCHQoLCZRZiWLRFdpLwQgjbLL4nK
Q6ZdqtpreKF1JQ6v9cBCV6V+3KX91g+rsQsFB6GLlxsz93S0zSF1vBKo3LSLZHrG0GsCaKVs+QpS
8nuqgIZFWIDF9BAq8k4HEeVQ4UzhU/yMMn9gasvXKCHvjJgZw92fXWrrhJgNcmpoowiBK9yV3zUX
0TsZwy+Tj16ef7V3fJ8tcq8VMLowOvH642kJxDYCrXX3IGDmpnt/E4qBDAvMBft1wDeYWVaDrJ3P
6uRkBm2SQ7Sq+qisVTH2rF0UKRNr04B0RHhu6Iueb5Lp/UqMSD6EplKy4+mqTe+irTH61ksfTWTw
qwDZmwnP85tv22Bz7Zx3ES1G+DaD38nwf/MSeVyq70yYkNImuEOdz/I5EJD3fLDkW2V4CnJBWPSp
zRseMcInAovVX3MRJNzx6w6PC1ZnQMlf75lBo9wOXdrcExp1nMZaym59LGTyyts6HriQXa1Hikv+
EGQ2y4vexQOvrU3yhUjgeo0scmf6SDhJ54XXHpFkwJ0qUv0pK6aUAbutulRAPXwiDSk6wU1QxNf6
Gy/Rd5MvLRZC0N2TgByTAb79JDhlf9wDOgeAkuob7X7e7mIQnIoE0PeyZtmtg1SgkkcS5KfnTER3
oTXZHfZFP4/1Rs1deC81W7LV2WkcYH2WAUkafaPzbbUIln5xAiJXRvF3l3hEcpg/zC+qretAe0/C
F7hdNcXC8mbXHna10sXKsxDx8acadiPBcVpAsBsqKYbhJYr3AbPBBxjj6KBXVd1kQMC1gMwSu/hs
3PD8SnB/yEPJkKEPKh0Z7wKSHR4CFecG5VrNKiEPwAwSjmoLrvarYKyPUbU6JtBll6YdJXUam14M
7T3I8VrC3gPqI8I002gyfYS+cFf3jB1hATvlfhpVKWiG7A5Ldd9SAl7vk6olJ3p76HP3k0jUqRzI
UB9P8iaojV3qIy3LCWHdXqIPp1lB+rJYJ/aEYLXqKOi0TmTlmHUoODVrWkOlM6Fl485ZF2Bhych8
CZ6L2ictoXUnQ/njJtDGCE2mwWU8E/rlIyHkYgvGUxm4uGKMK+QmLVYghwNzOAiczl99OKQatIMg
xZ7ZzJB6pm9WgASnTMZWZ2YTVLFGKB+iEadIHatyjgXnVjkldjdEX0vEpK8MeN3Xu5sbTH2EpsLa
e7oJnNuYu/9ucyOKQ9rfw0jNXHMHEbeLvfr7BTKBOM2RWNrcpntNJmHg4Z89VyKk/xazaykRXsp2
Rylb9G3Sn818brfiVKFGqsOqbJWmdtqHHc4pWKyJTxN4uFNMccGHBocFv/D5/yu5sQ7vmMKZzB08
eXsv0krpgS4+72/xg0jX0NiieYOM3EU/zzF1MZOhpbqmqX7sbuDQ70QrRHffFur+PA1HGgKb4V44
ElEair6pkCYqjLkaklmaFPJ9+Ss/v+3wdW4D2gFxv8Z4dhyICpUz8mTZA+ZZzJYKDbtQxkRm2bGp
SIS7yBCi8BgiCvcCJkzWsGjm4WFXfKAS4+xI68Sm/fldJuwnoTiRsfvHQbxUxczEmWKOC1hw71QN
rhjoV/sWmmWejrh3sRlw5Iq7nenUkfytkUI2Abjm7Z8EifI6HYP+GtRSH7fG1yT2nAeroEDcEf+S
WkpdDK7P+33Sauxs5p4lu7Tf3C/oCYX5bX9LHHF54cTE1W8m0szViVNzs0Gq0PfpbYCrh3tGDqiV
gXOLM9Zj/OixnYRwutY18GYWT3DQRGt53D4xq0Vge1Y3lAK+lMO739WQX8iDvOgbmCNPKk7y4EKL
V1l3ueZl24UYQgP+RW7VfLCgFEZtG3yOuYrV5cxSWl5e7zGlKmWwcm/YbDz07RVoZxDCkPwHd+/N
2R62VczmgL9KXFtrlX0HG8+yQlehFcM5YMqOAJJRHc1Iq8jilCfP+IilT/kcog/QbjgbKOPRzxRo
f2A3i/LbVoxvwliApdkBF8fystW5s6GwivnXDG3KKqvdeE+F6tVGQX1PjXag2xiLdNXNEwRH306E
XtpCgnBBdEB+XgtGhxGoEzfQa+WcVlrlU/fXCkhWALzkn5QKeVWq53U4JLam3nqqW3WtWfO8C/4u
xCrA5RRGnVlQSDDxETyVEq6ZvhnBsshe+HLCe3wKToKWlzIbHCZRRz0qxFLGX9kVzb34vXYQ1Soq
4+G4/l6sAmdl+FXSRJN1H7G/7ldCQND7LJ3MExkqMtGzedbrogl1oDk7hAAp4gj/7SLZ8/8222y3
7MM18v02SGxgI8fYAO6ycAETJzgrzz/+uIXWKAJKz7rBwvvjq1kCPwWqBUPUXVdsH6ol0j+o+wdi
CKjTuhohSC9fogjQnvr1GXAFaxKH8Wpg2So0YDt/b+QLuYJIYXpgcAxhgKXxBSwZxifK4iOSuht9
ThjtptC6AZdbJHk4tcH2ykFr3558xQ3HNY9HaKVGIUd45xWo2gWJ5QDlsYByVyTOuPy/G9HImttp
K07cSP/HqmQ8a2ins4RLyRhU2xJl5GUFEGqX6DlcaLXm9crvyyc4JP1FvHzjbiaTgy8Z/xmjF02i
CaeGbTx9y4nWCQnn2FJGIWl7isVXY8LH+oJ8sS4BnW5Q2DEKfJAQu71zHIOpntPMOxClWDPjAndB
waK2eU/jeoj5dyTfOQsdADdUwg0fYZ8M5PDGg2IUtLkK6LdyRhrsd+0cOeHKCktKyySzN4IohaT3
73vrpvVlGPWE3XXQXNk9BF+Qq2BSaLPUB71yU60fF9Bm/BW8DqbDwxbVVBJCt/ERYhdI2rp1LSdU
9vv6V+DHJT2vdCFoudJSXZby72Z38N5vBymgKIbMu8R40f+oKiowajq9zJaq8ZlTuRTJOJUebp18
OOIfuu6SJ7ZxSp2LroYjqSZkaOSiUyin/v85wOkgkScW23HYZHD1wb0bq3jsJ7ZgTvZ292kLPH+o
yTm7ql96KS3QKwp/W2ckcbh/cfqzs2w9toA814OJTlphiQ3/4pI9MPQXK9DFjV2AuO/9D8oGBOUe
kgc3I3RxP9bUzAz1uzIgzSzVgS+9f+yQzxbh7bIfcUyDJQfqTr5JeeABL9E8t//4CD4bSBWc9GSI
8AkBkEb1sFVzJljcXOWrWGZzdFoL/huuiKWyE9BoYSQOYCVVzKEJQAXQFOc1JVQo5XRv5UMFB082
6vScGKYKjZsVaKAJ9kph+JfyeFukLQDara4wIKWFF6nVni1PPUblCWzUADTv5CmbxMN/bgJIrSaj
7gJzCIKfe7k0zSaAqaIZE2a9jvg3G2SOuDcwqMfA+RCj+AuSwHlYh7iSfkyIw5TM1B8GFvPBS8KM
oF4FXaEjB+2x4faF4GxSjSgVu0rXvSALhB08TYst0JR/SZP7Wrm2qy4ldptamgIFjub9Avif8PnF
aR6czWWU5MstMsXg4o7d2LJAw3192Anxr1FJxvha7u9b8lh9kwmxFMPPSAdaada2hBw05Fgi3mpm
NZsSWFmnkjw7NRLCPHVeSXe+pe/lQ73Dqud2tGalsgKDaBu4CB+mc/sSdyupvxkSPeiCT9rKp7Kp
3CZHl+cktihL2rADbm5dRG/B+dUzK9GFCyF5FBVECMBO3wdUDOwPmmFV1X85FcVUQwEbrM6KaVJ+
YjjLpKtlWJ5BU9M9P6Ri+LwiEL7Mg1Xbcg9jXaRER8s3lprwtkjx8yDz8pcYrtK9kXmmmK5d4vZQ
W7FP/RuyRLzNVIHoZPYsiDQceBtXhDknS0vaWITSQC9BK0PsfJBRjdi+LVjo3zh98rrhFazPXb1e
rXafP1H6uVA9bzxPVlj9acoC5IqcT8wLcDq1D2HMUdm2B42Ir+Yj1SlW8wpmK+R4hHTXCD7kPHS8
iEzccELxiYkHMDDyBMg5q/d9jqsiaWFbJbpVAXKaitEP3OTcQjiArPX3nd3gjXSK/flCHlw5BxBT
JbLJFbCq+Z/Pf8h5D2dtBg+JXV63xFkm9xzq5BK2eK59E0ntGNObpGCLG5h29Apvo+vEJbOhYlAO
lDh2Q9KZBxdnDUgOtscypCEY6QcKpOZa+wxi1Mg1C5ZxXt40Nfnu8flmUQ/p2mcw1yTHURUVPJi+
klvfrrMD7SHZj7zdAguAhY96gEk4cSAv6Yz1GuZ49ezBI5kArQ1gLFlxmcjE9fnlPBkXN930cHxb
XIH1z54KSmSaSnxYHOIDjL/cBB2CwYH04Xm9Ev8A23rYYV/IPdAMjqCOAzwpUsJpwAvqEHWs/1m/
KTRq9gqTd2KwX2xua+c3tAjTnRSIEbi2rAYKmb7sH4uAiyFCoiDGXMv08SvFqBvo1gcyZ9yvltTS
ovxokxzoy1E6RBDAtnmWkfhMwkiYEpabwk/JobeCBbpE+I1TROjCfQwOf2uv8wWWvY+RrZVug3Vg
MKSFAMTmbXKQqIRnMXloDw8/4sZaaNFYlYjhojMNy11QYKiXqvPL1MHByX5A5EZbM2BVRkLF3LSQ
PmCdoaAXVj0DWqekSS7rb0OkUMbNgpx+5d17UIMt9nDZbwSOt2qE4dvE4EGB6OJsHi/o57QhnuOn
qUVfdQad+Y8tsdYzJ7hJn79231/5pWMsq/1LBRYpRuap6xYfjKxfwwLR8NNG8/aLdzn77U8GKSnt
Lvv6Pp9LRr3Fsn6bf5RjMySgBPCNpJKMTF7mBKJNKAlAnqNkt7tL5Un6Y/ULZaE1rt4Io/bM1Txb
eWkO+XB5QZv/sgAVM65/rk4Yckew2xZwqhewa/4WSYpApMNBF/IZqlCNV4febayIIzFxqY+Dl0DW
24Wh2mSvCTxUit57CvWOutNHv3FdM0GZpHjexhCz3SnIRoXpRpR1F0FPIdtXU9y6NG8GU2U22AB7
6Bf5EbywwmBvwPQEgOhpEBJ+3QFdepxoZY+zIClYMmeVKuENpYkLKs/PF/lZmK8IyRt73Kr4DTjh
zWlg7enN0QGJwahHNkld9exefSl48k9JDeTwyLPmMUH5fOH9RHTl2oCkl1wVikVqDZft0Y5RImYU
4JsghT1qPhVieOzeXXtPvXGW3gXmp7/Ud5kYwrr07ccvTQ1s4xNu2K6Nh+eity6NjtdhM4GTuSpn
iMLnfSXGhrdvFuqrimkxAil5k5cTJmRbBZC6YhFJx6UbAYLWIckKg5PQDxudcSu9x6XgtoVMvAq0
gb/zGM8HrEK18U347xsSODTXZrTA8xeoIiuwA7yDfPENVQlvTJpZViTr02Cj4mfLtE2tXOc31YLQ
XTDvIqJRrV2IVl4KYLoQnIKOtqamfBrXskbaLvNUWryfbLpP3u4DkLg+uhW30n6tUguQ600pmdKQ
c3IjhV0ZTc+ElxS2gw/itAkzE93I7QPQcqAawfbPcPxuOclLaXSjimXxGiLv4dAsta/pceT5Helr
tVAq02E2oGt61TEMi75X0D+ye5jt2JMauoqhKSM/TxX5HMwtYr50Atw6EN4Q0oW76h+2jtZ5dNnl
O3Oi64ElX+ebR9oE4H8tF/vaUnG0+49Mukijyw80rO9qeIUgSows05CrHEomFyKos3ipVGbbkhFL
3sHxZQ8SeVCPV4XGA6kcIuD278VKf6HDR+1JX/H77FubMbBDnelYEuHDy+mwSXM6FfhPdewIMS4F
ALAtLWrnMKv6MOrITBf/ozyT+3nm4sIdvRtGoVDveyE4wFXPKKXT8hjI89ppGk/4v3f68mSECF7t
EGU9jxyptuzkW13dROVznV9u8hx+/Uh3I1jU7zzGBTdTH1HnOYfNjATrGHImuqmnjLUPE2UcmqUa
CxaU5YaRWzfaslT/7gp0d8GI/OuyM5UdQ/Gf4TI7TsRtemXyAyFls6Fbu8eOwGVX3sfBhV6Gwjjc
2Xe9ogtlJ5R2O/8jhOzgqEgRx0EOafMR+/7juGRaPOJvM9JCwJxD1sYyshY+/qgW+3+euHNQtgTY
p3gM12PxaWNrExf3dGYoIIgXu0rU93JBlPwinHWwfRBuul2L7/hPEsm9+4xbzL3z6SlVbKNr3cn3
Rj5LyHKqxYCXSsVEwX4NUVKbXfdIct6Lp22LwZlQYoyt9X7oxg5/egwMQIYtQb0kV+hNYGt2MqBf
NQLvlaMXSXmf/4xtceia9YsgdoZb2HM7Y0dLsQBOe0eHE2/wJ7/VbJkVo/olxcWMr9PfK78153YA
NmHIXW7ACS7xb2po7KARPkriHhk1Kyv/rgpPvQL5Vz2V0l/OD1W/lW9lhIGzNTqjCCWdJb2Gf9+L
DntAejtjkKngbUal9WZ7uzEAh3+VCJF6vtfr8YG0kqUBWsgssky9jghVYhmjcj9WXXD7pJo8eg8+
ke390NeoWr9spjS9fjF7idj5bi8lCy1jus40FUup8sd5qOOWZZsdN/pzhE3m9HfrscesaAfpwiUi
gIDGVPEstTO/uk2zAVAvZ4eCt7dSA4bLQmvLk5nYK3XOxdWvyh3zUeEWkw6VvH58XsVC7Vpff8by
3n3Xe3LHJuWr7+OBampL7KpuJk++LLEw94/HL6NbrlDEk3q+8Coy2wKTz2giPW28w3+tbDXrrB4U
o24ytHMbqxrGwBGTsqAq1o5TpSdyrUtTYOBe6aLYsLSwU6X1gSNgHcsbg4myFCdw4r9BCDGgzqjG
7fjQ6z/WWFFSCkVZq2AQbLVg3PbxDahFiI25Jcf/AX5pKsJtrdQmSju7Utajwb4/YFyELpMou2on
/AyQCXT8sy4VH0mxARmlS3C6DC57xDL0flP2aAnbdqo3Z3k0FkKH+ZXXrY4SMMGrDd8ecasu/R/0
Hg9ZkOh8+wwTmWrZb1HqhWQh4aH/c1D7fX0AM1lh+xugI/QZxYnvNKvzP1d4QEtITkXAajYmFghS
yNvcgobBx3K2ZAsYk/umOepcI/MR0E+S8YHR1WBzn9dDS5wgDsshjCjgih8BrOxACLbMfdfbu+G/
8eXdK0f28CARyVY/6btkLcq9Li6yDLGUK9uCa/j1M86s7I24CwbNxqQfQDRKsR67PCsjDUbZMbnH
4GaEMwqmL3KJM8PpLqgABQ/aSKcaQrlkZFXnOBILYvxzLLL7WA8Xw4M6qMmrNEcW6nl93XmkCVQ6
oA1M332T3B0bK3y0AMG/oErdhMK9vafTzXi3upD4UC8OX6xjAhIL2tRMltdd3TXUPZLGZ2YcEbPu
2O/VVLhnm4uH5MOyTuIeMH8eSCX6VTZLs8eDXu4mTnz1tGIqrzrCjjFBHIopI5KpWSmdR3iC9ala
6WnyC437mKGBaCGAYYhjTlvIOH01TKEJajouSoze2ZgVwWXzz97RHRkaUOqIQ5XQJxWJSU84Lm+u
Q//6ZCnEQrbITbYNpuqPBLG/+qkcg5WO4+rmOjEel9WGixENR2tCqropICCCuWPD/Bn5e6qYakVc
OC32ViIqCKg8HgsQ3SNby6+b1fK/wTlS/7cD2XGCFKHsw1dhRtwO/AjNT5oV8OeK7DtlQrOQ7cTx
wD9SZ/32740iIwZfhoty8+4lczN1Aa0nd0+7qJ1uo52sNE7x1TDyT4a8J/WiiFr/Il3J/4xh33Tn
W3IraPKR37LyLMLYukCwvFd9NNYfL+ob5amgj/tTVTGSHpaKT/6PVvyw4YbWnG76U4RHzehhlhPH
W1qV8GPXzeeQLQG8KvscT63kvrIjszytRZMaqwCWIo1nxBMnKDo0RDHtCAM+eg3qH5m2TYz1Anym
r/kP7qyZ54lPh+y+rvRMEaU+b4PFRrjYSP+zQZoWIIVANUY1ir5soDwmUcNVFrLFcnjuUxrVA9OU
wo+9ujrFXAlNudjyt17O59UN6dUhpXNWAVKxY6nES9it76qNscZqxbC3VLHZvxrxUpCAcN9jTP1F
Qs1i8fAs3kLcqthgLoIFWlgn1z+oHJSrOpBGRrPFtiSkSB0z6/ruaVtMn+IpZFc0fAGwtWYHkIr2
vuEY9djmGtOaP6cHupBOPX81aypyYq29RDyFLHiGeYJ0uhBatYVimdufkeEXrE9kI2yAiabR5Fyz
dSByI3Ej8YZRW7OvtvP+gnTRE/WWNgOJbqEQW3mOP/1+JVGv+3IZKMrEuMZZUCvmxfpwqXNA/51g
ZHEWR/O566XKx6PWw2jltEdw8FiMNCyzmNmciLEIKZL2aXdqmrURjnUN8yTVKJBCZJQYjuibWAvB
6jXDh7d97autj3m68SkuEbM/GsqQy/UDsuEXOAuf5JbtXsJFt5C8+2hwEYG+iZqR31jJyvllp+jA
42cHOXmLNIVmBmw3pH8Mn79bNvuY0hnKJxF84BATZa9jJfTsFPr2tznzNMiApjhNeqHcCPHHs4ua
4SieVBzeTMlTLHUYHOOE0JxxymO4+rqjOtl2EtY36VD0DQFij2qID842FSeb2lDyudsZG/FrrXkc
WnqO5NC5OfMbogppYeHVEWsjdE719jkPHn+lmH4PLn8h3fukfJ00kt/dbq0GEOOKUa8E9PAHOEJx
sBSpI+8o8MkS87oMoHsueaBMQv2Hj82OE76aHDaIaenMqGveScagkVBn0g319KePcaEjqsxOjXq5
cGKOydcKdWJfEjKPgGU/Tg5k9pSQHemJZIXzMHBovOwF3dC9Nw8SE9sV/h+cObicB0w4a7qC0Qww
N3mCnvLS6iUT1g76x8x64eRpGNbq/9imX/cm4I5gIlXd1bsMF1ox5aCPFExnNQ7wMeQIKAIW2r7U
UMmV5COA51sgpELpnWYIaqFKyEqBc30aTM3Ocs/AJ6+O/+c43o+OClk1oAGNZoep/GiGiTOTz9SN
OSSydopItiZqnFCmcvVBdo4SI1uCyo9PCxa9jMd82AWQ0UFJxAYyJ/sKwpU/qb2QaXtzByqAqvoB
X7Qqr4sUT9nJ1Fa1q3aDR4R9z21j1VqaPeUoKYFak9w+cWcEFO1GjCKnY2lN/tuUOJxEI7grr24N
SHUEUhrf7Q1dSJME/3aCG+OZMMZU6Ji8Mxvprv/GULZNZDbzc61a11J0ge8aPZMimgCJR0Nbz4Yl
T7YfiuhMcN2FS0WjSiR15+GDgpfq4z1tGgHToA6ZTtQgVn7InG6jXWYAOGTGSifY0mny6EiGJa/w
rOXLMKJLSUcPg65U7Ck5vH2tgQJGT9pMlduoxKfTjNFq/d6ASd64XsNq60fQD1UmiuTpKhj5HG/r
jfSS1QKp+9YoKoW0aNaRzrjsmlxRL+Tq7CiJ+sQ+Ozf+Gc6+2k1Sz7iq7R7NjXxyXZA1gMVzBd9k
T5mrV3aIyn/z8T4nitcxSJdrUFGw3zlw4dIlofHqmcp88TycAgACXeQc70QDkaY0wmRou7hUMOCs
NjzRK/VdVHXn6sMDU1MQmieKm98wr7FDZszx72Gbc0A3wm2bgOBF3JIcbBEEUUJJwPbfbK3RavNn
npaZPfB8wiPFl0/5Lcg1Q/CLNn6bTMaWWmUTB+fCaRpw0kHj+jE0WBiFagfrYVffXzvDkuVM18IT
Q1MUp1GqO9KLmKT9gg+a0a6+JDPR53R3mBmTHlQ9rChyVQcMjlzyJqWI3csgrULkiBb7fuCJ1S9y
W4OWcacOV9rEBwIImb3qKZr3Q32xnm1+fCnuL2ezkFH/L8jsgJwqQ80/jMNh838IqZfw6bLSMJZm
xEzZb4QplqSUqqWHIbVLSdV+dvDr/5gkf2IPQeq+5BcdnREiXoMwFb1yYEGwwYwY6loY+ch1/NMe
SgWT0aACFc7RR7tg2eVSVrqf8p1rLdzDDCtbnNEfRZNOUdmSvovjjliimQftlcoAbb5FsceNkt78
Jqzw82I4IBxH/ucZq5buZXLfvg2ddI1TflaQrj8DDIBnbg1LRuslE9jReXe6I6j9N/WGAVnT4g9z
CK+2qG4a6ngdXQEKCyL/ESh8diklycazu0DMuiU61O62RSntvFE5c9yH946eU3cWoQmTOyDOK2ZI
zjcL3o6uIh9WhymrkGi8xhoTm1oUMKoBPI0vCXNVF/ZfQqUmXNgah/RJtCixc10316BB/oUEqlUz
TS9TG4C2LsuqGiUWea0M0wAYUwbH5Rh+Kbsf1S2BfMurr4Nrtq5uqgROjN4cai4k7ksfvfd0Eo4G
eTTKMrTMfSHjDzJeXdj7wXcSbUPT55+NoyCbKPV7Ed3u7aJ1/gn7VIPcQk82+6khpYiExfAQHBoJ
YBoCcLHRRG/b44aHndjA/7ObBpf+JauTws4hAnr7zzj1GO9KNRMXT9306GK9UBCXXVpAfGaT/duQ
G1wvCAXyt55rBShga7XDsHF2nmNxLOVTKQCq0nCF6HnUSlaCNHuLDWHkJvaJaN2DmyfwJXMLLEHQ
kaaFlLHTBo+fvgjVMkuHR5X7S92c41k95ABrH9HIzJkA/D3r3KkFJ5ajP471xYvieIqM+DW0QKrF
YW9IwIfrlnN2CnSYz4ihj6W2TKvPfVEevk0s2ef0P6A2j5VE3vlwePVoLvvFkV4b3uckmNrVBSDn
YeAx8AGLLAjUn3INMhoz49BTI89qSyIuqI8yvKI8sXuG4OIBm9afFytmXPL0D8sAEP1skzSCA5jH
g5GZNwSYeON/AqlyZeoftG6RBIfFdLN3mFgH6LH7z1KM6+5FtjVPvBC2M4V9rygewwlUTn3JwN3G
P4NpkK+fPI1WG3jyMRkQYjItpvFAxUc66nRzNF3RQJhWhwRo6wXaRY/glFE6JiD58qDwu1m4Uur2
riKQdoNyMMPSCYyDy9ReFXcujqu9OuwQ0aHuTkn5XSa64vj1de6MSA99x5BSX9c3XWwPhe5K1gw8
UiZYW7DYEp8nI4tIekyHzGRpz308GOqXeyOEBlaD5//AXPCJV7hg1wmMlEzMKCwVek7Z+C/KmaxF
+8bBCgaZDn8lNhNix7glzXY0tpxC5BZMwBcy90GHqaL/3ujCAryP5IJ/VRK2ZIwDtdfR/xtkuT34
SihokMz4v9zNFoiSY2pR8GXB7+NRfCyYV4wuZjh2NGqV0oSICdBaRSFxsq4UnYK6LMOpWJqeBRG9
zHBxeWvRDNdoS7LynVpYEzE0dVnIThfoZ2Eqq4UvSTaO5xH4NK79hC/s2bKsUQ2naspBz+uLc8ON
6NKTLLLALQlrtxWEeGdrqihY/IFdzpb886gAvbhgC5ymkezhTnjwWv2XL6lfK5EQVKCsL9iy6veM
Qr3qHHxfHWAhQSqr9Pvq04UDXS0RwqQ0ZarbZvXxL7zRYG226NfPj8HIA+ZHudgbc+q7o8NUFtC1
7NuG432eEKXUxygf/ThDcuUa7mVcZE8i6QLAukG/EJIa2tI30kHVoyHa9l4JtlMxWtY4At5wPJAe
Q+mvTwUDaesSkXLWAuJ/wDDDn6aOOX67zYbHukwzR2z2OAUcnpgYJb3gU9iY36JIVP5rY0UwM+Ki
TBPHAxByXtVFncd5mQM1U+ALgIB3y6y+iIDEnFP/RYnUy2N/wqa7cpnbYs1w3hdofz1wAp5DFZYB
uxujCcP0cKxqe2XqRyMaJZQ8nWe37SsOy0OqwGFLkM+ugKErn2ppXMAyonFsISt8WX5nBo43EQ7a
taSKrGpMUO1ljeHePJydREbyziq8NtM03fkXJuTVeQK82rXuZ/8CEynxkMzlu24Wk97TsTyeRGvG
Gzs20t1wZ7/uRuPB0fECpXCRAAEwUCkUO7P4H8TNpqeCqQfRfbBLoxTVE6wnPY15sFvHRYVeDb+h
AEtWk4TFWkp49le8hXImM8ubrA2z9KyrGWxptBq92TPhyZB9pFqBP3ZNJDnGdEHkFR8SH9+VlXDg
tEMoEktZAcCG/bi41fdrTHnfVVXVjat4f2SjMzyXysYxZCulI+fV/0UMN2O3FmGPjR00hrWTbump
9v+I3bDuN/wpOH7zH9UJi8Cg/V5n9lH7rIHd+jX8txnsY9sUEBCXhPNF89m0kEBmNO5Msfz7aft9
L17xU+x2lZhY1+j3+15UIxawXGoaoh25gIOUg5m9GWNPcRGpefMrxx3zBi6FreRIaGndXkz2G4Bo
d4+WiCLBhxdhFFOTQalzfhQiu06xral00T9TV7LMcDe69V9OgfwdHZAjGfCMi7qqqy2/2xYvzCom
A/DV8lYzhoyb6IDUZ4HwORGHc7LjlCZswsAetIyxs2x4gfEQ6OozINSv+RAWD6gVwFrUTUsvxsx0
m5zL/FBitbtXq8ScOJJLhQSjcQO+X0U1ZUH2fa/25DrdQjjmPNzPXS6CgEAkwS+Hj1uyQVjqAgy/
WFMpQ3KTPrQ8ZJBFEEmaSmxiOb+3KsuECdVQnTVoU04szLhRiklscevpYRDdJQ7dt3ShVlF9Wg/C
dkXDL9gONIP6gcrKWjV9CKlszHjFbfUs2RngyEVgSwAFlQhlUz3pIrSkfWda06JJM+2i7K37dg1U
l1H0bHpvH7JMZ6CiFbNEXqRJfOnb8pMghigYg0K1y2u+1oiroQT90sdJPAnWHInwIR63odK0lgHI
4fkXJ8j5ELckE2p9zUefq4Vw0FQRVdPEGFzlpOPBy4fkpXJ1xEJLd5VgCHT859hGd2Lkfd3Jps9f
oefc1V3Of824QkFOB8G1I70+ICmPMtCg9StnexoN9FU2+Bj3jbuC4uC7xkXlRlm4sSnrCYwb2OfJ
Mgy9KFtKmMcEafk31mYlihBoAiMhGirDo8XKTAJV72sO92tp2EI6uk/djKBxgDlbmfBoMmI2f8QH
xmzoNmTPKNlN5oFcv4RTGj97ZEq0wcSG7xgCYaz2McaRqNRjwZgjYjTUIf6/utBbtAZ3QdMF/z1O
1Ig8kbStzt88RExFam1e2BBbNfahKIuCn0es/972iWJR3LD1hAx0RBJZZs6m5VIE2KE8VHNkxlNJ
F1EK5dmjHniNqHJnEIAmcEYiBu8pjxenOWmISA3ClRfkr02c/tP9qo8ndYeN+zIq1c7JDIsApi9X
m2IPhZwwKeeILdkFYem3jbctQN313TCFtQ8Z/b1StX6pV88Bycd0j93ikRzUMiF6f8HbfZV/ow3C
65bQeQmTPHodEtqTjfDozX3serGRz4m5PLNUzxFhmu6EKGUQL5PRTgAKBecmfPZn6dcf07YQGI+y
Rf9gqUJM+RtD0RnRK0LKEAWX/oQipa4RUdjFpZqabr0nauGTKZizG8ILzC/WNM8pAnZwMdIJbMbs
vlF8SOsDmn/ch608uWmyaxvK5c/2LUiMy7+MfBGeA3g+hS5XEOj0CvWjJzqWAZi87DDRUCZSbUdj
QMtV7OZlOkqkj7EFQP3ibzWd78D4JrKXYVRU4UEdl+0EjMLorr3pIYBnco5nCGaKAE1Rlb9l8io1
gnvGmxV1Q6XZNAJbrdnzGQ358F1ldAth/UYaboggS3rmqjU4Kysbr7ZIJcosyIurCHRMjs0hOoRQ
xdJvyWrDXuO5h47cR8vfBYG5t9jFYBiAj0fNaQqZymxgUvWXxZ1kAtlgjXAqjiyITM0IgWxQ8N11
X1gKZcij3vSm/yipR3M3Rl7/ldh8QFjHzSPKEQzRdLB5qepPGn4YuCjmqSrizbRa4t/q+/NDR8HH
Y4b5LC9NsSM5jdX6/oafugk8FCCLPHZ63fvUGuwzOqcDg5anDHvHbEOswUi5whMe9HXC9pnqYiw7
4018wfWTrPXZwlNfZEsJOCKxcWmF2zm8EWVB1pZVEpc1u46W/wlYx0IiAGuSmELcAN8jVX90Q9/E
W7WzdX+LDm02YZVttPvo4e7eSe0lYplmuXDyPGT5QyugCQlWi/rCtVa8pm5e9w3jExHC2e1BA4zB
mo2O6haR1PNPoyzP2zKHxqCzS0nKIc1/BnSY4n8jaoxH+uC9eFgygmnnvQuBmBYhC6ccFwLnd56u
NzcCMt+2DHMmVKHWVmQcvK6BEDWKrlf/J8+nTt58PPtahnBuPLL1+2yzPE16Qigi5N4eKsEbIQxq
GUy0qgDOp8qOZigztvPNsu6a17ecCe1btdzD6gbvNXSciXmclD3a0ykJA7e+ZYRMb3b1RutUjKL0
Vms8R6KpzWlD4D6VjlsBRyP8e+ra0rODxN/A33qKzkC+5ev6lwKarLYLLiURypDh8D5cegs8Louh
jHKBEC/ywik1Unp3/QCn5F+8le1LgQ9aET5hHkLx1oycY3tw9FtCrunhssg8Kba+aLRyLtDFOMTQ
fe9lGhUM2w+0wqO9o6ZyJFAl28OJyeP8vvhn4o3jztv5dLUalGnynZYq19IG0dI4+f5OLZI/NRGE
JP/PukuUtB9CffN4Th0x0uAv6Ih0dVF809+ABZ0/ptD7AdYaez5ORpU5eh+aeFNCZu3PJacBHkNV
VBqFz6yTfqbXKjJwlXAw1DTJj5FJOwIQqd4ZnrIGB4OdrGnN3VEvuY0OK9egMZtzXMG12uFsqys7
KS+yfkg9nvYrnSzS2b80n9hj1NDeAbwRYimi63lqgorBN/ecTC/fsTUrxJeV/Vaxvl7P3nIIMYul
UkWYo5lLiShVIlhmE3EUEvONjaK2Iry/R8xsufZifQlmXXIUVmUppPwnOfVAJ12kcn0+unaytM0X
wPZsAl6MA/osWilBKRXA1K+5sAMIs4nhdimvf7VoJ8mYbsaWykIhStOVeQwGTdE0nXfoROyhY/Ex
Mu12tCkuYFFl0xFwvbyPBoudESbuc8WNl+hQb+qWtYHTZ6KLukSf+DISpN1Pb29lOAlAQhx41/JQ
hTTdSrXcnJR8s2Bdh/k3a+jAem8M3misrZb9m1UZC5ZnduObpKCAu3+sVcRA+o13d7OCU9Zmnf14
ZlRJN/u65C3QdenAb/9kmR1gHL0ZVVuBIDPDP4TEgZS4vATjhacRLoGE3SGxnNamw+0uTPo/FVeS
F6QhTEBUD3Fm671+3m7RTWHEELusAmADewzGcNf8L3Tdj3mA+vZTmmPRuVAML2gOp+y+KHF4TdYX
XgxAZC63o3r5S2I8dzlLomrJh4Z1rB/hfYtLog75iEt6opoV5OvcPyFaKqoVQ849NVTrFhxNstFy
dF+Hw1EFwy4uTzzNXvEhXhnCfbjm1ifMQKsx1b6FlXDLAUBaXDy61b+homZ5mehRA3V5NF5IfM5/
T078GKZzYqpkvtORw0cgB5ClcRlYbm9//eg25X/3ivRMmrJ7fq1/6bdmmU4Y2cE19DqiAiITGt+l
xPy6BRv/4FRHXn7hj/F+wn5I8m06Rxs2pAbX8WzRGhZp79dvxCVvtAAv9TQzI7N0ufJRroWQnJh9
87ihi5iw9ANa18FUow+vkr+iSmQ9+Ihzb6GQ4rnZbDWfNm1EBTw16MKb+H6YUxuRCbIJhwcRm8Is
79ZqsgrkdJ07ko4ceQQ4NOs+hdHL3LrFfagwyrBUC7B4E62qhw2kn2Bg7u8dFphJEaLKoW22tJmX
hdFeExgapZ4Ihjsuu1xUY6+oDcNccPLq39+WuN9uLB2B2GYqJ38b7NfFZ8A2CxbQyCkBhh8jG1cP
2kDpp2zb1OV669ejNPIulkIyixa5oCmUPrD3fr5+fXEo6KcQfl005N2jrSd4NuJH4RpNLcRt/rgu
/hRv7ZAz0WPFnGD0sedffHyNE+OEKYBhpd0lx+3hmjQFAAEXzD9BCest4YGBdTbQg4pQaCntpt7M
+0o7K1A3DiaNvgTBl4D1Nu6M80M8ytatoHgeXuVw4RknD4Ai/TCjYxZt1YP5vRq/ySeYWVDc7YtU
FeDIYIGppuig3OQEe08urtp21WCkW3xUzN+YXJ/53UnXSqvrguyMbjPDykdX3UFDVCjy8yIR07H8
Jl3hst5TPM/hMnCDiUqhpDUVNF4jgaRy9cSWkoWAfNmGAlHiJJYUZvKrszfY98criIzV0LU0RvEU
T7cUqi0dK0LD9rW4f4CQaP2NnIG6Jx4mlA7IiX9Pf0G+B8hfmePjij5hXw5XJMsmu93nA8NUvnK9
a4zJK2Txyf2DHLz+8CONM/GUu6BNYsJ+Wjb8xnhRLuYbC0prpbHrklTxKZ6i2QwKn2acAwRk8Z88
T/5QdLmIG0C/SJMIAbKS2GBJvpJOTK54WXakI1IDND4pWXLvco7Jp6I2loGcPhOGbfptXQBfShxe
sp2YLzAIqKJrwag2t/EYJSuA2BfxNYhssPEt65p1hAmj2e26ngulGzyQ7Q3k+rdhbsxP/ZfSDmmN
VFByYS+JAAVtI/fHVPMUcZUfZw6/gYKIkJtuLHmWYOSozLwcQExvfIgq91DMjx+DdWgKPCatfl+L
Si/1xNAbVNTgmmbQ6qIXDPN8e+RNn7ehHtsuBw9tX9WA385pf1I1JScGRuyTYQFeQ731WjkxjXLo
sEmXPFF2QpN4mYCYStQ7Idd+SU8qQxHB8hqq6Vuh2Bf32DyOpkn9KPicjx8jYtJRMvTdhj8GsuTY
Q+pbFmM6nWrSmgp2afy4L0+CVR5ZR57MOLdoA/kzzTr8/hZkM2jo4VuIWNAjBTfT8w623Xbcv6nM
fTtvni9pyeB3gaul0HUZfqaO5UZ60rOKsQQtWAWggfdxyFpcbBScek+T4Umsl+ELszQvzCRc//BC
rdUirnQofwknmpP8U7v1IxnD6WKJ2farRvOe45c51GO4JzpbNYMeNK4hK44q4fG8wyrosgbmakXZ
eaq8n2M82E/dgeq01eZ8dXGP2WfaTorpwDaCT4DjinjOFid5MToCST1497YHihgRjJpiz1NpjFy3
Hl9rJyMkKfTqyWgq0iR2G6T2sdJens8RTjLTk55DMVgOdyIhX4gAiLbsOpupGFKW/RKeKzvE9kQ/
NCLRUTjdKm3EIkZSPpM+tLTA0MnkCwm6NDRUZrD9nD6qd5nUGUskf7yo4htlmWLKndZjCrIHqRH1
o7zYZGK5fHEnZRuM6t07K7jM1kGfz6DZg3zGzIA1neyQluEm3kcdrtuKOZM3xJ55QqeuZksOgO9k
7wlIt2sIAELy0rYns4gfckFM065HaiF6aN/OylggGrbsGPXVKl3Gpd8ZucBMT7QzyMwXT6SWvzub
+r2cE5w1hCGXjN/awYcwQUYoep+Y7peCLs+ZSTfSZktc607OG0hAo6QMO1feHmiGBvPI5BOa+GPt
3ag6MHHoIFIhaA/g5o82ZYv2gxz5iGKOWE8mh/Fpt//Mp3727wbZzVABHi26a6BHiAfG4hcUTVYf
tCUDVgm38q7d5idQumPrtJ78+p1ZyS4LMtG28fdTnO+hx3zIw9cIsWLYkmxJOouXfvA+8ZmsKa6y
PSC8VAFKn422NaZCZO6AvntOjhD0rk51X7VatujR94j0remkF4+SlgyAcrDZ/HRU3OzG3gOxQkMs
fsXig7XQVr6MfHX4aAhPQ3sDZ6Rmkq+1ak+1iFKCcShv5Bm0t3y6fTICnABvrcbtY/9fL+GoXUf+
8W7HV+RKcNP4s5xqlbJGvCA+EwR4sl2kEdzah/YV+Ru/6ZnfzYUbpdrtOivoZEEQxCjUoVT5PSfz
/cirZorbtrP6aE4esbJM08dzX4HmtRRhUcyHSV1U861daiB8LqG5n6X8+RD7kpl/eIrC6DWHtc4m
meJBBiNCZy8sVJkNGh05yXWsZi534m7CDTYFV2anI5Gw0KtW0ZHLIswGX//UbN3R1FfiF7HO6Hz1
Wl4f5GoPd6qQi78D1e5f6OnvOmsD/Mdn4anxyRFJp8PNWjrmX2IgTwLUgtah3Msw5bZsWCRgpV4C
rzmC9zO4i+k/Alio+jW+m4e6rbfxbrSsLLVYrpcfe+lttQmqVOVDuqCtn7JRJ0nCYwQB6eG7WC6k
Ym3J7XAEKz6K5NVRDk0zEXLhVgsM2PBlarYcZOYivV6eQhT7zm60NXyxIbVqOCyjVxDAz/8hzzIa
2t19eLd43alxwhxu093K89cScCVVBx8NDcoWO1yzj8PfWLV3LqjJ4cxtgZZRpAB9qpDunkDkirNN
AMVy3K4tRVHYjasulHTkew07X7z2UHCNoRQlVeTTNU3rI5ood9HHdIPxJM0QWukTScQLtD0DAyvH
8zD76DAXENwr5jPOfgiwSp6cmDXMCLO6rFn89jEBOZw21PXVzHzjiZa4GXGqakF2q6tV5tR4iF9X
fvhyniFHrqWEXw3ZbWeCIe/IC3qHHJWJi1NfgdbIGexHPYGEJrewAhuOnZ1D3BEcNnO1EppJNLEG
1PMzFd7z+ZLUH2iLLA/LxSsJNSbuDVGBeXkOnFVtxSP/JidwNp6DjJTWo2Q6ZdxO6yQ9v1iQqZEY
7cU/v4CDtUXzpMNZBjX3y0WpXmBvcoGZwjsMlpCFY2SCRcxLPApRg4bAyIv9XmzG2yVb8G+TRCs8
X9Ene0aq9UO3A1Tkhb/aeIISMy6Wk94wR+yDHpPVmnolomFpIRX6kNWtzd1AfeE3I6ywrn+wIDie
pdgNMleh1bdN/kiJygsk9AfFNkxewjIySy8AQ529xO5OiSG5f9906ScnsdjIlqk3qEsDMaE14wD1
BccdU0uIxTHCJ4d75n8Q2o6XMbV9nNNbtfqDyRChYMrBNA23wAs3XbmjF5mkJGRGhBOQo+FJQWYe
DD/MN6BqJLz1iiysPMuNspbaef4Sc8N0LMjG5QOnb7HCKA6xuuIcwr7RW7Rcbe0xLZpqyTch4K5L
3oWRjQondmojjNAmC/9AE4fxg1zS+SvA8zHLOY7b8pp4sOXkMnSunJx4WYHq0rfiWsekC3WpYOSt
LWxbYNW6V3Onw/8a2i+TX6WeuweV/rAZe0PHD9JO03tu8emshR4LBoGmJrHZyisqiefgEFkdc2Ty
kp/rYeTbqSGbLYZzItgAkMOlN/fPfu0hfYhuiqpQZgW/aYPJwY5gyiprfYmb1PwQnoCZ5+6ux3kE
lbn3fZBzThOK48JbEMPX28eCbH7nh9sVppzCxu8vGmTuDlTfF29jfsIYCStIl4ujqJMJM+nfunrg
uC0BHB51WV24K8o5w+8WHc3a6BA8KGZQ/ipaJJvSTw+1IoeorYit3LKdju/JSg5/WDcXGBwMsRa7
TIOUfxkp4NQCLh20oEcJ/1dHNAxxoBW0HtDjLZpORG6XO1S7/aWY2JEfdAj5S6PMDc3GC73jYsOi
iidPwd7zfJzw0KL8jJb9eCkyAjcKzb78J7+8tI6mm/aozoLVIO3IQ8KDOcp0ZLO5TNZQUEK5bY6Q
QZrXryiaqXgkgM0ZH8a2lf46jyEL/Mu0YkB5CE4ZtQd9sQUN0BCGUYhjTW8VYvBvwJ6D83CEHVM7
vPJ0Tj2hcXQ2+w1FYwcHfeq+6VQ0s6jjY+IIi2dqEX1+RLYTq7B/pYBlJU8hstCF6wGTUV10PU2E
kzjfGSXzgsCJI+TGDl6z7fTh677xYA9WEs2s9hVoNvGYp7PmyTjisCbl3lYh9OY1BbkckUK5pVAo
T+Tv9NUUq1zHjIbTE2mznhScgGwNdsY5OnyVSiz+gI56NNyU0t6rf3fkFD9rKyZU4IVrPh5f5hug
SbF15qZE8ax7DsGCyQ5YC+QFWWnHFnLD5fu0cAJa+mWC6SJHPJMv2hYEBS6gwj4SLcXZ7l7r/zVu
GP2Y+n6FuEPJ8fFwOJ16aoJYLqL1MxXBaS8TsMG/CAplJJNZYoci1Ntf2wCWtVEPCj6OhQZsveAP
SsFgc4dK9IZsOchn1/U8zIOSQ0Tu1IsUdRATqsfP/hucYceFT8lU6KfaPAjNh+Zk8MYfMt4FJJif
QRHJWSn3nB4NH98gM8fUO8GSvGLCYW1h4hyHA4cGs3ir0hMmJ4hBMajc97nz11+mW3swuAFfalVu
KkUvE15RWypMrnIlvaCPUN78WgVNNT7OGWCa0NDtHIYXtjFuAFzw1f2soLylcsuoED6LqG4tqtm3
NNdfXyvX4qkqkKZVPYyprkAAzrA1gpitH9i4i8FZa40um4NW8ZRU3HbyweewkeX6AtLCS3Me98c2
gFBaAWKsNaDGwgC2+BWj/hcIcta5D01dBTQkwKWGcZsBMPGh2T+LLjuiXNbYKImmMZ0vb+etHuP8
RQ9l6gjlhmlEDqm0elSaHhrgKxWM0Q9yhHFQiKACAtTZIMHXtpFxrS4O26uOWOpsYz7+vBsXLkE+
dI7dO/YRGdEWujKKlxo+n16FUKXBKSBsxQ84qdQEOFYx+kDfDjihycPmxNed5cpuX63FQHFklu7X
BRBAvb7kzLRbWkqjdX94siZTLgAdc3cnM4Jftj4ACfPcOVhRfB3cXWFO39dj0evlKUx0UOYdQv1N
TX2pDmSsEhlZg7bBKOoEvgx86Ys5pxSB9DCY9aI888GPZfIRVOkLGvp4iEL5RTTh91PD5DtN5Ncp
n30h6THYRrCwzjqLdjILM1bTy3EXjnzvTWEaHb22RIyKQ6KTfzxlA2e/N3EoryRmSe/W9YY5x4fN
7BALpDlYjEo2iRs+DDWpViNle08+vH2DfdoWZI9H6czk+ku7ej/RJwI/U/JNOrUwj/u9Sw3Xo7QZ
mNJvg6Qo+cPQ+zR2F17+pvCWPkZSNmLkz8OW722r5jSgrL9XfK6NBt44RN1HmTuzRaoDg3r9DFZZ
w58CUGcTLywMjRsSvGqyivYPSi/uMFRoZ8XQxeRZ1u0fsvKMdbRx+pbqDQWHgJD5vMtSc8sMc9Fz
mP9W1mwXGwyJqL71co48ags7q/aH94pUAxW3DvzIyW6B57AzUsJllFjUEax6g5VJ94BlbIsOWtxf
+FHpgbo4mPWiUF0uEUDJPshHq3ZGMOdnCOB5+cCwCXxtXoeBSImZOTqx/8PLI2IN7nwq53KW0z4A
kr03j/8fL5ov96UzcQju1yiHAZTHKGnZqQduKjF+OVXb6UB5VI9V4JQ8oKjrsA/M9qwGH22Bkxod
Qxyi5afwWm7R33pRij8LlAxXEDpedwyg3wQUXCV8pMGectg+JFTQgDn6fXwf/pS3RuLFt9XhrLfq
9ifAezOd8xjkiNVI9ZPpErFYpTkhwsZ+0fw7sHDWtYzg7xJ+OiMlAF15SWcS9DGBXBsfzhTCzRKk
O9Z4NUdL+PslkQiSjdnF4MY+1dmvvm1vXvb6MV9HcLdStg0ZjdyV5RuNBNSKTLnXMitrWDTZrO5J
eNg6LiRsEUt0evi+EIL85YYTOxqInAoV/60R0e3oVjAnyVbThIgurYej42YVj6c4SqM4W7w2/0Il
Z1PkLd8S8D7y+/UBfUKUTme1WmFxmonottGv9GvQ5HtkqZniDAp9Zntd6A8uHsaACwYxo6JwDj/2
CJAwVjU9jU9M7sgLsaCR2WskY5T1rR5BLkJbTQk1dnRjFExyB9WKxYIWU4cR6l6yQ4cKJQAhOCTX
ipOpTsxo6qayJb0g6l50sDuUVnFr6raltOZx6YTbouz1I47g1kGO+DTuTPwiLzKRXiYljeoJI33y
H/SrR8TENwAYYnsm8hpSNW4oEJf1F+Jt4VeX9eyxo+0UJUni5TZz4BkIiEdH2+nsI0em1XqHGF+2
XKzfdHHskeM8AMHgVSAlFLmZ1oasoJCOd0TsKzU+hyyGaXlVWZYWlYxznnI5SrJOhbsJ376KAn47
IbF4cnmM0Nvg/XmuqLcaPhiaCbAPJ4wTeajPcPnGqitEBmi+iEPznA80NhyDbRhQgmp6fYfKBgR0
BG6BECv5CZpIPRtOw0B7dHW2OU3NgzTgcQb9yQn7Ycr3Hde/Vz174dK5p2OwVkhdTZfpc20NPpxW
NWBaVfcF0kyRG5Gu/CQ+kbXFaa7ZxFFp3LkgvV3Ny76NOkfOn/PwW3qYofAR0iUWMHcYZ4eKG4mm
sSzV0sRqpTlO+sIaXxhCTrBtta+WMlDe2VgeuuXAIvD+c9oS7TFuyGw6MyRtMVH7m2TNWuMmsbKI
X3VFCranYJzptJUCp0ysgvbXBWzUGd8CWbhV6IugFhGUfEKJEL8KsSlyhm/GC6KrxaHEmrGIi487
n6Hu7q3pLgDOy1W8f5tBUaejHQTDrRZfoGNLIqTeO08O3dCKGvbZI35E7nIgvF7/064yXUdIgKiw
z9lt0KUzbtzgjySsMlLM+3JnqUJzSSamj6hh9cL+TfGS/J6Ljdg089vfNt6ouZPMr0dLmCGYRsL1
Y6+Ylp+eBa2upjXFXhGUydfxsd4TnbsVXomTmJfpY3DW7biU9/c1p4YXcJQnKfsrO8L7uHtMQsDl
4jnyekaA6EJP2T6n1SjhfhFs/aUecigSjY7t3wmOGvCATO/B2LkxETEz2mtX/nMahx6FJBgxEVwG
snoHaG2nbMSFYqE4SbbO5417bTse4cppkuV/af26ib97UoSddhc3VIG3apewckvTUj9rRw7hgtpa
VNLdtdh5uRfB3jP9xpgUF6baobacLqewMKo3Hvv7eM5H/w27p3SkvEcDJi/moaxkMc55RU6vecLo
P9/4ScS5WwrcsZeJKpV4I8gk8/a/jDfQ8lrQ3cTopspNzfOny/826BAFntBj2HcgUOhT8AmtQDQd
jC8NyFSQE2IzXRMz9e6unNJ+Fc+GneEgRUOgzZL6+jzSUM9USkRdtMrJn3iebDDrJQmhMx6MDyzg
zgi7ftfoGp9Rf4eI5Zb85f4o1GJmLHoDVmBsiotR9z0x2CqCnOAp5YU/mJS7G5i0m01oObnl/3IJ
hOzml/rmqMOA9wI3kr26bqA31PfCb2svJhwRjQIXZfRnJNuFJl0H5HODvA6Kr4HAUupI6sDloCq5
xw+eURLpPFgA3Lv5DcSOXpnaJfK5RjWJjUqQc9BC5nkdwiidw6zjkpE7TE74R84p2NyEYJBNqNnO
FZ/PNDCl+oCesFUbaIWpn3fb/yBuEtrpaxw45JGYwz77CnXhraxqb6yavkAL7S9JgWDuhFQ+t5A5
r4IbO+Y31bzJ2/1yfO4v3/e0JEIKwQ10DLOdgBmdWqqU+RhtLbLdhySRXAVNSXsUwpye0H64Kl+w
KTOM2ngF4RsV4gqGDqNjpfI8Wfa8VGSi3lYuNAm3VZLSKv4K7c5/AI1/MaaNtaSxTrgPRXu+fTT2
Vbm2EoaHo1xeK8C5iQGyn4F5X+L5Pqi8N5b8FBlF3LAO4vkFjL6MMFwNZLGMNF1YvGsIRuYdB94v
8odUw/9bAIGa57nD+n3ExDP+G2Gm5hmkp5cvF0WK3WMkCE8vTottGxZV4NWeFfjAskZpW4zLgndz
23BJqA/f452aBF2a3lpK9g24KSlukqE1736yY7VOELfjAkd9qWocCv1lINAh7ZSAFcJ9oq1MK20G
ORPygPh4HpL95suHODp2zt18+LwYS7cGI1qOw6aOw7vu7VQ9yd+WpYW4cF9thrwjWUfnd+NpYom3
EmsgA5/A7DzVcCnd8zFPVS28t/SWzMg/FKn5HhqfJLVYlLEI8gTOSBVzlrCxdmP73mPyd7+hH05O
UR86RHujgStt/GdWltr9c9sCvEG4144ke64CnHGdZn/J78XLUZvJ9O3wOGLrzGNgQoAk01QLMgDU
KloE1dvtwjPnXnmph/P7jfU0Rsc/ltnpITZat7fImYRt25zH+HDF8PYj1YoNgOqFkqtPx3CFBnV0
ZkejtHoCbiSGS07sUAOfElP+RuUKGsZIu24bXIXoJ1CK14Zkwq08XpwwGNkeVKR/Z/HyQS4CUiRM
pf7jpM9xxptCF58bwBCTYbtXSEL6Nwfus16cKpK3hznRRuDlU01l+mK8Y+JaBtDzn6cmuLkTh4SI
f1bTMyeHWoBRcojGvARp4WAboCeg27ivYOMZeca4Ga5rselOEKYLKENiwqiY2PxNKCn3w4Hwjbkl
DwnyxC0ZXjR/nn+u5xAJhek8vANaS/G55cl5DnGrFxQILJvpI9t4lQcP9D2LG4y7rcUB1DEkrujr
KhBZZoWy3zpYI4FsMEmE4TIrecBQdTwT43alP7beshkG4OT68TZD2QBTTBhONMs/+Y6P5mJ5SCRu
Eq3nAlUYbgCIRZ9k/zpoBK9Mz1d1P80ASZqKmE0Y2aQbSYdyNh0Yj2UwwG9/aZr7crTcW5bJouv/
TGwWYgZzm7KFKpDC4fH+NoMgXnKwU0brBUqk06ZFC+a8HBCQiDofpUDGJK/cG9xqV/50NHrviuVs
cqD/X14P3lgdllX/gxBtn6OT5uiFhNOovUlgF6NwpfWmDpqHIi6Eofv6/XL65YQ9bvSS/XCJ6jL/
0jYgbGNKqE581tn/RH/3RJI/S2q8Fqcg3UnRch9ti4O1oQsr8lfdWlosFIy1jruLP2+w+9R2dGZ1
2FbFCG51LjortoYzsudE9R6QaVNrbo9sZYZJ8TSocIUVuzVTChfaoc9AZEOkgeT2PGNc9Obgc4n1
HrHFRCvHG3yAsopfrfVuYnn8a5OFA5PtrnLs+e82deskGHr9FCc7gbVKRt6XxKwHDGe0HaS0VXYF
+SPFVI7AweL60kGeNUK4uBps9t/MGaXoB9L21xTwCjySmH/QR9ugwHjtAPj4zmJiJKoRii0ZKjU5
hr7imhdePH7HZSFciU5Z5F8llTEpZJfov7jc3Ed1Q9hkzOgdG3aK8x+mVhZkwqGnwIGEPGgcOzPG
Pf0oEsf9KqA3qoTZVaXSOkGrQ17jByTaJZYD8au4O1AKcIi/HR6PLGQwOxzRrQWbR0HJvETDriPH
idRy0Dz4z0AISHYe/2TZuSdwwiRbvj7K/hOghoG/kKKPadxe7boXMHMLSJyOH3rz/yfsgxaauZHS
vJujrH9ZtbLktLAZcNcJPHuYFctlKedGCwmUxUA/y8EONSh0Jff8GTaTSX0hGd8Q1hX0y0ZmbaAU
tC64qLdWLSp6aQqebebFtpDlwW67EgrJUllLNsESFcoEHDJqOD6SXvSAGrSHhAKTirkDdKNA4EUN
45Brn6sf+T0MGDEZXjfx6lla+qrfhun2yPammttAC5pR5/L/WW/75EngV0GRnMgDjM05ElDQPn8G
LtCYQd3izxG0K/OoO/ZzVKdRyQEOrjzQWnZ9XdOJmolaeTGimZ2DGCCymHgWEdUyMUE5LQF9XLce
8oLntVwNqmUy4K9Ni7vVqzRbhr5CWaADFSA+NQSxLp0r0fC7xDSlJ36Eg0yMPAeMvuX9N9BJfGxs
ejjzm/PJYTxPoR274+r2gOhAN4I3BVF6UAGqcHe+KLOVz2J+vkKIp1+NZ2v5KsHuNC7Vx6F4IExi
uffBIY197gVaWboD+xtW4Hm8TsglJeDKtlg0YqijX/DeBk2uS4hORtrMMAUntKCOpA3Ag87XNy0K
owtugirjehegkg20eRNP12OVRSAUseIJv75d6lkjxmLXJtiED2X5pCPRt1YmYzdsjD1RzSD8C50w
v62AWA14hD7do3dasz+r+y6M+YVmrBG44pqMwrIVpPn/F4rUbkEzf3+qf/uMuPBELtLIOJTJpnzq
6QBmxiHkH9rbqA+UZCQ5h3on5zsMX9xsqvI+vzR0EP6LA89EOe5hhje/j1Y4777I9dsDB4wJf9NZ
2STLBHZspnS/S+iv0xeuKmPrNthHU09xpBEbbfvPBWpm8IKFnfTcP+uoqhAMzLy3gTBYKRURGb1B
sQWyapuxT1XnaYq9vhpE75mzDtTwcr9RzMBig2BRTyv+Jy3IE9sma2wQl8ffXLDWG4p4BsE6VPQC
LU7j6AxjpdpRju7sEybJ+7/DtU+0jMPOQFB8rVz066zboXRErPDCpdsZqRQPOQCNJGjR1c+BgZ73
tz1I5uTtykQU7Y3ORa1xoNgOnC6xfxcM981VaDQwZPUVL9cv8rX+0sEz5aZWhERWX/lpF6dRHHX5
9ISNdt4LsohMM84V57b+8xe8C1ci9+XKpoYEwY4CUZr8uPnnHj1cgdMtOPNnqRf3mxuLJ8Q8XezR
REdItmet1sy5cvg0+1ed2poGU6V4Q1auptNjqbKMRtw0+GFKEuPm12QlzC7FmMEqnV/WryQgKfgB
MnZEpKrqhMJs/bpAfYFycFPuMJYTtYpAuzTW17KeHJFl8hn0gfEsytYJnwoMnruQ/8XZgab4g/jV
e+9N00tkf6O9OKeCNJawncFQrrn+ufl7uYVuyM6KA6H0R+hn8MeP5oWANG4Y+hljYQVnoZqUEtjN
izRb3ReRT4HzWGwVULMvC7sqhoK1aQvJACFgrzH5smMXSq4iDrE+cB3Z2k3c5YD7qmZaDfNNpL+d
XwOMu+Yym7xrtqj2GMuteIwCP5Ksc9cUJ//SK6rK/70JbIEl5rcTqK6pI5ed34zNimIRsYrUMK9p
8OU/aVPXKUOX7k5zqkZSMSuZ0o7U63+a/c4Icx7Tpn2jDG5v55ZCsNw2l03cZCs4RKGADXKYI+2a
5DbOP9mDFxS7MkSBOBk1QZRX6pNff8nucTY6uTChtgsfpfQq1jkYyAmTAPmh7En3edOhRaryrg/E
Ixaxf6pnotr0qSoEV9ZsgrqDBRPt9/1FbE/s66kYUmU77lr4rw4tVPR7Hq55fUYlB7tItmr4hR4a
vmbqW+F2sqXBdB4/I/jFO1WLzqyPehftUgIghuZ+FdmGflmcGIuF8McnECyKg0t8mZw9BqEG1ciP
M4s+ygGbRL3veHI1Crj0WZqjObCRuXhLo3KxdPsIvo/iSOwy9qSYXMCmECQ/j3gwjNV+3ad+HvTf
ogtVqu0ogwVQJrsSXn+HkWwsbBtDoIk/B/gBEAWclj8nhm5EUpWoUDzIEyk+vSW9lE9ycIy0UtVT
mZO3d689Nj0yQyeq9S3g6s2ilQSiQX5NbeYXDOUosfuDTgDh/Zb6sjzHq2Nyf+HVKad2kkRSLpE+
D1Ab/vi2GidNyFAbKG736t3g59RxZfTCoX2qOyh5Cx4NOI38P1g1rmVgrdODy6q1jQAmEAy6RuJ3
0q/JMXemqyAT5fVaiSDejp6Km09RbK4XWl1oDUlnVsIK9RYGldTe+tdQ7mFDfSs/J9oI/P2k5WRw
I4YJwdOFKRcosYVW0/DUvnGEZRqPkCcDGarB2xBLcbtWcZ8EPQs1PUVI1QGfooshHe4mlFKvZXOl
0xqGg2XOoSZHpcjAzlllAVw8TyM34xdLVbN6Dk9o/V6S+TFMitdxT5ta4lXk3rdZPQGTs9uTQpLu
f5oU5q/Ecg0XO+1dZSwKh0cdTKgg9T4AvkYpWk3qelt4ec2uN0FufPi0YITp8IjGiRAgmI3gL9xI
36avWYjR3evBTvHxlTcpGUpXhhzL8gLW0YA0iCZ42hUZ2c5aT1iq15CdZ1sFECnL9FO/OVkny83+
syCuPKLutSumP7/A3P/iCWfdK2xtthaz1o91YzNspwDhYlrnrmTVkxlndrPcgAY5lb/mD/CuN2Ts
CSQLxcA2nCukux9pwM8vrWjl6TRzuw9b5IMPzRZfzPRvLk2LkIpmC5cvjKGRBPlt3qFGLZkAJLTy
z9tb8f+XhXeLppY9mFLYm6pHFZFgrIsKZm+0QN0vFpNUA7PNB6lSqYpPP8IMY5jxv96buCNg+OyU
IdLT2OFqpNyQL0ceukCE2ErOgBKY05EBosjlfa263DR8usw/Iv7fscbnHj5dWdiR8CU+iZIwYhjU
5cGOG5+jt2PLt/yfKOFhwADYGQ6g0sWW1pUEhXrhsYys+5L7yEXornk0n0i2nHtvy5Ij5YFnpuEp
DWpQZseOZuk6h0GolsCcBiMMJ7y70dZbdaho9XQFa7FiH1CGawxt5fCP7BCtn6U4DIfbgyJQJ9JC
TFXoCvKg2X28LIHnLsQFASMsBpIZbjiKXsRXagyOjblXBUTEl0ouNQugtHpP35/k/H8P7mlqF1qJ
PhRAYUHIwKXfWutmRf0H5nwfBN5uX1fiyz2ibIVrLIwutjE/j9LHtUekUsJgJ9Ac4MQnhzLYXVtd
RVF0wnEsMQMCAeo6iEzDmO2xQFEbcIZKBNR6EdGVuTw+tXpfrxjF47p9chzu/vXZc3B41eyEIOAA
AZEDlvbttQZ60K0QDTEeLOIudlKyUqm+W84iiLZ2hEdg7xND1sIMbzgq4BhDjS6arccLh6Qe65jb
IcM9wZWFnAqpAhenoU47ZS/+h1yNaXydNwFC3J+jpd/oVosdlo+X5ghvneHuvsAM6MORDzahGqp4
Ldeq76dTSRSlf8HnrtzSSrGH0V72ZD0etb50llWyVzF4VYorBJ1CtsFbBReXQwkzAHHeh+RyzUBu
RgYVNzXGahPoKCSzjRskVzy7hq8kIRmEf1NqwtYb60rCOYN0wtrE1hMD3CsKZeVX5igPVhE0QfiP
oM1h+u66a/B1ub2Nn57x2Bfjsw0cETfKBVV4ikzolppz9hY1DElVTjZk2ecxLWmtNCg6LYo2DD22
DJd8E5Hv8CbcdC5sOWjOjJqWBJiw0hManxMfxrrb3t0P3LkmFBypzXtut4wCMdokQc+Y7BzWVr30
c7Q4AG46hXSAdZziSrqSo/qc/yf4xe91CqWpCmaZtwvFkfFaEwbg6hhdKG3Qwf03sPDk6yorKHNm
nWxkVlD9W4D6VBnyWlhVyO9f1FWh4RzySsrt2p5BWO/Hb3a+EoWaaYgTvLYSBae7wyGw27ebiw/n
PoJpdhWzJophPdNM1zKeONKeu2qPjRY8NGRd+A29mTmjfoHUmNpT2My65IVvEB30ysUyCFpgeAzy
eM1ZVx3rGFmW5BvLIvmhZYvHNHu+srlSa3eeLB/e7rhWj8n0zvn70QT3VGBln7DzRqOWIkftB0I0
geRqUwHAKFnMxuYqttAJxxjgcohyIghHZEU+xuAlx6y21FTLyz29In+20k0Y3WmbPcWiR4/0nELR
0vvNP48nOtH3zHcOsX/dGrI0hlJMyp9eYVE8nk3xTMlGsoUbfDNKPJjb1DZJO8p9+luVqdkQpdfl
6Hke6ajtm3pAPqCkxrYOd/92ZB6HGDD+UgRRMzwkJemcjwkgs+/FiojDqFHMxVXwwKDG8JEQ2bzg
stpA1Li31uxQpYAkhzvf66yjKKRy84MzhF48+IndObL0dv8MppKtIrNChV66q+SpgIH4fvOVTHTs
ivZOaSapyPQBiXzkb8S7Ny89DTM0AjEqs5XLnH6Gc7f5ztGQzhXbee4e1ekpdAYOsjdFfV/8FFuv
42glYikjWavhHGigTxyRV5W16Z2ZwbQcwWmT1W4YQxm4vti3L48EgyMi3rUQZqcW0+SoKvzK1JJB
bJj++ro6xOAbj5wh9//kOjQzgfz+HFMir+nxvsy+ywXX1GV0mVewqTZPuBmHjEEelaQ6IxyltFbW
MbX5psGKIiT4IAATeBdfw32X35QGDwjgSHDbTYgLguWNKAl/lAMFkzUDnEHB7K7qNwmma/J6O/PX
0xYd4T13r2+pbHqDg6/2L66huFyq++PNIbGMQ92OHJEFKyM1Ypo3HXOWy9ylzb9o1Cr/RXOULUrL
FhoQhcjmej4rnjfHNSmjWtvAsAPLsLPBKh23SGF/M8Amw7PxA+Gk20zj0Ed7OND4/BG9zsRPC9Xt
DMBNhxRyjT4ij8+4QzV6tqsJbFvnWrBoGZSkn3kPgvg659jWznoGd+D+59313tFvGA/GycYvFWl4
IlrEYBJVDUJwVPEjQWyE9ltS4WhOTKilUzc6/aWkvggmqvI05h5+3l0q3Ak7R0IgXcRNKspd9ZVc
cCrqr6r8HdkkalNSEPJqFTHL2GdZiI594ok6wJ3O/ZtH1d1TDFlrtIUUWRWxHc7CLsRTcmszVlcz
YELJF5IZA6oUQdYQbM1nqGvrZREI12ojZOAqQnS8jgWcYQdgGXB+scML2d1p/QNYGQdR7E8BYxbC
6FOmYSJlC64rc7pgTubs5qqF7tYOIKkXZazCCEz49TbsXCuJisr8SQVZkoZwra5s4GOG7Txrn/gB
6s9s0YX8Rr/OWoUHHbP2Sv/Uz0DBEyucvwgJhWmXpLvVvEodiLoxmumEY7UNc7lrMZk00XUOrVRG
0eeMojvceuBM95R0bwdVE7mJreNVBmOU7DHUZ2K6YwUoT9grJalibQwWNvgHN0eN7DaWzWKpXdTe
IrnGcuxDtrux2cBvvkuESrgg4be9AgU1RlB6ciGzciUFY9cwRMsZ3ksbUS9LXUWf2sSSdOrtnoSS
j+LMmxiKaEg9q7jjUItsEkOM6QI+ZR9Sfdl63qiJL3d9VNRDfT8EtTD4fRs995vnXuiyIW913TuF
xagfINteBunqg7r+QLN68NUC2FTkZAeudRx25HZhqPfLEn1JOsHdRTMtxkNm3KQFcIFeGBaL50fh
oAyGkXAGoJ18oPMmJF0GR/CjJw+HdeLvf5cD22TXRtPG1HzRIfvzca/Vw1wHQ0VdJIpF358Q+8tC
mCXrpnHV2Qd0Ayn17oYpoiRKAfR4PXogvfeQTIBOEoG+kWM0d2fnci7jOkbK9hlutxwM8cud+inW
URmIl2H1oKaXZQLLY4dgmWF4AVBjiooq/E7XPRhUJkeuX/MZPboDviyb6/05NfuZGwBkBmanjYVR
t20gawcP1U7f5LsxNBDBLqD4WHi4VlYR+rNp0SoTUrq/U4jzIY2p3ymxy5TmHuIiXbUPvNSbdZe3
lcY8cM4feBfT8cYC/Cw2IfIx71f9Aa+2SCBYzeXtBs5ljRx71rt3MulCl/9mLHlMD7HqX6oadmYH
2qy2fgLAkQGk0lwx82MF95nbkwGMqgVD5mRvdFs5yP4Rj0GJJjGcecLk5g+Qc8kDUDInBlcHQWbj
2T1LKyrpnu8VA8y6Km9aH+mOM0ehWepePQFmV7IYekx65UVJfJTTTAIzT+ASjHMGvTNydrOp3Xp5
xRAYa1k06muX+laUoRUFTRf+4AJwxyXYjBCuD0nHQISPFRkfTlvPIjPf/Cdj55Pb4srJjRL6PbUd
d2IRVq/QMPOlf5mOUQ+S9X1x74W5ViDkFOggjOSaAGxi8yYHPEfZ5Ux5O6dnIez4USvOu3TOFhsm
O5pp9qmr3p05rJzOauEFUxBGa9jrDX8Lf8Ts7DweVErGEMYfNo/JnRN/pNan2nFMEHnDfqpHBgV5
UpIe3NLONIZC5letBp/fvW0UMKQeCelWUWvp+TVPIfeliplxW/XnwWhWzDkTnrFW5liDZQ6fWkip
+C5H/cnF4HaS1VJBsbWDPNyxHyOZ2+bX3zQp3I1z+MeIXoZbSlp7bEJEAyi5Kr7gs76VIm6bo4WF
AiVcvU985LDudzCHvUFh1yarUgNNAwwT76jqM1Ovqvb1az6S/fuaowIqFEA1+1e7PjJhcUA3LGuV
hZ2eFwpyobsBEbKOcjy4/QU4D8w/1dY8Cwe8SiciBC86P231gD5Rm7IbQjpeihy6mG2nRsMcsK/o
9q5g40Ny4NrOpXa3XLXWivfXcOTQXVVKLBh2SRBA3oUi2xKD6kvwQvGiWSgUmEGVgvQ50IHoO0lg
eF58QJ0SyPGjz6olEgO9SEO2LRF47pA2gMQBjO2k3LBdMLLY/oFDNgz32EXthFicoC8Y3MfuWjf9
xYCwNctWOQbBUnI3JuqOFNx+qG1RM2VP1rTio9+1mxGHzmR2e9hE/xGW2f+6xAb5RMZ8n6dIplBt
ZKWn+l09GiXPgsLuGLFpnAomcoH4ptMPeDI9h7lKnlWgpy59rhsGgKD0sk/GkwmZ8B/Kl+oa0xPx
pqbKk4/ZEQogwF3fknKdadUP9fVqLf3ZPDQqJ5gOkDvTFroy2FQFPYu8Pu47QtoUyCmn0cn3OkrE
JSTe57owzW9PGMR3FJZWX+PS17odvmhZBQ9xcyPDsAIPSMw1qxr1yh5NpSEzlILt9lqWLKtaq7Ka
xyjV2z0gvsXxdEuq9SxOi93qvl4KBWPhjz5275+Smw4mAeUlGSwSv57hzU9ESigevZb6QLcwWB3k
OKunBZ0dO7FzrwJsMnahJ99sD4JS76hFcSTGcJsFmLQp9UWUlx7KYZebS0F8Xzf/QH6LNZ/np669
fAntXVqXOo/+35MJQ/hBSAHWoNZDSGAAlsaQZStrd+5LuRBqL3hpWrSVqDapWzHPW1iTZtHJXNML
oB6IfLBFdf7freglAQzDDscvnwDXx4yoJx6BWbKKbMGcJFGmEQyNTCUsCysRthRJ7nnvTLAVRGsN
K7dZjAgYDIBzTXHcwT05O8OxhehgDZ8bo7g01eJsZXGYnXgw2IDwTIrJOSZNMtLfS/puc3SsVV0m
V9aH1QBXWdX2buSzRNC/63rCR62TInYBirkVgA0aJFQmS0xs0OQoBhm0uXui59IIqe42T42kq+RU
Z1QcN/9d0EPe5Y0KelhNme4U1BTydi6xBE0dhyIwZkqUsXNh4j39SPPtehBDquX1YKN2dLsrRE1Z
RQyxUR8AWtPMFLQ1hZugd9qSh+trLjiB/BW6FwNRvLIDYBUAbykIsXG0BNNIlrM2X63k/s5xC8s6
d00bwevC51I0kgD5qAXnmNjS41l9KxnTMVEJndFW+jf70OXU2x7E7M7ag8LGaMBOcMpTtK6bRoX7
8gSrndwH3CQeD4oUopY2yXJVk1yOTY1u9lz8q1850CxLckczn2FpIWtU74ldL90I9ZsoZ6KlSSZS
qnmPxxPl1f1qBcDPeTCIX+vbICEnMD6XLgsNLMVZCjrYcHPpf260FzWCFTLk364T9i+yhGQhKZbx
OvPsnDnKJ8xZqez9sV9knxGD5APELc0PPr8iUA+CkNNC5/SHWl8uINVzJpFDHl2qeYZF9cvY1D6t
o1kG5iELKtwJ3nhUnkSYqCtcsBv4dtnwvKyfmzTSPUHoXiXaqAlZvbp0cCevL8FvCxawoFT6nv+u
5a4qjG0NVQYHkMepUKbk+xio0nIksjzKs1629cXQMs4qr7RCDv+TNQnL8/iQP4g5IPl8uaqYmT3M
JHZyuxnJSyLDKDVNB2iE4RPElU0gC6AZlYjVfSdAKlzu6ftUWkl+ZTlLs+Lzz+rPf9BcSSlumg6d
rgajLXZstjOFOAr3hoZcJKV6mdRVnsLyFGr2tEPtPSkvmiXqsoVEMXPoqictMdDSkV4MZi2enipm
3xRApOYZO8YRK0hGlF/XAA8H/T6+sCkhWbQ/rL4pVx92oFNb0T5OemKShEzxeUjDRcyzJLCG3hMW
YM0UMaLHx+kOlL8jrd8og5+n3D1ZGND8/8zDxMK3DaDbYxWmJBh8CpGfEzKvh4TrY9kfxaQNMHN/
JXQKiJ8JXCCcGdw9bNZdJgGnc9nflaSINZVhcKwvmL0lV7M+q99YzCgFsCfuIfneHa6g0yE/llbQ
KH8MCD0NN9CTRiu8k7fK8sr+WUNGkJfTvOTLT5mua7BARBMtlE/XVHX+HLxDP+MLTSGJ4pqaz1vI
PaGFpQTkP6TnBYdHz80Huc5hHYP50Re4/b3WIbYH/N5N4tN5uS4WlLpv3d0lSPZ1+6vgARsi2Ok/
J5fUTYxEm01q9qeB/t9zQyrtloamFK9+2DYMwjB5eJ25ZWDIJhJ7JQE8L8pa450FggO++yj0VIJn
nIJ1jvPhFSmDRF20rak+dtYSg+MpYC8PVE+mhmdWaeE/fV+BPf3FsWdxgG9Ee2QXQX5Y5c494SBw
XNO7PDG7JAs5hM95vwLKoHiULZ/957PTW5juObgiy8vTiXwh5ZC4ZvvetVuOwWadWpHWS+pLsMjG
ZZka+QD0DTTYDZaLqEBeUpnIt0iMYQiPE5Zi2k357977G3lBxHdu64XbTDudW+oSOESLPEUaKgQ3
GQpdIsDW7wxbuVnJT3sAoubRLz1wEr5Dcn1lQfaqefv2L0aTMU908+PUpVzF1JQaGjC37zDzxyCA
FLu74h/bJLctQQbtxqeIzmhQR4H/SZ+1Z8XUBxmqcwzp2Bs5zGcmYQJHk0vCsZpeMgGUxDsb520Q
Bx2lanZ0w1NEiRd51p9PJKVrGlef0e72rtfzLQW+B7NyRB5173dEaLrQhNfS/f/nj73YNUK9SHF4
syZ/Lcro7+hXQaYKtuMXacSz14S47RjMyaGTucRThR/sAPtr4ammedxt6zKpsAs2P4gtO/XvGHbl
bzGzMhN6kZnhtfKLcGBCXDPbdGa5zLhWI5EM2TaTvBLCYnemdM59q61cOuzhMIbcK74t4bwaPOWC
xHuirD4wulmPeUTXAXLFN+U5T2ifihexzdRkNx4Scd8vOY7xnn7qr/vA09doBZGCWQ83GWUtE+WJ
k8PeBziHkKLBAyPUrgL6B5fKKVcf/cO+iqJcDXaq6hoV+fmqEI30nsAer46n81QZpkUOOj+8WeVm
mRvxVYXt8zuh7jT46XqcvohrImiKyeo4jKTves2BQ+d9SqKitolIHqIz9UTGZoiqYQeH6idiSk7t
iNb9Gs+WoEQnECU5EyfItLVCT4DztAuECq3a1zal+ThbkkzNFugQnIcSIBK/+7NUKKNV48ZFtIiW
r4HCbi4FiDrIkfbZDuSCqqP5DfcWoLp1s4Evj/BCDHb/5C5e+REFFkkDd4ctu5kdh7yHZSF/8kZ/
1HrfJWAJdACzNqoA9cr49rv5SAodzyRF+CSdYKanU+QEP5vvdq3bVm/R4FAKwBaGlI/Ni7Z7pkT/
R3VJXp21Y7eqYpSNOP4Thj9JZQs6f7VtiPli091qa0NWSp84mUJ77KH+31GGzdS3+vX7MhrATxjX
wCX413co0ZsgSMsnHKdoq8+lzfMRB83mKSbUX4HfX/w78WWwgj7sWqYVFwVvsNShpDn4DiSBqti4
IuF0A7jUXxCvVmXyewF5xCP/7dH+OCgnb1s9XbjoDFtjk8v6nLyRkP3FlVWNbNpDoDVV+ZM66HJo
FrfxCOUun6Z5v0GuGUjIq3JDHCHsmw5fDXJ+1j8ziCu6VoqJOIHtiZTMwbksa+Qy2cPpCJEtgGMi
XdhUVSpOYTz3jzv6wFeElEkcOl3CHHAJO9sWe47BhbuQMGm7F8/3tSuCXlBi+aWwmHrEYR9YefKE
QkMUw9Al40ngxLMKWrvEJFlyjZ4acfAP4h15HKI7IUfNCLSe2bKPX8I5DDG632d2J5HscMV7nw1F
vg41mvEB9igccS7b71PXqD0K5TdIsWmjqrMKyvJt1MU9yZJXiVwEZQquwfTR0+ki6kqlbsPkaCku
ZCzNIjYWJBSqJKW1GXUMp40SL9s3JGjueKkol5RwbgF45BCI0btQOiwgRP+D8ztHxcqVKo6mzeam
WMB3dplOR3/qzY2X4Yjs02Dpk3pzzo8niqFkvR3kqSXUoXBzivNGWkvLzT1QIjpi745BJLiaO8lN
LidQb5GEOttCx1/NQk6/qxGekTCC34Ag5pDcsN3jkI/gPhQ8+z7VHsf6T33lv7dHIXiOU8Hv/bwO
53ACFgl7OWmAA1NY3VQHhdnCcEgqoocRi5Cl+hcNr1L0wsxb3q+SO+acy18gml0TLT3uoa1IE2AW
kg/jFRYyXy6F9vOhOjd68krUyMvzScn4ne4o43OoA0fWaLtPb5oXOWsEyhCkPU7IdihaNlYQN23I
xq0uMZnoSaR5vQJc3XmDbBZHom/006YujCL8H33a03l5+RDFfHhEQ3uGpIjMJkZssaWOkFBMQ4i7
ggyNwPmJcZ/isMUjy6y9A8JSYcRABkxV+elBvwAgHb9pmC01D59oxto/CmysjFfk8QbbW0gWAfWQ
AUeuxyP+JwEzOmRC88t0XcNpXcXeoEkx3IIYw8xgmlhiN3TmA838GgaS5//eFMLVr2CrQlaSIcLI
yU1Qx2gpr7SUjoObl5YRWtYxuhtsB5YsKktL+z1bTF8mGAm8R4UXyfKqDx9yLvSiNTrjMbvnJh2K
UdxM/dH/kmt3Y/C7iQ+nCi3jc74g77MHC9NdHno689YfSeBsZWLcmvqgHNvL1X9N8pfrAYzmcwOz
GTRdXGKjLmFj816hF/J9w1iq5uN1Z5nTOup8bPc2CLzxuLlwwfhwAF2ZkBZEHKXx5pnxfy2LiCZJ
LMzsXjw1GBUEW8GnNaP+PNAkpR54KrXLtafM5oIdboVdnetXjtNnRQXvb/0J8tGuwIBap+CjQy4E
HVV7YreA4abou660G3ZLImpVKZmDDETSYoNpMwz50V8QeEaYS99wv1VW+Be3RlKY9TpE7cy/eU0C
+Pl4CTg061/VLa2CCxQXKTz+9HNWGkQAk5U/ak+F8HMvo4/MmD+92aNj497/qp5ZebBya0wu1W+V
kmIfvicFWkDLs1XdCkKw/pjkue01VB8mwbdN11mY/iiUyF9XrIaTfez74sTkrYpQ2EoKkXACX42j
CrM8RPS0eX7H3jd/EoqgcBfpHUrqRj1pDB+Y9N/xS72YXjfZPStEEPXEbhWwfTEMz0QZN0J9k7J7
cfm+nK2NJubJJ2T/3vzWHvf7s5r81S+A9Tnk1ytQc0NCuq2/qcnqFNqbuZ1o4A9qdum9jGUNAE7A
mxBAdm2IeoPkUqDgZFQ3x4mN/KI1t734tDG24RsdQ487UmQugc4GKVZovf6aHBVP34CQx7HY+mzV
gMh7hSWCsRh8+rMWTCWjvZki6iRPfp6M16pVSj85Htyxnfxvc0aDwjB18Vu4V6YizbBomXsBKIE9
ozmEpnfAKvUu0SFKz5B4la9fxAYG8su/udpyRlaLKkqZAPbQkqqKojT1s6FI8CskclBpQjEbx+9n
uJfdkbJMXmy3728lw2gQrHWniWUHbMzHBfnU9+sIQEZFTZ0OBPCucXCHOYOvBMK63VbgNX1yElgT
fqh/nhGK8rQWrA/jZokyd1tjl8kDpxGc37YbJlyqUOQKdb25oO0P5VqZg9TUh0+NIcDXbx9mlT1y
CqgbI/nMhQWPiwszUr/QGFudIZG7lhfyWIXx6mB+V33cekAPN2fKeYGAJV321aDg0wrIlhrrbTGN
KPmVcaWp7pI2j3x/JuEL8478gpJHQTVBY/wackmRdCMbbBTeGwRAHILjOj48d+jG4sH77D71sYtZ
fimItpfnCXDuUc9MWlu0tl6Z0glfZT9vVJfbPhJL0/DXnB+7xlHXENkRgLcz8xfmpT5Yo8z48sta
CewHCI3B1VvvhAeIi/68uy/tz8eO/4ICwb1jcjztq4SEPAcia9nhj+9PseOtW5xEGzPiKv+thMKI
Hd1LHg9zVWv1cCWFgykMUDnEAZA7CnNTnbXvwokT1qu7bGbpJ4aBx7iGnY4j7bth94aNkfUy6D7B
LRHR9zVdekB73rmD7BOLVmd5Yqh/FHo5lM2PZzewJCf6gzWUyqjMEqb2QkkEh/vEgqjoDonO6eLS
fIRUBab84h482XkSmMUmpWmcorjiINnBTJF11Awn9TT4OCRi+aOSQOTviuAPBwmnho3s9UGC7RoY
eTz90Uxa5OHSyb8cJy3tFV7Xv+/5/8sq+Kiz5jiUUtwxg6RbOQep0c6Rt36yQ7tAi2Q1bo2FTm8Y
TxNDNRDJLHwgGEVnzOp9UVBjxGAywoTHmLmljhDV+u4hQHeO7rOb6tJnUj7nWN1HbeTevfXy1Axf
eG7D+ZgdlQ+4v102sqhOQDgeFd6z+s/Oir5w483uEUcyHvmPV/0PlUGOTwh+FtkDOr+P9xUfc1UR
vNrozvTavNi1BaVTLZ4jhewzhuS6BosyYSOUKgVRymXjQSvz71OMChfpw1gjIc+GjfxgS7psesPt
8XxW8cQ/ZYnwneXAHHQQYsHQ5+NRFyKci7+FBP/zojrsPWJUKHXdd4/QRnwBOfs4/UOSidDdRF6o
/vUyrDRQlYE5J7o4pABlpdB/N7BZTC5SCBcclp53xByusnVOAKNmZc9duir1beJJrS0nj8VXSflc
ZuSg/bBOWOXj7F9/DehX0wUmMcwpLIeSyA2GPUUBXh7Cpb9FvetWNIidn4TRiXcfBZnYuQcfQVsq
/OrzYZqlc4Cx3/6TBK2e90Mx/gNd7jWjRqSyyrbdN8VRPg2lyz+dmo8OtUGsL2bgPrM0+W4f9GAf
RNdrESKUxzvj9pMGIXvTwcG6wRovy//uMCBEzq9UhcZUVLvTKB4xdZ5nr1amhy0CUcKOIsTPlEed
pmx0nG+HHBqpoheKlwgwS2UCm07cXVnKcilpJwdvLBrlHzfTjIZ4Tsihav2BuVIboggQ9vqVDSsv
vffQG6n/C0aMvVS3dEtkr8kHnC4kxY35BirA0kGxkx66ifDTFsPXqBDhUroroCmRmzSXewQT6yFv
yCVyKMMeRcC4AYTTSWpNlsbW+HtgUwmy6esu8bPUCg2V2hhfEuajUkAAxTe8dBPFiGo4g4Hh+M6L
6t06oRO1d5i4B/sr0PuZD8opC3oDweGxxMRRzbd5D244Fp/OI6T6ESGE0zGpZLqjm9ifD/8vBvE/
hRdWoxPeZY37H9RvAllDrJ9poRMepeXHXPrXt13YH0bW2ow/Snw/9FrVAqTL1fhjJyMqa0Skn6pm
5Us6xEmEx/jHXgC98Ktjsavty9IAflhchDojlPD5wk+7SfotJWxhqz6tyESZH44XwQwaQoaYeM1s
mxTmP5jKVf6+UOW3GBehjybofiLQvVoczd/4q+SvnX05AUz8UoTOIyzedOKJEy+t41B36Kt21M6/
1TaOk+kvnfzHd+UkrvI6/KYEXsCekGS/JUV7sUCbIF3qfHXVDvpP6X9f8rh/gHiUunUFPd83AktX
H4tLzmDeFs/8EMXelix3mFMPRb8TGb8H1OuG6X88OaLkrphQ9YoVsuTXDEUH6YK6JVEdqzqcSnZo
wwlaSC0duimu22fT9I+Dh32R+NcYW+kPvUlPhIyRpmWlbw+6O3bvtl+1b60KApZDYZbJR9HpUmw6
ewf4RCYHV61epXZT4vV4MLeQ1ugadW05B+7VsTbmBj63YcbJMCzA33/z1awmyiUjLbW1Cj0I8xiU
dQvwRQnWe8OMpqbN2RJidevbacwb3LMrwI4kmls2Ps9zWvOcrVvokSdaehlPQnb2i4SdZCEwTdME
8t64XKqolZb+Oa2+FucufkTYobIA6xQZga3ACp4vJ7iZz5BwSrI01gIi5UcFYQWPVFgmUNgxcYRb
IjJGg4piaUGBU77+9RcBn7LMS8CE6WddAav75Y2VGw30tK5OyKShIVtYD1dv8CtNdHFRNmylLrBf
bc2pwsIm3mwFCQFBQwGR8/2FxuHL8zF7vWJuaJJRPR2wNdgfguHgaBu8T5fcPJ5E2fnJG47Et/p+
Mb+LpD+1M6qAfqp51V5vLUwJzC/bC+wkSkwBwf+4jk0MyLOz3fNrnYtNYnsJe0L8wE2VkvTCrpQY
ZTdzVpL+Tyhe2puUPw7GWOSxM89qe7OmGWmAgqlX1SDumePJjQMUcpF8gJHf3lPahHsmdEL606+T
xylteI8Lng2FFeXyS3uq8rxerQYTLvm6On5iQeRVNZEiVFuKdMvkuBHAea4GVn4UYz28xbaWwTRU
q+8woxeeRxoZDwFOdGGtHxvdoNGs6L84nOin9kxfzCbxvEJCVzbVA2MucuBbbERhWJjaliKC8utg
qVfq1U3X3JX3tSzctoEchVCsb3kOCulT4k8maNnR930/JUDyqG98yGiocBskys12sVebcD4snwJg
XzBeWkR7D+cK9aRRofUdcm7OxgjHTAdfp3hbG1Wg9AM15Cz2+NdvGVS3OLiPPmDj0AbfhqhNQLJ5
ZYl0Cv7MDaGMjZ73BwaovqfR40LdVlM0N+eowNUaAkq+crKqca52I/RGQ0EYbfCHZ4D9HtZelIWh
W+Lgy3m7Vao1yAP0pBkViySmFIkaKXoKPi1M/QFDJ8gcThann2On4suFUx0FaHZVtt3b+31NUUKD
qgK4x9BAWpdyt7eJA6kmdiLLa2YNoUaMYw0T9svDsOGqQANpOrmHDBcaNxvYsBfXEqgO7eA+0SgH
a+4gdtwyWZsz11bVua+fwFwWMB+nPkO2Jd0hmWdXUC2lZdy9hDLz6eBhu2IPf0H3wBUmQrdhrB16
dlmacdlQuYyHX/kNyZEL5jPhdXww1xhdV6hKlNt7cOXIf7Ry0X8pFEoUAWVMO2rUpCbVuEL6AP2P
BCcYI/igDaKY0Rr6Y3WoiIKakfqSAYA7DKW2a9XNHqcSh2mGonONNDEkdMGvX/2YZDX5EuO7Ec0O
28bVO0XwjFGyxQWOm6hzCAM+oTFFgeXchLca7LDMeHL4JFWERqVISuEN4al2k5vkMQNrcVMj7gDx
VxzKlFhfVuVTJPrDSYFJbAFeNAibr+DREiH/2F5eaWMflI5YMlXDLKaEmh18pJorinQ0G5S1cDe8
ELseYu8lYqI+BMGfyrOvthVpnaiZw2ykmZWrFvDbVDHlBa5g70yX8iryQTe6wscgsmKas/72GmaG
V7HQ1GLTx4ToZKCic7O/quVoV/Ljhtot/fBBZaN8y8EOywxFE9GmikjSk5bSfjoy/krH05ne+ywC
m6bX9Wk170I+COIBNE2SV4SQsBNpt0iV35bLHwFE+TOIBciZfGWVhYnqFwls/JelYmeS/1gCv6vk
4sE/gpv5gbOp3Mdz0LUCbAB6vlqkSZ0/OktplU8+Blg4HiIqdDNegaPx5cQBIIWxiFEx11DxPXeg
nxIT0mj1jC7QviaV1I+ykegwVKvnBN++YuP3jDtJgKDsXkf/5ks3l+xUk4ZX1Y97/2vWw3LvjaHr
I+ktcR1LB6l108Kuc9Y1o6M1UEISOqhrV0LnOG6ByJPW/uVGXV2PcCYhCpL4CCI8jOZgmq36cDzU
dqcKPKXE30ITSITW7Y74kTFoXxLmE81L2RDrhYE1Qg6BaOn34azp+rvWVve8yvILPYdrJykp4Zvs
+C2bVv90VGU62uTqtXImjw5ImVSzD6Z841l/KmW7zIQFAQ9rPZcLPsbXpXBahenYl8GJOJzxIbSA
fnVaMUbaNOMGxN3U4Px5VRYXNKXdMTavoZEM+WyOI5eqB9vUNi2Im74xr88dOre6BVo6/rzVh2Pc
rZH/fCHvlnOHWx3Nc2NcYvKmSdMKiCQ6OsYHu++HzhJhmUJWHxpZSpwAQemQkOXJLxiV3qjdb8YY
wnhNm8uhQQORnIfb4bNP7hlxOarejgO0kcSD85ZL6wXZjNaM7BvslTjfwZ2xGUF4XlzL8vqfdas/
yt7c7v+NIgypgYjOWVAAr0GoT2jvFNeJb355GUYNCVtynKX7Q90SGIBiTFtUB8+WuT0UUw9dKWWC
4IxdOTPIi/U4XK0WOp2IiJ+WYANMHEc1G2VPl+Haontu4BTJWYIFW9JcbYQRWn28nEB0V/WZ//7D
lk/CKFBABWNEoptN2t3v5FVhcv3NGNhmG1XOOW4jUOZRfhlh0YpRD2w5vNmKpUQwyoASRH1IHjZE
26/nBT2hesRWtmg+Zx7M9ysDz3QwmFLEHDVNmF7Pq3okDSjwmqU/R79ebVvk+4nNYCUGy3bCrM/J
8277FoUnt1M+5szN5abFbMcjpke9SyCHozYzSPJa+KggeT6iTfNncmg/NkaquaAYi1miuIn0zuTk
PE8gAutD2r3JJMCqcG9fqYdZF/YOfYU+BlQvINgKg/7m9Y/XFKjgMPxLOGrPznMTgWFSm/Ae20Qv
0LUQgoRDH+zJ5pWQZhNBEDYb0KeUOOXSVIw74UsoiLmOEq4iFFgEXpfhYxRgr2I6ReQStX8YMzKP
OPZhgn9UNkU/C4l8Zv17/oTO3cEDNV7pr17BP2qp9qT916TcroURV4yMjsJPRBVEcl2i8BXxTQ4W
z5jugLwQgF/hIydeFai3oogbtEth+Ljo8JMXJq94x05VCxglA3iSDej+N0L87B/+uMAsE9wGfaLR
o3yhRyRwpA5kBwNMU/MQ+qaUcTWCISMJ2yWH4+8CGlLlT1UBMWe5zmtik3iKYl5M9RAuYKb8nFKn
pKergSyOQUV266tcqZZGdxC1Jc2sBR93sJxru+faV3Gtdj99nYq7kbT2GeSlXto4iSKzszCOIP/9
UJPwTiUJWDw/GLGTqUXz287rDR8IqsnhljTLW7zNvhiWfL9mDzvJ6xbjyCks4qtQ2gkYfVZKtjaJ
Tvw0YlJGu3pjZghZ7U9pG85DU3JYKdseoo4D+7Ns/gz6L6ZVGbiUk50IBVCBU0wntis2Gs+Z+X3T
NFhkzS97rHOyY0wraISjb97cbYIdsyEdI2yHm01oxpVQ4kYjpN4pOkTvEP5I0uRyKsHFw9HxC/AY
VATENO+HB5jRm5CpZ8j4xQ2x9L/gLHuwzdel4puPz7eXB4Pa3u/UBMPW1wd8X2r3aXqjTg1WRCOY
kH5pNvw6OLegrPO/T4HrGiWZsee8OBRY8N3oPE6cs9hSqe1tk+LdNq853sjfxn0bzJybmoT3UC+s
5cG7yHgzgG5LYaj01hLj8X5l/HhgMy4BbeoTKCyqohFjD7ZaI3LYiKHFt7m/O4VFcRjfObxg0EML
fpY9l7Kev+8Cnhj6ufhkgv0xfTvHj2+hBuVKA2zA9Vy39AK3b0JjBp91bADSEHoGH+AknZ9sO6PU
inNyoxsuXjWgB1S6+Y6FgNTZQdtfhvOtXzeWHUgSQZWY7WYiVAQMCUMZup12RvN1PWsZ2Zh083Sz
uwIX+Wjar4Sq1UdPuco5itN4v41a/nMZvdk4lasi430WMRjOnzPvzTdjaG73IfVNKShxf2vNyj93
LC8EgqUUth1Zx3Lp5PcUGfLxOU28QGd4Nu8IE4HGTwBXbuUXdHicz8WNNoFeW5qH9fHGLGHzngHH
rTzHw7gc628gh49z9UOvEWLcBg2UqmUFLzB8Y1WCtNBKvWYprDxjRcYCjFR+oGctXby+ukzk3hqb
ixMA0m9jspwok2NrF4evoyRuikQrQqml/MLthOvEvpY3xBFJr7EGr9oTmyxkS8IMwf6b/ZtXDOXc
KpANymBDEZA9260Ju+VEpomGQEK+KFL0pPDFLIFafAk8pJ9R1Xi0bK7zNe87slvgFvo4msYY9bir
IOKsVhGli9N3OXxGCBhkYTvvqXVjx7y6gFI9xQV5hHYB7vbQZ608QzahpI0+cHqNgaZf1tj+gyyE
SrX/nOElCW8TaKkgPrcLT39vXMmYCwlxrQeqmpccFkkYKXb/tbxVsFO9xOylNKZp3kIFhkG73Za+
4tgo7y6QViyk7+/5KYQX5MQaiKN/mP7smSXkh9rR2qe6DNNGS7OC+Zh6u2v7stlOF1MfaDo6+LMb
XmRf57HrsSrGvuRA127J4NIl5bnu6Qknv7FWOveS3kwaQxKZTelUFZs/mGm/TZtbDkzhxgB8BmNS
/IxYtYiapuKZ/AFuXIoIkEcXP9ATKzGjfnIpr2J2m9fHvNTMFJk4wV2VZd5CN1/yv4z5ytKZtHui
dA3+UCES2FKwMFqn7GCLxkNA6BsKsTppcLwIEzPpCkX8RhqCByDjpLBhY00ytvzFwTUDdwDzhlAG
Ruu6IrsFnEE5BpVu8lPEyCPgfRpwjGVusnAc2oZVT2kiEA1tfEfVBvPanqNIB9g+SZz2qk9+iP8M
xk+5nlGK4pcx95Zbsk9y5C193lv3UKWW9oM3oaK62/qiX92/QSaQ66s9jG8jWFDZksBbhVp6MOiP
GQyFoyJo2JWjaZJNgZ7/iMQ9Mx9TbH8AVZwryFpevQgSoUXBVSgy4MokERqBPpc9XCmA/kJO+Svt
cggrezJgQyUBpOQFwQz0gX2z30YgflTxFpj8IoDbr4uTBO+paGA2ONmY5jcpKO9igi9tcjuqDwOX
QQkQIaNvuquKnmiO3+MZ8nhf9+ArBoS1eXYY46WO9NwVzxCYiL88pcmlbXykla/I4RylSVzqH34N
fWOALOfqaUubNuS8NWGLlyMkABdfkjAPq/+/XzKLPWCiwez3RpmucRDUlhZKE7/MuSSfMRivzI27
Eb4zHNV5YU/NnpMBh8djgX1fTnVr1k4t7gt1RN8SU1YhDVOMn8NWSt1AStFonVuKrrhegkxrQsYO
Ddf8lW8UgkkmOAZ6Vl78O0muCUYgT454Jf8kSnE8FTb/BIbkNSijPM/VcRWlXCfIZeq62eNj5iMi
PVt8yIlnwa4V/ZQtH5aWTaSUBcdEdefRrZiZv3RdbBB3ksOzYI/TAO6AhorgwUrgR81S+hmDu0IZ
CorCJ4nETkFnO2mVO4auXlHG5Qp2Op2d1mqlDaj8c0obQ/PWlr2BC1+iIqED0PkrK7bwBVu556Ss
+rc2j9go0AUW1tP7gWM3euNQ0MiQotGR/m0moblZ1MH+m4xMUN7FQj0gUKhmDAhHAjyWUv/GN/mx
p3DYUjXIC590TJSHTFk9ZtC21ysqrArukzi5YVlaaLX9RaoYzV+KGtSbX2hv17EHPWD90MMUkNCo
nZWsrhiEU4KDEn3SgvrgLhiGdJs+Gd0KQcUGOtIcWMDzrprpbR+6hooJtPFX4FHWYqy9qIf6a6Ru
/jQdKDuyBwp7SGmQi73gc/Pc2rxUGhKCoikbRHNJ3KZXrFnUQ19R6QOedLizmEhy/P8WQyomzns9
oj2MFcqkTihOiJ7CYHQ8/Y2jWPs+fx4/jqZYjUkm1MC8xLuvaZ0DgyLvKP9opWA/tBr7yCG83SR2
F04JfixvVpZa6ljUgiEyXeysoShQZoPnasdJS5ilGLQB8TMjRh8ksXmYuaNmF8eb26Bza6k/3h2B
olqt3Q900+1MP4GWhBKgx3zHYQJ0s2G3ovgiZkH9JxzIRSzaW/8GI3ZvoQha3knvqArCFCe6iSTX
Mv7PrTq63Q33RjM6IujA/xfOK4671+2qiF+/Z5EvjEue1Buk3U9HwG9siyDWQ4Jk2VoqtFoxVs7k
czYCWu0+3EMyMLmGm7uzCtIYAv9wQhqIDbuL3XoGwoyquTi4a/LQjxtxEzyWqS7YvFqqxdyCoa/M
BngoYIaaR5iofcUMXyAMrslKRq1gVZl76QVoyEueMR/HHHu1ai4PgG38ppmaznJjvnjQebaRdCBC
lE+018apamipYSS4QcUoZQO51dk+M9g49GM1Xx3CFoXVbTDZMJfGOv7YRLa29IY+AufqCpzh0Kom
oYOQfpwpz2Ue19bAd9MwBc4m4B+/kJmxC5GXXfeFpDqRvO6REY6clbMfO0G9LvPd/X7GjowAPUbo
TKbrexhK6FX6Tq0IsuS8BIA4dPaBslrShjoJCaIDnrVs5eHqZ0tsI6YhKRQL9OKGsmtMwEAtDS0Q
p3sFbZLm07JvnOW1n1UL6xFqsSBw+V9Glq5HnLv7pvliBQP5DKwfRcfYBIh7og/jDYYavC5G1sI2
hQcbTqBRyazHRH7svOxy2AEV0V1teKOx5Qr4GV4egOchf0IJAiVpzDTpscMcy/CRn5A/Bplbg+Mz
lo23kqj47n6a70Ef7f8f2svi9eOvS4YW6B0BDp91PsaTpwdVyo4RgAn8GbtW9bsU37+dwD8bE+q5
d4Mr40XlD38UES7io8nV1U6cECzFNm5joEl+G5ns2K9Arrdt5oK2gYJJuy0fqYMdjbawcgrTvxy4
8O1eZv0eXdXdno6cNep08KcBoH8P5otoFczr7+aiXP9ZkcBdFAy4iP8az84+1MU0f4iT1sl0rnY/
/xdN0yHruS4KmGgGMhwFbO5y/q2Cdzw7WC5SQN3G5GpdHhgxLeBOHA7q4mddvtA6pl0LG6yfN7j7
bUhWweNdRPYl/NApA62XSuL/bW5IHfcF0rwsd0DOfW1A0fbwyiAJmIDb6bnz99kmgiMo2ageMk0K
6XyRhH5rFCk09J2WootS/0Yagd0ATHqK4iuU2zCuWDneQm/Tn/kEHdFDnXZN9YMne/WfvLlfNpko
LJdcP7z2AlnI30SEfXUr7AhvkX6arEr47Y3emlguTbZjJMHXGLn5+ch6QftmFouVNRszYRBWk0eU
gw4VDhnLDOooKNReNuTuoxHqzCl+2UILHTw/0Mp35K3SARX/gClmWbPqea5ew3L+K/Z/edzpXGkq
GHBy+etQluTZtk+h1A4nr33BxX1VdlWOB6CBr8WEBqSI9Nvv4l2DupiVoylgo3TyIWE6MyTOLDup
RD+PXwuJ3aG1qSXWsw6xqaE8b04X83EWd6aM9LA88jNxnyHZW1rrdT3RpFB1qbBWaN8KOGvNkku9
J1vir4Bt/ZHsk9HQfxDVJvfMJiMyU1BxsqOzpYmX1aCzDKRfyX5t/usKn5stiGn9gf/rqAC2P0Me
cH3ti+feb3Gcx235vIygsQwqe5FHm35tSXU95za/0d5OsK/D5o4vIWWR2wb6uaaaLUO3+K8PyqkV
fNMeBqxsyoU5ks8QAoSgrgoQfrxZA7wZh1r/aAJJnplV/Q2WEwcuz/NAo/F13iwuRQXZ4oC3Nthc
genrfl3RugOv6L1D42CW1PXghpZV/Q0nGDFIL3/0zqGI0COyZYLeB2j6Lda2dBKDKmkj4M0f/m2z
qyiK+SKe44rtWje1ZHXiAaZtiWDenxhTy2RIJC6fdQrHpEMCPoncyFoTeqS2GZ9MZkwNLJ6iEo+8
bqYtA0Q88mzkxSZpIxaneMs4SoPJN9hW5KrfzVhMr48+abQ+fEaJutM27pCHLtMUeTv+XHegJgup
UVKxBXILDxA6Jz2ktdZBcceBMyQ8CWaF1e6h4bh9GyeU95rK7UiEOGFQmUOce2UzLf5E73GGKtWY
Wz5/TwomMI5L9d4uqKkiZTIFMhKwwyikZ//iSe4BZZ4YKKP9hWYYBLEgZmJNjZ+LQMOYIhU8ueZy
yU2UVRFy5KeESTUnbzeiOgVaGqnaFIYsDjWaXQ8wOrA68pz0CU+/beL1e9bBbMkUNbM9zJhts/bP
8zqOdAndO1yoMpU2YDI1vO/ysbzxhYQtyjtru3Q4kWxge5G4F4J/SpFUSY2d9W+gtFkBFbkfRZTh
11b6Z0aERJn4ptVygtub8rjJSVV/FQeZUMktIKeJB+cf8B5DhiG6LQQnBzSU04KJnw9N/vNlKaFf
MvhjzsoHlY9U+jflNN4qoXi/OPkfFXKmswzUtgIbhoC7X/nIOCd3vOwazzwW+5G53medmsj2M1RC
Y1pHgc/SBM+kSTy8heKyxag4X+5p7bQaKORFVE6xpx2TTWDf2sr0qCKm/p7ZbKKI8wFce71QkclF
30ZfyB5/joFS/U9k3u3uGFdEtplng0SMeazjFXjNxlxbWLkM8D4T1JIlOpVh+GsraVJ83T5pmsI4
5Cx2He7lTqF+nF6x1hsWacZmgKllzmZfakRgV8XfVJZ4gZ2QIsG4GIBmc7+KofCPmIe7PF0AMsYX
tRDFZT5GWJM7Y3WHrU13vIVIPe/G9h6NzZn1JUjruBg+S+XMARMw+R38YJXWxgBzwEXSYIqbjpZn
gZhpdUW7JAGUWMiFdjC1u7bbq8Q84dDJ5LCxVIgQE/xLKX8/2wqGF8XSAVO/8fF5W0+Gy+rk6pWa
UHLTXFl1/zEo44F17AGrop1TjQ+iOX0GIaCWRe7KhInEq0RHYZ/II28JIxlAdbtNcAo+lWFn03Jm
k7lQVaA0prti7V+e1JbhkxqMac7wg9I50ccr3J11ebhAYGy7olxZxWGGIZYnuA3pPETxceucwirW
fE9BR3WGZgeAcohzYlnX0SMWpwHhRux3wdSYZb5GqmyBzQUz7DWdzTEs4aaezqr4+5GS3UEMzic8
XetBFB97Aox+OzOuhrGc7FbModK1ywExSS0u0Vkc0S1JfLvvyHeGf63vbfZ5kBtdhXKRWnCGGpYx
Q2DL5iHpEZfhR7THMGahKsbjlbds4RoVc5iRXWmQKpNJ+4MYfarHM1pQkd1ozZnMBGe8L0oiuRHb
HN1HHt5uigrWGEBjEgL/2hEGHxFbOWb5Omul0bNayDhA1beEaK6SXgP5uccHql1InouXHw/5WlkE
ORyI7vPwP3UTxMiH9J91wHMyJWE5FnVBdNa0Jqur/tMum/sg2Y0TXeg+M7f3zr9EPr00yhpbt7zn
sn2YY7q8ZiakT07mRVHn6/l3zrv0d4Idtp8JzBhhYWDn0Ufv/RtyfBgyqGoMuqaNCXQXBTlI5xlC
vbhGSogrdcwgkEwT0xpf4fTbqaj9V8uvevHq8wfZll53HVQvkvrJpwbZTjT9qCvmc6mpC5DmNx6W
fpgBIUcPw/BXmrQn67jI6HhjcnqpGbzOZL9LAVgaSse8S+tc4uwEJJJxGRLwJaArerzCO9rZMNn+
dEbbo4NspzIW4z9tlb+m3Ma/CNrdALcNMp3KzTc+kCjm8QMCC+4Fjphquph0+TTK7SwmawZTBVKI
+TfRr5GuDLUPdxRFV3103hxYZBG5JbhTfG1fHUQQhVPl7FV6VuYOKswnbA3rrTOxLuqRlmPmHjf4
cckoyjmRAmrhtPb71UKC2x72KWsqJsw1Q3pAz2xdS+aQTGuoL9cNoKYsG4aNNn2rGkvrlI+h+dvw
8AcFqBTeYjvj896ve6Kc9RD2QAO8sWiiWvSEZgx//i7HHTCk58yL06LC2b7a0JipcUUXy6G7+8nd
6tKzxI0HZuXsw80VKiDuYqm4IBczwhdoznZNm4aAs9DVHDrBNBJSDOahgCIdrAuF5r7QwedbW5/A
KF45FtWgJiffLk1P6nFRpzb6rVpwefFMHL1oeRNR70iFMqyzN44RIA0uGP9u+GskIpnvTDFc+CdC
nXSVfeuKWjbeOrYJfu89Z+y/njWTpYdO8ThJ+fVms3BFAEhjZ6QwUmo8RxmaSfzoKqQA2o464Qrd
7UZKfbZA1sybnbvnooW4cw8FXa22u5AJwYnhdqtI9SGyLHdWKFGmvMGbz7lJ8vCFBccsBAEMuwSw
hnIXYL7EiECuMfUjTxGXnCvJZokKjurtJKZ8bAb8XmBez/SAR0ri1FoVR3m+D6O+C/TgtrVJAE+L
F6gIBJCij3uVFw73syXfgxjWzRS8LPvSQU7fREu90dfHSw/qrRVqGS33lrOWRliqMNGExqHvQe6K
kldOWfZM4oXqWa/0CqJMt0sKzdIePtH7Y16sGezmKQFNc1shUCBwNwsRAECev4ljHJUKn+7xqxjn
xJnsSKXaFQBupn+54qlu+cnAV+KsB/xxicduOgMaEluDxMABi7iFjDHYiAH1W5A1fosGAUbZF5AJ
jHFOJBx29IhY8JJEKudWjv+0/H7+r4OVC1Iddw3LEI1DUl1KX2KxwVCmkPpYgOGAZeQjUl7cXa9H
1pd/H6qo0yXk+wDNv90lrFuiDY6r3DsZHBXrBd+HgkoQU1eMWdhSTSbB65zv9JQEeY+1DXtSpcUi
VlMiCaUi/VDk/1HgQm8hWFkyZj2x0J/7P3hBZhIanR7fbeMLJk/1pR4q0PCyxblMsYmLMwLkH50M
0+eNDneQ1wydh0J56fdSAIjrYJK3Z8cDtKtVpH9Q7JNhktXhuAPw/Kyra+pRDVmeTbvoL1tbY0G+
YiYRRIVfitmxx+OljYeS4IFXxOtc3bzN1BoYUz5V4uoYCOAkLO0ziD2rl40YWbs6eOMT8hxzqzgS
uRBWCNZZIGZEFcUIb3vd9KPl+kB977XobnCWJAPtFos9CSPIACNPTS3cm97f9r+n9SBZFVqpGf98
ecXijrk9Tz6ayQK/UhX46uqIi6A/N3nSmNncQ4S4cE3vK7URjVvhxA7JoE08fRAqkuNXkzM1Y5f3
+N9CDUmVtgFSaxSJm5bfH7vwo8k6iOc0wD5WPn6teuIGPj7ifEb55e4mPw3/pQhHe7zKra81QWah
7+yxvHW0Cy8sJNtR7U1ar0Ny+5APnnmEOzEgAbTMnr51UOQ+nPxK1T7VHMF9kN8X1G4yeO4JZ/KV
Sx0m+46WPNfUHYQhH0/68kF/9YLSEPQc2jyDlzNLpeJZq0YlImAjCRy4QLaOe+x2kDg4GpBLRr5/
AOqi+UgCttBUrdvZrRkpgJ+32SVfoyaalJhlPAcewGnVB2A4KZEeudgeVIcKsSMI5u4L1U1LybUG
BkKXUxkYpTEpnQwRYLzIbNnBv7UHtqNC0BG9bnp4h+UwkfGu2qrIwOj4NdsShbwb3dQvThiLxbqP
yeoRejRNa3W0TCDhjg0CFkBfDTvYHYMZhIuftXjKiWcSDKJZNC9bR84EUhU5qas2umqx9N/JqbkT
N68mTKfPYaeIhBzweNsEBC3NFcgy1VQmPZwhuFGBMCNIQIhrxzoTjC4Hhp6wQdamkgwIb+9SFRGZ
NX3s7bi7ODSevW4pfyK2MMO4hPyd94VIMhJg33wL6ZH/vJVzjYTFAI+jv2dY9wnxEUyG4EsyTQZN
dJm/Fg4AoEurQTC2CjQ5qU3dHmi0QhZUkAHElCG+crYybbCp3ADZ85KpCgk5tvuWy9IhAViTSH0X
e240N2ntXYISLlBuXdtbs7mdApMNH851KF8jDJSmY5TggOhfsgwhSQoruhb5YmGoZSL76STUStjd
nJlNWdtANeo2B935MQiMS1sopVfdDKg0Lu/bqwXxY+ISmvp7kffv5vkAZTC09QGz0vU0ouHQpir2
iIOIMONiJML0RF429EzSKAMz0YmdBEq5cSUvLHfWBP/we0Qtd30OuU2V6X8SUmtqGkRIe8+rqRlJ
uMfciKdX7UiD6NSiP8RjLzAW3mc5kJUpz6eKBJA63nD0rQp4w5C1grOPv58C6PGdItczPgnUSPfK
+tVOU3tScx1BbUmj6naadAKNU47c+xuIJ24kCwlcnv9BUprZJBWb5HhJl40FWoCZpd3Xn6lk05SX
S0opYW5QF/X2vb7J+uoD8K7qPjVY5zKfGVUMNJRZq3OLmRumNUzPaBDOfZ+JnusfADR3iko8rS0f
ltw8LVNiq+ZhGYK+p1oQl5RKu8yIhXsY+9WQsqFwlC2lk1Firmfnvy5EXJx83n6yPLOcrhct/Hh7
T5w7GVU9NKrMTSPlsw0dFR31lHblwtjwJDnscisyuUIe8Fccmq1VGHJ83r2vOnoLZyZXWyfGzKJl
F19Pp3BbumX60ML0huPbaPdIFnRnmHmQVcEfnE5Qzn+2VjR1Q9Hs5SxQqaObYJki5yrJrm6Yvbtc
v4V90drhbzaOw9cGsxpVmbE0iZoAJGOUE7Nu3gbwLPxs5VyXihxofjaAvHpNY76EPEtdlfy7yQfN
P6ZWwYApQHiqMTQkxilSTtlar8BZzS9ADsg11SQx2o0Q3axK57Zh0AT6dVBHxRp6MW0D29q6whLU
XBVQaHFq2ED/YF16LuY/RuXM4M6KS/x8/ks+Ly1dn7j67TcBvWqaDBdmqpLxSjdV5Gp+XymzHL99
EjHUfPQHaBaRTOW/RRT2sZljJWj5ccMwZhLQhKVQ5+2lwepzyjPh+v3HfYr9j2r/4CngFdr3wD46
ifLMGdoFr2NH24VdAOmG3QRb270R7+nPSwE7K4F5e1ciYmArVVZdjlAEYZhVCp2Uqv8fHX5xr46k
Qd9C0OMWgoHlmteAZafCr3nwa3NPeWvpfYnfgVHu0vkpyXOT3nZMXmVSZtp09a3iUTBMOleEDsMt
lIL6dYv9TutI3O9dZ+QpHHV6VaHgLQ7yhN1IRYXj0WokL0uSyd7Sv+IFB7N9ncKSNN8C3PE115x1
1lLDvkJywXUgvE1BxWVXEKoG3Nsejr8mAy4jwzvdR+gaeWNv5Wv3RoSEPGnoBCY9AGv73nAX/Dvr
fd3VSTq/XrMDHthq0Oe36R/uuMGkHdNQ5a2mgBpcskMltaRuEou7zr71Ok9v/I8roCRzJp6vI2iw
+GV3g+xGZb7jbWV2EWiMgdKJxbrxLR94P2skQN7p0eGdNJgaei5Q88UV9hzhzk0HUZPUITb4rIwX
CdOx5MYpmrQjScErXdm1JQMRhTgVBay9FhVVAM4cdPXheheLDQeClreV1m530JFzqe4NNvtNlntc
TFjpNCIFxX8Q/qq4pOtGMtNgZNuIPOAcRebErjhH6NqUNjLyhRtiCTjG8+wmrvhQtaZb/LO50bfr
Z1rVf2Kzm2v9Nsfi19admnsobyW0DFC9kG6RvjUefc5UHxi/4J028O8HCXcQzcYwlnRO8YgGZWfh
8s0UK4yrKc5VKMjVxipGzWJdfL4XO8UX08jdSY7Te6TUc2CNuesf6gK3kM3d8KbrSP3XAQUee/un
rp3wPSv4tpALMJmriMme/PYCjGpa2k+S09DmIIePE3JKWpG1GbwVRQKa6AlNX4wgNQkQ3BQZ9ePu
m8pChvE1umYaKVLXclWuLYERM/RqAILprr7Y3PNyDk6temIT2U0HjMJ3jzrwW57hYnK2WoqVuOU9
DgOwQZEmI50SDbGdiV5K5pOuBjMT4PYfk166muYx0GQ8osbokqjJqIheFkKUg1ipbuRfH23Yh3Hn
4L+TCn4ne0Od0cANtRLLgDI36AhiJ0bUYsenmuoLqTljiyjLcCRnwvZVNBJbUx34grJETzT0Jq5D
87kNPirGe3JIM8kbj6CJcoby7E2/eh+O5WixzQJF67O1L7srIwLby96eznEmb+Pm3tpGLhVbrfki
QqBB6zdHP1W1N44C4AdhRieZjMqowiJScEkw12j9Oj3loGgz6SkBG4Wmbve+tJ6qMeYlU/YmlJeE
QO9+9gUzhGyxtk2P3j7LzWmYcQZov3vfnhmV4Iq9oOoR8zj+JVFMo7nKF6MgIXKhjkqzEa94o8Vy
ZYxGnrpG/6FI/HaRHlp+4BE3rrYYyZHNfkRopCTVsPPwgRsDHI1uBQ1ICd+dgdqRahQu/bVG2vxA
fUVHELvN+8lLlsJctkw2tA8hEw1Yamwk9JFT+c1CZFRPo784uX1ecmSPCjnbtn0z15O9QEUbQytX
bH3TDq6PAdWnVdLNDF3YNrFiHGhw31LACJkZkb2Vc0mDY3ZBZrfUwHyddlJ5UOFhuefMuAEKWpcU
Hrmjv8AZMmuj/c2ASm77cBO5ibul8gYIjohOpYa4RWnG+bl4w1CRLZHGrY6tr3R4xg4kpmFE9rxD
9m4zC1vM82bsiQnms0WAII65mTYWcI+tV5+KMSvUVrjbaPX7abb3NGN5kznmSnAHvcX4MQ1FYlQU
cRcvmfp1NF/7EFsLbJ0bmyQ9mYoWsw5QNaKCYPsP1hsVIGvmx5XbvTL/cakpRBChYYGm3zEcgqp9
wzStWYfwmY1Jqlza60K8AD7+RXPhVYlaY2r6FJX7mAdLPNLvbIzZ/4zm+IrSbnJlqa3USq0AVDDP
Ycm7Jc6OMJmVosHBrIBi6T04zZHxF8ky6moDCu0RPdkLAelFlDx1OhHK31rAe8D0noBwX1Un5gct
dsesGxyPthkJzo/10egeCmD8yk8z6W10DXiKGFpViZ60VgYXhBBA6KUdCZ5wrm1mMG2+20MTL6oM
g+q3MnPIft4IEL73cGCCFgXwYdERcAjf+OVuHiVRusDeJDhGr4W3dGbEWnYyth78Q4wcQ4L1YmlP
O1wtB+lfurHwxywe5jTTn0rC26Ja6SfjVYXkZptMXmj4dPwA0MMlEysORLLx5M9utsj0Dnu/PbHy
e608+jE+tHHf/sI7XaO2wNZaQ3x+Oa6vo0Ipyyih+SHfVDg9SWrdlicao5dxvwApepJijBKnbrf9
B21PXQ2y6YRe7Hp2Hn2DPzl6a6tAKi6L1sACqG6oRLgVb9ImMPraBlOfDIjHenKcnvykTWiCsY59
KIshGj6i6dah33ilahpe1Llbk2sd5GA6xKeuKTbfKt/cY0fxqAEs7IL9ZXs2F1YJzDwCFMESOJB6
iXhyovoRNaA4JIgk82oVy7Tft4ratMlq4k2IxCZ0mIfPPK9HnKN2EF0p2Kpq3BfpVLp0S2IRtj/3
0S9y6eEuOWESYroe79/IMKs0Ge/npMWRWQLT+M6fZhrQOFdm9QvWm8mryEj8oykBCc8c4DStQoQt
kWsg3Xg8ORKfnHyUDLDzSekRq3cr56XGmV+syQB/1keNn5pCbh+gKLd9BRa6fScuV7QKUJTu4E2m
flQ0GkPudC1jfJ1qQv5FqqXntbu7db5eVI+dWaoeK6g0tSZLmGtVSgPFVsc/owgqr0Ue9dbbrgGN
fTK5v3jfKHbnuuy5zBVlnctKVZlpYDg6mlSVr5YrXB9p7JoNVFxu/SWFzOaMNHXEVG97SlgU0vkM
M6qQ9JOxHnggeE2BSpCrlvkrCok03HEuDzeU/CveyyhTx+8GYP44rtSwmOjldMaA8O92FMA7JA+P
R/1R9QBuvX2R8Flwh7XZEsMu/zIoJYWDrZZn9EIxgw4HNpJ96b50+92X7XHak7U8O1Kkx4tdPQbh
ieMQ7UYf3v6BzMNRnV5XUg7LHDshNVPsKHZ8NjJQIw1Ig0UT0CkYkN+Mv11kOEjQqplRM2/bxAmW
RBD+YAE8rdcYblawBLmqe1wUfKXH5yKfUO8czdyvvBB5MwB3w0JRvXurxdXCz3eRTrUvRVcSTRug
9VLtzDo3zRfRDxZ8kkfRIV6jeAIWDVTwcTFMVSRXwZ6KvCQ7QtwfhDr5c7PPRFI1NHH9EFghNSio
DIoWBIvsvrwKRL2UPlDxF0RDB0k1WDaiQ+KwztQ9HJTK9W9sfhe7jr1mF8R7mR5imdgk2UG+YDzt
5+b0v7F1dZd++axg5lH++FnCj0qrvL89+qSQ/qC7Vg9uAhnSI+Ogto7iiZ2ZbOhyUvesenOVFMWm
PSkJGoG+FI22SNwWsED9FgdOwHEUbjXRMQ34UUsQWR5fdcKotyHC/b8A9UQvhKndVVsNxJfHNB5I
aYDb1uc39ofQBr0mo1HtzPz2vFfpxbapx4CtjRSytCq2gp/j+3dT/SqiVZX6Lv+5yNw05cjCWYGW
gBb01cssaS9/81awDHUBUw3psIsXK5ueOcaZ/3b+5jOu9QRenraOo8H1rWp2R6PaHauYDfL+sphh
LfDergoganbTdLE4wOv1cjD+KLh10KByr6VmJ1jVY990b7tkcX4X49s31JM6J54iHoo/LkNHfraS
WAkilPUmCKwHd8loUmCu+hLzGSIg7W8kK0o6ZpV9iWb5OO9kmGiSFTLerueok/O3QOYlfV7CmghL
2bDyZg0LGBdEVITx3hG0NE5J/Xp6jakaNaJSxr4zlyB0pG7eZcyDKmPiVAzzvqPbgGMyzh2Y3hl0
uj9cZmqwqCXv+A15kVIMU6f09J1dHHRgxl6Wg/Wj0LChaHbf9iiEp2pKI7UAa50SRv/dumJGufI4
0HvioroCMD4Cqgc9NBcTupDLR90p/PQDb/SzmkXJUP7yLm4SIME0QpzQLEPyPFJK3hgOho59iZX/
MBv5p0/XDblJHokDTK9B7Sfsa2KH0FRzRdH7boDmizughf+eXQjkareSGME1xiPKGh4HONKCxNVM
YWFzfxcxtkKudGKPlbIYhs+2HRHNkLgef6vnDQUwggavA8lXdbQoqpTHSKiAv8thtxu5vsqU59XO
uxvh4I8Hm1Ha+PUhT7ss+Dhh1x6uwALJ5Ky3opYhzz+1K9g9kupze+Z0EdoIikRQDDysFUfOfuTF
YvRpwaezOGYhgzf2DzcCpCo9eKKJdsl0AaYFtbKy3au3XEHwhfEJXdJT9jxKegFYxZoMED3Eqxic
fNWfEAjN9U8Q6OCVizOzOi2nL/MqtE6SKd4N85zpye0qEgTFiuuR+SgjCx2VsXyl0wRDOiQVbt0R
3nzK3em+1zLEEROFUNUDvFNaaP0CxSOJvNu+xVd4hPPu7SlEhUx7beJjjJQyEYNhyWga8E78P+QG
FJ1ZvUBr9lRLXkytBFLwWJzMgG/awaxHyeczJlADG5WeEpMXzhL+QYAow7L2WlSdawLJx2YSrU5k
6rB+RQ+lsd9VoiNEF56VzRyikPOt+HgHmmJJvcUdr3oU1BzDJZ+W4yoSSvtHfXPSoz2mNztDAi8e
W0PCt2lrJ8PaNSGPHC9JRJAXbiArQsW76XiqpLK0ls2x7GU8hqVbL82TnEg+J3ZzVo9NEZZQHl0q
zW1HpmZMnSCjDUyghb20HvxwmJrD2Tw4Cd1/Q8IrLOr7yykUEETj02rCWUAFP7uRee099fB5eciQ
VYIwqRGof1ko2X4mIb8dnbwpuRP+34qFuGbFUD+R+yROLgaIAmkSwC/EHO6U6lbbP5yO0/DIinCk
eQkg7SUf5KIW5lNG9bwNSlr+EHLvp7aKoP4KArBmNAXwfsod5oH8SjGyI8uMi7O6Y8ETuDq23Xrx
vXEAjxJcWcIxeRIMYJIr2PEgmmGd7IdoDjPRVHqbq7+o/HC0snlS9NctEHx0X94Nkmp0q6i+8oZq
zYnAnYxwMBdm/7Q+h984e2Zbbozszf1FduW4LTVndi517FDGUo58hzXY+aGKywyiCtFSOKXOoF1E
w2xS8PqSKHPNsJJLxnbHsoF4bIi5Pn80xlnJkISZJ9SM2/kfp6NZ5akscC8qCEVwa2bit08muPfJ
9rgkBtUxl71v2R2V+Y6mzS4WPIgrQmQhHPRyLyKr8qBl0/hxDaW4Xaw0AaHRXKPan5L3PV4jqUmY
MTCguenUKk3Eusmeb21pDYMqWp2RAhGVxOIOgl+AE343vfm/xZytA4G2rwbOqMKA3CTxpcWgRbgM
sRCwbCmvIALcn3OHfBaQG8CO/vUYiZrU0eM9nq5Iit2z4rZlm3h0+u84vUzQ1UoYGtBC7Ceu1zE6
1F1mChFAFs1eSA0XMHTinMuWUlHa1+LFqbL/no2QtIi4cLS5o7WEST4R0/ZwGnqBND5kPSYbEwF6
zgrWe+W2ffJoUjrz0D/BVEpeudqeHLVedLW4v4gW9dcDo5Ccpdap4sOKzcWO3SbHbyfTMmEOqHU+
Zh80jYwI2SOX6GVn1XETKAkZ2VgxrjTS23xn7rsJRp6U9lt6FULFr524Vjh3EtbRckDOB68302fK
TeNG1Myqb7nIpUUTkTQ06+pLJZclbcqOcnRxWZRjifyTMfGuTEt5FvlHX0gZpzyDXV3+6l1SSaka
Ea8UXPKv2t+V7yNOyM5kEC7+6Ph/wmB0PRTCDV6L9PKzqeb2M04uJi2toW2hxOujB135BA+LPJJQ
3fdhLD9NXxV6ojTrjuaFPOWZOOvX7pl+1v6D8H5MopJRbVahzLx+LdyeTww466tfiWaT+8HLz6vk
VFgZcLonZoNbRApWKkAhnBwfaqEU2UYhYJTp+MvYFWCYryl9XiOAPepxoPT2HfmsjppPyuWw6+hw
4/ZpE1XUuXq5HmJ376PCojuvc4z5n6T5XfhfOy5Gz/EETVk92WMuQLlz/1VEprXcCyCEvXl3fDWt
dxpiol/LwsBUhijiAjr4uF2PpdoMvsTAI1cL2TSQCfpV8S4tjBE2xjPlP1pT9nzbccJdcRQkSUVz
MJzhxhXImxzpaMHUyoA1FDG2E5Pjx1ADZNHLdBnQNYnIk/oezy3OdHfeikOWZz0YRIdgxwQaZSF5
BCNgAnBIZ48YO2yCCga3KOycLdVLVHwfRmqZqazSlwPpOvrh9042N1uLcnLU7WysXCqP4jT9TXCj
ETopLf8rHd5hKTk7oip4fS97ZF0xXVOTPGoLh0BHKgDcGFX/heYtcwDgZpgXmqMBVOmydtpNA3zn
j3TYvZy38w+HJXG41oO5DBTtSCW3GnKMbAT9dEdOd+O9HVpDKe1skdd2gkzyEYchjibVKkItHaky
X4B5KD6F13D/wNwB9E0nV9rIIDe9jpFr8oF9/VGOv26rc4ZaoQ1rhM6Ra72XBRPchQaUGwrqqbgu
/2849aFo+0vMLcD+dpZeZQcfZek4hBF5TDrQ9tlzCQCvnZkXGBIU9w++LK+SE1CqGSAQHWkPhmnm
Dj6+WGhhQiVx5urkSRV9PUTICBaQVY2zuK+NGXvJ1ypw90g9pNQsMiOWFSNSwV2q7+/6fJ/iJm7y
sK5aPPKgeo999uHwlCCkPSwRFbIpcBaOP8Ai+pKBLomb0TPUtFnpbG8tnPG2xTvtzSgSWEq6Agc7
rvpfF8LdccDSagSA/NZoRHSZaDRIJmWbY/IS6A1UfCKcDYOfDCUyNqhU1pDiEw8M1pQ8RvwIJZAg
KMmAIM9lisYpMSqkQ+2M93+BVSZSlOJ/oAGmEp1ag7Zxd4/8ivWzrUepG9Oa0OmBvEtTcfmTmNuE
UfQgvXUjzXs4CQnpkNvSc6/kuMyqi6x6r6ozDH29Y4m7l4A+VPYW01+9H00mzeMUdr9hBsLrPUTF
G83VyI6R01UvyS5KWdX7rbX9YHcPYhdgnYsTWCqFlkjRnylGd2/Uv0r5nB82Sh6dwwZEs+jfYq6K
QdH9xZGrO9SyiHIDGYJFnhN8VcL46a5XZSeSKGwgvCuj0Ve0kpCObiDy8caYFpbDFB2eaET1Od65
8LEUBX2ZT9Q3g6y88gfDomkc4USdpTgaI87Wv4HLzX58WXks9iRAU1O4O1xUe93rl1pfo+p13H4C
zMq4MWesDNE1SotIPPe2eFljonrhcid3gLOlcJU4o9XUvugR14By+q27hyAMZJU9CYqHGL0GMM3J
ILKcphO+4OFz16AB/TZAN1Qjsxv5ivMTEEPy8vWMXvZotaISfYND2oHvTumRbA0FAtVmbE41GFTQ
g9bEKeKBgAb9DnsBCfE8XapBtjwLZrBF86RBH+ndvToHp+CH8Zidv9voTRxL3I+qujWTrwjxZ0uU
Zwvm9/XpicPKQkTmrIqa1w5Bfmw6Y7LsWNds9o9fAdrfAFzWST1xx8YSyj0xaVmd0LKkxWEdhSH8
vQXeVW/JPCOuu7wI4FNGEgiJNKqcz6JwrmvOvJGYCrf4cAH4YGjJMUkJtOo//jCag+2+puZizxee
l4jlL81ADIv374fqfraaVaTKYgf2lKPcTEIP1C8F4cKYOI8vxGljMpESOmIYQM1+R6jSuH9DipzD
U5PJ9zb7a25k0E56McXp9MNGGdSLIblswL3jIkh2F6/t+XKzmGVZ/530mAWiGELn4fmO7731Zqtm
0lVixmwxgGY3fWfOPybSNXj0w3MsdKMWjFDl0Vvye0D2a4wDMfuPQ43TTnUJVkbrnvEdP21z9vHn
LlV1B1zsW63x0RQFkDCcMzgN3shFLVhM3VgQXjW0dnWGgZx4vIuJ+vr65vAguWnZ06RlwvZU5w3e
44N3sFbeiQTtt6pC/bPh8pw3sclI8uFR8bdW+4uqUQ+w98SXi+IfjiCZ4ZAxJ71ZhxXLJnUsG3hd
R1KytLf5wcg0ADg1/fuZ+vO8JBEak6WeBRtAFSCWxggBn7h/G86M3+GzenDIwk95u4FUIyfpw7PJ
7k8kqNczmwc7ycPZ/x/xVDdov+AEKvArsLqszduz5nVJLHLlM7xXxiZf+Tsw2mMabZ65OClYmAb+
QwUn8yl4nLz2Trys8PQyoqxAGLtWvFgLZaNRDoVSzUlSEY59rZtTxbQGmxswR3kKcyDpk7RChWkj
TIPmGf6TCynJsyjGXvzJb0gVeBcaOAQQKcahE8axAolVI6a8BHQzH4UllEdDnTecK1HKbdgRvgzb
nd5aYLqde+u2YyDqJryOHk6EFmbQrwcyMnQ2cdPNxzmfO2Vc+J4vXXCNq4r1F/BjxAGxXT9laXMS
HEmEU9O2KecL9Lue03jCF8Fq2NvHVk2QLteFw634DJ5RAfY4Sxi3aLuU8cmrSoeQtESo+zT+mcWq
lJdAMs6S5RumkHniy0mpTNEmm+fLMTk8ygnrn//5rkXmClSvfggLdYrximH3/CUud83NyYyOakcc
hyp2tqiDeOZCaQ4RJQQqMEmu3IkvIX4WLMQGmqECzXlVwG5GxKG77++LBstzQclRlYh2AKMfwp7l
GSazvxskgY0JsjrOhfCnnJXRTRODskKdMcwWVjMH6NA+auaL6l/28iUv4E6mRN3ftpaClyDATvuD
da7ykIriYEy3N78BcyiOM2IZ/fz717IvaZS5/7PMGkbHCHBA5Yj4oHUhctI0wYGR5EUrC0Q2jcat
fmkX3+JgszAd3xjZpxtFWpCslt1YT0Ir8xkb3Pnv7idOeeuWmFGYCHx7FvpccU/bXy+OkOWuAApc
uAMVDRz9zLK+bgdydHf3EMFKV+l+DTTnf6HF19C7sdU5lQOIddYyUF1M96xchpqHsLJs7rodUBDt
7S0Wdp0xeHoxh0q6mgYYuvH1xGw85Zu5c3l36yH4Vq70XPm01JSnGHaZiXYpNKlTVwD8ZHiZpN7+
sfBsuLB/TtQgxFicLafCUJPCERxyUVWSFAmY3yQFqq5xf/jrX4/hfOX2ChmkmnHfFafLHp78TQjX
6aBVzZ5y0uxB4b3OCNsCv2f58uEE/m3aljS7Vsz4fYlXT/gDJ9f0ziqOIiV4EoONjzlW7Nncr1Om
VV0bhMmIsirbgnQ7RAR2jf6IdjiUY0aGCy+hojegejfkFf7nsBimOoAS8RNK0hDNi049R9lUbn4C
g0tbY6+StWjBF8eWO/jrN7uNGd/WJx619dXRjPJZplDAZRm231m+jeyK2oKRGZXvHzZFkpByF4dz
Qno9i5zir44x12+eAiR0suA9bNL+6I9d1iqOwHfOAxIVzUzsH8Y6vYQ6BBnX7oxBiYWeKyhifJrb
9RZeuF32/f3eaW4eigNH/6vEtHpd7zhDsF2++0JGmgn8NDSHC7UztA4KGpe5GE9hz2iEI3c/rZDv
DId1Z1qVaicby4sDPEAIIHLNLHSVvtSpdDqzSB4/cyJOtcaHx1fUaW8f5jVOvQIOsgQZhl7VPftB
8ZJpFfF1kEHPTSiRaXEmm8/Np3HL5WltaHwc3WJM3Y/vJMqHDmo+vSXqfMjz/Jy8SQHmZVnGvppM
RyTIsueGALYJSmH9NPfD5mfQItm9Cn9Nsb2OmNgtyzWc1IrNSLxj0JQRz9q1nBp+z5P7f9nj+H44
rnYYo0FSgjmOQWrvS1ElTuCTv9ER40MBiyUivzQ9f+0NaTiEI/gmNRSNXvtHA9NI3VlmSf9hbz9n
1AVAS83IB/ABVU9rDfDVDt5vvp5RDC74dtKR+/CuZzS0aNlpRLYYfjVk4FXanU+PEHCqA3A22uXr
QT/DRp2e8iFD4c3YSoGF7QvDQR8+L1YitnWc5v2dtVWvTEcYYKJsr6BFbiyIk5iab6weJwfYkqnD
W3C34e8QhSV+cUJvJXhFVuoZ4E5D8NmNwsuY71V9S/15EGy2tRWtup41856UBV/96pNoRBYECyqP
fBbPk+mhCWWe9q8v/fN2ZRgzEfbeeH9pGmWs7OYPTw0uYys/jr64EUkm9pJ1HnTMDg+ub1ONo/+2
uue6GmIYXDcviBpKSSEKxmtm207O2xa0akjCL9NsJgHRxg0RX+JB3i4012FhfgbGfBD694UOGYxN
6YSwcy10En+mL2Ag1fWEU8lq95dm5KBmFYz6pSYyrM4564RZ3W2tlvJINjRu2Dysw5fK/DGRbw64
vUSUHpGjSIC4TfJ9qYwzlbOcRr82YB6L9AR3F9/LwrLu0L8flc29JfKsEHIs3EUlL9A7hdPlOyPi
V4asgXpTxBDBCXzoYqeK5RNNhwsLZeKOQN4jyPkNuddOBlBqh9Zwiwew2VtuA/sj9sajA0W7bjL4
cGCLcTji1lvOj1ltShMNX5FNetoCuJ6A12H7Qf9C2IuOHLTWXFkCmr3z/o/ulTRz0QS4jtKxT2xA
pJqsPG11/czognUaR/EOUV3CV4/tt2M5WYXNf0b5Ihj9K/3ia7yzOSHILrNIARxRv7+rpJb1btwQ
WFqEKBas9u+lc0CJd/6WBLFCTg0aGzckcfa9Qc7SqbpEhJhMA6+T5LcWMcQI1qxDUSl3/S/kbfRP
JHPklhW91pLNgLlBlDboQILaPUNCjaNTNEdxOMkcy5d5fVlt4FoRjH5ugBkbo5ypk+vmZU8lwfDZ
DquxhQ0S/CMIM4CE0hZid0rHca3hEtzI3AOvpN8k/h6iNdkxUgOznCASGMYL6xVXdb4gq0QVNSdC
XgNP6VH+f72PSSdtmT70OsH0viag5ZXz7hYW/w/ifs96zTKdZfd4Zyu0MWJRLocunKXNnNA2bfyf
R9/L0dT95PtJtzeU4YVxuR2xY0yxVDsO2XKBtELnnEmXYPBd3LiV4EMEJbBidWCc82uU7JS/HIi9
nVpSZYSniOgiLFvj3B60pByMIAZKo6eeGHIDcWsVbkyZ+G0DBv4+AjAJ5P0fLw+6cWU4EXagVcoq
a/JTFULvaH0zemTEMm6edMoxMLM+r5F/Oz+E32pUQaeOb6uiFEFQQx5K1wqCvmYMJrUMsO6fr5XZ
hgpq53EK6+u0hCQNERQupujZ8c5JGgbPw1sHn38PoyqoBOMspdM/qcaTsBiFlDHhI/Ve4WQp9JDG
tXJygiO/+RI/gqXdWNDv44wfk1HFtmHKcgDJ1GjKCoEB/KmfBWadBGo9+WOk2WMuNLEluov3D36f
eS42Q/PEoXrS+Z8DS/hj5wDxhCHrlldVsA3vPE0G7BN8nSmAnwAjEO3KGXvnONklArSkEA5OWs5C
vLkzDaWbQultqMeR8V0iBGxqp1ku6cYotwJc8WZ8XF8IxM472mP+6J4xZe3HDRX85UuIbiSiuuoc
UQ8cxYWjrp68m5ixoRpafgxssMWSYAy+KJYnLhGjpL94x1UzqM1AQDqy0Myg1S95RColLjSvv1fc
ui/g5lQQIvtEGMj91bwHWDaDoZrXu2k+gJPM8KuK36RRuILWT9aX0APHzjUsGjpMCJS+7Y/MlFwF
QJ1kaDuvwx7AeqrXNZSCY/BtEqLmcnUjGL1G1nDExMWgobT882X685hDXw3hDIuwRxrXvjS7kTQw
vPqOyEoD0UIBFm9p48BJTo5/mnpNo4sXe82ntau8vsvF3IGS+rC+Nfv0NSUodDtXnPYKnxwf316n
/+buHscKWRO2hbhVP4RmGX0bIrhUtsZzG9ymZdDRjTqMs/0rDdmN70/lQll4cfiQbj2MHLgtrYgZ
kGeOs+7KzDiZaelzzfxxdrbMePVDoosF2yCJtuq5wf7hf1e0rzUB9+ssZoRO/bzFW/aSeuks/ZTM
Tl9FW4kCmM27xOVLM6hxGa1naRwZDWvsndUek2lGXwGziYXDiYsHKPpel/q8nZlDURRdgkZ/uvDO
IIPk5f703Q6tPsl/+tqOnCOY/3GcyGDo5CkV1LVKTzlp2oCeTtNPyxjGu4/o8k9w6EJGkJGJmzvO
xjeWq1PZ8++1AZzXtJA5qtJQgu29wWGs84UwwRTmD8B4QyJVEsJgOWbVGbOYx13WDh/Vsd//OkTD
6xjWBd0rr04OSWyiB68xUJUg4eJMa+whUfLlMcQWXDQ7JWm9N9iXtNB5bnvkZ0UAGJQ479nFK0AK
DltmhWMDEKh3kJL48YaOE8Zj23AFA6DujCQ3NvUUoUmSO99ZM5WwkWd2eWPrpgA6JGS5eEgFBygm
Llez5U12/D2P/rIa8m0T5eqyVXCRM+srFvrL4DXVxnQzpC5pNqcMyHnDTLblUYpb6UYEAS4qjPwL
2cGX8RUlPxDQXcGl6cJ7KEOqIn6KNQ+kN4FQbrDteSuWyYWDRRdS7/tFUNrzfnXJzk5MqzL19Jww
Je5Y0JnKv7/fBvKjfsPeDg5TjH9ZpiCJYqscGdz6rm2r5IaGcWbBiwrSgn/NFVu+0+NYtXdGUcvC
yGLXNTE8O1zWoE2E7O/2V8hcVxeLb3CdVHiYx/t5yHQzqg5omIufvOeVj7MO7soOISFLCtgj9t6f
lj2leERoJt+cQWBjJqxf9aBkF2+EC9piMT8KW9TPGQdLyh5HL1SMMZsFWW7NoAwBP+/hk3NBKqYb
50nnBJZQJtZuDCyWkCPngSknjOC9rwziVy1qbxOCRPsz1XRPB1/lTpUYP3aI+crzoO202zqERCaW
6zdIA1uFPQNusF/Q6GaOb/dMYA9WSjWx+qEM8nHCjaDeqZ7fkXeU/E8gccMAmbOMh3JMz6wh/XM1
VQKS6DRx34FBUpLakKurPUNgiTpqRzJSP0Qb4twmrBXNSNbByZC4kVtMhohdEgUl23H8D1OM5QDy
nv1Y5lyIKZoPM5cjFNaAUD9I7ejN8+L06/z5qi9ka7Egfpc+zZq28EeVtmRJ9js4DL/HEGpVybDj
KdfMdLsg12AGrJT3spiivePkYE6dLBK0x7xaV9lD/y6O0SKo4MBD5O3MMXcXar2uSAwb0faeI/eW
8l3RWmsIDaszRurJqaumEWHUvAViCqH6gJUixUDy2WpD2gr7IUti26yoTYHOhM/dFUOA+PjsUdNB
QPCen1HpQviBbJaWDmEpLeG3XH0ZA+sg95i7Tn0ebVdNfCujYAifToJiulL/hbFGKjSfafqm/C4D
ZMx4vyh1vCE1tv2CuP0LlAfH3K57GO5r/2kxQVFd1m8z6mkCckZge7g/DhtsttNYeigx9UztdbKP
HvTc/6kpCI9qEfQO8jTWDxgIHvPLNjj/OQalAZ33sn8ZdG56rAdoQQVWczudD7UHPw69ul/I5/9y
uygypfD0unwmAaI1nswW6s3VXIfIt155F3J3b8QnhNrmlI2DGlI/nLxhl8iDVJSeV7udc4WxBk59
IOgAv5hgU8lyYnSTNv22ZHCKJcBIBkEYUfZhDKLW3EW39I69sCz6khJjFOtOVPYjJVnzHH1iZDlP
kIeNKd+DmaBqpiGIx/5pSSqIpNW6jmXvXHDRdPtkVaf+qxbOWsUfyienxFAeFy89s2M5Q7Z6haxY
qOKPZVZNWvmAOyBumqHvI8qlizQ+VOJ4UR/f7OBapB5fuMo6XZVhBK6CYHWLrYfEZdN4zB45ICQ0
txO4UqwHdYAB4PElLfoVWDfJCIx0hVY37bGPXR+BOTeEYj0E8Aj+jCPSXdJGQD6U8ZbL3u3x3pWC
/O+ldErgOzzxLDr3toUGHqdmKTMZCIGp9ue4iOTZhcf5hWWPuKaBVJuXAM52cya0htLPg/mNrcpf
0zbdhchPuqH3JQkjcoxWedY3kskkSnOIK6jARfDqSAsFv9RHYGnj5irzuL+FU0Lx7wTrrSQ/3AVF
Zccyl1Myr5e5pLKmCGzgk+Nq7yPIBOePXO/yAh90fmeYzpC7QAQE+nPm+zdqfIEHs9LlkmvHo5cM
f/8a5ayFaYV9kS9/DMrrfO0GLcax6tQ78iC/Cxp6kANGvowTOKGXs4CHXD7ue84N/NUby+xKAW9l
v9ktQmjzQCboidgLzm78ivxzh/9MiJ0w2R9IOXfvPD9wVxLUl22efbz7Ig7UxSmuF6krX5MuX3A4
lYZbqvzXJmkVJk7WSlDk26FjVQ5mW8Z2QEH1sBcWZ7RdodZfY+kkvYNhv6+BeF9a63YA0fkAJRos
oFoN90mutvhbfW5nYAPt/XnmAYx1hMBlrsd0JdTK9UPWwXG1NuW23454rMiTXXP08JuTZAUAvOGt
SGiPPYUX/tC6Zy1EQ0f6DOznH4NZUgrhnMhAufz/ZpT1zHzLYHIbW3kYRDa0o/dcon9kDfdkBUYP
LY3pj8oS/A5rMt9Z/ISRLdi0VhDYc+gDVDy+Hnu8hLF/U+oKUh+AJZ3csmLhnoDyrVIsT/PexGXZ
16o7lAPRKZUvUu6UkdiQRbo0CPUpWHMbfZCAooSuDEAHcBQcUI1aMRDXQ4utP7tPpMrP84O7+VcO
9CFppcOCAaSi+puGix0CC3tuUkhrgceknva7QrWUQVvqyFI80Gs817FYM5FxTuf+vwLp0WwG9+b+
6TH1MrpjpEqSUCRqthpKsiGYXkkEloikVHTc1a/bpRA9ZOISWPx3+cUS4HcStafrBNAwmrRq8yf1
99v4DGntJUTGymPF/CFMXwQM1U363dItLmzhQGjxdn5YTSEfIlOoNMOWnDlSV6Nf4AKli2CtQI+4
FWRWBZfTNhA02ad4a8o+mkCSSBCFmkl72heYliFE1uFw5qF0u/PF2kaZfR3buyLMgQoJ8PeHkiPZ
WaILP3+V1P5yb01DVnvODVYjXkfFBkVx+EdSCOE1DR3frFnciiZhjXUysG0gNXLwMdptGder38LK
gbsAooGywHMsRMBlWHycDUX7gSWMD2/Sx8Eymh6VF7Yz3mvejJZhbAZUd5fKMaYG0nuNYQSqgP2S
PX0ktvjt6BDHEPDobbpCx91DUiKj88blEveq7nWWBgG4FSBLPqe+9hwV/bWx6RCl7/Z/x6VlH8t2
IczY3UhyLrQflOAG3g9Jz4SUmkeONXSfxoFUUqfryvG5AGpG6VtrCvR69kuYgPJTXQBcvatCsPJD
8ZPNsB3y/bu4SnKscZRS0VQ1wDS55ORR+A+CrJsKnP0YrwL2kgDGzJ19dlBMuIOZMCzNTBO3NFnE
wG68QXJqefaTrlimxAUnozXkWhYrywtFlWNehFcSc+yHpo6tim2duCLJSx+UST1YEMAMSkAQNFca
Q/fUhWcs+ERett2j2pv+gzSgljayCpWKxvnSdBKmLCdTuLS8tP2a/5T0RcqpXjJenTFiur6AEfDl
dRbBrb8m/oHmPyfgBwGrd5EQfNIl1nEEiMQS/ODz5Lb+uPHlRXz6Gg8fIKNQbKFIjXGSmk+3M7K/
GDGs3yhm/hGl/cDT8vQE88ATvjbOeav5ZZbtqO++jnmr2kRJC4PAuYXztfYJiZUCBrsrBSgsp0W3
psfb7hXVr6STvXxn7OzTtRT6X2B5V4DLdy/AHQ0x1/tzOMeL9gBhZfyjkn+1T2+wsafyaWgABbDi
98rZpc+P/mrCCj+flwMRLckw2FkMQXucrnLn3WP0+EkbdtOdvrILaQ2qgdbbdT9wuTnZjJjCynsQ
IbAkLTwxLjRRyJ6ae/yPNMZV65yQORRAaSlqMCscX3414EN/H/CT5lvQS/4iHI9DSWXRGodLkxeD
6JL01AajJFv96pJvwuc0L4GY6Sz47cboDg6xlxJht3mEXpi1EALwBmrLluLsJcCXYiSx1Jy/s/sf
+i+Fa/ALHt2enQW3DUQKksBJO3LtucSCKYJARaKnhdKZVUELQkvDKDCvrl07BCLuuB3bFN6pS7io
v/Ry5oMjOpWUuoWeFLNcvntaNgExjdSiroXqIhUQvj8uZqMgXH+xcvOs3P9aRYqVDSnc9YM9K9XZ
Ej6X9vuK6MDLks5M9o4/ZW12b95ReKiFoZbPoblTt7q9hlinE3rHAZKxzAPlYiSbwZidyyQ4aI2V
20UjOBPmD8TLzvZm4EO9lJ4nmV+xFG1Y8ko8pXXOB4vj54VwNZ9ScCkIt4QvpSgUvyX9H3S7S0iG
3Bu6jstmdwbjacGLNnlM4bykzReGco+AuV3Ul5cRxH+Auc5dMmJCiQ9nl4BJesHlEofD4PF0ndid
hL0bimTJG0XLUBnP2rrPKZv16g3uXXno11bZ+m4SBo7a9lR9WCWwHxoJh3GqBYSZsiJ7XL6WlH/w
jYih/qfUWpoTjF4TGsqNqZTrcOOhHZdAWlP7YwKmFiXFZGQpALlf9OtFBmtOv4MhqPyssLVSzYTC
LghdQF7aJ/iBDqHmZuOoN5t0ryn6GGky3GLP6yCnUlrzNw+m1KjaGlNJ4EE6+giW0/+ChQ6uX0w6
4zIC9r0KHuByvOaCiVvpWHqB7ou2m2XVvDp1cmcZqvve7hxRbhNKE869ZSvoKrfJRENxcAGI5p69
HfS7TVg8WphC7a2b+9iBY/g0zFQJ+ezEDXNEfFxE4lVypIV04jaRRQLNZcROXTg96cwmeUEJxhcJ
r9XC+EZG9ogh+GxVSOSUy364crlfGTbg9bpJaWB4YgQSwiAeNZKFVOkCwG6JBl3YMrsoPc5qlVfc
uKW+qV1nIuDsfdh1uVH6OL5GirQ3XiEeCMLrEAxsUQTD6j1251m3irQg/OqavK1f716KAtIRZWtA
KabWV6UEhPuSrIGrbh+3VRilRRB5tGeVTeJKNiSCR6heX0mDVUm+cE7feT6ChH2zmTv2nX/ZB5uG
hCpuo4PC8ASon+wUSyYtaoLn597OiiP8mv6L2YaYOHg2f/Z/NqMsjD2Prs6fdHUwF1Gk3iJkjIhz
Ba+QTA3i0zVsEei+6gveTnOjUuvTSqB/WBk+iWfWHC3Bq5b3mDV3kj4t6kQozkHkZi8EGmXj3yhD
69jR2kjnCX0lgJ6HW8DEqoqDNAbBLp19aAArCxzLnxD0mTWRDqXZlHnCvYEzPS/98ZqyaYmo19M3
I/FTS47BCakeYo3dNjBAlaBt0+WnWS8qb0eMrYHSOxNdf3Q2h1M0QW6YSOpKC+qt2wbneKviy926
BsbhBYXh8V/ZxB5jSGnJbtMyb6DJER6bn0/anOLzxplFLqJLmAFXmDcpJUbkzk1ENUBfq+3FDoeQ
3dQyI4hzvK/qwJ4nuISRWWQOwWP+FFjaqeh1yID03Hlm3A1x/flHmX9bbvheSDmprXmVur6acrj8
6bXOI4Z4F0maEWN7lsK9FgaUjvbLn2//j49DIpeqKnijscNEbo6x0O8HwL44xiIHGQtBGwHHywu3
n2gfkQKVx37wj0lvvwQg6TKN7ph5YaihuqUAapL7ANiiLKI64DNXHw1OuzGZEsaIzB/hi2tju4ZF
zDFC2H+wgmQW4T5D3lSIwAYwAgAoKcIxzQm5DQbucJ17eXEsNwxbqlbfF37y1tOpi0IWTIacC3NG
QO2PA595XzorJWAwpdRR5723PPR5L9iluutVbN719Om7CnJIEQSf7dHKOt7esOV3/KmWY57Bzw8d
B69/UggO/3/vbOzXC7YPgKPQALgtiWw3KEM1H786ClAwmGK1xbHE98rwdGcYzVcL3a54SJpTsyjz
al0BlVG54nPkDjnNMHj+8yKhekn5QGzxR9E8qsBlhu1SL3IyDdQkXylXbGWBRY+vjy051LfbfTZQ
XXtsElAMrCasYrh5pCRgQa+6FUZFpBWUMjTG94d2AhWIRvbh2CkcgBlNGVVkIo+PEMNh0MEB1pi0
eHUqy+wgn3eGhv2ThfSxMPOjbeszHIlsKnNF+xO9sc3WMQjGJIAd2Lj150Im8ao4sXeEFkte3edq
yZF64suu9hdzM6bY5llVJ9WoB1VZ3gWVq1lWpQ0sr3AHOk6fdOEKBHACMmYz3pMI+znWhu97Ipmf
Numkxs/vnSxFch1a1k0tUOaVL37OHhornQkZyJzn0cF58U9PVhhQjk+GpWif4AdMa8LqcvG5J0sP
PIDNWl8hQ+KTgKaXKx/BcCH3aO41XZRnRhzPC4QJVw30obYggQscEGdZ5BKuqiolyfub63lGu21c
godz/7QzlWw3g853rLf3g5cMAbqgyduRwFIcjhzbHNp2HFrlq6vmB5ihejHitT8pE6CCvwLznx0v
v3+emj1ooTgET6SZSzrm+/5BiN27WVhHRQUlxQk5Wf0HCItfSHRv/TDJr0nAij1W9stTXOmhGwEE
O4vLdhQ39w9SoxKxN8qdpH1w6vNrI3LdnD64y9n39LQrwVivwlq5ZMfuIgbb1fUE/qnC7nu6yj2C
2tTQaBNPOUk1JtjKno3s9Y07OafgB8UExWQor5p4G3j/qpsQUjLGXTTt64CL7BJRajVetnsolP30
tGr+HZn5v647vJc5+kwSrnAvTRtxf4ChSslUl9HYcoWIkLax9UrFK1DhF48+VYA/hCABQDRtlJ53
UCxdyJcQBc/hDBh0/5H022z4SNtdfeGYnH83S8kL+MPEtaBCzV7xO7TmOIUPBbj2wq0kBfaUw5/R
QtS2xX47GZacYoScu8HS7QDtSTd8eYjBhVz+c4fD2zpCh5Ruj4CtFyaa5pIOzqrBDAI2bDE1VhiN
TZXzDsIuPIbRkVMRFGeaz/t72nbRgprkRa1dOKoKM+Hn2ebRItbAFevAIgqqIVUsYlt+e6G6emwQ
qJIUDVzyL+evrP52EcCUHdaZC3qQuX2FGOoPdSw0zcNuXfN0hayX8S69H4qYsxokELpppNKzcB9z
ddTltap/OENoLqNSj4iIRgafV3eAsWzIyLoONakiSEYuXL6cnpIplwUpH8bubB9ywuJCZ312kHpr
V6EqSSvtscaaIOhbHvwO2yXej7IagAIYVNhzL8jzZhD48TR86r2lUyZ1JtV+foKqKCBqOPY7GAgw
87qnv9bKd/2gXlvuwx526+Ca5OKNEz4U9OwQ4lniOh2oAQVkpOmI6Rh99puVdK8yPrQhAmz5j2+G
dC/9ZwdyKziLAGFyiMR4gU1imeRNIXhOjRCOidftUi9DJYwhDfnNNLPMxicKyjRe7pQcTV29AAle
yUIjVjGR9dAK6ZkMsj3JJkrtjhTv2uB5xiNkpeoiyUd7J9y9SQyLwJjMqXX1jqrInofJOntGhBGq
pxlvr8qAu/hi0NbIrlY6z2SwQx0t5aZW/cYvXvqaPa/kUpIZEXppvKX506t+nYnPd1d9lFwLyW5K
5YdzxStNqkCx7zUkK34nBL+Ba7S6z7cbG78rx2MgjRlfSnfiT5GhH0hNzxlHaSgpuOi7PFBXcdLH
KF5qbIg0MI1eKM4ds7K84lipNC/svqobyNOMA5WUYPP1kGRP/qJVqw9neOHzM1ViT4JJ3/MGI+Xw
mI/txfrfEkngQLidSXeLGNDHHHpCm2b/JH+I5PDFJNzJXeyG1cLMTRDwM7CJndsnw9TePpx5pX/1
rZnB5DpPp5QC/jwMq838yRLTv0w5Wc0MQ0IUaIQ6lFBxaccr8xC6sp9LrQGbAIWR69zUcwn04FQg
hbiK42WqQggFjVJhqWoe9ymoSZKLlK6c1ftAHMjodezP9PbqTrIF/AxvXYilTFhe9NezwQXpXWrQ
B9sI7ji8IBaY1+314u6H5SmmmbUO8nowL4CRGvBIUsRl8Koc425HMaB6h9unIRp5vjsY0JcjjGm4
JzuBeRRK4rLxBTo6yJOuD7ZbtlX3G2bZV1uRwAQ6FJWgafShTUnqIy8BM8Xsvg4AmbtJz2aWCHrC
Xdd+2ZuKPUJYmaK2xOwFtF9Ilwqcb16dB9ETVlH7n3jGkUdw392GfmDPqkfl+jb+FvIdVNrfMgMs
KEoFg6Tlugx+TgobpxYDglJ3PX26dHqm4MXzP2DtphTbDvzSfRKonO+1c/kQ8756jhV6BZWPIa/A
aOtonp9dRzcHc9Db1/P3hYeYpTZgscSkUuyCF5joRicswoFzouUj5giHdh3ykpF1aOV1Gc8FzlFU
TfLWnXznOK8K+2abdI5rEGt+uiyVTOnVR857+fqJ0XruQHLImpfA5m3EYqAmXeq8bnQ3iJX3/nVy
5BX+HjArxiXKO9WMgKu2j/FpOm4H+cpQRwC9QUbqkjon6p2+Esaa4dRFWAfpnjMC22Vvsh5iox9J
u19G5si+Hqa8OBzf1Tj47NZAop9VkA/87xfbeQStaqIMEWuqU0l2KLwKEMaJGQwz6XzSmzn3tmhZ
4vuhCTWGsjQnsIVK13t9qgT4v6IvjsJH7YSWfJuKHvBqLV4/R6QjWv6e7RW+Tsjrk1bnQyVI/LmI
gE1/ltoTtu3b5ZUIVdyDi78vwRjT0E/Px101/FOYTHNbilqRhOT8USsfA59ek0unDKwmsmPvFx8e
5eDe4Lt2YSfNKXUwMGWosipkL39XQ6qTRZdsIJB7XPGOhAwLyzZces7xMOCubloOyKh3Zb/jMDfy
xFcyH6ne++Gx5Y83A4uvh0+4ZJrL+jf4iBJNzhJ40EOocgu5NJo/baJQYPRPXfLt4R7+dRNFhSu2
9DNKImsYQAbcPPgYvSTw0ePdUNnDu3w3vKO5aR1oe9u+DdZFVpNWsSw0cZu2sQTIR66zivfybFqp
sXTOpZGB3GS8t6pCX0IBIygVKI0DXXUHVao+eajLRkaguDE4oBzLx5Apk0TnydpnkD/hiZEtBcYj
h5sOJeNVmz68K+kHiGEU3J/YIiQP/C5XjcJjH2rN2AEy7BIRuDGWrr1sVSLnOxh4hBeXWavd3QBM
MBIMK97QTIRSoVDK/Cg09D0RnIWt/ImBka7eNX/RdjGzeKLFnIMU8mydG1iRDxDlhNLtYU2m1TFS
CvvizE7VrKbDsxKZaBOQfsn0P9/+6RK7UyNwIxKFseRyTzilEJhewE9atnUfuwaltXyWW4E89xPZ
90r8ydbT0DuljRid36N99oz/hgM4PrTSZVswgDlwRVrwDKTFclrQou4PpGSTLGlZr4gKUYBnt4/y
mkPaf5LLPL5CXnZfOv+cELFEUwR5hXsAZA/NJm7E16R1Nu7BZ1eL0OlczyPo4emSZr6jwDAca432
rZdNXuveDuD+lhMqFf3RGbbjsyOPaNO74tDCJcO+TVs6356jLQi15kCwRAPAWc0xtY1h/xCns0Pr
vCyUSA/dgkgI0vyYiAeu4/NKzpkKzrm3sb9U1SDLQDS2TRgRXflPDk7CLimLt4bn6fOX+DqRcGJE
d7EipOZbMEXQ3cLlovicQ+YuprzFtW6cwX+T7BTj7a+jJ2N2o3MK+OzmYIU1sdaXeZ90F+E5fmq/
gn8Y9ANVMy2NPGwLN41c27qZwhlAD0LCrK/F8bfWOfsHiX4/RlWYrKjOvD6QBKXdW41Td8OV5JT/
KKl+cFTfYYEwFa3sOLByNkoCwspyUwgqswTVMBiYdL5iWxbl5F3NmBoHorVbcHq+GYNELpQt6r8R
oo0VTBZw9xGLTDPFuzwxc2ZXSxlOAfaj7EpU/+byszMrF8PAxQpAVZXZL2NgV44abSyQ3JISNBv2
FGOaJZ38UBzM+1D36FQnF5wfPaGBDGhz299QSxDBn/WOdPdzYf1w8EOEM/cDWmgtyx/btXaMnSPx
vxdMuYX2Nba+Mzdy6alsLQPKbjbJ9I2/wKuP7F5ngqk+NBC5Ieisdy8QSV2fXNTPOAUm9Qup85IB
q7zKtWQB3i9Qb7/SB9BdsMpBMlW9v+xNiGhmtIQVAfj1dvyuWC2+AOkSk7DJPKe+fBLf725mM/sS
HnbZfBZ/S8jKQZX8pQ0som/LVfmxXzr79QqN6nS6MOjDRLxMFP50kTK/j/yJ1eJkI6z7/pqY7dqO
ktGfxSvKIyqiesQngkatb5/xRGjfI+XR1ftD6zTVRtrtGdaevkqoXDyi8afkFMGE1wOf1q9ZPQ/G
OY4fLx0EVQvW3vsTlU3eZst6u8noJwtJqJIisSii7hQbV1cxC1liMKIv2RJT6vQt+GNWc1yFy1Lc
AnjCMjxV+YI6OYeThDu7ElKzJ3rwUf+pHjwqtANjhRDpKqvY4XgFsmxwIg6ujvFS/F1m4J0mJ2S5
1ijQ0yfKrIvsRx5hF4aRy/QodCAgOV/IUj+oc8Bz8cg3UmqCYnY57K3EeJmppQ4o2t92mgrjoZte
u3pBs05NUBrDFcBFoy5t+cL8X6NQyatxSHzN/aSJGMtQ62rFNZ8t2CZq3o/n/fBwZJ7aMzkMikne
UEiCOnzfHuMUGXpnplGzb2MZr/UqoOX+7OnGjsRRx+nY4GZqptHZvDKK96vR1DDE3WFyXXGBTXCF
RoWG2j9kpNLrhl+oaB9HPWPvwJ1KvNZwLgEk9/KI6ZrXHJY330tPWGStZz+8X6fdsZD7C3L8f3wX
7x/OyZ+mKmcmSt30YDhgM4TFKwzgdPCOO8z0C6kfk+O/zl1xc25m1gb89tr7le5jaDcuNk5e0ho+
wmPbe/PmgFzaYoLZjwleYuNoGdXhxZ9YiTj9LBna8ju35RY2bp6CeXBiHfXr/S8rCcGkrKWwPS+g
dHTsiHDTXP3JqzivbZYQi5XK4PYxO+QMqyaBfLuKPJG1C5CZ2FYu/uaCmVr5eDL4iVemN3oFCygg
uJ8WFrhYUkqCaOpEem0nwx2NOqy2K1+dD9VCTwZfsJngrMHLl+EItMeh8O6GojgIBmtIJ/mx/nBr
MH1suUcgOcaa+BN0psTYVKOu5w0a8Eu9XJxr3T+wZ39kXPvec1ZPV1gt4V29gNWbaeNQnkP5RadH
v9MGoFVkeBobJFXYBDPWUEHI4GwEdQaLAtBKAlD5afIN55kw6qdCByh7nKGMoChBSGLkmmuGo+Kc
CzHdoAb2r1RD7CVQqMd51EC+K6IYt14KHBK3jK1Nyuw4G7TKWskk8IXUXKVylknvkQj67vgLHWUE
xmBPk40x6vxWrmhNhInnJvGZR4vg9P4zre8VqKfJgMoy+tKW/nYMRdhZsSzek/DGdooResf/NDJO
ECV64QCDY+8RjgbqbXUicw9hAhM15kOoC4+RpA7hPVOBYFf+hPFOD4yz7gCLPMznqbl50uF1mcyx
f0tPLd0blfU81lPd4+fM+Ak/tpsoh6HohJi6lCq5MuPSsj3DOzkq+2iA3DKcwZb01DvjpmyZvQLD
qGGy9SrO/fBhtrASR/yL/gljrhCOaoqdEqzlW1k5MPM+ZtpDDN5hZwzYhjoLxQHZ4exyTdFdaxgj
1JjArTyei/CyBAqs1XrRL+Cr0F+SauF0sP4lABCBDra2o1cME3ZGPT23xeisqBsrUyLikQWWIVwu
erV7/5zNMLdhekh8qyqrCbp9ZtO6RF+tlkeVSoAIu30cJv826KasLSDjhB909m4bSYMCt7DV5Jhd
5miiRPYN0lr32xnu1bwxKHRTpCmyWxTZpFIx1f79pXNpDSN8MCvBjOOP3xENx4Nkj6GFOS1YQswS
vIVE+uGY7kYdb8bqnyC3X37J29tCJ0AbVJYtL3R1Kp4l4hHraV5qmp4vQo9rgwuD2jBhCEGuTOGN
xROukZyKoUcj9mrhLTPmJfV7GUU1RJhue++dIdDsOM6LAq2UUyRSt8OG+jH7PJBJyAl6d+86cWba
/YMe3gFDtHolwVAN7aEnNXg4NzeomSU4EVyhrmo2uSJ72u3zDNgKZFqO5PSwsqZPkndmeDgEFkfB
9/tid1mIOYZiuY91Ky9FhxTWYclSiInZYPCNswUQcLKbTn65PAEaM3StlgQu+WiUWmNAPHp7GgeJ
VXzWxtOHXvKpApuxqB7JW9tqrJ7GYoxAnHkeA+ARUTGRlTqq04vphtxtsxmce/kaCQ62l6ucR29n
t5Jqm6+acqwCp6jGRZC8SAF8jYXxJ/6o8Xn+v9ka+t6jCKQXH9w3s/P8Kf0gSnhXkgmPUER8cTeJ
WhdBpONIjpFK7LNjbcRBycQSrnd9+lPjOUqJQHM3NvjQz8b9VZf/fClIwELk4eAb9H1gqW0KN7Mg
+nRltqeGRnCKNjsc/GN7p7HFTvDky7ANp9z7Z1OMnDkZ2Y/+R1YkAAxeb0PLGcHy9dQHa1GJt9Tl
yiQ32VvoIh4bkT8hDDqvpupcTUSiocKnciRs6JI8gLh6NelS0gaxJSAhuDjbeL9vW1yQCgJsEqb9
h7OHZcYuFmYwTkujSJiVjaoo1Wz23By2pIXFaj0k5e8LCzOHDQm/lGlr8Ll3W3w9dggI9SW7QzBX
iMOZl/ONzbaU+6Gs37zuox+knEMr/tkw6LOWN+eNFNSlxAW4xT9y9gTEnd8PdwyohK+go2cWSpg9
D8u2IDaVUVWiiZ47gBRRXvswT7VItDLRFLft01Ul7hFYpGMYqC6XaPOgcJ19+YTeO6ohqoz+C67M
tb6zoGrNi9vQwU+TleZrKWfkttqFT7FuPbp+Q6SCs3oyi7WrWOdoI+0JAFDY5yycdbGzlMlWN2qq
Xab5zDS/xCAnvTIXM0I5ZgV8Bhnl3Bt+mCJrmlNKf2zlbyL45DOawQWu73jVm4bwXxkGtHB4gdhh
JS0ZUc+sJLm73+CIklxHO3xRzwIrBEGHv78cyyDtGDmT8+eWJUuJwP/uLmoRH3mudAGQFkmADONS
jRciC8tYmlKN8mvWBqPiRP4HLVjcQJxnrMbWeqkC5dj2HItjM58YZmGQQAQf8mS17D2oOqvrc4Gx
8pU+EeUOThIlkVjFwYejlL8ZdNHcd9zc8utHFGYFRZ6uKUOwLcIYXSMjoRyTfwOubr6zP3tLhbEp
SfVPCbehrRfhTlfdbjNuxX/fvB0qnzwGsyeo7epGUQVmPEQSTuXSwZ/MiwahE1dsviS4S1ZTSg9I
Sw9PoGKl6e0fvpLb3WQcwwFvWGfbmuAz3nns42KR1jQd2R+lVu+iPJHRJLHtyj+5NqP1fJR5AvFu
6uG73k2Tvvibwp4n80SUXhdEpqP082zfe85wMBdrVAO28SAfDsMbvQ9a1xxq1GvYV8xzXdGYQgxX
mCBlLATgDMcA64CbHuSWyUUeelaHpGDgH0ktugoWYNtxAq6gUe9Vrhue0E/pVeZljiLhdBNKUxVu
U8wUoqLxfoP1E8UtVSHo8w/HtbHE8LRbxde86UCM9ldDBoK7zMkwbwzpkkzYgpfbwnXJIU7ejG6E
geBmN5yifRJzcJz9Qa41W7WjBDfNiLdE/UaOD0woLzSnF4d2VbmS5JwRPBMzlf5dImppEcnFm6ga
dxUuE0qOGuXQ4N9jTrZcBps1t5PYLP5miyEm0c3+2+IoZAv9basnDKr+akh/PYfEOWR5UaEDHaHt
shXcPkLx/TsGLKRE3055HvCEhhuOd3KY2U4LYXXz7jG6dSSXqXJPeKBIlz4iPDohPFO1dju3gjtH
DVsUfBR/zvUzLnqYHOzY1A6+72le9/EX6s+VHiq6kWKvVBTw81O5tLeZcUzSBIfI+SnwdsGtr+jX
IEUw1+b4mLAnj4h++KVxQMJNdbAmPbrX+oofvqfuLz15Z6V3TRoltvIjiwnmf0kVZlgc6JS1A3+8
3XYu9bugufRrN8ZPnUXwu15xIzMTP/WCTW1hDPW3+/OYwmXcocFT0xz4A+6lq8APiH/6J4/+mLGg
ut+HuHNGsSRIAzBksyZOw440g28rbZ7oPwwTtD9KZPtlD1tXP8khWJ11j2D4U3tz9pRZdfqbpQIf
loZPF4e5hmzS2o5AUTwuXwHf5zi0GFqDHg2WCIfjCAQOe1RCi3YNY+7tN+zhgZiWfs9klQnnIfsE
nQgIjicQAPJlNr5vbgGMk5q4L4r4uW/H8fIeBe7hIpBwW/rIoY6O5QqeoyVsWkc9jytSDdgy24si
4iMNxkYEKllEglHJJK7kLiEbUsf10u57+qmjQdSsOXTrKoSmPhAtVxVqrrN+4062UxzMwkzzolbg
1y9DqHxRw6ln3gzDJMWhX5prTd4NYe+klfqdDYH/WT0kFQDe6QGm8sx4QyFiOnvQ4ccPcPCdlaRr
oW/OOVJQszfly8ry50a3e+bHEIXnUCF0Nfv75xndafMnoS5IN6TsHJKJq7z8Eo44AyST4M8BDTRi
lQ/X6zzXdpyZ0kdRbfCidYpt86dO2f0FDAnP688rhQuWmdcib/tRoX4WbeHuoRqjL1p9VXKRdpSV
oebp8TuK4Aq43+te96snpl28lRxRjBAXmGDTCfOUTLUNv6iQIpx+mnbC+3+AkrDhZ4zGCJybIHDI
Cf8ESCrEFeraVrYW0UT1AKGwFjuK79cJ7EA/zzDQawe0+VdIzDHpzEmzoZtDDBuhgLjbHdeppPTQ
RoWCxeLW1lKl1w/0wsEEztP16955GAKMh4S1va1wUAdZEbek+JoIF7n7oQ0OyGc+cB9TN2xqkymo
0I47kQSUOFjcUEVw5FRrWwBuYJ6Mg1gUkMoS70QPB5D6aTlAllj2olBLogYyn6QOSpUqNlfoL9lv
afE+wQ3qBFcpdUREydpzm3jqKzqh9utjDxERpl6skUaH/cGgPniLNdgPCvFbXEHPgFwfkfMmiu+8
U/4vVO8YjDVjZGH4RFX3u4pOXB0MXXVYT24PXDPRiN/nXicZpY08aboq/rbvd935M8UrekxbCS5C
DNQI+7hYeC70DX/VipKQ6GaICt/cMTFrlAPjLjwxI9Y5cnm6dS1DKT489IC516SaAHZwIuo4o8MG
UR2X1XvikuPcSQn1waHI5q6OM1lYFqIRyqZRNx+gaJFrk8mK/mnHYOyiAJyRuZhP1r0r49g2brIA
i/pj6WBQCARApQBoPIixML9/6LfIe2Yrt/1eLS7E8oaR3r9YZ5cq2m4wLyp6yOUzekSNILlVP+Zc
CAir6cpx//P3gPs5xk+jF2TUhWDxX6S6ffbiQNbxPh7g0fjad0jg4dtuCgTuv63ANItMYE/jjf0n
svcj7GpHmY18Hga9FQ+46UyFRhlpnieTL0PlQONxKLOA8R+3f1v5QnNc6vzWBF0SsPbAWgxK4HNR
b45fPD9u9tivhC4cG+QoKPqky23CJ9M1Mpi93i93+O+jsF5RYctQfHshgSwJK5GkUk4opUMJ5tSS
KqAM3Vmn9M/TwWc++ovoPXevXiPPJ/+8dCUWWQreC8VOFlBlio9AKylkrvAq2XiKjc9BPe2Fiujd
bPqKY+KM4VbC9Oatz8YpJaKPCU/ovGY6YV1k9oG5YOwEQjHbucftVt9P7yOb1zNa10aWoIR8+W0e
xVBR6cKhusylLLmHxtx5uIvTG1puBpzY96wE/B3jk38L7AP4OIFnCVEm3Gx5AKl8miKX7T9SRAUS
KZBjmhGer9Sv9Mnb+85pjqaKNrr+89UZW/7lkPmgs+AIBJxTevgMSiK1PYmXFmUMTRyzxbUryAsk
Ysq/ms8x3pRBZHV3rLSwpWhLiEuHHaIjY4fXiT+VofNokz+7Ms7XNKsRSVBaBtCUbx5bnVEtJKBx
vtJ4YC1PPJpzKBZ0s75rS5I/0esFTQiFP5o07ltZLJnWYrY/6AKEzDfzmes/pIgENw6icA9789B9
G+m6LW7sD5CLoOXmt/MNwRoY+kn+mw/xI9vyJ7rFxzvt/Y+GBYbQ6MCXDThm5TGkfsqjwl9r7hQe
iwhAtHnY8KdqgkS1S3ZYShLYQw6M7i5WFczE1ZDASHp6xvc57QypfYl+QBO6L2pJbPEJflRSpPIS
QA168oT+tBjloYfWQYCgHG/C+hBkiqUP64HhRyYWIOMoZeJhaWwXCoZXJy3bS68srlWhL6lVqKIX
ELa8itZB094mA/Dyi5nqbnrQ5YzeMwtKDZ1A7HC7MUjuOiZFzsCJbqrI9diRBZfpwcEEkEhv/1KI
Z021HqKbCD+Em4IxaEwBH8WZJNBSQSgRdrUU46GeQ7RzHJ3N5SMNURDO7dhaQKRKHPdIIuE5ZNCM
XyrNCNHiVtvTZC/U1gBjoU3dYPYNfBQ6g9glp/aD7wJdKTref1bF/hpM1q39Xw+8MjvQBa46Aw1y
IsldJ/MyBagw9jlpOvwP9RMXdjbVRfUdJKmAFBjgDWeEZJdyePVe7v4xvz6qOsL/gFb3pucDitVr
DXhbQ9hcuARAuSh2KedDH80O62zKC1KGnwL8oXWf//oe8gdOJKDQ+HDQFPUC+w2zjQR0sjng+E6V
0Oo5MAZ5IvnoHY8sIf0x+bSDL8GQDVN9mm9hd/IGudZe+54N46dc/7YqyCur2La/q0UXhpryhob9
1yHXLlNoxZ1s56wgTdA8fYhkrMtxXHYCGVvrhOL6s2h2MXklEIxaeTV8DAeyUkwNRsLJ2YAjx4Zc
YdLklxNt0cANJZ0q9O30txwe5ZO+/fxL7v76IGOs9qgHcJUWLowWzjFJ1rUHgKux3GjFH9OULahz
5JqtIbcuEQleKetSHw9JcL0ZN/2r9Zvjc1djR5Jxupj0+DZ9ZZtBeFpLMzxoMbWhqDZj3oM3Bc+l
a8JxA+py7JATpRSa2kLUr4gZzWUmKybh1mLYa8bu5jTwQ0iElEq4q6DKPKsX+ylnm39JotE5Bcuk
mHlWJr+kGfTPAcQR7fkuEUdtePKaCPNOyI8Y637+ZJC3dieLtfntCexaZbmFVSt+creE8TfkBlOo
wlISvPiLn/ozauTHnW0niVTzDlVxj5jCE8O09xCOGK5fL7kf1ibKueVokbEaV3/FxO8NS8LAVA91
nJaHUHhYxvkfmGYuVPIfMJ+9D3IoY7YtisXHQK69cKCCF8JsdK8fVt4EHi38Lxf+9QRgw4T70hSf
Av8em2M6wqgHR2gub3v5I90LUpE+iLsJecmlUg+bnfiKpR8bDaTqmOlpEAVfzs/UriX5LrZqh9E6
PsiJC2eEA3c2i6sOQj9daBe3JYisPpIsmk7UmXWM7rzuBKBDtJL+ShQmVuRG0Jex99YuTnU++Ziz
ozgK1++/Q817frvMjDfiw16JshiR+MpphJlc/rweG2Bb1e4gfHLUkBuxj0aEXQpJeWX2H6Q4LPjI
cPbHA1UPaQiiOS7vFxQQI/SpWzfIfkYgLN6ePfawd86Y77tJiEIXBKzYaYjxY3dDalaik20P1+yp
oDP7mXkQPT65i/OcwG+OV4X8CJ8P9P2/xq6nFtavIb5S4XgIH6VMW4r9Vo6FpzVauDLTPoYIFRMN
7tp/5OQC6UV36F3kyxHMbsjWmd1HwW2n4ybS/88zv1se65CRrQltb4q1940v/PUaRulcPzFfh1yB
3Jg18mIMqSp72YGBMzFBrjm0AxiifXqIK+r02IvCLAt4nOAcZNwS8/SkB7xO1zy+AKaLlRhA8sfa
3IjRwwSwCWL8JvfC5/koOQrcSAzX2nNOTR/7Vo0mcUdAg8ge99xqkWb844LqlpGsIEACiaqbOLJr
i4lQoyt/2Hm6Mo0vjJg8Ls2oikpulCmDhBWterTNtKuKE0oykx3MPE3IQ3u5u35WYnCjtIQfIX9K
J6jaBYnLoiMtAVXZT1lpU8i2w91PgqRc5z+UBGCvreOIwUBi8MKW3Mu9y01dxl8KSSzlnwo+Hv71
EKXtRb9KW8qMNsfs31nab0EfE4ylEtMzn4TPHoI/Qle+MyyC1VU9p1l76cu13QqCPbwXST1onSff
MVqoLQlFT/tlbs7mdDRIW+iWGpOW2Egqssf/aBgD0RUKhF4B8OibGWrYtKNZCI3ijRf1w+tELXUW
nIUPeYyE1dBSs6I6x6QhSJhZ7rEKEhVBFRk1LyGN2fKhIEfKoHpD8KW8wdIVY78zUg0zev+dHkR0
YvEQ1MRmT54K5ZvvXynOkwyAPZ8gIVLpIUYBBQ9XGYhQQSEN69rmFXVJPUuvhmUy2q8rlJOCsDmx
LMoQ87edHmuIS5jt7Y5kARktC2q7Etgp8FMib0XFX4+8cvCgXBJzo6wCS5nNvbNLKJS4sYGdZ7uv
BiFBBkDhC7mPZC5l2fjCJNWw9eMTSU64xqPYE6JGu8zn1HBNq3WwwpMxEj4r3jo9ui87NUrz49WV
lfNbwuvXHUVQy5yUwzZCnEDUhWRc2I7Y2BGePQ0p016DQypyytQ/d2J92Ogl7nLzDlbyLxDW1PkE
tqEGF8vV2Fu0xf69dmsBlI4CWFWrgNJOpXuxs7sbb5LbRzDXNVY54cqfcRR9pBOVQOkfJojcRArt
BFxml/j+9IFQ9tvR0eZkb4h6pxbgipRELH3v6EQyhmZ7kKsQk5irEFuNQxFaYEzPJYEEWKnfZSnr
gYcMGBuB8B67/s7S9B7eX5tyzOJsGeGA/Q+qnFOHfpPwhdjr1+TrrBFK0fdJ1pnzxAC1nZ3qkt69
P/Enf68LOk8+fZozvX7JDWb3p/ZUonqqelxbVpfOnbTViYKyPXc/U9fHk16DGzAb2FpeLXiDG5cQ
z/Ar2jv0hFMJg8N5GMOsoXY0aRv6KFmFpgmZ0KaDvzQHQ3yauAhtAQ61l38Q0WXVU4l7mRQ4k1OL
M2wel9eqLwb3guJTSC7KUirG4aw8p5Repr3jw/2WGcvcLReaByjV2Ae2Rfr6mIDAJxp/qB4Bu0gJ
i4v3wpbw0PUv8d+Aj2zUG1syLRaGxWybgYJvwr3MMHzJRKwuVijjf3ngPe7VHo9RNqZ1pa9Z9ZgI
W/QRBW3DfOqOCGaAaX3zKPqmDl+iFSaN2Yp0y+c4uOVoZdXVhmNSgrX4Jn+bbLlklJ/ykVXMZk4B
V9bQjudqwBhra08kUe3ja77S/QY0qqHYR0Jl43kNZCP0SH5PaXtzeDnMW9NVxDtyJxHEV+TDtCVE
6i94s04h2YfiDpTIiMUohXztKm1D5FuuySl2iC0I/t/6Ua+rMYgCMUcBsynMwXnenJjYCcsdlu6x
4tIv9iWkkJRMqGFAw7LBtjaNx5RLiiO+Nk1wDHJiLsOUZNqfeaAXbXOflvzlvyVFUOODB7K6v0yx
OKBYvRUL9FIFMgvm3rqObErxqi5SCl4gZ28U5ZOmWa3wjB6GhibWcwA9exiOdQqxh/wh7TTaPAKD
qHk01SkvBL/E1zdIbkdMjlW1R/Z+dRohry50743oIiiGI5t/8KvW+EXlLfDBvi3LxFflLoClPuVY
CkAifDHGWRxSW32hEHyCM4MKmWd/A4Pqo/t99FKVFKGLwCHZp5OZoyHM6JNEVZAMSVKfq9NKEej+
1TEyN2Jcvy3xI06gKyzPo2WOFYEEq58uRu1dNfNYmkqxTlnOjHh4p8PEkHKY6BodhNM+ks4AmENS
bYPZ5eWu/8HYrSsQQss8Tw7FsTuO1eGgRTduw1zire3EjtrifYs53Z/C9HNFDVuUkqEzgHAHliif
AroBsapYMtabXOVcIK2DSrQgBOTHMyNfokrFVAIvuKUDRkg6qR2/LxxsCgFBwkj8wabcmhC2RN8N
v1fyrQwoa+ycTFopqzoegraTInXAd4Fbaiw/Ll3ERMM+FjD1RS06pXLGbW79B4n2psuNpfjD8HZM
N+ax14qgP1ghBrROiJQJ5uYayLaNUpQuD1OrDjeNH4N42mOxS5tLSMSmJtArn36VWtGZDe4z2Ott
+A2CS63BItOCka8lrrIR8ZOTYO8SR+YgishlNSVG20PM8Pncx7fU/FUURVYbrcSnYNf6Jhb7aFtI
cp0oUmseZwZurY6VpQOpa/QgMIMM4rGvCm3IRWMz787DU9BJYy9O8m/Oe83TWbS7sZaW6r4zHIij
jntlvTlz2QIe3kDGl1Edt59IwBf8n+5dU9gQeJgUoGRnrEwBHk+k0rlqpwngmxVsSkDcCBSk91XS
IDr3KcG1e6sRkplJHy/yp+3bGdaBAam7gHO2rDefyNwn8RklwhyUWSXhECXANeXRRx22MsZrS7TA
lSb53di6IB1W4CV3ZPRiEjh6Z3P516eXWRVqVcmiKPM8EORLso26stgTicHjJMa0BF3vUOThYowW
HOWgoNJ76Yh7QL+VQfjFVHy7Fqo0d49RuxZ7kN+TE9FU3MDwtNzsGMfDQUYpaMqW67htpw1VLnx+
2cUiRtNgL4p4UVb8Lj6nN4kjpLRygWV8+jgt6yi6QakId+liuR3T2NAKaLHhAeku+jLI3pJ/BzEt
8md+rq+tOxAyimaPYqAtMbt1nsPyORmKBnI/X0L2Z2xDEKU0q00X9gxGhtYhHrVxOye3D4TCbA9d
awDJRgBdxrdgaYRWJnRSV+84qZ8dTpnkGgaRzNgFOqrgEUqzYdtD5A0k85J8M8Vl4fWpdIdXWgJp
lIYCSNfV7k6EZZRm8TNO0uFxGwAfhgggpF3v3dZ1CcHc8VYb5Xku867UnVbVj+2hVWJerL/BBqf3
dRa3Gk5GBceRdy8SZQRUcw8ArXm4TewfiRov5xzEaJWZQgPR7oBJIlGVEx7uMrRQE10kpJAJ9Bjh
y694GYNCmZRowi6+i7yl/sVDOPhNVGp+WjYmGQSjinanehqjAR8s6uHKlQQ5jhrm2WDXbXCnhDNs
P9sF9IMEJX8EG2MYoU8SRsLxBjo2cpL9iETRomm+zj0chHfOt5opYXZYXoYuHMGbD/oOk12LtXuU
bCviVZg4YEDX70q+EHs0UXbnfBR62Wx5H7yu5vN5wGuF+JWS8j5jcntcQkGPp0ais9O7vne7m8js
YI9N445Ikp6KoCnQkKiG+ixq2IhyK7+EqRrXOunN1Y2gDQr+2VYNuxCzvBHdXf1LY3nKlZyxWPaP
1wc//d0+L3t4K2NWQb3vF3e5fd5cjmYLcoYeFhRy5tJNJbl7DTqCmeVz5tVZhYpTUT2NdzvsURUI
k6dBHaCqoURxS/kQVg7VpcICgVvDCoiqV5iHOHbPmpP7V6mMsGmRJ0c3Yv+G4gWeimIwskyYbMri
JPFIqEA50mgt/W16Xjq4sowA2GNl2LWS3TU1/zH6dMNDHiaZrR2hpvy4GvlGyPApWjhoN6Gl6sls
b/FV3QUMtO1vYtXML7L2pJxqbQbO2fTsnUO7K0VtvSw9HhgmbpskaIA18l+A+XfAjbVbW45cEGL0
QIvkI7v+Ko+jFii101Ty96123vuIZvuPUrhRbwCOofovotZdHPNP0cuH91yqtGbwK5D+pyxNTAFp
YjXLR4r9WR8o42Mx/AIcWXLarXkrk7BFy3Uu+BJSZI8JC3U9OfEqKuUUlRzkFuutulmOLLLb9yKg
qid6ZKYJFn1wL+MJ9Zd/Zphn14yhkqhHT19kvWsaMHmfPFnLZM0cvewulSbdDgfBzAkze83GeSQ1
vIvkEdFMsTUvxm21CJ+3TYJ6QE/He4YEGZ/zk/5xdzAKhiz/kMmTJ3QyrP4I75Hc8uauI6Jjn18T
p3VwuIYyyT1Skoo9v7BgpSHgqHm13U80eyUn6qQ/3HmPvYR+2R2WlndGrdO9TVbiBcRZrPflB/1x
4sLncmE66bYXhNfNUfWJQgjtDcx2BocLFrHbW9iE8oxZSTQiTCYKMez7W3EbBleXhGDez3MFKhlK
gs+sDwRXUslheMhxvgblpjVrLhILR6uITVMLYFOWWptt+Haotrj3zYjV3+OOY6gDV7DYbkvK28v7
yDOuZTSIahI+DEBEqG3kWwTscz2T5jhoEB0MYyDW3yj5Ct8ulqDNOgTM7WLXWUNombx1rladlsfj
zJm8GvpvQDoDOH5ysJANFwtdI1qDsXOWf1gGJ7yzPiAbrdccy5Qve+/0J7UyORHZEmmP83em6PLt
m6PXuypmK292XUfnQQu1IFDJcERFyXTLSoy7SdARkKsgblC5xcjyl+S9X+T6byuSh+xM+rdlXbqJ
XiN9ffw/028mYVAGPX24G54ZtK5W1QRVFTs1uAgowXfGjHfi9UqQaoOUk1eJe1ie/BKmyBJ9PXOj
prIjo8KOyBZSiQg66OPHdAEPjoSTQeCbfo7Yytx88Zao/bnHA04l+awVryF8o0k+fk5kxQTzM4dp
gTZZedpILtGGkpfc7zrWIY0Tx8caK4iasA0tXHO2QoXMYvQ6bYw6AbQo3IOyYQg6qMt7iw+Y6xEJ
jgPnbzQaFAaTfpi3a36N7fNJdt4fQ4v1J4dQpx5RVD63S8zJtcAMU6NKNEoJRorB4BX2feCGsUA7
3h+rsp8wu2CGWAK6WLphMdgRuRoMgsqn2CzOQuRaz39WRZyc5d9Fwk45Oy3YTLWBt3UL7Q/lOGRH
PEWefsHOXpahoqpTuzBzRgMo7GiVkIkm1mwAnVG9sxZbQmKVmfK+Zd7RKx7ZQm5lYxO6WVqGbDtz
gop6DdZUbVU2GZJOKEn8PPX755wRpN0NvZjSUnFvx3J7RYf750407qVkXCQqZCzZMM4staa+tFKo
hfOWmRzRuu/02FV1ie8HOhUhtrKhTb0MKW8XquVQrSQgyyigzAMJ3vAfUCZ3+rDU4mZogxcg1brK
EFeCeJIEgWh5N2jUrFrdk3LCy73ZdzcWT8L1ISoOIU+jVNZBJ2nYj5eYaFiNNItgEjaNuqoQKZ94
OL3DkX5PpPcY+B1fMABxKKOl4TBhNp+IkO8KHj8EvBcni86vTl0U5UbL/C1fVNqoQMHAk8FbHslp
yz3lXbPuEFd2LA+0UlQTKJJY+GzSMjD265P2r185G3E32u0UQFh0y4WwyCnEePN6hu8qmLIPez6r
LQaOtsI9Xw84T+akMRVXSkfIohbryQS4RUpFaV2WeNDUI+r6hcJVlsVxmX6s0+HxxTXpUigJT5tp
SElrVEuxV0lCeGdYBwoAurJ78n5Mnx8eFVVjJ94nuj+irrJT1g9iCVM1JEpfyG4xAhFrsiJHVkmp
XnrCutgldGnCFB2Msn1qmMH9Pv7uekWOTNWGKEQaV/Mq5R3uD8mSPG6RATLBFOG6Wna3f50KEqey
aUSQs9zDp3jYSKbzSqYdcGP7ve7Yo9MoaGj0cmww5FZSl+9zscK/UgwLqzfiFsjOtVXK97SCG18M
gvf3oYR/sJStYD0weT7ErCRLnalTEZUyGYd4pjrP0pmftk8gZmwRYJePARV5mN5B7PpKAVMkXDiX
amb7R2J1TXNCG7tcGknYcYwZGWkzFUlaqg0taYbiW2B/IxKhvaWhIDqIYpD3d3RGHtZgG6vvWXIV
e8PtWf1WbGlkF3yDm19p25uyQUieLWLO76rmIZd3N0dQJdNUhO5pFxqqFd2awPsKv7bTIxBEbb5s
VCIIYdEU4KFOXBUX3YHq7HOF4XY2+nCWkkU5srzfUcwoRWuEPHpKdPy9rYZCPQ4hp4zyA+5D0CeB
tSg2n0cSwrtlMCfpfNi5KRRkq/tkCZauU6mACcARp2O+veifS8Weu1Ci4jHxYwMEaGnYLDUITazm
DMmcDkGJM6RcjfsUN9yyd/2l+UHVKP88H0NXJnzwZzxuc2meWkCd/L0WzXhT/rT/27rO8a1meI9X
EC4JOhR+lA7YgE0VAmoRig/5NgvzkTaHsuCvOI4kYnPqqMkTygY/oNS2QaNKNJBEhlIHypFg+XZ9
2+41ASqb7Xxr2OR9W/d/RBi970DM4IQpV+dVdFmq1slH3ScNkYWa+y5lTMS3M1gewQTPGEqa5qGn
eGj0KKlEihz0OUpT8E1cTkjgIbSemCu818pKadCjdP6DfTMwh7ZDUZQjTqodHgPD/oT44UlIOqJg
BoqipiQ/3GWn3+mCbaf9ohGmyBtbsenyuE+nR/jLDgXn+GogkZQsjlXGOqw39xgp7SQDxVNL6UsP
1bd7yCJAq96iGs0Rh0gDQpC1nLV33bEQ0L5DmN4Z5HsXwlSsVzoqSeoqKwMc+2UEa7E3rz1Oqlqr
O9cgFjgdvL7fUl8utMrpUiL3BCjkfc31G6w43akDEbZ9V06JYza1omUyqbxDVQU6g+/b3PPkldPg
Zv9InT+m0Hs7gGMCSNRaLnZORTn8bc3USW7WifHzfy3iciEbZkaAkSx5gBT4xjfawYLvbcltp00N
uIsQH4EACWkPkZnFFeL9vJ/xOIDUuCoS8H/NK/PMa9htXrPwYdcbloaG4rsqIxlyRy5ePvX3Ao5q
+Va4wskZRJp0yz6rNMkwgQISA/nhzs8LzqfH5YujJcOUgOqpEyHYZJe1G8W0wwlnQEYC9sGZY5a7
38CPViqF4OzSNQZKlB3ugEDM87fWn6vwpXZRyjDTaIBjXx8Gje6qCsATdc4D5pRG5EmrzsT6NnHB
tCxTh33BpsXDNWwkqegVi82htneX0hCqBEIf/A7elfOCej5YvHxSdqm4zYRdEqkYYt9Y+vqo2BRv
Q6Ysd9qF4tOb/+oxlCQItBvXEdXl1aqWq3wsjNGsEo4NrQxPY0bA9z+6MiOVGY6lW44vWvlZgK7o
QilawvPLrB1Ubc9wQbXZxza6rjnvlOR+KdAHvllpxNMGtG5343TepTYt9IIgmas7wJcBgGws4v/j
zO5+I3F2JXyd+qD0G1ly0MClW9ej9NarnO2tr8P9f2KZIQdeZI8rF6J7BHWvF3dwdJydWveMdoxf
q6lifpYMlmbmeUlDAhXra4WeRAkMCvet1SvBCBDeh/3uFN9sNhzJV22usKfAlggSx7tjapy1NR8U
W4oRwSdz+y/56mdGGnXmDDKDXXsDwhpBSg+hmo/LeleKXP+kK4vOzWztBRXbmLUM/ixwQpyEAqv+
e/WWpJECwKm4sZz5iNbS/QDXr3nvWOrOBdGBkY1M/xns+wNtZIdEf7Zlf1xZ9XwDV15zsMszCxCZ
bq9JYeXxniBkXfwCRSzqtEjXY1g+4beU+L3Sc6zfhvdyDZ7uW0vUAq1pDLRelcjl2sLVm05c8Qmu
JyqRJh/6X3HNFEPcvq1wG5Bi9RSJVkVftQGkYkO63QHfPb08F1hiO8I9mEXoSHh0Aq6OdQmo+4jI
D5piTMT5ULfMEcSwFrrNlAbBexq1xx5TzBtnIotuQI5r8O/w5tRi3S4fpulGrUMoCRPvDZI3Kt5n
hPE9xkyKR1iqcZKurFjyssE6VG2s0zX//R3yF3tM5nf2p8JyEoZ1TsGtlGtBv82KQaLgNIQiQ02R
Cv7Bnw+jwPB/lo5n3sqsIEFSOaxST5rHrR/crtG+u9QoFeViA9xaxCZPwGtS4g02cEmTrYaH/ZwN
M5XzwtIvPYnPIEY0R5xN4byOo8QlaF4lebB8p9KG94bZt0txVQ3xiziJ72IynfQe2tBtibX/iltL
mJICOpzJ/6tK+y6sdaOIqhKjxfI0WCe8EtNqhJzeFw7MWoMyhddGog5QxpWEdPbIA5091FwXyhUu
d0Mo/Xalo8ljFcFOB+sX9tkWm03e20+V1BN9Nvk5+SPRrQaHLa53I7XNbgNX+L5wUZVpgoL2R+gv
SP6LDNx1O+23Iuennh2T1OWOWGx/vY1lIF7+GjYoQyfT4GMeealzPQUDxQr0ilM6N6NaoXgP6Bmu
CIt1XwjYHk7mY2/L9qeQgrFNwh1ddpveVEcNgGmQAi07MCO/k5qs6ztscVxgdqwy0JLR2pemEG9F
N6ZYZ08KTSEZNc+OvBuAGCqBIXNM61EucjPtblvcLRYfMbD2pHW8VN4mBQOy0mjxjHduD1hXwhdi
aFkqWXr0uKU2nYcvRLmmV+tJsRGdqGC3nYug/+HxJ543cVBKtLRSl6+Mg5bGWczQryrFsfAx7Fj2
R9nF3VwEZuwvjeUhZZrQ5qX4tnThYKoe72Ew9kBvHd/fKzuQp9skVYVPPa3rVREKc5y6wP4fZ9s6
xTU5OhqIus+I54IU3edIO6ty2miDdwqU9bycO00HX8F2IhHwmi2J4KIkmR4LiqLYdOKEDamy8LYT
OPRR23EEYwcKNn5f1L61MUxb3EmG2r6o83fWkETzIMmmK4WcHXMzzGqwZRnYi6D6hT7xRqMdpNYq
iVY/CqcPvBKr60Pigx9bh8pnJJDKr+6S2Rk7pdc6vScxA4HBc54W1nYOkHjfz22fCbCpJ/8IDgIw
QRFCMA+o9Jk01JvhXwefwz45SbLswmnVPg16avJPkNoDiucMaTIbsDV6fvCrRxNZHisuxBkRJsAe
tmTNPNRzaTyCFFwDK1s5CNLX1Vvcc99zhamsRSeViuVHcd6BkfE7Qg6do12I/Y0nMBLcsL/elMJd
biGyFxGnRqXIyK189t2Fh6gI9dXrzot7AoUOeIw6WjyxTYjY6msylHXZJryT5PMjkGoscx/F9v+U
yx/7w7qqX5yGi6Len6p8Ez+WTVweG67xQsE3B/DdblgwA+tfAebD5BWPE5OEDdLT0ybf7WF/sl5T
9TsMpcd6HhvZlY8HWM+XHAi2ZsFtR0Uq3PtqErdMN2r3K7uYVDbXdp/32O3khgGW/5MBidjahJB2
qJPc31Q+wb5cLhnSgQVkeWXXNppGK9ZWkfyAI+WF7kEMVC32cr82GVHVyQzjYNGbySWKOlsCPFHm
7ZCS9bLY31QYc2Z5Qi5Aaq9TSiV5kPXb/mrFbeJNhH7KWAKjts9gBKrkhp5XvyCQ/k2/ZsNg8F4N
qrFCkGoLhSKZpXCeQ4ZiYteBVO1SqZTN0egWUylK4kE6EpCfVO9m08BJm3gQPEqJ+wn88s26xhUL
VTi5GxGeF9OlGKo9/YgEtGfYvEr3tO1B/b6yY9nYoZb4yj/g9BMk/bUYQwUm/uOQfgkOhu4dMd8S
LgIb16GR1x/1qtfGOTc//i0XQaoStoEfNwWZQ7yuCtBKTzk3DbjUh12GQ3LEixWQadGR66N4dgC0
KSVnoiTbBSaVXccp8aBxRQUHDc3o+1wvTHewX0xa6taGO1nfLgVtpEC7De5VqJCeazo9hmGQ28bX
2SmiGE6CLcqoDCAPJZakX+NSTeHd1JzW/0pNNxIdUGCZvxqvWJk8qWpb1CohjOSm+xgH2NMu+eV+
EIsUpkypyRgS80q8hub6FF1sl+wPOb6jX69JurJWTiJlyddt195wK/kb9TmQAtGIb6JjxGw0Aicc
7NZCBiljco0gZyuyftGV3kyXJa6xCWyk1G7jdYh+RFtLCQnJtpvaANbYU53TUjjGcvsWaqwkO4W/
2ROi5mHcyIshFGoJQHJThkWElIdFDoOoULCExpkU004gzV8LQ/swPevf3E22X6cTD1KV7EuR+tXf
9dp66GQ0xv/2BQLfB3wTGFMYCjEuGsZNFIEpuUT7BBYFgvZ+Sbe+/U3grGowGNGBarz9epOO133I
oeaiTt2ZNuSB972/vbmPigF6eIy6sXJAXj/gn3ZGAZQx9BdExLvoDLjYMG8lQyShhxiKXUX/SJRo
iy8vYKgIKqGXGpYKSuCisoWDSent/9pPkBqTO66Eiw6NfZkqSghBw0PZ6jIOTPQiTVASZx7gtLe5
Uy98YdTGlMnFJtJLDLAMfSAAidPmrjsRZPfWcopaRMcfD8OWc2GJLMDIsdzg0a/IcBgg6Im8eNY4
lEDRQRIGv6RzKedxR/uBrnGmcxAKu6gOO3pSzUcu4NwAODBhm9AL/VidrZbPddgMB/fozBeFRrAt
ApyICLQcSRmX6AQeNqESY/YKAV3DtVS0igLy8/lW9bF+ChqQ+O3gubfLQ3IeqT3j92TPUbf4Jg1p
lyBB/d5EOcH3ixnQTW1E6A9hgabvvXVrSBr1H8VzlkKlneS4GdYpnJ7x3eFZEgjqyagf6NnLVhK8
S3MsWWBsG1ze1Y5nkQVPcC1cPdJX9uMfq55uDBkccB/nR4bEMIdv+ga/wQBw0AJM6uC4tBRYMU+X
qTW43U6TquKa+sqZUxjaFinQoKl4vGttgeSpWPSQRzwjQea6uqbfHOy1bi72AsMzP98um0E0STLD
b0vgfSmzwWG7ZUb02flMzSmdQR26SeUL2nJUhl8XnqKjPDPAxon8JYhduzUgnIiDjPhToYVFf0QN
BGJWVqhDHGR4w4BSiXIyqu5EP+2gJMtn5KBLSvRvk74O/m2ZncRky226p7FFdgOSPkdw7kmn/4Ph
1rZgdzs+Bz9mDmWJcmsgjX0z/7Ul7N9jKevYeI0Tt3FyQJNKb1mzi1sXXjXAYrWfTogf4mAdRLPi
hrWZ/swoGhnCQTilWg0uyq5aMY0vtpWPKFsE8lTBHC4NG622ZWDkJ0ro+YTXHmz8YdQOiCUUIudp
sEXCbhzx+0qT69ptE/il8g+nYvTftFCQmrcr2jWQ/7gqzITOkvee0BtU/A82MzluGoArHkvtnhah
QWg8PY70EXsvhMoJPBy0g1FfHLxAEIN2NtIYecKg9aF7Cx7dYg1/W/oy/ZnacWsBfBpku3ZVXqGC
dciHUTistpuUi7ofwglwZC++yTOGMqS8D46zTcdp9c//PqyIsQXTK63UUObdEWfSQ4E5fB6o9gIe
/mYtR/scMJki7sPpvk1bzlP7pCBCcvXUCTENYF2V72prtKWxvEsfmokVpbJPm5ihg07IyyQqL2GG
5FX1bK02LI8i6TkEBCRit9Es5KfZfd8hDYCQMC8bYCqvj1NVRTD7AnzFE0GP2YqD2QguGjx5lmo0
iaR8n5AKPGlWRC18e01pviqZzF9yCeB7zj64AxknlhfPqPs/V1Gmzg+nGZu2fTSAQZi9VdIZfOR/
kcqFhqc98e/l1f+ofBTBVV7xfGAWoTlJuUKlMiTRoYq9p/jcS3mDH4mDZ0Lr0RTLTf1mZLCifWZ0
HGBLTfMGfZwdKWanKwoFsSuTUM+/PwzVKOOcSeyqohj7NdwCZiAaUFi0ssj9bd6Yksv2KNoqL2vk
Eb7dYZvfBlROJGVlG64i4wWQ18KnZ/5TIeNToSFL6+F5mV9x/42DWIZW9YyKo9bKCW65L0QmARTQ
rWkn0/ayC536V4+/MKoFmnWExQwxDkDRVnI67InMjhEA00jvwppCmpDJAhc28khS7f2zmRAELG+W
GgaHTqB10KMeEsyTreWjGvqLUBEtePAsjxhDa9E7wMpMescLkEGKpK68BzKf92BQDcQs8ZhMiQb3
4mbamO0BzJMwr/XXRTbXfAOTNbgnCb0CWyvuE3d8rrvZpD28QS5gmvkKBQVzMgPuPJk/vBssc9Ty
wEfdZMHwV0513L2SlGxnTANP3lgMJioxpgR8+yTUWdIsuUPAoAg4UzGQx/psC9Rh8191jz0Ws2rV
+TEBQKPbzLrfLydkjrKblOSRPi+2jbtLkYoQQmjLHwQUH6vn0V/snf5gX21sPVNdxsh3w2AeuyTX
4tiatsvZ9g8iLopmuBf3znDOFCU9Jv3BAL1VJeMd231IH/HaQE+rNC5bTtj91gM6GdRlUj17hGoK
SgBgeuIMkze2qK4etXpOPxeXFuID3scq/lH3tYQfCUrjby/lAdy0ItCdII/CJkdkrXmVimDHqZCq
yRx438/GQNAXUppYOcSDvbaNLQ2fsq6n9zVFOFdwHwS/9lfP2i5CDzMtMwSBvil+u3bIp+KNsbU/
0I+4Bs1rqB0837F/lqm91voQmPihQ7JZHbzi2dQHmLksffPlzCi6y8Piq6bSQl6tAXa2Rmec9j74
QO4jihkKVs6vf4vTnpetN7bShC70A8VfERluPckHSZ14FMGeGLlNdXwNe1aTyGMnmuUgmzTJPEKz
+FxIHEbsEUec4ez1pZTyVgIJ4t5Ri4HOUPCmcg3T75SA2Rzhy1zQxUd+sv2aJrZJzJl/mMC23iij
gIf2Mo97Vu22O9R41rU9vnn/cWn1iy8DL0pqv7XSw2bQRX4yQ4j1MUZnnHpEs0oi0SMAYUC4maWg
K0xkL+81UTzy1B0hOch7JK+Cac3XmN+EbngymEG6iTuZBg4396EsRdrxzBd7S9h7YUxcuCBDTbVF
AnmtIYRVfdeFJD81bjKZu8tmlAzNjDUfqEyY3884rr9tvxq3WQZ/WeM/2Xv1MpOKAf11wzMUj+z+
RbcgCFinqDXxrr4Zp3Me3zWq8HrARGOYDA0bjLqtK9ELkBB9jrhzfLYviBulwJapoEjJf2su1q5N
u9swEUjJD6XSYZjMB7ikga8OEbjDpwQrIVaNVJtPvjas48hCVI5G2BLJTV0sGrsrUQ2AhxUnBJ5m
kpxbI/6CYFEn3uGnN9uPcN8dyJS9H1plHpHd3fvtvkBizXk87iMvYEEC7iAXAe/Z3DVPTjwAFOFF
7ZjYz5L/4eUbLvGAvFzIMm73cC/dByMotUh0clgzFY9ddLtbttZSrdiBV1KD7UybHQLkYsa1nxGJ
UyDCa7NRX38mjNC4v16JWINA3L+iadKDSh/ySKUeKK56UXngZ7hjcBUQkBFeeX0y9IMyeRjNrGx6
/bKrKqJnfOSxmIqlScSqGZdjYuB/U7Dx12o+RfHbuMh4uYE1bXHVb5ZlqH087V5zPhmEgTPKqYzE
3tU1Wb9o/6aPYv7roaY/6YELU+fUYnWioecxROILL0H40xCJNgos3tWznsm2Gx5qU3obwLyBLql1
cAxbLj+8sHlFRm6nn72rKvFMpcqUDMAP5cX3bvkszVWnBhoey847Cs1Si9rg97sbBZj5Mouw0S4i
z4mmasZg/J7h3JdHmqp4vdnc7QKXNavqaWjj30kA3oooMpUOok5wR3g/dLGYgmNTTX3rNA2ojsdI
3YLs7HoWM0MixKlNXWsJqNjx/kTY/7w/KVPE8wlNK44UfK7iMCgFlUkjTS+1+II1kn0VDEMIYLgm
sSVgrNf98KliNgup1XWdSL8XSP2RXNg9V0OQiTjiSqX16lqHCZfQu6kv2zNW2YTrrNea0U94eoRY
LBQHg79YFwuUGl7BfcO6bphFmF5IoHxK1O3PEqHUI5hFq7rOJ2wHSF4OERMu1s6q6hOLz43d1D/l
voEKy9qWuu58JPXT/+i/xpLqEr+BAEM7DPZr+8hege0V51fMpJeO0+hjTIdJl1Ftm3dJ1drgJA0C
zANKXvOr8MLZE5wfzJFFbTchMsMnwj+QnX5nZAyT5HyLl3FTcgoUn+Z3sVyQFWvK+afN8Dg0vDIT
Zsmc3zTeWLaoJXhn+wpDSWiNE4XOZeF03FvGaB5gL/BT0cbIuOU/+ixNj51br3IDWnPrb7vdR5tW
SHI2ZLuYaYQLXTajuG2/G9g5zbbwo8WAp3ZQnPWyCwha4+mX5yK6itb4cLvHhuUnQq5pqEerdR00
L5L9jJCK7WZMMB3K7tY+IImCVNXoZwuCYcYP30zl59+uzbDLXzMRmT5zFmq51mPVepgAhM+NkYYe
UXMw0Orsntww3dTMWopF8KlK8K2fCn0lo+jEWm4EExeBxQ7S0M2YZiaNSpCoKVui0E/+9Czve/6M
s2I+s+TZcAGbe3qIkRzB3Ruu9gyPmV0++tsMR98tWwt1zwGRPkhDeSmIk+x9m36AhBMj709dwPd0
uvYSR+xuYM9E05JzhUKAVtzmYYt0z0Mhl8w0G5udURTMXpESDTnTdGfyTtPmAfM7PrvL5+Ksy7r9
CRJn4mctbHtIjVfOVw1BBk/bMYf/vlL86DEmpH3IjIJ6wOm7DnOXQew8vW5noWfWnHRfw+v55Mvc
aeTE6/RTsCPvgbv3ClMoQbYdMPZPVUjxLOp1N+gopbK27LSL0T+AlFxLlWdE7ouRQX1pW4UTI2xC
rMCRSyh/ESg90xDyRCQK4Pvd7ttnAN5UggTtZTD0uZw/3m5mUATWxG5K5uLAbDeYdooUS5AHY8dQ
N79kTKsVn9r1nqh0k6pY8JSNkKIaFpuLnbabzRnZDyHMaXGynz//P0OEhhRGyWbo5LbbB5vBFhbH
Uq1XaOrv3okphNPsGcN88n7e+s0uHompGeVWR9nbRudXShtCzyd31bRVQo6RO/+/pZ4/GbDXME/i
e0F6vtnjnBvoBnusIRVxVPoQsui0L79f/oUTP07+zD47iWuPWtJvbAOWlpaVS9JjaF69ExwM2ucY
mFDOmmapQ6QC3LRw26XfwmzxUAUGN5OOm6PJ73bXC/G2wt0mkFvLijtCaKVKyClNawobJstDYnae
Wbm6xXET1n2Z+1d80Al5sNksgNPutiI+eDxBZ8U79++fxWTyX3bOoMVQV8MB9BkIouAREXPAKVC1
etB+qv9LM4MdJ79Ews42fxwY7n7lDcth2eOo2DY34YVd8xzkTCUa+rL5rp2wYxYoQa1uIIs/nQi/
DE4I5HsPz6LoSmkeuBc1a0HL4SWkosKtp7qUIb4BVHJUgSeIIWlXFfkXwTl0XPSpSTppQl9mqz/j
jSh4KPQxf34ug+7Lu8jZM8199m736EjUgj4ICFPRXa/l8EjLMpy+VCpORh9y/H/n3Eo0p8vlUFn1
c27jjuZxdi2LSBtzlZovvEhJVIlFu92lAUYlPFYOj8I4pBjO9BOR1iwC7/RhpHm/tAXFskocjlOm
HNwugBYU7DcR8nzsR5j6b8QZfg/UgmdKGpfTv/IW+3zMZTwyn+qr6SIXFLDBiFeKGtTt9KotfYEC
yFWzoAyzZkizerRqy+mFN4Z2LJH6pPh8BdXjHE0mAuqZ/WUFI+8B2Ay1OCopKS+xd6PDDh/qsVgS
dYfyvC20YajqqJnkLc9EGpTEZqheER/ZQp5rpOIMnFWN6GD+J73N2POTiN4piNf6WD51wPK7O2Er
JIJVTk/+0eHQIJo46EVX5WV9VnzO+Mz9khQpXUjJw5c60P8H8FvNOyJ+WWlVbduIjY1r1WxBIDcX
IirsM9aJjuKxRZJ6nbvRSw8sjsY6OlhuC7s3OumYWH73BwOaN8IfpptgDwpo81lxJ9RQ+Hp1Sx69
hOBS0WplZH0jwVSPIGoGOopKeWDs93YjsQUX4734cE+Fq9L6P7lJaX0ZupApFChCpS59wTjOXqG6
wu9Ry4tJQ5nmtasFUWcUNc4T4fA3Meumvi5mEtG6Oq/vecr1NUDpnI33/THlgmQ8CZJYuFq/5LcR
RhDjoaO8o7uBYxANNsN6tannU0yJWjpSKCEvh/GFXJ54Xiha0JMEdAkFxSYE6UzoIwsIBKfLGeLv
MorWjuYCTD+a0vAIVMldV8nK7Ej3gKw0Uq3mahjNfaNejFnr++JjZZ2aC84DqDJo8QjBqq/VdFnh
HfMsEja0IrzB3HxyPOT951qzX/NRGeMP4FiEXzXp3NB6GdZQn5zJ+ENFniKPuGGd69nzS/Yd/M3D
NzZ/sDDQZMP7b3MI8ktHZJu1qYoKzbNK0XDgHCXFyjB8RdnDpd90Kcxurs8/IsfH5QgkeTsqtjAs
uR4glN+7/rT1Y3IsJdkKdd7x4Qkvg9uoLUZ86zOep7neuFCtfZuGvFFYMft/HeEnch40RWm8QKsk
EC/nKeMAiuNXVCUu+gqUxSDvtWtKmB38HBM2Tp5QvzyecJyMhwoCcXXG/JFQFLnEoGLpcSXlgL7N
Qzn/M7MNOnPzh61stTY+2QOixecZr+0rKlyTFA6RxQm0D9Ir1yCR0yr3zMxKLIBtfPUoPHvk4YJQ
ouizNXcGzoiyum6xITwRiDmM4CCjv4XY6HueM+XgZnr2SwjErmpfxMd6YK/ZzvDGBslxa2CUIRET
l1yLCsb2H3JbZWP7RE7RpP5Ku8reNe8Awm1smJAd8+83Ronze7OpSzCBFShWo0JwxbPWzhmcmD9c
XzJn1J+OuDjAylconSda8Efd9gNsdwUl+W2jfWJLRVBQ+/XKocaTaJzReLt+8hWmF2HLNeeYHTyg
sPqGcGVw7JfAm5girWibMGe5TOt/52Z4ijjBc45p6dmnpQXZiBFZPv7KanmElXHJDLqJCrRiU621
eol//CHylVQnQfYep6S8BQqobwJYm+4eN28/uA/k//IMqUvYF1GNyy8TXGQY9xzjXl/TUPVHq1qH
QJhcJ5kTVi9Kw6ZdmCXDWv/RTxAbjEbhxZpf6zPIx4gXb6Jz6AzWFhvyJGlW5Qj6ont+hQf1P7xL
6y8poLIN3ZsifFArrV8gQb3jPrtcKvbohgfSzA5QByx+3pWC2kTfeLXYz870DzwVwwt6tPciF0Cu
uFAMopOjDbqCX3mwRUap4WJ0qNICc6ABxZdA3U0afR0Uzw+Mlq49MBGUHSxCsSpsqYg+uCuYIa1M
y5X36D4c/I1uQCXviErTtJ8ZnX82wB0gPwluhsAIsQS+9HtssnMFZX6ARrpt/gbKTDIjCDozLF7U
s/4AMiVZ7M9q4BEuWvnP0fcw7QJXXDlQJMIBqFVpu2Mfz+tOJzrluIkXtuGGaw4aHqN7ScvGvTno
P+EAOo3LDkeEOAv7O2vlHZdbL3RkjXYXFQgVGSiOO2yzWCdQ0BWMBtvNoC2omHqa0oYRVJX77iMH
9lnb45uappC/y+Ts0XWAaG3LtbipXYV6bPiU7Hgq+lUqzEhoqmi4HKt6ZF2WI+BVR0vXpohDhAJf
zRI7wcVmZTfLcx0T44cg8zFoAOoFkn4JeVs+eVK71js7SZfz5h5dRD8aBEC/pesKJxdWXtdiH6hX
gMB8aVZwzDJB9D6wGOGrLWuySQNitGGVtGGAf1TsVrVEYJiEFBfzYNIQW/89rO21EVNyp4m8tTPs
e5BRKRs5hd3du4V5aXMCVvcSbe5/uleOSBJJJqImmWy12B6pw7Ac4R2K4LEDXK7bYdgs2V7cyAVE
Svdi3QXWPvVqmurgujHbZT/+pxdoXclH2ouUekHJ3fvHu7UKUDPwpWKC3aa0syI5N6oZ/Sd+xvrR
iyef4J1jFCmb5y5a796Qu5K3ngd3KYre1mL0A6V8poso13WbdXCbntYch1DaNtX5hEzlkclV5FFL
kApNBhK3O/7xqzCUoNqgtHR/M71Y1nSbOStbXDwH2SDl+8AZxPNpiwwNBw6Lb1kcowEE4Wk5kU9s
AntKFLubMcy2QhUZfVerR3JLA3lTx7Uhsg4N5c08X51cprOWTDUUxP3s/sm7s24mp3Cz0cEYJFp9
siAvMNg3Sj711vM8OAOCgMbGQ5hY2fAKY62NyCm1gguLjJbbg19nyQ8UULATd5Nh4ya1QidXrMsc
bfEcmG/qiAk+0ON3nCtt7x5TJZcGXQOca/uweGamHo+7qylZc4hdEd31AZLZlUmZ/yRzvVqG1Jn+
Yyu7P6+PsNz0TY/M461jSTR6Af9O42JfKu22P7U795x2vQQeSkCeSRl+ykmxRzrb5/XO22zEgrjz
Dn+SVjap8/xY/+Anqvu8+NdLSLiUddGNuj23k3ccorcao79V2e1uAoeR4sfIlbg6HFdhM2Ugcx7v
ezxnzHMTXGpfYj58CE+n6OqCoGYNceouISg9dyr5uX91Y5aekV3HpjoFF8YFdaWP5YkvovIIlVCm
kmx5kNWV7AfU/vq0KWAd009aFNDAk25hRPbhHnLsILICK4Lq2zRAEAevbn7xbTI21OV9oa6k5rhF
63gI/OmWoFUZFtHx/GGnlfr3WlS7JwdxymSK/NK7D1/o1f3Fp/h/GrpFnjrOK6akWWVKPepGiQ2Q
TKIZabHfGLo/CpANshJhUX17351bNGSVeQ49Npk8IlJYSO2lazah7X8rxLlZpPDsr8hQSp6eOpAr
DcTiXdI0e2fkVtr3Z210jTbejlR8ullaJ9IrffjFZPgYqfadCMKOCZinK3O5uCiDDkbPj4GbkByB
0OZ1aPfdAcaMp9Tl8zItkI6FRGrbwnBW8VROR54ULyEhg8mKbDOl1uZW6X5FhuGGJ+UHMrhR+uhD
EShyV57D1gttsdo9FrjfaP+vZXP1zahVtLIjkh7Ru5qxEfiUjW5NwEY3L6JWavC6PEzVIpnbcxOt
Lc5QRFA+BVWjbgGfBDF1yQTZDxw88QccqYwunNQrajDuvchCyeNS6uok+mHMTgtB35ZaPfMZlNrs
a9GXphQ+EswXPFfVq5v+yarHxczT9/1SdQNwOeNYlO76bfT7ecaiZeRgN8HShSFJwDkIlU0gbo8H
C8molNQC9Wt5JEoJv7VysKtwo+cOcWP08X19iSgYHNXSEbkTGOXZoOanKRIuQBo+kAWBA8SmTcXR
zq1hsE/A69n9jRuIWw9eith2vyCi84Cx0KBNKpcU3EhwoSiXP8j+q5AJDTnT6ghZTvFwPIrH6Crt
OJQg/8xolXwPGr2FSyHAPHtYYTHrx2Z0Q8To8AH6TeMsqQmHEruxJVbI2XPQ61GMMRMWlSuatWqD
Tjp8/77qcODO3r2Hhrr1W4bHxg6UcBG1EwRv6DZHRP+WsmE4w9giBn9VfshjPOu8m4JIouc3lt5i
+svG6bVinj8wa/19AnBw8PRbcYF2uMyRQVJyS7+nVbBYt/33zrbDzrNNw98LHMrvZP9OwTzPNV6A
r9W5tPtSvGbXZJ05yej7zWCQB1WUidvC7j7yqzsgFBeeNdHhagh3OOB5FLBkSdEIBPKxxSMkgEgN
3zH4k6gnCcx2muFyJexWhr+ePQjwbDrRnYeWW+dp1o4fV5469cCC9K0Gnlhmf9CMigqSqccspbHt
b5vXbS/zic9Po2MFx8JlvdyKUI7oULvX1TPcdrw0wtXtQUS7nHz9XFhlbA3Jsj/ZE8yGXgsMXXqB
dAlFRvll2JZr214s4yQibAd6O8zCL5e1oQD/CE/HZqo8XKK/8HbgNdQWZ6V3kbYqzSq+MCXrcu2O
F2GMkzeE/DKQl8pa9cQJfEY6yNR4ejey7uKUWx6nrIFYA48/QEqE5gkNsYH4c+DR0EBxp0hwagGB
kgxjLBtKH5u5noHhq8y5HWqpPtrepvrX+U6tKxUow9S0lRHReJcNP/H7o/r9Fm0LWlupJQQlcrH/
UMRUd1VFuO704KvetLPbapFeCAeq3NhE3/TCEmayFaPR6boHPUO03D4sSLJ0y5hUifC+KCSDaxOc
XHLfMvrk11QJldJdELnDVeiUCJmBQHSqGx7mhMH7KH60WTxf/1TxbqU0GlerfjsKLHkwJqJX00pu
gKji67raQS1/RxjailrgUk+e+mgShm2xzfYJ68XxvURvwIIL6AXiZhmZYyxWjaYJikslK2zM6YjY
cqnGc/W5lVbDGlMkXW+NRxK60uDpoqzkmkv4PKBjNiPgOwyaTyMh4eRBaBt8ID2NOxn81ZFqMWpG
3h7JihPKiZGV6KOS9uh515Bf1gFZ/unIyGHQIGfHqJDRnwlBy0pkhQGN0DDVeFbgXAgsyuD8LKPE
mbdop5ZC9axvKe30pghGqUhOxt4BwHV6RPMe63b4qHwkbZZJVcvxVN0H2ySbSWnjcCTrfSt78K64
AP3MMQlWVBJ1y4t41VlGO0y8FyuL0uDe8CpwfbMc4DxalQiCgPKclpEDgCjhBHjJLoWW8oaHPKPp
a2K/QVt80s+1B5cfw3Bf4GT3aB58ZSjtUQf7YZVYkD+QyqWDtYdmrr3/WhzhbilTtKfiXJ/tv19j
QDc6SEObrLbi8xdaxUPOo5gROTumM3vs5vixFQvtR73w4IQo5XNj8IiSHubM0Wj/05mSe2mWqTol
5Ilu/KgwODnBgKlWllfwt14F6a0QAjRowVYRw1QcPqem75J1KjulZ+PrGipxEl8zMtFEN3OWcood
1l//YW8iCyp/z6gFXT0VC5YocNzOxmpQfJ18ZYYYC+IZB+qlBTnFqqYuOcdtlMc2A2oiWz2Rhlh8
n+sBH0i32TLzDKlf0Tk9U/HcvvOVoFygr1dle5+NPY8F3bB7cDFk0FulRQA5bjPXkQv/C6FxtkaS
0GTyBr8krd+FYpiwq+XelPfmlkYhxNne3XdvAqTfCtnKT3xwEI20BJAhqWrmnkyJDy7IuiDRupeR
svN6uzPSdXMiqVcvNgXovtUdChZgLNxGqEvaaZQc1NWaHHi1T/tQii3bMujrAPq6foWIiAMMh7Ey
7vlRWkTxR176fYrDFMV7jg8Pljc6FBeIatYlbOJTlLLjWBXWVK5vtBJSJJX5JtZyafOdN/jRIIZV
aa/HcvvTD/p/Sb6DZ+cfMHXHId1etHgRrgw86KBWwme63/RN88swG85btzUK0Zcpwecg3pUp682Y
YMmlVRmXrGolXt2kyJ5JdjAYaOWjABPD5n9YygEjmKuP+BWKwHDGNr7qVk/vI6eA2tCgjF/b1LKO
VMeANdVgrTdTHtRZ6CBhwKP+LKU7Q4nOOgn/lyGoERPMG/osxtJx04bpgjuGSOknxm3IxpJm1dVy
sOk5dLvhapWsgBNxdAcC5S762aKTQdlt5YkTBkRvrsk5lK/eDYr/rwDFto9BlWjvc178zftX7ezC
jNM96Gr6nMtSW/UDYeRRHSurWpeEKJJ2Srj4kX/+5VVwC71OVuc9E4F87eY8BxWK4DQdGTt9UOpY
PhAlQQQqw1v8z0pLBhrWXcuMeTvGbTHSujDeZb1RiiiCwT6GXitR1dhQQrk2cZ6Dw4kxtJO0ucny
hBJw9Tno942Ui6weDrqx+m/HSpMlGjAnpT4egA6o247TGb35Om033ZXJwX16c6MCZJbEF6aTp/j3
zk/uykcfG7KqL0EktrC2cth4qkT4HGzCvhgmocaUxf9NP7yLmkd7rw/P06jGXN1w86L/R+tbUCyY
9a6jX+HsB0bMd5Jf2UjQXXRHG5SfT1MlExV44NmjAld95HAa4RpB5NzIjPHCIfq7Mj8dOSdvtNOw
GKFpc3p1qYEy1wmpqNcriUB6RbU5cFBuIpyuUnvg+pLwTB/5X+L41kU6C5x0dvFhDxxMt8wlewUY
3AdEt17ElZ3MtBLLRqzlDsTm1/Zv0Gl9e7iWPg/l3z+/VgFzYcFmB7Enc5Fthqxgo0/mW2bsj257
NkP8o6XybVBxXOQ27ETQ0CkS91Ra9mAzcqzJlUesR2AigF1Q8TR9UPWAMRSuqOjqBTpWzmk0ifys
jMSgsJEi3/jQfaTEENAfPjBlYn58j+49J3CuwpWmesQM5WzWrE/w7bOKig2F6ICzXKo3tUyFqzwQ
Esr6DxKUYpryOR1zKaYQozP0Q9rWrlJ6WBuz9Ezc6rwqCPxXdvLqtfQrDzbD8XyX7vYyiOyA2Ie0
pIFmfRRQzhwCcXDEjaN/U+dY9xwQ/r8e8eyJV0IZ+nsUZNM+drttuv7gIDB7oP781JYtyjwnDaJT
RhbKBPNGbPqm7049HPsRkQnQVpDPIVItf2s9e1Qrhf9Ncm4mgMwRTvq8ddA9vpxMXD91zvJnV3CD
OSYQEeh0oV1z3lTqiQsoggUjf1hFNgGhiVLL8uBGYfOyEIDo72Lzekj8X9ZzZK8Uk2f7bbGOBldZ
IJLkzuKEei4JwE1sl0WkTIrgCd5ipXTi7wwGgMi0h1+3HcwNOclmXZJvZGHdxKxRs2oC/QGIAL0D
pU8dWK5pAdcbNxhesCwJ1tQEnMr+W9DgXvJlft+GXEEpVVuYI0erfCC8ByLqcVpK3vn3BxkCKqVV
390s905P/ihJeAI7/xWv2b6lMpcwo1bJSLWvSZCDINHWxbE1z0sWyhfPnYKlQgio0hese0V/khkk
DuF7+KdO3ob3PJ4Q6hOuMGgNMoEOAbCNy57k4nUBWcabMnPzJ5fgwhSGvljBhynGrgDuNp7cdWTf
g0R1qA7FtNxqC0KwMM0a9RnNe7LJ2JPYRE0NpwyHoscfY45V/C/vnWaIwv5uOgHudpPDlqsc2tdY
yNUz1D9PMSfSq7DLZvaYGKNZQz8zdJXkTuWJOqGAE3SCKWja3j37TFCVhLOk3ybcVxWLkJ/9yX7E
SAYYqGJ+GcJeDJ11WjVyOh6Pgd1Y0nSV/iJOsxeUAeShJgvdGhQwK9tJYFxpXPDm9NBu21c2izS0
lxml6dFnRa+NhRx9ZQkRmzT0WP9alj0k/S4+xHYZMvAl1UqKfBhQgf7syTu6/h9+T3y0ESo/YS0O
gRh0TWeMhITHRA7xi3isqRWbDAj+bbG3NmKQy1JEMDBYMuK6Zafy+8lugwOGdeWb48eKZqNkbcDk
r+KnVjE5j0u/3vbLHVt6iyfycYoXA/SOb27G2NPnGzlGvJd1LWxNE1UPQQ1ly10BGrblvcttYgZq
mPCAsJcc2++lCvCwkCUhAey780OT1AvzSL7IwmIJEpXwcFKEkvpRoOGO1weFkN6m9Yy/hUdEk/A+
enOSBYIRA5IS5oh31XL9mUneUsOnUo7FQwCuNnKDdxVIBotF1C1tD67V7XDV92o0+gTKET3O5CCq
wgiSk10y91aF2i0l4y8ge5fmW1iCQpbrS1lBwUBtwFlqU382vAagU5IrPwUQ/xXlfCYLJ6EBrpkY
A9DmxR1zCN+BIEn+ZQi2ZyfMy1ob2i0HRQPhvS6e0RtOHJ+NfdT2uzKTgIEBwxPy20CXAUOPa7Wu
cofFtKDr+Qo1Sdm+t/KPgBz9V8HZB2yrYIPswiaqEfhV270f4irykeCK+F5jQ5G1I9rCytvGq2R3
q56rxzBqJaWYZ1l84UZ1FuQSB8lE8Yd0eVMwoUjYWHRM4lw/2jJC0O1PtHaFtwJl/BePT9toI9Si
ji1vAn0HI4vj/Rw9kMgIcsG/5fc4wI9r/tjyPgr0RUNdksfJD1gJHNkCk4YzRSIrY/dYzsHBujqy
FxHqFtJKb28iXvToWQSVpxVAI8hrkdWvM+rtYxmysJrjJEIDTvht14aOZ85JdTDWs6XGhgv9HkD9
xSWkJdvceXNwZ6UQ8t6mTVrw5+EYBo7APzUZy/bsiugodQfzTNZoKbLnv4WxyRm3hGswrrKu3pmN
dsredCtBKvkFCjL9auC9jiAE3G6dni5ysyl+EkACaria4hWA+JfXF2PXuBVdxCFcDCP/FY9zJ3sB
IiMoTu+K95zuFxOPp2oUTczyiX8OxUaUIOGCnFwPch6FFDsq1qh8gltvN4EWDe4yhQEGCut4IXt0
WrWpo4LU8Ox4c+KQsiSumDjt0C5Z+b5iwCodY7A/SxAhLOGj8d1ifm26tsWn0S2y6+syFhSxTddQ
4sOksBr5FEbNAeVcbTGZ3WH8fDWtL9eK6hShjxT/8qL2IjKxXl62oP+WMu7zwtlWaGirPf46N4iY
uLcQPeSgBxeNi8so0/sVXoMyfgKuQMuVO27kS6/oHJEQ3ynHEIslElm8LND4VJqmKcWuxjVm7uGE
YQmY/j4wdc+5ut9dl8BN6jjHcwUEIW8pbw/7hedMyOUbTbkiv6EacNLeaVMgUXzuFOwM5ujqDNJ3
coXqtZyZIfNYONF8bIEJtQfty84Wt7BWhWOrUzg0LfJRQDjjT56bM6paX3awrLgGaWn1SJouzqlY
QJ9LUhV5JJoRSr13Nj8mRJAV2hScIqLN38vZXusPlCtmNEw5sZYpJOCo8YnFRmybEXW+bxMB1Gyq
009GA/O19DXTnGurpRTtmiDel0mcGF+PSEinCZTuyMRZvFmEDl/T8TkAbMnkLOmyvpB5JAO1CPcm
js8fDBJkXYB5Z0nu1kYvOwDYVU/P0h5oo9icxBngUEXlDi2R3qnbgseahItq0hMXw4rcRX53BjFS
Ds9EYdMvqLaClyqz0h7niX9EiKzM/vO4Rzs3n+zxcQjoNDC0WNS+5DNm2CqZRYZVfTewo0DgM6lS
d9j9TIOJ3tdvTzvgh64NsHbF5UhqN0qE9WdAvytW8VYerEbwXQF0ZvjH+y53q79T5CNOsmMDkldR
F+KgNjClk98HSw6wbmHTEUOZWKwMVNHc8hpokPmNa50ueu3+V6FdKE6JIEubRu20e/I1H9DHw5pG
9XKzMifDnSWWCnMH2+frCyybbMRujbr7mCVdlaH0HJBzk1P6bChgc5b24BL4VRnfbzHdBbzFkC3Z
KOfJAxQuZlNCp7+WIrFuSOsNtG1QeqK5moOzviy1EWFSgqmw//nIt9AS1remBZJplnkWb5a4xPQK
cyEhL+BFViA6FJ+MxXgOjLMEcyXEmKgWVxAyevv3EoxyYDpWE3Qsu194xRrj5Egae5gHdk3A6JZz
TY22N/XzzWXBgpbWLszvmh0CDJebiMGEDxvv6+bUJwRdjjKJlWM2irynaIkNClbTge44U6qx8ZPS
tivR0i9nfbt8OCQSggwNiJW4Q7P79jQN/if1cD7lomixYQCFzhbjcnopl6nhQQvLtPrSgIt0NSWp
TBjVAHSFqLEfuaLe+8vXI2vqDoDyVfsQQiKY1oCXLHU0Fv/u/R6MiY/omhzH+uVEC8gR6x8NxQPK
Z64gyFyz+Yn0Y32nSdASro/dXg4xI9W9jGJxjtBuMTT7xu2/amGAaOTYfrB/HWNHCOaf3IiSqNaz
wtgSyCaUd3PViqQWfmUPuO89CdFGdmqWeorzQIh/6JK6hPMCz/OOGK+KMNXRrBFgG1mi19fyPMi8
kG6EnsHMmfOh/nECU/BMpF6O/dosuwjXoGJz5B1EjYQ5vB7Uba8ayVntISUiRTfRddGWZnnYxx0b
5HpeLiyAP5nrkIWYMPkt0kJYAjBE2iKWRRWzVQaFYJ8w5kvY93+IWCiBeapq6EgwkPy4Y7FyF4IS
OXYLjJizQxy2rFwwV/+QEvAjyQIG07iA8MZrwORY3p7kBllKKDjeQyZLIZvrV3IuL4avb8JvwnhP
gaglQ541SfQmbECdpMTSSuxgFW1EFYXk4zH37V97WBLZJ4Ki8ROG0sdkvWOt9ZkIMLglLhT/2Q9/
ulXywUBZHnF4QVbxF6fnpQz9efhz7FSoWTVzpUWiF+qrOyfFMIwT8lqxCFizIIX+u3WpdX5iF6oi
C+R1S3u87qb5djijaPM/75CcGQbJ4xMDtx3gWryB40omMEciftL8Jcktj4Nu/Hd53bh4a6dkL1aX
FpYRs4UYtKgF0/6WaRomYnwXnoLPfhvExSdOVbA8Nq/a+nWm0zosb7FuOlrvyrxoC61g0um+VpBP
QfpgKiFUTo28RoBJ18vg+xIRabr34tI3+GGejUatQWnQK9ChdLkuI9MQuTXIsW2CuJ7JJGTS3UnK
SQr6xVMwfVn/B6fUnDiF0PKjysUttGe4AGaN4jf8AjoyBwpxqYsmeZ2PYojKnw29Z35TL58tyqu9
xukES8dwVlvSu4XxfMHVZNs82+4viQDSnY2zG5ueDLQdT/Bgz4JASts/20fW7kvgsGH/rv+WnwHY
veyFeW8PMAD2bD81U/08eet8hYSIhBQgIHvxHkkfkanpcoSmTnnXwk2Vh7m4E9xYDmOp5LWRhOXp
8x4Vq7W3DZNWviGnACFM+YOGZimwYa7am4Tt8WhfmQW9z6fSvgLeV+GJGakVO/HBpZVq7gSKEWPO
+dPRCzD99oYdYM9YUkUTU8gpz90tsQYnJUhIdJ3yNjplwF2QkrTlB3R1KNumeg0cpq9VA5wV+Zex
zbIGS0MOaL1tIyUyhGrIYpCNEOh9z3ehN280cyKtsSRXhlh8Rcv7UHUzykyfXosj6yUi9tM/A886
7hns727b1F6pcF8bk/evCot7HyJSPkiALCOO8uSUnpKb+2PusuSx26xo3nN717hCKZ/KcrZcMMRB
0vTZvU03qKEUgrNOH2qN9ROB0ocj+erf1O8Kl23C6XvRmSjxGye7kN/06iCkJCKWHhfVK14Qy3IT
Gcm31p5Mpc9+S37l8BJJ8wslmh/IHn/m9kCxlgqbD95RQJ8uAsbzaKerrKQKrqP+tA/HxFLcwxax
k6d4hOawTYD6WkOmbNiC/u1Lv5kAglC7zBXY6qwYiG2hNfyW0GrfXFkP/uurPfhSCzQ+ic1Xeivq
BoNPxDN+yy4ZbgsDlrdxfDRhNAiwI6s+KDxfTM8SOteGei/C8EBkNVYKb0VpsDspsKXRv3aFCGo/
pAKFMvQlC9YytOrK61B6oIV77e3tHeUeWqG4/vxOnZ93BNb+0vLozUGnIINyUYU1xTtViVrZQ7rQ
rh++lVBErPqmAk5/N8Qht05kqRdI8sdAxrhyFtCbAzpNhQ7KP9NKR66fpJhi2MK86rcqBA7FfEfP
rkyy37JhuvfZ9YcYtJOoaV74Ty14Wx9HX1RBDT8CfKugQ8bO6fg5Z4XFuWXwFVfQybDGavQ4dfSl
Km1e0C6kianv5rNkiglCbo0n/i+eDQAdk0u/U2N/qwXqA28JSMMUUtJ2UARw7rxN5bf6tbTQt706
m8VOJlXU6gyALWpEAHJebSe2Kl9py6UgtFa2nifHcuv8c6ZVrn+OT0Q1bsGxIvBv0e9asNBrB3wk
bRBwLngfaS7VTxChlsiVdDC+l7LzO31Hsqz+z8I4drKf5ToS8F5cmOY2l5uYKbQaGC5HCpLiZJm3
U3uYg9QNt36aIPreCmqzad+Jiavln5mWD8t0YYT5L/zfs1HjamqAcF/t/F3DLqiAvkG/Xk/aDQh1
eMaDdxBi3BmnI8FdwfMMXUWy0UV9cnIO6nXzhiylkdXxZOWPBv5gtDAxX0qo7uU0/0xq2xvglj1+
2U3gzDZEv9El7eoQoRdmamhVPfFDLJekZ5DaRSDVoRkYmA/E8Hn3KIY4dh7bygPk384YBJK8oITX
et+LXsyCEN4XiDUfkuHDgV/e9CwCj8pFcDXpY3y8u5uakJ1t6QIhaAp4gg3Mrap4nDbZN1Ru27lZ
r1eSOkJAfCKauZC/RQ/2bCoxSwAt7LgAc+lvoqV8bO5M2fXEoF8xiKaqrsIfyVSaApdftGe9u0vU
TvTePIL7/IQvxYPDby9PfraG1aCFRJeGzygEUI93CJ5kVrTAF18dOIuL8P7whiAHRTXYvtQJXL+J
J6Pi/sXwMPTrUBAclBVp++bKi7S+4zx4BtLVzFMSaCmlf6G8XXAAwQVRF7clzADjg4qlbonKubx0
BkraC9JwppGCG1kE3+n8fKYuJFGRukc/pWl9Y9d6VGJSprziB+kMODOBzpJkoT0TA2P1OTIgIV6z
HZbmYFVaUaZ8HuNQbpVIyZSpDYxket+ihr90GfVmRESRXdaFXQOnpcnTYrUB03NX6X4gYxkFtgq6
Ois7k4OBbZErLPiGQC7PVgwsc6nzwJYldnAT7ipEHTdzfjQ7zKQifzKfUc5XcS5q5GbBXF84QDPo
jLDuBgSzCeTeMzF4jDdY/g+8BbD4WEqxfvJeKx1jkqE4mM4fqWr6UiVaR8nHO+pVPtkrraLtaAJq
IeR/UcH7CYBZu3bHS4b14eKSTnekCVQ9Y+JkFHmUkw3lf5Ml9h7bkxzoNmrmjlwbH1dXNdcBBn8F
c86Jst54mF4zPpTZ4o5XYRthvzu9LGodjFLiO41Uj4tLyKAeMhnKp5DQ4XCz9IDQnfBo8XXKehO2
UkHJ7GQW0u+TVQv+K+N+btYFBPDqQDmjtiCqUjcVTPqTL9ks4TUkwdQmZjGbcap2K7NOKG+BIWKn
OyvQn0ArPbMRSWAra0yfHn0gkejB1P2IXpiMt3Pig22aT9oDcb0U4OQDlJR8Fb4xDnnnHjp6dmN+
VtcLE5cJ0T4EBh3KoBnRG8duAU10VN5HMW2HIfk0FrjobL+MWjTLCrxAQaNee/XIO45AIcsmloub
S46pR7zc8UdLXIpNjdjl2rxCFSI/6CQ6OzryD/XQNJGRSsUd+qj+LnH2Di+yrWfji52Y4SU+gOw6
2og4rZWN9uAoYGVyFa7sh50SvhLdjztsuORvALMc28fkkIa4+vBk5j0EBNL8a6OnGrdweKZdo2W7
YbqW8g94kTuQqy8MO0wScUjZ22BWClP4RDm4APxTspS9SlomsMF5BRCOUfBId08LDziQorrupuOV
ImoPdcvOuT8HZsE9jIRm8HSizhdp6Nq2LaVI8sxA3AARq8Uwz9FYAd7tC+IvpCllA7Jfg6IxJ8Eo
l1mcwyM7Yf7sUC6o0/mF9LiFID0DHvdcJLqvzenKikj9wqCJvrAONUqfb/BEJn+/CqZMj63INSJZ
UewoVb7o3PjwVnW5qb4hlHQVSr8hax6g6kuE+sstji/t3RwvMuX/OXRCckdpMpSDXEUfEQNdDm5P
7TzL8DEef4IB/0iOsTazUf1tERRrtNnXUAxOvFNhkam/Zvh1feEcRvCNb4MbhU1944/EVMCVwyYy
B8JfS3tBoWykGoqK2SyN0Yjtt9bbykc9r/O+B1sKl4rmoe0ktdmx73KizN5tm3Px8A5RjigegNJE
db09NbgRzIc1FAso1MY9RbQPE00/7j4N95jD7mHKKbi4brtNiq+h7/Cv2kSVRHGPFUqTCOjnUEYc
ciYvWMaGliFxnhlvESsnU0k8m6TawDUEowY5Raf258MAmKYWpfS4740XAEwzp6g28R/NbWoYiRVq
Hhyv624hdq5l2pARv1L4KKusyimd2krhnjGluYB6X86yGndH1GgWFfD5M7cqw6ej9pEWSOW5uHMa
gFyj2BX6ljoIIStynBnzN6wCNb9fDqBoxPhwHSZZTea4X59U/4nGbDE+3XbKB4NiQytmti4OZpyO
SUNMm7wOBWEWPJVArhB6J7WUM6MCxTHzHcVZCsDfUDFSsAvtm2KXBClJdPHR7M3PnsfJKacc05NZ
+FIr/g1ufWTBnTQDKbeWIOcAQIw+dB38cgnBdyw0DSgU+wklSlwKG2b5xhMI+M1HSjWXa798OMQM
fYasW2+dNb9ee4pvsY+afCxqODMgH691eMzd1dKiIXV6wW0eXKAmJBKo/AnzJcgWh4xZIqT24EAa
aIcMoxlvXPgQM0kV6BMjx5lBpc0vGxMtL72sdr7fzpUGfk8dSmjUM8OT/uaSi+kZKSN9FZ8ABgqk
SdkkZmkdHSVnvAbsveaXaV/sFUpvHHu0bIMNyKpoDvjd53Tq+PXYzwE84jqv//hTC70E89+RKhZd
3qMhH8loY6p6svuUpocFhDbfEw6cHBP4CyB3PW4SJYeEXKmZcNwxx5WjEx+JRs+kwupwNA39WzR1
moOqNOZQQktxKYx3B/XH7qIZezjVkK5EFKVp5o946NOq4hG5+3TIGc4lH4Ao2rTNR0jUsn/Ei5tE
O4WVZBVmyXrurIA+Xp20y2nSJL6xt8A3z3gEXnq30xt/RZHSlhFfUi7iTkRe63mOZi1YJ3+UW7Z3
h6TsjR5UyKajJzgBn+HWE/BRYKMS1V6TyzlGDdex064kDGV1eurwK5FAEJu7MK1josBZpMW1AI24
FySyoG9HD6z1vZx2qmBI/StwhHqIBvS86qmvGiD1Xz5KmbxQhnCcZOxPEXRKJ8gwOyjjXeyntNgE
RYwwME279QZvq4Q8iQGrZxQ9XP8cmBHLaISNJgGjAqgcrvujHi1nE31AJurXEx7FIW2dbN3V3zJU
UL3FcUl/vZihKKOTbRSRvPZbtPSAqqHmZW0iGiXzAJpvti6HTb6IkzgZrKlak0hNVE8fA6BdDNzo
u0oo4dpl6J1TejTgkiNQzmt/jvdOaUxLD9iexuFU6/8ryL4e7uJevP/4APyYAC233aclFORsuVNl
9uVlrqNQjwgNi1y4GASE7e5YCaXw1ANgTTjC1ZSQ8lI3h/9WppjOytQbZJNEzPImjnSHTePayiWE
M8IeiuIO3+dLDABlGtnPYjCDV/EnVOBIwGPcvsxcxCdGSzXIs7k+r9O+X6TPQWcWHCXghlkDOouK
gNCoKocEn9c8rLoSapdrWzA8NiVxz2zVklQLWqMwConbkpHub7FPX4yM+KfS6aPsQfTs/S+6PVPm
CJ1g+UFTY1eM+w3N+YbTGKL4JncvkJm7SAe1KoH+ptZfGMB6gdt+OBpunnnUpgNHBiqfLXp5HpZA
wZQ3VRC8v7xvShvpR/Ym1eqQgwTCf7ilFqY5vzt5qD6DA9MNgk7BRJUWtuRW2ksDXfnWGCM/jAsF
kL5/gYysewiyD5FPOaTl1tomjlPQuW9IhKqpY5zAEd7Y5mBXxF4bwSQsaHIsgbZzpeC6CE56z0O1
mRZVS4SPgX2masGZ3o+Nex3D98h3oEqrzKIrtMGUb/1jsDjP3yyoZzxKObziSZFNSAUhLV5b/mk/
903eAU1Nla8kn4Php/+eLkWMq+6EJLUrO0o8ZolgEYabGoEpwU2BMOBn3MLLqu3M9Ae0qW4oVxRJ
XK869jhNvVa6nv3MMG4v0cobfkLa+MUNHrpBed1qhfoHQ0xbK6L8pPhsL4i7xAJgzMtDbwyDho1g
48by/I2wBwLIlWFFBi/2+NPSDruTjUWIv5ev/1Uz+lMlRmI6qUQeW4iezge0ywb0L2BBGPFSlsLH
rF7zgPX4jOA6lcOX4zWI8s8nFYcWrReDJnw1Qp5MGxXI0jT7a9oS8+TO9CL+hemsBciEP68Jb+ts
2zO/6T9CnuRJB51IGc77PocrqtD8Nk3bXsK0ZFUbPsxMZmdtDBU+xfiCbqpWHglgLgFB+l7acnNw
amxvcfb1Y3tca7TsfxiOHuE/lbNpediXSIHHhL0tLjdIR7CFJRFtXzVcWy7Ncaw9QvIu3/uByKpy
8chXynEQRrhHhRGlhARPC5GtEVeln/dW7yjN0pELatOIMlVKXCHwfUyX4A0UnDJne/WhDN22/pSR
94JL/XUF2oVNZdKWNIj11k93zH/rcJAr98HDT9MzqalWa1HiChsxEwoaSS4QRXVUXodcgRwyLaDc
gJz4xyVVVPX5amnAYktpYW7A2ZuCsp7+sE2znSX8pS9M5FTTXp+CIHyw7oUWQAMZR7dusdlQHU2c
EjbBXBcecvgjZoY7pZvh4PK8AtQ0h1xWUkBmsNbJrYt3NX6znCapkiPbPKLXs3RxkWOys6/AkzbM
zNEUQc0LPCBqJFzqPnSqaeWdL7cFq92JlUOAaMnQqOlmoONWiMZFeYZAhCaNRFm3OffBbLGW5kAw
wqndLc/epAIWEPxF37FiiQXnqaCzzNGc7Nt0mgtbHEF+3ucSdMDnZ/vZw93o+T95G6XD4daoOl+Y
thhDSTC3UW8/mid/UIbs/EwttV/9oGF1CpZX2bmJP2fQhpsG467VWG1WjPzT17EIPDeazNDT04sq
vIA7ns8A5j4yZZImsQFlYdsML3QbDeBKVHMnItpnrixA2fln25DK9SiVRoUTavsDQBfP420Yb5AY
vQjq+e/7xjnKxrH3ifR/dwt6Uc0w7Ay4F3DyEFLfPgIJtUS8qyI3GPbUnYMoXt4+6WFadFbGfmCi
+Gd5rrSpFghMwcmOWGDIiJi2ELRRgXOTsvfAsuHLLlyipFceR+yBHKfAMsZXZLYVPskIm+jKcT5t
sG28AjH0KdPU6HuZuWg4H2sSs0eQz16qz12WY94p/oKHQ44OyjBqbSUFPS0mKRwfbcFYHyoR0me7
RzsTp1U+BK/owJqkiSPKb6XQ/VzR7hb3i1ODMx383mv7dSqsLuU2Lh0DdVC8vH9bDx4PhQ2Sw6+/
aWAvKsvw1ZeDBcfNo+AUCCBM4ntkkgk59eSfCSHWMH1YM4Cyjg9Qmn/6sSLS+Piob0Bg/rF0TD8F
aujK0naHd7+mZh3SA08XzE7KRRwQRJvUpMsV2t6fxGS0eWJbejx6KZ20lHe1I8pj4lW/x/DAcVCp
FlDwfNH6yVQmeYTvVfIy7/Qd6X3nRLDXE12FisgBFK7nec7E1xBbaEsk3kDrh9iJRGgRc1/lSAkt
e+krUKvhhLLRviW/rO0o/oT29p67Apt60SHIJskS85Dv9MKxO5OZQVb3gXT0OjHalpef76gJ9pyc
9vtizhQOQSYzCD5uo0ZcnWKTTdU1Lk5VCOFgVhPQkHdvyuD1T1C0gRGaSQx4CfO8WxwGuifO61K4
KeaeKH5sLZ2wiY3lnjRjfPGbsySZ9vfV7ENSE8svSFR0sfHQc1PwZngK6VbwRP7rQLjIM5VFvO/j
1cpgLrraMp8p5CU45IgBc9yhWSIcE0+kT5z7t7sQEsNpbkMCdOH7BA2dhRw4HZwUiG9C9CjPpYIf
vvvWuKd8omjnXxkj1xKI0lWG8yf4pj1SQcWkU6fKvVYLUMCKlmRpTxXEUYBHTxbN2HDkx4fHMJdd
Jfk8Tdh+WXw+JaXmXBpcTqwlK3Ssvds6vvFgxpxShiQVKbiKJgzBrn/piiKWsFR5lQD+UhUIzwpC
1/IvuWT3JpY5jDFYxauRErUAwE5VZLvsjUlyO1PWmxroKpvHWUFH0BhmMiUaAZ6AyLIJxTDAQI+X
+3DA8DgP0H/nTQjmrudNbXkfkNOIGX8e2DX0qcH0tcs+PtJsmUFcXuiwgpC3ChmIS9lhcANWjTlw
2zUFNo5Jw5ramdztAXbfMBpExcLu3jT+0JwIFyHSXOij7/6pKVT+3+LINTNW74vt6dtnpPoSYa9D
FtfkIVoa27urZ9Mt9qmx/xdOrQKLpAfPejQZf6dKgufYE31CUhNZkEbqA7HuOuoQ9aNKjZsCT5Mc
C9FB0t/cej2u6fz9Ob+TQU9eb9YCfN/b9wZRFH0PndG/9XKhWuHn+mvjFDqrwVpLUSWhW/vfb2ww
bBJZ508mlyrRPPIfp2hA7YgI9Y70bve5K6WZi0AO5YUwFK33+QNSmmbJNq3xofuUq2m75KC47Pdt
n+Q/bs+r8ShRMi8JTgNfaAk4hnnAdFLsiL6rxCaSWOvrUia2fi5SdONnNLQMiIVYl+3Rj1kAqLUq
m4/1cXitiLritqoeZYKhKnobU7t2emKNlk2kkawkAXpT+2Ey/FK0CtqYeVMq8UfwRBFIN0J1EPAG
6mPLgkdFgCu9wF30QHVC9KmEhCeALhEH00AUitqPjzGW4slAiPqIijpaWIIoKMP5qm5I0nL7Iq/7
8MlA9NgPOSNNfd3R5lO+F6eg6FKp4OoPtgQuu22gX0G65k3OeSOOjDbTpsc1D1/jB8YS7GkzDD6Y
CqzmA5mmD9YwWAvR7LTFAPzri7ST/Hl4VQOxmBvX7Bbg6SxR/l2GFVN9YcSnvqidMXvA7KK6AD7s
saXWH8aZd9k4yayly/36t4X1249TmvFE9PWhcaPIt53YoblGVMa0DZi1230O9VVFTVa/2RsEC7ji
pYKjJcQCgZZNnuRdQPfj9x1XdNo8KdS9IzMxhCzmJmiCW24SYtZLZC0ZAoztzDk07duHBOshvK1q
7RFOagk0/pS9VidbHz45hFePeCHoXwCzmbmKUOuthNIXU9QDJsfGEdDuvxhPF+bQ8RIWEdyi757A
NKbAnJtUMpN9WDwRzoMM1A7nOAQiifWy6LKwhwmuSEQp7G06U2gQTKp47d0pKCTiACNTY4FRX6H+
utYLxkL8hqnhQ8yjSPqikJhBq49gWtT2iO8YSIm0ILWosjsFwHZ3CtfhROVtdb4zN9IxMSmVTgDf
e1weswthn3T5LWa3NQSyVIlLbZMOj1ezJ5A6lQXc/qKH5XVr2epIJMPvJ8mFRI9YmPQ3HTar3qJc
y58U7JivtY562A5oZY2v3hXgmsGqR1IkbSMN9rTME7DcGml/y6XH/Os6bWynY2YoFwUp+Tcm6sDa
NPk+N3KV32CAc6MfaRe/wWEJ9Qmrbgh6OmBPndDvMTN0huUf33TT1P0epc+TiuqhR4AXHqwKQdt0
61OjQz/PqU7sdDyw1KNtipOiJwGtBytESvWc5RtOyUi0EauaQmFFOu/QhQCLparma3wdihiS8BPf
CSkLKXOQeTAW1+Ltho88SQBTH+xVNk59VlTWtfaG2jtETc5q6ui/I9AlTwm+KHRVh+vPrmdj8J5l
/Ys3g3D8zqKASUSfRYxVUK6suXocdh7SHRHggiWFjwmBw69V1/6I8Uf+IvsIfZY2cVos85433J68
46FFxFRccEz06ER3XzfLCs+1oJRVMP5WQm/AfMJ48XeDmb5CelztuzevRyr1uGrY21gANeVZPtBj
tURxCMC5lxI5tBkhygHvvXplS2L6wV/IiMHiKt/RqkppnK8Ake6DzB6GhF503ml7IZkwrdV2J0tJ
jzAPtA+6rcYPOZoJiYq1fC1ZRsJrQ9KTnL/cXgf6mWhjsJkzdUEHlijtddiyu9wcd82xX2yBbTyt
ElzBFb7daBSEJrKhekvzUiS7WJFtxUxf5HAm31+B/lhFmgJDYLhJZBDwiCCVPlURPhJB//3x9vTy
KO+qWJ+hanC5SNzcRQSLpPGYVuqv8+K+KAN7PB3wmLpPSQ8/g2OBB87bnfieMpW1ci1Dbg7KZmGB
HR/6cfSixudBWhiHhlj7D+jsKF1PTwL/rPTf8yFDhjQgScsfeyLYPiLKH+JpDxAmvWGvcgq2htxK
QKCt6vkJ4ojVlUBGqUHwtATja7YOT464o6G2ohayTloo3oiYoqnZ/qn8yStw5tox01oU+oJOylRN
6H5lex8tUvPThDC/keIMD6yuRMdXL+zqtzYC0Kq7TCqyN/NTooaMJCo7xCocVlz7fdSVRc2jsyJy
FGiHibAlWPa/8rD5fmrulv4fG5VovfljNoIcQ+KxE5EXMiG9G8ibkR2aG8X86PYooJQl25exvXAa
cRYagCZNdIP+cMx6Fe03r5jNDh+fy3dNFYX8m7n5378WTWyG/tkthVblvEg/ykG92uHqBAxbfS9l
EnaH6izmK1cpT4spStgq7MFWv0zqkKMMaudpwwtUjZwXP8iLQCAxBCpQ7a7Wk584IP6MsrvD/QjO
20utWgmsW+HwAIVdVDXcZfcqCRBvaWZVvoIq7+r0Yu+U4bE1vaW70CJK/zh61wyrOKq0izdHj2tH
xI/Xcck7wShlu/rpfKlpNqsRzgfmKHGeO/E+wqMZet/e4tkiOArww/8oTi37a51gIBk8DwMRkcx4
1aGpg7R6IBYGmOeWco/2Avo9vgxjZGqB8JMPPJrpQ6k8pCMXEvsf0gRdJZDZWlIgeB0+Fw3ZBCvC
GkZopBLSMBir0JJR9ehrHnXd6ZfXh/dRvexAJnPxJSJo1QE1hmcIcUbnqaG5rQ85TZOGOpbKK8/m
tqLDfvdTWFXJ996Uww+Tr/g1phtqEugJmDg86kRjCgTd1yK9Hf8RKHTedmeG1DmKhu8K6GCalnG9
oWCDlVjM2+zTCtG42eipwbkmAUbXiaNQng3mf83Ay8dq6xlugpxAbYb2XVk7YsjmdHoxChnCHIiv
qcEtNczWeKt9eoDwZMuKXpG1uKJjooO9JFlMRJvdfukwRGsTFQXWnLC89QLeE23efFc56VrZTEOu
71hZZjmk+Q4g6VG5ouwqQolvI6fWsMKUiObRJJ1HcjTzqqveEzXWZtWlXOdaac5iA8tEIhD3pJ+l
3l9SpGXS3HZSkJxbLA53jXtGz4KJR2uZz1eIeIqYQIwwZHN1/wDwXPITCfLqK1TxDdEH+OlEhLgs
i1eK0QvoRvnYlkKvdeHTpgUZgDMVYLov21cn0leGL1fvSvGIKsHPhHtWdNKeJALVrx0wvrT4+T5m
5HPUq0EHu0uemOP7zRYgh7axg4eNG9+d0zeSURM4JZVXja7hWu52HbSrvb4xovuRsqssjwnuQE+D
A75/0x+cZ/J04YEbXGA871aBJ3hfibPGQAEt8mQwDEGHCwZk3LapfO8aXrAzBVp8DAZu8r1a1FDi
4KxzBK4m7o35teLeOMkTPZB+nuMZHQgPMvZCsY552rJ15WH3AiTiKaII2FRtzRyq4LXLi41gHfsy
ipmkUcQ1TampfLBXu6/cifcpuBimewcfLKD+t8NNJQEr+naNf7WXjgIF0KqEul85EZnizmLU+XHN
vuI7SJFgxIElWwaaHMKgsVHAzZndhF1qRhOnnFgjz6EupTTPel5hyu3G19cx8HO2mh80dINz+x2t
mUIKcG9cFVptPu8iM9S/pztETnH9YY58aiAjlta5MkkAqlFofMHDHhjKJAH4QpNcQTxLoyiAcQbP
Yu3ngx+CJh1UtXNhlu0q60R5RyXbE8y77AYmqv6U1Kkal2vf6PaEuh4DCJd3AM5gsczKSIsWooOY
B7EdiQV/Zc2fk6tGFaUoUskfB0icQHYLTNpqH3Qmr6z94V33QnDxmKzgO85Hp31jm3XcssJ3Uvs1
GjRVYIbZKm31RQINlps8way20ygdkgeVPRBbFDlgQ2YGNLE0/rMPmlAiD/68ARkzsTwx/l1RZTPP
Ecknt0ukBmvjLvi91UJcNGy/0mpgKrJDqtufj4tP+ESrymB96s/6fRUDoDKelp0ERmgQ/bcameYN
81IT0155AHru8h7+JcaZY76pARoOIyR/EdqH76MBfQTF1bFsSlZ7D41gCEcJhW5An5f49eRDuggN
TtTvTWLzRC/smb0iRDEmnp84eQ9wp4ODrOnimaNk4zEBgqfe9/OoFcMBg4Jgk+ZpocBbNmRVTG5o
ZNyIVjfazYp1gG8mBdP4KpwpOmxk27VJN//EKjyeIYIVZBu55Vbs9KSWQdZiPfEnfrJR7v2groKW
JC2VjCeIqhk80jtJp6SUIfbptHE40XF2OJ77SJ1uwSPeEeRYJoY6BlIHHvRC+YfQlRsaJD9wCQUo
pLM6ihSvhs8LwnXBtuizdy2NUuerq/3lmwA72OVawoIEk2ilyDHBYuclSr48zg0Mgy8P0Hh4fa2/
5DLWz9rCCZ+vfpmxOC2d4/+1vpNokg4GHZUSnqIQ5ueO5cCTZ3SQu8ilwusFGyZzfRDwTr4pYyO0
4PM+3Jup+h2b6o6+n8Oo0BuB7SfCECr6zmWtweApCb6b40TYUctxMdC2ZY3DAVjLddwIDlELmg6z
hUJlKoIyiQATJb1o2j5jSTGSji+mETU6tV0BaPddW1tpU5JwN0donhO9At/UqOkyXWKCC4QYyn7B
nIacIkjDhz6aVslAmUPAAOinpkEgl26i53XodtBSF8kz85/EPex7eOc3oWqo6NK/BmLS8YWh9SuL
VyjAKwsbWR00aWrxXDJIGnxxSqQ5kKn8/flCq+y0jc1I56apCY/iBr7ThoyJqUp9or5KATshanmM
jDy62pBLp+mJ2lXPVjs+rVTm779zTR12Z4iYRyvfIlh9b0DnQRi/mrUjLeyqH3pJzdohcjP6O2kn
6ah0LquHBMQa5gmX8csn5nT/dynaE/X2gi+xQPGiHMp1xD5erxRunAk5FXxXMH9uw2Wp5KQBSYe9
GLj9YN483hIc2DkeMdYUPnTJglWqc7kZ3wevG+XXdpJitIG/qdzXTAW48/5W8TxwWW3bBz17xww7
OHC8JL2zhbQjsSOc1gwDun3pRxAN+tvqORQ7DT/NmmT5IPydr3430jiVPqJ52ZVJGqFvuHNXJ2Et
R27bN/4wVZwL/h1uPYTFsd/iUsPn++DvWhRstfazuTJcV4IX515mR7rrkCixTjOuZYle9k0jiEsi
MaIOzbwX3f3WAzwcTksTdxHMHLUO1jWm3nnQ3LqPT1nO4qfIgKBZ+aoq8HIDsMuVaO3whdqVYC0/
D4gv8Eku5FWKGHUYrCUChn1hLCRkV0u4+kfnE46Yin+bEPQgg3fsNkjloLx2MowehBvONs8UqcCE
OK2m7e91DyyxmZ8vSNBYLkyzZOEXXKaJnG/PnGQmxxl7O8QnoaUmlOaFdXCqBGY3OOMv7HwK30oz
03EEZ/JHBg7ZX2h+RXqZ3xx9LCgeeJZLsAqwh1Gv0TiidiHgC/3kZS3sRm1SLdrod3R/tedV8A3b
pEcS0OEOWTaY5bISGIl0UbkoYz229Oaedy7QmVpOhpzt5pFyiVDV82N1z9killtp634z/j6Ltl/v
cqxIZ1mOxgCxTpN+/QDoEfU+uj9SDonsbYt38IbTqrHD9EEzyg0A4z8Yhsi1IaR+WJDz+6SEGI6O
nx4FieHc9IKIPWNSqwBhu+HFL+BdOUSNHyRgeIo2RGf2yccNe6IfL2FLnkEZ3uIhcrf8UuPfOQbk
ZOg82yzycuLFyJUg3/Vc3VqXQnPqYonKNyNt5t7DiMP4zvd74vlVMsNMm4UdgiuVBpcT/X/JGVXH
1pqbH8tOzHtJqY7JcisYxmBlvtMs1WSNZuF3VArOfu1k9gmUWh4XYKJgLjctX/yzHvihwaJ7QAaT
ayMqLJoR95IbGNwNMnpFwTK2C6GC/zGLAFTcxEk2Inn3LEI6hD7hvo5CtA2ZQJrIjoLKsfMtXaO+
IgGQEt9lsyS/8oiPFDrbLbuwCVlvgAM/5I0NKJZwjetj7jjP+x+bWj3MWqC0EQoQl+34BSwa894v
7x48wXiPwo6sJMqnK+SoyEPxDtSjZsECFpceaC7uoApVvSLesL74NucW9OaHCPAzKNxOAexunbmA
wFBJMBtc2ffnqfBkT6KQfkX5kz1hOo3qdRQOxggWc33mhVcQLZSCTvqdE30p7wGQdfMVoYbRU7+Q
uMK3Hyw6GIxhGoptXaQcQWq+3oAqqmbrLFRaNvMfaPEe8mH0MfXXXxeP/3+vbq6mFxNOvnpgTnlA
G8iFcf9gO/ndhdTP60VnqhUCvSArW3RcP20M5NTDKsSTmU8CsUPI2i88yHOf71Tj3r9TvXTe5mel
MSWie2ao/panTaTP+DmH1nLkVrV1o6LUZuEOlz4Huxgv+VwNzeQhfxuH2Csgn4gUpRuIIqcgjRqO
afNogSgtsnzwXmX8dXriM0NVH002Kp7WLKGvs/J4UZ8HTxrxbpvxC5muKkG4aGgHDlbd/MqNKNDv
qOmgghYHtB7zvHa2v/wtTBwc9NW4sWkuZvn4e+AVzHnSUe/UnDpuqWRSBpcWLkFCOcC62eTiRXGi
ln8XGrXzgYtT9qBlheL0Yyk7L9A2CYkYmjFafGEwurt4TYUFTz5EK1d5Aed0WmAQTIIYcIw70sW3
br9YpsGCh0B5U+ZkfOUP+Bz5GaG43gGy80F3TI+oxCLNCAYyo6PQl54rKUxjdCb8bS1DLEEdpTaw
/8l1LLfQPCd9ubTK5zMu/GQUw37mJzt/B12JWOjjFl/vOsnznWHNWMozZvjY4hjB55SjMR1Wq3zb
ZPBGUUWq60jJ1Dod2sgeAqkjhMlXu4CsogswmEucw1A8nLOwQlNidkEVmqteLRpBbSwmGPjil5fF
uhD2DVGvo+onfKLNwuLcy/7u8JGk2YYJJSrxdZHIH9uBYStp7s0LLu/F/Jgg+MLCEfQ+TIPnkdkm
btAzEM6eZsf9cowTzA7nnfk6c0cD0Mmg4Qk8wVydwTgMDxxSbSkYT0MdqJhDBGf8NGNhLYlUtCpM
GHXWbHXxd7+w3Fj6MUlvbq24rx0v7ZEtnHyVCi53WvLxOAeTRRwzqh1anqHkivg3MCySq2ZqcbF6
vgLVKKFWeTVIQtFFrteBKKI3PlI1Z1gWk2fXPcXMtlpn1p567saFGuh5cla7qXCwG5N+sU759mgn
+8R8eJJqDFt6APqoJ9oLu0Kew8HvaVAtaAlaVbQnXxnq6oWx3DW1ys5jsmhUFwP2b1l1ddJwc1B4
8fVTGFWR+vd6F072Gq3EaGUFndpojMRHuNHXEI11cAwLHW6/Jklo9XBdO0nfPie5ExKWuyCZsYpG
ChoWplfmKfP/OzhrdD5crrDbttYReYpTPXZO5udUSfoBXsa3oT2y5Lkb2cZ7sSsw91AbtdKxUTdP
PmErekoFdjim3pRLzgZPsCbcUjnXxNGiX10FtEcf57Boz0LNjaVMps8J13tDqccRmPh2qlhD+cUK
/osY2Xh4uO5Mux/hL3XnRjTE+n/f1U59aoo/KRe0YZ3wwTPK41QT2mc9bwf8zdCXKZW7jXegJJcW
6eRiQiabgiBFOyW8peUtbHv5RcY1lLF9Hpv91gdMx7T4Lsvrm7kd+AXnfzk8MtviXgk9weOZvtks
qPqW5UpUUxbcip/x0ozTREwVfAO7h/sj3zC3HV+hX3s3/rBjmeIKd+KBbaXSFSd+fL/a7XsZ9Wq6
uMoYT3XImtpCu7YtpkT1nm+qsz9qdKKwaTdcfUVsMA2+ARk6pE3OF0RPGgR8CpAnhxZNgS+YYGQe
8atAw6QSaJsaCD8qkK3p/Jt8Si1/RyfHqnymYzdp8eVDnn0ZJaE/oZCfkTXxrClJrtg+pA8uLtEI
fRjIu/x5N+ov3wUwHicX2PlAbcxrtm3I54Nc08AVcAXzpaKCAk/LRquPoVp0l9u8qNHwvAGYPjKe
vURWL3N+dQStueg4731PVt47V5sseqGdel+aQHR55cVfEWTufLK+c9i19nQRgWAKAM97jH+4Y337
YVqegc7bqYwy2qYYt+cyG46xN1a/F4Cd2LxaNZo4PVstfW4/mMa4VoicsIhp9XP3URww/tT03s50
putQvzHgJKwC2v7lQSILiVruEj12H43KmzKonAskeGri/lqDKI+sWGfY5qX+0lwIEkE3U2AlCx7R
dMj5B+XaEFkMMfpFYGMXbT3xthDDaJh5Fphg67IdMWuDWzzeFYgV6FPeag1hWuDvZSR1pTquajFn
YJqzJneOxax6djPzd++7tkEKJknIfqrxZ61T726g4C31zWUonTDdM6d19ty22pa7esOm/2f1DGbu
oS7rFl5xNKC7dGkckaVdZkiYlajYWWeAHvcDhTc0ehmikkzEvQdHewJHgamhHe35/uBE1zgGFSXE
VcxBXpE6n3+IGeWyxeGfDIJJglPKhJTN04yWhzPwWsgBUcV5GZ9hpWWSzSr6hECe8EXMY/uAoY9o
ZV+O+VMNu6XLO4QN5GjvlEbFt4f0RgmAFhqRJBtesBmbzYl8QU8TvUqkOzBYeiQtqnFdH8V4vZsK
OquZlpObClfCOqL3HXF6T2ebvbGj76oj9ml/d85kem8hj05UkLGyX8/+EoJ1XQTC5lviJ7JtKs99
dAO8e7VWOW0am5btyT5v9ViHz2RL+nDII6RU++VzFe+k2bUChBbjEj+zg9Q6pEg7GvtrdtAnqoA3
g0MlJJpYxWuP41Kk+ceoI1d96JgdriTTLps9KrBTjEyx62qdH0zKqC/26BQxrD2oNLew+QCOOHVv
x3RLwBqlo/pUyLTENvMNFddAyYF9ZCHcuttXyS5cKD8WlzwvJYwY8mpWY/W7UO1ML0z4oVFDWN93
5ugjLANKvJb5FiBPsgxIIT8DHfah9OH+v1Abmjuwz1czG22F63+l5uyuA5fvnBFNFqXfWXtVj5WD
SpxaKcu7/bO2EY91k6fLshBJkTvuREv9tBeB5Vj91mJP5qBxWc95OHi0zT8beRGdRgY6wuxzOn7o
45MToEK3NRsrLYeR5WB0LBc0DGFdwBntkj6zuckIxtj6G6Qpg9MwjNEs/GJU51KlvUTEh1PUm+zO
bjn2xLvNF4a+XBv2rl8ffhFs9JDy7Hm+gm72agSIC2pX2rQfAm6ChW6aMPzLagw2guEEaxXM5KuS
doDHvdoZ2TFAzhzybEE6pFvWXUJ73Jz0FFf7SCHwdk/C3Ftt+GPanAfkYeKzcB7R/oXDhcRghfwx
GF4crOE8rJL3MBLcB83QIL038vLxJG90Z7SEQplIN0zhHpbS0Pvk6L5oHMhReatVWeqsjWUANR7d
i5Na4JAS5nEeuWGlOy1scyLZTbRqdPBz/mQOD+LURc9WTSxgc9/Ga3WEH7Wlrb31BLpgw1pGUAbk
1f/xGLhgLS8CAzMQuIUX5HUqOeqdc9bdfRMuanzoL64hi+RpCBAkReCbeSYziQgesfvI79GtMOuw
mFLVA8dqy73fgFYS9WuRgu26F3vSegZBsyMyjQV48BEYlDnbiHt21uY2SUMDwtQUkRhSjDlQPI55
RxZ145K3M4pRyi9SQfCsVK6IjsVEFqbn+P0PCw/Apw2ARAPznWLzvOsPM/EFMnAaXpe1nfm6k9vG
AYEWDX2entwzHn+ecd/0HkE6YmLiuGRB/sx9OwcPC8mYYZpJ6zoICAE3J2VocgF3tFfbGC5VcZyK
JDukz7CePs0jzHryGdHH8EJalwIhHlvJTBI4RLxpIzZIE9Bpjq0Zm4hiAFkt2UZCYJqNW+0HWb89
q6YElb9txM50U42R+VpwzjyeqJC2HGrfgiFZWu4LSzX+shMnukawggf3jrlKszID35HDBxLuD2VL
09ZtvrpRMi25S152jS6G88ekyoCw/m9uYTqu0/vDnj57dleCACthPnU9cPvbMm5oIuaEl52bKhkL
ec69IWK+5my/ta3sQx9+ljAw1reYnNARVhM4Rg7RUypto5lzlLslS/xaUbX68eUJy2IPCbFuIaZ3
EmA05ds76VqB9eY0GTuf8bacxeiSES7lHv31wlu7T5H1BcZ64WCxXpHW3R1283HwgPrEKFJ+aBaD
cxdY29Of3+b7nN2ZzFwmAVYiMWH8nLDHDdpkMGjUH4UML/4hCtxSsdc4yiu5F5+eq5owGgijuhdX
S8No938PQeVxVG3glEaorbsEgfygipdMJx4MbFZ7wikMBvRpZLy0nZpsZyTo3WEp/RRZQr4CRQqJ
8Mi8wZy1YqxGQBQQ1kQnXdbeW0cRLM9U1vTkJLLpass8e0vCDh1Hn1SkShelxq0Sm69CUVvpDQAf
Nxrfu571UYoihB2puUXuKo1V0YlNIYKJvAeyUi3Zzq7UMAzM6PAgT7mE1QUxWWyexWxzzS5hUe4J
EMv8xqEx3876vNM6cz+0dbvBYijL7TiSR5NeprGLWNF+czgOQFKyb7h0CGCTPB4VqiufsjmSN7pt
GhVu5wQmoUv4ETKH7nezi307YkunBtX8jyYEqPv165vLDZ3fESPUroxmbKdnq0FmFz9nNTvUBdYF
2LECLvwMWI3dY2XTLmaiiUpkdolzenxkiFpFgOSM/g5zlQQCSMPieLt1Q7lBFfbxjk5vy044Sj+s
TbiELg7Wt9vJU/TZW8/uHTV4Lw5YIHFFgaUe6k94C5w2bMQp21HMQQMGR/PkqJKEbmQzjqzAbw7+
uIerpC3nPlFCR1M1LqENyZjBIuht5XRWs9CYNRDoqXpWjB8IFtDmilryTyvDKwtA8OkgO/jehBx2
dJBxyIivNH2wudcwwOm7vIVifFIHz5ohQnjPIBptHYtoxePUu+1/Jxr2kI107an7hr215aBfxrUW
2sGipZO2a+Np8fqPZhE2lqzDRKWo0E7uCm4KKvWgvmUYkW5xwN3SQVQ0opL1L/SOCSCL+mcnmoFJ
b9WYQwbU8YRTQ/DaDjuTRRwU5cKWfoIh3s5tJJVjzu55uRxj8Ih2NoE70PF5/XiDA/j6fTqSh5tq
xf8K9it80uGvCQ6ymt5IZ58uZN0rMgj12n2VXb9L28I8+uGkq/2EsewPPccYxo8WiLLePqfTbI95
bvnSviPBrQHHL5nC5XsWJ9SozMW44TSZIi9+itwDL+odgcOqeTTrga5T4PMbrZP9Eot4IU/WGe4r
rF0ezGRqytJ/jEuATD7fGFGpmJ9DjxcUV65+0gSSyZg/EVi1827eP83WQlPJlygzfBj2Vi9FYmOx
hDyyXkXRD0X3qds8U3e30ifJUsbzeiiWqWIQtESE/m55xSoXk4JduNipq0xPbKtemEZP4C4xFZe5
vDlqEh3Vuf3nMpunjRBH+DfIBkrj2hx/dsP+xvZmjJNd3k7h2oTyNXkuPu+Rn/STQRlmjbQ8Njfz
tFKv28CheeVpNmyjbYMz0Vk5JN26fuEWHqDMxGl98ATPkHbrOV+uMISrvuXFGFSpM+kRraCxeGO7
iW2aLLKgsnS7i/zmkzBWCd6rSpQ7ysVU2rM5fExG8YA4jBMe0i8iV4SOGLAaXQ0tzRPZaQqb3qy2
v4Gl5/YfkqbVt27V8nr4PYR4dgN6ksfYaufPRpxCevIcV3/cLtQ7S7wJMyDhjScRFMd5VoaVYsFi
B2rU9X9aq/MHVpY9QrTVduP3GaReQZP3k7yaR4Fy/HqH7lERA1Qrrd3Up8FWGosu0KylXNbo+Yqq
xNjfvPFcg0LR9giOGGVhdRNUDCfke0iPzT5caIUGzJXLWIZqQEKZlFKWOc3GBVnWWIWMz8A4THPZ
mRUatvaPkIcCiW7M6jWuu0WvMG4Tetx0R3XzReTdOF8O7SYXYXKAYuBEqQRKQ6nAUB+vVhtkF8KF
uoakPdzEXlX9/FB/j/f2BeUgpyutDUUMgJz8LeDsvThEi+mMz7/vnMltQq21fjTqCBCTLCGp+zy6
9gFU3KHad/Y87bL56gPpxWMp6hDyLzwqNvCVSB00ZUIXw434UJGoENClnROm4/C0qbiXhetyzJEp
NJIXAQJX1hK93N8ZDYPFppjLV19/vcbRCL/RtxnD06/jHqMJvkMLuyLsG23iqboKEppbtOkFE4tD
kEiPjseEc4laRTsLDgn8UR4ovTuFhypAb7UxoOsDix2Jwjzh3JiF7pEkoCVud6tqaFAcDFHbHEro
Nm/xq6dbfC6XejlmpdiyAaMsOSu++MutoEBTGHvjQbc/1u3eUUT6Emp1t8t2ujbTFTXYwG3ipSD6
t6TjVWBnk33S4keN2+h9WhZ+NNfh1m89A+Ls4AZvo6fO2m5iLqWgMFUoAi/HoKe5x3m3SkiC0+nT
zLxkIi2WcRh5w8cEnhKxI+AlBQcNc/NxbKynRwp5cJBnj/illHNX6V0E7uyK9K2LyNpNn0eYOeAU
i1bZQAArJDAOlYqiMyBhR/PNMkqM5mWCdhGnC7UHrx92yt6Ytyj9ZV1fjaUJibsmUzpDnR3aCeHJ
uZk1uMm2Ar0RbyGO5AmdEF2TaiSW9/HAsdpIFSUZ3Hh39PbXV3w06VRmBe+qAeUM/i7MvkkvDOdy
Tl2NXmtLXCR0+ViwSZj5KNgaZ2smHFE4XJRA7f9L9KzaewJJKhRq/nmyBZWeBxy6oqetHFZQ7HUy
E04IztuepbGzq8TUoOuCSrLn6NICLesI9skDBEigccd4MM/EKOsQVL6s1N0M4AiX3s2XU5vu5A4G
MTu7yNlFFnQo5+olRe4NWSKBYQPhiJdHoXP5MvSb9i7Cu7MPhH88LZovDmtN958YULmhXqfRekNK
feZmbvK1vujSf2PYl65qvAGnBfLV0kBipuprwzSmod+iqhzrQzhR0+hMB85J1g0e1c8vjkrITbG0
dL0G+/4j+9rLbshxiZxNBC3djnBBDD0Vc4VwzW0b96GR7/uufGAHQRhgthYKc5LA1ENLwRCoPegH
jlxYSwBpKE17n2qB+ucO6EbbB/5RyNnhjquFEI4Z4AZKW6bJ4deqYJCzu58dGHMe/VAYXIYiGAtm
Gcbcs5DpQVXFanUO10slE6Y7OIQ/FvIQEd9s+22rMF6pGJXPr+CLTZRWM849YYH+Av5XPuPLnnuK
JjF47aE9vA5bCemOAx7CRiPesCxH79f0M6BarlyX0GcNSObPlJxl08hWlEEyPWRUx3KAW+MYw3WF
yqiMsH1HrLZcN4OVBmBXrtLIhxFVbCGsDd306ucWQULH5aBzRnoaxXQSWsnhhhJsMklLWNRWAfNK
zeexSqOIePLZckwr6u4GN4H3sbT0ELviWntYCPYCocPJxaBXgqbazpyTfeM2k1HePE5RcAlHQYOZ
6r+97pOrlOpAl9bjXruj2NBzKfX70/GOP9REFUwq+Y7QpjBOVTK/nucJ7ARcbb5L0YfBMO1D2pW8
jmNfqZ7oe8Za4RI/DAnbd2/yNTPuyd4BdWZtW4+OXl72yJuSYZyps3vqRLtBvHiuKJVcjw+b/aOS
g4u61ztcPw3shkYlGDbj/kRK1nPQNfB0D1WunN8ICdot4oX7NzGlWpUXGCf5n52zoGsLJCSuYeEP
Q6aotkme+aucweG76ObCYP6/yKWskZyht/SSfBpix1tO6vnVc5iiwZYWGkxdAD5HnBsSJxIEHg6V
WJh/7SzrAjkmifILyaAggYrAcSExsTh5a3u3smxc//yN8ff+vNNOZ2wijxpraI8jQ8UwHzswei9m
cYbBb9JjVfG5Qugye8T45ATw0kmDsaP/vYiBGWp+ijuqv1qXaS2KHb18019EXCefUYFvxiaQGj59
G05xzudb9LrZhguGawq64GCcqvF4BCkkI7l7gG0oTqEEkDBUoFGDsoonu1ZsbxKv1qlPcM20i+/H
PlcMnqn0lfGIo6mXYpLughmYWyySpE+gBYaLlBQHv24a56Qrd4+OQny+YYCmUfNtiW+IXDsokYEB
Dt9Vhyd0Tnh5RWsunLX9hl9TF3Cwkx6BoCltFb2keJS+gSl6x+gTAThsIbtQov8Z8I95HvdbYcMo
NR7zN3fc84/pm5Fl7LydOwoFP9/QQLmK8YaD5H2/jfe+cpSZZwv+zrpYQpjqeEGiVFYwFtT4iPp3
aT/TwD0BZM4IqqiUuEoGaKo0IxKD8XuYf1297C+LZOCY9YwznrHBL5tn+O+RNw4LanlfmpJVGoxC
rraYvUVujCQXaVx38HgobzUlS9oUiJjp1TGpK5pXJzPr77StpHg06lLean9TJKk2C93Jk5N23gfF
URM1+R+/IAWcuN3Pw+D/qDZKHob+NnZEjWSuzZ4MvplGeXqVLAHABFNwXGf8yaNccwtLW1+0i6q2
Y/uUlfUj4m/kAEDjGC/Gli8ZU7C48xoja/a3jlnsZ8lKmM7YcxWa7bC1IzlbR/7NXN3cd1mMZV91
6kdiE4RZY6AiKr4Y9qg2w7o4rhf9koQcC43/ieEKAPYk5d9qOXp1C032bL25W05hsC/Uglj/yEi/
6p3dy9r18Wwu5JWsNffQQcB75sCpq1aITQW7EaSLVt11GahaVnLGAkvwP+C0fcrMnAd7MK38ma9d
MSf9lpXQTZgmY5lCErt6dFsQZnnsXtJypnIakLFMfLxKWvkvhK0IS3yGJf8n5R2J/Z6hBLIB1P6t
50mxTKDWPBlCX+/v7ouJ6coUkr+HcGjYOXfd4FnSGFU9FP1NlGLCUcYZI8duSf2e4T0Fi5phzTbb
jdmtWThrFCz/BMdtlPfZjrLgUaAHEZOLmdJQ8qwBwn9owtqvCXleHlpgMhEpyHg2gZ53cYIIhozQ
Xh7m0MoUskS3fjrfr4BqruihYFqcMZOcF3gpMnWxPTZjkNrcsCTQ0PEWAZPfKXwVkhil+xhmKO6J
MBcbZxmmVkj3i/ZoYMQgtMCVpdOGavf8Dxd/dpV723MwxP9vUOFRU3Xin5jpCKt9VrekoHS6iPmy
UnD7YxpEANlGcpnzapBoRQ7jIpbEw03nbgr44fyK45qFS5KaGyMc8XYEpM9KnBgLiBngXlWUP/wd
yEoeEHggiZA/y9OI2JI/rWDFknUvlh0qdnjOT3RfidH7TyY1uPmWwwPTFqA9FDu4/D1ZsWYbaLxw
o4M+EDA7P9fvMLvOAmBbNcvZQiQpF/gpDqJ/3b1VAhYuspvJftuHkYXDjOAfDN7IoTfXIon98i9u
0o9pDeuOGfzgLrvpw2BSmqjtN9nsXs4yRHTWI4wQ7miufX9oDLKM932JeHKXgQDVDDFxPDpCmi3Q
yRQF5xqeLS0AdwlocUToXvKz51ApH4J5ipw3B/fzp1V52VVzBIiYo96wI8JjKtgFOkluiCUvLT8r
GFEovUIb8ifaGxQqB92YX21lwff2LO2JpwNmMNBo4cXNEE2FFzZU8sSCIET5YJR17SJTyakoJK+d
vq1QhJ3Ga9HQfnuwSFAxe6tlFH7PY6qgLABnZiFl5UDnl7J6OfN5Su0CroHKlstJa4JzRlO+H7eJ
8uZXSJGsS23cgjpie7eQ7r4cSwCiJQ3DMxTbpZY95OgasjbLiA/vOSe/cKxjy1htRJWeBfja+FVP
7HF+54aOEHNTRVukK/QGBAfOsiJfETLFgqUmYF+vei1STQIHiFwIK/QGifTdd+WjdjFWeyBsPa9y
2eEjrzDr5zmD3b5w8oo6dJwTuCB7D5by54c70rNkh8N/UILTlriMR+oDXz/Rk2IdBYt7avryit6q
8p35SwzJZLSyIPIhoJTKpjGaNprjQW1zcAW/u/V6ty8jUb7bpLfY/i6TCJQHG4UjU5Ao7yQxdrgf
j0QgPQXKXY79RFdiNlVIG4/R6N5OeegVbwrDa03Y02iI7DkNM4fXer7XD5921gVlhXAXapjsoTug
KligwcCyBW/0LaIbRlnA1f9oRiGdmwIYDi2Sh9x0RziteVptIok2FsiSVxMnP/+Bt9Xj5TbiYIkA
9nUdYqB/NtjPMYVuIs4lA1yVYHDoPLe1xhiRDtybFUJwenroUzLKbWX7vTUyIqEJeaNEjpbFWRwd
A9tG8cSildApXZKftWGNXrybJ1PDjzt1wDS9oQXdieXAbMZskK80bLDVDWN7NqQBRGdQzIM1dO31
c4gnLkHsHZ9nhWIBSt2l0XAYZ7NUsOkKeBTQYssuxnAGlEm86VauVkYuHCe44I3K0PgmsrpswHKX
7mHvu57tnj4hJm4KXnoxQHgGalhF82+FKDTFZSiWFTGHeUUAY6gPXZwPK1JUnvUDYGlYPsM/ISgt
BTteSMe3shYXqBSk0NKieLZJZS6368TPCsfWyTWpLiwTsL+SJTKqZAJ2mh7h90hYmq8I09GksuX8
l6+U7uznCf1Ul4cbDNz+Oj/Ytu40DF/euTF9o9SdWz3HvoaHFGxyiK8RQB7CA3F6H/l46GUKQ8yp
gTf1O3eZRhVKzERP5/stL1pXfYynSved76N1Q6u9RBRHd1Du3FM45LyE3AlBpgCSXwJvM0RqWEeb
U7P7diAH76FkJZeQZyASRfCn+hyJkx+zOCFqHAkZehVnH26Ev8eVtbvMK9qRVTfvmtGmZJEGYcmH
tVzL8vHQqQ2/MNXDM5x1haIej9IeLJY883vnrkFgHHXrVvsof56VG6oP7O1v7EcAStPLtQShVxQu
5b0vlO1JgMvgh6SslIWOmfvgGvFRVs0jwioxLlBKZDt3EgHM9qOCeRsJ9CFaHWOGiYE+XauNY+Zc
r4coE7xW1d5+A8NoyL5OraBn5hAJvCKDNVPEa15wyErMXSRzG+oZk7eih7KSvakHkUTw2aN00fo4
3h5i06hVt0La/+/bbBHOD3fI2LKIg0Xc/kJXu3NECUvBImjOKDlWeLEOXQNr2yJ9MQV+IISvbAMB
PbWbGlYGbXvsVdgwn1DLzN7Q7mUgaym73sbeZj8LnV26kxbmQgSeSfKJV4WfKiXuQVejHLDZOmWt
9/dFGUueZWDCyDRT3pESEu5hRvDNi5JGRU3oVTvpdDOEAmxQNb0p/iABy8RU8vU1ZpoOWtT3hil+
KlZzSdfzuDotW6nd5fB8gHnjwxE/ndfLBh+DIYja+95o72J/qqf3JtpElNnR5h1ejID8MfaGm9Ix
O5cEm8jaSwlcSjDD6F0O6u5ddNraEK2gwlBmiuzcM7fO+QGZUBXipEk5FttrID8+yVWvMpUwe6Eo
I1ndQQaUmUun4rcOLWcjNRq/72GswtRlCXHxVO1ykRt5cZVxsoMzQDZzPDujLHjK2atfQjwETawE
M7v4BBjGYN5EQoqIEwEn9XjXFshjjP65NLT2MgUVMz1OmSWe1TjNQ5Wwn8oHD3ur3BOa4W6Ibtnk
w5lw4elUen1590sPIFn22xQwwoWQnlAewW1mDC2ngeC+8IqiRX6q99dyWeFkWUCu1x+dv6P+jlWk
CybmP7CXQzCtKczYWL2+iQfK36ihH+vguJVAe52YoVpGsqAMQhjmh282E+IBsco76S8zPinOvWcb
avF8Ug1hrs4DWkftOZUn75kxsg8S6NcxP1p1FJW2UXQCMx4Vjy++Li8crbSiPIheeY+fA2Y0cgoc
w0rO8OaSJOyw/P20zvRyYr9bG6a3kYIwQsjzF96Kf6DkVE65s6yKb3KRepHHH7Z9ln4qu0orJAsV
d39kv/dB1flaCU9P/3TTAFSQVb5dnI5gARg/XktFjMluSs+RSyeK6hZiDDiFzYpOVZ09orggCT24
D421UI4Ein4VRz6lOHC8URO4Rlwo9L5gDiXNksSuHDJi/3Ydkv7dsKf+Zm328uadQ7lfxTD1mBdP
IcFBulOHBsz7uSqxp0eUiJ3/Q+hYcsFhGhZUVG9ZKDTT0SFsWzlZVjuWOhDL6g0ucvyNl2g4hiLm
xrqeoZAO00cfSiiNYgHtc3nDHSl+lAZg8Mx9kmf4ziaahItem6ILsRs28fCN44pn8yU7e+lPXbgK
1dnPLaY+RWgNOhEYrRaO90tzqmuWn2Oq4ZIaYER3Mw5GqZe6bNewYkIjgWPx3+uV+CA+qI+eP/6y
3C1IbouIT9g5TgMDBtlIb+MpkMUCsvLMlgZOfR1l+oKQfpeXvFTI/jxnL0jIJE3QxwKn9mlu5N/z
x0cChEHdWKHCl2DybeaUAbdp6CfP8FdPDTfyeLojxAnyYaBHW8R1/JO0MlyX6Z6mTnvuPGxdaQVd
UCa5WKr5HgTVyDchzHwXxtI39WJuTh2JkrCop+dK4MD7lfI/hL9pmMvjH4nyInc0OBSV7gTuqs1A
/O+5BYKV1SIXFzIcV+kZoONO+nodyjQjOwtTxco1X103OKkcgPnFf7boJTG6mQ0Sjzfp18vgLZbC
4LUNjAuEBlwwi5CAHdEQut7zgT63QA3VAIaa4lzQVIrf5QQ++HbSwBgk3Jhvyf8AHb+s+snSUCOJ
qwj6A6g0uhuNqFx95Nc224UVKMQhb7xxbuqLiKQKq5+GJOZJoEVQA0ebhGiB0j+hLg0gM7ZzyNeE
HDJhyHhNC3bXNyTrfzQD5u2iRwMB+8mEo5xXzWAOkNg62rloFr8IkoQdDeqhtydStpTXs9KLAeET
07TgiI7pEWZhmT0UaHi2L42WhcjGJcnaI7FuROn6Re4+6KBrTMsXURICke2InSaghH6hSSc07KHg
leWQepTdpWCGWgKY7h+agxtZtYMwyC/0qMnhosm6c/68wxuEYIOFfUeniPzxb0jt/frOQbeToRKU
Rh/hnFGEaya6kF6OACWyf70uNODrGJHT3GmrS1VIOwFmDgRovwrhjGn1ExjaE5mgyz8U+34tX9dj
kniI4A3FmMsWehnnEhZxvyVh0g7i3hJgnk6lf+zS+ItQwS5zr4duy1jnDEZ343VJ9mUzBSHAbZ03
SCEBOTX9IrMi+go9305ugrgai8/JzuoduFefJ11GI04+nGc6hKCVHJnz0+VK6tuVjWhSOiFdo8/o
lyMYP0ot0VJjdphxznUj4XU8IJ9WnbJCKv/wnmBTcMApXFHHgOMm5Hy2wANei0+Wx0C225y+ouom
YvZnZ4ANi1VyR76bs70/cGGJqgUNpC5fGtw7Wo7YL/k9jEX1MTlR7nYpNnjFGih8QK3dRcg2gmtm
CcvJmC2g+6oTp9CmzRsKQLpsDizKeYrRBcbJMNffsg/TPIRnrjUjfPz+7DctIY/z8QwsyR6SP5Mn
JvlKOy39tI0LliN2+JlaLjT7YL0GqwwNNA9mxVQQB1cz6A1yntzSz4De/Iz7TRzMfP091f+3ZrEp
J9iIX4ieQJnydj9MQvq6g9yLr0LV2dHn0KTxckfqxuALDXZwFlE0zZ5C0FF7q2CdXwemvlHmj5Uk
I93rNax0oKHJiNWrY40R3ySKj6D++kCMAhpILGK9XGmfEidmAszq8UKUT1CwPtbpKfxadfEo/yiP
1KjnQcig5gLLVw0I79tFt2ZpenCFY4SMsIR9KH56TQCbHR/0UZIfOs+q0BqvO65ztKFHqxaPnTSr
GiZ2f7LZbJqS4dNEeDTvo3W+kmrYOzAafkLgmRCY21ZChkag5PCAz6lZPcG+AoQZmSoihfT0FZ0u
a49UiRApbDxykQVh+13ug2Lifp1pgBgKB6qZdb6LUxIs/zbgarBsxoa1n/p/fiGTo6k/0vv8A+BI
EOJ3Kych62sKdp6OH2SzaxyUn7w8j95xa+5jJyTeSNrGNWSRh13RWsifA5EfiFxf0y8okz7UNjMl
UDfBjyHCFO0b4Yjm5D9wvhdE3983yd5w3fudctcFZBZogOJgdmzkuTrFC8iAS6cJerbxyKu/f5kj
njSr7MdFbQX8jcwL0vJUXEW9Wvp3W8/HcB7jQ/gC2QQWkR6o8wXrzVzz4JFNRzGqDTMG7u23ja3H
4pfgB7WTLjddNpBCbpKyPflzmVU/8I4e6JFadqAdhdshUgdx+zel6MIpoRG+U+sQ8avHdTbqN0Q7
el1qgkl2n6TNwXWA4t2rvxjWX3gEsg1EbY9gp2Ifq6VqIStgtsogXE1QWulg/2vdXqgm9BE+OTcC
yWtVM11jt380DwgcD7aWjoOV5oIY/H8jebqZstx5eKL9caxy1Zt3w631dFa9oSLhlx6LvjeDrCIt
YgMWA8vxKuR5WxkBiOX1fYpOHbLlJFk315x+1IxxDSNyGMupDAzssTPiorCbGHRRcRd8PlYhla65
Yg8kiTcSDCaHifa8xZteG3qTF26GOnMdQW2ehqhAa56OUyziiHzdjLyMKEXgq4mIYdY1JpUC4L6C
z1EGTj3MBjnd4VZgmkZ/McFmpN/Yn1/A9p00oLUfeBkiU78aEY3pEpzvSbmQn7WtTPzveXjvp4uC
foe668mrVdjcbs99NJEscHrbEX987fqwOG7pcISGJbKTHOy7qQzmCi630zqA6zJRSlmH93nYHJ95
JDbZT3cz3qhjBbUICgY8hSdJ2pnbi2fjSLPh9PYUZ53PXk2oNT/2yCBmdz4dcSZ1cPhymvUUC0tL
T6QDUEALCC6iMxkC4llaaFffWXEjc37jlSUx/drT+XCCIB9ja10Nyn36kGI0jwgh10MGUgfmMhJU
7lT9B0Ss+oLTX0nrtWi+aVRNQoF/UFx01Ld6dIm4MHIPbTIXn/Q9TeX/oU9hFayproRMjX5RBUFk
2leV7I1atr7SivLLcPKkqA9ngaUfvR5kFKMzijY0HeVuc68lyttl/Jw7hfvyr+7uuU9D0g4Y/NUc
0co4G9EJkcEPrvtFHqWkB5RcFTgTRz93CA+WLJTCfSkPMlp1MnsSUFUR1BYmq5OahmQtKmGoLR3S
fk50w+T4qNNTYh3dFX3rNcCoX2JqOAQUHS2ucjkUwN/t7uNOviGWdALho46TrBephjwEkp/yMcMF
PL/VHpMZqQoshlUUl6J7KVOcLojLLxeKO/dXlyOIHunMOMb5Ll8rdrV7vLJNiJHIqWwS1bFpac7g
zaTYA8/aXdYLVur66dKWP3bSPSM9B/gIip5FTuzh40DligFQi+jNlnhcUBsiaVAhqm3KhwbnzSi/
y/FBtmM+b+9nnvO/B+KVyd5L3mCLSZabAul4OF7WwDJtE8N+06VqvJ0sXVB3o3GgoJ/ofm8ruAv0
5ISw1RV92rHFQkMaPcqOrQSEeN0yI2KN5bJFscHfP4vnRpW7But5WqJ0coEt2Nwd9bgOFWZkjG55
AFWTMstwQP2VjG40XrVZJWBR44dMz4V+/h7HjAZ6+lWr4oDpbxJ8tF8p73kclum/8/FFriWSBJgS
6kNMW2BX3yBWal3uIQCmxFw6ASP5eLG0NZZdZA3nzbZ76Zsu49IVrcXyCoKkc/1epRE/euNuLF7g
fm86axknMTXN9pDcSyNM++hDZio/cPuap0v69qUkwyojfU7O0MMSeTRRE57hDt8vbjkUXxwUPp2l
re59tz49djt3jO8p3cgYFvj7VJSvV9DRpDlGJvUozQiEtM7KCoGQ+4/4lWzbEKs6OljjpuADb7ej
yN4kSmhBAOG9fX+gdNUR7GgQRushTC++5RpgN4r8chEHTVCOsb+iioCM1rlX051nraVqTINMB9hG
jMo/wZQ1uS2NnVkzx+X0q4/HcGnoaf8uvJNfMVHbSfN/zuDtG0i/op88DO8qbXf4aGvco5ZHdaHA
87ahFDAStIY00TbRk8Wbu7B3rl+03Sh7m4Sb6fkyFxhPMJgOCXe0Bqet4GuJevtR1/mTc+2h2bIu
8B5mxft2CvyMLNA7ZHBDy2fxxIk1ga8K/3o5P0Eo56azbKBsEcCv5GVICBI73KcFplFF7xKJgM7k
1OsaW8AR9Ge8L3jzwkHgC1cHZiqmrwUhg3YRJvHBATfMeczkq1NuxUL6gT9JTtPLt8fG2GU95+Tx
g6DbiRo3Mg3uvXzFLpsuDZd2EOCRLpoGPc4PKp+wlx4XaWu2937IAXU0K+MUOfN+Rblm6SvRR77w
u9hSbZjbP7vGdOJo/WQ7NAIN582T9Z7aYU/cYz5lWTeAzCba1TsGI0FrkN+4SxT+vMad5Ln/TpvF
dco1gh5blUQ+xp4f1OrIbgR8lXc5qXBkzS9O0GeOAu8uPPf122e0jc//TgZgyMi9RRGa8kFn9O7i
vwzEgDD21SFtqWp4GlN5+FmeBFC+9tBb9TdRdIOW1hR7oELv2MzI4kBYyDNld5KYqc7+dfQ1SgDR
VS3zVToE/n8pmW7qRVhr8OxNhGCnf1L5OyfcWZlvFpAO5jXbDE+/aq8g86mLiwCk0f/Douxic1ep
FfRt+2ppFU933qw+H1jVrVlH1x+mGpR6lrMGLjV/ANHe6CuOsQ1cw4VreK4nEAh+UDL6K+iL9WCR
yStYHwsOBAc9VoFnmHWhSo1XySSOuqwF1Rm6tAyNf06Ijqgoo7xMS17NSyrwytSl6mmNCIIvGS2h
oHCOCxdRo3Y32BR+2yT/hI7hC2ZZ87VtDdJ1ottcF0EgKHFUu4z732TMS/HbWuRJ/cQEmiKsfZLO
qQuzR0XLkbfnz7Yfk1kzfoi8g9RM6rdx6i1n5xydfBg5829M/hnFNg981dAepOY27hMN5wDFSczs
84IHWs5w4REeKmKzt4rLtlTJAQuGw9bCcN+i/QEiYMm2vZoUVBXFTEbEbFrlXdqrQ9+EPxmvMnkm
trapck0cJPsskm/aOTF7zfDVwJGPMl/CsPHU/iNb4bn6SX7KtcDdmeNY/MS/vHuHV73PoAURt1x4
Crzcj1xCGog0dPj/bcVr/NVQbUtnUUNImUqajrxt7QgWHehZBCW2cmiKW9PGT5kKzax3/hmvc4wv
wK4Wd+ltLu/AueGsfifkikHJlaqxxCmqIsjzzEY60XasuE5BmoJOALDUqzpFZRpKfQZyGRsHrwz1
LUzE3gn9SORu9Z+JH6hMYUgPOdsjj92mOyNMj4xv3z+zUcIPxvVZsuKpjQlYOZuBdfi1Azgun1n4
WtG2OrSvfiuUk4mWaGaqXhreLbVGMAmjFNWrM0xWvAfQu4OdEjZlK1YXnl7tUla2FUzWQhcQrpgx
57Ck3TIwe+Y6ephHWQ5IjyONVXbrYDKRSLXq1eiV6zJ1fv7yz92a4zJ5g2YCuHWxlQQFN+V31Nq9
pu08tBCE/aqBUIFKKagGozQVQx9s2Qys9kBPUqGo9IBstkXGAzHfMe4WFqr0c5lDRV/cIeepSEXT
AUon2RWqfB/RI5GRAZg37tM5jqIAgocW+bQVRhIZImJBBZRci8tPQex5MF1AbopiyXu3HNWC/Vz7
5aerKPKirETR34m13AR9zlmc6ucNYCPdnAZS2RyzlJDBfMkOxbM7ROY+UTJ8/Xv1OmfZtBQggeCe
qP8wg8aWNpBxE9JEyACCdfWANC55P9dX1M1Qx6AZsiwTPj2B0Qn9HwMIiiWIJWD7BTmfeDbaeJUj
PH+XChIsIryzXQgHv1KTZw9I4k7G/fCPgy29dXubTKJ8DbEeQ3QhkCi6F7iBkmYaeqtdn/NkluQ8
pG4Nwar3Bkpoq9wv8n/PQbTBBL+5rI+pzQLU2iX8Ub/UCjwn9a6NGqND6kNg4sx7Wgm+ySvxcR82
KusxA/vqZJglKuxISdo1YqgIS1g9bxCYB0A4XOt+15alHHfaPMgkhrVHEvEQYnrdvE5Kp6pVhKCx
Frv4k7BS9xjGg1fs+SNN2qjXCcCySE1SsQphayDPoMKw6Enm1VYS/s/vAFjBY9G0BQDldiuqoily
EjhDMn56fybr/tvg1qLTwVy9WwuW3qAdY2wchpuYzhPkVuDx/7lJhG0C0mt0M2yb/vOd5z1IAtLF
LWENGPoXAk7rlFOG5tSIh3q5YX2rvLwX+YvC/57q1xLLhsuUA/JgKj7kXPaEQDquEL7PG6RMF+aq
6TNr41RFAMPc5pu+2wXPp4viceZyfOSiyEorHgw0uVwiy5J7Sxv9P9gZy2HqKHvwTHpmm2X4A5bt
+NlxAIh7cOi4F5kn4Tes956Qqq2orgdJP0x4+o4KbQ49wcqmBkVXtJJrVAUEKBWEXxhxJwQPsdTo
iroUP3/jfhKtzpCMhyiCca6600mx7ChrFtXLcOAmqQUu705uXyxiuacUoEvQ5PH7OEGrCYH2KEkq
r43tIi81Q+qW9vwusoEdsxwk1BVhEC0zy9WDqReZRyPN4DyaxSTfBZBusZWzfWRc6K2xtiuTktL+
WMjxNCyy9Vpz4rehDE05fUfHIXWOU3DnwDYwQFe/bsYhGZ1xj9Va/cRQjpKdgPUB9P0EZr3OU42v
MWz9D/P1vgPqIzC9/vBiRVzE3Z/CKrCtx4l6jvJLZfCxl8sqvQ6hd7fnjJIUaLVwdUUhbuJbkl/8
KoS4vfnJ8lmb7tQsFSSThoDiP7buD+35W+njqtvHgNl3AcUFxPaXqX/Dbpeikm5zJoofQuCSZ6T0
3e2KC7bchYcyqeqEbFVok+tNcNL0bu2WH15mkiEzybdv+5TNjdJKc7G2jp8xIPqlum0nC4CkM6Qz
5iKQNbIyn7ItsFZs5knXaBAVHBQKlCX3a91oy4oowEUeGspj5UZACtdwXzFfjyocQBZj2bJZoZM5
wtwl+syptgoDz5wke0z4Oh6rmOfcSCzUIFI5/osDfEiaiyMZimBOXIU8UeHqTueHRlJUC9kypSOx
VuA1g/uRfoRYCKJpf9OTh+lgg+I3J8Hb0bY776Z1xHBilIraTFussNl/Ap8GhCZvIrhyq1FR6/Yz
RxHPLGrUYQqKcCnFVsMJSmgGjW5sAXOaJ8xvSAeIny9NdMgMWFLrayfBrmqFc2++nU9ZuzswI57y
n1UQALTWczVBYA3ZB07FLPMZEti3/DRVBnQNvw2qWzhjjXkAjgKra/eihDA4KMJibZWiItB/6X/4
R4zMgr1PnmU64wtYcU76nDlobfVApYuaTvLF6IAkMBYO+O2mVnGl3iJb5+/eX6c89JXd482ZqtVN
Y8gEuKAfKT3cZubWU/tWyyXepnmXfFzjvSYrQk95ItSdtpwoV/rkjLl/lRobGQKltUI0Robjs9aa
b1x1Rx9MNPi80v/9TdmsAVIhubkEc25F2LQbQu54qEBJ/6R47Y9utya5L1c38qASauqNmLGu1p8a
r6vd/+tZiIUdIYg7uxu5eHW5N/0uiHr4JuWfskspBWqYwAFIkTyU7p0MQ5b3qeSqrRD5+Gfdszs4
JnvH3wBlSFx2hmqgKZ2P3SiNudyHWyJ+Dbnrw3u1gyd6Mn9HkDa0C6nmliD9JqGs/ZXTgYmhkxgH
aeyPqiRvueXH6p6d/MFncVquNO5pXhM6NlsIR19d16GpUrOP6eNwtcRV6tPMlQmLepeX0KUP/VSK
W69xYvAG3WEFW4klyVHnO875ZkVlvUZ7DuX9xohxk55zP1MRY/RXpukIrQxzYRwovJeiqSuPccdg
aBLNGOBEnUQevCGjuxbpqXdi0RRHXOoepzNHE/sr7KsgrvIxLeJXLumiOmwji+BysYi+OcEUGcfU
gGJ+G+uF//IpaVuUIea/uujHAd/X0J1jeTPemgnTfJWOF6Buadd7RnPu0VLu+RxcN20fgcWognWp
QmwXdu740sF3zRiG3ToLl1rm4NagwZo5+dHwBaC7FLB76I4GK7dbIhIb9tMpbU/rq2Epu1JIvgg6
lJOxPbgIiI4Hx6ZMX0mI8vDqzeSbhsuwJzDCHAD2Ag6REV0mqug42h/liRvNDsiw2x2YtL0PIEMB
/7DWRJ4jkN6pMmEOlYxIAsnokwQ6crWCWVAOZnuKhW2yisLP8X5t43rRINRpWVU9SGubjkuJnFug
tr9x/Q6J2kCovMNmlrb4W6qqWxMddHXpMKms4JXUVudKhIfJ1BHlmTAmAVQ8z8eJFsI7OaMGEEoq
5/hlog0XfOXnWqxbWqrvFisl7CGJFRVCAZ54hTM9sAydM43blRiaYtZt3AymNRawAW1hNPU+foX7
FgPSBXdG3zzw2jUzvDdEiptaAQ5KDvOROq0sEImcgpXXP1NSP+7GTBmauKUbOjqgKuNy5b2X2IMi
TN9+9JJhwbZMyIBDqXd1JrB51NESZostmTTvcNWdofa4JyJC4vFziY11EgXRZGt4jgUq7mlI1r9P
s/m1FTksVCXFn/7b8BBzsRpH398UFQN/P1+91DztYdPela2FI8+4Vthq0+sGuvpklqk8+iTVPoWj
lj085LNreMqlrEmDgLeryyEXyOm3jMP70A4Nc4U9O3aogqNelk3zT/Zo8x/mty5WKYKJ/g9t8eI6
iLoXyUoOFLkJoOBsAcrn/TpQyhcxPsylqRgLzNutbPg6jKKuBd3u217x2GFiRnWmH5BNaQ5rf1ZI
ZtK78OhuD9g9KTzUBeTEVJQJsHtrcaXbHRZKYChqYJ7w+bYeFNXuL0SFxKAJE4PInZ+pfBSMv1e9
qWyog/p9X1TErWlm48S4fBeH1X2MepPbuIWmigTjn6zWrQ1r2tMwpCAIqOQefF80jceQjOTez9Cf
n1vc3c0nGn/4dTNLESbjcbrpp1eccihPhozzn7ctaOk0f8KPEGcMPqGNbbsm8CeImXTn6e65ScmI
lPxz0JrpAztKcUYvYsH1BVf0quuKiwQGlTYaDvKccKaAGGD7M+y3hXpxj4xCgThYiQgVRxQ9oix8
eTV9CKHa3HFm0Xn8RrjzcDLsgmWJlS4esEyo11pzEVpct7LpE6Hs5KoWXF2vCCeUFuI2YJJO9/bc
OKEg4h7H9RZ/JnP2MbX378nRpKqaMzHNNEAb+Rz11XdS0dVaizMM0Fbfk3lQEPSmo6sweIoyQZRC
kWRTbBu+SjUm31d3ofFFKuDh26lmeB6EfW2hbGaLSzNmZ1+dqb7m64pMUDxmPcUiHitClRzzpBQT
ehgSaitLHaXZZBggfXC7doTTFRDByG4+QwJDKSDqfdaoyKPvzrI/BPHsKkAEsaLUxdVL7xnND+lS
uFl6t7abzmQTfLPP1HAYLh1viPcKy2ywu5R7uQNu0xT8zeAcc+u2ZmZ2Oat72wSsm/x+SJ5JANwG
TnD8mK2EgFTTkxXxKnIL/wb7sFQ1OYwjhSPLmmNTiZSPYMJbOUqjri+fFsfJa+SzXboe9RZdFeSE
LxW3sjkOrv8FFrsXbTCAIg94rp7MRWMwPqt4LBekJEdi54W+Bx2TCxgoiyVAUhRB4uhaD4xoUsHd
AXBSHtorfXuHrTiBR74/8vDU+uJX7chlyVvmwKjCIo8UEh62aY8cA2jl8Z2xDv8b/X4aBl+qf+BW
clmZ++AdcAjDOv63EkCbCD5py1JJsQm8CKXP42t6CSVRxenr4vXhFRhFJUhFm4aCrspLSiXYj5vn
O9jEVk5FfVIqGjC4dwUTCxTXLwkXAMxDCqFU45OWKgDHMfn5Lp/ip8N3eRRcsL8nvPKovpunU3pU
PV7nZSTGAET1SpmO00muT46q3DNTqESEp+LAIyGq3ylDSKAuv9hmgkd9d1d9cgQ1tus502E/RcTG
32j4auYLavyomuDQE8JHdEVAeoUThU/XkES9XI/Ul0LniVRJV+ouhPtw1V64d35DYspDaS3RiJuz
V/zSjkf9Jg70bT4VfE9AqiafLOonFNYhVJu0hBORruIcDDRdYz1/xt24WWPJDm2SzjyBvk9gAxHg
i4q1L+XeXOUwSh9+9/43US0ofNsJX+yVSd5p4moIPk1RP/qVUJ6GL4zrpy0RdGScrQeZlTZbw6Ik
Rh/OKBYZ3HhDMUplNT/yqot4FbaKyA61nxXgm0MbFmgfFngLXEau0rcZsMRMVMkngr6vFPucvQeu
YLg9RaB+xjDL4QZ/NnGpMGQlYzxfev5pPlw/Md4ygNFveXDBW9k43OWQ5pGMZqk5FG+G6IBz9n86
6gA0tGJPNaWWNTJI3A/U+oTAXw0Ps8WGGCCoaqptRyE4OuXLWeHH7KId4usJaHfgyrR5yHb/fDug
emyn24MdA+9jCGhv5pkRdCLL2bSpmABaVQ5Qihk9Eu2x93mhW4D/3F4sH5Nze7BlECehabyWsJCS
ZQNBAg2R7q2B3BdFT5zjP56R9lR02hNSbGxU6mvIkrYT+40//iS86IESfmvkSbHMCuaCLtolX+cJ
D4/55/WMar8LYuVfihglHqJrSaapMKB+HFw2JbmGsRI8ZVhak74H3cPGTucStCJq+b7B6stPqOmr
Rw0Z6tch0SLmYMiCksa96FReLk438EjtW6vcJIg5hnjFq/cD1BN2u728kwj+4eupg2tMXxUemut/
L5ZAKmgfWSG3JpplH9vc4wCJWbnaeBGuh9sMisP42rRQt3dhz2Bdj/2SzH+jw1AzwyQP2ijDJsQg
OUgFkLzwkBwtqQPL/EUuRmYi3Aqzkfnj0enfwafWH0iFmfQ2h/W7BpnUNLdyR5UtAdN8qcaUxE7T
4fgaOAa0RSO/bc74n59GYgf/J8J70VJB+ialWuXrcgcWkzf0Q7RTZBZZmKS1/7ouFKYn+uY4ZvwE
zbTc3PEXfk3T1oh9IEwRjCODjAAlV+hyGRTFkQPIK8mXdNphV2E+/bRMZZ7J1Cfi86il8gIsFfnN
mBxyy307XzlOkWKCwVe/ikX0V3Kqz6U6z3S9SMesg2yAa95LJLwuQlPWbRjckYNu1eU8+m7Lh0Kl
mGXzlBWLuJOVElhYGtFBXfohLuMAIjNhcQCSV2xTXqjPSz/EqMHMJbvbQbfkBPrPB6eXCwjuw45W
7hvwM2WtO49NuYdiLo6TMSCr51sRT/CSwyVgswAVQqiFaxhTrDjYBaabZ6oXsa7HU+2cmYWD2oc0
buKm4KuIufnLQ9KVfgJI/K7uHOKpP3bW12IIn9orjatdef8WCEkFzJ/6qbW/MIS1fX38cQswbnaL
kXjKq23kjMEGS/vJfog0vROP26Xgt1kmn5NBYmMrDwxnACQNXDpQmOV7Iq8ciRzrUsJ0LSU2jwQX
YDSNtAX1eioKGLG1/1DWi1UYYDbsif7gLEFBkJ1ZS4IF57sPbQbLjWZDDxLCTfG2oziUuaP/hISO
JbOd8G44ymsabWZXR83sXZ2Zd9TToWosK/x0NwVV75pyZyAzHkV9hJj/0JdDgh4QUoZdwuQiMDMb
HU1C88/a3S8sXwStdw/dMvgNBghGTARhEYNePqKu/Q8QrpNGCRdppfV8VDxcNv/IBiJKC4ov/qDn
1NRnMu0FzMYQVLkOkC4TzaQWs8CydTjCtrObHfWKZfz23pcEbO7QMqIFAVQ8LbUsQY40/BH3vI+0
xaRTpAaMnLdXS/1qHTx/BqFHvtxOeapMOSBDEHe04lyA5l4scdTlXJq3MzX12vbOC8l9LudVPRnm
z2QLXjIz+fc9t9IcX4TibS5aNbXRsdeGEF6leyV5Qyi3WU5BAZdtRApCxe99HZDR3+CyCl8AAzLX
JM2CouQWzglhtzBUf1ZOefo2c2uO7nnid/tNcEKSARVv5beprlLoLhCqhuz0pjs/K0uzYbNR7Vro
pyxzLlsURTX4HNzwnW8OZyaRQPS19FfNbhjQ0uOAXFpuHfHMPRTKIGLU0oSC2gCrWvXLqrACPXFb
8fW7F5r5HyOZWtOV93SW+kPIPtkiP0QG5S9JbjyfN3ngr5myzFK00m5++hvnvF14wvI7VmAtKQCf
2iQD46b32XlR/7luMZjtV74qPxtoJ90K75NHeKp/QqN10StVoi7Snh81kmvbYIguqddbxm4u8ecD
gVr/P1KPRoziYrKdN4ae4HNTJWCU50YzE3DbaBWmyfRnyg8NCgiQPScYmqOtHgg0TmTBUUSfnGud
eVO+2/6Tv5MzCTys9d/quEx/hHdgeXV1JKRAAoun+o5T4hkgHNLiRQcmaTnyKQ4XIo0BHR31KXAs
vb43K2ND6TNq6nuIizrIoABrp0OkjU0aV4G4beNuyfqR2CrYh2lt4mrQMOMX/F4xGyW1FSeZIIFz
fLxDeHnSSmX4hdhCEZN6laeji/1OYlHEU70RfGiq9PElfS+aTuy4s/gDRq9ByiqBeSsM2eUJt/Jb
vul19lFidNT1SuLP5URgZVhf0UXdrG6umiLb9Y+aWs7rceEtsbqneq/mseoMfVhxWP5vqdLqIywi
rCMqf9zkW0XPUL13vgic9SGEUymK5KCMcmx5vSJbCHvqnfQUqI+RTWHSq64aIWhYE4rbRgPtPUff
6tA/Wyn2y/x2CAG0Xg3ZI4iLgL4Bmlyhujpy8QlnkSSbNpJwp/DXdXQs5AJj4mJmFyQTKf6E5+zQ
HEwEAW/HcvLPC2S7K+aeIPm9sbpEWae8jgEERSqY2kL9tMg9vpRfmjLX/9ecLofg8gDN2jXkzLGx
xPnM2Wq4Ft2UMlenp33C+Tdr86nb4Fq3bA0umm8pjXSDjrIT5fje8tjAefkBKm4MUs1X6BzLFUOE
OOJ4biEwzyWRGyWVdUOHk/ERxyAK2xDChEopcYk2bfJcllYoBuR4UUo25ljnqa8/thOrCYV/EaF4
rctlyYGQ2hfR01uidYciuIxemgCzcpRBXVG69vYrBJFrleoLnNGJfw3X5klKFCwj1EI5SucY+4Zm
k4IWsg7Gw4HW/yyw3Qqb50y40inOclHFVPFNVQTBBY/TiNCwGC8Z35FLgoU5yDIZ95D/NTN9lk7m
Bs117hNElQVUhj4Tt5PRCNatBVyysquNU27YQAglww5R+F/j4d1QjEhkVt0kd25I8M0lMLKygAfW
+gwhEP1gukizpvhuXNMoWDoPDjqUeIJj96c402+t+JAucsNqtDkCkw87QQSc0q9rABRTf+AfDYag
XT+RZ8l/Q9GqwOz51ku6sxxLmKGN1pfizbp5JMaGL2IKTi9NOAOJpv+D88mrG3nZFRECVrZN2gWu
CYObQbjpyFBf/zOewDV0tMw7m1uMjF1BP1RGueVmg/VqBqi6tvZw40agVZ9fXc/C2m5sSFQeHBPF
GTeakhak5Vfx2a68Q//UWHyKEfHQrZU7brKSAnXG/l7D2ZYJ9D95EhWOuwSincHg7CZ/QevBt/NC
h5/lxtrNoMdrZE1ZO9eD2mx9efr5ZZw4wi++zIcifeNhe1QJYQ03T2kvb2j6ykn6UtUVxoC3xtaA
X7ava4tHukMoJtnDxFOI5aGnS7S+lMstnaIXc2j4TiC20PM9wOH79Si7+iU5P21aR9YS6Td1yw7h
TDGwkCVM0qrBSu+lByCrg/eYRuIgix/d5GTaFCzekLB06BYcDBIxprpaZcuwXW+Yo6RLjDoBqpRB
a9vtc9NLJIkKOPgzR0jsD8/0HI/gXotmozv2Z7yFcVe4MsIUKSVyU8W6vpx9gCChX1sw6/ES3ZYC
3cZHm+54WI9LLbhKUBh9cRoikXgRyvNI/Ujrs9BFgyjHJZvZvOVE0oyffpZIOVz1EBktz+vdH5K3
VC+FB56q6y7jz7FIyo/bLhG0V1VeA7quVjhec+M29tyYeFkuAnmgGZHmduydCFM147e1GsCLN2rv
LKkC1zQsASW4B9Ok+vY1T1kpRfpmqhE1Ki1afNkCA7oCDoq/HD2LrCsSmgbeTEBfxb9KJSMV8YEX
u1jir16DNxXqPNDqitV/ims2ygUJ5Wb+3+Kq0WYw2IMqxPE5eK5pMUTIUJxE4z4AJi2GYkBbNuoz
XjEFA5bLmUJWQU3NW3xI/hrPJp8wjf4bwsrZzv3dxYe8A7eEr9EezwrGKKc/8bmSI1DyC7O5HYbU
B9zYRSMuGemDk0HYpGuXDEilBjbKBJLsnqiCIxVNeb8X0UR/WPqgHNe0fny47kE0AbiWjbXS09ik
xELnOrlbWJmD/hYATmQMp7kS0m1F3SG8XTRyLszUigID9B40yiBMnzwhcwSc3MMRQd2YDcDsPaPO
51HiOTfoWT7AJ1wyfhBT5FhrFKCq9K3Av9VVkm2ERj4FQs45U8nGV2P7Z2I7Es9L7IAsfp8bijl6
HM8Ccnis5aNMKTTZHvlSHuBiywjTJBE4Zsplx3ibfE37JzoKpHBg4nhj05THZ+V2GYq5JSUEiQfP
WxDhK0TTlC6j5R6Ge7g2Dn2Njd/a+SFBjRGAx2UyZ9bV/whvTLBgBuv+U2uYoqqrVD51Zx21eRt7
BDIn/M5lhc3tdJ9oN+W+YrKkVgaWE3xHENJroO542gX7rx1jmQMRPJBFBKd8LfUcU44lrb9YQxIM
InFUJ8L0+1jjZEM7/aM9nCUAW54NgeXQT/vF52nEGxphTqV9TigQjeUKo35Jam0y5tDZjGQZW6G0
YW33Fst5ido5PxhYp+TjmDZioUgUdqTutshbyKXFtPG9a0m45n6y11+eTq+q26RTnOjVOMI3xwGt
VEtvl5JIAkyEQHDCA4PYl4vR62G36WRfQC795AFeg74qhcewENyRvISsV51+3LSavCD4+46HI2tj
52CDY9hJc65It98AYXAnmpgcMgTxDR69YtcfZFuHGBJkE6eI1Xnh/9Q7HCxGwAfFjg0aZG4P9avS
uGb5oPhBen2dwbYGdNA1v53fpViZa1Hnu0EnGxbAXsywUhYb0ApD6b2KH5OW1g9rjWQW6DGiqoKn
/kfpI4ZEb+Hq/zWgBIVNHgEyxq/M7K1jv7qsPlFZ2d1fK1RcaS0pqBNbvopMzpN2cmD6v6RJKH+5
/SLKt7GjqoccZsz4vmHQZVRDGkXRUMGY9UGa4sGGA6oS/kPaaeNe3ap5nH75rnTkk0Sc7M2f2gmU
IpyhmDLRe48/s5h7KzrCdz2OtAwsQUr8R9vtvrzvrcjJioME6wFPMPWKCvDHbWcTPqkprqd6/TpR
betQ0QTGY92OXQ5eYFVxJC5TQ4riRpnoDopVsZah1F1WL6NbLYlnMXhI880wylWz0HJqUC3qcKhk
xmljOid9MH+ZiQ/PDvaHNP8G46LMaiEGB90QUc7lnDSMw8Yz7jo/pnQEq/llApremxePnUDaEGvD
qHcr18PFzOsLPB6nXAH2O6vQkw87AKboi8h8YJGtNdQW4LtgqfUUzvUkgTzZbe1RylcQC28ehYLQ
/+n/5pZAWBt2O3ml0PdZtaRiisSYqUC8RzYPeqluQLD6E9SbBDYHFfUxnR6MXDWklfxdiToik/LY
lm/7q4nNi7rRnYw9GdLsiA9b03aEvPzNHLyQBMeSrGERXmluhvBDg+xka9cuux7abqwZzRCyVuXk
dXdqbNb2CLTJEmZBNH5sJUbQ3CQQDwxP65Ig9et/BBtg3Kh3jAEpvY6x5Xet8+yPZDwyqByuT4tb
McLdF8CwYqdVFP16z4wlhh8s54wSi0NfLGzkiV+RY4usO8k6JOt2I8gF8YD6LGNxDz6z9rN3/C0a
fje5PyksqelLUjgbbR8XgRVOuOdo7gio565Fx5Wl60R5kP28Vh58483UfwEx1HFJNzCyDiEV3/N2
rTfVfXedcunIIeULalYGZf9/tCaJZ9Pq/fy3QmjIWJtliE/icFACMuqlHF77NbNn550PNlSLqkgT
UuVnq9PF6RYSN5Yz2LgVJQl/RQ5PDxgZiKSprV+yM7MKTr+TNa5U9W7hNcqFxGCqJYBdAgOK+11n
WZe3lUE4jVcGdCmFN6pbP8SpeoZbpkmfH8/e+n8MX13EaGM/95x4rNZHMWqRH0UB/1a9mgwq4g4Q
hbTxVeRREwCLok2bddWrcEs41UUzHiFrCaFBuNBSPRKynQ6RB5WQOLcZO1R2qj248PglUuOinFEl
km6hl5EQ95UdJjVqSsBKol8HfO9huEbRRl9QcOO1Pq7Fk7fTsNRrjpZsc8VLrWiGhd4jz3PvymX6
5e4FY55FwGmPzhoKEOMMVWr+14lRTwWkN3Fs8sritXtSbiiCB6naOKhuthyGyKUkBQc4A7KmZFgl
CSaue7OhNuZ17EwM6Qg3GNIsH6Xke3+V57naD9OSQyxi1IwHZbE5AyQxdXTDv4K35hwofBgUmhJ6
MBV9+xHBkauAtRpbEN5dM41gHNjDF6z3xkFEYENhmWFFqZ6LPGRbr/biBTn7Nr2jXcM2URgZI8yz
rhAZTRDteJmPnjo1b7lsQtp6GGeO50OxhTjkHhl0ene31KbPbFiILDKaVqQAp9uy6Yymm3lWIGQ4
3fjKUC5pT2dRiobojfIBQ1R+N0BuR2PyLgL5XcSIzIY2MlVMXTEb14NmcpPukrfES5TBMCcCO8QN
lc56igxH+QdMSJEsjb/eunvJKvDuMILk2jGzPKFYiHty3BT0Or3BYbpX1c4WCgZWRKF062eaF7rw
k4CLLnOt8W2BJmhdACddpeAY1jqP/FX7de21/ukNwnVHpeVg8FaS4T0OUIpGQu4RZHSpT1kFmotw
6tTDV3PDw4vOmB/uQbImorxnKYXDAyfLpz4u76EyuCYAi8lbCuVMmZJ9+dpqjchrk5z1BOK7qaU7
ip04n3SnwPdyzN5PTg9Q7oQo5ZoSdXGj9xgFHgbQXlGrZZpOyUbit18F9o8ULsh+IKciSQlFqa13
cF6dbse53cvvhuGqk87z7NQRuLnjyyVGiaSGPP3noa4o1xYFIAm2Q9FvM5wFW1JfNiHDEkslCjKv
YwDHk7KZr1ALpYDsu+dXATC1EFcrjNinLOOOFPF3/Udw+pjbsP1HmzPCoXM4Tpwp0DVSuedkYX4x
Fxv5PVs4CZ3wlesLJIcD79Qpd++W97h9mYrx7gEnxNgAIP8i1YqtNRbT9D+YE8Jgtl1WH6KKcZhZ
nl2zccgZSp3oyjHcqJ+s3puVSiPu+hI00nexPKXwoqhYtDcJQo51fEzgiATb8b4oHNuZ+879uWT3
KPQwOVTzNE4h1BR6BgLH5A+djCuxdeKsl+rXMPTcz1wBGF/87sQ2HWWdYEL+sOrG71+Hsb4OV3R6
OxfR01JbIlgwWMVvlBBqThWBTianUi17CjAAkGkg45fpbAMPtQLwYRzTWSo/tIYlZwaxIT+p0gFj
j0bs/FkD7Lc1Zy6I7yJp7Jw2tcINlSMfNWw3pyHehduLleLpPCNO7xoyHdHZXOSDCTXSCBGZWcQL
EXISxxMeUqbsSRalbvka7Cx7ZhpFWTd7J/ZyUThj45zwea9i3MucnZXoOMqLR/18ONm8OOYmsYMm
sxKs4Xmq+uq4wW1rgUggAlDwgxDgQjvBueVrOwRWzl7lLVYxkYsB8zQxa1mdrM9ixQjG5v8OUhBP
BQ25wwSvfWvrUzMeQ6/4vXZcnuaLXL81d7Th9r9qwH5WhoS0Jw9JEFklTJsPLWLsc9ypLZCh75Hq
726R7gN1Iniu4HkC6uBngXakg7jwAMmIa8i03R83E/n90b976rD9/BbXQlebtE+Xd9oPqUY+QFiB
/okRnsVnsMp71r6X8pRIFjU4lC6wNlkb9+Yiff9olWaFscBBioMWi8yKvZFETLBtQEpA6IZbnJFG
/yXfuwlvq/0AjKBEjzSlFEtUGuLKS+A9fesOfWtl5bUFL/oCQbyvm82+331s+5y180JC4fLbX0vS
6dwM1O5f6dhX57BDS054Zyx9s7u1xN6WpqsJEbCXMBwGhnynQnV+h4gh00YOkstP73lw5FzlDZbS
Z3vWW8tg0RCTmVV3d/Adkft7tcIpBmd1OAHFGBK5TYmkDdgKPOc/askxOv4IVB7N1aNAlYjU/dbq
yNI9mVo8PERPcL1m8ajdIy+p3nqidJxPBjgQ6bWC/U9qDIYi+Urlxvh13QVDCXFFxE17nofk+hjO
JiQPsopnjREgaiI4N/qbjPZ4NIu+mvv+CjB4bntaAkJzBbmGAdXi0WQUjFSQ0yfD9EkqvSzHTNpX
d1u1HU4Zx4TSObuBJKbwvfiifhyzHhHhoUgDLla9M9yn1u1xdX7aDy/+0iA+Wblq6wa7F7tMYhfT
ihv8NUhmbzQXFMQ2JfGZLf2iIibF2a3a+1VilLPPEg84+xj8cnpCBU4c6HPEdlWyt4kUMlvg4Jel
ZJiUOlqIDeGNLixTStaP1Sak8e8PVBnmhPqETG7oIBUzitxkO2tGuQORQHBOmUshDU0g6BxSgI66
V+FpfWsni8UVcPc4vIMR++DjVnglAWPKgGLL0aZINDr/VRvvikuBDos1raXOvXemNRm+CFSIHthQ
HjQpf+IZp934XLsdWdIEAh+7P0z3AGPOFxJZQrh5dIrn8tIKTbDKXViEyJI0hVsIxPqYUTfFrjJD
DiIb3s+5lp7+zxTxl3A+ctljCBq3kzL38YZtulmFuMNtmcvKO3ppJzyC5PfRNYCdFObidI2hWBSo
M9b2fMjlbhznByS/m3UOfit3qg9bpw9us5i2vooxxVhAdCIrCsOPxBU30xMcbnhpMQNDbWUPXOuE
qEI/mHNqf9rP6/lLEVusU0DMkhLVMcVVcqes+YSOzpxlqsnhhqHy8z8Q52bsF7R5bNbbxbKoZe6z
4/tkGC+FV8/CXM6sAUBma0iZ3/HGZe2K0CgeoEF4UVXh0AhBA+dB3l5qxkBownHeMZUAk+oi/Ww3
vp6mT4lv8iBzCx6zpvZfT3RpWbqFA2ik3QKRW7yJBc1tRamtFf0xV1KEaxYSM9Pz85wGss6Y2HNb
Ehy0ssYT94BA+13WcCHdeZOe5ZE/SNflZiqG1xG8zqYnAZypN2Q2JP+mOISO/KbblbCuwqTGLcbQ
rTU4yAefr8w7X6blj4h6aSAvSXw+Hl5Wbz30rHEBhP0ujGqDXk8DcgVcwcBdeoxu6d3pqCjyu+L+
C+s40hkOAgU4VWJlV8Hr3SKUWRwtGXmkGg5kGN2AmBUK7CwdUdiPzil4wYe9XyF0iyRErx+rtVPF
qCdpCDgaSgYHmRNFpAyjjVqO3tq6nGFeIGrBrnEnz92Ba74Pny2dNQivt1gWoaH4edF3q1h3mijG
qS7bEXa0t06Ibdyoe12TWF4phexQsKZm7Np+L7lPI/BDUIxO48eC4jZ8ItrpcckBnoI5mNkW5SKY
h7ZxVm5cHTQQkmLBq6S28GyfeFXZJ1B3TtYdcOtC55Wi3c/lPsNzppj9JrVekkYCwdSJ7JHfGz3X
0adUjtMfEwBQ+RoqTa19ZNExfl4LZsEtakrUHT0aNkQgRDUw4LQVqD9JFjBjWhOi6VkgZZj3dRU3
7yHDQLERdoR2wVgjBn+0G9w3TJPXVAS6mm6zRqpMS7Dynj/biireAhl6fPnkYPfEmlKUX6mnzd0Z
SoFuTjjuQAWtW5cgW38pEpEF/kSLIcFIzacnVmk3T6MKRhrWtk+FMxyzRR63xYoy2Rteif7eX7ZM
itdREDl33y2Lwru1F+JaMhxt6of6UEvfYyORI12A+qQ3+nvXAX5la7eskBXABmub4ljA1R/ORq9R
V0idmUP+wavbC8f11BqDtuD1ZyYvNeksQl8riUhqCa9m3JMedJYe95KSOEHrvkqlXbGKRY3v09bi
5r7L07WQ7mppD2AdoGy/MAT5PgXostLeor9QHY4Ve+DedcDwNOMtB+vdzzbKGmzXwzbsSkMa9ZqY
xxMl2YaAumWEgvVHeYjcm9PcldE9qeWF6QILQlwpTJzxajCkBx94gxaQtFr7OD7TFVS98h9FlVLI
UMut7DBoT9a3nkw5nve/f96A88AD27WxmEHAGQ06bSRv4KsiHIIkHErFXYXPOl45ALFQ6+ji/W8E
vazXL4/uHDuVxhuqgEd7I+iY4LcQhOtCYtbDrGDD7+EpQyFpGQAHaT1lKeuCAYkfA0t7G7kPGpLD
eOzEfMuuPJRO0NRIBwy19ocO8h67NLLAycWVeIPbRfLx5zycwjRfIl/ssM10utUHj+FlpqyLwj6r
QGSd+PhwDuHT8GE1AIzL2PHKKkJzlmaiji9rleQHAokhjdkOv93OuqMegPDYo5UocM2OlPVa3VdI
+SMXsg7wuLeqb7hoDoFwFpdy7AZvEG+CgJE19TZcja7c1Oza3cax0kQWv0w4JNxF5PE/RCIsi+OF
7kyCPJDAKGumUrJwPVfnHxyooCHvNejOiQFnKLmTZGXYT4bQkwrO68Tvb2+vFB6jHMyaSWAJv3LU
5TZbnMh+PyaTPRFUw1WWtLqaXDJeDle4Rpgi+ljQr4RKK8ZCn5KCSGrRiU34UprQqULiHmXTGYhF
OcVmEVw4L8PMHg9qwhR6OaD2zdrcW7v2M8ckrbUWVdm3Jdt6mqpTv0h0vf0o71FmkZhttoreQTJd
yiyiWqBTIBxSeiA/RZyYnrW9BcfsaRXEFnpaPictyV/2FRm4LDjZU6KAxXZmUOE/aeFQQ8EAh7df
K9VWDEnywSzYocS7rPgLINjxbysNdv2+KcA30HZo/H29cGpagho4mEf3zn3kSXjIJfQaron2lckx
5nFRtIiTPXS4LDXMF3rK2wcJ6d2x3xL87cEjlQZQqSH2o4/UKwwpymuuNsZqXs911YzPw/fSFwUG
a6kMnCmsapH9T8qT8Wu5IPsD2lgAhKLpMHe5XSsMx6nuQEDJyaRWTv97hS+LXNzkJjGpwnbesS/+
T1+1hK20RCtPmb/IPPhPTVuJOKlkhsbUhWLRCzdqzcH9ExgmWIgUT/PSNi+vLF9YwFRu4JGp7j3e
ivE67IT6isc9YJ11KjqOAKyP+lBX+9hjR/nzfphSECQjlG/dMPMISpEhEgWqVfpQxvaU9xVDjzCV
cdrgZA0bkVBZpVQpMrlqwMAOgWB6vykMF02sf82H6htA9YuLv1udvMWTv5IS7o19wnM9HHhSr2du
LymI2APSFEIRnR7W7gLOA6shKyRUybyX7wDyT+O+vXYaUJjk5NT4AZn2VoCw937af8DOVLbzhemn
Hj6C1dNEMHIF9LpYL0wMAKn+rwh1IiGXoLXT7bejLd96rEFwnEZKP8iglCp8+7Bpht+WNiWsJnPO
je4tIORKAGX3wwEQmx1sRdgLA+2Hh7WPhEquygDG+eam8tgS9n8Hk8Eubdgz8HFWnjSbRYnzSDla
DiyKQh9zg8+nwPCW48JODs22Aj+Ru1SthY2xiiY5oNw7/Xg1d7vuJ+2S7qp3zsltPl2K7HwPcmgA
dRHUlMQKdTtbaen0P0b19GkOx+ql4n9yDOHsX5qhevFnMz073OU2NKsNE+NVmAH0jg3Kl4AdcjCx
Aj+V41c3kc/uT0nMcUhvbW5cilPvf581l2+KmuPQF0KWmen0lK/+rLHjZT44s3JByArBbsWNfAoc
Mm/67LrWisbsmaf/Ke4jiMEZP2l9v5xDTbaoectLMI6vZRQfqaq+5iZO16PqfnAiHjErGB9fpTKG
j/++XsRx6C2I0H/KIdZNTQ6R9sbLK6YN/tKLUIGRB3KjZyw4ubwT3MUxgUSALyyzB70vznPCAD6Q
Aazq/DkvVfu/8HttlpfGwS62EiQnmP5jE6AO83M5onzCWPUsTlIxccaEf/DYUWvuqi1VZz9WBsfa
Tej5gkIQ4hhb3bO0zQZPTCh09t/66tab0V0xWJw8kCP/BTYJe89fXlCYEevOLc/WjLRu6zyehQpU
MgyhPlVy9cDKWeXTNcuqEqeN47R56pmio3X+9HkobFdK4zzVo/q8uEB7NzByKXCXkpPYBw9RHyCk
cogtPoBSHuZgOkZ7/p8SFLW57Bc0dRoe8rWhqByHZFqPjfGNOsbzfectdFGTJd98ANxXgxU3KLG/
Cxnb9rQBi+kQEFadx8oOfIzTEW7htNrBRzT7hli3gKZNVE+mOKlvgTaJWNonyT5pI0XgVLLQqZgj
+4jG2rwGKwJ88Z0Op6gmAK47/BET38jTpIQTPDKBtv/LTkQGq7nNdh4SSulb00KI6WaRmA2cA4Dr
wd2bfus+ro8QVVG0EhqI3CxThsTeROAvQOWCy7+dXaawhr8BJQJq2Xtyq10d52dQoWAKzBxlc1HF
yzcNTzxivSN2rfHEEkEWzEusEL4kt739Xl7BU5WBmEGDvQbDRpgAyLukzej3djNjw6IIc6cFIzHn
TwnQt22nhoptom7c8Z8wdWQ+MVJxxg5mcSKCusBXjz80jkxC3tB03CoFP6cNsu6RZZPBE6aAdLxo
Hip42fHTHb+XmLAGbYsUR3IGd1AbwFrVUZDp8i60Nfg53YiwuxPARiiDTrkz223JaMxmt3OdEDse
+SV9ShuXo4ovlaU3RXOpojPRWBptqcqfhqhD49xAn+4LK6c83MMxF8jc5pVYSfheLIsnbAxwvF+N
OmjRJKlL4E69i9/ygBBOh4QYBTFcifTNQ3srv4eOlNjDd46FHIBsNb/bF7TVzRtHUSjD26qJgfpn
/Rk7Mf6qTFOLniZFznd3+z25nQaY5k7FGBvADuqnR16Y5euRA1AmMEyXNF/h9zfh8g1FH1ObL8+x
kr8HSwA2G6eE3Lm71UabI3is/6ald2AZsnR65Z2wdC+UftwYanCW6Sp7RI0r1KmftpenQApC30hh
Umf6wTk0tCu+iP7y/pbf+7BNqIRjtZklu2BB46xvvjMLsXsyhC6nqqwZSeL/uXVO2D6KoLG+MGmg
NJCjkaVxGqiuaoH1RoKKKoaTD0WDTw1bXoLzgvSBtZrVK7PNyb+wwAqQEIeqz6t7hhAs8P2dfE9c
xpC0HNnbAWhs7YQrzqVh9rh2FRkNDNQE66WxI9whx73JxOiZOrgvE26N2qhwXGAF6nrdAtmb7loA
0SjhWOfbbHuXVTUAXRcPSSg0NCBPTBGeSrkwKaltM/8Qh27ZdSFrYrW+JcGdOjE/3LhW6i3Yabc2
PqfQInEzRn459HGhSoviBUvRP6O/d9tOagWBTJZwJjPG2IBbmhjWSJHDak5GetFlkKK3QuXVIQjq
++buDiaCYh1vopdVdWn72aXVy6YAL+kik4d6eYFUyiwjNwrFPhHzCAc0XkNGFjiMjTSwugxyK26L
B0ijN9MIvKY5oGbJ4PTHzk6DYKGmTrChxeZdayXJlZf0bGVyAVa4y6CrzZF59PzTF0vdlaKe43OM
CoEC8eh50E3nkmQXCWlwPTIsLo+CnNBRHjFE2JE+BFkUITydMFPrdJseIBgOv31xkvhcxMjaPEmh
d6iZFpgRcjwZF523ovQ2i/wYR6HCZvwYcHWfKa5QpScQzi52nnzE4BQcklbH8I9TLr+dCQFDtYmc
OO1+wRP6arF1rVCLUxekHbfypWSJGEWi9scsGh2kmHMjjBoUQDi4Oo7/i1gkOeNEx39lOT1GhOK4
M7oOIbXCux1cG0yEAb6Du6cNJ4qt2KCfyGAb5N9mHQrK8wy09c5bNvDNBeAqp3s5cqMCK3BLegXx
1zfWXo97ka0ZdPBaIT8XZ/d/TuewRnbSFeVo4pABdw9E8IvQ3zJu8cDjEvrTqeT1Nc06/RUOpTnH
pYJs2OxFjxsGH6jvmJyMDUKHthxlRwqa6avpWYFp2VcRqZs6FoizeVcgyHXMc23+ygKqMvzyPBrX
n+XQIKD35RlndfgjDtfEcewps0iJlfBQ2sxCHn6zSdibYt0gJ4fxMgg656VTeDYUMKGkY1e8GC/j
cnOP66/nE0PglsL+o5eVhb1PltkLG33XL4VyqFPFdSmzd839hSupQOrRoFVYBWWVvcjxe66r9CcT
+AWw+Gp6h3jyFAjt21m9LXGjRkqRbkf/UK4kA8kKVBU9OdSU+Dt/OxCibuxNixIyeDo6PcweX72e
kwDxpJNgXK8zITY8TT7SE97kpD0QAxJFvpoOe2f2aD2xHjqsKJLXvSGN2EcwwWQkSKduury8Y7Jj
ohw6CLzXU/An5G1Bmbeym7oxn6QyUcdz3ZnrNaC4uV8hvwdfismznSlyUmFHOHAlHXXvN9e3MqJH
4LfPCcwnwnVo3hgRQ6i9fuAZOoQvPlKL7LARQo/hu8AmHzB/FwcRf7sATeKKrHy2n3jRoQQmdLF/
8KZpEROkNL4dUG2KMsWWqVDm4YqThG2DHpA/V39Ar3G59sMc4U5IrUjEh4yGwGbVLRhWtL5t+arf
0wrUVC6wbW1F8JRH6pnXp5HkeleSuN/4PT+qQAjl9r87yXEOoFi5SBYASeHt0TSnpZ93uV5TgeXV
i2WcJs23+whuS3XGKGVvGWZ/ai8hhx9OfHztsK4AZxuE6HvJjzlACrRCljf/NwPGV7+rZOB/H937
9Jp4yM63XpL5dqczLAiaP3Ght8bTuM2Fdj9UC03Udj4vFhiEN35beJwbeaf4wwd3reFkvoexFs3o
ToBSqcWTEIGkSzqoe8dfzlMkzlTOHHnwwqDZnK6vtNGvPDcJSzgEYcn8GaTUXsCd9dxbnsmnLHqd
FUBq+a8ThMB0cj8HrP/BsjD9FZLDzawlri3+ITCwmCa6TEtLe5m6jyaHZAmgnW4uI8cBMR6+HjYO
iSWktjgbI7KJHvhiQOrPK2E8wFr5W3ZFMp4jlTlucxyTMcSQLbxZr/RROo61S429JDeDexIHkO31
RtoczfoQjXHhUQOc8dLF093GBdfZ/qBg+eJJXCkKtxTTX92imk0yHV8sEdD/bYy/GDhwZ/MFV+BE
/I/lUG/sltGPY2dEBBVYJgLGVfJllFmKzDxbyltuFriG1oa20P2CPe3OBDLqlhuYI5AAOmXHy2Rk
Dxccp98f17GCLamTJODmAxs7f8f+m01zmes6ZEx3byTV0vZLG/zX7xdFeODKVF6kLzKRxCvh1S5c
sTcoy5SQBsv4BkN296N8MA8Y7DcD5wDKzswSMqvUDna1nT1HNstxqOYHgmC8kdmOSAWo+ziFHVe5
TnG64LVrx/vYH/bIbIFG+5DYGSQ70PHCweAOF+SSMbIVgqRHnUThSQRfSJrUfjTXB73MTZZ1KeKU
uDnKRqKstH6P7X8Bj/oou2QTYU6FuSIHKQlAZeRRhdJK0i7YoYnWH6aiIsrWcVd2h+gjlDKL0DQf
+Ihb3tRdEU9lIfpP6hqAaxziQ6K1zC0pP79eG0MEBLujYxnN+jFkFvV4tQaIhCCpkrT3twILrs57
X8nVvzsj+LT2vJz74CqhumZBdbD07MdzjwLW7mXorSLzhEquAsqvF8/EEe8kt0el5olcoK+gV5jU
mQ4ZvcRe+V/fz5vFbbzTNHcpMVAq/2PF7ZqSOg9MzpX44DZ3sXkmC7ORv6eYCNLAXhEmki2SIoM6
HjL+AgT9VAESRCROPSINbc3knVWoCw/+HfT/e6npzJKA2XaS/7gVOaKYfPPd7g6LcgHE0vPG6S5U
5fyH6NSvK4f1yGSgL+yfPm+xnwAiAtgISr6DmXW5Ckwno11HD6oVuFmlP2V2GfBGTsF0RDVcEk6k
DbCa+NcSAUKokfh+g9uEZErPKRj2B6BaqbNwws5ddX7kjRp9SmICIjiwUMVnYOqNMlvvaWBDod6z
hBe/hms8O+JH5SzxExu0ooqmdtu0SowtelrZ6mZO15/jat3C5O+8CALfwhVK9qq4JPrGLcKj2DWb
rvLN/xc5RZ/zhIXkdRgGlbqsB5D1ZOko92tztq6O3g5PzLSPmM58FruH7xlHXf0D9gmDnnecIvul
4HM6OBfhmfkhX1LyPlAxjIrsRQ7+S86Oml0TrDOoKkOwgRanqrQuGEHFq9g8wCyhKqy931de3w3j
bzbbYd8w4wM8duMm5LMBXsTd7UZWebBU4eWQEeMVzNMFquExknIJt5qAsWxNmPlXvQpbl1sjKXTc
wvwRdotLlgTE33Z4iStp5dl8E+/8dRmGJRloXYxZa2yFy3ydv/xeaSeGn9jhLqbyVd3qH+B6LQqb
Kypn/ZYip4d07OIgESB3Z0nz+IKTcNraTEyYQiGjP1c0g088wuvn+7eIHU2/VH3py/spzmVAcHPq
Ay2aFTDgZ67YlIs7vdGLrlhGSdo4QPV9vbVsk9Pws1kym/0R1/6mFmvz19Io85ch0ihgra5Fk3Jr
KQMOUgvMn5YI70TriFnqmMidE2a4Lfv/Gye7VtuCcXbph6nVKIY116FDGUnGHIwAU+E8BbFsmv3K
Ck9YdJSMnsnrEhutoMaUqoMZlstW3CWsO2EKr1yflNdSnId1kDCC/DHY7KEdLcaxNIzNOigjXN4N
olgLFuiSDL8qjMmHKKiE5+0GoeOHnoDXF6vKk3EDxxJzVwB2kP7jyOyHoID2xNhrUcR1S/5q+yyr
d/R3k47RXgqnUuTll9nLbnGA1fTt8Z6zeddiJ/m2IHh0mxvz5Q/lrTD9M92vW7tag8bN4RxgpSht
vCty4sBJqwQ/T1an/Ticoa6ZQd6ukZlN9BTN1v9YkI3URykVDRRoGyK0LN5XmRj5M5U12ARQDDuF
uc0Ix+1wO9oz8GHsqLxMCWTq89M1TczFDV1r9PJFV8yWNq64MlB7k6waKa6AxsGxyvKaNO5O/J9S
9OxfTmHaDbChk/rqaIKJGEWzUGxK7XlN63ksZwE8q6CT8LVIPbl3K92qOgSCvFM39Z3qkRymPWsw
qig+k7malgyfWLXw+xGSyBFW4rMsSv+Y2NerclZldjTr8RSpLtP0aZLFuMB31yA8OsZu7d+I0wkn
rEBN8CuiIxTZyWbrY9ShdCU7w+u2twUadGyQA4GjpomabV1e/a79GIfFEc8Mv0tiHmTx5BP8kPEt
Yi/88rxOx3R4nOwiXGAZ9IqoW2V1irHCzrsHtrVRLSaqds3rcj3+ZJvbS5UJ/+Aepg5114k1V79D
IxLxq0saYkJYoZwx3slOSnTo7+lyvdB7j6o/wsXttK59Dl9Bmjd93q5uCRe22TbPUHDbO2BUYKcN
/860hN1QzICWu6yYQioQ9fM8TjtLgFaM33nDWsHED/zr7Aw7cyKiLr2NtJuNukw1QpAakdo0Z+KY
n8muTiXTH2LbAMkBeBlghKNU00ZitzQf1xSNZ9uKpKumvuUPUHi2bYKe92H2LaEooUNBYjJk7nJ9
Tps3FpeOB7BKn4os4Uk/D4bRvi94s+Ugv+mdlnYiUCmAyQpoS7q/cPs/y+49AU1LvQWP1k+RFK1O
FDaYMdCb8QvNixT0lJul3MP5WvLUZoveu2QMm3v/j3IVcv/x2s2oaqlo4kiF4yXWyHATGh9U9vxK
9QhuMSX54BEE5KEiSQpun1N6HbOy3uEHtWdg8YwQpf3rjv0fW9P2Ka1lQqiPddJG185GhNhHCwMY
iJur083Hvw1IJ40TCAD+sl2T/AR5XAgC4PSOIN9POKoqV9kLv4Q9uI+WRaa1bfGaAHxmlhzJChC+
mzu+MtfnbM+SwYrprVLFXiwhd/Y00m86ko/sZMXigopRRlM/WlhWmkmSHaKGvzwEt89yiUzDWy60
fXe1O3i7nE8dpcnzrDKs6aToSWxAPlnU9r7qHQ/8U+IfOf7NT6RN4mvc0gIxhSYPZ82VxihPyQgn
em/FnUZkpe8JT3rHRaMXYUwE8sglz6ruFL+7DbKa0aTmWR6XrHERmfcpbvmfbKfuxJ4gYk8OUofY
vu+wYHHi6EiKprPRszXp4S3ZNGDTm83eKPMbnnZA3OakXpSh7927sxNDkFlZhOV9SoCxZ/ttGxE9
4zBe3hmSn/MCP9Ww/+iSUskeOcrrAO4KVKrV8oUVR8j79EWrmR8T9Dq+0CfG57VF8gEnoFRj0Gqk
/49oVDWAudwQPj1DSRbDgNWZtVtbQIsF8yz1rUE5u/cHR6prcqcWQv5B6FPvIOp7B2UP3xEw81n1
xVTufrXvz1tNarPqwimLFEWOaH2Kq+NZ0G8Pj0TrIZQk72rx6ghpktFu3c8SqlvGKpeVKn69d4+p
/KbBMIvb72rkDLS8wgfGRpXlYuw2D0vEBqe7IHK4tAA7+eHaYm6yr93xh9XYTy0pVWHwIQSqhA2O
zRklYQGYJwVEP/oRzLI6R5ZcJoolnaLk1VeThKQTKwHLl6Aq1T27p+WkTADuFuYjcUEodxhQGZgK
0AHbLq/YtzGh4U4jq9wu5xxhDuaH46JA053V+uvYd1LZYomBIGWsHv02TbX+9BzLX+FMQfvQaKsj
g0oICDLF3Eu1yOLQPqr8Vbz5A4kV7OUGhf311YoZ6J0Z8oq96TqEIuZ39iXGyo9MCxAJ3DR0Jqze
+9u4/Cyi40qRSvueFCId+wKH8YU2S0zCo+t5xyVdlcBvr4Wlw2DvibSR1FFa0RW9shIImR6nCx2O
FrhwyA4EcHknHeK6GEQxFkxaDdV126Bw/IP4F9UQTj6e20luBYNQ0Wq7J8mYtxKE7RvkbTNn34ML
2Egla72Ibbu9HKzklE5LIcL3g/eji1gcF0ZyoQqXBccw/jQYjwDwrpzlE04Dmd3a0bDDcrNOE6Op
jFAssZQafIVHtyBRgyEqjmSELyC6ylDTREAEwPJ5RL+OkZXnRf1D5GXzdZ3t5vLyE3d2Wzzkty9k
5RP2XT8Fm0LauoOxqmLu58NoUtyYc1HjH0GnhVkwZ5BPnFJzMDPb5F3+D1LQvqEREGppqSIv27aY
Y6FpsHFIberOAv0OuQbI0XNU6jsY81ntNKkxRUQNcz0NSGsUcGJ6HHnlh0MqoItL1V9051iADPQG
Cb5Mh7+3bu+u0zisUwSzJp8on+U7pxBNNByAjQx8ywAka3bdJPdd/wYJRgdlL/WA979zWshKNfQj
SQfWE9MewnfiK4ucnfoztn8ghrvCIU2Crn6dUF4khfdXTT1Rcf+AVH4baVDew94FMy4ylJAxPcK+
R0ynNGVsjf276nloOlvH1ayFFfOk5t6PtEkYo5s6UXjWN9C4Lkpv/+NXH2tfLu9kEpB/Zsl2VNGp
mhM9dfAW1rH4RZPXZfcJa5LVSFMh6HzcfKy4q6DI1oCXp3sxtj8weLFGgoBIu04XPlJNYcEklhOL
k6/zl98zTK28KX55j0MWy7SS9d0bMSKUFnZnD2LARYRaNyYPlml9MYeZGodg7HgA761ym6kJnyIC
AfcijJYkbu7DouuZBOJQkneaRmJw/iy9WVjFG6qvDlA3RxUBMKXiWBuoH0/QqR+yLHOzSnbxAfCP
Ji8quGJOUQiE99Mte3rp6zokAvWlDnt1LpSgDan3P1VlKEmHbZ5UxxUIs4efvmHZnLgCi+lcLspO
ZWrw+OrEERyzfXGzNQMfM2j8jZZSttIlh4xtDeDF62DF+L2WfEmxaWYpsfDOFcgfmX7w1iXBx1Jr
/Mgr7uXbvbuAsj6jUdEcz0cZOA0Z3qK7rPf3zgtU7XsHmirCoubWKCrzaEKD5cXQrfeSQIRJUAXL
IPgiTnX06IGkifQQgFuMqgsDD/wRFu6eelOlCHLUD3qXTKDzPe26ASt7iKzjpKra9uBxza4rMSoM
ta3gadCMRqQ3ujNBAEJ8jAO6n99PVA9GZDUGQACk5pAUos1LJsmyvCuVdQhhOXVwwbpR1fuqTTWA
QLMXLhfxmjr1Vzxpv++BvmL5QHV4sI7A3FkMR9DsvKgWwnbMTdXRxrHOsaTgcZ2mhpt4AVTHSLIH
fWyh0ZVsTTCtb5QGYZXdGvI8yjbUzQsvkhIstJRa7hXFOmzqFcpxS8PWNLnjgGMZQod4jVKKpsyY
l3vW7TOqzy4iw7Z8RD87Ik98RggVMZkKuqyghlzrEN3EC6N9BQ/XvRRghYb1KxvD0Ex7X+aPESgg
gVIQbSaI1eNOjBOO68l1EAXfpvWjjg/1NKa7/u+FUmBqjPzw75Ce0/AIF6Ii8tXwSuxkNceqm7wX
eGnZ0Me2vmWEJLlkFsUi6BUL90Xs2fxSJg2s3kwWcAm8iFHMOcKg6aP9EtKzKGAlMseUYeqCupHx
C/8lqF4EuBiC9NQQSxBTRrRmqicyPJ/GcytR+han2omXMhmCdQcjEm1phCinwmRr+uRDJJ0WEQmW
i499jfK0EHyivwBSeiukjlD/BvVc3zf21YQfBTtVJhHCjlKAw4Ge/mBm5skqDPlA5cPGN0cC3Bus
9CLKwoIKMnIXjTEGlq57EbhVOpoNvO74GBQmJrYBcq5/aYhcy4jZ0Edvmcpo6PrDPeh/jB24i7+s
WoEkYNdVb6JEW4Do+e/NnaIIHtAe07L46j7Gkl56YnsuqRS16wpag9H/MMK8zVq3g5PAQeXvJPyb
sGhNFL9JUX5FG+ttBRrxs+oIgUT45gXVgfXhxZyUVcbNbgw905/fu0ug//KftWevssfIdNenNeKR
wmlN9zKoQAG9yyAHduqDLjDfP0dFpMSxsYFxMuwuLOH8gSqWDvfqZRk4S9J09YK1SuVw+F3hqc+w
nBWqtsQi+9MZ/5aMHMjTKjHcF6Sdo6X4Q24Gqko3pYey0RGF0DoBZabGOYeivUR0S13qNaXLGVNS
tHP4oQSX1s6V/C3O9WCy4m0Tr+cSCfVvyPjKRVDGT0KjTnER9fMZNsH7JmZ7c7QN2lHqTvSnR2el
zcDDH8xWrH5Sw1nXgqX4aP0o734lCOmJdRvG+9Drl3vDxSTAvPgoj8BAGfo/04wfFDFqVt9ezM8s
afuw84v1xkhMaMPHvmlX8X9pV+QU9puUmkZzHqGuci53+ENzXvonsa0vDNMeWqTVfbZCX5PwqnQF
0SelkexLMENyhLtrnpvFIFZkk1DAbElWErbk4Czl8zw63sK0R3QRHF3RpjLjOHZEUncjKzyVQfIN
aB/K3uHoZJwAE0wMFEYWpN2pHm4WDvc+ux8dH1mTg0lqnURlaupPYnjpYnQ3wu8axQrX6BNKLDa1
H1iEtAabt76kbbLvNrSzRA3pwLPGvcH178IOgnrCFmAFfxUbwbP00+3a1s0j/sh4E5lxQ0WASusN
mceWjiaxHxxwr2ylUk8zJjL7nVAc+4X6TNpc2uKdDba+QrerQahvdlfhajqZLnR/qtaeH6NIHLLn
H8H2T/wl7Ymsts4nrE5LmSl8g5yAYVR0w6Pf42/jkjPpg3K08Ou8WoGuFMcBf7cpRi47EDYu9zJ7
SpykPgLyFccsuL/Htcvr32nYORW4jI5dhT5Zl/9bzbbs2WluzhmcOHROzMCD/ByHfnkmm8KI/kp+
xneOppmVsiLBqeeeWSzx6ESS4DMW1SaMD51Mdtya6fLPqWoouIhb1dJEhk6kWM750JBPm46fA/Wm
OVqiO9m2oByCyxxzyeRTcc2fRX0MmPS8VHks0xPiKoB7Xj2GhgloN3K610INAHnmBEfAAkjFUfCX
rqBjctATp6zJ8SDc7X2Pv77xJZyTtW5bJ7ppSR8xqyitzrcfDzXS+uKT/51QOIYKwnF1bv4WZLtw
D6raEbvNEDxQz28XYX9aFtxR/m92LGblUUWUs/XCfMIY5lBJ0QKuN3Tr9JWB/1nd3lcB5d7GvSVN
k0ROXsmC+EcmsYOqF5ntxLWR7EgHaHHmn06YAQNasEswZGEPfvx4ph6IvKn3IWZNyuTQaftNrNC3
b2dEJ7Okc1DwcrrQW81KLGHWIpt9FziF9U99010L7zs4x9OSL5rw+BAbGiHa9bcKo83cUQhJ/6pa
8ACWB0rqevZHJx01zAzTsieIl6LFjLYvvxniPk0+iFD9/dEGVeP2J0uqK+6FTT0TigqqRLjBnQX7
HE6x5InHvxGm5Rkm7/hc5Q4Pl9TFwMFiF5/5XFSx3CpipKqPrA/Q1Bctp5z5yz0uF7QdZc1B4oon
E2aaKRUVm6OJndsb1XDrmY3sGJgIvHR1AsZQhV+MNQ9vyLfHKVqPVZUMtqyaLlz+Yl30O5OOrWsB
8FY4afpkLsp/7YluCcBimLeLEeSxq5oSw9nZ27tOBSktMrTMmYi4IQJjJepEokZZ3MJru5rS+l48
JBwcodWTBQn1JrqPkdYK8GMyt5qx9sAgxarUN3PBEi2KmI+rG4VIG5tXV17mgqPEAes6maSmbFYF
F5QXA1V0R9eOxHUXZ+6tJxD+s64gUD3uizT+FmDh2M8kToG5LTvV8TZqHfWf9kxTcgPelo505/6c
fNJsUmRl0RMWdLml9zngozlBfN6LexcTYY5baP8oSDw2VIGgctMiHDy1LDflVrxR0+Fv+mGYsQJ4
bPLL2fKBYE+XAIHEpg+QHJbLZyjsL2f0txyv9lFzsoX4gBH1pfngc2Dnu9f74xU+uJFcnnme+Lna
AWW3FlOKNmknPYwo9DSIrixkpoUt8ld+qncHyNdJ7/HgZ+NXpVVCvi26ChVdzKjspVdmLJuIGWSa
NZ/DGYBwu6ZIr46m57u0g1cR86BMpWOZpULeTNxI03C4NhyBOlnDjHMTxz9YHc4LnRp0SP+cKG7X
AalEkw7gcQR7DaN3dNYkOSss+goZEtTXSo35hqus/s7KPirL5Z6GoNvPJ8lqAFCJoJUnlPhtA/Dl
1OFWPypK7LTNIs7cSVTlO09RCujhua9+JIbg+6uEh89vuody8VQHjnXblKNZbXonY9pn/tnWnYmC
KSvjQ9Q6BIwlp0BWVMQKEvEieeuROnGIYnIf0KYVLjmYwanyBViyaBk3kTFun+PCeWn4rUxc7VgG
80A06SFoJJFBO7hGFIvqYPsP6JpX+0W3UJKfgC5LX/m2bYt+LrrBIJmrDUQ3Cu28uFbjwgSztgsU
JZZwCLE/RoUpBv8toAyaG1jQKqjwchwm5E6uA7yyJ58xZLgs9lysInihl/WUDrFLH03n9jStpYBQ
Tohv9KXY48IaJw4ktrEFdLwIqfHEqmWpovBSoIEliF6OdsKkiZdf2sv6t4e8MBjGryfAGlWe4iHk
z+MMaUxcyJNNDQQ4zx7Wedq/SN1tLYayeahVDUcyA+y0kmrXFjtYDuj5FhF/uDmtKZvckA8OmI1k
VIq9vh7Wc4Dz7UQixUfVvZKKKjkjyGhAv5irIfYT4nACZnF7tyOXoFlTuHulYQ5NQJ+QKhcOGX9p
mRSE0bNsSAO2CU0KSoIL9PnMbo9/Iw3q5Rdxav7jZeNnSAAeEqNvBhpcaoJz4qF9OWk1eDhdl5rG
zRHSMfHCMTSaCav5ID4dXhvl3KNUKBKENgkTVKnbY6TCjDSumF/b7bB8SukAb/0K//CDiiw3NszQ
95XJDAF4+gOcm+WlA5qoWwx85ePqgoS3IGD6sXWL7By7drOU4Ly0eXS1f+6FbmXvu6FTvmo435Dx
/tI+bGN1JntFIc3PslrAD2K4PblWlpxdzS0Egh3VGsHjxMnPA1jT8VsxCjjSArQfSh8yXjCB5sru
U4zeEf7hMysFFCiU/Tw2DruNlIHCDpPny78f7oy4AC9WZ8Tli8ukMv9NDauawvVJhjPHIepg8tPz
lOYzJXgzoILKVVeKKqVHysKqpdqG8kOBfjwb4QMue0NF5moImAKmwoc9K40aFETe3dSpdEPPKbHg
iy7TCxSz9dmDYPMfFmdM6osnJbhnys3TsfUkKbKgwj5lspGE6DCFzt2ukJM5OoiEuaTkDMegQdMg
b9cMFz8slMJ09aZPUKL3apGg2Lb2V2dHC95QkzrHgEY+PgH0qxxWGIqOhNpLfkufuddjukeBCkqA
aYT1tTv4QKlaCDxO83O2kj5QGbt75Q+rYlTcjCcYF3gHC5ci2aoxmgYgvlEXhnYIgMHdYgHdMf7d
Hb3hbH7RFYL85byhkb0OSEGxpQnHXXboUEo+Yol5hLZxRGp3UG4p3Ib0MaadPMAFLBD1h+OJQ5hE
SXdsNvSxO+ag0Fa+KPH3fW3jFag3p/sX8N2kUwnvO1ETH/CSjT9LDrB/dzkUqsuJkj8m+qrdOF0y
BVN7EYkQkM4cVPkxpvl2xHnRup1Lnvrhmmfi8q8JwAG4SeZVe6Bbx7D7gkX6EOkHxVi6gJ0NMTVo
a6+9/IYfi9ka+33DbQywkKJ1dVFLbY78OHDXRJkoagf2g4BVilb+CbiI+GNM6VgmOPywJEgDYHS2
XCZBuL1GRhTcfi0GW6DY/Zx7rHBnJEnjrawicwZ50TGkZIR06iyr868DIb1iu3tAdO453rGukfc1
w/n65SBN5zZqs5kpWGXek8hgHk5j8UiXGdFM8e7z3lKb+8RQR2M0gbolq+0mr60DL2lkGjhEnbBC
4+ped3f4nz7QMcgMLZR46JoRNJnWDZAlTgtYB278wBoYyGkx7foV6d3wAPb/m7G7He4PbDOyNUi4
AL4pUSz8xTy1P8c8PxRnLE5MACLbrqRbp7QsQccy36NlcEuCS8ae3g6ZRv7WMcKVPfRviSRXMSsQ
wacCIw8o+6hhYw4ultepfBFbrM0QwkGFWGqZAmXurDJpRZKyeTnK29VgXk+NMlX6f4LvsurLJa4P
HFTcAMYPRAxBr0+saVa9Juxm1H5bQKW+WsSbrBqrIxTC3C8suo9FfL50PtMGryhJCnpe2RbwHwjz
qnifUGudgCIMa2C/SUuSbcgyhBR3DAHCym6yWYFSvisyeF+z3s7sd8q4bXsBCHDb/Mh6fHPLTVj9
B8PJWTnoqUHIhIGscchfEUXORXzwcnvKQ28Xf8yKnHWzWfsYJMfaKcHD4JJ4YNmgVffaGL3cxjzt
FzpUsuLkgtaC98r5RiZ+S61T3mYXNslKDuV9sGX9pCDpS2+t7Vp0P9sJ2QKzQVcfVQrFLi7PK+OV
f3bekfJRPiRmQWDCRXX0RV0r6RXh2oIgiiT9BpzC/hp/suaZXIArH/nhTZmMFZRQnpbUFdGtnpWj
Se1T48TqZzjyMCJa7F4iMUUo3jagVD/dbbWoc+rBFUbuCuFyiBBvfX7M2R0Tea2B+75lIWG99UZs
FkGLB/DlVu8iLRkZj7RtRHkAqaywkRMnSaWejoIxewqro073CeIFbKmCOgbF6ffkgsHUTVMVPcbM
Asu5bkyxWagDXosAv0amcCsET8kGN+9PI+0xchpbCkHD0dLldwTgDL26crEy45zHoitUB/fqlgeH
8LDP52rzpbUnKfzF4MtMDCDKshwrewJpb7TfxJxr35MljWg8Wt+ZvJT5XmPzDsfTwktsbxNqZimw
SlaI0dCdp56/WFEMI/wnRtSID14xw9j1MU+xtiCG4aKkWaN2AHokLYX6tnGdcN6gYakYi/3dY0KA
IEGarGY/JFq5U3MUou20fY6ErjWr8/VYcyWWBYzfdYgYiOo7SgPzX1iWci2A4it0TvXruKFoTeTh
jKr9yiyNwLEnGLyLAdRKqhKuayhjWGvkS+sUe2BW8zRVUNdg8tZt/JcbneRAbmoocnHTFfff5ICM
nsg5nDKvCNBUAJ4IVMCVFCUrwZ3LvE+G2atSXs39CIXqGfZkiaw4Ixnd4H2TYXreR4FgGz9sSuBJ
M7ZZJnB2BeXUVb8NLFdGh/26r5pW7BnDTVU8D+O1CejcsxZw7S3blaXslgrKa/RsZh3NSH5YoLIe
S4Y/j1IBBTzbLfbdmgxQ0RymUZlEQvnFxf5+ZchgTwT3Cnz2F4+81iFjdZoxglK0u0N8PZdrrlOy
MUVtdPPda1Trc5TOn8QH88L3akjqnw+YblodTWqUEUJ+j731mjFs4WmSTuoDs1wsw4ipu8PdBAPi
ZhgxWfU0DKYIODePKFH40YJlUBubBwSsXYucbs5Q9ugryyt+68+aEgp+l+q2UqmdHsujDsOKb1zA
swIC/+mrjPyLlxg//sqs/hMIlHwnaeT2ss/Pyrgnlg0KORvq21s3ifv7zp8QGuX+wvIwk4EtkwZ5
Gc0u9214YRggT7IlIPW5rJZe10yGmrOLsSPw9xl1sOINX4Qz1tBLwn8/M5jDht+w4NxW2zGQ3Fej
gSyBSbckAv6LxMHc/y14m1dO+MEFywjiU2eQfyMlquKEtG0XPnePI5c/wjxjAKBPxeX5YEorf3Zd
T95mWVk5kM8wWgrXb6ui7393kB9S7ebb0IphOAi8+aM3cX+kLBmpZ1voy1478A2naUZH/2Y8PYyB
AxUnumdxBoGWpgHxA2UFzygCZrsoolaIUNkLslyClkcYGvzxnVn3bad6TmLb77kFV63MeQPyvLl3
1mOLK1A0gwF3ofkQRvQZ0cuoyp5Koy0Og0k+yaO40pfJA3JZ2di9ImXSbJbP17mNMxQnbQY/cmMd
oR2ywAmlMpB5++VpFbzS49iG9k6Etmp5imELKjvf/GX8/CeXySalke9P1rG9PMp5YgHkElh3KGtr
fbXZw8rNeMHfDmKauf9zT5zvqa+Hz5VJmn/TeoUODDjeLlrtOQuTBNm7H2MsSCD8CXj3IjHqZRCm
NBe7VTmYhs1uzW70BGYJfIGqCxK7rPtN40wqxjPF76eUZRPyLRaBVhmuoyRha4pGKGkfJrlQfyyh
hYUwxBc1kjGbjAutg9S1prB9KNpXeftIA62xyCzzS8lX92judxVwPNVcDtGJdzTh1nvpZoPivRAw
ReIt4ZFL05ATiAsiOh/2xwqEx1L1X7DIDokLL+QgVxMD3PVzl4Pc3mO54ovaZ4A63E37cAqYFj09
jXqeeL1cFKTny8z4OEzzy2xtmgucDt6ECmeymooDXPAWBAGnqwZfxJEIqqP4GMoXJmEeBvlQAs4F
yQY9oELAUhotUQt6WmfMJQBTB3+5HKcqlSNlUgsRmcvFNBYMxgqUgNZCQI070/oEATQHc0Ucz09K
xr+nmY1YzEQKkb7irQcxgAU/zpxUKztYGE7mfwwNuT2QOYn/24pjs+V5F/SNDqrpIb9JdIuU17BB
NQ19tQhH85I2EEYS6Mzr54XAiAwj1AlfbtFYGmvCugOAOZkZAmlKczt9RpBgu/Ar7Y9V7dpNVMwg
gzG4Hu8LWBhY8k5yewTXJBheKft0O1kvu7zwiAvwM9GLb6K+wLza9Dpx5eQeYhPsMYHEQI867lUh
aEY1dq8gffpe2U9jT2hN3fT5ofkAFv/u1dPSc1pVgaU77zoP7u59Q7zCh3Z+psmsCd91OnQgS5Da
/2mI1cdiMlY833nmefu+UU2F8dVNQJwjN+8egAiUN/MwBkYlbArnInJLdpuy1fvMG9tU+5fQfpA4
PFDzBhvOmVqIzMO5OjkmCGLlHlYVhPFnVznrJ1VnlLai0vwPRC41P+cEKz6ZAEAmxrUAhuiqlVmp
A/eEtCBiQHSG6ECezqDiSbUKyEuEbR0wJdw0SQBNbuMqJ3GtgvzYr5AdrUAC7GstpFlkPHmCz/rx
ANVKQ0xvV9tFr/8Wf3OGBFHBys1Ob+Oor9vqPwVbdHyZrfe5rTl/oNrDbCb4qPjTncyoph7mKVup
+3TYqjHMp6+ex5HkHRFKqTeLOjb5upY0cbgcxk/rN2N5HpFP7vW4idD0DTu8K+f1qPzTnpiRmnuv
Lr0tBxLrXgbubbac6vG6NCCqfQZ+gHLnVXl+1pgHB5ccX8w5Lqeim8CqKmzGT/jWVxSvkcKT3h8H
M5XVFgJT2qZwO2GeFDDOIdGsQasLwVvq1pRRXxxwOAVJGVVxVS8wgb0zK6h2idRzUCUpOzef6Yr7
RWClfuWJqQnCgKxFf4FYfyTTIM3WKS6/I/gieYwIF8yDdonoDycJqfZ1vDP9v4a/nPLbQYPQ6Qdg
vp9ZEqhs2uTJxjRVcNu4W5VvgxaUfBFZ7/2TFu01es5pQ8txoXVtect+ghFuZSKMr8RlLoSt+CSM
EteVKJ/OhUepE3jrm+5oo/lkG155IL6bBwEW/QAG2KqQ8T+CIa11zSINprZe1Ilp91DJRWYHgQKg
c8Vo+N+eCy66A79NM7wCsCLPHbKAPKihLB3XHNv6dsqxVI2JuXi8vkzlfoQjwN0VfcBGYfZIpfNY
Kj5UZaheIXAV0IWWaEQNErbyViL+HujaioJZQSDbHpafit3YcylhZmaoBFCR8j1L8U0qPwh15DJZ
akaYJdIEzSeDf9HPBcpecFqG70inrbdlEAzikgfdcj0ipSxbJug2flqFhMrhml8wqF4f28AlIHjp
SL+fK5TcXq2QwOvy5Jw1sg8/JVWI8U/RQDSR0dmKWdF34xkb8IEkJkXx8LKToxRITgRpgl3tS5m1
GfIiO37gzmYjMsq0uz7OeTCGWauctC8M8HS1/++jZGiyE6GB5igQXSUsvfwHQeMerdEVpC6++Y0I
3OcbXSjvHclF/gT2Vl8CLLpWhPOz5EzIj34oq5MlmP1RDHDT6PFo8ioDlRkcaM9nspj5m4MlKDph
oGYQsblzODnNj/LMHN1L27sv5dXT796axvUtALsOYh+48Z4qcFhYswC8eYUr8D6hPiPqP5azMRU0
P9FZgIfr2cDCKwHX3TRFfcrabCKp8EArEVYBdcVR6djKv+7v8oijRq8VfjtQBdq0Bf1F1xQIKeZS
1JdzkKxfgsE1BWujw05o5W4fA05zhZgGpRjZH1+E2WLU2WgEwTmjWfoLqgU2OVD2XoFP4xM8u8u1
IeiZgA5zywZvEIBZ83oclQRBSZ+zLPIdwh4SRh0wdRkyVMUoVMDbg3IS5Tkjo+VOVfg7nRjllbdT
zRU1bAqngl7RP7KuOCH9NA65KorMjSGvkaGz/3U9fFmrhpIKLKc/2EhktLuLtUgqmKo3sXqdW3gC
wXoB+N4X3OzrHNGsbO7hJzAcPY8FzAHS1b+dz3Uaqeh7mfvtdjdvyEGgUzsN4vPQjpBZ/btI+A3E
LY8aG+anHdx4MHTWoRbfX7JVDw1aThqMMZ7on6KKdhogJkF/KxHpZRJWrGFaC9xUXoYjZH1hkUay
CfJ9UyI28yiu/a0KE+MHM0wtShb/sPxRjnNa0Hf6XjUAZEE9uzwIiSHXolZXcqyRLS31bM1JNT2+
J399lHBrEiJNkpPJQZaMpdTRFSzNdGaXHzwTaJVzkHM8OOhP6ps7GFGK/CpfO4NwNY14FxUSpJz0
fOhdFsXtv+7ne7pyOpIKdOZk9TaRPtxrnCwcOBSqy3a2GgKqXJlJYu7k/1USxp6C30ZADAtiRDYM
urqxy3zb8bu+VhXMR52tAV8QzXFiZF4mFCKSZc/a9iMShZwSucNTMO3t1V9hJqGH3+pYgyIDjVSI
+CyhTIz0AZQJdM9+AlUcgmmktDZlAzETR/CkS8BXTmW3GViX3KwTep6SIShJeRci2xWyDMxeqRgH
i6mukImdDxaaqiL/tVwUFXv9k7SbSeNBdy5C7TfqkDBFoVWStYLYpHNRcwrIjVIX6Dn24WmFTeXK
yBc191MIstkpVwz86sDZSbLFkJVhR49wmpLrEPml06Q0yE7RSubskfDLbteH5CUexCxuuKfwZEr4
TD2Tba8jG6XGr/cFzHGA2QwADQmfbOsaaXHlKfJgWnf0fRvIDyZlxRBjfgLcXkpszfiUUcJCij00
2ODC6TyGgb9X3gbwxW4x5GL0XaExw+0Fxj7GC6V9RU5jHYmx1HkCgZHAU5Pp8Ma7m5c1HnDke3LW
y5EbQY73hfVhC89KcnlOGKoTo0nMAsbSJlUeU/oaC8rmIC1PZieHXo5wtCl+GyjCl34TLcZLIv0A
9z4fGvwpmBWlbq+IjeijC/nfeRljWtMqnrEiFO/p0mW8KkMK21jkyCvvv9WoPyWgaX4WyXJdw4Vu
AXsIsR0MfW81j0FM6rbFehNsduSFJP/7cchsQXVcNnKfdBZ2dewyRJ7pCHoVp/O5Wg4kD8ZFWhT8
BOQtcZRkiYkxnSKlwVL66iz9KJVE+jmzFb+m3BZ8+Qh++s3Jj1wvp0jdZS8sbRVk3Az4iY/30uZb
uaV/LPQvo7trmfLZlP5V3HB+FvrBMXffu6GlZ7WT1Ri91zRnFX2gLVZSzibEc/IsBykVcG3mB133
QRFde0sOcAs79XpofCYtchkg64fUV8f8tf/cKPTHPNNiAs6JD9BSVLo6Pi6O6gKevrh9u/M6C2+c
gfIrHob3rjO3EuTl70a/ghN5hY94O2mLZHfqD1jXAitELXuW6Zv6uD+156eH0ZvxMYY2guQ7Pc3s
UY+S04YKna5yAqCY1clHSnw+VSlVOSN4Gyf2HMMR381Ubfy00WAZon4Af7MkM3Ja2bw/YdYfPf3A
tAjXQTL6uRpdq8S2/6fMkynXRwF3aAgCSU2BUDLSmHNBWs7i1VnaonigAohUVcquC85H6VKjjn44
5ylmq/GWv0Wcp0jQXzMao8cQICqPKxC3G+uguDKLjLgJMjzoEnnImz8BtjntDbGCkbSU+6jWYcT6
mFvMoloPX5AV880P2ymbKnP8++B5FZzm2d0wM5anuQqFv94mbA1mfzHNfGBjOtrOPWC9d62F+pD3
hx8QBi56+ducwJclGzvB6VrgimF2j6dbZvgaTv+2Gdue9gU0ULbUhxM1rXfIiDT1GDDhXCggmffs
jzM1YsTd+GXSoLyhMWa7egd8soThp3Uipqe2wKZpXPJFP2qVgjWTF5nIBHu69cd/NZugQY2vryTk
qLw8ZBFAyVwdcAKwxeOkf37sFkALAB+gj5RteWPscaoK+nNfqoWVzlfNwu/QvyiavVHRqRldXS0M
hJSefnCtMW3SqSU4l43LLGpSQ1i4HwJpGahKXEOt+ab2zzrHLVB19EdwWvOA2NBVLwx5OAgZG8l4
ZVNUyB2JLT/EFGyuJQLCeoFqh7CXOnBKf3TLiyj0pwbaYjW+ARah4mnDX/TCnHBmNeraPqC+n9iT
v+LdCOsvv6Yr5OCQmrS51OhemdGWxo1PFvdmvM+DaasZt9ZJ9lKagVbAgg7fX4cWwyGOLnGzqtkt
By4pSI7sMHLCRrjc79X0nr/byl7VcYpPZoqivMgGpk0JLRBpm7yYId4BmnrrR65xwJknLFxVjPAX
anJrZJ/8Gu714z7ViftSUOV1olWmHrrT3EFTR+Zga5kjCnd0HJKGhoAlD5GoSBkareuTqrd/Me9P
m3IRMFpRgdrQMhg772OHHJ1M916jjlyod+6B41a6wqZ3PJ/2N9LzBdT3Xkp8AZw5RccGSptlE2v/
WHwOeMwdvVclFR3NcijFyaVfGNcYJ4vKNc33Bs4UKJ/AQZrMZQ6aeGZJ2yOeUmYeCAUruBdGj3OB
LAAG6DnluaSpc7kWie0QClkfUClLWPkrnc4vWbCqLQusRtbpADeV7gFBQ/3Axr+N8H5RCVVI238d
2dKlNfZiDUibc9FtuVL6k/8EdQskiMPpuQ7wS+fnoCN9nsqeRuZBoXAKZ4sgjWup51I5IhCLvlR1
WpLCL4BFtwzFTjHAR3Jz5q76V8e20WlkMxKUTasKAaxAI5R+J/Ka2qZJ2+RtI0UkruS+DKdyUvO9
+/S00WUsV/xZnUmB/w0MZ1PIrSePlmB8M659p36bdHPFQz33pvVRy+ySqBMxHePeh3gNDhgv7FnT
dghIYmf4N5tO5L5IYVyrvml8O1DgYXGJLy5pi4N80ZbzJ1uCLpNrDcTS0UMftu6DRCHC7vsH0DEV
devEFYdz/JU7z/ncdk3Wko5BlEoYb3I7zn3dXLBE3h1t9LqEW4xPbZYMvucZqjvyjgaxrzWaWy1r
zH5vRwK8G6Sm2+xT+iSeAOCAM6DuFdRZgBmDAt2q1c8OozieGZihSnXvVjFL0JA/Ya019OKT+2yL
fSwBM1TV1cMcJONxx8onQL4sRSY5jqHVPCxtGFRr2Pq4rk9vHzOdKdjn3S4F5dQ/133x4evskbx3
xOL8/P4jsQWbhto5kc7ioV1wI7fqmj5no9ZgqJpoJvMG8StL3sAu3foIi6Iy043ml9XZvnf77wSI
M0MhF0aylbd5RHVbSjjsFZ3YDmKh5YC7V84vKsGJGW7zUd6M2RJHxvYRXAall5AmBtBYAARsDDAc
TE0FC2cjk6xb0XTBnVF0/98NCIYTQuYn827bEKKRGX9+cUhWAHDhsgnSIpgVzfvHob1Umx5D8Yp3
AINcmel2qeDeqUzRmkItX+nxbWZ6v6Rhkmwl1T/s+4Q61LIw6aUpUNp658pByR+I7G3KfIO9VCUm
gJwBcDXtpAgtPyiyaLsMu0Ip4+uOH3prfJmxazL73X20GU3egbcehKIvwYnYQCn0JyGc9bvykRng
lh293LB2z8S0kJxo/32pQl8dzkIg4m5gG8TvOrmVsBYCwrYERtlexkSbgetDIs6+eG5LwvqcZrMT
YCie9sQE5bK1xzEouONf3HdSOtQpK1x9qHme5zpcoxSYxM/RLTN5FOcwGd/woovBEiWyx1KfwVrq
1wq4OM96GBvagXFc9rQk/MwXyNv/NH9bpsg9EVe0ORW4tUbR8nasZwcBS0K6wpWFNtZyMapZ/xiY
2fvLdvGgJSP2RpIa6QYTToGC7Y5H4u6zOUOHgOmhgEkVRY8U0/P2wDMbdBfaHKh3vYoZbB7zD6kK
8wd/hxwyZysKouVLiFMBoO0jzcYST4Qyszlw9mIoz3QCtkyHe7KhEJwlW8t/fCD0HJz7VHR152GV
zjAGaZ3nBtWVZFGtvCZlyQ56aJxS5RyVevywOFmm/iYjnr018DyoL0d5SoFZFIiYFxS2woO2+tPL
sx4qoG5a+m+ctJkIemWvsBWhdaqd4DlPq+qpG/VGmEcXQFPYVUokcAMDGXgevGpDtBEEeaYCm8j+
pUFQAm267Z2Pj6bJ+HTGxKDQayfZzIyhc7SLc+Rj3TO2um2+8Y7wjoV+Vu/FVdl5quopcQbifbb2
Ok92bV0UrZ64qvPFmqKbkfTsnUtod4ePeWagDeZzBCBcZBHPz4Btf7A0C/RwiwxCib/Dk66f0FCj
G5dDjHJ9p33SGCMyZwCBx19kCJ7OgaW3O5Yf+kJyRDdSwSBZLwap+NynRzS6jns26DQ5ZYYjbqnF
PkpRGxFDxq9D6cu/lo7J7UIgpH2O9TpHiUKRfhd8DCsaxRiWwk5uUeJoIRPYnbsTB5Ih0mJckV+h
cx7LmXbCLaZ3X0MltvsTf/hys9DTeECk3IRCIUdBxqR7dPih6GdNU8kianejAO97/ZjNBOtBPRjd
b6O8J9v/Jzj1tPakB89tBClpEtgT7hHxvf70GSaQTJRCNzcfsCGwD7qcSde4Hr5bCec5POppPsG0
P6B8xeL91o1YRA9FioT3Xn1CWVpK4GO8lWTPZK16UyakVgonN/fWUeJbLg5FnuMKb/ZDS2PVGcSK
VqGOryMcsDwW4XcLpBy3JOQXTviNIoSbz70xXjYSwem5MBU87zOCwDllpdAR+ilbicwzAc8Np0gF
Jqg6MiSWv7v/9c9UCeaZiGKStPwciKjcbiLlzeU6EM8ATVfJym1S9V2orY72LkufOsaH3NUioLOi
+7rjSb0okBivHwjSWtzo+IlR86LcQ9xsZt+svgT8p6mT9TXIk5CCP/vVvsAb1oGrjKaYCMktQ30p
x3qvSMxkYQcnAkqhD98vUHZz/q+apLqU+L4n4+QswgWxPyIa5XT1W7UkY8VCJMc1n8b5s8egK3tA
+ndIzVUyXVNhXv2iDzt7uc/kS20t7NY0v+Bv0w03IKbz5sx6oqis8wu1sSoPP+Uk5+u9WTurDL9r
JbGWfxrwaHD2c7GDBj4JScpMoxxmkoy9AaY9dAiPfoUwlKNrVMWgVlu6r05nNWeqbpTFNNPk+eMU
E/J4xfaco/2GD0c4lpa+kj6twwqagSZcce1MDGV0Q9u3enyBtcHNlJf/fZZQTPYrJx8jx8wX9dv0
1rtTQVxuGS5f6eVeBnsueVNzCD7ei7vnF5ZmWOR9m5pZ6mlgnVnIr7dpIHnGJzf9np/dVSVpMHMG
2IHlaIMgAMdeZ0zQ8et2PJI/az7jILK1NrZIl/oKwJZ72/CvPhl8JsAvfvvdwtFllvVoKOYf2tHI
F+Fb6Zx/Jg7e24sdJU3gE4NemT+XCzBzpmCmR3C7MFFKDOYdPlyaU4HIukT4l9HQ/I6Ax+0KpgHx
mOFDJ+kW+Hm4+vuvgeZDtqkKa0p3+a+RoSz3cem2pYlrU69SkPcjQQu1lrCRDC/2pthMoQ660paD
7r9j4saibuFdTPS9D5qUwiZ1ouETnQWAPvb7Qio2SABextiCr3X6u8UqXgNHi5ZG8p1XAOfnNTBW
2DbihbP4vJlTIi3nBMVJdXl8e26Nw3n4D7SqwL0P0zQUodJCRB/UjkZ5ppfNCRAPyZqzd2C3BmbV
xCkNOxhHV8WK4d3muBAByT3tHXXsJTo1qGddud596OMtZDOFooIWovCexgb7JOmFmK7RnlveUiY2
UI/wkC6aWSlOYg1nOkkpHXysQWBrCWiFqQ5Pin3IoQK7nz2clUVluuBJFVNHtiRhrGAL7SlWYtV2
fidzpJ0x7ciiM7ZCA1YwHegAj0s8JZnJvs2IHXtdgFKovYd+0OfgrdKfFvpIazo66RoGtZkAYtP5
5zygthoFCpvnqBa5GWKtu+fAHn0rqSZrd0mD/O4g0DtoywRf9XOnxCm4xFXQGdH9o69VrmHZcg68
TKOYaKOoWZiDY8rDNpeHV6UgWkBuZnUyWhyy+QzdxNMtIwwQrzsTAW/VTsp0ykoKL1zOap/1aEuo
H2Pls2ENJJ+2dIZIqJa2ocXtji4tUMRB3UMP0jAV3t3SWUJ6T3RRsgPq102zjrEHVrAdSTptFa4y
OZNi+hZ1mTV+tRKb0vozqoLkEfZhRHYQDdwV3vSuu7aaawATEwyKcE4WBfjtNMMuN2MQNi03MvTx
5cCvlubMrpf2ULkf32eVLSvkY27s1zUm38JENFMb/iPgygj2C9yksfCZjl6+bgP2NZSXaYf0Xhty
/ORDz4k0zbJ3rsSCjgllEliWeOtyEosjSIAOYYTpk1BDm19ebRwz8mAWmxM1WfRiETOa8nHaSRQP
SM/mLcUKxG5agZYGlpmdtyyqtncwNL9TT0uoABsQgj4OVXtNdDp78YXVrmShhNH9/ZchA9ERL1ps
07ue6qdrEbP5YoHDZRdQDO8Pgn66RkAMEyADZ1d4XuqKOLDTkKct9M3/zGkrPUhfQQPaj0AgYi+j
ryd5BE2fAXTQ7RGOKZ8XSMgGujvQWMPNOvnvQ5FuhCIbgb1KCo1uPy50CAWIxnp7FMWwEFAx5Flx
jV1rMAmhC3QAG/Er0G+07l1DiTJ86IgqVu2y3QwicUR5bhgJxbhRJSvlK/IRlE/GOSTXxZvf6BBv
eEI8uHuDHQyjSs2/fVyX+FctDb7wJD4WtsTHldDgCo+af5q8xOVrPx1t0Go0es58PSKJ7+4NDmSD
EV6tK9+ATq7fy6AALuGpuxMcXt/6UIoV+/0CBhI2kYYR8vKwwAKCpSkroJW7s8/zfKoyCsM31Ws+
AZtr9UX1ixTa6LWG/hC6nsmWo64HzquRSMQiK5P7kkhcHIlyOXUM915bc8W6jDYda7twaqxyIYGw
tCXKTRcNUkyPHadJ13HP82ZJ9YM3K/RyLPYVQ7OiDDvccouBZrvlcvvflRdLJdhv1aNnXGhjcuLV
gzoOecwhe7ftanWnYKPQQFIj9WBfDPTKd7OUCim0sxbsgrp9jwvZjyowuovmXCqtH+C2uTSQzCR8
cocWmGuc0K9I4n8tTLRdpuErf6m/phFrcWDW0FtuKfNnvwjQwe0qPdVwaYHy/IsrG0KSIXZMFgcS
xvdHPInkbW9NnhE6qcl3cKYiiqy9Ce2AOK4hQZX0yCof2r3JnHnLjir5IGFNr43K/lgc5bPm2RBW
qETLv9I3yB40g1iAHd25joy6vej3Hzwn94RgFuKH1QaZibtRmCdbmB1aJyeSRLsim/PfZLrJf0C0
PG3M6MFZZ+zlfmo2H8brU2ihl9RKi5pRvS+s1+Y4Lnpx+d4PdbgWAJtxO1YM4zceV5bW8fh9cyug
bs+G7UxT59ll6PecWDLKuMovjJKySwFv8c2C3QU6xb3uzHJNnNNV5XPYs/gn858Lf9vsnPkJ2sVV
LekSyeUrr7Zd10V5G5/BgshnCDM2cmMdYtYsSWMTlW2tw/+yeZ3vcXlLd7J5rr034MotLiEumo5D
A/LIGhTFBHF1G63V6YQc7IYp06iVCOTKvQDIYBafzoa60ZVD2ahB8PDZ2ZKhvZa0Qtn0OlPKn6Px
ocbBW9cCjMwqwa18Ufo0vNZU7TPHW7kveCsTKb5xPsnE8rp5QalRxuswma6tQNpFXHSlxNyLclIb
EtBwaFaARh+5yHfdTsZ/KPKcA3Y6q+uDjvbN6DgKGbJ8TEzKSZJ1Ha0lNHma11cR7OuuNBa/ZTJz
eNdwA3fIKyj2+yEj+oVhIsEzCzATSays1cqswWAC0KxEnAltyMneh69rNYaQY5ZbuMN8mznCeT/E
KWaH8E2BpNMLVAGREiAMsYrP4heYYv1/1XBlAoZkJFLVHMdOM8CwDZsn3WnG56Zr2dUV0z53WyRZ
R63G/3Za6ly68n41s8KabY4pGobt9H6rNCSOgG05aHeaPhjDTjDBwVjNNi8CErMoAWfxpCbIWpQs
9bEx7TDsHyCZhLM8ZEudQRyiTBKcEO3mLhx/F4z6IhRDHdzMSSwIQar06vWVv158kenQuE25HjJW
aoxmGvNbPscAr+/1kW8DxPQ3zXcbzTNDYrtnguVLZ1AxycnfjYglSyeAzHEXcTbgz2NtGkJ/4lTu
UlKlDkio1JvYpDvvRCDgaRKjq98i38EqYg2ehDT+wKgKoFZnOzbpr5P0F2DD10n+EmwUNmE+PWqb
AQpn7mEKIm1XZEVAy07E7njD27V8rTiUq/1Vq3SfjddWRLmzyoFOprfiXmMqO128rsO2TRmeruNV
DcUM7tGeNGoN9ZDpGi/jZ9YljPDQYHDVYFLVz3J/e3GOh909DfHb96YupQ0rt7zhFU4nmxTV/3h2
94oL/5ks/VpXw4S04i4BOkJmM0l8zo2vEH2eYADW7FdZRsbdprIDsxj1CCfL4dBFTt6vCsVGnli2
lLYm1+9XNe0iO2MRPEi88EeOwVpthwczPOQLHYsD4qLnlvhckAZOV3rs6rbLicWXDPucOO4qsF9L
O0koQUtpWUECQ6heM1KOlpSh8wQCaeVSEonPWs0AKMA5Ytt4eUKDEOp6kIaMwahjuGpTlrgPFwbZ
c5VqFPlvNmH1LPfvzEeRSzSov852PPtpEsGxM6p+hq9BtZNrcCV59aGc8NBsZRjSVxNkEAVJf003
nd+reAW9E5Wpz5EfGHpjEf7qrheXm/7IiuLzxQQHY8hh3UtO5iuPVzeXakqx0O+CYd8/nG2X7j+5
EuWPrJlY6MLtIsH7GBO93WuTCYWxip+UkDeakuevsXek4qVop11yHUNLwCBlBuCS4cdcbRgpSVpF
Eemg9PbDZKoIoDzH0kfYCepuJlAH8j7m/98Qx0Sm/ukZ5+dsfiKvYxz2WggwHD+UGuCD2IC0zzv4
ER+HEv3Q+z0xtk3ff4VBCRy+GoeYOkLwssvLQcMY/Ymajv/ssNYtKIh9EtqNXp5m8bnri7GZx5CZ
J6ANxp0iNCJ+3zyeTL5ZKOCyIBNmCNXYAkXETEyCl+tI0ediqfcKOYGTAOQ/wJAN/VGUjGpmxhpJ
pM+mdAPN2ChQDipdyDHSUkeWcJT3uFSS2KxTO8PbF0EUJl5MfCkz2JEPgVytyXLayO2X5MAyIcrr
PlJkYFjwBkWBsj5C8/9RigXG5t09MGRzm5Bf+JL3N4ax7YyVrfz/ycqwl4g8KtC3mAIJbuK5cHxK
Y96i0bVB9SneT3ttBpjqtG9zzVv3BR/ZJvAlb565L0fgyf79GU7g4aLK8r/B429w85Arls4X4cgd
1HIcnB7Xz3djtV+RruyVpheGxRsqAQH0N+ueOnzXWz1nFgnvLcQamWdTmW04BrBAddFSSMpS07Sz
D86PJha29kd4B0FRvw4uAbpwHteE0/cF6vTkLMTTsyehuzQmXvWwSGDrUlZpEglX2CGgvJtRchCN
sjBGujl4lyD5/xh0l2xNU6c20QhJI6ADOFVNxVivuIyJFyLY+TkMJqv/9PlnvBYkL5VLj2j+vJTQ
z/FaIAPl7ufXPzNEmuT2xY6zwSUz8GyM0aH1lJ1rTJ6ips8uh4aiB0ME1ax9NK6/cufwnH36Gkf9
9+RugyjvNhliKF8t34WC8Q4jx0lKezPdpsKL5rrCdpfs5qVDAb8fudWeXMnyPWhypZO7tgPqEd5y
+rOLVlbU3JQV30XlS/79/tb3kS2dcPuZbZIbPJStp8ZiKHUx+gBhlIQ2jigNUf7PQfW9jXG0vDbP
0P73B4dgf+m5Tt+qP734YSdrUxFLbsGos4J7CHvQ1vWmXF3O1wGb7YMh2eDJqs/aPSIjTJTxHq56
A7z+JaDXaH50DUto+B7aoKU1A2UHkI3hBUxu+9AnETk/XCJc2ZrtDN/jJcRSdY566aREePINHmZE
NLGtCS3ulZ7Q5W/7quIjEtIL0r1/d9sbSHaZ5gCazVrDZYTjPQpwLWeC7VXqhGdDMwa6nOpv0mzo
XKXnnr/g9S6pDDuA1efrARKhtBxnWQ5azkLSb2hd7qroPw825sYwwlrGpdyUDrVHf+gX8FGno3aL
HL/08Yjv0Sd1Q4COmMz2AiUHuDIfkXGAEzfri2CDImD1csLUIUQCGXcdG2WItG8CH9ZCbjDOU3RX
SrGv+BiiWP6lmOR4Dpf5h+RRumLP7feF0DNcJtrukgdo/7njX/Ry73td1pC+KQVvLzSodsPNddci
hSFonGAjIOTnVuyLZ1wXuWKl4JbvSQUAnWgOzCrMkI1PWKkQTdnqFsPlBJ/DL57MW2248EP5OKDS
8F+ASN6qFi1lEFv0D+ERUhNhKurd1X8mOl26B0ag3fXiQL0T+2f7FpS+Is0e7sFMnw+Rt/LJMWUY
EKBDNSuwvon5pKj1CC9AE/Yc6zuZDkTVAyPyIsngTEcjKOgQblMiteadl1gSlrK1vGocR+JNl7nO
bX10NBOWqAU3msL8nbPeGK5hIWnel4cmd9XAZYb2CGiyeif4LUJfdLgxSYQYJ6VT8J3+ixzKCrvJ
fUMpblX3/IWVmNrIewVCf4SaILHRYnbdilVjtQQgF8bq+/IhKY7oMX2WGmrUotOFvIXC5AkQ57YJ
cGaldrrkRmSnFKYT/VT9Ut60QM2F55PMCJC6zPlKqbQcaPIkeEm0RNy7Epk2RUBkUu3snKbJsZTQ
EW8AzFiG+u99XPrxEGAv6BWLaxDlTd97ceYn1OvG+ntl6HjYKRBCABB6o/T7a8W0+cdubkXlP6MP
3A+lTUnCVvV0mtQ1BaAR3N9+aP3oN9qHloWVsp5d0dzL7TQoy+BEUVbjdOnEuZgiNwGuwScgJa1n
wbUEh0oghIfiqjKkFS4gemKGQY41CP3HqkxEae/0aG+iHkqzPYCOW8kc1yLLs6n72pTHTBytZKPu
rHH+TTBBpKla3ezxi6v+m1HCvk/xyzj1KDRx0d+UjxTGM4kaAuNcdoPCaqOi/ZKAP+3G7fmyqSYI
Bxy61kFk/kdAtrdm+nJ0ypU+lrymtWP7zgEGvcj8Wq1u6IazHmd+kH12MGVUzsDgto58wh3HFheN
7q0SLUsQK5gOsbxiDtW13UjYpTJVrrhu5yYclDqI6JtJSj2JKPWagY478bMTJ0fYciQk+hfrLX1u
H6MBcXQj07ZICSpEiGuN+o7iWP+EEWkbYl/s8lH1P8vWmeIsjexvrA0z7444dSRnTPGGf/MaUboU
ZKajGJILL7HUjXJH8lOyXzUQ6x9UkjKCy8vPw7+p/CQViT18WrhveiJqXqJqhPhPvSR4rD2AcYy6
VHoD70v60u9kIqf2sPGXolX9MWAW7WnfFFEm3YNfQBi8Wi5fBEymil+yLIX5wtWrQvixNZPtmH/0
djaj31od/3np6bVyyrDj1vnfevCLvyz+p4VBVemKwBedfFhQRVWwWMj1hBuOi0zzuqxmMGBcHf/n
pvFRr8Qs20wQq5USBlp+yld+P/nE3eQkIjBiuEG1r4VQ/NElS80XJTpWS90ZfhrWSpZifeQj0nze
WD9vnxIndynjcK+dnHCjRSuXOJMI1GVmHLRstrj+y5r73Sq3FJ0q04blVK4eLhnJgn698hOmzaog
++2b7SkEm/VeAxogj/Z/BrjMEPkE4KHZHo4et1I0Dd15FY8IJI5p4WU8Ay9daaKvitVnSsCL6YXz
MhaTegTQ6vwBDLM4WK3xWPCgsDddfsYoYRjmmcJpB3lg6UmU37pOdBCJG8DIZnAQ7PyqOWqHgMKh
XWo14oKvRIoThE4H83+1Lqy3/k1k+T2sa3ekBupfzMStDCCuj2x6uwk3FKkefUpwwjXE0eG37uJC
OSAI+1tP6X34RGp4O3Dw9wPDqxqdBJbeyTtvy96n9PpE327YizZARGBe78WrOAhdN4VZfMMSM0Ii
ZL3IWs7KtB64cH+aIQV4UKbatY42yFhPbIYkooVdExsvd3KJEoHSOphF6C9XlTvgFE6mLHdB4Csr
x+KmivRZrfBt6VU+Q0HhR34Hcz8vBLqi2fqk/4oijtPC3+VPv2kiTGfIgcG/q0l6M60FFq7p2rdx
2TSriiDf8NfqX9TafSWA1dOt1bXnN9M9+LbM01kGbny6jNohdKYuksZhi/PUtEYRdkzVkQdxP6xW
AZRPKIZNwqFFYL4qYfHe0CgXUHfeS1aowAglLd0tar0wKCmcby29+o++Y7/Jxqs7dIzfnndzMmrf
jqIEeMxdLPToIcYpb42/8iSBpg0Ihsxx1GUd/ZgSzdoeLpxKdpiekcOnZRdYR+wen8Ogk+kLMAyV
Yi5iZN3/ssYBP6U2Y1LzJW/M+Szx9vO5AO9Y/nIAlzQ8tkem/Pd2pbCs7avKcyRSDlDIjBlCE7jr
enCop11nYRgNbT6CyYzvu7gpIfNWdu6Q556D0MY+OV5Fo8EJu5og2MrIjPhpspu2TOx+huGu2om5
9IoaZkPjya3oDvQGajK4RWeEgUk4jXOGFD0DMB26vWDd0ZzPI+qMPUaDT9yvli4jYQleWB4ZuIMb
ggSvJ4lvVPRc2BDBOScm9VEFj2y4vlxzWDNuPwpChfdhygl0r1zE9q0D5zMGogk5My4Iwg6HuSVa
QnL6XltsNG6ahUx+kk+hwOJHwz7Ap+ndzyBlbQRpgF2MChPV4BFprEQk4hW1vsvGCPEKSeY7KCQn
kCLs1A+W+grTwaFTFDs8xubhJgBQWwmFAASRaFhoccRq6vVA3yzTDgFgZT2HhG1/K/hmgKNZX9tC
mXaLG0zXgdhSFIWn4n1Z7HPsed2x5f++05ydJPxGiCc/iTQC422ReUtgIZgKP0ryWhCOwlfJ4nbW
JSaCbLDWIs17zH6YOl8xpm7NEMtjK66ooaD7uNqj/I7EORVFB0qSI3xAoE29S2W0DMKfDou6F4mK
Rc9YojA0b1AWJjk5yI+uJ9oNX9WMjYOLbtT6dKg98S2jZZQuhVjdr6XNAgGEPcDbBuK5IoqBwjGI
pqt0SZ30ssbQufn2GZxP6Vhl6xURnuVDVvRsTyGfe3Q1xQit6CqTZO7EyO1F+MJrDYTlzoFnkQLG
wfqIwwvAd78BQbHCyx79gVVhC8ANJ8Xi9kz6vgAvGqPJsMsaRtxmE73waubVfKcAez1AjEYd5f8Y
ti9/6LnpPVr5HPhinFJb+tHNTBFYoclDCoPPEx4dCZt7BMoSscBPa9WE/tEVTeW/uDMy0OE19N3b
TbyGc/CGuUZo2+qybtn7Cfb1BHfj+RA3zuLlYYc32M4R9Wi1QuJBDmbUFWod3krkHuu5aqppMFKf
MSrlOU+wIpSPIA7Y2OgPCEfKXSJj7eXQTh6dql5XMoTicuqbCmJ4ehlrI5YXeZYl0e3p/Bv9djsM
KZp92J1JS5qCftavqIWifLto8WM4iqNzVPVFzaJkqfDfo2pVG7I8Dx8SZGJ+qJVBRt4faS3QnNA+
yxSWCtszyXOPlv/abpqVKwMtJ526z5VFb9MOlcOKWjGR+IkxPhkPjPB0KkkoqRtmSwU8SCdUqFay
pKN20/fl5mdza8SnHEK9AXBBQXJUBQe+75NHKff0zTBqBs8BtCGEy0QgnrakV4qWGKLLBfuLtHnB
Ho+qEZ84LvYshcKjHo0KWO2k4HRiAwezxVIaN8LnKEZLP3419xxwubKB+3GvQTcto5p0McjdvSUp
x4Zfyjh2f+NUnIISJTAABRKscb3eK94Srczf1vJ3fQ2R2D94wWwoCpck/Hi10jyjC5M4PTKir1z8
zAycsslCOmf3oiMC4Cv6t/ZQ2g5GPmINj3EM0Hwwn2I/471zs0/b1BrT4Zvv9aIN+mN8r95hE0og
I0ZvjpclOI+za44W6yULQ/Gwc5wyIQWZSfWZ9csQyVQrQAhs0HeHnYd0nRU5eR9cmVTRlvqdsPce
Ri7CJTBnn/9OIzZXmqJanob8C68azRYz0KXjje0FwM5VnrfgOSDZadsxGFUTBv/hcBx3WBo2Nxi9
S3Eef6SxRQoh5w3mARt8vbgiQMXGNlCclzIMxo0hw4Wzm6zU1nAAofhK9tazgpEjF48sPDYAxFg1
F6bULe3RXEM7PCgnX8VpPJgmZD82bqfJRuT7rHZT/ZFPjLGGkkafzxHMboEIcXvHryP9qJTJSqS4
Xmq5zF4rwja2q5eY8TNOg8UrSdEWhe7u/UKoLY2xQAz7ugwnzl9a9r1L5oNtZ5oNxzID9Ct/GEze
iWqpZ48qaAVFqKJezIiv6IcSiZ5BNxJcuhFAIu6XYHd1ZzqA3PjQO96kVSjmhUt/hwokKV2B8wsV
8dQagSA19yv3DbCxRMce/e+Ikt1le14wtAFn3XrEmUw+Nap5t8l5UTq0Wqiqu3M89mpRSOa3x4Qj
RUxshYD9WJfdtblf74ciRWmeZtaBhuS0y7nZkS/VjIpbGD6cIeYfIHq4L1SJmzHodISsY6WmIs5g
TMtrW5IyhOssKIcgJohjtzSL7hhaWrEYOIVEz1cB03r5Ka6IbwtrznwpEbZjlZujXtzX+JuYVJjg
g05kSw4ONzMNzB7iOQsj7XpTsNkC75ZFX9TDcRFdKPJJb5nVtyB8eTRlTXzEq6oxcGtcR+sLkKpv
14bu2utoG7IbI/BQS0/VPbjCorK8u9tKG3tmBrBXDVaSzsIJ99SVoU74IO4e1kG5KHS4rGugy3Id
bNIKFY/ksOHn8PNQhQCq+scba7KzL4+82Rq3UfmML+/JFYv/cR8xEynFTMKf4jtonzFg13ci1X5R
g+m2214htv5jVmtblKvzUfAAOIOMPOiutZRSZdYkw5KmmISc3RtPuxpK/7oamdenpLqSvgSZpJEv
gz1fn65lQWlag78T3SCJak6mUM0Dv+aJMMRP7ilpEE7xHDQirAtIMoBbZFnXBhkEXjB6X3iIWm2g
0i8sAtcTBRZzOW+kgH3bKFw6QR19zC5u7BGc2W1Qi40Mai8Wz3SEKlvsRD8vsB8WOY8SvXhIO9JP
/+9Bvuc/mALeBKmjtT0UgTR8CywZBVktcS1uoUMrz+rvAzU/0V1bgEaP7rEg504yvgvxhCf2BSjD
0Vj5lR1rFwwJlkKhva3FKM6il57EEezjfChxhqHyqV3CzdNxEEhh1VhNsGmFOs3erF24IXtogvsU
mu8gwpXufoeLI2ZmgJ5V1VPEQ39iM0imenjXKFNvEqDAX9Z9Hv+ev3E4WaOL+hZaXY3OzjtRI4jW
63doLa3AGZDiKBNy0oNBxLDLsNxwBFh3P/HMaqeehoA4pzX6aQJZqkRp1MiKMEuocfiKjKn4CqCc
8NC05y0Ewh/yQ1RtnV6rFG9oloKvFtyxsulqFAvXBlXjpqHkArwfGLTh9QWboNmGBwB1kTm9PYUo
JdsPvYUepyK6OSAruPw+fsW/iUsipXWexQGOaJTKtKTNVtp4h+NnsGxIiMrKERNOO+kw7x/u5khO
YyXWGaUYQHhZHHQ9BCwYuGmTo8qAHC46WMwZ2FKIISAcy7mRSJn2B0DbRo2XB+JZruwSCzXRv0nE
b57aypsxjupYWGW9wAHMpfi2oMAoxNOZVpBcPF1vCyh9dFFr96QcAClf5avwhwyxowOupYXCto/2
Dqz2vi8OkwAjiBw6hAWvc/WUIxhpyn2G813vJA3hI3Y5G9a6g8vnKR5M5yUUgHXJ5qcplCpbY8dE
NeMOErq4fbVpx0dJUoQlNCZ1sMWpGj7na3iElCyi/YcCGn02oNIy791pkE23XIg27CqlRrr1TUsX
6WvUhJ9RsSvZoeqIUuJQdcSpDce0MtHsYOVnImZbAsXwLYrsHA1NZDTp4f7mg2FnX52x8lLAUkPN
N0CcC+zXkjMvwanbvDPxi2gPNj+0zFB37qpUSMh2y4PyUedwRxrhk+0tVxlHEhQJtUwEWDXD0g9G
zFAeJJ7jn38y8qEvNGHzWz3huWHr0+XV9RzeKJcBIO388WSp6eIf8RaOmiNYSj10tfoLIf2nhDtA
6EGsVXwhcMy0OqblH823Jo0z/xACjmTBd1NXKo/DoC/tlt5q1ibx6ky2av4C0YnZ5rvpc+/i0WwI
EBdDx9fRuxpJeH6nZfAHyN0GzM6VDuXW/MH8S35DJeOs6ivhwfLt/W7r7HgXjdTK7E9HdTBxlQtb
DBs+jd8zAFs2lsqbsyPxQSxwwZ0bEuTnz4XfSsiXBy+LujF+3NL23Q0fxlJ/w9Ku02MXuvL5W/GA
7kn7zfxPS6lwIjptKr5ZIm9CvKdZdKQKI9WfN+V+zxEqGaMVKMyYopxHk24AC8Zf1uSLDp9jQYpT
YHOLuiQda/AXSdR9Cfr6wErDe6ULR+MpmKgbEyJQGJ4j9UmrezrqsAI2Ix7M8IH0DNp3JqK6Ux9r
fzib9Uh0yTiO4C5zsE5xETNkggES6YL/D5B9kozis4eBBZPDNYqxiSSGuT4ePaBDO+4L4IRwKxbR
SRipwOSk2UKf94Ccm3Cljx9AWU1EkiztBnWYP2kDVb57ewzHTPi9m2TfFQKwuLTY4lvBLU2iXTX0
cJ8Am9bEw6mRfudLCIGDHJL60p20oyVQuAVGab2KmGvPeippCW8HfPNnyF/3XAEgObVnX/S3+5DF
1MpvDjYlo3NuN1cV3WRWhFLMgR/cBV0dfUqIWQztc0uvBO2Cjtkzq4mqOPtkmhpjWmckbuyMYdGJ
h8WXKo2UQJSW7WuVcqVO3mTqBYb5J5a5R82KV7WELW+L71rHlluw20ENWqe/xvV0Srh/twpxxY/5
Ijt2ku9HtSQZw4GUoIlW2QRv7SXcvUunQ+J+TUTdY6+zVuALuudKAjuHNOrJSY4LINdFMSOYNZ9c
/7B+/O0DE0VUnixq6pmTrfa1yGxeBFZT8iwvX2BlbfbGVjXQdzJj/jOjw6FI5xOsE0+MZGpynXLh
HpiKY42SrkP2PAASShajxlBeQbeUtFfFHaEb+EgaTxxcxXzaLrflZy5hQRcqiI2Rnc43kLxPPIAD
PEtK58y17UgRvXwhhssWiGUX5ybeDfbhGs3xpjuU9UfvpjFjUV7Ug5StUXVMd93w2QUSzpEByoKD
yB5npyUVc1T02ybfevSck1c6Ra7+WPFQPofzd/GSqBEyKKLSyvPhYC9J4kKxMeBEPJAFoQ7avZ4y
Hl7xO6Mp1DUlSobetMt0tUExqLZdEeqDvbVwCK/FqTrOll11Z755ai418OdMdmu5Ih42X7oxAYfg
WNIfWlujiNxR36UKn6qosla9Ynj0wiFhfyQAzwz028IMTDGkGZennYXMMr19pbDo6vOs+2FywELK
crc33H7BVoMOtPdPFa2opIpD6+RlEc4KbUpcwF8PlifLw/nkRULJ2INKICIKu+gOpQKweHSMGesz
OUhx4uBcVdUByh1cXteXXZjdsPeTSJdpEM6AtxEGbszJjvpn45Fb36Yrse8gXJq+JE+3W0AoydH+
tsqbjJnP9h2/FXyepiM5eAR8zfJvlc4nn7ZBwAqQL7RNBKTduA2lnX7uWCDQrxx1LnzdyMnivVKP
EE3aGj5F6K4CvtU5kmIQQrbXzCL1SQQRptP0e7ES1GkoJjQtnjTpd0WCbxAuLyuS9bSQcp6pDUem
XHLezesgeVPMbpJnLAld8syrW7FTDHAGIRVpGr7wp1FwzdKs6u7zti42pfVWCU6J6YBmHmMV7jLH
NOJlMT+4jWLjfnF066TWlxajO5rKWj1bfWx8zEdiojWpbopyKfyadeVQqIeqP5AK4YWO86pL8dBh
J4uGJdZTgqJTG5h9MCdfsYlNtU41d79l3T+5CZ56/aUW4T49ojQKqSCCIE2Azz03W1B5sY1Cz6yx
1XXnLhgbxTlia8TV3BsWRqNyHoH9shqKbVGveIouxYlCaTEGnIV1xs1jBp6/nFIlsTbtrkA3FJjj
PgfJhvbrQtcojtMEgmEhKYB0/iYVH7wRPvmOeTtYogrJfhgCG5htRAe7sZA0XLS67RA+P5nnOneH
MlVrF7d8UoyQv0v7ijW34+4U2rJwIWfRruB6admb7EVXNtXt9fx6g93k/mulHja//j8sAYMJWzho
l15RBdZvM/jF6VqPI393RhhNSk5o4kyFUnSGIa5rvxPe2FWodVeV8jf2bRu4iBHzb5ZoPcpPMU60
iCJABApoLw3YtWseXyhcrQe3nYjZGuwpKUZ9pTWD63jeKO2fSCkQZ1At2KmecRVfgSmfw+aodXlY
0nqJ9n6RKIlr3+rn2KT4yJi6sCv7w1cB75YyDD789j71DnG2cAgN9ysJTy9N8Pjvxrkd8MUNG5VJ
WMut61T9k4PnM4aSg5UAClkMhGllcnhz5PQTu/YdKyyG9Oh1y4LzElrl7ZB4CJibTWTf5Yef7LT4
K0TFNRXNELzJUGl+tVFH5MJEb7RcQiMFolOpt0Uvqq/drBcK18qhelYZ5QJm6C8GiMt6FuddyFvz
xxSxZTBU2MRkOzcGYMM86TGhZNyK3TRAzvA881D8q6aaZ4MPREGCY65OyD6qa1EdXyYR9k6qQqqj
c/k6Qb7opGRK0bh+hhKhQYyf14JOf1yrrcya0CDr2ivPKIxlig+9Vndyy99rojqL7jHvugxlfHBZ
xggCFQ7djG9wmMdsVhkWAH/bML1G7qM8HNtXsJfOZ/ZX5277Z+zeDXQsPK9hl0BPpPEUsC3Xqdgt
Ww+nGBgIstV7bll905XryPBgeksxf0cOFD/st9ClsDMEXsmwDu4L8O3K572dfdJCal7mZKk3HTtJ
cDCz3e8WbTRpP52VLe1cN8CcWQAnUFEkBqgwxOzGbW/HbVq0mpLFhBJ9KDSPBfWp7Gku9QDU0OCU
aL+JqxO/pHtVToMpwPnzCtYp6TX0M+KuLPSFraUFZNNDn4UTMfuRfSQbqNQ+DnIj/G7DYypSHp/3
5bnk/D7pjyYkqba34TXPLik977gIzWkr1P2Rii1N2RJ5N4EPaTUtTZO9kdEPyfwfcSvTnyeX3YCd
rTn7sS0EkDrpkTq7M1R8FfOFA/TS48bXzyb1c1sD6qBT1fLYH3heObs1SAnlIhMtz7xk00lTIz6P
bM/VlEqP8H/gtICxdeQfKQpjKRjVjKnezxDT/Vv8b9P5cWph6O0XGUgam+qkXQ8VVdj+M2xpe+eZ
sWi5BKAaFvL63seO2JNxyoNINnKbJ35d4hzJmsf0C25AcTZjOHgkiBXnywlJ5bQq/+NUVJgZmHUz
jBVq2CuNMuRNLGtcpCbuwWnYMzVqY8+Pu1hzFmjr42CxIRivQ/txZd/T+DJKUhRto5LpCtNnAsC1
vXFBc4nEX8ehc98jZ6EAjjeCr5ZvHsV/zQrOef6kVkLYF+RlS8jTR42t4GX91X76bxKNehchZ8S3
KJceaHSuYIJgldDuQyjtQRz7p9b8L4JD1o0pADfY7v60N8TozGX5Cp+3hN08afCPsXDsUc93g3vW
WMPY+wUhmQVKLT3LvLe6buU0QI2Vnu+MiDhh+dxfrHgudj52LmJOLlFXZalblZ8W5I5ipk2+NiSf
7iq7X0d2Jsx83qBFalHNMM9Q/2pklPIMsGCgCRhiGT2ou/WUMwiXtC29Y3Zq1ddUrr2etcqtR8rx
0dpZXXgL123h6DXuLbsM84iMpPpEuHmMVdLN3rNt6MhNA3L6jOzh43j5F3QRg/hQB5S9aQixGmQ9
gZQIgfrba/UVaIgldHlOgLDlPOXEjTD3A5eDL83MpXr/stPNg4npNX0mwbNHiqhugYu4e7K71BTf
39rgQVaa0TAZVty+RBDq3mZfaLJMZLiGu6R3A85+ETlFM9UD+oa1dppSkVzt/ZuMlh+eubJohZgL
skUWpcVzhkBFg9YORDLGJoJ9KsUYMnGVgymlEBbMpneL7uib35zxU7yR2GfnYVM9RnOhhMMrV/qF
RZKHgwsHq1f+fw6pabRHRce0JzhEAkDjQsdiyfopJ6XGPIc2nF8d+fedlnLiynotwjA16UUQ3v5a
xTdWOQFI1ELEBjeq74ARXmOTY1HybSSzHRfNAId2p/VVPXDxmbpzcDOCON85JZqsi/KhkBKAHr08
XxyV8JT2CNV04jdmDGvxrmX82Vd7/xKOOy/Co+9eM3kDfiXdBsWQ3jTPViWQuILa6c7DUvC/8mYQ
hH7BJiOr2ijYpjGfliynYX1k2r6AZ6M+0m1Tynm3ZE3OaXDIL3cV3a2h/t4PqHuI4P9GvqjOz0GK
OoXjCPQ/OkUiPNXJTSCA/pnvrnXXJUtLTJMIXoydRnz4eCMdOdOPl+kT0ASSbR9gQ84LeCs/x0gb
7Yhiodew2eeDE36TG4J2+soCkRtwY9+PrVfRo38wx6divnfdkoO4yYHl1Y8M5+Ud53xSwqyv1CBs
/g8OhY+1994ofX5lxhBswwbsWcVvCpOHv0zQ9oG/OXk9oTG7LPu1ATJcOo/RFQxg8cGLyjH2YbQM
bvWQjZJWUnuN0EnK9m+lN+YlCaAHnmvTVvuhEsySCOSxNaA//11qM8uuitE8vUTE6BczHql+wdg5
IwJ01FF17CBITu+W/nucM4928HwnV94DnlS+o2PKM6wkjShfr9S3Rc4icD8Bi898Z4TZ/riWgvjO
xJDTlfHFs9BbbvaFR/5CwOb+/cCWqTGby71txLqOVH6NBPEK1w1/87nLleQ4lHMuLcNp333l38pv
Rk2U8n+7TLKS9yqV2uW9J1hvzAT8Oecwy1NvL2jMuEnNyu52SUGvrSf9CkQmN6j7vNHO1isLKoP4
pwHPK7HFDrpJO4DbUKcCfD7wMH95Cq53zOjwAPAij2J0agZ4GkQ+GocOy6vIirEKfygj8wXCv4j5
0nXODcTy2Mb4eht4sXtAFHAUmIxhAF76eM5LtQIQ7CA4URDLrGWS/YkDtYMjgJurlITsauXuneip
fO1XWv/Pg28bMmhiHEq40ibFr+rktWrAA3uJoZ8dhD8Q04ytbC8f6c2yH/x2LSVhI0vP4m7FaJcW
OkTTRV+dO21ZoLbQAzAgX9Ex8idW/5dvHsv6CYlflAFW3ec7jZNURFP3a2+IACF9O3qwi6sp0XHa
NHXA/c9XN+1sMMpHYo7xjh5oO32kEtmzpZJgAi4rZvEMNl8RCjpTauDztSAwxoSeW/iERM0mJ4qZ
VyrMvKZIFSyB+XKg9X5OpU1vTKmTR2iov+tVa/XCSVFB5Iul7jYJWGaEIsKbPbOHGxrmB+tFsf9j
qowJLIc/+N4x03XD/omluQcLnzE2koQoFCrPOM7DUj5v70OHEBPcXAp1M1ZQBcrqRhNI7bzg1oKG
kmVDPS/R0t4CTk1lHk9CqWlJejeA4eZxai1mA6uxUSLYxBGd0vBXbjF0zrF3XHsE3ZRGcLDYq5o1
hAx6y4/zOI26IxKZoHO6Z9X/ZmstxQa+IXpYxSN3xlOtgtOgpKJ/8XS7jpEthwuf8zJ8rr3IqCeE
Y+tyoq40Z0vS0yruAVQp636N5DSTii5inh8sbjrLiOsJank+mcx/uakf4CqbPKW7z49T6oNdA6Ds
2i56liV/ibLW671Gkg/PEWdKktIYiXvoRQhtLJ4u7dcA/gRWOiGDOGEvcG7BGKrsAYu2xkd/DU4p
r4Bx86vsWk7TqWoJcmAmEqDWazKYwMx+GDqldCHYLfr4gCSDysLpsMaXH3LfvqdNV2Fgp+dG5vSH
5RMXdMDrVMcRf2i7cJ6Wu9hoxPL4VZA7arhQhtc5cX4mdF1p0iczRa9l5nAjhPJrkY2XIX4TWDJz
k/ibo+zG+L/KppCAaGuw8PhXoqOr2zMCyC1eheyrQjrL9WduGbra08U8Y3CZTYuyiwRjv5+yWrBE
Ge82t0eFT2wal+cAPbK0hOWe7IVwqkQPI8kDb1pfZWzshDES1yUv2qHOU64lEvgikOxyXNi7h3Px
bJGfcAhTjUqyBJevHV85nFZmMPt4K8I/E6mtnCqzyGGoD68kvlAT2SBb/Y/us8KPycF1POEeO/sf
o2h6Aa3vXsiOcoZvqHPeEZaN3J/cI0dX6SUYGkDOn+h/9IIOFLWateotpLGYFN5uuw8LPD4AG8ri
JHcf3bCMspYvpNu1iggbgeiE6HHChoRGzRjgvWiIFybqzXddYdsGLdUQ9zOGpxXPpJ6uhDvf7P95
hUIwX+nOCKUS3h8KckX/AeB7gLu0hVDccdnbyolmvmB4+QniaUJzOVf3xVCkyQobdF3iaApD+Jci
dmmQ5NPURa1/wuZPcBA/IaPFLMeohquvXbNa/atZNCCzvM+2VSUU7m4cUNY4DMgFOHSCg21axPQH
fPvRhDCVcwEWKzi9/8PCdUMT+a3ex9tuH7XQv1wdzmiMXLYRvbjPBPA1ikNJpF4M7TE8VLDY2dRB
xxlbrj72RJBi/ZdJPJlxvS1Gj1Yc0mNNSOPQrWVB4yJW0ySPSXCjUam5xAs/pTNveZ06LW9yYeg3
rHEoPGGXsx1yF827ltVpM9EVexeAVB94/LysksyKYDHaUKQPsmHflrKqTzn2aiYIrzvKeQexzGy2
pkLDQr4TfeP/ztf5Vl9rv0cdil+oxp6YVnz6TrSF5ADZEfwSPbeSeQqbEzjy8uoJpPD78tL6vGAF
ekrky52Ih6vXmTN+iR91vduPfC5crfR1gcYMbwGESjMmyT9OmsiKzr6tvd003w+OtAT6lgpiM8vx
SF1C9+WjQa7fGFVkk3rlDk5HsdFZehcJM8YqRScNujt0cwSSqpzW2AWX0iK2vr9vZsjUQ/w39S+o
l3jaJ5tUB/BHAOVNW/UdwSJ41pm4WtIASFconsAKWAU1Xg7NfCZTFo1EyLch88cO9wDCqbBwbY+w
YOECFvZ51O9iJprLM5WeNDciDiWSkf5bj5E19vn7ZzI+HM9glCv1PZTRazx1E22V+9Y4wCoH0Pkz
++0tc3eTgGZlLInXOwIMhYgEYhXStD2DTRMFdIfBt2lKxpbxckw3vlS4jAmTYfzr+9xkLiOYPPFs
jdsSac62MODWhG0zMhmBCh9besrkcJ6OYuFi/fuHypxK0d0mUqR8O5IOjnbTAZE5TIwv/VNal4k0
ewk79FT8T0kS1tYvTg6k/OEqgu+G3psxap4WGxJO0eAa1gjuicyqBSgfKB/vAX0h5QAYzy2JarfM
mXNmDDFI2bMaUk0OY8zidwjjhiZBN7krT5tX89TAA2uWP/4tCx1jUzB+nIEdLlJDrWSDun1I+fwM
MfDvfSeqdiNVwj+5LF/X4DQ8ymGMe3wv17p9yni379tXKJXP0C86McYAJ/hy0AGAHx0ndB9tko2A
zJlyE3kJIpEVSOghkmyvjWt5PeEDFJAxsUd/s2+w10QnFTPhkscHcO9d8MunWAmPpGW2kTuD86lV
3VqNqreBbmyi7pwHPGwWaYpg8fVTLP7Dfr1XGzZhYAq8Nx+20vDnPoIgONqKJjKT00ltsUDsP4gP
+NkKB5yvCicNfSFmPQ5MSArmkj8JzIFkkXdzIZ6C5RpLTYIINmbInUYyS5WZ0czuUO7SHX/MAcIr
KtEehCe9vOHcZCjHl6zdQ2puVM5HyPjyCrNc5a8MWRq/FwD2bI3Bk1D882pARDVRB1YlKvQmQwuf
zqU/5uVj5r4mhB+zQQZgFa4oFa3d7VjVR4xiZcN0iqgNjwK/pNkgbDdInXX5rqhZ8bTFzx7EyMGV
HGA0z9Db+7x86IbohtwnFxz4e4G5WHpLv6dHywsJEcmFeKai/e/jWjoNiZw+Jkd+ngJGgShtFqBK
5EAWHXM+C3+KPEsFbqnH9L7LJise/fV0u2HRxTKi+EEzkUy4rWqYyUpn5lBzJCTqIEduaBaJkE+R
8BM+7WfuP9Smz8nsvVtvwAk4BzQAvdPfiW4vSEvbWzHdxwNwvxoC8tvwCGjYK6Msh9uRWCwhm8oz
kz4+SYnYRqtJtX0ObERS0lHl6SGIoMq7vWm80mHMHMb86ViVabvBa6e4UWo2dgA8EnQf03W/vdfs
yA4swfSKG4CkxIJZDVhrksIXIaic4x9qfkW16CecD6o/+se6E1h5XYyzv7l14PovbJqd2eq/4UHe
eXQJ3n2o7iuDuHFKkYWbnPfL7zH0RbP62DTUqt3OVeGNSSbR2Ws+o13/yxewoIQ7RS152QStKIwO
mZ8DeQF6th125NYO4Fhvk9CpKnWgovFHEyfgcWqVR6OiI+rG3FIap5L2N+nW2CER2Rt0S/cfokPt
h4HfLLNhTk9m+EN93ULo5iFX9D5OUik1JKMs5dV1AQUwyqA+xyHdxen7xy3PfaTDKe7iTd4p6tlo
y+VXiPQ/RqLod4uyPU3H5bE+VfuA7C/NHeaQGFwn7hKimOc4zcLwmB0GsmXeFdmFSxzni8knWq1d
Xl6NLUqMDnZ8Ctu3qrNC1J0r1tDpL6Dj9gpO9JFaJL5zmttmu8X/4GQfo7ALDLlv7TbMjS2cZ/Wa
TqgJKy9iaUi9MuYyEHng1LvBJ5hNmA6U91ADW4Jufg0q1RDvubQsw6cfC+u0Wnqy8ZPjuITcpqau
WsFN+tYPPoIfKF036F75a7kCTfVLFhrPPgynHnXrD4AXD+TXsn/WtGcFhwe7H6hYXjnrjvTAf7WI
1v+WM1+Hg50sC3k3g03E6fKZnsvmn8mu8u54bWVacOeguyI5QP/LRcMjoX3a7+yDkzrRd940VLH9
W/NfQrUPUWsxZYprFRk4t4JuPEcpgoACIH7WhFVSPXl5WbKNGPN7pwhMU5Bz0xYQmkegnreltM3e
fPc1eqiM2pYU/VW8muXxF3FNnAXp4toa2bvjEFwqinhk5KhWcP+CMYKh39O1KHcMnhYErJi4Crns
AkzL4xRPoxqmsgWHEU9Hu7uJFhwLhn/S0AJu1BZO8QyyYV4PYaYbvHwG8E9fsXAVbMT6jb3uWdpp
alOuTq8mvmqut8IUMp6GRTMnjlYKuo4AoCbAzAD/QZfzJxnXb6K7xywArfN6rxgJbNboHxdbzq8J
4OrJPsw1wpyDEn0ImAV2i+IWo02ZcbLpB3pmLTS7iwUjnJzFVXYw9CGYk9uLELUd5OinTtZasKW8
OIGX4FwxkBvM2BMBDX0EVyrjkheHlxmGQP8fcMizjqZF4CgLs/Y7y5bq+krvIuHFCDPnH5gaVEMV
iIDFdP6x3eGUd8GjiE7kdaOGEy1kkYRYm7VCdStPQzCj0BruSvz0h+6uc7erQEB7YYlSMuiXpqSC
RVymoZlg8OdCzGly6HdJmxjjakztOrt5r23w1bEF9Vyl43u4ns9hHz3A91Z6DQ1qMEGf6JhaGwnn
YVotwIHai7S0EPrfP0g6+h3OnCo5EjoNK9DKsoy33izA8SXfJxt5cqHhuqdzGGIIFdshZcBrkuBw
5xCEkSPasYHViA2QGG1G/vsKIQ8DiW6l15XWZve94HHEBw9TzqAN02FsWMdMogOVIPi3IWgy8t+k
L9rTPH/u22IIdiKlrCHMbMNIJRsILoaUsWNyl51Lfko/XjZi+TUWeDi0UP2wFqrqZuZ3KKKSfZcX
DcnHSeaSG2GK9HTvWuoUVHYJ0DZKkKmG+/MrdzWFgLAm4jVyq1qonzRpwvO+QbbjUebcdKVXUHqW
A5Qzzr1i7RMy3Ve/2wJcd74prPxxU1U20Q8df8ij3tbmboeNx9uSxLXqnlyM4ekN/k1/Nqx6umV+
pkjpbn7OwQFYni96jVWNjIiKZfAuayTUT3wjA5pcfCXiaIs2r03ZUdueNUqcNtQDrBhygggXPh3v
bUPoZ/O25eqK8YxhPLDtb5mexFDUetm6oWUwxuGxPf53JSRDM9XrIoPmrdXUyWwMUpzQuUmVmv6J
2HhF2nNQ0/macd6uQiAGFCUu/VvosXjcgryy5UgRc43moLsGCN6x4b0kholjWD2O5f3MdMlBfUN8
DB4lAHao103ElkqYLaxy1Ay5G2e9W0QtmiD9vlo4JssdODXcf4I2uaW5GVMO/Gd1mERDAMRAv7YR
efMUC080EWcE0wYw3/7NODneaI7iUjCd19Z/JQvtANwLxFD2Gb/NIwrseHcfUL/Eiai9zXZj7NSk
BZXSLoWftFH0Y/1iZ3crjAIKA+XAC8o6tFqfbRuMvsrYgnaYoAqTy418sKstHhmMQ0dC6s1Sb/Bp
C482o39gBWj9BH2q0xBFawALbJC/UlcA/QXjVxwQPH0/WxVXBuSIzjukW7GoAlSJiFhzFILBP5ig
vEv+0z0+fPjmbTemjp4bSYwKD2vkV23SjZs2L7XxCvBEjLlvsh/mw0756AsFU7TXLb2UbMRKJDAq
7OUW0yxlUqwKxhsTmrlK5mHbfeS1EqAiJFmMd+BudTRMUYukWGsxX8SFSkapBGDKyUdMV/lnw88v
GKfPBhcilCqb+qb7v7vXB+cP4urkuohSxKarIpW1W0YI9Fo1iyMTnUTn20lxlGcTHAiZeSc2VnUT
QwcWG75PWfglY1T234jQeDNyd5h0wg9yXxSXPKG00wQ59AHPBhdsCMTGrUsItWdqQU55bPvjhOr6
QT8mxeCDAeeOfBWUXvIRNTxINYvvIC7Q6/FgonsseZobR/y6/jef5Hdxynqc+d3KX/raXZwhwvCO
va0PBU+KW70ndLlK0JrspKx/FAIu8xNoyozNDegqMzf8l3NGq5uyksMuMxxeMsQUCFPXcHe4VsKf
JcLn5mpOTzlydk87SId64xxbmcwOaxi1c2d+O4OJTcAlqxxbSNinMPPVnAzgxAAK9mAHDVVQOguI
XcCpNwzPx8op0aJDOdtLvKRlEiwmtqR6vvm8fPn+yLdhZR8OjVMoOzKzxrmlh/AO6S8d/N1BQEwk
9YUjTIjRqHv9zquYjB/vkxbMNYn0kiRkIo9sFuUrS9OsyBs1hGVbzVH9wXgopPgup9qLzi3Jh35l
FaQRTe4yuTq4IyBWJu1xd77TYYxk3o+CFNUv7Hvtp7+miD3NcEQ1DGEBlxcHThsIiRG9XIsAhWWU
CM2Q0mjC3RqvDGdNsiFJvIl+lfCpsKSD6q6ZxvCgd+X2d+g/0gX8wmoxONcjUFHVZuQj5wea6G+a
sOK6pzRxzQ+7u4LKdILHnd+EkIm9hEgnGQdo3ztn0V/pXQh6Bm1XYNaUKnIwGNbETnSAg9jX+taX
cI1ALq2nEV59u/8RVJE47fmVXiO7iSSjzsbzOS2Omg7UPl/U41vC0DojYoKPl1sr/9lj47X+/ACh
NjyncMq4ukIyLIC2lZbEYrdpRsMjxP2PszDPls41tj2HAMsyRhxCpYKryBlH35vNE1cI0O8JRJH3
x3VM2nvEGINvwHhNlt2Ssp93Ast+7r9jACUrnsn5qswxWIH3/P2K7u6t0gsgoP/RPuM23nLcQ2Br
m/g3rGIczCSCpy37O0b48vA3Uzs8nrrqP0+PL+Ew3JzWEZKEHsxxoQaV6eMRCwPfES+Pban++5Oy
MBO8D3tiqsg61srQQVm44UwldSl5jwjwkEhWXy88FfFGSrfIN/QIXj8dKlv5QP1oMbw65g8chNRS
tIcO1uGsKY05M/nL+M/9OM0qZWrv0Ouu1XqvhVb8UUqDpF3JOF9+NnTLx7JLzZ2M7gj/7UGlmQlY
mNRFqW6CVvDkgR7ZWlCjk2FFZsjF+YMdxlUo2QaOrZ9YnAdqTCrNyvx6bq3n1qW0/v/YppnU7z+c
SBqRnI54D2uvPkSFWqlfGEnYQVWoCw4fN4OfWQKoF1waJfXuHScqSiZChf/MjRGUQFbQAQeQbWvB
0UJUHulXG9YcVtYSpKYQ2/TvTwag7Ooi9CnKGdrn4YUXCzLBI+dPKjukIpXrQx3ruTL35At4m0Wh
q1Wng5rXDGLebei2SEv0gNg9GYQRD3mkedCHyOdbps/3kSVcdj+q77ZdclHRFD4+8+xrrGospaUO
3Ui09txt2SZ/xbKXhyO91GenEig7HF/3jzfWgIUI6SMUjqxBN28H2TyNNqnNQqrMNa0yuh0sWf9Y
bLxTFJyv0Q3t2GlidmWo/IAdlpd8KUnANevKSm6o4QYXGSlqRzXyUwleY7vF7ymPw73pNC6Pp07i
y6fbSYtO2OcrL+R+JzmyWF6uZWFysgIFZjl8T3zSglymWgVi/iUQd3tMDautKwaeOzJCUAutD9I5
vn72nNZhd70p5BGLN0kKnGPYHPxhqSJfUA24GDyTKBh9/N/1CGKdFCaDamwenTFGKtQa9Nvi1ndu
svAejK646li10QdpI4cG+2/Yefr4tN5Kd2fQkhp0Cr52qWLmHnuLQInPCbc8xU+JyXAcXSP+OUEp
UHtmGYOu0CgHIz6UpyNWGHLMDpyk7WE/6gm2nZU+Nvp01eY+QYbxe1kmwFuqtqKpYVUSLdePRN7k
Q8myUtLBm6JZsgrvM8hkbe3SvtJMHS+vVAIQNj+k2klBV0VWFEfabnBhis6tmQtz5UTqRUHdLRTf
BRjVAkBxY7Nl/4RK52hCjXtOgp/x3HtLpOc8KzQ52kvWEIafD/KxWXMO9ipI/XU0vKz4sa3fZvcf
tBnLOQClwRPCNQ8HsGno1Z/2cOwZnDJ7WBpVFga+qoWma5da1eb4YTrHC9uinsMIY2rJtDosJMUC
xTQgZ9esJXqyj5xL+H5WouGKxNqGnp22hJ0rAnCN+cmXCTFNkgEwfdl9594J97MUQpr2T6OkoYdj
SUsiP2wbYdu8gYFEf9FvEJS00LvAMk0Kx3uoNIjcNEgwKQQBGgrJKeomg85NHhVW4YOJaMaCtGWy
sZ7ehi1fx+58StK3ighdoN8mIl11eyfFVR0r0zyvhD41RmWusI8TTNnD6g7jqIRzPNIQ2nnfdKW9
RKEtfbyZE19efYHk8WvqLGjOguZ9ph4P+YjQmUP6o6vQKJBF6N7bUxi4WIjJWOiUJXF4rWWceBzw
jGILVV8MQTY9TBqE2hRzupSJ9AiSjYGmV1DHwaRvRnjRzguFIikd7gQKRuePQQ+ErdRvK9G15a1K
qZTb4OWEhPpgFfGuVa7KirhWDEucN5oJtqVSzl/o7ai6n9F13kmX6k5xhmEu7Cc2zliOAWC0yefL
dvwGtY4RPhydz24hU/JNKz7sUXPqCotleuOGyHR1VnK1x5LeRFfe/chhEv4EsJGyXqWRjZJhivrG
06ttJmbUfG6sYvJ31UsEZI07z7arME3bG0+3P8GUbsr46QVCYZlA8eu0qdCyxBERVDlRW3ysJjcd
bs4+Mq8GSFiHJmB+6jr2QNr0emTdNz5Gt1YT5BisMlNeogshKiFWNWImrhxVVVkhiQlK/HioUv5g
Jdy8jMW8uYrbR1EVfErArt6kGQT9aguSz8tazAE4Ckgc2Vl9cq0VZlP74O4GziUjoLUhA1ELzPdl
lTmJCUADIHkZU27m8lSfs6vf1o7KJ01Rt1CzU71CYcPcA6EU8fKTe2seYaQnozHA8x8lBZ+bHtkP
q3XqdaApEq6/TZlodbJ/sp/xwZZ1TKBl/eVp/fZAXOm/IfzQfxxk2A29XYBbIgG+Q3XozzY+1lLF
VwMx58sQlbWeDFBdPXYg6o1bcYYHiTqC+mIoofaJUDTInNyBAh4oSm8rc3GDEK8by/7HJ7gNMGhM
J9rF8dE60tP2TxTNjpZxifc4ScdNRlAAe3gFC4kRNLUed5V6710AhN1I0YKLcePJXJCw3rj98ylH
fFcOr4TEQAfnVwWYzRJd7ZlR54yQzNTfx0TQZpZXMGN8nFw9ClZOJXmyPHojHngK9G9ibC74aQ2s
SEO01k/KWE6i6bbkwS48xWht44T4hobCacYM50ujKDm25Tgj/XxXMFBeNu+pFeTFClu3Z2xISokE
WOvZOD5H/MAvrZw1QFSH8mj5OPxzg7/9+L2TsdiYUjf8WDfvhItrIl3Imyrfqttj5Ocwm7KtvktK
NHZdXY+Vz44Cgc9UiNBMxpMvDEhOczpOe1rZ4PYmmXbT1saAB8ovFF4UHiHV+uMX4VRNr9FExj1X
3iwfbk88JPwWMKTBzhZP8S6WzjEogNC2f1GKCBywulOsANzo6jLSzJXdDk4nEdxKehoHRFZ2NT+k
D5IpiVE/G2rBkCgufd5KZsIwCkfo8xKr55fZIEbHpcQKAi0+fxknpglfAaMM2CEw/XZjB6flUZu7
bMf8lGfjnWk+f2HAlJPIXAKEv7E6GFCI+p2aZunk9UD1cqTUQMRZNuhhsLgnAF1bCMaHZ6l2PG8h
0EXXe3/q7MUp/+hFm/xkY8d63LpPR8SiroRe/mymF1Rfxeizupj4nWQbiy8+ZzNz8iwlab30KKZI
YZNjKip1IP/9S82T0teTvWiL5CHZkczqB9Bo/AUqKqr+FUe5XzxFCexdxNfrUFiMKGW/Adkuo5mD
UR1mgtTxuqRC0ejsEdDZqNzN6fgCrc7eCHXNS3z3UctZYIMdLK/aB4asedS6leoDrn0ifBskpRMB
kdw3OHIXBh0FG+SFot6m1NHKaPQOfnBtJ9e7flmauxZEB5ppL7f0TNJYvlqP6shslqizKHgzszsM
wzf8mOnl9jYnwLycSDdUNoJ+ddZ4FC3ad1OiLY3bot2v5hrAD9gBUcKjK+cOBX/yGBCtNPnwOxFR
cqg2qjpDtP2ThBml4odPSNBKnfG7V+aJYyDMYP0h0T8QKdJshnu6IG5TllDnf0xSAOvxgiM9HB4U
cvqekNkkap+bXMi/pTmP0JHTWffA78qTuxaBQJY4vtnM3ipXPvnWh5gCYfLEi5a3TcmouWK7DZTx
JJthEJSoFp+2tvnmnb8G8AIbnwrojBT8h/axsAwpLO6SktXrpfXu1f2yyUYJWvFyNJM79I4lmNF+
yAKbdpQnrRzwHeVWI/oEPlpqxmNb0Ti+CJh2yrDmPBgCmR8+YDFJzJr0cgDNppodeuluO0NDWBUC
D6X2YQwtNslAu6yuuOD69HKCeuBCqINMrTnzO7xesjJut0GLChISHe4yMM6RkxT6jlN7ak1rya8y
qKo3HKBjfhYuMwHoTI4DUnDrKjU1MMkXrC/U4N3dw22LfEF8u9967jGrryn2YJrDQXbqSIUMtbP1
jDahYj74NLLo9HGKwC9uezQAwnZ9UDQ4B+vA4kNECAVNn6hxwyoQNQvQlDZzte/95Tu/2IaFUKyu
XkabobRxPrD3/To4jjLfrOXWQ6ZA44FZYa+cnNhKy9dnhYEGmo4PCsvRcypB6kIJU5T/jrkSiLcO
76p3NdQh6SjOVgRZCzvPGQQht9/ePBweG5cAev8FvSPNCMlV321X/Qf9BqeCRNZ2jdrR+k3VWRhL
jeeJ1o5Q12fpV/dRJHVKuas3wxkXI/pQSvqTelYpjmpl9j0peJZibkKx3potG3P/14z++rFyc8rC
pK2b4++xd5y28Pf1haFMViFHNlTrsmtSe+vblhkigglp8cWDLUZytE636EQjHm5sIAEfIh95+dll
p3N/ABUtmOhDpjUsFmExpCNpvNCXhgxDGm/YGAxF+a0mP4Zum92px3/Wx2/38paOIPBAf7+nZU7E
sPN3sm0q5d/8BnujYHZX2Dn1C543VQjqI9AnmsimRMvxBlUxHMuSAg3qUGAtxkfS+IdNNNzlr84m
KiZU2IJcWF+3JiQh/e/GdR7X4JOmCqIZ621ihHlyudeJH8vdP5Nhf4u9o2JTOrPeXuEzcz5O3Vpk
yH/xcOOPPkKT0iitC03NUuFTPYEc71lJ5AItktap++2uLpN034bI2Wd+qFCeIcA7qPkoSuydmT0k
/Xkwk5//F+z+WwNKQ6lAxIA1rXIoaYGa+osGu/E4PTSM0eG8NiMo/1FG4yNeqifDiI/kYaWRfdEx
fRw4rEC3n3BAa79+QT3nKJWSzxiKNMI8ewmlT3kHwQAd9IbF/xKRnFrjA8q92X8VHK4zW6gWAnhW
ga8YPkojr+Vqh+MwnENRtEghpSIuYBRybb4wmREro/ZfalIDG5we1tyHjD+44S6GICgUzSK/EUbI
o+r0xjn56OgNUh9I9jVF6AvOpo0HtKUl9iIQDhXr4o0RXUYeHp/fC+y/VGz58ZCVSaO8PnYg7qpL
jbb6eXmQ/LYS0Lzw9cHoPwASrZ6rHioaufo/gL3ZXXqijODyPQAyczPanIQbev1VmQt6aziJI1QB
VmVJ6b7dWlttcgEQUE7nPeSzl3zvn5P1Bv0Tw/G4oPnp/wOcv+C+0/0ly4YBn+pkG33zoJtdC06O
xiO0iTogPOwdL2tH4nOvmGGBmnrZcbpY6oI59eNq5PpFv7lpLC81P6d9xoL2mJkGVng/0e0pk6Bf
/WqXqP/XVZZO5Cjl4wDzvGKuEepJwTwYtTLZv2l4YgQ4+hO8UU0SXeNqmRd2rxBCbA5Ku4kLEKnm
+ycjLEgMcz/d/w1B48wHfeGcwMRhhwyNlPgzTeB98zAKiK2awQShCD3K7sPWW/WV7iKeaN0G3Ykn
ZNPk63KI2E+Ei1sLdwSFY79lat410xikQ3LsGbrqKnlVYqxaXu3Ge1mN1lqhc/T6cQCMqiCOmE+K
MQPoui61dOTjIFP6bfladYpdDHH6HshQbMdY/NcfV6PEYFONYgm28Y351w8ws7d4qe8P8SOF8m35
4jfuthTZAy42jDLGxpSdnz79nHN/oJpy0CiVmO/95W6EvVZfl3oIlIDOWdHoGFNxQ4St+iyWUcf6
fonz8zQOyHavuC02sp5HsCHJvxj/vwaVD4gkU7PND6VjF6aq4Tv+w/BTGMVxZnR0odvUUznnzEEd
yowBAM/9zUF1p9xgHS7bvBdPtdnZEZm25oJ/XiIO/Sp6gvo1y+usA5b6GeJ/VFRp31Ea/GMn5wgV
U7fsYFLQigosSBcRf1GFzMkI9RiU3kAZATBxb9f5cG9jTbKF9KyGx4X+28G/PdgRd4D3BTVTCRGe
EghlCU01nwEjhUPjuCUaKtv9hN7B2moliO1Q2nP944ucSyDZDGmaFbMPFRzS9mRKc8ucq4wG27va
0a4um5fYSZSgRvT8rcfuR5TOSluWTXRpvf1Cl4/8KGgFSBpDNq5R+NN2llFMenWzWDiGSfX7Vq6H
EbFmdBNCZUrbHm2KgjhO1a2yo5L+nQxl6wSKh4R/50Ngrtx0Tpa20DqIH6jS6slDF8fVA9/AKzC9
5pdadASlr7NI0XZCvT/C2E8ntk2hgu847zQl2Z5Lr6fbtKhu6/GXXV7kP76OtcxWNoumKZD1IjVM
a4JTYc7p0WRsC14CSbrbpHkx7jZYQLfTjovIBu3aMHa6l8wiCXyEZdV9l/YkCwaISPdcvtoDr3VG
zm92i+rgkvBxbX84SbJ4lk04LKkKg9y7OIbWuLMIxxR0tPL4h0X693RQM2KPvUKunRJwD1H5BmGH
VxZXvM6mx78UmmgYGdwg+UMUzRB7p5vcb61PD4VxzMvqkBRJkdBbnXcZ6NcU8xLSEfaSGySGRjvt
3UUZ+SN11CWbhYfFWEfaT3rgGZzxdUUSZ4UP/9+I98HGAIDePJ4yMzEkDFctecuVJXjd93DRDk6N
N8D9B/ndlnj+KnhmoX6UkK506mJkPpuC/7X9FNJH2BzoVGchpYtAJu/TQOA80Ct6FHXAxD4dHZwK
hH+VacrYgGg+1qgcqRPA+34X0FwOLlbC9dV4pnl7O92ZzncujaJuxJPLrb0y3Yfwnv+bSnerLRml
YsHjpsgFWgL2GTuqH3TFycJxre+vVNNSBWIkZ600mhpR08YRvwMMULuIf37TFRrSObNtc0tS6rmT
02huzIc3PbJWtj05nqvFyB9+6VgqAF/eD96kKSQpCHrz8MaYA62wSB5WRifzhitcxudstVmm9iap
YbAhDE1TfjRP5YwU34W54erjKHGoqXFfVrJpen6PvypUwrX1DQcuKYXks0IXNGq0bqi1vFZmpfNY
fl5VHtt9Qdc8QoFDyNWEXFc3ntkBa5a0apxV3YqdColi1/u/1SIeRAoS+ncmEdg/qtg5/Ql8+9dK
/N4REm0Zqzg9TpcK7UwHWArABRmLMjxhkYo/RhnECC1rGd9vC5IDO5w1IbOvI1fOJX6oKHuY6FYD
RDm/yb6zLLWy/hlRQ/U46/i35VAYOg1r3rLwh2L8KQ8tiGxzMI/cKlf5BFBaaP/jOusZ/1YU9oPk
UyRUQd6I5zsyKdjp41h2qcZFTnTclevtfNPl9WxLEJFXYTiICuBHTOspdXHACKTNCUCMoyVdjd/h
i7Qe4Rmw5nIaKMLDmPi0JW1xn9EfgYp3OKy7aRvJYjaXzE57pkJFqJykEmqKfdqlRb60ll3oE432
Af+4sINNll1qAgcMoRdBVnEKnPyE/J+YuWNRz2zLN2xuRclzAr+j9plBQzr75cVM8T8Td0Ck3Dg2
0wQqd9CnN3NSEUcNZmifaW3soAS7v1++WeoRqKIYpoABVHArN0DqTtvZqiQHQBO44Sq71r6SJrJG
Oa75C7wuKFrzJ4vz/G8BlNlBsUPU63IxZX5YknBm7pZOsYvtnObK8zUlqRWBKSG5vTycvA+LSWb5
UgKGLkohk3O8Ir/UeZQdoch0LqrN2jP/wWUkikmmqr39LJLZLwZtsaB0lQVtN+vcndghSp/uHqMW
cnzgbztKHGe40ckrkOJxwFTW62VexMRRGo5L/EU4TYu4yAhMzuR2gpERPZEPAj2jZhtnhiFqG4g7
fo+T1anOws8ow0oBneI5Q/pS4Unw80f5YFjtR7Mh3wzLZbYkH4mz9JzcOyME9r1haKIeeo7ZqIL8
/80SbeFnnQWR+mOIAbMGceF7UdCr4V8qNdpgHQar+Mmd7gN7LJWu4nZ0yq0Y9AuefzuXnDy2uX+s
YmzX8GyASpQFuvSkDM+OF4SwSUgERHR36M3scUZuS38UMt0qvclrDe1nkBTltJOnv/M/ErmZm7lt
NF/HTuM1JuA97Sghkmw8KNP5JLctVoSjlb4dTaIE43BeU3CtgX0XOgZNeWD57YlOy4VCfg/Q6fTv
P/sf716Hv/FTyod3il/HbYgjmz/f0Jte6moIdpcPladNPEHGHyqzOG70rdDBTp4U+ZsO/rrfuLND
9/0RREPEwlhzLn3y1gOr3S/wc66PGEnZ5dGlWqrt0vbAB2XcR01TpecCFCyOl8n0q9Ax9LbR7dso
UVCfjA37pP5ZFpZO/fPHHzg2DPn/QlwuCUxVeslZjHMeCgQnCeYlHhFiHDLvYq1O5sEBP6BKJn99
/sz7piiG/6bIRbTnQvPWs1GUvXMls+4v6qSpcPzXsNJkqC7ZKWVIWcgCcOfoxCybPrl3FgQGyOlX
AW6a6PcNHMxCPunMLhwES1V2UNvx1qqi+WsWxRpIE7/ky2BXuYZLjNlmH/ANtCapoGkrDhcb+7ts
xQVDsGCFofGV3MbApP+zR0ZOwZZV5lx+YfmCX+VNgS5h/gpA7iE9UHG2jcaDMj9JP2gHCXDTnDux
CrYivH+KuROQ1I1L95Ja0wG1bvyaBJzqJ3LTclc2gFaWxsBf9SSiuV2sXhDaOt7LyEGtQZbRE8hM
+8VbkZvnBp7+WddrtKaQCLXLuFGPH96dZGaUayYK2AeefQ0b+uD33ISU0PI9LJhFKQyNu/LZNT+G
kEXRp15hGiZDQ2fJCRIZBEpo5fK/bdFcTmjgNNvuldu4ZqTsVXUZDiNLzaWX+zvvjy1+smSKCwo0
7KaTzfoiLoVfLR+/EA8tgfIGVdgEQPReBvHRVwYw58La09fXfWiLKNnW+douukKWpjdT40xDNnPH
U6ISWx0vMiRZlIzyrDdlyZ0Su9E/g7PZ3eSzpjPAhcG7MrbZOivW9xR14AfvMi1/cx3+n3TYwiIX
rJGYDSRB/Q3u+OKl/QQmdiFAJiuzjwfiH/KHfYqyRdOOlUMDbgiQdPelOMNReib5KzBCzsAKRLuq
ltncrB5sLvu3utHpiNqjFZyQn3jPEjsrWG360fbqAXBtkXWPQv4kQLnGiKddpcLas0I8lKgdJ57B
Ft6at0EjXpOK+le3MnOhUHflh1AyNwcD0SF1beB58Tj6wuFnXpZp7K4eqTSxfLanACx1Z9loFGQC
E8wgXW/Ou4wmsQOOLhhi83VKODX2HZyqJP6E1ONZIEYGOrc6RqaII1b2n1ny1cT2Xl71vtqkrsus
XjxcFIop3rXxD4TSUEG66J3n7Ud9/QA82D8Gt1+DOz0AhCiNO/ntGzk8yinchkPy9iPWWijjdijz
ogNUygp8JLen83ghSRiSlGPUHl8lopb0rDkrgntn7EyrngYWyii4gIAp9bVBY0Ub6eYCkhKM1pS5
UBimImbG6z4WmVvqwIIETLVIUJK8/bdda0WGoXTJori1ur6O4kJta2ZO7yU5PMNlK61qI8Em5Ikv
2xHZW1Q6op8svCm6tidC/+KHv4asQyWuj0QYriA36QlmKxLkAz3tn7aMKZvFWQYiJSPlf4oRNIip
d/HqjNGCFBr4IGhSOgUf64mGXvfCErEzOk7nQUN7iAtpbCJ8/ulmjT5HUVKePwW3KUx5YebvgBmA
Z22nytYATy0w2pNcW+JOZLiwfUNMmhmnivvR3X6+eKLvRGo25z7d0OhxtQ1LgwaWFCryKZq647eN
INCJ6nMwWAvUk2iB3OxKzibK+jiaRFZuefgl5J/4Ts592ZHSRCOjBZXcEvIVBn04IDcyJnmtF/AZ
8HAQ1wh2cuqwsZzzKkzVjilOPT6KOCns7J/arrlDpgo4yvQNDIhj7VLzGcUKcf9sybMoFZZSjJRl
ajXthB1fVqsPdIzfaulZiXbolZTIw0bmxMBf//TnsUjjF+6uLyizI7AL12OKSB1gj5DQXdjWPZNj
gljVLWFmVrxvb04HuPQUlrCziLs6Zo8pLLWD3Ol22Pbr4xmMDlqRef3ALP94fq0kLkk7+jh1IN+2
zik7oXTMG8FTsBKufLcnm/qgE8mJW6PJZhRcXmIA4CTTYa5r6Em/U3HRcUcwqC+3W/eexNUKaLy0
Dv8n/HAD1UT77kuovQDuH6SQQzDlNNni1wywZMamvIi5UZU1uqQR2DHSCzN9yRMRjF+31aHW1C+4
hqdpbfzqwlbp9b9+mx4Jym6sMdXiN3dtf3CT9qzPxV3kABa38p0tkwClwW8Z/wEW3dvR/GNrBETD
16gSk6hUmHB5R5SP5AuA5hQoncYJeNNqPSt4vSPB40rWgOzQ4U8Gvcw9RqWTzLa/6rMjlMGb3tOz
+YFXvMruG9KcODVnnUeSLUFk/0gatJe9CHlBOfYiiLdmNJKuEM1zOVExH6NxIHEJ2K64VJb0NdRm
xzPx9cSXCTp0c8v6YQDkOHx2HUcjhPiwgj5vGxxaoa/HjrDejzv57no/Jli5b/2HethlQv2saMLL
3UQE1J6uSU75h3+FuaKsGrJLKDU4Vp7HWuyoZ8LTYISfoTF8e6Yeb9RvtRAV70yItGCwW14FnBdP
RCBhYOg0AwytXyQ6N3zp2pzQ9Ve9Ktu9VzlVx3e+kqqKfj2d0v0ZuTJd6/TfCG40jWYKz3SMaq9m
4y347E1FQpDD0d/T2qY9mtIqxVrPU6aauNbl9Ai5rXBYiXTKcS282wWOGcvOoYlsr1H1GwYFJVEd
yMm0v7Xwxwv+Fk4Mv7yoeyxGgn4TkgKca2F+4AYiUqa7/2MgDaCjTFGdpIpIOu4HOpX400I8ojHK
OQj0ver6C0W9YPLETxVZCrhdkMCjrA7s2o7verecjjF9Fprsn/MvpWjvI089orR8BtYZpM0YT5k9
Zu+TLsY8gz+/JwhCXI8uLs0isipfU+JX2eUr2+6NdfnqyEOiBebJpMi/u33WxOer0hPwwnR/VoLN
o22jkaJZqym5dlt1iHvKTNzYTYtdBzi9RGNC9iMYSl1h4Y0WpeD9w0kV0VjgT/nEXNc0QrG7qup/
qBaPVx77ijuH/I0zMEKxso/TXPnlP0ICTecibhYO6RsjybTyIqB+pcvTFIqZ5dCaUETok+QZU1Z4
HtDqQSCP5IQo4qjHkQeWFzKPBe+cJPiuPZeBLcDDQoZbygFbC0G8f4VxubHck08frnPxDI4jYKmb
iTZePT4RQt9uxdir+CVNhVqFJWI2vhJY/4trDkenbyC5lok2XRp0ri/Q+V6tqFtHMOmb43Hyd/1u
gD/lQ8oX7XC/mY9Z18r5SABbJ/4X/FukS7EdPAr85iZbJGSDPsea/VIdYa9ZsQ3J4Y3HwmjjssqR
HMgfC/d8kF7TK+i5Tb+cfSczphoKQ9Aoi9riAaTLOMtnkzwxz6zIP9wPL9pk9GLTqTS+8/PdNdQR
Efkjh4knsVEooKXJy9TrCdWJHoWyQ4OWNJPD4r6+sYse9UC+3Rse4JgyOp/k3irkgV3AZmul9K9s
kn5TgxD7B4cC+dT/+L5X/r8gtzlbOi0tX+wgjJY+BSyKuKH9F09e2XlzTcUe2PdCpEP4INOjAHsH
cSA2v2IsXpCO+uI8tMQowtWY2+ZoBGxEqUgb4CH3l+9o+B8c1BXIMjOT1WzwQO6CPPMMOYMUcKEx
FDI+MeC26k70fXU6+KYCW3L5xi0yksm4FOX0GTCt9X5dVXgBSOeor8NITk/5GLadd+VnfrESfG9v
Qe7E66iJZkwXLxK0lOJ0OJdPQOWfuGdJmf8ZcTTuN8hE5SOtuksRd06ZfiuMt+aYJ0cXLp+SfXU+
lQcnFPFvyBZGXFFIkRxY8KdhioVIDcmSUOv9XJXP7c1lrz808dYgTG0K+KQ5FdIc7W7Fee3ZvLsE
XpLQOMNKg1+atlk7/khlIcLeDMRc1fX5coK9gsf5i7y8sHt2avtpn0/9nrbWREwKP/a7UvkUprpP
6rdJL02G/8iDPzscZFNrNQ9VBKjng9UR3zIKoeWXJRnI3J9eVmGOKybqJCEBQnKxzNIFw/+gEsYD
1rzdGplZgC+2aWVvfRwS43CoJOAbAslxCCzl/p3XFqyRmu3+Gg5KoVXCRxaKisBJsdJ7wsJmcqlK
JCNASkkSzqXggVO/gVyo5822Y2sjHCtCp0l5obe1Pvuzu6OP3J1TJjRckgE3g5adgO+MbdFMM0OX
ME4GXRlhEjUX6UYmNIpSdBgTaY0LMe4tmmnojMo/SYC1/AW78I2BRgUyEp8XQZ7wYnEXZPaHVLef
9FBA3GXQy/eaOI3XnLAYqksEKWGLvsaBUtpqfqxSOFVYTS7nMMxPC53xPrHYgOgDGqH2Y88NdAdS
Y0I+QTZAfANH8OkaJpcYxuDGCpXbYg/gxqk4cOAR4zQLC8ac2N/WHLMaRgHyvD0oN//MyaoDKN4g
YJeeoafk7wsUzoYbBHeV9kDmaVSgoNPs9XZBH15cvwp4Mt8VISFVJR76oNu6W5pSCrSYb/R0WZ0t
05HMQkxzS6ntJ3VdVhUUqoo26ibXzlOgrdpcq0HkFizY9X7PMPY0hZV3kgrJ1Y7D8kgAoHwKeFvp
wLKzxYTttyiB9auQzql654cEBrpVNhme5dMpmI6gfKb6izCUAdxp2RoWjXTwI3ONZDDILKZyiVdm
VoVDI88sjScokzQsM2HiRtusFZjdCUFSCV6N4peJI2WGFmRhT7hIV9smCEVVe6C+/Fwss1JCqhpY
bgsTGi6LQyuuB82HHUan5QdlRCz0OXZU1y+jHXDqfkFL482QRgQgsfNCyex4JyZl5ibdPcnX1xUw
JcS/91DRYiikHyMuWJ9E1WFvZ+76fsQTs3p28GxwT4y4JvWagwxcDsPEDcCtmIEkggv/IcepE+ec
NkYkIqHN91gC05jfxPHEaQyIlZ7f08iH3G0sZHhM+ygEsKpO4dhV9MhrLt5Hre/lahsMMRcCjY5m
4sZZfYxvTkYQYTVyfoJJWrhyJfAG2OYOIFE8EK5if3wEfUbN8qTLRn6d4rPJacc3xJXwES//UfF5
Xn+9phRT4h6e1G1+TTIEQ32k2sOpNw/sAvFArOnT4H7hn4cUNNkHfRdNv/o1zsFypPzQbkUCWsfJ
4wYCRSw8lbMNIWVXN0ku2AgG0GqX8kQZPMTnZt8lV348upvOqG7oRblLMdL34V1lPWUjXco9hYog
VGEqIkZoLatWaQ2ThOfqyj44vX4D43pwJ5h+ay5EIMLpo6UWeso9pOQfc/T6vOZCKbDUUX+oHAch
lL2jVhzv03eyBReoGwSYkXNI1Cd87ecQP/mhZ2ALYLvp60ueFW7CACuRoFh4etUzpLOPH18rtr/F
0FLizhGWQv+nEvxNZBP6ox6hpYaxhNsxUJK18VdIWO7xYKnrjlGurW9uvU2UOenEmGK2WzpINLFv
WqtAtbd4o3bce8+6tMZRh96akb1gFH2AW7YYhnXGQRF7zeHZVkE06FaLU2pV/Bn9xlF+ONGSVFYw
DPmCTdQq3+EntzfSZzF4DQgfiZiZ+AWyOMHx5f0l+ScKYl1Pg9W2Fw98xzucNtHgf8S4zf3BRc1F
hPZJmPR/O1FWXAsM5JOgVFXbQq9iEWO9UGlmtNS1DZrhpTvDokI+T3sKtuGy5VoQALB6h6DOe/1c
/EGNv3JUg03KWnHwaYH6QfbZPRiewtjpKUmiDu57dmfsEmjH1MtTKe9bz7PTISIEmZ4r8JwsP0pi
CZ2ywZorM5WqyaftVQ+JFkNpjqUY9UDZdRewBjXYxWBorMzwlYqZtkBtGCefPK5EbSD/N3b+Q8b7
N/AWYYJ+ScAx9DPnSCtWxnWgObvogt5TbFXm89FBDYTv35bM180FmwXjJIfd2vT9JMKVLtMdm9PO
IKBqInhE6vMU4trrvk34YS8rHeRZ2QQG/y0f9wEr1W5fWmJHehOFvbgDNidjCDmrP48DGof7llXn
52v7rKvZmWrDaB86IDjLFFtD8UOmtdczEop9445iFi4mO+03tlwLY4Q7nLPugKjU7KA62WH4VFfl
DBEslwMpq9b448COqC7++F4ZukgTZX8EgPMabniKi6Un/8b2uQ9rUl3afItqkniwBeCWzKaKSY+h
AQtirvzgfJ5p8eBd2lze/O1dNQs3cnvMEiW8cFeyFexykFxoeVBf2Hc21ab2jgUtW9fJPmNsDLj+
tIoOy7HHfZejYfDKJCKE0gO3SLWQQH1U8AbvWTUiYXyPhO4IgNxx5Ret1KcY6ReSTv9m7AdgN/M5
6vy9BTmv0TXTrTKAi1nZwXFf7BJfMlP7wUGQzcwFAz+knjQJuttmbwljvmQRu40BjfMkEtvp7oB+
+6VXaA70GY5k73PHUnBrb7h21Pu8ZfJGMDcn5Zi9zJ8XO5c7q2Y0dL06palKCQhOC3w2sVJQlfeF
PpfOBEPc14zBiItY9iRweGKzy6CmKqRM6MVHPdr+GBPjXi2cz+Oz9iKb9jqB3QIOw+YX+jf0S4AS
+7S4gkXLs6WXKDoHpmHzWLYXjjFTh4OfxVBMePHzE9vHqbll0TnyFFT50+ETYvcGXIIXlMJPfkr3
aeLKYuMRy7z/OIYnMx3wJ3RsPb6fegRlV8w0Ezrem6eQMGliQPnLVaYhPFrFf+C0HemhMxfFnJNV
2CVhB1ex1jVltQUrUHWFIFHm15XXca+EUnYGyP8E9ICJxI1VEiAskF0GJBjSQ+Y4GlGzWknGglhl
FgzqPZP+pLTOE4qK4dZd741Etu8GHNy8SJxAoJMqQRUn0OnBfcy/bykQwcpfLKP8OJ+ahlqxQu4q
jStxAHpOXefalbDszaUlxiWqK1+PHVlJA/bfZErJ5zcj46ItMCLDg4zAq7jtIoRMtBaz3YuOPPqV
C9nnoxejPL2s6QqsjJFLrQ+nO5iO4/JjPykJ8Q6KFXGrmIvdY0nQKI8BOXUT5B4HyKmLIGn612JX
GI+LnYglqzYKwAMqV55fM2hHhh34qRIuC5PPhv4+Uwgcx4RKKPyLiJCRJ0xKDxySbwuZZ8dno1P9
UlRjvEUxkywaS1+ikpvulBEtFHPLAvT+e6L/lG7D6JMrSPw4nUAQ3vY6w86sHqYTr3SvvtFJUTf/
fv2bbi4ZIqzvUb/LBSU9v8f6eP5/rNK/s3fG/9zi0hY0Zu0TptxckRI0rlhH6NlozOMMVkQAIFa0
a8Ib9hs/pA9wIH+jNNY/HO1UDin6RZnEYVFc5FPsD2xgHZp5s4vP/yiYMrAx+vQgvFEJNpCtgTtG
ZFV4PMCYJDjafwrz2EKJCmYsvWMD2cTavUzIqR4KfPxrn+gNPeZipluMWe7b4WizByd1H6sZtYHI
RZb3hk+rT6MWbmg3dwejMOBK5pwm9NtTvs8mhOd9FcrKMFPffWucaUsNp8nKDVCfYqFxkSr3MfaF
nn4EJOOUBKuFVdBbSxQ1Xz3GTIhI8e2HX8gJTVYa6TzfSbBrRcLQ64Ss6IJdxEAANjrVAQU3H5OO
NWW3V6h5iHO+WUp0m/Ny8bGqQaQtD4wmuDT01WXKRFmmpamOU2EzQFTB/gbX/l/6D7klvLazsLhh
ZGMPBLKR4Yuko4ise2jhgpVrN4sc9knwExL7/iHMsSYUDxjrDU9SQaKLUqOFNYz2JOTy4VbY0U5x
hIYgm+94lNCfADXyXTKGA+7lV9fCavADyRmxGaAyEF+p/kAP1rjqDjezwWJ/Tc+bZ5CAmEtl6p6m
1ZCMBNSNEvsSanB13tayJ6hifoFf9VT4LiAKUU7eIZWgahQKqOL9mUaZocRbJbUwpTJj+h8+F7RY
BHibBvVj+yhRFYLs4lWJ38A5+4cg11YC71uWKHWLgsgz15+L9JmYF86ETN6VxpkOKAgd6elgwh+8
WTgh9/U5vWYtefBKjOE1j9Y5pSiLGSpu+k94wpZYNv8rF09qGaaw+KbqzouU0/eOEGtalYewpfCg
J436AD/sbvfuykWH3znXlz8hPuDPBOe8cUxDVmQ8SNCVJLfm5ovqRLs9nNpWtZwQeP4BgqDmSEM/
UyeoOQDJM7BYMFCIxMb8ccIoyBQMwVS51Kv03ZzQx8f9XyHCLIJ7TM+YgFVAj+8C07vuZQfRo03G
nlTIDDoDh1T/7yecK3OmlEi10vBt5XX6dRq3o0+Rdh23yksN3hms4ujKhcZ7eOBSLNuyG+cZuHB1
PCD7KUiGfbtNbf2/LXyJ3CLW7jKWGgARpKgif08mVJgrjWNWsGlHIfe231J19C/PqVqQKzDKGhYn
IK33YNeowB+NLhAs+qK1uIGh6lkY9uxJ26doWYRFF6c8kU/MMEY6H6yexd+UENpgg3UYMOWF4U2h
aCWBtIPxvD0okS2WgRZfGp22fwYg2UZ0A3JrIRaRgPvWO2jXFAWZlT7e8p7rTmRfC2xi9FPK6dJR
3bJaS4IO8uy9/fts2NqdZxY42Ppp70OHkmHbaEDHVcNgZ4vpW+gBUi9GZf556xV1LwWMtfAJGgN1
PL1RUFaytlVLI+ShcNH07ulvMS/1TSdcJg+wW+t0OMz09JfbTH83j2xae72fatPwwm1GRVE/xWu+
NbgK/5h+u9O5fsRvPVHqviHwJl5xatBr+mkvm1ITJL9Bz0BGY6g/DY4Mh00M6fjMpJxgDu5JRRho
6yjna00Hb3dMMnrCIP2kDv+io2CEfW+5fnKbukyyCkK5mITClSOA++6oYVC96YkIJ4O7qbW+avkV
46LxC46ra6yFmQaVP1A1N4TB0zMpjxwAZY36rpoZJgwWofxeR9o2XAB+N+Y5beQUp0MZ8/T0M/bf
AAgPMIZFcknyNuW+bZjsbWI6Hrvppwwab3cEDEv5ujCkmyRWcDk3fM6X05C9JgbRiY8LMwGJL+mk
rEtu4Nd99VXOVGIXE7F97jxvFZJtZ4ir0sDPN+DwHKWIOv9qL9ImRzIP6xDWiBMO8taSofR12Vs3
8zeIFRTfYeNOzFSqtmpWpF9xl7U87FhhGTqUiUjQPuza3rrOuqUqsMjjVV0KayatFgJ61rqozpWW
SjchbPQWuVVbkYdvzL6pXTgseBJ5skMZVEFpPNVP01PGQHvfeQBvBHV4q7XVOEoLvDRAl0Kg1Bg4
Tl4SSIhAMfu9fOd0+DGgstgw8tHfWhh8EC18SrelhKTKXlCSmKh000VpHovq06RORK3TFHRsVWz5
eyVra9EzKbH+1DJZQU0H3YnaB3PTUVPfPuqGAVvp4aOJjxSPdlXbW/P77dSa+LjJIhDCcZZpZ1Ub
l8XXeEayjmq6ufhQ9fK5b6V6YMx05RNSC9+UmnY1M+C7wioty77ZTFng8XeNFgxqSyQm6Gmq/4XH
mTECxB+1EGP3Q9sMKkWJ4WzF9SRRaxwkGWXUpj9rNbv+6VJjHTjjjSZPO9ERhdyd5R8agZbZaQAL
48lSAWeZ/aKHzYYF1Z4Qx41AKkJfxaYrAJWHIFcsfA4haMqSXwH+aGmX3NoNGXAKYf74KLBXxbLF
VwXOWQFBBVdL3vFmDvOImH5YqVL7FJabuvQtdDax48n9SNgJUrhGPbjDaLbD19ijUApCwCuj/qel
15Cqn0tOkv0XIv0EQlPx61rtpZhj2AJUwdPzp54RANGe55dTzOCHlVbVyqePWDutqEEb8DHfOoFa
N0avOM36e4YCMCzX/bzzzSD1nwvdyXOMwobMCRbt+KUdYN7V8YwIG3AqXFuffOdC5mmB7rU7lEl2
oTlItBYWiTVah+Tk4WUtbRPOrqSxaF+IUZhZrbEkeMW85CF+5ZloJ/7dfPPIl+haesA1Z8RcnMlX
H1VBlqViAWgC7U/1s4V26041JlV65nP6rS33SA09Ny6at283JdhJWYRfdy15y9oAFbHnBDKgZ5yf
Iv2UkfX9a14dg9wNhkE7k7fqIM5vmVVeyaZiP01P8J/w6qeEIfiYvA+4d0bNzn8YlfsmNKidXNbb
Jfj0EKixN5x2n5GwHzR9pkqAyc+Fm1L3S2bdJutix/DQl4VElYQevxep2Q7vL1i+AcmYzWBlhliV
nnzihSWTQljQ2so7q3P6LIaeQJAnpMqJ8xaOGdnDQq+TpgbewmfC4s0LX7giAHlXStizMu/Twspg
zAeFz4GuUuP+t4A8krtj6+yPF4FfTFwPNd5qLPZAJp5vrRPa9/i4OcG+nx0T82H9Yfygl3jXar7v
ppcrqkUdfQQiLDIflEToS3sfHvNKrMGJH7KeNnGL2puzLwaAES1jT//YV2vN14QdxdVAJF+SjeDD
m+obioJ3AP7ntlfsY3NSDxrb1xC2EC0m9bjTbqBRg4GLPc91TiPmNdlYKCdj8OJ+iaxYO4yVdi4B
nIWytSyUmVV4dmYXBZZzPi85BHjkcA+AcC77FYQyHUXmTSgjNR/tx3e8Ym6hCMUy02nePj6N799a
Hn0cHWnot2wpYT65KSLqTtTr/ulI+tfnoyenc/eUE44uFTTsoP7WYdTbFNN2jNuBp+qoXZizcJUB
gvz5h8b6d61AORuDcCS8B2FMDdUATR8BLMPzePtLP8ZZ1sH6OOT/gmNHGD7Wl7eIf74xtJDCWiKo
NXCJeV59hRIwioC+3PwQnJi+aEpL8s2/Gh9EQQ3xYLI53QQucRS12L1u6OzYd9TzfH4dHgU7CWWQ
/QCF5AwKHV0QSvI7lh9GsaI/VPIf6xxLUhFc1TO5j8BDVR9tyqDYVui4Tq9nJVTZiUUYNsUPtMhf
rxQ2FCNSuec5rPMHXwVQ7ReXdr98+6Y95RWdXqZCugGW+1ldNMf1GheHEfopnnEBv3ccN5P7lfRb
2CKv9tDQ2qpoyNG1klesjUUp7cq5kmP4OkoLpldSwnyrOb8pgwD5rSh3oxYNSH7MveWHFvOasbmr
AabhQPmPcKTpNQmd9AEIHNOICVcEFHt/bHG9i1LSDTFisOPyx1Ja10/ujkO4+YuwFNhSCKcgFZEF
vW5IE0IXeRq9EVa38tdmOyeZDUu37OJC6DPqsXmeQJAgsgF1/dnKMJOSZMdEj67KNLx3t6+0CQyK
K57SwiTAB5dvPyI/g1T1OTTzwcl/Tqzd1/qWEv/lsSNmxG+cK8kFuCfCI9167KOPQJNkJ68RkmNG
xc1AMwJHn3jl23eLtFpV57lGWmC0ZoyNLvvQ57YsyOsQG7gh9vCvXhLzQG7Ld/0lUwvTu8BwG5vp
TB0Dxz6vZ9KO+ezJBv5lsZKsAHrtRTiwbUFAKA0qF8MoZ3DxYl5PfdzFSOzGoPirSx2amHLuhRsa
HFUnHye0Xr3p+DAXc6ysh+2G9uwLZ2o23L1RVOoDXBsijN2EyoyHHpfZ3MqVb7GC7oQT4+EDZgm5
JDnCmiCwRScENWJyaEOoLoC+Jep6+I1VaLjRq2Dtk6My0uJiFmDjhQAbzj+yBU1H4CReVr6+W4du
YY8xTiKRmqNdA9O9f4Vx2HcaATW9Nd1hhazLLYM7Q11JhJ5FsUV9n8o1rzHssESnAdFFl5SDE1mg
nK8Pknwnqf3ch1LSxCgAWRsQHrn3Mb2c9uF1/bwCugkTjskz1neFqO447W2E+1h8fpEc5akbdZI0
nuE2kVGAYhcERdZrm+bRjjVk1Jcdy458uO+e80jO76ZyVTk9bVPKj3HtPGANw9gVz6yH+RJSNPcs
C70xoXZv9NhF8Js4XhdolftyqRlxp0pXyCoR8jlWvnFFn2YBFiWIMCtiGcawS+57iFK6XzSDYIDT
CWf/1duaDQ5Ijje8Gq17TnRNI9oGniOtRqxi6W4yLT0fgP9ob7v+XGx+8AyJIDwTJweGoS2miNHO
ZyADG4FKwGcJY1WcfVOnahhJ6Fa16egcClIVCRc1T3Te/E8jJURTqKCYDTUJcxExe5zNB9Lh3zH5
4izbPXKy3kmQWMIfcRZzcFPPatIbPCMC68eILZJRwE377Zf4OdXTvKPp5RRsWFC57moGkpSEFcVZ
tnV7wYRYQzre8q17GP+WKdg4DXuC5CpG8wMD6EbTuQqyX3AT6c4PtPEQRAYQeZHzK0h5XW+mKbBM
rWBgTbbyFDMPfGVCBomicU82Ng0MktCt9TB6bXe0EJBGz11zcLkzJorCCtXIroKAd4eisYxLyvPR
bnHBiubJD0npuH9pILGTA1qS0Qp4E+G/N7ev9e9snQkAJe+4QksbHr8O30F6TV2qSsaE0PCEjY+D
dzOyLPQiCIslxD1+hs3Vl4fkyUVHa6Oa8hgB0juyH7G/0GV5Tg3b+Y9H3zbN9KV4j8IjRGxSfnRO
UbpfNfUvbgMSpdKkPOgIJekD5PgTiLRbxMl1i+ZdpmtS6i+mYEEt2AmgJa9f980n2GqcpBEgQhsq
cPdgG1q+IClDjrJ0L7zckz3u3dHdkL3Jr0DfdfyDggtw70bK9TnHG4pdp19lv8w5d7n/ZC2gm6pu
nIdzUw9EPDDNSN7x5AT+xmOG462tfpjUDpgyV2fXrHBzRWcmo/sV+eTEnurD7BFK32m4Nz/RdmBx
ZKjb+Jkkt7QrT4pVesc4AUn/mmZt2lEeehcXCOZA24PNZq6D2h0QUoIFFkbwLcRKYYDV4AoV94Hh
nBJ9CX3SMgp1VV07gWA8G1K/4V0mNKX+CODd2DLWU9T1QxNL8FFSEV3fercZ0OwMC6UAQwi9KqQO
NkVq1NqP3q9I81+iU49Wy+vePxBWF0Q5/57NAtO3zSu0JPBiZOAZ34WsVmgq78y7Q6pB4c5tWKmI
TJJtQouYSxle6aM6L4Bh6e/5hToFGruvo2H2SUgvntrh/4HlJjh6KBKICLsuPXVJVgWdF8MLk1no
zpwgPWX8buEAJV/FOMLZP1ylVl2acHW5ZYB1uQsQ4HPanwMeqxR3elTGYfR/cA1ndH8OygtsGqB4
+QYvyN5FWLWpA2CtuaQroY3p/ujwjdHT+cVdBgHTl31qChZPzNNpyfIdqBG1tXJAHQmrbs0e6rwH
A1K8CzBO4PTd1PTqD597XEwMzvBZbzik1STsSQ1+piiFQRtP4icMtfp2wzXfrlc1UuCdZI6/WsGs
Zr05SVNBNqqem2aMylLZmOqsxGI/FbZjYbq3i/YNgBPrmXvN6SxqlagHPjOGqR0cFfG+qn/qtY0h
8oFgKCSqq/Xw48gSnmPKSaCoNNqf2oR2uZgs1rrYrqz5r+liVnrv7P/jQN8MLFdeEbEHbU2sCUM6
o9mxF4KuKTz16E6Aqwu3R1m5Fzn5iQzHGwQNr4b6mwIcLwc1qaZuve5RhXqfTAqzmQ0grHf48P0h
xUMFxYonANZIxKiiDaomYTUpX3MfRuwt1fBm6WeU94WUTy6ptlIxkWn+VDR9bfalhoiv5UhsL2T4
J/MOEJiQpI8QkliBx/hAa0YmM7MZCsf4dIQlb4xJSrnTa9RhvfmdqZcHV+WW3SfhxhebkZP0Iwr9
aI6+KV30ILIVE6kl2EXgugsa8W/iBiqyUg+YOs8KzL27kwbvaQY0R7RvOhh1H5fE/t3hqOSwkpyf
LUG7HQ5JhXlo9wz47ESvt8DsRrBLXsWCujin09c5pNHzF2KoHCJOZA+kyUCAMUn+Z3zkxHwZegIV
/Y68dKSy3RU4hwQYy/R40YD2ZQcIXgqmVR+3iJYY/ZJKQ7xZ/0VQ21KwLEFS7/wtIMHbs+A1eVK4
AGA2ROHfWftgTvvn90tApd9tcPzx1aoAd3Z25heBud3B/hpWuvjRALB/Yij9hvOJC1///VY5OwNa
9esuXnpRa/7UwvOLN2GkPkBgJu8igjXClEdpLPMSRT1WAf5OWxDTXKjwFrZhU5N0JtMqwHhMV9lf
kvHkMyHIzFned4p2a+4y+2MDuFFqYwmOk6sEsPME1f1U5rkt2wlv9feM/blz74XdK08HOP8DqMlo
lKJnfyQN15obKCHbVWJK/Pdb6g9dnmNdmRuz6qaN0CFeAIbmGOet4GEvf3zS3S9Zsr/N+RCp5dI7
qjoIKfrponzmGLdSTsJP5/kcJjnBt8q6ynTdlfYOwT4R3WmlcdX2Nnf8l8UlgoYX7gqs8oo5zEH3
ZpZVEbCGpiFHaAR/zPtk8jXaeuTbrfRkhV6UeG45NrdBPmr049wms712LjYbCOF6Y82IISKMRy4j
+hy2SW+FBULYaj0FVxKkuxVx57DEG4BL07LCO/6/yET/PjUbJ76SuBd9DrmnuYheh8aM/AwxTfo7
HOQYTEzZw9g1hoTHHPHyTtmjdseDM+svnh6LQPzwVAXQsbYV6iUzLrXcmHNhKgpUAOhskTiyUDv/
63tAiEo5k6T6gigeC31+VpC0p5vuJ7cZuW74NMEnqeE+iWyyhHS8JzNa53yRqxo4ckbWgOkcl5FI
gnKd4JohkeIkvQ/A361dyhYcK37WIbt/yEp1CGfIbgFdMXXjvTX1TZND6pHs53qGNzr2Fys5cHvH
2Rs7hq8Sep7o5IdPYM9yfFgr2k0LAUvx2FVZdMMOZYjRtvg5QYJyDruy2js0DBDwoQHDtPPgKjAA
Gbc3hgsd92PKYSBV50BIWYmhDRbEifSVNvlzlt59A7YajCmkXhbxNvKtE/5kUFV7f9S2aVBTssJi
MOfbx4Mab6IRJzIO1RIf1tS36+f+es2vvbYwSYniJsRVRVW0MBRzPh3ucLzVgAxJEhZDGAjvca0I
QHU3XIFdxWPOuAH6TuUmzy29gDsUI1p1vQ0UYI4SmIl70Yviz+DhRtDM4or1krLZLAlGJBWgSpvD
0ig/jOrtTBYA3gWWoGnyPofBzjJ5s4j5JsxjxweCp5uVLVmT79iYcBPaKcdOCTo31zGuorJnUaMi
rCTjDWV4j2w7CoNZlrnu6DFd3kDt/W1gqs3QYpf4laNPFIcBYBbNAtt7103X5ofHDTdPDm0MBFHV
NSJ7tPfqe666Tgev1FDAuGhp9plM2xBFJycSN4iq0J24hAN6ZIvlDCeoY7GqUajMMafWdoEBg5bB
sXs3nG2i+d7UlsftRNCJR0uoL+ujlWdijUY9t2c/CuH703wRNTdLNa5eZ8BnQTKR5c0HQ4Idz83j
htG/Eatxcc1q5Nu/Jo2atJS1bcLPsEkma8eypxfMC5YpHTtpooEG3jpMPFBgvAwMV2qWpFt1eYb+
Hqt/TuZKFIUff3cy6LWw5FUAAYYO0EwIxfzO4kXBcOlIngaqSwpWqAo9PgHgjhtbjvE9qClAMEe+
Cs42B0iEOKJB8bTnKsWsFPT6PSkCwjpbBgr70QCXMhGdoSiTwN1JTKf0yI6SsYEQk5R87vQYkJyW
cKRzesXtGq5G4hh7ctpnHxqXGuy+IdzCGZB2V9FoBnDsNgJK/7bxcF4Sr1Wq3xNEVPP5rDG+ad9p
wdzRifnQN9abB9BFVXJR/5Tj2dODmC8rTzyXPZ+MQA7ugt2NhxV9FgJ9DJsLme2rRZ0yrq9hG2mL
e6LM2o+4NVU4Tqkb1KI/Ieg3tCXjMWvzXdqlcbLJxNqis7yYz7pxRRq4T1oDEgoZ0IlROa4jthaH
3E4g644Nbq+2qJC4r/Z7mr36iMAWCUuGzNkSeEgPpsE+y++3wNgT0XkdsBKACgeKQqNpW7EXuvNv
5Y5foNj1Dwf9OjfD3DthNQtwDjAcvmQ3a6q8aFnpv7OUM151m5gH6t2+YJ4j74sjdp+09vrkkS8i
9JJq5sOnVBw+vYqpqoh70JMUmRxS1qHAzHV12dOiHuhyK7ZPVRlwXvXHR8GFSJo7NN6uQysNEwNn
Mevxxj21SHAnCBH7pgW01o6591Lir9w5l4l1Hy7iGvYb5lemt8LyYyNiFblMXRL6VFgYczKGGp9h
3nLOJ8EA9yYDgdM406i9MyWr/3XYx9PuEjyCY3xCLsCDzabgyIDimN7SYwfV1cHdovbQISJkvMiQ
ilRbJ+5F7+SYA4A9i+khX+mQyoZ+1AtJTxTnXoxF594s6qFnU30p/o6ovn4i7ON6eIGrYBb/oYiT
6HWtv0BuDJ5mNYVPVh0aD/chE+oU63EegJHCfGpnxGNTxwNXCXUTcAJYSmuu9a8e8FRVi8NGHVU+
4cepFpEaJALmxx+HfMXzBCqf9amnJdFGTwZ1Fs4T2in3If7OZDoBoOq0iNKvRO3lnh+uVPSzPwXC
nCJmbrVmtykGTFa/7BDyTfrr5hT+RVqYxY4DeXI9FTMxjyIEunfJ5urMI/ROYf8JQCskRi76jamI
p2yHEQEpjK8cvxqTvZ4noNrs/LzfV2T/UJEradRBAFB8xmOl0JrtsN/6bxgH8FVvGYeovdCe2ydv
CEhtNV7WgRBvZtAcoxMzCNU7Q3qbt9K74bmyEch7A5PT6c9oBAranJRNI10BlJQyF/xh8nAa8Snu
GzqR3TXTB1ig+0Q0Weo39kGi/eNB9S2tnxZWk/tOnYEyTOoXC+hntvFAWOGwhL5vUfkR1qXK5g06
X456pcGPQevTPnCbhitjFIk8LqNdERpb6Y0JTYbaK4D9mV2Qb4vy9dI/IlItl4/1d7Ipl3eefQQH
Ihu5JkaMRewSQLrvOWAuCyGY7tvi9SfuvUngV+rDt6c7/Px3k9XQ5QrsRpJMO2dxqH+TufiaH/7w
PocYJbAehSCSCvV8I9gxLufSeJdMxVa7fGCMP2yBgjHvj12Mc2CV4IYhNStWeSRAKdQp/N0++0D6
WSSpj4xNSx2X85ImwuW3qXsE3+BnBc4yrczumYo+tCC39WAggwhKBMTGn5BksodPA2KwPk91otJV
3L1taD5Re3NaWOjvMFYlqNN8Vos1KhMgifqVQHIWj0ivL/KPDuFIIWMPKcHrdhArf3Wu8uxMIMrs
rowIhNlBd0v+sdOp1ExXMy7nSOqtEH4bhl8ZFIAQSTglYPLaCy6LDcKSY07yMJq4IjqhHKOuLIWr
sBajt2PomnFWlLIh5EKUW5qwOfcJp6wfn+Nrg5s8pOxUjhQybCCbytrlPFDDRr2XNjrB1LKWDN6U
l4YRH+zTYVxFuISY5wqmor0f8GTT6HThX8DzkWtH/ePPc5gP/w1o56Z1JDIsMQ3BQ8tCeVALXgcZ
8ZZWLfcMx2TqXQg9G8afe3HIhiseb1wQinuojco94Z+Ymis6dbja2cp6VuNaV8Anzl4Y6ZGKEYNJ
/JkrXAR00OayGrdBwySjIJnO5qm3/BDRRIMHYUhgTIotqejMmOhifppT0e9ebL10k4ki5BxPZPs4
/Fdzs0wpZ8TU9jaGSuWRdrUGZYNxAlheBAZeH4WQVwqs8GF4u18slATETSQLL4vYg1o/TSqdctbA
aTSPcD4uqP2PILI/X/5YPGd6bCaN+B6LtJvSXVCKAjYqqo1N8fdHuEHqHXh+7RYXCcXm4xqe0voe
BOguGWXtDxFGzb9hJG1RQ1WgZsfip0KreU8ZEe6Uur9XPaqWZgYF4GiYQqs0XzwjErtUtBFaG+BK
ktSg8pDYc9eLoAQqPwszwvoroNj2of+WvuH+CCSGrUwX4iNsZcaUhRogkCQw9WFs5l1YUD5nmjxB
QxFuofJucwkT/gH+fkhEBw8568Af6I+1KD/+i7txnRbiBqDP5Ld8pWUWi3Q+0r0/dNuOrLZNc826
f5GK9gTXFyt4eEMvqYa33YK58mkP5ywaa60Hb/hXPx0Knw8NbVRkWsDKpqbZJ4biOXKW3eDpgAmA
iZ/o0/8oy18cGrIoUKtXc3IsjKexQabBhZzXyHsvRcUrFPjnyCiE9HW3zeJm1T0xbFDCEGBwd1MU
oiYxE0Gtj2ROcNiMmxA34ALpEzf6QYM2DdC/EpZBjlr/+Z8oe7UrW+CoIp4hzzwvC4J1wxWSA0ol
it0XAjTukLD3W4gD2VmyYvf5o3D9C5XIN40EiIhEaOzk3GFXlvFNSyGFTw/SdMBg0ZZViZaSPa+H
QBNHi0sPDl1JEfth99tEK/RQ6MPWk2HTC3MZPiE4/HQuWN/hV+NfJXuRPISG0wBwvUyxF+PsTH81
Oaton+n470m7yVS/Po3+H0bnRkLELwg4iq8ly0K+cIGvEyirP7AiGMxRYyKmGkFPoHzJ4njchuzJ
p8IKwvJs/bPcZzLmEmX1BqUnBfwjEMzr9v0KPFHNJjaVp9/e3h0AyuKVyj3QIrScCGoWDs9chxSK
snbwHg8RN2s7kzYt5gzARSkjJHrmEPJH55d4L5JiG8xEhelT7UWePvD3pMwaMR4DT/J/sQF2v51H
RvBcimbbCht6Prw4HGYQrvO7NI247XS8oPj+LfBUb3G8kX1d5jQ6sOt0j89rmjjrhiGaKZqOQ3PR
ldONn0n+hf+eKi5OgKz6rWsYqX1PSD0Zol30MlEt65G3AeCfv7YNyfYbLwuxm5RoUkL4Z92Jdlq4
PpDLhrLFqNb3mKgeVttK6o47nBpkjZJivx/pHO4f0Fzb7oSPJyy/kUDtsx+IpSWpRDdJhusoqU0+
CYuP1uslxylZHBPpoquJ04qJe5fe9tGI4U9QMoGHfJlsg8Qgy1f4c9MrGavlfOHz1J17jpobKICp
p8zgKT79HjzY2tGaGyqgedCkP934pyqi6askXwYL+BcdLzdkMyYJFVt6dtJClCVLdXhAQMeFiiIr
OrUqcM/48AymUzx+x+zmf2gLIVhkgXZHLvra9wgudoO6BIJZ8nbJ2LZyjyb69u/Ur86MaJcD/rMh
YOkGyO0eVRsbT2tZSwyvFto1xBvxL4BZPI0MYrAYs8re2EQ0iHnGKz6tLrqOvtxPcuUFnsMchWre
c0RQABCRlNLP7/zzBFeZRK4uhuGiSgjGdz3WkcOfT/W6f06B7JIGwqVtEEvX7SjzgMGPyXTnpyYO
1jyB7vgWCR645wzALLsKUzXG3tWxXLtVvEJfbOXZYwkVo3TgZcl1l5S12Pk8aCgJ2C2qP3qPJ4RO
pv43cI5QUxGozOmaUEgEXWwHZ6J1gKaMzMaUwLiP0z/2uI+ri++eEfpGoBmE6CgFcA9bsayonH0M
FggiG4UFuVc0Bm0tJ+EYVgg71kqSfJa0radBVe+T1vCaB70xwFpGsyycpEFbzyUzgFV5ErrN8V2+
BzBaANQ7fyWVMEIcfA9KuGpA0FuyL0jA7JslIC/xLTVa8LlSuQ1Zvh6nGdfWwpNMBLzeoIG7hdEh
XhuLPhoVhvedTdHMOXs2oGic7iZK8S8F2iGWghV1pStI/CtK4P1AVLoAJzAW5ZZXIVTFQbhxrW0B
uCc19TdqNsq/OPkE7CpdbDwESqSTjZfidYbiXAjBjAoRLkYbR1OT5bQTsGS7kURDNdatSsOGqcp9
V5VGchH5jS1CnoUPlxIp+uEfJm3XIiGIRVgkgiG4MHkE6NI0bcSGO0n2AliogY5XnhNI9YguLN7W
xxzpSSfBeMRcItGgP1iV5C0wp3hiibnih8pujjPx+Anu9RLopRzhn0lqKIecy6DuPLFStopcgM5N
9EB14vLVsaM5SymCYS9wlygzpschgjAkQ282m8TOjgLXtX81bFWx/oz3pnnaPqtf45TCzq2TeKOj
CI4K0eoyxOuEPFpLgDEz3P4JauSpaM0dwKe08/pjbiwkiS4bhkYi4gerezOObVDtLKsueWNE1jyb
eI27Rd8ASDRZr1yzhWPYyH5+nubLsfwhee5nxoeUh1hU6qxWpONQpIFRMilE9RP2o7VaCVBh6M9a
xDHdW4clO8NzZ/FXrWB8VM77h7CJIRDk9iAB/woOAr9A6vmQuFbk1ODEWTuQ3OoqDh4bPpIgC9Oh
//029O80abii4DaPwz6hk/itgGPRb1D2EhpaX+iZ5BY0GDn+cayRfHoJVXMiaXSCWNCg+FU8slhx
J6mndPNtapriu6/OJfzEn1H+ZK4gbxAfrgZD6Ji9jPY6U5dHVsF6ANcS/NQigYFfM+0MaZsgsEsl
9p5p8B6rTDZji+nSdYz8O0d2hmcYxXtEcl3Xp52ZyjANb5JuaQJy3xaURXuup7Q+VlSh8E+67hZ0
7R+nE0w3CHM7TVSrdbUPjzQpjrMuLdl/eytCryFSc+GaZRWKOFH+mw7YqSD5+9/qYz3MHXrtA8Px
4kIJcsVwGe+4ySvM1bXsKm8IXLh+8H6w0jyVBahSUrqnVz5i93qMGclfjdj9cGF4P5xKVgkq/rcv
PhhAtSJ9MwdZUn1gciFsmLsq/RUEGJIQi5hwBYTTKdlVXxPgqnFWwh9VzqjybQNO6hySOjW9CNq+
5cbLhBEcSiflsSVBeRuXgmpAcPwnuZo8KT9su4esayPwsJJTlBQetMWsW1j40qNQsPdtBhHXo4FK
xRyJxiX7AvGmvKBSqkxM8g5KM8AF95xoIQCq8LV6G9surhpCaylnCdedx9DDzjryC3xkSTDFfk5N
c7M5L47J4xDyK1nmE9tFOvNF3lqBKV//dwJ/9dJpJn+8ocdDr7hek8N6tJ0EriDxPGkpo4KJkVpf
YgDBXCKU70qdjJuMXFB4bx8Qq9R7zloaqdRJFXCxfVN9STwArThNIkS9kMzeV2VdrP5S3+XHMmf0
uy2GlOW+EG60sb+N5HPeFIOoUlr0Za+d0l0UTDCuIsvRiMxmWAgZXzMnjQBTaZbRtXesn5y/XxBu
c5Zjuj/Gy9KLEPT1eXGrVLg4ee9pdAcJKlgP6vIXTy9ElIB73edOguP+lfcN2RLcxrp3/b6Q8qAO
5gNrlyaiQ0A99QHMvn7gNdWykPEvRcxi+ZsBt6sFzr1p9+IZlpPT5o4QKESHjcDjMZFSzKJDE2DQ
Of8F4NfUU9w1CBVZogI1LNdr5VlKkYlDzr8GZkw/kMNHI8Z7MWx19j8QXx2aq/5V1ILMIOZQlWB7
7DqqG6+f3ggaLC6S0fKW1GcpRLW+BPrEIFjlYJdv/rHn3cF9PwBmc39rsdqb0anb2uFNEP4DQfLA
nUXY473sPn+OiKIDHcAh5UyWe24uEIkOS6jeZ3mcundqdt8Ulgqh2CLEMrx0TVXKuAleJmPeIYcf
Hxht1qt3TsA7xEthUCTJL0t0ou4Dga4nhvce2ZjLW1gr+pK8fmidSIaCfk51A9E8UemRBgEA4DkE
E0YEBawzQ1l+j/5yWKL4qFnPIguVf8qhcsEQC0qd8tnMOoHQtFyXhiFpv5l1ubvgNXVw/K9yv04p
2VjVmOAkip1Zk0uprkdvd/GuUQtzKZlnYq3HJykJqM3l3EG6GiGr5YM5qAn5znn/radyh18c2fSq
pOwN/D7Qpay4mz4nRUUuKx2MfQEjNGR84gFFw+HBq1E6MZo5IYx4bXrb40MTC5cmbNO1wuX0JvnN
xKbUm69RKJEcZ4eOOw7qA2j7YCaPozDxavwT3vOEXir1a5DYT8WZ4uqIUAh6yPP0pLoZUpDsa2M3
QpIy8rYVK7Tdnf6i8wNpoUOROh3Pwn5Jg7odgtkNjocN0c6NDyi3Z1tdEPLcUgXB5kmjes1iNAtZ
+Pz3M5VxpfUIUXvpeqcS6X3m6GhRnxsB066H6V3t66/5bK6IflLRvk3mHwgzvH8axJa8mQQQT4z1
GVX4XvyhJCR8iJEtskFYTQvUKfSsZaBTr86QKPsB8ulKAwQ4OIxhq5e6j17NimbtPUNyzvs00Kkl
L+MgbvshFnaXuPmvDSdrEdpnvICpUgKmmYt52DilbMnrqvF94q76NQIoF5Dg5vUnfLHBd+I4LBXI
i4tf5GC9tAcnqfTj36p1G+zZ7/E03aAM8MzmpZcxSgRQhvy5fSXHnyioRBragCGw24VNUB0Z+WQl
BjW4l55Xk8DQRD1OQWKIHwiK0Jyq1KoOi760uWnV+yVWcDNb67HSTEXR3o+Dkq8c+DpMd1dBU3JH
Dv9cJoW+2WsXTravwSLOeUxn5LbUdsRCFgFCl+b8BCHU/Pa9vF9SUWXAcmbkE3oEIKM+nuXu7Ymb
hQ9cMlCFz02c13avk1hwku/IMbRFU4Wnhy2yN2R2nEuA87Brxy4JI8nIiyiAGbXettkXN149Uffh
A0y0nhIvdYfc+z2w8njfPX+fafc6+4aoXsiDeq7VsboX/Ni7mX7f7DTuzDiHcahZNLMY6V8sRL31
Xj1XRJ30NXI/n0odHAkxukD2+WBBPG/TjwnJ+gprNoiUWyU1IdybsDVg+JXyyidsk/6pQGabFXDC
OeHwXZATCuLllxJYjDuV9ZFkaqWMQ6HTlNupBpk6VYqym8lOpikkjR0SEfNxBEQSC63oOpvxR0YA
G136g4CfhJnhhlmXE1v9N9xlM1fBdFE2y1B1CN5xtBK7hZPV6S9i7St17Tb9Ad+QDUK6TYfPrUd6
rTr3OvVPycjQJ28qD7QoBDLoJUieKl+Kn8hMljQkUNYNmKgZfGlTJZeHM39+lQp9Ty/CpKcf/pqJ
ZmNYbciW3d+p6ImxGxgsqIoQY5Nc/HPodULOXjaC2S3kIa3mxxk4rgDDec74N9ErLOKsAN4xGKzQ
KkNGvjVqYMQNGo/jc2GG8f4GXGeQ2xISeqoEYrs/FIy6dzoUEqOGQvnbXv+zrGjBRM2XJKuopPEf
RnCZnTo77+wP/6gEF15rq8JslwOSR1HOPB6vBcipsQ7LBfljoAG8/s81NqVwBQwPcQLH9z7J3W3t
tpwXHGgY/64zIZsrwLkokGuFij2IOCO5ITjt0TqyNc8hwH//qn3EZt6WbdFRlLh/tbO1dC0erKBn
9TvEcYERYHjLvSktEKhlo2wwdYKJQYK77//HKpjZMkj0H1ChfWIfaRxnuGBw0MOOi8RII2MetY+J
BX+unKuHL3Doa3QLIte6yZrjlb/gTeAQvx4yqepFBVtyslgWkpDE9XAdSMn2/xdgZEa/bGTBfnvn
BJNukbudu6pFXUY8XAarS/xWzsNo8vwXZ2n99ZpWdTmzYG/irKE3Q/1hEq4NXeuwYF8eGSl6dwRk
Sb9odIO40OKxi0tcHrS3T1zmPVbObHB+jhm1iNOvzt/APV9aWDoKWPOldv/q0vLQOpbsZYoydUge
eHERExijcqW2GjOKAb1lWIkjaMGqndpoa0+n7kvAzGiEMAKwkZi2mJc/kE5um1wPqV5lkzpjsaBN
uP9EOuHKrjLQ/tC7ggkZYnMWOc9i/nlZgagX6YXGIq+/WEZaEtLXkmfOojZyrbiVEcgmHDfw7wYS
bkJC+pS83GmaHa1JLrykVgbk7MHOOgAQ6bJMhlyagG/PT/ghKK8o+y72SEuU5WCgo2ozhyqJL6JW
I7FPy9RcvR/U77EGE+3Pfrqe/XYyXQ0/bT/ehmTFhe3BXFYizYUjTN/8ao5lbEF0hvfTHt75NtPO
UXVsFzRRTTcoemg2FoWLE+CjJ1bu4PiEE5nDY4+2/j2MshzOxmyVQ+2COHhKbhjAcFbNtQ28IqHG
cpmUXBoP7e+V3s1de75bkLdVkCTgBYc/6bbjhk4yAUq1EArDsyfkVdFTTl8AWk/q6d8Kgjineosj
q4wWW5+GSuK5B/Om+NWtE3BFIym2E3XNjjvQL+WyX2SG9mxyDk6+5a5yoiQzQ6zVY/+8lcI90FhJ
y7VIA8noxttK/5eB1R0N1w112ReTGHoF5o1p1hOO37XOlxbwhHJOfHusNj6L1qy1i/r5c9WmqUxB
xOlsSPQFbYY4D2smRDfKVFKMrRCY7fpTMj/7yc7NsYxe1T9sNz0JsgI1ebx0SebMuan0AZYUNGFe
NHmzDOfuGOux/ke2KzB9zB4a371erZJH9Oz0Z5G5VmxwHDpNDpYnafhXNxPuGv5xD0I5QJ5n3x3B
RjGHes3CGS3NolE5gehd1ijEJfTWM9QgDgiD9g0vSbFClSxbLKK19T9uWhZ700RJDfLWyBw0MQFT
Gpb7V/OJb9VwDEvrJL5EE4HoNvGovj3WTDAw6pLSFWKdoxi10IF3nBV7ot1nrdk+YJ0AhuQUgPkk
L+qczebOaXRzpbFAzyTNwcc10FTfjc8efjKSCr15i321OKyKpkbfRqB8VQ4EQLiE3h/4ZklDxshh
LVJWn/CNldzv8WMAozvVUy0YqagCqPOs0DaoeYOTBtxzLywcTl2tWFt728tV4o7VAuF/JhQxfXoJ
K8vUkQgdDMRBdUUjrxQg/8ar61OCxW2LfFDAL6qFpaKsMjRqVcUsyjAMHrvrUaqGvqFYT8Ms3HB5
Ow6x4fHgIXCbF7Pl9tY2EqOJgBOy4dmLHtKjutcuDXxbCo6mFnU7ytd2YlbFt3f4A5sqjJxM31hP
ojyU2UKdhLeYW/uA1zdjJVChfW5kPnzKY96DKbwmmNP9tdFuI/jF+6H8gjVflWaWZyjRR1dyib9k
KllvnfIOb3/OdL+yDxUFabYsA0/vQYLx7stjqoTTDLRRTHpwuR9WVbkqz0n/InsoC5jeQotCv3Iq
Qw5gXe9vYSh+gxwkWBDp8+iJGpL2YDRw+ix6RqNAxKeZ/kpdx2lg+d1JfMZWR3tQnp9NRv7l66W3
kczv7U8eA8LCeiZkld2CF/wWm2xTAyrwOvgfbEkuSyCQwkZGhJGOxAZ4H3WWO2VTw6k1R+ASjsYw
c4kQ7Rb8JnOGsE7KvLCD3KmHQcY+c6EjPUt8sqkJuDYyQxAirejnDBzGiXocBEuKnhriTBFCzpoj
EklAIMu3J6x7wUqBzzDbpSgTNrV7DSwtQjOfwGCdYQcOufbqhOJlmQQz4QDTVybhC0bcC8pIomu4
yhKKJFO+Sh44opLrTuuJaClJRiuGRTr5URtOHQwTaplAqojtV/3gY/P9YiWYUj6p1B3NaxF6X2C3
1D3qtrOgQTy3GPx578atEcxNy1m0OiDMg9XGO9ASGtVfkq9rNb/mBCpCURggCt8TsGaYHYa5nGGg
qXbMmvlaVTbYXhlRMh5B05jS6/ZWDv30wLXhDXKHkQ5dWw4VPAlLhTTh+n7eb425ArJiEuG3b7i5
2pKqe8TzxKUKNpqdilIF/j4eCoWj8kUvsFUSwLpgx7C3uwdQusCyUKNhsQ/jPdMTc4w9NDQm+0VA
Ij56HGWnvWKTppLLmBQxuslCIXNxS4G+8fAgEzOkl4hcn3iJdhG+CaTmsSit+Z3rAlRFzVqFp8EF
YCo2zbmBsBFgJAl7KI6rFtOWxv0G+vO8aasPycP/2AiThWPAEc0xxYL1LiD8gLX5Rd1dkLNhIAXn
5697Luvbky/uN8bDZcv7MK8c5uUQSOekOTf5CHW14suNq3wSpO/7TkVUdyVidFtBSjBBlk+uNPvC
9Vrv4lkwq4YjzBBmeh10Ao2J7IATn6ypMhKDcFpIMvN6iM+oQwY5Sa2UHgppIwYHCux9EdMUn1rn
ej4pCrgIDoaL4TPPWpyZ0NjCtav9GomSbkOFPHRyRtR4Fqljl1AqH07OrY7C+G0yQNddd9vZgwE6
GUkp5KxKFGVbsxC+qM9rat0DhZqKiyOLmzBwKs8HGf2m/Ceqp51DahJly7Osgdun++jyv/oWV+Sd
ExyCvuVI9RpqmEtHEMWSmxLxYxXi41wW/2eIrbjrAultDOtx3K1M99b5N4XoRHjr4v01rtVQjkmR
3Tv7JEBmkkFhm1P76X/EQ0uLXE9fZnvCUSP0aoxRoldaZ4jbgZWBHkE0EMopkQN8OjMAjtfntv8I
sPxAiEiflsS0kJjFyvIMvzVg93T4y9GqQVTN0huHPnCbGRe9h9V7IbHPPGNmsJ6p/+g3yClkPi+F
nSyabBBEmigRqNFwrO9GHoWF2wfZSSWCgY6JVO7PUGEsXMMzfG9o5DexK0X2C5IBdZ9O1b2hyYCt
ML9v9dex2cLVZTLc1GIAkJyQXyE5hHklRha4HOX0V+X/7KXW/ktMGq+HvELxstgakjxU1nUbAzRC
glmZd1GA8L/rKuVuhiK8ya5QHXf5xs/Skr2YRM7U+RBDLqdYGltlpqixiannjJO4qXXDVG3N2wgJ
vTDPvRAgw95j3TVof1h1+SVl3WZo2NkXszPmpdXfDG2otzfYHRXizA9Eyo32M70nM8W6+eE/GeuA
qAxtBk95ACVTCCxStekDT6Ro+J6BOXMh8dT/8BXXPjV+D6Kwe6FpwoccvQbXwOE1XKGXLYC9XW4f
0hOFgerzQnCVlVQdnGNqMWUg+Joa9AbbPqmaakltuF4p+/kNYYGKxuLar6cBkbTrkk60eacQbZBf
uHpiJnEXeYxFd7PAtr8kkz4CLuirCpyKhVbBUmBxXyZXoj6aMqewiAMjlYzArv5IXgFzRdh+moEM
PJhUcRqQGhnqAe30CEU9sRFiQW9xaYQVdTXub8Y72ftHH6sz7ck75uscIQi+kpS4IVxROeyNAz2x
Fa6EONLlDWXx58jfiTJiHAKd31w3RGj363v0ic1aVHt5jX6FtMklr/R2p0Gc7vEUlr3HicBEwVWr
9UOj2IRPnK8iQwrvK7+vU7bnsSk1eYnI706G0qCRnJQpeyqglf24rFdzzSixRnCcuHQ7gPUVif5L
U+ZE4jRsevUa/4kOFzrK96CI5QrkT5a0vWPnWVMUYfmmBcYhnNm7gCKzdVIcEpw5S+hinQXgsIZT
nOaKNxjJsWFBOoWlxa+3PuhaHhgQ3fU6+FWtuDYYEb7UUQHiq+QjID7pOrkzdAHt6Lp2bbssCz+K
WrztfP+j4tVTpDbdRCQhGVt/W1xabcX3OBQFUQS8ta0m6/sGj6qtmYTX8iXwappM9paR9Zo3qRI3
ygYtBZYTHuBScjfLPXc+m99HPpUqCTZILJy6HXuOMPzHF34BhVaQN1FsoTRUEVcUNxWhW1tr0Vnj
LStpMheo3Kxcez20QJ93YoEH/AT9pjR0M+9aUOkamiiCKHb9oeTrOUvC7C04Ia5xzGvookz+o4NM
Ykmc+CRN8/JSZgUhZmwKQmU9lRpAY6YYIPARmGmuQEMalBt4mNGnPaoCRi2R6xGJHTUWbKBKpCRR
OteyDlw/tL0mwsAlSq2frpLZNPYKdm5iLOx23YEUX8aBB6GkFkUND0Rxk+R84Z7hsVFV2DOgvDv2
InmY8MrFqmihDa8cNxIaHPorrO4dxYn+t3NVIgWHWRmK9FdxO24qkjIN9wRAwlHkjLGaZY3SE8Oy
RJ/X1HsayVTuZBVBM+JGzr5YBzY4VAYHgZF9n/1XwUiNAA6YX4oHLwVf6Gb/dCoqUwf/iprJ/I7e
YAbbjQvn22tDj9KoiIE3miafhygcaLw+l7TY1OQIrr5Mov488EJ1fkKy0wpsGXTobSUgH26gejJQ
3uiouZMYLpbCOVT79xLjJry+4xzAnG07Rb41i0c4MKhAAdLz4+dfni6XVaqpWitkc24TxpZxrJ+9
BLSdTwwfWdK4AaMpFrSOzkFGPTwr5QyVNdj723EkgP+DIGEIP2TmOuGWpIKVTusrXKsZeYoSOT+U
Sv2R0QIz2932jO7Vs6aq0bIiIhOrICAk+pyAYKbcvo+MZ3ABAavzchZoeiawrkHYd2eai3FK9Tu9
vJD83sEJ8ZuL//lQfSAFFKkK6eehWJAEAg/96Vb2dMvg2vSVK3fxn5keeNBDywTsJwLavmDdYiGU
fpbDfxefYgCN1GbDiRwW9GLLrGUJ6SvPA4FMRXcYRvPRlOBRB+u5E4nu3+8KfQLY62S6q9qNB8BZ
fAqPdP8w41uSQTdFhx8q6BdiR4gEIoWqhHuaJ5+9aEDZHUQC2C4sQkPkaMGNUqr7FbNknc6J9/B9
EXhVV29b84Z8rgR2YneB1rZXtZzuhvT2rbElsNfIOyNT4VJt51cr36DGf3L/sQKBboxIlcovO3A0
+mKnPuA8Ho+joflITk/oWtVLNZXWkMLfJKQOxlq1QA/QMr1/IqTumP85BEKzFUq/4aVJDyuIjCH7
beXNd674uzOpqPMUV6papW/vgIXLgcwthoS8H+BSRFY1aGp+XbkDRMn04iFFA1ixbGgCtRkdgeEm
EKyoyNK+uIjK5JEFFMtmI4phyKhbeLm7m0poth79QYBBVeU6yUiZMybKf9dDgGiqDs5vzW6VZ0EI
H+elOMD4EUvpQUGyjlkStckq1NIxwDQf2CvA8Z8RTvKM2S/2pPjpPzSNCTz+mLgOkwL0hjRgF4wf
5iwzJpKQOnzw2HMNQQ7H1W8e6ARxU03yWkUO1Mu9VmF6lkuVY8z2xJUigaIFPWkgdqT7O0a8x6Zt
eog99E8yK7AeRjHYxX7jMCV/8r8QhOfgHl3EGkbMnhf5KE34soyvcDeYJi5D3lAS5AHMsbqDdCCz
COiy+w8tV6rF5cx4zhFAqfhKkpX/QxhwVgBJauvjpN2YxXrD7QDukdnr+mnrneQErMmIbHKbAQ2Z
zpEMV+J6L2URuKoOGRlIkqp1Ze8kIKqTtgJMdUYsD4vSPL/Zief5lR8zhTJU7XCJ+agpmPXSr+fH
ftTSsBAa3fWO0VIvdWmm509/2y+ZbHmKm0FueY069vUaQAqwI2VDDN3DDQjV8SW6Qf5c/3AzhGFG
E9+XMjzuoQR5G/YiWSLpo7LSMKTYVD2nlJSvME4EMgtKrhJgPIOqWJDw7WYPptdu5ZSqwkLsVe3f
Dl5vg3RAA6/Gu4lxblY5IKWp76Sc/V4Q5zqVxFbl2FFIvNtyH4F49fMvALRIJVJiR/2dMtMxvTv1
xnj/pYXIpe2C3STcSe/BquH+fhnR7YXUbICIpdtOVOCVlu7HxsJAJkITnALciZzt0h/DhjZTU+md
eZOZj0Qt0N5mBM8y+OUg9NPXjx4taxYad26GBNR5KMoxHBjPXNf5Wcr4RCTOXCeu/Eg2cXYVHZXD
JUpUnWky/SXUTyYnBWZRosW51OwjqMzE5z4w9Wz03WT+R6qZBhdc2rKAYSpT36QzJRi8rAQ2y821
aMtamwTYm/BXI/YGfT/Pexsz8vuzUxiYQ4hITWueNA7OBts7UkZZxorBCtN/zcxlzoVQh0WXOJHE
jjKKhQWRXneOqUfoldTWXYpAZwsuA2nsNtrCD/Ds3eVffompYsBOVkCb6WODops0InPhznpQX8DX
fNsDMA1dR1Lbgp/SgWy4hmsV/qH6xHd1hX92lWxvDKfdryJ9rzb9TgEdW/TNxfdjzARa08x71a5n
PTvgG0Fi2L7SvVi53barcdzjwhKkz3tfNoJ8L6TbCTZRiPAydzGs77JhLc5PKUz8e55Th3fuWrmM
eUU2YtKWHIjCOgJvIVuJcqHD2G0r1l2XUWOTMArOO9aLBGp2oMxr3tbXYDFgAyxONQYtmr7+olt7
q3PBB9l0yvGivmF0OKHs3NJUHnXHHhmbg61OH2XqewTph44rZAUZfEWDVQVEc/JWafrfRpGkUOFV
IdMbyQH+ZyMj8zO/LOOPSkTA+QHQLnl2KeiRA7xRiYX4vc/1VnEyHZGu2xlXzbUs8o4Dyt7IaC0k
Hv7YvKA+b4cERZ6OUY/z9TzwhMpkVsQHqaR0SGOO9mo+pEbnMmn9rvbc5EpTuxAFSOWW33dyrAN4
EOpMMtWKhIOMTGt+gKN7OUrrY89fn5cIPQNAVjglXmGE04hlh60T4FD6N/YS+gR/LbrtFqFpQe7x
DquJtlqiJ8VIonBHF/6zegTRuZ5c6t7LAYMtsPQeUVGGsz5Pj+J+MAgQ5Awt4PamlJ/5RE1xWHfL
eS9ZepKHZ1v3jzoIj/eyEHMExQ5eTu5m+OD5hnBQoG4BlKPuaXAFuIGQB44UIYtTUGC+hyVHp3Kc
6rcpmPGh0Fwot72hmg7i7ZF5Y4U6JZGvX0g5CL32R4HUoeqDs3ZakEfyhfbqFPetTRIPRqXlP54A
6xPJQsHw1GZpspHV4hYIhiNE7b50BEVlMuMrdI+vtBjnZtRnDwTijRNePwhg7dMKBRZs91Nl8Wjg
b4J7PT6eNtXOj3dOgc50pZMA72FWqNWDbaZEpmPgc5P/GGGxCEdNaFRNLWUTYsvOzT6Veqor9/aP
O8YWhLAjbyWhKaGn3JQCBRz0xWjutQKmduwqUuawEzkERKoQ1LmnKdDhJ43TfueLF9fTeDt5Z4hS
0jNAgA6Qr6VC5tx2miaqOids8+KLICy514akvSFGt7w1ZnzCpdrOp6lzmgcIRJ6GThZcMAkB7WBa
GJKeQ14Rozi0Tv19vd8YrF0U0fU5P7mDdGpgNvYyOBp3NDk4IJgF7tFOSF1INgvL+g0WRCtdetA3
DZI9DPWJ4YxH7+C1m9OfGo5gXHYIEMB0XIKdFQIkADGNgcFgVwFR8fcG0CEDe4ymkHDnebGbYgWk
EReocxKkDJ9pTBaaQvU+YlZZP217ttxkubTfG42t7/a8/Pq5MLuf+qJv/8k1G9M0EZuP2YyVj8mh
DYXuJ+N4QzTIq8dQ6RBTZ5KAIMJ+u3uY+KXK7kDAw+oPqJUUD++SSTU3hGVgxg1l/boCyAVNpH9l
NV4BKkduvgOBzFXVGKiHqwkQFmQXklTzI8v4+CSqGtA+22S8Bnco2bupZiAFBxIPvbuJnvUZk8xc
E8OQr/qYcQgxq0yAnWK/UbhFvptBhTaoAVRkBoEwD/oDI/Vg6/sZMbQh8sAb74gibnCCWg2XTsZr
sHTMGXsxw/WGpnk2yBqZcVV5pubFpAta0M4fdjyCyuDlPG3KMyodkbiMnWOS8LNV4Ix6NCtlgVuR
cCceFuQNGRcrTvYnN9fC2xgDlamyt0nItm49qILDQ/zbjpPo27iSrbJi1mhENXLsichwAz9IFcbw
ZsmGyHZkazvBpZlhqTu9sNPPxAzPIagYCz+J4o+waoa/GUdsYYViJ2gW2zfWCnh6CkZRrJih+rJi
3/xHc66vkG1whkzj07NHqTF1ZFroXMKe9p0BSaDamBJjYfGFAGUe3ebsX3GhmN1sm4ZC7+4duHKb
uLomQJJfH4bC+T3iNSWMabgOMTAJWvJwOIIPMCdgB+zIuoeo82Arwej1oJ0aAcTFoetiLhBdbIpK
uEQk29E5Y6tiNIaQ1j/F/jlViJDwe87XrdHRXaeCYog2OUWBbkjEnM7nDqmv0cofjWjbzOnJbDHK
w3pt/Euno1gdLpTeDCpZkv9gpKXAxOcLhBPU0xJRZ0IkTIJonFngCYRXosnr8L4Z8vZ/+PZLab2u
dOKZy41tA5tpuTVP2tOOYMSkoJWZ2hWe95t+/6J9eNgiALq7oQYhCfMsZmpIiTcgs3EcNriOiekL
qoLUVsFAQonCY6DxUJ1A48QiLyeyVbNA+/qSsiFq+AVo7BOz/wzR/MY4tmHGQ44fZ6RCoMkEl3Nk
R3rz2SN90xB62MemHqOV0DRHpIt7cVSoznpqicpgpsSw45WzmnVl3VsQw+PiMYF/dT2XPKsNdmnv
KixkPzRUzC6ZTz1yxFPH6l9nGVcZBXD4jXkIXcSW+JRrd8/P4Z3rvmtfbTiBZ7hyG0yk2pLoCU9B
vSAzB5xUfrxfa6GA0ChnQVR6NorRhWbHVXp3AGpaF2fwxr7yauuT3nOQNZfKkmmX9lGapzZqCjuV
cpqUfHcXqVkAwQNzFmJQ9H39ZO0tmiN0G1XJIxAcGLK1tWHN/h+UzqG+f/xHwjNjSWXSVPH5Jp9j
pV7Yx2mv0fMvaSHngpxHZ8Acgo8B2Xx30THj5MO5O03Gkru3ajiJI8SNuirJZD4LO4PXmCZf9ywW
XlmsEflZguViG0nFZZPlgd7doEPksRpRfP92hpA+RA/zDIdsv5opsxBiOcoHC7DSk24taWg+jK1Z
ioLJD3EF9WjAlDJI/GDd4FPVkm7b9I7MNlqOcUZ0UKopR2rDSbd5cjIbrGGbgfdmKvuaE9xUsDvL
8nsuNTGGOj2vnm04g61pw6hu8gwl1AzqnRZlqZiZfm2mdFvaEq5DKjt0s4N+7E4Km9nasnrtilms
oepgSL6YC3E7fRV78KuQnJ3jzSgMb9HUscYldVz8EbPbib1pXOz8ZEYCD2nww0FMejVWluNb0mwZ
1+ko8lDrlou2PgWQugtJt03xht3nxou3ErBEWgMnYlvaybf0SKQtNky5sNhKV++n6816wXn9GtOS
1I2Vie1O1b3skQNRj8klJcIZqLCf0ExdMVHncxsw0QGtEJT0FVOpg3YkNKC2jIJIcxJqwEIBZepZ
iVOajrjUgyQX6JnCjRThlAZqKmpwugRB9RDKubppCP65IjsXdwgs/7tcdsGBkg1dfSsmPnpaw9iF
/X7j9ooZGjzpf6s4p8EmT7ts62zrlzQbdDgVDGeOdEi01/fmKsSupjnxEMbfbMjuNU27zPYkAifs
Dr2QUQd6j9FSScYxJee86y3rEizocdiQNjLiQMEpeoy7NrJQXoc6/vFic5qrkGMiF04gSNRaBkOu
1FXK032fgUZIX3MUeeXZ/HT6bNTF0mPj6XH+DFj4IAOC7rAnZy5GLRee+dEsbnbMQc0XDAsvMItg
5ZQdfD0XSrO+xP9iZKUnvNmvOBtviOc5bGMjOr2nKptv8YNgkTkbfKNCW2HAqLXeJFUobpbUTrHQ
O4ql4H47jdW97ssCBTyl5eSsmO/RDPBl9SimIHXqv+EL/YUPNauaoVUBMMcoYWOuTrbbP0WAFAJg
JF1itpswcPUkro4++GaohVHiMCQD562bW2PcnakCxpNTuDvVdNi+x34MShdA6nw7UsRi6tWjghsV
yZBEtguV+Zq3XjsKPDdfJof31M+lh34noeMizQIDLVZbHmt5/wNh5UgU7lDgl37QwR3/SwGRR3zr
gUhjzZeZgpRbrLvKJFYKw2FP2Y4PE7/pbbdzM9Ft2iwdRu5b2N9YoWRfhP9Gi2iBcoB0pPb5wxR/
huRJ3Qwjjm2CWaHxyNAngKdD97mPiy/+1pT+y67005wqYAmwj1smPfnR6+3rbRQTjuPoIoymSjI+
LmC5Od145Vit5t3pYNHh8kcrrXpLbRBuC8vtZ8cxjtCmpM/u/g7NGNKUms6NlbwI1W6PiifwjeVo
6F4z35/zp2OtZg1GbpK9dlv3Ka3hVaFHxc2IzO0D6xi/zNyjCYqhG9xREGWAngTyH7MuKD0EpCQf
jtl/Ab+Af93i6ZAZtMkrA3Ibm44cmcdsdvoMpA7pWIW5Hxk3+xpNDaaN7QZXr6LiG17dERpGALEO
xA7bbNwGbMP4HwOrj72C8S2iTofOmOMQJ1+WXK0p++YxirsrL+kCo0KOR/Io7PD8C7ZuXaBFgrA8
OzffFrkZx/hfPn6vb/U5qEIaJ5a4blgRz13QZOPm4OInwnZ52f3LDvZbvAHlTRlePMbSWnFI/k+a
oIQdbWCSfW+5tvRWAGYXdTmM90DQVgE2z0nIfC8a+ZDT3RV4BFQZj6NZqX1J744QsRHGVG4QhyK2
c3tEzog+9rjsT5an8xHfUJ5L+jjs+3amAYB6ObCQ/zzVeXgOpYDR5xa1A/hOlnbrt6FHRCyXVBoT
bCW9CkWb53nUWDl3yu17leE8JKDadTMHRgwg8QCJ0v6YY2IeH8nMcALRdftWNpuoBJw3QehUY5SC
KUn0eySyWzNVWS8IfF39keqrC+fXE37ph47IJg3CyuOEeyv8in/xuKgbyHqsRK86iWe3PbU9jQ4A
6pMmjwpDmuV9AZFJp6NwxHE4ome+HkZdIQW99BSGvc/aQ9KALp9tdDP1FGi9T2JMBehFX7ooZ2gR
jqX8+0+JgC+PBRL5RWu1VGBBjun9ZofNSjT+ll3vOmjSdsrEi0TmRDykBgsDsIt6ricncpLQtBps
nlYuPuWUoaQLEk+rmf1M+5ssGMVZ3LodkOsM3IrvJCww9W5OXTYEel+A3n+15bcJxX99aO+1sjUD
R9S6ZmqQfwzKBc0ovaygkti8G6XThGomogREEGPwRpTePudxPNC33IQfFPhusluIsqokDbFWoTTi
AM2Ml24CH3vPC/IfEzjR/JxU14ubFlqfO8wy4Ogq0LAkri1L6H4KuQq+voN4hPf28MUBKxGkeyqc
fn2/lui1klL/GS794pxatHs2fAovNgekRW5HZ5IjQxthvgSyjeYHuAxeB/YOevSLoxK4JFhEdPn1
V3DYSe7eQ830zlsM/k3rHuvDA5RpEYG3yzrLE7clINTHBE1hMZb8AHUfYYaGln0SOLeBxji6Txh2
xgv74hdzhGc7HuJt8krefxaEK7YjNIBMus1PLv0TsTSjdIOBhqug+uTD51j5PHQQMU3/+VZK6Gwn
IFojzkich0sUj+0O+pDH5NDIggky2+h0T6QJBcf4+o07JmEh9W3d5qnulQefWANwUslD/k+qbHAr
457YItQwd9awMoFf7tiJnEA7HgSkF1aXnWZOQWGILAbHzJD2k83jm6AuP1cncLtWJxnCotDBPGQj
2ARBikSkkm/FrdcXlvZ97z3Fj4hpooJeUNkhYqCny145YHSOciJNs5P8hqM/AJxnf0bpsfl/Y227
XvukLaY4TR3HsAqhT593E0uuWHdUC7AhPvv1OXz+Yr3QnxT2itDIMn4w+7K4NGFT3J54hs7RRe/6
eIf74gd7K3o8wuF5agMU7a9XzSatkN5+rHLsdcBHYT+XL5oKho/8TxgAQZwa10sjUx4FAD3E6aGa
rKqJdZZ0ZzPXeyL8g6aVcKtTFmsOs0AnybcLeT6Hhk0ZXf7vxiGKCzAj1Vzyqaq7g20KDsbagwSj
lJ5CKMwnfX7kKTv/b/bI9/oJwLgi3yCfTbM1Av8+lILjienQTFRibJyPFSSZiJWzIzE1OUIuBqAi
ZDPt9+0EiewnvEHsMCZ+Q4HHMPElQiYRibH/VP4LzPPtuR0svKhmKmVre+PvBgMsLhRC8CHvUua0
y9wxGyrmBpBWu44s3Qove76qMvXXsqqPrWl5i+6Hy6OtrmBuczpSLZRuYja2zh7MF1ufHluRCNUt
uej37bDJ/QFibhnLlMbjdclzry5r5EkX03iffTRoAoUpp5Q1SJZHQqDGtvMloYAnD+JVSB37C9Hm
iW1sJgdgHP2xeuChCliRgvb+whNS25OSozNb8UZqxKeP9BGGbijrjGMptsojTK/QJk/l7uAWTqmH
v0a0hT3TL42f/AlcajpjN6jTLxETB+6O+gIMiOoHnlnmgWgIS9tczxhEgZRm5SX3iuhaTpzFqXGl
XSvcayIxyrQw3iEh9qljjUJU8vLzADSEB7sLgpjV458xiU2xThZLwOtICLaj9BXhwjxLV6etLxGw
qDTwgxYBAwlv5yfDeIChOP0yrNUguR+yiNtoFSDYvU71cgn/zF9Yi1FnciMw0txnYtF8jHOoAlbw
pDfx/goEn51TWtQwd3V57g42XIBDDNLn/p4SA13rzBCSgk0XTzzxCOzOZfmVlb+xXUfWf0tUphRY
cchO4WdIjp5oH9qEA5sTtWi3p9VB3HDnN3QsIuoxYNdo8U7CRKf5hy229Lv2c1QIOdcuCvhqM7Bx
te5WyJV9zeDJT0KHp2v7lLIALlH9NNURUmL0udN/zbIOQM/A+jNvVkfjJ4/Nw36oy3bhBfuWSkyR
RT6np3Jn5GjMyJ+2KFlNd3CrUNAvudO+22NK3cleb30LUAGvWpmrPE00sdiCiobYNDYmFJAs0P54
OC6HCAImtaWezQAkGQ9Z7TFeXM17A60XqHkxSHcPsOyDFXQTEb6eC3B7A34XUb2rfyMhCM4yW0Wt
FVf67DdyOrEgBxnLFUmm3nv0+FXSMo+r0SQSnlN4Fp2hVjm1ZczBWrxlnIvDUhtLu71mr/bQ9RwS
0JbA93pzC9Bj8b3wItqWSS1LIfXnARV81r9bAFfrywBnnv6mT4BchnyikdjYUgJk9I+Cgb4P+3gD
0vLW+2i3c5Wj29tyDh05CdSVcQENEsGI9GwSEtZ7YEp06osQ/ym/ze+oyva86Y+rKXzheBSiAt8a
JW0Yr2I3ypYnGvBXTkUV0Ns142O7XLu6CTr/cAgYEQpHYceqAqsB8WuFx6AztBwSQVaNxvp0VZu3
w8TGWswTeZpNv0+VwOl5j0uYGV01S/e2uvQtv3SFWPXs3vVKNM+3iZDXJyrwvnd4r4CGv5DBN5J/
HxJA0Fv4bwXSp976A7wFc0hamvozcNbxx+/5b57pw28P5ZAKMv6gNQel4Ib+1QGvitHdGSazL+9/
Ncf9T2zspyjeD6jIX8jN8sclS16wEo+lSLaNlkO4IrTdI5QtmJHgk7hcmdo7RUOyqJKlXsHaNcy0
gfVeJdTmrrkkomtjJiTr5NCWbXGW6i8lb6aNbF92QpvGHoSaGMpNEMsY7XcVg3xp0lL8HUUC7N3C
hcHCFHIKmdQr9rqTRTK2LbnaEZa/ygmnwbMkxBvCtP4RHja6EO74QIOp+0faDQH/NNCF6F3HjsLj
uPdBn/rVn63+K4MR3G8xepGdHZeO6zE3MUjbIl5mKgHAh2WVDcIZKdaG9FB+G2ag3Vjo0XdLId80
eH1+nUH9PGV572czo5Zxj3PCTIr1ezQvN7vPNCH8WsMwGNiY2Pl3M3JeNCuf35mWltcsVnhuxh4h
o5HmYiPnxUIYej5gN+M3rFPywXtqnA3KpSYEJV3Ift3u7MOKoGTlb1fUiCL7JWqx66GrgevettDV
W4Jphpbilr/3hlhkhX4LxBeyY7h30e3HMoWhCLPyfPkLQh2K8BEXk4fI4n9M5fOy6sDxBlPb2Qk4
K9/SEWfFDzE0ElSY9gbeQkff3qsyXQvT3qJugjlWhlHcYGq+nV1LTLNpqV5eC3sAvesq4smXWoti
/um+VOwlfzK/YWAqsHC/vv/sZezFoJV5WWYLSb+cR4DiPkVKtVKdRAKOKZOLw9H7Nnzy0WmytjST
/rqezWtIXckQDx8of6rZQPLwtyl2C4K8+SRj2Ro/2kVGmdAx4BnQBr8AxW1D5qY2+y9CBHUNhmD6
1IB0XueBKGP1vjMU26P/cq8kUdFzm80DYWYlaAVl8odxXc03cfQAyuI5pbOZl4TkM41MGsTZKFMk
xoy2bRXKWZeKKO92dPgXq83kioaVg0LphetuC8neowLHzRL9wSYiDk1pZ+sOgmYHSTLkMuiK0MYZ
ko9DRz+dqYQk6O3RwZx8lHKhcdyDeE63fEsZCl6SAMhfq6s7K+PQKHxh9aAgVSIi4m0hmG28utaD
HZxRKaz5OolIfpza4iVXfiedd4t4eAnTY8wKr9JSOzhfSDApUpgTUxr91vfmAbYF2JF2PZEQ+tyN
3kZSB1N8cbHYiNY6HuWXFD9zpfP4bDFhTYNvvoEVF3kJ13Te4jD11pVvTUtgcup9r+gXREHdlMw1
C97p4fbWYBxJW4wDtrx9d9NO0gbc08giyRyqolwjFQE1S/zoJJa1MewQwaCcWXbS929Si1ilH6CA
s8fFdXUtYgjFhGoNYK7FY33lEDwYDt93VSAvqrtVOt092NcqS9KYT2WdnpBTpg0DuLavyou86dv6
v55oeKEZmCDewZH0cFoq7/Td5h40BA1wleMY7Lg7hN2raWhE0osQ1UOMwqb9yW/qG/CdzBBmapI/
I2UMbXIJnKNgQt/v8Rtxzz7UFF9Sm2irp9Zl3JRamI8meZu+UGusU1WOdJD2dQriFFJLhgE3UxUs
e8m3LEaj2CWvG4gaHXmYyHk5f889mN4aCB8t6x97uhAJ4ZiniKU4Y6hTEroePmV5o3OMx5q/fgFB
vu5Qg5fUYRtPLJqp55P+CQ4ZWKV+CgNKy23t333FR9786l/W6CsAP24ZrbQy7jfYp/eLUSABBqmn
iJMtzSSEY0W4Rzu3t5gtD9u4ELxUB2eXiYNAzDbDASwazRFSajhud+YbN/f9XfVOiC8N/tIHfXTi
o3djVBQE0cV3jOyvSkSVB8ymogeXX8m+Ir13ahQo/i+x+7mgTv/duouzunw+286fCRgm8gEFOtKe
TODWjr3YMFWwgd0BXDVyQcgRphWYb22WoVVZxzpjW9Sej+S/kZFx7QBpNFYGsfoGRahxEweM479y
kLocVvw/Lq7WVSPy3tKw4We5aI+3jG0YIqWWdU3P1yZ6TELrl0MhimPGDfmMUd8t8c3+xvhWAl08
kgF1wO3WiAMrzB+op4475QOp1RLSc59uCOyocD6RvVRflI0FsRu2ng9BKBvy/xaFObse0vf0E0Vo
aFndZzoOo0sMIdM4jPm7Oxv+o07w73KScwNcYetBB+hyfkJI3u2pgAVI4zSnBasGXz7/nSTCjwrR
4L16nP/86tTPjyxisnHBMbXpBu7I//AAlRzD76CL11NS9z92XdK8QtY1TTsCMC97nklw6nDjWF8H
Lu+nk/ctlwwk353Q+ckkJDtvjvB+I83MXCXkOa7mUU7Hoz2YsZDfHIqIpHy8m2YyqQt6uYznEl+2
Ndc/ymdWreyile5CR6B/cmYBiEHiqxIz9X+4k2tZtZVERO3OF0728KPX2ERTsf6TF4VUtRAYzTzE
h+VCfma5sRL02Le6fHwI2KXTwciZ1T0s5+Vc1sqy8CetbE6VBIDX7mfEQJ0taMjCCQJ+DG8Vt+ly
0HPI798jU1rGPHTH21RMLl8LFv8y7pkMNy4zLwK22L1eGxzPs2t51oOEdmAAm19NdCb80nk+MY0Q
Ypxrvol/TGZ89Fp3jn4IHt0qYxxvMSFJCj2eRYw5vXOFh8ZHGSf+8s7TTO20HqZNsPDnV/dxZROg
ujBNKzumufAVcLza/DPODuoY24KqYa2VLRRfaimk26cuKF+VdI2CcUb0TDxyQgvHph2QSO1LGftV
drBL3kETIZFtmsSj3EbGDcxbveKX9pkuAuzY/yZ3Fe1/w1uBzeRM/y1dDnoogxT96tA8hZOTwtTa
1Vgl+EpOzMVAdcNpQw0qmyTdujGFq9khsziJkbP/kos98sWBCZk7P9+wC849mhFRRAE0p6sQ1Hrv
Amh3W4pL5OFiuuvYgU0EqKVe7XoHvc6saPDBfoL0o3Nk+vU3vW9ll05S+PU5QIxge9h2xTlTgKKl
xHjFSRQI/yjueEfwwVXQpPmtVBudPoyAfpwabwP/kJNIpGepHZFrVeX/qN10qJQTTSwUWHyXwCdf
lpW79PVCYjOV3pzNyovzGvbnmOpkR6dSnsVZXXbG2Vm4aUYdzp7w1AciVyc5KiyZ3mpiBgQKL7zP
gCbRSj2mPWkaSKYj+/Kzm+cc4c66Kw97rm1Ii+2Vbh9DhBCbA16Ld4/BEuA0Q6rYRDZki9wGIvB+
DsY48XFaTl5LWV/MYtwniibqC3xv1WFO8fbAQG5mImP5gCLpJzaqadJOCmR+xgjBtPfbHTUVgkqe
3Jy7WA7v0hLFHMVNw+YbjpBOxBCXmxUZNOrvNUZuSf+lxsurM/86/b8pXVNBt/nDnMjWW3vHbDRi
nFWKFQZq0ZwR64/+UJ7Tq383AQZICFAWvhhWNhVZbyondsI7R5d/YPmoi9SB1ux3UL4N/ZXZxXlB
ZTxMpDJbk43bEcu5PLSsknmexA2f0LAk8ISSSkijZb1auqpqNz0/dRFY+pbxehZwzuMVgueNX3Aw
ZL0E+LmQH4KqducPxW/VIETaWTyKpRNOl80e02vaL9fb9KNiBT7mwG9mvQ8daowpAWEzbqQfC8Wj
rSbNM0Z5M+8BmGAeyr1bvyUhUCQ+20j/qF1th16AeRFCx5pmnSYSpmLwILaNaI6UuBdJA9SiRGW5
i/PJeYphBMY/D0h1TUa5iRqyYr/CoOc65A9U8/YrujTakmUo/PbRlsx9A+AV88RmnJoHb501PogU
wM2VV6jwoIWlWnNpHNqkMY9T2++SdcbYtshyslW/JPRzK0Uo6LmBIhGbwbONUp/1MNOaGG47wD6e
D8xflFjkUhZJKjYrsxuLWSzeAaw+x2aFlZZk0uxnZplDK2LsFBiLJa9ocPXtPPMzrR+mDdf00u8z
RPZFGdAMMorup09OG+C1mCrBzizN8vKxDez3m1S4tc+IUCw2EgNovgLNRQoXOdgjKDdi85fYH83/
d0F/l2BWaO90lZYAtUgsr+7Mhop1fX3diCVZawN5Io+AWhO1f+tK2z66NzaAbnPiNBEgRbHGihoE
TUpXUWzAK8EBswzFgNFRc5wZDdUmGGDwdPnMbPramkj4iq7Ie3366bDhMGp2gPKuyDo63fouTqGI
KWjWgVZe5MzymUvbzWdxCRGiiSZFktyq5lE+6QAkEyrGzR52SqpoarA/NTSGj8QGvuIy7LXvyr2+
cZyMMFbZjl3HaLWhZMRSpqOhizSq0AA0uu41NmRhiqqwNlNoTh+WK++gYIOMosKZB6A7vnnSA6mY
sQyKDQ3Ck/M9Q468RMr5iy+TiknnYyqL8e5Jp/ezNAdGvUwoikA6JYTntTqHEF8R/z/Ha1l/ib4p
8tfnDcyN21NHTXZYcPrWoA/IPnIUgQAKhp95ZxJ/zAme6C4BKKKue/KeANg7kNT67qdkcCO7+PWR
cNw4l7Vx7c8tIKhdA6Ca/KKcT3uxC0tOVtV7WEY0PgbqjEACyZn/jEosTYzZ/E3QsL5K147Q1/aW
cK3mWOU9n6S9G+23HV2uBHOhwrdzYQRc5bpszrlGSi7ut+OzpUq9L1h2eHMywjIyuj3rErFvS7hX
gr4+nOixpTPg8wFZs0pTV7xgC2BZipL5fdlan08WNI68kdlsEKNvEQELnKLOq4PfX9a+CyF1m0Gg
XkskFd7w2cpOE23T4dNqXTCr77Yu9d1y9ixGXeAjtXlKvWW3xXwLe6lIs9gNrxCGeJmSJjXEekZA
ndeLidqocoZIFLkDrT6AJGOXs81ynKl/ZOE863bw66qdBIOMycMKpR9BI2UOFcQHbw1e7yoBU37L
32PMECJzXfdsGzqthijXV0iX6qrZJrGYZTHV8ksEJmP2f4Qoz07b+jYU61+/2tXk2yuhMBa3NnsC
8eHvZcwGRDouajn+2kTSeHQ5GtAVfChEkl0JVCyPVF8DS4DhEsCEdLYdNAKBAjKBAdul+r2qSMnJ
uVPuO3QN3P8UJZVADKt5NB3JbcLe0RjxORwNqJiJwCv+lD0MQ4SiwyU8Oo7iboqvU0Kjz6FBgCf4
i08QUndRa2vkoqnT1YYNHo1ogUwkACoL+z71oqUSgLzp/ArBFwyHoZ76bUxUXvx0JQV5XEq43UmQ
ncVgDtBUuIpVvjBOqJWw9N48leiGTyjoWg/jE6HCRaTDb7uElw/mIzqKAqPTcqUcmLQhqrhV2To2
4iHuiFe+Z6n/162YFOZIlwE/kMsQRFc3lSEOxBXnScFPxbVBpcQmnmjIR9tEch777VW+CwrjZnP2
+6duxZ2mfn04/E5TepDCDsJZJwuvrumu6P2KzRjGkS6CrORG30vO8yzd4tCS1+RnGAj1FQBujeES
FoM72hsgHqM7121qgDv3ARbB74niCEuxTzM0Mq3qKdEJNxjKzFYGoagui3+AWDN4rlrNCHwZtV3G
gEZo/Eeoe4gRADjYrA3wLW5AQVC+VVW4c523+UT51Q9X6h5+YcufoCIZkuirHre8QYo10UX1oDXL
TJhzCnEAjiBW6yBHnL89QPaOqWC27qN7Sr0MfpQuUDiHRmizUZTIIeWzZsRY1UO+ngDmP1NcQzK9
A7YVPMWF7qfr85+9HjTDwArYJsh3GmWVFbow8YGmTNe2kP6FpLpX+MTyBmzSSCeUotY8s/h51eba
I1yng+ZLCnKHM3+/k/T/UXC0k3DycIjSUrYqrxuwwp4CeClPX8KtLf1obmAbdBJXPHRzZaaB1H1q
zLy+yy/nTno54Oppo9UKD1o0VPbX4KwX7aL2dMtrbkRkLYEJZqScXteXzOVVtAGo1NeCUOwQ8r+J
7Th/E9ufxb5cizkjnM5WUg5zL+nWSkluwBFpC3RauVKpwJqqmd0uCeYUEjckHE8IvfS3qAB6VBQG
bVXBLVAXEP7Bv34WbiAG1V2RyazMMxGYH5jfuv7ygR2f/fAadEe+FP2uDCucMOS1vICQbsa6gI3/
4eKEAC15CTAhwO9cOau8z9p3IT5M3KCQ6BHcTcx4ZFP5PPmyZaSuu62xGjbvEsNecw/uCahstUJ9
dNDDa+xfhZba/upMeMj4f7X8g75E9pwNAIbhKW5RU6YHDUeDjwZualNLGW7rlrAX6G9CRErDahya
95imk+Du0PvsgeIfqOyjCRKhi1MvZJukFKy73VM1JUPPKFARNZ91zOUzqqpP/8JwR+QZDoXUUwqU
7bpIYPkfQrMb1Xb3CF0Br1NAOhBTnbqzVijcsFw1SgazVqirfUd8tkb4EJMR1NaB/Y5aAD8Z/t2e
exRuTnr0PdWrbvnGkLS75vbi+uyFQSp3qBAIxM4d2oz2xj3H56WFJwEVBA72N93WgFji0N8CMVcO
DAmgpxBHo6OxF2XGnOcVqoyHH0Qri97J5lpi2oHELd7eWwlqOBW4iWXcbBdoMjmk/M7z1ELtb2S+
OyERKwMzeI3Fcnvz0ZeLv4ANqqaItZ+nX5Y+61f5XiE8kXe20CJSoooGHO+MlMZB9Rok9avX4Gwf
adZXxCaZru3zT3xyRRIu+uzxNC/yPXx5KwPbe5zR4Dtm54swegZRFaSEhqV7rzQzt4F3T4LPbzdT
OtmfRxRhqOmW86ksSM7JSACJ3M34WpOhmVM/jsOkDL/qe2nblGy4WuGB9K6onL1v8AZQ8FDYMtgU
W5gf4RV/EbSLG4CMR9EFAzOvpZxIPRtjCgTGY5kiYgEC3SbFQLjvf+Mh57hVO+2yg91/GZYKhKow
7vx4haENBKGrdfelCROCN0lWaM9DhiODdXbiDPGAobZbJ3MHDpV/GIaCXxO8vK4/mpp8J1BQVhrT
Li4jSB6UL7ZAySyD7e2tVs4BbSjCokfLfOH/Vq9vnoQlneWsAxQkE8VwcDl2zj6/d7G2M6dMkpyM
7OPFL0lQBB8P89j01OKkFZpiPFk9h2xfrTgQxpXB/rGkKm/EHkeVvaEbehn+0Npny67QjRqqYxqb
c/PS7NRCFhRTEGGdJfNy8krzsvCf9EgE6NO0RhgUfVLJ18Xp3AKAPEulfymN0XcfjpK1nz5udImm
nfst2Pihf27hSsKsXqRHgPY8jBTza8Iiu705HNYo1lKWKemfEdmBi4xqKdkvBrLYVTWuojN+qOSM
nKZGGdq+BRmGbyACil33U8wxzuOFu5tt17qw7NIXnSxdMov62ggqj5bqs0ZZWmsK9zz3LEGM5SRq
aTteWUzmnrOAVLyNtfjzFDawPUop3gLs6gBZm4B5wNiVx29HX4jp1M/ygSODtrpeI2O4VLrJYL5c
PtsvazAkpLeVeluZsagQHEfDgkrEJ2i9/+gk/kbYaZmtcPcmSL1RDt5kMDaROgqtRIZKQxyg6aAM
mv8HcyrPiqw2XbITs+y03T7CT8bw16nn6fWCHPn9Gq9HXjZo+rKltAUk5T1Cy/lwOuhYtVcKjdRj
ILh8VPZxO6lkzdfeiC3x0lNw73En/dE/x6cmJ+5n4YgN7OqAlybV9sZvv5+88n5DmcuP2OPVKsEE
YBJEQ4rebtyyxzdnvJlzMcOU41tlYHJ85TQhNqaFX15Jqma8TTfE8M4RxMt2uq4XM0IirBlUjFas
i4PimOu5R7cDn2RZAVCtZ1nhrRD3LtgnOYEHfWnG0U5LwYgErXD0UN+DaEY8m3WQl7CZXQiBwYbu
7/DOQPjy1ckiwCmHfK7XadZibpv47UDvsy4hEJhDrxP0hRoaQNy0WGyfLC613NaIf37vcdlNJQNY
XsgodAUaHRlJcSW1iebFpbu8Qq6ypvY1wnzWxWL5xWUANete8YpzONSMIktXZGWlqvYIkAvpEd1X
FVYzcvfxXOmy4Ig1sJltKa2Zv2G7SVd3UkRSWQBptk5aqF+ewzZoKN/zM6IEjn2ox3/cQjXOAwLn
P2TKbrY5YHqCMx81jGrtjOTTranfYUgYG8CiFxHe+N2ihEfLI0vjXgEWYPM64hioK1wsQ+qFP/kP
cmdERRpRv0ov8PRnSbM9NfHcONmcGIbbYKvSRc2Iz6pH9M61NwcKGQ/SAbpAaEjBjKBIPeE+YTmL
mSWlZ/IPN3B7evMhCKSancFgcDI/ULalu9nwsojaCJp2/yXLYTm+C5mcwDzZTvoaJHUZ9jkgTUhI
b8XKUb4wv5jpz99lIl/TtJyD1PSLr22+YmhaTPxj6IALzsi/6ZwaeDVp59/7BTmtkrYTfT/KofTk
1IUuZ/gUHQF/uUyhjWFU+mahVxO0iI4bf7wQt/EVoi2Ldh0XcTSKz5n8gAZlRDXvp4H1sVfzxVCt
QC4YTMGVwL3pJkrCVsuGnnwyulv21KP47Sy5XCO3RLDP3GBGj8viBktwojIsZhIRoEIKIPHh4Uat
4e5SwCNJAImYG1ddlWVlrqfj4hhW/l29xF9r63n1xVGo2qrrOar8WJRqTVRu5rvCpBuobMhA0j5H
QCkiBbd7rkaYMYSGu9TaFBHlIUJechAAz67jm6ggqFSBgok9Q04OLlXwhZat5EMzqdlNlZo7Eq9B
8pYmvOney8Qca+HtiUm/YsXP1dNUfelZzMJ4WjbQpFgxMzblTgBmurJvqOLd6Nel8dF89j8/V1LA
Ma16uiwNvhlYgUK7WUyg4oIcUefKJveg2/c3enval31QGj2+PyoS73fRggNO0zWksxry3PToNIGm
3ZYBUxXMD0fxGGzksKA/ZTJRk/IRY18lIJD190C6Wstu75maaVpX+twXCwRz3gvxWHPRYsYKp2kH
hwa4TmyBZdGcWwoXvwUTFNoFKDZ3G3lXRMDMI2owZCvcMnWHL3V2pLglLu9rzqzHcjwGyFzaEP78
SBwTRHji5Li2s5z7F5pJ5YbhKRAyAUeuhhbOnimaaV6l19Ebut+SP6AhRlAa/6C3kC/7Hy1iq95v
9uUoNEsfqapIeG3i5ZraqQKZWrPl8fcGXjhlTbXB6x2+7mm4kYGyh8O8Zja2s2J6tzBDuzKOy4pI
VYiJ4O2y18zUFWvoDCPImj/E4jEA30p2UlWCkkDw0IIOOM1oZR0H0fdin8ZvWJx6Ds4HZsqEn40R
86rfFElCs5WfN9lHnvBGz7uQalgMx1mtatekzM7koQxCEKYjEWS9/GmBrMHY0cd7daStzIERwe4K
+sM7hAN/SEOWu0DONY+kbYui7XdtkCIhog2Z8gMpkUzdbrbwZm68Bu3oKtIR3jRhht3F3HZqMPx0
ntd0KIADZ421gm/nvQe0+FIvz13V5UbqyQ2gp3Jv1BgeOmiRODzeCu6ZwUkRmX9i04FPNk7+qBVB
e9q3dOC0Mbrv3v+NzR6CFGy8bJj6rt8Js9ff4BE1+W/105cdOGFnhgbiE+/9zzMmypLY07NDt189
2454I8oA7Qbg7+Ju74njjTXNMSPI/sZyMS63uEs+qBg+R4p0kP3AuvosibvPR4at85AlxYt+x34+
RvrD1QZuE0ra4jngzhZ2PnPrRHO7CMn4wHoHTGu3uI+2nVTYjZHgBkOnR0xoga6QWDNVXPn6f3H6
CQg13vUqgQ/2yOqHZuI3wsy8ol8pr3VEg/F2YH4VYqdhUJlYo8ma5NeQjtLOMji9IsqtY5zurjCw
pXc3IKWzH9Tt538JRJnpnnXaDwZqTtTdcneRoAaOrv6SFSeyLJwRbbMsmyvrQRMILC0MKbzbK4qf
vUoGO9DlBNqjiMG+Luvntpm3vZ0hn+pR4tyFEvz2Cl/qjW2K55C+S9lWPJJWVhrUcf5KZDqRQsyE
KzxomyUcSaSgzymnuuZ57iCnjY1RE2XuOVt8Ox28IHjrlD5A/6u+oftAcjeTjlwdZ8AB1+UDugeU
uAbzAcQxB22YjLpa0OjVPADv4O6M3UzIrhJttRNRSO3pSuZlBHYGSnBRzgqYSnKjNIdtHZRpxZLE
pb7KLPd7u6c/GSZ1evBeuyE0FTZbxtNd3sQpjqrzJH0PkwPNangpRa1+AE5438LfIwSowT5MNVhm
k5xbzHpXGR9XDMWIqY9IxwFz0hrGO38TqXccJI8sgF0Ovlw6yhjwckJx/PJqijnR0A7SODUQIfaP
b2s0lXGgNKDrYp6nwz/+991xSGlHwLN+LBIo3daFw50I8Ya9dkROrm2IWrehUx8strK1g+6Tk+FR
r7841WZYxCfjmUg50tIusSfoHbZTrk6P5uLKgEVJ8jpJURhQ66xtf8tgcsizT624nIhuhNlIywrW
E4XJJwxxKDGl1nNb+hEgvUuLk1yTxuVTLpWNsv8xY8eA/u6B75Gb1NAtZlBE4NNiu0S2kcCG0yZr
q0Y2aZf7gkT3rDwq+Hy8Bsq6OSZo9GvAK3lUvgwzj0qIYzeak3onG9e0bcWjTHjiPu69ZTBnC6Xy
BFdrzQSmu8FNc+4s8niUvdv+OAS9M/LLeDls1tQwfyr6FeNiWhlyYaYvumcIznG5x7LlaKpGrToH
8AEuOaZSsKfCcR7NkVwy2kXwJImXHHLJzkU9xTSATHrSwpBmt3FCYSox7y7OPc2djjITJcVboQHI
fFoc4G4uD8T31g7khc++2z4ehdkQadSr4ju2DXQXnA7lcyFCriHveKM97bcSqW3NJZ0cuKn3xsUk
Ya+Dpt1+zoS3Uh4cwYUb95oJXbA9i6DmVoF36gLE2LKoHn/OtX7pAnJzkS4/SUTcUtAXnB9rYHaB
lweUFSvo1Co/UixxjUm4Gq6W3728tPPAhyeMkkqk69nc0Bp1sTv86g0X85TfDQ5UxnONexhoeGYi
oNCAyYSk8/Fc34r8YPQ6W92Qar1MCWHsS4m9/+1lKBah7AYXGiPbd0qsXYdfEWm9228F4OPrMh4p
1G4bGzcT15qCWpmZIIF8/58F3TiDEcNEtG7yB7oRxHBiQrLBB4r2fKC3jzl4IYrkfwjGs2QP59TV
anvmY0+w03O/HEkrEFlRFJfekqu1uZpxaQT+gTM5SL4zxcQQz3d5Cwi3r52xXKId7u2GFZvdmXiH
154JFgKM+q39BOAAkwtpHhoOWWZhUhNrE7R+1ek1KtEoiNGEWZis7TOs3KY2ioNCKHrC/sSSWQ3Y
A9U+U50JvfmJBnCSU+QUVUGTxB7byfNuH1Khg8csyEnShgxFP5bDhTRykfbnn2CK1raaShEd9zfJ
qQBZ3GbtgBZBfLyfD/svhq1mxIT1tEiMddXzl28f5qyMJaE3do+rZFGcQIecGIlyFvqlEZtbJlGM
7i2INfa2xt+lI6YDT210ui4FJnK2IbTA6QXVSsgBzl11oOz7BU7tXwzhDaGVenX5J9qeDNCsTMla
+dBsx7DB6UwCA/ehqXtIJdBtdDwRtvoeE3e2WofY7XJj/8mAe7Q7TPt8TR6C2KWdCGi0Gs7mBMI/
jroPvE6dybCyoDtF5E387jAx77tCgir+3kRlx7RpO5qfHReKOecvXUEKGJYwH2yWhM8xuCMKOgqB
Ki0RctWxoUQxxCs0yVQiY9EytjZ8UAwAZ2hM60iM/O8C2ShT+F4q7m/Z05GI2aGYePqRogDetvvq
34d6hRpDU3w0ZTiFx6usdRun2UqoJW3mJMSBVVbT2AfXxdU1krDPzQXOcKRWv6xl6GXYJikxqAEo
9XpXZ+VFxGRhwG1b8+wEvo2uHJfNiwlY93A9ti4RlSiX6XEzzQcFdMQgormHDdjhO0Jw7qW0UhNh
fQ+QsVgtsqboBS6tW4etT6Hk2LCjb3KjyisGl5xQzYxvy321wMgLkhGtb1ooX8qz/Ddyaz2Rmiw0
iLofnh55moJAbsrVQ0zkLXle0+dpUwRzikLFTxgJaiYVRNHcqthFvyuycXmIVfK4/Y+6RxPxUnz0
bsx/+0l9pCuFZymCDB2mR/h+cLbkOfEgF+tk2XHzAimqXnqKGIXKlQlssPAVtXLrOzYfrsRdeqiY
PlFume/XRzZ2+5xohXIHyvhG6Diak/1NUkJl1g928ymPGYT9sBMqInQZIujVWIbz6hsE+cGQ1E0F
83QBFqSsipr7sUj9wsJ1vG4DXXHs8PceAjPkzGj44CsVmm/twrP1xtAoB8oSG0Pn5eaGiNS3erq1
oPOY4IiQ0c2+LTotQ/IH+0xXRCjyiqLb6Uv9OOxPEG4wellQ8E3S2HZSU2wiYs/6rVFnzIgMdyH+
rQfG64w/6FCuZN26AMNmUTgnOk8GKPzbOkLqZdEiWaRvqtdbkoj/KN4FwZKKYD+69YwD4mOJyqXs
Y9hQUWgjdpTg0SvXAyf95DyFvDYXMthNzn1Via/xd+upFlVyhe+3Mb91KYNWwIX2o6mlUoQaesSB
0RKRxSy38+msHKT1y5TDYWsHenzAL9XEEUH+dsmNC776yj2/PyqhP0sQjn3xYk+X98pePWnqmTur
V9F244ptcF53GhbkVXJPlL7dvUl8UgMrARPt5YCEB8qVcUYNRuUrToUODVgjGwPpntjHI+DO1qtT
QfMQHl66n7ukxX4AmSUGnObK+MyoLFdgJlyKMryfndiBqIQg5GPMn1mJrpREbVb0A+rlLWRBa25V
Dbtx3d9RrTodfWsMTRHVMhc6HVogtoYsAgoEbF92O5X/VgRE19A137HEckOi0TLrQKiubhNuH3PA
/242P75x/I1+p9s0nDguj5BJiIXdrEatNCJQJJqSsHfbEijuliVJEZnxS33uWxB0C1eI8+KjJLmh
hQ4KQng/beAps3xuwcykWHFV8EazxJ8gqGXShb7dTkd/7bw3kqwcTgWZFAdrYmf9b7bhKtyJ5OTB
twq6Lv4ULU7K4rkyhd0n2qp+oLIOGjd4ki+WG4FVvd8Cwk8hzQEpOqpRhk55QsvrOIeGc5RdD+cr
ZWrvml9BlTW6ZjKKQ82uytffntiOyBkVQ5WXMw/Y9kBj6EoWnKpmvEFaJ0Vu/jTaIkzguELnz0Of
SC6/k5S1SGdN7ccq4aU72meCVW15Dzz52szXOkxNnakfHkJQY82ouNnB1cQVvxGt2So9AO89NC7P
AKMpBr/GkbSqQqbO9pvD3D/PPcsiieHVH9qiAT0XncdWuqocRk2BmRlyf4g74SZ2UhGR6khvpmL+
GOal0ZAzP1vtFAj7fKc38P6rE6VesEXXjKPEgTEAiB93EA2dEaMN+Vo8cA816/7mX6847nU9I5iR
RoDOz662nrv3ScwM15d9hGrdAlbZ65aIKCOm0KgGfvkn46LCK81d6njQplsF2N3LzmCWGz9hfCpx
2r5tvg1s1NNLTKluDK+aQwbR1+L9CbWxgk0++LG337TEEbiFieJhKGTUKksBL+0b4V/ZRhwvMUpy
nywxG+mAjPefOxNdCJtg7hYYXZTS4lb7hFiSveWZ2jtFYShAGCLwj0Awt79Q8yIhmmMg/PjmM/3Y
RYxwrlkRqekW0jIx5u4dOMQJ6PHXlDjec2mmoVNbTFJ3srcNhK7/EQF168FmUuRi7HencaUjOAmV
yLY40PMWapY5rni+u4uqVg2FJeyEGaRHPcdktYgp2B/22IN7DXysA4+EmkNsrDgjHSjbgXkWwQjK
DvJfsZtsKsFUntcM6Dv8+LbuEuq5PV7Od22pqyjAiyDerMGXTxPAQikDqkLKf1A0c+G6LPHU4jPG
hT8XlLJv1FY8KnI5IWBIotBTsX/qD7XWsywuHTS3ccXdczzou1LgR9a7DRIhugD8OWGgaE1ccSSf
SYnCuKrroWyrAo5vZuAsxKTcUuC+TLSDK2De2Y+F8FCJqlshG7dUZpZ8CeceDqNci86PmaCEDcZS
hFRVvsUB4wCO2tU6HWTnnjlk/ieRJc9fNY9RZmPLD8/kuFRbSG+HjD9NBIaaUY6hvbe+cxh5Zv+K
nO72Y3LDJEC4Dk5xYGEbEnIDwNtT41hHRaGNIlYp4aSV8k5g1UquLy9SBhBXibRCiyf6mL6kqCln
MxXoz19bKnJjso5mDwKSxDTATQPDA54pYO4CSuJnhQdk9QzEVkl6Jhp2eDjN0gEzWsO6In8Lbq18
SOmL/R1zaS8pbc3LPYwB9kmR8TTMEIKphd6RBW8K+MnnsSb8RV8EHOM5PMbV3jMUCEUGjDWqV7hv
vmtI4c4Rd+R0F4ZzgX79cRKdAL6GhuIF0BiAgvruVQ53WrVEb0gAKSOBjNXJV5feIq/1C4DKYuCv
M/+V/axIJvbUftZKDYMyIzPz3mRKxCkDyS3BxFjkGiyP7MbhkmolzEYCdSE8sfwRRYzn/W1c74A0
qDdnAVekJXzKHfFGxottb74x1us6HNBNFmMla3lvo5jjY+RoDD++06Vt7O8WKOOHjdveZusSaLy1
DyeQQHh0ggpQgupEXlA9aQKSgqMRwOEnXht5zxeI8lQBBHDxpl70dk3LQESosUnaZUU7k4UdSYo+
K25VHUdtQwOH3ZnCAhzKm1WYLhPyr6JKl1CvHu2pgv6fFyGwxeqBizSTheBaMRworw3BnrraMzNz
cXmjKllo4aftX/3fGW1WFYvNY2NpibrxqAx0qwQrReABSvBis7AWFkZyzAPENi6bdKJDgTwiEPBQ
l5T+WdnefWfQY92g2lu2BShdof5NvLceOMxrFCMALAjQSZGoeLUB0zGPEAZStSpLvPAgwIlXXYqa
H/7+XkfpWkkvtAzEZaeBXKnNRkC+wLp5J4bm+2Fse3ZvwxQseoOcoWKLpP4vf83zqoqBltnp/VlY
qHxUPJEoHL4d69ZGdYOH5EbiWBsTR7c7xZ6ClQd72HXad3BDsl1yb/VYWBZxKkba2sXTwHueW9vx
pxPerRs8iFX2imFpR1es0FHW3DJkcUVi6LiJ8txla6PpC8fLoar1LV3E79yyBGlPOzP8hbUWxdHF
nVBo8+hvTlYYXoxZMDmTBWRqVlWtCvT9z0DiqALtYoXM8vZEKdx+XO7AgdOzV3NPT0UFbuDZwPi2
SSxMcog7cecOpL4PQeXLfCWKeaqM+m9Pe5J+43VZiU7RgBXMN5T7Hcm/sHKC8Lm49vGJhlnQlbK4
p4+VVTeAC6iZvSFaH6I00tdwN+gThyr9BsuZqkbhkLtIUoHv9pJzWwD4UUaK52rEf6qjTBt17m2r
s09nYPWBfUjediquknmaJX70zi0liFDi5wSPCQqYoAyss+z/h5pn2KPSdQFbEt1+iOhTE7xPhVho
XbSsHcHHi8pwU9oyd0F7U9/PpXMBYJWmUZZX6802kLHrutwkooVGnRpBtjWV9G/U5ebTfHchbuRg
OnIZIl2izgfCA4w/J4Ia/Ff2q30aBZGExc3go3oPtvDjBWrlHN+8kYBm6yHNmIJysdyar1MlXhSZ
QCnbJs9UkIeCOaBcxoWuQ4gBE8siFyA0XED0kWVB5HmnKnk68XWEux+yvE/F7qOlNPmMYgWgKe4o
60li/+3e/+qBHg9Eg+3klcjTbuwTmvC+vipsvOEG8DplZ9hOKtxgiEJLNb4arZDv4GN4XC9s2VU6
0VJxqHOi/tN4Iy02BC0Of6GnBNGdIA38w79hpt/+vnSwX8fjUMYvYT5ZLWo0kY9kKYyaXfufNdJp
77pvOBCwZ0SOtccUzQgDTHFkkE8ltEEvTR9DaW+LBrhsnktSd73duYY04a+HpKdvAnngRQjbkr1r
gLFNqD1YfeTOuZxSeHaSSkwnWBT7tlnnhGyUpyAm+fTdC8kB/ywoz3at3HLacA9k8zdRSFbrQP8d
Mdbuvv3OchzWh1XbCR0NOC8PL22ccbN4tbb8lKLZZEY/ba7Zc+A0JuygsF6e72X6PRDVE/HdW/5A
tpee7hwI/1uIFWEi0Qnw7blSwyWTV2WCkp+NlIVIuQFfVvceUsF2SK64ojOt5PD6hacWhChg18ef
yxJ2Fsuk8BH5evPjRj7wAxfb9Td0pELfNd3CTofumdw6BNLp3jZCKJGka/oK9xI9D2Fjikh2aZcK
tf2r2DvvW6RiQfKzz4uslm5TY9CXFUikDwYXwiWyyDo10T2N66OCemKSPyRhrWKhg9YNodcgXZ2t
MH8EFwE9XkGMrlk6mWir/PqzGvbYLs9UgP86gJmMzfwQDXa16RqzupyZzTW1CNSPsuf8gAqPc/zb
q1fnrrvXZ5djTy5iQ7n4p5S2UPgerbeVSFNYCcKhWX/14yJSv3mdBQ+8K2b2Gc9FWZkRiDj/teHG
vnwcDmi5y6OCqG8vLHk1rMcB+UvmNkEFzaV0qOYWKSHq0ob0570yrePc39YnrfLV4nBHD2xpN/oG
xAzgzy/XLbIMeoF1I/g0mk6NYfYFaROvA0UooFnYos5IMTStXnOJv3BKQSVhs0Zml4zcbRjTnJZG
od3PwtN3iQ8x0u+xbjVk6pN21PGmhksHS01/wIz7tJBlo9cd2fo79g/l6/+XaG+zf8f6iX8Z0EFv
+/A0FEydp/QhyjddOC9ucqMdhXthDy/e9bKNSr5+hokjEs5rrNkmdajCUBfxIMS6sZrDH74TYG6F
mIjZkiVyRhGAjw8wzttjw9hylrSiqdTYU+VbNILAJk30wlfOo2blSFLwsC+qMTZNYtODWlvw9Isr
rsMQQCOZ9OGdx3Dq3n5CBdTLUFmQLvdNZ+X9ZXipCb+5nDV08N+3KhuzOZ6TPGnp06XT2a0nDB/P
Uhubv8Tgmy1cC3Hc6vCIOvmv+GgGe3U/WoQ7vhQgmJMFiC1RqruyNNWkZRb2lFGBoBzaMKaHC9Js
VuM8X9jGHzppWL4t4gVMUuv1SM44sbwYeFjHGhmib4xQByjEutqJunTyVyJZdMybEfotZceiSv98
2BGUiMbL7WUVXkWShHSExAHPiPLSEOx7C2ypNULCuFBAnk+hmFxG3cUYciNjUUwBEjm1P7e2RGho
bzNI/naN0wCGyFSy19M8UutBKOjnECQP9C8qY2hMHh0yg6x4gVP9/km3G1upTNr0Ap1l5mdCtBn+
Syke2phFUtCjem3sTy4nzWwPWWvjQocDftDyRDdjkdsZGfQ1aWCHgk++NbRz8CZPxw5d7DcTXkI5
smUWrfAZWwgzYYdJJBltIUetyQDRC5ET3ev/+dKn94PVnVpYOwM4GP276V/c/2vEBpRii6tiwHj/
l3gHGxv7xa8+K/dqcO84qVdqt1jArpI3cFYpMxpWwtZ+iM31XhKsMM9H4sfPwNXAxu/8mOqjF6E+
O5VxIaNvvzHyUzRrUv6h+WyTRZAAGqs8Z1fZl+D6d8/tFdbs2oqeR676L5/GmyymLs8Qtqd53VgF
qmU7qXVi6tuuSPbKVxRUIQUR3JP12hcGR28m1MxeC2MudCLjrp48KGOXBz7jN0pUZGS4JUejV1K0
8TRJzdb0OKBeu9VbfEje7nJNW6tzqTsfhAT/TrueCkImPwWyVPx/2j1/nJdOPp7ij6DOKMnZoLSe
Vx+smeCGjk+54KKSue7gzaWscLb4esVK07tc2Rt1C6BifDDske69s4lGGg6ekuHUAQpHyOTOzXY6
1+cJ9rwKyppNXuSpgfoCd6aPMRrHEsE17e9qT/0s3GhhUNDdsHmtfvHPoSUlTbLRWW0TmX9/Jj+z
+1b731E8n5U7sfBMJ7IYcuDjAkOT+SE0ymsetdmlN8wJZUuIAjWU6OKQuJoytHD0lnAmncFWkaX/
+ULpVZBoutuGuegFO4JQk186Fg3qKpqRJXlPkxjz9uShj3qO6biEkYWO3id9uWlHIBSlZh5iDdcE
vGy83LfiHJhBsrf/7O34Ju+hA/J0p5VzIrl0ITn3FNUGiSQi0FSETNM3zwl+KwoIyvL8QN8rWxAB
ihJ4/++lcamG4VO9guuJpp6u6eb99xvhMQ9U0rNheoEVvrv3Jly7RWGtJehSMPBIh0PhFDVoJGgP
uLX8GWUHhyOSiLk/VpWljzm3cEesQ0pV4ffYAs774imqZh0jTympscOzbQOC+UM2HlEtumX4exIk
pQEIDUk2Vgi4Zu+O2cO/gha0117w7nl5zzzlzXg/JRvapncH9MmE+NyJAPgAb2Ll8+5XUoDarPG1
W9mpY8fpXhzoEfDE2hbKdMj4B2WPW1/MIsAnrTHvdY59loM4y5mu42pjp52UY7PZx641XCD+PPQo
/p9SvpUOEtyr4Y4sYH+0RozQJDkDwc7XFIcqrgh5dHmFvyTmthlhsFQjvFzQFtY7dhDPki6VnGm1
e87+owmQh+ebfKgoCvR7JSm65Q8M7DBduxvGDLjPQu4zXPpaIw9bbiWaRd+48OIVe35XhlrA6QfC
YaIjfxvypFXox7rzbXISzUx1Ryab7GZtDCFcqYzEaUmmVzYx7Rlyw59k+2h7js1Dv6QBXTchZJDA
TY9RNTVGoR/SVVqkvI/yg2NIYcyCgHhqaUAd6RIoTFzmsUYHznAK7SZmnzd7TEUMvspboYiiGlpO
lWKKuqqaQhxzu7W/heZhwQ4t/PaE1E3cjBuALoUybFNlGmxVeHymY5xdG/79OsysD+340HvczeQp
p5+YjcN/Ixc/9OivToZzf3pCiOSRXlYlWuGqh9dgGP0ljNDDrsiNWSNrtOGAaAgK36YPYa7sooL4
bFLRT4IPsby+srg/m7C/4ThtbQmj6QN/QkCU5TK3tkGKbre5TF8WEBb7VH4kveZ5ehZp2T8HLsKN
L03aV8jzQP0XMRe2iT0+0fRLQjoRsyTqwVM9d9VKWS5FIMY//rZ38nwroneup0fKmykI9TcuMgrb
6rzFwXlTNcwmESukoheQcD4PaiPwrNJEg6L6TDNMJD2SVzlk58gTQROwVSTZ7lDu7nskv4l5TMkH
KdPRTsxl9uyh99JC06RxPmCcGTNIwQxIXjfdxBeMle4UJND8rNJ6ZzQdw+/uwWMbldtZL72aml8b
rXBZO802iiL/7qyfy/0cuD7NSejeTbSctT7En8X5gMfVvWaVOygdJZ12KEuwn8nx+8N0yvNZWZQv
wbWkrqFwSA6tOy4LDHVahFHib7XPq1mA/cWXuHxIVv1bSx7/5AQWCXOSsxLrxuL4CoWYANnLBM/8
YqjULpKW0MprRyRHzG5Kpa94lyC1v8qWNiXDL3oFyqYzKulJ0LJIMVMuCvKvPgwnhIW5VUFihIZr
f4y/6rK2H8nuz29ohMxN5vUtFSYUsH2FobZRifwQ9FyylTt4oLnClQr0yZ3lFU4B/wDCNtIZot4d
ZBwOm6E7XKF+I72qojCXK28QHbDOiNqOjRL+3QFJj/jZ65O1jsPvyZdaZJwResYoPOEyVJfkd/JY
M+g/tvJ7DbmlvRQxIeVf5u6e8v8c+vWtL9tAutnXstLMdKs71HLJKuk8RGUpWRp1qd3QD2EdfDPo
d+JQhBINQlC1vmvq+RfmsWzHQs/z3UU1qcHhymGzM+fGlGOKJ95jG5HGZkZe5o53lR27G9ij6ONF
OjKYo0EAiElziIF3tFTJSWqHsw4VChWhKx8UA3/znHE2f+w2uK1OQZ55OtBo6cH60cN4VkcVj4tG
mZIdgnfMJAs4wQrI+TRmR2JIwT9ocFRDiOMB9syL0dguS8SO73r7nI2v9oViWlg4IC0sq7lBQ6mz
JUzRDTeWpTE+eOTJcebqWZliwV4ihZSD318/Wd7sxP9QRGMUYGl/h1XnASrGH8mTb70fW9S8SLcr
j1lRRgArKvfhyiZeBMXONFX0zc1TT2zjbXZg6GhZaD/i5KjjpMj8PIxf4qRWVlmkxsrLAnVm9q4F
j3bQ0t9o9l+rXcCIpsxaxTF/WnjfH0/NmnR5xIQWICZpKvnJ3HDaKO/Ty5svNxU3ncXde1eWYYa5
GLPw99YFD+EsEdrkuDioI91LvHkm3oawvkajtUGeKOg6dTSPQAmN6X/HKiAaAelAowQ5xu5Q8Z2R
rmvnb1iWtMvyym6w8MJU4NQQzi4hMDICQ29l7sRzvqRFHQ2c85GWYhUP/4l2YMYnuVHFc0O6JrvJ
Q88VSPmj+I9DIFCS1AK9ayZMRFAry/d0mBhzulRwksVityK8A3DeYzqNFnZ271o6d78mZLSke40U
0pdS3E3Zh4aHf4ODVICePc7NWiPWEjYo5zJ9RGvj/JB51wb2nfrsAtL6Z6OmIXizc8MFSjP3kPej
F5Z1BY/YlTQ0TOTNoDDudTOXQXkarK/o31U7Gngprq42iN8beNlbaYiivQRZHnQwYxBVTUtIfYyq
AsGgJtBWiMffwYvZv3kzeJej0S4CAZE9eLuDzXa4Rz9ebEYN9actELpPk2f5mlkeCcyJBQV+0bkZ
AW670XrpPRJstq8ZhTMhF2/h+Sp4EKqkj3zk+KsItMwzsAsDV7DuO5bA5wBN4cm9/AD7kp4pDYJR
LMMYL8Uif/afzvlqj1iSeZQsd/dojbA1qAmCsNWlItdzYR2VJxNhJd83t9r4u1W3+V00uFQNLzaL
91V9wxJtHNAoJqF+99eJ2B/XYsfs+Qvot040c5/0YZRI5H6OORKHqzYqV+r1Sc52mYgaIa/p9TKd
+QhihE4jjVTRMbZgvCRMP/o/NoMGDiSPpBB2sulv9KUq5/TlGYqP/1WT5tyNL3eDnagT2D1fAGwD
TfCX2ZXsUfesQ8zl64aWgWaX8kdBcyNYjZuSPB4RvCfDwALKYdrsoxkNRsXYXF0YmQt6hb8Z3BHL
jcO3oVdEFSFulYOnOibV1wXnkLWpwECOoNsE7r5+4I5itZOlKoNEdFu27l6b4O8B7XkLXtY7qRFJ
/QNVHVDBx73x66DVz0sx19EGIiv+e18quL/O4jNvj3E2lYYie7+Ejj2dhKYTh5e18OQAwTinV3El
dssCewXwAAnXgXZM/U4VV52WrILJhGEmAG09bturDt/t4disqr3dD7iA2uHcn+7EP1c556ntbG5y
6Jr1Qqaf5UsukfNfCESb607HCpEQNwuObJ57G3HmajTGqpnDlvm7j5eaKqNkquJllFEna9oQJgcd
bMhfEoMjKmxh31DCAm1io8ePrbUTTVHVLJbaoEA3GquIE4a0E+D1/JPkBTGKer7CUa4TxfAVkfb9
5M8vyvJTEf7rQ+X37qnm3kZtl0T4cBjY9YJaEpC6/z5vHPOXmJxgNOYMJ3A4VF9lAIp5/d66v4gi
++Lsr+Pq8yvSJrZgyPXbjqOJ47uPOHGlJx3ltaapHiL+jDkXhuedUWFRVbcSBbtK4iHOpIaKoc3L
h7n/4Phkifvtvfkjzq/uq1kOspTliehZjE+2WhiU6qQrzBFBZPZhsSbzHUmHgwTqlyRW1l6wRVAU
Ve+KYZGpC6PPamX+Kib7kZEBuL1aWD2UFewXLDwV6zWvsaUb7BUmvTEWTYrbMy6JFHbNTGxQQ54k
YEU5DgwGUxM3C+sxrXxFNPbQv0lzcD56oE353ossG5mjj0laSYfIrGpa278oyzeI/WvgzeiPdCco
m5bsM1ahb8H8VYDn192nrgnd6aLI1YGYN9zj0GChMj9BH/sZVy4nERAMJoaNJfG/mLLnSWizzvgx
ZXoZwuna98x1wq32MpTFsCRi64hp109lcK7JQRQoS1eYQtkhCtmGyB01o+C8agaik0JcC2hXU8at
+9RBmaWpyYtFfj11nDgXqgAVzSYli3TpmQ/dBsIoXg6L3E/97lmjQPKi+xScE+id8b8q+1Rwyuwz
JrQpn2LJCAMXcC6Cge2IPZTiwNH90qN/3H99DCBukqoD+j2asgzNJYsVUoEvcUiHCfEcjpdpJFdL
6RzN9O5GTwIuoLvpdxWEII9OU1Gi61MH9M3vOCqWcKutmIcHezFT9bTOU5tjyp5pNKcvBYcn8+8I
GZ6Laqln3bRFL5R3s9w3DsjyB6DMLZDFVmt1Iipmt6DBhRCp9+aWRL3zhNQMRlxnN4VzDoh9aiOt
nlTelKpJY0URL15ByqZYcInv19DQ3f+ldcZQ/WiK1R5QDKU0yRFN7L1fty7ffG2z+GCg3YdJ2//j
fdLead1GvwjCdrLny2CWQR1MgikkyOW+JfH15GF16A3mIIBvs9OwyH/M4O6pc5vFd0SCb4d9o1g/
KtS+OUFrmzdjr9+5xB+icuLXJbYoO1iwR4XyigLdVgfkd4RUpid5305luYq9kCw8yIiNbd/a2pQ0
8kKfnuFi0v0rA3fJ0/9nnet79wqVwU2mRNiRkhIZXtPuPsoWELT3w7mEky8OjsCbPiA8NEl8SaDe
ob5WyQa3PbRA7N5zO4TiIi7dQ0PH9N9BX8O+BrUFzl+KqAs689oMofvsrMqhX2bxhT7370tuzkpd
6tQT+OzSXrLnG/SQY91K5i73fat7kfBNWxrPRzYZ2XOGGU2c6979EScTx38PwoW3WZ7XNjcFIoV9
GjLiGU0n1395lSEYuGo/AX9Pfqs+MXvzT+NHLny6kkcbmZswEffFs2fdj21KjCpuhD4F9XWnV3zR
w5R8y6WatAS1c8lV9h+MGfSqO6hdm8EDXJcDZ6JRaCZt7p+1ezhzWTgXBNtQyzAcsMNjWUSlOT3f
9xXAu0aTJ9015SOT2xkj5+3d6Xf+GWeWIa6bw6PTKJGnQXxvwf9Hdkm1EBVYrycI7yJR89qaIqk2
mdV3akKT9UOhD1RWfuDYRgRx4MbAeVOgISVMXELVohAp5yL9abuv3rMc5SEgl4Ya3KY/+FrRN+Lb
/f5rXh3Hb4tlYFrataejhh/8XJYBEI4P7ClvPGF/hGm1gyWAQqxtPAmpGqWkjFqBc90aNQP4M1uv
kh73VRJ6Dp4L15ddusbEag7YZcqtKXbH0Ga8pEcBfHJMeoqwo76afLK9S0KSAdxmTLoE+MpyBlMI
NHolhnY0qHAHSw6NUS+AM7/aRrwsBFZf+59rLW/JeMLipTHnOnDpgIBFVox6fG8bJzMon0Zkn4zt
AB9k9bYcJFtR+IpXI2r54h3YY8cq1bySjQ18/oMZDfaLDiOneOSWyUGus7Z0uMLNm53HtDRbuQLP
/Xl9V8qrPpp4GAgZAqf4SMrZuoOiZSDzeP0kwPG4lvS3gehOW0wEaKZazhZZrjpt0VXKhe9TOvTa
Il8B8yIHjNMF5GkNyqXQRAVJ4HJv5BFTwH631aZQpGj3XYHgkd5KALB70gHH3g1sDgAR8vrqmO/1
GqboOvDoL8jaOMKhAU2DbsqqJyYwOVa+ToutiGdadjwSbNiL5hFHuaxGzDf0zmRmWmKL87c90f62
/vzYM+1zgy40QiNZlvdnc6hzCwp3THJ8zW4wgjxsznlonKZchw/uh8vdMuIl+a3RWoGnnlFbEudA
G+/AlwB3JXFVzv6bqqclAbkyo0Stjmj20Djv89szOiIPjhAX4XurCYey8DRQWi3ttY3CNFNU0d2B
trzskNW7XoAZPaPSZ+9IKGt363h7Gq9Tc8Qt9CARFLtt0TWYRSfQo1+CrS1421ZxBlFY8fiZkhx3
DjMedc66pbyq7I0PPHqQUCAkz+cZVCUPLVC0Ef9tTp/VX8Ao+c/qzXKYFJsXDBiNFBT0wzOxJFGj
3120u+Xr6XgzRMCDV4IpfDtGkYL+H7clxSc0PTkdhK6QWCo/8P9EdtpdKaTlkGO1NODRDtZEx7BS
Vsz2P4EWOrUiZpLwSN6W4UvqI0OWmPPnuttiHDMM4JSSIwI4IMGS3FiP1U+emSAlLKwFFB7Ehk5z
7421goiAVrgB4gxgGFodEZq/LDjoajup4OF/Y1mAuz8Dp6cjteJGThWdCWN7yhW3hCpcAo4NhICH
gIm0DcXjWVLPjdjoPavSlrtQHdBQfnzsTDJU7oEa7/eFtFVtfkQamkcQ9eU1sVQY2WQ0TR1/qDgH
yAII/JBcaxve/D7cB1kTolyvB5o7ZtcBNI2AH1P0xgrE3XZnpLby74S1/HH9f9GDU49OEIu18aqJ
B5qZkKIN6KFjuyknhCQM8x65mApJ3hybCaX0skEkYS2Oh00axnIfYfjEN7Sj1xbuMEXTP77do9bE
fX/1lI/eCHHKAxNNYJjrsybcQJe/pOWs/CMkuv1RmYTLEtONBHK8RbvP9uUK1jjtPy0K4RYk4F4g
Qbu/5leMNzkc+aeIsQ8QTNG/uiFmCB4tjQH6S3II4KpxJhoclAXdiVtZJEPdbFuyI3hzlWYuyaIk
U0rZ/9Cne+zbqYKs8Ts0GeBY4HtGNF0UjnNO6IjdAQNgVGOyAvfgvGeaiwaPxWp9DZGX/TwaVx3h
8vtExQrioDjYIa2LNEVaV2J0YAb6VHwwFQREYi9/3FsPH9AaT2dZ8laBBUTvr26aSlijUARI2+3a
AB4vjiWktadsfJS3FCNQ0gtAkC39S1OZCb1I70yiN+YZG5qLRH5DiHmUjtxksIhaVBlBNmyS57Xf
AU5j/G3gMOy6IZnZtvI9lVl+tTV3q+xLdDoE9so0MWDNCbgnQFU0z0u1V543vm3GPjX3z48SaEgj
wJAmnNgINWgMKvZNVjsyosOx88XM6RdFBJ9SQAVlqEBas9oveaS+4SMZL96+oYUV47ER1fwmFB+o
0f/pveScxaM/Kqc3KD1Jw05ZXiVs2YTJXzPc7P5GRjxk3TbGL/anZLzDTXVo9LgQanld89YBFFTL
dTj2e7yL6R0aDSn2nA+MJChP+OsUYLrHsnX7w7LVJT0QsWPnpdwaicb8BbnoTF5NpdaAInEqXsJy
m2apqkKA1nkzYy8Kj0lOEdDUlAYQAP4b2Xay17qCJ7r8WK33ULVcTibwVMCH3ks7rtRfMKxPeVyg
FZdLsO3VsrtpQHa1snCibPnX1G1bf/4DISpQ/0AGzfA0TvfwhifxwU4DZ/H6xGN7xM/whfWwsVfW
3oXjfSQbcy4Nzofh3KESEW+4aLi6JX9R/NmDNgJ6JYrpfsb2X0FdG6PQCqCarWNRPxJCFkL5NA0U
cZFwIUTp9EvYYRyJuURHSDwrssi2olzPnWXpeyhQDcLC8YfBvzaS8A94MP0wGTRsr56ExGqBGLIk
CdlfhJn/4jyiAnQY9OUiEz4KYtq8FYR+Lf4m/6LHGAm9HZjL8BQXenGA8XMhtyixUOZlWKfbC9ua
pbZTjmCMXWmWQn7g09S4Abivcttgm8z5G3UzVuHXK/Vf92VCEfi429LeZ8UDBG70B/vvIkfgWof6
c3a1DJ4ZZZBX0bEXAhKCgtnONThEVO22HDlf4VvFSnTYQGckPZzZ+4c51iwakeNJ0lLgs25cAAxK
GaVfeR9sEhOVdCo3MA2qoNs88ftCfhClU0UlX/9FHxtqtMM+UcJCiTaAoPYy6wGLpp28oY+hMwWW
OY03QhM6/2hwnAnsWHAKA4x0uzhBRP0bmeWDApwkwyFe3cMtpwZf8sEFvJMVaZtvwT3H9yPT+HJ1
grmMJjd6BnvABP1P/cl0CFVGptNf2YPAnTEVCUzcwEnQ5knIa//gMWvBHanCgRhnON6Dmbk2DrQF
lmFyOo7nXctA9aydiokOrKq6dMy6kTNaD/YEx8l6bjjJQS5QmoJmleNAy4jxwD+FmGtD5p+8SrSR
vd4DdPqxxsO6bZOxweeRlefHR31v1x0BRG19xugBCrVxHIWWkOvOknnv+L+yYB/JmcTzNLlWSiCc
eA4o4WWyn+t6N62ZLFSLjw652LDKqpKaKw5zP3ZKbTiPq/l3MpFTagyQri2Xu6hmEHiOq0NWjfkU
JgIvRE7J9llylzTUqXGX6JlrLMea8qopG8EfCf17Bw75yT1U83sN1le7O4I4ZxSepENuqIp7uKZa
A3VlQ2WImwvlbJMu9ArNTf6mhh01N46ziuGFAVjrBBcRiyG09zz4CyFDwFME/52ogUiYxufL2KTY
g7hAM7jnFdvxxaN92EV7TxYgU/Vqg+P8pE8I+9JbBtTEfwG/I1h72wKNhNBWrqFQtT3TPmjYNN1Y
xH66uLe/14egoIb65P2KDr+0gF48zusnHQHJNiUHrKwkky0Tbv96b48m8JhvVm9KTfj5yqs39LDw
FQfnHIuXoZBJoKD+k8WdG2pzxBS0E/yq+/y4/WFREN25bvDEfs9jeaE+8z+8HkFSu7nUNlMqdRHE
n2LawXwbcTQM7D1XydZaT30coIds9TICIW0C7IP9f9E93QOBuBLzDzZZQ8kaw2wh/AEh3sCQS3L9
EmkIE7WfpbaZ3gre2aDT5GLnUyVb4s/92wJCEqWxaXHRE4Oj4Ko7QWRQFuVRAzAZqdtdYYbNkv1u
ZaQulzn2Cg9u7hM19P3NvS+O1c+wS3H2TZ47tmGwYq87Xt53ceVSrjOpMyvcuxBOorKFnV2fwuyR
VSNoLUPEnQbzBXDtNnIBmYifTDAP4418I8au3rX2PktgiDiCbkE7YTpisMKHxH0qyC2TTV6yYqEx
sM3iFCFup54aIZ3+fUjK6z86PB06Qqw9Y1vwN5TczKsTqhLIP04/Z2nOUnbfSSJrztR6H67ruITO
xt+8oE44glv2zj+AiWOX12eEAWevLHygKufkLvq7K2i+Ihk5v5CF02+0tRU7AgvbNYqGAJdK5ONQ
sF0h45FyHSp+oDCNaNU2uZ/hSaob6urxfg8kQbPuoqmTo1ebcSzA/Aeogv+SuNHqBz/bV4Ywc19T
u36tRlj80ZvitUDu+53fvYf/hSEPo6U4IDbphEhk59qzuUlSgsLcqmQ2B2eRXnO2jVXabStszQsf
Q62ZIITnWsleTz96JpZplXCbWhsE4pB1f06VhART7/1871v8Qt3qdE94cbCoV585sdnIg3awDjsk
a2D1BQZvTMr52pOI3+FfmE0FAsGj5zFAOZp0EOhWSQnYeGhLzd/dqlOJnzbrUR+FtuchEoTheU+J
tp4Cq+rWU9Ymh2n6pb98uotUNauY/rhvayqVmNynBHcZYsDXTuzwR3bK0RXHnTGbw4NT9x7adZa4
iOMtSIkrzjM5bRuWG7/G2hG1R0/gN6Mzhc0tG2yW8i+5brYP2qt02RnwD62dFEbKj7fKSLIx4McB
opXRUIGNpi4Veyaxkv7c5DFIRaZVs9qKUD51+BLRLGRelRRpcY485+7HZdbVmYfOz8Y462/4YwUH
2fX9dY5NrLRCbIUOQa++/TbysLuX8eD0ij7ZfUcuM/Hiks1Q7ZOTTOa5r7vkG5eYVDVK5wS1yZS9
MZ0t36tLU4Qh9d88Xu0tx+B8mv1NvRl7bM47+QKXjea+5l5orZ1D2oxg0yyV/TstvI7YP1k2KX7H
/Nf6u/qBU/Kv889p3Tw9eLPt3vHkK3KNECmfJb5cSvTxRuEPUGAHlOl+rWoNmWwLNMn4/9hpV1t8
x7D7PsYXzbTDG9tRrjubBn0wDeKT23dZ9LfgwvVcA5fbB3RnjIMWqgmJRsqPLUx5Jc489fLiplq+
wiXNldHSWRF8CvtOhTLB10MgtXFlXSEd+njZwIvI31ejJKoghzb9QMWVeyYbUbuL8WX5gO0oStgF
j9A5Zi0chTCeEqeX0KLUZ1ZBmaxQItrd9lHg373/z3sT3dOCoGye8LsKe5U9f/wQotYrNE7Nn3xr
82+esG6zjJQFJu8ol6ti36pZxFvWycvyKW11aDE3v3uJIaeXTpInu50oUmCW2izwf2ZpZKg+zQKd
RPT9wx7Ao4DFRyef8jKztGRoIfKxKL8/2W/Qb0O+qFZUOvrN9UCgbS13BHFibx+AoONGhwtGKQXe
Gwv9x37A+mUwQAg+sgt95Jt/hAnI6xSfdAWWnbD/BEpiLlZsKXlZeIiaagEqPXT9MhCh1Abhwry/
ovp4XCuFGVSkSdBqE9P8cvl6My8HI/hpE/E0SD834sTkyk7ScYemmHeNtx/1oKU7F8P+hfoishfo
X7K+xFckTP8Btj5MEAZCUv3opBybnyVAkCmiC3Jkm0SLrD4eeXxjps6Mp94euCakgLWEMyQ3tYFS
T4h/JZuAfZvcp6fWYRyglQak0JPxoHYUZzMQcqZjyCWRhMiqdyMBQcoZLyGC9rVF5w+3fDovE5CE
eCURFTG56rP1EC7lyFOu8dW2aEh9shnY3644xLx7iTNv5zIH2MLsOVxhWWX4V6aveiTBTDCcpgTO
vUhQU48sg1feUnuQ9dWT5ABc8gG7CbLp3k7f+Gs0A5c7sPjTEy3Tgrq4mp1J3tUdcv37RU8sDFXT
5V56USXcXiWEN920wFS8VxSHo2KA5sx/Ld/drVRUyNhrI0gzTENF49sSi+dCTSObdXt7o0gGzEk7
MJVcMMd82cRWTf+nEgxyP2O7Yl74oSWXhyJHkcPbGF9Z0V0MhFjKqAi5YIxSUYnWHylkeRRZNfsc
zKp4JM8YbdL9hnJwopdsHQraDwOqRvqxIu2aNViGj5KaZ1VzuwhgYXgyoEt91++z/GRe7p9gthEb
M8MhnlVjwd5w1Q8/1FstIz4HGAdBXbBjuFkMC5TJ5aiSuAO+K11cTxqaLSCgFI2xOrSZCttHjuqb
uheZE6VmxjX5PJjB2+Y75Gd90l5+f3LscL4KEbP42IhtiEFKj3HCsiJJxDuNJtb8W2VcvVZixgHr
V5Fr4zqXUtDEItcc79DDK6BMWpasDaY0ROC4FYScZz45ChvEBjyNnOuVPgMgeoEYACzWcH8UCyX9
1wzRr3XFvl2o2H7CJ9Vxu0UYnwPGjk8zOzzIVUF0Dt7MS17phNBeFIbIw9G5cqm7EEd+gUwzmRnb
ozg6O9x4PqFiyIcrOTbHrjEQDEV045s/YOVPxuZdNksILoaEqzAFQH67BOjtXOgBe0nW+nlsvrlB
hOFlig8/wqn2rhGRxngD4RA+yyzt47tP1AsOLui8e2MGXkMrdrYt7IrpZ63Ppww9ankMVol1FX0M
hPrsjWdm6EFIWxOoD7NC0U02NFKkTrmKT6KPn+7DoG3ZQTFUa1VhzddV/tPUx6v4RdZRR3PryLSg
PYXASBaW6dW4aGm5BXtzMIDE7oSaTATNasIxQC8/BxV9PpCiscYuEpDxoIhoUO3GtQb0UKTUd1Rw
L41+SbLc745YM2icpACvuVgb/L3XCkxJZbT3tkz8BAII+dPWn5ZOhDrGj3iEUBMEVLAQ18WQX3cv
buecFwyhn75V+btAgFDwQpSGFZpaFq/UJsWG9waazR6Q6e99n8lzhIACMxWO3KDYEB246AG2Vyp3
Mr9NsR91Wa98io+LgMUDquyeTz8nRlmvX2EGVNeP1Zs3+9a7PAXN1gZB79qDoxJ0Ca8mtsYNMppc
MPY+cshx3W1sFKce2JuL2p+GmwX/OoTU3CB98gnVHADzMhu2FigC5u3wFu8eJJxeYbrsJIEbLQbR
aM67YwkpR3KfK+c112b3tTYQZ7cNvfDRhuychK7JGPFfpGqep0ykDPxsk9OEydqSRe5Zgrkn5iL6
IijBt2eAdripEBGYHvgHJGZGVF4oGN/QVe52Zp3CIdUHRN/V0BSONw6C9F6zsJoG3whubwNDp0Lq
cxlNWj3b7D1j8PhtwjbKDn3Yhce1OjY6iK7mMLmi2hNAed/N2SnLet48cKavqyCRh4FjiAPE4oic
9ENaswVlmUhk88o5deffcgt1qz6BzScyE3SwLUTW02xw1pLPkxBKhBqvo6VdZHYqmQEJOiTmGHNN
WNhTlj1lb1oV9IMc6edLoPdqLNPkIMmgdJWCwIZkMvuZr2rZi4LSq72Y/XUtotMde6bGe+Sl4WQm
mYL70J9xOtl98jKOMvZdM4TTIu4CotNRU1qUmVFfg8rE5nEJs/787X3b7vrBAay8yZDADQPMnQTJ
Nbo61lAMv7qs3S1E2a0b32I7PJAAkz2fMadqTQBLYsHdgi31guY6PQaqXiGzIeVZ0Be3dOH/2U/n
7A2UtUFeXDbvsv+qjOamiXH9WbTn3IkCXr9mkrLjtAWHGIrmaN6BPODqHMLpV/Cfvi2cYY7SuAqH
Mhm7mLRGAKpjiu+Bqrd/8Veu9nkDdXAHK1eI7LC/02cUdAceEURTWECvFWi+pSveXoj9b1eLySbC
wQohna1C/NrG5m0GVOvJ2rKR4+WCyvoyVTl7/dUs0UqoJeJbkJFoyQYSGH8ef+244nLihqVSiD14
Ede7oePSPW1E1msF4FIvgUC2DA9v0+hTUpWQPeos1h0FNrB75ctYKQapgWkKYpOegLXeRivoxARH
ZrQ3QODAQYQc8zJi7XB9S4pqiq4D3NKWuNpntHJAlx9YlYVOTeSNHiF+jrrGoNVaRaRGpm/cIxyN
oJg3j0PVuQORraIg01c7dwtqhJOxlDUCD7irET0XwrcghT6gXYOhhrOWA2fIJBNYyMbtZa2MCjXD
rDo9s0+plLW5wEAo8a8XuTI80nPXqhCTNNVkHpAqG2cgDS+m5tz+tQgWM9ZUWK3q54B81icnPPJK
/WhHz9txu1LCxJHh1grssYEdgA1jShfckpUtzHxWE48izrBsMQL7iRQZtJEJVw6O6XyM7VqIzG1j
2EZp2N1DBwXvAQjKWnxBND1WV5xpMl/CaRDEGp1HWBGuwn/nqvFx2e8R5xCAAMrilvFaGXb8pZNq
GNjvwQ0R5w2HEi4Rg4Y9gowHHobNB3Pu2Ma1XXsBLv5A8l8Nix+ojMygIA32cvsZql0bXzNHEPpC
OJ+8lIYbMjSbMwHsv95f40nT1Xa/HpQt9517SFExfKCMv1jw541YNJNNzLT6AiHlnjlQkIlMsAa2
ykdHOhJy7GYyr60N03xzWJiwJIkyNvJg5yPMt/eD7ajPUGeCnBg+ejlbbphVjDo3fzIrNAlr5/St
Jh6VTm94q+rhX8/nDEyPbf+P4FRrqyi1iqoJ3/Um5vKQwAGVoo8ZwEqM2KO05P9mMoxbpDrzJgVP
JfzKyIB8JGV7A5UCq+bcKn/D2JT+3K4afGfcvx3XmauJwgBpqVSXFUS65Fl9QNS4xqeNyRUYbHVD
KMPBGA3f14ihZkXULET/YO5o/gGqAmy7xKTDdp66R9ptzW/rpi9EPC39gWr01g/jBw6hZdOYVqbP
ofRs9zjvr64jNt0XfRAvD/frm9RO/iiUUinh70zqbDSS4lcDeoILvsrgYFg1ukPcezno1wFR5cZn
tyrZSX/z6gciwl4Mt5U1Cp0zfhCxbFm6r3z66vbg3T9ERp3SVadNBsHOPTvSDlBziGjYjBQGV+hI
dCRvcROC+mXwfLIfRs58LEMVYzznvtiDgTr2GZAdWpxIwrc7JOwqk/sKfvgB21XlT6vpwfcEdgzt
1jLs/utuSLPxjx7hskW67L3o/VFL9oK4PHjyHlxOgmdc3d2Me1rmyO6C6g5fjpA1nN3HI8JT4aYr
xJg32ttb0+rwKGJn8ksMNVdCywBuyLiHiomZzOT7m0OYSyVPHFy7YVg5ZRda86KfUwI+/Oz89eEV
tVWOknMO7Yy/WUvmzVlsAC4Au5P+iNbTEvpVbjtrxHDejzlU84Mj3Ut7pPJbl5vo997wEnOb81AN
Xk6AFrtClR9nC0f5louXvSmXx1UDd2RCQrlo/rHu3G82Vlu5ZllZZrCA5mYoMSPR4044EBW1f770
8oUAa+m2yne2TcXCON+XkfaLrwO9+fSZuLQyE4jvRqkC8ARIlhdFmqivXt7K1aR7bQM+BRBonjmh
OiybDzSC4/9jKg0T1JB0j+YGfZyuWp/ZOjhfT9JiNMt5qolcNZfeEurtIlwO3oK1iXU0iaCsCWQg
9Owsc+kZSFJl1TPduDbWkAD3KWOFa37klRZsjkEkgYdq8wVZ52pleEx97HFa/HYlBy4Twa128QLI
y1XWIHFTwlhsCgPHBrAxeLMPR3iBAypeP7wHj5OVH5Bavierts+Zof/xObe+6mLTzPr68pjBnQyv
eGFqZCmeTxr8ugZjWf1ndr1anIzeP3eEBxNoowzZh9b09V+kgLt5z2M5kwmA5AxPQFlQSembvw8E
qw/zqKY6fvIsmxMY9kylGZDIyJlzL9MBc+I1T+F+lcomjDREMyOaHnGKnDOIERaHgTJIZYhd4a4t
n7Rc/6ubdQClwgX8YKtm6RTUw2qm7ozG0ApwDf7FnHbCCIcYh2KJAuE97T3mDKuxdhuiYBobCczx
weLFf0iY3AY/D/gb4DcRge+SjwbVDEAI+vhvrEmxo493CYSGYMw0DzY5lsgMzTiaRjfJSTKJSfkh
VqOIurhWO3ze2Fo3TfPHMTp+SrBy6HwDcT9RdDZO//lqP8nnZ0GGpOUMerJI35yztNA7Ob8gR+He
Xupn8mJzUmQujVruXp03XFQqQShNAA5fSoW2LjZXuBBNwoEmwljALVDjK7Vj812qp90jdA7BxHyg
jS3Spe9JFivgm9j20rx3LuYJ1ig1b2Eaa8tExIBmfPtpLmh/wE+L7cA6++SrQgFVTcDt/pE/jxHZ
46F0Pp4LKoO73d+S1k6jy5/Z+gzYYCihzJEGtpL536/pbDtSMWRvCy5Hn4fCdANaF3l35Wu/bpfQ
B0SQUSlDun7K2H1mQ/dcvUHyUMYPj3WsFP3LA/e8/NrLVOFa/najGjvJFtm0dS6U6oguFEUT3EiZ
/9y6g8xmwpPswoK2K4zRUZFPd/uEcRqwEditlEjYhF+6eZIxxrlEMYG+qxCvbtyC3hVRWtrSIbmk
h/GQ7/m+k+CHwiov/ux0GUhnG80mLZ8vYaTEbcm26LgC126vJ+ZKr+2sCA+Kd4OCkhonyP11XFYF
FuYKIoyjwX1/8i2G9OLH3Ydubmf3eeETqvXcE4Odew9zzD2bw9oNiNKob0gU39RbWISE1B3CdGuo
HpiSNfL/BOUI35gyE2L8IT70kxpUIUJZGxts7euozdVW8f5IAM63YskycNdy5i8LZbAsW4EjBFax
TN43L9MYKKzDOT1ktQzFCR3YTOlOhUz1pngihQQclryFAxkF1lO3ucZfKpeKV4bMgIy0MlGl8WxR
cGRL146KBWKjYZV4OgtPIFWmsY++gYke0lKQVQi8qPE3QsJAwFRCi0zx4eRKUtAHh0Z0KmxgVenA
iMjZmP+SK0xicbmPrcOhujYqXOVGNYZmFvMc2V6J4Yz/I0mNYN4ZzBIO+/sDT4PAGSIFUWLm2rkr
2eKvrdg6S/5xF5CcfTpVPUbV7lqkyJ+RM4nDWEIeItbyqGIpERkbrZju1/CylezfA17yBz2Raq1E
v0+XrxI8feAN68SAFrOr4fFsLu4W+WJ8o2W/MKMYdwT2s5UldO7Rb+QXL/QvGXAmqLSq1/FUhAzX
WFd76XHB+uMqPKc/oghWK2lhCbBxqsM4XBouPXGdrh5zWCbaS8oSLNkpBsShb1nXWRlPiFCFkkdu
gN62ehNFq68JFfB0U7KnFi87fSmS9FjU7c/hCPEf0RC8hGSDdoWdXaSn/fi92sIsG0iq2Yfl93PS
EJW2jnLYBFcgusANwc+fCEUdxmZXogctOo9IuL9HIqHhFDL0Cy2tW/rMEmnIbpVU/lHYwPQ+xLsL
m7DhXqdFA2imqoWsq8EjHERAc+Jiink0Qe3xulSDPH2BBJopPrRq4GtcxJ8JE3bwi7BJ2GgxDXQA
N4DuaeVIO5tqUGARJp0IDgDBtGd/Yg/IkPciP9CGfxhKZo4pDmQRLFFH66hr4Cf89ETxpX+vYo5C
laOKW/o7fgZOoIDZHeMwcKEHDDFM+8gAWvpp4/aycpyPpIn46aqHJ7K2u+n1+Ahy+HmlRYaKzqfe
R3ubWTb1H02UgGoa0t9igMDBgvP6lKhMK/EJP7Z/qEUZpoO6hZ/8Btyta8pvC9nsOfhqt/wwrx5B
eF0qQ8N38AGzHzX9Y0/Y/nQRFJJi0t9LCQyUPafM31bHPUjYeYxubcERLinqkFeB61GQVwmqmcUk
11Nbk3AwCiQQGgM8FUPJpWWip7elv/mCyYH9/wQHibgqg3hQsRvy3GYb0CtdDti1yIv6lqrTM9xT
FR/pWZzBY7zF79Or2QPiApQtrOzjgQvea4D3vMpSSwiMdikWBPMoTjkA/FpL+kab2Davm8v2BhpI
ggmTcovqdObpxYO+g6ovugdxqDjcxyQ+qEC7q+Pj0UvAmp2r+Xqkdn2fHlK/QWRLXsqw6iFNMeYz
uyWTLDnRvqkkiYM5zEhfzjeq35I0ta0FRIV9ZnjNRmIztXyxYh+5f8Ie/ONEtEVwkJLqvccT2Qka
LVxTt3/m6UeSLj1PjsGZwiGUMv+ydIZK6vJIegae3Ets2BNP0srmf8Aw0gaVgJ0es99Tmue+j5g6
GpCg+6yEkumOjYj6gnNVLF0fXLQE5GqtZZVoasUB6Y+VLU4cEqm+lHxwGoK25pV9in6siwIoqwEj
zhIGc4UhymIdgZpHb9jfz2b/qU/5caU+KtEtrw8BPcT3Sk3b88x2OHdd6t6FVmF9bUbXvXcfVCBg
GPeWf6b7V+2+RU8UT5ce9iFXKmh2RYdULqT3TPfZ7kJTHLFD2mghXkb/vucLm53TEE6IdneCuwEc
1j4vkhyl21jt2HyEkVq2G+MbZt5rGti59Mw2YyMpIcknvgoW8D3e0ixOE7UBW+hWPDpggoLxtvDp
TsdOBRA0U8PWhSyopqFzydqaJAfq0sNVDQ7D89BWbWArt8JfTyzLSZ4AlxpvQ9y/9u/NukRvLiTV
zzMxXcxIrRYHUy2PbY4KRyQKatIAz3djhBBpPWYDB4rkqqtMtmYzR1KfW0miV58GrO4c2TTLkqjg
nxwgJ/N1zORs5gNRfQMGCTPxp++RCQdkirQ97rVJpRBE3yWmAgxZck5MgUKpKYVITO7cQ0hZO07E
vZah/OkU4nM45QR5CK/xH6unev2SZWafH92pWSZCxZsMEh+NKEm4ln2h2L2tUghLf8FEcs+6/ME1
pbpsBgUxh8V8/vvrxF7Dn4bjf9cHTYc9Rq419LVvkz/UjVunElmb0NDNJ5anhTTqbLsid71HWIp2
XWMX/g3EyT7GX3Wd2L+6YmBE9ZGWsWrN/xPHJE/XuEDxyrrOUgiCfyc6O7QDk/ZiIB+RW9KSzcBK
5Wr3PkMZZhwgT8rzVH/23bkxtE9JdftdHtlCckZDnWeyBMj0hBOWuUrcB3t4p147Zven2PG/JGE2
0L+fxHuF3Nf6Hopilxq9CHXCq/zEcYJHPPCLh1dxXj2qVv2gAICMjEGqkbycxJNb9kRU1wffJrhU
JrR0OpHSUlR3KooykizB/Z1BTI1TXxkhrg3L5nkvuEsZ3c1JT8zFJe2/jyoZDXE29Rv4foQ3APNf
w5GNKNjwS3+WvSJwhtTbbCO+9jUgCWe4Ee7vkIWlw8Xi+bl5021D3MhBE/Dp1CEHd+y0Idms2okN
EdQEfqyWlwdF/bPj/pdDn5mCehukaFbaYWENlKs/lJ2aIi8HLnDE1xAw2e4MkePCSxgL9wi+6qrF
cjYrIFJe5aHxH37YKJVISqpwBaxvqMHiMgK0isuDWEpsH4XNKJQH6VRvjEzg5PGbKOHbiXLxR0Xk
Ua9B+o+B+ZNaXmk/C/7TIXgwds6JKWm/KmzrMutHkke+j80Tdn01TEKoZGqBJWP32K0z29pkZJGj
ow37JYwxRikfWxTf/WlVJk2wstAsmSbkiRZPy5uxGgRH/OxFcZvRC8aTk7oYOQBycU7cA+tZ0kZa
AQD5a564dG9W8Tq/Okj4lrScWcy30VCz3bYJbSxeqKTc1k+lSjNTB2wkMz+jFmwCgkwTBXi52Qn4
75BmpYSWy2QfWbsKiPtudOksHBNFMxlfCmIqP3URma1YcXlBBRdhBOZC/n4PygMLRU7njQp80NVg
cRE0yXCwgfx6ynliaw7uLtQlluA/opELUPFPPivhXZHUV27tzfAgdvJxjPDqm7KkQvXUF127Ns/U
t1GitYFwSDdJM1izrOUsTUq91kVxu2AfyToc4O4T7s9oTPofnrfRrDeWpWCFt4Hhix6u9VMNF3bN
po4bV3gMIELcMPpa1zdaN5q/Yq6wUOYLAqGP0rsWodc3ruNZFGEEOS1Ls/vMQl+CgfPio5QDsKUD
2fDCSjOtLi84zoKm7suEjs54iGofN94YHDpbxBDPcOmTZ/G88qDjDCu5n+0VsJywNhQd3J4I3EPG
ZUmCRrOdZ4TmesTo1D/SZy8WHnR4ZrMchFQwzcG8ymBwRf81X1p6UFCFfjlh6Y0Ph6goM/3fsPLL
WI4WqDDcYcDWdIFgOixJohJnoJPiQqZtIW8mN/sIUwzA023Eei8tIFMuUsi04TCJ+URnIvAGcNt/
EIUhx6FI0YIgGht5OVwM7Oh2+EZHO8okguHkSuydc4ryfWGrWRVV+5tu0xwnFccNhJprg3ZONZws
cM+37dUXtelRtsr1+VJJgUn2lVfSe7q+gyMm3eWPGXonYCLkmHw7k5BUhJ139++DuBc57fW0fQRz
4b9R6J1jOAOgkAS/wAM8Nqx75xTK4LtALd7liJBhhGkc4qCLDaRyeeaRvRGUUBc8J3Y1Qb1UWRMP
yJuCNf31g4bV31FSTmUPIILlciWIYxvr4zeS/XZhRW+qF80MhMK9LlFb7a1rJXWIj772JGoPm+A2
/WcTjCsH2dEzOSpttpZIFUyO6RxhiaKJ83914hAGhdODSacmjNvbpPPAtRs7AW2Ny/pJVH/ABtz4
ypEc3rLft1eGbsh2H//5p32GV2SBfvEVa70OCh5SyTscHWH6bcMWtPpCLWvwEB4gYuifUPjKDByS
AdxBuDOgv+KKbAcdSlIKKLQZU05BiLB08kAHsSnW9IhGM/m9lRXn/iw9CdMpbmNgDYC/Po4X7J4c
OglgsxMid3A+wnhDzZuztd7U0MnQNumnT5fJPbwHhpv/fg5SfRVadenK70nprhltV9NaJETlAjeJ
dwMJ4w86bDb5ucLgH9pgQgcimIBlIn7B8JsIFmsTzJecQCgtCemArxBHaPIqFWL78eaNguwBfQjX
RNudarX2ncnI9S8Z26xXXjdBkeJXnsGcu9i+WfVPU0RqcfJRSXvjXhC7cEPyJpFG3jBRFPkTUGPF
BGz4Ltxm0Hjcx+oqRf3aqukcohywryUky4UMT3U6P+9/3f/e7GZX97DNGN72r7JpqrWwLk5Mg0ku
Yal6dFnKWINtxuIgUSApsGvsjKOoGlZE62tdcAGCfV3VEdOF6/GXKJanBHMzJz5VlsKkC37x2AA0
FmSQttux8Y7lCr+UiUDYfSX8K9Qp7aJTP03MytLdLhYzQPcH7PyQvE5Ehwss4/MIAw3e5BFKSJvS
iq1vjheqm4jWCiIZoChd8dmz5StdijT5qNFqEQMLydgTsYC51nvzxcIQURFM4Wkxc0e+xZYfs0jt
iQACWPw3FA8O+bR3cvkXpiR3NAEf6AXcnFMMEiiLWL42E38SP08jymxxvd4qL/wOdRvXpU+TSQXn
0TGnKVR0JFOzkS8Xa35O1i0/3QCl4wNk5Q2aI78TA8/u1v351e8+OloKTTw++Dp7ytBJ0odidS5W
evoNJUAK1JPVGEBsuqYOUonua/I9mPTYxbaBUPGi6sKkqqHysvoaAVkS4xAKYPm0cztOPXXFqMXF
13okmnsQyNBYlXxawAQrQB8x9jSsSfbDWeWejRZ6BUl3SJJtXzYxrEqSNMn7/N1liQL1acG4rgJN
J4o0eEVwNl/LVrEMH1BVJ5IsMYoQBHogk2QeUpsbq1EFhNKUSFtKFW5iUdA40KSNA1uyJp06UeDa
rxugwUq74iNQRncYgNraQobpEu24qHy9x8QeadfYMBDqQTJEZWNm9hOBy2FQjr/clfx/Shcq4rgR
KeSqPkROdGGPVPXyNJlWRsRTwLNSAfRjfRLc+gBCza7lT/XRXvubd4Hup+gLNIxegQjAG3/G6B5E
vun4ByteyvHG8o6JJfb/hsRRtepI1Nqb5+9ZfIWCpYMzjnflfmYcwMNO2+Py4rO/8MiNTi3mZsZa
Or2n58Hi2OIzSo+k1IrZHE1NMMB6qCZJR0pFYaxrXhpB5gPXpEdF1ZNtCNBYgfhY0wZzHFJd9aWo
L0VkS+wjdWYS3JGNvPKQf+nPZZUQ0zKXHLdssbEVINJCbIgvcsSXK6H88GET9p8okoOeSHSIeN4d
gq70F9oDyH2XP8vkX++joFCVE3Ct6klGv7otFtcN3XcYVpz42yk79nmdhi+QOgBULk6FKx741wPd
V+rnMRxo4mXif1MhL21vJqeVAadjhx6mXTTr9+Mt4AABkinpUQKpVCDC3YXCzO4HLyYE8oQvlvJQ
Ui+dm5OfXg3knhZBkFKIG0AD5Iv7FUH2cgPrGcy2nSpybZYr0gezjDuOGly1HSdHohHcFty/a/Ie
jydghIqCwbeIZ9T1utydtcSWuafttErqfvy9XfxzpgsM4SeXxdIHuL5NCi6sB5mnS6jmGwRgt8vP
vS/4sdflSwmHVCrIponAkg6M0/CUsJ+fLz3Wz0s6Z6ELYxhjIuB4MIXr1pJSvemnho0/C50S3UGA
pTqATQFnpBy0VwFuBob5LvRnrcJW1o+SnrgotWjM/GT8KjONrMbaSzAdT2VvOpx2NKGtkC5PRDzV
wUmRwEfXxw5eNoVGhVV9XWvg6zpG1Gjf/sYzucE6fRXW4K++aFY1KYgQsrguFa06VPs9IzoClVW+
/sVvkPh5jo8Mtr0wpWSnolMIxUA6+w4DrpDZJnPh6QQdBFWrkfUNlISjKUY1kZ8xlL0aR0Vuu7fE
UIcmzY3b8vqpGUfzB+pcZiuQ+UvJvP1iB8xn8WeobTzE6gH7QOPjDO/SF5zYRBnqzlfw25CEty/P
Ao5VBzwePkTafNxzQhd4lVytAV4niSKqGht85GfGagFaPMhjaYfeWQb2f67v4exWl1Lq3xOahvMP
HNV9WRp0i7igssOt2iohBc7JenPPtTY3707+EgqYuyxUEfRc6fNUWGJ8TIL2TgaVcrqSH46dC7DZ
G3gfKXnWApi2KoI7QvPf7ZqYCtXw4AcBP6Kv+QPhZBcAiVf7NEUUJUI8XSUFea4uJv35EhJezkk+
GcbDLn0wNL7+yxQShE1ZA7FmnpZjHTimHKi6nArnUoQ5z9kynGpKrLhI73P/wKb8PHiQEvQJ7T3x
Y1rVZ8ACH4jf6yJTEpYdrjMfXli/Rh4gQMWio1Os75dw4EWoPGt2kXsWCQqzZM9qeHqA3S7xvxg2
mCFWG4DleBioODzI5/rlupv52rGxp97MB0M7LomKpyvud6GQGtuFHFHtiW1aregcnj5ONE43+yjD
bEChi1sDFO9PgkTHGjG+LNuZ+e2KcoV8rNmzxi0irrNLPQsmOqST44dpX5l+O3obI4k1z6lQE5iW
24JDoBnqrIWtxrh0R1RPCJ1A0AzCmhl1O+ucA6vYMhk/f22FIsi4qAPVMJ2KFtRY2VmmIlJB4E9m
yOgevJe1QZLh37fx0TgnVHuy1UXADsWWARJjWOzy91Wasck9vNQFmH7/yePMJbzamVhAmZPhxqUp
w2HK1TyQp8HBopKgbHoTL//lfkjBcG42PlRocJIXuBfctlkZVwy7N9OjvxkLnvxCKjHJvsR38B2f
IFuRpEntHn2MJZrrwZ+mvFu7Je5gIG8z9qiuSFysR4jhOpD3L4yQNAlxjSjx0YYcIczsarvr6jxV
cTx7lUqFUNRJQIfGMGGVRBRTLbU7Ezeg6dU3/Ufmq3P4DRXLydMY4MYK9ihqKbMdQliuqKfSGYJY
27TNb8DArOtIJ87eZPQyA54G27Eqb4LCVBVVixyJJvN/ysOluvjcgcEafK9iLqssLkMjD13FBZo/
fVfskDp6GuUBhQ+4Gd2vnDDLqGyuojRGnKouCp6jtpJNtGLFK/Oqf2aF2YlI2oH/2GpNFQcRWbqE
T490Y5VsDNIND2AgcIG3d0AscW8FGCCziNVNVCKSRQ1Ed8TC5Y1t6exoGT7CC714/rff8blBKAyV
LtD9QYIinawEWMOd2C3OML1XDha+cA4BvOpIfR2mXrqCekO7az19MI3BgDZ79IE/yDaN5ciT8HmT
VQeLPJaXlcoZ8ABi8b49YLU0KN0C3nK5LMIvOuKdCPZXVwQpTIwOOIjl+1je9BMuI2Z5hgAXvDi7
G4sFM1wA1jBYccvB8PU24N223LppM36odaHE3cLRH0Dx6cDLvq0Jd362OjxufQT2YEO7YZN3nkFi
BoI0LSFtSvzAwn5KAwN3PYmzaVJPI1ZSLlpLZK3tvtThmjSSRTLMMSwP4DHOZ1rOavorHRZkUN46
BmTrL7jCXT+Pb2UTofmo6TZxLh/AKiM8W5wNl7ikoXj3kv1pzbOGldS+LFMg9yaPD5uLFDR306sv
Q6XhtPjrsWSnrqSKwx0AKigL3AGP182IBYPaOHfsqQu0ZRgF0dlbfFWnYGCu40X5bXOsQXN+xP9L
bFMju90vx5U3s2q6DI5ZcB01m0CzIRCqvhdz2por1NoPXc75eNUEWIiYAh4yEuWPT+ttxnK+fibs
Gieopf32k5RScEc3EG6t5fUFaK1CpSbW3nQ1CTN9lxggkQx9ba2/q5hTNui4Ddeb6hVyhQiLZqg9
RdzPSScDV+CrV8jrBjNCc6OUiaFUB3VIi58TqsqXNOG34xlCL0Nq9hlvg3kO6oJxxEMccYTvwtv/
updMhpn6eHtbW0XfscJx5sfwF/9fpVnGYwrZ274hce9C0iTY28g0W5RpNXWcw4zEt8URD0F7BhsJ
sNRqvFSIn3V1ZPY6RgC6uck9CbiMJ6HY361LvxaZ5F/oykq39Faf86Ppm2EBOUtJkXC1OV9pEeyx
6LOnVCBSdwx8XHvIo6gwYjxdJZWH0ZXE3WMW3TOnbGAHuiREe31sM+1nOHPxBIfFz9nR5kg/wrrt
XvXleyzfeUU9U4XSDEq+2ET5eByRN18M6ECSLu8QN4llXg6OBDsw9rAmc8zmSLOnN0odRzmbcQLq
uHYNyFY/LG1g/lABTZYFYUUqLllTDJqvKYvG8sNVwX/ey9HmjprLgSP3kOEZeqrp02M4rw85+xVk
OCuRtosru4QC2sz/pL5noRu6YeTL2SX9aHvWFARBWTrt/GJVQKf+jrYNSR7d3oFEC5OcV8qT1qq/
9jxnbh1rNbgSNBeg0b1MgQaKMl5uSUNxjOOLBAXbH2DMmqxxNkCbSStWdId8Ii48B9917bRx+1SL
5Og99IucetpgBHtudoBBv0oPXysllSSPNr7Di0KZW84N25OPhCI/U6H9ue/XrnnU8qfbLkz3qd8X
SpUzEbsga1n8cmaZp2apkfwAr1nwZVHv4BctCuQRkGJB1kK/oOQjuCJBVQtJSX6gHLEzXUYJPzZ9
lHB9VkOzgyCSN0lCXj1/73Rm7kqvjBx6gtEUDJDzO6Vhi5Q5EqC7dLb8n61IPkl+Z8QEz1Y9LD84
vrqSAnPUcThfhzhm9A9oKH2u8fYEmP3E/We7sIccuvZCk3JfW4FX9IUX8M0wg05hfulSQDbNTu/g
dyFqUFQcVZwJf1mpONCUP/JpGvothzAo2k51MJCDS5Te0ilTKx7HgbZCc8654FVeVTjJD3BTzMru
oRm9dQQBB24VxBx9tgw74qzK5EzD7WiQuAfvOJra+MSeZzNwtaPInUJQ9DRnByuPmtlgbbDFOm/i
d5LrmqYZdz/+NgRiODODmv43tSsqY6UxLvjgQJ4xSIdcSknfcksnx4Ifn4tyOOqZoaUBDeBOI8HY
GPwGUEEZ1atrmwDghKnkmt87r/hsQv+uex4H0++1bRiJrDJPXLI0v03nYTXFEE1J0GrSY9tRzEi7
s5M8cU/Qvkyd8DCSwF5xb3977LFX6ISmzkEwM9QbCFGCO2aPRkuhagYGWOjNN9ac8bGkrRosgQf8
NpsafCNlb84EVzwGYvosWx3k8/Z3dKF9s5IEMGTIxWTbukmmA++QO/yPZbMcO7szWLQL+qkxgE3P
5MhjJ1eyvop1gxI2qUTxY6HZ8zsiwyN8aUfK2ejEIWXrn+Hntd9M2WkXNcWC/9YU4lP3kj8AaDtC
32BTFShJpLxGOoNojEb1EgksSq2zkCxgM1sQnrK6pBiDYmgzrTwVI4ADHlNFZpXH9tqqSEkPQGF+
xPSsagtLqXkqctXtI52V5L9j2/5A81JLnhpECZyb5ajKFf0B/gZhvBkpBsh8YaMa1dqLLYLk23Z4
zl2X2eydkYr/v83h1015uakDvZlF8SjV5HIu4N8kaq+U1KBpbISmsO5hR+RZDzBSU5hnwtx/SuHy
JAErCbbFlRGEe1Jpvb6Mbu1FiAGJr2TYOuHHhgcGTfyhI7Ml7uzPtoMlKxFaKYmrvbaWVls1qqL/
Eq9RNH+EnkZBmvzrvbIQ8t54znhB4kO+bJ5X5U8lfG24KQW6iqCGY21RdozCge8calT+xJ//n2ro
hGgiclzISOUzeztBJMKMcicZpGBZzPaA25JhJeGKA9ehrmuCje23Laq2NDLiSMAlB7J/MJymJuM3
m89fwhv3Xxn9o3hiWy/DVT76QNgFKrDNkAajIjJyeFKH/IH6AhA3V84y6CA4siNyAzKuVckzGcXF
QRk7239qZa4WlTAx5qWcu+iPjbcBpylzw8kbd/2cwqKBvXfckqqRbdtvmVrUTDds8F9T6ONARJOo
GUU59d7VT8zEpNZmLEk/FvRG89WDhs8zBSzZoZbYHutMt+f8JHwTkg568sU/iRP1y7WUccaDr5kr
Fxjr0KMDeEW9jDEFaEE/CusREuC5yAzVuMiYqWva+pScEUgtOji79nCZezbObnzURNwN1WwqK7Sg
CN76hW4SHtVd3nXMa9NiQSex+cYa/Kh4TjYrKw8AFhs0hkNfmbIgUcylWi0MJxib79rwr5PXqB66
lo7fmVEgzwdSNfA/6mxpezIy4tSxd9jsqtIfyx7JoqGGjEPIcUtra2yIhX1iVgUZhjsfZQwwU7e0
SxfpwA1cYo+X3RhjVTmxvMgv5LN/rYKaFZ4OYSGj2q+m4GlrAzLxS9QByoJl+lyw8efexKeT9DkQ
eJKduCI73Rg/+gMbNFLYGwYxBl3Psr8G8OCRXeQaaqkUfTQATqkFopJDzp8PX/n5DRuIzaS7OEwY
qwl8F03qOU3AKHA08+6TlzIEBiDk9Aoj3bfeoQkUjCwp0yTUAt5WIox9CePb2Ik05tgrjfWz15TY
SDEzCmyj4c4ylmr6bAmh5u6peOZra36VxaKqhPGhCqScrL87T6xIf2ofHpdB+nd5Y3n3/LNJj5cd
JkPAqy0dD8RrwFLTI+swb990bo1f/bh/gQE9PwCE3MlS0Utaif44dEAIOfV5HjeFcfGJSsnQQioH
CKTmH9Bz5gb3WzoLa6iXIItqSFB4hLhRCf3zIpY9cbM0Q8s3g2ufWhgPRGVmpgYcMrpNcTfRCgOL
Zw+aSd7uvLdewW07Z+Skl/0VHJbh52j4UXdz621nxFFJ3fEGcl5+tcEN1X90jZ9FlrD2N/xPLeic
PJQ5kyrP1HVB0gPmeQivmbP6/TAvqBhykmiAGXc73zVhm7EO+8D067N95qjjVzOHB0X4eErfE7AZ
d87CXfxtaVUKmpwtAgpHO/3r6/+V61e7CtUnWHG9m4QmMMTE1M8XOMQNoo81kGXiA41fbTMi1cHf
mA8hVzDjIoEg2y1F+bjQ5KrOh10P2677RePK9LUz4HHZVIKhIob66J0/4dh8JlOogmQid7oqNkV0
ey1hcl8ltsutgfjl0CXm/fY8JmVKbD94xWfe4pNnTrSQ2ZzSVl9ZYrVs2gf1/sNWTZe2lxHUzIaN
OEWYxG8nZv+QdpmrfJfIXwr9B4FkpnBLNrSc1HKRpJpT+5clZp4lvwVsoezxjZfGjwj7kZ+WgaHn
9vnzqMc91oOa93Sq652iQ0A3VCEIDV6uSW9Dptsljuq8UQFb/7hj6h2sHjUCMm8wZYWeu7cFVSk9
0TZ0DbAcUij7ee3IdV68Fu3MuRqrK7UoXwFgHPiDupcGzlKfpVk8pHnkDDNWFpfZ+bxDRZ5QWOjv
JFjnp706SfPyYoo6TQdqB+OFnTnNQUYzQ3eSdjqpe5rS4SYhSdAWCMAX7kxumRNY8DOiXtaqHg+h
2vTaKOXEDl2WKsrt55k2NlVhOmucxi0+8Iz4TBIwjmyA5yiI9uFDZFR7wYVw6LaNcPK16PSPXC3r
iQyDPUkuukXv4D905/xLNeW88lomz29tBO7AvMYDyEbvxyJra+o/9QzYw8rOL5qPUHN1S/vFoL85
z3bUQIQD1q1CsSi6PQLR1WDyuP5qGEiX87H+1EaV9/SzDvJZwi21Qullk6+rlGG+qnf3kbA26zcD
JRFqiPJOjK8ecgqh1K5WSZ42y4w7WHq6kCTH+gA/dos92hoqbt+UoUSJIn0DeYBSbDCgDuUFHqSr
dxF92fyeDNKEBEDb3DO9lU4FHKVN//S3BSRJbejeXeMLTsRpJLWqz1f9FfAaQhY4tUj2hOZB3nzo
5d2qz24k1LHDUN/T8mseB5aDiO6xa5JTGx6BeqH0K1bPDmAi+wZLP4DkRVYnADqOF44bMn04lffq
z8ZmanYfxJF+sR2CW2QrMN3h9/gGeNPgq6MvmvUbgtjpImWw6U0gkf15MhW2LyP8Dn96eNK/aEFH
6NCSfvvHIf5Q1bzdJqgywxyN7+FIZO65roBERWAOx304HeWyEVacHzDTGrQ0YL9rEDIHo6JP7/24
drcSmm0oKnFnldVSYFEed/w0BfG2bEv6Zh3GLJVaIciMyouwdnwmRCFOyBzcfp3tVnNahlCw6NqT
yqDQzILMLg9ehVWH4zgUCnUP0ouMn0Ufl7+Mp+uWZ/KgkfJ7UpNB5NhrTsKiL2+yGC/X0W89+O30
nyqfJtpD56+IHAv+WhzQzhf8LTkcf9pv1DwPRKdG1L7DEe13eutp53BPhXF8MWSfndkhg7DvBWRg
yWQIBBMAtP5yxgnNmYtWkavyG4TrdX0NjSQ2uSK5AAKHtE+JsMf+RckJkxJb+lyJbs5UK2z3IcKc
wCquXrJW9GcxXetw7kT3nq49ORuf5IMTjQdNf3Bzfo58lWEyR4OGV/YNLvzDcABcqGrGxO4ncYJT
JswJyPGl073emaLGeyRnSdt95iyxUbo7QLg/LvYObVQyXWsPlZvnlqTGfwKamAhTm6RphBDiYMhv
B9rq2pNJd9mYet4pSmpRZRaYynrEoLCyT4JgmFPdKe4BBr7Yo006cn0dUrrwg4xm4aE/ZV0woc1A
/8JJe9tYK0M+v9z3Rq4QgHayTBggtTprvPO/QfSTZwFDDZHfk1W+JnjyT+WmLVp3YXhutK+sAGZq
qx1JkSuCQxeLdKgSoJNbfc9kx4Uf2I8YtmK/TWNUq+nVAWeJqOkH5XjMksxuaJDMc7cWKnNlug8e
6efUqdVheFA20UWr9WQNnWeVdfMm3b3mhO5l8tzCKpdsYaO0KjEci/C5G5gE8myZajJ0eES03Nd1
z6KxQ99dop5OYbD72oVR9WnsdORQpXBSgup9UVbcwF6/ARIqIodGJF70AdYZ9JO/u0rinK7IN+Ll
3gDxigCb9508rwppEqIyW6sGPFOL2bTui6BBj0k6EZUUsHDex2gM/b4mpuoKoAViT64k/Ut/KVzU
n38nY3eaOqRmbcQLGvnsWQfsOgdaGr3JsV1wuGA0BHzyaoUUtYuKPHd3c4lG3Mtlaf5WbkqqXlX1
K3o7c2elTLgTsKa3XbIpi7GRHFMVpWkow91IHtPKAaTeHWS2n5csfuD9fYF6HgC/vf/3RXbZYnXs
B8KQIRYtQQxXdr52vpwHumTB5xsHHfayT6DWrd+L9iJc5bPzb1W5VcKisck4grZLxCYv2iOX0aht
wlwPUL7sOzt7IXDPKRoz2S/yVawQqX9uBOGZ1sTMJDuc7xBCahIcVfkkvGVQ037d25EwyF2sIN8a
7zU1Pg65be8oFl9qbFV2t9537iK+uC0ymKrDYM640pbZOkghCShpEB0IZl7X1BmI4g+kU4El03Uc
g3pLmDP7GXrdsis73yR7TWrl7DfeLWXb+47tZHeuIgNIjxZT8vJaEyn2UKjDDEw/XFICCCRcdjFl
w7M91mecVTjyuL/aMevszqF8HgoWqTtgOppV+E+xITXBRs7BNu7rFKMTJSJLGbKOqy839q39RDg5
rbLfNdb9wcGI2WwHTLG0I5w/DqFS4FQdHfClR9lIoakNS/VLeG3EV8eTc0cMthzGLbETRb3eow3P
6xgMqA4okYHIe4j2adwz2q9FMQL0GPqvtUPgCtedZAVrA7SGXRZGQQqH1H6Frp9Zb7kHsh8NZcHD
/L41+fL6bLzpOUqgFgpTSQX4mesimNRWZXV364Z10kCXV2WUY1sfuTV2duMSlzqhgf/bhwOmgl/7
l6Rf1xaa11xv3QczeQvKvX+fhy9u6dcx8oIdL+s228tt6050S1woBQHaLBUF+mDdbiX2jB1Jkf2g
O/1B9lfk5iUNqZ13NgGOmZsZbuTLp0GlAjJYSXGEieEKWTpVFaDtzM/Lwgdp3B712ZM2WjyWDOwu
hnopa/kFjfrZBXTWR/RqzaFh4bmmcK6IducwxK0ruquwt8o3Lh7SIfhh6YsY+DGiAK3I4rL6tO8S
Q2IZ05m2QFXcXZsPGWq2ZnxnD1ESRyRA22RK7JnLHvO6qJ1gyZoL4DTqX3zFFidIkP/XFwA/lk+r
m8HhVmOVXhMBVzRpqVDhqc8qWx60iwrjx4328YbPfYibIb4jQIm7bORwqinYDk2e+05bsFg1OmfH
2FBcCp+QY+36IpWR3oGdZHcCMhAzHvOKbzSvf8652nY2ufL3NkYvDCRZFw4Eak3XlbSFUAnzgYis
4ASngM8/nIT25kWyZsR/UYPy4EATr2BC+gvfnSIEXCNp1dCVpWQUi9WnI76ZMtEf/SswBdzdt9tU
iuNjQ80fFRFy46PoMftKepIqBlchNqm3njOA4qGz+9QhGzAkVBBH+WLdbaF9wbwyzY6XmaRDTPiu
KdxYc6Y7oGanGmwXUhLhp+zW1nhOKCaewak17YA0kWZk1mFc+wIjnPIsMQtjJFoLKLbtU3GjeDTo
75I6CklKwsq4+e1okJYCjjj3Kspw33xRu1qfD9qhzjuewnRBXFkLmzLahwIy74N1aUSWUehTPpq3
Hfau20q9AWNoQ8vkGu9eImAXyo5pZQE0xzrCev5FNOXK1Y/Z2BunnD3rVIyOHR8MQRUWoJXjiMKy
Vubd3LCFmt6QfNxSR19P8kV0opJDefhwKefu2qyQREzKlu/6xUvE49aGtl6gvUgpzXx6gC/QXR4d
BjIFSt0xHv2d8Z1C0VdqmP3wiMWuSfBVxP5Jc1ygH0kow7rYjVk4yyVUTCvbfxQOVffrWaty4lMB
CkeG7bjmZkx3rtssy6B/leXq3g18zTHQGhJMFTX2U7JlLnSBiJYAkS4v57hcAvHE8+nwmprceJCu
bg+je7JbMm7LQEnzNT1lD9DB1ocT8TlsadBLeV4noRKZIQi7t8Z1ZR6DG8JdFiBKyDQqFo4UpVfO
lwrOxR1YHxs7zoKLDDC8s7M7avL0q8pqq+lIlUsyn+YU835QF4O9YhgmS/m4N0eSZYbMug3Ykb/M
nbGzAPJDtHvN354kGnmI+3BQ98P8NJ75INIWYCch3TU7crFjlrCx/MNJFAEceV/tozrY7TydAu5N
ZwBIfwgFzkjZqusKaBNeEs7WXvTBIcj8gVg/EO/U5clL/zNvVSpmQ7mr3Q7z7gRrLR4+kkyXyLiZ
pq7kmP8yarO9DVM9ZAjQ9AyQeeaL2wgDzCP0zIYCDF++gaE3pFqyyMqsOlDDaaG0aDCUK411yfZn
e1YTxIhaViAZoNqLzQ4suEDI8iOaafrWWi8YW5Aj6njjNwaaLvQt/G6dyW3Z4Z0MISLnoFhCRTcX
ll5qipgr2Wa3E1QjU8zF+EzJIT0p+Z21Jb034gHc3q4+jAJveqqEMr3p0WwU8uTtPCpJ9KgFG9gG
g/xRtJgPQ8wLfhkPxnFe3vmAA7osVwUmmiT4cXl1A63gBNDSjt9aXjRO6WtW+msv7k88OxQyIDz3
Oe8oXBVLF+Taebqpj5/hHa3qaTNQvEccIrkvWH126xICPVD30e8/KcCMKe9ApdVln3eGM4ppvW9Z
arXuN5RF4SI+UXKxClysLa6EOMZp5kSEkZ27B+D7u9RbQ5N3owdjwKtnM3wt+/RARXIh0hJHXA5q
t47e0k5x95S5ijIbfPgS9swAFVQe8XTXhxixafsmVGMTEshreiidyDevtBp68yC7u9maudg4sJRo
tN6b66OZ5srTLLsBrHrHmlWjyfn23RXA97ezDT/rVtdosiLdPgi5TA/96CLcRZSnBvzKzFdpj4JX
xqvHqN6TMZ32CpRDAZJjyR4vXvsNsg37Jb/6YJ+3Oe7fKVsjRR22fFk5JjlVWpA1nYecxYrmQlT4
ziiIv7dB/EuKwMkhqiU/6wi1IQDGYMG91YT3i7NMSXrMi0th4khin9/b8xCCbFn7iwQc6UxpP/JU
4bBw5ghxFKjEKFa3VuHuc6my94lvow5Y1S+OKLY7wPngMLcsdPPSgTGXSpFsCOp7eXAIECDzlPnl
9i5W2661ODTLH+nyxjAyFROdDxd+qVbZMkAO6KnJonMrXp05ck/KmzJ1u1ATFTcn5IejXzETyiea
GCWOsP1e4iy4JoofYGxxdqZj5d4wkHceFR0DI5IwDdGIzjWyQgOAk8P4a+gEVOqXFAcRwB3nH672
Bl6i3wVBJwNVs6pDl4AciedZVVET2mLV6rGG+ppYBlqizMa4/T9p1TTeg5soOmPPdHm03na2te26
EaakeO0ZkBD25rmTjLdhfJ/fSxQ/4GJzWHxl5tk18N9V0b6RcklKVJdWJAh9tg/N5bZgrnKgoBwD
svGxc+HN1Y4T4OgcljuRGICRO53HW79STPaqo5hTDsrHIgAvN51U4rcsnSVd5pNC8Cp9pWbvIRQn
hHajLQR8FNJanbG2gnjCQVUauAenM0PN5XYaqc/285zDNmTI2BS3weJznTHV9dpS/KNrQWU5A4rz
phdkaZK0Rg3Bwm1XelMWfxYnwn41jkuRKnjxgJ3nhcnhs0n3OUIIQFiEVlkvBc7ury9Y3URXYRb2
w950MxkRZYjfSbTtwNfAjzoaMYTsVoCc8WcuBBOVi3yg5ISqs9NGZmXXAIGwk8oafcJDC7MarKXo
ETL7W09/drX2UQJj3h5yMQZIgBT8JjQA2ShibpYmSLdcO431aaMPXvRlhh+4c7HKQ1tvc43hgAqJ
K0RSJ6k1xrtaeBUrSf6w+MNTabsqx5XgKRazVIOorlLYsVcAbUmHeSGIn5nefory2hmvytqfro+R
mBIuHhPNHEaNu07wVBEKiykeOC/YJxZPgk0t2FoOEGMzj+Hik+U0RXi4Q4jvpKaDr46BbwPeyGen
8YPrEgxd6U4iIjYBmbDfDO1x+4/P/1Of3It6aFi360mG54ef7uD1FnPpTrhDlO1NTjFVbZq03NLD
mxjvz/ZOYva6ZsJM39BKpjMCScR0YNAiDxEopYiEQuxhujRv+y8NSVgvyfOlbjr0NYfGEWmGqizQ
2HVxe4Vjdro7MvtlXh9/xbrYZn//JcaogGWa8WSbyqxjXdb17OzDfuqQiHyL14fPFHffklX7J3h3
EH6G+CO9snmbXMjj6DUUy7wurZbv/lBa2ExIeElohhAJ1cBZpVqC3cuJwsF1Pq0klfp6k0K+JUw/
WwwMfItavaMMi10tNprl7ututDbH80QZRBhnyyvEM8Bvk699hvYeD8qcldy3XB+LsqjoWAOLSvTZ
umT9ASwFvFH0UG1BsoI9mJ1gHQ7r/bNX3XFhrs7WEuWOYjKlnLUmyHRojwEmAGc26xLDPiWOiBp3
B0yHDpdDsHJlrfehmCCflVnG3xe7A8jaY+mqsQ/bxxwO3f0fmT+HlaHf9Hh0v5Veagac8fTYNmvz
dOcrjJQsh44qxBKNCCvWe9VnQ/a5JeezYrM/GJBTuDMAygimstnOQOfMAUwgOAhHwd1stAJi2kdO
rJD368zZJ9CMKyWZ9JGI5+ufRc6hcQb4ezWumvTrdoob9myIux3tkTnIu4xIOUXHpWPbRHoKNqwm
F+wiul4bTzUaPkHquv8ZSkJJqODYsmjnLL48+N1TLXMp1GRPo6SPVsgr64X2f8rjJubXorW8h00K
SmrPjlEidx2WgBG7edNzqhyTAA9mScLJjlWGvhwWnqQt0p01MTWGN78khjDeLeTKCIHBG0vDDu1e
lfXLqlWKDjtQBXK2Ipl2kNWHX3gUd5gqsGZpR6C3bn50AY8K2uZvjjiMTQcq67ZLY64peEyICzAb
sznyHRgi4Fu86iSHKQ4TvGeyXx6rYG6j20dNohndxpEi8OXh2BWdFkjGDFIzW+N+FKmQf61KxXBV
PJugA1EL1I0g8EFNn9AF/PTz85WzXfpYzEGfDo48XJUTtZdi9m8q6wFQ/b0o8VWt/uHiVMEwlo3c
TYEeDo77Bg3cdqCEFtIa3LwXgXJFkDTlSWA2d9D3oxEJ8F5M5zZA8OJK3ywkphw4Qqwztc/Qxh+x
9a+Z3ackC/C7M+4UdFRJl9co7EBxrXdFY0i9mdnRSr+wsNKMi8Ao2XuPfZ8o2qJ4Jit/N9Ul4MfM
9S0DYoQL0ISo493qbdVwKVpBdY0jyjWZRwKEtWYb/1yzpfSn5pY0WnveT+Q0ZfSy+USjfgq/bOWp
dd2utUphgQxUDR1Fi5d0r1DJRfreKcbkIIKX4vLTPBZQaq36OxW5F1CxETgc+YaWiCSE5aMlq36h
CfrvEAZdif9fBB3rkm85cz7tCBVf3hrR4Ar3N++La0KQgfanmRytyw3LS264IBwJwB/a7QSFCE6q
iDob8V0W930gqfC0qY17z9uHBFq0yQO0MH4EOdZmSKyWfG8dTIA4WgzUttSY4SHf4TKN2poGsiBt
GE8+5geD4Hr9X56287hAvafmvYSP5UB3xebfWyJtQMr3EJGZFF/my8PGpi2RxqM0Iq6s+Twjh2Ur
RhJ+r5EPMkmStW+ipTvimYTelwpHAKgah61JJuLjPXLmIFhNGXgXJttf1QvGa2WiIh0KfcT3Plus
6qJNf/fQ2nlU0skFv/72I0lUwcim1V7prHpQhSNvCQJXNjUj3L7nCh3ze1vDJsW3/jrjHNOElvbF
a7ddqMW7/S3Wf83zguqyCFgFTwodpgJTZdFYniV7yXYoIvx0oIYjzFOljzkbyTl5ZaJssynGSnur
1l5Ip5M9jJkK2yrSEyBgAs69gx0GnR6on6CwkX5TToVm62aVhk6sDqAAdFKwfLVUieWvZB5yfbNA
iKFnMOOC50OKU1YRUZsgULgK+Acv+/5QWGhGr3XTxEih3/RZF415csYke2Cl+ifA0n4YZqtjQ34c
BKmexjSDHsPCapYJW1yqFXcLbpgtqkTEjwfbFKmL48pHWX2/HV44Z6fNmCmgsF5pF4eBVsS6hjuU
xY8XMdYfrLvXnx+/QSQq4dpjrcxB80hm0PHuGxOv4+2Zr2CBzqCJHjnlpN2j2STzD3k5KI+AXFHV
jQgqcHG78EvGCqJ9q+t+WfRZ332C+kqVDcISQHZ1Kp5y0lThNf/G+2YkzYWP1r2ZAcSaot2u9+an
wIm76vXeU0am1f2T3ABH0IF3oHBPCq9+22RXord1I+E16E86RtCIOSAGyttW3LD7uoOFYrPywfCH
bAeRd9Q30RIo0rm2xK2HGb7yeuLubpX2/llHSfwnoB2+A/kC0x9XE+v1DsuLnBQbIIyQrmvpWDY0
KStIkHoQWG2MrIgpBt3lWRslWxbT/j25V4bbX8bZwsp8W6MNXyrLNM3QduELcXaV2q+maoOj2mHW
hEBKlE7g/XogUeZHVpAzInl9wztiTqheZ96MlRy0ONNxDv589CZirSxJPCh5QWfmbnVcSnK89ZK0
VoGv+SrpYuo1YdFXMq3XFZZ8Kec6Vbuak8SAIpBwNGdeO6J/f5GZd7Ls+GdvTPcw9cuyY02JK64w
VWb8zHDyOT+QIUl0nUkNWJSFyRd1eBfCgfY66q9T1UnZ4d9jFE+aUS4xeFIWNDBExE3qA6j5XFS1
l0sNE9sl3w6o5s08bixDf+0AYizWNsfJux/KdAo+e5PXMo9/h657pmY2vnZph3gd1HJmKkyhWT/Q
FHnNpMwMs4vSxsQox7TYJVBSoIKTq4lzrsydAbIb3FxVYjJ/szGuvG0JtKrvfHmoxIELrfX0DeDD
x2ejhmarn5qs8OhMauaB0LSM2tP2EP07RHLgcQIMbTZwGOoAMT1b+4y+4xKL2Wujqo0KX7goB9sI
7B21Wi7dYB+ecFF0rOl8CN7s5jedmYF7Xzstt2tg1mb7fFz/F6RFnC/FBZ5JKcPw8fvGX3eNJ5th
PzrKFRI0qgqutNOmt1DeMqNKsnNepq/Pr64Ce77HWfCakRxFT1Pnl2+rVkIS6uOPwE3sDh1iPwkp
5arCF08dhq0v4mAS3t4vA6+RALEYqADDDZUlv1q+OrVrmDZIPRsn9zUxL/Kd1mydcfPc8fa1GDCN
CCxnmdoqfy0rDifBuPz8krAUgjfddRODJ8wJMP5kBTiaJkHlcTu8qVJLi88lY2TLqK7+JRX2nASZ
jGFdovwSRe8B8VCn7HpjKNy54B44RwAGPLdIss9GZqmtM5f4GBiN1lChcibuKvbY+kY2K6Rhtg1i
oqNi2z+Vrs2v0Y345H7PvtI8/NozmjnrrGNw5DYOw0gL6EAc77jDVG4ue+l+Y4xzF/QfVcZnLqB6
/ZfJjoE4al2U+K7rngHNmNIJ4d6bKNzwCTWfWoo1RRwY5YbOesERsKvIzcRlCqmpbzKno6QoVLuZ
qbHsrY0p6HvtvAGehhl3gIAHf6o3hQVzfNI3XFUKlZNE7EcqNoywlIDSTk5rKu1mkTeaLbwajiWe
aazoK8/31pXFDDO61r8vrGN5pMnVU1yRR7Qq0j/uY39WKvbkUo6vtVCjgEKK4O3QPGAho7VPsKyx
6x0+engDMmVsvdd9UBLweuTkdImhjoOtWD3DRnhwqNlCUKUSLcrDmqglk5p3a3Fjx1A7peTSQjap
2gfNpPvyrYCKsBB2TPibG1UtkZ6NQdZFVHx6g+hqNMyUaK8+p/2UxICBD5h0n4mpNex+b+QpknqO
mAgVlrZ8cBo9+IowBk6SJnGrKpHqc67H9hHsfjjl5rb3GZtgX1t8718VJLrppGRrVA5cBYWJcrx0
BTpvGjMxQ6TLJ6PXKfmS0SJDMVdSVNT6AfuuLgCWr93WUuZzGeSmsi2M9YHxarMNA69WVGBmPrdZ
6EorifbCJLQuevDDnHXpoKLuAcUokUR6wkipRSTHeH1/nVxdc6NmgVF7ap6E7K+VqtAnGFHzut/1
COHTYL8SUKoHva3lde4M31WKVjcmG5TKPnz2ppTMof01fO7YqADdCZm6h+FQkqgQvbpZWWfox/76
kUdjCP3mFKzFnVbYE6FnIpLA7oZpx9wyVZ7Xk3zOdRlyfOjYXRzrT4d6yujqfWDr3Ds6FYReyFS4
rTA8+MkCGE7YHEDvhuZQVoV5AjRwAVvVTTFIpu5/PoJK30yc3FirZDny3QlM04SbUS1u4jh2IHk4
TZU7hRtu5PPNHt44lttB9HnUEqkE3mld4t/jYfQTSF9ZD2NpK44uY737eniaHcYNCS9cuJBn1mKQ
vqRRTKxiWmyWucKMm/PPA4T6WN8ncpnvM4IDyzAp1t8EPxf+rAZs1nb313xj2YMwIlDp8rAel5Yo
Lso00FuDwHQixhJn4r0UwS+XNVeppIV954LXFm7VS/j3fRKc+oQIdbevxrGEJDewiqWIUVwajUSz
M4TiUk4nlD8w61wTuRRmmtn7OSS7za1fMjof252l4gJs+3IuLFG5aZ26bWJX4EUb8Gsz27C8XyX2
jh+XMrnMWBFTGnSnAO2IEQAfbtvq9A8YVO81aOUuF+UC11v284lIxFYZ89oWwNrXhY29gISZ+nby
2qk78xN1HIL18gH1UKQ/PsoATxFIebg6AgrVbEk7JNC4Kw2v4/MWqX/uOGYijS1r1pn7nd5RwYBd
KIq4HWF+pEIHugThX9PW57dems420zj74MzgxZe3b5vhGAIfwKvLqySK1A6qpY3pdoOmDX0yvMOo
TOggIGs8rllN7ambtgOi4WdJo8CJ2JW1qYBydlgKVYmDfPxQwBanQ8h4U1SxQrkq3+15WB1pb48k
7ASJyE+PjbCUjeCKx3w85wE+YP7WOYyATLAm88Rn4p6UPuICHjCvo3JNZrOG+IpdkOlod3Hg2Lzz
8PQh9BMY3nqJ48McXTp3GJShmBa+Ioh0y3MVfMCKIUMxzf4QsWbMQoVOPcwz/LIe4mfvWtP9zZhj
NLRm8pPt/29xXunye9e4G+e6C1CWtdJecWlaIA4zLKlN19/1cEcaKIzJbXzTum8KhekXqRQ+9Dxy
LyoHddoHA9Q/gKMgwnS+o0rk5z04HPuGAOukfwYo+MmQkduHKYYWeiHgcZSVV7+0AHVGPlaG+2az
1eo9JO5Y1yFTTw3m1xudGcPHOlMlv2zJfDeJqWZNjZEJeOeGYhMW8p0Ou1Ni+O+6Xv+JWJ9iEZhJ
Nyo/kTrZy//Epyy7cs5AEDnId2kpMEIua27h1XI9NOt+Yt9qRDV94OApdLNF6mA8YGGcxh63IZUb
7NjJwQMkgXvHq1Jq8IHeVFP3/zsWqMNwwRW1Bsmws/K4rMB6Q4Qj4FMNIG6t15rC4WLMeTmXOWb/
tH4+30BtZCndaqUKPdqpHcTbZ1CIM/1ia77B5HrYJQxZ9yKeHcEI2ZlvAY7yEB8PZzadRkJaIDwQ
33ukgT9RAHFhlo7ckKazHL7byJkaorh5D31drx7louYrrYvFeZS7ZJthQnrBWncI2TGvYurTcTNJ
gYGhHX9A2GthGzR+LOgPlH1qf6o1/Pd8lT0OBu8ALEOQE1u1P9sdrcAiwJy9uWoxJukrwRldmytB
OPDZbX1Hw2e9XVD2tyP3vHyUX7eAzwKfecmc+XY5F9CYVxEXxO6U0QfhCoAunFOxjqppRa+qXb6+
tfTROwHncrPhFY06EQKqUQJF8/I0Lv4Vt0l3zwY50V1LxaxUZywl4T6mnJ8ZBmaTJIlSeRuTuYm9
pj7/I92dbmLxqw3Cfv+tiuGF9EVuG6YdHzedJU7KBITPEXm29Av0odvOdTV2ydfUQXzB4AYygLmM
3XCZ0Qy0EF0h1MXXO/8Oo380gCz30EjrBZ+Ei0uh7Dx0j3KYZHKLwyHGvURoZlgBBkrizj2jjgmQ
p03EWgc5uMS63w6ZzjLXfUgzwsm8Ob9P4aSpToK80JboEJqB/TDfb8z6WwHPASFJ6VOoJ94sHxd6
X/NGOQfSY80G3A2MrcxXj1AP0RS19RNFqsoyh6BuduObuMzmzLs47z89XL2V5rHIP27PJE/f485k
gjfi+XHxibulBCiuHTLFI5JW9UBlqWFwiOOyq7WkpbL4CnamEHr3RTlZoZhaY0inVl+sY4LygQQ7
BkYcfOgiQE9MGCRv3M7DtNQjcO7aZMBw+apMxHCW9W0Vl6pWMO19HLM2F1hnsiDDOjSNO2uPU4f9
kcADJUEVBawqEhYAODwdkOzaVeR6Z71tH3WdVRByGs9gGvhWsxfGyfK9yi+kkTMKZU1n54ZqGD9v
ETF3txqO2bUSGoQNNnD4xON9wHkkGg2OryKBC/X4KjkWZ13ul9QeFZSVmXYZKiyUEfoIDUzifd56
lE84GxWCbITSNbUFZTEMVY56ZWYnJ6SZwkClWFg28d2yl0dBI/IK+p111Qxdo9GHluv6HLSYS4DW
PpkvoPANBZ8maC6CIb6AlSp6j5XClSwwz1lWupWKrAA1AJZmmEvW7NKewqga79rZyCgYvyqr+/bf
morol6ZYX+h/G2rthZjrlpI1DUS+IsKhd9sOvVjmD3GIWLWGURlA0DzbX5zZQes4EzV0c9zth2cJ
ViwglT1if0ohXeT99GjftMeB7VDj2asZqnRkTT4QtmZFFgxEVy3/nKA8MzYVKLYjJFq+KlWIJsqR
N8ggIURpIAq9MsfvimVF6kK3BwDDVxWGM4Ej4nHlCT4ArgKGpEON3YNhrwazF6Ym0nJqwvoK2SB+
wqqmVuiDMzLs3+MmkGh3epUV//lrbH6r6rtoYNEZIm2k1bbTMJtl0ohvfDVm3B4Xb5AGXAzfwULb
PybDLOTb21vXOlSdKJ/1DXEBS9QZSMs7T+JihDcJ/2to8g2PGIOz7HEWFFay8av9hrD/7uii23A2
nZJ/AeCEnTrL1l76HSMN7C0P24HSc0FtOMAFNSKmDkegKvoIZejHZnN6+G45gFJscnIR4BHs+Rhi
9Kk4iVEVaWCi0Slajh8kRiigiSLffCyqmZvoEkQWdL7gb58i+PCF4wW6xcYTRKDWrpUW2Dydl0CG
F/Yv3qXyD3bzmRglIIt+T9YZZ5hwqp6efTVGetyo/srHU8T7A6KJ57O5duzDw0lzUTptS4QqcKTb
SvBbGFmJxd0ortmmw4b2mpdMXwqZ6EmtusBjnvdJKvmpBY+b+3Qj8CyLai5I6lplg2Hfp6EfO3SJ
7PhZkd9sC4cwA67tRLVz2YJTejxpbf/taJ+kJfyV2DMuWA6Jo2PsuXRtVbqV10pGOhkZ26z1xyEg
DT7Ork0eUiG0u1MfIi2BMONQI6Iwol7/LvV6iSEFyrj6EKrNopdKD5NzxolN3bbEyd3zPo66Zk02
KYSw2R076U05uY0oyQIYYRmnZ1UTXum/sKpFh7gJOXpRIasXYsfG/vK2NzzH8TcorLXTPRGOWkJR
zaJoZbgwdIXaBR5ywORF044EyEP930uvEL/1UNPiPerJQvgxzjC4SJga21A2T4ukf98U5HDa4RWX
3Jawa6kxkxDsjo4SkwfEx/Ey0d4T/a8juf+/73XjD5nWQ8O2UEhN75yuJDQXnVt3CZMLnynKV0M1
yz1YTSjEr/PI0OgO+Kk+2C2oqDDeAu2y1VuQaxP81uCGOGDlKUTQnEnwjPBb1bOcpN+oS61MxiRi
YDLPyy+roTXRmxNTrcqT6jV2LSfxIIFOIbIvp5GXQXgSIyVb68zm9+3TR7nn9Unjpluzpg3fr1lV
dYzRDRFVOTpeyb02aOmWfNr536isBl2Nl/pV5pb7S0mOWA7uoN73KEkn7wR76bT1b5lyjU0FnFj1
pCIeSsi5f++q2Gk1wIMOmDiRfHXSmVd99YrmnHd0jjsty8YGENclmt65jIyV4kTZnkavXpkwclu3
FV2q6JDx5/S/UaaZVSOeZi0YoQB7+0oGUe8z1m5gSy2ClEajOYfWyIYvCYwZqG4Dzyb9/6KrGoOT
vVl09kwAEVih6NRAATaDvjKeJKTVmmd4h5aVoUmZBZBThYvwL35f6R9WkZ7tep7t0ekJw+KkwP0y
J4eLdK2JDkjygtSQ2ak2cqwPoWGRuuQd4VbiEa81ieB+rYen0aa4AcpUJm/JNOXILEZePZWNgono
MZpc2+kM9BcEAMc0pTL4F3WOJzexvullCVQ+clhz96weRe5jt1crhGOKsSbvx1m643iBQEkEKFYd
zOkX96jmCYdOdDeiInsGN9PVwASIZRQv31lCoIroXZ6dPpbYBxk8JZLGrh+o24nnKeGAOq5qQ/qV
i1tOFqCzKNzPv4Hk9SP3lkYGzqHLh/6gJb+I9IqP2QW/5ddKDrOOTXdgybsBq69MOzUDYIVMimx+
YxVCIet2KxI6g1Txa8GG1DnyOkhgVT7rX5VPUItBUJ987xS+wp13Kh4nrYE9ZPb4av9uXOarlVTt
ZgkRJiOyYpjTxerXIc6kNLDRBAVR4FEjhSmEP2jBL8vyept6ikVdUWKk99ir0RL9lBqlZp0BvutA
fPoNlH/j/8FDUNQUHGFMrDVsNHX6JPC7TBD7W+1CFjHxpPBNmOd9bqwN7Krk72O+0VRbWVq/Ew1H
tRrA39NKJTrKVDgy4QXjHUYwBLPpHXRrLd4GFeUyXq/NAovOzjfi0zXi9YxdEOKdwbTAzjkfwwgF
FeYPeBKI92/9UUJAh7In7nXaYaN8hsLszT0/LZCNkixWnQNsUtmknYlKQLas8ql/zr7PqVMTXDPM
0ALIps8iaPah3lt+I0j+zu6aQi/YlwxVtFaEwMRJXrphlJWbWlZ/EbCvnmxDvHANPuemZCHKpSgV
g25LKTggbQ63mHuslYSAAWbvowYHY3EM+Aa2qwTPt48x83MjisSyKFqgJupi8ObQQoUXbQ9td5pA
3iyzDjc5BJLetf8tRlzep6mgDJVNbwLcl+EU49SeE56MC1/c33MhUuEu4tSz2Epk+rapPiYJurHJ
sTxKJoAt4yroarSYRhHd3VxRAZiaJfty4H0EPXuZeU1R6gLlzOXDLddfvrjbjyU9L/D8bN7HfOC1
KPIMyXRG6BHdbIN7ldA0B4hbRVqrIPlThIROW0MY3rameH1yXVEO7ZR7ldO9myfoe6cu2yf8g6Uf
81sXeOqAbddcth7nKvP9RamQiKTONUSYxKoTT5yEMinJbVsU25HxlI3yh7wQLpFOTySSMJcO1LFR
icm//Ykk7lrwfTKmdSa1IQYRGLfaBCrQcMZ3C4HmRqDkbJOkKKPm8I9Ih30hH9kb/pamwBr7/ujq
2L1IrotSVpEP0XgTgLTl1yUENTOGmRLsYT6PH3hLuDRGHFjUvol8ffyOYYoK6ap9PLPRaY/TgHHw
N3E/0jmErZf1jay2B2cwY7461ZXIqdznhts4vGhyZ1iJaILL5i127ReUEmBZPJWiYTuLYPO9eB1Q
0Gec/xWRZ7zzChHC/BuGw4zDf6sC7X6f1SVTSJ3Ji1bkTlGBlwkeEkiUP2dHgx8/aM4MmnEGlIFU
CA0img/FZSAB5yaDkxqfcoZlzLcoB5kqjMPQ+1vpFgCzcib2QeHu/xefGbbh1sWP5pChHXeLGKF0
gC5x+5rpyJUi53dBVz8WN96OJqE1OLersNQT+AU6F/7fBX/Lq6WRB3cJ9zLWJhXLq8CEVTHQxuzs
0nIlz/Rw76CLuDVvFzojoOQiImDngSmBjMywq9L9cT2/GPMEw7okWke6t0BeOeUTeIZq9efA5+A/
Wc6kLYBQFD2JqyNVA60IIVCnFZkxV2f/uAuRcflziUD2L+jvUF2dhogbkAh6IPu2kTF566PMIHi5
JIWaC/fqOmFK0sxiwINV96aoP2lJPpy4RQ9Pj+sIilzJaDaW8G4870OTVjmPxQVPyQLJwB3hmKB4
bMmSaYTkDpypKNrLE9NKU6rV1GcAjbDLgXHO3j/pzrOdPKQR6zK5qYVU5t6sW/PceX+UXBGUEcXO
0SKc6e2Vt+/pWbk8gQOi6VP2pd3/cFEZj68dDuXIMv5soF6fhoqgMaO9AmjavuPE9rRUm4Z0ppjG
Q5w2HrcXYWQKRTorrVfFWFZKcv2eXDHGufGzW7Cf6uzDsSin2nECABqFSO1Dhyg694BAjgIDMa8b
EbWQ8ZWDMhHWly3G79j/yUEZcjEVaBGqOvIUZGvL4f8JdvK5+f60UwiwuHUKlihdFx4AvKGhcgU9
NSx/TFd4JArBMWaL5Kl8SBDUnVvg5wQ2apJym/ZhfWPYqAzHKgeouha6cyosALijZyYLAJBQGZnP
fT3Jp8UzgcvqaFYt8QLPinYbrBqqTNSnnuO8uqvejFr5cLG2HoP/Hn03Y3gk3sdjtK1Jeg3qK3h4
sm7S7OLZLBq/a6rfdeW+F7sNrEErVvst5IBpVeR/MrHQJZ0trJYqs0ujuq9vIL0/5Gv1fI0BCD+I
f9hGK2EebT8vj/WIva/77499ugwPAKQL/IsYc40f3uCc0d1di/pd94fusrJQpdyi1DnhSozNkVj/
p32xJaU0oN7BxcqywfgxtkN0ZGY+vn1I8Uxftzn7iAch7HCK+yCSTrtSZSnaduE+By4Vat89DiYD
CC3vcYhm2lEvjb03jYB1qwhkpPkyfqg3G95usY7kLvzZfLrPu1KzD1coc5qXIFeR1mzc1LZcQNV2
Wk+miox6uZB64mgA2vxWqoAYCKlufA01KCPf/QnOmeoIKib3QCa3hvAZ4a9YtPTJug0qdlRG1cKF
iy+BAJcmPM4owCyeJTf7yHQ30ZaW2Vo+J+ZX4rfmf4e1frYla61lyQanemBQfclIO4vlQ45bDJ4v
ev2tKkvRLzX7N+6cHWN34neUpbNG31bQvTg00BQrpLiJYccDeK5Rh9d2dFUYyYpPB1m20sCh3fPD
89R8xQ3kNGRgetT1VDjSzD6mIuSTaQFH6pO/cmIT5Yn5wdFJUEZmKJGg0R6r/bCdG6MC+pYZGrwc
UsMxm6aGqVPz8QzlwJwHRVIkS1HMwGJ8+8tOqs1SE6cDlPqd8CFN72peoFZdpBgg/F9ska1aa0kI
u2Wxbg+4HDU9PTmnVCLG8tf2HDIpfRe7gHWQI5SXzLcBFkVpzjZjtDcsFfY/25l8uxOEBD0xbmfk
no41k6qTplkRP6LNyr3+wUprRpP6amy7AijR046FPcaWLecSZz2J0BNLXwLIbEt+91O5e8m7ys/F
wi5PZ9yL93+C37xkKJaubBmtsLnVPvHpZn8WODfeDzushVjOTP8nN4sVMYnZCDRrK5vLrfWzkjsQ
HZOdLb+lUQ1S+0lI1UsIyf2PzyHBRQB9xNfmh1ENQNP4vut3cqg3VDqzqMoGrcQERAFMEvVM3WOZ
W423bAsnfOtu7pR9j3qPNWulOjY6GyIbshcYnO3WjLvEeIYj/OQtVtRs5A/S1TA7K1U4ZqHqmlfz
YDR3HrUqJ7uanmJB7Ls+hLXpG1JNQ0pQfQkSEoN3SPqzrzhMok3l/9iz8AqFE5bqYRzO58CpRcMs
WwoQmLWDNGLq8fD2+KApTJc0+S+6jbjfxMhDTxhOaT74KsbZKQO6jWWwToTTEVU3OzCFCkBjaQN4
zosVFNNnjC4Jl8k9VH8U7B+dLQBD8U9vrehG/C0PueaSFk13A7Rgmxj95t5fl4kuHP6Oz/25zuxU
5QKkH5nZE8iEQlXiJOsMl/HWtYSg1b5oAb+1w6o8vrd5QgxoWIlMQywIAqyOZhJUlYgnDliUxbgE
kdMUC9dMaQxJw+KzLoB7GVd0hBkF3wgfuEQvWYKMVJAeE/Iu6fw37Xu0IDR+9HwFdyiDEd0kUhMM
rkxk+J/tfoQPFucwh1JQngwM6kjuK/C3C+H/5VkPlYNT3zB0LoW8979z+aYK+SXKHgvvYjMt26C8
GPITdPsbJ6yM/rE37SqQvT2rNvpLZWrA+P+xKyPSauwNTWvLl3pBiWllrS9F7lSVk4QyV9hlOjy8
wEVqRRvpK9q7AgGlX9QCDuEQnXUvQpFVfvpSoTgg4OEloMBRaGHSvwEUt2sSsMNM7vqBCg41bbgm
RWYY+oQzNsaAxaFn1bD5PGrR4Y2yUv1XJGedUnk3q1axFsgvIum+H0qAP9erpV1LpdNiUFLIWrAz
IaTAK+DqxzyZsSpb0wHG+TsQdf2YXHwcMhLzBXwazJBiTcFAxo7chr3bFa8Bn3OVonV7Ozil5+Ss
rcKpfWV7NfX1gNaeWOsOf7fw77RkQvd2mV7GQaFl5ARyC78lCV8sldPwwmYDSPcr+2Y060kQAF0R
Bq7jNEiCMUzhtWg+1v2peQp16vhycxi8GBd9daQt12OroOEIN6L8+Em0jxQVeRuuXB5ul3zqH+3u
o1iG6Z6OST6hnH8uHqWILKG9ZiiEeBDGF1RKk9sTMrvRab3uzYfRn0jy5swYc5vrgkPi/42t51L0
/7a7x9YBBTeneGuBdELossddD9HgD3/TUJSzqF1IHRIININLMhURX62l/5pNIBBYZIKv89+dMvEO
PidJOMGH6JkY32nMJyXLDBu0zq7hGQVkcOtK9vfs93Yn7W9I/00MrUls4AzISRtogZ9yJc1wPkgc
l6iARvLR+yx+OllZNI8vfphycHiDbAezkyrpLULZmnDl+PeMxIcIckh3nPhbgKs06AKVv5rYA0eb
BdY47FfWaM7DJaJeTysEyK8wCVIVyuSLABwFRWXLYGy+ZmA28QfubD9nl3A/U9cBbWooq/A9coIM
R9+PiUJT2AbQUUydFn0sfCev0ni0EKtDnOn3olRrXMvw2R8c/dPzWfaFHozIRV9m414ROg14GoOm
Rk9K2l+q0gjTgqGpPnnG/jdpHO7xcmfmRKA/V5I3Alw7UXFz0qI3j34W2iuSUcM+14QAD73aLXXm
rEityAPxqpExu50pormuh8HkBEgNfj8lIHAK+atJzwKiCxzt27gt2dIdlXGV4Ceqn0K+JB9e+rYv
uinWDILRS9Qhnd5Lv8Bh+vfXx5gsC7vYSwM/CkV7y534UEiQUkmqWZoCtpSbuuG0yqPPlvSOZ0EH
cantJ4KOVs1J6N20oa1Mh0/t2zsoLVq9Xg3sYF/6ffFePtG0RazEbUBUrczQY66PgEdZ4HSO06rT
+1Ki20MhzO/riKKC/ZBiBTyu7xUolkOsCOmAvLbioMDfE/5F/nmNpbs9jVRJId6V9/yqZs+qbT+W
qUtSD/8iX/AySjK0blLlR/+EZ6KMSbh2UCC0JINxNYnw8GnZm5JCOo4ExyVV0SiVjNWLW2u8THOi
n59eoA56uzUCZ0n2NCxnBnotLy6bMPtSvRZhrOWs+72fMZMeSbX5Ymn3Pr2pv4LzFHInUwPHZ48b
Tq2iErP1iMCZhEp3535WQGp7FE3AYcy7O6VxphPL3/0iSMKbW3ajUzwmZxWC3URdQbjA5Gtqz/MJ
oJda79XZANfeOXdZjQlrbc7pU2Ab/qQJSuRHGsdaxm0s8RwkEQkJApaxI/GFXVWlWy/J+sNgCIsV
kkz9Y2Rs4AyMRESMU+noIUPzoTBvwfTYAf4SbWAIngGiJRm1NHoF5e3hTNz8kgHS3NZRZp94VkgK
CYFlirUx6OZb/mv6B+y/lHyFzaANcl3glpQz+cLoWinVEVdTnyn2C8CvQRY0mlpLyNJdAWHcMSn+
K87BBpogXJo5Z9xqVnrh9FfHsbjb/lKYQrAszomVcVF0yRMMy7zHeyFgqFTf+cq4Jtqv5y0Dp0Bh
PiuoRkYNUCx2aPj4ByRhhB3BlxzHx0IJdGRELqApE1oAEubPD85NbmpyNrdND/L5rueO1ifAk1oj
2PX9zTDm0N5f5XASi3CcXbKD3tNKvBYCxkGEMrVQYqCGl1BfP1irEdj61lVUfnRZ9fSrSTTbLqw/
8Dp43TA5r8N7fFuOTWxpDn2vlX/JHHv00HBpJPMcK/Mm7FS5kWxJEIzatb3Lzb+unDW85vOK6H6I
j58PZ6fwNxeIUmkEVhOg1z/Ga8BlHNCRDyZ7F8HKMIIuH/2tNAb7ewA+p24uWbSkGi9TgSD2rvGm
x9wqpaPsRiFFJGQgrqzQncwtEupJ5PzTfeb/QdpdjlabQObZORLTUZhrCAKB96p6QTI48sNcq47L
svNTTmeGtcjrhryfmoUavox+XiyrDlZ6T9iW8MUFiQ4VPf9+dAVaeCNazHjWdIWhbquY6c/v9eCj
cI9h7F5xzl7wStOC5uuGkxlTQPuIYkDkxu4H1PWHdH649g6nblpyS/rngQI5xQ4jgcSv2BcayvTB
JecO40kXL1/5JwdoyfVpY/EYLmzpSD43lEhtWZj3336YtqhfAd2WYr35tWL8s+2xpnlQ8j8l77xo
mHChUERnFMpXeMsXKikTYUVsAEtRb5gXqUTWVkjvnCHzDhumVyU0fOcEvQWQ/HjrZRhPlo0l3mxb
eLwCAwlBoJtQNwK8LSyPPhFRp3hqzV2O1sbzj9apfxySufTEeV+nJxDU9l5wx/uJDPVWtp8xBZxp
3b0JYlnwDigHBtibEt9gKo/RhaXuCj+9VUEdHcana1WAQ5g1hhXWZuIW9257UZIUY6Q47BUypqMQ
hJF159w3pijzu85yKTu/4BATG7r5o0ROkzZ+Gexu9RkdEqiionhbtcrOYgqW3zDplv/Hd4piqnRX
w9wcbu+9BWkJZYtpekAOVRAIH//+U8Z4EwPLKFJyaiG62uiatJM8iSsNNX+Q6wCtceQ/pbBC66d5
kina+CArpkGLcd1hhrQuCcQ0GamYxIMM99VAmDxKdtolGXdOP596R1Zn+6ML7D+doMhPa+Jv9R+X
yc5fPBH5+09ow/lveihgLXjLaqvNmvUwUvV+kTkcQ9OJcR36PENwioDc/oTfaCo3Op21eee+a/K6
+mSpai7eoEGHwLuW9/9FVhag0PI/W5zHRZxD4SWPnW4LwseZvCZzsEbHBVhKltbAz2VqX19NbR7e
hd2HKm3ULcp+DgmumKNj6Lh3FMpb0S/BJnUsCAOR4NphAGztRYXmzvo2RdU4GlAveE+0yNTmW/Q6
5RVpQcnwJhNFdmHAnk9vYBxoIgVzBP20jfcWFSpE+vQmwA3yQ1cHRXHlKqucqVg8nBv12aLFUUF2
Jb1ZkFWaE1mP8XHsJhcabe0OqeJvhL/ZJ9jAWsxVOkDOsYYSsjR9bqznoA5IMHN1Ahc/9NZLf8OP
LgGrVYgJgfd2YPjwLv33BqGVzX86c4YDNyhU2djTU/yMqXvj+wstHSM3QPGpe5fuSrZN2vYAAn5J
iOyliezv2FEr2rHBK0vQx5SuL6v4x+T1zJqSSXFuyCvN0wq5PjcRIKOAHGeCMiY9vFxAwx0ptIA9
PK6x6BYY7Y4LHmK+mjmMNcBQj1q6pnmVL5gkoB1ApsuUcMBlevnRCMJswfzJf+DI/R7u9CCRCoxR
0gBlAroIphQVK6t/b0MPtZxE+nydERyA9MYGLB4qIDsDoPIXGK+byL1WzP2gmPup0SwBD9FnoDUT
cOu2QvKz0uwRjG4IkccIMDGTegBeKm2GxawcDt4TWnyfD8y9sG9xSv5jweJ9VX2E9n5SKqeiNDnk
qiGl2CtyFcdsloJx4PUXJshCk7F7q9C+nNcIU6I8fZ36+VkAyDO7MxzuoH2GkDwxuPzL4hdE3uG5
Ej2g2JQgAtqJRBL5f7+FPZ4hX9SEr9YBu3OXxOuEsamzvSj1su0/hiZikSHNJ6wvOXyMhsohzQjv
Nq7MBA4QtWS0DtogjwGqSqOcMCiHLxmIpOnWTJt2SGEqjYo5864Yux08+Qv18Hsib7zSDGgtT9sa
Txnv9DzfAoAhPt2UKkYJqAkKfPHm5WRYyJRuPYbnhViYkeucdR/RCN317r6Ii+ig47QQDtHjCC/C
IQ/3oVoKlQToW3rHCQEw8U/uPZT7LsqCJLibXgSLUGArmtv3A40wr8aZKCL/RubHFWV0hfPVZAB4
GrvUq5rqSXyw7Rfw7de9xfWTgRBdbK+DXWQUaZvD/GNBs2cGbcOWvvHJicwU4tu+jN+EtQwNSTVV
MUgOuWUd7Pijl2bBafJ9PCPGDsMp94p23HHdmWwQZDxxAmi9PSieqp6z/6pP7tUy128ohDiex4LH
F7BmiaznbATHPZK/1D6/TR+G09epgsvIarSm4+UUYBBHwXw21pYnRTVne4dGAHFdZdgL7V8W/pFp
fX9SYg5R8Y3ieKTDWi1kYE4lDutlfqxio+UdH3goK7DOcXJgxP+BNuHyy5DOVDN6Jjw0rNqZi++x
GtqBcJ01ARCWjqqqL12zAYsfTxcUxhqTDK5lTC+X0GESC+Tm3NDIasusAgpX9zFGV4RZc9J11lEN
fXoCamA4YJupviUVhdOUOrEmVx811/B8rtV8pdNfgxGkQxKoaV80rqKcQJPfopHcCw1IVDOEETdh
3y/wIRZyLEDSyFSEnIJ8NGNs8ClieV68Olj5NsFpSK+4pcSZyAfK4fPjsDZbfm7a1m5Z3mkOhizZ
uJ2tLl7aO89raXxOlJWQY0C68qjaR22virjiYG33qf/7V+W/e96zxSmQeMGFPkbr2iStd6yuhx7M
NjqwV+XioRqHl9eN+u4CXVmKp0zP/TWnfCaSOJJp7E96Zy9ZTbHfLLYuAf93wqkIe7PB804ZhiSe
c3Ta1He8isn6hBjPaVv5OG2locZq0zY5WDNQJLPZfiJjOvWa54g5m89T9xSRi2NCPgizCxzDVCmk
MyKinXKBZ4vXMUKMZkpQPji5qOIiOR+ztZeQky9qFJhpCLVZEeHSxRHi7hf7Qtalw+kyoxOAC1Qb
G4lMzdypP8BdMOeYc7WeXHi/UBL9wVMnz61z/jH/xDoJVXAnMxqFMEU3heNAkD/80kK7te3fEUFa
7SJ9YFwr0ZW5dBl/rMupLDYIJKm2fwXJD9QC/AgCjeZgzFykOItWwYRA1M1PmVkh9++ZOGzfboUj
Oks0Nx8kOBasulOiiA/wdLF0nltcZkjAzKbmn6hpyFadZXml4yhizFJnx6SjJl/KWbR2QCyzSbYB
9Mx5gMW83ECGY6+B3NU0W1hBqjvL3ygQSokC3/lwcs/WTp4aotJnNnZUSa9eq9ZkZZ+ofYG703uM
K52kihw085GvJ4GhCRoyTaIDrjJ9ht8nvsgnGyMJsUhfPFTj92vZdUqgsKIQzx2uhyvSmaE+bKP4
80nOQEULo4PNqzB35ghEthmyn1QOpFBLFuRx0QjvzSn0vrCeE0T2Aj6xcUMTa2MISsdl6s+iRcPo
xRTABKuYc/SqIGp/fLTgd45KDiEN4eVJVXkTYExvuQudLXnnvf4NcKTR3w3PxKwPa9JwtfztO7I2
9m2RU1MBIPH74GpuIK5N3hC6skVR46d+MyU6iMkBYbx6NJ6AV/Jif7eueIShquXVPqK1483z5xII
zXeUe3RL9BKz3qOavavst5eUeTrRjT9e7cBj6hleAu9n2P90wlltgugOql+SI+ldjwFZu7q+mj/0
Aqh93oUcJhxUdJ/Kq4aM9W9uaQPPuV8IC1mTUqjb2hC0/O3CgF2V0Jf9Sw/uiicq6tPgv9dmuWu0
f9R4Ne5dygwpcM/VEPjcXgFFWTQp96cVM88b7lCSQ73zC8pWTcYP2Zf79bZxe9ibAeZdtvad9Drn
oxHzSbubQT7uTvJkvBCQE7qodrMLvJxHu4HtzDED6oiLso0EnkL3EWmzjN1mDQ6livdc1ZXtCl8B
sLSEqSWmfbAyy4Vo7E8UpYaLdXXsCmY7362HMwfRhEV96/hGfmO48zcHKZTnoisXZzT12P4fWNLc
R8tmphGx45kqHPUOEz26z65aZaqUtNqe2GdxvhvZ+wZCb8YfvbGfQZagXNBqRQUWyQByq5W+Femh
MunREc42ZdFk2y4dSQQvy/vgHykCAcb46U7Rh8eJRaRv8qOyZFlE3XAYkOufQkLVuAcEjrYeYFMa
VvXvtfDfAKApWFEVP7DWKioS/0FHUul8dM2hGiDnguq8gryX0I0JPSO9oqhUnQNPvSa4jbcdDDuj
fArrS1/6AXEWvGMBytWKvZZp5QQi/+LJRseA+iU46/UAiOsHVlH2UVHwGuMhIZQf2LgjTArGHBmR
mXWl4Ryf3d1y0KJmlQAY5WO8at2J8/+DwZPKqhgFxqJK+9bQGNQi9amcRudIcFQrzLQF8wSrd3u4
EkQfccSvWCmOyuhi9Ko67Z0XGYv9DHCEir60WjI84dKnKNZJ73dBR6ApqE39ERtKA10ut04kXeEP
VXTIsWkQ/XcyB+uAbizxsVG0vR0WwhLUh2EWoDAGnLW19eBpycsJFstef0tu1PI5L/EcbECiI+cF
pw/IjyTgz4KWhZDoOumywMzH/z+gIs5g5lzHMYx2RtRl83Sa9k/El74EPibu7XcDfYKRShHO4vlq
rZDkrTaz5pumHN9dtbkRU3SePqFPTDi0UcJXixgmxVUTCv4WG9w53EBYN9F4s7mkwrS/C090p5hn
ipl3gvinCUJKuxV6DiTYRGjtQDi00V2dT4DUuOQILoVlolGGfJ0+LVXbIXaq3yXulTzdf5WOuF4i
Tg4RXUF7GZKepXZXj5QWwRMogU6P+B9Y02CUnYKo1RQzDND6TaIN3U3wQQbo7UWvQaBB9dv7Ov6c
y2DYz0QVaLf7x36CLx6L4VJv4smSA45Rt1oLiK/loI7oo2vrix99zBZCcVMhGBnnnznEOZAW5DvW
ZWhs2Gp+fov0EJrS0IH50bHZ4wDT6jrvZJwtTh2BG6wRxZZJJO+LNgCWOD314j+PNtFWGLlATALn
BvF63cVvAad57/e/i/iHXg2gst9Dhs07mYmh2cWDIhShMh6DQnPqzJBynqVWHJdQAjHoY7YTxUAC
vuitW5ri4Wb+4AF3oYaniWPU4Kh4XxnjCUQgC4THzV0oDzCtrnKS5iHOxo4Ey/RwHwV45P0PAiwt
eQ3RVT2SX+cpIIExs0OmEXWfj003gQFH3aE2WBBf7uTDpPNlIv4WeF5myON+JPqksLyZNNOETZzo
KYVplyyIYKexJN27T7A4kdCP3BfS/g6p86UBdm0G4tZGvrZimg+6cDvVpkcC/PbkmIp0u4iBPNc3
ZoONN0Da6LfQIMT6kUjd2cOICRZI7DerQzq3RTOfD9qh8LhgsPlzb7EYkGqCBpAP8I8LMITv+Qsw
avrVHbS5Ib71JuWFjvRwuoeiQF+RisxmthnX0wpUXgB9LKWXu7CkYqwpTr53R2LwfJXTF0Xv6ii+
kYesrSw7rTVNCGWhBkQ7HbCg1TipG3x8YTGQMZ+3ldD76HwfBrAYoW2CX8QY+F+MZLx0sPP1abK+
9LFVn+k7eieuxBHycW+QIJnFNgTA4CEzAhZ1ezSi19uYB9jJ7CP45Hd4R3mSyrdYZkEsmgUaCOSz
azOj9TFiilScLOpcWP0Kx7+Sx5ZgraiWicrbsNn32C4U/Mn6PPevW4w+Qk6EGYWa0F56QP+xX6Bj
5+Fnpz5wSzhhWD30/UlskGsOABv2/hkpOrtHBXDGkjBd7ah2k/qjYVvXowuX1j2UUM8FHXxd1ZmO
BKQUh0wnjtij2wneZDMEq5vAJlzy3q1N0e1qLlxxNKIfcWPGzU1UeBcpJLsKJnclVmX3jJEbkJNm
AyOQ9Q3vPUPKXzA97kYfnWsNsM7PK92BvWBmbuCawclfbk8WHR5Qvg0Rj82T9X3HNAe9FQVpWqPE
6Cz3ISZ7CdLX4Le9INz90jqc10pi840P85FXjtaOHDzYDs9U1axSiObmwjdt8rGGxN3hYR0KaOn8
11Y062/qjVEyC8d+B0+G0X65vK7DQn/dArx6Z2m4dieJ9LoiYSndA2sqv/WSkdqzUPb6FujWOHiY
rp5pDpjkQzHdfzqByHQyPcRUNU10pMyCany1Wpii8+s6cQJv1glSN8JYq58tqTdiKkABSTIidnfl
OycIi0vt3L467q+wliNXsFOjNaI04HPELfos/L6skXHKv3mt20ZUV7Q4Rzuz8WNslUx/QVZD3bCJ
1IAGrpDCuLLH6qNel1j0S8PdsVOwbtS62WFIBrTXgnD1w4463OhBqFORX3id1aJL2nODRbF8wOZj
K1l13HizR1xCI5pIEAMIHZvPVPud1dEEh2nW+JKJ/72LcAzL5vcKMeVXk835v4qErD1gxdbI7IXw
tGbRxtMOB4AweTrAYlYimoQszmVPm9RtR6cv5qTLx7Kl8o28vgVUNR/M+c+u4yBBFK5nZH1vrLqe
ciDi7htErQMQkZ0WwGjpzx3i1c9Ts0Z4vwDyY/VW6i1aMaBqzkTM3gbUfxhs100AcnlGGksjeX3b
dqkBcK4PHLm4U2SEJRDZblLpaQSw6uRKdg3R6mqQyt3p86LtDS9fkFdFzOpSgyMz7YXZkGVNGs9u
dIpvHcfVnjIDkXeUGN6kx3mLp0QAn15UeLy/0I4JSt/11V+45blccM7HHM2xo6JYPb+z6kR/aLun
LUo4KkTxGdjl+rSbD0e87M+kIb8AKE29Fu5CBHyccsVJRNqRa6G36UkHiEqtLD+PsP71nwo8DtGs
qi0qPdzftQ5SdvZaXwcC0SE0if1zNVfTZOjMLyqnliPniIvCrli3YVa8vkmDedx/b/1hpP+fZJBl
1GGFESLiGqE+Iwl1VHIYxu//qi7NqK2gEksyAD5txM1O+02jacJXC+B7SaH1Gnzr9NsM4SWGwILA
DoYDumPO6rfhh0SbHW9dxRDOfK+aHh7uhNFfde7/IvzalscIL8mB/TvUJljkN8AmNYAVhy+JT9ph
pFwCtzRoFILP/1lCocz8sSp7SE03WcReCTNvTHTrH+BlSIU2Vj2YgnsG9uHtM7musj4Qtgp4nAjm
UywFIn2UvWEv2CNNjAtlfQl+muQv5jY2LOhNvsujeO61Wv5UZu0nMR14hBzKSfvEM8P366+yy1q1
5gyr4uhs2krs93L1b4IfK0+LPo6kjk6pt7bZb5zmmeLUAwNMqugQGiD1V5Qf1ara9FBxNwEEnqQQ
NFH1uGCUi75SLtHsiVtdbNHGVnNMKUVNNlfP4npVk8m+IZZ566n0B3s5F6pu1bAmshbQOz4wLhaw
1h1rM0tEsCw3488H0BvSwgkn08CW7ALDBO/sa+n2/gQtH/M4S+LV91LVJI4iXTID/QydJBQPh3cA
1+cVHO4cw3y8uNg9V0an4s/QbztczEsL7ohgow6K7QNouu0Qasn+w7HTMiO15xzoFSpoHWxAjAMd
eDiFdFwNyYedTLE/Ob/oURxx/uKXmJgvisP2KRM+ICoVtz7+QJfT9gO3Jm2mHaOMHwdKk38xgba8
BhtblsHzNdIv0l5Bp56UTSX+Znnhz/cew/X3lSZcuktiGt3bgEC1ul+PC7OFZLnz2vc8UcnFOTlw
sT/a9czShH2t3RI8gRjU/CHRYHR/T+KBF6OLK4YS8hNaZdf0NMA9O0AlW1EtWNwH5F5n/smPXMH7
Q1odEf2sARFZBgLoAghIkTQgJc9vCmMmcFYXQNw1IegzWNYJU61r8Mv5H8GYOHpi99j7GO5NyVOK
i1+FVDP4aU8uB3V05wbA9S4tIyn9AMfwfHH4t/RWD9K6Qu43r9g9e7HxRg6oJvvVSjryg5Q6XdOM
b+qUIeThEwjMt5roh3c7YirF7BIC0Xi4R8mk7/uG9+Sy9wPxxzjO4PZ2du3X0cRlDTrFF278KNfK
RSPgOvaq/N4oweTfpMqO0jkAK9h2nme+Zmi20GlfoOceloxnKmhFLH66682S64jx37mzGEB5eBuw
DpjhIMQULmmrCGoMlzQ2kSvINzIu3nRPMg/KEoq0iBULUz4GMSyiFQxUN/qDrwKRpgrYD28GZeHI
SAx25oZE2PslfByX59ejZs0GB6X6WeISV1Ur4skUkLS0Pt10LdGY2t7jSnCcpuP11l43AdmqxIPs
HCh/gCCiRjrj0j2xuvTpvGdi8Zf+ccj4y7HiI8SJ8G4VN1xAuFbenMrGCxedIDYYdBxNymSp/EyN
0Np0Zyo4/G0uJNd8hMvmXlWEOR1fqK5sODG2b4m1PqgGA1Qpiw3L6eN+zAUVqgUI6ZxJl6gG7aeh
7GC8t3lxZ14ckocHZJ6/qYIXs1juCvkCyaKzAYmcd3ZEucm4OxAfPdmNf9TgPrC1pwxnJMtCNijJ
e8rLRb/8MxZKOf+gUkYvzxlu04zqUGiaFtVCUgCtKBolWEVHvh/GhXLlst2dkpOWqNioMvv/I8Jp
IXrM/QgjWnMUByZ9PAc//RbCIiXSGYQGFz+3uLXdlj4JNEA/tMD8eTXRv5fhPgb4MIk5Kqul5xQ4
vhDcbEQ1FQjrvXQLA5zy8Eh/f2GTeRPt5Ba5H7KAqw5bGEasfQpMbZYRY4QADKY9fJyBUp6zCfSC
Yu0GymAvU3Ngz2XHtaCc/EWQuOhV0zPghNJAuSSlB8fbCqy9jvDJHbEpS8mfyz2D+aCs12nB1Za5
+f4TN221gYLdBBxA4uUYr3S+V23lOGEchw2rHATBPIgW8c0KqsBCsswST6f7Nm/y0kblT0v+N1AZ
+C/pVykedhaK7xXmqtZPnoz0qmrz8+8KuCn596VyG0uD0dpFKPg5IeZKJ5z85ICO+VNus0eFJN8W
OwYVYmrHCZ9iXPINERNRdw5DTM6RrvNbN/KGvPIJMkxOvaE6wvozZCNrmtpsg58tZB/mdrEGRgMX
DTpP5QMGZBxfi0+XZJzfcfTZQtyrbywhGu2Fjr79DJiBFfd/ecUsmgzVgtQq+coijSH78KZrEwUR
j8aV4Aa5eQc7vMPABSknvsZcni/RhHQ63Ki6v4GLKFsBzxz9owPh6FKwD4R1AAq2WRCezxXLvkSV
NhUr+R2XCrWnhFsabmUtcFkDy0B3zL1Gcl5ATG7YsZuWgopJj7HvpcSTSHCF79KISgHpr0VqNa1r
9AoaLdjWDyvw3b4olm3SXsZzzrvrdI1jf0tUM1qz86Lk5vusjLnV8cJd84fGpvhF8wUU8//naqK5
GcghCsEqT67igPMabfGmkB9JQ+D7sPLRGkljYauCz5sOakJizeMweZD+RlotUDXQn5vkS31QSe/b
D1E9fQ+j/aMmIKWCh9jO0KNVVW2zPDHmrw5lqowk8/YZNAmY43LVicsMEGTAWXl1XR2+J8zL4y5+
tFlhYXe2a/OtMWCXsBFPa3SRhE0f3dZOWfazw5AS80satfnTYa/5MC+qWaMVvM14lG4aqwJyAfM3
LNObgKNkB6jbePI167m3CQW0c+rXguvucWyOF4Ls5heSX8+Muu+bs+8/qbNTxLtgPEaT0hCNMS0I
bAKIDFmwSow32rKy/PsfX+G1aHWk5O3Z5qNvgm80MFc8meWttGFVcGKghaeXU79OVW99vn9bgfl6
KF62luH7yrIujyEX85KUPh2INtnZ1q32Yy1wvkLDKWgqsBx2X0cZzBMPRwHRDF2irqRmkyYftImr
fEZbwWDbQgyGom4YVs5vsIQ+BOi5wypbGQF/OdrxoKP4iKscFG2Qfv9942oDZ6WrPSFK4LXPT06L
jEeTf2khsSGtye+KOxarISnd1eWi7unOhZlKvs1TyhpGb23hzxnYGvWGbavRYEfZEdPT230sgaWn
OY/yf8jeOfHzvJbL7RSx7omO2/8h1UeC85OABKahVP5QJFUpBZRJk8o7NCjNupNc9bF0uAQaPl/y
yqNZLovPrmn0qA7dq9K+eYTUryqN+x7csF5F7xot9B18xWcReqmI00jh9xkS02hfqhU7AWBZZdmo
BGNyau03mXBzMAnvTYHHlV3R7rGrDTrh6YZ3JiuXEP1u75WT86H1b/OsZNCxxkPsN3M6dqPMcJzQ
+zI+pRLN92o4UgualVmSlvvgFqYTy2cKG+QoHp6iWK5OLZZQb9NG0geKGFSaXPmwVaD0vVfwADCV
LH207aPNxKEbf313WfEqvNkyJI0sjmXx6AVfK6NfmFV/NwfBF5Q54b/YV+9fMOL8fHsOn4UIbDGy
XFx+iHwaHeZNWelqt973n5vw+y64bJz8Utfx0cMmmDo23K8cbt02OBwAag9fEAx14/ng8x5+A1fQ
fUaSo2YkANFqx/FQ4j90uQ/wt7V0OGWwvqlQyri37SI32ydhsOYZSxdG54mWd8mmja4NcrMYseBs
70/OMczLrFiLk1ayvh5ArDgkgWDPvQAQUNYdRkQEjoX4D/d4ZLwo7nEaoooAfVRZ93GcC6MkVvPG
H5wDXmI63vI7jeijVwG58DDIHzSQuvo4QpHZ+1zc7Oh34wNGwsqCQRC+foiMcLdr7eLLCR5vgMKH
lAb8LnNxLYmlnPGEeLXD2wE0ORHWfNMXvzT8JHhEm6Pui1be3IFfEavkIG1uRKDQK6KwEDlI7m3z
/mShHVmHtYk1hmt4Hrvsffj7FKka4VZ04/LYXxUAYZU/eAsKEOf3ZH5U12hebnY+iKve/aZsKpXv
21xniqZvCdYqpZtS4uPSd1+/LAk4j5NWwQW2R8pZogxO9XbQXYCu5NFwfZGuTvTGxTD0Gnq/fEDq
poO3UxmD73pxR6S6XKrOtiN4xELSqXpQQls5ivl31v9EeIB6h7XlNNSueo+NQBcKNFJkQn9l4rBB
N4GDCG7jI/sxsy0M51oUxPmSIugpd0V/u9ACJhR3UT2rlJvd5mhXF2Z1jAF8/aCQJTspFIj0Erpn
7io9/VqNe7BUVV+rLQcI+zKTOD2wogOIHnvQCwf85koGFUW5okKQPwyPD9frwa2w9920CtNyul8Y
dbfu3laHM/0SbfUbe+i/69hjQI9xbbfCgBGXuNH9LEXDFxHjm9ZM09UPSSD6gyMAG/mcp7qEa7d3
tnJIHnaJK3J38vKmEVrBgqLKSjal8ewqI2Aij77rGjxqYCcihkWquvPZcFk9vTX9HsIZsk8Hupz5
yrN9ZjxEixaXP976ZZBxmdd92v2LSCU1A0d0xGmK8fILfnefsbNledaoCuL+cGlPQ6dTpevRgHEU
SbUzymcWRTop67nP11L/4OEbBUfC3kOYvkmQKpVOatSVAjdAdPJx6A0ik5QlCSIT647jzw4aH2bu
l7aiRU38sKns1tYwXLuRbcTxZ4p/6ywcSy3AtPaGXhAvj2zBGUwxIgiyCEvm1McFyoRau/XhiCvj
RNulPdAkDaNTB0RddXTwdxWcaBVe3UEl2bUyQ51H6j7Z4K0TZmOLOrKtKc3ch7Zzf3q2EkHl21qo
XOMgYXjO/YjBi1/WtylkI3oBTMx4+iUWgIZYbpNf1Ou+BEm492JIVZlws0IL62j3t459OMpkZyI6
FzU/MTyEfDnCW3NRBrUn4A0gURuT2SUQk/hhW33m4l9deUZBZsSbOK/DEKPyth2FefcO61prYkIz
fraiLWxirz5DkaUY7UJr355DYbzZx1D+wiHk+PuYazE8kIAaVan3DWt9IfOD//MF0yP79Q6F54c3
G7xJ574Re35f3gaVvoorb1Hpt1qLotj5fzgUx4Rx9vNZQA8jPssuryvRxhIvgzMtIKdsC0RGXoOu
uIV05aqSiaApDXWqTqHB8O5NBVGwZ1ATEOOGfmpSvGgvNyXj7+0dCss1F7PRYXoYl3bOpU9tHqKr
eVehuH2krowgelzXzv9A5/A2aMWQxGTChPXYPvIEjCH/h8eO+jwNSlsmLtCem+ipwaCLefTA8QL2
jUzejY+7VFYYnLWYpRKldQ6+xuwPWrLBqjAZNkPcjAjgInalFbMx1SQeDYvBSTxrs1fKIezRQcqD
cxfdODT1RnNastDNscJMK1wEztXdAHwk0U76HBJVKBByXKaxgJkoJ3iVAxgFsQ2ZDx1E6El0src0
h2bzW7Fh7xs1joHczFUQ/VJsMRN/dzUG6hUdx50WnOznr6cCpLxBEXthbvhZBpT480o7Nv6yDEuF
ja2kg+6IW6usdsfuNgrFFa9ZrtmgbTvlgzUujVK5/u5c9GIvgnZAl6CRDljoFerImCGYnlOr6EO9
tUG32+gqA1fpKoZ4A1kzLqP3t5oiRFIqCuZoU5ipj6e9eE6QlEz4se/RDMD2zFWTPDbWrcuZ3GCT
VncdxZgQopxgF55Hh/1hHWlz6VJmOU2LQnY5AN/NBdxMji59RTIjNH2l4maOOhID3VCNzR/G2LHu
zriEkzABDTpAJyK8nOoBrXc2CXHCdTYKWOZUR1P3Wkc9iYnJfYhYeBX5JFs0JJW2zAqTuzPFOmNb
GVSAz1D/yMWqMg1npjOB6dcPL+NR+zUrnAHpZCA8R10EuNN4yq1UQtTwvHcl+5kZPwBuO4hYoGnm
eaF6BEhzy1oY+psFh7M1sFnE9GQG5Rxd9/QFQyrM/LKU7iGwbyy5YPMDqVXEODeRyUyDyLv5Wlu5
v6UTw9Fy7JVNrZTiJxDU9YxOKtaNLkfO+Yk4bv/taOUFz4soC4FZXjybLBrrwH66frFt2hnhx2lR
Pr7mx+hSU/vBVi6Ryc/9GF30uNDVrcjG9tbvQOandmeCQFZP/1yiDLc0BN4FnwW3yaeCZkKyaOZE
X6QHw6IvbHnUqayHS1yn/zUjctV1EKz2KzNdQwZQwCVoxgcA/0TfKjTkq3kw+3O71vuAEnbfHmOs
3U5/EdpLSowoGAKAq58z/2VBoUAmD5EJw3XhJdIyv61V59znKbECdvDkd+DgbYDaknaInKD9h5q4
oB2Wm+MdlE1OEw7k6lWpx1DjCIVCW+Q5tLfUD80CQXHQF0opKczgCVrjFrop2tr4eawSiqJK7vuA
n9kIpfJx1PMjdcdFGVRZMxMBKEURfpkHSOoICSuw9jM/kPGjKxKNxWqbG0gB/suS/AxcvbRhpAL5
vMe1NBIokRrivzEDX/ZP9cTM3NJIQyi/IQbISXX72L+A8qiPLGYuGV05lefwVmBaWkxfE/UI92h/
UNs0fwe0qmy7Fts4Alermq3a7ysVX0ew+18Wi7CdFssB2WnDRCZD5i9HQWmtr7uPXy1AVUPbuNo5
niKRksd/5MSWvs24jAsSgtxFXX41vHRO3PwLOy699TDSQtXhszXWXjeDsnumHP2Uev3PmM/P0ptD
RoO2DyITzn++8CQMuOQQOatC7msQlvBw9+/mJVSqtAwl2ayUfpvveVek2xbkUc4cs4T5h7Z5Cuay
e6+gVZ44p2ueB6QBcZ1BmUTKvDNOPDMtBO+21mSylMj88Z0xVD23sp2vQcjf2L2eNHO1g/AI97wo
BAoPCqCrKW/A4GNgVaxfWAjAX+RnVgIILbIvqSCOhfcf+lDH5tOz61Ia1As88QK/oKoBq8UEAZcJ
tTXx2YI3UbLNz4u3rHmYSIumNgFcD5XIYhNelI1vo+7z3n6Hn7f1RlcJPczm6/VNTbEQEMZy66qt
NrLHGOQPBDWwfJ5+2se9V92y5UEVSS9diPYA+gR7/HLADJwtI0fCAKk0eaeDri9y+ry14hKk+Son
P11VeRa4ZXDlywdjLfr5qvuY27MNYA+xidE3XkgrSHcSXl7vxINCifZAHF6Bgs9EZRXE6gbcvFc9
SVwAOVe64W0W5vXfUEXbxzCC0Z4sYsQcjaSVogaLezCkL/fjliK+YmGwSzsGiDyYSfhYCBru8a7X
cqESdNIkJQK80eOx7KwBPvbX02KrcehbxvdOOH3EmdzgbGQ/SayAwmqKNO7Z5LcLQW4gmILBkZc3
7ddy5NV5wUDqqfPxAypprDK2pNWMDU/fEzfAPB2SUGu8emM5rtFBm3MNuX50L8qwYECDvW4k18s7
Yo38y/xCaqVi2igQU0A8yJdFJMPrYNWKuDXLt6CrjjiPZ/H8iVjBKlegL04Tt1McVaPHli0zQLRP
+HYlLSGZcZAtTGIzmKlbUPMlbZb5qamnsM6+WDi1uQKV540bkbnPjAcSLciR4cYNSZ2eMS/I0U5b
hRe+4KVjBgmIr/F76+ivxeua67b2PynbWOxfWsf1UWIQWwSzcM0A9uZWkHWkxTifraQaidSLwQGY
TQ0Rgd2A5vzXvSp6mzZ71izg7RzX3DPZdCgJqNIpUGQQ60k+etUK1uWbT29MkR8XAPojWNXqRpFF
SHZS+Kzj4J5KYX7QbZ2kv2toJD2uemKVolIJMpx2KKQKm3PC7FlgNLNZRtHcxzBBHYjOWhbZh/U+
RvrjUcabAJGxhc0avVfiNv7mL0j6IMFXFcqiC37gbL4qaOu3p9LncDjoAnVXBBNncY7Gj6jYAYK/
xPzGH2uzoTQkIJTU8T6YWQgbS39IjinlBZ/cuHz15Lm5biJgzKcqxEfOWDw+R19QI3CsJ0sSuH0A
m71V+va+HCY0H/rdCf3DXQuiR+wRqnveY4fDBKRAXnmt+WdrA/K2WWwVB33beqM9+wbiU1szejey
rOxEsQCeN/rPPkVz94u5EGxv5jB/URIGunu4c5C6OdQyJOa+mE0nTn9jTUp3ao0Q0fxhK4y9yDAv
nvEDdZyPcvAGmqYrUn4U1l7mS4rEXB2LjgxkTBfDGHlA9WtEjjKxiHMhHwABPjTSuYVGydtpDRFC
W0xGIzIUPIFcEKUcCpPC5rM/31rKb7kgjZSWLcJj3GbpADw/3Ifi4uw4L7k9eroLPeYzDx9+jJ3Y
8FlWiw2Wk43k1F4FaABwra3hbbvHFk6G29FuyRcLUhMSP1Opv9BXb7Y/aiCxiEZqbkDlHVos3GRo
+PPUdVkaHPQUgleQRLoIM3EclV1I4xgfXKoDeM6AA8v8BNyClX/5FFfxYtI8/dbw5o58Tt4iQkAm
/H00NutSgPj/XnW1FkCpfPR+bNd2Qr9sOyAtQniHpmobwCQzbK6gxPVHDiJQgLlf77FNfW5FuivM
+9wYiYaN0rT5Dmjt+M9a0J9eENDiBMRF+oOjoytfdELh+v0PtKAtdPJThe4sciiCsdA656s+ZGhS
82U7Gdd7vlBlQt2k2wbaWr8vLgrcVAF/UzRlR2k0wIQDzML7KloX/pDUb20prDzBeH/K7lR5sa7+
kmbI1OOqbvWqbBcckJKIzDIpU+hBIWtCvn4xn0JAnqGOVoNz+Ckxnc/PrCFXlw6tcRailHBpWwVi
i05WitpG7DMRLNt2i1TDQkEC3ZtQr3EENYKfSBpX629twrXfr0uBWHsDVT6WorgEilV44M7umAmp
Kg2zmVf5HRMfbHl0S7dg4aTPv646KL/FVJiNi07AiP/6CFHPHLFDiqVUjrVrBvUBoIo1rJ6+mOJq
8M9DbFxKmbCu1xt6m2BnVdglZvTHlHn0nzJcaABY0uayEsNZvHE5FHsKaOg3f4Of93jd54riNQIb
fJUhq7ZUS9fdyE6vZ1mNqy2vF7eW2p1xfPGvksK4KKn7are7QvGadOH9tt2FbERa2j/eEKMpD9Iz
kETHBB10c2URJKJNACKWTdVJvHR8JWHvBo+hqPZiyHnc9LWN6H1Wg8c6cFeO/1YFgxe69fK1HrWW
GOaD9Qji7XLKL8JKz1DEIUn7+txMbbCcSe8JN3/wbnj7OYQLmlmG47IoW4pOFpoV4js4WqmCcDJi
6R2acw/QT7MvK3yEK4qRN8CRhXdRvy+xUgpUtPdLtCbIR3BcT5zPE7R3FM6FGQAocz8ZovmI2m34
LoNS+nvZ3dV3Xm2qqfyCaIGm5moTJmEJCN22McFbCA5qhUZomVa5W36Rwh00cQ+3mKe/FiIW215L
nGECxowzhE9RIgcqSxJnGtkquNF7fA7QvM8yPpfU7/6Lcmt0px0gxgVDfSAik2yGaOIgC8xF2lqz
gnLzQffWXQQROpx8aZsuI5ho/vjyx3SyLBi/udkmUEEH1Bm2g4dA0z5yE0PhFQTzr/zNu/ies/8X
sEdUyiWqSDdcwcwux1+qsHxXxXD8+BVTg2HRHarQLx/BQOqmkmPpsWGRlhs1dm8oiPUrHy9gT0zW
tQ9/jU6jM5/EyM0f1tiMk2IwDxvm+KP57u3VpTXgo/70NGXQT7qOg0zx4uyxsPP8qY61k0rnXiXx
E2BCaKowgacTlj6F1u21/Euc8DjXKvOl2Mdh4vSqplKPTlb7KC1ehIFHolwO2EngxqYUk6ChmzNC
40lpe9dpbUtXH8kG3i2aAp2ZEXtLIne60vw1CxX2Lpu/D5d6wQW2wvwI2DCKQ4K+5D14mLfTyoML
OLNp6ksp0/D80Qz33ZQ2l4oO2c7E/77ULvXOxvBVJ6Dq3NDDM7Rr0ZzzL8ySgjjlY9kuDb5GEHIl
bulVVwhnZTNIsiLSL9rT+HrW17BsMt7FRw2wu4r0bG+KiJtXErGjLgjrxH8iuNHRGsM3rQQTWsVh
8OykWUJtPX9zuQyZrWHc0CSPiTzdRUm2JyB/nOB0xt8tKsY2Qfo5BMOxxHUZD9Vs2QONWDkBd0NM
1ZjG1qLL81XBuVN2lLFMcOClJs+wAI/maJciow8XRoaBD2rfcp/PGt48iik4PcBmhXRvbfsEFs2w
ZTLE7CfiSIUp7RuZ+d96vYDlnKqgaR6UulIqNI0s0YHK4FwOgmNuhmUeuW52nUQA1954a+WULspp
OR4zUl6Ii6mWBo7buRP6FLqZdHeB6UdfZ6RgQhAKmCWxWBMksbhQHRbuKYW32NvKH31OZjV2AO8D
EjQgCBO75EYwBpmAfFPLgts7SjjX0HDe27R+Sjl4AbJ5kElr7lco9+KHQ8UGT+0SRC6UrghHei5z
Ah/jSddkf+aaGuBaXFa+tkyeFsxcLV3A41oPxyfcrtetVFvfZjsiwHaSM17JQ3+UMegVybh+rTBo
9xmQ/kyy/IlIavgXYB7fSRStVLguPkVNsJbxRDX3OSm8X6YDYQ47pvUKK07lkYCQVQtXhk7l0g2n
2prpVn/peMx/E2yRXpQ9dtKjaOBY8VejjR2oZRg3nrghSr8+fU2u3ljLJl6tAoQn4JfItKkTKYNh
ELGx+S2oEtvbjA0La+YOBLem7AYNzvfzQNMJxYliYgkoaAjs6F3BKTt4LPdeWSmQ+ykuQxB8eAEC
1FH4lRH4qwW+CZJ424dF/9EcNidVRJJjr8+Kgm0HgEtF66+Vykyhu1ei9QRC2Pm+R2eVEpQimzlV
HHZEQ/IT5laAed1JOkEVZoVRvtvH+lckIzfcY7HhbUdBjUoHFFXjFh7Uras1Elx9UXloagwIwFYp
ssq1Nf78eT0K+WV7kNmzV5eg1uq/aaiuvbCOtYr0UgAsOs4c3ZlVDrsOhSWRodHiNUBsaEDGP06u
xUy91317u014OXAVCNUM1ax9QLir6jS3tXZFiXJYSmjGnEh1jt6IJ4IlinTJg9iVIehCfOW4xO7x
MkY+L1QJ91gjFJdaRxZtmQaH+R6Sf6PRGBDgEBg5lFFM5VplkyA90U4UKkvPIYrkUqesTLS1X9Ws
Z+IHtqYXE7mWGV9C8qmfTZwCA7aZz74Dkv35pjTkvpkbRMddbKhCNI/Lnsz2w0F0WO9Y7cWo++0i
uAFcx8BwVJa80g7Nw0bQlqoWz72BSr+FvN4ipcYyUnx4e3w1dPw0FZOSYrHLFh8KMbhYjW6SC1bw
9dSKi/6LsL9iC7n2xul1sLHFawbdwqbhyYC54nHgDeKkwhGFfMkWNQY++qBxf6+hz78I0dfectxy
tDP4hP3P9xQ7EQW+AZRQWC9HGziLR7h5Cw0QavjnLNgEXF2xFcj2pdm+xn1Esn4eLK0wi0Lgixnw
f9W/ykekkWCJQG5if0WYASJZuRNDUhLT4xzWNeM3PisLg2kRWt4WzxWIxWueHE1l9HSP5g+jd47a
yeXkCV+UMnXvrEgJyc2/CIDkkT+lNfO9LuqHlrja+w+up/ylb70tQ3am/0NxkNrVrIow6i8XutKD
fRxpLH4f32CZ9dNogxXAWWs3B19+qC/kQ4rI8+JTRBVCBlLsjGBDo5mjP1eJNH2w9VIbZMufr9TT
p39jITwNm3mQZUPm5GsnXTIkZsdqXm76zBo9E4DbNwjH6P5UpfiCfEWqEUSOqkvzOnzZftsRJuRd
SOMeEK+zPm/EINttjgtoPq+cYZbHkmEUDc0tqdASQssT9J+9Enu1UPPbBYMRBskafYFZ404L/OZ3
juJdOu78swt0tDiTg5fUDCuPICNouytRW2LpedvP2erq/VL2Y544yvEcotOBeaHZK/V1CV+wfhAI
WZ0p8r1B/iaRc8FsMg77BcNeByFdPLFwfCNFr8TzI8SOyCeNr4Us/ZVwVeKdRBxtficy1pW6isaX
bKFP3796An69kkdWdPUWv8p6imoFz3o3BV8tCDhBaMkGMzQAN5Tg36W6/w99d/E059/6714m5j/y
uM8KSa0CK9DtfpQMkhU8ZmFI1cNX/GLQIq+saTRRfw+ioPwXTdUfITvtSnUhPqAwyuRdLdYiCCgj
hUSpB4knfJsYIFXnxKnFFeqzSAu7fpSf8v7RwRJ4j82zpuC+lQap9j7uzEOo4VS/eC1v7YBQdQOK
1Ktl4uiWPwFsK3pdt7uwWIjnWBC1zL9XypeFWrz0tYwT1x36T2BwXzKpCx1WqzGHVKb4d0I/Yly1
CPOuGy2exatHBOaWHmaFuiNTcS3krVYr/5AkbIu0WeVpTu/KhXr3knati418/F6wRkYzfIE8w6Mf
0UmBfrfMohQwjvNzmzld0Adb0SRG6wL4wBVIrPoxfdt3/yzVvt1mXmpaCistxglwd5Dmrg5oOsWV
Xe9QWwy+ZIuiYGu6YoDDeadM0JUuY354cQauV9f6aTga+E+RJy1j3iljY3chXtn2xYOkotVUQDJQ
ZiIadYTxl43dgq475Pl3x2rppdSQnYrXtIySfUOJhXTZDhupvNX4Tt8iAPLCHc5y5qQqRlNe4CHN
XRfpBONQ+avCJaTGbmgqmBbZeUv+I8ikOPrEhCBquG+GRTWcsCN/uh8A6DsrvpXBOAcD6suUBD7Y
0TqHqH4D4E+IY5aEv8w+5XzcUEXqtwtyPaPhCMi+KT75G0m3D1AZSXTho20CQRvgG9l0KfhoCB58
WUQ26xNcA2pym5tcBKJP0lpxxe8T5Utmm8efXxkSZFgxZZp48KBdTuQ7paiaeB9jYzptsZg+epca
oYOHLiFCXx4T30O2KHutZmovPGdOd1gz0fMRS74NZnt9FmtO94pi9jh1AcAzqrY/5uSF4LQtZ5ha
HFVpFF5Vtc4nqmrJ4gkWVPo+xpQ2kc/cAl+Wig2+9CP/lnAgeyNcRcDmOGyQQnIPI7Ln03o2djsN
uFvTxNBjB8o9K6IePVYQ0w33WhRiyCuVhge8sgAS9dMs2yW14sE4zG7zbZ5+tiRs/0xxSnZM6DM3
H/c/S7tfnDUOL+t3vUoi0QTvu+XtEqCz9HVflVbqG8MVbycTpl30skQWqA3Zv442NqLt/Hr/a03A
yqiEj9Od37jPEdGyqT30WYxlh9XG19hWzZR85tKpJDVUJk9otPf4Dfdk7DHgtnmdsiWzd0q5cmoM
EgUT64/UZrFyah35FkhJO6V+bC8rFXc07iMC0f0056FYwLdkE5VMZHuR6aSvmGVVAcnVl8FiufNS
kV9iu7miH4xCCKQsDaxil5B38y8Tj+YJk5pwktCA5vQhJP5+CiTj5+Vj8R1wZYVQ3TBhaZKUJ3vj
KVXwAxhLHrbQxGCZWLFNTe4vLcW0S5g/wbc6rBCVD4el5mPEDAaoO14YkwTT6/s4wQeIzlZockRR
dRgGM75osRnD/QtaOPlLF86CVWoYTJDxPy5S77V6Wzl+MEHBhcVYJxdXV4k9dCivAlEBY9WHysN0
AtxPgrgnV4hiXR/7c3l+Ri2ea7aSaTtZ1NueJ1HElxXwLDuTyraLW7EOuV+DDa8Xzf6jkZiI/93T
U9wZHl5326Rtgv4KmKPAyY6xwI507I45LTFUncGiX9GEdWLSblZXlyYwodxKJ9SytIS2b6+Kz6l+
jZM75t8QCeDZb69KlozYgQ8ctJKEemfRpn8eZHkrOhlLEwF8algwG3e3OmJgiIa7tHbF/i60Ys2p
dhKdnkZ31K8vP9SvZTsgepzi59c6/LbTvgOS71qol7hPJWTfZzcPTAaeeA50FjAuEWs/t+eIe6ae
Yo9bSZOfmU4dcKtORDqXQPwkiC51gn9tKZxCsube11ao+VNuVG6RNnWkzDFLItABnM9RWjqAurUq
54TI3qaTa9DW56RYs9eOI3yWLwBn3m+NnCt+5aM4zNP+TsQ4zYBwzV6WRMuw66N3Ep/99YtA+vyL
fYuhw6Pwkj8Uy1AZtRgTyfK53IyHM3QheVQVcxT1AfSgCL4gH/m4LFhuy+ypSdrDqSiGFedN6Rpm
Z3ZKAo+TIaxILKN70gQfvh75FhPmR3k2aNi/1xNTPHHkEn6VFqtQ0CS3UHPgxI7C7nDdU1ayU/rC
qCHtyov9YUKkKlg3PC/s9RYvjAKunawYmyudpr5+S4PO1WA33WY5avT1znx9/8hzrXa1HgKX34TU
29onPbsonxmKy8LkJVnuMvVEQxr2AvP8PmysurmS8diZsV5arxS1HrFDaTTM44tHgaWAjCe5u6e0
twQUh34ssjbmIy/KwTmaXdbkgN7+M9lEJtqHstE6sWdmo0wmzv/IgkiJDn0h1/L8UehjIYoHfjxj
IWtuVhv8ZgljEwdv2xcaIe3kXFFzvS46KG6s/XaP/U8RuKAHjSIzT/iQRE2QTAoOn2D2nYy6EoBn
vYxsky0X7jtEOVfZk8QTGqjqBoAKNSdQBryK4yPg/GOTeK4x9QoL0qUdhl8rVlDMisC5FzY3zcnb
qa1pnW1h4jkVgpeIiJsz588JKBlJkvHqWbUE1EhlTE0KLTHah8MnRwq5FbhWOD2dw1NL2L/3s58H
hJ6/NRxDCT0Av6miG2BkvNzhWJg3JPWQGujx2kf3ZVzPw8ixQ9Bc2P/BjCfyDQhFNze43p/BdQbq
EUEZPObdtSB7bz8VHfuLx0724NwXv4kfX2QaEOScs6rBaCXOuiCIoY48b8jhvPesopzK0F2SfrV3
QdRBQC4Li4B4EXRmpXFVqSc4zO85u50j/Q3rinKWboIQdmoRZ1anb/dn/0qvw0HrATOgdAK4N1xk
5CiGLZwCOZlKBB6zVQfebwN7rLMy1INReoz5TEIf/GPqYsCPgwgKhOYCU71VaUIU523uII+rtDv0
TrCSCiD4K614gOWWJGccp/yMwX1umInDyAQtXta65jxz3XHHLWXBboR6oYsnZA5yin5gVIIJW39h
hlZ+yODimBh/WmN+hV4Hz64L5D2jAg8QzILdmsbb2JMZNECd/0IetBVlX8gchdgh3AkneeTxwOXt
P0EKfwrcgNN8UGT24DO8L8dAIwhxcATjyoTo0LM8LqJA0An4akCUJ6MYPCeNjSUHkihRNo8M2imJ
jwNMtsVZXkq0KpK30nKf+DabYwDxyGlEByvjo+zIAVWpQWbbtTUXSTtcOCWRXHCX6FIzit3M1uSE
apNE77IE+1h1clfy+pI2ZnvAk3gVVAsMo/8hVsNsz2+Mm9Cd/jRKXRR5b3Rri1qhE/zTyuByOvXo
w8Bnn1Rp/v9+oSPqqJK3H5coiY465uk2V+kNfKpLDxGQs44IoT8VapPph7YxM7IIfva72axox9AQ
o/5t4vSfgDIO2UIanWVCVVLpUjZIPDK0eazJxgsPvjBAg5CiCizvj3FClWHge8wEuQ4ZUwp9qmWB
y0c4ECFuIq5LHafxp0kIoHGmKeWfYOCvmfCT41+KUP4MUQLL3hSdO+VPVA0pAKCM9Jn1m/A5iMgv
TbRmORqaLOSvEl9/gy+MFIXvsKxJ7VdUXIS9LvmfL1UawH1MCLHqicW8A2ZAz45Z24CSqDCTQ/DA
77vBJJOJDbshtLY0qIWEmo8pV5yBlTZW5bq7XXfZELWpty1SIHIjtTUokj9ElQSzaR7YeZQrsQVT
baW9H1cghvJFMU2Ioi5vsmltP/9mdBJbzlsiXjAHTCCFj1vZnXE+98xeAZDTgOHB8nqbAm1akQVl
sUBv4APeoGlL9TJMDrcc6r5sYkS6F77nJrGf2unqW0xH1/dG3I43n1YJUSRv5V/Ux7LvUIC7jo/Q
nleZy4fvACA5ifVynv7zfeJa/JZIl6L8zyhfoWC2PrnFZIh4sQNAAsos3BelLDbG1Uc0q2WMWs6l
lQVwZTyzaQQC3gAVN12JIKlk95YP+Ga9OcAQnXK0RTjbRAvy+9cUFDXyfr9x5C6yuv3JIp0yMAwT
y0v94B/dmbSuHdGuQsadksCkbuphguYUKD2yOOQT3+tmHaSOXFt7gCBneKrhStfl5JdNcusbtraS
aQqJrw5vMtKc7Hgabj6lwGhkonqlz9wzmYiK8wXtj0EvapS/5Dv1tSAmsg39vxctHRuLGL4JQjpD
r3hgKlcGWviLrZax4JD6uiotBDgwS8FduKRj9wGgDHM7EDpqFI19+15usYkHTfvp8EnZhutC09I6
T/PhGxsPghbNT1nFe856Q6tunvtfJQmQvkBIxrPbQj8FcqwQ90UC+7SnocfY+AtOzfrLx/cRPKTB
q8R96+kHSATOwvzvI+Rm3Xz+vkH9CmzRP2wl17rRjeLaHxXnWCNkY5ftnzgeqQXAaAYZZlg8+UGZ
0ix4K2RThAqdNLCmGNfAL2Bv4UsFmZm5Vqwf2JW6Ju8oFKigX8NYuzjExCip7eXQcSdnphtx8bwZ
S+F6RYVud2HFT9rPE4Gl2y44xHMTRs8wTRVgCL3IGDh0CR5cHkKFZT0qlTZfZRfvxyLwTAC6aarj
6j0dr09jBqllytxpqU0TZu0yFA8NwdmrPVc9LWQ/R9rgXjyY1cv3lBKQQe7Pa+mDn9NumoR3iVPF
zP2MOQ5+SiyvGNqeP2Xy5ElYsZ6GaHKLqIghNhjbz73bXFfdFWmrUhJiLgL2T+Dhn3O8/U1YUoOh
BmhoGeXqxOlj/+E4kTGrajBhVBAXBaqVeh7EVSn9i2f/ExrdaDzanYcGcWuHc8mpFFtjsY60rcdo
pJuXsD3YEzS3ZmsWgZhiTinQk4nKznvHPjm+znAXblVHysUmdDVcw26dhxqXfHOdfdm7EQVZVEPu
ilUuqzFK7DBswKLYXyovcaKU2K6yVEMvjJxzvCnpnDpNSE2c/SLjStWPXPMSIXAxN3WT0dQxbxo5
axpZvHQljDFTEcDsdMvYaIcGaOhP7BHz22ICVNHTNmY+Q9B8kAcya6WKAMEaN1LNNCY7RWok425V
EQEngInlZ30PIJQYBKV/e/b5t/mYpGs7QdVoQ3fnYMTogKRTpTWOQwYg70rFMoXMXLIZAQ+E+09J
Nav21d8O7rBAdHpg9tjEBkmleEqGpeaSiMDHridG1WJYQYI35P1BsybBMvtLAmGIM/c6H1iVDFYD
aJ0JkN+zR+UISLmwac5kTpq7wvouF9VE2InKifUhfXwDQ2hyLBankGOg7K1nJ+1lzXO6ByNVfd4q
1YfkL1srXyrzzdzMXfAr9qMjn0STYCz1YbFSmBb02pJ8CC1YUlf5AK2BjIA2lXdQbVFnodUYx0rl
H4a/kBFYPBlX7wIJe80HfdN8BghsXNvcctPUnU6QIeW9sOf3pQoO2ot1fLWqkeXE6O/J3+8Ki/Tz
P4VNAfmLe2eMQ8OYg3YQVooX4lwA6thLIcE66LH2OPK3xik1nYlyCMDP19LJzTYd827YlKB0MkOf
6jGG8VKQPxp1RSwM47n+EbM/DTNGVZ8D1nCSGYbwPsYU4ekx62VeWqlMNCbIxbPHSrvS8zjykgf0
lUsU4nCKGxbIM6Pc9GAns1HWQuYCmnKe/VV1FlgrhTt7FMn8VjnVL+VgaxT+J/0SxNVesClNUO7D
My9yZwl5yLlGPq7rQWAlS43lC9kZimugT1JN7TiFGqe2P9XZWIuiN4G3eioZqcLhsTKoLYMN/lPd
DjQvEFzYkh5ZZOgKuFUvN2uZOm33PzL4M5q+dcbMB0ebxHoXU/Lvw3uyX1NfO6merNbtovGWv6Ba
p3H1Qz7j9SgEksyaJPeADYEox9zPNtrswc+GVBBgJdNT7tzCl/bkuDZKilS8X7ykyqN+XubabjaQ
AC7j9+A62KixoOh+mAsA8E98UMokILlyo/aRrcrihCWiVjQnRNMBOolONtVZ23868u1V5MrqXURB
/2bOr+nys51FciDNmcUg+q5wvDxmc7C9OUfcsmXxFqspZ7gETCkhi3hD5ci6ODkgkyLWcq27iB/V
FlWvgFpFSp6wWuoeCBgmj0Adqq/FPpp+mlCAxLCRL+TQ4FA3HitQaG0HwUJQgCi9ot4O6dcWXMma
1rmIyzoMIG3mXX5l/o/cO/zsLtG0L+rJ5XwRnzOrxn9cNPPQo+UyPm9i3PSdeyLzfX+NEGzan28R
cB0Dgmk5VijHfckUiweo7kBT5nHUF1XG2FnG3OH7a5dJ4bQS/b8mkBQKfQi5jXS4BucYWzyLhmy8
ahFAW1Oy8hfR7lj4hBk9x4XoliBXxhfNyc0k66KC03w+0ozmSS1Aji/or12oHxMjqE3VThsNSwTD
MTz860w4Qns0jmJ4r790eUyNBeQd57f/OAPNbyMkZQTr/ZuYTQ6WTX59NEGMvr45S+K6bC1CP4RM
HEH7qNdksl30G5oI6JM44U7Gcg7LG8XaRkqAwWY/RFEbVbwje31t/ug7ytwNYjXO8J/n0nuEX1n7
imPdw+LR+b27qBlPD/n3oXdW0cIvW/41VnQg3b3zsiWd1VuvG/T2lCoaBLb+bMrPtYcbS2wmtX31
nPxECOS+w/LB+PYDFtz+NfNRV5ko6ICIzoIGg5lrzXu4XTY9B2HM6KlBLavPjKuB0XCT+Z3zOKQ4
FtblkXHj6PP7QicBkk8hcEMlWexHpvEPBx7ZmA4zFxmJ1FmljxbJTeexbOuqWiilWJJJwwkssUF3
CdSfWEJ+a8UR/wsRMApERvQGeiko86RUpMteso7NVdpt1ln+TE4yFI8D0mMZUoZ/D71afFn4vinL
Lcbexvseypx66U6T0HR2bUGnvwBZjPVz8gTBLlb4K4cwI/h4XGHK1Blsfn7YmicUZv1PcnyhLZWJ
nHAeRnniiEY8365MReFiWPkfw+unIEche4k43nIiquZfYXhUrKFAGUqHP8Mm788KUMRdj/v81Tbx
Kd/ZwE7Wmrse6vA+IY1TJXZWdozpg+z0iaP6rR7HCE7mUiXZFgLDoEAk+ed9pMon5vcSFE3pyTCi
BydbBblQWbob9fCKHfzkUcSfWpzhgSw5JTEH4a1YFUv8D9DbmWUjdd+g4pVLHxYDzfUhQgNzZCLG
4oQxlPEgBG6CfIU8k6UXJwDEm2SQ36aQ4sRWFbC0SfEridB83lvQJ5NpiYHJPU2U9pfMOC8J4sOb
/BKm3GmYCObHE+pHR5YDdPAB7n6EzZRBOMTMFMCG3oCPbOa5Eol+neyBPcE+qa+8VQkxrXUFj+9H
e00uNsyZ9P0w0RljgRHO62/AKVnFk2LZtdEP3I56hT2hYXn2iYwUyC/F3k6NermZBMu8wfZvHvLr
Nnnevz5FKeT1QWu9sJFmOySxz116mhLnPGhtMaUXuscVYQjRNXo/0r4szqOR8stFEJRHSyfeWYi9
3D9i/cUkiK8Vx6ND0F/0Qf1gXmDv0emrqCW4m28kG90Dbh9JAoSNkAIRFsIFj9CJjC6oqw1b0Gfv
Eum/m4MLmlvovpvxjUOzUqc2NGZxQvbCF51np2hh+GptUJehcV0k1WOWJ5FgKYlMUiWa8Zl0CkFZ
d2EAV8kSj9BwMFbEa/D9YaF4yEtY+2zSXpkJtfrIS5lKwdO6tHSOm76vuP4wauMvaSwiwcd88VGX
/usgGKn17ZN8ekZo1baf9q5QwhG3lhrmdtKSsScjpkpYHQN/jS7P20j8bFERcP4Konmi4gRmmOzu
Lhmg3cECOKaHhTdDh+VHVRAzG2z0Jnrf6wdGEUzo/1jPTFYVQCucJ1MHWLTfrm//J1QcXOa+H0NV
Y9sNufxPcOeYbzy0kt59WgyUr+b1YYZzBo/R10IZ8ayCG1cHRCqnyqd/xo1U+Wi8kY6IC1HXMFCB
TbyjWtL8nlogN2TgiB1Y7/M/t2O3jwxjgXg4QULEpu9Ze9jHYoPTF4blDNaCpvaeOG6VvHASTXKZ
3eyXj3Mt5/XiFyn6TAmpRPQQ92sBawTgBGnEyeTXDZzinDVcdIDa7ue+iugVrjSBTY8wPnyfczxv
5kMf7mlPDZXhL9QfHAIJHl/ibPsuuHz0eIGeySg+6tbDqI0B0g7nzuI/GP7cLCDPcXz88DTbVt8W
jRnducoqofvHm2qawoHh/5n4A64BvRkEvamJO01HtaXH5Qcrl8ZIbXXmYIkGgi9RagWkHn1MHv1U
Xh08kKAOA9DUCCoIJMj3puYsDBNhUdJ3v3faw1IQfxYBgrF40X5LM2hZF6FNt6aQ8Tiuo2lOaIzi
DOx6KdMPRE5fLXLlf/lUrqoyYaowx0lausT5FWyUQilQw+ZG+MhCbBVCdX+W8GXu56sRhIgVJr/l
7kphazUTVA4hfNntCFFl5L8aA3SNcHpSzpveYL+2PxaMxhBi+xO3LC67LgGCu4pShA8AB1qan5qE
b1A/cbhlHETE/o9t9p9uSAAdqsB8GuCLZEvfUMZoh6muiD3UUBYT1FV+wwqLNWtYVffKfQHnJgXG
9sR4Pt0qsF7ibln+JHidMN/ng77v4F+59CU9lS+hxn38WVK7kvDiy9fYoqlyMf3PRO4K8Hmoa+mF
JXNmAB7wrlWf44C10t5XAxP7q6uKSnJ1l5twZmywn0Ps+579fEBumjSVOt0e6SDnIfuZNKk6456R
YDern4rjStt9k/JzPQn+s7uc7QERLyLIlzsUjBqPUY1SgK92uCeCcjRPK5UQ4uSaa3zf2xN/oDg9
sPHIagFW6BlrFUuAOerjFfkgYUw+qnSIhZqydGU1cM3nwHZVwCi5gynzs0py4IP3tGDGVGFi2Acc
1cYIXI/BMCWm+O8PffuwTn6CICgkT1uuJ6rcf2a5nlGGetlVsi4or8N7gpr4mx2Xt4Z1bmCcGQdp
3Q508J+WhbRdwU4WGLrijWD/ImL79A+jo7HLBVW7P54z2WLoD0/89pv1oGLLlHtBW8PSEsC8BMx3
sxnwhK88L1QhJSr/wM7cf4KQT0x9pZoUCU2RZsCskEpZbQOere+pNkW34IcD7RgE1rmZAY5+mRmd
ylRvQa+5o9PLB5s6DX69pR1zpgAAfFHSLNjfKy6YggKZlyUQCdG89KJAr7W7Zi34IZ4OW0fn3XOD
nRWiJ1DybQM8S+rbP0/ZVvMxYKMTEBjYo5TwcPjdTcPR6+XKqLxcqQEZPuU160hKGRSQ1oPTfd4v
lcM24K+83eIhWB+Yl8POKP+IOJ+GG73KhQYIWDCDpeISYnLelWcQUOmn27DOle5LxXv9IbFSNf/F
VW6MKb/A9Kwvhz6Vy0A6LiLQGLdfyowL/VZBZw2HefejIjxypdu1Z3TN9RTW4CQF78bmENa8fXF3
aPNDxyroDFWTwzpkDy7vg0ubi8s/2at1ust6mMUhqUpa9O0FAwACCCfdbp1wuxFwsFDOlRo43SNu
vlYfggu6xzpe3mN1nxkWi54BtamJNg4ZYqJIm6D658y/LYvikAa9vJaS/kSyw2/N2VV0U8Eidjdp
cL54UX7HhVB80k4APPzAqHgIWoLZeDO6gKVz+AbQs7SKLOGdkQiZu8kiMuYwbziy5ddak4fGwXN/
M0Fody8OrR2SX7P8rix0FYWtSyi0pMjoOmgcCN74WEO3s+K36bmGpSfnYBnU2C5ZxW7pHTKgPxxO
kscL7698T9MPeBQ9czl8fb/vVWPWbp4PcM5ezhVmgwI8Ebo8HwfCjenNSJDpg5cQw0PLCVgFKG6m
arnbm4eGR9K0kut2nW1edwjkkYQxO6zy8UhPfi7YEwuf5xyUdM77ySwhW9Sy9Ms+6sIvgREE/yvX
3K5UaWgLfd9AbBYmSmqbR7LVIKkp1IB0l+xw3r5KFpUx/+MpYo56FfptIkhn1lQ7QCeNs+fzc0eF
e7sy3y6tEvziTg/THE/CGR66Gudqwumc4DKPuBmH4bhKmKbFfB1nW7Ffx6ktut3BgWtXZM7HDBt6
FhQ3nq7drssQ0c3oeO6o7DHfwdGnszDdOWdFLSADtGVXBtPhgifWux4JzNHTN98kKczBh9XioDyL
eqF7yzwJh4B1wGIWe0vidyEImwKE0bzmF9jgTtOYKlGRCqZwrNumDT7ExAw/72m9yRUXG1WGXJ6u
QKPfwS3TkWHvJGSodhrSMr4+9oLVFazzVkHFMpHp1krpSaumPwB8j3LHzhr78bgRtFatcOLuUV3g
+7stCCDXtlpaC371tbKop3bGgorR4oBsmbAaUwaJq5rb+UlNN+1Zgi/k0OIc3lIMJ/2jvMfu8ND7
3SXmKd3mnlpRZoM1pHUjxduJ1u9bXPnWPjyGoiOTOu8KDBpzTwpjOx3RpgOu1R8PUcA1bTBLDQ0W
rNvwukwUv6HFH4NcHqwYb8J8+FTSyUWJyvKMspAkm08+xXNs0capMf0zr1sQ1MovTn8sn4Kk/csC
o/opd/vLAmPTwPwmgyMXeer3wShM//PM6QPYa9s05BOkr01Q4P5jhtC3YkYEO7ZcOLum2Jq1IHFk
HpFx1+I5gm2YCYsZMUcWRMBSn8nWRwwAqtcgoaiAlPPYKAXaYGZnw+JD6dj9VJY9fzbPlRtIxyQ8
TjQq4OUzEqF45eiUInBJTMatdvmdhV1ZTpsN9YSHhO9gUgZw9vovCKu521FUb1uLtIJEYzkC6dNN
dHrJdQmIecLQhPGGO5ofcOJ73+SBA5cDCB34g6zhqVHzR6lsBZzegtIE4jaZ1Zx0Vqq6S/4/+WaF
zpb2UVeSKRobCQAWj3fI+mvVi2Rd1rL8JlcsKUfXvfh/pJVnYNnD0fBB9/s4oYS70G5bHR+lr37q
oBVbUi0S24dw+U9t9o1eJq7G/ZTSn62rQECKzSVbvQr6+Yrnt3LPr2nitRj9zMIh1g7IZfP/MxhZ
OZ8fe8Dzb441WOXiVYaZAlCZKaQUEf9+srH0TADhg+6FbOFGy6irlExZCsVnqBFN4oUX+UmSnFS1
25f3cFw//NaQexSAY8aTg5OkzOB4NJrh2N8hypZdDh2aJfUkYouLqhvog9fZPflkzW2OnaDdqZnD
8YS1nZiKB5R4o2/vjDmSLKWbVeSluLvLTwwzz3Rvddnwrm0Ee2JGgkMRsEZHYkSOwu4MZVplbBDE
vJWQkfDlocMcqmTN4d7ZElIaeQCsvIpu2CBgTnnb1G2Jx88KBH7/tjZPktnVVquCJZoxwTF5ZlYv
A5jiaje/7rFv01A/7yPnv3OlqX1k9Q163lTWtObeix8xywHbA97J7rRa6lSCvrKsrc1LIlvExXVS
8dyd1+B+1GN5Py1S8zNbkMwn42GS15a39lNKMcY2CsBukXxkH4JD2qQ0ATiJrY4gZT57NFT+r5Hl
gSsEFGWeXHlAEMr/RzSxqq2/LfVnUEQDR3zyv5sH9YNCU55ebynestfIO/+V3D4WVTHNWY3mARbT
rFmSWs2r9osFcl7L4OVQOpqtqWTeenWWko1Z1znYde7SZR8gqDedrqqxRsPLQGGOChxeNfK3QsVG
fdGpk83wHglXRoTHrpGZjoRLUFfUphgHYKsIYLvMZ7V+M+OzPpFfpVrBvOBrXtP3IEGUjNu/Rssn
rJeUSyBuIlxY/1jbDsIpYVSqLcgBxqSgiucNDgKnta/8kGieTxqyoC8j4pHswV5Gib07rvTW/BRh
XAjI+SoPSjTeAijvkvI8SHan3Y8Y9RFB0YLe25ISJpOHgqkWc4cY04QqZkxqf10E0PtEkjBDusiy
cBEYfSDDE878gNdOuwXhxjCkFblhM6N22GkR4caTbfk7FHAjJJhWa/5mTS7aPbH4r8SQoKdxqE7O
W/yExCACL0H3wpavQCHsT2pXY5C3FyX4WRIfanLxHujjvpaZlo33oaTdPLjog4cjpd+3cPDLwT+b
DY0hgljqKGRXtoXTnZYx1Ce0L97MByalX+qNnivhhXhF8OgUUMp3l0J79m3XSIKHzEcRn+oLEHOB
Y8/HwhvgJzGDJmKIcOVBeX9yREtGQ9/bB7MXYQ3im9RBNOPpjY+6boiARZnTBuwNFmGTDYCWUmrs
hb7bmKNq7Q4NPjA7sHdO7QO40/PiqI96rxfslkpj7iH8VWd7Lm8JT1xEJh9cWoQWGgwnXnozSNXT
Pw6hM/RLLgZzPk9b6UMOBu0DD/mvWXktII7Yzkkn/Hpz0U7eE/xeg85eS1QZh1ZNQZyk07HgacAa
7VCPy77N1hreK+84AAWI6UtXUDVThtUvyUrPObNi8fEPa5fAKuR87Q1i+9wGtd0rie5rapcaLHu7
i6vfa7K8fq4YHloswQjH69Rsm6Z6ILvsL3gKpn7t/ev3W1jert1F2nkBAUXwoQPmiRI97A3wxGmn
wRyRp8hMZj+S5uu2gEZ0TabuoB4Y+g1VAJVL0M6xUydzVTLj0ELQE2tvX/8AVQmZXNLZVso7XFD1
WG7hw2qFH8+SMAz3ClCrZdBCwnxM3AvlbkbACaex1zHIFDcQQY3knO4JiSIsEyAnxe3CCSTXG4N3
fq0dRpM64TVJ4dkZeRjsFxKV1LEZrU5cAPFkvoIV7QsR3AYZqoguOLadn/DC4LTpF6aRrz2Ay+yA
8xG6yERMzb2PFMZm1mQl9uPxX4aaStOt7h0YcROV7gCoH3OlYDdx4PiR4BflELKGsbzRVz5wGSNK
NG8xEdfbEZt35bCVigegEm3m8YtAs2RK8HBPxhrIJ4at86MykdRWKZljHfsGRdMIeH4J+lCKpjBg
ffYjTFQuoYJjTNmrTI7SKY3wtuZ211P2wmKj+pU+eVepkukZIE5k+OOAfa+sOsX9+Nay81rhboG1
zrjjbdW0aog327FQEmtPANxIpl2nFxnwZ2/WOsBxBfVz6l4ajDOw/bHM8P57O53FrcRr23DQmDoM
0iEZ/i7Dls495yyHAkib/FOTeta1SQjDICNsWAwmX84kWAGfK+hundFwZkofiglLc/4Jx+14qxVE
KabG+Fj7pV8mQZb+7jQcpb3rd5lUTIHtMUgafKuBznBMOLQGvTdtPk++A5xeftj18ooRpU76gtSa
mG/OFV1ho/f8N+K14DxNkI9xaaUJ0+KoSzx7B7GnFUtE49T2rLjGjBtDAgXujV13BO0ZFAvo8YsI
ty2w7kDJlacLDz+rrVcHuqcUSxYfXhHfXSEXYbgtPFP7uYrSbf5EWPUrZkGZgv2wlugtk5j6V1Nf
VnaeEr3yFz0aTa/oo7QoNVwE9y1NU3AUwHAsIQxrwZhA30JQ7enmaBmwYPHwb/PX6aGaCCQ61l/d
NRY6cq8cxfG0fQcFgXhOcRtbdnOyqbvpu43tL8n+T473UOI8sK9T1p7FICB1ZFbEGdr4nviRByk9
0VjtzKx14DiXQHhlXQIpIYXWq4lfzyUeq2675ua8myp+DFYzh84g1NxAUzsddmjAwtM/df5ySWq7
Su5nM2FFnCYYTEEiERqp4pDsv7FtZu6VHpYf3shzuS6gIgYYIS+hODFJmjReIbUzsyGEF5X3uNYu
eUCmMGfuP3OljkT2MKLMX4ZL9UcZPJTyJulvbY5LOUkmf5fJv2KgqdSMYae5krCQp4xRg+h5+39Q
OUvX4KUK37AIycrMr5OmXev2P8IlcSpnZNfe8aOcdOEBCRN5f2XK0+zuoWxURqot5T6ksfaplDKZ
/xtrcpmN8jYoGv06AeSsAeWc5q0W+ZrdQUMySJzDANiiOxGetFCSEQ5XWJrrLZXdklypZ/YDavOk
LNZNWSa4QLfJ4hzqijeHsHPNX8Jj2B5Ot3QtdBZIIdoTVYLHs9RbWn7Up1n8Ej4gZacvawnV9jAa
AlGRbrcE65tTbX1wLGn/OcSJr7AbvZbdFQhSN7SDDBREELK582ZEsPdtqDZ5ut7cZiL9dfrFZD2M
0fEIOpl1CsakymOu/HVa1rJxnDkGifUlhfLtIJZSC2WOhKdPzgoNnRQDM4XCZJ5mYAHGcGzI3Y06
MxA1bhnxVEcyK+zSPJVqF4WAslU894daElze2tpedyPaflyC3zQrO07jXH9UyYMQL5hccqqYT1lj
SEd8YeBnweg0toF6DBjlKYxNfDnyKS2I66IlFuV/h2JIFn8yZ1s7czpqlQcB9KoQ7aZjnpiLigFP
mPm68LwRkNCGtvrcMc42Uira4Q+4VdfZ1JJR0eDBylrpp3QO3gAvKujxvpmpng7jRYgwybQhgC/4
mS+j4hgflHMNbVoJjAhJpvSpXjBKgzfrt0ANa08Vlme24qFy1AGKGtYJmk9JaSmmWxuA9+xbUzii
cQOKTMRxIy+VYVBlMa8TVYoJ6mYMQQJTRyhTDR/Vg6gY5htMwEXHFfEG31B3bcL4WTCGbMJbov/A
S8Im25n+5AEkd0Zv1TAcYswt29kSxCXI7xY3mg17EMkhWYvvbkZGYChFWmk3rXxtwyss7ZEA1MCV
wpmdkT3HhEjwKqG6Cls8kv7wbhV1WzG+n9CTKKhQqsQqG1LaNikV71n48ejLY4zNrD1D9DuskHN+
EgVIzB+9oO8Tpum8mLBnSm4/2dNa8HWE1eHbXkDcoDuOfPa6A720z18EMtreHjS8md2IUK+gf9j7
w004nIUOL5PMkqKUkUZLUQT3WnWxdfAIaH6fIm6rf+KHMhJqnXrDTcqC5e4g7GgZWneiHHniB6Kf
60/ffWNLADAWtc9bDMB88XhPG1Ne5SAwRGihIlj87G9okrQbX4iFUbDPxNjPlQva00ejzq2hqjB5
6zORMrn55ilTAVZTnGhcJVm3+G21QvSVDyOXrrZYelr0RFLWmQR6PGMdjxsRBeIteRg5m3jhuLhO
LUxEZWNMvfN5LoCiSeDwVY5X6huY4vDCYv+N273X1Kp6kJ9IxbBa7U6FucpEj9lb6ODoM/5xYXCQ
+nWPeZR5yo+L7ctc6ridncABxLkmf+RoJAxNUMgX8bsz2vyTXh+lFuxlSIRR1gNGGAjm6LIxo74l
7gLvS/9SM9lotSMaSX479E08pMeVJbtNDavwkOdjP3/l4t7FAJa+hG35NAcP1lugfQbSrfMfflc8
TnD88gwi+baeC7hkIRsRBWaZj6Q+TR0snyOHB6jIOpBHcn5Pc4Zv3rAeORQMy6ebwPvw+lKrGvIi
eyN2qCEAIm/zL3/dwmUB0BYDg8G4oKwXU/K9tGf938ncngqEgVlQ3mFUS2u+hkiOaAsrBj0mL5+/
3m2qCA1kJHyFbOvorT9o0qQk9wsBoJ2RoVHYwzGoXzUW8kCE5nzvbaBqgUfb2ediVm8BVFAielaC
bVLAhlsrE5WibPVXh2nqCGj3IL7Lq8NVSKPems+DUuvuO60h6Nc7Y4SV+I6bHnDtOyZXc2OPMEry
qWter/P/lRBtggFDf4seqhCMPsN6m4S36WNU7iogY+7mG50rvhknHQ1cB5OM+iwdi+gU/3OkJjY6
xuCSiBrv9boNHcDdZafo10sOtvP1m/Qf8utYrd7+pK1id2TNkrWe/NhgQ+nrEl/1+i1Nl3sDXr3l
bf3C64G3DtDVUKwLx4COeLa47qfEfwgThuHNiHP2jWoKHX574sNOUneUN8O4KxARcBpl2MjM3iG/
pF6SvBLfjx7RfEeY1ijdj/u+8lPHJhuYXKgB2LOK5d+n87XqYvWiLtgondhEJf5SQn7QfWxE2eJZ
mBzP+RFqC8y9HiJHeXIPgMdqcte1YG5yWGwLE+x4dTLLviO9gLMJOdO4nKW8WH8/O9PRhMGx6quQ
8ISOh+wFQYuE1ARwpkMSEtOYstxDYAjiyHc6iRFrtvKCo2AAb9pl0rQ+eyfsBrcrLLji2H99qx4P
SdTIA+++o3oV6x7tpkaged0rI3xCevvNrJr5MPb1XKLt4i/wVVYW/G69CkI/RvTKXbTlSDiRY+tk
WBXiRz5++ebKcnxVV0bTnVRoNHwy4dZZQmKYsutuiqLEbERlkxniKBqaD0sn1T+Y1J4AL81U56GX
3qD5Y/GWYfzTYWb3Rh1g5/Z9mU1LPxycIe42KhhvsNfkJq57yPNhIbS4i82snTLv7Z5kqvk5Lil0
5xZpsqY5v+7tG/E+1Sb7ruKRIP+QAcDTLMI8jl3MiNoSEy1xImEZgjdQgB/+CF/SUljKFgB/OH8y
dCPx7F2XfrQn4xLFULN6bOV5pSszTWahZucJ+QXHrGM6CZU5xt1UpmJBZRObESc5gswk1IMJKL9g
j8KcM5kFPcKmSjPwu4135//WmnCc2QK4blzLFv8xZdu7pN/rKBSRVW29savylIGwvUJT2hWB5n8z
ZDvFQgp9nWPUrc0z69RAZ6oK2uZ5e0YgccKyoE0eZoGaPFAFyg600Us6Zf/IyDGc7xLNoT+3dLV3
ggD69kcfep5/LaeLVO8BxF9IaEiz4V+tHsZ4q44iFaZKjoUxhMKheoDiL50tSo8QxxmdhLx63ird
YcYkS1LiZWDzjzzStchj6MtsoNaW0JmrrlUtyr+XI6ukGEfILKxi7axnvpYit2LEDCXPOIf4675E
pRxOTa31Tnd0/b/rcg/VvWi+RgrJ7TrSxILi64i9LN/XXQ7vs528AQC2sFrYWuDuG1Iol4yMfSBo
/x2wUvHkMCvxmtqCI10NdMLM1OUQJtZIXXK90i+4ztgT/ZGcfqR1SaVoox9S6YHAaeglC2Z1mns+
xMF+9qfMW6UK3QmM3vhGbfv9IZwEiVeWNjDK8xbtVaOIEH35zOzUqAWnZhLoHLXiQC3fTWimCoIp
3BuZ3xLAkCfUUlxe3+c1hd9WmviQF1Dfg2u7ADbeYHIRn4M5Iu2hQ7URm99E7KH0dj6DSqAedyxb
pdvA3WF3a/pQxH5lIsd2uiIiIsvUmq6nl/bnpuXo3JHcql7SXdT+tCMxwm5ThmjSLm0/mFzmWwpZ
cZKnV0FVj1IiG4MfSMkaMkTE8friO3/OuuyQfpApKYM3z/RiTp6buwxpX5QxKjOOJalhTnvF8tbA
i6GCpvd6FfObeA3+4DvGgNZmgKbiLfrBR7vci4ihtXhyNYIg06JiVh8o4A/kV/noHCLD/lufyZag
2/oaOfxaCMqThkkKYfpevcRbLndvAc53JhlanwK7ghKr8V3ONimrFaJQzDjxFX3LyDn+w023yKZi
p3XqREDtANg3uA4ZAXK7+wnExJwRyzJfBygtqhbd4Xo1sfgTY855ldBRrwT+XvjTiT4eIu1eEZu/
ztKguhLAldXzRvBnH0DTIQYFBxpsepC9IpfgoqAuGW1rlIHmZv3XLEDTkFnIMbT8Hs1GKuy65NQN
qLiNpGGMDdEhsfwjNPClN/LRCrxhzFuV+vxZpAbMM+M36VJYL2SZ7jKJrWRpVpymxzKvV734au9S
ZbXQd4hthH5uRFKLK40veddw0xIMmRBWe1ZDOJkDaAkSitFixi8VR0rMzPCwJ/My/hqBssaP39Jn
MVRNesJimvfJqwZg8wl5D5oL1p4h4/8lTE+yGUIBf9T7UNEjMVMDUBcVKMPv6Tdogk52Zk4JSEBt
5Cl85lWpDe5zOcECv4k5JqWTMD+tr0p6U78uG+k0SeRQmORvyI9p1Vhme+AXjNGYxakwhaVg1aEq
RaXpdMZufpUir50h4+klZj30TJ4Leut+E4X6XvynNO78iQsTeUJdjzFVXztzCZR9zq9wOYixt7SJ
RMiYX+AnOppEfdOCE0aVN1SWIzfb56x89zGRirhhDs/OMRBaM5vP/cECKqDar4806/QxZMhoyFvo
bZJY/GJRtzpAiAQEVbQBR8iCjK7HVImz1P2QchjORiGvn0tFUE0DmXYuW4brrvHywdi+ENikgJ7y
8BS1xs+rbMBGjfFhK/DHSz9gZBO20M4yO6Q386iXpMWYFaJc7MGPqZvIgtnvlbs57EX8tDEopinE
z2aPSsg+Q8Zxh2u4M2MRXSli1qzdsoBCWmyoSwh1bcQKj1ausMBymg/7zEO3S+AeGLzL4V7nZaUg
7KGL5Q1AMtkQc4PnVWtpn9u+E4yZNw55eWHpkXhY55eqZdCkgUiWAn0NG4qiY+Xa39oIn/tfkjbt
wyFOYmJ5IUgrP06kx3NpgIi76kmos+8oE1k7tTOuBhgYjYIGPw3cGOeCGohiGiRtvqSCMqOV351c
L1MiErs+EZkA7ZuziwvkwbbveaeA6CUOX6NxPJUXQCO+BqWo+xN7YH8bztfhfdyDCZWakZfRDFen
blHiHdqizEf658A9lE6hi2TDz+x4bDqwcG/1DD9fj+Hwyr07eW+0JYJeRMwldQKAEulX3ie/suKU
OUDimJ/A7V5l3EuiVSLynrsQB+x40c0QmbKLSp+uwJ7qalEqcX85oy3hRQFMkZEMjQjrJnVxREuM
af6xNf4kyRfMH+Gv88M13JXBRqIrNJrYIMbEYbjrj1F5elaK3HkE6Vn7GnArHaMwIY+AAp2E4zVW
JzerA3e0QaGn403MlgDqvibPszSGBP5WLmcIEM7P1dkd9/FUDTn32hYj4P9kpefH+6PNw1qwOFmB
Qj0BZEdV6pDwAsq3eTqUvfQIJYe18uPGoEkIeFcMXa5hgjOsGr5QGNgsDRZfK5SCy2AZajX+3eP6
sLzSrWl58OnV9Wn7aVUQkhltt0QhbXOxo9q+1BYfaYU+nDirIByOe6Y/k/hCNcVaVjfh7RKvn2pa
qpzO1h7oJUPDg3fTYmisZeWEjzA4vvyUo1IUffhjZIAHJFxejiOmP4dreuFCavfKYVmqPDAfB0up
lbcZ3DzOVMAiBPrniepEo8Fu3r/veGsH19xD/YmfYcY8Hrr07h9WxV3tUG5Zqn863kIFZNnkUgxI
99qPZT41IB2BYkmkw+jXDr6n7bIntFmnNEBceH+S+ywXVaDeVOuBpLXk5yZv6rRya6BxrcQcjgqO
HboMSKrbhRW6d1icDl5lT/VmxwJiQGX3kgzkiRve4cRjPLnP00hV6fzII71b5XIXzMBFq/BTSDMu
NDqJP+JFuQte1wMKPayLwUyXnTob4gTFYUIr8ESUTGza8CxrlOBGnCSB5nE9fE8k0GDxosluQ6Lj
4PF1wKDgTHCFDoY+OtLA2IQM0+sOoYXjICsW9Z72FokUorn9j5gL/DzNzqo29ZACNn8vUj2Zaj8Z
vmipwSfoRhKmnTbXKtRt3Lg1IzluY83jzqTQj8stLt1Ac+B8v9dcpqQyfc8l2HUsdlR98b6T8A/g
VBh1VeNpECTdI8X7khc8+d/2gkUC5d2hEsYJq88o3OpXYagDlgUxB4O/75hGTdxVUkzXDhz1Oh7D
oc5jfKp7GrWp0h66coB8l8dLqGlhevbmkrOYAjxumoS1MDR33FFZQt9ShMqH68OZI/wz4kgfnTSb
LFzgiBlO0BTjbbd7POoegXO5zUvo7HFbYU1VSoWu979RbtqVVWDYuFLaWQe+c0yhclu6uxEQkwzZ
P+TjTiOJIqoIk1Tb6dpt3vMhqD3liIcZrlmN0BNGu5///yuCyZf4vKKjInKZ0PeLXoHITh71h+H/
vBtdYmFDmDv4WOtMjZ6l/5SWES8UCUDCDIIUO91QoNNYO08uOf+wZJr6teQCBWOr0HeMLWMBJEwp
tmPLmHviBHU9MlcanZDtod7/r/amyrO3oBOR1hCEtcL9B5NB4leUt4XPZavPfXXS7JlZglpvXRLp
R8tNQKBRdjxRzDBqEDMI6LZYSU//RZtSPm1q4XbqwfuXe8oEDqiL/8ZKKCmE5lSy0WZ9enzSwCzu
BVg5/7tgVRKG/VqJcEwnRUROpyu3cxAdS7VZ1GzzIBobD+63/PFZ7oWTavp8Z694B3dzkJt69i0q
Og/zthk2OXgX2GinxNmpcm504coZ9gU1sSbizQBCVNkXvi3w98kKt+3MopiPhSYkAzy0tFNOJ/KD
8QL4Jr37UYTHiEWGJ0MX2CBIiwx46TmJSLOenN0zr+Nu+qKww/GQtfIAQLIbjK32bvFhIsMuvO8/
XjqfzV+l8tD5Lnr3JXlE8bk6u0Y+CYJOX1/wiIwd9huJjNLOHwtoP54nJU6EGxZn8oTzLLJmhbBj
2P4oyJO6bN7F111RVm58ZoGoYV9+1ID9QERbehZJVM9xZkmQ1n3QjJDZqB+EDwp4rebRhye+i+DP
hZ6WmGkAmMyv/Twh1+CXp4gJvGNzVHGjhgrmXr01x2wvulfFL0i3c1Z6as7wo976pPob/jwt9gPD
0dTIndcYKLg/ZenNYNHHoAitSKSjNbG6sKISulXOZuDZj2S/9oeA58F/GkL+Gumb8JCQJE2B0ICN
SsLBuzUVq5ZRx+QWL+ZOCQd7Oac6TxzNHncgs3rv6yJ2vjqWXR1NctHYGY2iRq9Va106lz+XjKD9
EaB/1PLGxEgdAP72CnQXbrhINRCq7Y8Qw4zHFkXpVjInsFfBB1QC1wM2O5WzEl6hfVOkkiKbo9k/
SIqWwUjfy7pnDWnofnBOZMdV0Oul7Did8wbCj1Qs3a3eGhAdMcZojoYb1CsxIaQViMhpH+OtBvTj
GTgt19weLBjbx4hizTZaoXdC+lb8jIm8Ufxi6PaIsQqkFdQM1XHrPuQDkKz+w3ShCImc6m8Zajot
HQxkQ8TSf0vHKXKyJkafd7jNwwOuW6Ssp/YlOw4te4o0R3CYmPY5+4Jzo3/5BnV0ORrLZM8hcyL7
VGbWQ5y21PARGos1y3HcKzd+/OSWHW6m2lYC3X9B7oVFyQRAjiHc8rMr8jn1BEYkCQb9CR1tlls7
WJGu1S7vBm4AZPIZxP0oVL8qXuHUv08bRTQGUR5zzhMlJp2L8nJi9JlvFa1wHJCcY0VohF/fA/di
0H6trAKsetHaexA6QzjaSbYIysv1meYSgI5nBjuIOh2Ox/myIsl2UAhViST6fuc0mFfbJmcnSfrW
CBWcQZk6k6LF2sc5pG7O7Zu0yp9osyMkQoIzDpLqYxe7GbJr3yrua14/izFlq7DBNXI3cgaXp3AY
CIfkvQW0stCIn/k4npGf0mRpiSkhY56riFKPIl4eTVcdngN80q1SajduEGDt7m4E+rGunyghuhjy
jSqk/h09XE9NHoMmiopSnojuFbWatpmtv/CBK24WdEJ5Sl+SxubjHZEvd6ZFfcsLH5wzlWUH3zmf
nS6wp1R6posioFbbdcivb0ky8vpVW/7i/6juynWdbj/3nMOANGM2IsAlNt8dAyLYXc2kP4D91S3b
DvaZOHPsUG21x3tgpxMqOYOdHio3ognqDxzWo5BagGTlugwME4QNqac18rcfyti1FjIr8WIWav+S
4k3cTFoCJ4kg8KgW80Yvo43tvKgn3hkHFWE9BJd31OTdA5a2mat0d2AaLmKGqCXysyqb6N25uEXg
cK+Is9Mo9VULNPqpsveUxDgBbly51P5MBrHSTzyG1pHx9neDl85gRZOyPgPVVm/j085hBMAw4u4+
vG9dRjkc90kIGe2h9AmnBaz+Ow8pVBfUHzVpr5RwzC29zVQVGCeW79Nw3XS65YbDtvaQaKtpP8T6
rwLfxe4SUUytaaQmYD0IMySaaoYF3t3KdoB58uneBG0tyzSYaEH8ZgteVDdFE9RK+GRGd9KFEnhm
qbs84GFJCg4viFLfJPKSNwuhhPpeU2BkwnkdiH7rdF5vPwE+JjIlxoFBEoyGaJknhztfxh/bdx2h
5BL5iw/CWkdw9vpXv7APhC77GC6wzl7Hl2YdTzZBAZxuh3RP2zjSJID4T6SCHCl00E8tEA8wjQeV
zFoYCYw/k9C/9qRDia5Dsm4EpqlmAPTakKFjSVWBSJ3ZvSAXsT2h7WhJjLRDNUG7SrLhDkWvDc7/
JgXU06RSck5nVvNHAFMeqyoBRsDLnDWIz6FItwPbw58MH8k+T1KF5C4YmogUavKFcu5kZO9bJjVC
TptA73FxjHTVLWMKnAJkGjD+xLGTXM/PN1VxQ7Kg1ZKSBWtW4GYNopz4zKbnfzkGw6w71k3RS40E
7m1nTa3c1101SejFU4UMw7Xv/OTZs8jWS/ng9hyngAK3XQ/vxejb+xp2hlVQixdY9WlNlZZy48Rk
mwSPP6t0zve/XzOfJ/ZqMR1UHkTNdJ1BCVbiQll3CxMuhKybMcE5FNzkz3aS4xXYYyiPUGZcEX4M
qzSx2mZzAA0S8V9bhSWHgVsFyYQ2q34V6hRO9hx9VSAJcTF96gwjlIB73WpTw0aPSJNS0KTJE0tA
mkWK3bF47OAddvmn6qsbvHE7k6SPMwXruVDxOKNJhe8Kqwa7GT2T+rP0qTmY0N9T3VnJU359+QBA
EV8KEiYbnuwoyaoQmUKNUx9woDqEE1kht8VC1kwL4/whDijoNqzV1v7JPbzXmluAIHoufa7N5ehD
GYUPIMFXQ56RXIyKKmDnxqn9j3j5BQBl5/Ir57tfM8xgHaSEC3BNlMtzZ3mlFBPQVtPC8SPOJjJH
Sjn7TiaS4N9l4QfMfjAFru26eD9Ft2ynQDlaJgVPPs4x3pNqD7wI+s6aQ9wAckBEzZAoxNOaBQPB
/jFmyI9FGpSUkSvnkWBRn4nIXNxmoycUcUmtX3KIlFa4oFU2zaIXUd1zHVKZjypWH6Ldv51z0VX4
GpGLGgoh6zvsH3ZrNNHRzTD7DuXBGnTGifsze7bXbfUNDwnolhdx2tUHlc6n6ZkTk0CI1S7iQFi0
sHGKMXQk2QLw9U+FwNidoZKUlE7FnIyR1m5+GuDqvmYWsK8S4Ju5szjPEH+8D8YivmE/tN3RHsV7
OyAYBT8NrCdDFXldfS5+hHFY4B6CGaL16a/v2WszxyHePPlYM/1vtBNmA8orfp8ZexYC+01JFONI
EpyyAcZuEQc1N7Wd83M+MccRYzDy8hlnQrA2lWFdHGcpjbibpHwJ/TBDIUX9k3ozY20AqG/BIDQN
uaLXalX/Bv8ebsmStffMFmo3iu6roFdctjEvpGJJ5oVPQYwLv4JtMqYGA90oKpfVQOxYCgQgOkSM
I52Gzcdq2r42uoWF61rVNG7BTF6dVIgM0ivjHXW06TrZxn4UnRkpsJF7ZdzVZL484P3EPEuZwDtn
Sqa36s2vVnXek4mX8ZRMPEJewaN6JWqdlv5eXVIur9NpjENO7vyId7Oe6d5JDrfUOO5C6MCkLwLK
nkFu/tiUYqvFQwLicoPe/wecoCZfCSer2h8BAANKyw4z1EUKVdhpomP7hJY67MglyEL3ATmiuEn4
9+s0Os2oNI13l/yr3BJONyvG9FXntKZsDPWSt3rUpvZhwuDDgFlV1oo6RTxUiziSeN1bh242MNMV
vYyz8SOdrbEZyRXtZ82YLFmDcq4nbnH5JsocT0Lf6cx1T6H3r/wTfdpt9xW/ea0GqoPNmrsSEkkl
SFivOKnCgsrABW0FWNDc9kuyc4zF6aTnS9yQiGRvbkPvlT/dWwZ9v9tvCESAQEqmO9aIDBZAsggq
/nNoQamtdQTm/+LX+KL5FZ8/vtNNKof5MJHPnauHYEnPPEB3PZQf6NhaGUOAcgji3t0PihcMa+YL
gUHycCvMQ5NGX762ct4va22wZiH7gDHJAhiiF7Nktljf0uzhpPC4y2JVbyLlo/uIOZVPHqyqChdZ
Kd+l18Fc7C9e3gjygjCnJyWssv0l9VKXbKVt0/nan1CNrcZE5nvOg5uRlW2OyZ2Vk5ACYpqxr6l0
TleG6vGxWtVL3E1LRnsAEF7JKH4eppI/uqdvzuMJF5f7/9O2bq5QitA+fJ53tyy0KN+CdKMVL4v3
A3AhS0N6eB7Is4REKOL94JlcQ/DvkMuE+Vbc/lGI72CQExlQstZMNOQRwTss6uLaR/nNigzEMOkD
Khh/5XtgXk7hywyMF+0FmT0ducG27OXc5bjSa9wuSEiaWLCmv31jvvzWGmMlnpGt1ateNLtT+yxE
2MTwRj+S7RKO6WSZmkEG0rzqnKiUw3cE7tIPzkZtxJunDXRUO5f3ZR/pFZi6tgGBrkT3J5eg4gVi
GnsgV31htgaCUeRB1uaJsq6YmAmdP0MC8xN/R7VxvnzfuvAsqXC2OhvCCaFcQMIFfdTLT+PG8XuW
y2QpYq5mEygHXOjYaNpJek84Oh+obznGCdPZWHI021ogY7goDIZCdmiQGCleSOH42pmu3PGypPOY
fWXsAgK/dK+TRNaJTou0AwKzOdesZlZjGx/wrvONjIGIYuTTPzKTxji6LpNO0Ot4VLavPXsTM8b1
CSr3IVk/fv/w5l9kYXavpZtJTgGSxKTcP8J7r1wJ29Og8CnKntWvs+sNO8xiOgCYDvs83EYbWf+V
xISrmKkrBrHwrUE54AhxEQVWY/qTpteii//lO22x/cVwbnzG3/tLFV8RsSxFbuWonQKjs/QVc0Zk
Asps0AJspRqnN7op8o1HOrkfvt/YwHLocrUhxwoZAVf2RU8ZGsuB2lTQmw63qryrSvdt7Z/750ZZ
GIRhWKLRKj0CaQDGaewSKVzGXQVECDhPX4tFow8JPkhS/fXNpy6GyGmVe2SbZYw/Y6nKGFiblVku
J4ZvLtXDjUjktSsAT+TXvGpmkto8m0sO7Ol//LLD7B3l2rZDgf1dS+x7IPlA4u+NqzawniyvnxGz
af05egbVW0vSjR5xVI9vyNBQiPoEmigT0MPKSI+UYBNdqNDoFtGFuwkqT1TcLo8omcohmkAOlpI0
aL5LdpvZpsN+Qvw3h/IQcG2XIDNso9MlViNK9qZO/jR8JnT2QdfGZONPlTJQUbfBKByylxQdpEs7
f8UkdFLhYcG8IfZ56JuHJEqL/lx4Wj4PGW93OCBtxco+1ynKt0lmODNi42qVct1q3jZzAVLaxMiu
Ln7IE0AxqjJ8thTQZxa19w78w8c7oNoWxhJnPEPCZuParo5eotBPqUYDzPAwD3U0uyTvL6nmlRus
zHbo3Rv1T6Q2m5ONU2Dc/mXs7gz7Ikk++bCESuTiexTyu1yLC8zKvHEhTtSy06/gMIofrDVZpBFh
nRXDkC/wlDZm+21h8hQ4hoeKLpSYDD+gnZuw7dDWkvlVNJ1PCRYHJoXDSpeBZk7laGyaGRJdEdI4
ZNILMsg6L8Fa6bh6DdJF8Cdd3MDOD6nTANbcmJXjQju4nHvztqjeqgEK+MGbn05QJtBkBOzsp7ZA
eNMCZd1F+SBBCgGpfWp5MlAUDnR8msmTu3EuJ1F5zp5RZP5P+TusArimIBEMPZR/Ci62Wa43BnZI
+L112xCBv28UYkv7vzgp4yfpftlyVj71LXAiGw7qTlXq/drC4qqQLhOmamImmJYC7sjmuat6less
ufnixyrVLL5P4iZQT6e8ahzoS/SV51BnkkUtLeHkm+ujzWdtvkG3i1vk4PMg2n+4MU5VaB11jIBS
cSgl9mDgemEQMNkknG9rLrzuATMKg1xgensSJZcnfkkK2ZLha8O7b0m7ZsC9sOy6SJY+Tzgyy/cU
8RFgcYp1QXzPzUrP6gljS0ZWsebrgkwqsRL6q51VAX9fzY4kvz8ZIbR3eN8UQTcmGd9IRM8CgnPB
Uy9WpybeV/6tFfQihgqtVj3BNXLRu5ou3KsXW4tM2iDKYXUNqyhFKNv+9lkOKUACVV/NDLXvANWx
aA5y+z61ZwEdsRia7Fxh/ZUTC73dmum1cHFKnUOE3yYgt67MGGCZ98ukQh+bOZiBzR1kvC0ZMDaO
2ps+Wd/G8LinFXmOvpAlnWh+ukJMa9cber4jQYjTnnGJmqlkydJ/h6eS7RoVoAssN/o41trMkrvx
LlPTZLOdFWuDSJhOtRBeDAD+Z5BKFz+xguPqXXdO/w9XXtBHepY+NCtPSpolU3/S2a4wltAgLP2y
54WwLhz54/0tK/Khkh/3Peaftte/QDZnyu4tRmzNmyuUMCoCgqQJHJdi9+lgRS31Es5wjc885kvx
nA+EgJt+qgpjZW3y7DkGMKj6JpcQ2dJNAjsgG1ivJJyUldhNrVtdFljZoVK2sRFkynClTvyT2Uzr
0GHxGKloHFPgw/K6K/GMZzaecreNYnawwOEx7PLgFJfUjzDvGuu0hDo0nYizkHRkznHkVFP2DbVF
kYReHu+Nvw+eB7eayt0CKCkz3YSggizU747JoUbFFYy7J1sHRviacG7H4StpipHpZ1A26pUhOoln
Mymo4jxbGsZdEjDt47StlGAmMoauCvVYSz/+7haF3dlZA35stSItimsapBxD1U88OBcOvFV0+iuJ
R/tFKGkU1ONRw4tCJgA8BWweQ7ehNJniDSffEuNFY19cyWSqAjF9qg5Dn4KxCuHme1vXVLYUMF25
TDyG7FfOhFuS6wKiaF9+ZkQELKPcdI1RVanjSu9TaPvT52GHPeNe5SgtpRXOYqrExslAtfSDEuWH
y8aMAL5pVn4yQmvEkW6V75J6JghFPDm9wIGB4GBlUt9VjC4U6Mxw/Iud3ltxm21t7ClW6Z2eiU3j
+Xg8RUaC8BL4Vc/AYypx1x4yPADl2cxfaT+uGmAdy5dZxvfz1+32vKaENW+h4+DcoMLAWuGvX5K7
tEkibIH1RAVcPa4W5LDPe4rHrl+TdB77epzTp/I5enSaV58JJ0HaLTTyqQx3s3StTLVCKFhuAXcy
j0PqCvsLf78+DsQjbu2PilWYdRjQ+QHLV6pG5eX4dea9Xov6I1GNSavkbjS+9X4uVV3/J8+7sAJ1
uxbsqNER15dmGYs61KofLQ++EOJinYqZMEwrpnM7VZDaO7VVJIyVuxppi4WRnxLpiJyj0fJOWDE3
QTDAPqiGLoBJYZgWNQly+Uu6wliVX8/a9TaHMIYoDSs7tvMVJ5Z+oh2upzNfyXgT+cYdZu8bxjrP
fRJRFXpAbpdW0c0TTmcOyFNs3GLmAp4SBnnbzGIQFfqMSJ/to5yKlgne/H4UOlDsxvhyO2webL1S
7AN0ffBIASwT5kNxIQbAIv4AIlvvhlOeaoTKcmgBJ2VjEzYvA5rLtk5dgLT/S3rKAW090lTnonBE
4Mu2nS6lGMobzIyBChgEYP1vbv9YOVsCm1QGMnak6fseBJR5w3h8uUtzpuwCaD9BZ+wn7ZeT0syc
sZmo6lu3RuMYePZ4nphQ2xkXu/ioaNplrVkNdAaBDQuwK0YOvWrHbgvp5PxnsNJtTcyA8aPdJLOu
nJdu+O3QGSPDDPowkGZ8uU+zDsehibeRt9ktx3dE9zxko897Rr0aDVMyddN1eyXMZND+WJfmHBJ6
8BD4nRPUGxtN+Cawc4dc6i7mgKonHNLWk9lV6FQjwjfHXD4ejoivJXz9/MO30+r+LsNKSeQGPIV8
pwbi9J1sMQQ4Z02ZjOUoy06OJDGrMFfaxWyTnrJYu1hDc5IQHE6MgarQgmy8huEqKnsWRGM23qp6
5lsvRBNnHqruCPSXvsCZ48iK8G8l6lj8ni595ylVGBTsNr0hpLEPBduYCRXSxXotZpmAkcrP3Jwx
XPYJTOuF21qnGkQL/U0ivZXXMzA5wnjQ7KLb0HwfLn2KYTR11az3olOF4SaheAgxk85Sx4d4jd8w
mVe6bcbTTC1BED0uncMILEC6OijmWqEIVnLj5+gDUBfZ9ZATTcG/P9R/Gje/o3J4PwOGwXbUb1Vg
lGqoq0e+jmk1YEy5wK7quIVHNOwqVxL2iyflM/LRSJuFCX64j1orvdS/2mi89LpEyCcF4Naxr5fx
nBYXbjLcOYyArjI7T6CUxhyj8kUzXJIoFBsvGSbOO+HvoUF+5PgXrTJvCJ0ZWhGF6lzW8WzlivY2
q1S6fNw5qmJynBvvLJmL9gmGeHe5JpoAe1KAcHDoqC75jDyJVKOtiJRDJhGnLmNgf+qv4FUn0oid
cQM++YVrI9sGXhnXlOVi4Hp327ZzhmhpFRFSyQQuhubCLRmKu59LhvjCGWI1NKNJDh4OxvL8TAUO
sPoUGrEaBELDYP60XAzwAWig7XJLDIudX6uw1l+Xzn2EY3ygOVlXLQ2RVjR7SWbm7cryBl/0Doxd
zmHbM7PMKNuY9UgZ9AMlGhA6UqIM1uhAAVThLMXHvIIvCEiLqvpLCP+c0hNifWJlxPXREXxBQbc9
MHpvKHsX4n8+odq/pN2vX54eHxrta1l1A2jtny/uU/KIlsq8ukCS8Z1XBzSdXp/Z+Qs1DSieGubJ
G/3yykZUBjZ0Om+/xByZaTwefUt1RZyBoEjre6p7FRw8gGapvduTYKTs+V2YOTmOZaW7zLLu62Bm
N/wlnwJAlUL58pK6XCqTdlMnc6x1DlknlueecDO/bMbZx3KFrUVR5POKxV7IfPKOTYnbnHBjbBTR
Pc2qOISKJeEPZV5cj82LhU4zC001TH6va7tXsouHoLrAGKqtFhsxstsxtKXbUBpoJj6W50b1cW87
tQRfOunjLvzA1JGlnv6R9AYCkjptYnI4R8ie6nyWe5T8hL0zGKUtzMz1o+49kSwIZetiWTGSe2lP
zGbXEB+QMjt4MTXl3j+Sqk4YdABryTEo1NqCqRfHC0OAXIqw8EL4r5+OKjQazYpyXDjoayy/xxqM
1gO1iH4MZ8d8Tb6klLTWFxG15qbzCoOD9fMsakiQVp9kO0u3CDX0ldL+FVKNdZBsfGFEa5Ea7VrM
Fr61A7Q2tA71sDfzExjvW+h1eRoL61XOdM+5oiHdrdE9CgnAy53Z9+M3xYKcokacMxbtVMs3ZKej
760lO6pkhwnnARssSN8um0NhK8ZT1ylsYu1Ebpt/MB2YcqQ2Ia5xP9qChfqT22AcyhdXk6Kr1dc6
TnxPMPp37hc5pyxRC0oPo6rsAZwJ+Y0HJQnEcBTuYgaDZUKyNW9eTzAh3IQjkcBg3eq5BZMqQAja
kZgkvLEfrAMrDQmkzynwh8/M1Uh5Uvs65r4YOE2zgwke13EFRamj5BvjhqF+aV25Gt5fxULdAGC2
45MrwiPFWXK1TC23Z7g+o+U7shuG2yAsZrUJBqsgzESrynps2Dnco3emREKnf84TXsTjMTp6/awG
Vcsk8I2ZrxgGY6u4or0o4nWnooCdKOELdHmYuc/xewNrWVxJkInvQfB4XNYvlPJWWOcV3g3jOZp9
rWqU4YGHOS3YyJCmeVr2Q501yiBktOgXgbXOtjiups+icmuH2SJVY1ypMzPRM+nx0fYARtW4oI9b
eHN1MV3hn4GQMqMMk6grFeyZsjSBYxXKIGrpIqV52KphrPgs0QYmttaB8U/w8bd3Dsfv3eu9T2o3
3Z9qYCRtrBR6Ldi0+ThJAHw0cEqA8DiDF312fk+Vzjo+xMSKNYnhu7oWJgxOwDVM7t2YXBFoxyg+
ekvcIXUVC8/fQ1GAf80xbiicuVA+Lpw1dxgeGKjPo4M2JYIJzEwM0otYsX0aLKW2OJnEHwZRVwmz
CyTUEj1uRu1O+tIkF+U/xwU1tDW17XVJxBq5nGyrHIYwN7qvE0UHvw1Fmk3wAAFod5tSwhxEmVxr
rGLU0NKXuZ6KZDPHNrGhoqzLnfB+oOJF6Ia/WjdZQNGSu9ORmEJA1pR4xgqyrH5ytWy3krnGMJS0
8Fdt3x+j00UkAmSVGGTvpL76gZaXbiUCb/gydkzCwKy4/jvs/BkoYJeRXcm0HBnhOAY69XLHr66+
GYUQw4YtwlLMgBtznYIrDsZ4NWJQ3NDYEjT9gdUUF0lDCiPRiTl9IZgRL2lCIcFP9Dd9unFhCti5
UWTfbSFQm2JX+57OKQDksxFHZPv2BH31MeW+SY9uqjnYcEcOB1HPtnxaLuJjr60lVOnWPrDEEJMq
qquJGuDzyNxceCL0VunIgMolBE5vK0Yae3OwNfmKUJNTAjyto4wxnsDWDr4/6KJ8ZfUJIrywWDs4
HIENMqA9hQjUTYAnoQ8JbegeEtJEa7afcAZmLnHiajWjxVsob939nW9sIbI+JWCoGxGuSSOL1Xi0
b/yl31xhnoyPIsETLzWA+a0Z8DhnP+lfOS/bVahHVTDczZqcWPV0xiQkxfCZdFlZm7FLag8qQDZf
cHjgcZZI7MR0usSsDbT3M/dTCDLGSkZLOycAwvvxcw7Cji04xOJXW2g8yayWhXasBaninCk6725W
UJn66zuFx/cPNxTketokJHWKfi6/Hf4bvvB4sQem4fyur/QS8wta5nH9ZndOMF5UYfoQq65E+dhG
LoftNyIfqsOgQZWdehTble3WmUtMh5ywhAkR+HQGursFLDSK4WmnHrHUdb7XZC1LNHMtjRd7FqMx
gYWCNUekwqvvy/tJO6SAgJ3/+KaUT9bhjrNWNjiJbWnPq1yyFnViRANkQgUHsteDL57LKjaRz64B
kBcu/L1y87/TbSwlXaZ753ALvImntnkLW8hJ4qKZvLjhZfVD8RweXtG7Fo6jzBYGf+Dw4wSII5C3
rhXfdm1tFimfCdqHpTElWu1T6Ik/xDYEMzS6UJ6hoBXXrhVeOcKpmkI/alEiqDXOwLAFT3iTaeh7
NF2VJ37GhqTum2Uga6r5AsJBnUUcLMkCBAd7Oyw6zDidlK0HDHx8PxcCjH4Q3flfxCfuALJvifhi
AAIcgUXugKu5cLj+6jnLuwZAiEi/afEFHk+qa8NSIQ7KdADdfQ4NAqjE8DlXRT7DNLHOAfQ6qaa/
UGovPLhGX6a1K8kY1ZFCnYd8X+fF4fnctLNCEe86zyfO1uu3oReEzbDaJ0Y/rgwhm7tEdMr75hNU
qsc/N1P5RI6HNMHCeFHGjPyuqMO3cw3usFl2hf59fehcl/W8xnFstFoGrngwlV28fWJe/4b7dcUJ
Nj3o8SL8p52QZ9RLPStcjYcExQ1maBrrFyOYgY5K27W6pGSexSoPWBJwqU/vpDRHPp2eVtApZBfd
mxuo/TRWPi1i96Ey80Cq6v/oY6xFxV0A/AEc++t8Enq2qtc6m0fNf1/R83v7EFhpFIbb7kvWbxLd
HGpYnN9j+UiHTtuAGleC7OzVZjWEqELJF4GP4NWmWjsAu2uDxFgasamJGU4e/nfgUywuh/xYGVzV
8OUQCkyAbBe6sR3/NWJMkG/9jKUPlzFWOSIKsrJNnNKpX/KrHxBkh7bzpwtfITx3xxNQJeIeJNJ9
mDiO1fXkiygdGAtM3zIAsMBd+e04qjDHYVmUqvOwDEXlY2X2ph6t3opMDglcX7q1BZwXq4pMq7cF
gXTG79u4PNg4Xgu2b6LrjnVB4I8bRAkraO3FqK415Gy30fKhNorh0BG100wUdnMtwRen5RrCCFSo
wyDBtADolP5ktU2YF8vHeW5Yl7r9rEZQoxfiXFjLNqTaAyb6Cj/YlF+HLTmYtciKUfMluglJPp8k
V9OVFj47tSzHY/JXDjA6oh+hAzuQ/Sqc6C9irG+JSbsmKrNRjWOhxU0y+N8/sBheVtx8qzx6+/u1
9dsKC49NJMTeKkIp+qFD23gOnEq+6mcXN8E5LGHSpmtlM3D2q8SoZAVqB4a0SzaF4dp3rNjQEAhn
q12PS3jJJxLIlDz+G9QMzV9y1YqBRjRcGAs4M9+OIUAsXaty3CJj+cSxrUZJAfeDUi0OUwsGmE9T
IkALHmO7xBAzrndQ8UA8Ypy1Mwrlvd71j2MMfNRLm8u1ju3h6Xi7zl1xGS/yYecOe80WaE325BKv
5/LaPTpVBEJmducqWOxLNUlMVsUXkikxMzjVEiKEqGGJ9x2C3//4H/2baCdVyAqgPEZnrd/IrP9y
Uwl35CPPNnjuN8Se3AQPyOoUshfnZCEC5TB23yHG5gSn+mCe+MSblTsoEY0wgQTcH/fd9fUh8FfE
IpRIdF9pxmpCScM+hS705JpdOhAqdv8erUZ2xsLaNQoU6k6OhmhCQcjgSYj59n0CzyrBHq8ei3jJ
ahg6hLv9ZPeW+99nCzAXV9c2zzUM+HbRk4PONDLVMLHK0VoYhiFi+xtmvJet8904YJHL/69SzIhS
uhLfAkhWR6T9pSN5VatCfxp4zEEjzl28/APbjGiQpYqGFmOgPduNPd1dR4JPh5mE0GdMR50X6uSt
2gqOqUFCxGA0sMSYqOCAyZgXaT0nZgKYVdbswhxvxyxfGFtxO3Jk4958pnPdtmWZ3qhOfPHPabMY
dFjV7cfp6RCBtX4TgLEGEX3gRkHrPjm3Q52WjDCLzyHiTvS+lXIoAtFkxWS6mopuN5BqAR3tGTdf
2el6Mio4bvvHLZDGn+xi1vtI+vZVRSaT3FEhDXHENC91fM1+Rl4jCub+jI2oPvloaP8/mlR+z1pr
wsAcloVlAnrF7stWwTycuHNuSe3uOj/txdSmGSU0pMX4R+GjyM/Og0aqRlBty//Q7Zf2/qcRO8eB
CSGn3vrrvu2MN+rl5dHWteIeignUy3w0GBFveECkRIkihqcwIYoVdymZovhkiwyNF4r9v6M2sTlv
vo2s5reiILhAGJWJ1wao4Hm4gdyWlVTrcvyrJ0D+eT+ov8T7rc6gt42BHtsW+iFR1VJmYz3toRkr
6F9G3fF/Mfzmv9Tx4quoHy4Bg8+QKNLfsp4r8R+pJ5UReasflDkBHwmNdhkwpLx590tiD25hpeAe
xyJrz1tE+tUSw9t6oNiQDHx6cydQdkiIilt6FGrhUw8Wrv3KVpkgsG7AEXr6fpZPORfqzpusZs3B
lhC6jbXRi3HI/ZZ9bzxD68E6lMPBmYSwxSqMrjS3U++hrtRDVClM8HG/jy4Ud3ANk5g/yyHePbbI
Agb959JzkJYRX3L6UnPpAxHXl8lasMcrHFYO0fzcCmzdjjJP2ZznMaLLxqDyrSnaX3lN9D4OY0CX
HrAcuVRYdsUYqSk6mr8Nl+OeU0IpF01nOdcA7/U+CsoymSZvNcv0PMNCHb1Yw10yET4kycWhiDKS
7O2isjtu2SfMkPJZdXHV9+EMGVEshw6t0rPytcZpbWo0WYHreFanGtM0EFyZ5BE+/55xKcAe4wTR
IfQ9b7wwlMoKOYnscz5os4sxInTdGKya0W7mnNYv2Tndc2vEN1aFR47Ki4m6vVcYQlDZ3NjsYX3b
zF8SrWHTUILFBSVvv0bTp0llC7jiQr9RFriga12gF68vxlbGDmzLCjzBGGtegojJ8knoHukS3MgJ
754AqObsLtCOgDkZxbrRNExklK9a8dswKGKgYQdBFBs5pDT9dMdeaUeY6zyTGITiup247DUIhEO5
XUFuyF1RV35gSp6WAmk6CVD4SE/upQwH1GU7MCO5/dOAskugbc3wr4ZzLj7s/qkAbuBjxWDQ6ZD3
6QdDHmpVWRhNXbT8cuSDvEQ+iwModMDrigIssWleU72/US0o9Lhz7uEygLx4Irg8ym/r6DjZbR15
80lfkRKCtbJ/Q1pb7Yenb6TKQH+d4JIwmokHuwTbMN76k18VwfAu6keSztJ2Nm8EQiS/BpU2S3Ln
DFsHGzM96InhnrUf1gNfynmEM2xoGD9kvbIqnehmtOeS8qyrjl1FU5ODEx3wYyHU/R/CUUgDiUkM
3cH4yQmRAwtUGdUpdSO5YPkWcXIey+FdOPCUmz635Ne4p3vhdYwMgCkbs/dMEthhe0VP/n99aIuh
ppem5Hge48R3f6axX9PS8IU5blgxkQLxJ+r5p4U0fZqjZ2wV4y9kt+RYxRVsQR9g2VjMgNQP2TjN
2jhLdRAlwTIaGfpvn9r7PDmiokpzbhsw64oOpmdHK3etT5U4YyfeeXqn5RO0n+qMoGeexYG1WQXb
WDsWi5t/WAGAuBVzAI9C/U3/Eeus3zSGOXULBFH0rOWNjerK4CNT/GRwjIwxqnqWFj4PWhS/VTyg
8LqdRHgsGEbyyZYofo6IN/vLyrpqd1PjuZf5TDPkFaYhECilZw1N+TZZwVYyYsn9++q3BMwo7ixi
daB5ePEX+btFxSiyDVYXKIEOvMykiHwrUevs9bQWLqQKB7pizsarzyS7nGavRJPHhfBIwx5b7Tf2
kOvjkrkcovXyDTAlZw1QFzp0OkSnmAAmdDv8wMygV+ZjRbsu26+wZjvciPgnFUsdGjUvm4W/KE8Y
Ty7h0CH1NHqKM0esNpXrZiOlNnWfo7VnfsgjXsaCkI0wBbAPJNUvanY1da0SfNfvZuRgsxXJxo4a
KKpljm5iY4xVmAnFJ4e84/40LBzpDMTwiijq6e1xnomV9rwkcMEgTkbig5FXOf+jN09ANJYfnJ6i
vF1G+eoh2e/kWc1Aq/t8+tz8WQLhWc9j5OA25uPaiOzVqPsaEhSMGl3OKRNgvXUb49o4YAGdTdvE
w6pN5D0Mbv1Ce+z0g4bTqhW4E1IFljml6U9io5AFVqkzrhsk7a51H7ea6suvmy76tsOmS6IGeyyx
RuK7ASCmsOeK3lA0M6F7bHx4hUIncnCDN6xmuujp4hkMO8cSg2UUw/wGyv1y0Kij9PPt1Zz0VOH9
egYm2u25e5GWkFeiTEf3Nq61k/lsqt3p/o0n0YvwdVmVVh/HQun+oF9GVgpUxzAxPnXZPD9p3gHo
5+RFsGxLYBHs7844ePBq5i0Zsi+8IU7EcMl2NaXOb/4/s12mLY8+qpBWmqdeDSChTgIOweLzJO+/
pZufMlnKarM4rScDUBeQ/1w/vzbvJwr8FOEvNnzglwQa6+5Fr6p9mX9s0mhxgtgceLNIBfzNDlAm
9rjJT+X/vtrIUDt6pAfPJPPC/LNxEion3vSRPZmL3jDVIOdfMyl1oaGe2MS7AfOwz2vqZeyFuY8w
F6QoOvT83qVQtl3n+KkkSrIPQUUo8nZxYhLGzW8TM+bhS+77ptwsYq6ckqEZVUIafq4NSs29qB73
2R/Km4UrQ9/MDTiAuKOcRBqB8FFh91dM0AVbL27Iw9+2mjF/HA2jfphYlYUfDNUNjk8MYXUyWDHT
KNxef1FVIUzRMNe7LDnvutVnTUc23QEMgP0CZwjIw4QeYpWWo37ARaf55iuuQqo04H5i57tmuUxX
Gei5lhv0sNarXyW4KrPN0q4uyQt1Cawp6tsoUahPKdyyDCookUd9fS0qoZqE1bjhuOnqOBAR+xB9
XSmVKEnwBESiimIBo7blQXTNulk2GBuy0BYKMeXmFgfYIPOrjUik3pgkyY3l0sd4R4IQUS4WUCyW
7+62ErUzpNgkMAKckIK6XW0Ytla52LaGjI8YdxybWr0IVjg6cnHdcGln+kVWk4kJD4X3qMjbyZCq
lcuMNCT2DyAgWynqouST9r/HS8opmUUqP1bJWz5bnZN0PoVte4o6E0PiF+jqOFz1QMHxVC8JeAqp
+MQD1tbpiA5Tlifo1incc+9unTvr2Ax19eQkDY80Ma8te6A4G4K4EQZxvY1dCS9nEz798riv7Suf
ndYh1b37fXCedYExJ5mVccXjYkTcxeomXWFsnXu+Ul+tBJ26UMu/4kGwJcrt8XP1bh0LUC8neIEv
pt8Hf3CUyClT89098RRpG6hKEOawddjPd+Ki9/eMh/X682Kn2aOpxWVQXO0QWVVidD1dwoJdX617
W/zjpVVVM8lksAuq0opKt38Qd1cobeaZKdETciyYzPN6WWMTf+Ah2fZOcpDNGNVGWdBwb78HIQF8
QIZzofzVeQbbeoLeSUnK5RUFGpsrANm7i9GRJskjjODUP37Ao+6PSawWiaiQE2TX1RhymC/2rAzT
5CUs8TuQErPteUkddnTGI9afqPZ0i9VMlRuq48DN4GqNJUrwqD2B5eT6JqfwCXLVB7Skbrfefx6D
53E77c/PuAsQRTWmzloeuwaE1Y1CEHEFfs9ElVFFZU04v4i8uv7DjDZsqk4njzvqftbS3H6yw2k3
KTKyhbeehk8TS0CGHnAwE9OagDnf4Nk9NHXCqtkHolzXUYrAPo/jl3iYR+uLpjseDh+LPSb2LgoD
W0hdq3iozYQZGINxftON+BGS+QubcgfdGZDsnRlbImSdmfVR6x3lZ9qi7izI+sJbJ8uX3O7jHAke
v7Vceeaa8AfrFrxXYNqGLXXfXYGF0EZ8NIE38PfGoT8P9VMpETl8EMwH9bfC8H8kn1AWmhV3VEXl
y4csEnrZBBWMwibNPQNAhvw4F16Jrs9qg5fVRPfCcyHFFOQB9GNYEK7Whz4dw7C72avTNmtcr/VV
7eoFOhpUwBbqdSBamUArYXQldOiIA4pbrw/PchkYdYrizOWd64mnjC59XsJPw3dcum1D8EFaxJ/8
eTEiI1hII94HKA72NlIfDI+tIW7D9HPQcegNG1KdZh3orqOvyghPhE20rNt0VJyygC8LpZziyA4B
cPMq+kix9dlWoNotZAXnAbtwOt7omyYJ6q31QcjxFHmLDf//inXBPVTIdTtMNk13U9m0zw8/J0wt
iQPh3dunHAKE60ziOqbHGr2qowc7v72A+UF7Ha5XZXyWit6hQh/ssCi+BWleoy7HLSiOU4AlvszT
pTYN+/f+DRLMc0SqAV63Wn4CW5oL5BP5/X32WFVj6rkDl+ojnZjUGlt6FYIgOrozcEmjzuJSmC5x
Jgiho9O53EqTAHzRTI1oFVBGpUDIBIpujlT42cEw/H8AwMh0qjGpU5FmKRbTP1Uf2gu6qt+i3VeY
P6J8UzPa1OjtG0rUpxsQG6SKQ0WDPhPiCdfrfTqKFGZd/1qDm4MjvTMZkdmi+Vh0QQ5VMHgSoNZV
iRbmgV4Z2PmYaoQaXnhh5OifQTZEMpE1I9MPSbjxKPP7Eq1kf22eIz1GMjkYacOEYJcy1J37gQWq
0TjirrjALVwuz//ZNKrKed9/8iUG6ga0lmRJRkuJn8636yeoOoKytOXFQkiXo9zKfY2yDncShgkD
w993HccDiiWfKMETzf+vvB8h5U2TW53qEcn+WanElW8/lQPcxsirslRcSiOCSWhszArLHn/qzUQW
9QYa6pQ6dm8kIfwYbtFzh+8WQrvdj9xiP+tW6Uq6TQ40TLw2qnyEa/MFuu+ojeJV7s3ll5Wka10k
qOZXIPfhe0mOrbWiV7lOTCwpMFvppDr+LWG7tt7wqt6dlQT80Ae5b9b8FwrE2ZCUiXpI1IsRVQkT
0UumEs10gtQpy971eTRwOqioPOf5PI9dJwitlH8hE+miU9pKx2lR3IxClU7OzqjyjZtonMLej5iH
8aYJG96ELAvIJvVzsj3/areH0OnqcZPf0+8cr4tvof1+zIKdRetPI0BQUTJh923iSyE8PreHb3ty
47zbkaNRkGN6Y001DUl85E+/jnsezaPeUtwKXJbOWt6+4DyS5gADG8xLZL9dEZ+vnrlF2TgpD9kx
pHeg2kvoHPCr4PIQFdDiRGi02rhNMhHzRdLwWDVYRWP+Z9Rig89uWaJcceysD6VnAKF+zADZdJHx
Y9E75h93PEUYUn6lCnr/PuRhWNwMv7LPWZGg6xYffpbtfihR5ZCD5AqioftOH2fmtW8aCk7zMK4X
HNsaSTP5njj5BPOmF7LOmvqJz4lFohU6nAfj/l+W5xehs1VkYK5SJOxAKp/ZGU1rTLytGc0/1y7N
Sr25bUx9ONZ8xBRDlkHG32AiCRUUPxavljMz/zNbcMgxA9E7dgPSHck9UXAUnO69TPtWssRsS05c
askbBLlYWSgl/czh6uLCDOBzWnnrdH+Ghx5HPNkx+DgHOt0ggBK1xl3zG+u2Ovk4vw4dsS2sKJKm
dRkgZXXa2fWmfA98fCNiSqEDgUofw7q4c9LCvfdYjl3KcecWQxEyG2btMdioRl7CQlj2i1C00uda
DtfeqzloEpyOAIhfYfFk2BrUECDNneIKfkcMlELv+wz2IT5xlVEC24mq5pb+vuoNv/CB3nOoP5x9
Woa2RIHoE6NSsqp7EhzYrqSkLo+fBCwMvJ7kqwOMDVY+8UbIr5wTKJMR3hKYKjTD5VVfAUnvVdPc
0rPY2WpPzdCghr697xpHv+1pCDHEUNL1uGOSmacwikrVcRnFIZI1+lQRfbriO3ckGgLMvr7b1kkJ
86qmhxp2BpI1f15KplxVhRs4Y9N+c2czynHoQtyidMdHIazF/kp18mSLvl2z9ZCV8xNzjcd3VPTy
SNW23aCFI3E1LGuc3IDa+/crmNEAZjBi7UeOyjt1StiOK4iS4k+mdz3IEuf9DvlBGGz5f/Wgm29D
nUXpfsMtbT1q/1DF4QIkQYIamdupv2wSNbHfMJnIKjxDjftOMO3M2cS5nlE+a8HYC56nXwn6qfKW
xIgJeeXtFgjAwvmohx0j9ozM42s5V2MDTT8Qwvo7SPfcmN3oMtnJhnFWMeXmJGLeI0LSz5QUe/Ah
QZ4HJc8m5mOnk30O1Gdr+u8yNyDINugtf/xMz8LXlG3OhsxsanL32TocFN+IT0okbLKnEL61lbAp
ipP+UQOnfAapn5rqdEqYzUr74Mi1ee1BCswQuCRlRozDWA7VgJNvCpcKXxiDPKi4sQIlNFeust3U
GOlnx3g+3JcNuvDCkSR0wE60gZ8/r4AhuQMCcjPd0OGfngAV/k9EzzGsDhQiOCdm2tbGsqbM4AMi
OVyi8U8xzvmxFW6MftQ3pNCtu7zyU6kU40Z1fkrCVF+TncqHTjyiXTaibsIFwP7wvpRMST5UnY1O
t693kgnGBdXGLBzP+79vG4A0Yhv50fSDAFSJdqdWy7ODavBPszSM2nemZe00gSmIsbM4LeWFvnIT
ELl8jlB6/wE7L7z8xrWMn9LKoTm5jQhiLkp9yYFfyv5IM3UhO9tYxvQo5kWwTjU0XpoGrGCTOEYe
HKmU9jtwA+XJAWXpuYQwlXy1kPmkdqYTpbNZ25t59z5ppM2aG2rGLcKOFwgC2W+MeFq6hcV9Lmgz
jk2Hq1dpE6qbih/nnQ8dcMj+yn9lv/PlMFxku3XfgZfjSzGBn8ij7pV/xaXV6i5k1EQAXZ6orTwK
vnKlfZNXEd4rUT3Hhe3jGuhPys9odmGI49zaEHCyB3D3UuvyT/ZqVQFsogKOB38p2qYf4q4B8Thw
SeaCQwL5lwb+AdzM4EgB55dqAAU6wnKd4PyJNbdA9+LlGesNw6xhUB0EaJeueXBhB1ALKWQR2NMF
WIvQiv8z0/qnIWxwbs71fNGmItMKRYeTiaeEzjAv8/XX3D8rsI/Cw5+lcvHj4oQfpPN+QxA/ahxU
Rtu0kVcLyEDtTkE3tzk6MgEBizorda/fufy2zzsu4uKSqJqfqzTQt98O1slCX5aUpp25Te22k3Ww
DvqVQgPxFYmlP5MAzHOzXaAbbZkYKV3eiZjl33A1A92xtiklfN7OjfyVZz+Xkq5126uzXBDufsHP
0xi+bEXZrWJUW0/kYmyKQjesiyI4Nkqx1D/rxar22Hl1GGzmi5LCyqyG31N4K3H8E4alqOu16HcU
fqSpOBq+HRQg46I59tqhB6xe2AA8we9SiceL15pTz+1IaWJJQoFv2Pvof9sJ38gJZALJcIQNhQSr
D5xsX1dUHryna17UgsnfcIr6JFgVeRwwWKD80/oNgs9OnQjEGQ7xWLyeBAntK13a5eKlryeD8DJL
3GzsBXc3IkFIUXdj75eaiy5yvE3VZ3RLbq3UTaLSeBGIDgPlG2plFZkyrE9z6lkEPpcgkzgSEZo9
X3+ioJc4IeTujJluJqZSpYV9bFUFiVgTfluNuYFZLqg2zVIJfXr6C+r436U084Tmq5jiPbRWEBVc
5Q4TzGLBxy3mLnONbybuP8pj4ajvAH/tOvVtjxosIbeJBySx8fvoRqsju12IWqaW6+VDH6YfC70L
yk86JzDG0qZ7d1z+chPCOoNEo1QKrGnZouMyCVVLoAqQX3jKKb1P3Zpbqs3P+IYnjeZRn5AwcEoG
aWI3S6djGg2BO28tkFBbQwSG8nuK0A0+OUFEHWRLN4gDHdLxWkWnf5N+S7t46UW8eF/sgEDw6HRE
1C85kR9JHK3YV7qR3+KQkn9e5JusxUlJvYhfGytEbUlz3y+1BTnlyRJ1bvrvAtjaT9gasMmfbrA9
M5V6e3MgikvUJyCdMjDxiR6JYxmoueX9lp5vY8U2TgktvoFrWX17POj1Cv//cFa6WRpCBqpH1sPQ
tSM30Sprs6zJuqROQdwnotpBksvsjVqXRA5NVVnJokmN/62IfoO7KkUZbmVFInKDu4sMZfpYrql2
GKwXz64EHbFSL0+VH+YFROar+jYfrnJBLJOpESpktC5O6aScD+PEaSCRqqWhQfG4MN6zbEbxVrhL
bAycJR+Buwe5N8dp0bsJrMiRrwe+HvtiJnDgDfd/HCRbed9nRsWzyiy6fw2w3rk7rZSfxwIsedET
LD4Y7idN7FwKJ603sGXD5HEAcynMb1icAxgFFXac95+nSZSULyfd34h197C1BpChuuLbZbpILhyo
vGIaXGU0kyvQWdJHrYkJTdPPfsAqkMNGz+vrB5KIOB2XcvY5e/hg/IM2Q/1T2zEMQBJc/JelkXfM
QcAQ/VBJbPHU4OkLw36awzh53G1u6OfXryo30InS+FVldBewCHXoKJ/Vqzdam8YRETlYlKdSGB1O
mGYnyjvkLHbCIhYDL6YxJhMoWKQViMtpGQ/6gYhLut0b5Xdaeo914r/8HOjg1zlTPFBAq/xC7NSI
sxcCa9mTw95fWMizuIy1xuwH9iwWmROqyPYl8S6wugocAnxCRsBMz3XIabKQJchb+J/Fp35yCl/0
MXkuRA4+bvF1tTXz35BDZarELSKOMYVQFc0/VCtVrZqguKgFjXutNS+EJbDxGAa39v9O33Dh7Yd/
hA9jxIN4/Ng3rqRwL/pN+lzp0RzOxcP3UGbteSlIWU/OdLiEpE22vjff3dyBWOTnZjZj0/Z4HWdq
Ik+sTujcTlPKkOkUNdP8id4a9k68B6OiBcy9ENcXYKaKJnu8xMdGP1Hif+E6KQMHsEdvYs12ru3E
xQNjIem868+yGAW3pzdNRDmsToQqCn2H4JBDqq/LRX22mzjgCmf9ehBjWswftdN+63C3hTCIfk77
56ALc5htgpDJ+4jz/jcyN6L7GLw+qo8Mn/31IrpMEj7frM4gkKn7NbpdaWfZqUmdAdsFc4poyUcK
M+WQ6LRopTiL6yQgrD24xTNGNcvOhK1O7+FXAJ00VCx/OSXi5vs6zTvuB1ixa8lJPnPuUBG5vXMO
Dmgz+yD+VrR/eyJTcGgH29vbcAdawZny+F8aqw3apkRF843HMQEvpEV972TgInsbaLzk8ikzqsjI
ftGReqFNPkmZEbVVWW6GNlvZ5eINNBDiJQrbKMMwIQkHhyLYKbwG/JNV0AqMM2mLX44RDaoPdK9Y
tAcri6p5G2mu1IfWC4ciF+WfztYKzSe91vPOsKEERUv6VUwvmEqRREQdP7vOB8/9bJuNWljr10Im
+1LrOR685WkIZz15j39omP+80LpH+ssEoriRjRbY7bxhoCNjVLY0FIsQG6GDaZUT0bMs8HFhBksV
KFp+SNTOC1hcVHSBDt0S8Vc9G9D2TvBtQvsNqn/osCTwsUiRCWkkLszvfbsym3SNwbtzuQV42MI7
e983GsQIKIbYOeV9lY+Xgr9hNkfzMYwXrsEHfvzf5JtFSOAUArSUygSJQdaIFXQe+qY36W+JZGcy
17Huwr/sfqBXUDlizBEAQ8yPLgqDSc1ouTPmme8p1rishAew03nrC5JAbmn7vDfTQ/UbgJD9f7i0
6EXXHCxD0yu5A+z4+Gz8Q9jOqc9uYamb2Lw+0Ikl8dXJBDQ72i9VRkGYC2/9SlALy7BUgCQgRjsr
yS7fCdIIm7MbxvUjuZ0iF+btTGkyCHvdqS7JsVtBaPnbftO5Qi7Hjn2vLQGifTgQC5QJh5wFlgsh
58dulN8C71Jd9h0AfFYwtfO1xkxv/lo/rKGibumrFnVpzqcJzOpjYtI53RKFxkCqn+jmpCowtkNu
s2cAMJM9He0ctSegi5QHMd78SwS5Nuiu2Uf0bIaZouKkZ5HKssMkZq9S1NnH6y7r8EoRyaAeKRFV
gS2N9sRZqyAnkAwJ/VzZVkgmYu+Ppn8NB2O7gQe5BWpgLCz1bW8P4YiA4XRSlFQzUYebWfA/3CKU
wwZq3epekibFLb4yFdZUZGLJPmHwENTfoLC5UA33XWXf/kvc12E+J9qcCaqEceIZABF9pl6/3Gmg
DdHDe5PGT28X07bysJTluXeCka4uZbMqcHBkgE1bOtKI5nBhjIbQWFTlGwO4dykkK6r4XtGKTGFT
3LjVA2LvT20/17d8DdL35mzc/vlMWu/iQeE1QojTNQebCh4Tf8KewZiX4mCNOubZNM+wVcCETKlM
9O+H40b6lEIOxQjl0IP6Jug3w05x3oEnNx+7CuwQkaDwqSZFuC2qaQ00fdwT0sXp1nz0/iWXj69Q
ohNWV3GgkbbuqYBRrxuhejPnxqcyofVdIwbYCzqcCt274neLlgaaWboCa4L6pOOmB7ZCysx0Hh8A
U8TOEDXmg6BDO+gXfQKz/ui2F2wheopad7cfmxOz5Y3r6UCXHV7wiV1sFY6TfhQVTwAv1LDNrxOG
nEiar8Inx9xivqEyRsywQhA7SELd6dbR0gfQ5Rtu36WaIlfjkxLt7y3Hb2NJbEfGFpQbY54v9IPU
WEnsRGNnwsdWBejq/Qe/BYM4PPe2SLooTUxxtvUqOFitgQRD+36DoLizVX5Xgtdr16x9RfNrBeGY
iJ+dIdQSQa4OWtV8+jpMe+xibzbELjexIVVYeFQMGFCXCCOKx/ffdc1T4BgiPKWJJLDNI86bSQ9L
HvfuXlPYGR5rF2DD/iYAv2tUtythJIxkkdM0RWHVUdjEuiCCoEm5GA9KaNtHEpiqUhcc0TXXjtKP
58Ap/dcPlflwRWgZzI7yUEirPTK9n5to5UIChS8WFlU8eIk4rwlhG3vCLeLLNf47kvgCxpWW70nG
FGZbGCONjtvN/fih7WX1d07SYWSeBckqoOSJDy8ZLIkwULqFHRLZAofk10ZfLIiMIDq7E9scc2oU
cO96trfO/Fiff8FJzXlcvBLy+O5BPg/hWPlOsam3sSJ20gHjw4F4/MarocYF+mbhs3WVAy35YyzV
avmzf4lFKPNbK1NGF/4AiCh7VrFeXCyGFD9ecDVNuXSKgnK/lCnBucTjR4QWObW3fepx/FbDHuvw
FNsJxXVfXPpML0tffItFJzJzSeNVjq1ml0cfpwy5WDAtzJTwqfwozsTgabYY+AUFWfxQgBV5LaA1
2/BC1+jYS4LAhPYsRRymRfWcxp3RNKdeJ4F3tmQiwAlcXNO7K+0Ri4rhP68/VoDSTUiAp+UHKMrO
9YbWGPfl+v7Ztj0FIGbXk1U+VgsO9vYy8VxWKFgEV7YWkKDG8Z7eN/w0RiWoaa32ZfT6UyaYzdFe
z44si2WXdhPkS0OUYCweKrSRrNoXm3bur044G+1GfepREKO3539uf4nMIcDAb5seacVqBGAmDq08
nu4LJwB3ZZLWfJ0b+SAsv7h+HyiApiBlzzNGG1h1DzROH6943j/Pizf5cliJOxVcmtpfBu6q/GI+
HDy8QlEjUyZaVyg6FClX3AsCCWWVKq8hpFAZfRkVtRpD3Vht9420mF8R7MNp2X4LFCVBjC52z5i3
6LXIpN4UfWRc60fQh0eIgpTo/9zFOzUgpLBMj8KW6YFNgr2asreSrjs2Axj9Wyrc2P7J1uEh+Rd+
gjcdhQlCCel4nX7K2YAxXMBh1QtoyBmTMAbfzCK+9Ibnst+36mmBSsmGPg5kZsqmvkoi6eacA6Lb
1HnHbEol3k4AhM6+pyQuolZ6zQ1xOHYUb3NfDvwlmeBmuymj4i5MiUn/eq30nBHNlC/1rA5KtLql
MDbcZeMATVJoPJw4QI4JHdHWLH+CRIHNBSSvtyqvFKcwXsZR1eUYZcT5tVwEzmMVbMvO/wCcY9wz
a3tDpeyQpO+CN37ep2mceIfZpWotBkvCzP5uOZ5rpb6Bf719zPRDJmshQ2s5fcjq0OT2QVYktRSs
nF2j7CdbYFgisIA4K0rw81ahCZO4FUBVEHIPP60YEm+W2x12wmjGf3ZfF93rvkRV8roDNTIHIW28
1Zs9JrEkUBA4W6f7FiMez7nSW/iHw7iVlazavS7Xy7xFnKG9PfS/eP2bics2iVLskQxVWyjyeGCs
p/Le0mXXp/nvue1nEv9R52vXGxGj1/ggL0sJ4Fn2Bdqv9RkmQqVVwGBH5T6fi1ONWQlOWb7Q2LKg
qBp0zrz2wRTK7aUclXMUPV/FOcYGWA371ZnhFWh/b76+Uc48y5Jt/bufunPwzjCO4EZAgkSZiPos
/WgcwuNoHZE5OiIYBbRUihdwXoS5dueRkVKpkKLOTVHeWFx7NicPjMFBigX2JV94L91vuJeOM9Mp
4We6SXDPOuMPgkpsAnz8Zh+8XzWDuzrwg5TMwTG0/TrpnzIThhdbtgSZJC3w1ZPOLwKfzm6i2snc
FY8zrLmp3K+2yKanJecZow+vakcqdGPlXOL4iK564CLNGGVTPuufPN0ZEHdUgNsd/SHMHJIX2gMl
+AGO6SKA16CIht/vAgAdH/6TtvK+B7rfeLCdXy+TgfpNp/Oj+ZwR+zoQJv9P3uzwdl2rjaEr7w2o
5t1rT266pVF7NrnF8TocaYIqQPFxuQ+9oSVyUa/CcMMddAG00/o0d5smsgtaxcgtcpQgDkQOEJIP
IbKIycvKmJjyKKJnWXt2dPH6H++KRNx0hRkndi0XLaqhmwrhS4tX7TH6B1cEfb50BfgqFWMKQRqD
qSH8iQpX77klmR5WVha+rzreUNbj8EnkuCKzWTt9vRk87wXbZ5cNx8Yo3sUnBa5lIguH11CPtO0Y
TZgcXyS89QqF9MCDM34VTW6HZ6pbRUydy4AFt4/R7ogHnY1bkoyMAqrgSEMUmHtgytDP//mcqZ+5
9j2fn0yxdtBnE9EucmbYj8FP2Fb7yTtuPUK0+Y7W/HsWAHWYbVehaWro/bbxTVVqNKkrPQya7ms0
g2SZ6ILi+ZmlLcinUSMsZ7eO9vQoBffYcdVfZcFkKpV0OcdtMTBT3o8aoZ4gpTOvJBBAxTCLSHs/
0G4oMIzP5ICj8PYR5cE4/wgbLhSCylnBatn4P134q0XQ6mgIVx/VVWhw4RQLNTfh/CULBUA53+F1
/VFVN9cGytO20ZiUFR+c2SgsOyq3A/XbiwZlDnGxaPyUMjzldLIzNvRUscrrGOfTvATzBBnFKL1J
oulwR+zyi7cy26NIpMPAQCKTbJ+zkhhZdwU2Me0WW1Pjg5We5LNAKZ55XhtYjisMhvPRp3oDfeQL
ruCBAxjxoxsip2KNhFevaqaHcye9URInyhq1dAP76TVgJCW2sDkQc/2cyrEsjuCsaKSlN0+m6TA+
iFnDergURsdwWQwku55126XoASNI9OxaiB4VBOmjbyrsVXOXV0H9Q3c2JMy74PJ1me8C/H7jLxIR
1OTpy7yJmdRzqDyQnXpluDky7FF1HgwNu8y9cxgH/w2tHDR7cuRyDdp1tFYj/fJqjwRvDLXefQB9
VdfyNeOIlYkJGl8M9EFPZEq/75NOnvxjJ0aE2LXXT95wmq9cQW7q33ujOk1rTjvCfRGqc/vtdIbM
uHZU3+EtIIdNZ/cfwAf9kvxLh081E9rhR76icbv43ewnN2QK430vOSvbX9Mcs09mo9uT10J+sUqq
Gi00QFk+AoUU1smWMFJ3Ei3A0lYaYxTGbQ4bg0HqMzE+w26/dAAIjSZrs2574ckz8SNcOjvkpzFo
5/KbtqHwvoL6jRHPs4dDRUICCu5C7OoFumBMWu2Ao1DaZqsiu5fFcaLJCexMXhEWbfwZKGFyPUKw
+P0jW+O/EcZUBEJI7yFP1oVTXHVy6xZUi+B9Pq3UUskLM0KDpl9AoIYp2K/Sp7Yyu+1OsugKcdd1
x5wiHFjpVWUhd/ArLUPfDG76E2tigGK+ONOhZG1HJO/RJg4fRoU3dEnjRhXdJdtT4G7D+gRoS0qS
6/+GhcbBO74WYfoT68Fg/UYjPPhHEi8ky4MWymNiUj2FVj64PB3ZgIzdqXU5VdCvQ7UlBKWMj/ls
7WWprlTbjLMXeN7dChIdWfXjoi47q8pG8y20b6w7m2RWQR7PoFEogXZkqaBa7iHxWHKc6Pb48Ax2
N5wBz8tVunF9k1gqdi+/6ucIe4XOEgCvF++ooH0h46F59nCiOdyUf/JIwaMWR9jl1lWpE5YGV2Si
K3AfxI6UFbB7RXBdHMtTO89ddp3hsECaCmslC6pyAKTnKMit/Fhg8eubJ5k+/Zy8qgJf26zGj+Yb
knMFYRECf1xGRbIiKpvuDkPpNhRBA5KIWmKBULyXzOIWkPl3OdmGBNO+d9LWlJHfR1VHwE3ok9+C
kTqAvZCzkVUW8yu+u9rWp5HQwRU4fWHjezF3tOffkbGnHiM+fkQra+viav00h8Ty6y/j+cjN8Fbk
uY/dF3s+/R9SN8gQ+ZJUoNE6jggmWbTMhdSZP+eN1pYu40G0NEuAjDY9Z7xAJEoVtXhlLt8N/WAu
Fpj7+GlxeUaERCJFFYrN3P3Ra/xy0pDuPixrTcCJWNZ870oLR1mqfc6jHAKvxHcrkgVKciXCRk8N
Zs8BNXFTSVrHl1hMk/B2I0rM6mbGMzjzovqYoP3U6LIBrCoEaa37dsO7bBWZyODOmPFYKg1YU+RI
39BTQ6DO7x4cK0DRSf17QUIpO+54s4FoYyeSNwWy9JyDd9gwX9x6SfAEAnlfuE0kuoPU4gfUdQcP
z8g9ODwhX2mt2SL2u6wr3kw994K/mQvLpg/DODfDTvwcAx/CHCUb3Drh8Eg0DmZPwRLXewTzp+qZ
PkNQf1c5qdyN284Mi0/CovrapYLiR1YTZ2bA+9GdKUp5CTNVZUeWXgwBsLI5ya5ufSowa3S0Ddzb
FxYN06m+/mv7jpMAphZGbKJFGu4jCIRu88zHgGLO7Ks8gn9LSXUSfAfMIuS5v77blqg4LTOYB3Ei
5kd/LdDv5kRMrI2pHmgbTcoKTnMRqDBCShHTQ+yJgi2DxE7a2Shqk1+2xmZh4fqLHbN1fRT/aXnJ
T36B+7PapPh2BVr6g+XhQMS3uE91Ol3oLFtUZtEfYZeoODnetb2zqujhXU+9frNopOjzyCFkD7sV
13qf+JIrbctW/jFJAFk2b8nsOZ5dmNC2vQCzIjAVmX2XLtFLJ6EjrtOfVe5ftTtDTSZlXlj6/dXr
v/LlWT8dVSxz5QlzbtaCXpsd5ER1YgzMGx37WMuKh9oioDGfpqQkhAy5xzOjdnJeCbSLCpkU+0C6
hTyWHAwczgI/AYGdaTazZSxG7SYoQ7FI8oV/IBDQbyRMgq0IzAzas/jjP9uStfjCbRFd0ZSxZR09
k2IdKO18IEhSfSV5RhaVFS49HcrSfDJAQ1NYBKURTnQmfM2R+DuNTsJSernD97+cPVnUG/R0kIll
mOU0izMpuqN6m63AsIiOwZuCYRdiKOXDhq1hP5Cl0dhefDvIdaupJVPxvFFs/9xGH64lgrjUhCHj
8U/C0KHC5wba/9PAqIYwtxDZO/wiWyRHI1YRGLj/Chhr91q9pPPeYQKCTUUkjw6pAnN5RmogagnR
kiQubwdS9O3vg5/Cek9o5H0ihcNL0f5j9S3gY88gK4ravTPCWpkbjKXxLv2Y0OM2yKHdb0x0C/8S
iXTBjbWVXD4oihzEtUh4ygkI1bckuK9J9/pyfJkj4Uzn1lJ3RTn0rWu7cTUmZ3IpKtjZBeXB0v0M
Wubbt6UdBw4fXrlxgjkNJl1p9OoRuUiqZVOGk0Y5MAXe6wIWPd5XAELMDo4HoAaAfPZcgA3aoS16
6+RvQ9DewSgTL2ScslSd1dUhbLA6ATVWMMpSUrX9WvTh+ZR4176ibLUxoYMbjHsPgSPJxqiwGf83
6S8KF7KUp1q6ilXFUZl3EO9VtG1oqbA9/DH2Wd0ZUNGAqc+l5i8qRvb86trhM2EZV/ylWAe2CEzZ
IMh2HgTvnWj2rw7u3lW48gfBrMe2ePVsxod0KY6pWdBHHL0b/kSP8/2S1iFXonl11BPhGm96sRg2
DM6j+311H7Jvtx+GwdFZ+ez+nchmLpj90x/sl4p/QPZU5MNXPLnNyL7BxI4Gom5fsASoJXYXWgFz
Sv31da9XI1Hp7PywHMNNEK0aHXd8v+yRUq9TwHOtqs62Rfoid0rBRt62k9B5oi0MNPTzCNJHKlXT
SRpdISKRpcAFFersZnC8o2X4jrwu4H4aShuA1BBFuT4CKqWUSnBb6f52WjAFuiambxrhzyNaAUEB
7jGq4PL7YAJsAjhm1ymdXJvD1ItxhBCY4pXZCI9Ko3efKnLT+TjmIgB2beAMY3zCD84OOVfBU2AS
BAirv309DYs8zmEYMrSPWr8v4UVvHp/dOQytA0fw33kPIEeYM/9Am3qTqAtRe7DPamd4VIGSnai6
C4uQ2zIPvyGt/JXt0T7AAlocP5glhUxEsw3ao1snCNQeHgLcJKhYQ0WD6d0WcRfE4UATYUOlKwVY
aBejYKU595ZHmGlmybxUHHD+mVAzYq/KyWgHk4pdlXzFQq6s+rCFqM4rWCM3AlSpGa1xy25F8DwS
OtncoeeFTj9RZvwhBar8nAdxawOPcqLEjOwZg3VWvEof9enZ9QhU4nyqltomjSOq8jl55e/BPSWv
Igm8GWGfscN6axCOzIWDrNPv5oC1LibnrLpgFblSu7sZjHwPRUVxFzooIil0IUUylCUI7AlKUe7b
Zw17L7xYeMF+Au8U+FtMG5UKPv8tK3h+vI8roEAAPieCEVvZvl8i0rRwDu/qxotEdVeoqq6QwPQL
TONBc6wsoTA5yYvS89FcFYXB2xQ+3kVwv6wNbl/20z27L47u83Ecqmk3MSHqPzWZOZeg5Nq7KTRk
sVGeIj8ZJZFmcBU/zK/7rClsnQPmAvsMpCRY/w7q1Pt2NXCBZv9PABxOj4F027ecBeYZXcViC5FL
a4VKgHfRFNl24Wy9EB7eu1BuSxXTRQJ5CSwmfZsUfj6jA2QVdqqfGFYtMFI4KlXVJ6GA/b1jWLNH
z7XD2P4EExk81Y0McyOogGyEsfYgwahstioqti39aNVO1VmSFYw9g0PooeV1CA6kWLOOVaYqoIhY
Kg2LU90LzxdN/ytoMiQp7Wm3CrRWDwh3I6DSZ4pdoUnhN5zpaIr6c5CFUzM5COk/rFY0SBqxjuUa
E/t6q9Va7ZQcHBdiSRTym7Wex1RkW1LFvTBYYLawEqENNYE7fiqQI0mOCNiq2QAxU+9gv0BsevuG
or1WKU28jt6gVQv2UebEKBmVoETWpe5Ll8RG7LHPTScnpN4Jd0+Tn7d0ZmBBfiPbJ9rQLzoYhLqL
TMj2C5WDYcNV8X8p6XcXbkeop+Nay2H+ITfBHyBfKfSUdXGbh/shgpEtzZF9y1a58zq0Y52u5Vy7
n32o89wlSa3rQ7Wn3ElamrcEOzVTZt4mFlzxnqek4NEYIgGUjBpdIvsbi7DAju/UPQntsRDObeA3
cY7+Qdf/tRGMXXWLK7HdGdsGahvsx6CKOuooyheBQOduVnPDb/KNO/x/CVXzGZg3v2+hdoKaKUTt
YKfmHaG29gBwLc+Z9NV7zZe7CV4bHuNmxkAnHi6YJZ07ku2ATAxIx+GBgkes+pUtIgC5Y8AigWy5
a9Bjkw2ESUV6dmtSRweLgxY9qc1HZBXaRz3/jKeqzDguNpQE0Pa3cbxhyMjwyUyj4ci0qQ9XJTZO
OzPw54//tSGo4JGnEzhDObkBQPUWvB0IeCCwhLQRRWaOtxPUb/wn3UFzYMl2Va5xd5hADP7IQbsL
cIXzDPKwzqEuYoMg63RYGfmRxDlnAU0yCos7oVvasDSa0HPar9damm7FYj1R017JodLrlzcdNVst
1csFuGJNMPeVthHegbarezx9CEpDMlDgqOHaDcaIrgTTb3ZfZ/ytMq9+3M+PIJoock+xpy94RpA8
hxMvBJ0/lLHtrGva4PiwPxDMlP/A0m5RyfCkEd+404vVJ9pxwvdm7hPO1a6lHF5Ues+8zrzNbS1I
Pt74oYWebvttiq5o7sEcNm/PEOdjBAwoIX7de8btHB6QHoew6IMXQeApaO+obPciQVLydbi4lXUE
Oaj8bDvX9QKXUkB8c0ecVdoJYwm9UoEbN0JwBYSRwf/EvE9LAWMr2VRtkeA3lr5xWcZ0KXdPu3Ff
JlUXRZRrA4tcebHFYfrXJiCyK6tjzZFtM5QmAuJjwCFdx+/2+4DfSlspLkLddMFFp07W4MEzTr0C
mx/b9y3Z3vkMIAVG9e/B3Pfa52pNwYh4fNcEO2CVR8KpYMseavMdNOW75lIaPIO/5imRKbA5FOav
byzFD+qGLLpvc1xP3Nn2xuRBBzsybaJ5Y5OksErFkmCQDjOmreWQ+O14zpFRj/4/z8u2XdtWWlHb
+YwCZC17S+Jc9WgKJYxWEqSpr1lYya7EBLP/flTBSxeyXL6cKbSNlGiuI+/n4RHkPRSXNlFv1zlP
E9htQzrYNXTBPlhZ1aryW/qEwvWDi9Aet40jroAtIAQEtwbcFoWntoAKBv50bmLELs5V/UX/6+fi
2KRZJW9QlwBiljDVVENd/cwwH6vyufivb5+mLDnv4iYh5qTU8rZYE0UB4e0MBdUfTUxOqynHZu8Q
zpjk4R4o7qr2tTOubqnIS1dnmNMIFxQmzm+F4oJU+e9DC6v/5CWBmjDjg8pxh56TU0KFttxQ3MMF
3MNT3xPdPuDxm7K1hLEXXz2W4rhkDawZYWezxTl5awnvbNfb26W0ACjQfm37iyeCrg7OLD5T9Xya
9JR7JhEvDN1irNgvpZygj+vpz7MYZeX8q2FHIWLNVZ51176yhzVaofZqyFaJueHXzpCjNUGzh/KM
4QXFGTp4ITG49rkRLwNg/BajQm4jH3eGyE2mYnXrKPYUyF7XYq5zep6shk2jOFrGCySGb7zLx1Jh
5f143fGpzYyTTGFqylRmweuthf6GAV5iFuD+3ur7ZYPmF5KXaZ0XpgflRDAFTFb5bUiFkj8DIeUR
3ev3OeJzMi1gAKigf5zjOXq1KB/vp5Xb6vTvKBjliNJe3jRVmwT9MSNeD1pNjqweCUSC6hctkkmW
89G2cRqjDay/2d2iaQqBsjveZaMny33NI21Bm2xMK6AIwoqMG9kJLjnVfffxi96rwYiXHP9Avgcb
buMZFIyDnqv/BLpkXkHSKQQ/7G3Dz4n3/5fWV5YjRuvC4YCjcQfT4H+GEgHXB0t9ceVuJqS+zT/c
DaHOnE8TBXxq1RFB6lgV19CJnlnBFSNLTeWC+6F83kN4l4INj2lrjQQCLwvlQ4h58VJsmcSa94k5
YnD5m0LZOostNoW5uonuW2bS6IpChbr6Car8m2Vy6Z+RDvFp9j940J/c/wW+72rhXBAyzDVGRCm3
58YfIYXR4+mMy7RfCyG8dOxdkTd9+2PRpMKjqbKyLosfy/3bdJpYcEeJwKtQ1hBaf5CZY5h5F3Nw
FKaXpkf9/qCGpsd6MV9Ct9oxkKbKOXRvwkTVBwUJvK7qlnuCfIPiq/llJYLyGkxiI5zRdRDkr7US
Gb1pK0+REZgycVA+Z+PNCCRw5GEyGSmFkAjXKF0bSfkPmSq3WghAX01BBF7qSPp1imvTk3s+vNjy
g5E11SX6eY/zbgautocHyUwF71BlVnhbHJAxVVa4bD999WwaKHJaPJ/P2UKkFSufX49KMVTEETm/
yphR6rsYD6mEfRd3tzaP4A3kJwAkASOLxenBPokRB2vWbW6S6e3/1A5pTrfJRpqrXRlXK7pnzwlh
sCdFTZ/AoiIbfKVLl2B4W7znefcuWaqS0KO+XrsvkkyfC4pQnuJrCmB5Qf328u7mRr8xtS2LgqmH
hTJBR8j8Esmh1cG72DnDufeNmkMViaDBuhKtxdzgvAMRqGEt00OTQILPLM1BGbIiqD+wjHczer+6
NfaXO9blVQDCrlbhbOhG2cHlGtnS+2+9Oi+t5OgFSKPo+39CbGeitu5lzXDG+7Ea1MTE1BHYAF4c
Q3RmST4GJNb78S2pnhYBVU8yp4hkfRPl9z1b2ecDI7zztNeBRTChDJa5MAo+2JvvxPhDhBgzX+Ah
JUeukSC1tZpBm8Xa4UMcDEeOPlSV8GptoWhmOY5xR7zkMnboqmV9vFldzRlS2JvIBmY8rEkw4XI7
CouhCOG/VdHVDToCn9JvTzBk8octbg3UTzACdmb4u4/s6FpJCAYe1q46FDyV+lm3kskbMOwdHq4m
aK77DjHeSavug2HFdEFzWaajulWt4lVbZmaLzS/WnlJcUP53hOrhIlJsHEO/kXx5a0OPgboTgVCm
UyV9283UKx/EtYtTOI/3Dw4C0WzDibwoxy5UlnIzxaBzFscmqd7YAWrtZzMkuD89j3+9cZ8pseGN
qlkg1caT1aVRTIVdvuXk6gzcvpLPVwejZtsevsJKFOcs/Cj4hiD4j9R3DGCvzjjBENtN4G14Iqeh
jnpY/Z3aZzlBDsngyLiqXuDpoe0IJd+mUDdPStHLcOvsBDysNYwSJuR7VoDsIVckYmD68e/suqie
hTJbyORq2dbGk/FcLfLZfQwCEoIw9ELLX8x5phnZBUh/vIZYD/k6j13wQG/KHV2KGacLjXlBtxA6
j95ytGkhkLGRpWJKdWZHTVn+peogB0qvf1fUpLuazap3NQEP+CDOuYoaQKl5/LQq69bnt6mn2Uko
ELy1W9gkdkQxjak1IUtzVfYl8W2NtK2nBS8NZdvd83Y7v1cA3EbcHzpgRx0nxs7V1Tf9NOO0ymfc
vt9DLXhVscA7ioB4H7PwKuhLukUils02D+NQo+NebSkvEP2c06iV2hs4CE3161hj9HjR+ZgGnbNw
h4XZd7LiDP5WV//wxBEJxE2sN5mYQBSJJ/gsJsV2yRJxJtifWLwXfttGiY5wpgy6a/AvLIh+gGzi
487Iy81AZwg1L+qAR9u1B/KHEhrqvWWPIxkjS1TzL8XOYl29lhGbsM/nS54K0ZXGsHaCqmTT3/l8
ymaInSYZNsQgzns2g47sVXu0ylCFnXzTxloUwob+/oKCIZSAPeRcXBq6w8XEFH7Re9AIveNUfFQu
HTAwcgkcHvFvA7JtkIlEy5bVRyloT7L9IdWXpRPu9jvpxdwUmjw9pLGhewap+b1K8cPdk6H90P0a
yOin1mXfjstwcVoDvsFzY8pWXVSEa19KZIpf0kfF17KqukDbucg79cpzhoUdgzdMo251oXXHP545
aPzN7dw5WtILQF8pyYQPOXVWUFjxecXJ74mxEu1oBS0AhZurjkaQis+HZgHBIazsm5+fxjru1Z4I
sXV4+CbBYSk2rYYueJVZfxx8h2egIfI7PMxQxEaXBV1L0H31IhnmWTyX9WioU9OF55/OStl6tABe
vqDSN3uLbaSug8acYW+JMYO+n9RI93oQTrUqJ5QAYCy71p+tdIz0vI5icu5wXRpuJHlTNbZOXWyh
bTgUr1hEnss6V30o5zwwjTOFxgcXJWdlossPBI9+VSwkEftJZrz8XhxidHILAoSm9udMc7OepZ0+
P/Zj1kpjDBRXbDPagBrnCRoYUKhmMT4nyyQHIigxVakDSGCv3bxh53zbdxCdZ3vNElpYMb5Qevfx
7o94DnpKIGeaPyMT2Ixn3ujxrW4IQ5F8MfO2wYSjmZsk1HJJBX5fGak1dUVt8MFuO547r8cZ2GTC
RKKBTVYIeEnjfqOk9HhB94uAf8w2cKkBKW6x7QSFFBJ1GvxeXMuAX9A9SXbGAy8aJOAxdf/EXssK
kekeSc3wKKm6td8OdOjyEcXUlZeHStTu86g8MX6r51rR1TdCYTBl59gjAaIT5ReJ+W5TXxUAb1qd
c3uoNWjS1mU8WjJsNbytJq435LHG3DtPAgyxiyy+HEphtlSkopnNxCgmCHr9veBXRmgxXwqLbLzF
Wh7EY7ioeaWsZN5Gpa/cPLy0RACcErJN/L+a0TQkiUcZm3gMImQlrYdXJngXCnlkqqjC0w+dZ8gZ
XlpJ257toXkgMBbsssF64MzEZOLkvOjkBtBqJlN/lAbW2/bpwqe9KoBp1tPifZFN9XRMBkcrxeNY
dKQtXM+knOAtAyMsQSCjEam8XmCU5wPPEZVJ0f9d6VZjFAHoJape7uj7ezkvVtv6pYc3GTG2CHcl
Q5eSIREghsk3t856SAEGSC2zkHOO6f3cybXQjYCWaQMCwoKf+V/wm/JdEU0lvpIJsXmu7GpiTyXi
dLef8Fct+xW8ob7c/HmUCOhEUDX/tnq3iQ+GMtJqXPf0d4KMtm7MazaHkZeu0J+gaNu1QN5LudFU
T0WfJ4U3Mtttd8rkaDGzLNZF1sB+AtoOA87BZElXDPXVcUBiCOp7XrKPP0TPmMZCE7eQcwm3TRf3
hHedztzR+Zmgm2T7xoKI7ZVH2hhHTPqeIbd8B8T2rmIVzb2l+DnJs34fcdG/M3W95zfNafehJXjF
EtgRdwTStnyz2YPaoPAfSqKjlUak8cqX4kdp1DlIuH0bJYqumb8+fk6z97HKsYKH0hfu+JEoT1Mt
bvMpYDLvCNPsKsyZ5rZfWGEpdxUWLNOkMIWoIhI/UycAAz3nWEPLnM5LHekCHu45WfdufDWUTcXx
yWB3B5Ggn9nXQLObpRD79jKtwWxTz2aDf6yTtHcTz2OU8yjAyUKgJ3ejS76HV8jEQQs/yRUY7xkF
dQIAnSxvXy9ClXxgwq5t1/rveAso5P/XCtngqxY54+SGE1fO4R1VkWEfu88RY8ZOWSAzNnxABbKu
wcka/NZdtfhSx4LRt8OQLxgoZt1qRNylX8P8aOu+BxMqKWwK6F804C41RBDpbAgwHX0G/EWiEGcx
GhqHJ2WpXPLkePfpDNwJFAu1Ph7jJrkg9+lXa1kQedeLK+qpiy66sgk6hbHHbwGIRKEE13PqYQLx
FL8ENIpdI7wLa4p5anStGTXW/ilZCzGWNL9g/a5huE7OlMSfbddaNWuVrW2jyx2Q747ciuFBQ+T6
VPv3wcFIKQL1Bu3wzqbCykCAbvxTTC2ePuIT/P6EwF+9e/sloju1Y0aIWlG8bvFSqxqQtX5FTCU1
2xfZLycOP7icF1h88ZH3k/PYY7/DgTKzv54yevn/I0E2glFABxNRdOue10Szp+n+SDVPybXXDSiY
JWCeakV7+IhkhNmV83wmrxkknc3UvG9cCpHjyHx1ukOxw3w/Jkt6HB9Q7AmKAlDQwsD2CMn9b/Z2
QcqajE9FAbqwlIEk53xUL1C1ITm93UpfQ8GJkB7fdKjXWQc2pTwtUeyKGUuHD4K9v+2ZQTCP4Z6C
5y+Grv6oBNZHZnFEqxzCiktA4odmhOir0NtRYg47jK21GbpS6gE5gnbJWSt0bG+pZE9g0onYe75s
dp6MhuQJZfB/DG8ouDJKRJyk1EgZdY6hNea7N7xLoSpzQ4XWPhNOGFaPHYVgIwJeX9Pg2kiicCwi
1c1jrvNdAgXJ6m06z/4vcHfdVi6zyBKiuokvM8gF65CQJ6QDT2jXjsOAogSAXN36f3U/Q7Tmjm/+
p0dQbZrPnnyrznzmO5dnuOcuhfJgb8e6GnStW0jks5VFTrlOQlKSN78AQQUVkL58mw+KM2j8byrA
rG4DrSkxuXdCz3PBWStNNa5XZFmk9lHxLvfD4TN/6e+SRF5bpIGZnUPQyAThOenoN/QbdZy55G+8
QGhBQMQDQDVlru6xm5joKTJET2NXDVlaoJ95hzD8dbfF+Fm5X6DaNoPb4BAZIPZKYPoVDNPEzl1s
fnWhxhXZ1m3TQm1vZjeN8xIXEnkeAfoS0JqvSYUVG+zyjRnTt+jPTLsD+Oy1DMcwlLrguC7ZvPO5
gWe+5PLKzzTLAVbpY8wwkK1Mq41KL0WasFe7kbCVFcU7uEnvaiS58UUm22m00J17bnftPOaO67MP
KjXgwpozjsIyxCwApuxjediDi0cVrVyDCBW4ASjZdLQx0Us6/NV2UNZMUWEIOuLn086PBTti2hj+
9dQNCsLNYDI0+qt2tabQSQwqe4P7VoW/6fqXOgvwC+FVz7xgj9PH4xiASUG3JMef7EjilJ/5hZCp
fv3wHgcfMe+HLj+P/cfnYkWfJkQxK+YcXyA7mHcBzsUrNlhfRV+yIK/gzORw9yJ9vu9RYCSfBSrS
phkv5v+DLaI41ytvaXqmXG0RDkupERuqNDqcyHVqhVbVw81Sc/FfDEr0cC16K3toI2uEEqgQgrEJ
fLr+S/uWZTO4QJwxvPPoVY8uxbl8jyAxdY4xlolsW0E2dKe/OTSqSh04zVCIOMghZvL3/mBeseQT
h7QFf0ljMgehFWrqf7wlM/25881hj0kgr+jtz1YT8+v/FOTkLnZz61I6q/uo8qHGC8pbqboXaurr
SA9J4DZHQY+Wc4nV3Hqomz+axvHf3DgueL7tOd3Vcw/08XRSkCtsj3CWuAGOpF9mPm3/3c6w4i71
i3dsmfl0pXpikM1yO4qgdzxTcTFldIS8rz/MtVxLUvZv3zTCfrYankF/1nbJrpDZCizGjrACtjpA
P/5vxX57/Vc/UghMeanJrJpquheC6IxH3mFGxQ8+rmIgcBFOcvPPK+W5lYYom6TwGbPScxvEarTY
ZzySvK/t4Ln1FOp6JIw7MTcHmsN4CwOkqhsylMK5sHpKK1omeRjBKnwRxlVSI4ekry7TlkS1AYs4
F++8pHVTUd+BcNR2hPtH7REDKAP8L9aQwUgXITuPuEjwIBjGLEDDg3KIXz/96tb71Y8yQZ2Vie2B
+UtiaAPdkJ/qx6b87ojQ76u9ELubo6EKOQPwY6XtWC8H1D4KRhoPPKdWpO6g6g6XglETHO6cI1Jh
uaoJiHBDvG5XKKNv4fFcIXThG5q1Q30E/j8BJMu4AeHqmuhFsNt1BSM3pwPHkim8A8815ITQiLSF
Ihw/yTK/NBGIMlApcNvig5INCrKJmROcdRrV23y5qm+vWLjwREzJTslEif+Ke1ROv8vvjpzi5Y/u
iO8+fVLawVoVz79Om+dNI341Nt6z580ByAAsCnxso0ykoMsVuYW/IRCpoN8BNI7560D834J7DwBt
2LYmOZC1cve4ebclIGadKBLWYPVFXSCvQIePeH9OJ2gHpKWosZz05Hw0oqFThrxBVg/5A6vxctpQ
5VPsLsLJpStOh4qo4aRO1U0EywnoypBKyFgq5nnsTfvLVXJIHyFdQmIKp84hnEUjDeenHdmWM4J6
1QxuwrQ0xQb7fHn7HhnVq7KsCOKkBjzP123rHCjsvzcEMzvJSOVKwvqNhTyxbgzPJBdnlOpkT5Za
vT4rqV6kHafYJQx0hMZGOKJ6w1tIp4BFJ+MVnb0YpgMpwJFU2UuGDFBxfNeBVUDf20wJO5NRKmZj
yiuBY3i6vC9vAFISvE+k2GoozmTGf7YnIbCGXJNHqEJgVm82KENLJTHhF7Vdtt3b+JCrr2qWW5WK
6W2qTpUxVoUKyMaZn4MS8uFogXS8n5N+mMPMOrbS90U+dXmt1wJv49bo8kpGmlZALwVeUNZNgAOl
HHc7euUq+/lHtYkpzvbmH+m6kscRRsQCgOF5hjVuSyw1IwYjnIeNhXwWYWW97FbN4SXYkGlhTUAz
31i6+5n7tLs1nP2njZDdyVPJPN2cGcVQH7kTuKGZZl9pfCS3cBhsfCVZbAl+MCsYdVc8x4cd/nbI
PwVclD3oHhqWKHktOhHV2z4sGqPMI2NrQAtlPvFnt4voggJdoJs1/5JsBVLqNgoTjZPfA6DbnCZk
doW0s8GVyPAUaJdzS1X85mE6BsQUp3FJGzjtMbV2+oWP99lhLZlzig6O+d4H+tcQte5Msx3Alw1R
zkLsrw5bnxfS/if9U3DLRdCuiFZMVwZsNx9qS4seduF82wg4KTp1mxS2HWqskIEmA2Gaybr8wFRx
JbTSS3OZa8MNxJkqLTTckGwDY+lXvRwwbRDPbtJr6qBxTJkbkXSYWLb4q66zhNCmGMhQsIzpBMnj
sOyMR10FXoiNlKTuUwN0zjNexWOrc+jDJHhQF3qseeuPqruw9tTLqOgJiy1myHs3kaVjUIuuUeRa
XnTeavYEU76v86XTMCT5X+/SDdcVlF9Bld6pkqW5PTgpfUTnupWt+5NCE0Dnp/cOkZkH/9XdXNHz
DZPIuaOceQrUaAT45YkGnQ5jJGwKx/6Ss5axQQVh4G1x/UebUR9TyWschd86R7dMP5QkhDsrJA2r
O86o7uODkBDE/XRraOjUcl5BWu7g2A6n9WTkq8XTvtMInu/W3PPEejpZo+3heqTVgkD1VMYMg4Fq
ow+MO3GKjsPKF6SJ6OIYefehqWE4cjAjFwGc7ld5lnlnhkL+2msPJ/63oO1aRI5d+jgimnm7/TFx
MUFJDYqdqcyEJevDI3rU2GFDvVa+0hToPa0kqcvEZ0sQi6BNMMJ8OueBY75H6patB+UCRL3Xyxda
HG5LN9nwm9X++ClbSrMUxkMIDE9U+oaLK0WcsTPGeA9h2jf2CTcLXpo/312GXLHJYtWOLMGXH5dm
twLqcFyHdnEQ0LJqr+cml7Udk1Hesq6BvwTXFnp/nLAS2m7TDImHnLh2qphG4eNj2H7yQ1CDz62M
ILRb0/bWoEkOgH1RRmdwdHwxJZ4gX3VDM94wxJijxg9OBx7InOAwCTca7gy/n5pikWg12J18qaQE
NxG4PrS1lJ/3BXuD8iER2OPJwyHNphOaF2KBXmyzOH58VIiRQahgwsHsZB3DvlsJZX7qC8LHD8EP
siVRWEU+M6RMF5lZDR3fgwOpLPTMt6Mg4dACiHt+KRSC+iczbIdSfBbO2ebb/buOBFxeco7Kn9gh
keJSJkG+23mZUiu+ZqQS4bEn4XARWMcwGEFWG77+EBGiD8kfbqtQYIF3PzCm05CeMyk/SqWo/Oey
/SXbnQ92xmNus5hdB984j9ILT3vVE3hEeCdi1DQHdrvN09FeE0yiWwP8FXq6tnw2CLs7MREoiQVT
aADtfhdu209yKYlGGBo53gTMBJXiiQsSzgVRH7idi4rw49UevX7YvkhHdw6MVzheHsLK49hOp91O
vb8aQnjZI4xkT4UDDqXCpeNUIU5R2CuEy3p4X7j13x/G+dTxQljQpPRwmtxsY6nIb8MVSdZK9K0r
EqXU9Q1rBJcPJTon7gXDH2e9nbKPE+Lla/TNKkx2J8YSnLkojg9VHeBUSOvTY7w4Ow7yWPw9XEYG
GgD6Lu4pJPpO+Sfus1SUO1L6ALgnGkGQi9DNCoZ9qYux8itlANlBd5pGiQINGHUiI9bzUZrw0HsK
DugmLVb+js531yvzkXCgaqnhXk7hNUEWQ4PIIQ+9hWfcz03KN1gUFnWW1TsiBLSs9N6u1Zew642H
qW3xLG6pFrGQMQSwoKap2IV+3bpx45CiPORE6uT/ElfaTFWw63yE6VCwgHrzvKTi7uVtOnd7HqNh
7/IwuW8p9KguNsoZMAMNS76pA9eb3gG9gHw6kPvDnZD7oFA6eYgf3JrshMZRZSWj+NhrCD7Jmf7R
OZouI06BXeb8ZQ7770urUIF9+8XRPSkj/PjEhr0rLeCJX8545nWcucQ40r+mxgQaRPeWm+qh2KwC
9KBFHR0knHDcZSmzejeHott1OkjXhu8pStqPwyl4XrnkxbFoEmsPCBr5iuxB3Rb27OAeInmCYVdi
XAP2Nt1czwHTYv0DQtMyI9CglioD16+MaQn4ry9aOcigrkg5lOEBi+agGoGAc1tWMq4iDZ/Sj5ja
tMnjXLAhyzvdlqNT2d0RfD8oHoFI3sW9sBj80hkOTJ2yKtNozbTmYJpTTX5Xtk/yHxxRsCU/BdmA
XVRcqnLlS5v3MeJPg8V0tjzw+rOeLrYnsDCrG9VvquChdi9zEuN52QP71g/FY3iEhdiYE9SmyWMm
opDTecgyavo//vVohI58zO+DyKaUQR6oT4qFUqYsHjTynqYMf7XziSzK3dTbRI8qxdPuHz8UzTKR
fAjIClW6RUaah0aZZD8XUw3+RrzOBLo/V4Z/Gvo4HzHwxiW+UtJGF/4F6TuCfKC5NyanHxUoxGqA
eWaJrzYgBaabh/akd+hfWlchNe5hoLVqp+LSVNaS9BY11HDeVsf98yE/ulBsZPUs0mIcjXlAJ6+G
CI67elazKlJcJJKSeavZyFRg5rdtkWt6RWLBDAArzWS1kJVKvX0KLuMhiw8GU/aZpsI/u1zhPQ/J
cvv7vL95jC65rtHfOMH0G5LFDrPUNsNq1i7LdJ5vm9SC/9lQD4vGztmIUOZJJTl7y9hBG6HQedCW
unagGBczTkGodPA9uyB6DrHSSlv8B51xi5Mu8DeqBH6i55ynbl4W2DEvPOCXSVzrLHaXacKBulG5
/G3RwphXS4AXNFvSFCi5ispwAHRx6OvydzClLs51tSxMT0gEPhBaZ/vrQWQORkZTqqyEtw+IsaTb
//P3W0h+ud/ulHrMzgh9qfeOKtSg09Q/Uz6aBNgnTmddvkbZD0wKfbRTa2buCdiIokCbyKEPkySx
5jFQ+visyOY7NYhMkYE0AZ6y79omKfbbkY0pu5sdUWLSz67Ir8LcIWBWQk64hKVNCLTP//wIgLCW
+BzZme+HQLwiwB0x3JAIFSfwObiZltmOBLDayN33i2OG8NBrf1PLgBO8M0kYXSggQQ3VfZqUv/dY
p+KG9ywSCEMTkHqa4OgIyj8EZrezkcsXGd2N+zjMq885uPQyEI3pPeKJ5KXkgI6WX1RJCHe2Lneu
9UWwiC963JwfcvCFr+5o0FCRbMaqr7LDjotmKsqdoK+t7zR1CNp8B8X24r07k/QZ/pn86jEHHFrW
jbpKxCdfgtmikpjqE3rWsc59Js/DFr/sMuDOOAWfh0Dmhim+tvbXadEcaa0Wa75zpUvJnkwGxoJL
8idFYOgy7GLIhe24JSuh2QRGJrgozFBDEB2k9ermXEeCnxFY8AtKhly9fu6OZBrLhlkhYQJa1Vi9
21KC/7DTpgsoV2Nfig3pvd5eodG+ms8X709zcW2riLGg4oYCmmS0UnIvWYuz1ruDEQoaAJeD+evm
0fDqPfh/TNku+FqomAOvHU/KdrZyU+HaZr9uv7k+dKD70XWVoof0AFAeM4gvw1WA38VT5bXETJ68
J/S7Xc/cTQZ0TjQyeUxOZaHqbu+bjwSb2Y2oNdxTnVK6p9hLKrYAbigB6bgpz9IL7p53TVXhYnV5
lFuMS/63gzWSDL4dAvZk5xnuqRV+zwIU2hTLleEJIYi9OSGMuOBxqj2ObKMNGul9iMPdXZnppybp
07TnusGWJyh1G5h5iGqod/ZohFTSzCJ/F0aDB/lOMDGvzBj16KneosDW79c0DDGFXaMdPeHYeNm6
EBJw/TtBzWCvdu94vd/FXFBMiSHTeY4V463G7NIgh3Zy6Ij7ODSKO8vo9Wgeu2FVKf5WjavQKzZI
qvPGpXvytSzFohvIEsS2dKxPnOfrUj6Fl6AgiQdyYdhieiHfq6nQTKLpa1NVj5KJNv1Ovnxlo3xy
aiDHtSh/+e0BFdL4P5RHsIPJnYUrbjjBAlsOEa8K5gm2A6hJIvC9X32xomsVm3Z8ovs6Ja/si42d
6ub8MEW5Lr3Je/xU2xnh917XRp0HrnKNL+Ylz4QNoCrueL6SmDFCqOiiwp2Qm8VZwMVtQQv30dus
OD3TnaNFo+EOEFNHtuFrDTQ1IkzPSlzG1XD6+xhVKVt1baw0MtJ/UuhxuYj3JZZOnLxN7IA0+FXS
UNreHjy10h4vBRvDx8B6gxMXc3jusJh+RlTnVh4j1NfQRBnkZ8TRmlE4EQU46aYvFiqP9xbxXAgT
31UoldpmmurHnSCoolJS/7HZlgcflS8nUVtMHQ6LH/UCSqs44+bO28mFfcsKbW6SJnq85Cat/hXC
FrALmZNfsRHJUJEIQB10OKjJTsj7SyshkKLA0k0CLjl+/lG8bPi0NiGeBh7WzhFWavZyAC4rRqRj
Jw+5zcIm/qsk3fKuRKYkMBetCXZk+dFf7rXLErA5E2gBiHoU8lvI2pxd5CkCpo1w5l8c7uTAPWiw
DsmyVjLwpHhSILtbkRcorNS9jjrDHDbkxpHNN4DsXB6ARpdWYTPoqdq5dnbGQbpGecf9C4qilcFp
irkuGJ35YUKKlytdtdOoGgQCTb6+JTJfmiQVTnZKWBnaf9vrCO2HQhIYfp2KvbQdzctIVDe6ultR
valMauziM2F5AnTsPNLoIfgvNkadjqHUyMhKGFJMLnB1ji7ReOqBwJ+Cgq1Vfl3RHFBpiUVMpngT
JeEKMy1uyh/+71AvHMUApAcGPCfuhSyDOWtm4s2H5vk37XghsMUPXvqQXsAbCSx5e4R3axvyBiAv
C9dpapTXnbcDiH65WeVN8/nfobh9l+cxAaKi23jm8ZeW2I/Cc/9swPGOBvTrLBh+qJlU/nFtKtvX
XCRLtrNwt3Ar+e5xgdmNuZqgevhF6FecOawlmvZ6BbNf8P9CspajZv5Htr87JB9p0r/sUYADmNoQ
Epg8sfFhe+lajqJs0dFKn0Uy39OlgQk5vNX3lr+x9WnXAF234UgP2JLpVd5B/X+WmXuz6thPfw/m
xc2Dz84QXCTVgL6XSMuec1rgITuy2lqbTS0v7Dhh8WJafVRoTctXgIrFmoWbS/dLDMSnWDX6kVGW
M0ILdMXrMjeWtW1T6JgRBHx2mNUvVhU/C6M3sWbCSetI/R4u2CC2Ak6sUgjL39UA/yNg5kC/xxwz
w1XMiezXa73xHn47hGzI3q1z2ReOPFFVFLcDuZNUHrgLxXTi7YdD07hdgyb9NG+QLeq8k6YBobAW
MAcOT4V2fumKG+EjCzuSsQXqasKm0ajdBwwnOa7GfAK4ttYlIxnSleT89K2oAqKIkOJdBlntkiYQ
6Osnr6PAuKGq/4EetcLAgU04BzbA04yZjWKShoQDGMOxrqxFAwUojtaSXBMiuUuhhUR7k8x9WHTy
eLR3Mj268My7KxocVf5JPQPwD69+qe7GmDEqd+KiUzyuALR+1jX9Ns9s6qTcFGfo4z0ly6C5pu+O
6wWCeDq9dhgR/iW5FHQ/Hwg3JlRLfT5PdCjICg4cZlQdzb6DpZ36ruvG8HGTD/mjhLjJ/7gcQ2Wo
SEP7+QkIRvGEM3ULw8AY5yw4bNaihQw7HEdtHD2eTm4mKyKiwLKk0N59vDvY2VZGDBxc7aqgKkW4
+tH2qS0FEaXTCimERX551j6QnZpNC/BVPOb5A+i707P2cB1t+updQAxb77yh0+Fqopc9svbqbroL
T4y3hXNayh15G/ynujav5fkrLYjhAXDPaSxFV7Z1UWx/6Ru5UbRV8W+W78t+foRJL4k7NjLFozMF
UEKOyROCAYrMFeMbf9+5VBOXKzxL9zdII9wTsKOWq6bt3UzZDDV36rRi+nITw9lgUNETa3fQ7cIQ
4yE8wxu60hGUzmUwq+TKz2pMRybMa/GKRDFAKtNn+zs1PJToH1v9USRnOPcmvQs2d86DHpAcALPG
t01ZdBL/Jwz6mLVNuoJGTqASeLgkxV2T3YlIbsy5Snybvv3B3dboVo8RSJsSYnVbR/8KNTTqA7AK
RW5OKKqsZwuygTAXMcE1fzEagkI6GhGt5URYxCFsK7jG3QPW7m1Jkc715CGU+cSlfW/+AUzwUS5o
6O4FIfObf6yIy8keUcAsosA9IgaaOg3x1/6BnVXyEaJ3HYLBZVmDPpvSNTIcw5P48DpZmMtNVjLG
IGS2L3yNLCu1/KRAbYjTXlN1F1Ndmzhl02uxYrCMoNxe9FiqZUfyEyhtJww4wi2stjtlbf3e9O/8
+HcU3PwE9NWp6J1gZFmsYxEDPZGwcuPKdZE7YJkwfsPUvJqKwHROaXqH+8w/ZgSVHGusPI3qBSql
DtKoDqIBf2yF3fe+BJ1WFTBAPzyDcDlKFZ3i1XXFIGrsjhpwpGbqkIcFOihSYaLcQvxVKo/mSPFH
3J70TaJcVCr1P0DcxiFlG2hBSxSvd4QobFt2xWZZrHxN9O4CdqMWnv/aYeqmrJgiCF1mu3lf/Kpf
RKoLCnpf7qj/9IY19yWULBS6Q03JSTGu8Fn2Wya13VhBm5v5ypuE7hMrhzYBxx/0hb4iX2fi1wjY
Rb7zUt5iT8YQeyheRQiCftTVjoxPVZgtSjZkBXVLMNogdsQq1eBWpyL1ZxeP3gxpsyne8JQV6AiY
JhusoDZDELprY3P4XfArO6ddVZjfl/ezjDnO9lAoWC99pUmv8h4NGqeoX07hfj8Tx+tp2H4N+6Bs
yy/DTrRYyvOzcGXIws0g9Rb9coHnz4VM9HP1KUvyVH+REjOd/Re6GoIzmR9lxM0+PSJq6B+BR7Us
CB9euB4qjk06N0B8C7F7YBWR+KUhEugluz3B8wiIG+Csq5PMzygT+nNyOsm1bTw6Byzc4LOpazCA
mCoileaFfS6r7FkVM0I3AfR5ker6Ew5p1Xx7HQ4y9gqPIJiKqlWVXWHnLXnO+mOKTPINLUHKrUBE
QeQajSD43Q1W+nad9ZHwLXYBL1h48jEkxOm3Jndf0iua7hSSdkryFJFFG/60iM+ucqpAyk6zx4ni
sUgiizp/F2WiU45nhjYO2wQ20EEn0szqrzb3DnCDUiaTyeEusxV4lPImI/qvj9xKB0pmu37SLoZI
+uaYbeY4SkSiuiKJnn2lFZrwxzzTshSFy1EvKLtrUqTLTgsLKhYsemdBXQNeojn82xrlR89SCgRW
hlDQ2n89rdFsFq1tQWRblM6wx8M6j7Bh0sCWbzzTBcFRxggwm9oZ72KphUZohIXCak0kKJuMZvdB
PxJHXdKwEZjmC6LTg3D2jhDul/RvZionkVBUZ4BdpCudVwt7LSHdOeey4Hgz+SrV6YFEMFuX0EC/
2roU6y0FHMJznlVSHYMNtabfN3oztu/UwwQJVltk/plCJvuuj4A8YzrFmlZNBJS0UXt30b5w71B9
3Ro7RBaYe8VXArK6gBGbscjJA09yeHhQLFxR8JKpv6fL6PZBoU5wmXbJlevEjUfVaaJ0TriD8XnQ
2/UebM+Fc+bsXsrnMZG+iwiy62kShbeV/NkuyHNLMA5chvIFmsOK4RsO14aFvamCMRA6+KEj/Z4c
5LEDpqF5Pk97L6MudU/3kgf8LkxhRjrCq16NJ/Vn+lMuieUGDUImZEI29QWA5ZStXsn8g4vsCtyk
Z7O/a4Y5/vp+f3KTU3BG8I78GQjzlvJ9B9e8hZSLvtBdRVDbOn44gGE/Roe8DER/YmRUg5eENipJ
uiw2iwu4OLSqLANiEjo4nQjnIgokAvTWtq3qtqAujR3hGIn6KHwG1jYm30mvbBrQTVX8gk/F87Xw
YbCQb5O5ze9Yzs2ttmzAwo6OIaXHL7DOTR0jnFvozp3DA2SI0pFZG+JQ1AHkjjoN2ORwAL/Kixla
SdBiyVnSs4IAAieZMYH6u1bAnOJt1aqnncXRx8B5nP83Lrx904ADW40zWkyrP7g4V8ua9HAIwSmK
XETUVQDui/uUW76uWSRpfnPoQETwejgS3yJ4HjfvAuoUsd3gSRaX5YqYI9Oel6u3pIalT2jcniW7
kP9gWfGRaKPx9MM7t99irXyzeVMTtP5R14gDnMVReH8AVPr7g2VcV7hUEZsG3ZaM/aZD3c6hyUDY
nKvW1EMBZ3UxauA3sS10hJt5hQCzeSS2aYbWZZoBQKu0dyaEZYkRimyW42PRL1a+t6ab/pakJiy9
FO88lRjIwwmauJe36/M8P3O1AC9aGJRDz4HoUV1lm9sj3PR+tOfyd1NL9hD5/0I+J9LLTbYjZsVz
plMjRWfsndZ43samebk+13j1ulruISp7wfejfeAUVAjr7XSDAKYewcVVrk+C8eRnmKdo9VYUAg5a
REkF2+S4DfPOo77cPSUAUSupRQZHGV7E7kpf4RRZFbtGXN7/pBXjoVEYXuFRxQqL+1iuTKtI0sJ/
+N8Qr/z5jxnpfJvTe68bpMAyFQgnuogixk5AU4SlS/1JEkjWZeL5IzlwknJGWjQ7+68EIMtdr5Tr
UH1duhw8m8WwGVWrFfEvfyhUN4ToL1kv7ZLsggBNIbeaiXmn/fwdoSL9w00CIbCyWOCVaGOOMKof
I6kE2I42uLu/di7bVoP38Al9qud8F35gz50fE3HFSRQoz3v9QTMa1r0+WlT3TOKmDy+jmvn2vzkK
AmjoYV27KMdy04bzchMRXJNqBGeKnH17GEvFqyqGEuUXFg9lFzgFmFnUAYKascU5f+ftcFSPcNx2
wLRJMIKfiN3hDR5tRy6ct+bU0rXxvsUHwxYKdImU2VS1EMJBwj5pI6xEIGoo64JWiXwhSj8KzxQV
d8GCQ2r2fYDVhaJYp3Hh5e7R96YSwHrxf1M7YjfFPRMxcmZW08Va0SjbX/+/JYF19kgruGpKcdj4
H8AQXk4DppCCIKIMVlYM1XjEVIhjPvbKNngp5wVc6jlWcblL6v72ZPIFn7UVJaxxAfgPjMOK8/PN
5q+dHzm72M42guvI0kB/PNPwYu9XW0agseugVF3UWYyPLnYDt+DXu6EKa8WXentIsxhngMGrwjMc
HHCKJvbiEi2UC3QfvkBGmfsr6A7gNwtKuSSMrmhwYZn9QuGJQXKREzlERzOiZ3oU78WxMohGgkjq
6SNpUy6bVxMCZuukQ7kwrfpgessimsAwqFnoX7OPl/mC4Sf1KLiTHnY7kVMuzbNENH3NbSYtkek6
pzuf4L5MJaIsZYjVS4KZo0vERHJwBOmVQKJgRgqJoWsYYqbJhhkcol83wkVeUeX/iB8gvAh6IrO8
Xb6daj5ijeWoW5zVXQ35rjDDgj6ucKgF26OPjMT9vy0jRcvACIbnoTidT1AhgnYZbPCT2TFLpifK
Qi3+awe33w53lVAyMLIoqZ+LoTfLogMMIHz8IC0XPOFf++iJvJiBDeguHtzNP69fcS7KRkXxPmxI
esaALAKFjhObDswpDeptJ3hb532+Zgfzk/m1MAQjIyIDKfD7eSxiU/9OxkjigNzH7LFhM4i3ybZ9
vokvJQ2N1tdOWQ9/T4X40Qilb5qVd/5hvCCJaDD6UqdX8CYFTDpu4l1BDr8wQ6j84zg2nznX5ji2
Y1r1eXG5QrXUtnucflRQifbpUHebpKplKsGOUVddmArKEqod4eW74vRhMYyORM4YFDJFIxP1V2Ym
KThlq3LKyKrSEeT54saKnaur/q+MVyv9gp/3k8v8A1E0LNZVllnlQvD/KZGLjbeUK6zz7Ntfu1dT
aLa+oh2ImISr9avHQIghyIESE1Od3+flTtLVdZmNyQz4jhNLmitE0zaym9IZEX4aiN0YWvkyzCy4
vw0BtWf7VnuY/IHM3E5RD+TzaCi45XPGe23t2C5nF0Gz4LqvqOtrTfFJOePpypd7mCSCxh6dN0qM
gLwta8GP/pJslrlkPBlTOUSBaay3w5x/vShjamhfTOtvJXzKCT0bv+y6I2rGCA6Uncj4p8pJJdLu
uSlk+0HARPMUfHgNYF+jJZggrdD+4ioo46LeEybtzMxWsY6ua8zgvNb6HacB9pkcgUXqAI6pkdd9
/PdeQYjrE4zVHt6YEyHpXUE2+Hi6Tgh8uJ9wi7hKrrWmv6WJeIWrg3U9KOKpdncTv95sKX3ZmHse
1zkZUYc4ehNoMpu8yI5r1HcmP/c75BCwtBiZEsHAneESWAxUQS8tHuvS6wfRd/mmaM0LbiqIN+LE
Xu37rGTigFhyaB0bublF09afAsvEuVtX8KzQMh5duMwcblgCVo6uAIUllN4JcWvTEdXBLW9LBBsh
jnAnthdwcCgaUJ428DsByGGGdp9QeG9zV4ryR+txXe4Y94Rw2a5lGASy57udsP8Ue7SvcWW9eq2o
IILXI0Pxvexs+dfygkQy5iT6YVPPZmwRd475VGV/0gVQw+wNLDFbzzMO219aZ8d3BZMD5JHSXHh6
Km2fkC03JeNf/Bw7yzBqLRTZfmSLP4WsVFqS2n99NSDiEmZeE6iNF5btrF6CUrVH/IO2fyVpmRze
0DuVjvqbD3JyGV0dfs0n/rafJLl67uEdbB/6cK3AKzV4cUv+SHTBTNFx4Cxw4cLqPkIrB8r9WK13
CRynj2RqxjVdim3KOgxb9tZCyRwA4KiJaKc4rYJmrTJfcSPwqTdhrr7RaSQOSsLoRNc3M4ZErHDo
ERMT0q1aRhKBoILoDzk1JfSsr3mrAF/PkhDX/SJVrUkV04WyGxCTcCp4ufKGcdO3LRm2MBOgiTVI
x6gr0ABcDftdB5GK/qDMmwqjfG0VV81hKJ84sDINd7oS+7gROrJdAaTJlhVdHc/Zu4+apOciOQNf
nnXGC9T14F5EPCYOKEYtpklhcxJeA1LHgs0RWTSM/5/L2s6Az6DpzzOpJcaDGemY6oSae6F9joVs
ZnKvxSzTk9CpusvEHZ2B+evrzxOyyBaObNBciG0q0pmSArP9uuG6oL+qDfOvdc1D9VdbhBSlffM1
Atg4TGu2OL6LeNxehmD1/XnI0MDxlTAV8Qpkyfhc8NJc2w/J6RvLhXGehfMqxLaEg/fwHJHKhfiO
n7ZOrEuZXkO/U0Yzwu/gAJVQTua6i4+JWsq6VAU8wWQ/8yBDma+2QbNwn/N0KHMQtqEuZtrdnxjM
1egoWQVxGD6NhQRtCJCdxXiFZ9YA6GjPEMJbURjpLdrdmhwR/JWxXA+LPp9g5cl53MQq3l242t/7
svGn1+FWWCrnet1bcOmzVbLyIPNCFqhi41xTdjwZ3/MGEEC1pDjojBVLP52VSRrHPUW7lb1yuLGv
8Bt8oMd/azI6dsymh90yriJULQ/i23XXYhbHBGqS41Nv1glFFcRm6DjhyvJL23UT0CHy0BwfpurV
SU/cE2lUs1TB4VzHRrtpk8zgvidHGbgKaK6DwCBOSlSG09R3T/W2jHGcBHPFekhOf+1vh0mrSXQW
xEke0NdsKZRyKA9YgiaOqw8hrZ1SUDN+uVsLGmdAxpZjSn6N7TCmKQ3AWV03D+fcOjvGEBZ7NTQG
yh8zaRNpZulJ0mzDCfz6jgzuKH77OWMXY3NqPirgCb6yW7WhvAscS53+eOt1KZZcHZM+Bthsg+Zp
ny3oARjz2ruNjKsbRYg6aGNWq0LMrDpJ/zoyKxMjpUk90IxqhySP2MLTtjg2npQ8EH5MnWZUh8MX
xeeFGLyrhHmtzhLHEnTXan/DyPxLT3KiaBZNsvM5JvTOCwwx6MC4fsvYc0+MHPLOEGGVfIaI6+R7
8HOrED2qR0pPFVaS4lBXpKPiY/rBGxrKbis1TVg+iOoQLQVCp5K+jrqaiZ2o/6bZKHdsL9tL75/r
xUzYYE6LfmSnoT6amp6t53M2ftPL9l/B4G3MHCmNvpLafrqwbyPIuejGffgeDU9IUDVAYs+ppz9M
S4sY9BMkPldsf1SsrV8gaPsOqW15j/9GBcDu49p+ibMv0VhO2jGpJT2lb5SfwggAziGettt7wxDv
zQ1qAl1gFhYcENMUSpDINBZhnRNrcSFalYPZzIYjq/ayQs8Wk6cbnmKMC1h0aslgB3FUUKaTvnet
6Mi1dP4ukD8yawEZg3nr/nF3vCy3v7sSY1w2FTcDWF+gB09EYLolSx2LRupURjdsqsShgXpjJphA
WDNz5oG8ljhUx8FiynBdh1MfL5A0EOJPDw04k3kBcd5P8jL2/5qwNlcp3sFQKtxTJ1pErNfltxel
ShfxtyZy31XIa/IEQlYDy3zXYMtc37ShVEUO1/hsa+cz+f7xOq57rE7Y780d+T+AnqroRKKrU2ws
8lUnm4qsvDVLFTSmvUK2bu3tVgRlSF4oEarFUrbgmzBGnU0oGNmS3WTi8Y859UNOPVxYzac3PYix
x7qwWgJRMSXat/jvW3kljTujBDhA5sC2AqH6hbWkExmL5y9erFesM9d2ETUOT/W1zgyFrdgOb+8a
iyPvuSI5hJ7mWa7dj7iw+UkqUq1V4fbnXokNOiU9wNtZ8xiGcA1d0zNw8lmM2ty4Rekntcloq31l
5mJXv0x2u9RuEHFTgHGoW2cgGlzrj3iaYz3lj8YR9A/2aEVneF3aWx3oAExq6xmwz2raiLTmHMTr
ERJQFxZMKJs2oX3SYIdszF5MdXfOlUX3kOP3qOGNVywwRj+KjBD5UaABcqZleY1Ui/EGHatOTm3D
ztqj25n4BNAAHz5QCZJks8cJA5JQBOcdv1+J7U+JPWC1J1mKE15lBL1s4M2oHNyiVko/0z1G73dW
zgozQXa1fAdsJZbf4PweFfXQXUP+cvyeUxlqy71vNgZ3N+gjc71hwbxnzefBVoZCOdD6HpZvqbss
IYpm1zi0uYcrJQRl7YWwIYHqzbgoAxjIw1+dfpRjwix1dxOqTjxpC5xkGQElpq5kMgVm5cB4Tgpf
dr22d3/rR2XJcttfslD9iRZkR16ufinM8fUDKEVOjfQ5r6kDvyDiwZuizjfWByGPeFpNu98syC0m
//4ibwuASIiLl1aoV2wh2c2D0XVOBYDawR54AUbIEEh0zo/FxIJON6yq1UFNYrIrkvUjY4DcMd37
ioFddUNmThcsgZGNnon1iWrrY69A8x+9hLSddwbuaLPlwQcQoLEjU+JT4acN3Yn2NxV5DyR9wM+k
VT6+47B22UkzvD1s6Dl3RxLGXGktk1sTqe5/B2uGJdLPKwEJAjcSwDGIYcfyj8aSi6iuM9ov0OOE
kPzPtYXc5E4VbIkU48zwrdDBV6HuU5AUU/zIAs43evd1wXQTpx9KybZAAKvj+b9TIrQmWVIIWhdp
VOnKhle2nMflXlkDTANsZt/oeCUfPo9LxfuENp7uZxrU8oE5QlkyWmvdCuaIe++uyzzEUFcu+66r
6Ri9h3Cxc3S+31kdlaR9ql3l6qMeuPlmj/uJI5ioiMw6DLeKLmwKCOA8UozusCjq7SGLPgQks/LA
yMtM//z1pNLecQhPacGYENjHBYmvav83w0j1wA+3mE0rXfocCBNZ7CFB2dknyb2SLBOurCHvdyfk
AjxaKjOwhRV6pqCusSKRLjVgsg4/FopjTAPb8NkLuortSIEeI8CWby65X9KmY9VgreDNIKrwETYH
CbrAdiJgvlHRNB4fWraHCI1SIuMv/e8w9wML7aoKdiMxPtTUSqcjQCHbGUv1/AI7gTdwtTyoZT7X
UWRZE9ruRBXs9PnsAkFajqiGneVEJrP7RFePm03Aq3+VElzbly0Z9r23QjBk3w19RVQ6PvPOCM6j
pPLFyv4P1sj2d+tEeAgGshd5W1mV8Tswa/87T1fMurjgCSZB+jmcdnHC8VWOxGBuaK3lgs5gUNgz
rAfcYHP+bU26Y3PRCYUKqla1J87DtQuNwv3twyZApz0aBwZ5A+Y1tPkZ2lj24aXpWZ39bGeqnJHA
GoBIgRlHwe0tAXJbOXmZ4U5Uspmr8nmHL3BWZpMRcuCmiYV3ai7sZmjRg5dMyEdqoy4oaOC1tdwn
Ik2sKM9q5ItwLSg2103c6nR8djNlJSNYfY8EFJ/7DYdoCOKFv41o0l19OhH5sDXsWL219WNIwxiC
Rw6BiWdKHXpliZ0Ni6btt5QKWWYPJfmq9EDts8SNKCLfnbErVPWVSVDxUsJQFchv25F2YqeWbxDL
r/qlJoWefBAqMs1C3cr0cMdi/Al0zMhcfsBxIdzmhfiHO4db5sTWmNv6zkbm+b/qsq4k/Kx/sqf/
S2WHem0ATxPuuxc2yICBUHEz5A83rIi/IGF/pGKYnPCVlSHGunoSPjcqzgXSvq3gmpRLdJrGPpTn
IAYKaUtJ7u5ryqgx0lq/b9l4OQYtlsnHsbgbh/vyiX1tXcpSyDE4MBxxAYuMqhRBgIH5cit1Lmqf
lX7ElvYr1p3kPN06tp41IwLgPUZoYgVMr/uBikTwCfzzVwCD2VxhUCzHRCPZ439jqei0BrCorzm8
BJ+BcSosznrEPx3A+cIy3PfYi25cMPwf9kHc5L8XAjzgSOfZnbSGidWSEbBNhT3FwQOFVO8ULT9A
m8+/TEtSDTv4qjS7ZzZlZUi8am0xnvzvA4mQF5jscZJx2A0d6bJB7a0cBysBN/mbaDzOgTOsnRlf
eiUgscB3XIPVcGbxHJVIqKyIHLJRxpJ8if6n9KTqJHdVf+DUFDyfXyN9P7YPvJ/6mtJjiS852Jd8
AcZNnYgruoVYsHOkTU0ej7SzT4l+aRQJnJkD2hCDjFRtVqBzT7jAP8stydsOx1Q7lPk8H1REU2MS
OMWnY0XrNNzg6dY6mko6r10wxGqTuky1HJi+LxWKlE68N/CtRbfv/7LFG67U/uEHg5bcU5+w1VZ8
y0laeYB9bQXhjR7Yc53GwX+TEGIWmgbXR77mVOD5D7kkgvD8GauAGWhEfNlqSV6ozUKEq202nCr2
8hHykeAn5cNJ9f+vslBDaYToQ+bPqwiAGr7q0nEqUvZPF5/Q0ENX49H48gMV5ypt2XPbhtjef+3c
J5nZjcq77F4/9K5cmPukXYCiz3v8M5Btp7gOCMfJ8HGdOGDN4H3cncFNE/6GC72Esu7Enh6eCGVa
6mErso4SP39A0uDHL+8M+MPOqIyrRH0wAX+1f67BcueEZ6aOIalQ1Nd7yv7UVDWH9gsA8DmThJRk
ijORzu1AN8EVyVYn5ahduBJ7m2712EBGBd9RvoYXU7tLqUWc3Blw4V85IdNskp9MCjvX00XKFGR2
cF1unYnw1UqNzKODhM2nFlQSnoox98UKJLXNgSj/N2IAxYDoSFqc/db8VKKz8fvH2oHB4JGR/hzv
18bniTy5jCDOVvYV7w49VTUKucgr/dwfiJEHaaySCy2SCSGtIxKwj4qTbwDE8+t56+GzMly02tVY
sSXAna10w29jPDaFrQoHWFGGsZyatQQ/dh04o6jNA4S+u0FzAU1IW/anHICnEtw22C2zNS04e9em
y4PjzC8u3KNWs5zkMyzyS69oI3JX3GhcaJdVicWKWq76FwjoYf2vcilDweoAa4OHoUfZvctEhNQQ
MmHY0QgzoPpQNoYOCFZm8Ysyl6jAO7XCzwiu3MyT988nw1BhBWd9u+FuG2O07l/zcoD9vhuDlvF6
Lz/gbG1Emq+ttGx2/ozZ6cHIIqr1qr6Zjesaaobg6eOfvkruRampK2jdK8Pw2Qo/LL1ze+IvJboc
DLHixjxHG1yLRpuTb/mFk1H3OesL/HH7eTEA+jpnLd62s3HnCRnoeTzHjS/NBlYKXPnwBhhIbsZF
d73Ig8+JLcRfY9iCsnEa7IZO4jGdSIDDg6S17ZYomic8hSbUGZNaY0l2M3AcgdXm4RLn2PQeuQ0k
ES5tSD0KInq5FwF9q+FDoIQ4ZTIdKgVjlt3wfUed3pFBMQzhRh0mvD4vA/knLn+LSdj+Y8lr58UH
cozUsCQZJsWdFzmeuq9tiemLVkbPoyod37KeymqWrVTOxBdVhJWbrGB+ay5Kc5xDu1doysA/U6rD
XcP2YNv0GXRVXaDEbhOm0M8IWxub+Ayb79zwACQBH8P9BL62Nwk60O6g0bhHNK6tn+za74qGFUdi
vd//QM0th3Km+SR6x6IoXVyzmw4Zfb3qgGsK71lordcgRfyTa4tvLIRToqtRr9yHFxrKqymn4AYU
gVoEAr2lMMTUPFWgwxiKdxLFmQfCZHO+SOap05ny4CuaXJCDeJNXVOdG+ETrHGrEvr8XXk+X607g
j8E/CXg37ME51J8Fs8+Y3AgZ8SW2kJzSF6gjTCropEhJ+Y7dFzynjrJjkAIRN4qgLGc4cW6uYtTL
DV9NvKO0nUqxLm0Wy+RIcdp/fcrIZXtk0BKlqYqrh1+7ypvS5pI/mi21eNaW6BG4Vbzb9sz8PD4O
RP/rKKXJeuyd42qUHD+jJxmLFehajtxaN5PAHo9zCddvCP42Aqjv7ay9HdS1PI3kXc0PE47iI7+J
hUdpn0u7EuvpX66bszUwlXc4fhKyXcuhaOvGBN0IArKcKGVcGAqiifaODfUAa6IgoaGoVuBhxtJK
uIMF4N1rECy6DC5BrfUbd4P9YTUEqVN5hv9Jg9UZEeURAqb4XEcqC0QBcT829FSlXmiA6ZtIKoit
j4wD650wZjkjGuQQ7RzTSt6yWqWeO8Gyng5FOgWVJhNZ4shRDbczWwroYl7iJQvJrWT41a9ksbS9
ms7HirboaMy0zNQEcyw5SgKmHJStQniHJh8GxMzvJtcgeXdXZVLKYb2+ka60OUyosnJYdFptD0bL
U7AUBMco+gOVLtOtrD6AAIVeOiDBRRzuqh9d+ohYrEDpjPf1I4ianpHR7P1NRVBgTuSL7Ts7tlEQ
JiWjK6VJspFr4fvc93PCJeqHvOq+9+j06R3ZOfeo0wOvlDnvMTRdsJH8G7xTVofxUAzXQ2/g/CbG
3V5SBrq1MsUD6/TETihXeTwN17A1TVwGct0efbLGkD+olewiEC8HtvJ3kk3Vg93GwRmxtZQBwaNx
eRmnMCY+qxnWtuxSqYIKxKmbyxnCQHcYyJ6CZXSDS7BAc8c9j0v/bZNmI7K0vbRPh2yZ4MVT6AQT
FWx032azGASFyJcM8bP0JqHYwGzm9W+1SfK9517tiuzbB/My2pIBFN4aoOxFytMmo2HO1Lx9rvZd
DmkqDW+eB2SHoiRfRJgX1qiTEl+r/SuFU9J0E0OIVbJi/pNMrFQr9OmPagp/sSipNgZirMC1WqDp
+2TBYAT4G+oTVt94HBKkSw+gvAwJCQ5HXPX0R2gl9UbUIYKzsPj7q1nJuVn5dwbUAoV1y1ZggGwO
3LKUSj0Xe4NYiHcgPYA/5G8wq3rK5/syhpp8sFqUf6iCMra9Ok2Z2i/PlaXMNz1S/kmie26TmUPJ
pjh+UeJ/ANfl5IGrlTD1mDrUjQ/dPUfGUWAvdcL5wcLXeHKGT0esI6qmXjpg99m4txc+ZrpFwb4m
4WK8kCXvgZvpBj3DMIMEFnGMbEVe5uJnqPnaZwZCnF4RzMb9++ysln8f4WY9e7xup96exsFVrjdq
1t3YrcKxzTQ8oe2Nmw9CeWjk3fS6EVTbaOx80wd2EaNKei9E/GRNuop1q8xikYpwa3QfBaoOUHrd
JX65bL7ykv4vBc8xC7yZKy1QTfVE+cAuuxkif3UcRdhVfPmBPJlOinTIoksMC8NExWDkkCVhpa7E
UUvplBIuQiwZKB89FgAO3nlQFRL2HWG5cVNdUBPbYWOq1nbQ1ZakcoZ1hAqviYZ2x5xhi45prY6i
3xqAvU+vZBEFhj8jCOiegbweFcZc7HREekpddTRNQgIIzXBEfvTGiUc8qbxZASC8G0g2Mgnd2eA2
rWVMJxwp5LfoAaaCA3Amxt14W1lqEfQJaJz5mP0aVkFkAwV4VS8Gt3XJuMck25FOrCHqs3DhtS/z
VGpoz+xn2B2hNGlE2j4OerQLHEFc4S02BGYo26n/1yZstwZs34TgzJut1H9BjQwydR/XQc2TuX3B
MvpHfYqLn/KhqoVoH2AILH6FRHBkKvq7WKgN+k4dLWTO7nnCiEIv/g829S3e+yI7rpQ5VhpPmTey
olDAKho4Xkr3YMo+NGNCh7VUCmmX4RFTQCnpyv3JffOGweR+appnyK7jBFC/WJCiAk0o7uA6GhWT
dwUkjEVa2DSPTpMOU6YpbtuXtyXdAZv6pu/UKRm+OvGsUOwfrjwpYSbR3GE7nyN8oSVyVuq4TBoK
w1BCzfrSi+uff1abZwtgnpYb7G7DV+aE+bwBr4ge53iSa52odjnGOfICOXc2DMZ5RI8XRyGf7EZr
TXWSNZxqu6Q04ZZI7Bd4Tj4ssobI96YuCo2R40FgfGItFte84BRJ/2cNIKYWPFKTj0YFk4760Kh+
wi5II25S3BepPhg3SLdRXPbCG+9TUPdiwZi3+e4HvMPvIwjn+C2RbYt4e8zup26B/ptXGDvuXp1R
NjM95rnTxcASlK/NS7gFOjogMO9z8i6UcWRpKTejbRDYRvdLGTuZmKrPkZwi0Pf8XfqdXBJWq4z7
dfJJjIYsl/CQobSw3U2ZjD/04YXQ1duiyJ1Gf0VvCU4WqHtUCyNsgOrUVhM0dTe/ND8QLqznxhTZ
QgpRvIpjwMft7I2EtA5RHEl6C3zh+Zz6ZeC8n1kAOtwJxBboxmqSNzIWnqIfcngh+jDaudNX2AQg
yOqCTqoDPn2pligYqB5JHM/hfIG5Bzss60TbftXd3ANBuUx45MnbS6HPlptosJ69y1smfTkj/Vp0
TV/I9daM8Iu8OJNKxB9WKDposk4gFpcgmRSxWEMXifstX4Rl/phWzTqiPg1VDgGIPaqb+cNFAKEj
mytSyj+++dTkyrYpIQX/W9X4dmQYUbYYzsZHaTKvtXM86awSjnA/KBwhBRby5qabiAfjWrfcfOLf
5ACDkJOl6c5wn00RMrAUn96kfxPKWvDsPCSBtC7MIZP9cUzimdvxsD5b5IZe3vKORhUOLUIKiyBf
t5t5sOMCuvaTli48wb6LJc6NU+qDnwU55VJmKYJ+0426sZUd+EWJ0hZ4j9t8d1iaWtp0llPcAgT3
xqr3Ucgqeb1YUvIk3+Fk7s5QQ77LLIeq0VeGyFrbUPPSV0x/Uzp4oI07QLPNahb9QrwlVkZTC5+q
swTb3Yw8d24XDZLlNDJwhlp91nTTVBjBOmTDR3WxDgFmfFzF0VFJaZp8iSyNJ5WHMjlKcBQfAE2u
x1NcUVLqyKQMJZTZYVEFfO59UDUhaTRZiBqB0GH0HgX8h5WjRKuSA57wpR4p15bT9EFWdyK6betp
AhcjO519ab8gJ9+a+ei56XVnTznO0LSB8RoHQJfzrfNq7owmzv/Oidemj67XdkReRRDnsURrxUcR
5tLtImIuoBSPgoH/G3DgpIvjiG5Mgm0/2sR2If2xMLu/21NEwYEhZW6T6NzD2FwpfQkkIrB33W3E
LoTI7p1YjKL1PQgJo6UrZ/Q7FhjZQdDXhf6O/YWy45qB9wpTA1EiqgpwmbsiGmlT3seGlETRW8FX
iUVrEXrc8HxL7AD9bCb59ZV8RLN5bwc7IYqihluyOSSybPHjIao6fQJtexeCh0d10C2+Qqcorpj8
CAJ5P+Vi0Y8Y77h6m5hEsYAQBJmg+ixsbhVoUmlzjmPaV6WAfUBwKs+Zjv0StAmkxmROoSGJaXO6
J3iT6o20HRKggsbbDeDlnpn3jDaMfdXLq8x4JoVqmQWmb8+FGX0nhoLOUHZNmJM9npPcr43yL3LE
qaADrPjneN9/R27p59Hhuz2nYA6NHpnLgE1lQBZ6qRBgZjETDZTrJTvT9LuvMxz886dpLV74sGrH
+7wgeDtsGQQjCDTcJZ8fwRbOqpqsWgMx/o+rLM6KDxw5VXE+kR2xaXMtJ+lBLHoVnDkrPzro6GcW
gNGXmOnU+hiDqo2NrRv4wUzS95gBuFdxSP7KjLuVZvgKMH7+BjzNGBczS1rU2uVBm4om6ACWXT0Y
DO2gtu5fncxhxvNn3R0NJCybfMCtgGcCceOggq9gjIKMfqqWkBDz92eai5CC+FPA0Tr/cUhz9NPj
kSfk2Nr7000ExlUSLpddjikEVOHlpZznSCGM2zOPhv96lHTiMVEEnPez91GV+abCqzU+b+a0EO+j
x/r6L2T6pkZqbu7nbMGgy4wtwoxOLRcm2Cofbc8G4qfgN6uoGJ1Y3rR5odqtUXA7R5DtpoE033UL
DqJkQrMyM7cLgn4xKmB5Na/q6eCSHzLSD/VKmWKHD9AC0nlzhzuQfaSkzNUUKKDnQX9RhjD14B1B
cAI5CeHgWjda8FrnuAWDadi9afCUAsS+enFYPRr5dvdEuc4P+xLTssResrmhcJ9qLA5uPYhGzc0d
6t2HhAO+hjAg6NBm2tWaq8R3QN/iyN7DkWoC+VmpzwPuLGIrMW1iAuOmozLtyfswfzQpiGlsZwoE
419KLSHiLQfi5hdJgP+Pk09qRZmngjHv3+XfrDbLf737qT4nsidsxjsM6HH4n8Nz4KQznSeDtKwJ
Av2XVIVEgqUoeHEBMD1vrqScaZ0zV/YKbtZ/XkX24wlWCz/RmsyUDKjVWPHPFtFhfxziqPfbPBWl
U2MIKJyfUvGFzOjjZGyT50M1j6HmlM+DuQc48AUOmI6/E3led/DNSwLWh+UXg+C0HOPFQhrPZP+m
sJb0BfgeZSNjrPJaJTKRXzUtf97Zfy/MsFf/iOFa1bomBbRqb0dbluXf74ooQOlHy2W9lcnilb97
xMtVJWv9/KqNuD7n2vQI/DozovvJOy+riQRjwAe0ilH7thonpz74X8kXVtXLXpxzh2uvRVPSYz6D
8VfPm0z2VJs73lTq1gMLlXDQxQsQjk+kiQ7nUFUYHUdhJPJOzZLhDXOaYzOr3fR9WsaD+h9Y1xAg
7hnLvQV5/vYsRFePgD23bcJHltSHPXpfE1aoADO/fuxoF936C30X42hzvRj84yGORNxQdTII737e
SiLpSpEWWK+Vg/BVhMPVB6Nv8ZFciOFnLN6bGuFz6cB0TdDdfK7/r0td4Jg8g8p0IITsFAaJ/kqj
UlPGTls1JfyNgcwCf8rXE8nFhW7aKpQOOnZgJMUHG5U1VfotD0oS6r9TdBwrfHFer+VBMcOM70ix
QwWpgBEYzkNGZPcfx1N1onUmk6KTpKnh8MNn7gTd5hue4QS39s6GygjCXsDOy0s6PbMDeyEV+UdC
7roPB2a01ZcKy/Z01HjbZrkBCz1GDSc7JdRs6MGhIktVTGMsnAi6Na9yTUMjW1Kshaok97CVYrAu
VO/iCoQTTo7buSw42Yrvn9LgQ7CNNP430UgOiYLImchZCNlm4KBkpXW9flmTtzKipFGrrHfbSAvD
BryFlWBKVGW9FKlXzPNbVWM8XsIAxnl6+wHF/hVuS6MqfJ/64S7/pgmUWfKIaDeWrgvdpsKU+pcK
FV3FVbd9thwTM+R2TFuV1ZLV7xCVdgzp8xwU3NPvj5BFgMdoW4JRM8tlzfYGIwmynL2pT7mwcolA
sa8WMMwDd4DsQ0O9T4TM1qw43W5VvYMVUP9JpipwvVl9swKbBhu9TODCozjhhKTxyZn24Y2tYMeV
7FRdcR/jF8YPdGh2gUginEm0kVLMVCI+L+WEBW1cv3WIKtq33K1as8aA7vXWG7CR+wBpeeTuDxX6
zRppbN38uL0fPy/7uCYbCYGY0KntMqOwd6ItCxv47sNRMlUkgyPO2ur3fEYLseU4kHP82R3SM1de
5ySDvZisEIPOOLe2lByLmLkrvAV/Oqd9u7yVrqNj8Dl4iQRBy/f5xE2J1chyJW/uPFUfFhIQVopN
gYSqIEy1nb7MFqs66m0Lu9LvYeNrRWE0HGG1iYgCMJaxr/LT7m7NsH5hVrv7sq8yAcym8SIGapuA
YHSv5E99F8ionTPxzlPMZKw/qnFoXWC9Pitdxxf4FxjQZCYpXv+BLBNQVloNGsnld/0gGEGGnB4h
GZDEPV0pcE6kHXS0OYcht4w5DAHmLxQiTRTGXIizJH4aTnjxE7rwaR4POieXkBj0dDy3i42EIohX
axVDYtjlm+A7VwWjsqHDGL6jwNH/ST66HwL8aDBl3He7UCf2vugo8Nt8d19kepD70XcbHT4Twcgd
5OFeZD9vIpr23osL19oo6H5NKNQ0+QkpnSlsXX8Q2ErH8otK3eJyo8v3C3Xdhbn35jmCmC94c4tQ
vb5Tk/nry/dqXxI2KCdk40JRkXo1Y58UvgZsnx0ousCnTJLso2+CYaxLrGQFwZX18yjKaeNb9nRj
oYYcShQDUc8bETQEe5P0bHqGM8XJIrOM0S7wdWlDtoWNGHavsgCRpOD3gxhej24dtmM9rWcy1yT6
2q1jXQNcML1SV0HePscOM5q+eRnD6UY30ePe6IMo9acRZj25nh/nyuIZ/6fHjxizM8nkrJfnMb3I
sH4exnepa9b4MNlhVeao1mXFLgALzuLTEwAQLbz9mAs20qlui0UhcE5rGrHwkmIRfSFhiYXWysNT
lQuhBEAPtMLtDZymDGp8McpjK/CaA8lZwOmAMWsEepSPEnW6bAEUk/pBBOwH1fBYwowCshvJ6ONw
J5FB6K3FzlkgS0pCzEKfNTAOwjEez9v9VB5/uPQlrbPJA1cB25u4yIhx9IRn5b5WZ8Uk80dmEJ8c
+Gt2BwK158MhQWqf17fG8zVZ18p9zvzhgx6uLX/ktrILJbIAjtfs608HcVIUBobfrsWp7to7Bquf
LJb8Q1tpcm84wcSSQEX7mzA1p7dv9rBVKAo6EgvioqYmVCCKVPIBaZlBGQZ46OY6TYwbs3v7iMhb
t1tbhJrcTVL4NjSXxGNH6BYGl/0f9usH4gANvhrtANOjsSMxC45dwEr5PIogxnQzTaM0qJJicwMU
a+2XPY9xBC1E7R4WuHiAA6wAxQjhWlzhyMOBRcY6SPGEStGBjq0WGc6p3AmAuR3EkJuO869tHl5x
ASNVZajtbdtN+HUkiJS66XKf4pxCd+54XQGtDC5U0vq8mCvAvRDInxtZBJMlzjEDLtJ8+VjxOIQV
PZuaol2pCF0QqrKvAQ7pspWFuGQC6F9gM9/HQoiMTVpX7Cg6bb9SnzgiUSBXTZFVpzRA3AY/B/QS
E0WAKWvdtLnWXavhSLa+KsIPxwinXhqRcn6f2vYQeRja6JY578heKa14RH0UweAr0nDH/dMnKZJC
XwnTY2fIVSrFIPKIiQcWVPx88+2UVYS8v9VcOnoJW1PWLfn3GMC1eVmjvQBaBPc1/K4jqMRTZFMr
eUDmtbpZgzhPmDq+gY/OijZSWDfMfcpg7kPlX2xqdQeMB6HkqM8OyMU4AUs9uaCIFxM7YG/dh5WA
o25XrWTtg129dqqdbnJggz+x7u8Wmt2aUp+EA1NW0qm/xpHt22dmPtdwP27HP041ihDMYl59OmnF
M8k7l+psvC5gPQkj37pUHj3GsNJzAyY6wHiDgwq1RgCQh2rka7Z8bnJrFGCfTF6yRU+ppdt3zn5q
2YJIcW9lg5C5WDjZCviBwFQPh3WTcHkgomAFSMDTNxeA3FFjIDtjHR3Y4uAIFOPorzTJZVcDqCIg
4szOZZ7oNjRMz0bRDpvNeFeadu29EsWFuAz8BUQWwLMDlODNVabL9XSiAV+pQ+uvfKmBeZUVbooQ
U36v3gKDCZYtf0XkBNREH4v3qgUqN2qQSBMQgSmb43uf1lZ/hWPvigVWCuPArTSYZT89tXaeZSKa
PZ9Ibb1njKuIU1NFa0K0leQOq1w6NSfVZkHdvoUt2dvH46uz0q4I63lKjvDiII1GtSbM7DAbm221
JjGBGPuasKk9dnVWCXJ1qzLj3jgZIMBPBwZguW3WRhlZxBeRoeW/Vu2NFCbDAN9CeI59udn517cT
ABU2ZlpvgDDKvFJ4KhJFs/+MHP/Xw0QinloHvusErRZz2EEZaxsh9jbovIF/3Uf2byLzAm1oFgTQ
d8FCPng6sjmrBTfoX8oVKpk2InuQl6WxwyUJVorrTR9XRCJZjSpE+e96J540+cOPTcZId7QoWUOw
KW5yUVkxNGDCX5ySXdYb9vym6NwOdGLp1eu5Rg83w85/Mbv4Q32khknI6mOfut/czLHphEBV9oC7
h3xbyUk+BLvij8Kyld292kCuwPeG05t49NEE7r6cdPPlvMDDZXxt7T/CT5xntIopq3biNBfg6AJv
PaHkuTi9ikuRDdEAQDHtNRaZll/O9vaTHg3B5ZJXS9C2COhujeLiimFkKCBJxNlDIgdPz0Ei1kxO
0+7B9SM6+cE057lCZRNzFCoOchw6qnTF4sNvzpq88Yytd79CwhEPsROoaAH5gUjrht7J39KDQqxs
eifrre8iEh5+dl4RUbF7pglPcd9YGqSCJmR77QBNIQmGj+HDXXmIrXi5QC/Oo6lUfzcpTqkiC66l
jPMi23e4klp5w++RZiyo104NJoq1B8Alm2Z5Tj+x/3s08MODOvYR4Qyu1sjzCOv872u7pw9b5EP9
6CU4pYA2F5imYgx8r9vueqvlFLBmLebWP+LPb62zBmyF+r2Z3AHcH5XMw0+qmglAOWv8AHJVIBFQ
U4t+QKL1oWoyCeQI3cd69HZSaJc4Hn9YwJb1eRkm3SD/rx6gbqLkGvxiXJv5gaZOpoQAWKWBJI3x
NE62YGx+/kcpNFVNd5guORUu3M/nKW+Wn/SmatoPKqHxB4vIZNU7M1hClbBzkUDKBTVrbim4k5lI
5X5Vj/WSp9JHFoyMn2BeRnfTlavTfcy85bBu0pJNpS2Q8aIuegw/KiUSPZHt36p6uDcAi8KBrMtr
xbATFYa9RPUv+iVkNJ2c7EnTbknU/Z16M4Ev/lnlb51C2gg97huytIHHJE9BtZUi35rcxF6hYuYf
1MhxpHQS4zZTXAi5CP4QQOwWyuDRsK9E5Mx4JPkprdVDZIJPVcAuC/UrcuCCCB9H7g/WHydqjEI7
2/g3t5K+O3R5rGqUjZ1PDLLifLZyD8NDjhFSMYD5Hc+LiAVTrh9YZNPqlYQcE1ureMxywFr9CJLz
P4WYVhSpe5qIuuTd+wg5P3qEGlFGXIKL9GpaHfPCrdS9+qdOCULPLJUxeAfOZZAW5aDCa7ZEI38P
Gc2oLxteipzWRYlof363nscP6X8xj3Nao6QsMKZ01QiCD8y/0uDx2SCU/BG6TnkOCSuWjjU/TEl/
2UzW3r7MP2DtMSIrG4/1H0qiiItYHKBMboqBZM9G+i7cgworVW0SIFWEY8Sn2WxIDU2kDdqLRjEb
9lLmU1KbxbxZRjMaJtDy43rsoiKQ5eaFstZqOX6rcH1UIzLNDI4VjcbXDxjSO1RcgOPh/cAW+J0O
QcECqO6/a1M6sojFNc30G6tG8uI7OEE8Yl6dwpbRk0JCAqrstObvTVzw8ogDFb/euquvmyfjXULW
bzprZCaSqGmSMVkxQgxxAy3CEMTIRF70sghUbPy1Gn3MG0mLaW8oIf1h8LtXeX8NHhgrBag0I9bi
nvYnHhUPtj+9xVijkqg4rdEJPFDwB+ffPBQjykkP6bV/rkTu3Y29YIoT4KZJ1XQ8xFKMn2U7vAcv
kjfFThGr5bm3j1h6i7ItDRnnn2ojV+T7ZzuMqDTZPGAFZDkqJXQeuN2aTgBYV9bCJTFXNZ58Ps8r
piXa9zLkDYRUdVqs2Shz15vEr3AgEFGU8O0AqUKrJwO33BYB5gu2z4EagqFIODoEux8ZYeG2eFAj
opdT8gxRnysB0uRHGS08Q8WFUgGyXLJiHxVDzeojocRf1KpBb45BdwGyVISMrfp9ca11Gm1G5pfT
BmsVGPnm+4cYOG6zEFhJ8shUqLLYw5An07CGPl47funbHKCvk5iN1sTugAkIMAHsukexHqKooKzW
Yz/MoLdXh5R5UYGPRBPDG96OzoefP49timh1vtSBBaG36WI5ZrwaIfseZTwyMjw1R9OFTAkZsEAV
vylElsTtgyL/CsoDyxnIT0VonQ41JF3t81kjudD5UNT1LMK1LzTXwQ3+V8S2nDA59KnluPfXQzL5
HWtnNFGXAs/j5c58/C5Qkb+/CHXpqFgNbix8Pn3DzceDXmia8/DCBiVUZTxFXcrNyoy5fd4n5tIi
gO5eHlx+4VsfkUC72yPg2WVH5fBu2Qg3O2L3lqRCSAEd5gYc9fRUlbqmANh42wm2TtwIJslWHCad
nAgrKl0fGdH7cLLcyoYBtn2qScMqMDDf1ayxdd0n176/lDYiklaa+aO/psPX0aFx88YctEYdmQ9b
1OkWGgm2aVsRXg4SVpC/ja+mMW97HV2LByOARWcSha5nd0/XESvbZ6Yaykg1rsRGRDtYS5XGXKuc
/+2CJhTvpkkQ9GOEzQaIKtEi10/1i2JznzdtpXp1GH7b6opC4CXvvH2N1dw9vKencpd9gBD+BPCr
UvvrvJ98xm23BTqJ6RO5FMQHNhLvvOIPKhBq7KR9pHRDgafDn9SJiqOlvzomSTtecyPka7kocAJZ
HVjg+tuoeFB3ObLZvpWXVlMdEvtjl0IBJtRVCNN8MREHfG7f+ORcl9X5GrZ47OOTYp5s1f9C2p0p
DeJxnAHn5Hz5lXuvVzfSxNjJbIgh+d0wLGuFD//O1rw5h24l9XXADRP55JApgl23u8kJTEmunLwY
e8h3AVWyVIHE/o+13s1sKkj50La2oh68+4Iw+6hXvAuWcWgsPZMoMiiURJRjTwuyn1jHyYVfXZci
/eRQHJZxuWRv/EXSz1WEyNdx/FeCUAr87Cq++In/RYDILDgUTkU12vQDWl6OSSsOalTQkCcPXsCo
IcwEdTpvjnOLJ19Egu9kdqvyYEmZAiVSgVhfPPvjeo7bGlRUzELIvOY8Azqg8JnHSRtstkJGOCMB
qTtdk9ghPVRlT+rMz7Mp3nj8R56AQVPOCxd/iIdcWQunlVa50/dkC+3FhpMm2PwYhcD2xLdLq/Yn
7GTLSpZ+Pm8fSGRCDhdJUQamw8He/0JzDspSOVyQq53OV+gSZCoWDFYk15sanPykZlWeAvkUluzL
brFWGvvFzGAbdglgwRRzZ2/AJqaH6DQRHyxVLbpdWUPoZPz/DJ+q6icqRKMUR1XR80/J5m//UsWI
zY81F6Ph6IKox5559arybJxEznx6PnPIXB+8W6fto7JzUtxtVqLtVU5mOPIemSxSqZD3b7Lh26s9
bAJ529FhFLm1dpCO7YA5U2K7CkAxmDnLCLPG8JME8I1AuIJEym4j1Z0f8WcyPjYMLr/c7bKbIWv7
ZdXGozddWJ/OtS6InKBxpUq45V9rOcjT4hQza89CA3L9c6faK89pSq4c7PNJvA6lvDJo+d1+Op3S
aBALLZYYPcxNhR06P4/XJ5hPPv6fEyAq3CSd0r0mm3rqsFjf0vJ1EJH9O1XHIuz8FONKPzYX6FhA
dVHnbf8cQULNsvwWXu3o+3ZQuscMcl89wqw6GvZC4mEnvARcnvg8sRrrPO1F4V5d1PahsiJluaVI
5XxrrqglrsNnSI86PEjK5uDdrW26XqJlNIE4nJzfURbH2RSEdiNUEVygLAxwBw5cCM1gJQPhzOAF
bgpXAhY+L4ZHPgq93RoCtkMiSENSAXzBiJdQFzBuomumrsKpy4nIncuW13YNtO8o5VpoWDFwPfRA
k7YrJ274aJUO3khyaB+XX+htfIge3pQJy4rjGoEGXi3LevK3a5sUG2XUeYh+IxUpVz4WMJNKFGS2
pvVjHA2QsImnFDXMvFuaDUUEFBbMcb86ibpuomlrsLiEnkzC7SqdwDniA2z50toskYdWQ1wTECNZ
lXyDC2Qg8ruSmHPHOjt+G7SDJar3t/9OMYMnlF7W9sXJJF2VROn8yTYwlZUkVkeI0epjfUePHmsT
Wz5LLTr186+xzO4SCpaPnmjwNUbGOBE4uURLND/NT/3gqaSYsXgs/SDMELyo8zwbeG90UM60CNMc
JS1xCCxHUKQdCw7pMCHLnOrZRx6EDK2qFEwpuc402ZmGw5XqBXdXE+yeEff8my5tBjh3xArSdSmt
4YMqJRmI4GRijSUksVClaBX9qxFeJG11HCH2XZddF397EYftTCFGph5B460q4rQ/H4MPCNHCATCl
SiiyxN/9GC3F9clt9Qn7qgqa3VEoMMEIzdRm886xNY4cqZsIlhlu9fRjIRJGmM5LIX8U9R/mUtZb
vgWBSZqpRPkUZ0Rj7bDGQcu5qNjV1jS65lBZ0bgxJERczejjQ0yvG9eMMB/pwARqxvfweNjHG9QH
uZrioBlvNzU7sgaypobH4w+GKfqT8FuBrSZpZdS5gA9puFAFlt82lbcHeOZZ1QLKTtbasK9uZYIf
0bATKihwmwkEB/s5xaA8RTOpcl/vi8Sya4XMzkxyioleB1sqsXIlEVwTLI7rfWXyzKZw+CpvzDlc
7T3J67HRZE8geFUHOZbABTNffLZPrpoBjKvBmTjwJzhafUvHVyP+R1djq93gIPCBCcK5QQFtZ8Ec
L1lgDgxN4k5nnTQ4CVk0vQO4Hq5e1ijGUIXlABU6kOK5ctQc+TC/ZPe+fcL4pKWyzEcuDFh8aQwB
UE04Rzf0KjvER+/kqX424aiDNdlToBVnqmH7B02f2SV4V36gy48/ZEg2ZhxIDONKz82/7RHe/Zk1
bTNv0K0b85ncqq6893zGH+NMS5jRm+PaKa9TsFb8wS8i5W9FXdu4pX+YSATaDgUlZXUfOKYo73Jg
7N0niMewv7yw94w4N/NZIM4d3r8gax1HrQqNvxvZC7i6IEDzzhWrJk32oiV4uO42HTRjTJj2Fc3Q
q+nsCFOQ7Nl2xC17JCo7qQO4vt2rV+yNzVCHk1aTO0EpREYbP48jIl0a/aXI1M28JgQNM1mYTNmm
wnsMQGUZpMGHZ9jhlZOJoOiaV4bZHUgH8GPlzBH5BKP/ZmVUq6xwagOl2s8c7MUGJ4DZ+5yuf7QR
FiTpf4DCwHNrUOLfZqtgoh/y5+JoKuw72OiUnwetlNK2ALMoDJH3MLK1eCxylgLJyHfi4wFifwZT
kU8FmQyx93CXZmEBItCsThyBNp5kHXhKK6pwscE3WRimm3d9ZdbHcULXIls2yN0DLrFGW/cbh9/6
O7gSywPpBli2HTvDTtMcRadP/dRR38NJ80tABGjXpV7I/xbN9Jl/q7Ec5/ohaaLt7sCY/eTAmi2P
vIMtH+yb1jmdfEOFfbKCKzzVON/6xqDNzJ8niZQx6CcegZdY5JiewwkSrIHpbrpVVcO8lh2zychO
G9D4M/+F6mGS89sLOgy9umEFgpa7urSacpLLW8QzOlEtBHTITIwCrN+64qvu7Wr10rbKl3qiwJK0
yVK3MLy8VCRHVg9bc0AexduD2ZHx0kzp87t6Aa/yGj6wW7Yx7FO4NIyTko8afl6VMUkF/d/dyP6y
BgxjxGsS49TzbAh4tyNCpWHeEmfjOkE5tkhcxYLcUYuR4N6aNEgGlGGJaGnKrl9SKxKVvmbDGhAt
84H05soyjDNW3PEuOsjNhrbWLzjp2GYtngkMqN9+sHL3MOtoNBpyF49NSQ9o18GeHmpTBdojI93t
P8DBxiXjp2GLVayhqAxsPsS+NTBRcXwurxq9uOOqxQ7aa+acjZViHhSfiqQSAzzRfET2eBgQz40M
BOw6smWHwypa8eQjFK6i9YXz4NcXllw466PgknfvnSHJIVG1+FxWiI1Sjpzschyt9FNpv/vLk+yd
RInDMBqnNMTiUfov9sFuJLablLAFsdR1ma94ld3u1qLSFWqAi6H2IfyIKz53eUmUuuGwtXvY6HLh
8MrZ0hybkNSKEaAUDGH2KfWjBSAJiFTcfV+ASCLzniowlBDAN28wYBdBlshn8frnlg1wDb9k02bO
MA80PhIoyon9YkLcJSZ4ycji1a0j1ImGxtVIXhTF1p6WM/syALWOmBrpIIGNp6zIpOcFFGFV25/s
BwEySvj6yxmyNlRBRqmFMLhGQqdugOe09i+814hUcDAoBDqSfdq5f9Koe7leX0R4slP0g+iLZLN2
ZXQULJa53eOHby6fc7NXOetU+G/OWCTShBzjw64+EBZ1Zh5a1lBvw25IvU1qUeKvxJ6odvNSLIcU
AootuZgZ5nE3AjL5SnTmtTvL6y0nI4L6yeWzf9rhPMMhOv2fEXITodnhBB8SBvpGHy75S2KhTmiJ
6Qo634wMa1sBzaWmtq27HXdp+1gps0lLnx5sExXiRnw+mkcH/OOxSZG6ZTHbImmZA7wrNi+WbVU6
0i0Q2jLdGATRNGok3imlFw3KGm5HV2vewnh5W41VO7dUmLIfWXOPuSLYLdT3PzH5bu40T6Jmru5c
wOHKt4lA2sT15gmfOXiPpseJasTYL5MJudLBX7FsthbkPbWONhjX2URsk+TxiOMvgiXQBfL/qtly
lmzqu/C5u+IDY4+ZBNqALL/7VI/lL1W3cVVTaoAuVGsopROsCPmEkrvJ/GeODfUUJjHEWpmjbsj6
/za5iugL2ST30f6thULrnhtWo5J0lH0Pd0yzJCiecZm2tFSt0ovZna1AWxjXrGpxfZpQgLNQ3ms2
MV3qzNw85MGpztlnE4tt6C+dOoA1zYPFKOOnkWKvcdM4ztS8QIq3OuRJAFJJ299Ke0+fZKivKWkD
gua0e2IympdwdFph0QfpKvYuXIbw8s512b9Hf7/2YgGgwL6POtcWZ3tKPo7g6atcl1zVk2m2d04g
VG+KaLcKTU4EbkxtAyDvMqBt9SuuVjXSBdOPCVC2ImaQLnLE6hvZE0vf3v6ubKs6kAK02G40pUr3
xO0t490a/1ts8QRDqL4UczcDH9vPKBF8oMN9SOh9MaImzzxsFea9CGnU1eE5z4wIVBNX+njwnHaf
SzKYL5cntl472a11q3QAnDDlDr3iIKo912LLxQUyXgjY7/Om6wJGXgeBE5j6zrp6s9lmVYSOJOdf
M3BXFP27kMgy7WrKENzcEnyBrypUHX61nWiRqYdLCr6+4bO33YS6xtF3Y5A/Ey+QR6nIkQuE1kkt
Pyq0vmPvzjMIJq6yvbYNlsEsx39mXFx/SNDntVQ4LB6+vdA8qlZ3a3Ebaa6i+sdO33l7l9gQr3VV
Dm/rfueVGJy4LNn/Uf4q5ayW/7E0FVh83pxVQ13DD7jicH/WIJxmBPexkqkge0pJM9zPcjsM9yYB
ZqLrNk3fIUU58aM6+KvYW5aXWCLz+iIQAyqVLFNyWlyYENMH9KJkYRvC+aCtcitbUVXkSWORw+Wp
Yujz7D8nnxA6Mt4VWdzGmn7qYH8bArp9BnXXCEUrTRiMhbTcXmSoghXhBQl1kfLFfXVkwOlfewtR
GehD4Z49e5lInMvwqTRILbnMQStwnmVd81PUbYjMZLlszNs4Jn+v3UgEt2luEM5zRZ3fKDyaHPz/
BUsx3gEy1+rNsnH53ykWs5m/QJLm9D600a/3+zlKfWos0j9N+v0bs9GClmACidPMrnxZLrHqc7GL
iDD3Ub9ewowC2KG8PM52Wux0CiFv3pQa1zivdGa/sT5FCpFkfvJpeZJabZ+dqhxiykHgmQxMW/AB
Rs+F7GrVMvB572iseSm+NogxuCFZvery+i+WV/6UEDBkLBa8PM4np2HEgV43W0GHjUrzd8yjmrIg
J8KBxYQQEWghQptk9u7oCPZH7Mpfm8+r69zpYb0lFV0z3fjq4RZUlzlamARM8vLC+OD7Cy5KpLSs
24VXQckVcOmNukDGsgEoSTJcSueW83H7E8qkbDWoURp7DFDdW59gte/JURJMyapJI7XAXeQmEo/U
x9p/r9Y/6g4SSby1DnklWhWSbPLRqWyUsRwQha/DsJaB/Un9unp3H2WRz6H7ODGebtfqmpqIQ0pj
m4UHjg9USiiAbQ2XZWUjA4unMJXWRF5/1fJ38whm9xD0nPE1FYyJ4xgB5o/F1zF3nGSrSnRcd1mT
LWmOVx/ywQIAHFToGO6lkkGUCYM2yb9flmAvVTbnNaGOJg7y91H39BPE0imCx6Z8wdkg9jT4alE7
ad4eVNZAwDXCgBkWjBsRopG5DutMHZVdeFX5X6eqb5VtLNg9YKekZhxnHwJp0cI7O46aU72BnRMj
Ty4d6h8ZVhGSGKYBCCm5WwhE/Qs7z8fxsHptCd30Q2zkMmaF9FEotYPPbeitNHZlZ1Vg1ouzW+Ru
BXXMmaM8EcKBjuGLWUjpS3xfeJEOcxjlsmyQxfzDnYoMGsC7kbp5vtQG+kK5lqYGOP4VmDCtmm7w
Au42l1jAMDEbk3F/twMVSoXCa8A/5Z54CIRq7Mg2ZM/esQnTHzBlYYXgr8Sxzax7+5isx98iPzBl
cBSc/wgR4UnjdgoMkpBfJ5YR5NsQrtQvGnxIqogwoMEfp0RJabNFOTFx7W8ogL0ZUvt3ye4obmON
FgmfrytcVKlclsoUMYeTB6f4efJ7EVL7kk/rv1XvHuqUZfi8gUTLCfdLGLErbqUnCcvM3405Qz9p
onMLxbNBHhR+zgCQfHwGcZG2pcU+g9zt0fPog+ecYuX3u7NlMTv3cgTfQs90tAEoPXHICGT2pcgG
NuViYPvc88TlWnsFgFwJlu1Pxe1Ko/WAZ6VXowQFYWgkYMIYiS122AtXKp5dURXFD0KRNheSZvDB
nZo2m812cCnIrO/HUEg4k5RHepGYDtEF5bhBtm2zJpnjuZxzJ0YjVhvKRybYVUXwHVBSmjczqt6z
4cFROXgAU6S1C1kMM8NL42ePfgTBT3Lolhz7wdj0a/xxxr14qtcjkwgNtkyAnQHKhXFZfxBunF9p
QfqZliDr3yyXk61vAZr/ynSY1L2meAmwvT3lKSLctC62/ZwMOOwD6KKIEqP1p8XF08XPkzFhk3ih
KebQJgBa7MdJZhh3FBWJ9lB4nnq4PJmaxf8N6v0RaDHvhnk5iJIsN9qj/tGuqKYuqr/MnzekcTXa
F3AWkL0sBcqGte4f2VCkFRqCnjdl0YCqHRf+9M5pDbc9nm0B+jP6zFHsBJRRdHnssEfC59JL0ejg
1NUtObP/1GiEF9PcCqMfPeawcAmhtxFsvY0GLRBOAnTzUWvHvbyLD6SsEp2veJordfh/wSH+NLB7
z9aSP+LaxN7+77cJGOtYrFU1J4MNNfSEnKLXTlJrOOrdvnam5Wk0FRBj+c44kIyxhv0PyWVWGQs1
iro4vCiMn88THX54DonvL5CAh0vPxSrlqqlJHGLGGDcCjNV4jENUPpmuURDTxI7sEk+8OL6MflhG
+WHAEZXx757FdY+SmZub0/0YFkzwKWdlUqA90QUiK85ikWLe1/8HAVXNPwMCLp5+qmU3Gqjtf47q
GRO949sYY8n9wE84ybnQsfn49tOMj4AAyMqv5lNgKRa3ogJbp2Zhv4qz24hvTsd5/Bm3vqUrd6Oj
IJ4aaJKLaIFwzUNzOsAOS3N7XHJJ6xG24MlZ0GdzhRqgqTKjBblri4XjWQQ5fgYdlaBvqqBavVYB
sZ/sK4/TA0prUeQfGYvS7CBwnMEShK6xGDhRxKE03Qqc1eHbPEMvtaMMWQ0r/5CUQZzBRzuS3wqU
BojJRwhyHQI5gPYbjsEdVWl6GJxljK8He/rv0KJta7IK8Ox74OrODEbXrNUXL8AkrmqUGT5IaACw
VzMnQuMU31aSZ5hIQy5xh3xtEnQFh9Eb8CrkTW9bYTkiyaxh8R731sxCYpkNk+lzDCLXVDS6xwcg
odckN60+6G/Rvo68c59uNZJ3WkolsXq8aiplwntmPCmL8SJwPhlWLGchjY+TkSj0oG3IMe8vfede
kQcGrL0b9IzmA+ljEHXyKD8xPunA/ERx53gQyyYGddBtL9bLtptfGKpeuBmA2FdayLaJx8h2jSdG
bW3NtBGWvp3pLVx3TTwFWNTTcX0m4kf53IgcfaUbZHOsmDu+C8yPDANpyzZSiJBo3a39RhnG24VE
ta9ab94rUaqCS8kd3a4axJoVesgdL5417B8m2+XNcW6rddy435wTYc8+w+KPyUd9E9pKFwTP6Du0
nhtJO23wYIWxMTiF5DnAC+qu6yTqbxa0RKkAEO/n0G4KkpH3LFCfywsfh1KGArG/xZpYm7KS9QlO
xB4p52zh4pzhoCRrKKzsFE20Q2SsL2LhX2BkkmDeGI8dlVavi8IenEWV1llN2h8/yXErW0SzBNsd
SEPAwp0BXR8ArAh9gR1m6uBRj+NPd5qqP/hALG9V80fu2aR6PIfTy/3Fi+LTSQCRAWZm0eSML9Ov
8fz1/qr0RkwqThoTfPIwZ2oq4Wpg/Tzrh7eLbhAHSSE86IlDV2z+/B1jRAsgvjYbQ4udi4edp6z+
w8AcqeErqns2QwwkrmueaaEvYr8x8uUwbaLTMK6C3FU8W+JdGx5rPCjIXWOK7FVWsvUHf8n0wheX
6v+4uFL+xp2XS583znpfi2cYtk9CPNID5W6v1S68yekLJN1pHUsL/pOdHGgB2AUX5eNX8m2QVv4j
s+jDv50Ci7WnFLAYwVUMljEGcpjM8H+WuKQ5lGYdnnffzCy1jF8w+dPaBWdYuNv2j8qowmUMAR72
2tiA9e+op2aBeJ5UTcAkJByFFzIvb42wa8DId1dpR9sTQpxG5UUbNrXS9897dgRDllDin7cVAxxb
OZkqhaltZ/7xhM/nr3AL5DvEo5UPeJyruPthfXWaWpSyeq/p3wpLISgnRVSAofusSsCSBR8CGr8q
kK5AIkUndh7PAarQhYpUGdYD8BRKeLaZyuzIeFD7k8kPfQeNZTujcBBXDiOgtGd9awgNBUPA1vOb
P3pHsUZx231mEfM90RyyDEN0Jya9XD9YBTIIxrpBePu3vxeHsnAJ+BzpgVD69fqUIWCdCOikOL52
Gs+IgWPgdyWAEIeMrjdXfoEC7148TWUtj3VEz4Qqa3AqbEYRmKchpck4yp5fiGdIBexsvlQxAuy8
nQUIiHoloobhG6Wxb8uvdEVUkjy7JB96XBgVkZF3kioK7eDrWtkVp0h4C6Mmi3+uLyA4qjLARRUC
MnsbnezKqIiOfUJlmopwWfC9CMJab6PwlCRvIDEaKtL1SwbuILsyfNuIUXCIoMGhKV3OG74jaD/w
73xgIjQMl4fR0ai2Ml5amelGFCA+LBhBcJycW88MRZJmVsvXe7JWzWLH/J1hlBdfdUC5P99/pwMO
HEXE1kD0fqY/5bJvIYZm7l+EKPd2xlfzSx6g4AR68BdxAy4JNhaNPB0yFhIctwBoXIt8gP9ZX+ti
DfsXNuwZVGebCElvxpVM7yrKEbh7QKSXHrkIjfcj7bKBUtm+iBHSoiMJE4Nx3ibkSZrX8DE7+gb/
2uoCUZ6MqB0jg5fxKGkOJTJvlWQ4a4GmnYRqd7AX5PUxMoUYsJdGGn9FW32w5J4aUrwH+ClEINsR
O5L+B5dfwLDX6+dms5NHzOdnA860ksMmWdP4jGbhdXR5wIZAWqXVaC+BvDvFOk0nAMaMAW28YnbZ
NzIeM8btNIAIRAZq4SNZQjlV5LctAP6EVEUPkSQCLEp9nJe6ZbCkiprj3v9ZRmxmJUltybXTOYco
a0sbN0z2J3oxzZVsNXwQl9+Gc1T/NAA+deKfbyvBTyTawJZbgKaremHxtDHBVWhpwnTZxxvP4a3O
dDtlMku03Zel9cznSogv1ABZYXWA70Ud+rtTOwPMJwNXK6nCcNv/1HqSGHCIfExgh60iO4Vz0zNZ
WlRfalx3/fYCxcusjY+q5AHzbuKwH0NODJuNC5gxabuzi5vQ0Hl19nirsgoYh1WAeuj0ml5HMXmm
v3huma7x2475nlxyspm4MwJLmcvzp5egdu/6ecsmYXfjo1WqgPVF16uMrNWo/MQtHj+4JXlvHdCP
lSAN2ew06HoCuk4kfn42C0SZvIL8htVMbfyCGiNnI7e3uWEvuSLPjs5c7qcUculRjPsQjVqLOLmB
iMHFedXtHL0rJxO14eN/zQaDQa0PhbZtPhdXk5e1DPiO0fpR0uHQzwJJWeqeyycq1vo9xAxDs9kE
PKhA9Uj5zLsTGYdBofDsXoVzKgekeeoK7+5PNksMRue66vUArqN+Y+NOqCHNNMIj5QwUDILJ2IJg
1bZs1cfsZwqpFPfthITDjgYXDSiNOY0c0sI8QH6Fb8lKCimM8phWKKPUJplbvF0nkbvkc3yqkOz8
UBWcjdMpyTUwPEhoJ87TSKGyCS1oeuA3OqKzqiOKiBPUwqVqTgH/STLDgzuBqHGH+yKR00n7vdF+
Bq/ibaWysdo38mASqAh5F9wWg8EUHN0RAAlnK0JGTLh3pcDBBXY1UWgNaeO523909VQGZQ4lz8TX
IYQitQgPIP/B7WP033hCkNKKmmxWZh3jvBDeql44ecbKbLAJUY9A4FNBh9NAq6TX8vd1Kswc4FQh
HBdMVh4fluiMNDxUckibvQJLdqwqxjzad/29+1E4ciIa0sUpatd+7AOjHa4J0m8pwzvPLmc0LGpE
j5jWZFEA1d4ESKDIJrwKiFIvckJkYSsLte1aJe8VSYKuDtW/cKyM+vItwEB3gv9CVE3Hcbex7G1i
FmJW8xy70j9Ei9hQaVjCRPtBudnyOUfd0YX7Tf9jtugWV/OXmFnrvAN/NBKwFDA1gJ6Anb2uMe1U
c3OTXu29MILqr8kII7PRWD75CkHWgSM8llE9UXVH78Q9BEw3ajs51y+0j3drXyxzZsPmOszjH2pq
rKg9FAZKmYctu+XzEs4JkL5/a36zf+rFNFqJGQZLMwnUDMlzqFi+raDga8Va86ZY6ORNYzmu3CJN
04D8i8h+g45/LE70ase0ZCZxNx+52x+0cUd94LVN1xSGp1vfAkiR4jBrKj5qfc+sDS+7GfWWw/dx
fScDHC8Su6p6OcRJ1U9nM+qA9MMb4ryHNvykQqe9/0P6xbp++eZEdSz6HJjh2VBM0iWoCZKZ9tPS
s3KHL8NWW1Ev0seEJQaoREZRBN0jnADuZqB2Wlo9sS+dcLiGZ+ZPK1CqjlQqRMYNiG1xY9DpWqtD
9jXRF/Hl2sk82RRi9+uzVrJlcA3aw3vVVH96SrGK+TGMZ3w5M8FErWKW2JEN5RunlqBzg7/DEzgt
lk+XkdtB1ieGsQUmandP88tWP162RfTnGdl08kSX2lK610iAuh/174prjJeVJE2kYh8yy61PAnla
XxTF6wLwicWdwNR8wRABAFk7+JU0MJPcZQ/QQDpCatU6GJtjxdUTqFr7I1PfxZPCxMY9B5gKu16L
C5Wdoi5iBEcmNsjkCrMuNQOkPzAmMiu+slM79vJxmYEQwUXk4ffmzSj7foB+5thjiLpYzy6u+PVm
fio8q8IHNmN0sK98c9Zd/q60MkwVLOtC3Ul6GNx34Xzd1xgcKHXPMb437RmVgtIZkJhKrU92DCf3
HpXJ1NFywVjUF2Ouv3qlKhwT0AB9zxruJzWcFNnN1Ebq+nExDEpsknYNB/juVjESzhFZ9r258Xmm
1OOvtG/BF4+oFEAPK9Kqs8zSFoRWKN+MG89Bb8woCVBASynQCe7TKJZTfwXoeNMilAxb55mMmM2c
KOcHPsidPKsmwjqEUbCPB6yB1m91b/6R+mCad5rNFOB6L2X1SPMDOVJNVxmu82eErgT2oNUtylRB
bPU3QHgtEOxYU4gitG3Y1To1SMX7ISucU+cCY5AIixPKjff2mhlTbA5OBUnwlmX3vq3d+lTs6vMz
zcyHTBRfWhv60rXK4hGfIwcgdSltgWDIAzAsIBGPh+CgaaemAwmcIxrqZlYy6D8WPWF4nOU3QrZp
r8r4s7DXtc3ya2eD0DjQzlfz3teNkTmEY2+gm1NAecEr62bUMtAt1YAPIlQ8jHyfCGPyPUaFAshQ
BySHSehOxwWJN/UWqRLxbyQwqGq6UXP9Ck46YTo8EKs1jMps3Ksxw7CbOK19bVllbcQ9jUJm9oLq
MDryI7uf12UxX2vtzPHi4IFgt9S25kWWJeOzmWJpXJuftDFmuRaJ4tH90cpmIr906UNTiKPHP90c
40u4cBgii9mSCAI8wzYGzHYQXfON2nrwD8rrwRWpTmUt5/e5NJBO5oM3F9cQ16WPoQyYRJ+pJZU0
BwRMvZ1pt2kyqyS8vPZ52zhvIH3dETzQKZLqZQ3nAUOTqEbq9I+OXNQ7jRaAxb29Bs8L23w5Tcsz
GG9qiksVD+exb0p64SZYIKufnB5zmiRQK6mH/TqV6F070kHfUUY/4lN8szbjddwSa1uGf5MQL++n
m8CQHiIN5fLU5Tx83Lkc9T9hRlCXkRJFh0+ThGzlp6v4M/C1s52nOcrkZK1T+QMRrQ11o96c33QF
g2v8TQgNKsr07U5JwTAi6TWQ5VgEnZLu6Ed7nhYkPrp9IjOxDtP3VYtf/iom0XEgh9BfqGwT6Qjv
IU9FX7APLxVtgSpbrwv0zaBalJJsuuK+uiiYzH7bsw2/hZLHbSHwhvqoHC0/lmaoZJKXzowq72W+
0RTKZ4PhvArUGExUP+XFZVqwYCjcRJ+pCoM9uBJL0ls5h9mZxdbx+Pu34N/p+sI/fSyQIp3bEadv
oyf7+0RN8tOUnKLwspTod2xfnk96jJaW6LobOP5oJJcyiACDIosL94VscAp9VU3XkHaIK8G7+Cu8
Ydf4tksCU1s47/B/eVfclwy3g6161PPr+9CVX1QrKAHK69rnDP02PRBBXKiY96VJSrwNxoNKZqY/
qx/OuJJ+89RrLrLDSvpi7/43PsvQ09IarI3OBRu9T75yeOKX2sy30TBv3mN5c76tpKrs2fECM1qv
huD/RdfaF3ZxB+XLMZ/vGM1x2S8DVjqlVL5lxTKqHDkEE8qzsHKYmmuFwChoXFBFrFxL9Vqzx4ho
soYxHIlpuIzozEFSrz/M1NCw/Y5J4Dw7rsporP2mFUVzCqA4Vf+ac+3fKhNF04LAOW1UysdwHMuq
BQPLLc3Vmb6bAZpZZx8I5zsk2BM5rgXrz6IBwSsnijjM4EVdBam8KmSRB+IehycnV2xcUfsJs7Dd
WLTuUnNkRvcujqTO1pkdtNQKiOYKzyDeqzAN97C3xprP/KLSIZD3FDcWUbwnpT7l6rHny8T0Iu8a
Pc8PYB3eY5O2282wu8TiWBKr5KKXdrUR1KF8yfrk9sLUglM9q55/RNzVp7NciyyKSQTIJAWH4VoI
BWd3ld4ZOMPn4KeFenTleQ3a2QESWpxKMVXWNM/eGFdauSTDZNTI2e88eJr3z7NmAb38d9KWt9bm
PiCVwulpVtPyh0no1uA8bSEP2A1tFTfv1WAjTOjAIbKM+VyzB5dvlL5HNhyWQGMQg9FMMM3kD94f
p0XRK7JKB+roY+XRBbFfQIqgHBKn18KZJrFzD7Ozcia4j3Ulq8Mw7suhRIs12T1eYuZqgxC1O2Di
C5xVu1DvsppEXdbOddjwkU4irn0aKKKW+J0DM6yxe2iFa3EHAeAOIRRwRTYXqFPsJcOj5xsihbxi
/Qh805S6IzJxcMsheQcJCUoPxv0pH290SWdYtDRVS1Kp8hDHh+K4oSHjUkUtGQek10YoisS3WvPK
WwW6OejR+Uf0DkQ27vGcbtm7smxPlkjY4L+e0Q4aajcZ5lO5pXCN2tTAgvxLdAjM+T2e1uemLQ4r
LCCl9IAO478u6mVvRMPaLFoT4yOOLY/wmU3HWdtd+xoLGaFnTeAKa11g0ccLWEtaADIU4xlp2a8x
wdQwldYuKlVtapA6RPPrqMEkADAukv9nlEp+Kybpvci8KMLRUP6Rm8751pHcTrQWpUeYRt46tGUh
D16sCQv4EG1EJWXBPNQOmVj3D69iWWvNmvna4Zx9aRRXXm5TCMbBiyR/WwUKsNgAC/LjsykYUcfp
ZaNISvxgrW1A/dtki6Bdh1NfCMRYZuAnMKeShe7if35rnH6+JnqLOEJiibEtTIzgfK5hDdUsdrSY
UUeHaaumVkC6NyiovIR3P9qBFo0Nms+UZCz49Y7/Gi6SdgzfvXxfkwwza0vqxXhMJ/SSBglGUt4W
aXn6nq2tWyCkonGI6H/faL1aDTSbuF1rjwdv0DdP9QAyevBg5J14qGaq0a2s8lZpJ1d+ioo2/rO1
VsW180DTpWOn/itsanvRYxBC7TDYs9J1Rk5oeJuVL7CaG/VANOCQ3eGbcOy9OxvDjYlbq5oVWjAU
RDJ5MoGTpU0bjxW1KchzywZcOTTO4mU53Qc3Ht04PBSjmp4XW/gsLqhqwc0VCA4iroEYmZacTtwk
hPU9CafxH8IeZBtORcnOIe02WKO8Bo2uWQgbJBmNnaLmKburzHLRR3l6BOTIZYREPIFVAOpF8EeS
0RfEVD8Pot6LQylrhm1jQ+SvSBfntwSbHTTCB2UTMkC9Ue3M2O34jht19ZWP7HbpJfqj/Z+BkSm7
aOjPXBaBit4bgG3H8MgAEsVDp+3ZDuCfQiYc9pg3QqVj85EXRZM24SUy7VLYZ0X6OQd8VQGuW0bc
grb00AILtP6V14G9TuWYKSZqX/9BDplxo6koybCQYyRF4DB20sK7UP6n93eiO1LNtqBmlzKbgjJm
Fs/H16oOwMSwlcUgsGS00E2Hpe/FT4UEClWUCUWJ0k8VJabzipuPNnpJ6Si+QbzZqv47uuvnJnxd
q+L1JyWEZfLq9pi5RgRIOX3xEwlhLt81jAM15Mu0+6koNtGgBj2MlQX42/1OdEDf6CAlUlb7J+xB
zSjCNO1W4DgIK/qWAefANQGmSi3QrItGcgVG32mjeNZWJ5js0jMJttr0G9fQDTE+keluhd7xhk/u
Ds32FP/hyQ6KNxwN09hmO/Kq7Awz5LKJzWZZgIJ1pSyao/HayOQZKpgf5JYsKwLVaPBOWCcxYY8q
UlZu2ImtvXWTCQm+l8I59xraew3cpbqqKiYQlBTGPd/3MWSGllbSiLQFuZGWCm0a4Xhh6qgmgvSV
b5FMF0c27fNYRH1EizraM+yCny4AbTEdjoQrDxFIhyFDC4wHpjcr2I85pw1qojz87UQ/IAOjgYo4
PtODf7O5oXE4xfJ1yBccAlpe4lxEmQMtAjYN5oEQhhb4Kfm0jrxshgp/r+9CeMe2jLmFMnbs8HTd
2vefLvkmzIO9fmqFIW1N3zfwGscMjW/KTkPfB9CDe0upr1pRxzmIYldOGkK3mzaNQHWtZKLCAhA5
3NWQzRkrzZeImgbUc2+9yCHb5lqS29RebTM3ZbCj08nOdmkQR4fazBPEOicsiwf8OPbFC8zMNamy
KQzYW5T/Z2DYh/2XQLIj4eaggd2IJ4/N8zg8Ajuq+a2yE8e9YbcQ9eC+GvFrzImBjooB/AEzonlk
GsoRYKc4DnHOmeEnNBuow/XZwMn+EJVVCWayZKYHoLevfAFV6x4i9zDpn7Dtg6KwWF1lSavIcHoQ
7hJQAjTIA+0bu9xfH8VHX01nq4Rnd5GEwTqswJiQOeHTLYeL5bm0YiqzMx6RalWkeM0sPIaUTjXy
iC12aRoqJlEzr0EFkVQnHZDFcmx8XkiVcC6mGv2ZBF+6X/U1yncULxB5idmXdov1yTEaMeFzGFpj
HWUei/3YhSjYy4wrTGUbTPmgRTDLJpLpJ7Q4jspJwC0uQZYDsBnEYXjRWszaC/BhLrztLip2XJi8
eAgpn9fsDyDve/p6uPF/LN2OUrSdV86HtkjUcZ4RreFJt5qe5yQtjbSu7PI1Uu0KxNDuPyAV9aeV
7d6Kidv/cDIavrGslNmMAee1gLfZm0RPaJk08vU/l2y3CnaiX9TiPhDpYlErNlT3FwNTYH9dDbCP
PN/J735j4wro4ZMMdCaPNQlOkI4vReYb42fjZu3ZyNrpadg6eZ/JU9M6yBz7iTODMk6lSGLq9TER
cb1dUJu2yRdRSPWxLooWibDX6fXytgibZIKRNkBw9G3Qz6UBiO5PcXLnEhT4KeIO4eZtvzjaBhhy
b4HkqUSL3YAoroUoxXp3fSo1PtuX0b7YwsA5GI/gL3hbKPkYlhz1vqwoS4V33BcomG3bz/7pIpFp
4geWjb+z7QXbj9jjRVc+eO3EOmxKuQmM7eP9yAJCc9sAvBrG4Tz6FOjrQ9HGEyEPXRQOKvFv5a4w
F0JyExNYXGLAw9LfrvYVFXBVEHksdkVloHBSvgq5ZK4H/iaLlaNUAuEWzhCCUT7nepm2mpPO7F7M
KzIY0mdD1g7lI42lJWeyEpVY8ITOHvSAH15Tr09pupzdWiwU9L8FkcxXy6q+uEospUEM6qcD/ShW
EIf21KP5Y0WzJXZQt4XcOPJXkD/VcgH7YF6keH6D6EABAMxUtYL010cl4nOsN3zynagq2K2PHD7K
AnSqjB/S81VZYPxqITIdYfCte2Yr5OeUKi5yK7x51FhCFL4LTKmzQxMtQtOaZl0tu00ZeRJKne9l
IbvsaFmoK9ME/M/68Ju4s8ipdNYK2lO1Zds0KIPK/s7ZuNaASJZ6xZ1oNEZFhtZw2YgBcMm+b/zu
5//bdehwyxw8lYNea8oUcEy5MnhCmIUyKmoJXH51IqsBX6f6oVJMf/8NAYj5UsfW+BPClL0u6wjR
rTI60GnO/w9XYU1zPEW3SU/Clm2CpVjhHXcM1SW0CBLH4TVuLwZxaqRKdCcr1foywJDIT0Kn3t77
A5gM9l+n8tOD/cEWh5gNQof7imAo3mdnJ19KM6GdlsMPZK37Ucqg6Id5YKUpQrnWZWTLpA8jlgRS
IMBmAO8+ufXMhmIa9Homb4TohtxdtFuaZwSMQLx7pxnHicJ9e1flIjqRVblci+dAw6R/T99JP+BQ
eNF48SKo1HcQzXqOpT/33XLHJw7Ii9afouDjMStLGha9hCeWmp0PnJci1WRiiQ1ipae0z6aR4nUq
5NW059ZYNng9NXssxrAqLRpObd408NqQhukAqggOKQDcyr+Qm2ftvP9kBWQB6HfB1e2tKS7SXU3L
lyGT2ynwwmjREqMKWI3UO50w1snOdQSh8TEYTa2AV/fXA6gUofs6XWYaqxurY/P3BjttgY7JncZI
+LOuKfF5QqEhlLU8otWPtVsntk1Xxz+DQGn26Ud0p2yAlnlg+B3sfC9QejXcF+QkTwzIZ3HKOA9f
tBaJVlwA9wEGeWcjRGwyUMRCR3FTFYOnzssrdBTzeXrYuc9ie4NvYLU33t7K8Iy/vGk7jjfMpIiz
GJh/wkffbQ0+Dcuuo+87/Ng0MfjgqVJWkEyZf9V7uwMkKuNGEyX3L8hOhKv1xrvFu4vvXs/g/DIi
7PpJYm/hYI1RmwizeUxtTct1FjPtV3XgrG5CG70JKa8nijk9Nar3bWk9Bi+4ZZLLwKTqWi7o6ewi
d4sRWqc9zGfYD4yolZ04y6sRhzkx2Iya/gxNJmWbjZwWKuA+1MA9ziODUf3Wi/0t98xJLUTMCb/X
LPsNDgxPmAiZtawAXyuMeCuJq5Ftgz8z5noZi3wts0IPcWXHnOGNhdF0ppIBBx9UpUUMoLg6/s8s
J3HnZm16XwFbGQls25+PyirqlNiHqIR+tSDmHLxA1bbrc5NL9PvRaUCi+MZWubJkjFoWFQFSTYBf
z0z83EYiNmfwo7gxJPyQWMic1xhoc6k48JInNZvg3u6hYawOxX/1iAgjq7wkKAO8tsDDMm7/f5R9
rDntGCcMGd2VN0EGTnl/5kwX4j8ECa2bRAqcPRjvGu99HoHw/bN1vdz6m2dwSqQbP96zuwptpLYA
GlqNgYmrTDO4IebGGNDkyOAnRrOn/Rl7oT4bsINkESIur6zuw0AoXl9PaaUTbxZCUJX36otGxJq9
KwCMI6s6yfzXZPWQh6dq0avSqs3glOKXo+vEQyFrcDOtsJNzr464LNc1fy3kbezFFm97TKLYVyKm
USrLRfjtOK7TNm8QEk2kvgyh8R9KcXuUpu9hiPb7gIu4NmX94hBmFlOUmWo4GE02Mu43eGBZMc+0
DZeL8N+zd6xq4SD5YNCEjzEwUobTdrBSoeteV52J9TtefXC1APaqE5MW+0fouFm9Zus6qFz8mP7S
Rt/zLE562kiOKPe8ix1kc/KyfwFzeI6R5UhoYeXKoc3W7VhfdX7CtWlcsGUj7C+sCwp6VAN0zcdF
ZDV0Ik6ap9BZiv9Atx1CCKYfyTK4SYQ7NKPTd4SdVkiVH9o2HKi5f2o2r/85xfT95T63LpETu8lQ
n0weMw+hup20RPbaaQqF1/RCFv9spYB8C9bi+ptqxvQvNfG07/Gq13tr2FmNPxYZQ5JMg/hrYmJ3
fLOvdnA47+iweD2R+w6RvL8LMC+L6RTWM1rQfi0ndhepnY6h+EshFFSbjH8qjhAzP125PX0afsIj
7ls6nY9Zw4Y6uKdsjgv55YVF45gOip44xbjiUytLGH6iqae2m4YgZs2FN54YMFSyhugA5qYzMR0h
kF51gbRVLuiNcLuNOjMCDbveN02e6XKXKF7E0nNuXRYluNarPsgXPusoucIHzd+ePK8VgjYZXG0o
0EUU6K8ar2MHbh3d5Ya7taK02At5J7u0LuEQJ7yLjEgvlluS/JsSQoougS1B96U1S8s4n0FNUbWU
rj6CklwgET41TN04r3ujG//Qc01r5LjQEZqjtNuqHT9MIduXhZYjclGMFiEVFgSAhpqxEkff6zjJ
EpxypkoZLrc8Uo6K4Sy4XLGUoRrdEu3a+h4Ssdv0ol//orgf2Tl+Nu7sbb8rF7jVrQCAukiz3LZY
sYmeVqqe1aDmqSmTxamp6Xb+LkTIFdiHZJt40uyoQrOnUDNI90n+P5IlfFaXdOf4XgWVfYCVOfM6
5wXOM9ufLR/rdyzS11Az6D6uDFLeA/KjpDcDGvl5dLtRLGuotVjZz5GxK3TrKcd9ND9dc5RWJ9uq
0jMg7kOppO2i65IHc183cVqHOq7aoLP2AkP+kVuIlD7ENrt1YtMQ5YeDxpjYm5z7yDjgwwLumHfL
mBc6/Fo95OgNnjFikrR1zyqx0Ney0E3ICH4hUcxz31vubCIj/P53FPFFD+3YWEwhsv80pnTdBEub
k91kEwD8CxptCICdr6/SLhzYPaWMhk9mj4o+tRDL5emZf9WdyypPaQbO0PnGgzVGj1+Nde/Jh2gq
ZrdJb20Ql1LJgHt+s9zD4bCCfxK8Ej9Lg3ykh4mizp2rlAjz3E2404I048aNWTf8afP+R5yp70ml
ShIQqFl3IqqN1wdlX4pj1VxAwZ50y1wwg6YDKMtJODARBIYlmg2B8woCqRWxsVCEFNTFszOvnDI9
o6ddFoAalYOQSU+w0o3aBLWrAl3vqmPs4Q1rODG2VNTZPk6E8zk+jdMTTmDipYOGds/pvlhNG70N
Xo3SPeBYP+xZqmExTiIiR1830v6w9RDTDkjTw0Cv4WRaw3e32hteF+EzCneRQSTn7s1LWIEdXTgg
TgOfsZts4uXYy3uMlVur7XVpWcHd1c2+IdUfX/ZI4ZHGYQ17nEnJPHBXP6ZFrryfsf++2t/OWA+N
QZA6jOKT8ZjHYwNhafwe2mDIDmBPtv9przUCtLW2pyc5RL/xfo5cwiWn4n+3S1dwqt9ipJxLeqMe
EqUPbdInhdIJt4gLbJacTtcN5k+7FTOuS/yYF0qtKVJIStLV9ZPKx/RdY9aCTI1xL0UfUy+ugxUR
wHSh3n7GqZggG0JYlZ0NEHbnbGoBnlw22O+i0vyLLjSfD+YMAAXHKb5hcziarCvpH1lMv2K1HuCK
lBHmDHSS/i1bJNrpPJCSVPGJjgMx2jnQDzpEx7LT+6Wy1vKnQHug1UbWmGUZUKrF2drIsZst27QB
k34CzRzcevA6TiLL/W91WNxepUHn4cu6ZZuXjvyiT1XgSPQPjU6ooC+cBCHdcQWmABz9yttkUAZc
O4XkpP6CLO4Zn56af/AtthiGO/v1O+m7m2+3rVeHsub0vDx0LPIWfqf0j40DbsqwtuPSVsyUW1x7
FSGlbWIzqqCBUyre1gsDHE3zqWz0/NyXBFt+99vTN6IUn/KycYANt+zwLaBq2a4rJpBR1QEMpwpp
bQEJ3Uep9U9PFFkLR0FEkzUWtu0mM6ytZ8zH2zTz1BIdOUKoTO9aMjrBCkdpy01WOut/TWdOa03w
oMYDhb4/xBxD34+SCXvFFkZ8jzuLWJQE/RERuRosTvHdRneNlBV+jRprEDiJh4Sj06H1zg80L+jj
xCyi/0WnLHmKXPA5RGSH2LlRR7OFkXBVz46kTsIpJCmHsUMR/oKwn5u+10TMAzvrADOHmKTfgGZY
ykIkoe2dcl8sEhg8vo03HxM4JrQQbT5ctZWqgY1rqHx2sropBKKwFnoOcYDZ/swORqwp6C5KGIUD
PTkv/S92f9J3eECZmUE+0gJd365QLNY17aQiqz8N3Lx15PfTcA3ZdjnaButiD0Ayx3xH7q10Xq9D
Xm6rW5O3m1M+k5zaupdKVu3/59yLEdD8fMCURfza1snzm41KAvO/L+yGwKWqmIAJtcQyqsfdlEIO
PQoQu8gZ1hVx//IKBMgKJHfwR32y+XdWZBObHr+uQKDV3ouw/F3oLsLcRjFmKyzwXnFYoRAioOmq
tLAd3Wmq1j5RMasU9e/3+SlYhYvZGg30hlbL9rg9txYuIKO+DkN/bohrhHQaEK44vmEns9Xy5mCv
xGSp6umbXvwGRqrIQWLKyEAIt0YdU3K876p7ywAeEb0vd7CXwph5R+m1iW/zLgw8qbjLHMKZ6hAZ
Q6tV3vXJfc3DGLS9xH0GqEDASofFQ76qTRvKrCuKPCzcNXmCiini5pjpjJHFMutEcfQW8P64mkUu
6jVjRILYLT9oTx0wUrokXOhtUYq1w97JJ0w7H9XgQe3wYnp1sLLl0akUfTWYvGl2Y9ae71AoT8uE
sGZUEwpCd5OkA8/Bm1oJN9eVWaASLznAU+z0wkKMOdSIxbKZV63xLVDYCfP1tI0dVTm25MNC/oFL
TUR9r6SPj/RpROgrQGU/srYccLfESHVb5Isd8+pcYZ/+pqTDRhckHAjNu7x27ZDsQPGvoic43JeF
uI2qqtCfcvNrV0Fq7EqRfI3dJfkqsY+X3SvCcP65Wn2mv082r1jXmWVgrJTTAdVSwssz15F4m7Jg
Liz4GjYeL4kXTpqlzaAqPj/9r1h4Bors2GFEB82VUr3GEbmA/EanwrVEgM6EGwMplR+jW2gXT08l
frPBAHERz0O4YGwuNUtQR6jbfDIu4Ki7CXreoAPwpKwPMZzQSzgw7REHs54BIvvC34L911cOAxUw
DvO7/mIxIX71cLK35ywDNjA9UROQs5Owt+KK2TqNuHV61ikbTdDrUQoF3iGSs/F8ICj5XMXawixe
+SxfSaWlS9GqOG7O8xFbgeNL2zsuOZVW2S0P1xg1hSxf6kVnhLnYbQiQdtDfvoHw3svHhXsYk7L7
1G6giBc11rK3sfQwI7nGAW4q+CPZq2fngEwcUdj8akXwnKAuhOh/FkO6Sv+HR+DNZftBnshRIj2q
TGPN7RgqaN0yKFiMKpvFX4+Aav43XLcYzNQhYxKOhM6ZT3X5FTwVhOq2vZ068wSfIzFcFQELCrbR
6AVnsaNUnV4TAZRZ6AVZPTygz/AiYkWj5ACsQ7ic7GUTF9dkAMChrLh6AigjxsndQjcTTDNzHAWk
N3M9dszSWtYi+ms6vqFqOuVHuTQw61oAIrrsqYdhK/6DnIylkvaabDcME+A6VevacFeO7zTqBDUD
306OFESnDBsfHIuA2QpMiX6eUqmWYxJNzakG4lZzHTEkZ9y33+X4plgee+txGms0Px1zuwbVBbNs
DbRVyf9qlZU1LfVOMKCauUTGQzIQPue76vJCHtUQ5zHBoEThGGqZ25qqA+VoE447PoPqHSVNpUZV
8fArsdbeg2Jev4IJmtbmsNfUS+2m+DhaL0/0JC275rc6Qr8B1uB2DIVRcdNH4BNvvgwNod1rfMyw
j5aofTnhkUyEVDsJsjme0M1Ng52QXTo37Huew4KfkCUT1hn+oiTiMGwz/FVLaBq/K718rfUx/KO2
jP03LLR5vnjHtAX+zrp7SMH4UIvuXmai8MUuPcZFcOum2OLdDtbCw1AQjTjtWCtAvTrAqRuWQW3h
pcSE5Nnfnc4uWzr333ExRWeGU1LWjqEvA2vhvPYXmFLPHtVq+zx3wwlQQsURCDD//ThBtXly0Ke9
JLY8hoOjEj5Ot7GNSUsdmqiAb/L2/zMAlbeIshR2UPawn0m3/uJ1UsrfXtJmX+aSMPauzwP3O6u0
ff2S31efDcpSS+I5BaDWh7JwdoB2QldOf4EdLXy5pYWVQxz+oI6VRHzyXAtlmDs6WCgVG38DZcTo
NkVeZj0fIbUoPSBKgR1cFkc3U2xKwHp9jQ5lmNDOurEsZ4qH7JAhLBDb2aAmaws1VVgU4rkky4+Z
ms2a80R5mwPdF5A7m2cgrT33CRiCDSyxnQRpd9G22JHUfSEleXo4tf1DmsSC1yFWkMSmJ3tELFqB
LDMuIOqMBz02yiWqM1XO6UmlO6K2FHHsQVpWCUafOVPDwG8w3IxqTpkhvV4TPzaKN8fd1hLhSlBc
6dhPLSlpPIAb9nptEKoxI8yGzJQRvP4U9Hu6ykWYwRuMx7SVOYHiUEo5T3XsLE0Vq7nPqBZl+cd/
h+tZQGYmZNqAnJeWciOOGJnUb28UCUDZLiU7+KMBIug0dWuXYvWNx99SWEcf2rVTIwtfVFvoWF3m
6SNqdL+CvoG1LKYT8pJ5mc93rveJiL2YmX1wY7Bkp5ytMPJFO6YmUdyXl29YvaoycXKd+K3D1V4H
bO8wWoddKNQ6d/vVotkEEqIpO1duqTgABIV5kuHbYgDA6mzderT/hxwrtmVXWT798+PIfd08+NiC
GV360mlR95Kf+zsx+a4bbs/Z2U34z9PxAMMcYsQ5s1i9A89wbFrV4jZ/Ih0Vwn5AVwilkTgXpHnn
82Yfvq7zCJA2pQsJ2w3P1umPpEAqp3LpUmkFvNWLVcOVGQliH9nVQyQLSR6fViyMqAY/JBXCZlRS
KXMQApObR5rSWvCFJX0D1pFmt8xu0I1woGOG85Rul6j/QRu1lbTXk6+lVo4f+4PjKR8Ze0DdC1Be
UIXtMcYO/vTAUXYcD9zSP9WhRdQ2eG1yxSJgGuxP5E2QezkkOBaThhUKg2zOzGbLVc8iLc7eJw3y
bL+pkTV4ezcqAt0NOY44cdkt5VHAcdUXfnPbU3ZJ3qRevvwt2acbO81ZMq8bRE7clLspthi4uhSj
iU+SfSSnVUfBq/Kbf4XYQjodthVApLtB4J0DgAH2caf/Qc3ZguWnbcshrJgx5/bS88DCKW5/Adxq
rbl3TByzVjNjhXMteuMdStaNxpe84zY2Oyf3DtFLOcFVjJEJr+Ku42P5YXrIHnoBYHmG6jHpKAIV
o7zGaYG5AVOBP2f/+okOHoBVNKUu3YXDGx+8MSmk+fer+XTKc5l1MWiIw7BOB/gnIfBsEX6lyNzX
RfyPByDva12Ap3O3GyWuWT0TzCV/xAdOjrDUBnmgNBY5iwaMKQCy72P2W8p2PByFCkr7OH0qFMZV
ggaYR3Y54tHuHwk7eCR0cl8iYNoWoMY+m5SE78/Ky3tYlQ5G+bbl9cGZSSPSAPKFBq425b81ky+Z
/y9uTu6sjI6pQHCZK3/Okw3mXQB+zPQDvxNzbBJPVTYS24sUKzcWX0sUC8/P5lwbWjMFMiPdQHhj
BCWJhRO+iw89c/Kiin72DgJiNQTGSV0DoKpNdUJoUzppHQ7wm9Sn/5Bhdiy/X7jS1hj1Uffg8WNb
PMhonA7oLQfgD4b+CgX62x7dEsMI117zNmTvKKDoKvAd+R9NnVpHK7/ZDa/HcIXoUVa8XoAE+IPB
+S09mKK7IKhoSSLbxGgCAXeZ9aBfcWnwQPta76vykZd3/iwKubO0+zD/aBXS0dNa+ODiYd5SOBOb
Utb5VaCSrf9vxL6MvNc+kPjmlP3FWvhErp/Fz5mhXgmXU1YWCQA3fRLWDiBqMm561Glo07elsIMt
lTkoz0ErhScTVVUfpXzVpYrYjoUJXFrn3LpMlXXSOxFRsErvnwPtrd4TXRl18a34CWltj36As7Fz
5taghUmqZoxvlVR64UbSHtEoInB8OPOhNYAGD8wwbvgIo29StC74HTRaP5E8/+UErjZ/b3BKv4yU
Jvirbe5Q8cVVPFpx9x2ARZyFZbabe85qjXovGunksP7xt2HyildDkz2+G9WBjcVYQAIEfTnVoy0R
npjsoXsMpk/r9ZdZhaXbvvRm/BN6uhzc4c+pmuNuBAcRGDXGPmXPuRwSsWZUTlVfS5N1wZMFxfMn
29A4zIXnS3uKf5/gNCj3VQSly3jUn7d+JPOcKwNFlT7mvmQTY4fRWC8r8R92Iehu+bwUm5/I9o7C
5GBDvL7hAO/TMPanz6ngZmXcT7ys6Zh/TXxG34LUyDeRnxrUszwDcyub3MwsAuRsvNaEftG7l7Dx
UrSKo8hKfKC2NjKEjH6+cPSvJvVMrn5HLZnn9lciP6jWQA8IJCq1O18RbppvuyWeS5QGrrPXCZ2t
cLopL4ULLSMzJneqysS2t4mO6++8RrvkLSc9+5ui4my4QDR0WSIEUSJGZ3KHC0B7Lf6ropvK0eCj
WNLOoY1kamiGDiG47E5wlgAJs9ms8Cx8XMKjeCO77hURQMVb5a+OUryj9Rh2IrvqCnXAoJtv/eJg
yAqTHNlHJjWPfkFohkJv2gj0IxVJb3eb956VdOHgn+cye48vTFb5MEtgm09WYcU1YoSuCQJO0QiH
hSS3SjdPMYhGW6KUqh5dqnXYqc9JxE5qcYCow3cQcoy2+D3HKKZpPYkw8oU/ORLnNJOsuVYNUvVN
nCpMvxRwVGsV4kv76sf9qrkda6leKOWNTQ2mgggLJvR1RelCiZPnSrMgasSukzureH/laUDlv2mW
e7FS+KY5S5WAQ5IErYwinmk9f1bGW9QleYksv7XVUqSFvy8apJtQOTiDneeCfzJTbTjbf5BujS6i
PkkmUPSpIX1Urw7rtSRrGqzxvA5//c7/NZGYIr16FZ3KnPYAKaZ0tRJinymdcRHQ63N7kbY9LIvU
8JO3Kp1vE7A+yTAnbfTw40DOoipJU5P5FtE0Rs2QIBT30cO4URpQIRh2QEomgbTx7l/0jsENbBXi
OrYKEurK9dBQHJlYnVNjn88x5+yM3tsCKu5l/5933M5CklB87SnicMIBJdnvRCBfS1o82+1vHGX/
5Q2W8AghlxC/1cCQWuEoKUVJNg/LxjOgPm7Z+/z4f6TJlURRbJvW7Ag6mNrYtxk8Tw7AcEq35ygN
f9/AVUYwRh5foU2MSTKmVNeF/Rilty0iCgtNN4ocTUNVppPM6Qu9gyVbLfsHoe95H6n2mBncokyx
J/HCw+zPr8m3/B6mzfv2Sf1KCmFxylwpH8liJxSeKtat/EJ1bC861HuHaTM98tf/QgDgixCTRH8e
Gh+lDgBuMNtTMSlaJHiwSuRi9ndgcD7gy6fWWtNdm1mveAtFB3qCN3dZDNbX9qQDQfG4xdzOaBCF
qVoYCIlVw13QtcqitjjQzLnmRjz7c6t6HwOpO+jSlJHVCs5W/oNiGhF4AjoPQQXdcHHfpiMez8Wl
6us6m1rqPrUpk5xGdli8wnY4M2HbQ9JZJH/oCMNvYkpAxFhBdYFIdz8RScIeo/cAjhU4Bdc5H3ih
8eaZPPYz4RISu7o+vigoA1P7OGAbdKIR4xaQXKgEBRYTmDZXgrdxCv9OdmyfCAJmdhffJIxuyBN+
3c7SfM1JVYtaKSHxHUVjM6NE1vDTrv2CDjYLeaNNhI7V4BXuNtDpdaKOzSeMg2Ti5g61hwhjyFE9
8Vr0la7t2Ri0xc3aa5clt1cp/csNhKIawZYUZgk7VC2U13Gh7v5xj+KHsfOIXCguZqXdDWMBqaXh
tymYGN549DMF5eJ9D4J/w/dryw0GEVlY05+g85/sGhLhcarWaINKSXjhVm23xq2KNQCR3rDXbY6P
ANli5m1OzSSQV7AInm36LwmoawbG343isNBD/07WHH8uq8gCsUPG9GPw8Ja8OrGFwcxwBNALWEpW
FPYU1wEH2S/RbO8cvpDKVJbtqyj0r5/TfW7IVzspoillTlOqoBYsI4QVk7tNv0QThhkOYf5Dl06M
yJxTLhRBaWt/F/rpPML+Np/Mqw8JpbMAploOZ7gsg+ayoIA7XYxqxNgZtK3u8xhTIPxNWEqP8nNi
KGiGXHJwELOdI8orkb36l2k0VPbC0m/jabYk1sMgZ5JZ1WxnGsSDskUsYEFUcHWWbAt8oIRue++8
jCCo9KWxNihcRwvMUrlnrFwaWBKv9W622nPDJgZj7QRVLJn6gD1lLTWiKnefczJwTFUGnNKod8O0
NTnfOomyXVvguaTNcJZdRjWnnyyJ/pb23xCdyjh0CzSClSW1JnDWyhUDNF2F36ACvaXmToFqhZED
v3lXw1dQRw54d1wchjXRTj/cFp93BnEv3x0LpyJdKTK/GexVwLRQQoHfVN+oa8QA25tYHBcunfZ2
VZUDL2BBbCmRPIMJNpJ2hyYYeEFgNkzTyYxhZ+j/9NYSA3VSFUPR0HSuNru0un9iAf6nn5sSac1S
Vbjovx08+jHD+qSy3Bs+fr25SfODhsckxMcokOiWROrVEeYJ1VCfV1skA2jRz3dUuf2JZSrHlhRm
M2Gnnn5Pq/nLRBrpzeLhC9CrLfmtAc9C9InyjBUSX4f9vsnYfu3yTwg3udjaG0i6/U02Ns4LwZd6
kOm/JrrDhKr2OhMI+CYANsMa8uKXgU1QZBJH5JRlPhb4OF/gMPPFHoCO0Tl/TJO5LjivRZhoGLxV
aQdJQYT1hIi31qEoxXkVSKc3R2nGA7mu2ey1LDd8sgs9GsMrye0es+a8qh7H9wRCxrfF01wcmqqS
NCktgZIVdkZmB9WrPv4riPiLhmFcKe7n2OXRODKkF4tA1qzOWXOfg5DGWZjxUMGg5cfLy5SjWRc8
dwVUt0cWbcb5ww8KjBuQk4B0SGmZpzCdfyIDS3ikv5Mm5p0UoESd204UIzSKuZRcfYZvxofMbdzd
YZH8/z3Kl8NY9AkJ/VwBSSAjq6Td3PKcN1d2CmebVfQUOiA1pJTSFHsnRx1dEIqqS7LInBrbd2nh
cK/hut1npFfDiArbzOrAPh3fSgfMrM9tFPxRYKKlVpHMk/2+huvYCMd0BpesWTzzicL6vyKC+Qo+
GVptX5lYxpw9H/n26PlB5VS8wCzqmjavOaNm0ylyMqjeErol3R12W2VT33xgB1cc3AOQG9NkgU8Z
6itwi4dx4/y55CcLu2gZVFIDuRv6abUf7NANX5xiUowLsDnkHLn4itFhycRONQtbQVnb90iID4RC
8hLe1EtoV1N8cuJMQ5K6yEpnBEdZ4xDVHPN+4htOdfWR28JObFWPiU+whKkvXkyNXjSiPpFn7S4Q
FqIDFWFjXa7dgaJHQtn31Aivb942S4Ie6LMesBV2fmr3F54/ZB24OqXCT71fzNntGNj7kywnDJw9
mhBjDZjDrJ2yCJ1GfRqZTFeVBK40+H9TMBbErCLKlHSXA17iOryQ14RDq7hB2nhjox7uy7J6k0Ct
L+KZX3l6I0UI9sHqU8emYiFSzWW2BgbCQuaCDJzR94uPjJr9wTZby9CZRFHHO+4bbggTbNRk9yx2
eWb/m6US6Xylj4FWCDH3+vOsGNtbhbObMa6/JibV9/dIobwsy7zyXtNmpz4F9p60u6uyZ5fvjCQ2
V3tqdvatdtgp5OMEc/qrqB2zFvDaVNKCwqMCfkXGFQTPoviEIXnTfv651mQtSWQcVyaft/CHSLr7
ZiFGOcy4tQwh1ne0hcDZdTVd7cslrkVFgJDX5PXQ0l7zb6uTSmUSvNzG635JqwSi9zeEhXGwL5mE
edC2aKzQ/ciSlLq0ve0Qrp4cdwi3QwpP/KSq0Eyv8ZB7cyqOlophamv4QEKEWA19VN2FjH7sPYmv
1MquXxb+vAbqcDF6aLDoEo7uqnL/g7tHW848s/2gWnyUEVgoBiygnUAJkCp7Aqcu5lwkB5Y3AlXH
mv7q/FsE/QIwEUZvhuwzTugt8XuynbLoxM8HUqof8IjXGf/eWrkWUmpO0SsMKTr3r/m9CfLzqDdD
RpqcR4Ifbx3OTvOGIk3ru4gmiJmvDaz2wF8g9FLluN7hNqy312Cxfmkkgi6Ihq2+qrvFi8Q7tITN
dVecL8lugqsJlb8zm90Jko2ZIaPnhtb6G2WefO0HpJyCGL86eLVKtJ4chXFD+ZyZuybrZl3eiQFw
Clgg1EswVo3l6ffJl50r1JC2digjZ8tQVKr7W6kEExTHJS6u9cnYLCjFtPXnk/GkwEOF75y0vhHQ
W/3VWJQKloF+tAzlSUFu8PWGkjTayHZNSiPLZkJSEWrggLYGSXekRanlHb6SVjZgCzE21U3vLSYV
3U3TvN+9Jaq0bKOPcR/3pJd573L+fPNVROTPlh+fdTpr/Rt3q8Eft2K+zTu/vheaCTKch9JtpryY
ZrAR2oeCry5cca2xVpPzE7x+F4P1v6BAciOJh7eKHOEJ59xBPjclDY0aqTrxoOoRidruA0Tdxkr4
IWLVFR6wfXVIKgwUBfyHDFRHj8d7XfpN+dKzN5D5BmMUXr9gCtKOTZQzACUSc1iteCZu0RZlw4+E
DD4cj+FnSxLb83dNYAcFZQkG2hBQNTBnbS2Q81AlrGB3nXMTqY6qt7NI7FhgG9kSn2qOJcltVNvD
EtxvSPaEdQS8cHLr16sZ0E+LWv2gfZ04mnfHuj4GT70QiQ740wQgq+kZF9YlZlpyPeHLIO8kKJUe
GT+UIesiv7+5OfWOTLPiHrPIPY/DfPM6WstSn/qWI1eSpnQwlN7aBVOPi1LYRmr6otaELqgeNo8Q
42zMABNdg3vOnpitBY447T8KM9c1zS2lXj7AaUJbm1wp3s85DxqrrDlfRg18bWjT+Vyi8dHURTH2
5Cd58d9j7sJogA3ybqb/FvQr0zam/MIsba/NHKZeuIMjfYJGsfXFHf9bHikdZbaVmRTwC7B+o04t
xJNrbbv5JSGlWU6/63Rb9v84rWKX8ih5bJ0/TobMW+jQJx/lDMVQhnJNKN2M4eOndNNbR824VTNn
UKaqh6v9ZwjTkTT6D75kv/eTnD246Y58qqWyOq4+3q9uhtplNQpMfJ6KjNdzCTPbeBzd2jG6v7L5
KcNV+hIQpa07FVklHFFx/2XRwf/k29s9E8UBZKZoTXw4N9dFdq+4dKWovs6kXyoyZPYLBwt4HKA4
bK8jePbtUBTD/pGFwRO6s8xte04TPo1afvIAGNtC4mgvYU7okSqSPCKTKjhvbKPgPz/iMrMYFE+m
+cHfQm6CNe4B5dFcZrNVoaXpIc9JRgH8KsYupxTKDxWJzaJVBy7kRzdqSXdOUOEZjv11takqtVjF
Tn6zLS/D7xzYZBtLUymZSybBx/r531uF9+PSkAmCj0f5SXoP6i9ImxW7jG2FahPO3CgpGL5hsGje
GfgSNN8XfXCMII46/2zpvQ2COxvwFlBSQOy1M4qN5bkjZI1xV57gywivgkYjiN5AgtYVhM418gPL
IvYtMEPq6NCQqYWGmj+fFTR609fymEQtsHoCNMHiztyozZXyvsYEEEx1XgGtIiNvBQhthbcLV6oe
IYfoB/lxG5WoVm4f5et0kRMYx5tKxTpogukRf3/KCqP+I4uveHOBrfTsOaMTYQakkZRBfrwXZuv4
0v8n3/xCSeLyIFmGQlHAOb6UjhQ2TiH/SOX0lJbW99LVbggvHIidPK4SS+8Up4c/HARyg5UvgBOg
H4VsA3S3ZdVVOF4gBMK+fGNQPodI1Yy7uD6yZDqWrHx8BCD/7CJQiACQxsl9+FLEcYvaSW/JtIGV
s3Fs3x3uG3hYrCgAuyDnEzH17v67btcuOLEteZqo6yL4Mon2r9dG85E74nSlvfiyRpcgqaRLd6Gj
CPGUkv6IYWTBso3u5frD3HjHjq8rAu8YsUapoJJ+7CITfLbsLlmlJOWcvvsEzuoI6cTRgoufwp2N
xPqvy6gp0wHoX93sd1/WP70LJMViGgIGU2PbFawkEJY17yt2qjSCbp1Dr6ZXbwqXweGcdnY90a4G
mFm72g+RBzzC9Ok4aQihSY5I8P8mMTzUkNFESR+WRZOQoFjMr60y9eH43Ph3yXj99L0Mc616VFEe
Z3VAOEQTaOXJDKWhUp0MCQeQyK6XhjhalfH/rGl9aPeQEX9S9oohPu8EPRY+i2BXqTPXI2Tq5nNW
bLrewI/9PGOsY6lg8r6aY58NTIWZvCYpcSCRf8iA9E6g6fmB/Nhv3urj2cKhNo+7BTa22eRULKEL
z+1AG7YBTN3RlwriXqDOUMU/aY+xOaBr56c1Z/E4RaHa0pbpOQNfoDE6MjOvlPyhAWsKOruf2AnH
HZMDsPkCrNU1KiAMs3EGl0N6SQgCBLAnwtez6LtFy0cyMKp49aiCMRUfn7NlzZ91a0Z0oINJD31e
v+8nypDyYo8it7DKDn18EY4/pI6ITRnZCi7rXBKKJ/adg96WJstvn3N5Cu4z/KKRWR5L4ynSz1de
f9gHbW2yjW7J2a8ramKdpE6zA4Go1V9zU9I0WUIKXY5igiJBQipiYM8JNZrtqOmwwGdiYxMcEYPg
4phkYS2pGChvOAXxJYg3u08ECmmmXEjnOmuXR3THv7QkD+8+DQ7axKY8rXHtFv7NXZu7mToTIqUV
6pYRTz0ubqDYIhJO6nuArTln+ebfU2NL0ktrLcIYOHQw7Hdhcez6AxIswOBOnwNaRPlQEyyGhujq
kxj7L08Beb3QG2R418vGBqVgE7plnTuS+ta4nW+yCkNP7VoJHJj3/amUDtek+Knh4xsqnlfsN4XM
gMTVIWIt8lZXOwZkR9Uz7/rAC3L3LQyfBSXP7utH0Krw4jIXWr2W97wBDkAbKJRRm1OZQKHUKuIG
XvW614TUXGbE4JSUw02Smzrr2/+WM7C8b4R1E2zfNYAoPlvtLT3tHpLe0JWVOHOp/gyRN1UA5xcL
nuFNI/ioYt3Rdbu4hhPAyrGOQfg3u/EB2HsJZCm5t8VH4hY9pgDWe7zImV9bcSY4FOjuD29K/Srb
h1cJVSAR49K4uuv9GsSVpHmKfV7JQomF7SnbC3WmPI9qAgABtw/FNsiAbG6x/262gUATItLfnxwZ
02FU3PLc0PvbfdSSSR3iX11pHiGzWGVzwQpb1XDFG0iWRo9W8FU543zTRflKMeYaeQ8AF6Mu5Den
zHtsJm8GN+pjhsEKfD2K0h4PXDIIKya+JdCVINoPBV9xds2SBYBxXCrVJSVzQcKKvp2hYWLMu5wh
CR1QfV2XTLgBlye1BDulNKLVFXfapRd3fbKiC/edOXjRex8+9v73ZccaPFFP074md6lWRhjCxvgR
yjkkRjGAhGwWWJsBQS5h/e0NUyWlksy150GliWJEdkZpHFecXK20qQ8sirB1Gcf4QYcR0OCMvhW4
1aI+LhbPUafIuLOx7xWsJkiCIPAZKS/S2ZBGAaAYvqCYB5XC/3l1qtzwTBXtmQ3DHtp4+TT+uIJi
QnplCRy29zHFSe0usz98gS3nrmc++vKjRspuoJWNd6WsztgG8BhrUQNGFFLF9crXDgrw/R0LZ96+
IdTb8vlZIUds7pv9v1eVYwXmqEGESEPACtzoq7WrprRfKxy7JdzT3nlvs575Aemaq6dL2/8HkNPJ
miDcPji1heHnq2+0Q2iVZb/JlKhPpQw7tlkjSXJO8L0wS7P0Sbr4xgYoGoI0Xqt/HYh9hJ4h7qtQ
CS4akoMgM0PmlDcacbnCIqDmvfhLCXyLVCAfXUBanilVcEtleVtfUWjan05spuSkScGZQarJlQXd
Z43uCMDBeUgY3XXGLoMC98JIYGBoiyTj8rrSSNZ02/BJJQyBHr8yrynXIoqS7nGq/wYXCI7tpHjI
9Dt6KLZG9vpvnBOHahceOLytnkAGoJ8lf4EFvR4CqQHI08IUCoezybUN4oo2Rnpcd22VXOtovFIu
glMbGPJZHYNgFGJTXUQNOVSGs3Py34q6wM/4CGqtzPyVO6Lmf8740VAqCJsvjvYCe5M2T9VYrv07
EHwq/vHdhIBccuDyvVU4Sb+74xlTXr5oLwswmIha+NlB5l/MeWfomJjdkuu90at+e6oYV0Zi/eat
aZdQXZD0Z+WQ7aLjM0E6O0ejjWc13ND1jee/AN+c8igiUJ6vlGjrU0d/yYXtG7EEKTvWJNsN9E8G
Vj5yxAxkU1vHQ5WgM+JdSl2ntAzMCXtO0IsBXt8LyIgpTeY/SsxRSLC0FJlbBfWyB+Y0R8+sDTdL
6HCCzvzevqzB4JpYgi+pTnx5M/xjDAvbe/zhxBT4qMwLq56aRnczK1rJgy1sCM80NZqesZxiBHCd
z0LCvHu/oymVfGs7f+nCG9gy2K1fiR7+gSFeD+zkoygJP+U1Cor6LP9w77VOJsCC9usCK34QxeIF
kSloqavIGYynO9LUBmdhxFOl6DZAKIJS/9MZ06LxcdOTmxIRRo6Y6h8hpIR4KEZkD6B+cRNULJTI
wZ2fCi4ngWdC3N/qZi1mqLOYxspRWZPtVuiS2sALwIqYptL3PuSIZZT7pev2A8ocjXPjB4BPWOes
88gk3Fb82+1D2tpjeAngK7wR2NawbCN9SH5OsvlcwvyNCOlAdN87H6hOqOVqu45yE/brJDBrg9MC
eUFyv1nta/MYe0ffjhjs3MJqthWOh3tjaCntZZelGD8I5xBJZDoYDosY2fgPkdUTKQpRzoecZuz4
VKKuIy6qCugwI6wrwkpGlr5ViorFy4WWtmtt6zMltHoAy+8WyX7Kv4eMnlRKdN3TlpRDtJe2Z/Er
2gRNV4RHy10u65KjozQdNrpLWrwf/qYStR4eei/onEvah0fpEKVIWNFxNn03/VPylQc2IcIRzQOI
tUyYmXZkYc312PyAjf65ydKs8fxMOWeJFIHdST19n0/WEbR4jh0L3JgmR3+fe7czMThRCRKGgJDE
apGBmhAMItYBAPRZt8cEsHSCVrf6U4n5wSJy+1aiTJXN8+mh6alSEUsrrnB03OWQb7Rn9co6O+iX
P3I/z9dbaKJCnRtn+JB7DJQyH5viOFwSrZdzWKokyyTdFBeIG9uO3LSxuvvSCxqEmM+Kal0SewAq
QklZudq1zepLQwmqVDgUeXyPysWJZ5EiBoerm8dU80NXEqfhu3ZH0YkivyiDH/EveGkK2/t6AL/B
j2tH2Qz5QCiPC7nD2bYvmQurR5a69XelzLhxO8OGR7CpqaBx0pJdGs90yNTftRylB5tUSj5RPzVK
AgGIuwn9t0m6zM3vmscV8JNiKxp4K8A2FZ3bp6L0NRs0sDo3vBVA3kRK+Ndq8D4umA7mlsMYKp2M
K346G2AuOKU/aN5rAgcuRTuu3Tl3RT5c4LSlBI3a/QwAopVaJbnYrexJ8PuZspqblswM259nb/Pf
qxiDkhTWVqsDwWUO1eiqkPHd6G8kB8V9Qd+IS2k0Yb8gWUHWJHvQsQ+ANIAqA1SnKXDeWvLA73+P
g3JuC5popNPfyXnagK1w2t1Arp7DqI5P/w2EQ/FZvVvr1167maYBgOkxj3IAxLDiuiUMdWbgoC5o
nju5QCfqWqzCbeG3Nc4PEyd/d0luUCJLB3Qky5vFuKVBOCrMSvPK+dU1KMf7jm93yap+YQIlZl4Q
kjd7Q+UVgNY9zOk6VL3hOlX8xwp3+QkOlgkRertoEelfNkaNlh4wZFAlekrAHKcuR0KNJhqY5n8E
0nk/Dsbs9IWuvVN1ksjeitlpHaYwdUSr6DxCM43GAOwpInzjXN8Ula3d6eT9vImFXJN+kzLOvStG
YAXGC6oxps+M0Hdg62uJaX73uZ2Bw5NSDVTV1T93JRx8Uo/mN19+aD11PRIyyC9HjTRYt3SPSKJI
8ebo0QOOmvIlBD9/kzJJ7LSRi3+LDEwBZCjPbhAUCO+MKPrSQwCPGjdk/ePh/XRsY2CHKlBMlF0x
TTc+ErMlwkD2CZSG8X03u9qw9O6xw2K03vMkRz+E0c5tcvKh7AePlTBHtbCwKeyFPbOrckp0IscH
riMebcTyaTjdx69gklYRNcoe22OxgyMxagyXR5jvV5FG/WtCBFVKl8+lGIQPpl1xAd3z6baBQL04
37xHcw8QDXnp6vP5gT+K/a9XZtN1CvPFBXGYeId6Rs8Q9PSfHTd8jTN3W3G+P/hZIDLvVnv6cKwg
A001m0Q1iKUMiVJMBFvkINzf1RiosZmcVhTBoyvVih1nLXx9e1u57n+fAlRmESOVbFW90HjfCMcM
7OBnet20R+XgEbulheiwBcHXCKme4ZTO8ss3zNN/bSm3c+Gtw0mrqTzDZF+/sbsNQcXZPkqjGA6q
uicFli/s2Hzu4j3leRdpx9tFA9NVKb2vpjNrzLgw5S2ZvHdJaiVEXj+orcjHK7XmmVSw8l4Jp5as
T7a08R3PzF+Qy34+tED+3EWKj68oWYsZcPHPsk6jWY34aXzniil3PCyvz7NlgoOLDhRXslYRYA2S
axANDHWEfNB9iQpX7nKYg6VkBo9yq2DmAgM6BwmrRvap10TrUo7GT020fFZUNhdaTKpEQHlGRPZG
IpYhS3OOI+9/FKcF30PWW+LA1Vyb+48s7QVSiDHwY/T2x/nltaP4D6Xy7vNMAanos07o8lZtUAmd
ry2ew8+zSjviuKH2mM+m59IC102q6ZlFW6EpBj6aCIOIZPFpL5VImUvMfsGRLYO8CCxAoJWXxqyz
dTwQMfifl9IjqukDuLNbW+dPmgp8PnY71e623kUAlEu5SZsSGASE2ChcFXRe8LvBEdyeGkwyOTC0
iVtpIfSMi+K1wYSriKnae6uhCPNpzTXlDQexdB/OTt41E/JGYkaO2hXFLuWPv4t9c379VlvYxL6W
V2OcFYFbAtbC/2wdVnttP8Z5G339oD+IETz40VDsXT2FxdhfhfAnhnlOpmhilcp+z2b4CEyn78UV
FGI4PeVyMogIP8VaomI5CmOTYBM83TWhFOPb2rahIgC1i6q50X2FQjUS10bgFKgKIVbguDFwZZpa
t/+B/9xCuc5qULoe6ZacS5GL2Gpnah/wE6uBnyQiaHIeyeM71BjKA35MYHf6nLaAkDXpmCt9/tP+
Pna5JU68tta4yjxhA02YkcS+by+ryyc40dsE1dvatuAEM2EKcObfTHebPKagi3NrlPw/hbcFy14S
7I12z7Vc7V026rm+/8uy2OI68557fMhq4HAkyOePy63ryi/TAMdwf+h6wQHWtpFwmdFdBnHWHQs2
JcPArzACWgF1H5kZ6yX22Uq5J/5vJBzUSs3Huc/B58YfZnBjy1+gcEmuHYD4eadPgJPU1tPS7Hjt
bumrLyMGV1Tex9h9WUiEw5CzNm9xtMMgkU4lchCvUov9pC0RayBaULMlaKccX6ALdxztC3SpP0kU
cNs3R0muOiEMOgcTf4T83Loe+1jVYWh7bAaDWjOl1oDLEGvLZBoVM1gMF9+zoAR9tv5hzEi4pyXo
N3pSOVhE3ZRVJ+W3SYhP8o+AAgH/R8+dGdf35BNgDSYI6VdMOmsToUJwgmaPuYvjWFIbCK855q25
1Ku79q7vT6svVC5Svl1S2MYzfJtsa1mKxx5TQs9ZwLNPofzIQcocysA5aVKsExdUicgMkCZKjY6o
pMbALmdH53ByxD3XVbxcHFY5XPPX/vjUruIXvCoRsWA6jWLev7DuGeRXFpCQrmoj57KsTVRfkOA+
Yo7pqdWVcEgX6FgWbDprHBfrrTIAiK3F1Xq1/1kfgWP2gdPmxl598VMWrPeVd3pdQqsODae18jOd
SPKpF7CYXSAXslg9r8iJyJHEdS/+loTA2Okjb1PJtyZqaejQYfTe4J5pQHVqm9wQrWxPRAV4S2Lw
itk2ubgR5pPjaOFDw183wMU8n7s2eImhaj3qABv5MXxy2Il38CQwyd91cu04YEqjmtk21g5boQNi
xZAWNjfQjGpHFcQlGvbbaDBS+y6iGr8xa7eoDnKZO6gGZI/PsVHakVM0bv6L7b7b1S09Y/N2QRpd
YtIVSsMYGTkuJf+LHkb/RLrsDfyHkT6yE/TTzesDW8mUM4tDxxsYz3i8aUklNwxe1Inka9KM1Wyt
oOz3JcPxIj2CTiR1dQKjU7cLBSpzR1Jutv+3YNtaqL8bGq9wj60xw6PLWncoZ2NAy7uVtB6rA1ng
WG2BPWknWPX0j/fgx5/mSGYyrP+R/N19xBLsP4CKPjVJ6yYROwypwVBpCodDy27PtMR4/Lvl2RGJ
hDxKJzRQl3/tLTBcodGTqYladyMP2SfuxRywlZbbSJj36W8/2LNw/mLd4Q6QfKCUzLUJmDBHuTXo
mLA2JSrV+/51wkvogc4gNU8hAKC79fYWk9rkhRBu++t36A+Ji5ntT0AMoXJFX/jlr6VxpParyy84
LejwLUCaKsGkJUL6enqaawkBY4mQtouNaQjCi/SOiFD8Ylg1pcxn3FT1RmSqdCnFsdlrmysHWUZp
qQq+IE4dA2J2mP5DfAd1gBqYzw5Z1qWKCtAGOLcOjPBQQyHSDJwQu3+cNIHQKs0kw3kidCRiylKz
EwYtg014qBn9FHgxcuLWNFfMQBO1pihBWmGl0zoViZ561DXdK6IccSX70G3BoCmW991R8V+/5LjC
cJx2T7tAThOw3Oy8fgV4zIkioDBctsypI5N2aHdqIHFPYSc86U751Qb2UW1J5qY7kaZR3SM+ZCw/
otsyjPb8SWG0ubV6nE4egKnngX71RbUB4Q6QSPN0psjIpSzogW6yMlewGqIJ4H+merFK3REvPyvW
vuBycQsa7ioA1iKEPcYoYqMgipYXLuAcY4FaFO2Jj0Pa+VmT0MzDKbgG9eL17gSWovbsYU4NM4v8
5HcixJzz69tTPu/6sH6o9+FCCmTv6cmJLW1Pjn1kbpg/1zHqmPDlw468AKyDujSYDyw20GF4knxn
/zPtvxSN1kFipszZr/eoxJli3+uBEf5fcdTUcMjLNignp8Mp24M2NP+ETOcB+cEtmc31ucSv0sy7
wFREdNJ5wu1tZJSu9e257D/UYhoD6bALbvwMDiZy6vJHzEixOjTYbhCa/RhTrdBZM7DaYtNeCz6C
tIndqwmgai1ZPstCvct9f5UB60RsEfLCi2FYYrz5Ie8cL2toW5/7NTBjKBdTYxWmq4yue3x01Cgp
EP7ty81P1KGa8VEeHxnj8Jb81rrHtkDhbYXnlodr+T/OlDWcl2APCbb8bfOOw/hb7SoGdBrCRZmE
NQAeMK+KjycNX17ahaZN0b1k14UOb347PCCAxoYYuHmt8ta0AXZeT/0pqATbfmQKENQO23VykZfK
7hpXq4FuJwjDQjuiMAuufLgNTD+o0gnby0j+qEpmNwTFKSUUi9JQHX68jkNg4ff3gCua76rmO6Ep
NkHnWsRcnt+XAitM93HBwe3jQl4/JKgLAnC8VXJkr3fHT+XS4B/gXCzIUBjfCzFEbsbkYY4+CpNN
kqBLuQDZOX9c8wmLhuTivxQMKWGjTnteIuNRnYip6RDlf8zDDXb+7TjuuVmCBVuQ9O79XeW/4hOE
xOzLMqXzAmb6DVp/hfsrNGUiYii/+VHVL6oxiGB3tsJrzPHScdfqrhfb0J4bAFB95J+Hjw3jq2Re
WtbqdGoXsPBI78+0CtfttKcXryCbMDRoHtn4j5BuFKkcJQ9yrH/DbdQEnsdPGx+oeanNQpam6FpT
Dnxkb3j/A/O/Tm4B0I/vb6ElQzBREFRX8xx7jLC9p/gJtHUfuKW2/0LftHi0be8VZ2wujJHIp7+1
P7gI5ROg2yXGtddMj20wPnwdePeOb7jEtN8mjXIkNFYJCes0k7DemsypF8eNWZmMfyA5Scsv9wOc
v9diSksv0YrSupzd/1oDOPB9zDcHbwLh9LqeigyAUn+TcO+zhKtf137j9+BsrG8QKxzaB8MZMfNo
Qr6qS5S+riVVNM6aM7dk2jq9ca1G45e85hoH+rzCPPzn8+SzesRwfUrrCLjI6L29KC8CCQewyB6+
+jsC0DfSVq1LUfFnSrXEInlr6/rwLLqveEQbWsc69n+z5MpIqV8hKtj5T/Tp1yokXlsS6+SUGf84
U+ezgcgDmhisJCJRyq7ggWOweOMfguQZz3239Hg5rI80/aKN00MvqKjc8xwZwlhMobsOsjOM9WwR
WhfjgcvyBFr3+hcol4xZA7wC0Oe5nLOIcAKECzn9MPwRkTrl92hoIfugSbP/tVY6Rkb+5GoIETKu
HkAyJD8Y8PjCzEXr1xEPl1tCwgxwPByIo5BplFVOw0/Ug20p3BLZCtLz629J0Q6+nR/SIAT3jggk
0+6WNU4sClLJED0jWqNhp7TIrxpkRgbK0RibPimmGfQtAIPu6vt5YBLfB+RqbJtFrI39iE8GwT6e
qNFlWKJQomyZVrgRCG0ILwE4SByx5CONL6CR+7ozA7B0fYu8RtzFS/OUg6pWC1IN/6CsD9HHic93
4TPaG1Ml6RxSemU9TQhIB76aFp4Ru+vAGBQN5478nhDwfYX8a6uVm+Bxtf0e44jFNBUJr+lK16vK
aurhrls3i01BLbxJU3r5IbkjeCvxGV2tS7hmA0bPXDzurABv6qn2zH47DyM6V/Xdgvub2qSpuZ+l
sbLfLWQGfQSEhU9ho66LPGkVn1Ls9VD0b0QvYMU2YkUgSXhzOW+NAPcgpvslNtEJGqV1wCffN91A
GZINiOD2ijT3Iq0EwMsR9JloaVR6y8tV/1YZ19FI737iz/N7zDZkrQMkBE0w65psAHkXqYWs11va
vy6WcPqQokyr5mTYCoGRZYO4S73gUpEIJWQda20M1R34wOVEzNaJx+UV0FznisNK1ET7VckKuS0Y
WAIMOCOpAhp5d+cvdyE9e1Y/Rgx6qd/3sZkNnn9nCyX7ZEVPI2R9jqK+VVK+R2Y26d9/7AKJkLpr
gcj3zOH/Rn1aZGzy4qotBOoZ+nygf7vDIYn8kiUmsskpsHyhIFsXx44filhBq313yRH7smD65qOa
ktOr26RiTv2EVd0ca9Bs8PYtgE/WK4DvkI+sxhr0QddVreWr7NONT2CtdHINI2RvTCGK44FLiznP
ywAMGLvnjC7Y87yPL+70rORFHk40fkW8mL6By8Mrdnf+xVceBMhqW3Jd3Mtj60v+H+nFjwKRMmww
2FKgrUxn+V8pptjWlfqRJ2BV8fkoBr/9uzMS5Uwbc1eu4PsfXvk08Osja1VN1ltNp0uDWKkGU+/L
JPchkNpiwe9S+LUiUZx812pIQH3GN5/mjNkIacngTsa6R7RdCScB8BcTt53beXslMuVNO8VX5nAc
vUbbYaUpqpD9pnRTjSP4ighilTEwnUrRw9WUhcurSOy2bidT+5GVbSmI2apS4F3WEnlqjP2CrpVo
8ApkW6IL8oyJBd8Yw3uChuwJolDY7TJ9Nyah/SArggCU//NLpIj58OkxB6a4DMpTmMjyqF8NLjIc
ASpuwJxIk2JtqZbcAloj2rYE6k/FjuDcGCw8+0XNg5rD4ZvluuFxSBWjBzB+48DJtilojmurgtB/
P6vCiRngHZRp2sJOHHME5T1Bg0aqRvXKYFREBFgZHu4MOhpx17RRdy96XPqwX4AWyGjJgQ1CwE2n
iwKUknqkNdPqPECORUi4j6MHlaAYSlT8F7FHnvgqjgvAIJkZYSqALXh/UKHCD3lHFUDMX3rZl6c7
IM/HCz7j0Q+9gd9iqaxkPGkicbNk/mr3e2fBuvxcCXzyqydDOoCpq7lgNbmt0POIvXI48ITXcY6f
VKDIpDbBm0W4RaKbPYh+rccQsMVF++Xt/XstBSQwcw+U4qmxrE3TtCKOEHYRTFzNkkp1jeEXlgyN
FG6SIFoGGxruBjU1Y2Apbj78TVD2bSATZaw9WwMuj4Vh2aJDApqz9fJ5x+blp7C1HapBPj23KnXr
Rm7oL+1iF3CE6vnSzH6HGNzyF9XX6yeK3BE0JdUuJ7lwokyX8MgIKnq84YHn3lR1wQTZsVG2cCmz
b8QTouDrzqUxcTutCHBDfbOKpabeASzU7/OYDTq/TJ1/jaKTS1MgjqBQJWmWoznExnByP9jp9dif
Np2rRmROTK82IrcWzpoGmaCdY298Vn2xTeI0FUtJxLoZbk3zFOCIZv+xXVPlKvmfJwepP/kdZyo7
1ElkgE8XQNBNjUIXpvEvsnnEE3cetcaVv3dfSGgBy8ryBlPtRly34jCccMl0UGaDjT1E1y8hPWOb
oEsiamcUUJZwXdLuz4GYSdjx7Fqt+KGBIWho8fN6lel/6nEUoC2mADvCvCEoepCqHSAXvfgpBHLG
oM81E6WUivhu/aQRnY2ZiiD/8WS/W4syldY7Zc0MFuGXgpByL8mCQ/5jovZWmYQIHz1Q4Kl+9LKF
b0ZXeGnA52PWWwWhDr6y1e35kp3EPxKA31A6yT3+c7zTCQuTLiWsqStuE5qb2yoaHbpxX30tCKz+
c1xn/whbJek4qZCug3e01WrUL97kS3FRChGyXLwcHPNCuR5e+j9+q3PUuzBxYvLb95lbUYTc4E9e
Jz158g3g0mhlYmzBzh6UV7V/bWx6GxycPlMCSAg/iDcbIh8oB2lDnTbsplgL7TyrOROLhTydtet5
x8nzLE8n7ZLgUwo0Dg/GC+wkDrkgiLqHMbJhiTzDTUoSD9NTC5UGv8Dc2NWkWvwQIFQrp6y1WpQb
aVQ5x6h9TGK2ar2kIDZcLa9o/ZriXgxZ9uFv1CHuvw14BLoYi/vVWCjzCPoLHHj2NdIfN5tdAbw7
lLfu4w3lTY7oI6rRTCXHQQDXILQUsOWg1yY0EeiEAQiujoSIZ5my5LaPGTJPYHm30EgoxsuF8p1m
lFdZmzJRD7Sl56zwTyUOYAH6spBd9f7MYJzF/7ZPtHb0lE7UL+lIOQKobKJQp42QZbY4rZ7SN2hK
eOGm6wdJc1E1Mr4/Q6blG9Nh4MNXs6ri/WT4CKFFYn4Mr1jCxHHWnmZzfx4AWs2ZYJcdXG55Aqvm
QqlOO9iqxKyV1N0j2LB30FcmCj4t4AUiwL/p1DRDahp0jHMCHzRSXqAhiRWNtq9uOrc207QeiP1d
JGDyg62ef8bbLkLXWaegqzWWVMurYYAdmfUxDXtNIoevy5mWdxrRaRlz63FVwTkKEXRgkB5XlHf9
StwH+HpPzHBVGRS1creI0U1GO1J0H2F+c+sA0OIXDTnGY8NS5qbQ2ahkseWM0TSO7qZQs43yW5Z7
LuCtP94OHMcaYdLwIIe88CO3lnj9UhrVt51nd3PsxlZd3kVxJg5baUC+pnKSrJx2l9Fh5LxTQMNw
KwmA/2T0Q4cS3KcafH523XMC2mPARARdhl5yQmxHu/WqPQT407vtPr7dSTWSsgm1kWksOJXSNxA8
kGeJMgTFOP/I5n1EHB1VjjbDC8buW9X8escpwvFVaRA+XBG3Qmk/k2gLvav/S1MGHM4xAKfaMf1v
qquL+KzspOTqDnoJjlz/QEETXq+ImF5O5YOsDPKTRsHAot6hAYFakysBfr3EDXbGyO8aCjbbTyfI
KdW40TK6bj/mvKutops8FtXNfYsTOKJIAehKmQa3Hf7ompg0/VZzvmndGIrcsoaJDOuOAd57e8lz
CnVn8eB0+re/i1aENZDHAlIvGyaIYLoiXBfyjxuf8E+lkQTldsU4wZ+kk7RXucMjCZpQH1Sj8bKk
Re+Ge15cZZrGbRfkoljc8pSh77ZAGWqCvVsAsqmjO5N+RmpZSbi6szyS3ZDzHoAmhlCbjc9cKZpE
ufzEyoiJrtg3vJ8GFaoJkKL04kbPtsNmW3fvAkgHsriy3kk9ZJyi1gCMdcLVw+QufCw4z3kMQuky
WvWhA5I+n+VhgGDaH4aJ7KdxN8d+zFvOH5J6Hg1B8hwJHS+ui8inYSKHqpAQOu6DFw4Y8dUaloOe
m5E4me+nkZEThHKjak+97EET9sq7ISrQhHaOYissPwV8zMLWmKaMJt5Txw2jz5b04yprZbsvAIVe
+wcDtV+JyuadI5EsvYe+daG5t3ACzVKYwK80LeIejTrzYa6jib4BJ1dJWXNk3mffQHOL/c1eA8Wp
srDo99ksWz6qmxbmshVuwScb6Cf4cRC1PTmJv5cNaes8wwk1waxyDhMsbEWKu/y3towMiZ0SYi8D
FKmOeM+udsLGy4PENBTpfpSwdrHFSt89ANzxS205Rttoyi8zC5xA3s7u/rQT82t4vLmLUjGnbZrg
S4bN9ZWvC3cQuU4dBcMLs6qfv5Kn8XJBcwpYTkz0S9w1o4GDWmPr+et7MXTUV/TNes+bAiV9++4X
LPjCJWQMtDK1t3m1X+vqmyL3lvtm79PWKpYy2DjfKtguzUqxIo+nAetWwK5nK10l6pqSFQwWL662
05GgeBHJvkS8GOrOLuOuhKStRDNcbjgbjWbU9Rl0+EOtgrkM3tvhmhyk6Aoc5nOKiKbOlrDII0vS
sw3e0y7S6s4NvgN26N+qMqMJSraVcxha/6CuL8sUioCoGJq2DkAGE4NHfUoPqLeTMtskC4/UxXSb
5I4JKF0u+Y2AOxZTlsOrR4l5ZtOzMlxEykU5HWv2jRtxOVFiXCRSlP3R9njdNzK0dbvPTmcncJca
2EQF0Nh0J6Hq7bGuYdiihist9QgzktYs20BnqrSSJI69F911iZMrDPxq5fq1CU2l1dYOKTT9Dp+f
1TmsWw/pYcltJrhjbhrEm3HSwtasoCG3sy7z6/SdF05v/k41uV4S/eHA2SajrkcKu+/G++qcdvXE
prOUlgSrIqcZx3MA1irYDl9czxnKElUeRHatvlZhL5XLQ6y7AtSgYeNofDwMvnTmIJCa8KpSamkS
CTyAVMJcmY8aTVONdcwHONvCCFYciGKAX+GNglCOf2dQLXN8xz/KzLhGiBhFVYF7pDWG5BmNgIYR
jSqWPl6N1g2U0zwkzOabIrq9075CpjSyiImIGvPaj3Sk2swDOr3JQdlM4XtxLSs3NTOwxmnscFnt
7oabWxOm9aV1LZPAQ7H2TwMEEqt9NPWjUdlRx88e+Wd9M4H1De5Iy/GT7duatMBTd67TQ8xcbpyI
QbSRTnAEofPAWKYtABl6zra9V33jcXFWZ6jtlYRdplnhqcHb5c4As+BuYJ6Ti3k/0oCSMwAMsMMr
CkaC7TIohr3JjR5HV1CF6dxBWbVogUX3k3zb+E2Scin6CTCF2egrqHxwdyV2IPujAmRQU2lV0aJt
gA9Dmibvr+9LWiV8Xh9as1msWISkVdjrFHQtY7TzlvZdv5AGny0ec9qMnXJdrB7UoYh2eoTN5VMs
QMlkAmHc0whsNgihYP2ci24b+R5knnFGajVBOw9XU1J4EAjBiFlD7pAMk1D7lNON6ohoPwt5k89x
khjgm0pnKbSnFLhCP32wDvw/i57WP7HO5SxnznML33A3/3+0vriEmuaw/oTwUBBEOEGXvxN8+C7F
jJwh9v5aERHHyKV4T71eCxPqktoqnth6P8VK5UWIEZfVPr0VCbQ7bWUKXtyDRRurd34iQDjs5zWU
PMFKXPUKXAd3PpyS94MDEJJGBLSYFB6YVlJ/bXNE3HvzdBAtmoQGkouZGikW9fwqqLGrf+MCcMPp
3uCmkFe0FZJ3WIzMANTLhSzT4IYesYlr+MIUDLLds+cSSL1fbOo+0KDlYfsvZvPJ0ytkqdATHIyg
rLWuy/cQm+uCcXFr/iIbsRxxgcdbbAC5XRQZFJi3NX67f/iZ1je4/RbmFLgN93+pb+FxOSD/YSC9
gnQJnpexlERAl4prpgBWEBV2ZvzoTqGNsticpbH323+fkcxQZDI1jLSs/BdlOKOtamPjPMJbxc7b
59BKie7HyLhrgA2QPDTXAvs8U0jossKjhEGtSQBNzIccNVNknX8VV+b3pir3k/RKTPTnuHeRbsHH
kcONY9/2ibp3iqHpKz3XxnFCYpIVhZv4e0wvha4KikADZ352STMHBli+EoBmR1KF6Wx1CPAWTkHl
uSkXRDOsGUzK3N/5qK/Lrg0g6CWVJAi0Jx1Lyd21HTnRat9iTXo8VyqNLgkh7P5jBdTXknu1+WiK
vulwmXEhUBiaRkavoVSKCQiySIi7xBy8W5bYRzgUiM1jaELUdoYcw2AwJK71UpkZ5d3uJzOInt2W
heNiaz/SBXmN1gSHYCSP6yIoMZzJ3kbnBMrO1t0zqjn/242BDb1EBQIbnZQ8BBp7J2807HYLvwza
JqHtCw/4wCpIP0iBNBcgCysDEsImFiKR3v0j55S2UHie1LafbvQOrRAbHt5opMYt3sI08cymh+PC
WTfDhe4D+qQfb1HTm6cHROAMKaQYLTlHhVmAQ710piLq8o2ilzLi1oC+jOdb7ktOcDVsCVO86WpG
PEg6njwe/cJOgVqXPrtByuLJWAmL/qCNDsVPTOu6LCH2sCtm7AfgV4zG77OIUWBBo9LblZ8QCFzi
Q+DmbUfobOp9Zs75jqt4jHr34qyHLd8eAESELcYXt7reNxE0oOQm1aR7uKmkBjPivPauWLrNlWHS
xCRcwHS2/w/Wr+BUVCdLXLGR+1aQV3mB3n4s6w0V/FWX9wpnTuBEDN0uXUHi+LjvO/MM8vqCKvYy
SNzvn2H9GFbrrtQGuUSk+NOM2ozuXmn8i9PTK61huRtUP97ftr2O/8P3wEKrtoQE+yf6vMEyLss/
zoMrrhvb0xtDrjMyWWKK6CHoCrfBD9jXAkk0GjuZxREJEM8yzsqEZDPFacopGPO/pRtU3LPm+Trw
eyYCtnARZbmKFEwVzIVVno5ANg9s0SWF5+r3R9qacVcFYFFMT/Dn2R97rrqCP9bhXxtaMi20wGCO
3ec6/8FCHhA7aZpENjT9JQQtIM/8/2fqzQxSGFUETLenOXGw5bHjuo3Rz21UNdwsiOkAGihUSoZG
ErrwJnQxyWb1XyEiCVg9ujQw/yVThe7v6dmJTvsteGHRTRBW+h03hxz+HjuHlkYn2IhXORhVdkuK
SbgewRKahrKP/cgXlqQ0tbxrJcJmK9vQpu/cDVow/610eTmqTXBi0Amt1xGJEbr3PGpNEUAxVN9a
RUr0bjS5zJRUkqSEFd7kDJhdKC8KcwceLM4XxdcqaQkBUPO3qV8Mq0QJUMKQy8981cr+7MROWwe+
M42RwnXG6NYVB6JkX+fwGvrySNpyU+Y+BEY655RQ6e1eg7bVjNlpRkBks1E/jEkCQLXgxcvgW0Cz
vqzWin7cmDb6FKi/WP01w0Xc1aqq9ItUcQlVph9lUEcoCxnjrrzTJ1lx8sqZbSGxDv4dUexJZNbP
ZKCI8Ri40nLAfhlj/Xg0e/jarlI+B93A52ckwsFkMRcK/Cx0NGFKvWY38a2tk9Wc8GArPQVs4MkI
bJqjjT80iRJTooTZH3uRLlB7RZz2pq7/Zy9mOG+w7f0PyPwNqmhXq2vyPs2oeXnVMiEUnZmxE+WJ
RJKYMjKmHdzFm3rovqhS+FAeG47jrebIghbP/0AKX05lm9i2vKgYdlaevnCqmf/Loz5mjD4akxBt
dvVq6Ky9V7OHeh/H0gd8GVuSLc469sIsRg3NZF3bRmh0aTija1ttgjYN4Ph9Jx2pL3L3Q8tVEVa0
lmoPnnWTuhHoCEZXqolxL7yVlB8cqIR7UZ/hs77R6wAvffAKCT+syc02zJnEkhjLrFb7C0P5GJzI
8V1doOZGmmUpNkdSU+pUi95UfmAAkdCtNpyVu8VmoBccT8VTGc7vL4qgsegercEUlbiW9K5aNPsa
Htn+/rxjHi8YF/440lNwWgW+zK75iZ+QGK5Q/FFjAcVySDDNWHd4EU2Bsh/PO7k8ZLtmxVUq0tMg
NtOlvu+h7ufQ86HR3smNRiBtqgRxUxUnmqX9qRbEYf8scFxmNJy/fhPoxnvuhltzG01ZuCSAM2dt
B9aWbiqvUs6XkI4Psg4QxFtVqK15rC1pIyym1cg+X+XaVKGSOSXgBZaekGb/cU1fxHDfPu+UwV76
sOzohYpTIoh620aTU4OI0yLu7cscLGY2AyRH2oazL71cZ0YjbA53V6Q01Bw1L/EMD8gZ6Neir6tP
8n7fNTPNQ+vM+Bb2X6PtfqX1HRWGzmNEayluJwXurz4h1yUXsbmNiId/zRuhXQ3IUNstvRAfp56+
0wAw9bYK1rLndPvlw4hUnZmZZTLvHe2lYM28rOj8f/tP+aeh7dvmdsdfl9+VqsdnqWeGNa04puc6
N3IyaFU+nlF5ff+hACowAbfsUR4d/NltvZ7KiprhSvqE0D+XzhBrjaksmQlfzIXG35k2Jcz7+Bls
+KUAAWS9tnsUobYmXyXN/tE31DsPXQc+K+v/+5M71Zgv5wkJp89bF/ou0GC5ehc0ejThYMdyhoJ2
GZNREClw6EANUsJnn3lg/AhsLDg4t5bmCzqDei/gXIj6rNxnIWvcv1oBs5iz2Y3OjmiHj+FpNFSb
ITQ3KHQejLMna9oCleeqiF0A+d+pLeY9X+1KTcU18zDSx36zuj7g5a1pf4qsTOQoOzud3qfOBeBb
v+c7NbgvsQgzeBePL86UY0iii/yKbw/IKe1uEwZrcZ7bbXlK/rbJgbrL7vagymykJ/+BtMUvfHy2
ImObgf8rVLHs5EC+fgiNHU2GcXQYy5ODxovMJyCX4JdhBx82stR/VfC2oN2IOXzDS4uql8E24IpD
qYRLdagXHQWD+IaDbPyiUXUUCeiLu+u0P0sjvroqytF3mYpD/4ENdrbu10uEIcVfDTR0o/YkZNTF
fZeCQxHUl6tKBdFnCyPWR9RJIm9fbW73RvLqARsDF2vsq/UvJ2T2ktd8Yq0xiq1tqnWg2F7gXQEO
+GlVY2QyZeE5GFiTPXzHvwhW1ml+sKrtCQpvRd5yo+pjy2hCSxfbQkup3x5x0ZRKY+Wcl64hWKRu
FpHo+GLiF4wk+Tz9wfZwrQpKR4AVx5tgZ8Fm/7i5sJoNkKeDPPuSIbyMk7zPA/gOyhO4xpqpjVVO
2zwlczHnPL3kXwZ3z3EqyiNoaXizcPFcxWRqEcXFEus4lEWjgPFTDqDunss3Rjvldz7tIiZGNUEF
m3FuQYQXbJmD7rch2+MrPRte3KcP7W6OaZSZvDpuq/5JZYcQrfupBJSNqFD+ncz4OZVDx94MDTbY
BObe+54Vu2uWkYiGMPOebvUgpbbVg2n4JyoZ9uRfmm9dKs0Q9n2/aP6emTH4G3AvjzJ/barOiZ4y
9Thw7z1KZy6HA+yDvTYjA5cHW4lUT1xqBPZWrqYehci2IL+1wHVJsjb2u2f3wgEo7lHfqFGj/N7a
rS8QCiEGF3oIeuixfEEfnTCTfo/0mOtf666GUAYMa6j15gvIC4VqUSKm+nr9JaPKMGAF/WtJWirt
EQ2jAYRpKCI400EliUcZ2KKc8aqg8iHWngISPpzWyu+DPEli4VYe2NDoaSQo+NrT3/3htCIaB1hY
cP2N3qA+hy45wMFbmi4hfFmbrUBJ2qFyxBFc0j33iVUqTE5AStryof0VeLCVu18cYycsi41dxMwN
0TDKuOfB2bPbCqt7rpSXmlPZDTpNUtMx2kR7mSfLN7CwwOS6rnRWzGEGRRxskbbnHdvqRJpnRRcV
QTCrWYhEEfRnMKujaGLjE/+N0nmFib1/qnhsAyjg0KFlZ7TT9izEMx8lNolgeQKHumWToUd5JC0F
kqF09T+JRKv8StnoKMJ4pwosXlL94AEEzOwkBeT1MiQyQwoUCjy9vwVP2Gn9thVu3chK54eP2q0x
CrdTUDNQriWpPDqK4WoaqMpSYZ9j5R5N6vh0eBd2A7cXN71CI8eNJmIDwvYAKCTPtTPRRn1VOdYh
/XwemriKLdPWK4184kLUcGxRe9dx4GHwK39B0dbA1ws3Xg6V73eu4A5bPxOh1jD1drmb6vPfUK1K
gf31GGFJjCPre3jzFhF3izkt0ZimnvBvY94iOtjACpsGiW4l+51bGsW0CPth4NIGejIITjuuFeUt
58PGox8lOsy4qyuUUdzSL/o4dcZzAdZA2oR1JQt+l9Iy5SuG38ErqgRFqNOXNr+VZBSpDi2zfEuL
v08Wlv0CjFEyEkU7PO6Je2wXQNVnGB8NbIZWvn2NVX9o+fp2nvZcU/YLCCyKEfIGKkzVpqeWlx/D
GCf4y0m+m9XjvR6be82tx8Gfg+u0H0lJbCcGQ5F49oAkm3c+tWJ8Z+hjFpF0vKjce8KbPdIKnGH5
t+LlTbo/7CCT85EygnozkwXFPxXdgZFrM3spUnuWt7A5+n694wkRwpr56YYHHUUKBKFgS+kXmfZP
jE3c2GHZcSWqrxR2BexJSZJFfV5TFH3FUSqNdNPlnCSYloMU7fSG1Tm+TtJjPZzAhn6J6d8qYl8U
uREyildDyzanMMI2hA63jZj4X9LLBIg09PHdKLVL/7QcSYG/KmZFGqex79525NqZo+yKoYSSyBWD
ibGnyy/MmobKQfappA80WzVoPu/3Fsbqkl+eo/KMVTLl9dpp77sOO9n/CGePg9el22ZNnBgXOhUI
1Woo7brVLZnnfKJ7hnsLmJkr+KH0mGQGrhTRRRazZj1xyE0BYYAUEr/+Tu8pff7S8YknAu+FOzU8
6FwH2OhkNeN3spuLnXUHBn0zzcoLb0NE30Iu2Ymt+CfiXALCRRQALmNiGYKrZ9ULZC0Jw9rkBJP2
6vO/+R26kq683X/5cnYLYj7mgCEYw8jFHt2sNnpDds4KApgbzjoy6/2WwKtdPgtWE5dVlJeMKei3
ycvkvSpqEa+5GjZ1g/VGfvCde3GyIW29hFFm1V43NLWrrXti6g14V4dbUT9rAxcpPcFtstn/7Qq4
wl7BYU9xqXVyXvDc/twyTbobIMpG9K9OLxPJ8uCBk7FAW3+XxaVvxLZs+o0x5SVf/Y9iuTesDcj0
bFRrvzxgEclr21tBn/LQrtrlLk/BLrqHJ7ZJp7kGEL/S0A2WKnXpBJ+cJ8fynSHq3trDoNsCtfe3
wE5ovaOR2ljjpKPkCzBZlNGb9b/BHz2t8zv3Z/RJLXkm8uZKo6CUASdmJjdLP3Ggew2SkGiCS/iz
lr9uQeCWG5TQZ6BAtYuon+T2pVxbCPlVAEyDwjDJJLQo3VPaaPsiucXdqRDneyu4e0jW3MjwvMe+
NovPyXoNhkx6x0kMSdAKLo7/h4fg9cGH0g+dhTPtOns6yiEWRZGix1khQlSAHXf7IQs1p6thYuLZ
pOAdpQ741kaDhfEyZpFuj9JMxvbgxcQdxdCuPykfO5b/sbO1ZymZpfiLE7pB7v02zJrt2UzmLNeU
20mnoEJO6XgFdWZo5qddWMrcPwSQOZXxciupd6e8z0ffDZ878O59A+/hqnMHa7QOCFeo8xSDb+06
YtZV9svGCtXfNaHM6BSx44uwkG1H8E4UlQ+BzPoqTAaiKfarpkwYQQXkkDqdpUU9x12qi9/xW+4s
PYCD2dQolqo6fht+0uw6PQMzd0LU9+ls9wL6yfU360vZsitZszuA4IcyGQHgafai/VXt6CMUkOqW
kUoAdbPpqob2iTeB/46ZQk2F0WLc5oGpwoMjvBWJceRSCL9tThG3/Njmvm5DZwajsJsGZbwwWt1b
y8mJTTsBYhfmTVbKqGPeWbGnXqamx++9Smq73C84/i9IST+TDsOEbTqmQLoemRs6y0AaX0KOAZt8
exgS46ig+GLRvMWph4lmvZ1QqGT8fgoYnefqrz+PnWrKzl3eE5OkkdYL6YyELiKPygiJjH+fsD3s
W9+RHJvjIkoikzg3KKqnm+BWDHwXs9arj+zhHDKk0l4eM3/0V/blHxExQsHaByUuRok35a7x+rjU
g7wFMUWlgMdE55AMMOVPtkBVR7pj0n0gtgrKXug2guvLxk66SSGi44urFLEic898QCMbQoHgLO3k
nAyiPF8PqbLV/gDIvCkBVC7l1tHRkYNwpCtEhq45qMIySbIBDkBmQC1AOxho3DwNtCEuq7GS59m/
ivVLBqkGGWMiUvjxIRcbnAwcwhigYCXgyxCkKZTbEjgzAkKhCpVhjkP0+1M3YTTAikst4XD+LtQL
ydUZS811ox364tqYE4vRV7+rczMs2MEVUdISS+IPWgp/R0mG9264NGcMbwqz5iH2KxOQmIRnpQeg
uqbUYhn9clgl2FQgb1VeHrRXCkMuuLRvYqchPPYq4iDJVv5xZ3Hl24pLdf1E3jhVISY1JiXubLIn
kgg72jmc3YHfg8WDVvmADTPG3P6zsJ18BsM/ZnkBZyslwM77Pi09VquZwsOI14e5Gq/Lnvuweiag
kZnmVFdK8jRP0By6wD/If0Rko0YFGCW9QFOCqpU0kxja+idzR2LZ3ZTwVwhXRwwV/qz8lfafUdUk
9vpkZLdTU8JNJ/NidJERP1CIH3QTEHMzvCIRYIE+0hQB5G7Jz8GONQSh6iWyPL0GlAx+hCTOU666
rRynuvbE1svKLwFj1sqlSFbl2i81umJu/eR8c8ozP8PES3U09S+hQkYYnBKAZehLre4paazK+Fvf
ARH7ulfrsPMypNhcoq0WLYI+30k8dvoHBveLKBLQZvPQ6jjAFj8MjcjSwZvKhLpxoZiwy78yB333
OyOumzycqFSs2qtTQZ5JPAIWfZPO6y2PbHuMu7U1aAJ9eC0BZ2Sid2xkMSLGttXyqGb9LoITmnbU
UnPgtLQ+zv3ZGILn7HrjJTwihBLgEMO9JpXMK1zUtE3n9sJyr6QE/rzFzUkwyipdb3kQ6w7apwTm
60bWW6PutDip48rG4dlMNT56cE6qIrm+b7F0kYOgrKkuto58q7gsFsKFaLPde+xLvQENcSO/vzZy
o97AY2rF72NznJFc2BfxwfD/FG+3aDt6s3ori2YouDfNLN0OyEp7Iy1g3IrOtCAupU1G89VDwvGL
4uP6tXydUufzGycXllxo4Y5DfwJNd/CHpwep3O/DrCXxzEKj9sDD/Iy4hAB+mAJn5P/Lmr5jKCRW
OIhaEcKItpxT0YIVDJ/t4jkgivPKb/LV8QnPf5wHwULPCfzdKC/b5GAO3yodZDT9bGuG3erLj4R3
6M9DkC2YyO4Yzcr8I++hwnnlLJoGctKLr9DoFHRtVuWmv37kZt9atHlIZtz5Whyy55aKTwmbQoa1
0OS2aPywra7QK0SkYZ08D0BbnA/8GeoZ3yfQTI0+2tUMd23jrdERDSWzFsUbhgQkK0J9hSmh/wB5
IkmeOA0Aq1iHrdyFpckfZzmNGyA+jyWVtzsuCIsgIqlHIO/4ZkBBqM89lDwSqrS4o1ZtGtvZja6S
3oHtsJ+u4CZONghxLcNGN1XFUG04LfXDpO6+Zhu9IU9xKNM+kLSFyi5NR0V/c5s+xN2JqY1Fwx1H
vgCDCzt6CBXAFc/ifZ8mbeQ6WtI0S6xUpgyXVayniv+lFh3jEAHdHTAsvyFzd0Vez5G6ktcumHL+
HrMLcbrGUeUoIMPuarpKImvRVWnKbTLnjY2Aflu0kyo0IG68q5xcxpb3i0DB11+MeJgbVRuyEMoO
v/hiY8PLJ6EPwTIg2f02/SHFtoA5zzyh94ue5gd8iEd1we3THYJmJFXbnVpnDVkIgAjTbIhk1j1K
Kfr7XgZOB9X6i7zGebcVzWVWADzeiFXiC2mnPZkDYXM9YFYylQotTzkx3+/81cdyx2UkSk89F160
0ebk0/57xJxL8LFK6ZCLNqO9c5H1zJec4eR+MmLy3+khR67Z/Q2rJh68nEmR0O8s2shxkdvr3g1N
z+2TpvTeDDjTXxzRVhquSWlszQH9cwTxcEhvqSjC4bocq1LZl83P34dU0T+qTh6xLkwvJvA45Ubo
v0Xyzo66xC2027ABud9ZJDJaX860AwCUGq6nR6wXY8ZlC+ubxe5HIkCtzUFHC86KWYxAnrSabiPC
uQMXF6LlcCC/9nQUGUkZI6NxMW0UmqB5ApsxUFnzG7O6wayVYtzp92Pu/yL68NMaWy6L6sKK1T3f
/IWWhJFvZNgxPhrwkbQnp+HFurB/LD4+BqvwDCUW/tqI5d8o/NAh6sJlgDFqpMteB8NGt4Fzk1xK
MZptuhbF+QvhLR4Xqy2dSj00Iu8gKBL/b2qrJM45/bTXIgj5avuy2IoXfrtciLwIIOEWHMxQBLO4
OefT840PZK0yy80felLtgc0B1SeZSv4FW7Pgjz/za8IfRGCO3zCv2AkA9zJF1CCtg9lPi8AJ0Gqx
ZjF9CEhh/0jj6JHXlD2xf2T01DoFBbgbqQrCZjOkcl3+u7QaP+1XELUe1SvGaJaFu2TR3DSH8Kge
Yu0Y1YkxB/9Ynkxk0hMOki8Xz52ttHc8jSrdjqxFPdKbqaMfkw0Xdp804o9Fsq01QGCfnqfPyrgI
KW/7tIOjRwEDf1YYsVv++PRe8Y0kDIHyEmYPMCtWaVR1OiRFgk8GUtDFb1S1IDWl2jgaOT6yRf9Z
J+Tndg4f6srkc6fTBlty0z70JWrTisk/Qa2yFdx/7FIDajXG8SaFyZ3c5O8bapjqWBrrWe3rNjtz
9wZwwgSyCkFlp6Drdi2h7lIwH2JKQB5n/Ng1UM4uNyvUOw7dHWttTAQ61VylWZxn2OYZleiGc8EB
2fGErcXysO7tU6CSUu3cXDu/nGT0eGglpH/iOKGciCG8NJnS1rh/6qE8mBg7uH+rmOou97EaLZVH
M3n2Iy6SnUBzNDp2L6p1AJp9bidoPtvJRt5vkmYvNgNkRUGcY9e56AGoDnuv8aeyB6rfOYfnV+rj
lFuu44nlZ3bHxY85uIKDMdasYfgnUUlWDxvS1Gqc3K+0ZCE55BjagI7P2Ef34VXerOrFJDmKUyFf
nLN4TvAGvizjBdsM9/ojvrms6ZaC6JBDEswpCY2lRfsK7nnzQxnxQNXlScVrBsCgSKmQOGt9Sy2E
zCC9G3Esla3X6DkAyJwNnYDVaarDSK/LslcLIc+Pv+sPI6VbCQJBG06cwkwlyBccbTlcuR+Wkd3F
syTtXhg66wuBVmZneS5/0k3j8GerJEwyzMSCndxYFipjnLHqhGdSz+wchXuEdoTj52B8eXwM6ErF
1QriW1JJYS0pdK0ReK6Et8YdIR2CzXhYCWOKqCWXIMakU5OK9dmow5U+wxKLdlJ9T/YJ2fmDHqUd
OjytYb+getOY+ZNDNMd+hHrpycibpnbgQvhHLwekb//rlaAqTwqB/lrjy/qvgdIsPHh2nJaT8zox
JteSX4d5USWXWOyOPv7zwX2jctGbbz30a5KLGljuG35LQyQbux02nqhPGq8eakg48i0OKlJFV1Av
c/BmVHHL4X0t02B/V9ukCeJvgB8ZARMX2QiuSGCdkjuahd4huanjyB0N/cJWGOYak4yTpOz8ylFg
NDePDW3HHJmq2ES2vOy86oXetxIyjJ6fVo5TbVidPsu4C6scIclQdUxKqGXFukfni5WEDzNed+kC
WIhDaAzM1UVnVRJlLW6xmJ4rQ3eoa33nbqIr15jcAho0c6XaSusF6VSo6SoNLYE3GZBlqomk06B5
Y7TPWeH91kjrztmc9TYLC1we1CyN0AUsA/kpxwQA4+djRys5bXvYqMai0VzT2BrqzpXDWNoMYF5i
0AobNhscGmp/S/to9OHacjU1ecJfm0BDCOrBB0UA7TIPi+i6oVUnYtGMtIHeYFmdmjAtcPCNw0BE
hmNUzSPSDEdS3JMs6kKkXYvKgVesQVOEl2fE80opACFiHusgGmRATzdX6hdwqzglm6bXpDrdXbtg
Z6OdhcFk3OSoWKdqFoiWxN3uy6xrgCWj2vQGJ4V7DdeeIHL8coe9eLVdz/OU8pjjuYjd0VS2Hsux
eRFCmfywBMclWq+/3P9vcqAYmItVml9Rmph1JFbxc5fE1AXYMheJ80qGLEaM/vgfqA3mGcJAyYb0
jytn0/9iTEDaA+ptKGioE1Ms5/sJqAsp5mzNaxYxQwph2IaUlGl4PHAve/tPlqBuVkXa5lApzZXz
9H9W/YJsgZLoewBvQHT41tnfIJvTU0e+LS4DoL4vj0R+JXTIkKG9MlDI/6NXkHOZ7TNA2fgTN5pG
tSpqsHigJPEc6NyasrW4UU+vzh1pLKtWoFwlVT9PDSSv0kO93L/GR4NQWrB1E9jlpTL+U9RDX4/W
TBB8SBNzFj5vetjgzVij7MXEXQgbrFT4fVxRb7aEsgfMl/Q0VUQx2K5NiGnH6zcu3gtSFFdAi88N
XEYe6nQ218Md6liWO6rLgxQRIF/lsKZRv7vjkhggPMbuc8weBi1zdy0AygGsrCPbvAW9PwCMcKRg
7+ioE9YfQQ2pSw6N1ImuhFOLAYt4zbRkIAGW1eSwRv/hapG5Cl5WEVWPsZUwcRYAkTnZo+FMU0x+
/+j3WEHVALxKQv2wcFh+hefOWsJVwKE8h6dZgSwdRJyGYSV+H8at1tH43weqfgJLcAHf8+/EJ1R5
r5xSqqyWWqivzZpBVYYjIIPxrgVlrwoCtICkAZ1ZdmuX4oUZR0LyYKP91BSXCIARfN+h4cS+3/uN
YK5qU2y+vDp9fYEy4/2kBRUCn6EuL5ycX4yKe3M7SAU5pVRM/+6fHiAOjgeBUWz4nlboIngiLSuo
sfkMsKE2M7QGx1mVQG4fpXa1z9uZbwJlB2Qgvp8tOQj+W4n+UiDSkvhEoZo9fUq9qBmw+PeQ+Ep8
vd1LNBOikXUrbeQL8wyMVJkZD3lRaKbA/yjpQRCO0dnE3zn05Zn4i4ZnlOrm0WohD56whODZ2D4p
nbCB9gJM+8SK9r9tD1SfO4SwTg5S3OvVY7F2YS/h7UnlGKvzhgnhZ3dDE3zzSc0dycHuJH/OPbCw
BECaIcmbZ1qpTuXzKoNOMhaN+QrQ3tznU59ZrjBX+WNIZovdFg9JyUcJbDWQpWneA3t89cNUIEic
KaqtXi582T0xKLjOGLAlSWpmv0Xb4kPQOJ0t7OTifGlnutPYMWr/sY8pJiNMcJBgar2NhR/Q8X+W
Ez4nQJ1hlVyukjt1d39mSyxkGz1NI6RiPsl93EUwegDTXBYkt2VbLqAh3BuWA2W6uBzgQumuQn95
ly9oCIzBq/Ix9HXXG+51Lv1yz5gMKGzztGY5J4FyY5dnw+WvNMxnLYGsEoRNfYlXkwBJDHnl+48+
2sQqN2M+3hqCK0WPSpy9/FKNiqrQzmMaFJYzFumxBUPXxJTDZ6Yly1kk99iDruY4djW4gid9XGoi
S2NzJ047LTZeQ4JLUm7AuTOQHS+z1x3KkmC5W7464+HWagdSUzpXGIP33RumWfrlZxB1hAxA5PmT
yXUUYHEMf2mPh7IL2k25ePLITVjNTgTmyLvG91Pnt2VAMeAhuk3xRcuegpxBsIB7G5aXhAbrr0pf
2VWJckPOHtPcLY/61tW48OGCK1meKpu+uB39ytok/dJRz7TarHONqOeNMeJwyFywyb2UKFzD+IU9
OePPu05vZfHKR7igfUYsj8nBHNK6/5Kdv1Bblwsysq7GIZYvntwsFh+nKgFL5nziPSxc/+ib7BTY
Bi/MkqraR4AvtiweCIX3wBTDBQ5vUsPgfBk7FVdlZeakV86yMfygqJ6sdGixBbcZF0tE1unrbp0M
NDKp94smAoldD+fvavRyXQSSti/3ktbBCEpvZ5lFeTnOR7VBFGo1J+pUDcPCLbgusKo+Ijm5PLUs
lPRu3vUg0BNKb69/IEc/fFmDBreJypLvHdY+5jJ30Kb0evl2b4IDFJp4qqO3qs1M/hNXwzP2cM1h
7cQuvsx/ootOtYtCeUe1npPLrmFUTdHy3VVi6j+FosZiMQRPYQNl1WlN7GV7PIMEC9gsZwDlirc8
lJtA4jT3ubMqlh9nU2oZTVsrnQDBsDOxM3/dsT1+ndqOnYm50x9ZXW0YmiKmyw87GyJ6wpfuamHx
w6pN+mst9VD1WKUUJVbqRDpGDa+6IwfsZgs2CK6upc5ZJl+vvJRgBX4FM1i1AYGCAC9SPJmYovCd
VPl9DYjO62nT7JuAQEf4YzkB6s1vwknDrqdKRxSMSY5RGLhYmB131ZJQVykTokDYZ4Hv7jqGPBTR
neQPpfzPKKgOh4tWUnhDD+MLJHOv8IZwzhzU6r5oNzjwdUpX+1T4nqBE1nnZ0wTjdTz4BwxBolfp
bapYiCDYA2yRtciAPiLqd912BvRYrJxdi03doZfRbz8LhKfpy7Ahc54Cuj+5i7SO6Krz1skTmdSf
BX5K5yl92CayelExBjJDiZV5I7dnnw+dlgw08MOoDWgHZAiFy/h2EHFTk6g5wMDfqsEJgT5uF1su
09dDSE2U5WRPoEZTW+CZtTN1UjEXvdoCmurk8MYjPsSroqhkETG3M8jAOzZ6VsD9ssA3n4Tt+qjO
qRwOhJQLsYYq2g0AF061pdumOrxVIw9zsu1/BvQ4Xw2Kxo5Yd5Wd5PwDFVw/IKFYcIR5PhJaR6AW
HrvQ4Kfvxg6oC2W8F1ER3dC4LDqC5SwYt7TVW4xYKQCPLq9Uek+sO2brhmJL4pmmOsSSc2Qv099L
GwdlXA2x1eT3dy0vBngb3JGKIXAVed9kO4JG43HkMSAFDt9PLvtFWEBNRfExSIX0rKSu5eapY5/b
NMob/2yjAdHX2vhpBgj5iNVom4Jnxu6qwlUyOorBzEvolEb6XAZiFegulxZUX0T/oBdcbmfy9Ab4
ay39fmfnb50NDb1sNidBjxBAoebngLjW0me8WYQ3+7LnY7UhhpLVOX61y2nEXeN0axNKb/u8SYjP
sFiHMfAknujqt9jx8+DWFjj0hmaI6JtyfYrGrW5+g84ntwxPGK8GPXUW8rPCxwWKd60LE5AGUhEo
UIAM0Sc9swueTSohhwAFIcIqgCbc9VrkCKjSZ4QJH3N8adC7RI52VGl+w4XtZC6tHgDzUxX8P8df
Rp7pginG6FkwLjzqYSUpfl3RroAwzq7ufYaxDAkowXgpcCSFCyCIBmuBBO9HVOsnpWYyVXcl1kvl
szcF4VEwFleNZZW3J9sY2SweH2AdGOWbd2ygFVRL18V2Ws2/16yhtyDaiPrzvqzu6qI1rpnYmLVO
k4ESNBYmAZ2Q7GqMKTa6oTPWkRh7utnuzmrXkqFh3t4PbjQwPe4+aM5L3KYWwckxheWmWP0JRv/4
UgeA7S3KJd/0mbm1kPmgpqOF2952OhPDa5LOJ4RZBOl7GGGZ0HdwQQUGPIGiEDB4lVA+wA4g2sW0
s9wEuNCoEU9Xab+6y8VNaG6ZoyWwl1PfpmwfO4OhEehHSlzbLkyZ7dUz8ii//Tb7tQcKMWzZ7X6s
IyrjMbPV2iIw+r369Is3wgktGl6TlrV+gPRy5gI7QgOulUnPgatoQxQGHDcmNYADV1OixacYxKxO
gIk/+G0TfK4p+O5jJHziP+upL201UBhZA+xWx4IKfy5vXTzLNs/3FR3tUV/dAVgoBWMbjmQigRPf
iALdmvGRrdezYHDNj6VUu6jNz2wVsPqoGRhPofQiSE54UkaFZfNXPxcuqlr1hsUlKqReBPov4DmC
ZA78IqE0QwZNuZ4l43hKYJO1dEKI3FVPfvmqaVOmvNOeZBEnLtBYstLmeGXCk2M0kp3351Y3ptqo
KvbUG9J8EZ+k43QALpJOpn/hxhba7uLFVUEbjQw3a3dzZxuz3sJXYqa+9/uNHI/wdE+aCqYFpyYg
eFGN9TH+s6nk2QebBrn35+1h4LVo3ELseMfyuNoUVWUZBDHREZVFf4oROClQmLq0MWC4oMdbSCme
TelHt6RAoOLsAx6M8YacIZedjIjtC2a4EjANE4JmfEk9nxETVHwYwLOP7kAXl85ImDn1oRJQZEzw
YlDA/8G4y8qGqeOWzaLsMh6QSqWN51XuMsyKFE/b1AOK7eyxHqqxp5UglAtbn6nl7uHWxSZMPQN5
gU0LJ3WfmpVvE+sHvj09TwkXgCmO1NA+TYgzn6kT+Cftsib3ZYQvc9ymkXEIZYVpYVA5i2eFINMd
r3Jz5rA3AhPT/SeO+t5FEW2Wv7pBiEISFDnZ3icWYDdeWIpdb4Vb2yLsfmYtylOwqB+kfp948sXq
Il6OfA5g61xibGv4jOpBATmQc7YJxdx+eHjp8dslKQ2sN0ZTTYX1iLpmoqVKVSFqGkky43MIotNn
66OuWi5Befbgiw1ZzhV5mFm0VwpTusrMgeNavS7bOtQ9MrZoWw9OqywDQe9+nxvIXfN1X8xwve4t
RLn9Oo3RmGRuZ7SOLyYwdTk2HhVeNigNNdD/j7aYdMyRUDDNvcif/ITl62OB8lJRZRXO85jihTP9
svnIQtnX8AMo3yXB8M5yCZf4g5ij3Dchuu0PbCRd3ZwzmhqtnSokPLNxQHW9VESQv6GAMBB9kqXM
z4ABLYQpPD4OPIQBJGgN8207qjcxThKy0yS/jqrbwbIRKG8mmnhnWqqiX0C4cyu+3nyjQsRsiXKh
8/Fk30Ah+fIb34MYyxQYKCAliZBFxJjnZxX8BPPIcMPoZMzt2lYWCIYtU5/YYS4e44df2paYvj3s
EU7fSjHUwcIL0ZWslAEe/KYVQO3NCr8DrzrJdGfi4KPqa9WU9RPyQT3vLsCGDv2GEgB0zr+CVLXm
81VBlHeuTjdGfzkrHvDKAQdtK7vGD/3NACGSf16W8oxFK9nPiKjzd5JQ7JLQ27FrBlCBpFZnZ7Pf
LBd+IfcueO7YRMexwaHwfsj2Cs4UhOPzzG59PXdEVMtlfGE2S1adgv5wywnfyYcYzDl2Ls9SLQrZ
CM9MjYmumZN1E1p2lb6SkCIwYkf1s3v4oLQTP9rPEIQgrupUYA3wQLo4exuxzQHaTNftd0+tyNjI
rMuyFCOJPB2EDBnn9GyZWEZ/ox4/p+Ffrm0p9xYKbCaP+WB/loNtiMkSP14zMYfEEmfqCpTazzpP
rnUgCV0uA6dZJtFIFjD4griJK5YQ3d3zJnvzIODUyPW025hQWi6nRxuCjENQrNMZsNW/612Zuqir
0B5IbZM0ypZ/Oihw4qne29wRd5MPb8+9pla7USHEaG7g1E/jKCG0YwjIukBaMxRAynp0HFLf2ODU
orGLBh6IOmdM1s1o95wbcAVoi4KfqfWjG0eJ7nAHk74is7meiyInc8a792xWoizCeghvyrUEkf4V
j029dgk+DcRc9cs9tfB64khy4Jr2joYji+X2+AxY5f8fu2FRM4yxJNAgmbdrBtMZMUzfe128U7JO
eVQpYSLSv6S/YPaWCpp7tN7CB/64RID4bniLuazFIVoZ7Hq3Mq8KSZwTEFRVoO9Dyk/sX+Gmcgjz
YyNyct8sLrLzoktDW5scD+Z3wsFs2rnM6/AvaH510eQzKalc5PR5LdlRwLlbq6CdnS+RlUeAN3xz
hzWLXQgB/qOyA9FPE6z3CzBQRVnwhHrp+eurqwdG4gq6FE3SA4qtr+8m9guGSs4laU1u1KgR9yK5
IhJqc8MTDIbssI7jC3u7Zle3+dHh0MRcdu5M4DsEu31u8M+3Dk0JArWdQezL3v06p9DxrYSfM5Oq
3dgnSN2pBZSF8pWgJ8P/fgJLluil9rYDMLyO214WbMgLJvR+k7eP/PNTFRBVkVKrckxhCsXlbagr
ArK9gDv5VXxoYfdB/vMo6vWr0xxHT3jFkxSijoZQa1NNsealMvqdQEEzam0P37EpF0P5Hq5+59q8
iUjen+KnRexiy/ZNH1htVv3XDsXNfGtUJTIMg3wM6i8BwdUWEvxSHlO1MQ9+t1EfUH+MseXWeTzL
FZ+CZSrcDF9G2/NtGUyGIoACyBgPGeheJiG3Ql0AghgjQECdxJlQ6Dq44fcgQBP4tafIFKk7Dicg
MNrXr5+OP0Rn3pFSUgwxPO0fJMoH8QsnvLp02DK482+pCyPsUpa2ZEQgxMilhNcuJQp+cPMoDmrl
+Cpkh3KXN0icRHMzXV0rLXWVWOiJI9vJIOcctGDTjWLW8lmPp9LuAEpqIXFTw4Uu7YQamhROa9Y4
X1TaoWzYW/o6M9CbFc9c+mbqSMFS/WLtBDaILVpcF8acicfco7NrtPCAoJvfOKD5RHfEJMngrB7y
gJCs1kUxWm548xza0Qix4THwl9rBAkTDdnHETpWiM5ZGQ18LgSgoR+9htc4dbaASGOuuWnzVgint
A6wfOcCWs8ik5L5cqjC9+QDoy9YKK4nFiZ+z0N5MGdWfY99nyQV14q4tWOIKECoCGJK/24FTbY6r
RMisAiEO5BTA+444X6Z5tTfp+VxFO4Uvm2KgFLbjcjSac3PGyZsJAXJTq6BE6fAPZoocDtx59H/2
kmhxRNiJBHmdPWTPLGNIlMd7lb2AVPKUhEUOIjeuz9uYsZrt1EDo2agB2ME4DVxuzd4IUp8Gics2
KMP2qs3xNV8Dgm3UeE1eyu3lhaF9XbsZHLSBxiRF01+s6qE7DZefNC0NBio5QcLFhwlUud+OsJt+
wHzmyA6+k+KPustpJx/Bbfzxi5+ZFTROGi7igh38pwMzPNMRVwN0gkESKFQ6bwsinDaGWT7BJM/K
17OQ5pIKWpmOTDp6gf6W55hCvmliJpyI7IBgksLsq0DbT2l9sTErujTCnWb6RkeKSP20CvHIhTDK
1cyv9wrDOYBok7R12RyGGVrfTSqBJR7w4JYkcel/AFwkuMUv+4RuRXYHd81U6KaVBmtyhBq7V1P+
ijlSKKFFvGevEy4uATezlzsDsfdKMEAszVac1wEvLrM7JnIbwVABUDBQtP3YxaBHUcmjn0G41zTi
VGaHcojXNNqvA51aienamZZBwKsDFV9PMfHogBuaJ4k3FVMiFtQo8NIycVCdjFBMCk8eJPgVl9ew
CyyRQgk+NDtdKNdePNtpbNl68hQXA614bfPl+ugnIM5eJPONIuTTgI/xRoWJGr1rhXFP1LvhIIFa
Tg7GexjedQ4mxwAouOlQBFTnc6/7FqVWtjeeP2Lrp0EBFTppKzHcRtNGVY/8zvG4HoTJ3ixrmrlI
ayyiuAUyXhJTaT+gSVfHh24+Zv4ffuChQKPuG9PyK/kU+CeSsR44WilLGiK1FOkFFVTEGfw5ZmNy
fMQY3wQ0m2BTBfyvDwp1dolJZJfNU48iQmbBiWJcvdyMKvi5Y6OapPgQ/1/UVpX8eQv8pD0FfhRA
uWV5jVsUPZ84R+ofNYjhUx9KRhOW239isfWLW42os8K4cZyplvZBA5UoQR/0ZKWuq8jD1HeP3q4S
zwFnGSkN0wMwDc62jsOFYhWIbtPuUWRQ3qYf99K9tBtHXHnMq+d/cs8FA/0H97/dkfQ+KUHx18de
0FF/WkeFO3h/03O+z/XbZVahgkdAlymWWsQvObN0RQ6b/9CmmpcuOW6lS25KPbBZRND9MsNYmELu
x9NEYl7jAAQ5D6Xg+ASvB719O20haXQejGru3d/wFT6XDjtH63usmA3/PcbYb7mPjxo424mkfZxF
SbE4ChxxWDn4MsJ1UF/FqPuGVzoo3jvLSUMMbwomnAHyexr0tBF42h1EZV77Ohlw+nOTT+M5FwKe
A4DmqqwwLF27t43O0+Tja1MC5feb8sAEZPnk/D60jgGYPs0QPb1hSZtAT9fTvsRyU8PtBPzvLdvK
yF3/cJ6j/qH5vL5vNryht7SPjjco5r+AO6YTyxshulQGdfA5+lPZzsq9IiPzDyjr93HzsW1/mg9e
fROZYXgi/dNWY9ACnfcDmmdpd8OKXkIZfk0AG2UQhrU4x561y3ttRlaYuyi8a14BoWettr4iiphp
Iyu5LUhZByTs5ve8Su+2K/cc/QsmR6HHCvQR7vN2lSOdINjiDAr+RUjG29EG5oraaOtczePxxEhi
Yl+95HcGCooGJxyfkAb8XZMZzrFurdfgRrPEi3wIg7unt2sH5Ukpn0a8+jWIXgWuonvEo1rNSDyy
P1EsGkSV1Zu/hhJjtVxTMDGKYZQzZHpliFefdIxtf1NeDmXXnDgD9bn42QOgudRI+Z1q/0DzguZn
FbcowQ8fuSezvm6FK/GyTjIfJxkSiqD+HnF5d3G2B18gZVgi8ItZgIcLy+sdqYTXeZ7sOHAmlPaI
ZEFJW2QkH5IaV+5yIX2xftPwr89XoePJgS2sADCcrUI7Oc0MSbSfZzdhSG1NPYQj9UzFJF8DbLBi
QCUiFXmmidF/13FP2SAd8yFXPzpcTuCJU33CHO2xulfXZmB2fkFyc3lqqfNOHCoTac97+MXWnv3a
Q0OI5wqsMEmdPrqHzU+UDIchO8QdGs1hrJHK4Xxba21Xz1nIwVEMW2ZGKMyHDgnC1ajEFV5WmZF5
pc00CtuDcH5DwoTJG7DVdzo4WJG9qzCX8quiOQCeKhu5bFIhp1BG9uuf0yDYpbNr11IXfEpHc1K8
RXHkhysf5uU22j8UlSEQuQCk/b0muJ5f40MwLfaYS9uwR4HybJ4nyeTpqwKLJapPvjcgVG+ufAjS
nZZCvMPzMBU93VBiDYVwatAsS6b0vC1H/AMdomH+UfHmm4ZYimwLbYyy7BR7EnZIw+BW3dZy4pzc
pL4SkW/8lo5waQXVY92x7oUOhYI0QOJ+/o2cMp0L81gTQdv6423zrRGHzMFwCjbW4L66tYIFj8Za
o678zdImwMhlJNu0J2xeSwnE8ESgtY9XNExOZlAnVX92aRwnKovhi5ASBuEFV5XBlWr0dZf1wyA3
0GglJQtAC2xRp9qIPNzuH3qK5Twf9xlNOy+KEilW8Y1RslPMbsI3qy/Lg7EZusZ2zq0jFHPtzW7g
5hVR9xMTH4M+KzV6dF0SDEUXVC8tjvNtItCtMPNdRJsk3CqqjuszgEEOiVzJ7pPZRUeqE8faFgxg
WjZCEpgUPLrzh5dPa6tYhHig25v1UsYmftTdhzCaFx88TVT5uP/1Nl+X8cQXjYbUrljbB+adk08m
nHD9QU19xsE46aOJ0C+v2wPx408phBCA2d7CqmYu78twZsbGBiyJ8wTiC20m7MMqZnpIDOnNg6yh
uANVREE8cVQQUKGgyQVYBhO+hvfaucTcJBXcx2AztcYat80RK286PuM0Yc/tVSWEmvcf+ViC51NS
btGkO785B7lUTY3awj70VElGZ6FezniFOowQce/YRdWbyUTrSMDN05mvP2VYqf5Tq/exVh1YmslA
C7ttX1+srnL2lIixPnd2UQrLq9Gc6hlruY4DeGnqW1zL3YYKPQjna+fdBFMDXLbuypk3EEmpSXgx
il/h77OxFPC4ce8LHUPGzOULBgkbwyLd/VFZk3k7huUCFCih1gFQy8qH8+LS7tOth7KlfQ2o9Va0
wE/N79Asp9J6nIPDcrpag31w2n4OMlMwuL0DQ9teAtas4WX1aZkhtPUffSP5pt55wsLmt4xc2yGf
8cFff0zbVReySg8DGS8ItHq87JRIyhAIv915r4Dqnnj6nSqP2p7wkIRCypP7bwMrKqPyIlCsO/HJ
gsBKpCr2jisV7/MzybVT5J6KsL/Ivm71gBG7BGxWae1Xsxm2AAzYuz1mQgHlIeyn62m9miEPCgGf
DnWXaBj85eKqit+jEfrhVcJuePPMk6pAEzkJ6QF44PxaXr1ZEsrzrKgLRw3hV9nnl5hEvt9Sjs2l
mUev2v08mGROZB+1WHa8KHZWVxDN2WE6tgn1yuuJwrB/iOlrz4Fj8RpaNIvhYZRKHvTep6o0e/hL
a79oYdrXgFvuAgnDVj0dY4ztg5KEkg365WoJC0g74NAAkkosc5AOE/cHef9lMrzCNaTtgUjADAXY
nDsaaGTN6rHuPcnxPibaCcORUJT7d3sKG5zJU5UaR7RdSByaFSWQu6dhdmE7DCb3bugIHju+iU4z
cayvjtBFtECD/pcZXtCLAD2y6eSms9DR0Uph40HRMKhvTZnH39slbp+RyHeB7Wlx3DZJ1J3PdUyr
TI2scfCkD6zgy+49feA46/G4KEwCgPepT5t8q69mKTQMt2fd+GVBjq4Vnix7xCs8mhrkTTG+xY+D
9E64C9NeHd8tJt+069WdidtTKHoqAzasoqp31D0ei/kZqFePgeiewC/wrh7wdEEgB5lBoZ5XJeSB
2w4XpC7IZqRmvoAHd6x1tgRZT3+jzw//PCpEp84WL50mn5AaVBcW83oZEEV263JYfH62wAI8hnnT
yMf76a+hswlKqx0DTgL/PXzIczHLpnXSGJ9zVQDLJmeOKhFqNkzU6d37HvsHyog5LHlpxkvWFRDB
q3KqZNjmliFVy/bKBdJIvl1Sm/Vn7AFSrnJhaBQwAqeHezp5qJwXCEoz/OpH+Sxz+fL2M0xA2NDY
WXoe4XKkcbdEvMCmphWzt0r5Ux0KrnuWdfPBm1skQviY8Cxe7Px3Yoyo311uDkOEawGzTwtclJmo
ys5RcXpgZC7DIBeYewyA4PIm87FtYHksnhPXfD2TGyL6IW9iXT+K1JBpa2g1zAS9KYH+tsdaRpRx
+ZW3g8/Uo5IyXd100D+iD+AIC6j0XKa0dDHS5KbSCWc1gEH6+AbG0WbJZZUpdEt5JH3ztyt+tMNQ
PpWUOOGKl7L79qqSxYEjxVNAqMlw4VjAkGdknWCPhPLjYQjqX5rTXojM8ajKsffIuCOhw+QyMMe2
itItY6sNuKOHcAIbVxRZxkeubDYet2Fm342+JgMJVFgoI2Ln57846Hsv6a3c8pFtrtJIo0ngAxGW
FtZkGenglGN7j7qGtxB2u5glAeqvijDne8/FYRpfkZqIgSWbfSb2WNayfcR3Huc6c/O/JVG4FLmf
3zkKR99V75HdUDZOF60xrFYBEBe9RFCka8f/H1DM8pqBrMkKdHpMhrl50mhQG4GcM9lhxq/VHF7B
V86VaaIcHiK+y33aOac2eHG6vbHOAhOHe+yYvlKUMaPJVeeYjxEjbjapFVXmxUU2l+a0Q134D0wP
pKcmRQzvCDwg3oCg80xtnzbsj2+eODzZaDA9XkrGe3MNTpdsDlvHSL+RZxjYqo/2GyX62UBA7moU
6+11UyTbZM+FPuwMViPAUKyyZiVwn4Vdn5nLTRnmNo6EEbhRXz2V9fUjqpxNoIACmTLsIyYnKwaa
ZFDxFQ9J8LjclG8ic5oyZTEvpkjZkeRDeijh1BnG9Lamf+bflscWraXgfnktqLvQM9c7to0H8Zov
xETZ3ysWNYYf1OhZE4bJ+aZTEq/885B07Cg9bTqM2SZeRWj1yxPso1RSRZIpZgvTGXfGVGtf1wVP
WNXQg2VgR7Zig7nu3mTlFdLilVUhavt5Kzgy0HrefCQ4rHlqq1DtePH3l57wASRvzORpc8nuVrF2
xFQWnA4Ck+CAaiuHw/en56ARlkxVWbFzoxAHVH1WDf0a3A1ukBHe7q8EZTyG5U3ckT/WdZKng1xF
qEl5oFzfe9mdJ1mzz0dl7jazQ5wFEi/Ew6wZKgztVCYMKyQNt3E8VYM5TpMw/e9IRdcEg9M0O123
oX7o6hxITqAoF+aHWzp6uFKli0rMk/U+2oWlJ0sFD4/xOeWeqM6B2QhQJgHqFbwUyz4mtp68KrUu
ns5ttL3QdUpAPbPt4egopS4VhTXZ9k7Hlmh2pEn6y4l/xCSjIaZGlZAtZanSEC+6olNn88NBLVXS
12lbsbPkZZWbNNV+Y2xsD0Cn5cQ0Ptr3bRZl0gzt/KrOXx3lX0QkxOD3JvFL+CNFNE8t1HORFb7w
fJCCpA+Q45x9D+ZNKWVx/bKXufuCwk68Oz4y5YJ63as0oadbqo1uSXisuIr4vo7piLmvmh3TYvvr
DafHbCOyKHtgQCiS8xFF5CI//cFyScuPaDvT88yyiUUD54+/iobK83bX0e5pgvriXy+hs2KXGy/0
f4FF7DdlGexYBId5a6G4BNtzi2yUmAS/JXMlvbyM7RsmjsSZ+5oQxJMgoUHLxXlbzrIW19hKEcIg
l5uqU8g8u43UUyGrqxVoiJXGbhE85cs1dLBQqPfAzcj3Yg2txUKXyToeiEVxNW4g+nE2TeTXZDyk
hes9Sx8qgaJxbL4TBmUnqvI7qO6vOdQnK/n2i/+M1Oooa6ErWnjb51vzOvsV5iBxRz7V8RSlFyS2
VFLwR1FGlzscxC00PxMxg9Ob/X4tACu5o+k45KTKJ1z3ruYR9/bJT2+8/t1xxWxlhXxqOQ5yfsr6
Xw31/YW9c/AXMvHWvYheJnJHT65lEmFFIs7JrrlJzB2EDBYXeBbAGRDnn/GPqlJxSXypnazOJ2f5
GJsiAJhTlSzGfKXRiz9rqhX0aPfrQWf8aNcZsSIKD6xHbfWpODc+c9HqaLQ+hS5MPrbj/cD2hNUw
ngHNBDGcY1ywgZBREJooRtTukeUobdodRm8ArvchnlQyVLqLONmg3ovyzsSfNCQ4DoJ6dP1xLMdO
wJlbEplRJtRlY8wwAV4S5JlDW1lGrh5zsW+TwBn54A6oIt+TJQV72GKlGdVq2tl7gEbm7a+EYeXT
CBV5NLXEHcUsS3Gl5RYMd/RRsEDisngXjIEUBXutU7ZAEK5fTRd6Kcw3EcGE+0OwnpjcXtI4ewkR
I9gIG0HUIVoDZW/2+2sAvPxOWvnt0BChakwNTa88b17aHnHA8nD4Wbv3JnJLDwSaYQSjPgbYZUFX
Dw3aEAiro6SDwkkQslVz6UzBfb5ICXsCA+uHS4fb/L1SMRm4IKQPwLgTXkifJX4YfhkKDMJO8GCa
eubWqCQxjarLyxonArbDodutDAIF47Px1lw8EAMjteRGbm24593bBj3gnBohvkj7uwTzU1RyBryD
ng6HNJrtgdZ3OMXXSIf7huW9vKGDwtGp3iDv8G8QsWD1tcXHKzs/ZBvtgJYtcDPJLH8HZvSOPI0O
R/Mbp5LTxutmQUoKwk+sfaN0D8+EsfWATP/N/RyZXXELHqEJkZvaaU9bftI0DUEKh3sl3rK7UzU1
2U47NXVh06KL0baWnQzHud8VUj4HxIYJ8r+rR1qVhQuRbvRBoohHu0m2yr8lh/qXhJrgKwJiDmNv
ABNp8RojZX0cpirTLWDqy6Xd1ZaJpMfF1bfekp2OEzCTwZ1AXFrk8uNEi96ju/VLYc3uDTDx0VY1
7KESFLsOM1rwmhwyDwCjcMHwFfDmjt+i9n/HL6lOv1b66AOEmrZ657gJA032zF52ZQTUIBRJV37o
zzU9cLX7ceH4gVk42XW7VRwwZ25Q3TpC+DYoRUXlOB/euGYEoGXucXdoQkWxvzxP/eBDDfn7EZnD
JElzd7eckaI1EXBwU9QruFpEqHRrEPvJ9IfK25P5L5FuXzVPqI1m/KLEGSvQSiWbcWZ6IUbVo5gN
hen6jO5f0IP165wv1SiFIBnBZMqsPU+ZOFSctZPgpn0zdOyzNgHFKVfOVWlpY+NNtDjZoQaCcQ9r
UuXCza3z5iilXdPM0LRNBG/IelCCJ5SyIlgCnPV1wzCgNOmQJxgQFFQYN7DdrPwIkBunsP4ICMAw
UKWM5ItgZd4qvK9FiXltUUp/wDIBzxxTYi3UJnkqqx3Y/YIKFtUMfAQPFcCAVESfk1+JFnacchGZ
Ktax9IaNVWGkCIcrc/5oQ87S5IAjadrV78fsL9ksZAfsNXBLOadoVLWGplmQMzU1eZa+AXmPE3zy
1f2HhtCkfwPXnV5we3cgJb2hL/Jcmrge2DhaRxeflYQLo+pKLPLvzJY8nq7h+bmjH4IgSgDvmB8s
edeRy1/DtMXiavCOAVaUUsfZfNOZTVvLuBvJlDCrU2akqqCwmFCGCoGmNcTIk5F9CnDm7REGK+dO
A0FEU2+lpthH9UfitiHumcherI24znOIaGL0/5vDmhN7PsCYbxf9i2RazWjWPGtCmF/EHLAvp24c
luqtTokRcbZfCW/hbGjkfRTzczsJ2o9eYpal2+AJUPGCq9Y/z145qHrIt0f98GaYhj7XW5lprLHX
phXbZAsbuRehJWMCMhPvq/ZLKW9eEMjfpW1o+fVGOzMsIlRkopzQmHqke0QwTeCVuj8mm1U8V7ny
dsFP42tdz567J6PsMpa5w3e1I0wR5VCR3MnDL55UqCNNmvjDkkIy5kDP2VtZG9MX32LYvysn2QCx
XiDlJaGTC3vONCuJsGNg32cC2tbuld2M/LG80UocqxwkH2B2vfIXeBFmvD8YJbQXYiHHX21mzObc
7Yh5yf7HE9aCDZYsrygBcez518+FnhyJjDec3NIxiQgA4mu5MCD6s4yEW0d1xsPa6DQbyricTzP9
ruY5eiIzusWzNy7K4c18IPTCEqN3OY9SWFt8VAxTgZj5qIq0dsH+5rXwU41uE+YIPK1IdT709HRp
TxWm+l62BVkrt7fUg1zHyp/axdy3zvim8zjTbHNzYXlELXVT1WOivsIphhoLQu7Pbg3MeGIHX91D
nL0C+eELgqCm5ebSK4M35CAfBgxI2guMa5T/NhpUlaNGM9j6du7Lu/q9yQID+odtp7P8NSN0EkOd
6e6hyxB2MPw7B0bMwi/k2J9v9EWezYymlTtoJTINnc7Kp396jd/4bXxP1j8toNdo+5IYjcSpcVHQ
ohyAzMxrWZYmJ/u88srUOHlPdm/EYuY+Lj8dd2tyRKi9MtHBAc+LPqs33UKfmHwtsgoBEwommixq
sKLhx/kP3TC7f1GJR/L7b+suf7aBzIEiJPRm9hK1gu2GW6p45eVtQTrFYQl70VBb7JAUXlstdaav
fd1bKlS7NhFQoDELKbtNn8aeDY2jkdEZBC9OYoXIeNzcfiocnodD13XmEABHjaM4UtRDFOi/kxT5
bGFAwGX2DbCYpw2CEV2TT9MCcdoFvIlnU92W+8lZR9MuHEZ6n09KytUFgrpA6yM1ngo60c/roxib
8x8JER3rFIwvS4Z7Nfuqzahv3Ffhay4Szgyli1FydQpMs1CnjPbOkhSOCNUJI9Pgs9bA4MIDIV0/
w5DuQaNrQJWsVriGMRl11EYbid5VDdoBkJteQw1IsCGzVPtxzhYzqvzQlgwD9GhvLrjNQfKuwdj1
ugdIBz42T2cWPUC/QtY1Gldd+61YzQB+kOcJyaFP4uvs0jluRPL7W6f023y8M3mYpLbDFw65tjcG
4H9WSat/i38gL0YQWNWb3E3qkjQxtJJEHXg8NzV6vceWCIVfkubzkdiX10ksX6GVAjdPdOMRDQyS
PIz0hqkqBcTOKuHDuzhTnlSrv2D3imF7y4ygpOVPiaiZjJKCusBU3K9NeTw2RyaC3YMRYTu9nlTY
0E2toRrKkIZdMi9e7Z/j4522zVuCblVtoylUmvJBAYwGCZSB8biZHaE2HED380Dav2BUtvtmP/A+
gqCZDV5FPBC8N0utTfCahGXNNLFn0pbT4tdzCtw6kQoJrfwVH6f4aJfkvxPPUCMlmCnow2DtrKpY
M7QMruBUQV/KYIE2KE02mOgR0dnxIIwEn8L5RPa2/9QMpEB/+VgU4hDcWC5Fl9C+ZCmUTa2nsg0K
KZSMNzMP+wZG33OkQatqBvOB9T2KXYJyb8qBe1yUeCG1giOTHQud+Zp0awkRAzW1XcUhatY0F9GA
uQOUKvJQ6qBVDJ6xC3oqpzZ2DIgr5uaNkCNWcQmyMXaPGUKVAF3+EalLqhBkHssMjqnLSmgd+kb7
mKixSk+c/+lWMVsb7/jhzGsaj2JQmajwUts6PFToH3FACob1lK04aqbnCJ3yS1G2iRKuHwxX6L/a
iN1yL1mr+l0JVsgEf6+Xw8BbmexFhHY/4uHc5Yo1YiEGiV2R/NjK2Y6ci/yYBNF/FLcLoO+zoP+I
TDDtV05JrBGu6yMdHZog/sWR8fdqDh/Vbl0cdEf9cblSB9FDKz+XgJNhzaN/yh9nb0I76EyHZwml
Zg3tsumd9zuRfL1N9rr43ITWbxTCjmUS1Io5dyWG+Il2u3ESUehC80acXZ6Y6q7geB576tRT9jnU
waaygbAMCpEAEZIeT/+DR/R5zqtOwRXRC5Vym+2wJSNgQ2v1LMJNv3/oeW3cyFCUZiUPDnY0AKwq
sfbmJM5/QqHLI82euQw+8ShsKvvMuFWZsSLjE1BkYPsfKwcG6T6XS2xBXfUAatI4ih6vzflC+s4D
qNODM0WaZom72fo3tHbxknUjiaK9VorwIJ5eM/6bYQoeV7vwro6s4paeShJXvptgtjVZF5wyqiH4
Uidd4ap0xCyrKWPYetrE22CJy01VFmxQlLDDdKAXl6dRW+cS9gNvfMoh9EaOnyji5TrN88VBGfCh
dZCb/wYTi1wydsJkX4obVb24GmO1wvOs/k+jmBu2TJ0+HbnJFPP/uO0ZP3/skTYXr85LkciVN/7W
XFTGL9ZVpOvLfD33g5ry4YCCDDNgIv3y9u0nmeFJCVqmj0BLIy5x00ncY6LShvYK6UfLH26LUJ//
m1lkL/WZu7FvrETK6wHiAEi5L1IqXFyOzyC8+REXY5j8r10eQDoPmsnfdcyYH9UQ4fMSON8KpPjZ
J1N/Jhp2czBp54nK04ncDyX1w9sTT7YkjRxO20AmMYNn5PGvpcbQ4pCud/7oofzfKb7WCC2wfLIh
LMLyRibkoXG9giDhRuTDAa/xURtk1swN5oqg+OJe7vwz/KRdQZvFCHNA2tsh4mAK93RfECi9tPbP
B+Yk4/zbq0zm59fOQJ+RON0KEKiTR7e9jPNlgK5v/Pc6gy+nXkmmD4Bxqq5S+0z6i8havE97kf+P
P15dPM1AUhpt2wx6DS02NTVbsuaUAw35tosh8Ndj33YlN/3vSMalfWw6vIfF6pFGMSoe9UuCUZT9
zrAb4W7kcjuMJczlDWgPtg1c1vKtBJIfFKbOb1SuCB6HgbetuS4f9aYgx7q+hhzEgqi9+6ADTpH/
Le7eEVLKf1zvmtXyi0GqGj/GCemClm+g7y0YAr0u1tF3Tdu8fKgcx7TKDyyzV1EpFdr8fq2pUYc2
WX0IIfremSoU05aAjPhN6+8nf/zEAB8ibRofSaoOGWJDdYF6tflqUj6KcjEWx3GaNcF10hqS1Yo5
mWWW/vbltIc0/pMiQV9tNixgmUbsT7dWVxq+uT6x2UvegDzlt0kdf/GIJXoP1m0pNFhik0YrcLY+
jmtPQQjiULR6U3nEemVkYleeFhkQptcMaL11JooCjLtUVf92O0FN46ngjnE1jL8+wMI3xDzpqc5b
DiHPs9UILiBs96M7zRCPUDUrwqdL2nHw7JT06nYWQ5Cvn8NtrXCKoz1sEOz87RD1r6sBdNYFv5uO
sHJQmXYjPYPmIBMjnO1tYXBepCLV3DENvqy/ZZG+seQ2CNH0ZOfq2PptkyW37z35eqUc8FnIiBy2
yCmd0b20NkRiVdg2xS0v7+70+jxUxXJRbSyQjZOBUMDgxr6aoVLHmUFbpxxErFl60P7FsG737TAX
eDSB6ke/MTSzIDIFT0hQO4q0O2F7xzFNSQ8LB3mLqFFvrOlF2aLKDeLizoUxiGn9eJgGqula0glh
5awin2xkGXnSiR+dSVYzAy1qfUp7jk63Ykl42hYL4TkHPeBnVyeRz0iIKW6TZ6SSjnr+XutclZcD
tRns4mD9XNjqMm9XHbZRcihKqRvH13n2PUxMVzhLQzzz8nLTaB+1h4EKuGL+PpNNzWiHiEr+PuW/
GL2g8HiPDFBwc+4WqVsl2aKHCoJdbmP8ELNLlyGY6qLGIVmNKsN93TrOyH0xzbeWAVyXgOy/eyzF
wdMv0sP2grhjZdriEDiCM2QC9Sw06AGWTqsN2WrmrQGwHDiZEby+Vk3vANfFwOUxihRFwZMFt8nX
KPQReT+M0yautSoL/99HypxFNFY7iLnyMQG0124VmMUTW8K1+4mo8Xefb20n0FXbsHAiKOfXVIS3
1e7Tbxwr0infdbJjg/M2r3zluaElgdo/FlDtaY4EmK+GR0coX7rZmUl8lO97qO2nD5A/4kGnABNX
lBEDJ7NBh6WaPv65kQkQfvMi98g5h8ij2rX8EAlku5qxqTZw62vmPlbKdicMx+MOUKMyBNndjkcx
LKWvr8NClCrcyJ1v5NOtMakJ6+zF2AHHP5NTe9mYJu8uTYpAj0XThkYa4ClroRGVUcuFQCyFPC+1
WbV5IU8fNFUPpUW32xXtDbXQb1461HxKzC1pWfKqdZv4bFABEojFKpukMmn5ZOovJyrtPPwgGvzC
PexckWowa9oxp5/oIR2jbn9Z+BILeuyY5ZA5LddTDO24hKOubvhnnvWC9+FuFlFNoRFG5HCd92Dx
wD6lvqXvd2b58w5m2h4uGr49OXFujnt612qMSvgBuVXprZUUjyEZwJYrh0epCGE/+7UOi7C9VF2n
84sINhFoJgA1Ct1VaAH82EsrmFFKiDqPmG8F1+KYRFqJ8dBmG2J4whGua+8DpCgjqOKl2e2bZfx0
sD6r6fCaQDlzbyzwh8baSpNuCofH2K1wqLRNCAZ/MFnyrMObl2s9bGyfWgsEvUWUkmXokE4RSB+P
R+JXt1NEx0PQJ2qug0nvMOL2ZDWN78hnyeYGhQP4U5HrvEmNpBc82OKj1Pe827FXUVPI7q7n5diN
/KzW2XDirPND//0PPgwX8/0i6m2eXjZsPRQIpk8JxUJ/4rfXHzRXhhtpQZi/7gM5alpGlZaHryRk
APZX+Ybupc6sq8W9ZJa23YgaHmxoIsoP666BhqMDebHiTegjoERF/8ygt39ylL8szrIy8usJTqSw
loHaTbsosjEdUub9m1vXpN2t5+2fbTsSUbPkTCzXr/9cQnRlxv+mqE+BGQx15DhyMn4YpvO3S3ff
VWXzyKO5vBWPfqDFY+EyjcVpesMXjx4LO2UtccUOivXpyUYCTCk6ASJBXAMpZawRUI5fOXmbZtLp
0818AIgLCP+vczzvA5/P9ZgMBxYdq8mpjdN5APqvWrSzuRsewYoVHBjmRF+8OY/jQqExLWXaHr8o
CP6/tdvCIRTvHLNQ4biBq66hqM6iV306d0Xs6lQK5rNVtLzqe4QSVsc+fEmswkS98SkLJZ5Zg0P/
JCunAYJ6gSPge1wfXRy0T+dAH3KV5Ua+IwtEy3Q3aJj+HNvE5D2i+w3zj6fISrUnRar1GnSVNznW
CHLsGRUNFj/hP5WeTlEi40t7aMuy1W//w60U/sk8tw1YqolVlfj+fmFZW5QdGyl5jLMGqpH8aOsG
Kl0eTJEDOkZfL9h5XQOtgVKdCJbvg+IsUz9dHkAWHGIOaWpvXh/dgW+p0Ubx9Bq7nPf9kmRKyaPj
I/KosmjsNApZDZsIe5YvnUi4Tyz8OjRGjDa1RTV8+/yq7spIy8wlYHuSeqaZsAZTAjNMbiqCLx93
Wl3IrfmTTqFvcpARjqEAuDnxAy2m5EQjwRxrDsOAmy6oLSA26UUis3/0kfYCxU979PwzOFeahkba
fbCyihzC1tvQu1lQM7vJlZAmIHkh/PHhNIr98B2rmkLCdg88jtv7YEf16CJ9YfcHxvGDfv/rB2+2
J8FoSvAqiQIN45sivW6f9zmPgRjxLvFuw36cc5hghQkZCb/LpbLNl7+Qb2TSkq1X2TEk/S6m2Bci
fneRCbEHY+9WoEiyXCJB5uPlQDCOj8YJiwxiV6rOBAxV0CtitdV6ZUq2/PhN7F1HmbhIIWEvnXB+
xl7ysMld/jwcoeneaKh2uKGi/KVdi7/CXjSs04DpM7nb0Smf/jKOKoFwUFPiPlvwcydirZ74irIH
s0VLfafnETbA4pMnnLCjovA0f8sct4DEpMkN5AIKiFvlMsd93iRjb7RQRW5yq2+afWErQzeXQnOH
ZsMNCpXrqZTH5USa4fcIkN+5vR0JpQLg/FiFku7MA1U0OiO9zpyj426dBCfMVCnuLEh/v0cvU2M7
N0mxPN2ruLddeR+W1A/cu6rfRnf5GuXAXsZxv5ahrpUf+truTpt2D/ekc8rTaANfi8zCzomaiKXl
taG9HKLfO3IOI+Tm4tMLwZSFtoGKdHqFJSNee6A62GPPUn795ZCtfWM07Z5VRjsNwl6QpYXlOIRD
CWF5Xox7Am1fIr+0x6+oSvtgZP0QE5P8+ZEiGkxGeu3GZlcodNH7Qf+PN7Qd2LaPgIiTF5sc1wgK
hKbXxl7Mqjz54flpcJEdgA4/SGr+gXZI3Ob9lvulVCNDT/a7TYqcTgSc0Ac78y//zqOpf41non+X
ZqGlC/mVBuCbo4Ke9vN1a/2OoxO6MUfAbvGKy94xu96tzyysNaLUSIqXNxOAI2AsOxuKcSUXBG7r
SAhbNdBFPOQFkI2mSTEAY+Oq+F3B3bDjsLmsoflarVrt8RB4TycYQrtpkyzA0gwBnMW9UIcH7gms
Vv+HardiIwpMSWyJF/prU1puZHZi5qH5jS/LrTDt2pkiPigwfYYOximDTrqnVl2hQ0Y2XiohDMkq
fEq/C7cB483ion8JP4OXw3RcoSkiD9PXN7LtcZl498123ASjYwG4fLomS+1P+g4ngRDD1zBIwFCH
EBP0EV07NwZnl6uf62QQ4OklMW9ZyGB3Tbl5HJADmI8BThNdN8vXenLqBNTw8vvncL6WFgaBFIc3
OcGE8yfh/62NNqgK7sKoNqh5J4WPzPIuIpoZyHrS6sTEJuMCs2IV4TT5pIRhFa/c4BYA9iZxOSCK
cw3VOrX4HkdG6z7m8JlXc4s4SqCmbmG3iO0vRqVItRZIkKIJk5FbFk+5G37pKw/EyO3AQRzGgahS
UAO1oN8zCxgbQNKAMg+3yfDqFFQmvA+C90DmwuF40oAItP+vebZ0h+VfKMgwcY46jMjb5bjYK1RL
z5JONe1v22sVLa1VE/jx3mnn/EgmMM6c9qKWfi13yMOzZSobdyB5WaP83N1rSpqHHk37/EUAj3F9
ygZiA3a1apyUQj8c6+5Gi4IgoFveB98uNwjXP61+qvI/QPy7NTVPDxaZNVS+4maEkAVjJQ7D1MYS
cwwJn5W8mMlcF9h6Fka4RuG+9xVbyJtgee768QQhdV1EFdLEjcj2+Um58Soy2RAVJaH+3anspbZf
ArPCUUN6GJkbtKEjIY3e/TyuqaYpTD3E2kHjLSwTdjfTC3dwVJi3glVci0tE9wtH1JF4BWq27zjN
xOTLEybRfTB9LKGYUY65Ra6Ze1Ms1cbU5NkQRiChE+rDvIJ5U6jxloob+Cq9aldbQBWeRYvo44+2
Wbq1VslYY+Jpm8mlRUlkhky1LQa3V9mwCibDgRd02Gue9PeDpvFCzAz3Sss5zgQxBae/T+nUCFIk
0j8iSESGKVSWuKy0I5XtjMLnx8Us5Hjuleiu3VwfZv9aTsMeJJ36vR+5/S2yQmTY8pjMF0UsIUdd
D9yWrMWOCVltNP+frzXEIaH8PClRVL4nXpvQcuDTRqLV76B2QNJAv+90rBbPC50dNbw1GqQW3mPP
0GFsRY8ywJgnaAzVBVN18JLd4G9xFMsvq0e43ck+KOSTHjKCFVhqiXpeka+kyV7oMgU+RKAdIC3S
C7UrVMiYA0diNlzpwZ9PMNXaU0FRYrHUqMTiBKgRtjhKrOn2r9kqT00drZtbw4T7jE814gOLOcwu
dsbrfDVheSx2zm07DB/WtIi7+yWTazgw7L7Xz5G0y4gF0kIa/5FObrg+inF2XAp5U3rdK86TowHW
wSAXX1ptQ6Tv5r6b/spuN/MuooWViqQQAYJIa1o8UTM4RonGXaNPL2Kj+k3JD9VAgsgE8lfduBIX
gWPU7Ca8u8ie5R+2rXIiMtah7jkOuttpnO2teBpIWYdTisZy5tCh2HKtZyDlwORKIspVPn31niM2
S2ptSV3H8iOAzPt7WGc3P5pXj9Vi8sQ0Lnrqmwom7NWT1SVz/Bda8dPYY779MUloBJr7HCjSjoW6
9Awq0ASpofKAQ5tgqNqvxeBiJ8KsLHmIm67KNxxUccp9FG7Y0z/M4gSHeyjPpMwPBEPr4r18HirI
vHQD7M0HE+qLb88uYz2IZglJKGv+9uUjRDM20Pcc9S5wp8FKDkDpqC1fbdcGgziQsGRA/oWKBH3b
OYdkhSIJZX5c5mXrsWVuLM/qG33CK1OMf08nZO0RhMJjJnpJWFgzmFENjPEpoS6Uuq1t+VWRqS0z
34P2Lk9hPBbDJDjOl8bm6MUnVjM5UzOSnYKj5K5WCYAmt0WOoQjRCYSLVbeYUdqB1rdXxiiy4cfj
s0S7bVPVLU18vMWc0MwyXKlliRVNg4u2po8e71Gn9stIYieMgN2r/FjHKff3/xvXa5KaN+asYz2W
Ah5FuzGDqt3kqqrQJjDri5AgP7/6kU9yc6rbEtx62/R9QW+GU1Y14BfHBZ3WRMT7TURrjKG1n4vQ
8s2RS5lC7wMmwNvDV/hnQjsfWcRx2n+359n9P9El8pvLMvYMajUOZN1l8qxuI/zaW/h+QEvyMmj8
VZvo4zXsaTTI7d13+aGfASC5cAhDv/P13pRNnbpo1ossFD4UpIPf9+b9Qp4DEXGizytvyXb+0iTg
cAru/V/7amqD54L6ldN8Xq3Tke0GoD+gzLGs429pHKof+rxSnsGRYKEWFLenfpHO/CnHQZdeLd6M
6vy1U59OTMrmTb+6HYFzeYVWE4G+FiWshrAfRBacAQ9wovUQyD5FnnM/+n2+0q7VJMG0jJpWHyH4
yyTDlOV0D4bvBpV1Y1+vuxaPhm89LqWZFRFZqfFlgO71Ozn3bgtzeH5B8eKEGoCcNGlu/k9r/cTp
8dqnrvAol9j24fdRpDVY9jkA+3wkitJWTNywC2izdxqiXUb+063FAEaOUhPxVjTppHhGqdDCGyRr
AXYbHnfzQnmTjJxKkVc79NCETWkhCcO5dIu/C4CqLFk9DKjXtoASB4eH1Z/xeBTeoshGaL0ybkAz
5j5FKWizzq6voq0vfVsmPKGMiCopD8VYtWpTMvAEt8rrldNLf8v0TxHsV6KNen4KuaTRW3+fseMY
VxCs7eM4W/lKY5ehPx4i215FjiQaE8NGeJlNjmWt80sizv5FaRK1EBiV2Zx1PRMyarBWDgJ70R6R
iTucocw2HbQRf5MnzJZqDBnKYK5KE9K5RWjbh+6xAX3mmSpUPdyLThxeSBtwFtfp9Oxjv9IIrRHE
VEC/P/Qx6fu+SR1Wcc/PpHndlGh0S5hBdO3Ktilyfar3OVaYvNWF/1IheqM71qP2oJ/5qN7ijWEP
2+eIMRMnXp1ZssQdj9yi1L72WfarFG1z6jByOAwhkM5Tqahv0q+1UUIwRhI+mIJtEsSh8wYu8jZf
HLbqoYS6Pqhl8I1IcWNi6xAHXhiQnkVYkSqYelVrWH5+5TIdok6wUOX30QXpjMzMBpVOVrSeYVOT
jODSgYClMwPyyKIP9PnyeigjUnezskixbFl4TBe+eMepbyV3s7tN7eYF8PXcX+I0PVYOXvXGRgJr
zI/Nq/6qJKYsdut9UnsHXTXOwEb8jyjMEFNPMU25W3rhOiqOS+X/5EvdqnCzNNgBR/XSIK5j356F
2hPLxnqXl2QENQThDN2hQ3ZLeBmwTtepPO3H7Pg4S78mBuvfJfl7Pn1B64MnpHJI99zFO7aOJZDu
SO9oFtlxRXMh45O4ND23VbpA33pXqEwGfddG6i5fbCv4yAmFZxw6iRU/L6AeFL3VJrw9/Usse1mj
UASNeVEZDemqgjkJS1XuzvoJOeLXByTkoSVQ3ngpI+nejWXg4QQOADQW9emuFE8GGzxuCqDH0jZJ
wOhol5MAkECbuaQvFDjFtCglGtRnbyhQTELv0vnXjz2cxPIli/zokWJXVC2HLsACimhPJGprD9b0
st4ddlTuMp8zGJXIK8KClMMMH9AzvYrmBg4MLgzhGdHqhvdNHjtRjzfbJ/dAfXL/XyCSJGTYIz7Q
rgjiCxuCWQ/narrdliD0Keh+b1a1oO8zIU/jM8lhyuiaDihaCgD3PE5lXGOTY+XqudQ9xtUHawTx
ghvHneb+HB4KjYDbxGvdw/z9GhSU/yeS08mjJLeH6rzdYG7n6iC0B3AQ1m/7I76SNDk0+YATjCLX
aLfi+LrqDTQfdOz1LKYoCYEFlxp/9JkJERqsbG/H2Bt0OwsG4Jx94NIk0DKSk6AQa01e0Cib6WCP
+DrxQievIKU2213lsGgOpiRBabbfIZ502eso/XlYwSDJqJ34k41WBtapw4RL9JtbhgF22yBnxlIU
xwyFTbplTn5G28p5aMeXR1JiqTH64DKMEl5/kBpTfKDqiCSZ4guH34HCXJYbqHiPLvH+7bdXv166
suICxHRhHVB0z8gBpS1JUaY6U4X3GkmHzvu6d21wJms9eH++ducWR0NkRqaYHssxvMw7GenuLNpQ
ob6EqoZEfp0PKTXfYd6teCp71d2TQuQpLj2G6jF54lWVRa8A/JHFwgg/H/K3ZUSc7xSpz9bqkcf5
9G4ziMPf5BM1Xb1Rr8B2RelI3eZlku+nW+LaCXA75H3ne/KVHe4B6qZX4nylIeYBxVUMppetsrAw
cSr9iZY8CBxqjefL9Wpf7rpTuNGbySYpkIBKw6q2VakANKyqlTWi9WxrA4iQJnvUMzNSM7Lq5dqf
+NSOmWP3PkX76EJ1MLTdCrkNWjqxrT9j27s+xFxCJ1kfd59g4YQmpa03UOZhOmmFjPpbhSfkmMcT
RaHIvAOCV3MoDUgykyIfxNSaopdAwYi5BLl51qmjFaPYpE1StEq0wkOoGTnGdF+vvbTnGSvlz3rk
dXLVUB4cWSytX/1Hxl0Ri7qOQRP7DVm/cSgIwec38RO4uM075HjuZfYTAWzrYZDXir8KHQNZmwEl
L1qFtE7GdTiZdueusldstfqeOlEatVhtsLL2oICKDZKywfREsLAQtOzoYHoNqWYyRV2PUQzWFXP5
3H0I1td7bJySE1/Qp4GdhXOdr06dmdP5VX3zUKNrhsMPXlO+LBLc2tgRrWy/WXmS2qq4oQKCCD3p
OM9UtexfqV/cqjdqLzEqoB6GnGj94ox+ioE3wxooy8aUYmEMZG05Tya5VBUfPsTSTXvMFnH7Ud2h
IXBZu3VagrydHDM3lnBpdNfavEZrSiR27NLht6cqEofS0b7VeUx1CZEbS2v7Dc296/1+xV5X7GEX
k9LRpAzTkDyGeymAOXxMbnynz62HkzNYi8wUShqfFZPbJtK63NOmqynry22hbnXRTWbFpr/5VgKu
Z3fN2TRLP54h2XxZVqYLu80i2UJtmcgb1Md6QBTROWy54AaOiZWwpLjX6cwKK1ihGh1Zj5Uz7VkJ
HtsvXQRH2GzZmYvW5CgFoMX9pD8BcdGKmxfqesAM5RE09P0ReHqGk6s7GKbZKAn9n4rBjCkUeqV5
g2XmROUku7AoLogq64Wwd691LURStrB/wcakVYG6KCIM0LVJNeOgdUIJkJpCj0gt8PthfGJ5E2YP
uFQ7Q/03AsQmgPi0f/Jax2aAGo8oNHG/E4p9QsAIPYrxNOtAz0r3heZ5KB6z1DLfyuhe8G5BgC8r
azCNHockLl3/W3vKyQzMI1Dpt03k60jRxIeOkO+LScMJ5K8srHNPNydIBMH9162Evy71nN1Hz2pT
A+VKBpz71c5MKMO0LEgcr6+15poc44u/If4PHY0ILU8uXQVfdUwfFaCzWT3yeDwjFrjlPTJQNRAL
ix2vZpsJZkeKCE9cDxV1m8VkqtjV1QsQ+D935Bf/DsflpMqAfMZi0Ik3nl05JpiTQRVxROvLRObX
Ud1L3zBztCYg7bBxv5JuFic8dVH2RCPOliNQ1pHclBnVHE4F1Xi0pXFchSVoEecXDblJ7zAbnouq
pRQAuCAnW3d3Fd94oeFBQmjpm5W3doANoXkTzFReqs3cmMYVRbE8x1H8+NLhrt4OLMYleLOmKYoZ
hQ1ACgw6UNSj/QGo9P3f9xqTKhEVTXzd6fqtzSqBiWZRsKIgOB4hyL0C+FJDU3yMeRlhKgRFB9C3
D/8+EvaLBOu9OYigP/H4INh9Qizt+2a9UKhYZ3EZw+vv6MMAVPxAqQ+jLQhorqKAD8UdRyb+A41B
YQBNOlHg0ByMiSv1NX2c5XRPU6VMQvQjZnqRfAoSMc06YHFxxwBbJcdOEr8lUDGAqVhlV3EzTpBR
6rN27SzcFIpFV53w95agGHEX4p2VpOUCehtaXBxIPnuonf9BLnRJtwFJ0K636ImOxsoukvNfcNeW
F//yCfpwxKojvJz03kLMaxB6XOsrHhoNMVxHmLtZVkbxIdDL+6nqJdygDkToya5+DzhwAFylPbs9
iqtNBMPr2M/7goqfiV7fggUw9mizUsFSwizEwklGYXxctF12ATXu/1kpHJx8Z6QGIbL9CnlycTAN
vIwEbgWMOXhqh/02x9Y/CG2b1l+i0FOmrBlaI11ApWdCpVNIc8TpgAEFQ5Rx7pErWntq21/3k87W
IOOVdZr8kAaLHX0Eu3H5esdq4U8GsUAB8EZKreRliFS2Nw9eFug9JVAi3Cqz0TLloAqf8TvOWCts
ZBQeSqtGO4KF5abJx0hcmTlOf73sm5ZEjxjzSZS+EtK0Ef6sGHhVZBgnMwB9+dTnLuMezT5MsVMR
wruHdLZ8zlIXw1V2bQKxgnSWf7Wb7l5aNJJ0m1zfaD2322e8VVAhTas+rR4+vDqCNersPfsbzCSp
8gAOXAkSxciA8/LWoVWPQ9KDQadBRGCEL1GAqj4/cK9I2AbXOzy6vjSWe72X4C203JLLHRgGsfRz
Bea4SkO1PETll5Rs8ZItt/ecVGofK+QLsgsGCS7GSuyZAu9K4BVF3xMD7BUG+bo+piAm5niEIPKt
z9u/cJ0Nh4uNbhkF47wWM9bY6vmMElDnEIN946lIDw2GWLBVR/SkGFrm98jhFdvqS9NwLSlfZE6F
Mww8T7YV12oMnjzmC1cEJi+x3+mAnNmgB73xNFMItJvUZyElSD2QUmQZlZ0Uu17vcSH3tmjAJutc
fDYQiw5zsbFjs2VuT8IZf6uhM148I5qZ/YjRlLTqEbZEYUjm5fqYPmFOTOo8qsI9J1lRxM1ucDxB
9CWR4oqd0MhxDavz82HnSiZWmO6MkcX10Xr7a5ToVahsXeN8r0iblo9KnuygOp81vJgEIvQQySy0
z9zT7a6ne4OKRxlOPyRtn2SQddsMfchiVKiOelxEFSShp8KVNO6bJpRaJ5wRGvtDTBR1IcAZUzjM
QZJDgiQqnnpfG6l/c4/zr3384wZDsgZeof9fZsiFyo6aVxjWL9cHFHSxuf8d3HalMQk4kwcKyaHZ
eLGtu/jR1nGGEn7xKddhwsPeJAq54pj2hD6K/uXcQq8X8yMOD4VD6fJizUwDMyrElY+VBMk+3DRR
MxrDPGUNH1QqYT0iWYpWyonCFyCPhj2yOYYZeYrZbtwBo9Um0rtz1QXq/VrHgdZg2QdhgfXLJI7M
wkZdYmZElvBF4UeLucZKmoV20hd0936v0tSU5PNYqd1ygrxKHQPMi5ntiYH5uwqUQjdJmPCi5ILq
8lmEn6Eojg5hP4eu89DLBheEk76i4ccw0crYul22UMDLE757EQOW0oAGdqS6dRuFoW//5cCZjzoe
rAaooObQJhy5igP1+PylifjY0UsyW4JlurZcUOftg70Wa4v4H08cDcYA3DboKxdMvqJyVoGSFHsY
hb32X1Mliz0gi+k8renMfOPf20E56GVbPXPHTFSdc8xGsQgV8dwjUtf8T2Z5ldGHzR4lgDeSwo6p
QmabxtNguyPveE/Wo9os2H0j9MN17CM8qRGbgoIbW/5v+W2Q9UREslSOALFhCKHVWzAikvgTP/jN
A6l7bmQAPYvp3o1ZwY8HEVNHxyVjO4gqYVyAmOx3Y0fD0N2U8U/bo6AleT6yJAuVoI4bXSY+dF2n
q17l10cVmt1TPaEZRarJEOm3ucYLG7YTx9YBBnb35cTT4UVC8kdZl+nWTq5JKl5d96GXP8DaLKqp
/W8m9wc61Da+tc3xfYR0UADvzu23oqSQP8JwRxU68WG+zW4ucHD02MGiFtQqGmgnByAqYOuFDhXI
3xOQmZDDJkfjeVCCPHSajaXGIxmA3PkyBqJsKrlua3MyXz92BKLfDP8Jouopu9trIAvdUYjiMloE
com0vNJo6CEHK3OoaSPXN30zM6v06UmHD8xyTGGDU3PnQ5Pt8SJNoEf+oD74+VxICr7SO4HVat+V
vv3aGNGBFpcw4fBvouh1iUbgYgt88M2SULR7X1FaKe3IrxY9xvKyDdik4itJ/3uix7HZKFjHSP+p
6h583eRzfJeBbWpw3YdV0GrrXMCPawbwJPWXHijZ7BcgD/2mfe9O1mEQAgPp1ko4uU0PoJatqe5j
PLtDUCyhJW8+1Mgzn/IpWoUrQVJxBqDPFrhGK78OzWZBzkPAoZ9+A1laPYyn5i8tAKAtSl/SUUCa
jLz944we3J9OseNo53xkEQ5dXcV3E1DlPexmo1Z28ot7tFi/crhF0QpYBHFm+4oUQzEv91JbX4HJ
PffyfiLmYxngFmdYf8eB1u9d3XzaYVTCmKlLYcMplmZTRqInwiGAtVFM/HKuxkcQOMpT4aBsTJ4j
gh0wG0Mjvr2WO79O3jeXhH1oTkq0MhLYUqp4COKDowCbSlgMawcUaISOq2pjkytGRRTsV90VCcSj
YNVGrwNF/TyAsyAtfjDyZw+tYiZmDP72TBiwCx8AGZd7xW2N2kV5n5HUfZWXU9bYjDu/Wj6+mTGn
4B8FSMDP/9foWEd3v/samZ4gkuM9Y3wF6Xu2lgfgGLz5B2bIIIzOXDL2/Av81qQL4Bg1rfOfQt8H
o14HTHWwOBRUVbVWbosxNh4PcBBkClwmdWtiSksBGn2chGTMhlgoechj3eIyM9O6InJh6xjAzDyJ
OqVtbMURMbINSfH4bhUxrqC+aNJSmEEBc8MIY88qTOaOyy9w6cd9W2f6+eHa0Ds0hsDIcYEFHVAc
VmoFaf4g7iG3WIwP8QKXnFhZtDlyDiW6UDOBSmqGhZZVPXrEtShAeGXnIf7wituXUI+jcutU96DO
yaJa2Lf++JTbrf8ZH1k+1VK88+mV8FHF5+A43c+hba0L0R7L3BbDaejKfo7ux0KROi894hVm3GIF
arcVqjW5M1s7nYZLQ8tmDQwY1ArjDuL5v2Q/Xr4mr61NYupzVnP+czMekwUUcrm5P56dtgcnnto6
TCuQkL+JKlLNbmYroVr8IUU+NiRo5QsucnPCFNCCoxfBwBD+fi8s8wSPfGjxWVPXExfdBJjBu4BL
1K0Mrlo+7ru+1WI1AeF7UKBZr5rM+Bhd0HCNwQOF0P0v/pwArNkSWAio083x1US7Uj1j4NkuWlI7
/9eZSHPXGM+4i3H/kZV2IHhb/+QH4kGx2PYdsbBB8yYATj/YwOG97lhHyZees0OdYH0EXr97ozzk
FEfYjC8yK2uVMUSiPpoBMop77QScddSk6/x/R8jGteNYu4rQh98ErIu0x+7IAPU2CO8hzafgV19I
/eks9bwysQhclmp74qXPsedch9nUIXRbN3Wfkj7Mna6HMEyX8Ng0kZ/5yO4Xc0r1vKuIg5ceLgG7
4W8HiScGsTnA6FyZ+1S4IwvUwuDIi/TRvYa98AgJy5uMVq9Z4b8ohaq3wAzK9VMndZTWJh2AzEfr
ipgNNsQKCMUjSt4m//WQY7VQOS34ih3bUUxEVPYb/RCFxw8lSDhw2iLPA4t0rK7hATL4IPYKCAbu
bChM/xSzeZIbPsDP7Oc64a5j8OaiF12qRtUMRa1Fikbyvh7+nTL8GQecJe68HIs2W4l+AB+1uZI9
o26/EZkK0k2Qz+fGKLAlY1b8Q8Bs5Ovrmn/OdBph0Wd3hruxMuNquoCyFR30NUq0Z1uzt2DgyQO6
hMrD7wUnivLGn5WprJ16DAmHX+9ERX7/aHo4K7N2g/yn8eha0CXxFECkxYxCrvQwCrV2NWWm2Qyb
qWlNB+DK6ARi10d2Z8smawq806l9JBMcSpXrdXTs12nTAUJL9x/GEEUxcwwfXwQ7XbNpMIerD0bo
SzZjddymVa2S1WOvLgK++rFX0XyivD1Ama8vrFO5s/smL2AdKXlTiMvNdaipZ2ZBQJ77n47FgqGH
S9HZlof1e8/46/Nc5qCJwbYVWjoHb/Lr5zaHN/2NUYIjIWy7yXHRjO62l7mHQth4JsIGsqo0smSP
5fKItqnMcyOVtqAFMpgpZ0oVmYPw0hFOCg38O7qiaRW7tv88gyAbrbLQAhw/tKmt1IBwFryZjdEH
2yqEkv7ZULVdQv6vquRvt7PtkBT22XydvSW05wzUhvHPh4Posn4ptZEnu8Mqr8zDuFQwSlQ7uLic
JJ2PnXN3Qyoj/3BD77s5o8/6I9KnuMDOQKnarbkex2xGZ0Z1F7iAjduqX0GSDkNmrYBkLqIDZtEz
Ll0UrAyj4usIzcjnc8FmAPnvvqXjpJelRb7Myrs/lKStBIZms7iKk15h58r6PEas9SjfIEWxuE1y
s4RD3hNl9xB0bdXyYK6YhCzhTqy1cbcywyi3lkPPoPRS6ITW05tC8C30BZv1vfwUbK1dRh19pR8U
hY7jKORlr0KkXo0j65rgU12IAHZAzAVX9DtQgnDfnRG+ueckiQ8kN52ctQVtRUae0eIo1OeVGFFk
S7aBQbJskLsRJ5TPCXNQs+mZ70oXE6w55Dmlq2xQHIqku4i48WhNJH7N4cUQ68BoCfY8U8yGxcAv
lT6ZvQgG6ott5mevTsdZtJYFHSh6TyNX3y7uO3D3zgv8WgRORFJCNYvRkGdKZwpqwaE0y8bufHTy
Toyt1MBMM2ovXlS41WqnaON6lLv1QzjEzmvNuZJJSAPvtzvi0RsZ1Eb2Ty5ut+3LXZBGOMAdfkWh
BzxCme/aVL/WtAS8ksq6r+z3ItCD3GH2fDSMte/qapsRDv9S41y+Wf2FBdshjsShvbcBtV/MoR4+
ysMqevI1uRtP3tgXKzsBBJfokNvX5tsJugZ/+Gt6LfNvc2LCnZeD5VihMPzVTqTHY7H+K0E8ArP1
GpDdT1fwThwxm2YfkaAf3cdFT9LHh0e/u3oyoEBDIlgxjzAHmGXJ6ktLupY4EqNXoZzkL5G5McZJ
grha4O19ngh8zl4lxJqq8WYbqntqnFHwg8QtiK2yvTP+aHlx1LzuFlbjvQs4G+DIZchOQt1hCsuT
W4wp0hzqY1+VD6dReItR8cp45BXWCz2GZcMJKPOMKTvZHQJ9L99aVRJtg35FluVnTkHzJPYBsmtS
WKPu57vFCGVG8maHwKPKFCxrJD22CaqWacPXs0zhOCnsIHwagztDX+adJXSMhTG9vKhFqTkORXek
7resNXJ8Q+5oYNi/a6hGiDp3fFpqYyaJu09x8wiz3OwXBzn9mNpgOAJ/QrJ07W4qEsKDJn6sVCa5
3xD5B5294c4Pxz2//LYYzEOPHSaTaHij7uWtqygOH3dvcmXwFC70uGQa8d3Xyy7Sj74X2SpCLt5c
OPwVG5YIRKc3dNhloSFAsfxhB1AV1fFfrmV03O/6qfKkx+NaIQp0ren0m19GT4/mjNTzW0L22HN2
Xag9Vh8/TSkDCdMZBB44C/37MOEEREdqi3vyFNqWJs23ud2uO0yx6tbTaE08Spw4EmtAgArMEN4C
4OUtKynRFiwBFNl32YN1/Hk/uIRyusKQir3A69F0NXzxu6iHAcSEmq5km5ma45ePv94WJbTYu2q2
Ftt3tptKEZBLwVOYUBVFPxlw7viWYmmkvfAsDX3ve8anl0RIFOISLoLYwIhKTJtkTM+Mft52cumc
Hn/fmcCFxEBj2FmoUz/aF+AMF7PDJW+fIiBLyANxa7MLiw1K6CD7lljzaXRDZ4DfNDIPbxyOA6TC
tJziuADhgD4Ed87qnE6N64tWIJ0pFZwjweEpK/44wAtKZPVJJyg4H0alO7Rz2pkAKSik4z/1qplW
Og5zE2+E2YKPhhczmIVteWC8ggfzvsyzd76KIMtMNh2E1wrRb8Ot9cv02tG3dUOsgV3oKEAF8cB0
3aJC4A+9p60EwsWEbUOjer8sxhy/8o/oLP0uHX+MLqjQEDNs3WluaYjfeapaEORN9YHIkrfytzkf
dYUZ0b+ybRUV5TzNqVzdC25RYiNEKjazENm+IlMIEsjJOsIOg1GYbMbaa5WjmWldbG+vzDKTsDjV
fv1j2hFa+z9TZePTLvm09jG3UWUdXSFwBzBQTLSnQda61TYVPdUwoFPMtrsLolTktVrGJ1OWh4KI
+HYZe8IZia+KG+OiYSdIiNsbRolBDq8WtNe81QoF1b377Yzz3/pr6a0aUtg2aHVoLkfdpcDQQNLI
HOS5x6i8UgOWMFzYmxC4c6yGPzPVqqzWlioWOrVEeoqOmG08+ekgjN41eELs/fgaHeogpBs/WD8H
sZJiKE8Hhx5CsgvneAD88S1dFqleRZgJFUkkZCMLzjNcorZF7zUrnH47nOfmQMU6G5mQXxRE2G6g
Wco3nkA/QVPeZVMfE84Lpw+IPW08U9Swk9VgMcAQ7H+OTMO3Un3/ANIhizcZVAszbr4MUSbg33ML
ZTpA8yUCOvrd0c9JKYpgibE4jWmlWbWtKb8Ll+U2JddeX6PNh5cmNNi5MazOZPv/PaXSJQeIelqS
7srOyyOUxSEi/EvdsVLzPR1Xo4SC7+B9XOjgeIgy0iutr3HzfT4/tSGNa8I/G2wQeZDB6jej4T0z
ytS/Q9ruJz6C49rcLzcXo+pj0/HIU5aVTAmqxqJxA54WzHaFe+OS31i9hW5Psedaf50mu9FJRp3/
lLEjSzYHD/Acv3RJcVPnjN21Ya3Hwln/sW6kxO8mGO4AQsCZJvogyjUMkw0zFBMioiZsXRLcJx9j
rARV++UPwamqAxaTknW12+er+cqnGJ/zJM9TxpsZVMwF5dHnMBqrNESJmB/oOVDDENRYt4KYhLxD
lv3+OcxXwBmhLUfcZXjWjgV+L5zo4+X0USR9wQASylhnj9odpBwTZ+tYAQTZFacvcE1oR1GBJxSK
KG3oJozBdZC7QPhcPOP3xEkbEGP7g8bgzADkTsdb3ItI0F/KzY/hoFhcsgdKd1RoPsbHOYQgVe+H
uopzSf6Iw2MGVjiOJCkwbWZTSuv9D5dlM9gDEldgYSKbNXPoPgKoUJt1XFxUUG4nJQNF5aP56QJn
6KmFMlz64NPECli0I5DInIr4BzZnOL0gWxMvwcS5PqmihQ/50Ep6Fxkf1rstbrBImLUklAq70j8+
LtVn6AkDS57frzIxpPswYGJC3aEC27PvZ6KM90vvCsqsvbcO6DmsFAZyxe+DC/U6d3aggAUD498v
OxVlV+OJmRvaQVsZvPfUaftwNmVisZEoQO8kPekb5iGqYRJxydNH1kdrkmMXn+8hAp5eqHdUtBTy
jF1aexbW3uX5BgmZiCWoSywqp9hnHV18N7ZMcnEMx+yVkFzQcsiSAlJEg0f1hWRoEKhydMptdOEv
bJXiSUk5TayoqeOIkAGBuls8MrGpo3f+bwFKwIy63QqJUj7R/wtt72cemhXizf31ecCCPoWDp73N
krNZTuyggw1khJVnODLjmmOS4P89/smc2EDHV4v/f/wHab6jrV5x5bQmTaC0918lcUEks1SmITDG
j7eb0NYTlE/o+X6ICZCr5GYFLoAd/OM+Lmw9aA+q0UDyeeWz2GV+WZEnqmNmB6iTttbSMwhMUjUo
F702WPx4mJcr1g2LNPO3alBcMKL7OzKcB/53uJwSxmtFvo34K7WEFjcd0jhMLLL6A1jx38mpa6LK
SEp5NsXHki5qQNgbVo/1QH2dO1GZFAzIWaigWvTiSWhgOxIyJpBFpZX3lw0Vwv/OaA6ZRLsp5kN+
hIE6QX1b5ywds62eGNB0wjfqjGyjtV7jd+irGauwV+t4yf4WDGTJrgziAuevzojMo98Vo4GVmv9J
/BU4BVCGsJB+aUsdAzi+tkPY87GpH58fW5PMwW5mHZ6ymxOpmcQBbL/EESSHXmJSC4voHPEjINfc
scAwdHvEPyXa55vBXLix4veUxoBHKNxNwvcqdtO576Tjdgq399GkMUnnxDD01/AzTs+Xt9COuu3P
cvQeRtUYwrvWoc5asCSjKwur4u4Ugk6r2bYaquY8DV2Xrh4E/Z8vubSOX3hh4KMxyAdjxn2IM/97
oIQe6f3aGG1U0rhX0eyXCTUg/LAFe31crAnVHzGKfrItbYzZOoWPix38+C+onvJx1AUkBdznB8ig
oXtkdJKJydlPa2/Aq+tfrtBCW1byVcb0aGr3tocdtzvLSAyk+f3An/RuKTJg1XkccWVsyIZAlWBF
RXTx/ZbnQgLotgMWuS77IO5NutAoQtlJDLyL8LSgak0GP1uitvlkeAW+Jpqrg5dvVjXC0S8x23Pk
XFXpHx2dq5C3gfYcUKmU98h8BG8MFMoG8U79RFxZ13Vph+KyxZrNcx+/Q3UhsoHEDlAc+4YOXHXf
OrQ26T+R4Dxt80Kw4XDB1IOQZtHZMYfrlN6/Mj0J1VD0n4I87q7RY7G8zgiMaGoCcdy7qs4auMT+
9ANYkzifp+9u3GTH+zdlGpxjXZxapcJFs12xtcOKpHYpAq0oaPueBSd4LMUNRvTzVCpOPFvNYevb
Q1KEdK4wDdcpmC54IgR/V1sIZr+gJTl1Rl/B0/p+aR3S8/dElAZEQuwrm4wTsWCqCzWz8re8Dee4
o+QzIPWMfFlg67gvhHQ4MogmJo1vTX1YWygih8/0zjylXC/HgMKXvmRChLq7j4gh5xVeinALLs+E
LkdntxZMc1Si9nl0fmAA2paCKchboOnKSOwvaX6J7wdbX8kCbYj1w7be4KAcQyUHHtDYMbat/8av
9uboq7NVkeTxur9aOGs4Dy8reFfH2osmE1uiaXmYHuju9qsL+mJGIxuLz2rYrHBByroyJCxI3qg8
Sm2ZIMTxzrFNB0GWzY0nTCCZ5rysO9d36yiKpq9lyEJisIArmpxfdQ545V1UYvlYoq/P6vqCvzgr
7Jm3aGPdKVZCzPOWFz4Hyud2dbIle2/dAoAlXpOnfpwi2EEuqp6sk4eRjZjsNij7lKb5VohEvGw6
CBOAvd9AfknoS5s1l9fRwZt7/8Xz+DyMb+GYgri6VsfqB5jE8AljiTOB1XAYOS91h0LnYgtiVlK8
A/SAG8CAFDuhHn2YjJAVNT7KWmOlmJHurfuMdQuqK/i3oddioLuCaM0YUORAb6mZGKZ9c/7b68Pj
j1J9NgT8OvIqL9/fNiQh2NztyifdeUnBneHAhtAmbvXmQYc9Vibsgoz/ai0wJOrt3rwh/BauagYj
DT4/nHpIPJXYxa9lMhyqmstTkCwJEO0ncM3g7SKwy+eoWr6XWEqWPE8dq5unhfBbtmNEA258tjoe
XoV8BLvr3OrPgtX07POlRu9wIQuqaquMdW4BEZfj3y5r2+eotrrLmH1ONhB2PJPQjgc6GIWUhha0
DEzk8cPuei8BRf8xWEQm5AVyznc4lUJcCm0M5nMpp3K74BCiRYF6pu0KqijO77L48YyhOU9rendp
Oqu40DvA+lbjTL5oM0fh0rvPYqcKxCxcw1QRUaGuQPiO3sHeUJGiKgUOtQqCAz8H225cFMCgOtL1
xXVuRlAqhcPcqs/j6U2+e6Fbemy3XAf/byTNRJpneffR7fPRO1k4KkZGZLknR+HjAbzfB0S4imwk
HsU+k/Ah9FePaDRrlxMtdv/h1bXuYipeVUaRCtEgcaPmRQWlAiGZbV6kTccbelkTSFomNqXYCQA3
uK0sSTJ3DvXVtrQrnpzAWtDCGW5EXC70r51FSSOwVClXXqI/Uo+aCenXx3G748ilOrEUMfPoVqTH
tsJkwJzxslOtiSEXQWxQgpAfX/COVfY+QdMp/yYiczTM+RDYeyLSWMTUlhrsJ55FCJ7ZX1fe/Xmu
a7j4xXeGc5ivKA48fCptZz9p21ghVmmBwuWSdzskOczfeD/fCz1CaR1tVkQ/si44xqj0YyazCy/q
3Jdwbcq7SnnrGSg4RHrVMDQMt4hA5eWJbzlIZKCaSZYPLQIeWkB01QjCHxP36qVVMGh52a/UTSsx
9AdfPruh4QTxVz2Mdg90hQUXd/HSFZZHe/a7G2TuLRLLxhNB7+x7fDZnEXdzimA8syLZ/MDdLnCr
W/7NP5IMdQ2F/U+81dXpnXzo7piw555RfiA7vsDshSgRuYRJcMLgx49560aVShPpusTYr6/6dIkD
actEhV98qc7b68XdwHT4jhlzw7+hODQ4FDKe7G4dKgIXPaZL1n+hwaVGFCVk4X13thTIvkf8UF29
IXeLro9GtcdU2eEwDGfkyAWUCSVFk/CoGCSTmTvF9Jb7wbJTkeJaMRTzQ80iJGzjPiJQ46t8D92d
RiH7SlXoR3NqUw+Duv+GN70lzwDf7aOXUHTwSRwm1HXxHKNnSjph+f2lVfxlXyXvRU2zo/1mkz9t
eHgxE87Ufm8uMWPaRALpr47ll5DGjmIQCKFph5zcvCRXdhRPTgLAShhbqfK4fJyAz2MGjBMLn5oD
c028Z/48kt6Wd3TSsYpfV2whyrh2r2sq1yx423zQsoVsF0OOsBOIupFMqfT0f6qDfe+Y8PUoxqAh
XUmJb0+x65kxnBAFeVhBB2bc0JeYlLkqJ3f9Zgc7FA1acVezDrZhp1XMRyDB4GPW+eI+BlDv70CE
72P5tQwNq82Pb82VyAOoyqRPYP20de6oLY1s9lR14nb9UHF9aTiNymo+1clKYH4HiKoWJi7fICzo
7ByfkS4d5HXijM9ow9M+USsbAsBDhCoycndhf35cabqAJYWqwKqIu+UfHUeZQFYAT4YhSoL3Z3Dd
bYJdNr9j2i0VB5nqaNidEQ4sh+cKmPIm8iQAPdVADhdoPucT2RwAGr8+QC+5BREpVdCyHId98ivT
1K7Wdv1GoTb4fCgfcPGf1Z7viOdHmLLKJo5wD/znZeUuA1eRs/QlMTId0xnOp13AUS+LDK8YYV13
i8TVnXhan++t6IlXwS4d3r7kYZ0+GOgZcEuPjwB4jm2+KcjnOOBi8V87k7DREPuGv9Gu39ssE0mn
EkdJCg6mcHaJzWwlT3lNqBXteHFEovF6A1lUvex+LHNvmp4Yl7D+8G3uT/ZvNg7btXrThuGi8bj2
dJuB6jvI/mlprpw2X6bEQgitTZDbD40mkn3rSu5e8/tz+LGiE/jo5A3pfMHF47j3Pk7IQdCah2Cu
deIucfL+HTwv95W8VaK7/dWnpRG7mWTJKgUPUv660JbjQ2O3j9FH/tZ0hrYxc7ire970uJH202Rx
yEMX0Ypw+oKmEECmck+XcRp4wVTPOsE8Dri7Sstylb/ROQ8mgHiu2eaKU6YMNw9uD63rGChb3rJQ
fkD0sBzJhsSaH7R1SZNTIGYHGwWepNPO/TxjX4Ci0gwqJIQYC31NWAKZgoqjuFoEKmrIk0rMmv7P
2c6V7Lf3NmK2GY27A7o5iIJylHheinGWpeJhrN28In8MVTV96s8XzSoAlVyNdlGh1UClvWn7+vuM
7jfN9oMN0UqkNiLzkzaSYnH3KsGlcj/FYNomQ1x6aCRfMPqRE8+fx8wvZdqjaWtUbP26xFNcBvdH
JH8cs2Qw8tvM2IvnTPnk/RORHIqRulkcZO+9KqWQiRDF75A+NZy6KSCY8eICe6JcmK1g1Un/sl/G
B/gscrILdr8a29DUIGgDOd4Y1N7/E7Q7nLzZ+A3gosGFLkJvDkQCc2tltLmO+RFX3pLQK0ny038Q
JUIvJbFhPrLFsqjkVlst1BZQPMlO8FoWO0pWerDL/uyIbVrMHaMKvoFyxqur9azowX1B0EpQURyd
iNfkoLSG2hjhGbnwzBUxk38nXoxH1+FOXO+FGDRzWbntGmwSUe+xQWtSK5oid8UMduvtQJ0iRvWR
r3l2/Fs4g+Zmzkd51IyVCcy67x41PbqEIOmFIERC7961IBXd714vcKXRYE9w7u/GjNEdxF/XLiut
Up7kjBH4KpN6q9Xggu4g9cA6WnDm95pAg8/CyCv1sKPw2TxWuQbfdVfu2v7qBVVtLnAm4Or6r62f
91h55i5jde1bMej5MFOONLmXGuAXZEsDqXdggxEL5oCykuYZo86bQWdmNILjIEYkzF3aWh+RlqE1
q7AgRSwEKifAbbo1OS8Y419aJaNmsuu2CjYIN+ppBaGD4CL5uOSe00yC/HH3XOToNfrjgcI7oPu6
uzbbxwwqUwd+uShmJJI0yTBBwrhUhvDKdyXbjXpCE1ByIqtr6zMFQxCQBcvh7xrkEusbu2+9zjMP
PMG3+0nFJJmV6uxBartmaZqONSoOTlf8BHuHcI4g3ZQzNRpiG/Sj1s2jRbPhC6kuommJU8AqbI9y
GwWreM181VqzwO/arJUJF4CAXrKMl42aPWpS98l91F5WDHvgWfPEYX+Az0cGZIkUBhkOmVw1EA8M
eoFjZd7xr+CW01iAbS7lwyidua4DhEUMPQWYiPws476aF55TKDFKvnZ9Z0wBxbvhoSFWdJWa+EVe
yJmjLY6FblY+ec+9hJ09vEIBkoasy9k4y3pvEv/YV097mngZ9WUcqQ9WDlOmT5Ku7c0dDz6La9BY
gm00wGXcpi+T94J9qSYDepZNC8Wb0X4QazWSrLQlhE1omoa5Rkp6g+xNHDWHJOaEUBsPmN9hxrp2
AYTiClhI/6GUFdSP7UEQTWzIfZt03OcBehCP8NcJ5u9KKJ/hLAqmzjItepRLLDfYfBJvDtrmTa29
YdreWEvbe4zJleu8vQ4cPKu9IFzoAWm4e7UEv90IKQcrl1+xxf0nhTJmI9btB7Ueu7FnaprOpj+x
bqlzMlkISE9ptpjHqRID8sR7cZlKKLk+2oC47R5J1Gz+qi6VQRrxZnaHg81orJ708xjsWoSKuO4H
YQHiiKcrGsON4FWfFoKqTix79qCrtrN5oRxakz7Yt6aVY/EXB88mmovYzAzZzxZv7KFpPiwnS7NV
96ptHByxvdbdvGiy3bEPBl7u+7UJxRBvdC+r0XJO7FJpliMg1foYUX0lTsjInPxOHHQ69+wLb4UV
44wmA4PFc29mWs5duTnxNjrVS4egmGKjlebiROVWl7ZoCgEuENMbaYFy76Na9s130haMO9hoAW2x
1gXHcycyR6DKpluLgpFZUex8kNJL6smA/KRWZe979Em1UwwhIeW0RxXNrwcQzCLoHchTBJipyKX8
TNd0ONqSN8qsxMch8lBU4JNOjFegudUav5HplbimMlhOd8R0svXvOBjMGudrRVQBfDT+QAjyI9no
dz0VpBwGJ8ZGXw9P5M4nEiEQUNVKhPm0bCnt+dNM3hI9khmLux5U3/oIkpuQgXQoZnhpE1z46qQU
jo2XT4cFAxUk5SKo9mQA0cPMiVPMm634atuygh1pOafZS+HWLi97oC5VoRG1O8lQ50YJliTSruDl
yvpDz4JKwd6oRGilhfyoPKVA0ys25OiVua5MiAo10WgjM8K74XCvyIEq/DjTFZ46ZCNojRDgPt++
vcOCxUstzmmxK3j6WER0XTjjYUjLaZ26A2hnsVCLgZvPI90S/etoAUrOCbJe+WofY+VaTlmhmlhg
6LHfdkgMO0eWyOgMn3N8YLlHlPXuiL/TnIgtngt+oA+W44Ucl5dQFqgFJeTPVt7zRviBj3qJIVu0
Akhr/WQKJJv8LHaG5E/wbyDWXDk3hQyen3K029QC1dOW/V+6eI3vpqqw/6h71lut3cZS3NPog5N+
U0VnehHqqnFKnznBJqBNtWasQHA7ndQ5hgnfST0q8JlvL6QNaM1kU3ZcThmoiI0x6Fs/5PqrK+xx
nfUf83DOme4vZ9nDSr5ViOWoDLZgev47CTjIfY0Z278DuiH//dPOAyECnTa/YyWLFGu5kRh+09FG
S0mof7Swa3XNzpZrzOyKdy6JLNHIUFljXThbj/mEYjKgRclgeYT5Yhs5Palau6vKs14ir2jaZBne
5CHNN6idbecqHHp4VobhVyZpMqSFevyV278Cf0UghyC5nCRLaC+QW5qj2fUTwhOxkNUPMmWGvkoU
f+y/mPAkahlYsQRBz0KV7V0TSxJh7LGrxG3lam77NdQ4OdcO1AukbFYGeF/AkBS35HZhpZyMx5JX
S0blqi4R8PStKatyLHQkKyQ4HWibJNgEez45x6TiPambqfws4w6tehtpo2Xe6uETBxxSPe/r0gx0
r2UZgjOujfrcAX2cg7N5h5ekY3sNaWsku14RYp7DuJuOnuuzAQix8+/9rPX4cEwebRNlKUtBUyCN
kkuc2H8eE8GiSD2gmFMoUFVjf5gy+FUugi4/045SdQ2Q+vsETjI/zM5Hfsq2cQIJbGmrjrs7B6dk
lt+vU5s/PuXBgETRYpvcqV35zFZvm8/eryGPZMvOAyRaW/nBANdoaboZiW0goUmRGPDysMrNaPD9
edxjf+wJ/UHxPCEj6muQT0koWn9cdcna1loWYKJdYe9vplH16bDkHjr5KpbWIIoDnx3QSBLQer/e
mI4d+TRxichkB66LxlU2qVOV7CX2/HwOmWfNYZ9rGlD0zGwC9+H+ajUVcN0rj+SKXi6CZFoRH6Nf
tVtl/zoYmmy/+T12p2MLhMS14PRrcq+DXTVKp+Q9ZLWnRPvMJGjXMx9iDvqZn2o3peeEsohnYofw
X1mFhe2zHlijyonmyMUkzIzPC/yRDPHD+kJTtpOinsq3WNzsmYGE7DrKs14c7MU2gcIqUyck4Xby
zVWqOWIabLfgwF6Ab/GoQni0tJe/uzy3x53bj0O+Nym4+4i/hXpfrx0+DwlO4JDhAeFNgaU7H8Xs
ds80u3q4HW7/BX4wVgpeclTcMmBpzcD2IEHqhj82CyChgK8CBfbhJMh5Zlv6pr91a5Abcqh245LI
yeefAODl4QyPfTlDltfifBFtzdYdB9cdAInyf9F2rEAg3P+c5zP+0rysTZPOyH8mqUDmZSSv3q8V
NNAsul+C8uP27HUci52tUvbXous2G2Z7CaM9J2sxbt1yrt6YdlAxMvpuCo3VaTSU4OBCJqhWVBgo
hQYg1HIRPaIqEUQt4Mh6eiR3XVYDTdcmjpU3uEELJAmra7y+vWaB6OsHOrTa7rOkH0G9I6h71kbK
aQUTe98SH1u5YhBCXBZoST/a5Im6KZKUXw3pKRAtF9rNp4smnyRSCZ9KSOX3JRPqq6kaH5vlsPCZ
YT8CaF5fyw3WE+kL/rT9yEUj/CYCxkFERX8Zgte/IdBuLfPsnm/jbBNZkmQ4tVx+VuChb73bhYNy
zwrEGFuevxlnUQmVEbmpw8+TguGiZ/1lHP8g6H6DDWJ2a4p6aJ82QOYyNNYYOZTbRhSSYx4ttvAl
uK4Sy2DdsFkR9v6wKwlQdXq+35OfgKuoq+uoofPd1nQQEiA4xh7KshgYwy1Fi8m2x8+5JLqwpzz9
cDfLDWoojrbvVvrEy3FivJa9MyJEAm/HzyxeYl5tg6R6aNm6x36TqIZ6WnyJ4ckMh0+yIMnoS2sH
957kkJCvzPPe2zRSKVreSwjmclUn853Lm0hN+osECOFtqGkXBsoiSTZddM2lkPPYOlTdlLII3buo
ZEIch3WD3qmbIJER2dgC+uy3n59mYUDkXEIB1zjV1nTKuIUucdLR5Xa9ti2wXCeBhJxzvebxaby3
YhlK+ZHQeGi09g2QcUe7ySWTVgQgnsrLbWmxvOfLdawoZU91RwG0awzo5JxbKXISVoYY5JtT4LlI
ZzuszeddE1wGPHWXDMeyGFSefGUPT+Gv3+D/33AkYGjXuFm1AtM8TXbba97z3b3xo3kED764yGbk
46YBhrqq6q2EQNbdqulWDsHnn6ff79FUia0fTyO7ds7hlGRAAkFdGa/JyDcQSRWnh2MGy3tyTTby
anUzVgpgCHihra8iS2VCo1P34/wC5TcKLxW262cp1Eg3a9zmqnuF4vHcMJmqXVDvB9X/mOxkmbA5
J5MZLVJriFc7wf24ikMbtkKbIKnuoILWWkuOD0ItuX8/DQ+JKuRdYiUTrbeb0X3jHKhyn9mtwhD/
kI389Cu/GTgy1OkLyqvM6oM08qYWvPHnO1ertOjyBlMVgOHsqEEgmEMOP7ceuVdFn3yoAk7HECfJ
Mky+XwX3isPve+8Hlvz5ip1UarkU1KAXuO/ouGcoG/BGhQVmeg0+Wo+YuLNE1OeCelVlZFh/Kyov
Z2YAy/YBRLhQTv48d7ayukpGBQCp9Dz3pK2lmS4+tM7wkYInCK0VdehRiXZx1MJS2EkxFe5gmz/V
iQKP/6jOzj6mldDPfjxzeiyo9kvd16pm4VE2jKga9n7JfmB+2kR/XlAMospuMyLB7GOlYupx9AK/
xaeEOJMkXyk1K3aI7bFWk7bfom2ToMFn4xPynX5XnZYrEhsenFdi8kov/nrL7wij0RXi6SR4+QKE
/0QYJGA2HIe0dSULhwpZJL0J69jLRmuYLuzMN8ehrV94lVxinRhCaqO79XNuoU+nVPyb64igFNEn
mNNloIw229mhhnK2odU7PqkNaaSTceZ8a899OYHUVVZq+WjTotzO9HDJVG+gRcdna50HAiY0Z8w8
11xY8sJjVRGTgV/SUme1ponPZDJSWHpQa2FR4q2K7fFP8hAxEZVse1MZ+QJJ+/qmquKhYOJYHVZi
wsLf8kGtHj03Uy0CxuwR7xVO3VyijloYmxY7oegjk5X9tsedi+Ad0FkjETaII45B/KSQQqlrQr0V
Qr3r3IahJ52l9BJsd73wXYhiffqNgm8xRbmnZ4+1iORqic2lKp6KuSejXiew1mhi/T4TW4/9K2nY
nqUjKwdV+c82MNcmY4vPrBMq4BDf/Moi0FLY7N9KzkjJ5YAn91RaSeDWxJABEg6n2fWrQpA3WISs
Lno3lRnZhj3bh8e3dUWDFt8ng+M5U93jS4GAQ9irV5w9BFWE0+ccBYC48eEvcjaUqltWFfkuzoJy
O6ZNrUZLpqhakzmW8bzpZ+xBecNSso2ceVL9Ueh5vFRhXDtplPtHME3xjsbFSmvyi/lV4lqNqAE9
RlLYh4BIrgrfiIwgXwXZTkcrZlLGihQhJoR+MET6+WroOclCSjHirptJrqYL3V2q+YxoQrsAQLqQ
MtEwpo7/wBNyR+Q/DqBQiz3JqUaLIrV7vPIUfLmWoNT9f18t66Hcodyj9GrzQV3QET0u086aadX2
Ugw4hMwjMeGX7kSvEfmxYT7JeQhzo6HxSnaIkDMeCK7uPQhXsI+Mw1xTZEWiFMKWAcn7nExZBO7X
hQyk2Imzky/YIyzfrnBRK2AWJtnchESkjDKnK87KInZmDNi7/qJ9P7zW3UiWF70DjVULbJAz3jv+
5sLnYUSnM9YA+OO0EoN+0WESe9nodv80ijiLv8AC0iewcQaHNaOnCmnw1mDxSsUytYhOc7SjnIFj
UXmU0OG4VLoU2ueeFgq7UNf11+I0K70hkpBw2QetRSyuw1NYBDrJN2Zijb3m/g3f2IrPp8xvdbj4
F4S7MWbcJX0erQ5fF8EQUtEzgmfRoSzUrDGjO+4X/nEF7ooOkEUY25Dz8YxKXT6trbC68DJdNZvs
FWsxqUl8KhiVLLnyOrv44ystRGfuH58kWY1CdPBJhJuKkZmpRnIIuWHQzZc2y21UP5M7Un0Dy8kF
qNDV0YbPjHaFvSNa9DkiXIvFnR6PRIz269HwctAgMjIJBIlnKvF/+myjfIRCRDPI/UlWAcPgo1Cj
HR/F+WWOmf0I6UlwXOYgH2wKpYTpU8kdj2tuTGZKDVcZguMdZGgVdm8UBLb4q6FNcQZRxw63eyX+
bt2psuUHom5/XyDIE/BbDzaecrjP5Q+7vIPlZ2wZadjViw4NJqGEKsIKUDq0UaGhq1kEYsAYYcm6
zjfomSuJvVMw+8e5Xl97ElBGGkiBBM0vJsEUI4v9xqhtse2H0CWRvcKFWyj85BY5CkDlQOl4wPN+
Bh3I3lG+BkaA44dZKAh6kSG84AJ+xbcc51tLVWecgM9vX0CsqNVeF76bWMj3X4FC2UNlgjRUPrvA
IAE6CgCrQ685ppaS48DMbky67Xp9X5IBoeLN7iBM9DNZRa2ANQBOUfAcsraxFmiSJUfByImrqTvd
gXbbXAVxvh7jNH4O2b+eqjO1y0LdIuXEU8HoDKMe7TToKMsKSrxgq+prmzyy/7LGK8ClIlKvTSGF
k5/i4SHlmQBaFssDG21iKitn3AIJhN9kagPcziddBDcjuK24IjRpNmEazYB9ok29FzgUVk3Co+Ei
Z0BB6HtF43+FM/lr0kPtCaIllBzBB8gsz/sya6yCiz4Y9V3UQnEEoEt3dBOwF8Oa5907+ycT0seY
2kiTPuhiV4fnACUN9TSlhEBbVSnDCqTkFB2orH9GBYFAz6hQb9CKK5zdCGy7fuRvz4mlGbkLvEcn
8/rjw5DN91Tn/bqsbTG2uU13UXHzHvLaDyoJ9aHc/Rp+mw3ijx7DPCotWsPVzkQh93PJ3MSZrPU7
VysUEQtuMUjliKKBORsfGrZcktilBqhQP642DyhcS8+vuP4UarUUtnstD4516EM9gtlFuGefzyhu
cYNtZ3osLmTmvPVGRB5JByoTEGmXTJ2ixoSTzud1VeD7bB1AZosXzP+/5cJHvLJyDsFoXqw3xG8/
lH1icCB3kupRIe1CGEbQGavXIdEO+9EzK4z9rTfy+v7AQyiWCIrzJpR0CjQyH7PFTFSN8qDiIsoM
AxvAFbGPXF5M4EgrJ0yLWLCuGj1leL5ZB6It/rvhf8Bw52Ol002ohaLopD8ESp+wXuv4G4Fr/hR3
wwlaETImJtWB1mFEOuLgmREPardElgEUmxWrP9saBUz6XU8eiBTqeXfh2O7MgQu7Uf+sEjwJb/aq
wMF4yon/a3bsoCCRxAhYV9cCLGp4Jf6axUKcAoIBfZmCHRAcvXZ/YIRrlFgAMiBrL/pjf1RU072A
wfLCEcbBfxT3bxdo1Mn2yJagXpdvJkOxRGb9iLXoOZm+yRrV20Sx6J1HPguAk6gxbvZOQ8v6PfoS
xKtuNXeSp6FltpJ2ZiAsVXT6TOEyns6s+MNA+Wc8QwPjPLAv/+Wt5bIXbrXkXxPgIyRekpj8aiHi
+5kteIxIm4xmszt75vTr+Go5UduphNROQC7LoThRtZHMrtPiXhmwd6ht9l/ij9Vh939arkAMffw1
e760T1RAm16TzrC9765HtzlWrX2EY3jJ12kJP/OPHBJpqWdEL7X1DET31mZG5kEX4M/n71VQrugc
1umAbdNw0WPEYw0COZux3X8zNkSFbG/fxfEgthTLKzhnWJurlJfzLSFVH5RUQeQnyWZna/SgevmI
QKTucVX9OqkKdgMtSBoNUaxg38Nku6GN/kXKMD3plwZLWSgT50Jl/ztCd08Tz2/ANHipdF0qhMcg
SqTI/+XmqsJcwHWm24g1QUNm+b8jdYwF3/mSwp41Lb2djz4ZfrGU1kjUIdzER588s4UxlAdg3cV6
pj9pR2qZVvGW4UV+0p0RyAcqfNRfSBfvc0GVOX66n/2+0k/HBgNsTqzB/wRqoYAytIyKW3wxMxeR
o7qRAP2vvdt3HKZ2rrbU3qtLXjVfyBRfDNmqjccLXsA+xY0B9GpBXDs8qgGsqNygy+hJaBLCAudh
7uYNjwkmxHPvR/8FWqP/bB2wJQa1UuJPb7wIyVP4fBMNIvA/9dHwJIYW2t98d4zxr0ZaAqdFW+Ud
p2LvztcCIQLiwY22/9InFbMih+BTwxJ4MLcQoywUynJzvJDyOVih7ELzdWnsJ1rRu8YQfOQ4710u
pmZnaLvTsq3cMGEb8AoeWhcm3ltJfhr7wiZyDJejKGbyitl7DNw4DVkVPyCmwvc+5NlpFCRmG9Ha
he53xk4dX0d6v0ftsrNdp15vOkqSR3+LRShS8FBMsLR35i/WjNO6uGNfnpUW42a3J54KjSr0cpJo
9atoDQBgTU2vcsphJ0vnIg2vV7WjHj5NPhEIcR3gvLWOXGzXU3sXdQ463PBnL+OgxpvUZ6Rw8jyQ
d7P26dRsNLlfivupj7KOzsVCCmD19lKMBUgsscvwsOWK9v1xOexQvELHoMnX6LLkjZbFSI7/PVrh
AZWR00JVAnDi/fQeOsleJBQEDcD1saeu4fAlPX6S/1vYtOIoUFGWOFtOZoU7287zgHP6XCRpt19y
bRfr7qIjDn/YK0GdvoXJHtyn8A4inBun0zL8mq+CGoGS1oH6ch3kUcVr8V4pqXqUf7chZC5cTkpH
YaBupTJ83l/LDg90eIHfw0A4ps9og3M1Wp3K0S8HqAJaEmePNtZ0c2vW6xpcASIj0j+dIrt6AhZG
BjiSXeW4kT3ylIhJDHoXqjd3N9WkFNX9reot3CA7yitKg6+GvhQNxhMNPQk8FSg9U9JSz22ob4/R
0bV7wnFonzdMCAIAAj4y5kLhTB7WP/kTaPSNvmwuqQXKpB9BF7DhcaB5v7JLCvCfskiE6BFiETc6
aBTeYK5D4zi8BfxVuvrSRlsaRcFxefPl+YKEuIYub5nF53qtKxWKPuP3VTXZPFwikRJzBufS9vLe
SwTNF2gEN2/hPKIPu7y8+OPIp4ZLBl94SNtUhWlJF0Jgh+UCTzE3xebJxx07A8d0o9b1w9Iz1FfO
hwrQFL/nR5Et0HWsle5++8RqbBQMDcDpMGD5OKUUa68ws23cYQbCDJGNYy5UYlW/EKGWfCZnyoeC
4kwLv2Lz54jtSbbqz3gHzSsuQBrOTpC7OCkL4DDOZyRy72c6k3SJEg00oP5bia9mi7cocngSQWP+
NBOy0z8K/y3T1G4RI1QbaEmXjD7GK/OahfUnNoiu6U6/cJLFABxYMFguwjKFuor4pZ6A0yDbR0Kh
BuhRZTDEJoZzLWQ+/pmRRyrbAnH2VauwgGYTYZmOH/ovaqKy9nhXVmhtv7BhwRRqK1SEvkfPG79w
33Cvs9Td7WiNiQwlOPS4+DLoHjeGAfhFop6SQV5UvY7CZYzqwIm9g6QsdQlIDjstyyOaFVbdDOQE
99G071GPN/V2DM+lvHcpaPky6EzM8neWtQaIKDw9DvuiSr6Zqca4r6ZRu1oTCGbLv0yACgSWIzOR
6q958g3XD4zAsZ8dW9pZDxIHboO1E8iD7L5+YufnzM9jRiXc5Stg+D9oWv6Ky8+vlrqDcg+4guvd
bGJB/JNeWzB/Zpuj5NAYYmJET6Vz6bhjjc5f0VeM0YH2tzAdvppzDgUr4vds/7x1WdFFKFMxGWvm
BWiWMvohx6BRz60rznDyXXXTfHFpxn06QwbnjeATavYLVoRh737jQ0O698kxrXB0mJaDfTOG5mLW
tEtb2nB/mBh2fUJLliUKwR3bM7560HrZeD+myzpnYJnuWIIMqtIsRyoz73L8WAH/wRvvXcQxnrTI
ww1T5OWmeI44wJCCVFEfQvM3ErbN+7f7OEX0XItZrqdW66N7D1cnUnsumaQGY37e7s8A6OFHasd5
DuO1rvkeBThp+xektYiryzSIk/td5kbqAB5KvjnKBq3/1HrRAJo+F2b6m5CqcBBQhM8tOnA7Zqud
NXXJX8KoFU5qTkWXvdTfwSEV7oRfkqWY3cMkEoUmQk1YcwHd/8AVJxNVQb9Df23bRg3tlMtmAcfT
2vV4DdCoVUl3iGXbsiFlCS3ygDzFw05w7kPVBcNsGzmjZajQDTuD5hgAbdsm2ISPJVX2t2iFIkR5
czAFmmB044pSQIa/QSv3pNBzOY4StzdkGCCZ3mSbFk1ZUXpMV6227HMJRyksRLfMi8JbBZso533H
PRBs5cBgKp19nH7OfmXl4KXzMZcA9J+MlAXMNAU7TRtQbYewLq9zhQt2SUNKH3XSMWh1CnHj9fZd
TzqgCm51fEazw0xaakhLiwwC8X+jGWUPdeh8Ptlc1burFTPPSjJ0s25ggnQV7OikSOJZaaIy3RT2
b6/1uDgkvZcsS52JGkTILQEhGW5L+xt9kSg/ubtKEvVqJd1xc0hh6W9pLqrGCc8DLjg3uUwdWZZw
liUDLP3ewJKhfm2+qPAiV931ATWazIPzMcWGXtMbVmx5uDHNlFuPQwWtCEDxLmD4gl96MQ5EcsLo
HpfQwYWaJYzJczc8BsVI9HLjjaS3mV5RDRdLOi90N3RCZqgeOFpEirus721Kw8Mu1hUmya+4HAO2
f/VsdmD9QdPwuZCpdnXSPMHCm4qh1w51yVL53TZDKfnVSLYnX6XPL5A0GmgAof9IPQXPiresailR
AyWZORXfV/uryI5pgEYWB1ECFKzHmQNUSNxdacG9Ce9j4iHfgzcHWqlO2GN22Rfe8BpcpfkNn2OC
qZTbkdk9SjJ9+ZsBKtvb765XSpE9bWTLAyZLen9Hn6ngrFBIoXe0YAnZWDIVsL61R9+n9AJD85/R
CsVwocQ+FYn8vnJ+BhmbtHJEFnSjk03UIVbi/ZIwgth2MRqDQaLG5iQ8fddkmneQsGO3+2M/N7Eg
V+Sxuna1ZmRALkAxBsKwOAS4CjVpOWeXro+aa51VgWjizSGgKgtiQzFFhU5VCW9+vWz86ZYlS+JQ
M5299vGVHh0ct/AkIrHfIzmu71x7V0b9fRnoIWQAwT+NoMMfPK37XsRo2Fa2/vz9ern5TiudCYfd
woy9oLAjlqnEzw+yQaSCLgfeBfdDub338mU5vDCCL66WkOKX47qYMrrnoyqpaZa1w4orEPtlRA4g
j22vhIMdr8sSZxtzr6kmzkgtLitvHHWyKeGY31KjbikFc48cPj1vtGRXUWBNDtcBXviaKPi+Z4i6
93KE3A+xuCjcpjKlvqgQPRYqCkwfjnU8/qLhKz6oYS3ikTWpPHl8CaOjjM2QDtCZfOKoktSf1Ma7
s2Ml2nlkb76TNJYicnLZX0MguRp4wfQTkTULns04dppk4+W+1zVGEkSYxvMBzhZRKfb+BiVCT7od
c4frfbbQ17cUaXfdztuORsRkaGEvFoEfqlFN/SiGPuCv+YvevARvOS7qtOSftNNboZ5s0/y4UIbL
YqZrOxvtklNAAs6s1vZw47fX1RNGDWRWRnC6ev5sWh+Bvpat1nVk6rF96UXV+j2wvGoEYPPtNdx7
kcn0nyjs7mqDsk7rz6xJzYm+OFP7bOHhd6uBDEJVG57+ndW00b3I5ott3reL/7neQb+9gsRN8MIZ
whlonFaF7R4lALxJBJXNDBcHPWizIdgGqrPcKahujX6NIpfEk4sYvOco3VS15NeF/l/OpDs0Y50Y
K5uuFt8aqzlIugB+JYR0brDNzCamWX/5026od53gZQvD+/2dSw0uzvgJo62ZzuEN9HXTiIskIYwD
8x2BIVkrUqiIGtLeEO6h5BSgsrX8gtclDUYrPYEpSGcSAM8poln61xOrM6qDOhwBKgD6cOv5nOl1
rllkXo9DlIyHYguoNbu2SPH0EM6J8Sz1ectJDeUcbOYNgXAIeruB7OX6KpHI+F4ObhizvMOzSlBO
jXiHGA2wQoa4+buI1tW39mX8zpV6J8xI7I81K3fUK6jeRmUqVn3qGNUH5Gh2DgFUNXr1DudfQ6S6
zttXWAKgzjaMnX9oxBaHd9eAC70cs4oA/N5oaycefugPJNNDbR9vBtvcZJWa5P4bsDdbbP5C+6gR
ATQZfKeAErTqRlBR3fI3kx2H/6icWQs11ywsYuMS+p0NunA5e0qLpujaEG68Pslxz9ic+E9EqejW
xxSi1VNZ8W2JIHLeXsHSemF1Eq0Czf43aTQ0lc0CtGh6UKFXD48RivonvnRKfqoZwY3yRrPx/TLm
IOmW5xUfOz6H67cKd+up7jJeREKbTedQQtKUBjpRD0A0SHQWZ0+srBSSBbSEE4rVDBqHxWbMH4PG
yAS1g8ASPlO9pSzM6bzRPDTjiQSdAdj/u3lZKZ4RLU9QVPmqROb0MOXTFZDcG6IPZ1hDvoJjiSRD
Mz06WK88TwwIGLvUjpkdFUwwNvXaZJm+SepxE19TgYZT6rOAZ9n/PZ1ObItl3COEkTDeeulDqftU
ECIWVJVTVMS5vsOijABzsr8tlxgKn46Wj5myZdc/Vw2X8YSWo117f8XTtNDLWdXRQ/op6ZSea3TP
wMxCeOj00QOb+bv1unhJSZJc7D0pUAc9l5pNlqqryvyBMwCvy0RG/pcs1dHmjDf0XwWrCZKvr66r
7ZsjF/oW9HHh4H2S5P5PvPqWmzjdWP02XGmhzdS2ivehpNxOhOHT5MDRBk1xHqlooEGetsUd3vHj
0Zv8geKH2vatpmKRRCyb30RfmAYkWzAHUTacwhx9i3vZaHcZGntbA7UqP6aW4oqiTy5NwoHRZn79
jhDGOZLzvh+r4mHitF1iYrRvsifC8rwb7DnV9eJnTtVEQOSEM5JxjbSXHC/UrEstT02JH7Slhj1F
WksVdOzQoUHrq5KEjXWVZar9uA2iu7VKCW12npBUHs9Lb/aQEI1wUFIM0A868tc+FJIKhUX6tBpL
+1VqSTYi6OoeyuSdcnfo/PS5H/02vTnWJpLu56FWsjNKjcWihg3piCNYzBvbWAuz2WOZyD5Aqr5g
jdq8Sp4EmuJCvRYOPiK79fEcmGBx8BnGJKssVBiV4Oux/fucAAVJzJ8+FkRdaWVePHN4MqimJmM9
pMNrnSSdADOjRlZmJyZ2nQZoBGYCHEvus5pqQx+2xbnRAuI+whCe0m8gKDkqk5XQ00AsXgnFASCy
WgwngogWzS4TMRnih0xcfY87qv/QMiFSZysG0bFN8w0psgxJ5WHnuZAyglEOvzlYoq7lhDR1lgTK
im9ZLi9fKcCHlqpp2AOnCetpaJG9Zg3skQZqQivHOMJ71Y4xzx3qSXwcKSlTZlmk74OhjeRj3kQQ
Vu53OiGDCZ07GLuphPl0CX/8zO54OI2gy6BndWdAZt7WjOolRiOwSCNRZ8Y/RDewN/wleQB1zuZH
gz4wf9vHlVdODEt1y8xm4B5ntvB+Eg9eZQHUNx4rTr58WjZB1YkFhQKUO92FN+8c+yGGKVB5D6TF
62GbxG56fu6Ww5cxqsW/cx84oj7eDAEA7usdt9KP/q4e3FRzEf9kUKveQkbgJMFQmtJcV97WaygK
tzc0PGHXFzkYFZwvZEtmUMb2D5s6KdsNvTSo9TP9nncv9yoUcxsS0nIHm9lFovrRk91Xwxs6svi4
zRQPhIpN7cAMZSYGykU8Bo59UbDYtJepZj7//3lPz9bsR9sBCSnbEX5wT7l/12qAhxYLYVEQkc5t
7NeBmgM86oMXsg8oIKt3u9LyQr03pbIR+wMiIn3GBrMhSBlTVfKK/ltQ1WRC7nhNaBZcMAroT09v
6GGjJKjnimtvaUBjoBhJB8X82Ei/0apScz6OJs0dA7q/8jLup08xlqi3LatAd//On6MS1D2C1zdx
yJgwxC8gGH8uuO8HQTcGHI44ZEVwMgGcOS83FFuWrP6o3AtYn5n3oFz/HZTyB7Nk39AyM7CRL+iK
Za+lxygdewzJdzOZIYksuRStZhmzTC81ivlwTnEGYcA4v9/bxazY6BQQBom1YKYtMa03TiK5OfUN
3uZ4SP0l5oVlbqgHItRwXiT9P5SVxDCjj5fTNS1dEgvJqylfF+EGrxfhy5COxlo8Pn0PSlwHXiMd
Nl7UN1Y8ZSfP1fDWZmzjbJbc9+IX7jOF1EqmVMtxZ4v1+2tEum6ul82lNNox2ATdsAA2xv4HKa3y
tpbQIBQxn7SjbUv2HQ8rQJtSOpHB78nqTkA94Mm99ymRBezhQTYZdWLEoEG/w0I7NFf1w82au3+K
LFBm7BKuDqnSOD5L6UJZMVuCF1ZVG1kyL+6WkkEwwE9XB4mDenG3DsDlYojU2FNh7/wBlbzp8opu
iK8JAGd3Lk7Srr/NAq4+MlqepnntrQ1/ieSftvdbauj3KnqUv40HA9UxeKjxVBsto+AdbPdV8+qy
akb9qDTbQnOca5oJ2sPBtZCwolwobjz01yAKk4a4xfZj5PSKg0VMfOf9n9l2Qu9DHeymYBjYf8X6
oxJWgOBxbnFtrsOarmvyew0hxRidZIziFFn4wfkTlauTvFAr/3EG08/ksmmCJaxNBCdSVVCgpiDB
kstCxHHTnRL0zWTCDN/qs5mSdue+DHwPwfyMO+BmZEaHxTZjYwyo5h8CqNZI+ZqtwG/F73TEypS4
/o30KxXCKTa8zPsEhb9IGOjx9sVsIzzP83cT7MZltgM9arphBM4Fhuq/413AX5zpE0ntZNkO2Lmh
p8+sUJbcNr1qmHH52l+jY+rFqlXsHjsbPHbidvvrsEPM77OBtAYFsMKlch00vFw9tRuAZ2wBDsgO
atk9zqOGIyrS0RaYDALAqxmyukccgDkm+Dq0pWMSHrYT8BqgsIKWI2hg+l3ia5xoW9Jo4bzz8Kpb
vuqSDncx1TYNPgBI8VCKeR0/g2kXcgCaxLRsy6R+w6JI/VccnocJfy+u+gVfRRcrfyAZvoxB7b1V
TrPrL3Ib6M0MZ0p6p4JdTiNkp7Ru5mC7rvNR6HcZQBPXwlESO6ALdIQUQUl18EdYEmSB82ysCOCc
JoOCG3h8EN0Rcj71KUSeZdoenMhECT1eM2/nU3Quuh5qo5eYDFQQXWUf+1+tUA7bZJ3oDl0uyjA0
t42dNmWXiC1xCgAb5YkpWTXzI1th874dMa3aD6sBA7OPU/filbs6j6wha7LGVyEbBhZX8ABkP/gl
Zy9or4sG1PWBDXVCgbkAJk0qXSKVxJfhHc5VfJh6kSqi6sFkhGLya96cXKhAJG1u+NFiEQIJC+7F
POgCDSZsF9R6m6dPYt5SPQ3G0VI7fQymzLuTUHkzyQS949rJj4OVIf69lPYaBrEgjcjm9FDPQTy0
1d9umbNA146Tuz5htpc5nOOQ6C8ZzglKSbnPu6eC3z88t3g5x+C8xATTcun7io+XDAESRPaurGu9
oQJ49lt8M800rnPkRxmbNQ2mXB2UzVPOfF5nIfaMrJ2pXEjWBfoyPwRr5qXD6yFh+eiTKeeONCLP
9g2HTGaePmaj4KzRrxXTKWITS7yMlGDd5q3okAdc8cJDfL6mn6QWbIT91am22d2Oe6SFoRiERCBT
gpn2oT29bbe2mEh6c9wNMAzexrGj5ZXznA4cTBEJAJYsX7ZoUpy83fdxhJraHpjEhYjjiplQKAiQ
WC2++FECkqSFhRWEeikm6sCWDebVYV/Gcgpkx4vaPKGqNTnH7hyfCvzzY6u4AvIjNv5FINBTslpw
Ji5M6mDvt2Uopt3nFvulPsbT2S4OdyaFm+KYmP4B3Ye0tjpWiVbYzyDwCtxcMV4hEprpaWVG0f3r
SExRVzi8ojoYzmlNmFlTKen72nYcSnilHii9EDq03bKo6L3X50+Auq8VaCmG0ysnoTfk4bzDN3Dx
PPB8brIdzosuLmKYNaYoVSkbqKhmdVv0uqG5Aqi9GgZo4RgbLIVDqO79CGGY/F4E8TpF7lzYfzgV
XuLKazucpzHfRS+zUlCSiQJeipEpi9jBASZKZxk6j6a7JxpCPZBS8fq49RkwJfFpfRSKSRDTnJFZ
ql5yOjUJdGecSb3bpcIZcqR0Uxp5HXPQHBYAV2xQwUBPA7DU1x1aPI6JJ/rxVfSqUt95H1t6AbU7
WUWqKUNzNt1Y63UuieJ/FHl0p4wLMVf9QCi8bYIEK4LNRnnAl8iRFZvTzXAVAca5obfCg9DQTOYo
AoVKRJXJpZQeY43i2Rt1ONr3ylGSjRQjh4BwwAJVCNImTLaKrhDIpHmotuEWt0nD96pVKY7N8bYH
wROHqs/W/N1oxZj7yREr7bDJActbP8fhoVZlZc0qIN5ZP3KN4cV+YlkuyXK6yc64FWhN8u9ZURrk
ON03208w+6rXsRo9vvN9TYK50+6k97F4ptFkNHcyhW32mLljQ7msCqQmMWNhUfGjPm1E/ZT97uHW
NRrMzmnmEi6D8KOfHyCWuk6D1nfkYOPzepfrhD1JYKzdkRzlJeg452mKbUPbAelKgY5AZ32OwoZT
gSmT89nqOtRm1Gl3bY2Bewn74VkaOwR05BaIbKGONsHqb2BtmzAs1AZVwW2lyiM/yjPIqPD3Dmeu
qoU/2IrFuFIMB9AzkN8i4gTC07e0hntFPKqo1SphtTS4fAMezJRFAaEfbpmy14zhpLl/ey/M5l5s
fHe4rQfbaZY3FmeCyaXZN7pdHxrKeUgvIlIsUZzDWcV+ENsAWUunuckyZLq2uD7eC7psaTRYHH5u
AFqj+cm658591VAhZS/g4T8spnKZbpoDrNfEkTaxu4Du6bvkaN1xqzsihhF7/CB71oBeDXroNeTq
n+xkuSKerzFDh9coftZt25+yQPj+njsCv/tU5NcFsxcNPpIT59CCCrNFeqQavTXvCkYdEF5mDASH
OQWQLRohpH1ujOrlx4o16lrJkksMwjOO+BRAajBxAOW4TH55otp9AA1u/rckxuYLOo9EyZrDMRuP
+FB4wy7iwa7TCjr731Rwa12ZeIHyuh3+Z/vWeUP7WBmFCKkecfSqoHS+7RE6+zOUlech5vJtFY9O
/6Kz8Q7ofjYlgQElX063SgnpPxBkop0Nua3kCkgpPeqXi17zLpKN8xCw2ZttPWlRN4/XL2CiIfGV
7AQrxrRDGATowsPrjT+rJFQfsAHjuQOyXVm0yetBv+twLM0VtZP4Y3rTpbxoDxFYJ/PKCVlRUSRZ
ZEhvJKlurP5D7wA9NIz/e2OjzLy8wOsY5DmEqQC1ds/Tbc0wPBqhYUZjXv9uEG29sUmQuAWfYYde
RrxzjkstsK8w7uXT7qQ83TzGYcY/Q4k0CmhqU1aEbHz09pYH6bW/u22Eg/O3uOnVUuda0OQd7gVW
wf7KYx19UHscNWyaTn3aXb4cKymINmRyOV+x76aSbQcmbjl9UUJiiahIJn+T2ViIL0VF5q1ArDkb
31YpwuJuCtQVPeAIhYYH46IJka5RDJnTCQKNXk8wS0jVGDhWk1rl0/rJILjfCvrZRZ7or6O9doVR
mUAmS9GsC+rxApSVKtYKhh1hVQfjNXC54TQr3DkpyV9oS3deycwIr8Mi6G24TSdwm3Dibdtvab91
bfylqSJ91Zq1j6JYEcmZlcNR2PZ1DjlwohEwbmyu0sysbyVBdnbI7zDc+3lTDVFbFUFQP2SqREn4
qFGKB7VELra7+BP8k8S4bsIvljrgZJYSkD08Pc1RzEULo91SXO5euRJrgmnfPxIK/OsVvykrBC/R
Wja6BF424KyqpbcLtKxC6E/FnTm8MZz/YOCaCqHv0rux7Eq4WMPx9UpZpwPjJ1F9aWrYy1DQlq89
uzyLKG2f6cJG2IrDi3rcvL/4eg5sdqpJcyuroLtlXIDyBOzfHfyccot9HnN0Mk0FRMyUIZbrF0xw
NOh5zHI0M9UtbXkx+PnmDHEB0iY7rycmUKV/if2NWs2WdC25yVY+YAN7BVv1X5eX+J9xj88zOhEm
mn780tbOD3geCTMAKX6RU7lH6+I7/+fOlXXoLm7DERu2kuh2r17GmETc/oah27oQ2Dbbyo7axvNx
FdnhkS1KnL+5+aOBs3vQ/l1mf8SS5j8R+lJz/hg2XsKhcpmSW8peohe254Ydr5E+VGv0lCG3jdHn
pBDEfvEmO5AokdSwgwj21FlOEZovYajoOMEMeSljTTJhlwPAg1vnbpYEi5n7saKVQVSLO1/XsReg
WH71/nNyN+9gB3ERVFvHT4I85MbfzJPC+3BsHuDi6R+CBmSux+dOfVJKhF1XvRGb72+Th35YpoXO
l7hxKvBxQx/HaS/AJX9LqOQFGkeaAL5kUpvJHXmWTSFz3WqvUEpwfy/2OPAuLp3STne0wKM0Ss4P
JNNSLEF1CS2IJOix0fBB8yN9pWmoiUMROwiVezO85L5dNfT2+PmU+QGRNIoYsBeR31ajmzQ69cXG
81yLsa5aD7y85r+6Yh7lS00xA0FqsZminjSeNrPCXDtkmY2J/1VEdS2un631c43loBkI6E5xm5zb
URvDTFS+LF2HakKj/OtFm4OKnT8jzTIrU4WoFX/GAl5Y+LUQyg2vtVJ/XXiluJZUNaULrBZTRRUB
TY4bR/qdIX0N27ekWGxfrx4xe6fsaDbctv7gSUZ0wW9HLRPEnR46GnLS5guC7BDe6ppMFmHTkD7Q
aUG2sL8SYF77qsbV+z8QV/QqTYtddn4GidntdvJBUksQtGNya5TWwhsaoDDbG1f15ukrs+zELjiB
pELKHuBcSka13iDajkwCSRCfVGMcMRGhs577nKkDk1xh/HGHtMTh3S/9d8WnSHIorPLJAr9B6OBX
V55VXzf5X8e6LrBieFBEVdB4tpbdmpSn5o8PVE50DhnK3AaPf1/gpFnfy6J26Jch3dp0R3bAc2ai
FCMtPv0Lk7obVptrodtoLftCi+1qiLBiKi4I34aE6vA1v7uhgA36U4FkmyKdphV+jNMXI+UHsorJ
LMYc/wuJYpe7IdqpDtFhr7F42xBIcvCSUPQsZ9JepAuoM2F6U+/8YmRd1ylkUOJSM6CpLvndqXE9
v0fzOLmIlAxna8Q7QJXShShhcziRfK5jSQciqwWQU1/me/YsKXvSFMnIDjVwJAYaJfOtt0/zCF+y
IuRyBI+7B6Ng5p1kCBkXwlHF8XR9XkUehtzFeKXSJovzIwEqgAhn8vxeDZ1hfWP75exfNdaQlarb
8m6Q6mhGmMJfcWFORRFsnDLvXHtRON2VO3BTEBHZ/0YHrSXJPSmZU2B6VeOjObAtFA3bqysD0zmG
mmryFbwd3JJhGiDu4yZuLO4lXenp9qm4+FnLIC2++/kXUy7wzxUOBJrZwz6Ul3y0gvyhE3rUr3+A
itAOyOzpstPKHxHljIArgzZYLbwrcDvoVO2SbVhkR7kmUHdYenGi2wBQJNucAtNNMabfLf2RrsAq
pfea7vZOtJ7DeWXknHI6iBARHhfGWOqZKoHl4OZH0D3aIl1l1Qw9biywOIyVIe+c88xeZ+y6aqI8
XR//uL5DUMQCCMxjBUumZWFukynjK5IjhB1512jpjMzg30E1wZ/5c9Dcriy5MXA1dZricCA731EB
U0kZCMDMMlEDz9vll/C6unCWr/Q1gcuVlccma+GKcNHPUQSmE7kInYV93qDYrH9eKCaxE25lhda9
vcY5itiV5GQFz4chB+35i7GHcaWN8Eqgg6MM+oG3/+HUF6UggH4UV6PpRTf6T1wl/YAmhCVZHSLi
R/3kkEX52fFKCTIEDA3sTw5AGpcXrLoSb/VNIHKcuuhX/RTHL0LgBghqGIkoQLleb43yMTKujPXh
jZ7m692/dJnKTn/Xq857FK4A/bH3N1gGycDqAe4Q+9OpDx9azfxz+froiSKmw8biUXXVVl0+D0Mq
leYBOuZhqeoAvWXs6m7l14CML3gVHAyrSANfY9jJeFMzPU8sDAcPZ+arYdnb/AAuoEc4p5f38wQS
xUpR5X+t84WuraXE34CDxhCF3cjhZG0L1dF9pa5mTbWAl0JApO41X3orX/8vTlrwaPDVkRPVaWOg
w0mt0DEvwhXfshAnbpqXFCpWaMtJoBI2O9DQRBrG60VO28uzWxZ1HPjSJZvK8JXROwe4f209XYml
t7vWNwskCsC9PtWYjwq1B5RzXHKKWKZ7/hWILnIWGPRdPluxthAAjKxKfGPNJPQErFiN6HyfG06F
9OghqV0NFo1fHQDLuVGydoUnF7MsPVqc/zxniNFtPBY5nxWr1nKtsdy+W84ZWFWO8ZnMRTzf2rw4
ZFsVGlsoJrxkJ+tb0jtzhrYzscZZx9GtMwYx9y8EewgLhDsRrLZFFKpfxJwZfyhmmvjFx7OjitgM
8zNAyyII+4qy48aYTEn9tFvwsSKLA7teAwD7646DWQQiOAJMIdnw61IhHXtEQAykQGkMp9hxqrvR
YTwRACA8tSleq1k/HyiHDS4BCl8HBOZhsJHeg8tKlBIDpuFL4If8I4LqB0jvan042lbzhG7BAQuc
O/j+gi2kdGMbRhRPMG6jq+3nq7pKuGPuSrt35CLScVdsu45P8LKDB5sFVqQcHvfFnJ3VfFsu3qaT
OIs/5WtMageBbus8yZzO8twU7HBtLG0kYIz87/zOFX8iwAEYSqhKHkQvQfco8nFCQS1/bpwg66tH
jRhqu9ORh9hA/acmExhTbHhIvpqYrC8A6wB8DZT9GAByhwDHH4GwBvklX3Pv8d/b1H0fCbp/aM89
Nxd3XUq6bQ/2Iqz5yYRk45KZLP7cEsXhkpmM31R3+HGCjzV1js/pzpRauRbjb4Ts4o8NMWWoMZfG
KA0b1WgMcNXQX3/bbfhUveiW97ovycVbwYPCaYNhLVPdnXQYJKAFgBUgKBZ4E8fK5OttVQcGrP3i
NoxY/IQloYCOn+sE8wiXeLDEsM2dz1VTJzbVexiELS1hj+8W01ZZ9VsEnQ1BpiseT3zpzW5bhC2H
VewQ0HVz/EZ1Pqamk2m4T1GcTk6gvEiGtgzJRyhM+xmQP2WaGBXuhPW9K/bxeVRMYlYzvepfwM+c
u8X3zSH+2gNi+75xMvfk0qUR/VrE4bE3ElZ3zg0tpxI/2xaKxdWRjs+rKF6z4rSoZ9A6QmnIJzWj
KHTjkdkELlPqJG0IN6AbUqP8C/VkuTeZC/x9z8KWNY15fmXFV4um2LW9DoPWo7TyXaw9xJxNhZJY
RZmkujuqF7H5CrBeo15iMxArltbHzfLoBPV3hhuuMaVyBH+NJwtkT+rEHjp2Afy9G8yyV3XmUtaQ
Y63xiQNZiPP6MwBrFp0mz6lVJlVWW2N5fG+oZvv2EI+ytVeLyTk7sl1L/S5DRqJyvo3b7vusSDx9
+jY9yAgxvHCzcFt48amm+r0Os7x0uUrmYdd5GO2TO7hHl+Ifgw2wqLBuDewWFal6D9bDHXTNRrhd
KutAcgw+x7Wi473/4IuOqsdj7NxqdFRJ3G9SbVensbpV+ZaJ6gJv0+5FfC8Q2BKWI22htCwUitgv
sI6AowbBASfJ9Z2wnp4N9tMouFBWYKHb8m6Tl8m+d2ghm/3J4BSsdwECDkQLnW1iG0/a/kuyXy3x
wcoYZsPlwOYUuULPIW0DhR6eW1dea3+w68x4sVntKOnCRE7/UE9/mhmGUQS2sRFvYD1xOrReO16Y
BJkri9S4WaSp+49hJwd4Sz1Qm1IabTlUWSjfUaowOo5SpvTkj9s2XmLHyC5wQPmGbMuOZxrPhne7
fnlzblMMUXBKTAovnNFr2YXb6o8/eRjzHGgfIZkYFZwohFT5hnau1uvhZjOVsNW68TE/vvK67zt6
KjRTtJBL42n9BDXkrjP72JsIWl5if9IyQVMiWT+/gopG1dst6FrNLpR8sU/qK5YM8SuK+W4YM9bo
mCdhdzExHN46mzzvAjs7BTfgDLuxljqgufSVT5lNjPziVeY1DqAcTMJqDZBGA/sJLIa/gm1ips4v
N+djxEWt9Oc2WthV3g9zAu4M6eQwJiQk+19goXAnVaPUFXkUv3lSw3P1JF+LVScWBAZ9ytAL1tiM
bHkHf+2oX82NCNTnl77OQCRSFs7m+98F4+QtQLubiFfsls1Shi4G91dtm/VC+pM9URxBd3+PNTxP
GygSx4YNtyUmB4wBZDDG6JeMPgPWUAdZaG4MVawbGLJrGpZOgzNQhUe1GfqmhwggkANT32VdJFUb
BbHPql9WxwRuH8BsrOAaakwrZ6wSlk9dQ4FSlrUNsb68oq8AjmQtcLSX74LnUfKsuB2mUzIJPAIQ
0uPv8qIJmCOu1U2KZTtoYlduiPpka5KlXdLj+TuraMT1rMZ9LGMW37NOPvA+3lceC6V+qF/ofCHy
pveF5me7k2qXtpD25uocScIfEj3nhCcYO97gwJxW/x+Bb6NMhEaDd/EqdhB5FziiQz+Ixwer+09p
AsgT4GQ6uMFFKHK34JaU7/KJWgf0NHEBvGCIuM3tA1XsJcuE1VSJVvuxAQJhyxWfYb1ja6HdDC47
hjqu81T3WSaPhfy0dfMUHH7Dp8JqH+UubgdIy5d36b98m2pzf1gvUpb2wG9jb6OVa8qpM3qbdg1b
plSCH1PwoA8aMHvqXljF8f69+0AbI1t4+s53IT76mWmwPXOifgxi/Neh9pgB6T6KvZrnHXPW49Cn
w9Eg3gtO5ho9YzHCyD4gySE/2z+mueHxusk4wiirz+wxkNdXecs+mXJLnJKonev6q7n1wY7xCd+F
1A6J5IOhbBTrcN71CaWcbRothdz0o1bMctmPKgv+fuVX0l0gHeUpsYKNwnPEgFlY+LUfRuT9plJf
/e8UoZ7IfJmugkxGUJ1mwhKJiVvwTp3uKJeMUwiRPt7A49JqTzSgG2C2423mGL1/ADsee/UcPPpA
SuXwWgHli2XW5BzKDKRUTFf/jRmQWXNTDptBIMard/6KXjh/d4+y6yPpwnfkZmL1LR4UgqiWqoTz
vnpUUHnIzBXgMnXKF0NNuQG/V/iGOiNAbRlJAPhxoYaRJeah9t9dqypKOqXIta8QEUlLKotK7wvp
QhU/Nsx9fvRcF3b4I/9Djt6ew8Lu35RNDYIkW637FutCA4LtVnC/SFBAxfyDMh+tz6NCZvAHTA1r
TkhW72L2F+aBQ2gGjF/Ew0kLsSTT4W2YTGkxl8Dxft9VRtTQVE0c7O7UFIAhbfKi/Tnz5I1jwgjp
+oXIrRfP4ZEGuMhYPVgX/tzNSumbqOuOOv6yUXUsO6+MuoAiXZ/oGJmuDQcPmHYoykKqxG5rCLkH
QTxQ+VZop8LU3CmO9NfNWohdl3pGusZsGra/wOC0AxmQ0ef1Knp1wNITRuSd3/aqpIygW2tWx6Vr
YCxO9L8XIgcQ9JPvZU11PwOBXe4/LwVE87ZcGLdCPj0XN1iJEocOOc43lROGEoTEjweVjL2GSFw8
LGUYnPRv4jjqYes3ABeXlRCC+YNV76kofVvQKEezdxk0TSFhzG3zzkW47N33La9fnAH65bTPTi1Z
N12N4iMXG47rRGGoXF6lA6FF29pSH2d+KtAtRelTmhdyVb3LhPTIHa1OaFKcAKbToBxTlh9jGYeo
nrWCjJfnBDDTi5P8288GtgzKsEDj5vmCJwfcaNRJYATbDtsu6w8qTT0v2WxgTfW/lBls263YFR4X
idzkxlUW+GTJnOFn56CVuyBaNoDmnPasmQ3vYxtejalDN2cQQYqdLkNrEhmtpa9k+HAnrWxg864H
rRmAYVZtADEMJqOZzdvbqmlJV/ZkgAoxqae9TymSr0IpQh0XmdTIvKAyYTI/lWc/DEvf9Qdrc0ml
8VHCZoGBnkdzenivIm36v/PK+S1rsphRgA9Fc+4Ny8o7LDbeKW9kjEXMUTAuVfXsnjXd3aAy+8gh
VvTHX8o5bSkd2ZiJH4u0q3kiTqtGKiN29FCpFfh8rNcOkUBJCFPhCGoYqHrh+nFv29DS/5GtdtEv
vNCHE89/gKTQSWvBRjUvqdX7uWZErG+sLM80l6ZpqciDESLu/XrlAkPP4qwkMarl5zF9nA7RVwAY
lSalTESzgUnCNpkYRCzU9rL3U2evJcqKsO8DXTt05e9KrHb4sUxJ2Cd8JVu8dwCyJ17dCnKeR8BM
mooFMNb3haxmqk9BTVBpSYNy4gmLJaQBtspQTmSlWnaqBgNhRe8xPIM1hY3zVm23Dep6UqJQfw2P
Ay0/xn5pU1nWUMMPDRL5mK1O/LSHdo+uc+6QjfkIgMU7L2JCFAKaVyZsfAs6aMVn+PJgVS/31AuT
a7fVCmbs9YwRsbDoRx2t2xZS5v4cVe4xk32UlnIXTckvfxGTnqoGhDwf1yJdk9Z3kKriOrskbUNo
osOTVEbl/RaeMdn8nFX9FLmjEMrj7jdp3BCGE19u1ABGGgKsjVaHUVqj4ZZ+FAQn1HDJ33QCXaxx
Xvn8fbhiVCM08iCJhHillQmgAUkGdZ2l+jtjv+8uPHo52c3Aph1VOdHsrYPdFOVUM8AbSEt+dy/Z
XsY3V1+HZyf46gDD1Cxy5bCr5WWIAKsI9XzppdWzzMMjI4eoQS4LsdtljSZm/hSez7+I/l4YrL2j
TMdmvH2M7pk2UOMv/A0y61Aw5Gk7J+CaD8rUKIkXFjX1x5TLamb6+K7c9MenN6s0E1FdwxDhZH7Y
EeOv4MEBfc6HH0vTtBrGrKgkCARYhs2y++HXp8EdYBD0iyL1kvoskN3S1m6KDNXDGWfpu942HoNl
w2lgcO1MXWUdHytrC8Wse2Ya4Bf0fPu6bp6WFXXbUm2DBawI6cPe1jl0Y+G53MapNLAou3v23Wol
FihbfxX3PyMMVHr/0XZLUwaj7LZ1N992+b4bo264Y1BQ1rzYJbvx6GIBXKFSEBYjhxr+isElHySp
+UPVxvbpNVq6Ci/MwB7pUCGmEEsiPM7U0sLMdPzvv1YgU8yk4XOo3RhXdXGdS3PqGchmcEzFi6h4
78ScxQhOXWUlBUd+xxcfbj3qEy1opsiuqa3TB+1xGlfcL/klwj0LW5OtEqEVzGvZW8QZXRfSTL4n
ZBgC518ErEZZh+G+II/Kcn6YLja11bZzzkkZaEHpyw3CFcONiT0fw0/LuHXW9xy1VNfST8sbWI7+
HoeFuz3z4VUS5ygWFKTa8UOfG1CsvM6PgfmQNckpU+23CSywYfot3H40Y+Oe3gTu+DhmN3t3KCKs
BSxNgzf09kp6zMDgElIGPt/S/JENCytNV/i6xx+VnQk/2bBMDTM+f8N7OZlFynulOQlAelN/KyIf
uGskv0WQNEYMyG6z3acp4wmVRRhJOlFBcqxBYMYJRkmZq1wJyvTAvyfkWTEdttK9Hw0gMIHMlPV4
OQjxp5Bk9g5CbXdtDmN8wP/DYJLUeB2IqMPaQeFzXR+7+T0bELZU+kV3y/5HhhqT3ivrLrMscOme
t9kJXT6q2/+tjOhW+DxEKxtx3am0lS+2VOOqlaYRmdcARPWVCWA2UHnGv44FYU+ckf6ZcvGnda9A
gqJVwtt5lqNOqHB5YBJMyZzkpp5fO3/eYgBKVOc8yq74RsO9ecmHmRSyUrI0VHwWM9pKyZPpXOZR
nNJKTMyWB4lbE8j3Sv+DAARGdDT9jHvT6KnOIHc52vasvu9a98dzrykl8muwBpWxklt/7Aj/8807
08Ja1nQDd3w7yyHrBFsRIgQ19s2rkI0lCxCMmxfv4zvVrGHbx50H8KSQgC//gMA4te6x9hBFscpv
MyuMpjB9YXyx59KF/IrD5iqt3vaNB3Nb6X9yVc8jx8zFzsgNHQYbj93aJzFsMDK+dqFzL//1y/VQ
OZVyeNR6px3W/e0ErpCUoOm/hWYX/0G3+UKBbB2a0xxdmEWc7zLzFkzyBND6Gi/MT/mNvscfOImD
lDTQiVl6JaXgTKqRq0fDCOBPAwwTqNl5RUbWXgk1IXaoZGzpt5E54aL+t6rGuw3AlLia2bHkRblp
dZCD16kn+g43FYDBoccAUtN+UrIgxi+mbRf9zkjS/+/ijUQQZgWzRiSPWwOzwdg19WCy19r79wBr
g6MHAr5qfhCrTLTYstOoTh7NFkAE2J8L/yo1b90prWASDtJZC9VbNYgzeDJ5Naoyf/PMViBaGddO
d6ZvbrD3siPy487GZvSemFUt7jT4+WcBe6uxj1nIDD1Xx5DhlCkKyhjoGvDe+RhXgqSk7BRCCzvn
SLUQMlodf8WxcnprjrViGE6KIChjCAWj9Jbb51B2Z3tgEAEvXgvEaUVH+d/2cf1CfG5QD9kPG1Qs
qGW/AWwi3VL4P3Tfi7W/I0ArQDBOrdfVajJAlKGe3np7nZxB1ZEDGW2wM0UAYoFI3wrWsYoE1Rr+
lfaTR6kwvpKzBH6CNHUowNeYt7+vku7yIw6yfmIHIhMBGkT3dGbujLAQNBhgA/lYjQda7rXFZLVc
JIEe0mqd2KlXP2Ec3zUkqXfOr01ICj0LwVA8tO59405iyb820TEd+9DEE5x7/LlQLQRyCgPEJeIK
RKNQNIwXHJPxgNmix2NNyeQdX3E9a5TEl8JHo8Wj8gBIyTsZSPxJ3lf3SQYEFpU79booewjW04bl
ohccPJCUSKPoUTewAyXAq7vVSK1bL6IgOpjXXPqwqfzfWB0tm25oJMkUhtffELPweMucTipx9OjL
nKe/kNsDlJaNT8WrOsDpuF29tFUh+/BwWUIDyp39hRSYjDJhEv6JE3m6NSDfjD2ihlj1MjB3EZlZ
6zEn7M8KPtMTa2R8OVwnlgwmbSouGX9B+hnr3bYuQ8mHtNsw+lofD0ePrJNPosSadpU09rloeBfD
0jBAxfb7c67FaOD4kinfhM1gwbCcmLvUsbIhlLVKZzQOsuz9g63zqHZc5M+UkcPcn8pAAE3hEKco
W+Vf+FnJ58NResvPUYKRW152fa22dYTSZkaatdNTS8Z+PbN6OCxowWVJT6qmQkZJjNYEnCyJbMB8
4YRbzkm33aHdXicZFyI/DHasrrqidF26jzW+uwqtGE3dnnx8D+lKP0GK4rIW9v/hCJWhuKauAFcY
Su9x9BWHFFTI0JG2bkbrmh3qMJj35DCw6x9Uv+Fk6mSP0Px4H6OHuuCAHlrI7v5PbJsfQCGQ9Bwo
xjCY4em0rVg8IlTz772KXekaXI0GE/GT10KNh9xztM+kG7pFF4joyBySsfBNYNwHpsE0yj3Adfmv
pJNDVw5o2GKkaEDLJSZU1Xf0zDRZJkVsKUM1dh8sUniWSa4VmmtUmM0tpsF04B+8rqVyki015Yo1
9fj2p+nbtj/VZLgoyuqMiETIX+swYqFac+n15SopKrjDgo97vfLKeHCIQkOTpP77dY8x8RfhTACP
UuEoiUF6gRIp0rXvpsWo1Ok2oZlVoRgOS/Vkx/fZWp1E8BiUD4n7FmqHELlBe+Pt9ZgvZUYGMjPn
JnH+zGPwBK8fie2XXBv6NgRfo6iGCUXKFdEjxhcXOPGboXrHOEixmPshu0Ma53juUqYf4Flrdo7I
ccJgVNBJB0F/mpYwbv+e5LnwoG7gAOguZmbmSWnRVmRKdjlgR/rqLaGmV0mvr5/PS1YCHyjuyzBF
7xQYrHbgvbQIwOhbqD16f/fie5QowkY6A/XIRIpNozHagtC6YzDZ8rzGS6PJ49p/k6Ik8WlsgZxL
aNl1ruBLr0oxug4ArjJiBrihUESmXz+uraQ+DWVh4Mv4/HLqUjjy9IwNC63thY/uteuu3fHN0G0a
+zjkw9BENG6rY47qZnTMEiJjDAAAKQ4gtvW44FVbLmWVh0Gf8D2oMumHTIme+wUFMYHR/N2FW8nj
XCnJ2L/pp9SGFw+8Oebqa7daGqXAk5VdqNSQtwfpl9MkkIc4qWkGLmKzrPzoMfv8DbtDkL92Je2z
90NTeKOLPynTXYX83aT5pjYBYOpedy7A0ynpN77RlV6XIsE1Yy6hcc1BfIHVMEuA7aqNPRgFJSsH
6cQWUk0AMrzvI3cbDdP9Oxo5q+g8AlmzlvP7PNsAbZWFq7yNocfAxgZD4jnqJsuFldvqwm8qqxv8
67BdHE3pQ7etfdRnyVzxhMej0TVR8F50wGl3dT8xpUE/yp2qFmgH7JZdnvjmTII6bI6STZ6zEwj4
CgKS/52gWxAxVbwIl672c3QGfaULCKLLQnc+oJAO/Z9/RVcMiOLFbFT2thgXzc1rI4ZsUYYDlJ64
HXLf1sa7u2uxHhv6wh7PKPyxBtSkdsgBL9A/RrOuvS2Amb5s6hYHRCK8JH8lHUzgumcCwE00R9+O
5gSa60e4edq7g3kmB/Ys1LXagkak287h146w3crg+tqQq4lCI7zRr36wwRd5k/lMuQjCq35pKShX
4y2y4f4lDYnlsuKJ6XngrRF8Ns/9H8CkO9hq8kHHSPzShSSROXAsZQtcVj+kPwLvqx/T2nc/YMRh
JRiqsjR1WlAuyfwqScdjVBjsoLRg1tgfQGcTxEZ7lSr3NDVPpGKEVYgeB4qGlroXEtjr8LBau0dA
bF7lBv9ME9zLh0+9qv/BhQpLWb0CmoDjLbl8yl+lXu6Zov9YvySUyMIYO4v1xf/iWi7Htp0IDW0O
856CRPV60UMlay0dpYEYh19aYZd1vuGMf6evixz43kpIRwhM0KvlXCFbgg4+9mxftTeI0beFwrUJ
ZtGZxCB0nMWdeS/GsA5YgD04xdemltM/hRkDatt7heVYg3Ylpnfx+KvReSgwjWsBLu0b+s+jw5zm
x2oVU+/tN9F2QbVRR4/IFgIqjowMd2pQlu6zEA7YA2UNCSvbVV8llD7yKMbw0EMDvJ9Aqfn6tGhk
M6Ta/7KerxulOdHtBHrldoyugNZ96OJSBLSDh9ExqqSlu9CtE+X94FRlIjgzFcE+UuXaZBDmOrls
VnYESXt6gGB0BUlbA7yDVymVy4T1ted0p0o963QBDDdMjYikJUAhdijTaDFxJYcuRxs3zP6Kgwfj
fFjlx4+NeZRYpPZpHIu9I4IG8hJkEOTPlbZGaVQKOucUuqKiteq4ConZq1Tq9V+UQgc6ReTh9/wr
T6Tl3TNTdqScqTj+Z+Zd1JCDqZ8x2o/74E5V26aNUEMQIETzH+5vG5N0i2HGwXptWkq1x7/ad20U
iDh9CMkGFkRK5Fz1yObSBMfP6t2+K8HuyduQJ9HYkNuTtzHWzmmOFe5CZRQDmSbcVfBg2d1Q0h2u
zNZfl2qXO+n2uY4kaD+n8AovWibygZAB4GwQTr0O/2Yi1+okZgIBkUtlhFFclg7L5jJiDtAW/h9J
1yteTnCGGBne+3WCehjNzlT8oc9C925xCHADgJenrEvOUVf7bM5hImrrvNK6e/rpHNiKyOmoEbUy
bO9hEKoYyY1D+7b45LfV5Z6c+m4hLZHT8n+gDMwxD6JkMJa/ocE/cdKL1F52Hr/VNJYIHgFXZyFy
5rIZx1w77c+3PfeYQxEavhwgwY492M4CMaJK6FUqtsbUBQiFytuiKYELr6oiN77iQse3/ZpUsEtq
b63P7wV/maqEWP78zMxsGPmcidYz0KzoS3UH5MWm8ho6RMKhFAxZWWKT7onBkK/7ZCKeQB4TfdGT
P14XrV2Azg1/kQ/ppZfDnjLSBfjrj2R81DWlGGJk2rB+roJmixTji5pLSZsWxpcOi2e6hLmBlIMx
sbjPGP6w3YBZbk+fAaePQ3vfcbd2qjLa6ww1eHr+p3he+jrsrHL4jtdvtSYt8W+YksaC4uizQN8f
Iq7bPh8EQrBRUGwXbHKw+s6gV0HX+WVNJVB5hgZ34IL778JCrgv1TLkoIdl2PV+00cCcwFP1fDvg
YyT4EOcjdvmgKYrfrQjNJgVE+S3AdvjBg3brHGjUzWuWkax3osVVX5Bq3VU+zVrh/09Gsm4y0hDg
AzLx3z7UHonKaVZrFMRR3rCYaERYlwGoCIUkqiDQdM4W1qPXfowUT0MoPt1639Tyl3OZWdOLLA6+
TctlcfOBHSJz1IzklE3xfrgwhEYBQ2ItNwT5ykh0JH53xwqqLTTNObnEaykb9LmsTbuUP5thB66x
8M4xChTBLHoDp6wZ/VF1vjAPf0JLljXb/9w4Kkom+T6/Cq/umWEASBkLZPtgXWnbAH7kvP8uBfMO
6b0+Db+BjbrRAPUMWc6MqssHXoXFBaL4w5Nud7a7EOZPeiDJby2YEl9r1s04SVolybDEBXJQTelC
K6KFnAUCHVwHnXgap0J0Ep3XGp/UgeH6CLJFYPmI4Fh23SrgeVD5ltUMTPhL/Aa1N9hqRozrudiL
9R6bcZz0JEK6O26Y/RkUVMRYnXGNPPTvgZWWNvKRHQowgD0D6PJLqsFyw1TpiiEMGI24v9ZC6QCF
tYVq0icR5v6FnsAyScDzn6USM4sDOQ8Xj1oIy1nn7n7Uz7/5vr3KuD4g9WdIlE97T2sYjMJ432wE
jB4S4SD5C36sTXb073Np+yQRoEZ/mWPMGeux3rerRAJzBwZNUtyxGziOOrJXIgzdfDNn94y5zeU9
M5FhDu4hSGHOG5ehh4LE3I8ZJo8LCNY8c2XDbdpwZzUnpGUCHhpUiIpf2HNnCH3fxy/cj7fWK5RJ
KJAATR45b/IillZXIr6pa7pzCQ9TK531lzWhwlnHxz9rlBlq3RSM3z9ILZ4lFI1sRX4txOJXzciQ
qqhXZ26h+XYAcBLNuKIXOVX5z8xYKA4niYN5a5Pz9HRizgNH9EyBdNPodpe0tzmXTYH6oO1y/Sbg
X40+TkxPp+Q0z943o+Vx8DmQmwwnAow6KbA74X0GoVuQEA366EaFoVgMmMm5YcuhncnDHKDVKI8y
EYe4DuXYxGJAlVGADncqIUfyHMDJ90JMRRsxosCBioG87jlC7l+Ny1OEJSmNn1unXx2Hhj01pIaq
RtkAi5pulGemqwHQQHhhLEAzsDij9rHljOsSIFMpZC/l8a64Oeulw2PfSdG34Qw8HR5gEO/pxWrW
ntzcVrVWgnlBT14IRqLn9CdQvM/6FuT43+Z/O4TDnaT2oNJ2ElZ7E7Yia/5qdh2ESTWiVWkmkEhb
b2a0MqYwtxC3v9RHthTvqcB7iK6gr32an6RqnthwifuLM6RO8tIwyDZFjYrVr2D37oPfEuqf8cz5
ogHi68BQBmi8UqSN+/ce5ZMdmgukzovk3PHQPA/Oo6UzH3cF9lFG/n8+c4vFLcJn0xPsaBkSj0fZ
AxzSOSOYZ7v9DjFc41llVCSycrjKn5M5HfdavsktfH1lxNtz+g0JhhbwyK4n3n8Pom2mT+Urr6WV
C3LuBstrJWt/IlNF8Pw7NlWu4hUTPKsMa7ZWXrdWQR9XYgy192UOA4yIb8+YGC41/Wy7YwDLPYy7
L2PqeQDNYJfAOCErwPzXyuhboxCLtPubdzmXbUhy10zCQfdzWG7XSnh68BtVnbkb0Fm/4M+SCRf8
jPehR0+audAp9mRlgO+C353tPT/G6746dXTYLmRxjvcWn9v0Szxgx2c2Upa5YhJ6zN5EePOyOc2P
NH69UMqApQyNY7ZSE1dNnADyaWpc/6ooCRw9Aegq2aCtR0THH9g6oCfQBVx8unGdF/9Rjt9ujkT0
83GeVRVgWvGuRad17r26nFV4VrmWsPGTrwl98ZHZvoPLEPxwG8gIxzxC/+yYHbKJLIlpVeyrixY2
NWZIbeLacY/NPGnjLILMV16OSjSlV70Xv8EV9XBCm9I1ufjXczFOWIO3+FeUQlVJF/Qlxwl8U04l
tFKWA3KqFq2Pw9+XlzqFwGpGQYKb5U+mSWZCsvqHgfrlt/nYDlQ6u04Q740euC7Niu4scYiecxIW
xFndTQEkHz7ZTwQ3pJjYGDCAF4Ew/9ueKtzsxlARIkQ+xh4oELN16yZLt9uavXL9ia8mOBdcP9tp
S4C9UJkJwrIaM0xLUhKfV3Ndi6ASeDqMxYxPpP5L8j2QNlHvriLbeJls3OC//PXdBVgN6HXwsa5n
TmZbfJJIWdRXtkyNix1+Dt+JRWpQAFlFccgX73Qb6V1mARNbaxILubzjTOQhrbDtKVCdCUt5INFO
iXWp9H1dOrCzGGcFyylC05i3vehu+uD8NfsteZ8qBR9/o+WNeTKca7URokLXNte8qsEQ6wod5YGX
YpdMu8o5luVZVrZf/Cg8KLTuuGvzjbBx6xWqYhkmI5a+WqiY9tiIwBQW2dQsMwzWDy5nbLZv3ZQk
X8Fnth2BsM0MeoNMrZJovG/5ddfV7OxGH4SC2F674Mgc/V90to8zWuWCu58xmbsIDuoDmNFVBBsI
3wn3dpDdEMACmaA5eevEq01QtGzzNtP6MOvLyHsWF67xKNDlLB9AshSjuUys+G+wWAETDQNveMoC
QZFJrLxjsqyNXjnpLIeAAfsgxcaF+OAROlnc58Xs0GZtFOBoYgXQVjlVB6BXb5K9aONvVanCeT7S
D9lhYN38rqlbnqFRsjJhRn0wjV1UvC07ZPEi3yVbqCJOTar0QISFATkzV83OSary3jbCuRBFYN4F
HKiZ4vwhhB+i3WoCpelTSGUFPgU9a7nvvpaPSVPOVJTPJX7uLK0Jn3n8ekWJ52MnkkU8KsY0NFCb
mDNKg8X00Y5+7DHL7br1Os+99BfzcJj21u0SwcrJZwRjjaoNAyCeYeI00ln17ceU5bdeJWvUOj/w
MCCXkZ0Wejynig6G/OuE6aYHdUyVB7uYjKQdqtun6V6WUg+TZd77TfP306q5SbUyzppYblPoNr6o
q8sdfOs8yrDdYwGWU7YjYL3dX1dopJoovezD9IJ1n1op2m3+zm2leEE3WDWffSEOZy/XfodmBNgV
ScPdebOS92BC/Me/auaBMGhpx9ryeyuB9yiWixmgTS+HtCJGv0GPXrfK62A7qg4sK3Mnyn29+PhD
Q2QW+nqd7URyMqTFLzlLLOUhucXONmpVyA6nYb6uZPvhjOllRIWyZg5UtMgMgpwC7fvB3IDBECVY
/U4WpLXQc3uCKPp92PlE6wikBraIH4sKPNIPCmPCk3dwxe2OOdsGjznnonxUsI0O6qov7Rrb6Urj
KCRunqX66L16wSDCEmCfP+bAQyhJnm5+2fup6COQWL96txME1E8p8AtFwgoDd5ozA8q14u5fjN3S
yr4Z2RLvTzz7CufsFY4e5EflJqdgDJaq0Na5psFDWSnbFcUMhZRa1LW2SftuTDT7epmDHQtPcgZz
MNZyvpzfDaDJ4jjXxNtOSgh8nhLvUwFnMskcteg6AsXaEn8AxKS/IDlubwIC6GDcerebX/EP82Tr
igCIkiOj/8taaqzWh24dvKu6lwKEPaRbTGjsVJkUOgtUFDiyBPQuW9W9P0d6CXa08vu51T+ZxBAR
1altKW/lOV77TTzabYcDqYuEzEh9B0FVzCzirr9Wu71MGGbjgyu8XAsj1HzzicvyT7bm8+zp9mft
mX+JEGzkmL4HSWR7N4VzCStgemYF7Er2DXYuTksKFK6h/usfJEioJKJaQuLfCG/KSIBtmsdd2sBr
I34b7IY6hH5Q3zC10kW4QxoHDR3i/RUYUUxZja56GPwsfiPEzlXY2HcepfTsxnvo6XsoxYC+NIth
zbHAg/g9eXpCC3xy500e5yZb0Yjzeutwka+MKiC4cbhV7gMGl4iWulxWRmQzjYuFwSIQ+qHELHRI
NAAf7dNjjdvH9uTwZPd0FdNgGwcji+cc/W4BIU7PzlME//07VhmsazP6kiB9AShQf/srPmmCHEQ7
FJCuxIk5O6HduAvI8S2I0W5cu9WFSoIBwDdTftCyBvtv5leCFICAIAB6tWS9oGvSxP3bDWDKMe8J
JW6OZvyeMQ6wglyF5MoW/bMiatoIc1170kk3D7yB5HtROXcRAQx8k+oeDwYbPPVg/qpblnRc5KxZ
UvlFHh7sot9GFBHn+oHwuoI/y9Aylc2ZDLqXjVuvcJrqVvBlowitGMIekAFhKx1ADgDiIxUplFlR
DUR1E0TS6EJMrbDAbMBefq+tnwU4ZpmmOr6BO3mkM9d/JJi3APH+WDKddNK9wQQwoFeTeOjxUqWn
fmQubiWVNyJX7w0PbhZU8RQbzlIvsIFYMey1U2yin2qWhKYJ864nrjh8ctYQJj8S2uLcx3mlnFMt
AAfgVSIhtkFzpxpCzJiAcf2+zpFrmVXVjl0V8P0M+411uzGkMWeDv0UhRW9n27CZ+SW8FFWZb58U
5zPNG8cKptPVhXdtb9HXuXcyqS4Y5kT4WIkRpK5gvSDBddPGYnqudF4CbRpimX5pMd20i0EPLWgm
12yuJkz5BGSACp4lCdy0qij7rjdEEHiIiXJfpXfHCb07iHk27XAahU5QzjWMlfS5XNj/smFsnssL
751lbqAqCshcEOcaRujH/u06G6vsAKHP/i5gO6EQnefEgiYUrE5pTXwp6SOnfHODdJ6csv3Vp4TJ
nSkGtQu53vhYchkWaZRc8f5ZB9MoT/AA6alrnH2hFIhAnAMW9gB4P4dJI8JFgX+0PecFIG9KgYRL
AGj34glUsnUgWC2Qhmtt5m+OcatBGOhKMoJize1uB5AewJAwWbBwEwijc2dakuHOuzDtD5CSnUxs
rtzHGe6VJIazh35P4SOw/kUwau26kKDLgWad25Nh4q3FMHlInEDtVo/7pnQXqjhvWM6XRG8sdHc2
qxxnUnm336TORaS3pkFNUPUG38psez6Ndicjf1vYGRK6V20u7G5F0dUlkhZfXEkL1VR5qAIxMJKG
mwnm6ESJvbX3dMs7Www2rsAZupTB7Nud6+1MWjz6oheSztwl3aB/TWadDSZjt1me8Yd9W+Okwt+x
qqoLnDv+syzJDWGJh0K87ObQoPoVs8QhcYX4FDu7d7A0DKOtMMoZGwb1DKrvmQWnV/rN+T/CNv8d
9xs8tVx1cVyMhlrqHD3Hqpso95H8NmKdmGxwBHu0DmUgipKP1abGkZSvnIFFr0IhWyIR+RQUOoaH
53PxfbquIKKV/UdvlafICCQDXszYDJtcLzlDUL5oyRpgDLxI9OUVsA9BPrxmZPlJe8Cx/bFufKK1
C5/N6Hy3fLC/a/7uNZDrmh15pKwW/sdoyebrTG0spV9f/ZazsklKtAXq/M1Y9UVwwZzzCSLMjsX6
dkA/5gKmPkQVX6PK5dPfe+DIupz2oArqFw99+q77MadBDo67gIaK/gD08ItJyBTIVitaJu9BGLYk
g5a8gm0ANIMDFZHfwQPETDqKrXD9VziR4X6/vtHI8mRDFjJ2VH/9SrJ3ILvQ8AI6WkS5uPW/FPLG
egIk+xRoqCWQ6YZhlveIf1K3J733fizXWvppl1S9FEOYCOro8yVw13Ny/l+T2W6vYHUcp3+xviQ+
4Sw3pXlrBuowcSOjdBz4tJ5ikWPpaThFcjAZWUmF2hjBjFdSguVDv5t4bqEfVk/Pc7FEnjdmXGj+
OaRpWWY48enkZpjH68tBq/uOXcDg3i/QUFWAp0236R4Oy3cAiUpcutxP+P5fg9y7+rgN8XICm226
VgtJc6S3YLw9P8OOYDHGfZfs6RLjo3fBdD5HG2E7EYVrWLJ9DTfhD4D0xvDUYa5cSpMgGSVvWdyT
GOTz7W6CcxuX+g/hLIU/5Uus6zw0Qox/kD8jvtGcGumRMJeAhJr4UfXbdMe57gzjaCF/X85Is/cG
Q5Q+F97ZCNGmUQD/LSd35d2kuYTA4aqBPo2WJg7KGihsZZ0ZhRgFiVO4DYrZSfF0npSZSfI95bOl
aeBriI1T8W7lh4XvE0Xfl4YdsopDh6ZvaJavuPYxZAfaQk3PKCKe0ST2JC0n0WY0EZeB18rW9AXY
g1wQtDqGRTUWLVaj6aVbUNnjKFwPRHFdsjmeCgjQMoAVV2xwfO6b4rUrxdYu1KejNjhYcKUIIsO+
eerQTRFi+YqwsPvzliLhOK9hBrPMne2BhjFNhgVPzywPJIkfnFNDZlIFdimZ5uFWcwKb2Jw2jniP
EZtGA2ZdRseRw0ovreHncb3VdpHgrksJYqBb9lFXGVy7rFJNWYvYY68MnuI597VQaUdXC53PUeUe
F4s6JdwBTN82XXu3P1mg2dur/wQf8WzQngkCvwiPDFW9tYQwq5Isko4dr4cxTpjNoekN6gcqxMkz
G5AccHnKpDSW2VDATu1qQGojvsgG8faCRym0ZzaP2CATIA93enxgJJQI6GynNEflPi8XOvrGHX1j
2tr6TSNVVRpFBNY2cdW0ywGILn1c1Fwq+cwUeX9UjrYqjSk8vE4BcD4zScQp0CaheZKRzmTOKZ4q
zZxX0NJRUWJBAIu9cRe007E9BdrbxxJArcW74zxKGi5O+mrSLjCBlcaUCGvGiDciQ8gKVvOLMngO
agKpczRsv3jZv8oswq3ywu1jcoMkhjR145EurT6OqIgWwXyrjtQtI1jgXa56Ji6Cbp4dUru8wsI8
dQ13H6buu17y4SmADbcIWWWzUFoTQpoD3NZeAtQekWjUU0mh8RmqhEHTGqQCQIOYssuy4zwvl8y1
2uW/ms147ijg7L5AqV9h0PyKitiiAjphijadjlnW6vKEXkrznUUWoapkYzSglPHTJaeXQo5L3cMT
+CVzmx3WcWwadhdc3agtDhjfujadvW8cpEc7VRvezeXkh0dOIJHCk/kqKPvoMA1hERbhheaCp6lS
gk9nBL7OIb+qvVqoEW2awNw9SDQ57N2TBCIU1vLA5AQji5m9P7dea1h0KoUWvZPSfhqcJww2ZIHg
/1ZBCblI4/3BRJq/Gzi7gCwb4pWPkMR4JL14+FKDOR5VjBrnza/tt1jt55pvIrDxzqKcF9OhUwYI
Pe0JeVS3oNVfWSqLrjknpyGJ5kN78Put+aB1tDm96tCDR+PlaZa/djth+hYEoIa9dFIZDxgxkAX9
PhGCm/I2n53Zt8+pMsWSTaxPK6nQJ8zU4gwo0utkc4Ql/ej9XICZG/Ul9G1jlfyJup22KxSrER6K
ptEjQBIr6S4Lm792MLvm7amkwHnlal0y/HfWZ4OnY3qYsFZ/Yl72d+BjkttsLLUDzVQ3rUUIOhVT
11Yk4uoR//SSF4vACV0XsQpmNIJbknBbpPDgGHrmh8DkSTc48sWkBzW1rzlgndrPsDYVD+0PavIz
NzCEJscp/V4JmRzhTshvT6Nq52lHV5ruuvtfDQRQI3de2Q1+cXCA0s/s5d7ZuhUVgkD3LvulxvBQ
RcSk+S9ZsvkrMaMQdMGdVxMTafo4p2CKkMW6aI85bdvd4Hh+K+hWWLvP2sq1dxKA0bZJbDrr1q6U
3tkCORv+A1h1hriKS8ZS8kC2KFEeXuGF8f8LG+kKmQNCyx3giN2yOGSgXmlQ2Yzu2B2/vs80yJ0b
jqTq8WYyvmJR0tWxwymlzAP/c1AlFmyIC2Z2BkotmP66igijt+VfIE/Qp8uLaFHdQQ9mSmT2TJg3
MKg0qYUZadsAfjkRHAOXeaXL3/N0mSJDq5xkXtMBWZtz/xSSmT9FfN5/QkQzlTowmyvfju+niwEp
vEFYdATVXM5ra3/JkIs0paFQ91o2BFL4h5EAHq31WRNIXEUUzEg5ipSyN8d8BYYqD8PpaBQu7Eua
flIBIquis8eeaR8JTLo/9jiGC2narMOeaSE+19nv3vuD8pp12CqqV2CgxqXKvoRaZS6TO4INlBjA
9npSp++McDpCxHq86utSq74rpBpuTfUXzkrJEBe3lxJFcQgUH+s2YSVF3X+JuaX40WRhDakHhzRC
XRcn25z9mmWVwsnCAkQhwPJUXkdp/crrEc1oqtgPz0EGsXQhEGq0XmrD4cgGKix3AK+M5KJE57iu
LtY5oGMGDA7ePOcUXo/qgq+lcxTPopWsgztCNXxC4tQxqr/bAKusiartOM8iENXbgEXtXv9Gr3bv
PWGTTrVRRO+WSzozWdDTXcxefLvdRnIV0rDKK9aum9Eg8keh5CWoy2CB4OeIKQXFj7dunYlVdF4b
r1TVCPlZ5XLCIArQrbPKFSUGhWYtXQnwV28pxyFZq7TMPlmABN8VrHKWi0vOagzwvwsVcFoJk+59
Bcj18YzG1oYIwWvhjc4lQvo0of5oPf9mCudQkLhP+mczepFaDWrMY1tpGp695P9feFrnv8pDtmNb
50WJONA39YUO4kd/kH5keMpKOZw2jhlpIQ69cehmYJWIoPuI4Ze5gcwIjgPgVyLLDUa8mkOvtutj
3FHRN5Bsr8K4+JxSvSJ5X9nSnQXn8CXi2wcmMaADgdhPAHYsmCZcEldpyBjXqBd6cRkIFlILs7bl
fQksgYVUOQ4OUiDl3vefGLTmJ/8RlR8B3kycMF5TDhIOeuvxSLRkzotLMXFY5JQHer7NE5Z5iK76
eZ8ZA9kE9BH81UtG9ucmlb2q3mR8eej5Rc/w5+kGquPK7mPquK3BJnv/Nr5B+XDkgsFsX52y9I/Y
UtrNUJvwPtbSSNBTAC/BOePeG61LWFX/8Qb9RVKloHG8xThVybX+71cgjUVc0efMgPYTEqZV+8/6
GzEd8hY1hfyi+kMe7cTX26j1KqsxOSz/RT0j5bhE5yRCUoD19m2DFtI3nWJUkeW84QVOnJe9G5se
HSVLDn94iDDTD7WG/E99zMR9UyWv6qEbROfbk8L8uP/ZUzDYjvJrryoNdhYnv+IEK9hbwBy5vD1D
J+6ShLIRXVWBA/GPdyT0xTBhr7l4z+01vtB1u0oxWwzDEfCxCFiAijlQoR81alOoNp4e9QGiNN7z
lQQBxw5kOFFZj2c731/46zERTQvi12Wy18rGavHHki2BqCbzg8W9kCj39FGHu9otXzF67/kQxsGs
QgEyTH4NLHrcwFvQldHEDsUiZcnhapmYrlm8g2ilj+xUGaPw+nSQPgV3rtVi7q910H+6iBP+Pghp
Xxv1A15ky94Hs5wZ4+5EHd3BvOdYMplIsXINm919b7sjYktKJM1ZjcRilTEyKKp4Yis7KxZap2iT
XVcqaR4GF1tK4NmDaO2LNPdasaOAZwsKlKfUWe41MyUYx60baqQSa7t/WYg20H9OlzaQkhX9ujIf
/n8mLy9WKLrWAQ0kvOBwVkQAUoU2IRG20fXXpt6zIvW4thxj/DOTaTjB8DZ779fEM+VeRiNZ2BfJ
mfSPVksJIuv7qDfGgbapPkBjaDiS9IlqTrSjQpEszt1iCAgfhlzjTt+Y6MivxN5p2wAgvGEUXBBs
a18FayDFLVXedcB9dMb9FN3yqAV+vN+z97F4iLaxK4LfxHTFU9S5FWvdcihfq064oyJanBG/wfTp
MACtp4RyzpWdNSAQGcnJH9uvQZTUOOBg38E0pDDg31OoCPeB00cxvY+E2hOc3qHN5qOMqZZIt7uf
XNTe96spxFJdYEwb8tvmkzUP2QFy+2598DSSuLlRkBHm7qgBUrWfWSxulUHao9ux4uJ63GiMd9vA
7qodcdUGEax7aD7QE7REgTdcfjXI4gMP8Gzxu5HT9yUQnIafxUXLAjHTSFyrFYLalPksuk2+x1Nv
HwVvBKRwOIZAByGM3Pq4KNGI10PfjP6KFPkrASTMICOojfAQrFmvh6ie0FStRSwKIUwGwR0cbu9t
Mp92r83Ysohx0bXNvkTXZtK8pfBjTJWwOAAQMP9Hn3sif+Pcw2JsTF7q4pjHK4TczWlrJzAfl9sm
H7SHoMiOM1/HNmcMY2hEi0iHmjYFbRE3a/0hU/GU5nVOpeYvlSOTNw7TznTGJJfWQDF+kZZsZomx
2K28hkar2GHmQzD9WHQKV3pth4qJsh7ppeqXtaAFKdB397vLSxXJxcsUUTNxItqwRdGT9Bvlu6+1
apdD9w97ddfQB4rRlw2Ew1cyiLF4t0jy9xse1M/aIlbFoT5rcWnDnTN4X2wi/can2EMsHUU7jTsD
2+C8jUcU1kbCTYPXr4pcwiG/AlIuvAsbdLUkP5NftxOPCBCIBjlYNc+OjVUWxIFmR/7/DwpG/218
vsZKcwk9SiCX1alACebz7QwDWQDv51ogbGb4iPO3908rZ/SOA7A4ZrYWqOJpgSS5FreS1OVmEWGJ
5isjTivtH4M3sfSlqsz06f/UVh11Fm9ppbK3GvJ7AG/zr5aJzd3E7CcWUcsZyrtPL54UbIOxRi1r
Vcqyz3WJUAVSoAWcWbF1u2tUjHuqPDZODeQJvcoQXe45K8isrglS3tj0fTSRglodaWamViitlkRC
rhPvy1TbSmgOxn0VMySQJYoWx98Ff165w3fFDeSdaTdvptAp6Po5hIMFaRD9RZijDI0Hx5BvI7vW
qQD3PXsQozdfhiaA9AcLrVvnG/u+8wgBWD2WrWUfojVCZTLoYGXBcb+4kwsFEEwpy1VAbe/Cbjny
5nEToLOh+54xdYQJjOle5rdyAXrhwMVYgTXekN2PzrsYMjdopRGvOjoD15lDgjgBPdp30Fu1ACFc
2lAPanoCfhJQB+tCFG65shUcMv1USKNmtKfVVBYnKqRKLq1Ki/BnOeiIGdGjUHeqpUlhVrqRWuOj
AsZO+MyRYHAYoX1nKz8T1dpZSpPqw2I+e6+gBdp6jj6b49y3+CBqmUO7FFETVGvLJISulmoZybeS
tU9pWoFIXxJAnFJAs+oVWm1awY1pcriu3g2N6Ed74CxdMzDqlTG9eJ6flkREBs8uDhGuOw+VxnE3
+4ZHNBq7vhltLC3r+qLg5WgK7Cov7zr7uzgtbm60Lo0vmGMA8iSXxKXev/Wo1dSN+GjimCmjDElQ
2wmrGbtjMVoMj99g5t7XY4QX/rTI/LjiszKXlAteGecT2gnQH9Y6QtvlJQJC4z36K3FJBpT/8aLO
T34exy4hj0YvxJDzkl/kfpFRbBcnwnDfQP4QowR1LDOIL+sgwc36bKrfOebQxvD8FmuXj8YSkLul
+nRYXpgxbguVGX0p9Y+gNNgsFPSaF4WbiDyFVeo0ZdDznQ4MXWylchQnd6O6cCIoICwPEQ4aCf/F
Px9t3Pm9f9pof+uKOVbsLIJjJTk31uJljazc+5gPXGEHPhsYTH7TfKO8qjH4GPgVvG9cUfsXvBp9
xYtRiTQjaDDHWIDpDRarVighx+Z4ULlQm+o/xIW8c9Df61qybPLf7cy+6gAbaiDRKaxwIjNfXSb+
agURNz9zytSSM0jvVXdrQqzYE3J07eVAKViwRPeLb4YmGiuOvz6GhoaVcmOW+hop7YGbyQyLuMRF
eVS59cH1souG9qvp6Ht53eD9tHiCVnBk1MqS/TQ7OmqcAnFTzKlaHPxHsgRAN0yo4us0wLleItud
y9KZsHF4fZwpwUYS0Y0ioUZUgNURYSq8f7Kgp6aQU34cou385o0T8vqWu5l/pNARmR+ZeKH9T+57
Jr8djHYcNz5D2TcGTIebVcq6pB6WqfvtPUTkeWJxoCELC/X2IaIqNZwJ+kytVM8tJO4JVhIjg1lX
teaA1w/qnwuEvJFEWQvhBs7F15zwzOHoQnDG63DL9/7eYchKR8wF9PRKrzLUT03HkEzIfq1u8Ge1
wl+AJjsZabTLCDDTiL1U77X24m4w2OeiMnppnu5oK39m/Qd5mc8ODwiV7ORRnMk18rCeZa0PUaOw
36rE3vzs/SQ1wwy4aqb9Gh+tacTv/1LbR/3HgH/STAeDKoqeloUuOJTJkgfhR1gdomxURBdHrnII
FcLsTMRi4zYUfHI4YbyJAzdkN4H6PSoLTzLeh/M8NkIoVHYnjHVT3fVenwgLpf/qaV4mScnA4NqP
bWvfTi3oNt+u2/7zJIglR2wffkpzzUwAks4kbX1I1jKVOvQUhWdeVvlrGa0W+VvP3yiHo2p8OOZR
wTTuLtcc07+/bLQluMhDCEMA1NhdRJIVK2adspzCGCmUUPZQ7JCiSfSIdBgRSIP6+J+KbXi3pP4P
bdWTAGy5AWQz+DZ863TcK8DjJdo9/s8OU14Tj+Y0yZLMepuOKwm+fTp4jVfSkiRSFscA2i9J8/GI
3w5uJ4ToZG/wVchNIX0vPNApFZD2auY3tq8HtZPufhAHIl5HUUXBLYOG3MjfbGF+mPZnNKf7DsTL
a0v3xKw92z3/FuKNjTBXuT5TwxJBx2DvhKwPX9PAYJ5s7HKWRBOpef/MKh7XgjchCskDdg8PVjhQ
LMOPPusOBPEZtgGOT136VhQxSZYYFT19885QB+Vz/EyomGi1L8iO7fFqWaIAJlOMi7ypvxofOJ7X
CFauL5U0dfaMFXn2zUg//NMCDdQPHX68iArE6SNbJ1grHkP3lhbgG98OmMPGPjg3iP4x41OeJXno
uk60hF3hWaSSHmElxHBFR077Ih2zqB6FdTQL+IdkXk1dmuPFQprWlT18NNoyg96yDFgGAntPXet4
yoZfcZQT0cqo2XuEswLqk+KQvn5Ey3dszUJ2sb9o1OD4ucBvP1ZL2jwMDBYkzaPrjxLAkcg/axlq
Ldoe6ZRto8NCukhiPn+qucJF8XB+uk7Ykb4ghA6IEZwbud+R5B9WeU34REYbS5ArKI6F9UrTv+LJ
Nl+ZYAwA/GHydRFM3VDreXnWHUvkRh6RhP73k65G8i8xu00amTme0KwhPHibxO3WOsUufi2Fsf/w
A9Xg2GYYeMICRIyhnNbbGV76uBc4ccqWTIWm/Kbr1xXo/Bx+qh6zJp5EZv44ndKO4EzZgModHCuk
b8RqtrUtGhuZv2ToaWMXRBWGySucGE1CByrBl0Vx+Ep1rWLRjT+nkzWoqvO54qqw7Dlq6XqMVxdL
+Gazj9MkBmT9wihxKiJ7vZgynVM6YE7rowxJ+4x6+Ri+tFWThQf59tnQPc5rV4fqKv9BQ25n2EBL
MKfXaNRD6RbJCyu6HpiWH+bZBXVlXlpBHgMX5T9tXfsY+FpdFpfU1QeiTZQGKfzudrBlyGyml3pl
Xw/DnPWk6VlI7DMvDyFuLXRd6l/4IuEoLVTEwBoiFbM5cuIMki3ZJg2zmaeVzxT/Fo5W1uJUanw1
A4kc3tKh1t3oXTNqwMq0X6PadHy7rBHaIANWA0iY/3Tuz/PdKLLNYmZ2dEOf+P4oeh4HRsnFzPaO
j+9j3iRxcYI5eTUHLkCuwyX+LJr/EUTNjnf3y/8ZvwoJ0JYZbBgoJvqmwpEv2yc0ECsUq3WzEAHs
IIZck5w4Wks7cwKSdVoDf6NVhWRtx/cNA+EB4WDV4XXmOtY66iTRLqeg4SNO4+YN7vr2l4OlcwtF
Sxof+7TD2JSaSiASdWJ+9Gj4nEjyjffTU4UllZHCSygebCMJsqbwBDJToMyAGxieWJdCmNd6PKX/
OOjfYvPv2ypLVl1Wu7zHQcEMGhtBPLW6sfWI6N7zQKhLGShnYigGZXiWkcwdhqmCXizvQ0kl4jBJ
sEdcud9LnDiWCFGB+gmTt/XWSlXtumaOY0kjqYyDJ4JoKV/4+nSiam8uqiN9+pDNNMDn7pcqMpm2
6sLF/V2WmxYBDjMfiEVr8zB0Ka2FiSh4iLcczWRtHP+UyTu++dwkI0ZoHp7l43GlKGc34hD/Qhzj
0QCjIbklu1rKXv3w6FP8JRaq+2QaekIY1TG6vcIe59WjrXZoodLFhq1LK9tDytto35C/2vPdGE4M
AFB42PsZVQZSIhJ5J0ctoXqYEAHNS42n1NS6TcUB+664t6UA0L3Xf6IGr57kxPshxYCi6eUa1ELL
jA7gpPaNR2kWygBd4C5t+Dc3PrIGS1C+EEyuIaoltVimwyllsUN3PpIJdjwJmLR9tMAtnul0sEj2
cib32PI6XqAySu2RKEeiJ4PpuGFCGhwzzvlLR52QEMR1kTo19Jg6EZWJ129SxETdFHpAI0gO1d/s
agpom3XYaRjt7maxOKRbUU3hELIzXUl8Y085i5G3ICJbzN5upvOPV9Mh8El9lT1Beh8J8XtiGixM
m8NSKAcu6QVXArJ21RTSGILA/oKPGc2aree6XxihNJgC/sAxmggUknCm+8RKTKOKU0yxvq44eXmK
i8cmdkrLyDULsxwVdsN7qtvctsIgc/PjoM8hDqx6X7L0jA9tuCpJV1UdWGwGpFdDEPsgcqIROb84
Yt+EHZPXnoLWuEZ/y9iWKf4oJpHUtsQi2+5xv19vCrDAJmdT8irzp5fzQ6OICKkZGlgp8rtduaTb
hyJ2sFFd/PBG08MVejtuQDE8qrCYMniDoBDX0kcSyRuCGMksmZmn6QlfYwBI3XajTq4Grrswk32p
YAZWgjPv9qRcUmuqIhqv8hsiROGlWMG2wtRG9pyi3sYBE3JXQF6qplzd3ofc7UWX31msGtlkeH8Y
AFooQJJl7fnzZ5ZYgax3sT2ftR0iKQVAZGnW/JrRrs1fwtXSjup2XGgf0hRqpvf65PJ0FS1a1km1
HoKm3q5AmvUbJc1QDv7htsmoKEXYLuH/JZt99JesGgaOL6dgh3n/66fsDy9bBaxFT0VusglMC0iY
oJoyy/+sA9ZVId/JDsy59tiJesJpf24+2X6yKHndZ9+/qnvcCKCoSYoiA8XOikgKyUCt0H1ysTQG
tY2ICg1xybxvprKroEBolBrKTvU/IdHfu09Sj1nkEPJ8Yhs8F3tM6hZPSsQhBSSFtZiul4rRGDI+
l/3mShSq7r2YEEwdu5bRJNcWvy2AZm1BjBdu1QczoEOXNuYUPkinOS+l4o2NgRN0vxKtLZfQe02J
LPNLol9pvNSToBr/LlJ0RKobJDts1I7J8ptt36VgPEpLLpkHzW39Wvp66aUy6IBN7VNe+YPfHb6b
FuSMbchbZCJ0g2ijQmVAAppoDooNHIkM3rYb1BAurKl1TwzI3oWwrLTt2gLEkMwnnLTN8j8Q9D0t
c8qYLwKrjLY25hy+o7oJd1MfflVkvEfSWZCJ9Cbm8GLxaP8Vk8A31sZidlR9O7DOBP7Qm9uoM9AK
jSd2qn9yCF05m3L8avitPdrh1kkj7v4dCaKDMkcqCJKZJbL4YmZHoV/j649W/aw0v9vrWJJgoF4w
Yqa2TdOrob87rK6s2zSTa4ICXldE7vCf1zadA2WO69g4uzerC6EZ/Osc00l8TZXL/wSWej9F3ZmF
r9LNKgrNTzyZHwjLV4QS+ywy89tMzy4XwNUWu6sWKtxEP+pZNiWDUnLEdFlkhGT8r+XpbI2UyZiM
c4i0NJSLA0lygC9lN4rma7Xw6g0h0k6hLFw5opt4VxnG2txLKkxWWE3JJz8qMVkFyD7GeVEYhVFS
gIfAahbb6L3u9U7n5faL/Pd/BRSai/XwiHhvzfcyzZ+ZmPgrBtOHPDBv+i/xVpwSmVXlzS/3EBw2
BV+w9prGIwccrdx4xM9WuG1UHr4V+IIZl4jb+DbIPySkiGLBy7laWuMAtkoGjSRDj6g+eyml4wyi
1XiZzjay8Hdt80XcFEuazC3mzTDSujiPCYyh7XGBqStOBjgnfwHguO2I90HNSCRL9shHcSbrY2Iv
8DWtxGuEtdW64mG8Q5NazM289wurXrALJ5/JoqQeu9UcqzD3dpHit2qgl0f1i+4SmcyIQHF/9L3B
rB6OYstPHIestBCFBxkgFFfgtlC85lGr47kg11yDfSTEr1VlsLSaImvnjDnlvpTytFeJGtUBi7rB
JMl3pjeq2wi0p2FCF50w7stL2LNG9Wi1TnWHQjCJbClQChp0ZIzvC7sWYbH3tUE92cRNi6n4brhs
gssa+Y+jqhlG1wpty1U+jvoioNF/N+1k6qg7312SFsAxiECleGWM8gYABA70wDcvGAhbOQUTudjU
JYfADBFLMyR7wI7EzTDupvJIaamXZ44qM6gDayX/lclTCdh5JAiir3Zmzy9pFvGgvbK2UEFWHjWU
t8jbgqeHCq65avDYcNQVzqICsq47oGdZ4rCMJmUqEAKUCcG1SaDlM4da/dj/v2OTsWkAhmcQ02Hl
TuFS5+T+a2PzznwtQZzODdCs7GhsZD0DjTjuglGtDCAnuyaSxXR7OajFMZMVUsMsgQ+ae9TWhGwR
Sbs2R+WTEsetCOn7YNCTz9dUUB6bvS5T6YLDwiYKJkKGw7gvqeaRasgJCo3AComMLMhx7qLn9T0t
GUuoIIIlMY3M4IEdqU/+AbEO8L5LbluLpG+TZphWR94+TosOXtDuig3TXq26AxaUD/o8l1sOXHN1
qpbC4ikXxiBsaGN33fu6Hp9UrwlNrbuoRht+7omQf35asd+0MZl78RGZ3xee1A5bSjE/rvgxyrax
C4S3rz9wnh7tLE/Q7Wde4sP3BrbGVnijyU2gQX5t+WvSOzWP0rhT/XQAKnP2Xxl78oIQjOpdX/h7
O5z5OpPOecQ3FlETLqM7Gw97PZraZaVZN3fl2ehmOejylbugdmnaL9qnrZaXEVHtiRzMvHnloaR1
pg5kE/GS7D4+shJTEmrRiJkn/MnyYxrbCatdCp/rvPJzhLzfXWYLwxvaMXWgCJe+xNnlqTOUP5+s
RkQ2XFnOnN5OMS/I4ltlqZdkdYirbZ9w/+1AzGpHyq8QT0p5vbFEW/zmVwxh5F3263Fo/5VWfWfw
GgiBsaqh/Q94FLWlov1ffyNQ1lpFa4xnazsfvcUzbVEv/c5IfmR9aosIE7LkasJhohvz7WFL5jCo
8JY9Pk0QjNtQXCkN3/CQzWR/rwbJlx8r2FkI2LnShCzcCjQd4d66IoxY2DKByrbVgI3V0HsHFVYq
L/KCET6qNjCW3QWxQRshm1Prz9+GQPWuskPDB4UISyvZl4NUyNN9rNqyWporUtwnaBRCvUvpDtI9
0BKA4SFauU+dbgGrr6DqHG6G4J06lPhZ4o3W2hZPt6nZ558X7iaVqOwwNKMrTO+uEOrFFKjUUlDG
JxWsEasU2i1DmMWKkjUSzr/Q8wz+UaEP7t4FlqurmT3djG5RiuPOdhxMQ5eJm/7op7EIQg4XNGN1
8Y9x/MUf6WgkreuSKebyUHGMCRkjn3Fg/Z4rLve4TgHoLnZjbfpYhBB10w4tuJT2jNd7Vi+sA18W
RwJ6BpSeBX2lpaIe/1guE2NMHMAUzr+crded/8po1hidizG8yK4AGLfmn7RZ7sBDyQLOp60Y/wZF
VCa+r0Qa2iKzKOeXV9wv0fZY1IkwKzYroiqXvivVGWC5pm0zwW6p2UWh+Y6GiglcwuMwatIpBUtd
fG1tyHkYB1rmllNmK9m5dt2v5GUBuZQdXZrtplskHvrWeCBsKV4K3YjIOJZv8q/BDe8OpAg9CcxV
lgH4BDCNRDIDWvM2mT22uQZGV1nCvbUMd2uHQUbCJx0Hc2XgKaJxP4AbbEFrd0rZ4eO/KV8uvsa4
4K1sMhL67JDEWMEJwLoeMgIGv0DhNpAuj5vlg18lOsHoUMSia9ibisGIqW/AbH6fDlw2k8L9iPnK
lC6q/OXCSF6a+42pVMSenbGlmVwVIk9XwIpbtLwqD9GjFPEytfasQcK6BAI2GtbdjVSjSLawrCYI
mntBh6DsdYidvcJz4Dt7MZsqWjAYu5UjBTjTV+XcqLREDH0iT0LCu+wcEnCsEfbTXmSSjm8IL8f3
8ZFOXVuBHPye2NNSzR3151rve9Ejd6Zes+g+F+FPIXB+E02teBRpsZTg9pPUEMya46vh2gM/3Y/G
5pRj3QoP8PpY+QP1sUMcw1y3RQY1zzokr1u3BzqLi2ODmrkz0y7bDt5NbufUD4eGqket8GNH1rs9
uy00mthpvRDdkVly8212rfKNpaLWd7yFHK29Q5fbFFc3GtI8MyVyPS93beLmjbJHIDwzkmbHMdVv
/EJ8fm8MrKnH1K2OiLD8s72rrq/Pu43Ewd3tiC48Rg9KjxXdhyshxTwe/N6Im0BNFFinWp+WX903
KcpoUqxJq+3VPuyc+GOIrk9kDEIexZMfFvgtpwFb52mi1qn/CsPO2MsvLglsP9bV56l9RyOEeWA2
PUz0YCHIqQvJHUTaUttIO2M8puSm926xj6HaLxkjCEkEujKOMSiwSW0pOUFQMInqynO5ThIXZxSg
3Rkz6FbEZ5i9GQANAavhddpsQ98UreqfYyY1Lw32HJ/W+lMcFSL4XsL8N7cyVTYyPhc5sJAfRT8m
t+tVnUQoVziPwKU7/M7j24OO0KAmo2aybRLwxvLuJXa8MQI3jeCBx3j77B9aG7PW/TM/DXS0qxkN
yfS1xRBF5Ok9VTXgC8uX8PfIg58tw7GRaJLMv1yCZvwU7XnNJV7/7s+HASUnSJyXVB1QZlCg9xak
nYcmXkWO6zRRLuADeaZ4ZkBq+pJ4c4s8CTsNa71HO5YU5wI3hXWLHWyLlQzS0urfJkWi0yWPlDFE
u8AfiJEOKscK9EYiuL2SBoD02f3jsTluTC7IvMg56bzrWIjtNYddngbDA4kOe3ZGvDfYgeF15Erj
/giCfwBH01ZKHk7JLW5y1Rfll/T8rDyjWEKmFRB49s13rZgHJquNKvjly6h4XlesQRRWRWn/pYdj
+c9o0dRht9Xf8w68LHw/cJtOpQlnU29uSIQVAxIj7Cv93pv5/8wHX/9qzX+caqv6DLKbQhTKdY78
rzzNS2UjCTaIgT76cHef7H6u7P5DDwlaCjdFmL+s/upKpkMyEjsMI2Xp+diCGiW7lPkvfD+b1d8L
UjkMcm24zKZLAvS6wLc/wUwKvY8LYkIX9PjI1P1zuJHGfdB366eYvsWKEuzYVCcU5LOhW4jodshN
y68Km5yEktEFQO3NvSlyfPN8o1aovJzJHZ94ECJ5QjphrmJnMqO5sscsCfTF89KxuVsC6KafeZm8
KglakMLQqgUbJLLw/KiagcIsG5kZH/ODcM1Zz09BodtC8WUz0hrocmvDm2ZitVj7t4dLD7GCctXg
sV86PCSw8FS9oER+5xCdR+DdwTbpqpIpXNC6yPCPXbKDbNPtPKeeDaOFC8F9xgZ7J3bSmKTq108Y
jf3tBha9uoE7CBDkhT9zTHHVfdXpgv8KJCfnqw8g6R0vuQiiUyiW1E+Huz3GqNowBRRilL4S+LvM
PPiAybyiJjC3uyW2JA74ic5XKGnD/34WSXXpqBc9Nn8pCrV/4FKeUcxE+GtG2QSJTWrQ4JbEhMD8
3FYTsvNiPKqpvHShlWNXP9lfzeNln6JBVTFQgR/zqjLqYlSBz+gQxtagbZ+L7mJp1qZ6Wrv/DvFI
QsYDCRM+sK3c7viU+E5eYlpNvO3t3syQLAgYn83Kf9+mJcLoGLwWxPc8TepijHYzh1YriJYqjrmA
GyhFBVG24iyIF1lWN5kmy9V0n2BtzUPqDQvF78ipv5XK7T5/NQXNOClpqdYNxe3dn48tZ8r5THl2
8hEMx2e7vHT47EjwFpQkSc0C3E+9xaXVEQYak329xMoZLEaZeZmS+ejuBYF45mDjHd2M0ouD2tIU
v12EbtlLirXnH8IFUpXSko10wyn2mqoOprh3cXiMxnztJDv6SR6DqbpVx88T1SBqrMPJ+NnpWhCM
xBOBT+idfqHVSC9P+HGKOaNqsoExRonxSecoDxGN1Rh6Mx3n0e+2LIJOhrDOEfvWagIEZHYRRdtZ
3A11y89efiH8hKaEEoHtxhY2sjPhsyWGvSumJWh03ZySvBF5mU0lqKefNpwuQ0o+I66/3IZxgHOz
DSEtk0s/hJroH8l9OfQpGLbGowOdTdo/LCOcyiGWvLvHS1d3r9Bzuqn7kk6EU7LUIINK1BkPhump
KunU+c9FuLIsJGcOY+Q0rJO9zclOZgwcJAazAKoScf6ojihChVw2QYqURWZya6j63oooLN8yeT3G
sZvw3xcCm7feJj9UzA+rLPspj2hI8myId8Qb5Y3aotJVaupYV6jW46aGWPTfZ8tGZDIdy9037CMn
aPlEHkypgWzfSDE/+96ZrAxkAlmZL7x3MV2Tql+psMeAVFMZDX0GLN0A4zPvOYsCWIb5Wl3kmy/r
cbMqQEbmn07wQAVe0PNWhHUJtCCBoEEF4DD6y0Y8CTCu9hOSY9DKnVnN5Aut0RGYy1/GXoY7er9P
qKwF10odgNV27WzOZFKVFFRlg8UJDAYzfjjXrL/xqjQRF/uo74nrpLULCk5aXXthKJ4xPAK3IiMp
cdr1qk5Ms/FDn8ONapv7KSOkKBQ2fUEe8TP2lYXPoClBM30cSIC8YdYv8rFahLNMtbQJdnxfFLqZ
GkQ8WdTquROyNWpJmZAG4fiat6wHNB/QDYHcjZlNk8zflwJumq9umsP67pevua3YsQcr7xm2y5Gz
v4+MsHd5MDeSYFCfEepSLe7g2vuctTQy5nHf7HrindLzwRLOKMVJ5TByX9KZDcw4smXgWZu+V8je
MBBsaPT8k9L5EgT77M6vnk+7acilA8G0hznxaYLoYmYv6GYxENkQReXu7hLrqRvuasgeQ4HmPPC5
qqJ+qn7VpSDRiSHQ0OAg4x9GyAzC24sIsBrSIriF1q7hFlJ9Lx9RfW7kBCrd4ZfEkCpSz27HaBZs
TMGaI8/Gfff93A8uhyZNZgqJ6Sm2Ad44cNS4k+jIiL2GWwzu4iF7gzvXFi6P6YiIDn1HUEFDzJhF
zs0Q9QSB4c+LVZ6L+JsJOjpSTPSG1vYiRsgJUHaFMEumGJ70e7DJAcH8oYzem43ZCsiJKjEucCFR
6wqF54rSZAVFJovsCUKrK+CppeN9wJ017GQGh+XruS/8lb62+y40D37XHIoOb0ccC4Yb1JzS7vI9
mORQ1yEN8svLVae24v3YPMD/TJnplbImEgDSx3LpPua6c7JZAQnkveLHP9k3ftAOPtzd118CGbnL
rYZHA948GQ4+UN+FbFHxWA6YsP4DNvQQWPzW56dthIQantYfztwmUWSiPPzajgttmDr5G/fHZ+qG
edLM+CC4Mg5pYXF90OBibcl5ZaByfj3Y95RPFufPP0TW4sZh0LR0DXl4iwhlYaadJa1lsbEpA+SC
pm06DxH+kN81oVpxBBLPQFKc9KSdBtNjaa/SGDoy9EUdcXcukQXcX5qC8FMmo/s3clzYRgpH4mky
U8A1FfeZk0UuQer4w34ZJq0rHL/7VDlUZtYmIPTtuxGL0tRdIRCdCasC91LfsrAOv5QM+3MpwE8Q
ZeBxmdv3IIbFJ/9DlyH+4EZSMvZEK2Qzj2Uxaj7ljWD7auhiQay9S6eWIjCPy3T70jVXQDj10NBR
okNtjsR7HLDL/gxs9ybsIWlhMbos/3YSo7ya6I5QeqZL0RpjfJO62P0P2+S5wnaYv9NHSbsP49YA
KHpiQ4bF86K+kYUlIyEzYSPbNl1JgK8BEUAfJrob0oXLcWzvwkrUYLpmtP18WqWP2jl4MpOUgtwT
XSv2dQRLiZLqQa+THLrC7EDm4NxlhFXNd2mh20fA9yBvh3ewPSNm8J2Blqd3l1RGoqIgHQgfmQva
IPRsRZoDRaCOJXLC5K9UG+d3zlvhSmSvymJQAd+8JkLcwYnFtNDYkvC/zs8P2ache/C96SbtNzA1
MrWJZlpX6ecW2LUULRVnYoIk4FCsKtlmXQA/RomAgZ4OmvMIb9xBJJBqIaR2uYvJQom+9fCBAjNh
jKuPDT/nFH5la+TN5Ow9+Ts9vJFdCoNuyyBx7Aw5LIBR2f/zAsep0/ff4XAmR/3ixmsuvRa+rlH7
M7a+oFEchO99bI3BOyD+tJI7lyjMLlAqXW9gJXqg8bvLoJDlXbIt68mj1VNdrll1pEai/i4uVJqg
zQJM2OuVICC5FUyzD10HcEClgoMBTHN3GIpgt27M8vQYtwNiQpPJA/J2rXa7l5WrOmCQowyfJHHI
XZslMomssfgcFBRl4hhwPAY37HkdjSmhl/Ca5B7hBhHnae1ZOyT/GlGRuxLthDk7Ql8xySuppJA/
a8YR9XeQaN2TIa41g7EOrfQVDyjs8dXUW1+ONEzus1TkHPWq+C4Z2vLE5Ptktx3I64pkrkQERJAr
A92D0Ma/vPIS8sgooWI4c2SQwpXu8Sj6hEvTIVKwYjfZbPS2X9R1BySmh92bfLgLvAImCeG4ETj3
coHdGMgTaLHJkrFGYnB+LpHkA/Mr73Z7aOEb7fwvaAJN+P9SPnP6/SPJUJmDwUZ22aYXX4zqrDK6
2m+z0IB1Cn9qLGQCce8NKeKLe2Np2WA+b9IzYXyWacSZt9dC5u1yl6AAzVZhoE1VXlgXsH60GHx8
oIbzUQ1KRDgEClGzWOwO/Qa5QdaB5VBPFj+9f2A6nF4+Gs5a/dGTfKb5bPJov2lUNEQE62oUzvtL
uOrFipI1Mi7ouLI977KbaWkhqM/rLP7leu40zq9SUutelvzGgKh3/XSyIbQJl3LEr5MwvaTVG+r2
/RFS717OsH6prxgiTZ3oCDhfrHotm/nzzKzdhCrx/WT8D/HwULcg37md82S4euvR24NxwLW2vb8Y
dmgp6XtZYeIHsUSCWbz2OJpcu4UfRJNwC5zDNwqgbuWUiB8KKWAaftY0zXjfKrJrwYdUr7274iyf
gKFcR3QN/LqwQFrAeAgbI97PgBwCragk0+iAdWtd9J6JGHaqCuSmM9+3MYNl6kbFLK+VMsN0t0TH
7hLgtAOwenwrJAb7+dym/qA9ks9kt1WLFngjKnD+hM1a8QCH5KybVnsb+p7iDAFI89Z8i3/jEM4Z
3tX7LIHIlrzjgGe+5y221RfYEV036RlS+M9r/VPJYLjb5DG7jla7lKU6eGLcsIw8TDeBmHzRZ/DQ
jNk89/1JjmDLm6OBby6C5toD0k7rmE1o7Vf3P3n9Gw6jHfAgu8eV4sBriV4OCbTh3xe1H19YSuwp
GzuhT/eW+DP1aaSaFG81DFAsVAffki38OS9N20OQqCzNTZRF5YEmxmOTmIV0OGziUYgkj/cmsIFc
uARK3knLWa+qU7a9k8iXkVcHkfjbm7wkTshuoXdfP3w4soDrsVFGn63NSZmIbQWoLiSNrWxhCQek
47OwwZkNhtj7AoM+HENU+eRGmWFZG5AKvLVb0/wSX9wleEoWkQYyYLEraHy5hXdn06TIHNO6Nj3j
oWOj9D2yLm6oa/Dp5vCh27oXRNTjX7Qbr7CS08OOyJB8Cm2wm4EBfUR+kWxGNvtVkMvxAwZG9gb9
CYg5saSvdTs1KcpHQAa+EcURV1AExYKsv27SR+88Bxbjy69+sT4my2UWlqItvgbBFoEDP2paG3wY
2Iw+2NKiGk48XJ6cmO8SHvjtZ7F2c1j/Eev0ZrvE5aigYcJiK+1kWJC58r8QPa7iVL20ltMY0yGH
77L2LByawBKmnKyThUsRr/7PUhnaxEn0xzhWkq+Ha66sDCCjXKM/LmdCpMtUt3HCn4rm5iHtXQDP
NmvyULUcf8kleb4dBmSkPt564G9CrcqewaDgliTTTL6+Xm96GVSaupw26UM43Qv12N/NXYwUYB7z
ryD1/M9xjGag3OduFQEWCpddOk0C2cfWoGbFQdI3DlXQPp3qA4kFOjNNK076KEhUvIUWAff2DkUF
Qw5uaxTGVW6yghJjMK2LAL7tNucSFwprQ2kfzFTdqM/02Nc4q/Oh8BmZITksRnNxxaw7pGGWZuvi
DQ0AOf+A+zwuPEn4spP36XWmqYUoBVPQB9PWPbifJImQ1d1srNsOx/pCbrhuyj9gf4OlpCUKl8os
lQ7+0FEa9GB3c1zpp4flxXYR1jMOUVHR095RZgpCrjJG2NMlF/9AAuvy4eqTGihXDMApIuN6xRMW
qy8YB4gzK6v+zRrt3U8DypHdOLIvMYWFPr9gSPDIPTawo095F3CgwDIegkWifxf2TQZlQUlkFJ3k
XE8tFysoALlcsKFxg0t76SKd20MiyCEroOdSw6KYSGI6Vvg5Bt6tFUARVsmgAR61lAhSPBX87jtN
gHL55Aw3WyMStMGX2J+5FUWULOgzYNAz0O7XzpUP/qP7Q8yV2yi+AO6p4QWKKnfaTb4c8vtyAygR
+KWQvenNpGwx7FQQ4S/tv1bSv8nekQv7hooG05F8ufzPz6da03fxzG67NwjmS0+OzbZ/b0O7nxUF
NSu7KHGuN7cDIR/Z7qkZYUgJiDp0lZSGPNW+BLQEDLgqAlNE1IdREqUH0tZ3DyIVLsOO5dtwuZOU
b5bGI6R6h1dOERMFhv92OymI1Wsf5uDsSUCp4nEaWCaU+W/ikgyyUfxB6d7uMew0a9zNskRacn9Z
ksmRVH0aHyF0G/dY5deHrCJw0K5KcUsfP7Jd6fK5ZtuSH/DkNHPL6Hh6aYeEqgHxFIB+Mk0OHWv/
+jB8QeCjI3AEQ3jPlPvKX8R4giAGaFO1BpggqNqBTcZTN8w+G2fqQyM/oBz3VBqSJO5XUwNV3i7A
DJm4JNS1Nu9vYlSbi5Foy2eJ7my1wCuNhDSHAN0LcC3p37aDoQkrBguvzS1JPxU+rQfBHZ4vf4a3
Q43flt953Yl+qGoAw0GTXbfJovcEBT+84y+p13k9MWjOHcTiiB42qjRIPK0mLMsKPXIUazFsp2wP
EL9jOD2rKKmrszeg9MkBflzhKtaP1LZ69AYSjKN62D0bndTmEl05rBmcOCUoG4T+niSjIbacZXBl
7i2dO8wpENYcKs04ASbT513ZRy+CrLvPs+yP8zeJPYUE3GZSFnCv8kM4VCMuEBTgBXcceYz5Nx0y
E/tHqb4beXdsb7+7b9V1udeINq9/+YFzXUa8VPflJHafFzRG6Qr+Dg/jpfnb76oyidz1N8saqcOj
5nfj/50J9rYCZupEMjmGS4CbtylBvfRR/0K17h6ysMjSjk0RDOJ5Xs/u3NdmbTsc9MRjAVNbUdYN
uabxBzooMuR1PfunXkJG6mccGnRQRI5LXd/shSqhpJr1Aq14mCfwkltWquT4964EfbryLXXQSNUU
7mLz3kP4Lw8fU1ovWMcmjzZWyNBe+h15aGCR3NXQx1e7oRyPmCdmhU9AYtQXHqrW9/B0+2FD7FTP
8RCZpYG42kp0qo0Voxhc/LyFCfiqE68R0yLIvLjkM/ccLTMTtIGZ9Cr4f4/Kma3L0oKjZP3GARpr
HD5sRBhq9tOuK+isTcc7u55E5+OJEsSwbiuwq0x5p+7aCmhIKJ5omYvmzjcA1G0LNVlQIxix/jYq
p8UcnWCxpZPjzJchW/oSGRmWteB5SApqDXcbzI120tzhlQnn9WuVZth9/xkoUO/6OLCSScmESiIn
NxO9iZY2VRJTgAXQQWJLTg9hn/lLdEMllsQrnpYinnOk6+23BlMNTmCd0x/qsYh207njWiEcuZjT
UY2jPWW/AQDB5RK8PcbKY8gg3shCSKCRoJYAUG1ifOvM7vjdepWKh3mGRcs4Wgy5EzHAZ9Xea8zu
fBobYM919vtsa3vD2lVApGDtCAAX/jw4wvzZ2CalxueMo08akZpz7WkGPHt2zHoyl7jizbVgpSsf
0trrheMklEh6t52D6F4rpxbB1LQAGKbq1t8Nlw6WKUsiGZOYPHCflymMCvchNaybXJkrtP4Q1GUI
185t2zvixhMaY+tqKCyR/cV3Plf7W5y3veLtGy4zD/lxZ16ecJcHDD0KWhWJy0jjuotinl9sUrRO
h+HaagEDFxiHrRT2WFUB8/5Z6wKhIwsr3dLD6JCaDz1FWoz7m22A87Zm2FuvGfkwoIrYelDD/laL
YSMzZt3OE1LMETzJV4fx9CLuZobzYJs5j3oaSs0GZgWYwDFfMlpa/6MQlGmSrfjknjHH1L7c0xs8
6RzSWdImcrmBt8miQ/FOhoNMJchoC8aIMarnh6uCvdzq7eubXb+VwmDYVOS11yaxPTk/3sk5udkK
a9EEyZ+TJU4cvGoePym6hhjJM836FDbHbr/WoQ06oa5WHjklj/aZI7IwPDq8XgYHkBJO7n2UIXoJ
hA3l/Hzi/AMa9vpG5f6iMEKFQvysZstL26GY8HXfWmHg+iKLwMPaGJ3Xk+Y7miCFppAN4Wc/vkYZ
hW7LqNYj1OHyHrfA7sB/ZQ/70Tl77f3+BTUCdy8lg4QM8AAIdLGEivD/Dr471Q8YZPcYe7ytjbLj
tlyQlSeK5vMquEdnLyzviNK9Szq7Uyiu7gW2vAWD+sazIMgNuRInQFtZHiqlV5RWI0ASZVSXKItg
01ubnTfBP0XIGvjFcrohuGmJdQVrLrXcDmyVTKc5rC5bBRsUfl8wXR+7Cta2aaHKozRG/7+RusZf
cUGAjwNYmszMDrw9VZ9ZFNHbkatd4yS3kU8qMEsEil5+43FifCKLBWqoujfK/IfGJerIfEtvv24n
0RYU1SrGS6ej+j60Kx9QYMpO1p2Clc38UF/mFs9wdTxJ3VE5Ic883/qfpagtu+qLLiy+9P6VhG8G
4ydBVvWuXBkpMUE8mgA4w7DKzaxgFjfjZOHhcJzjPxTAKr6x7PVU7j50mdGbtceJINy/7adGQjP+
3Ecmfn01teb/DpDwlgH3PqNwnAIAw5bm6swz1mfrn1t1NEPuOOnnwkXQ7GOEnIfK1agQNo7cXHiy
osXxLXjhhcKpx154n3DpYWX3hBqISgcZhqk/RZPNhdF6DJ5vRWnv+fIGFP6U8Uor49LrE/aruRUx
IoaMrYZaNB33qjWZwuc8mg2PArX+3bTWV7NdQ65FtQsNYTxLSFd4Lx4wndLjpbnEkv1NRQo6URfF
JXplmON4U2Ehoj8j88WSl5aYzufxo3N4vHnNO/TNn1M8lE+LKQQv7Pl7oSJoatwtOEPEzn7frJtr
4QFYVxM7VJREEbgQ/GP55Os2n0m9fL+vQYypYK+3TDs/3/Qf4h94S5ShcLY9IH/LiARRVAgrOs4k
JGpQ7V+wjIe2R8Knv5oNAF0xRKH26rBBI0J5I5r6j8lVCz98LntJA7BWGsyk2vTEMU8JHMToKxhC
v+S4x9p7zxkqotcsB2QFX8Em9XyzGQ3fKF/mZezZS3QefY2C1m0x5K8zpChaaK3qVzzhu8sDhB8Z
59hZq+8D8QkS2VQHfLV9J0hl4PdCUuKspoUDa8RYjaLl85NlUBNM9kJPzVrgu2+IGYDZensFyMw6
+wxK6/D/V0vwuJyjjDOO5UY7eRvshSmfm8gYTTjZukA7mtkyQcMuBqmhBcE6rj8exluioaOmZ2Jq
LmVZX4ZDv+GGLmOGpoBvcmdSIsF2QZonTlJkJOjxTG9+0JnEXD0fPccbqpMIdpoaT6dhWs8/HuCE
BGXGAodPaDr1f0/DjTHAdU63f/t5AXXK2hN45xrOd09/2etcQBxh8Pxiulg9F04BeDi5JWYEPxSh
pkOhZnyxWK7SQEE9ZyEGfJ8QAsGQxK+Ajz0NN0GLE6RyiZ+jJF+zn/Nob6ud98SCjgG0bd7uTELm
7MHcDzUZg2FgaU5WUAFe8ZRK0chKZn9Z0d47g4qiZCumZgJ/+L4T9eUpx/3oawG/W/cRFr0f/2VH
eewVd8N7A+HPWt5YE6b3rg5b7vuoKxvbh2Me7bqSYGUdRSJFTyJC231ngd2ngsf3GagbUrLlwDmR
EzFyvtvtdUicjn6IFcUdoBXe9DQ2OprrdVIOd2gXYXhf6vj6E+UQnzrVP29gXquvn2z20NFznZns
75MB5QgMme7KhSvvrsKY3IhNVmMNxg3ofdGmupRrm3VGgMJHIJD3inOKwWJQKh6rYcakdkx8g5bZ
Emr3tQ8bcIc0GL3BbnyYhEdR7I6HAZvX/dh8AHszT0J1YSeZnLvptINiYuhD0XY3T0wkS6VL3XHN
6KcECknCZQkihPJE/q4JbzOzQx/D1BkVoCMsZFFlS8daBZYV+HFMNg3TqeqFousJD6wuK03QfYqE
EomqFo8Bhm+pRBK1GlhiNH+6KwdZUv+DbjlRiom6sHvnxnX94rvVW0z7uL0j/Db8BXSNZxWrto+N
WRJC4L/Q+/GBQyuo5uZzWmbV5k7bmdSVUYMtr7rjoOd2nBAv8fDJgPPchdec0urCAprbkQjbjVXs
r7EHHVg7kmyLvxm8WZ09SstdzKZdqnK0+ulxY5f2MJevD7rbNtuJUqGVqjc+NxG8+YGKbCrxXQSH
tiMhj1lFk2vTX/IoTyP1qq/oUCrLHsuIQbE3HxY8byLnwYJfi88wb7o/8VAtxSyFAQqn+48UFzmg
iFA8O2FhHBe8Yafpz1xZEDBBSZMCTZwPCpsNRzju/btQOmB9KX1wadnE3yzElPqGmXC/+aqLnruC
EO1VGKn7JdBZu8SJT0y8/MBieQy4q8bSsd0OqnWwxSVyVyahZdm2F0ph8TWoKDXGBNA0m2BWHQUA
RnHSqlOIqgHLao6GtklAeoe/pVABfgB4bD8PJhh353KZ082tz9hSckqanQN/ewwq640AFvoK/MWm
M5lBjQGSFWZmqGb+jlmrGG+zs17P1FTCby4cPfsmhyU5Bv/gVxaC+HRss/JFmAX+RUTVv8GpM90A
Kg0EWrjek/utgs1Upl0Wq8iY2q285QdNSyqBWgiTwjN9ZAujJc7JlN1hAbq60t46LWjSw89lYnXx
rHtkbW0+hcgrq8XvBjdCJK5lvfixhXY6lysPlBfyjck70ntYUUMihJblJP3Be6JCs33YweewK/kg
t1glzafyPoQgSz67YtAsfP/Imv7f5Wi80T+dTISWtvOCak8A/f98tnTvqRSErVMOq9eeM1klj19I
lHGenM4jrcS458hrrpnrwaNZ4MXxlSEkNDyLIfid/pKRwozyqe5oo3EOIxm2Hf2ZCvPN+PyvFmuY
h8A36KOZB1U8laFKV0gN0/dJ4wzxoXM0Kowvy97Ws8xVOIzznRU2Urct3NtSyD2VALYa4rjEpIPJ
iT71iboVoSkfLlWn4AL4spY8I9EXyR8rTz9y5gpFOIhIShhiTHj48E5P6jJAGnu29TKpyb4p00XD
gsRY7y/m2h5fn3gM3w4zomVXQNJQnZX4TefBOh6PY2IRn/ovvswVbf2fxg45Nr1NJ10y7czTdCvr
jGFFU/ryn58A3ZRpvXZqaCQyCNrgeh2Sn8yD0BaljzN0FnNwutqH+S4/LX2dR5GfpFYbQMCWdssv
r5nWS2rIoC7RChEJoSGjMbK998HuVJR8yLS6+LJM8KMlm3/vT+u4+MRL34UM3GVAU/r720pC3N9G
XJrBELk/tuRpHkMn+c4PZyCcup6km2D8yWOc1t9Z0Wir0NxEyWoECSxZ0p5dF5+nb5BGrpTzYKqy
zsjMYI6/ktKqkvFXFcasaPVZaIah8xDIyZHvF8vft+i+tEVY4HmgRkpWqYUOPeoqnIQYqa/suN+k
/v1w2Kkc5vxZcqEZtVfTS1tTgAQXGoN6FElS6xq7vESBNstoV5TjBJadmy3sZbLtvapCrZan+QER
m5mHPlNaizt+Jvc3cSUaRB/uZ3ZpdVhoM15HbTB6Mr091mG9bxWn40OyKxGOUSQvVoiMTYyGuQ/j
hn/21+3Vz36phYRUdBlQMNuZOMdW9ygHl7F0ak1fft6epQ4uHERAhlX4YB8CeXsNV37xWbXKe05Z
KtfpI2w5b2e6pBXiiQg5hINKjvwGnW0F4LxgTdkJIUSMxiAWAHB1dgVSJZA/DIho9InKQ/gYUBRu
Bb9pcmnk4fKOaNQaS4O0Rmrb+aBJggXEdmDdijJyCNg+5JoQJVDcEURMswo5S1p1QxFz/GdmGQ/M
AbxP1ZKwENlexOWSHM9B3k2Xly146makgk1mEynXaFDozK9l3i5lGClBSQ2kxW4/udWHMHgp3hKZ
Jcv0+67b8eHqwVeLk+drCXZ0V/eA2WwnTnKpGoQrYeAjEfDuHN/B6Un97MfhyZO4ygOO563qpn3T
Mk9lvjF46H2iQUaaeNDa7GjrIY0h21lBiaJEp9qsaWbGu1Yqx7fX1AtQSurivAr/fudBuXl4E7zP
EXmWJomyDFIAq4TchKl2RaCbSZhIHNPI7jxbGwAKxwxmLzSAnxQsnpaILIEZRy05x03h39n5lU7l
Y1n5BOorVX+LQLHryaocUDz0rULmsAYXbpV/4r8fhJPFTROIlcm9V+pCCnLLzOo/8BG89vLzAZMO
cd7XH5zrfXzbHY9IWkbHVN3bOMrBe0kV8DqiO0YHTO2ByRfOdqMnZ8fpDLwHZW8zx3uPLng7tmz4
uAQmknjpl0hZw9rLcEr2BPtfVC+JuvrY0su0dMJ8+WC2JoqnZSFsH/cnHMnxYq2VuUxkw74TZpxZ
q9rxlyg10zv/SSLcaCQ+YK2LVAyySzHYC8qE5TMOw9ynh3z8Y6XHpR7CTfDzFrcI15Uf97DN19cs
j2IiECkALNq7rDt6jFZjXa1pEb0AnAh2PnDKYjzpmvete+GmRKV2dcqGL8+0Bg05rMZNk5TPJjUh
SYGcaUpx5REL2tsZy1FYnJldvkUfscjmHwqbiIrROjU3DG0gQIhdPpLBCiCdzDBuyvaQDV1514PN
6qRF8i4i4AH2K/qGHjwiyAK7Ppb+mCy2dzWfRy/eAvl3o5rn2MpqKZgK21/4fokixc4wQQ97iuOd
y0v1AgZMRf9Nx8lKa8NNRhVv3y96iGpkSNM+TmbMS7007iUyZdWFcekJRqodYPSY16FSXI3qQhzf
pBXND84R2xBFAaAD+/ZLAEo/UTzV2VySiVtewYw32Q3tTW8r3fmSdfnG4Kxk1MBhR15WxhdcnKId
fT0FZAezoODq8IKfTlTOu4aEfI1utQYYinEpxZgdANdn4I+kDIq5DWL0QDET9RJOsg1sqjxWiYMZ
dufXhvK940I7CKjgZN5KwzJDYr8odcl1FaVbi3OHdAUyzzGxr8wyplwVHys12OPlb/iot34jM6DZ
5+r/mJksOWcSEVc1cUAYcBTD5oR+/dDtSDt9hjxRcA8TzrzTKNwc8U1/6MQuS6lfPJhY2Yov+Qw3
6uiMQswQYTo9HZ83NY/Lu1ktUU/0KGbYo6H+2D/+zXxhh2b/OY9fnvCcUineV/sYo0kPkzR/PbCE
+59ctDdb5vzkOpaqvTgOWsYTbSbxNulmuFIDhSQW36F6B7s3FskjH2bgVU2h+lxk+WBqSCQzNY5h
s1YF9YDqkBZiOGQqaNGkD2hjmqDj2WXlSsL6ZvIsk8jjNoGH5M9woejSfFOsu7CFbS0oyFBezih7
kbBzdwhmImBRXT1gQ5xgC/nnAHN6ArGOjFfUTOoFZKTM7/KaqgTAwiawdg8N8SmDpfyFDPgNapEQ
8MdFe30wmzEeNxX2Pf98Pa5ecLntY+AaPK5AZLDVAjv0VVsKRBzRC8lse0zcKBTVjUxTQ9nIMmv1
53UjUVupSgBcsOCSkxx+JOKRJcMLEEf7qBdqWUepWsfL3yiNRR13Lb2VwAi3LuErrC1uPmNuPQ8y
4YtnFBQ8650a3yFspL88DBXh39Hts6djSKRbk8oQ7ciuGuAZZ8IKYbeF1heLVwvtVkNMjLaZHd03
P1duHYWKJSVkkf9s28QTUuO7s3XGbJ2lDCsDutcSOZE43SgpIX6JC9F8CDULHhExUdokNOXVfp8X
2BGYnAzaCjetnukfTd9fAZLMBRaY8Z+e5rukAc4+x+Lqc7mBFrUFAVSZVp+lZsS7ADJrPdJWH8Dv
8Ilm6WtG3eWiJNw0LKNoCrh9Iny0+kukUQuBAv0Kf/IhHRfEyuEBIzhiqtEAyPb3B/6QVSi748UK
2tDaow7wEA70XHjLoanKXEuNPF9PFHTpnNN8DGevHyo2Iw9SGui4XA/yPeKZHfsdB93V5UzYwcig
7qAEHyOEmvyelmZNVTUJqXvQHeziF73QDizaei/5jKR3v8sBabnMHIgG1Rb8LRzF4cPtq4pS33Y5
AtEb3Gsk5ohxR4LPq9+8SmoV57F4+ojNL0zSnNEIsFE0itd78Ci2reeoz/Z4legwz561UH6L3hd6
2Cga4zEW56wlWV1AzdYFkIe5OqkSNl994rtODLiMKGaF3ODoh3DTfnmEHpGHoPWmgj7qRhVZmts2
pF6hyHJd0NTxgOIoJqzJkImgXu7746UdmwlGVTZE9yXrTsd+apBd8nvSghYnobfaK8/csixKOnnJ
oMkUMgdw+CHNI+JjLgy7WY/kTEmKres3pAGiuBoTmuiy8iiZz+3AihkPIVDQ36dhPCQItdlHqg6B
sRFkMb6Gse4ifJtBlFLaU7573kNurpP2L287ZWdCpLA8CCHtWkmB2YczhHEvLMFEdoUH9QoKFHIR
3XwNCqafjqfxUtaokTCL7nz/UoH+x+LGXV93n6JYN09VqTOkKo8A//Im8fg9mSZWB3QChscfutl3
av3ip4sPmVSPgyn9Yori5EaeyV6CdjuI2VITvpn3cHSLKRf7S0R6OWRkEoNFFRPNRaySbBdv0Wi9
bRUUNRWD4YAUJTKRzk0BUwbroZXejvWzKi19/nLSZisYEFDsX7cRRBZ8h9OnIXuRtO2lhptco258
to67is/bEk5FSm7rfbHRxqCNgXGx0x6L64BtcUQy3XNvGNgqHBrwaTqCqqgrS3/nlH8ZSoJ+mqH1
24v8elmmY6Dhe/MRCsBP2+ZjP9gs2LsORa05dDO4qiooKBqS+5Um+e1Rr4vi8LswvXLpt9YuYCx/
vcy/2tmDwtXFFij/m4pXWbeAxz7W00HkcLvKhCQ/Qq+NSYxyy9VAYhPIP8BRNsPWPZjUO2pHBQzW
ZzDEJO6G0uZA9BQQbtPUDuxbsMO1o5d0dzZn5x3lio70j90/xQeNvWUohqU4hz+MsZJQVu8h4Drt
qDzYo3JaKoPn5gdAcoVsl431GKwY5KpPRSUj1bdKyAtw1mKk0xje2F8/V7YWPhMLm7G8xyrRp9a1
MSKGgCPYfN3ViNq/6Vw8kD10b9F33cxL/bYjSfX+or16dakLLpLbaLme80TJSNEglX6lchdr4AGM
ue43aByvnIGglDrzoNuQfMLaQHqw0jikaKpbmSqdm1qJh2ljhhtbYpsH/HjvtNTqif9mW2qqlSJh
Kyb2CJlwlTT5reJOXksAtDz7r05g5lgVEjYh4OvIb1Un7gMiQ4BqejxSteqgtQcrK21MK65Wd7RD
rqHwLkSiiJLj0ZRZ990hCi0cLuSoTqdTuXcsMtTXBRNLXOG4YWlbh9SdBceBpqwKzGyVJyKi99L+
KI0Fx0Qm4noQe9ZelVV2Y/RGynwNQQHK29+5SKEUSR7ldjgb9VeJYyiO3KXzl3K0X/8BxFyWhlpa
OLPmAjoDvkBJZttnWH2dT/0L6HQVtQMtUGFMpJSsgXu5ZztwK5PSTKKtkM8eOZ66Tqr7OIdNiwAv
2LcH8E57VRVPubHJKOiYrnR+Wl81mLm3bmXG2pgWEhkswo58Tu5lZNIopwy+LCi29yLQw7JHsA4n
pdfMZrcUid27mihFQ5aoDp5V3+OQ9YDRpE16A7i4tRGr9JgHnwhvU0B6QVkSyvugTTH9IF+YN8mT
zTecU1ezFYbDZx7xPOt1lem7JnPuaYsIg+17KJUcm/xCG//W4KzU/PqbBoINI6nuPZz6bJs/IBBo
foatiLoaGHKwQUG3gPRtmJCIIiRF4H8aMvzW7vDIitZintYsJKM5Z9Waq4Snsx09YbZKG0pKwBDp
04lKbf1AwGnlcaf2Gn58ZZdRPT2ItjXXPYcunduI6ft3GJI6Bu+0P1rSNeiXmSuxujiV2uMQ9Hq0
xoX+Kya6HVkG94tVA/EZdCnrWxSd4HuFmkwoxH6juPuQvMTM7FKrWkFRTxzy/mwzf8drhvS4eD49
93c6j8ZxTKWXufheRwTmrnELQV8jXyu/5OM/TZzytYfELVPhBguQilaLYwDIiLElbqBidc5VTQtO
rxmMCZytTnVgJTGy3So00BpMdHHGvIaAjzafXXznwbfOvGtxsaCqkPHdm2c5NtQdtq80foLTxTnu
TXZ+xwxmvVcT3AWBpVJrAiEBQs6JWesnHsVmcLB8mXsIWLUU2IVXFKXAGw28cKpSAbxHiQfyHXJt
0r+e3iIcXVhfAuCq2U/cYK5czBdJTWq7SkblSIgQc8ciehpJG9XDY7e7BHRO7j7kpHvijiLIOQqg
qQtSIwKoeny8nj2VxYC2fqaZAYaNu2y57KX1ooucF5cwG8kPzymKxAoFivrtSO7TaaKALDDsrY7C
OdzPLZH/ynLclXUojFCEA0rV17Eq5EG2vsBYE1ubBRtjJ/iJLCfTvL02Dyrzr/b2dGNSEnu9ElqY
LrpRqUtrT6EI67Si9gT8evx83/Wa8fPTZKvSJfWLRGS/PvIHOgXSYJJNxyAJoDR4cqFK18bu7Zef
e+YCrt//eiaKD4rrigg8IgnrR7X3uRamIQlNBEe9hmaZDA0l+Sr/tJ3OfyDqRTd0eKweyYcExMIM
251cxc0aVoVfsf1rSRAhjktNWj3IZ02HdRJAXrfXWoDTvsGGGhtWByLdSINuDJuHadGyszXhmuOh
KRJk8SW5yuJYxp597WDE76X8MYzFtd/UFTv9mPv4eLwM+B0HMk2+vdxbaWfcdslLcDbC/asoLrw0
h/ffi0GlQXoV5+wlXFAMq6Qu9Q5QQucIpUuwMdRdTE2yjvq2PBPxXxHBpeeu/HLteiKHfu8A/a9x
Y/8QrK7sNZvp3g0IbYcj0Z5GjmTZqnRGCXKM2H8bCBiM/vRmvY7mR6T8RTBDUCAq3GaUf6yRXNm1
cupTUZhb7qrY3YgFDWmhWd4FuVNsRKSEaqAZxUYq5TOTRSTZaqmZxNJqGv3F7kStVs90+uO5ooAd
XNTEXPgTiGV3S8wIN5rWo4iJFgu5soKqk/YXP3KmZZ4v+GqADENeWqPuGoLpRWFj7ovyGx74abp2
c3VaRLD6O3a+23GY7blc3KPf/eogMNKaR14G2ssMTem+sWeO1KsA5exsMc/hnOwKykqlkXhYqZeD
LXEsjJS1fueVAisvxbvAKTH7KIC4n5vsdkMtOXI+K6wFR1cNwNTy8AAJVK0SHwEurZNzISeugdV2
3CbLoPr+7l2I+HGEyazYkGqJO6WN4LVr7CP4wddidNrHRFqYzTeYKo0QT0obSUTgSkryDFYQlUWa
rIRX7QBloGKg69sxnI3u10MBy0vcnuEQKSGU02brJ/hORLyOWGovtNi2P5H71IJ7Q4EuBDsJ6RPt
rLuUDn+xclwKuFuGNlr1mG9Is01AX5fr4CzU5pMGvwuJXK30yuomtUI0mif80gy4Vo++LhG11EF2
oKkB+uMe8pQIfDfy70y/LcVdiAth6ACsVYfptih6Rdua9MCbzjFkN5KFuiEFmFkHhdjK4EYszSJe
yBxPv7fixRBle9ULj5e43k3hLeLCExv8tsywBAZ2gqZK9GIASUFlWRxf88Wtja8v+svNW3LP7agF
O/30gDyiwcETzHCjIsrVe0I/pMcNuO1Fa6MArtmcHa9T6osMBvYBDhHHdoyRBd/wohQONpVOTnx1
NjddU4wPbWMwy5OtXusceFPdrr52V0RscHU0hU9QE/Rh7Id18mAc+e8nGpI8h9GIECeG7yG+VWNO
InDSKj7H9lDLoceYTL6kYdyYw8M/lRw0CVmaBUIxSh1aUwhtk440f6acu8+OVTKVWEamtJN/ElSX
o6F/HYyc8iQbp4YwrG2iKu+lcLcgxnPLrKKBl/M1cuhv5xKFtH+G3zW1FOhVLAOJAjLdfLBnriHC
ImbswmhtUs7jBf/LzyzZkG+IxY8MDK3Z1zOp1fxNHtpnzsRx2njXCZlA+al5en7iLiwZENF97Fr5
Com5lz1YaiyRenzg8+8NosYIwLALUFbn07Ga4Xk98b4l0IXAMJ/aIShsyl944XGnSmXZB0Qlkgo+
Gzna215rUOQTvqAes+ELw6YmemRXqaAgFCIacAR8bTvFQdNzKqjQc18PCZtOhyE9qj5pTH+xRDQ2
+OS5F6Vukf2Yj6i6EaDFt57AL/aQTDkSX02P8dZZYJPdVIzIOGqI3F0vVS3lGm08xKkqr7/ij7VO
y/Q35OscTrS7KT9qvVinIK48kFH2/cvJf7+qJNLZykgTMcW9O2VmjjG6EvncbGQMOcO/p+FGS8vf
gtCX0t7dzaagTjBfTgZlFFc2XzNjCRTtQIQpWXH6PF/6KzctuPsbmXd4mk5sAUP737yPpkyGwegl
t0d0Q5A4k6azcQrXjuz+WhJXbOCvRAEKz/mV3vgN93qY9X2AXLOWoCL3UOSauoVF6OggBjkfb1aK
rgQeB/4jEBzpYIKC2wKcjVFaZ8gxKYV8KJgRqnamNxG1sJ0+4pHUDD/jWM8QYeU5c2Rz6ws/N0co
BdAgEnczkzYY727m6Kiwg/ItnDhbY8cNMMDqAEEbIX0DLsIt+U9hKJVGC4ADitQ6Y6jBUNNkBCz3
jSZ5OQUYJzZ0Zuj04kZLNG7H+DOOLssL6JNshNFO+AFNVQMY5STQ/JAoFUDcMoGEdoMhOvFMD8La
1jTSmN0Y+phHNIlY/zoxSnjvSBS9Vw8WCDZ0H2cLj/9hAx8kdAtTVTSDx1rwsFRj3A3s8si5hgnQ
GzCfqStpAbv17jqy7NyhWVZaYZw+Qw/MEYwIynemwpdf3LJwMh5qZglW3SyZnTWP6w6hzCbpkTO8
zJ0cnmdMIB88lTKpHP01dpy0v8r909l/DdqxN9dFDxhBKBU98ya5CkTChRNQ0t0HxAKgRKLSy696
ty/h1+BS37U0RoR56Aq9AAFiw2FO/gSo3NJ+iSYIbdHkr+Nefxswk2Zn3TmZXSkGkO4MWneGRnjh
ZTA8PBPl6OzO5HO1adFGrAe5XPDU1lxSaUR6QQ+Y4U6q/z8dcxZc5O5YcsEHhp50dkbKTjpVM7IE
V+jzle3TGgds9rQfYYwLvz1dmtUeIT+kuRTsCGtsUwQCS54Jk6UUSOsgrVv8moWUD0QYP5HTRAVo
Iz2TN5NpP52JyafiUMi5O7G2RJrCh12CJ2gQFgELTaWK3jA4P2mqXDPg4X/UfwUMPkbuHudwndla
/rHuY1PEAmorCxUhfgoOA2sH1pRE84Fl4WevQ/b+T0pzQ1OkaJKhFcelLgXu7lfHSdB1U4RhXygb
b3DWtxnEcANs5cKOISbzM7eqMxCxRKb7J4G1p8zPUQR8Zj13Zv5QL13SyzOdYMbABGpaJLW30a0c
wvsfFx7r7vztD4cc3tDN5xGJdCvkmmizVkz+e+aAKipH0gpVXEWaXATtMcR1jR02phLGFfDhhdVQ
LAB4+aU1lOkrnLgkoQeLrzvjPL4cQ6mWSFuPCVYr1Kj+iz2sPY5XTBpHC2p7bNdmaCasPFlzCYQf
u5u+wf+7lahMXDGRi/PXyZi/8WTqvC6Lbf5AtArZd1sfBfkFS6GYO5pWZG0eNTXCm2RBS4ID/iET
CkkQMkARpnoFSxtwduP0z0KYzVUrMnujW0UwtQ1tGrI2xtyoIVxTLvxkV4QrrtzTXygQDQG00Ck9
33UXc9sIJfd/1huX1dpjHExqFwxYZcZpmTa0W8gfNw1VomLbvKUZZpBFnYSsWMTxbo55fs/tQUJw
EV+0V1AlOks31Of8oejRXPZtUEAbpDyWfg0MKSReTauD0QjbuLnNrVkR5LqDIpuEg1bOF73TaLEE
fXXTlDR9sS7FxmMd+EzOepru1jA+a/0Akx9AAghzplMoYHjyKUl00P/CxXnUq14eakq67LD8TJ2/
uFA5lp3o9uYtguNVfCMTUcfy4JhFjD92J6jgNoofrisXF09cROZIU2tk9TPscwyGXVFzj5rZ3ZCJ
XadViCdzkyHMFyHbqHRW6WWzzBcUj4cKj6yntWPCW1DwC1hdHl4d7qlRQow7LdM0yBHne25x9vRh
k/Ufe5fvxQ1op06+8kXSUnLP0TJBa5Btx9bQqdv+fvVUkYn65A+PSpF903QRXO3Z0BPXXJ/jgvd7
d7oAKtO1vqMjyQySjBDzrJPJsy7v36khATARvf6N+WgIPF1YqlcHZxLdtqLWZ73S7xr4dwlewK2L
37/6EbGgRtCSLV5KpWlDHikliC9bJUTcQkUSIRBOnYvkECI9iynIUWZpkt2Xjoo9DSOUzTSFTj8u
DY4vObCUaLk1368GjhUt6ntYOyQVykiut//X53fmRQdFVyYWYl3/Mr4eJV9Q+PvMWLdug23gLq4T
QQb4AKueCSW0XsyTUJMuyoVbodpceBb5z2icjGVVijWFKVWw5bPe4lWfq2r8i7eJfZOuoN3amRmc
8O9m+/vE/432/xwESH6ykeqfyzV67SmDTFF6tYFoERnnxR3sGFp8BM+HbelVPf44MR2pu4ti0Ik3
cnMnPWlOcWbjJIINUBNl3U0EkrbOg3+A+A4Dhu2ggrcwv9aRhJ/NIjc+1RN/y4Gg4pCRJIBOFNBh
WzsS1Y9+oulc+Q5BU1UqVlkD3Rr5elFbtDwM7eGB5pttRDss9cGkfNA7hhSC35lJ3rxQy5xNpe9X
nEQitAPMEam2NnaFWdW50wZemBA2aw2exXTUQcyw0tCCAZ7JORvJdSnBunpXFhRz2/GRs/Gq0L+O
WmgilkTifagJXnOvcccyC0mPkJLGJsd91jUKLDOlXtqR2sZhmxrvfA9y37GhrS3YIAq0KKN6l1qZ
+wxDl+ThPz4LkQJmnf8OJzpsJinWgnHYXzXGb3y7/iXtbgc4SZRVX9W12bTVOPFFMgXO1P5Q7nF1
VIgup0JWphp33FT+iLLS1CwlejR/FL9/w6Eh1PmWzf/5X+r3gnML8kmeBNEbHiOryiIlZiURNEgS
GKofG5t4lZ3+K/Y6DxPIstdNDtE/AhETTGXWduFYjlBwnGiAl79akMrPRbzpEr+MnucmFOjzR+Dt
ytskMA5MHEfsrqVb8BCWhrN1SI+E09qNG4Mr2KqSm6U6V3CnqwzRS6pEydS4S6NbUdswd19+//RB
b3Wh2uSKxzV4tiwdd/9ljNVJz3f43ohqYy9jfiU8LwuPZ6/EleQZclXcrnyVfhrdvBLfelkfnWtf
0bMnWGgL8T7cvcwM5DG3KZ6sJmt2U8U61XZQOmJATdvlvAgTh/f9tcIwLou4c6IFf6dpVh2MKbE7
zQHwQlYHiouc2iXgq0wSmhCymoMuBNQJRRQy5DQo9Aw62MnqqgswhrmFLkVfUlFAKiZPA2rgSOcK
koM/kz1WENPmrvacDHg4Fm+3JiY2ZZ8x081rv6zlOCaCwNnGyzgySVs48Yr+oNXOpuL0TW634T5g
SBGFUq1BNIsqM2lMtfkViBhytxYiQK7EfuTFETOsSZu4+bxiPL56KIcH+e9tI2hOPiUwQ+ewPI+5
kfq3ei0B0iqhtWdg3j9sOtxlZMnrhRYspmhBjAutJvTFHGvwNkyEgApjE1IUBM2MdAN10n+hUwD7
jAIWpcaRNhIcUDJALJPcFa/Jv60KHL7Op3eWjFxb84FUlpgfSSnC9dDS1h8z3QTN2uwERbCXn+CD
mToKDZELpgTvfkULWJybqYZd89HoVjFa/K6WBR5Fbt72t6PD+bq3cLqUhIksEVIWDBBoUSLHlXHH
CtnATeZUp103aUOIuB55MNGqCPIVLoVTkSBVc9dJnqK+EUhHKWfIo6E2jmv1qTGLEX5K/wIiBVyL
flQ7qZ8h67yjW3WxxZPnohC9vhRGslpGaZhUb6kA/nnSSXIUfy8xQbamZwSSSHSQtjT7FSL42Wmw
hXjhbZnpm1oL4Ghi/Y/nd+wGH4FITCOyl53RBlE9pAZu12h7Ex5Joima+o7m3ci6FJBU0euQ0KWM
EJLihkDQ1J2nR2uSxm+Jdv/QGt+HcIkp/ocORaJTjL8YMaqusYSivR8k/u1YEQVHyy9jFynGIGXn
nJRKro07O4eRoyzxp46Lkoxma1t23qzd5WeTVlzH8sFMAKD2WmmmuQRa0nf1fPM7aaUZU2m1vBFQ
JkOSqWtr7DebmZB49Ctss6xHfdoOFMrITNWUf0OG34THq5Io7nkFT5/yVGr6eLXl3pLNNQWjvOC7
E4p/b138qdbYg1WduHoAELf6JKLp5UbxNIqnZeKruhuimTNxYo0lYjL+93+rHsXATJdXzwZAhkDy
LLdJamV95/JelcbkK7VHvKUJqoaa/psok2LZoTudEXKPAK9ktgKgmF95C1f9H54eGd6r+fGGntrU
rtcbP/yILTVQaPfG9Ehc7sRd5F54pQAgBEffTgRi5vslEszu1DOMppZoM+iwEZrhzxyAIrdLbkyZ
mRmiP3ApK0KZ+zGK2zFuhIUeBW4tq6fYysBPuaqwQlnO8hYyUD9JV8Eg+fb/aQ4P43Lh9/xzG8GU
E9Ls5VzZV/nvIFsbKddreCCksa2HfPD9cr938/uoxzZY9waEo+lAKfO4y+bgmuEtiO3fskWzI5vW
IKz2XiNH+qo5G6CsKMW0Foa6hIFMNMh55zlbDrJS4YSZcx2UqsKo5Amck+meDxL9sb9iOZQCGVeb
mxkuJxkpmHeVVaJINUNgidcNVf4NVAk5nX60uFLrUA1LG5rJ0VuqN0/MW+MeU38Bt2iqH/iL5M7s
vHmzUvqG0ddzdnlDtI9Z/HXbdpCK5hqbH94ptgsPt4e4VzCcQHPA5PAweC5OAbRnsd5a4W0N0LHq
NnyJGfvI8qR4x5HxfN6kDaIrD8VWn3jn6wB/XnU0icPLhfwRo6XjrpmSWKq2QYC8abzN4w278r+Y
dS41l+J6DeAwZa+PV9XlKITsEA4wXc1N9JBeNYlZHFNm9oQfh+/yNJ0n51zamVuu/OcMV+SQwCLZ
8cLQNNIybwKVkIoo4Az98u1kLRfTqU88jjWrWkFnDA31jEQHueNSweB9NuWi4GSYpUDg0wK0m6r7
UMd+YFH0wJLSkIkGHgAP6gkK+yBwa2kAYpl/I+7l+KnOhT9Mz0RbnOjUZ5G7dgT6NUN05C7y9rsh
+ZglYWps3Z7PwRW1fHySSR+3LvFxq/7LOVZ2V5dQ/I4yyhLxRLSyRem7ETfncQvVqc0+YcIT3fu2
M00UiyxYNvZ5GflZ4DILPCawo+IQ6L2zBiqn6wXHJsYD3JXwVuJgJxnMQTdcvKavS9MALK9IeQqO
odFPdns5oFeeMti+l1DgmiP2g8xRmCpHxQhYWKOklOSD4+2bMFXmWyD76VSkPXxr38KWU1UjdN3U
tZUC/wFvKvvcxUa7iWtZdWkkzRdR98j5jpFWVNrlc4etIcHWHLRlkvif8bV+e+cxTVx/vomDvBw9
jR5bKwZIkgiQeMVrCUyo/j3PdGj9WDrPKCH77j+PcLTi388/Rb6D2AOXbv5haWZZ0YkAkJ9Aa46j
CuBpFhaYVsZ3T20yGhzROYceZwgBpqHKJ8ZI32FK7vkl3epJ9dABQ59GqNG5XxkwLKgOqHw1M4ze
cBKRJL9KLkqzwu2SWS7FhJ2v5O+E1K8RCtOV8PA35eVvdw2qI/M3TlA61ui11FJd690u1F2eUaKy
795EU/6MJ6TF7kAC8gGaMO+y5hRVYCDflgX4/IO+ND+IrApeu5sAbB9Hkq32P8pChlmnkIvwGZsf
57fL3UAOnBpujMsf7zZDpmfXqIZQs62OfIESozHi9m2iKE77B7zwKL7nr2uLEKzY+69QZEBznVkY
8sKQ5VDurw8YJs3xVSWyikmGmCMpsMNLGz4XlZsQPQMflUqT27b6neK79QQ4yk9sLYX+coiIPiVD
RXrSsviBCaZGVurvp10rjelH9t0cFF0tFI7kbAhr0WPTV/1X11W9cGy4s9EMPfolPrE/gfJUIjTj
DuuP6LXlJOiv4J81sq7cQffRQWyMPYyj5Ijx8yDdAOl0MXod0teUeCf2iUPXonM7uXHhNT12J/pd
fUTt2nSc7LNgYp7sw/0h/KTfzxLywL024gpSBGQyHIo/6JtT8EPD6K38zuoSH43retoRuIe8apjD
71e7Wfahwjlr1wG8qGxTHZl7shI7HQoWwkkH41Ew3p7AtZo9mGS7PP28D8lV5FsSDALDfd/zxJQY
6+tD2gILI1Cwsa/NEH6KpxBJ+gK2up3F8ejARJIS9bgez2eAdOIk5PGzR30DX+u7GGRBIUzxFks+
OIKq5OZrM5sWc1AG9Zl9dzZJVM5GFIXHUh0rA5DubaMXk5sVKYiN5tzjdyJ8TVyZYeHMs98m6pRt
CIOpThWNuzyFxLQO+KCIUaLWZK5v8MIesw0YwszaApiyPwdEGgnp6xA/avXSjbAT5D8f5vmrBAXe
JQg7ME7USIajKy2Ew9Syu/m/+vEDVSVZ9PbVmDD17Ry7qCGuAD3oNc5hOQQfxJWlITrclsu39gLL
fQMxqUCIzWc0mnC8vOPyE0dOk+wDfxkt+Wrhz1ipGHUASxv/hyb/ivJILYNgnFhQh30k5KnKMwEK
cXnB+BZXdg7bRfRACTLt/p+E61ttUS9Z3X4i30YZKnHQoIYzzW7MqE4ONwAXINgmiSzv9ZkJYKOo
L+JScoEXq0rmH3mnoOgNq5dLkZMm7Y+n/R10ULOIVh8PK6O8zyRbI2Ywm3fJ2p3rUzdLm7uPAx86
6UpNxW9qTUaWlQHtn0gt2Lnstm2r+RuTJnSe3iNrU9fXIZAyqkC3ALad7bNKzVs3Fl0XQ7gR0iGE
9dplMV9ERygSNZzjhT4eDagfVWt4Z2iYQWZsp1p08UayQ1NOsPGUmb0PNdxxmc4kwqrR9/q0FfoN
cn76oLqWzQ8TnK/gWSzEZ9O7avtH8TDB3kjkIffYjv/KAtunCuhQpfJ+/O6G6vqVEi/u3yev5J6I
1ihV5iyOPBcP4lTdl/K7s+jgh5k4snvQBDoTa0+y/m9CECv35SP5dxATnduu8yIj0ZU4YJ0ljhre
5iPndg/rkrgAHAJYLf5/bi/lRqkYKSjtv/CJduncYgAEvMzhYTv4wqSAcQQMsiUZI0SP0sS0RQMY
ZokTioTIHYXvFjylfeI96vDFb0AasgvfZjx6v0L+fh2opR12Q2Dk2g4mmLFn8PDz4jwZ0UYj9UMG
z7a6kOTRkXAXfkTceVawCQuPneDLquOg4XYsDQWQsiv35liUFHsZSl5BANfVByPImqAiu35xN3Is
iAmib+tmmDkL+6PmVIU4a/qZrqZgakVFGsqIuJvuGzf0OQwLJJdimQG7sg1+7rFbuJiZ3QcrA8rb
C4s/uJRkbDpPdyOX2RdJV9jaKBYXdj11H6MxmjzD6dn3RNNWTeizWAS0ayx3f2+N94TB18pt4CCS
ZzObRfHukbKR2/o+MHIEMhvvW84v5t/anTILjmGF1ytPYpezNaZ4s+z4wS+AGXoFdJsb+BujP6tW
zHaoZXY7Xc5TLuIFlUrRk5o6cvJxsibtc+Y9gEpjaIk1RMmVGe8Qx/pkm1Am8NVoLkR3ynibt9Fu
belbluJiDenjtJzQmFGnzTrsbv3HcpFPP0bmvaPDwOQLumNHEdpTVDYDp01A3cs1J1sUHp9IFQOb
lfc0CLr05JDs3PgS9+TBXrAduYWIZmWH/tfjWJe1irP5OYHhTGeYwE8rtfBEWVAO2uHJO0dAyaPq
nrwlKQL45mxCF+IMeNrxbPgmWq/6NtAOfcTNjUR1jF5EfaCvETm8gdBE+GI0PweYQ+3AKgm6PvqL
Pi0h2kotXc5Jf1DeMWY8qe1vYpIIrHoY81Z4PSnfNFdnFLkBLn9YsykMRDk/uQ7bsUR4ZlIXhC6N
4AnONybmiOsE8Ys7FubISWQYUlhhZI1ud8VL+t2Tdj0cxzUl2FtZcsEw/nWLcqetSBJ0OgVzmmXj
UfD+rFh+ZsAUrNCi7AKQsNAbbEClVRI/EyR/ygjXiOAYsAbxBubtDbwy7ISZWt/F6ImSaHsbrRwW
nPafDjlF+wS/psqjtPBPXQUDwg8oooKiUWj4bf2Wm7t/4mlXRaDlTpXZP5oINegUe/pVVoQZ7NeK
FFcoZ69XovnmUt9g0Q+nkTCXd6k1RMQKl/0SSB2XWJjhbqmCeAQMty5tGAgBwrALS/STCaOX3rOY
z6iWHkXZLFs6QgoW+eXW6k+O85qW4iWySS9qId6fc7/uyHHWgs0mcwx7oKBI6tzlfTjSwiAFy9c1
IAAohR/WK+fH74aAc2PhS0H/mSwvHds7KItyVcawC9tW0lNX0Z4VsQOfb+hueKa4umEfEp4H6S0q
DDHJt9dtaV8G6Ko2oAy0jfux36Nfa1WSMKqQR7bIunvP2RVkSPxeGZXmfdR0tvplZ6WdFnftCIAv
9D5WTbcENYi16jRohzzQCNnqNfemMUvx8E58DI5ASh+K6xY0rSnkL3dcD/CSG8bXXTM4VBPqGH/l
J7znjB4mCfNQQ5/TRPdgXkw/B0XNY+ydn2J6z4jWztwJvMJBWMRB3a6WvhYWBur0x8ju6nzsXBVC
ZgqqFe21MPpkWZkALXepqT/HnPQnVJ9MbsmtfW8y+q/JUxCrTpyiL6byikEa8ROJq417F+Jvblh0
Db0XEqB6P7LJIqVRNtaXbNmtpjlh/GQXJ7K83spF0pc3emCnCvniF2zLAa5+7P8icnA/0w4YEDmv
JTqUNM808V/8t0qcS8NZiu1lkgwf/S/HZ76Ey1c/4Xi8z/hoNCsp7ga1wcJTqSi0uZYu7Y5N5aVK
BKIlAXfTPD1HQW2CbqJjpNpjoETahxN9/gDtLqfWtnEzR9HMqJqRhuW/eqYmZHPftLd9CVHxzUeq
9zjGd753B3xI6yPHVT4T5uUJboVDo7xzEee0fpfZB02rSNrTcoXt7/hRYEZT+3WsDRs/PMHG8JL8
QPbeuezIASszwDZvNHKQ/YUB9GEZHYTC6gnhkRkbclgIOlFpZS1mP5XnGFFjMATi0u3fQV4nPCF3
Wi8XEshfv20S1bBYI0YYj5SpE8ztIFPdlUmbnVNLVgzBwBxUoBzMys/Hd4yF49/9FwH2ADTrw9zN
ltZtGALqiNfYow+miUcjlN279PdcWRNvpi72qfO1TviDnoGSGo9tQ9CLSBG2H+82rDNhHfs6Cft3
5x7Oo10TSHfr/ywtgKIn5ANpIYf5Bw6ct06nBhDfoVyu3TmdQ40FUL5GO01WlU1Lf7XAKHkdJlGr
NdAdIo5GEiv+TfH5RGwdpdXqKQikOPlEayeBpofJ5nL+/D4dfXP5nEfw0uAUOgGizDRMLRY4gsqp
7j0/ktzW8nE1CS3N5I9m35KhkTajBPYjMehxfXk5EcZAjlPa+gPieplt3jum4I2y29zbhrOYla1x
tF3qYGnerliOU2+9qhDeykbmp8r/qww9DMt6EMaRpQVSdAtQfr/MEY8t7X7KJvffdx6rl+woJqZC
TibuXkSD/YCeU8SmqZaIy0wJ+ObRQ99Ji9cS7ndgha5QaMvCpyeZ+T6CvMJsnXKjc8whXnVNURXT
n2H7FzGwRY9um0eCm8D1WgvNKbjwktT9wJmXpkEM225kNODBkVZXq7F0bfjezSvb7kbfb6ehlNVN
omsZbYjAn9ZRdx5Cz/FtGsPj0lKuwkcwslx9dLAUXY4lA0pLt98J0ZW4wUv+e29pu/mOYLO2TYOJ
OSdLohPo0VyrAB6rwQa3gGoNeQMZva3J5RmoMNJlss1tC8ML/scvp2seT5dLTlTD8e+swVfdCLG0
PYiILIcA++BBdM37DV0BUFo4BsVKRI4Z2e1CPngNBgK8qTQL3T2mi9dXjEG8fBzHCxg4bO5TLlkS
fHER5Cbr4eocx4WjWzLQNF6uWql02B88bFApMolQaqd2/g3enQ+E5RuhZaweWUxoMzQvEsbw6+rM
VepEEiRPXWISKz6U3t+Cy3eS08PTjLr6iVniGxjLp1SChD6HLPwxvSm9w1bayZbEgMC/S+SyI9pS
bnGL0/+Bspnh/UHgyq6yoDqJLyGL6PWqwm3OpODQUSpuCc9a+wKuFznedhTlK+9J2n1bA0w6Szpa
ueLcaquqEFK3dYWJ3YMzqevIxE/7cRJJD6GKDbW8/slPG6H8C+6V+TCJLRtHAk7lIz0Nuqqy0wfY
2uUC3pYSODkufJ5SXVHC3zoe+Y6rIlUoDkA+FMZUwyYATrFRLMuWWQ6uTpiGwxgJrr7ARU1kRiqy
LaH17SYybdhy668aNd/StycskDbtcMCzvsrV0UvN1fw/cxw8JncDEe+N12C7LiQhe7ehjpFxVxWW
eIp/KhkXFcMmZ/ZrcJtDO7K5wHUtFtqgnKNvxtais9wsM6TEE5gcbxga0MF9GdFbsk2E5WPlVbgx
ehWQnyPqPbIKbYmb3wpDOb92BqiDFf9T2MRznLlj790xsa8yMdGVY/Wl6PGq3xxED0SMcx63q845
3kfRdIpYwkpL9B//hCubUee9K5fFp5MKcvOob1yuD847TFgQgpQKbqLwvbD/W69zzd+/bwWLVeUE
r5GyB193wJrlsDlPRf4F+tADkLcfYB0judECWu2KidR258azacCwz9hpPmrd1Qt0yQ04MlPOZGtU
xMSM4PXydb3KqkTGqmP8wKbjC++J444elO63KYuZdm8Ga+qjB9HPOZhY6EtwxHInWgHm+CZ2xide
KPrfpWYuNHmtuBzsux9pLHLoPxoBb5FE16+CzfV6BZcTET/nSNTIrXZifEWj8YnmtPVT0cHHk5k6
u99CnWhmECppiUpFTy83rZIbcrz0lVcjnZwG2kCafcOGD0ngGrqRPdXLgrnFYXJsoN0gbTS2gneM
lLlW+cM2nk+w+FxifhlOWZzrk/ASt9Ss9t60HT3TD3fJEn7zyuX4yYyEVpMSLAlhpPpvJHt3QH0g
KULGua4Ixt0I55aDyqHP60qE2TdaaXHHepQUI2TPSCI33DiMoXgM7L71iuBhwbmYfvnkyKyz0+R/
VXd+pwzhHC0kItpr2zzdEeuZSML3CNpdC5lQQRoQnK1pVX/Bgph72h6TKlGpdV5Kz68vCy0Ir2jT
djrJD1Ijf4Leb+Wbi7JiAxkubdtjYcsCm5awFj7UG6weGKS26tiie+ZDVyoSV4DIg+ZpmXtEnR/f
my28pEb6CeyZaFfivco8EHi7I4Mc9rcF+kQwnE0q3pBR7wlFr8JJsITXSorb3jNKd0Gqffeq2/Ga
Rsx0ZXF0cCJl10SH7SFypOQydu57Rfs/aAiR6myL1ct/qLk9+++u+pGRXfG+Es4kjRPp36bcpyEg
hzJPjn3+9Ztl4eY4IxX4JNhTfk6Ws9r1m242aROU+PHM+wUZkszRC4ly9usoNquIF3mQ6HjezDbA
GMC3hUNbqONYHmwoM125hr763p0IIoIi1NAxMTXIbQW1ckoCBxI/GZNfWd8sJneO5bLOGNTdBJgT
bKgXutTPkFBXswXsuq3MU1pA7PMK59rrTF/1pQL6kTipKuMCIqnWKk/hLtRVt5MLu8h8iLqDyM+i
+KVEz2HlTeHwJrCEfWLwka2KsjOJb+9U8DA8EhNahrQgVRXhge40NeQY7Q9xWxpxoYGEPjngeRLp
AbJpj/X9oRbxAz989XEnQMM2kWI3u0K8mwVARkzvSM4niQD9/pIISy+h6EoeopBN5Ta17ILd/YGu
xUgLCFgn5vxzkKFPBrISUETJdolhwWo5/YVXQyoVlXrmDDoJ+Y+E9B1tgZQctsQ96NxtZ8LkKmZi
DIiYj2Ue5bvK7xY2gn99ZZKwhZM9XVxgwaZFuIUD0eaepUl9hMJW1P+P8icYBq5Zfr0CfCZMWu2z
KoIdVc7Ctg+Vwi8pS5qiD6td5tDOfC5RY2iNggoxlBtAzis5hjP6OLifkF6HkjPs0VfU9KEHIDcx
/1Tx1UZcmo7mbCEkBdYVR2BAXLlX7LuGuM3iMitLAfKNQXvlq/iH7tVOLWceJT/Wo7NMRY6HsN9r
2zkWXAxzHBjAM78Y+usy+dg8fpCo31e1aZQAaXVjWV3uo6l1+WOGDb7ybe7mvQMgMlEI/grDi2Wq
3peBq+ImRy+3bpBVBBQXKgnRax+iINlO4mZ4Ff0McESkg5wvx/fnNU2e7dgbi0vhKb/FdQhWSZqK
JrdVlFXEqF3XZfUKcCnkY9UTiIUG0+x3olbc+OYxKLbG7JLRUlccHLZwTU4sfNzzsXTNghl/A/Yz
YArg/+lNNhyQd3XXzkqu3MrJqBli/fZ9BG7oTea8GbWoADzzZ7RyPgssGnC0fjKHOiNiJny6Hgd3
PQOqyZc2NllNGwoEkZlQNLMQcs/u4OrUPy1g9dbsc4vczcURg3GFU4ThIa2u38xCJBWVNj+Xf2Ea
cyPWyrccEROYNAOLRU1lKvQgyMIIUezVfaHKDyCMqRcmNfwFGPJP4RfkiZAB1yCVU/ftyezHmaN3
kcQFHlOmU0wvKEAZhagGdY3aew9qFed/DaX5ThEvzo1yJ9o0uQq+0ubC2Wn1jTe8NxZblWjPb5+H
XHiDZ9Sbbxub646ZmKgjYQhmdhbj3uPpzxbPgSxxVzPh0SKxyEaNWw6UgZsL5qaU5fS7gXH5WNzj
hpFRyj72MmUMJkT88/FdYdn6XpJrDjVJasB7L/IoZE3k4q4yogi/GwArFFMRxzFH2seAPjneIpLQ
o2hEnEMeTVFn3EEHySqvFR0x7Pp6/9GYL4bk6m/G6d5ZAjoM4unseNXMI+InSNYz8oPEK54qZFV7
tXUtvRYmqv0Um3yk40miS9C9HpvEAAWMqa7HuG4h3zMhhBOCivxHS2Fb/AG6hDn0W03DIi0WO42m
zNyQjomRDyc8/O19JEZRHnn5B3TfCLn6/HW1RcSRbpSxuNOqSudnwH6MMFY31PwOLjfSqOcgdFGI
v5tGOJTIOqjpwYMtOPA0G+V6O5w9jXGbC6eD/xzD2uEfkX1+8N2PbDnMggqw0HAqS+3YVHWh/UNa
91Ys42sRTH11yur480D07X3PYIHW1+G15uW2IJgH3xjA2bydu6I9YGrlVTFFBk0Tkt+rysOSSYCw
xZhHECtrN3PVZpnZs4C6lkhdy9ibU0UWNO5eBSUeayLK6FWM9bRpfTJXv1awNpCWWo97d98OFrI1
1hqOJVi+X8/Uf6DvfbX28NRufsUqKazgUuD7R5vnE4eXWwrO4afQ2QGNB9GEEIYyIqsnfs82eFgs
WFmZc/sf3dsRbN1PVroshagxJYtzTjQrzltzuKqOZkhQE6T/mZqowwdmLyHYkBiGh61RRyFHKXRV
duIzWPqD3gY11Wn1GLL60riso8+IJKib5C3/LL7adIO4uTDSsowJK7g9hzOY4zz+Lgm2cKnAWLIY
ZFL8A2jSHbwKLRg/ALtFHcOqXGCNhelgPlk/ZLWdaDCxA5Uj3c0FIeztVLt1OvGJ0bx+b7daOrLo
Jn3/P5Qu9ozfaBSP+iG5vm+7/s4tao3AkZlZcPQXnKL4TUqzmc8Tix34AauJyOwvM296lxeXVCno
lXfk8myRB6NIMHB6ZteoWXWF9cFh4AW36jTD6Qx4YxRSgZVTMSCaImqHPnZyw9QuTI+snc+/KVh8
kXWILWkLNMr9h0P/prMW8YodHpoIQagTw6zFM3qxSvLrAsnQkn41M8zsMig/0LSsscQe193FlIt6
ZiKBW0d/BZXH7fAtX35VAeLe0WUUv+EaUEUpWDagW8sjKZ6NLB4H4ses6ESXeuf+yWsLUUxvWgD7
PXPGA0MK1CdtWOuzO99WL8Mytv3MrHQFQPtdajN7N1HJqHySRaXuXU3YUlMk4eM6WfRR/tVebgCQ
ts9gzFlrCI59Fu2rF4SnZeESaWV0h/6sQ7cOh5KnnAdoT6l1ubp6W+YyTWjaTJeuXQhJkBZwJZSo
UpG4fmTNJELKs1zx2nbJK7HDn1LBQA2xU0Xqyc2QXxE0JmusCzhxg0ADF2hC4NtQ7QwhncQB2qNZ
sulCXseePHFIMIKY3tlByqvlgQxa+bqClZEk5ded8byPKU3kJmhYt05yopVRMULMFYxXGs0ApBen
z+3AMTed72TJKMzjr30ZIizVdgRM2Amiesw+m3AFtPdfcFXoPbg7tCCsviZSN835ZGjs8y1zhT74
2QVbVU9xKQCiaL1qAmhEfBCyKie7JgOvOgSwFS1zhpM7+Phlu1/Vm22RV+5zDHhNUz1yEeaxkT3V
g4bvYE30vDDpSNNnWOTP/qJ8PrIjIg0uy/17z/sj33jZyR5LwiIhmugvXPkhsmbQHc/x8K8oi1c3
K/zORcJpaW7lpMQ4nnv210tsbz4hTtjLfaqZrs7oRfVPYGIp2ZrKfrldEM+HZXjSW/Ep3ztrCdyP
C35VfAYCIeiy7CGjgP2tVzm/6janWq+wesNlooug6vTHQVEJHESs0qPBSifiEDkgpq1BrCS4FqUk
AOuzeNPDw4ZJox+gWitcTYKT69CXVtA5pYSgv6bfjDOYymlplhb5j2UDkx/OWjLw19KCnnKdAawO
Awa8dUQCrmdv1e+hJbwaNf/Dk0/ISox854kuh8PpzIxtnOOPdMJ2xbSS4OM35d3s2/LK7k4m08V3
ekx8KaKo6nkHp8khSdBSWBNJU1T5L7uGXFgEaooym8pKNZbDmGmcJ7ExK+QtidTlnvySv1geRa4W
xQhAyq1pw7jwghff5av08zOd59voZFbWN7isibewu93+Ycs6SwO43nKDQuNShJO0zPUgD/E+VHSq
sqAntb9S4/EH4XDJgkWV15SdSXlEp5+IFvHjk4Sv/55BxHM4X0aHiOPzpnfjRFBs1hejvtP+ToCC
IJuNYyZuSlvqIK9H+nXo5rnMnNHYtvfcbyavTNxJEwMXmOirAYAwYz+HqOGy6wd6kf8cNNrQ9Gcc
ofxx9cOES03lkRuJx1b1moMXfozDxAFFg9qLm6rG5LsGsxgu7QUv1Vm5osPHg6yzdLkvJhXh1Dpc
cIK8emdszKfpDDlgqMQYgPRdsgXiH69pKYZ3iadriasntXRAJEC/FpfwsYQ0eEQSspD3eUQ1QjzS
xoNZU53Q8rGThOiKE/mFWSPCwzyMMgLFHH9vFyvWeh6vlClv9DcZcBXkfKTMyy3SFEyUFhtS4l+v
/jmis4G3oaGtO5NLPHvhkRoOtrHcUK0T7/ZfuCRpGsbLHVtQ0pc7JD3o2p8MQWKev+dYGrhEX9jk
VjjW48K4iDq/L9yuc57z3IO4F0qyPp2ctVZFijxmYwP1mmWBlc1EYcwiNSKdkwgcH9wVuo6V9OXQ
TvCZhw/JYnF57igj0wKJ6pJr1Qkz+DEstZiiGSAcgzMPK75ndzk8Cqd4k6ZWA2WYeFvAknByzpqw
KaMoQrBHtKPtV64cDpkkZ8l9D+Xmcgi606mW/Fjg8MYz5T4AVela1eT6XZqCMK5GZJ0Lt6jvTVVn
UnwsjGxXTnX9FwTG1lPaKdY0FLg0R0Eo72HzLF6ORp0gbEBBL3oCT99bisSs1Li0OmM1XQavixsI
dePUxxWlOWpzdr7a6yDAwVzIrhxY+QOHajqJSODdIaJ3FkQGIxeM3LfL/ptXYk+M+CXvhsql9Qcw
BbH5dueBuQzspUeSNA17ILzr1LGFeyQ8ALOG5GRjdyFeEvaoFMxb3i2cPr5edRd6kecCExz/4Iw+
NPLbjycnPD52yf57YqFb6a5irPTw7aBtdlkc4cfwsuoNlVUgdpXTvuAQNgB9WwLZpx5FOCgOBbm3
4XmikLKpptMUfk2NPaj8wKDWBrSQKwZsGuDN9XKgDQi3xn6mrL7VLGk4zzKmjuScPQ8+fa8D+86L
5T/sRPKFxAtoNVfZOT3d/dMe1e9cDEzS5leQ0CJyC1w5I1YqM5/nKSdGfWJzlc6s/VYja2uH1vYP
bnRWtDfX+Ov9VDpxMWEK9wFEcXwsysZgjvpLUeADEvrO9eqXgPqkOqcnVzMyLSKNnRSKDl4P4Zuw
J6JJp6UyfDhQQMsIDdRo7U7T5AF/gd/s2TSxrfjoOFkE/cxk8Kl9xXl1hqWvNdM6yK4LNdv06rFq
KrZdfw86swdK3du6nypM54Vzs/MGWCO6kRLS6GYRoUMz7C4PInGCDphppL447Rqp6Y/Bd5nNQqr7
A6DoESByBmDqgIol+90qFbPmfpYU1tuiAJ9om6p0J8mXFXck0tSdvWt99QRF2asv8Brt1HWj1VFJ
i/vFydUzz2liYZPt3kOBIeramWM9hSTYZJ/nUB7iR4ncavARoGIdRxPzFV/RrwYV/hVDlWjT6aYS
Fx6tYmdJDzzzdOjIFEOw1ICbi7MmsdfqrhBhdpA4qYhS1+URFTjpiRzPhIiRt4OymUdnnc5xKo3K
275Owi8cSzLEn4Ff4B6sP6bmApGEtcb/Rk3nMXyaVxoGOAHZasGORzijnxtHAyRl7lG53yQ8UOx5
EWDMQRBDWqGaSXJ+XN2F7/vlVIexxSXXzvCHRqvDSJ+2YK6uB2SzCm0tV9VCdCj+9NLXaLl+yp15
JAgMKkYjxV3xTxbqoV6F97B9oT01+foOxA78QFbEUl39auYdnSOXvYL9Dj/zCmNjn/8wg4Cs/ayx
qOn8uiSGoftknio0jah4unvdpkyAARYcJOMwBTLUU555CKHChiypHzmME4YIayNLC6UWTjAH8Jew
cTFNncMv3/XKrtuecUKo6+/BqX8DXT03H/Z0ZVH7c0RxSSqtNOUEi5qYriV4GmsFq47hosJ0rHnX
YxnV1rQusMV3wNfh9rYwfnueegcZxrx0qg89rMRp8MRyWGJAolkcg0IY5jk3cgGYmtIBu2TuJPso
R5+ALEg8JngqzU/gk4Z+OgxmYxpoucOvV+dQ10o/4Dy0XERyGanjCYhEnF6OlPQYY3PNQvgH9JwW
RpD+vlvYxykk1VzY0qE0l0i1Wm7qRk19iAfaqvTz+NehZp2QoVITlc5/t0QSThPWrm2BvT7sETtC
OqxMNhks0Icr8yw34NR1ZzjQSFLtS0Xc+BsyCR/tVm0Jk+C6FBrXEUKCrgfuhBYuHr/sM6mH4bkQ
zi6YMCKVuj6sh2l5A8xnR4yaP9KtT+/owOicaEb5uoQ4MkmO0lPDTRtgSn9laZP+RAoMwUKtbjWp
egU6Q7Ch3tDjepYArKqrRScaPo+vd/bK2yH1jL9ORvrc96xPJ92Bmku6ETLyrR+agiBdAyljEvUL
rzJ5uTF/9LMU/7Kt5RODfjcEgkEOrBS4eiy9rdysS5w4yXswPM0CP5eCuoNwkjnwvRiqB1vw0Tcy
HwkYluBTw1aP7Yfyt1ZTXMMmLBPVZ92GWwQA3RkuNKv9+5HMNdxp9MSd0SNtV2Cab+Zq8MeybA44
DsqEnxyF+KcnXyNhKGa2+2ffYPG67dd681yFC/9zrSGnT5r+QrWnkuWx7srNfKtv1igSAqXG5smH
F9RgPGNmeYbDlL1F7bcnzPn8HeK1UVYzo2bySX/VFStv3sfTBBW7FwXw7slSGFu4fRqPAs7hO4ks
Mcg36jYEWGWoXlWm/zMx4E5g/MVNrnYwYASuihNXfCu8IO45DYK7V2+ulp7WMePQjGY/UJWWvLUp
mpFoOFcIprMZQy7w1fxEOFxkvIreVK7rHIwc90udMWcMtVTDncV9N/pdTuk0NQenDBtpOpt87oMR
qyyIMdKWUetUD4B4+aOGIcUB9p7HONCGKhNIv13GyHxYJ50PUzenIUwxslPZvZQgYyLRyTM85P4a
ZNtwj2r7om11xz3Ijw1XmlT/eaC3pKCNy40nD06wp3MQ5KWydyGA5mFqAIyHuORymCphZwmAfUfq
CTc/J3OJcLZubwklOL9Ze+HEsYsJWttkrPPqKS880jG0hFzMxto/WkNyefYh73BLGYjliQ0hYQoH
oyFFv7yhY+RnXu4/xFxQjvMLuKa9KvLQwrsqQa1Pwj53u49qDvohEEWvrNviRf69EsQOzEKre0wp
ATWAW5nsMy2WbrFakWoYtfZssWyY1LVYdns7p3nUTZIhMXZO2OFp2YaOKfT7oNRdqfH6g40mmMrc
rjqxzAOm7Q5JZDaaXRl3Ve8W0O6S7FmFYAdd/Q8ZGLjyE6aIy3v7kCS8Cgxb4rEvOCNmlFxgFZ3B
drckrjg+XXxJLX82vVOnK5nlm78XGjas5hP37IsCnfIfB8dQ1I6eFlS+S+vtNxTgSOueZ3AOZBZW
7JgUmAOsRYFBgXOmVTquHzqHxw1Dx1mA6+Is3ao7FgloV5PDzkHrmTB7aGqaCtnvf8RqUQBxqbwd
8H2s4HLPEwe4DAPz+ekaJobfhTrH36kM5zuaGFNgyipRj/NCy8t0ObUfygoIAQL1GsoG8/bU92HT
PvWT2w0vvUc5TPpsZtnx6F4o6/CBKJu5at0rKUzLpSLpfioZwZEKEpj2b9w8MX18LP3NM+dWAs7O
2VotR/w4w1eA/eWTH9Qq/c7Otq2/MiC3caDt0X0mrppQrS62WZbPMrB93TMoaH40BX1rqbsOqx+V
kSRDDySiJQBqddBw08jVQ+Vf//6yQo4sFyvmz32E/sZxgrlytV+V+u69gP/cZZmFHmrGDTLV3hHP
VlSnJSaY0RV04UcQJFSju3VW3B/WinjXmLGiz0CKReKp/FcvsiAJBbqIBvVNuSqNE5YQKYnspl7u
qkgciyxqCiw7DuTzz0M4yO3G9YETrAt9rZ2lPPOG5x3vLvyS60xi8NG9VoyvYQ1sybcS7csbTvQL
HEqmHvym0bk8xl4GFbGBoDDQhoYopw4EipdDnlrYk8CRG3ZDri6wtdhAgvr6UWJrvM38egRHnBZE
xilJYrw9ymZNnnKaGf25vG2cMbgv/V6K7W5+KgG2kUneSXcrGTI2ZRIa264U5xKrXeHshCDLP7kC
dJWzK6Zh72iFCT1oGIEespLx8A0WYfBFsXD7HqUKTW/QRvhNpQK5rPSIDjr95VN0/1ZLbfdXgCGt
1uaT86o7W47Q78fnaxxh3OxrY2b0z9SFj8EZUkOgD7+BGL/398hoPON0OUSZLMECac9GZ749LuIL
RRQdW11OJmzjBlPsE1ENdzQz8NI9a2E+l+xgEa/P01RYTa35HqrwamRhx2vWC8ZnO3d0qBPnFPoS
2NX33BI54xYZYMDQtgEF+5uVQ8Gvy2PnbEXlQMUjOXFbuXjyrYY/JIB845YqRk20qeamCNz1lzt7
dvQYjThO21zF7LQgnDqhAXECpNcYVMDDamN5GEJVLpFcR81n/gKdmZ3rX1ykRYDxtbcv/s8cH+zx
bZmsxDhb3iPzKThPkvKfI2XsKqbhkuM1RvZJ3XOMCfxWGdc70N+PwZJl+BG/a9QkBDqOB6Lj5RJM
aXeFEZTEr9MG+/HrFy1hkqDf6VT+d5WIh8FgXPmh2o1CFj/SUUV+v/XF7Cfdu8+N4pZmo0j/WXkv
RKF5eRQvkOTxZSqpjj7J96GMCu8VWNwV3un+fdfnXcDm5Yphs79yS8G3wNVmpNV/FP512dfu1tKJ
jIwGK0PDOIY7NvlvRARihS6ftmm8LkyFUf5dwq79ExmpuWoq68MtUuSNFE3fs9VOLNTl6eCSqOsj
CVGHr4GfQZ+jBIh+253WQIcHBE2Oca8n2PB39mnyRTp1UKQpblKpihLUQbgbgHr8RqOFDrihk3bu
q1UpHj03MMi0/6WQT0oZyhg1JXRroYmorrtIrdpbvc3lyqK5xHp2ZDipKruffJe2t8zg74JHoXmx
qHyDd6mhufPNrlbxunvuEfqp/Zzdings6dQiws7ZTCLf+w1pn3jsoRt2RNSTheeZaBjVpYOl3zJ/
AQrcEhmJRVcOJL8AvJD3HBnBDN8CbWn/UaQE91jVJGaj9rkbZzYKdVqqhsC3eS5UbsvPaJqd9ndR
x1R3SF4kjNNfwzeQIcekoGGtUPLv8LqNiaTwXfiiOWxbgNSE8h7SfpQkEBh1Q++oqVJVCcwukFI3
H6aUPl/eRt9sUu7EFVU5BZ579RyEzbWTCDyrXeylCi8z1rEZeJ9gM6W/L8nNvo5mHy+cLG9wIq01
fBImRxMyoyZhFuiRqmBzN0yQkveQn88h1UMEWBsupmNR2TzeH5v/Rwua+cR1jTHNVBlaCadTPKDo
51rN3iVw1vmvtY9nQl6KV305HfkfGqB+IpJHDSfXrLlbVoIcZOhxSemZP/X6tE2CE84zTxEHcdp2
xU6nPw9t4VTYKtMEQZddZ+GZRglRYG3Arfo1ZyBq5w1a6y+DAVlA4oaK76Ny01D60KA4m7Mvpox9
e6B3pU6zVzacIqm82ZAKpKCte124K+HrbBZaEvkR83xbejRy6J1ApdJUtkS7sRweJEjBQNgGRmdG
8yIHulAYUjXWOEf7rk3pvclGNasHYFqz0JKJIQfxDvPigAsr4stq33jsFbE9d7XimGYLPFELrohu
JPYyvrB83n613JE86OIpf8zqpF36HF98kMbgwqiDqf93HSacSTETqRuk8sbc3lVvaxCerFL1fDBs
klzwT4P5bmGIGOVv7xrMvZIWgKCMKjtLdUq0AzRtrVsNetXPyreJewL9BqGA/iKcqM4rGW+nq5IG
QjUCkeOfvpgfmAkFlo4bkOaBYjYJjkU4G3G6likOXQEZZUCPOwB018Dwlo/qsE5YhXWobdbMNeCb
ZXOAmvQygyXvZDnZBD1FRJ/UrhedzDCexX9kjHAPnDUwN9QI3lLGSmIQbQ3fIFgWmCT47YsU+Ho6
ZWq3VDjZzYKcVR2Kvrsph75JDkUL7CMIXAAJae/oCQOyHWkOveLSkRUsiYFpX6ig0mftbDLjOmqK
FhZKVutTAlzizeLiojdS9pWUxiLTs1i0O9Hc86tk61MHzQuSqAmq3t74Gv1ctY7WxAIHOu6S14mR
+YiTMXk2t1IIWjhiaYjPOJ3ENsSK2Ao8CcjyQpMOCob09E0tOKVnScuwW6ygg+htvJ2N8NG9Lv2z
xsy3RQbXMHtBSE8Vr3oZ2PJK+x521kWy8lFkKVJXOgpKhl2hLT83Akx7AutgN87M9a0juMf6CBlS
jD67wtOQHDrOA3z9yrzFbRcHedEKw/B1soddOZ4aPHKT5oj37A1YhlFL1cCXQsz6Md32yrvoTawv
pLnLQXGt8+pt4bS7V61I1l2RJ1HIGDNlbG7t/0baFXhCN36V5+xJUUNetNalcJIxeRWBaxBB+UeN
xFvRVGwg+LDs5LtnHnD3B3MjXfCk7W2qkykGJwSqvZUo0mVPy2953ecSh8GU8Etwydt1YVqQuFiA
tWTre17a8AZedV8TlVcrk6ZyPy5o3rGrEAJENiqhBWjUE3YtzTiKEwGd/Y8mhXcxLlEKmg901l+P
8a3ZNPw2xmJ5exLHVwxPN6R5tOPodcqGIt2I2fW5A1r5u93ayt+GZsdt6FiUZeSRTDWhTb1MBpwj
BDZX80ldtd6A2rwzHlMadIXbcIDtnslmRV6oNumwiY7xRfoWCjbL1qUcbrT8juS2azifsNtsML1N
byvIdRqYpjyUGWm7NHb55aUJcSAw3OhQ1HovyvIsEGKwNfr7xwYOfp2mkW9F9Ql1TlCxdXpnMDP9
zxDZXnBd6XENfsHWnodAwiKcA4wUtmLaOTDxT5yzkTrftb41OfsHA7HqdHF+9pH+IjzReCqO8fix
ZrjImq8BfU1Zv1H6e9U3qah9r+ZRf5m740+dQmqu5IxqbNUpIN5JFRllCh5C7GLgpXL/P4Jk2MV8
k92i3qbIeaxUFAFnr6D/0pQCO/xvu5dPAWzfKuxA1l8dS7GO96Hyj9WpE1/AmVFay/jGTwK/gBYG
OcsQ1mXOCC3KWgdaACyd3mC1BlZFi3zX37AXG/9X1TjkTZacoXJp3OxmTA+OzH8RocUC6i39x8u0
BwqpbQVR0zFpoUa4NlXA8SChzj9YujdjKX8lPalQNliavOt/UPxTRFuwC9kEioTNo5VmVX+eWYOf
uiWn8ni+a15SzsThjaj/OekX8PQf5qFhaL7WtGabnopQasWPNslIbfsBXLMfg9whaaQ3hLpgDFl1
G7IfGx3k0TmhoXkBi4Jobq1cf66pDWM01JM4tWmmfkYb6YGDq/bV7uN6FIG2dG96Sw5tBmo36D/c
ziVjxro2RPtF+6He3MGVEhPU3gGGe/anBi15TIJxH6SITGOS7D9O7iMICcuP67HUZaxiKT0TBF6b
wssSKmFuKGff/yO2Qo6YUbR1Ue/deKFnmu/upo//gD89yynU97K3BKtntMZX/xlYczQc3caDr0o0
4MhsLpDd7cnF/GqZKPFOJ+TksjZ6gORfX9evME8ifZ3zFbg2hdgTL+8Xn8srtNXcl5yiZPD/IByX
2V0DhPrIizOAYRT6xsAYJ462IYpnQoxtsEFXFxb7xqlJESB+SIiF8dXdub+2UJ/4+Y18bRNe7h2Y
mLa/wGzaWHGAwccu0VtCCsQ+84smj+BwTKlw9vGTiedXD5S4b6caf7qjdopi8b3Z1ylnJcc54XJh
QmzjS3Mry5g/DgNE3aBdyu0mkxkXb/E85ccKsFXT5aiEtK1lS8NKBIJc0yMGlcY87/e5Od2fVI88
1b5tR061Nud4LBNKEw/cwWaX0Poe3RPVQ6Q2u+WoY0M5xtwyivK8dSz0fiLoGpS2kepTJdcyhAXJ
3+rLlctGb1XHD5UAJrh+klp296MEE+SupUvvIY2jYL3z/zWNjzgvo1hA8InEi0JSg6PsfGJhppVu
dZu1IFPa6ZWbebWW/sKsZYyFHjPx4/FM6jJOTbqTaqi0DDCYAHWpslmpr47jiVMAVhohd3cc5xic
zGnbAZdzz5mYOKecfgP7PkQyFZp3B/ROPj/8EOYJCda4NxGbsVPOPlWJjZnTbN5zCOBj++XA1FTi
K1VZ9lRq4s7JxmFHO60nx5YXEl2dBjvkbix0XVC6J3aDcOXH8Qp5SGNMzJZ5htKTlXOfzqzW2fgn
XgQWBH3txtUObG/Tstm9IDQJXX55kSKoex8ZUmdA8ukgdLUz0YBHB4gfxTKzQeZ5a7cbXV6o61Rw
mA1nHK24NVkX0E6ounhTwQT8lBxBwmphQ3F3OKSbIwjWtEocrDui1TOThG0cFf+DNFkAW4MH9C2H
MSlS8/6K35u6JDKC4kLCOJR4pp7uSTGkfzDxV5C0lZEd+naRNVvdnsQ88BibIi55xA6eL4johy8G
lnElPKn39zxtsCIFDs8OOCzH2+2RUk8TV55IvRdb9iENsuYjzwaLYFLos6sDKQo0MgI9t2/alA3g
OvY/BY4ZQzSbq4IopNrFAhlw+AxFcLtBceSb57sH85Z6Edil6n/N39djSxspApDY6r8xr68ZzJVx
3ve+DuyTgZEwpTfB+W/BxlZu3Gknb5+Vo1VP1TzgP6cI59YGltfMNnPSGwI869BaN9iNy9eCiJSF
dFlGFLbLyFfxYF7TvVvZFVX1IOJlLvH9LEJQHiwZsjHkAszazWfDF5eryb8DznlhYtaOmQ+hTw3H
RlD4hn4OXwVD/yTvfHRsEF6kcindhS2IptSqWox0nj3rCAy/RA3a/92umH2VATc9zBb5mzuJvRlt
SP+XYdN/nPha2z0Wj2rmU7/zHOQrWnbIrOQEKPFuZTPysiAE6gIR+qMvJhjcHAVMj7yo8RYgDKr9
q2urFQ04aCosXIwoiHm+07zaKQ7RHU6LJh9mPfiRYuGGpiRjmSds8YS5eCMyFNkj1X8Jltg1dBaB
8ClgD24y35bR78HTM+uhGBjSisxeznR22jxn1GD9fq5dHw6cu6QdCzpItgcQaCNfRdJZt2qTaAmY
5st6OlDWH7yffA3bzZLsy5nM3bbRCLHsOpxfX/cZqaZBGwx03pZOkF/hhTkcgfVUN0ZhH90GF26o
GYVdiLnw2gdCEs83TP6bfgO5M01daPS1aB89joMbTSjrYTW+sr+jtd8VOGITyX/M7qz8iD3vUk9p
GngOWjG3T1BEmRCGg7HJKgSf9j/Sdhgz8lz3lB5BMD4m+zY/5OMEjQIOrV4nxddN0YUf64DoeIe+
3+L9t7BBVxwbWKKJ3bcFP2nWQQ7B7hzFL06tg9bMV1jl28cWMLK9XgBRsaYrVar+EHLIIxN00rxK
FAO5lhEB1pzXmF27njq+Cy8TiJR6leOnzDkNNLWszAHvwEphrOPTKfxep0TQvs/TI1nq2ZcGPtd6
0UZg5WR+FJfVQnon8Kxl9MlWOpydyW5OCR95mild9V3pLZyvIuUBUXpNiGaV5lGtxwFPwaMyukvb
pWhRFjMf1ojij1FQfs6PxCiNMWN8mWFPHA86TIeLK74UYbPUfY0adQuoclWeJoGRoFq9lsIVkO5X
f3Oql0hvaaQuIQKaqVZSCPJnFEEs8xoeKNYJMCcIR8WyZoohLZEobUaUw3SAI7L35tEyGB3LeKQs
06cw60B9EJae6KD8BJjk0l4xeLWiuikcLzJ+Rdmro8aW/oJEkmzaejZQsJHaHXOVQn8ztwZm1naZ
feyvxRepBmUp5YpGgZtWkfjVfx4WQ3H3NDrQSGrTxjO65m2J+XepwIcoasummKvbtVxTulcd9d8B
WnlFk037CUCO9unSZtSBpvq3XxXY2obpK977VDHGBA0XEr1QyUOBUAu6u4Vxdps1BZJ4+YFrxcrP
pDhS2U/cHmyDrLG2gXiuR2fODAdrR2vrrdsyZf74EFA5T+BLsQZuZlBSZw89HftOXrm7/8vAM/e7
M0Fdtd3+ff1CxV+zgBflZsnwryNPomWDegZ6vSQjx2LfpDXxXKRmQc7kuVoSp3eGzqseuTm73QXn
DZ9NhavVh6cblvVJwEcUqvDrWw/O5N4crNa0gta9cVhyiktHlZA6HHrfSnzuKd7SVvxsmzMlJuVv
UTGHh7WuPRk2aauO6AEA8VeyyuiGh1oewYy+ELXTx++NFe6wkQVBwS9QoemmzuApj12ELc7XCqd8
IbkipGxW/auFJTSxxRZF+RlyzhtCFEBDkQ+PAlnAQKczhtOSt9Ny+3QAq8ak5/54m91K8bNvxpcY
ERVTOYz92WwasxFuiB6rGizt5G+tgkGuYrCHgDNbQ6rytSl5USrbvg3yfw9VvETM/KnmotMvXI7K
+gv9mAVJc5xxMUOVVBti900/Au0vqVIl030inLBkIPID0SxyNvMUDicgt6VGNaBgtRq5pyVaHd8n
bEcTDop1Zs4RIn4xUJeKFHf6nPcLq9Bvx3ap5pcijfF/UYTIokB0jp9X6ruFYywfu6CDAZlfHmNA
lvxEA1xTewjSr6XpeYSX5e59GegYHejSkPTWkHeXCXImzNqwNFfXbnqIL3NUG84u91RvdJHmi9ne
ydSRlCGAEwOpGHOG1TV/znmLEmZle4dv2hCtU3LP9X42YfZNwhuy+OTZhLOlVaMKrXN1vz1+qQrv
A+NKtJNBM3Z7/yHStxGMilDWr55auus/GwUMSqxwxZTMalDDuTvk0b+nYiXaRAKPVgupkHJkgE7B
S0yjZhRKLrtRQuhKezNqlxNNWvhA7zgwGbq18G0ld/o3PficespSgiFtzzCGCQAqp/5MjZ0RJNzP
KnPm+2wYhoj8BNJ6eu95MEuqsQli3mdaSISAOr+nOKL1MF+ChBxOeIhFwCso5SIEI3rzrQAlzHJE
JDEROSrrJ6wXUlweZIK3dF0dQlGvTVTbdtciPgIZ4/KTAnfLpGNzcyOEdiAVNJgNup6kJRPONRXw
hE5mv3blr//CT4/uMWlpB4i6HJWk4N2Nibbjyo2oyWTys8uLVJmvnlN3/AsM+N6outuzWInDbILG
KUuNP3iwoyIP2ccNPsHoT9QR4frjlYBsZeXZiGwO8uTHYRbvoKf8Zn0ce63S5j1qO3J0BOd43xv4
fjqsm0bMO/weHlMpaSI9AbjTX+fD1T785jGAue/cjvp+yoYeYs6pSz7ydGAWnQTo4HbvG5tH6nvq
K0ndBNRJnYlGqoVIM1MkIR2x4QI9WngJldOkP+ge4OCXEFjaixKIbRvwN50VMwWygMKrl3LvNR/i
GDIkqFAXVUeER9urTMBQvuTr5tehKHeoh7H1tq/QQKB7HPy7iX5QWadcrYD1eCfnFAplaiCv5iHI
uVAIIMGsRv5KedSa4Tz6dt0reyOt/mr4aQck+qTo3vsxXbe8+yKN/xshyuxcTM2PWn46tM88PmzP
bWQZJ0i0UtDLYOaaa878p2g24JhWk2KbCzyNTYnTG+k/yBxh07UcORb2qZlmYfU+05+3SyspGhXF
CpN58GBUG0upk9GF8Tu5JSA3jFvHJbxUw2dCXZe7Rkg9fIpr1zcjDxoR7KzOShAh4YCi3YWXXo5L
NmFbGq0agVmWIHs2AeTchXt9D03Xl6BT5w2GOVteUamISf9ZVGi+nILcX9vbMYB+ztLStPJir16F
tYm/mfhsJIDSbD7Mam+pPn9kzwmoZJoWaHEu6Y6Hh561fjxxeQK8K216duy21xRkMXKOOGUsiYRU
LFHOzu/joa78DP0E/Awg6PojPVH4/xM89A4wfcNtjK9x5fjXe1u6iJGWrTSCoP9DR6IwK9pJtfz0
pjKFrLsHO4XkC697izaAcELdBWo9sVQi+kZP+pM6MqqlZ7MKKWPNAo30KTK4elcQ0pF8o+TIztFE
Q353a+ZLF6bhb8MYwemyr39IQJqoSe8+ofVk85yx846oQwbcJzonVe+PEDYLMShweTxxah8mTDyt
E27tiycNSCtXgek4qmf5addj19qtNgSdmDeniTah3rs+Ague14yEDRddODkkBffbZc42HD+jw/Ni
R3D8izpQqP6jUsT8jjnZmhJKlQjekLljy/innUvUm3w15qQ81YJOgHVb7dF30JMxqCJEYQu6E7wP
vFkSYLmyTHDi8E9ImD7yEt6VGkz78MwqqsadFKxmooulfzErf9PjyOkt+xLpXVJ2o42KmREpSUi8
peXmZGABYewF1EyoxxCcPsCoCby5EbJr56SwqisU5FfyUqCLlyZicCfsUvjOy/mKBH+JVfdAli7H
WL9JYQoL+2ZORKRnUlyijUBve/oJfZrPOOyNkfaZb2BI8gQkzymYQiLazQqfhlXDrfQIRy3daS8N
Adx7TmFy6RxxPDRghZ/Iro4z0lQEjBuxlzuSzVhS/1+qIkWOnonWqlll+UXlGl8Wu/Y5rRdQSlQf
YIvrEQD2CzABU145iJqrYs+KXvArHj1tNOtyYAycjzjROSU6nYkG6FGwZ8bHtBnplItzYPEQrhPl
fwL70PQHDcjwHRtEFtBqxwF7cb5KrzYtDFiu3/1xOWw8jC8Wf2LpXTQZdIW8FhvF77VaSUvHSs0q
TrsMWjGukO6OR+e2cN5lpd8DfYPB6deG3RZtaAgfxB0fbCPN8JPhYbjQLDhbg1qPJMiimTqgpPNr
GsOgARTuE7ad+vyXn/In3L7w4z/DOh+nLeQZkObUqdgC9kP77v7HvOie6KiuHac9AGNTlvIIV8OK
tEHO5uhdc3GNJ87YxEOna/q9o9H5gzJ6LdeDaALjugTqiTY6ZbGhynjtNK7TnNTv6vzv5rqR8+lF
QDTPJSx7TxnUGuool2VeCtJbJ+G7TGmTYuKbceVcGf6ipYfebkw/ftm+P2yn+OIwllcAVLb4gIWq
WJUzbGBuajJpBxMLhgi8xFeKLw+XXKSamOF3+uX7ZWnW6EwnmGewzNfUuMvBcwSMul9JRiwOyCx7
9sN3ldzJ1PDGGyPTeho5elNOl7Az0CDqfMSnUBQqK8xTtv/4oLYuMat4UO1BjYt2vYE4O4Bj04RT
wt6rfJFApq5RsG9veruIkEsh+5VXcSdy4MndhAzEV95LCrf/XIK6t7LP7uyovUZIQ5geUVp9zvum
rjZVxOC9AkaOkubsf3sl0EDnrZIBtb8X14zlgaxPsuWKl6h2iJuP3MteZbb8NwlrGIh9+stnSQHd
y6XwJJNfT9nrSKKs4+LdfHfypgHCBZEgWa9FrgSdjoddiEjoBsGmacWhDhzBOeC1esu9lrSjFr3L
4cMycb6mrJ2hq98FPhMpNxawZLBjZ24pQfvi60pqZJZo3dGT9XJwAQ9j3t0EQo9vNlTmIXeHN3BH
6meShRjJhku/q06lapy6NNTCNi1pwifKnG6ZZvpWfTJPbcSG6inknLpHSlZ0ZlluDN3wW0QmYCSH
oKMTwtf5nlzUPkKrChXoWpN1YSZr9v9Ut6q6cu5tlfZW4Cz3WcEtkPSNArET0vWB7jmgtvldO4Z1
b9fGKQZTwKfqUr5G5rXAHBIhmVXlmHd3ZHv/DzMYcXg56DL+PoA1azsOkNU62BL/mewGjDsBOi+Z
Rc6TJUboyJPE3ms23KPGcrP+NM2h5/hXzKC0vNH5e0lx9hAVVI4eD3Dr0fsaCkqHOxmn/vFVMdSB
Vw2A32rqdh8smNo/T3g3qmvqwhJoADPRYIMDsts2jbOkZ9OOlnRdIxx4mePwq6h3IKflaqQs7Ayl
LF89wjL8BWs0VK0HZfTyTj84yUVSTX2AKqclSsZGG+KRBag/mxrqyDWZzRgV2AMw0mgFRvzbRXEG
ZxJc/YUZYsYW4SgECgr/qZx3tWXyFcgFnQ+5VVQOnMkPueuqaL91tXvPMcZi2pKfnUo4CZelgnVq
sTZtS9eOoc7l434EVd7WQWj/Tf9BFKDIixmaEQrMINesxUEKnGtlrn4P8bDbdekepJ4Gb2CcxKX9
OoKeQJrPt95eF3br0ycO6kPYyUFtsR/FADU0H/Pk5lgE4uFtAtgGOpmxOvMZmOTSsdLBSzZMQ+jn
jlE51Mdz+cMW1Vc7iQjvaitUbV1mZo70ItGQ7CYVl6S4wbOSsnN7blkSrQdYMbFtiS5PhdvAaJiE
38J1t9+Fky2Nu9zeXSN+JmDVCMhAGrPBNXdZ+UP/ywThMQRNjooBHphMSIgsgu3XKcpa73VhAvoz
mixe86ToAbhmB7OMghz1vlUES2R4rJrAOoDWea8A2HMrMeHipTduKRADMLsbSq5kNBFXpzI6QmNH
1dSvaBsvlwSTVg/pxETF0Y7NhwOON1bnLF+DAjWm/PNjL0/OWvDip7r3w2zLu/n332DtOgmLvLWg
AeroErLwuTYsckPCIAtL3R0smmmv8EQLSiHH1dETmyolfyzC95yaTEZ8IotL4PBx+KTVCgLXyJI5
YFGEfGOZaj2IIHof7F8FZbNE9oBvZgbWFDZR6ZTtEFP2KLJRsf1VtNuH5fWpbSWBOxztxkgBZhzx
OKSF0RMucHtE3CRg7U3Kx+Lo2sfvjnla9O3Z02uwr7OEa8ZzBpxezyTe2UD5+doLNsOTEkd01p4j
gzuO/T8ROGOMwkSVlO1+HysZ/IOAlq/CRvIZGhwL8sGYns+iJY7N71z3io7sekEHYGjcJchrXbUt
SHrfcsE7+8AlF5ogM7yyfO9trvVr6npVG5thnhNYciu+U4D5Ubjg8bVaKzz4Bem3E3yfwk9rWm47
aLF8zP4B6cJKPmbWYhVAiY6xl4NoqRPDRHB073jDE1vLFjPNpMe8DBvKXyakECvI8/KNbe+oyfuc
b8vWkky2ong1eQ6M7e1/EDyCLzEE3BgWpaGwBc2TLBa4hL8CMq71TPiVvxT093FQqbt2L4cJ0GbP
o4jtnMLLfDeCV28HsgTPxKgJpD41P3FwTglJ/CSwOni/RkoDr8EWIww/nDACpevlW7fyPsspR+vT
w+DybouAe3Xk+KiXa32VuPvGcGuyIqCAovTYvr5TB3Q34R4s56W68Ip6seXWqWExQphjp9BZQeSy
srPKnVlD9bnpIXsNSbXlqh8Z1MvirNsaJCnm0J+Vpge5BRPWVA/FBTQcuKo+oYt2lRK/3gMssGeM
Hv9U5NRUazDQn3di1jZK4UUejhd0HVsIbwdOlDVyLnWGCoAJM8REdWJYR+38DTxwbTjAIQdsVLiH
lN88jBmSCBzQTbOiYthfzZ8kU3BG8PLz4zm7hd5MQFc9AqffEp9/Wu2VpG+ATT2rgVLgkIe6VtKb
gJ7VhOnRLz4JabQLtmlQB5C4W6KxTTTm826rZvZGY7YpWESXPd/XXVquTutV0E5veo7OvABVT0VV
NH65aQvzpJ3ip0B9A0IjwHtCvjhPDBLQRBkwQUXzhxJTU/vvANt3cs4xUcpf2gYdiqfnGfsyBr9t
27IAsKpFGenOOUKvyPXzfLyIZeYpVAkKNeoBWQnTbIczBY1Asd7jfUuS6YPmk0OVjTM+kTdbDozY
vRTuAgG6WOwocTjnl0f+Kr8Rpqm9uvuUagH1YkMWALywXm5JKEaSEsQEbaoudQW0xGUqbU0JuV8H
FrTV9sF8TrR/lihEaMAEhttXQUZ9kdDJiFRT4v8ANhBP3u89Pb0f1MlM/Sejyd7BkrKPLWKa8/0L
/LuzjL+9tGJT7AfCTdNWFGTvxT1DCOMVcMJpGcC1+bdDRuUu2QwaQ5LAsM+lPRo9FufjX5QyOqgt
CC0HdWzx42aycw6AXuPC5lBD9vnPUcz7Wi4rhVGtv/Bp4FXLe0Ex8mvSwlefXsNlFSa68mSzzrqe
Uzo/S4WISF5EJfZksr/ntLPHGknOwodGyXcbWWrchRyb54b/a4ZR07uH3PgnA09brZILmtmsoX6A
GVaReH7jLIhthq3GZVwplgsDZXF3R9ifRgccHJm1OouNxKCgCsHYzdzDIIyFU4uxDv2tpagToFn5
0YCCHUjMOQ5v1steRMLkFhdAn62VKGlX0hsq0Wk3vaFd3TPlbUDUatdC/cjwa7dfJp6KF/SezYFf
/CfZ7tfM34foYGY8wbN3tWYQqL73CaLwTEZb+ifbJav/ZqFZinSMu7DjSwkPrb4Ib+EZOrSYYGaw
MOCEUgJtwjM2okXR4ABw03PZfGmF6tp/AyF6L1lTq0UCeC5bZx8Wb4CiCIc0bMURxoAVZSkfcSth
/6L2HtE+9zYDXhm+vZ6xPnnKg3QtmnC+HPZ1DdaKt8+rlc2ouy5Dp8DZznJew2XVliMP42kf6nkE
jCR89rGXVMpUpxqndUXcMYn9J5lP9YMN1Uxr0Wwb2F/CH7IqQ0UBzLXBK1HG4C/dHTaHOanHyaNF
JU8MCcW7WTLf9h81zkARCL4oqFZlfiiklkXr8M9nOGkYXAl26lj8bjYLNc/cQJIkrSZhZb6CoILO
/1KAWpJtE78YMVx3jFafYYuYNhIbV/Is9sGP34vPCAlejCv3DTt9u2WCrW4dq8Re7DLujieKvEJB
ESn3UrkMbemr1sfYHOJhww+5TJrkoKeor1JmczpdT3X9D6j9TACpIDh7KefjZNw2AWVat0OLGQYc
+6qL1s4SypNr4nq4zj2A4gRRNkQYIb0HcFVdVnA41hGjRSd/i73wymZwsPDsVqP56cwCUCxlTmRG
UbyffcYpLzzEq6j1KUzUoSG3ag04tGONbbC5NeZ+bX0aC75EMCah15xEdghtEfDUO08JZhuX/K8F
hn51thWGFZr/UtO2vWJ+K31/o1Fn27zDVkNir5rPWNkfF01cM+VwzZLG3Bf0GgZx4qKFDZCM3KXK
kb9FLgN9ugRTJ9I0WI9y0/equp2OHQN01VJv2uFqJX5xbOjuU4gjt2hd2KLjA9qMVnQAdMHeaSVN
yC5V849GQQ4v5MWVVWAY5xnPqn7mTaeL+nlpMGM+g3M4GywKMKkrxC6m2+a3d3hWEHmVAeMZR4Xs
PmpgvinF+mKg5CI3Jt/nxOft5b7zvelsyfphof5TNRBpQpWh+384WoSagnLi/qWrSkQg9DG74OAn
CUBiP2uFAXDCZp84szfYG/ergomSe2zOulGKiAwWmfbOEmLmX4DIb+T1QuA0x2cWJlSg9nB+wqf8
+cUKBFJkGuliUTy2KkGb2b/9hNfq8NekxgG7tGD7VFU/Kj0m8Bl0GDe7izlG1ENSCJXzoOfCQ/7e
moWmlWHLtPnX9BKTD0Zet8xaVaLuvAW/RzuUi96uetH9e8IeJOrfvMgK7K1UwXhSS4LfwK4/z/AM
O7yb6keIEnqlOV7F/oq3rVUcJBrTr/mdA6+uq48mcY2JujD8cAV7IInGuRZ9lk3wbDAiIP0uvUQK
yQ5BY3uNnYw3GvYdcqmnO7rtCC1hv7IUlmKlp9kBk5PIUKpW2WF/vqhc9+EY63Ay03BrxS1+g3/h
U3aPrxZNl4sjeK2U8QlTh2wgXY6XvEXBcWCmD4iSaFH89v6+BCp8QG9PPEv0I5JL/NSEwce70TVC
5gAANCvm3PxxAljWusnmCspfIn8iG8Kx6vLdMFKbc235n4EJ8+BjaDViVsLaJYX+16TURBUjiqgv
G6g+TbF70R3HlhpZgRibAO0pRjR+X1mu+NXIMwjah+HLnBSf/ZmFsgZyDJEhP88UNHALI119ZCQL
e2nTDSvv3HB043zDj5cHw8wzC/yp9WeAQPOwdOJwGYciSCC9S5caSfBUFPsfxuxWGrm9P6vPp/0+
GO3G8dBl8dja4+WSpNMg+tkDsU7iN3IbKgyNkBjDmhnqdef3/NdlITAMVW3ZKNe8z5NwgAb4aM03
1nTudmGzmzSi7VAjPMZdbFHddVZNr3Laq7WjvftN63DPWfTUfcU1GabppQvFI+6c4RGvQbM9/vJK
ewpIk01vLWjsK4Ny4yqma1MQlUs9VrKyV5/ZbU+NdjrTlFpgbjXWFY8iGc+odw2VS/i4oF02v0Zp
rewKEM14qc5THoQs9R5oct6qT+UwqpX6OXkwt2vQbnm8NOU9DT1xoHonYaCDp31ifZ0DfHdIhY7Y
BF60jueDVU9hrqFl1ZOWhdZHWaR45gt29eiioWcje5gTrRu+W9J0JZCYV14b/BFroXg5LT6qQzwU
DsFYJeKrebwH7KYgw4pTAzJHMl6VPML8xbY5DX0M86Z34+oQDM0tdJxYYsz+zSFmk/K5XFobldbu
j+aV7LXE9gK9gSdiC+aJwHx5YnqqObsdzjeUiBpPLwLiWmvEpFb5SqFmprvJtDIfxKaqqikmSLle
G7PQ0qiQjZUzlcAlRgHNkBJMMcoz5G1bt4YSB/m1F69voKee0oAl6shIg+QXDNBFMbZz+/nZMLso
CIGMPT6M/jA7oBzso8h8YOEq1vbDMbEvitM7H3oravd/VBlhbUDDDLesdZweXIsOZG2fn4VyBS9G
u4nxTpQHMeKaOWdhHnhJ4ClRI/EqoJVV5+DWMt3AAZq7IyZ4MPsuy7zKhu/YPuawR5kuKzsgnmuS
NYq7jmxAcesXI0n8cdftk05b/AEtnwSJMF9L/CX/Z305J2WHaF8tKmAK6SSixPgulA/4z/iB0YI7
gtYbzGTB/i7taPTrrNnUvuodXvMhYooQwlNzIRdCzv0rxWQZ5eoBm22mqhMLu0Fc+mcFEndTRh8k
XIr8rQTsEZA7aWvmwfLCO8q73+1ODL91AbXs8JSIa8Yo0sGlLKVATPf5pgVaHSpzZwYcmiq97rIX
T/VGcc8EljHAo+ihxDeyGexov57azPvxBrXmoOdPpB6CDYePbI+Ef7UfiBijOYw8U3RiHxIJX7M0
CDrjIYI2h8sSWTdHyyGWspoB+sqMpK4FrC6oLGz3DBOXNUkfPOnqkLOvJzIl72wuK++spIDfAmhh
+951kqGQmpGzuyNBBmk8gKtRp2Jo3BgneHxyTfnf5abnAIKhua8plHlBoZboXq71Wq+0yP7hPuvB
4VXMJIl81jUzSlkKvnrnGl3dT5SeJ0yia4jYCLWMF8i1fPaF8PuSPATatVYJinjqaYN74GIzvZqQ
c0ck45Wi3WiyFEPj3sjSSyVqDUhXGX053J+tIdfol7oTeyaeoZ0gociZsp0QMLwDYpcSdAXqkrRU
rNwrsxQTli7hpGVS7STi0AjyUerlFmkLl2QrDkd+DvKKxU5y9MwS4QHt9tmpJlUlhgGdoVo2jgJZ
5BJgPZ9iN2lxuxBr8IJaImJWwdz6be5Wg4edSz7fvawfzLdQi0Xh8WycdJjIZKDXljNJqwPMAgFk
U3klTJOYaShtTeO6Kf3FkNHVt5oDVFV812moq+8/S3KOZl+f1UQtHNTKNxmCBgnRxSTbigqTePBS
zAmQXqhf0FqATyaSUqJHan10DHV812hCCfY31BKKEbTA5Ky44nvSEwkHMHNGa1a93I2P1IeGN/DO
ofidDkOi33TqydJKUKWVfNQCA/dlrrIpw4A1TqWxENAscaSudanQrG8ML/qN8tZL/5kLEYiq2qQs
sfuiLhRVsJeXBLnUAy6rja1ann6Lk2jiDVm3tWNug6/r+afrnR31KTopTQYXOoXBEnGsZ7EjLySP
dbR4sdZru3+sMCBc7uw4uLrfcvFyyFPGTSKWalTqd34Aj7Mh+rsbWnN28PrWFhYkBhAHTTV8V7sR
GAeHykbsGnsPF0R+f+hjbLfg1fXfwI6/4lXbspuHQzx0F08bR2R/mJrVgy2vBQ2Lmol1hoo1c+3m
CZxrZqGvdjbYqWy90+H9josNcACmRPUi6+SzO5ztzGXGT2M9o9x3IT+C/0qoHKbrgZdRHRYMQha3
/fkzAFxDHoOZ4rQdUWtyX4zJ8Dp0rAdJX6TEBeulX0bhRk5YADRxDLPrW3ld+VXdCl0gqlGJIvuL
gHTEilz7jR18Vsnx6DPEg4W63hGOlQGeez95nNPecZKErpO7bSuCoZ/RoodI5m+M0fEc6WLXe5e6
eij+KhVXi2PQgFBAFEwQyVBbOmBvmxLRTPXy6y4Kon0cjsNqkhGeViPNliM08bd4qjr0JV5hP60U
e5Bb5zddISVTKUPGZK8gkf09XKkTgTJL/1+vPl4mjwPus8Ulu1meOcxP0WE9yC76jBBKXVBF1cx1
5lAG8Nfn7UpV77sa77ikYpXF8xhLWilpYZsqe9RBIMhXnsOAIyHqRhWzhk/X7VnV84OM18W28PNX
6ZytCe8gOxnHKeoMBre5XIe3DtzWXXz1PrMNXhSp/iS7AWMXNvt7O7ypFT1zmANU19R0B2LIoMNu
TtcXKiATVP/HaOXAPLyIoRQIYkSm+mNg0EJJw5t+nC9BzwK+TGNssXx0Ax5R/MoJb3C8v81Orsrx
Cl8rfTIjxi+609d4mokivr8aEPLjC2ZBuj301spC6f66bt/eUb/eHv9jyo1o1WOT24Cyk7XQ9wWE
H1N9Itdty3he6VbAA9oeJcyAkYx04AzKPcUnpyEQXhCQWnmDJbjO+nuW2+FF8xUPyOEuEnezrUvR
Zhdegs+2CPC9np+513WKG6fo/VPr9s4tE7Dw6CnQNgw2Z8DGlUDYYkaHkyX4NrYWlVcC//fes2V+
+pYovJNC8HRMfsxXquq6r6g8kFhp1a66ryWEiuVBzcheV63MlEDbeP66y2J6cMuhQNHR0OAuROZi
1vRFMD82f9phcSd0t2aTfPUbYiLdN+Ln79ZvkJHvClVs86ibXi3OkWJ07wuZti0nYOSx5WaGODLb
nnI9t6i2I/Qn6rkzJJGgQ7/BAyXgFVDig3GRqZCKXwC2unaPehsMEwIYVfwaM5eLXHn0jIavoARz
Ng0gJpHfSQP+WPZdba0ysGkPICNPuN+RX8wI8xsvn566nTAiOeF9vjMN5WYNUdA2FR8YKlsT4BE3
vMVBr/cz6Vv6Pm5QOyHBPWZp+kQbw5PErJ/W61GIQvTR7w1v+eQNwJ3+ua5pSeE6VKY1MxbT8k+7
ZcK/r1o7u30Axv5lizenAEywKxmaCRhgrVBR0kV30iMC1B+OVVNeFZsMgwgVcMuwn0N5SwGuIYB8
3184brn19u+u5s9DFfbkS+YMkWc36hWZeJpRYWTLpPaD+NN93mXL0KxYdoF66VFIyEfe4JIpFcOq
QR3QB4jskIP7VK2H7HYTHTm4+n2uzaY+MD6bLrNNCWA7t2y4IHdiWhXOWzT6dqOfYZ9lnzePVW42
rgVgbK9vWeUQqD48n+kG6h31368ttbMuPs7X/xL4i78rqzNcMAYNqLNGfSH/s7/7dzPgpJrzyJPw
qfTWtnpWZ8EoVmjULC+IVyb6UPheDv4npch4Ej5J0OQCbcGVR/eFxux4aZGDCrlj+KILJT3Ciq6r
+TiEtXXxS1gvdfOIVvY/ZdzTnkilLIR3T71ntECXupYZUJswEiQVbKrevOVJbmF5UNayjvjJfkFN
8Y4toehiDJIKe8BFDhxUh5+rkwfbTHBXr6aJa7hOvZZaSj5LwLxs5djyjkgByXVXzt9YIowGgaPJ
ew2OProMEILz7Bo4Fm5p+AWy+Y7vxPNejts2iEyn/+es354QWqRjTmNklRv1Ng0prLx0vhAJasd+
HIc50IgLTQz3vd0VnfF5CLSzQq23LCHGJkpGyz6Btc9hI4q36+H0OpOnk53v6VZ6t0DfyHf1+KF7
R9f8MmOhmvHOAZwfGEQ/3fhJJ8HVuywwUCPJAiD4bUS8UiTgcCZPD3sRbchVP2QN3QSrjij3yn94
EfVIchskuowModKrTffGChyh9vEOBsFiFVk0DdiBB2t3XUsrO0N8WGA5sJ74BDuqzd8dnPbxWwoM
H14ziY0C/erO0wIh1mYXl83X4OTROIuN8ZS/Zonpd7MOot40phQ8WlMQCSPHCeuyLR31DhQeDKGP
7JR55Eav0s/ldOgiVUvZaOSAWuyxTlsJeKu5TOtY901Z2QobAU8LQO0TRSPPbXI42vjvZR8SRDvT
sM+kIO5+R7KiDbzycmfwm5Yxh36YUaMK6Yzd7qlzXHFyZXFUebn9tGQqXR5cbSVDi0gSWwtKfBEV
EAN0nBdHMjl2cGleFiMY/JOXACPZoKur30uO4tEPNRrLxr6XzlII9ZhKVMgVcC3l0IB365ntOqgD
ZSRORbgXry2Hm70gxUPrS60iSkxomwh5c0uvojsN9pQdcunathvnmVUS0jVnfNFhlbQG4pg/cADQ
k4WTd4BRTYaxhufzAMLZ5pBf9kUdKfnD6VF5KUwPyTZxdU36dp8DTUUOwm3RjqKTWX1hg6mq6aCg
fbS/GkY8NB3HFfFVMkOiXLOzVYqhcbVEMROchCKdp7j1wdFahzZoDYWNNN9fmHlFOb5RgNTG0ha0
OzF6K0XOKGWA1ROxxSkDCD9ZyKclVo4ME6ALkyrAISz7Yl08w8osAmfRb1JgXFh40YpBk54qQwcc
Ouv87hUh2eCHUODuzovZTfjtXcxC7UNLfgPRTGoxWufkXKx8DB7NhxET7pni5jCX8rfFf7EJB6eU
yN+hx+lvNHM1+nea8os7IpG6Pi6hIrk/KDbcq3BIdX7MDgoNURjoSTQ4NxntycCl4UwHtTJqYkLe
eR4NG4ytp7TmZvWpIL13DmL6h4Q21uPthr+cGphZ6lnFLLQyBeDNkPEd1bfyqC+V47V+pyM6iLBD
L+t6SG27ahSBTqYOMdrpB7tVnlkQyEMP6Q1FiFluAaaY6qs6ypzOTPLKoq7VJKyQqt2XqcAYytLE
DAkeEy+P4LCsZRiS5gXuyCBzUQALibakjaFJ2cRIZ81fupDQPIjgdSwEOflBZCMiYsa8FRdzlmaK
LPZkTcsptJw5vBJoVXp/1n3jSWBcMJPWUV49WsEU7OP1plFqi5QHUsxG1zynfYg0ohR7bvs1lvzb
ooaPQTPd4iRvNL0lsMkslBix+2l1gcLZZdWY9yqlEP9UazRzQTLdTFOEKUAkRz9HRv6IbHpaP9GV
MG8U6kf6bv0L1M8CiwF6Mw5vSQK28DFzcf/FUqQGMfhy1OdxO+MZ6Vwi0Qd9Hrf6b+7be6HXOy+Z
m49rV7tXH+RBCIPSeSse07dTBRGE5n+PF7WKznogU3knCp3nED8iDwj/ITTu5wd8Ygx1gcQzwAX6
hT08WXcmhpg3H4O+WumHlUsvRxaLW+Sm8La8XcL07d5Fr21kcTtWb0b3HgZaXd0sV9nl8eVqi4xP
W9jsqrk7WjfBQEtnbl8mpGrUKoXZYhG4GTgJMWpr8cisypsGUtFyRQjuT/i2m+NSe4F3BPnW5mG5
rXBfOnY3YQZbp4qw6D4+pDbORizKVQf90EEIgUqGcYN+IN1KsahAQA7DQHWrHDYeitdxcEKFncx4
uECLoA56cvi+X+RWEenB92zLHBwj5Bc6xLevTW5ZYDsySSyQ4Kk6a3W2U7J7PEZA+47BaDyGOJNI
qTDMftMvewENek4C5pm+kH3G21wVjOkqnnJdP2Jp58lRn06FM2n64fFR1if/cX7wZTnw50ONPAtH
JuQ4jUn5adZxWOLfF8YKie3ZlTSv/eMhsVBpYUomBDc3zsl2kwDSLgUpDblXqPwGXokG8OO9uK8P
o9UQpm/MYzAe2IVGhEvEk3VddrRtprE5yRB4iqI+/buwwJbPIauObMJpS2an4jrVdcRY+41vWB6h
WgC1miVKYRYt2QIeW6s8sPq/rZ8P4z2Ni+F36L0REJOJ42PyrvEU09ThFGla6BVDQo7/Pw7rQdW0
UVi8j2ik1+ssbHlTupB22iAkq2gLayF7T8yQosN1RWmEG4wdRjEtNMRfbb0jQahK7UweVIabI6nL
TcDgp//phgds2kkgkWvIXmDLiapLQb3isQ2mNHj1VzYCBRFgweN1yfRJb665uA1fzpoNDxpKHS7J
3de+ixbhcdSI8tvXD8mn7bd4AQX1GhOBZOkBlHt1i7866IzE1N8xZ8t4vJJLklPN7fC8L554sQeu
VfAd7CEjlfqZk7js88DvCfuYDVlHXl8b8W7InkC4AroFoNiUhIAIVy6KLoLcBDNyVljeIRnP28qF
nsA+cqJXockilZ/UnwZMEf7wygSBJTNSj8/1n+kCj3M2GhY0GkhiY9DMrWvpPOnj8nP304kiY2e1
ybtVgiGjf1ym7OsVIIeOLS9K7HGMnG418OXKd0QkrrnQIOi3uEVfEMgLjek66DNWsFnSwMs+fK34
v4BB4O91ZWQqLWiM3/DDLZN5He1VvBS7nTMLKyybZ2G44ORiMKGgW9xtBWIKOgfsgaDWtwSZRZQF
TF9R3aBFrdazzVPhTa/fN1vFnHzpN8wkE/y+mjXl+447mn6PEAsSPkVj+TxJpCCVYeYww6f0Eamj
Pe36KxhAUZZoU1Ad7UXRvY8OQ2QwNJ4ll898jHLL/UPDAOQVxiTV00QiYobIvJH6XC3ZlAteqoCt
Ppz4BBBErORu32MuIm7gwTko8xfDOv0krZeqtV6sufkqRnJDDT0RGo06cib8x1gx9vORyeT1J+9V
AYFKhcsCQLzj0foqx5l1gutpHGtUl7cz3IfQ4gOaxdPxAHkab8WjpTFsqqjrpwnTMbQks30XszS2
aUEEykj2rfmfu+22gYCcZls35h6HLJ3/KqHGDjBIiapcg12DLdMzaQMIj9WS1RqYJilhCkqEyKuA
65DZNbKzTaIz95VjfF+5M8ULUC6FkgUBPCE4xovm2vzq1JfEOnEd2rcn+xra/T+7ET5/5rrCnRwM
nfHNoMW1vdCBCey+LkXfqkty2d3Wa6VHhu1rY4338uG4lJzfXKpvKWfHBklLjBaXKi7744a4wx4l
MFET7qDB7PGaEu/p6dOMUeVJCPDzk3wBkeHbp1U/na0/MoNUf3HsQytJ3aUrLcOW+Lnyt+Abnos2
bvccyyMo5BTnqgc2bL4ugn+LDkTBfDASteO+hmDTfpLHATN/Y7Yhc4iFoBm6QB3J3NFjAdtIwMNE
mBtsFtOeaAwbn4l6vMiloVe9yeHBUBfcZ9L9EZuCCcpcH0021TO+W2WLyy2YHs65uk21G/KVhxPi
JYtIasjEh6O5cMozX8rX7pj2yJBi/IMCCIFnnefwS6ob6WauOnIINJ85STeFlwECkY3j8RZcIVdO
2Etl5b+liKlaJTleM5DcEc05hG4HSMwRqD4FYN0IOV9yGYC1poP0kZYc75bhv4e2Ts5ydV1LdMW8
MLC5T9to4YtK9XRg6FTeDgcejnDHYvA12ASHr8OTy/C8nfozIEBwmYtc/APG+5qOhNY5vl/dOoeW
TcqQJm9IWI9RpiOoMSAUcl0ofxDHD8DZMBcjlrWxVGu4Hk9OcaUhyB/05rSDiId3Nk/foreDV22d
aOHAj2n6SxeJrL1iCzvyy9lVIXD7PAjvoivz8BubB946hsoaWTA09dqU+v4PhfsgHa0wO39Djeaj
9F4hjqE1aPUrG6OSxscJNhx0jKp44FP5dfKxHo2Cy2Y65YzIKHwoAdvCVfzea47QD0cSyRpFVNGc
KB62tfH0jnpWYICPx11npsxwa+VcoeoEoObpst7Mx9EbHBA4tXI10XaXowZVI1oRbRHO1gEj4ruj
rRf57MDLWUFXZ4XiBm3KWXMPH3AX9NulyXeglaPwgG+JqKUMjHUjHIcHxRiWAk7YzKB3qB+DYOKy
QtlfDVnbaMG+Aaoe3H9H85av7RZn3VeEFU60OJuLwYywdSEGLFhz4S3Bxsdd8hPNgGMdy5PAFJZK
SmAdFOEFlNWnjpwLiHkT4Y5XYmvI8ibmizg6HYiLZfnNgGBRjyV+/iCw5PY35VRz0dGszZkUD7+5
EuKpQDkW05WUfeVIjNylxrvNpjy4BfSZDv3YLk6OqT10LN6aITt4D/A7ZIRtxiiLSDmH+kFJYwu1
4nBwYBfpPT34MGx7gvz3sy0Lp0/DWIJSLQmIUozjy8AxQOOXdbyVNx8l4nDfwT7QsXwaCQLXf4dc
uPVQnXqDBuih528w+pLSoFkfZOZUwkxj/JnDVulQMjQfFYwAlnbH3eePyb1Ynna53673plwgREin
X5GwUY6Lcdx1zMFK0gD1bJKqFv4ONSlVxD79CYgsRi6RQCGlIjtTcD0NhHKhsjuz5xFJVLuu8b4T
zEpcybHlYypcgFATyZB54g9xewz0dC2p7zv8nauok67xp4Cvy31+LxBRl6UZ4DTJcC2+9DGhr/bq
ASpmQBO723w9eVjrwH2a/hJZd0/Vxbnteajvv+yN1ZspKHk3FqnC+u1fDLs2cI3nYiWBFOAIbXar
31n0Wo9ccQmwSS7cX78a6wSsl2dsWxWTSt0MdYMXe6s7ezsKvLEx79ecyIUC67UZg1IaKKMRC1Cx
axatplnt9FLcs7mVac604Y9kRD2Qez28f6RUDWtQYD8JIi1L90+j61pppDrin59XZbccyPqPWAmD
Wwuu8B6C5qHZfYZxR4BqwxZkpUqzuJ3BesRepjWPsP16hcubY8ga4YWnPmpj5wrjbKWx8s1jVKvM
IrhEbYx69ixNxO05P5wyrEdjViCPpvlaKc3zKAipC9wNY8txId78gAa5QrkizVgY8AztyJsiNWWd
xqeJ//B/eYy5CnOhkYwtOs2h02ZuSWI+b/O4UQUTmTvfXd2yytiO2FuRxhNz9g+zI1EaFqBbgjnj
mf6J3m67DJ73tzp/djWQ9u+WrKUlY6uk1SsySFpKWD5y1sq5eChjPySbUfon8/6HyeoXUgRDk8Ju
ukodvxzsrKBBxlYSYCLvhtWput2bo0xazpb5CC84MvYTI177mgG4B90Dly9s102tD3IrvKTjDVym
Sd6CEH52EeFffx0LlFs0Y8F3fePEw0D5nkY5sOc36s3jYaQH0wFPHM6815axm6AiR13Mq+hLdrFZ
OgWu35fXqLEJ/mdEV4qSG5ajIkOWc0AgPKMoauI8T1TNQb0VVNd07irlDEb+pEpCysH22072+ypu
jbVfXzwKCKEcNqLwbxU/2VAlHDX/Fzu12mUv09JOcIqAuUxfu9H2fgUb6RkOwwMcvy/keOZjwFLn
qcYMCT1+F7jHD9JZcgf5mmk1jNL+6XQAE4JlI2R7fadco7U+KhbcHFW/7AJjAzVo/nXlRPMC4Ywv
YzRgf5i3ITbaPnoPuBExx/JncQ3sRCZj2CScEE+LQ8HLUz9M9eEwGMQB2jtNU2+rUG/Kd8piOFav
1fw2+tpO0luUnGxTwS0nwTxc9dkZCgAcAh+JbabDoMShh6Ax8bnY0VofHXHwzgcdpqcr0PJiTA34
HetrJpMCcoOW2lsXuAt+TgqANQgsgnmcRjqPkqhxezXYRjLsYli+I1iinNOedDmUQsdcrgoMmgg2
+ZdNl6QpqHVDLjViQlYWmGXdfn1fPW0JZB6YlwITkTiTDTtwNbLJodQ3YfXGqlo/5UXKHXKCpzew
3EgWYDWDc1/uFP5VzL+zM/MQNaMPv4L1+rhZWFFwy71BUkFaBSCnbNyEVWrCJLubhMVzQgAg53G5
RA2FbaJery962zn5QUG7wAInWx857TfGPOCYOHaVjk8FVUAIpBrgaoSjlpJWIX4D+qiTFs7jlFLL
RebikaYYFwWHZv6XPnlIMnZfNHZanAt+7vjLfo3UR1b4YGk4x6DtB3kzCOkJXH3lNP6auhtbdIce
R/Ge9I2pUApo9/5rVTBTDdYwssPeZUEHsZiaKqpwS3hLxy5FNrrw78Nr0EOT5AhFTcRpqJPXuUTa
e3VU3FIa0Q5Deq4FfeP+x9xKLeYO4+Rpj04bl2wM+jnaxv5OTdYbJJErhMYbhes4lFDUTd+4WRWX
I3yZdVvzlLnCb+ktiNJeOVMx/lrmNTXrua6YbCUQx6phVzjNQbNRUJu6Ggngwe/TdfG+Lw9bSui5
qUzWP63YyJisCs5cp8SVTUvy8eUnrMR2ptmtM/qgGVNQ8b5sxAvfmjtI87LWwHJ36sAH4YfTq186
FDI2qdhWKs4EUsx9lm0K2FNxVMNsGCOUQovP2U5UVSNct4cMv4OmN2jm3MZ9ab7bqxmAHoxR9fTx
CV54uvW7fMzpTBGxqVx//z01pGqhCRumzhuFI23up7UeuQHp4NoR+eVGkTLM6yLguOJLl0aZ5GpU
vLPFUo0735gEzYLxjRNzS4Uy0IjDukNMfBXSXFigIr3nM8xF1eUti6ujoboKnC8lyiXLgmOwREog
SHUI8J8+jzxr2M9UHvXfh8Kyk6gy6utuG4YOo6YHNcBdbEvkuVse23dokliq9HX90CL4bRJXZGhw
SC7Ra2KxObGi8HmhlxDjUd83a/4FFeYQtYGuwRq2LfCaJihh7Qg8Z6XGVd74F8a67b8WvagiOYUU
ha+wemfcrjDiAY+R5vQinO8n7W8roTL7mQEfUL9GoIseu2cak55cIXHhb2i0S6boGXAf5i/JyT7v
E1bMV7tmKgxUl/5RQJsRh/k6R2BKfOeFzceQ6HTbvr5d0Zaxe9+YZymWuHNMKOP0bDj7EFU4gAGe
S/ozmsAECZALO/hWh3Sm0CY7LICV4N/0dSVMq3fb7NfjD9gA8AIWj+s3wDPNgkPEcCUZ51apUyGP
GLIYY0UXiNQ7GzQmbb33xS5hPuIUb/w1YDjTofgaKm/2XTFzdoD/w4I0ozaB3UEL8YS5jx9bNtIb
lNOQmaIsEJWUtz17f5pP2rSAFS3mgjvFRb6U7pTthEn8Sm3l8qFhSmzsZkjBhbAv5hbs1ugE1MJ1
3W+Tt4ixtE4P6AuLvMu7+b0KaU/W72OxSh54BuS+UCuUImKTOqXXEKyF6VU4HnU50bpuYJYRgaw0
DFyUJ5l1Pa6/R1gR2D0tmPFmICjpIoqYiwrFBm/IfGlazGEktXsfEUpdwPxFDdqSt6gLTuZLcC8f
CuJks4/HP3+D1TJ9pnJWjj0WAVwDaXbFFReT9Y0G7qXUUb74OUigcpA5ypqF29Mehtg3sqcKGA+9
2tCPv7DEQEl6IRG7Q/B3ehh3NokpzDB2rF7Xs5fCJUHUQQ9+4YPR/JbKE1c+h6EzSWRMCl+rv/Z5
HGgXBUr3vj7YE8rsOw1nCpnxp4geXFR7tGWFIXiqVvJdefMYIvSF036bYRzInpSNBwcpSKFqcq8X
bOyeL6iGB7cIyWLLNJ4bWOnb9inAiRdE1HL+vwvoUB801IJVxEQVmzTYnRVdZGRsMyBkvLr7ZYlI
KQ7HIOXzdizup1vweaORbQ+j5tl8+6312jNCGtRFv5Vz8/fRoQKrognbzqlolz1AxRSuwV/C9ezD
iajHITOwfDxdXHdwe6QM1VU6tO5b2yvuNrsGHrf5mL7n/QjAFrQDs1U40CMJGODPA034NUp59o9A
P5I+WTI/Y7p9EyiC/3HYq22+bWN/IGhZa9jGiJkAlJ/0RSXbv8i7llCQaOvYfCajtsx76DIKm16a
mnDGRMl6qe7yEH8lu1SrktPoLuuxikBm1Hf+OxSG2pHCja1G1jIwVRcT2RkwGPeFec4M2R54Ixak
VVol3Q0czx5/SBrueSkuVp3rurFyrKlNa0V1pM5nFz8OgqYOH71wF6iGy8CyVCWk3STNboJmweY1
J1lRgISeX483JqX0cbLSRK96JudK+xfnCO6Z4o2CwO9qKfmKQBa5VvWHkZiWz1EOy3R3J7f0JeLl
XHHWTy+EiEUJA8hSy0PHIlHcMw8NA6kY5OnPfGc/VWF1bB946HPqgIVvefuIFrQ92L8NhlOiTg1S
+BsFRW8pL1XPKq/Fm4hCKRjX3fsuBNUxwc+tQVgzZOvMp76WbA1rUqOtxQ4F4yN6jSuZyPJykTPY
cMbusBpeZGPDbkjDfkI8lJfoyiiN/DGikrm8V06jw5UgtE9mKSsdfTy8OeYtoPCY5MUkb1KBQQnC
YmHw921G+Gk58gDntX6+0LCkfaYHqJJ7SVCGFFKl6NZu3LlKvXOGFMXoOe0a9bkvAPTjflfCY6IX
U82lp8erBwQSZsiYY/roBm2bO08I9JBMQjlHjvPml9F/3jD8EQPTS3ym+FTE+kKgoZOecs/7I5d5
sHxozj34SdXemAdNoTzzT7mkO88BTL82BvV64u9u4SNTQ2YAP4CLVhFYZBg5jgO5RLfh0mrE1KrB
+nr6Pko7xPcmVctc2j53XeQ7KdTpwi/cuc5dEM/fNYLGyRmwG9XnYWOvtPylfNjnda31gsm8kkK5
ldxHszvjCKcrmcX29rbuOlXaMoLGt8xURy50qNs21A5a4BQXWx5Rl3ipwRjR3vWm5+g2GeP0Y5SC
uGNDbehMP74wgukxDLCKtnG5x3ih7jhGHDANP1xN9oqV1+QCJB+YEplYGSdohp0BJHPxE7UnM/WS
x+2vquhIa85AVa94ZlTqtaXEiWE7MXBdvicPcE0R9DmZSaXmedNZizzEdPT8v7Qo7G0I7zR98IN7
JnsweGNYc9pxNxYKavLliBkV6JoflGtBUQduKvjxePY0EaI93FIrP+pPBBnZhJS35MTxsUdKUhwB
lWL5lninD1PI/Q0/6tWMb9OuKaVV5J2xtt0BRA/y3kkqhGJYA/72h+6E14XG3afjZgwxfc3zQlmA
ZqYz51vwRZi/mUWUK24MWrJoogqvZoKsNOdkJf2KxlHG3yq9LGk+xMm0DWazotLamGIkgFnGf+uH
CoDf1lh3mE9c7dDZMBVD5/2eHycfGeZM2+7L5EoEeI4o6zAkjD3JFIPg5VH4OopGOksBpDvZt9o6
6hamQo/etQdSXbUTQOfn24oDG10dYAwiK2dQEEZue1x8lMEGaQKF2q91SxBkLb4oehPwvmF02WR4
6Ldg5prqrEuvKh4BqpfelN25LZGwt40sfGMfQcJrVfo0tMYUOTd0HfzTqldSKse9dqm3QDeYo4wG
cIkGFkVlzw2IqPIpiQrjD908Y7x9atWKZmvNOKwBCPaVQD5PS6zji6ubttXdO/ZWEBv+gNOXpneT
jREYmgZ8kfLnrE5p6xrERJsNAvxVWeCKUlo7yw9KnhaCsAv1DPSaQ7bbdfAJyMVuq+BaDdRJskmQ
o8HXutPUmIm7v5YSRPBgGzuVlsWpj8Af7Ck00icT4DqH5BYsfyylTcWZt+dJxnMrBOIut0Yv79Er
sK0qPiC2x2KppQdb0QGCPJeoyNL+S50fZk7VihaRjTqVIwK16eF5UHcXLuc8ICBn2dVERLMPi88Q
f95svzZvvaFEAhRZpAYoCaGWF3VE1z6a0x5SL9OkCJWGXF5zIjsH68kXiflBGQzDmbeBEECBBLka
D3wS7pftQs1hMgA8r8s8CVmQRy9nIqOsFQc0DAFW9gB+TJm2vI9+qxMQaMkVzuVH6CGAywWNrezt
v+CuDQkfpOo0JaZSIHgkGaT0Ruum3bLZ/2iNV7Ok6nh5AvqQPGNBYbq++SrkU4ggh3B1VJcno3n2
ruGbG3oGv0eONtQGKkdgbZ4uB0ByjdpeIgJysClY2qA1ybElWPkr+gK22VU4VGxdA3nn448YoDzz
SjlD/SAA2hhuZzRbHJYe6BDuT6vl21ljOjRLsi3/Es8Wqc7vHtvBvwr6FOIDRiO7C0Ai2A/AZ1up
Xpo+9dNuw+8ra/6TNZK0LQBn8x1Q82NH9ROzqe0VtcvEzM6hp96wEuGPjbmaKfSUCXfEgt266JYJ
905Dwg+OTC5oRwH/O5C+i8OOvR+2SCzjsQsZy2E8GXKK0oihDtdWV6bPDkzQFRgOGJjVppOxXk+T
JKFoZMNsPVMp2yvUIeuWFXh3CkG0AkXrDpVnf/CZULR1lpEbfkJvmuS3Xms/eEkJ7Gz8HEYXYZL+
UcWT/+Ug40tg2/GVT/1iloB/RrGHHuTTVlO3Hko/zFS0jGW+qMTD60bIY59MEtvX91xdI5Suv2qE
pFnx9Ac5OzUunjH7j0p3ZKp/GqtEuYSlNZA4uDoc9u5k7d/MsKpGSmBBGKp6j04xUtOmEWMTeA51
nsWnd2d5ZO5q2jzJpeSdC222nGvzeUFJ1Nj4O6t5WOvheM6kEKGm2jihtPgMbLTPfy3XMIuFmRsq
NWI5DDe3hJ9/AdtEuiI49f12hx4oDZTVwvRvsLQJ8DwZsgwHoXpf96QKyz8vWO9pkFKI3KQEhE8c
DzKCXI1vgxYPkN8MhtpJqX3O2cY7Gx4DKibHI1DiVx731lOdN1B6/lhj/F3KuUaZZwJOO2/Te9j1
cmE9cL3UTzgGYlGsf0KqcrA7kxlu/35/VICIQpHpb6OKpIqP23ur4eIWTZ1w47jBRoWkDLMO6FPg
mITlbgCsXJVHQEh/2G5lp69hnjtZurWiq3b70xg+/G5gTF/cB0zX0+cIS6D052x/2TiGVb2kw7Sb
HGntyKFOtVWr00YS8xq9dzLLrt34vMqJYq1He+uuq8026c+DNHhw62FqCuUoKFuO/CfTYmun/jGS
jDdcWdjHIQ2zLuKSa6FM1Me9ziJ3bUkr/Fe1wJUbGPjVXP41AP5I5DMBC4nl0BmFPmZ/lwwiwY2h
7Oj/+UQokQdXmMZcohCBbtS5e9lQhrkhAv21JQ/nonZ8WRAh2J6PPp90WfR1FaldPW0emK0SbxNF
b4Uih7LMHaK8xEhDCBZXsWwTYKhRnO35qM9gnxDo0Gkw4GQrLu2nOH4Gx0j6cSUjgDmseFCJUeja
0EnwuC34tVxHF3HE604Q53HTork5LmDibYteYtvb5gdYtgRhdIDSXx8EMuzw5uc2FUprvZFcR6or
1QY903gfa2H18PKmLZKjHCXGNJsErMach0Z+xK8PhE7tVWdrbtE6eOFzDttkG75O5AxpdplLPuXl
CWkgNlFJFgV2zb3Ro9NVO+81jIGr/TVa/tdfY5kdytLfv2rNpp54dCF4VCgnJ0zVIBb8YYxvc6Wx
JaHLiIcjBzCQvczR8t0vyu+oDEQ8TGK7lq5W4+WP0Bl310Mw20OzT5EmUnmMYlgHBzTnZHjCXYUQ
B0CZvALr4O6e9+J/r457Kj5UPxU++vxXjWQQgGyPkqOV/Icu/ghaGwUde8DHrgdBFVL/8CCPa9CE
nq6YVGbobRky3wH/Q/b6bfnsj8LKob7N/0zrnZidJmjjCJYvLciRqHgeRNp1V6Sz9pGB5mg1MnfX
vu7UL9W+PkKrVPTHYLNH0Ko8R7O4naKqWyeuPKJisPWEVmSCOJnPEyRPvpSxrgVu+UGohGFrcTdE
h5k9v3JlAuIorHhWP5ZLzJ8psM8wYpmPa4ToJq9sQK3lJBE/U6be27sp7vWRWyW5JdrZiboYpqoF
bGhOcO8syoOQPCrTdnE7BkFVGnGzUJwQzwUmdRzMN0UUAiVBQrEda4+80arPiUQhNPnihiDIsBDX
knflaDmKnSlNIr2ImP85RZe/NaQmTYrAmiELQ3UTkMxv0+2vhB70oZRF0AG7OPAvpQwd3Yvb9oAS
N75VgZfs+OefZPupkgIayvsglhkvNcGNMRxCC8kh5Kgc1PRzQBjyuvIzGrMQn/TcQWlWrIz60AcX
fYY5IS0Dyh+ZtPgKs6LMTL7EVrNBTN/7XHXX46MBwzODSXCKBf5CowKT31UrKZAsRZrki8YjfUe2
kLHBb7MR59HPFhhdbS95RuzIljAYCaShK6tOcJxFYl6V8CdfGcoql7E8PuHngkBDPAIsCpjWzUHK
xE3w8SHkD9Xf7rNK+rzRzrn7glnfxD9caYKXYp5B5WNg5tIyWcesQVe43lc8khLunZOIhaLfL+bC
ibrNyv5jXxSQwWTn4dvuPA4EL5jqujNCAX/U5SPOK9IQa0mh2CPiukjFnPuBNAEujAVNAA83BppE
m7MbvrbPT8bvqJWDiodw07Qaag3jYYPbr5Vi2H7cRvDZmZcYziIGlRN/Fkfvpbi30xg0bLmkV6Cs
XIr9gpqFIBqzZQALVn7Unh3qonctCd9xrU52PIWKtANQnxp/cvdNJNSanxRVdyDd8z3whkqrMBdW
mhoWzo9SVonK+hDIKH4f+/pLisN4GxIL1J6yV9pLRHiCsKgzHSKtcdodUl9tPLNspPDo6TvjlWmu
ey3FajXQGU4OBB/t1gZyQ9GqUSqOooY7UJ/JFjjuFBR/BCP0bLhIOqGbYtfi6oYp51uyk3vR5X99
zsH1R4J2OMpHqjn7SveE/9ZVnBilzUUgUx3EOOsGbFhfoYU+0QXkAGYx3omBFHCEgdhECpETPL4P
GSAVlLzoErbyrnYSo6G/+PSzB5Csm6TriY8dqyV0/svJgaH118sPMCXOwtjsQRR6dS6NFKaMCPeE
ld1zWaVIrX9WdUOLmgHZHRLgtK2w9RCe8ShP6rALxzHUK0lwYUw3jczZQti+DI7BH0lehtiXnBq8
uSwF95M8aGxPed6IDSM2k1rc3glDbUtPREp5mkUEKeEVF38MF5X4JhdwXNRihNw/uc2vMmLmVzHU
VZgA0bdnWASCQFWzpz6WV+0/T1S8Jwlm0hgCIOBtEGtVfoTmDy+mRxBXymsIpnPOeQcaTZsIadya
NRTZYgNA9w+w5TKjrzfvJ2+UBC41ywwSV+kap5ou8JqVxzCsBNhEd7PEDnG/Fm+CkZiCQjVZVqHv
yJgVJ+rxlkUngkrdY2x9PjQwRvoT4z/r4RuVqcxxNzNsLCQFgfRLDLRzysYigx4oxcTRRVL4KncS
yVelFclsedrzCALxy9XeQ2rZutfT36r6c1fW9WK2jUSHlNfTdVRMhnrZ6o+HTTr5g6pgg3JLUFtn
IC4ysTAUs0Ar5Ac9XWE0mwL6zj0BHMUygA2Png2qAOksqcSp7SdMZo+W8gvu/qJ37WNSmTikL90V
z8MPXngjfKy9WqEYY7kljt/GqUQ83/g9XS1g9Rgya5YX/TTTbmvjaKvjzVXBAVktyLBZV+468jTB
r/WBzgKZbv/vP3d5zwVEuX0cz4qDno6yQzn/p6sdquwdxxREkW4Fg4ubyedwdTGf7/J4p0Qzq4Hf
uU0232WszydpC6tF84BU0iyaDi3jlZdL10Hmcb51AgX+PPm2U1aG8/qN3synWvN9qVWoLyYTEgy9
K4Ien2iHXqeWPpJISgNqfIf1wFn9k8wWcz7OEQX1Dodu+sF4PMwIM1tZPD1pS+0V2Z1/lXeWCQcL
Q3j25TwNl65ZovctNHRR2OAiaKe3Y+JAb20hF1iByMaFvqYLXT5dbOXr/px1TRI+WxA7EkuL6CWO
6QNLO0WEimuG3nN8WOO7QbP0LS1d2IufW185I65juQE3aldJg5kzCJ5+RbzBa0IxQtqUbGbxkOmX
1lYEjFkNu2HIU7eUfo3Y7tf0lKklFnyG3KYL5mnNDgkBCopVlTi2LhxyzOtxNJkofHLfGvsd/dC1
JeX//AzsUtqw/IHf9g29lvXMYJnruhh8qbgvfc7qXBkFaOx91r0T8Sfn2VrrgE9kVmaN+vRqhT0i
m6SfhjOSXjQKpKCqSJlLYkeMUB55ZJK1fFwPDH0aon+VUT9W3oFdOy73tTA2NvFwAUcQW7m3OpYm
Bi5jXFKQOTPFrWOnwnecl4ICtOswet1NroS95+LFYVPPC/1EZvXTymrYeMAFlOJlg8/aZ4+3RH1b
8jyYcSf/YxXYvKQMd37nK6QqFGvY+w0td7HGwV3x/egMrJqstwDy/U2KdvmKnQ+AMY+NSg9hpKWR
j7DjRSoCeFwYe4z4o9PvIaWJJl6v2IsVj/VQWhIZwOa6Y7fLdcYouZCPilXSLxafGtVBf+9DnmGx
rs9Y1aSSPEcOANjMkybFREoc3c0Jp5Bcfg1LnDqQJKG5uCba1ZzlAsBSUEusBq+DGTCUrD5PK6hC
dCYRcaypHf73cEnJp8QbUYDG94FzMqnfznGvpDxz1IoGHvLz0rvqwBFQsIuBoLecaJjnmK9NJj4k
MdVmvhVfJa+qZdLh39yf8UVKKBaMcDHMI4UK1EbY0eeQwJgpq0k45kb/ui9lzwoekHVBppm5LMOE
Ibro+/nCMseNjkhHqIur1a1HArRrIe9OqTyp5Cim723ul/LAne0CeZBB/FCb65k0/Cwuvbbw3Go9
pU/ESewyzNSbGuf4x+WfRTYB+rVhiDJrRLMc2oRSvuxhU1lTOZhYbeQqBUBu9aAJZ0zisjcj2erM
PXFHy9/QZfqqAofZ76+JVz+rBuN33qncHvQ3zOJTMmGq7J5GhD23u4jrtcRHB89h0cLQ1zUUqkRf
FC6iTEFEVN0sXbFeEfN6CcEaRB+Fg9/01ygNWeoyhN85EGKBIUCfGe46VDOS7JK+Yf0hpdSFcjQ8
wd7Wb3fVD8yeAX1/kd2bgN5sd7leKeVaQFU9IfLvCy2S+3ml6tI/+zDT0yVDDvdYq940KeFsT2LC
Zg5hh7KnDA9a7pHxZ5TxyTMBvjK2eEKU4BegnOaxT1rqemHlaAweDhqnyyni73lSKfYzchFb/2/o
DCm0VT6vmR5/b/r8Og8vq3KZrRPOeZVWF1M29cPk9soInBRdnV2bDQw54NY9ngYlu6WUaOCPyh0M
VjEbhDE3tlgm63py0AAy7wkmGYtj+qubAJt+ZzGIMg/YWy3WWnzzgo9TV6Zj/9A4UKbc0YqQij+p
k+O0Tlx5UzXLkeCh9O0w0taME2DtLOngq/r7e7fIB/YAvciTbDUMmFuCNDWIiP4RArivArI3ddfc
0RiBL5spIF6jiiVhln5P1LzB0QV26sg9ofK2rbU+41n2l1hIgaD3bTwPVEx43HWP28pby6Fz585A
IMfIHDDueYS2oH2HQFCRIZ3i0h3+nrV0Mzx89XPSJCvSXcdIIlKLqp1J3XmNlZZKsrNnwqYmPTUA
uvEaBqh5HXM3CcDN0IeO9ELLsSL3pxbzjKvTkkxQ9sNpqD65ORWATeGR4cvTl4HhUP4nNKWIg9yU
CEVKbMlTujED6W/5S4/zM8ZfSmMVIXXn8UsFVKHaKJmlK5RzSVUBocWKw/+9oi53sj+43hEYKhi+
rCtDOVxouu9HQG1ZnQ54vW667a28yNMbe4mir7yr9dOZSSWYYw5CCsYKWENDbx8SFaf5N1DSl+SR
s+Fd8K7iCMM2ncGSq9XVA7XWgdt5RdE3ebyb2010qsUeQH4R/mEAZ/PkAOx7TP7eHiiZEVn1RVS0
TvTngiW14ubfWkwkrOGmSD9WBamZawd59ttjpAQ5+vIqegFLpKRdwtmsfOH7VvumgjodkcqgmtbD
7xoChvWP+ZkiCd6row5KB1fKDEzj19bncQ0xf/TPuYPwwVbWTa0PMm9IHuloHhqZvXsGP4rIFg17
Y7gmipBvlxirT4xFVQpKEbQ3uY1cROSyKdcRSft5y+OKbpcE/4FtO7b48ZuiRrNBcV6by86bHrrX
Ui+3U3jp5BBEMXRQwy440jRIz7Hf1+SkgsqhwUyOZ9VHA7oxCz9XyjCbpqJvNZy1YHhezmo10/4J
RULnJqqZKYc7L/3QyvaboVwSBQQz0KT4QtmQPL00n7hbib0LpTlJulpoQcBzYQare8s914bSHvmR
TZcdPvfHZntYjyKIfssYBm7nYDCx7JtPzCvpqayLGnQViayesz/Gz2HW+g86MK+e7SvhiVjdMITV
F7TqwRyycLwaGaNmSZcBR9qj2hmfBl9b7H0atTuGvl77xekZU/PDMSUgXg196TD+sQJbabBZ+PYu
sAkD1HJzkR762WTxXf+gOnmAxEowhsSjcuHJXr0zGY5m6bgaAspBuLJt4P889q+voxHGKvKLIrOK
wO21RzW2frvbwDtYDz8CrsXOoDhNDCvZ4St986Ze2thHeaJfuR+/bSvP4hLIi1u7sJYGijPZAa/1
phK/OpAvEqAlUeHlKoMfivLtoziz9tJj14J83prXm7l6J1oBCy+GAWSLeOMeVTFj9ABKTNSucjg9
sXmkU+4JZPnq2pbBQRg7KHmO5h4R2GyuHpsaW4CpNpZNWa/YBqAnNoSqyFs0nqZvozPi89L5VJ4F
j29IxsORR9MV1I0FB6AcwLe6mQVYkL5V9lj+1GU2B/T1CR1ZHCciXLoIl/6Tdj/Zc7qO1fdxhQo3
rOoWkk9dSobQGUc2Lt5YHC728AKfUndn7mGxhpAV+8XQhgH3bv14EMkJuyNeCYZjqzDmRZ0B6QAg
I2b9yz8+Tocmkok0OTu/PptIZi/oEA1m+KwFlS3LBB+Cz5H0rDdIKetOri5gMgifxuNTPVr1Xl7W
yA7dgV1aHZPjOdfJwEYaG1run5euPtOtooxRpQaeeLuxfoxdhBVD2xX7e8k7+wfBqn17WwQMYw/W
/mLmJyalYzcpXhKe2hytI5fl+nPXr2vqIJz1QaSXrjve+reEF0acQri9t7TRgnFI5ZOk/kLqR3nE
arwO/Wzcrmj25sD/FHTaRgPhfk1Zg2WnuF44VFfkTdvwG+yy7FKgtOPtJf9wnnB4sJjFg7CrMSm1
JXiQMW4X3QTVCt+4aySeFTkeR/VsL1btw2J5bW95BBHbRrWDdeLg3rXaCTvSWczfSD5k/AA8G2rq
wlwskQN9OJ1Wa5F0KS3IDmz88/3yMSXGcm5brPBwo6jtgswd5Hea34fvoFYOIcAiCGZFwenBb0HS
hHlCajaNjSxFX7MUr1DGlpjDxV+2JCHqfchzEZ1LbV2qBgcQexEZntroPfYZ9zfPicOQr5QSuaHE
vnYmbKIeD7UergCsw0bFKQCAbKq1h8RPsCSC0PLuHYDUX1TTlkNCAaM+K+M/oOqqRIh1AdyLMxh8
2b4/54oBsownLNGAEhQzOIU89rWoCIIFFNnsnp162Z1OM0Jf5qXORv417yLqlAExwQRueilMTrAT
flGsKzIAnYANgdITUv4BVh4ZCyTZ3J9BHEnXOLLYtUt6Q/+4aeMBlJci3708VL3aY0fdyDqL/oQc
OffPJak9pf9v+6bEIL1qHkzGNycJTlDSqEYBJNqNG7WA8ot+j9vG8gWKJ/nOnYQOxriaqW3kItOo
rpsFkQlKxOinHLjdCf4ZTLHwMzKakvQW6+QT+EAUQEBCZTb1IdDVxzL250LqkJ4bUNAJ0sRAqWtw
t5sPOnLeNfI/9xL6X1Io1yQbgQyA91fmtLJmWd4hobdtCZ6LHK6jB+WJvS53TlOzFq66HOLbiRqK
VqXEmNsQAyG5fuc1C8/tNunvhXt1ic1GpUrqs/w5FGdkNkUpvHwNocgJmMX8OHpjIBDFiVYiVEMi
4HDNGRykiQd6ShTTyV7XRvcD+6ZDhlA9Oj0RiR5ZwTEwKtsodJqugJFh+XZmZTS+Y8B3dmb6TESN
EFBK3qetqlzQkQ4I8I5m2ukySmzhWQn4aCUei12IhE1oJwmVDbyr7Ig7nl0IIAiV91p1r5Bi043N
LDibQZwx7BebZN5itQ8ISL4gvTSOcDi2VZDB4v06KhzfuBcEKLfgGBDTbHdMhTiy4cNAMBGedF76
vdv223haNOFJAt3ApInOWuOqEa9LS/1bozv9r6LEWmzxOcVoO4014V3vm1Ad6CbnqTNQtUXrd61n
Cdy0kCxWntDy/BP7qRTdboIrb+9DvcaWuf3CHOTHh/0VVVtQoCdRzREkax+xe7CUo763vsOyQ18D
pd4OUmeYckLOqlE3nWseCF7MQF05R0G3U9xfFQ28VKLOAwKNO19igbjP7CEh9IrSVQgmgcZ+B6rx
e9hCx9hGJnrKBP3or9ZGFDbN4vMLNvdahmlBu+NJUkl15C5VuSQ/ZxI2EGUtSDPaWTfCWch8zEny
W4vCy3qNqFD+wnz5e6EhZmdlgGTVG6wSCiS3IrhOezI5xkPXoyxKw+o06JG1Ho7Q142UjlX8wqlY
hOtmRgc0iBRMB4m21G7xc2w3zuEfnZMlKRDMlZ2216F6ZHeAjQduvHn/R9zVhQEETF7yAsfpiGDU
cRHN8msLvuDeTcaDNLVDQoC/TIzpQ+VocVmqpOwIrLkUyeP6Q2l4a6dWtUC1abDIM/15Z2MZaRZd
o3+hiDGo8kVqw2d2FYWXhW7S7aTbxHDN7FVSsGSYpHTxGA3H08L+VtdU1mvomaVLIuPzB3UE9aCP
Ru8Ujc5e6Mh/xSo2JHvRypR/ck0B5BH/WMtF3gOR0RIctgIE3s79L9gnWcWb61dWXwsI18oHvo1M
cv3IWf/Xt6cXYSEU3iAdnztOUlYE0cQga11I1wuHsz1CHY+swUW7JmT4VoTVK6sQxt2sBswi1fhT
GVc9rNVs8SNZdNlWd56RDquxDC5wAlqC9Hfz/6JR+8T1svfncr1cxeG8HGZD0TVZYedMwT3mPet6
sTOSz1v9/rEhKhiDAFWiB2JOW0ONEsSOXR6yriQnVwly0taSjp5865P4uUasmpPz4AxXylUJcLiF
gM0y1PFW8XimNkuAvyekK1Y5D0KMYgweHJBwXZSV2bDs1i79THxvo2u9OAHAxW3ZKseGY7YqOdye
9m25sJ1mVMIt9xHwECAotOmamsSJfZqWWzq8Ke9aanCGAFTrS2lLqlbzXojrmWcF0l0phkUj7c8g
XuxRhtyHGprHpeYVag+b/Cbw/ndMDTFRA2V5EaMUuqDYml1wfbvdpxWL9QQhOQIS4K+xEKKHxxoB
YdUJ0fgb0oab6AKZ6x0w4BCUR0EJzUxgauhsEixAfMnxNxv+vzdxJ2+nW0Xd+W6z6jSxG5hvanC6
o7a+zRqgYmJsPDDehkBGBfclpv9/BpsxTN1SFHwmO39vj0WcKrS/MAJt5YaJEEUOaMzMJbeCZ+ex
/Kagz0Tp5LKem9QYnoO3uKPKy5vJgTMaXamWQINRrMbeLibb33JNWPslpo8T8XBv49jkwK7C/W3N
ZuMfs0AI9EhGHt1WH2HA5MgLYsaJJJWYnOtkMvStVFkiGPJKF9mx8LPHJldb47BO/LEtplvUrpom
z9x6aTdvpxMdkEOuutzgwM+u4I6tJaWCAXLgSRyFDAdd+pSO5roWKKjinRmJ0z21K5K6lsrLGQrg
3xY6tUslf5V053iktAqNBchr4pLM2zoDphiJ57CvWTmC0B1hkuxcVkF4C+YEJLo/t8CUlnOGlIek
/HcH3N2aDWs+TJYYJsTvLc7fDch8NEyr2E6LPVrucwiJaRXrx4FB8gZ1ThxofbbjWCWkEbsZ3DtY
c8gTMv6uxFvhCDOgS7WAjT4fkwfTrBsWBfTUkCmHRrGs8pLirQ6QQ5bQFqx2Khh2sWOkBZN5CYGV
5uSdzkClMORZY8ZwrfcV+vKdWsj0XrJZ14Zo0sM237hrS04/Bte2cuNiQGrRd1kT2GVNlJpFJmwK
noCo1NmzsvSZTFnuDZiXmx1rAP1MXGDCJh1t9j0ou3Xu93dtXz3dDKDlgTYgjNyKZPWAmlGP8qkZ
S5nnRTIVxU/1OlEM7phDNpdgJW/Fz/KFgtY5kYhd4NzlGCY7IMjsXV1NgOkDUaTykoaY4WfVuFPY
WvwqoRdT6IwRTmWm/EyAHJtJrvz6GHziHiyXatrfrf/8BlQVIQgauYE/4VGaXS6lQlCu+WVJ/Wt9
BOnkMWrk+Z0W+IvF3H3J/oCK31VoFyhKjPHo01LSUW36rdc/wGpL/YFyLNel6C12DrZZeyvEy2gV
k8ueQ4hT91LEXDcCivJiGkd8/lD1Ynb1z4ere07Rfqb9gtLdSsLQlm9hisOo8oU/8gAuqzbC9FJp
oXl5mZwrQWrb151RwCnpeOJLnP5jmtklFa9yJyp1pamL4RQS/rVm5uSHSG/gUrx0zRki5OqwjKDp
YbGWkd5xLprryI109a7fPU5Goi/3VfaO9DP1F7aV3SJgIcQXPfT20RLlokuoMK2WFFmQLKdNy4ZB
T7wTMT84tgyZlzQIfJKk8+Gxvs+G9c5w657PSfM+4luvj0ZH4S1d+z7Jn2D/0NZtsvqy2cLL/PLH
4TS0jkyTH615vcR2JLScGx7Gj7GEP5hm7afyMdtbFv8VuQEcWlXkQEqvy3wMaPkzXPnqX1gbhFPt
dDOo4LZx8IQt6UMU8o8KoT3qDBiwFc2TsZiRooW2LqG6HUH41kugO1uGjMAzSST4wqK3sUxkzSjU
QujUtEN74QpjYaU2MIe8euhVFLsUq8zrZjE12v4veULJoDp+PIZgWTJf6eL7JOeTwKaSw2YWnfgL
59x7GCW1TCVfa3NoCQYyfma6gP0zzSPeww5D7lxDFgYgvY0uSvh5pH4nQGtm5PzULW7Ernzj3Led
g3AyJxaitRa0K4VmhZEnzuPq4kyRpX/QbOiSee1csU+SSuoOWTdHvN1JUkutlj1wVrHuljERK3vB
HtM7wFrhhgu7hfsyUZ3GwTO+fQnxbIz+2I0ye78ZCtIvB8349sFFcdrtrfX7kOFVgxU046m0U8k5
d8bjrQN2LIncinUEmxjD6pqkRdS3MEPyMVfe2tnW0BWor1RWyx04Ak2rnzxsOaFa1oZ5GsgbJ6FK
PxybdtPtAX2amz7Ovwvver7Z4zpTEFUuQ3sXKXtt1mnbGrdcT0iGz2mjz8SMwbdnQ3rfIDOes6R1
55JAOkF5Mh4HbXatNzhA0dgCbhXGSZfRFMvBTYwPaBtP4h13A2K8NWM6dR7TDWirfCOVMUShA68k
X18SiV3Vk7AA6pcJWCmLKcmhSF2QN25UBplCCw9uj/OWd8Dql73V1Qx9aS+uMGXtFVIV8fFrsi+X
aXY3y2wT0tDnuqPCPmRELBPWIURQeqdBb78bfE5LVvknAU6jU811vdyIsbwguO4ezidbyu0M4l8q
f2Z6H975QP+W87hLqDOr728RR0XCctkcN8MjmIphrLtSuYlBK+jWEPrMQ8vuH+wx2howJzR87WIL
KKMzA6JgY0WcQaq4q45nC+wFohEcVeCC1QZeUFOv+6IUL9HrvpOFQSonqBoOX8kcGgV+2WgKcTKA
4hKLcfF+9JgZUArV3QH6amu83mjbT+Ww5geHqaXnmGUKUuJtDy23jBW9pvFYASmzS26t7zqj0MQ9
I9wqWDy/OGgutYGWdZakJbeHko94iCyCkUL/1tlKk/SHww6McPSHFO66CwFaGsNmQ+TmRImPkF6B
k+BHKpYPrj5NOET2S1+xYmKNZWLz4dyRamSHN7044E7AuQKWGq4u3K2J6QglC830KSOPvjVoN/Fy
mVVbK6p2xzmT49o4dQsqo3V2N6QRZGaZSiCMSZWIOEsTusrBjPesKwWnJP5X4kOGEKLIB+s5p6D7
ez+HybMhROlt+grrpYSmWilkKIDCAzFI+AKaZXg9jGu7SWkXDoGugz1okkjRas1/ppM4feokqWG+
MhSIocxHndmCrheeFs5+kEA1nHWcOnLWNWgrW6Usbs4sQx5f1ud/sqUwO8pQw1eIGNeSdj447YLz
Zsumg3BLHNtjDD9Ydgpe/SU6rVi59XWGYSBs/jWJM95JYzgh62/jrJK5TeRkRnTnnKmvONnyypvD
F+WWVHRb+TC06M/daVHTcYSpE0g9nrCMOIEUWF+m+NvRa9K3IY/JsigNY/yNox7c9e1yoaxsxxWg
wJCQ48X5s31W88foHosaJ4eqM8tG3v61sCzYbRpxSvp6lVp5hKtZKuN/s6xbDsQksmlwXd089+fZ
yhyfPfCUCBSwNGE2FMF9u2Q+Ddtae+OgVKl67z37HDwtsy9UkDdnNpeQML3QjSBYa18mXTD0rKQ8
MgKcu6W5/qN1y0VoBKKkeMIQMsEIUy6Op6pbkI8cG4NtQT9o4uZ9CnPaKqHoDDMTGv50ZPmvmGRt
2DxPOt+MvaqSkq8a/kE40vT0akSuc9vBHPAa//sdvNz5CuUqhE7klksHWc5Sbui90D6FVg3WPKNf
pgz7dJKrrkVg8rjGsDNU2GeurZGiKU3Kv2IIPd9qMfd4/rzqGOi4aQ+pzY/EEirfrVpt7EZiumgt
kFhwfv8Wkx/fSHKXPJl+B6nFH8xApo3Ikp8aFCIDkI53wc80e4eXMK0PwdAL2zOiWZ12inLgASpo
LlvZLgKKrV8A3I7IB8+iln5Yrpy7CDjzv1tQ2TBahiv9AGTz8Zzwx1lxGacq5LBhUyqHF3cVxBGD
KwRkiw+KkwhVRvqwWnc6XW0oFEbrnLjFDcLzgvpllhpNL2DdR4ohCeiODF0bOhIRVOisNvYoyHeS
qFBMkxtQ5vXT52MqpX6g/dvQQjALErLD1Bimcuq9fgvJfVhZ5IYdrcwDpmjDVI82L6pZQkHEhHMr
N/ksN0Ysu+UvF+QVTv79PuuXfS6F+pjN6irwT32hnRP0OnvgsEu7o+ypEboPn1hgJMoolUT0cfE/
3e5r8GbKNYwPtj0mnf6WNVtk4SveYcNbMs0a+OwjhxYZyFMw2NQWn+E+JGT4Jww6hd4+YMEpYsVM
qnytzZmirt+XHCbNydmSGxxdTkzSWB2NP3Wz0pNbRAN+kCuBxX6cMi40CNxEjejzBZYwVJOmbJ1X
NaOdg5MgrbgDQ4THHSUxpZAozfQ5Winu4wjVMb9vq6GRmNNbqjsM3WHZfsMz3V0j08v0M9T9Vcd6
8/wccEptF2nlGk/YcaiBOF+t9KtMn+h61XVCY0mgEer4V7/e8rObAfkJScdpLGgxukdo4EZy498g
eC4oHiWoJEefmBU7pt5A0uAgl3808eR2u+8Qisf4Af0rh4RmtFZrwfga17VbLOHA46PXgPZT1orT
IXplQKBR3zr2IVWNK4IbM5Wfg/NdiBwmB06euSqkryq55G+ZskG/UQAW8g9YvXtifoo5O2OS34Iu
IPmYvqVkKAgEbRbIPsli6ULGbiBNNIhwpxYuj3a1oADbaIIXNEU9mqBEN1bCR2pHEakiRubPRFVG
pVhJkDxNV/zaQ4qwzCTpghSWoNHcZsIFYZv38Z43dcAjsR3SxF30dI7MaPFHzQj0KkyWyxMdeJSk
KrTpMahehBeYYH9zRGyLPdTLH1EnPsAv25+BjIQ6RS1YTPXc7Hqcj5/TtDh0G6ShGmGkBKmdqI7g
9aRccRaR6HWqe3LEEGL56T2N/aygX/E5DqbeCGA7FZviqCRDwUy2o8+UmuzaY21+mJPEKZMxrxgU
j3DsxZ73h2Cew3f5UO72acP9KrSORSaLFzMkwRbl57Rain9llwOKxBA/Q0Er6HIOAXKwbBJDERBT
g2hfYYqW48THFLKOr13Yj13ONPMrHdmGYG6x4OfxkqoFbw9mIg3jXcn4o3xIM8XLAC69dOxv0Hhc
RR4pnIUm2HySpwQUmFsIEuFXyP/R0fUqXUReuFj2gvpXn46tYs0Y1r1IhsTRubE4h0k9IJC+KSgB
2w4bDyjEuGMU0Ub7sODNS/kvrysDzwajQkvjkwzdGMw7EF2YL9utc3N6noWhH3UjGjk5wyDM/wOL
NbRvKtb4WiY60vTMWlgoY434a0P+XYsnO6u6axTmXox5IONyu+SnsP5253VD8vvHdiUkHP7ZoBtl
IdH3Y684E/EuHdC04AYYZJ/ZP2iIyF4psUAVqh127bgqTBY9JU++J/mmaAADhMzvvuR6SsMYf0mr
Eo7Yd8R40RqtZq9AUktJnO1nb3rgm5gCgauiKRP2urLVo5WNIjgKvyyTTQlQT0p/gsZn2x/41z3R
2Uf8MpXxBNM3PmWSSDZGq1ZywXGxTF5fXWJt0mdPeVjDXhpRYR+BOFH1czWDZIlTH22sXrINNBH9
lhRAwLiL9W9R29MJHij5AgCPFYSnOEK+pzJsKl9hJNgTMVXkSU8G1qJgnH+fEAJ4JCEUJxeo5w0T
4+zyRIor2F4dSirKLxb3imbJSSy9KJjelZBGneAdz5cI9zkKaM/oIRJe8CqKcH3zhXqeFIbymU/a
9pqRwAhp0OP6ejUKkfVrBToAylE01ekUXzl8QP2JHUQinSQZ62TPNPhN8z4G7li4WWbQq4MV2haS
KNmAKCpXbkGMmVJHn9RjAj3t0JZO+4eQPPXOrE22bynFJ3xQNxb+BI8NYxJ53dRb+3ld53aYzytA
G1+Th7mQ9hamTibjot4CXvf+lcgBONgsK50r03+P3/jeN8pOvcwyOKFlbfF0Zp4rPe44EpmhIsdx
+Y3j0C+S/A7QYWROP5PGwq4bXEpIXKZcNDAaQcy4iKoWA9ht06SLuwceS/WcMFk/+94wGiW5nnO8
4bkK0ui+5xt7+xnldsgZpZVjvlGwDnuJ72IeIDS76YAA3DSZCVznxoNLbENbCqkUBzPEwPk55Qf2
B9i0weJ8IJ3uOn06AdVzq0WjnxaeVFW3BAeoQZMt9YaNlbmCVP+0eXRr0UHdAEzx4U1pl1V88VGp
n8wKxRuEhdA4ho7CxCvwQ6Vz/3KrcUljvBdMC2hm9FZ4K3c2JQS13XOkNIpCbfz/NeRlY08gmcQZ
/vms7AaYUKvHJahRKE/14RY5EidiKaT+QUw9WBDNRITvbbwJK0nxAESquOopdwOvEyEclqx+623n
0KXRTLsDk0U5UE3h/XuowEA0BmxNjPDNrQL7YRASBDWon8XdhPuf2zYgXMXGRLRnTc9lTyaC2FJ1
NlaLbgmpcZ3vjMb3dnypIfRDpOB+aXMwRrLLv6ejgHHX0H8wZ5ipG2kdaCOZA+H9fsyHswc5xMGK
SlPQOFyDGZM4pHb6sQ8DB6Qk2xACAzjngZQb8tEkTONgnv/fv/PxikkvyYvJwRcxlFJGAcFxYMcC
blam6Z6PSso6G8dlOP1s9yh1sV/xT/YmEXSfgAwt1RUXs2VKqLICAycP04h4CgtrB2RTPwJ7sfUl
YObSD53dO+VIQtxEHAgSyNKkGbyKI9ic4m7L/8wfMLxBLWL/Qu2uEZxNV3OisapyN/6oPrc8HR2O
wVMDQRXmvrvk0CfC44No9lokBIsUybmWGmYLV6qZ8dFkiUT6JOQ3YwJvV9dQVaj7tvnuLgT+yxFC
+m2tHjVtwjPf6W+v5/GYnR0eLtgehHNto5E3ne8nDdTFRF2+O7gZs61wqm5Je8/EFcut0zwkk4ZP
10ryYDU7IQ3AyIdnFWWme569eF+3K4cKM/0jNqCZ0aEJ7/Gyf1Z16CKOt2nWX45yzZjVd+SYtOW9
ItkEBXRkzzu4EYUeOJyN3Tw7KHLIhR/7F3IeplBsPnibA6v7kIIrjk7nkIkTumHkMxrv5Hlh2xyM
XWJw7OK3QYoR641SuYLzlHRSwL+4in6suU8Ti7lb3vjUnSL1eBLTBhYvWOUlFwahG6xlWw5+l54B
dk1dWamPyOMCWG/YSAyQmUXz1qOhXodhcpNDtjQeXStdGzWosAKas0m1qv1j5gRdfx5E0OszGyV2
CVIjg/TxrS/c7408UR2VmHs/U02v9OssDXBEvS57B8Scf9f4W2crDHl9uAXLKm6nHgPqHdB5zPFe
IflPcfGLtJPNCVBaR8dpYgXzSf1ojpQXc0OwWyzxu1GBRSdcxzSQCbQuy1ZHBQaJ8iquHshnZbDr
9TWgThoO47VSyTUar/gsZICCf2EAQlqwWIMT+if2Iv1qUZhGN3RI7Q8/MjgQXBBOW1y+0/zUgm3E
zFP9SiolHEpbrEcVSZvIrat+iN49neLVfizIkHAo1JY/VNuDCWtqkYJdRZALSueT8/zW6E9Z/QUy
oXtNuAG2RTIobMuJSG6EBh07w7Y51FN6ZuDxDKE5Y2oMxDINAztTZ4FF5AReLaEk1txM8QvEOlyS
xyA6tsclaZnEgP9j4LIJMuMNI5GPpIYGEvC1a/G8B6WrvZTG/L8IFLjycSOlZu2m1Q1dTBx+9BuO
OTRRDkkRxtt0GXFm6T6qxE04R8Wv1IIaYqTyQdn4bpWqaMWjnZIwzqWBRYJEvHlAv48v44Hnlpct
no/CEBsORBgWUk9HyZAe9VCr/Pdh1eM+99c+sCQlL2NGbZxjqHIkRTS1ScKA/8TLCZEPGj/0NjY3
1cyoLcOkRrYyuRRKGutrgs+k3JtgKJGF8K0UQyYIGDLQKuJJponiuaDLa97JkLR+PKGRXLgiSX7o
Id+sPNWh98jdO/t70tQcMLbheFKTDOkCxQKesavzOEHZki5FfD+/he3pI3UbV+6fe34ElYQCY6MP
3OUNNZ5hSqsXpbSf4VrlcRbbGKxHvUEZ8QsMCb5jtpu+tmABOhNvKswE8IaTMsG3LAkREk0H6GYv
xAqUhRwY0tdwDzALuGNrFV6WPLohuEvwbrq5Ig5mYUMi3OMtMz7v04Ca8laO3PlxUeXZeErw+3nJ
IfP4FZ4BSWElzWlnbii77FbVrRasQb3PM6MnuiLxwrla0JQmRbwmIm9TQ+IJszP09x8GFZr8Z1el
o72GOYuFDFx6Jo80XS6Cx1HlwmdBILiAtEC46HYtqLDA2rLcj4SZlmg2G0Bmdq0sSWH64kPx8aeK
lA5m7n3rakEZYTQrVITLqIgbMAZ1HXJ3Y2AIPGLbOHJgjsH446xszIkqtVEBjSoNCGeVHWwXH0V9
zvJZi+yqdO5YSp/ak2iGzXIthqAtU7JQeF4Yn2ciXJqhJKtdUsGgnuT6H0di+O000+97SJ6zm/pB
ysHnsVKlxyfyk0EQAA9ftG6mFCWslMSALPkV4Vr3Zjy67BUVd7rfDrYK4xO0g/G1SGPKEm5h+UQj
IplWYxmqWYGiPQPdqfNPgMWQ/PrXx5OkdQgIRHVeVFwKxVswLoSi6L1pNSXFttt5jZGYCEhsNNL7
lPo3e8O6PFcrzqHI6I0te9WOXNlN1PepvobV9+KQGZeW/4WnAQrQh9JXps7zn08C5MvliWa9O5fL
gvpG+ty3xHYriL4RcNjwTVE5kdFJ07+H0BqKCVtXDdxjyvjy51OWL4qpYLzWn1DUZbj2XbfEY9DP
dl3jeZiiIWNh+eBm+BHPFuRU3OuugYRhx/t2OhLI2qoQtB9sI/TMkm4aCv0MCr0WTi6za2wyQD+7
wmpN/yAw9fSHwcvPhwiFX+uwIG/BY69cJbcGDCvpJyay7TWI0mqfEzhYcqjHe0BfJTIa2SOVJ4W+
vQhKQCwL4neWKp/4U6EodjW83ugOHXGvl5fyfootFUUz0KjrgrrXq2KRhw6yfxFWd7ZKQBZ5gdi5
wq0FaOOSYTOeWWZM+Fplhcbl76ESOYITBWAcyQSGIkVacShURs86ew/vxj9jXxUqs9avODQ7SdaV
co/6L0TtsIKChQP1P9h4/jXW6O9SG0719n5M72vyjIna+OsP5s9kmlT4hSymsa8Bh4Twh9boL+zU
dx1PA8sj4RGCWax0yUap3Sboj7SctFkbS5DmfXmfl8+wnwybxsrx+b3MYGw1yYnThG/1Y1QVYmpd
bwaD0XmwMe9EdnUACVrcqkOt9i3P+OTDubfpue1tsPg/8Q6e08VQD+tFOOrIHphESl0pJQpLkdkZ
8ueyToQWio6s9fiShmFvE2mxMKoBdzZ8aRdWtNsyzgc20Hl7YxLDQc1I7zi0nE2md7lOaFeNxOBY
nd6SLO7cdDoRqiRH+FZ2Q+NKKkpg7IgivGPYd0wrD4MfSogXvlhp/NYJ8bX5V+sF9YtTDdKaZXpr
YHadwqqdOSzsLd3AHbLvlsB2uXKfm1eCipNMTNiI8yfI+NdldHA+hDV63dmHUgqwGtmkkMydJpp9
kqi8mrIZQ+bbg1nt4lymVXhqD4VgpDS4oX3Z5B9sIi5ZEUIfsm5dKI9Zteeypp5WWjUgjSRaYPcg
VSF33hoC+mM5J3/5tG1xZX32t6drjujL05qpgnpdsyuqhKB1qOTbrTA6VN6ZBVTSBrKZqpJ9APdT
/6bdb/v8gN/kIM5qicnuv3jSWG8809UU64h21qK913xf+uWAoDWMZi4aRh0X1JIufuu5o1qSQ5Ta
1TowrPwJJhBAhRif3DNtc5HEntOIo5sPSWW3874KVoHw9Rzf2eaJFYW/y1UgNNGv4f1/sVw5sEuu
MZeQf7ZDo0pbIy7r41Gg84dav8w1tQpbWp2BfRLtMx4r6VWKNjOUrPPZu43t4M59dssntQr3gH03
jw/Pm1ugP5ue3IhW+0bMboamNpthMTRtd50ypimQMFmbMLBI9+6nBCSTRdQDFsaPZ0rvfNWKcHYR
Byhs2JZIYjQjU61/nB2NKqEE5toulyVa3IkDjwg09vUA2yhv4UX6rlmKONfvQ5XuJcAU6R6xIYjS
mXt3m29Gje+ENQFBqhTAxw0GozI89jYLA+iTNgVBDRsJ5bvy+HmlAzVPPOTwWFj5T7MAUdaKjIBH
A6SznfgFKDDtRLmGwXz4fQvnsB9EAeIjhwJCJfMgvl0bFFIbtodma5P6C/zNFpwr8O3c36YRpm2t
q9rbPL3HkHoNR9vpAneimDOrzLL7E7eXTHfVldHGWM8DESo2nXI8uG/7IG2Ll5rpFCG8egSp7ajO
rb13jJE38uteW4eN+L+1wktZEmtKGSVGaH78MTmBmS6xUe/NskSy2WZjVf8BNDc7pRyGFR46/1w4
lEca8ZFefhmJXJzNYP/ZAsqfOcYhU8DTXp0LlgvQRRVUCEbJxH+Nm2H/0MYceYgy5Eyi0758ObnW
fVemV8pTNMIfLwSpunhtajjodTguyoFcoE2AaabPW6s0XRteITzlR0UK1Va3fLl9SLA31q7rkTZU
zREwCle5ejW5yjzb7arNDAT+nxfa9OKJhg7fcAHiywgR8TE838bqF9KzNKwk+4CdOf9NFOcwc5Sw
KJemxDP03n31YmTaeWDmsE7WT2TuhRQsPpOc2UJzVnA/9rpaxkWKGwZR5EAjDyEiGv2qPeYqP+KP
Jw+0IcWmNVnicMzZVmJEsNBhSNWEpCeKZPO141EBHSQ86sr3qQ2c7UCxfsCDhAhOBkyqEqC2C8mi
wWNybjO5xRhZ9OyFW1I1Wgj/svH2grB7t/lXDONl8bmLqgxyWGawhCihvp/9zb86mSc6XIJ/c8PC
diYmUxu94Zz463Jb4jY1iBeqeCkM33Al8UerLXsZIIPtFoG4TGUpTCrAUHuZMBiV2p08X+rI/d5g
R/qIa6ZHwmEyhShpmG3KvTmPcF2Gle32PC9Hygvm9QfjxzpUhIbaTVaIU+2Fsef4j1nnhs4xZV6S
A+/T9LRdUHPHxMLbBlmwriLLmmmfaMcU9IUzwoo4g3Th+w8GFsrTo9cgKXZk9ysSUqrHYv02XcxS
QUOwyGaxQ1zlcmiu8JY3dDkyyBjnQ61y0DgDLuZD+PHgbNh+p172H8QTBRPVh3qJXGOtV6BDy/2D
X/rjKEH4DHqOuEvo8vo30zOcjaBXtyzVgtdS96cTUNwi5BKNRPu9npQk0WQfyKIwlN12bX+E6QKN
cHpZUNGiHN3uyt//J7Nuf6laTnTDx2V05NIg70K8Y6mJAFWWwVC++JH9dW3F42NtIA6QpVHgdzzv
B1O4QYfUWAQHEJEAPaNouvk5BhIHZxHfz2m4CgR2K+/tuChYPAtvxM/nyg3NMuk81RaMBNh+W8Vk
5b/xek3DPJcKj3oUb5eYjnWjAcPo6e4wtrwBeKHQvFFgYEKOie27EbmXgWID+fEmy0AeYwjoQWF1
3fQ2zuBgSOcZBo1d4TXEBz0adhmZsR8ntMekcALEbDcYQvlBVl0E9/2eupUxZN6+ybDtkdB8D6hB
D06mfV/LZC3sNuTsd26ncq/IwRmyWFurq3tqi0a+O9QkhuItE81BJQyrCHZXTkEEa5IM6hgQFc7d
S9poEHyImZ9hdOizVj0QZIC7Gb55ciutjRC/e5WK5UwveJsSbUmzcUqa7QezwHXIDUlwyAW0fnGX
2m7Bzoqxcf05AYhhBykaJBLhORc9jfZK3PyJwh73UPRqF10d+XLoFcyr0+VxzIiOpiw4yJPeh2i3
PSOMXoDHz5Tn81a3ncHYxhHOzAavBEvSA0+lpMirhpd7gFt27VD9CHikzA+1ZFuFoj7F6FAoDhca
AKvmHgQnzya8OHXuvwKgxou7uHWTvzLeiLQBAsB9kqL5bwOGrSTC2R/EDJjKgUJHThRzjQQu7reQ
RP+l7eMl7ugn/A4QR4RIdEcBHthTs4Rv94ew2n2T6KAXG+1BpB1S+7a6WlCbzS3rbduydL+tyGJg
K6TI8tqYFd7ciA05+qL2U9MleJqPFx5e28IZ+ZQ78gwSZW2Oq25Z4Cf/p2L9cGFQ62+B5YtPzFJs
AEkVILed1M6OQX/WVTjEANyAVj/jQwMNbpC10ArG5ACotjuGTMqQmGah71W4Ku1aki7FXWLetsnI
D1zkRMNonag00x5SeF1zlWZqb4fF7Uc4wvO14Bu+cObUrAcL35SmhbV0ZY+I8L/r7SxMxGYqYAlC
z3nosw0Hgu/8GpBBVcJ/uCalE+Wu6S0VcpoSFZ87zWCETvmvgaCYcZ0/ie7tJxhEwwzDUDhcUiwq
6WfxQlvEX6eoNLNCLp7+OTzsUuKuVgXhq7iTLeUnza20J+xExQBEo4apJa3aGBYk7rygFUJyvbGH
+5192iUhkV7RhtsLKYtpk4OgBBB+RZs3rObW05Ne1Pj6O/pVPML3IY/ZNEhY9xytT/uPeGb2rckg
cZ5JJSoqZ85qezTzKft5YD6OrGosMMzI9P4ih+Lqz2lk+7fjCpENEWmZ7fdSHJ5Zr/dfyg39DVVI
dlK+uzTVWIzWmNrvhTyCH9axVzC/vSS0XKdA/YT7xfJoE/sBVdoQuu57oRWxgUvxM/0Hh2sYsiul
pbLMcP9q6P5asIaHjJhibwXgH6Mov+IHOrtjQ7Vee6RX4e3StcSj2xtR9DS+fNdY5he6U/3e865e
gJqqulILMQwnQNl0XoOviS0p1v4d5sR0NG+RxNgAfm7Tt9XX90Sk6ClTvnppBRMWu9O0TYceJlje
yh5QXrbbhaEJuY8CDSJciljdE9kEuZZFDbIvG3neWl43omZwiL+ZTEpZ+O+N+ZUnLKGcxklQeFqh
3L7NxV4QMeuY7y6M1Nh8zeGI88aZp/n6Bn0E/kJDI7qUEikymyiVSTLGZaj+klkSk1nVO0j29Vfy
eMqYvy9NUr3ysuLIS6WWGRBYDtwCuQHqNJRIIgpcq67kFO1wT7xuxa9fHbjkYyOvIYcHiNQKCsPk
wpJx7wOGanZuq5ijJnIV5yky7qOxqP0FAAmNuOvpGuyOzbRPhvc+Maq1T+6MI9ANZ9SxT0rxM8na
oJ/r8kgPdlafMk/xHwGDfMrnc7OCIXtxtoRX/q5vxIKqDai07tPkO/wtZUL8nuFFFvLTUsrUATCv
KN8oEtaG230Y77wLs7sAiLYxSskM1mnObFYRmp/hDi/QxATRBku+CHeLfvyEy13RuxjKo8N/TFq+
2Wy25sW5w62qwgsb5dn1TC/Cs1nLzsPBe2pcNYkKm5NNy7Zo50hsEA94xvjKessEjM+NEEcyWhTQ
JU9YDhltqY3AHBACtAezYgb0YqMih8I+VZWYPhWiYtdMPes0rMQefUg03NaT7qkGHw8PLIc939mc
mfjZHGh9f8U8NaKYRkFyWOHiYyNOWgSMBGrfJZgvVF269v7DHvQr3nMkwxMnortZ4EsO3hHVan5w
IewxNAnjhcCMXAL8Y0yrOmorMrPkig3tyV6+stZL5OeckTzUQ89eqYQSoAYYpO5jzlTrjdn7M1OL
IA+3FJgIORhXRW6VpA0czNeVV9QhVOgQj0tISs7Ab87M4aYIJj/Fj45M0U0L4KM7IMQPmAYV875c
FBBXqay8dX1jgK/jlUgzKYhgkZeLBLpDwfVegsbBeWI9H28ToTSJL9fV0wtjXJagyc9UtcPw6FGC
TCAiaJf5bg3bJcjr6E5Dzf1IIecxtksHb2SzVJ1aQ8l02aexSVAzg/8Yz1prvszhokR1zlYfDfos
HNdh/Cxq100/pIw6nzZLqJ6apg0e0lmiUFr154br6YT47BCHHl5lCvD8jMtci1IEoGLxzMVtXec5
1QzcjRxoS51fLhBQr1HydEdAT3iHS4UjRdlE5jTF7ODV3Zoe+TR2vzQ8ZAr8/W5rkMcnUubjs06y
Ud8ejtSpEH5HRcfIQMiCdUnlw6z7vrcIj//3gwdzna0RqcI+DUlLEjBJm3OQ+T3gbQmg5484zy70
rgs0ACIU+w4yxXh3jqp5WDv3WVybvuc0iVIoDyjaR0/Ib+z4aoMZMsQb0UAxXFVauEkTsXZrGrCe
rQW6h/T/6qydRoWEA29ENVtEbLGzc26XCAdOB4faSDNMXGO7+seblFuFCJ5ZBo90gw/AVdE8JLoi
uneq8QLJLQ1OzDph5ojBDDaP0xppjRfqs7ayPz+rUICa8wYpnabnlgYaQOdpObMaXOXJIH3bgPUZ
Wuwje2Lvs1aRvPXEaCUwRaypLKZTFT1WSHzt0uLY5lnllLMpdb8MxYWoCSBxvUgTOKZbPbD5RfOQ
nyhlkzVg8WFmtyOI8HbeRPn7eH5342LOakWQyFlH3vd8YARfAWbDKrzExQmhCmR1GwKoSwaWf81D
F7qpbvhw007puQsnxvyfUQ7TdFUfMTN3FIVTmN8olE7uMZY7jTpo9J0Hiol7PUarHEvQkwBN/rJi
Dc8PjtJfxnT2CuRGlomYyWBr8iWkoMhlyXjW1rLN5XHPuydiA8XJRqZaXlU/XEcc/rlw2rtPmpF7
DOKLdBijnp13Knx0fzgP1GlK+Fl5I9rkoU2I2gt9Spryfh8nwfL6f0icel9W8kVNKkRcPS0wW8I3
o3GQ3aSfMDIE/GXQhbREVuIKizvUr5xxq7ZAzXTx13GuoU+Gvxg5DYH8vd0hjjxDba29jjwm9TdC
jtG+2Pe3OaK38ywqB0VKtEK3zsK7+WaVEKWkT0rsRTLUk3l0fmHPsEuL1O5UjDmsqZpO3uIVas0u
dSO2gprSWj3Nour1Fce51uDrk1ohqfHGBVYQajWYhvQSRYs3mYVV5hLVy3wwriRL0278OdOzeqC5
AvfskLZstMaVgizlLEBKJXTL7n0RQ3F1xCEhUqEhad7WGoOwwhci1YMkDzL9pC2mDy5WE0ztTNXA
+2QTGhVG5lzHG7/VT2O6QS08e2eDNz7jVPWc73m8IxmzywMxIw/48oeU2JYuNtPRvyXERURnO4yK
+YIuceSnzvXVNR9RVK7ruSJrTx+46HW8KOubt57h+sm5jqNAzCPmc6AMIgj43ej1ElXKchy1NXIJ
dNquWvBwsq7+cWlGVLVIYnPbK7gZiPdk+GxjOfYjxJtS+o4outKbanb8aD3YYdyeD5RsVCBerqtv
lSPaH+5e+iOQvZlcrPxnLFRXXrV3h2rC/1hFe2v4uwgZfbQnbLiiuWh963XLd6VitnbPPqByMxak
9E+Iciw3iPyI+3TtcMdN3/cGwxYCM+jSuJPmlDUYX3Xet6cGkP2PyXTcjHlbsPHpqu7K1ci+Kh7u
FN8xF2G/x90l9PwBIaxcCWQCbJ/KaYrgPKVGpqGfAeK69QbJ8QF9rtRKgPO9fZSUkIf4e6J8cv8B
pKs2i6lltKrI6QXjNfDfT+aYnnnMk7HAAvxIhwzNkxAJovyo58esAKP9VJAGRJl3cob/XRqXWG8x
sHvCAMx2dtlAYNLkmWczsW++kognh5wLbWOD0fyZJYL+6b4nNgPO09yxyximeDxUe42mi0al0M4L
KPf93BBWj9v3frcjWUBb2eTQ7pGUtzfW+ekNA6cUsuBNKH/AjYuFHeflCJJQ+jm6UNevyhTSZCHC
eQgDo2ErlTwmVjlvL+bAeIHM//ER6ghNoda0KI9Fd2oZ0aF9Uqeuziz/fidNNxq6mEwKxMeWnuRO
xGeXHHXDknJeWP+iCd5GcMvHD9/RcRKJ/HpFkqYbEvNkxKDpz0lBGxFLwJgyShWY+Ph3fXdvzVvM
7YhdC3hLfO0abIJv7NjcwDUeKhE3UhM63RSslggFcXJcFBxyNHzlyZemDQZq3gkbcwH4mU7r/i8E
JlXDsz0PSEb71NKtOzi1VFTtDCuEXt81gG8+571RR66stPpynio3D1tWRDlQARV81xgkBRQyGwTh
sHNYVMJxpR6LCpU+LZsRlgSGoITX80L1ndY64g1ngexkn+ruxi62eMwtoGQ63gYZH+pgNx0pHHoj
62B63bVBAd/AjlJ0rBmqsf+Qe+BSoNPF//K9PofttF3qgTseKpme68y4auMJiheisHsVDFKt84Tk
PkNZ0AjxNuG2X608SsmyAXFwB5vAr/V36rKOo7spkleGOhOeIGKI1T132LUjuwd2VZ97sGtasmMt
Vo7patbWALyRn0yXtp1fWWdNto+AUAKh243j03QQX4B5wTpkhx0ax+gs4+0J6f3HCamQhUobyvHM
jPWoLU/61z5rP+17lTzDODke9BTOgncfvqX3D2ge4OgDt/jObvn7HnEloJE204wkpi2wbh3aTZeU
sUmdFWbG7PODtWAzHW626oek19Pn9MrX46foo0mFVXt06KD7PK934K4w93mMEST49KQpnqE9MyVG
0afhPvsXp4q2rRdoeTgn0D+uoitDe1ffl1j9jLiwzbPT0Zai8kqv4Fkg6r0xYRbDAE0yc6sv0n8g
WTBsG75c/IGKq0gK74BVpcDLCzFuly7FI2Xzwh1uxVPxjnKHm9x7i7fq2k7+YeOcGmLgbWfQAS7G
3thNWFgyJS1qx7gAZuPkj9SsPjxMxAKSmJKEDogoYwZ/WVPqY6i8eioiufPcuCshsMVRAV/x5aJK
ReWxz0Qs7wliWCSGr15Um3/Cz1uxJm7xK1PjGk1hnHMWEkGhLePE7JGgFz2mVwRsp8Rn/o1eJJpt
z3X6uVgbIHM8GI1HL76Su9Z5RgqVR5ReXpfD+ZJpkhWPkkgFYS9EFNsbbxiZdpnEhE4EXLB6QcKu
j8Oj7zOksdQkWl/jmPRehYmofows+g+MFbGAZb5s9XKHX9/O1PDSVJXTaFWuQhmca0o8wyvBGFM0
kgAmEYOGG34el0EBMQuHYWtM/QOZluZ+Xsn30qcEyDj8KqL/W1JHIKc/SyNk307DhU0ZA1b1SY/P
T8p8c8k7UUyur3w0daeXJWy5WwhoCjSvHWd3ykuy+vNpEG823JRcdqam11oy0PIkmsuluivwuqRv
patCfnFVSCpfI8I/A4to1hwPBHjN+pVhcK9C6+EJQz9Zfm3gKz4gtzOXU5fA28v+ey3KA4WSqAAc
Bn6sn7/8CIbHQroStEHruTXyzYXE09CStHQa2OWMo7UAVJtL3qVp+7bVuEf2PyzqG+XNsZ6BYr2C
pmVt4SqwzT2buSsdh0FfIX2YJzoVTAp+8bWf+1rqbV37LVblRwhHzf/jsaVfsQS2UAL8Ch40XTv6
S8NXygfYFNW9K0ATCQ2YuHMWLCWiYqHQFThrgigC6QX37SSzHAs+leMhiSCKHFzdVA6rBcRZPETV
LOg0Sfg3cxri9AbkZiu3cZvFI0jGGINB7tH57K02OD1mJxXILjq2v93cPG/5fhgeW1J3PE78PD5N
TFrMghYiMzpOfQdVmhTPOgaiHp0T0L6Yevnpes4ioT9FIuvL4kpTo8q+jNa1iGEi1sFRvvqMacAS
voUesL6NTbLj7h7B8Biy/v2LdsFyQFYnddHtschXrvpxfR/xIKkrWWvr5KozbB6sKkilH4i9d2nF
sTYAponqboFUMGPrAlgXM5gwa+p/kLMws1ZUEOY5tU5pIOmrupXp95onBnR5rAz0VRHuluHDDS4y
LNH09mWRfr7duGWf5CxXLZaY2HVHkVtxJJO+XmYI0ysIwN8svkaFUkNSeoB4VgU6ZOfgvAqnrb7V
q/Cn+JmmMtTDnnrqk9EyOsMlMcaMCEmj7pwenyEDJHpW2eBfpeEt/KcXbSVL7vGn/BWG8+MH6ASk
9LNgB3AFt3VuceI7EKWXJTmBJnHTwOCMkl4Q/uU80QiJOakkHNUmK7R+OyGw8BpQZYiO4pbz5ali
dNyV5WAXWIlipQKC+SSQXL5FtEr6fp8ab6s6/PMBDYqQCvFTcz6K/K7C1XIL0V6B8X7qBNtmeFsX
JzN74vlYceXGfkUxnbz4vCDDIFWAx4KzEfCo8rkIX3IQN9PG8Iv9XRwnhbTKwR1onNX+HmDFd5Ss
aDzE4btWeb+BVPD8bofmTzxE/2c9LTjYoBdcwIreMiyB+Cj+56GkzBOympX1m0Ji/mfg3Gab2xdM
46YZ49PWlpRX7KiUV9Jovsq4d33zo14ueNGpyuPd9SGUzJoincEbzSPXjREdGJEKTuONo7GH/lJa
cLX9rA2cRp39Lh2/ldH73L8bTkSe7cmsvwzaTfOvfscZr5NustIxZv5DMgn//zE3qHjqsR3fgDNW
LZVks2fn+TG8xBQQiDnT0kGayhTvMY8mdf/bos48CRhZESeZX6j9IZX5UKWYpu1Q5ND5KJowWxnM
io69uooUvIXeEhwI+TJRE1c04bUNtQFTRsZKPxGnT3hsnH/adW87GL+Ofc0RJmfXaP6n0Zn1updX
RNLz1AwxT32Ts0tOQ/mubGq+MXKz3nEEuGZ3aESxUwDK2x4PrqYL/rOt3vBIpj6wU05vkhv5XqeV
nmw84E41Spii8GfsDR7JcDaWzMpD9XIs0tYtxWcsrW5Pf2BcQe3nDDZ51vg1h2aU4tg1+lHGUTjY
npN0W3wNEoowqUaZ1k9+syFly1G4C0nR4niLz2Ekx2deVLnm0rlNtnPPfWFK7/0ZvbwqUPhgH2q0
Tgm+kAIJ2DnA1MaUeS3i28NNJw7lmnJQZ1AF/MpxPOvNmcWqjRXZC1iJiM1evYylQLLorGhbfk9C
B2rxWrzSRGUIDSvY0NgQ+oVqWoDiSBxyiabkKURPrsBK8t01Z6ihwkWGQ8INQh7fkaJZnUd8ADu3
nVv1rxqpm9ZeKCBFJtLKAiBRQhDHW0jZkA4hU86KVBD8/rkf+6moJEsi4Etc9qpWTiTNEJDlx2e1
Ywh3weK5vCd1k1opWNnU2X5a0cjiQLzqp1ZYwUKCJIBUp0g64meJSbZZsgjQrow6/MTvBPHC1RxM
SyxfAoDG2BEa3yyRSZPuasczd7mNG7QaP6idpP0sAs56lmTm2HjPBiURgvLSRxm3UwSqnQYG2pRX
S4cl6VGq9hS+5HcQ36MeLfmWtfFKFGwzWAT4LewH/Mfs9XJz0tPAFhRMGKlyHzZokeJhemPUteuR
rOS77ZsbcKTtYH174bpQuLsUft/UrKlRJ0M1ooE0yxhXDKhbyD5nHbohgx20/prf/zflAjhsQiwK
pgjWWnFKm/3mGLW9dgMdW8BTlxmvu8YG1nKColk8X01HaEvr12kmPxZjWf3x9QI2czvZlje2vIxl
LC0/2ON8AZ3QLounztbapjzuR9N0bokkk1dkEXs3iflaTin2yhKh8Ph0S3kPF2VOAThIwfbCRUiq
x+ipH/JbvUTnFWWiLVlUZTRMGKioDp3PoOoYp5SqJneOTwZ1jpZvmn8R2kTndGsqs7MIOX3+8g2Q
0ZcVq1XcrI8FXqycgq/eKiAOYlJPO0bjoASt0QF1K6VX8OaoY7lQCIDiIDY9WqTbtc270kI2ai+/
ojTjlzbiyapAHGtVZF2urwa94k/Xr8u28PHu+sEZUVMdoFmxLSw6CAIqcAr5OkLQDJxpJuW84Itv
zJUofxFw7A9SiNMvhxvAfxJcrLDA81o7/LHzCErKXjp2RXBsJRHLzya2ZA2UaU4taa8nMH+7Kg1j
DrC1+Iqns+3ZLKTxcRz3HwyScTGxRUi0sFvjYRtzfo0PJLPM1GNntLo1ofLe9HgrQNf+df/iaVwC
NJX/WGgRZDA1MlomGPPEcCAQqo8pDWEioWk24ipTMxN46Yyje/B2KZ498JRGbimcs5RuZx7ULcnp
O2lK/0wVblvANQac7W/dPkDHVUw83WoN5Xetu4zts/AKmTZjnr3rjd0y9TWVvkye55UpQIq3nQZz
Ncl+V0zHMhS+Y/Yli4MfmTO2rpF/sGjDS2s4Cm3j+Uv3MoltoxyYyXxcRDGwe/c4GUdTtuLScogQ
QG+/c0Vp6pcBvJ3JWJW0mQJN4xpQ1ZbuEy8LuShrVHtkPd6cyXEotwJzzgV5xtn4FIosjrVBphtr
UtwfI1ZiouZRi0v+is8i22m882nuEa3nctAap3mXVmXbii2caYXLhJ1LhdTUqjb4mesXsw8lzHmY
uOzU9AL6CLrmHh16X2Z8w9xWEOUDAuTXSykLd9DupUXp7ok5NDO7r1lki/K4lecBnP9QO4t8mjgd
vKpEn5f5B36CSYwb6KcVi49kivY+Zws+p1o4CoEWqJTN/G7JRybTa/Ree0dsOAGXfYpdsRWPV1n9
FsMj/0TbH/jCLhYJ3Keta+ye81PiGrTMcH8UUbGrbaFbZTTcI7Bth+s8QTL5F0TDSR5JTZlohqtD
2E0vuBRoMBhjRDqNXrcAINgJC9w3Gclw+znArQEDsxeO2Wvm2s/efuj4s9flyl1++wM1e19yZHwY
nbXcdqVZ8e+YR29S7K4yAzd1B5X8nXy4gOZpQww8n5iKC++bK2ogahZLfFq1vZ9EnPIaLcOYDtK1
TH7q3XDg/0ybF1lSd/dgFukxnqVDwpxTfvaxpnfAzZgUzJe57l6d9ROFbgmqXELugw8zP958mmFv
H0Je1t3Gn4SCZrkvBbFMUKX31K2gt7UKEME43tHj/lKuAWgLtZyXDRmZbArI1ru29x8UesihHPiZ
eUIkEelhrCFyz+yxHSjVeocZxmlWYmttb8QkCqt+iP42I1FvMXdTf+r9awz6v6Jdgl2+4QaEw5X7
WHcBijjMM6qlGak+XkJcj82pBxrt30b/HmOYHg6avaF4sCQMTSJH6JmNg9GbWq7B7I37C/pgh+e3
MYTNyKQhjI168mJxO46b9Dsra62nMFg+ezXQu8/OGU6GpG1cNcmsvFVY4TnusTUuMXXeiht4T4Ya
i282bcfj6hsXFTl51LJ3Kp3mpDrInU61TibrfvcT2y4VpsN5h0TYm7TgMQPvuW73ENfhuvdr5HuN
gV8l30FdoyR28kYfh0oEXtp5Z/KYwkdVtwUp5wVC0D12SU5KfAj3e5hQwcH6gtxtVTt5OSTVgq1s
pBzWddIwl4VFcu/RhefSvwqyMgb9QZwSTJErn+MddrPSm68QgwIvx+LqENfRKK2HoK8wUwTzVwy/
W4vWKJq+wAVH13o3w4qD+vOyWynD+37oz30CRb+i1+AiYMn1ynlrjCkAlZmEgTxg4zJhzbQZEJfM
AS+1ret0C67AZR6xeTSnUadBzvToR/wrTcOci7QK9KVeE8xtvxEToByWIb0RmLZMN49sKF7+JABA
PXygR9PjNOQfpi7R8ZzDNqak85WwKQ2ByBZ0GqoAGDEq8gMLuwnjOnQ03yJqwUug+60QZBWg7udL
EcUSpOaCZZH8fpHBAkK0QZu6HE/Mzefo3HnOdPr0ZRtbHgJYFMWhrZhSZroXjIxNuooW9mPsBr87
PRFWhwBgggBn7vu135wXT9hxzWcss/EEjZiMPLfHUJk2ny2z7ai5q1sq0DQZyUeYD3Mmpb9Nkp3K
uQia+/Dfzxo1aKDMmPedjDtvWmURe3o7nwIbIXkD4M89yvo06gJzuiw2D1SVyLUAzejsvrOfNkFk
CGke6CTctZmNAu/sC618f5/ECY93S2e1BDx3s2SBnDV9xXu60cEIPMRYJJPy3pTXAb2PHyX2/Heu
6TpsnHKNdWtwy5/lAYPy9xNR7DZI8n/yN/5UIlSlnBVe0+vMmxwAmx0RTUKeCftNUCPq3gOquIuw
W5jx9bSrJoW2dR/SRI91Q1BSidBTvumgQTnDwpSvAMjGmkvq6MbTQPp9tum9QqoS8vWpukyV/d0d
8Pnp5fztgjdxUfxPWwBRQ9qm4uHZNhDY5yvWhomNIeFVr+nRJ9bG7GMx5viaesEO4G6Omn8Hc0gx
JChvbLfdIEKwosgcBeo7nqGxMlJZNQsQGDQQBVbgjYdHJaD36L6NMRbtHWYjpo5HKcFx/0rQXcLt
pPYNbQ1noYCpx75G3vkSkapIx8lk0IY1LJWQ1v/8nKVE8tQMmYVOeHagC+HMJLB6IKMGTT9fnkxE
laPjzlaxDky4k+B9yc9gGIx5BpCwnZ0rBYuDT9r6B7B5Tyy/jWyYo1FLYRTH8AktjEfplZxYzPau
hgtN0p2EziLZT/Gl9777LlA+tCjbQ2QSUYbPshVDIT2k08saEjFaNNi740NsEpO/nZ1wijF1C1kr
YjaH+QPxCUoUvdCqzXnSLvJRIUAlZWn8cXUC25Pd+YA/4cWxbE4EKoJXi97qwu1bbk/y1eUW+3HA
pSsR9/xGoEHqKazMsKu+wvu5tcYWV4rMPIA0Y39/MZEbdoo27B/a3VqLJgCVp7qdZwY7zAKh0SCz
myuVuJMob1WuK9QJfL67kMj96RV2HtlsRVVrPM83LXZimJGNldtklwlzMSV00oLNNSHM8Xc8TXT+
3GmWOm54NjAaFxuN7nVaGjjMTaMt0QW22XiDsbejxMhetWyJkDsgJOnx+/SFZ9IAVlYdiO0Hh/+V
4xNIgUcgU5XcXUCfFsRuMjmXwFDmk41NhNkLa3W6692poGwcGrqkB2blyw+lrIQSbcrvs4UNTnrF
UYG6/LbHnyy5qV7+26pQl4IyTa30SQOvB4RV2J2n2BHYrxuHS72DxOr02iRU2W9faj0jOX34BK4b
hn+zYZyP8HEXqo99IQPUV5z3dl82krQIjise++PtswzfFycB2ej4OAxLqeV4v14TtighWTg3Zz2D
9eZEMVSlVaxQuZyAckYZZmXXsOfMO7c4ebcPqABORoVkLe8FdLs2xoyfRpoTfTYcoMKWQfd1HCEE
iqvHv6k9D1OgZA/gRxOcZfVj9+Ivzk0XRJGw9snUNE05vXzGgNmJ3BjEo5H+wW893QkmWra0I2ew
TWVPfM8KaRQD6qxA+i+FzO1AsFpemOWxTa3KEFmZYuFTmf5rVxgopCYWLj2/6l1aCVuK55L4Nn8N
cXYgbx2XQvZg610JPPYnQ+MPDsziYz7WuYs5CLazln852jabuZOCqZDtzqi8WRJZ6/4Wyyf6bU4T
NmFtWWcAlf29XRsfSmbKKorO4yhoKP5/gGjYov71FXPWistoGldTlPkCORxNQbtZjXu0i/hXO/iz
SpGvq9MsshNmVlnYJ5tiXIH58B/rVXMHnVCG2AOvinjrnzCmjBlPcPqgfQ972ACm4WlYhVhoEnUO
HsuyqwvZCAkAvn9BKaP7zM6AJsIXMWbDUKf7fzfKwnUP8hAobdH/9++PcIvKYOtSHhliVTECFwx6
oWM9EyUCEK8lYP+wLOeQPSanAix00Ao+m4RrIJRGX+c+gVm8kXtebDm3L15skqKveemThIOF5GB7
TOsy3KHFPl6LP7qRyVFlVr2LgTl+YR4p+mMNN6mg7yLKgdeED8h2ekFR7qV65Z7M1yWyP2y+9KyD
4+CyngkpPgHERxCIn+6mQJG8R1pf/M+hjbV+a9osv1fmjxS5EG601COZpeCNIZbxB/iBr/vS+ZMo
v3FP1UY8YrccV5xNKk5OWA0EgKo0RALKD54Fj+eK5jSIl+fGPtEmukFxXOAA5F0HDvHXWLuXYtKU
6KPevJmL8CngE8pLc4nsd02A34QZEhPLhPxQ1lTWGE3ypg8+PAvrteyImdEeHVIXd3n8Ve8Leqp+
h6NdLY7/Bq4ylKe4H/JKBjHls5NZrZbmMlBtTCH6Z5q0Hf57YmsvOkYWZH7zYQagN/926dyWl6YB
39pxrxflXssOIAszBJmHTJaf+n45/ixJTt7HEwvFChKXFCBc9F3z5JGdtF0hQZtpPjOOvs6DK6gD
tYsOZmm34ruXgUUHq8UhepUj6ugwSfdrtIc8i5sH5VWfcLiTmr8ZfhHVomKau1Gj3TzBlW4KfYj+
LKqJqitIaNJq62opUcLWH01cKPU51xfMEjiRu6xbZffM2bLB3TQ1HlTpOYgGKW3kmqMTUAAfLUXY
SVpl7ddl5E0hB+9yS6Uf9ctY14Rf57s45ppPSIAXL+FMfNWoy0ivBGoPAIZEfnBVSpAp006/d5EP
K89GB6laLnM3cWho+c2NOCwGxQCJMYlJLgjD1FeQTmHUqvnsx4np/jVNxmJmL4e6uULAOIs1oJhu
VhO4YYlsF5WIBi48Jx+CRK8hafRhxpC7jC7iReW+ZdqSKJ6w6W/xaNxdv+zTLufnSCOqLaG1MuDP
XsYS+okgc0wWVEufSQ3yGJ/T8V9gLDVlSRvR1ZjsIbLeXEvfTqICqUFfLTAQG7P4cvLyADWQKQ0e
xAGxegtmP1Ydcnj2CpxqGwVpTWqDWM2YHh6HmBiTYjeunVcHZ33hhDefrtmAqcTOsUDB7OH9hvSq
auQqvSOTFf2FUb8Bbv3r07JPfEh0x41jFcUmU7rfM+0DG7/Xz348dCsfEl2iqcgVqqvGT67PUoMH
AVU2xPfX+1fZMiZI87hz5ARJk9LBnknbkGHlezliyYIjovetWXjvsptfhyeCB9/vEGp7mSbxSTbZ
Bsp9eVasxKq7vlDUD5rJUiXj2MwXWyiHYqlYgE5da5fPsgIZpNgrbWikZSvJfpuUjSEoPjo7kwZF
5z62q1Plctuo451HNAbGuGA5ByJLCONRO8a8R2/JtSiFV+9XEaMNbY6/xi9rkd+Ev7bIuzRKXqmT
eKU2/g/uiK4LLuao7oOvJMIyKeOCw+4Ms8k1pltAzwiWfhYzwQtp02lCw66FA0fyt701FUEs+q1q
bAPQW0CEMa5q9mZlyIuBnGHtDWXxNpuGIDcOTOqWe1ExAKzEQ0KLG7fiGnTCoJUNDQ+ESsNu2RFE
xz4s0XV6OU/97NyP9ShIpiGTNrz43kym+bBY9J3QexnWuESk89AJ+cU/IXS5H9Lk4KPsqgBQWBRN
xP5nwS7nG6jYm7Y8HEZa9ooZZYibjHsdtHfMJCyD6VTiKI2t9x7KvRXKrDMNxYdMANiQb5B3oiXL
v9nqiXH05Wp7W4YF7WlTNju1qD0znfBuRLYhLDzejegtJgJkzyQaippAb7Vszq/koPg8KEYErGjK
9AbLyNwS5T4EDEudmMWbZhUS1B453cXCUGVllvUg9cJufqp7sicTlMvcOhyA9LDehMphXX8n6782
2EdS4f5ODYwsdPF01WI2p0Xb0kQV6xPmBdt5SC0MwTMBHgEqsX3smsmVQTtGzJ5l6sLH66UOCzLB
RL9q84hi1aTmbHyKNUxRdUIZBCLyp0QJKKqGNALi5ts3IXETKDakZNv4n+wcadfNqhBC+3sn2KE0
wdFdwEBFaywbkM3dITFehccm7v7KYkvUgyejm2SlcRiFUXJ0cund0ukj0V8+aP5SVad6/PTpXEOO
Ou6bCINsiyuOjJvjg7TkU2FflQzMUx17JgOEaZffbCRTtXKQCRMtb1EKeazXC+S1+eTlIrwCXcNd
HOltZlsYo0A3M9lbLT/eLPWpuBwZo8KIbWxctjrSnXMDs2480vfrunSBXFhm+Z3iQwKvIj8Of6T0
LN+sDsTH+S5FDOuyugp21hA1wVQZ7gsjgtt6erA5u+Y+hpE3q7P0SLRe6LLFLqlT9moXAQLFgmS3
cxboHD3CsM//ojhVbPb2lbb0Jzf76EU4FyCMM7mQLsg7zqhvKA3cAyxhgDCBe+kgdwe+BV6d3ggV
9XrHTkKe4xCAMXoCGhrg9MYRXmtUzWJmfcBlAhHhC56/suf6qcK4GprqeryWyqrI4nYu1JHTiYqd
13b9mIaIDOh6EFsQ1III046FrU+gVtB4/WCX8+YS/JhFQnLDtvjsMcxXYzM5kxkKazIW9SaqciL+
UhXZCRi+Z3pTW6WqkRbty25j8uCkZsRQtkW1odVQ2YqisD8YDtb1anEa2Pv9fH10hVYFAGO/PjQl
EbEx0lsikkO1sqLqZupRhm/TRh+34Y4ndcc8gQK7DOnWX+h2PTdbEUR7fNQocKfO6iJr0ZqFX4jQ
S7o53FaCTSDqWFPM1HQyS9XaoidD1vGH35mHEuoqQ6ilko/9m+yJPwz42/0keQ08LTkuajLr9h94
QXo12avlVUFh5y/jIo0r+ExwK3Q4xwyQyP7gszhXoMCxyhY7Mv5aAGaHccaHtXZGN8j5pwW86Kat
S/VvzZoi29XaHacrwRA6jcEto0s5HAtAb66NedhHDZ5sJvEgB+3BKDTZ2TtvFs3zlju6DuRMXLHX
sEhw191KLpjNTYJdfhc/HqVHtOmR9tJ8jsgBvB7iGkBkllDY19VNIhMc/0610ALtHV1uFt7B/M3A
xKlGiEUSeDOn54iPa2T8lB/rOxN2W/3yf9lweW2I1PTQKCdUJ/8nC31/mqllyLhNj49tBR8nWq87
1ErllylMg+YuxOWFK0SFI3n2+dgyoasfY1ZS9mdXj5LEhCJkFghMJEmSLZz683ozJ8YHjmyMrOQM
KBitaHF5tw6FKGLElQEyysGcVljF1LL4MUGYPR+7zAcL7a8L9ddoCz2OiY/hu5B/msug9nuHw+Kx
PTXYn9SmhXjQsuGFEnpUCLY+c6meMtfiBcFefOu/in7CRuA6nCNNX6v2PemBZb7LYuakNN1DUXuf
mrkfUB7Rh5yZzUymdKhmnZm6B/6Y1wmo7lDlBnb/Eq2AjM96hkV1wHlTGTVj1JysPVTKRiTcN5OM
oHp8qfiw+Jd46Y71f9H9oEiRckE42SMHu1rzj4IB3aH8u5qWDUWKQeqMl5RbGXMwcCYhtI5UaXfL
5lxHUR1WeYvk0FU0eA0s1qW+/lYkoTvsa1UAc7qwZk+K0LmqnfHa4bWgg8lZPIWzSSzo8J36DFzJ
qxQnuaY3CGLxRHRuIJmWZwI57RHzcMtf8jsYlOe2m2iJeX55648WalP5SxngOhXtwfH7MMYeE0C5
gaN7WWC9RCUXFgcb/3MLCIXXhsc7NMq9APdNVx2GisdSHC4S9IjGdNaYe+vTX0VHW/C1b0Ach1h8
1oQjAnqi3RP+DtnJGyh6jqnwM8EhOYRKK0SXbHP3WvuDxE49sGKx5HOuFchKN2pwcnUhdL/IQxO2
iGcLS55MIoP0ZQgkELzzrPYKfcDw/o/SboY2DftOyp4pxDxf4UiLDDdAKoETWc9pzQJq/VEebSSj
LZF+hfi29f6t9yeI3t/z9ChZH/58pyzWOjZLqI7RHr26Sxbkvvg6/yzvhudBWBYbz1ZPZUHuvvTF
nk2r+h4NnHGYlhlfUPU7pQhtGmXSqlYIpkvpwqz8NBpcI2iM7dAS5XWa7t4qYe62ClCWW3c/eC1+
IcfR16PeiGWJw4f3Pe6mVmiKJm6bYd5A52OeSImh8a3KsjP+y0Jm1RgMc2b8cxBYM7ciGCTlATa+
pANKQa+60TV3KtuUxi+2xan4gQxO+zv9R7+3NP9Nl4xFK+JvmHUtnL3hEc55FihDVi8VzyvzJnxu
zq7lbqBoZ52QgLB0NdRazzU22Ht57hTD24mA8eM/mRMKtGOMMvwinjpkL3zPF5qGkiqBkqWZr6vx
1biigGHY51wvHVUEfEQq1dxE/PyqTf1DSG/hqAMmPCLYcdUYCOwVm9j2BFTLASZbKgobq7HybSWz
9snNWoMN2IFzsswk8VN9jrxC0AEBt437Siq0ZeAbsRqOeXXRV96VG8lgljwWmFgR4PRPlKHJicHn
pVoDGr3KkDNBVkJzznZT8wSyzHP0mEgxAutb+63xXiTAOTvYPv3s8Kntp5RQ7nxIEVDkC9zzm67V
PplFdTxoNs5v8NAqYLfVZGY5s6vK2hS4pZw1v2mTCxIXVipmOjGAm0qFq8p68b46RV72Zv03iFAo
BUuc7/piAstG29LJ1DcxEH/ICKBCRb8hB0Efr0S3JminvY97Kx5QdTI+i+8IU5LimvRaENdYCXdG
YFJXwyaDJ5X1TKFd41wyJTu9kG+xvMohhm8MoiqHoFP+rDzX53JLD3AYDWHOFZmSN5QN6Usp4hkB
j9USnfxFlJk5w4YSrR0f6VFY6j4zm4FkS9QNALLEwmC4qDA56q9G+d4GvJZRA3lPlu7CwSecISW2
CBDEkLdv2DmiVgrdXlov6NH8OuFaV/FFIxzowne14ca3U2D6QpPzKyy4r+DY8FRTclsVBdcPL1v0
MpILRmTV4tfjH3ykqsmY7aD2GU7ZsnguDF+u1njANNXqShNcssqsVT7rxiMzKERXFrJbyGDbaKXP
mpezWHmifrMchmjUevj0YcBIlXqS41gkbMX/ZY1bZBIX912LyJcmiekw8bPyonwUDbl7UMQ26xIK
mKUo5YYJzdBvhaJkdXMAO0NfjHqXSic9ojjUQeOVgLKEs7yxNRELcR+OXelN57lraw3gikYOIXgI
SoTfhVrt9Oqlga2L0Naz5KSymq/COfI+3rb5bD2xaDQCFLh4n5SYBWuzMv93K/hmxHbHH25csdsK
Ua1iK/NLzOWP+wSNJT8I3/0A7qI0knp4MU3kM5H41MbSA4ivdK4DuE5R5qwdbWfXuCFm9s66EbuE
LmTbAETZyx8Qd3F0ytUJdmgBoXcwqTCSk4xpLg/relkXmExLphAKHtLhxKYQEko9px+z1ln9W6eG
+J6fC1+pWjJ/xXdldMtC1zFbCJSAmWfdSQn1ZxR147KhBlsulA8sJ50cWIEnYnlkDrucub+89xBp
o/bhgvdw1nzwlWDJMkOsdvDpgzcZPDzBSnwqcL7zHjMDLiD2WETdCQLQno3SBSmzq04qOndXOJYr
EgSrmk72qo0hRa2KLxe5ASnyaonB3oaL1hVnxJLrRukMx4jFhoIt8Oy9KKeG0WSnkvZRCJycRn9P
qSz3QNieg8L88vznAJ0di04cTeRszsZRgfOVV6tllCUxPLO9/ahdf4CAajP2yY05yWVv40BCczg3
S8RtwU0erQk8WN7R8WP8Q6cDGVov8vagRjQASyR2OMzqY5M7LhPF1RdgJe0TRwzops8n5pqYReZ0
STH4eqbSDBn91LtWYUmAi9d30n+SJBfVmn49RYIa0gD9vplVh8yg+i0aGrEgO1ypp5B2WIW5oWxO
rWcIKzupXyjT0QUDpjcle41/0U22gntzeYKzoZSLDfclPcl4jJqLz/E9+/apt0HEhlVqVy0Tm9ON
x1eO+TXneZfOjt4625PcEh17MBSaoL5UAGyf0XUIvbG63/xVrq3OYnEUkJwTwVzAZ+8ZR78foRgC
huRajrVwcjoA2uY2DxfbbvY+/MXAJyVCgETJOFJo9AbbPdByBTwLS/m7y56I5ASnpslrehR+Sycu
9kqf06xJK3TQt+xdVFfbxJdsmnOQ6lRQDyYAzconnr9emDrVogw/vsHUVbWkHiAFUcYgMqmHzBo7
XbC2JCX6tiQ4rFwxe5d6wmr5DHEqTjig+ggR4nDLCBJ6iijn6BTYwKROEEmXrgtzAKRh3IXO3qO+
rwppvpLADyG6cquBSC25l8NFMR+kC6pvS0pdkF8j397Em6QE1Sl54DDKJ1GzMUrreQFMy+mPrAut
/MikxD/zI2D534AkylQJwWfJyppHF4ygJ9RZgLfeUIlzAxpxFByukP3WFL1WvCA6btwC5+fKoVB6
+Tg7LCjvuZFeUuVb/eeCeFdnCY1Ex/9Gn4whH29wYAWSnGzQYQr7GIXw62kEcYoXSv43WiXTZhAq
XFocedU8Sm3ETtZng2aq27Tcw37MZd5N5mYKZixFd1V17kegvmHp84Rq3rifRZ/t7XglKlzVllhf
mTbzCvJbuUVQ28C7USUfuqvcctlk95hxBYPuUaDYz9lapDgOTzyCMbySmaHnHolHXrwbiL7DoUmy
ZLrRNgpo5PPPCuzZ4RsK0e38rgBooQkJN9RHrK/BlRvBiziWct6CgieSg0crz5Cxp89iCPpGEfBJ
HbndZLSfPw++f/owogFrUNRkXGXSGXQY83lpvEeEOfvMKNg63H2qcojx9BsJlPXoCK+6hjAAsmGE
pOYEPj2/348CbuJsD7guwCnCIJAbRchvoWXydDm0b5AG/1jtXuBjSQFYpGxNDwqpGdhiuHb7ZoJX
yKJqCqDeac3xEdggzn4Mb3f+olXMnAWOBxC2kKw3j7ds7DZfLw0DnitYzvX8ijm75kgnq0Sdzmn9
u4M4A7gL2dD6lBTegpzpE83hru+crl8RlS48b4viApP0UfEigcXedTH1vGNnF6nO8ncM4s4MnGAH
zx0WdAcf3Lg0HTWWRQcrTdfdsXoBpBzSQZgDDCRF2Bm9Rsr88B++t5ZKA44szrpsadQ6xqkVIMw0
pVjrz7YJ8WvfGV8mYBt2dmbL8P9aRxI5o4360Bi5WkUn/DQfWVFww79tTY1qJ+OkU+cZDmk5eE7x
9IxKy2ZkNvWSQHe9tqN1abufW2zm2yMTOMEfyrvW20M9bV55vdTKX36LoEKRqzKWeBQJnofSkC2n
2bo4b2QwJF2CTimmTWgSax07xBkTs4Z7m02W/e0+bp7MyW+FchD8PdKd3Uo0wq8w6NG0DjybR7VK
QezvPDCcZpYaZ7uhPh8d7cT06rHnX4JJStAAbwVGmyizruTzCtbEO45TfS8R05BepZ1b4PpovHff
E66roEY58ANp2Tia9/9wZWJIf8/XC5IeqPFEGEM5Q7JhSmeL2C1Cu4j77EEaatsMB0ALt65jw4RH
j5tfAJHXDmOFRadIs+pEzSj4sV7ZFUHlE1ORtR2QjNIsPjkrpcE7OxUuVJ7nhuO+9YD16n2Mh4Kx
CznUaSF44sU/sTCtXqSZOPEDxck4+3tOynJ42Sb01PzIWJZ/+lmBvANHHLtzUf/aO5iJmzHGJdXC
uooYYvRWTvWQBiyLgxPfIjVD9vJFaYjVC4ra5YHw1O3jTWj0S3gTlHmlD2hmIwqb4ys+Ec2iE6Yf
SmEZIqeAmgxZE71n0JY1UvjqyTFuYGZgdJtJWQZjdjzxEaHC6zLsIHh7HQ8xuzxVyMpRLnYeyrNO
1xGaREcqe3LXVQF2OTAYzlDwNuxlt8G8ZtOJl3NJDCyMslIPMCwJS9asKW0iDw9hSXbhH+jlvkKm
mH8DiT/vvjLz+p2yolUoSSGKLGOE51Fl2WpBOfnO7EQmX6jJ/xXGJ0dhRLDOgHNPKKnzD5N8Icaq
OAsu1sUQdOtg03KzTx3RIlaSuPsGQP6JKoNKLIUA8yKX1bYMKH6xFvACYnZ6KNz3lCMXwCLfmUw+
qfC3QFOid+gWZnJb8dSMv+IaNg1cX23XQiKM+/fzSw4b/RzpbZeK8qsFQZ+k3bdw6qTDBKjf7aHE
JbujXw35FUhVY0E4rDoRoItyPzgyZbObcjObmLst5ot7CYWPd/+OH9BF7/THKyHXHCBg+SnZHccz
kr7vAXmkbbE6V4tfX7zpky+2m5E2PUuE/I4d43yG7yKIlld8yo9CFSYZ58iWeHpvf03Z3NXW9xyf
kjXaF3uKUxFjiQvC6So17kosTqLXbrnYoVVhbN5dsFGgIDTbW+o9yx5lrqL+R8EYNrMr6wW7Z/rD
sk0wfOLTcYCy+Ht4uUaEbcztmExoETW1GhXT2djrKqL1ARMBd3EAM+ShOI29d5TH2NOWxRxBdneb
FTmRSSze67PKBNTH0TBCjuTbsAz2x4pu6x4TvMxRZ8I4ReH7WklkhyhTjdLqeKxGsp85uuNmHNwY
j4547/mWcW5KnuOpNY+usKjcRVwLXhJtTgrtbsYTIaOYL3r92mx/azM8NfVb/StJuQ9K0Mru5B91
bZwcaQYPextfvMe1QDW0Oimx9vkJzCgOUSc6jCZOe/Hnwa/y42vw1RTi+UpZWb8fIqCAQE8XL4GY
AZR8y3Xq9wIej19YDst9lyE111kYENtfJM/FRFTTFBWEewkF1p7mHumCIoU8DRaUU4iT9c0W4rFg
OFqNNRvYmW9KAGRbGbwmrfbJlyPOtctSqqRLhoYfhKsk89P6ksAGcs/wzgZ3VmaF+KjQvNzZoZZN
LB4W80z+V9lGLwAgM+N86uqZl9WrP5/ltkoxWjqh3mSK4N0e8xksMVdZ3pXWjabPIeWWx6Ff2eMT
xgQ9+KN8xSIT2AfDyGg6CSkuP/g8qIjs5fWfvQrKsN43uk1Me/velktA8hnmD+O7hv+zs2aErJho
HPBiX+2pTSZUuN+jBGEur4LA0FP7UpVEzFq1f+ay7G6DHmhEzm5B2WMspcNeQiuPaNVadBkLLdMg
DYzX4BdE5LfcOCeMoiJG9nPTpyjYRuA/y5C/RAwEUpF7ZSypa0l/mrGUDg1OuxmqniH2C7UjqBuF
HDBC63T7x6tIUP79lOAlfCHhhz7bYngZyWClNRt8TaPXuGoIvbD3sLDdq52Y5A0bd/l7i4awLQS8
IP6zqQwe8EuUbysWnIiysje79iLL1lNsCYHv9nAU2L1vG/l5TwhFaJKnteQNuNYVCuKvc52cLW/C
41IzyF8uJCaxTtKl9+mcUVghJx4o7Fwn70sZ8Pna84QvINcexI3ari9By3RIDOqxNvRFA+PmQaJW
hytkmPr53MBDCaqCNysB/w4b2vsqUt1bNjSysl5U98r87hsudraSM2d9c6su5l8XoVGkaCeTy+RV
q7NUiTp3yPLwQ3k45nM0U1qCLb9KEklgjAJmBSwYHmThWrVynazAfe3TvMwUzP2+6NHNSL3k02av
QIljoIHuFW6AkLkw99pi42dsPZJdDGwImYRczIrjrDiAJS1JKxmx0QM0ha5w7EkFwoP67BDTxEkH
L1GNh3J44MwZCuvRpQnUAk45XQNt4bGevydFNMOznlxQquaUGHQR6iRGkbN7vqwNUF9F2fAxsh8u
/rjFzcdIHKi7M9bjJD2k58G4YRxNCcxDVkI/ZgtZcjhnk7T8ar6brtBedFZk7ZxIMc4MkbRVy3bu
QvdC23Vg977Qt2aNKbDWHK0Df7857JiQseY5s7IMCvBirLWn65k/ptWpfOeGtmbAReE9tTTpOkeL
jV7HChmwM0ruVQOrx7AX3PTZlaB4ky7t/vhJUEO2nXY6PTBrgBusDAgGSuo44eM6sYNp4Xd1rrye
IL3eLNaQGLk9l6ZX6ODi/Z7W34FFESkSBIVXWLOyZyCOpHCh9cCigmOylwfz7XrFgwrTnKIMB9KA
A5yBHeRqfLjU96l0QfCi0hTmY8vL/NzLhQIfZqq407qQlOBBxp1TkZnTpSagVQfvPr/G53CpW18Q
vwbNqRrkQO5YpogmKh+669MT86BAxehGOGXwlrgsp5AXositrY8Gn9RTmoemSFRc/wQZ1SoZrBY8
Vaky5Wg3u91kxUfLZBeZqc6lJhKpSicSTzBu/JkxezrsdhGyrqjwxRLA5pSnLM1Ssgvoy1dPyGeL
ZL9QU2Zs4sXaI1xC/Yi3eCk/kap4GRO7gJ6bPeJcWlh4BXYWZcVP0gi7oxrGaq+HspLsDtAIOpoQ
G/fgVfFVWdbVKD/Kbz5Tji5dAWrvBYmV8nsZf9o10N0v8xS+dnbImFQ4JWchnn3oZyZOEPS2PouM
LxcIcwwRIR/yxh/+Yly8F0fyYK6f9DFUzXWjrUG6Npnk/1SMt/MmvITVig4VY0YnqkduVj+u9Ebh
pvkLCaVGS7qaTJyuoLbQnB2CdKbjiuyegnj4qNeXDsZA9u70dH9pSzllTovBybw9N7GeAlgw5H1Q
nKG2gdw6sMFL2woiemmFe2Z5hJgLyfltmrcsvQJLZv2VUe8Mz/Iv2LzzjVv9vpXPcJTn3lig61li
o7zjuVxe6U0lkBD4RCZnbNGILDYis960wDdJGT6abwUs7Y/piuBs/DarEoXLS++vUh6kC1C0sU2v
yb49dK7PSRn5eNxyFjy9D3cIOpO8UhBo3d1us7uLOyhvS9JgMD2ccaltLi4LjHPF3px0E3eYhsO7
gIMKI5ml9duecXJAc1fXQSKxcVpGaLJ3BGbJnmL7rEn+oah1S0piQE942X+oev+GMWtq5kA/M+mY
tgajBVQ3c3YhpIMtX3qeSIMvpAH0orNaAbeuUb3mHjaE1dRoalzSOlI+nhCvsbd9Np+ZLhJRC7tc
4tm99uwWuNNS+8AgT4iXlBIP7mOgql9HCeRax9uNrDdgcElSezn3LervH1bf+q28kZY78GCfT2BW
SAwmerS5Aid8IojzlGvWbVv2HsNp+qrOzwdR0G7xGXMVfs3YgLn2cogKohf7bksV42XPu+zmlYcI
+p3fR2H2bXcDBcnk/Sp4z4JIOvDQ/1MYqbgz20/4iFXOZwzRfMmlzXMvW5VTdrTzik1qWMPewQ1R
wt+XUHIKthuJegh5h6Yo0QhKmFeQeAOU17o+4j81M5c+X9/OD5pBqRPXSJLx0vZe1gNWE/sbZbDL
lFyRNRDzIyqMPfP87xHjI69NhBOHJLDhWVp9KFi8Pg1qDJHRQrpWY8Oy4DnQ76KW0GkHwQPuTb/o
2z891VXqcN17Sk+4VmLearn3bU8mvL4hn+0rnC6eXj1De3Wfli+vYCzBd1LiUNKAJpzJ6yRuAMZ+
9y0fCzoQQBzQqz4Ig3twNo1hQg1lv0AvfiOlLw9spAp5SIKfkzpEuw5vaSQoUUcoLFmstADG2GGz
7FtgAi5QqHMAM/hgi3u9+TUOYQPljzop29eSAcfICqfuyswIR8D//1SS0ChARVz2JJGl5OyvFxzz
cPWZ+nY2Io6QCGk4FYr0HwvWCEctIBaKTL6BmiIUJ+0c0PbKV/+9NHS4C2A2sibYMraF+RzqC6ag
pEB972vCcpRZEZTLi1K86GMRs+ETqvVohiDc0JSDf5BQjBAlheCothAdyJLEYmmYmwPhx2PWRHB/
M4jGevRRo0jPgf6XiRNc5jI7TmDkDEeen41SkH1pgPwtajxUeHpPNuADp3sVYMWRD8hKbRV2vSuM
+Dz9lpxHxhC+DFecqQ9HJhUDmjUJRYPOA3IB/NvNgbvVi4M7vCgCaiIsnR4HUQNHipNFlNxptiFK
+0S5jcbDGGu6K+eCk+td+P6yGiYolLDWPe2bnUpUtYpXt1jEV1sVin5+bclLNSj1LKTclrlPakWk
vTDgboSId3eWXUlfpoM6fQxmIetH0jVCgdrD6ONBU2UvfF/KCmmTF4GCcQz1wPH6hnuGh2xDNfdM
IKmS5BvPJl4+oABLjqz5SsHji3BVsX/WIhdb9Nd3aedmr46BpShcNJ8PHAi50GnCD4np3qsNS6PK
qMXNoqFZhHQoIQOtmKulHNJjcaKO4HO8cIq6yTGQ8REOKST2bizX4LwMesOh6fKJelaApoz1X3tl
h8cNh6N5RDqak9SG+JW2D5CoSHzOAQj7/eqZcWsHfRV8O0PVEQgQTJkyDqX3w6XY3zp09obzDe3J
tRcEzbys8125eaLkJqJz9XvSCw2pV9deg6ioQJIKbomY2Ofsq31BugqwbxBzUAjHCN9zZwzxMy+i
/kpG3utN36qkDZg3HpBAN0Kzji8U/HSwKLWW1ODvltUkNnBd9BJLnwIZWHQk7gt8PAbSijLCjODU
n6fJ7o8StFxX9GV/ajmRhkLmadqV0XoqWT9OOEqRAcHZ+HfLkS6b5/UVrfk5Qckd7LIs4qRpnpFW
rv8pFs6ObvhDeciv+lLlslnBBnuSllfSVirsnheHvce5FaCyvTRREINkssEID9gC/6vUdnN/Htq7
bad3l953NKWs8yJe41klr3P+Hgmdqlzb0vNk38rhE4Vo4RR0esPgSjuLTqO2mAizu0Orhmrf25si
tQZA/CRbZ9mLqiMksRnHt5UpvTW9ZhPKnh2zsNYd1kThIM9Q0A3FJdyZDyqRF/y0u9ucZrlV5YF8
tUEGmHNWOH5XWErfEbp2Hpuvj+igFUul8+ES8lg/z7PaVp0DK34F6OP8NSpVBolNajhFvt2QYCHP
S9BDYGiiY90FeiZV7TABYqcRUWob6RhNz2ncddKB306JTmLBuAAhjpY2qfmmlo6pZXkX+U9xTltn
X9agZXvF7C5kqWp3TtmnSidICUbaj+9nlc6ykh3iY7w1iRYYg3qL6t1G8Ck+QFzREEBn9qtJAbR1
C8WlgRZln+j0rQrZ3vSceQLfsFRAgHep3/K4X5Pz4bxShoo4DVNYkv3jcJFWIMaWEyEDNfaBg4Gv
0IvxwkQONyxbylO7KPS0B/SHU1dKQJQuIBIvTaN0lp5vQ/MRm2A9p/K3MvwfPzkcAuF15h19sPkN
CTx4+L3aFhOcuOB8VWxvJnmkFzoNV0fk+1XEMPiwntM1PlXst/Ei0Xfg61hO2u9A7jRzKtVHDAOh
EKjpITY4FupeFAZ9ltVazjQEHQ+3/wFjedXRZB81TUp4Pdu4cKP1Uf7UHY2zekqdeqSBAGVunLB7
XHx9c5BOsF6SdaVn/LqRBRDINMUwBeF6b5Swkn2hXbztGcX9QQ9fYZR1h6Ondea4O6MJ42MZPt0c
is7zB0lA0AckmS+e3dPi5LdrpMgj+SRrZg3I7A2snBKhiCQp8wRKBCJbUZmJonQ8Df+GCYfbUWEn
zlPxBSWaexxztYt0+ovG3JDp5+01DurXIt+4zfAlde0GqUcngSre60U3P61diI2VY+5rHI2bbdiw
7tGtsyg9LQG5e3OGcFNKONTca0nUb8r2kqmvuaBSfws730vAJhfGw/5m82IW0GjnQ6Jj9sDjn2Gm
gD7kvI7Yyc13YBr4KEPSbXW2MpS61eZAzIG5sUI9dHq5RxBVIUYNDQTrlIthvOFDYBDLPcAg5jGG
Mxefii00ZuTWmHKDKOlov4QDjf7mjKrdept+YExRHIP8aagIintJesIBHwPTPhdXbF6s12EIUNRL
js4Qhv4Nk0UBWFfQWnYk2c39HtjsrbtPblV5Obn5nnhxf2KQFxt0AcjUdDQlApERmtFIDVZKELQ8
NZNShYKfBM7FV5NTMJ+0cI755Pqxsl1k5dquYKDoQpzkJ4tKOsL5Uyb2MbC0WM/j4+0QqPkwM9Oe
jhc0EwiI/H1Yn9nQJ6xxAPGfs+Lxh53DV68N2pm8OHmgJpwywirOZ5jBQ7yeqY1HRsv8vrW5G5wX
LenPyXIvGMincRKe/aq4kqtideGOEvCsSyjZ2gwDwXWN22iVFsC8hss+PUgrRYzxhDmX8aw8PV9E
/DhBS8+aXc3tAZVRHa6+fMrIGVXsEqkgu8MkyVyJGNPXF5ccIAovJkpNjmghQec0IM+Vq8j5Rd7O
WfWhhsepWuBz4BwF/b1xdHRjxJVqnPyBFLDR8ELRdN1Su6kPg2yabrmALZQ5h5qK2XFA/vhykfXT
Jh+Ko2fpkwGRKAYZkMHL7+rjtJjImED45OzTwkUxMpDOFkX0/8Pcii2B0+7ofJoxmJjEdcllky0p
Nd9f8MVJEayMcuPJ4YM9hpJHvaaIAOLLR+zF6I/t1iuPjRtTVkYzwKgYXz1UAZ0EeHkOmCTNe55j
FX8juBXVj+UMQAaRoAQkzbQavlu/CdpfALDQVl5/Eh5Mu+wIJizkUygQWAarnmK6AGXzQzQn+T0R
ojHKu8LdVOchd/vmiiCFKcMZn1TTOhgSspUCnsp1BHqfWvagNtjX3qsW14WVV45zZgHGVTGXDFgp
tE/0oXBnTqMxwQ6VX5Lm1BaCkeMTCbg3iVeFDt95gk49uqh0a6QmyzaNSewxmokStPgzvm/s6ANt
y6wLBYVmnw9Vw3BxGEE1cC2jc3DfaD9LMzyrseQrwXxtACP/AIZCHimPVo4K1+8ZctJrPwS+T2DK
AoZbg0paAWWKhXn1PUf224rVxB7ac7VrHsZ2CI1V7sN46QzC55uITcAFBntG/GR0DbxThRxmfpX8
YwFiIKq4FkNjhaUSPOwVTxRtVYtStmdCTN1eBRs34mG8Kvihi9nxr0ZGolGEw0WUqhIINsSzNr4y
hFFzYnmW+JHlBoSOLOZohImLC8bn2EYcMvFbKMF4TKgqtM3bOUGZtg7xD8gR26CFFLafMKt4HcOU
bp9EWeYrvwBEIwrnMT0Gzd5x1qSX+0fI5YZYvcP8WwcoRQanzBqLG3WXkEf6ZdbTR3QH5yL2/DKz
lZFjGef9JDtSsWN+t8rbfkNJzEapG9Teo0Mvr2eqgiISqWoTU2EdE8r3a+ZqavXRr887QDst617u
k3N+JSMVVr0TgIrUpxbZBFkutU9LozoHSYUt4PRWsvudc193FMVFeb1OPjb82fH/7f4CT0HEoNJ6
paPF+qjGYVc/leSQ2O+b5soTUYNvWP4L2O434Qb9Pzn1scrnzoCVYCmocsIN7seYdijp8zVu2z2q
0POEs869bf2MsBXHBoobgqvMcqga/FK0duNPtVhQdq8p+XV7HAYyOLKSWPWYQDs3uaXK+Lf66bnZ
AzLuxxvB2ECE5wXRBKiRCSC906Boz6ssezIeHYOsOp1NK4jw7ZrH3t0lBfGyeVtT8LSBozaniqh0
bWD2Uxo1W/zIQWuLo4mmVHJujY0jNTtydErAStCfA/Gj4r7RhmXyCaS00/Er4Izt0mP1meVfYgqe
QkIMzb4yVWmk4GuyS2+E3cYoPIEOqGMka7skRyVGJa+Q3Hfs5CZIUcn9V3krwRgvG21R78ifLnAF
ifUnLokQZeF8IvFzjrewCHrPDptiCbnyqFVia+ko367CXGqoXK8fpU8mjkWCcT0YcAr/64hLb4GY
PqnYJy4cwtOviQmy0U9RTBgWRB//nPEt6VUd+4RJmxLCu1ThnSPmE95rLtCjSsePgviZQ8C4tYdA
dfRguLHgUFCscE/ENJ3MdSc7EPllE6XyuQXqfrg7D6W9v4AgbHPBZ97Y47jKwARtCpaDQ9QRle83
bU9VE/EZw9AJPSDyKScKCVHW3HzJLbmidq6GoW9WsfTp8Ms8BlsHj0xeb/nNVwL7i9CwFnCtgqG7
x47KdlrLdYVvOs3whJOsXhV3dxHYhYFWZ5q33PTBskAzYlb/VowyRyj9ua69jWpzaGG3oMZVEABs
i1q60wIj2zxYydhRJYdBmWqbnRUgoIEsxmF0noK2QLt6kPXLsmaA+SeXCu7+o/B0OxvHwjZ0x0XW
RYqM6A/VgcDZOAb1jIdge6x1+W75FmsN15LNhSmHW9/y5Nz+V2kQ+rb1miHE8WnsbQCogrsey6kt
jnlAXkIWQwKKAZkgVwSDTilaWvVg/wS0AcxwjgHgGTHTf58RymqU5zBRvZrUlGWFbW+BGbtAlZl2
6ALRr2Ti3oI8ma+ioHV5swUC/Y4uTKrZzylnQDUwwjPy8h7xIQbk22hgcjsry/BxnA1KlFyc9d1Q
xkHYBRMC7N3SSABkGc6gyb/OKecRBPHdNsZZ6v95anmpL7YzXdnyeaS8v5x5SQP2ZPjMlSfkmOZb
uxfg2wGJnSWX3+Si2K6I+eYdrdv3a7j9D3wI5KPs3V5GBSj7hbeOcIsVDr+hUoEfvatSRUmH5VeL
0x9imkQeX2KCSy3lAD1wjDdfu7XgwSwsHq7zSWzXtrqmo052i5eKW2F5NjVPaq0CbBulOiID+dvF
ipiLXC2xCOVkOtvcW+llXrBKzr4bhOEoeRbiASxD3GYTV7KKtc0yd+6nGmmkxumjMZAYieqHfGyu
7P+TBKlJ5MHcDMn+0/0RXOBdnrrWw+v4sJ1QcAEPq48S6AR1blRRUsCWoYD9NEzXI9c0/5Hx0nNv
zTn4cRck36Sg01z/BtXK1YskyWFU1DfQoxNtfGIuB0QlWdSESAg6BLqnAfLLLYNOAzQ8RtBAuyjD
kXfKj51BH4rmfUHMCtsq0CIpcR0RuMiD7iI0HWwT/ro1R740Ds2O6g07liipA313Vp9LHvVdEYpC
21hPP7mieKh/fb/Z4KfT+1gdpZxKQvgAlwEI+NbwJ+KxojAiVAMs8u+7/RCXMRPXmdDRjvgoclTN
l6Gyg6cBXHdv+WiCRR34iiYRpL/UmsOttuj/50r3FKDjv0gHF+f0bIIhld2b54PmRRDUo3l9jMVU
1G7Bhh1njBQpwo0w1wPSVNLbfFE/mUeasZTtFbV55CKOTlG7i0TtUpvnBcuNOxgjBws9jtNA44Hc
73ciJIlYaunkLHQ9/xc1RCqspA4LWV/3L0W6IjAlNyMxyKHzDiOpnlZKQBFysDhLT8RSMpaIg9um
mPUuEe/M1jo7uPa2+ZvnFLqs2L46NNps/Y7fz2JLqtrEDeAT0AXfSyCGcskxborkPkRM/4qDJZ3S
q89xLQKLSslQz/BMRfRnGZh91Govchos9RXv5284Kbw0yHGere+dUiVaaCMxhCQuNlS12nw6aYd4
oYsi9jztGrX5Nv/IVwLFS7xUm2F7kvKHRVCHBBhuaOe2JyyDGV+SgVRsNy19i91nU9+MyWEOLKwI
G40/e+N8IHbLFsxWxCviuCCowyvZvtwgMia8Aw+wAmrp80PT+HBP2uzc4C/d8DSYT92LMY2vsGQN
FJO/9SUcoGXeKCStmIbdYocg2KqXCvIz61afbftkMulEUMwrYjHLzISiCPiUsbX9zB17pVeqLN1i
7nUCkwR9HigWRSM5sneiPJaEurI0rgZzV1Pv51W6H0rgO1eEdKrvWKKqhwHZayvVfR674GQic5lJ
6q2W8Fliu8fXK0EaAS09rTkMIZYM7Cf4TWUPrSXz0iZVwvpTLVqXwvF2kyktyucR3dwThoxXvOoo
KwBQRSr/rcxRccj+/KMWfoX7lN03leQTrVw9NCtLibbzA8w3U/4JG9mrOgH+ezfpnKtnfFXGYctQ
MBdoY04DXdqyojjZar27+8542q+JoICcGGYscVIiyOF4QyUB0EJjiat5lZJU4U4qYexNtWmJM6x6
bI0ZHBXIPulkPojw6rfzgOW41dmn7TmyCEdb/Tba1515dSmrOo1x4KaU3YzKfBP1iGdoeqRYba93
+gtoZpgCJo4RliMKAy1e/Xsq7XPqHE5f514choFJLzqzIs+mk7AR/7Xzypn4rbqJ2NWlWVrpz6mC
+AFwxRCHHV+HZVkfG/hAuaAlbfXHW5JcP38n42jpK2xCLY5oH5XTSwksItUA0Hgn9D7u17NOMh0u
VUWKqDetLASXHt238M2pnG3wGtVFlyQqdXeUY716URKm+dNGO11SoFmEie95tV6Cq5cAfRro/CVx
WYQ0ZjkJcbKT0WzvX2pHcL89K80IgFuModvrt9rwbBGhQHeh4OwbEL9U/vjsyGKQ6SK2oab3HuAm
9otMu/D5m08fpcxp/jPgqxcj795cyiQR4WxT5/VXvI8GveiWwpo9AOdy+Lc7nJlfVVbeHctA+A1u
3KSnCIrdiFxSdQoPqSi6jP2S4Da1lnaQOZikQPBxmH2tmicZuz5yEqZ4tRhnELUtIG/CpJwrVsOp
meGVFrdwuH7DIxD54pPeLOvm6DeB1a2F/za9NBri/BZfaD5OAaDlEoJOhBAzDnxiE4FdjAFyW4xn
3YuMeSAiCHdqa6DwqZc21XzUycM7Azm4wwK7uxzsA3WTbYlDSmfFm824Q7pMvqgT72mnYJvRE2nB
4dTEOBMXonMipO69jC5FWHK0nSIDlTL60WgC7lIJ/5gKil8JKiuuGE71fLyxF9TK7ZJctPoSYb0+
i288bZ4umTkkTvVaj+GhYBLrwyHKL7//TSSKSVMNE42lxBvBj5WWs65y7yZsZReur0SCIKr+qMk9
GfI0uvoWxpwOMzoGCNL+jbaHYb2Zww98rZgflLnu9d2pg3wLStKv7DgdrGiUdV6D3D7g2PfJCO1c
oF0JrysIe914Qj6ToXge2+Pt3em5JWCzGB9qoO8EvWNzetyU8K7+G4kTlMP6jXhIzWcwVfYJmZ9g
JQlOX4ImJMeV8d3rSQ4SBLVnPZnqGYFUeT2C5wkYhNAWkLPAPeeaGQisaKVYomH8K6B58nJ6fqJk
qvxnoagpg4jwrQQYnpnVaVtsoQhc4QK0DlLzKfaQ6pEO0rTMZdMlVkoWZ2PVVXAWfpuMGUw0ZktS
XGtrZAC8+Pxx0iCe+7pwySIwFmZBzNHWnvdyh9QmUpEXWcGnzUk9FLsQj/eMzpEIeEUwMLHCX46u
aKjFWiTz5Ai4TDVwnt6Rn0IEjOp66KfJgpa4De93GZxIhVRky2scrakUrvSn8nEUyDCqB6cu2Nzu
CRUPdc9mapZjwDziUEztw66xwnHGy5lR04UGcga4DeJVqwjA1dhjG4MMRZv6lTKufLzqn/22tRRe
8PtRD4g+UmqYpKHURzZb9XCZd4la2kbRUx/eSQT/VdCAQyJsqfpzp+NjA3jzSUiK05k0tX4N4XKO
J1AGI88i4/IgfUfnZKVefeh3PpQKQ2X6hUnh24rLanRx6yHZetAHPAiZGupHICWlDdwa0lPDPlTB
5tO5v+Ks+QGKF8sLuLKsEhSpdonJqUDgxa5JIPHRrD1+wocSAbM/lWPec2l4TwcoGQJmvLtusf/G
gmJQ1am7eJkuAwwFaabwS+AUfz/vipCh+vEfWNCNX9oqHwOhqf8vlGGVRzOqLIZmlWSWRyAi15vY
RlwCbrwzj/of3sLPIIwnFVT0amDRg5j5mo7s1/K6DfEsbszL+oJ6rhiFxnDePoavpgoILhniLBMZ
W5kSsCJRKgLzOvbeJ8RGWHo9jnmtlNiuRvyqQYrHzaiQ0leumkKfx8TzZEEEYhtyz6vzdo0Q9iIk
cVYxuoPlvM+TlPvD0ld8c4uVqYsdBWX2cRe9YMgMjD1L5oGmVgmG465K0o1lVMv8MYtghO2c1HLh
zh2Syjs30F8RxUOBNF40pl6BW/bG6iuo+z4knvBf/8lsZc6GFcnbrhR7/1qVOZ7mXyYX+SoJGCEe
tkWPeTm4AEJDWBCvN25ANMXWeQXapzGLIEMJ4KV1oXDMPe1P/r63S9lESo3qie2XMxlZUS6euvM+
YOqTaxnA5BjlPDZj9x4E80TmQyFV1YKwLdHG6VGOxFHpSDsjfqZyCu5yscTUoF1YrI/gHyH0p702
rBieUbBW+JlYh1lLu7vuzTHTcZTd5DyXvGeWRFwZl1tabDEQAJywSNp0KH+aE/h/QOTQA67qH4pA
z0o9DLj6iRTiq2regIA5SM48hsrpCoCvf+qOS7/w7Qg3SXXPUJ39EFMc+9Q0wPA4tKK2qhjZum4f
21f5lUZNcbQ4FUlBQHN6LTfwOlVzgH3s/jxc9GBmx3y9GN64nuEAJ108dWzQFuurwsIqRo1DuLeD
bJ0N2XslOIvum5Sr9wPptJQxyY/bo8ESwvzCO+lVFHwUm7VFg7EPcY6I075s02knbxDgxHjjELH8
+ZHuOjlib6mAaWDnA6z7OC0L+7huWjSaMPbfh5MN9D6FYqDAE+kTr/Q/ufQxR6I7mY+62NszySjA
qTxTm+2chTCg2akwWyI4T8O0LJ+i9PNdsIJoNKFHfONSL6jDUX502HdZkG2LkpdmCAaWkD9aYXhD
QjeKnO3rbQXLEDqUY+yWbKBcvkN7He5NY8jThsNplmc+0QtJ6pTmeTY93fSelJ/mhFyTew61otVa
5nFVJRcxlzwMaOaQR+pqgc7MdVAgA9KsP8unYM7yNMl9QQLzES+nPhjpAsTsZkgoQG8dTkSnyOOI
gRuI7EdlyiadpVCPSOBWNLU53rRpWHtkyVDlHqymhglV6Xl3rxHZqdnETwHK16BlGPR+Q827n4Si
qL68f1Fj6j/LDCgAzy2MGi2apO3Qso91XB8LGXPAwYPg/Fy5ugwHCuMF/CdjwKG/kpaMdlKrQxyk
2Bi8zXjEFROoOzzzWhcYewebBTHV8JSQIlO7WOQatvzlIq2Q7gKlpP4C64ZHCD446MquQ1Tct/g9
tvEU/oU9zd+Nb5+3++FJHY4nbpJEJSiBYon061slepvJBKUyzsMCYLYd2Jz+b7A3Hg2tHPydALsG
1HMsAqc1/Xt0OT3sKr70tzx8zQVsZyy+l2+rsQZh29+27ELaty7Xqyiw+1T9K6msHIVvf+HXjzmO
2JPkjwf4ciPz+0TnvVrz2yV1Rb3r25GqbmlrTlhI6OCzZR9wrzDYzrvuFE1zPQWs7Vvh0WvliEXH
eOr8Hkiwj/Ff4Sbh21VjYlxCiNs1/P1MXar6gLwSNoCKF4MiRyS71PoAti7MSJ/ANQY6CJ68Rh+1
7aQoZlKTOvmWPQGsP2JS62U21V+3mUFHbJxdiy4SVXj13vOHKsoQoMCgNNT0r7yCccAY53YCNPkc
EhsBi0nfEz7HZQx+fAjLJvnGcojmZB7gsiqPmJpiY1lDm+LJUaye/omORAJO5dqwVgFLa/sj7b5k
/JlstJqvkWixTId5amwHUkIKK/7LEb3+oGx8kjoJP5J31XPyIjer7mQT+njFXJ9SyINyu0KF7Q4/
hviAUoZyyjFmv2djDKkLu0Q51ihDcw05VTn03Mf6C2dzbJsqOd3XzkW5muqsQyvhcEukddc5OaDo
/+dzK77D4EPZhuLOEb4o9CC+1eIHf9OvMxoUX/wyGiamPqhxyg135/AGeg+h9icllv4+yHK+im3V
LenhFjkqYP2JyY+65J5NH9ICUJRBZ5ws0m0TesGu65F18jC8S2i2Xm8VQ0eWiVX1AYtf0ZwMiOXl
3Goo24tics1HaQsawgEjhobBeCbfvAxc8GsWonoS4W32PdJtcoeE/pLO3ZdKMTJCu1mIx7LvxYGu
VxnYQ/Nid7OF4R0dr9FMzA1ZuuCQjbD3JuUVeKMmDLuGPdADxifD209kbhAF5CK9TNIWdipkfLu3
BwcU+SdUSVhB5G0b6coPnSt3lcCEeJ3mLYtylvmG3jeDD6TYFsZdK12gSWlfDWKo0SxZc+c0y8oy
ReUeWa4d03iFNP8J9sgRrAFAVogd+G7nO55rusPhCqO8ZFd+prv2Qv9HGlY3QJ9DOPfgg/qHg2UL
wF9PZhlyDxtTNK/9PuKiIgLGuWK6PGrBt7yj59ZXcDOgqQ2i9dTDmfIN8XdBwLPLKkVUDmuipzPL
i7fMYlE232WPuexmcuewJNXO4zQKFd1qemdiOG8Bkui8sdMz2BUVOWfUUXJyGUY7r8aJs7XmZu6r
Zn9tX3wywXwxAmz98wFp+Vt2sDIR0PlVuNj3/1PoUC4IZ/YnCRsiRRpTUVrNdGP/1rnc75WltIlm
QwFMi2HMGLByC68wJAMaTTtJQOyK/yh+PiUCK4kgF872+nn91bvXD5v4q5vvwp+kBF/lLLYwy6Qx
pcBMWHjYdu1iIu2xzApKuy7BpBxGbM+eLmoqRCP4M3mIGWyvdD+WteTQF/7pGjcKydkPMzrHUhQb
Vd/ExexolgM9Y8HVXIBSJi2itsiazskdM0xg0dPBq+rja+XN6CGtBOLR7aeorJSzrb/M6rY/g/80
nPYra5rgHztT2k0fg0ArgZDMfRcJ8GKVBM5R1qUk5Vg74DGFSdsziJQzXs6Ypxv+8emzhdHQz+m6
ArdXnmaz5l7lm6RGZwDsQcCIWQIEYAuQwBdqofUlX72GYGPyUgCmikBF+mWZXRshbvTOOBJ4ccV3
uMTLin5eU2YH0GCFZWqAUGjqETJ1kxpvCSSTEn/CLBw/tv310r8jHhz9zW6+nA4TOQdRCpKknxZV
82oTIwnPLBD5A3f6Z7TR96Bfolg3XtWd4M26COh9KiPy4S63rAjy8+uuxrKEPRcGwyQuAoIqeDjn
WmFg9KQu7fsr7ypDcYFatPNuCYhe2/gd/Hfrz98UdSqsymt2vz73CcdNxbN+ntzV5VhlBOYsNUje
2qaXoyA9WvGWYU5YDytM1dKQCj68VSf97wm2uZVuF0rJPcpqlwzIUcadezh5DepuoKNHbPgEYwKG
MZLDFJVLht+5SxFIV19lSwvV29AyJ6JdGyJeJ53xkfagrK0I1p5f4X/SiNlQIeW8ROOvxK0jepF4
1uE8xeWzYTb9wrtP52TJPuibx2tjeIfI3GHHRerDLnpvegAH8/l20xGtGRS9MXHaLvPii0ZTvRtG
s4ayjj4yatI8Uh6g6ZTc2Iamlu4jzuHlYTeurtTAAtHTgt9FG8V8/20JzXbk7TSa8mFzrnO2Y+qw
+iAJmENaa2icaGzn96XWnS2le/8yEBdYXKML2WDgnwAyB75Q7D/Vrlv/qIPkyDySDwP8D62OEyCl
N+M0DjpTmecqc50MFvw2La9VhQDQu7afTO54tNlHa+n4YoTsNJiEAVb74pkgrxiHGjjN9rSuMHp6
m1deRfTn79yE078qOP2opooS65E96VM92DCGjiifwz/60ldastS370UCDOMo4Gr432pqtQowIj6x
q9kCaeZUxhpUlYhy9r34XmMvPEKKFA5rcLEAPlKRFzswszNsNoIfVlay1J+/9U+7LoH2JbEsetSH
nKHHO1bGF6vCU+pYoA7kkYrjzPy+TrOUZO3s0UP9Y5DhJs+X9DdTng8q0/n/Z/xr5ROxmqX/7zTS
9L81V17CkXyrkQjW4nKezpdFFdMHnzbIlMRxxcDnhkqcQQ7T5/uQCscqjyH9fh9wx5fk3mRorlcz
mH1KAYm5/f/KR3u3vocUHWs2T5v2XZ3LeJwEmWIMIYpb5vHLGirJL0a9fw/XR9uEr138sX12vUsN
XBr8GPQpfUfbJncTod3nbQtZBjhB7dg5a7QqoyHQlxcKWHxkm8qIdEQDD/8Nmw/sBPeKpUYFzTTa
+Y+rmp1S+vaW+DIavE1TV+Cqo/rNnXd9KZkluPXCOCzMMHRPDVywxJZ5NmhCkefc8wMyowiioeoS
rrsupyqdeFRkACAW4j/NjkW+WobXIztYbJq9qV96+SA73y+aB8z0EWS8/h0pYb7O8sxBJwFATJKU
U8DUijc4b40b+aZAAFjZ1CdtuAPgPUIgREt2NT1FxhAqwDspbC/xpRsIZFOrC58/YWKsfJagStI0
nKTZieHgzXcovVDgz0EHHIX4yrN+De0JBpPHoET8IQAKPpuFzIsEcACC+s9V2AgazsimFSeEpHZS
wZ0fw37mXWb+IhK1uuCV1qJyX2UHZeIhbuaCopuVlS9zuC/TuF24oy0iPnRXleSimkrJ1BZkOWJp
WiylEFSiDwzgC6Q9kSwpgAoTnt47K7a2+BuIlM6tOswXstLyV512i5zYKb/fDI/T90h+uI5WU2pK
DyX8zLrsduKYTX34UHBOyeqjp0vzIWk/3kP+Xy/xBUT6zzo8njwS3XS/xXl6wDYWyPvAbthiRZxG
dCrbLL217bh2eNl7FjnUCncSkSwUGPlm5jQCcr1HcUBZxnEUZlT9V3J14odfxovG/lKfqcEZUrOc
z7pnwPKD8ySVaVqtVQ3jTR+RsIOM+FYdai2hJ+asrgl9oiQv0O6kijfSji/JvwPVz3Y3HaGU7J9g
MUkzQrGYtXzSA0bHzmZnACkdV+mWbs3cak708WG+PYIyQUdZFWH5951PnLPIvfaiQT8VzkM/1VSp
uzfxJwALniqNMy1hSquhMq/oEpq5LIpnK8wpA9XuhBNo9ch0cTYLGN2Pz50ZF4hYl6RfKHtTA7nn
cHa6ktST6SFiab7FpLg+q7fyE3aWVPzhPB+XeMfeIW46faUtvrF4YMGZaYZSSP3B287kg+JzesFc
GePMSb3w9hCpVLNOvy+ZV18Cd8q3iioWkeR/jalu8/qOj+2QBiZ1JRFUDfNkLlLKHjn4aZZawVsF
gOUjqOCbRZsNPDFhMIyPViwIQJ59QZIWm0kL17nC1zndUdwEJAIcu41PN1+VIqTGvxU2YyZeWHS6
O6f5rvEy4wTTnC7YoE1NdYDhI1gw+0ZyRG7HtbILTQPhnxULWHIM3XUip+g5yGbNtr8Vt01xetti
ehudAtdgt+59P3U6lM1OA0g8bXhAWgNx7yiFkJxYCncINrh5PW4BLXXbLulvSdla/+eeDzB4Gdqf
vawUapqlPxLN1YuXt9fKU6A1+Luhw34+1T/qX21XCgbMsQ/XMwPMVZhF0zrlxpQ29LYMVf9eKFMd
Vm+3nbgZE6DCaiImRcgfP48YenvT8bswh3qo4LEyJKDM6tzijaxffU0xks1wNFrsqpxqLeBryh7o
c5k2RSkYlYNhGleaaPk6OURq4ODzzNpDqGQOu5y/1hqY2u/gXvHGrGb8ksAEQ+hLXv2AmCfKREbl
drwe6/FPaxY44xQhrGirwGjd2V0uWtr32O6K7B0L32SH523WluCAG+WVWDeWUqGYmfAKcVu2bNDW
Um9zisWcBSxKYjsCj34O0QD1HWaDF0dK3ZS52082IiB3kyQRKJ5Ggbn27bzVHz0RTx/jQXu8422J
xFyTcPHF1Knn1TWDboJXWtQijFa/cFmdBYkowhVMs2huXaPgzJBgvDStk3Yd6deHJtO8iid9PV77
wh1sUh9NZ8yRGmP39AKKPembxx+SSehJM1LcYnOUMHM8KhMz4MYvkjbIahTdhhMz79XkqUTU2PXw
Ub37EIc6e4JHmBLxxrXcFC90opujVoqWp9VWEXAQIpn7lM9gk3nHa3qUtE/CP3ODMezV2TWKLCVm
8EruSFLeZtzqKhFGrALsFnBAN6K/VX8fBqRU9Td3je4HGrtQg+ZcA9AVnO6Abq3QsBjh2y8yQaWC
OUmOfF7KLIOIuftiEDTE2pCBiPqaUxNMSG0qIwIKj7oy0GcjXwrEC58zUNZllMX35zKkC75j72H9
8wcWvds9zphUlsQWpPDB4jXrp3Cjn1ZG6UCn6jP8idM1CaQ6rJVZBpSuvZ+YBPiyQ5JiLCIcbs+X
EDpCXe3YaOZfZybkiRZBZd2AbU+SHX5XaDuYpkkBeIADZpsNIPjrRX7SvDAdOKr5HfMia3J2vdqJ
65a4GuUb9hY2dprwCydV0I95U2NMNjD4kmPOMykVyZvXiMt7O21TloxF7x7ZZ1Wn6UfPRAQUOdDC
/LIgexZ3947wW8o9OybcodC6BTcLV7l06NHCbyHefhcMEZV9PjM4zHbNm8ry5riQsNfIqB4Oyhlb
jgSN9hhZMWXE1Jp78JvtLMmk/TKH0VI9l2Ie+H3j8sxtvxKPmZdZkGZGtGrRiqMzgbVsLhvY7Ukk
Do4p8PQ4FecofASaDXaQJQCf508ATjq5NlNSritePG7KkvWXwijWYSV02Gzg1mGpF2HPLIEd0WAC
8VR7Sh+4OjCW87zWUNgT/2GqqtCJrORH91inVb/sKo4lEWUExGcYDqXhxna0AiNMxkAsRzyQcQEa
m1L/F4spvE0jccxvOCQsLR5v3bamQ82XW2yA4dqct/1nodk6qUfnuQXcVPckZr/oI4ucZA3gjder
CId3je0805WD8DrZ0eHI3AcguuexTcZ8nJxY/DwEa5HBXd8RXwOFR1KGYEQbHC9/1HO4MG7JAGhL
B7BtL/KC1l8EMTtNKM8ZEgxtSQvZAWJklx3DDrMQm+PP5HCtPFIfg/1nQiYcGCTJnEVFfvFUkdxr
J5hB9N4HkkpMcMjxqqhrtcQAHnNASepflOq1uKysRK/hWOxAiCAnFM0LVJO7dbOJouWQTTCuuaJC
qGA4toeG3vdXAaw/dUgLOE+f3OnfgEIt5ZP4bcVeXQflASKp7zmYIMPxC6nI4DtW/B3FkRP5elB1
naRTLQ4HRBi/1i3VfMxQ2FssYfK8nTPYMPrG1x38Fb4YpQP0bSgAxNDlYVi2rNCm+dzhIzIuDHqR
jh5mFxUGafq3qJoJvyBU14YMY9caFaHYSbnJfOOLG3CRYa01BBaGw+HR5DuJD7iINFKuIN4Hssr2
wqeqv5BZPON/Fh9xaBdkz7UX8UcC/04SV+CwWn1WH2WxG5iZITQEcwG4cEAG/8cG8qCNGL36eodQ
a9L3OBbu17ys7Nt/+xJl5wxsfa9scqRruihvegMhCP4QeNj7BTBmMzTU0JA14hAZGuGVr2IOIr5B
Mgq9Ci1oQdW4LaePO5Jy9kT4LK1sJxz7em/CVlNomGVJnTiaheEGfRTcKWtFOG/gwzo9VLF69sCD
N6LP9Yi6XUoJTOJCem5qg8jr8skhpILDlGA3eyXITnlNqgaPRZYrrwmKsUNWImktB3lO7ZnBK6f+
xqEsnEYLPZA575ta4KmIUv4K2JeGP0OCa189MXxC/4385vaXkfJA7BkHc+2iwUOa8iZJhauSsqMU
ldU+HzxR6/7uz7bm3+TqlNj8oluDGOwrGbRCl/XsRNHH0K+qLWOmDDsTk276N4L4UN9CTfoA6riL
OkOAq+Ji/P/Tx6Lk6AeRI1gJKaM/NF6TuE489d39huW6G/G0gHxIaODnsE0NqWdNkgqwHVaF7UKQ
dldPH6JAn/azrX6d1ZwDoMtQOfEY+ho0W0JrZy1QrccombMIgv3xb4mccWjbi7xK7tJSPXqQFOn2
0EuAmacsmpJlY63wG1RtSVR/JVw5U394PLnUn9mPzEEQbeWVbsYZBkW2bp5Wca03ODxLspvZfK9a
gLGBkHOCaW2a531xhbx9u9vjv0FowvVWjw+IJ9Hnm0KJg2x9StduV8w16nGgksg3I39Z++z/yigS
9+OkgNo+76VYVO3ZDzdgenOeaRw6LyAdgoyySvmy4CrEtKRZWzvL4Byfs05O/Lh9cm5HsG5Y4csw
0ESnp4rF48MR+2e/fxnECYdbEePuIVhCoEoGiX0MkFmdRmh85csXGfD/9TICFkATReDiuRB/Ldv4
drsyGYKmWTZn2GbmSZyZZ3FgUFDn5TCLwP5dAgu/OfEXiAmWHAqUx7nU0Lnmv+ZMvw3Te0HZwsV0
k4dq/Cwrrz32VSSfSDJSEVma1w7HpPAfFwdqSSp8AC9HRSlhDILO84QhqVPFV/2v8vwOztnYKIDo
eC7jsV7+vbuKIiLUyW7OJe67jMyOn/MVBaN/900By43KRwDI1HkHCIRA3K9qbi1YA/VVybWJlb1j
EkJugJblmTtOjsecZEqVwa8YSpFww7VWJOSBS+JosGMmV6AOlc7Cm1Poo0coOJY8k6BfNYabEYiD
608wIZ7upP5gGuBY2C7afVf1C+jqPZle/x5LAz/IjUkvZzBNN7QL60DZRGcDNnLi9xJ1ar5WyCUH
hSiaIb6+iiOpRsd+ZtXsUebKhgS5IhK4EaR0ppZJyX1wSKwY3W1k3rdS3gBEHY6v8TREPorFBoZi
29y37JoGpblQ8DbkKxDmJDcEPWjzv7FT/5J7TKeJlYo4RpzoY8DCbcTnyOJjgnNEGU42m0NkHGk1
uOJ9fB1UmSrQtFLCl9Jq9oMp0XXSEvGbkrTT1j2ClBFLhNMR4ZRAT9Lse0fkVEc7S+sVfLkwndjz
6Qc+B3Lr3Ys2euxb5tXVmqt9Rt5dtv3q6zxDN7DV1fW8MGYYQrroiwKfzl6x3RTuo6VwMTuoe/15
rsY0JzOYdw8swCkk6rVLi3UoMBu7aUotqTwnoXX/FFzwKVGQ1aQanh1PEkSuc6rog7qA1JnAWf2P
AK5n3VtwciNs1fdSDP1UuoKMaAaa6xtR65l6HGfVy50X/lc/NrS0EvWHyy1JIStt5jANC7VQJQlk
4UgbSfYpZfDuH1vlgY5/FPZFerhWAdEcyzkEAzXdl4V6Nzz0whCca225gO/O9JEMF/GGpzp1nNOF
eSj6WjTmkpIVD2C/6W4f0iiqELOw6JlxFd1+5wSOP/inOcXDeeaznd12Kk+eZ2Qnv4o+xTLmHcOm
6jjQiFkoMpcCvntXRyEb3uDgHJVoAg8ztgM4BfoUOqnlOiB0zyKMjeUtzOLknt54pr+9Em2SkLYJ
NnjzUsf1hhdXiecZ4+HGbJ64kxZQr3FDaV6Qa3/QsZM1E57HS4h9BVKSVPlgZXmam8hUw7zdsiVv
BMB23yy8d1p2QwYZY1gzcC2L539nM2W/eDkpr0P8DggctC2r+xLBOknjKhDIZw3xMLYxK6fasNFC
zLIy/NguZK8TytUHL3uKs8TIBgWtg7LQtCB+kKbbkLEpdkahTUqYqc//rrSlrjn5WAvN5CIVDYKy
SRiFeJi3wSjmnsljtjN7pVCXKb7by9q7yjRcSYXyZeJJpytFAcm1uhC4EJpz3+DM9ByFARnvuSnA
ZNjRdqsCzijBomDqhKVy8/zKalR43ibX258mryZTAruoOAHO9tJ7r3PI1/gXnKZCxY40kG0gamQv
2a4LsKUp/RBt1tQzKZXZcEsXVh8KbZ+tKgQ0vvZLXza6/lLuMJPb4iA4mVnisTL3tjeoCxSqsMLC
ZkHGrc6J4Qeg484eO2cUaZtFtAyn8OKHbGf00hmnsD+IcS7qp02NiQBdBvKqgdaKOaYrLOD/uwak
GCn6kh0rmKgDbQPx5vgZQ0fbdEZw+fOHRuUhe4T4uQKyj0c7Y4OkzoZg/pA0+WRQjRkGVKzFHyvq
GIExvYvYzpqh6hAY6FsecO/gjIpj2XodajTmNK4YCLizVd08j+1Eio1yJFCr4YLYcX70fR0pSFQD
/nyDefcAIxAh7EZZKZiYhxeQdZOwECD5EAVFKsg6YBTJ5U5uPgbEcMasg7xu0Psz1pnu/vGdZgiX
pkIs+mBUkgK2mN0gFsT1eHEqtclieipzbe83IH1wRvLBlDRCL7PpLVxtrM2RyjK3qHl+TExOMzmo
XWnwL7IYDODfzGfa8uSi/sXR+cQ3lJpfvHfl1HgL0LjKREpxG17MPI3RRIbBJQd6Qy+7CgEkIQgA
c9kFwCTZ9HSd1IkpNDuj1zZtWK1q8wrqvuCtJwKIB9ysw9cP1e5g9xgg4PFbKgou6/TzKt9wDILu
seeCrC98GuAvSXmfT3uBhHqgjFoyD9d+qayxzkSbnTA9DGBXNxczgjmzEUDekvU64ZvhNPW47lV/
r0/au9T7n8U3HMj6q80hjZqU2OTVfFhCfZHhYpt0KeAEpdcOMpWOpJZyiq3udzYErsXlE37fAEbs
MYh0qB3PesooQE0DctFqXcwSgSmp4GLPZHkTqDwN/VQIZAlMafCzaGtrdVoICAg0noqUAV4qZ2H6
56ydAQNzHgjVg963bOUH8EwHYR5N3IzqZCN1X0zcpbSw61eSA4bPy5DtZmFihWvWtKZCDgyDTeJa
Rv82rxEZgUvTF/XuRm0luWUezPqkAeaOdQqReR0bU4hJqSNjakrCnnRvFvhN9nstiiSbismRgNXJ
dLS4AvvAigbuEo/MD+4X9EQ4aOpx+bBRqft2z41O/rzmPPW90oH/gWjsfbMz9w+0mpLH7pNvYnt9
Mb5dF8X0aQUEjDFzjyNhUkDMN2gfbSCvMZVfI4MPiBQN0BFD4XQ/kG+jEWmUPuClE1VOPJ9N/bDR
iPFh54OjKIURTURakgDR92K7EQFQIdajoHPwP1z2teOp9DR4fs65y4BEbb4Q1D+XXNtSAbdjEPOa
KGT+pvxHcI2P4QR94vx9hKzZunR12jr56TGs7V4Ar7+pVJRL7CZUhW8rpb0BHrpdt0x/tggTTbcp
wwH4K6h75wFIwPokn2Zuiz3vG+D+hK4x9+xQ5OriPPfeNToF06Xssl3/uVOOUWvr/S6muKEmVF2Z
0NmWAwhLB6E/Nk1demnGWrq4DcTmU2vbQRrdID+Tyj4fhuYg/k26qN3Q2gi06enR73myWdn8QXBO
Smn3ff+Mb/IGV83gr+CUHHNzGaiOrRPf18rW3kIzFd2k/agL0rastFPNogk1gTjV7qT9RuzaGgSo
JLXYEcotlf3rsYBvS2jiULlbphDA5F2KAvKaBBZcXIllzzSbJmC9bzkpjetV7R6/OEajwzpKY1AW
6dCQ/rxrjTPEIqn984Se+j/BGnOEpnlVZG0sQ0V8Or2YzBABFtbgghilNoG1slH6pLb7kTYW93yY
0nGsynR5fTQHFxYrb9MFrmtkfVxWOZnsLz2lm9fUt51z7omNlHaazy8IDkLq8/S8BxqgAbodCAc4
dzZPluXRy+g0X1uuT8b9x669ZaxdCixVDOsfB8WESk6UboTAJFcU07dSygamBFWXOnz7zR8cgzzg
8skf+jbspyRqUIdxyBtGSwdBcP9iUrghi0kn4Sn+aSv6tcy+DlOrHJbuDbDeeX7TiClA5pGSgvR6
TqD+ikcxMmfg7PxwTFmgLtAeoKZWfTDs6QG2GARqhckVTbMiem6T3BZtTBJNFKJ2/0wotgi1fl4m
CCsW6GpVJqk+aFyhMVyCYDg+yhQTO34WShsu9WNrgl6Pa7mLg5Y212zDny+bvEAHU9AX7bjFeq9i
qOrhalQ7q3q2N8deXmjWxh2GNudb5N4gxdLqSNNKr7RZo7AtRMRAGuwdfbEdfYYkYw6eGa5pgMyH
1jggyK+vdma5lcYBq8qJMv+2GomXBY6xLeApXv9SLbzk3R+T23DIqTyfAId8XPUIHb/ZNWhYJBvp
mEozTOS42Js5aYp/Z094tO4hea4vmL4FAOUYHnRxg4s3L9kTBE10+x3MvsqGs26rFF3em6rH9vVv
I2EBbN7dfmhUv6bJgj6IWOA8Otc4ho1YBMDkhCUaaZuFe//UZTtdBPyzHg+EXyFVqNlGyRos5kpg
DiB/oVqgsnWLmKVYdZ9/upBbARvZc8aGCe+ULuxPOP0lfAD4pCkbd17AYcMm9TWDud9eZQzMzeZc
Ui6AVe7gRL4ODcGe8Bvj3kTPKaSXO376k40+CEOqIxrqGEFyJ/lHSvRh9zz4xNHif+G0YA5S/UZL
iW59BZxhqeGeCoQi1f10k1WE75MgrvSq0TMD9ZsGDCml3VERN35Mwd2jpVN29lVdjgdRQqFFsQRI
cn5WzavfGQCfF9QYo2scZU6ZdETsLji2Whyxhbha5Ye/21+0903iZFPD5J3mV8oamjzS8lSEMdGP
U+mmJLg3nrQw1XgBVSIW9k3rdlYoBg1CHXMeIZ4/XrRY2QI0Nypfn6LEo+1Igkaaov9IlG+DQOCg
MQYXeXJIPMRe4anVVVFIW8p9iZHjIULvVgnQQxPg6s9zBqPXLYETFuzCoXMtIxl0T2ugedyxdThs
Ee1q/H/QVuCQNs5V7p94j9o9C5hkf6O0cxYOgANCzoIxRYL1dr8NVE64aBaf7cGzktD+4KlGFryW
EZ1zp6PkQIrKqKuQTe+1ztmAnFRZBCTyJW4kse+FT1LnRN0t9Pd88xrqhV5RLFTGY1TlOUH9Tt1J
Jh5StiVFmGNwFQSg4lJDXw0VN1MBehvC+Pn4HaA4ZYG2djdYf1dPdC6d9nANCQ63nmxP+ky5fGXM
VCwjk/HwY3kVz3dwrVR44ZGpQnxQfccf+lvibe06wMPeJIQghTz6ni0alzcP3vQexqTgSrpWRiB7
uNaGOVc5Q6c3JLuW5g95mZANyBZfLtBvPXFiUQDiYgTQuDgzLQUt5vUpO3w7NdktqmXYjqdIMxJg
ff5hwnYf8MmwIzsF11Pr8SUriywkXqS6kx76pf2tpeMVMTzZXQs/5a3ed0IsMVtgdtUtuG/UKMqu
kt4nVXfDwZUPglz7z28N6hE1bv0RcEjfXKrPJW97dUUQudt781wm/R9E0v2ig7QYD0wb5L/oPnrM
4NdURrUHr7H9IIrOXuyyLmMazd8QZVexTfpDFi4HE1gAPg0oCJ7ahmp3D0yeB+Rh+0NTzEaivGo6
9IAyOIcs3zgBSziEsptzw6XkY8ySvan/C/tn6PEtM4ode2bmAPaHlC4Unq4qLBt6B1qVUlTFwMgA
bQKfhqdx0qt6ZoUj8f16pl+Lz9Lle+zwy09AlAmMUWTQzbNXMIRK+2oSbAgTz0c5zjaTTpc0dS3h
4vqrQaaFuIRe987C/9liv6XxO5VBciS6niEn6y3AKJEUIDaXX4srUbbp6os4dEWu0bNNEQ77nVjs
RtcSf4Mrp01wT0hlgagLKqQ5IbQbJ/97d0hRlqWzZHLFh8oAd+90fk4cF+pnVEou10LFa4pMF2yB
eMKfn7NUZ9v+Fb/qf57Rp3q3fm0epel5+XRLC0tzDBIvZ05SbPS3D1SE/KOwFA7jpbe/AeTmRWQJ
b2IhJoEXEpqIVaw68TmU67PFYUympm/s4jbLJE5Aai4gKMoUFf4BiRY2zUJyPasdOPLHPkc1jXpr
p8NLuD6ktNpLOBe/IGdK0IluesYJig3IhjQpgw41fFYSeJ43A4pdTGqgYmScuErW9DCu4I+AvAZI
3nGlq7+RBBUaaNQPjSJoYpQEqlFkgVcGSe4uKKW5kSeBpfMq111koPEDtnKgYOX+RHSd/BibFjP8
aPj5jSdlG9yVQEsaHbbctjikHsVyt+BFH2Ed5lSslNEK4gF3YSr3ibd66SCWcyZ4SsL4V6jTf3S0
og0kS9D6lp4gaADBZF6fMSgeLa7ZqCoq015wNcjLvkdlFHs+q2duk/mjm1fzwImViNpLj+iPudiW
9syO5s8GdwzZb3Si5bmaxccTZeUpF4YsS/X6CQX4eUJOI/9EH+i1nKdQjaeWMRbC2o/cWyniYOgU
c8jeSEFQYw2qPjw9x5vYXPNJk+fKSkzQgpEU/FJg6z1ddIsqTtrB9LfjWRh//PlHYJjrXNmskKrd
KYfP2tb0n/tfA9OklQ83Cf/8TTa9aO7Ozk5Ye7T8j/wdG7ue52CODp4gOAUzLCAdbiD+mILDTlmS
vjDq0HGNvf52yP3akFyDxWNu7xwrg6E1Am+xIrMnjSH6Tgb7qZNxkxltNEF5JN/lOtLmEpvUHER2
KW7i7ncpJrIMjQeXHZElvhQRcNGSdLcnKWJMFQTy9j0FLijZrewr2UdPh2rLLdFbcQNPoF8bYuMl
KOq6C426MnpXQhbgT4c5ch45fkF6n/clM4YRumedwl/1RxzX1FHBM8lID70TUVLTLal0l0/N0Tu7
sc+/eh/ooD0ujrl8X5BdmDPApuFkZmHFO9T7Ds2CJbw/ZYB8UUGdKhzlt5WGOkbaxJs738o6JWVw
+dX51afGAsiNPA7kbzzIpHKdwO9Z8LqMgL7He4OCYqrZheKgwbXMosX6cywnBiXgotTrS5bgCyYD
/8y7UvoMYZWkjw47sdphwHq5B491nOgNYC/t2ABrzIrsjWuad5RgaVy7+OkYExO1dgjGpEFRlkVk
lbg/LMev0QwuMAauT24sVr1+BYYdktyQKVT9hE14HY07btum0NT8ZuV+gyhnucuSZWRfKPsR7QvH
+z3pN1PYPIk/9Wgs68jPDs10pChUDlZwyf2weaau4xSJxbJ75iEzz0qSpsXvfer0MG/XmOPe3CaP
1K6ut0s8hZyNZl3JWUq6A/4L+uAB7dIrfB+8owPGP2FSnkwiQ39RuyZeeo6ydybdysiHsG9TgatO
fCC1KH93FvLDgunGBnFSXqcOrxbDoL1eJTXySRvPovhETveTpPyKgzAjMIuQgBXA5PFOwi9RRYU2
G2Wg/oURXivonNLd/T7XSdTeqGg+6qXEG8MExvd3mflx9rFS+mXXKyTar8vMiIASFT6M3crhOS8m
dIJDVXbtAAGXoIly36fB16IzdCq4CeVS7gGpcbtCPQz8uwwCY53X5sOlYc6Z8t1KOLY/z18mIXFx
thwNO0iDf/jytbilMDN1axIMdBpji6AW596SyrWbtTm8I3GRspGfLI8X0lQ6B/uK8SE9cK7PC2rd
EwND/0Xfi3x7AB6RpOKLoZJw+B89fnKQGxst1M3aHreoRwqD4ukh8TfbH3rffU1tkYJOuLDzio31
WzEQEZ27osilI2sovl86SqxQdYMTdnmxnljBDzoMe3MofVTcKge94GNeJzeGnpXLMhk/INmKH6Cp
S2srtFUEgV2bdbBX1ie4mscM/oafnp8BfKYZAMsn9EZPx1WjTfUQJX96R9iRhg8YwH2DmVwhAN17
d+cC+cyeHHKjv534+HTujjq8q4TeR7wnoDaMzwkdtQMyfUznomCUOPnOpTV5NG2mPcmIPsRvgp4+
f3+DSXDCv8ZETLtog9BBPF6v0A3Z7VxPGVMMdyzPe0rHI/546/DeyMLRXhPYxhxdse9E37YUpfg/
aCxUAIQCedJiEmakA5cEpnWB+ncN2Wnth61CXnllbVlyeoAES23cygi3FegGebCyaoWYGFM6vKRu
kIaD/5bC93AJoiuj7PC/Sh1r8CIBfPKE/cy5udMzNT1jgolpB13lNR0Rx9TAwyDwMdzOYtd3xBiS
eDAnWJlmK+EVj6ZBSgrmBpnp6aRO3/fvA5NMwSPep/7C8naLKjx0NY6m2ymc+TvAk6jDVrCiku8P
LxzkGKfC/KVIX/FSvMxujUsdIHYdJxs4zofKKqS2eBt5Tw3bDhYz8HWTmEiTunQ1W6wuwxRelSrw
6D1alF+bmTE2uyoxwdYdAVKZ88f2e4IG8vh9saJztWOgVvgLZ6KV9v5MzsjQ+dj3UZwBWbD1n3T4
IAizm8wn6nkpgl7hl8Ho/O9wZUDLAjHXxKsenYoWmXTQmW/OZjMtx5CIZuLUAi8Zn7L0duic/Ie4
77Szall1ibvvv9b21mlirFNW60FY+x8Au9vveD4ZVa7oC2maP5K19jyA4MdNKrt9EF6vKQdGt/ER
ivEXyHF+m20I+IsWHlVGZdFjcbNDvboEVcGwTkePHnYOQNGaB9vo+tKqHppdCGcwrCNNPkgdNd6O
nG+IhV0AiuTpnCYz4L1XHgwAAgBXCxjWYWv/xvm5WeB3/QClQnEQtFH7zYxw+QBiY3qJtJBja9o0
JZ4EPbSS3fpLC5CcfkMbCZ8Q/cblSEhNZmFSje9xxldeqh+XyTK0k0eEqxaEkBo/bBQeAWBUYb14
DsL0c1rT/rvVuAvJVXEIjVHspDOMhPd+1HRB9YjCRi1PyjLm5ZApZ9Ydx10D5mopXeRNB+q4Oi2P
mGObnh3nXgCHq/ZTPqDDE6M1Fb/0opWdFqZVYvzZhkXk31oVhcXhMrqKIuZE7YSCRDqiVoXaFq1M
KE4WuQ5IZgTGvunMEwunsZb0+A7mLqYR0BqGW/2ZuqAKKJd1Ei9pssOLFP9nPg/y3V6mUjAjnLDw
W8AGpp/UW1ob7xScx4KK3eABxsMRMkYlhRiAPxVvenOoixUcVLYpT7sS+O1E5ed/mEjyYPx9waIh
8RzpkJmpoiioQlbKodSix8qSucXFucr0K0YKaPJQ/iIeZJGITBcMMn1URnP0YkunGcwB/xprGe2G
Rnz8aigcT47jpObYdBRJTG+AD8fBPumQlGY95TEjxVzrVFcoJBusIgdwL6E5HhsVja1xnOS0C6YM
oDyOgrYPjSRt2bzsbN2EYQUbylu1eZron3doZdrxit3E5x+XU6GQzv838/iJPgQu07iYab+PzWbw
s+4Y6UYC+vMCqDd89f1YBJevxkLDwkwXt3sSQY8SC7Ppgg68OdZka7446FLInPKaSEL+tZmAOTRj
K23bGrnMoKiPCV4hn8qFHWikWlx1xDLo6p6L9XzZCXqjjSasQpOuBEzBQ8TfCaXKySINOvjrk+2V
SfcHk79OOnIxfZRQvEu7Ho9kY1V3MyZCdeBzOEq4i36xaymxn9CmEpLFIGR9gfQDo+kzeIN+jIjN
Yg5RGjzJFXwwQElGo4ZesibPpGlVoQpcr51gqYU/g7W+fogxBYmyvNneoqmQFvxzWevXlmh2UcTU
P+5NKw4TKCGb49UXqHCUadnmwrtZH0mwS/E7FKHn0XvOIs/NgAyOye+uVTVzE8A+i8GVNuFLxIkA
yaQ1n0IkC3zAd2pu1JFdk+3F6VASZ2rIX93/Eg8Ay6WOHmfb4oTvhAPtS4oKe2L+KZuhs8KzA/xH
7MEY/xCIC1k9yNAPjIhKFPfaZLk0ZvSqDd1eUz55VHaKCSiOBS/rlTpk8cLPlwlw5WQIGCIaCNqx
1Kl6Ine8th6ldHobM0lCx5g88n5enizBahB+lFmMBGJx99Cbad9hgqx0Abz5LyuohAMopaqTC95J
n3nn0wAlFL2vXcsej4SEERoZgClTtB3Xm+Wd0iZkUfb+GLYDkITQ+IFBprDUsGqKGPKtdBc8VLz8
y+9Q7ikDRnGKiVj3nD/ErgHnp7MhNxqwQWWz0kEPL0k9zgItBbWOTuug+MdT3xwiSRdfTULD/yHH
E6HA008m1trCQwIZiDWfKRkJvONzMfEp+CQ7BRAQFHUYOplMgtNoyEZjoOUccmc8y3P+JZk5yqgk
XXXl+FmC4d1zA0aEiNjaEKAcFHPNUIt0QBnFVN3OKPgud6YOpOCtia38s6rfqhYzpHtmaih68Hjz
ME4tfwkDufgAVNYBQjXofYxbxpQjMKvNpfgqVg5+5S5JbgjeYzbIs7T69UNjYY6ZmRZJ+roSsRd5
N1nXOSZFWlvACg2taIutYlKIjUHb0rb0YVC5F5gMXWvKNnfo+shAprzS9bDS8EpHhI1W00yLhkB9
s+/yZmziGwdbCfhTSSWyQFK2z9UWcV1fRl55LCBsRDpjCz8QByEVl4bkwz5EpZHRYTW1rylv5+Df
GQ7FuZxGk7suEOE+HN/LUpD/9tUEJzTWjvnrB3Wi6GqBsEFblScJdDAG30LoqtCES4hS6l/2n0jK
1HN+nlYyTeLN/FpUhtugFOBf/G8b1/b41HeED4JxUVsjTvkjnATxQVbfsS8ehlHMBXQVTHOb5USG
/bEomAi2wVE1+ixn0mkcskrJRnSlfdNVgRNGG08AakPahyiQHEKu3Dq2XDb/6wPMK3m1lhA0RR3g
26Lfbfo6UR9IazU4T+nHbwlm13bOIn8Fk4m9RhzACm9Dx87Cm92su3+fKqSHlIAdZ52GXm41mDME
aVxJ0TFwgpNoxXbp1iR6fkMmMMo4rIqoTiuzHtyxEEi+6VgXo5jiRatHZSm6w+Q3HHOepbm1E8Oi
pbJzP8eP8BIrf+4raSziOnrO6WlTgU9+6yHI9uUawzQL1jNpUfK4S5cgsOLDaH9BkHeSInW6HtcW
2t1FlJcv/OuxsqOBs9bdlzf9tn0xb6MdSfkJ2mtAQP0L3al0uHbY1InN0KHjrga8ukdWzRTgwwW/
bE1Q95mLKdQt4WSLfIlHj2ki8Pfj3PPuJu0vyklZbqlXsw+IlsMQ7afuDeukAfuwzpU5UHqA8Ik6
pApkHdLChwXSDHROdEP0CLueRuvDosV0wnMnv8CYnkTqdGPJq3s9gnGOGAG9x07cwxb8KpOtp4+/
OYCwiXs64FauWxaKjHk00gky0hdrhHmsVACn8FlbpO6C/yh5F7ioiYFEQq2FqhXpF0Rgt4fTBGiT
oH5j4ds7/ovAekXy67bNvrSgqYx1TK8Y29Cqfm9Gk8I5OXwKGgsoQEuFF8Xydhi6RuvqqsFl/FfD
vGLNU5HMXPRlJ7fOgkvA1Xv9XXXV9aD2Xwsc2WcMvjmaRrc6PXO0vP6aeQRNLKFw7h1CwbK2HYqf
L2O8ov1Nw9i7xXhlfSXikGjC9qm7Y6CNDkDprXeAiCvN8D7FstI5JfK2T0pNdaEp+cw65L5tcMfq
U/P59kgjQxTwEa2zRI9uHTJmP94Y05Knii/cFcwf6cZbttAxtfFbc2yMS9KkS4SJ+FlBDT446TjS
TX7vZ4tu9DpzdnPXRxTsovNfXL6u9ze/XppY/vKRl/f7aM3Uzd8JgNDqvqYqPicEnVSdZ1IXZ+5K
X1kFb05DwLNJeq1xltXSpzKAww3r7TIvX4Dei/7wEbrxxg8Wmgh7yZ982sTKsyh4cV+bT1kAeQPW
+ki4F7t5JldQT9m63V4144rnLRyfczNfi5rTuN1lUnUCi14Dli/WeYADbbkiTphkx9bav9++YwLd
4p6DGvDby3buJR7nO3jmEAzq5EAVcaZEEeZttTSzZBswkfrGWYlUXitcTq0bzZ8Fg3zG/8Zi5ZwF
03YKgnO+DXRxuGOjcheli73zHf8Qcs530waGtbtiqhQaZG+BaKVRB6mx7rNv81NABKSXxZP5mrNf
d+UUe+DAa9fyKe8RFoQc6bRQmrMguWAtPJqlW2jpvNFEPs+fO7AVu8y1v9fPf1ZFsOslyZrePYrk
NgCGySFDBhqbsMsv3gV8GHxV+PT8dqrfewzrJBTdbjRQtUVicNTUw9EE5wt5Lj/XVXu1UG5e0ow8
gxMw/bGHkY7RWhe4rOSEwnXRlJRSPQ6u7EnMX7y/XUxJodt6cYrRieE2oxQdgT1q1BlmM3KgnB7u
qpBVVhTYumcDea7IpqMmB+4YFdHkKItpYRRntgcF0vDI0JBYVCi7C6ciCnc9Cfl6DQelVrd1Ue6k
VrNNiL/WDtOm+QVfhbD1FbbkJ3TBqu/0toXJBJxzexjhqO5sGf17ZvhpCcX1uey9V1XRgawjyGf2
VyrClZRJhJ1I4oloK5zqbrP4+/CTZsKI9C8BMzwqsFHOUdJ7H/JuW/T2tK8I7YU2eN9wbVWs2/je
kgxEUHV9r4cVf1eeJRdBFHD4PptTyAqK2GFrTqu462LFSjgmAPPISO1Z+Lv8V7y19w+/x6eLLOZp
8v3dAIy3XS+6Y9Ym8Ntd3z2ZCxCHAI1eFcdvcTZ5tAfGh+za8Nu/3jFaVYn0uIg/uEL7YJq4gfOc
bjT+S1/LjGml99FRCGbUaQPKlUYMxNbhsqk4sbX8NQxKfQ6JV5OLoG4eRRzxHQkeXn1BJIjHd+Nr
fOsFWBAGPoikZFC288H1u1+DObpc4XXQ8YJnAxGsNVkGR2SivxMyW1H8D4V872p3yUTDR8i6emSz
pAL5BUyLGDhsVZxQjINuOV5+eD5wQLuuekBYKWuFTKNhGEcuztpHyGPU+Gw/tZA70NyjiqF6SIjX
qMwknDGL6sGTVO3uI0GLXPy8erFkFDfL+0UZWCC4n+RdELzX946GxeFvzl6lxDq+E8JqCKBIZLhY
VvEAZ9/alzfzur9iNvZNp1fo6na3NAkWr8AebSFvw97eBosvn7ZwdFAAwaAqE24YC6TqjsGEewB8
cg1iG+YhCwNlLdiSZFvZybVoa7vHeKZhMOMABgJ8v7vHcIOTU/Xv7A6nY/m1TcR7V57OlJyxqCdk
CJhmMFNv+fgTJcC1Br7rG/mp6ZlaByBA45228NBomUpLasOb3bDKj3STkmzlaAsO/JwRL5dnbJTW
CL5jUV+6KPeBwzDEsmP4EBYd+xdK30kTu7Bs6qoItjmEk0uL5woNUDwikMmQoyeKUaGPo/ylqjs+
NjxD0IGtH4B40UnTOfbg3J4l+3UvmWo00gI4Aixk6kjkzl1Xnpuzzi2NFmI5CaNU1GaKPq8OAIdl
qX+TvErM28fUdG7CarqoM1OfcmtRskyFVsn4F/KJudEZ2HBgVRpbMnQkQrGi4tRN08YIKZ+4jrnK
2llXIt+4rWu5AIO32PlMSJeSbZazOEJDsCdB5f9gBzL7ygeIfx5ThqkbJp05qT2cfIz3aLSkhS8v
idiQACo5TAejaudLkR/VMqPhvt1fRyM1BYeZlW0+zKqUZ+h78XI9EFkLZjHgyIS5Z1/NdAGIQvCi
CPAIixRxfaHw6R/g9diN0aeaVDgtobdNvPGhD6l75D/Vwxr/6aAjjKHuI0MOrSf4qU60Egi33Gqq
f2jqgXCMSwmsoaZusWirBU1fJ+yPv8bqLR/nlJNqjSm05R8AvyP8UauZ5qfrEJ0hf/1TIu/0Lzvk
XU589SvKyYaAbryedK+BrjpOFenFjMnWgnqMBbDXI3MStP/OQcVD1WNpSMNkbqwyWBA4WlN18nYX
ID8n0SO1a1D5gq3Y6mGqCIV1+cS55AdCYAQQuDv1Q/KTg+eHsX1j4mJ7cVHe3E+AxI5AvaNCuNib
VNOdyB7cl3AI/24BRFlGUZsY96Io7xOYEi+EROv1HOEQMsHmBCwzfUBU06WWrxgqoxhlxzR8VpFD
y6ohyTHu/f3rZwdFkZnHtsar8gHzcdhGdS9Cl+aWm4+j+ytw6ZohgrwoWkv1LqaNaTlJfJsuPP4Q
bfZLAn+PP7ogGyUD5JyUTD6b9PX/MPNfzXy8G+qdQclOD/kt+WBFJ1Mi1j8FeqEd3+URcJzbM6G5
7xdCo9w6OPEPg7KILgNEnr+Abks0hX899TTw8YWZq917DocLvLHUvi27W6uKuJBJ8AAOy8OVqoxq
rLlGR2vlZvPWhk/oxAYp93aE5bxUqBxnR9GbsBNbnuvbYwZOHCjZg2J7PYWJCJzbQKxNpimioupc
lYmSQzubJGbChB3Gruoal7rHXiO2PiR+N0EWbpqJWHyP1EKaW7coFZARwnYdjvYjetkLQQ2VOvzT
0tfB67zB+VWX9dPmVfMtFtyxHUPOkDxnz5BogEhNBjQD6IRMqJE6w4Ukop/VdiFsbA6wqsJ4UA/R
lO/7LvQSzPRtU3mAfkJQszreJ69g4bMBqE0yDC1aaKqh1cvMyKrH3Qjs5xs/Lr7whx/GncR2qNpD
ceeAOan73B97P2A8HFP59ei+j4yZQc06zNyjCw4nSAld9c9l3Pyk4MGwNJLMkAF/z4i/JTMjLrdp
WQNolyH4ePhsS0IBTHdldHsbyIEUBop6pibTUfgosFl9oTNizu5FNd7sGt153KF+3gHPcp5I6qma
U5BX/Z/E6hAI9tNbKSKTujxQLVE5gSa6s/I8tj2JPjVCi7yLESBwj4CaiYgetwYtkhdBzpgHnK/f
1WWjJsY4Icezy3DuZAY4809FpL2o0GSx1iRpUpUt3QGoBF3hwS2VuEsA2cgwelMBKeBQTVqefW5B
3N+YJxC0M6UzzgJS0u3DykY/HTXyfTaA8GmMWfzxqXPNaJIWPycDOON6mksagoeSSjzpD0Zyilag
HN5zSVU3SujOfrEijmPviSvJzucvJfOOahLkqfwhJOHASltWggdt7ITvgtZ0qcDcM8MTp5Yq0PY4
lTjnZHT7gDGXLJnKY4HEsuAAYB/YDiE+6x1YJK4jrdq4uK5SiMdfFSXRWsOFUu5B/+n+8Gh6ep+w
E8IuD7EVcego3FcH08AdhlArbn/H9CcMl7j65gZ16o3BwxIj/FZUDjz5UVPAJkjU6sOb4NiOCly1
ffB8tjLggYzSmYqCGhwp8bF2+jGOh4jUYynY4eVVvMEmLbjEba5oPT/oMI/9vd1nQKOrOk2WqoFz
vbKmq3OWW3lTgwWR0JjuhN3n2ffsATK9RlpJKgwDV3t6zT16FdtiKw2XkG4+gYvNu1g6JxRau4+8
PdN/2nQcYumcFW5lhR84lvIkoDwV9hXa65tk12la/+hh7Hr/Ztx+i8zJrg9LwKwEbqRSqm03POZm
nAK5sGCd5xscuar66Ucz3EpzPNQ2rIUSkqi4ZmrrG9CTgzCgwsGNxhLL5dU3Apg5ow5HOvOqD/6y
uP5k/M+Y8C0L8jeyRlAIkgF7m8hStLPxsf4u2bUOaTTIjE3WfTLs/alRTSOIVcjTHYykvnPluuLn
/Ha9kUoLLDuv5faPKWm+n/t2ZBPEwmVXhQX/I/wXDM3fuqj6vcCn3cCb+KS7c8MNYMZb4+mkzaS9
0XMCUrJNN9fTYH5UBAXIdJeUQG1hC8lGvVXpw6NCESpxgIUv/+3dumzoX52DJ/PSPEwPjVkyrMYB
QiT+LjqzOxuVLqYhPTCKjp8Kr1jdku0oJAQWReLpFk+JXJBcDEjONh5fsBFUQf59yKgJh2Vys6d9
2t1FFohtiJzPeFLsyk0rpMFTFOEQI7aaC+l3wY+hRn8lhkILWew7f5zfiP7/7YcyYYiQ5uHKGf1p
p1xzHrLsvdV4B3R0xPa6Dlk8gDlBtdlRPibH2dlJND0KAfSVCLrutWysV2mHBRRslh4oyjRUwFRS
dXFz+g9pV1TH/9TPJeYmws1fhY9Mka7Dg/zFkQRTmAO5nUnoOAhVNdpi5O0qLAiyR1bbrRZst1ns
r/neULy4AC6ISQCYr3482rFsMXdOisNlYiICxjOpGEgfODOH+gjG9i7YjmLu0EAbpIIZmzPd73Xn
TJFphN63sNta3lXJvDSrYPbqy1YJUR9WbEPt1tgICaDQMreGoLClooWWRSlijIfSfM78sEtbEV8g
/mIXT4oXkTvkEDs3USKKCVClh2V8Xc1Ea/tENOvkfpcYjBOHuuTRrJ+vra7mN0wtdZPOGeQr27/M
f0LqlwKA+nbgHar4/+vQITlFDzhK1YIe8peU1tRgeLeSRD4sOqeaFmyTV4N5LpvV7ioA5Y1JjvLx
ySrl90YWqiJC4O6o3pnzq2C7pfSCLhP7JnmRZScHyBNvRBOKxBWY74zTRI530Dmk2p5Ojhx9iuDI
L40Tm0OaM4GfPqdcqCZ0kmVhxSjuGyzcYS/jgnkog8MX21EcO/HVzsNiOo7MYGzQJKYkXR6P7fvE
FqVd4cAXKMAVUmwz8el2oz04LMNxlOEbS3AYWUSHW081jO8C1Od1az53kTGhTul6pal1ErEKzucL
1M82Kq/oDQbIG+o3cvuR+8z9FjhYFveqmfIjl9vr8cJdrWBcVGUMWzdRcCX8b3tenKKz2BJz6srM
DoyCQp64+kkgY9qStZjK7rOvqdr56Z4NfMjh4ShCNL+z0ab1GIIYRapFD408VO7WOSA+Qg0kmaLd
K0viRDbl0BeDmgfVEu6p+f5wqsH8ThDsE1QkbAUF+OMicFT6r3O7neuQnZ2yeQYju6ZKww2jHcYD
RImcyrEcKBi6lLyf+XsmkjGsHi3OicivYxd7CerWghH9YS8U3ugFnjtck63vFPKWKzNCrFuRVFqg
sXyzPSANwYQkzC0leetMj1SZTJxx3ggnpA/jXjVx2v2reaj6H9beiwiCrcoIdWlmlaHTSAu9p6/F
pHANlHVi17HDUSp9Azgz99S6L5U9rlCjQTBx4VEWjJhNAOvBxrRzi7Jp6m55DvFnm6zOkfFHvhYf
Em6Y+xGGIYkcP9pwSDnt//LxGOkp4kRDeU2r6y7X5/xdle/modJddicwTUZ+n1Pr6xVf74S0ZYRW
EWHyQZQY3RuRpcGcWjc1+8P2va+WNHIqh9tuq1vPfSQQoeNetz+Z+fnIGS01tIMKKfU0ded+Ku8V
DqWlifBKbJG+F95eRAi5sc5cgpwegGMo/QN8Y5KoCCPXJG65ck/PQNFsflQc1nIjaQsQ6pB1xXc2
ekDLMYJi+kO3Cez3jbqUs8ps8xdaVKc4WYaqi0v8XUl1fmY5Hj66QWfAHFQ44rt8aWw3XJZaHoch
tsnUhZ2ikIS3kVfTFz5E/vy5nOmzUvXLDkDq/FXhgSRRssPRpPN1OYKvAkJxBMlI0s0UFtKNU+e+
+H1wdIy8DAJE6FZJqLfElu/HQD4UVsSG/L/HNdV1aKgm2jq2+whGGwfv6VYPp+a0q5xAerCrTTqO
n+XVKB7ClqfWQLK1wJGlQRPllTDBPDI8kzEqQy/ssN2wv32/PjT1o7srnv8HkH/IIxn7y9vkdamw
QeJPS03rZ20HlqeXuWGmyQ2YrCBayb0AMah9h0YP9yo6134fct2BLHpg/lZTGRJ4T0MxDIG6/9IE
QschYnOFhnERDuorsZLF5ru7xeW+gOigmEoPgy3tswVOSdUkO+tVWtF/5o7t+tudNaXcbMH/r0/q
JQ3rBYxGsf1dsLEt688Rnz2LM8+copJZxpFJO+6nFG996KQhDfuPhNw5eh3so8rMId5kyookJYbv
31MtRwp0yKL5D+Q1zCzMadXatE9eT5u5Ot53dmVCPI0zXIk1dHq1R52InYBIkrFzdZW5mhYVmpsI
So9PL+SEjQxEZhhJC487VP97xiVyFdJ/V0hi5ME8XelbeL/43Tm2uFiWSlApkidxM36sSP//XPkN
3U1koL+7tNbkArwlXXApcjXjddnudV+zvCPCjqrJMMHUP3k5XKIs2LS8fokIqLS5AU0xhGmY/pay
EPA1KUJNFFVjtxdnCCHPayNCoWuSJlxhe5AnJGQgMRsSHjVFKkFz51lajJvI/86IhnHaEQu+W9CO
Rfvt1Hsol2YgG3P/BJdNkez2iSxk3ef+qacH6r7I4YNAiaolKNBbWVwBOyP02Os32PtaByaegl20
IyI0t4e97gg8SsPwTwouuIeuGT19qGMvfn2p1GbwUq45o/4GKk36vCRoWFUR1nVK74aEr0Y37TCm
Igmodix5F7OX/tGLEiqNX6TZHyBdv/xtPEkR0OhNXaSB2m/aXz5oGZTlqylrm6/62toHno6VS3f5
h8p8eu972K3Zg0NMxtSbGuffZS4XwzrJXST/28bpeX7NJqsydlXUau63QnwtNkcUaTqZzokKToJi
5ByOuW2RyIoMtxjplprWxDX2x20k2dLp+b8XEi04dN/L93iCI+gBP80eJF5X/ff1hrdG1t0dE27L
K906V7zvrmdRxz7GvW1W5w1bQihJApCycr0QjH37mfEA7W2XN9n8yWK6/YrjLR5kLoVL3cf0V90B
uKIh1FGPvY58YgyA75fffNx969akSzjf60AN4kewyBiaMHESrrC33Hi2aY8EV0Gp2v7Ri5n52XTy
krjtBChWyj/dVLjpffNyr35CzEgWlMmLAtZ2DYGdJoRmNb0y+3KLNozfrr1cbumbO63zHW7Pfvos
SHJeMj3pwd9VHQFwcZIHvGenZFJkj6XKmjXJJuA2PWjhg6XUB4Wq4rPtKkZMOO0DBbCctgHAjGeK
FflmVtyPXYcTqI8SfoLOsIsvq0Uln/n3aiC9Wl4RkuWvFQQQEkSpCqRF1wg5F08ok8YGP1fsmjQD
tr8IzDJCUc568p4pZ3oKiUaYTyUD/ExJMq3WLFKbj87yH3auHS0YFa7JlneiYGuR9U4a3JcRRYNN
3nlGV4TGHu7jQH/L1Q9n20SF284jVI/Msmyd3xjHWnHfBX4PdjMZ23uceDSOixG5jUnr6tOKYmcE
6mvFUCgbApc7B5XTFLc9bx/uAKtusSTHTI+qsMjo1/hDKNR0GcGYxgZp3QOy7IVEy/TFuU+4D/N/
Jb0P6EjzZUWoDhJ2Y5k0khbh6ULz9Nxz72KlLAePOCYfesDuKmNkAfbuoh3QPa+7R1e7Hz8eA+7y
C0OLyZfErIfA+v9Dc7f/2Z9Ij6DpJWFmQwEGqrXBh9VtiJSGszK3ctPpTpxOUxC4kycxpfxQ0DcM
0U94YtFu/wNzfYYhatLLymhG7i43qET+sgQ218O5oUqzC90+idlaEd0GUSbY4SCfTz6OCZ9/lSj3
0AtjsFQl75BaemmqtMPGTk0XvxISAJEb8PpGSZZHnMhnp5/ZGCuNZCre7vzMrcTy9Qq97dQnFTRV
jDbF6ccd8rXBBJq5d6Fp5k62Cmo0VR7TPNRqsLPgI7QiTDIpw+q6+7/qGi7rc5nhP9OXescIP0I/
3ggc/SIAhaq7gaUor5raLqG+8mgb/UobOKkjB08VRm9dJsfStq6BVJKH3mueNcG+R79bBOsvFZRG
NC5JR2XvWvTPSWpW9zzxC4Pu/HNgGjI2nkKd9rfGGVk1yAkFm/38u6vHn2slYcaC+HZa3XhDK+k7
lolw/sUVYnUSzGhH9VfEgV2qUsaw8/mPag9te5cCXLM9ejsnfXGYW0PCOcKnS53kPFoNq4eIKJAI
52IFf71U56SrQ5Qyft/WhRoXEIgRo6XUOawaO2HDLJh6phKp8/OSBnRB0XTBRB7AXYYLXb0vo3qX
O+NRAX8Lgequ6oGRiXvCC/Lf4Zo6pfVsjSot75kmr5G8vPLqBw8EYvILE8TEX20iJcZkmi0IP1IQ
LIjZyJm92FtkSTuNgCdr4H7aaNl/cndB6/IRyeHkjxNnmSTkgR9bbyV/rgzPpEWb05JLrvuAPiRK
lEGWKvhlXXy1WkgbAWbj5vv7ikCIhyLM88CT0KRY+KwHL/RaLOhc8WaTq0Q30NWo3mJRle15Z0IG
K+u5504SrX42a3o0jdHHFQrrwQB9etWTGeM1kihjyHvFKhSbf03uEa/nIxwJpBe7tsqCEhCYlgUq
xv4hEpsCHrbmZwFngCCNg0TIzIx/ufaKV2bffn7bWyv04y3AvhkCSmd9gfyIYfQaOcDIJsEjIUY0
qZNTcCADN7oli8nWAGtYYKd2DvCEQzsxqny8n/9jus628xmct6LZITVy5tcpzQwELg22MMODi5pu
zecitc7aKGL6HtpDKrsdYemQ81HjrWmUl1rfhL96qWRati/fnL7WbJnFuxDrXEdwpZm3/B/bJqRQ
HMy4a+ABwdzxuRBS5/7jtujsYzsI6A03ohuLmOK7gluyEMt1qOPQebNKY2QoLmwqsgyN9CdN7ppr
6pzQ55zunTL0pZGqzr9HyUt0OJasB4csLVlGbZTj3gAxy6hI8dUMSns4sBcj3TkXWLlYzA6wQ+Gv
hwSSdtfa/9w5t7DEwS3JdNOnetEjNRhC6cuzymh2W5ZpPCCiA3ztvWMfKAP8IxjENBDD6oFEqjVI
DNq3X7DycxFMl+JRtnZdS0F6HafskNIJzsmXunVcK2aYvz7v0gvX8m4NgxS9pdx0CuE6Hnb24q0a
9rr5ffi79cAFe4Cl+/HyNzSF5n+DAxPCk0nuxlrw9MttkFp4LIatNEUGy7yTushwYmFy3tEOdwxm
xbwOFUI3rlHg8oQIJA993JxM6caV53VkJcbFYwVdsje2tbdg/UkOIvsdKSe5HSxu+tUjNW4Nejfu
gsLkz1YjZfz8yBz0OifImrRY7lQkjCf2qnnwf8N6X12e+ILSQMOyD65ojxg3vGr6G2+fUU2GLe9u
G0Gh1i+r0CK5VFjzs6mJcp3gPRVQIBjYFOz/AzE0dMZNrCGspmZ25Mxih4QEtZT6zxhjpwqU0FRh
ls4C7UOv96JHEIfZ9czjNfdtw5JMRYkNIPHWBxq5Xj2kbn6m722Jz2LwKAOMcX+HFxwZ8CMX16Zb
faYo19JM+diJjC0/jeoN3qT52+bb/TF58DIVSZQHlVEdVDb6mZfEjkaETQ6H9jgqdhdfMjmBgT1O
vifWsDe+e+STZ61huB08ArDUkrYADhtS8vtzw3QMNTgYVhe+fwBNec5ZB/6G68oIkdtQzPVbTD/W
CnH1vHAOch6mDIiYIMg25imw0n01zidwEvYnjZufnT0lJVec5ss6qwLPP91Ff03eXC58LUd/RlXK
M3FJw3ygV35DMQrUR8UiegZKkRH3CjhsQM5S9AKO42bI2ZsXPukpqeXKetMIuyRP2OCX5nHymjX5
FDHZDgGHX9au+J9NH5TpXUQwG8VYrh+VyBfbs7hu+4GadoDvEL2KVklC35t4SHUQObV562yu1Izy
nF1IXRLbCkcjZhysGBcZraB0POM+kIbBmU5EG+iO8VVtBL+qAtwOADE1UmSkR9ntpaK93s7VP4Aa
aBBj7dOMzfw7lbtkp23YzZjEM33CoKRSLF/A2ZYPD5cmSPnKdbxwMDqWkAnj2YBnSqG1hn/OGJQT
WW5F4SV5f+fYN0v/iRu789rrCblSGIW+AnTU6edFXXg9c+TYQtnqYADiYgDOeg+N4/0NAzCkNJZd
Dz06CLkGcLrqEzEghDmWtiIviuT4dv5KyKD0Cv6JGoRyLpWx0Y1twWU0J+1W87bze099X3xgDYmd
4DI8JtKwsh08FM6InA28xcXaE1MXe9NZfnSzpENJEGQrW5UueelqqgG6MlNW9M1QwGjW2wyaLLn0
w/k2Cov5Cu06wRg6K3pwKxBOZxTdjJqjmcvSX9y5KIojMaTurrRFjtA6n9O+m4rtxXYDc5Js8BAU
USdpHHcHN+DceOWQ0DNVd161o+APxpNlQXh03ffS/64KLyhWENIs3ghG4PZ9AsXBzSJZNK/KqnGq
dhkYR0+bqyRYeqSirWQ43rSqxYQBC+0U4FP8xRSbVKVSJMTQ3px3nnTEQWvBjAvqjGLifLWgkWh1
2SZdBocfs9NUkWgwJlqdQXDPAqYZQoCFMsywfJq52lCwy+lUduNc0A42uQiU7z4G9k6F64XTS2nD
yxV0R6/E4676/J5EMmDcIWHCIJR1LSXSC5/2d3xvaIqr5lBcxHpID9bO4wbT+suZCXjAcY9ZVq6c
Safz9j1/i3roNR3VLd02JfvBsosk8KfaqyCVYES3yqY41k0y7YYQholemA4ZnZkH4bEvrls8O4uJ
GqUaM6o7JDduDFbmFCw/R86aferEtQ0K6Gzm4rQELgAAIatpKUzxo8J4HJAsa24H1cLrlt3wNKL3
nR0bvnlEnT7W0aootXETtWmiHQUhe/BzGrfBWBZkHVhNaXNQxKjS0h05btYp55b2SAC7f8tlklUu
AVuZ0AF5FQkrkkSzU7gZ7rF3hkU8efOVj6Sbs4fdaR07UcYQW16LI/1/Js8IN7v+f4M02AgFKld5
JRtSSczps3ftpm1j+4G6iKxAPM6EqBXjhIErF8YsgOsJwCaeU6UkKQXCoRF5EZv/A1beDX0v0gpg
PmK915pZV+EknAPbx6lThUGqaDHDalDbQW14O/rLrtfuyjT5founxBxVFppKAadOz1RpNajccELz
fe9eEN/n0sAiQt68hPndfpS2AYyFs3Ti3uncVEstBT/2ONJDg8CVOOhwI3DOA3AKU3Iw/7jUQ8+Z
7vyF9la03zW7J9+vlfxmkFk2IQo/+B2KbszadvBmTEZhR/JvfHkC2GL+tBidAoL1+ZpSwk8+Edq0
nV4+bQ0pnl1YUsiHDmrsjHSvDz4gROHUjYqgySdxd4lDuf4bV6gs3qhvJTFrFFd4R2Uk1HfJJsVd
qW/N03TlNkGe5iYnK2cCAwm3rnc/6w+p2Jaag+HRm9qvymmIhUkDPuevnn8py+cuXZxf82y7wgQZ
QC9GMmVGi5cXfjzd70hb/P4TIDGfVhPVcBK0Wfd6cOP8DXuMQMAHKQWOstHi+2ePYoOYGArsu/Of
pd8IJ7gjmW/7Evs6jbEg6/LZ//lKM/ZBDMznGTcR+VPviY9Dch3o51ayP4XW2dmgrCNvyeZQfctX
JbWBzBHsVV4wURaLbGLz4UuL3jrVkuS4qF6NEolfzSjbL7kyNrkJ9N3ad5VKr/B4zz60BnN6KqEf
QOdHQBLZaKJ1qsBovO6BTBY0pd1YM/Crg98Bx7MoN9JW+wwF7Q7DJ4lD8k+uTGK6z9xmmuNfG4zu
nsKc132jTUfaoa68MzlA9s68bLwGnklPAtcLZHVpZ8ZATxhaxKvFsRotyMsia0IrFwC7+199os2K
ph5xNKrpnrQuAiEbOhgxIxoBp7BQ+LRD3sioOrJWUpUWgv15JaB/9l0IflOct0pvXjoPrgypGzrm
iGGnCLAsU+QETVGGgfajgGrTiTQXcnv3HHuKi5oNGukGX4BREqmHrr36GxY58/ODQzxR09qbsUVe
YsdBqNp+ByZC+hq3176vOgv8A97I/ujEl0aZ4rpgWSAgAupWi+eeQ1OzrRNNUilgC5g45hMlbIfc
AvJY9axVVysvOFroRMwpVa8SZaBr3GggUqLCMB0ngOuZxy1jeeRBJAbhyX6mjckMhsAD2bKo1L5V
0SbfU3gIPlTVS/uM6XU2mAQK6vw7augBZiEKYZ/0VySp+1DM+tkD7N5D82lTtIJ7oF5Ci27FNyUO
GdP84aAu5clfyrgJvbt7bJIo8z67OQWVZJwKGTxpO8r98qekiX1NjEVXO6zsWdC0yz5YGjJIP4JT
XY82m8PmI8Xhxmn4g2KO2LAn6oEBbcqdujRSiEhK1ZeKZ7HwVkgL00fUBaMl/ZW+z/vOPDNpWC8g
UoyiHVagt/3mg2qDQ9/qGg8PUmmFGJGHHsF/T5PBya89bNkbcSjOqZzsevEZL5+yg7dvf4ho/StQ
o9VwXABRjvRcnTdiGEDb8nc9QvPbzELZ5v6eWptl5b8Hug3zvfY+12UiIE4GJ1KEB1Syc76LlF3+
hfyQd+qhj6CgXgdvbjXWlpmjaBmABjJgyZuWGLS6VCYgkBQM30IV4xtTckNYmuulb9VDiejeH6Ot
kaZX+PXoMZlKyYH5V+VG/RjP98b+IK3YZA0bUu+bs7PUy4dM0KPeOptigBgz2oraACOS2E9gWCUp
mjtVBKB9izvfpyC503SQ56TnReIHS3rMAz4T6m2gPGetrvAW3mTD5sUvqwB4fPLvRAlgwtQu5JCR
aZqvDwOdiIizBtSyY8xnaL9kHLMwkFfWxhgr3bAJlQg7e9Qb/d+5vd9u7DD0QqTDbpl/S/hCVgXu
J5I0gu54nl1DdNYfy7Gv+09s/QWHUMifJaQgMwC7yxS4+hf8EcVDb69wtUsIU20/RMkbZw61rQDz
JfVbh5btHFE2EijPqsE/A3qJeoqm7jYtxrupYPFZCbkg0ogaTPCzmZgL9+7uKW36VhevQKRel9C0
AE8jQBjQ2K5vLjzN3/6Adunli1qN1qdNQOwGM6/BFZOO0scmML+9CRkUZaxxGe6eB7iKypQHUtnZ
iE/ogXA8Jrhrx4SIYnNSJVkxp7z7B66AuzW/5MKMs+AKLad4+E/T1OyzLUZokbbCXkWVmF8qkF/m
qz+/LtgexkhdSbyzaKec4SY1gCITklvT4HuWHoxwIh1Kaa4Kldv7Dcc4Tz1UY6Y0UAtSvxNur3/w
rkmsLEYm3/f+iUJnC/+q2om30P/qSmKuBJufpzaDBTlcM86LYHzLBiHUF51M8a832RPmNpvfxp4y
wL1GioxqHhjhvtdlnNULF3DuadjouonNAZNHhBjhlIH/bMJU6akwtQTeuN+sBOZ3x5v3QneWIZ67
khRQ3sQypPcHZXomggRHfv3k+dkjiX18UqA1sn/R/xtE/fIxn7eNW62mkq0FTcqOVraGFkMjGJLs
wRvhoel6d5x7fWubAJoY7h751gDPuQV3uABPR0/x9mrTYewojGT0NU4VG8KYsYz2g69CkasOX9Hg
/JzfSkHReD5XPJhjIIUPU4jaytfuH8UVNcN9WQk4ev9PjJfNEljRMbwhWa41QSVOwnh4/IbXpMQm
W9iSn/f43Nb10iVBARs22uQ6bLM3kH4+gx0h5XGS32uCSEvTdWFry/UzRrUzooI3o0aJk9iAb5uy
b4HtBDOyTxsCD6wfr+sYw0I6pNZGAZ5R7J3w2WbND/7kOY0/y45M35lBymFUmLQ1Fe8Ggf3D1+IA
4TT0rzgY2OAJ0Ld2eNedxAMRUWkiUOTmzM7/0JktqwoFDYjIHRu6ZaHZfzNAWLHYFA//R5OQPeY8
l+5Aa5W+4D3kjKttVZt92s8BEscuJNqAi1PGWK0wjdHlTMikX2S4HdlHw6yB9uL0c3/pWmm53SAB
x4Os8/tQFOxg610tWQuwPZe6wPVfvSdn8RtoYMlKR/btpftrKtfr3pyIICwrfQScj8MA6F1+7Unp
pVluGLrZ0hnTH+GVqoZEAcDosPZu3/MuQLmrgJeeQ5Zxn7SlBgZ/4vfr18jFREc6enZlEp3pp7Th
gcjJOhMH3J5zqBq0iD2X65m/5EWCeRvtJ4c1kJ9R2Yyj95kZQ2k3iIH9xwIlybY7Pw+k1ac+L/FW
d2j0JzxYSCw25xxelNcYm5IgLE5suFEJtBCCe3e1m0s+8RoCw/L+cYS5fmUDflXJM01wuPwSUspx
FF5OkNbaJ9EoZmkq++wFtbmo2Sc9uxzUh06xt15R4vHsJjpcWi0g++rWsmBaFPcYWk5MWmWEhtqF
tz8el++1GaBzwDwUhoxqh4iMwtEsilS6qML6mIxpVSQVPy6wSzVFmFsnJppyYck6ulYta5Q627P0
9g+nxoR1lr5D+nKyjsTpPk23a3+MRoNEMeP23aIspd5YIYY4VBaI9gKECxsxKsujAn2Q0fuV9bJy
GwY4GYnzjzzbKa5S6QvzX8v1/Rk3TUZcLfvuTLcgB9PIJ5+8/4L3pJ36ZqyL0kmVM019nsKg97C2
67o6Qij8pv6aQIXxKTdfZJ5SiNTyB2ggBObb02rRZc8zirsaUJvEqk4+VwWQ+pZy0ZaXWQp3/QAC
mn5cGjLYaHenj8Mo82h/d9FxXQDxitpkoST6JFCkMjge4enCbQYhUD2OkpitMSSPmE9tE7V3CiZh
MpjSV1dUqezqgNtV9lVovg5MlzD+mvTRXSjxt6pwodWYuyHL/iKU/GNaTHv2c6zL0THPjQVqtZYO
n5mxTpp2OCLgs2MggxytVfhBUgJvcIyTa+eNvzkbPtpOIu+K9HFOXeOHHg4kNiaZgF5Yb0kAm+ay
OfSGTxMcMQ2/qPvZoFdLCKe1cSI8l+8mwUzXS9qgxk4mnGGz5u+sJp9ZMMFKlfsL40EN0f7MJZtU
EMBy1XujCm9JnzX7rR3yYrlK5BEMUC+65xsq7pq1+wVYCiXZm/COjm8e8qlx/UreptESxIsWXXNn
0hqn9tSD9xhnPLJSWaABhOQ38Zz0tQiGcRUhgaFEKRY1PzGZUWvPNDAWPlq6xBcdAeK0EauwgGNq
gejbZLjLxI+7dpl7Qruj1cwjtM1qkYbWE2svueBbNVDKiatQ3u/eq4oTUmcTBExxq0OaldxJj56j
qzhfMXmoJSqdQn6XvvRSj3XcvpRKTN5VlMabDGgxlt1Dosw8z/QrljnuYgtc1+ijwbCk7okcPKuV
q2uPLA98hy63aNOiQiKC6UDvha3ry/Dl3++8/PFt7smZtj+rmfx9U0bJd2sBB/UkDFZK8Jp4JGKD
6O2p9c9bDYswqA34gg/mmQyPsP9epouZhSkpBdvvZbm77fDSVQeDVVa2oVOhdYeJXIQRTSIaYBPe
27h9Pv0kfGxtiQGe2q/Sm/Um5ja+KUn4EpveVXfVgH9Dfg2LCJ4Y8gAgXqgjke7u1gzDMPKtEsXB
h/phbtatXYwwMqQ4veYf9aGfCLbXNgZbpr2e4FIgVFnFs2PsovP/8eDaIuJPG08ul8buSwsZ8bV1
X3WrECErQUcbCcOX44OnSAz/7p4Y1fGhfBqbw5ZZvoPtLSmFpAN9Wyy4cRS3koQA72SX85zGWdW7
Hf/X0HeA9LOrVNoURtn+j8yNErTHJvTObE5gILY9hCDB2CQ42+bMfhvK7gZEWpPHpLMGshntaLI+
YIxzyggfifooptUoxVECzcaxEhsANTesuqPYidrr+Ej8k1QbNPAv3ffk5Jlodsme080UN+HiIo6i
vmanHI86MrXKfd5opSOCRbOKlTZJkXSJjMYU2T8a80B39kz7uvCOH0ZeA4q5Mv2HBMJm9jx9VsbS
IztN8DZGzRjJWOz0t+FrrKsgCNd9LmjEm0AMeElcfU/W+sGa4PSKBjDxYx4uJcWhve8O7xXH4I4/
O7iasl1n+la1IyTGfejOXzwasvfKknDGPmE4/0J/mrJdj46nbLOmHCD6l+9AHdc/lq4CELCZ5EZJ
ec1CU8zYtS5SbIXUGrpI28/Dsk/BfsSDGuj2nNJmUXB8cu2nUBCsdppukuk6DCFrxcDuUiFnA/6W
2s+3dPfShE5O+kLYQwZzvI7jvQf8f/YsRo9l5S8uEERRnXdg126Ji9JpcUwzUOQOmkYcBxpX8Z/t
qqrcbKTa15NHf36kFddui+XjrO04Co1jtd4eMfCvu1EUqcTJtyM1L1I5Z/kRUHS+9I4K6sL/74+P
Somkk+8uuv+sZ2TBhiOAe+Ypjk3gsFiQ7bUrQafZSSscbUHK0uf4eN/ZovkGkr5vf7BTQLobsKKA
LzgvvFJ6j7mG73tls2g62Nexp4TgmdCoOZ8WZqLkz3ztLgd+EXbx+Ki6dwocorAaXt5PySY35jk3
tmStavl3jB2I9WQi270rDXUHfuFTaoHuvzB9qgHK/RCRbY5wvSbfziypQt4lMNfLPYBYpCnQM8wE
TB2h5tA4hFu5rHJwf4Rue8uZgTYvNWCNiWOY1ZClEw/eHA7qPkeJGi9Cm0ic0QF6XCkPpzPRY1Lt
9j8dIoJjRb3u0wy266wlr7J36AomC6o/5LOa9djuXTSsohXOhJ5yxlZrT6XJo5yXy41W5aPGOZ6a
wMyyA/ivwyU3siJbOaaQo07P/MkT9c+WgSrbm+ridm+sdeWjEFRKwOTED0wpw3ckhcmEPe6Bty1S
5yGcMGE41RmYLQJce6LVm9Oduf+1ZfIBh6KE05CCAOo6n8o+LJxeVdmaNeGOGz0nWp9nIA9fKtsS
mewttjGEy7X77R7iybTZfgzX2YZeH65PyHIEVHoRU8kI8dWIBXoBt4SpnZjfHagoziVTTzf40UqS
npgo6ofNH9eiC5HuZb+Dypo/nF21fsJHebJIW2ULpHN6oeC8qwt26XLk0agBdhMF8nEQHq9+mWMl
xpup1zq5dUOVCBd1suaBNbX7oYtpqKQ2TObvLf4fzti+3esKg6jVjlZQWeBcjZcklH8crlHHNQEC
FkzwYYtbIhTGiTKcF2d9mlQYkv/3MH1JeAOvw67zj34L66Q75YakLPQr8pudZqcCEZLwFC2m21zM
F/6hJ+E7c52c6EwRcNMM7mgiZPVy5Nv+vjn1loU3UeDRkMIg1a+q9t5+1PEiArkJqTXiYuTSrBId
fC/sStCCZ6FOkH4/Dr8RkoQOeKs+xPwP5fjnN33HMoupZj5vJPR9aOiba3xaj0TEg/TmiJzlKHQL
GG46joCkYjoKlxo0eJV4FhHJd3HxM5mK9/lfNS2jJHsv1ae5C2Oa3Ma1gZFwOWz1U/932fZcyqzw
dPQVmw1YsSsX8Kcve3xQt+Nr4ZruIiDDYAAs/pVtut4aJVeTZjfShBu8OJO+Kk0EJ7XiQFo0Lmdf
yYIXJhtPsRXwNKUoSg6U0He6PJE5wIRE72w7NY/7yIeEbD04UZqmoyEicd3n3xof0p1OuVULikai
+t+UvJ+3aj6Vibam01gTICBWP3XrXwkkFx2PcjPIljQAojrYfpGi6gHaYops/ZTeZtiuMk3Ljdxu
r8cnQpsapv6zbCf2MQTjXMUVaLS2bWhKrHKFJSKRBJjLn7lFmyvYhVB/JLjQyt+lp2j7KSwZy4gy
qi9/bc4tXpHLzZ+eFY/7ZVjI0YkidNns5Y4aKp/g952TYW5BtQlMW7hb5jINmCMo/UjsuC8FHED2
sPMW1f0WWxSZAG4+IIstJgncY0+2So/jsgYtoqOtqAuIVo/iiCDU5pYBhA8wioiH2nOwZn+ETUSL
rUJnHAzQyC1ByNV7iMv9PuAm9gJ7SxxB5ZGaqvnlr62MfF7jjXKmpdzohoOXAO3BzswX8fftqQnd
GfwDIsI3nlwociURUjmXur/qhrWLlPuikC3Ht6Kb/R319nseDfxztn/ncbAzkomsg73n6TIFslAG
bblhuEiDM9jRsRN4LsTZ/n6sN+BLujk4e6cieZXPkahWjOhQ6HMhwPu9IfDruWQddxRRs+yn/efj
TiCv9AOdyZ1VltMwQHuNbN53L8PGfvhHtGS3NwAuSE4NGsfY6NiwZ3LnNNqe8moYx0hNCgrqk44S
xRCNhxgaUrPwaUWR0bXSYD5fGkF93KV9Rgy6dzrd3bCJUkh1wGVak42SI2YEGFIp8XBvjhjrCycj
QtsYT7zKRP3jwuQ9YW7Hd02bDNVP28BL46yWkYTk6WALzjwXsrfrIGYiE3FBr9BVzE62/lAKy0jV
sSClWFoltYm85k6H/6OOfapGQcKACUnOrAPAIYsemBbF4H4x9hmifXN4/Q9FFkXfilLOLUpxIhkY
ripZYaNELF/RPjQXv8sTxXCX8n7qmhST4LcyA02vGn38ckYoU+KfdpzRfKemH9hqTOsxe5aX2ZR5
SnQpsjfcbDgaqaXxekeck4C9EJ+jpOqiZoGrOqstCOZDqHbF0LDKtQKk4Wn7nPrCNghw8zr+4Sd2
BJl5gznU8GiPCtOzzPqssbjXTEkvO/9QACt+ouGcJ7rjrA4FrsiXTbiGxx/eht5M/joLNoFr6ob5
PHl89zVIOFDmTzCyILxXdhxOKGIcETCtET/pzehufXA/n2tu9A6An4KwRBpCMem4lRzXNm4Y6X1n
g445lGnqPV9g6CUxplkC9EmYTItRVoL9LZubxz3ByBXsI3BMbWc9njNSSfZEEMNT8StRVyZ7eV4B
aFWMSHXrthrG9nS7sEq5Qth2viI4vLJGQBY8Df/0h52FYztJh4BgCLhD1v4jVnBpp0riVpmwl5OE
oxmnTJaljffjJAbTW4CAdMJhKlf583dYWeKlTgEWcOqEI9Mk16IAlx4b9r2aDk1A2H/NovLcBG/C
n+Rc3BdrjR2mA/2y2TvlEYktOZQmA0oqF9rPQl6Na0ihxwC4rVsul40RaQ0psiUITcA4is+0q/nx
90oVI7LvbNhKvzQ2hD4HCGxSWbJCu83IAJi+WXg4TrM1barPTQ4vzca8BY0QsK0odRYFVWkznOAt
wKHcmDgDhbpeCRlnydBzLKlnrxrGL6OKQ778J6hjHwEtO5QhOv+cXY7FWagA7bYcBK0MAvgQKvVT
I9Ih1ySKGtGYdWAhQBYAdF7MFzx+jP4+FQ4QWqORlBNGdAHbrN9wL0dkoyfzLrFOxTd5SlDJNEx+
vIMVFlqX0kr5ADig5pB9pBMKBbx/IpiwHIIsnrLtgoa2E0N6lvZL4EtYYpDn+zu3zB74jCsHfieS
QXd2J7pPp56yhej6jJbuUECUSygT9LIM0EMH0aNbeoUnsu7pO7RPH5o/XirxSBxHpx4mc+FHdB0u
6yw90waz+mqxtnod3s2n3o1uIayvOyjQXcNaqLT4Ay2QLOvQP+i/oA/LvHQOmV761zqMLd/AKXyJ
COHs3glaPOICadJDb5D1ITPbxxzwgEwODjmhU/7x5aEmnWGJ0k3o6VFoCQfJ3RZN0LXSegEXqf/e
w6m5krv2izhh/OkjXwRocOF5GG2A2beFFib8WsobzmXUNsaLWTTMKKMMVRizktg0OxCGiTIFpHYk
ODa6OUFQKxsCKnkP0j4EDXniqL5ICTyXD6tCZ/uTAVBA/i9fvdIe2oTgF+5MMVaHZze37oOCHTPF
tknKSNSmYeuhUUgJEJWMCeDeg4ljcnpcXO5Uk2tO8c+wmpa+Jiffg2B98Ow+HpSzOymFaJK+RNhh
UXmouU8z4WRiXcduEQDT9dV+labIn29TdsfdaAqMowpE4ZOCbBHIQfPUg6efcAU/TjGfYu8m//Sk
XcXgeVRd8FqRmZUEnlClOxKYSsIlc7FJcxSSYmELcZypJnVbUCrXg/MuJwKQmckOuGfSULX18N7+
S5E7RnWHKFIShR+H2GAr1TSNye2omFOBlonSRQdmX/S3QnmSooAsRMFGeZTOjnMjjJckzXnW+EYM
RqVCorEaGNxy8HOVVh9c4I8yEvVN0K/BY+O5cBiav9g0h3DXETXAiJPl0jkTKtg6CecI7zNoF7eK
+R7gBnM2r0NvVRUZDABxddFzHdFl8HqlBUNACPDiXjGMXlgcrdtc5hsvAUhciC25Ar5YqcieGzAM
Qx8eVI0tQ412xSSGPuHvWIamjlJAatHBED1DfTB1A8NEJTSGhka/iPSj0L+aY6rDQT8eEuHsHH5J
S6fx1hJLEM0Bz6TRq8/vcbUQQh4AcT/pb6veoMFGpHOZwpw39z+Sq/+7pBdmaB+5Dnc0/vQlY6yt
VLAVSfVWeSpYDMzI2FtL1Y9PVTsMyJHy6w5rBdAl+g/VQb7gXzROB71rgoCicPsEP8BbOfE0nx5m
LBnGkbzrJB3A06KwHOXnzMTF8pU/R7BbH8nBRG+k/XexXzk+2cCplx1c1tuDYdpIflCJTdP6hrPe
uybXP1dWsHlQ5jvmbE+qVhrjeyHj7RRgWclETimDY52Zj9yfm88b3tCmNG4LF9wsYw+SHcGASFO3
M/7mO1k02oNRIfT2Pj/LrYz7M0bVPg1x/hU0vMPmZ8atxS6YORZOrV4EYbIe9gviIQDnIqdecyrw
GUsejqaPBZGWiuxohD8SUKnsIhon3/iQuVR/j2V1rtdlhICBy8OkVBe4jebwzW5DFDn1+7UYoDcB
azTJSSZdDwVEh+bN0ZGl5yOVrf4uEzqBGuTjd2q7zHHgovWNqcK+edQ0FI6Bb6hKIDkGQuNH8lHT
rAPmpFO6VM93HkDIGJLOgIFqX7PMeL0zaX/vlEXCTWV422A1mBehBgA1xDsCYKFjMRbGhRjTkUi+
IKPFxTIAuVERWst3+de9G08o8LnA4EC4VdLPM3uBfLtZdGCMewu2pdYrUYv11FcVLrbsEYHkWpCb
FxlCUBKLpODKH0zjT86mDyZwxkpvJzdxuAD1J3N/qGhv7ezYO9YZ4gYw8CE6/uXl89L16jAyHPT1
2d0x0mXcf7C/+aUkFb5MAkACuZuWDE1fKih58JexE3l4qvz8ZXhZTAVRq7Ujx5Yuuw0kwto69WYi
SrjBa2YBMIWDlyX6UhzrigV0M6jpw5HILMSlMtRR47NRFhSlq5tJ1zdumdPy4YZdEkJ9sodCwgfj
zW9YQ7Gyrzu5hqh1/6ys2kkva1yu3jMuwBt8XBeZHOLlwDks3RCN0kOhmwhZ5IOJpl18t/VTdUwO
fYQH1a5vAwySns+vn518NPmnKQAvAbpin01B8SOjmNO+NbYi1OPFC8UQ9eznCEtHIn3oDhxNMhPf
nNDiV4yeKDOvSbB+nMIE702C2SEg+VhJGzPET7xoEPzSCBGPm6bHinXTD4QuIvHGcs4CWicBo0xy
FfkizgJoCYqUj5nisKXHTRPLYkVgbB4Ba/+H3/l5E/9/J53cH81O1v3u8C6bgOxtW+ma2g1nUs4Y
vWh/3qxNxgRmjl1V1u6IPzFjjV1PXl7+Qg0nelWZEEg7B4yicgkrFnNSrwQZ3x8mMonyDb+j/FH5
b+uoWnzyV5KPUYZbrpX96Wkjdv29fFyOQPz86LIO/ZGK1xALWuqhFPBFEdNtLdTRVBB5wqW7Uigr
j8ebkdZrgtPPxB0YG4+/9OknYoRqfOcVlo4a7qNkFVAAiJpOstBvkWZBnUwSEzNyc47vGIdCINMJ
rAFnF7x/BrHx9LPczn5PYwEIfbMlnG3OpFZO3IcbcnKQ7NL2ErKtHagmU0FYSdhaiWqA4hE8T4Rr
fVZTAH9iv5bnweZ2wgbA9Tl6Nt840Ny6VHktX6l1mfpxXHYgGGz1TXGhIxb89N24Q5ZHU1204D+C
EaLM7l8tEd0CYzi2vTFBgPtZs1znYIwmWdUv85ll1tX0hfS7iB2aj9aEhqcb5SMgMZQRLnXpayFu
iwHML2Qp3br2ZYVJz+WRuTz6Um/ZOnIdEUN7FtCp7kMNJDPwToYL4uL/01lDfCDPjrIUSlZU2654
fiFD1zS2Lo24MiQf6cdTmus6qqV+/QpdX11znKRvxep0KdnHCC/u5xlto4ehZU1wlmNY6tJFgWYC
3HbJJqspET8ncfRw5QZPmMNgsh+YV95KqIwY5d3iPlwvIGcUCHP2ugN/5HgWYRg1feeWui2ytyDn
1JMrM8aTRKrSWleTtwdFzpMqO8EiymdIoYUww48SPQkjVLJL4LYGpHpPYDgjGNhUzWEckCqBEUeQ
J3O+muJTuqwE9e2blaj8yF5IADUYsNyy3h0eCD+K3pyAtGv6IA9kEy2DTwcsNyTEAUUxEbPhCG/E
bdpxDzDEu7jLI8shQzGiSZyNuGJd/+lxKV/8M7dsOzrrscl/B8N0f2mFxADGf/QQ35crRnq7RIWL
FKOKKHhp8cJZ8P0oMsqHLWHkeNYcyKBnktkwqZapU/w+oLuUOjz5fD+mTm6RaokPkaUnOmqVUCxT
+G1T94zl4rEKyZHvTg5DPzfP6fwtQ8vSOLxA25xxUeZpZymnHvOn1sPBsGiEFB0pcQFqybs7BUWk
CBCFhIcg7AKjxTuE1oe/VCAVbuOYu7vtIaiYBCFls5zlwwjKoN3Y7cvFGJjWM8X7E3nNwOzB6uhv
dnn2dDGYaPsac9XGR+KeOkh7hY+3EXigwenw9+2OZofxReeeAFNIVd5MTpiqVqekqx+lWREHznHY
5WKBp/voFHHjPlU/A9ijgaI5CcLCdDOY96upmHoYUGBIYYT/W2C2l3XklKJEcOt/oVd8fbbzYOv8
OemLpdtyWau+GYKmB/5VeBvoYNOErH2MYq5msB7DoA2AcFdIF9nlCEyqb9iGAl6TfrWxVtLRCH1/
Eea/NcT9r7G2an4iAQXYFlhZBeag1Vh0HdHvv+j9GPxguugXnyDZ6AoHqauUYE9PtdcUTaWnvghH
rluEXo6MNwSu+tp4TuFuPnbnc1uDGm49DFzUAECprPU5Gpq8sAxnabGNMNZOyvqYUOm5A2ANGNNc
F8fNY+oclmTWMtzneYafiy/a2AjQwWBvzwrmIILXHzjKhaJyFktCNwxXRZL7xUvh4WxbemRIby2l
jMpCE5Ok+vstTOPCbhFqM7Q0eKA8nHqyFCver5K8llFTbVgLykIsp2Yyj9MxlIm9Lhu9TZRf8Ep9
/kPGq7FnQwTwM2bYJDrmc1KX/mv1D4pZCmdkLUKmTmapiW5KJ3bHqsRjwbpv3p/zSRsbqcjT6nbw
7AknAQRU7JBY5eLt2PCIQIrjGosHSxNMD8N+oSUq4/QUa2190QHDhRte8ApcRe2rME+t+/eMsPdB
CxhNZXJIZTG6eQLd4mnu8JFyfvizj5JdZFRgYneIyQTrdlVhSNYXzk1c7Ro3UqjZCHTuRZ17lmG6
ABs/vPekWeLhpoedFPtZnRn7wYZ87UeqskA4E7bcO2ijDaQYpaSKKkNYQGiZXHU+dwgUdBMVji6y
aZKNwYrei3+L2cullnLJL/f7iOowttwsrbxjcmz7FTJW9V/Sdf9aWfh16Uj1OvUe4burUWd5CD+c
sD1TT4KAz9diV/KJYbdTS3iwTWfeA2iKAfazYC2IqbDJ2d4B8gpuIhfehE6and5wyU43OJfe3ous
I8CLrFqEUffR7C4dOdkdb57MstooIqurJIRjU/FcSaURaSb3MOm9PnIiCRXMZmCuM9QMBvvFxlrX
kD2dNl6qBtiIP1cCwAIM1gZ980vlJD7Hlrxajn1UJoXLGrMnMkqJmiI/Kn1Wukdzx5Q8d/AqJHoF
RiY74mBJJE3FWAgWy5WVRxDr42dlLM8Y5OCCceJlHSyOjfaO0oaB2PrJ5S3doTK5tdGZ6mibIzDb
bfdOiVFi95Kjl2R69cKy+jGQCDVx6u9/LqH5FbUnvcSfhOtWo8ZnaMtMFxYGLrow2a6dOeD52tP6
2oaAFUcCwoSVL3MYaPE6JupqFlZZ1HA5lyQUCTle/EEvXfasLBvzAb/kTJqQyLtQAaGNmUcYf/Nf
tE6ZXV5o0sOkYpKarUpbj7Myoio0+/LvXX/ykC0TQU+e2mJ4L72EzC1uRd0MXB+mHRfUFNZ21u6h
8gUiEDwt07/LJWkFXtoN2bvEQRIUZc3wtRkAsaxNie0A5e8OLB9L66ISDYJZbMy1KIkcwkCQWoST
zsacmU7HrdWiKozGMCnI+Y2DjPW+BNasv2+lNw2bsJpAbcSsFW/SW1vjMUbvwP7Sz5ss3YbhXrhP
EKMhug2zlBM61RWNMQy91+dOzqYlEM8+SgaBsfXtH67fyOaIf9XEkUgqsM+Pj8xxqewJn9S1wBu/
GHLKGHp9BxKi90tFYAiDDDPAkBBWmb7UiWsIOp9ulIEDbEavMXI8PPncsPzBw6BAL2YrH4rHRTMY
nh15OP8OcPmL2L9RqUEO/fHNYNA4d4PVqdyAxLRBf/mLalI/CrLzPbayTb0FAj+We03khsUFU+TN
MMazPw2PLoUvrzbi8D4f/o2ZqCg1P4iPuml1Zwe/XD3T1Mc+1Ag5kM4Nqk5jBoStPbKO76wArPpn
W6/AYuh0H1p9vnxqJar4MVS8hwuX4wcML75lONr6IODvzlOnLUTyTMcKzhcP1FOORbIhh/Cy4sPV
72Ib5zjpeO1I6MTd5Wruof7+cG5h97Ee00izd4TPJLSN7xTqj+8oGAJRMXzJwqalUNqXC+QWCB/C
NhMAuMzhBQaiXEDpfG2vVJdpMtJ2RkB4xZ0zMGUvIu2GoRlrs51pLzwqypm0z3h74gV6+yJrfyDS
0n2aO/fxH0JXy/mTmSZgRxew11qk9b47vADXcolKg9lCWkb2XyP8WEBkz7agnJjzTuanl60poWR+
yYCqwDOBKr+ZOngmUNMxDkj43sqqT5ntlTTegAjBGsAoY0dFNCw+eGDzch8UOyYG1PaNfWXsr8kw
F14bujcwayk5HIXu9GdANA08ossNr+z3GZSWMoMI8LnS8zXbmVZwbsUpvwaxZpOhWeDElGyo31+I
4OBlZIs2/ZrVYVglqtK118FK25dGOKqqxNpSHc1jd0FX9zHgwECSIHxbaT8D/fnTAYx6UZ0PHBqg
0d72eaBV0kuVFlrUd0iqUQzagtuMND8kuSUVuhqgK9Rar1LHmmb7D5sb8+3FCTUz1d1rcD/+WX99
9xhxttT0pFjCQ3f2t6da2M2Ec1yFoeH1lkcgYu3HoZltJc3Jud4Cb7gfBpJwDm3S1+RcDcZmJlKt
JYZx7JlAfniLXA23ykOI1s55WEGEypb1DPsW9j2S0drf/GZBtuoJaQ03nNqmJ9ScYMor2yyLp2xt
D+GWkdlCylCamISBjeL7UrGNrlZwQWUVbZZbZ6UXs1lyMqboVUYcqCYOXeABUEiKUmz1s+TftV5b
GawQ1CaJ1JBLKy2e28NK1Fw0qL9yctMwXeZRXBMSkfq7TQ+gGNQYKskC646gEGA/VPoAc6qbMxNC
I+zZEFHrv0qB4meQgiIIWnyyJiKqRw6aW4hS7HWn599rF+hypcgImjP/87wJdhApSuO4pno36U9J
RV4LFYyONOKLnjKAlzFJ6yHbLYT8j6fI7fAPUQysKZlSixlVMyzX250lwR6O4+xjt5+WVS/W5JR7
6Y2HIhp5qLRehs2ZNJ4j6cu74GPCgEyx7/OEBmqa4oZVpAePKJhq6xTBnibIAYDovNxZf7jOULq6
HA2tghItAV3XX8/LquS/Ktjr3QQeIIjUIA0pJADjvN0mS72WkwMOyjoOjFRSV8d7rh3wl26kh77N
+A67JTJPzg21f6tmwCKRAE1X0yLTxBL4kRkuwtO5VVOsn4zm65K+BY6wXMQYASIWseOSNLNbeSp7
COg48k8XTBK3SMwkeAkMJY5cnDkqMkIhZe8Rm80fh7lzI90bAjWUukoFhlwQ7k5pWY59fBfKv6UN
czrf8XY1D6FT68AUm8bAy/91e6fNDuBSww2253KikzN1gsC0XpWLrWwu40osmUQSCYvM16PcAuXF
gP9hb0Uan1Pbjnp7uhrvllofqnVjtLqqYz49xdkGKTFz/mqBU4WXVNFn4qYq4J9YK/m5xVt8lSYr
qJruxTMhxrCkxgymAfGTE9D8ob70dk29+uQEZGMu71BVwqDZk3ibfeRUhlRVpe5j41RGL4YmrYyA
A59D92O2GxjLkL87gaamEgFI+iEgWu0LpVnbxMEWN2ujNlzWyfftP3QoR8tS6Q8gJvpvcMjbt3x1
d0UVHRntMbsp5Ww3Evhk6ELtyi6l1f1TUBCRumVACWEirUyeR0HmNiE7ow4rKWtSAm3ozwxLHvj0
PcKlKMDt64QM8ZCK7iIZdB1SC3TZvAE2PdFrZUYRRWrN/9oDndlgo3JGxGgjrR3dUc5ofAIMGlC/
pPp0eJfmDQsSS7LoxySoFYeJjIlp6p1qRMBhPMdcSXP5tyhgdNb/3SDILwAYZgpajSVtesauQuLt
TdqFWEksimuL1g56dtjrZUnQc1rEuWYuPj9AS5ABN3Ni0ZI2cKMLTCJ0mOlsnmXNXwmL3tbS+Nxi
OYs9rVZMA4uSWwhb8/eCW3phDrpkC28/jdewqikXFojKWssX//V3DMK5z5bvQ52FEmY66qI3FeWF
tcTg/22ih2R89TrxOE7idaq48z5JbZt4+uvfeWWyPzTRq/gBYmxEOrgxZ5nqwEg56l9mHysAg1Mt
Co/YN9ickBvs06mo49ikBIe1Tl/zw4QpV7qSomWnqEEME1TWv0xG/vnCkg4wnLNd2pXlBdXrOK98
ddGvlXTQAdrP1Ltr0cHiEsw0iWE0ZO6qXn5O49XL/lCySciXbr5mcGnnHAZT0RDFmHAo2/FKFGJc
2MT07kc3I0zlUIDwZImft9H0IZLNmm0Rs6KrmEu5KroruTQKI5X1ieJsPGL+m1cMwlHgi7YdWNIx
xiFDr7JJPn+UugF3jtNCKJ31TlfWOQVUv2asoVgjNJuL1OUDscmBnfTOXW4PVf1/LOTw6zEeXBz5
mqa2GGUD5Z2wSwfWBhw6UoA+gB6RZPEo/M7+cq2RBL2xxDJj3bKGdP/ULlx1HmW2jyTVfldPVJma
U+jNlzvz4UXK5cTQZhbkJV2kv0qErsrNDjREsqrCuQIsi7XNrkUg26nzFHpSBQFsmcAhP19MHtpP
MXy9vERbN/4nk8rSyoZKh6a8kFbMCcgMVwlEXl9eaGokDE6dJu44B8MO1Zhb02yiXEM9Q5Qgcg0C
RPyyZ/QoUeaxDY72VrdpYmi8fc+R136LJf9okGq3ByW2Cn+RmI6WhXa48PD34Eynh2bYgjkDTNcp
PonjrRKtgCuebMRtSoASKnzuluJ4UPbWWCxwo/bcAMSnACIiu4WuYw9GneeC1qNGj5EYzf1zG6ra
F7mX11krcPiCdRY3ftBhaU9/B7VKzClesP2llF6AFNgDF2UUr3HBvyopOlrt9H6HJCevtoQrtaVa
9nRWMspFgpYhZELFENNc/N5K69kO0xyjR1p0tqtVsdtZjkr9WtBdq73EngAzPopXKmnIht5tDtcW
1XBJ0jtzRGzYrpINg04XWEdUWBSj7sLtmQu43eBYB8HvR0kSPpexVVddqC93WX9f1SYaf/E/0/oc
t+d3nZR7WTzFSTFEe+Q3hAldIzFf6DpY6GunLLzBoMioZ1MeRp6mPbo92BenxzHpnaorsjWfTuK+
J5GqdI3+l4led5gSd9EA9MX77fHkDskVdB1wHmbgY1sSo52l8DwQ9SZ0ArS5Vlst6HYj0n5Nj5uW
107dUzYzb7iWegUK1+F/8JJvGb8sBdzDNNhpZPYfUifsB4lgqf+4oykbU4+nuS8f/JMR5D947+gW
XVPdT0i3TpIhnH48LEfDrvSe4lgtd3qZMOj0cn1Km8vym/KLdo74EKV7+K0NBf7ZQrvq0+weZULQ
ypOV3QbSPfiCXstdtShQt7JxgWzqgl3w/YjbDqj2G9nVb1v4Kw88YrefXRIpvByiqDAa4RO2P4ri
eEKBVDZX7Je2Yza4EgmRRwG4pj+J3xYjbBESVVhnEYZO0nTWnQAzHYNc2S3Cax0jAGhAs5E7RWJm
XjaUSaMe156RGzoj0pp7EOiLD10a3vtv2MpRcARmWBFIe0OmQWmnLaxTlLAQ69YvEg9yrGotMlch
Y7yfNs5KG7arfDASpGUUOHiljN4yG+4qaqNgpqLlp7oOpRY2VWoxBMWuCGvwCO8YsSnodVjUXrVf
gljwtWtK83bu5mseMrWoYs/pzbUW6KV2wOrs2bubu3ubzvuL7ub+lE8HXiN+52suXwwUMmRjogRJ
GkufJfhCQgVsFjfxPuV+DFw8Zi9B21FzDOshQ2T4wPg8SuAtC3xlVy5dU7vF1aUrOFZYdBL1LI6k
IZRnzbK+Kx6xxPRmeT+Z0RdcKpZ6YrHoFnu36qOSpxzG8/7oLqwRYJ3L4J2QCB2tPJ9R6eqi5vpA
R5JTAGmPSkGRE29NhEgoA2jN5OYJdk39SBCOKfsAxmxqmmr0V+foNZc7I1Bb1MlAX3PjexCUXKw+
r1lHBVo5B5CqKwj66U2NwlX//519K5zNTHJFN+pwCm6IyqlykqB895Gtqpz0DjmrgLgn9cXvUnIl
9uOf0DEYEoZ+FJF2peak+G30/0xtSRYA2t4kGfpcQKO8R/wH9Sb/NUiFg8yI1JWrZ3OA6wCF6zrd
OoMdpkniAdGJgTYkYG9wsZXUPAU8OjPFnHLrAmR+uJH/Foqo5lnz3ubddM47tICXZmowhL6U9Nmm
1lUS2JtxFVP+x6OfiDpSXjNWT4kyZViFcOCIK6xjunAhHBBsFi7RR5IcwvwZjIuaRrCF89MCv5oR
iUNJOTsN0K9anLctoBJKxt7PF6A8MRUxh+aJUvchx/muKrxT/23VgZOTOD8i5C2CfDYHJ7uAHwPD
iT1DOSVnhKVG9NYJUNV1DMJEGgeXgSFDk5x+QhnSYpMV4+CmE26HQ36NTAW70rre9DSdKtYigOzD
6xL/aw9NpiO0ITfhLQBtzonjWQuJ3ujKoGU3wDFYCeamYd06NJdGzHrwDDzwe1lGnSWAnLJhtYny
bTelF2zXidfN7DscFoL956EoOn/6Q8gFopBnEAzZuUZgiJU4lwJ9ldBZfFVQAQpe11yJ5mNVbKc0
8MxTFUPRH4FZFzpS+jBDjnJJbWERuZTMTCfbUCAXaJSmAaU6e5DvtHaB41kG/W1je73kAjMDsbIe
gvARWvdHYdTzrnGU4uXBnl9WW+UyfSn6lmTOu86CUmNftL6XX75z+d4DLkbmSYJvNVdjm846RV1j
9O65+6Gdyl+HXlVM3nrHtMps+qwEJdV/tZDPVApceNiMAu+rSJHDCeZHElfr2fzs0AgaiJSpafLf
4oIJf5pjFIJtTfgTZgQMXNYESrJp1/tU4nERmoR4EM3dcMtyJwC2MRF1EaOEeM6eXCIhli/Mu7kK
UKp2wEoJDXPiyYeeAujwp1Rt/H9xlX95DxM+a8LJuONjJM7YVKDNnBtRXrwGPt/2EpTmoIyqziI8
l0eJquTy+KlR9huK3AqArax03ixSmLLKCqxqcLR/EEj7wc37EV0xcx26wRnrxdiyHrGKjwyPzE2M
/RY2QMpi22QV5vDqkfDE1+A7+PaVVaYVacUOWboF8/uKMZ/OvfX/UWrpwQNr/IIkCXwNPLLs60sb
DSB6k7zzTQtvuabUFeDPxBvqhrEmTubfAU1rL3NkevJKXYTlX/6GYrczya0b1/TgzXlWKp4vNumP
szotdH+Ycy5rXu/OrQx310jWSakugXY2w72MvOKJvVUSx5AOMoxj2dFxrl1EAajEo2OwRTvmj9me
oExoo7N6mwSqZy/1QMtLAM7VuTRQQ5bFwTUQAWZZwhd1rPjigWKFfiHHeAafb4KQpWqLMrD+rAno
+yCZOfG8/ktgVuKUt3t3rgB00iLhHbCFbPC+VLwQx0DOCm4Y1H2OZFwU00EsjMpED/NsZtYVWOF2
BBiVEPtR2BIAWZUPrvWpavzizh2OG8Vw4ARhoLZmSkhld5GL9ppPZR4z+D4EmZ03+QvvT6NHP0x+
QUOERoAxEbdSNimBJO+007TeIG2cadePFXYkyR2gA1SUhQYsnBIaqBWjSBYbS/wrDaPAt4BWyX+G
fwC8tG0y2RO1GO4qKnB5Z65JppZa6CY51RphkGBG5oqwS+T6P1GoFMrCnDu9prMlvGH31iVxDDvm
Em0TeucbXPw5ir3eoOA2N5IWnNgot2x1XpY40TfX+5C+e1tLzeEucnTBKn71JrQ9e1ohEbhn2AOV
tf+kFHSpPUF06ZRWQe5SaVNt5SAiFVgr9B195kGaZCZ/ns/GB75+5XJG7v8pMgXAHdkL3St1uoqx
E8ETHk+JjrQN2CXSlM1Sm80b9zjcNKSSDqhpLQfgoSduQDzF/8ZGM3Z/pYkEx96hzSfym6yCf9i2
LOlMej3CbA9Y2gq90IJ05/OjqR+bNtHesU4eFZ9ChKbS7LNNxvPl9VxQCNCVIToIi9L+arWRDHNz
O+g39X//BcGNSn8y5CPEQZdlYL8bum/9bm5RLnzCxwQTaPYU9UBAG7b/ktdH3UfvCeif5NQvmVUZ
hTQV1jd24qPS9yAQCNMXUxXNEnDRbkQtACSp0mwL8GTD8mD8Nuwt83NajkQPHhLZfu6mcieNzD4t
vjqSiQ4GlqI74BTehAmc27QpbfLfjzBexpC6hS4q6PItVl+7UxQwrcEFLbrc8CpoT3mmT1bOHjz2
TRPAZLxcCqn+T5QVu/1NRnXfkl4B772Q7FM3T36QBqph3RA9DlF4RtO9PkyoSI7Lqqc+vLcex4UO
CCLuFh5MMpsqOnU7ee3Y0V7CF0vtDHAH8+6UJ/dLcj52DKcZDUjt1htZYGAZQFBd/+Rvun1gmIO+
0mkSnh/OnBUatFkylJBe9+juWyS/QWzBRh4SKnGKMXOX6B93ey90vkh+V7VagXH1lV5u+sLya0nS
ZxbBdGPj5O8XHzHl+2SJ/qveNRq7H0S8TsmYmMFqmMteHew+ja4tN+Q28/nd0hEzonuI5th7BUrr
wuwHeqbzukZlnmFiVy2KbkixNqf7iqvGJcPEEBPz4UrEYy3MeiW2uILgkrItS9gHa7wHDCEbOtWq
qxKM5ZKnAMhp7nQ41CU4z4rCzVskI1IwtZ139oGT4XJdzGPyVhKYwF45Vg3YyYmX8zlJE2cLsHjf
L3y5X6eaPHzlXEd9x3CPvec+1CtzZHg3RUm+9H1Gh44OolqzPsqi2aTAm77UtMETt9DxLQ3uirmO
3IZAA4AM4uG3Ywe/W942h4SIbPnyAtpZ/hu2UZU34ZYV523D6HJjeeIhL9qdE9WXoI9S/KAcHM/g
y7ZLE1Jor5BRza27UQ85JePEaCdo5KO3rECeOdkaS3VK35MyYR/hLQZoAP/ArIOGREm2eiG3+Mtz
uBmdvsxTtueR3ICIjaCfDXyCqEeRbbHYtFwaVgr7pVLtBL9XGpKx5+Bsi+1JukbX2LjnhSJCX9fd
8e4BOQEIHGmasjkxEmjwZA7dmKoTMY2jKhWIGIbAfdWNNqHvx7snfOT8TUdDK9vg1ARHRGs7gf+o
nMI8u5VgdPZi4gAtL/gT+8KAzXeSGY5kgBNTbmCJc7q3Jkmy7xoEEZr/twSMxyLCX9w+PFLc2EfZ
y+xO7JB9J7486Zn1mUUhx+oKtujhTA02TGZtNuJEUs0RmW6k6Q4nZEwgcFzGnFte8terKdcD1L9/
LyO4kt8aurmHpS0MWD8TCRy1z0jb4bh7MV5Qr6TjvXo19+GhRzdhViLRIhe2QD3C2VsYXTENxi9b
mNQMMPGL2q/0KGTPkJ4MkwQRHK+oceEvkABLNm+6fB4qW9OywH+MPLrn8DWQyxlTPDexiWUMmrug
WEuNuNcr73qnNCWL5gWj+1VqFSkBHOaCWHmZNEpX7O2CUzLhIe5CkL1WATRSrK19ZisLJarroNyv
wf9AyrrDmwvOzWntOmNrt6JbN/raUSwsLxMawdRjwNnagjJiJIFJaAyeZCGpcOUX0C3Q6XiMhLtA
CW1UbmZiEjW3z2qnpX7EH+Ky6IEipuXKEUBowtMlQprhuCwxLAD1XAqNBsEGI234BgNPWvUc3D73
2cioO+wobTf2vEdi49WUW3ucbp4bk56L9AAHU0784noOCPa8QI6GCT6TI5r+LJB5+5m6zybKVKwS
GgHarx+/dcHWtY8sKxkB6Jtz8ZXr+MeIFPCQGLoWeKeh+0obI4I9/v2NGxX/3tcD2hlnAJ7BZk38
CSNNZezb19rnCgpIZ5jv2wvC1OfjYI6glECUeBZkXBoQol0NJ96U11sXuETuox0jGiYa5m/mKn7r
YrkRqsbyVbcIi1/j2pHtt8uZTulnkmyDtq5zT8AdeMYPBwaP6aChrQoKcOoygd0B+AZ553aU3RH5
8WuP1cv25lVW9uWw4k58IFF2rLZXuO+QTkm3ZxgaCVLQW24DMgJSHpfgb4cWoanppOce6Ab9M0xy
CDgN2iKySH1AOsdBVO4b8w8iSbuksGwyggyQcswQ7Qc1tTkwKYjGAlB9u5KexULk+NlSUgVahAzE
AWZPLnN1Ui6R1SWC4GXGCkGKX3KI6qLhnlU8tOT08+1QmVB4gnJp73o4gQH4JnG2CW6Kvf5pxduZ
siZQAAbRldG0ED+eEJEdRTsM1IkbsgiWfQ7LQDao7VCvt8TwHe4ggCp5sKmyz/Fray0Q+tdOYTEm
HfUx9ubdSq0N4offtDq3rW2/F++v8cKIdcq2gYJwD4aFgkTAfR2jM+q+n7Q59Fi/ZXapVIV0ZJiZ
B5UjtpKyjHmQVglG3aBaPtROOIGHOUeWTqIm1VfRDNq5s0cYdeW3KqCVPG0y1z6jnqh9tZaYkvWF
7YTVrKDJZYygM7AAcLl6glGJYjzHClysicjbvsfaBwODYGw7tBTymk6Z5MtcAiR6W+k5rwYNmTpA
FDJYdf7j4QenLsFVM1cEV0lNDfX/wtSFdQa82co92P6oEoebL0hE0SzxZD/xsdEAUiPdWtJAo6kv
qVnZLMlPMj0g/ADlbxnRDKrzNsia/7hW37Yc8zwv3pNVJxn4Skg+xpV0/6kVUPwBgWwuwrcXJLHd
OdpXP4pAWMgEd5UhIOWe9E6jqMW1yzrnRpyNmIHhKrKI5HJEi0SMAK/aw015bDDvGaOxCCoKKnvo
RQnT/Lb2ygdnbZszU9jhNVSJh3eOoaj6fn7Xd04KgOMK/f1iArRgwZhR5mqydWxgXMp7TeUSK8+W
4BGA1HCPKqLsMC8OuegflDHbbQvnVwBoDdnqkzuYN+iCaOABbIaeOpWiZzzbRthBYexq3PW1hxs+
I/6hP8Xuto3a2c44k1abbdUlFeuRN9j0L8N4+xkTah2kUNy6r2gvC7p2Ssgx08pk5XMu9ECmwktg
WX4jkRYnxUKn+iXohMoGat0LfSYyZqxVlkxcsnJz2BMQMsjCgXGyaFRH2ky4XerCxtaQV210BQyS
WY43FTljc01nv+jIlyTb9CZJWHNxYWGe/f/0GvAt9WW79aeCPaTeN3zIpS1bSLklQI0zAw7YlKi2
Qc/nVKXFxi+FzeeBL9n/WnF6uKCFMxWLz0UoRb3PySAfGBKxuZR7FWjDNHAXy+zwK2Tq/XF9860C
5EPXlQuTkscthrMmNZBjiy4VQhfsMuaiu3YU7+Y36LXOJAA3To4P53PT+NQZO8+HLN9CfU5GEoS6
6yOOidvCrBcxR45anN9VAfOR5f519Ny3PtPpTOsq9N/jylWj/kErZhiS+bKsoYgn/d8NEX/YAncH
n1MOIBw/Omr4edxKcpMfGQFIC0DhZNhtz0sUUMWaz7Xa3diuc9ZmBkna1C9o0aAOPOr//XOf01cR
dCumWL6TPEEUC+4hb7XSeuiCWRI0gKNftacff3AaU5oJiY2iKmqWiKOf2JzfwPx0OIsoTkRWC46h
FzkK0Mxv3p+gZsYO9hHfGGp+SbixtUGBG7eEBNVKEudCdFUDIkaMJVZkVY2Dn1XHMr+Sefjh43Yz
bU9sBQKOYuUwLkjuvu7MUguwHe0qKbJOs7XAJIrH2NQqbADJ14c//KN/+2qJAS93R5JwGjG507q9
q3DXqJvuy5iJURqIYTCC2El5v+UI71iEpfmRj9ce9xMSCtGaLYvwplgK9ecaQfaPm79JVrmYMYdZ
poYVZGVzyf4w06JDTCtL11SFe4wci7GYkToqS6WjXCI2Vh3446ClZj7dqP+ru12XSYjl/prSmVfB
R0XFcCBmHSkX3kk7Uoyxe89jmv3jFQJDg82LjbsvDvXeeViiPAzGr6Z+swDrn6LEI2MOfZWPtCJ0
xNKuoaphJkuHbcqm97PmB18T21bR/juq2iOttVu/kGr7CrbA8iJykYqERw/ZqGvX3Ee4gPD7Z8kh
RFI6ZdQC6mKrUQURhxHekv/EG+j9PvhWopLitAJpkbO6xYYUuDtXh/NqPbivwci/vVGPbrFcCAQH
feqo+G3VJTm5P7xhkjv/Zdq2VZ0S1jiyaEPnoLYeT0ZguXjhEh4/my2lsuM88VvIvofZXdloWIEb
oCLhKjaM3J9wPn3W0RMrUmLuzyMEdKp/x8SuUd8RSuguZVEuwHQ2JeDBc39GSBvfAs3ofiq+Xu6F
fYqVMWf1t4ETbKc8qVqWQeVx9mBmJ4PQb1utB5z3Nztwnyc4IeKmM0qIm0SlhP6Mcte1qCHHTE5Y
aut8efOcv0EUFRilQIZVs8prMABwuw44kpOCE9MHUa6pZxVpiEVwMhkDRuZXXV63pCwbBQUIj1xP
tipFDrmk3Wt061M+PkEZuVMU9cA4LKgUMyS+SpR30Fx4jNWPo1Krnm96lsQ9C4VYjx3BUc6WpPQA
J8EXUnXfJNAFQe9OS3bL1RNZPFjE65DF49U7mpYh9F4uSgR/qIYlVrgFwPP9DDV7xJI57CVkgh2E
4ELqfFis8FMlcwkXitiBymGuC9o/Z6r/pUHnHewSTTAt4DLQMWfvOgEzefDxoCKaqQ5waZNMPF23
82FYhkbZ481cuzdtfBYJbmYK6aULJClpll/L0hVMUKQ9be7yJUSTjmPAv9Pydd6liFt3yWpcpYE9
UUUhtfT6E4fmZX9HBnFd1Xv0i2rUz2VIbX1KV7q6sZuiXji2r6qXRzrVEszgBZCmUmeeyNowDwDv
cYQWIljVyd2EiBQj363OuB4MNbTyal5iawQ8bzaSNILDity0tHWsWt5L7oD96NpL7Gp+fCaG3rfK
NdavhwsY725bIdABZQRDS+M4azulmNxmPT94t3sf8LBbNmDH91J/rQfuX88kbRGKDfodku7GYr/n
YbBEO7pdLXmnxIOO7KAfRKTJc9pSYNWHD9r4WRYyXzlmmAEcUMA8LDlUpxXqMzxjN2itcUaBCMMp
S1ZMtjFhUGkKTdSKTYF4xX9RwJEUTQdVojYocMP0goP4A3VD+DL1smuzelC/TFut36OfIhYe4jrf
c/o9BceDwNAIRVInWyr8vbhqIWqIZpB7jZ4y0I8KIyva8Or5kdocIqaP/17m9CgAJdPPzjQPYZqB
IkMYfeos5Q9kWJkafHpScLyjUt4SkhDxZAJ/jEVy29G7qDKK9EK/X0NtdPcJ/3vMWmAtDChiW5VS
kAxkB33MfvVrTLhyFFPfMmTNOgdAjn6DY7HDh3krgnlVY6K8Wl36WlE/b4VlZ2mQ6hQfm6fk5dnN
IjVZDe1CT1jFft67kNORhgGQm4N4Epbumf/Set8J0+nPJ3EGVVzKsQefs4iB5fA/UaG15AD8rwN+
C9whzqz8QhLNMpifpTrpt8EECutKalRWraryKBJUK66C8kEAeRco8XHjprVg+nmEINY2cGoGGs8W
pbebq6izFkQonzLlTOESJKmRCKOzUdumMPUefXs5hqKimiNm39A0Zx5uyt1vC5YEoZ65D+1dC0fc
fG3pJQqiTkXq2hCFb9fHRxEf0k4OouSoCAaUo/o6/ptlgdxx6Fzz572d00QxxFRole8TztP4xJo+
fUNIrO6Er0WVSZEr0Und8UKxSBWn/amGWh21eRB+xSxZqO8CsbD2l8h7ZHlurpD6skwpz7EGVkXr
l72dgaF3dyltDZmNKAVh36AJSGrC5T9o2zRNCHKb5wkYIXdvc+76pbfX1NHPe4YTWXNhTWDu0Wg/
4lNhfMqFHOqFG8XFP+gMCDq7qRLwWvHa0KSMeSNVO3AZwf2Sb7n+fbHUSy99ze+ojYCCHyuLpp/q
a2qQC2XK6V8S60ambtnqPFtHAzezVcfDujy6glsAeRwVH3f8iHyT3AW3t1UGG/Dl5rJk6HkEuSCX
eEpdbve9hNO9tM++nCkft4F7YmrjHrkU6fjCK1NmYd3c0HJsSoSuIlwzEAmXjq9NEc8aNEfI7zk+
Wd0IkohdDX+X3qZ+TvLRug0HtIc/1yqwbTXLlAZJiwvwSEg+iyoCkQo4MO66bSMN9iMs1BAQzHED
FEROetPlGYF3kLP/I3eV8jnpUk727joCWlLoERKj/UFZSJO+/yrf9mrS4+CIKEAIf8VtvxGfCGQ2
pawj13K6XSuukURKslvGWJw6VIJqsqCn/vxVHERlBjhTe6ntKK1yeZRBNeAg8TS2ckkkdUcBuIr2
eT3aTo2VEI6M0WfofXYl+Dzp8gXq7IlXmbezYWRqqL7+/rKbhjdPI7np2Z9MRFXXJNU3eTFuasAT
laJwxr0gp2WO93pU0/zc/aPXZ4tPbcsDVLK+CoKZMQlN+LcjMBvjS/N6UzjiKzOwaeeqg4v+sMtb
ILFOFTi+JWiQ8rDepcbbQsCPby34X4M+LiLY/9i6x0tbvBbQczW4ZhWcOMt/u4UCz3Ap/47OposY
vmqNUSyXr8BqVR3ExpOyy7HAxcPWb89bYA//MS7ySXlDvQUWW8QzWaQ/nAKfDfN2U2GkOA9Uh546
6QF2+CDOPL5F6rT0wYc/yVqQ1PBypw0Nn3AM0x3bLvSS6e1cFnNXu2au1BEZBJORYYsAsMJfR050
gH9AmtoACmAmJAiaXWoaKguNXuWy7iJHIT/fBXqfeAAPryzCvJTDOJWiSjrd1mx+vKcflsbjdwaF
olpQI+HoYKETbeTpK0V7LZ5LKd/BOSBtYL912j7xGLSaz+9TE8Udl9TE+h12Pt6t/d1O13oteQTb
w684i2gd1ddswqBdt3h/7XDw04b692cS+KHr3aTlyeKcY866CF+6jOTiDA3fhY8/pmEUgDiEpzDC
sL/HVgbdva+NReULxPRcf4uhAHyOXgH42bzQBsodCJTrLpc1aLTGrBEkNg5uJiB/bcybaw/QndCT
MXsKgOFCZGFTrcTdnfVg+nEVpHtH6a7NTfZV5h6da7rdHfXIU48FFERoutsMdXrrwwuNoqFYiQ+A
SyviwTSkLfKAfOMhFDl+gIvyP83Lm6j6zEbVgJlK23U6gLn4omsda1gti2aR8LIPVgnmPwlgK6Ki
i2AFTaMyqpjVNFS7qbrrJ7iVy6lxbgmaKqTzX7lyjD4qxNtWEsr4KUPIiJ+6aOAtpMtQXuv/gOd1
WT3MVdKZIqCZkmHpdcx+JCzuqZKA4VcNqboqj0z6rJHpRb6W3tVai35nK7sjYMqhPb0jF+muuuEe
36V94p3otj56bZ4QxZxYcXnpQUIcyz0uSRlyvsGsBM7tFrzkL2sNm2BShUseQIaCTevo5oOt9U6u
OA9VqqG/z0HL8OWxMRyADK9ThL1BPgDB+3deORfRqt+LSkInm46gWhURmqHz9ZUiuJOhyNZ4ZYBp
kAsiE31wkvk5fqFxtd2DNHyCim1VQ7Nsn995oRFQUdyn7AfoCrVcYlA2syuxgRBOFL1+2WEAKPtf
W+9nYOj/x6tF9/jxQawnztvKnUPSHsVH+vpXP92FhMGeB9X5ErhW88+9/QkjAIX1M9Pz+YLuKcHn
86jXXsi0AygwT3yDAAuGrKNTgDL5N0sxCe9R/vLaZ9M4oeiYKO1PqG8TIrZwhNSYhYt2EM1uiKLm
p/msO7pkBPNs9B2gPvJC1FTO9TrA7XPwpYP6PeTfcQOp8g1ox64m2UkIwD0K2EKD61rfEKtBkuvh
V/0HidvNNXt2BMMEzMC6N8pm6KMETTiUmhISLPeUx/LxeCaJ9mMSHK2xvSLTT8xtNTEArRu0BKyR
e9+P/RPF8/KLMzAaDYWVjxIvTkrte+ofiHjpnD1bLM3eMwKEE1HQqN8mVifvXZLZlLMwQEe+hvl6
XNPgIdZLcUToK1ysAwEGDQykni2qhuYMODPykyLxxNfiqiUeFkLQDoMHc/FXy3AOgBjtnMH4qcwM
IKZiTXmSIa1xgrcCdqlQudjeY3aHO4AZMFK1tFCe19v+OjULEN1AHtY+AdeG7HigDAI3AiMJsmhV
ZHCdaM/GWqUY9431oPaAy9MOP4BNvIXyxtOyoDmv6Hif1eAyoBYemjwYS1nXqbGYJNKDkF9lV0fU
0kNJtNr2O95q1wa8KdWi82Jo1SlhI63qmCXzIfjzPcWNvlVRp/oFt9rWzny8K6K1m4YzKDqTFSyg
n17CUGXxDMNB2G6ODhaCc+sNyyUCn/rg+pLJLCxKdHM4Yal3d2ZjeJydxeTzCgcRFYvfWT86bMQe
joSQJePfp1zlq68ICTyuA+Dj9m38POAy1+h+/vIK/3Q50L7OR/m1RjPpti+pfNZHDbmVI6sga0xC
UHF3ktyhfN0sx1gtYlWheXkd+LQizikNabeDHBSTcKZpuC9AHCrZE5n4yx2c10TLjET7GRyhal4O
Q9tvqpOWh/VqkUewcUJuTmNBDTWk2aA7c4fC25P+4Lr8P4rAdgUmhtjP+FJnM63Qols8Vocumukv
VMUvPHVBpYPcLEGzF/vQbCAnSIcIqPH8WeJa4gGLxSWdX1qhwyyucEJ4YLCvQZX/m2AU+2KI1NQm
05BZCx0f+XSmJXCs5jZZI5Ga9qOrmuqsWX9791QshoocVzMjiV8ysjMiN7lAwMyX0OFPLyKta+0p
j4s2q0EqiKnly+osOyEggc0py9SI4YhOlf5eKob9SSPF7Dq9/FQG7X6EC87LNpNDdi5tBGbVj2y4
oBDu+R12aP4BuemSEJ7PFomuuBcq7yxTeChXAFYDBMZfnsv4tox9bdN3u/xMiBbyFVFhDFQjaxa/
jpAaY4bRf8W1Zg1tdkItN0LC/b462sARtY1KmDnbB309GFmGxATMFrbu7qmAe42ClbkNM6jxfO4e
8ME03wYhwrlxgavQK7EC8Rku2HW/h5Jp2rsnqzpR404mF6lU5lWaLbd1xUYam9/xp9IQkl65gzcn
Qpw2V7pC42lGanTVuNSX+arIclk5oOYVV7UB1rB07ugG2GT8/lD4SYB6UvwAWj1JREoxDYe5MfjZ
QUSkkmGQGfTDk0B7LtFMsvXgMoz2Qp0fLl/lWfQG7zvoUQHbZPNpTpiTJfMZ43DqpkHUajOeSeYn
fEMt+GiNmcn4iweh0jPuWH8lP/COJO92gasNQwto1v0QZzfu+Lg2JzpceP7RJbeGMYg5/6NODbpe
2mlW/qd58X8eMWXdLyJ3J12EOs44FYcwRyZ+eygnnmuwrI5wfTNKKGdol0BlV8l+kXFMADiEW6FF
fl1FQJaMVHK1rBIyEaELJhCK6GFm+tTkv0rFubYO4hoMnlZA65fcxSGk+pCOQHBpL5DfWgTG78BT
qejyhSsS7cyhdF1a2WRrgZzRvm5SXD56TOTn/EuWcrpqE8mrHSlm49/cViwhLBZZEE/ro07jfMIu
qq7AXOwB9fLKTJ8RbY/G925rX3Q4xRFyg2CUmTckVYheEDhpT13H/EMrogwOmYHOA2WO6+DumlOm
YSTWdf3FiW3NPwzs72+QKQsPULMVj1t5tFq6W+BLJ+cJgssfrnvDv4CybyPaNB32xWCWJS8H5lg8
BkMODh7i22sShzqTM9UxKaCXV7OS8i0y+qTQKhvCyFDt5U5GjJKP+JKiPRZzTRFQSQ7iR6F+WFxo
FNqw0Fu0CTonE1RJY2cVf1H2AjOhit3FrKR8scKWmgmoRwo3dbersEUS+kn/5W7qPjgTZbgrjN3k
Ig6M7EtDgk/YOVI3hJOUc15voMsm9FS/YVQmJXJnqroYtcs6Ctx6l33NkXgmoDeL3afMa+pjgu0C
1YVKBImDxVkKbuyc80ubRrHlwMtSqWwcjOx76/0/wfht59mE1FJe8oYQqiKdXsNxZdxAX3bPBRZf
1XVx6xrrbxf7/WLfFnF6jANP8jSKQlYedDxR7vUGDPo0m5TUwNVBCaY1lI/yjxzeCx687QYsOUZH
8v17FAZXRUrM7ThxKwbJn7etS0ZIjtIne2/TyGi538pfg2rudlXId1aE8cdGu8vBr8mTb1mjjxQ7
iHUpAcnooPGijSvuGDBhvLUTxJN9SRFVOd5hxfZer+10O+Y6TfBZ/IjnTK28p27GO5rzNxys/bKu
GK3QO2QUsJMJ1bOBSdimPWAMSVL8q/dIJzkPYdhTp6YBlUXWuTpFQGVaVgpnc2KLu5wU8RH62Nhe
8jA1PyBg70xx+N1SM/KqtEbfUHPslzliEZ75IS8FuinZwNyT/6D2JBwrCzggge1gsiHGn/A4MwO9
EJnAp/dVQVYhbQgmKVBDvPMnnem8iz979v4y+wI40S9m34lPZW2YM/vLY39SE1zrVLViyDnHG2Nd
O6M99FxCchGSNhyQ7MFZMvGwwwNKrt7fDqsZViY/Nq6jWkZ5jeyQ0E31xgohGa1KyQSDmYklBnyx
ELqxzSXKik76VJtlDv7TZZZVY2hFDkuyinSUw3EdU2eQaUOHs8PtU7OXG80+3SX6NQLhr+KSX1R7
lehVp60Z3GSlv00Gy9uldfegGWQGFX8vRRlKf7Ly5Ti4BiTlc/KSAoVwmKZqho6qoO7zFfkQpOZJ
d3oTthwqePHUwn4sZEeT+on43Wf81YTClkODQkhV97KgQEp82iWutn4767zmin8CikXcAp4RB6Ds
mZnR+elcTxPiuUt7sy0QEFruz5xgHAkzluVuCYE6UG9Abm7AMdhqYufDkdR/BTR9iNIWP7MBeHg3
FAISqx9IPXb8aAuUh6P8ejeovpgIrZ6/tpo67lw0AzRe8Zwlzc5QpvfWtpMkH8B7MIORNzjXxxzc
nyHZwpB3MoTCn5epquVLQZS0ilfIYWHRApKcYIBD5JE0Bi6fAGPBwnuL6VXpKXlr4leqqDfduuEI
mkjN8VT6ai1x0BAvth+SZaUUjoUJITvnV44UC09Y4yFdKaUYzAeT7O0yDODOMS70koiHhQozBDJn
VWrxhTGgjBLhd/ew4tWlJjy+vjYq2UzVQhp/EQuR9xl+c77pjred1T1VhZFdIOFdcvTMwNLh4PWq
vSUB0SPE1nIcYVQr4yOhh+tW37Fpi/E6JA7+UfFoEcpjiFNDkiLrv+SpRVI4QxUkqWn0eQv41RQP
Rthjxx/PKRB/MQV/EbypBxXFzlGBbsjNaSy+Ts0jBsk5m7roCQytiu4Uhs5ZEGqCVnVyXFNY8YG8
qQwkr6+/9GikVNmOKms0Fmmbk37x7qUD0W070IxFuWH9hC5/ewvF5Cj8dYg0zNumpION36ZLNTUf
c+3UkR4s/g+G5+6FMZo6tBbHeZqwiXWtVBD5+wq/Z24dR29jk19xhrhh96TOPYqMz59flWUi7Tsf
3UwawEDNyXyNP5FEA8o2wUzuZfFZ9OfkoHSReVyJHEAM/Rzr/ZCNvEHNRFYsGP1YCsTcUKFvJVcV
MhO9yNdCoS7tdiGHxN9ffpejsu/w30ksI0fQp0himxKutAH0zNX8idwragaspxHgSB1J/fxMpfBy
kMqbvM0hQrcpeWKXXGhLh2F1DHmg2ntMg1lDlm7V2DAJBdps0ZCgxupkQ4GC+fF2vZCrdlx9PUd4
bQObdYv6GEQzvJYxpLmZ0o94IDWSjt6rKeSqoP/c85o4OYDTl8I6auSLrE6hryHxkT5jvqVe2mU5
/+vZADajv1s0PMLouOHYVN9obk7lxGEJus+MQO1W7iQWtFX0B5u9e0Ha4ruVWEWn+++Epvs9U3TN
rvByKsb6mHkCO4LnzzHrJvfehteKUVk17SaIfFoeh54+XGn7zfuNUXw8a0zSX1nvQ+UHPpMEDxzD
ljKWl6rB1z4Dfd3ArGeiO98YiFTdx6LdBQ6DpWQcipALRhB6D7Dyvw/MtlmBR5Tawscko8b2VbzC
bZPl0tsHuexCWBNBs6+ExFcTJOYQmJE4WGwGYp9QKJ9FhE7zqA4f7EwCElrR98N/C6EYBrlurWPc
+bVNAWL8p35AiBOiDCeYniEdVI2GBJzusFGd58w/xA7lhPd7mKmj4c5Axvrcv74nMB4qzWtcjKP9
mfrBm8iWwZvimBx2z/p7pRTqFoLEbvOu8CDQTurP7RDHZk1VmqilCoOd+NzAOTnEevKA511cWhBX
mtMVMuQipPU5Nmi4dqt7VrRc0ZTolVI5f5cbUSNI4opgtdQ/v191rsoTBP5RvkR60lbxeEF19wbb
32idj9TmJhNWOuU06qbbbKeJrzbMvd8AS/NZAEbNQ5yieho+SdDu60W8qRCtZSZzIq85jBu2IFcQ
UxwIKmrKKtUkt53eANWKJ1QfN8gamdo6Ln6LOQvLkud38uA6DXRRd/N3uQo49FwgDiCLL7/kuT6l
vxr8cvSryMQc9Q27BR+zYDGxoSJZge1A0plQNnTxoWjupWM7F81/3AhkO4mFVu+PTkc2+Cc0VLOL
k6ntt1pUUw1298wWd4qAF3Z1LzTpYvD73WDI3+m2Y/ZavWF972QV/TbGHhYdSQjvt7py6+1K8Gxf
ENAp/rXSnopXkgrlp590Q48Fcd8emI8i1+76JcUZaHLPP24tDhM0BeL06GADvBJW7yKsUeK7U9Wp
P1t7uNo3zuPJiGlD1pV8e3Mr2gFiE4Khqd8eeHbaW2dTl5r4ZerxdpjwyTGCz4PDEekw1EH4A5LS
Y4ZecPmVh3I5RAarRVv+hwzFmUi8be7mtCKzmfjdecEa7o0JOgcAW3Gfc1fWcqfrwyOMyS6cbDGG
MjoEC7m2fWYlNV52Mb5iLfnhl0r8ylDb/n6U+VpYCBGkQKHEWYzqm3ZkSpuFs4Hu4KewznJK/er2
/Kk8KtmEdvaGcllqc51LIwXlFBlbZSbi7WPBeDPPxFnv9QtIoIh9oX0cgIydrekJUQkFSSsV8fvY
/jgCfDk4CpatEsfCn9rFwl5ux1LIcF8Ls73Wo1xlxzBRhp4qx3uWY6On+MYf/SlMVONJoal4uNNt
cDnywrO6W4WXigzRMsfAy6xECwqwXs2L0zPtvRW26ZuDS2k+ufOY9CW7DeztmC14VO0XwUyM2rp4
3n4Zc39K89/hjuLQbzwB+/ZbGL9cGRuELWnNBJNOiXyrQlpFo6V/Xm4mFk9IZv/3VexCn4SurOPu
2m1lRDmEEfdbxAwiIh1KH2IqA0oQyTfVsowa+m8msgLH6xzp3kyMtwWf0aenALkfpbxsxM+yYgOo
QhGGB6DaPYXf7CCNOMD8R+PEwuSd22e24nWVLbJNy+HaRdnehvSejY3Dzaaw/oI27hieTFYLOCHf
eqZvOgTMh4K9xp6LDU9cQB6k7AveVZo9Jf3rKcHhyyg6RnZaF0hq1hMw3rKqBkRRi5aajgx9Qx8D
CNPUIMva7gdErJaCnc/GIlVLHBVbMMLxnecZD2SAaFarqegGPbyEUhUFBqPuWHNIw0xba3UcW3A/
bXTl9eLsIkL5mvbMsTHeO2T+8GGuoAUYCkxWol2S6n92FJndPe13wp1zEwFSM//fOBUTG8GbXNNp
0j48z/IPaWZr7Q3PuJGQh57I+AUn6Q1KX/cvuJ/TPIVUwT9TqomUXWatMn4ScOBXG1scQJPH/zvI
jeDVKcaWKv2oySqZTtnmtn1fA5RtF2tK7305Qv1ooYeBAgscE6avC2eTCi7GaK+KUTyMXCrqLMTK
Zevy8ZTr2S02uridnDFwMChCl562PXypzq6/1TCG/YkMgLY7ZnAFUcECf+LuqvtSgXuab6PFlnMo
wVoi25GScrOhNLXALgdJmI9uOgK8QoPF0Itb3+/Ao6tknNjI3Z7m5qO5PnDtF9eJk0shaaliQvtg
/dvznJaDO9RBgeQ2mkirfo1DXwhcSx6I6DtKSdUAK4vnYWFeSy165ece1/x5OTfqtaWGopFf2q7p
qtvftKAHAMkhgpRf1UMLfSmeiuwla9o/Gt4lqqLOfL9uYLkP+eUetBCZXslfrbL6p7jyG+QsInAg
NsBzd6nw65AEVOEzc4vSKbTVLMKDpuXxL9IHE7ExqMNNyOYTA9JVUHnIoc/QUBAer2xgBHl0EDEI
snoSRX1eour7fNmxpd+ATYY0KClAhkgM60NmSO7rNxFhNPQFtYIxD/EQYdTXgbuDx7iQRaRz1jjb
9NM2hmwnvn+ppQOAeNdFmyf8B/ic0uGWUiprUCruuK/ZY1FVCZQ3FlaroNPUwgXO3tnLKjsLEnPF
eEjOVehC0XzUHrIvMo2Dk/sQH+GoSf7qHAUmhVn8Q5kQdrhesvSV9DtX8BvAEpXNGRtTsnZ5Z1A3
O3SKVvN7BCRgX/0/HGaOmOi9wzAkz9X8+76P8hDMsVDHS6fCinRs8u4tLEXkQ8n3/UYR1tSjYXIz
3zNAj3FApJpSXFtQnd4XE+Jkr75jJTCjkmANpugMNYi8rwq910EkydaqjYOmpqPkn+YEflw1QUzw
rGxDKsXbtSLpLnMCoxzlFtVNNvcTMcAsPUIyCPJSuFA2IqfZVMBMu5bxfONELki0txkUY+PdrWqH
pg9/O0hy8TGzB2mRPBzJK5i3UuFFC+5GY9JvX3bpl12ncEH4dD6UiNCE51JbTNUO3aaILP5w77rc
oB3aVRI6hvrgYiXmGfBNrtClJ66PgsyFHc78w6BUmJ+BJy5ZHAougAwJU3nZ1/jcd66dHGml/8B3
lW8OwjhbtINloIJUQHRtt5KtzqB3Q45MafLvQ6Qlm4rcIrehylbzV5BiVGkTu7t7w4Xtf1AqxRIt
tqUsMBluH8dJ4dnE4pZiJ12/njrB0QD+4sj3DqpApJvy+D+oAAd0/I53c139JP8KezK6BJ2S/xSr
7PXVnVuJ8CdOceXbHufR6FdJoDbNLLbWhKM/DPjSxvC1cpt9lgBQe39H6ivEfP6RcxtXccMbPTld
nI5B/nDFfmq7L6OL25OLRzMj9twDUa4HBy6lTLekjMxdEWU7Szm2dPShNAxkwOXduznsGUbt63/H
59u/BpwjRnXMLA+Rz/FwyifTtNX8UDOKZD306U3kwt8Z5uj488TdKPZu7WUKy08ly1UszNm+f4Xv
G780OD/A3WihaSwhWmFWTvzwd2Q0IGHvAnrs+oTOGTW/zmJke9DUzpXVD4dNXNkBuDObm8JDUe+2
69BHXsKNcE5LJhD+kQYR0D6TVOxNro2aZoNJaU9BmxkmYPS6pPc8V0xvPTGtQwPtFhOw61QxAD0o
DnQKs0zoiw83QLkd9Oui68ZkZYxPEOTbNNRzc3B8yn8XE+pISEZAIzggNC2Jee9EpvBKmHS/eGuD
Wtl9dj5wCmci38t06it4vOGvATG8wOlm2gV+Tf/md+SpDpJBHXWLbFWsWKiviI9Gdm3J2rVbxLjI
5VvfKkJRrfNz51s9Nl8G/76amCNZnuERFc8YbkiyM2WU+msdWwTaBY2d2fe0g89reFRuU8nLZjfy
fNa+JfAPMgn8yZs8dOP/VqQud8kzEUz9vuJq4uWuMFuJmH3HzIZbPoHSpD3u1nCqLeGLsJIwqeYL
NCHuPoybQUl7Q6CpCKsDedHvw0/BTZmjrzNBYCCasI2C3ODuRWcJUuIQiCrj4BpZZaY2Zb4e92Vi
UB8bOF0zmDET3bOqAaXW2+kMN5neo3pezDmjouwOCeBgFbVT9GFmTyTMwViek5FQnYLBGsSqEZXK
JdcTX8fCIfiUBCrpPk+UPbiWMrv1OWStUxv3hiNv9FRW8TP0AiZc290GVJ7KBdOkn/2vk5HEHcxA
uz2VXst9zMCuzlGHg68oYz4XwS/eSGJnxCuvVTMQqj+2UwoX4Z0kouCqi2vVAZNhCdgk0QZ5O4Gi
QOeLCvN5XeOdadD26CV/wBKYbH9RSAL5mbZTn00Hz1KZFNKLBV1ozukyqqOWxfABdu+Oq9mpef5y
Ovo8OabMglZPMx4DBUbUDdRMrRhkq3C46EgTPzDfI19HkWZ9Vp7pqssy9wAvFNT5j1DVyxhS9Wue
TGhYcFTetpb7ATKDPhVO2s/jOxAi3X7LAUPhpJRIgFKkawrvIuEDHRk2+GBGhqCd10f4YlJjcQSa
DZVRhX+/kEvkQM/Ex2vno/dU4ddMKrZ5B3J2KX2uQWRMq33RqR5myXPyFfKEk1NQwWPWtUHEewUP
4o/UHjwLOQ30HJcgWB2wQ2LlbIr89w2eLx2lV/vatPfcTKBSINk8QObXjJiV67qJudW/Rel0HalY
FQv48E3sWcMrqtJb+B74nyi3Pvk2vTwZMxI+Hq2nEJXcirk5kuoh4tdSX9XvBEHZ2+jUb7/EVDP7
sBjOJIvjmR15Ql6fZ4uDoGW7zGAP2nESz1+8Zs2EJzmGoMg6w+XoOtBnESAHwEAloJ5CTCwEHpa1
JSD/4whaJxcwgTOsOgJB86fvx2CAra/w8AtiyMQt0lrN5Tk4oJf99KZyUz12o3bh1F9rnDegyFYX
PDUwSpfIklmkF0cSi/pVMMUaZaKqFravys7yNKXb+6fWOuN1jeA18/wUt4Crdeh9m3xs8vZVmKKo
QveCF6FpCPrhmP/J+WZvsLoyXGPWz3hVvscQZpFAGWhYRUnRzkp3GgMXy3GnS9u2ToNzYZDdADam
fpZqg9XhPX2ZDVSfcgLesLWzgot2821gByiByEgiafynM8Kc1g7HCGgaf/iua3bxbzeT+WFNIJhb
ovIJCxzJ6cCKvUsdQT7cPjaCAXcY71a6rLL87SSKh72NDOTNhNpzrOgS9y9A+ae7IC29B7BeLATe
FpvNi/S6uTizL5slgCWcVYablodhZiHRl1GWsFMCW2MAH2FukGyzT3IelXJjTh1Nd8H7NbWS0lWH
vwq1ukkoZMQe0SCPARZ4+1bche/oMH+2Uu7iIJbs8r3o25DCVQXhZAN2M65m8c7sO+HC+S8DfKNP
rkHbWT99xt7SV2ZhdM6+lJnnQrRfe5RT2JZpSU+GGJ/25RYJATj+Fh5xPdFZMIcSiitXPppnH65H
DCd4beRqFQPOG2FM9hUlGhq/gR9biCJQzdr7r0hEzOc6MDgFpCeWx1BfmYP16R7rtb2ZKth8HOmQ
qVLScQj1zd53bM7j3FXvQ50NAEsbDd3d3LdcX/uTqwAm7MRJ9tL8QWXla2oODgnacNmH5pI8AfhN
u4ICa0f0R8jbMT9Lhw4iaK7ZEmvi/2TjbMtsea0QHvTKgf7DjGgHeO7hmPQq6zfiKeHpLwq2EfeK
0i9hd9XfmqjfY35SqGIrVrUdpcz2SIFrJxdmBVTjl3KfR33uFuYl4girDiIr8Ogq/1fS1xda/Qia
PBEB+6ZAZaSs/o6dLNGKI9VpZqfsCopmc7I6GLhj3zZ9vBNdTpu1gpN5hQVIXydQ89E/+d3l0rGO
pmNTS1k6CCMbEO4bIfcMmdOwlULSir1JCCzdtxTFmfV9U5w1FM/PXC4owEw9ccudQ2jo+i1tVDXT
Qd6VbnlehX6lFXpzmFla8Ay8kkQbDO+cthNHHnru7bDHOaK/600jFIx4Qdiw/gvWyXK03B+8Tn70
QqQIP4NZs7Yeeg4fAASrxtGnx2DWXjuyAFvP/sSj5QZdvrZ/jVjIFVusmrUA36ar/tzup60PZl6C
Bn5JRqdhaejpyeoKNrOOThLuwSmITlTbKUGjS2s1Jv0Mr0KPD+LQFKy1KijguqP2Ya4vulFcnqRm
j7RHdVGdIReTC9u7mH2YpTQ/pT2Peesgis+qKTF3K4UtR/gJCuDGsS5Olv/BuUJNj5rEDxYs5Lyz
UJhBfBlsZFlbAC1waE3gk//5Ug9PTBsGZCnQxMNiQlGETTdsdmCI07KPgmiPHyQq5n9UytX/XaKZ
RphdRUCzjEFPUkQTQ346n71kJ2LxbzdJIp1hrXcUiE4GPZWtDzMheourHOUXJpfuWE01h/+u1aGY
Xnql/0pS3NecN1rhm9nhuUZ2dAFn1lwDBYTT/WGtljo40M/aqpcTI6bodpsOfO1z+BE6pKNZ/g0g
szyhgsY8Pxv+mdPUkhP2P4fQK8HamMZwE8UlCGxRG2u9mluE/Kv2oaEAaL9LoPKwfzTE7w7ecczX
jtZld6YGR0afOhgI/fTizpVveULSaVp17ChWLZnYN5mcGBzRzUpyvOPA6o8Y17yOjI654QPlzOyH
brdmFxfFRGsdijvSkIqVC5xhbHo9biebbdOweI02UEIe7hk9diyQVNJj5hH7OVPvTPhZt76LrFlL
otdRAtqnLA3UljQS51i99Ui01IQ2Sup6RXG2wI0W/HLbzj8EDV4fQFc/btiAqY3YhLRYLRi+RL3i
jphcLQcuP2PkS/46adsL4wPByNWIVLcIaSiaSxainTqdYIU4bhuTfbpMoyZTUi/n8B10VLojOF5o
8Oli+ySh/Ef7zlCuR/rlis6l9sBX4uOr+MBadVdlBHeXWJecvmCLOaQSWUKnCrJ9X1gC/PziHIDL
/v5uiJXSTNum2OJ9aL3RWIU+6tNxzDg3frn1j87SBsoo69G0v64IIcunIHK+XvxZ5ibNiaR3oMd3
yyeoKAtNThJCExS5myyPzBTKmwa/VWytPeT0NMkA+aYRHuroLZUBGJiUdHT40t51hpBE0H4eOMSF
j8WC9kijJPmomD900vXW6mAKmXIbqZW0FqVGNGL04REpvBo+do5yDPNOPGF47T6xPN9Ol6mD2D/T
oaMILlfQbzooDFlhVGVwr1Pad0mFH8dLrA43TPoTIpXsc700BXoYHduTx/e8rf14oqjYr8r5GznU
3q1p17ftRIJmvCVrlnFgKYi2jyb02+aEaW6J0/qc+N4zF1yLv9i3XdGoqrrKqjz+bRVZHj9ONF8D
4WPwDTUiFifP17L7yC33WGy86cm/0XtvTgRwKHGr/t9c9cZkSlSfANKXY68BrVGl+JQdBsY9NauL
zXGf1zUkd0sDqaHsqS1qKlmK8eXar+4cT4kNCXdpK0Cbsm+x8FIhA5B+2qAGQA/yTJaeCkz6+WPD
RJ4TDXKRMbupr55hV8HFOpOcIM+iUS/mAgPSfQJWa0QmNG8PXYVbfu4POXJRK6u8C/gdEd8E9PKm
ej5pz7KFMJGT0dU17putzIjKU3qT8e4DWh++DwUX8fNfJ+MTWRcv48cpl35ZWN/JFz9kPepneWtw
EVExG2+P6rhzY0x01lLzbBVWDHZ44C2Se+MkJ+Kv+Ce+5jjH/auSfgU4czqDRGuPMqEyUT6oB5XO
FHoM8bEKbW7Y/ResVn9Indp4woQHWEM8Wm36ToPyEW64MuAa5EtFG60sd3XYks2q/DBACDIAMCuW
OzyRuJqmEh+Awpqxhv8CEclaH1re26GFVMUotayVEie3ljUMmDPyM2tw9F38RCNWP02OcdNl7U90
zSfPdanHMEACwOENu0YXhMOTKYe2fCOO/VGTBUbIgKrqDaQkwCPRIqI3Knd0Aqo5ULyFCmAMuTwv
KQMeWpLvXPdcpUqHJgx7Clhz4YyMD1n6HAOMqK7YWgYLi8znFh1l0lJ3gZMFlIdcXoQScgL5XxGU
vRUkZPQHRygsXzePUMbaUEn0eehEPeSGTWNknJY7dysDAIH0M/bZFUR3+UpILBl68/KvB4ktB5vF
08BVFKOcc+Eg+fZK8QPSGQwyiM+E8CS6wKn8s567TioTmuxfLuiUlSMTcO1SVGOB2HGBIoI9Dqsx
AzKtJ1USmmwyc7ycMb+LHvg/qUyirSObiREodw3PMj1T3AhgPtmr3ZogLLIDzU6us+VgZrJXYVfx
L6m4x1CgtaSMV5UZAlNEEjlWzvUUSf0/jAcn1MDSuxTa6IDx7sKAbRvY3I8BGZzCql4JOPqq/Ua2
6naaCavBkmejieBaP05ua5X74UTU7pOTx0/VGjO5mF1+3K3WNBqJV4oW0bvwYH1yHqVTQA/W6Oo5
H4BED7/LYyY906gzn3SfeM853k76T7i1eJNNOLv65VJ0gzsdTW46YstkcFjieayJ6JPb0BO1hKGd
XDxIou973fAtw8HiVYR/dUEXm/KpWSunqX/nc0T/ocNoA2sLWPS518a3jgxaiUL8Nz8WyErTgxJQ
kwna4/EBywG1RmjtJBu746QgfC52vVbsfr8heDYa+VwCzmjhCnQn2eOoXbbFfeXf8SeXP8p8/d3c
YV5ZAINmIKNUTHlX+BXJQ0fCYi6hiZ/dILE6Lyf5YX4W+wyaiA1kUTPNR9Xx9TKm7Eb80xHq1Rds
D9NZrGw5ruMMZ+ABuStHDIrZtWybeln+kcI/uT4yeC3BMr0awTivATSvTyAzGAeazNz2o0KPG8qh
ioxm2jjOWsmQQU+ee4QnTsWchY1MRviQT8Knas2wBoghFkaLFKpWOav8LV+Rv51f3CoIY6CNpWLn
ogtXeGS2S3V3bVQGTfE64wwp5hgwFtAp7zEeww8LapV3UfVEINTEYX1Y6lxxZTicF6IRX3VoPhx8
6ghr3c0VGJ0+8EgCsVgOuIYGlc/xn+CjTdZ9cyzheD6j2aX9ftFZVPav4GvyvKyZcvpDwAMfrbF6
T+dVcvkKm2LSEPkT2TocgTspB8OXwxF1xXOH68rpoV1cDCvY/nnonfkJkq5jldgbtTMJ37VhJBnh
Fuw1EJIRMBFuc4zaxb9nbpPRINcT7Kl/hN8f+FXDG+uswEbTUCZCeUGmFf2lxHp7aOcCheZAYf++
v70s4UGmscUkX83ybCOgCi4fT31QlXJ7duTdKiTlsXwyWCbnip9OtSReEd/3o5Z/xa3rIMpHqro1
A7rAahRw+8kMeKIGHRAMtxJwLhavp/NIe7eWU9PC6qOjcZpmRBSNe3S1fwzToFk7jHCZXeSAWddF
gF9YDkJ+aYKTXJFGSd5wfjFpuh//HBEdalsRHg5PCuXiTsOYYOkcRCsQ9IE0fyVTNX4zLn9fyWYY
ObADCDh831UpRD5RB80KJHeFWHnF2SZHI65MZrOzIO10dAqz8o89yGK/JMbSpLrGOp0hUeM/7nBH
i/v92UG2Zadv3m+S9OiTp+FwjgcOzG9mv4xAFibS1ax6mVbx3Xdi29PnNtdmdjS3nmdCRULEEdvU
mTEG0+hkPRLl194EJJ3LF6mDZyE726jkLw8us3eHqICVFy7cb7Vqg2TgSkugkJT9rrIvxEJ9WIZn
yqr5oKYoteJ+jSeTmtO0uynHawmqgHvS/qSIVMzBNyrcu19x47ErQnxhdwQvVY+pV/c/8hPYG+G/
nlIi1cuCxfUSdSEmlMqDKnlCOqM7RfjcvpE+7NGkPPZE0Y1cutr96aUPfUfDkb4hW9xHwEh0xd+f
0JAlzXRIZW6phsMAbZbOsTtxZosRtgMCS4LtuzT+d3A0gTC2GVGVRVgLcoHULDRZm4MOM5WAwiS2
WLCVgGNaCQCyW4DJ5Uyya7TtSLxSoXPW/7d27kkfrx3+QvfhIPrfhEM3nw76tuHRgMCu7EuSIzQ+
lLxJ23blBR2ssrpuksBaHCmP1CNI+10tQ8OWzSdFXJWFOXaAOW9czwuuSNPEImPDOkIpkSDQ9fKy
RqkHbiH4d+posYZM7s3qZzFNqZS1MNBx3hv/nSDm4aof75Cy374TBbRKWCYr6R/kRONGjH0DgL95
eU8zLyrSyqWoKYxtCVtGScoK6Sdp/fts9Pwh6qXdePpBfxjuDmpn0kr3NnYPbCGTEJYzgRKjGGQV
YJk8bMtwhrDSIeLpCE8Cx5MVaIjcpoNbkriowue8QORGSV+9eSSuPkGjN4wQPgJ3FsrRr0i/H2+5
XDFszJFP1wqDs10nAQJE98NGt5ooOf0MERBt/Yw8Gu9s+VozHbj7n6J8Vwf93f+weG77Bq+wwhQ6
XPhzKUG0FwBQqczBQDkt7/SzSjXApGzlrPqGBPz/zvzbRZgFtww5X+0lrRsxA/ssxx8It+wXnEHg
ESq4pDLsPdwNCUN5LV4IDw3vCpRFoXjWIBU2y4wGhBy2kgSogV6yyPExBtmQIFtmwQ2RpTkWSzUW
euNRQoW7GRH71oYNZ/0nJl8+pH26DhRt2rkN9yG+Ma6bnCizvilKuTi6Iwj8moMWagX8Puq4BBnf
tVCwUQtWJqe0EAzGRZRt5DyA/fPzKDvXj3LPp7nDj8DfOHNj2p0zo+gfF9HxCdwT1FHODhXRF1Hi
wl01cOdWbKjypjhxLoTlksGIFFn6vL24q/1XRqJcznJTS9Xdb+eGmcGN0t8nbOdrOQvl1T/0BZic
a9J4bRM/oJaVVxe6IetbZvhrOfW3DonxjBokePnuy4JaV9YiQxBN7Rw6nfM82KLeVqudgOsWDFph
007R32GED+b5SQcKcB1q5S+DqkepNDQzdqAdBQi2HMXl96OX86iTEui8xuoLSjYxsfgBK+jAi3gL
4J1HoMvFFwLk9FA2N77sazys00uLpEZI9G1Sta1+0Gpn0VD47rMjSdWOH6MFyC2Ka4t6hb6AGM3G
be7Tjy5O4U0ijx60EJYbjViM/F6S4IJ6hLTHyzz8T8Um9cS4HjwR8kADCWxbgHfxoYoB5nGmOUNw
kkaabkdtyp0F++MZJUKuqMLHjnh+M463TNpg7oN6AeSJoMSoNid+mBOTpp6sSzPUDIWfYX6nQ1cT
38ebTrzdOnCR+tIrHkwal8hhwmOAL4er/cmmsPMwg5IQIQJU1EdlMGkhUtQA8TBO9HAveLrq3zY/
7HbBJP2NbznP/yy+kkrWFlUPupD/WgoOnJIywRtP79YAea2Ke5R+nYpxoh+6yvKnc1tlUrGA1mhY
VfWB8yNq5H+7K8LOo60baqxo2WKHCD31cXBtfjHSOFIcuil4MTHKZCanu4D+JUm2Is+uAE0kNgxS
mYD6VSTWvZV+A0BkicBgIk5ohihYP0HCkeexgJcmF7Dd7CsmD4fG02XljOhIqvAYt5U22sn1Y/ji
6QsFsEGBxygd9GYYEOPrAfON7/2QVGBTtXXwSOWUI5FAvED2+twRgdeThr3AfKnvm6uJKozq5djq
OhDz1q7JX9eFDMF9TbU0/w0OHezFKAkAhWMJtcUUc3eFwgoO0mvbI+Hk87EChiQjKZybocT2OYak
AAuzgRoAGThoek2JNWA3UWao9XxTVsQs9TXBLzTUqRYzATofAMrFwQopH+1isaps857/Tl6aIIiB
MX/zpD3toQ+3MuF6MmT6Rdz4zLPxtIEtFamcKWUGpnwxWtQMVj+Er2Fo3nWldh50crBqyMpdJBOt
JinNfEaqXRxAxhXO5PbED+fKW3hf4lqU0WPor282Sa9uL/W5TdHQBaBqSk3UFXBcqhd/SnPe2L1+
J6iMO6DJCNJ/4W5vc5Snwa2HVG4A8vjFZ8H7iAQ6ahSlOWAOddPGjsALn577sTeIsO4z+bUxZ1pq
DGfuE4utIxf5+FZEEayRYyXEAIOLHO2yOXw9DBftVxQzJouf77d42VMHy/+PJUbg9VjRMdRjAHQv
+F99uNrDE7KZiGVBndwi5wWhxz2lQKfL9IXN6leTWR3jESNu+wsR80TDQDQLPxS6+0o7AnS0xpTC
1Wy62opsxxgV6haU9jWmxAGnDUEMug91IeVLL4LEfEQR03a590WFfFHXwjl7IKCmT2TF8AeopoLx
VUVgT+lSe8QDUGe4ses2I+h4WXOop/wGBdYln/0O7gh/pFfRrss1UxwcxkGS7C0vOw/hJgsw702F
PYRCyqX84cZalBVxkNohGiF3oUMkPUMST6xrHSA03xY91cL8ER3CdMVsER9dFWrBJVJtlS3XUHkk
CrrTJ8PXD54UEpYR1G1Zh7MbGWMoPiyXPOW+8jX55R6V2SaiI5h/MXKRGf/rWaapatpc4wwdBlbk
JGJVFlgzoNA8P+EnAUzD1AM3cI3XSfRPJRKikPg7aiwYt8dfJh2AtRajwzuXAUwWIv1MabOmFb9C
PxvR0cfCWhaEHZYXr1swdtujk3VlJpZVtpMVxL5RtpIkY+HMoyZWKGTcvxvkzFt0grEL3tsyjDo1
oIYet9WGiDiubqI1cLPRDGF1FghMddfEh01BWhRYR8oKLRE0mkAZOaKae7oXOVcgW/AuRw7IweAL
+CKy53JqzjCeJgMRC419qoi2XQ5vwqvqbCqAsMrGGCVRANHo0fan7TT1NIGSo0KLOm30qqi+DzYs
+42FfDrVzYURk1bwfjE8aEkUGYmCSGuezfMVoXPbo6sWjkSsaPdDZ48TWiivIgUzQJSGgHNp82Ta
wETVDCF5ZN+z5SJwwwweU9b/sFm7RjR6qIrjzT+skn6BmXBsUDyDxaaiAE8pAZ14nTOq69wfwfTF
4cZTt8CshvDrDhB8tmdnKcLeXCby8Qzp5Xy0LOcwr9QcnEEYAtp2reI+dpynwpzdsrIF29wbaF3s
tdZWZpyIomQYAcbBVikQvTkA7JmjyjyOleb7vjZo7+65ohOFVmyULThC6Cxe/mhkferpfjIiUO5p
WdJ1rMisOC//JfxZ27aMruuN/G4GruusTs6nCSDFBeMRwWNh31c5O79ZA1spq1cmP1rV4LY5sULG
d2DH6jiBtgBHHrWH9odMSAtCTP54Qfl2Sd8MVgddbjGQe9pXs8HObHgcbe+POvjqLJj/wzyPU3JW
dnJXCCn5z6xpHUioEY17JLEeYyS4mmmwJJdcN2WZ5PZRiGFomfVb5zMu7GK5HU0PMG1nvj1VAuQU
Osk0fkt7sdbFo7zYaeizFTppeFyCD15ZB4ekBJAclHQRkZXLJvdZdihzSWAIyDWYFo9RUMHZ1W0b
IU1roSt7TpbJFuLa1V2DnRp+GGL+NNnT1k/CUSx+P43qqiy6lxRlqM9oH6LfSHdKv4TiLOC+uXE/
8oItW8gAmS6p4Y5NaEu1sa+Ss8DQnzAbEcCUhZTwvNL+Hruq+F2EqvRw75i+IbWYtLS9+Q0hG4TR
+Oh7fyr4j/+yQiOrlyxYKJYSzvMkCbwoVw8mtXaGXvWvZEEnwPGyRJkeWPCIiO6Sy7hj0KvtTWd3
uiuJ6NhCnTsIFcygUKXI/TK+GHzBMcYA4aA7rEGIOxERLb9YFpkxbndT6WKX2OWQaEpUKUXzVBtC
MaWuBR9dtbhFNJKksWRxmPlt2jmoZ7HLw7MMWrS2X3Oy8Pz2E7A+CSF6oePrdAkzZ43oGcXf93Cg
kZEfvlsaLkRq6x+NzwiuBsIRYOxUGJgbQJ4MvBGum5f4VpyDRFfZxZZUVVZUffeNXK2oD4ANTsio
XOuctVLBLFakkP8CiSCxaVhyh76ZSyLOZ06uUzjhxxb7hL9mZiDKXP+4cgHKM9zVf0aGTl8ywGp6
yhKDs6SLhlm0rYO6mmXNDdglkepUbFr8yeM6BcLA/2Me0zKU/nO0uYQMDInIToJz+Ikg6EYfq2XP
CnjmKCUk7NVMRdDAp2GYhhO+EoKO1DdoFZm07ai1DcViZs65L2pT/XdQs+xcXJGKSKwczb+Qkhyk
6S7H1eP666gvWu+YWZw5kTsCbB95fEciCwwVvqTWGe6PGb6JeBalVIyDHXuIf8jjysrUIww7go8c
OR7Xp5zDsFOP4b9+lPB11fypVv/ogBOGcgBUWewjy4hpzc/yBg21flqOW04wdIPc/pkz5BuRjRDh
rjuj04CQ/bQy4ZrH3qA+nAb0W+SZc65DB2LbLkiEMcrHHHNz5b+UAWC/sosoQnjMipY9ikeDWHrn
NO9hTZZ/tQAGXwX+CX6SGlJgFecoI5/+j8l4BV3MSRTcMY7cHgsYd9d4RV59AtyYtsxrQ9fBA4OM
xKKY5HJamRkVb1UkJngHDnZuYWgf5bUBXrL94FPQrLXxe1krRRuj1BRiCFeZjrOqRGLbjm08iGHo
6E895TkzDQEPhVvZxg371OGjdACs3tjDyWB+p5Cfa9fU2+ruELMtU81pKe+X/Fw5BbYq6R5NPv4C
IM6R7DrDLZRRpAQFTyfKAGq6TvirXf761h2zYmZX3xnrWF0N+656xji+iyUYrRq7DOKVDoBb9yo3
Wf5upGvmNiDI1EDSChSeOHnxtAqtz98WWdrDKLOKhBW5q98Jta9SRRL5akaOyXIqsxDgTCYW1UPS
5PXbt5qXKra/XpjhBTKQajJdngq0PNgRlqkMLrs1aZbttcZrk/4nlrsubjLzMJP67KQKX5PQ59Nn
APq0wHGgmgCD7qPOrfFbA225ic5Rn6H92jnPKG/LcEHxo3U2icOdkgakGtmhFAzUJJMYCBt8nM8J
sBwmGaOpYaAGPGAUO6Q0tiLMQ3pbrO0PesJm4fbsiW0ZNem7uZ9A65rv5rMtM/Et8ASbAIbqT9DX
g+vVcwnAjpuIK4f0HN/bYR3yeasTQi/3l12Ei1+OfR+3neSYT2+AoDZXvgzaAPolfiGKvqA066am
R692c+lhkDmQ2TsiTVYgoOXiM6T5wrOlf+L37y7+pv0FdFiBzpP0QHgZ64uh7cmnc0Dctzy/7z/l
B37Jc8YsKYEOMOz33kNYEM44UhSRar5TwNnDssXiRTA/aYUiAKIj2SBtqhdJuXgtK/aL1qAkUZri
YPkoCrNaDkJ+4TQxiS8EyuTeXoYMYxKP0Rlk80ic4VXjQYa1x8sdxiQFW/4f8fM/uWnCJG/XX5w4
1ZPz4keSNwW99VGvmosKvfdizo40xP6mIWXohco9RxGQHDLM1aqpmUSlwg1NjvUETHei2MFKzKYt
BikaBB8jqP5SYoCczKG7HVeVKlJpZKSd7zRIzICqnnNSiB+Ann8Gs1wCtQzTAqIgP0OwWjtvZgtS
aWkXKHY+MUtLQ7P3XHM+6usUuNB2Owfb6weyLtBzqdwPFRYtdjooEzTNyjmCb/RQqNXegjS1ZwJG
lY+f8QCJu19jDXVW5MCu0v+HYvCEd/Ovj7O7uViHqzgSaGt/xE4IKXnM3FAtQaRJMB7xBw84pMQQ
f9z/+V3MRajZE2L77u2VzyP69w4KTbX2Vxv325B8tC1Y9WI6dd4kGuqqW8/aNHHPg95pJiUtsD/K
tQUVcjxpMH5lvgA1dd8Xi1VAvqyE46in6XqXYJ1d8QzkPbBQ9rjjAFIW6wtXJxuZd/ey+cAOGn5z
dPSfJUy1uxNGPuWnBSeHiLMHc6XN8qa5wbzW3oNPmaW9VRx3nP7E+/i+TabsB3Ys0JIYlqgLoMt0
cqcgzGfnLKxov+YA1JUFqjbddEZCrxlgzNkMYZat+zTRNR8kK1LvpOINmXAGckG+h0RZmtHje5Zk
ObpNBDgsGj9keZVqhpVPCLaTLajfAmUyhXfLei6fWGJfLy6TS7UZLphdT2B+tuwnEtQfyBnL9mci
CgB4Pv9rBwIGIawE7Z/WCzOYGjr4FmAZHQXm+E1UZeCtDtLWnFlnyTl1cKknuB57wwUB41HyZMtB
ZQNTmMgjquszPQ4FgAEIpV5Umab8EKKrgYIFyJMk8rCTkp5SAwbYgEh34V5anZNyU+Zvm0RcAIjg
veuuePgQ1+7dCF1CPS4l65IsM0Z4YqAMwTqOMtYFZXRKYB9RbYHiDHuWn8doHi3Tb4m69HESkI+K
4AW1NvD1BgqlwjNxlqH7jukEDki6BGceOssnj1HH1h5SzBr1EwTd0fe/2OaQYVYbmxOHv4T3bg8z
2n8NVduiTlc74vMv99+W58sCFUwsjRzU6KKmABmJAQoUilPZ83nAqYZG1tInMw0Vh+NdUXTXHAV2
wtNMynvnvZss8U7N1ynb+8tO6zyYpAKp43aYkT81rW/5TxzEEyHKeV2SPsPT4NULlSPJJwVhRWZA
LTuP72ouHQGb8O5mwvGC69Jdb2RCQeIGOUIHiX/8KTg1RvvT92VHb7qz6bKyWPYG3qyTEi64ff3z
r97DJxuvYcUjv3tDx3kHQyGhSay+83I1KEhU3SpwlFMR3DJcnRhLdJXZN5XQsAMMgezl+p0HQd4g
hNV2rS8t/cHII/j3JCWg2j/+RSedduvum4SGe61yQa3968gqRNv23NIjDpvqPFbXeBpO5dVVu+J9
bh/4kfrc5yWDOpvgoVPw1LkE6l/RCIQvqiKD0qPDERgaoRqMK3mai08PRsZnQ7etx7Eb3V2fp0Lh
oBbZ4kjQA/uMlWg8E7r3A7r0p0asTBIIgeqRnQEwIri59Iy3SIYS3R+OLmyj5VSaMhiLUL5An95C
s3VK0XzjXRBceYswyw+74DsNxzJAHL9toBF5sgrY+36pprqTu+jk+AsH8b+XMnCeHOEL9tTHufLV
w2puPLRpXMzlJPY5EwdceZJbHaIqV81Y9bohAJVMeqf0Uv32Q/eB8YvAWxFIrNp0wdUm2qGvymNa
ds12lLh1ALtA/OEWa6rgFXZPLy2OYt1eglZQvLC1z/Qg/ZfeFZniRve/78sHSD8xS0W4viQqJoGs
8PEGbNKu5w7vJWrrw4rHpWudBQ1tJgQ8G942tF3ZDBL50Q4eQNBjBLbjk2S0MnQ+bqeysEw8Pus0
k8Souq72fentp+uU5EG9DWABHR+V7AiyKUg2X6ubwHUfDdyXl5Hd+lnjsIzZqjNc4zrZ/uxwGiWW
iDSmgXU/B+QVjOKEhmdO8vBD/FK8gYynjKZBSDj9pkdy1uvIMsaE7BnlCPjPsaZtDz9s276k6TZ8
BRVXMU6ScXPQ/sKfZFeWEk9K1sprxmV+useoggm9MywH+SDqyljIvn/uCopPu+SOh5iKJe0Pzm2U
gLPc3UMKDrJgWckeyjEQ4YrHeOO+yKbZJXZpbSDAPuVXFBmuvY0eA5w1QCRdOBWXFnhMNUPG5/fJ
iIVNRJoOG2lwlk0OsGR64azz9Uo+lqcnkOAk7bx77Ap4zJFF3N1xwxCMzj5YL+lkIBhnco/v/qQs
yBcBevHNr7hmrHt4HWgNook4RFqsCAa9CHdAdd0ZUisM2FcwBRx/ebdCHzojiSdC8vnZ1gm8k2nw
yjWMEXzurLx/7qLVmE+R1L+/uS4qb7nYkCi4QZYelga4esuIYDlQFJHa9tqf2exy9b1EojOSYYL9
YAp+ud4n34pdYuIuTgU689oV2MFoZVF+x2REOLGujJfAASzqYCfe/f+pkNZ9kVJTEipiogtsNRCu
kDentjBNHQqld1nWPQ/OwipdxAxzJ6ceimIipYvskPFHM6mHDErZg5GiaOIrhzztwYII8Pwh9qss
sA1vQUHZ/dASAsdka2f8iuPevgsqO+hBQTlDHDpyvv+weqXB82cSKekOKdnFVGPyjGb0tbzQBuZ0
/mG/RSVi/0fePTDTn5RDvQqpMsoGOcdYUf5hmyoaxHPBOaRlvhTS+Td5AixnLJ2CkpQAvpTNOwPh
PjRpOVptiTang303agluZziTnqVT492+3YMbmeRTR/064Lam//CK460Y4jnwd56ip5smumt1pjfN
Erf2m4pWbCSuRwbYhDOegnuKqa6tLsw73s0rOQKmCAehXFbEmlyIqokm7zufSJl+lFuIOnr4Un63
YBq1LGabFJ1NYigVnG2JynvL16Z41ekfnszf9pjV0Rhfa/rww4qQsYuxfMn4TjVtDotM7xTu0JKV
uuMa88h8fncliHBAGSIwBAHtDgq9Yu8fLCkcQz1mOHhb3Q2MaO13BgqXmileOqZjXv8/Ou1LypaX
RC81kj0mm78t/EV8C1+AzQZxlZUcile4xpf0DYU4Wix0RQOmyIZbmlI75FguUGSCyo3IrCSexBhS
gEvUd8XLDqSAO04c7WNMGAobxZWmLzwvZEmmUY6xmYIPRjhQX3hXToITarz1Pv3iAQb7bHQV0LKy
zrQxl68IukDJ/MHmW07I5BIWikUu2H1TmCBAfIWCuTjuppz3HFYKsbnU1IgmRJzGEXZDTiCcZjXX
xt07CDvsQtAuq0xQXbqzU3auVI6srZM6IMEJyFC2M2L3msrio+/3zE+MCFPhUQ+cpbqMiqMSgm9b
c+M3W0yeF0ZZ1z8NzbEhUbfX29UQgqBW5XCNv5l1eyeR1W7wKK908dz/fzXN7zPwaNraV8bOkYWI
8AQM62HXlPnimTt/eo7pBEqWAk53TEHSfwxTCTiStpoSOgoWM7SWiVrNpWRdImx1LvH6q93pgsQ0
MJ96ByN+1YDnbcXr7L8fjOvBmKPcqTi8opvCpIrP9FU8DPj8ir+9SBzuUy5/SPxJPFui2APwV85y
JdxO3OJ+4e1t0z1Y0shdNpUHcxgHnjMLxv9KI+p9B4qKohZHFFEdbcX5K6Ks/Alrl/kCEIft8AaA
RuI9xjUtZsgzor6f4AMVjg0QtbU7DeTvcGBY/6/7eglY+E3szWWbCoauFKKvRfrevozmH7TEU9RA
toxyCeACNq0P/mF6XArYpU3cGQRXIt0I1+9j0Fb4u63CCE2nQFOFFD8Md1WAE1b1Wj2774b+khR4
uE5HgNndHsMiqR2nloxAJ71qmZDn5oYJRBwQJRemJ0yo5mkyKAa2p/yYzES9e2X2ZjFaoIH+W3j8
HPUFeKai0zlWyd6rKmWHCkd0BIWU+WaGnykAtQ8jK5k9VP7nPp80aj7UsDl2g3uShLlTQSB9CQ+A
KMlQ6mTKbunqSw1eCYuq6LZpdNTuIP2ldHtIw268QY4gB8aIXKimn5V9aFnzRVjq+oyi+F8XlTYi
ScteZ91cna5w7pqwQHmHkYnwYqrNnGfXNdFKyu6EeUAdTJlGjPi6syS7b+u+bf8Zca8qB0rTHY2D
HDJrU949YqboG6j20BLK6ToU8ItGxhBl5V5sJsXmaPOyenx/yDr8uf25V4OVOnUHTHVpzrcS1Zop
YTAIdsjSlrGbO2NmdlwSgt4S2xE4geey3nz4hM4hHsup8ESAD9BOhhD5vSQxB48egyLnW9Gg4rKm
4tDAOCL2c5PrjayeAZcNTcJxVvK72YCf95yXDjjUdwbc5oVnEqRUgpSER4jAz09yZNm+Q5JvZuNN
cMZyUeu2q3YJy+6emMfu9IFZvS5bRQy3FtZ8AMWFPibxqSaG4D4hyCA/VEyjXPiYmmpe63d/rhha
WhDa0ZIDCeO/C+5+LM3AwhT5KP/rX4HbL/HdNkNEcXiwQkgEwlMtG6HLUWyyznYgSp1D8V3ee2Vu
fD/kFwS1GhYwmfoPbui/fYH8Cjl3pzVVGZUdnMLLSx3YcMeqwVNOp4y6WHQoZwoas6I9kemvIIG7
SySwUL7n4MzecN5/wvETAnjlvdrxoKcsTNvOdTwsgps3kvN6Tq44rtIXzjO8HiNRL8iURPEzo/vO
ts75efexobaGy6f4zNehN0X39VYtQTZkJ0hCQoQ6s5IlP2B/nHbGZVaclV4Di+LzQLjwx7sVxMKF
UxlYT0gryPeHyaVhQgsOhledq7G+MFR5tA4XbEdUpafLlmD4xEo0fKdWmg7EZHI5QTNmtnZubfhH
r5gaAFnwBUaoLxGsozWPMIq5RLU6K8evE/rr+1pWJcykIcKpXPmr8lzTsP8AEvjmUDARev0XoGNF
P6fPyjr16tkMnqfXSOmLjRuAk6Bu0c+gOZD9iK7TqAt2TCDO2u58MurADD/B94alki8F9O7tNs8u
aRbD93e2g1r1bGvhRmN11VUkmOzN0NJGb2rXlU/ggoY5iwtlegaFnrPVAhwyhRlzGJrPLCpIigX9
CZeW+ceeQD6sy/5DM+bPtVbmoGmlPdZvm4rixi2B0Nvu7Pys/NFbPtElJuUvoC/TwEfl/dGPAzPM
WkrjYso/gxvFTnJ6H9fokSLrJ75js5hMIeIOpDByadLXMuMYJxXVykuB4rBZLTnBEih70Ehje4In
/qfhaUezgYLgPOHgnXZTB4LUx3YyJLf1AJzUiz5d90tPkrgHC0pGTugTVAh8zr+tjqNl/5qaGnW1
Zz9sE1iJlT8qO/IISxhUDy008MBvxe6bAB1zGPP0a1pGBL/9POvbKnSrCpQ4IRlqpA9wQMxe2vEV
zP2pLZXgOpJtY3jgeKAGtdM6PRdvJAcfHvGlTon3L4zffYAaRAh0oxN1najsC7C6TrQ5TfY6UFMT
vo9zDQR6/YwkHgRWvKOAZag7sEzAKRe9WMgbejY7VRIdTGSa+HHy429Eaag4ox1wWC72n4om6XEr
fcG+Rf5vCpmW+YYXfq+KfLlXjfhCw2lTlIK3WJh1P30ad/87N22ffCjcnWhoqO6xF9KCkBC7vm0K
f1OLca6kHwogA45VFuFP2lPx9lS33HeR0q2mAJQ5vUx7CzWRTF6GJtz2QUUwbRUzFX3uOS3Y8/XU
urY5alWrtRAkiybFrK0KHspj242cYvfbYN6VEXXucAeq4GlyDCT31aBUZawBI65qa47TssmIPf/H
v3ppJXlb5z93ifrmzmnE3lppCYySfAtopHM/3glDuNQ12QtfCTbilPYZVd6HdUPCvO3/glbawlxQ
OamooojMhsrnjBU4qNT6Nje/EYDMCgh2j0ygkQI6uDwOo61kPbWyH6f7RwejBpzDHhNAafU/p7YO
xPDrSPEkZk66Yg/qBev+mgm9SSkVxU+6fxS2RcnKXsLk4IiMKd4GxuQDgG3N6axELBWCMA0Jt5Et
qgn2ceONm386pIlqao3yt/m8dhSIqS3DDwyEzdcn4h3By5RBcXO6j8RYWojX61LMAynzJvdvME6i
A6sO+kkTv1eIYM9xe5sUPOZaYewMf8Mc9rg36FhgrgX17jKZ4bAbMCgS9g8ZEJHdxj8j7jdFFzWs
LIuEMhJmc10eJHsi2Myd2rx/rnd9pn/mW4EEJzcGpdelEN3mZSm5UMgAyjZLq5xoR54Omi5Zkzhh
XlMt1u3U1bck557f57WmRVs3umPZ89TvBOC9mWuNLzCf2wNLBXNoNTdxQdQ6qOP7uA3HodfxUXi0
59fPMKvQg3LsEWRKiJzoWaB9XrtZof1zoHqGpvbnL1iLXocBF05155hU3OefCH9C4AaYcb3B2LvC
QJwBoM58/X8Du657Rr2RPhjyHXHziFRqY5iYBVSC9pAEMY+0YJ97hXAnPOnHBmwaCyvunb7Y90jc
hgGtA1drPIPAolwiUYHJO/VmuDL4hMyYTiELwKsdPVf+j3M76SIhwzGP7m3dC32O2pX+/D0EEl2S
rw4PUpY+md36Ikagc3OjBcWVOAoFJVZpeQ/VdJp+NdWV6spPUuKJY+UE3enVraG1zod2/M37H2w4
tkJC44ArjEJMUAxGQQLA8LZNaEWT5/AKx/VzPb1QXepVuDWHDz1rTbK3lAgTRQjNGLMwcYU5i6PM
WMa24l9ssmsljMWsWoDQFFkeJ2DOw2z/KWBh86zmawfCcEcNcuEXcYbUvoyBtT1/bHU9ZU7Y3qTw
QnH1s3Q05azWEOcx8x1c9KPrOQAT9xibXgKQh6pBa3J6X54NusDP8EFNqRGBSRFqI7xN+RHP0wHL
WTIry+EKnm3xuYdPyB4bGEtN03DoX9FVOq+sqNSyRr8s+0y72P4CwjIb/72ZJwS0mG2jI1TNW4Z1
0Rja3ovueyBYfOSCUEFUpCuj6Rdb+0qVmkH3NvU9tKEC/YwdSs2WTdb69Eu5WsCs8pqz14DVzR3x
3ZiRW5pENgWTqrihdezX4DQWFNpzkmkRFVY166u+tT9pMzMXVnPCB24lY/Hp9bGE53rATurZBSpD
uZjDpEQ+RShRj+HGA8Kuqvi1sDV+jWlcNg0gm0X5xrk1nvuA878SGkHuO5/eHDXR+DhX2FxUlpDT
tXTO+zDrNRK/c4/PY1mFO62fwQAfj446Y6IRjRn4U3ZDMPqJh5C9HJHBx2iYUDt6SOfga0TEBwgc
kx1XY29Qp639x94rekuloIooDU/cyaBoQfZ0ZKkGCIS7/Gpd8HeXxE7d2wWWAtZ2oVNeASlNKy32
FUr7XHSbIg5BlW0gspCmIEx7Q1O1ecXbmCipBBbUwlN9l0CR1axOaMsVMSk2Ny3jqHeQ/q5OmFpH
ahRvUiK12K88rjwAPK9ihDiLn1V77cJ3kNXCu/6sKPWBQIB70QY969JrAR3TrnIyAHF625f0q/gD
FfLbWzYGcEIYrMqS6Mg5KLwwokKxh3dMPSVf/4DoZA2E0VwtsVEmi8a+MehIhvl8nRD6sB8ioY1H
KaptQv+l1uOsGm3kM9SoGKUQxIAcGcET8H8H6flTHUkQ1Cs6cfJSfo/43XKxsfPzNbYgzdh1DK6z
pgAvlsRhtzsy5RVrwFFpgTF74v7fTVVgMFGHHS5cEXAIpbSEfmpKOeskxWe5bt/Mhj5ejJxiPHL9
05PWxdsfIy2/P95cXgJ+bH6ogH/eNZ6FSo+eM6pOu6VtmVipbv9AQT4KvBUGJHwcKsAzYMM0+APJ
JaQ7upRn2eCxH3nxpJuEWlzDq94y/1VecYQjFWLNRNa0Rm5JBiHqRrSmQuZPfcrXaQbbVxu1TNnG
GhRMbb+DDbtM3ls/YbpvOGhh34VR/VXW+QcxY5Vvlby/2X1pZO2Bf//bmNykzo79R2Btm88bFufr
Dz9oRvOYS/RV6H5JkdV1K5Bi4UuSeY+2EKkbPVXgw1fRuK/9wQwyHMiO6FcvJTxqetD1dm5Ew3rF
R2b1bwKUDxZLm+vD9R2/xWuByQMLVctQ3HpaciUae2gnsgL7dwBraMkhW4zI4bHeI341hev6TsGD
WHtQrHr7y6hs52OWTyK6jplccRs1FK0gnCbKAFR+F/v66gsk1YwH0FbizbCdRpObAb3ARQXzZbZ9
uhmCQXDWCXxN0bhAuTcmbe97PkdC/EbQsFOmZgGKyAya7kxXTW1NtKUektBVYYx2WTuOGQ/vXnuW
lC5/EBFhen7+SaxqDP5v3iULJr+rbxQBWJS1lbUQ/t5IALMnuB1KangXqrBNWzUVOyCX6eciYF8b
GDy1Nzt57lIFv3VPv3SZvebVou7IdshunEbT9FykAX6kyw08l/Uza4cjEmpyJAHOH+f3hU2LKfWn
X5YRclZ3zsz1SyRLW4OIU6uqptIC5tI5nrq7gD78VAR7O9HsRd4bc2kyxapwKrgQ+z+4a23tyua7
985d9RdGe0iwH3TZQaYAuEloOtr6BnzM6CH2rz47oDPEKwtVjA0tySdlHr9nE3Rx9iY2WJYmFf+S
mC3px3iQ6FIH5hE4PzKVJBr5XQaVls08YulLPThH83yQtwBYwYR14g+qqFX8Wvulc6DLFI2mSFwK
dsCw+mMIezbIcNAfaFRB2HrpehBpkeDO5ZY2N+H4k8MzURIdIgs34F82xhdapdzNKVB3loQ/Z+5o
rkotfnjK89O/S9KUnlw/y7ZOg0Oyzb83t1EojP+D2DRLPoE1pwVzEhvpctjYxjwiLFY5mP8e8VHn
gAKxkriwLLF716VE8hchfQhPVfYY/8fxrIHfbdG1S8eDG35SE0c1zoASq242M1YPj21x069Mr/+l
1NM9o8geAPiZkEH9WcsO5SBtmwgzid7ADl4ywv/DVynjFMDfH/77ZU43mcj68NOOoS1W6CV4YwgT
vJlehgV2z7l2QZ2FJnZcV0cg2uQeolYrrUN+g0X6qTTHyEDQdPM+S+dpqg6Etfx7o71OCY5+5uCm
B0MwIAzKGbJlLL/5d27AI8Xdca1HsULY2mUjc+D0Pm7qpVFVGKVoDN/kEDpRNtU/VkW1RynfYxT+
gVGAfvEa0EH8EYOfmygJy+zrFBMUzatt//QTPuKIdJQN5oNG9992/HdhuWOgE4vLMIHQbuOKcAUl
s7SwU+ha8sbHJJU+ykroe9XAVr9PYJ+21Hw1s8jlPjVinMlC4bMnA3x8gDyYR3tCvL/ZWqsHnSPV
H9e1sENQIENkRdi/Jvc55yImheWUSppgLGMnzki53xaYU/n9zP4NWGlxrSlDlD86U/Nwxap+Y8Ga
ywCrDwy/nhBbu16J00PguyCX3xm4QVvBLmPcMWtkUAYO8Z6ZKPvKUy8d8rfybMgSMwImOLHYAeZN
dNhKU1Up+hBFbd/ZGaRcni6KCHMwka8fORMVHBbgA7frB3hclYkmCiHip39q+NaHN304Q//Mik6a
WgcMj+eqSyZbpGRvHBfcbhK6fpVYzWbRGlYL8pklgDPFeR/tjPlRBav2G4IOZgm1p8qgL/R9g7le
88bbXV7iXn2gQ0ogd5CFopIWxAAGYL5AWdjSgpPlQQck3yyYINPcTDDKTswxXxjf/+IT75g3mcDj
pAJZwL/tMF0ms9Mwfe1qDCpNYgIcbjTSb7sDq0dclPmeARjEEwf7J5ZdvtJW3DNZFN2+/+H7mxDo
BveBrBeIqThy3YmcUvzR2TE2VMCSgse4rjf9tvoFpN7YEKT64dKhUVRA0amxL551akFUW4qpsGZp
abtjGUJgpSCDh6pPvRUXGGq7zbXiLmNkBbok47OXFk22YM6XzgdE4yB/Ji1u3vakUrtQgHerz3sL
6Qg+oxdM/ZrLrg7UlR1ld01fEd1woLwY19YuIuwOsYA7kufBMpLKoHHkNwnxatnYCm3Xfdfvl7aQ
OVxOhIUL2I1DaMfkzu+iRjj9mlSptIofnytoj961UFw00yFyW4VHgK8M5VPv4wvl1KQj/EnqBQHc
xP9I1OZPBkBR0kF18KDLEQP5P+NikfSw0HwU8kHITbUyBEt2Gk5MA4UTJC5njy7rkr79mLUoDhU6
HuvedqOWls+0+S3EFcohvpi3ht5nIzfGy1jzOawNllvfCLNXXI6GWNNmdYU8hW7ikl/oKRoMi7h+
cQYtar+q/rRfmv5Xskmf/gVmgiBYYAPEZVTFo2EsKoMTi+EuW618ZUyarlNBGSgXIfnvF1pNW3iO
gPp7+c0FA0AXL+HXFrH89foMYIFoUYIBnUC7JZw8NO1DaNZd18jj+GaL6wZ4XCxiuBlqJYIzhqq4
E5Y2Y1JlBGsYITPcU/i4n4vRcKna5arwLVEdYZeLd6TbhEDyfNKGAsiSJ60kEhYBp9bnIz8atpOU
gnbNQZTNDSZ3z/bigQC4WL8bnyH0Q9iUyerpCnwi1nua+1Hf3nwkz2DzJwWkhU/BjU7dZNghaDcF
Bd+KCGNTkkMePnDl0AJ8coAUaT0Hytj61XUIsT+VPRJ+4aA7R5fF8jzGxG+jG3TNwDxD3wG4Qo+R
RVGGfQQcToMrWJrS+cIQlOmXheWJrR3Ht801FRpI/mY9uKwrcFzRQuKJfT/NLSBEFixzzigZjE3z
8SpA217VUva6GWvo2dPYofhWi6367nkDbH/VLtjPh37kVHwIjewivFw+zR642VIbCTQU3LebbL7n
cOlSzLgL+rZC/JPH5q7NtY1zma84jXdr2YIeii+937V31sA8lhUPX1GZbDrDnP/v05dwYXAT/GCZ
L3TeSlYkoMo/GwyIYXXZRn8C4mmymp1a1Pq9kuWMoTPwfEIHrKjjsuztOh65YH133Pid4hO2GWAf
xkDYZoPTk7/dvMYcf6bIr8PCM8ETiEy4lOYt+iY4RPHV4Cfmm8Vo1+ljmmm0B05OEemHympzfyeV
wn6pcmwJJQ1OIy45uAP9zn+a380FHVZ+2cPNZsXkGq9aUN20GzN4ah4LzOAEkF8eua5GJtkM9OYD
ySH6vx+oPR/JrqZWcRyjhZAS8xdxfGVL89gezPDLiq5nuZzVYFGf3r09jBARwZ1mXHhzaP5J6F9W
m2w6G6Mwdxfs5I0M/ROu0KNczlADghYhnIepeA4CHa0NYDGLFQW4hVNq4Gn61rvE+sGs/8dEHuVl
/00/yVXPZEaSDSqBf1/WRT7d9udaSy+ZjnHj72A/vRi4NfRRqLPixN3shRtUas8L2SuTBTJ92AJX
6QlVPnW9dGd/9njDGJRrID46Pd2pXA/F1eHy30pSvWOiLxVMPwc4m+ertvC/oJz7E5wA0Pd9GV6w
ATJKTlli2WPRziO/NW4/HIFKO+5sR4rj9O+8HMJX6YX0Rgme3ErkYIla9DR0/GIcUyCrRLLUSsb1
oaErj3Ieo8jE6FwlCOu5U11rBlB8JGKQVy8YlbDpu3gY6WoyWnyHey8R/R4Wm+EFbUjn9q5X0y7z
T0oNzGhnzyA/qibOg0xcb7+cM1LpO4rIahcKCNy2ALXbZ8QpIIsm+XHZsummvOup/8g6KvDXPuAA
JP81+HeitfWoKQe/kgiqKxbqO23iPtWNabNtGdtum4hXDNxRcLvfrgcSRcOnCaHum3mdfbQLhr3r
8nmlhCYO1wW0IeAhpUzvX7oKDc5oSHDdrliMg2cpeL2kPVsbqT5p70PFajfxscJN/+umT8vSM+HI
zT72L9iMWHLYagPWBAMqPD7zWbdO2X3oniR6QsJKQZVx/+WxS77wXZf0jKTzQHwQOhaQRldYVJxe
+uabad0ootlgXu1vzTc9M+0BZNWSr5jAgm93Kc4BG/07v/sVAf7W0OEfanBjy+jakn8ZcB5vypQi
pY/h1Q4upC64PRwvque8E3bb+RPF8U4t6QHd44jMQJTIKDlbc+IBANwzaWNL/jtix1+m+q8TQuVu
PpcO3mkXe5Q4yf4NoSIew4ogXWM1Ujw5mWuffclc+f3O6kJCy7oGWWpJKTQW0Rs/x1AY2YWzuPnx
RIPpBRJ2NTXVenmWnQDJufnAWv/xH4CwXYHrtvA5qcY8LhVrCPAAKBv02VKbvh4p8lm2GkTHjv2b
df3B7Fz/QVl36A6AALAucYzXoqLhIA9zwMUUec4aodyk9qdo8E/kPT5wVD99R9aUwVY0uonnugkg
DStFan0etVTWedg0h0U3sPYAVqkdoDAqj1YH+V2XP9BZhrOd9+7AjLHmB4Gs62PxfMJuWhg3flNY
hwBU8J6X5ScCreDWJ1uByHZTaIGSAsIL4APqIq1CzPmCTdaMyJz619m6xF74PsMacG6X3jpuSCRp
5979ubBCJHW6EGyobRY8A1Dcj5Z6vGmLL+vDx73AvhbdC+FR8x88z5yX1hnGj6NYqfmO64Wf/BSk
4j/2EC5T6ceD92eQLzWl+L0BorMffftJySyAavkPrxzSAhfKR99g8T+aLN6vRHIbiALEJHqlrbcN
iVPNZTep7E0m/QFJafs9CgGgkS+aYjxitn3Epdv82IG/irqyAP72SRtq8bpS67hclwFHEOm4ajpn
CKYRFCcVC0hjVhHvNDWTbT4ZFpJVhCqC2/uzwje+zXqkpDegxO/HgnPKErfER1TyMQaIwM4axQ5J
iMoKN3a3Xd5uDbmztnhFODrqFZJYjV7Pu8+WRDbgJWUmRr8HdhFRQfP+XuFNp+nw7X5KcjnAOPl2
/JeiYzUxV1isUWO+aWLHuVml/2xhU5Ft6qOUK9Gg/j3AN5x0jz/VHkD0d+jhH1T6RSrTzpLcLY8A
WaJY9Be282BM8WXtBITecRPdzDz/Ijea0nvHcIgtsKjOfKV07PCn/Qnu8nDgEchk2vCyJTUSM8tz
DHvQRkBk8PWD3mg1XFBugvOxFjzXLnoxV4tkJVaviink/RAwZaXfszOKldjAu7r5p/yTZT7BemIb
QehFEh9sd3UZoIKrU8sE1NX43fY1+o8mSXVxQ11HLcvOqQhNIFHAW1q0aj5WVKO+Brn3XwPGmAsM
mVTA6DiHHWSAEPyySrqRnN4kk/i1+YrOKA+t5R3APHuayxukZx2F3WrkrRbeBMPpIuYp2I8VuZeg
8mpHN2y7gY7fde+yzJqk4toD4ldhnrobRAfw3xMIRDqH8r1aYLQVmkD32L05fQwk7hfYH2+G6JmC
PSg9cKzbL/BDfVGkTNn/LQmVSeBvVlWhAddXj7tLYtlEPn/VZO+YFU0Pu06n+xXm88XUq1d1VxOZ
PGthkBnMc61KpZKWvP2xlJSXUuzskHyUemRKaZiZwvbhJl3CB0pwV6I6pIRKUiSW6jgDKeOXzQWW
TeYM4KhvW8mA0kaJHZ2dVBbOWeivEzJvdjgnNV6T/qUATKg2y2/PAQraFZO5jVDkLqI+sXJVths8
InIVrJMNpHnCQbMMsXj4CZ5QGiw2VH7FEw7qR6fgRY0NbzH/EMcSrCUYa72rQ9BzuFCK1iLAsat9
+L+FTe4JUUkFb5rqT7fxh3/t0qqVv+f2Xi38ZEH0DUduZntQ+QWec0vzNx2HLPlPoKFtWF0Izkw/
nrJBSjUQvbTQY2hLJpx23MCfuUlL1EGbdQ0uvRKsdxU03iGigE9R8wM2Zoa1IoDi2tLAtVElzZoe
LdT24JzTpda52KRr6A4mZepJt+7nmKUOqvb6AtJJzfnFZJFMwcajLqrZWI7bJ/LxPe5oTb3tJu4I
vOdBqKL/7x5gSWHhg/NUcgO9c0CoKxrH9VXlhogPb6Ff3mqIIfrVKBRGng5JgBgjMlV3/aoxn0Qp
NxjGiycwFIoUocBcHkoxBA0hx8bswutZEPKzaJVZXeaMzIbs07N33Qax3wKynhXBNIyBnyUzpUMX
RuMZj0Xc8upKtTBW5SmDxJfYCKpmmE87gDBglEmY3Ez3qFXZPbPipS8efe/hGkb3wR0RVDi/tA46
IQijB9yxjJY8Dp4ZChhfSgrvuSVdbPm8Sf9KiYgPG37wPFwu/qnC/vzzZXXaOpfxYX3/1TaOG1CC
/XfpVgWSNHGzZyxBNe9atlyiyn+6P0FbxU1safL6nGXly9JmF1qRw5SZDcwxVKYb+S5Nl4a7R8Ix
Ciska4rcDCioeWJd43XbJZlz9lrRPnuBFC0DRIfgI+74nWmsJeyQ6cq0MGcX3oOoYAJt9TJNjQBc
LU88ltVEmX6TGjSBnY4IMghWraU2g4esBUjkXVQauGYv1G8eWbdHldWq90LdvpUeYMKqYCm/coU1
Tnrfnzqa8PmSjExxMP0qZEaUDteF49xn1arjQJdtH+xJDkSS+Uy3vEzzDZy3OjIGzH0tdrzrWYYP
adEnaOSQvys9fOYYAve8XPphATF0hUoMaE/8KsZCN8NnnVWcNekprCqxiiYDUWMABY9u2MsM89X2
cSPC1mEROGqq399BQCwqu6G85fVJ3CNAFPmfM/4yOMmuM85uC/xt0shOHj/FOws8bfSfz6EyqfAd
1gW1sulfVxlXSy2LP0lIhUJ7zvyqZm2hzHob6NYhSJXIw9k/mHe9PqNl4j/CwIfVxlDf7uUeLxEc
U3dkCf32yybbZJPXUueSPxn1WUm6k/5+VEWAh7nf6k1FHEOu/dJXD38DBj/MGkZyLGfi4JVJUVrg
R4pGUd1Wjvvs/+Ue7CDLxYohUKC8W5t5zzjEX7up4B5Iq0XKhssmR8e0mHCSu9tBL73tWizt2pSt
QXWTWlZy254IyPKDTyDEfOBCaWQyLCvfA7TA796yTMAwZsar4c5XH3i8TV5bv1oekp10TMJ5vyxS
S897TLdLKklZGAt6zPgmbL+KfUCe9Uhc3JrR4kuKpICZ3ysaE8XiMTBYAgnNDuq9dcMBHqM5FmFa
5ePl5+UUh1djSiOrx0jYjYP75APwYo5rmegJzqHhskiPGaQ/Pq4XjdjdPrXeVXMawt72FBJsGEwz
Mz8hElsCotXueJLDIjvKioThFyt4t0t8gQt963y9OcvRPPd5VmGk2+DBsGMyQ200Itq6oNPNHit7
DBqaZwoJ1Aek0Rp3bwfMHROI3OT3TRlwEovgUhJG7QEsw/C1R860NINIaNFE5mZJq5ZV0FeY+Lef
H7sRubTBguEKmpv6Xc/zfGsBpkBZPLHYk9NzPEFhEgv4q77XjfmycWuf6feFMaWJ1OhJuuJoKYLA
JP7zo95rQbW8Sh/YFGRTqmRzZHHW491ioWx4yxaoxEtrM0HQ9BIiMD+zD5dKYR45M1Or0mdAEPhK
F0oYDT08jd8E3GueOOZofw/eacFA9RZ9KD57Nbkna2bOSqNrKWV4g7iajMUAyU42suBlmvcIyxLE
Lt0w5GeNXyVHgqBDt9wdp531tSGqNGi+9IDNtSas4oDa1YipbufyF4YKxsYAYR1d+EuzFFrQ/5Ok
bRSxrfrUjDITq9eBb9YV2zMNRF1q+s1t/eLCnfQAhUJR+iV/eqYQXiGA+xKWRzVDQXZG7/2Mxwbe
bdLYcL/Mxiinl/nH/u7352/L/RXIIr2oJCVR9JJ8koRdebZ4K8ri5qs5jAO7FWKLwQDJ4lZ0WGh7
F+FsTv74ofiElehRHqceawvh5lx+GctKok2aKK4ADBCqBLWjiFM4Km+9jqzYKp/BjbgppxvvRlvt
hlPOZPowErFwpsl31rYZ7Yw29P2+xijm+VpomwPlI8jBj+B6ZhV/oe9S8MgeHHw4FCb2b8CHDrBA
DIC2GUh62ydPIQEr30H/0htlu+4e7ewQg8uVWzdrEM1N1vmcFoyPSGm41uP+CcPlaLsufuZEQ3+x
IbhPe49blm8mpIlJPZZV5Gq0hM2kqgc1SxOpiyyude1JsM4WD5YrM5EWcu+PfDRVUaySZ7/HTSUZ
q7PTZl26sF1f2tlOOILNTELvJzXNgx5ImIIzEcJYxkELW2zAG+52LIQse7aaSAuQO903TK89kjXf
IBge1bJ3xnmuITwARXsVNL/b4Zkbb5F9BdJ0LEKkz6HpPf5JrPaKGJedUAKAhCX3ExM10TuREOkw
vDiny1xbgAwo0dyq2PxkHl/izkNyx2urWnxkCMwMFojvS+wclf+FQFjfnoUOy94issErTKasvlAx
19ia8qo2IAJLsxZtJjxk17hLcts2uHdpue60UV3P7BsA0Ykr7+LoThhDKeaSYTvGvMbojer2SwJA
TrzZPYFj8deVubCoOUwPzWmzROnUSXLC1MId8pevXPtwEHX0Zd81gkBxnMXq+odF0e4k9y9KhHiB
mht6w+w+z843zYrzQMAZiF8W17WDVhHXoP8g/a2SruKIxVkEMQHBl2D4XBs+HcfUufBXq2YJqcEd
Ur0+lugs68s0ycFBRFbaUJSpRUxNG22kmmXPZAdfpjZfR/JHn0aPJelSmSzgL7qd66XrrG1CvSOV
oftjNbAzlhT6ciMWWjfRbA+bZzH5kMvgZE8IBKNsaDwK7G1cjTuRtpWdfVRkmgZRqyhMWa9zByPa
8IFQMrvCs0u2Ohz0jamXNKGupKXQbqQY7+IXq5h9Q0CSiZeemXxcBH0CRTamEHgeVs4IRN5aIMm8
zSJwZXGK7CNuD9SymP1/dVyjtg1GnHygLV6bfpRfizlIP/wuZfmdAUKXoyNn5JOVTFu8FOZdxCjv
5XQPwysWQqra/zlrD4AeQVWUA8W0osUEBtcVaolfx8xpyOku0dCgTFHldXDftL6YSAJb9TX3FX6r
d4rYvUpctqNENJOFje9cPbup2ikDSg4giK5fFp0gdRQ+SEhEvqLnL3DgTwpHzJmDgILVwJjMoSyf
92E/zJLl5fxV14vUTF8/hsnPq/bHFLoZ6Mk6u/KNAom2xju4RBrD1dYB8gh9bkWA50f79OVK2VUr
er0DkOgwhC5Qpqy7VavGrodTijAz1sHC7wgWFZoxc04AMRJNIoNbbcqsCgylxA7mD67+2/EyOsxc
LmdBXzfXgBqKRsku95cDpSsxHmV28dSzo3qPadiTCPeDtkSksee4HdyNMeNm2B8zMZSjsD2eD4VI
isje025B4Lh8b4VVZknkzQRUcjGAJXxdiLQP+S+ur2FshJT7KnhTD0UUxbMA7F17GEc5UA5fypx5
X5264EyPPV2rulaYmb4B0WIuVh2HQQCdNICF58Hx2GU4nuWQXT11cRon29wxDKyNjOczcW4xoamA
U9+Anu6O+CpGXnM1cYb/+j6t5p53uqcqnOE2HksTskH6eqE5TxMDVX2imhdUDqXwjnfjZjQcRC1h
q+4fyUsYlTSE/Ykl0G3ZJayfjKoqfpqWKOIlBUaR1JR+XL2FO9RMX/LZnlhDVov82bJ3bMaQAxus
AiFcOEjz5MO1EASiLiz//tJB8f3nHJlWVyAl3K+DT+YviWqjeBaXmccmhCKKB2Cegc8z9rBWZgx/
4fohAJq55XPhdwquSyHGZwhKQgmeEfe9W9cue37QbuZrcnFS/Dz0fXHYyNgK2MtfjUrzxzl488WP
bDwcg25+zgKuG4Sg+tqPysmVmcKEdwhC7Hogp2STplFLUdtadoZqBCO/D+FgSUZaBf6V4RkO+EAd
YAxmm0AQESvl4xXmfc2GyviHvQMcehVFLJu7yDzLWN9uT6yZxWYQiBAp7E0I0KDnCaITyt6V8Yqi
V9rtYG+71pl8el2LikKwkLo0TDKzKC1RSieHxeTVyx0TnSEWaM8lViA9lgA7vbg++nBOgD6BdD5b
v5klL0VgGRYROzfTAz37DdwNKtGklTB2DSm+VEeOzOTVW5RTsmkub698N/zVCADsuzqCikcm/v3b
SSBpFtLoJ84QYwANsipM5yRmvXGTQxftWuplUVORZrqGVCkfU8s74P2yxc0WOHSkBL7qby6kpEVi
DdExfaKmhuEz84+DnDzyx+nyoI4P74utSXf/GmXsjNFum0ufAnp6LslrsHQzbgOlq86M2Rof5+vU
p3ZI0P2KppCRKzhUzdpHvmkfOnuSLRq77r21ZcUkCSqnjplHWNDTBMfPY7t2yjR5RhyeEHelc4df
QDHOy6iA8jtzDqXMvnUlCmTkRf6/Yn8a10zbjrETu5FfuC3XdUGBCOGvn9uT6QEEQcV/wBWyoZmG
hTFfkWxeWOZKGNI3wgfjeGE7wMKWDVETh78A4drQmm8q37T4SrgUJxBd18HmRg+vWBg6jO/xsBOb
xdxfOWyc7xPvvqm/BLSOGOMl6cVnu7yTv3kVGv8gTK16XqqzUUnUvCKtGoDvLCemhrnDD/coy2PO
G3E1RDo+vQw50VjwW7JGkrRqnqooJwI7ypMCDxBx+inQCY0clBlBJlerW0ix3XF1wJzcnRGC6XeF
gjg8IRi7NHyLj2GFkZWYVcImrUPFRQAHBHqJFs7O2xC9+cXyG+hSkZJ9pdcLVINzOwIzu2tWwplZ
qv3hmQYrk2jZ4XvwR0Nnb2+ui4gc3naaLj8CcKB3GF90IhDaC2myWTiF5+5md9y6EAZuh7p5PWEa
Oy80io3yaC0UgTEWO/5v6DAZxjQksB2uVUDtrFpXiYQntc+AVKxf5uoZjbtQNcw2CvOIBXh6Pnc/
oscTem4tTFUKcQSd8K+rHEQwl8mH1hg0bE8PBTH3gi5vWOPjUYZs0gJzbrTLCwBExtqyg5D8q+k8
2PnOGzhL2cLpeesbHqVChTHwbCAkNylrw3KyFMGoYZ3NWD9I97/fZIh1fO/VP92tY29E5XSDQ4Wj
5yQ3RrpYOk8h31AK1zvnQpZMzenVyC3rGtei2p17h6KwH5rDB/wID96j8TdqogK/HT95y6RUtu32
Sv+caBSMPioUMgjm4ycBL5h/6VviMZg0UtpUUDiguwO6IJxa11351TLwzupaKsD0VnWpNcpb8/b0
j6KZnNDTkCBFr0BEgRgyngh93LyePiDX1/dLGk+9ltB62Jr4eQzNI8gT6vEZbA8NC9/6apXBCGgl
W5wP4OvJ5oXM1r7Z44/7lDiiHVIB7JybjZQvqJAbq5eOhbtOEIHQlKTCDjzcmn0cViMzRPCb1kto
bKYCXBr2uxlUN/VSGFJN61HzuY/c6fK3h4LUTDId2SLmL8XptaI4istJZzOtUKt4s3Wv8dXccprp
0QrS+A+fqAABr6dCMuMcZascCVf1YYbnBtFdPfLGuhjQwlH+tzPpkBPyZQB1o642kEZRID19xCIe
kDvntHdWSdmmEj6ret7B0Gf8rJ6JRCqve5sdhmEt4GykjNEz5k7s7f8XXI81q8TG2bO6D9lRxubV
H+212aDaT7SCEczA+QKJ7s6oBKiwvjAT4X/wuCimSbIL65pG1CJNVwIdRNg9qQzvGBBnNWjDUEe5
wfZ568Y9lRxfxuvHk71v2LuSnBiw6G4iGF2OCc+CzQNdjImD4Qdmzwq/c189lAzQXzAy6qA/Bp72
k4h3T+fXAespjWiO5B/4ak2sD+i2cQZ0nIjkp216N+C4TG3DZCPRe0awpWBbOZ/TCqsJiN/gT2vv
dOFF8A7KbVMdloRcQe+4RW+uaiQAcoe6sVuGVGw1UXkeqQOIjQn9LA5/UbVF1rGgWlzGSWw3uNq6
cLtmAUTekfufHnSDrOeJUSxnAk5WZnn3/IRyG8hHoO/i9bNfJQJawDSd38+krfOny4OzJEgOgbpc
WtomS+xrFbgbEZs2nCcLaXfjf5IMEsCbuc5mZIYqsOgVGNgWfT5Z5aPed8+Irp1GeAFD+cX1LNsH
1qWZE964dwl1UU9p/d3+FHnGg3nV0h/RX5pUr+lj0RVVK4Qvvplsi/88Q2juhC4L81I/QtRmMkEB
ef/d6UfL2j9WHlBooy8qGbH0xZXsAG3GCJ/a3HEOlEyHCGY93zsik2mn8lGMxT/Tu/46ImdVxpjl
kbCI5uDYJRHN4cVFK0RYpPWgDSfxpaUVErP6HEMQflHzY0bUMr5UnR+3PHQcpR1rkyXqcjlJJgLy
8RYoy6/M3l34wIg7F93ELHUexEPq958DTld0lprRr0UwCEC5v9N5x85ktI99WLBv10jjuo6sYqxw
PKpMHoPaFiX8BtkJcMxDwnVg0Opyldf6s62F25EAcJCLYTfBC6+NFCEnnwF+BQx9iYnTZmIDOIQi
7TZjSzgwQEpvSBdI9lzd8L+nmaMX0nSLQ8pY6u5TXPlN5vAO7bOy6j2XuqJ4zS4NW4eV29KlLIph
rHam365tasXY6yJTBkXmqYkAmhH0VmSqritV6VZmIdx/8QNApsFZTwycFgBzxZ97GIQTK+54XPtY
jO0ggeMqv5bnaC848Gh8XkUjo3ZaB4zhyr/SIOmHDUaCPS8WEM8SLJCKDZdYQm97IZUHZSciSB4V
zt2vCai/y4B2+go+5SfYkPUa1KBr3JLV/P/+irLdcnRB2W1xqlAJyrL656unIeJYb/6Qk3zAfzfM
gP0vlazbe2UghZLQGdpKJUKlMDNs7FKNNSJpM8ScKpItUc4a0H5enyF7jl36sYmqMukx6FniySxV
5CcmPi5/j879BCb7zbSXG7+zPP6w38Ilv2VCVFbqLjgeBvh5Co/eL0r4fpXg/rxQafdihqIycIEG
5Ox8VPNre/mvqVvRoFgkOIAe8eWWt8TbhLPl+nh1guXIWmEB0GgrPfyQ4xt6GvDcekC05dr/+IU5
ANBq6/lZXzPYYuHH8S2tS1tuLyKYCst9FKvsu9gOtyMacQczGwBSU7NO0VIu7rfmCuYOlZR3RgP8
DG05oSgNvfUahQF9IENHh7b4uPufDvADZDn55DCsndXrB4aT340guM8vx6Wj143h9kBiisrNz/0V
4w1kK+3l1qmFGMEv3iuu59SMT6qGnGquSHymr0OYeAiJPDKQTLuG/VbshHjzFye+7UumeP1Eopy0
Qy97RAAhGFl1pFHUwLzdKNGAGOB6IvKBv95muhabNgXdGhBE6DrN6MQmhM68Dxi/BNYahNcZLDAz
AcVi3VO9sH3DVnADTS95c6M4FL0Yxw1ZZFEDgVK9rEKe1xcnTogEAZNyRMhtdGlmInfP1rCyBcKO
LQ3vqu7RAj3f9FFErhBbhYH8+IcNZHlzGIw4EOV4y/ieAQ7C/cvvUOMSYfEHGMQsjHxLgHleo61J
+IBwkwy7XX4DksvXDm26VVowaJnFkBkJDwHvvoS1InU9LCeY5RGWRet1rzqq/dDaRHUCejG5ftNN
ozemDPl69OfuTuVHGc8WbNBd+GSmQHjhusGO980QuMl8r65iRpwEHWAFa9/gCGrVI8oyyEhkItV8
iqbGfYLhukFXdUR4j8OhCqM/ICZQQ3pmTMGh9Kv3E5absG/jX1ZxJl54qc1I4ZNnwutsKW0ETCrI
VcpxNhR0kq7BWF2Carj3SRilW0etb3D3fOiQPK6P0LF8M84yvBbvJjq6dmFcPzn+MgSpfKV4LMUA
jHJsLcqt3cBCVIbOJvlPUDjo9JudADNiuKl7mfonK2NMI3xaMrtV8miyYou0HvaY98PR4AYMjIVK
oif1a5q9qon1NDvtLPEYOKhHU6IoTDCmjG7JGmMXRnRnpNZVV1nKVWzwyvcC0ZkdbeK29ZakDMyu
RSjKVA59vGaamsOmDHH7Sn2GdnMGOMmuL602Mn+TxI9Jodyw8RJR3FLBForIycR8qbTwXuL2jSu7
JpAOneDfwD3eVDTTZg+ztOg1yQyowhpYJbJoKgcnIx89nDg0fK0ThoB/M9PQpxHVwGV8GxD88h0J
UvJsCzO3/6c9r0siwdMutRSIpxEjz49k/lkL+sPtw3vOo7WhbxsMJEdhvg7tk6NtBtxwelLgQkR+
3hs1bxrTeWpWmdBtM2w6wEa5mcJRyBIg8HSRWeDGk7ghdVqjjESuVpAXgeuynvzlVIwy9kPLV3Yv
LTdgHJqLIodPBnQSEBzWjqp7smddDUVEosFHeu5QkVoPbz0Zk8b7O+0Bqc0OpLLDxgxEsuUCb8gX
Svka8PO+jG9FbufdVJFQDmdNUgWa3AmNR726auCL/JsPvJpwZHUioBDIyWhk7QBzPK/l3HbR0Gds
B5pa67ylzu3OHGpL99SuogvNfW9sf75GM77+sLoymhtGxsCEDvNLIKQBzD2vBtCiQ1/lw7NBbiNh
f0UlmBAvWX5bGkTAgWoA9dWyh9IwEHcNyC3yee4UmNkLX5PFj8GRqQbvpC00boxX8dwekamQjl2p
ZpdNLE7albbuGVyPlzCj6ViGd5S07/jWjFMnhVz9++rwMWZAimyWsJ4tlIMhVSRT64tjZ9apzf/9
CSU1cMGtqXL+dFc+IbmdfIQfJ4oISjPV39+onJvr+ZJao1X87d7UKP5ECaxRb/yGskgIJPLFnEra
HZnJ9AF2Y9lNK+ew/62aVc4ndZBDi7FHC/8o3HjC8JQKdCW6WPR1s5qHm1LfgLbr2pnQp2iWS0w+
XRZF29zlOg7qkHBuEJz9xz8v6TiA8fqcHND0porMEN+acNZaJBSpVNF++ShgMx0xODC38q2r5r/z
o8idEUnXCruYZ+ISS0wSJ5eRMVPUy3cnuvaKOJL99UgwzWep3h+ktX//o7ymoU7YlCB6v6pBEwrJ
gpMOEvk/0Lpu9fIl5rHWAbvUVkjpXUM+yXpPH6nWU3qdjbz4dEMfqmIoKPWANMMueLHAWywU8Ui1
uJvvs+EV+DowUJQHpIvUOdQXHQHXhSxBC4jKxnKZgKxYS65mFVoo++hm+K/h9XpHCU2kBUF+UreE
i4yyFLAIBYXgrm+Oe6TCRSanOQgobbIrAFDwgRynY6cluJ0B5FLE5YElif29tdZL4dlnDxe6cF64
v8En3CewEkEBlFKmncGXjBU/ljhTe8RzeiOqA7lz5Y0gn2DNLBdKg3HMkikPWwoClX0jaf6mIb6B
5YyABENB55/z2iTQFzonaTcOr9ALWmdSqIP32Td6OWxirrFc5bRkLn4nsEyTCksRK+dCcYsVNc+b
wqK5t5u47ja0eogBCnGs8bBYcu6nUukCJx6LqHDwJLP9Ao+G7fM7KTeVcsVdKjvEHEQRx0j2SrDQ
tfl//rtdhdxducvBqaRgPtG/iM4ZDYIPzHwLM0fxFCuxdCZXDWTOq/uXMIiCU/tdsbeu0M0uFoVs
0oW25uv4laNANcYGtxfkyw5d9HU5H219AF4bzCeKy4YQ0SriQrHwvKCjeyI3yJGlZn3Xc8MdqVi/
Wviz1+Iw7oqy2ydiD+BJMffuaNM+ITtbtXyIaLZhFpHIF2hH5k/s2qksMQQAUjnQADDOy5wGiNL4
lpsngb/gbUTGIhdSpL9w0VrRw5GHhVGkOVg1y2RF1oCh+f0PfYcckZkixV1/KAcJj6vj3qYReum8
CsgsV4dB1evX2sWUcLHvJAKX0Xit+jnOWU4x05ClVIFPcikRQG9XBMOoMQxSqxP/Z0pQhLctjUsf
nFWNQU1MiD/ahTRJM1D1AaYueKl5yiwuPOb+iMKNszUWlc9KEy85RXdocyeoaH7hfB/4btM89l7p
nIk6SKyPFaYvsn9gk6ahARFDP9tAWuUJ9utoM/hbQ0RNg1Kkes6IlXaqOd8g4q6VCGFAzoo10SpH
bTc4a14LNWMjCKD9KugS9LbRNvFGW2+fyFaAFLR9sF4qBNqGKw12nl9r92BoP8Pbzj7Q5ubT4I3V
Pnx3r9Sx8n4BqAqRDPKGRlfxDVIPgYkH6ZBzqdQ7NE0cbz3Xi3AsVgteoi261IErdvwNRfVdhr16
Fh4ljwVj0IdjGzFtR3c0BMtmpOfWlAauPp4RDnysicFQtYqyYOKwSBiqYQAJ05vanNRveR0fRbpo
mJ6Qm83Tg0fiAJD1fDrH0un90xYi2QCCabu1c7fZjprAz1vT9NFLJuPmcxC9esg5VhX4xWE2sLl1
+tJ1xppm1NQialW64ixN5h/5e9zpI+XPsQq20D1RPmFXbeKzQRHBcJ3hVCBqpG1r3DiHVRAfDT9O
0z3s6nrrLITcpz3WUbVTM89beyBhGj+Dzprig+Y0OwK8FS+4MdfePg5Z5xCWfCcotmWvOHmGvcoA
1sgj7T86SUbD62QOxSbIKOn8p2oYDGugrOOqaMTihHyyAEpvc3lUY7VKpK8DEj6i3cIU74e02AH/
dAuWvH9KFd5VDfAgEQlYSkcZaz6DCp1p5AE5rcj54isnDiRhKkSGDiy7CEqretgiI/VrUvaXITh/
9BRzY7vTedoGqRXu2rKxZyQjkTg3xzmJPkQaPNhHbvJaUQz88BE2m10x+19g4o12y+hVpbIq7dGW
i3Q0Jl4BGIZnN6GcID7HzeooaMl53fUO0RF7G0k0tGNODnM6Gju2t9XrU8dUxupkS5f+mJVtgBp2
haJ2JOJejWHZY2E3eMh4SucmC2zSU3hb/2n7E3cswrXyX2IUHOXaYa64ilPgUsf0szf6obBs7VGL
OJnegsXsE6iKWDQOvBuE2+BG+vDDkiT7+UC2WgzEclu/CWkodTrEHyb5dc857O3P7TDZeeJOQSu0
vD+Jvrnd6MXXKIG13QElMHcMNY1+uICzDOkIPzV6Ig04KJjrvh64xX1xuytZStyxivO0Ol1lHlZs
t1QRi14EA0RS1RHDEcehNO2DWY2yaizmy7QW88/zRmohasu0FiaQtWazOKPd9H8vyleX73/JoRuq
yYPva1kP1I1FZKN2t5cM+3cyTQUSQbcTZlwcMs7o+7RwnhnjfumCji084kWl8OvXrNqE9/1jMYQQ
N/uHSJadj+Q2OwQDxJZFK8dkPh1LeXhuVwU0hewOv7ks1NeGnPID8oS4+01aurvsOC/gW8/ac04J
WtMYD3daOsBZp4XTCkFIjiZzYkoES/wIECqQwKJHcqrRPtsY0MBJzLQhuxxZzRJkDagUJnSF8b28
ckpIuM+ZXHDX62OVIpLrSBm8WvcnmST2Fqh6w8Z0C00eR19i1wV4DenQYt6mo5g+0M0uyWedWzSM
WKdd1iY1mAbh8+lgDLYs4TztABjffB+4O2suZE8dq00S9kHlcmM3fGuflNQ4dHuDpWsTw8Hpu6zZ
9BmssYEjMqYrzb4SFlGdIHXGAND3/sdzjZ+koMqkg+SJmOlChGl54f9eRKXwp5iUSyxKBA2qRSY0
KIWOJ6DnHXocwbmcBYyQckzFVKSdcMoU3YFmGkIo80uDCjYHPFpTq/ym5J5od+AFywt/N1svvGyd
MR7Rdar8+kzds3ymfh9ytD5J5Bmy1YIh/hh8Q0GQbjOWARS9g+GTg/6Wppn7mJww6qY2MxREVpNy
zFLhxHTxz7vyElpDHCmrUqpl9RER2GWrncyMFmXvV/ekCAlI2U1HxQ6ykf7fhU0RLi7KHRxiPxV/
3M9yAiNqoRBRgfsQxRPJL6WdhDGeOLB6GJBJ1nJ3a3xdsRVIF1ZtUB+d52DPNLyZls7ejbsr3fsK
TR7qtd8GzheyVTkJLecNwukfuva4MJyg1MzCIQQr9f78aDDn1BEAm2ZvwWS7Vn/XOSQckTWiS0A6
lBwEL0+YfrXfTMgkBqVFkfhr8Y2u3HarXk389jwdPdV9Ek9Ca8d/jhk+auT598ULxRbMaN1U5KQM
rgw3UYNGjNw47734hZfnPFnzqkfrNbcBi6YwogR2F0h0OcjYr9QrWQQHrsZw3RapnktOVppYLnOA
UWjZErosuqWinfRiD/jDRT9xjGqneEntRCPTLdD2KVeXb4PfGoGMkOmwlvivhU9fKYGiO6UvcLrz
zI67QlUCRFIwOXoBBa7IpsSIM0Jd+ZwgkrS0xmEiNkzAeDAsqeBGVuRPva0OjDrg/WQ4lXLR2Lfy
MoT44z/UFJYAM7N+aN1laUQbOEhjMduQqRiPlOzmKqeTAGxUboDfAkbqmxi0+DoMgFLwYcd8FhFc
IU3Iq5D8bNfZH3S2prPPqTrGMn6/dcPDdpCLDrX+eJ98GZ5wrhVunDlbcHv8KHkEdIfTdsI6QRjk
lfduWd22NYEOWFd0BCiq1qfY+uDpG5ARp+ctltItcGXW4513eUEyTWz50Qe8xBqXXCcpBIo1WEK9
RcbEZVuGytBV+kKiMavWXlN2X6s6tVNJQQnDn8NbE7mtcBs1EdjiC/kt/rscb+qrDRvcDCLKeMem
zoDUcfF42GrmbNGY+VSkZQNADrGqgLsP24FJ25+usY5gpxVtxWXJ9k1rt51BACLAA0Y+ZLS2WC+a
FnkbvfRdoBtFaYTvWvGnOfOKBa6mxg6bbKlUlnG6sT508JkN/wTQNtOx9S/bMMpzAybHQ/KnqTg1
DcDlYVtnggOktWdLXApp5+wjdQ0N+0yY5N1Oki5mriQe1zuD49m5frFJpN/hS1xSRChdXiTF4Yfg
O5/dLvMcBskt2qDOoQsBDKoMQpbtPZMUD7JCWpku9EN18A/1R4h553/0bmY39FM2ubC08/IYaMm3
jty7oNAq0tntc5bXzDv0vgfOR+5UCBfvI7GFAxBCmgnvOy8aCDuYJQYgHNGqPmlJ6LmZtAbXieGP
PFlrBH+AnCnWqepj6faTU4Qbb9o1CxstQ5U0OxLG/2bU2HqzoXF+uPTUmJSqPjJ4sRbvZ62206Bi
npePS6cRwWwKrna6iJqlea1kwwR9h+JV+O8kKXat+fXWQTzRPCVpAAOR4VoNqRyRuR1iKrrXeRg0
AHGaO9CF4NwoxvIquiOE5sxLudMJXvWrKMGobhtQvIUg4LSPUt9BTVL/mvKNt6i4MfhLO81jPwlH
1sEjGJxgboiAhDJFPtOedKGTMjpqiXjrzHFaU5QZNk8II/139Rh3vtiNnLr9Np0iEuspIM04lQA1
Q/C573GOIXIxY7/sgkSeFcdeUhXzpKQwzqGFpoZJTunAxi7TKa0vsJG+RQYV38lvxU5ClK7VELd3
mJeiH7rCyACkrzq8B/IwdLrPm3SSNPIqHKb9ex5r6FBYa7A72tpYYU6LI4e56BEUiG9wd5VxFxug
8A9MQuOlYilmUPfP6h32+DiQUucmH88j/UqF5wgv6xYo4JOhJ8OQDpKnpCCdnY3Nax8ix9C4OZqS
LY0FTtpggXjd7Kv5OlIjFoU8NOtDxFAbD1ZF7fh5VFtdToD5JsunV4FGo/MPeTpT+1J4nxgUf2Wu
RS6mwcjSV1VndAkzrA/oVf+1kyHXJMC6PZlA+92Wt1s95goNxBvOjwRhurgxhc4lora/rAsY26nW
ZUKTo4KJRqK7TxqK2RA77FfTQ15sly4qfiI+RhLcGzkdHgW162l1fqGhgkeBT1D09LjHl+Ov0KrH
BS/qmmXWDsAVlA8eYNzJnA8DK687RxSlA8kVtULMvwwQqsxytxm18wG4pqxM6rxfY4izr/Rrcz5z
gY/08pfAol5Rr83OzTQcP5MZvDCQTJ67K9ntrp6PTeX+mvQow0CRR08L4poqaHXfZoNl1I2epHrY
6uqMlJVL48p7CAst4QhkIq8Xxt2DBwedgGUfbpzEX/XMB7688UaCNKAk1VkuOfWKjRKCIF7CNZA4
3ELBf72NKaTraEtskhVl+snTLp47+yCJH8uQP/fzK4VIkvQn3UTQo2JLJnYDUJungch4tYXODBmE
LsWBcyS2yn2xcs5Ek5AfDZHQkhUJ85MAgwQiIR0trLOQ60nQChQ6n5V1615mvfnoMG7udrDH8s6C
jPKi/5M+rKPRuF40R67bYmDmSzZz73TKeQjmvzvaa1azWXCwZPOLoNieyYU4hbhxozDYVUxodeTg
wVmWAc1/KydAHKhOQdDlD5GcAVNIwG3ig3yyYluhTf7qLZznluhXtx520nePcdDTVhXaWoJnnOhF
E0TXWVFtJbKxozEubn0JslgQnP6ZH0E6eLFiFy0w2Zs2VDCWLU6Cy3HxxxVyeE/8/PjICkdJzkAa
sI1QOQwOiXnhHzUXTL4lYShgIt+zGEo4hPsSrygXnuGrjbSbtLigOefUhXYgu0ZVdgWgsOmT44Zf
hMo/fkJ+sUIovFNt2R5EJ8Vir5FRww54QVP/ehuztorSSKnT4Og33B33G3MwI4cP1VWRMWUqQaN5
OcailSS7bulUU1FYJQ7uDE5ZtM1YhwN20tCIECgg4iQH3+tA6lucn1aGu/tY1NREA/fDz1EMRHZV
HwDHLiGYbukHp9ABg2GzusVFkXecXJPvnTQDWY16eCKc0voqyc4J9m6QzFWONv+os2y8qEtLrRHk
w7VMINawXSxK8/vs6wX4WcGRfPuDgVqmyHD5YR4QGORd9nCxt7ld2AUV1GNrSRLpMmDPj5bavr7q
/LKEZZHqV1jT/t+eBolrR/mEIHQQ6nFur7KvgdpMH2svQtwB3l0hJpVHGkIDS/Nv1F3wHmsNgjzi
D4vq2x5oxcLvwunlyrDqqixmTk7vrtT7v8jq9zzpNkyF/tn79nWSkkPZwHM7o+DfRmpJ4ZQmFAgU
esUc68uso50U4mfMR8xCHlu8eNlMJhnJoC/r12wwQrmINokriv2M70g8XcpV2Xb0+57CPr577dXs
IbAq3ORNNbV7a0P8i+EpBLpIAwcy9oIyvxgUnBgijizATZ2THEY0JQdb8MkR/2QAHevll59Horgu
6+c6IfRWaBSW6aR+lxnxAMXgWWinNN9kDvrhixIsZJ5INv3uB7fzDpOrD0ffAxcC0P+d6EzHO/+Y
c9piYIqs7dyYDyDJiWypxtBwTapkSaWIv+kywKDmgqBaqUseL06S3HJaxWKuLozIZhwSngemHD4I
hKpctPLG3HEm3L7IbyFyotmnR5lyuaciag6bPHWISUlz4bR7Rtj1PjHyULeAh/OMkL9wEOGBByRo
5IcG4qleeVGCXSq+O4BnWti0d8MpSLz6xDdiY6giMMO+OTuKUY+aALdgZ7MYoODN1og3hjumhKNx
dWEyGvohsj8qmhhcDx3KjW03IPYxRoJQoydG6lQ1K6L/pbty6abWH7KukQ9Ev96a/Gz7UZwOqMh/
r+hcou+C1qHW9HhNEB1chWy7zlETZQa8gJHMIjdFJjPgAr1NXInEvl0OR1uZqJPPLZt8vPcWOj//
MG3OPQH2rF/9xTQDoWArPFEvI3Ct0HBa8loLCU5rmQe6t+SXlaVVOk294XZxzS9RPABg4yrnj1Cb
ffS1Z8c7wxXZWeWzqrtH0yznG5izEPs0fvBsFZnp/CVGVCzmgQL+gRD/+eiKy6X/XcHPmV/RgEsh
DBxKcKvwhSrzomM3XVTzZ/d6RGRa975DMLO3nBrjL6iJ8kthlDpA+aAM5XwDncy7d4B8KF6XWXG3
lIhZHQfPWKoPF2huDYQ0V98hPg8wglpApyUfaqGT0bkz3fR9VZQjxfBORvF7rfZ2TQRHAMNRgROF
mZaZjqle6WGrxxr419nIb4/phwaHIcQqMqXxBoGytIeOSNoBte7iF8fQpwfVqkGmMbHOBL9LfRBx
7QoseIHAxg3BOgRZ/0J6VxEIUOw78Ip76xcKLZxY3PHt/VaZC0OZQWqtJVzA5d/LsVM/u0NyCGHo
PxB/iszIFBdh88svduTdvngX1lZFiAv4EQVu9deSXG16HI9WPvsYhaqygvQReIswatK5G5PoUEIi
MSMB66TQBxKL9diQD0ZY1aaBAXCoaDWO2DuMG7aNGLq+2BRDz4eQv1MJEMWxICfEewZxxp3npBHs
jJhR0cyUypCEaLo=
`pragma protect end_protected

// 
