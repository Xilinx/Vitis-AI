/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAESMdaIlSZ13Xx1diNupudHmTc8ebeHmKUXLSfSeqx2jk01S7c7yA/Rg
lvrTkgIj+ymuokyHAhiK1UtYtGqjo5NOTfpXiEcaUl9KToMDUtxkRenPZdhpBQy5lfc4vq1m83gz
qPBWT9ZDwUZxQjupS70WuyzVAWvOFlBwFVY+st75FUvNPq3FplKzbDEDxeJgT2vm13QUjCfkUmmH
w46xz+dDRF288vaR5uUKGmRVWle5cvmiJeoA5RmWZHCYsa4HEliTqWW6CkfQV0m8yfJEfX0ZKFid
/1dF2TPUFXlZHJMskgz/uMM33M3dEjClYNgGsBfYLsuHXbHUPpBn4KV3dRvgeyvN1FryPymCyEc+
i+E7vh1+Ql9qR92gNNSBJRcQBXdS/o+gdxZOtYqfnrXJWNVnkPxU5rDQ1gBwmhjPbhXfo6z1ngww
YIEdHAfJ0ykJZtGTdCxapRKek7pftyKuvY1+8yKw6oZE2WlvVownZBehc/oYTGJNY6p3kc/Jao+R
I6/u1PCEXSwFmf/3dM3PTyaY23tpgXQWgsYH5dvoadaqSnQvKY9iItPiBpNk9D7OCPmw2UczXsdR
5OxyqHgMExYUzAZGXxTdHAuutcj4rpoDk9Egz1yhIAX/r8OFFa3YP4FJ4KuLcwAPbaOR8bAkNK8o
J51lX4lOfEtjyvjuwinasjvYqehTROouqGQ9BOXPGb6iJLxZc3YCOk9S7LGI26Sof5IRxtdu6Nq3
hkZ1M0z1h2HVt5oHGXXXec3MTqC6bOVCXmwkQWIYpvp4cdzf8CFyyKnPbI5rKKxadIa8afYOnmXb
9x/nLDUIQmT4MsJeVamA1xriJlZzwfjrquVesrmsUXjyYwwdHvsy0VApsYMzXXFC3kBlbe1Um/EQ
PP+QZ/UO0xnjjmy9fVQQfzsQUrF9fnzUOYIwmFypgjAVAu8uViApnr9TfPhsams8aT5seZtb7Vjg
v+FZPGrmbJsKxWjrXWBEOH1ZcbFZxGAmU3V15euZtqeGjotUByaHi18J6ks7dQ2PmNiNEbOBlasj
rUcgkBnuEZTGhrRb8WJS8foJcA+6EFNM653PYLsTXggshm8GI2cTLBNwh3vXUI9+SxIgCqUtBsrD
DMiVqKHxMRtBHavlvZyAvZ38e4Uc8flxOw8hn2HGXl//iJrPaqyS7CjjU/w+IUeEq6YKberhq6xl
dHM9q5z/Crz8dlVwV2Sq9fwL0bfmC2GTciuGi/l5f0M7C+wm6Y1G+cA2R+Lzb2w8bSdmdiNSJf84
KO/dv1MSLbZrFYi9cs8fXW3xi/N2GwY+osbFLyhOA555ZGsiOUmPbR7tyEx8UTEjv7mp4oQ8rTQc
N+42JokjYU7LmvEwLhqWrT/i25rzgj8Ap06tAA4A409xRV154upo5nfgDhnLKve9ptGKploM+ISV
iX4uqBy4PCg3ZjCRGuiq1vi7tBLWUpoJnc3m/QiK8I33Vq/OD8Sd5ZGJKlDmRKV3/OyPnzP+p5zM
YVBVT5HE1DRfrOH9cD+spmRRwWjZwQvWkT9AnMatLc/yptT+XYMiXvgnM4hX4ApHc3FLUDz5MFUZ
qzb/LZkVDabwwQqikETaAgwEz4onDdP/x3eZoePA+fNucjvVVWiRY7NYko4krAHcFTtdbWZHGxhj
LjBaZvFXiqpmxWJvR49VZ005xtywFZ3Byk2DwH8LJL1op1b9LA7C9wGwlqmpKqO+wvzqr6uKC7iC
SWywftr0GYOOKRKUCC0EflAfL+/Dh3TIGz55Y7fth44QzXTKMDal9CfO8Z6n0LWdZ4vokwPHN4Zg
oJmYGKrGtW8ggGAfvA5eE6WzdSbduL2SEZaFBOe6YU4kZe2Vn8H6NGvIzymq2HfbX/fU9DkepP+s
DuZTdfqB+LLJGxLoZfniRe63mHlQBsu1ZqQJyvoDBganRqWNmXb70LIl8reZKetiwlJO1Piwq9P4
06Gxsw0Eiw6ARU6S6iPHzGUhb3O+9JXdCVaf0umGGisAI5S1KsnbLD2oBv9x7Y5reVGOgKIqmVfM
Xk+lVg4k4h7LS8RNF/k4nJ693Ap+suYH1fgzPz43tVhzwC5Lvb5WBHhozcjq6OL4KJW5EvN49v1w
u4KrEoJATKTY50ziubK6sOFQQxr890pczIKylWtLPTz3sEGMbCTjQBALXf28VIfARLdzzPzzMjkM
5n7sQj9/m+dTdwmeqq9jvO0oQ/5J6XhyudfPby9jWnwwQz4hlPIY3XcUteEivXByiGiHTb8IBDMK
6WQdDRXDLkXA9zkV+jqm3A8EEZ5sfzsgvCetWkUjtNBaHzqHNluby27YaBsMgwr6ia98qTikK23O
8e/qs9aw/oBJ6jKiO+PxA0TF2BQXJoZK4N8XrGPtiPHSrpg2WbWKSwPndh2lpsnKAmCp5QZ7wv4U
mJVWpvj8IIIEPK8GFuXH87SC8088lc6mTQa9cqar7S41iEQgdvyq+udA+wOf+VC/IgnyFi3y5UNM
tkJ12ISYS9/BTPwOycnoxHl6de8C/H2iOCdrp6wvlOCZ8e8BZnWYhZeZ39gSs9MD24oCbuWlWjc2
Hn6V0g0E/dkYIKq8SlfwsX+t18iky/78Z8ANrivEebPmDYwVa+7NFrRTVHzE4izlWVUKGrUDJlVT
zhn+/N8bZky0z882ony16B1h074ZRuyh6qwBvGveMNS8vP2+mr0YSjkL0TftlRhCcZiLBaFpWhtH
sVOuHkUNnr3E0QrRxxFMt5amCSQs8heSdjiKi+LcwIhlq2FHLAZ3Z5rdI1+sbaVDYF7bBcvAch2s
AGNuDAsw0iQNuRwgRbrcgA+S1S3mMcsUkw1lBE1T1dQBUJ7WRh3MPydOaCOkV6/QLBL0BwK7G/vP
eHsDqeGvHXPfveeQKzg0Gkhs2Dc2Uvudx1KKLKs6NcJPFzBWsdnq4qoCHre0+zmqDJya+qqUcDSJ
G/0YuFklSyquvtPz1Xs5wDnwxw0uJYJoRR4trwZGUYZ/3+DKhliNJZlZA4vjnVMmP1g5VUniRKU/
1i7krfjDbsl0FekUIcM8jR3k+JSvX1MknTu3VoRpvoE28aJW66k55XtyQH+ETh6MY7IODnJXiSd4
LCocAjv7C680I5OnzTAh
`pragma protect end_protected

// 
