`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cpmLTnckjJLm/GJhnEEySb5724
XCmSymMTLlXyajuUkv+nefl4yXy9x2yAhXfBlAkKJiYo+BnqQEh1UNkLqYAA87d8AoAB9ihUb8s1
IgM+IoyPR9o3uY+NiwUbJmA8+WWguyhwiuI5cBoSnntNWESoTGk94tPn9TbimmCK7vJ2fB8ppcY0
dzN/XzQx6rnja2k1n9Vpi5cSISAq+208kK6K/eOIeE3s7kpYpnZ1FcABWMhBsWlFy9vQNq77DLCH
vQRdlhs5loIwnFeoq5kU27voNphrYWoJPQfnGHOC5JAsZL5YuLlDup8nz6nz+7pEqb8bwZ0ur4X+
w7g6QJhTOPgcm76+LLV0hFe9+d3V2U/P3bFYm0AKGrCnC4ZngWP/tPINKCm+Hi6yQe1Kg2jyAWbu
oe+9paqULpY5oDPvW1MiDLe99cGM4nW3sIULfb01y0s09/4HRnQ/2AhXlvWrYAQXOoZPk0hk72/x
NfFfhB/WPoXEynoEUYsl0+cjzeFydbR6Rw3SJHVqWdVKbmDZNvoP315WrxImh2RSUJWoZX850M8w
8oSC8vpwoIv6t0hh1SE3+5ZQacq35OmqxEVBvQIegarYklD2y3KvwwZ4yH0OgEmet9wXD0Ip2/mA
TB5RgvUIruKP9mOZaHMqzE8fVMTrFyqwcF8HDfi3LcaQHt5t8DxIaWlSJqpmbIpxsFaS+leE+iNI
3zKSdwRMTfVaIkzU9kFuHAevd52ltWI3sXHw4SoZTNvwaQ44YPlJpgglTdcQWdMNPz9bkYw1rITq
rmGYGEffErgKrja3uE2dl7q3AtRMZu0EuirR7wAzbxSEQxsvxKIZkaWDaarRh/O0XnU6guQHkQnd
L+eT5Fzun28RPXvchbt2A9hMU/es+NNoEGNFRMK2tYot8/kQQSpFbXRI/t9W/iH33vBrF7PAOJaw
5QmZWQCLeWXfgWzBsiEnFtYQc3+76K5mMbyRKFHyJ35Grsa31BMK/1+Ynm/s3UcSELxHrE8P3kIv
U2fH0FkRbliE7RJQX4Bp862xf8PHngOVPJv7Kn3dem6eEOjfpXzJ6TxrJwYQvw7Kohu1778Qjkgd
2pplJVTSEkApvWJNRqrTRySltvokG35Fr6VGurE3jHJZZn6tzyaaJgT8aUtqFaktiaTgXLNJz0ex
oiEvegnvWs+6/AzjIBG97qQLP+CUvRLILiuMZ7rLCLXC4ePOZno6MP9ahw/pwhJNdO7b9XaXxQNL
UOiDePwJgs/qvk1Rh2JIZCarbKfH8sPUPJXpuiwfTImS+PSGRl30IBdc5/WZpi5Sl28CrZulSWtN
v30oOPI/yUKvkp9pex4tphx9Mn3nEx1+XTUlifxXF1ZSxkQDaR1L7ECxgFL8qrSS5yGBWg8u2HZ4
Rs05iDojL7mVidGBsOLUmdLNvSGon61H6SsSoeAI6KcspDnjb7LPBm8BKevbD+ALKfYeGGd6k3qV
Di0TfcltPiJjvOd3aqANVnu43BROGD2cSmgGG48YVFR3en61navSEKQGl2Oii28deIx5WDBuvr7i
+uj2Q8+mDlnXd9Fc0daGwD+vMQwpk1T83vA+dFoXIyBTh+li3/VCbbqF/TP5tMQPgbT6brtVHfO0
uo7wb9vtUfrm8mjmQfRzaz3iZWtQZ6s0la6jmsSc/B37qkuVWbc2gL3vs4A2ighG7Wdys1UcarIb
kDUSdb0bymooYT8OPHgLhITzvxniLVt9ZZBQ9bd5UvJcmsC4KVkXaHAQgQCzGY6Ksg38bs+ozapJ
hNI79hmigs2kTlj9ScqXu0BbuIu5F2IoZ+7ON0M7LIx03sdc285PzuG0gHfS50IHbJO9w+xqaFWt
VfeTGBSDL+ssdXE8rXL/tqTrx+bVpwcCtU0eN2T0TRE3kt7KyqfaQOWhgg3H6TN4QL38aU5ZyM7Z
UUnJZlJNcfZKEUHrXyAaIB/Z7Q5EmRqx0HH0Z9ZlHE+4r5/nTenCB0GJ7uBwSHJVCkej2cFWu5eT
QzDN7TONsAXa02/mCO0BRV3vWQkfu5+Jnto4qa84OjAG2dRO5CLis0VgTGF04MhQERw4AYKp5h/B
dq46dsZwvfr9KlxaDNdaCrJBVWrArQ/qtjQUfN2uJsckUJwo1dn1Yo1dl9koP46b6QgtY1phIO+/
Dgfz7Ng/hrKzqQ5l1+6viANmceOHqpwC2FnSBGnuY+Nd+LjMMAkVwx3YCU8CnGBm9hPa78fAdQ7M
YX1WVxtTHrJf1RP7bYkmv3ga10ZZakUnf6zJK6GSr3mr9KFi7uLL+w/uG85iZm64VkSlStyQQMIa
g2iWndofMiSqY5m0ghkM0S9SGhfx5TPRhSAWk3dbJKhEUaw/Fl+qJJvZe2fckdQNkre6NU2yoyIr
5JeeqfU8t9QrU9yW0RCptzhx+J+CvFynkKAuxmLGS9Vfn73qTv7NpwtqbTk1dVggxI9Qo0v7US7c
iLVxUOdDkb5RHxVCnocx4McAHhvkpj3ZJOAiX5TzHS4p83mE2UW8KOrPKhJUzFFg17oLkMTYE/Y0
vz8bv434hTp9YsUHQee6af1QtaRnVIxSin60nFWxYQlxc4Db8Mxxzf07ZzWr2vTfOvWmdXBmSwqG
wkHZIMRzR9eWF1gWTmFY/lQdTZPGSOncPILLKo3i9Zx9bLFhIee89wSOuuncHG90IPi7aMiJeE+V
SgTbkjzQHoVUrMoGMpYzITJeOyz5kTQl2letbxzQluJsMrXpiCr75SbFTDFHJT7OcTtJ7MjWA9nu
0RdImcDIh8QDZgNudREoMZ/eSmSHTuG73llDYSmt/PzLZ5sRLMN5pcDpsfXss4pXZQvMOUAkorxx
yFDx0PIxq/w49AInde/fkl36lttencyLlISV13qzamPhLNjJkdgupnqhCy+MB2fbWBISGdDu36pP
CGfoHMlcRgCSlf1vINGhhUuO523uszIqFUDjroMVAzmXXLtBicFnPZMFnxXY5xt9/lyVXxyOBWTC
ewvJWPocb17j0was9sqhUy7F2PGxyAtQ1iz0uJmKBeEHGTarwOKg/TyBRL38jsEsbDVcQvzEVvLh
eKYV9DYeBeJc2JD16RUyoo6V2F3+SO8dbwBG1dSMpQpaPiISfT/Ac/dsOERDcFS/aOYa2u0QCEV+
v0I8MnckHrS7r2ZTlFDj9+JXVWOXe7GhpzKbEhNZ0/nW+brmQzVxcV7/0tMdEqRnAF3ABdOIH4yt
Lz/JAYZoO4M5dumtNk4ivn9husse5WFnVfEKWJmOpXYB7Qf/8aCYh9ohHLHERxMmfeUQKSo5BzlW
qmS877Jg/nzQEWUxiOdj8G4Ky/hHkpuzVp1VYy5dL/WgDFe4X8/oiYFwybZKXfbmafcYappagWpo
7/Xjo2/Dmm/itqSe0DvTya9aSgFW+E/5iehFt0G3HcBS9NuBircqGmL153iNwbQTRMfuDmtc94gF
e4bMnRzhx0KDhq3+UrmpyKJLAyiSB6JwJ5ugD7stifOIKnMsJN4cHjUL5HuOnVx94ZgZZiKFN65j
B4uubOCTDFL02p/uZEgglEfhPzPGDombE1itMUNFpyXqIH18xtyKfuBOiDOqwkVZA1k4QoERoZK+
hPu9upGI1sABR90ihpUBpDunc5ho4HvsU8+i7zdON8Mgo3PPWWJ5CYDTf751l0kl2IfUr9K0l/2q
4u36U7W66yNo+Mlj54FTBzhhywohJPMwFCEMHDW4qgAVBb5dyBc6HzUhqmDmbHSeAW0IX8LJGeHh
/+pkTv8QxoGJdW7Rz+1gIGQETkJjUIc1DEoRMBk4bvHjriEQiBBMJvdCuYcBkKcXwGGHBIqbh/HR
Y0uCgrYPBNbMlHUXALgBBSKXh/BRb4raQpqFYKL32tdMnb+8a+MGv3BVrvJ82xlSOIC+RiEMMH4M
osDrbznYjuHCIDwIaBhPEvftZrliQnVquHQRDYvRBYcXZSfHS0j3ic/v6+VFqZlGLxL74cVJCuEt
GIZU/vs1Lp5VShphhajnUS72SSbsNFxVVaVUQxqxNyWbEm/SxsEMJAU1cTCVWBajBiLh45fpFt+l
+N0oXsPiwq9tDZpgvU7MeteHc/uTDm2D1hPSEz8Hx/jx43B2w0hXFTWX4mpqmVFMyIo+toyhXhi+
fOmN3UTzYtZF0sMIRVWLdvu6Lk8Aq1q8CTiUmma7XkHEtwFEKIH77QGpHpBA8jaay62KTEc5pUvH
dgdx+6ZLL7/IAWOiNI8ZPi1Hx7acZsM1HU1yLpGElKBd4n1qrGhR2w0jCpYlwtKSky7wSmKscACg
dio2DZa+vexphrsqZrbrhUNZBXFG1Kw+fAt07exMCsKyxgvOjI2+lP6Qah6Tsy6SckQ1FOw5jL9a
6JgwTPBhfbJ9AHagCaXFFOLZt9KuYSXrYDe4pMtYCWOMAzXArtDbIhxDohtd8TT3cGiC4CokVcOm
mq5MxSsAHqu4RXZbDvnfKO3mRMPdGkvVHHZ7422pwJ6MDokpUesugSpxogwgql70AwHjkRWyZ89l
6ty3Cn/mlJQYlq2oyF3yekE7mgCT+TzBkHP0oL4myfWgxI4QNczB9CzLW2FFPb0Fd6cuZwdN6Zuz
LeKaDVBKfk9nvPdwbZ9+EtGXXKyhR6G/QtHxNXXmWCqxxcSyAUKbUnnSV2u/xZpUtqpJoEevH7Rw
fPgpMiLcVYiRXxEhKKScZf3kK5yEzt8DU2bOvE0qZjbFtjNvz3ceU2Z8QnloXdvPkBmIsuEsOGQ4
urXA1AdIcKxHaSWuqbMoXDuvNbCmrnyAq2T3GqWk0hzwPyJwRjeUDNdQFZkgUpb1zPbyeNmRL2LV
8aFr+Udad+yrPDewnkHnd5MdqHlbgjAurKMFju4aO3poYxr3cBjm627eS2h3T2tdsTSntEuiJjwr
dFmZKlS2I+cvGMEAkeC5TaXvsAQDVly852GWJ+UgXMUnwwfqyg8rvJQgfqQ0G5nd/Q377M4NDD4g
ko4FVfdrc8Ws9lVqF/tSl76fud/n5TzQfV8n9egFblrsBX9t8Rk7uoEwVAMEJMSrnWL30165nzYs
JBnE9f0g+Czgiavsf6K1+j4g1AMR+qkcrdyeuCsRJbjOmOn6w67jt8IpVVebWLUJJJbFbW9k8/Hs
lw6lU91IEzClxRVAkPYvWq/CAAb9rbrDV3oS+lsCRLBxmjLLLOF6eJSvp8nOT0EZBS3wXexV7Tao
YNvCiIT+ZqamNdMKsHpuBNX9l8gtENd9VV01WBwB0nv92KWPX6UPXOADnw94LUfErBCRaHQlPo93
oV6l2fb1NzFOhermODiBJKImAPSDzxvhmp5TWxiSH8oOc+hMQNigbzoJTm6VnoOljcqyHa/yblHo
CouzcE9YfE/2UWyU80vYqwTENco5wFekBU3M7oUnehqe1rti4bcrhNRAPcPbz6s2E6SrauavSj/H
Ndohhmmt3IQSlIuUS4OY6TMQaI72BKOE5w4pirNUzTE/jQmdR+oMXX4WvsnOF3i4IYePwxp8OCvr
LwrHmhDMOWb42BX8e21WJKdxYhReooJC9D0PW9e29lh/FTdHgIiXIJyJbx2yyklV9eUuEernN0ZB
YLz515xCmzLibVtjpvwMb4OYHQ9D3L2hdrzJ1VE0le0YaJON8NUJ5l+bD/Yf/f6YRQ2sQL/GEehZ
NILAbVWvrZkw+MFqZxWNNlztjAkKF9ugwwbNXwVN/hqTvhcbA7z6hAbLUsYDZBpRESAGTmBITLlk
AArPO9ybE1ZTfjW4cwyfJ8I+WzsxoFMc9mabpBnlqffftEMWnSXpVJ5yCSEFD2mgl5uQZ42q5iVr
yy0qd6dTEi/uMnPqTzrzE+jqZRCG7iSv6pAdsC3fAwBMIjwmNgsiENLGfvsf/36VgWDZvFpYGuRq
iUf9YLxWEHPcWyNpuS0SGUrNBEfQYFUM4Edi7gugEUnv3J0DFTZ21TTaMIINhPo8FMobDWGdN+od
qvaG0Krim5Xv5E6L3mAsKcUEVIkkem/UWMOiT6Uf+9bndix+WsFgxunLJFmgCuKIL3xeMy/xoxEY
4+xdb0IKC7l94xFgvTWgsMh9EgsxrKWzgwjSCJWfVWBb5z2NvN6WpVGSbIAkKHR1KB0Z69Rais8x
eKkX4/aT4Nc9ztRk+xch6JPSloOTgJiZg/qu+tAErSDnWgOQc9CFBXCsWZ0DCDXf6gLWJm7H76OU
w6NJgiyCSdgumwVw7pga/auI6xNVyppa7Sixjnd/kYzHDd4ZHLrJetlFeC6SV6TFJ172/3yAzWx4
BL7q7AwsSEnng+EREGH4yTt+1Oa1CANEDHYx8AR9XXUrObXe9zbEdCyjhnZVNNG+9Q0xlG3rsPm+
uHer887v0Ps8alceuMKneIr+de5d9rXFvJ+/SSOzYfZhqWGkm3dHVcG+hRidZi9r82g2EilDSvaz
8B50gl1sMBVK6Rc1/QthmYtg80sGlpuipDJuZiINO0q7Gj6CObKLDnRXtRg4d1q23SBEOqI5RjlI
q6Oq4/FwhMOGR2WCfLoM7f7TQsO5jo9FyWQ0Pb+TICklz1t1/2TiDU+pUWU3XEhfx24bb1TnqJ9l
M9Uss1PJlEtMHxN44XaZhVUMdGHeeMmE3fOS4yM5GZJpNA1Eg9BzepioMOyjlxSToe50hxtPyKMK
R/JFPbxREZtKkwNWJmG268jNmg+5JTiIc0ugOhlvbMAzTCfiaVf9HUw5T5nt0/Nx6f571heP+lSA
cDtgPsFyqp2bm8ygSV4n2D0F29yKN5Upre7eQpWqsiJL+ACqQVi9JQbRvzh2WbqBkbGFJGzi5zN4
OMA3TKQbHBX97f37yyL+/vUFPLY3MblJqzlj/86nwPnFn1Sa9WPavPXkT059d6CZb1Thstk+ysCn
Ankhbup3C2utqpynUhs6JN1OrxTh360jSwsHVfxkPOfSzk7qxpkbXGLw1pS6NU3cn32MqFpbssiz
1GSpSasSrVBZrOyJBY/nYlr9begL3XTFlIMtgu8ywfHCSkX+6rBjnrxtyy77Wxb+1eBEFMHXk3ED
N7yBeilZCqC3WHxIu3cWTWdVKTrOqPHF1b5NKop8ftQ71zsY/Th4EbK0QC8HmNxzZwNG9S7OYdWP
ZwiJwwHsoTPylZTxqEPfFF3XfugDWPwEZi8DLXQAadjzIR+w6JKThqGa54T0MvBuP0Qa3WXUBqho
iqwaCzSwnLovuiE7dll7/6ZlLTl4j7z9c0Q0jox5irYjbXy+YQqMYcTis6HXeMcMubUdoK3uCbgI
kSMZ8tnhypIRlzi4bil+f5WPtaOrxoqd/XRMIbryTt3pXjx8VAbHUH+1J7BR31suJ1CD16C10er/
XFhmt3RU2t9eLxgF1Vf3PgY0tijLmtgYRzT1I7uviOX6TXXU8ukx+RhO1npeNrptMD2yV/Tws0RQ
g5nMmrGhkSEZ3syLU6yQhLgKAPjEGqa9AMsAVaF+iZ/TMZwkTR2akMrTb6A53oCLVYdu9qF+dJqK
1LtBN8SXe4BP6/9zK4OEOaHpBg0elz6GJtfx77SGPDRfa9lD/G7qtKw/lJk2r3bxvJrZbsOZ4X9S
KuPkh4r3E5lZPkNBUP/EtkjqHlZYDhmDLZhS2imYQVrjNkxe0Kk0YctPIUlIyGf1zeTOXuAfRpqV
dsgUMuk961nTGoDR9Ir8JgTw2NyPeHkpPM+eg5cq2nDe/kr32uzKB+vSq0mwhRboUiP992nK1RQ9
uVhN4YfiVkdBDSk4lf7foXtHt58fXWGw83TRwUrM5B9Mt0AewgrW1QoIYALzo+6mDPcFIotTIWkX
5MJf0oRdaUm8LvewxhVR72fi789xwARvBzcvdl0ZvBdNbXzwYLcZY0+Ivf4UC/kRKVysOTyfymd3
hNcR+Zy07Ze9sfCVY2TufzhrS5yKzmHkSDJL0+iA5JXgWGDauEvpYqNRHPxGj4b4GOTuCtN6hjca
Irl+t3WqgI48GNESsbbhr3yNdDkQUB90HDKhGMEaviWanjPFFc+UxmdkceYX3OJSI5Cw6Mwg5mUM
aGddN4MjloW6HGgAdebenn5/xfDKFJ4KNnBIg4tw6iDFyfaMZg7UBzlNnz6zXI6E2v/mqdx/QWrl
0dEywEOkWskD1HBpkCEw+lfQd/5REZ8BfGCV6Zu+HNXrbEK9+2ynrcj0MCQ31Fkc0MptMs8ZY0dC
h0sXUd+7Rbz4cKI98NCZuWNPxjMf0HrO6B4U/qFosBcAwnV1hT791sKXY/YRrNQUW9uOvi/W7U94
TIlziaJDLmCGcZboYVAzARDBNr4piXEYILTd5XdOanmMlpTaxdDQhXJieOrz3+TBifcetgXyFeMo
audICsBisa13iOaEmJC4rgS9WeV1ApCfc+Yj4frmkG5KQ8A6VKRe9/2kQSf3bGT645tuwdPNU8Am
BQdWpt/OTvJAMq5v7f7KtolsuGPKabk2t0SYNLdEbxs+1ANva7yd1ooejzp3AuU6W+Qg8B4tyJir
hbV1f6/t5zzfm7YaXp7rLZjqm+XLch89KNhCYfIBTC55gMsXiw09tWlROe/jyhaR+s5jiERZmb0o
XfqUXggtAj2r+74spsPVh9GrOCz5goYJC0odkBdaTOQy/EsUpag8obdzPwP3TH3KnjTlTaDPUzLD
zQ4S7KQYnUAAXCR+gnrpLpMnx1xR/jVSAPflajWzlCiQBQerrsutm2SeoBksZoNZQ6fqXE4xPAGB
NUCfcAzIkhej8yVrmPMO4AuBWwvKsWGVW42729tRx0T+g7XrnhvIFC7GKhhBzTUrSMIjYA3CQ/jJ
nrV8YFMzNaV5oFKRn+MSU7MjbihP8pmb419gnvAzzngyooaSB1USmPyfXhdUgqX4qkKQZWYLmAT/
2et6G5zc7O0BjITP4jhvr4WAFQ40+si2Z3LEcGRYmFYtHdBTDLRBAOo/E2JCrrZcjba1GUUGuWDq
8n1fQS+35Hc5TcqoV3On+qAN/N+grmxwMv5vuXOdJ0n5hEU89QzoyuP52bHDQdTtdjBqaZvvlKSN
bNrSRRXhcFMHZzAoLNHGw33WY5Hk36MezG+JM7UZsJofVypUjmtake8JO12HVD/H7o6oef2stNEG
sNAPxDy5pX3Iny40sxfA11p+Wb5BQPPSXmdyIWaYgcJOcu/9rkK0FKKEsCrpHdEDzwh/8hgBfqTE
4UL4vbojlgfjAkzMveWnFCQO36R0OS0IRjwLLgjNZOy7ufuT8UpZxfZGI/2GM1CZf8JsJCLzArKg
xgr9+0jm0FvjGzTPQ1VALCPvMdfsbpmRfCxYBwcZz6t+WsWjhVFXrrQXLdzyWuAvxUFI0dUDwsL/
2VUSsMDzS/FDg0i443tscCFaSYwSdyhwvyouDABLXz5D9Wk4gd6K6sPjeFai1B980eCW2wBelZbp
omjEJB2nVHEOwwE1ifyiZ6f6jEizIJ7IVqO+Dp00ksmQIs4Wvo1Ec4JrPSot7a2VjQPsVkt8Rmva
F+teAsHpEtf6zjpzpB+lyh99PW5IVf0xrsSWxMDmkyH+obpVYBft+NJTV+/GHYoEtTFXTsL4SIz2
mbieT7lb/d1wQO+BxUP4KHdShiOnf5vUOE0kBBTlIEx4oh2NJaW8U2jqFAr2r2yDnoUYiwB8jYBI
c5T78v2MRP1zporNeYi1T6k23PQQn0hmnE2jtui0Joc5Ne/yvY8rwiR717cGE0YgJhl3oK7/YTbq
bbEOIMtf1KbMS6k6impcl8sUR5KPX5+debYUrEdjFAIw1OwWEiQYE8mm8dWR6wLpekmSbhFcD+9a
w2iePNbmV0+p/4tVQr/snNMqKPG2dgW5bjYuzNigNQYaMGnHUG3M95zZMW/+YNGrgLkk2V4aclBk
H+hIpFVI9vJ2LZx6nJOkuYF4ywvEp3igad2vgXgJCrK2lcuUZ3jg93jTfxwIrPT3MYRJXC8ILGYb
+17pp5TC1RgTcqhJBF5E6IpGfaB75QCcAup9HO/Wmts+jOlwCaBAu2YG88ntk9sb96lr9gNB9oVr
hFxZN1RW+bj7aKNnT+oceQ3JXF/2CFLgoIk3C4PHABRm5BBFmSs5qe4txXN59qt+xkC+LsBtiQ9A
URrPJQQHbkd0M44MG0T6HPVFU+nnoRkQjsuo2JEZdR+Eoi2HJv3V3S2NrvQ8jcSg2ng/q3lpiD+Y
uf1UaPLGACk2DzypYD+hMRdW3NBsEHx98ICxLv/kQDYAyQtCdyWRsvZRCdMvDxx6d3pXt2N++u03
0m90lfb0Gf1dL9pz9P+R63cDWVgwFC+jQZgnxkAcbwDm9uEB9Wzu+qc2B8hxt5AphH3H6iDHd1/A
fio2eeZyFfjRdEVS5naLC2ihRouHeL0nlzJoi8xMa4NphwYuh2iGFl38Mq8J01iJxImCn4Wze5pf
08PtxQm5wn7KeId3kCdi++o+iTKM0VesNH2txswmTV5D97oSrBG44bj2L81VFJJvn084gM4eGhp8
MN3fYHwSeZVu7takcsTO1La1144IGQOSZbe/IWyYWv7cp8TXUbec7iVv2UH6JlzL7HjPnFcy4kEr
FnDtk/iQeuh9hyQbxajSv1j7fGg1ZQ6w1PAXP5gsS9oaaTkiW+q7M+ngxJGYDZNlAfLIeUnPMtUl
qItoHuGcH9Wa6DrT7J7nLUsc2m2iq0+jvHwNFE6oJeQy351YpCzFmHsdQuVpk2yV5dS2tye/VdSN
FJxZkkg/uq6RZk34QyCPIa/MZicKVSy/2Dk4R95cEeMoxTPgH+Cwj3YtB3986U9d4tNCaPzS6A6N
BDDjUf3l45N4AUZYhgn0ZftXxbVCvNLzN6kls9JOPBuOh5qbyjjW1Q0IWH3fPAyLjSyuVfTX4xD1
A0wKd0tSpUac52/YMEpZh7oCC/tEuJIGTg5a81L5DQtwPKkqSSxNGiUZHevXJQ00uKQ9hawfUJjR
s5DnOjstWD3SbxI/XvWo2mNTmMByOQmqbaA8Ttu6cu4OHUyabfYCp5XAllzLHrDOVsMahvyWYq+L
sloHu92SZdZFe/ssMuf7A47KGeETofnxRRkMgKfqGOoOtdA/mUKcC+PvAsbblFVzWaiZH6SDprPm
2nu6Ym6F/s/JhK7gHDjiuVJNHHD29K5XYxIuTzEM8aeSaCQ/o7NNkEkf7YuNTMlNiJLMhbJlaw8U
Wdox/GHLRZqqAFbP+/L6/sgFb46UaH4/X2wZ2yZot+ZbP9OtOV2G7kWzY1i8wXDnT9OWBVAhQmy5
N+APz/BWJGIrqqAcgdV8OhUP3hw90unUHgq59RSbDmWB9zNiXbajJxRUTQ59Se5tUjnqraAynsvb
1jldXRYD3XMmEWLKx+a72aeawl8Qx1zn4pGLA8adCcyH+ndFuKkmHW2pEpABQwRfUVV+2v/ZBeeS
dKfuWbMroVNVN4OeX0zvKp5L+pxDj3/ECrTmTxk1lLoFdCPxeHb1djJcmIucp8NoYZVM6o+N9OQe
H2gg3UzcFwNKaAtgPbebdVG28uQujzgT4XIKCI34Fg3iBB3vIWoqPyTKWqTJRfQjDQYUXk4P5rbn
+6Oa2Fb6SaHlahyLLLHAw9oFjiaO5xMz39YrM8A9IilpnoFUZSO62C1A+slBAvYRMqlHe+5yXaJo
ZyR8a8pgCMG6d06t8XuSFmnrS7scPu/RXqU7TQUYa4W8HYKWxIG5yZUrQ/cTC95vCDnUXQTCf6eS
XXq45zSzAR4HgcuULLpsZNMNNEHNIbVNRlCa/hJEarOCJ6riuWfsf3f2Nvgn4J1vInF+hCdoA8ZI
uMUCMed0ogNHpn2fPx5eHSuUbiG7VCuasKfFI3zzHuwbuyeD1jS3DK39V37uMDDxWULZDxRpVoNC
vB/UhVumllcmD51hO/kJgRo8sjM/ek/0/14WnzsOlSOicSr4rXwHqly+PgFeeYdSxu/LIYr+59rX
s4x6qLiR22D52o9P+xSnv2iFHjrTbaP6wi6wCL8NpLznK5uF7F9hVAa/yidPTFjPga9FLM+NBbd8
2ydWaSJ2CHFOYzBJZQSuIo77gfYwhgtdXDow21I8FOZcDkDXROKYRkYaMjg+u0JML+/2nDwNKO3Q
1DcutivXJi8x+PmvMAZwPXMP/+XTON2b1TyPPuaYaThPmiX7DUvwuvWkUrBZdLQRh0WESeu5/s+2
wjGua+4zb/5mzaumrmJeyi3CQuHZr0g2r/9lgtH5cAr9LgBGg+TuOAmCmddNJCyS8ttSpbENwUHL
y4j6lyjDuJwXV7wjpo5yaQ8/pBdYN0xbIsb5Odf3zNLf4J03JIIGVwKptL6CsH8QBOv87NJ/2W0P
YlPUfMhoVDCVVKa1P3b9sVaJ4vYyr6bNorSJ296zDmJtEa4lygL9mZ3J8LEpcemWWp7WS+ZutRY+
j3L5YWhNN8CzOzj1cF7L1m8JBYMnF1ES+Enfly0Xf6zJnTsST6Ey4vR+uWdbbtr7XjEYSVK/7TW3
koUUrgbYZFlurPyLQwfUDV3VXVu/4+Tw/47C29AI01nj/MxBiW8tKEuz4Xrt+WcnvHlNpui9xmSl
rvsOvLXJEFrmRAOi4LCNnU/iPWkh4YgfDNMv1Zs4EgQo1A4PBu2EH3gNkpCdE6CoURk/p+eYaaVf
Z7+M4WVr9vkxC1f2UvOseyuo6q43tQ8vf6lQNENBCNHZDZFBOUrxBdFN6PnDfbH8kEiEtRGUS+KO
EoUQfJd/UwqYueDIZo24yl/2UMl3nnv5Lg4CXeUGR/hpcIVznvgcE2j3hr6Bvru1xgCStXpULFMq
ua529cxGNzrYq9b0/gKjDCznnul3+6uOY0aOfBUC5ohHri+XCzSJJ+cMZarkup/bkF/Pi7+bCbW+
/o8MIvF7rnyeY9ACH6wTFfNNXKf+7JfywvwKoqilv8inqoPFPDqSJ8h4eXnVdgSm9NaomxBAkIk/
gENtR62Qj3uTxTVmP/zIVtZNRqiKnWu2j36TjchoJkiyZ/EczR8WBVW78WBIEnpqhiqnw4JZlX9Y
LLenOg5ABmu85CdGNSPDUH4CqDTYAfPwtIwXDLT891CbCNhLZukVyZFJ7hFwVwwc8XOa69HIVINI
3KuxW9/Y6f4HcajvNHyPSd/g9dbsZnur+RRbVwQ1o62LXkMViVhQRvBcAr03GlFthWkaoStH0deL
NFrZIuN/TcF92p6d78gOQp+nwY8VT/3bhyyw5LPWpTmlqbbYyolRKJZAjiBWwt06879scGPGphpK
bp3n9YfoDrgW/Wj3GexpViqbDvcv2XQaZDKdk6UGPBniAip+9wPLb0ooQqA/kz1Ehj2at89L2cf8
H2INqD1st8w7y/sCzZDi5iwot0lwe83omFQmOZTSxKaR3zjmQ8RF1wFc+PSPsZ4d/3gCKt6mx1Wr
HsCpdOG8tyov3GMStVpozL5GdW639tUe/JoWhxygyXGT5XzIZyLdoNvwcvlUSgc7BqFB9zgBstb4
2qxPnJVq5iUWmmnYJwe3MD7E8/WymiXS2DSfiv2RtVp6cmAMV7zzYvoHvg0OllU7MZpj5C7SW9tv
4OAjz5rwwza8PeKqABMzy7F+8cFwLIYeeVSlnYBk67pofh6xcf1ZzxToDzxJQ7fppZN2cYegyi/r
UTwxSFsM5196JY6Kw/yqMtSomP7Qq8Fpcf6JRbJRck02AEBn0lBhnuLIfOuH36Tcem2ifpMTsCfd
q46qwoAEC+ncqUioAh0T2aTD0X7PpS9Y97nrEp4OLMIK71eTLTo6jMxWRLVpKTH+LDLswnvjQMqh
afVdKuBWog2Lc9S1MSDMymWn21kWYzQvMtvZIbuYC/uEeYHQ0M3MrgqwooaLVGpNY+jCiDlBZL7Z
CVF6HoiA/aONy54x8tYXAVyLDicP50JNISndT8qm6olxY2UibCylFeLhMS4Yml+Bb0UmEoXadbeX
k9W3w++JPuIgGGA0oQFBtHnUhTpsGpCryYgoidlZ6pwMqMfLifuC62QvRR8M28y6Rcv1YkDAE3d6
d2KAh3YziTLJwnxAITH+B46XNgb2tms7y6dZefS8d6MUQHpbahrtYQT4ogvTCrHjo1RvO+59ZO3r
ff4Flg1oW1lNOCMjOyyV/9XoeuU0RhSWP2vdOHpKNUmqtN8Ae+/KNNz7cNWPH2uIbjianHoEYiJ/
3qYFfC9Sg5fDZ9gieLEHEAtpwLL57BnSXm7FjU+Az/+P1vEi+MU7W5poe/7tW/ciz1ty79Qjed5k
yyghoLtFIWWiQ+993n5VbWQd1WsGmipIhMM+n/IBNVFnCCSiU/2AeYJ0P1x8kLbl1XshIJ/RpzRA
NYeshG7dCpI4cqH/pXdPWHDqzIraBMpLB6kp5HgmLGLfiR8dbKaOfh+IS1yDQ/hCmZeTE8cKlKOV
+zm3wossX2Y2iXSyO6WGNTDGiDEVOH096c6qPEkqaxflLecCeuk+u2Hw6zNv92x+E8T2V6VSYANt
m7YiISnzerpXGMDF19BQzOaGFAlPnjHM1iyXNEw9VMGPkXx1LpuGOAOYONq8T+1Zn3452+f6gqYV
TlRxJEFann5nRDr1G5krYC6gXZ7/HRrc+z3QqMffk8Z6PMQZZ7l/kTWajSgTXiesAnYPDtm593v9
duN0pEl31IMJew8GsbYwpQh1GFniZ1raZeUrPslvlouMwVQNV4qZgtoeh8zNDQtS5Ro45VLoBRKm
I9tKfb3glYD7Hx1iHhPIM7exwyndOx2ITQmTp/uX435okmImx8ncRmoZRIYJc1fD1xxhvrAiQjnk
FU74huAykcsrA62Bh2iJLCfJCR71q3eKIqIFbvaHiHPNLq6lSuOuStkMS+E4Fl1fEpMprbFZGqJf
/GKM8Yrx39z7NaWHgi6cjQ7Vouv/R5LjifO/DD2ziuNK59QRogVDshi+OoMQSMm/jYDoHcJawNZ1
bStIpzeC5rNjPV0GxENrSnTR2bSU1tTSu8fMOwVvIC1eN0LmzeOWv/Iz4Pt4yRPtc5T1YNVzuXqc
dq1ePMqWrct+zBJ92M97iRaYi4eyZKVLM3Wl/1YfliMI77i5cfsfDmHt2qav+GhQzeviR/I5XRhb
pD6AYgpituH/i5nPmIJ+a+dYt1PWaJQofz7Wc9w34Wb9Aawr67oRVJufhxKmrVA91gAhTk/jvc2i
GKA+mRuDAYrgwVy6Cebhf9ni+PWbZZCPvd9x8mE/lE8ZkugJaM52HbVp3lGUS6rRKI/PlFGmhpJe
ojOHJVdo6Y+SivrOypCeZG30XO/cntQPNHZs9TM+fDZfo2xyipiiss0t97Y1X3vBs0srRRUJfwrN
aeJYQMpxVveUZZHStz6NMPtgQ/C0ENcD61R5VJC4uOTTG0eIdcTkonWSouQU0No35X07K0S55zpL
0j/6+3XGujBvFTv0DaZpNkVJUDFxdlbWms2FKwK2AXtfVifxdQJgSPfYGICxw3SeRjXrWvRYrPEc
JiwutfP7SUqpbMxq9MYiql9d99JrWLmCR+KB16hpb2aGosg3C17o55Ss9gG4BC1qIvBgmnBq+kIk
zmMo4nIt4fOZYcqZU0VTe/7ugRpDB2F47o2jZ6OzcbFv5zwHTDtneT0c4dJivwDtSpCHk8XHJfbQ
5fOuK01+AXXdXKzgko5RO1oL9isGB492WK/gMLCgTCTMSWkKkeXt0mZdHPPc6eBTHP3plZ+TH3gI
/xfVFDaRLph+PjUWXygu7i+upVLHD7m+GU5ln4h76KbtV08zSDVK7xnDofdlTHMWT5/p8ZwPVn7P
80jgptqjQuUiuULSiVpJ2u3DTPsb2abxNvz1+veqwyK9PZO3o8Zy7mvyyfNXL4WWTUqV3YG2sKf4
bICU6hOqgMPkGbO6hu94hWj5uWCL7FIMOD13Aq0yoaFcj/ks2xxTYaMW/TfLTKNT0CGkrCJoFWoS
i2E0/ssM1+xNI4A9Zm/bqIS7CnFI6Ninnr6+Dcn2+HuhiLL7TvAgCtxnwkU0zhK/fiul0XtgC5+X
M9xQR61opugglR1/R8Jn1BeNaqlV7VtcU8bdpGFhKNrR1iI6OAu3wsAcjhGkyckTryedpRJqXjao
HfL0kb3vWHmZqT24y8vDEGi98POHvmz6RMmcVIhPhLcBGJKFDIH+17KrmVYlbM8KEf0Pe1pli2P0
KM9NbUmghtipDZtOPNRTCgUKnZ4jhJwk2nTQTElkizJ4dmw5e04mzbCZr6nfcl+5owP7Wcmh6ory
2K/+WFt4oPt0Z/8dWXMwXNpXL79yA+IbwshCRR3yUNnETbSK6whJhsCSLF3OrmtuoeCfEPUtq4JB
zZvQ/6ppJ0ySPebcy9KYnAHm/HpjUrXdzhmmpK5brTO3B7PqV/XlPZT162m9KhLIqrvjhuQdpyyg
SqkdHf4MsQCerZ0XbaLnG034CZg+M5HItpKR9yeGLZFprNOJPQW6vU1Vi6pEggJLvuc5wooXSKOU
1zEKaZ8gXF0QAYR1/o031iXaznAKhNiYbL9Le3NfT8UvRDD472qryWRKELkOZyp7kDvRPpTrnHvu
yGXviexgPlmdI9Im/3yfi59QlYJ09Zf0kBSsSuKYRnBiqG9X9hOqCktXr6LJWx9dUtoWiyPw1QoL
c6iOakre4Qko3CFnxMd0agWW6qHLPA8JU6tJo8zZLn/c5g4of6VaXn6qT3P3xDEtDqQaXGbr+PL/
ylDvx3novOx4VRwiC/RU9yIf1ac+U+gsv2pjLfVvRCMUnABveSOZVKINYrvy1Oh+xE21NPYkk4rE
rwS1aGwE0JmSlEMyet4G1e4/6nNgs45OeHIgMoxstgHrw3BrJhj2DM5G0N729+SdeQ5fVZ4qq5JI
HPOyPRiuAWhky4im9/fR/EAz40UzjAvSxLRyTnyvo1tcvonUGQxLA8xF5gwjvFat2lOKCLnuALzt
mWqAp0lpxbWCADvl4CiQ2kIaqnBrxI7sop9NRWPFcdsXrTnYu3BUheFztoGaim+uxxm4CdgLKOR6
ALkiE8GkBmeG9ttgpI8NB+zegGxU9WI2S//45xaLQ5CD/cVFClify14kWEBR2qMP86Ikqkx+mCFz
qdSTKPC2YABkxdNF9cuAfNzRaXBqIizcybIrWrZw6cQlIHgzJQ+aItI8NZVUxGDqLfX7hcXz+qru
XIwkFmOlP3zCQioGiK9b8zsucTDHCj4B0OnQFXf00rQa6Lujf5qQOa0WK9nxA7aE2N3o9Znw5NAH
sOxN+VX8ownPi5wHS3R0G8jIX6jBeOxGFPuVb/FD0hgFHrKGhtazq9c8/UGAWsZfpcJlHV6CkS2M
Rh3q2UulU3orFLMUTZxkN1yf65R9HbzTSEvWil3kLCPBLDZLotof1227VM3dZyxCUy7pJAqirMqe
ZhO4RtNbwGmYQEW5VMXN36gh0uWdyrIjLS2lEA4Wb3n+//Ys1/4nZWun5ExisLR+Z7bKY9NTpGCg
ui8mYI0u2JbbaCVJjAcYnfFnMCqWD8FqyKn+l2ItpxBSO7TwoL0xYY76Kn/edqdqe6/zjnFJARPO
cal6Q+BCWJxog2yyjT8ralbwD1maM2zR3nVIWTU9n9gi5DXoGeHpq5liKqe61VEwsPV4BW+Lj2zZ
hrV03ByR46sSlBKaRX5sFFF4XV7eFTolLH00woLJS0+C650u4Zgi+pRUzc6s9pxR2w0urMR+oLqL
HzLu1u9uR4517UWvPUSncR/bpCDA/1YYu6PuG6IyCKfZgqCX3llFjYaPKXmP9HGg2XuYf4B+vpYy
NJw3FqGYWE/Hh1cOwLnJvYT5H5vxm3pR+YtGztzvIy4vrEUig0SKaBjQN2Gx0En8x8gLDkePRdeg
p+PlCvfkEhaQwPxL8crFeBsOk2/CVQXfcmFbHobgeu8k24rZlRCOX4X3tjFFuyPAOn9qZa9MF3jy
r5bydO0hFe84mfPd6Hv77tzElBQYOGr5bWzLpix1vCX6QwR91j9B+VoLCc2aEBGM0oX7UblkZlW8
skHUC9oBUK1op/K918firVwKhhU5WD4un7D6DcGDK42GA6IKLvHL+lq8dYKPQYGY7rSxs6XW4BCm
ysRVwx9KsDP9iTXjpRLs1rblJrqcl2SIQlDoajn81AXRkjQ/9YRTzp/zTCNvKVeyl3nPtalDP44q
0fL3Vb4/qZb2bgTE5v+x9PXItPBpkN95lm6cV0fE2PCCWPwUSApfIT4HqFvxG9oSjaM1gkfB98FU
d9M0c9Mq9UteyMKWVK2cnaFFP/K1GVdOjyU0644hqGRu+eLW2LQ7ieOI9kG6Utp9IEDXFdRLxDeh
7MjcDwiADNmOX4MfcAf+Rlc+/in84OJGxxZmkag77yllIph+3Jp0Gx/mmCcCpNnrc+BD8QpEzc/s
krYh5E7cRXyfn7lvLy4tIwh/o5sOKnYlKT8aY5JgLU787I58lUnoJ01zA9Ryym/sRejQZhTo8MRM
PHcJV1xo11cNNLVWI1y2A7oyqxjKustqEPaC9fu/UgC4bKLGO03AqloqDhDkubAEwBbHBMfGna+7
K0vbT/uTJqSuVYGN3obDqgD4cr4WADSSZfiqbgVt31uwnaV3Q08IkZo3xqeyfvn1EH/WRGpaZao3
3cnEWDspiyDsqtlyE4tlU+mt51s8CGOoSYyv8V4+GcnTishcIkSRc54cN716Sk9Gr8tqbWrYKhAy
OkrhZy4ywMi6Vw9fNtXo0/rWxLDCcgveSVMWBS+jAGndd4Ygi4LK7kvQLgexaikniXis6CiKKQES
4reQoRsLNKViTXJh5ZitbdY1PVK1u6MVRPBK3rh+yc7iATRGQi8LqNFLH1Eu2ZDIvHzMQ6JC2mgD
HOFLO4T6o6c7UQZRMR1Y+eE+kKn+pPpRAaCx+RKE2VnhqtvSpyupcwsHEmQtGF8s4hAU26NEa8eh
EqKvYYR00f5u7OLI+eNRonISzsnwY6uwz8SZ3Sgtm7HrRFB63IZ4/wc+jFVqs72/jjtDG8krFL3k
ZN++kHZ8okruZXyXU70Uf+RbCmF2deGPCo1h/62Guvzj5YnJzkvdFfCna3n0anizCE/NSo7b/VOt
Qcxoe139jErZBGw4Zcv4n2ivbz/U7dC+NeXAmZteeYxArymh7b8XSyUF5VRuvfklE7mavSqXeTGn
PGeo7xuMp+0L189IGUcOxAIXOg4SKn/iZ9C/r7s746rX59GOgrvLDmLoZ4/kE8l31xJ4vYqpunEs
YcutKCXB7Zn5/i9U1J1FDih+MhrtZqz1/tW92O+bsDXaZV0zyv2MG2DiH7EdHZE8iZPsppzbbZAs
rugbo4UlMi9b7tVpZkxmH44U1VKBkWfusUVzPROFhkLv7qPD3NLCOAq1vmjvfgqqIb59cZscZr19
5ATULOOCgkBVsaH2umHBsp54xJR9WvM6wwxcjlSWHsrs0W0QsqJZdaWO9gfYJ/MMPxBqROSzzxad
nte5GbB+hvQYSCIUXUpzVygg+aaNKddeUbhNqXAZC6TWsZc7D6OkKJIb6O1Fg6GPmqgdYYTaC0D+
TQYn0atidjPA5K2UCjxINHqz2Xa2m9XeNzsOS5Br7lRdeJ5S3keFqxl/24jLLlzXzV5OUq0sfyKH
hBZ8TPHzH+733S+ofwzbo1U9f6W4A+5KC65tVqs0BEsv+/yBGLUxmA4tdIKcVd39ufX2wlbF1eKw
lrVxFkqi83wUmzg72kAAv9AhPvMHMYZTjIzcZywHjrcXgaGXKw+25v7KlmrdPIm4dNWSCfrYiVhd
W66u6uQ01SK9BIR2hZQxr/0FlaKd1lbYD39PXQRaXPzmQ2kOrYOYJupSKZrere0S/FA1/CuCe2Ex
DiONGJ5RKJNwWcYdpKxPPK2hPYU/P4OaUGY5QuIrtFdMGnXV3MnERpxA1SQtNJtSdhCMBx4zVdqC
GCdzfg+pp9vdpDaOrXcdQwVm2ZLHUzQO8a8ZMAbysbKWtrkDpuGXE3rt/fCnFyPZU8Kj/LobjP3c
ErWh4TkzvTfWimvJXqH8F61b5FJwDIQonCwwGfJXUMfx6/cKqquBSnK65Q1ylf9mZnMibe+rAqda
sVtlX7pQYuoJcQbU8nloK/JDLdxhVVsMI1S4QgBEZpSNx6eML7bUoAXsU6Aas/BISqB3qHm4NuDO
IQ3W259cOxoyA++9dYyMS7LcBmsy+T/Kju+EKyRkCPgocuHogn9+yBPnLFyNKqN+nnvqZxPafxK8
ZVqT4B7CKT8sHs4ztkWS6kfmzNmNtr4zSxqDtLRULBVXJrk9PmiAoq2kgSlpVRgJgz1yTLN6gMDj
GuCDYkVOXEQbA9g+wGGe/5GMyPxDungUFYPcKtTYNu8gRpDxGjq56VlsfqV7f2IbNLrQ0ayUR67l
XUpmFqnWY8OkpiO8owukVZkVEeHU60IIqp+ZuX5iXel6QnpiTyL0jD4cWkxYmyx4k/FTEXyO8hio
h9jVq+lebww6MbG8t1TWSarJpwZSC/oSwumDRguxytWH0X5gv2cRVHu01t/o33KLQOQByJqQE+Qm
RXo7opVtOThTnEmMzvZqEZyld7l3t5z6s7elTUEPfQ7KOlsB66fRztGRWv1uHItyFCxmyFoTIqQI
QHOaHC1XrHJf74Z8TKoa42d2D8xfEUqyTAXmg5P8S5fuHSvbUDZk69vmA4wHiAT4ZCoBTvhbnWbZ
bTPZcJUFFUJS80ZQE8mWYRVnvmD7gzgz1pGeFGN5GUFuWXW/gVQAVL84Hp3vV6DwLh3m59nGyLCW
JxuwH2KcHqy9zUUPnCJIAhfncnktd4+IfRIj+LpxzDp/xzqn17hWcxD2+/4HbUddnjXIY5AeYayY
obZ/4gfowt6v4XkGsIlTGUx8kko1GBcjDGtlCABzkLWsHgbbNQkJN32zyi1ptw173N4RtszxB4LM
a8B4HnKEltGoZdtKpUToS+DSMjFOXUlnvbBjbico33DHrab+KU7DpKrXeacYQGDe9wHDQkthXzVG
csjmvw4BDAAv4okmfvlDlNoGlw+CEtQ/zPtPY4p9nxylC6u4hDy7tNf5ld5rjVDQ+fCsQa9Pxuwo
wsjx8XySNbs9j77Lcgf50SXyW7mWXvXHN6NEVpAiRClyK9OXCBprClplTTIU718eAXsp9wzcf1PJ
+JCRX48nxv1fn7kiTghWLvEr/s5IzkCdzw9I+uEFYFg1P2Hsf0ShxnVFccRDCocSVZVIIzrmmdex
bghAhbqw+6dZE0vB5zM4NlC15Eu6x/d7GKbGXFw31ic72mr12DgUvBACcULOnaxyJRDRLLIuNOn4
5sG5CQEde4nO4nFc9lzSgK5XoZxQW6dOAgcwSTIyyVNTvQI1bRDnU4WtY3OzMBLfD1HrQThuD/nV
zJ+Fnf41smZLMGVHaomyfLykP3fG+k3cNrIrFE+zbXuVwVV2kLD141r3soX1J/xB3FDNyAyODBVv
EEy5kTMNPwdE+BoNZJYXAn4SG1Lz9enNYRoT3dDAoq5aIUw3LmVFt3i7eAOdFP4yDMaaVXGPDdXi
G02y9ut5EV5CCilgHvtuhYc4MLJBerg+s14O3TdJOF2Csx06BdnQwWv5Tdhf5VafOCIzQ90IfZrG
ls4Bmjze+GzDKvI2t4Khu6r6JkfGaK5zqImc7SKLjLZ9uzkQTMtA6VPkEQfXy8IDbzGnY5FlKXZ4
jo74At9atjHFBzYUwA2kfV5NV2Y9TXXmiQqPBhqO1aiCSHq1/ILKr9TXGwtaMJWgdMcDkA/B0+Rw
AdUrHUdmn3eRgyFQjgb1+xZ50qhiKehg2Pf6SlqOh8p8qJPxYWafwPbXF9LrOaW+ZRE1Mb3dN3LH
kDX/4pr5QpDPz8TUrpEotpoB4R5kwNl/yTIUF5futtGSNwQSEgr50zvIcWVuHRZAtsHsvff5Baz1
SFuOcx7mog/DC9wBAJzbKAImtJY4+i6qYrL7V0hF5mUxnVubBbZ4aupiOOtUJhWciTz4jSQFJnMG
kO0fy8ldNHk8EeivmkejzP7DayO5k+yM3SYqM7KDU364R2DdK5xJRBSkNpAnzc+v383L5UgNMWnT
4wnfcSqWhpC5vqvY08yLc1cGHMkYujkNL8/raqr4/owy5EzN2JYH6TnhT17uKz606kS4nLswMnz1
Uqf3OoVHmJXf1IAGVZ3pnExxcWkmoxT02hMz24Duqw89kEr4jWyKb+8bxLXa6fKDAvGkJeU9LwQS
WpjCiIKwazXYxkQgA77YwL/Y9ND87mySseQEWyyb99z5ycxbH4boRBd7uECt6qK1YqvPwlPP/pTu
ZiVy3cjNGADzHSzD1Y9nFh2Sfp3LCeCD1yiUrKxi8KK/gZ//TyFGi0X+oIAP8dUO/bCNuL4qOTvD
Nrz4zNKFUfbPlxbYYA4tiyMAmg/EDwVCelEXCT74809wwIcc1qs0D1lzGIdxv2NSttsE15W7gPYR
hk/TB6X8HYQ7gtKufXqa9Z3mHmWOOZId30eIITIkRPVjx7pNCaBzEHwH8OntKlyZIC5Gudd1zvYs
uhvtoV0GQsPNPJ2kyu3EcJA0ItjPKUWgFSpzjooDar0hey8l7YLUeVq/eBH3TCkBJMchh0mvPb3b
FsoVUS8pjjZ+FtQ2NCpoCsAszW3Ii/VXydgPqUWKYEqtuZY5/bKD5COHiEkiIPVf0+mQoIFeGGEW
ArOqCA/rYTDqtMhz0Dbx1QH+0Ir+LfNyYna8aO8+Kdi2fJUnLixYh47jsz1Moov635zQRaBNMbws
JSdjoxBnoVACBshU0N+N11LeeYikh3SlZ38vkSlV2/uWGL9zvflOqmhXDF95IiQBsSblniZ3aSnz
MqKoD0Q5T4swciOLPq+JpfqzJeigucl+/o+FC++bSluMC+BrwG+U0T7K4qo2144TcyUeNn+lQ8K7
ZA1yby00yWWHPfVl5Y99MiS5+iDc2TzTgbMQXbHs0qbMLhy4eHPll3mcPEBi7R+grty++M7NgKqd
2G2ahRZg856tAMhjYgtgyc2ugh/6/P0lN2LN7cJoGs/Hvz6yES6bU29TYnYYihPftTkEbJLuMyc7
5UpTkzMMmwgurMJ5rIbg7lXU0KE8grYSSpJO5zTUS2Nv605ZbQvTmrKVK9Qm31E6cnScO7aDzvuK
3e/91VjOEJUtvIM/PHQHZrCqQxS5zBfeP7CCIf1qbKGv/7T6X1+Pf/N57Fv6dfVeHelpSqz7SkO5
oNRSYycKZTuwc7g38vYikRUE2pwBBqyAPtupBjlpQPEByj4ioT7hPlTUda9oI2haTnnc8DVfSRBN
+yg7lefu+4fOs30pQe6KsYjPFe6wDulVBmjhE6MpGV8eEQS086qlwL9TAVIE49anLZuWjeYTDnui
6wLEFsJio/H9xj8R8tx+aOwKyPZZKW2pCXSMbyU4q0JYp6CtG6P9ihr6LqnbJ8eTPcUu2a0yyqdy
J6HgN5DMmuzrMdf6+bggIcy4z9yeShjEVihFZ2CANquvbOrVFEYZXiYGjZ9+cmynM1N7pU4ZH88f
ToDQWf5Irlfu9o3dKzkTtb3DkYIdn6s/4flGpcCBNN/IHwXuNoBfkJN6Ccy/MmgYDsPpUCAzKp5H
4sQpsbPUsrJH6mgFai5wfVpM2jM10htWCG/zTS6kGMudQL8RWGUa/WkFm9QOzYTPCHODtNk3wZrm
7870xgfZrcupbzTCbLc9TPWeKHAMb+fpNiYtboWROfBkv39VimsQTGX1O+NZCEDTseQwOAPWVRlI
wMPze5Pr8dgqwMo7IzjvLPcbXmFt7fgAP8vf3uoa3COA+FU4FKMm6Fw1glxhoLDKls/oCBhGhOXc
94I/KaCee+VWT7JvaHZSer1nPKx7veA+egoerCoucalQc2sN6PJoKflItCGQ4sR9HdAcZznyaRho
xDJSvnmuQ8R5WytRfMtj49sCzPuQWdg3FEEIl7ruyd0sio5+dBKP8AkaoiDR6qfK+TNRclkAs+ZQ
O1KZCC3rVHSqjWdnchsHDYZwxtfr0rg2/Tk7ZTQdgMkUAzTYiygG4vFkmrh3ijYZfJ5IJ5P0wk9T
+dhVhG+Q3DMCiJxUAqV4/sAWIVptpFKKeAMbON4Hwuy6gr2K9aZhwkT7jFi7KGixzA+Q1aUkgsWt
V+QcBoQH5yhFM49VK+c17+o5ln1L3lxFYFNgl+K66qhMA3g5ryENlU2abY6Fbw2a0QyC1LhbdvFk
VqLevvFll9YK5YpSXA0SUZaJtsMfXTK5EiORTU+gl4l71iwKWTojoY7GhFHqsPQkbFrNKNpaSJxk
AG4HlS5DB+LoRydzOUeJvoDSoHaxPjGXK7aTpj3PD4/NGMWYUHZag7RQTF4WnSCwEJ6tWaA5P/ld
npzQOmHikwlVcBOQmX6wOXUp8RZKMbdGAY7Zg2Soza96QbIQPoEeujvwQ9sB8Zl/GSEewV8k9Q/o
H71qeidGpGPz7NaqEh831zhsktckkGakETZ/sCL+BUTaZl9xR/PbPoP6yHtwknMo5jzCeZzo7wY5
I/4wc2dzqhIsJkfCXkxch3m2ri5xmAJzN9eHRIElMPNpshsK2pdii7iEDC4ZzVDMaqMJqoEpG1t9
q1cjQ6Xb+Aohm9qg2NX9o6pw+exu4Jp0RWlAJKoeBAs/kJhTCkVpTM+jxtL8sZ+rueFY/SAxZayd
2iIVbhFvw3GXRkHw6WU83cE4/fV60VSr+4Z4yP/YTobcJC9H2C6byMFr+At7BaNZ/ST3iYIEy3UL
aBi3HF6aTOvLdFWpLM37e3jEgdiFMv1KNDyq+s9iKKDDVKGKWMIYDmGhXp4NLJ5EbA4IrlqXu4Nd
NknSQpIcVwN6ONtbhLdx8+B83iAk+9T+ADuk3Rs37wF+QilfPFgKiM4aaha1PTZNVob3YyuB9lQZ
rrKn8QR4P+ZSFYLOiXuoAbZyUsFlbUMf0bDig0BOX7IAseeJ7K07J/OBmeNUEBG0TAPbJnDGrlve
LS9Wq4KrlVle54+nYkEpFthlEWampC/dZ0whaaTxSvIUT3DRSOjfY6CgCfwGXEjH/ev43Udpi6hI
BgTiyebyaE0nknoYF0i07v47RxnARzlW3L8vOd39d8uLPdbYyqpTRqBFyDxw+IX5kj2iwDc5r6rP
emPDQb1la9adpV9SDlO0EG27MwC5JVeYm5xWCyre7Q9Pxscna8Dr7pOYO14knnYVFwYpCdxYB+0r
w9og8aKYll7QUWFqZCC9DqFm436YILHrPlQWcaOTodTs9W9tJfLdHQ7JyOWb8gZIA5PKkLCrwE5X
+FJod19oDf0pKXmGppKq/PsXl22MZaZ1cvYgqRWhzDUAW1iYr2wPGzAaVZ5Lp2PCrs7C2Ka92c0R
LSksN30YMAsMvccwVIZm3aCCZaKL0jNFCU06CxRbMP/n4Q3rFyw3jEBlfOcGgvDSYQu0DGZ1r2L/
iVZwap7xqhg/n2DC+N4WAkhqBOdKQ/ljC7DNxWZ61Eedyb+8HUN5inQ6MKVtLoZGSaAzzel4vDHl
bLrT+ls2ozcRHxh/NGcLqJy2sIWuBWEoP4Jbc6aD72e6GFiilJ3Hh98ULcKY5u4aEj67ZFzO5Jbc
2F+Q8oTo2hr8Vj23MStIiLDqtNTV3fHt3qrGWeeIxj+V8tawV+TDUdYYY44n0Vx/IB9XX63I97pS
JfLTlp8/pFa6HjagvkWF3OXCgP9zutbx6UTByPiCu/wFT30o4ONJcJQHkAj+MZ+lauBaQivKpMw7
9WwRX/fR38gTMv/o3LGxtFDQSYEybfGrq2FIWUckl79ttVJgP1M0cxQfZV7+Y02RI8o+C8GRvUal
QOzRR2Dtg9UpM1ZMMlUg7aGeO2/l1bDfDKMOKkJZGtW7h0gRd6uSx/lYDDlPiGm3F1pufxmgHhDP
58twnoqkOK4/rmmG8pCJOgP9VYiRiLY1FhQQkeLTS6/FDDRUJuqC+n5WUjTG3CgOZ/b9nNv3xfR7
VUjGKUjxLRpDJkCFBZ5dyReDVIqe4So/e/8AQ3kdxVD24Olo3QzbxDhYe2g5hMJ2WQF2Icz+uI3/
1yoLvHn8DE//HwaVGRed5W8efs9PcwNzHKv3zZUGRT6qGnAAWmU9NnlimmMVPPFEdVgP2yie5ySa
ExMD5WfgEDkBoMvutcq6svLhFCBpUOpiI+l82pzmmQT7dkJTqxl1dkL7eJrCKF82nn0Vzc+PYzi0
Ps5RTlfPlt/6iWuQDSHR4TWicb5L1unyB8lQ++WxcuRXsXECw6sb6dooabTF7e/uzaroKz6GqMny
4WPYtXmgJ7s1QUbCqBVifuPiUbDL4FLjeeNsu45VgHtbcPrvUNtcXl+/6dz0pRHykCayrIXG1rzB
I1+e4dQazZiDMm8A359rjOQLz0949CghpEz3kVCU5vAlko8AwCnc0/dY5LMPhStC3FkERNA0L5R5
KFx5P4/9wo7YSnAtrqREhhssMnZBHWLQMsbz51TYtQczyvCFwOOzUrAtimB9wUAwkUYTo0VKj4jK
FsNsRNMs1WxJTv57NmsfGGyKwf1YBVW8NJMqO+nYjLIgHkFeOp7SHD8/Qh3N0hW/mpYq7BDBz9HS
DUYNB4Bf9+3LW3GQvQAuelgYYvP+IEBkNgoZi9iCSxJugp8sHSxyLHxNXu07qJeHmX577WPBH/nV
KaLnJVdigKMxQDGGLALjXime1NhDHpZYMTVQeiNkSSg6qoCeoMgj++RPtt3+IvD8VxyrD3psqi2+
76u7StjhIwEs3ow25+rcNnBm6izglO703xwJo3MryAUQrl830VX2CEnkvJm/j13Rjr30mhj6hfYy
8Ol1/zJ5aYxUpXjXKAXCGf7Wtf6fFfwWiSl2YRxRKyOZ4or6EuXPtvT+4UqKZDpLWyN0fG53QGJI
DNLR4gfiDVstiHkEtwm9xlw927Lj9s96Mq5OydkLAuznyVfPvoxla88e9cgoZYbgt8mFj79sOygl
sQjXR4l1mSkLkmB8hP29NnvcQRf+N0LaSHjlxO7Ff+K2fxm/QZ+aE8uXBBJZJm3GXBooO6ROxj4v
j8pqQbXxRUxadeXvoRL/eLxx14gqqTZc6ZQnLgmfnwyHh4gWoRqTJgdSieoiBoGxbDrjJ/15qhzy
LPdHHUowEqtNBqCHDETgyAC0st7Uj3Xvn/zo0jJGVRVM2WiDZufdxznyGpnWlonYzzYy4rVJgBn+
FgytNcvo5hhH0FZZlXMbYU0vzkYYV2SdSXCKRnWRgbnajEWLCLFLk1GEd5kttP9ka6HL+4z0ns5Y
a+rqWNtfuBHATbpWmUxGcWZDdVQrg0VYXz7ZyT1EchWm4N0INTt1B9P/Di4qpWoon11+Uj2CzVpR
r1KCf1WB5XvZ9wBLITOxmkg0zI+99mYX6X3AQPJgsH+UR0HbYYZ9/G11h17uX5513YjEMq+fpzS2
dgBqaZhIqC8NDUcVZV93bUQRSWs1+Qg4zH98V7LlJS8CMPyzTuRMySRy3qj5FWRuW1+gyxVpWjmQ
xGrGx7XuPotRHHc8hM5J9oHE99gAQxREqzt0aQVyuN//Q08vAuyFY6q1BkBH2pXC4iw7TQ+8CfkO
r2QiP9i0kLCcO+nGI8i277DdWp1UfPDVq3hrlSDDWX0f30MExV/31WD2R8QcwBcXyt8Pzfi9CXqD
iqRrulliJAjROXgBTpY4QTJnt5OUCUNwsiLh7x3gdErapKJ3PeIMUhvkXnXk39MOVvnh3AEupi7R
VtH863tWdrvCr5cUCtI2Tx1ELMVj9sRqVaumuUohf8qYTRuGw/UXedPBahPq1EvMfV3JyO6u0jEz
473T8pIpV4hFL9amJYukgwj2MzP2v81WGf+NUF+FbkcW4sBd/2jbpLkNQGh628DYvCLxYofxReoD
8/eL1cdw6mq3o3QaX1Ddi5MhTHj5SJVQzbNmijle9ZuJVmrXuc13KaT8gmoFnTF115usj6RibE1W
NqWneptw0PIgSup4+Pd4ih8IpHaQXS9nWQTzF/wTO00fnfTMSRUs0vYwr+qNgo2DoutAqI7HFkPQ
27tFHdOaLFkWZ+LKYkCJyh9a0OuVCM7q+So9+HuieQLixZYaduqKHMeHnySPlUz2YFohWyQro55W
oPWBc7cIakAp9arMDpYAvZ90wPqOvsh+bP6TP718DaTFe+Pr3qO0/UjRP76OoQwaXO0FgJ3qYgFY
tDWkIvj4xmSnb2PNJs7dK2nZLjiEniKBP8oVET8R8jZK980GxUTEKe9/bEZkZIypdpOTKMjksCDw
dpARTlSKyFc/u1gS7+Hgh770WSJCAt1v1pdrS3gJQRIR584MC6pHNRhAmN4VqxbSrpj2f6saC+1W
eJ9T97ptSX1kGwrli7grZo4J9T+fV4CG7M4N+UGF9Apqaotqngkn9WEY6F9Jiw35B4w94pG0gqbL
qX0HB86Gs4zZ/y7wljnAhR6iM+p4SijJclNABv6cbwco3Hnq+79YYjOhLVIEMornfFDoAHzejkNt
WyrOzR2ld39Okk3+bB9GTT/oUIY/obhr4UYBmfhucWq1nZlOL8dV4/nEQ2IrAYfCWPbO485zwkwO
Fm1JCjHOfEN2fyBnnwbRnholcyGipyvARjladTmNb2ANlpGr+Wgfj56HPc5EWoc9F2zvIvpLCwEZ
A/ALZe7aQimZGhvhIVegUKVctUNKjCkI7CXtEg4ixAJ0sQCSqrJCsunPBm7tUupxzG4ef7ArFbOI
NuwDPnZmlVdVAnft9tOl1naOVqiznjNIOtjUYIV2T5jRN5qlsSeB3xScMhPniP63QkO9VUje5MxW
TFbm2+GTPy42iT34pAtkILivViP8cVqPa9DauaQSYY5WzXs+wsR0EELFK920aS1G8jn+ADVPhbpg
fwVRcRkITH10bvMiYR89YKi5aXT9uIOn6AhIvquelGMiAtpODrU9q4ve1fyvuZaywkIJW6oqUhEj
IEf5UGZxQhnFz2WSr8EPCFj/NNhq2TF00dvVUcYCrQvUS4jCOvWZG8WdbzF/KZIjNttu4L4G0P1u
sck5T9pvU+Q1lg4zg+PxdCdh4+C+NaCiLGamgygq/Muc9W+ekihMy3uM4BmlQLTevlkcn1yAEvjI
uYzutpDTaV0s3bwSZxkSDqLB8lUTSHEmfTAcAQzI+ZRU16RaeHKEsScQn2qKaDorCCetdhUgmmVJ
jmSab2V/MH8y1Rq7fxtRrFwboNcVF/lXjYTJui1jkcVRKPFfEq0l5Ab335JE0CvriIATqZd3NEWi
nWHMCQqgaj4NF+ATZN5wrEGmFPwz0QcwypQMOZoV/GHf/Ix7fYa28ggPr8+87lUjNzB3ioxawa8q
Og6yUv48Ew99C67YQB/tduZm/zinuRt1pO9bclfz37TyJVxAzUzwCO8ci12ylVj0cq41zFpx5jmY
vv1AwX7Yr2R8xnG/xkgRZ+PGxPypnWAgzV0dxjwIF2T85HeYCFTRc6ysFol/7lW5dSySCy2IeOEK
uu1kVNjcu4fztQBsGs4yI1zRpPlNLX9zbigedNv+ljawqj0jBaz6S9RR5C1q9N1XAbRdXB8kuMY+
NX0ZhmEkubs3+RBGdgdnjr3esAGdEdcKywB+ThQupSewS44oeK7MK0ksLK0vvHE4tiM7SfkEAgl4
BrNWfzlwvM1ss34c4CrclmLrzvra+Kcw44t+9SpeHwKBaiv2gIBS6VmHQaWrKUGZAcA0JyLPt9qy
UFfqIJLmFyITKdWHex+DNP8m8xHzUVqjQbkfH0Ewkj3NwXTxkOcLzSeoqEaqWHyqmL4JZAfzgJ/s
Zb1o+LzhxJNC4J+FxHcpmjSEoGfb4RiLUPSG/prEMk30xGUFuruP+x+ykV7v66TsAd8ulcACpSfJ
RNdx6hlQq4tJq9HHf+lyiawItQX1610Je7eSyxwo/wL1h87DHZ5cm4e6ubcDnrBaz/ZmSFyhxaMx
DMZ2Bx9wotOKCwPnOMjaOHMGfaGLoSSHeH06aU3ELaej8xjtDwR2hf/NEAlFKyVUIgn7ZKfhoenN
aLBkGxe+sobdHAKLe3Bp2aBd1eoORDE+nw7x/b84jr/cMy7WuhaOmdrbfCjOwOX/xLx6GRHnDZnU
zh8BdN4hqjHcjVHjsBYGoBPpn8+MRY1HIyeilFngYMgPcbzs3hBqHKXLhmB0gSVEcETKIEE8WFpp
6/5u/95G3BX8T+EMH9cDG7OXlvLwO+CGelBMCpZn4FrOY07zLDEA6h5HYcx9qCyUjdZjq7ocee5B
9JFD+1NxwL6F0Ii93o7RR7b+4A00BNBiQ+hBFag7U40VkOXsQXFdv0l2aUxXRkEywUDBxWZDwtjV
UoRX75jYlOc1Dho1nMWWThKTzRH10AKIrGnfkLj5GXh/paDkWioJcb0IUbr4BRoRDwMtHeevHQjc
gTSEHwJTvRgCkBcRhtDqSn/tcv3BpCtO7jKBKdr80OzZ1sINJO4LEYGR0dTYdXvuNOODR4KWx0xY
Kye0lxm80X4RVK9LXjxB2lCiGbmnN0zr2hjfQVd95oSVJPpNYO1kxx9j/bpCUaoho20mljDdeZZB
03JDTtwlOL+F5+1R2AjsonFM2oYGVBJ1AJ3ptQZB8Tyc3s93Ts6XVFFTuAzEgvMDyLlQeFmYvudG
mNSuj0uHUzZQr7Z1FZuPJejQwAO7KkfQgFdxp3yUYtaeVoedQWDfo8zWmPlO9lmz1Xul4Z1bfOXd
Y+Ge8GkxTuulqNFBQkpWYqcCEkFx7DhJeNwoqvrDJU6VmoohAADMRGytC7/as3L0EbKyEcrCBe/t
nt0LrWDSrIqDB8tMbHnJHf6NdeFNnSfJbDCyT/HDmQMWOsWIKNZ0KfoYPj2oVVzaPJ+UvFB5I/Gx
czm2Ry6y0BZYbX2AOZfDDr2bhGnW1g8ER4bs0Ci24oUjlnCGreBrzabLqIWX1DB9kpGXHzE+Yt/t
CBHIz6qTiGfiCQ8DWT4d5XLJzFOb7cZjEj6LJF8AYD0sOL/LXMVYaARVYqSy/vcuCfFKlmPtYi6m
MdceUi+rJOfLYpDKhill0o27KK5QQkGX4/3z/lHFlUaAJ14EZiJX1QmnJCKjniBm8avBgXN0dnMX
kjU0ikMqZnM+9VbqhMoy9rCiLVzm4ecVQDhuho7fovdcVMBaT0LPgvdcJtue8EiEo9o7nWJ2b10i
tGURB718gX184vWqNwHlnIzia3n/NPOaa8xw9Jy0yKf0/zBCioxnmLJuI8l1hWKd3b02AvFmlrco
KKUmnKpAhbjpkGTo6z/MGULT2QGqnz8BCUY21SnzzQu5c48EfGNP10vylId94l5xSOZS59Nw+CLD
ahGM123JLMM8h+EuS/wVPmCUbD20NwnIO0b0s/dQ3hvJhmqRWlbN3HfbHThda98UQxMIvOqecOVq
l2hNpXQVDnKRoMj6Oisxdee2fu83E/LvhDjaIPjab4Pjh9YExJysBdLc7zRcYpSXAQqyD15upjmB
Ua06douEuu7B6ExbP4J8wyfXmx7EjDBH0+OEimYZb45aidyqHmktKukR+AFhmi3WaEGU7K5adoFw
TEjaeVxMcXga9lwvl9cEzNj5asNkIDv6vzyvtoMsMeRU74NTORBU6ZqSEX6lkIAngbCkkmEvG025
XRVZmhpmCBi6+cUc71ucolKvcqkjOn9bnZuY75HPOri+7GB1mjuoearkzf+YQO3EEHIYs/6JAE0F
NH+VsLqiGF0EHuJT6KF8vGq/vd0J+T7HwKJYLDGcLClnolsM+ovjPLAMJg5SpKvHTetMaALEgy01
NhX8yvSNsk90nPhoOS5KFGH/DWxVz0L8q6vsiBqz6op5oyZWY/n5TeOACwBtSZibkXW3XVLTSpvI
PbX/zKDMGGrdxSHlK4TOrYOKGQY8yZ6FMS5ZJK8+PTK1UwRPEDh/XKQtvfEQ3LwM1hRAJFef0lK9
4Pdyo4kfaail4uWXfbVsyILBVDABH/aNm9hQ79l+b+niAcftoNhBZnzpVUa/PVFaFCJn/ho5bLdQ
lJuPERw4v2g9R1oA74zPaVMMktWez4k/4IUEL2ODLg518opkV7QSLnQ46gB8Oy+aRU9jTBT2Os5/
xZX7xYAohLH9QnCTcfJpwDvl9i1KmTxVeee2eOis+PJT27zTEKVQtAZdhx2NhJBnaRhGjwcl7sT+
N1LikS0PzmZa/krcbzweIgtsVfFm0PUslystQr41P/Fwt5vDM4IXI9E/nDFw8KanLX7OekF29WBW
jsAH+5vjHLdH9dvR5pqKMvsx4z0MCZPujCqYlMWm4QeTPVWFxAQul9nqEBVFsAZVjg06mqk5vF4z
I5iwuGMtjay5EQ0QUbpc4L9AxAOEJraSQ3ImKELC0+SsaI4IL9xqUiKHiZB+rL08k3Kxh+AFGwTU
1m1iJ/OIDFjv9i0D2BKP1VDfWeMF7vaklazq2IbFKj09z+dTBIh0Zz3idbzo1sNV0FNwj1LXUK84
U6W/hAgsuBIK7C9BQTeq8cwS5ahgJ+0e9BR9YPNZbZiDiy0Ktv7/o4KeadmsF7pQZ9dSBlMfdqqh
Iwxq85nVurHK6bnwHdpgD/i22JuTVvGeopRm5RMbJQGzL6CIsADAQ7xCw4stcA9u7d1AktDlsDP4
430P6qX7SFiGIDVbZHiVvuE5JI57Px8JmVDnvaf5hgawiagS0Mr1EPFygE1QI8JT8452CFjhELJc
F+Eez8JoSaRsq5NY49iAlH5uPOzZUpRgnfIz67ZTCvaSANOYoojRzmveYos57Ux3srG0WyZjXxUL
fY6R8RsOpcOjqYMr1zzkT6qy12CwLbCGhdTAirolurw3AxgJe0sNZ3shEWCNLlqLpNNqbenBgEA+
YxQT+4P5hx23065O6WfBBn22bfREek5frs2QJsDpIpA66K6pgrKguDN8+7ByY9PjCmF5yheA0Hzj
zN5AZK94/ByasD912Fj7XCjlKxodROkv0DQNRHQOBjYvliyqBs8sUDRfxlSANi6E3h33pzo2P1uE
6cVjplIbYi31LhlOHWpxuRCdXFs8VtmbS+o4vi9mYNXLocnPQn2EidP8hNcw4IvbQZ/pdEXDLsId
PctC6sm3YYzF26RUlwNs4LyNi/jlHNBPi03Dx/0pF2ruG7AR8XMAslN53J2Kjfuigktoq9n2Zm9t
PcHq1UVmBobRNv+u6nsv+HyEMKKKZv9tpZq4ePSLKFUw5ZBb+D/gqE9ErMQORZ7Yljuz7GGt61FG
XDXFnqv7jiTm32PoqzlHIA3qk049W//Fin+H5lkClNjHP5T4z3GDCrPYyeRm1qiUyha6TPxHOmK6
4u9oqcLNScQoVflvBdZ1f22sWEEDDNxDnCFpR9uz4jEa1cQtAnnjOyw/fQnwnwYa55/nnOQ7h1nr
0x6hJIKfpDHP2YapxVJSS+OC+v8+Rfakig0KScVniZwSjRV/eVzTdOniVmOq//uIri3+A9DBOP6/
/PdXRgPKDvNp30i1GzKiabzgmHy7f9rn2H3GWunYYCd1DJqqO6xKvRMXfAoTxvBdcspCx+/zUXXe
sJW2V734sIssmIFa/AhXoFAhLkLArsJ0Et3mNK0BZF+lRQKpbV8TmkQtgIRGVO+mkac/SuzzwhRM
wBhYGgz4USNlFanNEza4swSvvWN8WvBcfcqwuQyWCWnLK3dqPMSL7Bb6WFvXzUhzm7NTyWX6aKhV
z8qGObaownxX42qfMA6Et53AEOKXA4kJGVBpU022613XLJLU5FXTg7r0a3kGUlmNIaeI2MGIcShp
4aksrS0PXgogDdcnONUCZ+RC4GGICCsq7XVCV/va2uHz1E8DIPFwwXC7a1r3sabn5NrdaPWGTh4w
bZlSGh2UdQlnzKd2xPPYr7mdU77aBJJ6WYBqCNukebTO47J92uTw2+9aca142fJZ0ijkkUnAwMnu
QPE8HlBzUF9rQ0F6QPVMnMaVWmGSi0eUR74Z1f/7/qRAXfNVRxdeVl5rGvzAxWkICgnzxDXf1k11
xFIfW1ZzZ4A40yZ8cJACw67DosgVrKkUdaVlFqDEQEDhgKhZKvIjtaFYamow211H3t/e4/99TswF
i5wuEMBVcRcxvcAgzUosH4tm4Xwpz5Xx2bdWKii4Rgxxfgb6vtLroju0QHw+Ejpg4Jfmx7SUkZ5m
KDtdg5bCg+9ufrhXe/t+YEJlhkVO14uJ3XFAp5aBpY+/+knGK9J1E/aFQC8XtItECnYn35PDWs9J
1h2IYGxiSKkPTxf07dq1ZliPnQxMfyqyVXhe/nCOq7KNq4RmGdChnOr0m4OLxgRmKractW6CZEsJ
0oU66ECaFBr679IU4qPYrysdlqiAr9Ae1yWM0KYjR/mYaMqCQZ3UcwrtlkYvwJ2AlogeHvSAudP9
5oEmwJTl3Cx1ZN6k8K2sVlBkI9Dvbg+yGgo2kVlFeCzKPKbZP25fvfpOPjHvRKZYgC0+4Vfv4LZc
8W3+P6ANp20OWmOGW/CtQvGHzDesYfIIMi9g/bB2YZlAuf+Cs0i95iyjWKrCKgGlWK8B/PIiPaTA
IES2L3Ue9QSxSi/yRsPH+eOoWLq939iAOlId+adaUYXh5WKfs+RhfFR9YdaUfMOobWm2M9QHaI2f
EjdCTsynSRellm3LoqglJnqbFHdvBBrLa42kLjl70xLnfjayz8zGBNAqRPb5gULzrl/8keoAB/xn
I+OFUMZXcUAZZQa3Za9ZVn6PCnGG2E/5b2nRDWb+P+IXt9gYLRWeGahNxAqxcrxZ8TUur9ncWMnK
VGeQUwJP2wpqA9zSY4b9uBqmctaUyqVSSd150Y5cghLuHTl23kuKfHu3uH/7T7Z72NoM1vpQ6JbA
n6gX2mCj6RPYoBnfazjHdxeNVN1+xwfGRaWWSiRH6qSslXf/LRmbahQ5AMPhhdMPAFveQz6HvZlY
kGHBF9jTKSmznfFSsMN5aJU+Dl8oqi2eUXdMHQDT1VfsK4M8S7tXTzyrGLeg033C3Psbaotb692U
+IJHkkoaguVbv6c0numD8Hc3/EP6zOEpGhzAJAZxtjzMEmKDooBUxcT0QxAHHW325QjCN6skH6Il
4voUuX5HTQHu69TGqRxd8aAYp0hQQlGfBSYLTLxIzXA819GT6Q1piGoog1NILBr9ak/GJUmMYDU7
s1rmXOWarFwTcqUKKyTQvY3SaK1SR56kQnwh3h6+TsKRW+SrI0GkijVDr7VyAbH00rslG++JsRfX
Tm21DkbLLlyaJnon0Dsit/c2anRHdDVvDn8iteteD3JEthXjjtpBjO4Hod26HI+hj4H4Bh16+Or+
9LkCn3jxOckUPH+JJq0BH7vGhFTc9NPquBVhFnk9wunoK3m0vbgbZ7u0Vln50Tl9H9ZCWfFJ3NkP
v/uruu0PE0bMzml9cqvDy0RSWX5EJi+BLaidhRG9OY/11FuV34FxDp+2/4szO/hpvP/yMxi5Oat+
uZvmes4LywCkzj2brhrWjAdHSAP+8xvf0nm0UaUSebIDVvJV8sm0ivjkQH6H1t7wCVsbLK5jJEhU
qpYN5CgJm2hIco+sDkL1W21kyMk9GV38hAjTPPfzO60egVlBLsvkZdpjzfig7QOPGBoX4HmYPmOm
1rUGzEiYKYngJZXWmkmzEQtH2nen9VCRZqeJOzkf47QkQhy3wPg7cOsU0nWxWToRugCZmcRTnNUv
DFg7zz+hX8VHGUBVERNJPFLfHUTlf4GlmBLxwAFuASojNHyRC+38GmNmWu6PiBTkpJNNHcG3HQo2
BWMXWz5MekkBICB1hIeLGrcl3CrrDEWjjrjjPYrVMdS2L6XLtzH9T71OlEfDYTKsgaNauGw6MRWY
eEjeL5zcsIi8cxhcBJcXzC9sPCI05BOnopW1JMHK6Nu+CVf0+YR9zmVpfi2kspOxEER1pnV+pZPu
fHzfDH63MQhIjSzsR8pCtDZSA72oUMENoU/VVd6EHs392qWvtbeZzGs6KhL7QJ+DPvV7UlkKDfr1
2EFbuBGQ1tWgIijBcQs8D3E8WfJgLl836GnNTEOG8SSLfP5hQ5ZxHNGuBZ1UXUSqnG6dSAasvZZk
6QniWHCrGN7Lgq6Nrol21stfJZmeaSRAZoqe/1ZjJQM+ETCPjqLa4tpg5PoMlqMl/zOypB7KRa8E
An6z3ZSX2oNi7iK58QCWATIMPfH24uCKxh8yLcOBzoLFxz7oostZYa89X2RKQb+iiU/AIVL6RKhH
mLbwfgiVOv5Kdal27gZHW0GpZu6TpfSzlfQGSx7feSU4Dzmvvh4urThifoqmTRwrW9gWRYDJBb9q
1RJgkO+JTmp8z82LkLM9DFN4weIKZ5Y8t8om4flpSY4ynUOe/oCbR+qL+xQzQ6u+SqkSn9/GwpDa
h+eAQGwOxQ/P6vjl5+9bwS4BHyH20AwsNHP1+Jcs3j/DX43KWexVDLfW1vtgPGcAUyBjnsEEWKpa
5G10BjoKMJGscja/61I6A6ESrFQ7MpxfFlvaXDOjUE/UGbVKvNngNuvuD5fxlOdnlInvow2oNBjM
S6F+QjkVyOG69NKdG2hYzZ3VEbuh16Cu3qmUBxGHY3mpjfHvpUOwCssh2DJYtC2qTTNfvT1kXbfB
1GM+O2lpnVDlvZx4EFoWILIXx9SlkQExREuol1x8I0OLtLnML8xLYwPFT51pqelKFHbjPZpAPN7Z
rsb155GMyZqEmywUhK8f39pbqPgT1s1+6fX/0/bDrfgzKnoTw7XRvCXhzO4btA7DfVylk8SqmXFg
kSPzvA/baZIgaqP0SeHs31IlaAySH4exNOCSvg4++Q/UxvBQjgNNQu03DDDpP6fCB07ArdF30DjS
kS0dftpWQgaL+KM1z4PgDBlKBdYLl3I7493Scbdzy6giRNA/X/stkHESlLBQD4Sc2gE7KxmpgSK3
otZXxWRv/lSa1O7ruqXHlKGhdVSkztLoxYTseEHCfItCR1ERUGeJFI0JMthvw3t9az9FwYkzQItw
4LBYvwhRgLs+DUYgCry8j53n+koR085Z5qfdWIxkw46OUlHWyz/rABPrY0miiKYvOfnL9NwmMUqg
Ozj6Ag2kpR87bkfYjnjDMWxS0YjgIezhimQic1m20ERRXMjKsVPNTMijKN7O4EM/WmLRQq4XB8cV
f4JA75vMgr1A7qyDFI91eB2FJHeDWlYZCSEeJjgNIEyyrHEJ7LV67rzcY3D/yeNm+BIVGeBfEe3U
iMT7VoS/eGQnRGeGoSi8+zOQ5BaCcUPklVZe2ZDC2E92souIi7wU9q1IvLTm57A13ovLD9qpp4Cy
rpQA4KIfAztavRP6Wwlq3b1IflZQP5t1vAm7aHBoYTg19Xbl0UJmERpY6pI0Q9iIc7Rn7gwcczan
YfGnudw2pGIvt2WO8S5379a8scL/yA5IMjID060ZhPZUE2gsP+USSjbPDDHEHeCdWe0RN9SuDfyO
wpc3HnHtEuYfhfH9oy09xezgm66aZxXptB3PefDn+XlKTOX0O4LstBq3Xq7Bm5ue9qlJEr9zVhj0
g6+tTJ3dYnCoF0TAgrDsCtYgLcbSd4JEOoE6f6lUMcUrOXsjUIsH8os8sEifHH9B9mAQBKizUaAM
uKnLp1heCol45oKDUaRguCyyRKEXJqcq2mtsDYWbPQE29rdl/xOjPSMs4xTnSvxvkQvICljQfRKH
ZOzUJRo+kKLt3W7mq2xSaUhTbwWoASmZvNTf2g7FC1D++ndMMnCHmOX9GWbuIV4Wr0rbDJpwxtSA
3kPCV+Nwz1nnGgyfCx/VzjziDO1dcUNa3BQV8NXmTQlRRpOuUiYOJ3P0Z2g+l4ZZ1o7MQ9THsUbZ
ypQDdSq4GKJ83mJWG/K7VKuia8Z9bpvmkjxanc8ndhBqtUwq5BqlwF82oSQ/OT+mY6Ssv92HJy3/
UJXLgWdWs65cBBahSpesEpgMaMZ6xXSdk+J36KPLs1j+f+gWkl080xDqkbpFGNqRxzsTjjy414Ft
9QB5A2KE7f5x7UvKBgR+J7Bysi0sjP9AnXZ5h4ftDADMs1mgKaWtWmvT/qv8FBgbiCH+gH0k9ZHK
TIHrhVy29Cqet0A+zngGSr0xo6vkspZwpXt5TRb3yFiG35cDC4KB3sQb05jlABTITM6hh3T462XN
HPJSZG9vZYVRwPNCiexsyTMPo8s3qT/Pofk36fLxklxWCrOp/RSlT8wdsJTW9TDhtsnvel3SVAib
YbYyXTsD3TJxS6VKGw5BB5Neex7EGJZVMl1QcB2mj2vOEoJ9dFRF8FgC42Q75Yt9x9rSy9rWeHiP
9i35knhyxJshIFMiUcj29eGrK27ou7z62XLOg/Mb/WRPQLUgyIMPmXc/1TeD/4zhwM8JVI+EoIVk
9igdIdWmQTd3M/d25egiCnNJIM59LG5xCmsRVACqHL65AuClaL2dH9aght3U+VWE02vw/T1daIlb
0q0h2urNurcQ3RcrGk4Ms6Z7y6QjcwITzw9mU8WlqIv/H3Rard3XHbilRWPh5UyN4ObEg9dCjES5
t91TLiYnf1+6OH/L8ezmPOmIwx6EaoX2HeiKZ5n0WYB81J8JbCjj3BTRK+m8lKls4DhprGJm+U3p
24mLlmByI4XcAjn5FXB4BD098ADbBINcht3L715CldYGUP6JvY1d1C3doSkKmKcBAI+9KtZ5M82B
yFpVciRh8/OdSuo51lHcXCaBGWHrC1/ImmI3DgQYYNu43mhNBb4+aETbvBgrH7Han8K6dIJs6OGX
OIme7CLmXBA771BGomkggh7aidaEMzyejCA1fyxY6CD3WG0iWVqV6p8RWQjYYiwj0T/rEXZRKkbk
zqUC23f+518fCG2D9GbPyMnGY9Z2m4LQgVzKzjMUqINi6s7UXPCUs7E0ZwgKXIC7Zry6scSWr1FO
kVwh5ojG5a3c581v1VNckOwMEJYKo8br1IyMdTaRG+MWXP1WOwfiamveBjYWI2wv+zmDqNDH2tqI
x2VanFliHi1KBKco3MrlH4EhdXHpRIGM5gSbX2rsMWZfF5bCwjH/tiScp7RSx+L5EV25+GxXhzEH
ePXBGbv03vq3lJ9Rl7Ey51KyE79NSJv51lnHjvYxLgUUkU2o8szmvg8hSGwMZ4ivjEZLVaaHbF1z
2Dkk4/TRsB3yCGB0ZJykayDuxhvVLi1Xb2V+ZfQY05BLUobq1daYtMqmEuO5qkUqBm9bpgve68RS
To6KuRO7aKc/H59HnrlVomgq1oskVn5yc4xC8SgGisUMr2O6bKJ16ND4nQhsHILFBNZCvPbcOZ6t
ROCsbvatkq9leTdbjIZB35StG+jeBeAh2kNoqUWWzFX1q8m0VO2oid2bqkPiUgDGpc21p2t7mjbj
8lzx9uQNC/SKGi8KpqFttfgiTXPgQrcswZZZfEtEwNp1MdQpZizugezzoBnHJ5as6S0VZEu2eg7Z
Wop7LMr8aOud5JCqSGW/pXpqs3ZRMrwyniBENezrVZgH1fWQN/bHYkHFgkUotwg6DZcTT9KPIT2B
fGMo+b8RVqo9PvCYtB0KrB7933CKeeLST/Q7TfH3iKsBY4MtaF8JOqPJkFXAHWL8mbFnG5o3apLr
UA0seKLWAAMz4aE9Oo9GB6uUe06XAIr8FJOAsGTfJvxhgndQdgatBTbjcb1al9h0bt5gw0m7uHlJ
vcm1/uwlajgX5o+KCYMjPUGOkyx76KsFV+4E2SLzHh8Ccd/eXhl8DYtA9gOq8wxGRLx4RZVHgsJP
kEg+fASS0aIIoJ+2KCkhak2Op6oUYyhbyq/eNnHMn88C9JjXWI6406zLJDEFdKTCTjcezJeDVWHY
oDz33c+FC0rZwMs2ec2FqssIDQKqeXEuhLXAPKHY4IUrBHpfPS6MEr/xEZq2Ut2ZZ94HGNOOuqDv
Dv2W2Q2JRTJHTmOn85cLOk4yhZkRgQShzDR5UiVthXNuSERqmHLQlqdwFR8AfqAyjSnqXqvAxhGb
OZpvzIdaD5/vUzc37wtoqTfwLVTlO2SgE48Pv2v/jmNZquYl81X4SdEbxQdIqr1PYREQOXoHlUJG
fnk/MKEyTU02/a8ctZ1tTDJr7IM+l2AcbxTATYWAU4P86L4W2EQk5uLSwdpm6fBEYsZMf/BGAifx
V0RqYt8j2JqmnzZi5qyAZCAAcjJDxPFGkvB9oe3OikLNAFvXMMj28ACo8CRCAcaCNpxRjx9/Zszr
3l2CiDGlM+2Q4ng186y2uAB69D6mGyIg95cOjfVJzn6S3JC8mF0us5ngwcjnxkiAAzO3nZ4CYtTv
8+bnAyoVy5l+NaxnU4fkOJMZBY7WDMn7tgGYq2wbI+uxvq89lOJEP5SuvhS/XmgWyqJV3R2LC74H
5qPIby44wWuZwqbterONt7RMlx/1YOr2LfHjgevycyg6I8iMEaAwgrMO5zW4i+efZN1Xtyy9X1Lw
V9H3oMtFb8yNRLc/W1JjPXogEtdW7tC5E6VhQY8SffOhyqu8FRfoxbMiWEKm5Z9p1L/HaZAHm0Wo
cwVZC8AgfldBVXuFwocScSbT9a5Tfs0AoU1ClbPmFJHaw7GxdhNz4GyHLSbU8MX/4eloVb9eah8i
cYNIlDF84lOCvCha/xkP1a6r20CvLmhU8gADu9W1lyucUJG4WhcYVcKsWrisrflQzdaFjcitoav9
Fxp5QAGUNTenN75I1V3wxoZTVtAfYF/QWUyUYFLhoGdtOfQjcW/e56ut81T1EbvgbOLSSQqJEndP
uPspSPldzj4saSB8PBfPv2jwW191xExrsMoMk09LYFDTywwUfgJMIPRR/GjbsJFiuOb4qeDe+VCc
2nrk+UfqsmCWKyctDjzuUBsJsO1TgpcFiWAdW+ixrNODH3HMB/PrUN3tFlI1V6hjTiqqO1Gxlc3E
gkdHEYaVRDTcHn1TEZT6ClAnboHLNfZmmFoDRNKpp5x3kJlGz/9OVJr5t34SVP1d7b/+B/AMb34B
uwwYjPt3Bs0BPh0jWjomUlfD9iWMztepNEEQC2EVlDxcvCO7ZViMa5f8yYKWkQm9T0avi4Hc/RdJ
CQRbfKhEaLrCwMe0QCFgy4QAlHRSfrBCUzmTyMV+9/gJUbdBTtKy6ASROLEhjZB0sKiJkIcAyes5
2lr6BWJkdq50ngRbCEmxFro9iIPaf1JN9WNK3fpL14A0UHeTSDeG36nnfuCG5VaWgg01iDUEHea+
HiLTfybfaVmf4R0MwdPTluEGSR3bY9orAw+GZFIhYwHhlH3c3KNhxEFiafHdEG2Ml/cBp718qZ/M
5N6gcYDBeC/6zM59KR1US5xikSf8Yb06sSzJUH9mR5l5w0U6jmFakUhEwWrbwZyyHB3ZG193MzoX
niiegBnjuW70iiTdcl0grTjqC1kDz1KRaZt4SSgQwaE+lcW5EbvRXFl/jfh02ks6H79HF+6tUhnI
ZCi/lDuBd9pU0OMzDm68pQN4NEJdB+mz0Aa42MmfKhTMlZ0GWY6XzAlHDJLkEyfJfBfJ7dYQh95+
J4NusipXPP+f2Sd5QQ+dip3p1x7lDwmXgR6vRLCV+dHNcx6ODs0sHH8NsdlBZqy1ZkzXf3j58bsK
eHTAJohiM+V8n5OUnUp7e/FUDZhh0U9I3awTRv/87VKlMUDaWfUyhKRRbY7geZMhjwQcjmTuI9Fw
ep9caA/sUMG6zX2anSEViTTkNEeIW/eJFcoaCD4wJAWpi87Ua8SBWkOoPRK1ww64Oh+iyGmlzbIa
sEJQpyzMNrjwnoBv2wB/rZpOdIAk0Hy6o8XK/0q/nk43M6b4WGunWv6P6QA+h+HRyOho4g2Nmrha
MEpCIIDTPseqkwczbC8qN7p7adAEUbtffsXq9qhnqDj6yiTnFjNvlN3T9hmsAAgEYuB7qzorgLmR
PNhR/V/C5E2uUSs/QIOzUXA78bll6zkipwtOFSEPDUMt6SqHfTgwNvAs6bLSP21Ircj0mas5KYZ4
1uemCDtsd7eP6gq1OjHSbxFkFB5YPME6GbXzI7OxTu2/CVeCjEzUjOQc92rg1PwY0NJsfuVanJX+
6iUZTmI2GcKVfoLOJLbYbqPPamkMCo0qslRrBweIXHfo4CBBv3mey6XxZpuiytiX4MgyJ/rS/sde
5C0oXGrbIuwKf/W8v74IxWeprZVdtPIG3qBjTq065GM4L/hDihW49GaVyEKOFaMiUW79Sg1utTiY
ad20OVP4Ipm5u3JXP7ffdI0LeB+3zLWPIZWbnODRPhcysuNXWSzOXwDkV0bdK+CP6OGan1lneUdy
4+ZNW8Afiax31IYvvn3BgPxK3YL+4RbpL02uKPhi+DkOJPjWT63iTgp6fVng34qW++rF/WR7gE/9
kwEGTKiekaVxsjnsM3+mLjD64/SzUJlqhqgNjjs2m4TUOqnmxvf8GmRNB9D5sP0w37xK6nHg+VMv
BkFXlc1xhdhObXntL4NYfgQ+fp/k+P1eADsUAP8styl4JNDJySIDjg/bzQ/ZYCV/LrCPXauL2UTa
DghsrEWXVZ0Okfun8FJlzn49lfOeu7xAbsWLojrPPvwotvJUPSs0Br/P6jIQox+QI5v4F1VwJgZr
YzAm6aEfGP+x6HA0QrleGpIgJ/SzUi09J6s8fsYpXcY+LYKHHIWMuhFkU6zafxIgII1ARjnKH8pC
8YG/GAFMCCyXx0cS1hZmRVue1PsfjunMlmyzNw22yB2x6hpWd5wJgPH/qDwtQj+M/TGd4VmBFtwo
y+o3w9UFKqcV3+MppYAVOlk6MrxxGmiseyUGu5nODoa+Kb9Q9mtS8YktPQUrM6kaXhTBwqEOEn8z
JeUBJ6Lq4whQhpgZp6dzKM7f7n31Hq2CW6aYOtL64x5po/saWNOd4rtiLtq89In7LB8TyH5f5nfm
pKGeq7CD7/yHbUgZqZ8KFA6CeBkyrtvCfYec7uWwxCzA8WMzDrDxEOz4TRTYh9gmg5rYbYXbvZs0
i4QlbnmvuSN8sNUm0wht3srd2H0LviNYBvO/1WXcS2lj3xucfP+Jh4VrC5ui9gIhtHUYpQm2+QtT
zI82SPOvoJ1JY5IPovaZtEwdkWrodYrtB8yAo3sIBekJ/fkhMhfrbh9aQLk26OqSW7aAidSlWeqp
YPADIpEkR2lcTTHmf9JLsqID17HEkqBT6kdepWar9XB8E26s2yAxx62KizaHRJwW/wdKbClA7BfU
u9PRklcCZ5y7R0RgOttI2EpCTxnqIDZZRjHOJ3zvSfdjmzK6fDZOPfQWuDjI/J+Xf667emKrHE9b
I/oQwkLrGGrlApocTH2bEsJkx9R9RM1YLYpx0VrLkSjYSwhugFuORhKm15drjvO53qQc3NyrRxjp
X0qH1nH5Dvjca8Ala0Gzcz5iiYFIqa4BenaVeo57Ljfsyycy1aGPakFH70qcQysdj2Yf6OFocW1r
VnBQZdoeYxfxso7wOFJtvkip4LZBZnYNZabQvrwoHqQ0EMCmWRL6SArez6marKB7ZMyKKXjFqlXY
eb/4MtNG5j+MTDcgAXGCmfxP0xnX6z6zzbI8P2R4YiIxyMEz1Sb4B65LdC2QymAyFKm5/qjBAnt2
01RGH1b52UnKYBs0leDSQNPaqvmEIX4UFfjEqQ7huQxvP3WE101Ly6l66W3hd02ORQ6m01EZMizE
3hSazp9E0ztQH1YuBkm6qKjtg71L/aYuOGwTPPx8uSlJLU9+uYvVLbsr43kV1TOFBBcNTVKOyeFl
MOMtdXjwCthaSFmWjG85cz/7OLQ/bKSNO8ulbcx8gKVmYPTA8F/5TepxDKmiwtdR8ioNU26aZ42p
gBAg09XzA0Ec7ykKA8zY7qHiQuL1hdX9BtZ7lEGuTfpQuo1j2kIrubT7Ha9s4IL5JpJhPDpgHI3C
vooubFaTSR+zVqt8drW+G+OFPXuvV86RJLwkyyyIE4jHWYjJzdPVoUrqqQyIjFvE0b/X6HCeOJPJ
HCgOSmh6RGP/eHMtyyXfgUncqH869T6mLaJKfcqyxW11S8uDrH9DfWpilLy1GKgRQu33AU5KbKAy
gg+yq9dxR4IYAjU3/6WKqggtyCzT8MxxAyCmmjPv1IfOwAw0HqLR5VltKcdKlbmuXeSZnLjgmJwA
geOjUBldCTB6zuRa7IQuDB1+OSfRsRw1juU2eXq1P9xg6JfAFSQH5yn1uQ4cZBfmsEms2lcTcW1e
tYP3qM0WOOWP1tGzzBtHvhtjJat+AO8IEvVoxdaiiY7Rb2TxdeKYu97PrKpOpWBDt0h1yQXpfQm0
JsbhLSR86IRuWmbotTMwEUUXnXP8BN6aT6CUgGGQn/vEljRw8glZiU8Uzo+/BKDexh/Nfn4TRE5A
1pOl6cdkJVPLUWHxBE9EOMaD+RFx6Uy76LemLtuTxBUFyIStdZEOUOue19n/zk12yH9WuSLAnLaF
zbDT6fzTZIZsCKPGo5FZQNU1AJt18+yJpesph4jnHDNF/m7nk1FXyb6Df8+hkh4K/HG7RckRUL2E
2ynJEePUjzhiwGOIuO1Da+CI9XSn+bxxm+kodGiwi8IGYKZM0qzsGqE7JEhFWLt2toe+yp9a1pBv
6zz4QCl6xIOqtc4EYhapJgWIFB/gJsS/wtaCeRUeC2v5zDg7r5c4U2DIsa1UaVFS+jU6fCLNHJ1d
acGMZEAhg27w5fpyfoeLA7T3G+v+hJVBpg3XWbxuFkb7WuiUh0y4v3bI2GgvuuNtzYPfhHHznpJ6
tafkvhZ9SLbXcjfIrByfc1OcaQZU/s7tEjMoG3eUr7ah0iUPkGpgjDw7Qv475kzL9BHBLCNHptiQ
uh5biMx0Zexx+rcRkc2kGj0gl24FjcZ6/r4nMYGembOY2HNMmXZdJ9dyK6pRwW8xK8B+erpnRI8N
r/2VaGL1WVJsmRWmsWZymes8lYRmEXWdLaGI8bHvNMS7XxhuNLnR49ihOJ0uYBag7m27kQbaQzf6
ObZNvp5zEb/mMTvTUs+K7wdiZ3CgAq4nKRQVOOQXU8X0HIYuSMRUH85PYMm97Km7CqHfQK080V+X
igwi+vrvcTXOHIhH0LKQbY86IhRBF2iPDlVOKcCBmk5lqyhXrfSy63t5hNoW8nWhz3lT4jAV0/Fv
M55sNpt4GIxoWlHnIeSeUgbvnquNgWH7fId5kmLaDrkUw8Pv3j3C+2eH1FpXX4KwWUwYZ6R1lrIJ
n1gaYPmQULUHCNUwTFkaWDoTQ+jwmwVlRaEFQl5P8dzqCdra2ZaiAZX+gZHaklDRYxfr3rK4vwA7
RornmpDiLHrt0FxY4QWngggI5+9XV6Ln6jEVfPKetFbty6pqU7N6wlwdnxHTBa5pL0RlspzDTtCr
x1PJI81the8M4yFKpp0VH0qA+NcnPMrrinPdoyvMv349Y9UChTwmjHo5wqNPKi5UR8M6vQhbNdGm
Ovmb+O+qIUzBm5zFnxqnMNMEx8btVs53a82hZowAHJ93y7UMWlIzTBovioJGZJ9cw+3XfQRXw76I
veE8k5FqBKHM+qVrFZm5KN/O5XQFzwe+h9cNyms5qSUQTxqeHkndEAVnky4nvAydPv8OGhu90Mqu
/1v5rlfnudI4j5V1BM3fTUsQ0v5ebP6LB+5X+WvQHg9hafwKU+l9T8l2rdLuAi4ffFGiQYdRTx7U
ORHbdWep4TZML7qJwMqt5zh0FFMcwus8VsLUnE6p2rpWZk6j6Qezj6qmR1Ld8rFJw/VLqkhqkZmr
1BPUkB6QoL3d8FdZRpOdqwDKwJ6venidjvLBqhARrcS8Hqw4aLzR+mmVOTef85E71bIUkayO976r
WTNZki9ni2eRDmBtVbM1w7x69S/6PlcPgoHgHSXyvtUHbMKYismrMTD2XtGuHOoBCT4cCtGJV9kU
6VIX4+1d8YUoSLJ81u/QmyXPj5v3v6ZgFokpRDwabKXB+PiIQLrHBBEh/sxX/bIsN/yqNzhg67yE
O2i1Vcp+9q4EI15V8OznjfSw1rsJdVZnkzfHk5Rn8JKmNyq24ReVpdQvVMPO5RqEAL/MOoe5fRV5
JUox18bATQhNPl2ownu9bBucTTW05iIBfvQ7t0AuJmcKKYB6zfEpKfWnQXSzW2qvsexmTN7RqDWx
3oOLauxh/L/PUTVkEiYmUshwi5QHBXNYAB1c43X83kN3Vofod+mscpw3i4yP55cpopsGeOHmFOFN
OkpP4GnmMQ2laslDXPYaAPb+H4E2VNlzHuxbfqxdnhs5h10I1w4joX/K1Bxd++MjB9DLXFPP448F
OlSzJ+6LHVrZnzJ0yq7zcQhmo3gjOshPS+OqwxcvlTripTYVpb2UAx4NzeNk8PMSFjmUe5b7Y9R4
oiYGiSRLWEsKfd2RrZE8lDb65388MX3wFb333kIY4iy04N7rLXlVgl9t/0Ow4EI7+NYMbEIejgW4
qjd6D3hc5il5WZzUCxbveUTez433gMHnkha/H/+X5do4pkWYq6A++HZowMA8EV9TDn6MUaB1MUwq
+aJzldxOvvOFHOfazYzxEMvdYq9K9F35COiYxIaB7AO48ANteXw8LKVWQ/7kxXf6b/cAnW9RxUId
wiJAiPLlXNgFC+zj+mnrm+DORzVOV756fqUURMDEKAKaZV4hTVQU3QZSVoIEZVJZ9unnRNiqPE5H
UIpID18ISVj7ManQ1d+vWw20ixoej69fqBUdG/94gk83IifMJQQUzoFtljAZp/zuBrZGM+IDDqZk
m5wXPsCWPc6PCt2Td1MUFJh1oye8gpw8xunreZeoZB4El78kKtDdVLbKd4h/DnIMIdvw8nBby6mT
AELsGsMjau1O9qdd5sl/HP3k0zNEKjd1KTHvdkTqEnRjyUFil107HMASZwJEt0SMUKXyTnlZsWzr
nYFGklQ7JP7jJkwjYaIzw+wBrpwyL7Vwldvhqe1Pw0KO6Mne2P3ZKKwc1+6llFv4fFVxM+GLNQLg
XGTsG2xcCSjB/H5eAVF6pUJcz4b8yUwFks1MyqImys264IAvsT9AlUtEWQl4Aa9adIpYpHCTtLki
xefd8XkIK7Muof4smUL1dVlBJ7vZAjHcGmlRWCmEvirEYcmWp60WfkUuwLFDo21HCUhDYKTrUgY+
FF7Cp5RA34dYmfDYmZAkKpI3mVZH9SAXOBOkONblHm7ZeKD1bpW8nHKA1YRl6TUECdd3+3i8rmVa
IBcY3N2f3Nn3kJTmjiDS5arxyDRwZFgS5E2893omRUZk7X+V+FHcHk9A/EPNEuL0Lu3nYU95H+rN
/MeyRVDYQ0PjT+3ULN4ECWLvWVLJZq26LuassF3mHVsTqmwuYLytsm1zl/LAoxm4bRuA5l8mU7or
/4IcOYtNndauXQIWOh9Ya+hxNILbltaIkiLROCdNGUj/yzKUcSW+h6Qa5gyWKxx7a/HVmqc44l5r
qTV58LNcqEN+yJLtuDkX7pP5spl41m/3blAu/7cTAl2hMT5j6ayfP6LE4ZeLyQwHu2/Py/PsOhc+
BcZgEKNvBJXrBCs+RzoJNqQas2ofvJ3eiInLYX+UQETLEj2s27jMeko0AaZ8GNoK3xXZMmXpHjqd
fy24XDeI0/P+JsaNzS7fT2EznTL7lqmzQjLlDyUsq8X1MQk7kGj8bc0rWxM3Cm3ycltCCrHxTU8m
gPl2s9HH6BLA0rEKmVFaKOqnvLtPt/oXoH09qt6lAyLSfkMf5Q3Cf+ms9vSwpSJsFqzZdrlUH97c
Xo9+O6qeVVlbysgiCXtcZyBMk34XIdFpbLXwiKw3Gnf19kp8+e39R/nTnNA/OwMmeKbTAuKHl+qi
aVM3aqsCsEHqe1hlCySQYrjOPKaQ/JVtCVvGz5ttpLDJr03KRfWTizf3PDyPVH3ECXi9iQkig4Al
znCzTQwPg8lTUZ/iP+wPana5/QiTGQqgLNIileie0gY8+V9ODds3S3NxFctIRHde0xMCTf/zb2vt
vmYWN1s+H2/8DivvQz5XRE4VJUXLw5LD18ySYbO8vqEcuUFubErjjwj7KamehsQdt/dcB+5iLneJ
Yb7/G98zZkex+eWMMwxx7S6dGh3dLoNuRF/WZ2isY1ARsuXll6WB+ShACjOpuG1l+vcQsnuljvaA
USYcX0t23nxlWu9xAwNAuonvVumA0vK9SR8UOglnT99xeyA5hAfUJwuVQl+a2Xt48bXRwtFIJIAS
4qSVVcZb7LQhyBKLBGSON7ril0FwUMUqgXT8/q/pDXhcDWMbEFeGYIVpK7NZBq81qmEP3IGriEPm
6IFUmInWZHXAB5crWJe33DJMZZN5Vi3QjuzXlvJINbhRACqx7R9MFH28/0XMA0QUC4IBr5xrbKws
IufXGSZ/5I8BpgLEm5iMffeL/15s6Qow9yCEhWMG92XLMUsVu+SID62nBm3VBjjpoXLFkJkwk6Bk
yBueKXXioZHh13tkovyx8Ha56rdy8unoETyKfyq5Es4qTWFIXhxnM7Y9QVu2YHF5TEWQhan0/e2H
I/XIEb2n0wG5qgQem9vyJr7ldwh92giqBJE+Uc3yK31aCa5REelKS8aoxmQZpV5ehw6ek4pmiKlV
id4iKFU5IF1hZh4rsUmf1tgVOhIv6gujTfJLrs1BRCQ9rnjFMKCRpkpa/qJo9/793oFIeNJSrkkJ
s7/kgX9kQ0v3oH6rB+ZwxRZN3pfisgb57wc7Qofn9MZSVkV8I+BqrEhlfpPDElj8wAEwILbpWKFx
I2c4vJm+HkAbKdtfBPhropEbVHyjQNmcaUTdXuVUj2SVvTAGjJakYoh1XRxaoLFZnjXNwHbUHSi4
oCWpMlt1qCpNSMoKGST49H7QX/zTMY76NOOt9uThcY2TIsd5BxA8ojGrtrRw7bi4tuHF+loX+7G1
S3ZuNvy9yZHJj/CAOz7ksyDfTU2vrslKcE0SItbk48mrpZHZAGxZiKo8WxtMSzBWgt17DLHuvu9h
ArcjiAxHI/a+VfqwUJibBqgJsb9pcV9U0gAoMJ0su5iIBjsL1KEsx0jT4A1e7/Oj/ZtAmLdjK72F
cCkSSmglZY38MxuBUuXJTYjluXvj2PiYqO49+9PflqA/N7cBzgKP0lJ/lSFV/QJdcjKH+3mIG0CG
/oSFqQlQ5z6TBEpviIDd5mA3bElI7x72YuqNl+MqkLtsb4AtENkRksHMI6o7+yPuRwwGgQN3YtqL
4EKwr/1C2L3Yb12S/SCUxV/5IhToZ57Hb9TQdQT1KJIoNQyL4qE3r0URE4MZVGvDLkAHsyyLIKdy
T8AG5wLzBKYKvBkKFDaPsPZXnaMhMUpdJMOidHeD1iSSI8Lu4izOqY/RIB5e0f/dxnQ17WXkwYjp
v4JOpMM3y72j6DzMXPrBZGEsQAXmisiPuIaEqqGcjrxzhhKLWhWNTVOcvU6s1o3yuggfCl1Yjcq3
zr+jwZ3DFKXWf6oFpOZ4y4lVYQFOxxqXCYkkOVTOd5d1jEcr6JnhHJyAL9nN0Ye0Dg6EeD5YREsh
C+pgJM+1+K8Kjd2fN5YPQNWrccVzztifOkid8Ywd7R4tQvFxf8AcnThJHY0nnCyNgeDqCOioa/NM
f+NQpMMqQSI6nPoR5RetHyAet0Xq811QDc0q01dsyZQODevgWBKaFzWXscrGNRs0OMauwNKu+vym
8kxCPWrM0jUdxgY9gpVWkLA56JpsXHWhWH0eQB0wncDug2cwBDC9Jt7aFDpNXrQa1K8TiPxhnh7F
YRmdH4dtF2uYkO8o/ccCsUrm85/jDFEfbLWlXt37XeVqa+hlCdhdsQ/N40buUfjNDbKBdhCRoLcs
XO4F+9c2T+HoC8aGzb/etwn0kqTWv1E9Eq5N9TDjE6aa7WIRl3ALJlN+1GFAEn3ZTNdgvdyQ5puf
TMjJS9xGuMrHWY9OJHfj7RinV5bUOOB/Qz32xjeBuQRwQalXMvpJ0SDab8tswjZ3PJjKadxe2Kiz
8f8SXdm2h+KG/YvSG73lQeGBW25HlEyw//tWTO3i6qWw0Cug3dQSmxf12SZgshXfz0SDj5YF1UlO
B1IgBGOYvhJ/cOA1Vo4Ld/TMKvI3UMqfg/XHDsKp4Vmedz3evx5iHyCEL9pG7d1q+A4eXd0t2eRx
2XhH/KNCjDdJ8XeoMRXa4/cO7FG4YWaCow4mZSu7RT6VxIsbUti02NDWM5ASXPCEk5DPZqT6of6Z
efL8kmVDzAq4iWiIJ/sa6cdEfoCwL68S+rSf5/cQ1LUfFDuwPTqWVtpEMT4mQiBkzjBk79jbBJ7x
p3TgV2lo5t2dWG+wyWcLTYZ8QGdmgZWjVUrqcU6zTyJk7QzI4QRKBcDyDat56S21a9HEf/tiOnCH
hGnPf6kZDNZWmhyhf/GM40JnqV0wAUSZ7/pXQSbFv1iJ8XhJ+uPdn62z6qa/SAbQyJNnSbrwF5n2
XsB7GaPQeVQDMrlJMiY+NcDWytzQYczdePqkMLT4iyBI9zy3znuyPl6Ng/lvmYGz8vTW0XgqVHhM
1PNJFGni8y0YCOXSIDf+gG1YtxM9VmNnE2zj2AKmFDOLfhp89r0XGCNkAXLZkTSXqOTqLd4L4tf3
sxrErHpRhHqdIicBTOd1Olp+YHtZmIdpg5p6tpChpsonHChAMX9K2ImUMJ8uhoM1zSD/QJSYAWhS
xIpSpfe99OrWRmtM1TiYO1DrYCRAHWA95V/Uu5quLF2/KelK0NgNbS2UqDU78BQvSVGffYFwxvzN
odrLjjXqMreMIOecCeMQr14oGcx+QT8877mpV36VUPc5U9nY+Xfvh7dqGApPc/4hnVHuZszwjI5J
6c8O/9tyv+dmrtcG0stLKcr5bJoN5dtoDPkTuZoUZ0gBcvJEbGNZyZIF7TFfLou3wjf2fn+EuEi0
bIiOyepHSIcqH0Rw7AXaASuvGXihB0emBbnNOrOZ24hVVSjfLJZgG00vPVdm+SkuxvRsmFeVSSyR
iNZQzY3HTe7ccGM6AOMthkxXW8aK8irrs67L/Pe7LEC5AbgMBKrVlkHYsbYBnW9X4MwYTdvEWI+M
WjGyCIhBLEkTOCV0M8Pj+1lHcxLnxsONMYqnVeuObDzUTwrbKtfJTceodoh7/QjEdqGBSGu8L6Jf
iXperKCbz+W0BjWrYH9ddkZvnqR0aU6Rifg0xkjUvn2ZZKs9dYWSuDC4a3nCTFMinrp8n/0aw2I3
og/HqKyp4A0cKi/QD/tndPBEhKlirwxc7HNcQW1YNxrut9t0Ia3YUoEvKpOlVlX9hiPvioRxYIEx
u42ikLwZIdoX1KQie4VyXhYgx3M7wcWuRxj/7ZaI8KTAlz6LFLtJm78ny10uG5VfSpWgM/mQcuja
+J9TvDf7NNU/WeBSAp6u/Z8GXvKBPJVNzozVX+wlcjPN1YilcFEvL6Qx2fILLyK1sjOy+AGhultb
f8PXkpu/AxG/bV5K3Y7/kIt/thP7PjxBFVUrjCmPuvBa/sN1ZPrlwY4qThrQNIEyZxQpVvpt0JUH
zUD+N+gKHh61KUrSpimVD5cTQTRsz0/wKOn1BXgdc5Dm0Fb97Cd1ycYmictP9UZ9QZc4p9eW60i0
Mky1Nii/yKONx94idgNuakownVbvXvErdiUrDhz+E2K0RDvT54lS1JYKIgVBfnL5G0wqrrmz+fpV
EKub+y/vTFOcuYLgZy+/hYWZ5dPYG0MN6RWg7nd4Z7gZJP8QTqb/fa4iWBkDNGGZvfFYN4NIL6IV
ZHzvwwEkwYWp/7C2BLMEOCbkETCxzyouCoV54HfcXHK4EIwhP3DAq2Hk7b+56IfAgimwBMoRz03K
4JDDOWHJAOwLP22mB7f3/26r9ofxqb9tXr8ICUl0hI2lGMxfNAkPCkrRcBP4EshffV4KxPYgIHNn
6nOLZSrKGnzOlgCuEhWguPbAF/9UsZkRNexVyBs4NTF+eZ/cs5sPd8hXRqrGdNGaRGulwCPVaMoI
QRJFO1oKg2ZCnQxDguBUcPmoBiOPxPA4U5GBVEbSOKFzd8LaBOjvilBzONFckxtZR5tP3rCC3usY
jaZzHSRYPuk24U6TLr22R6s4+VucOt3FcF/l86JX2SHSnZCffr4H1u8vGAzUbu26IDRr6iJ3s+9H
NbHycbTXw/nkVEVX1v0UXtIKSJZo2pym4VVRKCiOee7pRRrP1hdfU3HvPOgiJiy2fEUTdI6XL+cP
zZJYu6jJSRCnW6oSJ7ZB185M8mIZE187/THRCGfSLz0lcoQ8cxX4CWW6vD035NnMhY7UOE/77JS3
+DLc13+QP68DaVl6NfwBU9hVqQlckj/Dkdw6s2FJ5Y5SdixMq0W+zUcdiH9bn5KCHkPNPep6d46q
hGwpUD3prKfNJ7gU3KYpfEx2XOUUpcLIkZRi6yWmAiQddAN2FyB77h18R/IBv7FkxAjwatwQ+qwR
/PoeWps5HpnZrXeEStMcYNuZTMLbOw7kNmsuZqXHWJ0gnZ7S4yaxam53I/HxhqoXdtm6IbV7YpGO
cKPf1xf60eDncxRsYwySr94btwUR7aMsMWMMTTXtqDb44tz+pm64NTmJaSJzhb9Vh42oib+uTtMU
qGDg9DMft9STf59QY89MPCRQ1JYS5HbgPh00WHvloKG2VuY8HnxKXF/hf+wk7iwA3A3G8VlJ8DRn
y/WLKF3w7LczN44YTT6dYEJi/MxqFnRoLIF6OI1EOaYI38DvFE32PcF0C8nt7Q3Zd3vbmH7IXOH2
LKSVsWE/cayNAyuF0h4adc+RhOU4iF1F5cshYze3+ONAcHRA6r9J0Dg3Gqoin81Nov6+CUojzJZ5
Xtjw8doisK28gtoAjXPnjTKxuc7y8nEh5PXfAnuoEHGylOMfvgNJWiFzss8I1g4Ar6TyK6WqwjrH
MbsD8z26Q7nV3GDCKwjQn7gTjen7DTFuPJ7rgS1uS8empa0t8nGGJf1PqzpnAyTUpYF4LwptxEhv
1atmJx8p+trIMlVjcoGEmCOJsyYLot50RDUDGqdAMF/WZW9nviqpzwegI0RixCwTylyW57XMWVAS
JQ/nM43q6Dt357Q50AjTYTUWATThBtRwHOA+NkVo8fFlDOBCFywTiMRVvNchXDqkAFXrtjss6jr5
oKtu1IAvxpj/PRnl93b19u5oX2N4y7EF0qegrW2RLCPVNUGuW0YG8IWWk6hxJwwj06h4HkcoN3by
Fg9KjjaCXpRLdphDN4RcgcDKOt+0fln2AyngSMfWYC3j1TyXOm8EtKJaYBgCI0KYeIdVMqim3Fp7
VxOn5VNxvIm1weAAxYTOVOHiGk2u9EIOaftBWR2wgJBmw0sCa5rOMBrN7QNQfRxWdFcq1DdR/ZmT
yr1FQDe3s/+Zr/+s7asnrrS9s+7qOKHDCOsWqFAMfN73F6Q1DGxfwLhhblJoYc8YfbMcDJ33fIDp
XrKQt3kCnQQAbRrdUypaRR/G5Fy+33NC2SXadpB5JqRSCRA2K6bAn7WFjlMGs7DAXnm1a6BrY9c7
wAL4urlU4n4l0joBsaMCsivdUpgCk/EqLHp7XfY7lCWkcQ53L7S/S1514yTnFiL5LP3ERUTqvf77
FhtjugXxQfJoMxuQEZcJgymCqDYysBoMStz94HmLN7IjK2g6CSDM0hPyRzBcoagCiw29zkpOJlPm
bXxMsEpDGiqO/lzcbB2+f+1tX20UlJt7MPGP6JvUomoiJO/ad3+jwo3XJ87L+18f3ScTJZZwimhj
3vbymbGXK2fRk3nZgwLAVLC7ZL4iyWiTWsoA1tf+4KHzgrF/L1djEMvi7gVbHffnu/iR9mFTi4x2
98R9wiCpzKFpP/zoHqgXZicaQfP+z1n4wzA4ExBCBvWWahx7AGAbgGWzD9yZZPhAjkxPS5DxkqVV
nGnWTV7YUvmS+ozW/x9aFqtBZgaya/KjEzqTWM8BLhII8N/4MV8ZmasTAkdjRT9zxs9qqpbgNI8H
ynLBfbpSmCLhpBR0oE5Omf3PXzXRQrZvHMhOhfO+vZrHJKWR8bDdfmQbgURvyMozdje3HU/LASQo
QodVNKp2+nRi1/kuEp1/wd8/IkFueSufASbX3WYtPcBagoZhRFR/q14g8s/48Nl26izMWQfs+M1C
Wvj6ZJsmVHpzszT3mqPH3p9j48OJyrj+dLeoGaN+GshHKBhzjxnRZs/uLrFsrQfV4reZdqndvf15
xJ7JLDDtblMrfGIpV5a96t4FZnna0V3acgM7wJy2TTDk8CzrDZVAhgF3umiP9HMGBwyxZCEwGl1K
Ks1D6fH39phgePcTQeNucHu2ZP7ITDg1zAF0XCGES1rndhgperU1XieIfeLRR31DhmTkcnFbUaWO
MLF3FhpVAchd0P/jnGTATF67TC6ucWjU6jMMzHmjhRLQv7HvqFzi+ZVzhd9sAqcfaTS/W5Hju2xw
pHu79hVD7MReNK1dPgHTdEz80L0+lNBxTQh9NOSTE63oNULRRbwatiJPvlhfGD9AAauYeWajE4r9
90wkrR3bFj0a1Se/DG0Nf3NAIgw8DQv1dnbxaME6bfVdJtpr00eFKQl4LZszQ5PKfNHhHgM57AJ4
T8xJog/pQOILs1iDA2qcVXRaizZIBjlz6L5E53zQxZyuEcgANqGtvk91AIeQ1YveIJ82ZHitHSEi
Cj0oCuISD7LhFaxX8g9aFaHQbrbcc5uCb/E1hRUhmlbRWGl59rRdf5soHSsKesb5n86bl2zsCN+M
ZfuP5igHMePtz/Yq52nnLW+NY261lNhgmHjUmue1jfs6qR96i7exHcUMdoS0H1nGQf7tB6SFsjcu
VYKYJv6Y3kAi1A2C1SxBCQ+/ywYAEuXqoZo3DdMV3zD1vUAEX6WMyjBRi+6ewkspV0KDN88TFa5S
Tg9jx6Oic0ewdvJdFjHHl9Fh3M3HgEhAfvwx/SaadvTZMmRMDmZyhw971sHfNq+52jvC3qohpmRM
fgmGEQD4w8hZ3DSzqO1grL49is04Mf+2f6/zclrrOgF1mwO8neN0/r3XF8DvWw1dqZRS9gt3SG+h
oMOMdIdKGI5/4qkwQOSLphXa1zIr+6G2tIyD0La4II9Bv7w0KXgnZdv4uTa8Zwsy3SJQ5Mzwgapo
C4YZc/eT1mUrjY5GZNs2Wx8ulxVbhYpsqxQxDbVFEu90Gu7Vq9cabuxCZ/mnVtb6CXPUrk3p6XpQ
pNClVrb5KuD2XlMlVhcayBE8QWBlq5dNBdTu1LlOF7fadCTNIHz8wvCDihMWA2PRtoZI2VKuAJ0y
x4Qwzd1uHX/GWRu4wpcpIgqxjekxASk5nl1M3Z09neszU3HKQkMUQX9Mr/d0GTsQm37uSsgkRfox
cJ5tM1hlsF+EkOB5q5SPElGEgaFBtP7n82dQV67/Le6keMU8Dp9IPD1+WGoQWMmOM80EiDkVRont
VpJ/CIckEVeRj9Rdo9SJtK00lV/HQRd1TSFVVXFw6QiyHIRbQ6VGIMWHM5Uw4NFb9CsOqe7NV5qP
85/tKH0r6wuOoSr8OzAyA80H/hOfaWj8xtiTJT68aaY1dFuNNULlEShLf5FA9t3RxddQcz89A1hp
HWg9dn7e6YJ+aaQLBzLylOUl0l3LjeEAOu6c9cnLvj0Y9zcpegO/oemXD6xB2sKq9qwhsxo75EJY
gUGyt+JuZ54wzQjx1i+kSnza2VsJXEoBPJcQyaqoswOwA6tx4qtO91eBzml55cSUNt/1DA5xt9HS
63zpGgl14dfo6Vxuvso6Xxnhs9kUpUXw9POy8aLugzWFlu0ohAG4ym0IamYQdWURV8tubUXP1Ve3
TepqCM62+k4lj1QePx99k+7jR6r+p03CqyetAamR+NPGt8TnJ1rBNYP2yQ8Nf7Wi6FTRRv5YVajf
kXMzLoXCAjgA3hQrt4HOFjgsuRYAKZWlNkR++x6+70WE45B1weJcrl1ThuhvAQv9h5bWSxagU5Eg
Nt/Xj9efO1/+6fEpbWNWfUjz+gdDzSWCLXu45nIl3yigs/95LNnlG+CTo7Cdn1lbroJ7jgGKQTiL
USs1jYpChZTo8WTzQ1OPoG+G1JcjJpjMM6FLM9cjupdiC8ffbewKhsLOl+likcywcrcI/BAoz9L8
tUI7BqGLHYksg1ytig0wZYl1PMF1BTnWUic1MSl1ib1fZqns5gSOpsCCFKvhCquK4a5eRmWMZkTs
OcmhBOX3fd4FbwaMoBi8yc7xp5sH5Dq3vlXeTzoK/2nvWyFZQueM/zEavq/1tjgPqVk3JVkGigZ9
ulBdNEddBqrfC4d2DipoDgABLk4KR2XPckNfVXsQOn7zz+4ITvKb7XbtD/obc+kSzi++iCiXvuQe
sNf4koArpbhS4nRt1ZEQcwRBohP6I11i60+HXNJ+YyMwKqFFwdGdUyyzc1kC+OmgDJ0o45cCloFn
N/Iwylz41nFJ5P/3dPYqPBkqmA6fdNixMv2SExIIdHEHaMCOf28Bk1hPGRuzIcQWJv3Qoo0fPtbj
Q6hIGr+5DctEen0zrWai41tE8Xw8w3OMudQqoT42AnlHaRaCmecOPPxv8yMLzMnWHeCq9/S98Rg0
LKJ6pLw1EKEogjX9138NBDS6rBAbW5cOhkmAxxDnVop+gkUWGiF6Ag7Yn0JjUQsQCKbyPm9hfse0
/yVOjZhWrbMUyoI9Y86vh25J3UR/rKUut1S/oRgokbBUXmjEi3/CbSKtG7QJOVhVF85fvg01O0RC
ljngg6axbdEuLyGMBtDWgvoYltZpEq6SzDy6wpiGu3teImIVGFxIQibNNP8Am0pmhHJ8ytS/4Lz7
Bi6hnu3t5liFhd5VQyaX1GzhvkKkrFByqDmNzMe+CdCaa5+id5TxB+BBZh5NFSsE34lWUPWjcp/9
9k6N+/V1JyKzDCf+kROvofH2iOIQhpa8s4s381TLX2Z90eLgTAZREDM7JCnEl7N3mXwH1iX27ETK
c8LaFUZK/vkGbDYf3xU95Qz7/2/R+q+MqlLucpBUJAd8wKQgD3kBF+Mvg1CcWTstqmKFavHoF+sj
ikKX1XeygPfX2H3nl+cY/RvG2MI25yEE5z/sSk+pXrbP0X92Xqtymqpb4aogabhLOMLKacjn12sb
57fhJVp/+n1AX6RGezKeMx0lVzr7lQimm1t7sy7y8rXQ8bOrbtqv+8StNijBO80QdKB+zVtmJfdT
vyL5ip8D1KHXaJhbOPKx7gNVa63lgcQ78TfMj6cxMVl+D8tRcpcqDzeV21voK0nEarCG3laaSIGW
KSWg8ByQmSxlrl7VadARByItpoJ8UBk5TzRMeUm+yARs9MV3xdqo2dzt5J6LCKYRa1MMY3HK7Pni
PyGch5uxUZHYPN1X9SDe4SlXjWXWWwuRscrNJF5wzmMjxj4WaoQK9tThajPjawE8GLPh3wm0DJCl
TqG2ESLsaEUn+xYvj/nNzde1HTAF1RZ+aOtARJrcYYizMM7lpyQC1IGJaz2qbVIBGs0jbBzC2UM/
Ddx1tGBJ9vPfQXsnePxHfhbxybBDsfyf3DUco/YYnUwbDDfovftSxokrpZjww35SldD9asBbgScH
J2Nx2nccl6cLEd8IDMW46j6/h7l2J2AOnAj4q2Tx2HeZlyUWUKcskygDrhsvFB++r2feQiVWdfqR
XKPqdNTTIP0S1vCWgjO7o0S++5Y403h+polantUm+HS4zLHV+vCWTY19lScW7D/ISKFKvS4b2OWN
hS2nqS4XEUrOA6vnp1x5L3BFkkRCYVd9ZdkBWz9I7chtcpvilY4q+JvI6MNHZtvIfrBubLPpA7g5
BVtGoFJ3iXYFpEjh/JN3MbWrKhhewAsgYikNrVy5rtYRSfD5rvkz6Vyf0curCJCXNcJPKm5uqPe+
gCtmqoNPk2bN4U0NObHipIlxsJweXp6ep598XFLsArZjW7fIRP02S9cV0Jk2hC3uNZ68BKf3GwCP
4zo5Nq+PJLmYy4f877zCxx/8udbs12SjOixPGcyKmQFbOOaGJJ3wPSBoW7qztb6fNYu66qmA7kpL
upOoHtU4ny7D1D3fm+eUTR1xREeDNzbJ3Lqgspn9YxMvTPbM5mwM+Q6s2hM4AndKrGCMMuW4QZFo
/mmCXUOlmFG2oYAgacU5F/+4PuEIXcVNUdrcEZW0I9r263miPKvwbpMs3hS51vRwecAcW1zCF7vy
nen/dnhgQb2uJE2FQ5eUB4iulu+6p446W9rfdW3Z8yNLRHKZSfcwMCsdAAJvAXN/ejep9GCC5Adz
jGTq6wAxdMlgpJ+HRiR0/xn7MdUUXsn6rUvYO6UKJdjLc60HSTEPR+RXyVghyWFB0Aex+1sgT4ui
iM/ZUkBekQvt28yyIu7WlObMlx/N41jzvEh7a3gVjXDNDb26c0eV9NQL3tuha3SamlW+/alqkl1M
FOv57PQfcs3VMiKPE9OkJcJE194+OH+U3IzYd9obbLx7kCAqa/EGMHdzTzGN7IIjTmMDfu49bA0f
ntjSsbEqp5kA0UQ4chwFF1tzVm0fMWTcBfhUsGghxrZxiYYWz+BOwipY7jOYxI+ATendmvW2vLRv
sjCX9O5dGazJpShPX5q11gaavD9BynQeqYU12e0b6rtUfuDHOApT9ET5G0JkKEFy8aHiW2CXDqMI
EeOJAp+AjkplpMU4CTO6I+JSY8pl/4Zwrz3Qklr4/hm+y9spMl8iLfYDoB+xeDcpQoEWJ9WnhHHR
0Oe77olSOHFkZQ2h4zjMZUJU+ZtG6Qd1xKWoa5T972BNMwwfZTE1ICVdD11sLVFtY0ojNIJhzes4
M0O3CI6lcRd+74vhALIdhQBmd4bJ7daPe4ZWvgr7cjILaQffbRQwJ2TvsLJDupC3pLvQ+zH6l5kr
EI4kodS504/zgwGhNc6LDaZZzQ3nO99udhpPI4G/mjcfOMUHf0WYIUSEaJ491bVLQp2uKZAwBBqq
9g1aupYclnjbaxtuYfHKOx5naAl6dtzPRzOsLuBNmgIZImVL9u6REUeYZ8dxNDOFh5BfvnKxBgmP
ypV//e/GOR8bllj9GtxgKgLM3wYgFOpba5V0poD3YMWT4ndyqNoRpj31uTaBW8Pn9df4+tXNNZ5a
Glmd1urmnt7Em7u/l+y0Xm9UTqZNmpRpldBonMny1LChrIk1Vs/aCt0jlatnGRY2k8ZunM8tJsky
r0O8JVlkaA8csmQG6wF45jUxBMdvVavlWSVr0UmquwTmVNuqDc48GLvkRhXODC+7u+QyaqJFmtqF
CFWfgWeZ3e+nGizu8bKA8RLBMLCh5VAG/UqlJlWD6AX+c2/X+oaNunCqL0ii69Mo0Ahd7PDLZ45J
tGEnwy3A7V4b1TEIrUpk5Ck+AErAE+REO8fb5o6nXsU+gK2DJAHx3qxGjzbjvbObQx9mOUKHpr8x
JMPII3xbuGAjLsPrfI3lIZv6RjgOD2u29+WPqv1F4uS4edNoB2zdOQtlxDmYWPkDVT0dshvCY58Z
y6pVYfOm3fNEcW+tPSDwe0ZZ2TP5GOQjEQcJ2ZgMwab0uJnhxqsjgC1a/yJ32/T7N37vOApfULAa
EuxQBqwUoQvWGgYa1O/8Hsxzt1hIU4/zcxzodBMIXt+LfNc4HjlOYsjkwdeOxqf8Uonb969Jr3vv
bmG2DCp5vxixq8nb4qkI86CJK+kDD+foFZ7xpgL7W3+dtPdWJyoGEzv1wuWXIhf/cDZ9EAMriT3H
FF9H/BOZCk84FTqfTOKrEqurTyzCOdwC4A/dlTorgl1Nlxsn81y7/yt6KmL/UFvSBAj+ro3E+qG/
lKlWvLQFkWk9izcfAxdNXXWCAaDvPDwYFr6DAHDBefW3+oSOcHJoju2O8yIacFqTCi3C9UanS9qY
1sVB+FhmKio7VIVTw2wlGRycP7X0PzhrfujJbr8dWoc21wrvDtFLIs4DKy8vkmybPL4BnPh/6Yzl
+N3RyFCEeWkhTA7u9I0h3wUU2L0TZeEz+TzrpRUmAu3Dl8mZ6A+BeNTmFaK2g3qKjZQIHfggrP6b
MrE/vqRMYAacjL0S0bWGgT2/obAg5pEZlYVQQ9wOZXblwDLL0hwmT5bzrVaJKh8uCJ3Yo8NEMwB1
IXuJzSeXV2sH09GIeDbNYI/13LBuy53cVB9OfXSbfqERtHb0yvz62ivcuaQ/XKzCRdJi+RmC8gr+
IjrN8GodaV4NelMZdSPY+5P37Vz2MxfY4U2cyGQN5aoyfrbMuCkEZUSf3G8ejYz9Hya2bn+bB9O/
BRZkvaSwb4MNlS5PUphbrZNzdmOo4SQr0Dj3IsBXJBMxVAYaF+HodaPy5GQdFX/mvwv7RmBbhoNz
K+Zxlae92oRFqhNFM28nbwq0xqh+RPUZyjVWgAWw+ogKbn23ujNlpaN/pBnv9uNRCsFFpd8/kfJw
ZKttwwAgZmRMWQuahtOJtUq7USZhHGDjj909dl+QMiScmJsgyA876cC8TPOX60wzprl6kV++Qa9o
yqie7KP6nzG3U+zzM0XciUShhVNYyeWFfzDsBVmbB8mzrtOYoK8lCsQvgvtZF7d/H1xx9bhwi1Ga
yW3BkGWAsyM+5vp7YiOGr2ekb+ePYNfFiJUQ2NX+G+TQXZz7yAVFAqoaBE/VWd2nzHnIGeL7zPmb
bE6FoKuxrpYachqO/Q6yvMAUp4CLxvv0c8+/02dZNth+m4PTX/8h0IcS8KKCOBMKJHFRv2rMl9O2
W5TR2K4gzQEKeYB4T/w2ezj9Fw8DPiDrVMlKcODwLfOCj/aS4M2vKj7C+iDa5a54mS+HHqP/McDf
AaD0Nza3a+SqM4N64UVn4cN8bbE2Im0+B6UG4JtXbonza5zGdgUKHbdwh7jeV1BscnWPttVKcN01
asx4k+ZWMt6dMlovhYuNhvOkoVPATIkY+W6tel+9pjRFjhRWi/i6YjgTdIjmvmmnAsK4mEf+NI1G
9RqdAwebR82qgzbJiESxEzljG403TsOhFwYqTGgRE5rP4UyMOXNAhWXiI4E++sqT/QGXfEmaD93h
unXd+ccfMRRZhqy9NPYSfs1BzXBo2zqaBIYlICR0RIwu2NdW8wGsV43GGfFZRlDDUNWaJKAPjedH
8AENyqS/lj4RBt//mWwgBhyhoWcuaqYDvhLpdNVjQoVc9Y1bOTc9uF5UqGMlo/7OfpWBQ0rfdH1l
mywn26DIMkTCOghIyebGqqsy7ROa51rsK1yL0GkVV0OXU1T5pw2Om/642OfTJQFz0AxhMRP2DPAI
6giWkfqWncTAuUzm4bVn5zD1kzyXw1TIrZKPWhbUOC4TaX7u4AYhGtnCQ9fXwyYYZTAQrHIgCn+X
iJbRl/88+rjelbzy/F7GndAGY0J7Z4iix9S5zfzh9HQMOdwA9y2KxyDB8cAfz4W7fPIDpeSckiET
xp1yOJ2NUHr2Gxwmrwn/LPOkCk5luPUuZJaEDuH6eN5fSunKjkiIJQEytRMMxuX6tpNHTmzxLTzj
jms0885+AnOgrMeLQQ0ibWAe6VaG/p4yiOyt1cyWKQ/OGG43rSdcP/8wojHm3bXEl0xB9Ci5nP79
SYvL5Vi+YhroZpBjC447eev3AVvtprYhFBMrZ2oIRkqSf6pRgQ+NNJF2iVRmLjIuCAqv25yXbDQN
D/VtcxaIaI5gK7fki8pYnqJDjh1NvrKdTgEf62ixah8KnT3fQ7POGd+5OCtVW+crxilWXSgc2HvF
Zt5xX1QEKb06O8KzTOM2RY4rGAhxRYYzaI/unzIEz5/2nc57dZ5hDXhbFn1CeB49gAhDahFnPSkR
FhbwLFuH6w1uLkRR7JRfe/OoFPUwleHp7HfKNJk7YRsrMrURTic4l82f4FMq5X8PZ6Ahm45Mkduf
ID48IcY/MHdsk6RQ+VZ2VNcHdFej47JtI4EkO8ladjJxM1cX92UgEdCTzd9Bg001SelAnJIBL0RI
4jMEAqfk8V6MrCnPrStTwHf1MolXDeVrxl2SSFCXJdY8vhdY8n1pTRzX+vd1g+hIJ1yqGUc1rRZO
/+zUrDUt6IeTgDxLYMXs9QKIuCST/8rTEm+0lk2q02mqHgyth/vuTFKIgwYWHJqo1W47b9x9+xl5
YasaGL0FQyikuzcvt3+545ELplJhdwb8onSicT6X6jB6bfDz+RQIpQPYzt3lWcWiiIvMOGGaiZY4
KUxZe8EPQUlyGptFasGQV44A/o8hxy5pvWVknthcV/qm6S1pBzV/nRez2Y4IFCFITuoAAh7VofrX
JXHetgpCNmtfH6posdXQ4ekJVt7u5jgBfkOhsQP9lwdKtGWWFq1nT1O7BjaEFe4UeQd7HD7gD6cc
4x2+t4lYuOXo7U32ev0u9CF8D8Oc3cGeHuEZYipd7f8ZWyexG5nN37vvzcfLZBXuqO3cLJejG+uh
gPXx791wLkof6NiS0el/OR06B0/dWYIJSiwjHH6faULtOzTD9uD+Hcpq8HgGS0rqVtR2TIyTm+IV
heH+l/jn//tg/t+w+rp8d4mUSYiEDlRAHuUyKTUB9BTxPBB+P3TTS6c6SROwktvOxlEznYR5OsAu
9WyQEx5LKrNHbjOuEFDjJtFuVpLvZU+C8Ru98sz1CncLb9UymkO6ga+VxUYRz70yT/7YvtiK35mD
V4QTkCQmvaOKq5MH2mfBTsvylbm2cU4imDf2ENdmvHmmBG0FMihxPVbgUhwgNf5Wangr/BkCh270
yyHoHI6rv/6UwSUf3YTU/lyxEleh61mbxgw9fe3FIC+TIRJJVaQ+njtYAlmxUodYxZfxlFuCpoqR
yQYMwzfVViNFBoLu9JYnb1a4cAx9nNp+L42PF4jqJ2WoYdH5XNzoIe/4bO0MupV0jy9JyXgwc81R
zShU8NEGGFYfw+DHUcmECJ9NzrKLQfidvdjQDFBmsTtA/sAHwhau3FJw0IrnanaT2dOp8bBiD4x3
1iKR6OaEMvM+CiDoVjBX/HP+iXuRyP/cXPqqNme8NNh/TuoOKEhB+K8wXcyTfsUuw4PGBSM7LmAN
4vChZNVRk0KmndND354OoaS8w5a2KUv0c87glGNHbdH06pL39RXvDuiO8B6877EoXPlnbY2PjQWK
1l3f4GMvcQyEa24rWuxP7I0oJ1YpLmLhDhw4+mgEzDLiYX+YeSSbGHv9DLF+wE8yohvlCKzzRWe7
MGEbHGeVYgIzuiUIx8nkXej0sewd
`pragma protect end_protected
