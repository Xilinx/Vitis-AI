`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vMl/F3Jn+bbJeZ6oONZAAPbmUyI8nO8pr+MpG6WMo4k8R34R6Ht3+nsl7K6UiWLjHiebbv6o6faP
VQSztkQsK3vfiz0mgF/c23PD8JWj7ETGP0YG7/BLFgTUnU0R5WStJbAfmyrJhPmvdd04Mn9jKgBW
zCiKn5dL/r82xVP0N3o5klZK/09H83hQFuU8KdEGdErKKJ5cwaFBicXxaQ+7qVLR9xqZt7WMrEMW
iBX/ZB8YJWcFZVHDielKlp3r1agEYaQ67LllAdiQBVI25+YX7YvopU6k3gtuHSZ6C65gIjDGiurO
TD57ihw0CDtYs1WbGFVXBvOMB1YDT/8fLpxv+g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H6JCs5wBp0QM993fMUtscOIxGEygcaiMQd6LzQYXmdRksszDiTXRFjkGdbzmkkYxrO09AXJIxJmv
OHYpPb+SCGDumIiT0ikq+4EwqFo5wpo7ZKS6iZW8uYULSyV+llzOEGjDiml8a1NyNGqtpXe8jicc
5hQvCsrJWdjqyD1Z4fG6LEr7l3cCowu65JYSdTLqGrOzQO0MBd8oZ3E54fgDZ4bDuRGb9AJFuNp1
G4+VeqpQNWxsrYseXTtdNdbVmc1PDnPFt3ghvfdXTUaZXaBfGuGAp9B42u8/ZnLh0JvYpU/0U3VG
73M89IkwSVikAv128djRBwrqNg3qmkZOQBBALA==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TlpXcKQUZk8r/Frltm1DjMB/QV34UgKJSVDkIWGmf4WGGchWGcrXI3uGxgffn4k2Hlk0dxVVmKZT
gBx8b+BtVjKvtakrclKcKceHvmtCTXr6fYowtGMegkF+DjmEjKTCBoc307lnXWu2l8ngz9ezOz73
wEYpyR68qSsMZfDvwV/x9I/bL8fxwTxFuL7fGoG0doxRn3jwmYM1W97BqrXwDLYe9FXk3u2sSqMj
qseCIHy6sXtgFbMwg0vMEDN+1XVBcncCHvtJQwmgfnlxiYpE9/nZCRWFZQq/CnlWiQgrW6XXH6rl
BzMx+eCNMz9Rk93sbAO7Z82H8PvpP6dvygmXsQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7904)
`pragma protect data_block
BclYlr2aGa66uztbYnsMeY8G4pkFseuIaJ3V6qeJuwnUhh2imxpDZvmBXZ9ogBInxH5nrvLDQsaC
telcbUSA8AMB/AYifREPkfddg7YxzwJJIcK22ssiJUU7EduHy8kScUKuB0okjZfC+CzVLCLac1jf
EuVNISD9gnaTWTs+b7enHzyezkBC4ETIJDKDyaKzVEFbgLf3PszOOLsMN45lmjAN+ha6YN/742kw
Z3xVioXWLae0DayQm7/mfZKIgoa7244BZp2P+a3mkuHHCdkCqTXNhAUPk0NK4R6u/6pw3hECPrqT
eDIrzZnGgNti5LTDwXFmDVfEDeGQJUNbAiB+t3tnt/I6BHjk9PCRAok10MxwkwRfpKDtltcDvMoK
ugEBbk12TCBvGd4UD4Mld2UGLONYc8WgVzAZ0L923NLD8zQEc+Yl6i2UyJHMRUR5GrHqg8y/Qe6p
A1VZQ7HpJDe6LW9P+mDDKo/+gzNIMOkDjGEqTuNlNRiSutYz7BrJftd7Mt5gCTcY1yIdWmkENi9t
7CThWrZWLic9uPoa/AWlom2tZr44S61YT0VbVcKXGjSd7yOytgad6g1ksg1zIED+kIiLgkbRmKYh
6e3FLMYj8ETFQJ9k9OVCDGNZ2mOI4s8P6S2au/70au9FYlXbOjUOQqZ3yH5E53Kb8yWqxsZKWdzB
7dTaQybFTQomtrlAsGLBwjx3ZN+zmJsfLNQE2yB+4iHJZQxznxIZjIrGo6lKU5mA3LexxbnG3uGi
Ya6jY1KEDkk3++WRMggsvxbB58en6pWqDNwpY58N5LC/o9vB0lGXBRamrwTYpL5az6PCcjuhzjOs
Juidbz+lucyzGF+xZZtXp7lHhHzZImRTij4v3BKwlChW5fUv4OwuHcJkTF6SUEOlNtaxQm+Lvkft
eTRPCNeiO34PwRFHteNKiLdsTGfFrxAXMgD4xhFLf7ucrU3b12AiCqSM0jJlpND2c8rFysmyxX+m
IfPeJ+8kEyhYywleuCY3vYT/2lZen945Y1A8VJHJW8rLfj1H2vX1+ee6esgI2RwWwxUOxCovBCug
GdfLGxhBr0mDGlQRmokR6iB/AunD0arZW3Koq0qg1Wf5LcN9CikJqPLXnBJZ9L+jlNKYefPTPfHy
1qU2ffZRBRn6GLfLrvujw60lcIcxKCpoRr22epGt/K1P/l4iQph1QLeH60L5L2ZaNOknNh0x73Zb
yl0jIKlvmQBR614jdqS4IgQryaSyXc/r8Xs9gMiYxwmruJDH4NtSu1wjjXjUK3dtQLsT7cw768pT
+qlFjBlAIAzkXDbObMgVC1yBrPdhoHpPRGRufotc+gURq7yU2GVlk++1gxXRPcGpIGk0zYx7kNau
k9/Ubvml6WvtLMwDwqYB3cdHhH54mJELq8TXV+LZR+W3o0gZ8bnhE7oSS0OiNae1KrQwhmfJKgUk
GbuggjPzazmAIwVO3BfgvCCtftOgt4qNKi2caCZxZm4/i31lgphexKyHrY3v4ZrTk9AcWi40KJgC
JSxZTf/BWXF8bugl7PCWcH9fZ4F9syzuDJZz9PmWQcwVxX6E5lH00PDL3shJz17zEA+YZ3xodUwr
eHPY49tHaPHd+z5CavFFEloZjGTkhscXMoiZpWeq8a6BZxApD4Z6uTK7i1t5AZZBYL/CkLMWRYzj
pprJqYkCtN+xxx5Ry2WGDn+Cas71zfNI2hYi96a5oBC8QysjhyPC26wu/s3IM9abKWoyE81dQ7ky
5/4G32tfXBjqvly1jfjcd6EyYINm9dTMchtzmEIqDLB4jFEQODrA1mzcLwTrzUaSEbC7H3J2z/6f
WUFbTyZCV5LtrcKg8m4iWpAB3H/E26A+8bUfpQJ4b3ZxqhS7npk54xzrlxFIrqdmh7w250NjVsA5
caxwg3ulEbOCqOsYauIcvzuLQ2CyoSlyfqWm6Y1tGtZwGtlqZVdrXgtytnwBgvm/jQiVSj72hAdV
Zp4CauEUHwTB7VQFZ66x5GcOxNNO/B6cYjdl0PmksSLgMISlam+PwrDUKMt2bgfi+bpwNbjr9Oed
ojxKBJ24f+gtNJoQh8IOz7o1FLdtlk7/NW+vFX5bFsKsWGoOgSr/BlRvh2fBBDic5ET7NBn2+jDO
9HJzkFRHJpCQiI2ophQ2gj/uh0mYH45p+wdU/gDvU3qF5fMQzgBsony2E6SMLhQSWB0p0VK2o75Y
yOenVKdilRmta/Hr9V1nHbvGvNlVnWQ9lHZP13YLEUxztqIAk6XrInT04qVW0fwylvysD2ISQSVe
LmmofrQjYYLXj0UO7LATLHDJSnhxT+WRLOEFxKPmudoXqaQXyW7gcr3wHpzAFge9jBMnZNlbBtj2
e+XjDpXPx2n8ri3RW2Yb+jTDDYGMR2ugk1Y39ia5X8XlniTJHJqNKbIAPF6uALtxrm22RCDFDWs7
B2TizT1EMu/fX4NaB8Y5R/uParTCtXVpGHtv0MJBcKwkF3c4Di6Tfc0S4I9EipOprSQYmupe9cmU
hzW7+52fMmFVkCDMq0IbX+vuXknK0ZqUQIL9fUtZCPCZocCGmNHQDhwtB83fEVacspk+Fxw45sXV
TLj0zy/qilDTWw/Wuz1j/y9G7N2P1CK65ewrjaqcATyFnpHL7jIxlRRUDtrpOxNcK3Ew75RBeO/8
ONYGcHokC51m8uULXXT9CQhlwatMb7ok2eBs4JqfmoVl829dIgfdDxgnXf1WNW02cxPNP7S1fx6S
5zNSv1X2nsYfbE7j4JIQklwGQgVHSGgnhwtMUrfn4Qv68DYuVpf0Hsg1QGFsBqAqsRZ8HEu+Nty4
36dKHcnQqtpW6A8ZQLDL9a8/gnRkBkeDJ6/SshS9S7fOwG34WUZVNrG4OwOMXqiNIx6v4wLjtQhA
qjdFekecxFlCDwuCfivEe4KjdF94h9BBsMLZWp1rRxuG9HEaG3J+d+KwY9ttgkIOXsstkj5oAE+W
cXx0iyjkIy9e+m/8NpodD6O9WTGrXx+aaBxg9xejCayfGhdXXdnrD76vQc9R8V20KzJ2yWDOIaf0
NM4CI+Ey7sPkfGpWCULHyJN17z9Ajlqjbty1Vru9bm4TTWJzk/ZX3GzcSry7MLZfdyslxe6zME3K
s+PXTLnydhfZy71GXpr2COI+PhSspGIOfUh56Ra2V69DQkpAjet6Jrqj6ZwVM1eEshDRrq7C9Td+
KPkrUTG2HzD3iqblhBQROHNXTcMsyXm/MAthBQOWeNLv6kCXy2rSMww4GnXNwriHSJ0IiS5KxARD
/LN+Td/VqODO7cdkgU6EaH1Lycivh4l2KF0NjwdeVIJA6ADFmZ8Z/K/Ac5H2IIMH5mh7jWwiUeQs
B4jxqctku/sgUj2/OLFKhXrO2IZV/YByDIRjRCvYXby3FRNIMqfc0EdcgkhAJRs/tOfg8lYJqSxZ
ojj4PVlVkqVycyKQ0sR0RCuey6kNF5kj+JsQvUvM5DBe1fcsdbveF3P2xFUZe4lA4WkwU/2YAQHs
JTg23ONs78Yn3TMaJBTgZvCGDtHYH2Xe4W5dj/Ut1yMOHxYXZ21EmWvFOkCzNJ3hGEwtYu7WVlp4
mzcexORGb19wnhq4ZWUL6LHzeotNp90TSCJWqlxTH1k6Xhs+UYL1O4UvNF9S5ib60GL5xieg05i2
yjHmgarHdU+0/V9vm/3YmdWD2wl1pO8Dwhi9dStBvYxldBNbonrQxqAbNKbdr0EVyZb5vF1qhEmY
OxaY5JBPkwJ96WgEtYx4LITqtBuKk09vpxSjgJELcXNlAl57vNltpZJyJZyNkKXXTr93w25P3xSC
sX9FRVnlW243bZLxzqBU/JR0rhlfa1SpAdq81iBQAtYkUnnd08ZceVEcY7mYbOKYKSXE//HRJH2R
EEFdQath8YIy60Pv2pLWZ0B5UictLaT2WaRh1ppW9BvlVclMJJGm95zDm6Od9zVPsZ0vfb8M75wi
od6T0qHuY2PjXkyYRkjeqghHq3tt5UctbsF8g5hcBmZo0NAtWo+R1q/hZnpRtLeN0rH90qq+ctv2
gdevFjZrdSQ2VIk+84Li4b/aJc0gzDSpN1jAcMsBMvKiKSGB06CpEjYPe8SpK8iumMiGcXWMSl/i
U+zLZ3QcBDJL5ZRGJthUefFH5SI/AZtCl4xs0uHSuP6F+fFKpnQTVeP8hzzrZBFYSggNgbi/HJBm
qr1CdVIFMMLKj8Nn2OYfZkD5hxa7BTlMhgrkM1/JlavjaMNlvX3y0leIJFmT24XwNR+gsYWT5orQ
S6jS/Txn+7PBx0OEFhAfFjv05e3ijD7XUEDNw66v9LGNqaUUFgy9bjQZ9V08oFLf/E4SjJw9BoiK
VVSAEmWDv6+hQbrJc1+thQLoBf6JQWNe1OdNpG+7LwYMx0EEmhAoGrScZLQzq+pW/zD49PQ5I1gZ
+r4UAD4gzVtIevRCFk+yDfC7Or3lQG5MHy3/R8t7GrpCsos8FzMKm6ct6Znh1NET2GhSnJ93WovU
ELfSZXhKGOXON3/ndV5Y7Kmo+1rv3oyBkoajf+exlc72O5srqC8kloLJt1hgGSuIUtjGJt2WmUqg
K7toarpQcfuLS0fn6jURUoNyUieguuTw4E25rL97wROQdK4Mcd/YQA1/TpXYzWUVrmHRn0cY/bBq
donvv+QN07soUmmaRrlmneSBb+YIGnS7DXQM6sh7xteKZr+wtZgDqLXu8ozlw/kntmnmD9hUrFA6
xGVkH0gbMDb9PtrrewT9pqs7vq4kbwu2PIGDG3/eRZJYOib5Z2n2khVoQm22WZzWDNFu/XyF2Z39
ZY7ElVb/T3mAtXIYJxdOLnEfmozLPFMMSJKJrCuVDjedVQcCvxQr3aZc0vT5YOsIjl1+jm3t122r
uOpHT2szRaH2MPq4r3adV8+bQD9mD4Cw4U4Qfh1CfSFqWQmscDqYgEnIVVBWe5x59lHQF3bplBCw
9UDl6YhsObzAo5PRkcIvrupJMWSSkKlJF+yN4VwY01kK2bd/6PbnGZ1xgzsHJS2ldMgkQ2JqAQom
NLn2aD789fsznqEtGi0i8upm9XFtWje9pN5DvAHeDk+f8TdkN+QGlLtAl7Vwrg5vYgow8z9iiI59
66vYngGcQ7ZIZw7thZQFNU38rzDK6meoG7+bDv3M/lsWJltIGIn5qBDajBf8HCMVXF2bEqDzcPlK
uyQXwQWQcUt8A5jZFFu/TTkP03WnX7vb/Nlm9drkExw/4mLpjkncQEonsEv+Y2sPYArYyz9VCmi+
7YW1VWKRBhFUzDYJkeb5fpHEwAN9wt+wxCCbl6wQeeu3jEq3InvWhS3BarRyrGr36Lt3jyVvdigO
OKyVHLaiebSsIMSrxCkec6tTnQR/hKI9sMMLmFzCcvRtins8Lb41tqaVoKFTRYNx7kGFIqTDDweH
/0gGqV3MIbFYYgetV71sghtv4DTROnKpY42TWOECbGHq6VvrYbPlJFyWswS40ZRC9p57RFC3QrLo
fE1z5KLyQ/y0FB1t8AYwtXPhpzWp3cx9By8nFO06KWRYX0Whorgg4mSD+OySmB/oaYLNoimwsTc6
e3dnlK86oI+ijd2A3iOs3/XhBekjvC+qyhGbC5mS+ZkUAV3VlSfMotFdS/LnyprlFeqnvyyzz4QM
DmkVFBIuSSo6zZ3YClhL/Df59iL94SClc975DdbyHOYtn49h0TfOXntJOzVcwEC4t6it+4Q1MsO1
HXtS4m2VYss8Y/Cp0Qs0fid3jkxRWjdIsincLkdW68CRyC7n8JTXud3lX3I2xTgJ0R5xFd3fryeO
rpTE3q14hOBqmJKY6lGTlzVRrl9nRnSB3/JweScE6FeVMHrib5QYWr0TJdEVfz1RquGxI1V5fpPC
3DPOUf7D3B8ihufosl/bV1E9wJlvvWCKSw+bigLYhvrdEOTVjC25e1lmm/0YcIs38RUZp+6V2RBW
tVaoj9oiNbwkZkvfu0TjIRQSdHVH38RNmBp+dXeDRaFHpxj80SC/sMeItJoKLNORJp4ftc5h7FnJ
dh2ff0xVDUVDxa1CouD0AZhg8hpj4jScIt6GzgtGzwAL31JqkATNGVJA+OPYP36bsvF1djK6iHbK
v3nYMMOHho9jT9V5pXh4sK3jAjLHOXGX40c1tq5D+uoBfqekfTzyNAzFXr4t4en9g4xNfz6ZdAhR
9U7kQYJWtSy+aKmERTO1zVMuv56nBNwVOtXGzwWktTkBCZV1e8jo6x2PVKgR+2/F/Rm8i4Bom/V4
30YSLxPwFJbe+35sR6A8lmhV0p3nZ09SxStKhJd4t7NqH1rIXHTcsL2EFibsq2CkHm/K8n3Y32gF
FhRiiwvg12YhDysA40XcU7mT1FFh9DFMVYIL62dLmgVt83n/qYOjAbkpBemw2oHLVeHEpUgkaBDS
DMx8safkGbDvfVg9HYkkPtIbq3EzLhVR4UNXv/K/0jiYwsg4t6w3vCUJ3Sa7KpfHmJDMwV/+P6sr
DI1bPI5rw+/CAgTin6tOtZXulxFg8vNxmWMi1TD+E2VzUQ89sAgY5tBhILzu/V2D87ihalYPNlVF
GNXT8ydDwI7XibgxUhNnkRghURiLM/aBjoWj4YEjZJWLhHs2p1bpNulvPtwzjXRVFZE5NygfFAaD
ZrHLqmoGiOo16JKnb8/FS5/UhGVOHiS4Ev0o5W9zoqBtwkv8CWVZl+IjJEU4GuuV36H/svOLYKkP
L8BwYDGYIA5B4FCPDOrkZF6qHrJHbLzmjm1/CspOpXPwCJ5T3nWjnhHMYJP/XhAbFPM75bkB7OXi
NMKEDKldmr1D29LclwEqjVwTjwLurRigIVDr8p6j+zvdzs56EgCC/KpT+cpg7pKHllRYJ7FpoMuO
GxQloKG/APwOWbHUiUbAMQu+2Hu7d4VFidcB3mxz72yMvP4xclQfEq1G/oxegBXmTX6IEvHBpQzI
+jNaIySoL9/IMDDULsvocCadK0T+0PYNZlvjIi4b5TRlXKIO81LgmM1YLiSgAUWeG4LxMEPqGhD7
U7iCme+QKJ4INgwDHV4jdTJmIcibAwjngyrBmHj4LSXNCxTGPe+JotqKmWrnCqoLTMTi2V5rr3ML
zbnMdKIHE0jOaHLn0xpITOjrvv9+xjo3NBsaFs0iAhXYx0+VvLAB7tlomF8E/BbmygBJbJE6tPMs
FxBSOWIenVHQPtReMqGI9iECIQQ+aV2GDdSZC7AdbKbNxArKN6mW3O34/mcYouIDZAS9rJipvNn2
JFc3y6U8M52Z6B7qumE46Ma0Hh1vRJpOtUQAtUmjpFGVr/D9fzPOVDf+74I0apxujXHXGZm70oV0
8PWEYKrzXdJWHj3kOsxg/wZY/HIx7M9ZhHOr+fI8bNYISkUuGg4bwLml2DvlJwkHBVygPYiKGS5W
ndSGndbDJV6O+BxBjP0H83lszmQY7KM/vA0Zy8hDd1PYdXzhIS/LO0O5abp1KUYhLo0eqfNxulg2
BVlXUQk0fuKxw6b+iJ629hg8YZaNqTXgOLAsXSS0vhxofYlXkPZKJovchZcYP2OavHyif+3r22g9
0hx6CCnNxUlfzRIpFtYI2m6OLTs9QaCwPcOxsYsRfB00eExvHxZgNWFvYYzMA+T4Gbcf3Y1Cxb/X
i+0Voa7aM3i1BPfES+bdd+Nh2aqE1sC5FV88ybJ55UpM21q7qq4H8T/CIdL67G8rvPd61RcQm4nl
bRUyyIbBE+nz9UnnBn6dVwsBBCEgedweO2SjzuinGaMvXDFZtMsngnhXw1QCar+dKZfLS9Q9rwnU
tHLuhO6BC038sG1v943Egfzm3TW7sUi5wYbQn9h66bjWdxGMX5u/HH6rkMGcH6S03yheTIrS5xuy
YkufKSrKOxitIEyMHfHadett8MKsNIq/k0lEc60HWw36tXNBC+07kc5DGMuKi382EfkPfRoRYfkx
bJ9cQ+VrB0FhRZABgInmhRQ2kO44mZkWRRRF3zFwMgE0egx98k0HxyHQoywozGBFXMdV2zWxdvrd
onnuaHwG1NF4DahHmTZUC2/ipgH+kPCYaEVeRKgVvdoVfbbeMkhWq8j4tUnC2MVrGUGTjUt5DTGV
vzjpIO5Um7CWCLpYLxJNcmkTPg35RGZrIu1ga/oW2ZzL654UkLP5LqiuTUccx/pJxUJx9Nh0IsB9
ETMFyrvNMqMTbLYmRSVJHZxhMRWVM0LhQRbJdgJHeiQjd8uP/FJEJ+6Mp0huOIQv34+ddYdE5G6M
QAYwZ3ZgirFzPwQ3+4ZCLTR4ZhmDNdcmm6zRAp5RxwjmNMKGx/FDO4FN9V5kAWIRUAE1mT4sRUyQ
YPoFpy/M5ytVF/eBKuSI7BBdEmcBvlt6Tfk/KaG6s97bIaH3PLyOYWYVlNPvAY2qPOGazxkDpw5Z
UrMM1PV238ZhY7C3KpPe6144wc9imMKTE5L2eZbz27DBv6nxO0eJ8NdWpkCln+uSoMSim8b89eC+
t/WS3TWIhUtDLFUHXpvKu9U60URzDVVSg7aOJiaGOEKluEnNUPJOlR/IOXqfKFsyuzaiunynY7OA
2Mth7HDtasFilxErHOQuXcoHwVNduSfECZljN92GorG+FjcaBOPpD8G+lIsyoWJWjRW2myyceEK2
uPYjOI8EA7PX10CcNryOornsP84E9rBYxx329jOl8xSckjTSCd4AdSZrS93egVhUmN9GTqrDmmq3
vdLryv1JnJqjMdwHTCic0owZgIJeMXKY2xFgJ69oHFjzcj4AAlDY0jceCaD2f/DSX2gEupPBAMD8
TPOHUtXoZEbZcJPJWDjyaWY8HSyyqTcgCmKB5rEPp256uSKE1YA+JcmXHO9r6EQc7l9VF11CgN2b
QqlAG08qYl/uoIFOOJgXPFLIj65VboU2aX/HSTtppscJWmOGpWJS4Nqt50SBq/f/yNG2M5fmQWp2
u7SbscGnt2RS4lDqcoTuOiKMscp4Ode4rQFYia/hL16bG9rwWf7e8ymgyTZOFrz+4+Owfqqo0Mdb
/5urOZHL4a2F976tJ51+aVF4Q3OTWdhL9EwmUIP/Xz/DXz92yRduxKFxG1jDl5ai7ElnXxwvv8e4
nP1m8Ks9W2gOdi7Dj96vi5HxHwa1r4WV4uub4F15k4lhIoKkcq+Rx7++jtbCtNVBGQdzX5iLpHnR
ZbbaNJfY5crihv5AKXYdjVhIZb8vLJMZiRiysymFaYfMSJOHQugfLBCheV8LOxftFcmchOLfWHtY
yEi+ni6h9A2pS9zgS1AAuxqvXRNVgMZlWZXsL5jSNDNQZA1snVRwhWZRCy5o9w0FWlAskU7W6y7F
IueTX//o4ysP9s+xVVT4JLNi6ZJ6xiU4beaVm3FOTWQYXkAlEBXF/NtlgvPMtPgi8pQ5nqP6CZKC
XOrfs1CgI/6EnvD0zHyJ4EdcYddYJlk1arRXlrSXv/AT4LiiJVxqCRLGFT4UzVurIL/yPAhazOGj
U6g9vpR3j78dgvSZmLH6oFqxmw/MdJjArk/xfNOVQL2sAWcdScBae6iaEsW/6o4LcXZNg2uDSO6/
Yph75HruVwd3vjByhi2llozcsYPQkEUwUa7Ay7ivd44ZyDZOaRzfkeC5RFBk8pmLGSM+LvRuDEIr
oAELNgMEXYm19LRSQNip5PDQSdc4ktxfkDEGNewARG1pZdS1MiitwgiCSb6PhgcRYBtEpTmiARZy
JMfzRTKRLd9srpRWXf9uJrTIWow4w6Q031tmqbkIDD+v7WbpBpWOqiqZP0wGbiNJS4uWjRvBm31+
jm5Pt+z7q3w1Vfzz1zaLVTNz6HRsZA+WJ0PaTVMLProDq75a4M+2Wh+RuZKPHRVuQSsVDFn7KjRC
yR1u+fZOFND+llwRDWfDMyaOF4SjV7bM+QwsDMCepKLiEh+9UvleVEDstJDHljLjREGihBXg6znE
e7hJvgx6ZBa6BbJaIBQpLMHY73LAhxJdJt7b+xB74ooHX8b+pTKs570up5EaVA4M9LlMTu9mAKl1
x2LqBjErwMjdGngeGoyyA77WG+wGr+XQ3pVoP8jevvHO/XYTkxxrx1bnISK7lnN18ddBvu6Ji8WB
lFBBioaOb09u9zG44nq4CT9+A6/IFEH1Pwks7RDlyqr+Cmzbd3CbYjCp2Nqc7LKZC2MhVNoBXDU9
qgxA4U6v8BJ8RDsQQMS0iLNld/pYCBZzFaRUptTxtBPLNuhTx/rjNfysG4VojmnEzTysddrnW9bE
edyIKIRWYc/cndUaISWAUgEFir3J5S7mv/Da5Wo0yJxKOl9FWhPx89jqJVlvgK96Wb5jr0i12byM
9iaPZpn64qvjIaALeefb/m0iQrgRYL8sW4JY1oiKRXLg9Svj5TO0OFL4dN46Fa7XLWQbvSoEGcDu
Qs5IGe29aDKnHF9UMb5w7SwqCsepk/befZOd/uC7+ee7xUXl0YQH5sScHZrtap+1B9IJaZuQnmkE
ehL15wOtZjtdLHqHJiUmXutFundIrc4G7dTXmkutW7AtJZIqOqVLXldOGYsBYS5kd7CCiA66nDXc
tKq70TVrnKNxmy7xf0krDGiWfOo3uVn6DHNErmbTJy/naJtTZZ8=
`pragma protect end_protected
