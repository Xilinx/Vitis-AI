/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzKH/Aq0XzINrqqhBdmPC8vXubRrBqn2uaJnhxNxRWaNkeSbqJH6ByzT0
fb56tDseE8g9RewR/6p6rGRVYpfzQeBbOjDY+deyYGds5RS7A2Np8XTNeX0mQo81+02T5tUbMi/A
wTQ9N2s4tLfb/ym2azfRjGQTWlW31JZUiJR6kSKJUOh+bOyub4KKsOfd1TWlrANLixPwigtMDxDz
QyJJQ6kLSf7Fon6D3gUcE2JWqw+CpebmxW5njKyPhF909lgop4Yrol9zT+Q1am7/1d7Nl9590Zwi
OK36TuyRnZiYpOyCQ5VekiMll019ynmDZpIyj5xGUEsk7wnQodUutMsWvcgTboQRGTQSwA/ekTfr
l8WEBqsefhspqKq9aZUiQ6CEvEwbwD5JtDAq7/EOsGOy2HZ6rB1ec4mbsj8Mxe9G+O6lOODiNndA
FaAYU0aDAu99mZUPRtB10x9Or+7Ut5zrSq1P23lzH+6g3JBrfcLHM4klRYyR7DN+4393qLwyEN/a
9uizHQOOEfNJk2z5H2Qr6bI2AC9Lg2z++Z1llszqXLD+Aad0YnP6LcP+raJ0kZpa2fyx4gOV7KQZ
I6ZMc5XmEbl2y2/eZyk/10fciZgI2aXTZD4PgOtcTu7r19zsodo4KoE/GMdH4maV4NaLTn2w/OV9
CzV5qhkjAhrGc5kvDy+xtf9yXcjtpB6SbtjVTP9MpBOKQcVsNiqbbQsQN4LMERSXHT70GLCPVCMp
R9fQraWoTaax3LMZklEdDnHjGjrRihrNxOiZqReEIr7aViW/ZSbCHmu2BCH08M0sXu/orzQw5FYU
IzAyRNLkqYDfQnZV0thDCXB2iKIZ93d1ANbj9AOE6i4iYhaI3KkYMSWDY8WXe4YJY6+xbmcD2mZq
pUi7oF4NuWUk9G5N81LqWIZOnw0fJdOQ2V0N9wUO+RMrgoHNpr/O8plFC8J6HTkM7PE2bQ3lXlOg
szKfJKUw9ouZbmqvoAj4VR4jHHewBbrI5OpTmN2rEpv6lDJiMJ/9AWDDSKZZIBUiZ64yWMJQDaax
ApOEgn301ZT58VvbAbwVHdXBO/D93GLBKpIfWzE0z56Y5B4i+Mg7a4FLvo85hi5kOd8iHjoVd7TD
D9ybFOwCzvshciPkXyFgc293taKaB3gN/gtH7A1Etgjg3gW47R8uj7EkHQGNdfd04p28dpj6oHkF
afhSLHP36HAzSMGeFORXNV6m122vkA1OC11P4tuw2IxgnnfXXto0lozDqpKTyU0pUZGk7aAhS3aH
Bs9/BA1vkMzDaVxDurjW3tUsar/e31Genz53Zmn5uDhQc7dsDs8b1rDKEg+ub7Az448fYTTSTHx9
CnmK/MzT+WyfFuTx8q47VKjcbGh2f161h6Iji0FA7zWKy1M2zhmXGzAVXABKX1KxyatLaT32bafg
7QILv68=
`pragma protect end_protected

// 
