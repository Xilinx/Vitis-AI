`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQGDi5+1T0zt/Jw20/MosUf/BG/H
bU1FHIdsAm6uft+7I5naFNkYDFv6fsxdnfu/MX95XWwn1vRNirzvgSpKb5hcd4QOYknPGL4xojGp
sZ/5G0qZehfOcSBTUwqBYwtM4gmLkZgrLiUWeW/+FNXWDn0NY2ltMbohM50vnoaoynLxGMkjWGST
+ShwzZPpZgxAGOV07TAjXi7/AwOrnFMZ42eEcNsk4cV/EWOJETvBK4Qlx5qPY9o0o6lB5GCXTCjc
GpWTJTA1zQAu4sDSWr6u52eLBALArnyjCSlPosz2D79tMDfaqR83+CpBFKi2HUu+S1bNR7Rnv/zg
2vloEWatUJnPzioDJ2oMpVumORMa9g8ZJgmWDe4Leob5fIvUawsR+pOt3Hj/QpbSO8GaAAuRaI5h
9yhJ/1HwXeyGAbTcxcC4EU/K8n6RyvlcFfc3ENjd2WWa2E1yr8ZDcv8BsTaecfUVqyZy+naxN/8h
uzyzdp39pOaNprLeB4bsq0h8QiuCX16jVEV4CoC585sRaCvBjTnbdjWQUxHGSDnyizvf3xurVk8U
XfPVxYaPxA9sVGnUPbSEGr4bkKYOWb1zwLw8ayEZcBrFmAG/r5q9oZPA9YhJoAIoDidmU9iJ9dzP
xDXd5tMrCp6CzyRsn+k4Y7SRMQPmd+qGDJJKF/w8qMoTUyoEwphnQop1HtB8e9Iqwt/dTXi3iGrq
xQaHj7QJXnq8U4ba1zGkFegfkItJtp6TfSZnRl0wMudEI9pTnc9CUVh1N2tWkZETqta1Cb4LMyPw
OhAF7rcF8NAOJlafDkUKsFJ31NE2pskrHiBYfYX70w6dNeDrTligkfrzlCLkF4RXbxeWdde/WC3w
bhscyD+HQoJ9Zqz39LdDSVVVmTdm8B5rkmrNDCdx2HFBsg/fW0XP7G1BoK6uhE1hwPtVmfWTmAzS
FpIr3n7YyaWizLDFO/tIrwg6b7PD+x+mbCAd6+1PYXt7TAP8+OSb1nZvz90t2Zbt9tLvyYFNUaVc
lwKmYflZ5OwN9R8n33FNZM8y+a9ELZLwOcbrScvN6lqbv0y99/H3SmMx+E5NNzIXUJescQs/Ccyv
xhsQmJnE2Tmf998H5EXkb/Ji2lUeGcpUMv0NQwXTWAA+SKwp3JD2RwNsp8i9Uw8twsEMW2k1R4jn
o3svSRBcFWJxaMNpHEQqX3OSBZt3wpqNnh0VUbYwixeEvYiN6dPXoOLYnlcZsakG+FvwjLLMjuvF
6DKTdt07claGhNzaRy+rTbicbYJZQD2UhgXe7z004Ix7VTKyIObSaaUcG6fvnH5gOwm9bbFmM/yQ
hRkvvR9isZPXSo370iv3LgdPbfgh/wg5+lzApFAegQH+jz3kHoZMCYlsQK9PV3oz1FZa0iOMgT6+
SjSyfI4XXAU8ya6/QXiQ0yAZHJm+kfW3FIHle7gbYwfqdFsaVIctRrJjkvhZvLbwIDfbcu0uOzNd
VIidjcm/Zlcxbd/cnlzAZX3GjJYT9zI0Deeamkg7hcb+h9GN05B2AKxAuJCRV01sxZyvahxf/zEo
MRdnIR82/u50isq1+pIJ14oxbxo0yu34k/Q3uQTuWERE7ALvry6W4tmOHXxIKN0fNuJYobTrsN9/
si8n0WABsg6DX0f/6udMTV9WnmA11h0qEuu7CK3b416OCZIT+i893fe8/7iOIsSUcTpTqMb3RE/N
jAJetk1I87wUvB6U7MbuQ/koxdsq282e06/Y44FiOq9solL8+CFJebaANWPeSDIfdmTI0tQWTtgY
/mNV9dLzbhJG7QQAQnx70lyjqREUNUnNrygXy2ChJlRoRx8XLcVjs1jzPou1wL3ghpFjywvrp8ec
cszCotg5bgPRyyEs2txLgMU02OUExsSOGD7YFiC2L1dQ7hda69sZe03vvGl7vHtGzLtrtzM4GnOo
kYDQ1AlyMXqlOH12+bLECBpJV5cLuYZ4WaOhuj1aKGCxkrhQkQcrBHM8JQmYknMU4N+JjW9cDBTA
HwnIoJtRox+sl6l+mwVf6KHiKY1MIh/ZADo6vY4JuR56dlixFrk1gD6Lr5d8yJtATh3WrlqXFnmg
ahoIFPdTsX/HYxUx9rbR9lzGmKEcEYYR9NDsum889fWzm+h5fC7qQLb+TLmxsDMFdMfG7RndsvZ/
IvPFVfLOnHKgHj4C3lARAw6WPxEPka72owk2QyO9w5jxnI24PnbTza4VKaIScwoUSoIuRc770yx9
s9s5xeRVOTiYbrPAGAAyYvLM09EBrbVDXuVd6vYy+ixDH1eVAqiQgKXuofaEZCK+FQTUWLMXu7kx
VcQ8HeiW9mV7XPJ830j1csxyXAQ1NqESR7fzmlMmxgCcf3K2M2J11mYIfy5Y+RH1AchF1COHVtSD
MrTymcTjqPK/n+wLBy7dnctMmvU/Dgv2tYuzXNE1f6OSw23RsYsV/xx3Yo/xdS8hp0sZTEcyIRu7
f/1ktj3lEcJfbuoZspfQG34Gn5QuCRLe0W1V1hZD/0JKBUfzpnnsapNTbDV+w46JbM1QxftBdyR0
8xwcmnY00JQUQ9VkyKRy8+r7YrFZynBbHmMIxWJm7XbCY0jGcnx0ltVBspIcZUoZEryVxCth8zEK
GdTw1d8TkEgVD/DC5FAdqntRHhsNSz1Gl85wTrhNH9rJsUj7bBrVXOiwpue1RFwfN7C2EoWSgX37
SdEF7jdiSmoCT/7rzVGeNYDoNfnp5BOLGwgI/YXQRv2IWUvQjoH8X2Gq513WSTRdJgIbCE7924OK
Ci8lQpB1zvqhmhqqdVYtw+89xQwe1Du+LqzyGfvjSqovs8wYESgGecT7p8yklOJlCTT+BMXMuTNA
y16mavrrWVJAmCn9v3c2kp7vl7NihG0PkT9vYRTYmixJlIDf4rw4iZnoYx4OK7vLjv3ZLx+bOFsj
nq/WtmYjBF6b3O1E/uIbP5PPI5IV9bP75OsOKKxk2fFfX4vVW7/Az+c1v1irSsiW7L6gUMXoThsS
YAYA8Tlu8Xxo/CjthvsDIy4zQeTiWqLDZpn2JwcINhDgb0r2uprJ0MXYiakU4eFgDzk8lMWLsjmI
9vsDDz80sLHyRLloEHeonnu9Jwzs2tvHBP3RXbJVDjl4tTqzQDbGHJl5+0F80JKc+lzqftdjccte
ykv5tOk2yQj+LpphTNPZ3KlllBn6FdQBHRo4XV3/ht883mi3yUsBuc7wzl56rlzsWWFz/sUdHLf1
xi058gh1zHP5h4k3j3E43EzyS7yO9ejTrLvdMIh/9e0OwpyHRdAG/7V7RoRg6REht9xFgoij9fEU
cG/tMtlnxnSIkEEWpeJVYJV2B149d9lSf1njV03MrfVtJXHQJkGNZ9wbjMLWMYXsIJbrZWXcHhF+
XyHSdG9JXyF1sr2z9R9QdYMu6yFSNJrMmieU4lAj7dQN4qTCYA8qZmpux9+xDu+K9YHA1qLJn+or
oKE/vCr96qiISjcC9GbhVD9+EsoU4rJASJvzWsietrwe9DsBkGcJ4/Xd1nxDmA67/0MOT4uBeGhj
n4KLo3lPscNifHYeNJhVBC4ibNL72qMHwPHse9ziubEMYEez9p7I0qBE2Nks9iv9dXJnYkMbsdJY
1DlVgKm/b14eMGdKaJe8o7jl3VyLw1p2d+WZoRUWX5UMH9a77axmv1Xl7a5fixsp5YT/nV1HRFTY
d/SlDg6dHwX7t3FMB/KpqyC/kZvjXwvx4txn9iDx3f29QEmWBVvTqOSLazU3rN4OcEWttVkWILwz
Thp1dqedwF8U/uq4XNFQetlg5wv1mzQepslaiVxiTDKR4DSvst4QuyH7DqerngNINeQArX7R0iLT
BwroRw9AAYj+mtJvOD71yrYzkOPXU9ivctG+JHvmHTDDQwYPTpV6zlV+yC+zCDwuf0XjOfRsmwFT
ydIPvaIh/pze90hR4fxEJyGja2QOdYTos2rQyOuNy3TyDvcK7qhhD3QhTT4qsw183FiwJIkb5Xzm
MIWzcUT0ku0+6VOYaAj8/aOpkEoZjtwJQKNAwtMZ2Gu1cBAU87tg+HfHbq60Wa55W9uE1DU5TEsh
oQITa4MK/lc7ZWkmRe6jFbA8v8M4GRdJsmKDx8ar5zEFp0pA/U/zms0BRS43drSW2+43onv2XsqH
a3gklxtuIZn16wwQOun/qJ+No0b1fX/9k7jg6oNmDKkSfmG5ovI1OTTWqdzCHuTP8DW7ttbA3pJW
Hl+EDymg/A91iXUarkzcuhXmT88XTMu38T/eVvkoHtfjE1GxH06ME9XvpBNLMCNvR7QLvCdexsQt
e46UjvzqfFSyI4+T8eOCCQu8Z3x6KAvtGX2f4bk32TZsoRdymCw8umAVye7srE7BZ29jGDHcW0xx
gUtI3F20wFKy1nyTuamnMmSoE878uhmiVlIaGVMLpJOpDF8nnMWUwzlTcagpD52mEFMaVkWoUNb8
loIm0AcEQVp2iQEySJESv4YCIsHstCZ77amIKhMuALsUOpUlyHDvxdW6IEMarvvOSERLL6v4urVM
fbxGD/G7hE55YXzVQgQOVx9T/O1ncG9LibhQoFPIbuztkpfsl+lRiT0Od5y/l/lfZlltuf0owZsj
g6gvO2QbjRpd/FFgRFLpG8FJZXlp7qMcYH1FWcIrVeORlfMYOmgfKUg+cf0nsU4GRed0Ap37LFh2
13TCraRdKhr9+P7BJsWPfKo4m1HHg4x6b6KpeIz4OQk6jCNA04aV2b/nt3yT/ke+BF2/0/OpkMEQ
9YO7gdJp9QwKkrk09rNKA2gOM2EB5ZSQhEYsPYs1v8Y35732ehnPxln9aJnxvRDgc8CgRnd6Qlj2
FesikR9QquVp8+AV6QRokSUcwXOMCemszLN80CfMeJimBypDTuhKjRodZFJnEjxnEf0dShPmckRC
kZ0UNUAdkzhSipFISFjjIIbdtujv0nJAqHeMH904Ms1URlNnk0fud3qNC3LZGDdGgG8MPag7ga+B
VyyDgaPNt0ScejHfo6Q2j/fdwNr+NkURBA/ZJvzqEIyk1nSvL1eUCa9dr+6I9uiD2pQ/eMCAPPuW
7GDfiWffxOnl153NtRt/OUi4T5L+eOreLM5s8WFBoFgpHW6T0DWN3FPUd2w/kGE7BuK7oFskgDny
g8DlQO+Ikux+HPjoPmMixQ1P5K7ggIXRlwgMubY/pYaclNuGYh4g9cisch6isxBHkqRZKUN5MCxv
gh8l2WsDnQ3VXZVWsXv1cVKRRBltWzI4BV1JccMjOFrzNzajwFxHYIHj2fgjfSZaQdbG1bf6ycvc
gdknlINySHAcM+k+wxvWBuP/JVR0q6KCMPj9RuY0rCfDyMNYlTT3Qh+UDeLpOZERUEO28TAPZwSJ
i6gEQZOpyJxB7AMCm/gjjg7HyIcl8vspjC3sPIqK2zbCB6CZxBUDv8B46ZOf7kQ7S1bLZm9IQXG2
SZ94tna1F2BOfTqovMh6UvxEEX4Q28eDhI2lWA/+wpVmfQ7+IY8a60B5DBIh23nvjCNsXsoAm2Eo
Em1z0zcZs/Q+6DZ15FDMA7nZ+gw1jniCk7uoWxollXgF1u5utfWWCLpI0m82tDy+FgD27JBlnRXU
t9VTa5A/xRlzMs6j4OzUMMbKEn+kzncguQKUmdVSmMH85cEBkHlATXaG6I5Fx7B2fkBCVd9Bk/1y
QC4Cz/Myw4Js8r/1CDOz4v2Y5lCz7VNYYpNXhQiLW9glKfCqBVMhh8ySfJw4xH6EdRU9cGc3pOt5
1vQ92k4yL3wlX0oPlQpjO6OjBTDfZuMuv23OntauNI/KHnZn38Kja1NM8VFJzItnlfaraygg5hgY
BOWhp1I+/Dy+huO1t7RDSbcP7RR1fZn6knEZR6d1W/Ixk2ZsvhzA/Hh2+YrzZxAT8Vb3eBlq0UYu
SyNO1wLCtBd4ddada+jK0ClYm5mw7lKadrMFez4V5yDdL8GoJbh51OUQIgscLHH4UCGak5p26my5
7EQQ4yC+Wp+fBenJdSJeNL84kfdorLPg25Y7ERzhCtPWbgiCif9iJhmvSjAhgmKBvcv0lAm288PF
NktSlTQETSSEDIflNl0twr7UfNyVw8wNUnkkVRgm/TJDMF04UnT4FTc9x79SAmDUJ+i32K6cSu8f
ZaTrqYh2yxtz/Iyjf8XhXUTKPcyNhV4UTtN2kSywEh3opJbDHT8PCxSrkEuA8rsdwXtl/A+/LqyW
iiuRtm3tVrjMKha8CfvjY0/qVv3mxZBnZM+9LP5eIpu6j/Rydl9AlrRt8/tvIqaWSG0Q/8IaMXGb
eV8vhWlRDEb5odfTFreYmxTyis8T8TwsTnSMmtKd4b/Rs28jFsMgZTfFJmOsPwxuxSKjggH6C65Q
3qgo2FT6POW1MoMex3C4Pae2kL4CAoavIcMB2uhGwTnpDRzjwEcNiID7CLb/J1TpZ2Vh/FISVRIZ
y/pF0HIBYNFwUz4GRNYmi1aiieGVZ0cuEsOyYNQBKknXuEW7ue8JF7dCTI91qp/zMnU+LuecMGdH
Ez2esZGt+sny0NyDKvXqfKL6xH40/mhVvRNecVIqKvYvbjivZ9VB7NTKvoM0dLne1fZ188oayjwM
qiPVIMzqrAHhzbbeyjrLS1oyMMvFkq2K3q5c7vcD/rkjXKgIMlWOqmtSl25wMon/6zOnD6SY2zjh
J7RSV0gY3g9Y8hWcgkUq7I2ybJeQA3h00HByPDLPXMm+epl3rNuwnSa12V9sUZVMxLaXOx6+ZV6X
yTi3mzFUG6qoO73CcO5ILl9oWDEVy/s8jBSTmfZ8Td9JVzsMkXWNAF3vZi0Q7RuF4IrF+YY4SO4E
TULeStSsoke/Qnv+DtZ0rQ+30IBLi9iDfRV3/noOMEtOdTa+lOMftyL58nqXaS0PvvZqPrmduDTR
9twjPnBvqIcpUeNDisq4ZaichiYL9qgoLGh7IoD7hyK2ZQj7WiVzt/79IyxXo1odJRRQ2XsIk771
WQNNSX0eeUAs0cSAqCoZnhkbAWuPOJUSEf95lr8ts+uyiTkv4KYHTL11AgJNGj4xMPQSbUb1uREZ
yjmX2t4ZrNcHwqg8FUfQMNSDReoJq+TRHQP7AdnJ0q0JPQbWTe2Zq51v9A5uH62lAguUKbyIM+Hj
XjYw0iUHv1MXc58LLK/jKEgsTohastcJP4Vbka/Voupb8DX/I3Bh52+MGk4SgBCi1wHhBgFxl0Ni
uaTR6jo+UIIhDm+mSaufbshDkO3mNMKRg/knNNJ2RX19h0SYHoisckgah7B3uqAhynFUoIvgWOVP
PU6dzLKaKb1ibtQWXjiKMaylT/Smyt3Ch2chsq54LBXFvRXHw/2wZCnJ0y7Pz/9YqeqRx6xrwt8q
F+3ciOT1aW3SVY4TPn8FO0g+4U0awkK8HixtED4Dwc3WZswWDTg6ltMG61JKbiusTwLPaGzjdxFv
K90Tz97LhxKs5YtbAPWuR1KM8FT8JMztA5Z63xz/xIHpmPqgPQ+54oN7tthe4Rf+nMZ4HCiea9so
V/GUmIQs8d6Ta3RTEWyWa9mSTP/9klMpyJRst/DOu1pzjKZDSOZ8ulxr78Xcym+rpITlS5qPATYn
21NGgB0zBGd7MYQECmbtNon5sFb82igwTx+oim89t90G9kzLCX97Qz9OK6bVEbZCloNb+nTaK7bi
N3a0duVkb5YudknF+h9rqLgVrmz1LT8D9hqtExLjr4BQS1YtksJ1ilzI6XmmQnVc57CxasgzQnt3
pHSkyI+4fQkZiNkjWwv4pLk/am0suZxeKKpYgqBuu+KojzJ23fO29GA2KfGBOY02BzehJfTjdPwn
HnkexxnySfYjBmEDX9LuPmVjxuHwp6dIfVznJ8Htg+j1tzwJ0K8einG/O15i70E3N7qeH9DK48Ys
r+QA0vTdgBZaQGsCbFuNU7kbj8pHRN56PwjxEM1IMX5fBCy9Xqwwm1ajjW2ZDe7DJWdllqQSaBAx
64MdMjtwDIcpOaLjEa94iVzoOSUPUnicSihP1Il2mcs8R4qkcfuorBSi6Xk22YGMrHhSj9OKjqeo
sQuou3QctCnSEdhdDgv8ZF8Ltcx8WSFKSyzqp9OCVek5UTnn2mepi3MBBqi4Ma7U6mJdpYFueLQ6
rYr68TD2F+EwYiq24MafSLY3ovMJg33YeFXyQIY5Tie4x22aqQOsDihynNwWZL1FWfp3bJPkhQ6m
7gvd5B/1rv9y3fuxeX4vz+H8pv+5hfv+hW8zGz2xKaDQFgQ1MNQO/EIxNCr0/hCLSR6U7nVg9iXR
fhwMoVllF/LrUE5bKisxhEpBmfMokS7XDLxhK7jsid5SINmRkaBaV+nS9l+Yq4c5ZIV8/Pd7oUEM
1Aw+BUf0ommv+r0H3d318RDDXfwBZArDQEjVmRqFZG+WT0UgZsgaRLgCs+1TojLY7rYLV1cPOGgZ
CBgp/HbhUG8TiOzD/JL6ZaYYwZTICb554cfeb9o2sWRB6fjkdKQBnZXv0w+Kxpl86a7iTJv+uF0r
YRTZG0JaSv8fRnYE3PIYb2Ow8+1f1uC7oJeUIapMoyEHJtBO484f6cNiVAPf69V5swxD0Ol2xKS5
meumdKlJH8GvhYpLWJ+3vU+AgmrqcpEPC/v4CB004DbrJs4zTHLasnYwBIbz1zaIJVOOkJ79bOKT
mAPuslgkXI30O3Ev6ZuX57wI6xnMKz77UDgzFNm/CgUhiH40tGG61xCDbb578P6Ed4icNpRB9ug3
BZRlVlCl5JHremDx7zhh/KESimcPebJPLlnoM0xbBySc/vyG4dNRv3XRfifPX6bOfUj6fG1tHVUe
2zph1D4oHhz/umNoymzEGx9m9NDq7WlegYqyxtHvZUAk5NDtifOLVd51CptuXj7755OTMCAWwd7a
Ao62nd689pntHMJ9+jC9LX6fH240hfB31wu2F5abmKIv+pmWYITHIpEvwnIiRBmpLgTRzej/npT4
XTdRV8llSU2TJ8PxGZxPJaYKB1vVI1iaOdcz48tXGXwJhzyhDuX1aH2B+FiMOx62vHxF4YcrO0SZ
/oXpFCsBrgVELA151kKLdhoLYSUZepkbuTvbqNRAStbHWCM/vQ2kNrIJtH3sLkCNANwcda2pLSjf
2MIp3+h+rX86VbX1dcYkMjfrTJ1LBLTDPtehEuxqrp9uykBWJpJYfGdoza5dcf6LZt3HZufSbSdY
VifHJy+b07HSwgp+yDZVUCp3riI+wHAuWYEuYSGS9zSvexXf0MmVeiSSpe3lrQz6riTKKmEFqThB
L/1YLUBFveW4A8o0nu4N+t7ShWmqdOsglU+wTB4SulgpPbc1QyN84OroqG62g+tI5dMvR5BA5LPf
yrZCiFVaBqaRp8tcSzkw9V+hQO4L1cGLPKDr9rEz5zUgvuUtiauikkutzgJBB/ZW+h8xiEBBUlzu
eHOOI8GoKZ/LYiN7RBMrAxWOZVi5HntrdAMkXpit44FSwDMj+5GMzBXl2XZen0bChc9bKoK6THBa
4MpEPBSgpboNlSgVhfY6XZJjR4Ur/ZVwTbVOXrxvyen9iL+D/2zcSP1sX360dCaSo9wUuTQf1r5u
6J2ka7r/oOW92W7YEH60liQ6gbo+Nk2vRXad43CmNA6RbiJFZ9bla4+zyYaq8QhjA5E3fiYPhzgp
6DTIsqkKCqWubOQ5dZAuwObcnAG3rq9qXwc2ap+PL/U5T4ALZ9+LlHaV9S7uBnF9L8gmMduekvdF
Onl3qs19l8i8Rn9kfvK+v3mFleqUU+T8PF1pI70f8n15GMP/GkS5rha6bSEIuty9E/9WF4VH/SaR
OCVC191IxAmlyPWpNC/UE93bQUQDa+oc4grr4gL5bn+lFPOzym+mOkflhU+6uTDL8PMWJLruiOtB
kWoc1kECiLI+sEf2PPZOrUxBnFQf85j8ayOTuMHn7Ehw2jET5agdxNAK87qQqaCggTMx0tKaLFhE
cbw5KP8aqsRrSgwH3rZA4TcBvdmjWBI2i7wAQuoI0RbYwqXjqBSLGmOf2eFNpkpbWbLb2a5iFhvf
Mb4HqQF99mXglhoF68/n5OH/J0TKwKd2HvY3sJunLhNnf1uRCgsHVYs0TjNbpNqUl7GyGmJlPwB0
PuQlXDVSE56LmRFSzxCYsl5X6YaSAsZAQVXWaS/fSmBYX60bRSNaJjQf+uNiz8ueoBf36pMpDO8p
lOue9H0rdKygeVEfpu4hf0IIrFu8TYQmmFjQARbmGlE3byrFL6ni96D89XyZAiP0KMMXeZ2ohmsQ
aWCPWOmvkYpncAEU2aZQYzPTJUdLjs11h1aj6OMGAuOfS0MOLXH9g5mL1gj31TaZHxRZ1E/xNbDT
oIr0mEF8RH3hjueEtdtcVyWuDTulrCqVg51zi+FKCGjs8UdTgdPePCVZcXy3aLkuO/ll6D3WyeEH
Gwqa1nS4UY7rHshATaE7pPnvwRyXt9IrjGb5fsc1OoYfKQYxCWYHdoUcG2LW4F8I0T0VE+NcxhhH
PXFzUbMZqDqgS4KOfRG5u/HaIQ6msrecgRLdu5gjIEY/MKenRtLpel27ktnrmSweYQ3YJioH0FFo
BKKdSgJdcMfHak56u2l5Btg+1ZDnz9vp30vHm5BfS985rLT66CHVjTfInmBVTVAqcHr/snZ3C8zD
fvBTOK9VcUOevpXD2QkTSzuqhuyekAFZbs7H8VGY4rVNCWw2Q9CQiYqznV5+UUx+HUwfHYc3e3tR
f0ZYWHyIO5iE0I2s4BJLQv5LlgDtlzaZD8ZLVvrljmS2eNVcGwC07FTSjidx7r71b5h8rpmQOeEu
gyo2rTSh+W5pz5fcuoDYLxr/p8KJZWvQz/0OXC/dnzXMMyWZ+kWTFCtBkAAvXOp5ja3DCBrnkBPu
WCTWcfgOCNjSsnFVoSc9v2SlUX8YRVF1w3EqenDu2P2VVht0LRsE3g1en5jkwH21ABz6p4ScQIf9
//kekGykNV7UdRZWR7ZG2G7I6xdXYZZvc1atoL/uVEbRUc54wfPVHxBmSBj2Y9zXEyW6mP39kRmC
SH7ex6rrZXjufoh+suFu3n+Pld4TGpgx/asCJz8Tm0wJd4bjjUZdV9k3MrYYJlWOaycyCy7X/HtC
xTgxqMZRTsEv5XmXlN8G8s3j8XUAyGGCOVWcFE+FttDhxlXDmjq5tqEAyan4ANcUycsDo4libqAu
HzIb1tZxUyU3smlcWHulwUPc0zuXCa3/K1EdSIM7yLRiapD4Wx2hlYvbl5KCrWNzuhaTzNq4Qm4e
zUoTGJZI0QnWbgB0B3QvLHERt6CQ5b6BZiPNdDqKl18WyLWUgguWOxuLPOihZgPN1xSGnT6wvuyv
L2/V+NKAW06SK74zuT0VFVXRthhWbsYB65u7TMTBT0jgEs+Pb85MBrvQc0zI4s/d+Ga8Tu87H2DC
w6QRykLJfjUaxQxBPyf+/IXrRP6rSfk7NfagyQVbQrujKs65JUKsxFeeeIYC3Cv6t0uhIdwwDkAG
r2k3QfgcpG3qQVEPUdkvkwfqV96qptB3wKHjRSl/LAD2wudoTEIsrMy/ssEMxbxi0viLoVsrhrbC
NkSS6L52YQDmcGlEky+sTfMjb0eITyjGORaqHWJzVCaMNFnfQUbgPbcSaRXEXD29gRA5XP0P3XEr
J24fg9zmLnHC9T/iE8ueXB5mG0J+AQCqor8EOaHrvSjRZ8VIxqQ/IudvWAOAnf4CKGHmpfvYL/UI
APpB90KC/KXALStfhuazXgKizKKtWl3yTBO0llBxrsFCmz/H0rTQDZ86BJXjOGOODV2KMBzR3Jt2
gbjftIXD6vvh6k+xzZku1X2cfTbfAhC0JXz5wHzV0xx0cuWyQrg5nXG8wlKIF9lAAKxfj+6iH+qr
Lweu2/zkhct+qsbcyHWSYDcaK4dMUnCC+bQD5zy8g/hBTPC+MMhGei4YO8QJu3BWGr3IAhXnDztN
WACm3i0FnczcIk47Ru3qUcT2vvKoUW/Zlu7s/S53vKpeCcnCnUBwXAvowJgh+t4jqW5gDveiE+cA
8XfFCfepQlg2QIYnhB/r5OsC+9Rs7zCg0aLXpttsOzMW4jAqZgmTcXfuacaNcCHAUYf7WEmCEMnv
UKGFLlXjDV5Zyp+0MoYtF1cwfbrJBIPoJsMSmRZD/uQhvLsvYs54jReWUAOQfyu22qb0Kizfibxc
mfFYq3LqhukQm1uoMQdWfwABvlkLIb6YS8hjiR380L2TxRrizruAsYilRzVNgj8A7+Yl+UhrDUVD
hYgXgzhaqVEA0+Ol9C9ycPlCEqMO6GaPPgqOWDxrz1OVy8UHmml3WfAV8Reyhkuq8rx4aVmye2N0
yELEAC9GJ+HCvuhInVhInTVCdqtT50NDxp7AVbgPho46Awd+pdp64VGa6rLDChJzIgbf+s0e1LK3
QFm2OVBkzlYfupM1JkbNOcILFLHXZd2aEYp5RJyeWQz4apKF2nsU/tJICxVECCmsvxnVdOWVpUwF
R38wfLtebJ9D16bdgHJtwyeHOZgS/7rdKo7QGpFH9b55QsthIzkvJMb+KNriISEypmUyHXrp2vnC
n17CHjS0L+MVI718t0T8d3Tk7d8e1WVVgOvC/qNbopFMxb3IRWp9TmhV44AEZUzK8oqNhEo97FCl
EhkaUeQQDajmUxd0/2yIMcIchaC5O4yN+6ZbS+saCcqt7+OuFzd8qZsaVI2hcE5pILL/klEfHwdO
zEfyOglpMghc8PoHt5C3s4cbg/hP+GQF3KCDpu5o+UCGlaKEvNgIM93HOgDbF6l4hg6UB2SyXXte
jW6VnSIxige+6IQrTqBWBk9yI6BHIoX0kAchCZg6Cx6RiLbzEW6i+gJ0kRmKfP9FhEFOAO3SfhRG
DHak9Fxh+dG2o8Z1mRB+z8B4u/iPF3Ini+pPSgyqeEJezDloU1qq4rp/KBtdNVVptsQ9Wz2zqXI2
jJ7KpUGX1iXuP4VWerwB2x1jPD2TPgCJV1Yv2QxxVKRbxEQdeCuBHDPM9k1ak4OeixPRiNC+T5Ps
QDNVxFnBtOFTDnUbVelkvfTtU3TGA02R84jmFqxy0KvFfoMF4zw2RzNbwbtXDg7zESCj96pAJoFG
WXMpMtTyesbTR29Mj3Eho610O35QVhwJzENJ4p6U8DzJUB2CCQiPabH1fLh9xOXs6rwIF02lUipX
fF8GjLXpY2ZWEj0hR2dq4i2b6S4lEU/aC73ZNurFcJm8rd3nxSleKkfkDw1cga/Iweehb3fEpnFS
ThAa/a/ABTc9qUpYUfNq5OYe7B70H5HviPZzWzMZMRZZ5cMEP7GPlhjpEuJLkCfkHVdx4O8Rc8Os
Y3PH6rEeRjzm44vy5l0iP+eX2TJKGYmPngoL5LUEa5U3Vs7mqvI2m8odH1s+pX9r5N6kFf7FxjuW
kExPfzIttWUMLMPNdJ121I3t2aZvTx1FG/UnYreux+NjZ4Y4XQ2vTdUk5xV6BUYEAsjoJItAzIH9
PcvVDd2WjgkFGcPir786p0ErP5PKD0ZuOASEHJ/5VPD2Bcj54lZ+nPX5HHERo5q2DLb3cD1M+WeZ
cCvrhvRjVhwpnfjX1f4pxnZwzmfiO2ArY9KUpwxM6h/lvwMYl2nbsXit2c4P6H6JDDpO8N/P1z8L
IfizzI72HlgGdXHg161T3mXRNavXA5N0pqOWsAwJG1MHn5ChRcpJXpe88WrGb+IQxgeXOjHNgVq4
2bekd/m9jv0VP3KXRXBJpCDCuYHrho/MvfS2XNf56wCHPxDTW8Nqp6bN0X6Mu1DDWQgwiyjCVndW
Z+J5zUeanMICaXUrD0ttOXgXZRs0iGC5ei709s/8fDj5U1y/ey7scPIEJeP7PuvHw8UW0Zsxe+nz
/8ttJbkEsRFAICHqsertqRlQNCga5QUMKSrqP2K8/PC9awv2Hy5hQYpjWHAT05kFPogsk6jNzWEX
c5dGWiDq6mDJl5r8NBlts3JiT/MbfiGeWJQavG7fhTLBpy7+duynnZF2Ng5kMCYymokl0NtItew7
u6Y00epUn0qhEIwTDL6JUoNV1iAGC9cp+nSWe1m39p9aJuv1btcI7Nc53HtI7tQzrFhGNfmuNzRd
5i+L/yBMT2eqqbC+ph7zoGYW/mD9ckveHc+BTeceNWs8gR8MPs0w4tGCU3mMb0mppJBpl1FB+7d/
H9qZSjUhr81zWJ7ioWojPvQCbBS+RM0hi7Z9JuFEHQANCxo/h8WfmOad+pF7xARQZA6Pe8+x0fAn
9Ax9u8MBz2G9mFtg3uC1To3zGhjNbzT2UglqkjqdvNCT049t0CpI2ABGrpxhPpXnmTlXH03WGbzg
9YLeFAP98MQNlHAXMiW3TRvVJ+t6LzRBMlG9ls4xEObcPgMIcesCdi6VCosgs6htoE7udoUD1LIl
2mZwhj2OUqxxJU/36JMQR56kBTqUiYidVzF0lsR9dV1ocMlAtng86Y3vWM2Odbl1FmGgXjWZoaoN
AHO+Uh86w6ejY0jDrlWKASxUi7DngnRthxa3Nk3YwFGTuIC5Ic+yBU+VGOhuHzxz2tnvY/AxL1de
xWaDPyGTx+2lACFXW/WMh6wswDSbREa+azTq+6vvc5GVn/LP4vYmZcXR9aRjsFazjVT9TadsLVx1
4zGgNnQ4zYFghDHfij+wnwGd4lXK82Ay27GsryvoipKhKqWkxX5WeMIOxjWG4XDR5DcW5TCvI/4r
wAe9kJPOihSpWExNTX3qE7d4+xIhQEaMQPS2Vi8SetE0f/kqgYBMp0Aoj4JGbq8VUFz6b6TLKERl
DaImNgl662k2pvt52tJxN8R3RIJ2vy8/ZInvUqtdbrkFhNWsOwreKSna4Kbz+MhQbkDgLUwWNcQd
OWiHRla7snPbBQp4h1MM+7cwOyuvW6dSFa4g8bnFADhYoAfiUDbnSc3kt8Qigt+rOhHYROnnaqRM
UHnCHrJbTJ785Mf5xOfLFBdhs8msOW6T7q0s5zEHJMSPhJH/x5wCnc6wR0cgw9YxnsYHiU2jwZaW
MlwnEqe/N2I+rY4j7o6MNh7Wxap3WYaMLgQcNk162jdmvK68qeuez2c+Qanyx8F+yrBWHE1CCPUV
97ecD0uJ8QV9XAu5HcE8LUedx/DDM1EJL3l6x2q/85VZQXPhQxpxdtfPFfrOqdqD2SRH7E5axfEY
cD5vkE5uu+ZqWZI+9eRgdzgWwuV/m4nbfmAH0lhr/Y2dl74WGRU477J8XrumBBO/KXHpZHjn1jIa
sgkJW+RrRh/nll7KoE2W6PiR+O8V1N+oadUIKi5GcgJ6QXuH7Nm8PYGjwQFNnwxzOwETI+NWrQfW
UGxXwazpFlAQVqtRLpTeiQe+bfNrmNt9j3KAuCiO75j5aJ8aCs7xQ6XtpaBNVrEk1+QZQWkPZXaS
vKevlh8KGUaUdHgPaJwnyxfKYvc6PS6zELm1JKHkwZczVkDuWmGXaNCJNxrzENKpoBxDWG9f5h6C
U1CkAFQ/lz6JTDhfBgGCAud/4NLlZ/+95yAuUc/e+UYIS3y4i4qOfEtGdiZo/dKM8zb+Hq1x1hhC
YGzfNHecop76FioaUooisVq28E2XsEHlQIvKv6BXIDvjh/HnE/xfLcWVtl+/W/9aOQiehvjEcEDi
/4Jl0NRSG3+NF8p8SktmjfSTyu5GTrr6GPWabPPpJEgSJmWKiMAD+Joz/TAxesizw+ZfjjTYupJt
9O1M1IwvFwqvKqiW7sD29w5GdOd6nhOjx045rs5YWs1hwi/QYOuig/N2b4vFMcoHVwpjDKkEFCFS
vvz5867LKcO7UWfdm1XeGPGQ0E8Mi6e2bV65Ok3XmYaiR/BvVvjZlJbqkFyeQ1jJw1HZVmY+ZijG
FHQbBQ+7CuDKAQ1bSgEdShA9xdhpLeg6OWDvb14yKMHZk1Ol92TsaeGQqfOJRibrARcphH6Rs+ri
lm79zyPLiuIMued7f6UDtO2czRk0PJzPmNDzkihEIOPGNsd8w+HCGj9oREEtcsjYYC+LQlQ7YafZ
IUPvyng6yoewG9qnHXa7LjzzZlJ3OGX6mJw906GPcx1NlzgyLp6wRZR4cFjhmADntfiLAc/PlqF3
f8BDf+tXbs++k3t3vMSh47rWBBbWMZ7dbUr0o2dqsgahrVFWN9lHk/bDSTUccCUxXODrD+wEl2fP
cgnK7mnpWPRihjiJo7JTIVbxeIc3M8TvKWFEAT1PgN/YZ5c38KZZ1X4t7TdkXnoZwzUrdrkYuio6
uQKFIqWpnZSidoGBZn8xhUXi1jlLk8jw+KVlPbPmSyPpspdl6G58YRymu2wgYTbIcwJ120eGeNXe
hlXkkn8itJZoP8AQQNjeDV+3ZSFAdU627JGLQs9kbIL6EESNTcVFAimxu8YG836NRtQuQTRu+R55
s4KLyalIA8mhf1pI04FIsmE8oldxHa2jmM4f7ZaD0t7/N4LxA81R5ZRyhTWIIIXTkDACWIwqA32A
FSofYicOOwaahlZtHqcd4oJL6CvzNUOPj7RL726aij8arb5GXx+uFC6ZTURkTm/ReTs7CjMkupOI
BvFe7C1CXGDFWD4r1eTBn0oaGtl4ff1YC8zCw6w9vCZNzrfK8pj+cMxfxSchyHu/77xfMq8aowPt
PfjENJdD1xuNM8eVasdI6GuAeUsClNDhHYE6uzYDC5PWp7SucTqkd/T3e0NxBZoh1s8nAEYSkVO/
WgOAJjzrpqm/WwAF8lsfLIOUsugctZvnWtM6YlW5ma48H1Z0p2eBA1yu2BfQiixL35utrouZeN4p
Vn/JvZOyD0PNcDPrLslE8uqnEH2u3HHVa53uba2ykTKl4PFOWUOvFtIJKIOUMdTz71NFRDWMP+6i
U05xaN7/YzQSQBc1kloiwyIMtdkpH+nkqTMDD6oBKRMuIEGSPe7v5W8wOaFNv+C37rC0BaujSv/O
ccAL0pZcEt8jvYLAhTOi4AUGAoxF65MAVxeHhPapiVOPjHy8/ZFIJsjwXGhTWlD7NtbhfuJPEJm4
rQb7pJYlKZb4g6GpnEDITYvV1uVAVc/jbkWKhnf2DKEGL3cODQANtodsGOrXGPUzG/wPVEMIdzlE
dao+yD/VHXkBekXxzqHoEd0P6QpiZYvUncrNNgkTdldJopffVTugLkQ2YDNUcWPAaRQ3pU5i4Nb9
F7LTcqifsCqCOkv1uMAQdgiQomO4EiSJABLXY5qQDPh3/vxFMECl6rxU70tCga7uh7Vn8j5Pd1gt
sCNYqetrS10GFUM1Dw4aVSPRW23bpyHcBJBMryFiZ7qHT1XBsLXetgYa0uOjKYGDVtKXmIU3EIP6
p1bIxxwVzwR+w0Y3jZHxNSyXBV+a+aOh/bAtwFK1KAyAa7h8Azl7ooDFYSS2pemviKDATO6J4acr
PSCfr/LEkuCRDeabjU0+pQhkYz3KJfJNwN6LiOZxtxtuakDU0seRB2VWdsh0+dwElIsefS28FGh9
uhY0yijF/zXicwirzA3uBSXrvnq5W/DqNtghqoOwsJxjtxT71zAeNX/+2/jbpiW9vwHflNiX2rrm
i4WisMxMUkmPZdxWqPZBL+ebwOgiC9GzKk6LM9xzAEfkfargDsV4V87JhQLgq1uUeYYEOENOhEDt
6OJ+4Bzw1ur2NmZtEe2s58+T81o1UnC2x+Q7RyogUMcSusxsfCzwuLTDQQICAMQOcH4LfOW+nQ1n
Xo8l9W0nqRhkQ31qRbWG56sy8tThYIksuDrb3XfNAJUY0cIVWgAa/Cdo7BvgBKEgo0Dl9xWPw0WK
AQFl9GkOFu88KPpbtbOfy4ndVyXt8yd3xX6Dk2M3cMLFgKlPKrBYG/lIHXACPcBlJBo2jZNnovHX
FfOwGR6YTHENa1cYLsT7pokJEg8YYkDdOjteOhV48Aet1BlNzzbI0Z4KaMy4YYBR0YcBf4auEozl
i8VO3Dwzx+DcK3o0N5v77BDlopYs3UZtCRe5+B03wg0LHPYfpUMBaXPVKZvxnjU5vhjoI88Ch2dV
fkPB2QPuJXDfFx0IwVm+JJr4+fscrr13qDgtwOS04ce/mKZcNC6xsX0I68SImy3n+t/L5Z/deUr+
ZFlKMYVf1rCvxy4o5bK9iC1TWSoGNOBYcKeDd6ekhHV8nWP7kHrZRbKs5B/1q78v2KWn8KbdrRGi
ZJTScWwiCzysOtcd+r76GgQrQDZJsQxHuLHipyAZvfb39t6fdTI21aB06buL8rtvrJWFUilhbGUz
T63wF+kBcStddu3W6nh+K9p5OnGtV16Im8fTM4PU4xNhBl/9dTrJODWQExmZt+12B2n9NPhMpkG3
wpv6QNhAUl7jLKaab6IWdDjBpn532r9os8eYVo5n49KKaH+EJqYpTYeQfA6+fTHnjWV3XhJ3VQP5
Fu6EQ6a7ia6IH7dWJhxseWxXO+nXXt3rafx7WPgli7eXbGxmjh3yF7M2BEt16250FPgxXwiJsITs
GHP/qP6Lc6ED+qvAl1aHf1Psk29BaMaIyQywRY9vJ3xFTetUqUwli3D8Q5MYkr7l5aKmj/ymZnlK
VkcwEii6/xD1/VNX62VwaZJ2uHRAtw4J2UTwnpqkL8ec+rMa/EUZALsyACWB4zBJeOLiKmoFnZ07
kujCwh5H7NhKQuG/Poclc0EWqAzddMnTj/tNloh58K3gVT3KMjhEF984HmfAJH7zBSY2UdUtELZf
Y7kgkrspnBr0WSRNkSHir2jyPYK/POzghZHvoT6HDKVicm30Vd/3Ds5lZPLo4hJzXHu6VTLNsTQQ
9/cFnNQwdXN7RAFUb/jJxHBCyyaaEw4k/4W0rXlz9twQxNnLUNDZeXBwddapTy5TOX5pjsQKsIyb
rI05nKjX9uTEpA0ctbx6VGNBtUFQDXuaXFeCk2KkQ8XNX2wTSv2fBsmKi/XNIMg9d2NGxsb4B3hE
awP0k81QnhZGvYo4+KOZQctvWlwa42g61TZaxfKlmgXePL3O4yylXHLGdFbi21RqD9DZS8qTn/Vr
7Ih5skfE06qxUVoyzW58qDzHTxxJElenR2+u3FkcdeeERpipRyrB5XikVWAuY/KRleoUqDqziHdI
ph2VuxL1cx35i/5n+EakMefOb1zxd0z4z3ams2ayhxMCWVUWhoDBpdvgL9kBZGfLmyYbsgOoeQxd
0rQQ8zpHGLFsX5YK76n1IfXOae/FzRui1MkNKZLKu5zZ5yCCFC0mEXwuWwWmQBaSAv6LLr3DQRIy
lSabSyPXCgnW0hx2uGqrJWVOpt41bB97tBoIh3tj/6fbbwBAhnxFPJyAQB21h/UOeOFVNHTEQUfj
BIj+zOrNgs42FiP064KW8cyMAu8JwEz6cZyOPfSZShi6h5C3quzS6LKhTuJ44B6VrGH0kHe0iwos
dypecyokM074dHG36FkDQFAkHu+kOKuUUtAZ5zr8GfTORQRkCt5ncVh5PC7UVRW2lOnjytGb+MgO
983CPHip+366fwDCQfMwNVUbopSdaj/258P3/H8AfvqToSdznMgxExEbv6lKlgshVT5I/OBAJ7xh
LWsBVnslPv5DyBAzV9ht1YXAD/Nly92ceSiON+JdKwaERwVQlJc4TFS4mFAxofBpgjn0SV4xW4kz
CzXwIF82fscPdD2sDZ/xbG+XAnZOi2uJmV+fiWBjBFK/+A2JtSl1Ofu63H1ag16FZz+ZsO2pXLbe
iTJiPjYTG6+Q/GFfg1yNr5zNEhS4JdmFMdz9tKmWa7VALoCtSt4KsuYnQodd7UHFQIUB7QZ32r1m
uHRCA9LJY4B/TJxXznDEflpZwvC2RtOt5KFtJZHVjVZopyNjQabnegPFy5KLKZdlt9E4/6yaPdeV
DIM9oPe/TtlAmgm6YI6MChlraWP78y9r/1lVPBuma0tcX0Sl0vHJ+sMerGOi4wPqZCb6e24B06fr
wlKwVHFx7EqHdLR1NR+UBt6fGtGO7ckEyQFPDfZggXjXC3kmdvE/y4zDw6S+QKjsik2ilgtUKAXJ
Ln5CNYbCI5upH245NzytRf8CviPKitL19WBdviM+xUXC6zX/miyE/+wSWXwswHTGP0Ztalu06Yx9
5dFKToPT7ROf/ffW9BHjI5lcIbfIlE93n1psKeRXYzTJyZbom+MyexUiY83I/ypWput04gq3b7kd
aJZysxcZVU0VlmTXU6VR/HhTGdvZOwfM10trGR56hdpFPTw32LzqF5SPvZigC76XTGeNwijgFTVN
JCWowicN5nnZMPlaEY67LHGtS2tjr62y8Pc2arXkCTG0Mn7VcTp33pvrWq4Jx+06oMmq60SXLkso
mkF5OvSJZNstldiNwbgz3Xma9KDNVr9WtjWw0/b7kqwaNKcFnShq0Cphtts86ANujna+pbgzlle1
sCxE9SxvvOoe+jD1KfEotB/Z8r3HjRA4H4fPqzGvU2Wvtbl4+4FvJ/a2q9kip7EmkIfHn+xjsmcI
rwQcFRbrs1JpcIVVEZTjqzH/cF420FfP8jrkw209RSKkugF4+1/KS1Tm6OvQ57/YzjyH4OJmt51p
muL2ff1UD7jawh5A/42hUl5DDuj3HtQbYgUulzO0rGnRiIXUnHJq1TIYThOkjePYP133eUpguQG6
fxsN/Mf1wYSlB2wsz3PT9+4b/EM1Y/hwzfPd1iI+0MJyDqfhCa/7erCvTSBN1G/wZxiXxLca/dbb
3hEgz7ROp+4F03p4CC5biYzHs2NwmnsyjmCEaCTNdELIV+SEvp7XpjRum8NpfEv4SQKCrHdn3jt5
rrdKL/+V1oXsc3iF7FtpITnbchVGaYN8NL5UOPop8/tJDCj/4WPu/Sf0I6fr5lsyaCBwTHOKc1uT
qPjkeWX5Esz++sqAXqWsqrub78bGGx7c2MmeSUvYKTUjBq2Ek+pk5pc3NOU4D3RL/SAkGkPFX34Z
BfMebNNNjxKKtzJhrNFkJfsxpR6IZUiTPZoI2Gl95//QvtQhqcizSPaC8iLNaqM6rH4tXNyVztj6
6BByUWvu4xHLr2uNantXCOl1S6Fc1sPbR01/oPl0HwQEbK9kGCPXlx8McMTttDe3Jz/K5vbsiph/
uSn5WVJWwepwhOyL0buEr8aRaIbcB17Ulc10eadusrBH4BdMlxICAfsOB1EYPrOgDRZ1y+M8PDYD
gZ5ngyCvdSbi/CcVrIE0wLsJwx2TB3OJTJS1MHR4N0/9SCDOkCqniJGTkGbXrBneRIEGKKjdzxWk
kZz3BkEiqZP+UCJfZZKU8SblfgVNQtfEMtoE6HYMD6FnOAWHwdMLYCqj5ZlbHxnDcYKEOaFzm+LE
HhH/wN8avNvqmoGxDKfOLWxKM2BVgNTBlJhz3w9Jfx76ikn6aIYopR0nkIDuNLv2leyE/xAHy+iF
+/pMoa9ShYjTehEUFhI9x+XkT1RGdompjstm6v/mRH+DHbSukQK2nKcE96+N+dytXU8YYfAEwyVK
jhaPlVUr6pjNegKMskzT2qVFnjVFpGZNGriSS2RAWM15d+EGYY49HbR2Uu/QivsqmDH2hbDlysJY
rUt0z1UeII/iXwxc8th4Md+ecaRtY+T2Itr2ULlP497V8duxbDTvnITnBCLi2CEGCHl2hTJ6i0jB
cu0v0Q4UxXeTIOFaXgbE95eRWRQHqIfRMWs7RR0y+tpXXX+IwVQUUl/3rQ05r1wBoPw5KmF6y//I
dMNrkd5FJia2IHzjIGmqLxI7lI7R93WKWGzrVIf75+/J0YdyDMy11JaMLe/OWlavw9ziPxzgZIbh
dCC+yWA7JDzmcOLiWOFqk2WvrMBD9RxaKBe/5vNVjpeE7LZl+s1Elql4QWSJ4cLsY61/MO0hels2
E9POGsfOxnXF1dVgtfNuHClvL8/L4iWaFOvpk+U1H42hvXnO999J0qZ70au3zoLinVcTY2Y5Aq2F
zZ3ZCKHBO0uaS2X/ErujiYChu7Pr95At1Qnctt7dqSkiTukizXIsb/XaiJUvAHYF0+NysijoSKBp
+HfC0FDML0ctIqg2kpG1O4JEBjdbtVaPcd4LesiaAqveOavmZJERKX3fJ2xFm2LHtCT4CE87vMMI
Gq7xv3SHB9kZO26qL3vq76PEDt9YJn6ct137TGWGLz4WN+vDgiRDc5IetfkWcrlJ2a6Z7zEGi6IR
O3xCl/shsQUUqfn55jBdYs9rgn0Q7Zb2Gnu0623Y0yOKnKJxLQ0izdQQtTx4tVVOHkeSQwoRzFGO
IU0d2GM9PYna85arGt9TE8bzQb72n5NS8GNnrN4fQoXKIHqiPAKFprBIDaCSbhOECPWvnLXiDWl4
F7JTdT2/WAstK+eG/Rc6Wo7dqsf/CAyUJ23J9sZrZ0S7/FF0USAzmnsi28XpSHtyC01M+TMCsEj6
KI4dauTvuHcNSFKsg8HY/J2hqwLOznSeptUSukbiMrbFpg6buKOGb0sQ24ZWDbxq6hhkn35pjk05
Endfc+3ac70wjIBGdW8Absg4d3XEbvFWdLZUQTNjwVSzCzW/S1sP2ELNGjQf0gbBG/yYaAFqbbSi
+6RklKw9beCVdGFt+p93W87372iSlJHIZg3CjSWTV7OKz7btuzFOF2OjxKZq83iBS2010Cuna0y7
zIate/ULuPHmz5I/OW8mcx9oFISaFiQI+lB4TnAJqWjtDmGgPl9WD4TV0tHbPgQ0HNu0vBWKMVmL
xkkP+eSe+2KMmSW15Mv/AjdMjjY50mItwDTZw8q0FjVzkHI+1aY5ws2cQ+1j91Hg0993a/FkMaO6
13a8ew+BGzcdd4C+BWupGCwEPv+ugs4DCZWt+QdEujYN1k6T058+BNL+sg49yquinxAbRPN2xoBf
N0cKf3Nsp3Icvtg0c35xMZAQ7zabH+wv9DCNCzj5dt3rh2BoLb+ncwhXX0aeS8jh/AcuGZ//swZG
TnTcgagruJnc1MadReIcRaTwoPD/nf5wGkUaI5UzVDMIxxrCyX2oxn2Q4zWdpK2IhK2ZuxHWgl7+
1nzQUFtZB95NcQOtaAku0LWi8UeVR68Y9Z5Hkzc/pBqlHINyroIADpOl/nS9THfWzV8sGiPUuH8E
sBGwbLMN/7rfq5ngocdLOy5dvLqoh2AK5ocBLHvtTGOH4wThCK00UStBbXjnGfprHlUw+Pcsrr7j
wHk5lKrIlOPpxOu1bdO1HpzGggSNCIyMOZ7McuUG44vj3CXE0TCyHQwmMApYBd+g45SqSHtvfZ5Y
Gk3ahNpguSvg6mRWVWxvheE6G874lyc9IRDeB+X8yTD7a4uzJDOGVAu8fx4Azk9RpTFxViYqkICE
B84EI09gqtlk75IsoUyHQ2ZR+z65CSj0YG+KCuvWFMgtcJK65Il3u6k9FMuf6dx1Y/CErozSHvWC
MXfP5sqMaQ1DArHe3bvdSMEPAlHj1yUxJAduZYv36Tl+Fl4/JL0nYLAuxoKHqzVelb/C+G0L40+X
y/9BpHjEy0FXr98SiREkGbly9qqV/OjjN03wgb5VmGwn3ItA9WXli7Nw6xuoDjL2mh+U/Bll+DHz
1xkHqttdBL94PTqHYToaniMSE7KtdvBx5XkIJhwQYV0C/fldneT/5iRF/TrpTC3dlibvfaGtRRCA
xZq4htV7oc38+dxtJefxjErse3KXyL+jFQu9tW0ahoggcNC7gdNTLY4jECHqozcJobPMEG+sNKEU
l5QlelPgDi9K2DvQRYh6gkLWxdgViD7/bYLp9i7JzOWIj/qtwVjJyH3XQroE1TvkQZF88lB3OeI/
F3NQoiU0vnZ2tZVKNxgqHnIjn3liO6cByWO1obNudQDs33nVrrDt4TjjJdK+m/xvFI71GSMu/iBJ
6nJXgnJzplaR3xSoyKLUFHzvqmDC2oB0W+vn8pwc8ZTcnovKS8JL9nYQFEOPDAxE1Ro4XvvQ1K8G
9cX85lhCSTkpsAe//niEB+Ar3nNnE/i1L8d+pvXDTQE6ePI4Rsvdci2H701LZMiGu1a43oF3gtv7
DsY0yMMx4P5PTEJs84y8O1IAWUglI8jHXq41xya8A5VBpLnHIE23wSfjnxr+/CeG5LNMDTDhuSev
R9E8gsBk1GZcZ5bXq5e7hfhRZJ2nkZy95u1ce+Nm415FzYbTSKUL91URGxIYYiTGhl6iK6rL903m
G7aEC2cPDtz+lsYHTv31YhESRc8S2AR9LcdNG62ArT2kP7t2CN5PGKwh0FusjSKnyrqCAMNL+KM7
qGNYt5/3xoD8kugOLTg7e3PsaHLiPx0YnR3v9kHWg7IRY7vK+jpNipGDyLvNg0GFRoM+L+OPajQ3
I0mz5jDK9NvLAsspUkw6FtUGXWUrHYlv++mBiM4KNb91YFYxKpgNc7YEHfeZHsMnx86a/WxF59b3
/w5BSk12fi/Kmglq+RpGH4c+x3taNQI93V7Ak2ZHa3v8mnUgfRvDAP0L9bsvE2uq08CmCkAQXEMY
qFTZvpi7tttlx4Fpb6150396caM73s/SN/LDILjQk5ry4wD07PEcG2ivntuoxg9TD1B7vK8coWAK
JLrHY2Mfpy+62iD992ZsXXxQ/1Q/ZbcBNjOtrl6ciWjNCyB/8bLqc+PnZSpfuqWoyALvpHi02E/L
i3z9bYvUhLFJhQfyK24WtvS8NzD19hi+279D+Csza3ftJKKCDMPcrkGBYqAOdk1ZqdRxUNuvEUwj
OjEQNetC3y5q43/ygl/OylLuUcAptI1CnmFULHl7LzIspcel+6ySiWg3PM5iBjx5zaiRZaJ2fQgl
iW5fZRdgGfCDGay5akYnvHUwkBrxsqqm7ryNLz4WyZZTsc1wOXgyneuFmmBERDd7Kbl9Qwizpiu7
BeMeyVHVKeFzTTEU+0iKok/9FYR6ritE8AXiza1tyIwgBtofFjkFOrtXHu4czrOk60OGKgfPMyKS
pQ3UWC4ZnJRgMMEHhOJ35RWEquoGdCUQ26naBQlK6eW6seODo37Xx209U/NYIpWjywIJPVuf561z
atQ9Dva4Q9J/O7/q9tE8cec6Y/aKoRALUvoczPCbT9+KxaoETfcYhSqLHo+FA3lP3cbNuinjUSH/
RQ9VoM4u3AqqX7JRRUvrm4+h3mULg3oIyaQUX8t/iGTSRUtl8pxJujgRPUp0bJg4a7JDH3V8nVBa
tjJdHNVTiQ3nTGnuW/FEo3sTF5UbCdJEk+/WznWV8TaV/UqbSCbyPLFP5lqv0iNjd1xZvBuQqNMw
NkKStD/I3c8lQxDtuWHmfE1Gqw6IXlE19RxpSjaWHrvX0vJ+MznYcWcWefFErhl6vWc/+IcwLVQE
fcWSf+A3xQOHN53pOlvYvUXtPcArWZdLue6b58KO0T9MBYP7Q36qE8pAbmsbNccH/bY4Tu0ytjjm
0EB7Aw/esgg0bVqxrIBMdaCHq2X6R7F8Dn7FoXrHSsenZaR5WMSkFhsiSftFSRrmP48ZT//FGrLn
nPdOQMjnmIeMVXhrdBMD6mQDoTySimPwVVmmD7plAovrlk8EVcsXFtZrxXjjqdSEm9C1yITLbBEh
dD/ZOXe6pFbHesBi1nStg/mWirTxYcYjXK7AkGzqsU/nuBlEzWfNEbYtOp3U48hi600FcX7ojvs5
u2ecfjz0wBnlTT87VZv8+vw4IlzKX5D/OuGF2llpx39O/kV1J383AXYAVcRqo2T7PYmCstKvRE3u
amBAAnkEZtW37dkaJ6OXHvvp88vR4ywjVLP68fJnHj/+CotBxe/4zOv2qpRFzT6sJWIio/FO6ww2
lGiYLzRsmFWhouEMaIgim6z+rlGiB987vKZC9bHGyR1RfSycDUa1hGinOc2YWBIdOCH78AG/rqFR
VN5yMeRpdkDCCL0zeMQ65SfaMACXpYdDUvC/0LMY4YJm5URAimVyelj/0aoYgwSSefLB526vfeku
Pc9AZgq+xMxwpz4g9amVsDoTsYab8XdPF8UggP2/4fFLv692NGElv/8COMQAYyw5WMdDBRMxYImA
hX46KuLfzCsU0u3HtNYdSdMniQ1ERkDOL6/ApIXLd4n5/Viog60Ssw7UQ9q8UhqbnfQK9hKBiVrS
a9HU22FXLX4OEjh6Nzdu+8jl6HXTDGToqQ3aWonhL4d0+3C5U28xI2sQkG+xYrTyIA9g+YXPVlkF
SVBRe4vkFSgX5dZXxttNiZZl9NTFIxaSZPPAz6XGv/gfOU1dkVNusqNKHEcSdTg+H251GJIwAzQT
I0rwGF1O7X1F3taOIMcxBFWbSClPeWC4jqR/3bm7GeN6E01TEslgAbYn7Od/nevmBDL2zzXpByqX
5feNJe8J+79JVJ087KXJhzLbuVAB/39qa14MvAVrEYfp318+I3/6Gqi640knLnQi5Q8NuU04BKeI
g9J+Effe4hsOfFff+O7iHj0iiJ83vrmZk5bjAFi4K0QPuU8CyBUQRJxETYbcqftYBej/pBaTWn+A
APdnAPAdCnWllqxFbd2nisby8+j6J6IDpKsJv0gAPxVPxda1hN7M/6gfWBgxDbK8DsZree6XC/d6
/oyqRlEzG92Kc5vhYmmcthYomY2UlFACDnJwQ7p5H59l/FA1joFWVaO6Dk59enJxF5UIYos7RYR+
Wk+K25ysciuDGQWtpyxI57MHXljqPGrP6crMkeWblw3hR3BxXEBqon/mWRfX4ZCeS5qfaheilIlL
0s4md+rqoiwQFietnU73j7+LoRfA8iSTLwVOMmT/PzVWiq1bQX7kqM/p1eTkoLDiQVchblR0xJAz
6bPrqS9JgcxRGcxgUBF5AhICP+HzLAQ0UqWqq6HWd3ha4P0C0Js0sRVeRiAtXiwkVXTdb1zu8eWF
vx5BA9bn2bu7STw22+XTFsK3i2u2hDXETjv3hY97IGti3DHyf/N/IGvWiljviQ7qa+HYB5CG7LLO
rwLFdlzawOATCirFstXOSnXSVDrrNpwBsBKzz/lu6yT5A5Ej1aVqt2A/8uZHg3hJ+l83fsh+sLUe
0sEt0shDxAr+CgG05BLXwYQYQIp9jHc3jLPAOGOGaAD8X9GhZFAMWKZcleom6XPGKXU29qEf1f22
DwPbA9D0fiWNUeBah/Nv+Q11uvSoxayZwcn2gLnjGqhz4VqCVqy5jr+Y9KscfT3nJBs6R8Ye/Jzt
BdEGT2WD0U6CCi1thZzO0kr/VxtzehYdVLQi05CkODUJvbVjGuhrsqdJspJ4hP4mFMIqwoqsjirg
hkyRSM6WjTrQoIFilTjXwMM9doqOKliCjbBFS6bIXk3m2qEDuOusoMvxVVZrLwcHYwf3fYs7WV/F
hfkC5poq00RP9biSBmFG4DsHhMzgq7+m7pv8I2y2kxn/QuiNaPtVXPBtSOO6MJy+TbC++cd43De0
dPA/NfpVMV2+gl+8AL0DAGtTWuGtbkTJ0kSEmtBlCuV8I+hBWkmuSGKpV+qcmpWiScyI9U0M7zmq
tZEH0EmGTb61dSkcZDMUo9O5/oN1V65Y6RvB9D1HBswi1UnyF16Hyoe/a+knLvYeH913ezUkkXUF
sIb1Ktd1sdEokBfZmIy8ITRByX1t62W9CC1Inq6HmlAOnXpfOQsKwdFdMj8jCEENtKycwUl/aC02
oqgE0c6y+Bi5LQNgbToNAGoEFC8O5ZurcnvyPMzsdOmoobcMbwC9uYyBcaOJmmA8lm/tZnNAbaCp
io1BY3xILnvhVXyY0kg1AFQU8thjlwgQTymub+0MeK0bCbnq+Iru1UvyLKCWTK80p3qcoTWLfyNe
0HjWLT/lGNCMJonFnev9CiSJtiqp+4C09j5vQtDahImWQj3T8cHWOqfF6W6/Ju8i8LAj/yiAt+b2
/MMBet08KSrrcIlxvlPCk/c3Mhqc5n8WJmAiiGYmD7o5fMiMRuWSnYclFToJbnyAcWOv2GCmVhdx
uGGBvLukGOyCowaRfE6BeySzm8xv++TGVU4XbBGKzVec5NJVcTpuXQLx8TSmAXlaOUG1f4AsL2QO
KpI4WKiO24s+VsJudMKasYYfkMcuhSYDo85Gnb01BEAWp6uyGaH1N6AFAiAbq40qvfjpSatMdgmk
DtEbNT22CNMTyS/TsOBdLKCdYAPSXwwkjak34b3pKQGs9MsTOFIrHg281yd0sI9yCq/+dCz8BG7L
zkGzVvCKOLHmCzLaWmqH8ttltxp1XHnTtistYHlg9oz7bSOmZcXXu0XsqtFi2m2FpgH23Hb0bS34
7FQxnklcZ+3+uS3D6KQ5L9ms1Cc8QFRwH92xtJQgB990/CLyKwrmJChSPcSaRBC+7kLXw8+92VOo
/4/GmaOCck6HW0V2fmrvL3nJr32rQy6FDCBBmxXRpGrjH9U+56V7l3G9H+j999eGKBY7PHcALluN
YPRQ/BKz6qTerq2MlZX6NwzlDTxybIvKKeZhoAK9sDrzZBvWPPBvoFC0s5gsBvwLxe3WwSMM21EJ
4eHujtJuhF6OygIQcRRj/DrbQuuk+1AtTthY+bARVl76difjDXSSaRD9zl39gxeg+qeERPcXjDGs
DOHmrrZRy2bEapCkzFqSuydK0qRA3Vfuw/Vur563qDMPZHUf1P3Qr2tgV6jScYPMjRjx5EvTmMbX
MswMyBLkmYk0uPUwZebjfJJTnKb+7TItBvUSPh5zRFXuIPjcrBVmFhpKJIiGUlg8bGto3g4HofzP
p1Zcp5OqWout+IouQbPnK5215nHhSOvtqEmXRzHFfU2dH7Nr20rejTUFAhc/eh55emH8aNukAI0V
TkjqPNSYvkLqEFPdqQDXrum2FKhvpuZThpaODq9n/YFUJFqe7ydGCa0Jq/xLxF7H6zLzLDM+K4Mk
hj6UKVQH6aow9BBg7BqG4CBEZmI6E4COJHCvDc+TR7qPlq1iR2/4k+0LSIjNQOqAg3XiClGHTaoI
br1o/VYV/d7yKgQCsLKlQTs2vcZa2J+hyOQXWPxCzNXL0SM4cQ4u8y6JXaKNMWpGqM7qRgxKNYDz
DXV6GkjK4LRaje7/V0Lfi+2mB5UxW52sAAo5n0LogWQx1XLZh5FfX/rfZIKwSZGTBWtO6x9elJ0K
KGrEiE90VzqQ6NOyt8QBCYH1eoBhNdZHWs518gIoS2vtrEJxT9nXZYGqqqFMSrdDDgtWw0gg73yd
Zr5dnLtCiS2Gth7fFQEiLg4GMMhDkYdxqUmxjVydQR8WcOmzn0v9HwZJQMn5Gsbh0sdsllfKt+rX
QYz8JIZd0sR0ZGKur1HZjClp6G/Uwvnxkn5Fj787kzvhxjcWjBPnSgqNTLxsBsUU1YVoEOVM9L8T
mxki+G4vI1b44eSd0EDkrOJNnVB+0uqcxWfMXlAXP6Jdm5kYM21Pz1/pNba0pFFdcazoPKlqTfRn
2g/zSTCo3YcSkgRTulvR+iZuYdWfaIYCFffRY39GwOMZ0tWDM2Kb5eYq7gpdli/hHedOAo5wnnXE
VameNqTT0h/cXZp2vXHgVa0vjOKUipYIxkBbHF1t1+8xCHWzKUOakkUv9tEnc5yxVBBL/mok34VY
xvgAD4Vhh7c5Cq17H79IFKU5181aVPpnveEvHXf5g/jqYn4QMvwBLvmqSeYpA+LCuZ9MmHmJefN3
UIdVetMv/Gs9Mi6OzFwcnfSF7Qk8YebJY4T6ma2aLZQYdha7MCM9gHj1MrP5TCdHyI/35OTB3ZVM
idnS4X6DnKdGu+a02GML7fasEp0fwzBuvI7JofDomONiDdZdcdbXnndrzbKnefvcvWmA8xO5CEF0
+62r8MtkuuFqwPQNAPuNck0/YwlmlVFDsc4gmLlbDiFtQHthEHvK8dYVjDBYJj2pZgiJcWo20R7m
pvz+tKhTw0g8KwQS94yj1AXyAWNy9HJo00+3HISDZnGTnxnKEIKik8XxFvWDmMxqvJ1j9oYkmdcv
307i+NyjcVG6FbdCwxxjEFnKV94f02xjQN4MkS3iwQAHF3qGD4bqzr8gI5INv7jpCcmoR8DNRaxm
+9iA4BUeSGFYJ/7/KDXW0tK4p4+D6IKee9BKy8U+g948zjn3pJYik97IAQRbWszV2VTf5LkvtX7K
sjUxe3gBvCK2B7VHszskuR4ApEACQk3b+w4zfbtG9k7AapOWqI2rv5fmhOBk2HK/C2BeM9gBfy0H
7sIdvy8wssHWQJ+yxXCj5IHuqB0jhN+xFkP8St43XmkXBgrgBCRQ3CYD9zGTw6bPPFp064EcU1Kg
eB3sBf7kuUmaeCpu5JAfs10jXVMlJVlE9/Wr+qVNK/UEApNLJwm1r2WMTMJFS/FwaUZGyM+0OtZK
HJvYYBhOce1qv+wqg6idgzS+8v29KzBKAcK5bV5vMiY9tJLwFCd1JeivFpq01nzV+a/dgZ2Yu/x3
sAk8Cvo+q7EiNZfCYz09RtMMIkUDRlkwsxyWkL1Vx8ZcwjCGYAPL7xYKuJ6F/sK7WcLRVFOLxKOj
vVrAhGw7zYM38nzNMF4bPbKRXa4NbTH5CTLx+P8t4vorwvjKKKjbF0gd8kJolHET4hC6CErr/1de
xZC69AFvHfC2ZhLnd+UdBZjIjWaxVP+DG3yw/lPz7454sA6jsQhOmSlgEpfqmM19+SADx74HRTPl
hMjQn4LGPkpYj8n3ekwNbp59iGQ4dct3Ex5xiate9oJom9P7SGSMHoZrBDrcFdU6OcAUueox7xb+
q/8hRgdflS81pL30/RKrHEdDeg/AaxHrriWklgORNjtfApYE+sOCbpyphK9rbMitV911Ggz45Ze5
V/I+XoqXhD0y6rzoz+opuFVjPns1JZ5FdTWo/HEnsyj7ILmd/oI05hjwY/PlXC7l42WBnIh7egDw
j6SLEvdVySaTdgz47lr+1sSyu0wbRsTJRcexSkWx6e12nhPt9yCv1HwFD8GPzaTRlW6vzR3bDdHO
0cqp9D+yua6MeVM8V7VWc1slZ/wpN/bQzpnbnNsTNcg8HrVc/IZHtHuM24RJl+51LVsfLNVcruqN
DH7bhf8u3H4vAMmiqwt1+wHvO6/9l0G7DmRsO+UIqGUHR0w72pNiiOh7oANMpUIGy9Vc68qhNZAM
Sc3b7ymJcnEHMgKXwubtZarh7ggiiDpnW9fGSbKxwngORcdzng8S4ovx0nN4pa8AFBkxOosj5yVX
iQ3VZr6euj2vXaytAggmxgPiG54TArGYrP0HATpiyMRB5BIgDDVXPuOY8IyNyHhwpuVPVOSKIJvl
21M5YWMrHtzihGuQ98AmonuqkfUqb3umzCsdCw/rPOh+NxzPvF1bP+UIQiSK8UTN280V6WNrZCyI
iALZhQr89Up6n/SfQldOvO2eArPEiaMyOHce7M9tv821tsNo4CO71QsJU4hKE7e0cfTLA0UML2jQ
WpF4yYAga722L9Om+qbMfHyRGdVA3pY7kF8eBySaaABkKoOt9P14xODGDW/XlDvXyBjfQfUPHlwj
DOAMPXV79RKGna5bZNSVUlFKQsMn/dO0nNpiMV384y+fjiF0AizCyr4tSyy1ByZIwr/YmRI/8zS/
3ywVCo7wC8sGnPWQIU8vwUg69EQCgY3l5r5TPk1AFiHCCd9obawQtYcNRvMHNmybaOF0evVy5AsU
4nJNSkSPEmCgFrEwJYM3E70UPJ/dGUWFQsDLvDFHJFrd2DCt7tSCRfAqXmYY8kefYiMKRdHOZUyM
fOOu4FYcjjm11SNhhJPEpTqW8w2jbUj5kBPcwbcB4XQnh1rj3Z9twEXy2mRBRfcoUMwQFGL7f7Nu
K/ErhqRGGyWnZLzZOypFFMYlm0KqdC+ieRoHfZWlbKLwEndcNuzQ2YcumVWO1zuJ1o2MM02LWt1C
98p4+08BHPj3xW7x2EuWNISMOqX6XFn2rrwVjvggdXexIY/flqaqK/sZrSv2UBysCDv4aQJWGYkJ
jBdKl5FX1HAbMeVM5HTlmIWUyo6eWXllUoD5hGGzBptH/GraUQIZH77t8cs9Derco5Le3dK48FQv
dbGhEm7YPTiNhq5H94wVBsIF8BqipieZDt7CdFWq+13pueYqbuT/dwr1CGWaAMreqfANH6WtflKK
hnLMEV7XMvKKYh6/D6hUBJhWvkKofahH6/oaUmDU5tUaxUDE2PN99hHhSlyhcuyMXNZVfPoPxb1P
k6R/ggGESmyynRYs88BHvNLTsT0DGceVqSfQFqscwoh0xarJH/RasBarRQzII/qmLErJYvEXBSLF
9lO25Ipq/NhQMu5GJC/JXCZFC16eJcvK1/rXFYsf5oqNxj7Zx5IJe49IfZ9oz5hxBAPE/jWavIP7
o4GIcPbW5iaKbejp1aD5RbTd5EnwGk5LJeK90lbeAMmCSo6YUJkP9nN3CT33PV+YqmKyeybGJVz6
FxBAOfsxpL8XzhyWucgpFDQomYDi21V+EJHjBnQ1n6lwGOxVmSbAFAh7SDejQwgd7kAAI5EUDOkR
ip63wsaEmZ4gHeZp490Mj/Etq3a4Ei33qpIIJZEN5eSS7N6i+q9huURoOUEGl/NKGa9rJEnduOW7
gdh8YpxBNITOfqdmLa4r6ZC76uBUD7RUmKC9VZPi5wwzbCjtccV54mLARAupiZFMh7wgkBC4ofR/
5R5+kJHnl1O4i4FEcT3o7aIeoEcTncnehmgM9U2ucmSSAd/ET3ZYXpKDJIGSco5iZWNNIUr2n9u9
xHdA6SLbkZyNBVb++FFkq4kMMDMgGdpieoWVsnP8Ic4pbr/W+kGBr7ZpjB5sOQ/ejmHRrEcmAmh2
tUAQgLomzYiKxyKGjJloT7TcyMrPWGaLMfZzqJycnC+0FqhvzaB5+Su3deRH0szX7H9VMgiGf0No
gu0/8qyQIwBkJjdkgixj03CZzikQoxN64OdRr9n4XWy1Vj0PrIJE5+MizfrHmLNLaPqPAxoT/SNQ
qEOO1fwVRBQsPfQEdXl+bj9J6JMFKZylLjr4Mx+L0RmPKbCG2t0lpb55MoQMRkqIfomEbedYwycP
0QM3YMmCl48MQDkL++uOc4NPlO/lWESNlyxlJibCdMESaONFq1iB5QWTVxmGG7sBW2lMoEvyYSX2
oL6dpW7vnWn02FAb3QChtKxLJSD09qsKsXhNMTQ85AdptYvuDsZZj8Q5OpX8rjTDkWqltFRbxaqx
DNoKX6migKUSuXIbaKlv7uP/sZH94aucA6FcBU/C9hTsBkJu3R+8iW1O/piMXpjMwY+IVXrrk/06
HpMLRHPy/a/CoS7QK/yp5KPmgs13mbKmlygw9yTXPCB22AXT5ZYBW+9xKpdLGPh8vzEly74jY4T3
SO6fjhre3Ahq3yjWWFEiy3AGiR2n/kKH6LArtstK00u6607SIRIcXLOcZ2cBT9nvGU6yIg3ox19e
6pxmEEdUcJtgLWBANZx+o66gTNJ2CG6cF3zNk8vPujg6AkZb7wxK9gZiMXxBJ8vhmBszyJMAaA+x
kVamQ0A8KsC3KSFFSm14UE6oDI7mI556uujvSoB9a9bZZu2kUZyRNmLTfkY7O0E7nSjtoEfOfEsR
Bktulp6hrn0TBE++VOHOJGlFspk3cohHJFN1lq3sBa7T0fJhp/TfwbTluMILAEJa7cpQDOlatjwr
bX7CjzHTk8h7QfwtffUmbpZbU05H0BOhcqQ/AHq+mALcPITNAcsOH4nc0rNtwyV6roWOMMDmjVBm
HObngfGK7QyfKSd/sbGgYEU8EBohcnAOoaLoIvVGVMLOSTH6PtoHtofkulsHuywT6Zzdk4wlawrN
P4i+sucVa7vrfH/FaHWXQIXcyUWh5OG8uXQ9A3dzY5t6FOqpqpCX2HB3BBoyF5nqRLZkhwsv4Hek
Oa3QII1Dqpk8DwgPxRa1WW7OIV4chNLZIt+mlIbSXWjuN5hs2rmuKQh3z1FP+WHhfXs4PL+JzdwC
4eLvvkNDw0VlFhuYd/UAr46bMQiSu1ObtJxOIJezwIPBDeqEp/RkGdzEQSOYVERjNEJ41EvBA8P7
TyhCPj/vfsZU1SX6n4A2fJebR0Z8XgHlXH8hO2gaBif+1/ikj3gkcMv5q123cB5eLKVY7EglEhEe
gXZXnzs0Vr5ZWzP1Het0FLb5L2sL/aLpJZWHJOdCdHlTRfaocgFx330tcYpZM3tphKT//sy9p7eG
GWCeRNxgMtJWcb/VZfBdBSvZ8GhGO7vxDYLKNYd1/vE6mCnAHmsefU6iWtolcexUMzht1Q0P/2Bn
iAbL7E5KzCIOcGCV10SFgTGyfP/WCMyI3Q7ch5MWz99inIyq8ZlmBWLgxclHDGxhqCY5lvLCHzEG
Foh8GnYBtu7B3+MVgur0U46TqCRfqP5UJre9qXGm+B51RVWIVz3Gk1V55Y1kNxM+jElFLTjAW1tG
tZf2FdsCY6TMtKlBhulUHc4J9S1MMfezOuQ82mGh8AbdSu7Up4OTpXFRi2uYivYybsSzLuZeS0Gp
WppdglV1M1kjQYvNByPsaTECw5awBhWziF7OJYDuwDLKSTMmCThCvtTFU6gzKH19occQWo/p0xS9
3LZ7qIswbSQPw6SdmSx84UnXBM6MGvz4fk4aQpjc7UFJxYlr/9C727R4IAAgqt2ElqA6sEcqa948
mm3Kuu8f/JZlhg8KmrlhRAg1eQxrkH2TO7SsG5PPZylTkkmUdLRTWiQ/vmSZ85vY6E94SvPLgxXQ
QghdJSP2bWdLjDGije049r63i+079Gpeo3NMfJVJz7T1DWvbTdzyodriqfk5M++uwvdKR1W3q3kZ
LZela7lKXFktuIzPNla5z4HnZsETmpuPLOVORgQduPnfA33TCyXnaeAhhY9kosybMKikMEVQWX8B
J1Ums0ZlTfIzIsK97qtMrofS8Pp/YyUuzxC3gBEoG86Kbu716iF/fJmQVLetSXkO5ztHMFbRruN8
SYgd7slAqEWioh6jwvB6RaV2+dNY4zkxvrt5D1rVXhSEs43ed+POD6Y+AODkV2CDw7s/whdpi1To
UnYtI4UlTDdEA4NExbxAXdfPVkaZBSfvT6FlBK3ckDBRhW1TIfh4nPw7cY5TnCbOJAXaHg6YVtRb
4JiG4iXHSIx6q1AmWFadd8ptx3QmAtiqQOcLfEgm4nSofFj8PwslR7VoipPeSJEIApOBTuQeI2fO
A6Ke3pK9KnmpofWh/+26C3Y95OsNykdbUZv8zdgH2VianFv27TjHv4c+GnZiyR9Q3jZynGhljtDb
sby+MrH5bzjNAjNBDEUqNP5vx/2xFtSIj3V/HOOQex+FZKxsNb4FRVN4853M0GqY0BAuu+dZAGZY
GNzkMpO0094WRoAU8q5EO6qsH4NFWqBCXMy79wyoXibhibjmMOeN8ho5i1nj6CnMFKDoCoV3A5mc
2kTgA5CZCg49TLaYIKxYeSKyT+wAtNWn//Iydy65D5tw78OXjB3AY8dQ2UhrUn978eiNaM1Z/YJ8
IoV/qODSDVhs6eyfZa3DgTrJDDJ/FNpiL69z1JOkK23rfKznvkzFacJIF/w+Xjm0iFN9tkz07o4/
jHlQ467TX8d8L3ETj+9AAMGB1SN66QU04JifHDY6ybO3cwrlI9uNQSkXjjx6kwO587c1pHgUsQoA
4iVlqfi9YYfTEYAfn5kJNqSPmJ+vlcnLE8Oqu8aiKgxxCLfqGBeZvbY10XaOj53ScLjAbcX5tA4E
lUYcF2qYxahHNwM39HYKc4sAIBS2ixnB8R2xHgJgvurnw1cyTAeevy2Yyw+iZBHEDJss/MrTaM0c
53wGcSnYGOHatPDtZNNGFM3U4DvMLfdTbX0XW8tNBrPPm+sNtSDAuZv0DcQzzkVpstx43hSfCGZC
GLLpZFqlrTRL0LSJVzJ+/UrJD3Dlzu/8Qo5jD1vqS/i6yHct3jOIloHDpNE4zwM8C6tyoepQDDOL
EXtXV/pLH/JaTPjRduD8XipfPjYPO3m7To49nVUuDNU2vjjRVdLbwnayqZ5D5cdrjmDD2cosh8Q1
a5hY1vdmyublcTV9YzC+W14/JcU4zEyr2D1SCyaMh8A3ajAIorWAD2iusEPNO0Rpi1Ex7fBxYwY2
UMwWUDm9hYJozVWrJ4rRhdiWaOkJAbj2IXqzYFfBK9T7Zgn6ihPTs/oxWIebKFfw+f0lTZ0yCsXn
RuGV1BzVMLrDLpolBzIkiv9TGf/BLNZ3MXBinmYnXOPvJx7FM3t07mk+lklwZtDFttaqphmTn2r9
LPof4GWmOIk01/C/IZEI0UQ5TbjlAquqlvztxVQet47XDR2/YAgmL6kPTFvnUt8URG7cW8wEk25w
bl/1pJCyk1hgOs3KOO5TmQI20Y/sX5DWKgs8fSkNu1mDVtx2nbiPGRuo7LKl3aEI2M0ZJMBA64ho
hLhIhfoR5T9l+LJkKOaBaBaEqOeshNO2gdyYui/3Sfary6+RSFHsUj+SNy2lXzLwJc9kUwJtexR5
+dyBYt3CyVR0Tb+X61BBOAxNN+IvIfbNotTQtLvOsF8XnJ4DGTmmM/Vh6CxxtvcoQuI+LQJuyEjy
F7btKhlDXt8hf4WC1UCjwctoLoIFAcMrpGS+gGUL+ZgaYuAn/0rtGfzhpu5QFA6PUaGT5NSh64fY
ayg9hE2TGQOqtsJJuBQZ33MPTaKPuSkTPqc7z59KQQQ2s/4yQc9cnpxfa+f54opV8ZzThTbZTQQs
DS1WF4oJBCWN4FbOg4QE+BeGVYoUyCWbQDsg5mm/jgVw/3YAHPG48O9PCWLIuhqrHJ0yfUe83zdx
TmXomumM2cjUp9ct5Np90eUp2ePdIqIyD4yVajq40YNeoU4W4uTD9cC6LhWz3EAjdv/CJyJsVPCa
/sw/6rdnq4p/UlH2nsgU50rvVg0I2aQmoLOLP19dVRV3JmuIYSjVDeXa3nONFBkLf+T+p4gEwrCB
ZBs2VCxNN0CpR3u6l9PRGYOvDqpvZ1CHMblQOZFuSx5c9erxOk1g4fMaQjIVWbRn6aymbWBrxLC6
J/l28Rz+mQD4mzpIPT3lyhQhmwOSz8d6vzNf5KtfH9Mo4qH/8JnzB9uOqEYXcpSLrVaVjxMNf5W7
ivxdYTECp0xmPobfBpX7Hrsv2AumGXT5PfaZ7gzKxf/HZEc1b91ahzxiA/mulHdptGsRqVnb+Nsw
vvG0tWhBKQDKGkU+X2ztdCbefCeosDywxW4FftKk6Dutaz9CeeaqNwikyj7S7bcv85gvyp6lsNjx
e0JuaUfgwC8bgEcy9OAVVnkutUQ4HgjB7e7K6qvjyg79Rj22cnpTtE5bYK93fxRgWn3zeX45SGI3
9Z0h3dKDi3kc8dUdBT5X7cfldvH7YBVgvbuDgiIT81TtV8XsgSYP6ha9b68CARhe2ph0vrLZXYBs
FZkv6cH1IbAQqp8Z722/UGf5R3bat7sD9APqPYr/afGkBA21/QzhKDm/2b6dX8d7IPco8P3uW0iK
tUDQgw8nPq6GZvWDGn3S+x2YBtMmleKRPNgd8psjDHyfRyfPch8yXm3rZRDOhTM/ArIj9PrTem/2
OJKhL0ejEq6/tOYCqU87yPEgR4MvsEWBmvBD9Gi3/8MhVN00t7RW0GhAdJzAa1uJhUvvtimshkXt
TQmt6ISbrD7ZW9xMJJ0c4UQ67al+IxVQlcPwR/jYMIpXZNGZvWu1XRhEZZAYrhQAhyYpuUM09rcg
n3qF3B5m0Ly55LfRHoK6xR6h7NMAW78gCt+myTgH9z7fLRXMniG6ym4zdODbpYM7xK/UVi6YF9Pb
zycDPQb0aIRD2f3NAlKktkpoWE3xQoMoTwrFv8FbRmY/lPhzt84oOUBVHYyjhK+3pNvm6I4WhQF6
q8j4d7mP47xBm+sxmw+6b+2ySHC1txIBOMdS6tKDad/Qq2FMgCyWFOQd3cqIaYZvnMXEh38mTZw3
AXP3PG+jExJOobr2CnYyS2dWWHKkjb78HILc8hgOBkrQ6dZ3aD/lnOqcnmxs0Zwr7PiDOpKcP9to
UQJuqtNjpbvwFqGkHQ9mlkdutf2bvz7wgzGLPrbQ8N7d1A8ltdwtx3veR6Vt23zPHQKq9rJ5eVjG
4dAyszg1HiGRHKoNpOhZ6ohASrmm5gPK7KFZsAzLgMeP755n/i5x8VlG2GV/mu7tlboiLVgjWykE
FvAbIR14nssICoVcbTI1UnIrDPP1p0tBTXttBICtII1mTyNoPAR3nAY3wzie3M4WG8I+ZoLqGU66
+x/XXezF6m1AmGjTp2nBi3rghqflw6D0TzJR1ZP2zrOLr2vnwcbqJ+tFrdeFYBBRDllWTZun2nzP
7TnD2lDDnnzXagjeHrJmy7JnEyX7XbyhKCWMb/QhIzmxN5zHd20ZTLB9PaIr1nPS7mHWqVuRAXZ4
ShUKIkggw5LB6kbMCyuZlbY9TyQsiEF20GxNg11NSyuOOYzwZ+l/eEV1IGAZrmvUQiN3qgZmrafo
DM5szdFH/lZ10bO4WThX2DxhNdA4MIQqsB7N2XeUkC/9HvBdYQn0xfTixbQEpWRQvP9/43fGJNGo
DZUMmAdETR2QOtWe71GR0JZ+43G/R3r7U4qdYw4VWRcVhUcHebI2hOHL4lmtKwItlpeBgCfE9rcF
j2r8bFspAtjYjwVk2Z0t+jRi51jEOusJfdr8QVFqdE/jSnBjO3oUKGrFOBz5Frm5AZGd6b+AQigS
GamHB0zHgAe9JkO01qULt2Tt6LD5KyOXMmsgJI/epYOf4hkwKpQQ+y29IhGoJDHauTFyK0zyraoB
MYHzzcFABa91pI7GYaNVHzC0D8/pxj7y3fARRxx+ZfD6KzfthJ9RNhoddbUKH/C5ULGKuBLgkL4t
6gL44FN1bISWHWqdNNRfWLv3qdiQa+1nnZ1nXvD7lWz4gPp09pLNJasFXgjMXTlTFaM+o7BNjPiV
Gpa5LT94F57ezWPKy9iulfKtZJPMJY6pt3UXBO9/ngGYHD3b32BM5/KniygK0wYykAGgzwohgdeb
+9v9EtP6p9Xmw7tgNCpu1L0DzyIFVyC6GM/GllxIsaaY34W0PX0GIr4j5louMkp3gZzS/hYhMMc6
4Fqyv9xZohz3qt9C6fa3/2L5Gg9ZwYu8ol+GKtZaAsan9Uyg9vIMTVP4K9ZM2iDgpXMalcN3Uoi7
LCh92J8N1aBoJR1yQ4W/4iYmC0y7tZxW5VXvQ3Ypc8ZTt2fC1dPv8V4HhyYn1FtVx21Dq4Wd4Hso
M+3ZU1LfQjHhR+JgCmZvcxEZiabAxH5/WPuNkcCIomXCXJK1oK1UVwRJ+VyhT8WK6o/ndSM9GG+i
1dURv6WrqNMUYeSEm8KoHx2DmAWn8lOQC4nKteJg5TXWpHrcZ7ckHeNC5Qxe6jMdTE/sFgQDmk3Z
dBV1s+t/GatvTcXVXjTigrl4ftnpbsLjFSev/+u8ZQEN5uM0tz8G/E2A3wceLwA/sMLoZ9PY8qgu
EN0eNRLVZW4VtdvWlrMKsPwKBdb2yHjKUajuiC3I2fvfyeTf786UPGny5QIZTd+u3wohOzDHj+gi
29JeF59cmUj/rSb4KaeNpGcArQF3n/x0mpR0n3hpcVJLnDYRyr3sWrLYY6ndqG/x6DDxUL++8u/l
zYlm8QqulpDKMEXNEsG4azyPKefMxl4P5PhtVrEUxFEGUnVGPE/eYA9r6AWeQG7yjhUwdgOhNE+V
/1jCF7jhjn3+TVNce8IelApjt/sSW3UItcMyYf2R7I1PlgbEkQFCZpbGm3We+Q9s9pt19Xa1l69E
iurCGm/yl68kt1akeWRiDne8bzfZkjSZTUOBU0+1ixTry797KK5yX491OMrPpiWWhVFtGSrRsmGY
5EIcS5pIIkeMQ6+KVIHIIyj/4f0hCHYmaUaByIq8xlfaTCQbRVXNk9eZ3SX70ET7dufu1bN7ajG+
r4MsBXOh2RzGOA7z6s98zziHW5IOKmu//nSMqgzTqkO3ia9Wc47JmOwABzGOleJ0pW8+p01/WY60
KZFGDTgIsTdxcR3SifpcKzcxJdp5ZcstiebF1gsFLB1G0dNR7mCOJzGkyZjVLCDrxJWuzajZ+u50
UIwVhK5k3FqWN15kKhOQPdU3/1JVLPPblNhmDs7Si4GHWZ8PTqgW4rd8RF2rs9LVHRxiV4OXzvsF
cRM+uIRTxXyUe23ltbgq1afGgGr43xNHUQF0gE2lcUlpMeTijzNjrVTE8MGW6FOHu1fVV7EiFsso
3y1THajBAcSQ6eWDqmd4RBqjjgKBruu6C2lAjNNysnHIocsFDkBqcsbuvJ6g9wGwG4Nq7QSHUNHQ
MDjAsuJ1AUIJS+JfTyiWMdIqCFwdvDhHTYoV1b5Aa007KlNEX96KvyICylk/YZWj1OOHhpk++Dku
/I/fYL2rXPDepouGm+z4AyTMvRGrFu/NgV0PQnWzaNUFjnUpANeZ4CqNzbzODUHSO8bHdUevlTa1
EtEw5drebyjOW1N7t5vZla+BzB8wXRMkDAr79BUfzE1aTCgWVmP3h+3ca6+i2QB0mJTbzubMnwN0
5N7617YRu/UrU3ONyR6vJPzmTQF4YqCqwvlrTNbZihIPiE1Kmvz2RxjFPwi4eArNvkacVeabSN8I
zC7AJZnPpLab3s83tEfBrfPW4PZtOXf5zWFhnthr8hJz9jbJLdNg1+vx/gMEt4yTtCkqKYWiM8dD
26+0p11KiodBJbolxCMy12Tsct7GSRfTHCa+eOK11HQ79eu53U4vHJ5Tp6FlbhJUKY69UtSv/Fgz
F+2UWUBhqAAKG1jUPIjrTndqrdIZKvORXfU8GwVLlMOL+0Gi5p7+fdG170CQeolinH0mLk1rPMaD
TPG/6hNdMpPX0Tx9FMrkOqA1gtfLT5qfLFa4c/0ZRXl5P5eFd+UG5xm+O+W8uchoZkfTDB/pQxDq
PM1DaLFoJ/Sny2/x2qhbynuUIHowxfOEol9qHDNSGAs8ibMXYOUD3rel30yd8iGgSUsKE236Gkoy
N1bqjDpjYLu9Hhd43NR50t33HY1GM5+RVoLYMtm6vN2jqLJph4+KA6mLihourRLWLZEg1uI24Alb
vjamyf3+HyUVa/qQwfWEJfTF2RvvAdOt4fOgGh4Kex8Sm8N0Wgir0Sstt64UXnR8N/Olp64hCKTc
eJyTlfWIafJypRzvsgJVpbaQbPCxos7rSc/0RWbFxkQxW6WRrEpqaY1ZuQb9tBb7kZ6ObZzjeHCF
pBS6C/iY69FP6gjUGgyyobBRzQjAMpJltzH/pf8XexZm+emA1QDk4q9mzzTRvfgrFSsOAEA0tRuU
HbHGcyyJqzyVOcPQu33YRDj5+UFXpgZXpefSwa+RpU1C6n6+YVzh6A94u/N5NnjwGrkIZYVc0vym
KSNhlFH2vaBapNmebFfNRcv9fVBJudXDUQDsqUUl4y3C57NeXUrWmORz7+wgmLU8r7ERiP9kH1Br
AWQrPvQM9M6m4kwvQGk/PFvJr4YZOBoAFnoDSuyLKKgmBEkOXvyeH4XWpYPipyrd6Fpt4bCkIMcD
YrEw1xupYJonW/47EzH0HtKM5vsph0rW3V8Oxm2NvHELjxcjiVXtFOLftoioGmw89X3V7zPSicmA
kFSYcBuL26fm/pYp566FYBpi49/qxaiwym8PuRZTbdYr8+YdcJCKpfWlUGbEcOFbzO6OZqHDzrz+
Kl/K2KkKPz8wEtK8aaWnMBupn0YdC+dRNi958lBW/WzeS7T8F059UVPzgQbZ8GSv4vmVleZfxp8c
IQOYXXYFFVKLuTcTQDT3QwN2HwQGaGX2W+TfIzzCXTLnP23KxYJwAa+pcat5Y377TmG2TOqhujOr
X4YQvZmTJdJcs5xUWROQS+fxxJDEnuooD5H0Vv1aaoBGPv9H2sYCkeYbNfTxwZTyOwt0mOE1Rh/P
s1qhvbTm6UTH+BXkgbwKQxBvgRvQ7Y5B4hOPtxGgRQ1ocSmeZ35plZy1dO3Bmw1nYVcWedADm6fe
RRR+akgAAfB6cnD/DmRGdyRQhesls3DeYTe9jikUeYUWzkQgySK5EUGnXpG0R+5QuLSXKki0+7Ml
IZLkBr7zFSqCikjcbD34ac+NJ+RcYiPeP9EB6lmBK7/nigijgsDDFynwGfVGjsNd9T4F1lxr7QnL
aIqxXNyXRkBeRgZTjo02+tsI4WmSxfkkPaMd1JEKNT/vbBsX8fYoObEdBc/MueEYm9AMujF/TmZL
LG5lqGpny9J1cdXAUbQFsJUPi0Yd4cEffTDBb20aswXyBqpbNTUqYINoUbW9Dmnt0Y58y/Y6Hrn0
tdXo4MIsRU89mUn/RgscAcH2e2M8wqvknniKKanqePrTxwl81SiWofJXbjfNeDp1WPTDo/8qA6jd
xFiobYTVy12OIToJhTaG4FptzigJimUscdLCepfFTFI3aCWrJTVPTVwGfLhUkiJ3Eu/oDXXspQAR
Q48A+eMZS06awx6ipMWGciVDL2Vqh1eGf9PawZYHosrb88+B2OLAMtkUsJzRKPDqQT6rmi8TTdu6
LLQqt+nJe/phwr32Y3Sse0BYwKLqc8pTTAxHLW/z5hehsmMK2cnNA+y7kRaNF0PRSdynkk0I3CGp
A5TC2DnGn9Y4CVoetni6qrTTMF7Kkv6BBMCh65UKceXO7c454zARFYwM0pbAsZ0VyLDWbyk4VDEx
5+iVLejBnx+idiTim+7M0z+yg41Gs3aaMQ0XANggLcX2SoRbN1y2D7oriMUD4zkHQK4ps6kXMOqe
6bjA8OfCmRlqpQJLRjzxL17hs8gecWXqSX0/nDujJc2dEfBJ1r6lkAxRBXfA3bapvLp9KtlbOWQc
I7axeAlsTg/cj+f3dfiXgnznqxyyGYSAd/FHgc5fytbv6eA4KlHm4YUDuoCTBXCa8wQOrbPnNDK8
p6wI7YI34wjCNgoOK23WCyzkUX0xPX0NTZ9WNtWj0Pf3MT2ERpYesXr7cvjsTZWKvIw6LzcalP4i
tsAmm0rSj6O2leLGhezfxo53IE6I981Sjkt7U0ArUeNm9aN7jSuh+fXDO+7BF2eADOoGphU3wQK1
UjAYN3pHoAWTBqYO1VZK0cpKM3VYUpxmgBywkGAXYprGa4taXeyv4OAYqlPSRjhFKvgWIVoLBsw6
wPlQb2zX5YttnD9+IIrHSKXKW48Tut5vPZ0xuD2zX7oqynfouQTKHGWWFXYeL4D/iYvyMx2BSCxP
CEwLVEnZisSdPxplEQ6cM28tmA1k9KVGs4gfMXOmkE7jfua7YIDTeybXK2OIP1B6df6JooTbrezQ
zd38u5SOtEIw/qQ2kyCSOKRK9mcrThoKWzLSiF249ySMR87qDlGv7Zz1jigg+NCOow/KsGoPVEuS
bpVXw9EpoVqfjO9bNjdMujw9Jgjz9ej6lu7GZECua87JDhdR10VHtTqqrP6UAKcpuYiZaeR+LSoL
HWTwBIj8/xeLQhaC3XXjNxUtQwlwPcaR6RJco5HnJKgSRJcA4YlnC7mrkmn1hme3+WLrgPNOp9eY
I81na53KyQoEcM6qwtBwh5IRhJ4XbWuMyrdQR81j55cWBj8Bi8c2JP0bWBvaMo0RA/pDiS45rJYR
jzhfdpil0YjsnRnsV3kx53STS4j7Ku2ar/LyEZ+FEYHyT97W/ITtwveTgiE2NMaFvd2c/Xto+afF
FJg0a7CSa6bTFtU+AcR8PSbW+8tWGEtI2MnTsdb7/2dYLDDxYqgcn8eHgBnfXOel3mCVVy220Zx8
sn9cNI5QBsmn6Iv+U+9oDRdOgogS+NhF8i3vzx7Q5U0icG+LEhn9tpdD8dUbYlxgCJ1SLGaJV0GJ
aMVL8kmVLADpRsrVTColEsci8Ikes+cyAtd1ayW6UhtwfB1NUTjzQS/prM/y3BmmC0RbcuxezDgT
3DaDrrgfWvOfNi4TxKonqhonNIfIfBDdZ4r20AHDmy+yJRIQ9a2SnSOWqIHMcJXGMPEGzpre+sy+
AfESuS3u5SuBwzEtJZ4yG0BsYN95aKzitQXRqNI4cKWYmMoPrILPrGkc5SX+WeiQ8GGLhVTemvcK
39qp5hOh4sNgE0lCYYhakEynT9q6SG1+5QK/p39QlSiKj4RdD8Hqag8O1NDAR4ORuVzlwc6XcvaY
YEuxVIn5nB7t4O6KXZba7zGa9uIZi/EtuGcM/Z6aGoCDVvtB2oBby8ij2fcBpJfXNRsMXXm6y+F6
exPX2M0yl94WI9Foz71gMkTDisqrgyKBb3PrNe9eOK1ZVpUFWWzTRt3ExCPL2K0Vn7kpks2g0htn
zYMwBy5Yf5YLQbygX0M17Pz7Dub86vmFtyVpwGvVUZh82aTSkrnLDeRPrLdDKzfJjAmrVb5HiEok
XFtPIj1P9UQ/K0OmW98Kg0Rjz6hXGWj3T7SHdIm3SrXKUxN2p70oX+NrKTppNt2ByHc4m3NFdItY
vobeRoknF4KOpSbY2IjwFNCciK6fQPgQ3Y1SgpZ1wExgkHl5TkR3YYSwY7bj8dePZW4iMSkjzMKo
hTxyOXsCPrxwu/XAE6Pgm3N8pr9Xu5p0MP+Ycm/IHp3RHkZscE5M/wJjTgBXJX6YUI2YDG2CSe7j
AvI+XX3kW6dB+fofyFyeBiCOUHiP+ZqDYmuqqcrAylYuThDz/XIcgFe8jwI1D3bCRtFG4YSIZnFS
69l5VTPDg6455gwYT63uuWnBuaBtoZnOjhpi0P6XCnOzT58/+3jxOCex/bXkXZX5ByBVHAszfjxE
LugP3AYEsSg3iv28HReQU/YGZxrC5cUCdHIVJT3vyHnMQFjftM9TqLbji1Nvp9VUT1LfOt9QWSPj
U6qVS/C5aVGwGXgrt/TiZ8ATWFQJ+JCt6lsRWG0xbjL3di1O0KN2eW2JmeFQGDIYxH7iYwmsZiGt
8/VwlAgQgqKLF5AupR6rqpdX5NUSEb3gDqjZ8tWrhcoy1BHI0dBWSotDfRvvMt6h8x7N2HDvWHyw
vhTVD1aJ2g9cd0/bfvCvKi2TChyWTQbPZhdmsqKTCXa+jPV+Aq2+xrnA/IG1Ee2T6fueAY9JE4M3
n7oYrPRVBt9pXCGvlSsgD6VObsuI0efXmLB8ms/wQTh3g5qWQHKMagRofMl8I3P47osTtlu6S19p
TYrXA8aFFRHoB1swCVlNvPgTRVN2je/XwtCAkb9lo2f548AVLquEqJiwjAGh5IN+l22dKVutnjtu
z16UWq2xBIGn4INoPYnt/SwKXIX5fFkbV3pwHJBXT1Iy321gU83B5vFVg9IP1bHuov5PZ0bPxMFv
8niM9vC95fhiNOV5f07qF6xN+/xaUCGpX86zRGMLo01XUjVDZAYrOXzTXde9/5v4YbiampYxvRqT
spEfYLCAEd2IGMBgbKasrYg9sTw+TJR8iNtWZSVpvh6C568/yGkeuABvQ5TIgx8ZOzb0HyXoS7GN
vbfkPF2Vql9/9gluI6vDgFaq9cTC5A7ssOTRk+de6C9ImV6ZhgUs/4ydxK9hdXdxr2fF5MmH4vZw
bMhPvhdA2Z4d59stE3ZSvOpRugHjvBSPrTTS6TcGwPFsb0cenTfl6QpLQG6f5gXA3mSAjgsw22I8
1whmvtrKj+bMyoycYC8T8clWMzGJLhMI9y0hOyCG1zMvDQBIUFjlS7WneQ4Pdd/Ofer/7ng17347
eAHqqOde/6rvdATSAGFdedreiwYp2U19wwPJPmEig79Ws+WXo/vQoUKaAN65TFZ9KFMNP6M6V5ga
QX65tyWb5Y9pmYsF4nDh2fJ5svw2RIpxB9167M1pXiHNJg5gM9JM3LuAQ8+LpY8AI2n2Rw4iFa97
zq+pHugBBJPG/ODtZRn47si4rXiyEP0lOKQ1HBQ9I6qd0VDe3cazirtfz4uoGlu5xU8QQTwbTjcP
MG4mHYPdfsiLBZkZ+4wvKvUP+nChiZz4Q0Ijp69t5IjmH27cSC5JDa5uMO1Tg9HWe25bBhzNxWTq
0CVKxq6OEBME7OciChekj4GAA5a5FV3vX4CXQtrovCY21ELqEahIrANrRQOmkFycE2cC2nc4vpb9
UE6pNf2hwZoNOLTJHbCNkUgj2FDxEF5J36CSf1DgFgFbMPDWSdbd5Ta54eg49pCtaGMKluz4SZ2q
cSbVff/6OTLioXdR+/usfSvA0+x6LQwLkz2IL/+rXGJWCd3Tmx1bgogP4sHTTROIhvPsqu6Mcj9T
Lslu5yVXm9jSsyaN4SnNP3SqpD560HyCJhjNJ2x5AzpTdTfC7wb3LdUgL15JiQRKuYqFn8eifxnA
CkUWfJJ26sq+J/O2F3QBdNSDT/bbYzLb4/mqtNT7PEQmoVSHe8ApW4/bIWONAL1k25t0/PWmfK1z
ncoL9vdxz0l1srgNh9vLvOWdTlM/LBsn9wLzD/x1etRph3tGlaqej69bYjHRE9fo+9lDovZxOG0t
oiF9G+eCZyw7g/9HQa10xbdoPURCDjtsUlx+25fxtiHGqaRDRu35D1T41hW5hax7w9eaFAYPdp6v
MPjNbhKRtJCTLMACPpsPQwHQOAkG1vlh/6Nm+YtCORw1u9TONNpF6Fz42UTN+AMPjgqY2RmniLXV
FflwkF+/Bur/LGGNIL+1I4WLrVcxcUpCH4F5bq1RtpTKDuTVkssWlpPpY5/WMD/kyQtbMwppbhsb
GxtYLRwtWz1ySg640w5YFhJW8yrUKugWJIc2zSTrscJpkuhLFtZOnreuJaFP/2UXia8KNwMsYJ70
hBJnbkQ0nSAzhfMpVkNfD+R9MKvg0N1b/pOZqMSrF9BCFtof0x9XeD7q5RqQxbM04jVn4Nvy3TMG
KoYx7ikkQPcLO/eQ8DqFJ5KqWcmA7SE5FfXqM3tdTvLflwulIB5/52sBYMzcFjJIe53nhtXM7hI+
0Hxn+igGLyQHaXbM7zcitZYIm+dvi/XdOKdvDkOAjNgI3hZlGXmeXOCT09pIZAuBZWrzX34XMWjh
FhtKyBHzQUcJIVFXgZRFpKZDNa8BH8GZC/cXoIMwirxFRya4nF/Xe3yqgDpSjgr4vDsEODdluzNa
zSt03vegNhOsXOCzf9P1z3Qgu53c9S80rH49PpdpmKV4o39D34FYu2TsELHHSSmHp5RqaLeMhEfd
Oszi7SYvtprRkr4n0QjUgZJEOpwM/xFtEK73RUU+NOF36XJQlLqDEkCaDsR28TiQusElgUeuiqq6
sdoRHkw9+q1GI6cXb3s6W4/+wDL3EQEiDm9YHUWicN3e94KzLBTt1wksVvKZoBsK6mGxydDo6vts
Phy/pMb+gl2mLarEwQe1jFzAX81nbPqbD0f2IwCpteW7LCOivkIegoBbaU3G04t74g08x8+ZP4oP
1eEzjjo1QC1DAo3w8EtRfEDzkF+94K5B9ukszj7zJko6cztJv+hljO7QHJpaKjRGRjYa8HjpK833
ekn4YU68/wj/VNo3ayHQ5KCR793936yNeCPGQGefTzwoCd5WGsqzPtDYlG/iJxPA8r6Y3Prw7gGw
EA10dKPchzoIbmKyzBsuX2kO979Jpxo6qf/f2WA5RVtEx000AZ2wRAIUPdwpTn5rLruXfnZP1Zjg
vcWfVbNvbPnNKlBN38uzd1o2stY4/4VX8kOG1fv+iu89E1lZ8LZN7kcnd84uO+oX2oTwIZqsAHtg
wcfZg8L0vHfyc2DUTVSCnd/UMzaVvSgcQNDYQK4wxfjlIuhn7h1JCXhNKxLkCeg3ajqik8AUxyYa
7HRtTtxRuAx74I6am3E+rF4sCtRE8NsBylRIqWd7a+gWOLGhviWNMwuZ4uaEUduCE/7oMUMrwRlj
bQPiRB17kqhYOajw3/Mo543G4UyExmZxfA+0iiKgsUepMCID83Gwtq6B/gpaXakyuTuuT5AFcivG
anmTcR/XUO5j+e/ltNyTj+Dv4Wcf+UYVUWidvFEplEpGYGQOWzdw2nYOB08ENJSpC+2sqsm69sXu
25oJolCz4z5IEWqXDYytEvkrPcJWFh93ro8/7AO77fqB4QIBiThqPvjt2TSH6ro6gn88hVFsEp7I
jxpattoek7u/3kdWDxTPchY/SVeorXJiajufBVgs1IOKOQCKOC3VMfh0OVFd6hjBd9OuuUJANsQ0
50QBbLAhmXws254vgwkzggMmywVzZ3OGGFRNYveoxJuv3yB8mBmckJaBDfBOfSNnZTDxX4TwVC1D
mWL6ILMYGyjchzbsMynO6OV0YBF9LX8N+F1rIU+zncjhtHXeNpbkBJinEA0RmCiTgsUVEZk3Foh1
NtGQJA/Qb97765fIZKjwkW7TY8MSKfNSHWbWdKk9JbprEJCbEnFFFbg9CIPgajz099yVLEX5nnzw
NRh5o6krPlahzU8hzOtH9deFViCzBfVp0MDY59568D3Mi+gbMlqkbB1lI/GieQuJ6iZ08n9X7UJP
DtIvXoUx3ycGU/cIm6+gQ+8yMzIU1rhUECugqqXAjBpenIRcj6S6bDWpw5goM063EhGd0yhMhtSb
T/mOAMdXfHy7w5THLOP4Nj0GGWsAA7MmCypkcufdppLIv6e+0axVt/2725AcB8WjR70PEPygFYE/
7IPrR59sI416iNkTVDPVd1lQGG68UIBfYe8puoYP0hjkriVjmMWJU5r5q+ZGLapkVoH3sJ7UcsBX
g5yFXQbkESulkcZq5hhvQbnei47zn1ETUYVgRASPgd9HpNDZTI/Nepb87qiZ2ax/fg1aQfWOEsGv
U0VDxcirT2GwWWypkmV9uViQF25d3EVpyDV+meiraPyAkTAdGmJNLZr4JneEkCaxE/ntcrH577a8
iIcIzKfCDcQhdS8mOVOBmoyy8GjrIwmBHAHFOM4sm6SfBc1qD0YjFI7IjBU4FgT1J2Aqvg1GQqvn
QZkJBUuejUIl9HKRs5SUmGnaSpV0WVu5RFXLmkZSv3H6QYrjBZRiLShhlGi3KYpD3sFz6t5xP/8V
Wj/xV8MZl9QY8Qie+Lt3rKHbJT7GkRXIYHf/hnFh51wSx8HCG5pXc+aHB7vw35aBhYVZ7+UmVxOz
05nhD6aZJVHd4UkU7Id8B+lsuYfxw5OKe7d4aK5fAintuvRzuk3rOhwvGTYXl49csC1V+3InTKwb
lz7DwzhLx3mi20aXRsdoPurl2LGcZIbwnUJD2FM1oHwyWg+7CZWbTOuJ7uD9b5a8rF907xVmvsFd
bA0unf9oSoi8ZJG2rPJeLg7rJ89Zp/2gsQGfjhR4cJDwt11PTNvJQyvP+qke3v7q+PK87Ux+4aNn
N9XUHJbz3xajwPlIsh144KVVlWrU2mOHX3XfV6QGODoxQ81JfdKIAltuyi/OJkaoF9p92lOgtc6L
ftC+LlPwoK4gOohI0riUWQ41DZAoFTDHz68wXCTOlgH/pPALU4Djgk7tGP7KHaWvJSD3di8OOKHy
ubfW2J5U4rkccbkcDE86FTPlecZ/ih2L5ni1Z5pdXZQMpmwe2OxdsaCuw1qCzvpvoxEjflt1Et/Q
syhfZWxX8uAUSAfj1VkMjMYRTnScFl65rcIAvdpjAqd3SMb41Mp2lrAcDONVzlEWhQ100MrWtUDC
EpFfBOnGGEJFK9Kf98c0RYLTESSgmnx0qULxaX0XJOttvUwCrE+ocmYA9Bl6m81IUbSyknFMp+ze
dmH8Pjp5EZ9sHCC3ClzS3P+QxDAOQLhzOvwX7OQnSrG4yCVKXJCwRjNlXwwci+76ftyumXhQWWEk
ECXeEjKfnsLnV0T5RPZfYP1/T+V1YFB/cf3NKRpshKGZNzn86WT1fRXX7suaMtf7+HmtAecDw3nH
9zRj4Q2tGMNr2E7zoE4epwAXOar6cRxHwl5D/tvOKGDNDyui+TQU2nZZiMsG0naEZcfaQnJwxSHz
CZo3YOEdm/OTRkF2zh12epSlnzKcWUU3lKt9HWKGcqyrba4n6+eKbPkP5cjrrgKgmLsZ1IMmKyqP
k7k/aqPhQ31E4aR7YYvAem6zfY/avsLo2k7e/B+R9GXcntrbhlT8E7bXnMgwFWwj/R0JDASxFxr7
CdOauIoEXvZkkjUv6GDNMz3SFArt9RBVshnBLyDCHxOQ+dUYcLjSRqTQzxrOdjC2giBg7GAOALuK
6Aq5qFPr403u7UpOkfpgL+I5sq+3zgV9YCr7D0vyGLEsC0+xcVqlJOgQ1j5PxlP+Z8+RJHHvNsB3
7cNBe30qs1Hq8jkJJMEcMgaGb7YIYHhaCO2YkW74LtzXS4oxr2wzQUqYsmxVw54g4SjGl+uiWiAb
4hA3Bp38HBF0wEYRK9kZCMOg3YCX45L/7rgzZ+RwzqzutsTqFA8c5UOcVPAm5jFSScMYNRoAUqJF
2Z+PKWaGATn0PHZdKtlcEwx0cs5Igj6TZ7Hz1tzpdfM1IdyVK4U7iX98o5J115M11++hVcXT6lMB
lkKmJB9hDOCSTY++y9pce+mp2GzGr2ta7Cw4Kz80y7delXw+wTIbSWRe3Z3ikKa/zXPbIUc/3JDr
e/9+8tDtOXwK2fvpPSIoECqCMeV6YKm2qk84Ou5YzIUmjTnIyv1XEl8aqmvDQfy6TabQmV4ZgFvc
BZl/898kcKfey9XLjeWb+VnqQ58dvXtzOWwEJs4aobA00MoRJXKtja3eK5jRfvc1AHDgmdfDXFjb
c5Ip+esStpcihhLjM13Khd/adOg8sSi6yHKuYPJPfaEzb5k5e1aCieyLrGXszz8E2kbj7Yvlk1jx
/GSmzjX1WYKGYB0fFDof/L0zRFC4qPbuRuGaFdw5mxf1poJ6y/Y4phKOajjzND167WVAIkfiQLP5
qtQpRdtM++1aWaY1ZM/K+oS5dzO5Vi06EAjf45SBvknINkkTPtxTu3uiBRTKuZeCa+U1Y+AjRFK8
MhjXek1rxbEcgAVj/BLUTgXtlJiPLF3+KqkGgb2qf1mpL0Ds7s7HXG73vOJmarn+R43xn9BK2dXy
LtjN4+iZWR9hbu5AUmdc97zQv51LPAozUyADx/+pqY/GhFEI/eEqv8FysJ8obFADxD0LAQgGgs5e
2xdB7ERwOmrZwLegzupyIHNyxvQFzr1zMyCTxRsYXVDF24iHhM8cKbvWpDUssYaoqICigqceZcjw
+XVAOCM7SyGpNxxNa0cbuMy/318T6+qMzXnUiknMtmzj7KB8DTb27VJWo/2xc47HB45A/0Pm7kAo
fn5oome6HM3Wc7yPaDVwM0qsmF0hhXbllNtClt3EZHcbrLIp15FdgfEljBj46SiEqOmyeaENyF0k
70yHtrOOwJtE5xhsUmCfn/DrBXOrlzNw7EH9Mh5ZxOOpd2+qRNnb6+VTJvbTkC7mDYAKgbAtmMWx
LrAvnnmwPJGyRdZHGr7Sz8ruGadPknS4ROHckUht1lhVHM/U0MPykUJCHBsHlcv9FJjbYgnfsTiY
NrvlmEv2SAvRLGH7UTUSl3/mm0O/WjHeFnKz+/aW4WqS7ugr673//cgY83RejEWlU/xOe59INUio
D52xrDTBklFSO1d5aD1jko4ln8JQYYa1xzuuSNYzbIbupskIa+GVWaEnFLzmif/TwK+EBR5P35Vz
fnejr0YyDoj3GAlUjrCdIwQ6vW516wrf2APe3MTm9tjBrsZ+YDyvJmYxcwz/2JC+SNeFzbY/esis
q9JlMpdmeBJVi6pRYWdsTHHIbZrQDKZ0wkOsDt+zzOimL9md03JZc4H9wW2P45IMW+zg1rtxjMVM
RQlxr7iYVwXuIRxrAvZVen/vmKsm0VYex3PfPsybm/ASpScU03y6R6957dgrFkj9QLBqqWPBdgJH
JyVbgCmNQfMYC0Bon8nZEdCRqQ3ynQ4LljnaDKFXvy34MNcKugn0UWM/V9uSOZtAnwcMKNS9C5dU
Ub59huSwRK4uTu0l1kjzq9rjjzFrSwPK3LE3wWP1OzlDHtT2MrYlvrqvqnv2PibwwSHMq9padoMS
/uNhvhpaNf02zboZYDOk2a5mLP816xJXWFjP6Zd2tlx0ZzMQ+fSJVhefThWV691oIWdGuLnzLa8a
hwRYRkiHM5u/ihTGFHGW6x9slGR6qN3DUc2TzJ/yWCf3U07Djadr66O3zGwJQd1ToPQxc46H15Bk
rlYdehgyBNiiMuwS/dg9+/jIq3g+WJEpb+zkAF/EBJxucKAK8IMu/gtBbYM5eIPk7pxFWUaL6irM
TQaUS57kKtZhPuWue1+P4sX3PBt7ekL1SLd1jbAb7pLLa5RIehovVMqxWG9kinSZV7s1wtVxY7LN
HlwSXQjd1zb625zs3fpvBMAgZ1jxVnRt3Kr01gviv26v70jcnW3X9QT77aPM9RyG5aXflFkTIPEg
If6CD5mNCLG2ZB6nROZqlzpJPyT3qfw2tk0SALomkfWyqDudVZ7A8mSNFz0DimfUKwjPuiceaqQG
Z5qK6VHerEscJ3/X/NbBHNCmxRsZwNwULi7EA9whSttqtzI1VSFCJOGgJLa1LLNukkHdj6nly8O/
/vxthLlcgryMbtph0jl5QvBHy8fHjLB1+A0BSeu6g8rY90JNCA6CvinPy650AHkxcbvmhSLTsIFC
WvBOIvCEltlMZBNyoMMhcc1WHG+EseyPOUGidH9KdqzNwYB0JhKrfuOVg+vwFNxlhqEtCB9wGMLQ
q+Pl1QJs9LOBBeKrg8et/FvHhp63Q+TedCbsV6/96MEnnyQyU7UcAJGfytEh7wgAQY77CA95GvZv
1v0TgTRaFykgTG+W8wklsbwfIcRkJUx9VK9/DIQYYXnMSdZB3V5JddgKTpvm06u0pTlATfrpp/v3
vvnvksjIjw66rPEp12xY98HXnWLM5MXk7OirO/oQ+jQnbA/hETakgr14+GhpL8CsNOdEf5LP2Uq0
bi4NzffI6slAIuvBlABGPlHSyxqsu1r1YqYu6LTij+m0ef26ubU795vb/pDK62Lazfdht5gs4Ok1
dtncflg3QF1jjbVmKa/oujg2WgPvYIP5vO3s7j84aIuUJyFF7WP0I9kHu8sljOFzmEWW5oB43lK7
KHFfT9gj6+9xjpP8jY6mESvujpQJwvCNO0wWW1BnYBlY2SeQjhEayGSBBT7+tkvWL3hUHnzdWfsr
nTye9UzupHbm2ZgAVBDk2RPq/kWITm6cjPyu72WIhfXq2awW+RRQVgADAzhypZUh57N+snqMPbNX
piYCNV0NyUQ29/xRaBPFigsUKQNphclFmDUHI7oxRjNATcrqwmeH902XDg/xBtfxLdB6DSF1/owU
wo9JVLGT1txF0h0//oMNcoiaAw/AvnaP1WdYh0d0gTfGj3X2sx5RH5monYRn7Xgjj6me0d2DW8Mk
BkskCT+z3FXqlnrQE4x3p1UcP7ofRPioX/WF7WIDQG7juNvFiXUT4pKKpiAZG7A33aN/zj9WimrV
pN1qNKl3R3uEF3Ld2/3amuawRCbpWwfMmbnI2L177xKCTFQ5PUbwQZ1KKm4JQp4JZBqQ4n3o+ygV
BzcuRL9Srxy+ZYtv1yFgeDlXTdiyboimHWndawu5Qv8DQ2wFEzUerDG2AuBijOMK0D1h0wdouBQE
X+U0rkRttSx1qpABUYwyjFqgH19Qft4zOdDsdG4Rh0mUDlIt84dX7cvgI1+U7oz8iHXUf0cXmDQy
ljQwFLVT5IBIgZMP2/PPRx4Y41pbx41P7zensDNt3SM3D0XXghVqDePz4bYC+p9mxmbtWOmiO2vf
NQsHNEpDSNNDWR45hhmDvsx+T6wkxVeWDKrK/KSNNnU1aF4eCQt1cTuWGDPtN3p4yFL2oqnxBp0s
UFk2NtzRG9Hq9OlRo1x5GL9GwhIvCWVTi8v6DiXsygu+vMHLYGXbomnttzPwxwJ5kfnryl9x2+Yu
WLYm/oFUOPqt8oj88ztJ
`pragma protect end_protected
