/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2944)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/4TZ0NRdFWNvvDSnGYmLQN8EcNyiLL9L/g2ljowHrRpBLPkFKsa2H4TN
ZSJYRKYyghl7NU/W2EkTkmw9iakNOzHLMhgM6RUepMtxMNjGZpBitdXNa4Ss1JDkvHWUdLumy9Jl
hG+Un+H3SgMAh9SBz6mQBm+Dc4Tcy33voKbFFnNf0yOT8RwWczMaMVL18VZM4HAFvsYAtsxVv/mE
rz+c8NYbwGdIcjgCEvBF0VPlC+MYw6BRFYZV8q2hWIEktVS1k0hy7H/ZLbF+cmsJddxdGMkvN7Xr
IQz4/W2BlfCyHaZcxdW3sjUEgy7M6RfIlu/b74OJUcvMJGQf5Xg1qmPuvkvFwiXmo0zu1R1V+N+L
2dyTGCBlNKPMXYo5qPlTglmHrwbiUWmeqoCrwQUPARh06zjXk38Q2iZ4mT8QZDKu4a7h9O65BBCh
3ykjS9oxAn6Xvc22DhOLYQrXSDgFZe9GqQwzaF02Ry86zNigzga/IwKRGXIQlNRuTem/YhgqG3/H
wqiNucIv06dCMFGF1nlnQXFDpLDkthnwuBioCp71PTfkblavApfT218NcraP5AYoh73SIK5dabbj
891mRdKipxdQMEBjtY1eAVRA8cvimVlUKBkpr5pnPuqQYWEz9kODhdZyB7JBZsw7hCLMZLHRQZ10
w3jmG3TdcwsSLdoYz3+U+NG7qpDEroY66IQqGhQVlxf8ibdPEvN0HPfwz8Why4mhwTbC0LHsl2uf
oKqPdU/rxEU/bDLSMBsaanq9l6pDbTr+PxVKElN9Xp6yWGxCmPbgSb7XpnFnSfav5oeXanLwejf6
VEg+WsO0LzBRfy8Elhn4MSx+Zz1iVXQzsecojU4yu1Cj0kRPE6JvHSEasuT8LAESCbSd+R5nhyYD
ADD1i/969MeVPM9q/kNiqKz2KMVU8rZ2ogH7RBjFnQjoYHt8U4iddyBttdVaJgSnBG70ycgKeZeb
bh65MdWjNc8ACdB6r+aP+fzkh26duyC4BVs6gomXKKuevqfQsdL0S1h+7L4alTTTK76qFkAIDfSi
gyH9qvaRfbzG45flpTd7ucrKMSTmGG3vewRkm1j6wn2W2eyuioKNw2hRstz9BXx5poeM+09/7P8J
K1iE4XaTlqPNd7Z3sOMn5ZRNl7d/e1OwaQxZmZY5QSKggVtcq1MxOfTwQzRjSvcpcbwrZEx41xzW
FKwCgXu0sQBWd9nS47q1CtxM0KYRJyUZ8YO8m+9jXyIy/2FkdUR0rqGu73mESP+Tj13P10rEch2l
W8Te+rUXXLw++XfZP6zbaIzFj5Q/MUmiFVY/t2bP1bYUswFlb/nITqFuo9PKhYhFQlpbxZ5p7CjF
q2zWKzCR3uARj1V3SMHq5YSIimqnw23N1vt9BAZDJ1rdJ1gmE1LE1Ui7FoBCJ1cHE/Ae8xooiT61
wuzXyJLDt8OwcjpSVXs6R/P6i9yrTzNq6cUWK2tDf50h5rLOu/mJDTXONNXwIqZnOQzFJ6vV4WfW
qluNE87Om9QKdzrT22iNrcdU9exwFypG1Vj9Ws8BVDWf0qSaKdKfezORlxrKYIi1bin12WVCDiUp
qiprNFDMcZ/GW3DVAKgZTC3fMWcDdnHUgAnJI6TLm0Z7VL2WrcoAhQeGiXdvcRxqhc9e3CABxWhb
tM5zWBf14tBWnEh3Y7eKIq6+pbzhIUb0K+M0aE3yr8x4WV2Gc8XA/b7IpoWqnVVn7lPAEM07g63W
u4t2sCVSm9F1dxx81fYn5DUFrKWSuisWPRzsVZ4NdzOOCe6f6h2s3zZQiuuk4CyS3bdKzjaSnbYd
BQFJ2mtpE8FkJM+24rjiMxft2DqyKQIHTdYegXtJeLOA3i3jhVqIVLg8Cz+iMMDTaVsUz4iTixuf
di57s6QHxhdL6fzSe3ESrntTq+RYQKqers0Hnz/f0Oog7z3+b12kk1v28fcjY5bEnL6Coe4yTv1O
TdthS33+3T3BdrW2avXOo9VT1NKzxK8tVlRsHjN7nCJpldY5muWjFYjxvXyl1LVOO1UuFSYIya56
2Yzn20W1RNv+mroPy1rCXM9AGlHMjE4K3FR9DDbU7rEAH2xAu5MDheJTpe16ub1HJDrPpRR+NU5m
BWzoXOwPv1nYsxSXDlpTQYVFyOI6smQapxJaid2j/7CbTVNCCLXdmtI+Y0H3V4JJrvZRGcjL5Nad
B8X5GVO90WLtftc335mwQolXAmm8MCo8M5lvg1m0DT/9NTs7Bevj4C7ougeahV3DaeE0j5EJySJ7
60iGHzGCqsxJ7fiY6K1IKtj5xA5QzMZSjxRfVextibU8K1YnEG+p3Jzs12ex3a23I4bFrbhdhcpD
Vp1AUkKa93Mtt8/KQX1axWtmb+ovH+K47ZWtZzNNzaIeeaYWXvuAly0zJV6u+4X1PL04EKtKLpXj
uIhxF2V6iiX4s7WdOHUJCZQSyIaX8mBn6LlAx1V9sikXbPBihNFN0wSOzsyepYMupP3bTRgDOB8n
ELRQmacx8i1osmTMm6ggNQAQ/IuH2GWd4r7iPjsMZ0wTGm9ZVGEvZO3oqLKVJnzPHQB5n4xh8bq6
fG7HFgg4LlpBAjAlPviSsP3oic13192pgC7CghBkF2s6wW46/5eUQW369aHuC4cq3j0/b6sHaXoX
5PLbb4w2gSMs76JKa0a+cgWxck99PVYk0N5aI7ykxPvlZKX443YVB/vlvivKvqTl3xTVDhbkU6O4
5xIBYomq22hWo1EyERwmr+wbvH5edTUX01a/fwTQtIE715E5x4dKKjJbwKG7bo+0JOQ5CY1OnK68
lymgr7dL7gEtBjC8vypuFph3Do85HG0JKXCayGiQvXj4iMdj1jdA7e8qHtDBKAre+RajczYmJtQ2
UD3hv3Lf7TzJJiifRADNC4UGhSIHIf63TToYz8qxLovobAHy28GTg3QzK1FuKY+w0+MQT7zkwF16
QAJmsTUFGd5Y+nn/20HUwosWJ5D3Ti4Txg2jBvw44Yy9hQVx2m2/Izcr4NSTMlvO79mpXMoskO3Y
tY5U87hPHEFqXHlZ2750BoeBdYv4i6yw39lG7/zNarN2uEuHK5AZgVMFY+UjIaysGHkT+4+l3F8t
+uXKywXMxezL7GRnUpOoqv5CmO/42fYbqoHzjMDOPQ5NYfAUyJcjD2GDz2oBbh3wbIIzDe6HX9oZ
1/KGAJSPzb2BN6KwlPkoh04i1H1jTY95oyzFuVjcgLEwBqpGx9dFHyiZWoZ9XRBwmomcTlwG7n94
0NWXW1iZeC1AqOtAbVf/SE6wn1w7anl8ChSwBXIVSGfceaKVrXyrVi0M6zQzcTeRvHgXVHpBftKy
WAiany8gJzP4AWB7agpspZ0CLcsUt1ct5rE95g8dzijFemvpKiNd+NN62vCcWfidq0gOu+DT60S8
8gO3dnv75giN/8mGKTvYKI6YtND9XXt3EZ1hWo4HU32slhn0z+Cy2KB8c3Ne0CFwec1aA6qRBSbq
EdtSsdKfzUjkf5vHkhvBJlxrZZ4shMBASs3gpeX63cTHZH6HfCdufz9Ozdpe4aFAEZ4EYbj5AvUj
DnBQXnB0SUvEIWCVY4i3tjaaHD4WwT5zFmmY3ZUUlKwU1Fa0ysRSHJVD7pKrojBlLfVUDaB0RprI
aMa2jO7GfRHGFlVrrj7hhSE3YsBRbybf8gwth9Uc2oEkohfdtAJZKQuMFrNHB79zrfFUOrNZ8N1A
QbxeaK1uf4RFS6myGOnxlXiBoFFEalu4sLSaB2jkskS/xS0uZXm0UskmBpnL6uMsMQbQd7qxVbzU
ju2Ispimxc4XCUJq4hH2FauYmdTF0upXJAuqOcKNGg7vd5ZRHFLN//uXt5Ji7PN15o+qS7f8JVLG
dw+7yVWyrbOYprx/QIN6rEPnxz90zU28FrZIh8irfCVzOc9cOg==
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
