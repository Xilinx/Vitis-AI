/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvl5PNnflJXE6BNaKWkimsNSbbVcFVZHq7rglo3f7B2Zv0jOwetugo8UoR
pS+OcAXulaMhuBN4FkBg2Pm1i1EW1b78MD9BennF1KQmPA6CKcubolI/nSTuayYlPNxPo0Pr8VPG
kIvbIYmF3eG6wxUOo42/CP9baYqNNpDeTtpvLPIgrbz7m/tlqw/JHujMnQ64sYXzrTPidyNT5ynl
NTMXOnZuFiyKcfPA+PWQTH26+XpFSzOD7l299N5cMGWh9Ca0hffjfACj+ubNgP3GZVWjCMeqWXbG
/pYU9B++E+tnTtxNnB6MOHDoEyMbU7jsH9ycz26Kvmf9Ug4o/7TUxqUfkcPO/XSZJIWxHU2w+8wX
lO7ra8k8E2so8ErHWAbCD+TB6n7R6aGQ5MVCEprsfmwv/XsufCJGrYo1zx1OqiK1QSfvU+xhBQyr
ewsfWeTCAx7L9qz6A2tTko725inIyBuaWGE3c2igLTWiT5j+FO01zBnkOHnxZVuoh+wy406YYZ8+
6E/XVVX/cATV50XtHr83In/7E81l7fgAXwvYcrq2nHzB3Jg97tY72XQjBbWwUrSAKTc0sAf5wKaw
Gv1wgCyJSph+BxSRiXFzg8s4rCI1OnIqY6EGQ8gYUkuvX68dB6vTzmKis4g16CwO5HAZe2KscC1l
U3Tj2X54RBI/sIM2VjFKsX7J64O0ZcvYOh7qG5rfVVf6d1xpBS+7/6E04ZXLpZ4Fci0/bhkI0Y5T
ABFENYFKuA6hOqBIs1xIgBrMqqCwSFvpCXov/MH4AHXrBHYr1YtvVkjBeDxOXR8ppYToblJFs8d/
r6QP9qvOv1cQDca+fqL8JzlDNXOW3AoK0OKHEluZ3DJWsFiuwHnn5BDTw//dC5relbkANN0M9CcR
DptN2jHxGJ3WbximbhziBFLDyyys9m9es2zgyhMn5T1MhmlU8suwNuf3rzUOadv2hpXi2/zAr0zb
TQlYNCfMX3j0h/igyR70nAgb1hQlzAJaEBL3mnDXGNj+XnIrCm7Kfzz1uubDX2CfP2fTy35Xn+ui
ZR2sryj+9rG7AKh3CblP4c+YiUzUYzstC+/b0Qk12JAViBtXyawNyy9xLXt9//jMZSclO4gE/4dk
C4LPrfbHADxSbE0Bx5YKSif82ukszDI+b0/ky7WsZTrnxC3/mm5SFPomQscnVwQV3PM8y9f9N10n
rmpSY5lDJfjFQmaPC5nRi7XmHy4eKduSDFcLF+gJoxN9uIFFaRx+usxF8rLsb4eMFGaZ2Ft8rd5c
hiw5VVX6E+QEjrOuO4pTvVXdMQZKH/0=
`pragma protect end_protected

// 
