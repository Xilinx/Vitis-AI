/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPS0XCbnF6yar4v3ZxvcskOGauKZ3/Kb5+RxzY4H6QsV5FrF/5NNZDi5y9
DwRt5dvE9S9IhggxQuE6kL0zEtTYlrik6cBB5nSGUDUCzY5uIb7jcebGy69V7phYQ9Lg3zYfaVKW
u5WVIdsyGCxVpOskK71W3xOZOrzqcUJ+m5a8/xh0pTgLXEZms1P8NL3kYzLpRjP5dnjgb2hlZfDD
ace2uJCoU6zTNtZbuSBkeZ/6he+KOvV6ZmGoYSUc22xUW+f9NsCpx///ra9BlpiAYbLIdruR0DgZ
hg6msOP33q8BTADqemCAnahGa/NEFEg01rc19AxeP+7QfR8ajXl74pkln2MZAPp9s3/S3pdrOJrE
PxeQvl0nGz6xAMtRZs7VUeQ1MA3N+/Ro52vtQJ0TCmPDk8KodbvWQNYk81rLtQOy7eSMWkCgzqjM
+xZhbCZyA1r3aaOfvPoI6YcrupF4F7Z3jdqpyQ+bZsvd2KbKEuqV2atJB3+ZeQX2F5pfP25p2hYL
NGfI59T5qZ4TNN0NgDfCdh9AKfzqD5N/aemCXf7QlJ7r8P9+k6pwNPauSNZsvrQhUWYIlCwYwEce
NkxIJkFmwE6TYtgje9UsWrKYk+qojsipSadKq7sSfva7fA0BnYOeG8zp7K2JPuoOocu8z/ESTW5Y
/lJUFqAi0edjB0GQOwXIU5jaFu3JsPrkuBXIttWkCjWMtY/brsL4Cw7Yj0OraCGZ+NLECGEvWV6K
30tY2EtFmJzP/UqND6CdaK1xTyKLn1NWdutEf0qAPwL4xnapnlsFzz093AdXW21x8X/hd0YCiCqy
PfSpgDWAPiNQZ/nObVnmZVxrzlWR2/KryqMhpGKCNi0YDkZVmgVG6ng+DiS/vBlao34K+nh7JVip
+14tTewK6rE1+IoCsZVip3Kr+ItYYla8y0e+tRhwysLdCabY+f1UH72LQjCoBUQceBWxHxGsqhHV
2t5yA9P2bNx1NG431mCv6PVD8o9qCjX38jGbXKASFTr4pJ+erGjgoZKd6hnAKmk66vuGjQScWna7
nlZsELL0RXiL6EALrmLP3ZwG2N8X9PyUzjVOC6nqvhsVcUZR+6CvIrrIRf2pYN6ziiBg0UIUSaJ3
l7kJ6C4Axl/4dvkRKr8wHT9yvD3nHCN8qOpClh1WPyQ67SKirjRek2o1Cju6UY7Nh/V61+dPSZgh
bx5+Gb7nEIfDtPri4en0n121fMpMRyywD1Fs7bBsk3dmph+B936jTIkR/JpNWlfllGTPmosXOz7K
JR46DeIoCcD6jnxvbKAZSIBSx07gU9iqnzNPSMAkeyVfrKFl578d7vwW4iwTQk0pKpxIQisgGL+B
xKXj+pnbKbn053GFu3UnFv2rO6fNmdDV1JN79Ua8+JGqnOjYVWGRyaN1n1Y0E3e8JChf0ZVv/enn
/59qkIzoULcbId1GYO/4r3QJdNvZ2UvzZBZy86K6L3c9LdjzmW13WQ+6ZChmyACk/D9spDbYISpA
OR9JWWWxdwCmiFO57UQVt9iZCfNrOGGppABPa4sq6RT9qtzuFQ28e3W1JJlI8h7P5wUrqTxkPKCM
2pxhF6nmjxxcfx0PPkIJDxQ4PGuEd3nmatygVEAecyXueMiq1LqKXNaSkGOLxDpzTQhx83I+vFi8
QFubJAej3qjJRixD/KTXCqhkmkePIMDvT3iNRWsRMe1wy7IXxcJ8Yl3nqjlR84UATql4ujaz4PJX
2wAxTM10yMPQv5gF1rD4iJy7n5aSaEfcfbFTXwkPjEWadxhT6fqcxty9u21lOhIYLynbBQJ7p75V
6BXCOKkVhlIQQYml8FJWYdxFryWfKeK8GpYkfNHFxQhxOKpprkAN3Z3j3qqqeuG0Aqu0267D85Y2
Mb7VLhSjNBqzCjFms43dt7JFLjRNhoH1fCyp+9tIa5E+U2tdXWjl/GszWRM3elxldcuSoaVDgC1l
+Ppeqe7/OdLCSkYuXma/Lo9o1RiMo0W026CZrMbZDLi354jhv4mWa8OS7HbNG1ZW8u1ZIXjNVaYt
o6FIQcJOVDrjgprPI3oUllEOA5SlkafzURid1WULiIBvcxkAuvHzjvpLyC5CK2B4AwYXgdjnfPV/
6BF0wXLK7IzIFhSGxYVffgb4vD2Z+wEcHisNGZkFpd1u9NYFg01/z6ILqMkZR+WVopa+lVENCkw1
MY0ShI4iVRXtCVDH8DVu5b9/ZLlmMKt8aa+TjMpM6fN9I+z/dSwMpQysZF/BmszMNIlNMKDkGJdH
jkcFmxv/fZYkelau+GhVUTcZhEfrcE3IA6HlLFRx8UN4lEJT3GKfNZiXTyXBpDQhwL8C5EgYqvsN
K1rr38HHhhXEU4Vhh/wtZkxEnHtjVVl+y62+8837QJNoq3fAR6qFskmsw8dh1EGqn4N72QJTqWyl
MPSomuHCpzlhYq1Ok2iW6FsVbhq9k55WhRyHOBhhxdgW9wAXNnd6JWIwBZciyaLOdhW8tMFtFidl
HVH5HxrVlfg5xxA9RNeaQt1sp98AwTeIn4X5tFoaTWV5FxZigmeJvV4tFRsN0ipRMSEdQAbnxphc
h8OlsGlfgwkb3wIRmyvCZJxL5fr6gmjVBM0XS9tsI1Bmt51BHtXLRySFC89NmrqZrH/6CFizxWWf
GZNdLmqGHDNSaLT0E9CS6yfCRhor1vLAx1Z/iIYv5UQG/6jujJ/dOn0HSA8JIGppWIHWhKu47Pyf
loHiUN00ABOLL4rYmSL2l8s8Ef1b/NORHb/FQCRxiF5wae18X90IeYrO+Fg9/YPqCIutgireStEH
Okt0pC9Jg3Bge5lTene2/6oeuIIw9hLCwH9yZUeQZdm6PjbYSqNaIcGECYxvmE2vfj5HAWGinuii
K8cXLCTU/XnxXPUW7lIGTpz0knnSKnvYLXEVH2+O1BWIb47jXLhY8B4Vtk1YdAOInRZg7JcScsZ8
iys5xbFBthDx763HYaTUc+SEfAaTMvLHYwg2HTra4qHoelQmZlt4JQEe/AYRQTbYNH5DbNlsAKpz
8e9BB1g4GPz+yZLjJ/rimsYZC5hHRSXaN656vcNBX1iVTQS3sDalZ/Cdb2LoSTlMdsngw7RDJ8lJ
jrWNkL7xnWt3bL5Yl0FW
`pragma protect end_protected

// 
