`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35184)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54vV/P
ofulVpU/WhvY+xpgCU52RqLPKYMfFff9yUOEehtUiUhZGSzUVF6noO4URe2dI+njg0tFPKiJ2vLJ
tctEjtiodOf6cgyop09ObjjA0aM9NUjzQL+Dn8gCzeJtZ68VYAcDVcpsX/dN/P3Um/1noo8Iv7Cp
hL6sMcUXcYeKnjqPEDc8fN2pSfQOG6ND9vMhT4dEXBqb4cjt0ATINzUMt9aOF926W7d1nc1pujWZ
qv2NBDqykabluc+K/4/d51PL5cULFp7MCKxvLpjFPvnwjeIEO42NeYn2HJ/6h4pMp3+h5q6qgejA
sSaFkeuzDNzR+D8G0bUmzqYEEUUMvKSQZ557vczMp+3moHsyC1P9jACHopI5QmXHwlyZGPwBJXmb
LS7VAi59GhPMPv5k5p9gcTCD5TtLRJSibT6muX6sx3FuKE4oijTQ/HFMWtwSZ8X1fZAP4JBI7IBi
uS9rUu1gJNI7djH64asqh+3nSsP3wW9ttxuAyCjjWuCh5QrD7ZZaYmoryCOS/IOurE8pyHkqmhvb
tSRkChMlQwugMVd/xuFIZrFpsXg2mkY7+bgsvxD/ljrG9cPG0qKf1E+ioCIM+kwqSyK2zAVs1yUU
bRPwA+8TNHcbC0E9N2om0Rcxs2qOZW6x8p0v2Vb6UGC+kpdt3tFdKujD+la4QLC3erGFjAmX8y2V
rkwcO++LZ83nYMBve9K9uHc0+XPEQmzc4Cw5SYcrln72t7c+h3zs/RmbiPROA2XvNuDahW8OSIBd
FTGqaPtRkKaRGUjbRopRA63+sLTMErSBzM0lWXHYzlyvQvvQuia6J0uzgDRSaOETFtyTlwMVSoCS
LmeyCEQ6gwHsqNbRLDylRCahV21JzzYjf/q+THDPcV+22wiy3gUsEQ+clMTohcxBaPooDBTlVQnB
8tK4pUXmD7LD5beRanJBDx/fjrF9BRCOnj2CRVpGgezJal/pnnHBPK1jkDAIKG6cHTkTfR9dT4JX
lmrtJIIfvdp84JXeH4YmbCE80GdslsRe2YwlMy6BmwEtCemUag8cpC7IbJcueQDYKZ3sI3vJJtY5
F091DyXZHVs3jKJ8dU3nA3ZX5MOdSixEREvlarFy4qqIix8To//2Yrp93iOVwho8gjqFWAp+Ra9C
t7u9SLxFW/jJW+p+r8NMamafs2Xe52dm9njxy1Mga9OyAHBZHIO4vKCj+Q0d497V7Gj6ZWzk6c/D
oiUhpVCV/oMuueFoMXysMQz0HZCA3tY+TIYTkWcGEj9jzJjkZYYecQQZUWcKe1GwggW/tzP4EXFT
jskDqXH0FRwdZZw0KFeDADXb89i/5Q7QLFPs2CFIluCU5xw/EKmJXlebMKP3c/dIRv/8Ev4MwzGG
HuFXMpcNGgmjFk+uLd3UUwCdU4Xdw8XQm4SRu7RrLoFWK93CJYJNKij/2jKju73qQFblGUyx3Gcv
cgw8nM+B+DDtZXF+dOGOr5mEpfXs9heRZi1D5RgkTkF3XuPqo+8IL+/o8CpK7XzuBiboceKljsQ1
94PnARAC3aN3xdpg4S7lcBbouzQM8Ts6OxGKvZJ4LtBQzdGPTHB8E13Ic6mszcqsWcXC+s7vAf+G
Grn6kzwCwRJr9moZ5PZcMBX3UuwCmfg4gfebNDoLJSauHe3J33vchHssF61GBJOOjLp/pTbpE5cR
sHBOHP0hLUMmXNpty5xYgJ+/CJHGt2aQbwQhrHWznP+8iHbYFCXFWRYQ/2Hs0+jCZX7EBx1GjBuQ
aVhS2bLAvZ3ltwmUvsNfz7pEoQcBJg/OJV3+Gwhdr5jejknKu/RCDoBSVf5+7uU+MJOEJSzV31gT
RyYfdOSt2F07QyS6jgvSbWj3/I0J8gtIxFn/n4mEfb+udf3AR5kyR6jhMOhI/kmVHDqePNiQi4j7
cNVXlfQCRj+7w2KsPN8Loia0Ss1TOjzTvhsm8/JU3RZCTlCn+80D+T80fAOfl2tfZpis22/6Bmbj
R/8UjPDiZwhpoEg6oLRnjAPiOpxDMFYFHNYKEGub4wXmhnqa4ryfLTwHYaOy7gLOP1L+Wy8Q1qJu
fjPs01ta0iFWSykREHCMXzbcuzRGhNKqppm3RMT9mdElS49RKIzQkBkL/S7KdX6KZOHLFPtk1P0l
KUCnkji/scvew7eJrNv4k0d9JGLx0HWKcBa3lkUTbYxnPYjMbUzj7yvZ38PsVVDzP8qYaqpwycf2
khh63i4bxehoVxO/puy4Zvz1E4uDcDGj3bz06OaYDAZ6/23XT7Q7tEMUtKTaqqvQfMcg9e/CUcAs
qE4wrqN8JC+r6nvi+MDXHJ0Q7R2/04C6kd+8IK+cqlUGfiMPmNhJqOUO90N+nlhCblk3JxWhjmht
qXUvfOFE1xZfPQqpEToom2kfMnVNscEAGybsxaVk5mV9BvYtaDGlgrhb5N4wP1R2pwU/IFFGMOE6
9l+DZr+/Kr7nKITOEIYXF78QHPwu/rJiyZ+kpYr0EVux5s+cFRDYzCrUa7dSwN0ZNMbhSfujJNm/
y8JFQ4hn2Ruspup1sSrMShAGzABs4uCifT65iKasjSmDK7DNrN+peIeff6Av5Tm5r703Y60lyP5y
p8y04cXwIF03UgKsNuVQLV6ctVEbIwZPuvKAsKNdR0Rwa0k6yAhnrXwjPsZdNriAopzRUfz5/3XY
WIEnDWfx6kI/Yj9Au4YE/F/EfpDVLD2ivRTBJT1asIJFxudxJeXob28nRODulew23jlYpWSwWpOO
tABicDGcY2BeHCtV2wg5jWUxHmN5nxPzN12KOs/3iQFRdBuJoSCxDAt2CYQOhj5MWZgwHXXpPvHS
9nYs0f3cRRWpdW5wplh8pWslLncj2vi7weKcsveV8fgpRzBGMeo1uVYy/q4gMQ6uKNhvG/EyaPNP
tj9tjN6wRTVxl35V1iwOSGMZjYM5J1WR1Sco5aX8e5gTGd3DK0xx5ZOXxhMBeTPcHeVO7FT9Iii6
3XFg5hh/O/Cv+yDLAgD0aLccaGwySC0AJN23+feNiCAclzHVXNafMRbSWFlys1KW/D9lGy1Dvds8
N7QRiQBrMrK+rBxKsrxfgFyefyKJfoWss4JxOhd17oJZcGC6pyLFNJEIXR39mCIhUvxbCpmEBc4E
MB6i2HIv/9XQecprZ3WmUSr6+MR7lV05KL3V+JixCa07sfqdHlMkL4d02Xr7Hx4QYU8BQUMW5bjF
0u9hSIgzMu9JMtpq8MAsNcAZ4qfQ9eXKn1ybETAMkIM+nl2lTxdeJlsp1f620Qyb34oQVav8nPBC
9sny7oDObRV91a8wWZ4Y0rDsWlPRdI+mUjRwkTWLmcVNnyeEuWalXYqYoRQdexP49JJBTMzkxbvx
Hln6QLFFMUjg6TvzHdjlvf1n08SJignqi7V58mNOb3U9zTXEkK4sNdSZl56Rnra8b+1X00nQHWGr
QvsodNVaU2pYQol9vxhY3PrFllqYQNYaG5gDOIDbsPOfjUJCgebRimsQ/JGKF+kdzF7YcZpgVY/c
2TRPPXhOys38YYAlrCNokD9oxZrHmotCJPBqeT2gds917MLIbqO9KziCYk/NqhsOQ3q0JJS/aO9M
BVfnYE3XI1ngazY5fmxHVSAaY68hp6MEdlQXxSMW7JLGxUEr+UnCtZKQZLDooJGlehJAN7tgpzOM
3y7IHZys+ykz6WikxSYzBpbr238HKF0VSv/5ioGEcguyxT7VD4AxYpwuhJOWTQDMWL/EIaiH17Ap
k3f1ybZwAURxRQdgrtmzs1BVzbqo6u57sS6aicnnv8NDsABlCWk9vMSq0xLJxtNOdis+pp/sWiS9
GaAjq6qsaUsbYDS6xRIdkrXNC71dpg3Qx85sCm9Kf5xaRNWBb08AhRgPdQlt1UKyZxeS3/9bn2DK
Dx6FgXX235p7tCr5Qi1MkrgzFDpyPY6cUabbHvQ/onitb+3NSev1h65MglgFZoNBRtF7eSW1tSeU
TO7MFZRidiqiALxAa+jc4lX1bW2Mu/XsTBS5nQgaHWcwSnyfljx7T77xd4/pkRhL0YuZkytZCc9t
EowMZI7zwIjcnPnE82WkDHvDOR4v9HqW2t273Wh4m/hg2J9NYsLOgvxuBYUY9wpEz9t8Ux+D0Sx/
JaA3O/yDlAq6SsE90pAN7dLLomoj6Lbm+LdtNPn/SlEz/QWI+3hbuHhtu++8IiQpHXws6kzZ9Ode
HI/bC+SeQefogheFgeBoinnRJ7ZH9YB8YLW27HoNhmas1eHKIRoS8zSR1AUJOCOKepsBT+Ey/+gL
RWfRXRJ61/Uw1LY0h2HyVOcFN7VTOOv0XYaAB2q6i4MlxHmWOy5u7Vsv0WA5rve743xCe72pteKB
tsheI5f1nU3IqgMRe/Kk1kzrGS54R9m0K322wduY7mH586/gGF5I5gAGb6ehz5Le2/29gpG4rFz+
o49s7ucuccC31mIB4r0yeH76Do1jHnwmekHU8oyX3DKhTQksYDbzOvzWhpfFy4cyk1jQLWg25vBQ
EKcSTlpNFwQct9Wo5NRvRXYM4iiKyLVH3fBVxkcVli+cEYbWTI7xdPB6XHpAeqWx2ymab+rDtQZU
ZPfx8rfOSQUsQu5ratis0edzr1CrfjKg/2HVxeo4OThnnTsLlXeK39HEzKrktgzV4ig97RkVx92q
diCGPBBiVn5VA6cPSnIVvre7SvDs5hkKQlZ7wsdlKHCO81Tsnz0L8TK9MwjsutBUDxqYpyXtRO2p
YMI+shCe4q69L0Y2uXfrMxPpxkB+34CXctSnfIHn6cAsKF3lBZxhFWwRpnj1yFe/3k9mWPCwvTld
M6xqJrUXXhePrlEEusDjy6NskDoIVL0Gl0CVLeJ9XQy9w8pSM5bJMNz8JLi81srESZb346kkuNpc
+Un2Wk4MK1Qqwa/udfWppON0Q2qXB8FrF7VQxp38I/ku8sLVAUW4Qx7d8kH58t9fwRXamrMHUtnu
w9S3dmfRN7l6XJprTKRjgGqKGmfopHvJCuLEDdlT4JY36G2zgr2+a9fG6oQsBSOH3q8JxRX//jLf
WpJFX2BJKxcOErYWwQ8D6fQnzyU4iOhyfqVN2cQM/0100QctCD/t/3BXOX1hFPmNsVU1HlQzmr25
HuXS/9i4sZN+0KwfrYySVCrfUabsHwli7d/eW2wLT5rwjdpl2BLUk87zFphgTVvcJlwup4zmaCku
Afje+ZLEQ1xGSXJm8zwRnu+S7OBPflTD9b61RINhvBSsPpwN6pd8lmZZi99WOh6PDVs9P7Y57zk/
TAGq7AjxWjuAU3RtrKhvzTe3QvSzSCv+Viq2zEojEGp83YHRc1BobI1PmSzc144cJBCdf0zagNkt
2KESte0AmOOpDHxpIxKTlhWsxjsV76qYI4sQr6HtmM4qQHQVWTfwVNZdatq/BuRK3OLRAbRTY0BT
e5+kN3icinpqA2vaFNLOZp/5MgNmDbCGKB+xrvBYoNYfTukAGehEGfI9gnf9IYDgQQnoV8MUmHG/
hTn/cNsfSwJU4ph75qykWbcfuIJMgvbO8Pn1A5OjxVr6E8UnXMv/KupE5WHQcvfTlTd1VYdEhNKK
8m+esfh+GJkgxFObJTO/ugpkS25Oy3IcpE9FbVdPti24wJpnNpCVcDqHSJu9EVxrNZctc21NFmiy
3HaLF2U9EHacRJUKG40PP2LKysxlGmc5kmLWs9X7dQiXsINKzDOxvX+ybZt9LASEfo1G0K7oPGyw
bnf/QiJrvl7jsmuHrj1QUnBq5P8ouhqS7LNfWYHHpXWKso2t14Fz7DbcB9BVUhostOl/ipWjm0m9
43y/3fJYE9CcdP5vQR7SsMxCx+HJ2Op1/6mnVyFRB3So1Gt5t+8wL/8BdL1nF8/pSco/G/9UtYoW
SmhEWFGNPpg00GpGRLcHVs+GCZgziLXgoi1hN1geAg3aST7B0ybqRBxyU5hnQiUG7Vg+LA6fpWcQ
uH6PzAXuJa/SgodSSPXhH6Hn1xP/yTlOq1u1IN65kZiJK7v+1gMRcDYTy0c87kyfIH3ph0ko+AKr
+Fgcn3j+ka+8t8Obp9ZWBKNrhIKKy3Maz6NXeNFo+sxV43/YfA95JTL2jpyT3XGp1f5HGEBvIFpv
EJsPecNM7sOE4J8WnGBYs/B9Lmg7m5oiBxjg3V3gSwNnUC/zKJDthvMzda3HNorfnDPpIg/oVWCJ
lcyt9Rnrk540VIrIz3kubZ2HR+j+wnugXAKlJ9j0IREkphZXs01kxdnYtBMn8y0H9lVL7yBcQuOv
vVQRRXodR+DBl5FXKdsxVs2mIa2bxtE0qjn1hs9UTa0IaebWS4yS1VY9f+MsTrhcXYUX79TG3GuM
6PIF+v5e+ZmaqM+t+onQFAuoPcpcL246xleZ9HZzIn1c1CqYbighFdWgQjg7uqx4Ze4+CaFA6NWR
mfV7pB8fpggJ4VFILsEK3s1CpqJu8XZmx83ua9YOBuRWeNotzvGi0dLmy0eTNq3mmxU3uvs1hBsr
nASIvIa68VSgDdZ9JhCSRB1pi/OOPrQnJbzTKDLU1+g+dnkf+seuubqTwu8tSIjdqMaH5fLEkhej
fpDqyvrLhdpdi1oO1cbsiur1ee9j/0tMd7KlsmrrmZvobcn1XQXQ7u78of3Y1piWF7duOuIMnxoL
izqLQ9f6vRT36FZufl/EAgtSjdWs74r9xZ2hsi8tvyFSc6wDpDBIII48kwhd9aG6Tx7xmCYYSiv5
OVLLczgloMTLa8e3FxqeeWmuOedahNeF3f491Fw9HW0vv4LhSUBqUOdI2MKmhJ/8MaJZhzne/Q+M
3j6pUorJiVEU15zx2iPE90fDRfhkFCUQnsEgtzFQCjD3mEZYWGaXHxFSLX9/NPsY98aP7WM2+Mov
KhmYKSHZXkkklbvF3BQEaPfCwJnIV9b45fuaULX0XRqOjv+ENqE94LM2Rn/Cntzivi5Pkb7xOlnP
2F1/VX+n8YkQAQyD9+vMU1E4kVjxvmHje36lbIfkAvyns8DmD3FQP+PPuQiaOvsYAPmYXOdyM/6L
sILPQvBiEG2qgN2akG8CGjCm/89nrPzK4B5LcoHz6RAE8KLWVjxG8v80lHsrDJpU4Gh7n1EJiVfH
Ervs3M6aIq7C+5r7BqZwUnJPayGX+KAAyGNLa2mVD7IPjMs99jPMy8OjnZKXd3w1pW+l2hVQfd36
8Dr/MauRB+qWppANv7hcZ9AKxQ1nH5UuWs4Y0Bru+PSdgvqErWg58jeVogFjV3yOA6NSzk54KLpb
OxZRZZnq+vQUnpJVFmRpgRRxFJWx/m648VpqqiDHydord5p9oLxM99QbWHA33jbpk3ks3alAsJeY
v0v7219p0OB8EcJJ7Mo9Z+e+K4M5twnm61Vc4JZa5Xkzvnj2bW0l0McOJptlgZW3fBD0LvwcduZn
68kjtabqKhIRIqFK3+xQzpRfhuaDXZb3TrNJB1SS7eBZNG0L458RpEbHGFc//SAE5uQLfYCf0p7D
8s11zQ9T+C3UIaBEPhL2vzXuY1ZLxYjEet64EdfPf84YP5lI4QxtC52SNATW6Gd4yZz5uPlulrg+
QKJWsJoFJT4v27HzDsXD8N2cuT4hqn1+xfh8f6N298ZcDTCbIc8TEVIwZGGb4hLkl+gbH29ETM5h
YdV5n/BIEN4RlnGuhA/M/MzRUrvOvtYba1FlM9ltXGPlpPn27V4/Hfm5s3xKNeNRuXXbE1Dpavly
TQeA53Y6FqN0pENjZuOcZIJAuaj/O3RU94uvgMyhzC2gOp2UvBVgfPTubLqdklZAfaU7DWP/YI3d
tIn3bFcYWAdG85/WbLSIcx9t/SXGgEqDz+XwCesSvv7dxcaToeu4l80n3y9QRMaNP9QIJpS+dwcd
HE0TrNOEoUNiRMis6BYaVS/O0O0JEsR+QPme8KtGr/LDRpdWghhNI2fYFctnEqVjaZvcpXumRMSR
anEX7h5io7flmFNq2JaqSP+u33c9HIWiLjGU36AAf6hy/+M8dyKj+VueQI6OPKNisjpDup1M2gRM
XEKjPCxozhj7fMt+wPJAQ386mHp7CSUrwcejCWNcp9c3+9GaQQk3NP5Nzy0ZN679owxhYVVKSJs9
bP8N7b2rmN/OFFohxcWRCwxeG9WEHLwdM2B6iHoSMQTfURsQqvMV7j1Hh7hYm2DsNvTgRYLpS8mz
TzBT6ZrMRN7uSJai3cAlFhTDApURZ0tjparpSiFOOPk5mG7wvad4qRMVldqTF3AgU9TKkloDQ0pk
DWVYDI7TdBxrAYywco7PtbqStWJBy5vRH7HbQXehEpn1IsNvnua66d69K0SVWP8AoOWDf9Fu6dGa
BusNH1xtctV35nTvKi3/HW96MUCAAXQjv5TiCj/WXjFLHPC26prcA7zV13PmUTbs1bjyhB3Oo4SI
W7JXAdEuWKZQgGqI6Yod85nfXhd+z+8z/c9dUq1lTdCOQA27W0CRPXGUYSNWX2IJqCeU5OeDKvNM
m2P4GMkwhPDxGcCPNJNDF94uel401j/08K3Bi1OzqaR0rALoXp9e73/gpUVCG96406RzFIO3dL4U
3HspBM3ItU0cDAIvDRwJQ2sN0e7PDf6Ktsw9fp3OXgVwFCkNd0fHAnMpUsKJ8GcOifawimmavqPi
AenFFZsiw7ylvz1zDD6aczk49KY75U+qM0jNR3WbaNpvdkmL8I1jW+OhZxrK2JB5FQMHnvfZZMZY
opHw9fL6EecApoLe+fb1Sz9yuGLBUCySYFaMeO5xVASGCrMnqGByknAtgEn/R+hK8btyMgMyeEWW
07n1R9JVE/AzmOtp4ghKhkReYePItvS5PWCvlHfi/4/o2sRz3fVKJNGt6Bb9VFlrrmU/wfQb9+QH
oHDCsAY8tg8dBCw2EN4/+PfLws0Ta/vY100+q6tkERIJw7PQSc0D2IlPEF0O8BwPr99I2ggaQjGA
XA8hl6FrG4UfdqxKw6hb/XeIhkJNiAMZ5cI/iC4SVdOM6IYdpvwWCwd60GLWNgpTTXg99BPKyG4R
1xGD0eR6mI+USual5Vl9nW6M4FKJIdL96HeDOUwYmQkYvAo3zGGBRk3XiFOGsHDwBx+VnKdqTiH1
gDP/Cpsg8f7qmxYBPOlQvKbzaINIWxwv+EOf5KpnQtystu1h4AIkZ/ri2pq60mFhLTMa4lPiNfd6
J0xZFEmawt1hv4slP1xWs6gmR3Ir3Y7W+sb9ZZsK0A5k1F/bKw0V1DhJIKqjVUOo7zzzTARCgjYm
zJd4jXlsTJ8I5tcZFo9g7WUzVpSn5tthyJba9keEIR3cnAlRnIq564l3odttuftKe1VLTk8y9Io8
yS/0R6EeNNNI0tVKldfpH3jKXsHbmOZlg7gbRYoczbcbY6Ou9ccjjfBvqqr0AGjR5VyrQMJa0VPb
pprvaPLUTnVVhVDGPwROllzmDGToyE6hNza2h8TVChdhRZS8sOde4CdsPnDE/xtlfRQ80///9KgG
bYh37TSW33Ctg1zgf3z+Z7p+RPBWzpy6Wwu/2Jn0uSl7p/er5PB+nMuWFVvtMOFqe4Sb720XTRCV
32yOuVIRIfzpu/rWhXE1/Pw585GEFF8MTTUNsgUTocpfhdd5nGkBeC9lykc7UkropbZaZQCAHr3E
aQ91IDq/UUCmzYtZNt6yfJBUyZAD7j1rd0NDSxM0yLbmYUEDNPcNYI/UkU9hvJD/MnJCbowH+TfB
LioUEwVN0jW3JOitr3r98OjimFSE1HGD8J9sUIViix7ZdxjPeJ9mOoPe/vGbGWLwXpIXnafWsMU5
TtEXSafcKTxxcoLx7uhB2NM3hnij1NB5DR+YrhOvU0NsOr6gRTCvXAOLMWB8r07UGch41JJCQig+
D4t1/hFvNQj+9trmmdnhx6v+R7CFUGUeNW2JBQphkc9CI2HlbhhFnjdPUxSlH5w5wWiNgY35jKwV
8B+OMmwGgvnqfU/KDLnSlr1pkrqDhazycr8MJEo1kkwTz3eW5mTIXtGvx5yyElW0Su70f3R4psId
sLlzs3Z891IBwUY7tYNp8Vw0DpcS/RtINpcmYyDy3IaqoirtisNawIxAr+7O/kcQRSjxCNyiq2U1
fM0VEh2iWXLncz45GVabe4ZMqSqgJGdnMdPc8TodKiXy012UdQDsezlWtP3H7H8Zx+J3SdtaWvmY
FbyEUMoCH5Ub/iKBcl+RQwSlg2w+4BEV5Gga0rHjkfdk6Vx4jhFHnvFWkMTzkfmB8iORRl+6skbT
JBbudJggqmApCMc2MDs8GLB+1MGqgY1VnjkKeHaQicQ7pmS41A+Lzgm2rOmtneZRyb3WqHOqs3tx
odWE44xx7/rP0X8ucZ6YI5jps5DSUzgzCkkUhSnM2BHjVMzXSjRw5AWZoy5gUW77YaNRPbFqTgpL
To0CPqUrkZhYwDv5iXi/YxnzIKV9BAgC/KMzz1zvmOW60b8XCUI+fbA9Dn/c3qOwRmB1Q+FOqyia
dwi/AZxSlI8HxNyStK12VNXpJF+YSiIgakN4Wfw4Bv6jIi8zQTUA3KYIbNfmdN1JR1GRPk8QnlTR
0JaIpwyhk0nLGCBwADl4DP+3NVrky6UQeZf4XZDqCXe/52ivbWMPaIPWw8VsIwL4kftJaOLiFG9M
wrDHZJ4zTDdIMKCgOU07b7Qid293sU/NvAOJVlNRnMt5c8MazJzcNhxYYvgdajujHx0EYMl0o+M/
aCaHMS7xHlp7KJ/KnXvSyQScW6oHKY9SPU/Q23hkCmvm4SiEDfC5A44/mkOiIa42QH5ZzRcjEIbg
8VjDO1Gjwy5Js2OY9hyEofZi5oIT/H/Ay/LpqxeiogwqH3pzvi6jP8esYIcOqLvbF7RBaxQoxCYp
hk9XFbVgXx5ppCCy3Y5QkwawqJTJkGFdP1xHkDVbBtMtK9VR/2D6zUGKH8sL5oEEecKqywHTZpu0
9TJx/5D7B/xlEiVimGgQHg9SFh/pA1O9Nb+o9X2FNwV80/QbxHwq0CWbUu+tDVHdP/4NnmbUBxA3
BfLw/tIvIkED3+n8/GL3DNt845wZxrCE1I9JnelKInjIqZ0SI5DKjUmNOo4/d8i2qsqc67GxD+Qz
j7eucHgN5SSP66rair40dEk98LKkQm9JFAEBs4Mzj4r3w6/MvtlnTYgIy+sohSe0CK2EPSFAsjAR
eklZ1hG7FqEQ5c2veky3fXUiVEfwhOTS9Gx0d52Hk4kkLVePz7pPpXLmMt3vgkrO5ShO6WvJN47n
kJewC5SWBEFBwJNEJWmdRoTAmbR5YUEmNNCY00qnJs40tcNx90hTw4PDJ42EGOZPH+kM28vUPc8t
8+YgJgrPMtYYYxY5VgYQuXnCHr6sEG1lWczMvTHYvVL0fBnaMVTtpis/hX6SpDSSZYFwS20t43TY
CuJxvejwFwrk7oHV8m6vRDjkRawiYoF5jWX0YWFaK3c/mUZSQK/vEsi1UrUR/ryWrReVpoFCqsKW
6ZxNZfwcuxHkt4UPxxpkzZMGjTGYexuGo8TYWh6L4jCvYaJe9e0Odx0qatXKVtwYt0areO0G6Kj2
lkypr0DeLATdQX6uPq/ijpEFa1IVpA3obCvIOw7JJsRlzUlgofwgg9Oy+be4wxR95W4zz4XpsZnL
k5n0jNOM+fI2Nm4O1bqD+wyLQRIqVCHkBlRwEF6TcsXmqDethGJA4TCcSncVhqtzWcMeHxHgF30E
ndrbGRTozXVNhyfcaf4DN1FmzQgQVoidP2pUPNeKVzxPIl7XcRQKb9i7RjjRLw9HceXWhe2BTXQq
Ny+J4cgEPR0NxTNo7sXfKhOxjuOC3lErnvQMD6USsb4VEc7LGPu5kESZQIQa7RtA77t/nvP/3/N0
8Tykh8vlIuy2uD+I+EMUt5CTPJKTbaBzPdmQeOxSWGvCmEdR4HgrH0yInasulb3BmrN3FoG7kneB
Dl1MB9E28x1J9c1PHzEJKblGaYGm4Z0UwQyudvKVhJWB91lujauyYbwOv0p22pKwel47KaphyP5y
ObjDaKA7aFYgX5un+Wfb2SzkW8C7kUXKizDjTw3G+630gLNI+RG5OR/CQxFnNfrFT6cgJlQr7x1D
5Q7h31qRzIKzT26j5Gk7nVjRYpOee/GDWo6gQqPJDkwRi5hPDBu+eiLIp10+fdj2nBapoQwHnEi8
uviTmx0Jpcxj2z4tDVJlGy7KpH2xGQ1T4bZNqcJWru1xebenag5kJr9AfeQRaUwpg89jlWlVMUW3
UL/B58NU1XfjsSTbx1iQOxp0l9XIfg56tGG4E6XvYQQ+0stjBTSeJpcwd8RP2UDxAAYwy0+8ORpm
YJgD1Lg3TKlDLMZJV8J9kyce+uomkDIJJozVP4Fo9kDBWmRRVJhr0ikmToOxD745WU2AWCnY/L3U
H87sgsDgKlqsnNVIAmf4i6yySNg6QaGcl1H2Rfp5ZHlEGg2CeUQwCqaQuFOADnTl5r25LrGt5Nvy
Uzb7jIcVkM1sW5YGwx2mNRjzMZ8kZOyZoH1teZK58tysxEuj24nE6EscxdPradcNDWVskO0yj4MJ
wszJptOSqefz3ox1l+Vv/v1R4vhjotEMz+hkXeLMnTC2qFc/pAefAnjRIDDSJ6npg9y8Su2qeseC
IEfmQEiX+xyZUzcBQtJHlbXxT7j4M2NZUBKY8435XHUXY/d7yjc2/d8Nk2bQ2Q0GhsnPUfiubDLL
n48C4qsytj3nYDpI/08iFrs0d/IW5GsZP6j8XLkTus0UuSUNZsPxdcQ3Hj1jeXG3r8uqIR6MrIVS
svlOW19LDGv6OGSRE2pW5OPGAPHDBch+jc2G1qH9Mk9G04QXQ7NWjhey7uKnZgSUxMZKPksw9Hnv
gjmUyENLxjk+SbSUZTVkXKB4Jf5iRC/w6aAD8TlMahiP+FTjVvBaf5YBEoTI38VB+ISbutvjfU9r
Dgw3UwVxmSznDIo8U9aYCt8NEBwoFaVJ/2HEjcHIOOTxWz5PnYj7+4pay7OIWKwog7iudHEPrXsr
8HwbHyZx5b2KF2U/sUyJ3JniO+lZP6+S+AgTQ6USX97B4MV7NlvWnQ2ov2kMmYoTfsjn+oJIv3/F
CeOJU3du+4gG8ImcqOn+rIUyhyQrv/Zo1M2SBVEqvde2lp5eoJfXbAG5BEGGqRWepm9RgCg1YbLR
GA67W1LrV5gkcMGwShoZoK3M0BZfA71w76emmQSFf/+HBBVbcxdjBp7i8bowQXnaRwCl7XrzNqzY
ueYnCytKeh8Ku0obCk7frzeLk7ykTzSRN6u58d8cEWTbdwKwB+NWrpdyknt41D26vxiLVbYdP+to
q5tZAAM7rNLonOmUElVekgToT7c9t1RnFSw3/Wq9g5GXElQgtvxpoR0IXj6QvUP+xavm8vZes1XF
WH4rj8J23Ivz3POOY82jzyKAZ8OnlpryZxa9rXhuWjF7RI1Uq8brMgI9niVjrRVTlwou1PE4Sr9N
eqYSEY5HrEfCVkiBt616ZMYAPZRSxmJmihmhlSV29NUgojCOJTKM2fWE7EX2kAquH/FSFFtvG+E8
8860rAFauTD0lRrFLG4GDmKhyAtzQ/viFiErgYRzwsoU6TqfUrF978ab9u27JMm79lgIPWXhesQa
NUGdwZQR6jcJiMb3XOWPanPlndsWM0mWIIPVySp1Jsmzbq4hkghxdaeAE9OkZ2jGIJzP4xHshYJG
wTnN5/cvUS0BI4cwXTcc7a/E9uuGjHFoRhKQcZYDJPd5EqXTuwhH5CGl5TDtVJccD3D221ctHfiJ
dhbdsx9XXENg4zqJLBlhDnzJVKzYDD95/AaOk0mLjnAGsEloaQ51/3WwprHLMfvQkma/1F0VKj9D
Pe+jlHI1Et1DHqodT4fNHXuey8YwnJ38fDLkjObfuCgybnuKk19T0uLwLB8EkbjqdxFnckX5cXMk
Os849s3pyuBXZVMSyZI5u0ZBa49vKFoEWef+vYTWTYkFaCpSKwCia4xvdaKwGLIa/Cy3BqLAaose
2m+S03k/DI3Gn6Cz6lGI2aLGuGp7FoDKpC+I3F6Sxg7QJ9VXaQr5tOOGeTiEocjVXX2rjBKZvgz9
Odrr1qMxFqa2NVrRRWUlxNOB6ZNzCPXBwrIRf0yqtQ60OBpFN+kBTSnCduHKo1Rb2Cj83ao3g/qq
dFYECt32p70y0Lrs9w44mUF1AxP0mo5YF7vLlUsXbbXGGQql3X8iC9+/QiUK7toWS5yJNUQtdwV4
/RMwiJmEtelIaeCUUxqFNoVkQATC5qWFCfWF1z5fP8WQ+o81d/P1ovDATCsQv+9Ypet7WdWUWPdn
c9vDmKnZGrnFwhU0zgdTf/pyzw+uig08XIrIB4uAESB3xYiclIqYq38Rl+dkKpRi0bck/BZq2riQ
Dd+KM+JQnMp8bBw7RF/0gX9hHHZV7J1YW7QpxkwMBYHlv5fZa0Bu6uoLnMSdwA1FmKljY8Rzj+rt
GJgCWOjrAnrkeuwGVCoGqbV7dSqUSsrqbexj52pLSSDX9QQDjGev2U8ZlFnw1fivqnhrEpjog/kR
ofA87Y1yok5r9LPAo7lHrmSCzmxJHc6/+dcAwjXQrmRpSs2Oj/0+Z0+MNS3W59TCw15D3i1QEdFm
aRKUt0tVY01237pjwOdGUqt0BWI5Ys/rN7MYSkTlsAZR/tc3qOwJGxoj6dawhkO9RHqBr8tP2g8D
iOv8Gcet4FQhG6oEAzTwCVsCcYHcrCR9eRHnPkFwOrQlZICTZ2J6IIkw8tiea/ylc4aOlkH9m5Wm
Aayv+vb3PSxFqo1qCRHsrozeK2pnXVqTndDPgNACbQFGXBawjTJ5OnsZno4PdWMSBmfKCwGq4Soe
FEu/B4iAHA2mulYu2ziSI5HUaUE5qm3tv9ADSyrEh/5AMhOYZ6PwkukbqHGGuqedFcbqx2omb+E1
2WrctnRyZrc2NiJlphB+eby07BHGs54/q34lnthwPT5GFOAyv2+2qAtZ4oRLLAstxbI0b5EUVb4W
yrm8gE7qa/5p6nMq1IJDic0CGgIJuR6Czc2BiUr3trLIlRW/E6zpNmE4Ekd/q/WdgdPDOIa6lf6q
QPnJ3mOIXXNENe2Vu/T5sz+IcrCQuGpkQg73oPgrRAF0YW57aEkkRt8d//2ELxc8FNmbvZuQXNB/
ymvLyFshRFauSj7j8zGdSmQmbq/6F9RzX+oVkT5dvrN+SkgMKIr4bkjLVuxOlIihYdaT9ibyV7X9
3DmqrXvhE5snt7cUo35YPvuBDr9Zf8BYIoNvimXD6XHru7LLmg3DqOxvpzqqVwEKTnOMQd5saHPT
4jD5rNOu7OB/LSfXlXNRwkPNn3avd0V/19FoYjVF80pYFik90DAc+Fa6UJABnK49SfUhJ339n7Cm
Edy4cbeBcNj9ZPrx+dssjQqtmtXqwXiH4AD9gvD1uCJQX+coNmGaO4dEuCydMweSMUW62BZ8rNrS
E5YCbQsskcGrGCAETbEZw+rVhwrIKAotiGfhq3lfTpK+zYoI7+gfEDi3Cyg7vmzOXO1JE6VgHefZ
wVsviSKrZoWX53/tOwGg4s5YiL5FyKoq6JMpk1saJsc+2UA67l0nwM83aH4rH8vJ1uziTdSNfZWt
s/zwidhshaC7KdiYPg7BGl1c+q5K60QX3WnbQzb074N9JECWdJXOZCARg9P+scrd3UunYLt6dvm2
xGNbB2yH/XdSpQXpivv1BNq9L3esrjpZNeytSKu/4xkFzN2ZsaTGtKXnZ7xl868Y/0QRGLv3Kp8K
uxznYEOrMttS73/qXeUO4iX5Ig8cQze4xDDvfzbYmEm1fUlXYp2jmYG3nAlz9dInXMlE5N6OjSW3
p7VrVZ81VDQKUw1KT8T4XJ7kAVCJdOSbzSKfWUczZIKmQl1joWv79hnvlAFXnr8W4PpOj5rsbbam
wDRebMVJPcnhPLMRpzbikiTqKFzM+fd8gUxw9eaQHQmrqlNmkUNhNvlw+lEfAVcQP3eRBtKuQh86
16NWsExf8P7M205GrGOKfEdWZ377+AG2v2ykOqkf7LLViW4PHcHfjivxfgW/hgnBBkgg725vO89J
s3Hq5Fqjj67Wa9YUbYnvjF6l5KTx2qBgOFT5HYzigdEkT9v81iw9VQ0hB4rv+WSLrAYaTbae/SFd
709KCupP8+FsI2j16Zv56KweAhnTkimO+ADdppExCdwobPWYlTdSB4ySX48PNBiyVsOus+TK8pDK
QbM86Z2YVzkGNhoXd/5w6EuulSvS5/3bs5CPUi1g2NeaefSNmeGzopWF7QFuOmEVmr+u2pDprPIG
6nAK9lNnP98gblGxl1OqK5vo4wvAgA+0TAiwSJ5NckNWff5ntPNtTQTdx4ca3pBNpGzT7L09Ilyj
jdLl0Ye4mqxrHLUow+oqU5C3cSvkrZj46BuL9wgrvsw8TDUer5bXfAY4fXn/wIJ34Q/a2mcGu6ZM
DmdTuDAmPI7a1mQDs80XRYM7J4FZrlqKLhD4xVwTMyQ7R4p7gAy7ksD85Sr4lndP0RY4B6pZ4y3F
0e6DRfKWVjdNJjtdY8GiC5cCQi4oEFg552xnBlw49ukDDc09gq3PPk41D0VqnDfKGV8B6/y16FFr
9Tq8EjBjUvMsydD6Mm4XP9YVwAR9bS+JD5j3yLgfvQxne1YCi7U/nb5+n+hnHFmYAdmdtAgBMD15
v4OQpf8g+ApH09B5ZBN/PoWGtcNf5/ou2YSZo1lmLHWQm23HdbPUarXaEDhYAxXIAY+6knXZG7QB
Q9+M7S5pSPePgtDEZEA/QBZ7No+tyqKQYKai/DSNZb+64uxWORp2KTVSCfq8NIafPruCBsGHhugG
km1kKTLg5ln80dx45tQt1B0NKpmR/WfcAKrW8SkAPd+zuByz4QNKmK32M+BPWJFWy0nBaJVkuQog
hXtTuF0ra+AMzSEPK2pm1AD7qLj21vrUtvsspicOyB4Ydi7S0vVRlhxqc2PwKp1d1TWxIrOPDyKi
nas8ZYhggdKCbX1UJg8lsFGsKTfLZYOxA7NTuAPfNn9h0ho77RM0tUtlmqyrRQrI7UFNOeXBPPKA
TEW3B4I6j3H0VO9TSklKkIzozhWb7D7RzBcSoQHxzLmvDrtmVa+xrWX5yshkg39ZiwSOSTfrZDga
5ueyZqE0odVCqmxFYSp5i1bDAg/bHSY0mBlc3fN253P77GPJTOHwj0VsDo/Pl5vV09in7akaS7pi
xKR/+5S9qEiW1tX00ltCqjpWAvydi9wPBUQA3i5AeLzZqwzH77BEBWrCHY8X62L3ugb3tdTcCq59
WMCeTsMPSSqaQngVOXQ6N3qOh0+h+KszQaYVJ4dikspEMye0rLqmu9qGjTFKQBU029xlBQ63iR46
ePCWe+bjtBrtBPM0cVjpmxGlpYxWS9Ps8l8HW3deMvQkGcM6Tq32AeOjCWGEKIDQpU7TRwOt0HCr
u3hVvfc5eRYxLFBcHgNF5QoFgUyDfofCPmNLlpyNphrH9wGj4+8U1mpdlrkcTr4OJjLGYgw0hPQH
b8ks1JLWFQmu2jg8E05dFy40hw8h16k3kqN0I+/js61Q45Ub/88zGqttfGHtGXtxybtTl+wmtcHe
jzTbeaANnzDAr4R1PrAaJCVU+kXDOd+FuOZ198nCJd1rQ6Ui7OIkUxkxsvkaXz6AdAI4aB7fMxDP
Z+wigPH8CT+f+sn1SxiiPtCK/k5s8cn7H1tpIce5diVvLoc2yNTnCvaRRCGqbdNOuAO6T7x2yo+d
DA3KskB4niW+7x1pxCAkzfVBI+2nSRDu7l3cZ/TfITCgjonPL6yPd0xYBo2Z2vr6zTtydwwrweiL
t39OCaYFhIHfZILmdmEriaIDUy5TRENi/GTW5YxZI8tug85aO/rw+UIy1Mw9A4eNuDJq/I/CwNen
QgfCmzOuCTIc5INHB0pgCa0v7c9YZG/rPn7pXht7hkfBHyNXKKOyrjDfObpNf4e2EcsiTXNxw+LC
XL5XB+HxW4SrtzdoNThIDybAAtshwJt6qVLKy7YMfklMj4QuLmlHSojDsF4qg6R+QdYgkfpDhTkn
elEhNepbf37AxTGbGg1KG/lt7BflMnjsu2S74EOq9ZHxEvffK+5CfUO7Rb06Q4/SmL5KlWiANhfZ
73nFOZ3yIhqd4ckCzC8Cj1FH/aHS7rfXsQeKu1DOxIeqSh7HfQqId13KzQ4JOzOsyBGAHhSaD6j0
qAQ4RVQVGVt9Hojfy7XBhS1gurJ5XgXinnhWVYkUgF4cmsH+jMIzp75ItLxIUWYmiTUmbuFn+ayh
S1znt7uKnWR7jWs/BlkzVrWDsUpR6Q8XjUztmAq6WT/3XTZBhbfqG2xGgjP8L4U3OtA82o6ZIv6C
SAnte9aqKhq6X7XTA+VwEVa2a5cAwcZhytZvA1tOx2oBFx4l9SGT5bNv9bwpQ+NeT025X21pNwp0
LUcLppg0GBJ6/MAnjWXlbqi134kq3nKeck30KgZR3UKNfTKZtbSB/AntKfi2fzls5v6CPNa/iJYm
TNzEW7yCmGirEdlxDwJt7+XpnT93eU9LZvcxxDwsLr6rWTOb+y5fk3r7Kvz7w5OVs7/8n7cCMDDy
spTfSwyB7nMI07j9AD/dsmNNzaq7CU8Si5SpgPM/YsksFwRYL0xrikXkodA+9RYMVyZR5HWA59XI
I1XUpKLBvANBypqNE5TjtEuyFUIvHxBduFvwPH2mTRIaTeESGXxZT3o8drGVtuZM8VfcUWAJPRgD
WhgK0G8aVt0lpcB5ZSVhmFty1Wa5bkGA4wHd+5Ho/+NafPuIuN5ASHzyIlShw2cv/L8me4lG6emB
26rr/ChoyMDvF82o2EbXA0qndNbNqrOkSu8jWdS4+NQtQf8Jib9UHHWaTDdv3PLqDQL7T0O3ke2l
TlFLG+RvPLoQfAhMmvTa0kMFrTly17x7yoeFsv1JuAM7/soissvzIYhkTeY585rHKfcST/OwWVOk
3BtP8EH9MU4MXjZ7qDbkZILciJHkuLczAVhIHeuQE4qclSSykGGudm1TaNR326JaiSVSKkPU8sRd
657DdRl16O87LG7VHKgwXtz1f+K/XP7aufYwRuJJ+zgvHt4ApJwC4SRtLRm1A73Fq7hmEFvUMKNV
4cCTW4I0Sf1AoqZSsck54cfNFMhYbKz2q3SIlZUL6rg52q+1dzIu44xNrZ5SX6t4PNt/ChSAnOP1
SfhOAs7eDPNUKeWN4wCz0JfjxhznwShmKO8yYts3iJMc0NX6y5PoBImBd6zJgXsFMWcK9EM2rC+j
ZTBMOJATCmEhld1kkUbgyd8q6LbogekXhZSQx5HyBKd3YVtLG5lTJXoFjQ3ERW/IFtCguWFcXyYV
G1p5w/xqbaoCZZBKm+cZsRqwjpJz1/NIc0EcU/MX21tNSESWd7yqLd8F14ceex99H8N58Lyyr7UL
Ec9ogxmxV2Yk8OAWvpQPlLJQg8Anz560dRyjZusqstEUs/QaxteC6x647K8MoXZmNNy7ssTzxix0
QfQJNs10rlb0Wk7l1LcJIBnY8Df2JS3b+X7NkPcIf70YdgIgaQRnGrvI7MfR3AL4AKpAUsUmvTjz
L5Nj4ctJj8lRK/vrl09tjU8i97lpcDxUADIG3B/VlKDyl2aZO5/zL1Q+T+cjBehec3T3eWGiEZZ5
FPzxSIuTvoYhK8/IL7g8TQSSb1H1nbd4TDSqcp0c+1L6Nksdb59YfYZcNbgB5nJFQRgQoHxVD9E0
TE/ojQ1YEkEQZlbuXw0QMomwWrEM9BtJMfAfoe7ztCqEh7Utvx2PTNVS3OKUznJQaavctb9PksUt
kr94fD/ZFnEcEKem4GYH48o26XnjBvSQKoomZHUe2IzVV4FuEQl/A1VMiRlLagppbmE6OUem/P3J
8MoNICwSWAN/jMNkmOKbmZOAV/Zr3+RUzl5TkDJdwvQo/dO98n62m+9CBYRmsu9Haa8XuGot6AnL
5iWR1x2eJmZMX+29byx1iwUsDgDaN9oWdiQq6GgdRP+AMIMaP5k8Jn1oQWKGcixLEh2K4DXS/ddm
IHP6kcgNHc4Z5+5PUW54R+83M4zqVtdVi3c6SUn0wsQxvrxqVY6mKM0sviVnRsHZHJL4UvX8YDni
vvrIKiV+dx0jNfuYgTL3bHYIGJjSvbX9yp2hkVYIDCnCK6YzqCl3uEgqPos3H+1vC/L+imUP24zs
c3Wl01gsDGAHdNC/yLaPMrqIzFrvWLqxp0tObX6v1ThSyztffPCcw3g3hkzkz3q068AubfxmS4rU
iehNuQSDTChuvSO5TbPA+Lq0NhsqU4dfzYzazPHLwuMdzwnPrb/LjJ3op+bqkYHVpBOzReUhzQyC
JzB8pw7Wb3LkK1OnBcOPiRL4wT8C38k30Eqda5M/tMkUwogq3j3lozWVstbD6MULs4uep71jOnTU
dGPl1jz5a7xkCY5HvWbIAqnmyufD8kr8TVOwVpCqQeJ15IDHvTGUOxl0LDnnYgTWHd17joq6slI8
jemFbouawGeDzCYjxcplYr55I5LpqbU4zeDDCuJQ1eIUsd5fUkoQ2+Zkf4W8IyZlhzpyPEc00j0L
53HbN8qP36EsSsZuj4c26FPwsPTCpY64B62NsBTxc5anjXj75GLhU2gTw97VjhMoYfUxGMkzEhJQ
Od2PGf1fxJCuWqdEb0EoiuJGKhk8wWbtH5eSjZ7UOdAJEQaGJzb084QJvK1nvLmFNXUcp6NzoGZb
tCxXp6nRpAIiEFD0Z5hTgUjq40c584CU5ixvdzDwvJJesq6U8ZAhVkFp1LDUYfco+Px8lfH78TYN
1WwNadKvFrzShLVFc+IWIRYr/hqaN0iTN7lviYhx4x9vCloPtUWOjzcRZmtf1B++1qX/DXRMlC1Q
ErMH4GSZJDoUi25Y4Ar7sSMQs5+oXlOyF7eyi3mVT1CIfzehHr3iBGGydocaMJwoKmxK/49c1WS+
xcBiBwZ0AQ/GmMrOYigfzTZeeJsHbfQKQR6vzOWwbyOrpzbyFp9JRUHgO/KbjtI+l5XWRWi+U1Sh
TvOwd1kqFosm19PgWXDOOFQYPpXGzxfom/7ELlZTqNXMNEAzwIR8kazCMGiuYCjoY0Uv5cG2GAJf
nGayjRDp3pc2MqCBypAZ5SUbUaN79t59pSvQcIgyhCnJy2Z9KDabFPKwV9kCUTuHbb/ScVZt7XFE
I4ru+HJlEM23VZLNGpjY+jg24ZIYkpv41T1dLrvZd7Hn+JPIJUT2zXKzPlilpDi9ZKr1iSmAT3BP
RAHVYxwETuBM8iQkSDxrvL2qNy8QfePZli5lruQchMXJdC4q/lYEVFH8J/IxJgGTIAh2LL29zntS
3c4V+DCbt8HgtpaD4VGWtD2LKxNcVwVszZU9gQeb7pO2OQNw8gOFcgUMMN0ABpkKHZaflofd2whK
SQThH4gF9Hajic7SYmP32RQ1NQHYJQij+eni9XzqclWUd4+9Vjubd1vcZylHMWexmV0I0dAJF3qi
s1nHOd5V9IhOFm/F+zRBrgU8mptj+kKzyRq7b3C0p13LPpsssYqjjmaZPDrQH/80mdfAqLPM6lw0
sYAsrUV+x6epYZZ2a1f5I7yuvInI8LdcZpaqQBte0yJ27A1DGP4rfTuo/HCy8Baggh8KzbR8zYmK
RQp+SdvFsFgEofcM7McrwEs2sPL1VcEYct0hRmNr5lOoIBgZWvS+4Sp7hmfy/JMTt6ZLLvOa29qF
c3Z1R0rWKM9nLzEGQWvHPqfTBKAAFNRPqwh3Esn5oD/zvyVfa6OBsbSivKbLg9i2yaCvzLq133Yb
0NnbFODSPixQkTB/CEbyG8PcZ0eomkswajRylyP98mC+E8+QmWln3gz7cWKy/X3Eu8w9u7fpbF5E
GjOruIFY1llyuqpZIXZRwALATtSx1HSJsT0BLCGtnLTk2f8DYaLlBap05lGL7NhkQsj5OMK0nUlf
2nU0y3rBww2piZoGKykv9pmg9PaIWht2zJfTOPsZcyRWYygqeil5BOTPiZ6fZ+tdIEzzlHYV3ew6
+JvIm03MVKSkDQqBS6UCdgQpssg2e2Q0bX+cSO7twy7NYahY6hwOxYPcx0OOoV9714L9OjMiYr9I
eBz/j9o9+wHAu6Sh2ys3asXMaFwXQGM8JvEQH5XtaCV+8c0Wnz29TBgAsyWSGYO83r4WVcdH/DkE
9+CtvIrQhklzjD4u/fmj/irqLnsmE+JqVPIIJWWXBqKwI1V6SYMsz56k7qx8tk3Y8jqdPgXuL2s2
AAHDWeAIR1ISP80mDNFvVBgumYxx04Kg9L3KVkOSTs/DsTxQXg1D+hX33lwZDyvBozjRlw1Ie0po
DpXwmCNj8KVq5GlOyIi8W4OKyfCCXxgzdcWShIUr5W2w70hAQb0ULbr8+OSepQODE5HflV0ju3Mm
x/XGfOkOh/LmjAb9xhdIw4H6aYVCLlf1TyzXFATyd5Xgz9XtuFvtwrXCEKFhWCDw8r+xn5T6RW0u
v42u4fGE/jk9+fqTgkK9gZvCI5Dprs2jwwsXKxx5au5t6bc1uPIezGS+K9C7gx4PNUb9LG/H9vYw
VGgrGmk60uHO23M2qMGYC21OUXnIB+Pf+TZkZml6pVUwHbjen4k7FYoVbT06W+H+jNlPo1F9SQq1
WPuW4xkE67QT+TT1AZXolXC2eCfxfY+8bDTtInNK5jno7nCEyUXuLpAkAkH7nLaIB+2LdXzo6j4W
hSm54ACL8qY9Gj8ucR0ZUXFEWQjsRdaAWan/U26kMmKL5GdHGlDyt9jQXBKQKekc/beU0Zxnk3+S
gfNRi7OyrA34cJP65fdXdMmJB8OtH59tH2Y6/O4LcBynEgEh9Zj80o7CI013zz/4D/bzErCOBxqn
afNozymy1G5KNHK2hwaEcMkWHpO+AJ/qA7iiTAVpgnPJbiQKh896ErPS49sGJheplhninD01k2xl
KUIBZvcNiFV2zfJCnv2QQ/RMkzWUdRQTWrrD2j7y4nc260FObZZejcq3ho8EuB9LJPINCvRanhAw
m1SaO579uBg3EIkj+1TYMVieZT/EqDYntD79qY2YbaZkS2bY92AAomiBfqY0Nd4wSrIuqGMkZ30S
+oUVCu69okubQhakUhmIawSZDaBGG3o01ha9QztzOjlvw/225iJhkGUJ94yR/dN3prD31E3TI3bP
3JxGcWpPiMDYyOWXbFU8numGd9VC/49I2ibrmiavAscxXjt3qPWMxxPRTl25gXVeYjoSKlqZQrd+
XKSp1Mrpf5axKV68BOOMAjm/CCxb+xVf3HFyhksb0BpP2IbtBLzsRunEC+NPE0dYhUZvg9MtGKic
m8tlcUs4qeXBW6Ic/YpE6BeNzgXUVC9KQRk5hihk/wDuuCTRFsT768VrEEfygGJG+d1I6qwitcrb
v4eneq6ieJSDoYGRjAMXLK4pBZwqXB4Ir4feSCjV6cvIlBZ5Wq05wpQP3aiN6kL/MT1INs+/phGd
hwmw2II4EhH4ghyiJeJv0Y73R9Wjdo84BdtFJOGn85BL4cUMqSJitAgHMdWuJwOfa6blN5v9KaZu
EBLttn8jVgoIRYl6aBjDig/b67WfJb1cEgkh7mz8CXRr9bdaiyh0fZRNha3s0+aChCSsoRPoHS1O
KCjkwOG/SoV1CCG+Gz5g+qC5XLt5ORxUfi2Vz86Uv5sOm8dnMBdVCp7tqHN7wKHaPUJA3L2Bv3tv
BZEULCUlur5oXZrI8zOx0QFr6+3il4OoYF7ZQpE7RlxjPApAYaR8tm3F3dzf/C9XCQ+YPj8dw+Xs
6grhCBaAZtPmd3N4+aN9m91KCxRaskPKRYpFwf6fmUEzyZ1Sw/vC0XOniYy69SEEkkPd1+lWZOnC
d7WxGGX1Haku+CzO0B9JaLV111zP/yZ9vGTiEoxIanoeMSu1HZNS5t5SUWr52/Xd+Abbf0KFSmiY
sygVb7J0AcrZvhVkzr1nHZ1xMAahW7fVjUfKJUyRA0VV77nstC+BaupBXoKc6UFG00kPlPyKM341
24HgIOWWOytijLz/MnhoWLCVFcXP2jK3AMzb83k0NpwGHoO/Dk9fSwKf+g8w/6r8efCzxm5jU1F4
cIZ5ayXE6qqxYzScc1wQQdYQ8ULyImJwg1jKmDd+uyTWezaXaZkRA6+pAWZB9k45kTi3aPAKHO+G
PaH+IvLY0z270y38iefBYxr1yUKR9GzZYhGYfxoLoE2/wY12Dbkf9ysAaY2pZ8MqCJbT8QaMTCZ6
qCo7r/emmSCu2DuSPoMXmCnelQLJx6HXuTJ2hjaTTTsSx4RkhWgHDT/eGvXJSq5HIa8HvUfiIzaM
SQsmA7QjgXMXHKX1TXEYGICcm94ntL7rpvDedj7d/fUazVdJsG2pyQvZOAVnwoLIMKrADXWT90Hd
WeF/jXydpDM3UGXh9NCdOPMtuJcn8L69INPKzBl+gVX/vVhfXIKz2OdSMgE9BUJjIgQCde1O0Qqo
PhdTP1xL2griX9osdJZdHVwqKeLOYdzKPORMBfQloCzjczfubeg+LlYDdjVcE8Wv8DM/Dsekx9Zb
j4f44ISpcNQDh8rn82FhzHP54JsPtO9TZR0pWSmjsBZS5SirihheLIvqEfr56aueTbKBlvaEjN6l
A3zvM/g197zH7PQepG3kgMoTCGydaY0sy/vnWjU/rehXW4TlgWJ/qAgJ2KWOW8duSTIR31Hsv5im
s/z3M8GdVY5Hl/hfBKuxv/AS2xnezQT1RUJtZ8t4WE96CGEpDjrm+GVoyoXI0R6mOx2sTqKPFiew
ECYlCfE0Ij7o+++MHYQXyxwlXrEkje2z5mtsgoHtGNYPnEzNAiOp9ImM7r4zFDI/qnm/CfKAJi17
qGdkE58g5NhHCqFN4X8qnCniC75TVLaS9+9joZd4Aka2ZFiKIlGk4VuqbLwVHyml5NDmcPC1/prg
hbk3kJK+bebA/nHk3d6RPCAPn1UnSbpRkCBUAJsWyPXlPDTHm6F+9umOrihqXdxPk4eFN5e/7zsR
W8HTJqUXLMhNd2QlGJpRMMYYB3IlfoprpEtjp+b7+l/8vTjD8RAW+u8jexqO9s7Kh1hxjGn+/o2y
ia6i9R+R7zLtPqvi9gCQsHUA404Hx6NyjPFvaRUxXeyViPW0+lCdEd2IisJ4EH7kB8H+PkupraeX
CkzxU57lJ4VKpEDoU+mDEV1PUhHy8nik2NzpupdK22g0QMJ2OFxg0qARqQ+TpQpUKEdbQuKw42iI
eUpFykX7YKQrWHiH+R8HVyM1QqdsVSosRE9djmT98t9dg7Lh6vNuDis861zkSUhtZfVtDFEyGg0K
uPJzzPMp6AaKxxGT5unlsS/4d2VDUklJv9CURNFVIA84c2Lcc0d4EubUO83HtXh0RAMTYTPJVQeb
tBg41OgoaRtZ6tbQuyJ/25+MxP895KkXF6CgU+X1Vasl6svPMQhIT8T+PXcaCl8yAzn27QLqsTJo
seVCBz7XXJ6n/FWyBGKqHY5SK8uVBtrhY5n5hf/YRqXPmDQqbp35tiFj+8M9VmbYDdMrrJwGUeel
Xoxa7LfZXHu2zesXQA+8mC6X4LxhvmLGzYwrmm3uZM88PU1Vlt9TYcP56YLVbUTE+icWwViVcoL4
Nzey+A4btKpu+2KhahoAdpEtUlBO5zfaBSFG1oLoLhja6eqRLB24Ua25QbJGwbaY/n3pT3jON9Kj
54Lr8ilFremC15yyHGteqU2lOygL0WknV8BIXPCZbzqxWXtB0J6uzOhPSTzHEkD50OfEYmXBUlg6
vimfM1ZVkkhiSxy8fajvyqghbn0fZLrzRppjPR3ThcKexHtuwleX4DNgjXGSi88slCQZTtLgdix0
5v70W7lWlfWhqMnZRP+LsabcC+AsaC+HiGOxNuNGKllAzkHvVDQEn2lKa+HNuIuYVX54ZH1Yzh1L
KMOSV+LCPP/mecxVpYzP/qHmFj0KUhFP9W5aIaSOxJg3zc8Msx+5Cr5+1Tan/G2QN1F2ZKKCVvQt
0BDMBSkKukXHHJbvhfXh1kwuSwWNRK8rS8USDBMxDI3zf5kivm/N2/8ejNG+FPBXDunLDte6AFEU
+rZFoB8GvFU3qhsDWktBF8CiwzaXVHdEFOxMlkpVeqUH7YHjJXuIAX2vhxzt8bU+1uAVCjJ2FLOI
9f7B3BrziBHI0KWL6G4e+HQ413kmkRMmGeyttyXLC4GJ1C0qZ8stSkP2k9OeBfbjyZphwi/m7Ctn
ZgRbN6rLjmBM8jtLtQKye5SmxR56XnECOYn745hrbJ16HzZDIsjsTGLBm81tnINMWCgMMl7I9Q13
12UD8+7o2qlSQl7VmCot6FUpnzOI/IJUTRlc35uisdSYecGnCvZrWkt9qAxif43msRK5gGF6QX9N
GY+GXKe5NgZsFg8QXDUCiw+1bWSNl5NVirOAqXIcXxuUoDI//nF6cYBXddpsE4oETHSzB7UpXJ1o
Bti4kqaIhn2BxKeQGDUVTTG02W7viO8cv+0ohpmaVGNdrPx3cOIvpi6xkl8MwvkAoUf1FKBzSQ+Y
fFpqHnZhVuziaIHke3gMZpRPOZd/5vZiGTL9PEOj7wXVbKB1hOM8EAXRVmh3lDPaXbmPO3UpWCZc
b0+kL1/XK5J3LtHnJ3eytMrLdld0llMHxWJtqDNxHqW/yxMjldwcsy9sVvvbfaV66I6F9HsSERXR
Hrq1vyGOqbMScEMfN9wtZQVKWn+fea/9VSGRMZvg/MMYoAg3q7Ef7yT1P8+zDjDNhMjo+PnGSOOj
Eo2lZYLqtMeNI7F6seXKEd5OsxHjRIH3Ekwde3Ng7z7GgbN3HGK1bdcFDJ5IcG+akE3Di29BQqvx
tDhU4jRX2AWDhRA6AbXOG4nA4DouOZGwxmHNf22bxExMAwMvu2N7V91Drs81AxSgHSRUO/P+S1p7
JJ08+sJ8DwF1boCfbSGdOzt49HZUDQOMCgcG1OAstPSn5mt7qJaw+bXdfpjWX+/be8nkdTz+k0E5
JEnUxb8L4Kk2uhs42NAp6gB4XeYYNnz+WIXRvYGAf8ZiQDVvyAGYrHOHmrItf4sc++wk+LlwZB0n
0/QMoGI7fQ6cLsxGnKPzB8BAJi4lBATeUNR1n4de0roLPtvgZHB9vJT6eZyJCdKVb32AeRoyuabS
FtGOAQ2Pq/xRjpSCxy4/9XpdvcZVMivV1KFADvpwdw0t4NHVnhF4PmgXl4DiZMe/l4zAPTv2aDo/
aKyNq22desFkEtcFtJps8ekys0R9nduDUSYuBIHP//GaCVASu9hZeGwmSjcxxVW2PgHIXfoeqYWO
sykb2tMz9kNrVRlCUuvqVP4mbkXDNo9dKqg3Ds6j1yutYChYXRu9ZWHCJIbaL/nZBBH/36dspKT0
nAfegosv72HdjyAIXgP8BATJtgYioqenosxgLVReb1smUyIoYx5c/PZ83Ct7n/yEPo5ehuiFVfMI
DIc7eTibRhYW/qiTXOJM+j1/FFE3ZHNclmqHqw4ZfsONr4MNQHjuFhGThD86vBPM7STXFSGNkYFn
rYNtYMtAkRP6ovx7Yxrz2+xyfFzH7Pri8OVhNrv8L1PfifSLG97B20Bm103Kp2XGD1h8cUWmA/0N
/G6pxbTIZ3e2UqYqckOznaCD+ebUDiMc94juzRkppzZgabHfzKpVDFg1CLnI9UGHq51EaQpb8Mow
CQD+f1Ftf7DhDczPX5m0/eayZAUEOeqinLiU2aEjSSpz4cEHT//Mui6jtqrCS/wFLJGBK5d6aEzv
ZyLReeXcFis+txL/ANqNF/ExjmbhR0FKvrUD/xRgEOREcyHAdmGAw73SfpGYoy5IQeCV2PG1B64w
0hGcYufCG+MADvCgeggyt0+0GfgDA7BYNX2MHQiXFiNSjewJfiXC6HsZkUHOU0noe3TIhl8OqFf9
aYXBC+CSea7tlnhrousv7JHcUYqKlduPktKF/lX7dKRHZo7XgoRM4ub2BJ9FLC+8MTF0S+y+AOeb
jtR5tza7ngAj8oRFlHRujPXtShiP70+vthXjdONkyFGVlhjrb7jSP8CQ3atKyxNIOnDwNzhYmUgW
3+3R0jSc4PZyuTYc7Z49qGlfptt+mZ/dazY2ifGp3uaHHUVbaFFk4j9rJtVdPQDK2IyMWzwZ6gSk
tgHFKF8TEBRg/d4ELa227/efRBS2Sg80mjdA7ZMe+gIyKaquJ2HBLE6d4ID30RGa8M9pgGaZxuE9
4Gw78EPxSXviu6bsITbtLfPCVUnCoaERw2YgPXYuHbRBhEOEXtrqZQClh0gRPy358xkoLhb1pUBC
zmZ+G2nd4i7ViYbONh/QOS58me/dyKWo1OQAZYAdmEiFFYXIzHi/DWEdwbEju2VhoiVhr3QD1UFg
e34UgZi1k1OT/FMy7RIPpzrZi5Z24HfLT9IJKE2pY3yf7cxwZ8rFbHXkl8FxnBh0jozSCh73P0vc
CNIu0L4gKAzH3Zj7D56kBX7EmtBGPMWGOfgVl4UrfKM0OyVAKi9RzYz6E1P/heBRL2Adq6pmVRGN
FvOi5JkYFihpmGDbJ7Xh27K+wL4+SrMbT6r0B1gEWo86nFDTmImnOmQ0B4KlQ8sEST6Tip/7nI21
3d6lCTOFfeXw/z851XHtHBxUqN+csKsJOVTCqRxMBqixOSl1bTW6M81CisiLLYxJvD+L5j32D8I0
PpQZ0p/EANVd/NnSYpJdi0S7s/BF1Wb/uftoBCW1uQYf132wbeBz2DACvdDdxUygMyY0KwfqJRY9
7foIsZynRtXNB84ekvlrbkJP3xZv7RzWgv47J6cfOfhUn49O6Q0wpihE3IdKc0ilgg+lm4vD21pv
fz4LWoilImpAI6kO+RhR6j64pO1kTVR9NOUqDegRUacQ3eirLTJMs+fJeoGyIcKwEJbzg1XfZBNg
oBVzEN3L/HKPbDHDnWnHWy0nI72CBMcu9iZvOvx1MahrayV+cy3GaOGMjLWR6E7P8D1rD8euUF9u
CB12c0/JOgn65kwiZFr1WeL2JL7tQwWveulAxDNAUbapDj8nj2kmxw80kzSGkOwwsHpSYVyW3ksW
N26IugapXpoINuecDKCV1cv6X0/ax35HO5RD8WgLhXWc8T7RbifLyOhNT1fXjIMda2uJOt4FlgB4
1SPJD+tYdYNrJ1uiGAVRCjd3Ag7MJjqMgsm3klSxx3lhbX9NnfLe397TTuS6IRG3MKkZnjUZkjr9
EKrDG+bBnOnibDlt6ZYM6qyoJccFIkmNKEcHzU6l5Fb0zgiitt93pBwjPXOw9G1QsaiML1k8mheF
FA7qIrJ430p3rYJLW81pFJZcp1M4X+8qjzTNW4qM7B1Ze3W44sC8pnRtbRUzramwrVBevq/eZxIM
L5OqYNQGxLdneb/7jjreT4tpt2Imo3rN84LjMuG3bcPlN/PJTiC/wRrVIiCd9zhFWXiqN40lZCK/
h9cRDTjHNh9pmcl0DukTQfl9Zpth3e8lCtsv21NcxLqWx3vd/Mu22KdGPCOUv6eXus3k5Wqaw4Hf
I28brk2GVeIh/ZFO/zqsilAOHB2BXAR9HPgv2hkPfqmpVO1alc5NTsryMeSnj/sBhIZQPSv6ay+8
2kmq4WJqToEF72uDJFEUV6nlQo8y5llcjc/f3W1ku0BZoku9e8x9XwZVRqUg2ldwX1+hyf9HeNNn
mhPsaQummMSMlwPNZdoDNq1AbFccTxt4yhUbGzEVxYjuwoJbKBbWNfXikccx2y/KPeDfsn0D+v3+
b/+geE3lbAXltTuHzjPaBH0ryLNrDpbKeUTDKccsxb3MwMY0nhcHY9r2bX2O5s1OFG6yWicBmf2o
SP81fz1dQ+y+YkiPdo/qhOjjKB2nt4LtE8I/i2nNXWaCzZNEBcE95h5ntZcEGunB150Z9PfjRu/c
Bwuw6sIUurcdhEmLmqt2zIMw01+oYJEgTTmnmanl9Eav7+APdGS1rHx1W9r8CKCC0F76HokGeczq
D0rJHy6egkpemgzr+1alNNh69BxpFhWfe8LuhA80nMDQ6e6h01+Jy5B+gciFntPomcjF2xAjVLYZ
0CSYtPLTTQyCkKo3bzQ+pXWBPS5lUe7rB7V28//tEtmzBPipikVtAXiJGq/R8FlfC/QcxFZmQMuW
UUXimrP9USsV5TtzamiWKAwtLiUM+Rvmu4IWJgJsvtnoOewmKs8e6yQVsld6hDUd5PxTINq67Rqy
L2laxaSwfW8yL/QrcCSYTyd/VmlryLRMZUOsFFclbfqYkepY94H7R75iY64CkizsMufCx7Rq8l7K
ZefyAko0ldqcVGSrNuEGLeN03QrO1ZgidzbcB26Ddk/acEXezqpOgdRstn1hX0S1Ps7T7HcXgDLe
oAGt80ffr+0l8okIlvVXHzjb9spGAZ7tX8LGQm9KXwTZ3ZmXp86Rhj4+aGtJ0vhIf6YKopFiaXi8
xy4mQSywRDjz5nV02RMlHa6pMkNSJPjGqJZvLk8snx1+fMTKRs56+WAhXzBX3vRvRtApc9G+pb/4
5tOMBVCBOek3XbTbfruy9cRAO4nVDYRh9TQQ0MXLxIsCwgkTXWegmhBTxw0dif/8IfLhw/FStx6K
2lN1P3dtNX5IUzlZVvtRP0iEoiKIshw4aRNAAVAVkei8CxBrW9/7NSTgc7CDQDXYwv6mJ5RUpahl
UspIj5WYA6G+2G18Gvhk6hlG3togHUZZwpw0rP2Gmisbn4IU5gAyNZYAXeSKB4FWzbS2YBPVyAlR
1wjPwwlucnYusleU2zUvS55EKUCN09gJ8N8BEzik5mLtpum0119jqIQZ0DxckJjKEmKfa67qM2ZQ
xr7R1lkuqO+aopBF0pj0xIEf4I5akVD88k5j2AxJ3kkhP9yG4RlWiSmqjnUmAKz7+dKlZgV36OvT
fhNYve7W5GJ/BMD0rA07h/3QkcXsaMHpjwhrRWq/wAORbGUG+EQlIQRH9NN+q3NXn1NlDEOv9Dcj
18YiUnDHOAN0bYTNkyinJNyzWHm7K3t/EWgL6ynQX9g+hcxOmK9rhFG7sybhjAtLZrev/7CvJbNf
A5/pfpJFu8TEnZfQ0tmaJW3JwBfcS9YC6JaVeSUybrh5al9WOL95D8WDIXCgtTSIT+Pi8bx9dpvR
DUkg3Z49CXfhubwbwPReeWTbRCgAvuj+TCmypKvXN+91XeTHmiNQq6xk77nCHZOp/MKgL1lN9Nw4
eNd3ZT3y+CTs7LbItMEPZM7KaBVLxnhIjn1u5lcohxpxKumrUS4Jks7xq6KIiRZtexMfywNjMo0n
l2qxlx7p6t9mpnbKmsB3PhTelLzhDzl1krBHRMaBv5t2m5E/hvIJOvcu6AU1Ou/324Vf9MNKDW7y
LQSe4odb/Lpfy7xD0Sx2iUuWVHH22U9EwXDTlWRaUfKD7x/gWbRO5txGh1cYrarlpSR8tVKqsQuI
IAA0CtoddWSYDF2MshwB2ES/AclA5rvpLsSdpR2l1EzD1mVB+1oYNkOYrQtRx5mHk9THur0lfZ5u
jjPVApeSu/xQFoIPNx3+Ew9b7Ggo8JYURh1BAc0bvo4AqLTxbnJrQla2btfqvCubjPvZYnFAWdMC
iAHdeIkK1+1q1U1dua857JmJaaOlx+Efg1R9NUP1XNptyXQlDbtlSmKL9mizJRBhREcVMs9pYonS
I/mwt2N9uW8KJL1om2sGDomI6QMNVye/d8un7gai7egotmgkDOMrHn7IHyTDupEi/2zz974s4k1G
7MljAcvW++MtfKd6gfE7PcP1pruTAANP9rKq9QDzsTCoIvviyjjz/1M0Tg1gQcf0ElbiWgePI9Uj
FDKSoQ9aU+EyQYthaU7IvkrzS64THHnYgiZhb6DcEhy9gQqJk0QavBwQvNQLcd85XOLOxdNl38+O
eE6MskZOKh6NoPkU5BDRWFjbX4//FRqm+eEU1E/vXQo9u8/n/FElN7sF5e5M1EilJWV5T1kQ2K6j
tluqb/k+vd3BAGPJ+GxTFrSayz0q06fgZkSO93w99TCCeGb3hj8jmo/MvqAy9IR/qviSlMB9PTL0
Yzi0t+M3W6B/CyCYuFjSEMtwom0GYBHK48WA4ANwmI6JSIs/0o8P4nloXDf7M+2sXWOpuGlLdgHA
AnLyDCBd7rs4dKC7KY102x+/dJQ4Vk9kRztQ8IfWdG+/rhVyLSu7TakgkOdcLEGPY79TJFwQVbcU
UCDm6u3egtWTklong8/HCxXfvodSNp6MJwsau5dmUSUgC4yqJ3YYMwX3Chz6unrYWt8ep5jNGtvJ
uIw6F9xmzXZBOiBP4DhPpFjzaEIZUPWpG268cB2nfw0kn0CPG11315l9/4Ud/74f9gcBLly1oRKd
0QWgkqBI71mS17q0+xfbnRQeZBxELDUJZufSOaYKOOh72JDvhVyW/T6oZFtWGKYO3tQHre8zJ/57
XesFRPuny17S3DTrrsVdbeDbck8cHQivhKGwT1390Mj6Oct3Dsf9QA9+rUgtxQOop4f9mL9/bTL2
MaJVCjtiai6TdWQ6Wn8hFGhGRUh3w3aEnKYrf7uZw25Xpw4O1PW/kd33ep2DL+DnTZKKVlX749l2
H+p1MGepacbc+Hfl6F1TqPL55zB0lGHJK/RF+P4d9gN3VfAFWNV0iGG0V3iyv1hsY4k+L3Daj557
oJb+91b4sqTB1lgD3ngDes8mQfStDA7IuPWbpKyfC6WU0t79KTHbCCA6GV6lMy8IgrxOmG+u1On8
aFU4q3KtCMSkHCDLuprPqfY33pWkH6cJYjTf3Y5Na9BgrF1fmUFe0sktxamglDcs2BD1AU3vyB3J
6oq2izFU5V41VgXvh3I4xpgZwfnjnKw910Q/W2Z1aM1TpnLNckZ+f9IqDnnlXwcaYDuo45Ue6Chi
+oirkNxGc6xmwbnqaikK2RBv6S+EzYbCl1VqUYPncayawNS4iniqIadocbaPl24i7MBHbiJMHovV
Pk9ihHtEFcciL7nAJciElqtDXfMZVne1V7YCxmOp6yQptdkTu8koPXHqm6WMjhktggz9IMi+CgQH
Dlu2vI4qjSXQmo37J5IFwCui7WZHwAfFsTNAGDPLgadrSZZpeTBI+rOpRCU0+oM9anlEJTcppzvq
pXvE/Wvf0E/rOaxLA4rsTVWjk93HNM0yT/IPCPCAAaFrgThSlKH016t5ze5V43YpCi6G8wP87O97
RPWFQwpdkAXo78/EIj6Hnxixw7aI2vMmnOx7LS8ugLo8bMxWadaNzLjYC7I6w3eA7D6LGxK0y9cU
rXJSS32SwtoWKg3JGXs6r01bnCitoitY79YbZU8GnDcPwCmlU7VScK6v2YMbEn/JYydvfZbkKE/8
Ey/L108d0zADnC7lq8udJobvw01XGVEJyWB83cmZl/6/KiAMZyY+l/yuioMiwsQd2zN2BJifRBm4
dClBK5khM53oC5FDYugfAvmwibsSlb56m/DdwCPWARf7UA3HRj7GHfu/+yRkvb2wYlIhWf53Ylqd
Wo/Dqhw4+H6K6zNkplhibeOAhMz+8esKXtkPYYcLuMNBF1zKQwgu6crVnxo/NtzKag8iZuXqhSfg
nMtL1FB1RwJPxtB+Ad0IGrs1NQgy065Q31Lodh6jZhq9a6rhwYCjRMXa0GjoY2NrOt8tL9NUPYrB
rEOr8pJeHXPPkV7OalP1TlQz7/KT4afyJXrTdUx+9aEfRojWYyM1AkgMybsFJTbZvvm9+t9ho5MO
xcFTT+KPbfV6s9PD4mZ5+ytkU6VTs5SoXbByxFwVbkx1GFniVUf8qGQ1mIUAU7McVObFSxAXUlwI
xH3KzrplMiE/+KsoWwR7/6f8sY4NxpPn0kQJKUiXltVgTMDqwFbG09gIgbiRYIWm3gLNa7AK7l7g
VJOFspHYBEh+23Vy2l8mISrc5vKceIlfDoHTD556xlq6zb0E+O1R7PCH8rgI5ond/RRGNujzbQLn
MqwUbo+GBxGk4e8jZRxigI49QIiUWuygz71K9xrKjTqIaIwBGdIHV1Eluk6jLJHfW1oysdMP7eg6
BFAD42lZ6NsBYBNBGxjo2hSgWPCR7pO8Wop8PV3uwPUgFHSPc9jiT/lGEOUW3DGl39144Jfg1HtA
FwxpOiNbneedQ7oZ2dhFz0c7e/43pzk8NK/Dl3OOL0Fj2J/48vsEFCCMg2j+N22Sf9U+lP49qpQL
yYWdItYSOF8mrWswd0Q8grmzNAHO/+foJtAvOoMJmbYJRcPS7MIH3febdNaHnEi2pppoaaxqMAzd
otrLbdrJDDnvbJozp9u/BaJ+Yv+UOyMyyFBOd9Hfx+gr9uk5tf07qXWiYLWsQ7A312g4ElERWPmm
t8JvG3d0SmIQxHJZXdNWDZhvYs7gzrYEwoC33fsHApNIiuqRsiTVg9KNoUS10VOitCZXYkDU3idE
kqkVR99B64QLb21hpTaZrvlXbmeHYIAhV2ZWx0riYwOfH300Nb3+GUjlPkNkVHaDxqRiFRUB7P2k
DH0fPNU4CplE7CkER9iv5X76NDCiuQuOlvvCoSPRa5TGNEXUzwUu0KDrs3t9XKwcSH99HGJfo/Xx
jdC4G8UCRlPBBizfp2EUpXhou+F50GqXAPjid69mOrnFSG4e/6zp8ozHsWdjjeRy0iBKGPM6nzvO
WWWhOVBvKtWLjKukGDwLynEeWcCFl0gSVgzXKsr0z3vSMj5FugRbmcYStLSmZREu99Drgi7aND3+
Q2LziGUSQyCVOUhFi8deiC8BYvtG9/cB8F+uO35P+UAk/MAn9QG4V/H9La8vLKtpqtVdD3E6qX5z
NZafInl6Vy4aGHjhUY9RPn1pxz5DJDE+X+goR6zdi5MFaEHIL2i0Dbz2Vnqhwesad67ERARKRzM9
ScuzEm1JkTQpQ6dEaFx2ITBcycv3aLXrkHrOZoSjDDSvzdpJR242b6WSIUTBbWGBxCUjdSjYxIS3
5s0dML18RqwX8W5VNsPAfJIHXPT81j9FNZFTss7LLI/TSI6NCwuFbha75QTHPzeH/9KfFismnZfV
A57ED8G7H8xsknC+GewqfS/OorZ/r6sU8XFxMOyQofC4wh0TaqS7UFYrIO3NJ0hdxkpz0zYV7qmW
jsogLjAcmCHpJHOEkTv8VBG5O9g2T3LSRL8yw4e6rf0trcmdVx5dQ/05oN0+Kca9nO5zlmMdhINd
qIRMiU5hhfOM7sv1i8CHuJjRYPnpwkKuVAdP0yUrWyCTN9vdmtgXfMHwUtroVIafrvDLA+lSeArS
9biNsJaWYkSMIeN9E6myh8nY1nrcGuFHAdWzXhSu/hof0JLjnQhH5T9Via63CqTFomgHI1mg3yTS
tjaZqmbntBId5WeefHud8UfDIyQMI3tA3mfLWu/V9lW7L+/hp4RkZodKt/RfjdkNS+1gVcUcIxsv
rbmTcrhS5LG4ROtAjc4ziSgneV5KsaVBel6pNPmtPTJJqQeeeHgsBWfm0kL4H8X3xfvlUhsLuxRC
r3vokk8xXW+5H/PORV2O+Ba3nQtVAfkzyHJhPsbfFVIPM0UoRfjZhIX6JETL/eqeiZCFV1PWpzBJ
CQ58wCewM6tpNsDzj+m72kjKSXX1o2tX7sZbzlXa/0T41n2EaqAGQV897CAXv+t2o+PtckOp52jK
AtPgB+SWXrvmjDie5IDvNic7MleQHxk3b8UDxM6yVp0yeJuC2r8E28+1LagFkeSGiAfnX1iKD+fr
/ujAdrmvcRDRVN3g9RmlsZImc3zS/SRTGsV6oiazSKTrVGF38csuzP+goIaF0Q0XfT8iw3mkgy+V
9z2usJ5KvJ6Q/AG3rT3tvnDPBXP6RD1y0M6dECMGHIjuqdTyiTfS9Oo8TVGV9GSRonvRSbIk3Dsr
bhzbkSv5DWniWjg/plgHNrneMI7AskiDGOjFpGCNC1pvFI0TuWk1VIHxmmqtdVqi2PoRAvUoSxLk
6OgssljAiQ8RRZchU0y4Rp60f36AD6v++y5CGeFrG0ntzwouBWWHIz+nQ7y31ietS1vRUKTUpHg/
qDYtSKYBqchYP/Ly5wLOYODMBWS9fG2RTnACGPrlW7Dw2mBo09G0muCgLxOpKu1kgkzqmdHRyVSC
sv5Pmogj7l3hpnnECzsc6Ujpvn513MhiHTdO6UElMjR6YoDDe2rKCTXN4XXaB0cF53nbs1HXMjYv
fsMmREYPos0RP2vQydQKG0POS9uMDzsahSoLhamN2OMtbyBVGyQe7CCrEmxAdPMlc24EBregKR+H
gVC4JnwTNmQN8DCgkBkq436FQ6V+i6DZiqVAfM1P7yWheDi4o9Wk1ilWkzcfYQNMnE9pbtYDkfXE
p2y0gOxNXofBrNPcbe24f42rmEOKkO67lEF8cFrvpQgAOp9lC2uBdlIQrudPsYVLJ47FL5BtoYiF
yWkPo667VmhoIcERIFcEqxz9Yt4euAr5Rrunkcak7WKUVZk6s1QXB/hlTNzVE1lJAuz9N3EpPL9I
W889wN0mTdAv2Ux18objW9ToApnWsuWlHbzoxXK2xnXFx9aLnwe6o+lsHCXCWqcq4nCKdR3QmsY4
sbyaEd9LxoRrUFsCSFKLncOz3byQLFZXKGappMLDWOX4OEHT46V+OtgRQAtmD+NKKZimcRVDqLrC
dstVjo+DnXxuNS00lhPAXcKSb1AmOYv6KBQNHuVHhg0U525iZSgaOzKmINJe27QRtRmHU4XVEAt9
2EJGxGPtBVsPLTM8IlCua2WR4EEB2zcnaJcoDzWKL77DnM1haLLzUFf6tHNOXMANLi0KI+2d0PaU
bkQ4/KKbSAGSZRqIqY/9a4CiQssAsCsHduIpJVfqTlMxE/5dVQC1GA5nQ2BEnGshJFxp19QhnJXO
YyuVT+Q5rE8YZ9d0D7TZXi3i8OuFduvc6ayI63tPuuA0RqscQFKsqPST3sFNtcACUZSUgpLIeAx9
F7FURC8OXZAYyLnOpOOjHbN9y+nsHJ+yVBxnsDS31/LgDJHq+lNOeM49Hld2SPQplD2Sp6Why0Dy
3DKV/slBJ0fJ5nST3wPshQ89YnRGXlvK/xGfXpBBdgdgx7NCKw2ZQHk+kHHhwrZAse4SACJGgz1a
AfIc0WdYBM8/KzOP4cDHg1IKM2lzQoUYnRawytNyKTP0rRESTtNgDMuDveo1bi8bcM9BBtzKK9Np
+5hRCEHtqctxEVzvSprH7otH8I+RbWMWXVs1PiG7BxQixNXct5OxL9x+9pVCU0d7UfEmqKVdmZhG
i5djX2jOmAXh6HWCO1UWkHAxKV6/6QxByz8V6NFGGH2QkhRFXY37UfogzHMC4M4stUxCPVEh66TN
xaTlXPqOdfXLu+UCxOn2LTT+g1xeeje9kaH+5OzB5J0pl0mia8vvB832Qgm50KDZSI+35Ud7bx7o
T83fbiisenviG0v1Jo6+Zh3MT68x2MpNmJ+xGrz8H3iAJjTsWNaR793UNnzUVnUnT0wi6Zjg7Zcg
oRCdygK9nPUPaQRKsvHGE6lapN2Xn//jHGP3D5lCMTazWws6wd68rj5S0BIdAQNBcGPJcnQzZZ3X
KmmGGLbo9q+7x0CaeenF4EixAENdk9PGJADZWlVwO866Q1Z4R9m6xl2xF4dYTRnyYqkQtSIPA0D9
EKH6ulEi5h5ZJ/aRg4WvYk3AxX0tsDUJ5vbL+IxRNjM+1kyhhLHs+SAnE+1L/A/iI5XSOcD/z7vA
MfwTUnthKCytPK0gpLktyVFQJG/W4YYALh2d+iHw9AlAN6SvbA8rfGPbz5jpMxHnYOeaFDwTES0I
vcS0U5HpsWAQ9WsY5gI4MXGBpzQx6kq/XQo28GP82eDujgBvWq6NfNc6rKQm+aD+YPR7ZVJGXi2Q
oA9yBbr5yWEXDVpJd2CWLCxzEXtSuLprqSM23psUaa/fL5onkBg/tJglgHTY/MZnN61ugWidH3lZ
sE6MW1j/kPI0ERK1WrQJsyDYsCAjRTcwoCwzMuGI0/lZpv55HuXEqYs3EUxZEl5fMG3agLIB+qr/
USDhnugoUhtGo7GdTYVATFtk5jx/IIzHvVwaetqwNgHO0aNFlO1dIjPdmtdbLKQS+uHhPmQ07pIr
N9PkDwtc9McoPXbrqdgX2+uqYKTU1fihCwFA+It/0R/0IBOoUWigluzFjUl5fXGc5HjIohOk0q0J
yVYDsxI/pdt79utLq+n7F+z+LO7Kc6WwSsJ4a0+23H8PrYAf7KkLbeDrTQmXrMK+bbKJC2zqV0Jq
r0/gGguIbpkXDw5cuvXqmk6UOmh3X9JcDI7uPdBRlW0GAdBDs0r09nC3FDAg+GvW4CpvHxvPbFyL
zCFVJ8px1JTeLzuaEehzlQ3Zrx2YEgxL2CLYNkvJD9p72txnALuVmysoR3fgG5tONUYMRK3geDuH
O42Bpy1TUNSP2rbqzDCRgOAbkFl3rOF9cXJFaGraJH/gJ4J7llt3LKGZMDegGtgwjPt9AI+K9ZgI
Z9DIlv3LvKc4fznCDCu8PaTDzPBXiMiqxuShgjGzN/Dz9AQVtBoNHyGlRW84ooU8gDmR5gAA93Lc
iZrrhgcIoTnpBrtMKbyE2Gxplp877N6CgBM6ILrS2ARocZTC46vAswzNnaPNWLKyQ2pGukowueAl
Dl2GkkfsybcwZgcMqJUDFIQPCP3EvcFZMTMQhPFx5J1O8WNxzCMPIpFSc1kj0Y6cjRDz5CqIXELd
fpyvx0yqgzcZvMH98k+E99BT+oDPXklxTWgwOoBY6IjwOKWWurKjEi48ZYd5TaGuBZoQTYHAls2d
PT+EzDdzr9PWCpaNsG1wy6XiGE2G60gc0wIkI9JgDOxmNHdRorfM760ZxTnUcJHarlGLYQVuVoPH
f/N1fdopU4EyUvP8qVqt5BqiBmtnooH7MGeFGgGb43crGKz3IjdB1b0nKFV3w/1AvDuFfwEkFFDk
oAQmF4iVDPJYpDT+mX/ucKE4ah60o8Dj3IdKQ+2Ak6e/csM252PbEtbenSgYKvUgFXesuvUO3+Az
fw161l+EEeGeJDndG1DmHLk9dgmsGan6m/NjIyXJR0Q97wNag0Z/0taCCJ6O2ZEl2Uffk7VMLOL+
PiuwlNXZNAwqf2AwmDvdbEeeLhYogolpLXqzHDHZBlFFuAgjrrAj+woDLZxv8an6piicCDk7ZNxy
hy3ET4Lq//5T3h6W5f2buVE8BCPFfzY9oY38j6Jqdcr7mHgWIq/Uqld4bPKKTtkpN41BC7fidpJB
cDaaRiPgalaDHIyTOjvrg4KjYJXqsoAlE4MldrQ3XOME2X3S32pbYuIcl5YHGBVjGQpkLqTWbav1
tj+/d/YLyRjq0rtYzDnIz0eimVjU1sKATHesCLV8YtSr5SaVInurmhzWA4gXMv9plEz30zfjiq86
d7zkkiW5ppG5jse0klF7AieoGoJMoWRQgPNBE6bYVAZN7cBaDxPK73bp/Z4DmW+2sWFsjanLqx65
ufA25FrA2BdYnUUtdR3SiSZKLNIQxvOMR9xfIt+npXrDh4yMEVj+pfm3NENiUp2L4hmPfJuCwlrp
/3BrjH1OPedEdGYX4qobetwhPie5bqDg6hsgp4n9GnpHqNOtbOCeo3p2kWnGh05jNieFY54qdpNL
gdmSe+aRGDHvoXUzJBsNo4FF2pOXUhlOHmWDkvDE0XwjZ90qaLRXCMCdlMB1T+ihH2pVHdyEW41S
GvZAgKZ/1JAMXXrYmbGgAWcl9jHRZFdB5TyTW6Qsn1MKucI+ORcJPD2rzanh+uvbnCkqKP/6NdoK
wD3QTPBR8E2cyNyavo0y63mNkMSJ1Wc+DxuGfVsvrxvpCcAiXUYTJQDyM6smuL8zemSIcrf8ZWsT
liq2cueRRovu3fkc8BvYvMzkcqmSccwnXtwl/2k4O8OiAaJmE81x54586vqFsUnqSACpl/YYYCEY
BpVaLjLUmxVKk8+RJ3reM1R3KQPndCIuI+iCfk+LX8I5eYFKZWBR4DgmefIfYc485sfklnxoR6sg
v5BkEK2xTYir9rs9rtcaazSJdVN8K/ZGWUpSnFMFxhb3a/y+REkc03F5auOE+xycveKkIGIyCj0B
M2GQ8CUHIwP3GVmgsvIW5yEHflXWQYs0Miq5twJvKxr4ZKw8CooOoKKVRwYFX3C/OjXiJQ0cW3bp
K4A7JmkaAnxgMnDsMU8QyfG8DAQ/dYaAitMn0AEJaUYhRboWhgx8D16KIK86HH/MYm/JU7N4bR5V
WLzh91WfYeyVCYTbhVVLcr5+y6gpF4puX9+bjfuMeVDTh7OGjxpwhUrv7sWuFox8Ru+9j4mPozsa
vMaCuhhJMuA7IjacCN0oBx/0QdWKkSdUmnoIFl+Xudae9huRrVbODJUfZgmKE8cSNUK6Mz5sZqgb
Q+s7bPUaCa7V7aIX+NhiUKbpAOXwooEb8Wai61qAmH1xCSUBsGzm7C427d/Mp6x8Pzm3PYLwifk6
p3Koy+DYVYmiq8YROeit10LfHfQRaCGzHxaJEYNVBVCnPmmELX2HVl8PE5kiE5YWw9kMlWHULGm8
pILPnm0YuScsn19YjhTkjaWXsu8HOg8B+b5Aaz82QCdLPLjfhnSyGpxu+sZj2uc7/72o4KG61t59
aVkbRoPVNDjpFEuR9KZ0tW8No5KkijJr+upHo8HiA5/n9oIG6mT2/sCwI/3K2BI2QkF9+wd0M2gg
sV4e8MX4pQPAyqX7TsGMaO8IzB+cBHcjYKXOB2no/8E2+pILrXWMg2xjOfqd6b6z9rW3DFzADOY9
wCTrBJPopkTucLjTNBOrX1l+6iTX9plXxyECmsHTm3zSnuNc30iTgCbeYzp3PiWuC0kpB6XOnxV+
6CVx/9unnCjDKp333rZ/3mDDy92OTuRlhs/P71KOBEa3nNQL/L4C8qPdy5b/JwQOcLCUil1JlAmJ
iiONhg8gEUpPKZmhDnpy8iU0was24uK5bihkN2aFkMBYIH4AL1gf55+4VaLbrN9NDtrF68mSo+24
m0IrX13aaYC4+LBeJl7k75WS+GPZXZk5cMVUHtNy9Worng8dFVqnVLn3gm3Joasz9JdnSes51r6q
tkBQh/C4ZdwbyM5DL0rKn8vAVcIsJoPW52xepoPFBuh7l/syPhhzXLjCjVlQQul0CcEABOXl3DLs
nrKvN47WSjdeFYpMh7bBptRm8e/U1k8OnKc3TrmxfyWf5LAoWTQLfeCRs/GM9qTKExXsnLLl3Hrj
qTAKrPv5lpzoxeN+xmr78RjurEoRXZAKPkY2yJOnfgSUNWMJs7SJx7lrp0wSosEGLQUvBMeelMX8
FCMEJImgx1s2CiAicP0cfx/Cxq5tYloVUL2zAMHSHG1bM+IP1pmON/izVHcbPs7nm/bSr5YPHRDE
qb0DvuR2PappsxJP2qX8TtJHILsQ9Z+UHMjhtkyut9s8F3QNoJZKorN9yOYC14nzrAaXGEU2wAtg
xYZOpgmHoYT1Ql39Veprom523aYfs7jO8qyLh4OfWrT5IGvn0z+V06GpWJ7SJP+Kr8PbKpK2Q/Kr
FtY2Bp0DYTyPO7gmIv/UKA6GKkohsurMERvVNBmrFZ6rVm89RIMA7KTUteHakjyfq08KI/C91WvM
GkXX0G9nce65rIg/dtcNSdgV/8KylHfg+GWbpRp/eE4DNcH6g8t98fHA4ge/LVR9mh03gkATigWH
aRxkwMYmdRWTnVdDk1OwuXmLm+vfuSzob74mZyd15NFiijqI/y6+RDvcYKz94opWIs2g6gG7gux5
/yXzV/NzzdBtD6O2X4p2IBXts+C2WwPamwoUB5yOF7IGsCAm3BlhNn3fFCN8w20Lmhaqp13n9Ozp
RxvGi7OaW+3yrkjz0j2ZuaIEFyIf+yZLlzZsZ9yNVo5c+uIfJ2y7fLy61b9iWE45tJaAlTbyvqrR
fZupPeOLXTE1ZaqgBI85P/pJTKg3Z6VoCKkqcUp7tv7qCl+hd+OcS+6m4O9BHGWkXPjHYxCRHabo
2cjNGgZsmjeFSdIq3/WCB4OdF6JoxoN1J+qhRMddjg0wKHGkf+trKmXeePJcaV/hZpvunpUUxptP
66TtiblsQ/OGdQ8rOQdmlAqzLKqJztm88S25+XwIv5sTqKa7FDPtzxQLj8f7ap4yuRl8uSGmft3L
R9rqEMHUCUdaTw5Z2Cz4ORL0dpshG3vAxaXW0A6LMntppeaAFWUIXbsW0yu8k6c2e6MDJD1g5YJj
MWHV9DbQFeqVZruVmG/CHfhPcTAdLNO6h8+2+DLSbYXAWQp1AK9cIx9Mpuxfpx6ilKnoXxDfodx3
u7cRaW3vb2ihtujSjj9iF/z4RS/APygEUKbpmXsKshbq9/ZBqqL9EEMx8H2HCiP2/oJbSIfh17kE
PLAgu/WNlZhB66K0xGWbHvujvd5/thDRwjCuwVPr8Lr9ohCbJNtgy+JwK4yrLywLmITj9tceKe4Z
Yhd5aQxwUSrPD+Oc3HVMSx0eM93x3bP00vH4y/lDiXnuRnPDx7DXtDRnCM/7PKJa6i4nekU/9QO0
m/Me548mrqnP/ejJfoB+PLblzLeLCgoaVu7v+p9yVfY6yjgY7AGdRlip20chWCxCUnKRfXcuWH/W
Len0LHVvYiEh+Aikka6hRhZ5vfi7BxSfM4LPaEe2PCGWcgFyufwp2eywyUzNpkGza6VAdsmkbhmW
QVmE9Q4CmkgAO724NW1mcIKENdanRKVyRPBeYVwEsNZncykDIgvqRNnqBe8k/WG6SwjGQ6l/KJ6q
ogOSWyVkx5zNWjKCCqjiU3ec3DCcuGS3ejk5Luk8hfepivMca0TbquFVX1495A/qyiFn9CV1dcDL
7ckbaHGeu3VVEeRK28ATAkvRZgf8XMOmiyruseKbYydE6Lb+uggRGiyi+DIFxfyHXkrSvA+pqZZz
Wn6pM03yVlXpW6BgLpWeErDGOGiHucI3H64/0NfkUUbybMwNN7DnH2WFTOSdMAtxDu3xtcGYJ8Mg
9PTZpgiRKs9hb42v+HuHPp5kbBeWJ65QBc8IyaWicrcY3q2WU5XnMBR30Lysz7fqkhTHxpf/4rwf
YA4l0sGTY+bcGLUKO2afiXnHRSAPg93vBLTxq1x9Y61QJGqD4dE5UV5sn/7nE4K9fyoYXAhJKDnT
5k36AqQdAWy9I0VF0hN1WM+PRQstMSoewkc+SAu//BzrS0Di1Pzg6IqU0HNDlrZNpMHvLr0ZijEi
0oZL5CZVYrVaRgiBefB1Su0j5PdlRN362TXCoCUug0lfLzadqKCldujBgjANDW2vmOYLpP8sLUJw
I27w5nHo1NZt+vazvx06dFG24RjtelhPS562I1ODoOv6eFk4Hf7sz41Drtezxt5SqAOHIeFF9P8O
+hEMcYSD52MVCzTpa40+ZvDW7RdaP9VkVDS/IkQJGYTCO4DGbJOPfOpAz36/lgCsZkS39QROROuZ
QMgnFV2lslZohpRqDJpsQISqUkchAPHX19uZL1XzxJFK99H8orfnvb9H9H0q81zsmg3CE4tgrgFa
lYkYXi5LOLxvintRAOotir/iu2pLMYU5PZWirVhWQdEVPNYZq5QgeTM2wcP6SQvsVSPegQULvl2H
vzHFjczLXeA/bsfMW28Km1O0B5z04aADl5/cjgL9vLPqD2F0rAIgMEwWHqmjZTn/VG+q7wwNlYQ8
DEufB0Q4FFtq5nzWrIeZ/dtxYgW+e+pwz2Ptm8JGpQ5I3BSZkhDa+JLr1kn/3mEdRATCHJqgqmP5
AmIJhZkMc+4chSnJbFfp0IJrN82LPDY956fhzmqdQQhCHjkpSBGF0CPDDnl+Q1tZ+Q8sFsPxuEVA
d7B34q2PzKeekQZ0L4a+l54gEk9V9S2kCme8VIKIxDi49/MxxnoeQlJIC5aC0W7Bx8/T1isHTD1R
ZclTErzdqI8LXdn2GWgsGuWtP5lAeTMU19KQ9nR257SCQmNDW7EgRXLb52rzrYfrBlT+VotQB335
p49xgMWuBSWCRr5wAl9BUlVOdqoCGEIYNTwBT36prjMaVVZRcJw5G0mRkSg9bb68dvBavGidQlUr
LxXj11Mb4R/xnbhbTzZsC62vWq6DfYO0HcUldYKtnoxhCse4Ao+mFuRJ9N/VRc3Cae/M3qo5XwqJ
RL0lbhvdUvLky2I9uw6rgavdSDH/VW1mkkA21iVxMIp19FHBfwMDGhBoZBate7Fn7UwfGC7dYn0N
/kafHh8s3XtMELcUFX6r2HQ2pe06QCkwQxXtGLoU+sHA+Bnf4SBv+1qYCZs+XdMUd8Ha+vKrbLM2
tG0cCO+l/jVW0h7ia7UO7S6pNxiYrjrT/bYN/Q5NGu+Eyzo/nfCY4MPRRFqDpVDswwaWDcbhZJSV
t/A8YCqpIP9+9h0RyNi7opujcTdCIYpl3o/vAjOIzMENvRO34FqEZ6J2zU7zq31kA01N6fkKpXSd
Ue0kNQ+aAHHQ4j5Gywj+76fLbXEcPf0A5kcBLlfi8nx1wMfNwJkYla0fTWlIiJ7DG6AsXcBZaDtU
HGAM6pea25EkOlASzXdPxwkDZpzLi/Yj/BmVF6NZYBphpl5tO7jwTKNUjkFlR6b7e5lUD/l+6gpi
OShJ11s6k8+tXvJD7cKisGRQoz5lVTRVv4GV6R1cCiNxpbpUyU+loyXgYWsAJKifJz7wYr9FK4w/
mkbKPEdSjSXdbkPnXrb1Q1yvkViGMHI1PQdGcNZfX9FH89MnijsVFTyYOxlXvIT+X2LyjFp3yRjj
M5ECdXIe/Tq3xEET397E6TOpVnsqPJS6OLcjO7Z1pUrl5cW4GfosvDmxeXzqGowMNT8ovUPd+q2S
cK67tI1aCJIW/KO23k+d4HQyAzYk+0GoEOsKlmKT0xqZovPGKLaG1fj2pgw/QcUkx2xgkUmse8jk
xzwfol5d4+TXOY488e9FF/TseC5tGQr79Cnx9VLyxyc3yuOrUKTEnN4S0pI2bT/N7h/xv2jSQvQn
DKeol8JeUZMBnU4JlNn0TkDz5lC7egDyd30h6TNTL4i680bLJ3d4psP8926QvEyi+2636N8SeyEX
d4SL31/+Pq5cOVw1/8wVci7PboyKuhh4MOp52qBVs2I5VNE1DMweEW8rXVVKHVNCQwhnC/NHx19M
RPdOka9502N+y4HejRhvjEvnwE8VONa8Cc089DshfwXDF+XJpwUozpfoMbuKJTIVO4I9C/HDNdxZ
+l73aHqztdCHxtyUtJHOxWrOuSkaiw0kdvDcXH4JhooCJEQ4LTGN9UiTmxdg3FBrjVSbhC5LwQBH
UEDZ8Ifqc8ppdcLWglPYON13mt+BXoG0oZbEp0RFC6EFik6TkUr7SnXcaK7ZgbGXa4LEs/WulM39
qJoDlfp7Y4MKyq7QMuqEy/68a5IPCtmgQOmdKbM2vchyEVVL7+nJwiu+l0vzBql6IvWzbjdNjoYo
00uylGhCgLAwcuUQ0Zb4wrE1SgwBNr8ncgsyQ/RTygISlnfX8RVJhPDKFwUIhLc3GzbfVk5/pk3k
RCM/Z/3p1FAsin+usVX9X8L5ag90ii7GfvETUtkhY1IFObfwlrQRo6J5VWrZTnJHQfdIG/JEYh8q
yyAXSFRUbkGX2FdHGiGSYAawS6+8AnCsEhNhe7g/jk5Eet8VKZvEstNXEYUbShh/g6J3BXMpdvv0
nFPg/K3O9OK+515LQcmolH7odof/yesfQv/uk4KhwCPsygIukPCAERj5lsxyRkYn9e69/qlkNDjs
x6TD44AF6xlLvmMylvJA4ltEud7t75fGHR1XRe0he1PwI0+LYnGlSAKBahGOrJrby0DXuiGG4rhD
CpO7weJ92dZugua+MbLlvM/gfMJReGDOO5mGLpM8otgS1X/liguwmUZapSxa1ZPMEV/MXzABKB57
/unkdld1pVa4JO6mk9vCMu7ldYMRQpwxM6sAfGUswycHNUwi+ZLD0KuaXTjATgfaoJuwuTTzE/Nj
7TSYqOIieOKuTXFjtP0wnORKf1n3PrL4JObDBRlmALpMkkwLfZfgN4q41ByAVGo944BP6pXgtjmq
Fzs3CPQYxFisxND00IIQ6hAeWVuP7ACH+1b2PEHcySPOo/nFuEs35BLhhxPFrV/9zb/0I5yU8CBV
CfbQUHFxD07po/ZWwD2KIWlbp0kUGW6vHbr9B59FyU83GHN5Vrrwa3nC+kR43z5o12TA3hjwtIcK
E4tJABeGgR3v3e5VVtGdzIRRYLrPbzDCank3BC1LQyNEP0z0Ws929kYml3EAGSqcR+zH3BNJxs99
NFJi81PYhuImkfubSHdZ66rAVAguiVocJIhdS8ePyf2eXVVsbjNJl8HhPjuItvNnn8gsljJls7ZC
U6YMG1p7AO3/Zw1ldFndGhtFVqO2A1XhQAbgFK5gExjkNg5qZrFTs/Pii08pRm8OaIpm7eole0rA
yfcznBkpk3I1Kj/lgZOzDIdaS4y3bhziwQlqWQRBZWoq51EG0XpY58ESZTb12R/WUxwBX3+DoPMn
MDtf7thuxmTV+JMfBC6bdb/Tc6ymltJkNYWlG+x224EGCShanGITONwKuADbSDGr6os0cb+au891
/5xuvwxprPAwMB3vF7AEDrhVRS+/c9+suxIRptax5on9wcotjwPR0TU4wRN89kSIe7KLzTT9Qqhz
gOpsloeQRcaGQiFc5vt3eBg9HFzIYGjE7ed2Jt5AC+UYoyI2M6nG7h/3p6D6aauK/eTrG8ob7EeF
CKTU/bNE1NcibxzJigEuMoi6D6ZSFP+GLCZYT4+tVylYY/YEDMwz9RAr94C4rIPCDSPqnAayeyNh
Ji4wyjhhlcET3lKohlw+euJ0GNYdSJH+2pSjnbUmTDe0pMdVR6ngHLNJVpWhM2AjPHaR1YQETtxi
oiNEeLYvLh6dSyt+7J5TKDd1hvX0S1TOehg4/9aWFa3pyy+MOf1cCSqIolG6ZfMyfcf2h4xaPA9n
+IXBc98CV49i1rMknRvQrIXEYVqko5ScOGKJnrqj3w+XocDMzmSQ++DWeOlWU56idSy+RTvUIQ3G
aEW3tTvrJUQ/jvCBh352
`pragma protect end_protected
