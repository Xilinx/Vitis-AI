`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cpmLTnckjJLm/GJhnEEySb5724
XCmSymMTLlXyajuUkv+nefl4yXy9x2yAhXfBlAkKJiYo+BnqQEh1UNkLqYAA87d8AoAB9ihUb8s1
IgM+IoyPR9o3uY+NiwUbJmA8+WWguyhwiuI5cBoSnntNWESoTGk94tPn9TbimmCK7vJ2fB8ppcY0
dzN/XzQx6rnja2k1n9Vpi5cSISAq+208kK6KhLcxARN1Di+/5T8WUJbGsQIEAp1zBaKpFTX5V0rm
Ql3304+6SyjBQG4K7CBiQy+la68VMxQ3zao7qFqLfVJYV963qTnSbC9D6VZ+A4wkc/PpDt5jLasO
SDtBN9Vs/Y3J8mK4ZGHuWXzIr5NuLyzm1av+8WX7K+CwfuSAKRfSaoxX/HRF2Bxp086BTZXJGHJd
bOaLjGh2g/wGj0aPSBCuE2BMcPzFnYfZ9g+zaknmAYKF805CbFV1UL9LWMswj4lYjXdlrkTRriJB
X+ty4aU1XH7cQFvy9KfSe8X0MYwUOB77lrBCj5HsfAWSGxAJohQvqGUd23DuzzlbZo7EwtdFwuPd
aDHSNlyXZt/3/TmXxoNtlAYmVC6rxMbzGZL1W7hpnof3aZF9bd5bVai7hS6YycFvcKpVk38SPKDj
htRAP50OyyJyC1LCvdrWx9fKAeG1Weh81CvJrNyemGn5OCsrp4LaxETLsJKdUhY78Pnoa+ZLtDsy
64VUmSESHcmI3mUKOtdyVHDEDQykOCp7Sp6wPz9062Px4RjTEWxG3sC0YJptsiBIlKjiBc7r909r
MUOW65dbY8MfHSr4y27a3KAzHcGtHQeWm/RlcF/oYpAXlBeQK7lJ4z+TqLbox4dwBRXsyViq9JkT
J2D/IIEgbdqmA3tQDBg/AEGi8IFBo5F7e72x3T32nT2tPZWjZIwFj9K9jKwHVST4/wrJb7RB/bjG
auzEA3BN5YslDsDbRRqeZfRmAO9mDSdJrRhr1R/ymAajBIUCQXUrX6bAFfidiACfUHHEh8U09hEA
1ZnhJAw7ai+8HyjMXa42+493qpBsKKyhcjcwk1SUWmEiVH7fCTknshdCHcFN3IFYLh5iB9F0xXOa
bwcmlWIptWVXuvUtmF8WmDC3iIQMszL3OU4LKSFe6QDhZFT9Yd9ydR9dL6sK05lQyJajdBVqqXK5
H+ogzTqjt+3mBMpl3OmFDO+9ouOYxBsVHJnsP1+rSnosRTSOSgzpzgcR7e/4Pwt04iOpX1f0zb5Q
Zr/5pINXu+ylRDi6mXtv38o52BBJ/PxzlliW977Apz44UxnwcOhvyR5fHycc7SwUK0SgOWCXqgeQ
ibKhAy/iQYLQZH5Iw08YcRQHkDx7pi6K3TLwp+gl8cKa+Q/j0YVVNAavcp6VJM2o2NiZ5VQ+M3kg
y42sSlhmFfPzUOXqNuDPdFenApgxllB8VESDg0UVYuzaqnGVwuih1gqY/RcOIaFiPh7wGPSEcxgX
U8yd9kq0wobb2V/37MLmmmSqxp4nMpKjL1/cPPwV/gN46KsUxuBE6GvxtGNaKbPk6juoaxeKJ3v2
Pq5uzNwqLPqd6QNz86XXV8f3zMNdY5T16SVj0Qttd1E4nIwm+lZ7KW4xOBuDtKe47Z028OOfn2ci
mL21IZFTjuXEFRBbPF5QU6RGsWNVX4kmePHhPugLQnErbrInfDHLqvL+jdpfhtWaJZJqUycodAe3
uKpwArsXvmVQA+j9d/NohedIllN7qpi6pQKgcuBS/Lqc21+LDWN0zuxyB6fzcfF1gCkFJHxtm1ax
vcXVDhTdCijhPDv4NkjmdvnMHNSn4NXuD1Uxi79/vN/AsOShVLNBgpIIFUezrzxXljBpOqgPmYLa
lLIOswozNyZTSyGRAVfUgSqRflcJog1to80jrj63e+qk7n8Q15BsvgIm0O70nNtZt6Ko1I0Yx64u
hw6EPAMcl62+pMnPBJErD3KLsbdX0CkNSD/r6QCQZVlBjmjBdVX1Q8goCwTmPtzlXoGMycWs7zIZ
OYeIgKIc2MfDi2brULUdSooDrVl76qI7h/RXnwmNQDF+APQ2SIfZ7QzufoPLY9zwndWg2zWSSbN1
/LA/q+6onQJbWPXPSUbqKvUGKQewbQQvhXDEp1mRbJxofqrqm3etg34reaI2s4T7ojKrxetkbpic
cZKAfWKZzsT5uB8a/bjv47W/FtqcPbG/ArdYpNeOxJpkLOH/MKJshQ/YKcIMiPsAx/xHBVF3SYIc
k4bQ+/EyS1y1SLwtUIPvGM8Gd5qj1H1Ev42VIJi+uxKLpy+WK7HarA4wWsxa0RzskncitZjvIj6c
u0lgVsDJHFblBpqoFectpCGiTUudIjvx9xucmMQU9KbTNo8D9hw/WvaQjRoaO28Exh5TplQ5WOy9
KmZm8ylZW03v+lWVE7DFLjs+0AUip8nK+NaQFbzRa2JTqPnl1vm0R2O24MQz1654cgxgsDmekZEs
3JZPPVFRHMTQqhgSQtaXpDRdSAP8kakxHkmZxLPXBGB4Pl9csrDJkUyktYmJqg33ynR8WeO8UUyv
VwEjI+Dfek3GK2VWXOmwb6lKqWQWw/04jhXrZlyeCX9jYxcdeujOjA38Fs8PFeQDslKftOHBkyJx
nl2rsBea/gvRVGjWlXZQVqfx64EgIRjDXuakLLxQ+6/Zf1wsY0LmUJfUTEa1oENRGLZPWGRD5RMV
2NjQE//YWaU8dX1+GUaZKgI6v69SsL0/k92WS0wCeXVGAPD5hchNztJi/RmHMU1M+4mrtoQJbERV
yPFsCnAX26Ls5fD27UVWOhgd968NOVE/wq+yT0uCXxo3wRfJI33Xpp7ukVbxNqGGVdSK8hhCtE5t
3mSje3cNoPNpnXvQT9Fc30ON+W8dCMV8/HLPm6blrhgsDlwjiS65HENpXkFBoH1f8+IsKuuz1/qB
jE6M6bXI8QEpJ5k/c5n03LJUuREuzU+Crm+Z+DZjmpqfO+3D7+Ng6Zc27OaU9xf7IjTMKf/JHHU7
R0zZWGwAnvCckZDabZGV1vgC6XtyzHVbGDAImu+X1eShiyXBIpEj0gaDsiBrAk+ifDzg8XZngrlm
DoqBKXsc+uHOw/4XmNySzxVHdN98bIcukjOVzp2wP8nxdkNUb7q5jUr83mE3f+zF7m6ysuUv9qrs
e2sHq2x3oBtyAsXwMwuBLN5XSfICcyAMuIzvO6b5VFuA7fVvW6S0b6GVkVvgJ5WDsC8TOpK2KCwU
z0NNK0PxnmN+ueFNh0GUCqN8JqtaAoZxq4+6pRAhZAZJTlJG0AIsO1Od6CKNguHw2PMMQizwxdbC
X6ro5fFlobqUitOJsTJDQOfNDOqmLE3+UakhHSrkHyVaNA+AI4E0ks96RqTKUUS80+1njcfnaZR9
fjAyo0wYExjXEoM1PdE9iFzNbpEAHbTjlBG4DrGsy511ZQA/X+ZbN2367OOxqCFx4PXPsZw0YvaD
NMvLlb9UgginMOtoVX70+kcmuRQzFa0ClI5YjfhgGjlbVt6m+jTv/DrALW+Qfj1MAx2EPGV8BVbH
IluA7Gu4amdKruYmvvrJXYULsidHUcBBP1zZA6RhSA56qyY0syXToD0Fy97r+bIYFKMjCfILGMC1
0BH3EdkMJQ1F565H+NDsbpJGZ+IIVkVx69s5mOkrH6xzDruOS3qcnSy3FcsYZgsxcvxjcGmKhPYg
saZGID/54+9GEqyMz5/uFOLgO372zqaDh1gNoNozRT2absuAA0ApE6lDqYJ1xGOW/CdAJEltKQKJ
ktRLpZljS7cVZPQjjXX7dZF3jf7DzaImwZePPonxGevGbhKIX9QEmFOUuL1oLeI5NgmUNkP5CUVM
UxX+xiVt9cHhGwRo0G9BdulIdeqcp0mTRic8LZ2wlXJy2I4V4YymXAui4ChzK7GHR+u9QdtBMMLl
6iVONDpTjSzP/PCr+vhgPrj1QREp8kQTK99HtZBPIjlW3+la79xuVIjmdyIsZpDbgwqX4pIpMrw/
/IJOUmneDSYc1/SsCeYWEmNpht8dEfoGi669w2NxJtyAY1cChuXygY/VENTMZpwjaPToZKaDxtV+
P4S1uyVmLmPUuT0+iccQFUURBxUI+lU97e2emtq/iChF2G1P8CpTA424NJP8ceOfVmUqj7te1Kwu
0ARvb9jajOZ6o+W838Mi0cl4i5DLHccaSK1aoSAKe2IGNI/SWXq6lp5nu4OcoD60ApNDyTkKrK5b
VnGZcVOUVE3TqWkOaZ31dfn4w4ioE1YeB7qlLQXyJCUAbwyuTexLHStgUBXKaYm8F1KjEgVixyVz
HYdF5i4HjUzJXzZT0VV3R3AqxuHc5VOG5J3ciFDwh2JZDzo19H8QqxXYaX9wODM5VwXs7f7Yk7+3
5F27SwGh4ClMoN5SaTGlMj1d2/Uq3bEgeQWN7a2ECLb2/3bYMRJXD8LWL5nyUm93W/sYk2VtYcCY
jq3H1FwOO8cs34U5PvPslsr8EmR39AGTMiqHmJ6hNWH0J0D+iBR19654MtL+QT2hfIDPeAVgkDyO
WPfLKKIwHi05ny9SN9NZLw4qPA8oS/+matU2lMruSNYuX+muX+/q66V1jHSGsDlSuWVVVCrfZ+1K
sdjZfslTzi8gs8JjIqr9KN7FNrkHcbHLc2+ptNDhy4pTD63K29MpR0A37ALH8ykhbJ+OVm+RGesU
NaAig2sN+U/lhpNwHANGiOftBOva/p+rnFISL39O3lyC5jzDf9aVxhRry9JPWlDWJunPWPNaN0lz
kxlbO0KAycHK32SsPrqEli/mI5m/GcQH0Z4V27GRwpZlNZbY0Bbb0iu3w3rX5MDRd4xMgQSpSHt7
uXi2NaUnmkepXgQKzbYV82Gm2Zxh0/peugwR/yKxYruKrbKf2TtcfgzURnxJAycMnCYLjRQ5qCw/
FGflG2n22H6I4TfUNCFoxUoiLyocdI0XyW535haVevGLO13Z/7EM1c8UKCElIMPKdq+YrRidqahE
xNrdrtxFWLyzht9ZP/ZNDTD10e+xsmpH1Yjdt5JqhUyAt+sEj0KfplefeZZlNW3suNrfjDezTv1u
6sXERsEnb7KJds9YlhDlzzK1XfQFt9cGHtWMzJxaBAc/BkepfxWm8dCeYv221ftbnNN1fEcXlvq+
3EPFmisT9MWFHziIXNlz9vCEygSHFM1YZaLRTMCGIasZhIAogeTGiqx6x69lOv7s46TLNeNTgEFC
ak8SR5BnSq+qiqZSr5oIFygeSBETV/jCwWIH3lsPjE11tvcce7k6eqnXvN75Z7I0CcAroAt7852k
lxfSYIjpPJyVACz7nYfesUB1QimO+vXeYwMJqAk952YX8e0CMFrA57ItKiCA7QOIUp5rPvYp7Yz5
WIqWeIBM+efRqO066xZaUTz1sKG/1ZNMKdB1h1y6/DfSEMOf2htzap0+h0a+pO1CO29Rg/SlVn8w
ONhLdz5OQftvTk6O2tpoRhaD2Bg+QO9VhnIlfPNMrFVPjS3N/3R00d1L0SSuuamKjdO5zE+VspiY
TlbrkOUStkm8lyF1NGKPtN36i/ZS0frsQ/fRQTzqq5gvBNzEo+NdwKEetczdsY8x54OW79OojYjW
me5TAncaNsPYQ+Mefc2FYm7n4eQuNQdPvU4oVhrp/KqRofe5kU+i8lfw85INtmZdzTAwspPkU6DA
Ma31UueVrnC5fEIkjsnwJXANxkMkuKNag/mQVm6ob+6nnhW6TAUdCnrE/ghFHJCCIcOz4HrFnxT5
c4+PmvzJRADWbKcchDCVaJNLCYgUox36jR4pZhFMiuOaO1eXWaTGdGkeSF/tKaMRN9MzGwvIuo/h
LsF3uhVy3ZDjSrXQl2pQ5nedHWXtVw2UncL2qGXxdVCbVsrlqwyOaRA+TTwBv0L2MAl8chFEXTE2
2XIRDv1ECEkEpR9gVoRq3idRnAtgbxsig7KSoKqSxkj5xaBYwflLQbWXMrpn+fsSoIfJ71XjxxWo
IoAYSD6XBLiXk93FmafbXbmjsIyYziEfnVa5a03aoKQmwMBndS+H26cZb5V200vpSgQAsIfMO/mN
3v4dRk+AygYWkUP4t2t17Nc+X+WUm43tqptgmu4Q93JXt4oGwUr30tP3QoT3UO7bBdDwAWXnfmhw
svaATqumQYKvJs7bGTzI68sKamzmaPT3Xsv7ikqzbxpK6nIAcR4ukekbXlAIH66YXxnz+jR+d5so
xl7sFktfh/eJIG5vCubiWMEO3I2He8Qt52eHEeH8VnVr89SF13Jywv3HJ+h0Ps+j1HQY4+i5XlSS
pymDd1ryjAD6LBOzW1u0rFIf4KEdMuLtvg2v8ben+xnQDwuzBwv7nlx2+CUcGN/AA/SB2z9b1URb
GHHwW+BGH0xh/hvaPTbYvpy0Tj+t786ygtvivUCpiZ3vG/VULulvSFxv/DnCvUcZ0ZYe9KT7UddM
fQUO0c8pK5/vIZSP8vf+bpr2rLFM8gces8vlH8B4sLWqUrVZQ8Xx4Nh9jfCNDNSmn3vvww2kX9OX
7mdOsvaO65vo9XIjy1KskXY/M8ADLZbJdE50fOZ2AP8otLwXDsYTFMAuk1dVVkXPNRL/WLCgRQxy
RL8hs/1LiylqbYj8v+yurBp00U1YHdaBAtUUGEpeWETFvWVEVNuua4JZrhHAaGjbIj5pE1TtGk+3
5w5XCklQ6EScbTlpQaSDh9f057vFeOZVvLB2/0bd/LhttXJ4MIubcav/w023+eE+j3VGHYVIT4IK
jIVMhCkZ4xR0SmpgVaX+VhQGtsxYJfa+UbY36SY3TG5oa/IKCNxGZ0M8voVqi7P6SwIY8HCWZUS+
VC+JQNmLOmnEPZ7XIO92F7JE/RtQIibuCerqq+Z7HdvSoT5T8x/FeyzFqEb0ff4A+M+GRIIS59ZU
/93U1J5TJ6RahXlafKMVv78ncDaa/3BkI4Zy4Ec1VvDqgyKTDqjdpe7x1E2wS11K13Qlul7UtDBg
XUbXhEyxwTU2FCJR2JMTwWFyXHpSVNMALGg6eDPeA9AGi5TIGK1l1doc9HFX9qN2d2JdIqyCItxM
QJ1KSVlBWsZ4xA+SQ1T4eWsmoXMvs7zv6OB+s0YosC7J89we/qbMQ3bvvZZTJtOEiiOawmAj+jHX
OaLoWjJ2TaZM1dJzYUOmEgHns0z01F1kchtvo4G7nhoJ28rBhEJvXZCRaFd5OxLIKsJN0lKlUPHy
+w1bTqR/Xi1n7b04RifnzAiuSn685GfvvLLd4XmZaLVJyGrY4n6ZdlnSVJMuJeiHNmj+p/wszNEQ
ZPxLtK6Ow5JW5jdB3k5AhlInM3YpnudmiJJVX/RPuUiDhMhfmmq8fs1mBA22X0W+Dc8Qe39eDJZI
pvxrLb2NhUwk5pe/C68mRE931dLzRftdtfXAMCOODvgO/cseP/k1GQObeXZhBPONRDhMCQMU4rRD
H5kNcZQbHsssuX9oeAk2dXgBN4kqfbhaAbYs3n6UxhCSctkEAsgC9jl4asT47rficcGLKWTrHRSn
ZGsJEtNiFJHaC0hFqxtRp7mTPV3i7wri3Trn6HeiyLQrE0AL5VLBbJngXAinN0N0n+61ztkx0Jvx
56Pmpj1DR7DZ4wA16f0xPpz+2RY8asM9P4dj3iDM23BvJcv8gxA3p8DRTMpw+79bUFZgSCC8KMw9
Im3bLdVZbZQYX8bCvlmxA/XWPL2Nzc4pY9hs2UVbQuNbScjDNTep6mpkeKbSk7uGr/HOPe74OWWY
TXmVuPZdkdOEALRJampq16aZiIVsKLmnqnvuqxgMACcX8L0sRoZfYgqVTGN6OpV+1nOhhloQilLV
7Lpf8JYD2yxqwjOYar/Rvd52EFKpbow7BjhphJ2rkB5bZmUR8MtzBfhaiI0KcLtE/5TB0RNBhFjq
D4pgO4PM1D+p12IvSjmznNQw4g4+sac6y1ImSmF2LFb1pu84+Y+QfkY1TlocMYkYY7pSjTk3oUzG
DJsZeZHMHrnNlwqX7xTnnMQ+Z/Fepjpv6B2bwkJmgrOnvJTwD/MdpESXmb9Wa/Ujhl8vESOappll
a2jtKP6Eur7r8/5A8si62beCfZSt67va4RJpjhtzINDqD63kmiWYf6i/ntSdOPwns6hC5ymF3M2g
dAQASriCvQlBwbvkJEhFhQK7nqCYdUoIblRJJg/esBIVqfxI8QdMm9BStbvw11LJC/0SyLhZYFJI
lENAyTjGEXLRRjpV5L/PewR6Q2mk95v1PfvFXh2VYWP9GL4beZeQGwxagiDSMkEJ5RrmYLk+f0+Y
euY/7hoBuhohKIiqEpzfYslIoSfoh6GhPX9Av0iG/wt/HKWI6RQJdm/3XMX57kIu5REDEtIFtAsa
okEQWAnKr8dZrNumpUdRFa+Dv0XKIJ6oVBy7qyLU//jp5GDkNlb+2bNVYgO+eZ24Az6KN/w/rItI
tpL0T9Lxf2xVfqpbxIDQM0AcGM+PBSUGbGeA805YOT/UO4KMVak0w9vJIJVDuLhZgzux6G+PfnUc
q6MxRBi6jO0SEyB9dxLla6cMzqaP8+hFmQO4e+YrNJto0E764JzOzDB1DnSsXqsBSR9CWOPEFkEe
IcGkPPlsWHhRoBDNRjr9NlLV43Wb31/sQUy/j+Hz8mG/RWyzJ5tmuJubX5SNp8qGTg2Fet4MXHYm
PHBCHXfMcRWcpghfmeo2ZBV85oTts5E6hAa+66EcNAz37BBNz7w+dk6IQk/f0dsn7i27g3100vUO
qgP+KsuRVoZe7O50sjRWsleE9St0/40JKIQiGL4sK/BnF045OGg0xX6aPS11QWkXVy/McoTPwK1d
Ei4jtCYM4sU9Z6o9Cr68K28LaQ7hVMleuQtDvyhzvDXwUY8TJ3Lsv0M5iOfr6u+2oW9Lrx+Lgu+L
jmuLoppqcZg9HmyglS0/b71R9C55IHkX6CQN11k9RD2sOIEIyWo3+49MhBY1dmXsp79ahKTjtdpq
M9jDeMsYcPB60ZDQ6JeUG/S+i9HOgh53T8P9F7Ol0LED8IXXcO0s/JC5FrqPR5qi0zoP+xa7QFo8
LtJT9jRlZcl6INflb0RBTvMzQorKMI34B0ElMLOoFgMb962DfS4RbZ4j0OuGrAih4aYluIX9/qRw
li2FQCfb0KJ/IvijFQIwxdvn8sw3LCmPZyz+n2R4Fmy6KjiFNwXnnwH5aFJaG/hBRKW+jLthg/M8
Q57WAhgysX9hjmvG2kUJLKjZ9yZXqxaPsiRA57SqXt0nJwivJnTntU4u7llEDMMoYT4pQRzCQFj9
nyTp2a3/Yxeuz8tUDUKdRjdza7/RWydyiC2VRqMm5PhscU/VAVkbiq7C4s1CyfHfdbZaBKpaNjzz
AyGGxA4qyixaCg4XzfFbZ77+ABSrA8R5JjvJZ93LkGxX5gOvliAZHOlNS36uXqaaAq/0WBjtgASP
rpJuHIBPfk633gx9y+ve+2WZn9XBuG+1BdR+gu9TdwD1Z2huOhBJYGkc3XnKsBsSyReWeaZpMm1c
wE1Fi54IZOngmOWP0DQQaOyOfF/2R8F1lL2zxP3CqOwtr6S4rlpn2wEhInKc7lJNXa1yJ1iBpPVk
HvN7Dk7sOF1MGS+nbjhDGN/nNnrgiIh0/PCDnDbh0y4IugudmfVpeK1Y/0S0Hy2C5sIO7Mzns+Sd
0q3Y3tHYFPurLePU5j1qk180DSJW4985+M3mtSRrkWlFvJ21dBtIfeY7EiZZKSNgLZ3ad+Dd43CG
eH85YOb2xGi73qzWdEAjxC0dgG5HDQFBzqwOUPrQTiEKHXuG6wHO3SUwjrGMtUdIQEA0UN4a7SnJ
ed95gGIijMWMID1pMRXCLYFPpiXf00mnqixQlp+eyHTXtAAB2mEn9jvyKGRdZMUrXS4OILq0pM0z
EH9Ng/wHDqnXc7AfJl5DXMZPAlZYAmMJGjKBRVLyCg+KEDzytGPFDF6RCHv1y6717LqNYcDiHb5P
qpFWv3gDi1OjnmGVWHRgg31uesw14qn/qNF6Npr827+xRAx5MSBqkiXw7WPRKTIa1qUh9f82wxdT
PrUBG2pYHDFFKiG6n6XzlzP7UZP2VXZx00I7seLo4H1QmhGxvzy+VkV9IJlrTRzpmuDeSSdiP4N2
qfJQswsih3zCchmfAFudV+imh9+wt0YWbcIPE+B0yLSiRHNRDL/g4vaqrYQtBnlOLt5AmbUT+68f
s3lw7JtOnumeloIvaWodn1ggZ1AVscIjvPyNkdjG0WdP8AhKYiHlLzyXWZbvpnmfwufLR9TmQ0Je
j3seo/J3L73ZftuI1RXFM0Yt1PFutQLXWfX2ZIyvNf/F4q7lpbA2sfLPeD9pmefXvpUhhXChJumd
cWsOxW4fMGeuZbD5vyGNNkuags3c1Fa0SqPIZgLSmECb/Kl4TX9FA3Uz7hmMGjiWv3LNEfFwJk1j
J3AdpiRIrs0248QQLYDvKj8+c7sNhepNH+VYInh30KUtUWyO7axv+wtXTPf+Gcuzj91BUmu0g+4M
o33LR6b+Z3E4m0AG0dwVMoX9s61gzxInVr5YOwZyDAHVynaqJkDdydOpgSGEB2dEbNWO8pr7UrVa
vlt7VmvNsK/3Y2yGfiQTWN9PeJNKdBuj6cZm4XQ6j5Yq6uG1h0N7lWKah2d2bWqgVjfU93zgdf98
rY7d6nd/EkvvhAInpaoDxRW6Y57Zou3qOLnmefUYYu3dEzJixNSZc0js984pH9lQ6FkZuXa5logi
UIZdZAEoZbJph+TvwsoKmzpNa96rDQ1AR20JTpAMb0vK1jgFy1gvABeowLQEl1yYFwVDoq2OEuHS
oAHZhExB9/LP+YwlTUDTdwi7h90TPgErCviMxQON/Xl1Uaelv+UYuTe6aZqZXpMd1o451lWnpGvt
+yZd0nZoqZP9X6+hXlzI3qcar9PnOzz14hhI03k/vWHSgFOKBaKYXCUU4O6HmkZy2CL56zVgsl6V
GBBiyrJRXYcC+/auImEJWLKbI1xgUTff0luf+l4p42pBnn/X63dyy7QUTCKxpxL5zHMRZEL5+9mi
33UX+Ql0U8NZHYbJee+MqktKhDz12o5BlXBQILuL/2WGR2S5mGsEv4YpYK0i79sTuYoFrkS+YTci
Ggbf7XCYJRnwNaBoZL5iwg2eTsT+2Wpr/KEJN47VIUQ7L5OddSSt5VGaYvsvdJ+vc2qjtP2hRUUc
OqE8Acm4SutDf/1WN6bxcK1JG0rM13ujYkhPCAQWt/7Ee2qMoR21ub+bFPmnen4lNnGFpEcSJnhO
Dv66c06uV7gqp5Dm1FqQVkEYDIVVrDKxyNu+s8O7hXaDwxsrouxA8pCW4NU96SINkxYEEbIqRmlH
ixJZw88EcA+tjz/LERTDlIItIlTDMDAel306PBjtX43axyqsC2N+5Z6Kr9WPLV87Y6VKI2Fc3FjN
nSNPlHBJwIpimXNSuHfv4boBMSUXYzN77TMlJQ17eQF9TW6LbX5GJL1GmRwQNKZiaHs5F2Xh3fs4
8iEFy4DRoo4z1ho4OtQupix+laDYosAI4+85KARmkatVLVHYsW2Hbo6ivjhbA5AoF8jyMU541d2H
5ob+GHpbabzUBG/al+YOavVZsE7T4zBVLFJfeaa0KyyTy46vDvS92hR2cUG7orCbwiNft/ziiG6k
Z0DQBjFYVTdpuCdU7e8vmpDgPA68QLt7ZWatmfeiv6jNOtYaq8X9KQOfgT/Q3GBtIA0qyK2LNAPo
wB6mHqUuf+Li7BH+Qfjgdf2P6lacWF8lkoGNntL53yrYTnSpHoRTCgViprqRJqCiB7hzcpR4ioo/
vH+TsZc3OZ72IquFupOa4Z+/yuo2lL34lGK9a9Od1d2UJjmpu+1GQyjrbDm9gapvg5erw1lYfU+v
RTzOl+27OQnlmTqGw4nUnx2nb2whii7qcaxrvB0ZzAxdNwRZXQOsWIQjWhWLDGJqY5yK/0P6A0Gs
zm9yCLhEFjG3vmGZGTYV4qrCiEMPhIYIV3fChKbf/stToqHbqXL6uuO+Fo0tppHXyDI5xd7lWfoA
WgywItDWEUETkk+/9V2Xt14vAwDvK9AtDqiS5Oe/je20Ib+jbeNCpKO/ZK1C34XIL30MJUlGmZ4o
DO9MC/kscXZKgzNe0ygaldA+HSVfOngR0argf39LHMgGeaquMnwvdyzli7tMmK1HLDGZwLl+eCXp
x6EfORQ9WDJlj2nX4SB8GGrroFoDC3YMLwlQF5lf/Q6qcGJWsRz7Fp43y6MSKVVLVLnAz9/G0TEG
7HzhKBuow7shMK+yP0rQWGnkGPL87sMqK4BaDWrROaaHp8MNIBhH29c4HetkoZhvOfOEYy02krD6
ApBQGu1LYfmZEH4LWR3ar/WuQh7Cqc9GukLroUyZrg+8unQ9MaHLDsetq+0qmIg5KM3U25sIywu1
Fu4zSuCM/oAdKZt0ZeYXkY7i69lvHOfdKI6/prKpxIOMjgghXG2u1Mp4XJGgOwZcBaUxrdkyPqDJ
Mxx5TJYz+otKpPHFH1nQ49qmrfJTyqkOGBGB+te5aTtO9BtmYIngrsjI04SIvf2ZDZHe5SUw23cT
H/2t3AJR3L3InQkV9AXAkTiCEoJfGfiIquSQ1nNO+K3fDoqNgKza+ee3+0kbGn7Mofzq339lPTOO
f1c+LLWxmxQAFvL2ad4GpO82asefQ/Y/LJ9o8DXKI6uvffQGBXXVM1Qss+8A83f7PwNromBLKEix
4d9Mn0BgPFPnMkyW9SGCv5uSAzPUWPgv3n/tgVQFLQi/mKjEyE60C8bekfygtJQt7YNP3ecwkkM4
PSuTCooo74O5TatZos5Tm8Lx0qKAbYZJHVuWi4m791Z0atBx984hGiXVIvzrXDcIkxywmWBWDxBH
x4XnSXNwtThPapcboxV9JV3YWzdFukPEsY69Rc0OvUoJkAq8xQEkg7ExcG5druEz6yZubBjDk/nJ
KTXLzppxrrEFSpRl8tanbznbHAnpUsJ+9XoPeF4eMTK7+frFyO4ln/X1iy3KYAhgJXmXXXIcz4T3
4EIOtef64QvQrpnB08/880ueN0CeQBuzgLd4JAEV8D8UDlEQBQP0Wlf8Jjr8qKG+vRSdYYWq9HmQ
URhQqWm/PyktSEdogQKHVutbKPQbOUPqvOvlNF8zp76JqCaD7Dk6SaYz1Wi8onNxp2T6O0UAtpo0
ocMnlV3yFdaCrU9r2D9+DCITFTx2jxlR/fdhUV7JBCWiYEXHx6867Dva+IJ8RF/ewtwbrLMcmZ+5
CAnVV+nV5WLXuV8ur6zHPAUpYvLjTUJncxlMemaKKw/WHriy9yHxWMuB07+hcqurcGH/gNa5fEB3
Ug9SC6E1hmKaKTh20OGMIQiFCpHig46TavIiI9GZ8ADSH9GHfdnTsXVQPDNYLPjmZoDcZdkOQa/l
AYNuwZOUG6r6QBj4gx4wWhRggqom4jNTMPpG7uRcs429zf9ombQkSsj7tGn4Uwup+SrbcnEzXryj
razujDgcluc9uddLndErpnLWNvXYsyP9sC2z/NCQb8fomUokrnqSm1gkwLUPDNHXNqQo5EWPcyo7
orqUL9Lo2xjeIWKwHnd6KSxGiB2TNok6Jj8YZ2nUF24hyblbF4yHq9LmXLy28GxcyQy1GhUoO+Ec
R4hctIPl6OFeQBJjbTwUVX9gMiJXX4ylcqw2ZsRWbXHm7aNaREQ3ZrFD6hvhhdoje7P3cayWvuZ9
8KWPCL8aHlADQzrFvdBcirTPZUITtZY3blyeCjr7ZXJcnHgCRPafVAGgoAA2GD8LRTy4wztNy/9/
/2gop4xORbaDF2pbzY6pCIHFOOLQ2g81Vz06kBMbm97oTD4oQnP4RMDJmyh2H0xBj+CMzoq5ajbR
aET+87A9lu2lADmT1QaDKHlpDPtJYSXX0sXvkkGrp4zjps63m4zYhOBY41gNJ9BiHR5dqbDx9pUL
neADLsYLiblw1xuqKjM1qLtKC/MkB6nJOl/WhsdRd1EHKA0XXfnVAcrr8EXmB1rFSeMXBxslivrV
Sd18W4BqrZyz5YWSwvgqVIq8+jd5izlaOyqPKDZ3fhrGG7CHg6tyxR5qljMQPMCOjVrJ3gsK4Eb8
ntoKRy4bX3VRKCanYTJ1XMeeywwFwHf+zn3ADTYxBFlAp8PGjEoimmsGClXIpJpa2YSFYSxRlHF/
MHyUX6VsxOUzAM1O9tC0X1tFCNnjrdJEVT5xUyelt3w84s7pwe3CqJxtDWydrCEs3DEMGbZbGKS1
tIVZYI2oT358V7Cjml86vOtDC5uP5eN1FnSURuR1aZPFxwDHFnW4khRzMNleGi9ASfOFl5zQ/tmQ
9VBiMzt9bqTBoxFtq9uu9PUqtyaAZgKRCTstzt7RoTn1XouEIpRRUDFau1/umQmWpZrOH54ARmkk
pQkL5u15iQ2/dy9JU0l5cxl9KQJNP3fs8rpxYI8mc08unUwx58zXiMDDWfGV50IyiHO6GyZJH2Jl
Q5rL5S7vOYV4ltrPKS/HZXAtvVuGw4z/qS9/aL+MHtwMrIzcougcHl5UnFeeI9Xcl2sH1b8PXSD4
gRp3z/TNItAhfxe/tKfLZ+cQuu6zNhcjwan5/vS5+BdeFz4rTBf1uXPX8NMyfdVbGzjV5k8dhhfg
KfhmEqIMnGUnC/RXUGviyrqG3/B8m6hveLLmv+dXkpFtr3UxOrKbCpAOpYDUJAXu/d28wmvvj/Ta
SGZzvWBNiAGkZnoWgKyyX0wOj2fame2bFJ07Zx+MVneOPpV87W6MA5TFVfdPEqyuoHQ2BkeIzBbz
O/Hn9+gdX845A1MaXryQl0quqQU4kfnSpn8aGpra6Zbbs8ZpW8NuKBFuuks1xabm13yePsOg6108
PeufFdxboEteHHYcWgbqjJ+9sfMFt5IvIsElQfQ+/sCorYUKYijWNMwuD0ZsYoSpsxf6Yl7h4c4E
81zjdQahDIJUIO31CXoFGesTCx+6+7LatHcYAaFeC13q4LFuSE8MU7iXPekS/UY9BxS5/LKLDOG7
xX9aSykqX7/RSSths3JwoFX87QhtQWKR93YKYVyjrR1Yexz/scZpfhP8o0MCgi8Ac9nREVBGp54x
PQ2umZKFeul+8dRgDp/7Br0FjVZQqk4AVrjheYUUrFUT2Y6iKYIgZ9t78tHiZhwFrItOdAOjmdug
wOD+eT4PkEOuhKlx+KcYVby3Gor6v2IuMVOW5smmObhlGqD24m96QoZjUj0DdWzoBBWTZTpAOoU/
+r/RNGQ9mZb9tKHcpaAAMbKT1Knm3jmolA6LiUHlI+umwY3YrosvGRw8wMTlJ3YuntTI2QABrV5s
t4g9hnTjbjaAFVSCh5wNXnyUvO6ET4nKrl9FEYjm3Pqj4496teXtTkZeGxYLzjlD19CPwzp/KW6O
MKnkoKRFZGpTdVwBp+5Va3paNIAnvArFMQUbrA1jKWm4KuRPIc+rc9dldwT/+10frV6uub2psZ2X
QEr8x8FfEgqNt/kiDi4kI/63lFdkOzZxtmkLXAB/Ql4+HEcdzRDWT7eTLPKS8Wtn09M2WLCglEbI
4XJVRsypGBzvA7vEKHns1kf+8TO4OqMWx6olsGTj/yad15MHRDFJAx2KNvty+ScjRfUVSMVFamxL
DgM50JmrrmIYcRGjcbOFDw/nvI26Pbr3raW3sgVscQN4ofzIiypguksYNbRDN8k7r1Cje6qgbxaM
8dqbKVXTDgjc/4xYjCS0PyM623lh38GDbyZlsBBF/8WOqYMyTprlxCYsauKW2+teqtWpWqHEhgWw
lvDJc7pFcxp3Q9ct1V+0n9pGl3P5vkSwSwSPpMpT2Xo+Xzf//4+OJiHx4NmysY0tz2QUgFc67DXx
SuBQnXJsUrg6bohrJMT7BpUoMVUG/z2pTT4o4ExbM052pODUQOzvumaFDnHRrebA3YOJTMULtEzF
U7vtIX36ZMpx4nw3Yk25/nG/jm8Z1qskDzNcqQ8RLjg8g+SuLz1CKekwhctUn3HiHLwXcjLipAjO
ZPwTRZJ/Ij3LjABpUPQ0hi8F0jgQzMeFxIjIfsITvwnM0WpcqhPLCWxXJ6/UfuHDbtteH8gVqX2t
pjgrsXVnVBcSh6Ymleu5iRFxs5q//GxqG62CLNS8C7JrQNgSCyUXzfxY6OduR5okradZAhSpAeQ/
0f88ewsmWXMQjr2vtTU1N/EsmfswpxjhrqdWBEeC2gpj8bsPp8eYJc9Lv0CkbSbR30/2UVm6dTus
x83NFbCSPiyVfBcthvhs7KwZr1DK/XRUGDujOeWrumC6S9YX0HS13rH3X95Er4cq5Rh782A87S3C
LvMd54NsujKZHoWjVCw/mFcId1nU8wKvcvWRTeUSmPw1AJvs7k2XY1+tTK/BxWKPjiFE2I6WiEVi
qH61Qcc00DfZpLMbhXDrY65BfqZU6fMJhwuA4fWREmyEzhnBsd1lmZTL+fP+MpDVPszqUzRrngJ0
lQr2CfuyL4Xb3Q9gsjavGduV8mlSnRrQpgB0YFHwaEMvVQ+CvFUPYAUmFP6PlGTTTeLraMXOyWpb
N55yeLN9c3/2G3M/3UAAp9Cv6+cSqZf5BpJnyue+Iobc2DNoVgVMGJuDYN+F/QZvLdwMbbO/J5Z9
WQGRC7Dqmr9zVH8HK+DPFW+YIABSmqnHjCo71QLsxmVo/oxXNYGmrhLCIl/2GD2eOXVIrHS+ZYoO
o3HuRCEEKBueXlffB+YKGKeE90NnfdQ/s47hHJ3QJWyI/3lRjLSOsaYrOV3Ci+JuZwWp7aLLapgl
gqjuexnrLLUoxvC0RXRIRPr7HgTdHnXdUwZTuhf2bgD1h9GYR0S+9M23xcevfXiDCt0Jcpvf2+Rg
eyHCjg/qkHdK5nIp/aDtWKyx3DUeyQcaHVSMcYrK1FvT0pIpZjTTWHj+q0TrAVnclMyu8aMw98eP
seHu1RhontpZjjCbHTtPI8+PcAdN7C3sF/LQQerVe+AXfTB/GQPim90U06o+1L+4XuxgIt8Mqoz3
rg5qO/8XWp8EsNfmfGDzKQRp5qXlb238SaBgBB558fXyc3yaTi4TL5USRlsUFxDZLrnC+gyTKVm3
Mhs9DxKI8+Y73fKVb9NF1E5VcfTcXcxsWgOhRyzI9awwrx+UuOAXnfpAgDF3/ZQCChYcLoAnIKmP
JM7O8TQgxb1Tolle/7YTKjsiH6dVG7KxpGvTQE5rljAbGRC7s8+Jm2SOW+Ck9q8wanzsilywevjD
JleyEceTPZFFY0d3QhlKRZhDcE4/Fn540Xvv8lzNMm5h4WTbX8anWxTPEeSqWQkKa4xw5JrP0am5
4Si6Wnm8/Rcz6+bUI1Dy8zDxc8uwuxuKGwiNghnJAapgrk54TcKhiKpvS4s+wY8K023Kal+o92m0
+csTCLREfSRc7drHkI7R9EoLbnzftveZ+/0PUahweH8I5QzOQTOu+XDhcdXsdUmf0O9/iJTJaY5u
FrNhz4Laf240gBao/5m0QooD6D0pGhVi/dgJwQuucCLCEdc28VQ7QSKYsIQ+GeyktKmYHpuZA6Tu
i0jeS7ETc4UhsvTverZwmOVnA0hOu32RMcg2k1a5XjTzz57wLXLVCUlcuFyVJRnxZyeKEPOT+8Yz
o8qQ6Ma0mdlevLk+oMBh3rSUF8p0sOjYc9/gdWcwoSqgC1Jit+0o6/ICq5Ic2ZfwTgmye1NBWWPF
rC+RjwpaySbOBJ/GGx3PrWSRhNbfWqYjZu/nl7WKtrdQ9vfGLAqlVl22pw1O8jYK/TO0zNwGFqB6
DLlMSiXSqVfX6sW5qlYZ6c8CqKVRP833ynm3yj6w+sCLglCoVd9nA5J7vyXJmgLlzY/tnxq2QCCH
p/yqKRNKNw0b69Be5MHIT1XSl4UlOUhP/zU8uIiCzRaSH7SIsZQ2VxdEyU2XPn8H/P2GD4PSLmkR
XQyj6A2mhpwKD+JxCzlLW5V7P9pPssp9CcveHTNZFRfWghZmhiyD3bjN2NpFc9HdNqZfi3Kl3jod
5VYrYL78DQGKPPyLJKfToUCWRf+c/ybnOdqIjhqJIfAzRTxFD7JpRN3LSviv8aA8YYDbmiVyk9yW
a0X/W0PI3yYkzWijZauZTrahqs067ZWGgNfAD2NgWpAgi5CkgU3mTpDbqTBjT4HqErsn8wu8dDF8
8orXpRVKbLXXwGjhCSutqZ8e119TRQRUWw3HrcqifZdFDiHZ3SwSIZde0lec3G+nOsSFPhv5n88c
FLQtNGrsrN6czKwg/VShyDQ83gmEYl0/09l/Pw8Gfw51pYOVbJGtoWYLPvqXcxnRLN77l7pA3dTj
uqfpXoVDMghDKNl8ZDRY+FDiCtzqWzPslWnmmzSTjy5RnIqIIov/CNnz1qYC0y6CkwyCgxn2dInN
ZDRWsU9q1yxTcA+/gIcrmCMeAubZn01cnd2LIo5nb9kGqyf0MArRsYsNBLSwp8Jpwfov4lAxAtVp
gqLlzcFAenvtGmKWF1zaG2kHzwk9bMijT5+iQxQhXCpKGo5sNLok5sEt8CRY23kkuvZUMmS+d36E
h1pM7ori7WI0GQ9CXpBEUWVI9c0aBb4VqcuwlxMmACBDDx4R419d0h2WmixsPzZJ6O2tFGGv0QbW
QGQIzUGff7gvTfSaCmNcA6x9LPATh87/CCATpXgrVoXwY+Tm6ctTbkeKT/cLHvq8iapTWR1JFGql
pjNoYAzCHj+BSwFf1g9qanIhPy4YFzDaLqDKLucHC3LIoI2+pwNZXS3JcnMR+l5xMAKoA7VBXsGL
bbeLHRy0RmxEq488eqAuo/oW4UDs/Nt+PEggt2cw4yurbMzFgQaCP6NG1Y/bxtjRoGD19jsKVU2N
ELikJNJqv8Vu7RFYLf64qMKKfZbJk+29OtPlpr44o5m+z7X8rF+4NLEPqUeYJZ1Hswp8d01lM1al
po53wne7AuKTUDe8asQ4ywQKCm9sm+hqV0DLlY7fDTQqzuNzi6t5pbDO9u3ydOfZa867bQw5GJ+l
zQfAOjTh0Czrj2MP/bpVIZH3SAPK+nnV6HyEM/OjnynMyrn8kwbbpzTTwZMVQQJR8NXrM41goXXe
QUrnptm1B7ESf7muqGAIPTIZVMYHmR0B76SFiy3CSLD6i1JLZvjpEQNr2/SkIrixJHwJIBt1K6vb
0KdCSEARxPtbFbxx+AbM6Q0nl8FcqduSDm1FWh2pG6MxtaOwCUake6jOH8KkD0MdpaNLC9JtzZ3t
jIc+ifDviP6NjYogGxwTcypeCvgX2pGDHovWqAFpA5oGLJ2PpanP5Z6nNl076cvE17i4pGi449an
7LjKrOu0Sy6zMcu4pk2H8g5Sm56Ay5/s9eKciFjKfvdPn4e/GHW1R7QSj87pA5FDJ6TGT8s69BaA
jUBGS6NOGZWHLCvqdOumQsEBcyq9Nsi8aIJp6bjvz4H9hhz3YDAj9cljUIerPSsIs7ZgIrQISx3d
xzL1SI8DjqmY7I9jy/LJbDB0EZXNCFup8Vm6FerqFyhENbuQdbPHGMNbWiW/Vp0pJK3FqaxKK6Sf
uKQPuDbwPph8LnlDA27Ean19gxQJreqyu3bFWlfXVQEq2uwkT8Sl/HN9kg0hSLKH5V0OYSaQgfBl
wTXZjiMwabNnDBBqwNubYRhRtFYkNlBgDAsBoUit9Vnyt8vEF6JqYrhRFPYPQxRCQjY41O7asHwA
NLwyQRMHVVdIhVktBFLS/r4xeqxpgfqvvKWSR27UXaqMaff59LHevFyu2Nr/hP9C88HSsYQSNmXa
HxSqgl65UFxSRyKomuEADGtjB4znHuRzSm/oOhlPs7MZQl2xgfG3FUkAtFHRyDW5Q8bwcX+3Red+
51T1jpvCdfmx7EwviVur2J4Tm3U7l6BBpzapOHXZqvMrFk9M8SoiDBuhi+lcPz6KRvG6avLQWumu
0p5hG+jp0JcYZL+ux/6xWDiJsheo082E5MknYZfCcPfLYFWA8GNMexNIkKelNKxXvfx3Z7XA4GMk
aJ6KTlhcscMYKp2VQWQACTUCvaXhFh41iWi8iTKo/JCg3NGBmf5kZwlLe9tbrvlGzjj1uXLrkTjA
xOAdNFJFXDw7kz9fy49FxQBHum3E4eNDLXOlUOXQGXBe+ycDk27Z6bzZ0Y+zOOsPTVYKWUFzjNxM
Mn/vFzb/qrd+l54qRoGubKt1Nv8BrqZVfvqsxxMEHcAlGU0n3ab103k12FJSZ5wyzL7Ymwyn9Axk
2zaUdX4fUvCKC6TtzNXUZKlNMiJsFs7wo3B8yd5/aK0W3dnphQLd2Qzgz5Li/D1pb4Q24bldKS6a
/bTeyNyiKvrmaGTTQWg5CUtrG8dgDiJvhKuyxEIuflYb6tZkQqWq4m9ih2UMRAep0LArKA9eA7c/
PV3ni0BcjkkRhbWmZ+32GsvfGvsa5BmZZ7Owct/kWF28hRD4E1sKzx3FeTzrTY6zNJszlFOPc7Uz
cl1xupyR2bE1h9PtmdY85rs/D3sGXaQzq9ZhG53A0tRIXlT+0gg2pF7Ia1UBp8LjIIeTYwggZxyM
1IDE116cfM8Ymzjws7K4aVS3wUAfiLXQEsrAPcekaH9urT2078NR703rSE3e1K/fgXsA3Uo/2n21
Sn5Ad4BNaXhcty8UrKWoE2fVexGW9UZ82OJntT1LM7NyOPJdYxmpD0w9+z4vMg44z7gY5o3M8Nlg
skiXm0TAgeoD5dLQqKay
`pragma protect end_protected
