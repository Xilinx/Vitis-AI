/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/0pQj++a1unPQwd94rBYLA1yDUvd2Tl55LCehxrlztxCya2TY4TDXQBK
sWti0Jy38JQeejI4UuY1YT2YsGwyJyO7fHtPSldPbLOPBiFMD6IYPxuNSOBNPIRlE5ehH8UZAw6G
p2n7cthTWl3M1N6pFh0tL2y6mmKyNPjz4j1WuR4STGfiP813crR2Vbey3D6qRKhPi/x+hxG2spAC
NitEsszK3/YaN8l0+n26LfFS9XcjALoMLlC9PyVsgu2W14Lr9gfo49jZRH8GwK2QmqtKJV/5GZyH
Y8pigku2Pk5NaVyHyfFIAZCG7X2lsR8cRCuuKHSrr9cqnFJWdNpVgsGH68CI6faLdR08qTyTdXgz
xZokqJXC7OCikMwSrAGXD+aYAbYnVgKZG1eIEwfIHsu0lRXK4eaTQG0pUuMcaxtmRENCK+gyfUF7
jWjF9Eeo6VEnK31Q5/J/sZA+jgpOJ7Fe9Gy6pC2ckkKni8jpYVHiP0PD2VHyJTjAzVPb3DaHoqbu
2sGZgcCf72CnG5UCDPseTZLUGOmwAXtFdaRStadW5ZWUSRUX0PsCjJDDvsoMEs5ybPOOq4jgU1rT
m66QdeSCzk3bQKMt1dVYawMXlWOTcCqRr2oUsAkzso4aHWSG4H1TOVs3UMH3HG4RHnsRYDvBuMIn
R2AldiqhImTXeG+kRCMehbPCaqjmVWGKn9tHlW22KWvEbhf4c0uLezcfA/vA37GFQi7M1P2VyGNj
WilzOf0ZJESIC2hNFqhMhyFGEadLf/9KqNJ9jovyg6mA9UuJ8ARI0siOlj9jp6Dw6rFrZTmfIbHv
7GBQionoDjWD9vaATYvUKCD2Wnh22G2H6yFn1GdCZUBokz+HIdmGApLz2B+lF+WaC02ia3fDaaRE
BoRzBqnvRLba41l7CcpHKpnc9d5kCDU0ymBVNwT8Yw+P6uPx9hEIb9WC67R3o+YHX9nrpa6cuPF4
Tvu3eq81sL9zTFyRMDNqVDwaQGpIrKJSDwmWFN6I3AtbLNLCSKCl28f8Phgqp0vZHVGp0ofM8Psk
pgvDIPbCmpBeqiizNTsl50jcViRJWZXBnzBc24ll1CQW97Dgxr+gcI9/QpI2XO7o0f6lucRvpxzk
21Yq/BD8NzYpwRNlMXOLNspkOMp34LRb4uJ+PBEtza2LLqQalL79ggD7672u2tVTr9hWvVFCxkGr
wPcNsIxY6Spas9WGq23q5VAn6K2OEN8ntEdcXuhwe+KHKI+iTaFU8uqp2Jd8ognNksjVK1kCep95
RHg8pCQ8eTQhA7a95fhfhnJ5vRezGJ7VMULsUp03V4h/ad4D62dl7EFknJkkEC78s5byb30tQcoN
A1azSr1aSIHUze1TWbBvR3arpnaDBLJpRL5sNIsN0/N51xtwrYQ/ub69kJyt6m9GSvcqLdOXqwTn
8PkvjNB/RD4hVXqsL5TBD3NSzhEdGe8e57k7A2TDNZ6YQer7rTpVVW2bYsMZIYysZk8ceynGqrnc
JSMLbpWD5qzQx8C6XY164cU60l1kRpirhywb82ktu232UATx3fZCeKjHEbpHkAueAQGwsrkeqg9/
O6bK1emyr/ay+D0J3ASqqaXAsYS6aWxHQiWUYx0blwzSwbiOZw16lLsCoXPyFIVDsGbRRe7uAP7M
MlVm17TYgnYyROB6qC4CtBe+QrWJWk2p9hjcNS4V03b26jIpbwqCIz9jlMoflIjBflnGztxUxLYq
vFgNv54b/cxsGJC5Y+PYMdDxgp6kJRckNPxvdBnSRnPppGH4G/kLQMjVErHp//lSGzmMLyx73mt0
o8scRrELVa8LJuKYKT0vIBc54BSUfKyJVXs0DO9YTbEw+AYNB1vMRce+BusbQ15Eru6pNF2c0bqk
aimsvi/s64i5c3nxR5qaMsGPzAXDShO/1WLBA99xWDADAzewaEJamo3NmQoNBTfyxMOC+KaaUqQC
em65enze80y2LkGtGHbmPdnKcx5Ace88m6IKxQxRxlcAF8x7JKOTj36eWqnl1+UlbvuzCJ9B95Jw
lxpYtAuee2inx7QuNKD826FWBgkJKmlxbC7D9y2Tx/U9l4tpPsS3X7xHexR7oMgRrXB5VT5N5p09
/oWJf+GFMTrmdLwNAzlSC5sckSMy/r/wv9VI1dO0v42p7hl5EQNxi56w+ZxtMjqdH6VjtdLu25kr
O9Oq+x3YDPeaKNxQuxQFT9zKoqm1V/xZ41VK3/lBXJOgW+4xN+EcXfHlndWsr308yv7P6PbtDo6q
QBcvrO0DEyVfC5TvdtL/lowpz+8LVsw9/kdTD2HmoOy61ecz5xe38PKPAMg1Zg968AF0M3Cy2QQz
MoxoOHejqqugx4wSnpIvC59RKiJjhlkhqmmdzIOEPdiPfSLAhl4rmH23s6Guu8D9RO4Wo1JYA8Ax
3yQU86kEq2hSr3TdzQwE3rDqZvcekPpj3maH+ivooMAJ6rOBAgGHY5ix8LYhGU5WCwMDoX8kYbLK
UUFRYLOpxk4mcz5D2VSDikivmQuTqCs5NMVRc1o7ZuEN393RuqVY7qDlC/ygD/q3C+33G2Zc2UdO
4+RAj5GFI6PN4Hfi878cHLp05nDuHcVPhTPBcAl5E5IDc5YKo0BJLwptEZpKaxRbVVw5vxyhDeX/
dDdfYG2Z/fD8kJxoCUiQnw+ssPA93LjFG4+6Xi1sLG7aZz3JXMDgl2GGhj7jL5q4ryQff63PMW+9
GvXINEQkBtXoBNFHwJza5O08DgEzM8AGM39EVDy/ZmTe6WFbnKO6sKu+tK88KGMkuBai9ptPm6Pt
kR5Prm9ysAFNgUcmzO3pb0S/+fv8BYhcQW1lv4qn+/1nRKLeT3Com5lyBycQbomDB9YbfjBlRfR4
nS7xQsf1FE5YTqeMLUL+xY2te28GEa552gmQCha4UN+r1tNenYfiNwCzSfq6BzI9h7rHHE9HWisk
jf8Tz+XG7myx31xnDsBhxCjOzYiyHBfvxP5Tdrf4tto3yJGMk6+NCEeXXn7fC284qhkSsY82lwJl
VQEI6XFx0VbEue5wG/iJJIby0Pd58fkF/l1uWtcOviX6pn2Co5/rzXEIwNDIyRWhtum/37pBUMr6
JB0DC08fOqDli8cSZ/51XmrbHNRTvJiYug8X0sEnqdC6lHp+6yAvh5jrTfUUIT9DbbasXw4r/1Hg
RKffbSJ/QheAgiNjMpN2JHKEcxs0BGShad3gD3/TV02NDNHqx0y3wBrVLcrgNaxkdtxeENRXTPyz
aQbPT1C3+42fHzAd1W7ll2Wkw3A736SrWUvLTH4CTHuxjiO4ePfkF+859o//LP+ZMgTz6iV031Fg
ldtuNe/P4bE/ITLTXYn7Xu0rvotpuM1Fny7CA4ZTeMNy7AoGSCFQWYRtkLeVpFnx0/Ave88YK3uR
kHveOF5TdlL2s5NjTzpZnhGqD5MdcaM6tCNEUH7ztcEsnJAIbFl7RuHmbFu+O5+UskS+94aQRbzS
Xp+QO+lofoCf1P/VYAJV0UzgHMoBo1xP2RegOPKGbOAv4dJtHSqI3kIz/jni6UdC1TpCexSL4gyL
JZbiVsztIiMCcA8nyQIUPSF9nnFrEJxG9KqeAX3TBdmEEt2TGNVnoJTQ071QevhaoE1C9IjjoeoZ
yNkgx8onNt6BKzE1EioA10V72IZ0Yf7s8kWG/WtqzxdYo8uLRO0Um9uLaC0v35HLfa0T4jxaHUSC
bivytekTc1cO9vnnDghVoN77NQqcqEotsXtlkPLYxbDmvaeUuVMtydApNZT8iNeWm9XktPNfEZlI
4J99bHrb7L2qj7sqkowhgRBEdjTCVE6CcISdGOEjG+JH+ECc4SpAZX0pFqAc74KFfSslrHOGS29o
C04pMpfqd4NAXg7g4vpbhlSEgsa3y0jCDIme1drp27Ya4vefMW1gj67G+Eh55p412/oGynIFbsiv
3uaU70v7OnIEXW2R7YoQZRy1THVNt/morHsh1WS0FkqaozXBwpITZabQRwbuOLxirIUFN9BrJfqF
aJ6DW/4XHwvB17P4O3RatjsHFddKm2CqB4+ubT7Gc8qXP93fdieSgjyI6B/YfUxTkbpAGwgqFJPD
i/PJ6u2LF2wkOyqnbOGUrACvZQEPmZRQGckZMHYbHmLOJkekreqOkrXP9vRIO4ktLpxXYrWJrUal
e/eri+MjMoX/qz/X31NfIAUXrfnffYzevoVZ2lJW3jVyJMZP8sF/rXa6ljgt99lBiqAyTsOKTzLi
t7TcJGAwE5nz4j+YM72SuSfX6vABsiTvNAJSt/crzqLUrkei5AR60lppewmRG+B/gX0GGvHg8xJh
3TRZM/ys3PPvgHUxmCewYI5YBuK1udiguqVwBnh5ol6rPMuBHz1jctM+kAP2uRn5nyan/uNozSrb
7K4yW4T2rUvdKY0vplqHOad380Dg95C2we4xOm4yyDtpoz7q2p6Xa16I+vge3zGeEE32fnDSSvhj
T0Dk1Xl8XYbvZ8f8QkBBb2jCKucBfleftR9fCh+xwJBt1EeCH7EB/9gr0u6IjaUdYa+vuNB55BKk
jSSX7OTYGBzjmqlp1fasiJuzmYSn5INSUeVyub2qGjei0y92rd6ljR/mKhFpJ5qW2MgTdcAbQ/p7
FwLBVYKB/c3HxQhCnaDApyxx/NyhtR/J0pe/wav25bqc+UagyemV1ebhwybXKHeMYXD9Lv4W4K90
sCAcWiVKPgeeVwV0FHGrAm9dSi3g+X4y5bj+f9OmBDAlOIhwf7accYg+HhkyacSfiSqTv9M6yzB3
fWFChDdWHcRhuMDM2Fhi3ZJUilpkPAxEWUt6Ez43EdgHamNssAXL4Md21cqiAB9cuhcGzp48Q5Ox
AXNjQRFjoa4GXSG7RAPGrT2+0Bz50O5bR5ZML2td/gl1X0VOOMflsOgbSK/ZOsf4aveiAhMoVzD+
fSh97DLEm/Oaa2Om1Lgg603HOJH8SrhRrNVFRNeoSv+5wmTHJj9XYQz5LZUQ5i6Q7oq+PTTVOqcm
ES6/WOkjRhtzBn/kQhI4sGYUXscqviJ6wxSBFxIhYdvA7nOV76+sXiVHK+eTJ9i5aoc8z5ONYCu8
ID22hRqi0b7QT3mu8mzkq5ixN92tvrsqdAAGfGzwdkYyg6CwqfPTWqfAyX5TPn/GUbRvUt8ZFSoy
aEcBlntIZ5zjIQ3fd8rj59Q2xaen+5wsoyVCSLt+3zxFywD9CILK1QHLknvmKAja6K/37kaDMH9z
bK6PGieg1MIwbIMRxFISs2bHpqT9EB0I20RHjC1hys5RyfPSnjjtpZtd4wc1jS3ErhDzNHIFxg3Q
+6q3Or8ZsMp0/h6+uipMCqg9vwW3twUzBjirIxQ2nsp1tn/e9v6yDfF0TLgvb1PS3nB/f09w9JC1
afJzY4ieo/GdcP35vvZP9wcl+Jwlz7piUEvC6sTUU4LOwRdWIf/ZhQr5tn69QsE3IKAJr1fIoG8q
DwoROpYKE3KCz0YH+pGzZo2YsOYmHpCBsq06dxqW9dnP8cPvJxSgYQGN28Mvb3U5s4hMx9Gdcc8k
0hFeefU+aKmzFKXxMzM9gHudUUTmM9rHZBhb/WJsS/bhde9uy5NBzZuOlZUOkypB7n/Rlt83/4zp
8u2s00yDh2elUPGr4EkoY617q1AGWMZghZimo9QRkC9y8pd9HjDDgQnTydhGgSvy35Dcv/rT6+Ot
hDhfET5WwBWA8ISst3eamkfu5GxdU3BGdAzHTTTXZMFEu7xVgr5bnmCl5blj5u+DV27mBdsgs1N1
0GIBQs9JdLqzAYSf9xC3Ulw5LCdgQBlwRsFa1U7+sfmA4qlQ68uYnTaiUzFN01aSEk6TUJbpYTMj
siSimlMrLSWGuUiQ9YcwkZWevMz0FZdD+xO+h1hIMiT39jsOjrTSyScL3hJwXVgN7FVk65ltlxtO
TIUYUieg4ndG3JXtOC5YR9dCbTnQo9XPTO0UGQdYzFdmuQh8qgXE5f7uRvKbGHAjB4+C4Z2rSQcD
BQttvVHfhOylFRMeis+UAL+FEHzFh0EdzVIErESAY85xsfhAWZLjxlQx1FQWUwNLfqjOSOUFizMJ
1jqgMdhcw1sOimmLJCDpMA4EP+mVSn5mg3+ZGIL8t6TdPitZHYOB1258wwr1L7D7jiIo3YmTqCdX
hq41ZGIbWYKla0Haycjv87Wrg9ol8HEYh086/BJHCdT5Nw3mfWl95f/WTPRwCfAzZBHYfqJtHsP7
P/OjJB4mL2FtRbz3mPS6IAGRYHOBKuRU9KFEsrckzrwJGo1eBP0LvzdeE0eALq5barlAs+id2r9o
tfnj3Gz5jfYyPXshSH6F7kEHdp4OtzlWwWpgHXx5ni0ftFqtIw0ESoGz8o7QzkdHQB4CExpNhGuI
8vhZIi0i8yzt4vX2gqC5zFok+ZyYX1W4AQsh8ZwsuIiQ4arWf3fZSBXnSLoR710kPnACn/C+42eY
yBj3eFvvMK81XR+9Y6fkox/sCpVK8xEaUR0x+xKx3xakHoQXlUc1bevvFMiyBPuyEg7Ua1ADR6eo
orxmQeYBs8NKOx8B5U2+OUoZebqbPLhQvLETnXUPFdQR0G2PbhSQz6Qhi9hCa9CplabK6avEc1Qc
QdTN3j6sEUUqOjUuvAUsPgFny4MNbjog1YdxVYuIEZVMyvV0RLCZLDj8/2lVo+oFZuvKjgJTXTxY
2foBS22ZNPvgmQK3FHWdr9uqDOfOu5Ru9GQVkZwF/5L2e9HRxEeX4wrCbSh71yJgr7RU3f897QEf
UOQEwDnb09YqrAy8mwRYJVORTgyCTEPzRpOjRvzYDjrldLjdhUhj6emY5ryJFAxyqX8owOgCE5f8
Pz38rJyRi37ZWbAYxJNNGhXpFdZ7CXaMBLWrEcdrtUELaILh1jsIW1wjrVisqAs2rTTq7k322kwT
U59axogi7XsDiAy/n+33F5lpJdMfLoYNI1NcVjAvUAYfMr2a1c6v8zxNdMqLd2lCHG0sJ4Nmz6KA
0+dKPxMi8cDpxt13J9/0wEXH2OK9sqXPLToC4HrjVUXWo0g8EXCbU+yjfRP7yFPbd4wT9BqXzKgx
Oz6OK4KA1F8wEm3mZC7LoN67U20VNHIVCRG75tx4iGP8nQAVPWdIf/3xFs61lJsSUvcaIUPEY8vI
qIu6N6WHRoLaVp3Q59MZNWgNQeyvxdZr+iiTYXRTOjKQgU0sf/szeI8cujLE0Cal7fy5rKnp5Xct
gsN1B9bq7CFfsG7/Qxc+IJoNP47N6Lpr9NVpSo8cjDBSRnKMrVIoSvR/gZeITR3w4PhEkM3V4qYa
LUvmrNoqYL3ZeycgCG3iYxLHE24So0YSRyoV8NIX32nW8uCQCj8Z1TJFGbhSoHGsjkYJXQwKlPUL
02dlROd2hS8vjErA6tcCq+PyIzPTCUpNXQAIUmUPq95F06puv0Dqg26+bXdMHn/KGjRbwAga8C1E
fzSkom2/RsXn1UbUfrqjLBkNjHaRsaU67TzzeYDNGU1shdu32W5XCCCZxuTKfObg8j+pzBkUi5Fw
Kp1ILr4qbPfIO5K2+8PnQeNmKnGwJs0DzEr4pSTm7G/tQ4pnA7F9SaeM/h0z/yfGwG0ORKKWIAqj
4dV9l2q3SlEU4GDY8SdjLrGT7eR9LS0dxLgolg7/ZVh4ck4gq8Hd0C/sBT0tTLDpmJkToxTLC27X
0NoF/pfW082owhz4VzbpOgq88li4tr6LijUgDhY2FCfxTXo8wOpHxeXveqgF6QaaXPgx93qOWh6s
/UBY3T8PbUz9VT1y1xVoA6gk3LUeWPcwBE/5X39b9EYea5Jdkif7CsL3E02hyFVoC8+rRpMpEd2F
2ud4oG+zRh92AwgOh5FFlM3eXASeEH6gHkq/vbi2gWegD6hp+PmaWJa2sbHSh/LRugI4vgWknykm
YFvix1XXgGkhsXKwVRmI2jDKX8+DV8F2aITuEoxSZiwOIU9UgIndtRSav0+6BhJiA6VfFOOsz0Fm
1vMS/fWL+rUD4u3jU2O5ARpfN8ayCoVTN2kQ08gIfBqYdITbGmqM7JHdM4aiPbg7N2ZzHo9n6rWU
tGgPniKb+6JWBNfXXPbfqKjnXlJ716k4aRVdQcHTBtk2OycAnqA9XDXnEHmni90Q/kONg3wxx1Nu
Ep09T2tCFFmSEYLsahRbqezENJeodxJ4vBT9Z/XVdU54pi5rERUTz2GW5aogrWLnrSNdXQyflMEX
VcFY9ZqJQhUhm13QUkue5t9dV+XTbNW1B1m/mNoBG37cbXQI0u2PhgQElosvTErZ8rp/3WQpI26+
O2UMDDY9QZH3peMOcLhbLRur4TR3/kHFwk+xq2zHMqcrJ7qjx5QSk3iIc15Ai+abELv0sXYnrVAG
nqO7zo/Od2X2hSmlpJOO00sqd1gYo2yrcPq+wX2A2DjM0KYEj1B41/NW+CriY8Ft1qH54B4f2/kf
yK/kErK4TbgiMWcI2rU0nZouOx1fr/TGD1XrDmgr1WVb0+Q83McxeI5likeLdvOdj9tSYJvzZ2yu
ZwQBg5sQPpa3kf1t8t43A/aEHPVu/pfJoJPCe9mCscE++zFRk46VOvKzDFeiJHQVaR82yrPwgDyl
YkfQD4QQKpekEva6ZaUm5/IokCZbapaBK0ZZBtdAmec9ZZgRA8XPMjMqr1awrpCxaACfs3sJ0vr7
FwUdfTABO3uX0s2j1zr2nbSUx2vAbr/4NcGCUUrwrPIvwD8+WbiA6H6+7Li2Wf8MJ/P26u17ch6i
om6mbSLqZllH+8UCW5qWgtgJ1WcX4etebLapzF1HT1V1Pm491m8hoUdDRRpozd5m8x5mXASG+g6+
Er36x7gleYjXjtJSjhR4IcfZG7/rHu7ro05AufsKMn6tA3k2F8VzTK8UWjU8NcVTnPr2aJenEtKD
elcfkUggXzTbj5RacVefZXCArtflEng95xu/NWr6yhdFztwSrD79Dc8ENM6LbS53Z8W/ln8DJoN7
HRg/LiyvkGZZ2RuI1tvqSRIrNLrgwnWGBrNgblq5xw+Hv5IWAgX48WgIq/RyWTjOe9pr0yCXM6N6
D/HxssKDWaSHZfmnK+3avJdsQae/p9ixCvnSHqSNymDM/LNhTfHHGyXbnzvPWoQdR6dmTy7wO8QQ
XC8NypbiCKl3S27VtswrEDvJ3Fi3Sz1MH2389qfy0/TcjlJfWLMxV7rHIWg7qoFJy6+84oTES4UR
1SRmEbcwI21U3tgQCJknxcehBeX3Vp+8uBufufCxpEt/K/NRMhPLfg2R23sMIkpwSxGCa6RPIljQ
4V8m53QggzEwB7O44PIbvlEopfmYTJlVbD/PLAl7dWeKNB0Au75eNKpRQMM4I3lW0qoTqfDt3LGu
utr7Kzcg1AHDdfQ1bCqYnXQ3Ut0PzYS8XdxUP/KNNW/peX/xKx7TTXDyAz5qSAL/s0zx3oXUKIys
oTsmO4CS4xM7R2VR/l+2YSfXXmF44ZgG0VgbXMmv55wR8JYnp679WaatW1/JAQ95/DcLkqncKwfq
+weX37PeXQC9vOcZ5erWn6sF1AQwvVPQoNuCabaXfD/7Sp5o65eszanQ0dMiIe6rzhgvEcnox4rP
aMsYTVjT52i74KgEbvPSlL3ZZx84+3uhGOdZ/Cie5DSJg6Cly72fIZ7X6xI8M7lEIN1U9q4lWmDN
k3UK2zDnJtIcy1Sx+us4gRZpV0W/w0PI3TnbDA/aGruBIu3Y80nFJNK/lztlmL6NVn2JE/R/XWKe
mTj+ZY9zFW+8ZPPsBOfq4GfrkjMTBlVV81rtNpu2CKIuWtkCmWgW4pJoIyQA+ehAIQgmgrCUotXL
1Jk5XRZbU4yHleebNt3nhupV36vp9ecZGEIRcWJQfaX1hMtcII7dZhUUZLvtZYRFj53QYSe+T5Zd
LS1ef6tfsg/g1M2N3ExD90kpWAgJiT3BAF9bBBmT9zip9GUgqHqcPlD1wgLBgyyAyciXCdeQ3/Ft
0ASKqfk6kNJfqJNnA+Q+uLiwE0JF9DQYB5j9kI/KfUnCbGlF5eq+SPKhDFc6ZD8XH9ml1/dOb1Wo
XxMRR6LwrV/GJgyKtL1A7kbInKY3rVjz55DOQ6RmSm5QEOrxF0qQhMSjA/U5yP6hMi3ZuxjJM9Oc
hK5tgg1IBCwoQq14NVWxvFcE4/6ZGcPq3cMsWemp/NkliLKBn9KLsltnQJXMIYU4GUzX4+z4HdY3
W3SHDYkDMxQYPHeoZ+5ZRdjNoFGv6wUbz6WU7fLRMGbWTMzhUWB9ktEHHr9YDRi70KntnB10cfc2
ErH+OqI6GUB2YoS0Wqp1ItlNcFNwyrJj5RhNtto/Nd14vb7cRMA3H4qB5Y6cPAQ33jgvz92WUdt4
GrnnrIyfCIz9e5sfFROO5tkQrOI7PaaGirsi6bm+c1Fyw9gzdPwuWR75bHPplbXvkqdK73mPT3Iu
St3uytKnm35V6fZg26zz0ZEaTLmsu978HrfYi9shcHLjqfHTAXJi+ycqzTjWz8EzhZMGIUdOGgVO
U6Rhle4SI7j8Gj8ri+tWPnGC//BUF+v/BNKBoFqzjNQqyMhBwIfC/nylJjA/AlT8gK13HNNbQc47
mUqGq/1YwXrSEtiWVGlDWQrsNQfcVzJ16G11QsaCJvncKCEVbxBz3fCZOLW3bsq87F48rTUpd+0+
V594nWoU/5UwHdu9Qqd9qPEV9otiX3RnlixqINalDnYOxc6c7VMWVD9LgKF1B5rbu8xWIsU4iurK
v1zGMdkOwjQvBbeOZW0LdXpfBeA/7AwU61nzWEEbTAHXytHQAFOngr2+/ENvcYdpH2XJ4ysWDu6W
YnUyuRo/LwiWFrrMRF/x7iYOa0LPwJBdATtu7LHuhDYM0fEOASXAeVvMpS+1vv2VSzdIN5eiWrwy
gNjV+eqavNjA6pU0LBL8PV4ujBNGMgWNBJwRPIVLlBoNsZdA0V+y9c9dw5v/ePy9P0d9c5RXZSZ/
acgGWnHW0SBtWwODkpsmAXRyEO5P5mhMICRs8fQs63xuiRpH60p+JL8WDF3CgE94F8jRsEaMjlN0
rIxCCRxeSenPgk8aS+PJiBiMO9dBwebCO6CKJWLM1FOVj4f/aBWdu5uh6iMlDAXQtmQBaRVElxL6
QXdXEHvncZ/RwUl+U7/s7ySwsXTqMsCrfWNIV1NVq7Blrte+oHNBvZmeNGuz2wWbOg+YBoJnmHOf
10Jhg9Fph0AK+umyerUMSuBFmQYkQjbt+TFqNsbjVR+NtTGxcX3juwA2U1AN+BsnVlq4A6lzWu3k
ZfH70LW+ztAwgz7ZorruFLd7a7CCErnMOxoA5mh/w8YE0FxzIyIYYM+S/CNeFXBbNvvMTcIqvZZU
QdUGzPcg8X2/zN6fwU4iDy3T+IceDhjLzxq9tTDNSbjLnQPV5U79ubbyNcl/TXgp9ibE3DT/slX6
cm7LmZtU7/0Urk3ZoL3imgbSYXERtvPX3i7hMIwQzpTmaJuk+IXxQBA21j2bTIclsk0j+fkCnAxY
xghLWtoSRz9frzhKujIwHCFNPk6qYvctCMIz444hzM15xB/blohQuBNIR4m85x/dZTfrMQZ358+i
IlD4/aTj1ymUq3D77lt3mPR/VNgMAK3CWEZwtUg1Nk7aRJOobOo+5O9x5J9WBdxHKwj0zLHYuKrL
rxY+EYEZymfEtya+CUDi8HzeqkS2K4F7RfL56wDiJWrkWbFmkMmtBvxEqzLIeCOSAzQ1JsgUGHsL
/m4cj/E24dxdP5PyDtydFqya4TBxfUCrMLzpMv6txNz6X2vNrv2QtfptMmLHzPEOjZGrc1T2rBkD
csytqIjZ4tcrh056gObNBWNF3il4VyI8vxtV9fQQz2BQ7j0ncqKUILqVYPBACbWp5xM44dB5H5+2
bOidPkNPs5UnIXe/F/VyazXnuKsJxjVPOMb39xAKWDNy0gyB5Hlp9z+jSjJDWTR5VlbBDUYrvRfs
t/u2ntgoVyv1CkbwupaqJ/DMw3erAAfdXAwqpy5dUWchKbNg3ZUMPmHIeiAcxZ3bSpowTX7J07o7
3foaCi+J+9p2B1hYHQjOmRj7HWnZJyqckpUBp5kFigM+CgcNwvwLXjbM7Zlcr+P3VvmQg7OsUbSO
spN+tM14LTWyVCGEides3m83s0g7/bfIBCNX4fUfozGqAKk2YVLkvyMKxw9QQuBja8Asr1/s4hdr
WP2h63FK5FQI2MM+wLC58OHyKwbTi3lbf6AJ0CwOLQxJ7rJNp8fQ68x81vrH8FVJS+g7Zpyv9qa/
+HNnyj5PxnwdCSQC7P7Q0efsx5sGyAMmD4oBW9ZVMk23Af4l4wM1XMixVbstwSOVZSE/Ck5ybN3F
7rq/fWriakmu/U4zOVcBs1px7m2zFRRMIfn5jgtLZ6VTKysmKSCiFcNYf2o05l2LY5bGnLLhuogt
k2n9dKzCKN1FFcCrKJCF6ZWQ4tKrhH3Pt6P1bC642qa2HjIUXoXfdAdetXNeS8Oh9ktPMp5+39ox
VoQ0tPAOei0bP94MmvUsXII1tRz9M7P7btPtNvnSsy+dY2947luU7NAsUQ2opMX8GwumODruQ+ci
jZi4YRC6WaVrGwtkfxZD9HB7sgYaFIG9ugICdEW6+RP+Ek9QhLhY+TcUXtqr3VU0g1CdB6k41b6N
t1ILRgnKZBRkmYh1q2sfrV5VaVNKf/OcpSF6/M9USh4Sg201xQc+iUSJPRYeFnG08zHD/GnLfsXq
uA4hExyE4mYf6/RNlteW6HHck655312Fv2b5kt4edUfRzZYYrB7/8Ehyk3YHWYxTaebEb2ixhOIP
bR7y0/ndSY3P/v7vRtqsizdraZqjKAcMlu/85R2+zANtmoBVHD3GhC6saQHZTviImA26hREcpY1s
21v9FuaYgQaXJFPNbUWuEtuiyifjFV1ZTOK+qU0/KCkAt1JTGv9z/tGGvSYxwcYjh/ihFh3ma39p
ekh6KEouaJL8hia2VVoBu6yY5I9NpzZ6KS+YDiomYhCxO6JI7drLHHMkGpX+lSoktmrf9EXnidjb
/gVRrEOj4MvpeSKMdpLjDQ9qeJ6DbD80kDecypqLkGSzUEM9VAYRXU+EwD2fJ2uvDTfvCHs7mqWt
dUGsiQVqMnKbq3iIGiFBXbecZGDaEuMFEiisSregnX/Pon/VSUx4nrbOZD6stPbFHEny0P50dgDt
TEhCm/8lW9V4LJAuEuUWlTGgWz7T+AKi9Kkl85Ikiz8UlwYeQqHTW4hqI7j79BY6TLcPYsm5BX8r
N+weJRWRWsPecdYTHf7HdVUlHMiir1Xd6jdkOiv83WIee1pjGwYd01ZdD9Q5Tv5WFLGXe7TV+/LB
32+9XHkSCrPXiENlTksmqlc7GXd5y//k9Lv2TUWeByZgoh1bX9P5FKJcb9LbeCmZHtkN+VLq7hm2
9kMX+OAB0x2BUXFLIdD3XvbnAwgQbLRdc6PB79Wm4gucMWx/aWdjpJ4Hxie7+/NhU91hktNCqdH9
ASBVNbCLJKRUMXnFQr0chNkTeJKIhQQsarncxAw+YKei4eritcR1rAcsp2E83k1vbV2MoXsmtDlw
eMXZYPHCZ1PNa9TSA/fd904ku8V/S0RTCbVbJN0tlUS4+70xP6HdCoYm8L6olOrf/XR3LNiYbKsa
EqzL3UmCYddwoIr0A3YwQv0U+dBMXm7/Vqz1DLnMiZLeNsPzV7fhzXnRe9NItRT/8Y7eo0q+6PSY
f9Q7orXWmbmImiINXYq/opHwY+OUmSzNiDUGe7Q5ZEshNLH1fPD/3AeHonXitB8/odvj3X72dHIA
+WBfv+Mwn//5Iio0seGiDg1s795yas9TRLdAu/ei8NZQYSgMXU3V+bdTmjABzxWLsKDIR59nrWyq
ocdPh9oK/vuqQZE3p90OFYKTYgW3zJra91iXN+P/STPKBiLa9u5UIvsC/ck6lxoc0lzf0ckDQhI7
FSj5Fd79XOzEtFxLRkZsI3Tx88z/vfXbAOzrMFWhnecgoXQjY696Jvrh5I1j44tyASEPduVxXc3i
ViHMfTCY5L7CTUNnLUCVcg89a7OHQ9Na2+0DlrbkC41b3OzpUb3LtY3vPmFiZ04+aI32D6sgQham
cg7uWmAjzn0wJXhDY+BM2pW9eUSRE6daCHnQgxMQ6VfaC5KeFkv+IHYc3yfF7kM/KTF7eueg+CrU
V9vTJGx4WHUbVKefFkr09n3wpzzr2wuvSqTAw2iofcrHA4/Es4YbuyHptsHytGMC1Wy2F5ZP5WLV
Lqsw76+Ix3kDqrbJ2RzbfbxwCovwQhdVvuKDfXugt1IY3lFs3Ob5d6OTqAMGKPT4E2GmC6H80D7G
TtKF30N5vo190LYwJkjXqIE1TzUHi29eznLq3bkNwKrr2EyF/Vgzh3CPfTfAtpBqNxKVRsp/ySti
jPNUilbfOT/izbGxsOdW2jm5gR6NXJKquv7g9JNqSGHBMdBZ9VIhP/a9CTm6dX6UjYSCFyKBOKJB
Re/oi8lBJvMmOC7woJq0NDe1l/DD221g/tSzdsSNK9WHp3HwDsMmba9Ji6ZVMK7rY+/AUeTCyK9U
9S2vmYZMQ2LVt+F+4lRPBfUNqpkHPPBS27grsOAi5xntzE9FTApJOw966gK4sIMnN08Mc1KRmJwH
oyk3LOe6CDx54C+BRC1AsbIeWPI+yk9jAugKqcDKDTgRTgro3eaEFjcjlLXcvpk23X50j6VCk+9S
4PJ3mbVc2ZvQM28vZnrmgPHQDVcFhKAXy9W8OeRJedxlp3pQXEHDMer6nE2mNKGvc8+wZgWa8nkL
04kVLgccessY08hqN6sBfpniAhYFp/qDuqou+JH/hMuPigNIFOjDZ/xw3IZXtszfXx617qQG480d
5BuZIrJyqRYbVy3tuvVtKZWKWOPs+mRtiJZix2HCSVSJtX4728+okUuzc0LXJ2Bse6e+pS0TpB61
Z1v8m+dePZ5vPxy1QlUSaONLz72cDZB7K4SpT8vZXSWLcjnDHVmMi9+q+JLlBg+DyA7TJFxvBcrP
mdTbb4oDDVDwIsxdIEH41xoAJNkdI3j177T8i8NrxZuIINGdZuuTN7VIpM4HQJl959B0D6+E4NV5
vQMZzddKwGOqkxIfuZjSzabe2Ur8Ar24Lysxt1Bwo1MEpg9FJUY2xOINGaomjMfMdeUMIpy7pIsG
qN9fwdeff59ODuyaouzyrFxXSOKMD7U3tg3BTJNiNPcaKHEh8TMhCeAnau5WTOFBFphqywcjCrnh
k3H8IUQyByTSdtXQLgMIXJsZ83BLC7HKUNzOskBEm+/yGp3inBaejtjg2xrSw+8vAfxPytBITlJV
+GltCINr+mpzL2vbQDXSi/4cidu4HFqKGC2yx7NWjP7kVuajOXpfvdTFNVB0aN43h5N3sqGR9/Mg
FHDCTgqzqm34TsW8dmHtzbV/ADFHs+s9nRYVh6c+exKOvLDty1fXtgFeFygI1N770+db7mYPGqE3
iBE8S8TLryIgdFM7IDoZxGQVwaV46hvg91oggh4xcR27xMyTLLBNHwg4V73sMcxrTIlfzPqWR0cx
rz6iPFrjgupl0ZkOtK/Jj8/7hMlV6IRcsJnHIoZnbAJT/f3o/Sb37dev/3kwTl/YUoHUxVGUjF2k
FKW32NFHF/rArk14vLM0PL7tdc7wkt4PuFcUwQQOnvwAT3ht+5bRuvFbVTvJ+6EKFJaBUZ7LYZ2r
mbW8XxIqiccjobWpt2NpeF5k7WJ/mOUiodmYWw4u8iW2kYZ7P7EgISSUh3HS/SeXILfmlWiMWFCm
+mx9NoltZss/BznEumE2e25JhVE43XySCDUA2vR56FnMgaIo0F8AvLKd4l+SrE2wdmUZ5MWYgvUg
AHAn01XpRyz667onjrqxWRi1HTr3qhPaW2lJwTrXLNszmt0WuP7BYC3jb/T87M0JMf3j5j18Kfoa
xlH8nBez3xDqTut8zzo9NfCHJ9Oh1+VUdBYeUDJg7082yRF6+lns8A2B0kkbfx3O6zhSFL48kygl
Amu9+OAGddprC6jlSvqjDp9zzos3oZKelMH+GbKiPWLEkLof31lWjS8jMYyQaav8M/anyvh8qJcK
n19QfrknftpSQHuYkubuaa3LlBJKMcj1bwafg0aCVGfTwePsMzmDSVkV0v+PKznwAFrJ/0YZ8GmN
6F6u7tet4azuGMA8QHoUUwUWBFbw6rG3yaEIpGUOEH+DTyxp8cvjwb05FUR+8g/8yaKfu6SMNqFO
IlSoMfiUYm2X+g9x9RuEDJwnd99YPlNdhXaVhItI7U9P0doj6Y9WhBuEKTA50TYi74sBeBd4n2OW
I1pwHaDO+/QWqrOw0sVJFMFkWLjI4UiUjpDTyrFcDNS1z48QaF5hL4WuWT1Fl9KA5PNizwHc1tJ/
9VU8HX6x13Oys2JSEbDGyBO+N4n1siFe8XyIKyq2iCA7CXZnp5sA6i0R2U3hS9qFVYXiH61M3tVA
Z6N5zInz5XfObvbmgpyP5kajOBejgwagvAK/35Ar++E9P6/hLf7YH1Z68OY2I7dxgwkm68RsYi2b
spfVB+ETbg1x/DMxOrQMn/hECcaotRP151QECir5Xzzs3g/KhsrjcJ2RmYlwc+FctRRrG7Mcje/S
cBIzjGyc7cDOov/Qo4DZlfmoCMKDFUM9SBcvPZow9/9SjsTIQSkwrTFXfe9Rt8G4+AotmYHW2Jxj
SDfQqvpXnXHuRwcxUm1sTnKit8oaQibLql0wbCZTe0WFo13zTauwzyfkRPJeFEJYhZu3KgMMY39T
r1p4tvHIBTC/Q3T2B4559l1AVH/PQ3vwquvSgcxhQ3uQalkMQEzD2GSMz7gVo2wRRAm173y+irWN
Zv6I3EZFpS3s+fjouqMQGMDNXPWR1ZufeidbYudgV9583xpVd+eUOMFfpkfX0f64NxPdVmgdJDwy
cieumEjsvAnedJkO0ngCDDKok5ZDC+WnypPxO/H2DXp+OEFh+sLp3AX+72TsE8wweYd5eTTV1GaQ
LhGc+FHkZ/l1Lf2tmHGLeyzBoSs84GBel0pvXNE6SxXyLVcq+IheGRgJ2Edf1IyEfd57ZIC0th+0
/NVeGXT3rSBnhNQhDTIpNPPkpehYsfNC5z+izWIpv0yExpG339W5S74l/BIWZrBkzNuQCwwHLa0D
1k9AMI/17koY/K69w8V1bchpwoiPwXXSU6Hlc/hYBuXdyngEXQOZqh3aH8Whaec8lgq5GH78gnGJ
3pcnoeOLJ6IBb2yKKoIRD8g7FuFczBRADL2yWb3XJbjEkRm/hM6uLyy/ccE4NpRrdHKV4Y4phCcX
cY3Orv5r0LunbeWbaPdnpQlCmJim/jxjlJZ3LGdbjLLb7zNI50wvLIGhBF6NP0D6mcAhOsVlgM3o
fSGjqLlbHYtZwGlvJwL/h1EjSq60kvHOWbfwuX9mrNnHy7E2CtyOok4+sCYf0jrnbbojVRz7udKl
wt1/+gzT+bE3HAY8K382hX/bI90n5NgAfiX8qGS1o+oDTMssG0Aj+yjttyd80Y/Gi/b4z63vR6Zq
lqBtl3+E2P8mIPV/DCfoFOlFxDK7F6fBOueGd0Uuo9LgkjnnpGuZaj9AAPfOppv7rIq4anhNmu0M
37TOOLdd29xLYTFjiszrFt5cVamzAxKBI3ZILlUks2rLqfFtiAStdFP1ROu5IQAc2fUvuTUmxenS
7qTfk1j2IVBlfRzpNp/0Jx/YwH44diGgwNJNYnb4A5DfV2cTa6lgOE1xyXtl6eqtzVXelAbiAbiI
lkjoawz08T90R4bCpkkT1Xx3ZKz89InaG4Qdd+8GbhO+BNjMOadACyRmMjyV5I3wmJ6s0FHYCJNQ
YV51OPvjL0SMNe0eC/KdByMMWqTvie9QnOnxYhRz2fvRdO1Ml5EVERXey1dvb3e9CZoeC8hP6tNK
SYXOUnr2+Jp7usqm1Oxu2BWrSjndtGT7cPrZqic00wfeEnLojegaRM9V9cyfWJHKGFMVJEBWWLer
OQbzpCKPZs3IrJfvAErHxPPsL2JoAEQ4OqBFt59QahcgXgktLD4lu/+jvJohklS7c/OIMCpk2KJd
4SOk/lMNpGGBntmFNufpvopWZx9owswR/Qg90LzzYTBACDP0NS8rKcmVTWx/qDopgdPLHnuh+BQz
lopU4XYSyKyTj1VQfjeJ72QcDv1G858GY1mwq82kOxQpefBeyV7diey37mgMIyg7xs2vG5ZXHg7t
oPsD+yaG9WrU40ID5ldvaWgbwnEqLaSl3qazjsbuhUYZZs+DEsa/BQDtHT/cUWP9I18fk57enUHk
brxD6R/dS29hPWyUxVUUS9fx37CDQ1d5SfdBpyqkv528Xb0ZVbdyoWXLPH+y76tF9gmb+f2FiL5h
3z5Vevn1SO2pzPLR2Y4NHYj7pkhew6fjtYzsnnWkiezmTGOyH5KL+r6WVjsac42N+6Qy8m4NJpog
0SSuBItqEpEdcDMsXRIgIBphjbf7YDbmlkGCjq0WzsqzhvSfoVSdgfCExZbUTgk5XgqXDodSKdls
D3bUbOH9YgjGj6o8QCgUpCPaI01B23JX9t5dRGDemPT2tIxkfrBm5XLEbim11jHs8UcdDH2MvY3m
GeoMkobrTG1TeXY5Bg8v6ToUJbvCfktNPttAOtcp6k7AWra6ELvIrNVqS9r5ORf9oJqgSovfirWN
veYseUQOzoF6UAPItnzom+k15dB3TXxxTRf5SbLMzwAG/kpiI3gyJ1lBhI5SwNvxnX10kWdJxmaR
of06PMfAdcPUZbEBr79tgfJX2ipG2GglaPbcbx+IXqebmNfqn+nVrh1tFTd5lJV4IiVxzI0XGlnQ
Z7WL+Hn15i/5Mmdhy8jle+zkyAXxP99ZyktrQ5Y9U4OdXpBk00yK5CrqtdM9DlFMmms7HLhnS2xG
LQYcbxw+F4bQ6o4Vebh3GeGA71VnT1wih/r4z8w+1og2XNVvQsiabNROoL8sL1hOulWn1f1Dkjtu
J4+USC7uEHT5PC0uUsWVbZmm28WoblGBupwOzfhsDWZlqzcOX4tLuqXjbaGscYsHZSl14urRKpZN
j8YRiAWllo73CdAM9z0j4QMRWO1WtbMoXtvVcuczNFgCxjvseir5So1/7OPGoPCyfPV2DBnISwFC
oCYMJto0yPIrpch+faDrvI3yH/dJ9upG2zmvD81/y9+GXyHjtEhk8vV69/wWOhVIIWK5SMnAFKOo
6nScd7kuF1LSNSJ+bG3BqEd9W90rTlhTSGi5pcZw0W2vD72CpvQfIWzwIRyUgmn1QTi7looi4caz
XRu7jAx568XeVKGpkOg+5tem6Tll0kQ2m0jVlcW5KkJmOnzzAfNMsTTLFGcEuJFZ4FnyLJSr0b8k
qP1FVbGYjrHdGNi2aEfcLcN061nKksAeB1vf7Ur4Rq0lCKK1MMJORTkoXCJ7mqogcxj5bZBqrspX
inJcviNQ7CdcAckqkPxnyMbp3HKSRRqOFceN4bCVQ8gch/7iK8LyeOjN03dbllJPQLJhSv3hxjCP
+Z0kADMs8dsVI9Ct5LvWLd4rAg+XmzMwT7ULBFkPoszl4sCsQxZ9zsUliJR5frkJvwihQUne9usq
2wjAPwW7QtP+V7UyaFQZ7JRmue6ZhGeyLtPILTXPqr19mCjZ+4GEDEXDwmttidiiQdJr5sIIFA9N
QTD1tyiqUFn6OD2IYrToAQdJ9q29CcZhRhIu5oN/JGx3rC6mwuunY41rTAXOIy9vWhBNAYbvrl9A
5KPjpAWwKZraay2BaKMFmsplQIrpeHyQhOuO3fENG3twUeB0NbyAeA4FNBnPFdRblTmMkUoqaQ/b
s2zoDDT6KNaj4tiC9ry1ivsdeFlHRWbc551O6wjeBlCJ9+2np8T8QSMfSNMmmuNJYKz0+I2F+O65
CAQ4eSnIHEot6hxZLQMsItFF02NJZNS+uJ+Fj7Mn9g43inBt8ots3BlaF35bqwwOt8L4eAcdtO1J
G2AbsKGQa8CaDHL86/4IYAn+TjBypvQ17r1sjULJmlWk3WneHj62tm+QFqs0wVEsx6JLJd/pQn+h
z4Kmuh9wTiwpL129A9jB7G8NoezQaqMgWsQdyY6voNxIy5spOWzjx77Qqd8SnynMtTnNhh/3+qHZ
TUZE346voM/BywXCmHNCU4Gtv/ODTZdQBOwV8Ql6wQgEiOiRjqr//pr6QbnM0WjLF3H7ElNp2NKo
YH5n7WF7RENM9lnVrAbv5roOE/wXbD4Z9GsmWLnv9gPtvEDg4SRWBTLXjfyBvcWm7uhUwViMA9fw
6wKgA3rJFoVIRHEwvTOaH7t0m+XWBVL0ePECQ1D90t6cK4n/bz+1A2bBxJzkrUCNx0Df5yLlLRY6
Aomcv53y6AObsXUxtQFVj41ofsokCM0qirIiYZK2JyxSokrirWfZr1bDjGWsQSchjOrn+JzHKjmt
LJ83zYHcWl2qhqQgHBRfCZ3eyDKWBgn1y2djMhUrlrOuYXSUthvre8XUYEdH38AnnKL1DJcji/4M
gIdVY6+CpMUUsGDxurd+3hEM77u5FPF3TlGWD8MH2LrwKfMrf+CO32lE4UTjusYJcWfSV9Q9FxJS
UebRAxXtkSCP3VXvFtD4KN1Vmzy71OaN6uwkRmICRxuX3PbNn5YWv/MioDEgt6ExQmMk124dDAql
Wy0M/zpspV6qRKg+/AcNu9Bv57vs/Gf0A6w9P5dFYBLNbJKY5KYR7nlLeRblGyP9iwHoltrLsNdM
exSEE/5dnt68EoZZ2cwMb7cC3aImw7bbW8W22A9AKieVAYLS4JkqSY20gb1091Ka1uEO0Xh/C0i4
uTWHQlGEWSBpEzA3Iii1pud7wHu8kIhCq5Kz4l4O+/MMq+bAnTI4kNT20YC6VdbxtbCdebdSchHH
5hbPEtHYugsB+HDANSLJ+COs7l8OSLuTw42sJiIwXsyeuQSb0LnIemFwxpqs9Hb2RsGFISjkODpB
TuS0q4GLTlQErh/KPdG+i6R8iORBWNP+OhsJOVHtyPt+r4I2tppKmmtEoPDQ8vsuFuky3ekVCLH5
0dxDQVtBoa8mVzeBSGwNven97UD/jM1Cepqy4Mc22VrOtu382l3krZRkHfdaYsAwH+/SMOygJFB8
tsxDiWkSmnMVtuCgtcSdv6VlKwSkvNGTBOdo4U4B9tqnH/VXaH5FnR7+CTyB6OWNFyPlM6I153Uu
81sBZzqNcPjKqM0kD6rkX7Nj+LoYnhhzMzbMKPFJ0jaLMh69o3auFf/ae5kG9HeK6PX3PpCocUTs
I2KUhr611Szd5S87Yk95+n7t5oBtYUyYqcQWXnHefUplpjcPKTdUSzvGh8BbvHMTh7+M5226e5n1
73boX/FX3kfDIvfkLaa6bqDycz1QRRwTNTfMAr5yn6e76V3ozh7ttAPu7fEO3jC/Mt6M9OCugp6Y
NDPYMU9gfOtDbqhdkMapBwKZgOgNUPo8F8bmJqtjeomtmEuknZw4RKR3/dW6zUaMsd+II6XizrZd
D0MANT36DDNz73MmEOn0ZAaG8nU7DAMeuoqKr6YKllbu9BKyoqu8S2UApWnRe+hpc9NpDH9uV4g8
ZumAPJlWPxtAqZwniFLenhZm7HpzXuEs3tyTqujh+1UukzkLb92oN19ImOQ2D6G5jeptP/+39A0U
1V/XnB8GGC66IV9nIVQpo6gVoJS3o80HFUmhVhZceUUA3shgmpVOPzn+70Ekprk54g5xXuAdKnjd
wb7NRkzm44VlmPWijwDF1so5JEZY02CfCeeeoo43BN71wI3qRD0vAPCwgwxtcwsjqQ4dwuKFINdP
TUBawxNjWuNOSolXxkl/cwN0aKVYqU+2oMP60yRK/RIC9BoeNT9fnrWCZfw2ixlbQYoofoCEtSx/
giyhjcdBoaLNiLU5cY+vhc3ylTtt2N0rwKKitW8TdxXtN2ScFDmqxiGi3PGyHEF7BQoO3vDAApyx
MVaOwyLMUmDkLzCLk8qk1lK+Wv1mvGps73smvx+KeOLKIafKpGXrRxlo7Th59SQ2x7JUJyrl8YYf
VPen7TkFMsEg0iyngMcWBYyGRh9XuXqq7dgzXrw5yWYKzo+RwLuVq9BTXaGqDKASuKor4c4IoqNj
izAfG6oFj2Nq3jaSf+DlrHq3pSVhnzZX1exwA1zNCcKITEJi5avtmhGD0+5Eh0BAjbggp2b2zkmj
d+otOcs+NFfSiIuzHPva4Ral69kRBQ/kkFAjvDuKmQRPkWWRnVqoTY9JoWpMdfsFFEeFry4FPimK
K/YDKLsUhe71l8Pdsf2MBZTDj6TxAcBAnOnr+cXg13rR2F9iaIeWrBHjXUQueALy9Miokrw5KULq
O5Jhh7aWEXwFbgrzHDkJxSKSFUufUASjO/R9YXuMiMVSVMW0/J6J0b2vpU2c2JhsBBHRn3Zv0E9I
kfBOHpj/hAccup8HLqVE1PuYQ9XH7bpH4VW2rYZblOZH/rnT8CYkcj2q3iD9zP/TCPeD2/WDkYAM
wY/UowtTtVe5qkKw4X7YHfQNQT2YAc+SGzX7sc8CVUB4PjLxCPKEM21zh0u3YLSq6iY3r3S4q3LF
PDtQZednUEuQb4gGye2b2qwVQcq8rwIssxOVQdAnyAv72q+UziPfKlNT8JZPvUpYCNbe7UyIQR9A
dNA8WwzmF4ekWEpwc98M+2be9G1XU9mYL/2lDSWW+rn8HIZZUgT+7FhkgaloxpzJ59a7ACRnc9JU
MkXE8ot7D8FncRoAZGEoKX72P9KLP3L66AWvOaw/IFKdqlci4WfujnvJpj0zsrOfKfHltvGnFt4a
unWN8Gvn4nzQsmhMrn3ejyRuVhQoTIYZaymnLSFy3Mdb/zUd6vhKnmvxIImA7un1TICfd65dVmQU
NEyOlhqa7BUrXajrgDLEIL0LmUIG2FMrzjggra+iOiS0rB02r9D2chR0wvPtesFqfgrrzaAIwA7B
JTTBxuT0jmHh+egGtPeKUqtPOD+hO5sQi6gxQ/40u35Oe8YZpuN67GhrEAcjekuv7QkSVMhBnM+X
kxHSXYef41Knt/ESZb+mY7q9zsdIQXuja6vfWfMGliH9xZ+iWoNHxi2vuASebEcTlZPU2tusw/a0
t8mPZ7QcgoXppPZi4pS935SIId7IFu8PFbhy/QfJUCE/KfpcfczpdaD/1DtGaae8P51qnmMNqT5W
3QCOx3cxfymvq++OuCcwecyAb5kkYSRgxnl/f70uHoyzc7YeFpobc9heTJe+F5JC8ej/0YIYAjY8
s2jMcvI5zu7HXP/heIfuC0JrwYlX8xzx3syuP0LIkgai2+Ctf9bAoCq152T2qqcjGiwzT3mfNXya
oXwF1BMLaA8MoL7gXXX+5Demqon7GTJu2A6XY0VBLPHtPHZKxHYGZAWghmhoek6kH+Snss7BlKdC
9+jt6tM1aOgLkznPK3KChGBGXje4G2dwqE5KkrRn+bD+a9tYdFp84sAkcsrHMmZaTAsIk7T5c7a0
WA5HOmWLJNXx7qM7bDrJSBus9uRXLMZ/MGWpRerel5jPe6fVd3jbjIYjsR9HoRRfNcDTXtX3r+Nv
nDPQhOL1SSL8xIpBdbVWSrid4vUu3hEUI3/lZKnIhKWJkoE6vUFBYxNSC5iLD2qOrtxYgYGRzwoo
BNcxnJ4ShuCJMGYw6zQb8JEPWO2WGrCw74MQDp7IRojNYRT9of1vAIHdAVWaacT4M32ZDuxD6dao
ikqZw/dCO51dMBsbO9mNrSPeqvOr7+mZ0zb9BcPN7xJpeXzX1Jd6f8D5acvW4268bICPBg0rIp1b
bAmcdKvU7UYY9RMelfBSK7MppuM/wdNp0V0Y75vU84UhxNLBE9Baxea5xvX6zypBjb5cm8CFGUBn
mCTjsgwTyassyPGVgqTyvgrrT4rq2nf0jkgSr9u7BfTJbfLeoVobGG9xIlZPvwHYTeNbhvH/5uqj
+Fr5r/9MRT/fr39vw/zS9i/MMEPRn2yvGxVW4bYcm0iPHH1lt4955isbLR9/hYgjWzdTAwHbtynl
kUMBrfCjFpPaeTrsjtSg+PlgkS+hOXBq3aR1IQQYxex1WFMvmCI631/ahAttOdlhWoMJT8ZWNIVQ
HrnzZ44IxnBD2Z1++IxmTpSZ1KFRWfmwRavE2aH07yy65AEYqwYMeZF7l0ZkeYIEcC6I6WEgOmGn
JsraZbgGXmZTmlvcKxz3AioeGnoX/N0ci3uHp3U1uqWJR/sWd9twi1bHuPvzwpekFCUCUFQuYSAA
88X0R7XcVtolrgnjke8028s6ssA8eBzGgEJU62VrLsu0mAZWzPEi76SnE/zTforTlAX2ma4hKGt3
g0oQo50LV11C0LmIYM/v/uvLfO1tadLJ1hyKhhO/hrQl2QrOuBzRMVROFeM1ll1jUy3kKRPqDp9R
iu/sqQ5/UTMWFRvijKEyW2l8uxQHbPbLK4jxGel/b4BjSdLYAOMwWHK7jth0vLyREjaXI2a3jP2C
1+y1pFPKjOVoWH7hT9ILxmMVPd5Pn/iCwMO1vcfrSPXnFNT+WY88aj2tZ34a49B1p2ZwT8uvd1vt
HneeYeRXdUMLM9Fse3Bw09btVt9/qcO6zTRmw03DZLoFHGj3sIA4DmR1WXZLNEsyfA+rki0L7gbL
qL+9Pittun3deiv4aTMO39DCC9nGSW8016Gkra0zRdVSLNK43TcclMIbPXngLom2nh8wvkGpTgY/
ElF6/0hz9oWL0ZsJ7SqGmUcArp7O8eJom3FUXbM0MUh16P9Y21vkMUToPlTTUydzzg+pXYPXxSGb
XJadl76SHhG/qEncWk80WCEXp4jQ1gRK5EtNu7j9LE3SUkricw6PxgtZ2wzvD3SIgBfZKIjfPvM6
UQ6OW2REot5bFTPE+UipQqMLcUkhtkzOR45IvS8T9JSj37MqQXVKlkdFznfA5cIqnngJeZz9osgb
vBrlWf1jF4fe0bG9d+KgscgY85Roau3ggPPFdl/GJyYv+hQl3TU6oQMaJ2vtJcrb3HnqdSTllMPT
NdybBKcqYhjPnYNB1n39jw0kAfil+IfefKiBU6RBhADHniUNFLaEN5pgT9hQDctnLDVcGTA2n1hh
KeZMqeEkyEn1nLe+M5bYqGl003BFrPAepzCjcniy2nGseS0+M2/4QqX6srBnyJXwYUjqk7v53C4O
mvuQzd1ZFkiqkGvATZMfAzWYrNQjJeYR53hQ41V7MA27CwqOBbQX6KXSh0TLW24sXKjo0ruu2K9w
gXYxT2AoeI9T0BiHvLiNPOZLycqipNevy0HTr6P2c+YMfmxAUhKijmzixsoCIjLPeSg+IPnTzOyM
Aj72SYGRYAhyEg+5zyJldL/n5MjPj03+6WuhanUX4FLYolRbYvymMJsktAgIaTQ3c4ixdDDDwXk2
0bjWxNkEZbsEsAW2jPW8f4uKcUUeUkiz8fWwPUE0Zkb2czHXOgP885XVjZzs31XKqrKMA48CRNjN
vZ8y3cVO5iFxMUz7/xiZ6q7/2fkE5kAnz9NGL1HYbptPfHlHJvAtcTfNYMkbtd0exZFFFVbF0/Ew
ncuPd/st95lPXseSJtbgOoFfaLu7IsyJGE9EB4/CqsUHWxkNyg60eu4v3pQAxNScbyAhYqMP+Pih
GPnh0W2EZEkiA3pNtyth5yIXUCEk21uYLdE7jetHzLkNa3jJcxJHIZ/N2dFYBJnqV5ao/s7WefKe
WL9IMEGvXlxZ6SGSwCgOGPl7m5cBS5I/nxNr4o2ygpEAKxf9LjNMYbrnjrpn1Y7MjbhbQzOqXqsf
hqrROR3N+rqhaLZGMJipBYXPOu+hAsLSqG+Nj7GTixzfdYvBepLAhg9t9pVyZ/UjERpLIx2yzCan
in1o7okhOh0vw3OAsUsWWDZaGuL0SmdF2qEzA4HlnUdYNwta/8tutVzgijKTzSoZ/rKnsluCidaP
PVxSgqnAciwES8k5SJ9qmhT7vRA5SnFgBSkBNtFlu6fobDFziha8+HcJ6dX++NOKoe9tRcXmJdWN
qd9uo57Xk8N862G+XZyFMUS84lYm0suvQH4YRVNo6sS3YSfR2BYLSgfYQLEV5/Jmy+8hlrXEdzDk
y/8Mqqwz0ndFSOMFEWLIa4AjF1iguvN91xbp2oXmEGpfUFSJPbwIoBouQTh0dlWePqwnSD5e7Fa4
rhFPVNyY5uv6G4NFc0lrSvkZ9oA+9nm0RqNl/PPoBIvTIPbxAJOZxEMXleRp55qJJ81YEIjxnBTn
vCqsIZoeqsZZ/mP81VB/nMXHSq+3Pa0JfQS5k+8M7n6auAuW1/P3VWNDd2a94ij/Csy9oUTRyiAc
K8OVB30cutURTlDjCV/T5Td0gEKsb6QaBpnmMCtOzAvO5DYBqAtb9F0kBlrHAILUzyUU4a3Fn0zE
FeDEPQ9gQThTpOF8JMGcJ4gHw2FV9uK5FHnpe2hEWDTO1agf6u6qyVqiKBrHae2maaeH5lPCRhxP
Ee6D2oIQ1mTApSm4x0hpBCEccBywlEIC7Ke6Y4NJYiTe17WDs4zGhBCjV7QQe7cyzEmeG43kK5Zw
Dv6YMTq6blKIVIX/NN0341gUSD+6FVKZxVFInQK4STl6eWe6gSZ5aC0TTobM1hR4A3GpTw+tLEmW
gbPFbcO5Y1mBsqVxTn/SXVluum/RaQZ5LR4Aqh6Pd4+RPL2iTMGZ2So9NH/3hBqYrlGHp+v9yCvL
xUAdBx4nAQElrxoKxTD/2QtEk14ZszaaA97cZNymVk9CvqzcnJ4jyAoCKVhUC6O1ILBNRFgHeMd9
faiRGVUrpk5NiAqhbTEtOEXGS6S7d0lAWm0s4J1pw2eOfFHJFP2gGBscAGYlicsvM2myJVnXaLub
3+ltc66pnaHU4xrmltN8NX6Qx0kxoPlHogVODrS+gIBaHAmmQ2onS1i6Q+e3iYep6/SdF7QJNr5w
E0U4+EbaNMYnOhme9a+dZEIGnmW5QZU3d1ZICCv/dfbBMDk6YWjSd5rbfrAzFDHCbc+KwC7/pMdW
5VOW0pwEj9C1b11/cpXK9ODF7dpvVIWcTtADyDWCN8IbhMgDklSdg3jDwgZVAyx8U8wjmdyPIZws
tQ26GG2j3eDy4PorHipOjPNac6yPByKxGg7KFiXFBDNNf5yWhWof8LhSoR6NOiPQYe1ljlIg8aU8
hrNM42TwLnJdmhlTP4e49uTSAoHrTnLZfXTdJXVjK1YgXvkazYuu+QCBuF0uNcOz4YL2rxlkgdzY
rZnT0qybut652fEA25S080E7ISirPQ64iXyzi10xnZzFrhAHJzv90IsyDkgyI6bgwbh92aUxCSki
SXZYKKAzDmteviwaV2UdI80WdY0PbQ/GYZ629wQkb7aG+urX631JUsMJJ8NDc/5m3YkMN2yiDjX1
NgbsFAztRYtpBHChbfXYNNP0pjH+1a9lqB2BYZOpyFzOT+SBH8qB6cFCXAUSrlnFAgV5cWNbypuX
GMiXIt5Cn4FLi+144aJCHt5BilZXmXZ7Cuy6Bwt38vaIzBX/Ou+P3gKm8r8dduKl0JofGkPooy56
j0zRk8WsIHcFnvPzjJrpzpo6g8oPvSlHMm9OdiWAHj1RnCmgpAg/qvFNmEktb0LBtqJB/e2+v5Yf
yrfKuCymkJFAJfzrCo0EJx5RE2WCbPvMp+MqbOJzMGRtWgqp4xOmDz1W5cHQh6wgTt9YAFbSX7/q
7f0VkfprlUFQdnMF/dE7Vg1brTXeEolXwki41Id+AV+AL1RTZOUP2BCDj0VZqOLf/VuVlKkgcNNj
ymJuric2gObf9l0FvraCPYZ6vpMfKEOnHANKpVP/GAL8JKI3HrI8jd2eVI63JGr9sqVEBvXslKHh
jXKNujnPL6sYS6rCpDRC4p4rUFaez7Iuvx76oDpsbjRrhCj+3DSBhOhHHqN6s7kJ/iitjt6R+7A6
Ip6e23kemA6It/LLhJy2gjDKIWwSQcSFvk8sYBy4ITaJPTaid+j7J+Nx5CdG+3nQm1c+RoxUg/xB
mU5IKdB4urrasn+EREwF27AdY3hx2AZIuzhZGF8KmYbloCSuJTPxHEKQipnVKzr7ze9PgnKSXjnP
N2midhmCrmj+5A0q/3X9D2xD4tgGIFfGGRfA06QOtxXXmnrceAXbzK4S5SPXAImtR5BCqVVyvr8R
cU966W5v9V3SY/ayVzrwP/JGQkltU1dHn8s9eKR9YT0+pd1XWyVIFiicEALRN5z6bf8F0wn2filc
CmFWDC6DiIphOcM0TMPUn8Lk7THRgDhGC/mLd/bMIdhrin7PC8r0gipk2TzlhCCInQCOU/Vyp5SB
o/kedXEktmqXOtt3yCa4HFjnwdHvDsW+x7WMVzJKBZw228uaO9VLn7WS5EYHPv9krCAiS02D742w
pu7t+LVZDiKFeDAUilz5xsyK2ChxqQ8U9slJm6aiSOhosXBfhdiyJnmojPgehVaz9IQ/rr3Y0+uh
YBYTQ+HvnpsM4yjBVpYsXOf4pErjHnTM5BUrP7fBb8eJ5NDCdyNvBNq/8LOsbi0Wdy9Gae1axS3T
6035sQGVTvnEg/h5aTfZUZRYUg/7626Zf8i84cuj1yysYKTBOuDXF71LghNBy/1HCn3q8IS8Xpob
LCuWiaGAJP5E0gvHpc8hW56ItnQcuw3IPkDnT1Suu0dW5/j4eLFDozZ6qM51Hku1ohxgj1ID4Lc6
p9748PZva4thGxcgnyT97YgxU6elgQ0AGljG3qobcp5WJRLwDWuWCSidaHPSOX/+arV+2H2qufEn
ZsqiO6k5taDRrntl2wgRji0sYCZQ3t8sJJLfsrDJkPj/HPgPC1S3dpNbW6fSp8snGy4n7f799PoG
DBWi+7fsDy9WR5fJYZefIkVnioM1pcSFOttDP6sA9CxViAvBxCMovdlsenFZA+9QJ1t0ZLgY7AUO
jcWd8G6rXxWrhaLp3E/cfjCeYIXqlnJB+ck0x2H13ctgv1u707STTv/VnAGGBWnY9++SNyLCNW3w
ocZOY7+2eysOKMvGcAeByxScDuI5ABmubIIrB+fk1Y+nbdWzxmJd4bc4IDo9dprRhoc8n1DON9js
mchxiuBBbEpZ4zOuAnJYBkbGGUMLgL8hxlArfK8qH8gcwZTB4Yt6Q2uMxvOm1VSjxQxS13X82IIk
XteLyL1jUvjdQMFtQfAv4cL7boTvSWy4JigyFgjACTuhM2ovCdGzlpwxc03PkhYFcIHwHMx2MSRM
Fmh5aLPMoGkK2O5jjhqi9WxMPOFlnEDkM1w9CR622CqXjoBg73QumLJw2o8/7250p8Nn9zRgI3uT
+lqwBjEd1kUy2N7yA0tyiJbkGCgYuC+3Ug4g1rrc0QQbiVAfygOL5mCN9OFF+FxY+qJ6uvfK1pnY
/K9kcpMSchGUTnIrHc8vSTlb+1JTLZ4O+2FYc1tF66X0eIjTJhbXjD5z8PhktakvrlpOr+X7IODq
DoTq+UQ9kkVkI9NDIL+5vV0k3OM+7UN5ou0K1GOIOn9P5ty1hAeSBofKHgAGSfVMAPlNCB8wwtRr
2R0B/1xYzT6yB7OTMHR0hg1OZvGH2wbR6T9SrrKjMaNcpkGEqIeyDdxKnRrjXkoZuM05bp+Et7ML
moMmyMRI9gJHm+yCHo5L818K2Yw/K/8kmSHAu4u913EKQcCRifCk4DyP2FOvw/ZG4C0Yh9H8DpZ4
g43swmSgzSGHD4/3efWSV1c1HS0cA0cLShCboPDwDJnLRxsMX5FIB+qeITzVaSecMuux8gWLZuR3
9vZqd+l9rUn0YreGfoZ+Kn0SFHdWXd7j5G7h31q2mQQuDi4I0OCNUoLQxihQwjS5XJUDzw/x+SA1
gCgIdhVIzKzEmc9eRbsty0KiI21QubKN7uZ90F6N9s1RVwk9TyYyBWBO6KQfXOmUoMFJZsp+1HnG
1GPukRz0iYHcWJ2zQcWIm/n2UamrJi0oNNXP8US7aal0/RVLWT8AWsKFBCrywmPhRTpOp3xyvIbz
l2aU1bFedfH+sWiD5AsCevzUv0KBBUNCsgkcN8uIHOTgOCdT8UjJyaLSDPnKcAd5IUi5efEvblxi
r/QG26MQJ22si6EiKHMbGcotPN89OIm/A1SauH0tJeEXPnmRGoKD4Y2RLC6SKAHvw0mzswuowyu+
iYipzsWJ5cC2xPdXlfcVpClUD8Q/tmRj9Jzv2NeHe738KLtUAVxpBFNcWTs0dvRTbat+6mV2Ca+c
P4Hwb3ne0mWiF75VbPeechb3pOh+quiG7+sAVEiFemsew9Wpb5l34RhE9K4yH/91LJDn6WCzOOEX
xhv/kfs4MzcY0ylj/gvvXxEHdjJX85hFcNLO0JQvYuFKQ+k6ifZGJQT3/Glq6e5m0Yw6VraHhaKU
dZ5FZdHSIC8iPIyI3AMjSCDImRTDzxw7IWTDhFzM3pBjz7XI1B0RVw2eCLKUvYQBfhY11qMBRdsl
vEc5DgELpIke0VUymFXIZj0A6DVbOQEJayxwmYowc/Z0wlJnS9ZsHF/yEkDN16lHqDiYgqp2fCCE
NlDnSdbycV+xeLwMTEYrJux+Jg6+oJNZSUaur7e8uRhSix72SBbhFeubwE5rgQuMgsYLsWNjmfMW
qWEA+X9Rx3wFsjoXggi4wcLNnT5bGAlGoYeYjoZsWjbcDxibWecCVLehUWFMwP4/N0gQaGKV10Ek
wTPkVgzE76AllQKbycho6UFflktvIjl2VCN6KdyfiEfLzn/8vemIKUFjRZznkOR25dWKzjz7L1uP
MTk4BEooh1wJEcHmGzlwa3rVJ9rtdev8MDxMga7PhaVlHhgelMTL7c37bvEL2nYviU4i5XI4S6aA
2nOs3NB2iphoq5tpt8dmgyqjxpyEht43bi1K5Ll4JgaUWeQweTVhttRmicozCb6mBNPJWf3dANYD
q6JgVvWRCY2/UuwGPd7J+9wEa4P9+YhQfemrbV3Y9dXGgbXiE0WTk3W1W/QwQxqdf6eAgUPMJEVC
HOG87NsZEo/lvG5d3qwx0O/aVnM7qdq7Z7rkQh4UIRBBv4yYi88lNr4k2zgJ4mOhAgbVFwyj+U10
upyFaARk5QWDAvRJUUCAYx7zaNgJDaaWxTsNB6e2zooMikxANHQ/JsSmxBRD4KEE5EugCCqk6WFV
LrMxURTP75JAo1Yg7OEma4zCz37Bd2sY/mVXXqAhSVzZXFngrY7vwzYmCSfw/HWfkBTzZfzEJyvf
ScC03gotP8MujVdSpJDFYo5qqBWKTn+WI8Hsu2LCRiGfjVcpce596RjkkSZJYQGLNxshHuo73/J0
yImMJu48P/gImgNvUq3hPleTt1FbseObPj88b1EaRilJW0g/f7W6tv5b+6nfGwHSudu3M+8uVzLZ
8tgGTf7ORu6oQngZ8LMAv1m/IoNN/sUZgwcg/9mcNGXG1p2lQ8l9kJt/KjdJIBZuMfhf3eXDIVtC
Od+T67AvGflS6gSMFWcHuCh7LASe4Io/lrU87U7oRRJfHWb872fAo5UOHGU22+mOEg4xO0AltaBh
uLn3xLPxzl97+Jg/io/8zjjpSBfftgmsZXcHxKcOztsKk7uGhK2bwPa1XuPjMMF05+dwpuV4ZNhW
1+AIkAZIeQUOpkouWM3/EfFa3RdzKWY+m5KJs+FCp7mj4FstQb0z2b+eB0Lht4P2Zd+vsfp0fs7s
14RLpNnGvkrz9+Sx/l7i2wZI6kxyyQhTe2iZdkWGX2yGTluiSN8JfNwais+7YOfNNHzBw0GzVQbW
TWCjpmDTjpEBRoGZOZpnQ1VhkYEvjW02mY+VSNoUuONELewoAjAZ4fuJ3lTWNWkRqgAtvdu3DpIC
2FmldH3Irb+U91LrI6c8dLIRvUusR/fh/iRrXgr9SJpJU0vk0G1kThp4/WYdV0Berub1mCYbtl7/
xRNIzcbMDIonyaJo3Xidc4F5O8Z+5dhJQZZcWbmSVXNy7TKc6dRDzGwFDIyLljGt8Kuord6HwDmK
66OZbySnjY1j4H/pCOauMk5I+nVy8NaDVxvUcaY2pMpS7BqofPxe08x1sVxwFARb6rnFw23Conif
cErX13BUpsrS/lqUYQx6FZOftYy4eZ5L2iRsGyt2ZmEYro99yBHyuNdzKNMVEtMVmhopexIs8zsz
oRZAJglMF0RTjHUb6pCIbpMvQJ3BDiBzIzz6D8sZQBTB5eE1sqoLH1i2dLrk1asPj2+AQst1Di5i
/8X+lodNpzeZyE8Zq9Gxqa2XS3tq1ZTsL6piySO6iWS3qFPBS/d/fRVGw5Sh/9CeWT+Y2QsMmIUC
FDuViqBxhLV/NDCCyWoclW1A57y7yl+IJuwOkyyOu/X5Eu6mJ7O1rXq93je399os4DWIQj8OeXoj
8NijCcv3wFN824yeNf5ZkHW89y3AJ+YW15eSYMaRxoza8Ca72ulZIJHgJnOCfrHXNgiGEbIAKQHC
PbCil9CI/y45Mvx3wL8eCHBl+FMj26nJoqgBKHB6btudic9gddML69HK4keo0SZXFLIn/BSF881e
wajLzXx5+j0T1n2vQnFuM6d1fndfhpBWcCWr3LqHFy/ruIlp0D6f6w1BzVZ46wWVAEV5TnEyfl0Q
O4li0AzQtfeWNPv++SyHBNLhGiMRPTToCYz8V/I1Yko3I3O/IlbVP//GBPSxd2I48YwNi7fJZy5x
eQ3tZ9ASkAwMIVRwb6o8nNqwj5B9+9isvbA9mfgCO8JurHFBfwN1G4cdAqy45i9O1paFEJuOUxf5
da+KeOq4HmNJmOjL9Y6jDixooayGs1m7s9iYRk5/bJhOhw27hOTWh9CyFP8GuGRxbKomUNwwc1qF
ZbfWE3JpPPkeh3cjhMZ8QBYW/HrvV+Y7Xfjtc213ew9ggk1nkhxbSGT9M0WdrxQsruChiP/oHFj2
tH7/hAG6ubqUXcQSXWNhkneP/KvuDy5nwfmU9qBhK6SR3P0Wukh7MjlXhsKj1WFs59G/5LySdgWT
bGHCzGN4TsnDXhx5sk+78M5F1Bv0GF09tXNZVIVOOteY5J13Q92PQuqqNOXwJAM3k6/KjrN45Bhm
Nz9OjimYD6El1uNDuRKw7q1xQtqVEXs3TLj7WtySrmV3pDHZHcTnXBR4BiJ4P8NI8fdDVRARx9Tr
FsZ4M1EmhlbnFJ1Qq09nB2aHhZxBDOSS4jVreZCeXTCXmiX2nN2Q6zQrHQbWKRyw/O/6DMZ6obzU
vb0sy3/lWRnppsLQKExnNE4c7pjYPPH7nzoHOqpu963lyjw/cnn2hsh7BDforFBnAv3+gS9M8F/x
3laHn/HK7ib59f34sKYsYxCp7bJKmF/ad8R2hdSZRQArws5XIrLmzVOG7/m4630zbAeYLqg2zXky
156uN7AEsFXk7qQVYuFGZvI3hInibwISGNvF+bXkLu2msM8wTUwZ/cYtoWjLgfl0e9XVs7l6VFn4
f8E0MbB9Q4XrdPey9IjZQx7I7MWimAZvk0EbPt3ekA42j2UCLF2q5ZMnFVh+0D+Rod/jw6vugJh7
WnfPJzbIKRkvfcq7w4Q1Gz8/Ee4li+YCCdsToB8E0uxN03Y7bSdX9vl0DCoCNTKUcFOVi4dyeWLZ
VkRCgkAxDQcLk5/kyB7nc0/6oiSzoA5U9QEHuoEofy5ADeHPPM5oCgDlH9312lICSHzK48mv/AqI
dN3PfC2/sU9Nh0g1dJgRzLSqd5wAAD18aAMIEeGF2GBaxtckZ3WeV6yyPG4v1yi3Vey3/pVoo3TW
/R9UVhpJZEvFGLUWqnk3QqTgmHUGvl6KOfmH/MZ1k1NvlbGjaGLWsZidSLezZ+XezI/oattqQerP
dTmTZNQ0o9xrFiO3HoJMTT74hlVWRKtt01dvvlOvWBr6KBGFsYv8l9WoQIqZa24NynTQyZ2qv4oZ
3ZXsx/+U8UiqYoA5kLYrq1eT9PKk/bpFd2proQlK5RP8jlMw/srBF/RLlRTQcoRBK7Ci21J4aeJd
7oGRAgtfsHBA9AgXIEc05pkH+Hgo0+kKcccW+xkdtnLScN9jfeq3uE+ygaAiRJsFZFsPk7r/Vd5w
Bnik21wciVw5hoFzp+//a7xg0cu3gNgJR9JicsZJLFKcyyraaCEYMC2usLWBP+0XUBBO/KWelfLj
olnLJq0MdPZ3EkJCUZhioYKx2X4Fg3bvy0CoXyd6tOfeHbhhzQaZYjaYq60Sza7boem3ogmHs4ND
I+CVymzh2eVELix9ZoUTX0W/q+fLg05fO9UDhnE+1atuHUqD8IEvOY00C33X9TRgKppzzNMVNh3/
DNfrNO8tqA4/C01UhIcguTBosB/x4RM4T/rvNRlxrUsiYnQY4DqziHdMV2Czpj1yD+D/wleeUf2n
1n8FAJi93n4wMQOrlwFK9fyVuARu8uRmHXyhxZjQOAELABpPtI/JINTPJT1BeW/hbiSP0vleurPC
FeWO5sSvShno0JCoqhfAcmAne24NAqn7ZKx4i/N7nZMKh22rg7jcCPJUcJUomRcVNyC60er3j1f3
Sqi7RmsyuwZ5jtnWyh/Th5/oSZF88+3x3T8+yOhTT9QgTAfONxI/2xOPsDg23f+/Keqz8P8/C2Z4
16WSRFgCF9LHoJqBcLZturu+6TeCQKW/HNNoMk7MOs6uUVn34LEKFqw9XrQlF2/k9EIA6WfO58JH
js8oPXsTa44nuBX3UJfM3gYBTa8PKoCkaoz6c5USvcPw1GVmBgn2j4jUZVvcEm1ZiD12qA1mj67e
8Ur7s+UrgADG+AfQwb+uEbgx7NPRkoJYD0C9bqmAa4F8x0vWlJCdZRYVHGHS5uhjQdLirCZaWtTD
Dk4OZbVtw7MbU7gh6QWitNmRGeu5rzZFiNYSqUqQSjy0agICxCBXp+U/Q/gt1YxVakI28pFxoVMQ
FmM5ydByUlJho4OiT0oACBBTBqx8H2ZOYBFPoyP9Ym5wLSgU9sJWh4w4MBmqpVjyuKU09tadj4hw
vDro6BdZLbFw+b+sa7xdrZMpbtOqmFiHqjcqQMKaTjbfE1lbuWL77QXKz72ed8GdFtKhXAYXtsTw
qnYGQdqrCVoexVREBHPGZSC6FzFnD5R1NU0hnpZoaTzth912RlSZ2hHuzV3C40/q1/a/kOuVbFvh
c110uq1C9o/YYuizm9BqiWZ5SQ7Y+hq1DpDOrYeIKpfbOTiZqHIYKL/OWlEeWnOHGzxpTFsTWpkw
CGPc8kar4Pz71LcZLab73sV6fo5HAml2l20hYOmB7cYsj560YPixW9f9BPTM1lXDZUyJPQvXJkJl
Y5kRWbaAmzV1tXXB2hHr4Wg92sTsQDSb/lDpnGs8rZiSpdmwQ/Kqnh3slPzBsF8171xxuPGaHapb
p3U2XrZm0nAbbIoZvBKlbrVVRcvViTiSCbB3if3dJTwtLWgItANjhr8WDFGggUndYjoH3sSlwS5X
zGWBGWaE6DQcK/5eIjSC4OfrxuUQfQEJ1fdEWV65iEx5zerdoocfx7DUAgewYCCFycp8GPjJXcpI
PuaXVTpweIgSE27mCnfzJ5sWwGL9zCMmN44f8HsufAKEmFWLWePxjXarrU4AfSjzEHmliSkGGkwK
n9Xwn/WygERE4jGWOwbDEEeB1i9eh92PZ68MvfdPb+CuiAvMpKpet9qGnpp/Vz6vBBB+VqONyclg
Vq88zKvInCPVpo15SfyddjdwKop2UPEVpK689NzyNfFXPbLFTwt3xu1vz+b3B40ZoRLk8JCSyCF6
VjTfROwUC5vDGMIkaiB3rOAgImKlSkKwR9yqI62GsmQn9ZqN3m6UcfHHhRyqet2mzcNIT1CSL09l
GZ1KaWkf8w4sQYBn7adiboEGm+6bifpurAe7NHX0k2g4IwfLps5Uf/Op24Cp/EAlMO2e3O8OpwVx
OkgOu2WcLwyaus3tXkMnWy82Ui2VO/++QExUWREgwj2SRE9zfgWmss2kKGBes8/pXr6ZFW8kBqpz
olTEKKvdy4s6HtLeYP+LvDK5Jtb7ov0yIeStX8S+KyvUcOsYe0W+tYUDjiOx64G8X3ug/ftXLkCy
99a4ePu+bt+Hs3D10wZAXB4flX/ypZO+tmqh45BgibMVj6c/mYHkFQngwUpY3/bGl2RiG0J9AYAZ
Kk+oGni4fdCvkAZok8Znyy6eHDHJhkpRI4vks7aKrx4+tldaEkC2K93t28ZsN799iesIplL9Exmj
dBHQr9+WuLsSxhfX+ZTRB+DaE+qT+wo1uBCbQkkUFNsrzEBDSVdR+Fv1Al3hImkmlSjE64YtoI95
jV2UtQRxPoC6kIO6kgKagZNYw1kRCt/rf8eaUV8Vi7dhSxZ7bqP2rqrpxsqA07g1yofFBx4pb/Ql
EV6t8nZJs1RDg58nbQqCUo/0wCcL4B/fpSOF+aB1wBuYkQuPRvXr/tC8LExtYZutOThOwc1EGtVp
GvVQBOmc+i1BVjuHPzTLikOlJAxdbcmWqH/Em52gMPTynG0zZ9kgpHXFn0oALNbvjKbPIP2gSRXq
IxjwsLdbRA7GaHIVbWPELmXU3EWIHecMHfhrQrrPGhqjVQiUs/VgFPtK/KVkX00xTxDwy50Ur+63
l3JD416BWMFjZxqlvFOnJZwXXTNOyb9gPcnm4SIYL9jzhWgz6whOdzQPEMyCNedG2nnsDBo8wcPm
VG0urAW1BLI04gEJMO9DbnfeG4ufAOduEH17dNosYqDpfjFytu9iAXBuArxx82juhwBcaj0a3ROf
ogukQQ0BqxqvhAQeqqbNnJ9+cFl/tDS3K16PRywNmP7V/vSFFoA3B2c9B3g1xg7WdBvrpR8zmu9e
7QGpB6yur99+6UkcYiHD1MFWc7yzdvVYSV50C9Hg7wFrxTO/IGMapisfFo/s+8j+87FeaYtNA2Q6
fQ3hRRbtbSgxBY70o7NcTzF3P9HpSK7CoE3KRRgLzQAtsMAuIKBwp3rjE4AEQS2p2ZI0VZN/wATC
MA12/Rt0QyM4lrv4SGtkBd/q8qtTMzGI6Ip3GR3JNYhfgLk9dtO2dgjC3/tjqOCLkjd4Am9wtkXn
qlGKO0k29jGlO/+VsPQEl94TBf1K//aH5urTejj9cRzv5+7kFSWPpChN6we6IYUMSmbbAtMBDV7s
43Bc3K76O7eN2LMKO8uTLMKbrL/f0s5ZezDS6QKpsDnRfOss+UjOVLUu//ECI77HW0E0vc2WCbwW
t1IFhgUv2UreoDXmiMTgQsPRZwF2bO7qjRpPZrxSyXut9bCtnc0gUhoMtmybd5AAf52LUMX2VAv0
iqJ8/ZOVv4LDbJX1tOIN6pUhAfHQHF3O0wCxvT7jMzS5Dt9YsrzPZdRXgPj3K7QIpIOJdZneVsyw
GMXPrHJPmBa0USHGKd0v3bnhwGFzGJQuZkwuI9rI52qVFi8bcHyLgtPgYivRoNZ+KCUK4bMMTSlj
xfZQ+yDhUWQcpqxCfxUpr39uSGu59wOUWs7VRkT9Nu1qqegY9+lxJLm/IsYRKqN5a7SUIbSnP236
xGN6uTjBbLE3JWOwiwNKF0lJP36PiiqrjO1bv5bg3v8mKx7iyXHmnhPSDODl2ThvUGVAqAB+qaz2
NdCfKTv9Ub+mnQHjWslT5BWtpmC0VpCHqrg3QadjVsdTEohbVe1HEV+886Zg2uTojrvf3XhsgdXF
Yx5hDOJCf3mEvsD0XTQf7PxzRT02m6aYlCYLYPpoipcJbqJlZNcFx2u2rh50UyNcrcIcJT/mudF6
tQ0W9k2Gbj5YllSx3FEx7Cl6FX0b5YiXeRhOKs4+Ey6isBqvhp0QJDRT+GwvmS4GjGG8Mst27Cr1
SJUPNsqrzvKeln1nGzyj9DzAGwK7DnWw+woF3zGZvWH6rzKxktFbujSlHg0JkEAhiXqE3Y54W1WB
TjTucjZ0dyL11LMWg7eg9nbN8AxogXMYNykaNN33+EHolk0X/QAAjB2XkGSGMpN1d/CuH+bTKU4j
uHV2XxAyAy6seXRvgVaSQaxNt4R4hFc4nA062teHwrk+FA7o+dzLsadnjx0nNxUqvliCq5Nyfciu
FLRnVt7TN4pgD7kyEwLn8hFOxvq3BgKUp4yVs2JmAEWGCJc1iHD92u/qAiHRH7s5jIWBjKXXx2mn
9O0V7EMNCkzxWc0r3KRe28FoF6Edfi2d6lGC7PvkjynYfQ9fP1UNOB/l8aWjNbk4lBgft5Vs5nq/
G5OsKOz+R6eDrkTOhMwFszsFrOSBjtF674tWpSziZTiJOzKfd397iim0yGio6GUnNP4Y2WpLaTPK
3jDilZeHI1IYFKaqcsUH1vFkdUzGmf7RSRh72wQMCOqNcpOy3SHjXIYxf8TwXdhODFcYAeum2uM1
qg92nojsVISLpYrp6pBrTOwy0VBqKo85Gm1FLWyQEXYOboiUOfWyyzhl3yvCvN1MvkMGsV5blcqX
8VnjNmuzlK7p5TSI+Ce2++gpCZ2iZbCtzchXnqdtIPzOz97mPuVBeIlBMcfKImVx0/Ffcw4cUE00
Eh90S+GNZDJ464aT9bVo6ZfnG/Zfy1nYHcD0bwBiqS14oRrcuM1LeMHtZzl1mSPe2CZ1S2bnQhPa
g0RoZa6Vtg5mqgYt+SHcoTzxfB+Xr2eKkymoatUSQP/+nXoq30vsNmDA6QnlKSMxou7QpEnGre2f
zfr20mHwxFI4NfBhW/661Q5hlBx3hp6dZ6HsUGlSRYBZCsge/pQ5vNfA36XP88IbD0Rdn4h6ydd7
6Y0CjksQZlN2R4aIrG8Rkg5YZRrZkZNzDpHr3NqcrDp23KcjIKgmjSzeLV7ZnWeJ5v53jOnWilTi
uN6NgrwyoID6UnNAE75kNYjLcvvEEcUN+APDSrntrFbzn4ggRaMAmvBL/MMDx0AW3FhzWByE+sB5
Y/+AtIMaEf6c06agnAD0WgkPTgePlQij3gAAZefN0QixabXwMYDE+/v0pkFxsSTu8zkbAwNly9AU
jyfot2uEQCZpaqcZxvK89j6WqduQJClB0SeUpnxZjJ+hnARh8AUgaW5LMibn+UhHzTg6UCYZ3Dm4
4zy63acoJH53cWEr9zwyW77FItLbX5H6PbssRgSEn+YLxF8VqyJrVakbdodA4jKgiNEvHPNPNay6
OC4RG5OBcqxrYp8/hXC55syikeBuS4A2gbakeMJsSuB3dwqaG/3FatFuYIWNaQ8np077ECeiCCfQ
d0HJuh1UZR+1y4VUc3aHs4j6G2UKfApkiRItVc5P3nN94T0b4mtRyXfZtvEuz8gdua3nuj19W731
7WxouvWM0Y3xXxZ3KDySi+bVo6Tfrf3WN/rrug/T8mKiNkvSc/S5rUONRcbNrbfKoouLfUyJGOmr
veJry1f1wIST+zCEVY0B85K+LfTbstwQ6v0m+Y2ySQOYXo6DQNag6x5Ro8pA9kM4uiz/+Q2S/Vj+
0LmsAAwRz4SdPmqIOh6AJSM1lalZkFA/UYBxN+TP1zTwPfbmmj5G0ZBu07qmQqM3qHUeK+ArYJY6
EzEKh+r8dgpwYREQuVD0qleMcpeEm76azjlUy09qvosFUmUCRwWl08EElGXlRAj55ELXnM4eUoms
/mjur4jwgamdNIawylBNhKXzm3NrPdqBRPpRsmfzxbkszwZDykwhujRXN9KQBKWVkc44InLvXtzf
CTcLI9hVVu7YOk7WK/EIxf2W3fX5rgfFWTJ1jvEQgpYH7dtJQs5z6YqM16Hp/s47lfDqaihx5jlr
qKuIionrdO4NKQ/FhbfGHcbTl5MEqR/o8uBGfsrSOgWjhxhQH+TH4uATcxsDibAbxPqouBN+l9Mz
rovDto3L7L3KdCS0/1IHF2GfcFjJNwMV92R4FxdHLhOcclr1UGVSzuQv4VKDlbOX/KseOXu4laju
F1zAmjzuzW7MMeXcTkK3/Cldhh+2U1D5IC7pqAaA65Duz9R1gjR7gNvsgQIxCEDo998soqEO4Mhf
pHgYJ6C2lYYB02epdeFW/N7EfDbjLiNX90fAEgbjH0MxA9q5tKR1N+NGvZo8kBmRu5DDWevIMhNW
GXzWgH13vbaMy7fLlc0Gj01Tldfic/wITFyufJUbqrQWyhx0dbQK5aI0Vhsh+B+zY36TDih2c4x5
s8jr7rHlltgp+MCRC9xCTtLpBZPbPQG/8zDWB/q4POvim4y3A7nA5UBE6+3NV2h2N+cWMHMYmEgQ
qWKVxScFjxgqkUyNilSSnqrABmW19TcAP4Z9us7x44qRILwXmTQqXaEx6dXTxHkVqva2FEXze7jY
Rcmt7W9eFeU++lSDMBNb4tyN6p6+p/tuZ1XENkbNazZQ8R21oU5cIMD6Wg/GKsCVtohS110F81FG
glvhrHKymuOtPieS4JIyVzeSnU5LWU6wRpK3wfOBPphoIMGpKbwKw6QUqPOeuO5xGOqDpCAZU/aN
Ew3HKlXKa2iFFX+68OtpphSAObT43JHUCCCkixCnRRNg1GKPDBL70vyRSwdAs2H3qEnYMbvt9lBD
LzIFWzfIOTRVjimZMmqZq1KGksyHpzhMUo5hIAELwtQzmlMCIhTLI/BEffmmgvXWI0Ay+frjfqVq
eNqLfe619q3TmvwK5gYDALLEBOi5JJN0eOq5nbBVBZpuCmgfyuLUax/dvM7wT6gdbo8wOwQovYzr
9UcYHM9/Kjv9SiJZ7+ATaybCopNp/fwAFoHzk9u0/IGG4lisNpkpbQyB/tK1WWOkulrNKPXX23QM
RUrrh/xrT5I1aHXaoXW4iZY7EnP1rFYnNTTJvGPbxkXivvHPDv2Q9yFQHjEKVcC9L0JK+epbiXci
jZfCcQBgvRTs4xsZrXTCa1tBj7d2bwRn/O9OVkppD5zDUEX5P3KHrcl5kKxdvmdcA6n9KTcaQr4t
PHLaoL8EdKGAZQwI3WGlpZRjCHMppRIdS1D0EHBNCOHCXpVuDsSQ8l13C0VPEIq6KeT7ZKxS8GXF
CrKo72CewtkE5HiDvNiRL+xm/JCqlIzu9kt1wZsynuoacIrtXnQy2+UCQ65tZG6xTC9A+hy4E96P
0mMTT25fFEwEk9l50ar02XPU1uXzrvJHNiYgcOoicOw81ixxjU4dRMxyzZ9LEApNcZTHyD5RY+C5
hc5SBAg5J4clXR0japHCldHD0WCbLFUKmo3q5r0YEiEZZ5iNF0Bp892lg5J8ytvHkZxQFlBTuLOV
GUyysv5TOr1GjZh7G7rvcnyvw8cxG8A5jMnhiOFAiI3f4qWruV98BNkgR6dmd1HTP7ysVGDmCZ09
axwl0cRuQ3GGQzCgIOirkJevUwHVMfBBZbaDZSR24TBl7EMTo8YCDXuphvRLMmIogNtGVY2FJKzz
hWsKwBjMSdiazzBCmdRFYSBionIzPetODi5eksMA22P37M392ti2FX23L/nZ6pM9fkeEMkQktZdq
/MYKiVWYidpko+V6r8rru1cOOgOEAA8MZK9TagWUD0PKl/RudQr88k7pM4iDoi4PJSpROYZvHzWI
WIXb7Y+07JHtUvHfcxulOGbJFcOdaxqv20xIFgtG9CHYIsiEvbOyI3yCaytiNolcjQDNksvkfFFQ
4KAAADC0eY7aUQ0FxweU/U/hozTIDIyuzk+kaXLJELGouus+ioXbRA8V0t+f7bqcxDM9JtM1DgyB
LK6y2KzMm8au4HeBejDLbzdgFsZuhzz77t6SudypicO48IsJ3VNon9m4jY3yeMpIujLny8UQ9KPf
ZNkhQqABPmHuvE3Z0x0OW4dc6uTkU477w360KCemnQR//ghD90KSZwPghPVNAi9e13iqHaUj8+2A
Wn2wRs+UZzNinY7hkYWh+/A90MHapIwfoxXkep8B5HVYLlxI4U4r47xyU19JPvQiy3FO6K531wY6
RSjTb3U0OqiWsiQ4agJoRDaA67E55t8tPEG+KOn43FgVHjhi+wFN1UeW7w7XKxTPOPjjwmFsMMNm
js9pazxTtF9DdiEB1YTtQMPR9ZoyRB05oFofnbJJHoVjDPP6kXjc1RE2f67wkF/CYonoS3+Gh8qN
h7IGn8wVqM/uzW9XpQRhUAmMNF9UHJPNarME7f9ednSFg9z7rdMleXKtujoWuS2TKsTQlmneuhFI
RD0gmace+QgM5RHikc01Z58H5lslpVg4yKKuXilwCKNBDOlCcLr9/z3fPNYAwQNXQBIVRP/cu9Tp
y6HmrKtmNqMcCKCT/+kQdRUQCujzjYY9hDOOXJki9xjZVNPXYm5rXzt3omMBAX0l/IMW/OBCQb+e
3GvbpCyG0dnoXjyCPixlkO8j3htzz2TD4vOPj1GcXpPJVO3eJoLKMew9ZsdddbnqT8n9ssoYZ29i
L8TIXNnY1kUiLS31pXxs8JySPMpVP2eM811Z9vwRMpUCG61UJck/ty2tjywtK5EKAVZH5nmJt8vZ
Weqqb3YyQF4R38BfwQTEJ2Neb+eQLra0zvOjfwgKYp9E3AV4Z+YNzT8fdkah2C+N/MCwEUNkEYAG
BZKirDjEQAu8vFqIeI6V2VK1ZCM/N2/uiZcBtTAMdu1/KFa4xhnuKYPU3YyFJAZOL/++Z6xba/8J
KMLVoQfZFJDlqMSo2jtazcZxuRi+M4UBj6LeJ8dCy/7wGohAafr42vNo6piojUvOsW/sQ2F4KaFZ
dKrPmSvt4isHXjD5jbJS/c4jEA1GKea3e1g9xckRhxwxmS3FEk7pk7xujwh3kJ686Vjlki4Ud3oq
i6HouPutYuepb+kfjl5b2DcIQZr6tlsNRoTPMZ66H2CPlfm7/mq0VKCQxG+/CSskQw7hRAsROhwx
bI0Z7ShlvJdvXv8Z1pOcyXaoAdXqCA+DjFYEXuOQe2YF0kZohpCR+OU3iWL3/fV/+HLiShXIK8f/
4jOBNXbMoHokK+ZhPYXdkolNBGWhP53CDn254QcczI0i/rfPe1ThnKbvrORy/BWXVDK2fHmrcFFq
kOP0JlmbiiMLI/RJ5zyzywUNwFEoBwl2KC5dGmjGVe+YVaRijz8pmj0lUkwbQktShDU4l658ZBZZ
Z1dLJOmzPG9sEis7WGDXR0OlUAMNSNMM26n2L2tE5nXcQPd2YVCRdkzFrvkFdW3o7iBGYKglLnVA
ECWVZu7mwocUYkWv8jso8xAekYUEBpgNutRk+Ken2AXPiA0FXQgpE0Y0R3fMUp9Lrs3znA39IlU9
KHG6ppRS3NKhVmufN54qL699pf4cdEdRg8P4FZ9uIbOKKTkf9KtCYh2HXjAHxklD1vng2NHV2Y1p
S/H+mQupUBsV5yPeJxTUyW5rKVPRpZyut7ZmezoUYL01JrVohvz04CCjxDRy5oLCOlYWOZ7mND2c
3ny/+zQmfibrI0xCusrqNMmRwsa6y2UxZML5aUa37eV5+Xk8EUJgrMdzYF83y+rAOWNsvvPywWoL
5ZYMlsreMMaqqRumTHgWQE3yj8sx89otAIFxWG0AK/Nei7re0fCsyYMr7oGtGCDVIrNt76sVEKGi
E1O5mmXmQk2MBJs5TqAL+jSdSaSqMNWZCfdh9DirVQJp32XL5XXiHjpOPeqfYIK8Wq8qjcgsY0gT
jU5hpHvcI/mto4siSaAC1Si8bQE2JAv5uxyOfm1sBFLuxFimq5tKywsu08m/xtSTmeoLW3FLpkRr
ctqqBYBPGCFTOpGWM4b+CHY76CWC4mDTLC1zIh1E6nOj+cu3Uo2cEmdrFEa7bywpf3grJF5sdt3U
oFwdUcsAa1lzCzisbRhOj1UqN4UlTWS+LRuovjoamGB/6rZZokPPWe1l7vK6MaVWm7Vq6N2kNkR1
wKUsatoATU1AgNsANOlD1nt5xiNILkDXSG+nnsPdDsw766d9mBxdKnU/WcEvEG4P/87ToLiTZcTK
xyLL5TZgbvjy99k7OT13pjE1uvTsf1n+wqKyRMo5Nen/vDa0upCTq4Klf4jVqeMUJ2BoCOO+7Iui
+K+vOl3Gu5vjsKNSAGiER6X+OIsIFkvR6HzMDOhbz7e4uAr+SfuhXu848hZ8LViDofCrjBW/IBTq
mcp0p90LUAIkx7hOyTqVPKJJ0YE1ya7HCn0KIil/gKuzyJUDJ5LV5oArKLECPlotcW+NtqKMVjZg
+KfMDD6rGRNJjpeTOILaJd5GqQPrvu8XZMsg7xgFgRbLYpL2Zq3q7Tg9XLJRkKzqreovanVmNUim
SYfi/ZnafM0pFVQB8xeIW2hb22WMVaK07Gqgh+UujZ4/4BnA9lt+jJqvWZ5FU3fZIijtMH5z9nuv
+R1DaO1Gyh/VSt/IuT1KjGJZ9Ogs84PF+DSJUDXMUhQaVug1CNwBISHNVmwQGw2OAz3gFvDS8ziq
4EBRK1EeshkXwR9QlW2D6Lh7V4lul5pN7IJ5Ypncev3kkX/Nmobr36NosBHDmuq3RQ1jFfxWqC5Z
u6oem/viwaBCW2dbjrZIGgHVumf7msF0XZhhnDI7xqF/y45/PCny8vJ4bKSg2b29N28aFl7ofmkG
5xNUz6tNxnNlovu7c8e/4FJ4DIsmsGpJZbhVAY1CBqw5Wx+1YDufFvlCAy5o7WDn2edmtzMLPFTP
xkD3h90f4/QDECLY+dwQ5aoBq/9yYfHqQwaPCdb8htD78H04M+4pw6cMBaqEQya6Vf+WOhYnnj9G
M0JtJ1257u+A9k0OQCgLMSrwMKI1d7LICzms48icLI5ibL/8y3q07Oqk2w7tU1SjNzu+iyJaQyDz
bBE8k6tNRjzjWzVB87ajRJxTn74QFj5P3ckamtXTC835vQhq0zEwaYqqr30FSZH3GWm/6brwTZYL
Zs60m5/416g+PYxN5SzSwZn2unk1GpKaVyFlEgZ41q7vODo1ANOa8+Iz2OhiXyE/yySuADm1x9zC
RRazUBqO0KAtlcWWgMQ9CIttQ8WBu8Ccwdw4wOKv0ftfBunTZBYv9baaJY6+JXyIXdIb1he7LVAr
7lTTjyvshY/tazc/AeQe7Nqco93ACbtJOT3a6IiHjmW//rFWnd9v0jGbl7LDJMLVBShVR8lvucTP
QqV5ep2skhJ835D/z4lO6J9MNCFT6eX0kwIfu3A1BAZ9ZzA9V59rJ4q9VsdKy31lhrP97QEq05bc
kSrTziJfQjRh8IowOSzdcbuYkJxU41/sdI7aihM3U/ii2jNTE9bANdTS6lCtlnHIe5gW3VMZoOuN
fTsc7J49vqnBy38kroLEvESa3a4B13qmEMLiu0+dNgnBe3ZV2phOpS62ztXZl6NC0SIq+UU4GtY0
tvvdjuJCjy9ltn0hRWPVUk/aDlZ7PAanXEpEa1FJY/gLYK9yWj8XQbGcOzQ5RSNJI2duwtS/uzzY
7q1s4XO6OoOHK6xxcI8k/8NPWQ645T/+UrfXWRkDU6O/3Xb3Kd8rWhytub2L5/obHU63dRzwzxkM
C9yCTT+bStobyMh+xjXy6KC8/4dT4BLKtl88pB/OkybFcrSIKf/UFRsdHXBoIX0w4hCeNr6SYppW
YTQFxux9DkQ57kFyc+190BLgTrZkO/jMWvA83EPUr20XILHBn8Ww4JxTSvFFiRAUlZNxyFDMN+BW
Tiij6YMFoEl46il5RY0mP18HsOpsspyNyYI8H/BaJ5XlWInDOL/o+mz0BVCARFg2rmP28Fgsdpll
I3u3wpc18VEedTIrgpQLXq3U+/BqDO8O63+6FC4wm1UMzfx3pS64arJ71Bq/OZSOPxUHUyvfPv62
m1jGyDLK8Pu/rFOuqo4ruf9bpyZ+00hq2X+W/diaAJH7XyTft2DzMTKQllPSun5IZZ+hgH6T+vVz
1B+33DhUYQ5dsnlrWsfgi9dQZWKQG+HRMCeXvbqkM8wf8EG5lbEyCBYgv0SGjmYeU7g4e1QCkRlA
DQpe7qprX+mKyKzK6FYMwNWxEvoGy6SHT/C17/TkWB81NX10rGFnhYyBck2fvgachlaLl/BXJrnH
YtlGAcTwUBss9+0AdO+qmpwo89Nk9wK2POEQTn649JtpK9bhhekFlXDGQDiRuLUwmiz//2ibaD6G
EB0RdtduYKLe+2B7KzTf4UAfWykT+eVirQ0eT01TuTSpr9Y+0VGhvqkj7s10gHxo9wir843ydJBc
77QDZXHv7cYOonb7qk1Ft9qV7hL44MYqiWJ3bA6kVV6EW2Magxq1OmsqWHK2e9thdOgYq4s3o7U2
NLcXHHNwVoSxQlG3F3LDgoPMaoLVoj0EfhnAqdjkyl9bIeEv9/rjPUR3lRar9Sn8ZFylmaTRx3mj
25VLxEG5Zyykfi/OSSvFcFwIi3O/HMkrIGyYE8ceXGQTB+C4yXh2/8pj91G+DKFqpwj6ZkLsdP7Q
YRsgPKuavTMdnpFWBpo33WPMMaGVL/LJ/aLPxIV2HYslRMFiJs/Wzx+SG1TU6SBKFUTdfKiSrFu9
ero2sLjHJywfoGshH2UflsoD+tdPeKpXRCaMp2Ibk/z7akfUMjP2ptKne6UgONxb24Fosb4mek8V
4Cgjdh2tT1knOF3+q6X2X7dSn18+PS97r7qyCs3frLLqwJjiD4ojkrHeUFQ28N+d2ML/92HwbAkh
va7JN+f952Hli9IciNDhj3zfBKHed7I887QNOyH41ZjK7R8fr7R95aF7bXk5InucClpCxz+DxYad
dsmMHWqyQW56b2oAIGCHmcWfoIU9wh4eStCQY9kj+fTh5wromSMWPqtOmPX0QBAkdfc0xf11YjB9
y+pXIYKe0btDrqJkKlHoaRQwgfx+JHom7x5F2wxBnaUK4cS3M1FuF7twpzZzyZQulP/uhNcuw47Q
EO7aXLVaZfMFGTdlnekwpDHH+rKCbUAGQYZkoH7LDAranGHmLU/gXfgLBhMu9jEHTBroB+jB0OJc
MUl5jPaSl5OW8NTPDSsvLlQIRcSAHuPnWxkQorlfaFqY4TZS4khwCt+h/76ij0EfNkCLKXPnKiT2
UFALtSzVLLZx/JjB6fwSYwazAl9Ayu05YbbDaNadhLS4U3b/Ye8OJpw38bv+rlti7rCbno1qx5Et
fkJ0j1IghTwTaAqsdXfiFXBFQuK05Sf6+OAhQpMAwfT0s0vlu8QjmNaqdZbK9Xcu/tHH6LHervEe
F46SLByfB/GrR5LjLznfs2G16uwqc7nFjRmgkfkuzmqZiECqS/hcTAQsl+jrcLCSAKGL+wywTpzE
4Do8f0C12tMd3Uw74c2A2KRxc8Qb7yKrW1qwH3VmBzR/HOqR3er8rm7uFM9oh8Do7QT3W0Y/N3k2
5DFAFNJSMNN+XpRbCR9kmi31GimBicabTkagcwwOyZl8EjqtEVL1ewjsAWuC6uG8C73ICUFDNC/t
ppFw/u00webe+Y04cx3f1AC65xHJh1Su9SI/RsS/YmdhvEGQH73aNw38Zhsn3wXDmNlV3Szlu+Wx
Nt5gnGUi4eHBBtSFL9nrUnmPo21cgj9jkMHo5+arl2wLSercJDGls4zJmpDp45cOnNoSzRStlFo3
qZlqmzixMpCNN/rYXhwa2t5SAYD9tkn91DDIDzXNzzngAz6419HFiBp7WPIPavKIsHQGPBgKTYA5
lb53R82Bfrr1hQ98Hz+9S3p9FidWhjD+cwkp+enaY+GhiWoWD7kj97REKKHleg63T8jpXL4UWrgD
mik78sdATNcJNlMeDGDCjanab/rM5zX/cU/ewHPxEnUIObZky2FNeZNiucHEadKPo1exSwNGxWtK
xJsS0Fpir9sXssniKiB9CKiBzeGA1L6BaAlsleDvjwJtV4K250uznWQ7EY99st75sxUhN9U2y2bk
5batWynedXD0U0y+qbVQSEzi3jnyz1/0c+Kw72Rp9qjGUqF1IwmkxuGOu/OI306zKHQIyyKKyGUF
hyWDAUvf3HQXCyKCcdm4rWmRFdoMSgmj9Kd1vT/LtwXh53lBBQnKKLWpC9pNGYWVp22xoUb+1w+Z
nzIanNgp3aibVwBNEQpoAPYy6N01A9x+dgfRyLsSTd/xRDYkYGhBP6iQpoFH3NNSBwzI7PlTjbkr
wpCg7EH/o25uVYLgXR3090T9olGli164s2ip8abh3Gkia2sew6NcC4dXIl/6Ypy1NaunWToSRVAl
2t5B8PqcldpHO+OlnqiowgJzh4RhJ/TdOtHDm7Hhcn6apc3HKvNnUTHTn95iGxEeMqs0NuAbIaVL
LYKrFWFui83rJCMhCufd5Y3WBeDRaCTDIA2qgcPxiiKKsBrEw5bREeuYDvr/18cB8nlWze4pIaTA
coO0lXctT6xZcIUhQUwobb57L6uJvLPF8R0tBQTlD/NtGL+UojwnmN65lUbVz//vIDfYRWg11btW
3qJbqhaC4CYwAZ+Vwpg9lMqhZlhqK3Mr0QUN5ZBrz4aTcQlNmHu92XpFar16PQAkG7yT48bBX4V9
mWE3WlWZvPdLEnFQs9EvayKeW9vmTDP402VUp6WniMNdQQniGXYQTFUigH4JEFIqq0I1EFr5vbdk
gjh44iczo6w77YQwo5VP+S+g7c44h5acSoLqrCkVH+HxE2xhzCn/6um3lcFBvcYY4mghkFWVsyC8
/JOEQ/O1221tJk69yZ/ts2HjKCFZ7IdXKY5HAFDnJU44EikmM5eaSi4gn5g9/Mc2QGBS04XI2PKG
ZCwka1O2xi1gB5ZFPweEM6lI/ttsCVE7WW77kSV04lzFPzJSE1mk29tN+kkXdd8F9reXqRoCHxoj
K4fcZbI5fg0mbyDhHJ3uP1DHeYF8A8bk7j0JpbpgzEGJRJez4wzAU04HrSdgjlx2ytu+dNDDippj
gsC7jUI/SA6gwC+1RdYNEl4iTnuvEcIW6vBMFDmVPZj1o6M36gcE/uQ5AuvGvYr0DxClW1TXxX3i
1Fv5p1ay+uKbxV7i5u0QoXGx3RM/I1R9RBdIzBYfHVigXknxldtqNeoCieDYuJbe4WkaLMZ8C6Pk
QYqqnYdIHFkOMvgbGyS6gh52gHjobhV8YbDoFhiwCSi166y45+BnF1JWHPraw6QXBfqgIKTz7uPN
dyY2HhD7rLjOXZH5CyXhmKjJC1oPhzEKOtvP0GYG1ESxUqhSEkDCIUyNVZuOmUlv8sZEqVemC2O1
2GsJm25JrtsoUjK//zXi7b+rFrKDpO5tD03IlMXPg48tJ/pPl09Sw72JQ20L1CBCIlg4ipeiveuB
jEj8/pGLpvSCYoRf7H+rFCF2fvRitbnQmI/3bG82Nu1zT3SsnWr7usHRrTvG9wf9yEjtc+dre4QB
FN1C/+OhHAZEL8fUUOaT9AOi2LgNzbKMJhkrYZ8Zb8PYjYq0nEuhmgLO/fsAxukXOYR8Gz/Qc9f6
clvvbIAwCsu2uL1VqIyGRBMJtxGPebT28rUfn0y5Sy3GWUCm8WYjpwYw271zaXgcJ+WSdtT17CGF
mxlN8V4rRWG72PdPHx86DkFNGNPHcHidPc8UyR8uJU6m37A74jYg75QaVefl3rkzW5qZ8VSgcqk0
yoxTjDtVVFfVVIIR+Xoh6NQHAVgj0fiP83zhILdDauYmE44GDN4oCv37cc7GVNP7ucuBYTGV5vJ3
rBsuQ0L/EYpC+CK9IoyQuAQ5Y5CB+9PQkxsVXxvRsGp5CdHwZb6gLHrQdw+H4PAeN71aCamexeO7
BOThbtodcVdiQFSDFGOiTUB0KobUBKuqvJD30UlXmFLIu+2wQUMQWT531fPCqJ+YQmeIP9TgXp2V
pCwc7TlBuVV8VJu6WT6n15h/tzKTUW7GtxyiYhz/EmDL8CqHkvmkZ8mGUlpASQH+sibiOlcaHsqc
MxKcoGNxBOUDe2kh2axUkWNyc/wjpZaybOude5bzgR9dKE+4V43ShqU5Ql/2o/WfiS5P74bqrO7g
4PsMZFhHYIOabpesLUEJUY8c28zj0LXN9gyNfRBytLjsHt4hdxqSn4apZDIz00MB5oVStTiXOPSL
FH17qZjSQq0U/65/m9fDzcQEbLQ8XJrUr9ScdpLbqFj2u4+2lkguODpXmVkAtgwECm5WAFf+lHeA
ujFuYswLjc1myVujwUM+UI0ctiyQiF5S2d26xeoJ1G88YwrnZXXraclXzbMQvQteQ1TqLW610/ms
WXJILmXEVGTYW/jGUZsGAlk4/UyM3lESQWrMMw+fMCk+D4jRRhyijDk3NGkFYYDCMQHmiwxqBb1h
vMwPsZz4tPmsmkF4AvhQ7DNuOAxfysUfXj7xq0udurt+tCoFqG/CDSdrqgjdlD/EgTh7QUhyZPsQ
7Ey5xh7xLLXqNv2EMDXyPIBwNa89Dq59KZIJBrmrQfuk5ZAgfw6C8I5jEEOf6SSJZVqQW03Ow4Vn
20jKIHSXUrgj7i3nFvcDDfdl2Luy0eDwx5Gzv0piEHw3w+CHRipqCTxMK9YTH6OkCexhmQ8dAsXI
vkCMOFrby/dbQRxxmQDLBaf7yEkJVBVzpECyJyGgf68ZSTY4USx3zDqB1FUIYL10TjUDag1NnsOS
1R3KAsEVbI0Vo/BDvZHRVmdfNMmS71Eal5R0y65UbaZ1nB5mtgZrX4mw2JG35qy/XHNWytYSThAn
lrKdeEzs3WFDBHQ0Ck+Q4h6DclCCbwCdeuP7vAvuTwCOxQ29BH8UDAWzJ0rA2xrKDXc0vkAro1nH
v91EFL3sSl5JllcNHs/w9/Bcji/6Vv8U3nuOZYnOomjAjlQXDYck6XjgFRw0LSaq43QidDybl7p2
pbYuYgeCvNYcyqWeOerEzk1bkv2HcjEZU7nU5e0QGB3904jP8ViTFHR6bw0jtoqeTcm5qODlMU2/
NcHvxHhIWOB+4iThgb6O8/MAGGSVpKSkWQ1hDUq4so+R2VidCY+YgdzQisqS4lQMV4gjN6wvnTou
mE2R6IvwDOgaIfwNPyWHaxBf3grQy3Ks5XSvyS1dazt3y0DokG0brSe8QawHCd6l8YXnC7wsi+qs
L6FAYP8jVOXu5vqZv3TLFZjT/ZCadXvYrQfA6tb2JBNsNhwFPXsCI8bKef1JE/acYhBR9Wx7TGlf
wkm53piMfow6xeKBwGXy6czERCsY4GktUB0bfQS4XMFd+MgEO/va97HSCUi8R/+T2qgvTDIMn6qF
mchH1N9EjNzpzk0Sljgmu6D17nEYZyc0kU7OT2kOJT8Sb9SAGuphfuJGosx+G0hlZavoYf6n0Hm4
wxwx+Oi/7vg4rLxSPa/2UHjkiwLoe5XZYnTe+0Ntswa3XqH3lkUbZA7h1QX6obD8zNI2BLISEbf5
2OpDoALRsZnHY7dwpLeUN0sWytwx7VZp0goqLKTUUG6SyCcj7Z1PL5RXvcVfm0FiYc6VwCoJL4vR
3QNPFOw7pPwFXEgXfnzIUKQd2JUT6opxvctJtu/qn+wJDM8W/Vlso4s+dcNPzL1G4k5FThTlXMI9
WgKFSB0TR1jzcSg9sADzoNcEtFIYKWLpMkYeHxaYCJ7tS8wY5c2F0KaH3kRl1HqBYTy/hNCpCU6B
mQdaT6CLBcLUBWISDPzL71XxTCnYAltLDP/Y/z2FvNXyGFI1LW8cagIUU7f+QP1lqeEkps2y8QVe
04y+yZkEW3hgLKZZdZzqHkdoZqGsVpWUA4Dlwn+r7JxoKF51VdMbk67Vx47uByJIu3qkf9stfByU
0ZUtWxN5Yvq9z+73qPYyJ6WITXO4EJPOBxneHR63htdKrAOnHFqE3e0idhsxXtdkvUmFarn87zA4
hgAA59lOKCcAvaCTGq1lA7Wm/B4M08v5Jzih87lEXDs0j08cwhPEeH2byuHpS1W3itltJZCFLaat
a/fWHCEMIu328hld5kJIzM0zyvVCS+iHLTCTrUfuaMuSSNHeiRgtKfd2yXnGOUlBhUqXaFtsCYIP
GZvNNlg0IkF+2SY/nlOTEe7IYyG+x8NqB56Hg7GtW+89xb9Th+kxiZvQwWiXaoE/kSfMRhXcrTYN
YOfyUg1xjITmbhGnE6hLEPsiNU9qjnnEaTn4Ga2W8x3XfsFFXRdjyzlSaV0Pda+tXws0qw6UHA/n
qu4gtmVZqFDpv27OQK7EGTG1nzZ8cu0pmkBiXD8EqoMRCz8jfdqsHWq/s5fGr0PrsJzwPRzCpPLL
smgXlnxNGybEFP91SMc96I1fKT3ipAEFIwHA16qOhbmjKwZC5kQdIszzDrQ+5ZDSfRHECz/1khH2
74VXuNLhYtFffItSJag7/9UDzlWlq0dgZLApjHaM1zruUIFikRO6ToaTD2vhNKfkNBGllyU3YBP2
egeVNM60UpnN+ZZ6n2L9wJun44wpIwmzyNEB+e9Y1IcealGkfDDGk9NePSKXXmEvBb2NHsqXx/E8
24REeP+EwcEojjlaTwi3KHmwVgKZ/THaTcbE2AWz/rEK0LLEm0TiTSYoqatK7iDvEYt9OV5sVUCE
2CikWsfDKgA9labYE+hj0K574iI6UTnPanShpYvDOHhKp4drXZaZuGP1f0JBjgYUAp+KwmH4i4wj
kwhjSW5gHLaDg8ZsBVK73Ta7Cz5h899AEyqz74DXUDHjfFhg0m9aQw0qMjE6pF4/McNuuwwsX9C/
M0rwgabR440keYNy0YDS3M09Im2+FjUZQAQ/4YoorLlIjbsZ34TlSptvTjpiX8fwW+6cO0OIXYe+
xjNYzdQkumTahGVOCTSnyZ3p313S8a43/TeDI7DJWy4nXW2c19qovjtpeKMiUUYh2GMOikuucikZ
WyQ1eYuJEVVGVgY6t0zsTMwX8jvKBMUX92tjw0LKbsPWpdqMux0D3Cn8mWqfTaoppcZ/GGKkrDGK
70YgfYYswEuXF+7dStDyIjVhqx1ixgmBH3wU3snqolljb+d/Tb35j2Att81Qqof+dXS/pyCKgtoy
nztjeggnxx3gytYU2l6p4ABmaOxN+muw26RcUaBkmLqB7A4yCV8tR9QcClBqr4ekmZK2+bL8tviN
LS6DUvCpzW74hUOXx6dIiSOoQmJNC2vST144O1Z1Ki/raq5oHR3irOrlbrJvTY9bMzhKE9J0M3kS
qIgMqBkvGW8UkduexzUuTuZ1yzqfzwdUHDfXcmcyM8vR7Qh264FyPddrPBF+bVD3kVzuOF6fFxCi
U4pWrg6fRy+r7fEkr8tsuhz8GTHNVkG2aR2IXErAjBN865DdW2IhibY8LQcdjcbByj0ayw7JaZj4
i04vXaIdiVtnO0OUfVf9NoQTYpMsTd6dCWiKrpq2wPkNg7aeA/yGwrdmvd3cbJ9UB8J1uWZR/n7w
MDnz8+uYxG3EkPg0vNXzqClt6SflEPGC4nX4KTegWpxTCCnskcDAoPyEB1IB2uVAhPZGYNRGmMtK
0pQoNyNupakVRxzRb6UjocN2aSphRqedPP+0i6Je6YgF2TtQjc7JpdcRUiTykIo/BDpOFK3BORHj
PXickbYxan+cn1lSgG1HxBHppNwk9Dyxt4qkhAwydvSfxAhBXfZQzrBssN5QcmCnbamg8y9cHiKm
pHUpz47uWtjdAN1GyNciLWldOOILia0PB7rVb4+LP8w1QziJGLZ0QQ6cnZ1zxe65OMBT7LOjvw/Z
Ps1II0h9FWHUFsLAaAeRrEDuEFAu4VOG6zW9KGexqa6L45Qo6mry0XdNPJziXgk0pf7d87S514QZ
LSufEKZUnfTdhXFNXiwquP4/FEnVplS30tiHXUtFNJSXrBrwYEZW+Cg/7zPqvepzz1TRZJEaPT3h
QBbYHziHN1EYyhwF3OrXjWbRRJM6HV5CMbyDAlbH5HRBU3tV0oVOilL977xDH7wFam0pOzLTYLe4
45Y98xmpjFH1eHPQ5ENC/ccSpu9dAV3MfIgLdFOY/q3NnWjMCuLErEzeCQKoe6w9rAGtOpZK3UfZ
0X34VZ/9oI6WBZetCZ097PZMhM8LtRkX/DTPt+fOyrNl77J2kfXJ+gOdEE53IMc7bhO3RNGpWyoc
+vE2ZMIhioJTErb5P3MEIV8TNj9EoHqrZToL3mfv2yA+A+AAZe29QIjFyTnocpKKut8ySMu3TBjE
EQmqUoC6gOZaQH/GXzY/N3xu18u2Sp3+7oYrtc4typojOlAcEDKNkB0Tf6RLrdYvB2sVHcrNUHmo
Xvam0ZUGM9hB/F9vcPB3dWOhv5hWAYWcSqP0nExcvV55YI/BGowZ1MJdvLnsQEOpbFyoBOEviazA
+Uicnhn8klbPdR7kn2+waeCm1KtOd2CPQt5/bXG7eeU7UuupNH0V2K8rMKddGnZiuBDcP493hmnn
/1uzmZaBRPlxF0Etr7FOn+GVcM/fa3Mm/xBqMSs0KmmJJvX7GeF2xeHpHL/Ug7ATvxl0D0WcoiQF
gb4N5bWxcJgVhZE1g0US10UoxeEQvU6GkoCzvyBL//OOu7KZ8ciR1eRxUU7Nw03KO1D98PmeC3yi
YQrvQS3/S1Xr0np7ybK73FnNIoNZ/kJUPrm352AH6uWQMEU1pj53H7nVVb9ITTaTW29+MjYEXm8i
5CzKw3N8yLYgIyfbBPT+auO3uPh752ct7LtfeIdZm3z0QSJt/wZ5/6PZP1JSRNseKXrnG7pk+DkH
g3JMnBzpDhTcTvYzuAKRL46kqDB0F2NJgpDsrFj+NPgIVr8KJqvuwn4+0zooZXuPCZkVbRvEVwdV
pKMTFyFRsLY2zM31O/K3As3AS3NIuRTboaQlbXBovDQSAp/ccwVXdWM399k42m47H+/SUHebbXrI
b15WLDejwnwnHWJYkUUUstf+S7BMKbzgGAn3fJikW3pwpQmj/8Bdo8IVC98l69PHCo6v7s8ZsOFf
eLiw9vpJVWDqQto8GUvtxAUSg/mUWGaaxSl0HJ5jBA6NNtfPKzk/g8sY65gpgITU0MJaXpKM9CP8
N+gde3x1U++a1yMcVcRWF7YYyLIo0Jv98G/rwx9WIDkstyBErL60eQGDk2BgwMbLF0NxxcIUt3HP
/p3DIFBejOCoaZI00H+Zi1CG8KXNkizTBjenUJGFw2eMZVe2EdawZIAIi0ChXUKZxmETeuN7woQi
GuI0o77PqdZWl3IJjX7nw2I+mttoHsQ8UsASkzbM4FUOB16M+qTocZQJt4AnsSagHIGOD/IUMUGG
tzEtG5euPjylAzLXFtGxuI07uVAOl6RrGg8ZyJTAACuQGWT18Q2EZDw/9H5ZcRRSSVHbkfqhowBA
eY1SCAfa/q6Ujh5WLkHRUsmu7kCnB8Kv0gVwlI8yg6veDVChHamEGDmKM6XuzMdBhJFfjFg6JS6y
ztHJv7HHKBzXNxYRdmyrs8A4yePJB39Xhk6I3/4hdGWmVIjuz6SX207FUR3kuyHN9PyxVSOR1sX/
Zmk+MCcRWelbCTZm6BpTCa2KZ4tCRF0kaMo1wmDBrf9KY191ZlqGaNqc+aNFh+jsQYZYirYpaY6H
Qy1rR2OzlVR/tr1KhYciZNr+dpcojxyn5fGFfwUZ2f3jxF4xE9ecxhMYprPD89d0YMRZRqAxYGCK
hFwhqPcyP5fP4nB/pMNVVGcFuoxib/t5UIk3FtUK4QKhlsLk+j8YxsUfb9rftib39el/MzdHw4zp
nahAIjlyjLTHO6IRa2zyarpFAovyYbIQHiX1pMSlE9uNo3FIRvZA6nYpoTrcqfcLvGPsHuv0/Wez
CpptbusIO4hbu7BjypGQ+KwV4PQRHOuEXphdkPN5Svmks1wACK6ymDaeR3Vmc0cEkAn6pg2iQnKs
/XJpAwRyUpoliK473Ixf0eloHSQeXm9WIK7aIEg/hAKu9EYLqa1u/iaQHPh/5iu7RJnWxsq/bBQn
v72avdzgNE5MJ9o+enosS7bxIaG89Z1X2V7UBE1egiLNIJG3ZixI4vhoIOLRwcGskBnQbTZoFgu7
ItaQb9rmCvfSbxyarFMnCfe+8Yvo3D2/aatjF4Lw6nC4OIqWYO7s0+Mj4ZWz+68nh4Bu+Zf1Zy0l
w1y7dPbIcmNjoBZzSGHUSaAxY5pfe7uClwE659dTnerAwgqDSUGBmJn7ni2vv+h6U3Drb6uvBifE
N4NJbb1/QBwzspqHXhXfFP0Bu6SGPbiCOH1QDm/5xMICQak7sp1N2NLQ8nlvEvyyJ1NC1ZnH2cPN
H7rN9Y4A2Y9Rw8Pc2ZWzIRMuN2Jz87Ls5lNSYZ+c4FvyY9jPDJbn7zn/FLuJ+xgLNg1OVWINSfZl
ha8huMjk8wH6/StFSqMZEMqWh4si9BveX0Pv1eICopc8HNP3nZwWa8DomVw6H0vXnEoMhSCCW066
KprKGty8VUkjQg7tfgisxwRbdMPcRqJbpvsy4swrSlPHkAxp5hqUmTY4v0+uDUgeBNOoWAAAW927
cssPpX5QV7lLP2aZMDz4wXG5C0XahS1198718S9PBXQlTBa9//m5DdFy6UjwTTg45PcOD2NQm6ow
TFDOrpSTgPgAg5VcNZ4XNoFGobeXadH33bSTOuB4EWZd3ljiCLDnimpOXsyUriuLXt+gCNrvqmut
L9/4t2YPny1GW/IhDl3jH1/tNHD322e2KB/TNneVfDOe1R8kEmCoAs7rL4183ORMEyKD43NUssiJ
m/Sql7dr9S/BVuTzC/io6B1CanJVcjl7hnkUVXNc1ECBeRMznWRplHAFerJlOsKL+m4AdjwRLEzr
caIjkvoJNc52cwOeuzTOXs1e/8P84cAvT+4IDw0FjIdaGHfX8c5EhMpj1YfFJfSwiqsIOfHXl8q9
uhEjKDnVwCO4Xv1U7x6U5EamKdC+U7LIcDIoOWQESKgJUEG5rLVv+/39Cq9GCAO9PXOuRKnXCdL9
bUGFH1JZEapQWUhu/HVDqyVopxaXNW831Qh+7UkH5a9DjgJH63qQGkfahu6VdPerFO3yYzNHjDRO
uyPeQgy7pjjPLd51CALakir3/cabKJ+KJSdXCw793t5w8rqB6HbMUGPfF7LRcoaJiddHUTZYARB8
FTBTLvjEVUtQ8UVkyhtkcrdcX1qx6SgTSgHZLzWYt8CX+LcdO/uE9bqoxZ3EBUNEuiBXujZvyYbZ
i34Z9LKVLD2ffTHzelx1ya/Psa3ay7Es6Ra55dC1nxT8B/r6gSQV6coJYuus0hfm0Iut2up+Fx/f
AkuB7h2ks3+m0xjP13wi2Q2IukVxNLS5F8bGmyak7yr83zEptI1Vf0eOsbpef7sDCsjPP/XDJXFb
ekymD6cPu6Eq03KL6nO8w9SvY6fomD7u3Eg4SsWJ4FY9U7fvWWfO82eg+nT4VIhYgW3ki/Jd6SyX
WotPBixHlmrFzjs5+mdojPbCPWlJIEKuSCllXcJcLpDxSbMM1p2E5gN5bGIS/6m3vE5WC1XOxBdf
ddwwuWan5O+bJKURWgAM4JVJlz1BDh7gtOmhr3sovKN5t/ilItsHxfsZxEq9HBGgq4+bT5iKPmI+
WtSgaF0eX7TfQHegGBXGlXXSJKfjoF3hCfSkyqP0wlycPl1Z1YmbYt3z9J3d6zRGwNubLYykQUiR
NPLh+b2+OrMJwYcF6jxnhtgZsACYjqBJUPmYRs9EHIkEBwGELKS8/5z0Zqz/+IDf2cvY4OLMHdao
V9Q/tDGrO64/wVepR3ojIejMvJRKBjrJAwXJnXM8BHWRTZgML39ZUSVX81HJDdKtaxDf2gLNbUMV
Uu8yUURl9G2RePj54bwN/N0bFHKDUU/WLsHH+UqfgTM8s5tQKPW1Jr2SiZ/bwj3Bhg/2XpIPe45R
VYRDt7DKn/zYhxtcXs6p4m1G4qffJsgLl4AZ2MnxecJTMPPovbsUHNILwDZHUEfhtjnmUOySXwEn
9jrA71DScyNPIebvsNZNiDZflkQFIYI4e5U7BxfNQj4o430Typ/3c44c08uwGsBycsJ0DvgAAgsT
sDHKC5ul+gcPNo1jTWFwDWQxUiXhngzFuWMFU+XKwuzN6Tf5qjyOxDVdDhqPnftZpCvIKzlxyHQH
dDuBv4mWcFPWrtOdxQakoSVmDItdW4qd+Feul/4H33LsNUp3w/I7mxS5tSxMN8sgxktfQmgfGIft
nWSuVxoqmLutMbpJskv8LXZdsoV0NSvrwTPZJRY3LGNtALeOFbfOiftWB9rRwoS0BAnrVKnwS64l
+5wLyKaTaVq/YnwDQeatKFtWtczwcUg+BQj+eLwOKrSivqzoOxYmD9NKOCzQaeSs6ar7pvHXZRyB
br0ZL8kzw0QLoKUXJJZnMXkkG0lNqyWTbxf0MP4FUla8wW/Oh/M+HWvCMIxMfwsw3ovIIoQet2UD
QHrX79LgruiiBE2VUQ9SRCUoMN80DLvsEA5GZNiAq4+wYZS5Z862V76C97MjYITjoQWbk32arvg1
cbqqnZmVreROw4WAg8hG4xHT2otXpgww003x9F/LNvuXMEq4rtPYZc+IZZDJ405cqXJNBXd0Ijd7
iSeYeDAn2q8fKEHEh+QIcOv1bNvVaFpYdtGVa2Bx4QzIFmDtIHzc8TC37V2gvcu2ZAq5HuvswbFX
yKwyfUNICCZoTaHHXzq28wceDKnJRTAVNC+0t9BQZKvqn0V+S7oPpHnjL8dfbxtPWq4+xq/QAPfw
cAYFT9rYuqb472MlludADZTDX/cA7Fh0yY24Jy+FDLQXcIEK4estPL6xbI7D3gRVZP2J+/YlgAHN
DuxrOJsj7Vgq4LhODDhUnxDW2v7WchLbtnAzS1hy+JTSl7iMcNEqNi7BqhQ1QxG//+b/PM+x9MWM
j+8JqHxXf4vTzEmUBvVoQ5DV/0W//GronaCZ1rF/ERLbGc7MDK+IK3Sih6qckW/KhLO4/O7xWCML
w8XPM+n3xjPH3ZZVd+uBGoNs1Vlvruj8LCfBTa9ZkEw6xW3kLImpfXiIEh4hiv+KcQDIvmawC/Og
ILYN2RymWZcOkwHmAVN8CFKQQanIBWu19xASC4bDASflCHID+2dPUfw8aCl5v5xA0BAEILWz7vIc
LQcgdkcvvfGAcTeLDUXIJTDPAmN/DEkzM+mOcpFOkWcdl8AMWbMA0mkiIqs2geyPSO0m/5fCG5s3
C6KPoIPcS9ududHIUW0trfiuB85hSyZt+x4gqqxAZke3vM+xm9CEnu4n2+RM0kLtuxIHyPoCH3a8
IHrFrzZRBTDL91vtDoo8Qr3Wte2Dy0T9abL65ss+3qZ7GNXr6v+zcLOgkvH01Rnq2SuuqJl2biII
380sx8bTbb3nYTPsjj+kXPhU0HCTotzXMi23qF3Js4LDKXZuz8JAdjR9bLZUdBa/RcwmbeUV2BMx
7i/+PxAvZf0tFzT9mY6fFO1sigHhKvUx+/2/daMGyhWWL2UY7LGrXk6vJQLECfTF6l047V0xTe9c
6Oi4v9rQPOyJaqpSVYSTrINr0GOgYYJqkWB9+jWeM9AJywh8/3t9G4luGqflakDu5Z0sSTMPFxby
+OwkmU7sHZrSxr4MoPrRJNce3c247yj4L4/si6Jtp1jk+IKsomO1jEuCjESNtrccYbpZa3rBb+NY
LricFBsgykTE9Ylc2VYnbRjmltrAlyq4gwD5OIrvEFQmuDyLPYviwdE4DnaKjYbZLK8YDXgh3WPZ
PVSl0pw7Ce4dDHuRZ7aT0he3eeZgdBFDTnTJ0pO1E9yrMxh8hsf3EISaPMu8g9QWsRGJvsgZ1CU/
wJQGHW/b32+gi5/dJsdoGcn6TGuHuHtFnkcQ84Fq0S78nqo48NpWxurvv0zwUGx1LQBIuPf/Q7TH
e7TqwVKdu2wb7/fJKbeBqlBaRRA9tSn9tAjC6IULK8XnazKIDJMmP29jAwPXppTo7i3ujBOhyi/Y
r7v87gvGTnBgh/oh2UHjNgc5TJNa3Xx1KUvfK/VWCszwIQjcJsoeJiXs6nzJZMORAIimugPg947G
U6t1X7cR4/8M7BAlYVN7XCQlri+RcXdn74usogsvjPfb9DeUGPFxDva8ghzR2yngtl+ImJX46Rzc
8TY9G7g7IfWp8IGugsqOIzwa6duUt0LpLvEJ3QQPj0Nh4iMH/EG6uoD/sLFMy55ft3wnGOJYbYdw
AYyv5qg4W/a9hfALyjmsHVINam3OABr+uiz6apq6bGbLXo7/j/9Jw0/md8f0VDDXasywaiiXJ65U
A6D3voouyGtjorgJfitEnjRlSKYwCKaziIi6JVjk9xsFyE2Y07S9I5p6S0U00TO5cO6JSqaJvMic
fHERh2JTUhhBjGDIP4CZgUsGMtPd/pO24Jl++z9h/b4p2DPGvJARdhYNPoeS6kowoi/yf4haBKpW
fpdK1srweaq4+ZpmgSAHuuyDWZORq4VebGpQPceDCIDLEzPnSdfonQUvf9022BxMZSbl2O+oSSXf
2F/F6FYNZO+Q06qRj4i6nVsQ+E9tqQEvYItr5k0l1yqxEF5v5dn5rHbNiNeg42hJogSyypf9votQ
h1CSnwf21IQTFTFI62DVw4gs47QOLOIzHuRktbRRYkLFCwOAlkbqYNdL5m7S0RdinQQ3hvqxg5NL
elcL+puXc+eL35p1/6y6jk/bgbyfvmEKcLAeWbZqmbmhfBPDpdoFpUR8JyF95GXt/JLDUJtGp5MU
nKSwPvBuPZQfXklWnBTWIG0DvmLuR1saBfvSqDhDJlM7yXRacEh6UrIcYjFmIWhxyLA0mfZ6xHEB
f8uv3AN+Hj+ty4qpe1BXXwnditzW8+7s8cBSFmB6dS5ShE8YeZuexuKt3SF2qTwGx4h1N+tgSNrt
SX25xaCA6HwwfV3ymSO9OQuVMNQQErK0W7h3E1XLj5hmkkZdXVv8j/PdRsM7F9ew59KLTdqZFTcB
9EwJQfKuxFWrSUelHhjzaojD3IzxFMNZ9vHwohgNFL9AX/G/VMDDGVZvJcXalpgD8G89v1mEVAZR
usLxmGJuv3egpOh7I9A6P4cMIwEqe6Ys5isIBG61Hlhu5S+FEZIV657IIwe+EiupFAOF8t/Md5oq
myE9Xwf4O/OUhEsSC5ZdtEzzESHrWQlzvQn+hhDrjMFiAL9uQUpMzE/DaJcDt5vokV1mKFjZQqnT
I13g9Mb4TVdP6NPGhjlAEobh2CaRlnEEa/z1DEQTgTnN4T0KL4OVBM3N8cMMXAs8M4QcnwjymurN
IaPDXvbpqgZUbPIdtsFR/DMSj8oE5kaV5L1Ew0Y2xoPL724DfSzur7eIU0V04+KQzBLp6JUg1msD
XQRgOSlBvuQkJAtvJF/oRw0ZQhA6z8hPKfhsPAeHDvDWXpJw8nurlDIRSBSIugFunpATuyukIKG1
dPWXrrSYSg3mpVHr16/0ytIPrOVmmxsyqqoQk6utjY2Y6uqMQhe5kCnuJvg8DEFbRSi6L2VM99Be
r/UP5wmuizm7wHpfd6iQZp/PeaPkBOwtCU4DxMSvOAlznmo9gNh0cwa7g8gIJ+BR5HZr8Z/ZI1mN
4rc2iJiQpoAqz5SBVoJQ+e4PvK0EY7f0YN1zDJUi+aYn8Ja6wTqCHPiGiTHy+gS6j1YT0apnnuDw
C9qVebdXeZ8MkYTGxOyGV8igjSS60BX8km/bKGzrPzZZ2JBFOVvHHfbnODOpprYSi05LveFP8+kd
Wp8fZrGi8W7ogvCfCZNE607Yj7KWJUx7YV2xSAW4QFKlaSu5y8sfpcWqNs86RzBc2Oim17cE66Nl
HReAWMBq25woRFsWyGBupI5YXVeyzjM4y+5Fub/qQIPpRWmYG4iaLN8jbTCqBRpI6ygWrnPMo8Aq
BUog6Y4Ccvzem8HThwghSVDoxSwrbG4pjrUmBSusSSEwGJZQizIkkK8eFIRri7YgueyvUqMW43/p
0j5828tGYHn3kHQ8TovOPzyV2AP1MEeCn7LjZEv1EmRkef4EAQsJfWFy3pAbWHza4qt9icETR7dG
olgL5GOlSJTbTOQu/aHKlCXgno6Mw3s1kYmhYxxNmaHxsYIWtGni0jN8ococISRBYgyEKz3/7lbE
GjPX3pPbLDF2Gki+w99Y+UqR9FshLiDvoNVUYaIJyPFh2rqJkKtHXqdsCUzk5Nl7FBkf5H8J+5iF
MtLquQLt7bFc7ra6HmWsatn0pZH6fQnc8l2N850jXjBfq93qrHqxBzr0uPi6ZqzwL0xsoP1RO6Ia
/sZb2mM+6l0SdEA0iFbQ0o8pvcci2hmI5Dg2fkBPEe2D/ObbfVyNDNBEubziPzJ2joxh5QaraR76
rBT516A1lSjseRXScXny73yGWavs1uO6iYGlYEHppfkIeowAN/UcTnIYJPa7y5MBT34A3y6sd1P8
r5TPdV6km78yTR035ON78IYQsq9r8CDCS/dfvBypilv6m2erSgqv3BbkcBDohFT9O2EnGdVCvtxD
yKgDq6Kxffrz+pcz3Zt3OSbxZXmmTGMMhK8RK5FltbNVB93zBe9mhVJcUm+FssI40JWyMZty2LPl
BPcDMhpTUqaNnA4JSTnkiM43aiDYoneTWS9xlzmSWH/y8ufHbB3BV3oHIurdfYyY/LhyfD8Hb/xf
PMZIi3trAsiI84RjhEoTUQ6bJFvbga1Dq2r4xM+76MaZ7KniSlljyWUtARSt+YtwWmDYPsTrgn4r
41i79WtaPdR/Jr753hkDx2jPkOiElMuis13gAiMutZiP9J+rWxj9yuh4gAS8e1+c3FdfwpJ8eyeA
bBxoFUR4c96uPD+wj6rEKugs9kNa+3hKAE/HdpH73dzqu/cXfLr90d+LpewfTMMmkZIqfJGr0JbH
cepnzgF4PPBkvxze5fkE1kTn3KuvkQCnC6uBbfF1gWG8I+J0wfN34Ads5HTrPwVmMelDWSfnFo57
CLFLWi1Zych5w93yt9563AmvnYvR/ML1JR8w86MEfYfwZkzZpjkvrW+dTFMmWB8KLv1ePAqR9FbH
2FaBSEi6q58DjqwwyRrCOAS9Q0YldIFmUoFacmr4zFSVnVJ/pzZqC1/+UbObuKqtIPImaQncUkhN
T/sBIUZXchuoHtDmjpaSzBbUSxqe1tRz2gY3QMNq1HE7AxElZEIyu/KnZJh1D5fmLAG+m6kcFJxW
VSdkexH2hFWYXT8jsVuzfZsyCnwYKr0Q3TyROP//s93BburcdNpsKS8NBn+RpB6wv0T4ySdaWaTZ
ztl44p4fnkr2R0K+HYXv5feeELNqTwtfJ1to51S3T5bQG9U5xlvL4WSwfU/gII8KDQ79M7/9uK/0
QHTYpJZAS5FUxPxzXVOypue+n7L0rhfAXOSlmk80IHVWx5nTMB6PsUzm0gWjyUcfFOworcruMrI6
HMoh4ZsbhodPwTXJoY4ENhyOCIDcYZ0PNhmoJKdoT7Y4KvwWngV8D3BdS2gyGDscO6JYyMLE9vVO
VDmK157k692eF/RdPUgR1tVc/J55HtVD6ZrUEgGQrwVKhgqL8AtZ5dH2+1djBLZs8eW9HgG2Z/pq
ZkUGuonwQJJEEtQyxwPaAnl3IyBQRY9h9lhm6e9y+hFiOIwICjUv9GQImW3IKUSql7SeMjKznU5d
EA4SkfiSHys19ymAHWETf5rT3/qaZilF+R4YB7eISawR5TODTo/esHGVUNgT2Gud+NFG8TQUfmLC
yTw4/3is3wM9MFgPXI1nRh4su4Pw8M/VLYrg8bK4nUd2Ca4R6fGlQfZ/+nC4B9O9f6YXwJUcU1iY
fq2PdKFnsDK1QgWQA2EIe5hMfer3UrZDh+QVTNVtLsqda7ZKx+Gmb4bJVSI1n/8yLTKXffmF6cxP
mnBR77pohM2hcm3djC9P9rSy0kURgeqF1RRfFH/OVv3FGq7zx1eQZBb01oGVRblHffiqupq/FTAX
RUX8Szk7zuYsAeGWDy8Cj1EltBPGbjSx5ueZ4rdgUnTVUNmR1jq/0M7lHpHfgWcSSNyNBIp9HkNX
2teH2ROsIfNCbNbwVJ4CT4ZocdEErHzisp4mKsGRgD6nAOm+V/cy+hMOrglhdJ6O9zMV9upja9P9
ENNIfnsqLQVxga/t/rzOqoN7Bn8jIRMrmDLqVlK668Och6Zu3fF5+TOUpK8bebNxLtwDXghQrvbU
yLHOa8wum7+l9uZs5KsA7xGpKcXV+sXi/7jIxOefowl28iG2+8mZrhs+IEH6P5oW7EwgS0fgPbJ+
qldEX9+m9D2pWIkIJqJ7DR1FN3AjUSeFY+b+dj0WZbnBMVZJPlRhpVFPISOQ/PYE0fU6n8jlaPvj
8/rAMLlxGzQELt006D017N63f2u8n9ogBuZNrKhnbCnvJjJj7gY+t6adAbY0JT1b3NrZa5ejKmAk
w95SeSQ2X5NigGCE62pIJqtDM6/7Jvlgx+sf8rhF2lksjRHvWt41RI9WfREav8vT3FCG7UCPpjZn
wHn6LvI8hHSDXpaGQBry6t5falfvNyutmBECYg0rFKO5bKIxHP6p6Yf9oS6EBCZDATwoG2cfd2cX
63l6BsS57jvZndPD+DgZQxSUKYk4yQVIcCoeGNcZKwx5yFMzPb4nYAv0jQyd89NLTv+3i6rDckYo
iLbK84vC5W5SaS1n+cYdqJgAX0uK2jWdmzwJ/VAOrDvosPREkkK5MhJJJHg/HLAGruGrQXU3wGju
GkM+PyxXIj1PfxQAOrPiH5T4Y4LeJ8nXm28ZRPkjlQiJG4xmWnOmut4yGnYz0BJww3tUiWCUQGuH
ELmuIThXBHQItWXTP+1cfwDGUWiaRJheTWeuTyTLJWruKpprCXJDf7g18Aj0Eczellzi8PjGuBuK
l+kSKp8Rygkm0I/XoYCMuq3hxG/lO4KISdeqNdduua/WjRGKPhiOKq/eNH4ZpA9+KAcVkaVxGaqv
GWxuTLuq59kliLCKm/MwtgpKpeZXbJ6zfSckiQ2CVpa4Ys1+9f8kGoZWcKgyzuoW+sKw8H8B0n4T
u0vD/qjFv8Luv0heUBvOsm6hrszwGzS9otq5or9b/0RH7hWozzhI+QpzxyIc/j3kFPxP46ewr9Pf
rlz//ggn/+WqFUjJF9ApFPeUipd/T6oyKKwBhDG4T8O1Z++yPaWOODAsKltY79Lc2YCcjNNDlrlG
wMYQXUMPhdPbdDNbj/zkHg40rU1A9P4pdK5VBJ9DAyyVGYqD2KIxvvq+xTr9SKvnEL63RaQeSAuZ
oLOITT0f0+BhoLjcmG1x87jkr97ZHyarhyr1EBSJ+OUFAmJ1Pl463t/pB+TS9/IA/089gwV0gVVy
AU64Z42LqDZZexf3HPvBP//uZDwfoxpTWwA+E0AHgVTjj3zdVCSPRkrfHtgb0GHbpNIZv0dgFyiZ
mjJBq5kHZZv6Y5gY9FDNFTzxalgaTSIK+16kPgCDMkQmUSj/2NU4QO1LVhRhPRH4+YAqQGCs3lqQ
v4YGcWKzVwnlxfAp6PgAGJvWD9ZkIgIQO2csJZmKR416J+RtfkwfhNF3bv/iwRLX/ye4x2gxqKvD
suyax1Qnd9UXI+GDqu6dwP5WbAieOLLqHMEfqEgdBjqCu8sL+Ku8nfhGTDQMWdIn+G4uUXBOh50E
ZS3gNP/1WGdRuIrZbWvTaPa7j0QtpKrXMDOJ4NtoiTaP2OadzLYRaMp/tJF9Kc1apGQ+5LqswISf
3NKsL7+9sVrWQ+6P/xiOlMcbNqFS9xaU2xx9UslGsjbCnzhXYepZ9W8stMeilEF4jqtg1qJLKqU2
k3w04+dWIWcnpNIA3OgnpMuhifYDEUtyiaMAIfPTNGRO5UqeQSGyNkqW41rS8dBKfFlLzart/Fmp
6mjPLDtDzcUvHECB47/Vnh27Xx+GD5e+uyVIdif2Xqd1UJiiDDdfzhk0S2MTpKaXvfV/wOm23qkT
fKLHTR0alUKCKlYTDDEMINXIc8v/NiMikbGgce1m+JKm/buvWKt65g7ltQlOjLpEyrqfr2zkoPAo
qVkoAlKSpAN0dU19Cr3kn9zwtphhKJ/2161hvdhC87PrlenpkH3PMRGRYa7TNfJPpIllNvr49+YQ
1SRU8xd7DizlfiPS/RRa1iAMleqBnb0P9BEXuhle96NoVv3ezz0ySbpKlyqbYupYlPtHURneJKg3
h+NrubLILWOhRG+ZPl1n9Rs8h8c6ImQTTj2nITD7PkYYVNEcdk5DMFpMioUsA+P3owuIcXbxIrm8
clak8tAh559KOcrEiVjyb95KyjRPJdwgBpLx8CFdnaolMv58nwYZd+YAWfljylwnBYZ0yaCaQjKL
HEqreyhg2CtPoi+QOLqH/oCyKR49uxyBrdE4fhhYBMJJbX4hXssqcksOEImEo22VEZK/xSHbnpqi
xEyLD+Ld3S8NvXreMhbIaRstM4GhI8nhdyZrBb3A5JvOrE5ytdMKWmcSuCx3tVjF/+5nqQST7K5t
btc8uDHHbH1TauHzfd1qFUUNXvBDIHeWKSUkyQOfm9gypZSdTT3Cklw1MN1PyWHw/GJcAu2qOTeJ
in1LuFJi7B3ELElwkGkT+sbubKx0zfx24wVqGkUA1Ot2zkS+VLsPpqg4tNT7spZcApBl2ofHwRK8
nDYQtPvHtHyhBkhJyv0NW6jWTLc6yzm9iNAj/bLJ0pUcWlrtBfJvwM8wnVetxRCoqkSoKEV33Ta4
IV4+S8grT3fCfoZx8J3CdGoFThesNn0VQO+xuM/yQcOCyOPxkecVqxdSZavERyoq/sGm6yRJqaZt
Iu3l76TQzSdLBwgiWcsGpYjBvSdLBDHFrXYXlVMWOtXZuwZ76SAAP/wyRWL35IiRVzYTGk1B9RQh
V0lg1ft1CdCUMEXJGKWNPr1fbByk9pO9hH3MwJClTRJkTp2bx8OyhG6/iG/4ULcm5gBVKYtXmCOK
/P0Hb+Oh1foBUbx9TVg/mOhdlQi3M2VdUnAqXByPtFYiBYyhxEPpi06k6g7D7dy5nwOySn/id4nF
xAazYZbNJ62PBxgW0n1alFxtIPHcTqQUut4eUAgLz53xDoMtePh5t1SCB5mRdiXvYFK4fTVto5n6
08uT5do5Oqo9CJP8gdheXRlDUcXi96YxhRParwe3SKR/rrITZX70TD4peG6wGfmiVrmjmqfTUd38
DO12gYP8ik4TjFR50gDsPBWPxuvFfKVNKhFbYRqUXm8OYSaFQweGRIOqfHh6kvTBxh53NWxEwPyY
+hJFGYs9pqSG1tA+5uMNyaFNB8nHmOKphsz6HfnSBq3bUM8RalVZFXniMsVp/q+72JrKidL+Ud4L
QQm2iDJFAAhvB/jM20Ty7N43rXji86zRX8khqWPKLHUjuPHzPE/exnldJBVUq4Nwyp5Z+gXkHcLI
HJMmNNtxqmDvM4hbsT+OnAEP66IZqHALLmeyRdtq4iLG6JRA9vSrzBxAaXgilw0BzCqLKTsLjpfr
sURx5juS+THTiOqGzaC4fIJ2joxrxz2Y5eVfkK7Nj4lG60PZlgoNooEJqZ3JhfpLoTH8vOQ4W2aQ
Tekdm1nk06NcZ2ITfN7Bp2wJxN5ukhwZf7KVLP0btH0euovMZA6afjjlSup33InZSqV+w2jQGnuT
fY1SBiSeQx7c9KvJP6vGwMQxG4vNUbry3qHZOD1h3yEWx7slkUkfkuRMU0rcYDgYV7I7CouNdUFb
NQI+pPb8jeF7SxU+iRq8nJK6lvpfTT+oOGgHdhkfYWN4JTP6RbVK3CU0Z6MhULrdv+49TLa6d1D8
1TdILl4aEa2BkiYjTVNkhHwdh19Lch8d9hUT2TQyNuFn8VzzCowJYfvqgVu7uBzVsscX/pngr4HA
g/z1laKx3MBBO4isLnMH+Hc7x9G+VUDsQzfpsa9s2JxxSqE6qRNNRHNStSg9YvzAqDIhqJMeIQ38
aE7l5nhEpCwE/6tIt8jascsx7VcSqBYilrQszGUrYCAUiytzxR0lxoVRRg623jc/PGGMp5VXHwni
HFeVKtgNaaRsbgeKZc1JfwqD2dQZW+sih8Miv17NaOWoLjik5FM+3dFrvTHj2aHTjd2EIr1Ml5bi
7Iv5vF+q3Edr4ub9AS8x4NPZf4a0dBh6Da4gPhkKdsCNkZn7UL9MEQ27BeZ+DYwEi+5Qxsnaujxm
CueEqNHccZP7LfplnsePOsWgRutj151lJ34+9OLguzJEZSwLWu+EK6Y83tM5zhdzFwGi2Fi4fJrN
Gh5tSh8+YhUpU34PctWtAtQQiciXuTzknNU86t+Ge84opl+XsYa8x4H+4LlHW5Tb+b06tyWTn2LC
qf8XkUfNpHxFOLQlQH9Zbtn+KvYJEZ9h2TCmkbtBcuAR6LSU0tx4ySGa3PqQsBfjrD3226XwI/jM
5FDOflsn6ISkOSqvZCxaUsIF3FHu/vtUVBfLu7ahNjmkGhiFPzBU12VooaCS2zhn1BEvV+vxH1IT
0w78y6U2m44HKhXcfuIvHgQ21cOulp5f5tie6vgms/rQ/hd1uNB1FTga9sVm/vSrvmJop3+x4fao
EqL4j0xUn6NhSXFU158Cr32UR7umaPIP8b1KM7l2J/n5U/eELYcJEvwPLdrfaF1zaqRlzVvpd+wi
Wrn8PzojvA6w2UOsNZelk4xZ/JkBtISeDAYNV6Xd5kwACKuuWH853TbwhH1cvvRROLwvXHGUcXcZ
pO4bFEQRc/E6mWDTa50pxlxLRbBqhUA6S/vh7x9GCfPUIyBgm5vCRHdxncPHaQgxwCn9vV37kI4g
FzNlKP8hUm7m9Ps8ly+qMvafBVTcwyfz3TeZjNNgwhxsEB/8Kthlg7Ri+ZjcnL8JvkUI6gwoEG7A
UVkQFnwqLH0YFgeYjpQ795KnB6XfU3Pxy9ydcFPBxq8hGHNka9ATisiHG24hsF1QBwoK0CDsPFtW
QwazNwr2QW4mTaCwiLPbne9q3EX66nn/UoWCtJX+DRKaNwAIivVDPEE6bd7jIoPIiGFTHe+m4JCm
C8y36FOuDeLXD22A56h0tZP7WUvQmthAstdG/aU/q+k4AQoLYOcZIn41xm+/YvwEwHpBFIuSZLoL
oVmnjcmJsbS/5PiliH2WwZZinhfF1owLHmBtIr831Jiy/eZ9F8u0Obd7yfvPEYOwxza52E2/1ZEs
yYiL8r3SC8fzPufNvdMfapw+SrbjqnA7NZIodqhWfYSoOwnbXc2yxSeYreJ2dWoOgm0pxAhJoGq6
0PjYgKf9Q3YI9I+i79CwHwnJkm22nyKGaYeqk85bzYaS+zYLVksuhKe2XF6w9OZ6Ez2NwP7wBvC/
jaTEcPHnT33jyfvUd0FLdV0H6oFlSsz7D8/C8IdN0o+nsokZq8D32rsQKl3VEaiYQ9ldr5C8WgGP
ulu+nRo7FYAk4OP4mhqjVufonfNg5tQJLa+FH/+wf7bzCFHLbEuof2WjymnloUaGoGVdrNVH+ayP
aOLOZdidNZa+6Zo9nLMn6t5WnzWhxNZaRYneoWXA6pxdTR/MpUl55NmAK0VXi92mCo8bnxD74sSy
5jT8Lqy+il4GGR3AKsi2kxwDM+NnmAkI+433BVIRMz9LURW0xVWFn9Qsyr+uOxVGwf3g0NwN32XX
TJrFdOsetbE7PdFdrjUHTl0fZ0BW08DejVPK0Oj7Z+H2L1wf3WmSGI0KDC7uJ7sBc6tuSw3PoQFI
pDDKBzJKARANPrAW1+GGMQrSQ8UP4YxfxAc7Sbg+UYJuTEpdrcwfCYX4SJ+1sKxwWbr82yuzuDUV
b4+O21MyZKfrp9tYedkQpCH5H+X4tgV2F53Vdvl5+TkYKKBmymlgy6sI1ptFC/Y6ali3D1LBt65w
dlMPiTL1lXeYJyy/UvmTc5e3fO9uQr0tPBLiWucltTfGkZuQInvDpL8iVA8YdhnyX+MRtVqrkqQf
nI6rSytBkKX4zpBLU5h6m1TxG5qk0BuuBf21Qb0kPpEYYq9tQP7EVm3xhkEFR/v5mxo0eGcU5xCi
Hu2odQ68fNVeCNBZJjePAIlqJVMf4iZe4ooQhF+jZbE3kl9ES0PTqDBtE44m+aUNFmerPzWF2uz+
fGomQRE037kba8mbz2Ilak5pIjNmYpL5/80ad/KYKdW/OeH7/ZXg7/JnUWkSEgajZQajZhSx1Ekz
UPa0odmlqm/QxzoGpU2b5ZL1aoTGamUvDHn8igGYrC2AweIa4o2b+F+DhtXWMUzf6XyvjB48ei7T
+ENDwXR0T6z8R2ysKLCDv4ezg0H9E04+DO7AIs7n0FpvRoO54cw9ff72kVfh/AviwNGP/sj655SZ
XZBZOPVdy9UJOa6tRCQ/WrN/GxjWYhgbUOD4l5ac/xCCuqC2nLkorbPkM5vdVxmoVdCg1iwT+jMK
zmgexz7kYhI8kpdUorN0GWeRRh8iQNTtCw8Qtvah5ehMXBidL2TxP9EeDfemBZp34b+SLy7WTkXk
dkmxMdaCIjoWALHsSMHaiK/FiXdUkqiO+05VTNRcuAH4K1JadO8h5Lb7rf6DDwtdw9jkPqe3RGnW
/soVT1byr3ozBPCBTay0zsRtcs1gTEtMZGTNAubE6YprxZZ/r5qaNhJiuUWG8Kpkm1BQu5gG45dh
KCTgX3M3PocU0u871TODJ6cfKj05VWhZgkf2paaHiXitd877Ryp2kc+gHRuPcY+o7t0ZWVJcXLfU
NoZOCOntHPk82BCWsvcQJwtxz53SCanNjKTtT81uhGAhKzGjcymv74XkJGem1UqErZU/SGM3HZ+Y
bOF8ImJb9XfKkXTVz5Sp+340ROFBOf9acLIUieUVjgyloRic8ebNZBFpZnukhkGVskv9HDcRJJin
zw13vOkU7BMC9rRBFOZoulGsMocG4uleruac1pets5wPgF7TqxW2tXXAnIAylpfWtKC7+Iv31o9m
41hvC7zgsc0qtHGGNPgo9l7QajWPHZVMK9LeoUW/0LJqPthgMze+fYB3Aa54g/WM1f6J9dYRUqEw
GQsgLliKjVCklFeUMN034xLnBe4iNJQ85LrpuqUD1rzaySoQaIxatBYOwCt5EoiQnYShtUsqIP+d
ZyXB1mkMga4+GkNteuqc+11ZRq0rgrBhsFFNnulPEj9kKB9wKeg1XLoddBzWCPOZDUwFMXniYMSM
QeDpRBuPHu29B5bLi/zTE0dJ/jHqF7Ph8Y4QwXUH8fSZdq98H+djQl8rjB5ig0PbGBmjFBJ1Logg
0GCq5Rw9U4iY7InPMTylO+GW6IADj2qUvqVX1TJ3J1ntwQI0OmbjEIh1L49u83XjauExXhyNTnb6
oKYSUBsdCkGaZ8Cxt75MD1YaGFHrkI0A3UV9Rld5qHWQl6WMNwzqY7W+N3+JMwDZU0WRtFfZmcCB
YnQjfO3BvMKizn9tZhvu2d+5EZrBdI9lGorje2tUcOG08Rq08hJYJpv8VQGpAwfaTLCvfiGOIE8R
CtxzvS6UIFhMj1Xzg/kY7uV+uDaGi8PJZECB4iStiyc6luUBPJ1eCTuHKOwqMDxNi/VLYILwOk8B
WqRqUAAtewx3QLK3v2tO4mmDkBxg/1PrAokwPSveWPkFMpr0xT+Ed6R+2ONYZvoZ49tv+LI5E64K
9Mfop/hTI9c/XMmvNUQ6fUen2f01uB2L926N4djl1Fzer8kXlimKkd+FcdlajzuA1FZ/xdMOQUGB
i0SEXoWbRhU4qF+9+Q3NhYlHeYw0qeQFSIzXn1Z7Q5U9IQCqy1FFgStIahAOQhY45AoAwd8wUzrr
PE3jpSLdmPkP0/0Q0BrEoHvd1hIoskhOCPFPmrtj8BdDOGQCnKUwQ000PGnoXnMEywU4I7nvIHZl
3AK4V4bx+fjM3bej69ZanBj2sB/ctUYZKrFauduYBMe0Zao5fw9fF9CmETXnIser9Xwb+e3Dxy7s
KvJnBswkXh5UNDaY0InyGxzXpmOO8yuN8TpPon4n68YypnJ0Ey+n8ujUm+GLgdgi/BE/Jn92M379
/p/U/BUBVz3jsF1ltPtz4JrErhl8ugOaRkclv2KMK2BIwSrHBXm0kKkAjjrn7aEv7Z1TA/Cx9P1S
0DiTioe0J5h4TLLgYh5/WxfVEeVc97x8Tom61tu2px4RpFDld3EZW8dU9BuGkh0bo+tsaQBC6Osd
KB84ZeKIEFduXk7i8gVQmZM6yrCrmFaBO4kTOTAp7nwL6mmshu2BXEW57tSpujC3YzWoomKHlIqp
i9AGofb1n0dzsJoWsqZlawhq0WIUWhuVRshomlWgHGJ8i11TCLkW8z0Uygv9DVK2iyvUmXLRS6+x
qq7Pk5K9ttPb0X2Ntt7Ja7quPyHDMba4GIQ3SKACUKK6U8eQiaZwKVdwc8pLW1eVa4BMrE1ZddSp
d4HiM9zd28NvYout/FJI5CfjCmPDM5VZBLWgSEzxEnYTFOIHCYQfW5i4PALC2T5AaE4my0uCrq+c
+Xx9bTXGy6YpipL+xlQ4XfwvWBihllFowF0GbucbxCiPs4lmrWVl4vETmGzbWaqEGRc019Tfwt3b
aM5YlwxMctKgxfuUN7NXYkKw0QQKGWL/kwAjAGU+SjtTYPHEzYjB6L2WrNxqF4JlhwR7dvrCtYL9
DVgs7JJ3P7miMTmtGR1IN15SOmYrQxipB4Nf4ISRf0X0PrRKsDadmSzATzJqfrvMediaFs6cMaMt
s/UmRzWKLcYjNKD6R/W7xoK0T6Flu72aKvKjzHXDylRhJy3VfaCdxXCxdPZ/igGZIJfKhQwe3xE2
gdRsrSuDSNvQ+gExyD72hbFSwcGnDCHptHnN+DQ6p+oRU7DlEG6x5BLm7sP84XMog9KCabIGJzNw
5xRXtQz5E8ydcJa9LsCyEn7e49SLgAOj2S/S/CcnTZ4+YBDnaeedAm0LjwDZldRQJsc2n84eLodK
eCo0iQXDA1IsdHgL3qz8MNwzTWheOApnGhZzpj+XOPzRun3bvJa9tIHXI1WFFB98MuAOig/yWtzK
v960ounbE0Dbj8l7/noahgzhzvjp9v4V9lxXVfn7ui/SU8j+SNHDH/xbggpfOvsbHPLsKty1vcxd
YkJ1l43FjmZKEdKKyumiB9mF/jtA8yDCziId6wBAMoYcaZCx9j0wr3yX0aNDECouqXv/Br4eyb9p
bHAPmZYEabeYhjdPz6muopdDV5L5CpeJ6GACAeuSYas/4G6YIiXgHc020JeR6T38HAGC0JYgXjQQ
tin/6unpvZ6/uDcVdic2bws1963o4VJYlVueX0y4Fe2h73+tWDudtSMdTwnUVSanktvTn+d96QeW
5eWOvwt1xJlq1v2GtUgasFB+8EQ3vdpGsGZd7U4awcn5ET56AvobdiLMh6pGardfs186dInLoY3/
H2j/vC8bpN+jI9btQsLcOcPOfVHh6bCwWiE5wEPYzf1qVjdft1eTM+nfkw0JeRRFaU1t/mAfnzMm
7BRtIyYlcPdojgmEQ2U6MQ6iNfdOOu2WbtPnG0ax8zWoGeVI94LaQzFk5/bXxjF9ItNE++UcOJQ5
lJz7WmsNX7YN+liAEyBM4Y5928IceJwTGexoFosDcT+yFHWHDEKC6H4l8258USgofEshlXirvaEU
0IHai0bMEiAlfxTXk0da2JlXfXXG8g2sclymLxSpnxaKTYVU0qSM63b74TjIAxQg0x4ex8GFmH8D
+WeEXvVCTvW2MTlUWGBO0RrlNqcxCKgCCIteQcf1QdW7/s6r2UZQZ2ajNVP8N1hrNPduD1yPo/1A
cyK5xvkLBra4H5BsL4kPDTHMsBviEUP4yHa79VFJJ55oBloSNC7cne82Wz5s2qm/NYGZecxvM08e
tPgHJk2ujcCJZ20pVDnzLeXlGWjdXxXgqyeVQEjERuFGjdeg2sgebOkRB7dU+sFsJ4mPBXpkNDFl
uGk5e7QmJnF9ePwBpUv/HqPBchdbZpkV+cY9Z6JCxR4w6Q7mc16O8gLnWVPymsHs7/xsYbNfRoRZ
8ce8j1T+VolAAHMU0IxF6c0vSd631Q6SgMkKFOu24IqW6ovojLK8c/x3NdZApkzLlYYymwcpAAK/
5a3XGTp7iwIoh1OWaPOW2hfXpL/4z+ju5t1r0yl98m3Tz8M7ibKNdWIA2ilbaVRD6hfHhiZ3V8NQ
KjSksyPAkAo+NC9IKpQYWIcPYJ1V4PHbvqTxsUEqT0qooGHxMwHHVjMlgmu5VcQ3RZd7N3GLcP+k
OY0+P6zTCWKbkY8ieqsUo75SyAcg8QoOUKTPh9KSU5pzWXShVdaYk4bCujatneEvuCfXymUj6vbq
p04RW1hVXtlCjibVglYaZCPUAEW8HWhVhmux/UJH6SWo1qlMJn9u4XQ4ui3tv27owyGp5u69aH06
siFcZjtYZOoQbdjtx1Co8sKMyJasycFCkqlV2dNCkCuuF9Jx9AWZtnYPTPeuMNyz9fUn8/CikMv2
55aQSeclejAU5xW38PoQ4kKd1PHRRgcflv+Tq2UjLrQvAJ/bcHD+wNkV/4FafPcAbZ4groHiDR43
kN0PHT+Yf98VaaWE6OYyLgvU81UFY46rvSARmxK/c3xSs4tCgZTmad/XiDiockyjwFy8yDorUqtP
RcubsSz3KauQuoKMHcfs98DT3FNcdyW0rZHr4Ai8CP701hSrchsmiGLvYjOykAB4WzNpro3nXFUL
liv7Gr7eCl9elRlYZVXB++VEDndEnAfVwn5U6Hl1R1p4qpOV5Bskl2KI9wqoIwffa/uVGCE1/p8/
RcmErhBTg/t87w7ZnXaPoDJRDicTNCDCGgiSlY8oWBnu8qmeYZJ0q6rJGo4ZmzUWecmFbwDMhas0
I5V0zHx+SsJABTGwNa1FyJtYe6s9JH9fUhND5HKrnu5q8J2r1B8M7lxWbttmAnr94TA2NVVPnam9
2KD3bT8TgnDl+ORHFLwe5s1AhYZ14slcJaJ6abDJTfyS2Z5hxK5TGB6fy4E+vmhbPdpXytetQEx7
8mJgUUOVQMpA/S1jPe6FaAeHrSayO9VoVKhl2VYWeDh+ZLYowsNsLDAQQdQWougKOFyZWHsjrWVl
G91Rn4LPuSryKyeLFxnMvLHUFC61/vK1YIPLfnhw1q4lpGesG7MhAvvVhoXVg2CfGUdFjY6Vu4zT
Qtqd+RWDNt0AAjMz4JX0S8X2lkxwZEchBhGWMaYjRUDadSm/yQIfW8RPzu6ByUMuqvJO17g4zDHA
Pd+f6Ff0V/16gR/uJvGgRfqXbzaseIY/ZLRt8HuPWVPxN4sQHNyyKfp3ArSybR2y79ykWKOt76bQ
A8Fesmx/C4d6CbohKEq10QYzeny9ABn3IBH3oKh1NYeD6eOssLXQe+T9dI+v9aYg890TMv7mcCth
aqlefgPUXSMvz/0BBqZ9FqKi4Vb0gVtYG2X81jdbnrEC4Yx3jyfgLHXBNV1afuPVYDpeG26SYo+y
rnlP7QyNyaCzY2GhLxxx/06SuXra18+O4Pjjpnm4wfIktzdfKTVpOtye7vBeJSXwtpoIZeCCZsaO
rZg4llXfMnaK/ctrnAVvH+fCM6EQTnQnoxgAXPtGYonyWKYroowQpokv2a522/fJZF/5RqIleiqn
YDwB/6fibgKMPEEDZdN0y7fTneyMfGxNsNcoJxnkYmWrDG/B/kOlgZfCc9eUPQq76QxkZrb9oZfV
wo6mfNUv4WbCNSz2UivwyKHwVOLc/Yl6VAEGW8DV/xCS3Oz6SxHHERe0rmV5F4XPx9nglv+0lwcH
sPWBpNunLQWblKSvP9VQ6GSY1iiEH3yoQwjHRZ0N0grkvaaKdznuZuRc83RmjNUMis64Vb2JUKye
9VTINCEFZbldf9vheW+SkRVbXzTqV8dNMYyHdHQzOiwCOo3ZlVFjO972YCroMriyOwEBUvnoz1/D
0Q7mo4+KcUpsO8AVF33gDxaOiU9z6xpLnNOuEum9fxEQ8Gc56QlubZsEBCDwJYU5YYWxQRM4ncfJ
D1ubxqcXxuZnWdr9RepkzzamMD62kjXjflQXbNPfsNzLvAVMoC/qfsdjUPXgAD3kfgC3tOmAvDk6
o9zDHQEWPNNLI3iGecDdzbKJ1yJJiKVjiW58X7zREL+CTPbiCh6gIEJ3qhGKi5HCd1Owj3sTtJkN
IG3himApKqwLbr+LtCGdYX5tO6cj5EEZWwxZL023fSgZ5RAWzKrurCdOpvM9wzXBEcwPYwGU+Zbv
4AiL7fthl9FEC0ef3hROttYRQfDQ4Ss4/CMQg5luDbuK7cnmzAbQubwdYczO+k/ZsZBAP00NfyQo
04LA/wX+mvmF/HbIUttvAHnTspxELZWrP9u0vR6hlBN2sgAOKuNxV7WCFSoJHdzS+W665ayfML5Z
2ptuymr0b1W/JmFdUeVYhHrbsHEtvmPEBT+UOp7USzbxKa9R1X7JAzZfAyqYq4BeHKAYga3LC8y2
+UIOqo8g64OAJennKuk9AHeUCxlMNiEc3+TW0EGjSwMdcynmBamck8E4fWMsi2ic4hmYrPMn9Yle
PXk6dqENGEXU2Ym/YurA+Rtoo52go0xnTjlwDFDgEbxKautzWmx4OPX2SVIX3UjbrDTG6jyzLI4d
6eRCCoMUx875sQokZLBykZnj9i4s90rahz3mz3D9Ne4UlH7V4F1GhzKSseUHIBbQ0+s0bRY59szf
Q8zdyJOmshAXVWkLYqWY8WI=
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
