/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 880)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbPY2B6DYkvw6uoLggeRjkFvbSIdJ3AwKN5WarYxppHbXVKgIqP1Rldi/
ZotLuGok7l7vOlNJ56ANIOiR5KyJY/RLCADGNmuvlPuXurTUZ33KznbDCjh2hQud0rhLrCUaJvr9
c4phAkVsehV3uZs6N3JnBLGCpn5EVy9pGuOpFGMe+4wNe5P5JAdBcff98do3QsPKgmcXc7P1ZiAj
Jr6SdfBuzYaTBqASjjlO7XJXgAUVg75sDFHFzXyYZutA5OKSg11fO2ZRyvyM0ofeMEhx0XT2C9aM
tBYhEA3uVly5CDzU2eu+kiCMndMUsq4qcJaveaERFdivD43Ja21aiuWtGtVELAlS/2HgfrKjrVnJ
p+0daHV8cxIz0liP2NUm2xumaTg+WZgq26FDDGU891r5OIKp91eumt/vbVh/qMLEmRq+0Ssd7HQ6
cHQOsu/LK7++hTaWGgB+1xuIs79Z8c+dK2Gp3+EkrH5rDjwZTV90U+YcLfFvHHymQ6rhp/hjxt2E
o1BfQ5/+rkC+zyuTgPRNaQ2OBUBIlEDoU7SR2HBrRQEMLfadCB+RYCyxmItR2KU30YjlUY2Ky0LX
PLjVHu/LUvHjxfRMhpU27U0KB6ebHL8wgvVd8xmHOvvBu8c++2gkDKrpBfC4JmR+PLmsScDoFXQM
WBJT29g3A4jGGn1YRUtX3E3WqOkeQBylFIrlHhP05xsPQSEwQdN/oGTh45r+1mpOH84WAv92e5B0
2jcz5aued1P+4Se1Cg15+kKWSxT6wnmdaX+knL+pBpwt1hXVBhkXNY3wsROYb+T2Urx9VLpTKT8V
+tqQbQ9WZctrZ9CdWJPvge7vFWmJSD8V74OfXvX6lSZLyWi05E6fyOzcN1woF8ORY87cl5NjQsDU
c23bruGIJbD5F2Gx9RTggfdqxOYnY2zSAT7HQuRpGcyzr3RkStpJ0DK92X4jAoVS5sQ4Npg33pip
KYSmX78TRe14PqJSgOO/c5aYaMx0JFETM1ZB1TvHLwpY9oCDwpIO80ZQaQNsy/VAzIWmomEcVAAS
rJreAN1QBqb9rP3lDXupQPGxPPM6rRnLv8QCVPGwPle/eh+p9A5vPytZQiPdisRN/JHo9/tiJ3T+
UpAP7RPelUmOm5Q8kZcygMpkJoMMQabF/g==
`pragma protect end_protected

// 
