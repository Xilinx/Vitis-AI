`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQGDi5+1T0zt/Jw20/MosUf/BG/H
bU1FHIdsAm6uft+7I5naFNkYDFv6fsxdnfu/MX95XWwn1vRNirzvgSpKb5hcd4QOYknPGL4xojGp
sZ/5G0qZehfOcSBTUwqBYwtM4gmLkZgrLiUWeW/+FNXWDn0NY2ltMbohM50vnoaoynLxGMkjWGST
+ShwzZPpZgxAGOV07TAjXi7/AwOrnFMZ42eEcNsk4cV/EWOJETvBK4Qlx5qPY9o0o6lB5GCXTCjc
GpWToZVWeO51aACjC5QGr6bD6A7j76UQZGLZ6Y5ISGyuM5f6RRs1B8LcS5i54fbeyb0dwKE+3pmB
/gWHwZrOvjslPwTGuMGscadcs49x+voA3hy6lF/4R+DjhOE1c3NN7SAQiSLjFirrP9Mk7AD3+EYX
iQiKVfC7LpKJYFMFtK7brlqasy4XZl3px334sysBkdDvgZs9m3j5QiSkrVl4GhvIY9i7YanMOdVh
ddCfLoc7tZFKbQh4clZ1edxVV5QXiQTaWLrfxszA3WToXsFNRbtOi9dXfLjDvbp/Dtt+fYTRkpS0
yPGTjNXVae0Cab39cDq4N5rPS2zNd+VcpPlHHmbgJU23Wm3qFBSHU/eZrOCaZu2wZkZwm2r7tCCT
eEwfaL1J01zegU3J0nia/y9VzgkezPzL79fdmi7RqzzicO6fxMJv9XkSjlqCvfMGnnUK6kE9Hga2
gFuKr8xeM/g5p4iw3GaGqgZB4ilhxcw2l5hjjlp8B3f2hEKJPd5B/of2kkJQ8LvPpjdETJaUP9e3
OM0vYhN+lK83NYwW0DEXd3wWRrHimfXDigZOhq6PWQwgtA8Fr5fn7yYOLokaqJtBJkEVGnh08iL0
MyZq1Rh0XzdNbIB6tSj5fIwnTBTK0MiXuB91uUaVNehb90fUZp9KwFQ5gslChUG3rSyh4CLkzVjA
JRQ2NCLzkdYB5WVa63jwjd9lPLj5A9dLvUH3m3IpY0YlGrKoPowVoNUMLi5gSj7sVoKD/HS4WcMJ
/7abaCzu9ja456PlTcJNcoKAdcz7GmDpA9sEdoZMJiviTz0F2pmqRANBWGQ3bL8sTimOSOWssLBX
/h6gY52VSZnI8DuWQhjpmE73Un8IXptrTq6s8yRl+PAYQSftOHyE0frf/l8P2sqinE9HLCcDkv2q
FjrOonaBt5KwSzFh6U074PSwcB17QeJD1u+yky4lr0a0OavZ+MYez3mg4OOXlDNcqX/43b+kyVTc
SKQKqyxjT9tqS/OzbYDl7n8ISGJubE5ZlXBUR2Yur4WuNCbGUVbeTTBJgB5NhV6AOWpdieDMD7Vp
ooM3ie1fd0jx5EWE/nnPaSaqAitno1T08D1vrlJfqalcudfTpzGMejjxj5NKEK3aQYnHQrzPOOIz
ZoIO8K5Y9wkaNvXFiybDlyjwFL17SVdjQLBygo4yozzzGOgcTSKsLeAw6HT7dihYHBTowVFP/6lo
kNHq3qM/wcueJozayXc57dPsykFp/Lhg1DCuXHZwgwGIcebE3CKBofNRQbe2k2X7BkuHF6Gx3c2c
Id3M7RH1KOEgMZ7G6tR5LRqeC6Z9exUUw3mXlECkmgH/TLwKtYmGba+NTIsiFFslY3p9Lp1hpA8S
C+J1WBUmBbc5WNRgQXZ5c890hSLhROSTHf/042hRYM7T7BbDWGfnpi2Ok6ix0lZjdjEiZLYl7XBj
3BIZc+t8nS6AjSmZj4Tx3NTvLhJJKT4Vwn4CCbxAL+oQ3nXelCF3tiGgO/J1zVW6uvbyPNxlk7+w
vDeJs/bcbyt9PUq2Oeu4uGR9GsS1ynZNlGiF8N1GOHaUWDVE9WI40MEnXMdWdUqqa2nZk3BuJvRA
YXDwDtbO0W3tvLtu2ZzpzJ9bDQ1beoUCMs0mMkKnlI/G8TGni/HMclx/jX95sXVSTsZ5+IN1U8X3
Q/phvqohf4qVqO8fZzvomC5anXuEe/p/rRfTTRkjiwDTmUACJtbJPbq6PAGWYxHqx3F/ADyDGB6J
IJKkjgCi3KNL1+3+nB9f7CZpO1etJ2Drbco/0qNthaerrPzGd5R4WVenQQqMaNrcbGouXikd+3WB
clCcZIf7r8gD0DArc/liG894sQbaJVXFqQf62z2hmzR54R7gvrZ5USOOzFlvpwTm3Aa8haUznzkx
dXkNp/O7o/RRF3aEyGGQ+xNtDZfCCR3xpMKvKWfE/vumHswIqaw6Y9NVBFwSThKw0vDgrqmM83xc
bsxwkyO/lwDyItGwiNYpAk36fCaz8O1TD66oHzq/4x/kUiWeSaqJG94yffBG6X1A6B9l961atM5E
yiPTtxg29z44z4AEp+O/ZI7a5NpoeMWElcunf1Yp0h8kOvPZVOIDkoiX2lGOmzbEQd14rILcFU4Z
jIh4IVxGfbnld1GGcp9GesoXLa0W4zbaCn+daM+1EB3nXmNxtH/Qvu5muaDKWj66oAe5PF9Uz6dc
QmX0L+ZmFb8u6opEnproAzBTRL7Z1B93LdiS6/BC2HfyA5SxOEUyIYgT4VVLF7AzpC1t2CTVQea/
RVneAALCj1yhjBqVpLmnCxSfqW1unjihCcUoTEk0Bto/aqB8inyyT1UEkQxvapzQDyCjSTzN3lpZ
wvmS6k54MAXHSTxreaxjzlViumu4OHgSIAjJDx7JXqVaDcl0n1WVAn2AYSX2gyfHuIFDFH35zrFD
nXG/D/g0nxP80dtXD+p352Tqtazbq8sSEya0G1afcl8b7Wb9/AxinW+ifbAOx14SMIwAYR5Skuy2
p7FVHLvYMiDrgJdzJ9wMNS9gANn5U0slq6Gf8OTOHrpscU3BfFeUDxVY1Jiht7S4pV4m31fvaPg1
cMzrbABzYLXvVns5m5B2AhWUulQpixhsfBZtFnvjBL+ysCRhJlfnHFnSIu8CPhigQhm8FeaSs123
BscV+bd1qhS2N7ng70hMQ59ayt98+dLg1ongjxGbQpMHT0C5nMv305TIJKQ+4fI6NL1nv3JuY2Be
mSnW4ffWFyc6nyyCSpAcwqcamcYITfzSkLJDmFOU7SgeVB4WRQG+KSJDVoq4zvpKtp35m70of6ui
sceZvgDDuwAv6vgzIE8F7asE2pGBLaSyjXrJ20OXNaXMu3IJpu8QrpMJ8EvVY0J1dU6rPBsBvTfC
2sJOh2WR0M9Jh+PYZ79VrNlZIMZyyoGAlYzVEwGTEErhXSHs8liwsHpTOtbkhQJx/lJ8kj/Hurkq
h0zn+JYyEV7MxkYk6hkK+9Xb0YwGFVuFJdx5ffxBGZ3VABfESCuRxKQwdy/50wLNFZS1GhAe8UxU
uO47XtC2BAHgURqYknEoXmjod8AL49qZZqAZ48xgOiQgqTU8tY0q9pL4/r7mvhI9WsQR5Y7tpRFc
Vrt/Xp6hlpHg2Iga7FGw3lJVwRRm/SGWOM+HZnjVBxz9PKo6XJSPjjDjiW8zVfP1EniDCBfpA75u
mQkIiNmeEYhtE2Nqd4E7oPx5oVPdk/JYeXJQk862N1ky/Sq+k0O0e9fEyWx25LzNw/ANtvbT32VR
ZPte4Xu1fQXAcemvsTbtvqNazwT7xxR93Ye48R4oSCSOMiTXZtzBfUxmI/yAO3HOVK1uhC6abF1k
51MK0yR+KqQ0TQ7d48jYUqRRnnuKEZSrlgwzfXR+DEx+6KjHHKVcJArfZLJb4/PfrVbwAxKWHRYg
4CNxdwacUhTtrWM0mvh4Q0XWyAxHVyema7REk/T/bUukW2v6ZknhCPHNc/X8e25cFsCopXn6TXIR
PRku7lMF+Blc1VlpUHnNaBvXvxxMSzOLCZbKSvVv7Pzg2v3BKdRHAGHvBeDTZbWaC52Iyc1jwZYl
M/kjKaAo9StU/7nLlwDNPb/hJuBcGo6z3Tx+PZkwP765KdUmipzkymbEd7tAQf1yxGbBkUUnTabs
bdGmw5ho7nUyB+3iDZODuU1lOect0rWi6K0QIsUiYPW7QPjeJMNh/Kb6Y/en40H+PUm/YxLURjeD
vNmgr+xgToppW7+d8s2JDN9u75Vj/DwNn702WEPPLp5+k+7KVXLUCr7/1HaxR+iuUyCaPyc8eC8h
laraHP1fJI0B944PbdGFCb0yNdiZWsNHCM1sPjYj5w6GDz23x9X1SXZGZyqYEtiljGHcGCYklyUT
tDlpsN3G8Pdr7JRbo6Ce0kRqSgpowq/3B2pskq9o4Yv7xCKXsW2ek9q3+LA52tGgjBN8yet4Dzry
G5nX+npDUAbGvM1gwdwSPwokOZb5LTTEuhe5LS+1VNoBQFuIZcaPb1nlRzLracKVsKFrnKaNnwQW
qXOrbWrU92uFQOwARagXJvqbUxgPTO+mtr4J44ECSOM8fCkKYRpGEaqEHslJ5Giu08TDEPOFspkX
c5wlAnaaCsTgFnrSuGmvr8no6yzaHrMPhcvYGopKDIFMA3Jkkzs7EEhMYYUfFnoHttZt6GheEgNq
sKOn2oGn5P2BcgpyeBeJw7cRRcQnWP0IBE8FzT88WwY4jKhIKZSRBv7XnTFDjiWf3qciEDhRKLVQ
j2yYk039bm33HfHlJOIjdXlrbS6vjShdXHWwc27FFgZ+JiQK1U7WQxRvHs0veOhzXD/cBxS09dRq
cUHhbNz3WkPOfUorkxHhdVuPAh+i5O+goEVetLiciRcG5PF0QOPEU5eQFPbXZ+sMNUtIGiDUwcaS
lmNC+locMevqw2ierU8k3L07j7wELUdnvobcexro7GBp12A3RJL+PURm6YxFUzrK1WI/RNIxtrmN
xLhvPA7u0UIhNDWjOyw7lxsRhBt31W7e1m1p63irQN6i3MgrTbxabvEUkhWJTNKlnlyAFiPIveGs
0ZGejMeI5pr6UIhsztYNAk+EeJjZgoSxHAha1tJXa/IuAhpR5yxDn0DA+UiQ2RcuTWDG+GP3M9ke
fxgdrNX1mnqjW8yPkgoM3UJspEq0LnYzspYbwBSd8C6vtf4iCRDEYnWNjuJf4C02vN9OsXSQTZdj
R6OVv1ZKdq+2vzHvvEwHDan6Pdamv7QLXgUCxPahcvL9g3Y8chWlbnkYvz4VF/s4PhlnZN5XwAsb
2LLolG2WY2iaIkfsNoOBAO8auX2ktlmJ+tNIU6oLEauLnYCBxh3O/2jMirNbx/5tqQQkyn1gDkFY
5Y4sMpFSoPlqeZMFN0i5yUzBG2cDE/qLT8aN09mSBGJW4nCAMy0uMzqTtpHMIDWCASWFUKmwkMH9
vKPT7gRrE+MEW8OntbNK87dBxjOvkTB5PP40MK7hyTudea7/WfVQAtgpJEn7hQzbfNxBL1WPI+vH
KidZLrc98Mshzwak7Cd0d+6DK3AouBQPkPtvoacWw/9bpy5tC29wzifUxQxA97fnFcAGUMqhLFio
gTPpg1Pab7LtlKHWImijEaZTnx2PaiYZ8xjXQD2vuhpNZr+S+/vV5GzTy+DY9y7s7aBApOoJt92j
7CufehBPKXLkoZALJWEEhepqiGEIilu/fYvSpDufgVPXZ5tCGfldB8uz5Ipto5jfDhQGCmQMw5Rg
Kwbl2vNmJwt1bg6WlSRQd7S91737aRRa49PqxMUuwQ1o7C6TeJIvnxyRLhlrQ5PnXoWiWKlGunDW
mTZwY094hZoEchdyZqJ1w9iblhfKM9pNz7PcvAEeteREliPHH0hKEeE0JiuDCEVZDVnHskFDyJbg
qW3Olt4WOLc0fp6upybjOK7iPOsKJbSTOpAg8PN/oFfuiVWmBv4oInSmxdybPRXjRleSAw6sm4Xl
V5P0Hf038evpmzvel770M9BIijT6+FuSc4Aw5OUuPr2SPVwVruWBh2/alozF8YBtzDHolO5v2Jji
BTLxlKgwOtIZH41FAHaIaMTeEwewFVSE+gHEGlKak60woReRDXHA1DZguWNbvMgefBx240C3hoXg
mXlVbtDGCK74aTstlL4eHAFMLes7d6V49/7qlkzJR43QnGHLlAzTkhXz2fXkzcBAFz4b3L0+jgNU
FML2yAqnXy6dV1/Qk4hrWx3XAbcicLZHtRzOAju+EzKTq8w3aJsrQ1a2H28VRkuiziW4sTX1mhiV
4mb1JB5R2j1fNIxVjlF7IvbJODbNIGdAajrOdJd3bnNUof7DxrK/ox6N473MugOmkl/Us8VdPtHS
aGCsKrTdMzfO18zTc0M42b1cJYhNwz7DdaKvUlp5rA3fvGUs4XVgFA/jkFdcj/W4L4Xxjf/xQa0y
hZMMcDIi8v9ZZ1Le8uicOrEpMwfbIIlq2I7U3MTMBFayVNiEg1jplGgRlOG6KMrGbgBruItMT1l5
u3zqXlXxrfXuH4XQRSZKrqEdxEkcfLU4Q5NcvTxUxiGLoN9+CBsaE+FHnsg9LoEckmjarOHI7M4S
/DT04/0EvRG4RLu0lZZ69lhAO8YE6zkauKQH/4JUfVpANvtlljQ0TXhluZgCmJJ/1vJAThiTYURW
qWyapX9aFQ3Tx1mGOHHNlv5Fx/ojsjyNhI5BvqjQhgX+ryNKWRJ9OdiXLHEp0NwELEHCPPXGk4cG
JVxAfCdMFMxCK7XXieD5Xsm4kv2X0bmmwlT0HBGntXL6+mU7CnBAS33rmlP80UA8tuhS3E6qaBy8
/jymN9A5ni8zo6yR165UkOqHdozFSn3odfIzaW1meUWPXpzA1JBzb8gLSdZkCLYeSHCMTXpJh7mC
L1fTT8KhnCKXRIBR7f30m973DURo8IJfjp3Lpsu/aJSxCjtJM78gl9Vv5Kv3eZTXebkZHTD62iLw
4hvab1CjD+rWjGIOSxFTve+MLhP4ZUjAU5URAgQOEQNsZGHrKrMSiCddNKpDv6yO7gUDSytqPOM5
BeZyub4B6NNQBmkF03vL1ugDoVIywNyj9l3xLU3FWaHNBDDRLgr6jNk3bBWTOopY3NS0FFDgMo+E
zcBXC2hakBb9JFR2qa66xKCwgWIKhzCblxxVgaRPStgIwhVv31su4Vs1a7xtLEL53M4irSxKo1WS
qTwUaMvsL544U73uX/8tEd+GUu35s/rOk1DhTtAFL3786JknD7Di8jZjLLhHP7VHL+BHJ67kYn6d
QjZzxqoz+3Pr/Pqv5hpMULMHocLkMPoUewP5ZYqSGVBZA2WdsPPE02Fnx3SFnFYG05RW5+dmBc61
ApGZTxI3iSzu8zp3rdg6KAzIdAa8OyE1PhNXHPn2k5glmYYwB1mlP9Vfui1U5GPNhhdp8VKu6iu5
5htfDs73YvLgZZOD3l7+AA+ognoFKZx8ZCOgXeP/KF7if2OxScBcxm9ET6N6Xj8pD/EaaVX67NaG
clS0TCct4ObwNqY6O07YTfT3+9xgMT+PpZ7qlXPQuNPIKKISdChUcAF3mVtLYWLEvELxw1569VMs
+23gV+uOqZQd4fMpotFOnHThi9XEhL1wnNBeBhso2j7taZxU1ZMXOv9nU/9Yf9M3+ssKV/kiLfuf
tyTN8KByWTOWZU1sgOlyZi7emRiH56upxk5L6UvpQ4aP1NC5iqYevT3qV9vCaiuNmzCsIbnBXpps
xws9RnmX94+fw/ZbMAnUzWOFUf7RQs36Ux6whiclzEOhnyQKIxjwvbl9se8cb5Ld+4evrQHkIzNJ
5fqI5iwqIXEfdmOGLwMK3yuqRUIFWrNCav9X5BxhfDdB1+/rUyrtV5YyM/fwpdEX8DYDn5VnyCb/
Khrcq0qjQHuyAT3hw6mnSPieEv1AfGHZ6RH2TpFZh3bEGSZCnBPh7b7+ZZVEU9LRKNmxp2xJPRM1
YEEszvJ2uH57Fif+SbDDXxx47pK491kEVN4R/WoDrB0Bpvx45ZYONNoeEzPPmcae6hU67GmD/+TR
ikfht9KHeBpWQXL2do2P2xF4CDU440qPNAWuxdBxhfa8v/Z+jmB1mW5+oVbda9gc73LG1t0zM56Y
hagcixhB6lva33a/XxNDNeV+khLKLwJxPxE4cXKmpxwUF0UrPM19Sbp3ZCQjy1UU+dwMUrL2+X9W
ZSuCiZZBCy5N1SCPb449dQ59qVk2N+6EPbqQnaWhmwXaoboXphK5OpsoUQNK2wZqOBmRci7sQKzF
L9C2fMOGE/gGKnV0weGmhMy2CnDfAJ4vqhl3f7AfceWlLtRQ79GBHZC3YMKeekpAbcwN4A1ojIE6
WuHx7AU9QwDXr8R42TtK+HZ4Aoz1PrIhAPL4irB68fktTZMkRSOZuzjjFr7qva5JmE3Abo9vIKyD
2XikLsS2ZTQ1mxtUHFJuj5uyV/z4I5lmvvG6l8orl5mlpD2xz0GOGMmhTEvpz1yBfJQR0czPQTVY
o67QYp294UWugl7gf87slsz4yj5VNfgpoK1fZd+P1Yjbqxw39HInumTNZvHrApmgqhhuTT6kbnVJ
pQ/lzkAEqSGUGaDSofdlfMSwcjma/iBT6Xj2USLWfj5y0dbuchyqmWAIwmAUC0YC1m6FQGDHmlZZ
YwWqXkiQu1A+T9BB19Nh90mfxSl2WQZERxw0IF9meoGX3IIzUqiThGv5vgiiLjbx6fnigkLEl3Vp
ScoOpug2VXLuVw7fLJOkwTTxZU2TgJIvrL+FbclBBsCqQUQ7OgzBFgYdK5ARc7T5e0d4eF9BCzLs
l01I4XzTYC9ivBfOL4hWWCwiW1Ukx0S8THaMXY24DRXpZ4vlp1v5sy791teYK2fC7gjzDm9E6iKj
waK726qqn7sFnTVVwwXgJPMOC8CO+8E8hJ/23WBNmc3pDbZ/JntoSWvgaaXOVzJlDTRXgLoO9ZFe
OBAXNL3l3L5+gMCUisZnD1vBrzRCv3RmBE/nJa2Yqw4egEqjjmF0ofQmxs7MLlnBjqL76NItk/4T
bqPpPM5tI7M1MnILdx0MeZ36QKIOtBPPml5zDAUvRA6IUS6nK4x4tehUdcJWxmqEbVpYjShKssTY
LKgCLx0XDVMsIQnFx1/jFlwPJB9qLJGOnXP2kBoDGjFWmr/dcxPaVSe1165jOcI9Sr4UQzDJES2W
+TMciA19gfvartO3Mgdy6fTvdHHnHrkGWlpWAcaRVZWMKItF7Wc6k0kNyQqlnY67qouOiFsd8gT+
yGXW1uq8bgvbgcoYTntwxJjSrAb34tc0r7oLV1h+Y6BsdXq01G55oh3FAAWG9WtbRqscMwO0YINe
7agFO7aEJA3gMZ7jioiLQJWpQzWcbjNGQ/nEEYOKrET4vXKMcQqdAfqDuHfwgM4DAR0EaBZws2kW
vFY/GRzC4Um92mdVleJGBFnh8hbmmo6VQ84MFj1dJWbZw4gA5LSq84GULdsA3gcuOY8P/xqx3LPY
CA0uvoluNCcs46APcud8WBkPA7xykRvdJR8UQc3C8h/yiD8GV/wqAhpL6I9uVobPHzbfYk4o8yCp
9xFiJr/5IwLJZLAhZd1tIjJVhuP/dkSPk6vmBP1q3jyaA7xrpkiVZLKvT6xSAh4iHZLbBvT28L7B
U0zzq/ie+g+x5Z3y32ngZPbDIxwKM5mKdlRtSUdYW5cd9LUZXh2rfB+KKugtmmj2oWQhwH7NULDv
SPM8p7xyJ9iFx1u0u3RaSSJ6Wn7cZ6MmTGSrrjiiJ1aj4bng4iHOuKUDXWjr+c1v1H+VYEuba4He
kFzLy03tHZcLskCmi3AXIdHnjs7KlYK5PoKiHWo33LR5ixLJOJMunei+eE570Oq2Hd6TmiNZQO9G
VQ4iRy7TfUTknBtQPt2h0YnGdHCxEBvUjbbxfqoXJSDdszOBPm/jt4V8eH9xaM4Udk2GuKbNMkO1
1qxgn2G13MFtHeGEyVw5wQCwxZGeiTP1KGKGosgXMCiEHy8mOdi5XV0EMyAkWE1bZhs8wxypHaOI
ZCxfm5XrtRKxtFOyfTdeSkO/Jv1Qx4M/PvdXwhwxWZXF7EX1H2Lw4SX32vgmiU7LzXl0RSebOrmb
341484N0qflcXrKldC53Ku51Z2mQTXX7hIgQJSP1511H56uVwbeFUp+HXS6UB8AgJNKyfAy8dQaI
xIz9n+QPzEvZXfeJw+1glPBarzpHyDLeeoLtwsjRkjnBxUQXTHp4TrlFR8mqc3fU+ysDDknZ+/57
ZO97Oy1TWDYpJKhtonJVRvKfzExM30MLXjTwjPYTW+nYVTR5OZA0Od214io/ZpSSsCfPTno+EpRZ
hnjB2hT/IbcIlRz9MM8BIxvW5NG4Ell+L4EPS3KQs1y0mfWsPIMWIMCSaENfwWVp273f1LoKs9h/
i91oARKtK5WGxWlqqewVRaMbrEThPqw7JeTeEDjQ5AkJxWFh/4nsESud/RRaQX99puhlhdrCn082
VqcnxOIIMLfPhdMmh2N06scVG06denuYHF+yp6/Ox6xd68YLMxT4xOyBketha4ov1rwhOGvtd3/d
wVnH2E06VauIrTEEOhhna8FMTlzxWDruWDWSyfocJt6bp/KYww6rPbSncrjpsdoFZToexPYWIckn
YnxQt3u/jYVB6DYIW3qvhWR3nIpvRgJ6uiTDW06oLAebQMwRsoySHjyA9kp/gGXw5zJIScMkwZNr
2pmfRwqgkMnnAzhO1Ihpds6ewZG1axvwpn/LTdNoUaW5/9f6MOHj13gHh+yrzb4F/SsKF4LAOzMA
PHIqRj9z+iyoaClVKMGXxr19JKNKbLmXqh1D/4m/ojp3+WjIHaeEbiOuCIjEfHpstpIDATEDbJ1x
7Fh8u7loJ1vBfjztJvRnNoyZ4kyGWmYeZ/GHys+a7x/i7T2GOcObaUzxCB0Jnw85KNiGsuQVNUz7
/WoUpm2HJAppphiLkypsERYuGFD5l60N0wWucufepwlX9hywEV7lLjz5L5bjQyLzjigpfWXK+u6/
YGAk0tHaaRDtka54UUs21DYYo5+OXRpkLvSYCOfX+gvWRAD6opUyg0EtihhD+fmz2SqUjqzVk6k4
qJDO+6mBL7o0ekBi27+UJJvfCxnYfsDlVJTH+gc6FeLl2HYsbsfkiAgw/uW2l4ljqtbVuFKXkTsA
bm/W4L5SAr/OiVbIAHmkiZInGw17h6qeSnDpzQcstVjtLp8Ozggckp6j+uoENQpqKewyWr2CkEWi
+X/7khybaOctHuB6LoHhAJJbciGnRdpdw6qvJdk/a3lGez95qieOhDVmyexknC/GArxICq3WrLyJ
/8jIpKz+J2gelbPHhs3b2sWdWmgOQ35BX2K4xrU/H939fQaSsVyperVc9r/Jl+Xrr2A4ewGTfyAP
Xw7uIR7SkFCDeQ7TqKicNa00bDE4gUfHpBYbW59Q1z9JHWymFihcAl0B9ea6vubICU3Y0JsvvB/L
INkzP8lnF81qxFpWbuqjypNluYYZ0jSKz90JHzRvnJrzWDgDSYajS7sKyyZyFxvR6bsZFNxGSsXR
dnLpAXY7eEfTW3N1NBwbkvf5ANJV6kVfdjxlSMFRKrLKPxvaM39TIXJR1IKrrLjrVyfEjzhfzFCq
fHjrxOURvpGHg5aSf2wYdcl0QA54DVhbPywbtqEPz0VvGYsW6CMafP2lSmCIHZi5YTmphduo8EBm
iCDY4usncTG7hrR9vivEtvO6tpT7/2paWKWCcxpXE80unhgYaDdMygUUMfMafw5q6kEd2ly/+bv0
yvwyA9SFr3p1cHTvz4xOj1i/hG6Wq0W0Au0zCvqUpO6q8PVctseEMP9CMpypG/H3KdQG1djQFCVf
qzsVsUlxX8GnG+irk4gGsYab7JhPAICuEmekLQ5oQW8IPIIz7GIYmhJFPmGjliCDGKNsIi2nMdnN
3HCjOmtwTmc8v2PJNW5IN2PX6ix8Sw2Rd4yOjljEi08Qv8cfZEQD92EXusIGYdSbeBDa5fjNw0qY
Rgd3lSJnScn9o2GtKuQUxXyCnMTUnaEYucSXju8MgfFIKIv5ZVDOqzSgr3N8LYw9e2HRW2ljJCsx
WBLx6vuHsJuGB9cUHzjzISvvFkiFGMuBsJ4n4NgeHfNjnIQyOY80ZFnoPV4TSxcvwlE9egg+MyDb
8/OReViNY3IOP9QQR6VajZz9cqn3krOziEKbn+Cne+Xhm1oTbJ59Tk9XrX1O8mEZrPTOz/ku4mVv
M4yNa7ibYohEAY1Gdl0+DoPiJq+UwoNQtgp/Ip34eOTKmJ0xyLsM/1bAM0vKurJNzik+9r9qBb+R
tfTbyEu35+MNrv6iW045VYOovRz6bx1R7vSn5dYYKAlbkSJgRrpTAKGcO+qrD/HaXGI/rOHvXZDt
B+4NYb2uKMV45HChERKgVetAUYO/Bh7IK46BOQ8PuZpGplwAXSrtMhF2f8hxTIJ07FO4PX2DBMtk
A1v7BJWJ9Sxz+09Ks+P6Y4WZgXqL1h5ntdC1Omj38W1UIJJA3xPIAzzHqHCS1GVcSUjbvUOIMrtc
mssshYGJl3rVL+uWCCxj1XaqCr/LEGQni1NsN5flkKYvv1Ex+zoCbNtiaZX++XPP9yINFvXmGWnB
UdS6D4WUTftpKmm0b8GxCRg2Qto21IIngTkoxtG8yqS6ojpKpkQfgRfNS3NNmt/XsLGNaCY5r2Qw
qj1e6mN3dIkPQ3qXhHy7C6UdNjCqoEPnLi3TifJCkCvcKGW6UH6ypP4JBenJLWz15y7xUEFqdmD3
9hEp5V0UupUL7nD8/3PWqCTkvSk7ysinWhZpKpqMX88u2xhvAsJoK6PZuN32ApVLWGgOP1P0CFfg
n0KtpFKQzxTcn4cg0iehUlsM/ZYYJyzWL3ql0dLGCiduMrzj7NuAcJkRfRps8pAZMSx53HZ5RiTk
KqlwocuQixnnxWZblaAsfInq6/TUuoe8KobJfZAERzoc1PzNYjolqAhTEq87DCeA/4pY2HL4uJGl
uytMZruZc9cH3LacX7qAnVy7ISIlfQ5tLHYWSkAiYCw+7/N9zLY0k/I0k3kERVZJA5+VK9AU3C0r
Ru3sdNWhU2J+liezb+GFjmr8AzjWly6fg3cop7ANgsSBdIy+CNR96A5++3o8i6AC+x9shXrcpSfE
HARlKQFGNPcO6koBGOvg8/94B5hJEQZD2srh2paqaofA4SHEPMzQPckpxw1M3b2oSCEA6NQp/svI
RuTu5WeLHYMUzNufxFto+ApZcfyqJ8TAxXa0JO9VJBkklv5T09S9/Dtut2rot6lDA6rcNIn2zhQI
wcH2jYROEFM0o84lc0uGKTjFZf00zDX9hywVexsG2fMaVoM3IlonnHuHfmYPIufTgYgGHeQzGEFk
casHgpIwVOEuIonbhZ6WQ6uf0p79Gkwz8MuqCUtoRG5srm01jrI6NhGmCCsS7jo7A71lFkloVw+P
dQ+TffQufs+b71Hg1DWP5AKxCoWTVcLCalMeX01RE93Tm54LBmNpQJzoFLrTeSjHUeiY3X4wboaw
aUwJEEuE0whVqGZ5nK9qbgDpflgu7jkRC2e195XLhB5MR+fDOJhPOHCGt4oOE4zFnVptGXH82BzG
4Wl3GJ49eAKurWcg0SDiOD0KN73SDwhqAcNNBDZFfptstverjaO05sJJaOBE6ODYcYMoZPFfUPDM
J/xkunqEPD+7Wd+uPG6Vh/8wIFEVP7wvTQRY0toYq0SjI7ZmY/+t8xCc3hFc4YIUqe7hMcD94+qu
6WPD8IJiN1a+gIPMvPuvSV7q++fXdJMAC5dDMSNLC3VtXXEEaato6vevV4RQBtTf33Qkhei+oIQB
xt6EiDnGUKgrN9xS9tvswc74uU6WYi8dHcKkPF+fHzt7HdJgGQFwZ/0+5NcD/MmqwhQUkmkFfgJC
4i+q5e3htx/YqW4OXrVQgA5daGIhuC2WAmnbgYqfrv6q7KXARXkRBP8f1kQCo8Vd7JBXwxegazCE
lg4W6SnJShrc+Bdw1JVW8L72rbJdZNJ3wwHdwW2TSotDbzO651oqAUshmdqgHf9NujzUdIDwmMNI
HSYEEnUjw0s8h6f+bUo1FzMV2CIvUcJxU9pGlrOA6B3gkp7dUv22EQ4hMXibw+1hCc3lvg7lVqBo
W26KeOVD+C53Z/1Dmxky2H9JbfaV7g/aV2Di0iZAIO5UqY1BfannIzAyz6SXbvNpY91ow0ozKgTX
zYZGrGF1rnHIL6u2Ggt3zYnyQs5GWekYLKlTwZAvXBeVF/9x8eOj0AwIKs1smtTQIW1h6M5lMJIQ
roULt7TcDEBTTXeVvPRRYb9CBzl3Gbe42+Y5rMGDzHGynqBaAn0bV0u2rUCbTenwyQzYL1tKB3M5
fc4EVvRQqc9OqVwohXZrHlACEIO3eSUQ4KZz9WVaRX+Y4ZWe4i3iHj7xDJftL2a0ixDPKxdAu/Ks
KVYfWs6ICRskQQda3wrupudixe9L49vJGVEIOY3fPC1DPGAHQhBL/2cBFYnWExVakAeysrie+YRk
MOFf1RWuevzaMPrBNg+/hYzV2oYPg4B18JCqxB7TFzdltU84ix7RkrCqgZYkfu2GmN1mm5y7Rkbd
qdQO4H6IKRcKyNolm1zA444PYIvvlGQrjA2jG3Z15LcGM6sxJz5TPe0qkRsTZWbjMbXNN64Rw6Mi
GteRBqoizFDTdSgGKIzSBYkzzigkdIqvNWq7SEqcuDnjTOiF95jyVxrrx/dcYjd1rVcKx5MYR6Sy
ZVmdjRA2bRGxht+jyZDIqiQBCySJUxli/wKA+/8oYmkqs8xnvLd68w7qdDhuuWP+mfGBouU+z79Y
FQZ8AKazp6rrjupfRzIBQr35S53BypW/plkThqrHxHyY5/ptDpOtis197fdODqzUNE+MLw1eC3zf
pdumx0TJrWc/JdDYLmCTJSua3t1K3YZ9W6VJWrhCRlu2CoxrzPH3V6tcJp21MmqnmmDCL0Ak453b
2RAMSEUG+/+yERjo6H5fgEvAP8V7Hdam4Cvhj/y4cNlHcrL7aevSlFljd/7ij91gvZxB5flgJ9UD
9/34tgZ88ftJi4GtMlGy/63YX0NHLHeKH3HeQyZR/1FUzTu+oUEW00ylDwCkFVD7/HGUohGM6eSH
h94R52x06f9swpgrU+lkcKe+FD2qMP0WDNCxrtpCmhc83rmCYr4n12KylgC7pAfXFfqCWFbzgIr7
yO6Od/LMs+GLQ/pYCEGfV2InJwh+m6WWMfTy6Xzq0rUbLKIrQzwOEdAoN+UBLGhHgPglQQEJWcQJ
xjCbUxfJtkIo6wy9T7I7SEdWWD6mOfzRtZh/8SZ4taQ2/oFZ1DjhJLUISmMFfRzmjaSrH8fDpjLR
kG1G/FavmV/Ur1lXkfuczxVqap0lMbowyBZrZqKpX8i36X6+yFT4NYTPjCztx3O+EDNRAxP+mN4M
BGqJEhlIsRuHvBT1G4h/NrlELwKPHMonQokAYyv8xyrkLvauyg4YA4phsVh93TsslCwE0vpmWFow
XvYbAdYP6mJF7GepY/AtRqntH7UG+0r7cVNYey0nrrjFylbIQ/CDDztM/tgOBN30k8i2eCwigY3h
Nh/tugY8dvRyE52+WI0W7NfBfbbergMs1Ibvlr8dI4jDB4qd9W/rTeSduoAbrcUT18ylfkxdVi1g
wXeji996MNCIvaV15lj0l1XgaRLBxxT6ncrDOU28WpjVDV8r7V0l670HpJNfBXzv87gzsyQiZi8k
3E0IdyQSXeDpoehZF9xVPvhIxuoM4frJWvfNLJ4sA7CYNlCTAIS/XK0e5zZcYfcVni24kDPsx2pe
JBMzTBvOW+jeWX4JLHlFwoZoUnode7Nhs/nIr8cPanESJQdD2ow9J/ayGo2sW86/CSjhgtwITRw+
UjXz8YPO1Yx4qwO+pgGhOLYaTDQbHCQUGcFbV9yk/sKO3llcovm0ZqOagCrM/cE/DfcNOalnaHq2
ctj4EpieCOQ4M5ExQcIA/+mOTwJZ05gbkIdESzlx6GYAPCzcx4T/cYToRU8LNL2YXentFyQ64e/b
XlrY3T+qVUBAhGi3HGbPTkOSOavEPKvH8SuPCtrzhMT2nb56Ea2bDIspBNQNVl/AL9FBbp9I54O1
ckUIXDsPovYmA1XNSNPih1XSknqSHb2yXuBUImzch+NUy2TAG8/XN+8IczBP1nlz0NaWPaJDUZuN
Pac9WGhSNXzYruWION9ajDOfv52dEuDaf/TYFQfZUjh8XVPk1acYFFg4lJsL9dq0XFFbU5ITTq8k
dcLz/x8zliHbhPeNUWbj5DCaC8cZ6K6/d/2QFMw7B5Cywb+inWdpCemosFcEH7+/8E73I93brqCt
kpuv8JkKx3OrW4qqqRxkZFpvK2artq8HhSu52dmMn8iNTmgvDq/4qzsRAizFMq9dcLj3AfOxfMBh
hXH6RsB8S2NQzuV30LqI5weYGFBFqr7XGAY7bwhz7gkB56Nb2jETIuHgrLR/rA1Q7OhU1TmKRaiY
QD00FwJUIlMxR9Kb5rF38GCYy1l4MFexsoLEUbwRcf78naG0jOkvotxvJiJMnsChbu45D0MC1jxv
0ssXny5WV8D5fbC2S+24nDuxV/cpTk4q0fXX0perQFuAwfWySBCB8laJMFkF8X/PjtD/Cs0RpLYE
doEOnfSWVKkC3jNTZTTbxCxQvDPXnwY3PQMqcSlMexo77r3EP3V90B1TtO1431vXsNyBzL9+7N4w
OmGK/FooqR4h7yUnAzqIzjv5AxeBEpR8UoO3RjJkuihzwgQy21aINtkQh7dtOLwdcsax7ZZGCgh9
Q/8ZX75jIpTSc/KmzK0Y/4OPNmAjbOEUJLSTYuTNCq+eq4xgB4NRDDIoHE4JQH17vIKxQX+CF7jg
cGR4Z4E74JGJoAQomPTokLrBBHPjZh9Qz2bdbFrlbgFiU7epL6j/42BQkxQh6OgmilTisG9O2rBw
++s0V6tEbUFcU8HrxX8R8v2C1x6AqReEmII15PvB6BWAEWKL41pNHbVO2EcXeNUVGfI4gsxkDHsJ
0tii8bB6XejhdQ6rsfvtYHEBSWRzKl9PbGlFN5VxDWoBjeSuzgGHTJwDbxnYkTrrBF2NEkNqbNJ1
Fw61nSNT9vEL8GSBRXWmCMMCoFOQ3WQ9N6lXqVjS4bmZAIUFNGDkhiGnsBfK9wCRRCKlnNzFZnqr
bO6oigSPsSDrugiFNPp2wQAMrx/BjlnkhKDi9F7tcUi0Pd55aj3VYRbdLhYXnIp6xp+AH8mspBXd
k0+cRBTvSKqHJFSAEqpklzC31OmBMCB5xZ88plmoExhS9L2qUe/ENuL+MZ9gMD+fUj+l3bEDYlLc
ZyzIzUCwtGeQX0jwAOYlE9aP9xN0bMdiSu/iAf2XrIHU4wCtr7AQzlfEQUac8xQ1E60PzWLbQzTq
l+BR6CTt+/QJB+LsTVgTN7z77orVxo8++n2ziTdR15Svb1pCwPBlywB79UiT/TPhVo92VtbG/yRT
GzVMUsqBQGb4cde+lTpBz/a2gGxgISZjN6tiO2z6Nvqtno4mmrATNDKp+jJErC5w0ddhtVYUw5eP
8seY81xyRRzAU8rmvsOMcms4ntEgLF2AjpLNOL5bXRCHb2cMSOAgWDlq+V7PQhmPJVKnm0s3Ncmb
nW1WnP13pbXd+shyZIn1D2/F7CbQ9EpH1xKeP1k+qm2QdznZ7jJWCm2OD1ocmYDyXr25ylVhpyHr
sj+wlSc5sVAReiPAPqIvCygA1gQ9iYyZ60bvPAZYZqrOxa9kmdHokCtoSw6Nzu6xgxlJzOrYGX1t
JilHEmAOFCqADAjxnL24B+/kNNP2ZiBr5bMg0wUQR/KcwWp+/23xsGs+xuXg6lafmMmiqha2KRL/
41EaJ7k1wC/wH11ZX8kaFOD3HZsTvtyCh9D+NTOiEWDUg4FD8VeOcjQN5JDGGIt0Xm87MjQ2EDTl
4APMPLoaSFhKUBDGX0waZ4L6slKNVFQgdjGOL/4/eC3O/m2f/hSuCxiGD4I5NeHAHrhVdXLYQKDN
E3ATCdCMR1OERDEHAKwTiiBUIZtpGUIpAQXW6AGPeFSdDlTbJ/sYYS7eWjvTGYbvCIJgg679rMjA
i9xH59ScY06vgUQOzaCAPOAAB3+EBYbQdqNFFh4eiVMshUr+tptPAQo5zwV7pjsCQbY2QBtdWbBl
mtwFKWchWMziSw5vTIDWdKwPcbMUglZ9WY5yThUj6mGkb4w8XCuT0TJnbxWYOT25qQsAvih1xZo8
9SvRTWsZphPHPvggk5iJePUxJqwXDV8HQVouvCLdbWwd5A/JbG43zLqM9GcnRKO2GKNJqiGiDWzg
b9N6ehGYjj+xMzaBhYmjJTjSpr9SXmi6CvaIMZVCQP2vJFp4cZpZxPbByM87WYWQ8aNzg0c9I86u
iuHqRU8Pmmt8eztcm9vhs6gVZB1kL3zTuHgQC4NYyKNh72KpX5CEdHpfXHkfo5fus1Y4yGyYbeE8
Pp8CmyI+LY3I1cTFEcxmVZAkpq/zRcOqMRSXdRAwn/gMCxkHHRlQA33BjIvtIny+PGkXQ6A5LCHD
icBBABulBGOWnQSTQ0bqs3o5FS+MA7Baqi3e8T/kmelA3l/hZRVdaFC806z7NV6jyNTvwTruMEQ/
BFiKLOpRoYhe82Fzo68pOtEfvdxPaBW0TuNrihUN78eio0EoWd2N6nqM35Y7SsmKYi+vDRm2LYeT
mwEp8PfL58fENf9UL7t5S//FEHI6kK//EFL7K1wiB320VLKKootnHk5UeVwvASXZP6/Px4nEB4Eg
T3aJDkq7EDUtvI64ue9Lrr9G2KHFkPCcMs/kzfyrIo8yaYyolyGwdhOb28kESOi+AREyUD3+YsyZ
B22NQorS/1G33xq4mapfTlTdhFRRuQ1xbJLKJVawymjnQVexckEZh83wJ+9SaNDXgw6rn80UsELV
yNOWbFe+84q3g1UjFwICclADLDHYj64OsTlCEb0Oz4yhHnk+NzV7F7QylHqr0Uy9/3pb3y3tdAVI
SixfDNarFOipdQh5GOzSvBCkYdCFpo/bIQeKj8JotCPPi+0jWWZT1l4LTUa9annyzYGgLD9JFx38
jGk2X1fLsTWsG6asFzE/2y2uch8hzuYqTBVwnjmAJV7VMU0J21ExQ4qyMfGk6ojCz7SS9gTQsz5e
NDGK7s8Dby0IBbM2JqCvscmY/GisYYHiiPWZnrmEbVsbevVV6s4dLCi2UqXQa9HWZeBzFKG9d1rX
VxwGUxrah5Y6/FDtUkJx7BPHghvutBb0qWB1ctxGV8pZsgsZffuaeGCMBtMgdWHYxDzroAKYJ31e
pnlh/gpVhLgI5iXW828neOpHlWM7CHK53fW3vUcIeJlBFgSs9fQhJUTz2MJT3PC5azH1arMixf0X
JLIoFW13uC2njPd7cCDtYTefFsYq4duBzPuPqBotCFzetuUNeCnzWxhTVqVlgLf2ziJWHGJKqd4K
ZWAjLFQOPgsAGfGksxpluuY+5/f2oKj8r1/dEb96Y6S2OJt/3NZkOpqZSSfW8pvlY+VsBuGvtwBf
7RjNE+9MxhWLGMQAZYvAKUhyGZyM7n6wOIoTWTTXuktZIqdeKXvZeDrVaq+Gpu6LD4KGmuJVdXnP
78t6gi2rzfDk/nSfwDO+0S4Xw9g0uZ6+lVUb1mud+IG/SPgIZV9OOs34tOuqzVyLHDYOrw0hp012
oIk5Av/i1b4zdxNZNpMKgy7FPO6d6m8DOds6xb8Bj5/dO0G9nBzQUk5NQFn0YNhmfQKdG2so33FW
JCnv8kj9dH/l0bPPkqCnSPoH76fL9zwrt0IlzAR0mAXam6BMsbUNam0n+AuHO1V/U7xEAQQccL79
hh4DY3Wh/AH3PIUMORkU6VsPlDbNq30UE8CosPvJqhD5bmx5aSH7ioLNc7c6Ioe1kNWxDcR68lU6
WQAkGtwUn8y53edDqzpiRW5snk1TJpMD83Y1KKjekNpabriyN/poRTcnDNhS38PsewL31m60JRHe
U46owu9tAKOegUQQ/Gp2Y+sjSJOSTTjWrW4hq4BPsVoaF86NTKpcYhRgAIbf9vV1FBz9eobj6esU
iAWXjiE31yY+vDqlMwiMbdYiq49q9uNH+zPydLOFkI1XrnmaaiV2N8Afb5Ys4xBRGs5EnaLwz1pk
Cggm0XwQYeL+Vs5SujwCjQs08YuLdXmUxSnZDEha8y61Jgx+lm24cXYgi9zpliTa19dPNCEWEpzG
Rd94uHDt1aZTlk7ZJZG1qUSbl91tIVRXMmXkk2EG+mUMH8m1GoKCENjy5vcmobLSFkDDnr1OKCSg
oCWP8mkTQh1AF/zCcm4XR+EdzEX7uNwgi8PRv2x7BBpxP3CkxtnSlv7qCUoLPu1Q10WezvyoozMK
PQ5M9elBKzROyp71pC20YOR5jnIhs/JTQecNkPDZS520WyIFM59kkWVM682IOImAenKAy8/NPC6b
wRi8COH23nnrYxmj//yoj86oPNQ592r5Btk0nH0CwSKqRo4h5s9bW7eXlXMxRE0l0jOoThJm50cy
r9HFRN2WlhX3ywKNwbIdlJqEpl3JRnFbd/VV3I/qDk8LFF+dvNe0AUEt5w/oOiddmqHHWmZijVag
U891/otzvTb2OI7RJa+bU6jRa10Y5H9ua0VvNKMq3WSeg8WmRvhtZVYr3DpS3elXcMmhQCPYz3DP
AGaiH7NpvoSS2Ts8vA7PJNiGXotwvMFmQPGfAJ/22wUbXZKn0Ug8RPchXjkJis1f6Ln2KPRnVFIk
zi5HksR2RZ98oBaeSSNQg5v98N4kFm9k+ATcIm1soYiQi82PH/WlqRAAIO+li/Kc0+3lkozQRSAl
ay9fBCS2F1aFn+d8mu1j7W5A+MFTKLw+UFIThXUseK7vO+5DmKe9AQWUHujDuoGw9CTJ6sApjbKP
E6+eZDl0dHLYZHzD43FPKBgCsX9uO+Vxm7v+GVD0qofhTTuQTT2pTZMQhIPGlJkdes+RRpMUSOoT
QlWpxjcnwfCE/fSJ5TbT5Oh0MB5A3ZhJdXw6wefw1tRj4YrAKtWfKBE8sBAiFDOYiOpWxj/0neGV
9veiu7AAXx9Z9kICcdWQOKP1TLz07LtgOSeZiBQAbEVjwX3u6uhaK07GJsHVmd3F0DJkKlanalLT
CzCQDCpPzsOn17NRrnOG+fo2d2EZQd64E8Vd1hiiU7MwxDvRqWxBcKMN7O1vOlIKtrvy+smGgS9f
gU7EOPirJDGlWztMd+2oZc+VOGB1tlmQRzpLxdNlNP/Emb5TvjLqd6PJiKhTJ82EhN4P71CSQ1qZ
/gWWzng4u5+LhVowEMOQvbJBIwGEqr+VlTcIH10qAsOJD7r/mnqyaovxsXmTKy+MF4Ohp26QoZ1Q
w7PQOJV+klBhLLG3XAyLKkIk3C348xWhbPB3l+VyMzi9zRwca6oVbeOIP7U0dr/bmCz5RjLnw9RA
sCO5F68mLEKHKGT5ZPpW0bcLd9f3CFPkcg9pD/pacbR00/gDlZ0bnv3Skv/T3bhvMl/5qKy/XQEx
0zMgJY1MyCQtWwF1rblMficNfukKQCZl1wVZbziu52WqQjdY7hKTb4h+wFrfBTDmlyeKUp3npvZd
ToebQaVm1j1HXp/5vQQ7psQFF7bSU0TeaH3w6HYn5QfdgMLp9I8Sp6lVNmkNfrlEPIllYYxe7rd2
H0fVw1ugX5GipUX11Du/sKNYc5FTSKOABCteRw23ieUaroiwR6jq8NKpr7fOIJOYCSCaXFfFCL7r
E+x4wJMFMENVrybOTcco6zxlOzmzOpbCZb5bLxkFpjIflUEXxqNE5WfKXOqVnfYBtdmY2lujYo/E
aGJ58yhm+fe1UaC6kAvyMWhczxDoJT2G1U255mhhDgAmaV7G3tNAOHMOhNwWi8hM9z0ngm7AjLhV
bbN0DfRgkd8qiPsmSkw+zgx4eFIpZgOa96Uj1k5Vs3sLPFdxXRJZn2dRFZ3Hf9IUHKCHD5jUSpgN
A4d8joGXpEcp7qfTjmVEZB9quWb1bO8MV3g9UuFN4l6mhflyyjixT9a3P1uapFYXI76eKUfe6KDR
cSpQyq/OPWvUtuB0vfIlVb/OjKXf9sjaBytUbLBsxXRmZLlHyCdVvek8gSYWh+VhvG/nraH3pjO1
wdO9cYcT6nmJKcKexXyGkoPx2d6Nh3bkZ26zEXaqbO940lr89Mwfr/E3PAtEyDsEYx9u+DuyAe4X
TU4oNoAegPi9FIsVJ66SajUQxR2sszh4j0eCmoIXnmwZzEUclpABy19CeqgNuJN231VnfNoq/Yj2
sPSPGZdLYCuHPJqzG3eq9LEAyKBCm5YdT0pheAyRfkH4lKYIqTMJ+9KA9pCl4qo707Tk/B35Q7By
t140UtpcPibvyaAYyfadpS4XsPlBTcFwIUZOAk8B6PfhOYgvJnH1R/Cse6ZQl/YRnQPdP0ggCRoj
bbcmcAK6diBOh/orQ4nAswsqDHQpNUIwyoVWhH5t0AGNHWna9qZVhq0BYQNNb2J4Cg/kv2qGfiLf
+Vzi/nJjxx5jZEJB7EuDbp8IqabVIKZtn7SOmtXmt3jNdK96L3SjfkTQmernQSWV+G9K5MMZ5zyk
kONsqJBhXJf8VccYwI61sE/KjxVjFH9QKKNlQt/NjMEEh4x8KRci++BpEkoaa5FzWOfJz/CNa770
SJOpK02EL5RI6M7K7aZcPrqumzBOIcOd2Z1znOT1VLByb1Z8agZtMg2pVMUyCogdqAxGp5LmkINs
zY8c7x0U0nhaP7uvKU4CI+YJZJyqn/wA+ZAIjOiDShI9/PO9b9bWwLFF51f18bFyo3l9X5/qNyYj
HjBY2e3AZAYvMTYbO60Lp31RntlO3hxsUeB2YHgfCBs6Zo0EZ+TtjRU1Tx7EyQd+BqCvHXfwwI2N
mMpL77Gpmwh6WkFbQ5XJDeJ6pFSFBiDARcP2I6T1ziBio0BWNpExId14um+fBmvGyQ8IVlAKFMsX
e+i0jbpE+kOgz71esy/zfu1VniBiHC0Y+TxNCfn28gR11fsg8N53Q9i211gHiHzAMUQsokYhDTTk
ekzURhyf/wIruOkpI5be7Llti7s3F2nQfZYVc25tjy53CbFWEOIrMEU1ZE3iseFoilDX/IEwh3GT
8aEVID6cRX9OwMyz13S31hdqaLooxjTGio8HEXEacR7UoOplf+po0OguiXQVWL4jwqlXZlNowxv/
8dib0R6FiZJCA3THXWIwWUqadCMxZGXx0ucm5zkPws1Tgm4WzvFZgQL6+Tqgh6Q+eRVb27NQ7kY2
vUd1SOIjej7ZdxZgkBdiNhBbMCDFoR//BSlpWx4yF3IK6lTYsOjelqWsbTfgIxQj7O/se8TEMGqE
siyINn468c8TM51NxGGFHKcdc825wQrht0n12BDbXRYvOx9Gg1pef1/XLlqQ2NfbJww3xDa+MHz8
2We2VlbqZiyaF/SvIpNf4EbqQEuIiqKgWegAUC5lr4E7z9qwoAO4cOL9pGBr7fR6BREC9anXvZ1j
C98CADpUD+ogUfLG3IpAl8qfb9x1FEq/3IBsd2Kf5rQ+J1+plY4CfHA/AfIFG+lYtRRH0do2R82o
qnfA1aZYstK9z7z4IWCKa3OnZ+OEKfEkjwqdLWSMn+iXs5ch5562xumuTFa2ORoKJ9PMDAYWOQvd
Tixs+4V/ss4L0LNawc645d0BwDOE1o9CNDNm7Hmm3uR8X2VsryyoZ9BFLw7e33tUW6XzcPB7rIqY
pu2tX2/5hvKQ0xguZXIAxSdVkkXFft/xsXD1cMN4LSwrNQzJNnaJGAA6B2nHtnlZfahY5EcjzBHP
52N7GGFK8TsyMzUpQ2e+zVsomLkIKXZxBxi/lzKF0+KK5T7WJ9cgVn8tQfX9HFc0rcrI+zMTa9/2
+MtKYQULAanm8EfIuB7XAZC8mNm+/WTdiQ540lqD6qt21m0418OIg9pkWWCNP4nHnD2Y9MvK+iOQ
6/Lpw9MKzAOByfOrSJQUmZugPOTikRqT7+moYQjUEkzKeJOdZQVQEKx9RcwRztcCbjkmRoPixEKa
YjizRmbCHW5lyLnhUFLiHC7+1WoFIUmpsMd9AY4Uz+u3eUIR0AIyNd82Atjt5srG9yR93GyhqWEC
+u11+kWENAX/vgoUjh90QqxBLMOlMLywPEULcK26wM4gFCL7LDE6KRk/7jeGdT81K7jlgvWWb8k+
njMY5ccTRbwIlmHsOauF/b89VhtZ7lYX4mYZn3eHdoliPZF1mXL7q5EP0lztE8hKHWZex4ekKiUw
56XHdB/FEzzSKOJERoJZyE5YFT8TFlV6YpV52R7wI7mcO6ggRuOSsUqFFtIqxJAmfrYLIpCTq62d
9D+ct+4jChvV52NWwTQ90r78yoi/mx5Zg6pDwNsP1amUsnjjdkUzdF3BXyTYLAyzO2TjawdZcOWK
E/wmfFn5F0XrbDhuJ/x9Tywqt0hu72KVhl7zth/j5sEef7pZvufjLyWO6DI0et6aIa0jdGkSbqUD
9ziTJsjbeyDfGCSysBGyzSu8Hj7uY51PE272rvEWvadib2vIotwY9wFZ2xeCrYqskoRqeOm4A4vk
DwBzB4291tLam2aNtZ+4ijVFCfh1zo0vNin2egfgUKglh34JFuqodod/f0CY3oOoSPy8nAS7GhOM
LHdYAeVQUPlWCQAYpw4//baSU6dbqxmDtYoINVC2yru/sM7suMV9kgzSDWOLbMsnHfCGjwEg4sQJ
5+etPcaBSdNyVvwk9aWRIbqsSvhUAXO6eBJYLS5nQRNoB6fpBM/PzmbWmrbgAtn7TB1kJEOCvm46
zvB1wx3q1wJ6N1XKv3UWmRSeCUxT3KwwPqFxNDwFPUbfiEDqOGhtm/RNvCa9vNTejMegVXJhp9rC
MQxBD0+OB/gzn6LLy+FlEWn6C4u9HUB6A2V8BW1Nza7AuPDrVRIX0lADjckXbSvg97SUicZTMjL9
LIntKhVHhRgI4RO7NZI6A6fpLo5qLEspqe7nUGmKFYLWLCmrBFML6DY9RD6Zfbf/PDpYjbr3k14A
/vto2FjnNTKxIwa0gjU+bfxlpAzRoYh4xt3HAtzvck2tZyejcJ0g3bds/ls3IKIijwhC0PqxdLpD
ZoW/meEwmrXKFvtiCZHihWYfiOjRohL+P8dBfGM74jso9zRexrk+DhsPwLaj2fVz61q9wCXqdg1H
w8dCGgMLqdjOD25mz6WvoYdQayE4wmdEw2M4kUR9cYyjoWGStwTMio33YnJTU+3+XpjOcbfva/FZ
88roF490rUPYcA1eFwJyM1jstZiRj0x5fWmvEF9gxuWXDc5x929mL+vVcSwqutjl5/Z97FgRlTx3
mx//Hhc95AD/J1DvUug89acPz+9CxykME4Wk9ZLsREJdEZC1IubE9jdT2yQTmUK9Al/+adR/3WHw
W86xSfD7oDHLiX5KXisgiVEgO+SkCQu4pl5tUysO4FnlnxAS82VnzSTZYsSyWX1x15tZDhydWSA9
Qk8lEXWCMtXtzU+nggVNL8ayIgIZOb+aVl2BkhXpEK34cNcO5MBPTnwwP+93lhE2qLFiom7OIemT
jp7LMdzQylNccFIs+KcJKR13VLTUUd0d4ec229BcunGv6TrrsIUh6Rzcj44Xt8N60GKe7+G2hvQG
Od0z5GGGnTkYUm95BBmthA9m6/4GK2q9ntZL8SY2Vmo1wU6h+rt4qnGleIN5gOHBalrJSSK2f3uR
cUpQ12sCWtCvS5vLNbIGLlT5CttroZOic2Isv2tWghZHTDd3EUPzLjKDeqmnUHoutOia5vqPgHDo
UHhHkC8lU2SHX00yr3fSipuY8jNCxIgcyw6mv737hiocKdWYBgi88CIQXI+Zks0zzvyZmSWrKFkQ
yhu2LvHdc635RxR9wnW4v4ivwG4aTIW3Pa5ZD5vEa8mwAfijQyGURNXr4PWSGDPxbDZ4c+iWNkuI
RgIw8Ek9GFwZNjcBuDFuQRzaIzhKN63gSIXUmnSPK6E3ExPqBsAaNBqeUuNlw8ssKwg2sE2b7gJr
P6ZU11n+TBXmtP3Npi6UaRDMLM+8zJhGF4oRCLuzH9OclVsrj+Ldcq1so/0pqdZY7/fXmsaMDsby
dJsmzPYfSrJR/dJwusC9p4MyaE0Xodn5yXw2p8FR70Pl/eOlyiddw49isCoHCjsFxbVwULJEyVCu
wvbfW7g5En2hHRBd7lsK9lJ4spESTcdx0X467gmhCGJiXmWj+8wGdbdK2q1wckJu8r6LHuYc4FwE
Xe37vH/qyRtMMJerDjWQBWM4V6wJEIQMcFM+dcw2BNg62YrYJeNcn2uD1237prVeCuO8nnEkn0TH
aXb13GNaWMx1/GUzbQwMqd6jjDE/E6Iqu1e8/GrcTq2zi/1VOym/CMckBA3lo1wryGdnWUEGc933
ekG1atSp24iKjjbYrVMbHgKNXYOpH4pjTpusjc+dpsnH6kgEQewplfe/4LYmci4BisAUotT6c/Kn
aidF7JcY1sNZL7HiEpOssf6B+eRSMBam4R2zKZGE739qFedH2BhtEicD1tvC4UcPzjcIrmypYY36
LBNrKfXAJYLaQMiUlTxZzf0F0A1+0p9HU7ogjFzCBsVahlV8LQ330TybCVFcfIbl3sY0cKKn5HpN
2Rou4FCt51LtDqzkTcppJvU6gVbfg+C5ENqYvB6bOEAQBkqwhMbWFz6B2gEmClJobb4y0fEBWymS
9C6hU3DjZ5lGOIEM8mCt1o5MXEJYpjeCTRK6bbwAyd+ZKgfwRQ3c4qMM4yfkHh4Z5p2YgeJrekNM
u1o728bYLNXNbbfpIo2wKGm/1UO9brYzqNDz0kzw5nHsexxEf6LwrH9BVXImpRiPytiulKsJMib/
vELJOw7QwyYpe1QTklUmTgPjZVDHRUzEjI1UTTj3f2DHXBW9bGefNz28l4PLKd5m46ZP8ceWTt6F
oirhVITcFyFAkwyhp7utyNEceu9EubrfwnQml5lHH9af8Vn9A5/aXq0dxh5MtkHp/dspEEfi7hz0
V0K3OggNJDKPMf1jbtRLDCj0Tm1Fzp1FrD1VzzDCVMhUXgS3RF2TTFHSPkPDvFTltV6FlF+6alZI
DOLvtR5KzlS/W7ZImKHaiDEaEjcnYeDMlGswGU2uYNzgh5FUT93duTERTq5p46kEDsPV8l7ZClQs
RDWP+Ujh36N1xAEadV5oGnZ86gZeL5TeXTrKpVw0t5xlt6qtHdzX8s3F8xYg2V03TPuNmhH6kmer
vXjZI3A5OWYkWNvcOYSo0XBCqhFv5sBnc3TrctyTEct3lshmXvanZXuZWkKLmkXq5w1VKoLx8DR3
oJReRQtqAyvLIqjbil6JrI2pt6vnfQV5TB8KqCl5knd/D1xWENgvODNEBcM5XSFqe7Euzud54aY5
oIE05vyIwPoFrcHH1wAyAFuNHdX2BTGwiUXlUweJTTNDKdegFZfAYOK8GFZ+A0cWv3fHYfeFzEj+
rvwoKoxwf5b/q5ByX1Jn8XEJbbgo4tIugJedz2J8UJHDM3VzeOIjAzSRlkfhUTezYAahtvoOH3Fz
3LR+WhaS0VbZUoUFKja22IU1RqffSTE7hgTkENNUiBXPDZin1jAuzBM+qSYeM/imq6ugVHzsmwpL
PW2FKnnm/tBWdvKZVu833lRmbSVt8+LNGXdp08oJCqa0YA8RSHYBB36qU7JUM1ezCgRBLWfoxHK+
axKTeglXr2ebvPSDe0fzKQ8/dz8b80c0yYFRnkop87Cy2mFQ244/OM9C6ur8435n8YFjV3ZFH8up
F0ZpUXBvhtlJJL0QKfADMjpcF+XdZOZ+p5kvX2UNT6nZPta1VXp4Auj0NCcEGMg8uTd5zS3ZLOLQ
Z8OJygNWRjaFhtFCbmDsNoCbZy5RaWQyPe7WP137657NCKIA74nVT4LQr+tZV+Q4fuDNrdX4EY5y
IyAFr0i6ahQTNPIPeN51nKWEJR+Wp6Syhwg2ra1QZUuLTC2n52IaVTs5nYw3hO/p/rUKf3NiIRRm
EepBB73Bd05HhcDyIoJ8hZTCS2gqy5qrnGEFk66vDBqeBJgM560Oyk9UdGrtTOw2bTiHOqkVKCKh
rS6C3rffdjD0XsM5iCxIdBw7ofIzCx442xoNinjlGmJrf7/PVOg//AwXuR5RmQq+ygSPFpiKzNjV
mTJJVs4Ura52gfV7oU8wL4crjhOiFJEsJhIUCYRpQJAJHGsfw5rWINymmKTVXfy+HJmbhv0k+uFa
NPnrFpCT+ej9yTS3yLgQqjE08mkI7acFMCl/IrvTvRciDuGSHBF0xOjvVfVne2Ww7Z14ghz8/tjr
Pbc4C4xjQL3M9yVPKGksiJGp+tG/jeRvwMfloZr5+7v0edElzS5iNe2uNKGixoluf/U3y6hxC9K8
cYXFoLQtuarb6uSt0a9C0TqeJOChGqlBKKjpx3MWO9I2yOWIHg5mU6i8moqlToJh+Leyl55eeLXC
PhCPSZ+PxOzZEeri4kwsEQjmz7pz7v4B+PzvexPmHsCUTBQx7RF2S+YdYiUG8IzH/s/Rv6PLAMKt
p3EMKDWhyJK+FJTGe0ppY/LPiT01KEQohItiYtLgVQzqxYpFm+WiYmx42pKx2ZtVe4UKaxd3323e
qMOT4MAoeswskFAN8mv3gFb3lVPgl4qGdQPB+8Q/EygvJcXu4zNgPj/1MRjUVpjekN9pJpEOQgVW
Zczkh/Gnulk0wTp89f1pkFsLhIk77zfsvYVvQd2Fi+J2Vuhz8fvgWQ7++mix4pZuP4KZbcRcaaqc
9izVXHEUWh2m3I7BSJgGYPJzcGnA291Z8r+JKQben7WyNFa0uPW8OToQXRtMyueWFe1hi0gQ4nBQ
K7ObMqghTTYyU+4GhnwlEpnXr6walUYc8IUs+1B5Ilje5lGuXKSFiNBCBmLYSwo+2LDtp/cajNqp
9PlJTMFmOGlHFgS0zON843DkuZEFgB2NRDPprUyQ987lbmNrS0/bWePlUUGYULDizWbJP/TthOz8
JyVdvutXKxjCW6FkqFiheTB165JaD4LB/3GHxeL6M55fv6NGvK+POA4aP6f6xXJJYdE8g6STZpvs
BFiXpSDPSvlTOQTHoSBrk9t9WCKJUZb9rhz7PFywR5sDzc/Ntv8ZOwKKYm6OLfF4hQ1ZkQue1l+R
WhKU7mTkfa1WBurUDxs3VRdVsH9ZLoqSLNdo9tHjgbJjURzflJisaGEE8d/ZGWOr+nv0OCLq1IAb
XLwkOHi8u9tsRX7sD9XKg8G0WTUu/nTAQ5hjuSO7ONCu5yjlZz6IHdUcringGL2bOzyQN4+OqQO5
DiZLpc6qfSoj3Da2L5dMc5devOKDsonFSiOAHErVIhebpWPNX1bDeqvWcSeLq9OAHH9u/H7LHlaB
63jmLVa9Io8wiNjw2QGaL48UPugiPBAGhhUAP4W7uVFp7cEgCMGc7Vi60ZqrA0EshOnvs4Zr9xs0
Oq2wgp9reX0k6CYkHOxe/nzzx7ffdflBQ2+qR1MMd14Hgxqf2it7VM6j4Fj7RHHZ+C7tgj9SAYzN
r3zceRI4kfnpa9vEelrAwcTCuLbK9Uq5A76gbiogrgnQNX0SNkhG7/ixjdNPRTxyUPoDEJlBeo15
M5J17n5pQF/k/CPxbW0HaecN3bZh6CGOwfdHvFxgWieTnqI2hg1B2UnZl2WEYHaRBuczXdjBPBNe
0xhUgQxHAS9eMDuSSzDZqKx6wXJX+8kXBKf82aJyKQC7vNKqczjweoSk3rBcvQyVdk3uEI1tPS+W
g2sWQ8hJGuQqE7yjiCTtcrYUdZszP1gZFnuksfbCC+nPY8FAey5sIIbSh4msm+x35KbZajCofodC
ywXGlcxjO5jQKZnDYdJEVuqom9DVPsuMf8DBjfRrqwncyDuAvaC/BfhH73GcZ5pEb0eB8oyFo8Nr
OvHo3NQTSddzv2w6HLs0E4oskvhD/OxWdlfKgP0xrE6A7q/Z9m/fYpTE3HBkCCCnwwWBOTsymen4
Clvt2FR8jLsqIE6iW6cU/UlCO2tj+LUX/a+To7e5JBdAptHW9fXTGHIHFRDUImzE7vJCF85M/YcD
sV3roYap1Sl3vd/DK4ermaS3XCt/I0upJr1sd599kGuFiezZkMwXYHtFatqkVjOmiqDSkJ2XCyr8
1LI2IB4IGZjky1IzjNYWk36SGpgphQsPGq7G02w23bKSDhgcjaCGuucg8tMp/DHjLKkZY6DEk/N3
HIteoZBp7/MDc16HkhVexRGf2IGBqiCME4cTv5AIL7Y4W1MUvUKQmu4S7pSpMiZwe7xld37oFm4Y
B1U+s/wU+jF2aXSGOZwWY4e5TcfTAb/OOb7gavq0lH+HysosH2WdDpmjhJU6DBG3L6AGEz/xqrc7
lFiyb+Eihb1CsdOcTbuklT4g4KpQD2JmeUqOoI8X2WkrFRCQWHslhfizpM8zl/6B/RrcxosLT5mi
fpHl/Or1Frh0alPukirHMGxj4rMuXMab3yspgoF8Z86aa+/sr9yYl2hXCIghYq8dG6wCxPOSd9tr
6vNQJmMLBfKbDZ/j1pJZJp2NCVfUGdxSuCE93Y6J8Y+6LVQF5/NWABBR59qJBotUVlCpG6i+raOl
xAYj+GFTW6oCTXESabqvZMdpgq4WEvWrRtL24VxFqUURu2148gfmKHMzAviAYmp/6SFqeYnqKm0k
tv75jFXzJAUCn/T1sa0vDDrZflIXDTa2P8J4is61sVwByEap6//nNlPpOfa/zrwLSW+FPYZdvumw
rzJK4LYbukgHYydYQgzK3v1Yaj5oFROoNbSQpR0wRaS13lNS7r8HOKK8wC2LIJ1ot0h61BuNCm1p
xm96zwAQ50RgpIe5GpOHgX5vLSx2JKcg32yPFQGPoye9ApoptWwCeWV5gXKTv79Xo1YIvRRGODeM
TIpHsRW3bloCYnWxHoXSuqarxlDckUN4i8ySB9VA4nGSPiDIs2mDbG0rVhebjh3HzoxCGZGJoAzx
eY23PW3kGuDr2kSZ6ayT3S/DuadgiqYfxMbRA0udBbr3s1ZJgsVRXDczL7sRawCL1MTzk0kwFdFV
o+xHu+l1XO6kXQBgu54h6yXMeUp8AMV2ekbEEBox6yMvSq2QFfBWz7JixTO2aykWGfAND2wjwexe
YzwviisSYbos8g5j8GdsYY2lD2DS4UHOKBg/JYSGULtrvqJ/VH5Jwl1DHuLtkIlFeCfieizziEHj
pQzSPrInTkcubq9VtSWDJpiLEsnEfPkS46B10jsLpos9x1UUcPBY1E40QBYwc6C1hI4V0LRfECw6
qMyVFb7FQy7/DCS2Hwp1XzqnjPXC2/bE9fMLUTMju58+0TzWoN7z3gGl8AvorYCKiiUjlenhFEOI
THbRNJJxo087xWs/NGdvffjUp9IpCkpv7sa+wP7ZtDWuK2+7ee0dpuiET504BeOMVRsM92hrt6sD
fF3EZgJsQh3cRCOcHZS2gyTJw6QSoPB5yjgb2rxz6svW59PDNHbD/EDp3l8/oUyw5a0CUd4EaQbd
i635tw889lRgnzZIhPNmXwnHnXMX/c+V44t9rD0WgLnuThhrK+L9fTHEhBvhPerQMcyuy1+6yVpM
/TS2MrgM1n8pOndwihPRcH6DFwY7hFDVa5eH7N2fk6viSop96qKdB17GINYz/oP2W60Gzxcu+q6/
BUFLn34Na3nHIaEw1eQHUKms85mx8OYFrhr/pxYOtQbFxOha/PIp2EwaMP3U514GwQZc4yhDmtRe
xzyLy7TFYyo7PkAD1CssqSGmtMJDZMCZf6SW6Q34CQ4p7UqWF7FVbsbb06/hxXQgbgfs2J3eHu0y
mCzRH8V6x8ghaWI0eVDGjaKzWZsdRb316cPRwPY08JGwMsogcMpotg6iunMCr8jqe9lKL0cmlsSt
pj71YOca7Zz9eNgdkiLnNLdSQ22shksAncNaAJot8LV8OpHyHvXIHptvcyPrlMLsh1YMp3eS9GE7
WIk0M4RbY/GboVXqy2bcj29xJJIB8SauPXckyYQiccCTspg8CRLhfIw0r82kH74oZB4viYfa4B/s
Kl6b4rhL/dPBhSSXvb67e7CHrZY1P4seANyR4i/HeVxQHo2D4MDEs8UMp+6BBEq8W4L8pYGHWc8P
3ygKDdEZ5D3h53Qg9bUl5NfZY3xqHS5NC1V8gl+sZUjr2Ca1h7UzCuHG7hNVrLc+ZY5/h9O6upa6
JkCphXnsaQ89otvWV/413k2DnHxRacshsToJ6UvHiW89NG8XxavpwZ6Si11eYrpV5jb+w4ViJFGu
N7figcDceDWsFtMLtRQSu8NYBwPPwDzPs+8H9WLrnNOg0bblgRNc++qN8RcbBWE+A2PucgUtqOdB
/1cN7qVReJ+hprt6aSC1GokoKoA8RI0upyxWG/pQ0dLG5hosLhGhkk5aGqbd8MyUayc8fgiKwXuy
Tf1hOU7oeN6K/b96O3nNKNMCL/e5SIB/VgJGa8sZpqxcn1gITIGtuEZWcMPx/Q+XfjXWhOwcrWVX
0aUq0MNpBkEqDMd+SaunSwkJAotRnKD4nYu7X9vf7JMEdi2CIyskG1YZW3Ct+nHT6gPcNkmqJRa/
9vmUJLi2EgDbx/TDitF4tcLBRkC4IBtsRXBWTP1MhqEjW7eHBkfdhteyfZKxp4IQgjaXXz56cEzV
X/+f/UA9+iL/Gah7FxRAek5/fxwXiHiUMcz2y4XO+qNYYi+ciimx+4BL1LtD9040phlKfDn6m4R4
d4Iut0bSzBFTP2XxDJ0jImS9dY2U2jTkxHFMS50sIrQCGDGuB1XotuhRXJaF5KbIr5TPHkHouPsf
WrGZ1elp2l6qz4xTbGyFzIyY7lrthYaPnA/qRJdm3BwA0ZTF2duYwOBQEys4fjcDBloducQ8NXRk
a/GK3SbdlIuBs2f3BcHifprZ7huwwEUk39pUgA8T8itPjPMc9676IcsE49iCdCy0I3I2KC9+tDoW
StzLCwIFWFCSRKF2SuGoPu+USjQPvZB7wCZ4Bh0S5wTDhPvpCQjQbnxrvwBVPDbCweMGII9Mr5yC
XCx8YRO19zoIKPkrCNZUcQ1iArT+SgbSoQE4wbAJZg7+DWT6Uu8bGj3xA4zDRVGfNipZClSXhQSc
rYBaKTgxwcD0oihdHKguz4A6fpm8WSfCv9bDsRYviDfJgMW7MHEn7aLyBrZCussMr5J2t7ey4rfW
QV95llKlp3KGmpgqotQIDVcXwdTPAjGIkjG/GiE6LLEvXkhEbiegk5lCuYOqBoXr1je/u/8FI1Cs
qlhqtGe+BEgYkW3pB6EDsaT22zp2meZwFrgHyglohhgX7F+nvqsMyAAx4iidFvK2KDakVZAtP/Sc
Ipf5ADKmSSWdxTVA9eLAd9GczAnPGGHvBJ4shMJFgyZiYuY9jW8Qs1ojOy8pjz1wej+4seQxaTuU
CnhYZPgji8VqFrEM/TS84rKkHEsL+BZ7B3CM4tR8UsBVa9tY1nmoSbamr+PRnxhzvdxtH1VIBhlu
NrJ6MyRoRIWU84bZKsA5yTF7GgcuEhCS3cVqoPkbJKWsutZMwau0TtH4spjWC6QYuyOe7DOwuI1/
kFMw6300E3+boqYNlQgOFM9fMj8tj/bi5ws4OEuftC1tQVyhxCIfpSHA1wRc/ikBbhrk/BxoafNJ
lrXmSUQCmpFWC8tRXpXwXA2i1yKLxTUEeQDUhkeC/4WhA+iuMvT6UWdq9bT0hELp2yHi0ShnS6m3
vtQaX+sMrVHaSubHwVkPA74qOGDrQ7sDLeb26r4TyxR1riTlcg5zjHJhxf+GMs6cgaBCbR4jloci
j+tzpZay/5jUhcxsiKqPOsfJE1F5gCchi9H8CzxDEobAfSmpRfNREwWe68QR0kdXSkWgBmLRyRpe
lCHVmML01YCbI8CatAoBPWnKymkioaOCtI1o0Giz/EwMfkTcUcKK/fzO3u1zno/sVRFVgDi2rGta
41Yr9J8CvZAYafqZfAG6R/mPlRGDyETm07QE4zDOnc7uOnQhj62sbQ7JL5TbME4aP50dipxn2+Mu
dwWCaIzpgL3H9dZ8Jtfbwh3T8Vc12FIhldPXRpfEkHwsjzEH/BSYSsZ9rcVGgGeAshYih5T3Eoq0
H5TJpUppuRAotJcZCukTClK32eq/+eLJMteBnW5ddSiEvxebRCpmqSxCT71+29VlAUXMGClw/DBD
NZCSnTmDhuPJvX63q4RhEzkrqesSXW1OkqeSVoFG5MyQp7/GeL7vwIqza0OMsv1aBjVOau6Lq+Nu
2HBO6sNergCDUPJaqc4jl4X6O6Jdl5fpcZR5P3Vi0aFhXI7UhynDSSYWcMLM+XmP96tzaWlduQ2m
NNExsdErKhyx1hj6nT0vSZuTpab0HJAWZWD9PulGx52cACHF2nTPZpY7Nnj0L5zfiOo5i3p2S6CD
4/EBvnvLt4umhYgrQBsMtuXqcp9oQOs8NJCWarjlJANVGsARTTbMK+EVKZ3X6cAUB3/+f4fdMBjc
rWnk29h9fHhaAhLbBGH2f3xN8pePXuu5Fg/+kd6nHoBTphvtJ3nVLKC+P2KaC4s2rCeD+7Rld4BK
HXqVfp30VvUsGZYsJ8cl5BE1gZ62gu8mUDUKA1ODK+iA/j4Sox1eGwCtLJIUb4Aqfbf9ilDiVoRj
EOEAPwsLCRxc0ZSp31D0yrlVtKuIKeRthCU67Msqk3vmWBP7LhV0VlCgPYQJp+UGIb5WhlzOJzj+
Z4SH/yqLq48QAHcHZRPIqJlMwkXdvCVr9cZgxtun01mijGp075CtX62hKkObjgO+OFfntFGvd8rp
oSF6OUOWg3Gt36tOFCjbZnSU0gWsaaT83JSE0S8fjEialKJFtD/2rqgXBIxvS1XFHczs5nsY6BT+
pVhz5rlIMAe0XtXttQ2nwGM7fVGBJrC3Pqy+6SrOTSr6hXNd2Dar8l7joP79X4/avJobYQ0TeR6u
sF0h9ir0ToAq1lqV9qHB8y0o/guRzHOPY1yovebnZc44nnOZfvOIUJW6FQ3n4iP0v9sQsgnXE42t
+riEudl6I7whfrNAN5DySRL+wVPFybtxoRvlp1j91+4Ale8oO79gVAenIg8ryuoITyAahDmwsyfh
pjARUxk2iieaoaDJe6Vuaer3+iT0IkDP/TVaPZ6RM/AXj2dRi9vyy2SZwLuSkC0ec1lfKxT5YaXp
LmUiyl2ZxGjqnWe2o3i/Mv1HpgTixdD9IcfMKp3aaKlkigiwvJKoz118fdpdCtC67p9fr5s0nhYy
iru/SXAJvQlX0QcbyFmBF17ihbzUEP+NVn4+wdiwXik+GjFSFwW9DEhQoFprLffEflVMmMeIPGgD
Y0fULSRylX9pYghRH5eoQ5Uzx6YndXgA/XiTOSpxcPIKuvn+hynCicdaK5/jzOLyMw6bKY3UyAuF
Y7tUjJu+DbKkUPebfOntW1iPfxizLn/9ySoFSvNiQbB4ZoqnG/X/D6gq+pn9ZhqzzUKWzjVdSiUE
Zn4dpnoVcwXo7ykVCH0Y0meF0341xf8VIJ0UJEyUAKgKwP8PxB+js1c3UkRwQj77649mo1sLjGmr
/B8GUTJ0qAAQMeCPwXwBMzanwpVT947pmwHWs8/1lH+MbhBI6U2WryeYJTLEGMSMCkEyrKlEJwe2
RtvstB40hFibSXNlU20Sqdq5e3Ouocs5KDiOlPG5JCrL+Tt4Lk48xWCufHOq3oMeOi1crG9s2xZm
6odVVFWeQNFDBKwmOueU/1f+N7ebAacjWmWxpzAtjQupUDvQyyGUMG5gDrNBfchnB4Nd7TXRD7Lc
3Gkk9C9r3baEpMyYgvsWolRxmRWdIS4xGIybPkYltCjVrJ3aeUDavRuTVJwQcPSHRHcT8SSrwTNy
a393icihn6UOCq1zaL4/c9F3X1nHEr3kAk04oB2OnA8mM/hM29796VWt+iXnfH1/ma9P7RcUJHjH
IihJibT9tC3O/Myq4k1o6Vtg9M0CnS3WAuljuRIB28/xehyWY8DmEtmGX6x+RahbkT2Y5r+yOXWP
KGIqbWKkuLMf9jSSqgeF0gzzFuvBCee77JO0lUeqo6cObQY4u0rfzT/5Lr7QuJeoVLDGM4LxwZkI
kB49aqsQg+9BNgfg8aMANIh6PIPYuOgt8lpU+NRRA+roYzuBz+z1br4pLCfa09ZmDqXogJHfKUZJ
mGv7m64iKxxVZd6VMrbPwNp6P9MxizXFLFwHtkzR0/eZf9hiuuGz9sZY2i41g8glZ031yI9Bzta2
0Yobs0VHVglDcPbXujKygjyofmDB6VUDn4EDSrPo5HQuImHw1sTIagpfvBGytpiNq5XY2CxCYEyy
9RCEugOAuSfkaoXdav/0RJZ075vvYEvgAclZT0+ee5/B5Gm7oL9Ome7qYhof8ttClbzWNpKxq1XL
Eb4656r3zn9Ob5FZe8/bnP6o7rcRnxh1GWdN25nQ+0MwFY5mLhfAhSzI9ps1IyQVpM5UpohzcjwT
5oBuei0rpAJHr30PfuVEHEc9li8ukiOpVjGYn5fHET6UD4fZOk9T8k2gflc/Izf6rz02Lh/nt84x
XAP6k1mWfHQoSuk+WXHn2OHNljTl5tCZkuOXC07QFK+4VGhF+6U/k5RI6MGtO/cklg0X9lEL5y/U
AX8sdknJI9SBS0Ix2uiAJ5NRim6T27RMTCs+Umh0CRSudfRU0GbZK+Kis0MHBM9yoNwxCGTtcR31
8EoErE7frAo5Kye0fIVtZHCTnXgvCZ+oZ3EzxNUl3GaOCKnvMHA1SZvbmWcPNkMz3Owqy/W2QZKr
o7y3Q2JxTuXGtxuL9NHe2mX4mBpl7zBHq1DvSdYhKL89x7sYpi+n6r+MxAQmDc5TITdrSRbP2Za9
w/8a0btIZNmK6J2m9pz6/LnebZb/jbgDd/B+aBSvYehoMpUQdICUH4atNw6SDsFxb3rKwJylfF31
S3hJ1XhWRys4MMdv5/3xmXct0eKxDwIfXWHMwwegpLWx9pl3VHNrkrzg/XdYw6IeJaJ+pN0XCq8o
InQiKSJ+XdTkbq8Mltgsev3E+x7f2jyOgPBY44SgN6FEbtee1Izmr6/uyV/kbEW1ScZyvTiMU7es
lLMlgingD0mxkeF3GVMPFXFPTvieZjreSeVRMO+jRzUelXyUE6CtkEyXgdDxSxXhSZ26wt7GGgfX
2boJbyKlK41CpAtW0Xq9hy9amQqd9tI/d7ed5M7+Uh9jSRddFLoSYyGuvCMRYxgc1PcDT4AzrSSH
PLro/kT3hhOC1kcZOwEfRXHAnhsjrICkGsfM7iDJnN2EVH3lb14QCSMb5W9mhjHMeqtxzLVW8N4h
f0zy6KMdjZjLDxnvi+uzjm+oOikks+dekPpq2LfzWrwk7dE+pisW2G833+m88zhVDCEYTIaormGl
wWQDYXmpOxqarbH/Ixz90GwfzNPl9PH/jA76KIQmKo39lMxbgC2pDsRkXLvyUbvryufQuzdkznEZ
cj0uswlWXpkceh4GIC6S1n8nYxFzLfZMPXATJlA+WOLKlf8/dWjBiIwVp+fdsCocY6xPFCh2zRZ6
2SpBwlznbItC6arCRX+YWdkOrFYj5WnplwQKYnKxLekV8CKtuWMI+hNUg7CK4poMNpfaX75iywvB
W6bmm33CnDqnVKkQRCypl6hNmC3ukxcpf1cirTyreXlk/nTk4nHDJ5R8ucEd4uy4RFtNokbL1Lo8
rarlZTUd/aYqMwcivPamkeT9MiuPb5xaMZCwbn9jJ1Nzvj4U25ogGW90snBtpgxI9G3DYfmD1tDW
MI5gj63iEGGi+pl1s1kKDGhudxuqslVQFTx1euwKU6MfjawK+Bl17qu8wLYKxR9GZjoJPYM2oWU0
a6PQmQOGwomgfqU3Ytv7jSdbdvSTvvAqArNkt3EaXXMQTLY+mdriKWgT82ex3vDpnIlDikMnUfD0
PlgRrA/aYQmnGFlRT0w4xaHH+z3erKIlhaEmmMo3Mfltxn/KaeESCZkMeCtQ2TPNH3rQVT0YyLdH
38xr5/bOWbnd1bEYF11MMzCt4a63bwVChfTLVC/nDw+0lu8srqqt9fdvrAzB5KlY3bV8bQFTTLFV
c4hgSwtU2hx+H6cBqyNyKZ5+6SZocWQHft5yc+lT1juPEz1ERGx49SUBf0JZreT07G8WpAa+6V1I
SCOa1pXezM9b3Ol+EmwiRFnm6tmEQLx4mBAdbS++5eYVxQvxrm65QZwESS/MCnNkCk1pGEE2Rjtt
NGHJmcycK+lZiyIZWRjcejsQ/6nigVJXM0y9DLvPVTBmlWR6sWadXwq77ZoVJ0a1WeFEMrAZCrdo
ycpJQq3GLJiaJvyysq1ve6H2XpHinDZtrNNiz0iY7AwCoG0tckeOetVJnUt+qDsj4Q0myZNGMuJO
kpIaZDSh0NvYEimY6Px0xBIwPLlSWenj04Po4k9dwnJmJvSx+/3P5qo69vXR38wFz/mMixTeHSsS
rrfYI/xUFePdMHSjL6LSF3qaMZR4OhiEfkqAeRypfkpYBXAW1+w3NSPB2lNoNBeZtFubEimocrhJ
u73ml4V9lVbgJO8kACnNUaq/mbjqBHLYOcdmufjla62t1jWhw5ZZR5axUMKMZToXiD2/KFqACKbq
8UfuKgpNVfFrtqXwoV86mKNNlVICytW95BO6vP5ckW4BBjBhCFUZaJLmU03SlqSaIvVpgjqj88rO
+bIkxb15Cg0M82942I/8E26YRGe+UxNEwY3cJ6yXyhflUvA3NHw1dZDqb4GUXi6E9DTZbF5wwZM/
9r/ihFl+Xk+0dq+HQC57AD1YhrRNv0W7kJTOQeYK2AUpsQpWhJO1XBC3IjpCCX5xtN2aEuH5ERC/
HMwdhetmP0tNBBh519m/Vy7J7MQ45oZLYkRPwd7yZp3jvoyOHYftX8EU+w7UubxiGW7u6Gf4U6h8
jP5ECLjn4ok+bAQEGKLieT6XSy0U4gL/Utv11bFi+c77LNMoqhwU1RhQ98AM5S90X7b3buta9Xfx
NgXwapXRP7OVc8yhK34o8p830szF+aDRvJcBGlBokRspHluG4L6kt0C0pEi6fcb72bQKRlEWej7E
NifN+rdgjNro2pNDJCAPJufAi5TaHSB99JoMRJAoeFrur8j+s/2g9BUE4jQdv02LALx0HQuVGRf/
X4xRAHizfutULInoWk6MDjEfhu0e68RsNylhyyC+MgVSKEEoKgEondCiw05azZmPvR1lnVhsT6kX
7OBuqhF51uvkcx2bC2KpvIoYF7j1e7bM74Yo4d6HlJvMRyrBbGK9PR6gevdWsHxVgEQI/ViGeCBh
TQBm46zxSn9aSZI+OyZO6yybIwgYKx5vzYMv2OHaBK8jGeYGQ2roJH9sRiWqCYeavb63EPNuo5OA
wvHWOOYBUK5GtNWbQUXZGCiF5fcw7LPtS4zLAUY9gz7mwTqsrpSpUBIo/GV/NjmpFwf23pPtGXFq
intv/Nf89npyckbEEYt+h8SO29iscnoamsUgABdQ9PR6SAcuJzbBTqIvVfD5nK6kKfoVvjO6GPo6
b3C4wx+X/m2d/xBWu2oSsn0S7wHa+M9zUb3jaTs7B252RHGvLKPGR//hJe5G+lmOdXDnZDGyaTB9
uBqkdJ+cIQ095DYhBoa7n8iRllVXtFfD5Oc8wepopZBgOp1XdSnEGhrXT8Rc35kNj7lxTW//6tdW
HeC16D0H7gOrvSHN5HhGMpOkeJmaBRRV8gtHXXFjgCtH5Mvo8HOFeDSPJJzUM4C31ESt68aRsjgX
aP1VRPkHmF/ujGO5kZ+Yh5LeODCcq7uWwdJwylReDNZbpTJyTZfwRNUyX0CAhTcUwGZ/d/YghhhQ
kQGAHLN1UgBNq0KmFgqsu/UpdY2cPBYeoJjtOu+tvMJURsuhFVIxMDJtq+pMm4yGJCdKlyn6UGaQ
P7s1GUzPD4KUKuMGoGV0yW9iCCmcbvAH9M77nZhdoSfGm3dyl6Sj36debbkrGOfppftYkZRz8Iv6
YFqOy2gLtJMi4qFLCUnP3bEamIDHaBeDZzA5/MsPKYsDZfIC2Q0jT1Qxr0vVSiLC8rel2BcGsAuk
VT1iG1egrz7h54HgVtwmjpY6KDZGC2laoBZETKrn/vyT3dapzUBuZsliuc1maVZdJNmcLCN+5sSo
A5RVYwaJQdAkxgvZn6e+h2VzC8/7uSSs7gAIlRHqPL6Ujo9jjBUKNwvG9jmehJs3Pcdw1uo+57hS
aEfp1xkQETKw7zMiIn4/HWOVvTzfh5wGYtITVictmPqzOly3olSZ3frqvhkson+AMyj4H/+dgZF3
sL9qMownZ+xvlxaQKSKSTU8MnJuV61rQ1YKeCljlpPIygJw5i3W/E3AG1BMrp7k+WU38QUQF9v62
iZLyhefrAytbZgA11TQjKYrkX6deaDPWsrBU49Uk8HMAVZtZLvcFD2/FiX3Df/7e0PeIaTv3KST1
Q5a9SE9/rqFLkwj7D7yIAmOvjaPc+yQWZBUxuFGvUqYaHtoH3LtvOqCR9eDloho8sA+suR6Ernbm
hyM/ux/jgfI2sl+UAdvRdkWz5iaXRdMzKw6TUo4GJ87gQ7HY51GqR1n0xGJlqH1yERZF5fPv5RDN
le7ObqVYFALyNdq/IlxmjAKMApj4q3vq8tPNOdESq2f8o+sxli9jp6tHv4jDK+eu9b6kKIrU0S1s
yhtFYd6OiJYeA72Pmkx3YlZ40R3gWP5z5Uj7dmsyEajKecp2D53JQsfzCuxTjOpifDsZFkIBMqG1
pshukob3m2eOFyZRQEMF4zhOiHOPX6oh9HM3R1pALTNOxyhnKLqxgPCbAo77fD5nUOue06JettNN
q7ogv6TSlthA/KaSb4fn0XtZ/DRGlaEMTL2fRZGFtAQgwDIyx4Tt8FIAxhY5XKAkcSOk/PqlF2MD
F4YXLfVbt+0NfTOY5vhviHNmIWpxmin6xq8z7y6b6nvETqyT/coH2AiprvrngljLixoah82ihN4E
dJY9vDmTffJqDdpr3+J2y96MgbC3RJpJePmO3il+rDfk3ChyddiANen49tbVd3AfW/GMywq7kPL9
pgbittKoKZbeT8sYEe+WJ1Oo+hQGybNIsUcCMgcUtj6atdFnKwkX2Do6n8kh5O22R9RRZPV3IvGE
cLedicDkerLfYy93m/G+B93pODw6ktL0RVZziXbr12Te0pz4xPbfwG8Jp3rHRUeo3m0K+y1zRl8i
klUJdraO+cjGE3yhqw0NATmT1x4y5q8KGM03lUnFiEO08EoK4fPTAYpycw+WojZNNtbTYROTGvh0
CedN4q9+JgJ7Q/+elzwrs5488QPyGSl9H0n+Z/whqdYecp8l6AtRQW+yVS+qS3XMuz0WtWIn6ihO
XHlDgwifiG+b7d4ETR2XEKDxNJpG2GZz1L39VkfOBoGtNiwtEJGt7bwzjzKHf8DNU5WjZHqeYtos
UMslYPMeRPLEMyQMzGqBV9BPzUJdgDhOjMmt5aj189md3ttvG32wOZYA4pCh4snrwG9OiRsUTHj1
K/thKnMFyX3aPt3Wccnb7iU1TgqN1KkQXr5ij8NwA5OdxilaarIbtvdb/moGSQU4PFGK9DKDTKLs
tJH+F2z81w4+Q+zo1HhR9sOFYvxM4rOqOub2RKJU0fBNhYh6EZJ4Bb1oFcsOlXPgvxvNC/iceOMg
tLHbvCEJ4/aox8zkg/eqyfGC6wAIFkUsUNvJZSug/0HB3wHRZAFAlPxuoMIKhjpn6VOSYGuNwLts
6xbwlwxkcV2k5Ls+AwwX8oBa7r6a/H/WrH19oCVDrIr3qUmYTf+YwthbCmEKxaVHE/AtaQ4B7EBX
LGmGE5LOHr4kYqzFJvRmT3ZryK6LkuYDdEX3SUklkVcfXDtp3u1zBWL1IblZieNhqvvPyzyz9iFU
G+hjjsB8/hrpOQLLlq9L2E0A7F8vqnwWrJmD7dPXKJkK5FRBj6zNAE54qTJPPbpPPAIr9GLagAXt
75D4nOga+aZ/MCzGT574xhxljA9/n3oCKQd91BkggUFA7zBbEqviWfHcaPtyvQf9dJuCvhOxmJOM
XWXQvmfw3hR0Gfma23tqVJNl4xOFsWI2V9Szzl3sY2QA2XAHmfmPuJ5zW/Gm4CHJbQHMRMMLPUBm
SMyI+SxNlyVKpPGc96rsdsmlelGMr+mlt5SGOM0x7jT00knuVfushFbQUZaKcUU4Nv14QW7thgvq
xkhF1KCjvHSI7sZ8zaZyFSrojNy9szMkRSRjfbv4SBvGsdXhH/6U/hEhfo7EaXfPcxrzRXKofJLU
qMMAbe4J6Gi9fKW8p6NQcfteVcUE6rmaK3wNXQbMYIwqRlP7u24BE2YQdAzDmoD0f7bVKZlQ/uNj
PBEFMM/AqOa/sT6YZ4v1VDVphu5Vqs5gFGTAU2s+7SJ46BaGg58g1uXwNY80hnPkk84Fj6NR0O7g
zFNQAV5ZgBPfx/uyUv/7W1A9ihUd6Bc85TmOBxo2CHKLdVk0+z7pLZbQvLf9eLcTAFmEZB1PDgFJ
FTdtLOFQPcM6Z8CTCErjp71rprbtPyowamYdO+6vZzswxuPwrc8QjxRHSGoY4qcDgFaDvVtHs9hb
XRU3GcueDFNuod/0IjjiuPh5xJ9Gd5KDlMq9duFyCim+82XETRFRztIYqPUzcgeDDwf4Kufc84BE
yCaW4QGBAQayq/B1Ev2lr9uTaGM8gmeYt7w4YZcpDRAnzWRmRFeE54L0e2M4xuY/K4L2XE0O/VBr
h6BMJtU2ERsYVpQ3BJpZjeaDnIuH9SH0YDEyqm1vQ8C1Qeb98LREXDBfkPcXYCH3uZnQfsastbgs
bpvx0Gx1An99IUoC0m+iC6hulMQTn9F1Jrkbs3Uq4/HZsZcCoFjfHvQpnWpHsSEsGEUDKv4TK1y3
Ln/RMjvdFoB1V2v4sRuPiPUl+3yqt5MCg3F3xfWSP1cOCNl/6w1UwraCv6O2s0+iBJSj1B+qPo0g
L8BrekjJ5DKKX0aYfs+rkeoCLk45ON+DGxPhrCYdKBqGB7V86nB/AKbOgxf34MaApX2SnZk5t1AQ
6oG9P6fYeqH2mtnQwNrvcTcJ3t6EmK4118ufdJD9xi810wOzli9XUnl8yOsXERTdT4d9SNCohVdJ
Q5N8E+JX9LInBMzMj9tqWgKa+XLEkQu2QBVusV3SclEaKGf8dZBMeOCOmmMkbaSJiksJTvygdHBG
cKaNjLOm71e53zcLfcNv+wWZxQZ1Z8eYP/KfD9Q1GRgZJU8WI8L4TS67oee/QOztshbFhEBeOdmt
lVKR5OtvOWck15MJOs7qHkW7MtxbGq0u1Lv8TXcroJtstxM9E59bSpkMh0CnM/OU474C0uNLIbQ5
jDqytCGzjk4/O4Yh1fOvC2JMUwWo+/6C9XYcXcbe4Pu+kjycl+1Tp+k7wIpp1q0+wPwGbczktNtE
0aj/qnkc54ca2d6urPA9gO0xv3yoetlBnPAYf0ssS/NYGnTN+5gNcJAEN80BR/TYQ34C9IPSo5Bi
90jS4AEuTm0Wp0ldAw4f1HzDFGg8m0GBnirWgC6bI9FfhxJSTD+5NRyYIfgZYt6quofQnHa/uFNR
y+NJzOSbf+f0rBUtrK56/93r0f7Rfn8GRYJpzygb4nxyGGi+evNhqxkNwB0IJeTe7ABKestGh9wX
oRT2LWDat7U5efhg+UMVpjd2SxqVVNNs4Mohou9oa9BCokBzQGPbh/+jMwwNkllEf0uw2o9qEuyV
xD6JkJa57h9Tq4bQ+vu68H7e4E0tfdLk7XqQNcMRQrw1PpOGZDLAg12bqVpNrOerjtwGKR7nRlFE
x0C34435tuBLZuY3sMnwECBLllcCTZqAY8Vca/2k2nOHw8HgZnaOdn4ilZj2BiRzM7dZJOuEfuNh
uetI90q5cSScgr02oaaFHVeqMLMU+esoa3NEe1IQ6VWTss+Ia8clLHpDh8IcLEGLY0iMhCwuLAl5
911KFPqeexj4wC03Zk86ybTDu07Efj7WWTU0onMaV/YCzexID8ImHN9xKK9KPpw/C6i3q7/afwKm
d6bGUcTAAz/iLRwMpEEQfWz1EKgbQX0ngSIpllChqqyAdoz1Rm4o+eIjsytMkuTNE1BIkFQb+8DE
mLJGBZrYDjS+oaHLCbxCC19gQpQbLH+1xbeCv2gYEJDZz08MRygZ14g3/Ba+rZf+3IntmjYDdvUA
fWCPDKJXoHH9XfgOPy51FYWWeeRnGpr81vhYd1uoQQPc6QBRP5zP9OD8JQein++fXA6CEDb8yfKF
krgTrXIfr2yO+wQoQO93O6kdcKk3zDcbkkbZgjT91dkL6iLRNBHCXcY+MY1fu7Ct8ZqIycbbsnNN
nHXJFZ5ZkHrY6bv8BZ2etisIM8nbij3aS+CDb/ixqjgRiygARo+XUirSiXYbqqN1A/D4xCHn/InA
WVY+yd+FCNhxJOjoeBOL3AWvcO5RpM+bRjrWFL/k2UdQ5YWtDvJ2eIKNCYSdeLkKdjzQH41FQrnA
wt9z/CpCwgr4yQ6JkkbrdDXUvS8i49IT0XKzQgX7GZonWbxT1qGcleQuoGbt2XoR+fXSsJoNjESt
fr34vpdbf5haPA8/JVhUEu1Go98FC03ZD+jShgVk5v35ZpUAs7qRT4Kb27XKJu8IqSlmYd5/OrZ3
d1Gimr0dkXpWgwxu0n1FJvcP6xPXCC1HLzgUkHWvJKFppXcnTuBq+N+FbH6BP/6cTuPkSzaBlZ5n
GmsSaG66nfUzZNIeuMwWTJqEoBYJVSzWSsayR6KZP3tymyxyNU56/hvzGwKq4/N7OSdG4ziuJ68+
Lps7tLlV4nfnBtQf1WrNKFblpGil5UCxVSE+dFEtQ54hlGpGCo0WeJui144XKsj1tuiAEAJdOJh6
7nZ4DgcaO2pvBIRghuZfIFEJeHl6eC4GCPvCD/TyYTZZ0PwpjKORElvrtWowileOkmFUMsRIefkp
glumWlbO2AH6yOdW6S+C4vlgVmNe7mhStyiexFlPrBmu5YhJ/n9JhmSa1O/ZtzaatAQ/bNLw9dkW
gFCavf+TVUzoj5r4kXjeDFAC/lqSoIQTNv9/mClFXc8irthG0Kox+cVGa7rXtvfMz7Ufl1W1x3LS
eiS/vtXT0gbZVVAVHIBYXCh35Hw9kiJC+hrkMpmxWguvvwiVi+oB/7ZvycpsRD8yo0rbhke2CEqp
D8K/BsqpiI57sfWC0eJNI35L+hY5AOHqQyBQn0Pvr/IRSQ7YLhUxVg3twykJwA3YY9c9AD23sKgr
tAx9lDxm3SUGxpYcEUTjzqAMrHCY4tTAkB3PKf0w1P0JyxYiOJo/zkXKIiR0tH/3Rzigd2UyGvHf
CWngyw75iHu+HCOQIesSEhkoX62o7S+pU0GcKPG/1HgijSyKlnnLKJVJdMf5wtLRLcC5RuhcW+uy
WdSQgZanS4Z3i1Xui45ioi2kyyP8yCO0O+dVktVY/3EoWcJ4cXfyrkK4awQTQzO1N7fvcaA5Iu4p
D15qR9UUZzSar6W8clTMV89GeeJjWy3xrYvw+Mt5wqO9zfzeiU6YSR+Dqe3VxikY4mhj5ovr0sEa
zeVpB/C7/Vy9oyWBCK9eZmsUt3o3kp/phUc+2pvehDT2pmj3/JjDubj3+EDuwtewFHnfaGvb6oPa
6dMJoJUo17q0JXtC0sjt59ajFLbRd1H5u9s96ZEJtRPX+ko7gty83P05xnBgmqXru+wigbH5j+2s
vQbYQxxoqCVn8tLywwd4K6VI38yMMS+r8F2hhopIeyq/ZA25lH2EFtOqg+3LZxlZGv2Xh4DhjpOt
VcOm51bU1wO1rGa8BSoeCQT0GGtyoVl5Dh3rCo1gelQxoVW5YVuo++zZ5vY3Tz+JhgHlega05ALE
9KCIcBTiho2Hzw1TQzroKaE0GJxSyMgHUDTzQjjpMm01OjyoIEjgt1sO3l2/NHsFbTcGrpypzBdy
23B2s5psVg7bgmHbmgL3QGV9dCT3LkmPWtmI+GmkTlDLSk0CzT0mO8wDQx1mj5bYI2t4LfJuAyYw
lc9u9qUf4nGj4U1iwinMZ48KRlneWX7nAx9NCekmvFCgZ/iuKV0oZCHnbNiTF+GDzK0DXHX4CrS4
7hNkOO+yvwF062pnhhmSOqnmKFBkcToMPqm3X6CmkTHRoUfUiFZEbXggWHWNb7YsDPKBvEOriOnr
7mnlO7ReMx4OgvkI8xmGTaB0yzkoQxDH1Ahch4Dah/+Jyy+ZkqSNojIsH1F+bHEM+qS6J4iCSUn7
l7Pr/xkA5q/0X/h1RdkI3YCGsQEY+mGM8igYcFGwcoF1Le1gyhKPrqeKLMv/hsRNpZwQ5HVOg2/s
aBruoquNkQ93z7Twaogk7yJmuw1v7NezZ11D4Cwj4dWkVboNBMG4WWz/cKPkCRZ6SmfFMLoUr3DP
4J/uRb82d59MfAoBTPS7/0cWGB/hHZn1igVgAO6Wgn79polXKBnVnet5qefhbkOkvoViwgp7cfAb
bsQoOhslPUzDHFT/8fM/AhYXDVgQnKVW3qRcVGFrcf/XrQtHO++nIfCuzl4Kh8i1xO7bp8bGUMuN
85n3yfeO+MZzUkAAdY+d2pRaZyUvsJr2vMhcDasZA+xhV1hEB17/jrx8BUMW9tfRuIpMX0XgKpQ1
DhADi4hWNL9MLQJsczZx1X2UOXFDg6Ph7nTO3ePYnLZmftnU9Pm1vmki5hzgwRKFv8Dk3TxH54hF
GWPvbIHT/6xNKXV14KHRYeHYUxDN2miiAIwqUn3Dy49+5Q6/yu51OjRWyTT8CczWrVu/GGjuEHkT
W8pFxIGpIgZZXBFoj9Lim8+um3c3Fi1MnybPwp3aKLUvumaccJ+rXe8hQ6JvTl8UhSQDtVawI+la
CWhfXBcuM5SePr94iK8pL0b4thEYzklFmXaZZt2tRnHlIb4/2nGh01H3DFeF3o/wzpTdX0MQ6J9p
5C4dxzKA1hcxMB/6x6XfZOtDNixJ2lcj0WRWW13osTIWuhvxuuia9HwD/VehQZ5Kdq0MUrs7zA5l
hERY8Da/yq85sMQ02wQbAb8iVnoBSyJnahBa9VkJN8Mh3UFzYGPSS70wqf25XMeWQKm7OgQ3hvws
vRHe4kd24DZ8y1HYkbXnUgabSW0KTyvMu3RCaHWb346tsrOhNUOSYrwbfvAYs4246Gd6BP7JYyfw
dPa26ynO92TZqXCu1NBmpKe8ZF9eMKigG+AUnKYHYVoTCnN8TXaPDYP14zXrUayTdhXww2GnT1Qp
3L3+M5tlLGFmp2rGk/lmnkQZt8ny4nPvzhes4k7ww9xXFPaA0QKyNtRcmC9DLUIgHOuUV9bo6SlL
QfQ/+Ce89GgI+5G3VdnKexSbbLN9/+nDUeNdARl9Osnov7nE+sZfAF6k7Z16/cFcWYgWA8xvYOnu
/JZNz3tw9wVXV3l5j6/6y8bsUq/VDVTWHCAEvLU15xxGkkagDXa9FV8umWGAp8jqKi6pQUJz4WtD
nWSSpoia+x8Vx4CAR0gw9+o1QpVxZ/A0CP/igT4tQHd7DMHDNBLSbWBywBHQtgBXlbVmpJk287gW
E3tN5xlS9tM4heQ03G++swvXv15Rr/LhNVjyhyrf27/qnHtKv+YGLdJvffpTkPDTiEa/sC6tqpmY
Jx8tYEkAwZFzBvDPwmOBykaHEaLPkAKGRgD2CT6/3H+XBcmkKQ83WkJ3XOrEtDi0m9QHzWvGrSiR
h+tisY0fKpQjKZkbe4FwS+hSmo0RVDirN214t31vLYvwNciyD1HNw2W1QR5sJsdLeEQh9osFP4n7
Rl7Z63aJbfnM6BPzWR73InW1ksqZHyyQFGVSO2Zu8HTWtwLLAtUpXIhYKLlB5ySnIBa3vwzqC42t
myZFOTuH2xcrwaxNSsMEwPE5rSyT83BKQyzs7bBWQ3StldUU6kcse4UTsPr2QzKKf5zq7qquaove
HBLJoA8xej1WCJv3db6inSji7XVfHi++1undn58VIFEQxnfJ7B5tGmDGe0T0xpjBk+5N6MQ3l8wz
y8zB4AkXEWOGzxsrnSg0IFP2TOXXKQa0rwqMzzCqUUEsC42+hSwVbo/e+045sQDYJVx/v0VuWDYu
XhzxyBdWutKg5lFxe5G8VePlblCSlnZSvGU7o9FNm9R11h66u+0qTwVt7q+y//Ie3iAxqZEUk5nM
zOhaMpimLlJevkX/U7TsaopKWa7/ARK+8QxNOVxjHkrkj0cOY9Hx0KM1UF64gZK8WivROIo/ByJm
lwyhTcdgZsbd1L92ck0LQ+iyMtRA+L6hMNyX9BA5YhjcmIXHnjfQgyUGgyRtIMq+e40Yn9JEptNG
MGHR/2NUzinOxXZMYephOalEnrcTt7YmW7KyNDCjOdYkmOvuwAX6lwO3HP3jPmNB394evleiv3U/
52l4XoplA5RcPZbxQubA7alirR8XXgAlQ8NYqUrjWGdyDvVVeMpuSO8buXsVLj3Pe7I0HVwRa/rh
7/kJqcMyf8uTMdgSC6A55CRfffVpEsC79gI4Ti9GgnSZ8jko7JajED/U7+4PCddMxx4NHDiFI5h0
V008t5IK1azmdv1340ukVi+kqkE9Nb2DSc+/umDYhsLz+CuIkGDTc2OFlt6iE9LuOLDoQ2jR0wSX
24HVZV4b4O642IQjq03YkP0JwiKvDn0sR1cBpwC7KTEen0f6x+YM/d6UFqjsAobnVFlxwtUrVeEY
dPxdfijm8t0i19VlQOlcGFRMPXtIYOvQfeEsNErWUHNV238zsvgmmy8Tj+3zYnVKBZQJvANMBCNu
AOkCMc65SzOIQG/K8dtISKvl9iE0UW0W9RE0Yu+Pxt7WxH6+zq/4g3qq2ShHaVwHuxvdw3xOH0yz
y+/dBfBkPSmX8Tx8oDSvzaQSbh+IIOFD1/Yi2KbFWR5Jf3F5qwWfKsK3eBbxkMu9pBxxuO8mRVA1
xVr1oWfoCiz2HOyH6moISGze16WfEUmWSb2fPozYnY6/GdNlk0m+yShXqiDy3/i2VrtCrPn7ip7M
RndAopmAnjAIAoWzocjmDvmxuTw5PiWz+SCx0xetR0zgofghGPem6BEnGiR9NGVB2DeZTR6DkGBb
NuUPliJVt0HqO1GQKZBtN7/xJQFnBU3VEJCGzJXNajWHS/iEdM370PnWsHrCHj92nlfahPDr2Z8k
IRj/DVnXJExL9YtvGTa4jPTVNw9JFhxxggWb43yE+9pBS1w4qUWeG2ZZ+9kagOsl1/yVJGSmjxun
mi4A/CHMW0mtcRaUZNiLmVDYuvIaxFVUBWMLbUYoeU9HGlk9kKu//+pJDzxF3efLDkzQtbSFGMLz
BsIbUIUiFiZkkR59awQGmToJUXRjsQiqQG+g89R/M8kFHQNw7huz8aoW4CltPJ54FTPdaTV5s/Y0
n2kTAPPlpn9x2xtaPceojRcVwZBU1LWNLOVovwoX3Jf9qyo3A7b92m76XsxnPjqpl3XwpMV7rJHC
EyBrzOVIhR+4OgBQFwDbIX+BV8yuu6qwKwUCfhLxevH02kZAsObsqDxTHQIG/RzzOBjrKpbj3WtG
1zL9rK8wRgc6eRppCgdDQu6+ZKctnJvwraFFSqNaKPdPnG2+WWWvkR2TSxNbDalpI21FqI2iIlQQ
WR5w5x5PPKduosEfDzi7yZRVAjJVHyhfJEjmmyUdcZwZnxwyqpHDGU2cEzOVzvDypZ9/x8TvF9Sn
PIuIDRqNlUWzIu9Mf31ZdnOfjRKxuEEzc+gKlLLoslLarbwCfXqtc21jngz34bauXqi94wLCmsAb
Ojh7TC/khKoc70WIp0LUtFZfcdDBNxcJUmLM4/AzQMQ0zyWKjHKXycbYjh/x0HATHaqq/2WvrB3O
9Sb+iVoPhLK9BvGTITw4BIlsQSJThaqmZoz2fKEvLmJ0cFc+Xq/NYjjHNWzNV7CFosDjFvP8DNc4
YpKaYW82oAFjZaMQjAGtr4T3N7ToKLqKFfO30LdOKnb9IpBXc0KHD8mZLtBO3x3X0wiUNQEU0tWC
DZSkkEDsemSDsVD4LnbqXI4WCwGdOIU1EFm/hvOLzDp8pq1ybyl/RijGjvx8H1uY0qeVnSkGOu3G
ZokJZkHKRCcVgx9Pwbr1h1hmKob5Ro7ArqHf2BVE7gRrG6HrBI23b641IiinE/bGcg+ShHAGpTWV
aoR4vp4k6p5/rKozRjoAqSHQ4HyWzP4wtdVKpCORdTM0Z0nErnO3RYhrad5ORVoZs6zmwky7ximK
NXPrb5V07LGTA5ml4P7ElTf9Iu1DyumBEsd+QySU7lYqYbplmm9+Ms52nfdhH+Nx7p1ohVU4WhxF
q61HtTS4+NSYl5sRnPpRuCP8+b5fHXxAzpPxA0TrXskxSiTIZG7rai69kwD4+J1RnNFNlGZR5RUy
iAylYdYptT1sGjp7bcCjZA+2DcStylnrMC4KTQXbjmKLJ8L5rRYeRJs2eVa7eCogApoL7oL1meHd
eBk6haDURrwBen+OiS07UwJPm1D8KdUUgBHXloRufADTgD+U4la5wJoSTsll1rfi2T9kOlCWvIU4
0Vu53CzPBNXcjnjyC5/b+EAvkrFTcrui8C/6oP/WGsvJ33VdOchfixNN9MJNN2ZW4AjhXPObEc5d
2iUnyApWpdMeAh+zJs/988LRc6oj9y9jMBLlEl3D7Xu1TLHcS2vp2ZMQcZys7Xaa3fS5bKWtsFT9
yF3wpncwVuote3BLx0oFIZWTpxwnqjW0qqEYTg2QsI9e/EQ6PS0E/mEyVoh7Z1G1WkX3L092JJfK
LN6rASz7P7p6vrNsunxivKweGydLHxxhsFzEZFO4IBv5tAB36/wTBxsU4BYTDw1FjrnOER7j5h1c
Xd7qbvDfEd2qJzIgTdT05lL0oyCjVwybAvZgUVo/6my4qlkQ+cn+MRY+BVoCTYe1txUY2QW6PiFC
0Rs7hO2ByYjcBOKyJrQhIMFEnqSONecI2RG/Wg/JMhneSPNY+mZFNmc+7NWdyZiYB/AbD38ctVfg
OBxQYbG0698Wfk22cCHJ/AKRICyYSxWiYvsC8IuUQ16lFcqWDwSjrenE4ngQSSGPE9dk21R3j6DD
4P8aAc3c2uEjTlX8T/9naXIXXE7xYo/WV72tKSkEv5omxilz4bXi5Cr9bp2AmX3lFviD19fKCXUm
pDgBZZBmu1GOwp9HvEI8udDK+Zmvbr2hHWxyU9Ax1b/l7ocSOAITM+TSjPAzPz14Aeev+F60xSFI
LFkGORuSMmHfdo3wqnz7511nyuKYZKcONmriUtg5kdM27pI07m3Uj5Letvf3U9+2PaKc982SYGzm
xfRpQ/4LXIqYSzaEPlWemQCTa+1ku5bH1GpQgFI2bcF68i8nk3JpTEyyraSJZPcT/EhMY9odscpz
gK3ZXST3sDpUpDI8OAg5HYTA2a7pQCCWFvi5Mt3RDdzDZ4yKJXZDXe45lmZqpvrprM6f6lJN371g
3xuNBYxMllQ6jvydDQxYYkAmGveNdxUF3yHnZ3LY0+G0YJC4svm2O5F7wybJYFvQBwznXE/0Cop/
YiDauoeo9jFibY6GIqDCIvfKE4c4wvCMjfUBeqMfTvHR3q7EUw8Rwq1QMAQc4lY+8xbWzTQB9o8+
r+dI6GBGxd8s9W269zy+B6P54sansvt1KnK1gKubfF7rAp9vcSFwOyhCKALY841cCkBclTGtRq6/
xYKFkVO6p3fr6yOx1/yM8sYxXB5IcGHaFr4mZNBQzeWlcZsRbuc3nN+M3FK3MXcXvYOlAOltmva+
ABpAH8764WBUHR9yk51vWrmXOWhuCJzWxjRKXrATq4AY6bnyyxQC9VkGV2wcs5PKCSh42Iy6LHfY
p2+0lYKEhoQIOtjEVXDTCXIkoDJC89v6uYRqQLyre6dv4RBEaYXS02xS4l6pecMgI8KvQFNyVMOr
yf7WWLS2aQ7G+Tr9Qnl/sUwkjLQgTlaAheyYpL9GbIgzGdfIo8S1N+5b+W4TX/2O+0Ix0ud7VQYi
GSBLALxf075pERlhPiTEqChbdReN+bWwDxYHFD/Mjku9+Pco6D7IgVs2C/tg63kdgS3F7KufiW8m
BQSS2YIB3QR3KhB2wl/NfOwA5BmqoFhL5TZ8oVCYcSy4LyVg8u/E3Odzx6oJNqqjA3kTpPK7iBF9
6A2M+WHXwVYDIA0NQUFW1q9obAAJWsYagY+zV0q7h0LgLp5JusJWMJj6Hv2z4EnZMte/UmkusQPT
QG9U0w43nth6pdUk0ftizWyImh5FLLkgLvfqIdWVredYEURY4NdR0frGE1USEvLXXOXeGaBzhVoX
dkAIDStOUwWyQZVffiya2lFGQmN8dNeR92ftNoWYvG4yfJGAk+JOBi4MQ1pLgv60i2SaNxDmd4XY
9aChPNLg9KGx+4w5gcmftS0vnNyO8H17knmc/iocOsrtyYvW/bTRZe5qVRCWqnbJo3v6fT9c0Eot
Xy2V1Hp+mERlC0hKMn7ajpQWM5EfQg66XxIOOSXYUWyUyV7aQQXPUyeAWUdxmKQc1hTBBBhfH+x0
B+UQkrHbq+na2vM2bkGk07CnXXZTm1Z/dP7IuN5K9usC2YyAAsnGPlWJPlWvsFR2kxbWTUF8xwT8
7i4tjWv2JWo0Qw0ZsY1dKcMDvDkFlIwOPilzrNgG7T+1mdLFvB3jBp9t/8X/J7CbPbRXgvzE7hCf
E+u+wOdLhLJHwMpFKeRNPzfFykfN+fe00fhmU6nWKg5nxjlGHD7ZN9UWdfMckR5gtPLeemqPNEGp
b3HBaGJ2uS/+vaYNiaYfVpGkEdg5G2Pw2nQ/Ly8P1azmIlXgxPbzFZsuYissjAO5C6XFOBH9zbTM
bSISXm/2ni7OALE/8pIe12wOuj0gdPgCf7uQN+lB89H7/rsKVkMkQ1NdizJfjs0gDHXLqoGXEqnY
Zlmk/s0OkIqqKSDb6xvKLCJC0Lw4X5c/ZM254wOFuW7b7cS4rdCm/COb/i8sK6GkDNVBAxHKcIsX
ZnC20iIpyWCXD5uLpIrjqWJGqTjLYY/5hm2BPrhAmToQ4ifM7wO5s+aLj6mk26zKyg/s6SEFK9Wi
4T4PtL3fcK97EiMVQKL7f8bzxmpbj1/9wg9BamWhV26+4oe12p+B+s3HDQk6bRPos87xxzeO43MG
CT3BTfzpgem8mubqzBGQuTrzqH6T7Y+pnuskAi4ypg1Olp+DJkIdS6rzPprYFFS6FSkcVU1Aujg3
OBoUVBbGiCfoyQQwBpntq5aBgPJ7VBqdmwmhzh4qO7g2yWU/2vl+CNn3VkvytNR9J67H9/w4/chf
vDRIjf/odIeDzX67xyzn3luqov+KYwJm1qjnrhP32tAOjm2m9sSbwSoT0NUTAABPOvvWoBQdQBCK
mbMlVA4JiZdAp0q07gh1oVRWYcVnf97P+NGD6lig8tDlzxYDloxC+jM+HAU1Ovd/R8TViwVDijNL
SUYXlu2agTtVNplffRksuYnWVSHkVHw2xtQlLCa/tOvXNexB9M5TPRg6Ai9bcp6PoMor3dMCV1Mj
XuvzvhM1M1NbDXcTD23t5TDGHJqa4srNgI2N4Oop8UmTLsGN99S/K2Q2Sy4OSzY7SnqYQtl6vwJH
EGcGELKefL50PSAxMaGeeIKRVDXoA0ZQxrCJ3Ah0jfreSktVo916dPOj2hYEAZTkj/tDqGu/+eXS
r7oNkdiH+KyeSVxkadyedxqx3vTCmFCh5j0YrgrWg/gD/4m2HEGecei0wZEh1ocdvoPwm0bzkTxX
S5PnxRcaoK+xGXPK0biZ4P1Gj8zquTwHZyXvxYxQlbUD4THriq6fYfqh2xoJ4SfPf1HAcyTwKKeD
ir5sqfUNkAW9JRVbozTzRO5uK3yVvaA9bG1K2IRFuLNeI4vpHrKTtKX6TIW4+qpAZKqoJkz9T/EN
DEvavwAZk6scRKcv5kH1UAep2YdaAvZGxEmOA0YYX0W3CjNPHyjMrmbQSZhIrGG9aj4Nj1CoeO7H
SRahHqfmfkgw3rPXaVCCUolBhyTROlXvsHeuEle/dBk/Bxaz+8IBXXOd3zC7lkLpK4AFyJ0X5X57
NwzOGbX+Mp+P4GwW4VTgbhdOlDbE19bj4unyMMHOUWr1d7RRddfQzFwS0u6hIZUJ0t0zQP6okvfk
eTo8r7da6hktDodWJc2wJqkoSPnuisTUcXEjX6hQtah9oZIZ8qxOR5X7wlHNTrUg/hSlHKIupPIT
3TLddszxEBwLD/qu7r4cmcCVHstayivll3OAwfoWfKiw194B7EvJ1Gy3DM9ox0lPvLRhr5pegv2X
Ofu9AVqwiWNcKozmchujV1NOVl0jlBAO2V63fj+yf2HIcop3QTWWF2EESNwlsVPgvgvoSxukUXOk
Qm61ipJ7TefhrXyEhXVZaisuei3mprfSjBomVl7oy/Il4Y9BaJ0aoQfcFhtCr5N9dTePkJWXhICS
5rKg+SUYO4xVCAuQ2m5oMT8a6Ir65CpeZmQfTvwX4Zw8pnUo3YULngGXMiaeYz2woN9rcCQ6RUIv
I95UBUhzMbrWeQnP4qGhkGm1U2nKJ40FvjfFpLQBamygRN8BChAPBBZb/QYuH/CwuSXFPXMJCka8
OXh7m0Sjf/WkZKSdbDuiPL2FVmERgBX4Ohz/b7ZNp+x2lwBYX9U0H8K+5EVKepKRH6AGmn0mmMaY
IK4SvMGI5Jfz+/hpoGKTv5T8IpXUerSH91v5vv2BDsFm85ns9VPdxk4aimsH8/+73u0qdPiLFR3e
JMvul3hOKPaJ1Sur7cK/ZYEC4g84RYVXIRot/91ftxioOxMEnKt8XZnY/9PGiy/kz43c638QwUy9
r6krTkNnZ3nQ3Dw394u0FFM1tk4kvrI+mQJoMHAa8D5J7sSkfH2YsKhWbtpx+sCmOY9nbRylvyE6
ZFE/MrySZcjklUKxviIezcDWWBROLXU5vs7I8iVHl0MKq3uq1eePDgtJ1xgI+hZGWpJ5bh9NZx5K
SC+WvjMgISVuqbVPLX8uUC6nYw0b1MeMfLxyybesqSN6+AiEM97gm8d7+Vxs/rFRCIa2wfvValfD
cslL+65wLBADNyEzHj8fYlEYB2+7CJxjYvx5perIrmBAAkxuAyLejytxE0gwwDxoe/q2GD+wUSBp
CBYXSWEnRgfQpkVYgMk8GFBKjcjgwj7SIcnZjUMlyNyoR0ZyRDwTAH67WiYZv3c9OQYsJRcCGEgJ
pq13VU81jXaLJUcTp1bgpQ+m5Kh16m4Za7jjGYPsLmKL4A4dFo4uD4wyPRLZlFt1CgKEz4hf5N9e
Rq77jSyBwzj2oDuUn00cPXsTKPXugl1eIGuZU5UHLBxai+NbiNnMdF+9vc39ZzMknCS2Cvz3PP74
n6k/OLrWyvhofokWlmTwMsii3JzHSptm6RRqPwQxAzK9M6j2YfmvaUlNtfEH4BX3p1Xy56HgL9Es
lBqAVQdenwF0QDTnt00XDKsV0r/OkDiJ+XOx9KGQo3TYF09pe0MVsKgfnneW/opOFHMwzjkvE9v1
83U+oog8nw3vqsW9CWNvfoa58vd33aBQJK5IoCRLKTeDJmxW0k7ODPh6n8eZ1jb/YNcYW9EBOu7U
Lwj645uRQOSvaVByRDQUreXFNpIRoxv83k4iPvlCPDfO2BqDu51d5hy6h0nAnB6RdwkZZiCDxT1T
fsuD5oauuRCcjuowic2k6pQ+qiZ/Z9s+xCIwUc2aLr6bjkGsUniwfqYqOyAZdikKfL409Hi5g90p
cYwEAX9uBDpBXwPG37gDIc0lmzFct4H+rW67HwZd+U5ukni0NlqVlp47Ugc3eJysZfof/sQMtNxO
xoOHs8y6+rH+2JWIfRFPixHbjJr/wTBwKdRhpe1LgqWWUjksXyQIFSkFKJvR270Q8x6b/NHFErdJ
ltt+ZUPu2RyrvcncAQSDCLT9Nwk6VZWyeULh0gtWYnBXseHe+9NIA4554FW3N37BOvF2r9IqIviH
ra8MDjJoHICj+NNmT/EfkVa5W5M6Q1XKuD6FLJKmyPOO4Sn83lZlq4TC2lrxp4aTJ7OgX/Bgm9Jz
LOUh/NX7w6hKQ+XjP8CHCRRIFg43VX86+7lTdItI6cKQcSpSbb8ljFj7uffngXP0gbGiCp13RI02
vhdUDFKZqFXZsekYyzBpoXG4ONfX7gjSoIon/P3/j45JrT67BWEkKVxX4OlNB1Ot2g0xnosUQlbs
cIyGDyueGbtYezlRR4FCMorYr1pBDAx8WdS5ErXxsyxuEV6HUjvg9RY8H/+jnm18mHGJ7TIGVEYZ
xAJMESXkvULWEB3UT3d5BVvzAakyxeDmY3kZ6PApTLwNTYshX+rqYN8VycmicKkf4B9dBopK/FKt
mE0LezZlR+pT/MD8aDWojdUcOLONq2N+gV/E1RfCpxNzxJyrUQh4z895UarNpOLaWjtMdaOh9PXi
o790An0HpYur4MHEsFnWRPcOtnuizkitpr9KHQf4HaCgaDuScL7+OvcMmLQN2LvdGb847h9Sg47U
49mUykS0fZ2CjqZEjz6cWABkx1HAhGEh2zXnaRZ0b5Bi/PuNKFXwULF5GYifRmCCA6n6g3KVa9Br
vlbgi494m92uMsc8rtRK7lbunUoTo6aMRMfM5jIKsT2CUp/+QKQur5GuRtE1kAfzhCOPrBNCjxLu
cAMh4pmJ96Uk//iK6NLMKPztriTBrTZHTFUta0swmRg9+WJFABFEu2C0xvB0ui4YbirLgiHc/Ms7
4A94oiD84wf4KU5fJDRlrCMrz9YqqpgaIbMFJbOC+eOcoYySNKjT3LLOcL0qn1qgTr1IdeT3YpOY
iTHQuy0jIG0PJO3cM75u75b4akLVf4xsrCHbRMPlV/Zvost/NRZHSeHFOYYgOPBNqkVfwKsZ7rF2
I2QlJVkqrNHAVvtAYhQCsPHvmDoqRruKGH8p7UidmsmHPwhMGTJCnWNLSWxX1jAb3fU5+tdJw7j+
cA5eScipggVKhpu2vsRQxi/w3dPRQ0vp/bpo29ZViT/tmbhlFn33165X8ql6BPGaCLXsOVWl+PHc
JsMDw/BMJFtagyjCyA1daRGBUcpihfPM6+Gv3z8rY2b2I51MttjT0oAn5XdKaiRp+kzt6ekrshZ2
Q83vNOtg/1xGwz1xqgl2yeKisEho1fVt5F5ddjewjFMWvjurNTei+FmE8PrNoRPvLk/2Qms6jjPC
ScM4rwPP6TMMykXO99/Cl51xIjLYVDGiyytGyZcdu/E1CeTxY+aDcAR2MJgbfzOAyEtY7i3k8Mep
QeUMw6okpG8wCcYQ4rjsZuF6lBZf9VUHx22ZM3/pnmQ/ces9cyIyggoBDWweKV5OPuhKoNmjmQ9X
9JShZ9HvFEpLaFFYymozzBd35+ZN2gnpKY3WZAVbAyza03ppNn7bb9O09C5zpkiqMAGt+fTuiW74
qAAd5luwXlJauOqskpFm2zxHg2aC5tjEXw605Fnc1+4WKWZgtp/44la5JuTI0eNBRm9piW2X9wTV
q3jLjBzugCYjp44gO+NlQWnmg2rHqwWRpiz4YcOf980R9jo1lK5RFmYQ88IpE/Ri1bjaeU5JkW3D
lwk5JduZrW5NpilzdMcx1r43vgz3SZFou9bGEC8tegsxJfzoG1KOSTCmE2TbnDpanAugbu2QYAd5
11MsH3p/ksvAB6k9zsOTgvZwssldBdlm8ZIvitgwHwikmOcQgbtydHXMnGtECpzTxQ5dly7Uw/NQ
sN8CkoW97JZWlbi+rL2C49H7y0fjIJvyEw5goOgex1rjhPQ3he/2V0nzPoYvrpGy1S8hFzvwsHhK
PZW4WCKo1lF2WRMk61Lh3stM0FStA4PPrnCtnhRqJw79PJxMZIsX4+JVWuZyb36WFGiNCgiqsvwg
4G0XWLnugnY5qJbAhwpZe/GR2GZbDnU8mGeSFMuNkFmfQ9uDiGdy8NLDtKoOv/p9MD0W117VOQHw
lfj1r3WvrTaMBVDPiTBZI3fbmNOcCHj0RRrocwAIabEH4oM+upOSGGbsZKJpOENxrE+RT2drXPjV
pPc0zYdPqm7VlDhZx1VFHko4VVqFOJCunFndb+oHOr9JzpMAaKXFMB+zZMlfnPYTOP6tS7njA8DO
fylXqpa7sRDfMvg208BE5W0fP7SeR4bzvG/tfG4UicUcr8NDmYfKFp+ejwuLSglF8S0SET0LGhi7
HaqWh8+pLBG3VMSpT6OEoV57Zkjsmmt8entkrkSjuDoxysQTiC3hp+9MvOFF3LZcQpKVLDJrE83/
r7VNoGuAXY8fRQD5R3pl0emecKlCpfgNz6pkCrtd260Q0n5Uc+ImGIS9oYmDHBXKp/02XFYEhz3X
8jFlTB1jeseY13YSGyaAY/1uRKHrQ/mLxXnDejSM0O7wkoYeW7wo8gBt/OWICae1XbRmDj2/N4yM
rKjCH3wnZH6elA2XOnGZ7Y48dKXyZUPhcsntXp1y5mQjRxnzPTxV2CJF+v9PconqJ/bQ++br384e
P7RRXehjVXDyXesWPDDTeXhLNjYtqUiMc4VHxkOkyfmGfZ+158ufAjo/Ij4L5IGs0ialfVnhhsWD
bG3+nfQ32o9t7YRarkEYXpc8uLM7kooBRqF3VzrSwxFtlZWwqAe/83hIfZaWQQXFgDeZXZlIRBlb
ahwh17wlIBww8Scfn55Ha/oiBk+9J3FE+6qthbKt2x8Yk5onMAo8P0S6rAUjxzAUICHHoKc0Ldx6
R7VVc9uWMnoo04cr1zmLSTpHwuy1oyk801bteXshtPsfaMNaf/isUCALAvyE6e3sk8HvjPzGl/6j
eleeeIvejgNRrhWOm5N8b4oa0TUnefOo5gHhHfSAfMVpUr0MGizuD9nc9spLpk1DwRCp1l0lhtgc
MLnc/JEH0cqlDmk+1y7qvvkt2kmkgI6DIrkmb5fBOc7X2W9I/eZ/oO/uiIZNDcOFqj8iv1nc6oR3
xmR34bQJNK/qnfGzbfO5jenuGHGSekcPjX/9yX2joTUia7+hcoaI9dcyaUnL6WQJPkaK3AMuporI
qFopXlAmvjLNXRdeJ+1K94+/IuAG7er6hSsgnORiX/67QXmP4FoFfT9XBtUcKNDMTUAd8i5S4Uo+
vgDgzqA0+95ZQ2moCeBmhqlEXCZmNP0trymJJgKZYPEPe7nD3Uh2rM/Xn0bucD7hsAao9GTAxqTn
0Cs3hDJ/LpJDK8fVDJWv1thP0oGNnGYg9mdEzosfJBBFFC0ebXk0t6zQV3SUTA1B6BaFYEwg55+i
b5lgAXJ/XnmPFw0OySSic+XsU8pyEH4srkFEKV1TyQs4GnjfZeTO8uj6jiBze8WPfh/N/+h173Lt
rpKcPHbhkeB7Y/HgYsjZiCpH6DGIaLILCY98A3p7bdY6f/hykY9J208nhdrmp0+9LO6CaGCw39VP
WuAQRLQPL6Rm+e/VeQerLSRFBAAONo9IhGIvd4dRfur6ClIZaGGhxb718n5xL2SQucApsOgrJfcU
OJvlT4pvS3wpoNG+kTkTYwZxNh5SVhMJL7zx3tVFhwPuc6vVd2WmPX5769uI7XAuYBHp7JATSu8/
rsKIFGI4/95HNtTxMGK/+ISMccNcVcVKX2qnkYdooCD/VlnA95CKcOYnj2EriLxwKKoRYK0muhIn
UnyXmtLaRn8NH0QM62Iyr0j89JB7U3pgNkp68T3Zus6ZJdhIXmviYQ9NBsr5x6UVIPP9RJHBsq5O
Rl+DUc3XvWWZVX4vkvpWFDrOH9aKUr4ZADJi2/cfqWpxizVWOAG3o5EcfJ7zcd89nBbDePCS/Xb3
Q698ojPZeOFQWgL4YnFcCg2WH4vJupXAMixAwH7ajV3zCwGJq4V9vvPg2VBEUxXVB/Nt14oyMROP
LhCOEsONgeniQldvcr54StNY0ic+jVeaqTZ85Md7ihY7NSlvW+KeWPqHaTz5pN0qFIqfoltGIY6C
kzLoE1Ww84m8UBtBsJkWrvpJObNXnI6qgOke8UxvVFgkUh2kAoxFowL6o8sYGUfj+9nAj31xdzU8
QsVO9iZCANOx0EbKlXH634Y3hKZuCCGygGR0FtSRPP3aDqdGzW7EfaAvgcx3K80/GwR+aJArJS75
ZlbUCQKWoAG270j7vQVDVzpS8xhTa21XHV6vI049kTVuwu2jRqJ9MZkb6YE6GkV/mTsd7PgtGEvg
U1Ru6gZ1v5AB/M3hdJOKPVjjebw++SWNyqsSd8N2VcPoe7qkTfL9nwnXasen9jI8D+5WFnHmrG1X
sleY3k7yd2KBtFGBo8Mo21URJY3SsdI9W1rExPeeZKfwSspnYKyXRGUNSKPVt6k15UZr32wfvO9B
KJxQVtbhmBH9hYabdE5vstUsjVZkBTi+ltU3ctfFBZNU2ymeq2g2jGBrJtFEra5oLqO0EIn/svuc
j6RE9iH6rBEXAfHX7XSq1cGMyi2i1RWNt7a/a/tnyaO/4ICAAcEDDGeeIbGmLk1hBpNcMMclZtM2
bbBojEFeOSRImItg4fGoxlY8JrQSWVupFUnROPO0lKlf3H0KM4EXiHPaYJXxlKr+VPyTE1An6hwA
DAClqUB73Wd8q2SAe/9HezZLRTAF8HETnQ69FxlAB7QU4UrWx3OBKsRDthrsj5Hwho901KImIilL
nz7VUtJjqqUdiHkDD+n3pu2NggYqGNUwSA5WrQ/WYc3rrFn0zn6tTknPuE83SKBKvduPT4Jyzrtj
0UI5wv65zHdRb5fTFf1wZpxQHXkgVvi7wmpWfMNbZ4ccw44AVwhNFoxbDw1KQe4BH2kcBhGdcc1d
VVBaTWX6D7COpkyMITBU/e+DfYZ1aTT0hCGA1OMXL1Imdlf3hPpWwnl47Fbhz0DbhC3cWBstOApI
e2YDBhufjFyNcwymx+kOWSlg2HbgwFWoZWpGddQ1hNCLAgagIa+pEvjLffc44UYu7Dk6y7BxV1MJ
kMmzYkd8pzxwd51/Pr5314WEBLtX1w8WMTDXQ4yCrRQo2TkFavK4Rnap5ltoUqEh2+1rsj9j3bHy
6I5EXp5qRVZV5kg1HuYdmYHXGTdg5J2Y1CiIdPKYljDoZRojvByK5vh2OqAy/z8NvrEQc/aOGRDl
LhFagtBzVGpEHA0Tjj8TuRMiWiYxm9Zdv1WSPUj9v517n4vPPL/VsPa5SBB6h3r/cUbsoBkIPvwZ
qIwarfTob7WifKH0HHYVXUS5d+mOS73r7nbn0zLYSWWJ+zCmrG+NmwhZN1iLNaAY1hGi5h++DRSt
6x7nY1ELI3YQod3i0FkX26tgmOy+KdJrmwUz88aw4pNJyI/kJaci77BrO0aaMsCEBsXcVxPaiNG6
r2pV+v0nNpwIb7OhNxy5E8PVjL7BMf0Ey6kvEsnLw4nQhxmXRcK2IINaXwKsdh37GbNMy8SFm5Bl
qXyE+9Iur8EiEWpWp4JgUIYIs2Zk0hHqIPs8KtbVXguy1zH1tLZ9OP0JUK0Gax//DGgzLq+3kAPm
RF7v4BuoM0dhgYFA9ZP9AOtiSb84FMqPfQtuTokEyaAZgfyHHH+RH09ZGXh7aFoLZk3bgSvyzzpm
2gwrt8+PBbTtJVmMQvNYcokCNZdYHt9/1nY2vSmo1rfir/OkItdxqWJjUYOf9qvhFLhf8QwyIoZK
QaPvDSfAqMkY/2w0x5xrTY50CKHGviNBcy5PFRgeD8FCWwEDQz9hWoa3wAVX2RV1x5tRPU2BmCAl
h9mnK3PQFhZPUFxwb8LmFg+cDBmITLrO5J7TeTnKrI22Ny2cbYPmkvBS4q9hiKp+cRRxj+GnFnTv
CHNClqfTzS7gXJ6mK4Sng3km12tn9ouP3hN2b07cJr1jv5S5tIN1zqohzFj55b9ZH1+IeOtVo29E
drP7rpF/DC/VoKOaTywBJpS7NaPbHjbvIt1fqUGiTD+7mErVldb0zhLVaAf6JmWXjLtkdg5zUBDQ
smoDgE0VFoqh5NR1L9byiqHoAl6kOs10b00rV4MNbvtpRQk/oc7CMLxWmoXTOt/xDGc5Cf0XIoua
jxYhj8+uydgq5RPLD2z/zxve7iw97x5ZwJYpgKNk84uHCOMs3XLMU6y8yJ9eV2uoZEJ9ERsWfyPe
YCYjvuDX6iYH1TLUgZnf4y7nD1Rti1RDll4+tRxfCLqxVRHmAAD5nD7S2qKiXz1hSPEIf/lQDJ2F
8AMtgrJl6nRv9fVkHuR6tEt4fzq77kcYbNqRy0lclX/qJS1PozukANz8MB4fFXVa4V3jn9WrMnRO
J/VKCtI9LS3A4E0WJXTGNdc3WtEsWinSMUFoQulhmA1JEWlPi4Qog2KWgqhFmn2EHbkV7WdHnhvy
klDol44egeD+LAtQIIvpkYTXsveGPr/s+QXza8TCg4rIcjoEWJvpCFRwnrEJaOk0vipWkv3QPQFX
UxBZtm4QRG0d2x2hC0XaH/oFpmDU48g7/q7XYWh/km3/VHDmSCXcbTO6Rg1LPxOonNQMbjkcQ/rc
tSV+czvNmF/jQVJg1eaq9TvpJKKyr/JJCNSUuOVmD45DVlRN4jou6gHAjXr/GgXio0611G3P8gcj
OB5dPD5W9j4ObemB0Fsf/3ihJT3oVJp+h6ZwWet/yLiH+yphIXDYCCSbCfUonH22kX8wGpXZ3Qep
+OzThG1SjpqufKEVp4dWOGU/PqnAWKDuoRvUVONWX1cqlUHKAb9jeuQ6BduA4TTPjx+nRaMZcp0u
Y1Gl3bLLp55EIviJBJEWc93slboDQ1pNDZX6HVv3Wz1qFJNoEVMiZJuxG9RyeYjMDkIXbbhzf7ee
/7xeLU4eNWwFfGzcHf6DFFwWY/jBfuuv2akJbzcpQyrDpIx6AbjlABCjiMTWIFdapNY4mOJS1U1C
GWZ5kAHXKjqhv5QAEK3CS8wYx+UdCf3YECmQ9pZrJ7MLRkMnkdrEqw1/dEmF3mm1yUp2Me/vOxW0
3s/ZuRrMw0e8o8/KBp5HGV6GOZ5Yy46TIk4WJ5edht+ePryKte4je2wSn+0nSNdBp6246CtJF2wB
4dvjicft58xJj2xGkKI1x/e0/SDpma7aaMgan/7Y2gWN/fzlUPZdf9rK4dVMg+5soxZAvM4Tcdf5
tryA5XLP/EHM3TsXgwYkVSqToVAvpH9Ks2vcJ6obJW7+73D8S5hHdCDo0mnGjPDMhlu9+DnfuICG
inzw5Jn9JeGocUn04MNzFGgaUa5H96t8YyYu/dCG2BXPglf2O+uXeyOnrpkDfSR+jbZt7Ddfq7Pg
L329qK8TB+0ppFpEvZMET36sOdnD3mo3mQuYMOLxumXUUoY6welhI6ujSdxrbCCWIIKE4cR0zfGk
MPcU26b/cNd66BA6ZgHulFXxbYEaRXawZwImy70h7N2VPyTD32Fzqa9CCkKI6o51OlFh+ccI1595
T9l48MolBaimi2pRaydg0uObrNZoDCiw/Pve1Z+lkSzg3lbGS9Ug8dv8sdtI9qm1AtQmzjIzE+mt
HpLLlrqVk5DaVRudj0LuSdH+i19R9J22A9k0VYq7fZJpfE7KCp/x2UkbPqaBlRLf+vMDMQpSzGt/
kFTR1FumWqO7tkyo8J/wlXWFkwLAi4/w+x7ka/nahm+HElvcczAc3JIICKU2fC5qgD6kYVi7stBK
OtWT59qrAo7Az9sT7L7gNQAfPSKOZ0zhBSiq/F6E1eB9ZiTd9e7uLZuLW6MbrG1j+2pgKcBGmsHO
CKDZMt8v+TFB7h6/QKjsb/laGHWJL64wyfVK4PcOA97y4DgpOz+AY44EbDumh4h7/ZhJMHPcP4cw
CtCsJlr3mBXmYa8OnmLkk624Y9oN01ZSSe0NaOMF8DExrHhOaRO79r7rBD+3DmjbNV832yc8jbke
n7L4mSmeqq9320U4URRGBOOdtpxlz+tWBoo3d574AdYjzEEaEyKWVONCUlLwuSOAIRwKanKA2qcH
mgu9jeKxHHA41qfh0wp3q37d74bFraDL1pWnmvq865zenPao6rkL3bh4+4cVYj0pPn4122kEpAGA
Hz6QTVCLK64pfgzEj+k46NiEBCE12y/uBJHu6oamTSB4Ib1MzbQZp9mkPozDaEySnUlVq7lnyCzT
0gm7EAQTzt44PzRmpsPM7RmmhDjiFMuBucS3OOvAKjrJX7xNpArNh9jDihI+ha9Kwx2PzJeIs0Up
ESDGoGcaZ+JP00g/382e2cq6E5SB/r8UVbfQE0HjtsAbFa/NxgVvoiXhV/6TLGq66VJVaM5drPWt
NlySW3leTf6Hac9g38Ffpnmwt+gSmAeDkvzFQ+BorlyaoeNog4OEnh1F+4B90flBqkNrvbsjiO3Q
4wBou+6pnsXKccYQY7/ocgv8S3potDfIXwFy4a/i1CamkChS9QWjB2yeyfQ/iVu2v2Q/Nn7BlSrJ
fBqDoUEBfVRiPJ7hbqFM1Kx8PbIpxanBB11e9J+Z6f7W6RQb5aKuKYBg2/ZgHOt/qKQVcGjWLrRI
LPmyuDEg0bbUinhEqVecbXBD/Xe4Wa3YPz32LrPuSvh4epXhujs/wfNiU0wOmUrapcQutHsqfhNt
mm4giMsVvh4rcrSpiahPWnqOnPBm9FREg4g6fqA/Xb3udbQr2g56Kv7vdeZylDuo5rfNrKzl0AF3
ZeMMtI81L0dqyZQIW0LlcwrS5ymc8RdfHFCcuhvuQevF61Pz1xQqOGoLKxRMU8dvE0a21aHsdbef
1X9NAnLr+JvrB4AO33M7/i4I+9uOGXIyzfmzaYs8J5zdQFs94jvhi2wyfgDyVcIIHWLDCuAilo53
0IQ/yMJwWRB7+fFyBK1DrhrmFLDW6+fSV5+NWjCTAp2+/kVMr42c7GK7uDNjU3ElrjPs/o2TDoz9
7UAjifeUy/adzS79Jbm2ylbVogaj+iegeqerXcd/M5rZo1jkFV/0fnFvzxdPVqcgq8jrDXO4qO83
E8TsxreaQB6y/fe/syF8bxfe6aC7FjBu0hdh+FvI/U8Qk8x+K6g7YoPYNLILeEt6CFpgxlk+tcT+
HXDD0HrRvkfGSnNprqvgGzd6qAEM+7R6XA3+KUZltUyR82nZwlw+V3EPDtQgzEah0EnkDxzyMAwh
zlhTvFa2fk0+F94s7fIb58tGm6dbmniEABHGBj2cmRnjRQciMbqr3D8xHOcm+s+T/dPxkRBmbSu7
89nqSBHpYSDf920mtjraQmnaWQXl0GHKZnCrRy7g/RQ2WIXGTQrW3P6AqhUps8xlEXiuLHoiqiaX
db9HS1P6sA3r3w+dCRTcBWEnCiGPiA79iXXCjtgqz2ofsl66+d1MRZaB0ZENm8KQ4QFAwDAg+NsW
G+YqmMZeRMNTqVf19JfwUMXSGkA8Z7SKKc7ZLhGjZnQZ1mRB7aa4a2nn6qpvLhm0z699JwjWXDVm
8OM6jv4xmrAWSCtlAoW2qsY/pB7qloZE0tSonc19uJopUcyjd+8He19KhQkt4A7nnHklumI4ByTF
Sb/ibZtvx3o6x/CGA+f2xvu41LYET5pKozwW345acS3d/T1Qoxo1sUszlB3uB5pWXzse616FllFQ
4INAjganBDvozAcEcLx4lOJTbi3FeJON9rEFHYS2mC+AzT68zFdB/m8ix/D0nH2I2Rmi6Y2te0uh
wrQbA8xUWIH0fPWqf2kdWlXF2lf2Axv8LNvYsp08NhzfbeFw5EezvKHqRNvm2XbLNLeEnbNKwiqm
3juVgZyq/5smwo+MPWYeyaPzOSsOpqSSJWGbZi76PVP0q6vzeNmNoDIIUL/H47J2eNxa1vAdbqEz
vdWTuAnX7wbZDY+XgoPSU/9X8I98LcwDpPgJAsLA8ar8HfAAgIflx3WDv7MSDbelsAnb+aZkvsx/
/DwQsk2eQndGixr9N9Hm+GgcDXWlA7AHSLUmwHs3guLZnKyiwadNSWkUNTTl8lfCInjwPtfG0Jur
tEyoV7ilgUyd3/Jr6RBmTVZUzm4cEaAN9DwtE/pAPvaP85AULFPaGk5GjBUqvipV/9XFW7JkFUs7
pVAywgy70fFr4Vskx83qw3rzrx3XEPGPvvJpCUj0b1Q5rKJX4hMN9EV3lkhwQJJMAzjjb13R+Ia2
N694hkw5AgVK5dSHHnMfYztNyT6DxMvjVmA3fl89wIv64ijdFvPFZrl+ErVWfnaZwWuiwpSd5cjh
YWYUTe/RaPljNgirAjOGEsFTJ+7U+rqt0CEcWo5U1SR0nOW7l/WlpZVg1yj/KH1aAR9yUzzj4m20
LyzPWKjDNOBfvAnmQemfhvFMV0J/K0VIvnpoBZwpzHiusgjHEh0W5FJqLh8RhiVh/4D7wn4igI56
cNsI0fjNxfMTjw2zzd0Sewo1VkCEv42fMAhWiUqSGIRm2M/Ztqr0W8m3wDrWu+Gy11D7PGe7R6Ji
9WHiR1WyKoFuqBeGCnto0aOq6RRFopWAPNI532XsIjOqBo2ATIx1zx98TqE7D/HHcqwirVBFuTNa
YsXZHFLXQx3jw+O4BB91XhxpB5DUb2tao32yNfCMjuegeDt9Gej5zqOZJPK0vhYB3ATGRFLlXv45
ba3qAXAsBMtxa6vmbO775QM2l6LTDK8jcnHSEOJdTI8lXVD2YkbLO2U+tD9qEGbHWiyfyaJqL6mg
LHg3kFO/qHbEb+9zYO6vpnz/Pkb1ZvndkyA1mIka1ChmbE5r0abNy4mUvTVRQ1xQfbfM/XRppAkL
D9KXaUE16Rauw5PWgCLCRfpiPuhzH6SqjL3cnH+l7XTuJ0fp4Oob5Hwso4SYc1kXKP509/mj+7lT
GjfPbqaD3szsKoauLe3qt1mnR7eLh9JjgfeOEvjABEJb/Wpfnhj6hjQfuB+LCEi49JDwdIcXEWVk
LmLNQwx5FRqJDs79y6efsDCZf1a2cLc2sWIFx8Nnz+masuBfBfnHGns8De6Lh5NIvmi+BZXvuyfM
B2i0vRtRn3r9q8Q+zaPxpMRXywguiS5zaPN7Qwdmoq3/DY5x7Hz32Ffc8HO/Xyb9pIfl+ty2Z3AC
zzmEVuL9H+nP2sU4B5NGXRQP/OWZlofatvKGEAIA5lJ1/CHGBnytnPnKHOf3vkQl5GFpmTsOhcUu
xzU5IfWDJsM49GfM5yTm2BXgXmOXjtyqxu3v1Q+M90cYh2pPA0CtEFlkrluGtq+TWIOMk62kM5cY
YurK+hkpPQQGNnFZ1pz0GagDRcYRpHizWF0Mhv6AqFAgIyOOC9i2U42OZnYyxgG/PbNmm0Fjsu1p
USffztaiivT7jiPvnsr5JCzqGpkEFNnJiReLCM077zJd+/qbUXG7WALvGds5Puc6JbCRt8wFjOXU
DtVRMJJarGDdUQZCPfjgzKh59DCzf58yEG8i/5CEUyMx1GzE/kJNwqbqL34ueHb+kUS8e6kK71xU
ACcv/EOHyVmHaDL+l/9OmMY0Iyp/07lDDeCEODXcXTOPVzy/B7iNecQ3L9wn3KmBY0J+LaBLFfis
vBZq1qvJRwu/3rA1LGlPIkcj2C1+JEwQ6KpD8nnqzQCsbCvoMePCLIFkdDJfYFL7aMtit7sNQriw
aap6y4dXRIVNhKfoCkf76NV0dzJRLLC7KyOHd9Ak96XrhKXJ3nxtCDANv9RHo8W4oIssm9M8ngwh
NW7eI95RS2drJU4OJP1BoI2prakn2xkBbCVwYpkYQgF9cJPowMoZsSlltaHjy/prYnL66sPaIVKN
GJtdJCZaPJW3qP67GTphJbbEx22VZqcuRN9jnlexUpeVkZXTjytfw7bhVM/vZE8v1VmmcsvY/u3G
wr+R+0jaE/kUSF82LzuVeB5V+M5vjQVLNsQ/wHpktHydDU6gTCNQiX/J7amNYpzpAHglaEM5IO2+
NnZndBup1pRzYi3Xmv3sfmM3IZxrN1RDDXhJYbCBgU2DL4Sy/kJ5IaZql+T/2mhdh4jDo+Xtf5fO
B1kZr0wnkLnVo/1JwS4Z4fq3c6I9riHpuClMyW5rrR4gxNH8s2YwRZt18wHh/Gv7Nw++qUvoqQPF
nPIUOLqoDat1q5N7XCRScVIFDkDlLOwUjSnjB0I3vLZd4o69XDZ/NhpG/b2VhgQqYMPABAIva0pT
w5U9d5LMOtiZeGat9ImhVlETZMCl2YkVYeOWGH44FlpYlol8IuqAMYLzwmk/s/4eGQ0Ru2jCLoMm
miyTbOXMcITyqgFaNtnk7tjvHoBKiNSNc+3X011NxXaCyO1xh8LKXjnCHZG/TBVrkCsPF89vyP7e
LpkTKkNlj3KXye8JEa5oKilsCABcuRRf8fZA74vbBZb522fR0AP339xxuuSirp8kHi0xzi0/BeUL
dDG7geQbOnLOKoYf/FIq9yYY3EqLwPXMCgxWJk737r4u1HUUt3ectqO1Ylo/A/AjSNFdF+KEvc6s
hsXWIShmRn/4o9rRMxM6JiChJQXQUhYakcMBCPfTpr6ZCeMA1Zf7AZqBLVbAt9qfDRqKNtFlVktN
tk/rvW+3WYilEZp6aJmEJ/nQFa7kBZOkBVWKPEWIEC2o9MQkGTd/660Idkk7FC9Dn4na3Te/PODG
eBhLXffbxHr9GNG2zR4j8IbEEglDREaKmKUyRqJ8q3dkYQYJEfK+uJVbQYDR4mJXoIUOAFYw0ABV
e80HGpxSn1+QtF76ZOcKi9loETVMzR79a5zG68J60f6fqypcadZjZVM4Uy/edX6ove2HMS89ePMA
jQN5T6tofi3YPOq6yj55Q11RArwpkO7Zt4HCgztZ8HurIzrZEtO838lgy0Cpz26jcG6Knx4joTQk
TXVVkC3LvqVcxrdxt5I3tqkDWv0RyNV2fIfX0smchJ6Og+QXzzZfZKZCyLe3bre9xXwIShQmgk14
ANigIElmixC3doRXiJEHJw5sOJeRjpYoMhUpEt3caMGJC+odpPFIX2d+Hb+bQsQRDkDXOeGXmkRC
1zwD91AvTZyp7PBoqL4SYI++LTieeVmo3xBB8wNota7x7JxmLpT7G43wxwVMSMyuWTnL+wMTf95N
HNv3wLjmJt8BeElUc5Pln2MzOZkp5Rajj4zG0oAcd4kpRzakPziFopesfm+p033NLMjqOskETPJL
sEwsaDf/gL6zubTNVY4anyWzMa9rs1LXaj1xsFhfc/UCD0VXJNZr4tv+SAKZi2qD/2e+uYPiU1eY
2818NPixf+WnVxrtTpqDfK+lke4roOdHfjcqoNBS8nFbGzuaiIb95m9WIAx92XSEFn35VGiAFmNp
cGHc55s9uhioPctq/omHutr/FGTfE66ltjpxRZmHrKt54vUDOtEJ+znfFN6M0NjRfmJB6IADbuox
AD9+DrgCge2D54GeFn5bt8/oBFEmsQunVW4V+KyaP7KV6csWCBJpM/UJ8U9uJW3PJ94W3t2kitAI
ug0TkE+78zPnCQzICQGBbTXMt0+fo9tIU2Z1/hHaNmH3EqN/k9GePO7wgCIKQGGIJKsGFwMjCH1L
pofopHzPgUWkQ0RJ8E9T8X1o5K8kfUGIrx2AFB+BDciIDRuh9m/iMOIyrcOS11eOhdnUDJbH3f3v
2lR/CSHUFy1P2sX8RZVt1YCfApfhqfeSGn0gK8sFNjVidBU7r7kGQjxN1fEd8H5xBrSW+AJUP2+7
aCV2UCyfaPwyL8XXrM2pb48ujBWrgMputtTnaYvN9Hj+a3eE2WkSlNK9pt0GiBCXbZh2iQrl012Q
QJKgFDrDj5TIi4J4iYjIJ8BRuC5H1/+rreFtbuafKmiQPTQS7toxwq96mX/WCrkof54mI5VqbmR1
agSGXBLhZ7TCtwjg1QbvpZ0pVGqorwNZ9krYQo8UMLNLAb0qtgeOerYiHusAsPghJj2FowlHTMBh
zPtmHc5l/hleqDCSCNvOx5XvOfRmTA4Ewcb6CKc6xTy6Clm9jc6/YToRzTABFjSepvOhVEJAJd9S
RQe/434guurOJUSNu4PUYV6sz8k19N0IyK7BeurE+mf6bUdhNzpzr8YxPqaZnv0yc7xHqMth++DP
i+29M0JlIsO0qTdKKvY7c3sFreD4CkXBw70AiCuWz4nlTqvFtfaw2VDVFLJ4R7LSluNdDAX4RKRB
RffireYyVWelmZszYrLhQgZdUIYrpVQy3UXvdRNi3PPa7/xAHPV08ytyV1FCsr+oBhZcewfwSklV
Iog+mdNbVnH0zta0bIoMIj83tzi4wWmzuAux1gESpFO6F6MtBHU+MHrg3/vA+TcUNvRHldrfyLcX
ZCYb/s1LnqBdZCyHpyTZKumwyRRV9DDknaJOBiWi+Dv1lMsnOlj0uPzQ6FG6V4MwQ6X5DPBS22K2
dowRoIXsKJ2mONLY316tSzDViC8ctduLMAPBs7BSZN4J1QPj4SssqzRsPeYzf6mP2jX2+Nca2fqa
9k+37Z5vfvN1f13iJV70KbGwt5FXzzCFxkmwnpNlgPlTik+ZpNZepgLAChLJSGZ56rR1dd8d+XBn
xPVanm2cDC0pcj6+sYAKPri4Jrq0KSVAg1C0KQ5jHA1n4iNPB3i4Ecd694pNm6G/WhpvHfH+3/Oa
ETi3sl2EvwaM50p4y6tJSLmro/qg/iKwZ29YEOz522TnVFABe0G1588fjXbWh2jrqoTb0ERfu2Pp
6z9Lc26DHarh3uPll/AJgbICQeO613kB4eJ4DiD9ThFeEOwZuQD9fuebhj/76EbHd7303sg/ZP+m
/weh87CObhpD/IL6LuJWw4jGi/vVWGqV1D5LjnxvsCJ1bFTjxpnytbASrC/iMtpY49vRrGNX6VRr
NjoBIK6ZwgVl6PplihmYbc/QKtNs7ihP7XsN+3cUZWMtlnFyJVvUG+70ShTRyIoczwBnHu9lmS3f
UofH3sEcrLTsHdvTyDcZsaAVmqTjZ6Uq629SI2y6hrW0z6Hu9togN4Z3TdhjqxplQnJo8yrVjzUk
x1TI+//Ugu5D0UMhgCddF9PYvZ/zVQUpDdWot6t9Qe/pBkLXeHMqBeX4fcPyHXHJvNu0yd9eyQLH
soJnqxfIbNehfOUPn2LaY67V/2vQJvmahMm/svRUpjW/5B/deafbTRoIbmostSG64Wy8WTgKSFV5
9mqZl8j67iuyQ96Gd+qsrtZhgeHQ1PHFNpUSrdtT3Z/dBYXYQO6ZXyrAzGrEwkrbdt79YH71DiMM
AIsaXYufBGh/EIOmg4Xn5zzUSukmX1fPixbEIv2y2oIJnhjtgGKe9BJzsiI2pndncjlCGT/LQ7zs
NvW2+fjMXQjTFb3EQ3vKXGtpsjQui7YHClRgMedyaqZvpFqPWGhcPWnc+R+IHr7m+QwuUP5hxie2
49aoiWkZMv7fNcGoKe6U2SW3JyutvKejRVsIBulUREx96gkg0iiRWA2SX5+3Er6gmN7VQ4ZxIXjq
nGV8Ak6u+PEQbVHUNXHt3yoVl3iJWyswzMYSsYYoXt10Ds0QqMw+Fb8RRV/UADLLUlujMsmhTyQK
yTAH27vEo/hoNDrNq7uQN6j/IOxyr+cMTh654U5p381zl+1e2oNbbGa2ce1qVy9R6Rvq2G7ptuHm
yBJlhWqI+Q6vZf5rmEJcIuhsA+T/dVtKZDoRpzt45JeMRTjn780DzkBc4WqSDDlsno8VmZX0H1rg
Znvm+IiCmD8/aqeot36Uoma9OC1KRI/YEA5TdL2H6UGC5iZsIHOeWvwG3bQV2pKqoBMvMDPToa+1
MnrLgLdXIcbCMxDxHoCGTInoKp56K7Uw0MgVQ0b4tItZBEnjcRdAJqQsvqqmqX7XKVjDpAkv7sbB
ifXkrFZwHmnq9umjhsiYxJlR/Z8bAi6bpYnVaXjxDoPPaNeU/TSXL4MN+xis04UqLS+4gD+dj3bq
IpBnMig9VinCVB7mHIO1qC3bO42MiY9ka0z2KSOwO7UibzYD5sICGckN0gy4whZ7a8PwMm9xEFME
Ym/23a/ggL6nx7in04SSRSOmgP0/ol4sQxkMZohbX6hp8br1MX5QiWr3hmbV0FwOmdvEsipw6B1D
9cIDY8IBUt5YWYpW3A4A+IBrP6OJYrT+tCtyktiiiCo7Ar1VgwUoHsj4fe4Ei4/AatiEnHA8Tcls
F8jgQvs0MAxXOCE+2KSh+lPdtuCObJ5GFy1NNyfPsb88LUVdKP7r5F+eE2pHca8oIplJ+OD0a1n5
oyvpPcoDxfIJ7DX5LsKVg4/twIKHoM4qfkEaBFJHpQCMced8HyJiYLtaZlGLRy0On/EydriKfzZF
YA0FNDgOeJNSu0Cp1ybiBo35dtGpP0PW7E/PgPacMq4fQU/UjP9S8nsfWWpKghI0Eo01bk7srbQ+
47ydrA0g+FzTo3rn4QnJBWGMCjru8q3TFXbxD2klGegRlSHJBmXkrcxwCNUWEYlctDY7ORzgqqqN
Fb0RVP07GWSfOP3m/TDWk8LUrX7lpKwW+hzgG47cZpLWHBsbWwFWxUO3StNnmw1w1YnrhS6dn4gc
tIxNKGpgV04t3jxqtUyNrzSjpjjzE6XwUqUQ7jKs/4YewXTQmVlQ6MM/7bI55ivlbToAFFTVRazy
mhZSQaAeBh6+IhWNdVv8DsYGIWbSAw1iama5974fGgrgzwe1tsJ6FZ9UmXiWemspCp8PL3mL8Xxi
sywqa26lIsLrKZ04DMSJR0PV7wvj7pew7x3XyqaVKobHay0JLfVZtVwTXh0TGtLfSP86cnlZAiyI
IPRQkeVZwNpOdhPOJVh9oRdSte4wtU9sBeR9ZtOIUP0NlXVYkLjZbVjrgC3TkSJlX2ggR/Xn2usA
ibPKeHuZ2AMbRLe6qvJHa61PUt+0hFVqEZlKSsYVpkmdc6pK45qUVeCpTxaoPnjorUdvOO0FtpHo
7+IldLZcZCP8RthJWX7veblehutmXKsC3gcMlN29HPTMxmplCm4paqOf1Ro2ibysgH+e83zl4uAJ
M/lj4sKBJM5q2K2WXE9UNdZy5lTmjiQQ4grDA5zvkotinb8A5Jay/kywVNIACAtETbaamH88m1DF
ZlvjrqdqpGkdcWiXkltrWdw9uTnuvIbmPVY7lSAjVxhtloBsumZjN/TpA773mWk+yVxsETrcFWlV
joJGOM9Q1HcQckVgYEIVxXTrGllfG6Z139Qw+CeOvj9vF5hh9nYeHv4kqbZV43qgu4XkvbfyHGze
1lqYVmo4PHzQOkRfzv4IVUU/ngXPDE+ESwyVvuy9Z8jgF3IyFDUewxNmhg2+0ZmUzp+VkPeBWhWF
CVmxifD1/RP6/9bpnGUoD+XIodMtnRq/zEmHrrcj54W99BjxnTGRODJNNI3ZUt/zbV3+1Ur2uh2e
fkE5Wo9ZlD5IteKkCrPOsipjXWIge9du82656Mh7Dxl1JwYNrabzRDuS/etva8vIAXr8BTcZaRCY
LiUjWwt1wBF4kds4xAJYYPzzVgh3lvh+I19KjJDle074VN6jAUI3BB4q9FyPkZ5jvHqAfN+vNyMZ
kXUhjJ0/vBeWM+PSjn0Mv6d2/gny0L3yHgQDzhdRk4um9DozWVc7aOpMn4aOXPMTWOMHf/OuhUl+
KvEzwZ3uorG8YhlEKmINlFfAxKmF6bPGRxU1hm8q/mllGtP1UOFCqw8u3cUb97acSUGpV/InuMb3
GhB5VboB3NIMt1mmFEqGqp2oABkSow/PiYJcwhG2fDJbNlAMyK76GWSt4j8fQJ3wOJxjQhKAB2/n
AWyP1XotmUSciBVAFngfmWCBohMmGa4miZkIclem0H6aU1ahDPQ9IpONHX6k6axuJY/YaFiB915l
+vDkxAtIIWbAQ2dyWhC9HhYwnhWer/mLH2cV+y8ZpHOfOO6livpPNxL1PJ38aLnWKXiDzTMslukL
X8aTbEHRfYHADPLAd1OArRiJcFwFHSN2nOkvrqz2TJU9nzIUoQLS/6VlskbuLn91bhQMnfk4s+da
k7aRPjPS5PegcO3o025dHWyN1HWekMsHAPa3TA0HA52mVx1T6tpKIPOioEb83l8bbVT60SqbtHDO
0j8bRxY1YDlVcX31EELZZewCadwO1ybxRNdr9+6oPk84IljPyPesn8M4dCb/tDw+HD039ol9cp6t
0utlCgdfZqJ6F0LmhqquAtX6ksEViZOd19pNtBJCSHWpFajADvJuaWrv2DomH+wLidOjejJ3f+U1
broniBE0LaVIGPOAS2DZ9BL1OjBUw2o2yaSGoN5RWaOP0gzXQ0+xlUB+ZrEuj9YIlF+/+uhAhW6n
UJ60qYpVK8yfm+tWif0aGvGgPoURPpYA6WofaNebSYYFfkdxzWhPWg/pGsLJ5494KfPYAwdtpkQn
kHUoZEMYOXvlEcXKSLJkogsTlf+BbCQugtkVaLVofkkG5BrqvYWjh//zfQO4pyDqoYvfqLrcmbfB
pXm+kw7n1E2wtLTusYTr8HXTK0ZwTZDDoLbtCiZHkgKIwQeEkDtL4wgxVK0zCsHlZvMBohT6GQG+
MoJ1Os6Cav8WhusJR+mTTNplS9UpSdLT5v3uSNAyRf5cG6YDOSfH70dQQynV0kGTgURisecAmCdS
jLJt/xwZ/90PJCX++MuD9Dotm2/AeoBsdvc1aTRGFJbvpJMzM6JdKiQImssousppvmm38rzVgfSy
ygsPZKlNxTSBHXOraD4kjNVeeTU2zSJXpxXLkHbys8VlqsJMIkEWMfJC7e3DZD5+hdhjenzrqEHC
IrB2+wWTU5LiTDk8KfN2UVkyCeroGuWMChVy3W7+6IDfPytbwxX49BmaXQjD0iBfgbiWCqZSUinP
0cdC/tMzj53eRHGpNlwAeSEe65brADcdhxhPtVe+kDxNh52ZYPIKkfnG0WT/DvPgClByGHkonwcZ
jcaPvaMzcGvyzTt2JJ3oCfOmLk2VkP6lLPZwhr0iAuZtrm5oiqcxCLCjv34A
`pragma protect end_protected
