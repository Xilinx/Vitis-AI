`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15440)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT9rrfVTtnv6Z/atBuUOrnyXqzLBAxGGYaY60hwY/ffGQIf0wbrKvthFI6ZGEGfeEUu3UTTh
GTNpQFyzwMmE49+wXoPi4G12NiVjQVMwOWh6g+CuXRroo7hg4ABvLFwhe7sbsfM1wsFxYfktq6GT
oQTV67Ks1LBMgWonZm6eTy4OxOVY/7Rvd3l4YbNsZKucsFaxU0Ge6tTOT2ZnPyQl/ZeRR4TltErW
TaB0AaDlx710J57Fw7xa04t0jtE5a/UDWP/oneyOsQUPPGZgrf4CbdY0BpBT1rjY50o+5OkiZ/jb
peYbJkVkNOxYeWnQ2EE2zY+xu3ktSDKQYCoUOMSFmuMk9g70cZpPheK3Xw4/LHjuktd4iyNSaWAf
MNujlSGKMyWYJaB0hrUPcwLA/HdGWyQoPsJUW9MpfxY9ffyEeBHl7NvYVGmyE0vkW9N4bT8Jzje/
3GVPEHsH+laV39yIpOkIaAJCm3sL0+RPK8VDE9lWhZvxEF1j37GcPHBYg+vgviXZlXZ/pyvq6pwj
2dziDsDett+JFerRZGNaYsUb6aiXQdcNZZJ6qn3FsVTJEdBprVN9CEcYYxtZEc4TWEdafTwxSPTI
GajjiAZXMGy6+DvG82G2MRLIdfF0IvgQsDdyYRbGTEH1OtPmin9G0utla4ctfavH8TcaLHtS7KQI
D9TdkLy+tFDKbuhdgWLOWCzNWqLZoiAWdUD/lKEOAYMDGy/1c56AkqjvfrGCh1BM92qRzjCsVyib
CGl8QRYNGHAiojij6E7ReKpAhWjoN6ucRrZen993JF+uup8oNqFla+9wDDIT9NdnA4dMNAXaxQfz
1f+fwVlvKnIRkI4ex1dYNUcXP44u5eZ8JK59+f6VqAvfg4j/jrSKfFHyfhYv6KJYOVAlQNyIreiE
1ugKi+jV+SkNkYmBZZ34FpezWwZ3c0RkDQHXyBMEdrfiPCVHjrg1K8w32f5T7nPKMbTJXTZf9UyQ
W+GT1TK5f6WRN0vGB7opu8oFIvS1tNorV8vHsnsNLlyiMFmrcu/LaDR3TM1Ktgq6lwD4tHbyFsBf
AGe241KorpAbntxph3qf+UunEw7+iqmjEh8bFWNy/f/S8Y67hoxuNPFcAihKr7C2cIj/fAjoRHwt
d9SnUZUGWTR3KvWiFHpx5RvutT2oRVL1GYdGfY0NqdCWFgIZsg4WkSd4QmLoWOUCspxyADq/7lu6
paBv7NqbJx2cl2YPutcfF/D02EhkJWunZjlkaS8xTLOJLvqAEBZBvqakJk5iHJpk2gnWgRp56KCA
OFD+bsgdZj5KZzr08j/2TUze3LcOfxZmb15+Osi5cJav6yBuNKOdESStLrUP1zmr1Q8GkJ1143gi
V49xwrDAC1tDyHLNEOy/N+CnBmoCA8SJqsOVlHOmQRq3IPmakqn+SpS7hSDVV4teo2TQupASk1P9
l2JPlqVInr45FNAk6zHaJk8UwP6mmdF5FcnEhc5SlV/ZLIxh5/eOaCxYJcKUVIiVogApe0pvt49t
E3NXcpBopsnPRUm7vt8pZ/eV+QLOE2K5kAQOIxSmUkDEtfelDsj+CfTLhrUZNy03GFD0GUsoU6rl
TPRnfjBLi81rfVWNKLpmQJgryK0udjvc5lz+dXNjYPVOKlsYcjOtKxRrhEzw5O2hurDDCHhrr23i
tofc8c454M8HwoHDZAbLhIy8De+bGn1VlAyQPc/Ji1QlXi8MBSuIdCWW+tj8vFYeCpK8uv8d61qq
9LiVBdCamlcBMB4aVnMnx/gSw8aY5k/0Ua26MiXTPvKHTN/FlmrrTcs+wkDtqihC4xRC7OBqyb2w
ED5a48oDMZEAoQGVbuK4V0pmGAHY7/WgonAMBbfZ8o76nk6+F8tadJ8/HFA+mwu2E5iNjje+8vcp
43UkyxOtzqzJr3YUyFHakEV07hv8tb06A/i7iqDa4o+PY4BQB9kpOfgjnCn9Pmtj02NtfJnFQzcu
6zUnDCb/81U0EVRbEP9yF/idHMerTfyfdgvqxxcIhq2R6ijm5FHDC/r2oWTW4//BF/mKVtvbZX57
dBqnseoekxgCIM2n4KYrIcFmfXI2RbFj3e70aDE+T5fOVjJmjaUGi5eBoTj6F/SX+r7z3u0yqckt
sc85WIvnXTeXZUZOUHauzLJwN0fhGx0i69aulY4DNBftHkBNznMZ9OGH92schbUzDJ+ZPwUS4J4h
GeUaogoE1ktBJ63bTjLz43YDBaOo9EOF2rITfY1myGMGLwYs0a2f1v0ZpsaMqYBR86nFbOWWaXDT
rwzqRGhlzYxBOl6orVd5uJVLSk20Pjx7XRINF4Y/4GF4fMY5rmmi6JXN7Vu5ZOJ1zuVwQivXqoSZ
b4fMcyMTatOAph9xsn4Z9zJf40b5fFPr/0bryHxykLfUHDkKY/7+cu06Vpx6dJeEbAIQSTleIYIG
Jqey8cc4+TlZwog4gFIrv5QI17BTiyaKGszT6prqlYH4N3KNXi/rLU7mvRx4N08HYxm8mvqOFgSx
J7PJ2iN15rbvIkf5B63KYFOFo7SzCrG+Gozjp2eXVpkH9z1sBE36+ORJkRfZL6036fuvZDV4FLex
/y2yXCZqhUBv2fqRGc15V3oIJs2x67G+OdaODYelpbJloZxdOwZML35hdqshUazGWmIGSupx9XgN
hEOzEm2Ke4KYhKolTeGa/GvajWfqpIfTH7Vy9GTc4tviSgAHrUHsaAoi8yfLc+HAz1qY2vXIqo2X
PwrDT07GlG6+zVc+tSlrC81ZWw6EnO+7W378qWinQreQ8vgrhSLXNon8WPMSphI/tnNyAaCEPq+f
tZpbfPjnmIb2isdr5dd85cRtoUzdpEaDocT8+PQ0vTgoL9wsNRL/8GMexGAT7tb/qC7GtecHJ7a7
osqo0t94Og6hV4+8IsqP1XXBmGenzVRZALx7g95liLQVUDP7FkVT9FMfqMxa7bsPB8VrivaYXZFQ
R290438AcdpmrIHoZl1wcMB5VzY+zhjWPcPjos1ISVJ99EPq3yWX1NA4mMtewEtfmrPyTNJKd3G5
b/A0fGTgMkqsZ2gvJGmC7KGL/lwzF+FrgEddEWpbmgkYloweu/9+CT6FwipD/6geQ6WmQTxL7MpL
ErnGvYNRPKDAeQysz6Wv1oDJnfCNNsb/6Bx2ny8y8upQCsOYZ04UTtLhFmEzMItnz1l/yEg4fdWL
OUezPIVXS6HOiy0+iv78e7zSopCwKhLX5vnGMLstL80G0jsh21Cy7NJHLbhl80DTit8bZfoG7F8E
zCKQHLpsikYyY98URtQPa6B2xNOT3gXipQEUlp0As7tXYo3oAIg5h1F7Q6T0wY7Vo1yn2AkvOetv
X8adrnkIXS5dqP5Odc+AinFIYZe9fly1scGoZMBQpvoaWrmZ/pBPW/DrlQD4n9QAD3K7sZXfOLqe
diEr6ak2JDa8O3s8XS0WnQ80LK7/Enz5sZ8a7nRf8LrsrOHWk252TBbef9+n1hft7wa957Be41uh
oSJBlY4YJnwKbRIizw2hoGcJM1UmsHy08azEmsLCnPQlAPdkSh2y/l5U1Va+AhfxYTRRnjLAYhfH
uib6xZGbB5Lt4sFtCMOulFEpNuAjc3LIngz3gy7Sliokt0pM1FxgisVbxVJfERxCfLaOWe+U7k7r
IXCcfj13J+K6fzAFtQeygW4znpRctdoU76sBlLtE+AHvtdBLk134CKuCEjwR4sntnf9s/kkHlXxh
ZjsdNIipjUvjaxI4pF0mLgOO86Qj54pY3TbdSbs93OX7Y13kekQCRZZKdeS1KYuIcl9zDoTHhf6V
/tIxN5feD3M+MLs467a+/c3Dhfa3OWRF0EW2u3qnVOyQc5mhLmn5Aladtrd9PLw8V+C0bXnsZ0g4
dKvGf2BGhSCQf/3obfVAiG8d3bA2nw97ckTH6/zYoSZsTMpqig/m8ypkxx5qF8XVUIhnw5k5LtLY
Rh3Uci1rd5IiqTu4xEP2E8r7377Pwwi8I4XWiihigT/1h8VVOybdA4rEoN02G2+zCQMQsCGYm+fn
KZtg/C3Wq7Gbn7tMPdv0dNY+YaHOoW3Cu+/6ayIrgHrR5Qd1y3tNBZWKTGuvoY8FvAE5eQAmfcgk
ztK/tVauQWdq1h1OOFjFoSrGcR0QmtgNrDXiKB0HYEX8wmv1og/87yTiLkO9KwOXnX9scuXCCc+n
kuMP42MUiQse6RRstuagj03J1VP7UGT+ahzHe7Z2eaMMrlI4cKnabYz/ybC7OFDlmhtXyg9C/89C
AyemjaIw7tW5Auv4YRQZgcA+BfNz1QEQJ+DWzhMeJkVMkeVI6XTSVrKHQ9qRbhJDZ5Y/2PzHCCwT
NrXCFGonfrVObNZ3iWUPxvvvAxfO2FRFyglQzQfqIFK2EQQLK8tgOwLROTtiJ8+FHGSovuHT1Gby
j6YGtX0OLk9w1376vKA+vrQTl4+x9ZBvSWMk38AjJFJMXszruCE8R/ZlDfPlUnUneGFMsHvaHs2/
l8vV3X3CGYBTDiyo6NfEUX82v/XpExUUj585VduO+UMmBqnnGnlRirdpeRtbX9OYTb1T5nm5OIyD
KNmBCGwA46nKuwAf5jAB9+0yPHInLDDHBpx3jbKNTQUKHqvBPt/BEdqaJCJAnOwbCmwFuuJErYui
CFJzxSWzEFuybPGxKvkgls0HasQ5A6I51AurA76bkBitGBAFE9yDOxWjitEiMsE9Oru2YE9sFAO8
/DjG/GRaFSadOqOw8bJjnSqnxm6RTkkjKj7jUdY/Uf4//vFYBj0AzFCTBBEEqihtSS38RzjXnxEX
vcDZB9ydqt8wR5DW0lIK0Nz6eclM/++KhDGz+kTgDbLS/h9bOwUrHL1xkqJ7yuvPuBgv1TU41xdl
2xAQEhhnx/3FfWzGjJn1M8CwBUDqta4txNM+n0k9XQ21RXHA3JeCNvkgneQjSVhvBuWhkED1theg
rDgy7B7IBJhBLNaIdyfq3hIazz4/LqGeRIOGUHP7ItOLg1YnWvaTfCkpFMrh1tiW1ad+DW414MhW
pEXI+aqHBnB51i0H07b7BLufPemsTmAffeFqzcQKEE2qO9PD2fHsATVHrioh3gaCmwTfsGuVc7HS
UJKOMppG04YeKWNsX30I9uF0M4WcIBUtdC0baDIoDN0ufT8Cg7+bTDjfi5qlG5nUIP917u9E3BV9
ik2YkefNBFT/41lRKjfKgUYDXwE+pGdKGH4J3qRrLA+NfZ/uD9M/lzVoqNV8XpUCiRdDn8kQamWP
X/W+AkfcSYVzi9zZghYAqRC5byTBHrz9lw+N2FiUM5wAP+u+3P9oXgxh2lMQ9IikIh2DK0hNU8s/
5m0ZrsoEWg+j2CpFJWbSd+5Q26KFlEE1ySkURn6YUTaxQZ+R//dKr7Agdo8LWyITg1MiJSpcgpMD
ZQOgVSVhk4+/e0v/q/CLFa87yGyJXqjnx14ZceeKa7ECau6yPb3HqnZ5mxecM92nvjbTjUbC7pW1
NLB7li8z6C7GM6Pv5qWYZqwmEYZZ734ob1q0IRFBB7AkGOawIkhKlVUOZ/gkVwF7J70HwEhkFz3/
QoTt7spSJqDCnaevQ3tulwovGfXLsgVSuUAJF2f/qT0PAbcKSJw5JxcSyFEvIuGVWPtkUY1cdslj
JNUjnA1DVzO8zqMQH9eM3ZHHJxHe8MU0k/2EkXkYHLNVioTbiO9iuDJtJWFGvOBkO4N2h+0BQMml
HYXfFEYoGcwrTef24e0RwjCwonSfZMiKqKPHi9hiVeV5Sw8vpMBlQfGKjHByYJmirurf99ClSXKP
d8WFnDOgmj/HicF8fX+Aag2Bq8apLvQK3brf4WE9KL2mRePwJs1DRmPt+sSZ970mIgDUl3xFYCg3
VXijr5PWumZRZfN4cL8f0mh8OOt4WpLCyrUoyXKNMJc+xP295ivW8o4qSWrhAU1lkQ+R4/x7jWk8
bdz0f6ZqbYK1QDUr5dQ3/1LmRoULnrnL8rpjvIMk0OyV8ig56T4CH1flmGAOvRys71y9zOYw5eGh
c8y/sutiwxS7H1x+ipl+BOqwIUBsTjFYhjiV8sb5DXJJesOFgJ4zDKWIp/B3+Ys5gRQYhYLevgV4
u+dN1EkVQp5bst6UTNviplLsVdbcrRIAcsbZpzYa0hpZqL979QG7PdSkKElyF8OpMKmj9RSH0kk7
pdLPn2Sj+DVMXHXC56k59+pcvSUSCdR2NtNjog3OQdv8Rq7Yngcldk92SNWPVa15XUww97r8RYtp
pjon2/u3uHknV//leSG1SAc23IcnYfkyXF5Jt1aLHLpS/MedZosBAUILFNiUV7nDJOn7QsdHt0zL
mRbre5H1QEsvenCWlt72J2Y3mbr4zj6LMnZaUUpuKB8scfh76HsV1Im04Pb1+duEQB8vRZF2HGaW
/pzkbZSYILnjVF/uXTJE9Wym94ZC4w/Roh88dsD4U2W16NAVeNB5OmXEQqlZNMG7E1GVSVyA1iPN
B9vkL4G4md8zIJOK2K/gkvbvyoZiOmL2/fEl+sFX6eTRO5pgKmiiEUJ9lUtW4e1q/c2YZ1ARpZrB
LxxPHimRRBx2hZenO6Ku8WQAS5l1HlzaRlsx9aCUsUirM63NwjQgBL1TPdruLd7xZoxAV+fhdtQX
WJE0OvAHUE3KMkdjlhGkLwX4sq/tPsgNt3zpGkYME2bj+SKkKWDAQ87zueEZ/s6buSWBN4SeLYsO
ATN2rKXxGQ8cVlfXZoyCwJnVyrD5ZC/mncyNxyxdBulNSXXt1BcLJXd9HpRrgLvCfhJZuwZGAYS+
kVUDXEcC+aGn7uAXRHUJf+wMZ6PBvJrCWdVHsON3/VY+RWQbwdyTyG2JWuSdP9pnNWcW6fG5wdNl
f375tmhtBPiy5DWmwsWYGV7hhfcZh8i8jBUYzY7DcKJ+YpiBOkeq7D3GrbkwN8RcNNV9KAGlOVUI
vXxGfvsHLNsRi39/qg/+ciHKHI8AuOrFb3xVLEvUkzH4CIP9Cd14RmAPArTk8PNu1TVMRohXS8Yr
8AngvJ3RGkhBb1gPtm2/h8nFXL8BL69CP6tBxaglCCShw9y20G5Db2gzuD69SryULj8Js6II+NFB
U9Vkvyy0jmwCh0ZNLyCLiPh3JNo3yL2u9qHxqvV7Hu/OFO2Z399jr0Wz9yFaj+FruJXizu0GsUdB
Drtgos3LXKfq40XIKRnQl6NTm5WsSA12u9tj8hHq3vzI4QbgZuCTrLK15l5xf1FeBkvTnoS/RzSU
0fof3f3GtaqQdMsD8lp/BseevYH3ZwEZ25mgKgm+hV9ZWlEzRFaiDn0cApql+vjZBjgtZ1LARctG
1UbIGjZ3Pk57aoH4MOlN2SLAO0dhQE1Z2PbHTPkNC/BJVgt+AUF5imAT4f4DkCqOJawr8OK0PH2K
atfKVNWeT2Ys0smjRHnCuLa52jPD5B6uLMI1BkDKUqgov2Fe1lMO8CeaiQYARmIUTjDIpbazx/jC
X5yV7EMazsatO+nOym+xFN7Nqev1+l0hfAxSCja8/nmQt3EBxx6zWMacL1p0QTARDLU9Ricab6jv
9Mbzohhx2PWlzo/5zQibteUzSPwRwZSO51KwB5BN6Q47PwY/tQIDe2O7iKXYZtKpoz91i7Oqdy1P
brm+Wm460FfIRNKszEbFRdiEbQiKLLnD8E61GB26M7tr/WQ++rC7XxygEORuINOdDkf72olQUrLh
Am1yA2T4ujD5LViEZynpO88z1s2fS84M6LpP8aqR+sp8LGb6asL3FaJ3+0ZKnwCO6jtM9jT2ylqn
kOthItubSzAsVHDEJ2Cpf+9TYmqbZMlINaMJA1sl76azPLbQx5bsPmFkAZelNCqCQjHw2UBs7eaE
XkEQeGcN/5H32rakShCdFU5hR5JXxF2STP8Q3H5XYAG7/4yDDNgxiJ6+v1Tonfh7Es6mlXB/4Fsp
PaXk0BTD/w9x1O9gu3+5Oxrx4oFvutbI/JArAjqsZLtAKqjQzp5nfe2T21cFDd/U62oAjPERLswC
e5yJGZACs6Zeuh/BHTZ3h9rHygPocMfUlDKnZgViUtAcn4AOVqxcYJwXEHNQFH7YnJNnxMWbHzc8
IHvLoZyCxEtV1H9A2M4snNgJr3zzrGwDRe+OmTezxL/un1ZSydaRKYPoxr+ctUNyNSAtz2/A3IRZ
97VvQX5KWJria3erlkahQMfEqQke6dz5kozj7Z6qXKHb5iFx7xpTtnjiQGEeWHW4o8bxztHtMF9r
mUQ4DxXFNXzn4Eu9SQRZhUtzQPuY55lmY71Pl48Rv2npL+ltKPowa3XPrCw2X/uPRMsArK3nh6iz
0ykuSNGQgDA48TR9mTTBiJx+Q70LHSF0pXPQBsIme+IkxvoHYgSpBkpd09dzh7mbvmhJ5Z6+Kn7w
7ljWGPATW/L4+lynVfWtHmGuppm5hfEjsvBJwzslddVgk6BwiPPM18GTBiB0c8oY8XEgd09PrIwL
R1VeWzbhrrqRCY4IDGnK2zRjYdUMg3PfVBz6X6gg99NgtUl5OADdX8pyUK8JR3MEKxSxzZo0hneO
17dCSZNTlBv2kvoETowzA6j6C3kc491EziwUFnqIq/hK5S8Lc4ZQIt/NTAr+0Ja0EjBTxEt6IBC6
SMP32qlqCcJgZQeLm9tHHXMF07UU7InRD1FZsQRBIG8IIHBH1EN/F6VQKFt/5fW+sbu7+ettnmDr
CWBTqvhOkNmHIojhMzb9xi+HjlSlScXZ2EjL4IfS437RD5MfWt9CvUUgqst/fEm2x6DfSqYISiv/
eAwKIAdQDTpjtYVCvSQXGMwL0oPwRNEOcOlHHk1XGWHotNOB0r0l2HbCWpqEt7RPuw3Gds/gq0p7
QRkVKo/LIX7w3grY8a8hZhpoj0cgRppC39g/lHK4mKUmI/J9kqrz93uWjqRXrQp/zGg3KRiDCXKt
pjkLYC19SCIjWlhzpTlBKDliDrcw7lW5TqCF5nNXwUdxbIdPk/kXhJyEG+QxGa1MXBDTzcx3B7T5
hV/F9ycQ/L0AKHb9SeBeStjgo+NqkpKzp5BXkKpQxfpaxpftA19Nv/4xU1LXYcdV52Qqz+MDulY0
5p57trEmAktB9VRqBRFWmFZhAKsVNynJLFoJ3u4dY4+FqtNflUEF6rL77f3GDNKXOy8hEmxajdA6
JZNuQE2Dh9jfKObh4IQpd+QEtGEMduYGmRxLI6kW0M+hdVnvi4jDQirXtKVVulAPh4kSHCnaneUl
eJfX9m6atR+phMMC65ANu8B9I96KRVAKNffpg50QEgoTXjuKKxYKKNln/APFMOCk9NVLcFAYad6i
QmHNpHB07bx1slclYhZDkndt5UXoqIqlK2DflXX/DH8n94x6hRbJASAANZAZ9mHPbsMPn5javFLc
EEx94sb5HwAXMEb5ofWGhMmU9/2BLEwzNJH4MqLc3kerLOZynyhvn19VcL8qdp9tFUVAL6mPH4J2
jSn30cKGfgwVmQ8hlPsCILmt2FZp6LhvocFAp0ZKfV6akBKiTUmriRryiJWhly0PocDZIg3cMXCH
dLoR4BZXPfO7krovFNNVOKd9Nr9hm6itrdGYGWg7DppsIZUQRmTa8IPyz1t7PHP/5+fFOuUdAzAA
TWMjghL9eYn2Ptg54Fe9JjHScx8gutr9UYcFj1thCrO63hP58WobeAd8zzDaDgjIMMYsDS6zHPgv
1GCKpvpIwI1tGEFs9wC88JT892HbyrqSp7FsmRdNvKX/IVwbXzM7ks1wopDdj+vij7xgGGweFUPI
A2KbEnP3Rc4Rax4BCCDMm38LuZ0wM5cvuLxw7frX/hwE+2vf11HLbxkf13O7bqoBga4RL/Y6hAtY
Ms+Jx3xUNd5ZN0JSuD47/g85J/NJUPqxOQLvusnQ+8ax4LhtYmT+armiuJQe7K6Oq4pCz0z02vvJ
g4Xqkv0oX0vrsZ5puHZZuQJyzz+a8mawBIFHBG/NLOEJaipw1r8Xsx5WKlNF2cRaEEDQShqh/aSW
w+AkYRj+Yjg3j7bXeIj8dt/MXR8Mm5Nz1G532sbFFTA0x3WXmK5DriqqVSrifDREDn3A6BHB7KZ5
ly8EGYPpIuvWlelmFC7uj+cVYCKuyoDj8CDGsaaGey5efa5xpVE1Xnn0zh04TmjuHH4+0sThQhA2
HK6ti1+BDEEFAuiXavAICrXjtloPWhvXIwHPcbwSckiCoXkCqwnTfVPuyqS9O/DAhGr1i2MRJKA6
sP7MZ726h9NzHzPBadRKL8gFrORWakWPAV+kzMfVvPTcCxCyWB665HHoEeunkafuX2OKvnzQLSyN
CItSInOQvW7sDGdtcm19glyzFmQCMlY0P6bwHINdU8ne3NAGebYTwhJBoP8QUmE/Ckww8hITrayL
PvLFjy2JFbUvm3KviAJyNVlDlzljV314c0g3EluVU/GxR1WtMVj+4M+T49VZBSHHTihipvCyQpbI
MSN0Jtr5o86dX8X8tupTAa1BNZ2xqeap911FasijZ4f9SJ7yskWB5xSmX9CK/DomLcr9ll5w4hIf
WGmPw8GUHdcNkD7YGLtgBhgQmMFcSxgJQ1Hvuy3mW55NvpqQkaYUNRaHcEtKvQ7C/PzTKXzKhyLA
emjpmf/5Exi9IIaBOiucEELmpGQKXh5pwGVhNLQD5dxh5mUXXk947c5TbsawbqZ4flaiAGZ+Daph
zscvKXQx/U8jUyaac9G0ZrM6gDvGU5GNTGsPQ/WUCptsPWOzU8BYLR+gxUdrabyw7OD60cet5aMS
XGxnOBZUl4iyfmiRy+5WRWTw654LnNcfBlOAgMzDhJ/KkaTNGrrfugNsvYeA+Bo7q2OHGRgPLqyg
Ji02cEacxt9rjEYsfK5C+DLNl1eAufsK1WXsprnZVzDZ+JeVQFaDqRo2u9BRIxvGwWRsVrkZoVmw
kjpseXO7WfMV2FBbhOXIxgR5kX5tR85EvfAqolNxehb3WnYu0/HtGt8WuheAzRUiavhBtyEcNjX8
AogE9FlTIxIH9YA3DLQDov+HN4lT7lwfFXeEM3rS0r5+KMWIhKTQCNS6xLm068qWy+twNttLg0Ru
Xd8leEYdEqllMUK4Bk9bl36s6iMSiAFDDa35Brjl0dClD5HlCJGOUel/fbrikGDWfEasVP4RTtiy
Ui2388KvlhNBV2JaYBTiWrQQbVlxrbUKBhVIAXZcZRGvtqbhH41aER7032QNmAihKUT0PEq1qoXb
dKns8BF6yd8nEJ7HP+ThoGj9Y4bmRFNheubKJiy2MCeosjKERg2jthZRYK+79/ZpI40TGR/VdFzv
FjDBfJ+7qKR6bLmkzzps8MmaP1cQONrkiRjUFCtbKxSjlzvKYI+8OtNdIN0pufoE84leAsgf7DKg
7I3qw0R56jqT9rlHASTydFQeKIeLAb4fPoSUt3ozGAebvW9PcbpMNGP5ZF7Wuq+pp3Fatk5h9BXP
M16oI836zLImuWRdiiWw0hzv4lVhRSaeFiMa4Jg/kScxEpSxRexNrFvmJEK2DvPYjU/rShrSjcl2
Cs+RkyLdjTvOW68slswKhtyRYYGM12CDLrcyx2Rv/aH7f0ZvTksNd2uPd6erfSwx6IAt0jc903Ro
QFIHUHe3kmTHhqSds2F2NejHHuO97YaqiP+4v4LjydO31Hs/nuUVLBN0/CRtAuOhCeihzJKEYW8N
lKcVvpj8VlEcJdEle3V0u5a9EFw8eFVG8N+15owNQUA2Cb1bcqibbQXtNjW2g/95ILCzKbxE+pXi
mU551zvgFyY+mzqTjO+xbM8orC/8D38sFLzAsXj58SBTXCfAaCgxNrKjMI62+xTcpbIjS5PIFwoM
KtaKGyOI9jDPYy3+BR5ucIMs8uIuQ/+Q6Xb37drXpgF3+NS6sYP4hcrUiZLmojMR3F8pY4Dpni2e
f0PCDLtzeiMX1xn4JyyWp3h90xO9fpVDvfmmvhLzpTLWPco45hqB2NsJmTuuNT1tuY98r+3umK1a
xuURUlH5/XV+dmJ4QkuXhfRnRRTDS2rCqoLbHTnKFaC8TR8/cjLRfHExF/IMzOu74RaHkUnnSH5j
5UIXIO/xfWCwn/QDlaUQJXIQzhMJgLoAg+6WVbDr7bEMwJe7p/qVWTuqUctDqKYya59cCcIdgkLE
6UjUavQPU1NM5T+TejWTkYNAMW+PxdcjYuSmsOr8DDJw+nIvqxicYzuNakfmkeVnw0bZ+5D7mLSD
SG2PLzR/vTAyN6YJQl76LiP0/z5JVE7i/AGs33qNCyoLazQwVd08hC7vpyICUd1ym7iSx3zunyAh
K4C5Iwot87Gs6oWnbxcvGFgbegX2LPjQB9YwGMl7qhw6lXLmaSU+pY4Yi9JpX6yWDkKhO9kPenWR
Dm6uH/Vo7ltAyJ092FGz+FdXBKoY/yaJFBmsDYuCUAZiILvebotQfCTcid3htbRouUKWwlRF8lCn
gIrX9VTEonncjVynUI8biXVEtG2IQE4XLj++JQ8ljL/m2pPp/TmdfiC8amIQroxAQt0oM+JYMdE6
1mjNAGjv7qPGYqzTpQKwwz8sYtG01vWgeviyxRA2YVCuVEp8lrF+SCrTEtjJ1Jn79pJCbAwvDY5+
u5lt4zneW5xdh61Cb7umGerlPa83+5aG+llYOl1FiIerY8WQiHsa5UOzjGcOGIIfax+b4nlIA0ax
Hd4amevAu12hW2q+myHgYNz5JumtgGhmbxMBC7PAF1S0UuRKavz9QYmKX54wu+KAiidPez25+Q7l
U3iPN+5VuAjsoszr3OnaGdJLTtCJZOQBvs8EK4YvK6vb57Zp7GfRmWZG1aQpPoqSkZTHS20XmP9p
dzjYHLBk0uqjDWtn0XCVGMUYa2JPf/A9r/tuTfQgUzl37QYAzzQnv0z/AmwFpoy32kf72L8hh1M5
D6cwg8GcJIBkAuyfCNXFL/kA9Ev93uEX1lqijgOzzAFoNOUX1hsPjg9kLQog8vIwukzpDC1m4A09
8FJv0oBssyjTnwmFaowFDIgAiPoW80cg9sIWEhXEMP8mU61a5Dx1se+WMXwtQZ7uIx/dlsefznwt
3sJebZk8JCHSp+qMiLTUZ74lXgFF0Jq9pcf0k3SlcB+bNufLWNOay7F74VKVSbpS46pezv2qtA7t
tvLTLX6wvovno7ZizXy9yKwK233ANAVxxI/6Y6UZPEA6UQpgl3Rv+heiwHSd86Jq31D9jBaXGnx2
7g4FLB2umOzJP2t3X7xnSSszorK9IgYOfLGmfN2w8EA6xusGm52WpSQJfN6frcRytfdy+iJ6aot1
YR3uAEwuqsZxoDmBMzE+Ju2EGx8aoIuN7ZKzy87W50NsTahxjTaxMVFJKQr82xRbeluShLJIRpDN
xHOxr6hUCatELNE3OgTsUsrq3M9QZbrBPwvCPG2P1wLGJNVFLo8hrTGznCmGECmSstLSy//Xjoh4
nxGSczJ7lQM3MLOL0589ErkNeBxGcAXoD14S8LGU6rHJLaRs2WO+J3F7Y8pyqFz48JCYWeCj2YO7
dR39OOktiQPRut1ogodxwP0eumDQTgZ/3W/FWaX07sACbAoTSsCI1XVMEVgDlLfJwpG8QA9/lHKf
+prEy1noxDUQhSNjzXedZr2FArFka5MM+mfdqpv3ZyzM/1AVIgDa6VbMYDMl3+S+FyMgm4r17QC0
lkHfesk1LypEk4tkHrK2zu26c9NXx3rHi9U3ZJNWd92HMq/1gLNQWNQjCKSO8ZnuSUv5qeD3V5ut
cggN20Y+mUwIEFfnD1xac1c99Dv41f+WI+h75660KQMwG/BtIcYp6ttwLReSliDpcHsY8YA+IY3p
+xf5W0E9fdSUWp8sXkoQ50sgai5qFAz0tIF+ybTMrs1nqfMjKnY6Z6wfHCAHIQUuxeBQsiKIkRWV
u1RftElLS8UOO3HUIaiNccCSoVsbNBn8Rdu8FO1lEA2GzpdHrvbBR+fE46EMy9GQnaz6QeFc5wGR
AhySLUTrpHHDpF5x09zw6qIuaqJqWpvkQrNpygZM5RzZREf1mkaH3W0L6B9gCFCC9qOrgO7OV8zI
mhAPq1ucp6R/R0F4sa5cy4Yi299ygIZgEiU6lN8LnVLbfNgF2YGlIGhG8IgQhZZkLkRlXA+5vStF
Xnm36ZDkscrLDTa9cp3zri9LUYJsOL/Jt/ZqSXMteSxHpIjP6bPv7M2m2Gw/X5QOXKTo2NZPp5ri
SzsrJwGWxzT2zyerrb6jHOyaKy2ABn30Qm7D005dclwuvKa3633oPVpccG0XC1XsYnA9Tn4CYF+7
wvMPKPHsrByxcrmePNc4h9mSxS/eJxM/y/diWVzItsgrZbnkBdmT5gQmSXxZFgkBkzaX+FhI95b/
s5MZYt2OUsiJ7615ykHVNmuNqdVm/ROy1FdydmDnhL2Sn2E/s7I7Nzvm7BxAU41R0IjIUjefuprP
QP/629dDjg9PlNppkmCagPl1HqjYcVe2HmvJHmW92a976LX9DA6hRl1kbirq9MbSUxEINwxVTMdr
cP52KriEnqivPuLgOjIDVUittXDx9ignoRepe0l96UnxN16cozUqCoKscUwIJhYZCLz5rN+idQzC
bKqfp9F7nMeu9y8g6Kqo3m9Jolf7a9+uu/yy+j1s8D5yzLiPExIWthh2fwXaYiMkqeBVMiTWOr3N
QDkEQ2la9lU+GrH3PlPhGRN+Y0ym5o1+4f3/oDASIBf313l+tXzITNiNPz9K4a4yNo0Cz0Lh8K0l
TLRleTjoQhTI5lfL4zFlEKUWsCUePXu2fDF8C/hqVu4MhD2K/sfN0QXzPzzEMvrOzc+nXzqnbyqH
MO2Zj5jS+e3ZKYUwB+oNbO57GXJvFH0ot2D+q5QZ3odRCavs/+m/oyj15kallLv2/vrmG0CWIYbC
juvcxdiHWdBQ4awad31ioLiQhPyE5O3Y4Fc+m34lZiCzjpDlCBLlcpnRPtjIU01VA7N6yNWAeJnY
am9zE2TNJKg4vBznDeJ7f4WwXX58WOYEzpq9yiyfe0ouJ4ItbPo3Cs8iu6GkI5AV29f+QTRAeHIF
ICTasFZxBVci8GGsamFlMF2PqdFBLsDl8nNaLtNidtD5sYF1WpjevcCNLMRNCR7ZW/S8tnJiJsvO
215iZkBHaJYEetpl2TLx86KtnMsaoUsQl5wzijXgZ1U9o3bSu/ikPzcIMUwlgkq6bp4AJEiuMrgo
ezEBMzrlt4HZQp1aCl2uKOsP/Yo7Cb+4+jD3nr6lM/V3TO7a/XA8dry1wefCWuRbwVZQJ2kRI/e4
+NQSw8DOX8saDSGe3HJVp6rirT8CdXIvgHV5yVTx6+5lQYkXyCxhak/SoIZoTgQ/WNNRpogZQ06P
xCkl1QNIn7foMspKNg8kFdyQj+R26BOgb9LwB7IiniRo8omMru5C0r11NZGf5pXDO/JTu4zU1Kv0
1GWuWaMHp2ffkoOay5eEWBGvM0p5ErZMBQSTTskYKjupuVmLx5zzoBmJmQ0RGoMmgOZW7nQfawpT
ubDuqaIqHd5/1GyZMQt6Y6/W9x76d576XQBsx//drLQNQImUEJ2i0nIoVUORrBw3bWojPpQG9zQ1
NK16v2z0/soK/ShF+uMg0QE3N+kn6ktkOUAUcWbW9nXFEoDlRfp5OLyXGIXx8FtbdsbE4n8LmP5f
stZ22xZHBi4FbvAOawOv8sVl7itvklijZlnGJVDvvXnBa2zCNmP+D18ZGLQ+5ceEF1gTJGaPEYJU
T5SI3MV3r8XAh8+4kI1Jc/nxiNU9N1njy4e/SnUHaurzVnQZlbNKfont0FULwpn1wJp3cAa4TH4Y
mS32IYEaJQ6Q580TKh+NpS+MNCjGHTKoG84i1z3sFWyYxdEUypwt2xy070G7PsN0U6iBL7vBvCCF
umeov32MHWhfSnReSPNl9XekrCu5b3n8/j2hcR3B5T4SKS8ECOcQcIti17YJHdiYg30HxDAlFLUE
LSvISOC6Ty/e/BGYY2Er7hhKJFa0ivk+YfoqejzbpWLDEj6uCztQk0usrRutO5iVVb61g12f4aSW
zSQUvFIuzAfXLTPhP/llIBc89/wHJzABt0Kt6BxAgYAMHSsXbsUPJT/ZXMkMv/60+BARUbX+4aoS
hZyazJAfhb0FhH17NtO5XUiZPAXO6DOPhCXbuPRkzGHD9oPeKXIVJ+BLMp8UbpDfwyQS3ELkMSGo
9kTZE9LD+Clh46r2IyEbbRG/r2qFJOTWv/RQTmD+neKIEpHqMDFVx9dZ7R4rVtyW8rhsINRUYJN8
xBnEcUhnPw8So5MXngp6P28Ms62I/m/dzhOBt26qA+tocC6rQJzqkZLNaKKufmVYPRx+yj425kRL
peG7ZfB57pQXsngkhE+g12+PuM/rpD5CDUSE8zehwAv4qR58zmIoN+V9o8OJn0iT0tgh0/jRzHUG
EDa/iPiE7bRAzmgsxcERagX+ju7r8jRchQnjEtBGgGULXsJ630ZABfwRvzKsRsg0bWDgsnodmyex
+MwcFlQyF+mP0P3Isu3Du678jLifeLB8ro3KG4QMOUr5q0XsR+HyHsNxdnXgbwhTT5cIvolzQGXS
6xskO8nVmJnbHVJUGaglyEXJ6dHHc4naGJsdh4S2DMYPlOL2BiFFOeRoiBGgJfqw80vDj6NcGltf
KKTgiMDBWxydK2q5b9nVKT+FjvycFojadnpVlMmt8GozjeZe7R4GV/Phiotg8Nn5d1Ov2ZIYa6k2
Ki8tQQxmHPPpc0GkRjcMp0JchIDUevPznqHrWBEcLjABCN21uUm4E6sXjXNECfttMjRPeU4oMplF
wOuouQvaJa7Sz8Fi6rB7mlTEa3tNAJIZJQCsRSU9rTUIX6mUr+m0ecLM9seRecxmmW2IXAy+0K9Q
Jl+BVJsxg4d1Xlcny86c8sJq1UL8fGVus0h1It98XExI9VvXO1z/eAXoRXX7qC7CzEazvSkuGoVz
SM6fb6lXbWIoNfGwQm/IxLTX5pgH+fQeo/ni2Bkapu61sacf19/kLCnkYugeIriWQ7XQJiD3vPyb
8Kd2sllAqDjR1xvp8lWE10SHtfR5YiC9U2sbmXvWhoAPRRpScxY6lJCg3IKsNFj+oig1nxv8tzbC
QK0X/rjUKS5i36JTKOYO4h2D4+oZu/c1Wx5pDlDJ4FiwIzr7GLBHMDuOSU2f1ZUc+Ek6+RRj4I1U
8TlipT8VJQvSKirkt/CkpZcrLSrljjvC9DG1YkyusUecv0VZKPg3odo0k72LFXLNDIL50qM6vavU
0Qb1ct1Vv7M3YIJiUUrEkc246t708+wx8BtpSzgqdtJlJFKsqOi7B+z49JHZNAPrJfKsE7Wpslc1
MwYY9/WgTZweYHKGS8MI1kxRPMOvtSTnH8R+kZ1X4nSCxo6wuqHwDYUEsnXVBlk5jqC3H6T7T5AQ
Xyt2M3GPHmJkYr7LqrzFNrZVhnx98vBbgwTSjBIaFjTqRQxlHgNYbT7PQxA+1c93y44by6U0GX7j
0+g5pifYwStTb8jkqMd/LBwI1AaNc7KA5scjBpUEo0ARyjD3ZYYsjR4jczbiTkQVSRFemejnv1Aq
aZbAK+GCtOl1YhrrmpMrbH/7e3p3RDhJ7xEeGbXDOHto4BNm7seBM57hQGkzAo0tiR8ttuukT9mc
uAIxIGT850qFiYDXUryqQeao4SV+GRn//tzLU+JmXRLur418IjSjhMjg2f1MvApmr8BUgsWo3ZfT
8Mp8ola9MQghqyCRxYy/vErVLAAIO28DugiLblFKXdyxlzT8MX0m4QAxTgliPXTQchwV0bAlhe5S
SdGrIB4uFvZFcxMopnHW91QOdmm8h7PKfAoSA7Ec99Dz68WorwgPdvAtUI8XpB8THn+OxsSbQBKO
uT4H/zzxQV7BAgsDaqeJXAgR40XePzquu+ExjJQKeYRYcr/U2IJRKQswzx4VOoJu3vtmBqCpY2ls
JKHdsPONfih0LE7V4ilvpohd906Kl0qN5UDT3mto68GqgvQpzkAjmrxQmUQ7Y/Ix9vvyHL24OK4M
OD/Hz4vXgEIhZOpXOlJOc9orQZLHnSwIgvqI28PMa+PxKbiPxy1gvkXSzL7qxCLkOJmYu+zI9CAu
ksV6cXtyOzb6Oj6Zo9tcDeqXx6ZY2KNI2tKML9ZrJ9JdVvs2fR5rgEomJvbXf1qvnWMaq4Koq1co
H1o5V29oaNqK8OTt8gaTqi2i3s7TAf4P7Le6MyuH5mVJMge7LSUD2DIfL/zMS69HLMF4M8eHYPcR
vCkSziPWhYA57aXEj4x3dbQcIT5MFsagbZODjIj5EUy9v/en6bs9pDMCYMMcb4TX6DFg7RIZD21x
Q4iJ79b8qakhh+XcmhYWWodtei983nnR4EWjB0OqCpVnWpO/i+2AZn5N7jhf186yd09EWu/nS1QK
VhyXllvHaHvyOc9EepWOsaX/4r2Xu3Bi3b5FbafXmBqInL6aZTD9q5rhKBuYgoxwe1odxRZ3xDFz
vXgB3CA2mrcy7H5oi3HyBs2s0JvzXdEmmNE6TLN4KPyC4H1uQsLtPLv4nInYJlvIQiDnu4LbitBl
Hafj/Xql1gqL5qGl9qDoxB6W3WnVbyrt0tRD5HcKOYRmDMf6xmcoFbRJ2BAeoEjU+jBd4h3bVER8
OzWX8G15KtuftY99I4PzHumttJojCAwbsNr8gri/hu9iFtqe0eNKdFgVwENBuY+riQH1DZ+/o0DQ
g5wJjCPrQasZibAwu7p1/u6tvEBYTtDQtUwTHt7qbOAoq6kyr1iP/UvWq53HTpI8V8SirHsJaDQ9
dJrKfnk5nL+1qX6tjy6LpgpXza2+5CLUh0P+t4t2RlDIIq4i6D8zRIxBJBq+cXzgQDUIeDCMSaAY
DdU7WlvVRPxZmBQ4cBm7d/263YKlYdjyv0cSKu/hsGmupWv5EovfVzJcnBMz4KUy7mQRTsvyg0bQ
EcSKv9crbwtRl1jHs8pd7bhx48kA5J9tzxnWSSkDPxxLY17rN8i4zRhlbaISSSC2eOjhfMyRTTu1
Mhjqa4kr4DzOWPgemZX0T/wB4A1eaHGFNNLyS1/2aHjmks8neL3yDJGXPjnC3ynY6JTMqePgE5fK
Hq/5ZwPaSyZXg9NLhq61vjdUbe8YmIt6Zx2cEAiDK+sF42hmpAUh0FCPILpFYthY3woQAFqK67e6
IUib6fzypETL8kvMIFVUuzlwlFeNzlkItPLadsVqutBENXr2IyiAcp4viSvCJnj00kYRn6q/H9I/
VHjMfb3zBDYpGMsxyAvnT8E5SjeOoZAug9hR3OnyBpiSO1JntnRaoSZrh2b79gMAAnoOR2a4vw4T
ZxRkGzCHqv7cH0nI2AnJP59sKeXhBREi+LPk8gGRRI9bQw11UQ/59lznCX0b6oCaOhhxYvjkJGro
LzPd6moxvEF8I6W0DtO5sjm9mTmAGSu7BtLUJtEIrilvDB9JRHV1e32ZeKU+OTWn97yaKxqTu9Aj
qaD7giyrI+NTJh6BDUhyWKRjJKTNJ2RFNbdl3sPkdu9vngYMJyzIwMzJ5aSHsuwVke86fkufhTSy
MMVAPx+kgZicBn8+LNLQddPBI1ra2dFIQUCKwEZ/bU5ZWpwcv9zDXGuE9OpbjRhhlfTLIoBrnZI5
f+5OpkKxTQ6S8s/Lsub1XJ3d/aF6wtPI8SPEVghM6wXmY76vM9yHIrnS67XodIWKbKURTZnEbuuN
YlIi6ezOjgnDV9FcQ2EGlZ8BjYP5IpwJJ7sU+9JNSGvS+b9p/zTSeguz58Vq1GaQCDowXIyJgogk
bI7rPSWq2BeXANBaIm45OQF1UXahaJTwZJ07r1eb1GGJ7rGhX7aKYyUThbbk7vePzvpWMn80r/S2
ys8rlHcX/MdKkJagsQhehgMecjZKq3hiYn7tTa19IMJNe+Z4LdfmPJtjYdUCfbJJ1HHws+3E7tqR
FP0grNL7fsW7NATpqstDK98limu3OZiNFZHO7v3b07o2ejB/Odqbo0X581U2C7I4CrcIJGtYKPLU
+Z/O4aydRUw253EnaHaMTUCFdEdstQh5hjNXVgdeX9AYj2E946MdQtHSOPYpdXdhUYvWKBy+DF3B
q+VmgLSomOBDYKVJnD0WtRG3XbcO5xw3Q/iLjwZFHCZqWB/CE8bF/xDaS7FrHUJ/ntvcLAZEzr7m
Orr+goI3x29pdwsgwbQguyh077gP8QtqDb9tP+uCre93r3xisf6VIy6A8VnefFNsMLTsMXdu5nF1
9ORzhJvmssFg7QxNh7gELH1bcxsW37pWN+twPeAUBEMARbpxKvqXajZFjXvccd+QBmjeqazB1dfK
mTXW/8iXChneJIIq2I/qh4ewv9TqaaQXoZSXUX1Rg/wabFEKw8cxWmMLRchnlPB77MB/qoUejZ6X
HQjSphQq3IJwfJsBiI95UG3upDm4g417htyKVfAviAJEBQjNr8MaSUVcmP02KvDa7NM=
`pragma protect end_protected
