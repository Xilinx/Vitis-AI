`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13936)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54vV/P
ofulVpU/WhvY+xpgCU52RqLPKYMfFff9yUOEehtUiUhZGSzUVF6noO4URe2dI6XnCVkoePRjsKTb
6ZOfn17QPnfWT3Z2tty0q/EBxUNzJAk75yiPJ54WfbN3xPsyRAUv1yyPrY+DC96LkeoA84yBIwhu
Y4Pfej1l2xijDAt5yPImyPYeI2KaoJvDTlYgwn47lmRzxVYJWsSCDp8uDCZ1WTuPwlzmGvQkEe2/
iegzSaw89h3y73Im/DfYCOl525uBDWJd22hX//MzUuWSHys4DRcY0c5dPKHVppBer4e9ZO93EOpx
8+td2bct09NcrI/PvBI/0VwdhEhC4y1ooPiuYM528wK3LLHLBKzQSL1hOWv7JsMfllZhmcSLG4Sk
zmSX7CJyDBrC0joAK2Let35sxZbYGJyE0xKmOfsmp5vugrLW28woKbA4etZVT+gRpNF3l23tXJNW
U2JbmxDosXpxQ1f56DEzT5C+Y7mkEtUsN2nzMHU02CcxJ1h600grUKU8WxbKcDSKNKMGdTpnqEX/
ADT9BPo2XcsAgqKSXVV0fWr0ZbL6NOVMD/fmVu4q27NSNjC+0XXR5r5z9d2/znaU/VtxkFwP6cjn
Mv7wnfniRaZV+SRjQ2aPiOnD22hNu6sr2XHEHPLaeF5tonevtb2hubT5p3EXCgmA5SORvCs5RKmS
ksK3rK/nkEz1P+JZUoyQVCCpWspQFs5Mz3CSM2M02/9Vndkh+BPWkpddhgR0SkIblM6onx7ZsQg6
tFXCFGUZS0b0kkobYq6qVfno/m5+KtIE8XG3+wvpH7oh1mDG3yXaXlqraq4UwR/i5jBFPmctxkbQ
SscdYOYOzt7xS0f2uvP2Iust7gMzYln/b4h3yO5bbIxO+ixu5A/vHOW1ScJj9fY00J+B8ifBQu/g
sv3PpvqivsnOV4E2XhUpvfwUQ/XA/YQfZOOTUQaF9+A9jMD5b0derekweQnkCMNbNVslbgW04uS3
YmBQmvMoAcP8E3vc7Bp9H17cjAKU8qOrz4Y7JjFhsH8isWUJa7xIY/RnMbyRuRgtTOQY/NsKZcLd
uj9ZsV5ybE+tPMfrXxeIH6inUZPqbFJJ3gu8bEmoXSmbm6JNgMHMFKc/CjlV3K2KHttg0Il4FRnP
ExTe75nl5mTZ0dAYGhwLuzgVobu09OCflyajUnLBzo+em1Eb7wu1AaTUo50stS3SccU8Jc/3ckFs
IiqDwAMgL44Xkm21m3PSvFa+BwN7H0hUAqH8ZfhIGptcziG7vEZ2ubcrFRUC7dX4I2K1SYe5eOq5
RonzZNfuTZKSrXy3EUBotkVJHw4P0HDO0zGQ2GvkufceIynJIbIjibWIBi2xbQorNC00tYgaJN90
byIDEQlNvJLdYraRxJ5LWJHaDsGTw19Rsrd8P3Sukr0K8fNHv5yt5TbNHbknl+FlgDYjeWPay3tP
aALPe2Zuva4zSiSVd+v1rS/+FFxSGgJgOZlAvSbxUD06abUQ8wU5lVNC161vZnua08xdMUffmelB
+z6rif8ZS7zEaXP2TnTuHgctpgUgT8LB2XhcXnN9sGdDogGmDQMLN/+RAsku78/Mo3aZpZ6H84s+
xfkAUSnF9sY18Lz1nv2lbcnUUXsBRNkiXfg8YUCvFR94/qRctSgqDoi0sVDN9lU7hHvsqxJOpeSa
dtMVoTIkC9NouzWKduqEGqQh7DU9dQSso8UA+zuUYKk4GUiLTZTNNhjAur0NluxHtPcUFx/qUhVb
fjG+AcRzIUNr9O/nP8kpEgHgRMoMMNY8vnanaRUpXkYQtFZ5RsGs53oyRoU7U5+DeQT7ZLoI08O4
+RqO0BFj8IlN6q4Uh5f8IQ26AQWt1VH7+c3bHDqg01fhu9+t8Ae03rqKemC3cyT3OJlrW6cLgAZz
uznRVOfAOvErwn9oZfgRE5QvhUqpgOSr+5DZZzvgow9pb3VkurBKQfqXfe/l1rer5T0IOvoxSu3b
UDkEsbPWEozUFVT5iErXZO3+13VYWgIAlXYkfvsWbDSguVxquQ5xCIS9NsUPHw5C/A66Au/Ufj6k
V4ZnDBw6mPxN0fgVkRNTEsb+bFB6QX2F0e+uAgodE1TCxzhZtlUgNL20n/fIwk++xEI7UkUIy3cP
V5EYYt2k/YxQyZi9oJwPT0JAVdsXQGTJQBRo6bg2AfXrOuHmmw+TQM1vplA8nRUDvnGXWeAT4gNT
/L5f2W4/G3T6/7Dkq7JMxU3Izp1qovsj3/c0mMKfCLdhemL1P7r6hK4+w+ZNmnp0TBrSNPGHJm+d
yuCDuyLD7HxxG4eF3VMKFu5xNriOMr9JrQPbkrTPLIue7nQifSBLQz/dn2pHMbHfuXXKJ+NGaYNv
p03ks5jQsWqM0snXxUz5kU4ClhnCauplPtcDx9+f6txw4yuBBzr3/BgxVr2TW/wp5vPx3SsE7l7E
ojNtoyjCTluvfw6NbmRxlyTlS8q1VQ6CgTLfBrDCBbQ8Zwm8oKNDetAirrROCjL6ifDh+1wiMXLa
ggGA/c8+FdZIOUQZ1yQg6PPRLLH2UE9tZDRk3ytcwYjACL2pMq9mRdQHC/TJmIkvmf+Xue+6AXsx
dZP0FAX/12PuMsBAESFliPd3Bs97SkkRrGJfI3OEWQjMl7NZX43DOfazxuIyH5SBQPVCz4PstLEh
a6WqauuyH9HNe36QdsyE+C7b0vglgH21VjvmliTLef6sZzL7kR2LHtGM2C5YAdjR9MVWBxpiUxUs
2nsT0NWprOVNqHX4zfWuO1gFsPqho7f1kREqxqBzYZiD+H4sUh5Is9jXIIIFBnZc8aOp3gtPM4J0
rgJ2tJlDX12iMamWbKPzBo0JCx9Q5QhkKx3qXILiF/lpXUIahOYYFWiMEbaIxwdbJykFfn92RY+4
JbwaoUuKnSWHgMqxoyweAsBYgjUmslNS6uOr9pHTfxpzO3zvJIF9rqfFYJ+PtaxhDTWCcVcu7jSd
H3AJpTqnHK+D1JzGmCDeaF1bZi0C3HrCAqK1zztzTgsA06GE3LhAXskz8fXiGFcYAsyzyeovxUFC
9CyEKLL/WoDgVl2txTekEYhO64TFfQYOrxnfrGR2aNlmoemWVuZ5p2xFCz9YGcr9JtHirTLGYsnN
wX6PIeH+SfRrTvzje05xQ6UaXuUx182RapkNZPPqoBUUKScEneqWivipOgUDImwTy9s2mdgpQZ6K
vp6+6EsOkCoZyQpSOuEqNPjYVunQBC7QI9dhfH3HyIlf/x8wrII4yARD8/bXJgyIF5fv61LU3ZFc
JaG4aV0I507dBMTfch/Tqw89c5aEum1QXXXDCddxw1voCjTQODk3ZCbLOhT9AWahs/hvscxvNb8W
HCxR6zTcBQsjHS2jWLIriaKDqBKPEprcTGtvdjIddoS3FN0SqXSTiJqTLzyX07khSKnny4sAAh/q
dRrfYCAB9LA8pVoUhNFwJTjjnLAFZBd/PP6H5sy6mKo7I+wDAFPWjGnv7byOjs755DrEBO83j6Jl
46dq8TG/UvDBtMF8lkcYWslwE0IQJU/j97CC7BudrDSGHAOkOA66C0Tkiz1QibDXmgBedz6s+vcq
R88NjaUKl3Z2aeL3Cgl2h85h11Q3FKIyY4mR2VpDDwa9SpWT/P8Vg7M/elFsXnVEF1toE/AYs03z
Qs5uCCpSnzmnYui1nmCBZ4hTD6uiB568WXeyUHnBZDERQ67xgCuM5riWpcftRpo1uSEqX4NN+92A
/ZoPt05rAn6c5qW0IS5DTt/hukhkM9DLzsGtChBpSTGBsGowf486ENwrQmBGTJ+bUgRrLMuB8D2n
O+Fibl52GLa7GP0gic3ogRv0jmvmvrsa0sOJnfNmQOmZef/pgrc5DHL1mH5BM1Md1kKU2swXlwYO
rPsiHny01c67f38d3R0oFVXpu+l1zQVeG0iIaTELnUSuMSPTSyCbgQIhf118Rkca+H9ZU3dPfHtz
j44K0xuzCawrhpqT0r59/9bTMadLx9whO5aJz/SUzAr+AdFD9aHSB3IuWdmTItvmYwHWnSEKzblq
/uZu2Ij/JFGBswQGHJsievPa6PsJawRjCCd7g2rcKplNQIthv0QnNyI0PFdYVlp0irpTq2SHk4Fx
fAV/vQW75WqIbfByCK9FIiU+bconWLmXy34dSShsAyUfDsNg+kh7o9toN8ru3YsDZ/1j7lZf45hp
FkFGcqPnTEAXKupgTsta6QZ50Xoe0DJq63vg7XpOuRYRLFmtqhLZzov8WhsDfYbKgTmjjcX1P+1k
p8OuU9rGlitzu1f7ilGB4SuAjwsRXc0Vjzf7VeGZzGne9CKRZxl27/lkL0cmuY/UQYMb2KxOFNXn
/MO1l6hcze2d9QLB39xX2WxZV35bXEgUXHn5zUXsM2v6UQ9v+aWEQjoWueo+5iQn0Y9004JbqP+W
2YHWFCp5W6QZy2HTgqPPvqOlSGSklwGmAKyP2/1vC22YXi7yB7//+qboxh/LcKNLxJ4pIWdFD4J9
0gA8G/Exa6AkRFq74XiAdFP1eCZfjKFgSLlelAeUFzcwEF9sahF6Um9BNSlT+3tHF9g4EUjIzXES
y+1EIqhhxXgAMRrdrgU++Rt4iU7n8kI6OnS2HI+HUE7empqKuKRLAmdrVMkM3Po1uHdltWyrPqYk
ljCTu1mQ5ApZFYKVPuXC+Io23JgIHz2iscSjbacdTUwtiPGUApq/cWFEVoguDxssy9M7L8H1NCFY
SdakYcrHpekMcHOiQlccmisrp1Ju56WEa13rzxNnkFIDoOvaUKdFcGVJ8YXg5Z6Dyy0xnb5depHR
yHAT/mKS/Jco4Kh05HWA/N2a31ahu2likQJOjBHAV5cSpGmVRVPLFgspRK3BdnfEEH+35H4tW7PW
+4TJ0ir0OxDif1GSKVLu8Ew8QY2e3LZ0gHgdMGBE+x8huVywnpzv8VDfKuLX8Otgz21JJBrdqNza
Seh2B2G4rLAKPfcH9rFgrHVX9wFvnI0Bjk+82p3satdFB6FCN9bKtLIyNQOTInWe03g8xnmw4IpP
aqeqoBl7ByLDYXlO286nirTkl7h+NgXKdytDXmvr6WFm5AnCovKMNqvD0sygfRV/wXjnKBzrQVFZ
x6PZkTBQxgBn1S1lzX950aYZDv91lrfH3uznEK6Sk7oiuVL6F6eMgPwr5JaQ8SwKYAeA8nYpOrfe
RuyLl2EZynz4lCeFvm0FM29lGDUukEINgDBHEV8d/ZBsvirbx4vZm/g+3CKo75YyFQ70Bxcdb8YD
YVKj97jhDcha4wz6dOx9li7WHh5TZtxVn+NonBJSD1p6Z/VpNPw1epiLX/L4sI/f741sgEx7q828
+iOMZjbz/z9yAt5rp5PjXG6NUOgMsY4cQ3TlHcGyIT8f0MdAEh6zy4TbPbwaHdMo/aybdVq9x1N3
h1gSQWuJvMdqKoUhLvnc6o5bqZBNFy4oSmio9+LOsdBAc5h/N44L2fNGnugP89muWp1E5sMW6nmy
KIPUuaQLvykyEyHALTkHnufUiEQImReKEiIDU1cDALU4mP04jb4vzSlAhbpikEPb0EbuIStX8B8s
UxIEqX9Ky/a9UXtG/PFt75TxpMZUmzWaiFiO5TGCK1s1YrHRclwqCUDy9Kz/rRpScZGRC5BsxLKv
O08MIKSYyyrM6eUchyrKBuWMmowdGX76x6qsHa5Vqvlb7wSdHlt6qbzUTbwZyrbYTR1pLECEkQ5b
8TPSQe+0kAyLWVPa9u/y8ytN4m4k1xFaXvJEFFOQTeOkwljqgNndypbm1IPPUhz2KRLnwc+Sb/nH
cFtisvztnrWsBQ8gC/EDBURl48tI++yd/60w1+foJcV8uYhI/VpYR9urvD0lYVv6CHihloRbcPMA
48cy69ODp7KpuWOc1fd3Sozm9UB8EPOchHU1hT7/DJ74eO6oxDYXnxQk9mxCz+WfEBuXaT+swrLL
0Y5v7BLVhvmOP9O3l2sNdtWXisn1KyVEsaLfkFUH4DEQhsOuLuUsX2w0C5zxO+kJFlgUU3pOdbSN
qehXlNKCBn9ZH8bBDH8wCF2rzYtaheDAHu+QUlf0+ZgFmEp5DhE0XYVFRtIzc8s6573NaLGlYoMr
Zxhww0Ub27Zbu6tsl2oASiiVdRj2Em+mk0kGmmHcV8RfR7hfYOv/opqbAvXlA5eX44m+jqDkds+3
tg3EmfSChDJ48MJGEhwGDHufI9028/WQn6OCKf0DLP1TnKT2nhAYbeQDD8msevNpZxdZ/jF+reya
phByxW7pKSty6gGpPU8Cx0lyfRYhxd09ZHkhqwJrkXetwUcP5iklvfEnrDD158Em/KuKicnPCipL
iHa0G3moMLIriWK5FT/Np0MApVgpnAZMenU4OfWFCSUSvs5sHJoEzdCML6ZOQ4dchznregR6YqIE
YADawaElNqBSHKbTFlwpU6di3ILQhrDjFzqV23b8NTOTvvoKomMh/FVzqOv23FW4uVgjRGP9IaWb
hS1A9bPNSwxwdhhSHqd0tS4VeP2vafRypalT2k7GBAGI1w/R5zu2JGH4Z3z9IXYBAMj6u3HIrIIv
sUej07kOn80SswVhsfSVcNfWsQWsK4IhtxqRz9HPubbKNAKADbo6Ezzmw1Jc82EUs2ko4TJ92Gk/
VfyphDhZJNRU8L2CO5WtEbzyBfjBTtW4WHtmi2kKvFbBVNI6Ug2KErsQmaHQ7ieLvT6JEwkcgvCj
3HZg6zgp80wEt/13YTV97eiv/5t/aW6fplDaNpBbjaU1ZwJPpYGUJkqU2M42X7pSJfypKxIvcmUm
OvNSTXtxDrafeoI87akMptCnRHvwieOPLW+Q8GZBlfRyhTU6PMfMmmwC7ltPB7KoRKJRuIHMqv2b
DoqWHrH5JwmoV0pVGG2bu1r1aXrSfdLWqfsYmIP/k1s7ccXOpYRvGNRaQ0j9L0FzJA4mBJJAFnCp
2tgS6EvP/6IvUgdX6cd38ro56D2xPlmpiq5EWUafXihF8RJ09J9tUWs2r+0fu7sLaHSG5RDMT7Z4
2U2ng5nCyuaT+VjliwKOD/VAScIlZ+luYcWEki/GJChybOHTssQBEUa5CsSn7kN/LAUnECZtnLC5
+sM/1G2Va/+i7KvAgFpBXZnGkz6nTa0AAWOBYRFs4PnR11x6uN2SiBCrgvrvEPuXr3pN9r0wzs/6
qwENraL5xDeEhNr50Dds+3FEgOCnYLB9ovcTsSLEwN+G32Wi0gQKAV1XUNu5YSCo8aV5gOCrclfh
43I7DLMiXG/mfCAmiH7easInkocztslY1EUxnHbYDBPp4Iuvm0kOd333LWWjXUNsyfJAdJXabUe4
OrFPPLtSurVwX+zDC/nXiYLiSmgmzBgGrs33wn5yJ+hE0j0g0sh7ycx6B9h/F+Nqet9vjWFG6bjW
VJ/RMDBWsI+b7XLRTVqZ1OR3ynIS/ae/JGCIjXveliaMh2xJm35LX2Px0AAGXCQStk/pE+fAHoGP
7K0xOU4byZ1KoTlMlNYagfiftRmIB6poL0bSEg34dtI/XhRx96AptWhQ4imPE+x5+2bDRgazixT0
6DsFR7GGahSQvSrFn18DqF4wos1McrVApRdDfKmGqhlNvWx95qaSJQ1DERy/QsecgT9lig0POLgI
Ul3VE08yqcYAuFrNYVVn1O6CbMDuOcF6CsT2crSbUQQq96CxG21SrQn8dkqPWMIwtg5EqqfYicRE
amyky++qetxrHG/T2v9Z8vt+GNv2AM3G22xxL77TLly7ZqMly63mVSV0rQpgcRx3wsP7WCpVInGp
zEewLqmI+FAKwwnLRt75DWdo/6wTz5NBNAhJoIejsNnk/yBYcEvWaoTsns/NMiHL8pkgOMqYOAh/
AI1U65CVkxe1nJWebsLweLc6jE7vWhoAFiWlp9f6VJkihG5E5k9XSy2YKLniqCHsJTOviZN/KBbk
JzdX3/TLcyEsL9YgbavKUqaLiqGrSD98J+5ZLTbLr21jGtPo4w9mJ2MRRbnCVQxECCPxzGL9Knt8
pRSn4mDE3d8RNVhdYTBCIjvhQz5geKX11dBdfUhc2Ej66XutUDXiQElHRxNy9K3gQRsy03jj4NmQ
TZB7wVlTi2U7cUTLAXeIijkAeWp3dcBn1N3dEzA9HBhFZtrRteVC5fikfKmaRyaAOVDAiZeCw7Vh
8tClvIOoYpoPkyCpNI2NwuaMuDBq5YzToiCZhSMHhaPwRK3ELwqgO1yiF1tKzEpf7EwF2XLU0mAj
XqHnMDuXYe7nVREd59UsDgw23jOWN+iWW9s0TWCJjJCZMHirhCLCx+Z+6NjOf+d4LhEthbmMOwHB
8qZqkk2iwrphHCPfGw3/ZxK0f207mecm07T7NeEkByWK4IICCBzfVqk6UWOEgpZo7GA7Tf6tDF3I
DqKeLrW5M3rwKifcV+lcEZ8BPPp6RHOdacZPVLfefZsMxZLoXnf6wmGakZ7JPX76M9B/7MH8A8ok
lKQe2UqrQU8XwSDSf6LGVYt/qWP9Qv9JMxORMSHWB03Uw3hLfTAC0Q3lwuZ5FbfT9NIsRJC/x2gf
Do9bhbCDFGCJ+1/QnFAaQhiNuMtMiOFZq6hqH+aOYbfT9VOAPRxTYPJFXMukOetkISUWY504fzI9
OLIXIZb/2cLWRERuSjnpBdSl+cgMZv5XYVaH2Cshq8mA0fUqQ5kywMoHLjQjoOUG5o0tsnYAif77
fy+EzQkgCstEq6DoF569EfYLmHRjB5po5edupfMgM3g7B6TsGrs8/w0FqCJ6v14AV097AIOnOfTR
hSfpkmZL2v2i1smMi+4o8veP72f1Rm7NdrNHfB3hjYCozCIjSS+DhtaTwPOsE+Tz5zC9pUQO6E8u
KbsOLiLyQXREAaJKUhgCuYxCEtxaQsuzUpUR+RPTd4N5my2Y+ZZMXfOJx2dx3Cz7/WDOQLLCf4xH
ZrnGLtyBVQVC9LxGoBbvHYijEKdH4lP6XSmlaZPySdXvvFDRjbVNNrX7G1Xt8seKTKEFQkvtsBtC
Nn/LL+TJehDAPtvs9TuY6iq3OzKlUT7lT0z2vGafCRdYOy+Cu6DK2ucHKEHb0zn3u6CNnEZd/iRH
g/WmDXbXwEKT0x+mUdbP8lDYHUIA5uesDL6Pe0baZdM1wk3k6Q/LwRLbG6H92omqkARtCvPwX4aG
QFcD/NqjLyU1V+/vyfKmomAYTLMQ1C6zt8zLpwbyunei0tvIm+RXqgc8QWyJXjj9qATyvPV4CyMn
NJ9sAWqTssti+H0INEtC0MFhWHjBAhfxtH17cl0qn3wiZ6jpc7BqKS+t0LL6xH+Q3zhd8aPiQcPL
kOhUrHucFF3NMhBIBFvmCvoyc8wo4yBZxNYz3uAxSqmUMJr+wNMbNphTXELj584h0oIyZ+KD3HjI
3ELpCt3OrykqlZy4KcvWdAC6ysXDQAQ00zHptptNOHt+y9B3yVKnWpNjVZiIzMprj9NegsTwdU5F
FP9Q+ivSMrZfTLHE6ij8ptnLWvFBBSGk8qlt3utRIgamY2XM/qpd+dbuHjCXy9ukkkL3OJEyB5sH
0pqTyhlumJ07YYWHTyK3Prlx2kglRNgSKXD92CoIa45pYRsIkj8teyO676MUuRerkijFvDJMuTCg
MxtaAk2gPvCHrrLA5YG9s/H5/Ob2xEzs6ji++0LrjrnhexsgGkjxL4SMD/rbIUe2yqkl2BPNz7XB
tc5chvR6jL5CSoiEOxrts903AofJ9x93n9PEro7pRqQzPMtYTrFMrBIpUmztU9qEtzQLWRZxMOvI
DdMvXzkRgHK5edKqG2xRpgN9P+bS2H38HLa+g0PIztAZ4WAPi7MhD7IAHI1PZWjREpEuoDIpOaQ5
EEvi0fnOL+NyHakPO808M12vawF+iCz8CKBtgdB7uWZp2fVOgyl0kq5+aCOjyMNh4GNql94fm5qs
BWJWRIxgkfWCdFZk3yNRRhwQ/tQ8jKOVPtoSjFlzQ2LZgVLLPXFUq1gTQf1hXnKtLUpzL6AeeXeS
ngeSz0swWmW6h799ZSE7GcJjDPIPovfkK719Yp3lQTS7Abxfeo4RmD3dt0U+eFZSXGRD8WRDjnNg
DI1iwXxx4nxh9kC8RrFIbDWXd9fkn1vxRDfZ2mA6CK6NWHgrC0O7biSJVrQJ3WBF9iwMseCw1Jer
Z5TbXrV+R/euAQyT2Sc63+LNHhu9+y/n0rhBFqkEpXo35ZrJUNfVv8/dbnBQoQwv3/pHGzUlTokN
l4d/QbJjzOHiRHSaugYucuJ3vYMNEUMLb+SGV1E5l61KnXgEGfZbO5dvkRADV5pAlDxpCZYi3JqI
uQExx1CYuWpGGBaXjGm6VnqOUCOV8NfBQunouOpVpTUBe9+GK6jF6Fh15dvKUffcOACSfCu90vtn
00nU25BUSQn2lewk/FANmKqvweine0atmGD8QgUN5egN9gj7+Mgw+mDMa3qSvELIFC6ShstvvIQH
gaiygbg4BNSqLkFJPa4rDinsi1tnyPuWkzJEZGKazIYgUn7dOP/FyakREmeE5h3/9nIMrc6gr1Es
gseGj7WnBAl1TlOEVSH+WbRuRPztJnosN+kAyU8sv4hr5vGODzlctIc9gLKKqtgdiM1mUdhWlUhV
xPOGu1RN+38PftumOJRX3raMXe9+eVDOSUMDpRwz5ij+p5BMj67UlDgYX06STiV3uBQ1lMcIHcpS
RjfJ5bPZnH0zmJv35Tr0JWTgtJUuz7bLPFDG+Qo+wAF+a3fCO9KJs3t5SdpplR9f/As0Yv+ftUEj
MqIzFSO31VkWSYlop+rm81nz3zSkSJWI3pLugW0Xtv9KTpaFBjB2zivyHDF1IdJE48t7BCfB+6b8
OoE0mKhZ3HEzxU+qmSp0hXqgh4mGUnewoQ5rwgD+HYU7WWb1oecpQxecuygsofrJUInctIm31qe8
81oxkRuaxvOjvu9Fokp8shUSxTPTBi9TVOZZqiU7wP+6P7Zd+gU5gqI4/+bmd4cDd7wydGZQIquY
rei8SJccDrqY9RpHJD4JVQV7Nd8d1f5VFBU/IeJib4V+GCj6nKRmhBDoNGRozAOOVkqVm5fhcFSp
XWvil+De5/u8ja/Xb03Z5Zu5b9syrw5bpGDJjItgek2EC4pOLbtzPyiCm873FZpBlhvVIQGzQjEZ
vLl+ordabAADgHF0hoZBvM5gsQAKaFsaceZVsxAnIyn82JVjJ1LKmJcdyECEOX8qS8XfwRykivEU
zGIcqyGDFhxARSeu95ekhsNG6/+yvZmllpJwfKKoLq78AWTR4BQ6mbZGxZiVYp+Uj6gO7G1Ag6Db
2s9rZXQQ7wbwm4yJLwtgcRVNvfTkr85u6oZyeq5Gzk1NNzBiQqtuW0TyUbQSA+bHKjO65efPDBjE
NXJGuINezBdMoLb5wBgOPnAAMrUO3aP7UVBZdm8eZfGU3kUWQuGL/Q95Joh61mFvZEepHBioLxIn
YEkTVeqZYtG5laLMrelVTRrgCVgKKkI3cTz52k4ph6cbwMLk6+b8NYDoRNLOBKRyv/sOLtru6KzH
eBmth/9ZZL2lpuQd9AT3DtBr9xIEDs3WMzQuH3zlMcnpd3E7z0E3BmFJo5oCiDFeJXxLvurd7VAT
yItCjSeidK4i9Bf1CdNKqcu+CT+GsK0zNTejJJky1DGNaCiiG78nhE0ho0mMVhsqTMVHguc5Fsic
3aPHfTmuroPKwW97gwm6r+k2FsTjA/9rIKSjNRdPCZiZbybjTfT36toZTYpJ1LfIKLLqGeEjKYAt
S4bBDi+8u36NOJQjPyTJtrMBNkQxCOOkfKzZ6Vcjpr38VGahPdvki38jMiCU41fsMon5nA/x1RkW
fUYIbT+J/7KzFA4wzsyVGKAmdI3VkqGYy5oCB+r4feuOWXjZ8LA6TwaaTF52adR7bm0cglCugr2g
I3ZZEh2sUghWMKvNr9IdMMkAHtm8zAEgMjkj64jft59Cfhpvctv1zLyZUp7NGgvh/zKucJzC2ePy
sDUJ5ZQoBkHTZRUfhW2Y9CaoDRGoDCX96AzyPkbXl00MeHSPU9s098bZjKqegg9x68wy4Hd2RNc9
zj6cscZNOc1wSERhzuQM3+SVq4+ofJIWa3dInAIxCl6by0HgRdJIrpNAf3eu5PpQt27aMIeEHRV3
qILu+6peW4WRQUPfOzlD02J5wWnRwdIQAYnNlS1eHQBGC02wktxkHNkefPqpmh9Ysxi1QdZyGhmI
FPXCyovWERRGR3Jq6PUHHYNoB33JAJOAQG+jyWBMgM6NfGlOVen9uV9fctPqaJNwKqvpEpV+dGjK
4ribVeHmJLSImfF4q7+eYUiHlVcdEmQqjeh8PwLE/TCaRCozi8s353tnuEYQujirS1t3BQY9c9C4
27xhN60Zk7zcMpBWTnyy3NeLhLHCORrNkCnWMOSenZirsnB4eO4lZnrm9NwfN/1yrOmzkqU0eP9W
PgaLyv5h2hyRNVEP2OhW+y1sNW+rVzFFl04FBaYGAQRsuUV2W5OZRrc0120YpqTiJT7XeCobBLUs
V1mAZoZsj2K/hNWSAyTm7QmLOdxjg+06oRC1dAmL9pMv/u/H48WVfpdwuaMk6hZh7IW0goS+tPok
iu2iGHOniPIHeZCg/WwfkEq59OUgzY0rhucDUf4e/2KdbeAg2q9Wj2ZVHQyPwlPOyWQqZbVbFQcw
IVAybQcWm78v9/h6ixfW0fal3H5ruWeOo7oxEOTMfbroaC7PIgGjHQot3aqxQKUc8qK2mGKleoF6
EP8xjibmgqxYFhj53CJkyByt38JCZMX/G1fhuDTPZ5GIJUermn9B1zU9sUZum23D9YTprSwcUfmA
jsMMmxkXszbhE1jHRMw/XUX7EzSnrwhrVJ8QoUbFkXBZAYHNcFZM8xCSjfrddg9KvPrdbXmfJ4G/
g2z7kAHW6wuoN+O7B1B9kScTlbmezhGlc/c9FNEeYk3Vm4o02Cn7kkT8yhgTAK7/kOvXkexQpuMt
cSRgxS59y4I18EZFGwyHzblDs94SQq2XGAzS3VGaBCCfzYSmMvjgrkedQtp8PpiHNJxICDXfa4bU
5eTxIhAm3Z8kihulilkxCQwXQ4Dsx60cuK8YTlAU70aPdmx+nHXxOX9Ydx+CVXliZ1GZLA+rxDAj
6YyKVOGSj7BU5gUXSqFA+/8WbGa/UqgAMoaHO7MnL5T9WjgpfBXLfqFjarufLEA68fVW/xzjCGEV
cCIT30/h3A46VD8ifHpZBVvwaeZQBHoCeZJHA+PaFFwmCBiKyuXbqQ5/zZXEBBu+9JjWMUCWuXf5
aiuP/AJeagd4frTxt6nUMsBvyWDfk0RpXNVwcMnFvSIVUxKta1+0D+PWh39Zc6ydVkvqMFzr8EMp
H30VdYar2UfQQe825Eiw/+WEwxs5JmQ2X1STIz7KHwCkvyACOlCL6VaBwH812+Xt+pHobSAYjklV
VpYzYazD+CF2C0sVbzsBgxNchmdQgDlaBZDBXj1hRh4DHstTeGgsK31cY+BQyKtDjyc0/PgK1zW+
PqrwtjpUdHpU/nPjju3Z9CvKREj64UT5nP8ZieDuhxHE3HJHgtzsaCkulz0jqrgV6uA2BralmOX+
kBJ2NV3UFrcRFs95idjzhR+OMWjm42cZGJ5Z2M5Dhb78LFD+1QgLJchXC61IT1y6f6lzNXC31jLs
FfuVuPbZznfCySQc6uo2aBxN8xGaCqsxPmIkAFqcJ5VpsbdNdTx1PdrbsrZbOJeIiks0jwsCFwb9
NdpcPp+fpGk1M5HtgMToncMeRBMZ/IHUnmvNRlkF4jbwnMJ/BkR2apER8eHItqKN2bqpH43a6Wvi
A+dCNLUK//kBgT6MQKgpXeuvCcOqIC9yekE9owGTZt51fFHqNnjOt1B6DngCxizfOw+KnqAFemHR
4qhczzUckOkp0y0VQUnzHQ0PIANew/6TbWsALsXAcSiQtAKDtfvNpcUrK3WUZCAy7r5u6ohIFQlu
sTioAVAO/Q4DocLyBbdEEwVUPPLhHOrTSh9+VupRa+LpA4J5fuuCeyGgDsjE2uaCD1LUP9qnL8Gn
6SO/gzioziVW4KHWA1zQceyR9N6Bh4Oa+5LoOnlzlnpEfoV8oH0DDmqgy7hM3tnD3M1nAjH/IetI
9++/aMTJfP707Bgly7OGBvJwWtrVMNadGxjgxU6capldiXQwLP0/AJAq1oZy0bL4JOf75+RtSXYH
KttC2plG3tUkbqSk5QQ5R8QBfYrxNtIwqXFoodcnx9OCx9i9g2GH8AOi3az4b7Kj1EIrdFDDcdWq
QhVH995UbF1YmOVcRyf0xkzsXwYey3EcKoEsJeaMkLIv03fs2XIq2eAtAZJPzIX3QBYiuXHb+F1T
nfhxvmSnBeFKXt4WrkEMDeADj3dLkuZOviCyemxQS08xF04S04rOz0diYiW+XuqlS5PNw1/KVdkR
yN5s16x2A2aWj/JiNTGI5OP9vHLxDKvIJdygMigSigsitOdsriWGClcbqDduCsKAlhyEKSUUziM1
ME0uC+tagDU2UgUcsfljFrfR6rUTdPjMTC4atPJerxXLYXGHUUIXOdEbUT+GeV1VhQCaK1zS5jhb
GDPTv9RZayUUsVESBBM+Zb6a6wgvnGdd9cpLC9oNMZAMQWFgYkeWlP2pcMD9J4uQnqRETQRqJvg1
J4e/Qr6lvZn837puBPGLINPo0TTO93Bdsp+r8JTsEan7bIa0bt3ERrP/8OzO46yJnxC3Fso3HlNK
oeoZ7y5Kc54TMhSINY/4KTqhiIDyAwhmhBhPM/7h6zS+s1sAGFkmTHV8CQ7XkpROuDNR+eQh9oEP
RawSJNn3gNB2QiqBoVzqpzlOLMfqXom/8eP6O419rsDE+YtAIU7KoWVMuOr7yU1agTHVfEeY76Xk
EqVbtIe15ZznnIp82mz74ZWDeNGcUha4NnEUJEJ/zVoymqZMsczu5qgDdd044c8vHNzeUMyGgicr
TErU4AuXqH2OUcUBa591zVcQhpUEKMLhSBRlKikiMpJmbcEU01QaMBsGqAGVay7u85ZQW3a8fKO4
oa+h1q92esVGucBeRMOj4oEsaPgPX1v7K4yCfefv0CBHKsq32FmLxTxOXPXLEiVwPwxmmgnnqj9d
AILFJGXd0a8g5aYx7/GtjFBs4Ndgyhs8Gfrb2fpL3kDTLltll6UsCtzyNZ+cLVVctNpxtf1MPww2
jdh8+pZAayvm40TAlQ+T2NVfEIBEEKlqE+/Xqh76xG7F62DpMFJelJH+Xw8XH3CzC71rXnzfEDLF
gDyYhpnrhv3et0JhdTuXOPKp3iKVjn3iTnmZTBGnYpkY7zb6tnBn5j/XfhGP0JUrHgzlrbqzkH0w
lUsjZOfyqmu2mqjPrEqRGyowwqR/5aezfwBpZ5FelrJ6+0GRBEQvFS1TYwO9uYgLT4+XWkYDIHZc
l/OwqJ6Ur7gRERDsfMSs8jZM8ZR15aFdaSFIU26eClBtrNdf1zW5ppkW7DbQG5FIDBUdzg4FMjR3
4F93IaXyljCCSMb2EbVBHIZMJ5gAF8D8FaPmrZuruoYTkmi16pjNsQs1amm2aoS2diHr0aWuWQlD
UItedrB03zUfXpl6luZ9BcVe/SLgXcF63A1un+VJzhmMMAiqMbJ9RYPLWUlPLKb8oIAyc0h70HFw
KJt5H4mNWdtFMzVFd9JQznj7d6GoRYWndPDTnTrOM/PH/vu13pEKPL/fff2EUSrMYhr5zXNJpf23
AQJHp45wjiT0nuZm4UXocdYo7YFSPXtwDsu9rbYL3cdbrqb+9CW7qsDTx4lkWfTlNvdPAmqXApuB
b64O4D+nBassKnNp2G0Xo5FeCjx4T0rlSS+Pxp1HbQiy0LMJ0JZ4uu5si9Th29/DVFKhRTa7MZq5
DDW2vH73vJoSQm3GADMNA3g/gMk94VN1f9kd5fM63ftbKY14Grcmfrrlxjz4qjuoAgwxGcfiX359
gdJhNM6W9gFpUHsoWoQKw1On+pejPKNAAfnF1+aXgI5NebWUnYFBV0a071vp+xjx7ttxqQZMuvid
iUDOOIE6EusK5QR0EEkON2SCivtd+BzcaE4oCDW7EII6/edc6LCTK5HxEaQ9rHz8/dEm+8/C9mn8
WQ3T7ORNW42okRDQkrii5qUR5aq4ror7eO/7ssi8eNv8jF3DEjUrYbCX36c1AGuVMa5T9SEr50tZ
7HhAduJ1IGsJKKnP1a/vQP4Ier6uRbro2ChX/aCiqYqQsU6PkAR73FdYS/AipUbWqP3qpyQuwHBy
oEWi5tikSLuFN3FZIBv3jf6kiH3vyL7ESgSLXTMThxjchL6VN5fDpE25wTGaKS16WdmSxVc5w3aS
Gd5rjLuuJzDDFZptIqGg48fzEM7v9DneePLYCKL3Q+or3ycBZVmJYpIZW79Va9vAi94DSfgyu5I+
siDmSt9IcGF78v9GknADe7hZ4WE4LMr47KImfbFI6qN0XhkuFbn7p5eCq1FN9ATIWcYuTrCX/n6M
Ws3sRIqlubnB/IO0xaqKZQnnYMg6T5LDWrtDgZCh6rXx69hET573fQ5BKNlmNuzp4xKHb5twI2eV
S9OTRJUbwLqGqL2Lz5RNm9og7uqXOXIyola4JTuZNDPjlpE296WipHTEkeicMhRcSAFI/oPWpfik
X++NBAX3uIrEUy1QcWPRkzDWOzp/qqKufnHLzxNP+NvVjK3u1dgNn1IC5CkA7hCIc9qQsKaEx4wZ
qYhO7y9x9Gcgasv8+ooM1a1inryDQUVMuICSqq9B6ZcDa3QPox3Chdxl2l6VxWtZs5IE3k3l9xxV
vMLsjWeNuZL0fELzdnagTWdkeTrITrkoiFtc+aQja5TYVvMJXs1v5TPUhhxiXpyUHWJs75m4vJw+
OhCd8ezHiTdo1LAkpG3KKhgeuBcYmFWU7bDEGbB4ri6Bc3ifCCbU+L5NHQn7g/8Z/5CYIi3SGRB5
ZvK3FEJ5T1lNRVVMZy97DmuFbv131emBefeDWI2rGJkOsXNZWum10oVwbpjKWaCaYqplU9uHlyd4
Ob/OrLMxEs5No7F2BebHGyemZO95uEX/FAwgXy+2zkUq9/A4w+eKqdNGpUARLKAO0nmNhEa0X7Ka
E1MuByJkygm3paGKxKj069bVyvWF7tDYR3ax//Xf6z1oFYRsWiK/9t6lvR5maP3XgU4fB1eULOsV
mXvfgwF7TLMYxm5uCbTiuNF61AipbO8WXMNZgi7Yex6oIa6AXEjd0PyxYiWn5hPyqBXoGEiAEZFT
jNK3zUpvW3LUUanMCDrVcx4bJ3Q4fKca8d2oA0dAlilYsXvBr0iZIkPZz8AHWFxIcxyVk0meuUJI
hqokTBr1vr3sA2ZCrarb/N710gYgHFN/7QDr68gWnj+PuSd40ET4yhpyuTz9BtZrzK9zP+DSzFt/
/0oSd+03NT8IvcEhNiGXwWf8FbsQoLd28YWzpcjaxJ6pQoY63h7zku30/EOBZvFYuK5MyNPEhO+2
r+B1Wv2vg120FKVi2SXq+tMWhntVIL+PzwGSdsD7TcfB4rrp0OgRqII3Vgnfy0ctuXovTJ16M22w
pri4JEbdM0TU+Uim6sPSTICRm8Iwf9L/xpeuFVs19bv143Ju+sSQPSIAMhvKjstdOyyRTUg4kz/l
Pe5ezbupj3ouVlazTOuI4+y1BT2k3EqP7P5Pm912gUntrDwpFza4b+gmv5jknkXu1kZve+8mxpYv
l8mRBUTJ/5yMez4jh4nrfcf/mYnVO7UXhYG6y5D/2Yp4Gredl1Fzg3KPKMisjZ1uE0dx+WjCa7DJ
eE2zb6Ng7z0HfqetYcX7st0faFI8ZczR12mKEGgHDNT42g5NPneGXO8Ot7tRg/Ht0bKe1EmpYfGb
WqwfSvKEufDXhZYniiI2vjw7hu5fl8fa7Banru4ejwe0QTqnTU7vrlLWuK+J9tu8F3aN8ohbV/i8
MwKEGeNQ4VQhyk+zCLjJ8o4+rSIIbjggUJJKj4QyfcX6MOPbBiuaA68PIVEJbkHNj9rKLyc7SsQi
nXOyxXFWqSotKyM6prAn0dOgQ9ZiYXObuPS1wY+w+HywhO8jDNsvjztoDC4P0reLOREENZdaETrE
370MmOHBZe81ngow+xas3NP1AkSuIkJtBfpUqQJ4u2qVJmzv6TMs94AaJuYqNm07dOI7U1gKn6qw
y/IArhUL0Uaya+AQ+iX3G2+jWol+1rakLtS71xrdgMqVLrf3bkCR0ZFVXxi9fF3SQlredt5xAoH0
5SFjQtoARMOjocMNIeaaJ+zI0Ug37ID55RgUaaN4A7lSOg04VEdOhHUlnmAzIOnu1xx6MWpXgcQ/
7CPYu0US1XPm1Oi7CLdNPsZwG9fZcYE9SNUSqFZ5cjhg8QJvbCsQO8iM11S/qhbOft6eCQUvM9yn
Fq+ZC3O7Ml+o5A4pAXU1uLcPrwiKx2SG579FRhwCtT6jd8BNh6IuaB/HNQbNGba/bn7QgbULNxwq
DDVGkEGNbXCEPdTFzf232cFggrKXdeNNOEsp/A==
`pragma protect end_protected
