`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrM41f83zxdpq7B9Bxc+63s/ThO5
lR4ebiIUudrMSnsXzTRn4negwrrB4VipTwcqyfoZbX2gIf3gPwkP3q41DFrLyf9opSDFSsyylvuq
0tfuxhMWxI0KvORiuv+DLG15sEi9Zilc4jLqmJBgxaj93813ixDm3VBlIU1BQYAYzQ6XobruGhlp
W7l+H9tAQt0BvNuSDNd6KHRHtkpbBcXPwpTyZJ7RstTWqPbVIiCntrKr2mKrXFSxquvkPLZLq2tJ
HYUQSXagRZkQn71RvCHiKPsBHgpDhs1lYN9cIncR6Tc//qtAqb+PfX/OSaluCOW64Z++1c0Ko44Y
FMx1QSIQbLeUjIM4+0SHrBLXvS8Yc3JN4pTIc7kIiDprvnG+wDYT2+lQ637BOQV06DruFF4SC5pf
sLXqjj7TbChmrB/O2AZRMhW2i8WMmJOhJGWeX5qy/DPdwFi5AT5N5SU5ZH+WuAZM1xt+1s+E6WIR
wMJsh0UgitcG4jfRsrbeA5dkQ+CE+f+rIjCHaAxTqTuh2fGcMJdqVcaSj8r0/DgWWJdsY9+FZ+Fm
D/WHwTTOn5TdQAzGbxNdWWCzTpfxRNINCA+2M7UiXzSkNK6sk3qOU7E+cB8loLYEB4bntfrL1wyv
2IywDX2BQBCpLrj2mcH3c/RMkswGlRtLZLeTKCJrTtLejEny/cN41KNaFET1FLeNp1Vk/fioHFID
yX/EF0eDmSvugfdE8lJ75LudUMDN2Huvnp87jwC+c6ePjS8iI/z7rpwsvw8VIApwKynlELyS7kzF
mkx8AwoDGqzXr5d1WP3eUxLE+NYnd2+svtb0lYf9TIYCuX2C9VfAFpB6Sl3iYSsk/agb6MmsT2VP
zgG+Fx5OII6B9hPA0snh7UmmBOyHKWo32QX/hasJUUVowVJEeq1R5fHYuX2H1Rz32qBRQ3wDap+m
y4kpQaWFlj6Dnf8pBPZiNUQy2J3W/9lsF0xz1KyzNcXdZ3yjRLnItcbk0jfeHOyb0ZD0Ua0Q3yq+
HT29eInAs6M46WA10lpu2rlNUgGmQwpYVY+tOaN/q6qH01zyftzGAfYKvEgAkavXO2oQZ0pEngFh
trEnV4EY6u38bYbbV0o7hBqyt7Zz3y8HlcNtCCcKezkwyiMAtDyC0P4q5LOk6XFeQ5xSCM0XyVdq
+QUKp9ZL6kfACyPquqYl91XY2dt50STwnLJ9g9dXbbTTgRsLNNkYd9K+/Fg7WQs4Bh/1xKo4iwYC
Fxun5UnVXOZW2tKlAOHnPlh9VjFFF3CZW+o3yrR8LLQii+GawsxbXL8gxSx6I2E0bqUmVfOYB0Fc
hdNoYiRtVZC2awSP/nB15QtmcbzpEfxa1cXiuh0E4FE3jpCyrQRsq/1pyJv6dWpHjXzBK1WOdqEV
Ofu2YbO8C7MeD3gTPewo5mZ7hIAWrmTMU+RGv9+DYtTmb91glYMKVEQQ7wtPhgDPERg+/tp+bBtB
hKyEar8C09Ew9kpwbu2IvKvUoT4VFliEMrKuMKw7aLczBIR4VeGBjCfOqnOBMjzMuCnRgtFLbF5p
U+PHaM6zybQtzn0Cx32IoK6b0z40R7U0G2gJ06gSDu47mJTyPAL5qJUwuRTk7s084HVWCxcaC2Cb
03r05nYCm020YGX8iiaAl1ua6IrocqWbEF4PiPnd6VQXsCwCo69/TR5XO4t3syMXWtXJGLspyJ+Y
g2tXsHAHI00/JS/bTuCG1PSgkYiZXPSweQyER8bdS6vIj3mCdJoe816F2cSvb7D2m/UAsm3tWR4G
fXyeI0L/RG7CmmYn65z+fnubeyqSki6fe5HeUkEBXXtscbHYD40+BQvgRA21N23BNtZyrZgl3CNI
ItfWr/+XkbqWeojhOQXANVJd1lsrX2v60U9Q9x6kjm6RE5ScKtx5bpltdoP3jFMefdeqh7LiQ7dy
vcPODc+fiVpfodUGwAnTrS5uW56+EKsPgqpr5OrbuHGjlnoQdUmkEUJikNM5dB7KU/4zZyCJeSos
wb4uUnJZUsp3Vq6tnz7mbBfYDTn8eNiXZHswppdijcsd4IIR74gz3M74FxKbH7c3t6m/R/wVkhDq
jkbdwtFraoilXP7gsjQ6OmUGBf1rW3VIwwVr8xOv13MdmN8Ak8JPAG9cKR3oMvaGfyXJSIeSRRPw
HitiI3B9U8XvaWDdiWOYq7VPqdTEb65EC2NrKg1sc5kpyOfkJE4QJaHiVhe6elZ4nQIA5HfYJnJ4
11CtPJ7K7EsziKnEfnuzvObg6wARo1+X4R9DCno2kmhAQkEWajm8jeTb4K6DX6vWtUUt4qOfVcsv
04GySTV5tx8hY9xF+o5kpSdR0xOPsLztIk5voglUJuo6mGIO6MluF0w8g77AW1ck6TWcV+88jkFc
o1OLLas/O5Lu9rRnoa/zfcFRCVihWqX/aOLu3zK/gipKQnhjWqHZvTTcvt39UtHFK8uA9YgqxQYd
Ygpwvu7w6OGwTq74QyK2v+ckmzKh2ogbTcl4gzA1kccRA/KdKycVz3mawtPkvufcZ5Su6KxeXKEq
gBNHF+U09cICNvhoIa2/oJKRG88pJegUyGuIek4Bvbm8yUoCHiYWvtlGbeJgiHYRsPdrzVlYlJnV
0E4dHA6wpcIwLpk1tBpksDdysGlBpKrwxod+Xh6h0wRHcscn7E2LM099m0hIG3y/qLjd4irHW5/D
lK8UsQ26LSgILsRgkr1mZDuHrdd/9qmvkHSCuUuZLJzrmoXNGYKfPKwD8PDE7IK4mz/xCovs1xO3
hpeSDPRQTiEoSK4WT+tmC/6UAjq+EYQYiL5LUdE8gKVrRu2F1Y4tcYD6g7g8g8mLTblJ+CWnAzUW
Dvqz9UfVw8c0capJ+AEZ4R6urm+Zavnxc7VTsXeIWnWrKKyF4lCOTlRRtMllgyqK/5NsxLIRuUyu
TBfMNjah7F/C85vaYn4MTIY9lMhOyrl5+qkPV+coQzn6TXjERCynaavh7un+/xmYcamEdjJTz4NS
wmkvSbgjloePuk9t5R/+CiHKOJK17nLOMma0v12RUUw4Js93fbAmth/QxJwdlAd6FGI/mcLr6Woc
mPO3cckXnc3NAUkZpUkSp4kN4O9QsE3bwuNAG+l9HYPPf82+goR70Q05RiwMW4ap82ngcpVgatSK
0hgP8U7whfbZe0OWDUAYOcMI7yHl/5DQ2bp22NjaeDWACzZLsmrAiiN7HSBubkEg+M84hdH/ODEV
FQAjgfDHes8D8ugKS3PZcAYl5xTmp8ib/iChdlYwnAH/XR/EjOD6iBXH6Hh5LJdUpHUBe8KFLiM7
R86JS2OXbF58PK9Yx/Spwqh8d8YL7HqR/UZlLcZU8nSYEGRBGjfbwqx2n8+ISx6Nua4FD19EFHv3
Pe7mR8zmAz8IgiqV7xKdM9KqfcGKclPf0CCGbcoOguSGlBxGwVamYYCdrNFen+hDu00sc7iBmsPc
v+ZvhTzozpzgB6XRrceAnLi2c5hRTWJIvwop8AGlMa2DC7s0QFAn0/B8yzrHMmcm7BUHF9MCpgsM
Clcm88smoBYKxCxLKBj7mLEY486EKQj6vsNJ5DhFS2wO1CkVOcMRh55P3J+L6yZioDO5vLDkT+F4
wKSgFuBRN9t52Ordh2hxeBBMoPMdvMZrE0LqYz9U890rHfj7k0GFjsLz0HJBX7iHclT4lD1sZ3Lv
qHeBu33ZU13MG4yXAnIwlT48IeheA9HK8Gc3nIhL7EKQ40ExnzmoYunFbZXMQ82iWJsgzhcTaKni
gLYaK4yUT2T6li17cFv4Kcmd5/3UFVOQzKi1yBVcLjA6rFf875BbZWxC/ctSHCGo1CET7U9nwdQD
gRfMGGVR5yR9Vm1q1EHBVpX+1iAPwiC60G31mDCweg+YA/Ph3W5grl/JXuVIc+1cYnIGkOUv3zUV
45rVVwtYEEACrgVz4EelbUkRdwQ47/y2/v8MXRboavG4/syUPPzoSXK2tqbzWQRMs0QVBPDTGwiw
Kka1dFIubkCKISWi6hhWK19I9amcLHX/Pp4whj4wkw1aiPXz+gv896qBReV9cqP0Xug06qMpwLeN
WIAr20ZksJz7brtMH8eTZKnR8jxDu2UVrYsel+6FTUC3hcM84frssN/NM/UxL7TqZzRI5LPeJdtC
1xen3643U8NT96E87xMWxPzsj0t4GVioH6CBU1YkfSXka4vlsKEs9NIDPnN/ZUPFzwwIvYAxCHWD
SU3uDVjfqt0ZdT1gndnNhlIkiujTayjspYZXTpzkbEGUcXbfXLmTuNq3YNvzz7r07vPEaYuK737v
OPeEeyp1R8i0k4+A1FG9s30BVx3sslulMjMvPBHG66AP2K7pTQyFQG3RlAPbQbh3X9DAS7vXhWnm
cRUXmJV2z0uXOuf0M/Wrg2l1/0H0Zula19t9gvrYSyvye/c7AW7GPyNDjCNWr0XDna1+bg14jTI2
GT4HB79NY8wDv0cGh8Zffe1i0Hjd2Fhqq/v7NCV0iTov1JD2n285xyr3oSD1jFDx7KwalLCzkX7L
q7XA1RqpLOlCJxEK9ysvibqibpTB4fx+za5JOJZBDtKzZ0tB3LG96H/nCswh6MQUVTLENIMqtsSn
6neEmCWCM6HUYBcBDP+hlccl7Vzwi/ri+tjCUogudkGdihmWuxXV+jwPXfn50irvnwfwbF7ZKIv0
de6jy6hmY91D47jOoRo9MOWBQMYNHuHot3B2O4I59N+XqEhSTkXjal9Zjf71/6OpdIzwFQbJK1dJ
gKVxyFN1hOhCH/LyTRLuNnI1Ivf7Kze2324M2O+c6hZ+cuPli74uXBtftN1DVNUGbo+noBwQ3ddP
G2o6ZPdNmLA0iE4f89oRal+PNtHjR9GDz/kQH+/a7XI6e8u+dt3wVC1PD0dVonipIJnZQyzYWeSV
IxfJTzihNr7+P8W9QZjSf8pMVtSj7qfrapfyXmvKIBQvHSSv0Qq0xJt9cc/C29c537hFU3PREI/v
Zg/WbQlI18OKs4VR/PKReoEhLwo5eH7FhPsq/lf3dV9UeytQU8DVi1dhG1ymGdFgNo5WdTEI581f
3++kqc1xG25WDErM7gbDGPIR0UPgzgZF5Mtm7ATN4/VH/ym0iGOzu595vJrTVi0MTb1yt+6V63gd
u/DYLTX2RaSooNqh2SWBVA484Xb2svap9gKBaiWZqSoINO/mC6/CJEuEYes2TRRDl+vXicebQoYj
jnxLOOnHWiQDeMMnoupDmlvm5NfKC8InzeZB8mb0Xa0+VKQ5hbSr1aqcnG4q7hyiQsZUdRsfteS2
AXt4a/5bx+aGXI9lz+wi3vlZsz+YWVFHwedlPLxENRmIBEtFBZBH/DCCxYm++JFgdN5cY+qg0Jek
uQKnwuEe+u3vkTy+3fc04/hakRzcp7Hy07P3PcVGp4T2pJLSHNOi4eX2Ln5F5YQ/b0GePhXCwnbK
jJdaeKHFMCplNkE6IFsRAe+POazpkYAJ26jTtVXoWlkeYsKUAKYjXJ45VzlBY2uXKeJBeV2gAtwX
mpFu241Ty14s5ePUQI6ooPgk9tUPeIaJWAsGxOvgbB8rwtBGKN5+s9Jurl8kf9r9cFM2Ht5FAGLO
JNUNkpXXViFPymmSuAcsMGktevDALrgmBTdrSZbNkoBSj5VxgwdOiZM36E/xPEcssa0ZFA2yXcLO
3HL+81OS9zsb0Qq5V//Y1VsIybKOgYrw2O4YFE4m72oWgXgzkWJ3JTGNtBipt+g964YOhjd41Moq
+EI4XQchuvoRlEWC7+aQLpOAgyx989CuNF/4TrI1lpowUR+qOj+aKEVldBvnxES8svKv+SRRcoRV
9tRFPrAw6LUOkr3fWpnkl4WzglDx6kXVbC33KKnaYpH95Xcqtr1BqhYtD3yHUSQbgOtHOqqJHHam
SRyQchaXpgS9jgmmicVu7jaPRE1GrzM4ged8DGboqF89slMlF3LaBmT3/wcC4Gm/Vy8yUAWar+z/
PnKFf+fj2jvUMji36mOWQCqWxDXufhpDyZDE61bFBcdDjkQ3ip4gWPanONSyQ0BTwmtsmy8wFGlg
MhNWzRYTcIXQS9ZQYXOFHkpfdmDY7jxN0O2grm6m6/R2Kx/GF6JiBDbeUdueiX/7t5lsXJuqyv0g
0Qh6r90MMoLvLZPTSA1Q8fzxVhXQTm1tZ6bJdsZxb7EK37N4louAsCKi0D+criHFrDjNyGuAZj2Q
HQCY5uaNsLadqzd82FTI+E61agVoHsbjkqNBniurIW9ddcyoZDyF6lmz4levdHhNxFKCB7FW14kA
/27HFGgEijKXlqu97nYBj6T0Rb/3WXc+lH27YQqwgKQloeFxj77Ir27TOchnxoKcZkvu8fhwzW74
NC0GBYdNdsID2HFVMcxZsGf/P6p4euCYzdExG+V3pMSckuikHats9droCo3IS67UBh4bT9X4QM02
VJYNIw0O9uI7n99S43anm4z19IeqqIuKeWVY9ndXksH4H3s4tRqD+KWzi6EuFuCx1fyoLLvr6uLx
lwU7GnoSuws5K5vHYp3zX4tL+zqOyz6Qx2s2VeMDAK0s0kOqIwmHkOkRW8lLQpwBrsYJsKa+ANq6
4S1GUWirXGYyuYZMlVn9TExsGnYx76twExuImJ+VjU91+at0eC09I70O57dL2k8PWhdJZey70RhY
3NL/pzWFzBwSl/umoOkr+cETbb/e4/ilw2gjy6C2wm13rHPsP+dcctkVeOmoqZais1Iku7zvzjT9
jRa7V11V2fjcY0/TbynkAr4nzI5LFHNrW/DUA5/OqM/5YuOD6EKVIgT/PR+Glbg9SNK67/aF7DJn
z0e0VUtSU5Cka4QPP0WzEDr5ItLWgsFoeeOD4bRoaLQoK0QaDQZPZKoyAYy7+X3GR+qnttZsMtqc
yqB1vV4tHalILUSd7PgFft5YINQLj+wny9g5e9vaYu6l7iJjZY4hYJtqzaN0KUgw4DtBTmZyT4eu
WYG++lGbcjF6CuG59HCZtvcoplyByw+jueHaW2LplBnPd1PFVZ5LYMC2IopvMjDHA4QauY+fTuZH
l64XPR4zl+PbPVrSWeJNSIPbudhESbzLiIBWJ3aGVRS45lhbvVJ1LyAOePpmqG9M7shFf207OdxT
m2dTXNDg9fEUGpLYYhmqfm6O8YoEtnAvZVU+Sr3PMrZ6FQv2SYWnA/pZrnmZyZ1KHNBvCXRMIoc9
2MwGjeS7s0CYkDUEgTkMeh+RanuRwkGSXoras8+IW3UXU4hSeXpG91t0goE7oQ90xtRktmNZRvk8
7dvaK5pnfzBcBYjYBUynvfK6Mft+R5LAZhzd2dyRkP5RnfU9bju+v9GRTawxzSwhbCFPqXz8Khbt
xYms5unXYyYHRts0eZi02F9A+WoC10WWtvN1qay+cJfvvMq13VLnFgop6GKMtM6t1F75FcoNu4Ue
aMPvaBM5gYD9StjPqLLOmLQRjQNe7VtwBMsdg4wDcFq2FYco0wiBQ3HvPof68WE1YeFxhh39WIpS
M5U/lxbBCMNLc5BU44Q2l+piAI9Y3i89sNxcZK07Uqty+eScDmRhxAX+4FQNIuTicSGResLvsnrb
QS0lngtp8xFhvEA36/Malp6/2oYCXc2I/qI7E6GixkxGHWXN1CrrnIuhbe4h/CxC8n8cnVXngrXQ
y0QnJnNjyChuirzvFcYTvdhqeKIaWogVvcHqLbNsrJHcKwvsg5nhuIbkAOKABDsz6AaAyBcwrAS0
uCJjkks2AKUcKS/Fz/wxDEBgZDcdcBX5yY1dgMZse/iAdbbWLj+Ky0L2hUAwzK5wcjcMuB6BDk6C
tabdSrO+xIB7+q38Xb2BpVtN+IJJAS+m06L8kKQ8QmzPnywfLkWnoyrV2dL6i5AKt5JPbAuei7Da
A8kQKro1qAnkWoHWWs+9VBHN2REupo1tHhuoqDJ5yIfs5F0Ybr/GiWf/M1Pd0qXQpr8V6uNbhyLi
b7jfSL2JqXlOUUZZDUx4EPeBAvxFkvI6q7kzD5iMhWU5wFUhBAOgqF0xv9wOb1ExC+6h/HCWkeut
SCy7ERvCO5E5hTspRCFPKZFcAA1VFCWaTGndnmw1SPeur/QTo8FiLy20SQrpcG0xDM6+xiRIko61
3FJzQY5OpAEz9KhnhEvgMRlpaObAZHZDSVTHJ9LjukCtYMj9V6cw/TMtTW8CEqqCWf+rPyprCEDc
hQRLzgilKt833Jps6eEz0pZC3Niv5tb46W33KTfmD469alIIJMDmI3I+CKgCdlhzsn8vIy5GqHwN
G3AIITjz9eWUp0YGOWbmIi++9FW00yKJJ13TzQQTCi1VvFgs9jCJ/Cx+JVXj5QhTDGlpgbrH6124
kqJNQ5gRSTtrGSgtmxOBYlw8ADTNRoM/xjF4xQCBtynqsoi6kTrmNoVTFYVNWA3XFTbIf8+igq4E
1DIN65NLyqjx9Liseg/w5bNKuxlPiTbPxuOprZP6Qab2QQzCNFgPeWhKxvHFiudkb8Oc18MRU4Uf
UJ7OZoAyTfpRe6umX6+ujczHKYVyywWUFPF31GKn/HGvfAw18AMv6czsm0hE6IsyjYnTd0eZ+zub
VSl2P5DjG3EvAcCfgtUXeBZh9jZ360TSncHzNKugoxvxujpdzQXjkQTExbmI1bmySFEV4y3MAx4M
WCGkzVddyWCJnbgWWu0L0HUbiaBKA2uNgkve+8PJy7qPz7y0xUqhGClRhmg/92VuDyNVnjeoNmNq
868oK0iQfFPJczSa2SpzVey2pqKLaXDdJHEi468Qim+vh5W3WUA4u7H5OK9Ege8soRm4hsuhrmPb
uRvX8RG8W//ql2LdeN78zygpA42AqigksxCtH1+5MXw3Q+Vtc2poNZywEMaxAGwzFt8p/yaIhmvT
tNrfmPd1WhUdQSEdJoB6FTj9kf1tWuLhyUZWr30zO/uQafKuqn91PuwyOsjOzOtly1VE18AFkRs1
obDWhm9FGoj20G7/ZKiHbY3oMuKnfKT2TIOUa/18mwgF8Ir7QL7MFCWhSJFxR3JQqC8usSuf46Rx
DzM0VRMOLHz4hlUjJFteZCx/B8SkDM/Vvdkre1/DNTi7L7A7Z6a5wjQEeILjRwNBCuY13odiLKim
xFd+dGCxZL1KTMZNrMHm3QDOLD2PV//JRTEV3oJgJOZN61HfR58RgwbFXoSBH843J+9/Z5uKmS/1
iAGE9eG9Ht9CGdOcp2CDVN4DBo2J6+A2E+U2tgT5Wk8S2+bulzT61Ewe/mVYUkvug6UQBHY48UIp
gEoGR4Pf7hPvjIssyFzBRhuXo2EhNBPvj892JN1dLeMFMDd1QbcoLFqysKz4BGwtLsgNMitgbE5N
ZicRglIVNmXWImH0dPu8dGBFPNDcbq02UVP/wcYHJxm6JGzEBgClumi1AmeW1gGjbmLijALddvJC
mE99I5mtCNeCtgNVvULjll1sduCDJ6TkM4TwIukcLTzj1K+qC7TIJtcDVBj6o+ZGvXcCxP9WV3+C
pxJ80EjakUcwjL58XamP3dn7kxJvF6TptFGBHfZLhVXEkiidhv0LnUIAfR8wGAwhfkrm6CTKXF29
q1VOjntSGSi76NCFzAccSurZheynbG7E2CE5PGdMLV60gB1mzDmI438bXeEh4o1e6gMLfaJbWeXu
pIN4+myDP+60vw50RJo3kn+NLUy57zbc9Ya7dyqm6wa9SdOeP6O5//bdqODO2iKeU9bVv1C5iox4
TnVPXlYgYWIZQoOCNxAXN7K+tEdSNkCMfbxyHaT+5o1oN947FS2eEWpRN8MgtPw2JRNbcgpLXMpU
yeFwDCCKv2cJ0Vz/7SpRrNlj12EJJgMnpzo7Jj9QX1jGwHV88F9k06w2BrY/tLMw2dyKtsDiqJp9
hgtzH9jZ/cr8kaDU3mq++M4KmRmSjRj5Fr1wVh91WWnXDEUUq16Jisvwd4RzGvNHKRhRA2NQXG4p
Dh19W+EaMil4DYTEuySLlksYFB14tXQbpSKSAH910NNK8z9+qbQdLBV9kT9dAIBHRBSGF92buQrK
jXvSflHe4DkVUiRbtPEBy9OrgZrLV2D2TNv40izlzQgB+FypXnvNrMqJd/7zYJzjglT9wLzNDIoW
kTR75dhF4pXZCwJ5cRBqy0PMhE97yY2PjYotBZeufxtTmpxh2OTljIRXW7w+XAm70KX/Fovnjm99
Zt+YD1YpK5huGngMCzMRshrkF7hPcsr1W2/AhrTxsH97hs8jdQoVjyXo8MR/jBfQ7kLZkraDu4mA
AUkJ7wPZfJNpNu3/H7TnwB+BwZbOQKfe68C5SvPdAD8cnmegbSjcAdU/fHdkUXkCYI5FYlZ2xjOC
yT+6SKVEfdk4tKNx2zXfEX2ZmlDiQJsRtf1lvzoWWR8Eekui2a2E2n+8SoX6lSyNyEmhhIsp2QPu
FUdp7kAol4Qa3TwHk0C/toHKbYv99qg+4dbJ72gfYSEgKKbdWlSIpJZroWYtafXeXN/brUQh6G96
ttLHnbVRAAU/zXRc7oCUAHSTz8ks/KkA7R9R+lGERBB1lt4cGkNWzKurD1Ggi7UN0HlEQ1qno8xs
XpS/sVY4a20dzu7ZWRxLgvpX8p71OXiBRQnLp5oY/QDWQ+iefxIoHdw2wgIVFpOiVl3UOVkIdDjJ
JBDsitXzF1mHtb9C/4QriC8d8BaZz/EM/l9YkrhscyfeN+AAVrHzU/aUcYbB7Q8NsECjetcMdm7m
SisvgLm88EWDi1EaQ5fjrEypm54sIDZ8dng2l/0sHEhIK0jWDOrzawsgTIZXKpB35/W3B2TWHzpe
ayGMAENptc52xy7G52Mwak/k4APk/I3JP9Wt9IfP+LDi+fqBq2Zsf2kO0flgMGD3LnO74/4ZAXN+
r9Qby0thP41UuXL9MjRXjjMmEyPF3gFExiASmqfYPo6fj0dzcK8IKKdUyQVMJMdrXnSmPhaB9XV9
40LY/9rmZ6zDM2X0LN7qte8yRoOJ7rLdvb8ihv6BZlhTsUzOa25iSMZljbsz7NvrMFYLq2JayeBe
XoX2EL8UsC4jcQHyz8qefXsM7eGXdpp8knfPaLOQ4Z20Cl32YptVoEfv7jzVebC5IFdLIQQmawka
719WOWAS9DJ9p4sUVzvYsMe16K9I95nBwUkSZ9C7D/Lc6TSFbKiqJRmO3ste+xIIyCvEEdLorqoU
WBqUoe2eKNY7tAE81xXkfyOQOqf+DCh/JqHcd7DPvPX4riSkPfGkawrGzEoJ3SOF8bK4Uqds+aI1
jJB++h8jSzEu/LZYwl6FZb0/5roAGyOYwU5zJp2pwyl3iF5QkhkVCeqtkJ5GuZFbHrihye2bSSb1
1zxke6LcviXsv3Leb3+aMJCezuiUQAsy7Bz7UtwhcvuuR2aiXg+EaIzh0XEdPrsKVqLxmMI3aPUy
jTNe3l6IAbeGGAJIwWS+dAj/d6dYZWskzqXB2AETEhxWv7h/rh9+xUeWusKGUxxDykljnsBMEzai
g2dADdtg27xCmld1mOJrrh8wogtK7eATvdNyUfLVs9CjPglynOROI14MOlyFh/Vy/X/vRxpcybDp
4n2sDKtIt0QKyRpH13iBdcS1188SB+H2eBT05Dm4yg3ttSZZfo+a7YuHoX4zIbk5nyx0eSCnwxx9
YmStV3mX8nJEeJV64YHdBNraEfNFEcpjakX+3WAKihXGvjvH+WGHDhJCGAaQiTyDX/CmpgjxDIa0
DT+D1guSQY/EqXd+ej1HC8PJvCA0dLfp0yM9PrKa+wuQl/Zlxnyko80S2yv7oxxh/3p/a3hlENau
nv6nbixxPsEqp5OclSZT3e9B1mDnhT2EDRnWCPFJOuhv07TL5/8r4pwEZaKwD4z8iVOTgQEN3dgd
BAeWkvZT9FHggQ0/AWp/jALKFHRNiCMzJYNWrFSL95eSQnxqVjkRRq4zWO0UB7f18RPT2tuIcZ6u
46XVg//dXhGEMaoP/eMfVRL0996woHDb73EQcpo+tBuOJB57Zpb928GHfV18AwV7+hUO8QsIJ7vU
wdIyM7v8FkBYsSyIaVdlRD4hgdzB0ZnQrUeBFFdEHVdOhqmmc1Da79LgxK7c4isYUpEU0wqlViVg
FaF8XsE/7+Gx6Y5A+LRdF3sQzhx5Cyusbf1nD+N8VlRyknvSlkJGx8KGSmF29Tvahc7bzG+Od5aq
wL72Ck2XEv33XTfn8kHmhNv5giyYcSgmnPiWGMAbVBZH0m9mBCzHiguKTj8f1tIHR1lQBji4iuDG
Zsl1qNVPlLeQG7wOK3iAn16hiNoR27smpe8GgQPvEH3NKxhbUqeooFzkNmyaHfUp99T66jjPEBJu
wULnfd10pxCYzvjYFip5T71tqs39Ts/agpmhKA3yVzjJnYeScZCpsOo16QUJzvatL4q7HNJyIb6f
rYs5ELYiUeLofVw+FFNFSG3iPmHL0jWplAZ0CDaBZLe2KP/aDEIyoBn/FBeU38c2n4XeoncvvrRD
cN2CunFlghiqw992zR2fkDpL4SEKj85fciawqWMNkJp2bmKUL0ReRHpFkMRxNUBLmB9qa+BJgS+D
+i8qTzABnvAtQ2SDBa/X9m+dDBy+ls6/HFv6igrX8rTksrqfw62LdGunkDmdltOmcjfqnYkxV7sC
LbrGePdYk2cNpxh/OCZwNLrFWGCzQ1RxyrLEzKj/pq22T7b1MEYTT/AWSNBow5BkQDMbYNBD58CH
N28coqS62rroBnQrxo446UyNre5sSkPplm1Peg0fID1vX+IOiycm0Jg4jgJ2hTN52tndjqLddX1s
txJNlB/uvkjdVhUWaEoyZJBOUrBiDu9jI3QhPquvOwBVxuCga2h5olGTu4hi3ijQVLdfLm6NlImC
rxR3gGwUfg24Gz+iEYgy68J8X4YS+VC3+HPyjsxGpMVT9eLKhyYlVy2/HXgLQ+hIxGhDvZmqaOye
cgRP4RlfJvni1PixZhrDLND0Z1rP4kx8XUtZYE02JbkOZl5UV42ZLI2YgYwh+OxZTDwLsHjxgx1z
+EH5yrmO+Vf27f0sTXUmBRc7TM9yp1lQDp8p5e8JgfvZIKXETNeC3Nx7XGBvNGGk3BQQIFGjH/ro
9aEbU9OA3u+yr7GCoB/k5d2xVmdY2/j9+jlAaePJJDUVYK3SuCdORD5IRcF6ef5QkOH3EVJ2ZfeI
UGQy9ksmPM5iQlon2DgBOOM7c5p1EOEVvjCpQMcCrPKZaH5LH/0A+0J/E39cp6nVLdPjoxtG2Ica
bJePofuxAutYhQ963zwjwOZtFheMo97d9XNTruLNXucyP2+hWYpQ6i2UnXf3uNQ/Hm/C57nLbHNV
xaIkcDfoXzzrAaG2QnhdhJfy9E29XiSxBQcJcLfngQje2kujnFhKXUlnjnajU6hYPy6Dj0ityGdR
xyRC+uklAoHT6D2lSzXgPYMANk04YAy7arZN84eqKrrNLAxEs8RMC3Onr/iXa25vnQFDQbLhCtLB
HATbqHKjgl5mAVIouEyCEYtVyhItRv4fXPULnaQH9fAnscinRbcAu3GWIoMPpXuMimPqhSF6viHn
IwE6xXUdFJKkT2x/r0mAgoVoLDgwcp/ap5r6Aj1b0EkhxDxHZRsB7ArBoccWAOXsZsWr5ETECm5L
TdOkxEgtILhcXCfNOD3J42IYsVGGMPN6fvj1DLJXdZpQTVaXKMzKYcguCm0Eaazg3AfYknuev6rJ
z8konSy4ucWzPKdKY/hsXOq2HALLVhms2bEQjfgNp18mzzMbqPqfaW+Xd9VJ8EnWkLf/q2oKK/Of
h3vNMmkm+QpA//p9BBv9S2fHbSKvSck0Uc00Oo5bkbUDZxeG7152jKv9SFk6504dXhZ/w+DylXiz
I1FKae94EFYrkQ4MJTCYM3OvU2pKLKM+NcE9pLPCvtlNsCYa/BpT81LF4l/rcSR8KvbHu7+9kulV
lhgTr/hPxs9FJxPE5ZGIP0N19EL63NOMM9R6fIF7bTOPQrUkbB5ZbJCgrE2NJiXX7BbQ0hs8n0od
FpdzQ+v/tjiXh0xEF7IEs9pJL3ykSwElmnvTRfAHK+YTMcvlhYo6khy/OTRkfKWLJzKaWVhcinjJ
8mF1Vp/3T9XMLa7y1LjM1ySkuabHpRfE1h3nkI8TnkohWb5qeSXYdfEBuYigq689VX2aexj2FE6Y
ppqm/TX+6MTbaTIYoLfqVoA+16zeX+fRRbzpNy6Q1Apw1d5BdCBctOboRcdJwgE2AglDxLqSCUGK
gHHMdelksIcNYuDkJqxtwzS4UPA5UIVnSUuaC5l/pxx+8du3SbUGcIHxHLcLyuDy/3wloMWosKE9
KtgTEcZLjC6vMTeh9HGVkEzhdJxJxBaDM2fgdd2dtDDnuRwu4u32UaLDNAJnKYau5P1NK3nXYmz/
kcadPpoRz/iyo6nNpmQB7CTEprQgzM5DYOwm7IvOyq32f1pS1TiBlS8Gc+ewTmokjq94hHa1HGYA
GVQLkPdgoS9zcCZ60jqUVlZg852mdnlaQdGP4savMUdckYPpy6HL0ScEzBWv70wDpRySK4h7rfkY
xRybzvIaiLlp/0+RIUp9XPzJxLLXiOmLvJgoLpGwuIS7LKDDGkr1GZMHJdebRv/TB1Y5eoF5hFhb
ol6uqmRAv/fJJFrQa1V0V1/OhXX5A/YxMW+aA+mAFSUcJAABy4RSwFEgXZJ4dDtBdoe3K222zFy3
wLJseUjMO8pSqE6me9JZfTr0we2v33u6mXm055n53LZYc8Ac6P3jG8le8UQLPjeVZv4QIOrvIyZQ
dd70tkt1VPaQ0tJUP+WQXzufziWBTHrH9RfSX7NXrlk9QRx0qv+vfauKbeLw5gd0B8vuzZThxjtp
jC0x7xhNj1YPfESkpx8jEaY0FBjFjnaaO7869g9U5rV4m92L+3F+c71bf6rUVyeLTSq2DXP3J7Yb
MSGZ+rIUogYW0M4W7y4dPB6qz4GEB5MSKLaExKYf3Cfs95+0M8J54Di7bjyQpHUGeN3swpMB7j0Z
vWPnJRJ3gKtRSJq49JsPbytqm0IjgqmxjBKhoxsNypZ8y8cjoulraHJ53oG8AYfldStg05dOadp1
lfGqM7uk35GWnKuPQWUiHKSdE+nM2aDCuBp2iOzE2B3eVfa3ugz+zOww+JRAkD3/DEXEQz7KZ4ap
1DyIQDrN/f1+G4j70Pve57aviNdvu6JAi1xp8JImITN/9owidpdcMYdX1fYMxwLVsAAFosxzmzqQ
PX0HQ91Y/zCny1Qd8BpS69w34IWWliog4790/c0J5Qr2z/x4bIL5B3DqoiDzT5N9+0P6RBZ1GDP7
QZ62IinvamUa1uAGS8PM8bi6zWZkEQNOqZyoPdWl9D/3xSHur5IY7ZzLRxGcsVkltpnTeYfDwKmX
wREhAFfoKcv/oX3akBfro0jRvjg64nd6mWikg9Jc0n3gZQL232ZcmWgzlA0ZhbxbboK1hOr6fpQs
OhcDLBK1qSDdrKHxhbj7I/UTjAY+mYkoHZIixD59UVMqiUX0MfwWlIaU2V/TlwR8bQ7TOUnZvlp3
8yugVOk3Tu40f/2bVVlt52ERmhfHcXE/nVNixp9mO4X/UudYHWIDLatpnbQbgPvgUfu8B+NW1Lmh
EAglJR/3m5VfClcMLRwhZSANjWYRoJvjVBJd0tYlgs7AhZzfO7RhFLonn/oz5ttlY2lu/jvhrwRz
rzt7wj4LIq+qG/F2QtyYCeUWIZU+jY5PGb0M82U6cKrQssqrXa8rehf1th8Sq/YsX8HhqaWGlXm0
of5sE2nLyZj+sIEQXr/3Sq5iDacRsDr0PlCYnoijOjTv9uIqYjegdjOqAgrNEQbxINIB/M990RNj
Ietmn9vyVqtmwQej6cgE8RUymJDqlI0KC6a7nUgUHM/t8h3WA52m/AzORpaslJUbhiKzXlxDZB1C
FEvJ2OHLPSpm6dL/pooFBG0Qx1mJk3q249sWDR/qp3rVfNMxzeIWvcaBRf4mqyIZp98efKYDHEU1
7dnxmqfxxMIvvGXQ1Fvti+sh6gjtSmXoZA/qZxhmACR4UyYBLwrxDODAMR+afQd0DOR/4IoV2JF6
lDYBuQMwRfdlydGnix1HNVEAesw50XoV6iWKjWuB2Ah0l4lX0Yn6Yim27VrF1aAeSE4fvYor9RM8
IUY/BbnMuiX5qRBxqG2Mbj1ukyliS95gdc4/fVUb/PsqcMA4B0lwqSb5qyaEyBgZlDm28kJ4IFZ+
ptP4i15OQFsvpup/3ZHlIJQWsbjmrBMOv/JJdflIJcziJKJk4+AUJEV1+/xg07RAG4BpiyV/CgO4
jRWweE+TzrF+96d+lcRSsCBnLfVDeHrZzn/v6HYbMAIBN5cXWctJqREkYKYevRu2ni8bx8lKvU2a
jpeeyEg3O4lAkn+kBdv45/cRP9JQ4gX32VBBk55wapR7BmMMkTFPpc+3QtP+aznZgLahKG4n2uhb
fJX84l2dL3abVwynI/Y8L9iNWpVwdV/UDSF54xhx03rJvAHuMSd9Ae6mhIwN+AEFND2EG7y96z+J
ypfVM+d8VYuAIK3gyvOjykNBo29Q1SrQxo9Q0zk4X+OtEp3vBs7VBUPggAQ7zPSbNLI4EVBF4JJg
DPoOWWKveiHHS/xA9iCuEidQSj82DPqLB5EqFtUVdf5xtcAo/eYH6K+5nK3ggzrd9y0xyynBgR8x
yWYyHV2r141FLdR/RFwgfDA/P8Tp6C6bFefHLTbk7o5wjcGZnX+z4GQmk+Y6aP2tkSaFv+NkjB7B
id6IMF7AvRDswO/nJbTXDs/fRDqfLLSFDSGi/sUge1hqRy2br4TS/JRjXflDxHW5xRf8CknG+HYs
Wb4Gq740VLmquuTSVQzDc6iPwhe+CeMo1JGAzqlg5SpeL5IWCJzPax74Z9zE7tdfunkKivJ8iOvv
lFYQ62uMzfO1WAVZlkEeXB/6/eYjYrc1ErJIsigsC35TbNO9re4TAr6Z8T9ngQov9W53eHpQfSvp
BaY9ogPuV4MD0pcICVmxq68dZZnKvXT1ZUHvZKqUivZjk2xb0S0KIjmOJYp/lunGRRi/p/qD3Lz0
V8/DpEUrgGDxdW71d0Z6WcIQ7X3/3zBaSr9qmiSHV6rCDdC7ec9YReviNmoX9Q9QMhwaIriLahO1
bI0QxVjomh0ujwbTy2nVUOj4L7K/Lb6Ls6RGRiKiXj1E8kLDaHQUi8eMHszYPQVHREFJfnwzk0Bl
TMcb8ZpcDwAyzobOwIp5dTAKgdHSaIA5wAgArHPah3wtAsWJtdW5rduJdT0cHInOpPHwvpaW3tT5
N6GZMJYXA/w9Z0z9ay0p/ZsA9q1EwcVi9iMIqeFWTQf0cKXwKKgymgXdJKDR652l0FxQrCvDoTEV
0xCtRKr+qqqq8PSfnaIG4uN7rSbKtWdBViPDb0fS0L12EEykgJ3HlM6TxbLD1nbVUZkIemhxkfH0
i+PGDG+yFF4gRZJtH0TtizM6m4Sdo4SfEzgjPN61CAfZKzjJUgj2Tsx6LE6dt8wzRZFEqbC/I30Q
boPHuO6c9N3ZGbdqxGG7YokZDQaw0hNgyNct/FESWO3qQdql/G85QtaAiDhInDmn1zSCfPBPEnMr
0rmNLP09+yF9TPrhGvtXpD8KLKzocm7EqVfpmpWRuqpnKNpssMpso5KBREigJNzQe7dQdzpiy+ch
vJ63kgCdTbJ0U41qFOmSz/0jU53AcooJPiIza2vqPzpt6yN0MhZir5OVMz9kBU/6mXJ8gVPHtAyA
riqnJXubiK2ukP8QqNF+XiDgEK7xJRbWbKxNzTkKMj6E62N+q1xNgVdhNR92pqHRkH6QM2LeyRCG
gEeGXCqWnDbZZr1rGsgXL0OszFmLcZtQNAPMZAwNqdWVn2+2gkXo1xT7RmTqLgcJ6rP/Wr/ykmPt
b+0ZWxV3sLCzUzg1G0IDWPjiGoP8IQzylt6Pwe18vIxtVGnt44xhyJsSm8UFfgKEaQp/K6aZ47ur
TZqBgAr/bfYDqeZdWGpX16cwTU/9wzJlwt4jzv/NCdndtlVWYdhYInLFaUqqo5c+iHUqK7KGfacN
Az+4jh4Pb7WK9Dohamm9U1vgsfYLl4jQfAu7WlRcNbFoyNBXJ05dQkyxVuuGwZzYC14xq4TaQt+E
7h1ooyniRZVPfnIVqpWnqJasBk+roDXorrhu5xFyfOtdMGPJzK6SNbBqKMCzsQQxy2z83VIAhn7I
A60FHBk/qVo8ig0uC7H5Ph1vQ9zUfr+JUtGksgFvRv7Nu00XVgnBO1xjSDjap5A2vaNxsZVSe6E0
i895eeSMy2h561kv8efpl+2rNyxa5l3K9uGNcDoBg9dMgk4XAzBe+A1WYy18sFXfIcRDPQUVTB3g
jD/d8sJNeA5EjSe80r/uhc6UVvAT6sSy6kl8rLc6Os5Cx8hJzWpeOduT9LqGIFpWhPAw7UHWexS6
cLNZQDSPLZf4WOd2WAGeTQ9zYVNgb/heJcFm1bYVCZncM/J0diiq5mJmHH7HryJ+nlT+oCa+t3m2
Je7JojV4aFxPw2N9bthQlD0bgT3r2cTD3F9iRT8Czird1e47Yz7cEultYI1shbSBEk0WMZvPPeE2
F+f7M4FN3d3Zo6638vQiWbDz40sJnfmW/18Hw7wvQU1OBKtVKNq145GiGjTqc6BMU4IQ39FDP/Nl
8XoIk8puzypLZcMsF64yTvcFciEU/8l+UctcL8jradTSWCVNjNT+eNkHUCDswfnGe8iIJ/LoC/Th
O8MtNwuUCnNOkLz5PMZgBn9CHPxJUpj3vDTTf5ekf1EzBZk1hX7V4PFpR0VNmeAGds7VDwy1T2lY
IKc8xy4mLwZaGe5wkMjYhHlGixzZe4a32IRNrNpPNLzRyEcHxoWzcGzhyYiPzMaxKLL80zfPIoEe
V+KDCDLh/Hk1z+VgFUktodwdcb0MeWtbDXlbbeNGIR/yGhP7ad6aa7HnoOsVsa4A4/k6cv3WQbJ7
s1z04XXDL96dd4bx2pPFlQADy19CVOuFhcm2pqXdR3mAzFrafWVFRzhvc2ZlLgyt2vzqZ1Kq0vyT
R+dwe7be29SemSx2bChjjuqH2gbrttR40f9YYfMRLLoBDWb+elTBpzeGnEqyOoL2YZ8Uh+wIjFRU
6qPFR6nuBLcGZkFmHkKA6PFMH2ydjrsEWshWwMcTvIaE3b7f4dM/lhhwX4iPFfLqIaHeOK/Y+o3j
mLnG94fw2xrCSwuiLbRZLxtQuTVSx8UPBivjpKtkvtMPOt5D4yT4oSJQown78DGCIoM2uyIfAy8T
lv7x2ClLcoM3HOfUAQc9Uoq6OxhmPUdoZGhzC71ED+Da6xdpNLO40oSg/TNoVyjb+TviLbdVsH1x
WKLkOJRVQ5B5b9GObH7RxLdrC3ON0DcfBKvoF18dEYTJkdVAOFDm9mGBEb/7EwuafnR3obIaIqTn
LZ6HUWAIeRvgVlDaDqzcJlGZy0DbTY/X4n5vqeHD1mHATZHVrN91PvUZ93T9PKZ8ZhCWsrhSKyvY
J2YAfbwjl3c/M6NRFnO0wGQLzSxgL9skkOmtRDYodVfZXR1UDoQQJN8+d0hnJlBVx91XAdkCQIg1
1N6Q2iiJugOZkQl3ckY98mPtIocmSj/6d9fP/Sl0bczMgLCwfXyJUyNKlBz9OYRzSfDKz3wc1anK
1+ZFR1UoJcl7ao1tbCDnz3DiFwZi0uN3Se550po7AubyqUXXWCnKt3EMg+SEcOQhBvbKIGmEPwun
Heu2NpLSsmehlZvxwAMLhxisiNOoI4lSsVzmGbpB6FBC4vP8Dnd32agYpCYs+Pn3QU0GANYQeBJb
ruvU+aPmkImoUDcET2590lEQX0NT4Ryx0ZJCwj8OzyQHiq8Hklmj9H/Zm3dNEoERz8EyWgJ3nTkX
NnHc/ogvGAIDjclMLXte0vGcm5XDaSz5rAtLwfkD2Ph2gH83ERXsczF4B7GI4wGkYc8PhmApICv1
9MP4+XIY3Ps2Jsga+EQkDe5KRwwebuoVU6HWP5x1wCdvFQNbbsyQ8MrLzD5j+q0WyLZSLtW32x3H
SuAL72FAne3cXZu9u6/VPsVmcwbpIjgbm87GEJ17gNzcNcLEKyHYLBb66XZAgQDqT8ptqWwGVm4c
4rcO2o41rOlwVlDfWI6JTikEB59NmBJshQE7HLppvCpDkYVP6pvvdrpxbX2+cK5D2P+tWJkWCB59
pObxuHGdsPnlMdJ4ZYiKl7iKwaqXIzbLgm/2yzgzI9OAYiIQc4IDPIj79nZtQODjcyrA0xWA3lpJ
Taavg517XBzTrFQmSHRZQVJ3EevlIYS9KGW30RohAHF2cZ+COn8GQQkRWvcdgvAk1QJHlD8BtUIr
VShzTPYXzfjMVTGYcyUvR4DPvPTYbeBB25+x9uLTn1IUbEK3G7EyPMQw3e2B7qTGWJm/qaBjAHyf
pgErGHkCE03uoMw7iOF0rnd1yulD1I4hrG/Xh+zxaRUfuLqtw/w1KILoIdjAydcqS1VFZ98Gvkfp
EsR2F4La0lsIvZ/vy7vpn8yr5yiPV2C6EbSGPvZxJEY0wgwJ5c5eY/HYlV47MePo1v0J29wM/Y+z
YmAmbeFDXpTvDywvdbyxJfwILU6oinlFERSXh/kZP5tHMcufe6OAZGCc+5hPS7xxL4rJx7k/WiAE
37uURmdUMr27kd/KEbDgy4ZMBO5RI5V1TokZ76qzOtgqlNf6bev7YW6sm1/HP305cIy+9tprGxT3
OaS/iNWmj94NmYYaVmlhMnEl/nQ+PZdZmeYr0LkvAdmxO4E1lMR/o0WbS4FjrhbYiOebcLbHS/Vc
s19NkdNA7BFBDzloHkMH8Cy/J0NQfi5QxgTLfYAy2Ys07jM7rubQHyr7/SD83oWksOU+rIPk+5Nr
2XelLmT73gkX+JfmQlvSyfBBcrXHvADpgfTVo2X7Xs07HSc/rjVnXUMw6es+0ViDnHnfHHUywlRv
yT6UgQmSakQdECl1Z7cMMKcXAVXOkO0oGErTYQ0zN352d06mbVWIGkrbSdDR3Kom4pcQ/WI/LHgl
I9Ow45hzc/iSdwmBFxvd2+V7bGZnFu7VEwptY75lVH6LcZrkATUMBN/YL8BuaxM9WL/HqutIDRMH
c3PvNPEsOUxlM0zYMdylVyn9kj9uOWgiC+C6/HcvRme9GoxE/dKKG+Ps1TBsxk2nWj8zLuEP0um1
MM6XEXC+hr2+5+kfuVpaSH4/yv7njjMz4a8GG9b2zUrQayMOxSgWwHEgrN337xiAUsi5nL5g4xD3
yqSxFk99ytHlSG4ZiTRtZnmHu5EunqxFDPJvaG+gdEeajtBP7OQ+/YAfJvOvDnMMnYtvMUMlCmvF
V7imRf47+YfQmLdxjim8IazAm5TeUEfN4AuRv3es10/E/XFfbB7UYTaTvn/Sn+sq1qWI+NgLOSUE
Mo/KFq/Kft1nAhLKazS5bUFi0LXgq5eEE6yGa+XE+HsrCsICxSh8MGVY4kDN85E92c16Mj/VtTzK
IK8Cp0Wwh598Xaz1sfHSIKQDEWe67tWGnA2J9kzxRKIkaCuZiTyy1Ds/p5Ct7tjPK8qVAoFuENxB
5k6Te3tlMsWu0z+9x6jqDrfVBxk828bocuIRBQ7GRUZsWzBzLqh/Z5olFcquR4ODHG2UA0brr8ut
UEcn4Cjp2gb+CH1AdmSrOxUhH4diVmEkn8yl7EOkkurh0wrzjbepHR9AWB0WtmrHSYe/WxP1GHwj
XcndvcB4cpYcGm+IxOk+V04y2YgRno0qr2gYDW0sJwtFR30dV1b8btxIMKebvBWfaAGiNM0+fV/x
TkInDSU5qmSTrVeISYz8wstLIfs8TaXz/6EZFHPPPbA4RGCcrtk3nRvwRSUMAhK+yyslrCP7AqHG
+UTMdPOXXFGDi4IEhsxmO+6ojxVOwnmCj325TLKKrecG2VkhBE9SUVoJo9xgWPxa3A/jIFF3WV2P
OUkIuQqHGWzw8LuEnpSdS3/7bDCgDl6BbAmGbt7koTpGMnPxAKxQn4yWjc3nYHCG+p4lRnjkWzWQ
qHqYkDVhpRThLRkSB5Ec5sU2eEs3ALbUQwp3tgNEz1Cv9qWqjgx11M11BPOMV+y/yeP/dVFKVF3h
n46F84yR/Tq2jKxyhlIkhmxRTRZzPndiRndrmAtOoU2XKFZflxHK4aUSo2CLi+cVtZQB/JyJhoN0
dwHh6mGbAK3FvMeIV3OYt5bOrXunWWDhX2+3fNnHSp2vthR/8McOZc5aYeiyOQxwoJrqcg1ibhr3
LxTCn4PBxoGT/EVyijbbei9xC4CZnmoh/G30yRBC36wgDUX5D8e4rtwEkJrR/x1U18e2qan0Ssyr
O9VziBdFwHTkjzGZ/waDb6by3ypcptyAnEoVYNTHiBiMVLcE9KfArxnoulXqxESm/gTWSN9NG59u
YhNiR7/ys9jXbwg9BK0tm6VWNhdtWB3Do6sc6GSNYSw0f3JNS5iFXFjSoH/p+jQw6eUX4CsVvjvj
sv3Y2NyS7t0Wi7pCnGE2V+OxGyk8EmrNZEOieDB/preX+F/typYEO8aP7ZsfZNkOzz+nqXkeHkb2
9ym6jY4gC6jxruYeJFz0iFMz5+mEHfbjs1I0sgdKNBH8Ph+6OFLfmeVGDVi33zfGqizXgO85oFoQ
VK01I9azKFs7QBOzNjERwgCC1HJBhF8/1P1Mw0c8t0Mkfu71jApFZtxWfIYq2wl0zaxuX8Y5zhI6
WwiKSyb86xl4DJvvhKXd/ItOoLcfKpGx0ZtaC/hfMBc+RhzqP1u/xyMwk4b2DCZD8UgoMwKvlJVM
M36FOkFNseUYSIyZYrnL+F7px9gSQVUXqChtu5KuC/aUHrMwDjbH8x9NfkBqt30GcGbA3YL6AkL3
Bc1gpWckNr1KzM6V5HdlRpNwWNrv53EAp1PAhjMp0uHiR/dazDieVuq+bJimD8+H8ND4tNtV81fj
f72JN9JXxw+m5JGOwJQbu3V0HJJTFXZxmIEdVTGstCzqrNA8eLpJ7m5iTD//n2c7q6LCRZwy+gDB
6u4MiUOEIqrKxdulOUinbyretkFVifi2FaiU758Wb9RJ9goe8IdETnUxRcnrhHEBCsIs7JSSCz6X
ITg1l2KOkyXvjXiOsWBj89Zg+l2VMGkyn+0WoGJa9eieXyc8vc6Z23ivpO5eQizlBNKBZzGeHZiU
tCbcUvg70MnO7dzSgdConVcjzWHCRRxSWYuJ6biREwNpWfbBcH2GB/6ZAA5oZAQDn4KbBuIhU6OY
83mSQRg7KV4DjSBJIk7B6Q1fc4ZUvgrX4lLSMvE7BzsFe7Wyrjn3dOmW3Mu3Pn713ksHqPUtyUdA
cavRJIpTH1G10e4UVS/LgpL0aqXWzb7sDzli6WJ6kR717GWIktcT1ZLL8HdYSjv2NcLh/AKTJ5Ba
sk9N63WoQQuTQRJz/65nMivu/EAoAbl2kIC9MaN3CjQTCJ3xqw6BHqOlX/kPifh6kE6KEWy1iyTg
jN4MtMP4PFDuaaTF4ohXN3h6wnuEaMjgNff8FDKNemrOkpusZ+nk7L6u6fU+ywJOqAMLdA24+saQ
XZNItqQiLLuJDOJO3ajhCu5nMrkfcY5u//gFFhjm6dK6CzWsF7ygjGr2oJftNlIGFsqM73gBh6+m
Fh3eabPLXIIRIFwVCv7CkU1dKUyZ4s2NjKuAmw/KfzXCwJD6z1SJ9Em1XTr5YZeU+Zrpe2f7evFL
RFtka8kyv/4jl+GeShaObWZGZe9Tyt026l6kfcI2m1jGfMW8nVEe8pOQ17TvTPpumexjulPVboH5
6d+wfuqCBfFm2lnrjRQPAWf+pdLq9ugWQuOUQBfKDPPo6uOolBMfL/+o2zSRNxi5x8AwZP/frTwD
fa2ScV7QPlYevbDSR0NoSIe44v+uKKHZdy9PRWntK0i+7gHkM4BnCFZLG2dyrUJxnVcLkw8ihQoZ
sShEWqYb/rMxkSV7jSpiYAvQkkVQguvPGhTp2bidr1HGkxpsiLe0POW4e5bZgrNsMe5Pn28WtWo4
ZGFpRHDJj3nn/NdbOfK1fJmZ3wO5u+FYFMt//4FYeDRdvmYE8xhR13HbhdWEpYwWPeQuusM3JTL7
1r9am4NsI9LC6EpGuKaihmF+LH3GhVwWtUIA3mDdwHkHai3+sx72kaa1JCz/fkPEUlbLIVm4lBB6
qFYWTEHZE2xyk9/sc+IGhQSqlZ4hZ4Jz4GagVvij5XYb+3zZsHs/3yVAZrmvB1X6qzqeQIsAKoLl
n4GiR0D4/hz5Qwx4TLifss7tr1e4MsMUNarS85NNnGhGzdyRsbOn0RnE3ul/pSMrIOJ49r2tXsGz
ei9blikVfFeNcZvyUa5x1AVnRdgXOOck+ulA9a5acsPbIxXYwhyr1xk+q8Rf5cOL9r/kUuLI5btF
d/EJSc+Z/nXJKSkKa4VAsBMSHelxTnaMYREplJG3oOjO9UT/vqvR4mAFDSErK5mKlCOEexZ6K5Vr
/LDMamcjc8dleMU9TmEYZ1yqxZnHbkh7jAYXgkAyXPVpRXwsUTSnNZX66kWk+gwjtcestdobtnOU
frcXrFuMsopQquxw77adCznDIF6D+IqYusY3ZwvbHF08XMPBSWJcWR7uPLQOaGET4w44NIczVDnH
oYvy5msOQK2j0dN5J/Ra/1pQMdqxdfOJihGyoZbI44mhF0BggJX36DDVtpnFJlJssYqTlzfzz73t
atMcbhucYySLjm4KoUXZLn3os1nBcmxEdio6JG/VcpHJIPhsQZtwhTggKiQQUhQPK4gYD7tBAFc7
8azzSFmBo02Y3Xyvuyrqox3ag0ZPojXcqMYyydvI75RK6KsBB1+CJQ2bLEbaHJaPy2B9l2MC9bpS
d15Jl+VXxte52B+Xeu01K1/T3IQsGZm/hFTNxB+LevGFAetvyMcVgqODFzdIagEL05A5/shjrCbN
lCtB8A+ha/fW1JvjwNe2rON+v9jaDIyyCB+bOxd4m3sRicJTvcXlByV4d2LSVuQZzG25k3bPB+rP
EdvMuH88/uZKPdrL0jhGnDx6yzMxh0Bva2kPFKcYg4qwiOxqP9v0Vr8Px+i8xpYTeDAIIQIwDwnV
Qvfntqw6+Tq2zXQ9wJYwudEeD3PvOUQAtiCLSVlS41u5IrcUV/cl8c0ky5YEA1pJwzrbbdWwZXOc
Cb2aePD/SrFUGZTuESzaxBH2rcoMtM+kyqvf+V8XWM0qTKRlc8JHkygpOBUf8g5L1SKUc+h0DghI
UoBbsUHe9OaCRrctG/e0ZvvOr0sLN2zct6N5B5G7Wo4cMt/oWRq8H2773AdwJ/YyujkXSnS1LVg3
hBF9XUZBjj0YWevga2AbTOzn9tcNgPezTIIFYIDL2XKqC83Q+4E+d1nQGwZkMQDQTQPyo6OcO9xm
P1uS5cXi+WGoJ+srvVFEzoa7EufGwpGRw8FIdZotWnmfIW2Pi9AiEOXvSvh/a9HNHqx/dS2YWJ2F
zJIUPIK4U8C+gf7S+UG5RHcbKJ4VVaLN2x5zP37MQt8vuj6A76qePkhKWShe1XjAbdUhrhTIzqtR
Rs5aY5IeeZAgqc/L8PVbdVzlU4KXH8zlVXLDG/c1TdyhC67l6LWs+k97x/P30HUeazxj9VJDYsYV
CKXx9U/y65PAmpfRbSdKwUsPB7sY97CWXRf9K4tGw26qPT6DGh5+WcAqJ9bvf01S13f+ooZ5nX27
GTi2wFDlaTuuwnJCQYBVtsoD3kMLwSxdswZVjMMKUM1dGbeYe+nGiI9NtYEqwqaXYoUconWFLIbj
n1+Grw67pdjOAw13dKpPDcJ8QFrB1lyi4sXadlBScr52Kc0XjqRjGaDMIJis7GZbn9Kk9A3uMU4C
g2JAH78HruUVmib2O+tvrkywbk+h9isphvQ7kXRgp/JAaJUtx55VO7y7GJWCNZOFBPy6DugxdlW9
3SUTxL3YgLOMWX5Lwz7Csc+AZhQNhXonANI4d6pOmAc44ut1aWIEcAbYoNbiXGwJ3G27CquaMEds
VKAUl4mAYaJbQnTxYlWzazAxN/I5vjyyU/DN61h/lzvrHU/2Jv9CAh8W24djhg8nTAKYoAh/amke
KfPsczUn1jiove/jwnF3u0G+9RT/rnDcgIYysgXBY9vZjaZLZbHb+UrA+rViijDYrPZ+4f6u/FGJ
+w/gKfThGPY/VH/SLoMhgibvgfCvhlG075wIk/L5DULkEHkrjthR9eR3R2TXyHNvKA8CI/JV5G0B
WCadn3sfzoriYEkuYpNJiIz86S1Ka5pwFMtq2FqE8yn0WPeFzYhCgezYxm4Qpcm2JTrRvkUmao8E
gPqWJj2ceXs9yC1jzjAKKb0fwKpt4AOpHueggYDcZM5ldtWw+3WOagt4OxZjZ5ZtBZvx1PQLJihB
Rl1hFcYhswK9TbKpPW8LFiA9nZyBIwG0KmawVcoYclTI86d9cR1esudJDez78rIFzUvHtTc3djYY
LNQ7plq8ntfm/enLRAn1zzLHSze0vRWOMoMLpySZVwrwIjaKWagUWJnX0LwE8jsN58LICLw+cCd9
XRx6QpTQ0KD57ZmuVMJA8Se2GXxW3BKasHckZWvUPErb+sxa1vLxsxWnOey1Z+iuL3q8TdRUfIyE
EucvcReg+DXMRsbWV3XgFWkalvpChJVYm1o9VBYrHzRqfeQa20e+Gzraq5zZSWf5uhU8JFxwdmda
P8xKa/9jO9XhxPNnPtcpTqyoKwYZcVXf381AU2mNZeJgeOVDD6piG7240ubTVIfcHadJXrKMeQfn
9kp+OxJEK61ppwerF6OpN/1/ood1SG9CTOISxnEVSw63nY+zE2lXLvo5vTZd+cKnF4p7px4/w/5s
HokqfAYhgQQokXQWFq2ycMXueRkLdu+7ui4SdyWvlXwooRfvMeyx05O+IaAK04T3qEpKA6fMeynM
zHkuUvmmvxymCOa82xtjVo+amVuJNSnX5ZMIxcd+j41Ku70m4zAnMLgWeAoSwYwDP5ox/paw6e/n
hQOXieErcrIUVBjhJ+7u8mv4wd7kHIdQyZV16aBAKbL1T/JDxGlfZZKJukp+/4j78m+ZORaGHfzj
6Dz5X617eO3Cu63msiKj8hKG0YiX6Y9K6LZ6XwOze9kCyQDSjhKwtw2vBwZ+HNsoPyszB+N+bzRa
RDLdHA4bu8roZR8X+aor6yaQ+vxUSMWoU2VKfK47Xfp/DG8cY+9a3sXJ9s3btYSc1guzoIWQpzzo
poyGDhuvbd6sKBwZ4QrzHqrFx1c/A+sbS74xBGrvDHZfNA5r0oId/Mso4IfzFRf4p/5fR/+S3Lol
0SWtvZreatdfEqGZAiLehN12hZ1RacnZNcSsfEF8khVwp1UmiqKkWxgrMAA4/+2IvhLhDUs5k+Xm
ycyLnRA3AAf01xDyqdAy/LXTWhyhEyDYVPqKuj+AfYDjSBp7SHYVYTTEvjazzH/2dhJ4lgbTqwev
eJxg+JYWoEmYn8Xb1YI8W7aSNQhXDwpHODVN7iJejvWPkmX6B+pIW+ip95qFN0qjfz8Xlly4i8N4
qgHK/ABnlH/A087bhpIp8utWM6zr0wf+oNbfbVGUIIvNk4ODCAlMznHpKqwxjoy+hq5+Bg62M8nn
10gAOkWaBSKXEc/xxvSDPU7xb8+ruFFpu5SAr/VxQetJI2ktei9aNgg/pe7T4lvQ5paBeo1aJUoC
bmsWNGxnKXcvb9jtQ/+0sRRNDp3Wmti9ZPck9mE3vL5mZOAcMUqKq5vKC7umFzq0N8Dl3XuGlu0n
8yZaXubfQag3lR0PMhK/kZPfDyKQg3PoiW7YbJ4ZVrNZtevGztEpZqWoSkR6okSrwYsKsEfgu3T8
nvxtPxAG3eqVl7L6tbjN8mUsZu3Ir9bdKUYx/88dlXaCmmjxpllWUQQEb6lvc0S+Xg4/1HAe5Ohk
jJi6qoudRr1sLpjDY+0IssZ7Fgq2hP6+lnMsl6+0JoBTaJCY/1sPz/QJo7D78WxD8c6yXTGOvFfn
Rkc1fIPt9W61G2QogdOj6tSNKSPzjD5C2B/76c4zWLQrWML88bkhzNWp2FCC47lHPl+EKk9Udd4o
PwV6sD7A+EhPZvPrepgGb7Z2FTE9x+GQ/aS0W5sVNC0hWsVsxWg4Ql+rrEqd7+sDoxWYPb9VILEB
fjgcw0e1f1rPhDj/lTUu0J8QNtmPqoWZhP0MluZW3gILqqaWHZIGdVCjGS0Iv3indPWSy/zLknkW
+AyFZUGUS5V2BmpUtIwmAeny1vaJ88uLIxFhofBSBae5XtxhLVqwB8Hf7IFJkbVTp8T9B94J1Dbw
qvskeQaPO8RG2hRB2i9CgvfqfxRDBqP/5n3krhRpx4QKvou71iV/j1LWScj7pqC7i7yIXgO0jxso
sfloVVLF809O0Av9azEpC9HeMCLXAXjvmr1eBq7jufJ9ft63/wTcghivnU1Nmin6sdXZ9O7d6UHH
6jCfaF4eELE9vptxeCrHxhD2zJvG0WPBshP/Pk1XfOKh/5dIQwCmpZzvP21Xnt3qw3cqtLo/2G6g
6e3xL9ZFgX2+hGg4AncYGUeBPpcI4A7unK/tWwPejwfHjNZDz4Riyqnhqu+TpySSW0iGcLUWfHAE
yJ9OVQ5hEc06ld4Cz0NgoKkSgQZI3hF0Xxsv26mbCHw0ulM5y/OKd4CnsCEBEbMUkEQiY01OaXwB
lHIHBfqikddAlYl+HHL8aitwHjlX0TZOiYAWYchdkCTWInjG5IhuGEKZ9AR9NbDImtP2TKQLP5lh
hjn7uAyWZYr7wYXY4boZDQIrCuLpLxgqKxXIj6D3P0e7gby61nBEGsOmtEXOd0ipfpp/AF6gvLrC
eT8CnLWe2Z/D8lxzAH32ZtRp/xPUU826UI7o8dKiVqCqpwe8HVDj5oyNu+n6cVnDd/s6WTQCMGN2
qeHMOtu+mG2JrkKiRCSmNxTTdI7dHBYhe1JoDba7KYJuwOV+WxTGeWjAsosjOhPpwWOJQAI06YSu
mfMsWOBTG/d9IS+zj8wA17A8XD1soC4UJnhXzXMz4k8ev3IJW61VjdQ5i5stIWQbYjZZt1A9Mw3k
d+yO9NIcYvqZ3nYSetlwqxis7oRF2PW6qMIWtcx3sSZrCT+yRF6l0FwTvrWT3qKsJ4KHIcIGpF/S
094ZhRZOjdwNEyxbmoZdxKm+djcb66IUPLc0wikmPbNgR9iV0a7ygHJtYX/DgHlcdUz35Lj19FKO
PX6p4MyGqWdoowIcxdVHP/zyR1gpZQtt2RPqddKm12UX0pFSqeMl/zmVnxF38b0X1gGqbx4JgySK
eY/Yuf78mxaSUifgDyvHb/wzcQNTTSoIbDCbB2aKs4jUvQZIHLveP6bab0Nv5a92duqAL0e7gZ/G
rinAR+78YeqN1Zv1tEysaIr3AROSZqx4Z+XCy5/4KjSqyKjgpSZQp3LSJh+fMbufZ2+qJVHt27h1
HxrAbH8YQw0+W4RXrWy8IfXJ7RsJwSYMhsNRLlDAufPlFTW2dyyK6ZSC13LiwgwwUOUgHxJ7Shvi
t+BCyOHv3UuA10dcPrTzj0jMu9sXrZpKszjLhQGhrYD83l+3A/19hm0ncD14GOL997ooui91dwuA
NnDCCjSkcGbnp9P7DSwC/icRBxNTj+/V+V8LvlFLdIzpSb8KkSuKjdVzvlxQo7CHvcscN9XfavKf
I8hwcmftexv8rMnoCCg81qGzLgxKtGl0GSxIawZc8+aXju81osyEm1LOSsVdXcJAJBcA3t3gpePP
8dCuPRCx3ltz7UbT8pvGb/J1KYio7fYxEASqlsmT0qShU01/PolJoQt+pZUu48SCal8HPuBniZq1
z8niS8cJbikcfvYDPUtmpmYaqMh39mfThhvP+u6B1nyjRyfVB+q/kZy7Uj81ki3AnXF0ER5MuUTm
CMYA3vvscdKud16MZsgCVqm3P3oy/G3GBHIcjo7aE1z/gRybKeREUHZoGzMFMRmioFMcPtvTkAzY
L7WMD+5CKXT4+qWQxiziMb1xc5Jw4CK18gcWonZYVbbCnEigv3F8/2qJTsFw+Vd1/bZj6n5uBAR3
R8zx7vz7WjIrVk0Zoe9FbEAs2kMwvV4oW9WJnfaWPntbdv1LE0WLvYZC75poLSY8rgJaJfP6uTzl
F8mwQJanhCWGrjedH2AHxTfoIyEn19kFJOv7r3d5t3JR/wOTnHOgW/PEuaDhfjLDA9ISiBL2Z6wm
96Q3JscmxOFQbfY0fPRXQ83NK0u5S8PNyhEwke3YK3UlshEFwPbkQQym4KpdirV4vj7S0grI/toq
L30dHe8SGqpIeaARmtl2fPN/8+8VZ4WC8aelc/XksNJh02Gg5jcpNSrwnSqBw4r90MWtQe11aYDP
4tb17eE8oUmGW1uAo6XOIFuAXog+O5bgkwKesbG0GI8fjFv75a9r/z3115uHz+D0fEfjINh+uC4M
+sggg2g2ueyHwNJ3P1Nu7T9TIGRk6hdwPsI5YIdB8pXOl21PE5MFKS/RRuvjYQ6B61MMYMsol3IW
bfAR6JVEAUVIfRrfsHgwn4mxhPpbizucsm6edAF0e6nWHhmdtSzNBdJZNzA8XaxgnUiTX6rgCWaG
rJ4joK4Psenbjo+pIRZgvIF80JFRKY7KQSRom8cJ5mOugQf8e2u1oaRkis18Stasw2YAjzznslor
3urwjqYvmvdskiUReDtG6Mk9E2Rkns/9U1wEbIEiULiu/LSSN3ZmdqtZxMhUVYisxYisb1Oypvtt
Bf2dpPxZzNc1RYyjviMqe6ZIALQUKuLzBsvnZaXmBuIqBer9aTOkrNlFJbir0tOzyIEO/WGZ/Avr
JWMOVevhZQCJV7iTRzYayH6d7HUkRerrpRB85rkS49H4o1+KQKKOfI1W/2hN/mswMBDM6a5KKpZO
LCiarlcW1cLkNbo2QjZmzlflooKI1QVDbPnlNIYS64ebjhx4U3VvmwMz4bZ81JpFa9LxNzMdCr9I
QHvINw15FRnupeukG6mySCFi0cIYgwNB+Ji/93X+SQRqXjtDn6+OWjqHXOU0oAoSzy9YY6kLJyMp
0LdI2Awz+XDOaTebjfOIKDgIfHCreNTqZQFTNkykkhdAB6ln9CL2cK7wm+CuVOzvJwIE6aPyoMeO
jNesHGpx7CTjvUi4Pq9Brb/KeVDUuwocZIQLb3kEiNVUr1/fEUU1fWgP7mQUAKQzGDJNC1m8j4da
2YHCa0VTEDi96ouHN+lvvONglWij+enKX4bAxKxuRymFMUvaWGmciAkjZZnyhqxNZAqvF0SIy7Fq
cORMebw+S4BchhpweAW3PeimL+rejhLglUGJXT5v3xOqjuFEZo8hw0+vntWtvCkicr9SN9xOrhHt
mFe4+1JHf8ZZbbcxO576G+GPtByj5mvLRe2E/oaSLHOZq1RO+H2ZMpPFlz1fGu5CMrnPe7b6hw6M
hnzw8rstPxKdxBrFTm/ch633q8O0NgKMtuD37V+qoFnD3zG6+taVLqDpILhsVskMRsfGN+cQ1MQO
nB2oNT6fS/fuiwUnAbLB34GyjX0AawYSgqQqOM6tBQJtIccH0C1XQ83mVYI35y1D0PIHd6rGGVQw
lRU187r1HGE1DZ6JkpzG1Kah52OxqHhS7ZrKAVGWTBokaQOUy2uHjKxz81lwC0BONHJAi5EHKMGO
9ASkWhvwdoafhCiSHNfXKDLDL632ktrF0amLShfUhZ1vQe11utf3aNgNi223INujdaZzZkUnGxTb
vcalItA/3LM9cm/jIRnI2U8IhzzV1Vzf9kqwU7muzKIpo5qzwbiia9J6HQbZkwjcQIvNw+QfVj6y
4YnVF92gY7AHSFKnK9XX6k8HnAuEZLWMWWTHQakjnhai89w6Y1/mEkk8cL19lFqWSod3lH9dKlQ3
BsbpGroPUtjUUs1a+1W2P5aT+cPS7OHDIrNvTw7uY/q3Q2N6pCEn4ehij1ag0VRuN/EuMD2XtDuA
PKf7GrfosQwV0S2Pwskp3OiM9ZPIYUlkmssqvue1UsCaOowpzb78uBj3ge2b6nyHuCORUQItOGEQ
/CwvDtqum4cPClt+mlj6tjJ0JZaf6ZwNf7bKobmm1wQIOXofClH+MX0y1iVa1o26hI9Mt8YrbEJh
1/VcVS0WAEtONdzdVBvFfnQOZiGTy3k0dIS7e4k4OSRVXDb+82qqJfTQ1+O4MBr6l+wlAEBTR8Y5
FB+TnoTiTpJDYba4chNE/Or19+jn34/l4Wz0Z0FxkbvsIzvCzts+e5lBHkJ30b1G/JG7nzUq2Kyb
Gg0JnrrjlHBhWkWGxkqi+TJ1Vt7oQJ/8B6sogOk81StytHX5dKnDPTRUvu8Tjku3iC8ov9ZMop/u
PVTyuQ57thjSv4GMfqNuj+413IGut35MG2eifjRqr3+4zBSoauZKC6nHDsbWaT2OC6iOmnKAW0om
ux1VG6Ju+yQuYi9stqWOfi5BK+25gKi8dUeqvpTUsWgzlZMK4m5me1PaOR7dM0ljALPbWx0tA/eF
xdyO+RzLVdeqLItnRfQvgbpr07O6rYy+03gBiQiaFZxzyxtZj2wL1w7GmCULE86pnA6N3IHQZmWL
jwJN0IDVzinVJkkc7zEK/kkGV3xVgzrE+zm3kDvAqaQnM/IsidRDa/SMx/bOUjEvzbq7LecipnSH
atYeEKKL4PIEy9wsv3aim4JCRmQpbrzx+WnFTeX3irJoj2M8a6GxrYi00u4QLtdQu7nOIHf+zLVJ
8WvKGHLep04Y5Tk4QUOVBe9OAqsTqhVQyMCQ7ItVDgn6wYAdzDCNd4hktiRx3/1nv8IMXxT2gjIM
JORgJWFBUTOKwD/aL/tKB1xv25BfXRcWw81/PW5J5br312VMGEhLB86I96Tw/iJMDAU1H4Ry0qQw
KlIalrL3zTq1NrQwWUYf/g//NLzuWcXXwA2772szmjHeHbgXLakCudSpzbOro47ciDp2Ue5jinHH
9IPoSIU7v3hf2gQvrQvUpsDjZZMM0NRg+sK0y753UF6UrJQZEKQ0POg3NTPNoLMbqGr8JouBZyt+
UoH0/cp4A6j5cscXTHkpg10xOUVz49OyjyhLuhzJ7QY66PPe3e1ASsnSH78ZQ3YgdaewQ/X4NehD
8Nx649T1U9re2YUXdK2hIPoIzodt3E/GwNYWBb2wlNox8lgzktw7jnm8rlGOc4GKytNoDHfkJllj
g74k1P9j+uDUVaAyimOLxQ2boi0Ag9jM1xCXcTt30CaYexsu4xkBj4S4/TKI8vjRk9yuW9nzVh2M
wU2klKtMySLhjqJUBC9IHaxYlhnMOIGGAoVgy0zSjR6jOgq1zQG9vSyV91Z8zWSKBaMDKO23rWi8
80ioILZHUAWu8tSSNIAO2lUoOE/A1hdrHbtnfSA90Aqa6TyzYrBH0877nlHhPKzqGqRklzI7BTGD
KnL1w1HGJvg+cWRjEmOiYnENN9Ufmn7XArm0P+CeFksnGYSoJV9p/X0NHMgXbnJp2DGxe0pJhRLe
T9BeC3BJVdCmUlN/g72W5O5w353vsKe2fiHdAkHy608zqyodCz91CjVsRs2C03hEyqttVj1GmFQ5
QBRwJDUIa+8qS+olpkAdJVMGiN5sUAOOPU3jSjIbJ3vRK1snnAiINfFExCRRn2cBOlK0ymV3Tuws
Lx8zeGBC7Y6l4wCyIUISDVa/Lk7R7LGfr31xetp3+onAsCLt4bE/eRSW22L5jknT4GosU8+cwZ/E
VO7rZ6Hw62WW+HyZXswct44rMy5dLTldceRu3K/24xT9nzn3gegP0o0N7wEEhtc4RMhROd1RgS75
EgWW/3Ld0eUZ/yTgyUMerpKDyQxUrrBy3mT0If5j8mu2++UdLqUzZYT1/nVQJKsIsNbT0eeIC0vz
YTWWaN8lbPZkmVTbzY9n+Qqh9YH4uMBGNi1+01EcKkvoVuvrbDfGY+f4Bpix1ym4jHeYwJ/ZvjJO
jyo2GgvInTbbgCKyKlYnR9454lrUG9LKOj/JiVLtzJ5vGINw/7eb2Zn4eHVAV0kLcbVgZpjER9kc
QZ3Um82crqPZKwwllq5pIufFeUOYC+0hctf5jHLeS/T9rAzdOsc3c8pW796FkEYaNDlOotI8St1k
95TlLMBqyz2zCeN4hI36PwVhZDUFRv2NtbLO9hFjRdFYRMQTAZW6QFifzf0V4id1uVeTVNuGMn3c
zGQe+76Pce/gipivdBwb0CDqL2WFC3Grx6Zv+9lY+mz6VI8ZcPOCwxek5PBD61RumJr3UGYprPGp
EUx1+e3zADTHaFJGQaiiINIyQqVfb06R2sh0UZ3ZNZdF1U94yaIMwHyl+jXWXDgW5wnjTDqewHjT
t29w6SDhD88ZgviYwVEjecLsRP2c/P6SkNzlOZRhEyPHpLgAVcwZvj55UnWo+Z7sOqN/BDyfbZ0E
xtmHeJPSd7+HO5oXl7UqDcH+tUDDzQVsjgwyXyZgVDIoYeHjrsphnsSaxY2zNjUoESsLIvDRaJZA
AAXaCSFu/jNxX+XQEjnlfOBtPeLbOVsmRrQZsktkGYTprmoTfudo45YiLfv3y2J5VD4aBUI8YNRd
FdPrzO4/sNADQwI4peNwzSXchIn4MJr33cP18Prw6f5omztjrRMlHAGDxRziyN3bDau+zkmV3H4D
U6Rn2Bs9mYUJdH3La0dsH38B77W1KyDooyNo483/Kwl/Ihp7QhFCClrHHdqk+bSIXxODXZUDpJ/x
cHvmSErzOcffyd7Zx+FqViYME2rUK8MNyc/Skb/+F6N0vJmIVr9oXFaomAlUWfBx8yY/N6KNPPhy
vHCZyF2zW+DHj51VOl13OlxXdxb7HJqp7voKeJeU1RVo5zfchmDjnimv+wkCkQGwJ+kADIKrfVvw
cVWatVga3op0YTK+peqWQaB1eVLDNrAghKO+4QZ+StI7jkPXSHBR8irlTNx2Cv2vy+TE3WGQ1G3D
rHvnf4ovbk9KOqjx5q5l5/ZwcASw5hoKMvlBNLWL5eLSc0nYhM3UdIRc6slMvtfWZlZj3MHzBPH/
CFy3F/pqqDoVMLAp75OdalJA7e5b8ghDs8fB0mFpZX7qgr9XummxBHaxHkwqlI5EkBlGQOrWzFmD
/UyNms9GJR6t+NwPthkkb6XjoqlpWKPaOyKHBn3xwwi1UDwIXcZwIkRLareD76C6MxHJ2UyMlM8j
CDgcOMjDl8NTUni71CYQGWbwqMqQrLkdBRBjDWFcyUziQSRmBdeOPDgtl8RT9xYY2uKfeBVeXRlu
ADb9phagFyYAzigm05eRUcklh7wbLRY8h7lgfaJiemMz2H0+ACNCI7hUlm0uayZbss8i0Tb2ncoj
s+C7R2z3wYbfCJslD0P+QK9R48lQx3dgpYYuMnPvq1V0QTuhH/ynw9tqUR6HQPRlAwu3SCC/XQTS
SK2sdP0zBmjYCUQY0fs8Yt0bPm2wtAPVhAfpGucIvM3rcMBbH+8HdOseCLg7kjpb2e0WPAhBTy1q
/JaGawYoT27y6sPO7eecC7Bm77Mf/UhV+F88H+srgcQFjqP+zqVR5JUQ3erT3FwaZwFh9iqAygE+
0Hl0ySqh0xGTh1KoD41DRb2XFFRj9RPFnbKhMzh4LNL5FTBYdBxrBWcsFJlFEBMs/m2dpkIshCF0
o+UGueBFpeG57Kafj52FeIYkKMy+WNrj2LtwI/oiFu6dFbt6m+EIl7MA1pqN+rawOVq2qHgi7gNP
Lwm0QR8b0axiLZuwnrJ+taPFDeDd2YgUqLRKTpOO4fynXm5MGdO849VM6GRGntwJEdrkR4qOLOGW
47ogZy7D9UlbFBVS8n9aF9v3B502J6/aHb9fY4b4Wgefhd6miY6o9Caa9kMwuvyluxZV5NTR+t0J
jEzG7EFkS5Thr4fo509CvGUv1jLCnci2/RS6OZ6Q+hOfOfTT7P12/S16bOIgoJKpRjgPQw1PxoCG
yLCFsLqr2fi6sw2H6yIlYCHNTEPATC3XKHq831tWMKrPhzPdQMXpMlJMXpCyU6MentG11iY7oCwU
jxEgfb3rnljTDhnqgfPM5xRLbv/nITjDAXIQnJQgDSrwWo5gPHgN4/KOMG73j+GWlEKtIk4cCrzB
1PK8ybeqJOvIfQsPn6epiCl8yuvoboll/3wHH9Xqnq9klDDCN/mbNyxPZ3lSFy83lozbfgLnDzch
cN2BC++ERFWHGfXQusqQjrfjiCdRWIWluXtX0GQOd3R8mx9fb02e7jfDoqxC9vhls2TBmNguZmQD
ppOFEwWdodGNNACv4M3WYeN2ufKNTqU0Yh+Rd7G8EV8LqmnQWRduwI4fZ4HUc4/8Y4kKzhh+MFKj
4Ym1ReyxmHhNwFLJGRkJ/5xtZ8adNfqDPCAeqPJpYSe68SlxX5TZ5OPvecfEtOxZvEvLn+N0R8t0
wkxs3xl6R1yT+Lgt52dIYDiBFO3bcM7P6WwmB3oN9lEN5AFaQdTCuqLK2p6KGSXFQbGOMu83AhfE
7iK2VfHLSsSQjItQqRvJJ9Pj7Jh1kOxN6i94/LR7XqAmVGu39ieLDtekuEUWD3Zt26f51DD8UjDj
oNEOF8ttmNL6WvyD9h1KX/oH2DvLX+BQIfID63Db/BVoHHKxXz88Od8jPM0ISzsx7NLz6NOQ3OaL
pmtW40v0gooDzUz8RuCbkCzLIiCxWBHdyLhawyguv/9jSz44YRP5n3XDi4mvx4yEXGkYNBjzpBpY
LDJ07N/v+TwRL32SaA2m50Hsil+zZfWVn+jOhRZHKwLU64NjBFMM0Le/g3isWBUqn0K/XWa6FYE+
vOReuC+d2C61Ph0u+OVkNNZ90bhLLAEi40kLvjWoi//JL4TJxZ6kjcG9r6GBS+gwnv0fy1aqh+vf
xBTXWfTG3HCkVi/4SuggjSWjQwVMnmnkwHekpf90ECYP6Eaxa0QgxVmT2Zc6cdGI8t717e+pYMHN
s2Kj/cbDsZ9IxmX4H6D5QyPfDdlAyQewZ7wKnTYIvERcT0Mc4ZxbjVVnuqkRKqIIStkLSUlgm4lL
yPDIwdmAx/htZ414yJRDPzsfRbdmlBniOB2E9AmQbTuqFN2GpgkDXyRkwEmr+2aKrRYja6IqniO8
QIHODdo2zYDZoPr3E1/OmAMp2a/qpcvauetV2jSshcJWN+PmyvqfA1nut4C/NcF2yzK7Ab6FSWI6
NF9o2ywMCnHEHnpwWnYDqhD1iYVzaHas2ncN3j6mjg6fLBvMIxQT1D7XrOFuNiUus6jAb9k/8kRt
VikASKYFYVX0B8obbeM/0IF+VCkFySA/aLtqbEH4mz4PByFBT5ShkQLTdAYZ2S+913aZHTCeJWa6
Wc/Fpg5fSRTSyhHNZb9fSIENhh4RdEBqXFu4YnLAOvc8KdwK6Y17uMSdVZ0ujpZgfbkqO6/oymfW
PBsaFynk+0OSKhKc3ikoqejgMHBq8Fav9MMqRu4vDalmjMk1/Z3XeMSo/60YjcG01AXE+NWTa1Ce
53bYCpEg4sObUb115QTjHuBeWpZZtCjFmfdF86v8pYdI80DLD1U6hO2hjlkuN7jLlRxmvHnMma++
4mSP2ZdmGSUw/X2xCstQkK6pWerD/g08DzqjTLEY1L8JnEzeLjoFtmJKwpgxDu1IyUFykcgl/j3h
3alePghMGJvVIMYbFFz1iyYES+sJc0h2A9A1GBWQx3LPANCVfp0xEHa2ztxIDqUrywMkkBzeuOTh
9wNKjLUhJoYueX0wHjvXMvJlhLuXPlRlsxGs6xABp1S3M82NJI8YT4szkY0NXonHmZdAQMNC/9RH
8pUcKgzdfWvCM5H8ShHRsTJAgRq1UanVTPDC7zYFmvSxcoxv5i4arJSkLu2+HSOAFjvNPaTNYamM
1q3cAM4UlJo0J9i8hXV/wQqcq6Mkl/AXyLpKuZ1J08lJM0HSIEqmz2lVUxtOaR1WMDGXTJfGGnky
yph2c36ZB4janSJFKU3SsE/zP4UKK68ArIzgF4Q1TYF2MCbSvYrOoFVGBeEWPfX6xC5bZV6GLrPe
JDzohZUtyHGyuKsNnD/4yVwFmS0a9TY7GiDSk65AIXIsVXOnQQoebPM7aSlBa0Y/DGbwdBWJ5Dhh
Qg6znAXDcOqVS4IGo+UAuRZshMB6N8x4yK46MNn9mPebPPqldLIgMRgHydFm5gVat34TRSvbDX2G
ReB7a2rF9xvg0NZzzFK2+4KrU/xwKKQnooacDZ/WZqAz16lGFalmOuQy0gj5qncfmuJqagF/uL1e
l/i403q7xRfLcJDHONOFwdvVjY4yHfJ5C5aQ+km/IOfg849F+Ei+ba1PZStJ94qjUD4/eehaKMVD
ckWoYySbd/gGwRsh9YE8mUABJp0S6P/kYO7Pgo11VBrf6rTb+vmhZ7V9jshocI+YjmSFveVXmV2Q
Gn8EYWNW0WiYgfpHSWKwN13cfjle+RdjxnXYQc8f+R8NfmVdc7Tz+PsJ3BHyBIR6FMDuE1ihJgOa
r577xn/uY1Mnzgah8fJ96QT6RubaGu8DRSxOVZyvgijBQ3FId2+AYFVXAyMUMnTH8SJoGgdy2ZtM
y4elgisGv5i3lVJ8/nYEGTeOjngefS14LXNGXCmshYxLvUDXH22ppmP6c2U13BQkfvr4UI6pUjX4
UwhgSVl8W83EBn/kU2yAUFYLMg6ZqxMMVWcQWjDBxrT2m8Hb7FFiKdcnAjr+Lhu6aHzuIMZegYM8
C1MgsJ+qyKE1DuTTejL7spNdxbSZ1KEIGlUBHV20Ylbx92YQ5pJIXiEozCsV0w3VyATeYg/1D/Sh
vU9w6MCO02uqQdpqZ+1xHQTWICGYdfaYN92h4YK0A57LBFvMD6s1T3ey/qQo7JK1liXi2Uz9ypBK
O7cAabUa846MWSNyh8A94+gHfzGH5OJ8oF4Ss9TOdf/pF9ibJ2BG0/IG/x9iTkc1Y/3SuGOKJHDw
nf0hPuSzc6iOMADO8m8GRnbbtby3aUvFmLL1EEHLJNem0opyRGVtw7CoWFaTGSRYH62P435OEoLC
u1QYsQYOROjQ+U8WfHWXHywR25D+bG4OP2IGygvh4KAkliUFyP+yPffAR/aQk8yilHI2c38zyh86
0SuLBCSmkZKp7p/+kSP0O7MdgaIabJZ/IjpBq+hODNmGRyRhlyknSlT7Tp5UKDAeatvaBza8VbBx
jqpS73ZUASzIsC9x1z4HdEcWep0qQ2SOEgB8Cv97PT+68YArHay7zuijA031U9Xkx4MXk7x/ZezC
vHKi+gBTaqku8uFz+CJPRuQfj6kuHQulIseq9iSAdsUa0kNZdZxwYCYtpUb5sFjvKGO4m+KxxfNG
OjT/GC4qO683jpreAs8EVDNKcrVuc/FXOghy/52CZSo8o/6dp8RNMy2D0rQ76kSowDjlqy2PPi2N
NEWIeQyiEPgSawln9z0jpF8d7tohhtnnqK1nRAv9eb4ctiGxqLmrBfSVL2HH/RlHb/ZIwWux8RbJ
q94c4DkfysRamhcv531+HZD+3IsLsRm9rywBD1XZXMiXEOa/42tP8Se8NAn2B5s+jWWw97oOjFpi
KQRfkOrMnR/e6hW0t3oIulZXqZK2UfOE8s65K3wksWrpbfKJfnIokgCFx8WswmE2s8wIZkRmgXUH
bolw8VB4iamULYvnrZ92XFDIQW0b+TE6uMuWlO5Gq8ikOEq+j7PL/oUgDg0Wu6F2z+5sY0mfux9w
msPuIJd0dJBkUsJAwKaCSOiyiuJLBBBGazTEPzsUD0D0FVE/42mVQ1vz1osj/UQzFk/L+ScTmVS8
p50NcV/GTGixPRgyr6X5xfOSI38run8f0rl2UEkj/tj0Q08bI6JlovMzS18WcERVPbHj1jmnFTH9
p6Lcug40N/FVUkeWIm0C56+xDaDJq+GttqLsJUganhilBYo6PO/Y27BSjdCGsYHtgBfGQC2TOxXZ
DFCJ0VUlbj6qqeKBmFgYVtOcBAIahU23rJvFWJwMOguG/g9SFtjzQKJn8WmkCtslx4HVTfgNs2/z
yC0/m/zSyVGGG4IoGE877m2tOsBVZI431+d4MXrYjxD3wQMS9UNnjXGKNx7PBET2zwO9bZKcmAUu
So7T7V5bDm3i2rlX7AnnJRlmx+VTVDRt4WGUWEYUjxYTfuMc72Qxm0wzcbWOpu3nP4tl/37Y6zik
+5Ts3ajOp6OJ43oNu/fBOnQk5oVRniBEKCDUTy97Br6hwSO7OROz1iaa7Am60FttQ3uJ+UFwo8Yr
3O+gjmViJYXdRMeoHfG5Os5Gldyd/nvyeMpKMDcPI9m8zmJDfsZbDKnys8iUeeV18PKgL8cEIf59
L3w+Mf924AJohVnpcoGxn6pE2mVXJMOpq2xE1MeeC+gC+j/Ymz51Wug//q6MalzfbijVnvfDG3pA
umIQoZqLWqAxqmOsyCsCJsNCYl+lgBOIZvFliZWUXvFssCiRzJOv3k7UiIY4CpctDi1deha0YEU/
TwxWBaFJqX5uLPUTHufSixXuaQk/kpMUWCXIEFHggJpHorqANg8Mq91nk4/Yr0fiqhv+mDB4tHzU
gUWMchT0pp9sXRBODWSzNvwIRCqD8Jvs2I93FI8WRTLsQ8asw5CWfah/2DEwVJap7Xvy487J3Kgv
TbbLwfiR49QGCZQkFhxzRJW+Ue5ZI2LZ5eHCuI+qQdlNiW3vcYsvChRnxoOPY528EofLCZKBvDLM
hDgv9JpAJcXsQjIHTRNs0SdbVWSXvrq1f2dlBgP9UdiaEy0vnBSjyrTMQf65+ObBoGI/ppFBIWMI
FJqLZpwE6x5EMXRec4/hQwF20XpQimL5T3xi11aqbKwQ1iboKQ+pwx+cHRm2CUj/jSqVxuEsMJuj
7hTdZwoAUhP5SAJ3+NMTRWwmw203vfRywF0CijSRxtfFU0KLMsY7/CSTPHUJRGdlX+Exad9S/ee7
1WxlR38EK/XmPWbM+6cfrc+dXqBXxAR7u/63hzb8gFJmSAdVxYYKpTSMebmluC7GMSQtRF0DJutQ
tNnp6U9TSC3Fq38F3NiOVskfdXW0cNKp5aF9nOKL8zqo43ep1FMTuxZViH3U3z6Y1bKCjCO8Ywol
LEpRRpMo5I74dzwf97ZhNh4vrc0YeVxYe29rvcuxJRaXEnThFUz7CyEqxgnsk7j9tc++TDfdBq10
UQf7n9YKqsJesGTGHhAg33edJ3p8XT5eyBBdosklCWY9pZ5BNU2WE4qYXIEc6fg2JKMkeSBSBzy+
ZQAgT6qszuM5Du54/Sqw1l3na5O+LnVI24l6VYT5s0qIyHpruGqYQ10OFs68CysFdyBznTVgF27V
HY0dPZvvDwgMcfBltJexhxMBITCdY3RGc7mA22mHAMg+VXt9JkiMC3C4NG0imrD7vxACVkilvHan
3C7OPnYhVl+B5hwrIVaWGT5KjrTfoiJJuEMKw5kXFGGhozbXkhEAcADfOLvoY2b1+/OlzCVfch+q
wr2JruJCdC34pOQBfN2Jh4bNk9JlZsKho/7APTLb5HIN5aUFE1wXRvc39TZHuz7JkizP+igTzy18
VbP4uv2BBCQzYDrh/SKK81XiqahkPD/qzS8d3Cy4tsZXlDNiA4Mj2zjfd6oupLBpXi/bkJQBX7VU
1hKeY6ZJVXwOdtXO+BGjSWURXitHQj9vD7eReLLdyjqqEnn8+DI6sP6StLcamRE7ddsLxih6RFQo
qmrLG9pVdzvJvbgnPV+JD7S/XuHIHy6eXARsYesICV/cA1l9Q0G4kk9MymH8KwBu8UW+Y5NStu8S
Oezq89sSNtAx+Sg8TS9kXyRIhiDDs85xj5nDphS72MUO73Iz/Fcd8lPZ1BDknntlMKMCMu1N39o9
QRWcAQwf2GwEjYOstdKMWLBRqm5038KMGDUFOKgftMfcZjp/yKiBH4aop7BcVJ5TKG5T6kdn9x1m
pch0GqmlxAu7N++vsa06eJALQ8mDcdBtSCWLsUPBrAtvENcLWJOExefv/xxdaX38Jx6K7Em3JEo9
nQY6TsH/zWKbK46bApTFXb53QAJcIUIoUxFQpNsa6hxVYQ9yUNG0eL9rF1iSXOGf0G2u2VV/L53T
PENzP1sxZK9NP78s/ri5KsPPLnHf3AG4lggVbIt35MKp6rcyQiAuHNpZJIaPAo62S656hGWwNOZ0
CO3f3isOXMltAGTPxmp6e7aEBG2rnqIhjFMwI2AMnBKbnvGKZDBp956HvViIQ422+ycKV0VeN2Xe
OQuKsoeuTkC8p0hRPZQCETlWe7zlLZu7WbfyKv3BiULapgpxkBoQt/2by7O4zOS2+ahxxc2f/pzi
Q78t5NkJDSV3XBK/vDh7BM58ela9DzUSXvCYUYlN/vxhKKnWKEFtIKrKy6P0JoHK0gYIJfJNp9hC
Iv/ZfrS/fCzOirUs+EXLP2LZg/MQzQE2N2Kzp/ViiG4ZtXD4wAhhtZbX5Od1JZUHYXIHeEwfuzG7
foo6HS431ByPHmO+x3rwA1h5ui2yIOPOLwCeu8inU9dGXNvxGdJOejuVGJuQ0QayaIu99MA95D48
98fwcey7RCdxwAjEmaBWuzbtCPqVutDgu78xSbFwQ8cTSV4Rwn7hCuBrqCmi42HhzyN7OH6UAccN
yQVqPU7C6vwuQSJ0U9bxrCTQ8bGOhNyGZMRx4t4+E6cvRRkrhlzMm20ungNH9tzkeDfZoYBMyVDg
f5z76R2VU7tIbPZKvbeQdlkDNZNi/afYjXFKWo9wVhaci7TVHHwsNxzIZ5B/8PkI0jBiO/ffUtfo
0ggFyM8KwrWbAqzGPGoP9JdQJxZ9VCqYE9D5CfAja+Jp1AxrhHZIeGR29Rkhs38JdwC0KN53gmcH
TOY1LQ1i9fKv0RhKp218nsCZQPkdGY+w5Olcmw6Zn+ks/jMy9SMKQIOtZUMr7444Kg+fNzkLr4LV
OPkcIgEZ2QLETFp0k2WJvUWaWJUSjONn9SGAmleLIhqMaBhOhKNPN4kuKNwjU3f+XPZG5yLUH9Wc
7BOlT6SolG1nl7eAWvXNqsLba3yeQ9aYQXlba3QQPe/QXgMBOHg/JT2OWktSZLrSoIjYFKoLN0y7
ua+ouAXj9ohU9YO5CYVPtQFNIfemerEqYLNiWDBZvrEpXfyH5yxmpqciHyznhqEwY1mSmunjhuxT
YBBmVJUQHFUD7gVEUs2xwPxAiCpxiz3AmDPtMxseJmcTwNadEcAP83HHVpT0ADDyrcTNrZ8YWqjm
1q+c0dDOdzuE9OTdPO3wqXjLljZvf6hPKXOO6Z+KxnzLmvNkv2lu6VDmO2GMt4sxyCvxSrLYCMAd
DMan3rVmRlQnij/PCi+vNwnya7S5wS/ISzswh9XeyQn54MG6FS1d/OXeX3SUFWcdYx+wKPAlZgvI
8G+YIFyTT3/mvFmjq8d0dFOVGJurt7boUjscKdMaS9XL4x8Mc/sQ6dta0/NBPTBJbTDCbu8Gxvdv
23wEKBDbimLRQ6A9HF94yF7dZvbypth6eVk1VgQxMVBR0MH/hGswIw4tB6sxs22a8Ml9RjbrvMvR
K8DnrP8rHVvGhtRIUqv1vQZOj/eMeretG584T2eHVWYuhuQDBSc/dzakJ5DxLVWMUOU6CWC21PZa
TuuzuA9EeCM/l6chSLtSILpBol+hDluKjF/XLEoe21/AFVbjjAnT9+ZNl5UmcAff9t2AWTRz4uYL
Xpek7mt6I3sKjeNBB/pWP6CUi1O4tTvNXIPy2ftRZCs2wwg2AsIXPi/v9GkRaVltogh+BheAd1yF
8w5/SMVcnhWoB9a8di6rsSrM9o0IXbwQv19iySmY4sVw7sqsI+sUlBGPPcbrdalhMxtLKfHC8sJP
heZ04ATIh2PzXReen7XF0UmEVWqo8WKsy0DNk3jqdlBlcC/LLJPkQL3Wf48tg/DELK6ndlkOrU7c
qTmZs3lbeoQ+zKy1NGGJlPbvWhrVApXIz42sZil9L4DaTBfOJ2AOrc5bFdktbOWf/FOmqdFa3LBH
Wf7bWa8zMBUnhF53xpr0l9YuxskUpSCeUUetw3tbP9Nuf4NzJj5C/aJhl8w2gd3ZdMaI0J+xryxt
aYhu8ZTmjekV+KFQbkhANDbKlUbXjhd0OMRnTgbhH8XUjvMqgNHBdKTmJATeRojDEzOGTSk1jUS1
KBMVjKvInOROjE6ZCxZgHOweO/gCD5BW91Mv5tWum3Iheki/dslT3gWMfxYQcJFewiSGuAfgr0fl
j32BDpYiESaXMXNspPVBHN9Sx05gLnJowm9CC24Uw6PfasRJvaNwpwSyOcKK0ythN8NPwchk4Lrw
epUTFYOnn4Xq2xPOG4p0B4LvQ5dFlFRjrUpSCryRq3xHh37hdSgyJBSbRT6aTZUCn9YSKWRpB+Yn
HpoNtEncbiY1il90qgVZn9hIFUpuFE9t/npvQZ6T0LfGrQP3GXeqBjPJuQNe5TZh/eZeGHnddf/B
UI+f9RcR1MPRmlqYUV4g9eV0HgoITvoAQMKTmJE20n0qJNQdc3NbUACu7CNRSZpt/x2yfGJkOk8i
17LYVAtbLIg2wQGI5gRHvfHp8Ks997e3JWoRYeWIgG/E/UwFW0wmfw6x8RRbgvni2ew4ge4GyxsW
5dpajqIm8TtoLJTOrDFurt7EHOJ91BZQ7sohnOj2f7Ky/xc3GWMsCkZkZZKJ1J0sMo9W3eimtXkM
zh7yVMswoFtfyMOFhCVuMzh/MJ/aihevr8w/HTZicTp1jZYa+G756IHvMxAb3wZ8vGAPP6NW2tq5
35U8QmCqrkHuvPPNav/IifLFzRx9xmOR1+NsHQyeoYtYhmZWqzaVtoBEodVbpsQHOW2yrUiaKayL
ku7YjTmN+Azdv940douM7z7jE+rKbqFXMqSqP0V/NdsL4NtncJKX3aEBdSg3Of5aWGGCLQs7m5Au
IafoWJ9VcIwUVP7gdSGoY9kIvQDE3TPLBhGnu7mmb+NwO24UNLEpdPNB2NxTwhZd79kATIw8V1Dq
2Dya2ZgawTeooMMXXSCoQpZK/dfa3udPxzCSEG+SWHrdW9bwthB/y3zfkW3m/0H794D6gnPPxt5t
sbPrK9S6tHj23PhS876gsKBdDWPcWMdQ6eH8E5DsKDEpopbvxNlkeQDxfJv/7Sr4Q+DqIDam+I/S
JCD0GWCwDi9J7zKzBg3GOBIOn7+xfrwPZKiu5Q7EYyPGcoaz4MqSGRRAjHAyFL1g71jJheed570q
XgyaVQMnbmtiDdxn1U98FM5tyaJWGVDYSxx8HwC7hON1+prQmOUCDbSuPPb3JERlL+lA3O9SAC24
jfcov38En3Ze2wdqfBIUlchjcc/hNmBiLlz3QEWZQpLu34aBszBqZlmxNW/4iKnv1gx2iC306nN1
hP9MmNvqBcBLoDMdNV6t3PcWI3P0Qmm1f85skkhbjemV/cYQAYzCQDA0hk/tilSRgbH372nNh34H
LEDwekZ/KQMMGXVzON1ogfEkYE/6I7fkC2lum9P6Gwwy/j2+W0pl8zudBaifXWCJHX9s8mQT8tcy
bd9S4R32YSZxeiRLVN0t/5XCvR5wbDX1cpu6OT1rxXaH0eQYluqDc5TS1H0ikHCOGj7p97zJUG5s
t06jHlPUm1FEPESyr2ViF9POdU2gU/GikrguRSBnEXHam+wDXsm9MBGFyw/ey3DFW5vdOXqm4u+s
PK6E7OFoWUgeYyF1WaONGhQPUbtto79W3aYMd+H1Dxbdlh4+4S8ycs8k/REUr44OII6edOwS7xQn
txozT/k8ZQpDxnYizphUO0wGyeeyb5Hu4+WPwo2TtOLkl6BYh7e8EBlwRevEYgxwa+ijUsxJUu6G
NdVBsRjfc+dLlgOHQYn/U2wxU/Q6wFfKGC4SPf/dH1yyeF09axuu0b56hiAZD+3LxhJ/s0UmRVUA
T46v578ppxBhByCW8yj5prFW2YpyHxvAprdcmp/zKXjUDX3kvNSC8HpyGJ1T1XW8PZVtkKM0nip8
w1FL+jjxnmxNYFBkXpbo9ViUTgXUDD2p5VvMy3a5m2O4FiBnbyjUPif8EL4EvO4NBX1tpbFEHHlS
aYk/ncYTsI1XdIVwxmfuHPqfttfFcf3xqaWJuHQM6GA3OUyBYsLgrSGMrnzYQzF4qSJE3aCCgGk9
NtPSvLPjqfFyDn+f5QapTsXdxEnNq+C9qID6rxkn7SmznMomMGx3biPfPSUf7tTPe29HqKiswmIN
eGn6TeYsawFE8v6ELGUOsKGNRbnwxZ4Oz1d4Ol8Mn+1YYAFP9UePnmXsu7/QaklCBFZR75NFKo/k
Wd4F6ZWqj2xH3FLxId39K4tphHnaMAFrfIM3O/4O5tQvKHX0TWX9J6lKHEkgWXy9ZikXaBjTbME/
X6uj+FiC5dtSNqYBNpiBpVnvV2LF7RH7XoB8QzyISHFUz+16NH9nvOy23NkMCiCnQxntn4QBxOwB
P4BUu3jiUu2fIVRkoKJ85q0OWTE/0fhGW9r1AmYhi1jSqNdREzctwo0BByetespr7v9vckO4PLiI
2yftmvN+j3k+mMWUK5Um4YK5bECT6a7V4KN/nPTvMP8GEz/dJdZ0Uev3c6+kXDt80ckZT2ppYcdA
rvnZZvFGGWH7A7YNqW21kJrOrbiD6XtHHX9/Dqa/X2Hu3B6es4ALsjcaN2or/1JKjai61K7KLODh
rHXUp3vnRnNeuhq2oeuQkqqBkYARbzPF5riwr3i3oHTbLNkTJW5PovU30BWEmLsUXw+TFewPrnGL
E3Ekxci5RxdxKRoAHTcoBFOHFP+9bl0O9waTq/1q4Rpp6TKY0mFTdWDq+EnN8AcAmHnARd8SPWoH
xsY+fVNmiWs6IQNzPjEVPtQH5BOyPMRrEE/usRBtSxDjNg5XCfDQrb905zAsmXCtTiHWyoTM5sht
8VCulr0rawKkMVDAt5bjxWPrusrwR79FYZG37nMdYMARoifZS1IAJwVjrLbLKzvcCqAWjVmxpwj8
HinHBWv14ugDII5ZsITi226Cl0qNXR4z8DwharhcCos9Bo0J6/4EuMVRA85f/Ak7Nj4spB9jiYEy
QpnDYi1yQgFKLhzAv2MyDGmmOahc3XEfNJLvl5yak+8AeDpUxm3m3iDhA9v2PLJ+qDRC/ODEAYtP
R+vpQjtcZ2lMcnJXEnLQupbGi3aUtj8Hmdu9Lf0vnPiv+gW2QEkbFO1NLBwBG5MuSp7XH3dnaDDV
u05jJovtek3f1y5X/k0L9COu7I0/PMuqUks26dca3gc+/GlFnDbeS2gMeFdI9+SQssAqgex00Amf
72bcaSvztHpqNAZ8CC+U+Ob1FOnrH/IbCDo5vooir4wyVWuysvK+pNYoI2LqLxOc/h8smnRnd6Ce
P+Rx+w9DcmgOKVDj8G9I3TrCQ95t35LBM0/K1sh/g8klZk5Q045h5W/yFkLZDp+EAa3L+pRFZHZx
74jnyvrMYV2e2TwNcgEYX3IlA4+qoNkxWZDSF+2RCAwK2DVGZncLosNhVV+/xrMJT97yX7hAtEJu
pQdIny1+LRKOxXlwwQAIwNzK9acvod5pfIjQ6qnVo3kYMw6iyqUvucd6Mdj5pvMEOvXynGJsOFsp
qYlwn41/VBNIToXaV4cl3UVdqf7Axs8YyYhfYIeZAn7Hktv4oIuEJ64EUM5REIr7pRS9TwYkxNdX
VmaAJgpbua0XeDDGLqV3EcDjo4CCqFmaQ9ii/mzcjovMo0I+37pJxAgUQKGHcQaVfGjV05o2gMLQ
XBg8p+MnTMgwyAJD3Q1dfdzmA5HESogYnHT8UeIzSV8+nebtiQmoEILQsEkKrRQbFwqbrHTpnQFN
0nFCGQsDuVQvL3arXBnXGjRlC6BXEt86T0YLyJ3nigWL0b0b7UNk9ZzEGtWQ6BrnNIsyFqdDrd1g
u+LBBX3Q7WSFoVjucVbDfozfyaGH9eIYYtY6jP/Z8kxRrL5P2T1sHksHJze7NgWZzFVljOt2l9/v
LL1lcvrlN3UXfs8DeF9/2ghW0w/CofY4FvBcsZrASzf0ofDY7j6jgBmGW2DpbhQlAqGo/o3k3KK/
+7wi7gwd+9ebVezaEVrGtTRo7gBg6FXTfJppQfNFZpa0wBE4+dVbdqSmFiHCk+crxx91OmkjFs4H
fB4lx1eyqc1edV7KyMhemyjN4UbhgllTAgVWyRu2QndVyYpzLjPtUnqBBSPPp3JkLWxKVW/Rtsqd
wB3srXusTkGCPX5eHKt6o5rVFwca+LXPjtI+GOhepjGurPr1uA3XSVbx76DA8EYg5P9kKbv7kjq8
znx4rU9pC2YQf49MHgJpPJHt0Qk5ViknO95cM7aC+aRPx3k91LLW99YR9qIdqmanscs0RnJVpA8g
67H0eiHd7mJlb3z/C1mAOtkyEj+iG4sHs/ZeZ4FhYYyLdIS2HyhOC/jmqCngkDr+ARgKjvEyl6GI
5UrHaksfKnIQLXsA7dugz+V1F6MVAv/cHlPb8oMMTvg8876hp9clCv0it8Ul81kqejbUjJKXXJYu
dFYTC4mMsI4TMoGLsMD29wfkr+UfsUZG6qGLvhhE1GOeuoOrZ/br0dvcY2ctKCfKvAgZ3OFVrihU
/khuBp7u+Wn811+7anT5c+BnFuc0xJAXPFuX6hrMuo2hB614izOzoiYAYAwRVBxpjnR7PMqf1Ora
wJ8vzniV2jfddxVi/tqULFTMsR/gBo+0UEod3wk2px3ugWfY+ZqY4bj9vZva15MCoal3Sc5Cl3rY
oWuuOJbYaKzuOerIbqliC9gWYc5lw6/11O+tOIpb7Bba88Hopa7R33f0ErPzrmJyv7cvIYVtIGJf
UfJH23JtEf2t4CrPKiogZQTQ0bHDcEV4QHBfNvzqVFE+Dx/Si81vh2dvrfsxjXbed4Ir2roWSb6W
UGoDwnhWxXpWXKZS3hGBT8ja1aPyI3g5xdrA0fxLJq8HME3pGY4onCON+Bq/ZcQhFRA3lggrUhEd
RSiMc34tnrN15evyiLFAp2SC6y+7k9s4ik/h0yKEg3o3UJ3NAz4mE1l7iF5kw2o8KZSgIf/BxYNL
oX2sOyW1e6Q2XpiI/Ps31P5i5KraeKDJNZsOQ/iwqdd14RLRxVtVr0i00OOu6ibmaSIbIBO0INI/
1K63INIVze1LMvaqReOAkfHlW2OjMuxM3G6AkJnwlzg4RLfcZHImegJBJ3fgT9YVGKUW1IX4cdxf
nEXhNIP3aRhyCiEL2NqA6oeQWm8vkYqD0AK2s6OfSWmPMZf/hgIZcJdaVXBc/ON5X/A/uFQ0kNc7
MvsmFkyZQd4cFPkWtkcVFrCCC7a7vTmxWu49L2J/WUsBw/uBGDnWtbSLCnzOOBpmDqNDgaqrozNS
A2DxsWJfsRJD6XDmoq8N/8gFqYTTvefd3vVR9WLE7NabDC/Kn+T4DnpsNGH0yLGc3FETYktaZDuz
HM2z1EdQtHwSqHtukVMt9mr7TAJeti7oNAXYuH0b8qDV8JzhwUj1CWVV9/yq41P1DSuuMUwhuMUF
b3i4VeYkenT8E/82/uquZaBPSc3gxBBUHXwStUH8dZmsgGIFQeCzZ8ZappN598D6A/Cf8kHoZwT/
kpJAEiQiE/rzJgPjieR8HnJ/VN98Cy06TmILjZeL/UIcC7KFS6HR4/VzvAQmGuWCzyMLN4haUOwT
L+75BiOhGB240lleCalcE5SR9HP71nYGO3IIq0UG61CsUbn8oVBUsGuUpRMQniMOwcqj8ShVO6ub
8+VvVRIa71Y6JdP2R6Myy0oa0O34GwRK6sBa5ouN9wHIdZ7voOmONI95/BidRTKbM4D2KO21orNL
AKQSepAU5uXEu+5dJJECXee+oxp2y7GRLP1YvSpx7EDmnnjuNVHqZYmW+mv7oIwty9X+8LygWjDE
VA1Wt12qWyjz1ftY1JnMl+zk92/KLXga3WokDCBYjbiwwjhiB4EmS7FcfvT9ZvmCm8NtQVh2mqge
qbgc5Wmdk5S7xCq+ee2BZ39wOVf8V1883HfLtHAztVcQ2a04Vfo5J3iX9lwIBdnhl6HWvJZIXjH0
Yj5S1BYRor6dQiTP+esv4M5CbKaX3sH6RImhyqQzXEUWwFvms54rpjhX8dd1ue5Vy6djrohMyI8M
NDZowwnHxrfceBZLYiUUoUw3uosaYZ5h1sSZsGdZbjA7eF6JdFIP3hA6eT7slgGtUD0wrAYQa3Ds
RW1G/q8miKAl3Et3OS1caj1NsbU6SE5IwzvSgijUIF/fMu5pNeye3sdFrBPPMollF49F88X3+WZ1
4n3Q056jogovs8W8EwAT/mW9ALS1S+ZHXzOtg0r+OaNQmR7FkI8gkyA+UHiCZU7xvnw14A4UVvyx
hTP/gRfFXu8FY4jSAjQrs+yQ4ViB/BuYA2UNtE88Nq2PY/6kFjaJNeY6EQ6OM0GNiuAUGaXtZhWf
BZZ8UOJiKAv5CFO/F3/11JH4C9es4qF96iHVQMDUjbsF6Of4XK/L3VmBZL0attSVn7Pg6arsrO/J
Ax2MMxLEsKAX7FPBYaVgS0npI25AEGSq26ceyQMY8TFfdeJ0RKYFHOdOiC47GUGTg53rgeTRgvw/
VYXa3pEl0jIA+u73FOHPLpl9FYAcBw18Qz2HFWUFKbaj5BhQ0XdJXRPwVni2swy1oz/xnGFtogMG
V0yVbXPy5IurF/n+t7oMFqUKeF9YgCiEvVg9pow8qZOYraVD4aUDmphoJw/2Xr1E+gW9NSd1YepG
V9x4bnp6OuZdmmTW94VjzeRdTMomC4Zv1U683NbDD+rSoYT3vXGRhbK6CHkln5B5IMrndcKpR4kh
TP+MuUaLvboE74yKLaw+uS9w6R69Ct5PYPeVnQypwM7yEqwP0c0AVA7sxpLfH3SXoiSh21rXGPOi
YDLBTk5fMzHpNBvlL6UJlRVVhtT591SIAAI6xTIUypdkBbuivsG2IECLfoXRDhCGZ1yA50qXRg3x
Bzw+oqeutFRKU0Lr+UgL/UOFmWp2yhHqaOTpXgt111JJsDWmXqXjCycl2NeiS5HVu0VMTgjkNHG6
RXonaaGi2Tjd02hPdhCA2UmUe6xWYmr1ja6QtWsAtakNgNTJkIQvlUMmSryHLJhZCmEgU0/TR60z
r8YZ1VUCv4asP0gmN0dbxv4PIyPmlmN5UotYAnAehgSTKxlORW48JzWkpyQDraghJq1pOeFV/CEN
R/GCMzqVpnC27iRWY6euKLs/jPWburfVvD1QAGZ7tzMCUQbXaEmRvbGQmKmbxtWrvewFtKFv8pa4
et4MuWQoZDwen2iq1+n/ewDLSb7vsNNRI726XFnsp/ky/XsEGWkNY0nkO0KweZyZxC6butL+pGco
CUb+VgClSDu0FHG+7gPuC3kxqPyE1jVTnmM7NJmumnOEqHqPgOZe1oHrrwfvK21XrXuDZFz66gkI
OKiJ2vFqdgB7+Az5XCjJY9lN7lI77TuvyG1tDaldA5jxA7DvkbAGkSqpN0qVJVROsgw7I+67Cuoq
FIpw/iw92rF8rGLecjj2F5ETR5ePv9zCPVRb9Tc6T6ICwv3mKYYveQbjCIqU59Fv/1hSnEcCL/PR
pgBT8m6KjE9D6HbngZMgTDCTRY2d6OTqFRL/tX7BPOfJp1i2hw7kWwRUAKEspimU51BWAvWQK35C
XTMEvFQfRqSEiE401LTCm1dc4e84t1UFl342E5grDHT+Qo/LecGgIGjKhX20uK46dcKfSCXI1rmC
OB58xt2jNl8X5Fe45eKAMr9WXdnAbuhz/UyPd79aR4AAqJSh1sTpfBFrgDYux0xsJLGDcK02fd1M
X+vsD+oR2E1xCVuCStjqFz5oydUfDgYs7WlHKpheImjO3JpaAg3I0oGI5mCJn8i4n0Df81aT6328
dAvJ4lHwh/5n1CaodTibJiCJYBINcsrfU4ZHtOwMmUUSrwN79R4Zdw+z7fP1it1t+PSQ0LygFSGg
mxoCIIgPcSrP5rw0o2y7JBD0oNBs9NGFJZSliL19hk6bvPpklSLiToolNYN1tIelhA4d/GS3Tt6x
C5xdZO8xE4SjlCTlm8PDJS+kdZfgRlOjmNm0kdOA5zZZOti2p1L0QK7J5nzxzdqM1eUdyz+sBP9D
BAgIoGdrsgRsBYZYv9NQyBY6RNRsX2/z+xWmMgdbd6uKy0q2wjzyw3sbxuZCAuUHHH3wc6JM3mM2
Yl0+/49ZW3tt1hP5ovGNt6ryHKHn3sNBfph/zon/fZbB0/V+aNtBmxXkXo0JCWH0B+dbdLripJYn
BComqRar088eZ5I2nQhjLVYKVV+70aebO/PkIUFfpj5kv+KgDbftFNVRv/ggPf8LzH32VfjrB88S
QAwe4HrhAJAo9D+yn9mREjgJbKcL8AJDFG1kYrxltDRcH/MtpnNcHCKWlRKCOwxkk/0946XCpX9+
xesrkU4cjVJMvKnpD6rm/l+xdY2nwrFyvXrjYoOtSk8OYAZ29vNtHhdeBY4jRTHmOczWW8tvA6Ux
Xow5zSGrnWyFbg72Gm0K1Yz0Gy/vjV9gduXGrxiN/5AVbye4oZ9V0YMizDIeTs67xsqHvvUEjTX4
15pUF5vJRDPrxA8v356n59vkL5Ne0GtKU26LtB3PbF9LU5NGhm+pp9rwczUHJJy0U2PKoR/4IMhQ
/EFsI2IbkcuadpMWq/PyE870LsQwBI2zHhF3jQmcBXC5tCZyFAqWRWt9Urw5Isv+ip8SYTMIchL3
n0xeZxHpUFfmmw3HXOyfICC4LL0HmM7drWBl8lxBLWMbiojMp/HZpj//nDqYk+omR5gN/xXHBUoV
bRYT/a/Bfw6o8CSTSZyBMzoBLEAXZUGAPKpJRnZ7do9fAVWOTt8q5VFzstJMSTeCefBQaNreaFcE
SaSUeuWx07hNKtyUXcyA51E3PXqEQpolMMVpL/KraBihcUcEsVHJ9JDDnV1Q85VZeu9owojfZh9u
UY+yjttzXwAfz9swOVgyS0HLWIeKy8QFgHdJWawLBYOqd4LszwpS+iYvwvNxxTmVfob9UF8hh84W
mnSP91l2whKHdSiu1m2SuYBzeTxZHE26wJ5hsSNpowX8ojPraMIZb+L0QHtNAuUFcGV1oG8vqOOZ
D5GClhmoKzbJZPl8mAsF+AAV0katR/uQ+Xjxu+bd9zaWHn8ReSfblvO8WuZTJ8K6mfM0U9pbJXM8
D1382VMJtnhKd5CzXM8QuC4L1x3jWvLtC8ebfv1PE0bgQdfFhZti1Nm3xctzOlI5SomXfA2gTxhm
WXiwRRUmpekJvT51QEMzmY9flBY0m/6G5mlVOg+3SmOAUb5/ddBURIO/Wq4I9jIqeINBgSihoyZi
LiBgeNZoUWy9rQ/eEI/Fj35klOf+trP5BvyJMT/iQPGhPb9UiPBSJjIIZ+yEK+RkxmWzkUJCRikj
N3JrRbHt1wSWdzRC2HsVny3l+F4qf7AOOIucHawlAgpkHzRsZqDnbXSh9kBMjFlXqbMgU2fDDx/7
a8nAnd7X1PjTXTZtQSlzCPmroLPoeUJ5ZqF84P9K56dT8t0XHl8z2XG4xp1j7Zv/zSvxl28akblY
uuFF5LDq3IUbt2fzYpwOt21omzbhfT//KSD1602AE9ucXi2xSRk+FXfxRgrgXnE3rRLMT9F6JWF2
TtHEjKHVzB63uDpnH76j0SCI5qQI6lUwR/uj2HQgEeoZWcAfKPOnklbnjP5hyfBdYTBrmgk3a3IU
6KTSOJgs3BRa7RFQmJyaomuEu3D2VPzekUWAibVMvybZ+6OEaK8rd+pocrPoaomvAvpxlJTjTJPL
05RU0NFucPTF6VjGR9hlEb2B5AWoTtdrW9aj4/8hUKvgkrUzLkH7PJV8yJ/2uBBQRmWMGb3O8KU/
5jQdVUcytVLJIzWygWBsAh0mRnGW8YBFhOYHpheB8/yWgbhpeo4iIRmAkL3Pu8lyLlbYqtcGS7zt
HwSjCu090y9Zg2+LomQ9LbOyNYNj1afz9VTyFGuv2F9EIr38rY/BKsdXhX2UonQBNnLwkp1/t7gX
BSnmdMmUeeei7BLgEfdmrr4eldpkQz+1Gz9V1AlRCnoP4E6jlujaPkgNfUyRgvisJOQ6m63c+7rn
lSobSMV7tryVJ55MuMOVUnRkKZFGxYKB1ACL/2FSuoXeLIbbdcs00tFfY4PB7/BFKJFxX7R74KST
qJfcnkXV83rt7zQrmOBO5QFntOPNkR4yuofGuvVpCix6KQkhTNSHUz+e9W3r7WxFF01EMkQXNbBT
UVtC05WgYpptqRVNU+jgn3oLyI+xZp7w7+uDm3pmUG7f87AG47ShR8jz0jV6EhXpx4PJE6/VQC5g
y4NUnQzOsbg5/f/TvIq0Mv0Srv8WsuEnujz/MWVbMA83GvBY0qfXRiZB14TrLMLjtnA173ED6Zlw
6Ip70yy0+QT1f9XgO3CdlVLZ3hcAP2/hgBLq16uRVJJK7LKbMABiyKpNXNgrgMhTtkVnzpHBBvNj
WaMEr1FREJmHpWuo9puWOuB3wOPxccgvEfymHvzG+yvceBeESey6xpqFcrsgSO13wqF1v+ol5wFn
tVzfkJxekvVjwwaDbHZ48MvZu0t6cTqwMaYGldhPZWgDUIdQoUTQeFhfWySIerc2YUXPqE0wRLUl
C90ceCoxaVZICkcidVpNiZUSNcooSC30C75pdXgd+T6ql/oh/w/bTOJ0bAoioX8lcpwnZjknnzQj
9AlMH6UBW+X6i4phrzhRYazmJde9U38eJmKBhSe/zBFQbAjDQqMSR47MVzsFh6LpNskHDXpT/VR3
btE5SuvZzPQ2fTFuUPR4Sv7zPF8xrFQ1bZPrbdqq1p4oIOYAzaUYoqQtbEclmf+nqx38OazkpVF+
iDWwscvTzGC+wucQaQ64wAdNNYOPxANUd/brk0HaLsAR+5/rK2rwuZ+/ee2yUvj6zPqsuWs0wy+n
bJQlU8RyJWq/VzLMrPSxrMO+ZdZaEHuB3anEKhZgBPXlM2+gtS5kkH17+ATAaFKJ1rJvvm1frt6Z
EENhbuSv5K55DBxxUGBaKBULtG0lTvWaxRL06z5Z8eJqOdS5fXRHglrHBQPe/3haqtoTo7Hi7Pfc
BKKyiKPYWR57rBx1OSsRZ5OXxyh7+01iVOxY4+YzQlj426voqaHmns47HsLi28DI/L+xqZMDLbsM
2xDH0TOh+XOQP1Kr+nGVowPYzw7kjuj3TMTe+qg7DLhpM3oCEkRMs2uME791yX8IpzoxMYFWGPtC
xb5yFC+5vDUZXkGydleCmBgkIB7QVwMs2h4pkSOGLyoq2bW5ZJigE/hzX6HQhdwSuChpnV8p/at5
gy4gOkqQTmUiQPhJQuoI9JiHOguMQaKJiahktxdGRtpc9V+HSpV8dQGJAAZgY6Kvwkn9+TP06CKj
cG1oJC9sOOvuNz0Z6Y7eGOqGzitf8dFbkdVnD5SN329T1UmNgZRfRfLWTtCQBIPe2Zz20tulJgas
4SVjEInhw3XddOmzjqaxMlZEO8FrybmNsB88ybS94ZNhSX1RZoQFzvmOtqL0JBfns781LPgKyKbg
XEzbAYn8yeXb+CgT2ndk0uKACvYHA4uOH2OjHyYgxqGM9Nhkr5geGqFczBwKd5/USfKf+UvfiafW
de73lZY5ZWpA4V5AG5GJbddL+yDH/vP3LKVSKQfUYjxaXhFfJxb0SCq/aLK6ssR80Bu3GcLyr9WM
dAXLMy8nIVIh+ijVxDuAclw7PGfT6lLFIUd0qt1QFyUsoa4eriFEr+BfLSJTXlkgKZFmtia7HRXK
GksRPEGGI/OyjM3wt15GKvOtlP3pYuPtxTT8FrHjSTcv4QCQPbr9jzdDcsVvW6e/eNxHxRtH0DCZ
HfuWj9Np4HPLgr3EMxscslbQUXEIhGcSkN39tOHYmAvPWH21k5Lg9bCS+AXqXI7VzNG8nkpRHvAg
4zl1n6vFlpu4XBAOTHppdRdPssTfIPTWXhUKYdD18YRVGIlphpco3/k1yVjOQ2vz73CFqZwlHqZu
AGiD5j4CIJi/iBskZLbDE//qUnIhWR7eTGjB4Kl/TQ0JLKLhZj73nlJuVZYeq8WWat4G+JIJu0/G
qaHI3SHm536VeQp7/yPKaUIMgnPNJcy22PZII18Hzr3g4p24Gu6Q3SpG8p0f3rqk5b8Hcij0iEik
1wXZZXGTA/w4qbsCTPg059TVlCmJy1LqkehdSF53rGso+VgFGP8/bi0fTAefv3BhtVTv0VV5EVjP
YMH0rXcGYjLLb+JpkGnpJfGdXSEbAuxK8fDIlQcao9+fc2Hbco+DA5fNv2vs+qOg+PwdW1vXaAhh
5R7r3hglVWrxWFnVR5/9H73GdKAb9+687o9e434niJqoF/LM63vVSEmQgKb4zdHHAtey9t4WF49Z
IhfIyBY43s8wzLnljPCj1lHgH081FdHi3DB11jcfi61gJ9OyHIGrv/RzPomQUDXZrMJ1YHO1Yn36
o8D3JpMnHi8y/Dky7q0tQR5V12JbXf7qw+axwhGyyZfqJZNUXWxc7uaaQULow/cnqPZ7O7MWzy2V
nPNdE+yGY2GaCznbw3UOprLrfrU3vfVEp+6LsH+ney5ZLKAf9wDgissMuyDLVO3uTi+7u/CztSNy
UTHSL0LITNkilLOU3R+Bz0DkqWbgkokXb1xSwVCTTOGQBj3KXo6WOGbYBR2WXkYNrxg8F5QTpCwL
9RL7ArhA4m3ZN1JDj4EGCxks5WgM4CYsZNJwZa1QxoBS37r3LAuA4SfPhOBnPW47J7Z7YaW7waEs
40cWgifyoCXHGKX+G2r1RMepVTs0KjrdqLjk1MO4FP2/9EIH5srgtoYBA0cNI9gpPnl4S2imHJba
tOoa4CFFlt2Tgy7ncuVxATtnWukAP/stYDdNMKPBw4/y6JXwCEUYU75kXd2Q4rcF53NN66DDrbgH
+oLFMp9kt7j5XutCjnaS8Q5UJl5488mZa25VlMjqf89YFSmooRYA69+FAMDqnt9fxtiAlUw6xBz+
RFtqivpH/+C1Iu7NVAHoJWgo/F4eDKqkKH+kZlqwzkTU0MM6eBYVpb/0esa8E/8XvvApw7cgdeiJ
1SB8xV9Om+tTqSP/G5Lzyq83R7lQ2iXv2psYhdbdXZLapVLB7f81Faf1o8lplw+ivqvsfmRbjEr3
AyQVSwRhuhYvMD/FknMpmKdPtbGCNxqteiXtllnzIppdvpjLDMcXjUAwqkS3+5GpWWxgmV4TStOO
AyTijut+c7VUyObnYy9guK2EYAvA1HW6jDff33+ibg2aYF4Uj+xIu/HVhHe0fkBL3R0gbDYtRZER
YoiT/RWJJYngpmzy0aON4KWDiqtl8iT0zUjHmov45W0sjtZIlz/HsuBgyQyHozhDcobB9BrfFb9v
Ds6Uxfw7ErEFKjB8BsDki5NqejK0rhYf33fqFgx2QK821wBo1Kd03lbWTAfE6DvBgrtxj6vA8vNt
iPO8jqJW+fNdVUX+xTa9yhSka1HP9hxF+4vf7qHh6rsKjZJ+LCm0+oJpcrKD0yBw/CquELuyZUB+
J27yftpOGFA/mDB29vufbtfyDGPBdA3M1JIbTH/bIm2ptZJzjxF7zPDn+LChgnETkpnGuZoouFjG
5ePyvrEXEl6hA4Wp47ToMfXEaq2roN1m0/Acel3vo49GJhnFHH204f8ekd3wvKOvpmoG6+jo7u63
OqnWQ5LwrUjpCd4Wq8VmeI1Ewk76lNkTjCoqPu4pj49PCalaFUEt1Gz7lBXXPMCbGwGqwK0Qr2Ov
1fMl6x3MZWHJTMT5nO1yXCfxQ6Fqo29vUUIJNN8x0nnf2JZvUI1N7IlJ15xejHBBvWNnMeAL0xYt
pEfDfOw/foIdpSpfDxq4UdWrdNPq6o5l/R8Mi/zf1cKTXDgroyMTdsFDNCMZNXcZ2SsB3eX1hcCb
D/oR6OnuhIEQUhkPMHy8PASn2A/9NwFPXTtA04LDYCbJKIqEiB/OR5MH+w2cHizhTnIkDYja7ciq
ezq6y2sjZ8Iz8AHYQwK44VFbJGRteUVhymjsMHkDQctR4Hpx1UIbEZ5nnC1ueZK9X4GS0UDoZjc5
9Bp9jB8p5HNIE16TJeoPETbvzAcZQ7mEyAn82yBCB6ljFMS2Ck4f0a5DEcOP2+CivtBZ3SW+rmgq
8ISCTAHW1RRH2Zs/nHsckWInsITKF5od3kc2OJh3hqgsj3UloORalLI/4I+9n2KcO8Hz0E8+sfnn
qEOLsLciU+5r6BIxLQur8L0BBdKJZ6K6+lCOP7H8Y2MSZ6Guw7qKqkuIeOoKVtfGerwPuNiA0SgU
VEoDAEe/H6s8/YMMfb6WKJS8I0BhMohkoCXgaoEUm8LcsT6TZ7zkO4yvwLZcPCP/KyMypd09xmw8
1rpQbdkgrC/ZQGku1YJQQah5ijDiuUE5h98/BHphlNmDPajZ9vOcGlj54QHJjQyLJgPzfxZUyMB9
xw0RY1vN9HJ8reJ+Omo14Sn7ENXpkKK0vHUtimeBr8XCPz4XUzEi2YX+nXTMlkvbwE7xB2w7eN5o
z4wrwFV8HTuf3s40fAL1zACnsOhpundrufhhgsIVB2VR3N2bU3RgqVvjNFWqfgd4H09J6y5lOW1q
pemfHVa0dp5+mVtoQCWNmZ6NlhHSCgYUWywBf5ZQJTcNrpx3l/shy6UTbUhnM6GEOi4bKRoHGl48
dTTsIPdhFWm0M0EirycPup6b3CzVF3vBpWtp2XZEdAgQ7f15IN8zD57lvKjwJKeE5bI5Yj/vrIbQ
NF9NYRs/2GaGsrzJ6kTnVnAtWjI8E/35UN4tj9t2vJ7c0ZCOJxlgHcDy6HPM015zPxZGdPhincth
PPNFhePmk01WKPQKRVbDINyo9mfEVdA8H3XapJw1k5N+tb0KW5ZjbRlEhLGzsOapzdbCmIXNEjq7
AhnF+wSUc7a7slv4PIrFttPsLPaoYjE3Dw1YSMdZEegUl3aCSz6TtWclHmg0ebUW+ymqVxlwS04T
kI9TRgoeLCljl2amxuBXCRai+j+ndpAS72kaGBwdNOQRnOB6VIDH616sD9VDM1t89MfD90kM09o6
C9d7TUwCbhK5LkLv6N5q+ZGx9hBuBBE3RFysYMs1L+7rzVcDbzNUk1pqf06b5+yGYAzbmwN4go+V
UrPCwwsmptSZ4VLdjN8G+pSAaUXZ414g9otes3fqh6l4Mw+3ujSsMINP7lxNyqOgU8UuziKh9QcX
N5/dF61lfJ3DCEpMF5/afkQUZUJAt5bvV2x5/mh8Ok8prdkfb0slCWlk3Jymqyb7NYTEqGpWqGmH
qqKMxayMaN5Vtzpjz5RWYHDVPMGV/xiIJyiwNHltE1KUPKa7ygtBuBpoZai5jbLYjK90k7PcaXmn
0OfMkv6PB25MHTef1veqfURHyw2W1+lFDFa69epU88czeMXAyJaI4yqfB7YIeNySGm8Nxat6SHby
PXeGl9rRzsdo9OXIK7/z+rhqTntb0IbEUlOG70zmStZ6H8XBxJquOuZ+V33tcDGmW0mcTVE/+Gwx
LdfV7VoaL3DfnixHXuSCyBBp8SJB16F778KZb44mNqpl95/uM8E+PP2jSVNWP2B5628kD2yyIpeI
bxx4cuNvDpzSJtvus7sAtKrwcYrbya/S0B0HPlpK7G+5ra8JHz2WJFlzlycRiwl+2wIEzXTz38MM
jxED1k3QWWaavgzushhsw9ds43E+tEvK3f1yNs9WmtuTyZLaPoyU4oscgRs68mvDo5Q++2f/kcEn
umarUKgrSgFPSbcQr6QFv6gMDHmwc4Idxy6n12fp7taJeLcA8RLNezs/0UuXKxYIEC2YoXUFkA5q
FLyPHBV6g9OHulUc3ItubRJw8pZvc5hkLHW5GSY0NxuGPRCEGdF5up5BFXzpsf3T4hxdB1SrSGyu
wpBrxVszo6DQzXIYlLjzcwWauig9fCrVK8O2S6RDruzspesVSpbqGOd2LUgsEGYytII6L62aaqZ1
86bsjYL/gcydATjJathtMsm8fMt8iJPkhlPUwY/pYk/Ad/3Pf59EECaM2sHoZ8rxokzAs7T7Qe+2
eQuqfOStTQQZSv2px6RGFCWxY1egAQAeQTb59vRqIfkGk5mVUL+WcR9SJD05qVVhJzjo0uJ/V2lk
nMX2xkwxLYeWGjAr+06B5ZOm13RTQQ5zKmmZjYJ7qY3FzzDxvIp7I8wvPJSH0sgjMe3Pg14RKLbg
5XViTMWQecotCabg0Sws5qQVPNPuQUFuLK+IHrXBVrkRbHodY6b28+5q4yMjhdL8Q7kawOhE6+FY
d5f4By7BOaa3RSkbn+Q+nv0JAVwzm7Cm4lbm97mP8eQ2eu6ZWrCo0Z4P9HHbkwLABY20Ou6S/oas
/qbUfikFDizvu/GEyt30uTZ0oL0otBbxJ7QeNKrTV44FmQJSP50qXpTprsrd7ZhS89+iZ07w67jU
YDNcYvXE1JdYpRg9eIVnL+GdUFWDIllF6IMJ2nSyPhyduyQryP2Eg4Zgnw1Q0juOYP4Tr5j4y0qH
MEHNa4sC1H476EiMlE40pma2i4ROhZiBHFPBdUBFGdfQWEA9b5Oxtb8p5gxi2k0YeAm1mLDQbvmc
D00f68b2equx8OwMpxNq/NocYj2a38quTGFEStbmiWiNkzKbE9dt0Mkn4w2VL4ZT7ZHgcNyMmX0Y
l2+AxocxuLAnXt9Zuu4VXdKeyY6k1J432O+a0cDYHjkgH8u3XFIzTm9pzEYUgm9TxcuSSMeSih/8
0sY/ORDvzUarWySSIThlpGH+a0qMWrJbCTn+X4xMJu15yEZdwcKUbDDJiZkqp5NEvWQWmmkLYWLC
nd/lC+bCAugY2L/xRV4zArP65vuMpWDPNhonJ4FNKbtqcDQh59+WtslETj2kaZCec/4U2JbIWMyZ
OIXzahWXdceNgxk3AM58hjoSej96unOD7Rs6+4cgQ6lowPORYGt6L08wsU4n/YTybIgficXarveS
Ouymi0RBB7rpAr0oBWY2iocillZn/8Oehhd0uD0BiyvZxC5at+/GC8cIlDOLK41YsATSoY3n8FOK
0WuYfTiAnkp9R9Th7FMAUvg9o9hxNuC7O7Go24O0Q7KDwMaD2mweCqoTZAJnuUeSE9j1W7Wu/23m
NuvfieL4ahVKlHh73tN80Q/nAcofrFi8puorCYEixXNmCYODHz3lsP5WQCfANmF9W3EuPX8jil44
75JmYLCo0vFQ2hPtjPtKYXcgBUW5YDPl0X3gfnzPKXiC7PY9OK6Gu1tkmirRPrJlJh1LbRZpPA5k
os3S8nQjMyTcI8Rkckioi16nf531TJ/m/Oh1L4KCr41tZLpCJRQEbogDmQPNhiGhue3UJqVZEayl
fiCVk5f4e/XVqhlSF6wCcWZPj6loRrSCITbvh9Eu2WMq4Y+IjYx5LOBUVgM80g/zkM/cSS+tbvG/
7krJDnQFN3LE0DpdEVqhE24ADO74arZt+TopbY3O+cC+aW3DylGi1mvjf3wbUnGJIwx1laAaQRUG
JNl7Vp7nwPhUb1Gxug4tQKg4UAukCM13k+iH5xI1fz5t1f8bGgOvBdGyIvEemu/y4U3sa7XfEqwl
vgVa8VVKdxPenpGQSR4YyqPCaisTFoVE3PeKwmVHbCHaJXPj0Kxb8Q5G7GBJ3rTEXsAsbfiJPxF6
2rZomMWkrHQ1SbI93PEnh/hJmOM6SHqWhb1a6U0l2tZFfMnAJW7prihcpY5dzME4XavrWuPXwWv1
wcbQggeLIZYywXeEAXmpDt5wUmQ53tOwXNuTlIbTufSbFFehkjTe9LxKvbP9pEVG8czhOx2kA1cq
+72cKl+64281dfTSdDztYbDSLqPhgpTettqkEVTPnBcV66B2xPAUougDeacrZ4Kds2n6zxM691Z9
KjobDcE77xHbfMTmisTJlP19yov8EKKzynlnpuVKgZgG1cLiSkAIqUNJhz4h2k6d695DGuBbdRSy
VoDZzYQKb2NcwAHrhNA510Ktvbhc638QJTRhQ6J96KFs0YrhfrF8dZs/SsqDA7S9VMvou70iO8Is
f2x/z/t8HTUH9U2c5K3nb0rZb1iiwUyqoyYtmrQ3T24nqHmMVC5NKo7A7Tvl2f3k+/bto1G1FohT
T0fImkbvzJY8NFQB1ddGCb685FIPmrEGqCXqEJlJdGIX5lZIJqq7dCf2lZNKHelZXG9d99hd7miG
PPqz21KFuTcUcH/574jTRPBTryJ//DdX54fPDfBSVT7fQqYLR8mB6rzMADGdTgXd7SAbb27BD5on
7Jr1G6Cssb12epc9WS7MBrJzuK32lp2Bc/Y1rxMlnLhtnLqSjwrVw6h0k/LG+rzyeKrasgIelh4B
zotUERkqONlweIYq3iqk8IxrDefOxoRFr+qC9jPx+p5nQVwgGNlikn+qMTPhf9XW7STQJgpXGUqG
Q2PIBPk+5GeThcRHqNwHctsPeUahodFbgRfKuzAFu6pDtPNjPPuFbcc3+w6r4dUSBfJ2eboATafE
0V7XPp1a6DlNQ1ogtuvLCyqOoHhebr3wIXGBPpXx+1S8KVc3yHAN6zEbZ9uRsj37Pf5GIRzGu9FL
bDIA3tBS2R1t1TEepYPKE4J2R0qNK6BGVgbLcFgICmnHHCs0rvAbY1guj7b6FvaSCOZZXA+wvuK7
AGskBPZ6HL1mKTj04gyTfWEt4e0rxCvrVTrZzQiMVPVVckdgdRuTmXVay4K7q+oOqdkcuuk74J5W
BAHivTHZPAVsDsEmd0uXjnDWQ/5WUYtslCgTvuEQXCBHRKhsaMhEoD3O9oGVI62CHxoOD7A8Yhor
2xSfYBAXX/rBrN1pEMggzjzKYth7Sri8mmUTyucFuCShOkDTKtd0D+Q3WFCn/pOtoUjYRoDUdhVc
uCZRs29JYZZJbWkw3nXS9wg4MRKm8Xx0DfOsghoVNO+4r8aQQUPXZOQSGfOksLKGMjN7Zt6orPtR
sjRdjSAa0E/2PEAYDXLlsrepNAHXptkM1sl+e2t9mA+e0CsTdAXYnKK88lmbm39t8qhTPWY7gKLU
VOMVLputfYiGdzi+X8jCH7qrxEee03mO5CUi/UnrYsTaXzNPSuCKXWEHWnRdix+As7QBrrBSZDQd
BqlixPWJ/YSH1yeZI45ScyvQqkLUP7Q44mKvMnREM8VHbRQPxDffKRa/ivQ8O9luK+8Qn8ADYYhw
6D8FNwxivFyOAml/fWWb27+uqHuZkFR0Zc37QUCSePRX8S1UfFYaJzex7saMuMLyJklNf+7gOc5i
BFuO9t0I3vyp4Bz6wHjvOTZq9Fi1kpOA11cbRs8spWSlD9LIrH/0BvRt81/EQBu1y85YcoYnGpTw
vz3FD/nD+GfheLPmi6aT5UjG5yFqnFiZjB8k57m+diowQOa85zrIwgPe9pNbSg/tx5EPHDQORd09
NF2qiEvqMRYBEoWwK6qAFGAYtAzEc1LbjXK7qn39c9rZdoIHjXM25zY9k2y/uo/gZSIr7Vu+wWnX
b7lIt+2kipNlC4xD2Vzqbgw5m4Zg9WlBOBoGHBba5RIdKRcWU/SDRp0/IVN+QN4FlGHm5z0dRP9o
6NIY8zwxij7N7vmpjIAIBOLMFcjqeIBFs7cPBrLM1Py7Kuihwz9Uc2ryuIWRu2ie58YTcJm73VsH
pq/a2dgvrI/ZbMG6tUxchOCKGvij0X4TuCeN6sSbQucwaUIMRhnD2PQNonwvxg3p4ai/fMsFKWfQ
FoWg7ztRtHjDZlCgyIJph5FknvudRtP8Ww99C7VVlCbnOwwkXxYE0m0MNn8s7EFkW8/DA6/bfPc9
Bdj1j34J6fbLEQnsR0fj74s+juEkaa+rbOSH0tLhwinXrgW6nRRSsfdf+r7FaPEErX0wdZbqEAvZ
N9ejrfHl1DJR2ap0E27p03qZOBqRIMdezCtDqp5kCxuo77M85I4jgKvjOn324F1bBxc0US85WOE0
vooSiRzHitz9j0MPZIqL0eex63ZnH3e0NQcuLEAP4lVDKwVBvINKPI9NsfrzVsdmTs/jdLI3/kDL
QSensn0hyXwAH2V9Svz1tHQWs2qHdZe81tOLaA9hJ8N0rmeTmit16Zz61dfRfZC8LEciRGPpvI/R
w94EA8AS1IfroS7InDpT9AwM6vORhQReZYSOQaENfXCTxDz+ofIK+cimbA7wx1DJF5I1YDLqtbxT
LqQzOz0l95RMzA0CY36T+uIvXvltiM5LB3Ql6DFwxZnz6IxbLCbznM85nupVdBusynd4ZLgPXsvA
2LSqLRHOEbPnFGpu6Vqs1odKiK7pec5YIZ0z2cZQsJmZsV1CticoH8FzDpK/OgkbcF1GFGtR9Pk4
/RHSaZBilDIo9A4Tq8cObG9WcGBLn6YVaJn3LxRjtJw++6onXKOlfZRPmLjl14WbIDdws8vFUlI8
6V+TTv/a41k7dHC9KF4DowEqN19d6wbbdimYD0oqNKsq23rNhKktV0KGsuxTjtD3v4UQtcahfVce
QMmBzT/1ElY/mQjFx2bgYqR1R1befqESvX+Uhg/AU+H+MKdO2AjEw/zSDklLfPbXBvdw69stVqc2
zkPQUE1EcLWoqfVNWWFYA37Le7OLeo5IY5P2hXo1cR41u5Ibj4vDv9JaTeEaHLaJj0gjAk9qWbEr
VW809TJx7eXSLZCI/mGkSBj368gYqoUpu+EAvbVD4KgJl7rbw7EccrhiMvC1LeKR0XCEQmnvo7rc
WDcb8aTOGm8vDuoWW3OwRb6M9DZMsiRc8PoXW0WyzIzFrN+4NsZfd5fDEGFJ80ve0E6J3jUNJ4dt
fLVZaxCT4NRUnOEt1+5EKOufiwYb6RZ2ijgvRnWSoDJU8FXv1oDcqYf0eGfV84OFShdOwMGc+SPL
c3jT9nfo9yMnCkJeRCL35iNC9+X9CIH30pSPZLpcKS2jjLgqXoBXKfcfr6t4qqibUGzFduxxIh2B
drlTVmAVKx2pHO0HKdmr9MefmfElCS9IIpq5shB7mBgsZnuBMCjDuTTcLvQFVUJ3C+IoIVIvUWWx
mLhDZGN6Lhp2YIrytXT8T6bItXNFsD9jAXfh1yhCMYYgfWddJDuTBtjrLIkZEam00QMVFACfW9/z
R5pOevfEiQGbfN/PFg8nnSKoygSG+Qhi/9AiQBzlZEbdQuOd2bo8HsYSf4MAsyAAYsjTJeuQuWUB
HNz/VRX3fbGD/0PeUQ9t8AqB+o2kee+TT9Rrcf7vaCoByyE3dFHkbY6YwZ4YGL9L1zPOL4Ajy7Oz
nZwSvai+dymm32UCNAsYuC6aUKeP5dFzKBT0WPE9f/JYNeZrmLXWHZcPw682W98nJk/y71Vu7skD
IlfAV6hPrgHDe2owP/r8i8oKnv/s3GfiBqJ89wU7PsE0QmsCzUnbxHl04/coDVkVoWOobsiKe9RM
uXcVFX6qeSA6scb7HcO2Cw1Z8L9Y+MqkBiwgHNcFoB0zp8oVEwVcvuRI7MM9WO9OO6j70YhXGlgL
l3VLoYcX5iCEdNuy3sMh6RbZvuBYhxj5SJfgwiFSU7NZ6Z5TfNB0gylarYHyRDg8sS1Rxc/DAldN
0h5W5OHn8RNbr2ajXpnoQW0HTKcKhvMhVNTjcnHz3U3H99GGLsTAUt/L8iZyFbEGCDaAusnADUx7
S3pIGgXqbx/gKpAcnJkBcQekhfpA+X0Nxfvr2W29mq8vkyuy0eXgoTSVj+l/+4wU5hFHVq8S/gfk
VXVX02hZk5ANyclL3y44rPo2WkoVKzZOsZsS997Y96Pme9dqDLWr3mEMfXel/j0PCBvgKELlxN9d
hQnM4CuQ4lXgJFFpzg4K/2IKbuqOflLKhsF60kOr8ARFs3VyeEwbUgPJLU35ZR/6XcspDXxFJbt7
rZuPwycQ4bVfppdIdiFWh3KrzeHWCJdm79bRCqmSUESwn7awpjfuek943R8Bqebmk0BvNTmCcOhG
t7qAJPBo4hsVs6cxc4j6ztDzTiiJ+PKZ2hl/oANo5GNp73i7m45m6rKW013KnTaPIULMyOtFPsBh
36dri832WEzZvMeNIi08AiQJSxjwW1FryanKOU/M+n2R2l8rYkogX2s2Ck6ywFnQ9mG5vP+nuXR7
A3ifvmcjsDtcoPBMudUoL6SORXf9bQ64avzEkfnZGxdUIllF4S0VnSemJKH/Ec9PDDegPyF5uH2E
vTYd3t9ksqsrXoFV5SMnIG3u1WMDYCmwJexmvmfEMjoHDXMIL392dCs7oPdX0DkOix646BtY0Hst
GCpVZth274qyf7h9WJU/unrGvXvk36Bpl/wd0F5hMX5n1liQGQO/DRNxuknB58tYAWmkLBZhBdzV
fncfoQ9dRb4QSjmMg8vYIW4XeyLkhINaL6AYBckCjmYCmgEf71lgVFwkK/ajKZXCv0u/Ua314Qbw
LDObtNkYJGFGRnouW5El7zI7i3I5vS6o6yWyJv6kHeKf3ctq2ZOBiJ5PjB0Ebqsf9jpcXAlWvwHZ
8zkJI9IOJYXytrjzu/lob6Cz82JOAx+5K0XfpQvH3y6W3CuO7gGIR0U/W78M01lV7Cvmw4fY92CY
Q+1vyIEoXBsKtnMi/IdqLInx3DjzkkxkQRgkWCrSTih8/DBSl7y5BMUygL+APEXT+Wi0gb35RT/L
OaJfmV6RUkjEKSyB1ajTgKUoPIfi8YtWCzTrjMfYyxmQThQs6PsnqulI1dK3cGeUUbU9H4VD6Gop
QgOkQG9KD667QbS54KH0rkBIiAAxxM+peTp2UidG9QZ2Gg58PZC5JEIxDLCtjjLFRcIEsTEgcBiT
0KhXGct439+P1fmViIbB1jMISE6Uhx5uJrhz8gel8/Dg9E3YJMgS08pnEeW5xaMUxqQWR9U4E7TG
wFeIo26Xl4NzUgKtKa8NDS8cJIapH/kI2edDoreDuYS1s/1oSUOFOGdT3ZKKaSLAtKKafFJMPVGf
4bKHrxUIYtVEEACFDAj7fswfA1+UcghHOGUtW0sfj0GYigN7NgpiMYaBLrDhMG6Gvm9z6XOsfmTy
eCzmseFP9HZeHNT+uelIXZuGgQRrHXfiEeF/f0f6mUYOkShgDV/XUN1eAECYI8NkbtJJAGnOJu/v
EgpW2SKNFSKUMTZkEAoh4zNoznJf1KA3fvnYK3WKh8PytjnSaqYmzY+fzyt0QUAe1JUxJ50scUUO
1esQ88BF3BTr4gCJVp2QDAuAme3PhzRTi1BOEbjRQi1kAqtpP2hkvdxp1oDNmudKGUIHJAbXkr1d
Y2Jme8xPI4c5DdCfUsa+s9cODgcvn1KLfnNZ1wCNYJAD9mmb3b4jT3ox89oU4OcXireeWUgCBkZo
o+bBevprvp6TEYXflU6B97XSghIsJ+2D0JNzDh2Vb7QvXKN5qpCcTsrh0igQDGajckMCNZQxgwKt
FF80mD39u+ZBxe5rC0oCGudoVTC9M9H883+O+FziwgLKPW2cKT8tsJEpDghtyk8XiwIt8TAqdlOX
Yu+rCFUC7ViIO55pOX3I3xZAltwGktpu8+He0NYrhS3NPNtLWPTIX2YF3bhHZbmSiAL40KBbRvt6
kUSw7Fvb365vbWERaxYeU78Lm2vbjXAYiGqV9snECxSe6LuwNIYvdygHUKoaE762Wh5LoOB8mANi
IvCrVWGLq2K/vnLUujkAKH3DEZWYvEfSHsRtOZjAOixKvCjRPfttjCxA3LZQTVk/VOz6jsTApNlH
QjNQFa/rOofCKaFhJlvBVCPEkpryxBpZT0dTdgcCqlj6JNPJfBG9EfvwtMavYuygYhaFPmhXDct6
P/1XJ2k5BB6gk6urdoT6oIA6nKAyFbSAwKhKFjzStRA+MzMpAlAef//6swrIx67gciwyk4rmKnmj
/p8kX2ZRCj4qhd0jXzA3KLP6/u4YA92qbyn3ZXitDV4kxiya0XlhQzrELsIPxXMcjQS9v1nF9knf
IZOzDlEGoM/adPpc+c5lJ38/IWvHRT4qokX6Iq1zDuPbgAmJzhUHd6QGeDxQWbPb9U3+EKom6XJf
L+yV4FjN7+9JJIWe3PneI/LJhBN4TB9+cLoYbF/Q9PXL0Z8HwtqqagaUx/7KL9qV3erdHmHc+w1j
6aAz+tFwD6STTzRnjPCXc9clLfoG2rnNsNGQUeRNoR6QWEbS5huGlJvjFXAY5SbkFgQr3GJUhanB
zQS77tU9RTXULpXm8gQsQjYIX0BxTybjU24bBng2MRJ3n2xfDxloDdsel70wYq2fInDCcWEAIglt
ONvwXxxirZwFZ65NCBMGGA/EaV3CrmpvSjTK5Yt0FFQpxX1US7gg1djlCtdONQPm9IJdP7hNnxzL
7scfI/1MhP8pGlr8/L34snReJdNjrb2ntE41EqqdVvTSjq9LDJXa7FpGq7xv6ILjxhTLGWMrzyzi
dtEgbIsbyzT8mO+dgMSfSqJxqt9aTIms8OHUh2pOwYmpRb2QZPSzA9z5LsVMbyYZsV7HB1z975+1
o+6bb4ZA7ffngPBz8V0f5S/lBlnQwtDlnvaTQtt91tLM3Y12VJqAv23LaI0yURl+BoG9gh3SrpEo
KGLEOvr29Pti8GA3Q0Y8M64HdmsFo3YCYzNFLGDtcBlAZQTPAU+s8nlN/cKfSLz9EKVLqQp0QZe/
OskLe0fMMvT7r4RI1Gcq6xe3FUB8M2o29gG2y3r2AmBq/u7P+q5ANAeJ48tnfLkeSYHuAUEsJ1N/
/2KmuZh48PRh+CR35gBqqZoBB+eJjd26jOJaYuwjxQY+8iWz8pn873hGhMvgHSpyDDW/Z8cpjGgf
qKVh/8Nv1frs7FK0tHXxOhzf3aUPini4okufIBSzaKNk21rJPNkrZCj8szf/rN9mEhKGTeySxez/
eGw+63sTJR/Y4527LZVenDnWV6YlfuCvX4kLPB3XjUk5IURTWebMaUmQRD8VsUbZsRa+SeXfTA+U
xJrlA+UaMqIaonV5UgoYDry1WhEvjiMO3a6HgbRBljrp80fS7V9XrfYrwjPPvDf9Olm592xw/J6l
kIN15/hP15QTFbNg2uO61CrahzsLpF2ye/1sKoe16CYccyUypOzOURUqIF8SQF17jITcp0amrMye
NSSM+GbWTY0thdGL5FSLa6AmADTqVpKojlU3QYJmsj8usLkNYwxDL3m4+5o0pM2kaTWUaOqWR64Z
niWGPQudCaJtwJqMK74XhtLaQZXA6YR7Tr/JvBuvwEWDDhHsCr1fOIb4jRSH8wGMxMDUGfYsFuMi
Kzi5UjCOCWCqb+cR5/Bih0Jru2kw0E3azwjNhXbvICmVvbED8WeRD6DD0BwiRrH7DFhEZjrcSTYR
LoXQqBWtt1HufJ4lUAvVf5NQk730F6euLRZ8MkD7kzOyldEX54CCw9zUYxf85svH04F1RDq9xZPN
FSfgF3MQzaTP78UzK91YI9th8c+C+2zxGCUtCXOv86d6bH6dowc4UJK/s7PbJvy209Y4cXjzUDeG
XqGYSiVq/+WsAXysdeYBMIGC9++v+Bir+zRE6C/bmmdpYFYAFeH62Hfo0K5Oj8F5E8u6Ji1aK7/O
NBXpyxO7q2x0OWirwSWyQQAas2YCDBg0ICNfwwZfchFkVF7I3g7FxbgIY/rDnEXCzOf0+PV5P9hd
QCcs9xykegXLr5+51qS/kEBleZinObNhWz1V4B443WXRksMjI9E8OcUqwPnCDrC1LzN1ugWNnAxD
BWC+DGfOT8iiF0UiEwBIeQqFrWgT+aEnTWIQWjAmwTZIQeFDOyQExgphJXzf73c9Ob5Ji8hSctZV
WCA83AsCxwUcFmwnYLdXaatUk8AqVDIuyYpjdffGGNpnO3mm9ZAoCsID0dMEQrSUkWBtoepgnhH7
7QlRVCXx7E0gsJjTd1zjjBZt6rx6HMNu9S0b/fslkybmTsGVNGiOVhP+gI6a0rqWt9rQc7ZprUT7
wMuiJzvnt4UdZeExeGgULuRVgXBVw+wdpab+dq414NH25N60XWiCtpnsNfUYPGQZZXr5gcB6D+qm
KK1H0lrOk+onWS0/ClN+fTgBnbRB2qOQ2ZeVC/7ll8Sm6G4sJUzpaI7wZHW97mDpWrfQHLwEeLpd
zcw6mD6K8BVmqfAnOSjBd8rQd7JLr12jVt54Pkig3pt2ZnfHMYEzoCNP9mgsAs8T9sNFbi1qnLjD
mkHl39wRlAoBmRgm+VyQfvcTPG3kjXm8POQ/GuOgfH+b4n7tfDIi8J73Uqs3+Iuc3iWu9dKF/tLF
L3A4m67QMtXbHmOEqhHv/ILTHQug/ss8b4v28hTdXNSOuRA68B/SVa/Sf+DMp2UmVgfdYShy437i
kKiX+RsOxEHhhVh+czqk4JCx5btJWwEhugFoL5odMEAQ68CCvb1Eb0anu5xNr/j/zNCSZV16VuD+
olu8ywsobPnsHCYDaI5Taa2UCLCnmgvE2AMy4WSe5pmZGpQx63s2ZRoIJRIk9SNwzCeNyq7AFTG1
k052A9gw3Y2thjWNrzegAy0rO8ilpwsDLrzkEf2V3WM7QvN6yzuPyoe4FqTDOMrbXkC0njK2sQn4
NSxoQ/HHn2XHtoCX48Gi291iIuDe0mi4v4TyTSsUbU8gFSf2bEuG/OshrUzsXD5JIuW29rZO9Rkf
YABrdPVwG9KM48rozvH7v6kZ/lz01PUs5OF4Uyl42+aU9SW3+MtSs0lx0i5kiib2ZwXTfsp6uC4J
Da9lOkE0ryesATUsxgJXDgdVE3svzCaQZuYJ8lUIkaUxTMjrvJoWnQFqVq3mgX4sXvu1wsnEXsr6
W+U8Uz7Ms+tjj+XGswvJ6ZWXUiAGtWTExV18mbs/fq1SfKsXuhPCbeE4rgxqO78EbjJJZCgBPW3o
K4HWeoIFt2LL3TkfY5F/Gunc4Qj1fqSOwhC97lu1By2XbkGO5m+zpJSI+eCZ1rNTYullTvx+ziCX
Il/pmGYFw/ybKYkuSbh+XwtWC0kjXzNWL8N3jAzrNubpiFPE3j1UGqWwgIi7uQH6tWcWTSrgDopS
SORDc5IpMqY43GV9U18WYgeEpu2G2LkgYdzmSHNyX3cKXahqw0Pmb9OlmuX3bXMu1W1S5+/wYN8Q
V5LTutmnRvfaJCG1mekgEKqevfFW6SAUrojdWURbcXN+NgWcBGY03i238u+lMEsc7Rc9UD9TfcJJ
1cple/ThIU29NRx/kAKXqZ30FYAY+CacEUB3VAPALNXbpglRG2B3qMLGZuqC5hn6yCAJKELki2i8
wUaNes8VKTwziBT5SmmvBenSKlQWia6DzY1xwQHitgKJD8G88Ts+pd8qf6NeTFw45kr/Mj1b9Gyb
zdfMnYrMz5Dv9kzb0qtPj7kog+2z7W/P/SbwLxxKkOkwLFAvEtO2XWB9srI/XYgW/iMImJODeAy1
/79jJsP0P/JJRl1bElO1u/SgxfE8wtCazAmpQJOSYLpT+nAWMUOsEkMGZsn8cfTi6VVWDha0cjs1
yfVYtkJ2DDqb9lxqxzVGSFT6Y86TzwTBC7r1PpV3ueStS2b8TCrojmIUgetQtYZjK+t9wIjNLHa9
+DVJIyYcYxX/jxlq/6SwxH0NtUAfqCZEguxwSmeA0PuZX2bg30bbI8l8928c2TMgCjrmawwLuAw9
ECW83ljj1pSvG2SiPJzo3hhKuAcTH0JCVlTP4/Bf1L5EYYwLzaMeco7DHfxX1qBYznEouLrmbbJ4
DNnZEvTYEd9cLH4oLVldHlIKX20qSaXWNEbj5sZwHg1B7o1bLVvDT/tThFhPFnQynyDWJhZnJJS4
182CL3LeoSTE2St3s8TPcWYXa1h9jPvoC/TeVKAd1Fwx0MOqBl5WZZlX9O65p277OLheO72oUn0r
dcG5Qs0Az8FmDJd4YsACejRAdoTKm1VCkNBQIJeih/fMI7IlwfujnwzoT50OctVj3XCImVNbD9Ws
IRBX7CDOVIfm9Py+VLduQFtGo0G9Nh5XPok4ZPe4RzOcN28xGxxYFrGK5tutt+IPk1uM1dhyPKvy
6OA0IsxZa92ydFsAncOWI0Imn+4NV2lWv76Xz8tMS9PepThSlcLYDWJdkWjhJU9pbOy4abexSPhM
c084Th+78GcX8gJk760dl/x9vi3SaDbZo8ytHtl09tWPaQiyVJkY6X/b0F8olY6XyoaaI4VQgdrm
+lgBmISx8vgYaG/mVKsix9KNPv74HNCSaUbebNQgcA7RcN0z2swIk0/CBtBX6AkHodrFgC5D7lQ/
u9fobT1uKmwCBpHu1LfCfrgnS7fnvil4XycuU+0s0T8x4QKcPGUsUbKhh96wIiDG0VAeDQJ8hbG7
3DsCC3zUxSuLibjWC4LmrzPdcyANXmYCwqkv4qDEZeNtSIHN+fyHg8BTSluzbyCQAaicmIvRVr9q
tBWf9FsCDXyxTxkoFlsCs7sTIk2YQiGKaeAFmdMpU6qs/qEvawxremcXIbocetzRQoDBfZl0yhNR
sdJrsEoZ7+AM/MNTtZXROtn5ZEQt1MWSlYf/MO1xzvb9+WXwVgL3NRg24gih6qrDLcEdlz781RVe
8n2DzVbo6ghy7ltW6cX8sc0v5vpyRyi3305eDmvdEDLopjXtzhJ7nKaYHepS/ocnakHNlnDuwBsa
VUn/ZePWYfQDHbP0vwppCCvd5dP2FHhub/GitOuQj8Iq0GQcuhdDbUsYk5PdlxjlOBNjsfKbeqNt
ot+9aCDEijvDxtj69R9UbbiuQAjJozfUxxVB8fk1NahGFIF8CxiR7KiIzUuYnPTw9DZZC3gEv/gb
UgYKJSTzYV+3GgRcJHJarQ+BJhvBGtKb4wvs8LD/flAyyyMs6FKjtfn5jFdP/QsZCvQU7xOk4tnw
qhV8eJFS3qp/CHDUyLCK0clhy1Bulsko1jR0T0vLVV/6Kvjh5JidE5fVgw02b37M6ARCOX7Qapsy
haHGcS1KEUez/hdhYh6i0EYAx9Yfj1lJbiaDj/SGTs6PRVzrTH3stSlJARD4HCoFwynFkZsr2F5K
y2JkMmoeyG+l33DObU1gL/lsMNm7DdidPgpD1jc8D9TlUzLTtTb46PAloJH904Y4HpPKMMXw67HK
PuWfS2rMHqyvj1jIo54Kq28KRomOJHZp4M8ZfvOANt5KUk3PV+29NVxb7eFo3XlKW+36+tPV/RYw
ccssL9/fWkW+UGEAwL2AakzMGSEn0sApTBuiXJUEJg1SHr/JDqbNCJRhYZKD4rNMx2mFlzKTIbn4
RzejT8RRMGoV6Rz3QZXvrUp0BDXGGdbMgFKm1mhEOcbSpwHmtKWt8Tkz1+ykl0Y25a48rVhGl+GV
OxlQk6yTEOfXI7SQjbBLeAKxbY4vfeKT38UDaTIBtkll4jMYx72a6ioC4lthwfaZZJ4EpKi7oZ6S
Q8UayExOmr3Mcn+Qw6Gw4HTwSJaEECNjAPlmD8OtUtuCUt4ButjK4U6tdmQLp1lrERkgPyD9ep9x
zil5vVEZCz5uYVLKZQ1zFbJbIww8Opn2KNFsw+hrHV0kT98/w4rGE6Tycex0CC0gKgm28T4xBxio
2VjsUsw5Jz/YuXRo8Z1uKWqMfMlMo4ypMYTI4k12Re0Vb9vsL9XbwTCxFTbCyn1se1GQGvvJdzHT
cErj/wBXC202X+YqefqDCL2T80rKmqpEw1YklsmycdkKcd+G7AnFnGOIkPn3UQP1Up7SKqptaULw
7RBvapIGtn4ujzQOinlf6ajDrblhgKH5/iz4iKp55EYocSHselp2Ql/fqLPpKkSWGP4/CLFhexFh
3WzJcXg37DK1pPxYbMOhKo6NfGw/DuJauxqM4G4Du9WHhtqOWdNQtc+Bfx5uPM21FGofJY+mFq3R
gfR7fsbB8pbV4LejxQ45gtv9eOT62/c/0Gu0NS8Bm7xiyMujI2FnRM23LIm1GUjMWvAQ4Dx8XvYB
Aq63kIOiGuzHGSJgfhn1zhzJJsGcEQWL2v+6ifS9Ca35pKOLAzHrZ/5zajp3cxWCo79ctjvBiwN8
VwFoLmPA80C/MY0YwgIVQixRhHoZ9b1f2oAyFq+nSnU4/KNvIe+yF8LLJh0zlk7/eaplFowYQxfo
hk/y7NE9nv1Nu4ugjl0SooeTJKy+zHIhU4Yhkg1DyKRa9xJLZ2fuY+XHOytyflrc5919907UKALE
F3tJIWZkQpinACf5sff2FPibPd0iE8zmojjyXzeH8lLXo32xxMWTVWQ/c/7Dhql0NLnW5BMWQF2K
0Cp2CZzATzb8W7kMsXNEh+KSWDkHYaCBgPpL0s893fdNGo01j9+y4iVeGNQA+oIhOJ9759QGKGaz
jFameZxw2QFlGHIctBNxKnm4q/gqgmW4+HmnpbW0rwNQR988j3XZUM68IX5SQSkX1UTbK98gwz+b
NWxy2fM/nfxPc6qZ52se9m0NV1Wd4bXohdykWXshRzmmfY+qo2UkM8HCvyJ19lPM/YHnLdJm+OaO
AxmzQK7POvnpgrwh9VTIyIpWu5gVscf/EmF/Kp8rk6x5ABtfmQi+RWNkthzpBh5BtDcCUUXL+LpT
9aZYdrUfu0u6p+E9vYH5JUBrhyEHJCJlJCWHS3d+Kh1droY7M9wN/hBdzr3ZawdMJUR/b9z+3xUB
rJ8MMSuyZGFYzlg7M+zPKhr/Buk9PRBiX+U6T4Vuu7wVK0hWCg5wrgc7EDDlnFswuYhf88Rh/mDJ
gOPGj0UtY4+4jhTEd+lla66IT41ZOdS4MIV1Dxs64mj965q70oK8JmsnDXVA
`pragma protect end_protected
