/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 848)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAKw7bPg8uJ4cUDJQ+re6DaDmtVc57NyHbhGDnoz59L4ALdxqmNfPY/pj
qjky355QdDQ9Sox/8QhN4qS/ptN/wLacZFtJTvUZAoTYg8CD6pnKFWQ9DQDU+sJmG5vST5zPhKF6
0jEGt1MGBPsyhMU9WTKe08VCZp1Xbunwxjby8PVNFpSLNiu03t+UYZVrpH0Wr4joVbUCVKsN78uY
mQAiNZ6yAv3ZVMBGcU7FxLBw12dCHU5ppB26EmswN9PzW+yXeP/zO37rZWCQe1UGbg50nC5nydZg
k+gIBZbh4swx1VFPUveTPAmC23W8oUF5mEIPTSPLOlAhfMYlohGzZEjmUUBOc+5gU4t8XEyfrfXS
c8w4+08pEf3NqC++c2d11Qv2fcGQ+1o8b+Z9YIWrUB2m8yepnrmAIp0FUtLhP2DY9Xu/ehgajpXr
nAEyf7RP+SeEWTNdEdcpczwbHfbNaNBPW2DEmDRs0VTt7K5Qh2/5xT7xwvv87tO3Ngwjx50xPXmK
Byct4WSDoOCAGxtiXIISZPPsJDVOhpPRoRJbIk7ApSX0DHCjlqFfy4+P87bsfYP1cRyCUUfBCgSn
MQ5nHyauubHFZA7yWoudNs/L2s50cLluFg/Xki/FBFnwwwK7dsHxAdGcHtHGJ/HrzUN1ISVRvP+T
07aYF+FUwmcYUhBfmmPOYXyh2DQsiceiKsRetX5CXXQWXIu2agutbftxfvh8QTLP6XgOetRTBejI
gsjt5SVUb1QIYyePnHRQDbbdEwpYe6zMHeTBUlXQRUyn6iP7OmivYcWIRKKM/MMfa02tlfZ+3Zrq
BmJjSZOWtw+sKnaYV1KqZWmCZIZ3SPy+jAz3fGO6AoSYPG/xMXWVTEKk1lkcmgR1N0Z1Zga3KZku
hGMUHZCPPYSHVAw/F8qwt7eKVZXCoTpYnJioFWZWZt8OgfPml0FxqDE5DhdYwrzONOPdlD+ip4EK
k47AGdoMRzfvq83RXT1XflYsDJBUln66f6kfAKCCTfInT7r2aCG+vmwv4ejVly+kq6VK2cleybRw
u0ozWyaBbVeVDrvvDxqKhqnhijMdGPvMIxFkxttIXcwBJDqZzeBEo/0cfQJH6Lye6YU=
`pragma protect end_protected

// 
