`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+HL2qqGaxFmavb17XAoVq1038ZV
4IMcaU236hM1zTyd6WcW4g9OnGgqmwme+rjc/E04aXdpLViBO5twxX+5UZC2F/jZpxW8jaEShO+k
/Png3aYH7P41Emv18mR6+J735SuQU1J2J1FsXl1ITUWAeaWK6jEWiyI7nxDW5hJzJe2yZzfYOGGk
PfPhv4VJExchKK3KkVdQA1hEaACj2PFpuoi9QFxj6ziHmyTuk44b+VbB/TnRA1wCHy7xuzEaQLQw
WhPrrfsIJ45/FFbo37wZwEHBE+yc/DLHEr2ZwssnkUH/EKZQkUqca6n1SoibFBisP8hdihHO79dP
TbVL9aM9oikAlrMuyYLtwaFh2o09sn4jYhcuVgtr31qtN5bwTsYpWDhKINuym/j6fsA5IRqPO8ZQ
6af+4EOwyoD/KfsXKCCyeDd5yaQ3NjsJ6umd7GkTYNf9qdvdoZJZNzk1duHEczcrgX2XVHP6cmML
Ic1+8NnemtIQqrZ1k2861Ia6Zzgd2+rt5jszjBxOlZZ4G52qpSxIfYE9TF3EHZgz9GCh+4uCXa5z
4R6TV03EqtEjApD9gXNZqgWSLbKChXGht92dIBD8EecX4IQio1W+mLZXvj6ZdYbHoqervlqjPpW0
rScVnukE5beoT2Or7/2p6YaZrql2PiQYZq+9J0OafAySXApya8SR3L2svu/tuR/6LFpamae1cbBX
QAnjva3DYqfYEdf5i7hOAYoHigF14ltZZAD7P72h/eUL0SNr1a8bfkO8o6uPex23DhHmFCJb0DiH
0J6kkYWHhhCj+C8mGnffZRwgtsLVTXplbf4UZgXoZX/kYE+zu2Tl2RiX7760GU7K9MAAFzvWU94o
5ZQX4dp64kkZks1Ln5rBOLMxD9vUPCLCqtlyqr/neC4XZz6VEL5SIfAcB1Gyzdae227Hcpq0han9
1VssNqfcdA2MsxcIwWs1f+nVt7slPJ4GEsMt5jHgzXW6FEueanqvmtu2Hp7A9pVgIJIvOAWlm8hm
iZYYn6RwjlkdVHxdMyc2D1zoApLY0X6hdPZ9uB/cAKyOfeAMB/pdtfAH4N3ZGK9Zk32KkxhZCPdq
Xz7U0zkd02Q63chYRlhKzAwGmxtvyiMW/eHExGcALJqdBacetvDjDkKIBuO/o1bMEF+zpw1lYxTg
pcofURUgGVM5nYOpbYTlXbCt7owDPu73Yx+HDLwi779AgRLoCmnqRL1ITOoEOLIkl/jRMfqmcuH1
644aQ3YMI4gfWmsQ7nqC0UU5YGcSYBbKJlGGCd4a8EgCw2Fj5wORCUmpQ+gnfOwvms0Y/btYXQZ/
XHai/79WboRblmhtbiCdJVK+i5/me63Fb/DcdcYNLv2xThVKhhpwjwLTV/5Y/q24nOmKK/txIov2
msdxdfwpQGmT81k/tZnkidVr22xfBoOJfGtjUMzaiIRposkrc29awgtYwNWIOJD2TCfqogA6svv8
YN/Sz6kyyffWFzE+iyGMULPSdAvpkjPXLUcVPeCjIyJrXEFjHeDREFqK8nX1GiCew5pk4EyuPfpz
Hkfj6zwZNGRSQKAzjhpiqYk5sZWQF8HJbctFpyy2guWRv7FIF01AWGkxhrjXAUg0lJJMgw/E5vBv
1lMAUqkr5YitJF7srQ3bicUWM6254g5myQwyFVQE16ktmnL3pnfEwD/T7qGTTNJdEoRq8j6rhH+F
DA+kC3hbo3w/IqSx8OWmYEZTkmsthxpgVyIGQOo981zhCfmV36qwhapbDq7jiIS8J/YC5zQOqLfW
tRt78dscn2lGnvz/m/jGI+h8+ceY0xHZj4Um0fKFqDzXA5eLiYQsWCKTX3qDSBBgytjwoJWJvK4E
H+150A64VTXiEVBiujmw3IsduCsBhwtJJhYXXFcZ2kwpu+y2zpuBNO5KM9+70vJY2u5OGJkOlNpC
t21d2bnb2zxtATeD//9nKOH2q1UL/3lg270DrxOfabV+ZliLz8QSlNoFdOxMpeBztwESkAWhpS5E
gxaSEgicDjHaYoL9pW+GTXAI4xjFNx48HTgSv2AaYkrl0/lVvckZGm5yKl65o5n8ExQyLnlmZvmT
8gzMLB29t5wrzqXsoVklGEEGP/0Vldm3Lbl4gXMPsLnAETurVwjrFcWoaztIAjBWh0aJRopBMbX/
rZUAXhfBn6BHgUW6SSKwWFlKsq21fvwEHR94GXAeI8LZi19qYv/O9EpjlStuBGP92MlH/Q5Mzz1N
YDGqTl657XGfICjcT31aT6tqDVRmoszIWQBvx1l9JppmLyVStmER+yJEC05aH7rKF3HM2C0VbTXN
0MCKrAtdY6RWJcIDk+Yf2bIUddlXuU/udGn5wDrOky1Ig+MCg4azFVPQOvHn6ubqI7737He6z6BO
hGMvbl1OuuxCtj1Co+Ul7enFkeOKPUm7wGhjZvFkha2IzRRE682VZ+pu2F8oN2IYoJ31fTBabR0o
TKkcsuQgPVRbPg2cWs6wBv+fGPp8Q8hULNF9SNJd5W5a5RIjiBNmPhRjI0RRK3FgDhmOAULGMSXb
ny5SOkSwjgeSaYylnSQqxjA4HVphhHwbGjFBVNUz/3AgB3iirSW+1m9XjFVOUtcL+VJ7uA3VSE9W
bDjhb6FSPGu0dVOevusAIdoFc9/DzzLbu17EMD5JjPm3prF8enJ040vpcFsIGIV8Ut573DeVT4GC
s01umR3gexZ4UVP3a9Tar5ZM4jJ3qyHy3V+Ssf38nvKurdSoXS+OZfQcB1oFHwU0N+/PHh8O7Xe+
O1pZUXum5bSUN7mmtXuuDCbtzxekzwnTlO/TwNxrvTwKNx6eJLKua3Xo7J8Hkzrcj+kcn7PnMr5V
mvQdwP+7n4EpkzYeCcryIPEg9vd2ve8rSv+9xJVr4SXQR1ywi56d6oOvKJ+eaNE+QHyzMj/Elu9X
WfvrYpZSMvWUpo1L7wwb4eHaChCZCk3e4nLQ6CN4yfjiNGaKmXYDvVky+6jXXkt2EmTgvRPGozFV
w0Gm/d65pZZ5PzxztXi3TMBeWjvkh2+NN1STqg9HkQ5xFo1ryfG5N/3yboupTJP87zfCMzXyxecu
DtzSzTZN5nzQhFVHxmXgJHiW0kl1oJAU0nle2m80ffMnCDeCYMlaplos3NRgLIOOPUFNmx/mphh8
T1GX7qRmO2HKQrho7/CUhcLTm+oikYhEUQuw3D5lfSRmCeT2lM0wq3ACgMNA6EdOIqv3vRELCUI9
ZMurZniKnUobkwrRPn5Pxts6zkvNiaZ9XqhsfoZV5pr4CjR/DIHzrlvP2BEb3F/PADYkILypXIeP
5JUMxzHozlIybfsxmtWVNEku/P128gm+cbWH0UFtVBoBfCajpq8VcxQd4yjhako/ghz9aN1k0ffP
ivxEOVwH+CUD9b1KYll0rkZY3MgMzhe/aLgx2Dy8w/DvYIENcWtd8NdgcFBrAv7hWivsCIoN7GwS
sLXHJVGaMRQZMJ/gtJgMJ2h35OGrruOdEe72Gum9jTdySJnLWRilZMzdMWzvpNUlLdfvMmmtaEli
aCLh0YAvDNdCZoZTatZEHYDJI071SUDYr4M1HHQeAfN+5xP/7CPSorl0OXmJaN035+MnjsV5IDqD
v1c9N6ip0xWgO3pLV1Lruel0lofpgK+eIgefqKN6ZPO2lGHrlubVDQ1n2nzO4lEJgdpJcPDoj4ou
TaPB+4VdE6sYvVFiGCQBbd5CdGh3FHSTtG7JvJWoJIAH5JC9KneQnOrX4ZFcs6EmjNZvTIby6gWs
83/yOAyUohRDSPSj58zqQ9bH8SBZfx6cQoJcOdGGmGi7pSCwUYDdFipxPP0CamUB40h5A0HWU/nG
UcK3tFwWTbharyphlT5TsXNWvbcBufIoIV+JcYaAUz6LC+7Ox/SDrOrBfFWMc/luAImp7l3e6xR7
+rXE1TJ6Ft7bfWChZvmBkJOgrwVQqKfFlY+8oVD+nnU/aCJ3g4DqNm7cvSzN4xVvSGbAxbmkTLQ1
VaNAuEKZ1rpv8cuht656nkWQo6UcdiQvxdjMhQYXrPmsDAZy7EYA/5fUtf15tBAqCdSVgSLBHjwR
Q0NUYVYenpNz8kNQlwMv+/PT2LawWq/G6wzPdn8HB7ng2d7IMyYF9YMDN7zPCu9Ucb1ZplGnlMgD
11VGQQcVAQ86EPa/On4ZdieoLTA+HrzstYaW6PjMuXdNnXElZ8CDQeaF3yMih4GfuJCWCSewP7Q4
qUurbekxAtxwl6cMcgikROrtIiZqzk+pki2vrHc5CRlCcQOnEUdbxaXf1beO7n9xCHF7/ZH02jLu
PBTbHhjBv3wL+MJiF9GKOBYdEWSloEnwXoJWEofKU3/rQLPaTawc91jG8ivXgfP/f9ge/61NfzBw
UrcuvIq13nDH9kaqN4hZ35+80L4iKyU9S10J8qKj2msRKx1uKss3mBmX/D+I06Z8uDxF4I6Gv2vW
pikhjXLSQpxO5iHXiIqjCcJ0LssMdqOWU86ibhicConumHYF62WBZ4Q3gmQlLECfI9FavYr5HgHc
HSooxgvoOw9t4F9uv2jkorH7azcWC5ahb4+Fksv8tqk3TpyZVO0dIx8lVF5bVgTHGnSjOndJa06N
qfAYV2aonp28hbV2llSjGrq/vuDAsS7omWEUmV5TOTXblbCzDsMj1dFj296WH0k+9rTc3MJiXW2E
PWNVgsCcXYyGWwplRqFIj4Gh0WAP3pnudfjpP2NlxOuA0k66bj3AD7CIc/gqhJZJfvZpHvlQr1gt
6a7llk32iHA1jUWfn27kKB6V32leTDfsFYP5R8ZEKlqvnqn7GA8ODBnLBL2bdsHNpV9Y7EL9iHH1
RHx8gzMOInQllrLw4Q6jzRJk73RHB5/PUWP/dYHwQ7WK8x+vm1YNzlfEHgGXz2MoIlxchIhj5Wy5
lZwuqv0VTJp2nvukFH8zCrS4x17sbn3S73s78jezEPQuQ9u6s8dYo4x9WCkut10M9qJkFfF0rByD
Qw/a4mQ/wPjfbSdsC/cyh4fxTtOG10oG3SA9ZmP2N8LyNEXfhKLB+rpSlFSPhcNe6X8zRGBmYmB0
AIyCc4CzJzQrfOtgzwYWbWgdgkKfEM+CN1gTGbJe5TFiZosnCEWtqrwWYQokWrRGe7yAt8YLY8Qa
QqEeTqiK7P7L48YkOJVnsDY0ZJ5tKFqlm803yXvFtQ/06SCTmWIxVBLmkOIjNQ+jYFqCZavtSHD1
42baApFmFJs2osPBebZVjxLiLPWdcC6scVmNaSd82Ot++Fa3dxVwvsZ2A7NOzqR105DxBEN/AUd0
ecl3ZCslTkKQnPTzkit2SAbFXHg0bxnoKGWfbkhKn/GpLXC+220XO2Q8v94U3c2oEDxLViGGDJPY
Vv8zdUlcNvIUc6HPCZUJ5yW2LBZg/GaRr+MElUSET3eVVoz0plIiIVFZZ2axNj3tXUuxBfWU9KXc
k3b0Tu2ThdyDGYP8BF1WWhrxbEPL6MRx3QVvRi3vMp4aqHBKbUv8nzgUP/H5qb5llmNbQS0Pgrg3
4kxjqzz4M6uuEJYE9V31J+tdXLz4Wpvb/Tk2olTn3S/N+jV8OZjz8uUgWTozZs3hnuDkxQ069xQq
CB5yHjbNThliHhxCAA2aDV7Z21pOa7xnnxkUHTQXyexUBDJyuqDvdIDxj4oip5gcY5k+fLKgg8ku
o/vjPwr3+IBGuMByj/82jMIMSG9YGbRov7UFuCYIzgfgi92JM199GGJrmnIX8JTCushLBdpe0Vz9
nozrPLDbuPF9cF/zJG3ORzA49i9dJCi5vIkTdu5qO7OygNw5atM+2BVC9TrncUt3a8yrf26Y6k2U
zLc2XYU9S4dMaM+HRCmz3idEVLYYjVf4sCoT4Q7nd5yfr/PUR1m1wrPBizP3HAe4yKL3IYrSSenl
F7D9213WR+UZmpPwX4kd7fYTPAoOiEKrZtDuMhJzVbGASvEzinWYzryJ/LS5Endo0WDqRRWQwuvK
bFmuM5tIM899rIW51abcamX1vnrJLp8SGuvsBmSDop0Po8XmtcuYCFR7fuqWxt9MZiihRvOzRENO
sIrjU5Cd3hnvCFY7C+rUKy2MK6CETulxHZTlVyVY/APvtrBZpVjKDnCI4GD4axPymErtITx44a61
Riw7Rtp/5x/zBqdgNEiTX8liqBi7c53Ny1Dd6jfLU20Y5aFrc+C9CQCXzS/5xwuue0ZDGkMFlSJs
d5WoQhxUeDhXYHkDTJ1wcJuY1HfTOayBNmLu1A4VCuKKYYqygGjCAWK0uN0odjhnnSoHn3i1O3fB
uXQtmAaF/Fc7BADmSBdyk1gti+wJ4zKBz+Zg9cXYm0HiF2UuAFv3erAe6SpYyWdkAORV3IMoWWFn
0kE7K6IBftaObVJqvfDVDRkz6coQy1PWnGuZfK2wBbRSQhVSkdLtAUI80OcOwNckuQYnF0UoGTvL
HH8a02WD8BfAdPbFbRIMROqE7nIM0/MvXnh/9pNermGBiNC6AJoV1Grlp6913uTpRKpuEE4PnQSx
dKI4pJoKZhou2kNhDmQ7P+b6SkjFj4H2NR84wEXFmM8UFmQmJnKjOfhnL/p8FKl1ItWdsoqYl4W3
c49ytRDcxIJWakjnjZ2GfyWcnY/AUASfPd/2FLQ2xHngN4bIbz8O4UwmiO04ST/m+I7SvP+I2EPL
jA71cMkqom9V/XJCjFe6Wm+Y9dF+YlOsfuTZ7nBywVR+usd2YBSMHsyptjlDWugrvymeo8AeK2z7
mteri9/1HyXJBQsKFbkWmtrJWMUISFocua4PAgpsGcR6KNaYXPE5r7kT9BEY41Shf6jpT3CGCJgi
F65IbamODxx2hLT9kZxjQKmqD4uLiPnWLho40kkRVtje14mVwElLbzphfLVyMII9u1uibnIM7yu8
UHFRVkF7gODskp13Z4RbxxPEHS3FXiOjbzQn4D9AR4+ajUyZTt9Bxbh8S+IED3nkFenO7ZLJoUC7
FaL85HQ1R1JhVHDz63FMA1wsm/QZa8bo9NOZHR9FR9dHeAFaq3Hlvu+MaPXnfZ4bs3usxRF7d2OD
7ardk7FL7xdMc7CeJDfg0eIpGGh26hkPb23r79+j1YAu/fRHGa6hMi0GAGNmcnIl49pGpo3nmfxY
UniXDfckCqNEE1uO+Gifsr6j0GIaLoRcKDE7gv1YOiLdKjJklI1Hu2PHVw+yEoMxdftn57c7utCQ
qzVGvBQl9RaMYLRzbCCHf0xsUJ5Eic4neQkkIYa+/1tJcP3/4DGpvEOycAp4WQVHO6HF2vh8URMq
EclIREnaI+ekg9qFwk7lww5UiD+NCMSLaaS6GTKFJnQGor+DeyyLB3C1+V03DK6+Ja9DCtyfacGv
rMtdac6zMD+ZPu3M4+4Hz2rcZ3jL8xtNR0dwYxNGr4X3rXTJcu+pE9CzQCZwRHXINCKRtn8oWXRc
vIHAmw82EhAQO/8ujTJsZ1CoVm1OmkxQHarbOfFgaF5B0yk3eH0N0T0/OZcAmkmxog0BZI04IEKw
j5pagJK8D5tDYZoEIxRDITSkf4gOdAF38EqZftA1HThowwRYfnnH1eaNHsKCxP2RAG9YgLTfjidM
k3Fa1kBf9vOdIwA8ZT9znx9So4bcPvGIAE2oQ5wnIm+LjsS3cTcm/4xyJVIsWubw4UImT0I2dEYo
/zBvKPvq0/1AJdTRSw5LFI4Qn1Sea3hj81H91rtZYyPNA9mDgpziojtK7QBsiHB/cGrvPxyswYz3
wcOKjYI2c+5U44dpRxuEGnhgNqyPlR4As+dHJvXJCTdouZ9rtosNNkj6nBBG7wYeV69zIB3sbRy9
Hee5DQXiGheB2uG+Mp0xMZRoBDtr+xuziybq0BE1B3UyNnaN/pQtpNh/pGIEkkOVZGoU3A3J2Xy7
0XCEyXwqtioV/vqjU78u2TnfF1UuD4+RqNiWZ6hRiVgBOhZNaNycZ55Dkv8lJvRPTaMXwsIRPNeg
t6llYWfpVdrus/DlqtG5s57AuQhJ7PYZagsmtT+QppsXda978C6b27kic1zGSGBFgkQ8kAld3kUc
ptx26Hgd+X+Mpsbx6wn3q2QbClOfCXNSHWF84Ncyp2+5+WFcgZpSC/S1s3pHbRZLzvMUuFLT3gU0
znOOqiNp+6/ntdX3JW9wXwkBk884mDWK20oernXcJ6Nyu5XeZIxHI1s+KeRul7uP7vmwn81aftKa
jv6a9Ac2JD0tlEN2Za9UGHzqlcNy5HFgHOr9n76emWPvkXiGqEFxhcvNm2cRxPfXqnSYvEktBrLn
gvN+FY2NPu+vbPPTe7ObdN9Nm21N4Nmgok1ko8x0cRFkFoCbakiea3wxvA6KZGp5gzbPQ/qtFumx
uEf3mUQPgUaVbutpLEyHzyjY6nuJk2A2FBaRzRbewiC0e2Oi3nnkXzzh/S3N8c3oZQfc6VLCr2Xl
B8VmaATJFeuiAB/RnQb7DKRhqVx7qG0I9K5Up7AJcMr6hCB/DMTNcIGBJaKwhJjHhY3zHKO2IvKc
a4eNTAzZADILmB2QpQrDhdvFLPik7oxiEVD7u3m0a6NPJNmMesC7hTNzmjBWYxg99qJHxv7PRmcZ
Fw6Wf0QkQukrJR84eQwsoeGodO4qh4wRcOdIIBVl/WwsltglHmWJUE3t3DzZdH068NDX8QWBNnjl
8ftW4H7VKCUoNYwTpf0FwXgz8etFdmEBLi/aZ2gxipthaqCHGLZqxI45UZe9svYD/7a+CsN+JGEt
AYiieljuTP3AsQzhkaPDHJ9cCnI9Iv5jbz5fU4t7MtT1pG6WMYq85MZnuhgbRsRfDPbOgf4SKwKQ
XCRNdLLkqCKYLXi0bzpTdewsmeGRoPO8gA42goa6Rxzp1z/VEop5ywo15cuC8REahOrryfzM6rGT
38Cj8vh9izTYfApuJpsjMaUB8peNnl9rgqadJ10bSfAapIYUJzKevgSuE2cfzq1d1p/cCgSE1DVN
mQ0J1UrB+BNmOT09D5suJQPG9xhf+HNDMf5oFMjQaWlE0HqSvUX1CA4zvq/3FOYFdSefFXHIVL87
zp3EOzILd5QlLYwYiQeykjaOb00i0GnQa6H/8kQ6eSbAkGWTfrOOXP9Ru5s/6QJp3BMPI9jpVTRQ
nCVXS7v2T4ElBRG6SEnfvKI3W3IeX+MHmruZ4JQ+Wytxj5BJJ5U5SnRJQW9C30YphjmK2ik4mB0y
xEowEIy5SEqXh/FNvPPNTX+JzanwBSfQm9DZYoGMqDWfFUP3hYfg9nNwZqs84brsca26do9iKEzL
nZ7964Y5PHDZB1slrv/A/J+a871kFHzkSq81aux3MJiRj6j/iWJKtWodAACOvs1OMTMGeVjLo32o
XkM9Wh2GGMVvGJ4vQUztphIRey8cI7AvXQzcnDWxxiOSWCcNlulPAjb5SsyIq3z/FRp8m0WD7XTq
RYQHQoJK84Ztc5LKHPTjeWkbmStqOPDfKRNuFSNFBsJq+JdiU4j2AT9OHtHHRpy4joJZIemliLg9
vfWLCyCGT0BSYWLHpYA/X10Ac0byiQTXs9dFNPYld2L0a+beGKbAbFGCF3F535NxWLVkOK51D4XI
ImuOiqShjNEYHUAIiuG77ubPXDkBOGQeartb/9UmSw0u+6ySTWxR6M6GEXCYvUX/s9koXwGvOVrF
Dvou8ReSTVdjDDQig0bnwl51c9PdE1F2Yk7A/P5Y450CWZ9ch/Hf+U/xdNl1dyCCDpQqk59ty62b
2vuc8uJxH3PyHZYCZ04sYnfzWGsIwpjcyVBnD6GP41OF65hFuJuZdUJlpCxfBmdNipsxyf4QykKu
K7X28MgSYBwnSP9sqwdqhLx4epyWB75w8MjwykMsa8XE6AnQCI/TMqVvL1Ieq6qX1TbqOrkVa2W1
tW9Mh07B5qDA5p9QtjT6lso1gynhcRJc9+yk/30IfnroUCcvIjQDJVbn4hFFdpQFLjbAoq+geVE+
Tg2vGFRdA87Kx4XcJ2D2YoBpxVy34nwY+Eew/JrtH9GgSOjezz886Hzd3AskHWUTFG+10Yb48lCK
YAUj13gHIV+PBxSJ8so0UTbh82TFzgQ1oNlIKPDZ/xQsmZGK34vMvjEXibHBGGhpbHlje7n1Ei1V
q+D3KJeSv4uBfusqS6lPJ7txSec/kgCnDD87g7PyCl9SITznCBITscZKiwsrD7pCZEyW3UpFvDsX
ciLkHLRw6UIVgb52mwCrtieQpvQR2TFWIpdlX2jy2lUdx+jeMbXMwRj3fIuBMuBJt1JMGEajpH/f
hGFy1ZidAAL+CZ80X8uU3yklKtNApAQZZi4cCkRV9qAhkIXQwUwdPCm+B+Vxdoo0TKoREF41p0hb
InvdWRk7KOelER5AKYtShzn/qsqjDEUHdxn3VosNeq3qGRKQe2e39e+OaoC5j8P+vU1LGpcuJ7z9
OrcKFjjhHtPDbBbVPNCsmhaHbNhL5N2BNJwJF9gvfcU9akEeNP6/MuxDyjbcyob4BgNlwfzKwl4n
BC0iB8QBVl3TshLEGz5jAcJt0BvCUD+AYYmpj+cTiCE/+zsWa/NDFnnsVFSBpzS80vfpgrjrSA+h
Pttxqv28tnPZpEQRYkywau3vdu+H/s6AaH7MRM+ia99oo85BaaI78pa/x6tMDqMzq7s0DTuHIMuY
7hA3beAiYd0FCldqkXU9pNQsGvVSt2yK0/WGCBCIxSVNMwXlxv/jPmvL5pNq3MQ8wHWzjHmRzylK
+UdudiNJOC3TEhzQfaitxPg2WJHYCQ85O79AufkInAEAcdHFq4ss1NoNl7q+yd10uabZGc1DDH+6
z39j2I5qoV7vOFEdqzc3EfMqO9wN3cjNHNyKcM0Jdubs3hpgOuqYR/xo0zyROdLImEzReYZBvPui
gKZ4pt3Ut2yo8hE8Y1mn8+RE+DHeqvwuLyvwi7bclxYOwONi5x1XtgQ5LJVdusSL4d9zx7w1v2GK
p8KQYCH+xA+ys0IFYVKhDASgb1SrPGvK3mC3GPX/x+0spTgWyxJoxwhgYmJtfDHdNfkPqynUqmB3
c29dSVpkb9NUMNAmY5snhC5p24fSGSuraB2tiEW6ZrzpY2t9yIiv53gNhmDioR7WR8fJ2aera1LI
uNUFmUjUXsOfZ+pzxVMMsZGcI8l8KOCHcbRrlzhkz2KNf8nJIR0hlzTBeMDTpBj2Qw+XX1tK/PS7
XZk92T0iJJTou3G5wvLVk/iwSq4AXFFb5PRtK33PXswjOEWaCUFYTb9Aeaqm+FTH2/Zad+r69gvx
OscC/YZwGLVpbb09hTKLG8zI8mayyhzVJdHpWVaCBvWvMeAYMtpCLsIMFwHyh8JPr2TDbeBdHNPS
j7vWthkJJBpwJi4ot7O/5A1hmNV8JNVGXAKAvTsST3fpaFbwML4Y21mkAQ4qCq+137WrDyN5kuX0
BT/KXi2e7q5R4oNsIMBoGZkt2QzWNwZnEBbMiCEWJPJpjobrp8KpN7qTH2DVY2jsuOAe8K7qb4mj
SVNmSPBJSp6q7AOxdanHr9aDjkKxo0uy0HBR8Uq6nTGZnJuAKYSL1iVeodJUOABEG4HoGNsIfRVB
6bwat7cRU+DWtjk1M3tPYj3EeIspG+n0nIzqFpFJ2e34wnwClllxLLOx5EEFzPpguK3T5VO2Kz+e
lIGVCnIIz9RxZhcjEQlYG4EJwaUV82Eg2272In2nYbKTS0z0tynykiKxoYyyPJqgTI3dmhjR3ydI
EvhvZnJ5pfoMsgx/34vNQVb7F5mNXQpl3KVJnx8hJTRynRit484B0BGb0NegBFJcr6yPMip4jlTl
KcjsGsR82v+VYnLj1/G4myHuT/zuFlBgxrmHerjGm6s43eW+ok5Stkqe3WSMrSgPSvHPks9PB3K4
1yt/Cb02muRjqdNnOz4iPGdweON/pccjnvr/xTSya9tBHQVw1ySgPKQ/zxRqFZr9M/LEd8VB3PSn
o1F0m7v8TeReIVp4OffdJ0FgeczDME7Ui5lAnVI8eg83BPuLQ0Ve75mGrnBIWp9pPKgomIxqnwzs
sPrXdX8Tgc1kU7/6D0lS1WrW7RsUzkNVQ21zK1Ldu037eib5ZcidZ1hOPFCT+4G49S8EAkSZbQ/F
fFU6GyGPkzo6F084eLT9Yv8ub6qBgP2Q9uR+zP1hDLlumBrH5Of6Se1t2RU67bWRQuWQQFJt6rem
q/Z50HSHn4wfyIzXM61RIL2V9Hz1DtCBf8BoimlHzn7PfzkV2dDlTMEN5YmqkvPMsrMQzcybub5X
1tKR9YPEFjdZQ7wqly44XyFIy73zfr3o4Vfu6JqOHKGLBhWPcE3DQz9UGBxkDI7DZTBsqouGRzE9
RDyWOqstYoCzC5MmdnujrvdS0L9Mf02Ogi4vv59XvNbkN/pUxI/t+vnTmYmOZPxb88+AT+SGY0U7
nc0KjfMYZB4FrUwGl8e6vVLS64/3th9Ty9Jac+yVm5XtvPToMuH9Zsd/D/wDjxoDliZ/Egytk6ye
6TlYjf3RwYcI8WYfbYpi+ctIeYQXqu89z/VJD97cNJioznjAv/Kn3gOD8czbpx9GxF88LMUzzr7A
B1uoSWZCvNICt0jw2yMG/fw+0bhLeIdQkBeoHR56Bgm/7irkOs9n3KKUirI00AoWvZZyoTH5pVFn
EG6lk6pdyWceNUN8IGHlsQl03BECrdAX51admezg8LGPgvR3WEaOgc2PDL0HfkEL5St4Fkr+6KHN
J7Rwus23+BeNR9Q9LIIlo7auWjK8ZXdVAlsylQUbjeVkStFpCXNpTTQ+otWHy063QKYH/Hig1rIg
F7Io8S2B0blnsW8DpthUXJBMvuhREuC5648UpXgoiYqBHgaHRmwHfbmwE+KrEBULppAeE7KEe2mK
PSWcuueBlROawO/hFKL0IdDY2BDC8S0lgYgYfrPsawx8iVvo87KPolyaqPRANakdTFXPQQ9FOZut
s8QbSctLBmuRwXjUE1+haYm6T0faOGW3mr8g38GGOYus8+Hv+5AaYIX6Vc90gvBp1CX5hzSZZNVk
Kl3itZ7NN6bZ1LGY615cVj1tat3V/7LkTwsIpXsXcwXzqTYZd+Zu85CVmaZH101ihh1w6u/X7rKP
bsULJ898iGqwqobfiTOEsHdZFvG+r+f7XR6wG5XoM4Tj5H1U8FejvZ+f8YQvUDrI3B08CVLf+MNJ
rnfbMZ4kVpAGGJvqVz0S5DllZZKpJ3JV1eLB7Qg3hxyE+8VqrdiGhSGUSDX8le+l3BF2zL41Ej/F
DSmkMUSRMcmHUI3QE46coPny5+iEYxdTTimdEDt56+WEPQ8ODjtHcSnoTbzlXvaCRp20EPtZ8W2V
S7zkgBKk7AR5JczDwSYpHOFmc4PrwmNjlldQQUl45+vtDYOJBnV7eplIUwTbh7DMRPayJTbtASaV
wZ8vQoYt/dDAJHBOuSJrE2peMfWD8SjHoiLHg5WLShtLl7xz2fIqMx9BvIkdAiKpA2Xshm15A4EX
Daiq6S/VuAJG90D+pCQHvnTlbgtAw9mOZEKqwDueknfBJV+EXtohYgY25Viq5WXa5BCHCHZ11fST
PA+4aBbZjqPJCNpzEq5+5ibKeqi/DwtFmy6s5nl6FWfyb3Onb4No08lax7EkLHc7OkUwda5JAA5A
jzdr/cFYx/p+A/uCg5diGvSfGlH+M3DqHqS5uQz978WbzWTT8sHHS9q0jqJNFzd/DyqUOKU/IOW6
n/Ko/smBHEWM8FTuXvqLwNkftDAXc7tHmG6sPnQXYpcvnw0VbmtI2cERCeeVXwDi5bXCJXpTn4da
MjyfZeDPCKlDS3BiL9nQzygsDIco9h8GOzKOFUlxhcBB5f1jx+ZvWZWu5IDIu4C5ruR+6dR4Gr4Q
+wI85J32Iyyu7w3oYLmdQwOjhhUkf9fSCTvRNoWtAWXHockT9oZ81+DtpTXey8tYs7UVCnpIc0zq
8zWiiOIobsBWGyS3z3AjN2WUmUDSvF72UK2NW/v1ldQyLHgGHjNkuAXPfrcp/DTvy5Qqx9Dtc9ux
HFvMLwvbmd+QgYottAEYgEacJ9eGH5Cdpcd/4Q+B5JwisUpBQY5hcTjB48E1SlfusQEaQKesqWxT
rk4IUe6iVnNUCanXpNy93CNkZTN2O3oc9DDDVVnCFTfmpP3l6LTL/W7v/hQar3A6P9uKs3DnLvY0
AS9rm/u6BGxTasB2Y7169/wRQMa4OsmZUbiY7bbOd2EWiffCcwlTC+dwFb6icezXBbjE50vuIE97
EedUo+C6w4L3TFAnl+FLX9f7ERTMSUOC1HTpUqZlWVAJC/xfHtjmEVzksoisDBn69LLw/yc8d+w+
D2ln5vnyqc7ZsUat05IP19QFHPb30iUV14D1TbIXsAHAwqWne3dW5cx7W6qqAkAM/AoC16ayWuiE
Z9ERRgnI5wCuIQbYcA6qm7kGnj9b6fGRhAQ0qkrxZ/TbTAuly2Bdo3G8UoIgETBZV/CB8HlXVPJ/
jryDV5XT/rtMrr9pJYWi2b0PFMm/ySHsXYtV7xzssc6vwIvrE1UuX+ZkSdrxrdYwMIbCqOs62FrD
7qvVzAWh5Fz4TcC4j4vtcoE+bZJbxa4u/NG4mo9Btu53NcEq104iizfMR2P6EO4tXIjUaiQidaQB
kSttFwaVrak/tsvwgVMMU8hgF9tQmj/heaiq57zpEzhZn/yMW8q8fBK5d4pah0azf6XiLnz4c7t2
hzALdatZCXaS4qn7gt49AJBnsA/J40WxqmfF6OXUby32tXeG4teSqznJ9F/atvcegnp4u7kajiNq
J3Fxqa2gWCqmquTdp2JbFUVQrY6BWqKKoXeFK8AklmpvxE44+wNEbic2P2y0v+Kia2CybzUygvDk
I9fsrVB628NyZjkI8PSjGQkCDwwUuymqNKu6TEkUCivROjJ6F4LjiV0NhWZgtal1pPbpN37uOzW8
Q4WcgY56Gg96Nx2SmnTPaLXPmk5skQG02OV+Y6DkYN3Q/XI1UmTCWyLknc9Z0K/Av2YhpgRdCzih
VBi2AzvJ5ylPt2bDi/ki8hoHDGE7b9I/WKAJ3nqDGXaZpqSw5CGpUQ64yPYxappiqczeMZbmtjib
PKa2WJBVdyP74+jX4kKsj2Y8Wlgv/AOZmKpUxf3i/wuDii9uEGxFw40KCCNghNRfl9X0uCEyoVXS
Gg0BBFD41J5gG+T5tzRBPLBYJXQb8rPriRfhNj+jR2hkkerA3iXljXRf+Z+9KoLW//hBTGpxoAPa
7Rkd2Q2/Cc/BnfOQ7dz2eFwyrRBe2+xe17lwUEYCWApkTndJAlK0oaxUQ2SJYp4MUdL3/aWUVzYS
KSp7oyhCuRXYnSy/jFfsIMDXXBn2nYGal5A0UhYN9CHnG7kjuJQcLxEEyOzL8YjOytvP/+yoz0fi
hSGvyOuKCaB/Bl/ULD+TzQyCtlf7w5yycUKPhcz9X9MOqh2gy+s++pA+bFVYmyglNSjd1JYDoV/u
wNpzbkhbSZPpPHeuX3l2rgS0spC842mc0yn13VOHyIth9mvr3RAms6WnlzMEF0iD9kw09GwxkEpE
5w7pzeg6hkuIGmQ59KaSs+kqly/WwLOoRx6ISI2dcsNLJ1VBpIevJNeuvKAyvCWWoDvcw57hZd1I
o/xqKldv+KUUO/NURrjmPwnTS5kQWCKzacI0Ht+FCnLogJb0eY3r2T/MTSYw1PQDrqV2S7TakD5O
B0KZemH07iWtQ0rtzyHNS6ZXRskIKJDC9Ev8g8TTNjBo4jES2pzMG1VxUT99xDGjxKsB+vKlohVP
9ACcFJN9eFVv4kq/xhRrtupOOnrhPzu2gVoGFYeSzJjPPu/sSf4fcMO9+01NzH7oyO01vCjU93jV
NluTiDTlM3dCQiC8aug3dddgNjyU2kcTp5cAOSNNq5EceHjWFZ/ExVOf9zsmF8Dg5Z/Zd8GZ3Qro
UxYh8eBZik+cW5IBCFEBMHtkRyzsaQaxR4Hnac/oJxrO2DMnK9kb7r3pHWgYhlZaPyXCk5V6bs4k
E0fPFxkwH9OliBoJUP/kjuxruJvdnxn3rZR7qCA4RrBFlSZNmgjfvS+7b2xgxpJc2V5t64LP2cyC
1S3yFpolwBP4ZjtYAHgsIQSnDTjEjvwYr2xNvyWhFhGLBYJ9LIQRrZY5qokVWjOkxEDF2q05ZPK9
SkIh9a1Rfn59FUvqHKUiWTLFiz4wXgwPEArd5tCSg08IAoU+o2A7QInLPlOHlvdGrN08x2LbdbIz
+KbZFLauVEViBgRs1NxLOQTKNWgXDmzNa/XKXxGbXO9Im7zkXQXto66MDV0kYrb7hr/ASHKL7kdI
6wNHfTx2qiFhSl4lefMtEW8TGSR+Uj6+B4OR609JRJk2mIliMpisaNYxumNuGSMSlOsqnjxAEctA
M959lB73VmfGJsImrwkqWRQvmOdFmSd1V68aJBIgK5VjgoVy8BK+p9VC7IGTPrtzsAmM6TAC/9tG
JmZo4nIHcgH7juZ9Segijy9INVyOlicfX3uLjt3wftQ2O0Ogtoo2HdhvCKx0B/V6QTbq/oYEgoXX
3mgwKEEVuOiwNkFM9rczaR6tvMbWsSP6jW43Ik/Hmd50sFkX4AFlltCYx/NBdDSJtXoGJv4aoMCg
0O6VWaAmMGPSKbANxdXSLXaZ2lkDbYhXMmZry4X1Al1Dcrdr3yR/0TygRGOE6hg8pECzHvRWIrwj
opr3CWnA3kAguZZxdaIqbWfjG50ltBpt2b6IT+wMZopWziOn9NYMLH0+LYF/w7n+qLPCYCz2xFKh
6KPuijzyQIAwfFJklKBiLMHGffIvCzkI2hd5lk0QEVZOQx3SFp7ceba/qEUf6sI9hTan8Ib2iySg
cVxH0Ios/9bUnrt2akUUQr5rICUHtyAODdMWjDqddJWkZzdHvlM9rFRW+7dDOgxxhboBK5+SCc3t
bZipDgfDXY22KluRI03hTU8a7iQub1/7rRSFWStkcVwzdUMNMisIPRWDPd8AV4BOhq8hKtfBhlYv
LTNbJ+Wvs1tLilPD5Q3/ipXHKcerFrLcZm1/KJz0Z9GQBvba8bZv0VrrvObJ9KImWeodRj+MlDNe
zPZGDjD2292h1mx9saRzabYG8zvpkmtcclcpQtmEa+GpUHSwUdOchMfVfOZp5aZiJSpRIGTjptPq
EvRnmqfntG29D9JX1PQgavzWJIHFvBFYH2L/OIjs5cTGGl4TqoOjGXW6+98HjYr5OCqC7OScfR07
pnO5EYQlieJX8+SEyUi8U3r5BXEyMnnHTcmSxYKMjHUsWPOKP0tp4T6y7BujjQJb8AOeN+yHCMhd
HA9wnSRzwy5sDgrRyi1spAZUzizX6zmpoNLDKTpfEsR33FFgear0l4fq/yHE8Y72E6CyEzzvJKxo
CLSxZ6AcguLMCp41HeqBEHOLbsC1ROnj6OvP02XJVi5dARJ4QbO2aqC5lvHr4hAlV2UDw3XcpOIW
/pWBp0/nlv29KwOk5gffTXicjHYVibJNU8rtzWrAcp+zsGi14t99f7RWWex1wemcDPhiFEJvyHzY
7Pq0eeD0krxiOyjh5mdpNinBJMZLBxbLEk6mVD5bkJI7RHW6/XK0h4SmcOX4f3+kb3tzVxzh6s3a
u5R95F+v89Sd9/yIlzbEYz8rIqFLwO7qh4vJt5YK0szplx+YWTQ4cn3aNqXKGR8C7maJI/9fVyq+
Sqv4/Z//SRMival+5FTy4nY1It+EJI+5sEGipowUe1M+LVxcr3Ti8luOIjxhuSUPdKmcJTTxzcdf
+5PYqoQ34467TeFuudX2zqV5SxRUvyURXJ1UTip16IciI3m58CaEklyU7JbD2+6wnCi5mAMDkP3a
W/zRalmiUe8QS3h2bMjWJvLD/LJ3NArHS+ZzpS9fUsbCMovrgxVDWZ33En/5xmKfi2O4bw3+Sx2h
Ua53QsuZQZaUEiUndBVuf+XLO2eHS0yggH/K1nxnsn/SSWT8cPUXuQ/tpL9QUg8yHlL9d0Kx3TVC
Wi6DGO1CKGLpD3GRQpgk/BigY8s8xPg6zTwPIuJBh3KD5nc5dBVvuHIvp0rv6OHgvoA0yDXPZ7Ta
RnSO+oZ+EjMzh/LeBFVsdJPmaK/jZa/ldDwGf3aDM0SvXyRIjARqx4mnc3BKVloXwvwFU/QhLflF
hL/UUdf1jX6dQub9OcypZt7N0qTJWNLn8u5pyF0xgrhKPkxsZJuFlg8uMh0bp6ej5+3iTxCcyDG6
rFSlD0E3g7bL7dyrBIn/9AEVr1IyLkcKdoukGexEr8YJ0HH5XfdAB/sXgt6V6FWLEz1onmxE3NoE
v5kEPd1LGaqjZf5cIJvqPU30OG1wXlIhEekZapFWBsmC3qZOG+D7WcD1nNm42dsKBcWb9umRE0DJ
a8LLntlZa9X0lpKyEcoofkwZdx+uNScbZdKLtDMXLTWjfuh+EPCyzTWUgqfkWhS97PRi4p1THDPO
2cHyX/AWnO6KJvaHI1opUvazYGgbYTWnkoXy9ABhZjPh3usKf19Q8g3yhl0qpan6Em66IqIz/pAK
VQkts9YH8SfZX0tfgh98zGWe5zu9p6NNrmMGxa+rPbJUJjyIEMbjUHz46WUQwmOqHMwXuBYkhyLy
+yXYizCqTz/FFbVH9UXAOnq5j1ioIp2TboFZ5t2LLPvHjWProG6h9xyhy6ZSX1yGIIFRSWgsjg86
zkXgvJvXz8iDngk7vNil+KwqJKGMLkvSUDPkxuhH2TyeQwGPAR4ci10EZQ70POpAbC5DnOL5PN7W
73e4Nvp3nGwG5OKATWL8ow2VngAYUoucWp0N7wRi4fAdGfLcg+4oa5j4OluCBhNiuIbMjojABCS9
GOYpo3lPwfallplHpXziXM57rVYRt+/7lSq49y3EQP2muHH0ub8it98X8I56v4CGCuOtSZZIOIEZ
sVIRosFUP2PyrHlG7Tb6+KJeFCRHhamzgbmO1lYxYHpCQAZWjB9r9x5tYSD8dh6XYnKMzgF1obMN
+WAUKM6zLni1DVXkiXVSGxGWKONrRu8Ws/DneRwpMNQvEt4bsb8YQ++Br9eQ4GTRIO73myNx2v/p
pHMoydT0LXSOCB97BBaCudatM+ZLH39E3Xhw2u3FTq6b3GoQ5SKfX6W0H0mgGw9NTL8GZan7Dk9C
ecz3QfUjQAMO/y7yvMLy40hxq+keD9168Wr/MV/EHkq6O98hqimSCGwvdKToYcgWGnvsequygm2s
KplA9p4lU7UsqjEgmcW3h763WB0Ppt7ps0AIBrN+EWukULxBULw/n2O6oPGbzy57uV+AKw6GywmB
xrXQUfKSdClQpV9R3tTL4+0oARzLgzPNWDjWG1AybbNjHRRBD+g+ZksorF1FpP14if+TsoLLZYRP
uGoG/w1pRE5nuxL/tkYew15bgsmmFpeBzoTiN13ccfl3q+F3Iocu4jsFQYD9pBggWK4A6myph0Qb
wx4vcJM+HL5uyUaKkkzI36xFS+SmVv9U6jM6kPyynvr30jSSfwrZYmckXLuZsTEAo2A/cQERo6yh
zHhStk2MGqNr7jx8Cgq9GUbw99WbDzbiPOxjxwFaIeB49GKAN5NEQqp/RF/oIoUR1iZgZCEdWgYI
0eddiDGyvBvgZekpYY5Qy/EUANxYus2Q5BlMPoNEvX2GwzySBXf7/miziK67+DwESRyOAhUI8DHR
AKRfbc7SiUubTlQ70lQw33pjtKqz7mjS0qGpPv5l+b6/+1NbbG+uARQ2tKDaWqI6w6Y+1gihFvDU
enq+limsWt3dy18wfeMX7w9C4JCHGrCyfRi8u8ybncCXoCeQ7SpeDiPXSrciycfj+fefiTb1Iusk
7V8ILB6RfjO8xdwgBNSpuwgFt7KbBvzj4nF+2Puk7HUVvmAwX5UVCKb8v/Gq5VLJ6HZWrs19pLIZ
F0BlXQdj9f/uNS6MoQsM5OeAbtz3ga0v8u/amPcMiVyzjLZCZ+1Cly+ySoWPMz+vcQlxhyify+aI
DHG/w//bI9D2YL5dom14RB0u/SH2zjHoktxs5YfAJAUlv3tVWk8LD27pwTppJE4OFl2HiaYP3OKq
8MtCGpQf3U4DaX14tA+r4TW+grz+W96hzdyhWlUSz3bzMFwVVi9xlAsK9iBdhhM0qlIaJlRaRDjg
GZDkJTzzX0jqXdxQa8RqRMuwPfyXagXGb0dY+kj/AITaVaNDM8muSsoZO1pc/RFwOX4A8aJznmvK
s0fzI9pU0r3UNF77BaI55Z/y3NKemMnsjrgSo0N5lFKAoqkhiSJW43Lsu/yRZhpDojtYLR54zgQY
9s29yooisOXQSQUGWx/GobZcxyZL12RTpKPTr+/Wa1GpLiUKexGSJFpkA7EXrdQHZnE0QGxvJmw2
dnbOtTsNnHEMDih87cM8ZkUpIvBkczhIAFGNIsT+0Q/h0hMZ2lEYZrCiil3o156L9KNrrCj/BIao
VWMyDG3M1tSzCdrFJqM+jsnfgcst73VyDolv7MN34jIQCiKj3NHb5UUhga0MWbsg3YH1ZxvekTqZ
MeZjgu1fJVOabag3KVN7hQokMsLxxkOu8LUc2WHHExzs6xtvWKnyfM3c71roFpEZJ+OkP/T68ese
3xXYQLUE1FcxmjYaXijMa4/LEN4NTeX5fX38gMF7kne7VXIAsIAP5Zl7IuG1+3ySRcQnQV9xAuxU
DxN8BesiJX6IppgWrB7hsshH45KKFZttooxH2ovxVOPgJzE9salSrc6aR90AQbzI4RX/YMjs/sa6
H4ypmlsuvisuiS4/WEnp/hfOVzA9aPN/BOpNjOu4RFvq2uoUARxpM74A35Uw+VBylivSDI2QfljJ
Qc5xccDWRScE8aahPXE54on3ITNiKIqKVRW41OpIkGLrLyIzAeJ0fNWOfvlh2V2IO/hNlJ37qXDd
KVw/2oORwdRZodJhrge7wFZ90sKjwGIud9dX+E1XQAo3LsMbDTSaT2QidfN3RLwl8tEf/PHe3tyt
U2SoOJBEZ4tjn2hb+BeRAPR6yr7rrWiZiRpf15wy/PTXanqtVJyec55fkG29iE5oDyawwXE0sPI4
7nZReuarRJfS8HI+LBNRYd6h6mDdFhfCrMEqv+1AbsvI7OAX8BKg1UKGhiX3/DBQpd0h9h71p1lj
QjytGffkzQMhNu30jb6+upoRQSHy9tjuaQsaelKqCLoMLw4PVm6DnjQ+ZzmfOsk6z9H8CD6t2Uph
4PCH6CK/7yNDkOtlIuoGKc2Wzp8UgqS+2aj0kMkS/ACkTjNr51bIu8dF/qBpSsGV9bMEy/09YOao
ymV9UG3alh/SSv6jC3vvUCyIy9xILJxsOpke8RMAWa/wiLtvI1ZKSyQq1k1mcqxVtDmuGr1Ut/Zw
NMqmbZwCSvk1FCjrIdS1lK1lrRPTvV8fHKn5oEOhbFVCSfgs3E9KnweKgbkDKY9lORpKi74kDDLI
q5zxHMfnzucmXE6o75GWiG9wry7d3qpa2hGzOFCNUxzbPJUzKLmbFGEb4uz86tpaBAjf0bZssdrj
LW7xBaM4hbGit4nHgL/tjKm+90i+dD53fc0fXsnBVv5r9BDi7tc6r6QZaNxP9Ip4bETefEEYkbLS
tGAOIaoHUgFbnjx+CETnkFjWnUc07+o6qV+v3HVqimcye4YBklpesG+jv4NRBffYaBJ4TjPmrlsM
PlulJbh4KdRPwmk+agiJGwuhw9YKrJ/uipGgRMr9ArxgBzFGiy+WVOb4V49Z7Cn61ucAmQHko274
smNYr/sveUjaF65V2QCywy2KnTZ7utfpfSVxCzYWgkLIJaYo3TTiWPLJus8Pb602Nmim4WvEfYv0
zn2FKp82RKJztwNNWoRk/mRmwNuJfFGaMrpuEpTG1+If+i42RzWa6v6NVdzUb54dWmacU/Yjwfh8
+SW94457z5h23w6VKCdnkDtT80YmTA4EQ55aWZY4L/3j3fzi5S311+nBWjQIuP94u90AhtCTDuVZ
k+Qt1sY1AbBu8ULwDeVouWoWRwfTDj/OpnUHBZv08wXR18FcutI4F5s8fL4ZBMpaBVJE+zIMMGxI
95+lWN0e7U4fwcCH5hec4/VUjpQVa0qJanYJ91xej3DmLgOCrFLFub6qotWOCr90wWibDJkz8KEg
IPzUjfsDBc2Hm6sizq9DjwVoeNHgn6JQDJPybfetZraEQVl3oSiHcyoIIML4z3tE47iEP17jeE14
tDw6eGKx7+NSAGC0+ZHD1voRb5iVtwSXe6UQY7M4P9f2SnX6DSz46xVvh2Xw1S4mcfjwA74pYUWy
E9ihWnRINCM32SaGydipmDGnfPEH5mDA1PkYfPqsna9KBV9b5GGwUwLIbrHe+ELqKxmuqwliA+dx
dsa7nGKXP3aniXcR5cLNCu/vhHlS8gg9fzq/IopwD+54ZwhoXvuHlKbzyW9m9TCP3QBA9eQeSDCg
Wut63eihiM+WbuLl1tGWd6tUJ50WFxk01M4dP+weamOc//TNx2Fbg+OAWw/XdEcxP7ad2w8waXXl
19DK6TDCWrpU4ANA5LzCx8pJPctd5I0UehK6J1B9Bp5QiGvSfBKCPpM/B9Sllsi5Fae0JVAVcxGj
BZNZYiMjUEwUYJzh+ONoUAgXVe126Iup/JdzmqROVKoVvmyQIsqlFZEMeOeCYKZI4O2dWLZKg1Pa
UKUDUlJMZcJ4OTlp2KIWNFQgZrp1nBfzm+/QcmQOH41H9S39jcNW7MzDkAWQ4KcrG0nk+2oFYpb5
1/hyj9xASyiFDXhxo7Ood8HVWTrL+tdhYaa7+9v16aDoylZCSQAb6RZ/aLpu/6l+MAL0bCc19/2r
9zg4Wud+igqdSYlglR/iqiDeOXbhKfj+RRDKJwzZBBbrSLQHvgx37b61/Lp0UV8ZQSUm3DmaR31P
aGJaOLkpcb1o3dMR3BNqbkbRGVk83/GOWPABbWsReK5xYCdANrid0W3OvoFjg40i9+8Pk6nhW14l
lWBhTprqRKdZgdbmvVZ1vRqJxZ9qOrscqu/VLFX4EHZEDY0SaKxwToa3zILF2j0aGa1wqxSee26A
Rno5p5D4ExwjIi4t1v9TJpqTJgsl2ioGK2akN1+D52IIPB3yP0k8ce70CGw9w2qUu8aFlhNuwOz/
3Qzgd3S9Qhk3VPZCpuA2HLYNktrqdu1DHdslh5P3nhD9CYJoCereAm0OIrETARvt7aXdFvFAsWZc
6UpPr7pYk8yyCYhnUwsBs4cGBg8TATOEufjFWNNK+apGLUxQPhzOYRy1Z0xfKICmzas3tc+571Bg
E7ij5EE6nOPvUxMKzO6J+i3UTgqDby477NU9/sneW37XZKoduJ+0+iMaTNCDyZeQUOFyPosEUZ44
AqbcF1eJo9vI4/OyzXrSCzBDfwL1Qw4ZwhKuqheLADRUWlZUR4LZ5kxo3tZ47IL5Enia6UZSnbnT
xoe6ODkL7F8Vlb0AWnAyT7fu6bboo2E1qI/GGZDNaAlnnfuYtHyYhao8ZJJ1EEmtVsJNOUYcnGZ4
xNM0v0cy6hhfF+5klaqb+8k4w61LiKqXfU6fyZFp2XIm8lXiQMYd8/bDkCQpChttaQhGMdy1Dl5V
0wtpBijNhhr01HOABMx9aBgh901RWYEfz8CYLU1VFCJ+Hqy0iRq+lzF8JBReMIprWwZnzjr+3ZaW
UGdaC29OVpvfDecJDyoH80wOJR527FYv78zxvBBhrWrU7pvwBphHoEZXXmNn1czzQY3AIoqTKKz+
hC8B9x5c/t5Hx6boDEiM53U0afgqwpXmIrGHSg8Vr5hptMwrHrY1GV+wlEjvAG5AwX1MEhPDc9TH
6whwe2GtMUgSnu8iUnYE8FvUlG4Z7cG9DaJVaBrjDNel3htISbVyXvAqwZNuCL2MnYxZH92/oOZg
+c0XFGWb6N2SEnE2Noqqu488g15Z+fSsPYZAQSar76o44tTl+zo2KLfNdolmWJ7SpB76LfBOitG6
1ameseS11DTCObK33wuYZjenaszl56vaYGgI2Z0/h9YGyLoR9ui/JJEPF3beaHRAQv4NV1oRdnxS
h9WvWxrnFHfZVYgEvwIX2eqWvKPvMVNHuMG3kWgDiBb/o7FDp9N3yJ4eaKtW0XWvN13WvzKBsvmL
92hcHoVwKVo3Z2EPJYIFHONZ6XyZbSP5C5TJ7BpfxKr7LTgjf/GsNo0r/564bzeuW8Z/bHaGdjEr
cfL3dOcvN2tMgOLpqX0a7Ey0ThuALAZtAEqRdO+GDzwLjBdYpdtJp8o9qpEYxtzwnANh62yElsAx
jwoOaANpVrXsTBU41oRLLTXxkG8+mlC2tA0T0OTqL1N3Y7y5wX3rnVCJaSSNv/bEQN6W2lXf+j0f
xjVy5zBM4GssbXon7FzUUqJHn8EJDhq5Qca3fdtSBJ6lWi1OGofv2YLdOZrPlTci4FY/ZZTrdF2V
+BBxgNDgW7WMDmu3ipt1MXKOlZI7633W1I3qX4MKdJPCmWngqJuJOSxTo2mw53/x4GbUCWd/8+aH
Gozz8maYXFg/V4lTZN50Y5TN9V1o+THrhHz/EosBb0p69qscaVpCcOua33J9zM1RbNP5VIvae26i
9DSVI1yRsAKcAZMhNQDiCoc5M1/8Lw5N+GMgebljOtqGwMq1LoVlbrKl2ozY+3enMVl0/7IcQh+G
KfpZuS9llBjm1Hf4w1p20W/mi1viQ/qOI0jqAwsq0huHI0Sug3gCVfC7I3L5jrI29Y0B5sweLMhR
Qsi2ceZ8kyVHVqMCaNEkts1HIG+1AKiuRJLSNUpngFArs2uHTF7pxLWqh8sqzFCAabFquBGJZomZ
OlLw4Z+985wPFc260vsaHJJDXvxw+MHTho+FCdc7g9GesbyP5dtJrMONv7PjrvSFYZdobz1YZ0k/
NP413Ul4IQgbJuh6HdGLFurZzmt8mp5qLnVaRIBI4qVNYPeGRvakbSd3vbnI2heiCN5qLqGB4eO0
Q+PlQPicfcCjgJWoo1BFuEyr3T3lTO4KUU7hqQQdq+1bR79mOgqWn4gXjTG5AM6NDchj+C0G4ACV
RlDipNxQoat6SrmVI2OWCtTBBKByNZKgnifxAXoBcqNHqr1NsYOFuZ6bxV4LAXKKMyLIKPSQFPMe
jlRWWINbf/elyNDRoQ/ABFl5vRJKolcKg6ZE+6DdYRMa8iO+6DScgMqk+9z6YoKjro60PrjuCId7
9z2NIfclh8/Mv+BGgSkYwBeg5GM3Q29Hu6KPa83Gs2Gp13UVIVoHj4UUw8CALlhBFZeK/979RMTI
R2c7R4wx9kuGCnIRb2/TiXikPBQzZc5woIjkgK3t3Cx+AencTIDmjrvUPuB7sp0h3UTKR4JOvlMJ
gdBNpW+ZIDUNdSl6OeE8+NCFtcqB8d16qtCMToDohWr6FBlZkvISH1Op96pcU0yWtIFZeRN8doDw
Vo1p2ElMgZNq/ajCWyx5MNr/rGnNdBd9JiIVRAS6hPGPByGey7XLN7pJ4uFYOJ1+UDX48536MFYf
jGcQTjVG8LE+TY5GVdAbFam+1rYFTolRbMdEz05bR4Qd9+u3C1eTqQSX2H7JnYPBCfvOXrR/SnMq
nZ7QGUotwkQpoeY+cPU2eK/xFukI8Pl9FoGNW+EWk8m/Sg16DE0KS6wI/DI4SfWZEmDwfXD1JrWk
ISVubOednH14j9WUyZVxMyXLolIOkNytFWD9QwZTSFZ6PkwM1AnKJiL/5ykCavgQkhwDqPdrkYsT
zCh0Xy3EgqdTxfajtgQQJMwNH5RfIX6A867BzcURndsZ3wIWZontbktTMxJokcXpDsPrb+li0a2Y
ZZ/7oj+GhRr1Ug9QTxzrEX85doxypyKZU3I+SYCgevfOyPHnbcROl/tjF9IVEPwRAen5koIhZ8ek
IxYQQuKPJ+mc2FZHDPU2INTnsEEI0y2UKQvAQ/yXqWvNJxpGe04ZliXM2TmOWtcvc+HYAp3EYA8p
jZ/Qtbqx7Q6/S9l/zlgxnA2zgDU2cAeIOrahRqYe4bqHo0Ds7Sg41E8TbmlX+tHHJ0KKUbM++TiA
UXgnO/eaw+Sd7p+fUpsq6toyyWgY+5DYu79KMPqhfJti1quKgOFXQDZmAwYmqd1aaDyr5zYOFK9B
9YS/Fq2YEaa3OYB7/dIVW0DlG7+YuPKhCen5RlN2azWxTvBEUCVXK9OJWuPL2bK/LEtBSAVDg+et
BDauW/GnkAMsMIxY25oKLBTdDVMw6ZDOrKP1sSW6fGdduOiRyk8sAvnsqg1q9GT9uTRC6GMFKT3b
4KWdwxFna90oCW5VexIvCIvGW2yEkgs3xs/bIr8vTVYi8XykYOzCTo/IjHZYdzItEAV1gae7/Nli
jdQvT4GPQZU1vKD/htE/Ae13nAZ6e8TdfdIS+G0BH2lKwAjgnGajWQmOeZ/cXhzkDKwZUBCiKm44
uR8e+A8/G7EzfcDSFrtjxSLbXTLTtzzoJMzJSUis/AGWhDuFUu3rCaL2Uh3WeWBZ6CVjwgRSd32j
a3A8D8a6DWZgmNxQJJu6P4yAJii5wr551G1lE/cA9kHT2e11zTfT/pkkACZCfzGTMIi4U8qsyc0s
tOGOFKH/0YgJqBdDuH9IUJGZk04YTWBNGqXK/RhCFIdY5D+ZW5+3S/4PYagPOsK1gWESg8gr44eX
3X8kJiPH+v4L0AwgYu2Oc7zcWjOirBX0QzOQg0uYHzWdFTy0rhMWc4ezfajkCtaMYPX8PdlwDULv
m3j8HJmJTxvY9gauXU1KlkqlGmAGFZLuKYHuHePLL8phoNiFAcISGEImikXVa//9seHAWftjdLM9
6VwoEoQflFCENBH1D0HbagYxGsOpx5JYUtNkA1c44h/iUIr+hSJXPXyNmkD1jFDVaPThC97OAZmh
nYcU2/sDDidaEpuOGAH9tu1Ho/7TJnphtUje5tPELkWiFPH2tzIqs1cE3ScIaiqOm8DO/oxMPx61
N0S6/K2R1IGf0dkmZ6iYqB1tOi41d7iLj2jCqam2jsQodAYpE5sUQJ63Ic4qrXwO5pfAyXvE4qqp
+SmMh9CiS1fwS32ryxOFTP82F8zNwyr83dPk8PZfyB5aZdjdigZiy+SaUT3KwjReo8zIXlJOwfqq
mr9BWd+KAcpYZ4Kd3g+3hRxCNaw4G7OpH8KnebugBVv3R7A3fGZBiEub1qUzEG9YEPFSPJ4znN8H
lNc7WxxqislEF2SG1mwUf/roKITcuQ4txAPLb40qyN4FBRxhuNLYLE96WmgfizihFqp2hw61cGKP
Cbk7JlTRsDJxA2SGrVMvih8shLQjbEOsmbIkxPTlvF44d1FsLk0No+qvVZLbaRRcxFc5YF9KLOQZ
SFQyb2fRLE1kOrh66V7U1jDXOtXpI0VtMFWfzoNd4rUOORoOe2wL/MfZNhkbpbGNXlMcmvogyYHI
b3KKspjSzswkrz30qVHxb3Q8Z84CGhm24AiMqK0WQarODKJMcyolJrTRSIebuaw5YDiMNmmcj78a
EuF/18VZ+uJMeVNO9oK4sChfJe04FRCVUJM3++O+9MJccyoZqQeIENfzN3ocss8IyrkdjjMr0oJ1
p5TE5v2kc9Nckpear3b2rCo0Tik5nF0maM4CEf1guyZrSwdKfVTafnb2C5G8+VnFQYSPASDrfDcQ
RtILhthjx5qWOcVtzde0sWTTNlmIdw1x7E4YJEL019szSKo7pcT6uQXlszsa924gAbRQP4ND1ydy
oc064PzQXrZrwVYZuWMVv6rIwuqmUJtWtu2RFwCFvpSJ7YPVNmQ3MReeRkAOPGIBR4KUAYxDXZ9K
k5NTL5/ho0+yYsEyaOx5fTMjq9XszxeBP6lBxjEj2XRTEJhxAwr8pqbuyBJQJzzrScyfRqk3xKt2
lxuIIpeaT6byBIutiYtsGZgG7ACYvFCwAXlGXsfdy2ORbosNSq4N9DoU8Om/dK+vjVmrLg0T4Yd3
6acS8pRjxI7C8SAFgcQ0dXv7blRFpPsSIZ8SxxPqXnrwiid9DlK12NOj/dn4b0N6UhK59B5usGIp
tj+2+Qx6lGy5Hc12RaC+3b6U7Xmn5PaLLaVLem2NUvOTe2m4V6PZeBwpJl45TT4AorhcltbuZ4Q+
Fb6Y5tYteu62bAFuxq+XlbG5PHzmiiMOqoRFtwOEynn/lNRLvOxpK2wcEJbfi3gIsNRronM7NPzm
TwKbzmlxhQ9tY5U/xi9BkXxgrU8VJ/QbFgM4LeEW0fuIiSt+WDIR1CxkCQXnWUEfpFSJjGUhnZUD
TksVZcyOWr8XYj4GrWwQucQg0HGxMJBJ1cdZuF8Wht0sB6+q/da1druT71kqjp6uY3rv8CyghOMU
iE1Ra3aCeUseY8ecIRwFaZfCW5QMYRLAFuuFvwAB1pbnrKmpG4op08VIkMeVBkzVnLdWjvdnI+eA
Yg+f+hyeZt3bkIC7ZMhLdvAULS7H32r46a6GX5GGpyz3jlrPUSuiFtCTQ/TRF+UbS91liZEE0E25
mV7Y3ZAj54sgy4vfF3hE/2/nS29kNh3dPtGSEhUgxzoEIqJuHcsjyv1ZqLjwJkuSTj+wQHqPrevu
o4yqpU2Lh3oJEEX5awhRfgAQZ/y450YgcsZKgFgvDd2VyylhRqSRVBE00FNc7qfb+anA6UyykbIZ
hsst1z+KntWqNDejti5+dFdEfhyLc7tOAcVDWb29MD5ZIwmgiqn74Qozoa8upuXW9BBAeuoZ0Lgs
CZdmlMLcklakgx2Q6+SZI8iCPkIyX+fdpeRBsEb/bIX9/Moo81frWyHXAMx1sfmiXVshV+xL2773
zZOQbHqUrk8ZyRAMaXaTVr2lpojtI7tSNjA1dBpPr9ojzLEEdBRVgxVqat0qDV+JdCW5z48A5Nmz
i1pB4UJldeRq8T/HwTnDM6AEc2TcteKH8Oa8OAkXHjE+e5Ld1TWWm5xmkAxFcpILvg1mdUVRtKoj
1WTvvIdma8AOFGQwN1/uLhgzpckg8g9Krd+0wpiTN5vupjEHJrs1nhV7o4OOUvOv1XRN54x/dFMG
X0Q/Pic9kxG59VP4MKjuke5qmXMbuZyeFdRFMzPcLfKEcdOVc4WiJGqCJAXRc+12fbvbbMsrgrs4
tB92mXi1YjI8T6iOV4GieBov4hmWaz/p4r64jxe17f3k5guHH7ldah6p+//rGvwsJQ/5jKJzAqLY
Ph2Ut4fkzbJsMFOHC1FcgzELPs2nyBR6VAM0umEZ1ozP9RD/psPeVY6QuVqwcBkx6KAY6STcR0hS
XFTR/RV3AHDb8UvCid1NsuypkRjfly6OvCXk0R8BtpbxpvPSilVfK/0OtAsJ16zqUGs8N+2Pg9ZX
3NXDPoYNaYlzxVDTH734NFhpFCpwbXW+9SbJonHC7637mwPxGQ60QeKCLoGVAtpYFDdCkjadHYMG
SbDmJh2If8IAgGkrH3PGs9ZoJhzI8Ib/e7537Em5oejikNhsDP8T1TycT2QOSAFr/AMh4nNdmwxX
oLKs4n4eOYnqOMC6vhNMFJDwda6oIkMeqB3G45OdCQeDRaAXThAwHxuopD1pjRyrGLdy+tDAmdc3
WVv640NtZoXETpM9b0coc4Z+BEYckNKIAo8KdyZBHW6aJor1VLuYfFTVQDIsJ8NoJmf+slSJT/Ga
HbXHONSmKzY1LiSSoPEm/PuNmwguXcbhc2/BAqlMUSxpQfeU59wyVZjC4e2QIm8haNuFnj15cRVn
c35lG2Qp/nO0DJjc/vHQm94GaYpNOxhphAWdX5Cn+lhm98XKNO0HLFbR3UuxA2BE74FPiBce9Qh0
lqb6Jl8hxjDuK/TsMzDYJ0dFTnH/1xPBssZGUPCv8uKqNALcwa2iB3r4HuwrxVkrJNUtJpwY71ux
l8Y2PRE2rDHb5ND7csnYP8YDSCkeN7Tcp/L9NPiZQdEkTzcDSRUXZucO+jcivKLNhLkIuEHk5vZK
Z9ifhtvznWKNi+1Tg3x0Vxh7b80eZZ4HGpkcxnjDkkNSDOP9qF47KztGWkb78zb8DrprPSlHxdFL
Z4arpJwU2yR8GL9wxI2hMGkL5qej5tsP4uj1MMPGtXo6FG4iwByeq8ip3A2WdbXX20dkePbG9zn3
X3Qu39jzQqrkGAJlogr1oHKGGuuOWdoBq+H153VHzeMKNYouNB0Gv7po1xxmo2CtVt+G80+pyQie
WOWVN+vn1Sg1YWtpnX+izSYoOfQ4oC1DIJ76Qjr8UMgku75cVgQ4GibJhI60lxYHoITDG0RGYr9q
vHMTP2utkF6TA7ARztwfqBWyIXLUZKFNHYKDRQmoOxakEIwq1P9JyPGQtdBhYaRTQrEyVv5W2i3d
cyZGBiiZMZ8JwFCSLP1zAMNgRVw5lKb4yy1W/qrE/cVru/0bh8RJTmCXAW2zdE2wPH1mLBKfKJnd
m9xFC5DbKiH8LUhmAzQJlPk1XV71aejqJ2ILQ7cU9etoJPvgJkKMEmgz+LOxOdLpBGY0fynAVGDD
7WPACiirSCUWAWdPNcXMKOEW5LlAcFQR62AR6OOswO2cJe192XIt7s87/XuTe/DuUaEhXqFnQh35
Awu/JvBHMvFWoZ9HC4lZD/M74wM6T+3FEyaz6Pdu++EJiNQfVW543SWsgLFQYx76GoBO94m+TG4Z
QM5FLnXJfrG0Yf2AT8zjHtFHUfyMWCQIf/wBgknZJWxekkwfySDMSesSpMFDa8sv7UVhNysV3CFP
/IsdZEvqWsby24W0BM9/3+Fygvuje5AFusnf4S02vmDC0csAyII8nt5S6R6N1qzP2MKiHdzYVyxS
uWuhEmjlL0ZiL64XdMGDSfRKRrG+lHZBHN8zv2MPa8vek/In886zR/UXW2F04K+2Ch8GHO4HGvoO
KLWJU8S9HEaJrKGTJbwCJ+rxEXlMHa3RZKjXWEofkIqt316GV0pDjVAhIGh30jqeStWn3Y2e0XPL
sud9X4pmTKf9QFPpYYKkn4NaCijlx3o/TeL8u+dU1duJDZT4WVRGL7+WAbNGiZzEXUDvWxvlrzZ4
n3ZlTG1F5wXTGPUPqdMVtD0viVRhFlr+02uqKuNtltK14aVqWYEW3u/MSqNvbdKz1uq84yYn7zyA
Q9n6PMw02e+WQqWuUogXnDKC2fOW7a/KuF5q36yiGeJH+rGJff33ecxqxbc8DfjJxiExJo72Vp9O
nCwHKpuSoIflc7bn29P1fyyuuNbpqW4mlTRRyZK13PWi6yM9Ra2aBdmzsyjud//aQEvpvNlh7Gxk
3+JJ9BZKNFok3ZX2jwzkapxUdNBom3tf3pp9EFtAst4hzgM17ibx9uO5mrgNGvCKKsUM9PqtoH2K
4mlAePWR9IMCUCVnf/tsw1KKYpd/Nm09IzfS6vqVEBQbLq4j8thFgiKZ9O/3pL7Pwh3fqAadFMXe
Z6hURegbDOkGwwGBQQHmQU/VjrfaFofpXNT60eQ7BSixHyOmSDdV0v1Z+yPe8sPytiMYa1hD5eh7
SPBqYQgsfAMMxRrHkFwslH6Usahuv8N1QArhLyXeGqyBVThZ4X1BhLeIchl4w1IOrmhB19XVgtDx
AWq3sRK0i/2/47H1KnUPAKJ2Gz4WIcyjXiG50N83DQDLZdhvFiMVSCei/x+67QGYhWcRbcyAVGvh
L9P5AcyFNrXOcxX4AejiG+szhldYZAWIAY96Yhn3oY7FoMZlEJb7mBk1GBtaex3O+rkTVRfhrQD3
15dNz3UG4559J0xuvpxRA7zI6WkXJL3Bnup89/pHy4yTJErGp90sbp9Rde6yjSJfbW2yZWar1PGF
WKseVU6Mk4Zf6Kmyku8tExg+7WzW8zEFC5HMDve6Z5vyCIo7guFdzUnUWYtgfMFa0tXNyGUpJRF0
dX9+dmreq+dRc8nIwVHmrZCRN+LHFA0EGg6gicn+Q74Q2V8/ktQFBh5HHOppkxD2K1kgtzsSd6SW
7ChXlbnezTrkpyh9sN8EQZFVxCBq5UMqz7XwwqltDayfJEvagOtmWDbHniLfeYYXfnGSc/Cvwxpt
dCtm0B/qID9bVZORMXHQP+VJ8f7ZaVDB/UWX+1SMI1vgdRFBTwX+owmiGRfAn/AjBMf8zRpecljv
XtLJGpAlSOrJ80O21QEN00W0wuLvZgcnPaSGYldjdFQMW1oNPq6w5HsHliypF9ZSzncNzfrIhZUF
kOkbI3Ve7k5aGlM25ASL7w97znFKh2LQ3zMLC2DlcYJ8apxdzXeN1o94/FhC5lOKdtiWcq+KgJXx
wj3lk/n3y/Rt0HDNiwwDoL77ux7u0AKzHxk/rELjYza6VeNKA7Zd8aC+iAtlH38H1hzboG5XVnoC
T64AnT5F6A==
`pragma protect end_protected
