/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3296)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPS5CGEjGX4+ULwveQgO3KBYZAxdb1tVYsT9vfi0CpOwaCMTfzwkXc2Uoe
D84cZOmUT0TC8mWvkTfLf3+FacBeb0U27/rfOmcA18ARR0ThB90dUmUGmWBe3ImrjDPaNiAf68uK
AFZx4SSszmHfpDaXnrkiLWMUcnpJavjBS9gddyLGhXyrUEtNNsUSkHNY0ygJ+wUdSptoWotAPJFe
JBYxOvjmhexsou4c4/ncOjtG7rxi5qSsOuNmdX6xZSdhc0Hpy6ad1lDD6Y/Kl681VitoUfINdnqT
s2q1NdxwHBcFmgsSOZsTvhcgW0pVFAcmkAggHJzYJlwcCkYvtINP5gus1BZxxbc9yrKQv0dZlEOI
SNxj1R3s2TzymiODueKzEdW5hc62GaPLA9HqFrbBmcJAqeNF11SuckD38m8nC0b89BkVRIZEA4Zm
bvB2gfG7yr/9QOO+WFYqATSbCNfLHwTcfDMPAKt7DQtEoFXrbON69qyqaXlStxKjH49Incc9BQLk
O3QDbcsejtJ+aV07Jg+6KBiPLIldO6b37OBU91sucJSp3k6oRpmmSmezfET86kAzvyMyscqXetN7
xinKaoDyGCsiEHwAtI3FwG78qp6dysmx59H0mwFYvoemRE17k4Q/lkg7IAYW8sxxrwrJxjrGU4ef
HM2QH3h2H0OSzFlesUxlb8YKmQO3B/h01Rw0gWhxv49KUZP7dAMGz+rATBVLhrbQVfz/ywRYi+JI
tgur7JsoTY+AvkOgShJexJQOatuGJ8k3x8P4Jt6onvi8jpXmRb3ofX5754sYvC8RIb30NEbePzaX
/3tGeTb2MjOvkcYZuVOLzLtcQgj4sPWJuNQvRtj/9yEE4VeFzFduhFhOit/aUQzKFLXgN73v55qv
G8sWNh9zbSH5WgDzEyUwJc8l2SNLqQQGuNRNSy9Eu2w/nntzCJVot6POUvlaWZmmNgEZsW5VT8m5
Yzepx/4lXnP96F4royO3k4D3CSQQXwGqW5HuiEuIztgT2RMDgJyhdP9QIcWlAbhdHS42G9qOeaDP
HZOweTdAoFS6UdbRcHeUUD1F4hIZ8xRghfbZBUBGuVl7XACXQICpAct2aoLcJE7CWDRSm8z74QCI
bP7VuwfqlCtIIVkYI3Rncaq1vmU0dUD8dV1DHukhekvNw5l44skxU/TEj6SGBCXGn4d6nyseEYtq
rY7ppuQzPcaBDIKS3Yw9dTbp2ZtdWw8hpbs26HQnhhvIDt3v3ycrA4PhORZ28FA7MQ0Hk9M3FvFt
hL7BYn2xDLEHG+qByiFh/x5gVPO+bgjZ9HmDWY//fQuW2hCQg10UOd5lQMvnOZSBOBoVQtbpMZTl
ZOyc1FNPnrkLUKT/kQsbq42USI0WAB/Y+A12oLpOtUYJDRxKwkZgrMBsSQlBcW7OHIzvVhwjCRJA
nJHqDD82ppJEVa4/n43GCDTeuaotRDJ8BNVVphWHKRxD1w8yVnYABzr3/o3ByqXrahA9AqAGKUhc
8leiQy3X5ji8HZCZMxYkh6d2a3hfn9tvEueiMcWxmDe4cyoRQcvKq43th9BXowO1JVcQYmhBcJdB
xtsUOBPM/VQcUc91bYnI/D4oyRM/1fBncv4/38EPRRqs+crccKLQBEzpBbXiGDFPhC1JRCnMSY5t
R4mbqIm/PV7QwSjHTVR8AI8IbXGqVumZLrAbRdFbKz6W7TPYcr2CezCbBZUHuAjiDdQtz86CtiDM
AhXYN/fYr+6cOsBezvvYOQpboQWb5puTjKeYNgw0uIxKyr6pEWo4wuR2HfV7H6kYKvImDCRlw7kS
JDQlCAsSLIPPyO20bDRbL6bMz6FGKQCFwUujmLL/84wYzsGMFjryUOCHqZZtDHEos+6TpkQtNqqp
by3LE6S3UcYM0gdk2yzPo9RutGnJncd5++UayxQDkaaQ9FRmnkaR7WB7FqQ7TCLSSGO7gF0y6zhr
FxYIauF620l6sOGH5JJz1xVE7GwogW51ot11j9RsNZqeghAUjxJceRXkwWL3jNIl7jNjUyonuXXk
04LTB+cDCFEmsv1pTbDQwMnRHvcZ/+NKhbhzyM7+oXyFaJbDQKaUUj7onDgwobtWwDEXnubtSVuk
ZJ/85XLoqBN4vSI5llRbuxzRLMinO1zIwd9kjohxXRHtaLUjwIlyBIGgl1z+8Bm+Hz4VluNcNmUm
e2uf+YeBWU6q39FGaZ/MnjsvtLTs/E1qFXM7JMrwNjyRfTMtPwZmK/tLK35B4tvGs+NR6YnkuGBa
2MRZkrDvkHk+neIDFUOLvvjcGrQx+6aFuj3JhzuF7edpPRdrGu3xhSsgRwtxllo/4rLKGNvWMAf+
n0t8lJqVs3GkffdnMmaVPjoQyoziZxoWSe5tf2B1eO9ra8D6jAFpffypy/6MOVd5U6bBOAfW9On9
TCPZNljJnc5gfH+irZiHrVIRM2qzRUVR2XmeNnvCdT1fQvtiTOt9+PRDLUGTsyH2/wEel+g5uluR
nXI11Bnn0r3S5aNXLm1+/bTu1DlmGoJfLE92tiElVCMvtLGL6WZxnxVL0NJSOPxatQ0/vwmVv9QL
tR324qfMzK9plt8PEYfj57sruup/Ng/KLibmMmuyauZMrEpgPvAQ6T8Rhg7rCIiKfRg4//b6dG4E
5qxRHvfdzmxdernHYuJsl5fen/p8p7f2xY8Xz3A/ymtZTq+ZTIY611EUy0kHn2aH7p41L5jid9yQ
O5OboVLsOEyBDYWod4w2ZcEPbLF8wSKnd3qDBLVDN8kxu2yEHCnxLh4lNqE16XT4fNGr1I36PuPG
zg19NxvtvPnwDZxdIyWrNz3NFzVT35ud1dVNHHe/VH9fIpbBDbsAYKddsHtHmQezUZqH1BfLzf1P
y5dnvP4alTthLeSWV+SUJJ0Ru9cQdM8xLAbZv6feBSOybKyQbp+fa7jXs7ncSuJlDSZhCHqMcGwB
6JbDAqxju/ySEcpCuMsa6lc1M0lUil26/ZtKlXhsnOmmEFxGpNx0/j+dSkar0lV1fEjYCvcXUpTA
OX+ZySb4AxJvfBzHSHEhVYCRbClxaVBE8pi6wlAtZA7c+mXZDL8zowlFuhZ9dg7poK/8OXricBAu
Ldwcm/OwEc5Yl50xtKbuDUeFOAC9SmEowfK0cG78JyQI/AOr3ine9G5ZwmntmN0UTjYb90LH+o9j
tIPXvQZHvcXmJjGUXiewqLtRoyyBPfRyRGkxsRkmfFMcrL+YGrgIXap/auYPVVUi2dE82I4Aq85l
TUg4imms7uJYbXEzY2RWtJixeZo/B6gJ6cwmDjS8pnx1WUXU/yJCHAZsUyNa/+ia9ngouFBetqtQ
SCyePPcO+c1ahzZEy2CwiuxSBClGJFMrdx/ITIlM8BizbNbQRgJQGP3LWjrdqi5+TaMlujs80/wa
uSxugR6M9zWR5R6+PTHU4ejYj1G1vB6axnEc+rtbs0ISuhudE1jDCT30MRqPJXYRsenjFuBHtFz2
/7iabyEAqTbmfD/V5uXX3O8G+jbY8WpI8wvr1o26C5rp79o9TZpkYvJSIyYy8ulPIczjIFWCeQy0
wvwIgMfHiz6OPDuIOPNQyiaOP4X44/K7ljQZMo+O7xF+6gqRJeqRobpgQvR8W7J6yTFqo4yjbJ6l
0dieUlZ0CiwdClvqgAzKR9pVG5Al1xCYM/wme3b09SrNh3sLqKTctNbGYuDQkyrqFiP3mBfn1poR
DvOZwCZMjyJlQ7e7R0sEclP+P4AN75zyG5SCMQXJRdFkyDM98N2tggVkmEjLZORLI7wZmJApd8xk
3eklE9qSI6802mxOXkm3zcBX7pdc/+V8vUEZkSJM/ARVyDvLkIOahfw1S9zIcLtMG9wOrbxptjW4
9PlaOCeNv0i0byNJMdbKVDle0LS78VqGm70JyzfAeWF42rHW5tvPsLrDtWuZU1pLv2ew6k6gbUdB
Y5EcKFFzmyjy7ASktFsRDxtlQiR8mjDmtRdSFyyc8bIFp+gHYHE64dJBNDzkSCjt6YsawW6QuaIL
2QypMtoihB1R6vH4Z4BDHpH12Rp6YhYAL0GJAS1MrxJ77sLpbspOWIxW8QgxpkFjf5txNX65lGtn
Z0XPTxulU6JZ4ctRrfpGhnwNzjD1SeHq4dSTTfNRLP1EgBtSujgrNVfeOvbpdcpglA1zuz163J3l
ERBBN92zLxsAf0GdaELRLRhPBJ4ckGr4ua7mKKD+BD2+n9EgT05dXhuD4UyWXH9GTgi1M+d/jzh7
O/XHlzMscPRoGuiY/TDXduJNl0ol2wyth9DRLQNKUdOCjsu1cUy2MWm/OUoeVnwMkSRc3LA1G7lg
rCXtvVYgHM5RFOl6DbegxcEZ9uWhI+3Kg1nuPcvku7NmD/PhTrCZ+skspx+N9sg=
`pragma protect end_protected

// 
