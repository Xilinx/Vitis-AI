`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+GzawGdEcIuxfE2xohKZ4YfAgNY
udze0/JpwAsGtIi3JEG+f9Lc7KzDtVo+7e0axUtpWWG2zchF7YBRjZ26kg5u4E7NrejsKmQn4oFZ
2qTRJZGb5SJ+gdQBQzowrZ6DlCm5Ybvng4Y+fKORBe4O+BxCB8HAkjiHJvTxpq0VwrUrB2IS9/yv
BT0mW1nWT9cr5BxcHY80c1SIh2SWvSjyo6t8/Uu8goqodOeiB13w7hFPS0GPtfT7TgJBs7CKLsW8
/udu8oU6DrbuaGIvqyuhYDLUdvSeTbI1yKjoRhQTbSZsmPHD+BhP41ztTmXP8841D9OmucONcw5W
nz+qYscJFHjEhiUKhmUAqYkFeOx6gBtDwl02bgV/Ehx+qeNvEQTnNUoIM4joVXJp4gaoplybaaqz
WdUgHp7E3LhMlCdQPeqf8Nj5N9P19ksN5wBbu0jEHnSrjht3WaSC6qPemy9Sr43xjMhdDx9ezJ/1
nufPkpxOYsI7sQ6EQjS6u2TVYeZPxaRVbT+3laEfCq0eAwdSzrW3CJGDsWwthmo6lPbJ8Wb3/KVt
R/zJ8hNfQTOBfvDGgTVQ4g423oV3W2xKWKsSveaJJUqIW8WKphZAdpDmegQNbKQfmpQd35V54l0q
LtUTWCmDpsvFd9SGBmXXx8kx+8wZSIq/ivgqw+e9cp7gsau2q+Rn4R8TYRrBzqAPhlKVd7853295
32SSmwXW4IyftXavbWa3BnI5g6TndBfBwxhWignqlcTflqrXNpDoG35+jWPs2bzGeZRjvGa3KqLx
wPbZaixTEV686Que47d+YOKipqEkXstIZG5Gyel/ZHCK+fGhRmiW0vjlvzON+XlLa4l4P+zk5VH4
iytKfZsCHl4ula09h4TkZpDpy803UBSkDIyZiHNntKfRh3xbB5Hc5pjCLWwz9BJqFjcr9O/yWipg
V2TUi4HwepWD2YFCLpfL86zlimqlpM9kAulT04yBJROok3Gst/AWBqivWXlHXuo1HTiQjr9RM6nV
RFm3jcIVTi6h4HTn6+X9/syeTbiz+737c4dgzJre19HG8U/LlwwnOV1GOQVwAWMUVFaGPoBO3Zbd
QREvHaV3gWVdO7q/bqCuTPhOZZILMfTPAaHgSaan5xMlur7H8DAIScuWXtOtni47FGgwRohGB33U
4N1zMwRN5Gdc9cGyyb0ySUVCW3nm/tNWeGcfneJWl6LCfuMCu/1RU4LTngesngO6fglj/b43l26n
h1m4CjSeEN3tsnF1Y6+/dFs8VXWQ/CAVtiD3Xa48qdrd49gNrr0lHVNz0gwsQVQiS/xTcvz4myek
nFng9MDPIkBtj7ZbmRFfo1UgxDsgjcwdSAmSKqZ5ZjxwVF4wDNds6Eu62oB3ZUi0xNk8GJKFwrtT
xaARO46B/DyKwU3OiSsmhyB9uQ/bVYEEoSn0YAUZtq8WkYzuTcjk0SJx4sK29Ov+pHC3117WrOD5
r7t1mCgfN6nqxUzbKjcLEGC52znv87xrn0zfLUISqvhHsopJ7aYiWSUtydr1YVBDDc642eE0Jp1D
5s8lkdRykhqqR++0JtwuPPdNqtWCEIdD2roxcSU8h3shLzLR4o1Qn1HsLJ2ddksl7e2h8sHLIQT2
WvXzSTV0PN8yonDtiQBX08n4SQt9E5aUIOmShElMEhP3vAvit3bSBmOz88Twz2sc4Hu7PkLwbzoh
6kAOwCJMKd9eTC+ABdTzdkrfYgEwbLq6+WzUPJRoFx8jEq+cyiNzqINKzb+uFq5wjLKxOsRbSb6g
MDoCZLQ18oqptNKqpGUKvScd9/Ka8YQ+Mg1G632oZFre2esFzXSpm6pKi+s0rVtoXGMyb7JoC4l5
4zPO2HRJKNwjI2VFXQy7uRsFqJp9+VVEEeVDCHMg5GVjIhFPPeemCZv+MQX3o6hMHUaju92rMpHG
KoyhZyqaOnZER2vrutNUuM3E5tIsIRP1o6TSFxvZFLY/ogeoFIAYDj6y/vnGilW9zdBRFO0wbeHj
yW8fCEt0rUAkE47Kba+O7QenGn85eFvTRMsyqKyqs3aSY1GVGUuKCNrWOUs8LWY3ArGjJu3ckY6h
YFGK6JmrpJpxXKnK1TYagT09HViwVVFSx26b94SCh/iCnMBLAZ1ZY6QXVvEPoIaOpv3EktmRkODv
S/LFDzauATlgTU7y2sImrQGhmpsuUxZs0xy48MjopeWmcE70j/wOXm/0D9BwBUl7rjZ6LU56uSwx
J0SN1P1K8VLVBc/cuQDgz4+ZFjKY+FlwbwjaqxPG1+G/c0dc/M97o6QMfg3YB+Zi5yt8ePTL8/IV
R053KqEbk318bYPKJIXzsrZ17LBgyZ+E/yBD2vjzLxPHtQESn31/wzfivjqcR49UwtcKpO53IQqA
eiTV04SJKVd8OLEa9nwmPQK509dhmNVXz9DR6n9SxW+2xoamcWyMxEgb7i3QsClVZl+vVyoyXhLr
QJZ/HH/OnqRcX6X/e60Gjje9x2EwRoKSPNW3ABMkTvh3aPR4stHmLdzmTQzt44GM6TIUtf3tAZwS
qRoSgC500FjciLOHq3a5J8pHxyioiOcsXJIpkk8eMmI7gC5geVnFC8xOZeWnX15JHW4+q5fNE24O
tXE99tY8FXlJYxYYqFwAiGl16TNxABVJ3bGs2e7In/UiQuKaFtoQztTLbAM9Q7r6s0m6EUd+uSQQ
fuCGslbLcf5c6ddEi1sqlDCVOTOce4li+aR4r415N1Z4pwA++qBqelSNr3wiaW/4chbmrMFYw36R
Xfc3bdygZdipEjWSYd0IpKAvojZc7InJeH8ja4qhwnKGTFIZ8056u80ImND3294Z4v5hSSHDza5y
NCXuFWucltzibM0gE7yHEIkADK0Z3XszFmznlop00Om0/bMO4xp1V5mcCH2+wmQb7gzkcZWhcSqy
6SvXA316iLzYfylly6g0Ltpi4J2ghI8DG8MY9yMLSXbWAOpWNG8k5rCPpNiU9C49v5Al0XHOFBsQ
ZUvTGVSeMnfyFYTVvfaQizYnYK5D/KydxB03Uso9E4gEYg2Q05BZlOSGxna02vFN8pMiKwrZ48Jx
BAO8yAAKiLTzEphKZxaSHowkoHsc9ccjWv/aMaiagwEo0caCOTGdFFSYVBgpSRZo9bf+7EdLX9X6
8rXT4cqL4w1gkkBOplla+jyUdbwjtowpe8i5mfTQaDcXLcMul1Tez9gGVwVHuSu4Eh+qS/hykgO1
nyStmuhW/IfYuHWpPNDtA9twd4G9owy2PE52YY5ZKhMldBWKGtNrZYQLhsl6+lvFqXsgN/vDtZRT
Z81dMUgQj/RK7vufsLsQicUqLLVf6bKdW3B/SHN+pzA/os39tz0+AL0Wlp9k1L+/v4I4eDONImIK
2EEmH+vzR0TU4krF7sXNjJUlQ/OVEz3jAMzh8d7Ly/Y3ysXAvxc0pnxnDLHcT6H6AKGOKWsceIIp
odHxBcmKbV/pLeTu9BqrPd4pjuF8+Ds/cVYj2PSiOHjZvc6eI3tS7jGW2au7o1sUnY4KmhwLVBXI
BAIxCPB/pLYmW2mHhLilpsZib/hyklLSfwM1VnS+DUFM/iD6BxX6OyUl8jS0Rh2Cp3fyrprs6M05
hMPumSL5QqkRaaw3iIcjOF2psTnw2ysY5wMfS9rW9vJ68u37FgiGN+yjXtEUXjNuYaC439scIHC8
anWcxyuY+fCCbSNajggCutrEmyRzmfiZgPyhJG3BLtfC+Gc7t4Bc0AY4LQ9LcHmQiESGATdBkXdq
s5XnvhgrlvVV52znpn8ZD+QiXqA2wE5HVfhwRnJ+NT59mGglaFHcgCtCIOPNk+n3S5AbcWkMn9GG
bm0WzPjklCqPNHJe71d9Nl9jMXQ1ZImRCm8J5/YkdP0yoeiUGDEyit8Uv7kvbjEpXlKEqemASdv8
mfdcK8qKuXS8hD2Sj2f34rBctH9R1y/vf7PLjF3JkI7nWeFtn0eiPP9S92GUtMP9mxr5WCbCWFkY
L4frKQimoi5TBtyR/g1Vqvklo0C7AxD5/OCKDyQFo7dvG/I3XVSurSo/EZNtusZQPEP/YuSK0AFL
2qit2pZLSFMP72XE+FN+75LMuiJacrwKh3fMdwIi7eZIKbDn22xE/BYmmopH+ICMdg8OMzVQPZq1
Eaa+UOiT8Lp7Bk2OwRkfJukFyWCvRMDHDoF0G3whG+lbGAT5tf4u2X5vdoJ0TMqi6tr/g2H0dHEm
U8Z6TM/pjJLTEnhLJ+uH/tpYtEcfxHJqEbxlN0179SBq68K2V2M18/Ix4h9adrS4CHoJCRzuCBtv
wb2/U+P3btpcVDgoG4lMxPBHB/pZGnC/4lZP9uyqP7cfqudU8glFEfsoo3NE761ax+zARpliW76L
aWz8J+5DL3hnqieaxuQq4TYeA3/2qhbEaPqk26qtWRc75ENv3CmA0mWvoJR53S1CywBQmYhqTtxQ
ye1zR0VyI7ahXinypS011Pc6fZW++YeSHgysLdNrdsebAcKHcAn1kUWuKA1B4FMrRC2MD2OOkRsV
H1Czr2BNAxIseu8UJOGa3fuGtIzw2NT3APDS2R4K5DaQ/MpL8wY0JETrqt4jtLmcCEK9hUUTS4FM
ZO3rTbYnSc8jxL1YZ6k+DZlNyvoqY7AAvdBq/L3zsSNlwvTNrPY9z50tx6NJbP0FRO8+PshDOcEO
WKTYwltTgNdbmkd+xiqB7nlts1GYzpQc1N2Mw6OgU9h1+9kUXgy2dnCMSJyMFHCen5wrl5gKIm5M
6p6U2maX8Xgg3IpIDFJz8Oq9k60erykZIuTokVBbTzNPwYXbbhhjOG/Y+SvhYLZR3aXKeZUv+ekR
MBfOzqey8tFLRIfJsp7Rpo0LYwXCYH9QpnujOatQhZeiUbW31lX1DMmvVjWCueo3IpQt+9GCncLh
6XCp2GqXNGw+uMwweicflkrtvBgDXRhawamwo07Y1vNcnqz2G5wuleiJFXcD/1wocAmEcf09c5yd
lX35aig0oSyLCocLhbi8woTC9E/yMZiZxYAMI024Q5ErUuxdqGZKBg/qa8KGlGPf+2nk9nGNlSDw
EBeunSnmqBkJ4gafCOj2ocQZtavopE5t0r7B6RorrP6/laA6NXANNoznxWVmXtzjfKCtd+nvte0t
PrGCgBzIdwRhy7DPCLaXh4PskH0BI2VUQ2QnHkQfc4Z22uCtaQJ0+rP8EcXyAkGcpyQkxU0RAW6B
2rbylpxlsiPhsVI1oO2aLQaboNBejT292m4QtEQ4rxVPxAH4JaDnqnPr1MAC+mo5FntLoImBAjn6
wl1MN1mwwykGNQSUuIlTafUFMsJZyxp2T1JRaJiS3RniGTuw7TGkJtJ4BF8JbnINWpb9wMbLd06H
oHzFU+nCXTIvNznYgjq7VQrJPy0YPATc3ew+YEGYvGfhI84ZTaY/w/URkRg0R5/NrGhuiREV1YRH
jTdi963DI4xGUU9b6R7jeEiGjmUBoPPNXfDRhfNvH5n7OBq9cvPsCcnE6g6Ssa1qD76vSdFEsIlu
gUxhMqpAUJlaGfZT1zL1FYG7aPUIGS3deAJ5hvrXVjV0g7CepelHWcE/aKN1m1bRV/4EMrXKzLUT
KkiaHDZqBFecCi3AfBuJJ6PIWBN8mmEasODDgxbg2j7k9Qj+Z/ruPDUV56ybm621UB5R3zn4tsGp
EoRsgbxkW2Ml0Lzi2ITpNgqFw97OPELXi6HDMOZ5uPXODRmmMrJAN0TImfbsAyAe990ZIMWbBAoQ
ywVI0ql4T3Q1h06v+nLrteDDUX9q9TuyW+kaHm483kTcuxgB9BuV/4HWJpnXeQsbtbXSkRE/MfJE
44TY6K81q9dOSKRwpgIgPzY2Db83c63agcyk3ZmtwqFHw8nkmgXTLYSEwIQXwJTUSuJEHtilNDgB
p6XGVynp2KG0WfoiRwCpClzU8N3xQXUX1SBj388mt0nZLJZM6Gykvbvh/iF3utfIOwumPjiCYuYx
Aez8tVeCxzg2i/3SV2i0ZjJz1V9GSst7B1nglrhQgqW8sZPlXWqIHjTu1FQaYPR0UH4Pmivg+dbj
0SNaS/Pl8vE5F802sUajXhXKW4Ukl9zKwtYBnpZccUarAMluKmV8aqrm+4FnTsGmEl88SSUiv5PM
oLHZ99PdcaqEKEVTucDDTzhRVl7g+bLACnbr0+dtrhempjJJ2zwonQ8X+i7RhkzkQQRcmEa4Ry+4
+v1T9UfBbA+3rjHLTlUFPjbRlCakjcYB63U5UqR7aopuW5ciEwGL0kvlxKwdqVfk4BqiB+lumuBD
iiMBJC6os7++v+g+IxeiBxlbRmQl4fazE2XDiirARu7Vz6FOf2c/ygdEa4A+8+qtIZI3vDlBMvcf
DqsA0wEHTQSELrP05iokfHgNnweOhT1teWTL7GQuPsQUVHtz9OAfT1BOzQVYqdgDxrscJy/HCXFK
xpsQbcfr1/DV1upc0tG9eTzlNt4JGTbSxscsg4NT8AUs12z88rt+sArR6fkE3Gu8Btm3rjkg7Ik1
dK/Kf1iNmeHpUk+s50977FYmDyvL2UlbjWUge8FS45peGWl80478TCELhb5RLkYfzuVVZkA+2G3/
IDunPA3reHHyhFDy+iHe2/yUgL8AR4Wzh3Zzle/QGakd2pO2DEw6ATUK5A6VYwHeyYlBZXuhtExY
B8SQaFaW+Fk8oT8hR1SUa4P33SoZAjnNUqo2ycCaUEnJj6gV2anP77+bcD9VmTV5ss/tVvpaF2V3
XWH7QH8c30phzJwwjVA4QwacCdwQUSjBM+ninw/6zmZG3pynSU2bAK+m1d8mitSVgNVey26iGrTZ
6+8mRbei/VbKctUzBzRdzAOCUvnUa3DneEKivQCuZ32P2pVmaUvFz0xx1CZR3CO9IT9FcpRZIe/Q
TmEQJzvhpZqw5achTwGU6dcmADhDOoweBPQZngxr6TGbsypsK8ZtIXo+y5hLwVm2AwEWqKhAu2n1
nqGPSn4FxTvkbG7C46ptwqIQY+TnZsYxBoNQC//i0AXkPv+GSl/6IfhjNL2n8fqnfb0EIsjRa7EI
t49g2F++gWPQPK04jNhtA9RMD6FPxlGCfU5S5XPjw6u8rfqb2CjtXbsKq44mKfTLfGbLVXBqhIG6
RTRNwLVtujQXi0W9qFW9Gb6EmhJDPGfHdCRBNDrzDdMNn3O4Q1eT4aBZlEe+0O3DQ0LR/Wls5XVK
VO8m0o43G1oxcppp/Urp5SnMFIcW+3F0ml1LXvsgOJRdOngGRllCGq5BcBXEVzSTlzt+q7WynvzT
SU5bgNpVZwrebt/h7TB28QNTTet7hyJAh9+3ekbAxpe3ImSY1eHRjuwK302vNt6PBu2gIFTNUANm
XlHsaqs7hMPTC5egsoV7Z6yEf5ZSav21eG8ER9U+X2Vfu5FZ4oLPIb8FUeRwVjVTbZBq/cVLm7JQ
XS2xAYTVFpBdihE67rHhRS0Js6slTzNT8rQBE595SKgn36I5YRzLiu8mZhr2Hq3AkxbZDfi/Ch61
T0Q2WkDg3l+x19Zz0OQPubglBix7YHPH+elewlgvEGktyTDUBoWgifvkk9Dov3NYEOEzcQRLLP9Q
y9Dk0rlXH7dKxNfn7NdJdl6N6YR5nTqRllrdCqGzCDFIIIqthhnBzzb9qLGWAhOqWdbadIW78q/v
HNVv1e5Vmxe3xcAcVcAgqxh+SZO97eBK16yxk3vADSuYTOun5Znue0YITuBaFG5smFOHCnaTtcF1
b7EzhUAENThOCY/dwwdzg08QcKQTl7E8YR47Nj433/LlFp4gBRuBH2AZm7W3P70Ua/54fihsA8EN
jlRZJzT6yrhU4M8HolFd9lnLGAY7RdUCGm5Y0xezpeWGrVE8YAn6NnxA0motcuOT6FW+HJvUSnKm
BBg56PcstEWUYxfJ9sF3qqAExqnqM1uFbN92DhLKLyTRH/mg+UANSGta692fNiyKG2gGjwOk+dql
VVwm/O0GSsXgFFlhz6yCqHofknmPBDqjxFWlEFsL8HV0CNGs2RZVX4TUL/3PoG0thXQJ7lpnjEwh
WJM/o9V/2KDIOETsqD0CXyHUaxEXMYAMT9xi5V2DRfyQ1yFR5AUeBwdEKcGzqwzpdW6NLJ5wby6z
bpbYuAzkjTVN6MxxznQN6u9R9p+ofz5ec4GHgm88BARx9c0dJYoQCa4eBjRc6dkDps0+TeyFj5lX
srCVRpRDu6fT4d5q4OQKGR/yKZVEa42C+cf8gbR+q+deahwzLVXJJHluA2cfXEVknmsfE/iiBxOr
oOZbGoB1N71Q3CSw+iuRvnKMPcyr0Ej4HDtyBCsUc4rzEv0mXorkpy8lGmLI5toqE7IVaZdJYylQ
SdI6kWrm9Nh2z9GuKJqhf48LVKYIqcwUbW0kuGgImhpI7Smx16z7cMbzDGdwOjJOHhgsGCb1Af3x
Ec5t741PRkCSF4NW91ta7AhxXNynI+d5s2a1D+i2Fe71I240y49QyRr1M7WT2noXenMicPPRUi9Y
UjAi2WC23SVO1bl5bO3rQkr2Y80N3/VumyLS4aV3i9wjTmBpo9D5U4SQwaaR2Hl5svrvO/ny7+a3
hjulX64m1MXlT1wHgS8FS2gY5WIColTX5uUDjwDawaDWNw9XZ9rH2H3cUF0vbR9xt6A3jhSxHlD3
wUEc0myJNjFc3nx9zk2istCAbVb67iFRysY1lRPOo7bEE9r1fdHEbtvkgNp9j8es0Am0phKrr/Hp
1SxzvOJ7wRqCgZdDG/TM0YZUEdOKYv8Dz9aaSjuxmeSUTpcfmFs14jtgMFAI4xlAksrm4DefMiTN
TnKqyK6d1PbmmsfrDoeOTgGmKPjl9AluFil6MYDP6ihfIpoXBI5Y/WfeMRwCZEeyYygm4D6H75IK
QLa8p4g9Fb6Xi7RS7Vd4PCui5xM+2nCYbK3SlMWv68N//qRszunupNgPIfFe10/XjA2Tg9IIcXfh
aYbdNDdgWmwPc2PfcBoxzJbKO8JJlC6Ars+NS+UDNA2imegY9kXfWAiDL8IER7YbBb8sgEP0PY/Z
2JdfvVITAGBEGAgMr3sx/R1RpxkaCilDBUMizal6voUkEg9SK5V4xDd9aaN7Qz1KKwyeiCdPmqc2
ZC9i4PEOoL4vaJDfDi+XYBEB2nUmVvOKv6Ph/CPFIJ4tPjAQg8JQYsS780b5B8u46w3UExCntkIS
uEr6HcWicE56gRB3SFdApmIdP6UjPBCDyar99CTA0QeoqheiGlgz67Wx32UxC+NQroffpR61thAk
e3HaTx5m6oIDBoMGj7AJ7hJ1JKBKho5p08ecIyUnuz+M77zvPLH0ooq9+rfFsH8djU2Q0faXB8kL
uu6o17DmSfAwMDnHK9fxZyytk56WKgFFHAzxz50ffpB0JVKHxxn8NkMFY9W5bzkoeGNprP+5AuCE
XgfI/dqP/2MuNWrMEosKoNuHlBhKUnT0YXRDAz5MgogOmlo3KP2I9dqBvjiIgq+/LrDOFZ4K6+JN
vBq8r1+riqsA+eHAJGdTjeAjcnEy7IHkRcZDr9tgHXnY9+nfnjQWnpOpBrPB5Jgw+OnGwR5FWs6L
ToPxc7zmOBdDlx7ydJzrvpVjY6fwK1fe2eDPOvVZhlxmLo0v93CrC6qrWDah9jqdNX/UeUgSyujd
B/beSUzOtQSBr1FpWzH2fRMdxmbqWxfkYokbszW2Ei1RMpOhr1YMJJXuKq2SYqsJktIq//K+HUo9
jW1MgJvUTfUYSzXkBssyNWL6evPGp7sut7VKcsJXK9GYTB/n63ckr0vdPyJ7U/D+f8J7c9AWuwsZ
Ug0c84sQZfX9e+z7an7jVcU6WGW7uMcVpfaDgXTXprg1wf4IHAQvLcus3qlmgz8FTbkA9n3IGx/D
Yar0XP/JrQc9DxXuQu1y2WDjVQkbWZT7lh+2g1s9BehqfRtN/Rk1J+ChjBzcBFm7OvsPGu33uRga
VxDyZrkCzudZVytyj63CXnnEOaC5ylrtJkkXi4ybkQ2rFL34IapJ/8+xxPx/efGpdszioGmplu43
TeluK1dh4LWWHrxgkRkqOQu0Snji5SlrELmmVzVekBJGc/ZY2SC8dr8X8AIMqde7R4EtglhXigY2
YvzGIERFXhaC0WREDGdiHXRU5aLOkx/gM5HFflGUTjC904/u/NfT/wIKSdjdIlvo7CS2Oi4Fc5jg
WfaL3W9Ld6C2DPWgTg7S0CgoTFe2VDRx7tsoeoZ4fMVbv9Il0hLSFdBbJKT5YvnV5I2F4x6LpFVi
r/VRroMyLLSBbBzuVoIOyPkNd6K/PQTiOicb1ys3m0dUyHgxYecWSs6//YZ/AtxX+SXjiK3dc7H8
lwi6FNOTYk9/rVImCQZtAnTmIeHZLBvJMF4gq/wOKshSFpJexO6WnWuBZYwKftwDEd1El4b1t5+g
1OhaInH97Ct8OhHkZpbXFcmfYru7YNnsc6f4yGeLWNEUYVWjtcGi7tqPWd5EvvbcY/GI9WyV6mSE
jH8KiPYH7JkHVYThPo/qJfmLlOreP4MLsYwbTfpAgJIWJ0Nrecneh0eMrvQcErMi1GrClap67d0w
K6MnyRauGhGQhqtCxsV5OQsLc+g9aXEqKyMe1QFgidakA2CbeiWcvp9wNq/rh9jXjPfEZQDwBCQw
L8WhnqN7SRelbcHrDTckQx+r8dLwojfupGBN8TusEYZ9CvLGokDd9lhPv1/Hv+C8oGegBAs46fbO
0hWaJXoqld2qSLG6gdJAmd1UeOh195ktoa8fPS7VQfQbFNb2hYQZIYjufRPxwJPTzIk21I/TqVqg
MooDZbzQPkR/8o6VV2QDmJ4QBwKEUyy+3bp/KFvw0FlznuJxzIEgnbOAKYhiXxOv3Hl51BBnzcsm
k6naKH//SpdFWjmy3YKTLVZpsaST0m1H0rmxQuLfvXU4T46m0A8vobMrj+GVr94MvhFMfSNgiyHs
aZfrOh1/nlWS55QLxwlN7PrJAob7xECafRm61uV3+azvTjGjsMFoHixzdiWH4YDqzg47LE/jaF0u
1GYorYCpc3vohomSiGhev3/SC+zD3vqZ92+qg6NP+BfqbWsv1lHwl8hfpzDbg39Mbu8qSmm/kUK1
idiaRHjIu4RMnLGMokwlhw/QtN8RWSwTncrcNf4i8w0ufdoonimoyjscZZDsLt+I0D7txiD1iTKr
I235tncnaMNn8hDO5b/YwCyTebPr3ZVAPQO9uG3ShnQMeeSyOKQeEjojDS6IM/+8qEgW/Si9n2VE
I1qROXw3eUXBdebempd0tYbqjXPydP38sEn0g5csx1w+AZkJlc8IfgUjVAyAL2kUvHmjDPCf7LYc
31dUREzZ7kmABW7ZrUPK7i7NEvY/51ahwNcGcKfaoaN6QzUdT7mllmYKNgANNpJH60z9fJ5GmtsU
CX8s/0oA0wR5xxuyHIGxXZw1cDxWh/N0CETGWyU9FA8RLNi//obKwDbhumKu7A5/sutTApU5cGk3
i4ZF7Gj3VDQrfEtZSy8b4YotLtOazY9vgpiLNaMrNaYodOp53z4joGaZ9zkT21/4rlj+2mAWn8pb
g47JsgxqwPTCcxrJFWBFJc6rXq1FxW7232BwZSh1UTTDzVjYGuhIKb9awN/fGntHTTdEPZlkiCIA
5/KVWqwvrPn+vM1Wg447dV1Mern7UJ4c0NH1vs1e/UQ90DkGIpMlFPSg3COOrOMz6iNfFwn7VpqB
q67dqDQL8KNvW1fQtnmHoTlEcCk0khBPo/GpTsEEKr3ldJOjUzT0g6UAhvCLHPBPCB5TBCAENgku
P476sZy4d0298sHhzqzUy1JDhInlnEwHf54aoIm3tYXJQGDoma+12tZfpS5hN0qByAvMu8JvwHcH
2PXRDoP6S9EEi1Lw7EuDGEyqap2EQCrSdLjHBORvtKgKZIE8r+kZz1GnzqWXizU6P23diNanL9BW
mdItxtGDPjc7+7TvFVdJkamnHVTCUrbn8q4ogaOIS/DcD87wr+hzxH2RgUYYl7K1zqNl/u6gT68F
GafM1dRUh+q3uAMIyXffCm0SlcFszra6uPCxfZGapDpTOeCXimh8QuTYHTzPb5NQbAEsCfileDTw
pHalXQ2FyOmACAJ9XzG0t6Z5AqKpU1EAVh0Uc31vCcUZwLs7Ha5ThTm37xIZ8vduonJ4FFIDDKDD
C1SWIPdmowFEnG3H6GhgeRmdaB1F/RpVBhowu3Mg5shwWY4xyepXFT+ryQ7it+qlEKOuBrdEwcEW
JIhfDnwq1a/NigYEucahRmtGrCiAmqiXvwW6EofCgzM4I9e/ohF2UMdJ8N0iC2CjrDv8BzCSoPw6
WL09ioRY7Um6RxcAkDvxxfRE8FSnE4/mhmbat8iDOM+XTAzKJYLLeYFlZji+9Ndd/K6QCUduBxeQ
iUDelmJMrj5ApVIDOoWPrXD8Sv5cUgiyan/Lq0PPpWQLF8F/LY1WTvhBn54yMfT861nvqNDvyfIx
48jKBgYFUg7d+gON7vGC6hySrgnRA6MLoPHj7I5rzlREJBeZyn9M9owWiLS95kRZSa9w4WX737PW
XWRoLUXyW+idcz57G7inNB58c/+KkQpss/T4c5lW8M6zcbDYJiqPeMWk9KTYIoAek3tBtBWQtOH/
jIWR1iL4z54e/IUE+po1/6QpyOrRtxPPNf0vNZebtRqT5ryc7F30j1s68WlhgOqVCRLsvP0XlAOy
Fku/1X83rbHuKKXYBcc4V9lCk3d7EqpI1DuKCGW29kQGsz3BUUUZrojbmDBPXyG3NPpd0Yx40qWo
6wAD+JTSbzej6/xJFdFJ0Ulza8Xd0XL05E+83L3SgwjajiuhGEO4pOxfvDPTga3qXq26OXX0d1eF
tQ9JORrKPSFJN3Tb35z4xmTUhzHCiG23F6T/qYyMoeI6CgrqhU1dPCXy+1dN+C+/D7mbV2Poml+q
9SjVI5GyqyMxPoFWto6DFlR2bmYLj6eueyL9LtWwMVjZnEv/S0LMxwy/qx6aa7w5tu+WLp9I2AqT
x4PAEIYRFDOit6irt3z4FxSsAumSOn2Ei111Q9J0hRd8ORlgc8PkJSn8AK89jt3MpTM77LnmUsIl
YcGLI72RSmC1ssqq2OYl1pyVdkcAYsfWybvpB6+5jE3Id61ohW2IBG5EyvUp09ML/8lVBJ5GqvGm
/cJS/tvwzwVxRbdkBLfZSp7WdytTxVVTVqA9TaX+54ODOqEUMSHPX+flfc79BNjiz5/SxJdjKF5O
wWVGXwpYlDn3qPhUGwDT0R5yt+kxY4rfKYS5JDX7wsPNXmnUaQQEOrIy8TtWOiz8vQigRBI8iG+W
GcYr0fXl3dmJO0tSZaEM8iv68ABdkQEFncyHhDdUgfqwHYWMNN03/ZQEGFl47xri2M41cQKZCgKy
R6ZFsbLs1n5/Ob7m1v7jkmhfKo8yS5Mia1LfwmUrg9dsmHqBzmwdbibFXhFRLM07TnMVJRJtHEiE
bV6RdirFubCcKmu7xM6brHrgfk1JgSu3a9eLcgmwHm9dI/6hyNlaG5TyI4Bb44RduYk7EVsUHxrO
kqwVKmYmCLtsnH2sU9N+UUS23MtwRO3BKRj3KlElxOM1R/TyBbI5fbyU/0on2eNRTQUF5Kicigxk
PdXNXle293hyVoOy/n5EdXOxgtyuuAt0oVkldnZxreihjxfIqzALtP9A0bvxHYybEIHlw4ZTMZcd
+F9Lvz/X+oCWOya7BglJQQtBSk+KP1VySFM3qnCJ67Ay2D4xT5NkYcjSZgeDo79cQWTM1dB9jW2m
9r4nF5ejZrQkEtPpqdb9VMltYF/kCcg2K2qKyc0ld/jJLw3C4QwopwY65Pbts1YkoPwHJA4vYvyr
yWGs8BPrUimp6YKbXKGGIeFNhVAOf22pxhK/5UFBwV7e6NpmJcnxxInLxIMOSBfw5onZWMSnBAfQ
gh4z7LXL1y0RaT4YXJo0P72R3PGn7dEC6CmQ8JvIFZ4Tfpfeug53hxv4dL8y3zglXoamwaqmTdyd
eb+wQF2HGArdMpl5z2VYpLNG/EPygSa6e/uc13VD69u4j+I/vQdMh0Nc+4y1OMwEPgmdo+JBJQXJ
Ypcsg3wJg8UfGEuDvfCWsoEnWYcnEwGmAbborun3h3Sx9allEOdQwRC1bm5DKFQfGLVKBqPZJrrF
E0V7p2SXXQC/X6aVT8pk6eV9AO2IM660ZivLJiKCp0dVj1ynTyc500d8ULTZBoJxN7T+zzRJUyKY
lhhox3AQNqt+lUNlGhXix/f5mXgmp+lQaWh1ksj2a8m0azNm8gg8mskfxJiQSj953mhJ95trbmtC
QHm47eMtI4xX6SrQEtSVhsmba+36AdGLw+CHnEgF5VcE0gZzC9OwU3Dam8qBWF5werR0Y6Kmtr11
oKJ5ruDWtX0aq9uCzVPseEEw0UZfi4b7HOgof2sMrYHYuwwdkAq85KGHerZ3nbRe73j0pkNvge6X
AaJrqUL2nueYWYitvqde1Ojnl4WjjNPJTpPJxAFplbdYQNANwAGFnoCwO8bbj61cJMVvQGPrpNsF
ddrspgonEksVoM+j07g9gnQVK+Op3d615XgNtOiPwqQptFGkHnNrk3nDKQhCIZ4ajKXjqynygfXj
bl8kdfbJWQXpnAxNDTXo9JSagf4OJsJKMVDHJuWCojmYhSzIQ+97+Guv/e8voiA/BA9+g0B4WRPc
O2d75fkv6efgswOq8liGEoVaKmjhkasB7PdPRNZEypMVpPDxow4I5mWpQgZS57BY0CW26yuKgbDQ
ArrBWbGK99qCAwnmDbId11nQ0cLxGI1Ttb69iWAe2lQOAm4ML4QE9xdcCPcWxqt8JCzTwCTgA1qz
+2wVWvAJ2qDmisWFd5Uy3RJLGX+2OkKWJF5EbNo+7nNf/UNIKOfMhT2RsNKzDYlo45oZpazcQvC5
zBFTs8jzd5lS9FVSXpdn9oIoxBQ9f70VOSoimVHEziqmaDCVnK8w7TkpsDSgXUHlJUDOfGtOCGeq
Av+WxAgPCjOeZN3GCZk38UEhhcg7jhOEbTs9pnix9kSRinknnSMJnh/YlygwZkGu60k3Vdiz8Oj5
+jqQZIO6HDlEyXzU3SJRlu7PswHa7fSeO8fBbapYNiPE8cPuqSLUKDj0l5Zu41Vm6ONC0grJec16
oCsZqdHN2W4Ro1hE9DcrvVgzT7T01Xvh35ujwkoemx2h7dsB9jrfBPQc9mf4cPrVdlPLrChBC9Ek
H6XdN/LsrLG7tP6pAoYPnAPE5MejxILOjGBsH1Pu0NL0aSrjLpU6vkx3ZiF8tD2dPa9R7sr9pbxb
/wYAmMTW7i+ok5zWsKuCan9q51WxUJRN4uMzPlrCYk/UdnzeHB9SUXxMOBnHgSugHXiLUE+qmbCn
5RXXA9BBtWRFlKx+Dwfgyb1HDGh/WsqRG7IanT/nZJK7Oq5YC0xE5WsRFd79v65SuOd+NbsaOMa2
3/dxy3YWockmFEsJIr1x7Z9D/uDKvtkNfnPysyL/2K6eZF2SSy+DuW1zRp+0PCjvhA5APQ4IV5s7
vskKygmApVrMSk/7VI4qMb8zGi5ia88o/NzcMPPVb1PMC9WhkAKu5PnXXMqz2R4qCVpRTbmNqvTu
3Hhrss4hxrcGsPGUXrPz8syh44A8HnvP19aQEfP1KRRYcvnD0kdVqdSllzSFpxUkkxCfwBPLE7xE
+LsAHp7sgr2H5tdda1dJN/TIhN+qT9Qkl/ugT5Ja+5W+gYYGhKWLJxuIV6kf101t4LGfLCZpSgGC
LFjDQ5Mi0q5v+KfXFJWANu3cUBKRGUiFDRDsbQKHs6ZD6XEYw/8rFdRKGx2AqMcAT74VjlCXuLjT
LZpl1F3Baplp+iF+hmDm2h20NTFFT0SipDSKlnkBni8G2t0yNOXdABsZUbRuwlts8Cnzy7T9J/lQ
ngOidXkyfjedzfdO9V2YrBW0YSMFpr4NaFb6SpR3NmRkzkR3hBArKFPX3Ttyw4TtwEoJVp6auNb/
lnddC44rnp8GdmuUzcrC8p6xOd5UMoRQkLKLEx5VpRzhPr+HvJhlMy3++Jyg9fJxFejZO0ycFW6F
4mvQA1968ZjSzSfAoc68dYAPRP/SAj3FvXmcnYhHumkWCHm250yrRGrtURox55dJUDjTMIWynMUJ
Fu3Zuj+98sM5j4m5CIsEgRCwToWgki+QDbmd6FFoyFKqnN3BW0Rme89BX/V9qJ/OsEZWoxWcnylw
zIvgXd7gZrtvYt7CmO9QGeL84EtSuJF4KOzJRPL85MhVq29E0D8nofZ4rZomtHFkNrgqGNXAkQH5
943QzQOnC00J0dDPPczCdfM8MN6EzxSXMZe8hPwdCmTAyeHYsmWpncIKGQg/MOD9ZzMGNBFjFZso
zgC1NQR4e/V3u5Lpx66I1dGVD7Z/MtvhTiwwYJdm12W/DaXxHuW3uhu4GTeJj8VQk44oxVMNyj18
Pi8Z7P3jvc3C6Xbfkl/JNz4zlaIIEIuPjpQnF172IsIQV/vuA6BljgIGT+IvShowEojmxvFsw+IX
kZgwYli+cefL+Ewi5hKc7xyLgPysYtwHshuT9XyQLSnAdDWaRKgUqqjvXbA/FGSNnLI6BgJQAM55
BlIaawFosjoZuNAT2yqKkiUzqkGKtDGtWMg7K+D/zUNMqR8vRK+WH/U4CZ7QL0a3V5kHOtUDWOh1
w2F9USRNDbYQFIaQKvxunjArGq2GijzJ5pZrtgCA5NnNyCCL0cP1XcA7SnmNq5Pro7MqXpm5MgNY
grCBRCPx1hVfryq9xHTZ7QVRM6RqLsYrUTkleiy0UiTFoBTb8s28HHCP6zFfZD6OwmZRSywgvjPD
DXXS8BqJFp9KckCombRrUF/pX1EOJrhzC/BQHHyNc2mx9uYRgIb/A1lZzhvoYW9DNNHwCxA5SeUT
onM2/SXbm7r5ZFoBqMY90tFzAPc4FOg36vQlhQ3/vY4bUFXG3fBpbjIonI1l+rnfiZZWM4MvV+T3
QQlzlkYNGz+4spO7z26IX0RMKOpZe7hAUWblhdwVRMFAOqb0yCh6VfsK2HtN2GLzR4TtAHJYYiF8
5olRo+h1qtZ1hrfcO0Ql1/t88Dg6Bb/7Lr6QATWa8sWEBEDC0MasmRo001lLyqAizb0TU3XfPbwq
OWiwJQAWwS6UmuEg0Ck0MHkuzUv6er9qNdMvXo1Z5t8KKzlzb/wpVfBIl+RAw/l3DFSMXIUD6kbu
BA0Fd9ieIrXBv01nqCNpT5n/YT4ZIAGXu6pcTuDoCWpW8I9Q0BPd3JWSbwWCDbRIKz0KD/w4fjpy
rw6H6Y6C5/KhXuc/49DbAhliKSyYykoH5CGRYq6BiZfZ+Z0Oq2KqRUwmspiaS9H13A1gnbJoDbNG
BgzzRfZ5F/InBJSnGpNCdg6D+Y2nCfnPymeWZBhNduN94z3jyk480xsQ0LaRAVnuRsBBuZRtpYyR
kPpuOJ+znlLbnBzBlqUZ6RtN4YhTYp+OgcdGC+qWvBExdC08siospQ9epLPn8UdWlWv+WblZD+Ky
sz2Y4o0vrKFiy1ICkH0dwgvH4i49L8q32sxnV2bDd+NL2jkDTSLIQoJnoHUFVXt0+6/tXmQbfSm8
BeBkVGMOd38ErTRSRYYrp3bjT3GJELOuQHoOJxTD42JY/6qeukVfDchEv6oJtk3zPVuiFJde5XSG
uBjLNsDfNg4OH/8lEn6ntftA2UjrFWkXgRnCJQkiQ/UN6ZQ7QSmErZe7B9+AguRk8iEfbSNO1BVC
FIq53gRMsbRjlTGXkC5yeZNACKVgjRVTsimsbeHt+7AS+nYWX55t26qH9no6YGYjryeuq5mlv8yS
R/uvElUIUgdVtUnhTNtG+d0GuRXv9IZvoO2HaIBM8cpqjjLzhYoLP3IwH8v8y/wM/88mSVwV5kJv
9qU6kBO0VCPUYbT2HL5pF5HPkTZMiG1vs7H/v8Ble5Xlt+l9iPey1E6TrJO2fBiHG+YelyAid1W9
2TkXpqvXzjoVuUMkM5GbtN/Yu6HMRwpF6nBKmAWT/AkemhtE2ov9kRAdXGS3+GHIjOtPjbnVN8tf
pS7KAIUq5K6atEBU1GpY0WuqQoYI7B+fSCRGub+BA2/THYNFOj42D4PJXiaPeJDExQbyjUt2J3yD
AuYLoxq2xJ9+GudC8ytngDYdOY+m3o9Xz45Fc4L+yo/Vqq9aaMBFovVZFm3d5w7hgfzJ0cZtsj9c
bq1/ZuIIhEyhkzjXUIgksuze6fJgrFbk9B3oupojWFDwYNKpDN+6od6SGyL3bxIk2cp7yMnzeAHz
fNEL5lrS54KzwJhzvGdzyhFukLf1FQ9l1qjaLFJ51dK9fIdlCv+hvZIhtJRf0Gd7PTix7AR7WWnW
982VS1FFrT+rtn88jpxuDtSjEFSmIzvW8rTTTGp169xGD2RWK20aHJcHt482cNKUnUERBQ4aIbkd
j3NNbF81ORqq+Cccheo3p8FX0CCcyUW/0UgA2EI/c6Jo7U8OoKhhkOqkiiihnJ5yPMYkVB1v0KKY
62VVQiRXxYhlsfyi2A3IgPteUsY8SyLt01oQfpXIjfN7tVDYE3pe1HxjxPI7QOxLh3d9jkZ41Na6
J8AxwzneVPFdnFclJoBw0XNmHlEJdAdpOz1uqALlBDZGu0PBiYXSnJsw92ZFKX6/KIpbO8xI975Z
JhGJ3jyE/NQyhp9+Auw7q90KYrZ5FIk/khNl+mN61OWqXFT3JNT0ATQYWEClAB/rDyugo17BeSnc
h5PL16Noq5RJX69a8C0RCkFo7sU55m5OVMpOJw7ELkXWgLHHYvLkdmJNTEvL2aMJ9TjOiVBGT8LQ
NMEkMspYe33sTfFv1UlyZIMWmZ7bZg+hpjzOk2UZ6ChUB26MdjcUTQNd1/ta8HvfFIH7Kuy7m47x
IbWJEECy+jL+r+DHjyHQm/pvprzGu4Fv6AgJfHsj46V9bPwZDzZTMqt4Uk282wTAe4IpmhB1Mtix
xSQrSBCL40gBTs2g+TwSRsoF5kJy/W5X43AOJ/hVrHYjICG63ikUltNTQUlJK55nkQoaBJ0UlNwe
YaqHE6cefhI/sMkRuulMAjGmQW0ARTYBIPl2wvjxTimDkX8sZHlYP9qL8iuIyOFR4HSRayayoXoG
svmZ1KsH91zAF3a6nsuJYp84agWtcDAy/PkggFEXPvJVWkL+rQ5KWgrZKdDrawnww9HU+R5gfAn5
DCPEDePEoJGVgbCrytVcGF0RM/oX0r4HL+oiyEJWTmjcWuDgKZIL/keTbqV9IuMqe1KNvcD1rXVy
gpCE1a0BEwbRDioBgvpuLStjjrWyDMyX6/kcVX7tD68La6XuZZUeHrtRwH/+tsemMUM3lgL2BDLn
caR7OTbCVmwYLM86C7WQVu7/0FZEMGuJnvq5CvQFFUw9DbuUpGaIKFsAwwgxnyzmSlZltNRSg5na
XuuNoUXB3wJqMU7cayonPiscxo72DhlaftOmoKVZmNykbBoLTK8FF+x8rg1qI8rb/VR1r3zF4Ain
xoEaBXosFflaI7Dxi4+5zlTTL/SkzTtRRRykJRWmKZdt8EwbvH7Oyev4w6KKKHxOnUzi0Jiydg7v
ThFRh/E9HXac3JLCVNLwMgkffP3ej9pURioewqVetq2BTc2SuHL4KizX2klAUaL88vvqwtyAQUsI
cA31xVOzziqcWU2FpHWtmPUf4URvRZ74dslywx2JQnfUpD5a1loRXsLz4a61AH4zbWRobm1veD5D
VMrJiLdNgRNNYOAVIWL6XnUO6jmk2R8I2nk5gUZN9nrAg1JeyfoMX0utw+SMoBTPlJFtJ2NXxWpc
ucxNrOBNuUJ4lmJcGjdtTzd2qGY03pKR/rVdlojeh9faB2U/H3Oy8s7sSvYy6czMFJjmdnPY48+m
IRrdZvGZnloK5EnxLSU9kWaaBTp3eNocOMur4n5ZlWY9baRlrmgLfP4GTCjEKhGY7y+SvXnYrfyK
neOGOYLF069Libp5/fp1xX2XxYAlA2ze0D+n3Bo2QMDRKYdZKsgJYUswb50wO0xM83/IQosBHV5V
+Fdn1yk5XtN8O4WRPK9SL7Ai4cVHM9e+oHuYMl9nZyKmYAPsimVrrcKTkLz+eElSfyzii9D7rxR7
ot+YLxIOwdx5v8MsuQqeOBo9MHVOCDO6lNQsMMNdqLaMx0yTOfGxWPAVqIqamsOVV298L13eF6bF
My1NZp7Fh6OJ32J/+R1t7Qfksin03yOnzyiAGI1xn70kSghCduqPjXyqwgizgj6bayZ4xaVBgTpm
O9lE/HTRW7rqrcHCy7nyLLyO6nboeWA4kPL8iNXbY7Nq1rAyVDbLT/+sP0lAuOuPEhsbx6d0CVPD
sXBMh9PcyvM3whubmYJzRvRXR+YtQNkpR1QfxhDjTZ0LPF6WCFqRMvq4BcksHB4rEXOyUTm+GJjz
t3A2EDinJCgHRry2B+d1t0yoz6xlJLTL8eoj6ODAkAArlP8wDQQ4TIjfjv5yN4u4FGypJ4PiU3Cy
b1HgtR68nVHTytoGzdMqkgIGJDBxEGwRpeT+7PlZ+fy/bN1/eXqwXyV6phxeE/nE31WMV7Ip4kdq
dYHMod6+bWeGxbUznH02/xXiOQMSm+/iH3/CYGi8teQS5NUQgnanx8UHSrf/6mzmdAHaogufkTsN
25d89hmLjppzc/cFcMSj
`pragma protect end_protected
