/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbKPfJfo4jNVPLOLEZmuD/9YFJsCXHb/vaU+pQt6TullM1ODOXE6t6j+H
PWqFOgXR/As4eoYkJ9ajGTnNdVKLi48OwdzbveCFS71tevKNW21aMq/Yt1M0tBg331V4cLHcciju
HRmQkpGF63HGTY/hX3FTSu17wCcRyGpeTAFgYxnkqN0z7ipqEniFDfC7VCUqchY/Lm+PXuJckoom
rEuZP7+zpjsHeJrC2DYlqjyJAi9XOe8jQsYW6VeJWl45vo/HE+Naq3WWD8b1Q7MmvE38PyHZWbcZ
gwItvTWx/V4p2CQQ+NxcX5qKIRDDTzDArG0ybeU99KHW9YCY/2vL5j6aH91bDwEjkFXEucSDUbm/
Zoi+hIddY9rJ8oz1ZolCPohhVE3tbRVjfvoxxeTuPcxFw90Ds886mSMljZ/B26xVwPINklq0XPX4
QpB6cPYfBfBtbTpJ12m6cZFWg0IcrrGd6AcZKMDR78u85MZJ38YdwiO4KzjDl/BrHF+fIFX6yW0l
Cr/+KvhJejk0mqdeEXwDAWhGESW9VVs8Ymhkcy4bDSKfLfiP/RG1mwKBK/hPm+hMz9M4mBIXG83z
pYfKA/X26AzWzikSWiuhJXXxN76xNdgHW9yeSFhYQSF0wYhx2JdcspDOhsPwFtMeI86ASMmElJRH
SX36a521wwOCp1OI+rgrw4VJamirPYqYIwjIxisP4iOMvlx2pnJ8z11PJezQIWka3jSmpy1nP39x
i55q6Gytunf4vOSJsIGlKoI7/1+fr0qHSTlYlTMcGT7/zV5j2utrEnukJM2FSxdKgMu7MlRdQmbg
NsFaI1/XzZavMBs3M9tczBbgM6PEXIiyQA2hhhMRT40G+1RIDXt4Q2TEi9LqamaDONiaifqIMvgA
W3JwoeP1dFruQnEgdP8DLS5NsP5jgkhezsdeHgryUcpkp2kYArBrPKcz/EPaewZc3rtAMPdoKxBK
ZqKPQayK+Tg2n5hdthvwqfNSxqWIaT7gP98U5QdhPA6ZHKRLblx9U0rqhb345Ruc1qeE94KWc+2t
C6Ulg7Z/ei25Mcc/8iSzd5AjuAG2YRRKgdAgWN0m5mnlU8kstujgPI4FVdRBVYY9IQjI76qPF6cm
mzUxhWTuoLlQ75qUXMken+twoJM/b39/uEzBwG23BgFlO2FTrnPEMDmmTj+pm6eS7oiw6gjrcxdg
dsWGPqpSNF2OL8q+JDRrUT49G5ZC+Q3RIhkoN1iNqPcgq6VOEmDUM29HBiZBii9TrbT7ogy9QKld
yaCM+CqAERW5i1eyxPyR8cvFsK8F3XDUqCR0e4DcasvpWKTzzCT4P0e917DFyPXLZwvgZ72gZokU
KXqKEj7liUAt6Q0xPNjAismrYujtwypPTbVuHaBeiGMiJh0VFsI+AxZGGpuh7pmwCnCdpi2RcGml
uyjD7gzhxvdkll9ln0sA034qgLQDhGqiJRqfXO2KpIbXMLNiPCDpm4T7WwFLXED4UA1jREPNQVla
hv5/6dBGgcm9QqCOorimlGLWMhYxoHvvQo89P8+bTFJgo7kIGsAi265hxi+DDo6zSbG4zfxENfO/
6JpzIBgjqey6kZqAQ27bEojqhD4ATgemw3fiqFODqscRazu1uU0ophR4eDdky3X7iQh1vfj/+TuK
q5bDAdF7K0VB9wG9ltPokppwgD4dMTrHB9Ev+YVVygLAUwQUM7CLTZxjRk2MW/UtxzbbRi7j6LIp
/ThMOA8MieJYCSSayic1xBN55/qbYddxyL31yR4SItCXvjUxMsV/Ad4kMA09+npCb7Pz5DWyhcMZ
4LECTuM0Bho4xayEuMH5C1qmLUDeu57X8ZctuN94avSIl1dvIBdJBv7UB1XCTJrQxE+JmAfhnvPx
HR37GzAGnak87r6xEIJIe5qTS92Qdv1DJy+4+9tkaPSXxIc22e9faqlBzq5NZcUFDwkJWtXvECYO
4HUt2mFuaifP21urgzoN8Myaz+Pl5KIFgXKt/QjSMtbJ4CaK7bWG5DoOsLSXTcVudyCthYAOGayE
LHTHvkk2anmaXMk6TPTgXCn/ZKFJwZkfzyy2g/fWEFlMyxG34TkhpINmmrTy/bUpTFU/JpmusngE
j6mbhLmhlYlviS8mjldlsJok8YYsXN/U31OeJ3vniKOaZ+7tHD3YvP5Xinxq+cjUoiDQ4c0+33SC
ADVLAbtv6oXkEm4oIYUmckK6NGep1IdsDTqWeBQEjSR0Af1JHacDvmaUnXFOqZhYPnapZ8emieVM
mPotRTC9YQ/VCZvdOj0FjlM4FFnxyQMxhgZQ3fpON5955Yo0F4jjVk8KJWayPjGnhPnhscSbHG91
Ma885HM1JbLSCeA6+ROQGy43M3oXJPFtIQl05Jwk/IGi3axOd9FQmFjSKWeOkZbgh1D5BxRv2CXy
DoGHS6ihABohUY8SIIftbDR9nY1pZ6Hpg2DkYN3tqH6zURSdA2IUVxsfqvN0028xBTPCTvaVUQsa
+T0nUnko/TDUmXJUyWiM8sQcArSb1ku2LJm5bxrET0GWp6c6LFVQiOBg+vfwcCrGuDfS0Qw3ZG31
1tEJO1qnqIJZoyGLcRxCfuohJFRFnHxR2COLKrdJJUNiMucO1bnnzdknr4bTAq5NMnjqhA7T6EAR
bO7R/jBk/kOjrL/VctK3bK4QN6sqPhL5gvZdf9ltcBj+kbL11DvHa8Z728Ye6NvYHWqFBRk0Z6G5
APaJ1TKO28DOZu0AUIoTeRlvTBkyc9An4+m7oBIJsqObgN97elY6SA9RDdU6g4kl1XT0aG8oLAds
c2jewdf/rr0RqZJTpne0BWTfjxHi89RtiQDfO9mAdELg608b5ZOIulZR6HiXDaKxNtb+Lu/oPKVV
6fFWovFOJJzbNTTm5tmsEY+Dxuggx7XxJiahISAAaz2D+kUbV44QchgafZdsuBvdMFVT/0bmCC6a
aHrp1uRsMeqZyuGex9oURI0zmhCe7J6bQDpxAKM73oSzSSNFcNQzUa4Je2342KHDpi1kx8+eRyXZ
hDPX43VS7CPOLJsqTHO4aQQB2+rw03LioReTO3EIIsU4IAYoVqu9Bnz9wqmFmj1EqkNQJ4A7mUNs
LoqNn6ARjr+HlOzeFy5fms5ArpoPvzJzKN8v1SZcqi5FPN8ZQNR9ZrESpQef0wyisThWgvjEEbCF
88wlsOTAx7vGVyyPGH3Skx7J3W6kexHbK683shyr+DGyv1jVOm+teXbJVOJ494iC8RNYIx//xpj6
Zdwmmn1pjmSMJvsrV3L5EqBYlzQgXyA/8rUThiEBZW7FuZrS+PIR6oHN8dnFHpHUoe6MHZddm4zb
zKwhZMJasJIjsZ1ZeszncxqA14w6OwV+ntYpiQS03c5AJ8T7FFomgoorXucL4sZz3BXOIQI0HBli
IE1z+j/+tJvI784XBnMVOmgvXrlqMsR/OzJIuLvB3+hWV+RZmsPQ0UdXif2icHv717aU2/Bkh5KN
EaCcl56ds1wu3Nz8U9yDptSjzwqB4nqkqUP4fB5pK4c+i1pX8efYMthqLOm0y5bH2nv21CF631ly
rLoiEr4GEfo80qDQCbzL+eg5yiyjaXSl/k1IM+j637S8y75tAhgHWu7+Z5C1XD0/8Aw73IsdaOoL
WMIicL8w189w+czpx3k7//tUdTbocpiUo4KDn4gs5/1etFeDuIqzVZRk/2+siMLU6AguBZTrLatX
w9e7tVOk/siM5BPWp3EgdskkkOdQn9OXx05iPZHzeaIDKz0E3gCns5eaeY8owqbopr4wES6Ncxdh
rwnpXr+N8ffX3ZMiKwQZhgV90R9+W7NYe0l/VXgPOueLgIjBdDgTEWsdb/cSgVFZujiJ8XZSdnc3
4SRLR2IsMtA8ytHfUGE358vkqHrF9TM5+mfiqE/7xI2BuyoqFqjSEY95YMcli5n99aEThCWer5ec
OFRthEarBsqt2SUZRQ5uJCxCc3y3izS01gNLvPHm/ggvu64L3VRQ25isO5xhvZIwj5r76CD0APN7
JbODVloY9I8xGPNviboGFHbadi96v+TDNhs3Eqx9hs+VxSxlmRX051tmVJ6UT4r1ydAiGJP5PwPS
qS9VWFA26pYrlISaioOCz/b5GfKSorfJpmBfN/hRGVKysQKTKfuPp3z+wauiJqWW+GVnpFygeumB
xo8OOfShJyjYoEHVqHEOSVazuPHPQDLnQHRLKMDXZ2wfYJF/7t4XI4HrCjXdFHwI1xnmo7bAC6MZ
e6CcyAXZ2CAGGDmmi4RXDT5I7TRIk9xmoPBvzymxrlmxSCX+Zu6ZzZGaY95JnMwOHorUA5/QwAil
TkO3dKq46UyyfXMMH42mBQAWq3saR4/4d2rAx1zUacN4tMnerz5r6iiJ9D9i2jKqgnmL2sWmQ+qj
8gGGYlqJk6nGKydm3yp+tbZNF7Hwgop5XzbjmgrMIXmil3KBCQWM2ragOS8vAn0usqTYnrnd82fG
aYAGb6KiLR2VxvarjRTkwU12Ev76zv/T6M0owSkxtQXMp0uXhOn465/1LuVq1sDaIJ/+rWdUFo0y
DoJ55bAnTRHlZMTDvyj2Z6dVUEmJ9zaVWtgT5GIZe8JIL5tIwUD48YSXj5Aq4NdzrUORPBGX6k9X
e5yQDy/hndvyeDJLVqrFJ6471BSZ3hluIklZGBLWAXy1Xs1v3wJG3ioHmpG/0VKfXvTxpyMceqHN
nEcjKYaIx1A3h3UXLBVv9l34kkDEHyG4r23+NDsslCRa5l7y0NrQ40uumKvZIkuaWExtN0HwxlD+
iKNjOj1E7gwMA4oMQnA+s9Keeg25Z1cnyul4rIMizJcCBvpWa2/R0ApfAAPb39LIwwnK230r7VHv
Y8JTx2zQ+lyuNTpUQWmsNgEgnMFtocIBJKmH0BzAOD8UykDvFQSabSfzszPGu+XFRjtyD4sCrh1F
P2iLKF8mrBj6ldB4VBTebo91ZHuZjR2uz/2zCtiqBG6RmTeN4YEdgIAF99y2u6VPZVu71tjrsSNh
YTpvlGVCUSNAf9L/R9p9gSZk9aadr5zqo7IHvFSii//vvvty/CfYsp/skLvd2bzg7ZF2TFQeKlbH
UxsvRiC+f1wc8ixa+XqYtmtXGA5QvNIX+xCN2q0+OPAt0k49xpptXofDBv/5bN6RO6uI5GXOFnk7
izJCdesyxn21LxbKEwjLS/UDJaZN/LAueLjHd6P/hHoQQCVM1oLco5Z6FSlwaE3/mAh9yn9yq07D
3b8z9PaZ8NYIxCYDdb7Xh2ulAkkBwkSG4+8jI6o39W2IXT6qdc/10W3cuOYDgpRD4BHIjhkFiixZ
s2lBUZBUIzriMXOD5QxcxUOBZPbC3tgrAA+Ux7GpSYwNUGAY+12PvUNM9s5yH+xst3zrotRsoKD/
uVNXGr1c/ZL1fwYx9z2IMd8hAqquw95OQX8x5WLIxNmpMGgoCm18fCS0jJA8trvw6FO/1nZMN8Fc
EKa4NGsZgeTvfnsGTOP5ytbMkNQTilD5zveDs3P2Wq7HhtM3T8ooHXPjCJo57dRtl2Z3Tid2S1v9
kOkOdAeGm5l/Apxp3sMHY38POI415VKnL2YguJiybqWvNAb86wHxLC2/wY+UmHMqXP/StqoLhW4Z
s2Zarwjj2b7WtaOerfRa/wHRZPxchfm6OU8Hzjd2TVc466iaR5cXKO0c78hQ3ofWoXjAals70pBI
9lxy/aYhSuC0UW+viO8zJsrEFonychlSAMK2AbU2a/ssZMqpCG1aArk6cC+1N3KGPlkFXmhwe74Q
dqFJxpGfQdz3LZXARXUoZLfVRQM4yrNB38/e/I9eJnRVwGClyoMUHLekd0YL3ylSUPxlD9mp1Gr/
X9SpmULWkZPJVeb6xKrviaibzXCnezV+fuNPwcuH4MY+nXYCAgZzj+zW2B9BXh8qgm+V1WcLVOrt
GBNraS0I/+WjaKMXg9TyhJktbB8uLnxi6XGFpS1BUu/eOtb391vvuNg2acpCZubGXmYtnDFSQ8vg
dQudSlHC0SddLmO6LNpbhnsmUrc5wqFKX+KTFLkNQuI9WLBNznXHQxFsF4hxYOZDGHAwJ/XLo0+b
tiDoVN9/IfgVis7NwGP+pda7yDymaJ5yci+CV9MtG9bBMXgS3VZDF5f4S3IPKOb3JAr25fpz58Kc
8PvuWAp5cPrkWiKgbEXPibqDvyX+XBr0Ue1JxSCHe76Jp+HWmWEnF+cD8KBTvpE7o2GVrOVOvxzS
IWr8M7fARzQueUQKu/JBllNZcTQ0/MZU4mJk/QHFHWPX0d4kp3Rdzg0PkVtc+kIdNWRRgRik/Ugm
IImyAZteN3eIQkn80XKvBZuKihk3upk+IJhUPsST9IA4P8CUYqwx6xWwJfOdWPnunN14MWsIya9r
CKqcE8umz4a4nWalxU9EtfnZQD6LHORCsHL60Y+3lHqucFH72R91PX4csYjy2js2NJSJt2qqqrf4
TPhM2WChAt2LfeY4lgvsUF1xPdO1WcRLC2W13UugAL4zADe6f/liqv0kI2hY530eCwHzTTFH24by
iUE7cy4XcYbTQutYnp5QnzbVLO8x34eD73n0SxSdSYmcQFZ9FgsNo64+r6GP69O6RMiBq4sORoK7
CbCeI+FJ4E61DGO7edbsJ0AxhoSim/rn1X7cyO+fylOpp9PXgD1qU/8XoK1bNUbBHT36n+puwPgT
J4qSt1o7cFA44ldM++j+QwEhwqZRauOXqpzns3mhUqsZ6UrB72GvJ+KZ6CoxJpoHrz7M3X5w5397
BGk7ir7Xa6fadu+GQpiCVcomEc+kjX761hN9IJl9lj8rr/fo9V8ixAcAyis5+Y0zYWs+vFjgekLW
S1uFGjtXoTmYvkNX0p2wvrA9urIqlGp+iAAaa+Nk0ssS6iuwTDU00PaksR2n62IHvCFoq2pXA7gX
1Wtpuhq7U3V7ah+6wiaMw2KpHnz2VqTSZ8J++zaD3SXWwmc52S/z8QJFPUVYXluN/PuHsVnTNg+y
yjPGzlUlWLGJWmwMN5/VmCpezwkDTYDcrCZeOEWlCaoV3Cc0U/cGfbesaOL1PqzpUoP686t61/5n
qbLWuaCBveoIXSc0PpgZDq5igDjQRpUv58SAKws245nzzqyCCyhjRIc9yoOFQxtibtsjbeoGzkIw
Loy1JQr7BdJFBWT58Hmmpr0W+DG+tR+t/nEycvMUM1j0ajr9VvZIgZYrex+WbI2ueivCO5iq5aEM
6wocKK6gu75je4Y0Hw8TTIVhGEO/PsC1NmrGjggnoXnmquiNngra+nbng2c7x2SJ5VpXvICGOHpw
8ZExjn25n4GSVrBXaG9uKWNR0gJHyapi8h3pJKsUzQ9bxJ3u/Hmo/LiIfzaHd3AjaEPbWh+vJIS2
rsQLdhNfVtDKkkOVzDXEmkimuUqcYOY/gDOVL1nRFcqaNcCQUzrNq3evLuLdVgjJtuaOOFvPFjZP
7xJbQOiYPjlFgfyF+zHtduGBcu5UjQy8mKf6COrTm1+Y3p3oXBKlPNVO/faqXV/fXoM4EzLXTanE
vJbQZk3bEa6NWV4lxAtko4u9IQx7I0Cw3dxeTn2JkV63L//it/bJ85OalDdn173f149HhqsS3wHe
foKJsXR7New7FDT3Nlvkm8crs1WB7HWNrZfzmyLS9ml1NAmhnXOA9wXT6DLZBoTkxCO9KOr96hmj
GVQNbjWEdBXC2cEEzh8gnK6tRd3RFuXs3C8mEKDtyhMeI7bzrihtJYZUJAjuHDhKjXzF0pTKGNsg
gkSvgt/3FX9RSrl2cTmSia+RCoS+ID3OFv+EbOE2tu5OuaaCo8mmc8HpIgzLEIw4UrTAoqqhzY6k
NgDW+6/wYLf6SkSmY/qIodxE99/RfLzoqJVS7zWNcIMnOWy/RV6SVSJMqDp39delQLgZkmI9dX4q
DpV/yndqEFJyfFqxIp6hLbZrce0/a5zUpwPBD0o7+3S9b51k01xSbR9eJrkG4JXH8esRZ5GrceBg
G2/77N7zbRUAILA0r04wv/OJNihvC+rM4mwbM/XYO963yZe12gmsO4g50fifRPUR02LsqNgcrwZI
/VEZzijSFBkNi9QG5SjCXcCKhEdyVFi7ukuYby5bczzZCgCDABONdXYaDs3vdVFw5si6tE4vN2f0
pcwYK7mVQ6QQOZV3vvuFhPgEQZ6PMa4lxrOxs7BwbwA2Bm1+1ezri1WYvIwd4u5SIxkzxeA+XV6T
4nkef5aOE9RwnCPyVsiZzAIe/ENOkkPXOGyXqbBaZ3pwD5ezJ9Aa6HXcfJMHWZCXT0lFVdF8jqNg
3W1612ZaaRykQQcjHgfZJZMuaNaUHYdU9CJX3kCPDpvPp8EB+8VN/y+HM6VvWJremBWnAYEgefG7
Oaz94XR0rrqr4f4OAaZFKLRm/zEfh1sNliYZ3fhraJAlhvkG1hr9ZIaWBlFAa8w6sXk8CXGrEebO
rPmq9LZ+Hys9h2WbrP1DIx8sT+/R9qv0752F7WgDW3bcOJy7iBXPbyfDtxmxAWuK3ZmPwb/XXZTZ
IYkiA5Q/k3LM1WbqWsAVjVs7OSmjM01++N9uZc1dwLrbQiuNdLVFkU6D+FesjO3BXjf2POmWKjn5
I9QGO/W6uOehSA4JUow6Z4Zcx/1KdILRsnrDrj6kkjqeX46qp6E2FXydyHyA+alVtZx0RKQdoGsA
EeRmgxxuX64RFZY16n2oLFGgXvYpbgAVfWw2zCS0Rn/qG1jKMVQadVdbThyVbqomFrp1uEmyPykh
/1UlvuSM5jnVxHEJuQQFRPSLGB4QW11iC1526Oh/3MVUyGPGj9EYL0rHfpGwXhIjQFFCZJq40gnh
5n0lsRo8KkQ3AQWS0Du21yVSA2Limv6OPUF/UoQIPrfJ/LeQ0Y9GVh97ZqDSw7J4RkJlYsmQb1IF
1yGlZthi/iyzl39SNgBuOoz4tfzYuesyJnWn04RNLzKseqA5VMb+gx+A9neX8OoZQtbuVPoIe1vz
01TDeLyZHWJC2wZnNwvwiNEmF9Ne5QOXkxb2hkBUWY/ULV7bUVvGzQk4NA4gPbKzXRLmTN9EDhYc
9SqZRUBbKSJ0JSCPjtPPB8+JQhyR+h+yxB0JIKBtp3B1TZQAw5n7D1o8SaVuGFDwclpS9BRnMTzw
SsMsDYQ7PL0OY+bp1NOZYPHTeGBC4MfXl0SWTxVjJJGBp0yWmt4VhuiSEL9DYb4La6iaO0hnmBOJ
cxyTuhJ2zjt2OfbPuSUBfWSj2lMGUqP9HAq8PEngbl/DZ9DorqAgvIQy1u5gOC9SjyLpAXD5isB9
TPW7VsrDlpu7ugh5mArgKiowpw51dbAvv3G3Mx/SUyjB7h8YH09bpHwE49/DZAFvgS/9YHljQzuS
hyMYpDx1nwmt8JpL1Lkb9IpXjfriePUacbI1GRrU4uFvYuSJFb/ucB8Jp3KqWMUY4dGM5AkMsrI3
3IjNozhbty7HU2KDwHFMbGBcqW3eL/BwMp2vsFMpg89zSPEFeEFsa5DEXihHch+6ktk7YIMK7P7e
c8VkDGZOu2UooDG/gCijMrhlIy0GYkbQWut6LZvY4Io8lcLjJ8Q+knwqn9Lm3TFovRAvj9egHTn4
IFX6DXzZl3ygCRV1QMupTq+p91YlCnNYAG/L7s7ASJ+GlTxgcJHCWbBqgL1NMPRL3VoCZmRB91u3
TGxkpwTHXXbuqQesNg4zEibZCdJa+rbSqNaMJJAXjM43M2sz6Kvaa/J2Y/GAY3M/FJkqAHY5325G
sQ0pSt8oJwR2K/spzqqhtMu77EK/fu2+OTCoyOccUmvHgUb3nPdI9oVVCyrl6ZP9PiYnUMaihdLO
G4BlNu8ghPJfac87zRRrkWmt8hgzjKlYaa/q7oT2rG4fP7IbLDneZlX6GdJXIG4Fjg1T1Y/VmQ4a
2f7li++eQsqvopbB7cpe6kfCjnqGUPUKTGYghJtjdqJ34chjO1HS7OZJDh4OoJYPZqXx8jAszdE3
I+F/jOSZPupVRVH1qhMTU+RxQTxzA+hxyUneNB3Gw56jiFvgkgbXlK0VmqF68DEDEhVnr399vu5b
pm3LxcPoLS1DBs1OlapBEc/urquUg/nU/OU8Z+v1g7p2qsjCVdJotbcoVQ3UkwdGaVFVTkZoeXzC
qxi6QmNkj/zWEA3pwK2qEQqof9MHEcQ9MObILTG/SnDCGHRnKZblIPMjMimmFstX4PfufwjILkCx
QBChsvO6bgnPXtln9gJ410sXofbpVCafGfICxDabi6sFtE7LkBw7382UutshGhQggeZ4lx4pDizi
/shDTSDluaERAd7+CSk1wzvjIwzKCnvMBSbbmpNOiLBKf9U71zvllMgt7aT7l/JpvQpGDSx9qUv4
CdenvZWGxYW8WCAwwD7FUuGjMBiFPHwuGWP5EAFX/qqSmnOTIlbuWgeyZb0un63dvDE7EgxZvoNR
Z+LCiViB0b2kBSqu49IoKYUrFWapfYl/2x76P+h5xZ/lxRhOUzzdISz9WeNcA8Y9BSjNJ9V3UwAY
SBRl+wJzqrG3V8y/mK+vkNpuffmkF9Prl9N80ZqGK2sVpkWwO2vY2O/O+bnmW4W1ueF76d+n6GCc
6nmsqdyxgimERk2Dx3eLZTZ27BlACxXPVxyxOAHOir6m9DI0HEDlLlIEfUvXDvvohDLYukdY+Cqm
UUBDc+bn7RCIow7hmb+LUe3v7o2LFAN2d9Nrg1u9b4oclo0kzSCYhqwuzP/u1yRxsKSCLqrzTjJ6
LDa+U0TTrq09aCHkj1Y4v6hr8lsfCvC2DRw87OJ1MK/Mq7vIlI7+VeUp+zBkXFK56hxICCSfZXbf
OsiCwrpkSwXb1GFe0DbZXZiMZ/9nAnxrw6sNepvstRDQSamICpnGOMi/w8vAB3mLbNjHoNAAVsXK
wmZAFktOWr57MOTlCbu53n4SRasWvPc17kvHr4MX7XQ4+NY8djJERPIt4tp44SKltszdjiCwzHY1
I6CLB04bKQ6mRBL4AY4ZuwfSwC7cadvtUQt653ynQUp21LVipQZq8YrMSS6Q1wjG/8F4drOJoNp8
j66KiBCx0zHS/5+Ey1i4LSXdfU2Fcb2OdKX2BnLlMS1KzcicYgXcVB1cGuz38FaEIb2GPrm432Bh
5pfzb2g0gX8NscfT0QgaT0Y7byHK4NgvsQ1YVNBt7bu3e8oQajehDsv6vvFOBoR7Sur0ZrXV3u6l
PRbkW+t5Hsn/kjz+TpZoUySeMgmfrkF7VY0kGqMWRmyXSxoOXG5HXJZz3W1+NI3fC9Lp5qAGs9dG
FUcRxGNllCSRk9JkY8KLVL492sGaKkmaHdbXODae0ZnmoV+YLwQvZ11ufSofZfyWi5enE1DW4xrB
s0h8VaU7RlOSdNyk9ktn6Fkdg3Af8CqVPuAP1bG0vmE8uY0Q3cfLG9P98onyd0IwGSEUhDnXDA6U
5ABpEgtRFy0yrUeq1z1km/P0ZpBwMpcFEMnMO7cP6CvaE04IIYHxO5jENqVQCDAU13sXhpMp0F/1
4iIKTDAZoxZWz51f+lrMTPMRckH5TsVzLnqH+c1Zacmy+FwePzCf4ma7/Hh9YHhzXGViEu19BCDa
qhh1dvoiY9dF9PROJCH+rR0Lu+rQnowLJrLOAPZRXA8S+I9Afkz0o1B8H0YTekTLElYySB6aaZ0t
ht0h/o9HLCJaHJo4GaUCQ+KeKBeo44KnhfFokp9JlTAHsVi2VuwO2LTo483ybdD+IPSv81olsihj
a4O11viJejelCcJd3xj7mhm9W+nr22AQ/edaooTIkDSQ6HpGijJDjnaTIObYNevFdvqPInMlrICm
3+5DH9iYCNlb6uWTJXyQ7G7TO09+cXsQbWCsN5GJAhh8euU6zLVfThnlwTWxzt1uI9kIvd8a6+d4
TyqgLUdJpLT9nywkmkeRHO2HGZv67ssk2mcw4YIaluvyHFSTw7iRW6JsAdVTg9+c2dPCxnhsFAs8
BtDxpGtKyaZk307qheET+HjXvPnxZg8Dcik99pqTxtBbvKXMLv7Qe8jTE49vGesobJzz2JenZMUS
K47iFP2xuaI5yoWhACiIVJCsdOXLW1OwCHsE58gcMzvkyonHBUKYrUzZHzzTKg7jcBjptzV/D5LT
4g1vxJe/62ReC/lAFtSmhzHJD8EgCPSQyCQ79x4G2BIl/IJkAqbTO+5JiKZ7d1T64pvDhoyfk37M
mJgADJ8O3R2z1Ubgubr+/Jb5RVRPiSy5QtS243kWFdx+s+cTbJeUV2G1993X20VS/jvSmB4GE/bk
OVznYMd9tSTP2P41pq7q3up9s1hkF3AJPqzwfMESPrqlW+QCxcQskE6BG4xHSowaosPvYRVyZjXE
EbtDsme4iY5LFQqSMn6XGNCWgvzhBcYSnJCyh53PdyF9jqQTPvsijxocOBAmeDX+AKDCO0m9DYHq
TU4ZffFpZw1ReihKNINfA+wVCOa7V/EQDu1SCIyIqzJBFZGd6zykKVoKDx6TPzUoXbKYG4s1anSq
dnp7sOyHmM8inp1zvjst2eOFzAK4jDmAwxnlHbZ6E2tzTuXdbsAguNARwPLd2+njg8JMx9Mi2la0
JrmkYbclkIceQlfX4YXHtcvZgJ3g0izdFOh+qvexY8uVbwbMzBIJ/1RIUuLizD5VM7Li8ou6kgZp
lXeAImx7XAGIhDV5KFPVAVE1NgjInh1OPpfBZmwyCedmFry1JWQVLycVJ/ESbI7qvmRQeqvgy7v3
z4h1Xf4/cq8JL89sWUD2pWSbf/M1J8MwHKgbe2DGlk9jCtwOxyzIiQJTQySimd51wX8zTDMi+Dim
U6HbHMK4S0bOmHYy8bF3xDj+tGhfvk34FoZHjxUrGwyxMdg7S9H8E9QFTuIe9fXru0dOM446/2Sb
+RZDD8kXhGWSXj6mj2t2rtjvJkqpz0E+D5w+1TtX+6DGD4H8nMF8TzwJX3tcDqf/xAr+PvAtOTOZ
zlRuah+aNzjwzjeNblCB6dM2tn1IHTSg0HeTTB41QX0OyqkYvnwCVUKaEneDZuBDgDAcaZ3IQ/Ge
0nJInmrYcvCpkMaOtX1apzkZEy6X3C/5KVfurnEi8Cr5WONZZTUhQ532+R3IEvPBP6XOfR8Ws2Oi
ePDTZSKkFNJgH77hJEgsb8URcIJLNW7mztX+VpFvqwZS7EtCNCsAYaxEVskAPzyCI5uBrfIwCEhq
ksL7xU+IU+et4+fp/P1RN8y1MqIM9RY09tHePYbrcdw6+pAzO4GdvdFPVlBsFNyMF+Qbzf9bomt7
L4RMGGWuXLViPcyYva10iahuSYrM+8mf5EAW6U/4z8XAXS/w9/9EjseNPErJilGdnIM5Ftp/L7Br
OPjfP2xGxtOSzOJtw6ksvARt2zPmDmC9t0M4dPfSqN4q3nTpkr72SMCD87z8JhHJvTBhzj/CSZcR
Fn3b0PMPtPI/k5+f0ls8Kwb1F9CwMJqo1z2xUB565tsUGxx/qeUGyQYUFl5yJS+8476EMri+BBtj
R0WppkYleBv18nxCRRmCs5YRsB1SuKMY5BvfQqNhwQX52Dh/F9c7uSbJCzhkEfXTTJV5GN+PhGvE
bDaeM2NmBp00r5pkfghiZGho9QIZVJm50hQWsOixYbyg5rfxdfDDkyuty3ruoenf2dJrGtrAN7Pl
ijdXDlKXtIX54XrbByc2oNi7lQqcK6ogUMEmae4mzYDnDxUSOVhYeWiO4cL6EI2hD7r9bG1i7pYR
1t7srvC4BdJdFh0FMwFSdCq5kaoD099vhrviPQS27kflnNlFs7pNuiNpSEb3Cjv5CUa5JKbMOpIs
tBVNnbTmerYcKMkVhx7GBOpj39XtIDI2xQusTyJdDpL+ZsXCW2FGssSwCWQY0TZpmHHoDzOCW4GL
qq1S6F96T79VW+HcojiDwI+4xnc33cG9V8ySDw/UfkLrzS3nuzHJB1w4+vz/ok5oHK+CS1NIRMd+
JTLQoVmOXNeh0sUkkCOq80hcFxL4WMoi4ysVH2ChAz53YYlJgbluc0B2vfgVzqAV7dsN0QQPU+sK
uo1pZe95Ym3ELr/wuL3cTbmcyPxrUeXzcvcsAzB0kmNsf+GP5fK0lo+tI57LBAmN17CeosQhHpfs
go2OlxrESIYzRGjmIjYzoeZaVY2+Z5ufdVasR4kcGPM5iLABOXVGZzPuYjMXOTXvdPgGMzB8UFiJ
Rr8HDQtDvW6svUVlvyEiAK1u47b+BJmaKWUStV0tnhAZxL4NNwxFYorZcFEaiPdDcRrXbZA8rtPD
RcFFRf8xJy36rX1u1rplbiOjd0XC/XlLP8PX1QAEIbUonh3O3cE6AmOsAi3df57gSw0EG2xiAlVC
w52+QhOWmS6pTPXosDQAPJ8FH7YTbOCejf685d9qVKos+36hcY9wqSAku5BSVcnckhpZRCMDhoa8
rPa4xgRcriBgMliAn60RR3MlIVee5TnrxHYYpJnSM5qCV9f1p/F1L6eOYBC2MNbbL17qQUJm70lq
moGqpO/ixD5L7nZtK16xW0PqZ38KV2bqVLKhSexA7KLHQkpd3IcA2NT9rswbpsv4Eslw9loS/pq6
Y2veyxV2la8GMgUI3h1qrq+ydaYFKjWVKnf9Tsz6hPqbRMnuyHF+7JIqo3FP1zubeOgg6GArvG1p
GbA6HsfgCGYosHxwSL3OUpRZJLlhMr/G4n6mXXuP9mh0tup0ryrxFLXexdB2v49UnARfNK/jnjDA
DliqZ4O1aDvm5bzathqZb/1Q67NSTTuIoOC6zpsC5vIHjT/ohdCPS+g5+IxFl1aw6E2BcpitHo/V
hYDcEul9CGpKSDAy8zPbVlymcej7YMzCDHv4VozYQAWFGKSt5TrLf+fRXAVqesUh1U/3ZaiaY5aR
KBxx8KXFUSYqie4/N4RLClxQkPqfoWl5Oq+OW+qUf6PCs4qMFvPk/OquagC6x9s/sVtXQbHNbbbs
wE06XLxUa9XdQeKstM5lsPbwQTSmoCczQkC3B3i5mzH2b6QaS2EqJbhIPDBNTRmIH7Z0wkvlvdpx
jlXei+qIVu+idBAMetJF8XUZDdNAuwhN7KK0oDXLX3cL7byDq3ktgYLp7J37/ReTxArJhzKiytMV
VxWPyaGhUTHym2c7FI0KMeK4CFn4bbdIzqu8axtl1m00bGhohhR/oITo9Krr5YFr+YVUhHyNl3iQ
DGvJ+4Kcn1AfG6zryY/M32RP7YVgIMXvVpyVQicK0MWJ+CBWxkg3oGYJZaXSPwnqKUJvWvkCybkr
dfh/gnf690n4abxzbnIabtuwWlXFEYVScZDNuR3/fyktij7FWlmf8bqAB4i7glMigHA9GeQrRT84
32Mnu2HtytwbwcmMjWeYtuF/6VTBpJyQgVA1mYTatim4iQjyJemRP+myhjAGQbEuuvoGKM5zgOVU
IqlhOJBt8sCX0vlC9mcS4u0VwJ73iJ5zyR84zj68rMXT6dW3sL27cM08HNoxUVdBCQ26XV2a1BkU
3vu/2+hU09jERLQILJyKOhtHGLaIYxisuq4yk/nUAjI9SsV1hbNcSMZsmfXbfoLN5bEFRR9Y+wLl
0MLrwbqv7YLmh/Wod6JnWTTKrnyjsxAz8WE2iyUUyiMkotlqlpOLUOY0VWAs8YkeWLiBtCJOe6/g
lS4RT5dpofHji9KSkMr8a7EYMaE4cS1K+5y4y2WCN4t/wA+Fu6hZeEJ6/V1wTZL6UKDguHVXVp2G
NJ9VDCFwdWTe0zmZhqi9Hz1+Zc4OLORt1UpfgbfUEI3Z0vyYxzbWG7Nm/JqPUtXGvOLMo1sq7X0u
QTILhBjJUb8t67PtEPCW5I0CuAe0o0UuSJr3ra/sjkay+hyleNv+uhNyYZfOzQtdI5an39OLENuC
z/o41OVh6a51Wp67iauTurxoCgQwXRvnB98qxDhYkrkW8VQDxiecHZ2njES2x3/JWKfBWM7lVAzK
cYNurO+oUn8T28jqoyBFFQG5YZC4Ra62asHS4hx+Wy0feOX83KX9WPwuRXWV5dYmrg/PBQcdb6Zg
BXZXeM44rGnCDEavc53doN02UdQaCPcJTprLKLwoO8FMHIpu6PuaarF7bJhJ/ZWsTMzbQszMd1UN
UNtRDETXi8WskbwzkIke1hQSwi31ITLSP9oT2C9jqglP4oxfVPcPnia4hrwDupu8LSMD9hJA7u5M
9y8BG9TgsxsPvQakNeDZ68p5rMBBQtUHwXceHyecOQEkhlQQfvnwnE0+8Es/mo0p3yhZOmKe3NmN
DCyGVBGOTSg1/US6GkZszNjEjx9La+zNZJYJ6KxUa1aICvyQtfowfFVWGUKG5wcdfd2fPbu9qbwk
W7JLnIuw9wbdcJ4yn2iJJlJXIRv9SXgsFPVr7ChO3fx2P8oHZ2E1yQph/rQUDxtYG/uQGL3v/Cbt
2sR2wueavqJUDzS32Ivx+958OrTEQ1xP+HaxPmLZ6rs6FeV4AGSaGfiMnwwcfzH/aWeimmD0J7I9
WLEJAr10L9UF40SZBwSScEvmBStqGvkOZsHiUV93AjTSbgSCX6quvQKWQQpEJZzghmp+FZRRhOeP
/yme6Vfe0kcq+6KvtmQBNU5H0TO3p33NzMoU/xX2A6A0SJYwndEi9nG47dQZHoSOfzOqUuzSEOLD
gFBik9Suzk4HX1W7hUXL9Tcg6THHxPEyPVib9wUyhnHeWMJAW1LuI5D8J/1SfENjaP1CkdqW3Gg0
04n2++GmNCF59BPInemfDp8zF+4UJ5zzTEeXMgTX6LZyDFGVPTr2D1OOhVaMIdTMP4kL9b+6eO/S
Ad85Iy/tXyjcRStJFIUhLnkFgEUkLU+3FGJh2QCNBXiC6aeKnKHyWOvMwLhlkCtIQ+wDmrzjOn7q
2wHGIzQ7NEFYN1MG9Sibmc1NHi3Tou2gWVcnTNjn4nKX5cuavRY54hiy6m6JpzhOjNtLvZOBWFX/
Jsi03SOOqJuwKvOHlw+jIVZDhPSk+MIk5Ma+PCRkentDEbT1yNVoRCp9dC6dUVHIEx5jUxE3HLId
QqE2YIEG09rP41GgoAq1oRHkrsLXDRvqW8LGsD+Li5mp1iZQ+pd5YVicgo+I1iH2KlWdcI4DKNMF
UW4sfWgf14RyRrPzH6hygCqhpX9exIshtCdBduyfvk04JyjzTCg1zneiendaLcTpcX89VV2XHDUj
fF5g2Qlv8eTTGbzBGQuj5iK+ne+9tv4h0s8/DG/37+rk1a267MwEZ0kiVEZTH9JWL0QhiDxV3GZ0
RXoYhKLp1W5YJWQj0Dqjm678A5UUEgmBgoFLPRE2OIUzhXRCaZ3UyPRcD1gaLLl0Uzkyvsyc2ea4
Ha0nddBffQuJQSKosyQ7L++pKp1Xu7I805o6eugzIX2LFC/UVHi6b7U9jSQl6jTvNiiMlTacBd3b
VXS57Grej0gQ5ss/73P49BIuvDr9rnDmIK7kkUdE1ZYeDSLsW9Bl23lsr26hkWW+o/gO7jZuh2LU
OPDSqnzXuodF33hh1nXhPlJXcpEpBN6QTXhSlogb6NpGwd0lp6vv1qli0ouVGB82jNtiUOI4PxbG
TA9VPArDyOI3PvtnNnYYylbvN3ixkO2t5fmJYXKEfS9YUyMJbjvqQMSKn4ASdCjZyHPtSstJgqM0
cdsBcyuXHVe0iyDZ9Pnbf15+ZENfMQwipeJfwQVzAb1/1nw2ryr5EacQ0GwqO+2598z+pBJprtze
/kuBv5XARoXnvVgNVOUgFxqJrdDldJwO03lp/7u5LY25KMpc6RZ0NcTca/LmT6Di0zyLBTEtYY1S
X9QP7zTdsnH0PTugr0Jk/TXLKcRMSegjrLc+FfelDUQ4qg3tt/Syuy7Q7BGfHAhqnXJi2pihX3G7
CYvDyGv60xM5nEXhwn14d4FO4fGABC2DmfGqYq4KHBPgzCMYcn91goMONLAyU6UKwY1FGGNmoM6x
ppUzYb5830TidF1fW7njeaWWI4d8HNTpxQD7sGfS3kpQSrGZMQn62q0C+kAapz7r3DzvZ8SG8YEG
rUJQswarU+gk1I9sVhMpfpnhclkKCpP8O4pXsbLJbImqyKFPLyiteLhaVwAO/ltUXZYl3cJXzzqg
rkS66/jY1m921KcXjV49VROXsX8l5rm6cC1U4OuurXQHRoVW1HdDmNwFHxM9NXbzbFSGogXb4me8
0arJrP3PXpB5AR9kDIXbqAKgAOqhwPUpPjE45IwENv7ilXew1S1xwzLqPD1+lrl8NXrVtGT1vd+A
Vz4NtocW5vjLtK2TomHg+GDu/cvGUQnCIa50bFUcoEy7/TUnTrQIXwJ+O5BHW6pV7EEhBtLx1jHw
WL4Ab8h6uuUtOW1UZpu+54oeImi7NOMxztwvYlggHx2ecENZT2od994rtDxEHTDVRC6nFHXKD00n
EeVOYgHRjWsPoiHEK8p4HAbNChhDRr0JFPso816d0YejpIWJabnoZEv8XtCfP3FYn38CNzsid96J
OZHqRRUMZ1zgKMKPK6RmDtw9/ard0sGU8Ggb9HA6RRp3GGNTPsqlUnjuATO7odHffNL+WGm7nfmx
d6A1k/10e48xgEq+sQLZG9EFLghdxxYbWpP5YkfwRX6S0lMg0XlHpHd+uEAH0Ow3Fv9Yqt7jnI93
snuvFegoLg+oZPlqgM41dc5nKxPxJkq/3lqmgA0SIji4lZgtSqyfwWgGJsZJQ6OUGN/SE08TsLOw
Kw6tVnguMOJeYjlEMqQxXt41Y58H7vlXikwklQMgSe7+rC2PJ/ttktVnt/PYGHWIHX5172kfxZE5
Xu2OEQHXq1COOehIcckXFAI0S+ZETOB8ENJvTiQFGUCa56oR7yrvwVyw8+ZW65d9iXb0MkB+mBEY
tOCBOrVBbmICv22JC1lQtLlGzaCZXh6ui4qLlj5gdMDz35pbYnhm/BvM5r6EL1Nie1k30yg2oO8c
6/wnFIMK0i8xelVeGSEqsDBeaC5hct5cqTJzj1YqSwZ1saiMR+ZakYp1hwfiF0bmoAqiKpxyOA8T
93XpQgDfukEkilDV9YYZQ/50kZ+kxPrtBSFCk2C5PhBUSMWskZ+l14nnvKEC4xe2CwrfLVQBDMm/
+AWroweHlceGj2sqrJiCIy96i/GmX4iSuSnESBir16lsyqz/IUX/8v1fba28W+qnhFzv8wxPWL6q
3HjSSltyj2EkKuZYiFQ/BbzxhndzY9KH5ZfmlQQaAfhAlswM0y9eNkWgiJFbS2kXRJEwj5iOuupW
yMhPOY86HT7GGIj6Tc2c0TC3ewA6ruo++C3SxyWYHWM0lVR0VO+e8/AHLZDqJ/VKmGY6VLGBSj9z
qBzNzq9nCnwc/CZHOKVA56SlKGvMyU1hm4ALVieF4sOnajUTgDjdkJzyXO1JEPgqn26iPXnoDI3y
VDatGT5dcnHHb37XBGupo7yUEz6T1oIsBGvRuHaEUUMAja+asOk/YYPUaV4ESJZuWUex+mmx5ndk
O0731nKFyE9hHIP24LBhGxFgNwPLICmbvbamd7aZXekZOjbaXTB7QK8t/7M1GGuLeW+vA/msOfgb
vnGbeQXuiU1ndigGnMx6GdbOMftJSuiV7kDGo2oALcjKYfDAaxfgYfr9YgxylVGeYDqZJ9tQrowu
YCwRwQA3ygtvaEVIpnE5n8Ed9ydedtdKuEbT1cxdanGwHzEYQ/Z5fPmMSp1DMp3dxzFzPP6p3+rg
bNIrnSRsz+IlnXpcT+3GiWQSYzrniiSqpqyayjo+LxbI2uYMIo7hqWWLwEl80SKsX+hfZs1w1vof
XeS3bTXS73aaThN3ZgKmviooJ8cUeQPRy27aCyfaVnjHl1ockyXDBOJXg78YJTj1UudH/5LSeN8p
kTA8JtCcpUM3u6zVHDVDfaGK4MJ0BTN2SAMSpQJUSPIfEnH/x0aVI7tNM+04qXLq8f/sLWL/2kk2
5JXDoQ7bCXg7uFkru5XvpBeuyOZMa2ekx8ac6kxPk8/ysF8Me/Fjp9dUQsyesYtqawHuE5xPz/GM
l5ao8G5mPt7bQoB4fmJfuePGSYZsOl7oLRHDwFkAwQoLLNy6NSLz5A3oS00gksZ9HCOEV4AXuMEz
YSDX4ayigeT7x30gy8pxfJa6ZdCHdza65oOZT3B2qWww/9yMfvXD3fmqZQmo/UhtznZly6eGKedq
kRCCyZ5G61dn59rRarK1lM/As+73LyNBZ03fd5mJQI03Wf3Ogy67NSv+O99nBIa1+blwPcZtijc5
Ibl01Y/wy8iYfBd4A8xLhBfsX4ZowwZZ9TFWo0B7u3U5s+vdiQh6jD5yBq4wG9Ix2yJxDGVPqWcZ
PaKlJsEs8/FzPYwujJEfQzEhm0XJrzrFp26SdeOobp6EyX73z+my5lVM7OPuScOhFoU1+ZVCcBcL
gyC4XFtTP2VyCLB0h1FlI9j405Y1v3Y3XjFqcWcE4oP0GuwlFt7iZrT04YzK4cpIN2r0uPKNAKA2
6JJ4dOw6KbfT5/i66PTdVrwCPKuxM7nNHfOp2MDOevFT5uX3M/QUF8k4uDNzR4VJJ3wNk0QAv3ao
2B2IIdpG9KPNgrCmRUyYOs8ePwnULQo4t5TTa8SeqclSbtkJY9WYr35z0VEauMXa3cTtP8rGAPbL
aGOVFwV2KlJRmfDbnh+zdehx7Z1vStvaAJSPWKMBRaibYkuVEC8KPyniUJ8r7/zvzAvLBFYDGT20
i+wUJomCRpiBZon9FSv/ExColmf1TxPlxvrLa/YzATYOCbnHnuKe21Ep7aqw2WKpCTReK6LTN1SK
8WLwDl/hiWaSygDx+irPsDqbVZ0Z9RiI7WEVfxqHYl3IXk16r6Wuu49+4tNdwMNamcI1aftntOLt
Ud0n2Mneom8bN9rT83mde7+RTy/qcuzqf5eeRBhFvPGk5JndRG+4pCxq6ZXnGNWOGNQQYNUfGDSh
Yq/UBx78aOKJ6p+UVsm01HP+jtAB+5vBESI6KJy9vX7K1OeMSobJ7aWE+T5wnEyU/QqXohgOpnom
Rsr/WegiAAD6idJwVWao/TqtUDYpmOzrZlxxGVgKawKXI5NH0S/wfl1OcfNikC+9Q277OTJWWtSc
IqTpnoShehPbPk55uMU0ZL77b/uRWMnMgIXTCf5gtSTUzSw5D7ISl1XS0YoBbLejfnQy9hA8m3ra
ZeS+l6M3PGSSGtBs8hLpmMPWNpeCHA5BwFxGwmEUy2QYJymq3bIdDZcxwdDQ3aTNYt2Ib+/eQNsv
XK19Aw54hmG6z53jBjiDddXWeN1foMIaFFve/sVJAJNTNF5AtCU4IvD360Vq9+fPfdlt1SSgrlEU
ZYuIOu4D8pFErrQ7O+lE/2oORaiHpUYcXUEETjfKW41eLoa8hvgH0dzWxwiVuhigD2CCBWCOLgya
/r9xYZsdaut1xvciXeOx6CNywV8S5JyLIWs57K0opon1TFMG3ZGTt3r2B0tYCSARS6c+DAvknhfK
1vihvU1M5uhaZGR5EuT40OimvePDpMA1rx1M2iaLNlUuM/+wnK/cMr+fRBPB2MbeQiIcEhOKSATt
LrlfAmknWkTvHv9VGQ5y6Br3pfkOM40VKsKt7zsYyyi+HEFgdSIgTi3DxwcQUzvNOy3ljyxszXGO
/gT3VWKo3Zu5V2RN4XWvdgczgN+sLLuihIymnEbcqc99nryINKfzRaumaortq7iOO8Lfph0wu22t
w3xopdkb+wCON3tmaD+7aattD99dKHEw5UyVDbzrjHClPgTMpifHAZjdIErgPOHZ9vHUGVAkriT+
AnGHk0fCGgrdaB+S5DfNTH7b/NVEoa6XwYot5p4jwbeVlZ15jLWFuIaPo7IaX4OhP+GlKH5WaCMA
D36848pjj6bDiG86KH/OObcIQHa6/BhiPLxYtFbFskjxGpkm/pqVgZfLmjg93eA5J8cbIQaDVM7q
nebZsOSx+0afNZMLnc5PaK1tP6zf5xyqcndKBz3p+qkChTH+hpiOyvGOewk/rt0J5SqPG6iV/4+t
U3DOjg5qoTAo5L294l63uaxZanHkMxaINMTCMwpIAKiWfFVSwCeS9FURGC1WWJgbKiNXf05g0z7y
YrkiEmrafcYbP2qIVUahdqHpIVDCyeD5rxBIqoZw2JuRqzRumbtUkvR7phYqoOzY5w8yqmjsMsZh
/1papCkukY2tOndINJuwyP7ocyjPJyuvFVk2iiFPAM5bUlWnko2TZB7Bawd2b4GErA66rnglutwf
2KgQxC9iabpkhQTBb0MjfQKN4crbQf4zVOTJjp8ZmWIhLyca8kD7yj7whWoEVllpz3nurmkYlqNA
ZPYAE06cVrdxa2SefYbYz+xGZ1M4lBUApD7sfmA+8krzKnEo6SP0jHeneWwhQqizCIcIuVWP6wnS
r4UyhR1k9O34N9zwbsJLtGxdIl1XrMO4E8Bnby5/PehutK9nVUqGSnwVbmYys7BvEQqaRSkV7M3j
MtYzuDNcYMYE2/iIUR2h0Y7I1UUBgsTREKfCj7ZGoSgi3D2h1DZD0WTBq4Uo17oTOSeAX9JKa/5c
WhH8TnNLzPzsnSXGoxyJRRuhesygqo/8Aqlcs2KZbY92rufhnn4FCOQx/UHo4jwptLIW6M8ffAM1
qbtve+qUuWxGfMbG2bK7Qv3dKF3rHXD1PsCla3afPpBZ/kx6MEIRmV3TebNX8Lu3/Hvk6XYnsF0K
JMAGp76O78ceyNCcVTDXTLsJt8k+Ng3bb/iiBXpXybt3U0/4rxihqpVaM94JwMzwI0kfVpqWsn3m
JVmCuxRy+BR/rDSZ3IuR6i8adSlOimCArXEb0SVaa96cK6MQKpClgomxnm3jSkBNiG98Rx6BD2mw
7zJBYO/E3xE1VWk43G1/D0AvgNbBKBnbMVeIBDdpABXjXVm3rh69pIL5aw5zAhtb/IeAnD0ibgmm
7+cPoDUufh58lU/V1M4HzFM7V4oxY0Vn6xa3J0HZvbz6300CROhs0AdZL0kQ3dSwf14LBmFnYFFf
biEAs2B4c54wV5HuxRkiU8eLwI5G7b73DpweP+bEcSKuZLyqbBMgpkKvHahp2wMLyzvkBFmakyO0
DKo+t6lnQyURcuTxdDS4/PPWXlflvI66mw7nHehZSz259QzljiO16dSRsJZwSL0ZeHrg3sES16Yd
RpC2pH1s93NxMP14JJs8AclTbLJ+fGk1fAW2ayVYXTX6/wmySSfbsJmeCpt7AMP6gU2D1yvUXfFG
/vkMk2oUAFygimMNLvxoFmGORIs/y8yGXGKHXD3rt0JK95asudUdqpEEPZ2Ra7g/3jserfFnF8EW
KqTBPf28+snp+nDC5/zXae2PQ6xqQr6wSHoXLx6QVbHhoPolulVn6xZA9hnooirws83fwoIFa6ar
KsDyNsh8jBKn8RqIVB5+WQpQgFVVCVieUbNJIG8BJ9BGO8hRcdd7QRzuMdxH5tQntRUSxJRwv3gi
QetnjUv78OA6zYH5EN9rpTqNwGiDcSia6Kc1l5PmnQ8jEIttHAl61p2P9JuVSGw5oUFnKi2p0vg7
oNnA1QDEc5ZFbNLYMWcEaX3aOwv4B4eWavLTxpradk3qQJtlxUHAhtx919aWpDsk6HuUj6tmQ++/
i6OdaU3BbNbwUhP9OCNDTqkCTQyBO7CAX9ziqtnwrvAHCFaw6Gx7JuGz9V4j4YuPvuH0elz8P7WK
HVL1NAUMGqDFpwLwN1z3iBwZawGm0oKx5hY6qvezkZ8WMvoUFnixDR7iDeZFu5dO6BkWCOf9IHjJ
QUzB3e0kNRrIXrdZyn5HeRbQgsPX6htC9YxomSeAh7GxbFJizUBg41QCAO/fSc8FUmMp0M9LTFBq
d5qfa+rZYwYd+6Ns0EsGD5AMf3gG1uFqIo5jBil5h57FBZlQMMRh475SNsu7VVSu8Xj6cXISnRX9
uhKoo6HN4yCFEceL8Omqa7nng04D/MlPlCF2qH+z+hpBoZwjc5W6kadoB78of3haM33S4Kw6lBPf
y0xFjhEVZEZL6xKw8L4nWO3e9tVG6rD4EOfxARaVeLvK7bH3BXAt/klrGmuv5qfRobUyjgbJWvO4
0wG9TdB6sXgPeaIUKP33GQMaU7sb0mYLq+DeWUJwRdpQtrebMCaINgZ+hGK4FFK59/fmY3LTxWE8
QGeNHIUAGz/EmTf8TNsp5TM9ce96dxqApdLWkqrWLwYJeS/od3HVPa41I28dLjXs8aatnC/NWxMC
91GXRYeDJMIU4JXFTBBPOMHTxvXAOc8v13JQKOg7aHvwSLNrdytfv8p1NSHSf760qBpoBSbZlleb
dZDQMUAKwJxJkMu7plVoXRZt4LS21KgdPqKCir4PxWUfxz9qKPay7kznQsM9KLKHcT3SP0WlXAFc
9uUDXP+qh5u0SPKfvJ+WD2M0NVoJskljUHLTfxIndrR8Qbp0M10ubQ3Qoj+xtDhv/gp7fsOSmFUu
ag+FENq6oHOb8wN7I54e5GUa574zz9FC3Y4TkDPoXdWj+Vfq2TkY/VBhv81UN9vc5gGsjbG8dtKa
o8h7ULSpOe72nk4hI0B2ZUMTQwDar8ogXT84cCNq9CUGWtQuTHPt71dx3PlMDVz2WCHWAoNZS34E
wXP5RkIbMvD4V5RqI9HyJMy4+ThANUHUc9cV+2l4Q9jV56fAAYPxgdf5iU2Vp5gwwVaxXhpmGt/C
DH983Su691saHd5+Sao8VkDlMrrZj+Z/+dVT+EYH480KNUGmeQfNkw1dnoKfTl0NuTMPwzQiH/GV
s2kjiJNPLNoEvhndiOAfTDv55gIvCnd9wYaWa6EZoan/oHcnWpk59ZG0luaSakheN9N2TotBnVwq
R6lxVfgRhJqzUbm2I0iX48TxvXkhd2U9lIQmtGwk/hseudSAQVIDZO6fcsw1di/p/h9g4n+95ySF
QyiMgT8gQaFAfpI9Abnu06iW3ZfOHVbV26IRqkDo7iyrBH1FVE11pJym3jDtbAQ2xtiaw7nXDRL8
fN+v1WFlSeWBhScohNXIOdU8PHle7rAHW93LIiATkxepKdmreqYFz7uSC8dylaSgl9C+RcFGvl42
QIpN9s4M+hHmunaAZGjqGq018Q++AzDmUyFO0zSGFZovhkPDq2B56oqfDNC7bCQFr6NndLZs69am
CR0ybUv6AN2Sfvn+jfuu/10nD7KEKqq38nSkmWVgcK0KCT/w9i7v/B9n5kLCZekS57Ym9Zua+59c
ERyTJF7Wdq9NhdouLFJkmHedYq0lC/bGpf/pUkh15IB6Xjf1Z8DT+4a6880HNZp+cJ41t3kT84Y/
hHkhTP7Vno7/bMNq3HoolMBqbB0NbL/ajcuHi4OMMnZ/MTKhYZxB9Hme7E7JWncYoaTHFkM78j0j
TSs0trOfyEAyVDSw5E+5vnkvDMXNf6eFzr5LmI6f4GpSI133OqJvdIyNZ9n0lBUhXoWFzGBAzu2G
iAiAZRhXY5MjFbOXl6b1ybtOx05isbuFvAPJLz+qyPV88e8n261lMzPTP2mLUnlhwm9Tq1fQmzoG
F4ZuibB3udz2Mnm9Qn/EG42LBUYQ/TO6KM1+Lnht4xfeLBpOF/ovK81blwfgG5voLdU7eayfsyWX
r5kOBJ+JemB1nX+JW4nCZxD51YDcMzegPkAY7U0acsO4r9ZTHaFPRTImElgeNtMkUPXhllGNrWJS
eMY1OZQjg023aZjaQGFWdcWnQaGXMk6YpRFsWam1kThG5eUXlgk5C1MhM+pTxyMLfQNCWeVLn+FH
yxCyOmEIRdTK/OZnhulQ8Ttd5+9EW7Z5b0bkJclRuUXJu6EKsKnRzsSYzZvZ3fmKBoNwsvjMn1Vy
YFxL6QkqBPBKzzmBmvf2wI9tng6XTxJQLflkRhtGO4mIWyFEbyxp7FgruTA/0zgYO5gn6wefaea3
GZQDG55K4IXZTUfz6RasmTlGJAKZQ07iOq+vbtk2N63PisyNsOIwGg5ya+OOjAVxW1RC4+GaQ/ks
YmSLVt/GLZ2yR4G3XeDoxbi3bvgpdHcw6vhWBv1xpceewhsMbfhMnD7sV0ffEi3JEL88zyiFJOCS
Z4lVMBDDVqm91uJ8VmXM+7VzfPMSYVC9E0Wb5jbdM7IQoGB0lai83cF84XY97kFhYnekE1WNnM0S
LT1EK4ejefdyQpgf+ZuOYkQNMbrOWSEWIR1pOdrKXMCqI60PCFZfnIseQ6FEpSZyfG8HKNSbve9q
PtxH3Mwlu1Pevr9rAorjIPQ5NY7rx0c/WXmDS/BO3KBw0yDpsSleG+TlGNG6NBVMoDMTpG2d26S4
F5SnIXnCTbgfZShWwLLMNuUu/baNXA7YUZTGOJGBhd0YnlW8vZuq6qzWmXdNPMbLNgloNxHimuu5
JypuJ05QW7O13NMLpWvv+AY/AgHDyx7ync1id/h3TR4etM7urXjpG71W3FM9BJ8cs50f8KD5xlK+
1loGwsgGpdGPPuVidvpOFQpu48Dxvnd2HkGQsHQUc2OYhofzOnYXllloYRs/xR/eMvjWnQagc41m
emg1qVEUZUSS6Wl6y2Xn+6zZi1BaFFw/eqm9Zg0eD1Q6KAq7bvZ48YAazJMeYYKJYnPhhDaepDyA
71QWynMgH5vYc1FD8UbhLHzz/rrB+6HFdsygFeTA8Bg4XF6e98eR1M/wVZ3u+Ep2/Wq+90/9Bqfl
1Feq9KbCM7eqtDo0UajQ69cX2G3mpygi0KkrCb5KIGrJiqA5p3WIwsLopaud+LEJ9n6J5/dm/Rbw
QPgffKISR1ClpzFtVkhZ2zLvw1ALbWIVjQ3+rCt/GxwUCttcBccxrvT8yusaM5p7zRAzPr/pupLL
BIcqT+KYPqBNSERCGGcNeTHzu/l50d+l3A7UZMz0WkVyCV5Ieoxmjm9nmV1IcbackB/QCrZDcgrq
0HWQEnG8RkWiv9AuGr6YDxsZj+UrGKy/phBFCUAb8UcK3wwKLJac30jvMKIuW0MDdsGjinC2uv9M
n2jkBTioKmjBpH+XnZhSlX0ejxR3ZQqy/E2vJGnqfOx/5Vh1cr82ANHEHnhaEMrF0EgjD2OMb6rz
/yItlI39tki18EbllvNDe0ndRH6iovwyAHxQQwHealUh7P7Gy6M7l3hpZAaylsAzzYkCoxBypprn
NWbfNkKv3KyxJy5eqOqlY+TtSmw741C7KRrzmZEWtQNFGJurXqafyi/aB+6hXH5u3eAsb+zQP5ow
9UYD/zUMDcXa5PL4mB0QBXmWbSwsBCJ/4tde+NAojaBYtyD5OJEQ3ZEZDMOPIv5sth7BtMjEYEm+
9Kkg1lT/aLgbHh4YF2HDvn7ApwqLfVQN0M2FQSAXd49Vk98X44F+4Gd/x29GhIUhwjWRc9Ua/leY
zMK7Mg0VvCOoZu9JzY5MzHDYoDVbCRgLEjqJyg9hAx4eQubtyDNHOqBzk04sgjHtMKlwYyajLMej
9NI/qmmm/XBnUBmYr36aRCsa/sxxpaZBScI4Q++TXuIjWu0ruueRGyaBsiifc0LPikL4hi5nFC/a
hgI7IPqxFeIFvOHZreQoObZitKsZfbHP+vhgl5wBb1Xv9zpICNzacwFX7AKRli9lEtUMUEdvNURB
9C3QbgCglFda/TlvbX96blTrZrljIS3n2UOJ7iuLpQKrTSELTe1PCbDgjUL+Bkm+Lw2pZlTDL86b
efNSoOXuqk6B+oh0C8le6WTURCJkWa+DBw/SBCH+8GuvXKh1Jjdh0DMoed/+MhnYe6si1DjOH9oY
3CKjsFdR2HOngk/rV+HiXl9CLIl+uz1ZokaQ0Hp7P65SeH5/YneQYV4tO0FwEA/llCRUXLacCVEQ
RR3PXvUAafV6ndSH3f9ea/kMyZfm5dL3rt9AM7pM+bbCYjehh+zYQysiqAgqdmYn54RwyTZ4R8YJ
xaBncc6v6MHr82jya9oLqbWSJBuVuiW/NN9or6d8erdwwXXURJVSiGx6qr29jwlHYvXIkVoIixlR
46vajF74GRuFjMdAu2KBSuZyEf3HtRJVAjaor58DcOwtwS5Li3zyKageLJASvrglko00+vnHoccc
Zm5pEZilLhmW3D4aCL8AXTdt204m2G2W+IsxtLE750HYHZJmrR98f+aih9KsksVuT5NGZpvtXbEV
b5THe83ZaTSTwoqKBVE30yTjQ3mm0x6tJVIkTckpQVjLPUMDO4/aHM0xbkUjWB91441nVVUscRbs
pFOS7clir3eB2LQRBzLL/9PaIwD1QgGZNwHcKJE8n7wOCta96ntTMQ4mbpyyGmuEBiFte3ylH1LB
yOE0JSQbM+uY4haYoJbsKzzLSMqzGrsWTSlyn4DqatXDG4dfDK/A7qTNT+vMSJJMP0JjCcuMxPZu
K4WHZXrn8/EyyYizXIrWmFWuzOT8E1adW3ntXDurW8GA7kgmkSGS32OvMc6P5d6DFZWhDJNIAWne
jIz+gOGuRkeskF5BFULjtYTgP1i1P4RH4mTyHt3C2WfZt5eS6DVcF4RqDRIAJ2B3jCsqXLjNLmeN
cht9HmBq4R0vJmBZyZURf4R/SNUKNDBz5BRYCgb39pMuaLjx+VfT1/104WS3jJhWoTXaeP11N2ia
/qn2mTwHtvgfZyukzMK2SbyhXF/tWzt0qMTNoUdFAs8Hp3UdmUEyFDF8yJlsKffNALPmijg8ZdG6
OQ4TPJpgJtmQa4/8LcoIKhL70dO74YUzgwu28SRxS/bjJWex6oldLFWJS3RXdGY6kXeoKUX5XbWG
XRpBiMy/rJ1RBkxz1HSc0jbGlaSUwc98N2CF7EQvWgKf4LDA74Su73IraEmlUVC8Sn7o5a8+9TI3
YLFg9MDX6Qm/+NxevhyF2WQUhbLGxP4vD5t5N7cQH7thhd87ToK0yk5GZUfPgW5WRt8ZqN0lHwrP
uhN+goQtG49pSGDMAnCplBSDyyr1hsa0weR5yEQfBN98uteDQiTT0YhfTKV82wRD7go+FCxMPURQ
8W43qQvRHFDrHsFnbkCXVNfMTBMNt+84qEKzC1qMfmNMRMaH+JCxuiV3B3ljNk98sRc4LON+g/OG
Ipp2e5TqRfN3PtxyTAA1ABBsC08lR3rLginijYHThCGQBFzXzP3sX3KTgQoxCSWOQBFxKUHcFZwG
XXKNbxNXFL9PqL/e3XXaMhXXg9R88X9Y+id3xuxCNdKnKEQyNaX6mSc5kBaaUdlrzRB0ULewkhX0
7DCzPDBy+UctfbLRuDOk+kWIDwIx3VNKnVNEjgGq42oEHsR+uyKEOFOiv/xn9jYidv2yT9GkBTAr
yaCJhOiFe+u10kTXydUNExDgZQp8+RJnc/OhOKxgdUeg4ojSePWQo68MPtdWfSCFUXEsdWXNnQca
B9IFUNuNyOqngsEQ8gnh36o8RwjtjJO37QHR2AwvUIrL8I2B3uqSsHQkBPNriwf6zcC6hxOmo8qp
m8AwT5UvmuDdkIkelKWUbBMJaTxiB2G1+GqA3qdUCxHlZvlji2sCOQjT3OiyizO1lpT5hyAWh3NY
nFmw0gUaB/X8QCdcSrCh2mhm4KxQmQqeOaY1uOObHCcPmQGi6xZ04mpUx6B8C2gX1pVI+ca3sBLb
deLguitZNff+p5HX71tzqG4TzZxoUEWkk9a6aTf8RJxJLFUMtoHf8/igXotp0cH0lzlVUTXinaUv
7n0R/tf5noEHb5s12H9NmKT0sLHqk147CjifamluHp2nB0LDe1SqV0bCJKlBXuiLEHjs1I5iLqas
apALNclEFqW11gJ3jztmrADPCOEr2Am8XRDvqtOys4vlQZb7YYQdShJQv1/C1gGbh7d5gGe0Cs1d
iL72LBLMkLjjHRQI2ABHPokiRH4WbOmt9DNwQ4CD9SyW10g1xSvwWtChLe1xax0U2GSUSXD7eS0c
RrXHCgLwiFBBQjGqY+elYg2JLQbaWzTOvl5VLGiv23Ce/kIJ46rHugW28SU7Q/cL7A8Blkm9D6YU
Sc908kOR3BaLgHnDXGyiUPVikF99TpjPBtcSczF0plkw2yuoFk4Lq1IeYYGhrbN50wovf5Bdfk4D
b3p460V2S1+tn/u4sg6BG+WnjHAgr+brx0cQdB9sRZLiiq4DusMsjcHM7ftgvbqzDWvOQDj/GqJa
jWHgz91C7mxEEnKyWzqtlXI333CwjL6gi+ZuZOi0ZhJiJuygTYW2k9e/o70SAP1uQrZ+4QdQClQy
EV80wG1Jlnd7nnARy1xD47bMy2SpGKyWReD1/Bnk0HgOivfHLG44oMJGvS2IaTxjx6/CO4M21Dnc
DuNQCkELoAb7X2c+h4KikogBM8QQlUO/4NIDFbw9LhV7MVdL0b+tVFL5ZthXNAeA7ENnBAcry5x7
lvEZV3K5gYXG4B0vk8uOISB4zUpSlg3s80u9dTKW2UEh5Jh9cJN30HnSTVK6A4JfbfEogbeR+uIM
bQ0pCb34VsoZQPDgcyoWdZgsQBoBrOtXO+DQOdd2ABn67p/uca3J6gYAlepJZDWL0S3c6zEZP/Z5
YW0j2CKVLZT76nKDj1wA9k/pKLqhJeWUMMF23ia/yEyaW1As6KF8LY/b/o1G8zPDP9XG026W+Jba
MsJT5xgVjNvCi36WkMGuecMN6wA2LOG5/hm/aJNCneLAGKdu1eedsFMzl4kH6SGq7ccUlHFmdRsj
gkVca9YBoOacfxgSKicPClCD9e/HHN9whuseh72VdQnX7r/O+AA7y4FPqEfECjPf6S0gBtho308m
YIUYKi51EZNxk5iiWMYrIP+kzLnyM4aTB9pV46BUtYYk+g9Qca/way3/GCL/Qma5rM5t0B2rnSem
NJvAqQRVAASLD93uZLB25VW8fBUCP3xog7pXODmIIWw9JjYU/WeOoUsK4g/LspYMgMrCJ8k5cOqk
JdY8tieTLiO1N3D4Ows+o4TgF8bTC2nvLpCn9x1ekIUDwRrbF4uJWJ2OdKS93LPdR4lVpmTPhafk
JXDifH1PNcsCu+dnKyYVLlrSQbQqH/HSdf9ccZhjAGMvINUXQU0zCblrvJ+f0er+4nVtnaCyJHIm
QdOYyBkOKeDcBRVV7xdtNJ/eomWYuVPZx9S70XQU0Q7PbOv4/JXzttuSb5hYJlMlc7Lt+6DndRzl
6L6OgmpLtCOhLU1Oww0zEB8D3vGGmWUsJLhgeszJGIQzyxdhJlSFwPKDXJidlRlVFMmOC0yT+KV1
ojzVPMXAFldiwjRIhCPTL4OZU0PfxK9bhkgoepwqO0IUt84Ix93rjJ9oQGJ6e2JaB7R01tuyiHpr
K/RKpZeH2sZhgX0KnzlomQgBxE2LImQifig8LFW/Btj0+zbJiHM3wLKBkN9Dk6gGJkJs1FqaNoVP
S2rRJ2iQbeK/a2w8y+t6CuQbYS0SIIp7rAqSDjnlYLWAkryU2NwmEJiOGWQfdM8CS6eKyL3T+1WN
+S+6DiXK5m2r2lzTr2s8dJN/QTDesGbTPLO15bHhj3f1P1yzZcovxLFLN26T8LWutf1Uau8PzP+p
+7q+7BuibosVQk7m2XoNXSVI1a+ObM48E8ERxJYUU1+P1IEGBAQ37ON6yz3p7kGI6m1XJyDw4bHk
4WvwSCq8BDRRVUS8D10ZkATUVd/EbAah2DSGS2IuPz/raK6NoheDeAeEwZ+MMk/DxqwH7KOQcUU4
B08AKPIzVTjO9okMhcZdnhB6DHhurLSzVHZGiF321u7tPhWGxU8fPawEV9azwY9p5MQFtdZqNydL
qZc/KDKse8JyMmWRx2E/kJkCzgAHRkTPsHQeetfzGa2vZCyVAH4BWWzMl6V0QNtQN/8nr1dwAzvQ
/5Uj8LdffTAKenA1mb1PuhxeTtD89wuzCdTm74ETcRxmu+iRFggXlxpFivVGX8PnJpXkGztzSHKk
i0TZcyrZcKsHIi9uClXGjkPivj/qe/6HQcuU2fb3tY9/D40/T6XlGs/LBXEQHtpTt3RHbyMd6DJR
knNr5bZd/Ad5Np5R+2JniWSKJB3arKoR+0kY2L5ehnXK1ObmRCjJG2Q30pwC2Mx4rv3MnOMUe/Fv
4SC9eMyvP1f/7bEZypzo/IXVk0lpcnl+BJLMOm0PaCinYe5gKIWOdL09Or6+SiwL8/+1lzLbY2ng
JkLfgnF6kzcLv6F9lgC6uPAsMubF9Qf+wgMxrhcNw+FswA1cVAiEMhzsB/9vcAv5k0sWrGQkDYMC
vDxhMgipfCF+W0OLF4vmi+3WTkUnZ9TgEDyzajiGjtcWvekdc0Of7EoASudMQUwK01/geeIfJcpG
o/rS5K5mtBUdvCPxTbYEISAxMUdvCUoTKpweCKqII4qUIPVdqT8dMhmZLcdEFAYiwX9x5EVWg/j7
lwtNciZ5AmZotzBwlfBr/onnpG6sMCr2JCEO0KS3jQ01g+JCnSl8/Qi+KScI+t3IlLUqHMK/fnE8
OknAdtxnGCMv2HQlGuZ3JqZkxuL6pCCi4AgGnBUmowB99r+Bep7Y8uG6vrN5uJy8SkOOCNROnbmf
E9fK+pPoPsxijrLU+ZkfCf1C2GaSprRZgJ/73bAqhZDkJe40EFB0znf2aP7fk+gicHkD1sMbYPSP
kARCnCgMUgpcZuhExgrOux/WOUB11Qgt8Ch71CzWPSj7bcagKu98oeGpHgF2Eosh4V7qFPB8ous6
wIUg79x6hHcgpUgQxWfdjAIzvyoDdTcfEiGbMB9i7DzmdNnx7lL3rAOucQUJm2aKTG7+UahKgR0/
Heu9RjxSGPd2RbHDcVCv6D/du0kt830gcJ/emRDla4IUd06Nptw+YKC9kDy9mzPGowIjjDYdsLSX
yg8593e99inS8N4Ej+xkkHfx8qDQ3lQHiJTME0WEA32R2HuW9YE826bIFz8wzNC7RX8oJmi6m+cA
gxO/+t0S8TCdtI0jMM/hDCyfEOf/qYYh3PK6ziwMFsseRdNeBpk5W+JjHv6cKwNSPYT7s7clms3K
cYoLOLSeycwJsphGFh4gGBFCpmaU0B6ABNYgViHGr3ToJgQ2zWj8NgN2MmC86cOoZTokSa+XB6mM
X+uLNiBJ9lvOWoFxIMryE8EiCK6i+8PTX3NAPKMOcWcG7sYGCizmGqiKj4aqiDwPSqAZrIaBiVtb
qw2MmgQcxdDs3Yy1O3GQJMHfhZdRLub14LYeP02LGaWMMiGRSY5TKbxOIHARwlAg8zZIgJMSWviv
oortkvO+ECEUY8UW5MotHp1+kCwQ9uBG8JM/dONuhNx/7fK5fh24Jz2R530qyfEdwn44ljT8kulG
evBTAj6WXaf4smkByS6uC+vfdpkudxzrjUOTxhXLrjAeghUydDTkwPYurbhynLK9guq3ducgIfoI
KsfqICAuUVUWct8IzNnen1MjkCNAViLK+Nhg00MJOd+55kd1pNUwNVypS9/fOMM6eqkocmzat7Tz
NEWbXsOQowOzeK91oliuANe/gFhl68dO+qlS/0QxePVEtPHcJxKwOBwdZuGZOEAdiQz2kUuOcrkp
Oup7Vs7R/NdEBTtOZm3v8qTW+vA0y4gGosbggpB7UloeEkuW101MMGIdF/dbDLhZHtPurg6ON/eC
SiTngzEgds1MVfBVBP1IxaYk8NFhCrQDjISsefz7rwXT7Qfb7TQmF9dZOEVpNCP28mYbwsAsUx4T
QNCcj13rV7RlvSeC7IwVvlzJ6BUGoDeodtB7qYWrjndAT9eKpBVn6bK6BO6hNxrX1hygt9QRiMt/
yUaLV20ym0iTkdPDs2JEdf6LgVIGwXJSwwtod8Pcef96AEKxP/pqUWHqRY8Ia+uPkZREr35kYbOh
j3vY7KfvTPJtJNC/xNwP9fUOw6hNkpN2XYXZNahCQsrxCxXUWS/YQSmhDy8ze0bijnbJm6TdqeTf
0rNjmZxp6nwYKOPMm7N7PFIa2olSXOK+tYT5CSv4zNIZ0RW5oXDHXB1TdeWymfZxhC2aTWdp2FB2
5xqCoDvv4dcgnJvhVywdjkaiPHriv2emkun2NzyvgtZLNIbkNHuDk1QNtkPIe23YWB09j4sbjL2W
VHhmKrkqcrdaAA14PnKTqBph76/r1qN48GpF47MVqr8v4dkYryzdDFu3YrQ7Cheidpl4NESiQ6r9
gsmzeqsM52ydBYT9avjZ29/KDqC/Q8QPZ++P6XB4AY1FtgvGoRHKOKQ0N6kUiHnJMVf4RZ5sO+by
NQVUzcEaaAHvuc9qPVGNxzlZLus3uedaN/26xxGcUEadmTrS/kDO3cw243r1YKH7uD94lov4835J
xPBTtA0TVx+61VtvYD0LMxLK8kncWKJ1T9CViepgwx2uDVItN6a6r7AKAI5v3qPm1AeIvzj/gHdx
ZVIECRAlfqeUrCi4LfwyRHHjY2ET7Nahd6Psbhii+wqNeprmR2/uUkWytHNZ+/CD8k9qNbwoVVPA
yP9bXHXCXctmU2EiFgcQDFBsJgbCl9Y2lD/D3bRmfgjxRojAQgT3FrUvGsNEfVLtx7RJGT4nD38D
8x0FyqMSpPuWxNh5e5gUGvQpwHs2jtg2h6Uch2NUP3xWmC7DSk8QnF5EEOeqBtbrXhxVlsXlW9J7
NHM5KMict/V/rtqsBtEJx8IvwRoybZTNPlYs4kz1EwLLlsEEP1f5mVZi+L5EfQX0OtTJ+nTglFlX
LI1ctNYhhplc57+eDf8OEupBw8KL2vaX1eFe3M00cTPRpXNCJAQUIA3mYlZvJe+UCuljhf+WASz0
LgTw6Ul/yORF6Oay1/0ghvw8RDNLAPYjeOo//aQ40T5m7jSrlXQD9999dss1Qxeim4QMnQrjLdJ9
Orqy8qTDhuTSqIQEap8yFa05v+6QQHhCzpVw1ujZcJ5sgQUl75zp/XMAT+GUs5agu8Ac7FsmJwrs
PmeQXqI/4k3lF1BXRfzewArTigz2F9etOpv6KW5w6zKVhIIiAl0NTZ9y9+xEdU+62yVP77BQaepj
B5+M+9BUMIctxcLnfw7z6bwS/JcCe4+xEIPxPJrYDiV4gES+5e1pjyvqGp5+7Oda/MN7XvB1mzpN
OkpGh6DBQW7P/ajLztUVJrR163Cl99XgacLxZTBx8duIB762lJhl4R4CVFjZtdgR0pP7R90hfqr2
uHUOyUxX51AgYsx22LbPQcFdboW+lCfj7RjU6dek+nmWFdvpiVzuMN6Cdz+KjXpU6duaI4JUbEp8
AVgvk60ZN5XNoEnEBo6HTuMENddcHkIj4vhnlGUI2ge9IRb+6rdGIwPvGzWD4C1tgVs1ElvC292q
fx+YT2JdCZTUhqpthgdWsCC6n8DoO/Wkcaou109NJjvnSzbGCWVFgEDnxVtMLD3kzQWrtZWPTVwp
ROEc4Vmzrw3tllZ1Hfg/nTjKa+dbYqQfAfQjrzdcNG5Pf//EN20u56S+vcWGcWYPbG/cbvogqgZa
dB3/lGXGwNyvyb9DK5l1vyyKZo3v9xxSJhrb2XMpnqdOfkQ50U7HfnoLPscNgyh3DrSc3qREGmgH
RLJdMezmQ9JP/rSj/AxOoeF9HH/DvWbwPQosj+7CgBVyN++X+879n4zl4YBMncWvjERmSXbeGHOK
dWI3bAymCze2WMX8/nlfQQ+6aCG8NWhrRB3ZTe2+VqZpHvuc1fR41CYVO4EiqBPz3jkfAsyHPL/p
3c3jAYnI/AmjEKT08pE6j/KQAG8MA0Tkzo47xPKSpJid+kNZqZIU2oBZXiZoTPVjMlctpFGRXX+m
V28XIsJJNaDAlEWyJh+gd0rhNjrQv+KwSc4GqCBkmFk06Gh5FLq20j8zmgW2hCVN16lx89Qr7DRx
2Hle4uF+XzakUodf/SuKlOwJKuw2RJwNlYdnvQn0RwBlcJ5GIC9hGVU0ipVAFXEnnENqcAxvdFSZ
TRRpj6uKo+gyXMo3Ns6taYZup0wV1Wew4xcZ4SxOQm7nJnVYR0cWEV2E7j75N9jp6QUtHdS6gPqA
fSKZqTT2cngSPeNWP+XXhywSAW8/HW60S8RT+iCCiOfmlc7T9qY/wSkKUtRel1h3oxHtw0l2Pzpy
qcCMN4HWgY/1QlFwYO+DjKw6RN3Cw7N/ZDNSZ0+lTvfLzfZEvo0YPFkMO+9ZB0vtqfx1on2Dqsrz
ZVf3tCXjIT7zPUVjgR0GkmsPsRp1DTg0AOLfvuaOYaZIeJ3JDyNS0S2i3D2OBL5mExnxo5bLCXRz
mKW56fP9cNsVHpwRlgqMW9fuR8tfjc1cLCVTz0JE0G5qcbDELQhfYhZUuvC9XBqOiOupz2CRUZPG
Xqg1eOaAvjjyBA9IMuWdWKPBhoruIamNI0nRDuh95h3SluIHcdwfC7GosBbaebL9FvI6SWbwSbGT
fCZo4yIdujwGN7jiYgsCZ0U1fzJ0jFXQjr2iKsJrlo0kC59u0e4mtuyZB5cjmvMvrav/bQYAJxU1
rxn/7LpMCyhRgjrzK45AXNjaGbQHxdZ9dkbUuZcB79cprzZMATrHEgW5Dg4m2hoiWrMh3rjqfJqd
uL73eH4LKbkWGsP5hQiCFylp34Wb74w3dQvjoLBy1xAbis29kaifqXSiR3CrKytuWs5uL3sbxdn8
CIPYYZ4V7GON3AhtRllW+nshISKVgu8AHJLZN0i6tThFVIfynqPUc4TugsAKJfWz9gvrZr+i+Toq
48cr6iQPQsvmDGPGGsUlv6dgpizhTnbMhcqxHu5LiZQtYdK5W6xvhvBe3ZEr83Y1FMUCB99DCFua
l8K/md9bdJPgGlPiyOJSoGmKkzCQdxnqbNnTgVKWO8e9nnvM66aZfroQ3lTjeVRBfxjR3ewbm8wR
0ZM/2cmk68km7S9I4/Z6c93iClCgJci9dzVsoX5FzXGgv+dcDIe87tNq6ZVrfzHKVAtEMSllAz5r
Xta2N4P6tCxq+tzzqiz4mD/jFMcbjrDYcNpl5YuludGaqGyjNVZNGN568Z35Nc08dW5oTDhz9bDX
mLtA/le03MC0ZXhQSKnNfOppG15kAUgQtx9d3TgWkrudq+DItLe1s0K7tC/G5vfH4cPyEdsbRXC0
gccBdz8g9bMAfJyy/fGdx/VJkN1pjv/T12z0wfOvvwrHU3hC3ekW5GdKnPlSLnJHLp2lw/ha/Tqh
RBaOV7yb+REcpeCDPdwcSGIP8ez+Nz5sgcBnFKppM1p7rFkrw8oqShDxoTmTDHw9L0AQS5GmZwnh
k8Lj9pUN6L4yNKboXNs4hBJfAT3TQHeP5aXcsWyAVkWz+K5ki1Rz1nhtdJ5RkuRI+UDxiE944fmE
qDzRYbBPvIKntV6DNJTgREcZxH2wwjMkdMh//ShgvD2cazgZG7sbqlExqzf9AieRL5VGLHKXr1Da
B2yXwUijZz/Z+57OVUp377x4IQV4aV0LiC6Jj5uNfvSuHopgVhvtuKyL4LdJGI4e9edRoxgau6nf
1RI26aTNUnIFLdmNJA6J80ixK3poRozdcQctrLoemmBiVnr/hkhR8ZkybH+PEUEQV504WH63zYVP
VNyqCGaWH0hyL+r4X0IghD4Uq/J+L07W89aSyE0S8JOShONveFYMlq8b7WXVP6Be50+czPS/4KWw
JFAItXqLjLV7zkj3hgTgTxR21lPxpeYVg+0qNjTrLnmrm+6p299JIh8kp7ArWuJfPGuOMIg3EOsE
vzMN56CX2mwUN2GBPvAm7kMtZARV5yHE4D01IRhKTPNdCDEqcxnHzJVHxtMV0WJLuiGnhe+xzPvv
2zw/yxwoqrhZvJQG++hguzt1ujXnAjZX52//LPDvIWXjQmHsPvsV9ApEi6cAlxFhB5c/dEyVUGbv
fmTrHgLpFvfPSxZAQ7KjehuSwaHZNWUvmMVU+C+Zdka+M2aKH6x+XE3Uxz5+lqMgirRYGipUbvTg
uB103MTPnTrc7MfaQiFaLF4OkRysbWF6NYEjYD/uxU9kPSV/BQVX+RRnkLX2moji9VvMV2ou7Twu
vcJy7SP95uS4qzB9CMO5cBk6rGzuedGA3EV7k+nIhQXMgQNwLen08fzVRio/80/GUnGa0JYY72Fx
X8KzFxzretYMxpo0i4JPcUuK7Ra42dAWUz4xACbnqPAVcLCvHe3GNMcN7G3rhug5KU2RjXlesAoL
ABzVBYjPTk11s7o7DwkjO3pq9ebOXQ/6k+79+I7It6MDhwC8B0NWw1BPYCb+HNfqLiBocXQKIbk4
VRcNOZR0+bdoVO+VekMvpEMCF1bta97X095IwRaSI3i4uFc/5zfPw8dHBBQcgMMXuSKPnY1Z8YIb
5c1gHCqvmuP0hKIV5cKqjbr+PmuRSN2DVAu1WchJrAUX7VO0TZa+IbqYZrNlvho0vJay74FjO61y
qLos4/46G1Zre6+sfMeULCP3cYV/h1pbSIdPkacU2i9WZuCsELdDZQ0+XICv/A0VU50KxWtC1cdG
L+xApWE4gS7+q3dwuMGGz2lTeTBTdotLYK/3CquX8+3ju632/2OErJau96TlIMHYGJ0I/yMyOLqV
FwJTQ3hgGvT4DPSPTwPxByWAjieo+HcJBmjgbRfT8G3LfHA5HJCRNfuNbZqf/hpWv7jTxQ4YRlS4
CB/c4AUAHwNU+GWi/V4lgrOrDCpI2kmR0JbOnjC53iEARFEFwplQQiLg9WJBfZYicobaWGEZs5JN
sMPFo8hhF57/aQQlLLJBtHXdCgTFDPp0Abu3lSbgT6xzWSa15JFJSRBOvkwrPh2jy4tdbvxjUEid
Z03gT6VK/16S77PSzIJ/79NO3tb6+iNTQMVQmYpnT8maPzSQaKBwqz+EydPvDc5n/ecGAFIn23SO
c4CgfcLwk1hNHmeXmSyaPaBRCcxyHJMGHMAaKaS+st/MdeZzYgulju/xrRCYH8F3j7TYAmg43Jwa
C5D6NpjYzUhywtQLxxxtcpjB8I+bKVRq6P7aAjorsm6YwChxIHkDeqP655AObeOpayISYrNDoiMM
qwiahuVBXsGh1EzlLzo7kf3yf1Uadf28LJb9tQoGLjMFcXtwi0StKJjkMIjhqCCvzvYXI++llaau
u+orHu39VAPkAPsh8kDvbqC1ctVoeAoRM6VvA0/2zXeUUBlXa29xjWc1aMdwQkNmPpyAf/Ul3uD3
SKBsHsCfr8TPpsG+sEuRiLfFHYBzTp0/rRBwS0iM4ETyeuL+Yya/4thbHrL7RFam0NooK5v3OEbu
6d/EN4bV7++IL1XkO/gV+5daG0pj3G4k3P70JYUU+ikC+EFqToAfmbDaUF3fIywkW9FBogTiOYQJ
blrecVdEMDqweoPGeEClikcOAhOmr0hVup/l+JsoXNLRL2UlTToBjdO7a1TW1nPC0eN+dmJQN0Ph
GgDYPbYWaR58LmjZnojY0cMv2tn/Mt+8SBcghKpIxGBu8NL0BnhAFODFpYw3VwJpjgYSjn6VXYvW
8qOaHKZ7LLF3v8zrNKfzhK3vpz0Y2DU2VXrJxe0zMEy3bBy1ScGu1rFUh4Y/KiJ+vz4N+KqWzZDy
WVA+1EX5JWAeHRV81Ni0/NmzOnpBKRvVnIw2HvYEP5zJDx5oXfiwVjT46siH2eSgutb3hQWKypvI
tiwfcHmLj6Sae2QDHy0QkhZClPNtKgSoYBNNCHi26qajC2Zoc5TfxRexH9epZPqUZobWqjBaYf3e
O0bqWSVgTlTswFC79zR7yih3kz/Ml71tu9KVRBDrlHyWxL+QmGYi3Idhuy0w6WkCPVhotmFi21HD
1ZCQ0CIipM3LbtOhPuRd+WCH1SIViR5pID0Kk9yAkH5hvQSgEMhW9iBxrQ6HEfVP/EZTnyat7VzL
fwxIb43YYF7WNut8o/3DJ4OhL9YOJwblxATUYkMhqI1E6yI38EKu3yPBL1kNlF6yEAEU4pT8qGRF
1oPuAC27YpAmfJF/IYBoHAnIVGgQL8HPr07X4dZJbvGfD+2XG75BiocQHXTjFEo/ZoUF7JsuGLKa
vbFdEMq9NDwiQ0hcuny4ZbbyBvVWC+92+NNQdKmJ6VjKJOVsKhsLhlF5Np0h6ON4qQE8VsDv0CSE
rown9ZG+zZDhzYlKv8W9MlhQK9l0SviZBcWDKhytpHPv2TyFYjHebYDBeIHF0/SNB5pxcuNcGDqp
QUKfspqQIghukxR6R0EleUHplDXaOM6yvVmphuqQlB1kXv5s09FNqb3OZUDRoxI8vDLXMrJ09Cv/
WSlWK+LYk3djzwlFSRkwyfVi2VfvMy8FvZxO15ktz4EbooGJFzAvikt0gpLCE07c+webFR4YaE0u
34jNbjJEecmW3P5nZVnSd7ABzOLeeuuTej5fOMFJX8MkpyQtcS0fxJOtUEQr0qT+gKhYnNTY8aOS
6/Rdv5ehUE5u+hU/EsUoWv9/duaFTDIuEC2vrl++TwWaC30UXL7WkTF6Kw3OsgArUEtHBSMgxy5S
MRjlMEb2anXPj3FwaAcECqj+29BsGk59lQxKxXIY9ePosagVuOgaBodXe3dGJv9cQB2CS1YFfBXf
dYT2BNYS/ap8yNow8cztaS1X7jyd80308PyheMUXvqpLZy2jtCmIgNfY4rkmK1psJTPRpNJPX8zG
c33/Nlp9291FCHDsJq6HRyONu9Lv74l6GJA/ECpX190ynleFfdRvtkInBlMKfb9gMfvVUjCBKidB
D/zCm4HYJ+RCPgVl1p4Oz8qdIl6lOp/XiTKcyPdoGNX7ug2eiCQXzcWF+v5qClkPX1ECx7vC6g28
P1aFsIw7vwPUbp5RophXbP/N3R9TEZgnRegZ17Y+yc3R5HhKL/JS4M1dEEYgwiDSPj92gGONeIPh
z5SnAEds4fcoquvu+RNlJLH31q9uGFrAL84uOR5yUKBFnJFYapOUhQx825ct3Lydru5NssCNhK93
52c6CtT0nXMVdlT+9UY//wEZkUZjohcheSJPQYq9zdOdztxMCmxamziWItbgq47rsxbe52X3zjSd
rPbo0wbr4WRHGnqQUGb60Yus4XlnydESnJr4T3z4YDa9HXgp127yODLF6/Mx/JIopa5PwhBrehhn
qc6MQfvr6WYPHd9igGzJ6HH4KV6+aQBwFrDeZsuKMd41jGEcCwINmfG1SxwILoIoa8xXDJl8atSy
bZnqACO3ih/zV3jCNP/QQWFHCCnBOQ9k1RbERj5wz/KDe0mTDt3aS9S8CLcxi7VHj+lyxrdKSH/F
Dron+dZbuUQKHXKZkbAhNmr0BRolVKA8C17zI3C2ebHaYHQf3QKnhSq7be3DDTTsv0pSEnzQrA0G
oBV9+S5DhmDwy6nbeI6rgE/sHqGwhdvrgnNl5GPwpcPT5adrl5Bwys8/Q8VVFGPeFQ3eJeM/FmB6
nPgn6wWAMpF9DxQnTyTsUajKgBsp/gobzkieyKKMlPcsK9DGC3DEzGsFJxGH1egQeYWBc8PYnZFd
Eal3K0swFn1muuwIq9L826TqsD5/m+Ij2tHfuWIMCE34donO2XBZRAU8eQifR9R1iFsZhl6Al357
3wa+jUJmp1Aw3gyuYdWzJjkgvQD/tv1psUTUULaMvWCg8+KAO3Y6xv/hQDytm7NOSOPrIrKSfDPQ
B/n4Hkg7wCushdS3MSIvFyscxveym1DHaxm4KTs1YbcYn1ZpjMafuNCVFKPPX1ZUcIBqjRZrHOCS
a+WYVtrkKzjhZhqqMWV2U5m4yMOJ9QMbBlNoe01lTelnJdGpRWIotiBh/qCl2Q1AxCazMxDw43AK
ZFtZB214v6LOA34QHPPxKQUdTlK2dA4K2h2bl/77RIxZgT/vm4URYmbir9Mc+3q4m+TXjuFTahMk
8UUOP/sh2QT/FAB9ba7K01RC5YTAgzDf1DnyERvzVxttJfFyPLF2061N5PRREcDmJz44mcBaO4U/
x4+wHkbB0giaANjo4mKc6tsuQr4RgGV8Wi7zWv+hC249di2V6NH+KZtP741TeojwfW9JbPMYXQxW
V9aDb6gcSPaP3YiyQ5wPfz+am0gu2Gyjijm2DNbinpJct6JzbIfsa4WB4parDQMdXmNj2NQlJZN6
xr187t8TUr5dmTcqM3PAOMlhzD9qiL50/U4tO+hfvHqQMuAemYAdBEVbMDIA8SqTZgXCZ1gdlwtE
pCWBDdZpyeXmyDrMDOy2nleLNcUz8i82Y3R9ZxCMEN7SW7ymSQKy03QPVoZsWzQkuO/Dbi0x6weo
a24yaI8G+RmKY8UNz8XDKbp1f39MNNB4YZjke9GQgS8qJHcfh8OzfO1w2m984VJdEBWXSuqAz4fk
dtL4D65X9TbXzxNe8K+TksX+3k7yRjfr8s8Jvbuk6OiJg5W+suzLP2NQOCQwFr2W8cwFhY4fTY/B
eK5ehT4uzBOPg6sWmkpa93zWLrpWYJdVD8UCRH0VELIbx52U+Kx1wVynRtMPE271r11GV1wVrcB4
M2IsWtLy5e0XYL0znalQTya3mwNCcNQPdxfgzWasVn+Mr6CnVVVX5c5rarYYam1libcsT5PChBVI
LcAOAoInBATe2F6Q4ia5lqTfPp834LnDPBoAtN7VFT14NEO/fvA+2XkN5uX5wzdepBbcu/WvUbSk
pAO/9mDw+Hgdsx+QUv1ZT4Kg57PWmYfkgrlnRLhBZTFCMbXFsQVv2i2QutTS+SFhdfOYEINrv3MM
FVNluaAmCsmjoB7HwKVxWNL51bFQ8hiipGp6bbd2+Azchfo6Roj22UkwZ2ZSevffPIZrCPVpfeMn
m0TZolJcyT3kLmzHUiHnUDII0HclE6O1TaogNOSsCN+P0lvRjIxoiyKhWsrFp9FoRfBxvInDfFPb
pJhZLVGZX1FKbkMrCaGbbc12ayGWgNF1m5OpVFw2cxI9uQVtKMIubEBfP1ehGBmwFu263ebYUZKU
CQTgjs7Jvqoj9QkQqLDLkBBEHZ8wF1J4yyhXDfyO/zRCtmmhXxo5SZchQk/OEs53s6yw6gxOaX/R
dZWWc1HAgVsrODRmYH/pVOvtDrkI2yGs/2hIQPU3UB+UCg8VKEGtfvM7jPHcvzJA58W2+Ea0CdqM
ZU51v5+wre9z/QKqNtOtX5kCR3KJuP2Sc338vvc4nvzZ+Ot1znHxeWpGi8kGPEs5bWqtGLAiMGEu
WBPArO09ixz1kpMEouLmMvfavCT6KN7HUqnCnckQwyUp72gTVKw7mJlEJi/CNojO2OXtLcrkvgjN
mw6LRvUkPsvnvdU7Vog3ILB7Fttnd14wiYa4VZTKhcuZ1puaCParrA6w+UUq+M/cAjYrWcIw/IbP
RvlP0UFpfAYQU2YhZf6L7H5fHytx9fP34PHZ7ykT1WTVW2znFhQjJ1cUuq1+a8mkOmkKDFrtiPSO
ABtnL/R2XzpMkz+i6k+jAvWJY02HAL2VH7xlFTRFwmXW0OPOS3kfIDH9oa0T7MZahuU9291+40vz
XKk8XHBFUAtlBfUmKXvPSDubKWP2BDeGyFWeWuh8JzupDhNSwP5zBf9dEOWFxR98tIH362hmH9xY
GAHlGlMWtv8cRP+hSTciwpS87LyOfltOdIbhqTJVAhebCPDyv5zTs73JKUvNsXAqeTQ4PRL0qUa9
vSAqybI/EWYxNZOOzNMUdi9mYjTXoALJTf6mbY/6LOzOZ7wXId1g13nKI0kNXVEzIbUFjLrwYGsD
PHkj7fFnv/j7kdyr/YTlb097kTOIkUBfCQzGRseMi9vRXsYVVnqqEiJL1cjlCnZjJkXlJDIH5IET
7ZEN05NrnL9nqejRvNerqY3l/csqsmJaRF/V6jY47RHwvGakhRqkCIRL5UOBkqV9t2aXySl59yr2
AXWQ5kq820BQ9+l2eL8IUPpJGvB6wcYMPm9J/22+0ocrb37Hqkw3zGKJYD0rl0ll8v7vPyegm8GB
fa/XmDg/Mq/bmZN0HbXvd73sEwi6je/H++nzZg/Now51R2RWP9hfop5fYqJn6Nw86VNptfZ0TqSi
uxvjkoCAbEdwacnrx2l1JlQFe4UN4C6ST+VLVuI6YTxApp3OGcYvoIdJ+8HPm5PQI5217PLlaB7v
XI5OOL06bvlQKLVTf0F6CL9Par4sQU9zVQcqmzfordgAGiXrWzsfiT05kIOyxIEhIDR1XgGlqg3E
AISKA4KE6RjfyigAYt87N2fqeO7PL0/GyfrQOJQmb4MCEjAaLUB04/V01UdRJSNCd7tp6wjoRSlh
F7zsJN9xABbkXe3YSLrJNmpKCWQonCbMhiTZ2/0P5tux1OhqG2KHHsf6zny2xmy2NVen8AUGNZJM
juHW5WVeR6cTvMMbwQtMPzOY5fjKhboHrELqm9EQXJkZAZzPVv9xEnlq4OnkuNjsXa0674RWGkEF
6JqMFu/fVtrxf8fJ/BkMz4JbrIUxacCVxPxqW8fXP/OUHDUkTcBJTUhfQ2bXQNsmJ1r3g0dkvAg5
isS9LMU0BZYTz6IiCa5BecHGPFGiVH1t21i9TUdyY94gEmXn/D3yFiA4jhAFtwv89gY/uxM7I4ar
CRCWqEUDJQll3A5D6ybBrP9EMSicekJsdKya/CaHqsXIOCTzqHWycDDwr/zTMcJ1sfhwsvp6t9sk
0oqg58CZ1a7fCH9yic4NOa07w2JS2S7fTQwYt3qz2ZIVQbtidSrNVGQ3tTxZ1rQJKGxbZznG9fLq
2dIoBfTFOLjeMtS0l0vG38H9kK73UxJLIiV/sdBTb61WwWHJLFxNpn36z6/gl0F8/z4bNlFag25R
UFa5EmgOEAhxMWXuKgQnlRYFYa9kHei6ONpQFDAQdVVjkr9Oe+irY4u/KWzOZf8ykFAJbrAKfWSp
GCNZHO3v8v+nfnw5BTVbFxYyUkSmlxQReYR2U1FVYGU1TiERfv3VgPgw0RTA2B4O4BVaAjjwQ8o8
pMpkBpFamqBugaw1fbTD8AUg8zUBlM1b6xaTyOQHe1YEZnBHB+y10rXS7FUiriMCKzK8G0lNyzsF
lK/5XxnMnvWp/PkzcHcVlUn3M4rzz5sn7N/Gz1mkPydqJsI/86msCEEDoaECgSmOOAB8HYTDEYlS
qJ3rq/QELfn+F2g0Z/1p5/xp+YpCasCJ7LAZJwQSUyUN/p/h0IN0SBIWMXwRI16GCQ+GCBqmzmcy
Vj5Ho2DXqkKFCIfJDzgttCrifkIorILd36f60zU9poXkpq7KIjFta8FOhtDuVuPwpb4GNLalgbBQ
oZqDpRiKSora1M3uZrFX40jG2h8eJhiklbpqGM1XmTvc7aVU82uG+5+ccJXohyCuqnFk5DAuc9XN
NO7P3p9fLhJzd9kjK/lHr10fKaYzuHzgZof0rZlBeGT+yje2IQouTJB5hUCj66NYa3lJvFXBtggX
XUExhjChHvWhlkhQ8tcZF+dl8myp7m2nCChcteyqfgkhpI84Kevr7KOA6SlisleHyaD1WEyBXWNz
yPnAwQ5qohV/gPfR+IYE9zP9VQfed77wGG8ni6Lb7jVS3DESXTBe1RObn6uZ4UPFeTErOq2VvpKB
O0SqyD5l+OG0KRuWxMlYsILFAvYjzISS9b5TNtJy8hM7VJnGUEhmiwPKY7roX9JeY2xEGklixzvt
RIicA5bel+gfIZxgVWlDTeu0sn7gkNXLxf6cplNp17LhAFU9UFrn5JXqzhQqLi93HCPRPxvwgsMe
a2PeJLgjB8EBYrYoH+BiRC3gbACWJZdCS0/IWn2Q0rWQKfX2OUq7GnjzJ3656w63d7r3HeCKkfnW
4xEhNNMkZhrDbcelTdDl3qNE8kEpMV6ez+YJ5x8PQtzTM0CqjhBo/Ex1C5fNyxMhJrwfzLQgaZQL
VJuITQ9KO0cAghYxcEVmQwcJ+W56nkCvXCJFbmHwKAgQT7KjRaYegT0YDI59tv8qwU5TZsMHW1ng
jjJlGGxZMCTIJk1DhRaKBdjwYxe4uHHsJImNxEkjsnYcDfWHRiWBAbyon10ORWVAuvgzDvZBDTzh
/6SqbuCtqB2pBqk96WikjejbzKjRmT1bsq5TrAPJdOkbAZ7cIEe0H2xvNJy2xudj5xRjxY9lXvE5
BDq0VG0mLAOShPb+hjNn1Ne5HXJLYkVk8coa2OxIaRZ/6U67vVCB/uxEjMMwDJ9KihZd0/QPFR8C
rycx32GnH1ub+qNIbi5tkhwEk6kM331x5yTR2tpjxVPJWDnYGcRLvWTQIUKWnLfwoLMR16+wz9ze
JVl4pyMebImauA0OGe2QUBNNBcen36mfhy30PPLupQK8WVQcGi9wtmp2aAeWf6ouWpTqVNMw9MZI
/DmCrr9zKuynoabfxJfRLeYcs0gb7dLxnHgFISaNoFJe+xzOrEmVmelLNAcz7XeIZEoJZ7quYwvV
Elj4aD/JbdRbU6Mlf81ht5MEvnrXT9olluO3b3Lu6IbRq7T7Yi3BCIPN2hnPbJTxtVKUteo2dPgk
IngTYfBfSevKpgbvTjqqnpI27EHuJL5OulJAugmV7MjkZ5C3cR7vkjgZTrqm8//PT8XN8m1SPIPw
bO/TsWNJiGnh5vyU+5B2gFT6lqdnqEtUF5O2GDCqc5QrLdmra8EKNglNloGehBwvhVl70g4YVH7F
ah6l0kjXaJg94kCcAFB/rStxoIeWP60VnIT+fX/C8+OBa1veQmle1ls9aEZPQiPd9mfs/EU9BcQO
jGEYGU9Ztvdtc3QI7d1MXYOJCJ5+MdivXABYHU2gvSULC77jGJM2Xz5pY0Ok6BTC7EFPfmTM8cJU
Nnqm6NGA3uvgFCSLEt5jxpp5/VJiEYsGhlc6joJYYFb+QOFShUgOc4NqEkLu5CQ28AfgBspLnHGw
3a1dBKTFCLABJg3w7itPid3PWRD98uxNz7+bWNg8JqCBAY+AdXuiFv9xrFloS31MUOCi/VAJG6Dk
XopdX64qHvtdSQIbUo08iWW+2VLKvPsLG8YJTXx5BqgRvFsE5vyNzft6a/GnbU4K/gdwBmnCUijg
MOUuccPWiXc4iO4qZtx03jEPJ42ENwbivptCHAic5cHQG01n/eAhs3C7YE/87H960ue4A1faY/YL
Nwe2NkclZSfs+BrNBJAaoeUVImdzIDWGC1RS5h5aZMW+NLwZGQUkeEKu0zYhG1+qpl+DFE6lUG1l
IfhUKdwzA0aSUnAfi3JC8RBSf5j30KUww260YC6b9MhdwG9Z2Hv5NEdZ4ddJWKOqZ9MC1oYFZndn
LSNC3v/D1axNvphH3M+ybAgn01zplo6rVtNl88bJHhE8wBllMO7nSA2JT6miXLE8jbtL1SivlWO3
Tc51Xtq20AxtLjbLceB1WaWWcXEyp75EQV5guR6g0aBGGgyF1CsIZmw1wuY/s8VO0T1GvhaSHgMr
38a1va147xVSA+XFywBLaael1ZGhKZ2oOB4OoaHxBiiwISxkQ/hUIZ5MsxS0Rnbzo04qBRMsK3t4
XOaFDU3hP62cYVRdgxgp3GVB9RNGzirQUpGESe9hSh7y+P3lqHhvjl3vsh435p5L68/rVTu9Vahr
ZSjxJwH+YpwCMcR499JxyCpQcGgaYgHdzXU24nYyIzRgjiRBwoOX919XhRF1tJ9Jz7MGTqGVaQlT
Bh6KUgbBgHSu/t9B1j+k5Oet1S+62lXQFFQxG2wLkigvn8MT0HVTXR271z4WnJkOSAIRWiynaEwE
UK9uFIk0AnksJuhkoZ+LxXb6M3wDK7ICl5b5/MCs34Bd7jO7HYZ0A4PqRqjFdi8sHYWiCvcNhJQc
TQAySshVANUm9Hy+2kQvyJ5BsYK0Kww7ud83gAKOCNvV5lmSMtMAosb4iQeJd7i/OSzMlws20kez
8tj0L95jYvJF7PkCn+rDY6dY2308XIYBlCmCIhC6kA7U3ejRRDgmzuJDcsfkUJ9roD3Yp8XkvGac
Ehjp31EedgZMWlb12H2m2N+3kla4ph1k26a+d1GOPayhgSP8BqN0k8R9er7VgBCatf6BBZZWD9qy
Q+tk1DtGoPAYBZ3eUyEDmFBkB6wJ+v0I7h13RF+MlQkj5j+M9VSyznwBSq4Jf06UB8apkXPSJW0+
8mxWW0XDksBnTUAWL+scpZmOzKMu/vfYI5b+osKPeTZO61Gf43hYMNRXuOkCltdFNKKdNUdLtu6B
It6rWSadSyvoFYZMyNdliryQzCe3PujtLfLssOfKFcuUoBQ8Z8ut0ZqXdZAn9Pzr4KoIJ5GmszSo
wDEvA0Ttf+y01dR98x3qacUaxbBJCCLmZjN1vw7FWW4ALP8VUWYeF2l7jXTkWjqk2Dimv14U4Od9
rjvKrAxsbnT0otpoxN1FZH6rjOAPs1caXwUf0AUislZSPyj+cWWSfIVYubmR1PsMmK1vM7HbcQaa
SicmlE4/6hB5L2CsXOfGFZy5jt5Ra6CBI2SBVIRDbQaYGxYJj7pJe2rtPdi47I6a3FEUpHyrUzVD
lUCvQTnvwxnSlJNSx9tgSanWMoQMe4NENKR1y1pVnyZlFWH3AwJv+EClWqNOg9i8AbEyktz25xcO
MkDfXbgONTrMVglR7v+DW4khReOuHSXpQ6Gpkp4E0xOHyIpbVYHjIdUFZwV3YqAqTA6twh4UBt4A
ZiVg1fsTi1dbdktIb9fpkLkqcNiCIT2W1slK5niMgKO0eRwRKxjgmicKTmvzPBD7Cw9XC52YQjWw
iNx7Og/1iFdrelgW730ZqjQQ4GV0RVcuufs+lLB4qMiqbYOPzeCSGk4lCWxxDvAK8ZYzcDs56eCp
nWH8s9iFp4v/0NqeiVka4cy2NXCgPWSicmrMdU+rlVaRqwno8r4B/mUpBA2w9QTA03n1DYx0YgSI
hb7k1fy5+ZOBTOAnGK1I9BFdOBr/NI8v3tE4KqUCeTYqERg2u/3/lPoqxZguDQtT8N7RAJ43wjp0
KJFaVywj8Z2UZiwtCtQYat4VpaLdGjnh5g+p8eXLJq+tB0476Ld40WggQE0SFyQSER9CrI2Mggfk
6NwgyuKFRzGUGogSH/WjL0UIkVGEvO7LqwJ0qDL0tDIFyBZ9Koeol/jzXHNF8gEBLTEvh1yPwJd0
r/LAqRVoBvmX1d2o2G8jwETt3KZI5uPop+ilePQtyt6z6hPUmIUwLUdLt2cgH0PVWfl4ewgBrxZZ
udhRtLzwzriZ7wCGcah7+gG7BJRiXuMZrYiVnpnVFuZzAPDFJXOKCS31vLPINgJ1JRSJBOgWxty6
RGu7ePs0HgzfQxKjVkUcOequrTvD6/HFhKGLL7J0yfERY0UXsGnAdQlIgYq8CYXAStGr+Kti8Jz/
afPJcCXCe13qvvx9BsKMs4Q6S6bcjz0nlTJIPd0JKDqgwAcxxMDMK2MOS1GcZ/6sEeROfjnTFhyb
ooWzoHRa0jylk3o5HrPlmfZxqeG2Wk6tUhh0NiPgrogrpeDSD5svUblEmTUd22+xXIhRdez3r1Ne
kPHWVzFqXtA4IAvbgJ0LqFkf94nkIbFLVVrkY0tNt5Y9QqEzVqcSsLbgF49+oZK0YSbtMzXEJ1WO
K6vVQR4ne2RSM/HHsoNQzg2Unm7wjcKOZ1pDbMiX4gBeugzA+m806K9QxRbfBA2ifm7TAmZ6zvnq
LFA6UhQtQgNtmqrX6Ffhb1zbJD6iBCdz57MPjNrBOgTtyk6YT9wtN0M1PF3IQlpH+Bu3JtMIXGQK
bsWC1rtuW+t+KFJ08VuRdZ97vV/hQyFfKqRiRc3N8TLr8MvAS6pdP2sYuS+UiFrMK2I/yG2RVBqJ
uLtfBruH5+vtHFODOA9OPK6DPCz5WB32LpRQ1u5MEhXXjQ65z69HHSka2vh5nsM1yuh/+hFmFTLY
+cUxP39DHKMFGye83J6TVaeOpP0EFYL68Cmu6HVym56KsCiKU+enxl5ETonN3UWP0X6tWR3NNnLo
zmP1dVnNkmq6UY7UhlwnNzOhpQm/BonPcgak1m0yaKk5f3ujTeLMLqof12q2PJqX/tyMLTCaQdOt
L2TA10yqu6LlIIv9zUzuYLlr3mWwl6l/f+VpjTV7EXMYa4zgzeYy2QbAMe1Fb5/8rslsxUoYx4ev
5wgN6L7vGRcYqVhrrTGif7SaeGuN7yXnf4tRoKGGHKQdvuNIkqHJV+C1ykqC30sb983723tKVhrG
hwjPQUaFgAYZmJd+bw/CNtcfwHNA91D+MglsxI4bRm/+Xq5CmhoTGVHaWSaCGejDvdRyaLZG+giI
nV73Nwzx6eH5cwPiBUNOZqSqHPwm9oOfKheL/AtO2HGGPhLdoLdSIO07BpP+tjOpgjhD1zvB2wZD
tP8KGe+4OjgA+gH/mCtpHoBFRf/+yR5G8BH5uEXFCQWYZYQGBP1NdPIbIGn0L/x9opzx6vY7tRO5
AvIWF0ItwiQcvw/3NFgykZ80NtKfceH3c9MAFZ8A/8tJ45Ul4ol/iTv2QaQK7UgXBUjmnISsTIbV
dkxSrGHVPd52aR+goAjn65p4ZnYHuA9MMWqkLmxVTZcwo+BFtxf9apzjsEBLjhnMdYlt4q+Wfr/I
ADRB+s/GoESpjqXM56AHyvxc0TD4AczelMk2pYXicCiBlKrJZBZhLteAd53gmWksc3EVbGYndXWk
Lw1G4ripC2AbFKAHz7ycvi245uYo+YqdRJmzJkmm4EsfRfqQqHQOVPDs2YZwKPWt3SP6VkJ+6G0l
NnJFamj80IwksB5Gt2II2ALNl0/33rAbCOg0IpSQF8HPFjOyuXkQ8dZQXdCdzeQ9nLxN3wfmOJz8
XqlbxznBAr3rHMc0Z1ihXfO2dAO7kOEe5tW1BwBwS0B3DFNECuY28Y9UbrPud14zX9CR6el2psdH
fjGOV92hex5dk6lBvF45CmI7bZAMI/gx+eMup5HCI6bceVn8lL92iKZ65ngkmP5hv3eiqPBIO94l
vv37t5w2XswsLyHrXw1v4ci5sNWvPQKX1oJWxK2fDsTVzpjPpWj5deVfc+EhLe51zqpRHC6mWrRK
TkrBo5kKW5DrNEV6bVwgOA6TLNPu0EC4sEVWDI2IVH0MVLDvUlb3qEUBE4Z1UGB/iq6pCeLZ2tJ5
76TOVrpGUyoNTof3ukfbviLTVXOETEuXK9LCQgXiQblB/xPZaK0HBnDvfiqqnNcy12qBp709NGYR
WGBcNvMpM5YGT377VCp7Vt5ivNNJvXErBffAWZXWxaPWF1pcFxaxGLwXZ/jhpHqlIilVQmmWfb0/
iDNawH5zZGuF+snCi3rC3rY4zVtxnw03K6zuBcaw/qeTQxmgsSbhdo876P9wQe76+EgPJ7HPPppE
RBVX22x8Ik7zKrE0PdcxIEiUXLg3EJyKFwkFvFaDNRHdLCLarSEi0E/ikbu4bylKfV7YK654hvJ0
FInGGMN5LalZuvYfEhp7t0TOC9CrvYMESzQJS1oVcwSuf1QdSHAvg/0SosBP0koWNczPoyTgHDuO
VUo1qENJdiXmYjHWZlg45TuOPv8GotHusVXNbs2QjLqAFMY9h2XB7ymZKvkAIN/+mk6oCcSuiM4m
vjBHk9B34RU0AS5ee6hsKChCICLTs4gqhl35hRrPMB24E9lxTYb758TzWO/b1TRieOFjV5brYnEs
El1+COVvoN0wVHhGfp6UIVZdBXxHr7t+MS8qD4+ZxNm52NE129ntTwl4QPDEX2fJzQ7kMnvqH62W
+PXOJ+QAV8+97SvHFfyEXYSga8fBRa7H0xh0qDhMw8Xch/PvaW86Osei8eRMLL948fN5nJVZVDnZ
UADriOUv2GCxl/Wty8Iqyw0GW5KwAUOEgyPWV4Fp25sU+tUNLpVDuraCnZ7aa09hv3gxHYFR5NaP
MAsE44Cd1aR8hTzDwIVKoGtbRxwPqFzcaeyp9oCdL69QyKbqBceWkHW8Pmx/rgkEqAxShjCNmK8V
w7kHi2TXNXOYEEYf3iEdnofpVfp4ic1caFIRLDuDWxaQd6zo6C3oRnYHXlXLXD6ApnGazObNafU/
ZXNuFJNyeY+1TlreZUUwtJFVL7oIdgE6cLnieJnhckqtEk5Ibm6W/kxhpQuya6WPwb/soO/20ufR
th7DUH4PCPjcJWyXQ2x40DPVjJ4lvwGjqA4GZi0vDZkgZ8s/JNkxqQYzpbmHi6XM0rElHeC+7poO
xTjN1tUvnjPKbmYomndXeoQ32adQL0shvTyfnPo41CCtiquaFYjfk75UiGvyXOj9w3idoNOhkIMu
j/RHVZ+I1gmikvcbFIDRxIu3B/exxUDdCb6iP8G7nejuqS+Tvx92c/IUxiVaZ6mzehcMdpobLLce
w6MWIFMCR4p+JTC95AoWWxhGJLBbNVT/4jUs3ejiEP0JyINQ2M0IcHSWVvnIX/NzxsFOHW7QnbHN
Pca9fmjPtCE2ROSZym1wg3sUaXMf8HLMlVCg14rkJuf8d14ZbcA7rsrPNm0X924r3IkDDSp2CzU5
C3ueVLh8gWP5mkFZsBseKyLXmIYA1g5hIK2O4Ww4MH7XnphChpSMpOPyRUM+3kfSTiPMbNAryyA5
PPEm5Qw2OPOAwOrxRxuWFFbETTOJf30gEmtnpP5RmR3l88Gd+0sTWTV08+nG5qem/ZqyiTG9DDTc
Q+EczQAK49t6rJi1XSPDxowfst+ViBgYWaR47uasyN/qmSOSXJ2a8xn4d1CR9vlYjKdZtxCPOyBw
HrJ1UdesAIWyvqSThOGWa0ABgT1vmZOT2zCg0DTvKIvvsH00YGraEfUr8lVwL0V8exvxFqZC8d1a
aFiEE7e8XKWmgDJEZ7Fv9aPoaRnYOhVls8S96X8VBvbX85ca9GYwX4L2GOmdOnUeCSiQdZpY5JkU
AKUi2zG/F12FZnEBLwVe8TkQHhuPtO/uP2IwY4/5W5yiFbvY0NlGPYfHFxZBiwhIVfL4VR2u2+gq
Cxar926pU32spNlPETSJz7/LzvkgM8gc5n//G0V9xI+LNG5cj+B8iVNtxg8fYqnY7GEnofZXK8cj
UkTCNH0Fsmr2eYT8zYRvIjEka+Q+gPaxn7FOR72XwiFh2A4QJUfi36EP3h9sRHpn0hpia06Vi0yS
wJkqvod0zxfWb6TyKn0o1/e00GuopPTvmtI8vMQ9SKnYYxfWBTkMZhG2qarcchMkX+gZ+ghLDld/
qgSX5x7kCmqK/zXa2xpQ3tc0xk/3i9KRhNS9M58X9OsZAcMVA1NdrgFjR7q2YqTZsOxEswd8oP+o
/ouIxW/0SDRQ4bIInMHQOkLY20L80Blu8Z2PCe/nahZ2/gcVyVZn9QEiv3ziSpqH1F6X/etLohCq
CM3BykreywmcZoTPvatZfxaU0TzADNKO/fyb88KhjpB4kunjL1ml3zcQtOpzeyqWG6bzRnnN4YYl
DUXvUT097FWsNFBNQla/5w8DRs6TYaA8xBEtCpkjnKc/uuxeiagITtQSfxrD1617j52h4XOic16Y
OAlK8/NGCcyEAcmoYopxf9F9+D81MjcW/E+dQWM2trSAoeuTzFytQE4mNu8yrzXe0g4ZGwZeOYAn
4nCRs3dsstWlTEifNuzCHexBI1bsltWADLlsB9S+ydor/P2O4pKV5kAExS+JSxmVdUoDkBgkP+tY
DTPpNcg+HClLsEwOBz6urLUzpr24DJPR/AaUnEbHtQF9NYXzHDaPsio90886Pe3M03vnToS/zpJD
1ZCRRlpgjXuLJB2NmuawVZD4X+6LlOezLLKCmDqGyB5ybKWSjBqimoyCB03//KbA+Td5sQ6pZ1M+
gl9Rn6RFjRp3xgcbe9BLMicQ8GSsdN8bNIvSmndth2r+rfT0hS8sMx+6T5EWM1veH+4fILCroT4S
taxU5A/6tKVJcNTx5+lD+Fs+mAeMnZA9AoZJ/f79MrS021yzXPuAq5ccV3draMMS8OUeqMEVjSxx
GxlKZj/PCOkIAqGueR7zto4gfVSXIrj3FfgJSobOy18pjOGVSWJ7diW8qzyNRC9QxUalvYbe73G+
baQV1eSSMANoqzcYsfgoxr8NkHyhQF5wE9O9q2vT/+VCr0BCQwroZkhywYRRjoQnpxBWlCXQV6SY
EvIz70nHbY5m80tfQty+PPMCeMwdHBt5o09g0aBY6bqARlXG8aHnQpUjQjBE6oJ9LgHAM+nG0caq
vy8BBf+vewIsSaCxxNAdyP40447SLrbKNCjpttEiVaowP93FMrmBA4kIz40Wn5dhy00HoEr4FV+L
A+fQb0OPEM7p/Fgkxlp5IAJvpFrPleM5iKNe2DP4TypzbFioujTvGC9HoKnmKE3Vz7qrShZufszr
374GPC7nmq8T/8KYzfmNkHwHCapcdU8MtWSEijDEFg1KdIipRjOW4QmXeB+K4i9vnCTOKSsL71qO
gEZ9axcxmRu9r4iNJx9kkSit0YGzCFSOTczzj3YWRZ55o7LSv2Aoy2JbRFj6evNDVbICJ9IKbA/B
l+Ble/TrhEsAQM22vHJsSB5guWaTSzqvHgR+XYFK6NFEWIdn03vgAxoZTHe/7mSY+eU8Otq85K9n
4x9vOdD7hXDiTrPMSfa2urbC+mel6wFzrSER6a+ltcWsb8hDHpQn208h4snUrqIobEAuc7y+ua8d
onfr53CES/3bQL5Nv+c74Imfl7J0FQiQznsnwUSmwhHRuJEz7/wkbKh6iqkGaBFa+tPQLNaYx2UP
dUcURhrFFAQoovep7qJyaQtTKgUwnHO5mPH5MloTZkD+ERe+kVv6ThwpjKcdVwFJHFlRd9UmFzor
sBSYzlrCWIT85dBxiU6xmrJSPlO/xGRq85rFPCxQ37jqw7WC9ShI6ZC7c0DrNBc8nojBlauOIYMy
ligPsv+BDPOKIsNBq50B/8u9LjdjqdLr7uPrTxt98MaZZ8JH0IF9JpyAtiv2VA0SQBeNtGT5FIx2
SY/8hPyqRFAu2HBbXhD9ba87UQYnsdzuKt3RzYAoiFusM94gjAYRAu17NDiabkwAGywaLGr9hmpZ
/OlZxkqQFm3f3M/b4Y+C70a8+C2BTSgiOWE0ydeyOaaK9i5mvfuvBO9D6+NwxH9VT4N3I4HgmKxV
IOU4pWVADSFbDJO127Fv6Ssw0U69UnEdhsKhG4QSby/9wnk0NYMaeEhvltKsy9Tq8zK18mvFoPVT
DEa8phIZtDEncrD98BMcjh7W5oUL4mO19u5j6VkTQBXpwcI9vfi9Ip8gllCZDF6DY9ypbdYDzL32
l1FKybZmfr+uShiTDNcctgbvOAJfkBvJkKDbAOvC0hGCFNGi8usE2kfhfikPd5IzzRlfFuDZ+6fv
vb6u6vyl9VtiRT9eJXqRph70EPaplzWAUKObxJeBKtL6pVKlZ+wWnSJqCx1IsAtubpw0G2LIRqWw
l+pw67Vqqk0U97mgm2zul9BTqmdWzKOz7FhF/Lwn5fwU4TgoOUYVDj2WVpNTxNFU4YN4/FzN65+J
Ap/K/T8RALVmoq6kZ4GYj2kWQfTBk34zkDfLr7K8LeVQVG/uNIRswTUEI/DeYrznQCFEZ+btL5qb
lNLeXhHCCWTBXw1WPeJCg5QHXlezxCJcBbc4qZxt1vVgT7vUFz8UM8lvLIAgMx5BFBR2lI9IytwD
N+dx7i5aGJ686yTES9YOOI5wZLbXPEwzF8FjiCvlxEyEtUGxZGfd8/1aoGHZoubolo+f+mUBPVDw
WZ2Qyd1e8/SbayRggNdyF4ektsflD0sxIjnrmws5UPa5HJ/ranZBc2QUexYKQiijXsrMqNKbFtAq
H6wakNDAydHxk4f+E2x3PiuudU5a9Y0AIyCq4tSvFSpTndPDYr4QWkY7+Oy9zVGeIiUqth4VGMaB
52YA7fx4sl+HFFfinOW+p8K3PeTvdNSnykzBrdPt00n8i5W3y0u/46122S7VCRW8mZj71bE1AiH3
oySlf+yWFSjR466KtBzAl6wLhaHkLwm2D7oyHTOaJYNg4bsQzbQ4euJomM4WE/9uOPdhTG1VJFYX
ifLzNEYWfMaFHkTYx1bbEyqY4qFgkBLHOJILn+lRTD6i+1wV7kjAj7SlhbBz3jB0zYOd3HUO3FbT
vriPWedNJ0ht0TbQXS2I6EbEWY0h9cds0pTrbrE3Gqj3UjyuobJFvzuDuGnR4h/YaYmdNjHZsqf3
eA77v9/hw3VFm+mAOaln2oj6PYITk5/EboijCg7I6RYZe3hREMo3WXmxKiHl0srhCVv20l+lqJXI
8ByfQ53X9Hw+YD8lkbN5ZKi5gTQsrytvzhVSQTW1yeUOQF0GgQoQCFBtdS+IAfsgsIbPkzRKGlUL
jsUvONApiZCr1hGBzm7Jcm/1eYWGRv5mdmzO+HKBEIiSXwXCS8257HGwS4Dku9q+Bou40LAYEo5U
zhbvRExRpGaRwwyn5wG8wktjfymPoNqacH5C+OuvQjgYQIKu2NkMOzhQxKqww7oQUpSYQdl8ndwK
zlZ9mK3eikWQ1fWz4JdhA6pON/R76BmWp9M67avkZu4RO1KVs20dIy8CqAqDn0h4oQLljXllTi1W
4QUQdmMIyrNv6xBT/P/GWUJPVeJy6Ddf4NoaYM10pQfJobItnN5ZhoS2Eka6vnWfVtFJXx8l07Rk
cMxMFL9vNrPskhowLwYDXAEpveJGgrRdZ6XZVKTOaHCDkxQeRo7OYqAlsQhKLtxSUpClg2xPJZzy
sIykNsEwVAgtP+EfALG0Xp9Wub2zPrbucTwQuwT5q97Z78UFrSlrv+zLOf2ORAjOun+4OFU/zPcl
55YpktggND/K0JI5Chj5OrAkkdbiSXiT0q9sJdsSAjHhg6jtzzNCyw5KjwSvx1g9vgNlXBGx4e8M
Gz7h4TAr4pZTtkT6iKwehTd80aUjKDNA/mqqzOWm7laI9k2eOcRTiW6RZFqqImTzJkp7qcI8/0s5
TNBc3VmwvHbpWGqVuIkzfttkYXSN/Dz9iVcoF8QiOkwtGByMzqGxmrSLC1q5wPxOnv2GXIhlAi0v
8ACjtQTU76OWolm7sVtkB16hdF7ALqmJ1n7KfDpb4PiEI7bTkatU/PhchwmGgWKkWWOb7uV2aYdY
fwbvdRAbAVdaztnQihVb/XA2XiVjc+m2+4VIe9m/QpvFF+dc80zwRuPHDlo9fxh+I5e6Lfu8iSOD
7hNoMGH80bIG40WPTrViIt9LfCbypOny3/Rda/q0usJCWVng76Mo2y7zis1WzbOToAf7+NI3vpBS
+cmHwj1waxUnnfkE9IlTBsReK0YThxHRP4eMyyE1lvDmyAWFa46NOjXeeZIZ+S+0nKfi55HwPuzq
OjLY/e2xrOsKPNsdDMGz2z7WGrqh1UOUW2z6Zv5agWPySV1I3IOQTfTJFmMgDa+BdfQpLLHzrhKT
qVG/mZOV2BvJYH10AtfRHotzjucTcmlBFJm2nZ2Y9Mb3Y9zUmKfiOMLSCpX+c+PcpTtdATGGbCA2
MvvANBkwTMaRU94BHsn4t3+8YqceLZHAYBHf751jn+Omp4+EnawoGFJ6RLh2pKkimcU5g7lrqM15
UAW5xVqTZELSyb56pROxMwa47Uq1IWswxQONf49eolFQQ2R6pHWlv0hwzdTl5o97se4veXqySiUa
4j7w065IzjsycINlnwpcB1pWOpUimTEPBWqlr+1tMcBfToBN34wlCPHAtbTaNL8XSYwxVW81HJlk
4Ucc38YZouaagLdUO82z8EaiMqQhk1F05Dkeh7CGPhTSvko64/fJU2mDZTZjEIgOw9Vtp35tMdCj
lYz3fRJxKSGmMb3O/vH3Bz0ow5D/Yp7fji69G+OYUIniE34igX9Ywh/7xvZTvl4kjXHS5vfwf2bx
uR4OWQaZ2EKVbqwVXTV24TNXv6QWczOWQJ7ltZWJMcDz93BVun9OGDuW+FGu2QbNXKxdtoFF6IJ0
BVy+zrSduNDaRSh8x1fm2KtyS1bvpjSYFpNbxmWq4zSaVKGcvhCnBZIyJqfc/VbJyXUb34/ALEO2
3ym73ChpNG0biNvsW2Y/5D4YxgTb9k1a7xidUC6Ifwrtpcy0ck6e69LXdl1Tgx+CwPrSi7tjWG81
WdEdA/DWbB6wmn0i8x516fvkT2IthPzYdUwmurrfULC9zn7e+gRSczhdAxcyWHEgiHuJZSwL+Uwg
hOmEff5m5TYxKXAOyuj1SjJqgSfERYpb5x/bjF61+MgO1Q5zLc6puXjBI6n3JiUKqVUtyvq4/PbA
5o6UjTMCJ6Hv+FDTk6prbXrciJqpO1drVF072kq1Ht0lPfi1yZwPAeYLo9jN0LDqQUsk63qT3CIv
sVbLvt+K0NvDa1kotLbTgl3wvyhosUaOIRyMtql5iN81+Bh37GLLExrpkb2MOeZMhgvVvQZpS8zi
2D89NH+r8JVVL0QLr1mfbfseyloAvfiBwiDLR3FqeWWfLN0Ru2WuRxIQaCwDsZ+rpTsTsX7hfC44
KUFso1u64wI+qfAsJw2KwYKRV9XiJG2kbGGEGOkJes934B+OH+y6Fys7XvRB63TPPv4+CB2Ss2c1
ZGCtkABS8pQiwnN7GOvKfQgfs/cNul306BjgmIdzO1evCCJ7V6kZq4n8sxnmu6QObtbWHzSrVMdw
wMDfGeN6h3NOMdRTIjIMzbydYvGuvZnmLRZite06zs5sWPbcSJ3K2wADI4WQcAuwFXwQDWBoCUw9
C8T+9w8FApY93VgiVk3hFiU2vmfeiYxHjGJHd39OTwCUtqPxJfDNGZfrcg7bb2r2qx+xoprG2lN/
JKZVdcdfpR9T9Laci/yJEfJUk6RshmWLPVPuFw2VVrCjc04LHMxhU80O7WWs6mQ7qRTmVrHXpYto
SI10seX+zWhwGyXnEI1I81eRJp+vd3FTD+I0OTFlDWvLz+8jU6Xg1dOP4V+fi7Gn8MW5PloH8Fal
VecStJFDWMht6ZjbqDSXOEcpluf7Ylwetab5tfLs3x4nerDuW4szN+RLukwaDaDDAme1Vj83g1pt
F9SBlBcKvLpaqZQ7vQ9XYv2ZXXn/jNHLjWLvvqziaR6vKj1F2DcnU5AYU4yG3oQ/dsuoRPQeFFMn
Wt+2oCxA+kJemuLmZq7x/NrXsI0luiRtSgifaR2a50X7MTuea1tQFSFwejLPMrqz68mn5LF0oHuh
ffEWiNvzs+KUD5UcJwiZe4EAlFwD/xyMzoewl5D8top/A9KRT/cjhhkAY5LRDoneWRuPskE9Wqdy
wsN2e8cOxu5gTRxpwZC1K3aN5es8pU0401aeOpaTo5m/3FfTYoCl8mqET5kARhkxaB8z5U9hgO+d
+zsyWSTLKNUp9KqY7nFCJq3PaPbb+8gVPj7Rwk5/I0JaObZLxFpSfKwnfbizJHLtmYPG8UUdvBuX
YeMsX1LDG0xaYQuJaiL8OM3ljOrUHRCYgTRoXYQ8/zfDnCcHsJKhRM8zkXzvvMLhrEsYpIwOzLYv
pAL0S+kc8y6p0i0TzcGNIFk3h9RXhOkRVx/mXSOUq0MsaMBGhePAoJxIM8Iqe4K64S8MvVbMmR6m
ED1SO/alHoJOJVgMrxjL0Jfp3m6waKLabWFmU9N7bzC5x8HglyU8q/+UhzGNY3jMq+yTYoJBPUgP
Jux5PpGYC4W7HioqmhE6Op3oIfSBgUv+kko2WXbX6z9jiYGyDkzgWpF6ccQ9xS7OXeejfqeWeRZs
X8xHVb1qRINOkhyeiPofXEehFuCASBonvhb/cKAzLtgqlrZZ8CN9+/6ABRfZeJIuD2tQU6onwmwB
5xY/a0shfkw2TrFekKHp7Gms3QV5iItfjxrP1EMDLd8EizjGDH+is1TSIBjWQdve7mfbBEXG//QE
Pyk8Gcczn/Fw8bN+zjaJoQKMMZTyvoWL/25c8+oIZ0o55MQS9wy44oS2zNsLgvIqSfurDvjlrPbe
NoiqI+IrNO+wEgp/y8iktJTB2TPBzTvmoh95PDqmwyL4jxWHwrtLradi+X/CiksJDyRtOAv/nO96
ztADOCMRoqx/UAQmwB+OuDCRX8mYAhwQcxsPMMUh5C2PMf8CkMwSwxlRkElDmZPKe7kEKnLVP2ER
ErRqXRDgHGon4ZGEibM6O9aVsr5hI5rcuNjAaj0+XpSAw4GrGycA24SzPYlbJ/eqiyKkvzvLaTHD
Us+bBSy3RB5PIbWxaXZNbOP5SPTl+Ztea/pU0BfC9fb36jDMeWxiCW0OMeT+rRXqVJJfgVwm1etV
QpY7lcQEbMisV48pjwyVzx8iHEfU+OUTU9zbYqZrqVzkfJYBcsFEMVSyw2pASuUjpU0P9+4uBos3
3zoI0PekRYhEW1u+WC42Wvt/MYccnTCadPbFTXZLl9G0pm2JRH8UCNA5EUzkzn5v4oG3PTtgdMwo
/uQJTaOVLWV1T0hU9wlRjG/2aH8myWI2Q9MqZJYygPbQo7y8YKA/K/kaBRO6fQEO2AEuFHCCnIuO
jRiV3HNmntcaYxQ5gIzLXZpvfaDyKSy+M71LveMV6kosOGoBZ1Mq+L7Fsg0NS9ZAZoBW5tUEAHqP
XRXkhrBh7o90XabG20RiSJO9wM2ZSJ3rKebIdlRrSgHSB5fMOqXlTwH+UHy9Vx7nI9cL2dZW6F9E
aS/yne1rZw18QQ8YVpnVNXMCzJdJCzq/hWZ4KhkRCL2ZjEouiAlc4pmJnOjoRz/OczOWL8N/bpCI
GXKmjYaTIAMqEPrOaMrGadLzBe92VnKweZWpKD5QVNVoCOJ/nXb1225xjGGU5FhLAsAYzpEdwPbz
i4SUNkhJa9UGi04EIVz5H+mzNpmLGffoyA0LtsfQHY71XoYN8LqqUBj0kRJ6Gtczhok5nTqBFC8w
f5hD8xryVUsuFyBrZPxPCUbRawLrexs/pW/onH8e1hBAjhj/jb2ZixAL1BDIPc+7cujWBJ97D15M
LFzCQfBS5xX9KfLPuyBCvBtJxw70nu72x0uuF/q+jkeuO5gtjlXoH7KDznNg9hHQDe2EDSgyIUSA
YY41TaeEDnqBtXnu91lLFKL4xjliJR1gI+mM2MJ2DR7/P3ozjiwOOaarHv+fANln942vbu5YIdID
MFx0wfc3Tg901X83o9CmKHNbdPE6m1XiwkNOy81Fn/tlYgSa3E6drDxc/mohOuitnPuOWJgAGaCI
dkUeeOfABtN8mT/NXZ5brUREy106gWVZ2lU0je4PvESvy1PyKNVmzg56aKh7MBgabvZBqW7yxSlI
SQHmqcSvMRfOzCiNCHeMGpk1KL0sCcquL/pNg9CK+mdcCtqFnXGq/KpYOEuYNnoSsxrJxcEHMaHs
a9elw1MYc3YQgi+J+DIGow1rWn+3ieXi6O39o3VvEh4mqj07Sr76pfjX96+AucqfKPuzAT4q4rwl
GXSL2NfsgOZ7xxzlgINI37wjMzG70WogoKsDZyLtWJAiyAafLGLNDskM3tpFs52K6yCpNCoTw3+N
pwGfA0pAHUzJCS7FoMHxuRdyxrmsDLE5o5CegCoyNUcIZM/zUOq8Y8s0Y+Udh/swILBwf7Sw8Cxt
SwST6eCz7dJDslE1WW1GYhb4iU+GjQRRIUPqBFqCb52D+wAilziMuhmxdio8ev6EyQIdmhyMzlZd
HMY56hINTbZ1FE2Cs/w47+pg122Fz0z0FZJrxk5Oz+yTKZOT2dOFmFl33Q2+1zy6c1rgpFNN+478
jMTmJtkR45dWavSreof0YmOjRZCupNcA8o5ZFFKtK9GvRB6c4A4OPSPcnbr697WbLvPALb4LANGA
nI3V4FnZf4hCn2pU+Gd0ZwykmqCRASBsHqxUtBJzxyGXM2EEdLFPZkS8GW1Ebw44K7lvY2Xu69Vq
Bm0L1z172wlt//QMcsaA9S31xxRknsrS567vX/W6cmOkdWT7HoQooN3bcukYMIJeMrXMMOoxJ2HT
UpAZ93gvk6UR4DLQ7c7IhOkQ+qg4BASoInE2VbWbOtXMmi8WvYXR3PGiUftavux8eDICOwGrsLPK
Z0zlkjJKytH216em9U3crwQon7LJH7V7U1w4mazPbaABnUmSDU8bj8YowJDp5zBlVjzdKRCoWdOF
+8Ai7DH7bf8j4+br5D8yYZ34iwwhBH/B1ytQeWFdaOgOOwynpqdrHNr3kjDxpK2G0Sb6JynhDzWp
CnEBSt79oWORwbszLqAWRSdzqCqcwXw6HY/8Y71r/EAColCofhyZt98/mXHeXoqj4BT/cI427uJH
cnfyJQpdGjFgG7vkJ1e4xwpGnqtF9w8xZsW5r51H4Pr2PbY0j1ZFyqRZPHGVzpCJAy6/fPLEtiGF
8mPeQoiheY/gnM4gYfMvnuN/VPkQgak3xkzoOuNzGUSjsnVXCwsJiQhRAiwph7AC4i90y3If/mxg
MwrQp8HQBDEUSOPEOP4L/gEfoVMHtTT3Q4XCQ2wXv8MJ1yPvhLAQmjTRUtkX0hectDp9/x7XGFHq
U7we6gSaqO8786LK7c8cTu/A3qlYHclEv1WvQ581KJ/vI2/H6ZWkcGWNxOjDas+i2Q2KdviII/Eo
z5A/JT/tPIAxNoSmRm5H2jolsgHNOmPVs4PUw5em6b0VtBmGfo+K+oR6F+mB2ZcPZT4aqpBKgKZe
sjlsr76wPcfcDt2A2hLN/KFHE1QTCYyUWZdrpf4v2lJ6Y56mVw5NbiVVYipn0ujYvjURg/CuXGe9
HfCv3fAzN7g9saZAnuAl2qHMyDBZiyyZjOvUVXCPccvnF8sC4Ci7SAybli4uFH+xkXxZ/lenq+ui
Mx7OxUOd5DPT1XFObOwcDLbGFBvtODukcLE9SMQ3zoFU3cBckLGEBSOlXK6Kv1BbPyHI+QlPMHHZ
k2wjclrDJvJWhb/BDYSa/NYASgsCWo73gfcCR0kz94N4kP062cPb9qmS0KnoDEe44BZHO0MOB/Ca
mKkdg4TdcvykbNrRvVsdg6BseW4uCuI9lYt5FcprHnbfsuA57MaNNXAD8t/UKdlA8XVZFaCTZ1+N
tHKbVwQk9gxMsQGM4whnKs+zNh5c6a7rmIoB7YB59peArZHML1a9M34TohbQn188g2mQnzWkZPEc
oh/Hp5yvHPb8h9XgwoQcziqWScHmnqgJpKvfRj2kdxAl/RJh2OHB+tQ5ZJEJkkH46q0nCXbM7w3T
TzSzb6Kou+SsXje8ofp1paMhaE7HIZO5nITcn0kaSuPY1rNOdH9Ed7BvGQN7lIt5NG+eWzsLuZlS
qY1PyfUuUykRQbZEE47m1dBJcP836unEhZEjE4lE1FVmV39M5VWIwcgnIPPCrBPokoLcrVFCEv5Y
C2F0LcXqsaTtPfaw44uvXXic84InweN7s8P70I/cEUt0YRn7ggX97zeayH4I5VZWtKWpdguohDfE
fj6nwI/jswaLQX0s0TzAEwVd5hyp15kD9HtbpMuREbiflXf3cHvnBstbZ80gUYHtjgma6EiD8BN2
ISX95QmpsPCOXKIFJG6p4ACRE3daVw7a/KfJLV+aJf3X+71sMlYKztd+ZTx8oZ+NzqLQFs3uHu7O
AoOV0yC1cSr9LZZ6onSr6/C7nD5BN5Es1T8QfQkmO1cStlmSCma6pPjPkTx/6uEMq1mGd5++dSKI
GdMwslQRId5GpWM9OvGuGn2xxN2NGCIS3MroplD98ZpH/0mPmXFhsB/Zc2S7Ki27I113i3HalaUZ
OZpjAPAr84mB0qfOMZ8VOUNNMGCBOpTeKIJymNtNwKVDRWC5c1tOZymrGcQJ313KzMpt1f4i/cCP
6WLxNSpBPk/cdxhTZs9jt86oakd0Qr18md2TSfrIG7HIP8JBbmNDHPwvR6ZJh3mHk9Vf6q6KdpRh
rRHeu0kP8jBx2s4azrQmlBpg9Ajw5ZiLwOQcdm9qTEazVWZQMrfbhklyg1gd0pyUbSrtGKRDxGvu
dR9QWocC3l4ZKG3yvZDMygMWro92t+1iyAsG4OG78B8FJLw5oO37HhBxDUgzeSqylquRHrfoJ3qn
BWNbR5XZO8b6ZPO2owMfCCThVsDZiMsYFirm1iBHd1Vr2BVjjfOZyFhiWTDeKDbaox5Ksxa929Lw
PVafJlC+hMypnD3LbrUY4o2GZ97Dmblm0PWH9XYaINxJnPQHnNYiQ2dTyQi9LIYrcXBIpEnHthDF
Aj82PK7tMQrzpVE18fbry0R/f32AOxCQ2pOXYeQ8sxqt/SHbdJdWTCcqgp7gF6ZBsck340D1s4bg
/OrGdRi2SrHP+vNcOYHhGPpbeB5eYReHJGA5yw7BfnRQmHszm69pH9xZZdPmNNLRU20/TtnYi+PL
5k4FEKJna0bpylsIh+VG1PSKy/+/+7DZrrCm9hPDEcXyq9Zd/OH9vGFGpCCRwNc31lnFgWOtsLNk
VyVYnF3b2G7/4G3dOBjO9fTc9TbHiu6eYz3xR85iZdyonxZVVBJ3wvxhHzSOUKgKcGf+TaKLtzNK
t3Fkd5dHFLPTMYq39MBcX3Eilmvz5y7uXB1p0GrQgxfOcVG9+/uzyGg4cT3vSSP+vpUwKjyQEUCb
aNGcopFQKiqz86wnXXGDMlfb4+OsWq9TirvSoZaMJIg5tVRBAugNFHLr4SN0iT8gM8Q4+2FuGP0z
8FRog6gP1y883UQf02mjJgEnnUuoYcJkVwsMk36AOzCrZ9Q/OkdvaY0hRSmB35qhSEB+RLDGldym
vpo3v99LkS+KRSbhoFd6V9SxIALc82ka11TMpEGXyHyU9ivJHm4At6Rq3OfGpfC5GMUAeO3v1+hT
DLEnlYhyRSSYT5hL8YS4OcvyqDdCa7SV8wlj3DvCosaaYAIwPUYwmnfHGilav9YDb4xILuIzqAy5
iUYhPlu+0sqnAevebiucKpUXExGseYSznhrBN8VmtGcoYHeieUvNdVUp8PX7kgLweLT3Cbs8ETgB
Cv9c45brZUA+2QKfSijNQ/sTG3Kt8l3AkKiZBLncqgO9dPwwuxC3UroprKzHVhxVrVccd8K4QYq4
E8KkmxtIoCqb/txGqSjpTtIij1tXvtZeAHx9ZO0eNyF4fA7cXqaJMczJn57ljhj9f5bpqbd5fS+g
P63c+ZLtqXhFPeewN75e85Q8II+ZElBf+NT60xYp7LdFCC3EPC/LOEPn43DEJoEUadARI3z8iCyW
XAfRaD8dvg2FPAYxEfey6t7QnuK5Cf8RdnwrEJ7mN98JYMvdXrmY8++Cza6g4uGTjxCNboQ+tEBf
FXLUW2DHPAO5X3RzU3LXk+UoCA6f0F5skkCo48ThjFHDae0fou28hHPfn5YQj+8IZbOZenfSyh2U
8bRpdzq3M7AVpdPZVxOqivs5l1rreOH53Zy5+TXSr3I76QgeHEqt+cl8U5oN5Jtpz+6acK/0tKqw
VXGiISWOWOKOqf1dGQogEdpXeg+iuzpht0FJ3Syb19OwoUMoK3ejFhJ17Kc4It/YXYJBiAduExq9
JZtlbv2x0ZkYObfxwwAPAXnrWTnysit0WrQf6nbjO6thhE/nvV9nereYMgywErMTVXve3Xa95Wak
fsnsQmkp7HXSAE12UitdRBT1YlzR9YTmwDe9Od/93ACe0RFlmgmYeSveEyD4gq2TH7HdZ6FKeGXu
t7Xm4ZQnsV5k4Mo0h6JEmsRbhbnjHcL8eoOymXQfQPqG41oNsX95+gRvED/68kHV86FQrBz8sI0q
aosuovBKJ7K6RFCgjQkvxlHCalyoFOotXs201OmBLu9LZP6CzA8+Dn+PZUwbDVC5COJb/dXXxYJ0
Y5Oc2eLCxJhdmR74gpMxW56JIW40wExHvYWiiOHqjqrNeRDXrGkYvljUIVMk72kigi+m1Hu38Lfi
Np7XhXWaRqWiaeCpMEBQk9w2G6IlYUFaXasU7Q6p/DbU5hbO1NnX6AFMfUSBFZECwM+SoC+AcnSJ
XtUbxDq9vNuHgJmWDCO40heTbS063VhhhOJb9/DpDxc21WQvxPmLc5aQ6dRjte8eUY+UhINq/juT
/AKVfzOf2n9fWCzZS5IWhqOxLJcORp5JHDh23m1yuYfhPzPbWIHxQkdlMSQtoNvMxpVTNP8BEHEm
y7j3w9yaayl1gAL6LjbnpHe49gUfs0G+ic+Gn/RAQGkyaVxK4zPyOQx+3uuuJDRvyBkN6k/bknBu
u+3oncodX21mJJVICWUMpkvsZEoh1NdUNiR6ZdUKTItMCgOH8IbGcyAJAozCgzNvRwbKWbL1DOtC
s+2eHs1LyQ52ZNba2LpF0cYVW0GXCG0tKQLy7GnlFkpbyXvXosp2TMOT7kTTUGHGif5oerndhNeO
dCf0EUzo5rDogaDk6pcxi84FHczFIMKZzWPJQYwFGh1BunDRykndiyB1IQzSCr9z97Q2askdvLSo
1BJY97znNQbWrn52IlPbFZV38u2V7jG2XiBsLoiICJxmDVSoueGa17tK4XmEObRNoydnRZxbQ4hl
BobAxyGJWZMQhNMtpW0MKPQD3oDdSIHpxQd0zKtde6+5AXDTNZPlFnHetRN8HEUiTDXlg0zyPewV
iUXDZatm7FZRgiFzuS9+V5WwjkwBPutvYk75ge+jXgNZOixLRmDA0hmfl7/AhI1lis/xeefe4VPq
J8xpp1ZxXEuU56b++hFAquJZswgRFki9BIvO16Ohgpaeqm9bFbfIhOT6slO24upk4WJ1gSM+YzMS
LL4I3YS+YLhU/KLT1iL/vHUgU6oXZst4KPUuv0dtEacUdFsK0OGfZz8jh1V1ZoOdnfHiEQddX3AC
LRt1ABrt0uGMlie6kdITQv37vRb2UPYlh2MayN9lxAOns2Y8QaL62DQAyCM7lFXatdGx20oqge3b
tD/LRC3EFn/s7RzusiHTbs6Ogqu+IF0yEbhu1mqcJVt3mWThNB7QHL+26RIUDfdn5bAbo6TfwfwD
yHajrTkYgeKZQB7MdumILW0TqikwskjLK6JjjoyeP2PzkrWaQZnhlGYeVIfLfzz1oHmoyOi2gGqF
n+lGGSGCI84k+10uQ3Dxn8LsupPFetEgtbG74mtkPsmIZuTsQOqOCNuRpaU/Xz+kn8HcqGzwHrmM
/FKoICDO390Gb7+PMBTgXTTp5DfOhytHm8as3jVb5QoJM5qTO3CuafaXN7Y1uhbANoA7Eyi74KfD
0b8Tb8GZKpWVHP56r4OMxI51M4MPw8eZCetKr8dXw+mxSi8w2xPKmp0nBdVYynVJhZe9PJyl7zh/
A+X1SXlGjNQZUGFHmiTGrKWJvi4VoDqZ57rGJChOqPH+zxfHlFCaVlQZ/+FZ1D3rKpjNf4gIO0hE
JG1F5J2zOrkzNWKUwU46O5FvfCYreQt6w3HwnTTlXcKwTjL0Lx6kAY84Wcu1xCDa7GYizRSazoAo
yCe5zH6xeFSJAUDZbs9rh/MuR+Ok94oMSIFqVgudeJtw5IhdRCi1S4gaUmxEJRNrSYsXal+p/3LR
mUPxfKFDqmiBPig/yebXgHVsPbKtnGBInJWJyWZ9K/hxm9h7wPtHMG7Zrhlsp/soq7JCBS8/nrRy
SpqVDDK9W/+Cvzxx2iawiT29qlfQJBMqvt3StaCURjciDjIgLfEi5RjQn67JNmXbEYpMIuAE5mHO
pWG7sLpbeVaP38Vb3iMi2wgA9kX75misgx93FXKI+3DxLzH4a6J9tbTagqbp4fBEBwYYqwpHoCyz
SAohL9g4iVq2s2NFb90JIlJH1i2hQQH+Rvr9Bf+YTuBWMU/oQSNdRjBU3mEzE6WMBH9fMPM2al4V
XCryx9rw0ynliV4kPJutKVEqZc8EcguKjrG16K9V1mpfmybfqviW0mHcbboQJhKHSqNLXKo+uogo
AO6ouFooPhhqBm+TkXo+Ye5o0KMBf0BfGnlQz/if9gq139r5RQ51iFC71/MSVSDF0DKzG7qm4WMr
P5q2JEdZa8b8QRi+ymyyPyQUTvDiqCBohstxdFExCjTIyZGWAwqVE6l/QlHhtYYxVt+9KjQ86CAt
cndUkt46QiryBpwgFNvuRyQ4pK7Qh5kvJ4tBD0UDofU2ufoK6kKyaa7lTDtbQJkkGnTtdn56BEoY
AQGTndGbjuxtv5f95T0D9EAj5zX3zFrjHEEAl2418pWnBOr+ZNVscWs1rSS+5hJc29Dk4CyZtOqu
44RlrsheeHVHUrDW5wFKWfrXRm0wgIpIxljeUwiyoOt8sCGq8e0Ugyj1UqfJN8dAHeZQ7g39pqCz
nAgXKVYFyK69b+yk3IAVjJ1B5uCjdedTL2/ZNkjf2XANFK0x+dPwAnjaUNvsKedFUyxX+MEXKJZ8
89i+rei+qRrMGrotzsRYF0g4/a2mnDz3YKLAJxv1rL6YMnZXfzB9wDMrjlmEbgtvCDed/e4saAZ6
lfWZVuZrhYbCnzoBbWIolUeFhmLYd/Ascr1Cj37ww/c0ZKjCyc1rOydOXj+/0eEivtMOqI1DWn5y
jGVs9c5qoS4TFdSEvqY1KCbpmmy3LHn3KO00sCyiON7INmLQwe8HtblJrR+iWSNTpcuW7E8vrCkb
/ighmJife8sufxROAbMKhfz6zntvCzEuLtBUfzRqEsw1nMrYO1N+GbhgdNzu7MnbLceC0sVDTS6P
3cLL0sLHBxRL5U4Dc6Yt8tr4fi2os6hxhQrJOVbUQU7crXTrAyHGNZTUg6xjDG0Pycr8tWgSBPkz
jA0zjSXL2kmdhwKfQJapn+VOVblu7nTiqgq5iGJn4z0T6Mj/OX2KZY7sYAvN8OEFimKrOsgEnVuv
qHpnsXgUmC2AHVrlgOaT5dpjzt0sne7sND/4ReuItrwbPzt1TM2VJgeQDLi9h9wrJnpXm8sDbVnw
E1U8+47ye1YF3MgPb0MCreCZz2zFHnWKdzQ812aXyzxNwcJo5tnOxAZrNZzyPusYa/nbvcF5JHZY
61CNfTTtWBMmTJZ/N+6HWaYW3bC2YmUeM70L5Vd05E54l51NJpf8rF0CLFXz6L0ijmjV4k6r9g0Z
Vmzm9AcEMC+6MQ6629jMKglh9b0UKKRIXLgEcN/kdw+7z25xtzXGonHcMFZ2cLOjqQ4xzcbARwrW
/ujze8xMxk3pFjIK4Ws3Szq9OceJygtJBFPvvgtkO3MpQYO+r+wDllCejJk5zSXmjUtF5LIHV6lO
zAVd5tBnXxoSnhFo1Tfa1oqAqzVL8Sd/iVxLnI0vdKdzGnUFRnSKm5+ScD2JOrkrN1G2H7wJ6fK/
Mx8GsxggOf43OjSuFt4JgzWyHGdZWFX4/woPDcp8Uoe/pmpIqUrLgd1xIFa2DXyohja51iLjrRVy
2Ao234E9pv7A9EMbG9iK1QpBjZoySb2HKrYjLz17hrxHlVvzEtg+dZyQXgYYv4MJBBRSphvoBs+8
auPKU9EKWewsAS7Sv476qgkOj7HrWs2Ksf5dbMtk3z/hncoFlOzjNBV6OTA6nTuyRRUGjkSr0hAO
/nyRrCOhrNfr0c9I86RUxVfbpCHK2ldQLRtFVcX9+P5owWr4axBN/pcQacGa4znmYcvEuyBGocyW
fu9tWQYD2RR/aIwJjMkCMn0VkJLhE8sxmYj4m3ptpUiDVBBP4L8vaxKRCFwVJvMjzkgkX6C/Uuwe
qTehbbvWITGoJW0eBil/WlkQRIkgjUkcEt5xziH/j9Bqj58fNEycUuW+65KAg7YqNN2+Aq3dKXU3
GGYJ6txjIdU/DT7woG5j8wiyoB6MRR5AOoT7NkohXAIJTpVin8dI2f81b1VU27FeZWXm9ggXwDvG
L2E7wBGVXtJi1Dg3e1VN/AXr9hgwgFZnU2NI0R12cBebM32tm8mV6z6NzR+IV7zRr2IwbSP6CQXO
hc3NGg5UsPHvzu4WPUOdbv70fS0AixdOw/QvCe/caG/YyNlTPU3XbMqwZBFiUF9wxG9P4zNHx5yS
AHtEq3M92Ay0iHznmK4t3WS4old1WHHcmJRVi7qGOrxQwDGeLyrcCB0ZK2Yjq129xzTBqAhhDdJF
4P+v7m1zwos4sj6egyTWJuKCJ/2ssH5/RAYCcQnTxHO1E6wfFoAYQqTeiIeYOOUNcOBRcFCy/wE+
7Pm1UokRP8rcg1l/K8KmR1Rb6FlBSX8sSOd+8ALu9OaD2oUiIfKO2l2NffMknzlyCq4PAB3tYXLZ
rdXfw/yD1OCd4DtiPp61H64DEKRbpIi/f5cw4+lDC6fsTjyvi+7tYRshIl85e6sd7sMGXBV3ei3e
Hi0jeGYk0HGamJzZYoB8WqULcFTbVpznMj+cv0vGr4xtefgQDyE/Teogbr/Ufd3weDOin1uKJQeu
fcP+HuRdplj1KpQUJZZgCQq8Y8lZqw09UuEuS7yeUyo6fig9dz8fyQx2YH9YtClw6NDoOZRNRLAS
LJF4iwdkDV8YBRX+F9agL98UVNoNxRVeRloPE/NuAjMnPzxEkxtqrxeFYpdjRDxh3pRkUOoK7gb0
SDbvLAShOLdpLEPsTl23lGS6l3jMWoae01NPellw58w0cg+P994Rfw79JCAZtAroeWZoH0FLEqLB
C3t9jt2B6XVM+5xl+kPalbgfaL2OqjjxMdr+874JAGS7E2aX6QymWa2tmYPGLOVaUXmk5P6zww+b
PM5jYRHXZVMMWtedvDl1mWxPQT7IUmD9CsdPkWESvBh4VsoWIg9UNjOWXJgXmno7iUeQbt69HzGp
sjrNwh7FZZzcflMn64cz7PWiJlhDXlEqJN2xxFoPOGaGMz4uhnfn9WUjlzm/aXMOief2eMTwWds6
tC7VGUN5a1YANgj5G46Bj5L0eNBy27kE0p9s1ZYJpOXN5skXiPOEBq+0xDINb2Kg4zey8NqI9RIw
EK+5/fvzIIIL3AlAgSdYbnEaFlKCvI3CttRnvOsfd4VyaK+EsoZhb80/9fp4zFHUtf+fu+rFHjZh
R0zqyAGYXZKDuGjJt/yQ4z44oj6pV+LkRW9EoWzTMPX82Q+bPIDV1H2weXEZQHhxrYcSQhv65FSZ
XaemCmrOMxF+enC239xQA+ws96wS+mXHl7o7+V3lnvKcTtoak8uy+R2r/XgeZVQ9HZSKs+oIzTTV
CiJqvpdaoa2nHPYn4K40ViUNd0rF+vO+szpzOUBCu2aU4iYVSUxh9sPfwEkQA27PeC8Xb66lejOE
pD1XP7GjCkFycZxYNRr9aD5A9QAuYiXMUOZKqZoJsPb6UmUdHlKFDBeMKyGjTnfWYAtFrgYVy3U7
wVq+CRRPBBleDwnTSr/Y454qDMy+1nlwf3ZRfNhMw4GZ8gJrr4R5CHMdiUaeLT7/H0xX8MqKtEgx
cQaq1Zq/jYQdMUAfsC+MKDfsya77UUouVL6a9cpXbot3ZHxRHlCQGciaXmkuP+JkvS1MXPTD8a0W
MWVDWxUutbJYFZbbq4EsQVijUKFlnA+YANc7VRSrbkhTybqRs+HRCEGTUArjhZMjCGh+SdODYgNS
visGFdkisOGyj8/CjLJxFT3BxVFgM4IG7MBGOZXMwtl55J95obci7Rnp0bcoKVAVm3AHSyUEi6t9
RD3T4PANC8D9U/J8H9VcSEzMJLl84wsKax/4p+JqPBc64a+NgX1lE5XVRJ1I00oXmCqPO/KoHUi6
zsxl/LgOd/A4FRDi1Vf45AxoxY97l0hOmvvBoIb9spFoXDMAmUk/57mLP5EPgZPFfJAgdCzyyhDY
56nZ61NuD0+A+U30FOQiirr61NU8u1wIXKJgOQ4JVPOIKs9yC6jdlHLp5x/XouaQHJptEZpblW5b
WrO/pObBjIotl1VO03JJA85vMZabAH0EaS8aX8tiTbUJfaNOQgfD4F3HQNOY9ssFg3qiEHyJzEAz
+WuvLUStV8SweQEOG/SLmhkzIUjVueT9mfoaEEX8SRH3jbImHn80DgfRwrOJLFrB1W8wh0/3jBb6
72AGK5XLA3dMl1TdJTfe3QhFeZKMu5xGV2f9N8/INOVAFCJslCUPsYETb/ej0C5rwQmXWBK9EVIy
eKCmoKrZNU5STtIYet4/XkA/8H26jo6CsQYSyPOlqySG90c82v7dXil81Ieqsa5GsAeV7322+jCT
ohdfQ1ZjxRbq9IFM0bT5CQAENg8ElP+Q+cfJrLa9LWdpMyMtjq/OazaVXlHpaZZ8uhKEYhTfS9w4
JQ27jQ7njfd4KwZz0HOwfsbpIdbp9Q+Zg2R7OzSN0mN+Ywci7vPT9YujEbmMxsJru49e1AteQX/8
FJpnnm5OsNnxI37WNVxe8+KJKXN+k8lpAlFjOkuI9hWFEIdm+y5EvsDLf7S+qvEvw8VkMRLxF4D0
E9UxMf2ElcFG2R8C2o0ssvWHm0Nd3JGpw1vcjrnADXG1Vjkpzea/tdibEte8KbNXjbmUBICMsL9P
C+GpHWocQ/qDE1urYzTiDCmumgsB81jrqN04ICfmsjfiqEND+L+9ASr3B8Pw+3mDhMwGWgKTSYql
+z2UNWRU+XfFD2XihnNv3Zm2zu5d0cSrHS+UC2cu6m+20rpWs1fgymTUcijwIq/rnrPTjKzGqyCN
TwXt9a6vOnBa9HNI7y9dog8otKftGlfavhtJYI35KHxDam+FZC561KGNpQfzPD6WQVhAOvTh65+K
FffYOqRm6D9ySdbD51Br21L3xR0K0QYvYQMPwfyb5W22qVPjMcqlqhOS4aXPP8KboNgxMiL/RgTz
IQCn+uMKePI51Vc83cs2YdJHajETPmjv3pauKfqx5RLYT9tyikM41cpZn9cf6wQvJRYFwzs5jqAo
7sVAwUVpzXs2aA6lIbhW60/fuPrQe6gYxIy2LFH0CuWsq0+cYIk2Jd8pNWiSqt8CzXOEzQh56f1N
VT0Oh8+Sbqn84AJE5MiFc7taC+utAc+2znfQq6qlzinynJfHbrkBtbdlAt3Hmq8x0FXN9dlaeAw4
2JzFG8IC15MLHO7/5aJ214/3n3+wzNu+clAmxSMhEQ1MeEgLkIIBabCmTDBvPJjkLh7XjghJByXy
MRXHsjpyEpV3lZMUJeE7WFnh9ARI/UBDJ7xZjeRmPBlrdwP9f/5g/BqIEJW56WwcW6scoeOXVDKY
hsjJWtiTwcDoi3wFvEdyci4cwoAdcoXAt46fjPhuhRllWiRLGLJT3r7EtiACp2mXr76yfODfMGCT
69odyXpaF0xZ7d3ntgMUdBd8Dr1IIDfEHgtWkSJjPqW0YMPoZL4n/+Euy29bT7RrG7CsCYzqmZUh
Kg7LELL1tErMghmK0hHQJDl5IuqifBFqZr01Yw+B5ibr8lRoMsck8ST9HsVz4I+ZIMNHLk+KWJp9
r4G3uUEpbEs643PvO8Nl1OzM4cPiqtNg7voPhPe5c9d+A1aKF4cflD+Hr36q4uubyoTzAfwTCRqW
JoiGWiURQLIEZXKVEIYfQJLYavcY+3H0b55NMVwP1tAO3XhIymk/TzAujZLHGn5CMPdZn/Pm6LRR
1biuNL8DWR/E8BUD2VBxGwL3UOY3bQUPGF6MwBZ8P3mEB13c6qONSvqmTvplVGRewmE5h7Or0WIi
twy36AU1KTwJsAEfNsbf8q2+vU8oVnAhVqwT/GjdRpsHpAsz7VqHKXbGJ1XNFX1MHco+jwyABPCG
bBUPiFuvw0GPju74vIo3V9eBTapxi82Ax/PNeMwjVr+DuYa2/zq1g/MjW/yyn+ymkuilsdsYCgnt
1LsqaniHL/u/iQLCCXxjOHybfCPoG3JyBcxmQGZSxoOI0yvSSb8Ehd3DXsR0/Y7e0J50HHqape2Z
f63gu5UzQibK1T1mEj49VvjWzs+XD1eOUAJJE7o9gUVn1NIj/HMTHoKO4nPzaAgLVS/Q69h1Qr9V
HInujZOT3FYZtpOx/uHkjS3MBkphWwHb0n8CVre0fsRJhk6LLpk8sNOmr3UL93WXf8tXZjTovIB2
GpdHfLrRSXEei8GCHjGNl/sAwjThvJ1XL5rZ13SHwSDW28uc6aEmdlJWdgNvttJkhafkJGfsKCcE
pw1B2GqJVBTCH5jgIV3nrI/tqBV/ugzPVIzPapSkjuB3wdEb8g2EVmieR71vm9xVksAAgWMuBr0q
6kitFCjitzN2QZp0S1+lU2y7HqJOVHiDicaG0fjFabZRHU8X+c77r8OfDozvCPgZ6/IaJiKwzIJL
1Qd6/pTZkU4jk9+MVqUY+t1cxMjLsrk0gGIDPOgOs2dmpOh/+queV2oy2ctN7JZMOCIMjA+ECb58
DZtNEVHb0UlFGpMLX0o6c/qBFvzZ8X2RNWEY9OyelOacOkK2Ik8NPcpob62qqQZzf8h/d+OpqpXy
0Zg00OzR6ae3zzQSMfocm5AbW+jXsdRpv8djadd78TCGEGvor0vtvjC2hKcFyG5L3nMBeIzrzbkH
l/RM1OMEZe19FD16THeJGsBRwhAOY+gwwjop+rB3QDY8SrSjjgvEP1omJe6+/9cFvtLKlaPkvMzt
HM01FBZJWQZ9vrPNrY+eoyA8r7CDwZEzP/b/aOTY5MUhTFZhgl3Ae7q3QK7reJUOEH69kYu1NYhb
QTnzXFHXG67aTyM1S1XDMLf9HdyU5gkEdycB99qtc95Zf1kxKnEzf8o7E93lcusfR5MRx1HBF+la
49mBbDoFC+qoEnwfQ5kETN/cUsKloLXdr00mn+WbieJLFgYQR85uQ8AuhE0OW8diSrTeiCfvqMqT
agNwSN3QZyL7z4mpuzpjlVTZO9x0NA1EL2W44b4wwBauNV4y5VCd5lsy6C9Xaus2LtCfR+klyhAn
ERQaDcP2wuY5ttRIH2Ci2p99ypFPlx7kHRunliVlfQ8VYw2ocG2Hm4/swePXuZa6ScYWmmmneXow
avceK5TgWcLvxGIP14XH0kldBWAOqlMSFHFwOCDU92hj0z5U9y71iZmVI+3+b1Iq6vbcextI9aaz
K4z+tOaZJWFuHUAv8dTfFpe7YWMzqg9G6s2qqtcwQle+5la1dwsu5aw1nay8oeLzdn2KBOSDt4gZ
xeKrqTcheGCsceg5btAYr9xTA235k8vr9WrvrRNo/38p2jCso9TABl6OJrqxsZTQzelTlQsCW8Nr
Na0Lkul4djmP6i/w0iy/knbBRnbtBC+BBL+VzAUglZH5Arw/ClIbv9KsOhdWMvhSkjzihIMdcXff
VDq4D9cEXFlm/SQ/m3eKYjiJtShO3QSedLgWmQ+l+nOQDvsMG5CPVXlmwG1/pOF5CI9J9SdRbMW4
liWrm3OMJ4IA6HJfk0ZmjBAGSNaElo+HNim8IlQoVt8Hh41O/62rIj57puT+UBUZmUTWQMdv1Y6m
l15fXGleAx+6aSerHGXdJKb3L9ZaYPep/5pVxapRLWN39861i62gkkVhn0rT1G8dkmYsiEEDnBt+
ECGQZ6YqNZNgx3yaCelgMwIytiBDzwj3S6wjkASIxw9IM0I+H/PuN9QkTbU424Sw8fR/KiGbTw0z
Ns/9Tpjx7FabnpdXhOowLVzHMrtmp2pq3B36bVdqC8LJ38IOnL23agg0XIqLE/0q4a4qTJqcclyZ
d0+uTTVGa7bPqLLWckOAJOJGJK90+i6o8NpOKADCl3IwPiTeshTk7zb5b5DGb/4YPHwCg/2eUIzg
QSUJItDLmBUN7ASpcSlKDRaqYma0bML/G+2UBx7yO7+ooMfk3moUGWcQFxQyx0cEzXzIFNS6M6SK
iMhlMxNmoxnBgQQMZbYcsV6QRSYueQguiJIGdbImNcBEcVDhglAmbp44sIJU+db1TEYEfrUwAQNs
dSn7YgLd0eGNTt8xVvUIh3NGWkCIRymv7N7ySRUxgchlv5sBkDoXoLVvEo3riKaBtVugZiO97fQL
4+YyIJ6IhxNQ/za4J+R0bAyht1SFnSyCeUzw4OBGYWwidhzy2Qs7mXNVe0rjxKO5vBg9vbN2gbLU
mfnbFXACVawmmscsqh9H5Ad04HLWdTS9iQUN4hndfbTBw0Qu8/xNBtEnsgQSRfeMTPWBojHFwVoa
ASKSkA/8LQFld2Ne5iHsmGiQZGsLKQWk4aFN2DuCTf0g1AF71tlwfFDMINM4olNUgNbgZu8/ZdKF
Dx+j35HB1NwJPSwN49QpFOQusYT8qOClEf2wbQ/pAb2WDhnF9JKjthl3zGKd5uI9nLBzcCnQhtzr
p+vbI8yxN65bk5f22LL30f1u1E1yZ2ExA+8G0dUmYrL8AW37evwoO1BZK6UTWRm8syoroqbzh71M
3anEs2TwgAkNOrebXdie8nF7yWvFoKnm/P/0f/Tf4slSw3LZRAkBILUgz/lYbCtSHZMUXTPvFgHx
PzIwZu/zZKLHB6cKCvRyLYLIMCYo2bY2IOkGFLSd1pKxXjA2hB7dUKLVLujohe+Y0BlprcRT2+sJ
f1ibLKlYuD8TFJYva8OrIRKJEap7pt4OQ3sI5pLN4hIoB1uEJGocJcL26rTCbffzDsKzBKtO0Y6k
i/YZLj8MpRCp9pV6AI5nP8zA7Kqo3MXPjmb2J8inQeFTK06p2M3yqT2EjBHl9zJ1O5EpTXLhB/lD
uI6qetg56sEg/7IBCbSOS9ZzOTOgWMHlM1PN3wt3mPo+GsnWgw9YlAraQt81LMU3QThS3buOwoTf
WE78G8IR5A3cPzaRlNiQ0kEAkuIq19TDvZgswAoRfNyn3C+ypgfTIm4RV+V4OoSctG6seFJLC8tk
dQh03pNaj/5GvuKM2RL+Am8=
`pragma protect end_protected

// 
