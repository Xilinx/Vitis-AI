/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3296)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbGy58VxKRxo4zwlY3X+djIdjdLesuuKC9JTBqvbq8ducLSTYU6ivmbDy
9XK73CnYEwD//LD5HAr5ZfBaxIueXLag22W/kcdzn2gLbKyeWd+tbXTv143DJYST6X+2qNP7gILg
xjlLvgczV5Bg8chBZgJO27qVPaBDoLKpR+kRXmn+2pwzItBbc4Tvxlb+lYSeYfrdCvoS58oT/hpX
/dBa/x8BrYx3Pv/wm0C0Lq954TS0FU2Gd6JwbW/LTPRc7La4uLdXHUy5d3CajtHESKi3TMERmdsO
6Bw+zaaIJUizIR8yOk+PvoKyvfPfSKpoE9u/XvE88R9fUR7sf9/RYJ3h3zS4pQicSRtDD9GN0dTU
XADKFLXPqurhMVJFZaoCJ/wfK46aM0LGLOsdqVnayVoq+Z19vgXahMS7p7hyXqnepOf94wBt0mUG
2zKAmJMJTs1sEADV3E3du4XNP+KMoXSUB2CpS2HcPvLS77Q6K/zX4Kc1qGVKJijT0omhfmy/PvS6
GWZJdJEZ3XB6uwKArIwaR6QQ7WOytbIF8e4HOg2KnEmSrvM1AqrqFmT2N+4WMw/BiEVh0h+nUe91
ZP9Cpl7/mhusgBZfIzzclrGJGv0j9dOppCeecNTrp0xn1edS0M221WRNdYeWPSiLRCiY2BQspF//
TbINOxB0fyMgPFuErlaVMik2MiwRW460jINUpnuw4piAwvJALFl7z9FD3+osYzbx1OU2iqugEA1U
k3/WAvdDcoCJ/rMnOQYIIpzrsGSwTUTrWViAzdlLXskIP3VsG+1c73Z+knEW585jbA2nJvLmsDXP
g5eXQlApBzxPJcjQlZunRUk+I0wpHI8rJKjavt2c5yLBd+LDA7YkIQpThf1Ewmn4ki++l9fAT6J4
qvo47pIu6EMMHXQuc3QwxCMdj65hyCyyN/Sf0CJ2qSudXCVo4+zVT07hx44m3Hilux/tlsDXiPUE
o5UfRNme8DXHWnJ31pKPkFemqVNud3xz1nd6pFKChB9jyj7NzjlGzN2jABBUtay/ksVtghZ4Wpt3
8+OM6TSx9qZAhhQlGtHqM6Suq22EQEGAhG9XGEVnznAwXnCuzPOaUu9Vp4L0EZmhM4OGPp20Ztu1
bW6w0WBxbxI0v4NF7xVCYeZ0g5kdjpPAMewOqSCStUlN/ZE/aHNzPygLNdKZVhEoZfPu8f+9z7NX
WYenmB0oyZ0CUldyMKkWBs7k/ra4lGqo17xR18CShESchdXd2X/ozPpXO+28z4vD/a6S9seUaqCT
cTPnaXiBgNgf8+Go6uASe/kKiBt7WL3msBd4DTFrPDPRCCFN2ATtu6dWZQVv7CVyQJhgO+Wn/pb0
nfDTaTNxkhoaSX/4fnZKOq731UeBLKY1eG7iQ9WiNLhplrxzxjKCB1oyg9Fq5woNSIOLoqgE/YVm
6Q27WZy9NNzt5Nx9Ion9rKpB6vGwL2TGFGEo11U+u5gGceyhZBdqbs7Nyx6zmLg7duYwrw0UH3z/
VUx5JT/FmMORskh2YHkvtmBmaLcJJwcfetefi46zg/Qsz1ZE3lP3cUftRQZjgiSoBt+2eme+whon
6cZub76E/Y/lLOBD6vNofjRCmdjFRhNt+TQTtLzxmethDDGKivzthKc1Xfqb+SfUobFZ5qXgWpKB
23NPO95KMaHa+bMyFlcYBrk2LgoGU4kgTSuqeeuYzhDdL1NC+3C//y4bWBlr0OBXIExgNrrKfWsh
CB0Iy9K99YqhCg0oXCWKOp6n5bxk5ddTYnsTD5Xks7KCRIsPa9VATKAnM8vVr508x5fPIkdGAElk
Nqc6wmONFe5aFVoyL21KG5yrA1Fmm2maKjDjVIDH6NCunuaDu/sE1Pw9COS2+YAnifGhX2ruPOzP
AspW0zVU484cYTQcKk0Ips6QmjU4b6ZPgjxnd/ZI2aomO0EfBsRYUiDXxsgUOpFrLktP3aR7OHBI
ka2Qx9pNesenc8Ls7ySJ8pN+a0VG1Qc2Fkjwuc/NiBkQ7AolfYrHIXWbQ0CXyRSSTJgngh2g1pdx
q8AUPiPYOCquqCwDpzHf7hKJmxVOjFoz/RwgdKlzP5kj/F+LvTT3vLO6JVT2OED9azfvLkVdZc9P
zhHUOJ7PeIRJTHFGFreKWAXyZW7jSzapghbMAFlMn+FvIBe8giBLD8Z652Fly+0cY7w44xeKDwm3
Ore1PmalZLcVnjMgEMB4KX97DAhFymfIMapzWT+HwftJji24O8x4eZ8uUEvGH7ywBe1iOEk/ISdu
A3Pmev1l0JY2TBvbI+2oQfbhCKFPXF2EauEkbp3DCLIth8qyGTCeNaQ6w6SPTQ40ur8d4nSPUU0r
GANRdEwneki5eIbAxbAH2VkKR++/TB2KTcvJS/c5iMfEs2eKE/6gcigCGB6TZqJj4LkLWtY8jcke
xXCDvPQVBO032pYjkzKQs/I2OVxXm3FqiR6ZUPhi9cDwyJbVwjOOFOU5aXh2oa9XzXkWZ3pK/H8+
MDgeu7et2JB0p+aVAYSi0mtO5yshI2c1tkRVtIAxg3HM1sxyUiyZLlAToLHg03Wtrisl279gGt8y
P2qdLfPzeZ5ddBFGO+vfn09mydsqLbP6YM8WnY+IycsdAvjnex5pQOdf3s0s0JZp9QCJ+9nt/zt/
kstuxh/qHZ8YILA4R+fmVeoytd0lq8zpVJSSe9jtK0laYJeSF/AtDeW02OjxQCuxptug87rsfXxu
R0VSho9vbPfPtzRrj7hgmZl7C7mqrZHfYsbZwzPP1nG2RNAS1kfVg+ZByh/Q+URAZ9uQEoGVkYad
VzGlVS1UZNmh47JF6WMP3hzhgcWjzf9bGdyUNcC0oVynyqlPSlzpnjQnXAlpYCXu2hIYuQBH5WQx
Gtf7KWIx7dwCozo0AADk2s6jWT3dFGQzi7B5okpTffxDVvBe9et5y5fo2rXmI4PL0sLq4FnZNP4Z
1TOgSIS1lIDEOepC4dR05oCayxKhaTDhDDn1GyMfut0wgLTmpL/JPaaT4LM8nLdrfLVbAfwfr5Rx
Ow+1w9MRllZeaCf/PbHO1EkM78OvjvR+miM/Y9rqLnAF8i/pF09eh0H7j6cHW4Dy3uyfpezq5Rdw
xfxNA6KlUKrrwS9CNu/wTJt3mZc1dDVknwjVSFQ4qMqgIMRv4O7y510Bx8K1xhcP4/nVMXmMgrWh
gtjSRjfMSTGpG4C34Q2LZgkTnPYwk/pmEO+EEJLnarhROkbS7USbzP+M+kMOxBaIGWl/k1MBA8Ab
zKpB19tRlzgsR9Q1n7g0ISd3BIE9tzfjHHGfSINkI4rSizx0ymjOzETZ2Ev23sCIFGgXMjxlRRum
Khbh4zCMBZ5NlR59ikwZmPg1gemel3XbckV3U+cdxvsHnslacagvmg300Dd8MveSuV0v5rznzIYS
icsOiSHkravs9gw412mzblsDG4BmjaS1fbyaN5Py95EpUGQsQy0kdDI6m5bAuW4zpzic0BUCeGIl
klahImKWVPYhd/xFy61CJd720/5aIgivIegN/LhCVpAx4Kjpw0UPco2Iau81Zz4yzi9gm1u3WDrU
Qr/R6P7QQai3d5vTCuZk0bmeWs7iSTcNvRNeFgKwr+z1JRkKEzpnMlvhld2vhM9GajIe9YVWI+n0
T/TmBg9qPy8ma2dQqPY2S1+URlg1myi2EKHq5sP8X9coQdffJlHTagqim+bdFXBAl/PZtcUku6uP
nYBPvpZBtFg0HFknU3f/0FwVi54qi89qZSUzpbsVxyE5dH3Q6PWC3THP62SSE43CnjctKCDh4fCE
EQSPB+4frzMlEQkPpM/YUf8y0pTZc3PmjNwICX9EvmYXDFGLUn0aVqsRtSHKh6N6xlDrYhoK6tGu
/XVKXEt0hMDjzQHI1LN/Fqu+vOU5YUA9kA+NQUaYXS3LHopR+lGwLJ6V2DMMMHA723fxH7GOUkFv
hVBNOMtReSbTy22CiZiZgGwMC74ws4bDa1PzXihjCM1CYq0wr7/blpsYlAkFmzNMZcN81pm8d6/K
3IHRGuRYDueuQSvHqnk/52XyhdgT3vX+pCRZtMDyay5i97/lO7FteHH5j9B9W5KO9bYQyuWBnVKt
8zU6Dvi7Ju8EKeXuHO2VcnRewcp0v623ZZ6QMZyg00kq5t6A56T3IEljRNVsYuAl1PVuu8teUUZC
76tW4xjjgodjdXIM1CEWQ8nFxg/ycSBtc51cUHPut7QydqJoh+566Be5DLUAj4Q95eqRQv3zkN6h
qOLhj1O+oz1DLgExzQmB6eqS6iNRdVUWFfgGX3ENCT2kOB7tcx/1DqXWRxf3tTPUgdaIqNy+vieh
dPTbTJAlAql48tGg+W2UvFX2XCt9nj9lc03kcdNltqszOqSYApsDeOY3Ycgs7og=
`pragma protect end_protected

// 
