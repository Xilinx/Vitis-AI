`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+GzawGdEcIuxfE2xohKZ4YfAgNY
udze0/JpwAsGtIi3JEG+f9Lc7KzDtVo+7e0axUtpWWG2zchF7YBRjZ26kg5u4E7NrejsKmQn4oFZ
2qTRJZGb5SJ+gdQBQzowrZ6DlCm5Ybvng4Y+fKORBe4O+BxCB8HAkjiHJvTxpq0VwrUrB2IS9/yv
BT0mW1nWT9cr5BxcHY80c1SIh2SWvSjyo6t8HbC5zSeDNq/HCBlFXopiOaiYhaqw47uoKfrNcZxV
H0rTHABTaroPjtWH65lcfVq2q7XuKEtNxAZHZd+IysVF8aDNUa+0/1TDebmASfxRYR88xkW6yUol
9BsnRiDjoHKKJ1dokEDxPMXN/sG58MZZa7mdJT51pf/XKB8wFBtrW60ZQyLywtG4v1luLKYpLAuu
Vlho9aV5mGurt92qLy2WPo8pdiwySb0BKFpP5F/DGS1j4d0qW66J3jGqfw8dGTTkozhzgCmdiQcG
z4X08wIuld9Tcf/eIlUbQDKstBdnieaQJaL029CiWQYzETIjUJltuBy4YXVknGIjvQbUKCPhMW0d
wOmWv96Jt4eU87yGHEKzoJctFUB8vT23OjnNrgtWg9W8I2jVIHt36lDM3mY7Encfnwmtl7Fk3k07
WC9/5K1o87V3SpAlrYa9vpoHEWCnVh3MvX8ZhlayYXlY0cPm3BHlK4NKANJMxD/dzTf/xGqyzUrq
nfTL4t3Uv98vzAP0uYSeQb53dMCmeBopYgOvmKSLT2JjIR87IlhfRXRDCR5VG28LYWBKM4cXCxHA
Bj+eRr+4TBZNXg0fhoeUb41SH0dFMB631AXDE1kiriBuRoGtS2Ck+xYsQlrTjXjbLblu5M8V/6v3
WmFucQRZDqzTrEYgTn86cPalUF4tYXvW0NaoXBYhavtsW1TxDXVyUo1Td3eWUxt9w1nnfeVhpk+O
5xvnuwPxPdzWV1GdnmD6tx/zxRQgDzHZ3gKFEnMvk5noN86dX9STBYeUITojkndsDMzTgz9eN+d7
LEgqfry8Q5S+/351Aor4pD/WpzCNX/tvd3ffdI/xQ3H/0ZQGc6RDkdkDtLHESN0z1z49ySn0WIJe
ihfPlAemLnpQU0pdam29mUxgv1qAJlOuTfsHLkiQFbDX8w+VlvWyXWpCiQsnNYyHXdBQzcheuv9p
55mcyvxO4d3kRh/kF7RiiLjlpfgPBiDyvIigIxZ2hZPUtl6aQPmTyaPMoqfR1FvWLuWfkmBWbHc5
Ps+kTR/alyXt/l6+4CODPNeEJ+woXJOa9KL4+YpGlAD7Wf1EMGDT/InVLhDG84xeDIFeRIx6GMFF
c0JNkm7PHC+15MEVReQFUwDWUfyW8hSrle+OQEHet01Xi5Z+XG+BfIVQkwqdGdSjpLXfUei3xODC
EkzZ0gVN5RIe47vxyGD0Nc1ciFqYg+3P5ac1qxt405wnoanFMQUAm3/l4NFHG4fW3BlYQFiQs46f
JE6cET+auucyOGhwUbQkrXpGJ5Pw+DB0T8gzMl6iFKkrxyEG+ebuww7/YLPNyB3gkmwxww9QB62D
F3uAVbjXT7DGk0PMZfHKFbVxAoWg/8ufNG6x6HM+3K+vySNxq86VtHs08rCOaXG0/qopkCYoz8ru
7K+qbCGcCRn3UCq2/EuOdCFHBv9bb5TomOcFkrf9LO84DftmW/Gp2Mq3qMRHVU+ITGRhQfLUJNcW
2pCtBxwEIUOQf4B97ywMcANCNwbdp8n0EImfyecbNfZcftl+/KJn+6n4xavgD1nid3XsHGKHo9Ax
QxBT8QLTJ+T1p5AHB/r5SweHdJEfEyMLkYG6KKhmtZnBsfrQb0EgxVq4NSU5PGQ38+BUiwKs3iev
p2IE3klXxAk4RxzGYXcG9IzuhwhMzb3ySteiHQ7OkmwZWiCxOvAItsrGXZfoA7LM+g6EZQXAmZAq
PfVcHC0w5b64pINdYbc42nIKTFuzoJSRKBw8ryw+4s4UtZzofRJ4vz6D8NFgwJXdvvgsuNoC0VbI
xC0XNBOYA9518uDcnNF8QzFTOxEk6DI2wXwxK5DY0dMGUoelONS4Vjl1BA1DTWurohlR14UwEdsw
Ys1d7mnRu8yeXjKruEd/WWlISrrpx4L0+BrEeLnlgoevpVTWwZLbaRbKWE/VjFzOccaIs6/OmHUv
D72kjZpPQgBb1yCWUU5as96MoPsHtwSbuL6PJUfGOYpm7hsRywtaWtJGmbUt1vLq3BBuuKWKJzhG
Y3lUDD7HEjwCFQKeeL0C9PFF+vujTNtpQVDKLZtVMw5o0wIRCFZQkLUzvCh6Ofw6v7TWBubYW8cG
dve6CXkn1SChG7eTTO7u/VmaamJ3dphbPE8EN8uxZh1bHDXbcfqiBjtQg9gp/XeYnVvPEvDWy2HJ
3tO/gLPO1Zoez6bf5niYsYqdigfA5JMH2BUt54YuA12IE66wJN7obK/Hl6Z1YlnuLu3pzsHTXGI3
ZBHlNFkJmFPVSF8gZB1YduDn4t/eOKcN/U6CzHv1n6dtdtyRl3Oh6GxgR4S0SEts84o0AiZlxUa+
MFlVbiGgSHwJqvIDHmcvjcb0qjGJDn/h12RVLF0J4F+wicaXyktGwRBNpT4ZraLo7V58utw5GKfF
zMl3P0V0XNkfoyDriMzcInpNqh/w3p4XK+hftHkLhxr9ARb2kogN8PKCE44fbRyIYQO9r8bJDL15
iKBzEMoo0eEzp0+ynetbGOMF3sKOlDIldJ9/79EXL9r9y9jBQYnJk/s5ISRFLQ26/0Prnd64DjG7
YbW591vVVE7yjYr3L6oSDFXsMGxoqA9f8pu0N0+YnBa+T5w/eMf4zFDrKpoCJsBo42vJdPIVMtwY
xhJAEjciQYP9/Ggs3VM4AX5CHZLRYVY0Jb1XUnz0wsG6xowFnVIcDeSWUYBd+qOM5oZVLoqJvvjh
hnyuxuwtoR75HqY9UknV5GX2bAqps9LcFqy6w+GefGchv/Ftuju1QLSukV8lVUmnaoJdF+ObnVaO
t5nw0IglePavEikGUoIKLo7SyVIxCDrtbIt8S6I6DhzOpC5Kx5X1AmLNq+7Dnr790VwfKnvb/58B
8b/Z9dGgQnmIQ/FECLpHXGQqXDGNkIq9A+EfPjHxWEJRgSKZcUgW7XUAb9Zkag7nvOamKDhUI4Gw
Bhn9GsFQjNDsjZnEWtAd/Jk+1JpkGtyeOCdZRNpDesPfqJu/XelxrGIl7qx7qzDWb0eCrCRshU+N
mEEqGJfkjHJv82gcHWZ/9fA9mjA2pNcAjNfMMks1GoFWGOcaYYfZhsfk9tuwnYceLjJGgvJOkxOn
e2Hl6gM6r6VW/7SezbYkbSdoAHkv3CqwL4y/mYtWl2RhqU8Ndn67oEQVB5VHr6WuRj0UHq9KORAT
ogfYDcyTObNnHCRDhFFZPqoOtHcts/rBaE934p/dfcNuhWObNsNLtgWe5wcoZ5/cPSGVBAx4QcZT
QVPh1GnTolW4alupwF+jyS1ACJsqm8w7fjPHaISpbyet5GHN+v4+1SKiv1raK+YrEb1DImGFFAJo
T/GI0lcEcR/Ys/Y3JKHMRR1zx53oUU468XzQXkSuy/eV+7s6/xOxuYnTqxy0YWCXnw+opG9FkYiY
WRMOmi+FvfbPYFJMDks/P7HxiOWfOJwCJXHPKMV/roUOvdHoLmZyLpzBxGZ5xEU4IwUAI0ZwQp6Y
ynXIrJO2ILo9PA/p8/PyRRdxpUDOsrsfSfkKWSozFZKQyc8rVkrBKa8ucrl5L6JOl3ikZ/lK0pKQ
ohPbF+GSW0b4S8hrW9X9hHVV2OBjpJRZIHpIT6ISMpoJk6sD0Agvv0PPi0S6l5EyDS0/FYp+ZOSI
dTnAXSZ8hg/tiI12GrkU+hcewkb8+tlbZSCrBXwdolwchiZNdAnbfV2ZqoTHWuSjMDazc8flThNx
ZLJYvj3Jr+hipYiD9O+xdhNhkkbuJN0c38AUkA8BUqFDEd2fiL/vnHCV8nqa8QvAIab7RCmQbrVU
7WGEF7mnkR5Btbkkf1XYFMd4oAM7/zX6ohzG4KpdxyvAfdQnM3mr5cpl87N3Jpue9NSnQ4yyJevW
QbviaCYEL70JFjlh/Erf35VzQYXdWfOznu3vxey39cBLzSxEIzLvXoy5xNUpRtBIr1ajjorScBUs
7GIv+/DpT21Sd71ifri7mtErtVD6Bs95P9i3LP9AguwtAWwvfBPiy9YrSggx+Ffv9XU0NNR9sVSv
nBr2CIBwhz+le8V/FThlJwWmX6dYK2Cnlu4jn/UjDSLE2QhUq1hLQWx7Q+0d82m3HIL8ppZCzumJ
vzdd1ytmTOI09BLZKNX7lGMOa+NGy+8Sh4sqKAHn0N+O/XmR2/67h2IVRixAD+zkMVjueXXSR7Q0
kKW+5O2zcp86cVWEBf9polAq0ZrYrRFQWaOcmMYq2f5/hGELSoTDqUpsQldbqiadPjYQ1YkM/JJk
jZKjo4LhFpAp4zYW2GPXUbO1qtQohTIxsub0MVfxfOtO35qpBpk1EH4mWMBxf/mDbvBM1v95tJ2J
rev8UrioY74BYQjBO3HezADtgPs2Je/8q9UxaTxTrGduWIoTyrMItJ/G+vxBQ6Qd0xNRDIo3yS1G
VtF3eYMWP0KJuxbfhI/WTukwr4l2rWrt6EBx7HkO30wnC1/rUu5L19QtvETwZJbUt0GHWW7pGeSq
jPOqrqVtbyY0NiZOV07xgCSoy3wo0/bUKrbG13zfHM8EdYH+1PbMVMf7RynBlm0VvqQUbnq8+GjF
DsQ962hjY/IqYsAa0HLeP2kyBagNV2KHrrsLDN4QDArzT+6Qvl56BDjRI88PVdgaMq2upiMceXq8
BoO8nd6evw9KODOM+MyTcwEVl7CVNklmlDsjSR6g7tOinU+8SynL36WtbD0visus7quZzxvDE0rb
EFDYrXmWBwbwvstq1nfSZnDbkYIByr5rkJDJ9awLDsfpOjeEcLgpmsefGY/kXoN0fThVuHpRDcW+
CVJIsDPwjdbp1mm320ONRE87whlbxpiR/4m5fYAhTpsb2oZX6bUwIwJ4dzp5thC0KMpG4rqpqzta
LzMYtOOeuhJ2OzZ7B9BFoZDD6VWvHcebCj/hY5QqFh7nN7uYAJt6+fbqXGlapH466QN+47edFhWZ
SYMd25O64hujKEdTAuYRbIQiQOIhoIBdwOLCcMgYpe7Ru95hLi9wcekD16+A6XXlRtJ7JDNqRw/z
txNSirndAswxAbq+Xa2XFqtHJ2URPbB+coJdD3ebX1APpduUnt+cbXRpVTGCGxCMC7C/KAPZ8pwy
ZvoqZxTy9WMtncc0VPvRIQQNjo1FiCclG6XzQ7TLSsks5mqOmpr/AAlDjyRkI87HpDmBu2DbLS+p
mt1AEevCsAzUdtvYhwWND64spNlBi+66962Gsmy9ZSPbbWEibnCGJoBkuEd9l6Ra0LtLpYgIonG/
DsXInCQt4THrDmGmyjmtgY5IrjLAR3mlgJV8Oc9XXm/2s+17JzI46gjM3EcWpZXdbxXjwWd6jQWl
YTfTH75z6IfL6iX4K0vYQSiU5d9h2sbZQK2Zg4eireYV8ZjEntCvoaMJqJFpYeXvseH9Sd9pipXd
Cb9uMSv4Z8y5zz3zbWiSqeMGgEdP/NdocSp1YfugoOL2WPwkXRtqp1vuEdOr5O6YxBpBxQ9HItk/
tp80FnCZrZRaGv+7v9YOCPkQjKVcTC2k1cuRJMRpqKXuWnZ5m/79URA9ltGq6EJ/GwQJXWGEBj1A
NtWlXefR2p2tdTTa6WJWMv28Mw2ULTFHRln0QtZ11nT1Su19suXDhw2nugbAVES8zXFIj3vwoaBD
mfJbXFai4Xy/CgNkqyjD6QdEjMYN+xaJAsJsXkCYFzmYn53pBlDf9mwp3WIQ8riIonAqh8Q2tJ0s
aYjojwqVdWGfv6uelbFg1Kf/aRgmxsIkxS6U+waNMqhcoYUBOqepuF7e1jadKUtF90puS3vG6IYw
blbDsHghLI/yT3wVa12OZxh/Js2NY8+Hnf+CTNajBE6gN6jz4BdMCxY5e95p38GXfKnzQIWwkajg
kCpPE0TenXbFfFhEpIjSl0ZT87GJcOr55pxtnT3fy5Ho4++JTfn/2CYst4KwfrcTN9A6UFDNsNbK
SVZr0FHnDCLTNFjDl9MXVcqQhCQTeOKK3mw+Y9U7U2p0G2m66xZCmGyEOKO/9cNMpGQgvG8uXrMU
mtrPD9G0CqnsxbTp8HhuHbg7qWNFzxVCukvxdFUt7fRlaU0vV5hjIF4cSjx8Tc1NzWCXmu8lcjI8
Q9LVm4GHetz11NvD8GqmEmsnxpH7EZTX+H3bJo8QoKdpd4rmONAJVAETEqLyc9v149avq2rxQzXp
nIow2umArfX7uGTGKwtoqPwjbi3JiBP2XJp+BByKP0CCx75XkXGgVHLpS+GWYZM6m+b7PqjoTn5v
rBMHT7QXGRvdmIb742AVbjfBFNr75+wONGDo9YKqzB0N05WgXvTrVmo9oyoXc4kb1u5yCKeiJOXH
6EJDs6tmxTDHP21T06akJ17Htv4bZW6YZXzhzuedKXqBuYNycAZa9wuCM1FJYMdgCfKjtrEVe44G
CONtUD3YN23oFpXQ7Z5oYCX7m6p961N5N0MmVJXzGJczcmTT/UBuOFkFSnbz0Zaclufvfp96pq5A
jtp344vO8KCmXQe/UgNwT9NKYQGUhZkx7/d1xJDT6UUHRwNAQk5n4LVeCRMt/MI9TCMhyI6KKMCO
wqZ8ro+SaEz9ittIkgvZFIgxk5DASDF7rL3QonKpKYlXYgY6ORkn4rYHd899HS+YJYr0BVZl4vvs
GvKAFyjr/0eEeYB1ptCIo87sBtPrFN/QTHI7YIqn0zm0DxV0JT41jj60EMVnQ52QaPaJguHQh6bS
Pr8fP7j4Cp0eb9FKWTtcKYaMUMzwWLDb3/QhYgtDred7RY+f0POl1XKBSHNsHkDWycnoIRJZXiYr
lUVTRAvhnduw2mXkRwxP0E3E98C6lqo7lAUwqrJ1Hzs3BYAc4c0If2FnV7DZe7bHLJgjvspmLomt
IYq0Z7It2TlfFWqDuZji8Yt9zWl9kUS4q4l4gnukY/VbDqSeLEbb/rbsFKXvoy2YUPNl+b4uO9pD
+iQJN0KXR9fbvQLlpfgTFVQNC7EzupsA+HkSjUoATOElCgUAyllnUqBdh8v/BE2xEGfcNxnq1NRs
IK3hH/5QTGGMRghh/kNR4YW0wdy1MHW9abo7klGqo6zOwzvOiyleUPf8dk6eqZ4F9QsdS8WbGlgQ
Q3U+2NuavM24+PCE9LBp9DiK5TgEMLBmW6v15Wndc2e1RfIV5zErPt57c4Ic04ZJF/Ez7q8IPZxp
KauwJ4PmTQeAEfS8TGWG3tuuPM7fpEYuo6Xpx2eSDzQte+GwRJpK9XuiOmMnICehYedQyCuxQ7zY
N3Xeyllcr70tMUYAhE0wb5jQIvRCquiFPnHv1jNJLF3lQ3fj0qMBr/03qZoAOHfGj3yiXWUmiVhv
3wp3lAtwbwDJlkqBSNaLTkMPilqvX+bHlIbX854s6KpQinRH0aLXlrhNgExk9Rn76H6K1Q5V3Cvq
lr3004amCrDSWJe4czgWgSKSsWWZoTkOME99PPa8KEztQ8gVf9kLiFPx6qiREfh6DdwlJiXmuwrQ
MUkL6X02+xvO0YX+UCYDLEFCpBllBSexMY7Scc/dsSr1TM1dfyxiuHgtY4TG9K8sNgKOIYWVKkd/
/7kosTFDOkfwb5qvDYfkazZ/IQ2qqJfRNdz2D6Pn1APo76S6D35WjaWQ8zPyAENoXfm1tgl2Qs2B
cio8DrmJr33BN+/1URsNrL1Q9llWFMQHlcBGx+/YoNhWNsYcZBP4HrMH/4MALUwA82GwEJt1a/BX
dD+SvUTP4Pr15SuPCPvPIqDHsKr/5/1e5WoKRqIxzuvGl/KWZjp5xpgB5LK9lWhL+3282SCIQiYK
GU00o+YTn1qJ4iuXjNmUtsJpUUIUYsxrIkhTHX8RgM8IVzha9n4TogK8L23GjQF2kmaKAXvF90ES
O8WQfhlBKbeR1g7QDE4JT3WPY3/AmaT9CmVANTSPc8L9HS5irIUluGHaeCX+BJEtEIYAbT83CIvL
SIE81/A5QxxDxo7gpJ6wLYFC3boLqgoDhAPd4KvxIyrQgiyiGQ9Aipg9FMyFedb87dy5wWthpLaU
X6KVf0Sa11udGM4gsJqAiDi1UJQYaiWuh2aybWLI3J/HISOe5fsHwYndp39rS1hdNHK52EREu18u
c+IVUNIpCTZSIzLEzBewIu81/Jlbf0vOE9LchyzPs5Wz0nP8f/WiDq1XZ6xkLpP6eHoHDUnp/q6A
PdXIMRoo9IuLIBB/9duoazfRfQxhoG3pwx2q0Sw8jWguTwhzMhWQIQtyecycuKjmznfCxzAtJh2N
3NC4w+4ApySCoYlRdnXktJBBlFbI/Vo8f3mVJAfR02dV8laCnXLulJnwLOP05v0ht8i7qCwCOB6S
V0jf7xg5wE4pTtInmNGBKIUNBOCzkNAxeUDUUv1xgEU8KxGOhq6lvGaccgOTvcOSalYj8o69DSh5
s2AFB4NrqgkSw+OUur6akdt5FGQpZVxBlGNd0Vi1dW24ER/kJhGRFzifJu3eraLQfN/zVInEVH8j
QJzQPD3DWslmbbi++oUYoHMQ0yRtdV4Jp75U18HbgbGT84X7ilK4rWQWJ0IGvXzy2TnoDJEQq0NE
EU9T8swlFETCjYRPkW9127dMnFZrUnxipNnuGedQG5Zj6/OtrJi/YymmRy/UR7o2IasD4xlst1k1
X2v+vE6peIHR35nwB8fyW9pZNQOnXnsbjtljJpTwBOKEOvf1JVmWkfa9QsBbuUHwoXo3wOVEMRyg
aGz0hUZ8KJrDORTtzKReBmU5q4al7BFQ4BBAJ14FyFXedzWrrhoJcthuL++P5awHGqGi/pItGU3Y
uN1JBBk6viCIfoslUAMb5yMtva02+9wT2MlTaXNGD6M45JZWzROxOpcHZ107ekpackfso1pzqQb8
M5xdmE5vYad72cLUlE0w1wiT3VmlB5ElgUcFMvILAP8+N8BzR9jfejbGGINw3WoP8eaqjK9EAAT2
/QQARTI6Me36WZRMz+atbt28ombVgscSAlTw6yuh3ELQwXTbzAMZpTux0Go7sWHkFuqHT4AijKVR
7LhgV0+nZCUG+52OTh5TwvwJtGirBIBH67XQQA/kmjGkwWcQVOydTwPcNnfjJLVfzOQTR0hDIBOu
cqEsoGS7m/crwYxjebRSgQco5iyCVJ8dKA3gYKpakQa94ErXpP1aFdECw0v9CWOLM3ob9TO28NU3
d2dRZ90qkI0aqtNOYK1RzvKeS7KG5Dl5N/4JmUgIb7f4hKTra8RN0B8uDsXIog0Con5Z76hPoC23
xFUuE+ilgVeRQL5Kc6fZemMWU2Lif/OEB85dF+ZaPui/ENHWWdzDCcJo5Xs31XGi9TpjtM7OBvzW
bq2/+SxDTDFvKhEOs6pSYCMD/abzGMhPles53V2BiNbuY059jD1+qbNujswMjX0ULKiCw8bDbSke
O5sN0Mzyb1t51GxmPH3/hpSpd9AC3u6BnFdSPCBsbbxqPSTmS5T/pYojBQj+6Coq6noFBZE6h/kO
qOLk6HqT9q3s4Qm4P2xwnckhGbWd4xsUuwwEAYaF7IESL//BKoFnybDWnL/ZvDCI9kQlK34nLIUs
Z95sAr/ZZlvWiLSyqQTtvJ8pmS+aMCCK3xqcDmHC/QueXbrh/CUkfBo8m63RMdCKwNyV7sP0zft9
f66Q5CqgcNA7u4OhbwCKCncs0xWaTzezkK/CEOiPfpxflid+XYqlHW4EcxbdIfJj4dsStGx6mLdm
4HoZAi3d3SykjfNQ8IPBbt3470ngPgwmH4P98dP0UOjiiMYiqvVtLGvxDIsz6aHT6p43IhjaHdeY
P2afp1BD8lB/6ESTXd17IV5FWflDyQ68SC6RPz8lo1JjfiAkDSJp9bnwgozabpkQK3YW0tfVSc0b
Ih5t0oaTJbl3ZBgu7xMwm15ek4eIMM8bc+/5+RFZEEx4G8hVGU1Mdta54osuP6XEwnpr/T33zcBo
ss+jHMse9gXwDmYTGfbjfQv8qtjMu2zHoTCYolUTq64xZQuHrp/YAIo7pmky02E7dYJWKM2LNA8o
Ns2Tl4bF/lzLO/SWMZN9P3UW/adr0wNiftYE3/deQnK4KELYcBCiy/TnMxXx2hdxUQ03ocp5Mezl
CZuqL+Th/YhzT4q/YHGRXsFJAAJeYwCWF83CdhyBvYVcBpYqBX7wfBq9VQ30NKAILf4UOkN+6XJv
ps8jLAfVOheiLvsKUl8c8wJW9JSI1qIcCczbiIjjRTzfenDuShlx+4xZFArhO0kjVAqlcAhFh6Bk
uOjvzhuA9b73Y/aRgap4430eiL4/LXemblecQUQqtbgXqWU4JBs8kmIJEnH9/QMYa6JFZSyqygY8
JmH7xEpgxAKDCYqO5LAfAkHJs1+Tj1VADRjsLu+pqI6xvmC9Gi819ENKe+2Xk7cI0zbJpU9b6QGQ
CjDpt9E9DwPna6lIWLjZT+b5BtL00Y5AyKpwD+P+5W5W0v5+OV8TMzeP/cABykaJlyFiVjtcGXn9
27StN0OOPT8lWghwTC0zlJ51IxF887UG79ORdixe91VRe+PImoCQDIdgylfy9hnewi5oeiJS6gg8
HzmWvOcLMBPL4tx9ByYtyJ/VWv/rr/Lh0xVbro9q1X+BgkTl+jZUOpYFGcg+yo7tRwzTq7GEwl0p
CL8WVXJ6MiVzS44GW7FNTuXs6qP3R3NcQnpozr4WAas0/sXf9jIoEUx7NW8vtn1/xwTYNqnsyac8
214REaBziU5/+BVezMzkkYalfSJ9Zqi2Se0a79UPH3d3TLslzAqH8UzeyS2OuuAA2UaTR2pULtlI
qEaWSyi+h/iQ9O83oRpr5Yh61DegM5Hwa5frzCF6ibOfRa2Vyv5ewWMRJEuSst+AjZkervX4B3Ob
NJhtZDgm+keFwI8AP0biy7JiivEdaQH6HUsAi9o2Rkt0BbE6V/yjcq5HJT8oH8URwHZI0+XPyD/m
aDP/bQZdyr2snHs/cUMLuPtmiRE3aFc+rCgFhhVb3NT8tpMcCjniQt+56IkMLQA6NblYeThpSn/1
9IF1cKrSClIdbDI6r+4hQJ73G/YoDwnZemsWyfEp6S6vomvFwamVQ2adH9U3gMIP4MW+sLlYDWVj
yAXlKUQK9yr6qeng3GcBpvVjV3TyeA+iYJ+lSjHsXtawTtgYFwI2UndsCpc/fNgXegK/nL9NCQxD
EmYNZ9gLDDs84BKtZeqOuncYDq0EWvzmh9OiIMScYcnn0kjudmZ14auikou3HkYW9Jj0jTyByZg5
AEE9xbZAjT0qxvlh0A3o2/wL8jQRODiL9NJgmTVBOPWi+c88rFCupP0MbCz3IXzYpYu9xfAteZt3
rdwoo6JsuBx2Uv8GD298FFRfUDLoCZDAvyFkEisFUDrFtQ9RtRC6OaNSR5UrOPADQGByRAkKaWzP
NM2FNm/bVEzhglEBL7HPUxkgZJ/aObCo8dhdM8XkSQ6MGykkByqPKjQDqUmVjOCTw2uCL827gaVd
Yrmg0NQlVrRXuU8t+6SIKR4ZAKILlxQOwIoM5Q34mgv1zMMJcvCenOGk4tzROsKhfHnWfy7OrWh3
n8tOwVHsK0RvjsbgwgubdiRH49Y0ej3IDpz6oDEc0i3A4IxGRgiFnqYobOGIqbUlD0Jq1BE1TFXq
UahLRobcqblu5YVpA/UirrzN2/k1b9VHm7a1QasxXRFgYzIGF15x/Bglrta/yCx/tGW6e9XvjAUG
x+l3DBkuMYtJHrIxjLyt9q7bGgREpqeTmkwFtpgicYeLaWqwYUmPRwv6VspV0/bRKffQwgN6zTpr
4aY/UOLLwKrc39DnD8lCdXmX/KFNhDlPjcPBk8P0rizN1XAEYzvOMqb2YY4XeXsx80gqyYQbw0c2
V3npfZ/0kxJ/pIhXMVu+PWF6XXl5oT6Tq1+o8pS9k9drqRxjMRur/+RT6AIsafiKGopyOUwa6oPX
3goSORhvajQx4d8Qd3EFvqVP2XSTwy+3cYCRODbDFiClfwdtYRffFMZMrrEUeRqlEwCJ1FekW6KX
wH4KW+ZSNtzgjRlu84tc2fTUxlHEdfyL+gL1LZygE7i05TF989UoiAU0I/R+D5FdAhFF/OD+8/rL
aOEIlymRy2NpW5ugupWyi8yDn+mde17rO/7i9MBwmoBM/6VkqBz12rXjxVWnggezI8bqav9ttmkY
Kg+pwfT80dxWPTs1LtDq5+2jBWPx4Z8rcf49KyfOucxtSdKGe8A4vtVEXp3mKQy40sz6M/U0tdXM
2Ro2uuhrnkMuybt5AnZcIHVNAHvBTNrgRb2mnkCLf3PKaE/n56+guoQ0t5+gGlZvcK5WHxDr3qPo
juphrvU3+q3lDCxODDoJ52ruwa+SheORPvdZiMIqZKFCLdqZ1z7XQnEiLtBrl1zsc50LVhU7bRqu
h4wjMtyVzcJhFa/gTNYgDspsO6swMmeiGJdpzAyN/piPjVDALoMFR8bhNr5TmXFyAuvt1nzyHGlO
moqur9kDGgAdhZCwY4LdunI+b1pK25MxbVmX6BH9HnrOvyPRD7jTqoqwVgJc6bss+xO6pKGdjiha
sFduLdPXxjedw18b0MXwDjUGr/BVqrSL3BmOPJA2sFxOOR/1pqzTZ5KVbxLm9udiOM6xTMNUSEad
5U4baYEc4upiIBVpEkUtn1G4zgp3pu2iRGjOPARkuLfSCpsosQoN4L/iJhvyeaXwWk2iM+mdtScx
hU+ZVWy0iPsgvlhHzLqHIEUj4KbtrhSfiNqwdr/LlD7l2yX7XlvFoMZkKYzD2moJi5a4+W08Kq5w
Bxd557lPR+Psdon8ChpP9PLYf6+x6vOPAAkRjlHdY+dpmkc91PpSGv+RmUbogfeIWqTh7apwAhE3
40s3Pez1rvBjhxDYpfGuOeSU5ZcWT2ZHtjnB/MUOx0G/AIb5wPWewdPIZQTFx7SDYr67OWmD/m+w
m9FH7FujyK+n+xNFX/zk/XngfspuCAA/+gOg+yyJiBJxLlt3EoXWJ77KZDJwQPKABPFsVWirTLy/
EnQwZBhUeyikoV5WQFZsKa9W0bHDXlLC0HYMEfiqKMt3tulyZDIo/95mpGvmFEUidZV/1O7REpiB
TLPG34vYGvhqay6BIgsxE2H5bC+ANMnsCdg47BsjLwx1i5kheyNpxB3CIaRhcrHIX20lnBZPxxVE
/PyFuYmUCO/V5zLd2xuvnn1Yeya/opBiN4/Jp+rt0NYErY6dQVmdK7CFLaI1gFwiUltvD36mREHd
941jnmhD6RrVCWrfgcVFW94QHkvSOvNw4fDev5IhpUDOqDXxgrOlfs8uflQoF0fpP5eYLXQLUbC/
dztIX725erCbLdcZC1Ia5xe7uWwviI5egDpFPLI/QXbzz2bBQ4ri5XfSF1Vayq9/RoMCvrUxSE8I
+RVusQuEUN9GPVeqyulFPOarWJb303eG51Nrssx/UE7q5uWbllLemAeCVigCPohDIi0tHhXQ6cck
wqA/8A5kjM1/Qp0QiEjw404uv277Ie1CNhxVTC+Szx9h6D+bUyZ+pUrURd+P6RP+mdGsrf/PGrn7
zBwmoQoGVJ3vPKKlbtcfDnFr90pOKwf/0BFfQVfPLwVuzWy+u0uk2qmIKr82b6fAt+jdhDVwfZvx
rhh+5UngxS/pwrKoHHyPt0FQRYEugUkeeTMtVV6KG8c9OzadqlYukgWUotIxlH2Jb6919ji324E0
TBvasAYu3CIU8K5jSu0Wa/Ynk3Mleig1sOrOB5+e3h907kdflCOyWuD+O/F/WrUudPEt0R8ksZ09
+VgvIwxFbbUyk2T04BVm1OFaw92vsZIiD/rgVKdKQAVijR9ScRuXYw4ELCPsZXkWIUECgWhsynvw
uVI5EOufQxqgMpU86JgO1DVtanfZISiuhlj8RONdk2K3pOy70CT0nyIxxq+YEVFMMdYIqa+cnZVP
r7F6wwQ3NoCfoRFhkX8NUSMtJVJRzXN2aCZLqVzAN+v7DaBIPOWbOpxyMZXqtE7cRVR7mDbx898X
fDRWZWDR7nSFSJndAV4D7bbLPBN3/Uc84H2C0yPCM2TMdyjacpsyza2Md9xGbMmlwirJ7mm0Ydxe
yqrchjJWa5v44Rv5Qy495/9E6Xxgj4JpOnk4L7JekA+QRl566JCwX0mfK2veFv6f0XR0piVPZzta
XIbOX0cfAqAIq2oaw8DzFlPSGfvMqQfWkqJauLc3Uh3KRvuVS9760rIHi+HcixeuJ6cmepTbtX1M
jDiHz90QcSU6LqZKStEuttMYXVdR/OjYXWg2hYO3CyV0RXeh8o6xDEd2Kpy2xS/YXgKCO7FDGOuG
q6U9ziRt0HyImEAXBUefkest/T/P61JYhz2PEuxI/q1icGSb0Tc7zPj7wykiEcNb+c02IXW4ImCD
AOrZz6+0oigEPY5UzzAb0uTKNdH8xFi4TJqF2QMb5uV2n0vVSGJCwdKebSrcHSGfua2eJyppVEzs
FCPdAoYizMnkQxN06XIc4RCy4TE0WbCsP4sAhBNdl5m1XnEUTuOXNxXWJB8u/X9QbnlXeaR6siWl
BsD/P2GMfbRurtxyZG6ipy6gDhePkWTV6meAePxBYwIQ3eka0jAu4eSp3K9fF5Hp7pUYQXsrIfrQ
87XY91Drw+zaMuLv78ur8yHknmYISs8TekffgQX+S8vaHHWfMT9Q4SysXsofZV8CvfqVXylpvDtw
NLmywVbR/qRpQcRvfZtyWDQpBThKfQKcbj2NUDIlgpUJtvfSOZcICXK9YKkkQUoCk3aUlHDL3aNp
Js3TWTKyQ3ic5hJNiiid2hjCa5TDARIJ5vc2R56zRhIQNEeGys2GvBYH8JDBs/NLKczQ76e2gGJq
MS4uTXMrP9Nco8rmFrJuVNPPZtkBsy/A0J2IpdTLHuyNYZG8jB6mNZIZjYjr4IwLj9T0ctsL6rFS
6+9cGhf92PQyS9uMRrcfj0GFnWJxiIdB6QJMXMssYs4fdkTraMjEHpgNl2H0zCsZiNwFbXLkxFfq
soQ62iQjvwxyr8xJ3IkvLbiw48u/xTc1uPwffH8vgoD4QWR7CWtE4T0hJrcJS5jKmcxboOraoyJS
7I+6nFb3eYCIOZsY6lu2/YTMCjOHGZMrWnQWGdMNGIk1x1/zodDuX2Qng0pXiXM8MI2Y8dFx+df3
/zQiv9enjYrb/poCV2ANdZH61DzDkYd2ZlK8qYtGTnKOsrt/ODQwB8uTOm3KtOKceYJw9448OF8V
5uh1EP5zYpdVlL1w0EU3SKFjy/AlEr1vIjk8saSpgDhEfkGOKSfyrRuu+aSHRdZJ/Apqb4y65FHe
kXXPvv3dPMBCItiecxuCeBeMhsJhP0QBbObb7Q6UHct1LHvFsN48p10tSvw2L7aTS/+NDwTIi0nC
ysqM5PhpHKGJJfi1/PxtIYoRVjoQtM4uxPDuArTQc2dDfXnTL0/QAUd0c6oIW8rpE80YPqNROstj
H4KqUHXalovMeelIix/XEkl8yq0kdONoMN42BOc5kD6jS4WFDWzhmnZdUPVoyga6sQuOom3Se9n/
LV4ziwNpzi9OScYt+zWXDHWhopWTYsdGHrcw/EXotWpfYkyVLAKjVAouTs/l3RCWk1ycD8y48UiW
62zc1H06KNYRi3vxTkZXQfqd8N23qXLBIq//+N54/5ElaDTcaiO40z7wH482RS0v11Y9rO92xw68
vRlXB/jZsvXI4dodDL5Ex4BLaaahl9ZFzbK4Fg8ZNmexSNkAr0IQhgJCVQZjrEFHiI3f0qo3jon6
Q190C5cdQswZ0tRJDvm9+AJJmEXq50/GbMQTxqHm6Tkj9592zKX3qLJPBpnQbGQQAQnu+nyrG7Uw
QtcGqUwQdjqOhrPSkkvLMc81zs46I5yGLNisAPheDkRtdHcT16AmhdRuxWW1VCar54Vq+lCrSWWT
gRxBj1E4B5u3AefdbN2KAp8ehvz7zWV3np6fLXXmJM2/r+5FxTcO0CX/mS+INDyWgkGQ1KErT34v
9oFm/Qptxt0nDkGsoH/kyGcIQ062AkxkZ4dILKIIK52J79En5IwKU4BRg53XzAmw+O23GfsuGC2f
H1WMKNwep5B+P6ecmsS86oVopYjPqy53uCS2kOxDDbnLsldpGrwU/BNabcs40K8Q27ohS+0HTWZp
UiRznqjMKBvRkQlnyaCx3q3QrrjyoKHVc6j8BtE6TnW5wnlCu7k+0E6WzxUBRiiBOjwn8brulQ/m
Oj3cGpQrZRGW3g8QWQnmdTYl+18SZ5pgrAtOtnJwshfi7ZryJVGEIDT9o6moiGumz1e5LXROnoiV
ikv/0GWfSsK/hVNJtpBc95eeO4lIetTAXK1lPKDotf2HypZDaEr98HqGQaqKuBaYDZzDUq+7DBep
cJlxMK8Jd8em6oRIyV71mXR9QuBnDn89YpyRPrf6RLQHny3XFX1HmXgiNWpinywJxTuFlluP+c5U
LToCD12f+YTd5H0RKUDXU83NOBG1E06Y2jWsK6B2ii9wzyj3C+ykxrKqWZVrZGKBrT+mk5j+lFBi
IgNhQ2zcWJ/4gnK65ISl7oucCaVQSNZK2ISn9DRW/4Wkmpc7Dwv6+Fw+lHLVoA4GDtpdRi1xSAXz
f3xXMJsTT8VWMiIn0RqXCIM+Um6OkNmVPk/5UHWa0rxktjYKCxT9YSItOpLtKF+H+nXCwayPNy2v
RCXDdMH6No/g/x8jvOKjtnLq6nKzIIgF+l37mf3UL/ajJfKwBbonMul4D6Jyvxvd5Lp50hdrK7Vj
2rce37FKj/e2RElQE23bJsHdyxIxJ8nX2mJJUlP1TxZfzKc3D/Fytlk3ljufSULTzcCbruqozjLf
XXlr6THa3Q46lZLGre0M0t2l/8OJZVSY5mlhqbW6/mRYHCB64pbCpTJQ1Ye65tGdj4tJ/QNbQUtd
zYvjAzuZOJO7zJh52htuDSwY0X7CBlTEEdhFZP9UjQprXcQET2SDDLE8mtu4D0qb04kemdHm6qd+
CbsweMl/xBggykOCI/0DAeTDndquH7YpapxdpWlOH2maQQbag1yzY4E3+7giH6RtUi+ofibOsZ9m
i/d1LA/YUUNtJ2lfR1BVIufJkahK6RCUp/FbIbzNSs81H1yhoAcFEW5UEH4X6PbwkCO0+ys2ticU
fmUaAPPXiXCd5lnpFhIKNojD99T9tJx1NC5ORyafZIbqQav3QRrNTIr8UxjsZ5PfQVzsu2Ob4TBq
qq6X4NPp7Izn2nVqzzhJOh38QpIvQ4LkyPtRmTZNXnfobRwdvYp02rfMFKg4SKMnrqWLxlurojVn
28B8suVRXBz0RVXic48mrooQPGv41woBuRGeX6x47fI5YgPunqozDdBVeRPyfI7b+msWlj8MVQIU
SZsiimrRZD3JYsD/K+S0aAg5DuwBAlb0IK5gkxiOrD4UIakuODxptC85qqXTwBBJSLchNoeZYhuV
uQqYsfO17VIRiNCyHrTgxuMQ7Y3gq9TWtv0q8VtSd+E5VHhWOw7OKnT0Omvp5ykqslFM8xqEbC5s
fHfkVyF5AXAl9w0eYSJLglQA+5Y0g7x0Vj/iCSCxbS+s+wSoQExB2+QKt+xMspFVv9/2H3Gv4E9Q
AE/UjQboQirSHMULSZFS8uBC+7xRn3sF9Fs7F5P/ewGX++ngjvLPQnii8rN/4y70siiMiMu+WnFv
cUKCdDKhvEdxRRaJIA6GZOqhLKlqh8RwU4Uk9JG/V1n2Xv9heF/HsKngjJ8PIED5Ow2j32CJ6U7x
L7/DF793P0pAYSKsavxsidEh3c/hbLrkSjSdR56NbDTjn0M6+RCXMRul3AzFs0vPmE7h08+eC11S
/H3dRL/eVOD8Eaop8mmbu0l8xdckV9M8MBqoCWKpl7IkBqM9DQyabqcnXIw9T4NNE5hSOtA8r129
tgQzVCjaPxvo8vvdWWcUSPt+PGbT+q51nYrk7hl5vSveTwpgHXFYVrJwwqGfRLfJMSv+1z34gvW6
S9F5fwE4yj89SmzlzKvOCOiYDrIw4ZWGGdNY5C4mBdK6oE5zHnlpG9AR+slfBA7pAE60AGZn5dRi
urwbu9bk21LiqQFQLpZ/LAQPZUAsu/JhqrhsGltm5Ik075YqjKlfOHWt8khHZ89jp5e47zhq5xfM
O0h4SRhS9jPaVHoVbxYNTg58BJGowsmSZVzqqLmOJxBG7cUyg3QMTPWy22Jhnwxk/t1InbyoxfUF
aDX5NwSvgIWWVXjYY0+1KLORyVl/EaNpkCEksuSYcGcVvBLTx/rUD/ImNbgvecZxKYsk8jWl+tmd
Xld104BSHS/BSdcD46vmDWxU9f5rtys+0yd7qxUqkZNJtN4vemrQxgaFMaKKspNq4CVXhX61dtT6
xcZmBd0AOSNh+eQPJY5emDzZWd03uKj5IoOZtDpsH/xd7eaZsKI5P0Wuou9kC3w+7OZtNEwmzdD5
1zpyNpU9r/spFT6NL78XuMCWGiBg4Ww/zEUjEArYyw6wcfIiIiZfO6Cv5uVP/xNhkMtx6tiwPUp7
rE5oDvNVXgdCvJV5vwHmfxV3sFpyltbl8vmMpRXXhCJ/qiiA2CxEq9jVuUC2uS8S3mlOjNku4dcC
SzFquMWe1n8fWUCqQTWPHlGM5zOTko1tCNpSnJzvo62pSJ3cN5AjRcBZIqd48bAyqsRKYgOKuGSW
43ongHEnwX66dWY2CNTL7uMM1mQjtNQvy1daWejlYbgOE6dGLquUiR9sExugQ4nP74Ia3JNLAo5b
clxwtuGSdBkSY59OSDZlyL4t/QSVtMj3MYNKn+rS4eCTqsCtRNpubB+zIl5rmQxmyBLIjO1YYJBk
5/ThKPy8inBN2XPDApLNTskc25xktLJozVpkZbRP5LTifP7qtiIuZ33hgyv6t1aSTuHulx2PkdKF
njgR81X56/j/qDIPPk337H0gigpa2yy0rzF/31WhLuNSFBbzLM3IFrzY0+d/yW/f94YeI1ND9th5
P3rOQK2uTwNB4d2RXznCOqXozxyPt+333mgFNVi6p3v2RoyrmFMHK/pHdtyFDJRcejDqVFvcGcdZ
9Yr7E4ZUqkMGp/H2Fo2DGpIuTQOgc9jiLZ5z3T5XMj4gsWpZdY6KN98pY3IJA62cCPVdGqPKTBzU
CWzD4eJMrgk69PE3qrx6sOzHyitkLeZo3inl3YSVZwKW+is4vSYM7OsUPtRLO0KJa06szYW5gG2y
HOnQik+kOp0ybWv7iN1wKRbFUR2pXnQLMiKAc7wSoxFd2J/59qNYXqXnnJf90sZ9fLu5cI+F1cTb
ffo5RFDgaIOqKOshJ8ao+5+VGLrCODul6/xpHclPxrh1MTlAkzDSWw38lOPSjUeUk4lqik1XubPr
O9R2ecQAJ32QW2Y/hHOgoi5E+54ysWKlgiecuaFCJ2HdYXe6utwzlFLoAqNO8ODRBBiFg7+TlrrB
Ig5Xqhc8Vg5jsJP/cXRLgbxYIkehvqrUDApAqRKI+6UJr4Cxb7wPii8WFcGKpjGM8XaUVpdNQVm9
bxwBBlyfa+lOxo/nc4F0nWq2Wesf7ILLCn27oETZH8u9KPAdycDsuAtE5R/eTvjy4aKlmp4g7arc
Ia7oc+GvdTGtMdlfUEU94jop4CI2t5EDRhahwnwbumcf0KZYpWT7DH/0sE1dbi1TfTbnMENMUunv
naMfrwieCIRKoHBIgTqp3D0vJ3r4WiZMwmyzgHfVFg8hONpflBR6ER6IEmXnxuzvHipQ74Vl/eBE
IlL/lb880Hj3wc5efb+immwat55g6xQItJBS8Q4PZQWKHVNa7iGNVApuMz9MPkV1jnJV4yQScm+V
oiN/psjCAxepmIyez8nCxj+OdlAI7joElqu9yUj+vlmRIfnMcUfaTWO5/AIjN0L9ulfs1UItevmJ
wsKdPxymFDjb9H1VkP8HxeO57vsu5+LN53Pcz+NOiGJc3qGy8EgsdRwN/TO7fd/TWO4NCebXZlhI
a6aRK6jM6STfYOOQo+Z6orOyPHOQKMcvYT34YQIcEj8dLKeFgzg3BytHD8RNTTLvkpw1ZU/xJMXE
DIEUE5PLy0A/PYXFp+fJxzCBODhgOivivQgfNHXOianrcJWLFfa3aweEVhJnx2nsOdAldAkhntfn
yjzTsqfOzl0i32RQgVkyxH74Hh3cEINlSEXFSIrR6N8DhaH8unPjsskRpRtYjOTNGVLC+6BMpFPZ
szlUAYFGr9sK6w3zsTtGBN3IyU1dTP+/chZ1gIZsgjvecILZONzFmqnxFTlayAuWAalO24VDn0kf
JIh8LpPtPlQSX5E8dOr/2+y/CLOxLdTKjcNtFGzWCMoMuIAFUvQz3IDHOwtKI2Ispmd+cS+flZJO
ne8CWlN+GwX90l8H8kC7Rkb/V+KbkYXggkES9xcbjyiLXkwwyIwqMl7BnCtcpLjLMed4jD6Wg4Az
8cRWMZiIeW6AbFKAa33PxKiPhixI5nWsrgaO7x9j1lgnvib5lJsXYRxShhdxjwEYrvNjruAGN3ym
uSmnEPDtn3YK5pmmE15Bkk0QwnltFzf8GR3KY7WIizFCYpIuEP+TGz7Q2lNrydmubIDMfdGcapRa
iljcpBJznIks2d3YA2ZYYL4wxC8EEAvbR2NVELhcbFazvBDMbnZ8u1HCS8YX60LdgyTFeioR4+zb
b3i8z00f58MZwTbp6qyYMIxY8EqZz0T9VKsFCrRlq2SdeCemvNAfvHf6/HmuO71K1rH9pMS27oe9
hQf2LC+A+Xy+UQE1sBnnzdayRTp2i1LwJr4eYJywYIj3OwsDyrIFh1ZodHXb+8MxkETxzuNjgEO+
ijwKOPvQZA0wU0R8Lu5G5aBtetEOZaHPScfAhOgUZfnhFjoOSMKuPIRQeeVojjLtlKa9ify6lpY6
lUB/eNqBt9xowiGWosrcKneEZv6m+NPHXC+CVbvs4Jetqhh5pXKxdGGDlZwcPuc7pzZXyP/Ld0VL
GzmDlatHQ7yGm/FDIW185MBTmSRkXNTIskuLchmwoxoC4krwN44UCfZ6lMRLbPvsjtUc+l31bllI
C1m/TANqrilp3ntzJXCrhh1KgOrppMFln09vCj2kZZmP62o7NrgKn4vIDJecwTqK3WorBixJLF6G
9TvtN3Oy1Wprj8AlW0SarnaEyrxGTbUJI4L8gI5RKvp9IX1eAgBY1bB0MrBARMZtE/UuDqDX8SH+
RSWCNxaD7af6MSkUspVnk33iooRVZDt+jpU/ZMPKtzHqO4nz/66mgDqY4ROfFUzPXp+X+Iw6MsmP
dsLQRpsIC1jRW+pY0uMmCHYlw77RT632wySX/606KCuVtoficIUC5En7UjrBzXAZ3DEeOBIjTSzS
cHgeXLsoaViReFurtTiaqMxjxRP/4x/tMK695LKzi7FdvyvwYcxumxTHYnT6Nsz4H3o3B0I48tj/
aK7mzlDBVlxIzT5BJPNabGJoDsFuniR92A26HmfL/DRvjFcYqBlQ9hsDeAV0OFLL3uD5jF5G+6CY
7VUclbb8/WEdPGORkoGjnSIOwNPPSE+SUgIoQtcvYBLwl3BjeIWCOh5FJJDAmZz/Yxdfqem1H9/m
bdLnhrI+isoazx8UzwKaLUEofv6FdFBAMNUG8z3KSSRFi7ufqP8fyexpGbcgjdpbZJeCW2B+x8+E
3eMIKQbILtRbjXGRXHYJtiBrR/aNnTAQtfm9KYLY0pc7nQNOS4+uImUToC3l9XyFKHdRyulw8b5e
7GRedCno4AMkE2ZAaCGxN6lj+jqiABnztoeGGMk8aozpNum9cxySEwGRrm9EL1JZZHM7p4uHstf9
sM2XAr1qNRzYHw2fmCeijKK8gZ7v8hmtdM87mcXFqzP04ikkZvl2nuugm0RkMv3uxW+XWQ6a0ZS4
eyEkmvYVtKMiQyCDO6fXOvBSMiQOFPBlP82tx8XjVr8axb/bzXvc4A0AJ52jDh5Nhbj4K7mjeHsZ
OQXxKUOEPl9OUYJiSOdL/i/b03jlPpv8eAExtr4K9J27JDezsetLga7HsjxpTQyRlkq7xv1HBKSj
YsQmrNLM9keoYJ6zf7w7t8O19Ncp/q23y4euJ/PKqE/QfuhTkVxtzFuwwzrtAJViAmQ+/0h7G1qn
Ew+5JsEbBDHZExWC73aTKYFWJIpYSu3B83VB9DNa4xBvKJ6o0BSeHlMnA3sobER+BvwBqEaN83gq
YCj+hKZsKs6YyOrsEEVq4bbCpqfg2H52n4cT+xnRBol41kiP4pCsVCKc8M5wRjlBTUUhWaOkwyC9
vvzSgFqlH74IiYloXDnOThogN4kY+hKnwevww3bTcmIfx73DQMPKWSEFdL8S/Uwx/bKybHhtIcU+
FJc/AYo6+xvjQYf0GiJNkDxtnvM/2F9yFtM1SpGuSfi2wT3D1Z0skxhC6RX5JjURNqKDoSopKtR/
Cn4gegYQswLJ8vNlM+wQwxV52oD8g2EknGPab0fX3+AhjEkYKEYnNSYBIych4WA+AqV2jtsSYpI0
EgS2ALOVfFGKCEK0sDzKGYiE6KxoZVnUWlP9BNouhr2m9bSHJc5bf6MHZVuKPyjbLk08jiqePwph
xHs5HgCxpHSXnj5LK+f1OH5ftiPSOwBXoFZQM223M9+rhvIhxSsLgwirsAehBHvpF09oN5WhGgV0
xgk8wZOZ0FW9wHhw63qm42MjkaG9xCUH9dllGRSAwYW7qwxq/XwfQC1uhD9vyXT+LAAiIkShLOlm
634AS2JycRus7qGD5iVjGCe921EzUXW2Y8fw5BbXzNaoMUDh2H/z9ETsokdZbrNQtngunq2sMS5+
UFCBxiE6uH+9ZZw8BYHoh0zZMwAVimHAWlq2yEH9TR5GnK/bRuYoUBtSH79odT69ak9VJ0GzKHGU
0F93ITWiej6SUzL+DEtgVS7poC82ORG2j0WGSy0huSXsX+F7CMzfPvRczRNzhLKueK7/SMNiWx6l
01pPRSsLDd+K6FaLfB6veUAz5iQOvyGzRIjxTSgq3h52k75h+M1hKN6IYZ2a3R8XdtzSFsCu15wn
uZP57/LjOf7wLz0Fst8gVaboG0XPp6c/slfL52kYD1cUuWXsjQ+MT75+RT8P7MeosdRrxAV49NS5
KZy8AzidKsbgapgW6L+6gOgZIzFnkDJiLs9vNKAfzlMEExrOeCb5XnhQIImX+lxsbXRCEPUawmTw
TaEpBhB02PjX0tx3FidULFlERKZ/JT4TMgnsTRw44mi2g2GA/+GHX6IOLw8O/tjV+uRqYJ9FDC6j
Hg88kpwkU8uqYyatgAk+31UQp3U0KuNId67Z48PSW7OEOuIfNhGDFFYbsZeCxjUZXOoKNY3cU4WD
PNUmuTzEeSBKEb9+djPNOhAFsM5z8aES/zYI/4CJN+0a08HLkqwgP3MOwWfyESjHafhvd6SX1VgI
H8aeIQzYwQ3WoTvvO+sa3rqZ8J3LqOEchm5SUaTuPlrOogQH8S4tEOzcVLr9O1+icqHbbtycD23y
bgk05yojw6rSHpInvo14QkIAKCGilOTR8ph0htvo1h3knpAp7terKJm4VR7P/JQ3olVNbVqVHm20
6BNwb5lC5+c66JA1NLEfgC0lqDasllN6j0nZSRF2nVzUiWjzHS/fxcsw5ZvCHXll1M1+Y9AK9FBU
7fmegqfYeXegte0URGQlqwV64Gn1frcs4EJF1gZveRizBr7NueMuMWVrmFvqBVMqEg8mqj7s806p
qEROpx7ssEn/E7swJ9diITQu7YkXvwHwcTz/IgnrmjfZCkp8Q3/rCqAFQqgYwZdwasG/AB+fF+xU
61zwOypuWS2RfE+ckFfGQfrd7l3qzTrm3v7q2yosdx4SaDk0/DMMfP2pXD65XmHeaIchq//KJA0Z
gsu0C8s7BtEGb389/xSSP46pyRYZDAt4nSIivUHfB2VTwJT1BAgPLqELNIFcRtOMsc6AgsV+WpPo
THB9mB9aVQOnyZUBDgRuVzc9DiofJPrfEN0q4o6StUrgQkUwZ+kX7Qou1Dr6Z4L2miTJ6Kp0UNY4
d9EJqM26C7IegieObf1fNnspC5UhbZqdDRhVQWM5dMJc/wSFzIxbAvl4mvhM0X6VMVk95fHHG9K5
9w4YKn/JKyykNUeUjY1Hu7f9LmP1Iz3RMLEAvZ34pS0swlvCYetyLW5Nq9lKjBQOEoXMOza1qwPp
DAhy9z5QJerswj1qibMMBWTOVMJSJcjdFH/dvHO0cNzS6vr3Uy/OlFRfZY/8TVUjl7Ujt90dcAUX
Dp+w2jsaOhKFRUamW3m/EnLDYYtC6tOSsfpbjqal8KxXhadNXE1YqrkEQEwPTKcui30c2NtcQ9np
1AvxUhas5q1m96nSU9RoR8Oyl9EjvO77FEV/w9V+oO4VfExL9WjXWr1AhlVYTRflQgmIfreV6HcN
9Noh5HWqsYqCNWUReSsVvBbbhs76P5gSwbPvPEQyfa+JwEpr2ajgNyEH2R7koyo+MXlnLYSnLQ9X
xqOuShddqpO44yTLvYZmd5ouAxE208LjLIO8tL7RQCyAMI5gIxVTHNDxpRV7v6ZwLwS0a2OY68up
6ipgK34tc/fxPA/fAB+TUFxwh/DvFXT2RaUZ715+Re3LC69scciry2MBWWocvLhnVCbND8Nmf2bP
liPzWYLxAnnInS7sqLm7nVpOBu9EemqUc7EYBbFT6WqEi2R013Bti8vDN5st75hOnMyj2O0RGhZ6
Sm/g6nH+Lj+TBpkUbVO4tuzpTmuU9FQMSB0tCT9+u4OBq1Fu41fJ31C0RS5qTiP6iaZtUDdsR5eq
OzbekV6P1oM4D2JYHd13RBwuxJ9Nto8zQJJe85H4SihGFu7qlCvW+UIOs04MiVAFZ8wexX8pgJLW
pg3tiApb0ab3yGCa+FCq/7NufNyxQJIapYpTJscVQ+hb17rsp15dY8MOVxV3mTpDN1NzcSsNnKap
KO272hByGnASt0WmGA8q1jQZuPOZpntjtqwj1y4fzP7MN31Se0O66e9h4scrW4X/7z9e1mdKjJD8
ljF8ECoseJvwSPgQUXO7020gQ5535gIk7qd5HnalV0VWyih+0xTD9aglXTUSjxS1dX/E45uOk1J/
KofYKGxFafbPsYkggj7bYPbRb+wN/rOGGpIdNehd4zdrRpnKugyf1Bptnhosn4At4qOZFzkAUpi6
gJWcUipHedBGRcRyOZFlyZjPooby6o+tDcGVvEjM/hOfWTGcZISj4wvjcpLCYZqfk+Eb9ah975gi
9Bm6hF17uFEUGIePKheFXgVV4lGReT9zZnORvnIVJLHNxy0s5Yut4dktkNizH4mFxZn/e7gcASLj
Ms9wESod08qyvpQyJVJwc1kW/BICeuObSpBw0vqOKlwwg7kMo82nawOyyaoYadEEeZCGmQfV61Nd
FfB32LHVxX3ya1RjOz2KxnyavdQj26YOk9bltZzFhrxpWLkIqameayPm88u8FXNSrpzevykm0nhb
PApMJ3+DVYZlmSlh48HOZx1mSewSTgXPenKdwC/i/TfpYHH2D7n1nkXac5rZbJMRMlBPAyPLxzlk
Svu6Te9emV+oP+1zxDxLOfywPe95sz6uVpIPAI7OjsL127TFD4pcesA4LkojrgjAud6bGsCYbTme
dvJYdY1y+PoWA9xxFWEaen5fAbvP97w1QZklGv5G77RKVw9ERa8Y0wom5zI3tbAakhirdrNcouZG
l/amWTlKq8h6gdLsZPBnPV1KoXbfC6FAdrRB62Cyxxk/Y6H7t0sSdSvseP+IQKVp2qhXYN4y+w+m
E6ugIT38Gru5UJWwikBf9I5Day90qdE+qcTLGTxZ/EACNsLTMfELUTC+UBp5R45IVRvSAdr/Pd2k
fbqWxQjca5UIb2rpOsCiVt8HEU1hZpfZ+XwS3ymx9DmqAxgb0UASLMPoXC0sNdzLMd8YMeqRNqeA
xn9b1t/4H7XjlVWzW6fb1HhH6NrBdeXVBizV/iOfJtHghHlthH2EWhuixTignxPR5ilmqL0uT+Jv
L/e4bY+C+23dkNdDe9JSXkuf8nggoPXp9aL0LpJL8GuroA1uIMhi6gKBxsz7SrwuEhs0BcANVlWJ
9H4P0QAD0tnSHKrp0MQvot52EFOreR870mN/5uscbBSXivDBN9PFdTN3gWCRz7aIwKyI4rsHSWCs
DIisvh554oGmvrEHFgWaYnwsXiuhhJpI8xLyqp7aDlkVgELkNM6n85zjUFqpRIRjs3StZM1Iafya
PjtY70YJ8Fyl1vLJeNXsOmjXYPE+1PAKJShnWS2cP428vsdcHszdAQsj60jpoJjWSlwc4ac4T8F6
JPDE9DSxNArMtYSifCiu+sNb3SgMzWv1S2UZ3FTqAb3fCUmmnuf2HuiSCPo1x/dIDmWFbwBY/xaw
oqrf8+uFuPIGCIrg/8af1IkYC9E5UqaH1tSV9DnCGTk+K+kU1AAwygd4UFiVoLrPbNygxsnkTEXx
JCNw6uG4IAqdBdBwsxyMV56LpvDH8auKbE1F4Oqw2F4/B9+n0vftG9cUlpU2Fm2uobJyX3c0asq4
wZUzv/MEdqqRdcTQ9h95ciy7Y2Y0JXMwWpzwNJus5bmfSEuGsSlM7hTRsyUTMxXMKzCsUPaMf1dL
QHmrOagvKlRgy61BJFyh5F30E2S12U6qJt2/euR/nHroZ+0chH2gLmk7t0AMbuKxH1cLrABIDJdQ
WTdSvUljo8VTtb/rSEMcjQuHw4xVQt8qTe/2CzCnrC0mVzy59GedxDj4ZzEUDLQCcw6kdKC9XgzO
bAsVnezurdqoT0WevRL/7zHUYajwE1a9b8FdXhHAuLAAPEfDHT0Xhw7HfG3yNWyEUWU1062z+a/K
ZcNcUak0lmOTzYV4/E1U/S+JLkE6CGJCqukmxRzued1tJBNRePqn9vyHqmbAm+UA7h8IHG82euOA
95sZViq9hEHDD1rqeqRYOTMemp8lsmr4xzXxtW1+7a5oNvVGwWKT4IsU3//5XBbeBEDSglNNYz6j
+FqsURGpoNFFoTWZEywGe+lby2rRz6cIqaP+3buRqdD8CP3kMuZIbBgds6UxZCZkUs54bIsFyeT3
YY1RsUd69eYt0RL1hlTWDP9zYqNoja+mmuClY86rq2izJcfKFFTfjmZGKk/FKWyih1LVnNt1f/2d
xw6AzwG3Hrn04wdjhwgImmc+Ly3moWMWx4MK+AL3w+yZUwTwo/kvgT5sxQPdAjSOYDpyjGc5YnG+
8L522TU1YP1nxHYcJYns567grMmIIe9G/R8gW6stBaFLu920alYbLGF7Pqkx1X6iDQRhn15jp4QA
h+0uhFZB/AuS3sh6U7PDeCAHnghQc2GOjLBp50aq40jlIun1lahJ0S8KaAqrYLjYC7q00ZpSp9/O
lKcR+Vrr1PohlfUR4I5uD3mgEgoHnRjON5KUmm2MQy0JHkXsZ9Kv/QVQIrLDeNh0ulYOsht3HAc0
NG6OxgQ7eDCx19b8TXK04KpFQwQYwiaSHZV0XtuJIcvtZYlXMam5y0vTMAwcX5geGOnOVzVcKa2f
+3IoXKkNCW1U1BO21PRLSHt3Jqp1zfnRnrWEGq4bxo3naxQFQHFZv6aA9IDJo3UID/V+hekrXmee
vMxA1KT2vdQO3yJCNLvEW/xsQFR2KWz+W3RQHdoF/NeDfc9zYYm8U9QDOhZRG4/vTm0IlNXryCH9
l/r7NbZwgCUDNtaNXOwhwb7MfrlnonHqUXsPlr8moxBBjro6aHGZAId9hWEeCtrY6/r4+pB60xtX
0ubU1WN/AKMJRxACj8mcoIpLWbxwuklMUbIEn97IExhM4xWKnmnKHCvHcMdgTb+S9M9k2OxGnZcf
MGzP1oP53jOGDVzOj26k54I4tccuLZ/amgsC2+kZ7Ae36veJ30nvQhqVN3p2l1l44okU4K9abh8+
YzNoEAj4Sl7Hs9Z584AoGZ32Qgj1GDvu7BOvRzDXz0b6zpKRBbFYiDX+m678uqj4gobNG6repdMX
sbHS4UYWa9xjCFfFqJjYoYCTG2mas7pWP876D3iR8hWiPnKRTYMWWOUW9tFz1Cnd2/asIX9e3Lap
/zRc9FMmuUwJP1wVENIRuOkQKk8CEqzdWhzAoPO/1depE8RFXxTEV9lK3ysmLQWBolFk42rKlRTO
Io6+s0jw1i8xEd4JSfabl8AqmnCEmhD8cwRnVfXpy/xdNtRyvZOQ8hG2qiP2YIlho8ZhSaxMae9T
BK8MrIfnSnVrLOYZhzhptrDg8+0WZCHLRnXyTEqY8i4VzudFHuUeFYFNB96IRq/obL7ALcuwiUq1
JXOAJtdOL8Z91YU2elc8/ZsxybdzpZwfVegLz3p+vzkmFp3NmbVannr3xKlAG8K/4L+rY+gEA/MM
h2RL5gW59+qfImgPDb30LHlivAudVvY/jyIVzLqc1S75UkBt7RHPqM6vs5Orwsux/gRH8ANQ96vW
5Xf08LDZAUm/mxbO5Jdvk8uwB5aW2vEuZXqGbrgwD/LbQIDYg4sfMGbpdxQBQSvLGRVUMxj0+krW
VF3cDCc5+bY1kLqtS77dW/ev778zrv39fJGNjis9Xs7+0hjvvc29Ooh4RgUcLPPFklpijpighahh
yZTr2Rpc92g3j9FVhqUBDXMNon7Y/kMOporOwUGfyCx8LQtshfHhbQj1/hIZcSDU1H+otZv/JuPb
PmnJ18dk/okV+h8pFORXi7+M1HVXPanqc6Uh6alkQqHbKqe5jBRNV2TAOXwKUm2PcZrQxXtBrTLX
m7rcsFhqjC/CJ2Q2kUR34gUJaHUogHA8eZlROZ0z41mNyzCAcaxHmXZttn5Umevy7Sqa+kijk3qf
RhDAeFojITNtEgq2kAJUDCSTtPGliqnM0vcCfBHulfu2UzNbF3rdyd5Gy9lJkwetkxGRhJ4m7iPV
Yk5PcweX9N0BGG+1h4kkh+wTlQVkEMno+oHT9rSMV8Rm4+5tTb077JcBPIP3UwKiiHlbs51RuvkB
ZRZO0jxmKWIDaCa0HlIiA5tSayMnA+ypWR+WLulSKx0WcDFyMKVAOMfx6Jbwd2MxETK1oVgs+lQq
jVNmLgHSecXlVRKJ3MYggydQZxxIlTdzyvn8bQXdZCyDj5J1Vl0GYW0KF8yuSJJfZo14PasiRr2e
dqt+TKpd9sIMgvA8YaVPdT29xyPm6h2FJKmWMGdkwpTNjDLybYN3eaSj16Tl6fVBoonNmZZdrTlZ
okP8kYKslnTxmzahCyBhlti2aBbh3d2pTZzUho4jlqDKBEL88zoXZn5l8XDKwbNqcXb57OCfECFy
pTONTo1KHHMH1yjyJ8vBt4KlPxc4Q/y5U9xj5DF2u1h9zDjwU6n2CC7G0Downr9h47J1IEq8Ffs8
w9DjbD3Mc68stmEfsOgajthyoi2EdemuHdgUPGkbj9Pd4Tn9E6FwZfkqsLyqYL0AUUn7+outXGnN
helpovjMPFdof7IpEpBb6M4JeI+hJGBUgdTPedDIKuEONlVWuPd4g9ZBxStPs8KL42O+wfUNImE7
DJAIrXd4YOjWn0QtRyV2R0HIfmCjO8P8OtwJMdwlXdt0npL4oXRmQAQaodP4VTW7Zk6YtZQTJFZC
pc29peAW1/AC/Mjix4o5PZNHLQ3hzp+hvOaZF6cFmPX1I8jh1KCLaxKCJSGxLLuLQ8qkWYTtpmsd
qi3U5ozUtrasUWyhqLzaHnKgAG6+xw5pURwpPnPEccdpZKxyA/prxcueUND49F8VZpV9WosOIajV
kEGkJrxWWtcpcvJoRgX//vCERKCuI+Ij4oc02U9xzLqCgXFrkA4osLgX0YnhwtYgNXluewdG1ae8
O4o9ZS95+iunhhZzuqfp2F9+yCB0HVrvzWIC22YR9LfnyAcmQEEcr5ta3942zHvXB25z8kyVMHIL
tDAb7r/4s/gMO1E4q2k9yMHMg53UY0/eMOaU+2jOR0W90UrupHj0cuvaSWy0WqT4BvXy8hpsseu9
DQOvLbL6ZnUJ8qzqSB4gQCE5EiocHu5bJISH6QBZtLa9ZbjQmcCmpZk2X3raofUerhYbrCKFDBXg
CPAeDZdgJrfo6Y+VHO3dDWSg58TBetWxAf7Z1Yi96ru4iRcFNKlTVjI/6zujC4fBOjW6on1xbeqG
OZID83QIAhPDToTA0rLhUNitEqccQv4PkKajKOirYy4k4R4jcxgmEkbHQdlDBXw0497WC9gR/XjX
zwug72bryH4tmdVZ/FNOmRUoi4kA7JLejgMm6QSRTbfokAGsDSARz3la0B9iCLOEJDIU9fI1jwLc
Ny81tFm1kzBk/dt4K+6es5aw3ULa3SmyMHN3MHHmWpUy1B10xFP6v+z2W7DE1echPgcn2odBW7VI
5oQXJ/URsOrZWsLV7uq3mFUbLCG7Or6g6dv5/KZjZTfVUvhqdsJ44wZ96TIGVTvXH4wWhRm3Anqc
syO4gxhtlR6bimqUps+vEYxDSPWtajyxTUWPLE2CffKcEH8XRmO+UwcVRAd6MGzpYIOEhkFe5pvk
/OYaJvPd+cYqUEybXku31V0jh0+rPU3ry2+omWImrhTv7nvlKnx48McoyUtf6t5kkklMyvOzDWp6
YeuP8x3xoOlq60dec5OSGZguM4RBfGCKX065rYhPVmOfpGl9lDM0iZwVpdiCTF9eR2Rs1PkGHBjK
7Z8MQB/5jqq8Xi7Mq0sU287MjJwjPB/KmfDDKuKXtJiMjDpGFMFC/Ig5+31SgAgdR/PCSRBpfyhp
+TiFx2XDixHXLsBx7p+13RnGzx0895d1uTyexp9/x8vsZ4JeXnYinq11nQZkzJQLArgNe/uhWNVC
ucm6qh5X40E91cEs0wtxvdMEUq4RCCHIgAvhZtTtrq3FNfajJcrR1GJ5cN5KBy1+UMVUyryumgYg
AV/KpuVkqZd4dDyjSA8lAt9H7rj6gGGQRmG56TfH/KUKOAjM/79eqUfUMBmORWAbMqTA9Jap1VvX
ejnsaWrB1/yt2dE7gpX1vNOEkjhhQ3HxXOxhEax+bOQ0AXr7ZYbQdF4+QUvbBt921innyLckSo0O
Fkm4cUziuYRcU6anmII0KFgLeB5StsSxn6hjL20UY6WABcXUzveIv56MySIo61CM4L4gH9euQUpi
AmyG6zMy03iMkukAaKCC+Rwki+dKPbaH9hCe3B8Wlk4yShIAgJ+Hvl8XLAe5OOHw6CvEUBEYCdXF
qVpH/sZXcaaXTUx3Y+Xdse9C5uPjVbaaKuz+baekwMyDtR6TaE8Ji1SOlliChRpPHVZHEzSUKXbk
qupZn2XPCwKvHHXrJ5gKFKzCbaOyCOAYMdKL7UezXLTUy6+oyZRgUWdzg/zJAUnUJruxoc1it9U3
qkHxb4E1baoV15wrS553P3wi47qqamRht9SS9vlTbBofvU+iiWfIbYX0DtYYELSrMlzKAtlqXq9K
83qc/+SJRojF5n4N/DWlelclwO3UoZZHognp/0qWJvN0ftMxvdT+OowPUzUWZ8I5PNJdsMkLUUWE
NbY6RA8Y7KbevamRYLeXI6EOEABkfbnaokjA5EDrri4BW+WG2gYN0ozAG4x5b3+kbmwgFijCANBK
8sbrIyy/ZSy4kIBgwPSBgEEONvNPtyy0XbxBGIpFEtX88LsLlU5F73dEg0PHDiYOEvFLUrcGKEtl
VY7HUmtGXuk+pLMAH05/YlYLRxezawV/uwS50jVcwtgwS0DeSPmOyXmCKwWEtSbc0mo43Djuu2Jp
iFFNfN3fSqLDWblS4N0VcEkpXmjamLsUFYrn/0PD83d7SqKxQ1LVfoJpdJweUm59bNYP/j+jQX12
V0JnRR+w9Ovq44Zxr8iiwsa2CJyqtsvi+ljDFWfWyHvOajD3BH3gfIMN7nJPV++OzH/IBrLkLRS9
vBN/m58zPvoyY5hsfVVWgIk/rwV7jiBo4ibohF+RpLWQtCt2Be9iASfSb2CIWWhJzEk2mI4BkaPv
CKNUHAwOXTGr6/Sz5TqLS4W8XzHPmMOPJtwncbfPa5pgL9KSMQtuhzkhX+8Klvg+aVUehYkfeM2o
5fs5iqQiSVNGT1J9xLfBhMHhhgYPi+d7qQc57DKMCeFg663zGAzmYWsX1kJMDf6dqen0SXBp+ugS
QjVP+f7Jn5ljSslP1XPnWMPyX5f5QSERs2x1o1PtvCCDA7V5XTQclO6Nek6re0OCRSs25WU3fScJ
TQEx0JeuJc80JoAxSAWny6d+OFY1vjwCMKwTfoaLp/1csfhp8oBvVbiIulWF8VeSmNbcsUPaWbt+
gsg9qRv7nES+kwlRHlpzstEEo8oqbCLxk0BraKTGWHmwynXiQk3dYhEwMDoc7o1Vl7lmCcXgOy+8
eF1KYcTIdy0cP8ERELo9AedNloYta6kkqdLcFY1QLzUg/WF51TryKcNXY1yxb6lAvC9SWsDYM7Cf
oGEXOTpfXIEeV9fubijosT3/9Vxbd/oMlTqgU7101YqI+4wNtZZRNT6QHWg0W/ukYhpGK54/U+YA
PydoZ4/4LgJQvnxhXllMHFqxXaTedp4Cj9Oe8A8uGyrur3CI+Kmp5iHcTos9EAs5tdhluEoy/2eF
tM3te+qNV3qrwTA+/NXYadg1Yi3O6mmzv3/A97sdOWvM07O8b+M67zWEpsWZeMVUBuipk8CtjDjZ
0sueszQjNcqKYEwWZuscFaj+4SrqpHIhJwdFRso3Npahxyd09fOgxeSnH8g4Ru5JOEprMQfoDRwR
wDcCPPiLvijFoRB1FiwwxqQuwU2q9kQR/Accd07nF6smZ+peYrslbkn2TjwWpKc6OjyAKuEXTzVs
swZRwuUq14xkG3ZPow+613zH+UzAtKXoLUwTPi158/6IIAxpZ4BbnfoKazQNcJOgJpKvjuWe/XA4
M5Ss+2RiKYGaCC0YtHQEHovCc3jn5wPsY4g3rW8mvwWTTaEmm9LYrSEYxtQ5PN8aCL8CbJa4gnSy
qhgvg0bjl+ESF2dBZI+1AvvRss+iqyz7sOtM1TVhSw41Y/F5zg/iIAD39ZV31/1SYaw4LsShAVAW
fuQR3Yy08L25nNDcNGXpgNM43HdwLK1RrE1s7RVw+tCMoTMqRK6BHaYI9P2EtraTbJr5Y8vZybwl
US6RUNKDznpDfmGHllS7W24uIwHJiHXfLETUUbJPtS/WQz7kIemY9RgApR7FmQn95BeqXp17uN3i
uiCQntEaXxWBcUv6uUYbMAiJacA+8MibL1FtMsjc+Rh2BGtEr904d7OB8YXKX1u2y8upik6DUwI+
UQumCE5GZpzEx1ZZAOgOOWq8e2jP/lkq+y5PRZMeTnS4T5qFbVX02tyamYA3YLpVIhgwP8HfBqKe
FP2k0JN58fwzXe523vBNJNalGJlb3Wl42yN5Dw3J43OO3v/alcum/QxAg7JAEUDEDZKQVDRv+0Hq
yMqU6lYArGpKgBH6DZafLIJVMyGRSX2dbw+w7n0v1fw4d0ZdoiYREnckYrsb8WHrw+0XgKaayhSM
VM4aARNkrYHv2FNT7tCSzAVjGr2Gje8ci10Zzhttrebp+JZUGtcFGhemdP+3dV9l+ZFp7Y7AeovW
YzNVfT3MKh/lv1BOKCGeGHP3DWDXJG/tODVg3HxYR4JEj6ZwXlYtABEdoIdVEU5ac884S5REzgY5
4L9W9H8N3Lgxmmbozls+3hhaqCd0KW4AztP11UjltNX6ISCax4WwLm2XXp/EOKzxoxMoBGnoSs9z
AC3suYr88RJxqWIB2wcfS4FQPRp/Ad1j2R2s0/yURDOnEQGW3Q/mdhslHybVuzQbTcDFQ4AfZfOc
60T7kQIOC9eOF/V6Nf9Ams/tyxRHgEDqA31ylKd2ZqvVsuKdl1v11b3T0fP/4qmjQCg7e3Wr+ClU
50Xke627JOSH0kcIkzd5DGtfwmdO941viGVXMG45juxH1dY6ajI6yurW8pyJ27bMNbTl+WQ5Vtpb
LQ3oy8BL5uZ5sidfvL9ai3+axPsEe/XHfnIXHEAGcuNykttkZTrjR/oVKFpe0sAvaAeQSGfVInbu
KGjAyf3UUKL8io0Nn1Cz5k4SkBGN9cM+p31k3eYmnISkZAnS031kxzJoODpRw3b+EPX6ymg9jIOV
HcfPnFrZTy1SRUkEKwj6BTR3rYo4KbB20017DgXNLL1viYwYxsWu25HdEWHJpRGBcTth2sdDrDSF
RgjTSNvYR7Letgp95O6IkD6P206PrPtUw+T1foCPqNS0nhY4VFX2Vg6VipeWSYdzHR24sslJV+RX
UiwF2/l4xUIpmzT+ctCAryd1JE000hKNTW5nDeP/wQuxzfjlvUXdJknhoOIYjeizfpW0lBfR6le3
SSLhT4KekFRBiXVmqZ+FlxIJAT82VGC8yS0P0iZqkaS9+yt6H1gaWUoy94TrsfUoYg8OCFDGFRZB
y14FxIteYlQASbueloVgtiFrBgrSFhBPo/EbloswRLUj+lXYgQTkNng3e/obwdMRxLmHF+1Jhcw9
PPpfXIt+UCXB5ZMLdW83S5aB9t9AuhqsJx9dC8ojkgcEJY8QN0EJ3ibKL6CbbJoGbpcX79OKbA/q
/Oyke/haBAEVRBcDEwsLLweOF1We8REk0ZpsqAawRbea9IxmMiZCrQ6SYUha8UQvb0b16BEsJWsm
DQc2XTDyuJ3cB0f3Xw7EUwpfh6QDNalXi3y0Yvvum/76Ze7c4/691kDVLXIHbdt7V0JaRSN+8+nH
csbRt5eaffJHpnTDXnGT/O4t2xT1MYgd2rz1/5OfjVitOdpnwB3u9Tzzkdb9ws/7NQsMKZQT9wU3
ak88TBH7tfRwUb6z3f6ff9h/SKGAn0NkS7bAhHSPla79B9Ou427le+jEYw1h7CfPJkBGhzhyXVA1
fqH0xrCBC2JO9OK2E0Q4S0j/jWx1iMGOVJQ8KvjG5znDFp9nCWyMHc3jky5bquYK4ICLnwaJ+4Ni
UXDisV1BA3chxThazligFIgpJc94cBjKAD5EoWlTuUHvFSHh4kU7RYmzDxUls8isjj1goi2NrptH
u06ZISQK70Uwix1EF7uKDh1JHvQYK2gmFfJbeLeuXsuPNUUz6/ShpdANpEUtpSJpynuR6giwPKhI
fUOxYE7I1ZxkaOGVaRX872DVpVnFFXvRM05BLYT9BcWM5C3/zfTuHBBGATw05c3EYVAfx1DFx2KK
beAorWOOUn0MHJdUSU8QaJgHob4FJmNtTyyVe76HIlMgwc2pYIL0EpMOlG4vfvLPyLtqreWMS54Y
vfZkT62TfZYEkLmEID+XEoozCFcaAKMwoajY405JQRdPFxHskDVIrziaJRxbKQM82NYgzGSK5vWS
9EW15QUUX2NZlaKaZEW5akfpFCuWf4PS6fQ4ciiZOYyDnmXl9OSx3GITBu2kZw9kYJIv6/6dZMcI
ATYrLt9C19uN8hLAVFFal1Y8i9U4+et3GyZwVLWwRtTqIoEQFG1OgqxFT+Uv+yh1LPqWtmLUMdGK
JHzoqFGQulrMYpaFL69zUj4NWtN6mqNgnhioqRqhGcPPvJd9tOA7fKGVx1C1u+X3Bw5vfumAji0u
8SvoGNI1hKypJw7mFk5/vi2eWvTS+N8P1H0o6cGeszKbFCnz33c3d2Vb9ucq0aRaoMwYvS8lxcQH
cYgtNEt0GjwKoRnMONJ9eMdRHrjHQqDg52VD+ZikqGMuq8Yt3Ou7dk6X11rte2fhCb+qt6gQfBDn
aQFTMPMwwPdxuhP0OrlJx/J/mf3gaIpYY/AVtQ+/H1HqF5EbQWeWf/djommcQr42QW9dw6zGjMfx
c65PoZiKCQcqGK6fCYvnRS6Qpa1/zIuKDabgpOxjSZxlv+jY+sVHRvA1HDr6b+80ZTWDW/+BCgXb
dANZz/wh/lWPjMWvpIp/kvYP5ItpAsWW4r6Z6A5d+/EIF39hmuXnpaz3G+yOYkREI69rUymAVV4u
ePyB/XEqxFfKEOqqtaqFETZ5cVyDob8kNMh0wvVYS4dOh5AIg6sbV3GA+FfGVKsBW8gVmhJCjJ5a
ZJvuGEMpOhCfHpt+LL9Coa4BvQ+MSEVZfyaDYsvkGJyCUJcwsBgOm6f1gJemSpWbG5iuWOPssuJW
2nG6tfpuvn0SIH1daJ/ULT2Y9S6Rkkr7a7l3M0voHjMVg6Li638rWBwZ8AVDyVUw82dgyU8DvpK6
WJwSw1dzCVRg00UZZd25ztCruzQQ04HZH4But0D8vDDhBg1nA9aKfyRQkO1/9+k2ymN2owMaOU+l
KOuQhEjZDkfvCTKvydFc8/n5jQmw5FQOva4lbnP8IMy8DX8n3M1NsRaAOYz96qn9pLreeuNfDHn+
m7yCV1HkA8jLkjEmFd9QqKY8pCozYkIPMhVAbjFSoetP0/RxLs3ctT3cwVOMpzgbGDN8d7blKZXQ
OyaPnWe0nCAIoowDmkuioecRMBr56Ctt/Wif48g7oTnBNyf6MdGwnw8xSBcMipBB+7zteJ7pMN33
y9c02GOUVZMQAvW9mX096LzjkwhQ9b4d1rgOnpQXt1u5cjKP2A74dB9gU5en+eoo2jSJGmwDyh4e
YHm7gFoHLlRWpKoU6NFc4V4HcMB2GTM6QXknA0Yr49eZefvW/o+UiGgg5ttt93+NQEPDtciDWWCU
jhf2GWulSDIENxLZe7E+uijB9pTKnjQS3HunQqNCJusv7b5G7ojbyOZeAN027c1RWohUiNooHARP
QcFpK+NM1GyMVqOrEJFlfQG+3X7WdqOYtyDIDpdxP7Jq5kE5BbxSVHotWLoyGjHsrpMe0Trvp+MB
oA/FYpRswm+qBoOXxZR5ZcWL5LlhdKf+24lPLR1gkRLB34iBvyvSqiG7ZSYkbFwfYaOl2r6hGFPv
v8qZ4ed3O1TgNpWr/vbdtHHd4u41SE7LBICWco7c6QsT1vD/oxnTxFQHPoHg2v49VQ22BxifC3wh
1XYHoUNpqQyD/8VvL+6M1q4qn1p0q/RNSULFURdMIulbc8P+FfR20jRBT3AWa7rJiTY3N08XOOBM
K5cNqx/tMrrgdhb8OZ4HWXWq2YWA6h06XnaJ1fYQy5LtGXZo91AxYpJXIj4AHaOcgUQNF5PsqeLn
132j99ytvm9KX0IuqJqCZH1ZIPfOIbbOxCh59CSR5DD9c8itM1v/5o1Qiu/Kou2lBTS0sOJn1kg3
kIHsTls+rgdf9aQ6WXnVjtJdaiBnhqXPSW69k54G6MzChCvaS4XIp5gG1+bUONtBWP6BGnNTSNEg
zHd5zStszQ/yI7kcjxNqkrz8l8yVINrn9LirtAILYZXgCihewZOL1TuXe23JqnLgZ6ycpr0mtqBa
QUexmxAXZ7WzE+4zZ5c+lcXvf2sdGWuWVHEe4OSkAoavpn1YfsrcueoQjOq4Zw428LIjAyL1XXiG
kDPbCEcS1cWpFhZklqt1QunXH2G7oTuWMpXzn97PfDzGaOv8pxtNhkKOZ0w3Hw45LG0M1VnKylFK
MAMmZIbSPtlo8hmn2hh9n6uBwZgvQ6iHh99XInhtos6LNFpD4N5j/7GF8Z3X6JVzxWLFiFbEg7Gu
eF5eF2u5JxpV+5K10LCIuYx42jR+/Il1Y/QOO9bjuES95c9Utx0WuX0eUmT3DfNBaoYexp9ibkk5
eW2fIW3IzCkbYS+juHAfSma4PAVxQCJZ4lmSYmxxfugIzwRUlIUCO6bT0qJP7CvOAwXQ7IYLf11e
PXsQ9qvRZB4N6ZKOSwhg5VUMcvxFBFju8ZGbs0AlmoMca3vIEh445tgBfgzVXW4Z3b252k9FgqP2
Bpjyb+iuLv0AZq2FRFRD7UEyLi4/iGO7A3E3p7/4agq6lVOa6ZXvO7jG6l2ybXlJXClULefguYmC
CXZitDboA+msN+Kb7HkBvAe8GNbSmo08v/9D7kUvsiH0rlXin6ZZgqUjXeHYrpQIMV0OMgTyO8c+
zOQCRsOXvTFxSn3DaxnY0YGDfP29/Mzuk39WhklkgXGvoN27fK50LQ7F1G3i9yLHI8c/qfpKyZb8
ya1evhpYKRIfRS03mFvCuQbUtswzF+t9cZ3ZMKouSLK3aTklOT4UGVaTgi3KzJ6n9K82Y9+Rch9i
0BXFgwMcsTJwUhlk3RdMtgXAOc/gOkQ9wjQ4iPNpVORPD9Vx0A5thjwZxU0yHLuBi0u/e7JcnGZR
9yRczs6RMrJQcgdGXh0ndky3BQP3xs0K22tJNLG7gXT9826PNavsjwcDmBwM4Cz7NqSZMxj+7vET
98lAcmjKdeXpmosLEJLrpp2yqChp0cjVfTz3IyfTfSimr6Jms6CIMRBwHMsMbNjef7QxmKGPTR9Q
DH2C7NOEqESaVymb/KyRWi9xiqz6l6wtU694HgT6ROtFgdVvzy+1qx/gB6ISTLjNFeXXrqCQXRoA
KyQ5uu3wy9MTogJfr5kML79cIIdXNzBIEUR1GqOpf//eo89oUhmxIQWcH7fHCFBj5Yo6qIfoA+2P
Xn79/6Ztb1iBttIIMytiUgxfHvkSBMA9p9SKSpifce3lZZj1r7nDKxAesFPheyXCWlMuwu5bOTMS
c1LRPVhx9NUJQB2DfmBv84wcV5VCplW9YzbVMWKqpCQ/29HcL5q9JAXqR/+MnTaSJPPZY9qYmL/W
sMxp0HKHTNs3wbLqKY5RakRir80SZPGOBzCdl/yAI8QvZeXoecTTjOgO1KpFDFdrOUuQkEuDk6+y
ubw5RwWEYuSpEXgqo+p25nY4d1+C9egfHqVsqkT64gdHK8W0WpQj2BtlGz3VP5la7cpXHR9jRVEe
z1Mk91M3G1f4uWBe+RGGZ4ZrDHdsmvcMAfhAQBsuoUGORscfBwWJfHtzsnSkpId2pTMUosdhVwrk
EPtfJyQZeTJhq3xBRMUkOocEIumcAjqeR3/awNN+yF0kJAKtmYfr4tIOiwjHrxtk0gNJ/0HDEFBi
tpPmpmw8LK3ekJwQbOLWb9/2TC8/dGtGKAk3jCKbG/miCxVHHzN54sJlIhv7Ih68fJC7zZEpIymn
sSmfo3q8tU+ljVALKgML3MujJSi/EZg2YKHM7GTJMWCFeuh8dRxF51EFjkobs235upluK0IQfdR6
iLRPXSYdhN4XagU/wmuPYSAqIluHftMkx6qlD1f+D9Gm7fFTxOFgybeWRcr/B0mOuRiE0yL52lg7
i/cs4OPKhPj38klvBW9Mk4KNyFrFfUJ/4+anmnHYP7iwjKa6l4AgfbImZ+bKAeJp+zKh3rFVnPFn
QvlvWep3G2Kc60BwzTWZL5bNvV0CB2ohUvw1Mca8waPZWvNcbN18LJ+/S3svzYggWtOkI/oo45rw
r2JFASnyLuT/bxtpiUrM2Bbm9oUr/danwCC41QNU8cvns8kP/r82BiHOd0X4kwtQ7hvMEFcY6FZk
24XjmquN2grAuUDyXHO8BRzX8ZXs3QtTGM6vGejurTEXC047bPD2cipsG0wNEf1veL50oEnpwyVQ
YAn9rOXLCYmWEM8YXZvaBKZrWcNJ9UUmC9sCImrlSng6p9getgTgdnWF6jf4FWjUpSkaCmSu+pOD
aF2GqgvgbcoxYlyCt+dH5q+WfHmZF460QHc3AqB2iepcWJugTazV4m+LGbcLmXpQCfe8OX0gjwev
+bQmG0l4F2GY/UcErizZWlBIbAJ8Fxm5mEp5VVT1Qos4xIGa89ic8PSCPXkDmm59z+qtopxYc7x1
igFBfb+zPipLjBauAyy50NyhHpaptem4Nl+/C3SDn5VFszffVpjGQn4OMXnZxdH81Hc1n9oSZzLO
TfBPNcigp52Rpq2VIrjiGXu2XrxZqOxNkE/tu0jQl8VM7XXHFqtAynjNsSBTXXTBbrJjZw52jHLa
w5cT8+HejpqlJYdeanqDglrHBZVntYGJJqZoB1D8BP2ms/7Llw/s7IvGG1gEAxxqozJt65xOPF2D
9HAWOtuuhCJJjM+8szE6Cvs7r6XPizoPmLPc8rEPwZ8L3FyTj/vTxodNJez8IO3DhzctwO99Sn6L
Xq7HtNiq1GyECtfwc5UKhugJAiNojjrE20/wZYQg+DO+ISMuK8fSm66Xxm6LuD0Ck07WlxvEwE/G
paF4zkTybBzzsFNMXFtTWQ/lOfg11sILcao60usn00QXfHi/j7E7FcWFwffUDhBkqBnlxwJe2/zS
yitvEHuI8V7a6aRQP0nzMshxdLw0mvvlOJttzrBJGJH9FVUsyQpHxOMY8Cnb6iNLP4eX4JrDOL2S
DujGKL9qplgmGoLUGmZd9PMGj1QyShQAN6rKweD9aNVreVsZKb77bLG4GxhDzILv9uBCQmB6YWME
8caPcoKmMJkLI5rjSLmtzuMi+QUpKf6+4z52RYH3NlSA/LMxyEgymglWlCWwE6i7RglOoRBEGiij
YeIxYy/ekzaMNhH+Y5CCxAX0BScPDumTDJTQ7njomNMuJsY9bxsUkJ3S0/hUVCXT3jfaOeCIcQPk
M0EqMQaPs4oSn/07G+PdssoK3l3OhmCIa/0R6k4P3Txrm28aAElZvT4iapxivdZIAOViu7qzca3R
r4M+WxjAB5yIr19brrb1dg/36XsDcZQ7Z3VrrXpMWB6mbXXSQde7tYVKn8qLOuyWzY3zS5BT/5iv
Cj9npyq1DPVLd9M+ay4Ln4Gb9wJQltLeLGG21yRJYEcn+M2IVc2E+j2Vpa+mDjTaz52NQ79QuXjK
xC7oLRRxWkTqcwKq2MoaROFnCWEhR7qrd0zYPI6CWTvJz1Yv2VJjegO+iJEsNQyar5aiwe7E6G+z
QeOG+3z1EF8UNVzm0oq4TCENoj6gdYbFGmvbRxXMeanoAHIXjkdEPLqEhqzHhLN0VrDC/GG7KufZ
MgEgcB4lKPii1znEVPiHEsAkDNbKIEzsK5a4fqgrQFJy2FMeeu1oP9+M2kzgK1GV3YZMCWIuNLkK
2ZlO6QcafVFRZacjiMiif0WMYgK9AaD+1qheivI4RM/w8DhwacQY4A6iJEWwwicXDY3/lZX/DTdy
l3wmnI35xEg+lOUJzUUq/y6v8hLZ6HXied0RKH3FAfVFZDsDVX1AUMeESyUjQ9m+ZaA0/tZXqBAk
7lu8Pvq7f/NCYY7BlKkT/vW1LT/OoJuOUCkgVVNAY3yDphhofRRgqMxIArcWZmI0Hjn2TH4iVYoe
96GbmEEm2qxKw6kyoUlIlIKpF4WoP0DDqsM4nHKIOG10hdy03zP2bEXRvtoT6Tu7s2hBZZltJTpU
TlvC9vB7VgPkXfNhJPKgEnUMguIM3BVEJ9BMiMyE1fNEn4xboUqJH0i48SVtVBFcRKQMGLNM42VE
Ng0J+NqNS5kXWq39tqXxaY0QQwWkjeLg7QQjFZK4575JeaTFcXo3nnkCYyBEgM5ubwdBiY4BiBVa
PV70FNZ97tH1NbzE7667Kjt207jZ+MU6haY086PKH8NkotuCgRCXfI3rgXpfMVWRH+MID7CO2MdZ
5BQh5jekhzZM1s+U/KnRZkJ6FzP9U/msnahQOK0h9uLwoeO16A1hePk6km7nPzU5HOT6BRN2L8W6
xXECiksJucmR6eZep1g1D2gPoYOx0LsU3DfDAp6v8xaK0HYjIFauxAyzGkoAHY5/mGNE74jPFW3d
Du0fXiECx6R//2/N7U7Nqr9B4fVSny3FWTPXKJHkuaket1mLrcUOcnRBxsYwerD2JqBteYtFg2Ba
WGF6M9x1gy3VieK8i4fyITAAvIgUifBRxN3WjfCGlzxyj1W744uLArEy0t+2hnbdIF4e6pyfsbHr
ZwoavjO7QS+k4Dk2IR6nnr7Hq8XNPsoc812yBpxrBmaCYRS4W3JeWX6OoDBppDOObX3tJ9Q/q0CD
45lYIW5bCAmnxUBpLLbW5W0Cw+yWDJzsE79BxJbwFfkz+t+hoexMB47fH4SQALOJg31pwvQzEIDY
NCa6mKaovtIIw9XJ5E9G3w/8Iv8idbAOnjkJgw82sNw9wouWhLkYUfBG06+tn+nFhERACxyBHs7k
tWUAU1HpYIr1vv99qR4V4CDA61siCR3BjXB0eP4GT2ZdINEgRs/XE3QYPo1hwVpFlXC/JzOsubJX
W80Gz8+THktTAcqOCuDu3IljJcku8COzqnGogUVRNt+iBmqUm5Q2u936gycsCCvrw6giCnqoBPJN
JHYec3rEf6psKtO75YuuaCFfp5UK0AHyZZiKILOo4JUdXG0SG/0OyiGMRqfR0m3on3ehXVBxe1Re
6JcMaS+kQ0wZspWPCH8ePVR437jxrEv2pbSzbjCuCZ/7zgUavTEAzl/rTvfse56M4i5riFf+MfMq
1lKTZ4i/zBcubwUfQTZz1ARLuRIKhln4T/U0z5E8KlOemmCFy2X6nd+qMqqFvmco/ahsHTr2ghQf
bIm6QS8GlyhdJ4hDhF1km3Mvv2KabnpGYw9iJlMkIc00hUEn8OrOvzfUEL4TnS+VyHQd2Uae8VFO
V/oRsKn/RcplXfhh6qtocc4g29+V+V1/JupnA9t5CLjq9Cy/nn/R6Vp9Z3RmWQaJcPy9yuHxa0Yf
qgbPeR0QWbQ9tpZA134E/QvS0Zer97qx57Nu+VpttWNKfDCxj0wvSxRI8YEBZdFvMDCRAYcz/VQu
4uFvYA83AaAT+U2aDL4fimulHKEHD3gLqaFPdL+hiE9LZ/byrPpB+G8tEUwaq59pCmUIMx8zP88V
NtBkAWr1dBVCMom/JzKUP9rCN+pYOLXC/hMofJfa5KUyHHpspQotMdIjOFoFPsococKEcaXG9LzN
1ejRxwDx2mt5r90n/zAajReX+3LE6s1V2vOpkxL2MBy+9uC6MNBpEGDvMLVh7MnV9FRTL3+36V6J
AoED2yRvznv2j6F7VrwzojBdT+zQ4dUzTeA/UgW/rEBmzbAFhQLVFBmrunpQfXNQeejs1XcSuDPD
ktXi5u0l6mO2m7SRdEJeVQkd7djqjwB7vyg4hkc3BeSR574jBaMsUfvlb/8QlE45AQ/KVBc2tuc9
/TMWtfO2JZ3iZ57FwJTevd2qoZvTCO8hn6cvi0YtEBdtrFu51YbizDHIZ5JaIBcQ5zmccXIVLCK5
VCtN1Bc57UdphiolbSEI9Hf+mGgQOM/Iafc9PXbjxIqVcudweSHB5N+O733WitcGrYkU4ZPCWcBh
719ENSp+BpACgbCXOgqOr3vK8HDrfI+4heS+oSt81cKSGpXbT3MHFQHW8IhvAZsgKFeNTDV0awM2
HSTfGvI5OzCJGmgVpEw7Bat2wT8Ltht/6V3h7KeFBDmg6dghhel7Z9LJouhb2+RQnV2NIGJNlwzK
ygOUNxuPbIEM4gu0PExwPt80O73xoiLwSM6LdQ6Qberng/hD2PMCnj/SbZt6eiHXDdkWhP2/WmmL
UrfHmkgJu3zFgj8/fBVh7ewt71oYDCd5vSc60XbqmQwea3p6+RLtfSadubhYEWwZi0o5HZnWllkw
oqVvOnxuU0VSp0h/UZg5G9P+/MalDxXXCP3TCCFJYHEVw+cDPEiBr8QKv6xnWebT1y9PneH2Ipd4
+PdejQcQl1RRxCn0ptqzkXMZR9ExyXeC9wfPwhJJJqDwWK17/FCt6RcX47grlOq7+hum/2YFb6FX
wkV+aWEek6VKPWQQ99w/jkyCN4xBFLdbsFsc6+/pOSyAAHmt89mNyqVey3x6SN7UpfpI0FgnK52k
ew9CErlJyw5E/zIr+rvgsyHpxqQaI6bUKR6/oEMIRiqQiZu4Xz01ak/k+Tr/NUzITPWHFYXLF6TF
7j4ruS6h54E3Sw9TpOva731aF4Ok4YuE9e/qPHolNLeYNGmXNXNTuR+MnVSLau9wUAsCK3B9nCWg
j+qt1rRTKNNozLf24L5SLny2mSZH5/aghKSWvRgNw2/brF6YQkldGDAjh8spDkNUoKIAra/llEGl
DPfrqc0LgvsomT+1BnYI5WK4XKRgrCmMhvC9XwFXm+6zpnfvv/menl63L7KCxiv2DW3wtJK1tp7h
NwGKM+tPJFcyNNBTHxJtTo8qfgzLzHHBK7l5hJq7ulj4m3UqRkRnDaeZqweI3yvOwQ4l4OmW3hyE
Dxi9fHfe7/IOHKBUso7c3RSaQciwaG2xoaifqZ7UTdAs/Xo7Ey7QCErg2xwBauhzAQ4LaRqBYfjC
6kqDgP0+6s2A5xGylAz55/nhfBorUb9zWEvWhn5PDU7087dWSwEZKcn4Dr7ANczm31Lb4y9rQ3iq
gg77OlwqgLr1beFUoxtqq3NpeK9x60++juONtA/yvauSRv+K9r8EEEUf7v2bkRG8KW0DO1o0pxw8
ekbTmqeTkcy4O27uUxc4IaEG5s0VK63/Or1sdGMHZODlxw3cn9Y2VcX0ZfoVMBSdlPOhe28gv57C
7WVNwupP1pICO/U9QNXM3lceA2lHWcZ6mWkCXSi1nkKOG/8vcJnA0ITNMtBAUnKlSe/uFIn9l2BK
MNaORVoqV1lv2Z+JKxSxSLkj+IpedYDYm2u23Ip+iRucayEeALTQGDZFkfBwXSIPYFfLmUUmGBox
gL1LGRLW+M6gkfNUKOtW5rFmerPzgDd+QCieWSdJucCw4DLgZ3PRoXCE0bfOfVbwx37gfCDVdngn
NlKQLkOc+bJw3LN/zU110HY5btCGLd5a4msfk9vixG0wqGdVhZwVvosb9fSXKH4s/QodMT46Zaam
fQneWVj2l6F5cI86IAEE6zG9ZtSYpQkjU1gqTxstrHBFN/7ptb5Y6UqqyEFUmEXDsoufq+XGiZwf
qQMMO2QevX69Rd6oSq9D+3wYmOguO93Qq2YNIuoQfAOGu56GqQp7ExEh7AprHgF23cbo+9nvMcTc
nknNB+3oKa4sp6/WhImvhsTj6U+HxOEWsEiIsVVaZeGKLWnZ0Jq0zCNNkM/1vAK/xr32aoImbSSM
R0KHBju92W+4CKPZUfBWcBkiCrhZ/vlKfo1M2kdB4Dv6Bgiqst6FWCX2F6kcUcxce5JeTlvoZA2j
OymEzaHm7S0xaETVFvB2pWttD6d8Z8Q2MLBMNfyNNhare7jYOwGhkqX6qWkhX2EOpHHP9/0s9Vq3
aLelR6uGgzL567rccYSF1x49DmtmL8LtjcnTt9YVLYOhm3ipMrNI6sHRqBTrPh3QSd+au67XLHOo
j35rTbWW38i4DK3nWFFqvrc3s3wSavO6cQW5N7Ppnixn3fSn0E5ZuLA+BfjhB82Ugnx0Rr7KZtOb
cKfgIjSUtm6One+ImhcigMu8M+xCkDUwbVX9zoFpTTp+tkfZhUmm4b10bnyirhaPJPQN34mI0Hx9
SXGkdonKVPc07Xx0pRfUbXRNg2W9WSm3ST2mypqFBaUwiFT/DGRukvHjaIRnt7/W4fhhHJk9Y9Ii
C2KC4UXwkzzCmG+ATYlHxUW2BmMsPAeSk3bHrMdMfQW9rY2ZwcUNqS8ViWumTG3eHUf/UbAkeCyx
3d5D9edFrIz8dKtkA4r2X74BRRfDgsjghAqLSa93gYpd+55EcSI0VqAzZRpFLJD/YG8iW/WS+h77
JzrCTySSwz7+HT5XhTsBhlA/5h+z9B67tGic/SX5fYJYJn64qz1NWjpdQ5OTj+F9OUavd6orG6Ed
gB13RN6vNC4ewxkCwPzp7ficYMqZNoB5njztnVnsHQ8cxLKKhFxZMyJzmnthr47lHD3q34VEgVzE
rH0LK7SIML2a4rV9hOP5mnbv2CUOrBqY0IKtP5ALu1wlf8Shluk3iDz06pOgoSYLBQYjGVOia3qg
qFAcrRXbMVnS3ONm3MtkZtuanWcE50FyzOYkyPcUZWwQ92tUvZuxvXs3By6zMK5XbD1J0miuCGHp
lidXeibP5Z7wL+SLL3UNR3VCAjPoS6hdmkfGhl/AZ2Khn1rNodQTNjEabJKoF6mVMCMqbY6sEbuI
VGqy2LjSaPFiqnbY1xhFar0XZsi/GxDzoVlODKcV3vPYYE3prjcSAVO+tUQbRSxINVvUMrNRxr7g
N05hG/S7UpSuiDa5+JJ4T/kNzpoeCZjR6net6LXeU4mPRK3vl4P9j9bYdVdQkhaWSrHhsIv0A5iR
eJpz8XcXuIXusQFHbuBFKs2Y3bboewLyHcMW7SzWJXPuc9yAD5Z+eVXo7lBP0TnafU9bBqCyTCbA
wSA995kuzTTda4XMj15ZRy5ng7V62ZLTiZmUgqxQwjarFDca/opPPhcdCBuNrRZtuoVw6wlVovQY
ne5RTcUaV/XvdvcV5rV0d1F3jx+GozQaeW/hx7yWrHGu8O4McRq88Ks79EmqH6vtmBzBf86mbQSh
AfoCPLTA3OjicLQgzmrY2khWtt5tWx+biL50QpBCWKAbJdb/azKe/IdqERhJh23f3fhzzQ3tPeLt
JrFDzGOzik1rDSanrJDTUPPSirP5kwSJ1ezninRK+EoQjqKAw4NCrf8eFaG1gR7/qor3ruWzTprm
YoZ7F6iBztzTqMp3eXvVRsioTROlu6GkHmzQm92YQDmFb/tZC6mC9a4vfNSDNHc2Sk8enja+mNSp
7hGayoU3MQ/bMUC+r9W+BDr4JHbGzW8kWlqMkIgdlNtWWm926IoqJkLDx5voMer6lORC5mKtTgy1
AhOdyeHrrW33PYcG/O+206r1wOWRUYMftwjCe6WNeaXECQkVsl/6qNacKyIPmK1zb9UXmh8wMuDa
VWdnLEhGMmz7U8yrfqz2V0rUU5uuIiBrkoFptTtONS1rMRrz+UoSbamc2edsTVmCvmf2O9ZBpzYR
qqaFuyA4mdBrUZufqFeY7Zk3jLL5dBfu+xk9HlIgGE3x/Cd5MqXdcpAUdN80pVjb+3Glem3iIc1a
c/uO84u5YxrDj6GLjrLI5AVBwibr2g5umnd+ZO0UORESF04rRooYeIgKa33ftRFtljedsd1jnvs6
ZTmF4CV9Y2QBqii/smYwFeQEAoytinPptqrmHnrkPrITkknHMNPwdXyRGjLp3ZihfbrucBu7Zi2K
F9IGOwhgA4ZT2rLww5Js7qyL5CmEQSh9LK7ZLYqnPlA4/iwrDha+fPmvCWEBSzPG6Zf5SFfWVNOx
iNaZrHOIHFrcdy9KQSObXOzpH9PR69qAqNTkrxYQRCAPJCWPg1CmzJgOS/IrWPMThgYwvsaxMS/j
jFv8CANDXmWzJreNjMKd15xbqZLGYLsNYCSmDiHCo062zthx0d4zuwzs/EEiTh4xuEokzeEQErs5
xFmCamKdR0XIxWFtL9bjyc0gA24FhB/CDrtl2LdjM+IynvLM1B12n5whJKgEjAQvRcIztaSBA0BW
K0htkpmO/xklEDv+vA4OYTlLTWaaNN5+LE4QTfHGWSPDVqKZbSSSKfffrZy1uGzMLAKYU4CciSUX
zfdlQ392+L55nH6AQKVBdvGAs9WXdc+BYyGAW7Rv1MpCunKANg/Lg8MffCqtLJy6y0PIi+xWNaY2
CNIMOkv42ojuF6eOY276brGC2AXoj9O4gzmfkowbj/An54UbB3ULpQNWl1GsPTdlSRvd6VbaQdJM
MA/WOMmZe+HVp5sCi6Qs6N6qGzb5x8N/J+rbr/45RlIJi321SuGSxzXDJkqsKy2kLl6CI6BhTVFC
yTjtN3KYNLi64VmJMhz6KJjXko1VBMYAZCLh6xaSCu9f8fcMQ7UX7sZHoKWHgYgQy1qBbqwRBs2w
MNuTHw8HmRISw2QAjPuzP914wSdEcLlPF8uTCLt5O0It7tbmj75GiB8shaTtaN1gUZ167REaL1BP
17nJh6XVVfgm/PQypQzvmJqpCLON/y+LCZbLYdrGIh1NCW6M69OsKOqdbjSG4kcBdRy75YF/+VZf
lVYzNhT8GESW/FKExQi/8hLHwSrtCPKVE7OkZ5Js2IhHCHNCtRgjBK3bFmKyJJIhSVQ/aiWdHsrT
3RfjKSrN3lOD7UwMCoKiQmMu7lyKh5EZLuC0KozfVu96TE9rbk2Naj0fXtPPdie6rMvckgaG/Jaf
L3JRvnwEF9C2/D9nHfyqFz6OpfqSMdgxqjdoQNYYdSO8fqfm5io30XRB5gwdmbHLmBaDzUfIahf3
hu57SmF08Ywb+AwVwe4SpIuyDC14hIpSffRjw3xjWWwWuTxoM95MX0bpW3dA4cLw6e6nT3O/kCR2
pNKGfkLp/lNXQiXEgvdl1Qlth43wqQJ9m0Bvyl/ZBABQ997dN7j5C6af9M1DFK82Y8WFEmA2K4WZ
5kZuvzGMMInNPIG0IWxgMXBl9qLpYs8Id4WQOLTH6OlocOma6BNr4etHoeqFymX75yv9fQBxk2mA
75VpKA0J50YF9Qq2ZJGaoxZ2rmaXpMut/w8txZ029vZDQU3Nk1w7R4wwwaQ+t7ryXk/avXhjUoS1
xx3Z4xbr/XLSVqCbzWpDKV2NWB/xKMuXO8lbq3RsThsQWtEfz4meyw6aH8ChpXBEBr2QFto3pjVz
RNUBIIQrX94CnA/xqtC5updk8nHX5Wxs6YsknvDsaQDboWpGEjgDPtQ2bgIVdnn0yI/z+Ao0FgjX
49np7PAY4WQ1lsb2ML9UP32QULS/eOxTBJ702Dxambr17M27OeUtLfBsIQ+wH7EZDX7o57b8PR/6
oMY+m1mV0Py5F/c1PlKWxXWI2jDC+jERw4pV6Aknkx39q25db0h5bAIimxnkUtlM06ZJ6vexpGoL
2FnzRXovLZdd2e7J95tCCW7RQQPXmtMOqdesSQTzE2BOZbmsHYdO0yO5lrmKleNNKO4xRjsYq2GK
D78814DEZPmOpfd7e+hvvBsMXlVZ+LT6m5HX1j+fIovWX0dS2/t8geJuJWmNNJ5G5uWhe8MjKyu7
hLQRngOcQkSJdesc84pzk1B4rcw5peBrmM9P/sU81OeNxaEm7BWQ5/pSZzSkeytd7Sl8eByDE3mc
HQEyiB1tzgcYadv/5ohVeQIwXCWmwR/YFmB5TpbGUW1rrIu+HQ/VoHHbYJx15q9SkIP1OaRP5S8G
WU1pmkwy7LSAJS9pz/DOlD9CpvYheKlwoFEjjiO/GJAfPOqz/OEvsFyjm/xF8v+i2tdiOhzrLOdD
Xqey2Vg5TTmOaa0u/Li5NFwxbiQzjjQbcY361DkQaWUBIAMSijPLC0rtG0VIiA43KPQriAJuKcNt
twm2ok+UNYKGpvKZ7qaAs7cEqY4UWGlFpz+KT5d6L56hLoDcz1OF3llHRHaQ9d3beqohA7Tw7yUS
VNp045cq/XIRpoz/CLV3ECs6IXW0GB9nAigxnnl/t2HgLzNYHRZhg2OnRgUIfIcGj1nn12yCyDd7
muWyP2rMMWJKMz6s7TaAb9nQEpSBkFUf2gVEmxzgCqSt2E7Y75vhBXgD6T5NjSYAOPPdopqIqHQl
AliS4P60I0lQu81/wnCSc16oPsAaAReXRrnmucuRhtTZ1+TyBUnSIZrhYfb52ScsDoEw2/3GveTo
EIx6MAi6LJHTUEnop2BqeHBrHXins8Yf+zL3Q0umPJlxeNKTb3ooEbVZ/cb1gujK6lYTBEu6IiAE
B97Ng/XqRhUYRbsE8HT7qCCICHnUSgbHzAwWoLXyWPeLY/xJhK/HSkdiqhh3d5K54FFcUsDA/0kG
YtlLPPT8atmRR/clD9hKdqaKj4H1GDJ7iJRU9Cs2vpwszdb+TgYE/F7O3/mg+gh1vmJO2wIf6zIy
QptANUIO9ZO/7jAalAyEu2ER7YZ9ipVO2f2zYBLKg+HHOEbxRW/xp7rs1AWaEueG0QkC7QCjdJed
YFE24Nte/U/06vGaECyAskk3sj4z7olxwrkdxRUy917XSpXvU8fruzl64s/EHgYt2i/Dg9k0hilD
0WNE3P6Nx9sqtnaq0A/mmps+Ji15aRAASfgT0abbz3JMn3r+27svzkj5nFf7lXjatox+9cf5s/1x
pSidMAyzaCQRkfI4mL8o5sLJhDDe0tr6fc8xqdtlvyKXCh0OfFbFXHtuk4TjNKqmyudtf3KlK1ZM
1RFU4Ul2PlNk1DnWwGJS/AXNYq9OzY/mfevrJdtrXTEYA4K/8pFleoV0LDSCvy6FurlFM3Kh4CTJ
9iLv1VclbowPHlkcMNQWg6Nfd1yYHgKtdXSZDOuw67MpDF4vwwBdwGAG46xmhUpTBWi4XALdkc4l
M2WW3C+MTtd64CYqLJxPAFf38psC48U90dr+WM55aJy4jXwCiLs/QMcu/N41/SdqLvAyDLKXpQOm
IN6ilC0zP8a1YTJ5J/h+IxFE5MWCUBF+u2d6PeMCvg5vvoyVOyJHTT5YdsWwXHJlIkCNxDyZBvs8
tEmmHYLPHIYWgVLPcXD+lp1a9H0FBY0EnJnaMwOQgD1m8220cQEH6SgkScxhmXmYoXuWnumVfLkm
L9eH7ww6wqpXK9MK9N3fylSLXGYdVQLKy2Ge1m9XNpQ1nEU/gEGtubBwr+NCaTQ4ga3jGpaSHM2O
U+4+5Ch+7FMavsQYVGNPDMq033NA+pICJ/QodH8Dh5s9EDMY5IlSCyyVFsxPnuARmOQ6W2sP6CXe
5n3+r4ymfE+tSlHJG9MouFxXicCfCCIPvC4NIz9VW63Z5p8923qICE+oRcuYB+/oOWz/6xZFVtMd
CtiTPGN15A9XupLGrVGonlzfq44shz5hDo9eBO6zQWk+4zu0R9H6TOHYxNsYIiFbO4tqRiL2lvs0
U29rUrv8W3XwfB8my2M87KhjcXgy5JOWGUhf4/E+2AYY2+1+2hc9+vorWaTKq/zmJoJ4kss68q5J
JMl0FWMXEubTihJDfNqqkwVgnH6ghnMWlZhN3Z7B+QbXXkZ6IXmvfjzt2vYYIgOqgvcmx7TKtAxq
hh5V96zVy1J50S8wy8DKf7dpBWxjJ6MCW3DSdTHjcz2YaZ7PHpUUdF96J/WMn+aEODQxVwuzRyPK
eyFZXeC2EqgSpW6hGXfrAEgyB7NXayv2dnF1KiwxLl5tesEVPa8nGFWraLgiwqwjPmdtoGcerPkq
X2dIfCGNO86i8+SN+gK7LrRnR4QV3Y6nidEHRR4kI0LdtqWjh/nSxuUGWkjbtemKt1AvDskcFj21
kaNAAFtUdxE9YkNg4huV5juvz6zNPpqV1I11fCBDH0ChY3hiIdnifZX3sF47zla5BbtTAokxhy2F
W73UFNFE2Gl33i4vGWxEErOxujHY8yM9EeNqL64zBUSO3ORdNBmA0IKPVx8HOdBKyp+b/Mq9fUpF
AI6F6JK1d962ymri9PuxmAdxWPgYu+/7PmGIQrf5b/D238z9tjOkNfAqYuVbrmuBJfEu9Q/L4suP
AaYHA6Lebfvx19+S9eEJa76zQG5xhfr9vEEh9xBS1BQg2mibMeIlfnPD/zUyX4kmc6C/5cEuQ+nL
dIpqmY/BlqvEqEe5Yy6CgGl5fAEksWB+5LOOuMCC6CWmH7yllTroaUyNqv3r5U+VCrH5Pu6oY4MQ
tG5JicGn1TCJKa+M0MCH/4AuQIxfGwFIyQnC53E3gKROyxE2DjyxVxps0L+7Mhe0XBJPhVEp2jzN
dmE3Shhp1SUz2mb7e6fu5Y7kLZmHmhBhMZgZ0XI3S2aBahMO+xo9dUPUH3u4sKDZKA/ea0JSgbGj
aU08ZkTyFkHvycgrkl1Jl5BsUlbjtqf1UuYGXs73BN+3wwHoVs9j3CUdQlH0NAY06lo/nTlbBc4G
EQzJeJxxcgQMvF7v4MaD7fbf0KhUQUFOQ7/JsguQy9qhSKlj4rd5AjL2+r/qQWclHqcXoHsMOuhz
PaEjWMIDcxFv/3DSfEk5DXjlGBLgUj4qYKrL33q2Bx2ASPN63h3EnIJjsLVT9Geua1j69DYmdnmU
CS9W+sYM4UCO0iAHuPFNs+AjhyDF3JRIe8KcUKFQws9NrcY9gZcXAGtQnkCtoESyEwQSY5lg3tZh
wZNxE1wPHKpdUq3uAz1CEfuzIhEK1sFUSwNNckC4YHfSSKk+qq399TDfLS8lrj2i4/JImJctQ2Gp
5AhHQx5thBDrWIdCC3anXaJxssSdLJ7AnejOjDHwdM/biMET2asZ9i51mNnqegb0goksV9r+Ktf6
Ulnd1EoEt8pr3nzx84H+98+u72jWm2Ye2NGtkqORxNdLiRWm0YqphPuErp0APLtvaXQ/wSQsykAi
LCjqH2MQyOIkcdPCPYKUWsGXMEBQFypLmQHzfXync4V/QiJs00biBm1Rts6YvCpMtXvGZmRWBpsZ
rOZvaH2+f6+331+b0WimSBBoM29ZmWQXn+5le87pFeuHxNUn01h7+UfrIWEJ/ldUgW4ofC9FxODh
Plh00ove7D//hMwX+O1awzSIgDkEQ3gAUGCJ2GHgDJQdeD3HG6n5yx8u+cehaLNs04lZAyZCDgT3
RvSI3BuKVx+252tMbWvVhluTsOd/3fEeAFE/SkmlLBY80ezi2lz8ctw1fgkudK7jSaP5pLuJyQon
BZvv93hi2CPlnbscLZkY84NqGhU59LLZsNNJruNi0nGs+hl5/kZbdX2bi1TUvcm7KvBndYOrhFPd
aveGLIUwXILWkyiC2Hwwp12AZ0a7AwhERlorEr8ag3BpehgZ/xEDz5AEaLTMDdMNVjS4p4Nyvdjz
+9sy6j3uL5C/KrcaGI2FK9EUsy8fMbu8cXzIZLjCeye+oScdF4EzUWV3SXousnjRQNWvWdWUVOmf
nRNpTRejwAK3CL5UXbi7dJU2hiuYkToW5aupnwQxdnSag/sXrgdg6VOIJ7bQ73wMj5llDrVZT4PX
AO8qyG/5Ujz2MnjoPx1ZdBdJCQ4LKN15Vam+O2KUQmA7FBPWC6DI93nvbTqPwyZpkVvfYL1GlZQE
C9GotOSTtbxyn9ZtkcEwwi8TtLtlAWwvlpEm1KuDBT+nfmsp2mwmPPHpUyLijphXN2I1LCg1I8cz
msyNU1I1hEGFhfDVJAuUMi1vXYg6i29pJR/GI1lxaaAt4vEvQdwlsnljr1267sMSFvbdWm46qotR
nC1I18hV6Co49mjqokaLWdlChpO7c0PQcYse4XaMXst7nhrrFMXec64vNnyw2std75QAp9igiGbD
+KQiXELuw4DL99wIO59VGNCC7qLjStXccV//HR2Wc2TywvgF93C3vyVbt6fedZLzPKBN0ndas5Mt
BTk/H0gDQ6eGqw+cLZVCp2r8hSp4S4I4QFaCEMsfXjE9jWfhOczUC2M5r9c4XEdkd+vTgxamiQ4X
GFgGLezSEOmHTd5oa9YCsOZ0DgY8zftg9GgqV/Ue9+7AGHYBxt7ysjgJAagh/kxDG0HyPRvARiZ1
F2S6oAQAwHJjC2qI8/i9T3shwEQplFcKFoqNO9dSI+Ykwi1QhnF0ybXiPM9rv6xaMY1lpPkRt/3z
1nyWzFE9T3K7BWwnpujHrqqk53Cj/GMj69W3uYbXrS5sPvKncp5jKHjsP2iIzcBJcbcDgGQeVQxm
/voxGA1pNH4qODqpnP0GyLe9VEPvaSD7yp20HHhHaH2BBk1Sya6j1j6qPkOKJ2CZo2AK5cYBNODD
5R2MjLU7uBeIUfi/Zl13Oq1Zyso7YhiH0SFB0fGllct9rKkVAkhlCaPnFdJIKr6FV2R0756wCQHj
QSLicoCwdQpUHkvxWMVImvIVDoM5hS6VBE7U0Ji06VUSOSusCX0stcifMsIvcrYXihCFzFMJAjYl
FssX/cYLZegYklMEnQ+Eec8OshNqexgbb5QN5+AhTcMcWfwYCe6Li6VIEkRpvYxF8zUhMx7i/CJ+
n/X3ggdEsrBHwzl9T6EFs2bUDuwv/lRDXEZt4afLw+BDxx1OAs1ZSDnlsenC50Lq/e7aR0bB2HBG
7p9wPk6N77/LR6ekESV6vAGFD92AKCHcQcQ02pB1mhgNFXMuf7FC9E1NgZWwedW2WwOjqKO+EtJt
+94DhacRSJOwY7MVPfIf9cGiiD567CcYHZejTwc37/YlerXNIAlhJTQtMwnmdoz7xLPuJbFm3tOP
wXbNDSrniPNswGpuvNy/xp5YTawr4taB21pfrGaiRGRmREyFYtkSYPgVAmUCHYo/RHbUBt7mXiGP
91w3Hq/2YSEv5hy+J2vqeWYK8o9gYzkSVw5uSlnmH6fpTkHO7n7RowlcU+UOtCPgVedRJ7fq1m9+
0V/83YAOXmyWo2t4leABQJiuJXh28+SKLPt1v7h+gHB/Ru8+yg2Y5YRVm+r93DyhdkXFu9KHT8Ih
01h8r0KCGcpkYWFaf/nYI1A2qR0jACchWYVo+dDUGjbZ6jS1iqtuctr0rVBwsVsBMp9TIlu6iScC
RgQvfaqxBI8RjGrnw6v4wywFbnCXh5cAPwS0nee7S9/GLqfReIPrtOj9iDvsLreRD5gdeuCBBHmr
6exyeuqnd6xApilC+xdPgBLR84aY8b/okX7GSWmnbsxqpA0ZQBPdawTTDEDVO716hhdgAaOTtrbq
3+j/wBueq+g/aDlRR94HCBkSIdk+TEWmAoaAR/LRxGot2EsoOyLggNY5G8coSTFiI7jAegKADzSh
P+pd5I0nLJyGLdtgCVRkWRSSJf0AqV1JFpJsOWKXotFND3xfCOvpn/xBVvOUzS+VElqwElynwMGT
4yj+ZD820d05rt8Tec2vFD6/BQQL4GRum6OuSZoupTTdFALbOS1ATX1Ip9w/V5yqqu3u6TNqBFST
2cwgpkteQP9WnbwBrxrRNKs+bWEI7csJvjoj3KSpMyFuKOgfrTMa2EM/KxcMyS9B+myvboX1xocY
CLFiBf1Kjp/UmN3pTpijvIqvCv5mZbsvM+7ruNIYTJ4EAZzGzyHCpSIsVSGknp536u7+rG4U1mNZ
hoVlVRUdfKjsvQEZik+e5yqmUQ7vyiU3GXzKkHIOVRsQEkxiRbCgwbQwLW21N2FZlYo1HzBWlYy1
cim57Y1CF1v6fhb5y2p1mcd+np3rI2bgrUOuXN+rMPmapXli5pExAKZ3dYUj5FziiJBi3yzJhm+J
EOwMJ2wsqV6ihuX49N1NT1lbvp+CluZvhzDu9ELcCVdd7hwGMm3THRU07IZ1ME1Qsg7qiwq7Jql5
2yOC1SQ0cBS1oZUbyO0kxclrD/vF9bOik9ZakSL+q82X6q9+Z9EYRXvs6RUohmwA8Dyo5RqH0Uns
joU5jmqQmu1Pc1v5yyZ8JxyiW/JHYBBtI2fZP9wxRjn5IFvj7OgdTRZuUJj0+ABn6KyXpQlP9Z7Y
1RY+M7C7S0NBCjwht7klgYuuYApeoeR6bizefAdlDf/m0oLVUgrH5ueMBsO7cTrhJ0/JEXOxJJUu
fd5MY077Je00XFl2TKscd88EejoWVRktiDFxTcOAilTGcpQKFW4myg90IYo+U4StqSsyCb/1LnHN
agof1zx8qYzY747/CUO3wRbS0cYw0MucU8J5S4DLT/7PrY1byqz9sMoL3qu8fYjAYN1ds0S7hgid
7qGIGPhI+Eg9U6WVUJo6PujxbI1pMcfmnCVI9pMXC5dz9BCqwWcXSZ/E3kuDHEOhGrFfbOgwlkfM
/nWD68jRDUz0v5Hhi7OI6OmpXs8jL211pVrwiEf4Nd4O2d30E2WcyAoBABJlW0IvHhKwHTCpHiLn
u4RkdoySrLa50FOak4AHC4CH30uPTbRS0pdAIRhI6qdxDQAhhl97ZhUF/EsbYtvrWpPnm4LFinlf
1R+jxM+3WF8dwHXJG3mX6W/FLKrZOltc+bqdIRlpNbmWqcmF2JGgRPxK5jiza4djahoNh6gatKKq
S94Ru2atMkTjjyiO+i9804BKhhV+BdFVAJcnGkPNy3gXnxY9ftx8OexBKmgGMitP9zDQMbhfQNuW
WmJd8XfIp8xIcxg9McBIrLXfTOOwy7aFTnG2Y1X+/Vbff6GVYJOLc2fN8Jww0z/r9Im+Uye2HzQs
PpuNFCMTU42rmt7tCs+FiypXII/El0Jr5mKolXFCJU4P9IgYJVLR76pgvnD+XVncu5JlO295ePe6
zpmsh/xEJKArU3HfOVwozfW3A/XbMTIQw7tSCv6mFoOJ4mLWeaKqqtoKw7Iy9XTUpokho/RJRXuA
zyuQuNUM9O4OD9670z/83HF52dJkElAeHzucJGa7Vdic62cWTn2lq144/sdjHU2NGPMFhS3YyJRn
SXjyHif8C4iF0PzrbpzZUsqqZjMSvBmfUyzzlrKXdckEywXe2VCeH2zceKNUy+uA/RFlYK21N3FX
u0Qd2Ux52I+juCBDuHQBkiQeaDxEIxMxvzq3247nv1P1aY6KNam5INiLjIBDRdKzdYtVvKNMJou7
fj8hCN5c8CeFVpXAIQi8JvtrEC9XN72wrdOoNiR9Tk+ppqDK0W/FqF9FBVfQIDs1rdXPxU0uj+DV
pIh+av0olSUVTnzKpu26P+mjfEABG3+N3f/Lf6i2DOGfBowEAIzDlB5luNCjQ7oECVqsEQUQzV2+
yokT78OPJ0Gpo7Q5TpueQ9gZ+Io3NI14aMn+Yu6O06DGMeLkujBFtWtQ/z5+Kx1ojs0T/OiNhmHN
/yT8485n9poSQFJOSy9c8TEbawvoxvaZfxqhErZL+rzE5GATCvojFtABtgUJiYiob7aSmVwvuqIb
Ipd8MjIaKvbBk7fCiuEehLpIMR/O1nDZbQ/01RZF9TCAltBNmaYmFQJzlmbSfEranfZs2I8ztYcJ
9t+fuXhzjL231nkZ5Mxtphy8sRfCAfTqQr4znEZfJ3JSMs1K0FyX9RDFHEIwnAjrupPu3tOwDu+Z
SEuVnzMsu48UzRik2jAd1OP36gRSskl7GvvrLsM0rAVYqudocEON/o7ifOs0ijkU/veyOwtyG1Vh
3Rs+QpoaJ6hWre9tyjc9uZEI7AskMuAS0fw5lyAMUKWNrqJb4PponiMLH+JrDheCz5qVxpjna8or
xsCNMOGhKFZvEnNfa2WGw+5old7C75Hzz2BbfJo4vCE9CurCG6mKEMOjz3lGovaHiUl6JqhodxKV
/8qQrw3n2P1qFCXYjVt4pU/AXYwGPakFLG/E45B9lTWTMJQ4k/hAi/P4OQvwlD0H618NoEh8r8ul
+pCI6noLNv/2B92+qF/PL4w+VlfrkX8akmsUKPpxS7vkq9xiA4kiHJ7Tyvsw1ulIE7WwGxoL6oaX
F5m6i+98sYayxpbMZWdvdS/CXSo8mG4s8tTW1BGMozxW4yiL7hhBWegLCRB9/n5ev66FrFy3jeM+
q11d1AuFXaqX4KsRCR8h6AsElGj/1MSaIepUX3xCNmK1h4Mhd44uFIWNIrvwgLU0euLf49mWkjTo
00TZnpsdetsj/H+7FhdTmShRU0bd8Ir3HC5A538MxD5x+T+ciwFwfl13+NAcRQa5Tlsdixh+OShN
KmZH2QHUMgKn+oirSfiYQfgbo9vJCBgQe2f1pFV+q+y7b7FPDHcI263LTuvEMuyZ/xGK2X47dtLY
tc9Hg+/wjaYutqu64p1/PVn4BU/bhxxTd0SGyxQJ54dmr1NYQyT6L+Yz6rwGbV+0a2CrDu4Fmfri
RoxNRoJ83tm3ozs6gZ2Em4rdbSM10a3A9OhXsryQSOeNY/DkyxTG8lfzjmuLoNyOyt3gs25p2NiG
ffAyPGebEb3ngSpfHL6HXXVvsvRhjBhDDYATQW1mAXHQvvHMMV0zMnfgIJqdsDPKRpENWP0pgsos
IhLql/AFu1Un7bFAnm8q53KbOBLhOP1wfDEXbPpqSAZGliSMLKzySRN4CONO7kPoykCrzbkxgJA8
lxGa826tCIHI3dEcvOXN1Tc+SVhpDhJV0FBs6ndx9NIBWKumjV/h54WEinP/8OlKPqvMENeZhtXk
OODXVDNht3dC0YLCvDR3T4TVCW3+nVu0DhdNynIatzSlt7rYtka4syVqh8Uce2nh1cbSWyuwFsip
w0gLx4qIHfDCQbX3PQ88HWx8uV6STJU6mtSjNup0HxYU7WKlE/2lDf2iigZGES7n0+fDYhKDRU9r
zrbKoX0EMAJFqbjagRebqHWd9f3aFVnIDr50kEMQ0W0uGDExfYOFz+H7EVqdpEi45iWWz1rUxvo0
tRLRklQSY7DFm4jX8P49t8QbbqYpUjA/nlLcQ7dkUrXQp+4eRG62HDJ85ZD8K1Tp25e2VRrJ8qfC
dDl37RV6eFkd5uxZu0Sm3SG1xbaNOMydHlCdLUsRNiAtQCzpzf8CVFyRVv/j2B3P7fSHW88mVZuo
5CMQ2fmo9HhQgxfp224dREDDmtKhE+lAR+wDGwl0KJ7cJHCpUuzf+rlosTrMuRY7MbLDGPD485/z
REGlc01tsh1zWn/EP0iFxwZv/zFGoZsTMy4NBUj5lhmKYeiKwHxL4wLb2qSvrvPjJ928hvU7xIpD
zWFpNq6r9sFRTOOvPusXBb658e979r+G6D3RW/Mvsz5fYLodD3D+mEb1aNYCYJm906sJiMtJKT5P
gneVZvxo5Uyhk9yxU6wq9uxQohOd3QTpm8QcHHx6wotStFrTpoKS9nzSOIeYjYirkIlfS8TldYOD
W630IwkaNQTrqnlOZiReT8g23eW4GeQQzLOJflisOrVEMzpHJd2N7+oVV1Hddoqm8D4gSp3t9iyt
O9toMg3X48J8W5hgQ2tTk6FMPTM+wzXDBntnh2SClEv79xwvP8oA493AqbvJh6vQa2SWOTIkkgTA
CHmLt/QTg6EHaeEYO5o3PzBKpTFxx277w2TQqeeJOFl2XLPTwDLQARXUXuhbYhb4Ycx/mEPsU/HI
vNtn1olyMhD4utSpJ4OOllLh3fRGuc1acI6zBWSK1c38mXV0y/KP1zYsZ7cwomPa2qKi0saEqSJG
C5f+6ePmtTwy2f+Mb8NL3yF9gcEGS0B+Uz6nZKrBugwMNM2Meu9W1Q3Qp/ilozFkHzTHVW09LyXd
OysNvGJ9cldSx8GqfdShdSAiGUOScfn7j8Z+L/AKFuTTeIrM0enXLGler0kmpRbIJL3pNXDVvE+c
P841WYN9REGVekC5EKLEpVYe5hwIpVwJFooWMUKCVXfvJMjn+aXo7uY6uBxvaitHGnuyAdge/F2s
wUXKRdbe97g4OQhJ9Jy/ORzOiT9jIQcoD+OHvz9dYVIwI58dxJh4DmMp8AbIiNmSQbnu0VqaHb/D
cQDPVe54hL8YCX/l0rmoTu8NRLp/EG7SGnlAKiM6czXJILY/f2+i0egtj1uTjmdjtxo6klmtXCMZ
GiTvRd7rOKfMX0CABaHTmHzCqUqZCfbMWK6nPTf/9aRjGu0R8kdCOWVqs/r2UmHNuOzsNS3P4917
7SGo0ukRidcuj6D1CTP0OIsoePCRiA3tBZ2ywjcBH5yr6IFl4obf+sTA8Y04Q8OQtCW0oYv2oQpI
pRFShKT1VXVqua8yRqgBGoy8BTBfRwqE7XbhwjWEhJTkqnxBe5QPAvPK2tt8Gnc+EjTHUsjgqmkZ
2Y/Zq6I9YqxjjPiPRZeePYQuBvLZqjaTKd42yelYcljwU3CNCNqQw+QvKkGc6JJMBPgR6pQvWjTe
P5mLsPXd0jS+5SiWwKpCCXjp25aAuA6GscknZCk/2ZGbbxkV0MTjE5w7hXNjOIDFwJd5OVcfafvm
XrjoJvoGRgQUKhTTder1UamilnAahzeEFOCV7dRrnf+0uVDitdoVuvrm4NZO8Ah6yl6y3+zlxYxp
+q1zIj4sVtoyUfK8ygXHheCDsEuKKKphS91B6HMFMt90CaQM1xKzEa6CY0NT9c3c4glvNSMGpYT6
RiRDER2iudguZvbG2IgXVJN06Mkn6XCX7yus/oNzvhXIAF8fpEWv8HU6Fea1GsvtULFhgiutLs9H
UiGGxIl4+0xwP8V0M9k6u3CI4N64Zzi9kPs6TXR5I0So/mRdnDD4CxcgIkAv98w3s9Lfu3c2szGh
mFzdDyDcwrc/nmz4XoVf+aoJ9nJ8+FlJTmI2qWQt7Yiw3l0Ro6OCAoI7Hx9OH7ImfN8zqQdinpPi
aDRhngqcgIY2zwQloeH9bqg0wlp/EOq2Z/LMLvS5FuOSV4YvgC8PDeSZZBx7rBVRfC5CEyZf8wQk
aWdbaUP3jYdbnkp1OwgDlT13tg2En8VKxo1jo85r+GMHdLqxW0KoQgcV+uEibrcfIb16FRBeMdS6
44BcxYX9ywxdIbGISZxJkO4FchhjRMQLCV6xIOZ4xV/8y2Rk1bWPCl5UjVaK2GETyP7euNd0eXWi
xt+tTegNyGrup781eL3WQDu+Pyy+QtsVIFer848alQEoIcuIZEk8chdvBONchP7+ALSfAqDgVLm6
EcPtdZ5H6tIRmn9ia2jiP5WbRrr1nOqxCaTSI6i8O7PBpgmfGuHAmfDRT5oIJp7T7C0w71n4SYZx
QwrQIh6s5TN7HtPbuZv4Qi629lllURyotT6FirwRg31+OPylZYE1i04glxjoH9b1ntZwcy72Tds5
mkWOWBsWsMBEXegzbOyDE3ZQjdorJ6IGcd8wo+Av5lodWQlim800KlbFguz2shCuoor2aSE8LKeU
mIZ3HMa9pls3aE7QH2V0fGtpNxsMeRHGb55LtpLTcaRdlt2ZCjvvHJ6JQHVZ5sffvnCsnb7yahvF
AKnUep9Ff00makljpk8TVamrn70+0GNxWNx04NYCxrO2lIWHXQZa/GAwcXABg83/wNSqVALPxpQa
Q8m+XTGrq8v6fDmm4afQQ+TtwkEtaM++cI3KSQur5w2sZ3V04jjYG03vTh5n0+qRt8kdA8bCWBHR
WKQfrqNw18TBSeEGYMBi6ff24Je/ddbI8yyFD1MOs9OytdyIveXMcjyw1tbbmSbweRm1dmywdyNt
FCXVtkZnL1DIMclOvxmqV9BltEe060mYxLd69jAdv/eRkjOfR7ZvRpheCfRRrCY1Gb1XEqPXrMkt
Wl896I6f7iTJF0hxoS1Z80uwG0FDqYiXn8nklwKqjulfekUXHT94h1VHWcRUQSAly2flOIcmuSPF
irbdxeyrOp+JH/8bNvooclFaeG4QEZ56rIStqCao2pnsDoHqWWHx4JZvya40A12CVakMXEdWv5Gh
b42dhykrV9jIemxxfkqEtDekw92xMo2qsnrgnYu6ilajup4PJeENaYP12UV0/FdGhagvNiYOp32K
u6CTsU78UX0RzPvQFxD0GFllMDnu2xw5nEhFaEDy+a/ZErfELZK0qMO/2QeptfFTNheBT5Tl7wcD
BRK3QTVt9MsvRyIsIAYvxS+ZB2CN62uqiRp/oua3ThjWCKA3s3iV4BgJwxSKJ1JbBU3qb+2L/VgT
f3A53RPRVBRB7wpfRl9PHMT/vN21DO4VHilqrDWjfVc8BnSf55uj2of3pnNUblzo1burQaaYMHgm
RekJXKnHUB1P8/HGJH4zt35bVOYnCGZucPI3VWJbXi8HmfskpJFinRcM29Lyo3wqmrLqolzkI+VO
fc0tWzmOiRAb/LAAqOpa49eH6V3ip1NGDyniHRyZxvnaFvPBw7of0b4HDX2ySl1XY2uY1+I07uPc
YNvq+rqrcJpUh4P961YzzJyzXRT42uuD0g16Wf7V3EN307TMCg/TxUb7/htn0whXA/V4WcX1IPjr
+eyGKTWP5Aj7JUBOzU2lyVDEc8XUvBcHDi0pAkR3U0dvpnn2w6Tnk+wHP8R1h3ZyyJnr57te7BgY
XkCkmOlmsePrrz0talh2Nk/ytrvIl45CeA1gRspcwzB4q23KQR9ldYX9g+FEhfgiw+WVTR3sD87/
TRk82Nm4rr0jh6mZMaZC54U+BawOhsgEev2z4lxXJRIeiNtDf0nghnqcJ8bmb7ZqoIRVWBbuUe/K
xua+w2tkRujp0/0lE0kocHTayZr7VI5xLSssz+4yHpF1IWKYbES1YbdLgJEd6Yla31KiER/hFA9I
5iY6wUkfh2qdTxhOU0txPZmpjzuYxsSLj4ha03k99/9GeZ5Yl5zIxP+VW5Xa9aW9tq2Th5ZEXQnm
gZ8lpsOpRXu6C7aoDkdk7ke0ffxyPNkO7sXyGOw3OECh3aWu4hD2tFu1BWfbNvKaSannC7DPBykD
394kX7QGoAB0+wjXEOE9lN6Ai0kg7SS7Hi56RmID/8hzSbUYs57k2EPAjHpBWuQK/f0ILGMVI0SS
Y0yeQUg3aQbPk5sj6+VR7VwpB1WH5A7Gyl/ve9uPJMVEtgR87s6sEe+r0NltGSo7M/1hakegZMT/
pE+5MhIHr9Vpn0sLujmyxK/7tsd/cQngSY7umaGfbJjVbGxSERWe63mN4I1ZGWAY4SU2Dg/GaSK8
4XZ7o+oIZMgGK7WknZy0GYYimGLrCQgsttkK0LscwszieY4D244H36ZEbH+xlpZE+Voh21sMfKIj
X9kXL1WN9i6/QR/IYJ1VlQsoO49Xb8rZiGQu1Z1Rj8ydPLiP6KDdaVDQjUSZAz0X0IOUz7yzRJdG
XmkMttb4HPUG+Kcm8PbfDI76gvFFuMWTClE0NSCgOmv30b1bZlha8cfb/ohxXal62fBhbXsDB8GX
OO95IeF66M5XPmyG3D57asLv72CQ6zfXwIPhTBDMRY7mByd0fCux1c1lqpdZlyBkeo+Pr4GVLxos
oxMP9SnT2hYp9qrkwAOuKPrTV7BXEh0jB7ujGHJWOTpDlFR2uUAf1mVLNVS3ZkoNxXI5ZCazb8pz
ecB7gACny4e/AyY+vVSyzDU/bXCao0cM1+dqY1sA1iV7jAeNkSCDViWYDy8aFNv+q514pKmDwFUU
05fubWdT88n3IO2KT7TJQN1vJZD2HTPhyFRuqecAGDwxwyds5jhx52yxg9cmy+/KB58v+gXLZaff
FA/chdv+gitouOJkmqI4x43gHjGmJsRpWL9c/tBQ7mV2ROUhynBF9bNuOh+98gn/34P6PivWrFRF
P94zkU8Nk4pZFR5K98gVP1OvvYKpCwjBbuzVSLvbOQfN+OQRjNInR7UwzKUgqDRlMtNN9SbptXlq
1C9qE+91u4abjKQ3xCJfI31k9PUzzO5diFgqSHSvDGUqClN1p0BuZvvhqN8rdcQ1wPZEBQ1DqbvR
2mG9GfBplrppW8PE8WQG2NX0221I9t5e24W2oG4xFT/Th/Oba8RVL+5h5w5g37GZdMFclCZMW8wf
9KDISzgQYQk3g5bfETNfJgPdMuJGHIRSkdrF0XU8SZ2R03ijaw2XVo62sNM3tVnDZtpfh1OL9dkW
SNF5wpIkkkwixSJCL7ygGfIFtQGsSmKU73JwJEKzgcSg4gIZDnJaW18yoTQSozEfwOwTdjwUM/jd
PwbVHfKNgfNYkAPp9ABIzQwekjbwu4oXgP+1sc+k4Wau2R0taXKDFu3LsipJnexoFCvw04X1IoS9
BqkIJuWtfEJRAzSvzACr+fvnCPtsNEt6LSOwFtEPim4Iy5IG2EZThYvxFy1CMrha4BYmCnvKiTZb
TNuQlB11HZXkoPNuYoTpvenLejz3dXID3hb0ZEdC+G8i8dKVXIbxr+ajlR2pRAvWX53SbAdFVdaB
XvXEpSHpCMhMNFcMQbyyIt5/0fhNKW8utdEWpP2vrayJ0SQevSrkAVGNjc6VceD/uMHj+NtAziPX
+gaUES3D8hAvQXnKnC01ak/dTrJrSoe8qVcNFNTAP3GayoV+wyRWT5+OdEttdQtfJMWulTlSDHtB
9k1FVAv13dS5/6LvPBS6rJZVB4grzp6XAM6jZOVYhFItm4rgovTeKl3SaQgv3p6ktj0uB64riItw
0N8ZuaO2tlGDR6nLA/x1vUwcnHAEZHc5lEq8zF46D8lAkAumLMgXo/BfE3uqpk9m42PDArYfF/q4
Pox7IimHJ5CXRV25gSOJWrYksV/r9UP6Xa240Bc2WaUEqISduStqlnyxllPOzBR9v9yCzlwA0OD7
mpwEJsrOGmq3puV2QvJXqhYQ2IUYsWwpvzA7KOYpkASCO7lOGtBearccTA3Ku9wos37FI26wmGtR
94Cug6zR3HNS738nbHyEblnhMBvDB3NoBI1F4xryQzT85zfxiviR6QtBdxIuVToj14Zk3sKxI+ct
SJzvact8+Dza7h4+TV07AcMNXD3c1uR6CvWT2tHY+Oqi9meHWJXQ157huyEQc4p+WNxEUFct5lPB
+1fnfL5tZ/l8LFaTHLIkEF0VtWSdiQgdb+fZ5RvH+dqTv5GU8BVEJI0jiHieVLfSG+J2/kzMkffd
fPqz6EFtsBF5GDW1XUSV8AiAUfl4207O3dqHWDdvRLa6fKeLDXZ8DDRHMJNQ63CBf9x8KhYJxXu7
lZFCHvotcHyArWr8YCrW24PJGiIKcdVWl52EgXwQ4/NUBZMGjMr9KlQvSMqHerlbyQfgW9EYP1GK
+CM5CRQzSF/mAaDtO8lCzxzf+HKn9pMk+vA/GZoSpihpkIwlz2OMw9pcwIQfyMlVtYZnRe6h+iOE
OtRghWmNJwxkUMnEBP10PdksPbU8T+dw1hkKreJPxib+6iAjgTZwriH4t+Qe2Zhwi1H0Z4CMC5Xx
EXvetwUt7XXhbPM3Yxl0kzIKpk68W1MGF+Ym2JQLxtTxzaAnYmjPda5e4wnjxGL1psnNuQASmLes
8c1ieyEPkhOA9CATT2v7YyWeALtl1fl0+HzPh+wlyWyQzNbhUaM3mBIq414lA4JM1yd1upm2knvg
3EdcYzZPAZpV7xF1lttoEeq/Z1Qzua6xKxVTfRNv4ppF25PDt1gYEf7bsK3k1uKtR3+oAa9nBdat
uPq5zvKHNED8T8h5l1lembJdZC9zqSXcPUu3Whyv4X28HKjUSsOWrcupwzfbViVYyZmI6UIUTTEa
oN88bpidf/cwhZ6fEC4+krfdlm9s7B7Xo43qThVXdUKt72sM9KKKmUXIkARmYaDrcQ1oHdDP+N+q
ptC/+jnv/+ageRdMxejI6RR2xezItMtX5X64C+iaeXHHtT/MGnLSRw44qavE/Z4S7hnopllfngmS
Xi0SSkGkj4H38dHFSJCiYslEulhqONlkQtXlWN4RRSu76Qb3d93tHBLDeDjQIv5H9J9x3RjuWRMT
yq4bSCelrr2F+3BRGKHGHLzHXnQwZj53sLjXCGf/msUcb9wLub5gnfO98Bs2jXLl7UF+n5VvDxBJ
1TgcuHetTx33dV4qtqVDkTuxpoSnmkU6ZFtG8FHJbakiNY1ddhDecwuH3MXtS3NItPBaWo22O9Zt
K89HmD7r8E4eccsILv8/Z2Jcp45zgSdaMBEvGWRJ0Otptx5aU8ITo7ABkBbsqutOV5W4C34mZYME
Hb6UFIsTomZ5gKPlDYoaxF0nxEzs3RE9pOs7eBdcPYbeabbXBdr0ZMqy3UiFr4oUKl1qqoNhRId1
PIYlM/e+03s9rnIC1eRnu05uIj7OdIatsW3rAQnBylhocUkVb11B5mHtloEvoKnf141jcR9jl2AW
vVOfAxabFykGE6SL5+G8vTYoUIgk0AyEy0KwMn0sBQHF/C7QYyQmtqUwwr6tGiAeYURsvgY6Fzts
h7/KwRVzp7JuCisPL6kagNPNpR2jQVCGSP437NsDXqcbGT3V15wmME5oWQxF5B58Vzz5DNF1dUnO
I9fMIP4aJmUslYehF0TI1ozwjvR4DRbSL2RU+ulGMsVm0EU8S5SItlTVFSr8YT4qjfyHwLHFFBsP
O67YYiElpx0M9DfKKc15mpGl81EKwaHdXe12bqoh168VXCqgtwOBvXKinktQH7R6i51HKqH1raRy
9GftO8aCKsgqpx1UhXfwXwX5BbRu7d6BNQsz+0ekTcvxM5vVZYGhS3U619y6vSpPon5fSPIhlGGN
z9zlvT9CH5T5cZzbj6fjq3L2N9Dbr4IVuocLgt4mu323cDcJpO3qBbQXUeeRfwBQuTyrkWq3/2UW
0Viix4Pg8jdcUhLJ4U3xsfnBtIcJGh2iNuTJR0kOmRM/TzM1zSewCkUFjiTe1W9u38YtnIAKIHNQ
0FFGkSx5l/r3yz8EaYMS4+TrcnSXq2WNLHbw5l+L8E4M8W2wBIWzji4DNUGSOtF7FrkxC1ClO0tH
9+arZ2qGAcR+kWTYewK2Ar5zqD0EHSThLFC2VzN4MtBrfR8QgY8YgDc2DHO4xebqIu2ZP34cgG+e
OE6+PDFQmd6HnnDDFzdbxEahItFlDyCs1cRVwwsW/IxcIMgDD8Mxx8Ul02a6fX5GtqXfTvkuCHhx
xHMFcMoXz5Iq++P0NZC8nHGE7JKJHtEJCn7ggFwmvks+CphlqD+uhtiqXUONuUb7Q7/TLC7zS7/9
UBM/NymSJRVFVPy51KONw0phFUlqZZ1KKVeeGbHeFOD2F6Gr/OlDELfwXokFVU9oDNG2KFmY2ijF
xkViEU5VQTqqOO8RHU29ZXGU5rnL4Jf3J9lU02HiPSTduZBqNgwp+RoMES83g8CY67wDw+8qsAaw
zWLj9UMAnD9Dze+qkjLaIChc+9dnPaYmfrIWySJf+fKzd9dulsZ2NLIStaQhyeyqTb+CfedRfVE3
sUnW61pmIo0SzxzDfhEmaWkBSyq62RQirc9h/0gT/HpGauWETqMv9PJbnIR1WAKA/nTpLPmTOcGo
/pjP7hEVaQYfJh9mN104kxXu4//qUmInIiz59a7NW71J3ckydHhP8iaGAI3rMlCN+tAant8FPIMC
DyD2WHIXOUcseibTbnhk64B5VP38MHtQhR8o6OBaqo7dv+UZkmMyTuoLd4p9wPSuckT240wTjleq
ZQ+8qfnK9VPL5c2PW0nQVPgRM6dCJrBw0gT9RR3DHFjo7Z6UrZ4qQVvwfFZKanAW13z63AfMwGgf
3SyzDdN5PKBzVM+GIp6JmPFX4yCsjmbYKX3jM5fywA3mDy8TgAxJ72ja80RB0YZoArTqQG0C3rBO
qj4LNs+ufCgGd/m1SPpimMTrvGH02Azym750nxMrlVZcPLcmVHKR/GsuSOpfUdkxiSnwbfJY5r2Q
IfDHTOLn50phzwWh9N9ZwJoUHjqMzHZK0e+C8lFKMELQfVCvILgz8b5boJNEPLb0XBxwF5T3kHAd
QBf5EACgCvya3cMx8yBJ6hilTJX0zVOwzFBTsgHIq763cZZfk9CvZBZmM9/MsJlGxa9Us2RKQEYV
9P5YGFUyHwOlWHlf5MnzNmqcPd7Zuy1n1vcUXY8AmOXX0aaMzoY5spR70x9zyh5P3Y5DJkx1L2xT
8vBMUiZbrJGffkfhndg13cJCXUp5eUEgMR8bTw/YivSQpFEFbQHUmMaVxoCU8zbJu77NBKzf+brL
PKntL8p3MG0VLFEG3MGkNpLzFzJOpEZ7fYZ7ezpAqo666VhnDaPQmb6oP3B2bTPZHzAPvCLBe26V
zyrTBOFp9WJEPAiBopeiaFv2YZyP6EUk4X1wDxGuDTnn7qnkQpnl0uojk0viqLPnwhkCU8+AMUQ+
RdXB4FJo4u1dRcdKPUSQHvBRoYxSkVZpl9hqJsylaP0waQRx3eXXUKxo7Rrl1AymWBMf+Km0RuuT
avB0xNv5jLBkycTFs9t2L9tIC6V8wfp6kyfgYFmbzDclwczuxteiHIMP8wjn2wwWevLq+2LTUBbQ
Q9L9PpjqXY0SAgRd40zQD121NdTo0oHzawy0eORZiPTCagmPdK1keCOIiZqq+pAlnKfXHZjLILjz
Ud88cg2LYQVYBjRY2ClKcNGSjx+DD3JfwEsKo/Wjkf5AA8WK9FSUBWZrHDk2IbE9DFftx/LouDzs
BqO+gx5OKrynZbsbzvzDez2oePhinuz+Pmzr2W/OJZI/bHa+GOeNRjfovfwjbM8UJ5SsE2jaO8O0
WYc12RDVXObqAYh+sUibNZ+QwsajqPcWqJHHHUpK4IHUr7PPAIUAI8N+JBHDf1muMS6vQyKFB4tL
9WhJ4xsNPiTNkchdRpjE8W/RUMU3omNaFq2ICOLqUZjbIwa2qvJMzHsIp8Lo3kOazeuo2bW1CNfm
DLO87icKbmqHTsKxjqvjLQOVylSOJQ6g02Z+0Ok17ft/rmE83bIaEvXdUKxEBvZpzQlqzETij5st
WuuJZ3Umphemz+0ldwc+uvKLFQrR2ZFyrQRg33HLE6QiXMtr3NPkuDjPjOjcfaxrnt9BsGJSw70H
RJoqM/5NEweUc+oXgOVc4k8a7SbhHjx4sfssm7PaCGBHW43ZyhWMWR6zCbh0ABhIi7xGYkhrwbMO
l3kF3WNYKbyoOCWZzG8Gd8IKt3QjIifbJtzy3zYx7/y2Xu6EeVRl3s2A0pviyjN3AnL/aDfcIPUP
zFN5qP1r1V0nuGadVsxZbAi+L1IISvFZZOAlcVrj0TgoCO+VQw8K4ovEZU2ptzYgoEgs4AMiW8+c
Q0BVoY25Dw1RYK+plmhuikm+cMNSogFfX9xyzrqJOgd8ej76912l3pnFy/VqMUJyc4bx7VosQ8RX
l2wdxCBgkg0fL2FER8M33pxr2foX2nRsctV8w8QbxS/7hVj+3Od5j5vdbjsVwwvqWjMOG3nKy2DK
imJoEK3i4MSrqgk1OmsLtV5K/te3PZKG6FvzZGQPH+esqUVe56oPwj4s2BEHOY+mgPEr4tHxN8p0
l5qGXlkU7zBZ264GNBKbd5h9xzNybapgPxz3lPTBeRSyzCmObqXHYG3fdq/wiJDRBv6SBHYoNjHQ
/KPbXM2LquT2LAKLKhtg7P+JEFrqDrtzTLKfDB6g/mjOuyKKNntqlw8qZpi25jLWVfIMORZzARzI
Enw91orww/ZyEC4J/LwY3YiGlCgu7K+67bQ844u0uRJZgwEeNJXWgAlBwLNKyh/CyL9v9okG0pcS
0jJzNg2G+cxiXexyZzMEO63v7ANwc02ZS8aojFQTe0CgOLUwVV3AdfSTI6t3ZFikd7VQF/Xl3zVf
HiVd9TV3PFu+h+E1P8Gd+sq/CNdVJcpebJ4O/zNpoRYtp4auZtoQeKHsnEuOpV7u1VCszJH+zt0n
pDJbSNUbQUiUiWyNee1hlNsjvQ1ntIw2DBOVrHleo89vRKvNPSqrU7XUkdHEjKsz4pxLIopPeMyP
oUchW51nq2R7WugarKAQiAU2d2lB90i6YX3zdpuihJezzhUVWWCf0QZgXN8ukDX7o6i1M6a1KKif
c7A28t3/cu3Ww856ynepDIl/iTqc4gfSmmeN2v/M21vhFvtSc02p2suCsQHJjbmj0GHeUCAX4GQh
sF+YF8SB5g5DezizIunVF9o0z67BQAwW5WpzcZcBpiSzUPSyioz8OONYPaqQw+gsPuCvsUHDSNg6
TQwfIrxGEknkgKU1Epf4NwcYNdRnpzlY8xdHpz+GG7wPysNuG1zSyEK4UqiFn6q68KJPI2PtaIai
BRZ3DJamH0nT5snAGWxXxc3YlZPQIBHv75mqkUF7XxTEKBXtj2S47LvpZMWKEd3gzCOehyOxJ6KO
1rUJGJtMjb1hZutdURre1mGc5fFietMZVdwazKInKl+Ct7D7OQL1oOP3jVm0+ibZt1kNvAd5YTFj
9q5CiMWk2MJUrTZ6MIQuARsDDDmmPq2hvUVDMFBBfD/b1ShbvQLd9qBEFabrc0Gmpz53AqsVneLV
hXhcJ/RzciPOoBWjErdin2M2Xs0wiiP0dHypwHWkbyQUh9wvX7t/Z9zNYrw1ChrYV9YwvycCZTqx
7pZaCitNkpsubFoiF8U5UDgGQJfem0AO/jrJCNnBARc0uLyFI0UiYmr4Kv0VpeiItNVK6YtUbt/+
/L06QN/vAcFi2dx3chRv0cJ13d5eeI4Zo9jDhCa0V020k8Pi7lM6AGIUK7gcioNyBfxFIMBVXpxU
IlvtizluMmpOReBfofMiJGm3s2n+wjN+aS36L/+9jbVFXQFLl2TmddZAdQhLC2qfMsaY84ecxasS
5jjp2OmzhKR1POCTCU0HH0WJu79Rcw/ZQrtcwbWLEJpVuuz1WXQvkbFxrvZN5ob+AuKYSMHJjwT4
NRD4sTVgBJaNK5MqTmFiF9nN2XeHAJZwF51DSC5SPdq8NzKPI5fTU494obNRVQo6yawt00bxZZDP
zijPbdYUQrMZjINmtTbJ2lrFAdqRAquBVuAdCv7S2lQqHumURXU2OjrwRG+S0d5ZtQHnXiFFagsS
dA6fiJv2yyeSlhrsMTMI83BMtPHRk9tuM5yNO6WkWaUsNlBpNCodlfN9KRdphSQFrNX7awOldi0f
bgJCb2kelA0H5npUrskuCSzkR6d1fln2rexSn7KSULoJw+QmU1LScyEUJoIoJ0M23pjTvbaBvwSl
RUPMnEoEI6VcJYlKUZgeRtfV9iBpoJy57oW47FflNgFsa/vkhZCLmJdTItE6+Cif4fI3aU54Vd18
c/rKmolnX0sm64FTdu0qz6GnCAOj8xaZtFeuXTyzf28ICpSHQ+kUKygfD7ZvZh7gJr9kNJ3tBvC9
dyanrmMp2RaxFKKsKSZKQQGDhZuxlOcRJ78riFXrpFUR69GuFsYeRrrJ4XD2wahZdoeKO3k9k28a
KWEbdz2RdXnJfbl/T92+Yc7kucwnLE87b8dNO9f7V3dP7E9LpZ1tPqAygIQk52s+Lf+bmlW689iy
UUnDwLbZ+MI3n8yc6fz7ArESY4FsNsXrJQvSLSS4oTgkGS8B1HYfD+qFeYmjKrleGgIOjfumyiPQ
pe9DoORvUZ01LzVxHVRlXFJ5MmzEZfrGVsn9+wWN2nnRbSTDRNOvFnYhN383ud1V1oxMrR3j2xUr
qvDY5lQwD0yKOls4uNG3ZjEdjrHcN/c+o/QGv/eQjXYRcoRJssMdkdFA8JEY4ewitTw35H7K4Fis
7f+YESptDeNndxRMkJHID8qXS92DKxnTn3281Ns8VfrgCW7qwKIhiBpq4xSZE7vD4TO98RpQ/FRd
iBtV3lA3Jt9+9+rZvDd+jK9CHqi+1DJsbgyjJUmkrGortkH1bnbqAKY2q+3SWW4+5GnEkv6UxSRn
dvrbCrzrFfqgO8mFm8RKtosMuhfaTjovzIRu+Zv//bay5i/Od6nQPrUOj6Botw65djoAZ4pKub2W
SIUlJZpqusOPbvOBKuPGlqQEs1TTCizRlb0b8e14x8ih/7oHSz8oIHDyzJmQIhdCxRzQ9kghJRQ0
aEwJfdVwVPbSgn8ErfaKHSfYzqmnv+iI6h7fFPnbEVwhhLn/jylioWCUUgLJM7De5vpolxey4A7m
T+Dvr1vHQ69TPXOOarpLJmDQVHlTSBimQmxAC/aZBhfdNggQ72GrDaJ3Indq33CgORT5/ctmxzKR
ig8KNRKs1MZbflppDupRxjXZl05yaAknpkCd6IDGCKt9wYJTaDNiaBN1uZsLfMuaF0EiBogsq0lA
ca6U5HCcNejpVTzoUC7bdRC21GWQlSba5xWEuePBrMpTEfu4S+vpEv/VGRlkDoWca4MF8P3jLmDe
U/8FU1tjxTb/yWM/JTXcuh3mu2NUiH6cqHc+P8MM1pWkIHSyhHSaC6+JIH5mJJJ2NjKMRFblo9Q4
0ZxQwHqKZTwcBS8mXsugMKEqblDJevCXp9yHA+b95dyxxEdlRJLTT3TEvxtSV7Bt/WUxhQR/HhX9
t0srGQcuNx4CgheZw0If3qN2qkZFKVhZLh/QooqoqdfZIzJAKjP1+F9VMXss9HuNUgjSMG8CQEgZ
a8DLeP9PHApcqNpXjgXlcXX07ws/6dIAM4H9wVTLNI7mFdJohbCkbx/z0BSbmQe4CYKOI2MURXwn
80rqA0pFogE8AAhxb8ll3ACfWMeGTHhXveQAkxD13uF9gFVvHQtW8zdGs9WWCMpZdQu+rap0hT6X
q1pFLdebLzfoOQ+8nksL8CEhGE3oDrM1KA9hF839UtQaLYhrPVNpLR/LyZYLxJm+rSII1aNiw8mr
CF2mXkL6pfmlOPIUlbQP66Va9ocweJPAn0knTLYXMRfg3MAbmUrAvwrG/2M1eUlTOQOt3g7MP8MZ
K/hVYzLYOt4K55WQGSYBExcEGQlcbu+uYVRY33Tj8V/xeX5FBT/7PeP3jE9uYbWY7ZCmKCDdpfnp
beJK02o3Trm40GHoNaLhqerXTaJQ1hn3orh7jrAL+G+iyc51ldQOUavHxhawozu2wszk8ajc6dnx
zheCb2dgzFGfdzFoAktEV4ygI7j13CeDMVRflB8B3yGH6iBKqIKaKvQUUmZ82XAr02X89KQ0i/wH
gkqh1JGWwuta8nSy/HX1wwkD76TXpj8FwXizS4HOPftWqMWCFJVhUNRFlhcwAAab6O8e+jEKy/+1
Db6ZheN+cVqv7fF6pzPpom3pPPpBDcHSp58Who7jMBHrjDG8yzJvr7opml/rrVD0OTKOcQ3II0Yg
Jqzv0/ZqYXLnd7tU+pagDycwl+mWE23CtxSIDqBlKjx9NI/HkPNfRNDughX0sQDlgy+48CdvwNvx
gL+70pjKrz6jAOc+o10d2LfpDgU0G9LwsNrvHTsKk2FJ32s6sjkS2nkfrFbvqPb64MNOjs1EfHEv
HO2J8iacvF54ojtcC2tgHurPBH+96ZFt40bw2reJRKDH9alkZE9fE+8ICWZMhIGjgiUxt+VCmp34
q15bQx9D9zrirQ1b4MTkGpdG1LG+hyZTvMegbrES5XSBr5RBkDMNW4fflE1pEqzLUKc+RcxY1u5s
l3HWc906iwdSCeOlLhE9nnpETHsoh5hJKnBCKJjR8mXL9AoODDh/1VgtGJPgtv0uFJhjBu5xcq86
a6jOZ2yV4runYaWkXcjxnHDhUVndCXqmqQkjPssYa42iL5xBYNDS0YgPqjw5cpcClfpJW2+6xGPP
aTkBnzV3+EhyXlKa9dN2ZKiJxCsCR0nQRSEIN/GDH1uRl/Zd4xvI3VM/kV5Ubj9Zux+KpdgmF+OU
aAWOnKtZvwd3jahminPkOHrkDrZtAh+oT6z90RrM2PN1rp/JioYgSucXFaAi5U5+1YKlxkScOwn0
Zg803+RlO1Ukaugy+dq3VTE+IDTGsUZe5v7KPCl2H8ysst715AABxeJo0Gqnz/8h56icpTWcw3oS
3cMKCzPJMhhGb7Vb3tUhL0iFKxVhNE/nz3+wjdXF+0CdNpVPXF1N/aH3YL7exn35Ket0NsbCfwRW
60d4qb4/6zDwQ519gO94UnCT9A7LHXjDoLAfZ8I5OIdqL8VHv2UXm3lE424p0iIzjHE83cyxJP6P
08Dpf112P24Yy1J9hHK3VQ44ggYXHMmMlHtygEJP7uiE6ocLJz1BUYn9+6xIjlH49UtL4c188ClS
dtM9DZuLeixc5XVct/BfbkMl1w5brvvDaGbHFjtRECn1KxVoFMn9Un95PSeK8EFXbRW8vwJVVG7t
O4b7tptOrSOOPaOS878F1EyZFFnNiZ7SKcIDBGHmZvkzIF1KYx2PQixP4gE1zoG+JgjZLTQKgIfH
b4+40OVrsSepZTnap847R96XluHx5emVVedTlH9j4lLB+ir5zRdCQALWYeCZKKXyoUDpf19BuR//
s+STnDeHZuoVtRlGaWSE9FyDLK9/H6jti72/Zb/MFtCUuqskcpahdFW87rxpV+sPssu7zIHbCMG9
xbrF7xP7OEkrV8HzjMEidd4mdJzSQlRfOAJgmI191t9lOjHz2niBRNPHx43dSTfRfH3hIuUg8/SW
aSrtY1ZUhV5WxP1xaOn0KCuuJioHM2kSPuRwzzBmP7IOOfP9VLJRK4dRoJFZGWxqcAzczUcyQSEN
zwMlSi4zZ09y+J8ZE4qIjhZLkHRdjP75o1jZzCrLTBYLPNuXFp0IDn+ZWlzyiAZhDnoKZl+igKko
KNQroWwdUMz2FYKVYjc7XRBiOPamoem674M6A+BiKzMSw+8Qg5FGvKGcmktGU9sMn1Uq5lXPqh1d
jBla8fAlLC/j6NullpDP94+tYhImLOZqcFMWUZxWmlxrLNz3L0JzlgwGdA8oi/pEGxE7FX+9CoU/
mxRCIma0n8stvh+xOmK0XKee6x+db/4o/lG8ge6IGGFJfGalqu1r44iGfoMNToEVfza2pzFNr88C
YJFb//ASp/7tS7lNLyJILt6S/E+o/iby4rVNPXoNMUN1LEMvtAf2prjfMq8yNMwTiHkVDDNH4Zka
kI11t8muPoR06HRIoTI+BvZqaftSv0Tik/bdkXKKrKgzKvG4ZD4srFjgNL1F0nlMFwz0RQQbD7Rc
HnN14/yZbSi04jThID8FiDOna6hJRhmhRPI1GK0YFiL3k/ZfqWQoFjqp5xqLUYX657CXyGiq9fbu
xNl+Xb1kv9gGxVPSA5L70la1Ux0qXmFwHwQoJAcGk18/uz3+K7/fdqrOAK/fex+L7MwG+Jh87u4S
jOQtQkdnpptAOMKAWc89x8IRc1ge90eK/CN+xe5ryTPoZ7bS//xgljTE1NPxpfXANled4HLLwSRu
Gk/ACbdyyvOZ6qFt1BJ5j/uEzkhykaJWbd7jxCjv8NO1/ZgzDIiAR2fBI3XK2M5+e6Gz28PW1viR
O4TBb8SsMwcv0wbWBiS6n6KC8UnAm9BhSnWHHPUJY2EgrrH5G2Oku0gvBJLY0mEAz4XNMXO9xDwl
mCWomk7owYLK19hJA9jNKmwHxUljUueLvutNi++JkMcHpcWt4TXt1fKI8gOkUwtcB0QKds1UAgbg
l5Vdl7rcBnI2KG2Byd4MmKS3OrSaqcFAvni9aI0qbR75FaytjacvFdntwgpK
`pragma protect end_protected
