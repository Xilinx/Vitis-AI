/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2928)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B695KzjSFwUzAcF8d39dHtFm0SIK9mPLbuMvjdjh+BJAz138S/bydsjvD
F3qHONzEWbPzXX0geTb6nv+Ge9t409l4aPWYHk0NaOnUvvkhvtoIjXAEu0b/0Mhix/vIRr+/VUIl
L/RBxMqCk6r1iD+YnPySrk88hYM91Bz0HhIl6EqPX4xMVr/IA/fZuvQDigzM6UQFMAp8KYT8AdUk
7crCvMY2UN+aZZgzqJgtD30WpOwBdiJ90vrU0NkZabkiw19yc1r5LK5iGnz3op7lYvl00Aj6QYk5
cd3QtNhdzx6IKcDOzx0MEDUowAu0AQkUUWzZYCWAY8lTJUMNUcPgPrd4qME9bBEZvttpaIAoCBAH
uBL3ASb4W4EujELnSNyvjTDrU8nLP6XR4jh56wY428wL/I5LPp6x82ENiiXjr+RBGhyDAKcSIBAE
UbTKSgAoWk6r9wxDMwR3L8UpAcxMWD3bkICkAMw2mTKGxw9mi3dWrrV0GjeBHDdDLRcL72kjujZa
8Fo6eGhVxbDZy27JrCAzrJ4YIiQBbH7jyL4+BsZLKVRHgQrRV7TVW3drJa2aGuKA9Vkj8zU/S0Ht
wUW55axiF+srEceuRGlxeTdr22igRuhut8RMuG5QTUkQmJrh1CoYZTeYbZT7pVDGlt+Ew/TrNdYn
aWg1WrRRFbsEnvFjWzNMfhOv/sXu/J+voz9IU+pMgjV7oLwBv99SZOW+9AQgsMyWTtQizdQOYEOz
miyF+BiImZ951Iya2/A3zetTyaiYwlNOZNcsHuBPTRQGYGJ9GOEoKzC3x5GDNo/S/YQaL8oCKt2/
Y2gNdTds3QKFbwChUk8N1/2T1aDGFJjp9M1jf99RYuSPCUSE4V/VN9VKHbI7Lv9D2eNz/ygNlJ5D
s49T4eMdmXrvVo3/L7ZizD1lf72RNlFkusYHO81cWHYUhhlg2CgfNAATwhJV/TuUCcPTJb4qVFLu
9rQvtsXrf5eSURnH3No4uTWDpCUFHMMiec7ZM50O479AIq/QIHaUsvJtIOXKIfi3Zr70HkeWh61+
Fh4VfqmAwFnDKUWxPCeGXjYDgxaKXgCa6v8g2p08myTRaicaxWI3wRBlvyVwuGzbFBY5UYBRTY/G
FDNsFhDQ6rBlYIfdx8kSu45xGmbbPFBsbXFMHa9gEDWT+AaBBJpOyqDSS/dBE0pAuFMOZaz6A5te
u26UKNe+XjeR3Y6vhYwLro0GNZ8xHeCacMgOk1rwsptKNGj0wdaEEjk1oAYnMHOThYQe1WO36Gmx
VXOC+JfeZSzfeOUrPv8cf8rOionUYw27wjwPum/aUWmvj2Cl4u5l8xiyDwd7sVHG9U7C5FmzHBtA
o5kJWUO2tCsSl3qHaaBmOZv9YQKEOXwnF54OcWlBu/6tuyGWJeW9HJCpN92Tn+k/xTDd6lEKS0r8
fcvT80VeL4iIEmOTT1xEzVMmjzCgtuAPF6ueZ2ST+BmT+OEZ9uy2un+PHGGcI5XPGk5BbCDQ2KwJ
gc+tEAhOl+WttpCzZC32s3w9H8O2oVNdUpoDU5kVIY2x7yyUJu0cdKB0L0t7SuDXnHCA1O/bOrkT
CfjjDQT9PJDmrCwiesSwbG7d087doSDVoM0k9OcySu7nQuWggI8qwqzPq1jdpUGR0jvoEDE9o4ZZ
PSVTD+11a88ufSzPQapUI717FS6KZlLRLXm+JagJnHCqlfMNQSC7gXpIekOLutTBNEH9DNfr/RVm
mVPdWT947/1RkADSkX8bHmUVGc875tF5Kb5uQtikvVZya4+VN8CuVetxASkycQQ1qwVfuo8dCZVs
G2MWNZA0JPC7Fuf96NYNJTuNJrci7hHXk/HHuichVhvDf6lAjgMmYcIObhksOq/bK99GW9GqHgyM
dFi3qwYomlk4QmInQ7pdKRiQ2/uGQXyxhj9ffdKiMDP5t7mUN+czh0g2m7eraZx5UYV0H3vTwUBH
85xgUulYaPAq6qh/YW4k131KfnWxJZfBnyX4Tjv+7ta6/j+7H87Jw8L/x86lrmuVKEk7xGsy/Mgv
Gn3Yph2wAgD+XsLaK6JnKUnyQTPR6kLq0BmfNyVTpJhoi6KRo1U5taCyBED4fVVecef/ZYCJIiAX
JXWMKKhAUbhtw2DwC5+uOHW8+kJ1XPLQv/chqR04QIinKUl4JM6KQp4tezmYmmDVgkpXxFnhjnUH
dSnJUHUVwlc+QrtZv0mV7bBisTzRJlVqcK1J7e6M8GUfo8biP6Q6vm8R0kPZmu0SAtqiSQWWrmur
fUoC21mZaLFzuYvGtRCgtErSiSg15Wy1htEB4YKoPHMyuwoRfuAkZ1TxREjq4IaUslgTk6QsUMCr
w0/CKIZiAJW58O3ulBAyzloVzhMs+VLiyouImYLt4ukeob/y0dyGXGdDDuZInDSPgenZq/3UvA6V
+sk//DwSg8I6yA87Zqciwq6CPkyDK6+eHh6MStntWpgNr/Wg5Jo05dOzIq6RPtekv5rbFlGjvF2A
ODYdaOK2ok5w5HN/ut61mF0PSzZka27y0yMfN/BR1uVP3uILUUsEs3OGOdxAQpXhXXtvliv3XH/5
cJXsxsezTI2qDcbRJVO7JwocO5ZTnFAIHmLA1W4+r2TSu/uqR0D55sy8QJlCNIOqQ3Z/Xs6EaNLL
CB/UAXh6zMGjXLRdQ7Co9pmJbvjpjMSoWutSfmcYkjM3MDpvYQH1JxOwo/QkUyaoOdwTthUA5c2F
Qzdp0p5CUw0bhsaxsNzfpV7e3yBJtViage7yHLAWVS7Vb4nLE6ITh5WdCu2Vly0Cj1PzcBheres/
9FDY33wnc8hHOqL93TLMVqzmajyWES8YhvIR6SxG792Q7c9FbuSaf8sHIRoGQdzEFXBoVugm1Iie
iloPgy3Uj/fzNYBTjnKftqcg80XjLivr1rCPN/EjOtQSUFP5rvYPhuu744Kdoq2D+t6pHvFy/0h8
boeMo8Sg1acfHHL1sOo+EpggXLoFTZCwVFin+s2mSb/xStkVZ9sj4bT+1NVJhN3TmBN0My6YMmV9
EtoMib+ncf2pJebuB7Pr1cMOCH7Tbbi2oAt7x6X3ANYVqyLs2Qbyc9bBFkyCNKOuI4cBa6uQruXR
4Jc7LcXs8+fSnqmtRv/lEYq3Sipqeb3PUTdlyLIUWLU2t+U8GYdPxOHh5EUtpD91yp8iRSRZOvIR
IXd0OmEP4vzMFqzTE5kddi5pq1c4jB0/d4lWoJ5pJX6OeroCTU2at6QoCPlh99tn+qBtH3jlo7VA
6gIVkjhauIRiQXhicR8KyqBNWnq9k6r8TKjSs55Yw74C0T0yKizKYCZgVhbVkCY4TX8UJ8juvaX0
te55UwsfzT5JctuMSt52kT+N60PD7xQoIp7fBb0wlGS2+FqmJf6yKMUhTlzNqsKAUWnaCjarLm/z
4Q+9zEDcqjBSUe4kVUeSAIf7NNHZrNGLsSYOg6PzrdE4tknpoG+CFo/ETk+SwE1iG5G/i29ddAoj
llaT3/asI1vpaclMpD2pADma+eK22Jjs6c01q8JH0ZL2yjNTodnRdTg5q7XHeNvPQs8C/whPOuqB
3aMkceKNUAFobtRBVI9YQNQs1Z0XOS2e/czp5RIcSSuNA94hv64dcBe24QE0PKmSzoWJrjJhoFIu
ZedR+yulaEuaG+oDPTWYL9neQkOziSx85I6HBqO3b5UZDhKQNuGcj5rNGINPG8Ps8sYmurGXUH4y
o5PIrpwMu//aTgBr4xAtjP42Aduh28u8eOrp3VEboiZuqC+FGJf7mBMPVZtptZWTWeAedzCTsucZ
yEjYXuHFb7N25pJ3herhlv1Zsi5uFXZwoC6OTF3k3ohBI9uMcikCmr9xbKmKK/iXLD43fUV5KObM
da1y2VHsDI3Fp5zyAnQEHc7Dl7pG
`pragma protect end_protected

// 
