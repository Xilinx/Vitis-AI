`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRkcajQVnMQxKjPBaLZIaR7/J7zs
kEF1+54ixDuIyNX+QBxUIanAUk7iqIQDed2hUG0kfoXoL3vuow/GsZ8M3G4iHfWrH7YjpZpxAU7u
+39ASljNjmhxyj7sp43zFjND7KB7yDk1EnS5RQNQKgSwY3fvRC0feceeFHyy9eiKM0+E3KW82xi5
RDh2XoenLekPW3PgKxqpPoG+gCC21CBlAB1jyVhu5giqGNu4bAVf/Qoyy4ljAhFmoJLCZWCvKUsi
ICv2MqFHKqIij/rlUrw26VvJqgt5PBxqKqEY62u+yEBRNPG6sBwAtGfbLTstjzbQx9RGnWetL3bn
tduTwLnUXWim02JwoBrLHqTyHfGqo1ZPrbw/rsudPnmprcaDCdabcGeL4SAGV/8AvSWW1oCL2nYB
ezoMlPApKZgWMAS8XHtxytYUrmcXEvn3gMuaYD1UCVzw0jm74CbBuqZecCGyE+iD+aQQxeqi9Ba/
dvff1DXdP8zsoS7CupsEnOV2zeNlF7/+OM01Amq81zXqaenFJ0zkRZg1y1PXmj5QCj7V6ucaT4Ut
7onldazNSYfG/ENwXbamxY66wHxdxp0YxKJiHQJAOA6/TSzpzAWbvPi2SQqlPI1lphuJ2VUkyq2k
TREvQbcbC7sGduS4DfCZZJ1KojOD8cYNdedhjTo4nWZqp43QK+VTlLiAw7kp4bxjDS84dhBBHPa3
9ImMBOlkPPqJlRbcfTlaQiCiQvfNxbK1h8ixO0ftq0lUQQxiAmUmMwXIyADQJK2ZR5UPGr39t7Gg
mOtF1c6pgpTqAn/duzun1T4DixN6Wbrdfw7UxXSwWm3q200ba+stIk7IRLRSYPBcfezOrGonhnrb
OUJJpYJBCAQjZDe5hYpX0kI6gn8kA+uNoeEfRNwLXXZe0Gb95jZI1xj1cbEw01bHY2Of2BE5LJFk
2NbIQcOgY0SDcbF5qU6OBu6PjrzNd54MnwuYUetNGVEzv1VX7TLBVhS37v6NydZqJraV0JvejdYG
w8f3kCfRmArswcNfZ7pJIhas4AgpJHIeFnR3sDyZ5R2N3TF9CUD6O4/+nmWIRl9QsFYUAAwpMW6p
iK8ztzjInBArmXPcHxRfORIsWSnxfiDb45PX6ih9HXQrjuJE1hDsc2/H83tx7fnstNgVCccd67/X
lzr8n6XZnaiDIh/t0ZYkT/4CR7VdTj+ehRP0ViIuh/eT1uHmSsEJ1Xej+0Ut7l47Z9aCZn6+yknd
ISZCV8QZkDiVQWyRBEO+i8CJhybf3VMV3cb/Rw/u9jJfZeNzVJlR3HvJBRbAfhgRkw6vncidtKFf
lVbvtlyMz4YEZAYmEMNK2T/5u87DyKRtWGaKryJ5vqpYWVNt1nj9jVdD6NL+dL5MSs7w6sLqakEB
pttg/4KNfLTNsZYe0Mf/Vl9cfYUDH/1nY8nVteZrf1yB6fbdx/cqgsddxLS8cIj04xk8QwanOrrI
WlO705pbzJw6b+uvrem03rd/Bdyu4VCRkq/DovD/WDENG2n2XBmqgOKaYN9w2v87+lMrNdzoloBM
PpnEaAkYOqvCIzYcZnhI24n5TNe2I1Mrw2/SgMdHbdCIfs2cIFqVDkowKBkbZ99nU0ZSdGVB8YWg
HDNeGHWCT0QDxDEp85KUZPwqpKnWY4cKhZq0TkfV/v0UdOO2MrbTDNBDQeDpOZvrhA5TQXaGTSCF
Z2kq5GUXRx9Ua/NSX8NkfqKr6IjYEAIvv6o9fSo1dI9cRVwD7odJII8X2BNENQ93xasuRfH9SeoE
+I+1MS5RRvi1/Vc15emgG5qP4zoQR/sOkcFET03B5cHLt28+VtFCrV90Y0bjNbfJf9M0zctGLe9a
LybyZxUyWaZuIDkJWwdCpBXth+YIV7JA6abswTqZpFPOGlWNQ5/gBAw4ArT0AHLrA3lqw4YEMugu
udWlte8CzoKJOiancKvCn3LxtNSb6rKuS0ESplzto4TyrQOIQ1lbsD71/ZbHAG0niHUZiCjsUY/O
ao9FtFGub9Pbxg3dmRO7CQ/SIXpz9+9BpKWxqH71Ufd65kEKCKf7/iBQRBE+Q1nt7aLUsrHmYCrb
UpzJdWTtFknm6KX6J0D4xWfqGYhsz16mV0oESv2KyLs7p7lv5K6M9ezg+0ZKPJca84sN0lH5FTiU
znvSOMwBEW4w+KGPXMQqjk1ntM4xJ1eKqbdFshTGE/KfrfZUlH6dgpUy/So5f0AcZx71iJ3wG+jN
RkwxJou5ybyrDeMxvZk4gm6MrOfGM8cwuTQRBgS/G+aw7rrNRxaGIP2B1ExAOViY0IHPFbuswJiI
gYWcdQZ/D4U2m/ow/ZcIEJFWtd9ApZ/dlHSvcYqmFgueZXpNN6bImbfREsOKk2380b3NB/Tze+eQ
c5UeEOZxMASjkKOYwtj9augsgcHFTF61CtsdIK2f6vQNCW8OtnaxmBJr3iZdEVcK2ULlu+UM4QK/
eDJ5E3IYN4MiH6W4luvomh02/M5l1EYsr2TrP+SrZq9tgxuG6nmHNioGLQKCZI1gXkXGorLy3o/k
L87yad2q92xI6EVbfE+o76uvi68kB4NnemmU4BfaAHTkEqI5dogc2pQ2y3QceNZ/c2bZN+5UEiVU
MJ3aLDazo4p8DI0fZFpyJWm2V3xC/Su50wT6ggAw9zgEr4CprRg8aRofCObQvNc71IaniWFE608i
BqJinEC+MRFy8HJ8IEmPbZvfuhoWWPWSTSCPibnY32vewcgdV7EsuVDdZzUYz18dxt52aI0/q1Lf
wSGI/00oohg+XehDX/JsQFKlaX3xsg2jbaKA1kUglh64pQX2T6xfdxYA+n/Y5UYavEN6VvslMnCH
8jdMYmjk9UeHeM/CK1uAAnkqxQyI42g62F/KIS17y/10HvPsDeqkqH5pDYaTaekDW2jKjg0FSD3E
x7oC6PRjZ2IceCv9cnwVVJonL5fr2Dr3cIyjB2VGXnwTiHaRqj3XwqwMsIor4auOV/8godrMUOAj
ECuoNIiUG8SzPsMuNOZTo1zqqi61pERoXtcOD3IQMH3gAlk1xpf5h8gbb4+MvV01KjVaiqAZGnqj
Pqr2BAhN+24UWt3mEgaExr5C2rUby7xY+Trdf3kyOBx+7p99EZsc6SAbsp5E9wr282e5bQwQDWiG
on7rIcUYHxk23YWQb/v6a6DddI+jUi8cWXu6eTU/GuRJCJ+/TQq1DgKnCMLC6fsfwjtsIwSfmG22
RCbg/zBQKpKiHudqNq8lOPVbr9uqsLxMS0EjWM04fUhe4NCySlFz33hrBisDG/h+XA1gu+IBU4dL
WbCKSm0BN+tMOM8hkXc13ME6zdv/65RecoNMoH7meoZqY+kysUk06UFwTRytjk6w2rcUYWWu5ztp
qOtX0dnh4tzzDrqjsm0MbCacg0+cxqSnnp1eztG0BOkEESVrNCCMdQLl3D6eWYaQ3iaZFwGCqu44
lEJotM6DzeTQ+PJQqU6RRvzMQxPp+SjAmYVIlp9zSf2LlBxXGddlOrE7oZnnwyAi/lmnbVOLEwCj
iT7aewP1PHUm5SI+CPrdcLNNUVDLDTu6cY7ktI5PV/rUWumf+crofvx+9kV/v88aoOJhu5O8fGxk
JPUglA4FFv+fLlTGZi6Vb44ie9gXMF7FlAryLorsi66TYPDkR4frjkTBEbuXNgTn1JHEzOs1GI8H
2Wslei+efFdRLZEIoqfMfxWcPtcPXkUOVJMfx+5zzW4sHGvh2lYykaZTVNyWNEYINaklrTPqg1h2
/3a/vZsuCGWiJmtxhx05Kb5CmxDgPiZ5r50WFNB9oRWcM4OuygUABJI13P8z/T8JSyfXm0jl63wg
nbNnCL1sbo1Ic/DeVoWXbJ9p0ATgKm9oKliLEuuEJw8/VypQp39j9K/S5f7kRi8O5g+eQ4KZ6ivc
nW22qVATk5hAQvbmbdWJRI0wmxf0VYfdOuMgUyPj2sH7BILKYNLHe29lnr3ShL+PYyvgJRGO+CLn
wvV+AkCpXN8nuZlNVb4Ju8utUHB95VIYMuu/t8u+ZMi/MCWMRgAvkcbVIi+3o7iKz3xXj1RFcIsw
XnoKDpp+k6fKvtItMZ1xpAf3dUCygRyLVz0sH/S2hacaPXKUdMZFoSoXg97EzaEXqFypuF0Vafxz
fetykquNjnX9dxev3KZf22OLSRlJRLTKhW7DpJhsYmCI3hEHCbbyQNatIdr1pgaqV3cNiRlDc4qG
vnMUeAMzG9MNWNumOzR8Svf7MOGlnbKiBkIVovH36oLzxoGIssiFDC+hDBv9t9tiMcj8Tru/JcIL
iBk76nrF0Vuix4dcXfuK4l/jVF7UeTjKaQ8lx0ofE5eNAv1TOTHKp9y8o3MgeIDYF+m/sMOh4Dvq
2cN9x/9YSWkg+Q0YsJWHSSjl2ZiVcGFW2xJj3b2Vx5QA5BvMNSZPs4AO5IbVClyi2tE5SxLb74/Y
Fe5whfrWxh97VuJ3TET+KG5V3cf2oT5FcrgKetkHMQ2ZesEoWpnhyVUTcNxXjEhEymfwO4Qlub6j
p92kYIaI7rjEAx+dz9J2ajuZAYf8Opx3fhpvMRk2/eU8/qKA8BWTrJAKNC0NLzHmsLnafB/SK2Qg
o0CUY0R4HYrtetDp/1nXXZ5R04bQZ63z0DC8TtT9EtT2vXEMD6Q2KjNUAL9alzbsKPGzvVnbpAKN
zFd39wkpNC9Fn8Gqo3UylVVZGsQqwPOL8YdQiiGABIHb9jLIq2UEGLsCIzic+lwKoLZNr916nI0d
G/jVM4SjULsluvuoL8Ls9WpmE4Dpjmcehe0bKIsYAfOqapN0v98EUHZK5LB8s0hNIc4IOnSZczDU
MRAFa4wZ08tbI9q6FplN9XOXdlYw7QBYJKxcDiRIOZm1uWVrzF7p+usVD748Ij/WKFhjL9rO/EkF
EExmHeXdIa3D9I1/u7zTxn+ydv2pP+35GPPxY+mvJo0sR5rQhUfBBDh0MZKl/wBjJcoyFNgkmfKi
HZBkV6sh8KvoewKVJpI+1UdQx+gAhqb12yXPAH8KuMt91qf+/1X1Yda+w10HovmkZJE0Sc8H3INl
UdICR10U2iE3/dhchqpcc6/v96e34RKVmuk2HISEg6wBO2CU29I7PndN/QV6BKg5Fq5pmcdajxlk
5+C8PZo02nJhBImF48y5GMjiFjfqUno2ZEQlpokRhOmjKcGOLfV8bb3QyKXavq3G8LCmfNLyOox8
4MuhKUO7blWi5K+5vjBza0M/jWLFZawQUXKlvLc2AblO7ZFJZMmMAOljWyO8/eSusvxIRcMTaxCX
qgjzjZKo6INhzDr4RkmMCGJhllRtla6OScMx3FDon2Mj9Bz8m+nTWNdjggBOYB6VP2NAjQblAePO
noMrOPvpCDT3CDUk+mgomPhxcq2/dBtNF3seHt9LPazzqbadxbySjVKDp7AEqzQOeWZsqiUBv+mE
7YzavO47/HC2E72bi/0se9l0BYzZ0xyCMgVvWrJbN0ggNdbctxnCgDedQceHs2ZT18r09n8mdBqs
F4OQq13IZBQMwyXicG/CL+JrEg7eUg78F4GWOByRtSCXSxeKHJe4dsJaLNK1KJwXfuf4zOGLY7PG
CImxZlSfMsQ3Vz8Q7aaxqsUkiGhguGtr3D+fWE44RKZ6PckfmINLp+KLmyH0h08QJKpO0zRrXuro
PsJWsALhWvu4IV01MX/RBJp/wpBkEWMdZAKkHhrkcYTTetY8V3ZYmvSb1Pl8McbtGm7w8gjbrmUh
c27/laVrbkXiM6YFpHdrptiEAO5PDU0OylEjYO52Fkdkr2Cetho9bXvmpcgUsdf9mqdBtMH+qXvc
fFixhh1uZF/WBHYu21JOIPNH7LFwyNoTNWjwBOQYDNk2EL2cRW/tDdmM861AQnsj49rLKMLxEZx7
TS8QFkM3Ek6Xejz49cnDr1LEMIYgFM2M6Qz4obyQXg1aNdKTsP1tZR0JFxnpoy6eQynBgmUI0eMx
6u48cInWmU2/rTQ2yINFhBNtmyAWWPqblgG4lc2yA4wwr0PMCjnZLEPR8WhNyI5eJrlZCuWJjQ/L
fTO/zjKOMS+t5z8fpvPspWvoki5kiKGS6GG8aYf63q1RwvX8LiAsN0oh4fJoJS2korM6kx5WpOjk
FHTypETG3FCrOM9lSjx3N6yE0OawD1uTjuPfqCGjDH2anhG5+I86C8/e81O6n0O/OVwy4sgHwfdA
uqKA7jKnbiF1JehzXwWLYAjVUkHI/C17fNWjs7nQw3QqG177PLnc9rMC+np4/4Zc0L+7hpAN14q9
eqg7wNZNB9yNoXtok/tbzBthRcGSO4kGYP42SHbUPinQ0IUW1KrEgqcQHXulJUIEHRQF0tAxEhKP
DQRBJO77c5j7eVl80X8iVUIZYTZW95OmUSScvPl83bbfIIYngHDzrc/mAWlu4DRjDHWlbonygH3t
Plz/HQuDqU/+WnwScNSOVG4nUWFUD7jBO7oBgyCd91igCj4LLoiPGc5asMSL63CLF99igA0Mpl7X
blCcPd+NpQ6Is1AQw5B3NK3G+8M5WqJSpohYRv+mv6Kx1H/+a+7l9FI0wsu0AqYXX7ggYwNfawqK
muchJSeQIlQD1MWK76YFLHpugNAOC0QSGLdpzX+pxzmFCt2F8mOLVNZWxhI/SciGRI2p5pfR3K9N
/rDzbqED6gvj3PbCkMi6M5cA8si3os6RSCOVY5cIS95yylh0tdgdXJ9kpgYPWj+ye93bHmu6c+4V
HXn4McbUXCUXrQkzTeWENZVWtCLjnhM5Y3ZITpvlJHbxw5y4JDoikfU+HFaGNzARhk0rysfyGbAk
OUW+htb4Jy/RbqN/xXImK8MUBssffLlPWQzTmOEhKl+h1vb97OE+PzTEihZT/VsbP7ytBMmvZIPt
ObYasiAKZ1kaCEN88PNNCGplEJ87IJD/tWwCNuHtAfPsifZroYSqwDnVoZisS8CI6jLhCzfET7W6
HqF84KPCcMzHI7gXkF+UIgIsZ0q44LdrIhwZUNfiSOnyGYSstwm7tYp8RKZNEK8RuCKpOvCH68Sc
JU1PLlrsH+d8aRvVMrS+uJSyzM6ezg93hKa6TZ301hOc4dZBEIqJUVZpLtMAqFSudiWbbmbBggvY
JYyK2FQ6JAZUx+LuuM3h+Fnp29o4VJLFlrVHNsyFjrBxC4kinZNmi5dCfr5JKUIXdgmi7knNQhtK
dcuo9vLyTnM7N40oeazx/F/66AXgHvVOCydCFo3C3oXrdc4zqkI6hy9yeTHYRRMNReHTWpALhEWm
Ey24lIM+K4nk+2fq8UYEg+3sQckrwmRSnPQh0zc1obqMSL/LdoHRuTep0Zq3veMpJNnd2ngNUSBt
LAM0zThkR3SGVjSKK9MdIaBODhZcV0yyNgnD+REcjRfNPTRy80dVCFKih5ThvcRpgSs7Qo/eGMkc
MTzhzl+XsmrfrFFo97m0bdECWxtb+VjPRUxWuj/Z9xTXDZUYDbvr7l7x+ojTUWXK6n1sXEBX6286
zALXkTDVvIh4FwD51xCY4xXeIgkn0Dp+gtv7Jr09SIZdtvhn5/5uNJxBua04FUE3983zdRnRL1GC
lwhOdKnM2TakXbNW0Wdun/9DKSd6pzS1Q/QBUYH4jPfrP2+fRg/SEIWdggjWB9c81A4EFYuiZQD7
keL3svh7fGWmuLgMqBgzFMbwB1Pwvm5BdOdptj0ioOiO4x8GlFaM/fIBXBiJ03jxO8VZijTd5bxg
1gWyx7PdUvNC6jyto8+Rm2yKuQDz+zQPRWgBDE5y+Jm87as/0DPTh4wAc7u61aBK8MMqmXGAPTqv
aBIRlWphpJWCVkht8Cmi1GN3H8O2m7IXcDBklR1NcG3L0VF00boD0JSS4maMjHiZQxPiqg6KiZ+K
4T/U5be2RL17oXIHLAYbgzuicxBmdzCOgWvDdOKqBVPDi3xEQVts95BAHLHQ+srp3jkniBFOnkfq
nyC1oPfK6ism0fC6AuTCqaO8XhfpnOBeCwygVWwyqX8PFIgRGfmOittjPyhONnjKkbZ+5lPrxtC8
DWPlio08sn3+sd88JpTmU/t0LcA8N8z1zokFqva/e8otTS7XS2kePwE13rcECeHjnwkHEwtzRbqc
MTKpJos65tnXLZRbx7Z1VZWcwVjumFzRj0myNA8uzpODNBHoAt1JZiwSAkDG42c9QtTXOmOmzpX/
X6GZGV0b1yhZ3fl0DjkEK+NlkjbVAsCEkyrU51/shczgV2NQIIaOHET2/Zwmw//ndeDY1L9i1VQ8
xuEN0m7UZjQ/Ga98CrPqxLhmMbue4Wy0JTqC+C60ioy4UQAZMGE23u/X65OBT8wcHpBfM3PJkuex
35pDdFj4jiciwM7iVR4eRN9uQw9bPOH8Dj2Og5G21GSqlRj+10q0aNHADfmBKczF7qRfXSzYqDSk
wYeFJOo7hKzHWvUYDcRWOgHfXD7TnCbkr27Djxy7jUt31uoB0nms4FytIfv8Pnyxy899iDB6Qm/1
jOnIadfGbi7Dkd6JGrL+iSvL/uhmrOUXC1AKI49pCUJXeZKIUN5IdbTtQGuKAt+9gl5o+eeG/kAu
ounqiCcSfjNgnLeoPJdwwYMjkryJYid5yltRIFUV7cF2LswosVTfSrn6ZMJzwAgBNRtAgW+o5vY4
zLc9bz5ucEKGQ+je+9t9GgEpMa4WObf1SUZcSSGzMTS1gJxXQ4E/vhCZvSvsqOTclHDcn5RyvPJd
UWVA+4vzRXg7m7QYXDZ91mW7ylt6J59gcZpsGb62fLIVShv9z2JfDBPiWAFrDhiDiLGYDhQTwpGv
Vbcz/4bRKIuFecyFhXQmGaPAGYL1JR4GXjHPWreFpyBBjuyWipM3u79EUhQtTmx/VmZ5L+lV7JU3
3WnOOkoPDzg6D9MqC3QBO221ugxOrADLVZeZTibFQrnqYD76RuLsN2trLIlpWl7S6/l31tZKpnt/
aXQ5K/enBe8nMeGqHQ9KnOcxqeru9pjlAtRLaT/E1HSHNWYS7ZZbrZdMvyEvAtDqM6vU5DPgfK9D
cxfJMkPcYPg3yKhmDxsGK+yJSgTX8UzHhxjJZp+VLSQ8XIWISvQK0fPHNUkrIt771a5rZpGIXY/r
4cNkhb+pngvC7O327Kb7hqmQcnb/ee8ORVpOIKMWfWAVbVmL/ljrmeeEshJMbZmzW66HNytQIt5R
58z+xZpVhmPxocr+75hT2QLeBPMZiSSZQv+2H5hSJk0aNgmWdJWcbDWEVOS/8oWQ+zC2xMQNeNwB
1SC8mnI+eWvjGH1snvrMT4zTGx/WjceVgSnqhMBukmZBPOhqkunrPLRAPnaeRa84G3QZXmLwD3NW
5BMw/o2J6Aujs+bJCT2MBDIG1kFSv19/hmVfKsPfhG7VljJ7z9CLMo1q3Ki8SNNlEyISzvjAplfs
Qo4bXLf9icWEYC1QA3xCrGWhKLNF7keeq7GMDmE+8tdSjRfzWRKihzEiV8dTAuQYh5vn3YJ++iao
abucbCE9J7hv1FQcBCaO/yv3sDVgYNWECbLhbwZIPr58yUIcf7JOJ9WNEOWVbq9my62KJ/ALURy7
8dtcVdoIUU6/KuLYq36+FGnpGhWWFq/YcxXrGuUa9U5CMuqbDVD178QLeLsDvyT6fSJ6VG9Y0CCc
euIR21pF849B/Ntf91prTMevafCYyKnVEYdR3KCYWEag9gWBRfseVrIKHqJ7kODAfNFsj/isO5lg
6SRYwaTu6Ir7cf+vDogNyyhd7K8ywlnw6TMxBx0wiiniN7ETphEk9EonewWp5ihovc0c9D/xJhJF
zfB8to7cZHamtBbKDitAV3DAk8oIws0PSwpw1omZPsPKI9HVFe7ONiinjTRk+ckRkhyZb4irbK8L
WosLexO+u2FFw0n9oSC6UjXNQ9KVrO7X/0vcJMi6QVq95owMJ5T5L+a7zAcDPrdCJbyeUWu+yZG4
erZAZA5O2PgpZR9wH1L3JlZ8ojh3XHIqoAU9elT86h0f70pUrYA1CDgU5sw/ZBG7MEoi0B8twQJG
NgtDPMNI2Gp/gmzNtOtkcDnEKgJDNKYXCec67dOf8zZwnmClZaZcwXpwQNUYH6cR07w/z/2HWMtv
kSuPASY0Fbmuvu+jF1N9dG6tiI3EnIaMN1ZNpq1OV2UCm3/Ck++el2+4N6QAdv4sYzMEymXX5+T2
L+zIaPkU9r+ap9t0vMb5Ab/RwfLeXqYo64+KzVlK8lz7hAmGzPdXHwXpHecHY/toSF0k3YZWv7PG
H8VpgARf3CEUO0mLaaWA/LE4o5NCFdiSo+ucjFoiubAxWd+VRgphAfoTL6b9SvJovv8cmgqrl5Go
wgcogJrWV4a4/VDZaDM/RpyC10klUVE8ZTTfSzVK7Ytn9M/kiItq0WfyoIvLVW5LHflYGDe1ifuG
PJTu68usra8LwziWaIgCInAHTSeLCsp5LGNJtUeeLZ0a5pvznQsRjU5AAqUEGlU3L+wJ09/72ftr
yw4LGXwzPnMP9cjAog2+9Qu8SOp2WLh7g/o9E7GFpMBjeFHcB/jXzAjZGZuByYFqvjK4qIGfjgGq
El4Ognzj8OLNtm7/pq6ToXgZ0r9FmRA8eA6sY6yZtxCzTAL5izw4zdRrTupuK1XbZxaWB88UjGYj
N6/LrEFns4FA/ElyXj7tDWb5NbUsc+O6PPFx47kox1efxsKcogwbctwQx6E7ZxgDVjJRhy1G8+Zc
PEc3mpxWhA7n5E5zxxGEcV7Xo+VQkrOPrx8mHlJ/fj/Y0qBkwpkNqIiVIXJ3FLul+CPhdPMpzeVw
dqKfpNzRkMRAwEeXJPgFENGmeCi7cb7PSNhnfvQAmXi9ReKwiR+QfHAPMtOCU6aSvMaTTvhO8Gu8
A6hfQcqgzZntQTcJrx5m93zbqJ9qVV3eUcUW8bHFyekWOCZem1YrLQMlk3Y6oL4Uq9By037qJZTU
JaaMYVbQkMmHdycN3A8rc3QC9aSzdvjrueyXQnrDROvTEFoByLr82qVh25NDDthd+2mnEZ1WkFEh
W6AkrpK4m7dscawjBcz85vIfkkfE4cRg5ooqZWyiangZ7MHei/UjVPF5b9TEifc+gMOilcoX5GGp
uLmRQyHebzGXDc+MI7ofbErcmtITebjCHw75OlDf2n/sPZFe2NGLlMZ7uFNaf6U72T3hB5ZCIXtU
UXOyllsfyukivK8/6zhbJOV7BHngDW3gQW/UsDEiZHP1MX8i+x8ITMXVhsXyN6Gw2Nx+FLMrhz4a
b01A/BNti/h6MCi9R5oRJ2TF7zbApXqDTUnWNYQYGH2SXjeb2qVCmSKK4MmfqgcLzQruTpDDtggG
559KDTx2auq/ox4FGPWOf8wv4BmTGZJYJPpPVZd/DK9sVfTbrwuplNc1+hUuAks6D+Ew2oRGt+XC
c8PF1x4lsI8OeKUimckrk7OXlisRV+T898HcFgcKZBWHqk2ET0d1A/TiKY2c8/+0iaaEKFfOiAHo
zbL9mxVAW0QToFLsTd8/fF/TxvId4kvpl93W4nteshvzoSO6S7Ad3tZMBTfO88/i66L7tVzzqj5h
noU/3PIXN1ic/UwnnV/yl0qCtyPa2fzFigKRV+lTsBFy+KktPYswr2SZ76iL8tE8+M18xBwDnJ1/
rCl7MhHt++UmtWGK5PTT+d71rtqPaMh4pnL91C2Rt3B99zPqfZrKl3+cWwb9JiMILgSCKFZAhoH6
GvdixrAXHF1ikU8X2RkiildjAx0nUJGB0bHACgNnCdcxhZ7YgNSYBC6y23baoJZ8Gcuq7GfIqEQj
m1yzIT2eG749Nu2yePrm3WJbVNCWqYJRbiUY/WEziz7Em7tRZ2gukF+x7uSN714/IMwbl2CsJQYZ
67MXNHlUE+lFNxX+agSSv9XyP6jvJa93nLeFEJjrK5uLpd+ggVF88jfTrg/CbbKlAE6XcwkWlcnU
WbsYSeBOnh5TyZctNwLyNH5ZwYPtJlrnziKNOvJLpOTb4cWK+wGTlNou5Om2asggvuQa1HjOmauI
31pyxN2GyD+3Td1RxSh/VfwTNGfK9XwRX/l+pSic1ZvzNUVDp/vjF5crfiYqfWjbmqiD/Fn69xkz
TicWD0keQ9YTjTzoHMLFa4YLMGXDhWMKW60L4qLM2ikZsHdWtVGzZRXYV9Da84m/eksYkXqEiF6N
zX1kw1bPbcv/SS7O+tNLu9r02PeeWLJENPxlHFICOP4Hjn4gWUa0NGPBIs/lPqSZ+Xn3x4EAsCjz
3Ve8CR19+uxjNjMteqwZHM1PxGn10AW3Ui6IdVHAmu02V9feFu8/Ts88qBBnyfPd3ElJJeNZpJXR
r4clo9MSInJCp2RPiFjqj6HkxF+SNv1AGTEtiBZD1NkxSeWLYeb787e3eDZt+oi+J8G4T8CSCwwr
eOpzB5ZY2IJDo8vtvj9Y/xDWghxkjbuRPxRYYEalalBPFtfFPRCMZOaf6aKO8HysVOZ/s5pRsRT4
hva0xPveNtxd7Di06Xtg8mcEkD+hU0bV8h+nc6aUJvXA2em+0D8OReuzgWgJ7UmP1E18p0f3jTRV
tQH+fqWPGbcD9QvMvWcQ36wAElLHhOJ2yUrjaE/yP09R5+4gnVt7+bcsp6Twj60kUmgbCKsOipjA
NJQAXueK5v1HTuAmt8tfe8eSx7sHWRQcaQm+v89FhnN0IoghGFUsr0tXPvp9np4h2YPOqqHSj6FI
d8OYMWiy1wA8ayVZDaDXFOYwtslOYqSzgTS1QbEeCsQbMKEYSIlF14wc15Rf7zHo3lJWNikcnc8D
F/56bAczZRdK2zUnpyIu27m0VGDoQ7qMHl/ZCFY6IisNo5HyD/HIBYX/41tlODzZqRN7QHjZUGme
UwjwKJ9AUI6F+ntFJs9t/tiQbajgMWf5F7Ks12xrBLn1EINX6UkMAsyNJ/+pL6Ga0aXIbxbheJRF
d7iFbXcGE7m2vWccZDV8keIeQ1cNcpag10+kgPHHdOzI0oWQ22W5HKw/9Y53T7IE5W2GPU+3OR5Q
kzc58nUgXPsXXsSlTwel2upwRPV5KDjH1psuUtL5qs9+DeTc4pJRBN3dTK7gTn1gnm+IkDWt62s5
m7NLH9KFwysgKAtAmKPmnkMw7thA9tJRnd+V2+IQa+c8fEQ9Id4W86GQIsCoajfPYeVaPNDZIpri
bJufSH83gGbr8SNj0OKQiB0ovE9GBRQJhtBu5AGDBawNfDwUfZhjlgUV3gxhvBxP5wnfJKTe9po2
lvWc+K++nmflBc0VEl1lgw5p1a0CmDRCIe9ytgpMXe0GC7dnupn+lrBTfuB2SSmVZb3U3YwxjLpa
1j/SSC8pXtYTb/xDWHoRdEC9lvBzz5roN/QlTgdZJFP/JwJf0ao9IetaSfQq6y95NwAWhrpnA4ff
zcAR9yUMYgJq3iWzrmArsFG9eAXuHHRfArQPDrghrC7k+Z5Av9obk7Yb9Zkdnvp8QhSQ0/e8rr3d
jQfKnvehdujp9WS58WfEy1gAVp2TfUrShIqzraPxzaWEgXAKia3VgQeVf3NTb8oaZvdZJmCxvSd4
C+TN8CkDWgNso8zkzbpIWqcwiMnje0mvFopxHIZdNxmC4gLTqenymfGF1ZP00nNh6S8wpI/E+p64
TNB2mYB0tuzLk/zurfGMwNlRepB04Q0mNGWbxYrWpSyzLmVlVMnDRvPQb0DQD59yypOeT3Pup/o5
Q6Vn2waEYau4hHr6LqFVzBUdwrlEgxD/gjdiCyYJCOHfCHtO0RPmetdcfUiRdfysTDz25yA9EVno
QePAzY0Scbk78EeVSE3nE3SdKQULLJ6Dtq8YVZTmfGq/1C8SwgcG6yUGeW4k7UJ0o1Gq4aHC+kZi
rtUvC8ToBWm7aDMIYOZ9wIzKIAr4dmiLFC5/6xqXRmshxBbEp+W5OXPFbD6Xpx8NtyYCbQfXFY2J
p6e6m+WDIBnZ/hgi4SqUAu3QBug3SCfFrYVCdyzuZZbxpOV9qlacrFKVwPh8RH7BQDAmfRd2/SQP
Rl51OQerZC4CKGm8LY+fG3lOg6p5cOxByikf7Gdxnz7tGdL0SG0EPBXP0FveSOfxUcCPN5wpl1wn
E0AdQjsKSV9GO0kKM9MZO73YMu6sMvqSKR0V0osC7YrmwWQBL6Uzm+08TFa8JF25ejVPlMe+NUxn
tBAWut1bEP63rE/FrNevTB7gnPp9frnl0wSzuKzeLmLLP3Hym6yrikvxkV9XJru9M7GvWj+lCOBq
DLu4b3vLQlspW8gQMCp9aMd/TnOA4XvHvNZnO0fRQ7UHb3vci2coPP4ujy/zTXg+ccD5PFScXmuP
XpsSBmSoe3nR+pGyvb6unC9Tt66zKkmZdmRnREmkSKYgW8fd41qznux1JU4JJatcBRx0T8ZsQagS
DrWEUow/kb/Y55rKFDfgsFEk3F5fwDSXBnXY6fmNZ+1+QKuWSKJ9zn31uFltjS5JdavnOPMf/PP3
DQWPJXL3XyGKMbX5Z00P+HsJwTaAoHUVe7zWYmfjSQzpw7GiK6YGgUpgrEwdmF9n2iWViJxEc5j0
+VHVsmx12LMj7LSSZPtr9wa24DgajWe+Ds9dMTHJRyznKhYd8sVM0IWlMEpqeluKd3q8wkA8P470
0l5S/j/PPVqgc/uBtd03OB1Uu8gwx9+5I3D87nByhyIKTo3BniUv1kNqg6DXJqrldGg4Ot9DhoUR
XspBJdwVIEyN67Jd+f5kbRx0aVyw0fjZq1ru1jMxEywYudusJk5z+ISUmPBI0XHb9MJYz4rj7ipa
gGusdZbYWZFvugkyPGyPRHAzJ3nMuy9LV2S5B3bHpEvI8IqhYTPu9MMELo8qU5S1RQ/F9FAZhj/c
EWKu/5ABCLFCPCgJTo+CkLTZU2vzL7vt0AmOdr+b099u5P3wXGqzCOOQ/EIjT9OY2gYup2AvEGDJ
7faJLyIRHOkB8HlNSToGY/fVvaNYz+P2Uw0G/8Ub2umoBWst5GepHakGeCdMOGJq/yI7PkSmdSiv
XeSDEcSwHKU6cTIaMs755gINT2kVO5UYs1aExHGbI1MYMqb97kv0TkSPjy7vBDVgodBqOGwPx9mi
M1Fu3j/zE5q+8ZwNyiLpUCcsR2QyYsRnuTTq6QotJGQiRBgL+Wg/2jte/zSRHUW7AsVX5iY5bl2J
EiJKDNBNGGJ4jymwfxQUoNGxx8j3okwBmhTQ4TJ2TVo81sg+1wR9AmS5d7Kb1FpPGjRdRfSN3xn8
ANzAYOqFL0uYY+ydNKEIjCWoh9N5rkWXMIjChrp7c9wEA5xWnD+Lk242wgVsfnQ3kI/WFs8DZwAA
D5z6e5im78V36l4ww5MDfH34ljKT0CLLOnqezI9a45rLRxLE3i4h+y4Zkqd2RPtNE6ZRLhfBk7Qv
vRKR3KT6mRHMREOQ21+xx6Zh5wXd578rWn97QoT1AqI1VO1j+iimFVxD4iz5rObNDUrjeIZwitbf
U+LGcPuKNcgT953ahdF7a2xWvFRisZ+rClM+5DHA+RNZMtRwrBSNDV/bFnG9fSGPoOW1O+dT1wXR
3t0cqPffUZIgkSfSz/MRTbP24PStLQES1tLskQJM0IY6rmOS/Dd6KooMb2xo0DfcBOCbIFeU1coL
dr0HRcBDC8puYFVlB7eDShsHFc5J0q+U1BktDG//axcGb9JOQPzOayAPRsCdWWonZc6rti/V6Sdv
tEdQlA5xrXbu7fyZLv535kcgHdC6Xxo7NVBbeNs+VcqXbpQ9LflWxF81Gsu32SoUQPl9ZdI8g0aO
XzU/Zk7WKX4EEtJ5V2xf7/JHWdkwlkRL+nPh8luGdK/1y/vASPhl6E/he+hBfU56JGsecsw+7tv/
JHDurWqYbzeM/M05QM89AK7CYLd+h3KHYlotD8Gu4mHoGvrpWOVbHGjLqPU+cZ8UkOOPkEmGeaMi
6lD+nJR1vzVKLwpD55MBDazPraOokuodWqXZS6Cpk6c2hELkxe+SnHd+iLSRKEKJMNUWqzkmRbaV
erVT5wZ7UQLf2MqsmVcQTypuS+y56+iJqQH8DV6sY5bMcFfL4b/LunptUunI2cK7yOVV1mqaDZWi
jlHlrUss0Cu3JNbHZcpfqqv9fyk9d7o+T2fHpW5x8Wo21QROJJAzkogS70bqLytoYWtEiZBzHSJU
LLeEonEpJEpbdDDNxPM7Fb3NnC+bwSDoLXchhKD02fdGx3Rr4AYiEOeNlY5kpUZoRg0uGv1tvGrl
nyhzO5+qSr5BCrU+PqXci8qpZHqDTNvobqc70TliE8uBP72873I6qw+tKPNVyo2jAO1165eY8+N1
BabikTgUVUsM9D12FlUhWV1hrrKMSSLC1Z/gspRxjCCT6r2Ew6L4r96hhwcTm9PNtxeb82IuwHN0
EOPGaBRzzn7N+AQDDU21h8+cQU+kRLvSWzBBioCm84iFJoxGtFxT1ePm9W2pXWgk+4Y1nsoQZGyQ
2ogB3P0inRWCNB4PNZNwl8KDJM63EIkszu8JKY3YaJiOrWNFfmZvE6Y3o0rmyv2U5h8U+awWZEeW
iBYRk35S3Tx6XhVE6cs6HDonDXt20JvnXD9UOHl+kkfsd5JPDmg/EZ1SA/95/TkyRmvfJ0NoMt9r
lSvpVpi4TC4bfpFFfU0Bwp7T1QUWAJgYkv/nj1Q6xGkfXV7WDLSHLWvNLBelgKju7Qqh281mwnU0
TvW/SKKGEBrXy00KunFSy/aGQDbcxo0CWUz4RisLfcurR4SI6md4ejn5n4mkmiY1RK8vLTtZr/4D
LmpFqedfgVM6k4fiAWMFMomMl0zkbsqvXIyFe0vaDUH63EHpra7DGO2hs7t7wkJgnrsV1RXhVm46
gUCzco0/CjLpA/dp2OAgadH1XD3mooFUuoLbBuTOlhO8Q6b6CWzqsuehv9jwIxO11pqdigwmxNno
sNwJs0Ejx7Ih2IJaz5HXShGFUAcurHhDb08iRS3pHUjcDCD5RO/GtmRG5NYn5/M0naOjmFa50F5k
fyl62CTGlZt8lTkIsrpYESYvrOC5oyTHjp+lEzRZLV9MF36yU8qhkCMRGEY8I8vDEs72XJO53fk7
KV6SwdYZaeIG13ojolMqiwotkL+RSL5Hm8X/tPm8RHD96M2hReVQ882djLOnxsvV3GgvfnGTkoSw
IVQ9CjcY52KN7HbqQ67QLFBbZi8fUfgVyUhOaSlCBWtSJShv70Y0H4/TWpgpbbJddjGGsObwVc1g
bhhGOmTbtDQyPA2nCIXceqyaI7PQ80e5gX5GICYAFQkwlCGx3dUZ+cXQ2R3rkpIAw0F8rBHRMoVm
BLZ2sDWrAwkApE1exUCN7oRHPYw007xdQHfvtr32XM1eeZY014gOJy+rFP7SmpRoI1nqsaeBvJnt
8JK6zsTM887Q8/GvqCRnxV4wgMVdPzoD/QL/B75V/XeqIP4GCL7DGYRkEnln8ZIj+QQgiHimNJPg
s74fQrUoyDKbSbfksjM3dNOOCLqFLtYaZXbjJPPsLPLp69pFkph5RUwtjGbBEJQfasm8Tg75a1Hs
3h9OSXsJ8wbo9m7deAQ+fVmd1zSfv12O283CSUrWPSADjEU5OIjFS7kYFeyRq6ZUzg/gYtsxIbjS
Cv04nZ0QQ5fVf2znTEBwKg9D9ahDSxOKROUL9S/PrIIzhUgrQHNZEbvayHffOkHA2irdPkapC5Zg
zj/c6tDNB7qNz+O3w7mDJwTKP1H12Li+PJ+1mNFYdQ/M43rOw67cDbJ99/TVqUb8WDKU31RsLSJl
FIoHvkC21OEOxWV8KUSMiEaIkPXRNrwmqA8q0fOOB+/MqLAh9b04XjMesNm7BAUJkrr+dpTXiLWA
BHtL0y1PbUg5oIWobJ074THlZJLN/fM8Kt4prnH09BDlxzDFW3CyWkuirvytR0HuUZlWwlkaqFeu
x8NV2KaXE/97V3QnScl2NbqRA+AX59tAFznRgEkXMeHNoUQJEJ0R/MPihgWraD3lsH3ar40LtC3F
2BhA254hQ0qP2lNyHvyHxKvJ3K2PE3D/ScJgQCMqerN5nc5R6uwqqusGLO80/CX1llAO/DqVrr8v
xyvJquLnj+wxRIImSbet5+UOktw8ifn0m0Uf7O42K7vootr5e9S7ulJERmANexlGbVSWnvqsmro1
QHQ/nOIa12ihRCnzy8E0i2gKX2As8SxoCM+UPu9UNzvurh99Ai22rueRwNhPutulMLrqSLEbhHQK
Jk657iMHrRAHoYPrrzMUR58+em6sxuGWQS2dNx978K9jyOEljiDPCTLsNkPvytVQGnwPbrHBt0XX
orOJb6X1yo5DYWl4D5fA+3PrbGoogTqB42KAyHHX8IXQ1Jr+TkQLMGGKuWLkpmA0NUUph0njL4e6
T7GpaS5EI6bC5A9g8e0l56LAQpY+6PT66BaJwdTgEHIZ9LvUN37FUOz069mkntHHbN3xNdfskrVY
CPWsEKbKxTMhxnco9bZaXtBE4LJNZk+aOfPGcV7ZNByoyvj4zgMRchzrrlOmb6vgUX39wtiCGk7F
yD4xrxoa/PWIx/dv8Sg04JdD1h2AWgojfUuLp1fPssPz1APvCo7nypQ8Wlbron1dEVJtMN3AYke2
JEbQ2T4aUZwlMlhPFNthr1jA9GDT35CvaZnQVYOLCTEjRyy0PIi5CzBA37Q9SLlCp+GCKfMefhA2
thMTyMS73tiD6PbMS37yM8xhvNceaBND3xUTyZhxYEWDaAxx1ndniXvuWX3M+dg1iFnZ+4jZrMax
hpb68HE1/l0rW/EKUYMsz2uI0a5ww+wBaiMrIVw0CxR3FSo7FVsVb+bY0Im6UP7doY8V9oGt8J9e
Z2225y33dIZIx3eZA5Y45OFTDbVeZAX82TfIBAjXLCkI42M5X+U7VwelwzMiUDN9z5hy2ZWKAQeu
3saXiICoCRL34DyO0IwysLHVn3yboZG2011/U3Al/F+7O+dc9POQ2KcO7hcafUHFquldzwsZFIAs
/Y7jo7xELFfbxW8Kxk2c/sP3vPjG7z3XqYnTRD5rrjY2AqjMJJoniWoRwxJDr1t/1RiRNeP3AN0Q
DZByhP4AN7APqsB5Z4Rs+xQtL66hPqvIt7BxHNijv7ALj5pShMF5NPBL0xH5TFvJ/yAB1pmnZE++
i7PySAmOBKk4Bmopm9bwIAq3zymXGYKnSywNdXaMTUTqoPvy9N0Ff8IZ/FCc7dnLHAxGk7ARAoRp
eadPix2NH32e5bfC4VQXPZb6815i2uFmM7UVwPilPgd9tHH3TqO+VeQnYotV+jmdEb2sN98Ex1nj
M9y8UqD9JIe/A1/+eEkcGHDCKuZm87kHh3IA6I1W1sDaUnUM8Aygf/ORFHte1/mQuuBH85oE8nWQ
foGmAcjXbS0IhdPDGm+HLA8Iit+BsyRyfJXFvDgQ/v2n7nK7UXgBjje9bDmpa7CDO/e/+A4/D1qp
52Pyo+uIADNxWu/LCyxz+ok+lFE6L79T0a+wYqBSYcWll3z7DKchVNlGx7GiHfVDkRZEnNPoBbWz
jpoEilsrUkKgGkjPkA6shSKphGRwtholcrmAUecbbzmSI0sKo4kLXLPKl/Gw11I7VbjntZFxWhM8
0ALBqO9wQHNbmRhAPCUtDjOaNSKcFIsWtXBrdJxLSvpAosZPgXHmYxlRqYqHwpFXFB0ykQxnM0wp
XwhfTPMMbgPASUvaEL+YLUn60SB1Z0zxrPlZcwLRBC1dpzzGzcjwPcwtVMeeYWz9+7/dmF86lH+Q
5Yd2SYeDkxyP/01Y3Vj7HtqTFZyu6koWxqhSqAE33r+x9fi71c3JopWtCWQJhGQTiNrQK7KZptR9
HTZuH/58GdqeMuYja80YvRBb+dGJCmeLFLZOVvzwjmfdINWvRFFDxOTm/v3SqvBQCCnlGut3HxKW
+XEyMhiZI/BaoX4uYSrAcarVgmGa8ITkxapbGv4uAOdFihMg+RPfT5jCun0mbxRSvXgbEi7V4hDx
vYi1b5YIa25tEpZqtWg0vo63UV0yfA//sz2CdW8Pv5hy2/U3JMr6wX2xWHj8Zx59YtYMXus+xasB
hjXKGMH4J7QF1FeIA0L31/sj7DkJYudW0TLAxN1IXRXxI1wyt7Lg31GQQiI1gacHVHbIZff5Dnf3
IdECNMvUuAxjuH8fzidfJCcWvzSJtfSkeFtuqZ4XqFvYQ89AISrHh2Y8P543oQnVdS1M4dTmW2PR
Yg/1k6k/qxwjurQCrFYZP68cb0N/HkzGHmlkgxCR9+X+O8JO9ZzFOzdeSWESkIH3z2EufiOYyzJg
7/K3Z2GywMI5UTRb/4JN0rv2WiJLJ633TrRffISeoP5x6QPVLVuHRyAspNjcnquNznkoZNQ1VcXW
6SI/k+vwCNmmpzvOGKktScAySUb/717oesJ2z4wemYQEYIM3IepZC2jzX4fyPk27cGwoSfVOql7i
5SPiWwZSGcu15VnMJ4ut1o+zRpZjUtcQ2zmFXNnUKkX8Hv5Hj/asAzZYlOjmTW3uF5vN0gR+QWPm
OJf203plqt1h2nmSiGT3CfDwXDb12UxF+St34o0XZi35WZ6m1Uk0WavY9IP/3IDiSJrf0g8ZJQm9
W5aSCdT/EylU3CkmrXlYZYpmhH/vEHnE3VeCzkf994+/570fTjfuTDj/D14/Ly3H51g19T/1Iz4K
IyCuCEruTclpPz/LG2Y2
`pragma protect end_protected
