/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 848)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B6w6teBKHMgmb4jFN2NC86rxpXTAOh23JhHEbmjZNkYNB6HFSpeATRIOt
QPmNY/bzjomS2qD5CUWuq+cvhM/i3oaevy3DnMoLjAj4FeB9iPw8RPuqUDnWPb1IBN/e7qWDLQE6
sFTe6SZuW7juX/ZgcehS8lseKO5T4hNt5NtU/Km4lHQo0C5WaUp6z/woM5/nXB9DCAXAMbbBgtpN
KMi+ENUA01TpgDB+JsrdSLbWO27X0wn6kfef6LWeDWEZRSeTlVNSXSWS1Pm1+xb1Z8oWHn550SCN
mCxXnhm4WNv+uCvbB+DIkR9sNKw4UEe2lazWP1owoKEShFxhawN7hF0vEdjh3wDM5WCuYtL3ZO+y
Df2K0LLyokuX8QTKbfiDHQttWmucyaZRVGRCwKiyy71R2G2Smqxalu/wl6kENEWzbq0qjFkUrEt+
if+w5A/1MOfblAjQXw89+3qZp9qDCbb6dbzuf5X+3QAOVn+03R6aqyEQbSGvZ53GJmNpTrZXzX8D
I3hi0nEobEf16+4CnxUf0VZXEBM47cHzd+A9hr4eiZDtE0VkgC7qjOfHxdyoNn9xaHcaIbwOtpV+
958KgX4BUbVZHC1fjD110CQ72TGKp9BuNHU9pg4sw9ep488+BxVAaXc89QAlM8avKQJ5cAg3fio2
OG5kKRG1V501p3bafsSIJS9dVkyrE5u0S2YoEENMtjTntAIKZhFwj+XXRlo69xX/1VCd+04GHpq6
fBQHlVJTh4xkXMH7f3CJkllTwcn2YJtc8jd5OCZrXJ/6oVpfrWIknsBGtq1FH/bdsUSNfbIjn8aw
viJYCQdONvAAho8rgD/gyFkZjFjlTWrYRIh1NNdwd/YJH6xLaWZnS81BwWiJ95kt1c+m/Uvr7k5A
8aHbC6hPTKSnagxun0vKNi5EAtEvnWU2Ao92aXnMec6zdQGqC9MXmkwHjpSppH17Q8A1wVT1XjLJ
5VrBOBIXjL3/53OuQs/GZ0d2WZtHbMmZwGv8Qx6tDukZPeE7joxPvrUN6Gb3s9j43g//erinVUOm
pqyoiIRuCHZpBgZrd0PVUyeui7t30B9PJFNCHBLbE3vj5cyMIkSvNUAq9wop/8ALw70=
`pragma protect end_protected

// 
