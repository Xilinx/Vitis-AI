/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1102992)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbIVl7Qr5jP+nOJ63FcVColVe2Lik7uB76ZDHEtnM5YW2JeKxRHR0ub5J
0VoI2UWFFvQ8LpwvMT5rZMUMa8fFJscxH48gcPutOatrMnMKsKi4ed8Y0Vc4HgQG0gdrgYgOLPdo
k8FJfB6qzIyQLcdPHpE96g2nSZ8TQJKGZoJf75J1ODfD//138OV1uRFmhu1x+xRH3sUEde6Jrmix
u7I0VxUkgw2Al56hSD12PNVBt46/SNq1EUsc2L0mQxAgrE+FC1zvbNdLBLT2Hiu42V+KWlupBVxU
2+LR1vKflE4EOwJcjPq4/5Yr6Y4RGx1mk9TfWOqPdIlkTTFJ3RppB5Fi8lKxopcLzPRfXkzl5FwC
ME6Z4YM/JYYVNyrG/qtUBEY2OHTzULGKyq5g20/qP4aepnSQ4IQGhqDwOsiSrQdeN/USx2WaIkvL
m1FIz/eE9MLJmC+L/Q1jP129CZ1XD3J4PwiYJXpcmqDprw/g/X8IfH2GNFTSqklz6FtNzU7uplH7
28eUGUBXiGcw5lRX23pdSUvDFl3sEHFC4xWgX7x566rFUTSqPCvDmRiP1pYBVAKmGp2FusW1qKl6
1ind4w0PpS0CASIJfhFFQ1yUHv6FKF9M98pEd9zimxKFDHMeRDRY8ee76Kmuw8DgY7YJ8c4DpQ8b
yx+DUSHajes8FzXQGCRi4K2P23Y/EDSxiJ9TAob7k8MUw94KM4nE2YiZaPswqkjJ89wRcg9Mmzcz
WF4tg7z6XryKCw5NLP2eYQFQyJYU6eAHjbw/FMJkT+GbWxp818JeVv+fUu8SHJ23piGsar95EgYq
aOcsp+CraqkT8ObrMcZ9wWdOv6dP6RZUj0rN3LCFfR/bwb30N00pGHRDbLa3sIbjfSXMtdwYSLjj
cina1fBwdVgwCIA9W5pMXFGIkuCPPDQ2AWJNR149Aykh+jTzPvkRyZIH2IYn1vWY8Z9IJDosLH1H
uiVgO29Ek701zFx3rJS6rFUsPRYE4TvMIFIuKh+qwRcTFGx8dFGseEIZWrfF4/XouDzmhbQazFUc
K3GPiI4plL9APXtOUQN9J/ItPK1RWwC6QUa2H0u4OwHduFc8cXMsIE5Srfac3D74LDmL7vY6S3PZ
9six6dr14qGgtyfQRn+/qEpj6dzjlVq8KrtaFL9jsrMi+6H7vsIZkB7645q7DMKIuoYeqHatl0rp
mogUF+QPTfO+SLi+QW8P8VO5gXjPxHSzTnLpmdSXHD52BcRmDFXPS/nTwceZg28m2zUDwu/z05lO
Bxj1n94YHlSjcnvLeOksNmc4PsspUxfiB1NNwnDQm5AZrxohoI9XGoaVtKMW5fG0aYBvtw6hxQED
IyDLDnM7flwvDgsdhtqdPHP34iZqmDnvF1F8VKCtMFprhIUZZMUd23ODK4DcLz8fDJRHCc1VQ3/P
ZihfzNz9l6cyI/axRaDhouH+3m1M+FAKufVgUGtZ8ykCtWy1T2s1Okc6pcljn5emGVaMcDGdQMy/
sdTfw1a1RQXVlxIsXA9GOCGvmp5aVfE7fIazx8Xh2gEBIKI2200FSew3r81sAGykqlk1hJQOz8Zx
7BBWimKGwH3dbQgrPCIAQ4RuIOWvGCY5SiWJYK9aNvNiIm1oiyTLJU7jNjJPSUgAgSUJU4wUyHfe
ZwmqRF9xaljIX9AyM5B1QvIoavLJUfAlAF+sG+4MiowwiUtorWI+bxv1VgX683WYsAa4Q86SMIx+
KQ8ZAMbmGrzJ6pjJ7kCGy56zQAKlhGD5Sfvd5C5WNrjDKVJ8XOqeXLDmJjTP0RaSNXebGPbSTjqX
37YeI+uFHkcG8K+TC59hCvArsuxQBzohm6j7XB2pd0hTbepicpS5AkBfSE8nN6IbM6OUD+MQJyUY
wx9Hpy3gJZza0NwtJIKmBwWiXdo4uH9MHiTPH/xDHe/DlfLh7ecZAwmslsia4+qWZgxyIKWhaDmN
OSYDvC50DcESvI4G5iDLUDaCj70dwCksE/aHejEE50qLa5DL5d7xjP57cSvggZtyM8VPFjtkFV94
1Vf0PBdANyuerxOJQgvh6itkkrUh+8GFukRfa3QrtnVpGjpL/x1Wtl3X5aT+gr0zf4F6mlCuWuEw
DBO6m4lvBrGm+2R6KsthpZx1XrROg7KH4aePrQSOZnjpuk73ZRngNkRfdSBajnlUXTmhWSVgEFNG
7ogeJF7rvFx4LyAbZYI/xKvjwuydK7X6qLz8n0KJCFSruncUFp+6p+QNh+ypwha7kQbhRmnNC59f
CebYNkRY1XvLOFHgChKWbfDkwe3h75yUTlJ1SMnc2LLnSWPZMJgiOhJrdafw60qFOEjdVazOgvRX
60vhvZvZ07Fwu48YSGpNoUsja0QLgCV/inOyh/dRhMALJTiXQ12m1hFHMEMuawrq2Zp6BL/tia7L
eP4LiNjmHlqwcvseyNA4hC1KzLfpmHWCOTe+JoO+9/WsuW/sYwXv5cfZPyAhm43CK80MPV/GJ7PR
+RJcCSxyjbs+iTgYeeoys848pQZFU6PlAFRm/bWl0Jovx4+GgUWhCp6zidthOJo96BKtBcd8X1DP
0E9snSPL3Qxtdp/9vE/FjmE3TD9LT95UrQ++pS7t6IiOQPtl7eRffijij1C5Y4grFwpb6+NyG10L
hlKlFVoTp6qse47rlf3fh4bN5B0JG7/FdXw86EcLpmv/hHWZ20/qJ+VdbjHmKo0935cZhKp5T/Es
4og3XATp6ZMBleY/G5/isW4za7Be1QYbQm1kCCsLN7XMNCoFAEo5+kZT38BTr0AiXEvViIMkdi1R
VyqL6svdbCbzdP90kVphTffPSjDk0FgV68D0gUA09LE1nE5miDsSNVlVR38TFHgIdb4PuzZspI3O
avFcpIy/HZ6UGKVCFe692SPiY51BKTKLUOrpaJhBlqEIhm3/qC7KHyeaOyGGw/v6ChD9KiFAmX7I
GBRfol7EqOHfHFqkS7zk5KrxyiPM783g0eaoY5ippGzMpbkX39N2h8d/aXypJfsU9gBffaYTWkPr
DmC/E0gBgwbFi0VeMY3dDguSH44fSziwVT7r7GS1GSdYVxUjCW/T7c0Mxp/D0+3pUS8arxAiFXA4
KL+/2V1FdwC3VGJB6N4gcJNHVqQ8W0FvmyUioFnX/tfSq46og/TpCJEiiy2TInVGZToAHcVJzakC
4xHYbsdsWDkDJQthdKcyGeJPqERAi8DmrEcotWC3KJ6iNDijPeCcTHmXmKZ+a7ltdE4zjprfNIWR
xQrtsJFKSKk0YLC0CRjqBtRM6QucIpV1b0LDHTBMotwe2G9/jzcR25wldxrgulBseJqio0CO+7fM
7xfqIuWCw+XAe4O8V6N30V6vWCAHrbO9TDx+2A3aw4mKFZxUrbulS/L83xu3OLKwKb5zaNEYkfsY
4T7UW8etnWJZgW+8nyVTI2mEwhQg/lB0wDv4cvuURQbYIqSKBKpxDcgjCDQLei6FzEIfZNTmu0Ts
SgeqYTTJXShBfwKGZux+aJ12BukazwPASmpmqMWJQxjI/F8RtRtgwbJGm8Gv91Bil73RRl2L4k5E
aJu4QdLtuLcOcktqCl4wepH3rpGtwsW81ctP9Fw/4E+RV+1MopPGHgaZtaHxAZEhvn+gQ2SUTXGC
3+YMpEPHLS6WZre/4J+J1RnhCajWs612OlYyUhxCB/aXfEgxvpMZ0csY/lMhsZd25Wk5UX+Uy9jt
hKSLddFvBUOSUOlJfoH9RDqweMlgW9ufPJljAWCHWuAoSB2RJdEZdhUDTJm37KqXdmWouYHPTtU8
7PbnVkx9acjYrcx2BeNETTuwbjtY2nw0eitx+WMizm+olV/PdcQKvAo0IPDvfh69OZ4raNNF2dSJ
iITUrrh9bg+pPFLjmtL7GvYSfgWg+wF0OXFwKh2edpPUru0D7Pg5gXV+dfWKBNXi14xFYzesdECA
MbMWw3mf5Hom95JoG75n4tZhOSlW1TsnXr1TXXXiXyX4lZ/gt1/SO6RKoA4QZ+rDoupwU56rd5JU
eO82/64YlgdheZ6fJFJzBGL1mexpsXFQv9TSyyPe72NzOSdtit+CJ0qn27JrHGZqcvkB4Q4imszC
wV9UVlDhNnMo7PBNSRAfQPIJEDIOKjUkG4siSJTQIQVkv9wYc8jZh0iTFe0A3uMZOgkrpHFNznX1
dL7Je9mKHZDD1jKbRlMnO2kGV1Fl3XrPbq3oaTXo/E29g+xleyp1L/muCvCK8qvI/j6Tire9JXpk
vMKW2JCXkdsnA6HVyORToeW1r+YiSVsFclOfjNSbiUbUDM3FspEwGrir/HVPe0IHHuV2w27C3s7n
7En8TPhqCg8Dnpd5hcpd8sstCIIU3ebhHMR2tzu7oihU9cE3LaWm5LlofnYsDFZVpiETD09UavLi
jdYu1Nja633Jm/YTAtKZhJr3ycI5q4USG8yAUekPoDWj/qfGzK0nV8znkcWsHHUPuNGLhXVznfYy
EEOeX+yXOHdIkUIf+V12p/nOiQIg4pHYtS1HRsGn6EF96yWXcgSXbwCpScweJKWtm3v7hVyCvmeC
u8c7Cwiz6p1L69POqMmu9mFKzu7v2Qbx3V1LJQlMEa9QoJlI9YeVOdjQR95xxZdj7ZGfjlwhvPiS
eC0ELguxuPrTNzBrf3EGhMpMPy6FwLnwEMVO+LSX+zOgQPEAjaklacSt6HBF7CdjEujNHoKMarms
P22qXgvbye7V2qdAcKHrJcdyd2VbXibTjVu+iWjKiF8IsGr2EEQf26gBSvxhf9okeYmjb5xv/4A4
xNu2Wj1ryQF0oa2ZgI9dtuKt55CyqXmP236aERYyolo+olx9MqYYYDKJLFQzX5GzBqtJgMDbTFOs
ucthp2O+XbS/W2H/RF1WjHClCaqUzzWtqUZ/VoswI4PvCKNPT2EjGv7QxXjWsIEFi4a3YfPAE/9E
yBWOnWl6nyUk3qro+v+yHWsaCEzVxeFrJm4X0U/KebBO8YrKMtlZkWVmbgENXhDGfbv9NjCPsjdr
L0530bOE3Vg8OQnQA5TZALg91R09QyNyo5ACpgqa1Gj5afwG62Khm0SyiBuWa/HQC2hgr9FXN8XN
xs2QwofQ8cuVsM0d10m8oS4TqyLw1nGMFYyKbTC5AG4nf2f9bCZb0dGA67BQP2tfMTUTUGzutX+B
5s7LAUJYOGvD/fI4IJsxBmqOqvDWnycHqdoHsFq9/HWWjEKqcVEtDFCYmnp1j1CzJoisbnGzfXc2
DU7ndIhvjG/61gzhNVPTubkr/lARdpHFTHf3M9xSB2iYBrKogVdXNFVjdwGllazdkg4/Q6ID2xPw
zhnrSRaSsgltd1shTxAuuSfNmcZ+jpoYSX8aBowNo9wljOsx2mmFJ5LJ4IRETKY6fLkaL908F5XL
GA0bh21N8byxnM+gbR8ED4c94wEaiIePBW2Z9rGlQYSiduvH8GORIml0NLJXljWP55b5xWZ47ghu
qAKuOv2oIJ8aL/4d2T9p80dbmCEBkAlB4uDxK0gmAfJ16q3hd/52iGdRYu21fx+a2tglCFMqb9Tt
lKzDPJ7ibsiHW+ycmG5c/Vz4kIVV54Smes/l1moOc5l0J7ZkXgBoQfthVXRQ/ovd4Hvs4AkRZSRA
yKtZF3D1EIS7yV1LPHBnZD43D9Ti5raMLU27kPg0wiV+B1MHD70zi7wyp0wYo3p9ECWYYeOrrpkV
9u6eGsTUWdq5PtkMmnDanhGHr7x0dm1SClyZgBMr7h8kixDQo6U80M67Mk6qufmJFxBO4TjAMep6
+ShknJBw0uumRIZcksPmzeMdi7wHZhF/s+yjMka3+1IlniZerF6s7pvWD1q47pvkH49BpHbPjan1
ZM58PSoFU97EbBE7w6hV52ydZhEFueuV2/QfhXv1q93/7teIJX8hiW3RtiTzxz2NOSDLsxxvw2MC
z/7Q+eHHQ+EAeOCbfNlb5bpGDAV3d5im4NIdlYaxzavhyXRyiKWXK5tBEruEZdotsUqB0fE+EyR4
UZFPcSkxZtJGzUQIHH/t0MoLZKNdsqyrJfhCEcFJ8DbgJE8DxLFpnf2+lAC2PdpTDraiuCftKIZH
/UalkGo+X/ISQ6y1fDfVrqqAh+msvOTqxsAziQ8LOd0XwLgcd7ZrDyv79/+PNCldqv+IpFpEBi+c
HGMBUKGQRl1Sz4sZlEIGmscLylcNR7cjywoBCA9dFjOVvo1W9sh5VCWUev5YCEMFGbjM8qiLV7rY
yZce43ngGfuIcib9AgDWPvV9y1uLL0FZaoRAIqSlJlxF2XdPZF7HdInEmqnQoFZgTgJfRhoVrDSO
Mn99zguKkbAks7mT0qBK4cavBQjBp/8tcyzyFImZnuSQM6tDZTH3ALdIWOdZ3cY4UaBtBnQtXKh9
EEXtX3WYSofSen06QWu82vaBbp5cTjNcPiVA1SctyW5INIke25Er8hMGxuS9NxDeOqG5vxY/Smfk
jfUbkrzmoigPkQoal5olm3OXLrLmfIaWFawmzeUqPfBLGYw2vvaUslKytBsZ1VVrllc8ThZVnUcU
gXu/3TXpggI6ngtkP2QLjKAeo5Oi6ByCwnY/uQ9fS+npsdlGHXnsNuEU+aFWgHu63FtiZ/2pR78S
xlVkzHmcHWSXM+zfwpnwx14f3icSEfMvI879ZieLD5UMluKwDBIFHUbagh1SSul8jYLXN3r5FbUA
RzwpnYP7XM8raKh/MlDxmi0hlA25Zab9UOlhDWxx425mmzIqlr+p3+jLH7E1136euajS4v1UI3jM
kc5NtSrclB9tBYXLhHefJymfqC+1+GE/uybRSyt6NBiShWtLPUxP6UsQzy/wr2O51wnD1krcCyxW
qic/6itud0WgobvDfouHAcGHyXxBrLwZNjGvDwJtEPwOBCV7J1EAgErNwTnp3x5Ra1O5GyGI6KWf
XTZ9tZdre5LZ3HOb529xq6rsn/aJeRojZxmWxoqXcudhzwV4aFyeIyXRdWjqP1iLPxJFGaPCBzWV
InrHETCuCyu0rHCWyZ7FcawWey2ArkPzaGQUtaGu0642myy2XWV6j4q5uuQy063wxeWKjtz7wVY9
eEZCqcFCndVfFDvTCr981o9V1RbM4Lpr1vVsfCaPs0hveS4q5cepV+aeBLVneBYIuk0O02RyRMk0
m1B3BpKrWAqjhdaIl02HqyDpqmgtlZ56Fzx3/U2xgV5BTMa7wNZXbmBXbuL/MXXkVrcmA9Pmil6s
N322zVIuX7HbJ/odTOjXMhc6qMITgAkAZWVkn3dylCw/Qabdzivh5ip8PU8DnD1HvDN29XxG+R6i
DLmwfVvC2KVDclzfsMbSBMsohk5Kvlin4gOFBPga4+aSH1rlE6bMLxMNooa/s+efuHA3siqNWgGw
WM+DEEWiE9ykKbjN8kcf/4K/4+DMEWWNpl9FN3AzN7p6PeU6lGnFpbqxi4HQhEGCHTQWuxrBJ+Jr
mKFYpKY0nKC5XZD9rBy0b5oc24HzsyC80R6FrBctLgYGsUSbSbE92Zhj3k8Uw5dbb4RcyUgdnGLr
to1H3ABDTq9teIX2CReLe9jYgQlNh8tV9S6lJajUmJ8DFVgeFUa+o4fpAczazxrhIzmTE72VCZqM
f0J8LuGvlHWYiXzziv3K45oZNdKTNTZidAskdu1bG99iFn8kSbmY80y4478BQwMViaNeyPGY72C2
EXI+tprJ4zHutW71dbXF5oQcJlwM8/w2Rg0Howdwsu7sP459whbWdtnwk2fW8eeXyHU1NAw7Ny5i
sGyeFvIONXMVWIJWnsaKtU3Gb6N7VuTMIo9bp6yuq9qiqHqawddZtA8YCvLSbcEE4xx5PWQ8Qv1n
VKIH1xCK20G2bLA92i4mfZvgtw04I4ngETgkalvYE+n6LKvec0zBLEpLUwA/16eSLdD8mYm+G8zS
imx/f2ncYQRPvpL94ddwXfLt6u+ShGr7NtskpEKGPMugF1CRAr/haKW1EQLzYowhaQOgw87iqqv0
oTV38T5KAgd7TvSiP9aWFyKOX/An0K3/4nsXFPyqmiQ136BRmwQ4E0ozinowd0/hVM5m2jpxmnpd
kLyu/9V52peko2P9w20PuR+u181Du1DFctUp79lym4WqtTolqsWmwVm3kOfvFHYHpCW3CmlC36Cd
c0baW3kUGwC8rpn1jJPnDILoK8w5vE46xQtgciZiOaA0twT9KbMPTW8ZAd59CVczzoJJo8XBRusi
cLWZxjT33sSHU7/9vIsmD0BYOZYnyLApbQXTzWT7KF1aulpr60RQ+LpB+EEt57wOqyQ4velzB0lm
GaS7mWwAy0HhsYYMZ8Nh3GBZsjHuLF8ykdzUHdCRNMfl9dw/pCDugxkfkiHFntjdfHjdFg3mUqhS
VuSCN0o0G9t3zNRmSa/uCYDL08J3SE1ycRZ+8z82WvTyPLrdjsXD063Y97BO+xMgjZlc08Gbr0G1
+K7RJnYXu5nUQQYFDslqEjdaWoEERmc2lafX03rKI+ZFvcA9oYdY7859XuZ4vcxE5+YMHT8/E+TI
wBYT0hkZ2SNceCY2hmF3dE2CJ4E5JdUm+ZgBD8G7BHLQZnq23vwRjAYbDG+OrvBjH8XyojRtf+4Q
MMgaDVnkxqp8SM3mNAN/06VVsnnWwrdB0MHedxKRpAvg+MtZQIwcubjOs6DElEHhe1k2hEdwyc24
ec16ft7mzJFJZiZb61A1jDqvAZwD78S2tcfjmK/Lun8mQDHSExeIdKotOiu+fScpHkIiNVW8Ug+W
tC7nYAt2yUzuwSpUsac2iFOM+BP0qTxRO96VHJDHJQHDP/YTL9StOW52HTlRAq+IGhXfMiP/AMXM
yfHOXf1Q/dWNiLKa1cTJE2bJKWnzwwW1nN8nItuZPNhU6eODIG/k3jc7ja0FeJdu38zfVaLEyPDG
0dYQIeNOEuTadullayVR/1vKWCHG5kmGH/CsU9qi2LaIJwsQ57kUP3NyZZRO+WzenAZEQZvfoapQ
nucxfJz76wDATV9Xm0hlfSBmTNLtNxBzZKqbfTTI6FH/gnWjXjhv1idEqrFMqYWv53efE8jZJlO4
L+k0B34PuaNEO6s3bb+Ot4i4lTuVR2arX5svw5/4bTukoOawGAkihi4P7ySI/AdMEYoikr/crxtC
3V/QB1EH79KXo9YjWHWx6MgI7IWBRSnWIuU9mEVQdaslGmMo4RKBi1cyJ2jMNq42Qg50tpoo+bJV
IcnES0FARyCTA/l+YTjyPIgvsSfTjELBaTV7pyY1MSQg8IBiiP7RUhivoKdQiG+3LM3UE3suMw20
P+tMi5UtcDwivzoz0eF6g5qDx0sQzcN1LFPmPhqQGz0YmEvo8WzDFky0hngl0vU2H3uBgICveyfh
YCSq6wvNnud96rL1QCUA3xL6adbrt31MVeqHIaiY0jKq0+pNIy2FUKQOFI6xu1MM7aTuBKdvAqw4
e0J+ziCzo3V5B8T2UoYfaXl1d0cNO9wtC26/eHTndGZzGfm/MAuHjb7Gp1XFUMmvZblG2TdAEKYX
V+OeJo22obgqL6ZL01fLrDBcTc1U+Rzy3DzoDAgiqYK3buuWJlrsxrx5aMuLBv57QJ5KDni1SOYR
5XCadzvby7v+9iS8oZwSuWrYRu5L7wChhouiP0wT2xGtNX0efZLjMDAB/CFVNmEffOIg1eEgm3Jz
HBHTAvZQalQ254yeny70Qr0tDbJMgJIzd4oP1cl405+mgwineqAi/3dIHRKFSGHfShbBkm8YdhoT
pBfHE5CJfhS4ynh4FyKjZwQlf3eJkq++VEpIv7c5kNMFaAR9I6HrCWHrsUzaZYzT5RjC+RrOr7o5
h4HXzpJg1cZCE+E/2W58L+BUcp52NtuzmSm+0HEKbVwltw/XJQ4G1asfhgzrc7AYt30jc6jp9sDh
BBq+WhXR8sUG5sgoZqyusOhELIieTr76+IXoRk2Kr6FPwKp9AHlst9g9q1IEGwMHn/3yYOqPVhDW
TUQi3XCT40VqeAw1ZpIAN+4rE6DKzDmYPvCUjqcahQVUx9rfMeeH+THyhsySsCIUMyByH2ID/9TE
0GjNZzLuHewDicCiWLzeYpmlvq+4mEgB9buvi+zpXjIP9IJNYnS3AHsuY2imZE3Iz4z9PQKx6KCA
HiD4iRTMSaumk9wwAK1+Ehh3D2MadG0EtuVDaZwnaV+nVAVNHUss7Z3H9bZZ1QhwaJrIiU8J+IQs
DAwiI/CALX8TSGw3zVpxpTcKhfRkrxWVh3DZtK6av2wTDb9s9ZjQVLP4RP3hVVxgyrBQDd2jYqcc
jJBKmGj2FF86NY/ZiRSA3dNZSzLY4b1+EQZfcnR4iXl6etx1FEgZ4XWB3qtJqoxOQodACOQvq5uV
CWKQ5PpYgRVPOfm1ZV7F1hlmiieBmffTdW0x4c3IqSfwBhL0z7VpekVFQatSr4JuQJnuylqT3WWO
egbYVtWOZrx//yPWSVGWpizmxLThKXq806FHWluwp2Bt423YfkkoTFJbl1Lc9LyBuN3d7yjPGXbK
mbdTpvIzJ3dGeNwV4uWi6HoCZtDDd3fT2uqpkD46hQe8qH11ntzDC8ExPiqi6KKd1XJvOxVGX1Ww
AxQxV74SqPOSnMLl3nBTClU7IcSC3hd4KH9cNYSC2V+2GTPMkb78qhqiSIS0TN4E/u0Ebk9IMDcg
3WCf2pOz+MVbZqe3F7F95f14Lsl5e3if+i8H3cAi3CLd289j3yAAKvWJm9QMPpdJzEEsqWno7dUZ
yVnrjifV7aVJLGEJXK5kXMlxnRvGRIMN5Kr2revs87ffDwO7+31KGEswC4lXAvKwlJUVTcgV28at
jfNfEErUAIn8X7W7MTnlKkT4KeEswVw5stzpxQwBGMUlgJlDOPYEYKOlKH8azyNBNhM9yILjhMUE
opxFqWXNXqo86wmRhojwaJXvwGi/Kv7J37y2OyDjHYPE/mbPOA4OL/GbM2pR5h2eWz7VXClxnJMP
p5fdZpFO27KSUbZzygl9ZvEiZFBrun1XIJX1FVPapxP0oos1p4v1tgFWgue2myrZVAhTBiN4nJ7U
S/ncUOcHoNaDvd+UDMYv/rHSXUwKRK8cCeHpdwEPtbvMOWXCjsdDV7TkT2d3PoHEtHF9R7yhGLiG
GwymT+sAsGr7b6ssyWy40oCawl0GRcM1NylUprJtRXWp29SKTlnXy9sWUqbYt8WWOYlPjFoWuh0a
sdVlZW8n90p7VYD8+xQ7R2VSqUEusAc6ZjlJ6FVVum6BrLm5L3YnPS36hbQzumTGiuMQQVJ5Ni7k
OcMpzPy4BfViTDtnmmUPqpl1NJT9ntrPCEEYH2wG7Y/nMz0WctMEeuVBkAkKMCfn9aO4j1BCYqdU
/OW5r4uroy1BJu2AuTl6i5vLGzmIRGFNBZ33w/iUQyRPPIWeST/Qq3jqAxqXVg19hASHlcgbd5iS
YmdkXImi1yGeazFGSR9no4orrqc0L7gHd/g27WQeDFU9J9sm9gXKRAMHInlQ3jG9QpCgf0NFlPOJ
Yz4POuEckc/duHPnCfzLhMbM4au8IG6GtYzSaAGYdLbDs6bKR6+nT5ddvd2BS04IBkSo0Emctlxl
GGQ6274RFmZGfa7NGV5Ax2do2ZN72EziXfGpqg0IFlN64s99Ikhn9/ELZ7ZBE1pAOor+pwDnuIyE
Jkm+rjq74P1+ImY+rTGb/8f9pyxBGYd9hvwPJQBwcORYQP+Bv7jP+myfMio38M/5r7Y0NnRLCrBG
voC+cPP0s1XLSxDINV8FB6s+iuN13Tv7kcMYJL424mgjhVTp8A29zNFskWw8h70dLLcnvsvyO4Mn
ZrclHrRmfFqUu1PAOyhtnb9CHOf6J/v8iwo9ht4eZUaGQtNgaLpYCvH0vuyxdEVRhjiyGv/HPBLI
oOqvmjIqOX5fPevD0nUJvOguqJ2feMMyYJAcrL0ecGYChTEDFojHa2G19r6TKftFKTSq3AWRppPx
0nb9FT9AKFvn6nNDWNUnh1j8i9T/ewggB1h8fB1S4gCqWcvO78zXBAT1HP3Zoaa/V7C4OjeYZsuA
jzLD4iXX8MJZ7Kfz1cSWKuZvrEsZvQXPTMm1EbrHlXnxyuJ4t98dPH8IXwqQ5diHNGUKieu9auVz
R6OHLv1Dv4/U7AASTb8DlpTzjn3blAZ3bVU+eDQ2Cs9Z1TxRttH3F1HUPb/BaAq0n8STQMFkHtJ0
vQc3/eBGEGM85r36zzfdufb2MuQyXjp4ZS1yOXFyrv/LjnLTzBtm7Aqh2mqIyOyM15pZGNIRddGS
f7y5qcQj978BuHZ30H86KwN3rrLcJ5KLNs6SZrLjs4Pdz/1VrRNS3PbRMjpBdIfTqKU0SwTCJQra
pah9xRubRqYPSe6brnA5CHrGDsdkZjQh9RVy1xzCHKKfGW+B0x4uBa292tgK40ZA0n+Mdq5RIYGu
cCtUcOsKkvUOCd0PMR3FIki+DoCIepEs1DqifNJ8Yqn71+M/4LZf8VOhRmWs2FByhNWTqHLeog8P
5/QpS3VK5YMrQoF8bPb3cpy+ZtHLpLc9N6t+2IwL3u1FMb39s08LvXdKWvZgSmGLbsAk5k/7gKXc
v2Yelz13Dcg4653i22VjRjjhjvF9zKnOIW2dhQNpP38jO8IkJTMFL9SXnBoI5WvBsJ/TdTVX/nW6
GHAfx5Z6f9viyJ5ldP4HaLAwUHnWNVRfBfmHTiCzEi5gPwQaN7JklKg276yO5a55CK31BjcTzlcZ
EPLZ1snYkssuu2xRbVvDg4bixkG6utvvgErrqhBzYG78zOaYqDanC2wGw/dzY6zCfgE07B+R1o4Q
3/BDLgOEbUX9NIlt5ZAfx0aV7ho9GU+Jl/Kx/mtcsSzp5UTll4oHYJp7tg9JaQGIgkFVUh82CmcM
xGKSbWvMFouTdameWz4SmjlzEykv+vJfZ5Oeand3pzVGHvkKixOEKIhy6NYEvW6WcJ3EgkAziyoc
2n3pQK1oR6J7E8Nhno6IOJJsQ7ME54jVs/Dgd0jacrjmsTaERlFsRtZ/ABVo9yvqTDTiIcuplmFF
67yHN8GcnwhZ1EPmNu64I68o8uA+HGxZQJoGr9IWSst7YNW+Qyqu1f//dpMWWo0YtgES7dfhV03J
XeujvYQQgpeYiZfwLs6Oy/GSrlbFrAd6y778IvZQGmN7C7oWemBY9sgTlE77/4VWYWi16gHA0K3J
s54EItikhtFuOIWFrIjdRNwlDgwoGJ2a6pkbsRsiR9lPKPZ6IWXXCanCY/dcDsw89vUQ0THhLLJe
6wyvTWEMGUpgaOnKPE250Dm9m7jSSS5rDUcK6nhphojE+zq00q+jLHFbsOQhdbmU7zDjDjWyNnYx
YKPR/SthIgz6lwUTEdcvqH/jUq6COykqDMCVoQDABdPrkNUFVrPpL5Y2YowmGlYLnDrRLqpAu0bx
0Yoe2GCE8Fon6QGmKsbUNdXmjn/nRblty62TUn/fwBWwJEybIdCoqG+KuEDZ7YcN5iIdSpQ/btzn
+sdNqKGTO86wbRFvo66rzSB1r/BEQ00Kg3l8LRiHvVeNvv33+NOaishFTNHDHHR+JF115G1GcwDI
8ny8DRq0ChP0KxAWYgK52S3qIUOY7s7QS6BNKhnaom4twBp7K4SVzEsRHDZoyfDOg3i/SRuhhlM+
a7R489lRwr8JUtKYgGc3Z2vVn0p+hJqZOXw5fmjdhtZYVuEwPMztl9ommaDV0FZwgr8z0o3R8pQo
E9Axi2R35TukLvjOiSo3fzyrsQV1YlCK6zLRX0T8H12LWmpaQ+xkcKImkx1ZlUwcZWP/quMU29C4
nGYo8tzZcRu2lakIbmBDLpbE/gKnHx0IG+QtuKbpS+AK+TktxqDxJQhsqhqsTQlgzeIwsYBKKanC
aNHJbnAa8xrHutT21KLUJESuCEAEOtlx/O+qs/Chos14McS762eP8Aihg2nmpP2QF0Z9B9rsu9Zn
3+0zPysDjAR0eatXMM0aikmJDGgwaT6mnEKp1hrBRpb+gaj2n7qsP41rkpvhOl3pthyoLsiictG+
Pe618xKWWNcsI/L52VNMpsfqxTPgNJITiB0JehrPtRy1CquCBUJQFVFnEX0T8FC5M983yrLtuVqT
TDj9SrqA04PIvcIWT4JG0pe1csA0AeVMqDqn6lCmJk/ySNcJnyvcHoqovsbWTynG9eV4scl8oHMm
EAlCZs3HJPHdvJazxyomh0ML4NhhWyJscZNHWUhs+SYKZYs9mc5JrBjOipf1fUC8qo7WZBE7Jtqk
cJdyKecDaUgsalz6WjUKaHcYHsKOWZVi0FQznC9VI1boSy3F4lxDkLWXv/x9GxIUxzfPptSeUSH3
ngmTcNYeUcW6PKaUCl4xeP4+wvvL1tko1aMxiSvMwQOvvxqog3acezGyQBDrSYSiEaPXPwywV2JK
wZ9/La+SlOGfI/ewKZtUT8WZJkb9COs9c88xTh0xW1sg4N7l5/JcvAp7zitbBNxwmvpkf+4Ah3UN
PzcZaIRTmetiM3igU0FQRP+7WmR2DtVz7LBoI4PSIs+I82J5NDJAK4AsA9FY66tvvUNdXp+aG2+y
MHkGkTWHrbciMsiN+Ya4sCY+hF1VciIiqsPutgtH9ST6fFgPp3cx6LxY/YJzAqxlJOHGfoEUKjyl
dDumabuvJScgKy39wKZT/moV0XjjglazctPRqWZSH2EU/VqYgJ6xk+EOGMOyC2UEcp49lopUBL9Z
vaBo9M3+CG6I4mbBcDWUQQUPo3Ur2vApeR1o61iYBiVeLS5wY2OpcELIBa6jGHOwlTTz6LBtCnZ7
cOgsssr02jZCjSrrA2hiFRmqIuHIysTU7Fq2t5Dv5EpgQZ5uqGjBbn7XcwwCB5+fDyOue44YmTvr
NoVV97yrsj2sFNFSE13mylGN8vH1bPaV/53ohHET9Csg7q61MvJO4hI2q4Y4O/UrqAChJXjkMCv/
bfK2Z7PaOSAA3xStsHLuYWus4T8VC7RtE1KS7vXwDwK8mtDcw24fpiHCsxPDvSM6YQwdWaNLp+O1
yx8ZPO3GYuB8jAuGm3hbRBy2v+DywpN8ZfYYDeohB+ejvtBASUENxrJNtrm2HncoFNYgbj3nntV9
D2+Pu/R9RBncDBgdSMVRGYgFyHJ9rls3Iwz2mmaYKte9PxuWdlMs8rzsT96sdkONLXHkikAjXZur
bmlOnuKRGPw2QDqqXmgiZ0dLbkSuwvNWewvKZbxfiUjv2L2GQpUEOZf6Gs6fvaf1sXmEqfMlFkn2
4vQ8StV+EVPvSnEqEm0D41be679/cJFNqzdoslbG+LReDEZLVjn2xPHGmYx9/lyWg8pTuJ3kO+uT
TBatbpI6bbzm/0eyu9/bzfEeAmSCI54sSih/49Z8HTY4dPfgysNiLfVS0YBPQwMtqzvJDL15kE4m
MbcKEluY5NOMmniF++nHsgbiqG8iJWttwHgVYv3ES1PUvzQ0ce/GmBjsgGLMtfWxMu+8H390AWHM
Q4ETdxsZiD2LnwE74s24+8ANJjRpMeasHA8+/XLd17rPtNpHl2eK7UAr0TB+pK3kUkjWjEIaECFe
wLL0aG1zVJ46Y78ZCqbfCj7tdBBTt8u7t7m8TztlI6oGf7SSNpAOAVUqkRxHqH2EkDJObS3XEihI
3XIkAnSQIH2dPJziI5SfJ+Y+PWsMBn4pcO4rhIFE/7LrBiGxqLIHjEJytnU69xpF9Spost1FM9Bc
Y3ZO9ZsWOqpZvAVB7HMVWG9lLbQVMB3gVRnGM6V29lKvHfKcXMwq66IQ0+I0aetCoqTGyyDlcm7d
GuiMHaYORNapSrA617Sy5yIJWIxbNaPUr2QcPgFqEAP8BcxAur1DYu/vXuYOQxb+8IHF1CFIy+At
uJj37KuOVmuxh3k4stC4b+dgAtXKxW0JmNbG1Em+FMZZJUkas3RdULJ6AQFjeOVXWcwIG1kr6Quj
WxxCQCUCLDBGGsQB+zTDXpUqnHYuEO7cdIh2LfOak/KCFVc8aqenPj4i8p3Fou+hs206d09AXrzq
vJcj+l8F1O7u2BC/ozsv//PD7R4c8AeszzaLfFSk/6y3qv1s6lVn77unBInInYs7I9ZCzhKxdlAj
R71YFPhuyW9IDEnkPAEJ9ncF48A1ptLKnRgOv9U3EphWgEy1c0GLFTaISbKLRCqKSa1QxVWWQ67n
K//E3y65dBDr69k69rkvVYtVlk28NoC4C38tuTsMTVcY/n7pbPresNznRvXwot7QQZKwH47MAz6p
S1fa+ANKB8PnyIY7vOLPj3mHfh2T8Pljfrwy5LfxHJ8b7aN+75/cx9GQRsCmfqEcxxUNngVp12Ny
n1DjDig4++9Ba7T1nBf2XGHeTJljmnIkD9ytC6REwttdhOUg2V2FQm+dmOxPYTSSoEZga8AEr8Yy
P7Qccew7y/RDuqKIC0ytHiazAsY7HDIyoQ5VONUHy6HddnqXJaczBE6etogwoyBTl8YMtQZT3G+y
b3QNnrf2DBVxVgdm57mXvFO1s9Mm2L3ep224zSFaLmNKBR81NXdw3++rOjSGAARxWmQe00V2/5P/
Wi7uzPny8RF6tM+hEWjR3OQYe1V44FZhn3Y8JtXvfzdrZqfYRrBKXBYk8o6Bk0hLaYN6DH/QAnwq
6mJsezVyo9sngSFNCvABw3aSb0Vn8nYhI4rRZlh4HluIJe4KZvsmShhA2apl3Fq8QrJyRAez+O4C
le5lZXVQOpx0wsGd9rnuZ+d+RJVQ3T1r4piG9XILjcEfq6qpgUQ95OC9HfBMFxW2Sd4dyHyWaOpw
CiHuTvnnLh7A8cHo1j1KaeuX71u8FrMO4sBZQTmLB48Xg2hnxE3hEul++ecbz11tShQJulRK/0+V
Ssj+ow4tw+SV+QmQBanlGLNdsxivN94bNjBpLyzTkk7sqFm5Zl5ifhCIQ3D6844NKhgn2rYPghVU
/OFBG+/U0MR9xIRuHl28k58sVVnobt7xFPJRaHfRhqo0qfFWWZDJToIW1EaW/jMa321dTsJ6uXmi
2bMpSXC/IJAQLyQADqmGIkF4c6eH4TOpUybhHDHIR/37qJpaiVhUHeOvwAJH8v33Tz9iwPR6i6XT
+5ZpoEbAlPXJpOLoekNODiDiToIaS749lCMcP6wmn11mkAVTo2tNY4RH1fJk3jEBZrOirG/3a70D
J9LIZBLFxMqcgUJEkhzNpmgwEFTmZcZHCdMpCOVsB7hx4Hld5WsUiuO7FcAt3DxEWTbuKXiMFefl
ZcQF61IZ4lLyY7kQCqFGH/1GnfmDnWh5CI5M9iG32TQH45QvtdMfu6hm3fCwqe/HaJA3RX5Zqnrd
NpbLR2zAjXcpzJiTGG1twtBTB6nnoIVmwYsnU5onRvX/8xO1eqoHDf49YvaXfbIJ5zmb/ShMbdEH
FevQDpP4NCSc9gBrAkpcHA7Wh+eWW6LMFn+6cGMYKuPy8dcPjAKPE/Pm3pL2723jMmmFILzgBPNI
p/kRpAP56KsiQtglXeVKWadBiUhkFZd75kgF241JxYmK9XZnAIp48Z3epzkXl6iocAMQT2R7LE2i
JB4EXddOhMyD3ua6nn+y8jp4laH0PVBgbPrXRGpuma8NNc60yZ9fe/cIHQNiNGC5fb70A3QuTk4O
oBcfwofnqxwoNlugwQkXzPB4yRd+MnqPPdNw6XD0K+qOl9NZnSWzwuwxhSyCxoxYN/JOrhOVB8qe
ftffaaFH8LCAO38NLxBtcQgZfDzajTiE2IJMj1cpgR3IT4jjGtKXQPYYf3mwef7Ydoaj9gbYQM7/
4RrbBk0Y9Ef2pYn8uXe4mM5jY921QNWGwdt+WZvkYRIjJdV72YWPnC8aV5HBMmgM87i5KG6h71jS
/86hmj1RZUHx9NwDWum02ez7v0bDFsU2tyWeVBoHuZXJMHa+Rz86wHXO5qXdaybDixJ2ODXlmxSN
awuo0KM0KH9tiY25i9J5LbErBlUhVTkx7gG34aM9MZ3aT3wAmJ28ceiSpH/QBlLCS+zB92IWubWJ
l0Qtjvnr8RmkoZudGZqS0VXmS6CVq+sSD+/C8Nj6cWDy4QEitW5kY6LF3ifGGC9Uj0ptMgPCVO8W
4oTWpJvPCfgkifIOPgGfUfNLCUokbKEpUmDnTt7ddJo2h7t/31CLL1Rfpw6gxZh47DXvHC63h0c2
meTpT8DzrGPWEuvdQ0THXXhwppkerVesgHUny8aBqtyk4HB+UfV1fGWiD6pSiZYxFZkfiq2Hdmj7
ixdHCt0Iz4Zgv2vrrs5baVP7PuEB/FkEIFebs8ZRWIYRptrotPCKtdX3kTlQ1A+t6tJEXyAuBbX7
FT6zDI5tfDoGT03kybiI5lzXVVbPSa1skogPkndhBVm1/N1oyAeDoDv2SoXzvzuu82AswBvzC4ZK
Z80qs+t//gO9EHpScKwBS5jWrLZCB5HQ43GAHpjibr13TYm9qsnW4VpONgE/rrfAFdO5mQcIqUg5
PkagzJYaFl4MSjXsmZHy7LDWLS5xTZpYagXsMA/lYBX+AhlFjTUWVLeuhYRvWwlQnB1EL7z4WkY5
H+rbLLvabDsrCCKC01IOLIPKjYji2/kmbHA7CnZF0tCt6s8WjjbjzjtCATYFlIippaXKJYULq74m
rjyCyKlpND61t/bzcZEe0m5myP4Gleq8f7Goyx1NnHV66NldmeIHKz3bpkILm9Ef87jLAOAnAflP
SPtc1UJY7Fwub7FHJyj28XpY7gUz3gUWL7+JlakBkQSfa9O0z1wt3iZ53Co5ufm4rUWRo36Ujcpr
M408djY6mpvz0WbdGMkcoSJlu8+uwQsaUKPxexD1AXh/dAUUYrtq1OxiQByWaGr3/b1GJreC1wxS
LEVNXpddxNRa5kcf4okABQU5bJ+6kOxZupqBRoK5UJlUp61cqWXXNBEeYHHjU8+MKCEut3yJxa90
KZHgqDAP7gcgLXhkBnGVc1m6TnfvWpHp7Mml90VS83fHomCRvvKhCVjEi++NgqCLrIW/jjG5G24o
BvjCmoKOxdtpJfaPZB5GV7TWuJIUK8D+HDo3+0f4g/RBVgtd/ntMsnp+aJrmn3EX4utlbJNhfb2L
8QdeUBWRnhpTsXO0halxvY6q2dVllOZmH40oakal+rkuh/hkAkKt8fMjxzr3JkTWB6IjhU9TweIg
VMSMM5wKVq56U+CdjHH8hRzdk78phi9TJFealYYzlS3EYNQ01qDN+drm9TYc3jc8d771xvxT+1dY
Q3yZBQJ9pgrDQlcg9SFpMoElBFAM96c/wNXxyhlr/K0+nyINHq8iJv7QaEbNs1NzlrPX1xnvjtc0
bk/Jxp3e1ajsuRB/x8SrdtQJ9+bPxWLqSRgJARPMHklBV04czUDw7qJEKrCnzQPbUcYngRJrJjT+
nI18DZUCACmCDFW3VpjnSyUlRoFqmfa6ayhgz0wkXH1uWHcv/ZTf2H8ksttJAS7m39lqYDShDGg4
87K/7t0HUkG9SDfevzou3WP1mkcCQH3K5pua+DSafy2HqN1x5VM1UYSDdB/UlZw5wHL0GohWjpMZ
sWQVC6IuMUJbEguTYJ6XLnreh9naxYgGWigyGORapYYmxyQw+Rvago4OFGYZJfJQaSpaGX5mFOO8
i60e/UEBkdKMqRSbUz7MZtx736i3u+o9GPyNlxBUtSsfhLnwnKObpmg27M3G1jNNB6/v8B4mxeF0
lWXb4/7a6s60UCMVSzDZzZvuV0opJwpJFfrC/T6IVL4LYUWGK9/Ep2qls4n0NVboyfOIgg0oo9AD
eS9pHB61J/Iym4sjpV18dJNZ9avGrQieKQ3AuZSE5cmeH+w2aE+GatIJiwamLkVx5RUjZvfOAspQ
U1W2gr7AdpLcbckb9VveKDu+nmLTw6TijPl4hj+js4iZ4xPtqjzCYv2qr9uZxmRyvwt73q6zA0+m
LCnuM3e2uvmbiNR8DlvWsZvNWrDS9N6AG2xRqlWJ0l61IVHF7ri6j7vvXhAUk2wZtUdLafyXWZJp
6OTwWslCs2AigmIvYn8N2QrcP7TrTsDYPcY6DZOO+mMul3htUMxhZtqYXjUmuOFxGEfjqfr5Xj0W
bjMWZs9w1HF5HLGzrkDpThLU/WqSPmNneXepBT2YcSmvBog2loHXUNhxbCjz/rh5G8reXnL8tcgC
NdCpaj/fSpjGN0cYhVtxsmEmhOnTqBgMs5SzBcOtHp8WPfupgpH2Btn7cAFkfeGPKFjWjZgBY+Nk
4by+olCZsMfKnbgC9yuKPBuQ0fNlD76EMNGvuSMl4SXon6iQcKciA1TvTEEzuwd3S77XARInzlnE
qLdq5aYEpxs49NJcdzzc/c5hVGPg5wfHF2OpaiGCkaDTj+2V/YvPFNtJZscaVNFHPd19ak+hIfgT
RSTwa2Ae83PORoBc7hMDr9Qn7Iqa8m13JoUf9QpPI23b3EqdvtHX4MB8KNHM+ftnsC0ToNlMIroZ
aCq35jJMsHUaQAsa4UcON9ysRkZHSPepGYSoUjhpcMgh/kZeiYkWRu51lBdNta7zUkMMBCduWKqb
y1zKW1BLTzg0Hr/4CL/yBsd2WLFAulgTDpV8R+F4nCod9wTKrYFKae0FG82EUXpskz4aPwyl+WAT
0QqSIWSXvNh0edhpPf1HA1HfzyGg9HKtyrrCe5sZgFZS1MTFhyelil+R5K6eK434KJRYCvYMCvGe
hhX5NG14E+WZLWdwnHSlUiM1hKgqS9wRage7hYvTQ38I2kFe/d3X8+LjS3rnOKO+OfvFrsB/V9gu
b4PwPVbGKjPg5gzCqZbqncRAHMZI4GgGKsecUtoq/YncMCdbclZhlADpq/j+Ea9IdaqEttkuFflQ
U2gc1hpCskSAM9CTzulgYH65Ix7alo5vTHHBSlU5SQtQqsVWiAlH8VKS+36aTJgzYlblwtdpG0DU
tOITifHWY3T9Mw6dyU1Kkwqbi0F8IsBvrPy9HYsY4BE9qWrW5COfAeG0ohYvCYfTmzZc1cU4bC05
LZHGJdfZuDDDMm9qu4wh1grftbLr+C40ar4HoNOlwu7yzA75c709L2MNQM12K6G5juB/7hW4IKTN
OWd5aYjRMckqYwvv9HxPtgFnKBz78I3WEd/3MWvvEzD0JgKKsfgPYZhRHb4iX2ymuk3S2in9YZWL
dEcMIqI2tjkZ7UfthymjcgCLsOwHtPCTRsn7ZLSAfvqYJbVVbv37wTNo/6LfgfSRB867NfT+4pkm
gwRXKJzG2HeqiET1f7trd90sFCVPE+snv7Tl4SsmiPD+K/EMqCMiSGBwxIolf3LA9r9ft3QubVnM
0alW+KApI87ch8Ph9SBMo9t228gE0IMKIUj3VE3/E+INMfN3M8+mh4zeSClU3RVgctevmQfbLP9m
gJTNnYmZsDLE4BU569Auz9y37wJynrSdL09C010eXdezZJ04PqNrzm44uGqTp8hDpy7bIWsJ76ih
gz2s0nzUXWbUk3K1VH1hGSOm5d6KCM/8GWDw9NgNoDkO475fppmqYTgHdizkWbOE2DBXsu/B8pVh
gGNpzMk5uDZRifCND7ZBwO6dJG39WAwvscmMtVOfoq/cAPZh1HBXjCXtHpI+U27R+4UWi1CwMzZq
3yH+aYvsDOmeRng1GWry6vdNHpJEXx609rulyydEBwNm8mUYmdY9RBaVKGmg6eWGCcBKMJDvmq+x
vYOj1wzoZoqaf/avDRZFKxuwjbBi7P3Yt+YTKzYpQ17M0miAFwPKS5H7WwIYYsXaANYIsghHMYNW
mxUCCGLpP7C+c1RGcpt3c+DjRybjx8+a27HNMq+LEt2KJwI+J2JgV+3Ab8xJiHnMn6aPRC9RqOC9
GlZskYEbSzG89YvIGHea9a5WIrPiCcOFkZeu8BVy0X79YyfBwZNDGzWp8KW21w61iVWNy+r1NNe1
QcIGBq1jPzk1UTS6N2ywZUVDXr9Q+gbtaTUJUsmW0RdPZmC6cnA3W0iqQihFGozKJiCbvFxwsn8/
45Z9/oa445B3sKtZVsD03FrZwSGxTvaBgEBTYr0HDVK5rCkGMbKOnO48ZA2Ojlzpm1LivbVDFStN
Qqg+aHfneFhRbKdWFJHEUdMTqfereWZ9nK5/Elr8Lvq0FmnEuxspTKTI7mSXVK/6T/Jw3GpnEJXt
CCSXTkGG50n5Q3KosJFP5Pj8mKMSgqLaG8T5OaEYq1fCyLKVycdAl7GKJPk8yRrMp7pnq8UOs/yM
pI5GijxlwUX8oBG6mwfKUSU+SkFTZOeh+vjC77qHjxjk0qJVsotAm+2FvpYfqdeflcGaZu+C1CVk
Xr10291EHBEfvbRbAJa3w4jtdvYsaBeBme95n/HYZeEOD3PnyKZGmEns089xyPW+O/BKFoholqVC
nbDC4Y8S5vy8jF/m43eJBepWXITfO9PN2drKZ7xEu8VE6uXfkh21nY04/0gty5OpAoNgORa36T8x
oLvd2s8lA80XGFNMoFOxVSGORxagemW/lzQDoLYk+z8sn9+uxfvV0AqGgGs+BO8/gVXmiFyx4swO
FMek7dkABgC5SueU0aB6w69tmUtAmK87D7QS+uaLtc89WTLrVrmqsEh+rK0HoV/3IG/N3RvrGzYN
evAo+4AEhG/f35CnTG5RWdLomdwul0gpTiLUUopzFWFlrDnajyZuO5GUFjeGpnMKUuVFvPK85p3t
qh005aU4Fl0R22yqJPhMIkv+KawxqrVjxtaiqdm0vV7d0EopBi/YWquNw4Hufix7vTeB6uMP5ev7
+yWcUyFUZbeWY5NEJEZibMnqSoSjH6uuh7iPUOUIzvCvsnwq3HA38UnV9NVDZTlwEXsMjhuCAsne
XnRjEmGalr8yw42FiszvSV2MEHxCdDQ6i7R+xlyTScqIypmKJNiJfI1XSZ0KsBqFwKCv1yKXo6Mm
drrFV4f0CPYj820ihK/zAsHdeWSkekjXCMjyIq3GtWbaR1W33aBBqqiSbik/kX9PACVsE1OnOEx2
NzIJvVUmOjiKB086c2/kHtZjajIixl/SG0q6go+jfvKRLuq5bV0X5xlaN49v1tvNfQuwPKV1uio1
xSIOeOBXpXIIB37xjRUeOaTxvvASWqKJDydbuAdTtRcMqq/oYNWPtwbNDqmc5n4oWMbCHkV1SpEF
BDOQ4w4LKFBM4Ncksrlb25Xi6DnuLLECwOafzfD+NYAqGNgtKQE0zs0itzRuDpdUBPgSdak22MmH
qd40tIwpWdwozGo5ITfvNyNaJqnKgc5sLy46ejUNdlBhRvkrIN18D5dORWAag8gGp3mTRxP1swkN
z0baFIs3VXqRjbMirtoxZNh3h2grgoED5v3MbxJFlGcpL+uCjJ1t9edzNCwz/iHXtxx7/OOnopUR
Nx3/xty6wKnL93klu/dmvmX/TkekwWkHKoSXbRc82F5XOVME6C4lCXT+aNSC+Xcu7RSbi/xzjlp4
x5VAZf/ePLItBSBImfJZ0To930o1ei7+/OVN4hN0DaSUk5J6sC7oKe5niR9fP+xd+JvcZo9V/Dgf
RnLjoQf4svcXFUBtAJSGTZp9Br0U3q+uBDRHbfwhN0lg0nPOg4y0E4x5nqd1Rz51n1i0ApUUYNMN
G7IzqwoYr+4a1AQN2uDXknzW/43ClMBF4dwpGjec/GcI6Eg6noSi3Qw/gDL3eTryUZ8MrU9RnaR9
P0umgGpOwUeyoiI93LEF3MWK+U0wYa3HmKMgefLAg6yvZSbuTpzmCi/uBxijE8EWTyka3/yzXSz/
Z8qArhE59ecn8B1VLrZ1WhjLx0HWP4FeuRt1Fxdb83vLCsNSSH5KktLALrZCGgeJEyX2D+wjrIbN
lz5HRKrRa4powWq5GGeQ7ruMAUCIe1SpFuP0rplL5MC6/JRnBSnPlBdLdvOnPeZlIoiJFXCnlIwu
zctQLcG77F6g2TtTHJNb787OFwFUtlv6GiCySfmf8jIsEHGkJVFtV5ZT62lJAfpvMZYqdXcjpYuL
KV2RUJjWebA8bj4nnLhzV4bJfP58Lo/ClMsTJary2NrqLhh8OEGqxFZD7uT8ef0pCLs7tjs+bppj
Ehu7zIqhaPZRZDANkfyLkYmJe9iY097fg650EGKnEnM+ampmZVQgh4Vmojh6JQUQqW5lX+8mHeos
vANOqSEhIGJwAeZxJUM3K9yK0NDgRVA30X8EwZLjLvts3sceC+LAc6CzoMTQ1eSN0CdatFc4g0Bx
0X42w8fYBsTY0PSpW/x9JfOh612F8EARectnbhc8dIRUrq+UPhg4eIWVCaGAODXz2vOByiJ2cO48
9dzvmcgHJPfkd+UvA4CZzAJTcGRTmrO0pxxxFSuOi/aOF6tI+yFvwdaxnJz07kkoxr3DYGHoOhuv
j09jJ0iVsEteBfhcycVSp/SohokmR+zz942p3JGOXhdQlQqZ9cC1S1nwSNYxMQ8FSJU0dbcomvRC
rzDAPzr3AqO2FIgErwtn6ay3Ta9zSFRRRqfiFgOZ0sirqNQYVjxoFbkenPjNSaRw3imVtdjYMCj+
lSO5CT5A4MCE/NowedJezB6Ku71izIE75ZVbz065cbMWJV+NDbbFJRHIdnIxrmjOE28Wm4Rf/zpP
6EENe2ZQIwnqizR8hndciWdATzmCdJpVr8uWh1KgVXFyp7MZOJUfh5GU5JcEb8n79Ar+3qME1VUy
YcJ+Z3SAYGh1mUNc6ZYcKNMtpqi5pRmt0Yhnc2umRJmeq12dMdf2Ii9ADCcQOqaoubGad0phxmR7
YfJheIjMuSETbqIJOrBu0sAUYmWlrWDb7dHzhFpPtOslca2rMemvoIsDxmyCc1xDixOAQtBB/JpQ
rgqKyqUIyjFPVRFJt3F9Wd6AzPkQI3ZO8Tz7krAtucDuSwvAtGPXdzf+SQZrRlQwbenXwAA+24bD
v9PhFRIF5n9O9R6SQeaEo0SL2by2/A6bRVv3MGetXS/eIy24/pm66mfu0gVJfiCiggDZQFE1yRiY
7difS1g6qwZHBgeHOdkggRNaFyoXr4KDTyJVgTLo9foO9/7gukUyp+l7Y7Wu0SPtJl1YJOGyh548
8sPt7aGwoJUcc6lSJrSOg1GphSnoMyophIsOs9g40YA807RMAiw6DyteGx5u/iuyccNhallsnh45
CC6i4j45vgyjyLVm/A+kw/LjkZLdZHK0J+JTYWa7PvQVymo2KMtCqXaGK48h0DdKbICEyO5/TrLU
PrE/y7qtHXIEXKnexXe1H3jrWh8pB9hav2iFx/Qnpqw/StZxH/gRVsalSGsozPgf3obtP2OTg7Gx
w/F5qTGB8073O+1f366oUpntAVMTXLJZe7PrAeouTdBbfb1PL25ws8tXImh+ENsz/zonugAvAoq0
Ae6KhuI6IA9h4zm5IZMFh+ClE5T2k9LVwVQxkExdxKncP07ARI6bU0WTcGxJaHLCbijRR3AagtEa
mRfni0SgrRTO1a45uEX+/RGHxpd80bgkR34C2w6F4wcSiddWpX0I/KORcYSkheV4MEQmefok8bH3
icyLAJ6J+lSgOsIagpoprTS/Ucer6H5xrV7wDruttxi7LQKZkGfcWXDrNFFK8QXjq8hyoUlAX689
HAmoxHi3HAfSe/0BjtruoSVfHULTGATYPAFh+LgbL4zd0lunHDlvklDcta9Mphr91kb5zgoeQAPJ
HjOL3wV/27ov4scvOUC5BXj/m9G4e7lFfDC17t+Ba84RKYnZS9VZ3MqIwz7xCIrW/oHXZz0qHfYb
2RhRbykQM9GBs+KNmTQuALMwgQALl+BioQq0QaJ9TBTZftKpokUD8QoMqYVcGbDlFw0iVyFht0R/
xCHwYfR+8l9EXKrK7gmZYb9v61PgXKqY7RozsZzgGba0AacsR72bY1i8SX56drto4krRFh7p8+lz
ndCvhpmPRJ+liR313gHgq1eEnv6YDw+EVSX2JyQ6ftH3ofOsZWEmNHrgNWlgrAdgs9o5tvU1gHqh
dA2pz4gJ48S9BWm0JUGeN2ZUDuxL+ejtEkyN+d8cYRp5mSSs3eaojk1IS1suVpwUj6p1ScfERyQg
1tDvmrVW2teyZcuPB+LS2Ut/FJM7JH0UfGUhUKVhil/OM+GTq/FdSe2ExNYN6zjSt0K/tgaB6jWZ
q2nqO+Dj4rWZEBPyV6tRBJdmR5Bqmf4EngQ3HXThgs2hYe4CHPiUsw+Sr2+Bq9oHcoKOYG0GnbqR
LizH3LU3lRTFSJ3jxawsoB1vOiHh8raKJqszLTjOdHKJx6zqgqN0xnshn+w5s3/bZUFXmNDoWyCw
U5LLGAHrHoSa8YHA+p1awpl+o3ZAGJKJQl+16iP4WN7mxbP9UjcD3VAFFbBx1Z9VPzwgglm0c08+
GRXJmPEZlmq3WEjmWJfafYXU1u2H1gW8LpdybPHQ4Xz7TAjk3R4vXdds7J8oWQabsuTNwKLppANk
lGzlLWl1vbQ8E7HSKJO8JVcy/mJJRKuIvRkTKugfRT07ae1cN9AiP/X3pUaNyaldS9cj9k7EHZju
bwysdFufXXIrlMllCqe1gE6nKo0duDVNOfGEKq7nDlhAfFoo7G1FLeDrfLUgAmpapfDp3/ebA4Jt
Tu6GsDZsJIIi6gm2I+Pq7JmZzTkSh7UlC5e3/7g8QbPHgegjTpW8kMKslCzENYPrvNnWEJLJUnAf
AaigJhG2oI7/VhIBvXWioWnIA2jLRKsSmnTIy+kovi42gqtPqMuufHstHiF5zM6aaSYBMmkAkniY
z3sqhS7XTSA8EnTuywWrFec/FUGIemHiOFSu4DOeYApUtm2WiBKF9X27uIa2c8lSq9lpGC6wOF9P
oAU5hJYKL1YwHxqGFkfqUsjfRXp1F8NAHEtOi/kUoJT92fyx79ywTm62uZuSo9fRlRcEbkO77m0u
kZ9JVE2E+JS96OpCfSUByBOX4kQ5jrCCtbrWrm+exZpfjwdof9LkJT6ydgEe/wqt+bcnf+TQ+NRD
aq5Rig2OIG2nu6Wd2M6t0rBO3BUpZuLxmu6hQASwIHDVQI3SXca7nFLZIDRJt3Dv4Ox6OfFD1PiJ
AM3RNwsh4uG1bbCXLeGH0m22fNsnQ9ZclAumvHTSq+HRgwEY2nZIukDfH8YkfwjSDwH4hWXJG843
8At4CXzcmldF+vGN+xnevQdIJ6w/2G9YxZAJTC9QxPaAAL64HkgHTk2kFoYmsfMqWtOTdXYnw2xD
RPr/lq+Ifkj/yuUV/phi9ZR2pmZRu3XwUat6gcJvOIS0xeBTn6IPAB714/7htnrh+Cj8icSNv9uN
sPdO5jd4Qil3T2mmv1oIuX2gn9lYSj9BVOLdiKL5Q2wVrBTh1AOYAliXNNUGfrByKyKGts50zkh2
amhVSAzqGw85bkqodT3uMttAkO9Y+pk1c3GUgzPi1ntK+jhuUH65zKUI3clOlTbo+X+3epNP4U2G
QmxwKyboMNsLXQI7xQyMAX66sjTzdJ0g0h/mdqq3DGodP88aHMe6a6C4fh0jqwk424t4rNGDf5Ut
Dvoj3QF9c9EWQBEHLt4sXCviiZMu9piBjjFwM6rTt1cx9knQH5NyOvC6w+CQjbg6tp2TamNvJjtr
F1iwN3h7vN/+vFtoO45//FZwOmS7qTzLey/4w+AoWJ6ig5L+k/LpB7j/oQ5dBMNSH8vAdJNwhURq
fjzLUJdtLROTMzO2Io1oC5qlWDtBF7xyWjyGbdQlNGi9/12A9qqNkK636hGcqXBZCwnMfchZHGJj
WBUH1K47oEjwFgZEIEhOE4HKqvxF/UGfzMMHYq2P7Ith1cIpRosZURtS+C3lsyDQ2DEvlaE+NP1L
W5BBMgl/W+AOVdfhrwXlLCVlDtt1G7FPus7TZucH5Uh72M1WnMmADBGLJhEnro7RUwHgAFlLgWVZ
61Fu6+ai/L/XqNwIZ67Ilgo4T/VTTKRsexf4O2fAAWv1B8aUBaAhgKSoMM0M0PjSH5yHOeQ/Dp7i
8ewl9yVNjJM+45srnuXatwcZyYBgkaxlGgNbPDgvUw9VIYhl3h7POQpQNJ2lpMA+D5pkIDGGiPC3
UPzmffoChTNS/ZhD5r5RkmGwZruQBundKFx0UXmclWhDVK1ZE0tzEejJxSOHgxg3sr2PshCDzFd7
beX1b2q+2RYofEZQ1CIH5Gt1DlGtcofiihZM0bn1l5mPUliOuRSglGlkn1X8gr/IrrQFFpyz+hjk
id1wI9ovE/49tSJC/Y3/O8K/KJelbIFLB0VS3rHEVulUNBz52U8SdwwcwbcsGPCpMe2u+KaoD+F3
rBtEqnukjzjwd1nTawfQ6IRWYIAwnQo+rjkyGjPpBen1dtntJipTp/JDNz666phiWy5v/AjgLdJB
iUeHPQsmnX39jcvkvfuFhNUXXIFSwG+Wq+bVyfUx9ryn98nJfu6Nsqgdir/1cj4KYaKlalyf5PQ3
JUCjvYVlh58+ahGtrI6lfbNG0pwNu+A7eyyjxrFdWpYR01qdx342rYlpkk4Vyhny/6F9TYgoTudc
E07v5Z1372KaBOHu9OZOlVHcBN/Ndz6UVyffv/6qhx6h1+Go9s7Ek543LmJemkr2Jv/cBrR6Zdu/
Iw3Zo0c/484+2YgzrOXHFOgxSYC0UJ9fV0juAuH6/TEVU3/EDV8eUpH2S1CzMa5el0zFE7QzOz7k
Q/80SA4uKprN7LL4KFQG/Mn4J0q8PvqE9bDVt+uIdhA6e5drjTQGZoz8f0bp/3kG7KYaAgCdnlOW
2ks6gIDx8d+cGvkJfOiVC++u3Z7GktT0eiSD0fxNUDrF6mmFzgwsPsMeQS81+E5rrRJSKuev2aIq
O28qOkRvnkIsJ/tYVTdHO1ivPKewI4uGhm+sdx3foIBy6oe4H92TqbTEbU6xiNkbvF86bCxf0hF5
CF1JQGcWqniJxpkfr5uCjI8MV3O3U4nwC/GBY6BJZaq1OXZup3qUt0tztMdGWb2vC/ufSCq4/hLL
vMzTj02FpUxcgTELRdGd7rCfTcAEAqd/WyprDhfsFSkfit49UuagcRkn91OEEGW+OjbLJQgmQUQH
csTnAlfTLkV/orfKnziLctmlEgEqYcU1v5BeJWqgsJudzbd+FKyQT+1vbWWzTUYgPtm6quKeKWaG
Ju4ndDov+zIIcYS35i0GNmPbZikRh9vG7TwJg0RWYRQ66AkGDMngOoQv9ydQJ/FD20hAjcNynkeQ
GnFSymOezwE8cNOP/eRbSYw2IodzgkJ0ZUc2pPCiJv+0E8p0fF03SIXyURn8CRcoKJvVPYZOwzpc
na8OSDI97OjJlCVxPkIXs9EDM0uF5zp4PjNolv6fp4+MPqWIk0vB3oKcz7eOxR3+If98dTuXlWuk
Hrz033drQRd6GJLjNEAmUnPRKssIk+RXyL0iBmKQZcHE7iYCj7ztfXr6YRngcFP39vGb0IhJxYsz
9UrfQP2vEWvAaNg0PVlhT6ETiJNsLAk18i+7wm3YuW56A1PM4mRw6eAI0SEKAv2YhZdSlZ4D4i6r
78k88Ife/J4pP6RBFcMD6qthVApFAsk3xxgl0lT97cd8amOQ0EljQ5TneM9fOv6uf//7nToucyX/
08jo/ArsAaD7Oacqbruk+ALy3jRpqiNcibn4G9/gMTD7zBAr1f2jh9Zned1nnFDUGaaztwlpuAli
rhuEh2q1zLFZ5hNbqbr7xzvj+MdbodN6dC3TVY5J461ZxT5NRcQphebULQFt/ZsWCGWSG0AhQ7eQ
CWiWMPr8uofSXkgtpfJbgl5GV/Jr1VR1RJhIvE1n2TXw6swK+ZFpICqaD9Iz7ML0SrgVYpW7vvhr
CQq1Q4lbywo+GliiSXzpGZAqt8b+wvRnBX33VTxo7vDcp+cB0aonXj+ErasVGFHFQ1AI3sDBpzdK
xC2HsGPV1h7lGrI1jMHnCrGRMvjjlAg3JFGw2n4cMjcI49kX+aO2xMPcIzmJMkJFrYsZGb2Ombh1
lP0MFHbiqfC25mJYPCOqd4lE+iofCHObMbzaH30Bsa9pTc3hvCgrq2errkiC4iVVmJHxxhT2j87w
OJKoETltWk3UXoPOYHpvN/nMtBms8pXo0qoHxooSL2SAaSQwssI4YQuKdRSK4fQU7PZY+4boBSA9
DDRZSL391HDfyGTToWWOTMdL5y2Su4zUnPbBzR/tU3t/Umb1k5mexNunYUW0yqFr41RJsVsktxvU
jTO3XY558fTHY+Fb8wv3MlJM3Wts/ao1MivrH0ZDg23aNh2I4casB3dvVeiycPaOAOyTqnv1AvBA
YLHQoN3zxts2thUsRXQBatNtl+Xmhj+DvIoP2Qj/kJ9BFpYMsdxwWdcdZUojy/IXcFPLw8Pwka6X
gNh0h7q6Kyhn2i0KO0D1bWB7cwFN5gS3BRzlz8mPsUsqu8721eyc+1RPnQGrUDzKe6iQ9zYvu4RN
1eqjbSt4xkVbWutpn6vM/IkWvgIOw2c3gVdIZdOiaHfr6G+21hY5oqKafDyPJCG/4L0xdf7EtX0A
Po/YG1glVuazuBtgh7goy53aDFm6sOScKY4e7rMdw4NaI7HWYaEgOl4PfGmxGf+oUDqfzkeWRaun
PF34zXTor2wZUM/ephC7xHYXJ26Gomrx695n1pwYPd/Yk/fIzfqX0UJ48fzSzY6rV4w4kmdLKm0v
W899mjLGq6QOKMsH5DIeU0r7Jlp+gqJWloQajTWAF8WGSHJjGcVxrjmWnUSRqXbHvqYKXcO1214/
JYvydYT2htlOOPaS069AhhC8eSrCZtEMw/t8OHHJdfuum93NLsuCg8emSaSCTx2SQKSH1oWL7pqt
k+yKs3kYT/hJGPukkucHcIeauahz5im7EtYCp6HZZoCUgtrc03mo507Mm3ZAt//OlVHp+LJQ+PAN
bA1+ZKmhBA/ag3Re/VIGvNY+GAVS2YmU5T6UxOVZca3aiD+XwrpsMw9SDDTr2n70ZtTydh2svuOk
R0FDbk0OzhxK1UazYcATWqaFUNEGCE8ZzPixO4Z3zfJs6bbNwKnY/Q2/Gn7M56qzaN3s4U4SIyMl
PXNKyNsguIuKw2xYu7iPlRZCN5FBZEGBpHiLgkD3IlBNHXRjI5jDRL3L/WdMkQGOcVAJxJFKva6U
ySvnMOdra5AEXFMfu0QCaT2r38KSCr+IbFJv0TAN6SZAZC3UI17WOoIF+p1iff1ypy3oL00Fcvnq
1HtrUdejl43Bond1ujO9etwhuF16ei12kNdc61HLehUiGoYoFhnDunvFLVy/zZ7d2TLLb6ydcVuz
7KqT2J2+gVq9LiXeO2kBdxYsedXjaGb84FVmOdZO0E0LA99LilLtm0WE3b7CAb/IHf8YHEKDUtOI
9aKCNxMIGrPDeIMmtX7qNrD3hfaL7tWdfXGl6aGyA3vZ11FhNfant0phFDbBgWeNx294bXqcudxV
7/JUD1K4THcPawZ+wYhjSUlB00v74zAP0Ci4sCZUG1O0eBS+76Sn7s6VqGp5JDvwbHEXFv8hHqD4
GbTYMNe8CfDffh5WELWWkrjLYyNkahhPq6QKdOfWoTnZAhWs8cMDUCJwooKDy+buc4ylxtDja8/7
fKW2ul5AZKg0me7ExRfVwYn9uOU2bjCdX62V9JR7Lk/CIkwziVpBBzy2Y0L7THe6ULvD22oWYLw0
jqCJtfZL853aKQTeyOFivj94xpZohvDbjDhZNFxPrpWtS1t7Jp867Vw8LnrDmOPdHH1boeDBRC4U
Y3FAFnqY5Ln0lCPJb+ZG8bDF80VIlJBgrOWptk2tiRzFPhDGtUS8soIx0GbPY9HjHCJ4scNpWqL1
XrCzjRWO2oMPecxNYylCsspgKMj3jOtb8S5/dGmymtKlWQbFX8/p4SbhBGT1PBAbpNiXFADwktF2
lyzaY7LtsbeJOGnAGfPnApxbmWQ8vXaqL43iHHN3tUv71cqEkxPyJfCqqmNoZuZikRfYMjLaPf/a
m23+QgyRsmv9bfmHWyL0IvrTe7k8K84opOrkMGbkDOLccbMSdcv/IW5DZpVHAdFBqnrbhSDFA3B1
lSzvxxm0UHcn7NGs3M69Ff/xS//TdvsPMIR5prL4DYMjHCqUvkAO47FoHNWQgruuqhqucsRGWzHR
eQv/v0swR87eCuBEI+X04LOyepEY0cKeaK7bFtlezyUADenwimbsvfU16xE2E9lb4T/xzj+auYv4
MDXUNbRuej2rNxIAa3JFGxQysuXTliZwoCaDnZu/yqFzz3j6WHNiEs/eGjIka6pBBG4nBGb1J7hs
mLtGb2KzxTudXa4HXBrqO7WMR2Kj2mKUFHZ5ab/GFcEwt53S0HNg/yQMTgiXYpmEImy8xUDYuMjw
zd9y87mAQlyfQ/AjVgJaovdwpCXJV/4XRBHebYCPQtT+2JFvmCRotTx/o1RPsC1tFYQ6eAaXySKZ
wUGyb6uv3pCE6soQQ3RMWvUYi3TAeiSo2nEusHbKskURCCqLqa2eDw0j/ClGIiJCeJmpudtw54PV
uEOjqVWUdSLxFzZE7RHv7lC1CDFef6d7hBxEu/YLvnXQZM8yoD2V9Xu+C6OjCjd9vg/2m6ntXBZ5
OcDlPHlQ5T0N8MYvtzbF8kZV+eVh5KHdd6TAQzvjp1BA6L5jHKo0Rzzy4C73ibh0p2noNJxKUW9X
h4PCtf/77wMbK+rJwc1eCwdVIRekVL7sg9ltBgpilZ48Y0d+B3BvENJ3MF5BflEJ//jdp34J0jX+
otsydULA6qDEMqvF8JAlfUpEHy/LxGfhLAL91ibRhE0+N0iKXDdJp4RzuYrgrI8WfUFXbNTIOOMz
HToCE764S3+quGm8gVhf+ZE3br+LbLCtno94DqTyr03khFluWGOTT8UEbKsS5hLRiVOaoQCrx4ik
Iep/StUVQQDIDY2k3qujIg1bcGAH9XK9ziJatZV/+bQ0VUCS30QUUtLL+aNN1NRq95YzJIHWtW2v
hL80RCiOH0bFLA47yh58v1llMJJ5lIr3lZNBE0RrLxI85MCmsaknRQuI5qC44sf3nnT7KeKzcxE9
Ru1t85jf0+DJQ2YrJrvY6tkBsKTjgKVX/WGt0ZLvFFfpcV+761BAp1NhwKLGeGvyKDI7MWnj+W0A
46I5x68oMA3uYhHcvMcaoYL5LzyawyHlGot9rn9Zf9RHwXBxB33CmfLYKSUrwJebQ3TzRbGG6bBi
MId/QMilL4kGyM9r7cblmMTWQZ8gDUwy88uuntGHelzek2T1agO09Qmvy7Z+vs0Q5O8SobUr4CTE
XTj/J7VFHYnAbfNONMkUmkGclZRBjDe3wOfskLsaPBYYmQf4tt8OInz3MN3PzNpvnhfWfeM8trHJ
gkmdho3Mc9agWJWPYMR9Kdfwsu2j9eaPPITCzZY5CE0HY5cFU4EusVw1PavNLX7y7VMpE7qiPtce
CdSvtRRFX7vpkLsHRGrHnnnVDRkbgdr1oajFGxwLwUyESD0lq4yt8GWycZ3JEwbpAO00S+409KNb
Jrkziy2vl8Zta7Jz45Yd2nvZvtCNjib/xqg2yN5XXvX9qXej33IahoknMlrPxHHOTIpMaMP8YZ9o
2bRRXvSvRtwywTQqtLOtLxfsuL9FujtKLIags3CP43A7k3rU6NBQXtsgbd+yHmilkLhvwQPeWakF
1oK+yNU6A7NGIywo6QDuZ6q93BtbX3jGw788a4y6rnK+pdEJYLqauE8ZLpbqXE7UL449T3kloYHa
jjTBu5dWEjl22MkpqRL0ltkV9uuamJZWGKZwcTgghAD1wI3gjh/6AhC6bjzc/3XCQksvIIXzRJSk
XUcmAWSIwHslLPDe/fuZxNBpjkyOCJUj8vrvtoEGiMrnUCKm8j30PKL5BgtWsUHG/AqpY3mqJeV1
O4BbCia9RwaXjU+MEoa9Uomgi+WK+VPfLnubeBeqCnvR8bHaRaWmFl2xY3Q33yrBKbsGik/LWhIa
AMQTOlRIV9+hH4N/YfpDlhzEmsrFUJGoIf++edzqaR3Qp2WW+1adDoWEwEnUbFEvezguaa1eB2gY
CT707CRO5e+K38mUuRnvD+NerxkHElaaPITUi9IGJeI5pz+8rre2Abi1D7fVn8PTfPzFh/4FsYjm
luPmgpqp0pfLhYVEY1vk7uMLgKKgspHCAIHgd5ni0sxo5YqyoytWz+ShoGDZ0OJXMQcYoI+QdMO9
M3Qm5tztV7F15VW0zwnLjVmKTDck/L1XSwNdZzmVixpeEkMYHPifx4IUWCJpGeDaiOZ/nemp0pjh
BvRE3HqyKz5X0e7a9qwv3qMjeWCPd8cidPyj3em3HnagCQYJBNQ2kuyMWVeeElZ4Yp/akzDzJcPG
HGGYo8hbh2AOmVqPbnLVbqFvz/RihkL1KvQqNPzeRIzzn6V5/O5Dgd7p/LEffhfSDiASVrBDd1q+
EB4FPataHxC/8QxMNlEgIVUiXRtlUG27PiksDnoCXiTn9P3MZp5BZgRSt9ZgvEXBhz3Pi8zcl3Ew
gv/C9IsQJikZD6rk3xCoIkbiFhasN+465P/lZXfjAruMDiJrdwXdBWRGlkfXoG4YPxf5MNg+UIO+
F6KNFjGrtga2Bo2De4sTJhl+qfKLQMB3iq4RgfVr1Y/aA5ThPnIeMrH+c9y0yraKDb/kDBGMXsaA
6Nx5DQYVLVLbJF+m8FjDVNYpKYMgqgAtrBJfnQkzJa3p13L/0Pb7f+Sm90bqWGl02y4/VTqsIPN5
RBa/iz8DP/YeR1l7pMMB6U1MrCZwP/nFk/rTL+uXEp6Y64GcREfUZeu6Aaj4Fi5uEpGzG0PaYlvK
ZcnXrsFunjflUd9txIAQi3UeciBIW28d9HVvFoofKfQGImCHUohC6zaifwGFfqlTj2B+CZytnnNx
I0n0RlGJ1JhSLCh9NJrnC3xd0CJa+l5zhbG2/BbNOvZEEpX7HSPIKb07bXgiiY5ZiVuEqfr84eYB
NnSP5yObj4RO9UTmxq4Kc78n3deU7Rv4e8CSkLKlMpKP7TBw3WDmgqYlfIRAH7W8Bm6Kk0wJfzw4
0+ri0+Vw2k0hkTOS7OWBawqX3ibZVLy0rDhXEtq+6HgixWu9KAI8h+mvn+I8fc3WP8px9eC6RC/u
VwQm9DrRjgHaXJ+Kkz0kmS7J3DTRZlAxh7PRvbZTlJnjh/MmuZffWqXn0EB5Z7Pv7KTJRe24DMbR
DSaxfrY3wnzzKh2II6q3VtvfBK16FnHEyXKAx93Gh6eQ7sZ5sJq94bE0wiFZLaD+jHn81Oc00NKy
iszt4VxuvLLyA909fr7+WaaoTne/2lwTsOKMEZ4A7YDdvLbanaGuIji5AF/lRQVxIOxSXiBgWFyd
p6DJPTFAGGxIsrSMPA7y7+yqKGmcleR0D/NTYDy2LslWqvuIkxketu4BdpEFipvkT1K+00y34UAn
ZtXS6lOaYTw+XJdRUGPD1pFTeWB+34qURfTiwSkueX7KrWceSPZoO8FBtixeEi2E1vChqLn+dsa5
94IVa+J8YRLA5BXcrXXqmGwH+nR9OJXsisMANzxUD/Y+0bKA1s0O/w9LJ3RmCkEREyb2KFh6BXsq
e0+9p5wJXqsPZpvUo80m//6WsrMlAbhpKatZ+yvVgZRjHJdewGbSPffaMiEAbxa4eKEdrsENqmyq
gkIhDH8EKo/kKNRVEM1CtYNfLIzYhQHCnMGUunHfL1U1eLP3c5+zA9bwux2ML2MA75DyVtYtebe1
3mWxzorio36BO63G3achDEp4+2SeHpCW/CX0voc+Z5QCgeW9ljLfQyL6qQn6uCbxL8jJbGSPO0qw
sGLn3bVUAl13y236IqTMFbmDss/qcjdPlAiMoVvCTFwv1Pk6qv62kr95W35Kh9aUGjNuMReK2fC/
CNCYe+Tux8a22uBJOsAzsdZ2sMeOHZYpTxDqafuO6z3e8oLrqY42zMxwCzd3Rp6bqzfZJVfMUwUF
lZiso0gmjBkNnF3WT6AEaVk1DezmAVGtImOtr9ehDjZ9Iore8DzjOttuAuDGaaVLQnNgpp6RSGXl
XTEXgYMIgjylpSrJqgxb9Zf/cayKVce7+3sN0P5Z4dl860TShnq0jra2o/vwjuss2d+jFw2UcHiq
w7OS1UpKurZsUyBypXKMaMFDk3rgb8MN44Sq508erggXZFvb/pRmY6y0aqHWwEW/XaII/R0X579L
Alpfxr3MPt78yRusyW12uBm17vhSnTePcukzdF9LlB0pAi6XOvQesoRcB7OphTVGVanKf4rQMFy+
sYP/fXDfF11zBlLmuKfExQOPe7OnuOZyvLamuO4BH53/nmPXPz02ZpeEudYyej4uACoNW5F8r3rW
jh8DyP0HGcxFybxTdQrqceJhYP+oFUS5MDJWiWznm545vKXvuhmH4mcl6oVQwyo5NQoxmOJLeWoo
YYixaxicYunYBKTBnqCRVBrqoloqnwK+IAyxfMLX98necxEYBudfhjni62T3SETfI6AyuCqU8U/U
p/L7Up3NLHmXra6C7tQwLhbRNm3I6OVhxdnVxe7B0bFCnsWd8iP4JmAjLYmtA6/UHNDFOYkCvKce
M0+wjqZtS1+kUFv8aOMuWTQMHfB8Rm0U/v/Ac26iAfvOCKzb1SwgQ8AuuhCkscLKW6fIF2fMMwLt
K+NMsTimPANhIl/ZuQnrB6mW6aiGyegLmgJtFQnJFM5GCjEfdsOePgRFHSNxastmk5fm/NTSGu4k
8reSTYh5ymy37nxYCDyAPDzZdGT8WEC2wcgP5LPUJ5RSfWKrmV2BukWToDmLkwvN8SsRXj1oYxhT
/bKH/ScOPwdj7hxfVp+LTBN0h7BQBVBBNMlKn03wvtzpYJNYy4s/m+3wS2ysgtXph7938U1kVr6w
EtZquMdSowpxWJGwokUQff/47gmTqAhwXomITH687giHyziOmIelGA/a4xyBS8417WVlatbwRUuM
TT6F2ScQ4PO8Izu3Q+jkJEEchimarRsaI3BV78Xlvo51XJ8DXNHDK42c9it0fk41AUEHbS11IZK2
p3mWaYJgVBKLo0sz//PxCm41ResxW8RPftUgSiUv3HQh+/eWmMwBYMB9NSJUyFNyGIWZOimwu4kB
FLLsBTphNfuCOvbmuptaOqVc0J5dZeZqHjXc79VlIYqWStqb/Oeld+vLZQydsH8yLF9Js4mHMdbI
4tHZ0iLB4fYOGFoHTliRIUDnxmfTmwUQwo0oUlUZtsnX1UtVG9HbWiU1SPWiXmBX8Mx3wPfRnIu4
eo/XHasm5nryUwVGzzGtZoMFR4Q/LZxJnTc7Lqgc3pM/EPIZOQTVh09QFzJYQV7o4M4Q+WfVeHeX
yRhFWI+BxQdHZA0iL1rOSE8/H77ArD3uHVkU1LU67kEHtW04f290nZFt6iYsWFWBUyP3v0CZNMHr
kq3RhQCqe37HMutcg3Z6jE3TOvaWJKr7OLQ2vo7J8nz8FPfnXOuSCXQJuZDNihrLyDfWOy6m5QgX
bJ04Yski3FLGC06w3FP2h10o6l8iDbqOn5qTESFz6j+Cy9jImuekkZSV1UCmbeAdjKJ4CbYre6Iv
/CWiu0qctAWFvC59D+v54gi+RN1vE7/LGdWY2arXXDJHO2qtojv6gvJh/uJ/KdyN9MsO+3pS58wf
fHO2NFj5oRNqoZMvvKgChapu4WifSUpYfQbPjjA6zLUiQMhwpZK6QOO9TUh8eIWR8Dp9BQr8l1vs
asIDhGzahX2C/b3UgW5NLo6gFvpUlf27AcrKgM5zGzgeSxCLx5wXCmhCGQdWVBsvuEig85UPMRXo
Rf5v4PpjafORaxs4fyRnjKjqLX0ZNElDjBWn0Tv+lXuMYOeXSRYcRlNxlQeFHXkfA1cYXRO8NfR6
PUrL9r/bavjeC9sPvh6cMvd7DUrENH3x5UR2yvTNR+pFSjCxAcNVHJ7YALNVwonEkXPOSPKohbiW
ZkXmtSPk/kW7R+eslDtoh2spUQA8U24bVzmmhj1zTAwAhSJbtLmRGOhhUjzHbTca9sCdupmzxJ8J
d8LFpJPfrwCGSUE1TJeZJmgkLdIC10tT8WvPMwXKzQcGktNcXLGBitKhdrsSW9A3U7Y/5Aj4Rl3G
a11kS8WqI4LPybhE4p6lnGX56ekauuuwLynVl7kTw7j5KZbq8sGF0dHUw5zbdA+tT0YqVbJMVgj6
aZ8PCKiKdFPzJGBpfMgtaRAvk+fCUjM9DtqB/8Ylc1rQ7V4ae3HB6RYTRaxIvKE6s8rxJSrfK5kv
BMe3WqgwqAp0q/ZvcJBOn1K0W8QScyFdJzgXubuTM0GoMrbnmX4jwJuS29nJ+ub56fon5pJgzPR3
lwKMOxatPYNI/p3GHGxRHX6/QlDtaSliVfKtD/DU2NZwYePGkqHIAFWDI0//Cks4n7A1hmAGKOKK
JCExe69t/4qnwBgDuGKlh2ZA8jmBBBp+m8uT2h74aSN3SD5OpqZq/Yopqf/ZHbtzMEjINfV19ZGM
+kjttoXb1N2cPZp3JIGUq+CSc9nfqxtuigEprEFOpe78rccfwplBrhIsQWt5DTVSrLl4u1x1IC5O
Tn7fxBGu4aEYdNmLLPoRqIixhm0u4/B78ruQZWMDco/bM+5f18Fq09dYUKAM6lx3RTWXDVOKEPgW
7w7FyZDK0yZEW8mGu+0h+bipNFOhQ/kz7ZIOl2+RkEYwjHrQnuIGSRzJhK6TSDwT2/1TrtsF7EZP
umxtnzyfHiyT3l3rqP5Ypk4AuGSG4sNsO76vUZdm+GMIn8POvq1L2qBRf80MTldMaeN7eAdBHEP7
3/DchJ7x4D0o0/nwlg/P0/H33H3/S5XjTEc+u6HT3Qly/1VaSghjmCFts95wkcRB5v/IOz/5g/EJ
sgxxOLUFDEbxRNfphV7+1QJFit5x6zLrazu4t+SLv0fuTqgOsOBnfQGS18teXkdRGk5HMbFFhIS7
4ScaNAHGOMSZn12kBSRXCIEv3Yy9gz9VlGh1SVR7cDp4viuDWonYED8QTzjDCRzr+YJEl5dLPhgV
t0rVg2AfYEgwGwP/VQILe1ecOOCkxzMdI6+98g4qzhXndJdsE65SSp3gYAlnsmVR0gZNkI/G2DXI
5NxKwjX0IYkEPSevU1rmKSy2zSeaLdFZrTv1kdZb0f9X1OeBLrI657HcnJzZUGS/4o6L2p4ZN0YR
GcNC+L7CrUEfRm6/EwjofFLXFtfamaH3m/Ls+aHtlk/FMm0WDTzSgNT0Ivua1GFKLkiX+ZDZUG84
VTfdM2aP5MCD7RGv7j2LQL7FLQhAOzASz1DkeT9cFC+F4QdqI7bnBqpAE8Bt7P4C+WvnjuqHfGwd
wT6JYpKV227UYLFDGNNft8T7qVG4KdexlXsn6qu9fk3ZoUHgvnyTMBTJRI0Stbs4uNQC5xI+PovD
z8KF+XELnx6U4XpmbVQ/FF2j2nR8Pm9mMrQ1PyfJZfpQzwVN8ojetbLwZ/O4nYRoxYN24CxtArmu
rxdDpo7Oq07g8FjJklb3Mv1vqaV8mnL97eHAOXmJIrZOmMke3vjCSzStu7GLpI5CUZS0jLtFhsxe
lYqKfuV+FDMtB9PAxtyAvjuaD987oaJWEMcfcRAsgFiPcjZ5jhG1VozdA+uQSEOEs4rPzZOsZydf
YHtpdOY4v1bR9un0O3NWjBWAyQYJA9kpW+WJRnmq9KmjfKciJx6hJd1N6eJRzuhour3strDWXdFi
UjZcn+FCOZXyqVEqmiYWs/srrdpKFig42W+g63Nz2AYnj7HnmlXdVfub/Ysc1beZs7Lq8SVebcx4
ezleGbkYhDj36u8mEgPKea3ch+fNmw3d0s+XR76z9f3BJx2txjboc1EXM5rnOlJmdmXuYTaeDTig
ZJkha15yGD241b04eYSpySRwW50at/1iNFDlf2NaIL680zC1R8i39z3sK17Av/TI0YumLJ9Zfjxi
94/PIzAPTulOl8PL9kT8EbTFMw6t7+wwkMmYvijbPVqb4jMBSaB9AnwYDw7aFHXZ0fHIRytVRMAb
rSlAbuxg3666UjZJk0c/+y0xh44DCSAOk5L9TOp+qeYU061+Tzjff9sYR51OmyyZdoSfgmZnjR6R
2bk3TssgTEX6vJVAwrmIwpZkhRex6DXBzACvNyI/PBHiQSEioZ+OEFhNpSKBUGN7UHD+DpsOpURv
e1PwB0JnYNj14i1MFH2jQKeN0oe/2NvvYRU+7qoczvcZGO63CzgnWgRLXl88kdyRHQ4tNuwDYGYp
0d2c/Oyp1cPGdD+VFB8k69e1bAYxaALVfGA9mbqdDN3HgF2yZC0Y0OxdxPdqv89noqCJGER+F9oL
ceWj9twBy/5Fjv2NTf9rjjZPuNvSDjtZvuXPJWYWjN6htIfJL2/2SzUK+AgfcqsmYEXb0o2dv3EG
2EQSZmkHpNxd1XOPIhTV5JsuSuIWQKgGXi05G+Q/k9hIgkTYlfsF8RkwsdjV/4Cj3QgLpo2PlG4o
aYS9Rt9mKEDTc6olDNrtyXP5KSUdmZeSG8IqtSSzJjYpr2RHSBA38VghCrx88bx+rzPTTKVGEWOz
JChmZ0keko60GcFwU6mExqifI6gyvSJPTYxJK+Z9YJ7P/pqrQO0VCDjTGVy7/wMukzY9aHA6WlDD
/dFuQX3/mXDURID9HXnvxuz4t1s2dByQb4pIuTQ5DN4K0gcmDLa6eImm6aCeAGcwbW3ZB/s9L/60
M5dHz8tVRb9H5gorqlLii6Pplk2czuOGOQGxi95Xbd7hcpeFPqMKKXO5qWmo5CkFecYtHSdpZDjt
N+xFc7UZsJNrnqxc/GhzFekrfItEOqHU8Ok/zSE82oqT22j4svf8ocUSJML9JFLZE48yeIOcKTXT
+kk0Fc1L6mLbFIJ5WcCqYUdbtd5p+z17uU/di+JDLPduLU1CUswk13kE2tBaQUAakE5q5xj9bwDG
th1rtDkayEHuy567wt8yCAtX0TtjrjW9vuEupnczUZqT221DN/hspyXfJhQS1X1NBChLT3GtFdIE
dv6QVZfEry/XBpTlBLXbmtE9e935b7T8Yeth6kAF3BAK9sW26bANRUb17Wtc5fMAPMPySM/rRLRB
LrJpHSqmxFG3vi6G++5w+9fOmfWvkTddiIpMgJa0lgkh/iTsADbS33x3by/sp/uyWmF00m0cKijz
WkYIKXqWwQvkK/DbeJv+ZLJQgKSYjOQn0tjccncwqFjiO+EbCgXNnZgL0vDmit8rSkmzKreyhtCL
pubt6xsbMi6phEYF7RhIyVut2nEe3EP6wxu1GmFnpvJdF+FLJZsppCgNiTBPnBDpKxIQ+6FR13a8
MdSQv98cAJVNitUjZPEBPg7+vrjK0xu0ccos4OiylO5M7ycxFm567i57tt7UWMvJkBdth0zoOdr8
mFN+w839zBGVL1PrQ0Y0s1BrGlaTaJbvzCrAR/VVCPhijGJ1sai3bS41z/GeJN+oepw+q2DLrKsa
YeQ3O9uZZ8wid+WM62lVuFG4SvMxPgGlCKyOfN07XZLEAfp40D0w09q66uF821CT0JPoBIGdPfNJ
3oF5M7IDUPgU7j8UyfpLSxEBY0QkkO9NmwEPO8l7aSSs4lmIpwMR7tYq0rVnV9KhHllUSDENaQR+
FsQXrwezbmvzPMvh3maFL2ER3b5ahLbcGFoVtr7jjuD6rF+wREC8JxdiBAxt0SuDABcqPHBUi3Rs
8w8oCtsTjeQa9Rb47RWUkSzlcPy4PBnGz/K66X62ylC/By70f36e2J5IJWCFPiNtgH8ALFspp0G8
hQvP/GJdz6RyysCdqH9DaNLOkuK/dTrM+ZsEfRxkWF4VLgqOOAx8dzzHcRhq1Xg4rAYDNefhaHsL
4vYpsGc17CvGxdgLHJ4V46xxTgRukz91+CALUrtubkEZJwbPzdiAUMQc3Vq+411ZmhEE4TpeN80S
j9scLD8DUUB6WAs2DZMghgCg0j7IFhNTKMYVtASN3/AlzbclNnTCI6ZGhRp1zbFaBDFssu+0Ne8B
WzrlFdd8C1SZ4lXwpgm3oh7RtWT1xVBWOlQjH2AMMmqPFX+VX5XRrVC8aPM9awdEM8Ik0kexHHE6
QaNQFWH9LsUQUC20I30+g8CICQ6nyhWCEoRohNz5Du5vYxheXr9eDjawtYZwCGz0R0ZTh36UqopW
H0Bdr5wSznGjKmk3pGHqUHfyoaJ3/aSILLzGwbmADJyrEJJ12V6u/IYfrhmdza2eg+Glwk6OMsro
5wLr5BSszhWkKHyhAwJSmvXk0XagCPP38YipG22VTjwSNRY6WfGiHfkHk69kDUZQh21jS2d1oBfY
SbqOMwLpbWEPG1t0jl7FGCUmkD4wddSufr0RXAcF4DExgXvX/o4B0fGfSFxM+w0CoouI+vXQzmo7
FsnhZ9ZB96jk2pVmBLi9kPE7bjMmaVVN4mH1sgGO6ayw1cZgouIV3IC0pS5HQAN+iPeMjjf+Ujl/
h5OXPL4+y0HibTGRYRhqkcjVfncqII5Jj2/tWoRsKFr9RKae0rLsOpgNtxPFgNXfU8Sqz9mufwur
L2W8r2i0FDN/SsIDxq1SIM0jhGxAWkpihg3bg4p0cHJwycZxDip6t50sFuWp9F7e8ejguX847WL8
Y88+iwWN5/YGi89qYNIy2/PKLMSlwScnZ7tVwxKs4Z1IOWuqX3h7NOD1RdvMfWfpURNJsHRRGc51
qnMU/J+282ObkkWy4g7xYh1Es7hwtAsKinIhBsgEoBUIx+8c1WjWv4BioBKaz66I4eA3DqVgJRwv
GRmwl7HS99NVSAnKbQW/NMX0A2STN4HzQBK1cwXHhaXekYptIFhElWXk/9lUmx66XPMsFG0SaoYX
GtXjSpP83HVX2JXDHHXf+vaIEpcJmhCXojve1CeSEkFVtld920vix3GoYNJR/gjMrfntOHimOxmq
DX02EywpDur26E/8YKfablV7emZ/cfU83D++33P6Gzdp3yo9wguVH/MK7MAEgL+3bnnueUTZOgPl
H5cMgTQ4aI14o+966vhLqHd0VehSTYWjA0Vn331OvVHH3/NQTAjlNvWnF2pIi6W3as5J335CB/ES
VeXJU5AKr0MjPx5nJLE46S2mchl3dAscD5vsFXYSQ/sqU5Yc1txjkphTpZCXUNMF2RuYFg1fnSBC
62U3I9B8rIvZDMD1wkAxRsFT9UGRRsZDI2uneN7WrDD6TG/1vV7ZhZC0UDA7FQFBbZonC+YtgPdl
ZkSoTLhK3oOvPpVUuo5ep2UJvl+jSXB2vz16AqaU3e1C6aMmlLGWnH4bWj4yOE9K9Rplxgs+9fhw
XJn+rmizDk5SMm4wmZm2mPC0mUA/X+TMWrGSAR9oFNTeM94J9lAB/YdrHuJuw+uWLsTORa5NuDSY
ndKAUjVWMjaQ2de93bqG3Ox+iI5JaoLYFeStqeNfqx+OhgnV6R7BLnQwBwv7pGkrBhybfOc6b7KF
MNaTSQJ9RIt7YoaSDimpS31LcVd1bZy5WEtCpAclepMT9xKas3JydKSP4WxqIzT4lBqFlFMYixoi
9ZL5TVFk3k0O6P3K43c+KbPVpyaujfSM+/gaIWw0DfyCo7QK2Fnd8rt67t/hHO9jsYFnigfUb5j+
1G6Otuf8Aj5twMirgqdrF4N5i3mFrnJUmdW8H4/v1+jO6zx37nMmmOuaa14sS07LSyLu3cmu7w/C
FCkTK485BwEfmjGU3dOgG/LEcbU9GdPLXFNQVet1LOPwVbDzqaBok/hBqXMcxC31Vq9fI7L+JSvv
c5Bg9c3bJMOL6IxeC9s5LCdvp94NztP46wPvOU3jFF6A9yKo/PejM0oqNLw49J6yPK3YR1BdAiaT
Azo2gzRaSGbMEloVDEtcX3pg5qgEzfmbKEUWdZUpEbuMemf5VZ3yxjae0CumYVy9SqNxNix4LTg7
Of0mCZ/eC/tlKIJ987JTk7KD4yFzUYmDR0LNgAkeqUtpIURvjKZTVOMZSpQ/ldVgBp/QZAVLMwAn
r9Xdsqq+GUzloR/MmuIVod2SjtH4K8F24/Nbnj+e1Mk4czOS9oClv+sd4lbr+esaLkhnb9YN5hqT
/wIh87MguFSshuZ/TsXJonqv0zje4XJxiQE1Cs//ip5pH/vDYFH0sTr7C5mizIMBm9a+qiBF+w0l
YGAgbDanet5F4h250hzMcN62WKUX9lmhZ5PNRAOpXaVOmzsE5axpuPYAd2I5TmHt9EljVY1D/+Sb
3Jd26+ePeAi+xIMEBioSNzekzwCpiIc7JoDVKzuJPZ3ccLAnwvdpneR1nYgZHXfPrzKMuOq64fxg
M72IhI0PLLIuB4JNyICcQUuVSfAqGp07f/85NqDfGWuFPtola5bST0Pki8E4tu1/ARMbDlerISoh
txEdmbP+LzeKGU4EuwZAd3ZDPL2CFZNfLQQGHQ/kJc7PMB4gQJJBnBSts1qyzzFcjvM/SfR2N2T6
4Q5JCefDtfoF4FBVWKev7Ob9uNrVc+SoYZokaJHB4g4XUQd2ICXlm5u2dj8p5GBEIdAQ5FGyeScY
SnYtrQfGiKJELzdMEuT3yPhacQOfYeNmx4A5qqERHLQ7TRK55s1TB7hcmognU74MkkEKo5Jasj/E
jYpTMVIXIHNKNfnyhMfJwap2sZtk+x5IWIBK80kn8RFFFAX3/PfPFb3Q78g5glxSqLRBJVbPxeNM
N1ZJgKJxrzV+4VI0Vt2K85fmqZMV3WzS14Y67HgafCl8khFh5fFNh1gti+FpYU4/IOxx+NgF/TsM
Y8erY0e8Y//ZhTiunxRhwbutsZl578eysPnfmNbg8Bc8KXhO9sBzqOY88JJ8bCUBNJsU1vXWj/Sp
UaqRjR59viVmzPmnXHO+B6vc4Sb2DwannAu8ZO+ekFbL8FTVNAFtT22DgkCSiM9oy/7+47jVGUG7
tjGX/U2ZoFUOVu+ZFGKc6QvLWeyoOzBKL+swseoqM7D69jiMOi7rs11uljsOqAP/3qjuKktJIlUX
xAIwzlI6ODFuVaQb30w7pAwCgl4xmzl+zfGPMkYrfB6fpl16tWpRYaVbYm1AGgYei4CjOXPWEn8f
IDPdVGZCUDVbyrY03W43EBI5OesTsjBpopO2Q1K1TppqZxwfB5hmlabZW1Krc5CpcdOoAZRarGGg
aC4AYCgewRgyEk+iexUUFtM88dQNi3W7Fj9umoVxgNC/qV8Y1WqVFsomwWhQRZEraDFxAkIldp9J
ks51chOr8AyAbBknf91cwaZvC6wXgPJECY0gtPGbT3t+bTakYIlgvzthepwj/Mszp4Hi96gQZojJ
/t9TbaEpxuYm7RqAw+qZdf1u5Pi2l5HNYVWKULADX6hL3DUhjMU8JNILYKglO+er3yBdkdDJht8G
mM/RG29cRVWhr3iwrZdQ1w59Xwl1ulVEtMmrX99Ysjq1MXNhc2ol3pNg8HazeKTaduL+z0Pc40td
/aFCCKJnwZUDKB1jPNT5lrJ9Jntku7nhAKoAKxsZT464DlV5O/IyWGt9GKdPpEsLayO1GK7MGw3X
PB48OH/LZOPLE8u+g2WMIHwkefPEFjjSScB7XozWe5A4hNn0f7FMWmeLsCPBO9au7TOpvexAdMzc
grVxdpU+xPtOp6Zi03mSFFqb1cY0ecggLr5aSmAaYlCv17iRmoeNSRJ1wpSFxKpRlKmegOob0kwE
HK04xSMFMxh9unD4pOet9LprgPCOtKhC/Zs+w6z3K4bctwCEnMiGmOaxXW5xS+BsxSu+Y9l9mkp0
vkI40BgzfTX2LUi47+2OQuVVtIHl1buYVyFpoc/yyEsZlKgriOuBE7ed0NsJvmgzL4flo4Xm4dSh
Lt5frxyDqQLVDz3ZAO8dLFFMlEUGMNQgsa0i8eXPTW4TdLA/OzSNqpi5umD0XBOejaBhnI+RyEW6
1oZDxYjZxX9AdC9754hPOJlfkVlnVSsemZVFA3wxhR1PLc2Bm14Nu/Hb9E2glSbobUw25/xoLjMZ
MS5NYofZdfOejfknwbCi48GZi2VKHBur4jVqxgqz+7k7MrXFi/RGJm99IKtgEx/0UClu7pbjhFpn
S9i8Of0KFI2IHIKMYZ9IuJDoM4FJEp2+gRCKFP+JF0bIpOwNjUWCvGqiuZwjnJF2umCcPGWtgcGx
MnPmobXG/DIMWr13K0irR1V82v5c9MtpKldYBte7mma69RnM2yhcja4CYxzqc0ITs57cmJPl4JQh
CStqjtYr/ob3vkVWurMe782QWFiTT7ls67rq7cT8qY+SsjbdjZ1R9BZpbQ+d3qiaudCEAMdgGZxy
jMvYBsyasEy+vaXiCGD/K7P1sh7YW5jKeYmc0+LlNKfLxFN1Jh00MbjuWx3KIa8HdTViPhj+ao6a
2I5POPaAFepUTuLa27MBDgyxLPyaTC3qzUpnlc0cgEhEymD2WvAeeuTWfbAF7c+q15gqdZxxnfdE
3whijxJQ1hiBecoCB8NK0QIV4HxroUIPrEqKca9f5wILvqB/ids4ADAgP3WaPI149xnpBhCFhtf5
ixkalUc2c00MHywPU2Cg7Cxu74wv8F297t50L0QsmZZsf5z9gw29cDGfVbxPLCN9/4jG+YtqlBn6
89KZUDc2ghADJ0cm3ZU9IMG+LCMnFtu91mjlnHGP7Xbr1oouQWZOvQpoXP1mP4ibCJrtY0aTsCPq
WOE0fabKBwmOutfiVeQvwGDb9ceVMTeflFmGaYixz2xMiHc3rtuw3OezC052AmQEd62kpszL+f6k
Ow3SeRcw5C0exjb2T2wE3k1jhnNDOqQf46vsClfIBzCS8gXQHQTzYIDpIk4ID+dClZcmV+QhtG89
lRIdCqIjXzWM5d0KtqjX47hsXqm8wNjMWh3MrZ/K/ltLYH52fXIZbU8/7LxbVCnP7An/3nczSgNu
mXrk2PmZaAoQ0a/YopWFpLT7xYZzfC+oxasAaU3nUuD1zdaa0AjpQa1N1XbkQTFlOom0RnctJCXB
L5HhFWQ1CbtpVOqyeQvgbDIc8lHVyEf6KBOewv5qbg3Dc4QgI7A+LefSRPJGBJpjKZZea5cH/8GS
OvLKrtc+8yHvpYJ3KzmkGvl2fbvK1c4VsO8UVoQWpJM7oH1J4FJXZWQnMcKGBTlyLhwch/QesnKz
ex4wHfdNsnAjyqQ7tlEOrMJtLmYwzyDpDIs9dKp/6AFY/h1ZtZ50xF5REylALzt81n5H/2BW8ZOP
+5d0ecdvItf2LPTmt4BkRqYdTr4h2DmMfoN7lDPGFufsm+H4rAJLcwid+NfjkqHbkpcWWxd0P5Cz
4sO3v2gSNz+bW/+o4EDNgPqTiggTIAW2LcOQkOUb3hC9rh/5THdsARnXotSMOjgG7UsEOsZEonf+
diLC6TQXjUr7ow/rPV6FjSjAtCOhFA3In4my2KkEhJS1r+xkEBX7cHyl1hlSh1z0d0C1juy8zbKI
PG63CexW5xfCYWCS7+Pngokb318gC8/ejcP4JEZ3keaF7HzWq5Yf2hmC26z9W7ow2JENIeHLGGEN
gHBBO1+UDRz/QxeiBM9kagkeNGzNq5HrNp5iCr07mg/rVV4PJGbWU1W5kUvQcG89o1T5epX0WUky
W/3dg5VgARtEi7svKOh6IQCFqqiOEjacpXnFGshLToJ+UcQ6IooR8ilzLnPvaMORiC/YXZJWXKSv
cuUiCP3gfAyFNi59EOpcsJ53UToAi5brBoVCU5JCaohkqlratyIr70hpwG8a0bdbYABVnELIJGu5
hzRksy9VSjLhjc8NLtmiBuOoF5j9cD3pOPQ6TdR00+XfJShEEEdjWJGynURhOLDhpyz+ZhHX00r6
2Gu5j+0UyvCLd7MZpuKP8XR7K0vanGA0R/zAWT3UpWfB03Yq5WCCfYfaeT7DDgz105BtqcEZdXdk
K9townkHfW8OxHWB2Tt+Hzuem3PMYqHNK4dqv/ewotfOORUXoptSnzFaIl66BNV6deIy7oqonqXW
Gtx0msCjyvU/uJeNuiblSaD8UEtBtCZ3Q6z+hyBQrmHFgM6DNIBQ++h33XeUeK0N2CY6d72FNMvu
4qOBcPyDfR4HDPRpEjSL8f6tat9pYtIP+uHrsNN/n1KE43vH4yQRPdrAKUTZy88zIiH+FeeuGUGK
xWbfov7tf4HuiM6LALWyuRAO+8KZl17zMI4RVPTX1rbDaF2YqW6A1jdnST4ITxttis2TVn66faFM
P2JiuUW7q756yNDw4eO2xhFdLYHbz8u3eIUJf9ud0QpxcPNBDoqvQ1ndq8SB9rDiRtu4ERWbTVUD
FKVgc/eLBd4nySvGgHte2EOtzlxQizZ4ylrQRFQ+wECsRDY4+LesR1hzKzYBWOLdhKVtcWbMc4EG
fSJMpwB7V+N5mStpjsjnGX+xJtuTcbe1jw6y69rjjkTCnDuC77z+4aecIN3Wqxly9tjN3hBl6wQz
nuaVwo/XXJCNPNxQT5TGOFuCO1ji1IrS863W69ddj7Lm9A7p4UmkPmmL51nNWg/IvCKuf8DZt2Z0
tcGNCG/QBO96ZgKQoNA39hR88akujKMa0/s8hoIBRNMpbP2x4ubRImbmwWQ14h51da7hpHT9cSSz
Tew3deIY69mnU1x2p/FPAhZxYX0dY878922A59ZxqMsLQh5p9OyWglCOXx4xcuhT1T6FKu3z6uPE
UF57Z11zwtqeGFYRW1d56UA3oLT1MH4wBlpnznfBZd0VsgTmDv/Sbl5tDLguYLp1lxmNg+yqA/Bh
jiqM+SQeykiLsMmitt9Kzk6ywFtEqnBr3hkJ25GaXUvHvKRMozJXRZgv+kS7Pjw9/BLFCagZc9tj
F1RlQihtjoryucQTjOdDXXljB0Ruj4finqhfQ8VTYsWbP2dhySFDD7NeqGg0yqH9TUchpzWwNRzM
9jfWQDSjJq71fvaDOJvZ69kTlFx0jy0I0yOAuZQgN1AKGRw5Gj0/KNSbyZYEDqVl0Ech1QC4fglp
TqEJALO8AsHpex000I7DZIfsZtP2chOdhIAteBZqNpVgyXSZjD+W98H7YvR/uy3JJjBCX0qDwyW0
4O+gGP1xukgz+ZMQKNiFexMvsk1diQmWwGPO3Layqry7uxIjNVt73MsV6bY+hbGzEhH5L64BLqHv
kCCsEYWWtEFqyawQbudlIAIYm92UQI5xqulRZGpE87WxnzcZMmFVtV2AIg3SNguYK1N2UXpkAnoY
/6kvpKVa1ijDLiPuopADPf7OH6tVMb4Ufdp++uH2h+Ms13wVJNLNZ0Ezrsd38pTufQ67feBuMnp9
pmT0SCBwVfBuDg8g3ImYRmBsKhTmz99yFgHhCJXT9BiA3rNWhV5tjXKdkqdPZ/l0TIE3SLPfnj8P
DKGvPUQmwczzCfG1Hhlqh5hAcfPQg3qT8ke3ryE5otOJ4c/UJVPob+pZGHTrYhQN+SHwzQTLHnYx
chVXsWzEMEh3LT6dS13YxJQVJ2gNnLpHEnBYhbxKFp+cZvTjfEq1fR9uOoUtESG6+1ia0SU6WbUf
97AIvMOTPx936WnSERBGDzvxreywb91rLO5OB414OzfVf+SnQKedbasxh0qLMP6QcugKi/6sfyqz
s8UpKg/vLJFqG3QfMwLMtawcbYuvLX85Dci7Zw/CZDTGugEM4Ex9YMhvnZlEaPzDmbXsodEcNcyc
HuQUkw9n8hiB6CMooRT6Ww9pCHFkpiHoEDC1kEtleVeaAImVbQGiSP6V5sDAFLtS+dHomTm2J9tY
QRNQ+GwIX8xyJkhcqVV2eobMRuHCTVwg1f5WhmxhN1/TaixgmvbdvJMhJDtzJZGBRtHkihTK2vf1
+yHAfsc9J+WH+/VB0rn3X4X6ck5um6jfg4OxcKgk9ar9dcZZCiIrZQitBnHThgovA7XeorlGkM5d
cBjojaBIJp0ROG9/Kygg6Bk2c3vYmwB3Hfin79ZbluBjOz28oOIvoHWpeW1JIrqC4XV6jx4HYwnP
7bhztfJGTQpddK5x1H3qCN+8YQwKFoGqEYutKNXT+7cZczEthB3DPppfa3MNUm34JYcHsfGvuDrP
Cm6j83VIhG0d84S4oAV8lJnRRNu3nl8XFULwydZrGO/F485Gst7syxX4zfA+EkS1ahDkGRGW9bRp
avfyiQCoerZTHfDCgrY4CcZWl8WD2iBqVLzzxH/Q7tQ3KaFm55c9gpDTv6i1xpa7iEHSEV/8BGYh
OjQoiNZm3LAOagLTwErIbNikThQA5TRx2QzuGkJAS8n8RAV7352/jDmruOtMPTozwlKH4KHRi4M4
GqpZE6dx6Dmel0GJ9J58iWPJBLpPSiLiT4cUljz5c3cD8Fn9gLiXVA4ykaHv4W8CkRjX8VAYTrKw
2csMwF+YG/9yLxe4LUxfY56UI3hiTP7pcE8zqY6rtnX34yWZAhVKL3bWhkYF1ScwEg4Fk+SFXGcg
W2Cpcmf6fnkV5S/wAsJfbgxBXfszXwEAAEz5+vAVXFENQz/MIMKvAKNAT8AdOtB5nNyabRmQkX0S
+/k6xHYRG9eD3KS6JjnXeN9JVQwlpEGGwlGMzHm0x/BkvnX3zvRqSoHbuspenWD8aUjMpstWsRlu
mz9FQbBkVXJdw3tTE2keOQdUMkBkXHg7fhKgADmppGlP8oSKWbTYK4TWGH0TaysxLbSX+xRQHA+F
tSn9jRrmyGhVWpBH4P25LTy6AETxIO1uKm27nsKy63ZTdGV3ewmbzoz56IXkjALOQKcc3hmUq9Oy
dNoi1ONH2+h44zOJjHaUAucpQftwvpzDNoFT6mHyhit8z9p7cpvnQTJmy2tMAv2Ng4M1W4DMxRIq
FbDlMCD9u7v+GqIAfZj7eShFjMjHxtUFFmZGvb4xhRvWBu6G5xS5xMQiwSXQjWIqvRItaWfBc2AY
RsoPxvfHkDXZaIgwMc1CrC+snxMzP0uMIjnYoVu5Jjts2ak9bN8Wh619b4XFq+F1hBqUrqCUI92C
rQyP5nUhdIjp6zrnROdfLBI6IkOPl5K+f70fynWk1rwh45vcJnohVj9PuczJL+U9HR5Puxa64A+g
7NSo8xbPiW/pZMO4RSU84FoQlyuypVcxSbgUCGTiyrU825NQVRqXi7YmvBm5mb2+FsYhWO9R+UQG
9k8zzfVv8NtJlMgGkXAl8XW+/U4RKaG7Fe4lj46bwO0yFRdjjzNs9jezkE5vF9FhfthO91WDAyxh
5VTF+XdpjzYm7TbFSGrCpwzxIdDycteVeTVK9gvBYLLYWCIfRLz9eO/5z2fVDei9GKWLQCtjW5OU
gSo36TD+PRUeN6xqUQwG71og5vmXZwQOcKI4G6BsrMJWbctBGOOL7D+1RQIeqCLF2Q8XHkU1jwVL
TZImB5vPjbzdRVjpTz9EWPsrQwRhfWqG0B7xrWIapStgjnLp/oBsXdkkT596TkxSZ1xUzZVkshUD
bqdpHxUQbx9upTZG6en/X1GzdeHDqZdZUPRyPTEpMBaBmGZ+RrFnwpCU9fXrQcbyoV9hds+25tMH
1+O9lq5IY8uXw3iTCSn2VfIowoCChzOn+n0hN+aYBDouer6DakZ9+dUNMWI57YFztVqB4bVrYOlR
ue591Iqo5E3FfaxwirouhNB+PRsU8ijpZjgdT3O1w8izzCoNRNtKgV5vfvNob5kIfwHpBvTX8Hcm
J4WIKtpYiX9OdmT4hKAL0YTjwmI4SyWp3upLcvNcWLB28IWyL7IqJYJFiZq4Q59B7RG4AUmFs2+z
VV97HTpKA9HYbrJ+20cIkVygDcsXucWOB1FsRgJMzTI7Lblz6HVMZY2g9FeH4kqLTEnvQ0j8M4c3
PKpbYQJT6xLZ8/8xPPYfnoXW7sgTZXDDNaFqxkdwjOL7WxQ/0a8ikARxnXhBwAzXtupmHab9+3nk
goBDVyz50p4dJ5JlevPAVup/MCvJ5z6pdTp80N9eg3OW5X0nH91cUg9h/qTR2YaemJXDZOX9005s
q+83XVJMqyeeQfs5vGINUpVbpyhE2jz0Cl5eVWasoPXayygM858InKfY29oTKnA453rbJSSpi1U+
OXwHDDw0QxggfQzl/c5zDxItb0yuph/l65swQyiyXMOaGmBCWCtd0rdKMUhgbj77nM21T/LJgJZC
ByTQv7sUGFFcoBPMuLkBpdRbUUvmKBWkqN9zU1B2wq3I1Cf6fmsUqLx7GVHMNzW0hfMrhSK0MSnT
spWfcLkjpI7u+iIajRHD5USAgB30RwZpIbcVimIkJ9dMXNIsTvJ3AN0C8Jk2s5NShYqbOCb1OVbk
y3HlF4sOvRnc5yoAIGDE3vq6LLD+6+FR5tnn6uzhlXBHGLXnkDKb6RHjwtIINItUOe9bHjd/PPOq
8kDBdWVz/kgFIDt1T+AHEq5Nwkn7KOkLssGF8h/R7nHIut340boJ0IZ9GP3kAN5TP3yQVzNk6zo5
Si2MnOP3QCLKFHaEmYYAUwSGokSbPM1AdkNYdeMLSYsc9GVzlrftJf6kEkbB37eK4PuNfTsQIjyQ
DFfi9z7DjmZrFAgO3N/acIb+5RZiAm/EFIkPjxWu8Dis2JXm0WMoE2QIWqlFSt2L6GdPWfiZtRVp
uHg+r7v2grsbJjsB3s2DMRzmzcFxG7DNhIoYeP10j5hnKI+Th7bMlylizDmU5Fjib2qt5Y1tj+BT
67HWl+DC470iW+DMhyzG9vydjz4Yy4kXxK8M2cl73uOAPZeuIu8Z60Mf1LQGZeajUzOExpeSDl3C
ZFYvoiVbRKlUo9BL3thFLHTomx7f61SgowbgeU2KLz2sqYje1q5KRpmw8ZffMGKAy0UuY6l5atgF
K5AEv6Qzb2w9VGiDQS1pfQM1aQ8yigxoRTudcvZRkEP4fWkHJSFJ49thhjE8BmzP9ML6r8Q0JRm+
/I7ttjxCGc5Lv+znYVbqBLtOmQnQ0UJhvdIf2LXacc5iOgZ97jJQ5lBF8UBhy99pYSZO+f0y0cNq
r8fVWDSfQFazkUNvbYGTOnH9jJAUWD+iU3MeHAbTBC0mFi5/23jWqkQXqj8Ts8AGLNx+w6p9TD4x
CSbiAXA3O41TYgakaqZNVCpP4TJ4IjFlsN2fS6HwUPxOkKooA1mdHDOnfHNWC2ZvX70GJHZAYZ96
7Co6729o7LozooRvVarvNwQ24mtv1xubgZbh0stlpCVgEXKHiCHJ2SMRs2CEi5x+07Xs9NcKNj7o
dGK+OUExvduSxVw2sdhLVnCF0DJiliKvCaoDy0n/ADosSzDmQfO0O5NVXGurpWiOF8a/1FVHDiVg
n1+U1X7574+KtpV34XhqNS+l943AJpF2PzPuG/t/98VAvWyZvr/pzifJSNMATUfJctQ9Y3NJZrEj
llD9gc9azRt0Nu2wokCSjXb3mHXelw4F/r4mmRWpDklLDH8TECxePhzFwtBw90UHtHkdeph84BdH
tCydm9JHyN8MV5DgDCJFbXY7XRyhNCSw987/XGh1Z/Q5fahBE96JbvXpvnHEoEoq2yLFBgAUcPDX
YWZYYsATuIJ0KM8V79lISoY7ASO8qokz7pFNPvV7hMPcV5Y6aYqRvB08p1OQmQQNzPIuCOJzuzQX
eh8E1hU/6238KeBQKnkIk+hH/BL5KzkrFXL6JJ22bVQ9hMbyeRQlqGolr2hTkQcxvHXvjN6tuYEv
1T0YxxR4oFbDdG59KwMLTFL7yteexOqROtXmfuHWCnvmmnC9VqRFX+OsX4QhPxIjxxCF9ZLMm+tJ
HOe2jzhTk39s0bjnwDHA5XxjQmYE35eZmtJzhcZ1mSzzHVRYJnf9L19+3/2BWgnIMBEjU/uoMBU1
Fb+2Zxd3KQ3J7RMZND4I+hHjOY8owVAEKcvwa3efwdsDF2V3Jmzb9EOCG8KlZgSzEZzAW1rBqbaf
fqCYnXw5OR9/rf8DE7pxKTDqLrEZ7JQJEo5REcwbAVyMua5QhklVFxUiOQxejx43DHm7wvHMbXQF
MS6iT28NsoTMyXmbWwz/G1xdoIe/tlkAMucnHNUNulrrrm6l17VpfHuRXoRujAJtS6pD10VjtOOz
4a6ZUDvOQ2P0N448WoiDJjW5hLfXNZhyNjjQngqKe23JZzrpwV1sqa1V4RbZBdkVN4aMqu74xyy4
x3ohh8QMDAS6XRl9p5ShpNANrX+xfutWlZttp7BC2wIQPdcT0MVLkBXkpVSXqkhf7Dd6Kd7+sD33
lyyC5Hu/Z+Acyc3D/FXWvtjipKawxrYqFWTZddWxT0uhHHuyZuH8LCkycTnqWze9LT+L7/qgVpHM
rsKYoHuj+E1SHGYn/qLaoWzqC1t1fGCSIF3GrH1cpGGFPReeJXSPllBSOH//puyrbHMIyjNitNw3
3H27W+UP8CmObuNqG+7pU2HXz5QWmt68lqPS2ycaN3Ke2clQAPcE1sSHQW54FBdmu1nc7v+i/7x+
gMD4CqDjZAM86g98CqSI2AiGrM5NuFYWvkYEEJyNZVRXjz0hoKdCBqxHqhgFY377rpP+NF6A8kwQ
MecPS317AznTOacaLruNXxsDZ3v9GpxDaEICSF6v/yTWxupmPOVeqUXsV5ige1S8vIrhkYcKhmMG
IoQdhhzOpuapDMv9BgNKHSiNj/wnD2cJ9SMmkT6MUyw18l1VHFOOXoo8WBL1IXTWB7kJjP7hHvzT
KWskPaKYYjV6poFPYVCKPD+CGLPslRvWm1BJ4VE8cq/3quq8H3jCyPa+eGzScfEkv0376OTvMiJ0
VgX0RbPoMbwNlAWwvHO+2aqxz77VWWkWiJoTFl4SN2wp4VwWmLmTdo6Ua9V02Tx3JT9/GfEiDWla
KDdnoDKxKlISPet1kLe6WvMMWNWkibsh6g8mGwexABf9/GkjG3jReo5Ma4lFh56UObDwiUvrNsIG
CLKSwFYwXVzrPc93TQ8S/LWyAz2lkDZTlwf+WmrK/BuTw+XfXhKxC4BtMnREl2X8k7PtPtEBjdNf
yZxsrJACOiVb+8JbdZVr/OwDRq3UNtDzTBzCR5IlPHJrwDRsxmVqcVnCNKxHnoHCRvIQvXpJR7id
HH1sJpQVH2heGeXe0xluYmxPBSjHyfAj4INGIh89juOufDATbyEN2agLkLQRmAhJ4DzOV2EU20Rw
K4bL3xNFnaZpsgI4L2o8PbS7R0z+XsQgu8vWoQLnRsVqGzZSrkjRGSuawh16+6S8YoOU7cgXj6zK
SeK2cOsVFqPlJVSwbvRt9okEpGEdeH9ClIPiMv76XHPekOJqXqeO3FSsPI1iShsfZ12GmAibA8qk
mFsQzpYwo5nWNTzxJlLfBEh7pnC/lArtqG8DXnxlSD3xbtAssW6aL3GrsD3JU4/vCPMroTwTqLtZ
T5BCWlLIMxnuqLmmgoa/Zfq2KuccF8ao1dW2VCdtqrwbgxdAuOOX7cWzdxXZC6elSvygFLTOUjDB
NIcVBPQ6FLdfY+eWpPv6IOJRZl3MVRM2BWYp2NFDDHSstccTJsLtHjyfvtWI+6aF72H5ksEXDteT
FHwa+jP+hZ1TMgB2h3isBx+lXImHtSOcC+lxGAaoqOuRF+Rn6hI4RLRO1Lk2kwE6DUt+njzM1bKu
kaqzWnBPHfAJDrnamDY4S/HW9vrT9K9u50/017UW9CgQeQGkZSaR87GwTgHM8XE+Pp7jT2SlEi25
FYwzuP57DeSimICSk7X2JnUwldHGgrwU/qXvYyRs9pvDrihRb8k9nKgBQyUt3wUhZi34ocdycqV8
OS1ReFgNfXunNSjQbSvug/Z1BDGadOHFrEZwa9UmWlaaLUl4nFxAPgkDwr86XHU268cjPp6v3nVJ
nPfWx1HI9Xx4BDDcBkt4bmh7G5m8DdHzQ7XeaYNSRtEpM3YjXdDDZoAAdePs9E0/RTZ8HUuGXfD8
B/GB/v2RG1/wtPnq/iIjiY2Jk3/qqVK7LeDwgNsFhnS6EMZafFhFJQ4Q3r80WAatdA95w0rI3gUV
yBaTkliKkIShoStjgSIOgoi58F3rOBBN4upoLEgB5WwIgyzEdRkcss5PHU/FgMWz/yUxNc8iwLEp
gW1Xpnue708eRwZyarpjoXlCmvLlCIqjjm3RE+ITowEi40zcLuwmxM1ssKs+uJUo6DQyY198uQAo
KbUfcicFWiU0Wz8TDtTHO928UpaPicizwYK/hrt+gtnWBDwBMYPpOSkbr8lSDQrE5ycoEGCkPs84
Ya2W+rDIBFV/Xsplb8XQ3HK5TmdrdnSx07XLDlOnM4QRcawDhXCHrcWpz0fKw5/pAJyJ+9IT42R6
MUzyTXFzPl9V/QCs/D66fHHtn6p3e7H04m9JQH+Bjbnlqlj4esuKpkE2pp10XuCGvRZFpWBatJEN
OBRJ3pX+NYqCDEwHxfsj2dCPTyXeWuXHf+5YBjOpBZqbSu0/IR9/fn4pu6jthH3Cr/21o8jElSDe
4R+K9IzA78QRA5k8NuheY2pLSFlhzefAQBVLxbvT/7UlYPDawLPxIjJt/mxwdJGWgV9jrcZ0tQ0l
xjzJGM/lAFJYXdAxS/8DaSsV2ohgBUv2/b5qeh09z8CMkGj3bUyGx3XZ7UqjqNzq1fvVL+SA/w3c
dqsGdxAwDQ1fvKNP1bLmYNLdAPDJ1sVmKfXEWoZkLWFzI1gIyfYQ4Nw1fUzeYJTfUCZc9N/uu01M
HGrcntOCowrT76TYqeA6ms/obNDkC/aSsS2LldK9TKKpAr/v28vTMwenJEt+H4SpAho8/47AcOWt
L3yezM0jhGY7VQhz3QogU7vDd+JYRzT8o0FFrZ1IdkCu3TO764klEkGZM7zzm+h81/jnez6jtotV
oobfgFz0s9rafJ5qctyY3mqd8lTCxT7slazcKoMyRsEazfe9/GA4AjrTjAs8IdbogyTEK7XgS6HJ
3jFdSy9MRicgoXr5NWlZQOlWnRSQA/jBggRyMjnXFedRQjx2WqHyMyG4ZPblBva9yjtxiUaq8fd/
XgwFCeqsnv6ZY/xE+9tEmnsAdESj/Fn7hg6VOsmW+rF1BeCRNH9nrP53WlMbgKAj/wg09cRgWdRA
HsqE/YAkgX/dcBjamse1gnmJ/MKogOl6ECWBr/eZHOdYqrXm2h+d2EJ9TfBYxugtCL41QlVyfsA8
uDJRLDNPWLlHDPrlVlxVfOMt5U5TvrWfgQ1oyqDi6DU6NHjkoeOTMMqVFXndmXkpqvfizlxtdZgr
bjaljg4QN61jjgmQKbHXpBcra0pFJYjs85ruJLmKlj0uE7f+9cvW9NxSA51ePAK0qiux6btvMgss
RuSJrYFNg7O/fLKT0uvomGDH/c6x/DZsdC7I1M6zY+7RFg886JMP+YbdLEI6X75HAd1beyqjzMMs
8jWFxCSj3Joys4b4X4l9wTH7/ZGkqd3lnSeD9NTP5+JjbRlkbavfmlkSCeior/gdageQ2qnau+9P
uozXFoguODS4LJTgLOmdhYDxUU79X3WVRMruvQC1IHb87cXTbKlZ35lRn5iY9jcHfP8S1RR37S9s
bAqUR5zmlnE3NJgLdOAg7iXNBKe08qLsXyQL0ZrGo4OGclTGuDREwQ01IYGHt7pBAbB2O07DYyJn
zN2f+P0xQNpKwobvHQgunX6MinGB1tX1feQR51FTDxdqL9qTfRazw/phViYCsvxvcJYobkv9JVBR
mHq2MRFlppLnPwBY8PinmwDiGBOfYADtCLJ33+cASGMB0vfS8D0ajp6mGV+8VyIuJ0H1bRJiCXge
XeKZyFz5q5ZDRlM4EQcI/K3y2wxGXWHOnr/VeoJ3GPkraIfrlq+xMOqN80uDQj+j4tGhLdl+hGe2
C7nl69DfBoTuG8JOx09mjQuf5STKjRCTi4ine0HB5bghq2LdJwDlLdlgnxIlB0T2BovjzfrbIo8Z
aULfGIArsGwmGFAi5tv4bvSF6KVeaK/Ua1fgwew/KYr7iPdQEoepNeSxfIlXh7809U8l4+ALNCx9
U61ANGsGLiauvRKhpuOndtuTZ3pOXW+nmObxtEjG0u2b73Piaxw9i7JSrTi/Zb0AzUgVfsWlB/xP
WPvHPIg/8OI8rqaZ08780LEJk2UXHbKSN4+hbsSwFEqAZ/LXCUT6C8er0hy/rjiyAfAGdGAtc/v4
7RjyLqhne5uscR7f312L1X9DHH0g2ZGF9aLvaGQD9wKAE0pxrPp8TF5qaA5qTfUYZxyoG4ErJGrx
RjTBfDIeFXq6hEy5bUxjiad0nyQioHq5yYvQtUkt2UYskTvcvPz12OUvmb5c3537R+HphJh9HuEA
an5oEKP0x6EE2My7nJGIQi/Ek7MKIr51K5424sGaGGe3SyT2PxZPvzsRQKi5WmOkNSJ3+ZPji6Ms
9uCcXNjaYfL9xc2z1Ij/iVqu9EPGcpW5FVY1f04buVXTbSx2XBbkhidOowMoNrmWmv8+R/tAg1W2
EXZNWaNrcfN0OMQraurHoF/VK6ZIMXpcOEN/jvyiRXqky/iTGQziqk8RJScK2Q8t9rgvHIk5IMIa
X8taAYtEK+VVA50jnxRi/K23WoVov6LJNxu43zt4PTj2mrIU606J6ugTpCSZygj901sQMt7D689Y
yeH2+b+M6yFzxfWpaSkT24tA2ikyR3B9Juw7T0D0Cxm+vvfpOiZwOJBNG+W/+20l8d9BlxgTm5l7
Eeixe6gm8WKooI7BBJwXfxgyLDQA97uTh4bmNsRoe6RDk4TNFX4EoHhmMBw2wLOljZdMKZmUV9MA
Zq5dnMRGcIm07YH6Cm4cwI3yKvVRLjCJho/Jachj7S10kdg/Ckn3lGTib8A1PP07W/wb5SnoJTLx
pGc6yIvnEhptrb5fzq2hcFFrdqcU53VoYtZ8vQnP7zVZ0uTuwwDSmwPxCFtXTeZNUJIZ32cY/GQZ
vDVWWws/E+MKyvx5EYtv19HlMsl2PXvSU6NqEsnRvu2EAYX6SG7XqvxieMHBY7/6hfi7td7FhPIY
MIAJGEaF4Ju5JZs/xsfgQcNqb6abhq0MkUHEQl52/L2gY0+ayU4+rhx/0vrusIy7cF3fG2Iai1fZ
TR3x2bnZQWorNf2TVmRjtHpASQBm0gP0BlXMfh7c03acKJfg6PhDmcQ0tpIrMyvpUOg0ocbZFiFI
Lkwc+yw4USRHipUzdH7bfteaalGUVYEim4mJyNcS0XUEiiBjqOSCXn8ie4pUjDHOJzMEwkeCzSzs
ShbYHZYd/M6Hup8Sa+VhMIqQ3KoRc5R2q3DgCaq7xM1MC4X/aQc0x/6g+C9THh1ohASsXY3G+iGX
NJF6MnQMY3e0CF/U6mHsNaYaRvgmz9rA7xfM/9MKvHDCUpF7KjMD/bIH6aEWr5v9lwWy0Nd7OibB
pl3CzIqN5B8okW3RTNbSu9K2DvAW7A4Oedkf96kyCQBjlykK0iKoMJN0/0g9oy48HbqdIeEGQIm6
JqTU50mvs72XJbnl7402mObs7/aSfk51GF9dFXlhneAjbbroJ66EwbsTCDBda48/7qGIRPixjPX6
CQxlvKzi4npRLQQUDsFTGTDp/w/LRbBwjTyi8Sfuo7Gq582u2LN5oFQzQ09FnqGkKZ7m8TW4L9ea
qnFO1f1qiH/Wy6mdJ8GVCusVL4+xLm1YBV9jeTzdhpBEfyLE9LlmY3CwWh59iN/rpb0mHxsbWzmV
XNFPcJUh1qfWvkQDvXQPK/Nx+D9IgpBuIqmAC1Ddb5Ko5N5Y7iyDORwGY7hNWy41qFfzy8A7lv7N
Fp1JmhWBc6+nwjfjiHV2c/YZZB2Rrz4t347YRdBSbT8BGuAVSfByDC+rF5iQIDjOJuRXUh+5o7f4
G1yNxby/Mu/aHuLk8j6OfCpweV9LwoMY53+oJIefLcpW7gei37S9F6jfHWoeeHn+XHa4ex3lV7eC
TzehFpDKNuPtSa4qZMtBM2/zKK750t1y5M5bfbPWp/G1rO/xoPb09BnWNAH8/lCwe9HBd10USq5h
R5bigdvyy+mo6/6zTd7ySUcLmxct1vxPYdEaSNXeOWKF5scEE+itJMZ67eJpvwFzfUzEgUYkHGt4
8H3PMy6Qs41mE/t+QBr65ed2ZljMzS8SzXCji1JrZ/iCS3ALXI1HFG77k2Ul5rQaY+E+fRP++olg
3gk4bfPg0m5d9HHMPCyj/akGIBjLNt9ycLz7gXYEe/u0r0vojUMoSnX4EBk7IXOD2jzkmNM5p+aA
q/4psMN0EPIUB25kC8C2rfAEnfg/WiG33kjPWjRVyo3RhwAd+0OpkH4aw7zOTUd/FFfLaq9WFZuj
g8ZdTYaMkjdE7aX/9c2eB5NqQ5xdndw/sIlH5FrYOMaCouBke3KoI2Z/j7LEQ2V0Z6FCHFS/RHP7
iV3Pxi/N8vDdd7O79s588XwNal17/1qdwZhg4f2dtLoBl7JrolO0E/9WTbnP0g6rgxO52MHVDMDc
WHDtqhQSkHWhMGKcq5T0+s8uns/YKE/USapmx+g+a276QzSwVYmZGAJylCcSoRJm3eJvpwYVCMcY
3ZAzJYb2uCc7HF166dvIeNr1nHDm5FCPrkL/8UgY2PXlcVuaieKO1JLgDbh8ciLvSQAsQ0s37Ynm
cyZOwlHyve3Z10dLPFfx4gBoPwMhWkcqcCrWsq0iE+TuUCVzMa5DoGuXV4Bj9FZk6HF5wlSOBrn7
UWjGjcde3PYYKiz6QnP5OL8ZK7WdCy7Br3m6b8PRM8oOKETYJfb5BoY9KbxQpvMSEOygIunpZuNz
8xakmNi+MWkE87+nj6kA8c8H7hSmFwV4lgbY0pavQq2niS48zsmKFyEJCwg+zT3FSxYkGEK9JAhD
OGIkhtkfos8I7Nmja02Q6XahS9j3h2qg0JKwVQXNgR7WhAQ//gX7tHz2d1z/Knf70BuJXhU34py/
3VtBI/8YNJ5GeV/vmWUgkPO+9mKqmCFktXVTwJRDoacTNUBL5ivqGwpZGwexTh2BZW+GI0jMhtcq
GPzkPUasNHaMkyVmRFO7JeGOgGCu4pJPCsOA5k5trO1Hgts/OPMBkRFMKhumz9qZ4Edd6HTo7F4E
8GHvhvj/kwjajqzqtOgENT8l7qb25znzQabYAdPxwEU4oRUsARiWgrTNs3KLvQ9a65/fUgpsetHf
ukqevb+sltKd0Upx7Z7MqO1Igul24sa655GM21KoNc0CtgwnIYZ5HG2IArKiTMi5XfclcFjo78ET
F03Y1I3D0ICYSRHS5kAbQY6x8jaP4GAF2nK84GPR7vD0y7gQCyFtCnSEww9nDTzjvosYCEePJiIy
+UvNKdjLBkksVLL02DM3ZsQWb7rvwdG8zDlXt3z2kTHgWpRvziYcqgyxjKiGX+rFrEtZmjtT1YWc
3qTNyB5c5Ua6Rk0vlJF+AxTvtjWgg99NVdrLBy7cwSWhrixTlUBgOFM1OwkfoLqdFEaBa/gOqdkH
ep5ylTysBiyoPi0XVQ6BZLeHxePkEOwLd7xkxe9UdFbElkZRMtt267MndppUVPo5xHkqNuRmKvu0
2z9hsggVUW7pz5Ph5sUNUBW5sWy5z7JybZAUTRZ9uGj+Ne3Q2ntC2xesanOMt9vZp7h3QHrvbH02
+QmNqw1PCTOn27KDk7Jw4N5lTXh0JfEGLLN0RQrjxU2X9SwinVOxPFpNZgLGIaZ77LK1fW0p3hnO
VaFPr5w8ctheR/3qik1pta3pL5Rq0lEM+qCBWpYSl1dPJYgdS0FMu8swNL4Sa/yUQOSHbBZ4lu5o
RjW9x+r+qMaEPmapLuMUyo3WbdA/HBEO3iW4U+cPT7lS8LSACb+twQEhJakdE662snJs3+JdaXlx
AELgPWp0u5ysQNJy2h65vWZBeLDGogOli+papQDJ0Xsy9VX30G2xU1Yu8gvFCrn4QNDf8VIG7pXc
BdIUmANi3qMS+5HAgwPcKTQPo8oElNEgtSv5Qjk5piM0fWZsE2OR89iBW0c4p8AD3iiO/HVkPb10
BuzcPCeBBGOaNLM01FVZg9YvUHHoQ73yITNzPWG+NfWPBhADhI9W/7CmRwy/FMKYNCD4o6uh3S64
1uO3hmSqmsmt2cOYxNyqm5FfkWLdSmV4rXnIIgstmUauiNa+aFZZ/D4ZNoCj1Uu9t95XI5KQDfo4
BKPBDWHcYsB9P2Seyqmc+xNkJ+u//lBKLq5yWq8yfwo/9wyNe2M+LuV5LKQ8nd5Ta0MyqEwQyPZx
OMfCvGJyyNozXNTrQv9zLnmjDFuE8Xsy2jfoN5hkOezBkERAsQ6kdD/vbzPoMQsIROd1OvVM9Iwg
QojA2xCKQEerkFcOcvOWNtmH1Y5xJt8EMtatB7jWwyHUvasUQDEQehoI2qJyQBngyQuNCyiTSzxU
uI47TKcjAysCZ2A2oiDtOLTMDlydLlNNDrpPFr42Cx3uRUzXbvDfmzvxHO6qbb9ppC5xrrJE/wrD
TMF2fe11lguTZPX5VKU11mzNuubGhx0e4AD08cb+/BRDaSAhk/LDEvdFOr4ESPPisDu2CBQDdrN9
0gxUoVlfn5JCkDl2vbLTVkkyzbZBHnWGxrWixpXz3hkLQhIXLVIutR5GQYaJRHPyOd0idOhkuPQA
axAXC0/DQXTS35adKxv3XXGq5bxWPox8Q2AWgdnMx2yDPIG60RPuB9YCh6kH5SlxccgDQioyQtmJ
CfV9jE0fF2yhURPMYqfkJuS51pA848Y7iZHLK+DsoHBxh+BNC0gZnARTeNrFYhHkEjGrxI2qeG8Z
Z0nk6fc9JQqk1frKM/frRgDT0HnYDLx18pQiqUsLTpUTxy67btvafRrjIRdP5a9sIv81dDW7rsXt
RLPQajfM9gBbfT6crWsFdKfSeYwyQ2S2HVShgTG8jCyYCKC4gdmITd9rUBcmErCzlpAcC3GJCyam
cf5G4vi1D+HA9E9s2A43PYDQ2TztDggj/VVLjqBjeOYNB1w6/6Nnp6nBqFGfor26cK4C4ehqw6aO
zGxtGPR/Ox1eHEyTE+Spda4WL8ce7nKg4v6buprAuIVgOg/MxfDMieWsS8IWkV049TnJXHRLn6ht
gFDNj7/bobW9F5+TxBk4VHgPKPs02AbNMuSWXa0FoDA5BLsCPQEr/PLChE7yf01YbrmTK6FDgBcp
ztS/FLpKl6NXx5XhXyJbKwfKx1MCUzMLYgbYAdyt+zDSsXFgZXDeXyzV8Rjs9AYAa5IioylNsOnO
PT4vF0rSTS8fK8p0CVVDMIYu8oRRlHTQJSf6WzAxFdwlXL1c7W+Di0j3er0FbBUu6xaF4Fu3tB6I
TVSHhCcVoi+4fOz28koztamjoaibEMNupBGsZaylHGrJr7Cna59BGY0cdy+kcOhApT0FGjzNIf1h
t9kY2ItDPl2I7yhJOTMGGFZXaWH3/opiUpeIsFaJ/2rsUKn1zYEPV0UMJbc6B/CwXXQTZK49CE+l
SJZmrlGhlCUFuenLioAHkaA9sn3P/7FgrtWYjHoqCPB4qLraycRtrGgQIXwm2fJu4Lcck3CBRVKV
uMfGGaHDqdwUDLrla+SEkPzOhoF14h314/q0OTdSvV06AluJ4oo/5YiwPPMZRdf/HDgY/YKbWg4u
lKYw+wG63NCT1Un4Jm+tIIrMuaRmhQx78gSU2H6xBsiuJGwYcXtqf/YcrNjOKSgkX+1SPjcY8gXa
TyANpkIMN6XvItAqrJTLfg090RnXqV5r1EB7XP1VmlkiYQa/Ah5lNTeIXONHlYpBFerHrpc68+W3
oBWeGEn0wWZq93ZXrDgRoFmpcevAKrSOOpaAsjHUGtTqwkdxnfKMZYb1qdjsLhm/0pkdtepcdMMm
XxPY2df6RlARIzXvCoog3GIdrxeRlB3IhIVeWGPGBz3RWd7fl5h0uM2Fvy1JD3l6lWghMmIOBI+d
3CjPQJ6WYRSr00//axK8yq1L60dxotd6aXgjVCmMqE7gzIow3LubHiLHM+lQYC5K1rL9xfnEjH9K
mB9LL2ISPgPl/VKBw9XUB1rk2RdIIuQXn9CAPiPTqy3BIpa0nXW1RNbiB1/A8HRt+lS+Bd/czRpK
J7QV7zYf9q167sy1Z4anXJHpKs4ac731ozPzkPiWBTGcHzdCCqtiRifynvHF0cPVTgAOK9CIp8SL
AGXAGYHdIcYqA5l1x0QqNS5JEgqS5sly4I/0y0yonVXWeg/or6z00xfut2y/okIEVxwbQVRn2Fsb
vvVLEDuBAClvxtDs9fzOUpLecLJauFuP1uxj8vn2cMAQ3oP8bWer8JfmG1kPV0kLbsabUemKBibP
VKSor30EmzS2F8yxqNSY1JVntGABSp0dOA8TQM2CCKvgPC1VZGrHfGMMy9LpFj1sEFeGvuNeaQE6
5xek0KPtZgMvxwQ04qg8PS/JFXKsniVugYPWjuv3O6iZC966N3pG5wdHt9yIcQWIOh4TW2nFH/DA
npSGzbD84C6/BTJMcl7hZvF6m2q12RQLfrVg5wHrY2oq+EbSIYyZ0gA75arBeL3UgSiipIiGiz3h
LxCVHIMBoMaLf0/BmYmbaW/pT5E6AaNqVFQ7S0MW5vd8qcjDF/izoLLBOyyHfL3Yu7olcow7HAMa
HHYqRKx+M9RnSie70mmT37L33xAIBIhGmIGAal6QR7l45a/UtNBbDsr8i+9NSMuuKp629JcVXjN7
9OTSbMYtp54UJx6wXVSDnRkYbFZCAuds1v8AWo6k+JE6zmwTEMfrhZXnldcmv5WXZ1pRJEsAncQo
21qouN9mdw+2qFK8PXcesaYwp1F2bszmcCf1rz01g4/x93NJyX/of/hgpauvzxHkSaoP9ZParOtF
6XiSl9/TrlEq3AIdi1G7khA9LKa5SDLOXDzpFtLZSlTmODkVIIWhT0gXeNANpj78D/EpvEwO9vf0
NbOYGZ8uUmrP60zV+t1PkyYpzKHaelA2mY2XzJnEGuRo0R7i6YSW6VudtKTLxrKN/u4NKETJgYG3
RzR7Wb1GU4crqP5bhDYH802KUGflXKnRCMCbofM/eEU/5d7GHRwlNMFfwkJMgOBm7PPkiwlLen7l
leftXY9KJmz0GecZVwXrMiwrSKedmrvzIywE8bDNa0bV1Ld7sWO+KM/0h2+lvUp4V02DyDH/2ljB
hRwhyGESG/AqWIOowvPNNWy/QBM89yl/3uRCcAgDVJOCy4aMVYnhZjemtIu1smuFITuaJ6OlHaZ4
sQepZXVsOumnNUrcqhnq/Mbv9Qg1JcO4ujalD79WySnxfZ0zmZg+o3HP4PETm09zAYOIG10qEtzF
DIbGDlx92aToEjIBgGi4SdZ9iBPqkCeBh+kkmiX3DLYcG1+zvBz0voWHpXpvKuMRB0pJEoLsdllm
FoNxYoABx33dC6y0TlFJLlvoj7PAUQbC4uzDkFylD2x9SlZWvtjm9faXjVzYxSe4WUZ+4FP9T4uY
5PAWdLF/XCtzzAX2WuSsCfq+JGVkfhWlkkDZdarKiyH3yVD+f9qgm2y57XTBgS2whf+HWZoMfxzR
giUu1irdksfDSFWWqZ7+dpoEJT/CKiMjKOyqfJGBOx4aV3zx1hx4VmfhzkO62Kf+GpPREsY2EHsI
2F7xgQjXes0VG4jHiczE7sCA+fO5nZ6XD20S2krewqginYtw3rjklMJfcl6/H9xGIBNn4j7Q8OYu
Km2BUG/N+GrVcwrIqeY2obr3NGBOChvg3JNKlEa7wbdSPBMc5lNj5EStHT5sJjR34rB7ThLICeBg
lvg40DRhZtLLOuJXush7IE9hCuqNPSGo2MybkJY5F2JZb2uZekwIrDO8HK8xhEHiVpIYkEJ1RQXK
rFwI2sedPIScMdkpygZvgGxXy76+w0HzHS/W9mC7rEj4/C4G6SGLgtlZVWdLIIxbpB5++ZLTEtoF
z7bzIV9loLZqPz5KT+FbUyULyhQSiGuGyNsD6DJX/jqoGm+vE+99d60cStZVL8J4DnzeJbRpAq+f
IddJ/ITbwsvWw4j0GwTCl7Z2osfd+zTZNve8g765YFGjWztPqosPkG15kKkugHer4/1IRWUVkCkY
hKUTP2DDGwrU/D+BqJxnOQcpDs27mwGc81tl62cqeHUwKmsiiY5ZTo5kRCyeqW79CKd35/4MWxUR
PuIjRNhpVFFRP6QsukrWERdlja06PEMDu1w66hBLMVeJwjvIb8w2pV7UnPOaLE644L86eK9f8nDi
X0qP4NSTL58g2Gsfu/mcmKJeAcN5uYUn3n9ohP/1SKvaoLohUSGk5L4Fabf2cMKNAUX6P111cH/u
IXeCsgqamfScYehYBZmVLWBCoPf3oyL0VAmVnEZTZBc46EA3Kedmtg9PRpoZT0iC/0iy7S+DavVf
WocvGO9TbYucHA14//Cg4pi3KN2vw3wB9DP8h0yKAz+9+f0QsbUuD4PwVcANekkd4Da0spBTP+X6
bPVwIk+s56PZeJqBQnnBzQxHTTTbz0fXWckx0TXLuLLB0JQB7CzB6KKvRvQn9eFEU5O4lI6MXfti
woK7YEmqJF5Wed8vg6ifXLp/eUnEfxkR1tKJzlEk32Qb7Xnso+leOzlMH2cB3fwig5ppJjWP04I8
6xIf4DvVzJ5jll2bvZ53tVvgTlekH7j23A6ZYJ0/A6aEZ702qO11ex7tzMxXAMqld2owhbl8bQhE
c8Zu6v0IErOhQW0zamcEwEi1DwV4a+jnypTQuYWaOgJCOrRarourWIrGb3+jOOx4hCjpXQj4Zu0/
UZd+2pzuilR8e8VINDVC2qK+X3DVoHIWZz9Ypr9Vl/0j5r9WTBU6qS55Zai3gAsLP/RZP7Hbd9Jd
lbEkJp8A0ECwn7f81H+FX3hHwJiuHEHohYKaWSRtRZNauZXt8yfRKaoCHW+T5pw3LP2e3/IgGfZm
Pg7WRAAqlaV86F/vHd2NnOm0X9CTMyjRrKjiLgmoz4CDqC0N+njLS25aNjkR3qZWeMgCR64+pr4j
58/rRYK61qTbJps78FAtlr5WuzqSatYfOYI0MrRvViAuFeBghfeL+f7xQ8m3rARa0OAKZ/5bLFJ7
QtzBn2LN6ovSoJU025lgJFHzdoRMFttEAbzH/zcfak6OdSZUpOy8JRMuxusQ1cMvqpRrefTJPo2n
baV0p6HtwR20tA8bYteLWLHsjIhDeMbvno0AGQUd+ZLA4o6QRjRjPcX/kNXpcfXLzfFogeyo6r/f
7+v6dohwJj12GCtc7Er0k82cO+c9xVY8Eo3RcqGMRdZQ+WUvJX51B+7SUML0aStBDeqAdKrmi2vf
B90aYeVBiFMgJ46o3RCJYRufDe1t3qgkSmEHqzOPlNXYYuwiJ4TEK+2sW5CCyqOJ6aD1tKJfj5Zc
/N+q6pDQosfZ7abu1pNu7CzPPSxv24cQEKiz18fFFq12ReJ6Ncl7nq/ZRe7BOk45I4Rneueg+q5S
mHk6K+9NaZncYHpBJMVRF5ZqQB4OFlQmr/8BJMq9ALEFwouYVuCn64JUshfVEUPygyQnQQFRCiZT
Ft3tRui+o/qeDgTQcuXWA1KJ6FQdNz+c1AzmTredW4eVIuavI8hFdYHWdXYie90y945jt7YZA7dH
m4ue7wmWKJfo6r+UpZtXNwbhgZOcl1uyv3y1b1YQw901t6v+1qRtaYMTjp8yToSPDM3tFUpt3T/j
huKGxRCmO/Ht2qU8cTfk7Q/8LcaJEuhWxegv4JLFgHtGmfMclDyXDPDhaj8O2eqsDR3ak8oTG/F7
y6Ocg/Pk5Gv9t8HzjUkoqeCxvZUjQCCu8mj7bNvmSJLjNcdvgQ6H2jf+dxewFpgk8MS+a5VC1UOZ
wD4pSmvyeoKmktGZTxJfhlGADAz7At61Y3kee25NgawDAgoycyIW+VNZKJgWBJ3cua64AX+VBQ6h
ENEzjYQK3zW1sgdyI7cs/KhkhfIA/lQvifyxrxZRBSVVblnhPPfznjc1QPJuUYQqjmCqxujx4Uib
NdkzviDgnykClXfNeuBDNpI/OrufqyMYJMSenEvDwxGYJxiya8AaZHPbWR2a/MbHSesVIEtJhBeT
abF9fWJJQoUftYgpLSD9/6TxIAKy4KbY+ieWDq0R51k2ft7ZodX6zpS+Ox68XnL3MRquxZHN8Y/U
Sa6oaY1Xedo9dkxHJ6AKCHlCf3pU4UMG3z7CwgJZNlobvIDqvOxMIa5oDwZds14kcT0GBFohKsi4
NMfXv0VwzcKBTIWlDvi1RwbwgWwKGzgXBzZjc3Lm0pdMk/OSjS0fkJNunvqeWFmamA9dhUWC7092
wbEaKe1VVKDKNwSDJerArW8sS7e6RO18itXPmypOchVmOd50ihDxD1APxNU0WPzyKbAmzvcvxuUZ
i1ENftt5bTwV+HJdIpAQiyPyEBDXVSB/qxE1yahzYoMqZbUujAM1K37DhqpONv0kVDF5mSL0b7h4
FsEoIDmxiiXw4tchVcq+eMkedoq2cp9lMYGN/aLpVLxWEWT7bppjFxQjfz57uK8iz78AAqOYDP/W
k7036/PsLoFEWySfw6tcGkkD00xLVUefppa6KDOokKPppnDGJVoPuulfnsUGpILGEUuAdCzw1dhR
P2E0rK4aiZ1RIko+oUeQrfJUv1X/GBMnaQNtVeEKHRzT8ufIYLFBBkQaL4Ehrr+W238pZlFWRWe7
E0vKVZHojamYz7sWSFnhHcqWbZGbkpisfLFLRpLpDHCrzAaqYfCtJ5VNYXazp1qq9Yfv0svGYIgM
Vw1fPUer1//8b5CsS59vlZrQYXmpFHtg6KJhbAVcFhGDkQllS65rMypt3Kz35j7dBOILCWqtHl16
AQirtdDy9gg49+VLgoljhIaiLBUWz6MPbq7wiheGOfKwLUCCKypi0Mn8DTmfSXchw/0/2xv+LCy7
/mk6vlMSTYXAKMZTACK/Q+vstHqVbKWujwzow23B+XJJCX3v5TXTj5AhcYtI1DEbZuWFb31aYo4z
5sY/DjWJMnbUBZjQzxzn1W7hGtXJl47/dgEuXdmbJ0TxbUurClsowwRdl+bkc9xqJ184kvIEI0wJ
hg2u7LGo9fLwPVYe+XQSeEr/bVRXwat5Fyf3M6oneyH6cc0rSPh/BzYwu6jjn3lGjjWEf5poTrEY
hVo7/ATGvGCoK6f8vvWZ0rDtqAqkwI6Pq5qi6BL7MpTvGoGByU4PsMPKJsFGo0M1DaLNWbH3i2mG
FTO7uESFgCLPTPbiEI5Zo7bHEALfBoNTtQxp2R4QXXgh4l3d1MMsYD7tCq33kezc6iv1NYlv+nmK
YTmq4S/2X2XbWrsireoPhou2ZNv5Ej/9phbdU1GgNuyyhbs7VxXzqEgw77USdtTta5s38LgWM5Nd
dbHCwPkyFLFKHnMb1gj973P+TeuabIApb0JQhOJh7sSjdgDue+H/N5zcPB3Y3UZysTk3u+JOF941
fH+qECtmATO6EEYUmjUkKYh804w08E7O/saKjxpCXy1IcmtL6O3Tei5u26MmFJ4h8RnM0bB4FkWM
yWMg79/D1+gbJA7fWEs1vYmZVZ3lTzwOdGDRrg9kngV3aNte6sNellLVE/kqx0uI8L1gviE+K2ls
YJ65DBrVeMoPmiGOFTXJGkFNNNOj44i7i5HHdksvi2mR2AmUEhjd5fj3UI1h/it8OGbG9sK8BUk9
XmOZbLwbSf1yglhLVFkvmVLNA8a4KkIwmoUJBmTxSRzzvEx2950HbRxBeIfr6z0s4gtU+vi2Y48v
PpmCy4TQ+ffvzRgrrin3n+NeTFbX8l0S7OPDjE9TIdMLn6XetQ12bH4OwSByzK5XFjSm5sUBC+0D
lGPeFjC0tj04MopfiQPkhA2tIP+B/9QVqreDP987yQgpVMdAaTG6E3PTO4QmCWVZ8PDxjoY+7SxU
7GJZy3eMf+APywPxcSkG0d/zx1KJmsv79eiJmCu2qmE3n0DxD1J8JeIzTeZc6HMsSUQBIaJ41UQ/
e5jXoKFbDGhpYHubJLpHJsewnOTnLf6ccgZocn4awPDJD5tPqNh1cIEeV8OSuO7BP8UBQ30sbjva
6XV2YyTj29Tg0ojU0lQ6MITtZ41/7GaZejPjEh0jshBZaOxKmCsOzBEbUdyraxkcHREhE5bqus3M
znpmbIip10mn2blfFZD8xT3qyLXlKjbDjEOp2vV4JqYkX9l6GKNsg8UA6vIRYXSD0t4/YnArAlAP
O4bilBcbQU6Hm/z3cfongMnPxR+p3ZAWauDEDBd90VPHLecGXF4JrD7QvaAaemhfzQ7E1CmEknZ+
jC8Q5eQzPTvvUp/HdpHSBoH0+qzm2BaBtZg0VK5bViakrUWBoFtHtHNtyiJmFEGtKGkNe63GzOin
SfSsyCeIXfm5Yqa+Km+PYVlJMnZVGbyyGFSm2LiPmyLbU32ZqdpKkgxZbCQxNgiBCZJf5wq3DNKZ
Aokll6cK5yx5xhKYPrvYz09wrrQvBL4lbZvaVq9qhRi8QiGAPpzMKsPbGGAn8ODXq1yNERAsRltH
G/UgFqa9BjMYK7lf5IqXGHW1OTLO0b0YdmhUYhTEoajQczgvVrDpvlMi5hhQrzyqd+xxjQwclbGD
O9GUM3UZDfGmbca+a5wZAf4a52n6/yBAVGg/STfdGKtsZUdwoitEJQ6uXu96I+ihvxhNdkRGrRK6
EwHdxsfHg/I7tZ7XhDuzEUIuHcRHDIQmzFxByyfyD1nK7G0lgRpb4lpt6dG26hMBL21LOvBNaiQP
Yt0PKjhixK/K/RqbLaADcrbuLQcNuxz4yQqg4tFRJCnv6BOziLA94okOTNMzy7Wme4g7O5TTTJM1
hNzBqDpt3CGvYkqWoDoB/xCww78L4WTm+xSO+9Xl9qUQqd9x6BGQQ3SJadpMOnuEtIQELUrZutKI
5L3xGJ/iYlaGoDaAZapUjHYxsiFIdE83Ynf9VFF2d9keqClxPQ1jl1FHyZGH85CPFBXZVG1mD9h/
/u3Id4xoPdg4Pwjf4+3JIXXLlc6TtB/OiP24Si/9qt8uWZA2Pa0ZqWNy/IIRrYcrRUWUZEK+i7OA
O5bS862r/yO4uZJb4kTYV1D3oXqw7JK82Lz3ELJxCOZPP+E9+LmW8gWXPXcH8YoX1uP6Z/XGBYpU
35rzzxU1688Hy7DrfXKEcf52SbK1H19rMhv7TOWb/kOyFXwUdMD+qUlM746jkfgWytahrgnVvRtj
UFeRAuXNUV8UuXShL4JCk+WEoE/TBWrKd1Wza+forTkdfBmNXDgIdxVF2C+yggiTU0NTPCY6pBsw
+42GKUqYpbOAd3LuZn+FY/nPcKg9I/cW4ce5PgG8em3s9gn0ddfbfCkvpmmBWXKy8aZUxeJTQW81
G4Dnd98aW8Upgmaa6w3zTCIjtOx0n51j02Sq+WWhubCECn2H+4WnrosBj1mLVJ0LdtOdENNd0s9K
4hHiAbuIpDhuJR/zQI1xB2Q8AxB6RyIKaLfGyeFUTw/YSv+1WN1XaghzFogl/g3Q4AxTM80lKPDK
J56cbC2kse6lBLsxYYWVnBocNiFHj2LpDkZFeajB4hxgCVt4q/HmkMqxvTrl6uUaNfzas/OwrRYN
zji+tjHJ1A/UWdyUpMPUxjeJMpxGuH+vURvXfE1kWrgZ2BoSfLJk4rQb3H7uk7/JaOC0uqsIOVzG
6c6OKL69X+M2UB4d8KNgkRwClP+EmDAnQwqw5GMyN7zRKCfbIsjjQhvmtfRBkjxNq31kUCfEnBrE
W+Du8nREAtww+/0wrZ9hnDD3H77B648+88jWxnkOHVOaY7UeDhfsOjK5w4wTFZETE9NrL775Aawf
M7gcWtGTM/c5lGGgP8w/5A2rm3c3vphaJrO9C8AuR4Ua6jFeANUop3PcVyOBEfGdxQB2xASK2Pzu
SyNpv7TADTbfRaHx4IhFol+ouwAOn1/rtIrsz5k2Am6A2Mda//gAx0B9mEPh04/WGIk5qul2pIIZ
zzq8ilruaCiCuvVPV0SpGRDywR7qM32g61fW9MYHO9sRlZr5xHYK2QVhOwjYnttjViBjflpqQOTA
TO0iawfiVpCBmIF/29+BqHmK2CqjQvJ50qAw5YWLeTJszTva0E/h4ferMR3m8Yljz8jW0oPd6TrI
m06hcsA7GWpNq5g6163cW6+mO9w2Znv64Z332j4DA/wEhfChbxQYLeSiTHOhE4I+UHFVY7h3uqc9
IPxc4rquDatDhKMoFXwoojhRMlyFIaWc3wmneilKLPC5qb/DU4iyA7rk0dfdRuiqiQENxNDR7AYZ
hX7hAAKLeujfcVxekHnmAXUhOIbBeNCKsbZ0vRrvUjYS8YI601G74IRU+FrdTHNcQP5y8vzNcYn7
SAPHvt93eWQp1M081zhsUrHoB/EmGb82DJO1+GMwW0E0OF6XiHfKK2iP+0j7ytx9ALIo1lhWqDTj
BeQQSiGw+9vT6KyTgV+MoqG3qR5kwS1EFLYeQk4g4GzIAsjwAc9ZrelWxZLUbEdF+Ddg4SobDdBZ
LFg1nDvbatwf2UrmtU9xBzYqcIlQ1DfDeueKfHfbmDadBZawLe5v6gn5avltS4CGIQ1jC0ajsokH
7msjdg4G7/35g9+OCxliPifRG8/aPtDL/iUTdAwwLYcV+69ozmEtaU2T7RLTNQjB/H7Fv/idK5m3
izg+lTBV6evc+8BUVZz3HIEeYGGwuv7QVjN+K6IdmnkxVn3hWZVR0bdlgL/+VK3m+JQA2iLGF5Bp
wmrBiHK/pGloTdZtxRHd5uDZQo3DIV14UPxvF2HQalJabcvjpnM+ozxYjK/fx6s4fFe9EMZP962Z
R4nqsoKNB5AfaeBjvvLuM+nGRZMf/PDXGq/Vz6o6GU6otsgY0NNv3Askb3cEyYN0XKqlSeoPCfkl
NvuCPWvLCBaoLRgPA77ZeAyRE6tgOH627xtXV8NWShwFAZErEi3C88vM2hPqhxXdp5d0Bc+JtgIj
FNxpdz1vo1nAqJAGlUgI7zUPaUJ/C+qFa6R+Fpw2wFcnwrbYzQ5l3wD28vWiVh2w6VDpeUftdID6
TrkynBJtMOMW6CBK+G2DxNvWyglFLXuMJeX0v00Yw12ukwGczwBf/d+SCtplMNEVBqQyq99mqz4X
ZI9f+GoCiimMGIEMyV/SeGsCNd+jg/owUUTKJR5lEXKV/rvXodng+KpQd80DHlkLvBDu4wfF6wny
k20D/I+bsTJvOOINsjomZruvw79iKVnfdO6oBcqXUlfJRdYoU6XuGlp6FKVUWmUgtS9OpYfrOz66
pjvoOz8YmCaNwNcJhM1ArleOjpdBv2Htfxb1KlwKS3UgO2gZP3K7r/h5QipO+vRtGsmDZBAlmxzq
g6d3zOP8iDtYDiuP32bM7guIb8Uvhqa0rF26XgV7GB4peMWlJKstQk318PhkKuP8OmctlWhvImsI
qzVvf4SeIpnhe1dy/+6MF1OMyl+iXOKC7OMOGlYwFFshXmjuubYu7FoRv948Mr6MlOS+aM47ad8h
G0q2C+Sy+M4icKcgPPWDkZ9X+B+ArcxA9FYTh2oCfo6BjGKMarCq07vxnJyANCyVLiBly5nR9zdC
PXvMVteRuHf20JzlGG2cbTGwRRFegV4X6GTElJCWvDwfiVkEqjYt+NYmc2qM9jN8674W7xOv/jaX
UYD/5w8bHLz18vhbF3X4lvN+xwzB9otGYjHLjXRgcPHDyOgjaXjwMLkkznx4M+Jz9BiHfEoFPlb5
mR+qoRMgkpgGS3AF6J6OoQtHyyu/3jWPc8AdKut9FUnp8oE/1JQ7qfTF7F2C/So9/KX7Sr2DPSgz
m2KzpJ1r2F6zNckQtM6lK5KrjXZaGs31XqyJBkdZEGlPagahGbHZ4vzdcjGQ4TSYZ/HUGP00rlzx
2XGVearQDhdCZc1qJk7TLDabpvHDEocr+FsQhktnekXx+71eXRM8fyoENe0v8gfG0HyX3OIE+JmB
Wb7UaO6usDMobFMpvCma8XGMKib3TUUCLSWjYyeVqtkkwFfvXAfjyRizVRkMwFMXWmIRsUk3x38j
z437ReSX3S7CV7SA6QSLHTxX7mS63li4SBiKIrWEOyq3ypQ8OszpmYI4pI4DBSqxXFjC9FUv49UV
/+214FoFsRxziXgq0328ziqjPrjxyNOtH/2VVbCdD9QT8K1K2T/jx75qKepOpm3iVJB0gK/74QuT
em7DU8mes1bBGtE3b9Shxpbf1fFMCVJSgJgdB7XG4vB63wkmB2qtw8UTkIe6npmczXM1GU3eCbMp
lHQbwEczn/mPibz3X3rlSvYdWvc8RD4p4+/2UUuByCe3lLbDILBaVu3wUW9dXs5S/a7w1m6ynjj7
Qoel1/emQRwI59b0ZfJDQp22OrWXzGHUV9Q53aapp+z1umQjygBXy7CuOnwpi1e8C+62kGgzzC3u
ssbcYx1GqcG4GVbCW1XoVBHluUub3jdU7q2gZvknC0b3osV5zUhHEW5C72KFNu0tp/qZbeVos3uA
SBKjHtKmwwEu55rK5rZIMYnfufpf4m+E+ettcEZyxxYXcDOailPlkNm9Ch45xEVdTTgKTww4F6L5
CTb4xZjP6J4gcm/KJStvg1bhh569G6fcj5DkCKay2cimvAi9BgXAxi9/KNqNwLN1WUtQJoM6/HTt
LIuIadiIPxJfQEW91EYjOw1M+hOU1kiwHpk9r92yoGyxXF41VKp53kajr8vzNwkUo0VGltFWd6m7
9xjLZiTiDEKqPgH/zm1RcmvMiZkU5QxEhnmWTn+YeV1Ehtucciyt1964UtFxKSP0hfiUXKyO/syi
0Mrp8iBQL2XWD5PJVIO+hNOTL6MiS+U76Z9q0VptjVZqM7x4p42FEtj5JqbGBdGO9RQLgVjg7sWr
pNj1sQUWS9efpfUVowLFVFoYsERwO5rOv2XAuq6IBAmjN9rEWsxEvFsOpLY/hoHTn1BoiL8c+/S+
H1ciuNzoHYoXV6u8S8m0adj66JCthEUa288aQp8lGkYz/G7r518F/slcrQo0I+ymrekwkVRyZo/t
LSBJNtMgBk8nTN5QK9pArrW4RZtKZ/Qs57SCiR/+HrNiDduMtdu0Tcwr08XXYtUxWye7jZ5eqAx/
GchXaFp2tz3GqNkgFo2WO3ZUI/WehTTv7jC69hOI1atTJg09JSMsO/gttD6mQPW7r86qYAtyrGeb
v69BaDLsSfaJR6J11Uq8D7l5Fh+BhTnG99iGGwvLsrgndsCsJUUMMK8f9XH9ag065em1qkB1UYrz
MeZ/UxJx+YUhKKiwdNNcvl2Wrwpnmpgk9RmKCId1k0BvLEEpjQujorxehThqfThn0FzWRccXjv1G
7yC+fEmYe4BKn3kwnZA896wQRykfCZTFf/iturlxb5Ww5lcQYT6GE4QYo/OenV+X5AKl1yO4fCdc
1GE1osjHjav/flz4JKU+DzW6Y2dombEcQZEmUvSMo4GVwhLl6rFkkjmih7fgKgAwYBmGPJT/pNr2
kSoCzUOHy9O2ZLConGKEMDCZOAP8KFi9sFDT3Xgr2EvISeIRCGEfZ62PE/bBUWsP7SGdPmh+JWvl
6tpmc4wLbBw5PfyzJkXqQS9W5pyNohADkOkrj0W7GrfMoDlLrboJIoalEim6Qt63i53qzf8W/wvs
zBkJCtU9uVfVqblv2vRPpYSSw7//DFp/aOy6h+gX/jKaenSFJVUm/RXhckB4ySWz+es/zMY+nLtb
tYdATYfO7pzKpPweT9dWvcNMa8ZA/j/TJoOThxZA+174fXY+cIyPukNmDm5ep3oONrPy0lecqoAY
2wTuImYdw7nSCg2U3ekuGOjhxLs77urq580XjzSgtdqoCxPc2AqksapDsUFRxCqVuGhMKZRX/PHc
jNitiMa0GaIeAJcL2BbjW6cOMYBkPr3FUoumitwBUt0YvzmkW/iRxQ1vFmCRNgAZrMfrnllIHf/4
LD+b+1OKd5zl6vbGukKbzjBmUMEJyrUuE9m5qZaK+ZRt09rMm8ChJRnWuDBzzqK/gynSp92vLxr2
kCy7UK3hn4IIiwhls7UYFx1aWcbZTkZA8QneT8PjbvnlPtj9tXd+BIzGf4UTei2Cq1tmGrFAgu/m
KKebdQgNKbDyaT4Y9r5NPQX8uGwl6YnYfGVxsGI7UP9LtrvqbOgojNFBtmcXmiEeaoB0a/QnMc8Q
wtuj5HQ6Rh6lZNO6Gt2DpN65i4DSE+Z/o0UwSMaBPY/jw+7ZAXq2BC9bQltfYgV5vjEcui35EgN1
EViiMWjQlDMXYGeVUhYPAA9cBCzZgoSnS00+G3vKMUZWtLzbbGujz3kM30ixeODfGxnCMd0kDiF0
+3Gs+5102iglIwacCEm/ZqoCbLd8iiusjW1DDHBPpOxUK6bdXqZoq+WpqVQ1H2AoqOXy8nP0hoSZ
rK/4Ou2QNqofALvzwZ8oTWp1Juwvq3kdKL4sKtVzXgzVTAAubVug/bzkjCDukhOpTa8xfUJo2zPJ
Ly2P2MzpKb/yK8NT4mXTOkKi4Fd5NIfE0BkTJkoekI0oY8jAZCeETLeZ7glwoIuWY5HdV1NpTLAf
lcVyFAns19u+t166gk0zPQltRGRS745ASrqt4JWkPIuLAxCa2wogT/xz0V5S2/eD6pG3jyhs7fAC
ytzwnsHFCoEJTTKC/qwBlmcpkJnMWdoTy+E+46Xk3+/LpH9IZgFPxRj+9WQWz1HHIJTXfSvhsXVI
voKqGAuG5D0GFJkmmM01ExzrbzkpAMDMztB/FVb6RKHxBl3zBs/4uG4i/jmnMAZS8Co6le6Anu4K
Ew46OBoh85IqllC9I0+kmk0wrbiho76OyLi4kLbZgMvWbPyRw3P6Te7R6DhN/w/lDDs5PEqIpjh/
m3NreIXf65D8Ty1X3VLPw1qfFqqlwbUruaXtwJi2Ij45AIjx/dW80N60Rwsv6/J/+4ZsbJTqJRqt
f2tXIh1QCY3C1WPj/BlNeZV7TWt2r+nb/al47qPBLUZYOYn4OyhJ4+8fwYyrQFPH0tQ+n7pe17TS
ocHB2y+O44JXBEgjxW2vbqWkqM7uNOaDUVKP3ybJgg42NXtCVN9V7y65HTm7Pme2sw2eH+kH4DYa
ilmFoI3pTKOtJmX7Nzu3BgZvBL4Q+QIrmpNKIFF8HXn3ac9NpjG4rLMTAaUzuAcFNb/F2iJDF/bZ
oar/eALywoAVIUXR96ftj4LzgF6EwWntEjuW1CxlJ8/qBRAznBSaLFmssjJmTEZwLCgeObvixWA3
ec13mxXjyLBDFvAGz0WH9hH+OSCMO+waUMQA3VF6kipJWvrbuRNR2PqtZpvtatO9nrPDjVG83MeK
4GouGUhkp0Tbxt0ykouFZITSAGvOfF9zWginaHPhwIHUBFiZh0CLJrU57ffSgykS47iHoeONaVGo
nxSH0j9NcCApeJI1qypSTbg4mqNDPXaqCtR/9xbMPNlTJPkjzjlPfvWIqCKfZZSiDx4i3V9+gna1
eFBGE95nT9JuLnsryHHZLTp2QRiwFG1P+38ipFwifFpYooinMRgwxljleBM7aVkrhuZoGXl9+d1O
BEuwp9ODgCJzuSMHfOb6vE954jTc1TXJN3YSoLfLoQGkRUcrJQ+ADgGzvJfTgiQElyUYvrIenwPG
e15dBj6tn3H4GjBw/Xx/IJNW9DqGT3a6fT+iMx05h8ACK0o9Njl97y1iJfp714VAxSinEu5BPYML
8AkPfhYW30BNyJkGXAGJ0nDXx0g4pWZJhuMopy6kIhlE1+jGiD9vAnY8MBT7IdS359XjwnS4FtNN
aPjyYyfdsuX8Bt50oa+D22jEG+TJrIY/5QfWdICqDsv3sd/1Ehxp/rHqlgHExJPwI3W7wgFGNqeL
LX/fD1MOcQLvXAXpnU/Rcy7fJQ85ghb2mR45YUSMpEHrwUn/uno/YNcUGoWFjyFHtgKDofKH/6NQ
zPA+KGyDUBf1BDIBxEV/S6NYibrutCpcabr5lPNFnLywmAle40roiynnBvrFIQWSHg3pptqqQuVs
z/WXg2Ek8Uvbv4h2LonJbR08dSlDVrKNDa3qrRWEY06SNYNLLQm7ph3F3KPoii2B0Kxvf5bagM1d
fSCOnG0r5tp/8amVyL45zjcM4mQp+g3zvb2hBMZJG5gfFPIFcd8IyJizlljF+K/2BTWv4KS1mNKu
fZC48PXy8o4uISDmjAgokruXXaca5osiSyE+w1losvzarbWmQ8WeoukaHRDchiASQHvjxU6GZWUC
d78ePwCXHOdmq/rHMpB64YUMNFpa3cUzREogVhYQcFtZ/9JmW7y+jNgAlZVlgkbNCgbAQGf6YNrO
cilVwIgD7d/Zs1nae5oNgRBPeCd7BvVREduL0zILTYsOb5nqQHp1fZ0OFq//zV/ecJlQCjlQJ2Mj
0z1hUAuZBxfKM0ROvSH5zcohDFChK4I53g/DdqOfc/bePmEDyZikMaALF0PHN3LCD8mu6m954CVQ
8zaH54cV594vAeC31NCSWRrjL8db9zc+yq4ufMr3qvR69mmBYQ0TqsWANxDv/R0A3ImjTKGH1qFO
s1HDsf3BRCWQif6ulaq+01Isq/otyvbwwTk+DuzRHKHgxjrmQrEqLrF758t+UNpwROlsLekpRbh6
n00PFScJ82wIyLmkbxYXXfYEtWMyR9uRtmhnTeO7bH+3RVc5xmbXixZ7jeFRmGt2XgX/STuAxrgf
OGLUp2DMCK5jMib8uAKL+J2WwSehT1AJpAGcKHDrW4+OiZeVtUz9GXASTZn4jgoxcvLHwbUq6kRs
dLHb0/RJAdJbpYeyi9Em2k81Zk+JviN+jNS1qvkoNBdmvHsoRKB6HkXzEPe0y6LBPO+vVjKYdIqj
+e79HPnUuaPNqfWaIHVOLEDulItakrM8w6fWnvun62aKYr4CYVR6mqhtZYcrtp5eYFjwmw/LSa1A
yQkZl52Ld0ymvNnzFWQ9+ZPqcst60yjquldmymw30o+J9S5XRZ0KCG6GrcQYGS/yZoql4zG42n25
Bxzg/tsqD9yNk0xW1z3r3M4A8mynZchyDQpq1GuuA1h00XV9Xs6wti5pclu+uCATHP7eW+Y9WLX2
0TxsHPTVFV0QSxRN1OSUBWMG3SivCjhmRMPXpu23m15f8F60CbvYNqoTfLDKABq0e8V1ihE/nqnH
d+keGqP/dKwTzHlacGO0jJQcT/PTCGfWtfCLCn4AzUbNEFxmV0d8XAWD3yfbmNpboCW9SB8XHEHj
ByvPj4AfGfG+JGpKQSVoVdpy93ik1XtVWu8dz+HcXkOp9A6KGL6L1HNAsvMQmhdQtLcvyYwA8fgE
1sdLW4T8f9NI0LdBPFgSQ6WbAbkoCWOhGxib/ciDU91hKL9IYNFnTjN1V9rzTaDYe/jOhXG3TsQj
Lj3jr3UOUgf1NczwlANMpoAbBygAtaaB4ocXXZjO8ZxFly1iH6nZs6WFQwYIAmmjjR/jm80vvo4v
HnigBjj0F7A29nRo9spZG9eDcphoptLYRDIp/jq9li6drgpqvt4VWgL/WA8EpiStp0xLrlFab/fd
mveXGq53VvCMtGP681BCf5EmItQgxZP87gp+FlXlrIwXFsuAAqskwsJv2OjXW2UgJpx86mjmf9cS
vhC/3uyZfqY7bpQP2GVFYJYlyySoB+cf3BFbD6CZVKKJwSIm8a+/z3UkKdl3fW+QFwDZ6K3lLk3l
Nrne8UyQCtS6xM5y0gWJskGJFXeDuXKfH59o6G4TKz46pFEg8CCN9K6qNhsc7lGKf2n2pmZtSxFB
pCH7f/EU6uSDWfPPSNdHujMBF4xdMV+MST6sraLoxin9iC7P/hHjTBkruAam58wrd3QUmtyZKtEb
t6q//zB02x2Ddv7K4LqFBvCwrx6uDmr/tbNmww7DwPsF+xhAg5piDMdtN0DVynHdFKYgjxb+qBOY
gkJOHXemiKTfkg9QUocTwluEhah3LBbbvvXlQR+E/nm3GRGnpPMId6nR0rnZkmh8yHuDeTBpHGld
vEwaGY2+0ANg5cWF57QjqkK5ydCZlz4p4sT+INDycrfIhQQXCyzSO8W2CfcnUJqUhit9AorKEVaS
gWq4qLkhrzLfQJa0gzUGnc+OoVVIiGKEqjExhXTHU9GmW7KoRV4PmmfczzH97hiAJkU/rYb+f2Se
QLnmXWaqHCFBcuHQb9jczkQwcPfSsOvhnJM88UoSTXeJH15QGa7cTXt9c/hACC5+/3vyhsyJklSs
DDnAnH4+b6b8prOz5CjURkAFDLbgrToJYJD92MzvlXo40iucuB26GuziS6Hiru+1HDJXMPDp/f5H
lkGB0kEQ3Oi7G5oo5lK5cb0r/LmilP1FUNGcmqwse00uHc9A2ZBJ3nDTLKlN7TcKjZNOep4/kV/H
WiVo6ei0KQQ7F/kM0Blyzk2wrtONvQ0C5EyCxwnj3bQfGkEHAYE+GNbthFzovMUdzME0qlNushaJ
cXFklscEaxE95HH5JLww+HJBvMbMWDRlzMX76cAsGJRCo+wGomcKakgzuenldStnxj9sscvkvbSv
/1jZ26PPSsaDXHGPAHQV5Jnc4vs9xJ95jvDv3ctXMOEv7BUJ0Xi7PBxpPqO5l+nViCRDVigtUeVB
mAXWVEtWp/sVWboSQQSOmQSe2OlxRbKvAs0iOf9TVA7S8BK23oYlqyMjG3+qMUpr5Y6iBHsc3RQu
3cUVlNX7X3IGnd5RBs6vTddrAtsBk/9owhTRxtuPs69WRc2phMmFi+OpBHblNxKU6FQWjfOF01J4
mdqKFSUGz427JRSoraVOdj7UvzCbEyJpFYyvpyP9T7LAn1FJXcSyUAAF+ZkZaBaqpgG4TxJ30jHT
PiRU3FvuYCuR3RSPMXvmAvgso93j53gNTAKIIzmRVhfX/fOULn8LwRwzI+ozhc6p+xNObbjybGoF
jxdqWbBmt1zrykkVLTuv0+LGfVRn2DjT/1M8mXMsOjVh1iH4ZKMiEpW3BKwZDyGV8jg+b59uQKQN
ydjL64VgGrH1uMSb5uu9NAkfCxI2fFuAfpsVnv/0x+DWzN57L7FoMXkzXDps0MZ438Py5rELb3IG
qRAWyB0isMLKlaMWJtGnp7u9cZe3i74eHDSd08ASpNIWMZrO1+6/gFVYwnf27u/O+15GSPnu21zJ
GGTYPVW4v1l0flf8fMUL496DWwtqkA4xQToo0Ild8mxEr0Te9RReTuC+haKlnbOqNvIWL++ChQ5y
O5bqJlL52SkCiEv6a7NTCvpeovV9nTuqD59NNUG8FgPkk8BJTnQzYVQ70AE7urG3Fy9petXqug+V
NV411CuhWHZ50C9xwgffFTv7/sVHOgB2tm0BSPIY5GA/kQpPDxh03maVEUJd4bfbLR787+1u8D04
T2w7gKoTZ0MEueiGG/0XQteOmFhUwaQnCmFBWJy7e+BcDRZj161hBQV18VXx/ry2tw+H4B0+NYYM
c4xuve3OPwBZVV+y66YrFvmEBDawlOGWRi2Wpdu1SQnZe1NwgRzE2+FhrTbbejoXsFqgsCMJH0Fn
EE306wPAc1vz1EIQftZdpBE7DLRDBV7sHDt4Ca7vGHCozLp8bWWY4nfU1JefalYLA5+SijDdWOrj
dO9xOQMljEPP8DSsRslB8dq23S2csF6loyEPCDMQ06IJE/3CDEpM18dbI8+7/XqMJ1mYP9nqpbNz
JD8bXKZaBQn+CfRFGweAf9Lws84e6qhOXAZxTNZw100jVDM52MbkpTMkz6dysaUuL7okGvpbZibq
t9KmWr9Xu1JoNKaoQZ7JavfLp6mlecB05u+icc9Bl4yQRcTUNRc9I/q3QLTA5iEUMk4hGq0881Ft
oXfXOG9o22/FDDYCLzVABRZ1UmwVSb8rSiKSTTHjkHM0WNaT9grbb/igOOTnpzbW7EAWIUevZBNH
QWvT2vKf7ly4oAYXeGhVphg8WOsRM3TsehfvXA9EQstEHa+q02Vi7GUSeVMcQVAqH16J0t6q9YNj
+TOFmFQXMBr8JOcySN67CRpw7BmWptK6b60KNQdZkZq4tcxsYIgfV+3wrJm2ug76lHXLGwG4VNTY
CpKvR9B7sU8XH42oMibBcz6U9Si6gaKbRF2viLil69r8cNSp8eyZfejQu3aH0yaRuLwVpqbKT8DQ
mm3H2ZY3qpW9fShSybwVdKs0FCHH3AavAHEMwl80xYP+SKOJgnPGlxYd7/DzEhAXjBpjVMsNda1R
qIqtVHxoSp8YS61/yWVKPNY4paoYdTS5AGsWto7Kfa1N4Pd5JavQt2yLXfPiP+kmPPUky9F4hvRY
WWwPXHK9JYTML+VO5nH0Tc2Ze2OXzZYuPl+5LpYDHkrN7yG97NL/foRruBw2NXixenYaVrTiwx2v
hOBl7hEYXm5Hlfe0LCO1ceS8D4TpksTDBQnGzbL67Z5e+YFulnta3ryEEe7hjHfyfV+GBj0YGwQV
oRSCBe91NJL6W2/iO9LJT3k2ToMd2tg1a76iw+BUpj7f6jLVqjb5yAf6HyYoJwhE/jr8B5EbmCTn
IrOmqTQEEkh9unVZU9wMURFHcu01v0TLWYr3yDcqBZuYyTw5WphU9/rsIkaxN573Ws+3HPswmlYQ
q6xYsXRYelgsrzn3v6EsGCuPpLB0Q/TPp24wriIVukZVkETAsxHcvbWUqzwJltBfHy79h9f5Fhsn
VEN594vbVQusyN/IwC7gtYtoeLsGBx/pU0LVnki4dyherb8gk/XxyTKowiR5EPpBhHyRi3/orJC5
RnNx5cnNV0SZqDhaGxQPxm7ICW4q53qBtGKVogZ3nbwgvKH30mCD2qTpiq06T0ugG14Kz9WwsE85
dBgtrEYIRcn+FyUgvKRhdz2oeI5DtlRhGAYhDSyDfFzOPC82UoxZ/yBHnnC+dzi7yhKuHp3vX67I
GwjQKgd9ic+L5Ye++MiWxMpPnjq7lA05jf9vqNIhZ28Okcql0Xu21diZf6bidF6zmCox+ooCtvp5
rAVi2wxD9SGVffBcHazXeKd4pXPwH5UbGA8jz9CUHV0c57KxNxCR09sA8lY+w2TV4WrXPGlGqiA2
F7Y2I5MEDZrYBrLyASi3awezlxfRUJZ6pnqbi8WCYuNkJutifHtxm0PU77s1kgXGjr6X3gASSwrg
HIRpI0gXMU/P6LpV3PfVh3A67yFX9xXP4mctDiOoOmI7vBIIv2RiKO9lnrrjPHCDFMeEHkHda6MM
lE661ELIfBAJ6iHufte4+SCTtvGc5Cg00+7Tb7O/XUkTqZ60oRM1ZWWUVx36X8OMh0w5vv/0umxh
/HG448CwT4CRLuuj8BcRGKGOJangWC/sGOU+cWhamXgisFYd1/5wAnevlqVpOjGZ45Eoeg57FOVl
u38Bk7BMK1QexEzzm9jQjycUxNI1LHJH/KN7vcNGzqqjgKZq6B3iL3BwnwX9rfYSrW/Rv+hBPHEQ
8hzW4uZdYYJXwTavRWn4wYO6EnDUVPs4GyfFdHSLFWKV7KvX3z0nw+Rb9tFPhf1lHCpU5RLoqltW
rJSZ9SoKIO9zkmIiICs9Ep+y/1obvPUhtMFjl078c49OlV5jlTaUElJc1i1pu/xmGL8i7ehcHiHu
XRW1qS+wRPPUBtYur47KQBI8a0YGMOi1sayAJ8vG0+2UIuMXVPOlBFmnoI+6cL62WfZlNEBpfuL6
fvHp5001rC5eehGgD8fUcZ7FPC+xMpCnEePfzKd+kEQh0xOUfXdYBXaHziuBvVxfU70B4wzyg6Wu
D0EC2OrSpTE2/iW1O8sR0WHotr6XfquwO6s28oWuxVNGRfH0MOEchc46PTuLfMoyqD5SC+9g/qv2
w9A36kIs8Yymr3qYs7PtbjPUYHnXx0V9T/1sfvlBGrl0hpcZrNXfs6ePE9MdttS2zizXGH2D1Cdt
DYU6PMtt1K4xhiH4DgcQiu34L72XvEEnR2ovbm15IQkTlAihLje9z8BJZ2kXEU6pwIn4AYQ6BFIN
BFo2A07TqnFXgOxLFzdWkpJxULv4YLLANG0YL3G5m9JXeQl4byK1b+QewRNiiB7KB6+lZ3l8fmSm
fAdLaWwJGDdBHU7fTLOhP7+nKnd9czUyzXdO+F9383z1duEt0vrKmGk2gj2hjDgngOkHhz0A2f+F
5s0UoKSmDwPUDLav4YBQt7u4NTcHXnSYF8NVmkrQ6MaN83v/rLZbOO7jtfluHlJQHQhz8ba+nd3Q
Fs9mhmm2j10sBzWMZqdxzNdaPehIrRjax/ymmC87U4vQYv4kmzp2JYykQVaxqRZt946yfG9XVHtj
Tmc0PsS0wdAirfAYBA3hZQpchpfPJefmh4azHOYqo0Z5/7g+lLwo9gj83hPH2KKlYtCoRBogqteL
buhekwNAJtwwpTxAVQN6mofEORFnCT22lZzLHJ00Lq5uj14EtthFWC46lA3H4UM/7QwsocvXiwlI
+8ALWikDPBmUiupHLNqRek8d2mwve5EV6V4gXnxEIrsCg4x7/1/PIvSyMTg8YC/TvY9eP5aZB9Z3
plOl8zRz85GBNFcyV/feO14sWO/FzfQPixne/vHRBxm+TIhN1fjUkb+8sl2NBgTHxIcF1LDKm89W
AK6LV5SVxDSpDPJBERsJXuR0qdlDz/WxkEp99GFj5lmrOw1MnA1THnrm04egGOzuUXJly1snfO8w
MIEe6QePkcjSHuT/i/i7OYlL2meZBZEEjPrK795gxzpvPhkSIV7laEznOdM/uDDl/taPcwcFD+P4
EVfGAl/XQe/rjH7y8AhV8cbj1qTyPO/ZY3Dfy0IV+5AjIMlJY5xbK/76nhoa4pYwTJ4exzp4QCAF
xTQ3n+Pj9RxZ5tL8mproBMRbCjLVwXC94Xw9+XwJMlgryLfycAGBYgk1V9OriTfxk3kXWqS0ACNs
ePyLqFJF1ROq7HkkPj6SAyjh7Yeb6MpIDtFAEwQgpfUzDHN/aYX7Mu/0JVVclZOvysDDXNHQSnGO
AwTh1hoEH7f3i2FRGttL5m7se9kean62dLpWa3sZSXoKdFGAwIetlEB0P9mThNqt2jDP3fcA9Xzp
y07ALtGp+bkwvOJfadYhBfW8wp/9YYgSNGiDWj17j4OMjFc5QSJRch7UPYO9fTDUqRyVGRLlI+LJ
igf+SB5vg5fp/W3ZVWW4knh8pwMaSZoDiVPMjY9GnIJrQbB+PQe1cJRty92YhiHpjtieIOO5KtC3
RAcVC9ppajM1ZR6oqhc6YM7wVlv0xYwnw010u29Kc5Zhf4TqiZkbWBtgU06fPx1mwprUvBYrtD3T
21H1+/LCppNYjGwKuKktLgKZqZ6Y3vbFD8Lx9Hz3XE4BANPRmMdOWYmpEAMNsR+CVTcvBa3s7DbY
nCkdUfoi2dbUyHOhA3OhI0ni6Vt4VtH8EGn+8Q/h484hUNrVvd1ujPYr3cdKq0fdS26DchdQMXKG
t9ZXjP+v+wJ7DSNnS0HFRY2d45rdVoxDK8WRTqC5H+hlTRbnBuJPsl5AtpfobgfUE8MJxlDbpoOn
2P++xrmt0dNtLfuRD1SxSHNX2EORgmaQShcVi5WicXTh8n6RXOOA1vsezcbxXzgGlcVQ221RZFOm
xQcUP35F7CpEyznozmlcCkGZINlGz2/bw8dqtEga1C2LnfrwHniSihA0pXJTy3DW+AkTkkK2ZcW8
nnkwsGFoCm46ZQct21DBv5QpbFL701kC3NN+py1RQxNeBkLQlVcqBfO7nD2iqjYT1Bnq4yJdIYlq
KaRrb49ikusji0VqWnYqsPuDF0oaYK8KVv4s1aobsQGH296QDHUv9PJ9eOWq9+J+I/3S90yxNLWu
6TJK5becPfBPMM0PeBJOx1OWJQxTTojPYsElk93k9s6Bgiei7aG/o3ywcXVBHch3PYpEfvXh/+3y
llrvE0OQnRoGVlyNzzvO5wXLboG9/Rr4I/QWfI/L2yujoOam7j/9WBCEf8r34Ch7jivrDGXYy/1X
HVj0jtjQEHTqP7cw+G5pOpRIH/aE9w08CiLfP0XbIriLwNGLZ5Bv0i/d1VzchmgjF+UNDRAOvaFB
qr/4l4S+DDp7jLGCik60Y9WyZLSzBAWpwTxtU5os59LEHft/CWlmbtjiD8bOt6CcOQSkNaL3oVfo
ICCGcczyBM4AEIY45ULI79SGPbw9jgXOusVyhmBIa7VknsR267R2V81oLPsuuEgaqiT0gd2A66L6
lIbIWUe0nAlzsm/hdIDOnqXsG3Izx6A+HH51L2X9du+MjRJpKrscknmbaKe+rxj9ehbhiPsxjcr4
URfKSasFNk+IhKiJ39QR7bg0LzJhrW3UZGHvo8I8MxEfp06wBuaCXawgLranqxV4ECdrft6EqFMl
xOKyqLf3Q8cIFBQFgBxLOX18jBGNzKhWaygfPhkyFG9NyluPt8OL87uEamnrmN2kxVP+hX6BxsS5
8fAmngKJ0oFLXeFBSHHrrGlsBIslFfLQ1MVA8b+aYmUMARBooBpxfWsIzuTAonQrt/GEM+Uog4hS
rQm0UvWj3OQWXG5KajjQgvXaEIZQwe62Bg88kp3FEYWXS2GZwv1gRH/1zVkYOi0avtj2xxhZV/vU
/oBMstOAoTAAXqBMI1wtMkKXwNVY/KVagO3dkV7fCnHYrTG2lyact2qtyP2iGBN0Lf8UOEwT7W0t
NjO9v4DqZrVB38TlESigab0URE4arJi8Jy8Eeefypn8lUWQwb5V1jWE8UKxDP693NlL/DKCv0Ll8
Wegw1Za9ZGnduFcLXbzEsJmuJGeyvUMt4Vm5ABtx3cVMfr6pfNcOL+V6SoBP1kHMCFE+vcDxfvHG
K5ca5hDikowe4CFd0l0ZzyoA+xKPlV5vwgeiA4uhFaBmLja7/xJ2KsemHXJSlj+a95VAKS0n5m5/
rUnIvbVoNoXezRCcoPDKvwCqUtYeMAyaXCGvuICXk2LoKPuC64UZzPm05m1OfC2CbPnE5/+u/CMt
PR7+Y7NskZixd1zIYt2pwUYKbG4c3c7V0iruKZ7Q1bTCaP8qztBOkf9baLVYrO80wUYngHEP5iT2
icSRVwnX4IeTZgv5m1pE60Fombr66NFKRsZ8XCjCPPoVM6+IGdoddP50MEINKMcRwsKx0IXcUWs+
fQYlKfWjKQMqgvOaPvyrhiTPiGOJhFdog90ibV3FPx8XuSip19G0pMYjIC1PNQI/B7T0ZPDb2ybS
D6WX4GNMQVvvq8/wncw8ksqp2nBpzbhhyneXSDY/bTka7Jy5grJjOaqWNnFcE+Kqfl506zossIvP
w/9ld7XftjIvDpLGpbQFSYfFFEjhckxGa4zqy0G6nYT6EMHjSQo2UQ8PZyX79K67Xd4wc215USBO
83qGoniUETi/03509Wi1gEIWqhDC6XVJod4nDXQSOyIdk1J17eHCifZHv9T4ZUYA3hw8mGXNU3y5
JYMW1jFCRB87PVKbdrhag1d4FDdkTiSAD8QOGkmIIfuRPT+whioBM1ToVoAK2Oow8+OsMHN0aXLe
NLqj29QwOi/khjirxl1PbCj5a+E/joZGy5vA0DrFMTkaqHxcP5qYrfZT88xF6VNEqEu71RTaSGFP
OA+aGuIEWHXgDRMKoXm4XotTzhxmajv+EV1Q6Uqik3fCCX9IqNn7V5mj9XZOEX5M/95vH/O8X5VG
Seb51gofp5vrwIsb3nOnGiVZDGz+Fe3ByAyF5qzBelIYGXmlwBaEqh6RClLiuj89TII48tpuGTd/
V4PSwjYavcUHk6ZEBt4Pv1anQ1fLwv1f6IE9P1K005i+9rJytTfjkgBtHM+rTwl//H1l9Q92NJJl
TtghJy9Ti2vGoSg6FAI0E+ZhDf22yRgOF/lvAJIm3HLdaWL4bE48dyHuE64UBwoTWQPBltSFwCuw
EeolY6gMT7ND+5g75l4lNuKfqbARjlLWimCHBQ0Ir6jgUMZwNhDBW6X8yQdguGEar588gnZrgY6U
j/2UzVsyl/SCgZub1+cUhTO2NNFivSekUZI19H9oyGXaqQqO2xvpW1b8stWaY912NNxYKbvylMdu
LeydL2hMJtTede2nKNRghVenej1F6Uj1SOt02N3mcLPcwIPPiJIFEJdNQNQw0oX0uJCuu1lKx4rZ
vVOlH8uwhZkthRrD/O+HGFAndF0ZyH+Ms3S86Wyy2seXlpCDIKFFQsz6CZbKp33ig0fGYqrNLP5I
nxhBq4TvH31sDwkqPEfVtj0QuaY/CUIxoUgrIHf/+qvRLod3ChgaBmCwnRTyMMzcNmRlYeIeQfyM
DlUchHbmdg4idXzHUfOiH1X3cI8wQahnDSrdSQKu5lMmpBV5D9MUwb9bOaOQYYWNZKynDJ9Gw8f/
66owtMP8uRnm444TQevgYa8osrSi38gtT6oGrehifBnEhfxNHGokGQPQJKGqdbyk1jJoVNr0sAUo
ICChfZgAP4Vq/0f1ZlV0Z4Oz7CJmdGRtFYI8InvfY0Tk9VWTpr+AYYnMOSsIdn+xBJJ7hlesP2jG
8k0EjkuSK0sREs77s92uc46G3H2rP0LudCHZ+1xkT9qcR31b+kdhnIt/WYSHwZiqvIYONnVxmzFF
HuxYHwjAib/D4VbZ8Gh3dz/AkaTbyFuiNaGJyNcmoYUm8f3t+p3/DvMTM0sSkfkgYVVbYOYz0YRH
Xmz5XgQqqwadQuCKM+XZ/naDEl83HM3XTfrH31TAy+mTP2cIUKDV+qw2DNPedCVgVDgDbdbBMYgf
kprxVbXb5wlmrDHE3yCj36wAgrHXZ+fwXEP7hcwZPlQMyRLu1i2mMDcBmtYHkU4dSYNTGtUI8S3o
yMz0JaNra9H5cH2FJvMKrv1TYRMp/M68Nj1fNKaatAlfecHkNKc/rfnuCogWI6CkfHRyS2Gdo4pX
Om3+gfkbfHiY/S9io0f+jDjwuMZGsMkow+FlbuOBIb21dCF3U2hcTFIIFYuy3nud4PIFW/1oSl2X
Oz1NfnnlqhngMrq0WswAgCvZz1sUxTc5W0xkoVZAvbMTF3bOvkvIzHogp80QTjMfA3KDaPNqJmYb
F3g4Nk0XKWyuS9k+0KhpvItNG+jkQMHr2hk5nw0YcV7X0JI2PD+4+xKC9kkVfkiG9irgavNG5eDd
G9XT1m5GSEi9/UlJ6WzhABwt33uMVp3tWYuCABN8WW1MIRlSF4UjVKgJs3MNiDQksTZeoRpycxT8
AHTsSB7nL4sTFru3gdfr6mdHpIWvgIQnK5Clby5w+ahptfWXkLroi/6n85qVB8maBUtV59dyU5G9
5NRJv9QAvmdbcbPPrtWbMPtaaCcDKKV7HlbXBjfBvENCuHFHzDdgt5Wokfjnpkru7aV8cjsTUhJF
aW7NYh1NjX/pmsWnVGiFFCoZB7cfCPQf4wDw9GH4VdpLXmj3AdIl0jzcnHABLmKe76+ODhunU+3C
OMZgN0CD4qtgqoSnIHR0jkzNvqDaAxDKIzDvt+TWI+xk9AwWkhlVjAMcgvLIFfCPO5ne+qjmb15+
Yfla9iTc3MDSEHM3pPIbyfZylsvauxLm58+G6V371VAlKk0A1FE6orcNxxGd3q4gfLuvXo/mNzFK
7vfkYLsCcxrFxF7P22A3o55830HklwthdWtu2uNZYEzPkSnXDkNnWsjLepKKZ6a3E7xFGoVHJ7hl
M6V+nMOPLfj2dsYY6+mJ5yfz+ou2nxYNkYP2LbtVYi8Hsu6Ah1tPfrebFBZv6ETJUFgWedKMffY7
N49zC/yS/U4cb4z8sDqf3exVPNZc7VJPprBlD82BFTJdnjwZ1xSPQ5iSTGVIQDxW7XBJuvqzSdy/
get+QdOCSvWfLcVmwLXhHHQACo2qw13XYPpE6CfYG+K3U/VZUyJPf43Lt9tN2K9MPIT6xF6227rI
K4kf1rt4eIP44U3KIy1QNe/RKvYrlDrjulnE0LYOMGkvFeawvKdAfImL0KavU+2+3LBaryJHMmwB
PHUZD1Z4mXJEGybP2NADBNdZslI+NfgqMdeTRAmRjy/X6AyFXA9oleiX8Afz78+cDcsVrZQzZn+D
DuqHWCgleZFAvDCGPW/e3J+y+0GxPitLnX2K/UuBbdculCiStqfVOgG8MIBe0vke2z7MUxUTYKEq
//UgsEHJiWI/1bBWedgJLMxBR1IOccPXJPSEDkBYQ+CoLi0sI1S/8fsx9fJS01SLa8Jnqc11HU7w
zyR77PYeFbQe5aKTJr310ESjE41qtRhaC0S2GtZfdXGOjEGQA4tZHyApi+XeHQuVhFAAW/wNJiST
vdF1di8oV0vtui3JjRbRSYKhbtNWmm1WYFX+SqPyUxWXyeusmzfNYl0lLK1teoxZIZwuoZl+ARyu
A46kxdvElET5WivkUUiqrDBfQSfsHOzS7Chh95dzd5FN6IkZXPYhqz+Pc7t5Ypddi3edcR5V1T0b
+xHp6Js4d5lDkvQqc+8Nf/i6yO5zB3Ht5NbIjGBLaqRbn2G7bIxiynq8u4uDLc7EoRp4KA9Mi5DO
PRfrBCpP+j21GPguyQWkhfuUWJR6xgIsPc4Z8ogD7TrIiNpM4C5y5h3fYeF1y38Qh9F5Z2PIJjAx
8flWH4ZEf3N4dCL/kZKMbED2MSu4H/pFAyNouR+ANWnftqy9iR6gNcFgPOr3dhfWop735gt3PfCo
f1h3y23U6bAytwQ8FBriKHACWkAzUOoo4HsftvYV+MaSxPoaJmFwltsjY4skmtzRFbw2drz5bwcW
ZVakufTBaXIKHgzFtBA641LIHsanqdj+KERxyFniIniCi7AGGS3mlzY1LJMd9mMDXDY14LvOlz8M
BA76LPtp++vosMEE/ohPwvdi4FSjBv3S5J5jVhujMlpexj5BeioVCAFJG5Z3+l+N81xxmnC6VL7h
po7mk6T7qg7mpdR9A+tHHRfEwkderctSk+SuDiBWf8W6NEr0eID3ZTWMvQsWcHdokxO6UzgIgII9
7y8z3BwjpjPpwfOkZ3KE9zDZwunrsqaZotEpOUD/qcjo+sc1xizdOtsX2xJgt6u7LJ+octx7sMiK
t738Bk1n/+xZnmxS8QbwL4BoKu1F+wcvBdFgqDRykbD/on92pNMyKma8d4yZz7UVp+YBGGiuu1f3
Sc2mkk0O4sxTuMSuZ3NgmchPGayEjMAxSDBtc3sIBfVSlwKDcTjVafkWHM2cRTI+cgk+pgiQlxNP
VyJA6B9v3nYyLs6a5OnDggcsnaRnd1bXzPsCiQKQFk36U+oGMXAcUqXqih5083h/ml0K1AtI42o0
HvQdGmZAz2QvW1RBCvop89DZsXfC2vBq5CdheF7reStNrWlf9xxZGBBwNe4YVwvZ8bHXGmRdCNqh
oo/3iCse68fbdLvrWxiTdXZucw3evyxrpNUpIo4nROrBbHFB69tKSEG8Ax3btUkK/8S9eCK1WcnN
yyxtP2IANt8AicJEpzdYZxHHV1La6V04i3bwFBbTnRcH5LXHLVUVPUxKLy9O505owyvFEwvMtPI9
dlmzHDlUHDKgu7KB94+Cy7UOfVkhLCY0hdLfYU2uL/3JG842y4ZRgl8m2h2zKGVf2hjhv2AsCFqG
m/n052njb7PvM2XJkRGXtBoc9sH+x8gUCKRnYbEoCDcVPymQ9LyuDbrBnXjh0HNWuMHz3J65bQ3q
FJf+e2IaSuX/SJngjaZyeimeWuQmkjCUMFjtgsNzcdbmTFw/rm+cSk/TEZ1kExPwJfypqklCfS7o
EPUOXjXAV+Xdhk2yjVeyIwVzrekOPlrr4eYstfQ0gynyOEdcCKWhllcz48GoGYqvag3pH8yUNFcu
Lu4Hs133kAGWR3t+duGYf+KsaRuFehpEmXKOIFRNt6F4Q5CLjhvLwYGjHRZU2j9zv4onEPPqG2Hx
bFEFrbEGlnp+G4ZfRqkDIX/jTzwS4a1eZVaR54yAPybNMEeRHupb/EalvwUsqH+M7Abeg/G/vCTW
WUSvbBB8O/IXvI9wEMq6/C28mve3WxannZbcCoIixqpJ06veETv+PCdPOG20BZWDoeCOjyU/EwNG
sgdnvy+2zIbw6bMBVH4wqOv4HV2QgRvA8noFn3UhvuXj69mfDhnTtQWjLA2i7ddRjVKuiPF18CYr
0QD45Ye0Yqyg7VrnE7/YXEUgDNDXSGgLgMf24QsqAondBSbi9lCGeptdUaSn/WU8+difRcRIy0EK
bOBZyzFl7mXCrfl7rsR28z6JHZ+odgIG1cyOrB8//cgnsXhUX6EWj6sUf+5zdNZZ6F+nofo7LEfv
4+MoCCOUkomRCc+6PoNXViiF1a+GDXPtFuESSb/iImqR5eA+LRRoUssdy9h8fg16kyJOY0hodqd7
DJV39lFcJGxY/++06LR1X/ahlR0gKq25CYD9JpGrfv2l3/2PEcnjtun14j2qnqS2Tn4Dt5Wf3lxo
wALcjgN6edXKYExxL99aPEcNcTRuN80dgEfZocYj2JubEgQUOriCekSw6ntLiJQOIBhyA/Qk479/
yw3/Ye2hfQlriTev/bRcjFyYUgN3yfaci522Al2UJvFOEFLudvdy/xCbX/ngqHOYa4J5+Biyka8q
sKelh/Z2ZE0BR72V8xDN/MUWM4XMXwMW0/7pKkBOASZMIpR2cvh92arYmFrp53yl1C7z1+IjmyZ8
5xiUjG/bi4XFUXGaK2UX6aOsaobFABC0XT6/5iSBdXaix1B4CvvmDR110iQL2TtirqgZ7Gipqp41
l1pUaubTJb8zvVdrZbT14ibFC0MTWgpX+ocoqsw2fohe3p5ckQqry+D7UFJd/sjpDkxkDJUNp7ix
mxhc1p9VpdcBCNAe5CgLCusgHwwTUrrCtjD8X83Pn5inKXSyld1pB9GsaArQ6HFlC1kHDat46prn
Xhu6nKsVolscf/6Lfe7yGN8P+EJA9n/1waJhReB2obqJHNTEcnuAcMry3LHQ2IwA+hql99deudV8
Xy0uuGBZNyojSY7Sv4oOp2zeRuYNYeshEzPlEiJHxLxQlD4whpJj7ChAJJdgcRsF8PhSgUOwBG3p
UMjiSaU9/xg7a5vQlZ+hLArtM0EOokpC08SgD+erEQjbkuZQe02/3p46o8t7RkqVwJVfpghCKb+Y
FLr+tD9Z/5eijpkYWvoyZ96lzDuD6v/3fQcyHS9N3dDziRDhN1cwS2LLBq9MIDJqKNkNpy30qesA
26aafWAVQ1UM1iAl5al10xJPGNffjFPKId+Yk7UqXIQGWZ4NYtoL/bYhGQLjbwgrcTRBnMA1nGuD
pDfqhmYsEFgVPfh9wftZSgQB0JYSiRqPy3skL4L+iUMwKc5tCKfssat3NB8YcRznn4dUSIQbXBuv
XF6tdZRB88QQUw+MAHv+QX8cw4qX05vlyiA4uGQRyZb2L1Op6h0u+C9Sizdwq1NA7htOcwqPJO6D
2BE1ylvhlBbau+GNPGAASvP0jbdUwwZCiseJvhzt3PljduBAfKEzu8/kwrGQjhFPmYWpugSy1/G3
AH33srZ1daG4WXrKnZAmYoDzRlssKJdy7Pr+0KQqEVZ6+BpB9Jc1MCD3wQduvwoko/rakd9Yv9lM
5V/nti+arNXGmyzagv3/cp8D8QiNJkWgZvMEKTDuAD8hqDQxUzTGhlzOBlSX5JfHN9HZsgyjjkh0
3QKEryaiiFc/Bw3lutJWMIbZyO0dncyAYeL1RyiLKuiQDFR5gcYZwIi+W0hAKPaHT1nzpeSiPu+0
HPKKriJIasfGUjT29k5tqXX+x3tzdhpDuIBfRSGiR3GezP7ALMYXvY8VQRW7YHoQaa4fD4jTpUbL
tjFbIyYEkUWT7oh0OoIPUJZP1o5QmjujiiJLEpC0a43PitCFxwLr/AhcK5VipK3y9puDH5iyNgLN
zLr/x39rElE4BEdF+/Jvv1UcE4/8wPT9KeLqpSVZOHgRh3EcplLhS35Tzk/wC41i1dLTo8hNVuXZ
1Ei988rNzakQDOMC1bA1sTe/0IMtPA7eWmYqy57aaRzHzfk4ptHTy5sj6DUtpXCxhtcjgJu7cTYe
dWUtnidZZPINmO4aLifkvwWwkKfo2duqR9I3qncmtaMm2/YZBbcF6FNFV3ZuU+yTzRuIKn5E0DnU
v/IfY9pUZnfgCVKLmoXQnz+QS4jcSpDo5WN9GKWnAy9y3lsGYh8/2XNYIFMPaNHYiBZ3pjhvOZg7
+h3MVCwqjHZOhx13HfPI57hnrmn2tTvW5z6Pb+DiSBEVetsygcANrhN5MJw6rJaHbZh5IM+dTwb2
ePU1oSfqVKg2henenfMU/CPziagSyN0onAf6u1IkJX0tX7NwvWJWSq00QCfmPRr81aBTjIa329WP
oaStcDoJagg31fbq4lHY7GU1ZvZP74T0lf0zGJe2C38BkhoFStNZ+CpDypOHUoQJytcDmUGxPtjW
p/mSTd0DmPldH80NMqKPZfMjEUuVMbg4BIns5z8yXwMamlrdfu7xmSo0PTcX+zwGHVRSc/N0hZpa
kNhzBss5sLmRoJMM61wj4BfaY8DlpMUD/SqIB80NneTFKbyG5+bZak6iQcyuvi8pTgqnrzEpX1ez
4diIdxnLVCsifib3YcaE8m6sEf1R/7Kt/dLfM1OI2P3dWhw+uRGm7Qau+uPzfhp3K04qfQWXiORS
BUuqVY+yvougvm+ufF8KyPlIxaNhB6cDfkC4znk442+hGICUqqaJPPVajiBTi/WH6vS8Qb9Y5ocq
Qb7aUZm4XKaUhQMK7sInmjxgtQ2Ty1bNzWoxiLYYmxLmCRyWJSbnzLPIeRgggit4vKyq+dPnmTo+
VknIzEqfKDAIwzVMz4AeGJWQB9W0tAs8jmf+SJsLIkyzmCtu+cJmeRbYLLGvvn0bz4FhJ3Z9sfLB
mGZKsJSrM+7esLPhl/aCuxE/YLiN2x66hYQBI9AP8dWteb9McqfsFwCpbtT5CdzNFIYtOmMeaOUb
u7mhvVzFPTqzom5hWSbw8Y5Qdy1Wm2oJTlDASXF35Wuu0MEwqkHH8Y6wMRa5us1CR73Vuqmv2a6a
kLfhneKdwUs/LELX2LLwU/59gjNyhHXHYbqzuU18Wzy25XwgW9O0tqMVPOtPnWZDtfhoREea02/O
h5nAwYz2Gl7o7/uFV2pMkOKvgWxh9aqQFmCt4VC6nc/DfVMXKPtw713rWLUjMVOWX7YownDvSn2l
CLOk0AhogXV9KSX8YLD1LKG3Y4/9dbcEmKn37dpy0IaVNdBFXwgWPXz2g9F9ASU+GxhoS51vmigm
NqIU081CjsaII4wDgOawqA4f5URNg0FQifDC1zyIyEMS7b9lbx7Mi0IKvN6V/6TKGB7f/JA4ETaA
5ycaG2bupYd6/na3Fi3criRVfMHsTeX8ymkAZcGsNUwfyQ6kbyuXD+j6c5zOgEQ+NzFkFUBezaG1
ACUphZuBdmMYdhLUCK7+vMp0VpSjdBrguJSS9ioxRZrugsZEnL1ZojcHT3OUAEKgE5OUdS2HDHA9
h5eGW0pRZiq3/YrTmgDUKmaxNBnQorImO4Jy9uFteldo5ZBGujJN06CLp15LAHT7CWceusan9gOD
/XSEI06P5+b+m/KpGrdkftojqLcrsLEcQOTEFmRDrqMDDcchD+f9X0XaCQwjI3IhLin0NTU8vgyL
eags9PeyntBQyW8wWxSrj+i7NUy+YB2/A+EUCNB6wLexKSOyy0Ft8EQKNWTeOc81e3JkW0uGNhF+
VZiZR5nBDGGv50lFj/Olal35cKCmDDPp1r3Owh44d7vAHXqyiEREwgWS0IO7S395mgEQkOWxAcKw
tzv7oc3lBOWjxsjjr+yxw1+yNyz8dmJRGyNiaffqvHocxBHKJ8JhNmmeYrvhSPM4Ct+UMI6bSlZ9
DVnX0c1b81wBuH/zZnLPS0Jc+zsMFpHte22GTKzcGprD8f5p3CZIdfnNuXwv3y758VUe806VzL0F
sX2fDml13V1L8mZvQlK9dMBzfvmXQmFD4eDThNqqayTL0KlplHcBO5TVkNPnu/5cz5cxuRNle8/v
HnCH3vlWZvzBeJPpyclZU9iQpNMUDcokR2ULePI3R0VmmruZf6pbhKEKWQl40YmbQTiUqwOeidY3
4bN5ZOy67CcOH356AGCpr9iZ8cn5OIu8TefKxLmMTfKVrEykpdSB1GCxMtQdPw4t5xqRd5b9bRr+
kGQu+XhMJ8ydKn76yeQHSw/yWezzCkhYEA0PsGEwVZIO0cFo5S7ZReq6/KYQeGpjgSngQ2ok9GOy
Fbfrhb0mz862fmZ1PFIw1XhtuffIxLwa2h5E47vHaoJzdXmyJXflMMp4WWDWI1+p0mkFWY5p2xpe
H6R9bOAq3b9Spd2NqDbSjA5FlS9t2xX4DWDyLg5Li4XVIRgSBbLgI2L11xPD/iTJu+l94Sju9C2p
OdQXQEdQ7P0SCw11eB7elAm4ZkUk/xG08NDF7ix5p/0Q91VFdnWrdySVBj89vu306lIrOxHgUjxw
cBi9dxq1RHpsrXQS66qhBUGG0xSijkvTmJnTIiUU0NIisLsOa2OD6tdmCIwZQM64XtXm3MIK6d5q
yvvDdcldn/Ee47eZBeFucDEbggwVKeM5RJWaUdJ6HlaB4xuKS9BcCUVVpg3ufCyeXhqMR6xsQdZ6
ycJ8NYyVteFFBa//GvB1Sn/3zQnKwmkjYHZa+sxETzyFo5Eo2H3u0wGyDQls9ZKuA2n00PPMsPfq
HP3p2GqiD2AvT3f4nBlQSLynHqWsu4f0Sp5+aEWT1g3HLT5qRMIqlzmh4nCKLNhaUyKem5ZGqXKp
V8/RoYJ5dI/9Q+hJsFjXmBiTXe/3DxswhVrc3fMs8ONSYLgM+NPvQI1xJ+ME7TdCgSLlUATfgFEb
KrwD41E4Pjfip+C6x4qQwJ/6+6lsEGQou/ydJroKjVvaZ45EXirsdGtCp3UrLiO7+ZiUwtwlHXZL
oBdHidu9xFxo4Od+Ug7u3b756KL7hXHHyqqboGHd/GQDznxDdcnMSbvaWJkuy+cEp71sCKP3zt04
xZGKZmbGs93s3jbRt9zCFgZkkxta0fcMmQk326B6cfPeBVsfDYHuhKq/UX4NM64WZp3xmRvCLwwU
Q8bXjiEmwZZOUv3cBVo72tl4iYQYZ4fLUrQVZ4ggbsxVjbgZJvQ6XT9j2I/XZ8iyGAfDwKLkjCY4
PTF6YeIRAt+HauCTsYf3lqC3RLp+rz4WbaKpxe2X9yNCUP2H0GNO5L8XCIrjlf80tSv3I46xUkoy
rChhOyKlLnWRf+LlQputo0GRUXrJqiy83W8I9GiclrCfuuSkApiLVlKTg0R8hmONRyjZda4gm3TY
gvDgLeokqECCbDf7ZHoNzYAlQq5CO9J1zlzs+LDVB/TNHYYZekthnIeIGZ4ykxea63RaA0oORS+u
9k53Rl8JVulSnl27mesN6zfOJpv7Hu+K74/R6+Xz60IH4Q9TEoudlcXLqjxHoj7mbb06J2xjdJak
OpHN+75gwNOSTj5lXqVCQ5PyF+z9J2PXaZyh0OiXcezjDMrC4pSPQ7qCjEt83ANxmfFInEVnmKcy
2BWd8QPnpOCxPrizCy4Ezm1pqRKJlIUq/BcW/gqBvkpyp9lt+7RJ5IJDRPgpxqbvL2SATDio3rEC
o47UQx8T1sbGHZgOTmKe84JkOqe8z9iIJHp+rQyqf0x0o1OMcLHpU6YJgLZClcQgfkgYBjiXeL1S
HOCYOzOhkwc0gqtYH34oufdWyUrbRBd8Mp/ADgOvWPyc2rfWCv891ZFZaWGLWS2pAA/tyZZhKO8P
rGzjj3B+QF88kWJUzspFUC/cQA7zU3j2JTGzlD227PRQwIuZz0zebTSCr2HbGhYav4SRGSRx5Cww
rxJ+KPqR+x8Uah/mRMvxMpjbYRHdn+u/vRS+4C08rc6BffKu4w5sfAMUGdVGdbHYRBL7K+ASidRc
rY8syr1dyrRV5Cfq4Xwqcy60Ljk7o+YC2GHGuFgxJVqJhqf+XBg/SEhhs88MAEaKhsl0Jjvy8e2D
k1wFpMsP81HLjPvRMQydSoJ7kf88Qh1lMGTioWm8WQPlFp0Jh9gQhIXnSVD7+Bwhue6TXFrgpZl7
hy6lhS1018aCJjXqi635wEWmC+T23M0PhJK+w0F9DBRnZr7zsEcj3CJiIAUnA/znMNTidSnc7CJC
1ELg8Ikz/hBwv8/VhNMe53yfFSdOo1AMsE8Dc0EX023gWQcnEtY+IAueEUeLgifvQET/jsooHb/V
k69XTBjHwkr57kB0AtRYAl8hcVnHthTlG8t4Op+qNL2BFH0GTRzANPqPGHSYoGPnmCrpdjmRVPfa
vHhNbf8oXJF8iNCr7vNYuNaX5oLbWkQhmv1AqhHjor/NaZLWwL9ZYaiBIg19PudaCsxlaXpLiaB9
0WqcwLhvhAIqBKaJUKFVbZO3yx24wZ9QU6v4YNCbCiocdyvS6jkFy4YG5xg4S7j5R+qi1IY/dK1K
PTEQ+uXZtKe89usdfdOp/AjXiX0kvc6EUw6WmtwrVpCuTQMUf6GATtXalSnQ7vwH75m5vv6RFBV0
2go21QjKUQPWM6iYMYo46qmjmWHLaIamZ6B0GO0CJcsAxbp5F2LNrq66/gZOME+fSmtMO6EUWyUZ
EThJIL2qxVT/QY7lvhAFuKSqIZAHK03FklblBGSvK3FYxTkWm2GhsQbGZgo29vFIE2NFs0EOr5Fc
ew4qoa1DsHHSYZ5M0SSf52SIRnGsrsxx4zjtMjZsqBMLv1jEeMARLlOpZEUYiPHfPVqQkCIHrTV1
f8iLM0B8DbgDAdNLx0Q238Rl1fNkR3dj3zVnNVsV4MCUkY0jgcCbTQSBPwN3PFWEuSWm1T7xVvFN
QDRx2YyCLS+F+tNSA2Zwfe2Slwf9ATD0QJw0yIZ1z/fWTR0O9I8wRbLIGCWCqlhVCggNBZuFU7Yo
uaa0iBA9qlfEkT1VYU7RsI2kyxn0fbdQdcMtYBS+ZgA9zdw4Wjl0u6kzfqvSbKwKeugI13v1QTOe
5GxI7iInras5fU3qeFg/wSLQ2Yc/0JrXj1vMSD9nqdrJfcwvKbmSYh9cvj1b4kKfl/UKyesABDBS
R9mJv7lbeI4pES93WIjc3gx6s1DZjo3rgPcU/ale4SyUImEzAM+twQKGXW9UllCdO3JpphsPlXct
kKSlFy2UubBtB3mZzWJ/uJ2yYtHOSmCdtnYNKyFGGfagrzqv1wkghrblcC3JzS2GNLvRKe+IppmU
EPMBFmwuWXy6SynQqCVaR85644a7QJrD2MmeOMjLWmAMm6WBtyfJyRqxyTGoh0+gcNGimNV1XX+B
ggrhnDqstv7uWvs3yGYkeEXCgcRSvxgJG+BPGCUETquNBBUxJSp+F4XaJkrIYogLiIWlwJSEPPhk
ag8ZdHv2WGXEOwujLuayuDAKTdt/M5vxAB4pILvXb2m6il2HVtOxJBo2N1Yt7RKvRtgG06R06TEx
C7RqlABqawJEpEjy8V+rCKm1lhYl0jMYlm+MZ/cwrkyMlV71skilrwf6vuyh82pWiTSUEXkQrSxN
TRVrZpQoadgSioPjTBx0ATsSZ5sWNsLkqOns24Mdttk1a6KQ3h369KKDc6oS9uindcbgknGdiHDa
zyKIyx2av0PJ19qR/82EOmMnQ031CFhMYKZzmCaDQCLlLTeqeoSachJGxLDmuSTM5xzNeuwM0NqV
ziEfCVOGLNvnLh3eqGXBOMo8a44pknQg21FTm84lxKjkPAWY76I+wqB/5ZaUdgq01SjBrqXvaTW9
lky1Sl5L8OJA8iHpRSQJL1Zaj8MqeAFSZEVYscKKm0+EYZh3FuzrvD3XxaPHD/WKUP/zhCRWWNp+
zFU5dTyjPm9/b2JYVxYybfeES58MXPlt0dtYn07serwQmVcCMSZxCHdZnfh9VDEddp6QMmXcR34+
8s3FqGycUAyygDRUFuTJ0aWRIme23PTs1oHX3B5/kZlnNQ383adjwTwwlOpLcu37znNQh1GzwFlN
+QhDRvuLN0IJDiVxyQ+8xTNvpbGzBmYub4rF7szXFRjslrWNfO6+TpciYiv5lr5UsIH8fu/20tRI
CK5/kpN/jsKlV48aOQlF3L4V04uQQjb9LRRDD8SS7Phf2j5evVI9oS+8fmT3f/DKkvHMoKMvWdYK
w3d8yktZyiDhYlJNHLRSE1so5UlvEMlglIbiWzHuyd2NrDt+VcnmkXt8qKwNYfXHmnUGXAireDa4
6p1HHHOI6x+yVWhJH0bL6Uwej+mxMhboFdw9XZxwYz6j4U6I5TESAHGgMnKYtHYJlcZcUM0X9F67
Kb3vPNOrS7pfmHeddPVcIl9PWxvdNTjEMs2UmnKi+Bkee+I/m6lNz9W0NpgQDtEcZAvQk7gSqFpK
rSDrXvL7ma/ZGhx8oYDAWPqKhET4DEJbvW2H4TG46vqsvdDgriVm4m3I2p/Cs1fPYWfcjY2dm1W9
BuJ5Vbl6d0dIBVbMFpvdZKAUVzl+rruXE47n9JjhsN22ohTxWFzV/zy15lMvkH5Fwt8GwBQCuxGb
UcwvQgQoU1zB8x97jYKk6O5StHSz7tmKYXRU8F0bKcPrKAmOSy/5ZFScDzLmobmcRdofzbCzKc5l
llGfyFo3BfJRMs0W2bofmEaiHy1cbpMW8d7muf5Hp7uWDVSEydJWt2wqpmBwNtHLG8gmYOd2NWKZ
4OWZiUY/9qwBbeX3FG1aoetptCi3emH1tslgXUinmfuP5wc4XFEgIe7gYtGT/cRmJdAl0XS5KJzO
1eWMwlXTYfMOGBQE+MjEuXCrzwC7QQ0NEdhFkBYm9IR1f0bav6hYMAnVcki5J22WZGhmQzwbbOaA
qqV9vcISmgEGJEkAJz4CepxnImoCOcH7rHmnt9nWoywohN8yHm8abs0jSZikiLD76jNyjjkS4PsI
gFlU4uT93oeiog8p3twLaZOIS7drDHzP5a2X2T6yRDGllIj1ZLLJyBP26x82miUE4zYLhY23OsAC
i0i5jckisuBdaetgGTPtttEo/aG8N8WCeRqx6QRL4Zsmia8c1Bn2qvs2XEEkxgrwS6JmVdH8rE8s
HdcTRmpmHpTtgippB72NmQefboOt1gYkDbHHXkyC4Wenxp9+8nQTV7fmS84dsk4E45IEicOSXAIP
wfImhu+I18byGzhppt2upn1MRN7BtaeNd5ANvSQ/PJUPUVvpIeAhqrjNUrkxXSjQgnCEwILyMRAE
uSCINNxRidMqsjT7bnwr0H8L0mdpbkt4GoGtGMHk8Whj214i3733pqjzRv95R3HFa/HaPv77RNpp
YqszkqDWJFCoNL208QBIuDqnNrqrBeB9FSTJjXAwEYulz5LZ1ORoiHuKRGqNsHxOTA+sCXOqEcmd
1zE+Y9UzL2Wz1zZnhOlT9gELS0GmrhIgRzOkD1a1rSVsV7V58YPk8uRXRj8fz8E4sQbkz5k52DrT
rtDMdGluHR/w9j7qYg/kHpIp3yMU2gssOIl6Sq/rbyuDdzQpga8sckBs19bHlShL/YBknsITTHeB
U/EsTrkGmTyE8s37JVDMA38VJmF19DyPIsWyDjJRPCT70EaHSRycBZsHhUP5q2255MGR3kY949KA
DBjOJcSotL00kDNUbTz9h2q2MuW3umre3Lds0A+Ca9UTuE+WYoZF3IMjxcAfb3TcOGus6TuPSrA4
bhG0R6S9bJ0t1suerInonBErwm2cXQukWRRFHTsXMxRdXeU8Oj7X9d/HH87SIUep4PKGaFTdiVZ7
8chTBFC5rVkS38X3w4NPlTFekvESFlIGbhSTiYaSNzHENLi1SuUJgMnX6GE18NdeVwxc6FVJWFwx
jmijO5B8XbUBL0e6elSW/yRNPPWUX67qz+6k15gHRV1jVtV0HKlEabkweyyRoVHs0XNOT0CtEAZk
3uqACd4rzB3yeOqnCzRjP2p9/KxVj4yFAJzgQSgK9Nr0pBlLDRpI1wtgcpgB6xoydlWM0lP7vmJ7
qghq/H/zugA3mw2Y3sPBluMJLWb2nEFJdajNjEp6o2Qn+tA5JYSOq2S51L7K3GT5hvWiN7NpPAgj
MPBIE97XYxlR2VNhd9da2CzFYJhSluY8C5J/7gQI5AmNG0bagKQjLBVirKjzp19steOw+jTBygrM
Audn5b0pZ+GrIHDDzrjko6KshfSjNXWE+KIqJTdDxw7AbXAnu+iM5nW+KHoSfkXS63/lNA24A9vk
V/5VBe2eyeg7D8gOoBLEmvSmuTCsEWW/WHFN0CM/jNvE0SNTAAycOocGdj3/x97s61/JnJ0M98Oy
xQzSl9LfnZ2CxlJF5unnvJADlxNoJacMZ6Vozwu6mE6nMhSGtMoXPCIjMyVZN6MXKJmwdQHS9tD+
9pcR/K6x/ETzIb3bMRgXhzQVmf0DqLw52I1PGIkqHWLFWikYjJeE1WI/Q6FzjZ4YrvLNRe+lzWSG
9U6w0CqwxtlTYZNJHToE8WZH6beqP55cnbkhHQlr1ECYFoqM98b64si2rcpdLo1RQ0M1TpWXZFkH
YAFFma0ZwXoMNgeo6nbfYg0MwiRv5F1zvNC5YNQtF8+1U7CNLPuN9Ux6AdWFXuzvLLvnrJ6lr9fq
5HNVr7t7GMj9tE9ZxWdak8N9QzKs0s7xZe+LkXU6/FI94BqQYge1f0aF4SEvjOHdyS6hp5IBoJtp
KCC5wDJLBzBqkDWGLqedGwBF3eEjcAfMR0aVb4bv3R6mBAqVNog06VkUgPmYJQMKNV8LY7cmXK4j
IXy+RBVfwPHYTKv75kM2ePB+8zkw/4r5vWL9ZnOhV53UWu5y2/mH1YzDAGGfrI4Bdr1adHilwxOU
2sxMaRxRRAv8MG6KhYMKnsYJE6TQ3WQ6+KsQEBG2XksLPCRZSVhHH+cWjrbuPTIlLfIxEuQCGgof
Zs/rD97LQMnRg0JiDn1LgNf3fzmNuw3V+jtd2snq6ZQqPR+eCJ0IEJ41Odlsk+OeBR/NQjPgp7j7
HbB5YK9flvdmMbC8dUVQqxsGpUBsgMM63Lq5/4Jq1xPfBj59+hRDv1UG9eIo9RiTxYtHYp4KFx9M
7RY742a97FleM1BWPh1RhwtGeeOA/D1f0jLCkHrOG4Q2O1S6KRCyavnFvPHPP6p+zvadUWlw5Jtt
IxmBwJRPoO53tY6JGn6uRVmy97x3pKSbTPIROaCKxUiLFJI39gfcjW3daD58fTbugm5bz7uITRQp
IKTqGTCx2V4/sL3PyQ0as5boYqQ0Fs6HOkqliy8tl5VNacBpz44MwxIrRYvpKgucTzAOYkBUv1m7
SAt4tcHzZxtEg9kqAY0QsMEz8gopUmz0l1z/E0lzLgPOfkq/kcUaKJS7u0ScDb5JPLOjRruVVQgL
DoKMPyhaHUbo/BG25FCF2pNRn2olwBC7a+ziiCUt5JL5uVi88H/VQwSd/stQ/B7ICpDU5UePJWmN
ojhGnrYcsMt0BsUvdXLwDLxvlCx9VsMMyHQFAzpNCYscd5xhhNiFY2/1CGGRa2+BG6SQ8V9upNPq
xTtToS4qlS02Xss7AwDYiS2E2roItsz8b5P0FZ88c4pTeZTIllPjEDP2pcts5QCcIdxRYbwACTI3
cZiS+2r5ZPXMOdM1YbiA82T3tzbrJBupDcb0vPjWj3UTMMVJ5blqEEPQifQKkzEIkzir5qbJ/PcK
hvoON6Dv9A8L4vR3oQGFYc5DDvqsbMPcbXFFgRA9I1daM5j15mnVcu6jLVLzPhbeLjlgEp/Wzt+A
wWYxD50debpy+LkKxuwKtJ+Yr8F7SZ50dUPODB9uCHf3hRkSpKvoRwak6JJ8CK+f9HFqN0Ce9tV5
0n4daPF3buinLHrCUGIulmr+jtj9KtMZDBene/uNOkqb4p/+NJgDYnl9i9f6KQ14mVPCCAs9rX7+
HELDGGd8270d43/vn4V+zclu7gEu9HGl+mepbNlwir7cZYNs4AzG/88vZibbYb0oZ0p7jm5OwjdK
zGlMNevGNsSYOLlA5yckIQWaeSvAVLk+FTgfJKjuaGKMmDgUrdXPUIQ8NkCIzrv7yAKnMc6Vt4Nr
Tnjk9U3PO4djmOcjx98hUSurCDNDK6XHDHpnDkJWFukeg/f241RfMmdmqXKIRTZ6ENO39VrCTgdl
1v9NPYL/WhDYeLTGzmsBBuXo3sJYhUBdWmaYUX1GjLWTusz1ZZ+TM8TntI/TyXyAlTfy0NAa/njf
eagJJzIv/Ms/v6WoT8rs2Fi9TgE4sjIjeSH5PNzPtEw+v49swYbpfqKNUllUH3qPSpdYuPv+Ma5+
7fs05pgB0K2qgGjkRlRdxbVBoa3C8kMalr1uc7lVmU5urS8rHbFcBE4BDpndn0MOhOSFEapGP1Sp
dQHBZ019pZ2OWqOfO5kleHpEoYTjiBXjnn2J4uhg5hU0QeGK+JHsSesm9kSuKKpl9rFsmafHCYUc
ALJ9dxVD1wh4BZSO0uqmbLWwfIOks+kWcIW0pavODWKUNCVZ1CJjgBsKUJ/KVQOR+VhBP9hdV8Af
ypaQXCyqpGSlBWmC6Lq6m66k/e10vKEI8mhULvPpjLG0e4tu8bV41R5swv0ad8Nqc7dGn67NJyJl
kIG5X7nOD6hglUh7psheBbE4ZA3nglzzjLVBGtHcenWonEVNzqGRCCV2PzlRAdtTjDDg4szPWSA2
dzy8QA2TD/UwIXJKeYOmuTsP3QJHxLQW0EEhcsCDlVs1qoLpkplCEEN/AZyY8kLXKn4cssvtWC4H
1z7VjbFbFSmQA3fjkDHi0VtID5CfB5XnbvxB2eijx9YDygt3SsRx9L3+NFElXu3Qktw5egBkTEep
NX/OVu9SHQCdo6GfdiC3H30fWUgLUvupbe+N6rH+0HQaN2GFPCrSMtTudzTs+Mlge36jQTs40kjS
scmtalokE+APZN4n9f50FKa9VwsDef89eocIwp34wP+nYe014a9nVaFMY0zERzzh+oPfWdAHiwwY
Il613WfR7n5/fo+NC8p88EzhAPf7Y7386g7hIUaCEmEN4h8SG4ZxNQSf1NRhc3+ioA0ZOKlsByNd
5Q1cl/PGqBho4d7YElNzsH+eUWkBzjQz+ipKCA/9aBZnv5sp2fa1Y/mi09hehTKQuROx+SUusv1d
7X8PIoPq5uV3ZTMS20c6b36g5OyG5OhyIP7Ip3GJTmU0zkEyo4s+OveLFRAg/nW6MNuPxqWpIXUT
Ku2a4c1UyIjdvmIvU21fgs0IhcBnqyO+FDQqzmrTorkn1DVieg007Gxj3YceTLGxiqWUnPxLZ85m
dzT886Odid1syr2ibn7hAiUjViKnnz/uR+DrOC3lB4zAQ2MqZoBicIHjnGqUHOLU+o2nhRgjK55l
p3suTzv+C+uz8Lc/qm14JalWxCItas1TOb3+sAyXkGtKfciuWIdJadU5/3SracI/tK24yB63+SNm
pP8lVBycxMi1Ub11UJPVf84tIfmxPyM/tn4YUA+hu+bgmnVAu3ohRvsBRwr4IdtXGLmw4EoQx5kL
JYWNkQuB4Oyj+txk0esQ1DhjX54dUMY9JjQ87Lr3ZXzBbl1LUCqcAzSTzhvBhFhBY+6L+6wdYxIl
pO5Eb+bMai6nKa0gBrQlpLiHvEs1ID4tTb7xEelsBJajlCtP65aDlH0eBvVoP1KP47AC99oD1xek
Z23ZrPHgCwSBXtM/sCfvmBBOJCb8jgAnTvdnl5C3fVZfutwt2VcjjVbodw6tQcKGgA2i8xQ9AG8F
1g77vIF+NzbKW2bLn72IQPa7DP1dAspvyZdRhDID2pnV3C3nE81hQPIs1/2m+9g83gKsFp6mfGBN
l3zL73PRUH6JthRgYCqw9wT8Ioq+h9UByxglcyJPm+VoO3IcKkm4onhBpf7DBVAm5nuuvP8vWiHZ
PqisUkC8gJ+8Isq5a7JotI8dRhxsYhunxmHF+VzsK7C05Kk+Aisml1DpfozBGiQ0HvCSSmNDNskm
lcL9rQaBMzp/mluGsunzPpUcIVoftgU9kM7W3h+OozBDNLSLcFW/CQTj8tWDQg+y9DVbZkOsffIz
hi7vO/rN0wMUz7xlRuuePV8qO93HAHWl/0cvFnkr7d1KyY/yDv8J+9H9nFJ34n7ZvP6K65ahVGvP
I7eEsxHQVDfmg1hPVt9tRdqMBlPIFDRqB03/Y3MzIZvaCLPNFXStZyGxdoaDRrJUa7WtaCN7tC4L
IyFoIbh3RW5v+MwewGriL4JhkLSwp3mRLx1LvTq0pqxd51SPmKAm1hJOLD3C+oOErxJa7PdfdqP6
gyKF9V+BnYOD0W28J6fix6ElTDMpCwwFGs3KZ5JG5BV+MyoDeDDWvDX9z2zaquSBPmgx4bBaZed/
fjvyCqQWru6RzLDFyYv0APInZ/0U4HR38we43C4Kr64T91InquJDb6MJTPGRohIIVmY32hgpaxjR
5i5+m0fAsm/N9tyOmEy3EBSzLuMsXkMhzJwc5r8Sl8CHexpmmNzuAdYH7PiOzJYJN0zthnG8V62J
tzH5HaZyYK+I9zeSkIuIrCtfaDc/yZ3pGImi5BzJ67qaxSNQkpsF1vXh1w0+15dBqoGFdCZbkeCu
+J4ovj7AB7zzdphvJpVJdcyv5lkxUkCSnJxvwP5Zg2Losiue/mZ1gTh5y8Etdun78h3hwdY0C7Q4
9Hw9zEaHYQddSfM0JWGC3A8SFYn6Nol0Evq3sf0ehu909kPu7xTk8mJw1/8drKknn6R1Zwcs/o5A
Ev9yi2cSgeg+u1TBkveWRmHfDBIba9aykgfxvy+dcz/hUabRqCqHnkc02C1p3i/GvCnEjAJfykYl
+vfoxBgs5Wq1Y3hpmDFCN2IGRWVLsknRPYTUgrz6dmLDiHjg5KqHuHO2HLOpr1ybP9C8nkXLIT/N
WJ8kMhIjvXthJ+iFY5F+OpCC+fUadzNWNojAdP+l7c9vUlE1/FWO8Sus38EJ+hbmopRjK74QvcqO
lFRjMAdmNgP89PR2zUVtQ8Mt4fnz17EQS+/QQbzpd0MSubO538eFXKMkdNjpZS1ReUAmJIsUWQBr
dhqlER2r/EedHJbSjwcvg0qHkm+GjAOuN4Tun7oQK5TWhg8tJuS9YybGT71d2dcMsmETqWJ7v2da
B8QFTYIFog0l5SmIHsenRH5PbLcI8R0PZxiLvHXczVwiOYSPCR3vv3XyBrQCQcIghC1922+isSW8
4RILbttSTQYgPPphpcDLjN953rVRsPpWVKnSBh7f61PcTjNJBftEnaPWeVdj/6dnety8+Jy0qnef
eE+Qm/6btLRPc3C3R/7WiwHb3GM7eyCtxdCVrLcfzQf5KWRUJ9ZzeX4WwCbwMOayM560MW+ccTcC
0K3LjURxZ+jnWfqLLGG7aW+SfMYGOT85S2rjd6h87grQNsJXEg/pHqKM3dZfPKWWXe7SPUSOrAqk
D60ewBw6DDtP/hO8SvEk+0ogTW5WwpnPFIU0BNArYG2FU57t8g3dq/ZUVVIUV2Hl1Uvhz4fJxmNZ
luvOgB8Indavo3FuHOMcb5xLPpFntaoigSdqpA0TX9z4cKnWc3b4VVTNnTdYT6zz/VAk4Xl0zuJK
E/H6zSiRkPkjxWbU9OTMevC4UYBTbECSNhMsTTDPBgdFNNHdCqFfhqKCyYA1VdQ/U6p4e3mLpmsE
dgM3eGJWljZJx4XzJR1d43EefGXZmEm2xxr5GDS+UESZT3znY9m9dsAW4AMX4PAVT8p9GYm+mHiw
HdsR/I6XohaLsqR4jCVm5J8cVrKiWYz2phaRxUw26yydOzBsYjD/IjOum2QM/zBmjsZmrC/L5hJk
eiXrZ0dsA43VviCDRFJibsxTNHpM7fWFmHsSkjaxjFodNxBPFghUznFFRMy81Eg8YkJOwUBq+sUO
nA5Zjwpo3r05Gtq/Nkpku7ciFYpqjacX6/B2hpmLGI+jsayNT9oFQsy3BkTujEQ+ib711tY7VUTt
kmyd6lN2z+ytGdsfOIhuvnzsVsWwpoR4xwpOaYfMvGFvySqQulWwhyOCWN2CDN12y3DucXi/aQQj
frxxtopuSCjXxMbrLobcwRsmb/0LjorCO0CpUqMC8zem5XZoF7tBlHx4EnOU3WP9nt8MrzZRE9Kv
otpejQh9VcAyEPmh2pfaAF4Xv7T6xnAVwCLuzsLr9A0PuoKXIsiKygEr3o+bCaPiAmTHEdtqzj3l
wT3BcoBaShlLeVtx6/N21LkeksyOiPxsqBbIJepcFciRknVL9Rrw14gxVAzZNA0QnR7Sl2D0ebjg
WxD2yv9GvLrrG+cDAAN65V9SGTwfQEBgl7RH/Iq6AQVbaan3Jpcvji5/5xsEZ6PL3tKE+Whgwz5F
I+tBhCDWzVT18K3e7vOrJcGCq3ajkI0/w9csF2kvkfL0qV97+iB1RNgzaqgDKiAYjU+AJ9oui1gN
nYZxrvji/YV475X2FGaFuVSMkkrRYymgtQ0lHnSxJBmfgFSi+s1T3Wk/xGjXv4LQ6bVxO9CTWw2c
BWzDEGNOw1Wa8UK8DFC4imdpL0KGx8r24S2bIBt5luHEtZ6DRRJxYi449MMG89MOT9FNTohjBc0m
JmTbjJgvvQfwE1rILbT8tPKIPNUUAgjVIwukcPxc0zR+ASwGlksWXFcG5IwOeJtV4uhumX/YhgZV
nWdF2jiv8c2hzwEg7NfCnU4tduibYzdDTSSfoLcI3IxSAAElqmCeUCd3Al52pzbavinj+pjqnbRT
S/6ZePLCP626PGqUo4IbdRTgQns5WxpkAIqEtAv0oFzVrcKkmgI9L0qf3DfM1KrbfuG2ShN3pa1e
t5ZJaxr6t/aVcDd882m77WEW9kLUAtnPclL7yLWWMK/hsXS5b/lgq8cMZsh+ElXC48clGOTJWnBB
bpUq/lYtKN1lpLyKmbuPDM1QcwtyllS7WbNSBHXp2ui2JSoU/SAA1ksK3IBmSlngnvL5P0Q6DVK3
a6heGufM7tAi3xq+hoJhcnSimlwsxUJNCdjT3544IuidPSRHwE2hiqRXgv11hHuGc9x4aZ5EKVGu
vuSpokcvcUVfctd+7ZkyJOgc2Vz2fBaXNYfGYMjsLpLQ700ImbSWBLhevhgyZJoRhHKKpThXi1XW
W02DUmKR1klQLd8WPD4h+uScHNmngstU5DTq+DoQWc1I/ue2dKN2zETVbbLmGtx8ySHIsZs6KNxY
g2vhWe6+Wcs4oMSmMECXZsZ+p9RUcLVssydGyRa5N8JItHQK9OIjZu+GoQ74+KGKM9IGB1605zmo
mph/nZHzxWu7y9mSkWH2eusJQ3Yt/XlYmwgFD6wT6dU1EvBGYT0ynVbGZAvaN1DGobq8qt9ZC0Rx
70TiUZLLlXPjEFuBLrz1W8YIyaLJIhUKMkIOhkvQIUcntFgMaIN7W0YL5dqTwjPZXDBJ+rUetmZ5
nY2GHhSt5La+auxMTV8oSV1FcFow2gvVBa5ZudgB5jHqCR+0DnFOfAQZrK8fKyYQsRnWQ2Q5a7Xg
WiEoEmTlT667s/E8HEm6kn9nU6Bi1ZaRfJ7dTg1KXCrky/qH9TJx7doRAeMRtBjjVBjWIftKjTG3
v98j3AKMFGFjSbVKD3Zy9+QNez+yHSD6E+1MXQgWM8u/83MPC1lG4TZ7c/pzCPzD0gMa/Z6/Mmmn
Jd9IFkOH4rd1XzrsJaiHjOP5F4aLI5tDRXqsoFHxNwWStSFB2CmRODFM73Z6R1IV08dUzbHVdSo0
4qfbjpq6jnz8HKLI1h/c4jY2WZVjF9ShpCfXnm1+FzsorYvp1Q+H+NmNtiuDbSvIubZ+ZpVKs8fn
ZunttnMZCpDQFmocy+u5CjO0VeiQe8XEeITM8IdfPnku754dFGhAUsfBwAlJDhdM5IfGZkXixlP9
fl2/cj3Mabi1sQCV4NvSVPte7wU6mYI/Hf8IBTo+qDxIi8osXQzdxr6KULYEqSPHuSnqgHBQpF5N
IbCh/ZcNS1nT8WyXuAzZHKbnRtFZa8zeO8Ou/VlzDLTP2UEh9yMQbjIWOe3zKT46/wtewT7taYBi
iol52+q54xB7E8/AnweZc2zFn78O/pqkx3wQRMIXEzPWa6desaWCl1B9uRkX0suTJtfpDDWa8kBv
2er0kI3KfIlNZ1KYM+CjwZEL3qJFuzQeE3vzYZ7fG4UT3X3TkePeCl0hy8KdUt9azYVXq8xOwAVc
YMhDeO3wEXdOrIehVj7OGdA6tmY0h+NIQgofo4I2l/dCwrIEumRH9GNExBoJ0HWe0qoMmrUjvI31
ZuZD0DKST7OxLTzgCogBFBdvBJe5lr28HvfUu7b/13HJaERW1PfbxHqvsWTUr2otcrbu6Ic0vCMQ
yrpZfKw/I9qSurHeaoFWYDb/aFgK6rVXb6oSk9mV3Oh4x4HL+z530tu6iw5Fkw2lrjAMBdfqigRj
ruH6mdSjZBX3E5B4GPgz8/9XndLmi6+hdJXD68j5Cu5pJmY5/TrfJ8D/vTbK0LYbnKw7B3d5qoJ6
qhCCq/+qE39W8k5Ruk34Axf341PTJgx4UMk0j852ytqhebe4hI5Bzyd1GguPotSFwzICrvSTFJqy
l0L0PxAo3/jjfLVmRzOeTs6wd/XcFJ+IyvV80jYRMZPU5dmYBRuy14ljvfE0JUgy2QMSkWWPrxLd
2EkligByKENx4yy4+QVvuqxLpOZzdoB2RRKgjHRInB9Kish/Ouzoy3nN/R6tMiTHd9zDdGfcTfsg
HP7b8PxTSgYbNAdR7YLmw0DqUE1HyuQj+7zpq9w79fmvawdteJIfvG5Rw4v5UrUFP+WpzfXEQvz5
HYTkm7pUzT4GEJ6Zh95eq+HbgGNsI/aj7F1TGiWQ4bY8K/5t77C42YiHwI1w+nUYYQk0AZGagoAg
EHyFq7wPNK1swp66VhWgeYh5g5PyCk5t/zfQi5UteoR9/MsnjPUaD2Uc5wRBNv7GD19ZgRes8/+Y
n47bAuacHVdV/WrW0Sp91WoEFu+6MS/bcl0x4r8lkW4SS68g5XwL3aJTxPiQEBtIF7nmXiRZHLvO
OEnTLMcDMs/4sbzmrCvUEC+ibCSX6ObPazGZEUS0//MI8DaFzJP96N3hmXLZNHWVXcDCHUt7LHHw
yqL9JpemgOpDWrNOWuNqhWfgG8v88rwLdUSH0QwzeuhggMw2n9bmY1dpv3oCUPgO99x6gsAbVUmB
6FQvBScpthhSvuXKgg5qFogtZX6dB2QUG0PcRqEu+LZs2VZ9nnIRy7vulQupr6Q4HCkV+j8GBQQd
KUIs8UlEw+aw/vWFLF/vrcQ5DS5RGGx03YN0P2+r6eUBqrFIRpyjoyAhRXdWumjZIGQzxIpJ2aId
5shX1kJaxwKIphn6b3YTxHhUc/6t7QNPLiUP0HLadONOFuaLX3NpJAP3eUGbOa/OqRlU0CBYWSmh
BGRhkxf9UdB0za8bScIDi94y1r96rClKex3Gd6IFe98GBK9FbU/mULdhT10n+RQhtLenFO6p/Smw
Y4uzw89sExZD+Tf0CHwXISYnRWN51cf3G1rLLmBBCnk1s92zU+ssGSyriZZU3o1JPDJhrTBubnIz
Dy+5Ue5QB5wBD3Q01yr83TyV/D6tjUJaRaK7MVs3yTL7zatYzx/dx+srDYUousG7St8pqulfHEI0
PanCDw/SnDbVWFJRp/NK7kTUmiR9W9oNGssUyKgX4q7FTZgkDoWSTbvv+dTzIkdsdLtW/IALkFJN
w6YGMLr8B9CYFcNDgRsuKocCu2bPfwLErVu6mo2VHOFJiC3oThKCmthZTIMlpBaKIvH+IgRAO8r5
BMlHCV0lblOL1Fm95IrzQtjx5aKa52soxWp/17Z09TfJ8nQUpW2sllTd/6/dP0HyiDv5CJhCILpK
5saQv6aC7UtMFWAbgvM8x0Z4Op9kkCVYCH26YVQq++POtnDCJE4+GhdiKFCiG7YKgLc0nMbpfKKf
9pTKveRJ/6ZW6VBfkDxwIuTuE/Oi9oAh0QK1ZVA7J7uds+S1lutWuYsasgmGM5yGjzqrtuUkdxuu
tEjJ04ykePv+8KBzlS8wSgt8mhn2zAtTojjwa6mLRJLk9LLmq7N2AtUsC5vZ74uYuBuk885mB6vi
jWxQYhEell3G4VFANOmzCkvtgrFPon8x+uTtep20nUKOMBgTmWT/WD61cHLb9JbWFF54os7gcTnU
PQFnzvMQysTyepZDL/nnKnssMkoLCuyQMQz0PN+FocN2XTfSpfMtODawKKuZOGiotQSegQH/6dkF
THgZXMF5I4Vvki8OwJuT8Q6KiZQ1c0kBlI7s4JUB1AjNyUu5S6yDa592x8a/ZZXd4lRpXZCvAV6/
1Ujo3hMzPzrnGZbTEdINVwm4tAE2Ij/LmcpUyQE47M+SxltbpihG5Q/Ju5gPeAXIaAhNV4nKHSt9
dDawNOuXaWPACkrXsmU5uJWUriUMdvSl8K6/7poxtwS4Pkyqutw8insgF87kzCIrHTf5ewXhiFbF
NvZloCJMknS94pBx5/jSxqJ57rzi8m9mSNhKbRF01xSDBnGUISALvxxpzIg+mrsFfi38Fo4MUIKq
Vs+4ZUSgD5wCW24tqAFDxF0rVDjL13i3AaNY21qE9sQoKpDMAuqLwGeQ3UpUaAsR++g8bGfEIq+G
XYQFF8kdoQKgGTweMZ2bdZSbSv5pzhq61xGafhaTYxuF6EwmUnYN9KE8K3flDaak8PqzzXJQm4sz
pOR4ZzK3f+s6mJbSZsNKSUJoJWVOQtaALtNE+LmkN07TkhjlmhcrPxucUXKzkiuRxteG+qzZIuxF
pe224oa/tYZ9OhrXLMMp5AmV/XNmoP0vSxB//0n06ebphXv03MnxeyKdc7Ilx4rZF2/v6eYAE17Y
COx7+fIuDsz+kJ5KRAz+Kw5xVnjw7RsLtJVCSO+jGPWYWVkNjCHXW3RKyu1lJ+6bqDqvAZMt7sQm
GCMDP+k00xmFs6fdSkZgeI1+BxNzmFJIbQy21B7cDaWwvZv3BFT0eQ5ONvZdxplaEGCrKAl6B13G
i09KTwx5j7+EmQiyXmvw4LdK+3RfMWpJj6qutj5b9Y8hif+tbkcWhnSpXylu3scOhQ+Q6JNGqHxV
mJIYFxjmzDCRCuAMvQiveaSf+HEKpDltR81kInSFv3g4WQhCZJWZL/gcjuwuPawRSsX4+YSHlyeD
J4iOG+hvd2WV7TDSaL7OkavFsqo8SjqCP1pm2puwV/wmTpNfteJOlfu6dok0CjfnRvBrmyGo3ikj
iFYbapisl289VPXvknFg97k72h2ioP0ytAOGoezRP5k+LGFtr+oSI+hu6VAzS3fk+JE2vEr5QXtA
EORGcGIKjos8/h/HsWpNFcx00GRiCVz2a+EkhFJrasuO7N05+PVYX6VBdpsWQ+xBdddMBAWfeIll
FZ11qAfpOI406JFKPqYA69ha/NXf+hIGdaqIqjj13dEEyxTqB0Wk58EhilmTSjejXaZTi5Y1Y/yl
S5ActCqEuDn3kaC59HbAN1o8tYwEKIQkTAky4sWYl8sCQbINRxrUKAcHKZt9x2fMdv8JAocDkN4v
AARGYVYL8J5x0kgxohaIJGN3pvyk0oKzCQzcJPM9/8XBrFI9LyPYIb4GPR4ybK3rGC1zj+1kHs22
Dybd7uI/P498GRGmla9JWZ/bsroTPDVcczGEK/qwriuDT5TtnEvCvDCj3Uoe098uNGezzG6OdTJH
mZYhyVmcQ/AC7YRRNB7QBrzskHQdTDxuc/F3MOnwbK45uo/lOJVQv45ITdQyKzsdDlobcK9R3QEd
2wgfdJWL6bpusUEcf/wjeSGzzTrHDs2jmVaUCkk9C30nEqQUuKizE9GFUkWnnBriVeEllfy2pTxO
9ti3LxVI26DCJ5BvJXoNEeflJc7drvmC4VB/ms9GoZv4Eha0XE6uqYQaopD09fyms4j63BwFqHfU
iedjnBjsDWsSGI9C38NVjELXU7klwi+9lGODiOhMKWzaGz2SsUp1VyTv15xNEGDccZfwlNv8nCkT
5fdZWFADje0Y5YcsfmpI9fKvQOt1CJFdScIsFfB0s5mZyvAK273hMioC4mX735RR5vMurri+ygA/
bEzKtxKIlQ9PG9gJ3UoYo4hUV+HMg1Edmhgbmo7AsX471j9SMWV6N0B2wH5jOgkhSSIcMo6KXELi
jAdh5dxT0IN5/TgVEv6KkjNu+IrH3bSS2yjSsQsblE8OkGUmWcTxiQZKR1IyP7Q+jAzc/tBgMqC/
G5Qsy4DonKuR0yjKOz0aD5DypBQKe4WxVJQaysBOVD/5KwPBvOEGm03zMssycXY3TGu0yvB7oD5c
ZdhzV1ejA/Vt1HfjNU/4ov3nam151OkKXjMgSxNJQe9OM/J8UJR4FoiDMadpHQnVV9CX4Otho0az
P8CJyIZOIclmKlEOtc8AkoDr27n461Oa3KjcGJb1zhcKNAvIzzWMvW6iGgU3xUg9avGkYAW7AcRv
RHZejRvNFupK2oHd24KmAnZWYZXyiICA0gxg1LqPLie3qD+Ea3WNuFjlPOEO+YuMcHzLHtwiMcAo
oiXcWA/xhNOyPX74cExMCKaMdEA1ONmOzPmWXE58Vw0+1wfu276b5MjCc/T4W1tdM+swAhRp7ucu
kwpn4gLR5zeEwHpNhU3RyZUeaTWTxxisAEc5WkWA61A6mN3p4rvL0mtW01Eql07/PIVtgAguNR8C
Xr/Qnt/lOgHE33/9aBiSZ+7vadV/KtssM/mZvTDkcl3Xv3NEN3MdHR/Mo8QMkUVqOh/4YsnetBhR
TZEab+5K2snHb/11mALpHc4uLCFe3dXFSs6u3Bo+GwOwzEjUS9zPMe/sid8zRhXYdCC+4OZY95gU
+lupQHM0barn9wxxQyabMvtMDrSbXiAWodg1CfSN8IDxomgZcy3XPo+l0C7ClVfiiPszWAt0FYEt
OMYKaURtMjtYqSzsCKHZ2CMDVd0Q7P+Q1u8hm2sBAQ8DGZNJ8WDr/3LYnM5C8f59RdoVOICeqq1+
UdZuySZGaNXVl5+XUEO1gw7Z6YjVQpy1+khGD7MpQo0S6USNzOxfyKP/pdxRNjXPqXJa7XEiI/rm
fNYDYU9oZC5OoklWEiLFVTcuiAEnL6JR+BloDsQ+xUQVd+6Ra7lZ6cLUm5dkdTz9d5Oz3BWMBpUP
P6E9pgyOieVT4DVyHt5HFtMPWpTv/mUOajJdHAIJBw9C4WPeD1TqHSP77sJ+j8VT4Yxw1VXoUCMC
OsU2WJ4r+L7reZtISNSRtI0wgQNFMLLIOHqwB5O5PIarIBoc1CWACRPIJhwKMEI6yjGAOjVelNAa
ZaHC+7uWtGi50eQbxb5qc5oUwPXN0CmCE6+kScebLUXcBLolSBRinG3a+kQ+DdNvmf2apqpfEoZy
es3ul8UrqmbuLt3sPmVNscIKHl/1mtZacUr9PTaIsIHI2mDWLuG1q7/rLb7V0H3AIlzPLa+bZjSg
P22bJvrE524IzDy5wK8w4CFhVSG8S21fCVZoMGYyvTMV3+oqR3Ty4O9FyTgvqZlmJluDTLNQlTI5
rVYXUQDI+UoTN3iIW1XvmQHISay9OgcuzoPunRl39S+APPFxkemwLTS+gseamez+soXzvnxRjzGY
5yXg8E1vCmtDm+YGXX/Azdq1/jZXURS7/LwN+tZzC6D+LI1u3zT96pmj/VFQgngeimF1bN7GUrhZ
gClZQLC05HzmTIUq+LYAGKQYNseAeJObv1ZgmSs9cd30ZXIaCgNhJCF2wRpPtzDFfwg8T4SovJQl
JiWPhYVvb7eBflduTyKcvy1t6u9Ryj5EqNYtgr82nSzv7PGJIkHSHMajcb7UnEcKW+2m6R+OY2B8
TVkD7w6LYB2kMmcsSFlCfUkpJlLrX1fDXGUI/54M6FLD8IQyPepZ71pBs5Da+cwBkgwqQRVT/Z/T
0OfN37bm3ZOwqKpqi/Reux32AGpF6zsHFPoYGXBgidnk3LLGiQJY6BOOIFrludZezlTOab/XD/cq
ffWCmNE2TqQ4wP1Xx5wRb8fwi8IaxgBWJo5pOkNVcDE93VA2e//WD0xNnKEnCKpBkuFjUnAreh2q
/SU05LpUsc2T6kUmvrdcRZhCAk9n8jeiOTZxBN9GECQ6+3a9Yt11QbPdjZhg3C1K38dfK0XbLtyU
D8N78acLdR/a9OfYssHk1g7zl7I9LmydpXQTcTjOYueu893hopE0IUKEaUkJ0xtQ4DmTsVuWdRkI
YCHv2wlEK4fWeeyVaFRmlGGVUHcTshu1V2+cniITlSY2Wr09ljMoY/9CsJdjT+7yheA04h5YVksX
8HuJucO42jKmV5R7XQaPV9a1RkTAA8g6QdHeeIJZyS+wmTlAr9c28Glt8STeLycoAPxE7mZOkPGh
T37NxSro2/iGSn0W36fwDV1VOVC7v6SSU9xuAw0vDoG57rxeunouYMm7Dr33sc0+nGLU5umrLuol
4uUgF+SFZJPK4PmvS2n8jv0vGQJVsMZv9720x8gidnckii2x+JMyD7Adth5HQ6TVFwlToXXkuZoF
27De5Ejav0DisVd2iZ5GMJNosccDtE/puz+iIN5BYBxNe22JSpWY6thzgdTZJOkzljScupOeNLca
nQOkD6EPepZaqzOjbcQiYrIM4Zs5kfPQd58pVpR5IY+guq4cj35BTyv57efBwU5NuIQv7XlTey8Q
Gyhk4/rHaiP9vX256rNoypRXPA0m49sq3T9i5G7J+vylUQHodoAUmISk1vel0A7nYQzehFRiHL42
HkebqyBmDaOLaetzyAmaXzfvPanrKh1m/bFyJUpZ6QrNYWldpLWjVuBXbrt7DrbPT5BThJZ0VJTL
uv6FZ8qJyrYOpm0orC7jqbwV0g0vejr1rova3Xje+6blkAdMk1cppbaJDegx2NT8tAr52HdqOzQl
rVPfON5P560ebYMIklX/HHXRMaodjoTGzKTMA214TxkZKR6fVX3XyYab6c8jhyKpnRWpJUwo2PfK
LXvWEqPfZ6bBJ/kQcrtxn7X3pQdjbKYnWKCHx7P5HqwJGwil9oze8juBMwTiiUnbZBNZAkjeXBfe
IonQv58wxVQZTnqtutxY/z1I/P1WZREoBHqLyuQu/Y0XUq9MxxMvXuL2drYbruOw09MW56U6ibz3
kptK+uSodCkCdKAWbpQkdhyiWND3OGDA6O+NJznmQ1W10BRStWG1y7pWm265d4HUBcLdS1ZPHYk8
ajVShbeTx+xWXDpuvRqm19LRsT2ouSRgGiFdoYW5fRUObbb7Q9HLlKFf6ZIaPpWRlkY9Lrq8zmBx
pdNJn9khaTeTiRS5xJqonYpecBJe2/NcHiaAoxjwIxF4m/JJEEgU6v8KNn0SZxz8pDeCbq5gEqq1
E+MlNR5VZzu5NC/0vo70jpRGjbPwVr2ap9Y0YdFX7nJWAnZ1bDZV05bd+PJ0MDKWtkBc6DsFuUdU
50mxCBswGN4x0tjOH8Y9MmI7NNHpiNupOFyJ6Oq7+QZWImSsaqg9IL3Ahk4mSYzYUBpfBcGfEFTj
F51Q61eYEl+oqDBdOZW1M6IjnTa2uFMruciF55q8MOA0DE9PwVBXhvmvkCTZcaZL4wmq8Khl3hUY
nW0OkJMmF12S6eXYtrq72WGuhQH89o3GXUrSO1mloJ5xnB4uNwJwoW/zvVkvoxm2yCRWuG/3TamC
mt7ekv5ocAitu7H8rtbz04t8zR/EBmnb7AtRuAwaj29Ey1IFyDMtN5YQ3xO331nhqGrYlIR8+dkI
Jejmj3H5DakuT6pey8oBSImbknm6uAHnAayhyp4dv1+kxraQE18VRiqu9FX3gkknDTmXKo9cIvZf
PnaYSPiEWa8i5fiToJ5Br47f2U5AzYG2nT9JiPnRpWi0ixVnMWYBdnbtJT5d1Tepq2KKg9u8UGjD
eKKgEK+vWEqlHMh01QNme4ung9saDdN81wqastfYF6KMQL5esW0SKyWxtB2nW8ZPH+ZUhcdFAiuX
W1wmddiBdPxayXRGUYG7eFdMMKXRK6uqqMMbrzWQaiXXiNhmPUGJWHWE7Mufgu09620MnQJti2A3
jf41oEPW0IF32TLMLkXlvpXdVCSXvGnUEkRq2odN6LC9SYzjP6mPt+VFeXCTvQka9BIPS754km32
igbUBHPbfdrJcvKzj5CF/GnACLq8Sb+RIU7Exaj2SG5Om/Id5nVDaRLH3aCAA2XLyOZH/ILiuzFj
HF8Sjf0QhYzfb8M4kb302Mn74tluEj7ue7N6dM+mxGuLurQMQoUlQYQvSP/bQY/El2dcNHv+C22x
PKjXEU/haOBNtLO6cPrUg4YHGffUP2nkQM38nvXYP83BGIuSHtyWI9rFWYd7ujNoQ5OjoWxkKE2S
4sdOWkziYTlpJTBEYzVwvDJYd19aN32SeNJ0y0h7/SH38jJb+GFqfF2mo0p+GZXGmIYclVb61e9Z
72svMSrPRB0GlRWHP5Utal3SqvNZ9RBAYMUQdBkHdYH/M/WGJEYdp7518N85pwF3t39FBK+fMwTW
LHfrRn7U2pS1a7pNMKvC2ooSWaVO7Gzgiap+xjbIqLztJzIrzkMRAsjo3AK8uufcZznhpCGLc4x+
nD9i02aSw8WDKPKONzM0TeVF6IGgbC4KelJ6gKb/W2pUWyWVdjma8LkJEfLoRamMd93hyvLwyzVB
aPzjbHGS/LwtksY4cxHPkuA0OAnyy0bsBt6SWxQLzA/9frLMT/UV8K5oldFmeUGvW2HENyhwee1L
uAnJTRofRg//6GYlQHvNZldLn1HbKLChNEe6YKb7cs8JNenzJVyQF5nEfbzr2YjF+GMpnQ7YbV0O
U19NSBytcy0xAfjKJ+eezkvJ8mmB+7KwSmk0NOQhQGOQQgpKYw3PJQfVzIG+1BPFPqd7PwIugf+a
XJIHENMQXd5O9jbhvmVz4zYB030BdPMGLFwH9nNO6EP10W2XL3vbBFYVGTZ36F900E8c0P4wG+6R
zAFkxr08qXk/1hfY7eGJiA45zF6o6dnNdmeKbt8iOkFS8LZ6sR8SfOVlP8c5h9LgmCfH7ztvjHYi
Bbtt+gYPA5iFIfOGdkCkcMWBpQF6HpuKQOdlwqMim8v0+6yUBlk5eenT1YsSuaWcoimPjt4FkFvG
jdP1T6BalzNo52Lcwtp/xqnUs1EC4/B8gUv5E2D4f/rRQgfXwQnRhhjeG5m/tfSIZmUZ0osQ9+tC
MAqC/7COTiUgxJvnuk5QeuwGL37G79LzL2RFN0UMTLx7KxpDhXq/RLsuGXQ6dYxw4Dj0HvNgx3Sv
I/B73xzfslDtqSkXQYvwoC/LeTGpAgP0pE7SK5rSP+yUr8A9S8YeVIA2A7E6FlYTePBvGVGeyyw+
c/IFSmHHprIBNi69yGKFNFHb7K1S4pHCNKkh6WPb4/xH/Mqf5jL7pA5RsnxwUed/wEbeMwFlPyep
z8w87ZTjU3w+iltKU9deuOawBftgklLwBEcB9ZEMCzGLMFHZBbuP2zDdtozmju6H1cLyFSrAyheY
PvZJiDV1Cs7NRPKTmr8jUffoW++4wffyj4VYiExQsmdSx5/BlgzH2YQ8YY/KCn30IutMpfHs6dnk
WFqfti8EtH+nKbgJu3wustDn3UBAthgOkTJKb7dZISUeAt+H7sD/Ip2KV0u2oaTHK3FfszXz1DiL
Dec/OQWTFl7OYKNFi1U4tKbsAOwlkIC6cWOcbfA57XsV3Hh+lBOcSiWnfU3A5T7ClWqORE5ADHwY
ClqeNniTq9Iekv79G6qd6GyRswCtUtpTHbpqb3lYUws9qv5zDJ83ahycHF91ep18Ar1aHSORYHWi
FNxm75AO531tRlaKgKP9auu6nX2yZIiuJG9WW5cEjqsmVwHgsWvhBGsQcik/ieEy0tHPF0Vs843C
1gNtifJFq3MEUSdvOpiILz0z4Z+aei6zKOTcvT7ymSw8g58xHiZwNmEyNKT16RfTtgHvcejk6B3e
tupKQ2Za7LB3b/DLZbrNddfONmZEU3gGcu5rQHSP6JykqMUFvC0kdB0Uj7VI8DlV8DObV47X9s12
F10q2KtEJqytzR4qCePyxEmZpGUIuP8G1nELVt9ULCxnnQ1Bs/fHxujp9MYbqaSLwIbM9sgilIrt
BFyFSaYZhfAek9BrNpJ59WpnfbYAvdhTr9TXozkSzbTCFWXAqhGR2nmVYgRDB6wuwwqVgVIBIyEk
SFHufsgw+LDywSK0o38Xbe3Y/q45nE3FxjvvTYPoI0xtJM0if9Hiu98ejCci7imkMDYIMlhspTB0
BP4ibI2XR6dTGud7zyGMnE74MiKjYGKW61vkclPdeGAZg1XCBO7vPYtobpZ+LyPIzTkXt6Oq5kpt
edaV9EwmksyuyBZjE2781rYb5OB8mzvAxJrtaI4udLUSw/n8smp2xYpAsm2sC6eEkUA7KhuTd/8a
U9nW/KosytS9sWGsjVOqsYjev8BI2nDa5hx9zq3+NXIbEJIMZ0BQPHdULyvdyZGUGLU6ufMYzFI9
81yzjTlwpCMxgUUZWcEKssf4aDz+yVY7BhLqCtIcQHrY1FAhDcVDOF9dt3WL3AqQDhw1Vr0kJ/3f
58Ep+oDvSpQWYt3glOJ2o+K/WSm0OTWhPz+BBVX9chi+NyV5xAQUEAZjkEZF2JIjSwgqUlckyNtx
5QNTWmhUCBGGDixfzlu62yIkaPsHU1K9J1YqfeiQR90/kS0xvXRqi9Zt723PmSAckwlHQwZZezNR
QYDN/Ps8YPUKIAjr31odgirEQSFn6ERX8AZAfePPVrILqo+9CZp7vwn0b1SyFyaUgus/vgoWo7rI
H+3fnlsJvy1QShPzf2Ogl9MBh37MLlSKvoUgTd0xAG7n9JVrD3y7e4HuZ+3k7Skxi3JoVU2QDaH4
TCPvPDOQjzLK/udQc9xsRXCKxtiu5r8WM/wsbZZb3ZD8+NrMOm3NRNuyb3wmxgu0fOXiCY4pE81t
suZRGbJJ/z28b2lApNluYcW6/DReKfy1gJsQ2AJB6tnK/8L9mK+bdz4AC+8qW5W7APa2GoZm99K2
Qw2oG5ypWwI0JEHS64BumTcw9f2Kwq4KkXIkTohS8FQsBI1eV8wZHZ3y78ug7YklO0lk/eGr0O4d
gafMibQCWdE8EY2k6Rcca1YlWS3VvO/Do/1KNanhGHv4j/BFAkqsNEG67D8J7E4Pf/VJ7T1WbkDH
C883MN/sgvcIFCC63gj++QmOTK3aR1hrRtMG+LzFYTfAeeZ96u+U28/hICzXdIPCCA1TGdTkBAYC
/4XbvKoEhspq6qtDhSeA5ickX8J0k6E/9f8obirkcykb/wVWsy15HRBt4Kfm3BKlaid2BK5/bM92
C0f/zwkNDxvU3CCQeA4eYnr2+6Zl+tIhKDOqkEfF8wMyz2DGANvnaMuHHqwU141Be9O4izzbGzG5
2e3jcnFEqVyoWY2lo+xdy4csw0+rbM7hR/SoB5UQW2keqmT1ogFv3sXjXWmupnQpPJJYsBiEEfEV
baK1MXI70QzAshqKO3BeGg2mSLM3iQz0P2zcgkEtE5DXJNc0KssJ3AyCDjUvH3uPW1yMImrQ0Csa
GaDOPUG+XDkwiCo5QMP152hix6RbkeD4YDoNGRMzDpHeEhGK6z8clL26eSpNywh8wCwzZKl9gAq8
1UsubDstBpLCPThowCMGj4ul7TBKxQlp2CWhqhdW9zMY71KRTy1Otvuw8t6nJ0WcnK2orQuzrEK0
lp5liqr/Jw/85QFfXa9LMTM+qpCVyCp+mMooAq7fUYdBHCV3VbupF7iBHzosec4l4gZBQTwp/A0x
m8AaPufXLYF3bMM2tVtDvVFrolvSFN2ksH3MsWOJ2tiGrMgF09j/UrYWcOzRC2GU5t5YcF0pnCTf
m0JBWT1e0s36vIwKRtKYcULLTK0Pycdwe7zRB1zr2AWXikwm9Ut270cefptZuF7qDoOqOaWwvQB5
KnlNx9Rolz8UM3xQ/ciWEaITkMbCw8fJNbNj39+ZOjG/vCFd02aC7cHiJybuFAPgFU3Q8IZ447I4
VwXaAIzvenwGiINPLGxuE3CN4/tp31Ney/ZiMuEXU2HTbEz4vHcRuYavnHM2RzEa+zFwzHsQ1Yq6
KlqWbLOp/7yOXum8TmKH4N/KDLwEaP2n6eWI3gnks/W1z8DuPBmM35bL/IrlecTXCMVxxkjhtkO6
UBMh47K3wo1RbbzrYg/OMQh16mc8ZIbvmVdCabSM0optjagEilXqCBvMpzBEnLMuLbgwrhms+zhJ
MXSFbi4LKMCSpkF1/nzVwFQw6PdCqveiyaheVl8mUHj8Xg/CgKEm/aEqfmIHh2Z/rLrQae7CtY0l
jeX75EEFyxqvnAGJQFoQMqVVcF57sTxcmI88QLIPj39WOmmClaybUsLAtRa+kKHgMYNrfkR8dstW
LBqn72t+1/vBMnMU2MTxPNN6bJaLTu8El9Y3YY4M614sLSuKdMNamKr1Kl/9XbpHD7cYgXRDqkZ1
LtGGQx4uQioHaP/tyWCieiCaYj+UHkpfPPC8DbK1dcudAVJaks4KFP40c29L5gSNycWeguXcxZ1h
wa+u4ySh3NJH+8Z+hT+UhB3R3B2LFWT0jmsshbIJq8xirm85MYW26kNaBeFlrs+uUuFdMMGPAuWs
rB5m9AyLP2zW/qCJ1Q8I8wq+zp6hy/iYeNEPq4bATkICdmxcy8wE4q1kUpXXge1rhMb4kcD87AFs
Y4ENg/2aLWNo6mZBQti5VVvFwukmGKNCtoZCZFgRJ6Klw05BI9py/aHxDQtBL/DkjNoHAZTzPiqh
sidF4FbNcXAkfC8PT6Rgwcue/x2Kuno58anraMCrQXBVdVAuDBEYE+kjo4wzEef+ZBlIFRXEniM4
X68Uzj4ExyPRGZJxUc45TU2jZzVQnnpQAW1zfXGIILboQcNywZgwKFx7JhdXpUY4Z+B+e6Gc7+N1
a3wuME+rtYk8RDaxmKibzpWWqbL78Opm+rcUBnzBxvHYDr6TyKZvSTbd2RyuYrtlfAcflNNwXNnQ
MS/Jhhm2mHYg+zi0kD1OPYKg2khn0rlMadC1htdiNcoo7zjOfyZn3LCuvdI/xxWL6A7fYov+7Ocl
j8BmlZl9/F8jCd5mIT7MuPLbytU4MxqvWpFQqa6VJro4XgVdS4X8mWxJvlUp8K9G6vzXO2DvhIxo
N1datkdtJ/3NRpjy68vVPteCmwMrVlG53+ji8AmpD+R0l+gtBv8VAjblo1sAiyUKws7Yj/VAcUfk
8yTiNXHyixyLObvsK46wLyb/Jb81ulmpOyyfuLRoRpJN6SPCj4zL+slrVv24wGtFKjVVpl+wIsUE
LNwLYgOzIBbKqEm3WWT5WrxggwFLkGpfzbVhTPlzm33Kh5BPfPlkfCQ7Kh+hgx72vdFh+VaWRl0p
9ACJBgLiBzk5VqhHLD+c2VpAfMQcbQ5YnQ2PBw3X04iT9TIW4vUOsSbhIfttOBhLXVM9lq8GgVC7
7dtHl24gR3JfoxA11TlEYx3Jv5Yg09Tnjb0bzNL7BI5RZnw9qNDOtFTtXdsdyTSFKsnNg2j69ryb
9cUs6tyC6yWX75sD5kDFhNuw+ssFoIr82GR4qbDVm10tgnqkYhhjY/ru6KlQPBu5AaqkIgE8ds0f
/KOEjR7CYE4VLzG5iptjS1sRF5mY51dk2xtaRSGR5LbfshYm+ygQP4VHfDJlCEq17ljK3YKfRYzM
/c7JuxNM1hefmTTE/BVoVcDy1i56Y8xNtT1F9W92NhtdVzX3vf1isvYaVan44cWsGMQCZ/4J8k1m
9Tjz7BBA/OVA9iJChiL4BbjwLCEjRTClwW3tzSp2cGFq5ovK1JheErebC1IyjOfU0v2l37J3JuXB
Lz//ObRFSXtizW9ory79pkSw4QX0lAqhKQVF6iUdGKt8I7wrPeJ9GSpaMTKK52dfQr3m9hlPJAwF
jkgFKQhtOK36czDnwD2PNN+umeinEImOmTDx2SswPie87AM//iGg1uzaRjbMeD/NI+Y6Ivhiguhx
4m3MvzkS5ceOVBdCY7mLV2KHD7rMWep4oTtGk2wS2EVVEfo8H6zwOaCcoYPiwY2PsiUOJaNGm8Fn
v4tosS38MmhfMcmkjGdtFnNozyT9Fvn2FbItQU6x1TPhh4RdanIabz9HEixeq4UngEZ1N/AEqR7L
X6peZ6ydnAcQEdab+NuU9pVSJHiwAOEP/X7sAjEJ0g0Du4Qdq+dZU09PHRapAu0yoDKnf0VyMmOZ
L/KZMwjUdhG8ynrSIN3QpVT3vNFjlF0WBM+iz33u/RlpKQBT0niGNwXXUNo6qHF4+Z3lEKcDQpU/
fhnR/wxPfsR1mZOB4zGjFPItxFPWt1IO1nVL48TT3ItHDLIJrV/jdnaovEci8PFRBEKrJrOYVnQ6
SxE/XmqiDRS2FuJ3ilPWcrJQCzhvYMsfTmBFifs7G9R0ClomHRfaKo6atefvVK1gG1vVydxriTl6
fB4xEl7K6PWjwtnyyYLhHY6W2O8pRgjlmHFIxfPKGdiNvgmE4XUpKTpUXT/r4FbQO/U8U/e1e65g
KrxY98wyxvucnzIYGHlyTTfs2/p3PBpcfjzlSzy6fpz/TmmlaZXIXxGQxio9MmKf6ee/xKTtgzj0
AUhiGiW1su7b2LU6TYzgF9RxRU1Z7+TuC/eOteImRwfDQVZ3Zsp2WE3AYAuE5cSEXtM0r/uO1b+T
psx70dPLnPwZpyFg6zzngXPhoySzZCnXTgOohQ8GNc9V3ttZdbs8PzX08xOgaawVxHiCpPue93wB
7Kq686s4DB5dmRAxxHWVQt2s5eufe1vsKhhiRdAnFZBnYnKQKv9hQtvGlK4JMPVI1GHxReWWWal+
Q9DbC3XG1htVE46O0FNDHqqb2jOYFxK787f0dY3xiaycSlOXelYt98651OX7uX4H9kHTVjjsJUta
aubDTu2gnrvNL+nyQPuh6U0ieQog1tf4JpgvXHNCzGLsLVeClhXt2ob4G1BrcGzVvzi0ouRYO0zR
ROuL6WK2aIhMo7iQWyirh+BwKLMMwwUPcM4yU3tAlsfM2oqADkW7d0tWTXeDzF4wvDrU9b6Ozbkh
9VEraOUiVwFFFz8BHYVbJ1bLxBpDtlamoactu8u87J1J7ORBvTX4EV5emQETOeblGiBtLsgpi2uY
NDHugDbMx4D22MvdQ9SuIpgBpjFvHd87o5hrW0XkFisrIaGz9wNC5CMcKKbJCo4sQdPb1WOiR9AE
JsXSiHjhBrHMxj8UisIAgr+epjd7KzBz4YkLBiB4rkDn1rZNOqoj7eASKl5IDnRQfrJAeVmnuSu/
GUIWNjufZKFCa1JcBwoQnJ4LdG3/cZ+Et/HINK1yJeWXc88ESKHAKWXroiqnxQI61Kv9/robaByY
IabuUrYRBEBQkdP4CnO36OokgEYlnnfeZrwWmATQae9UX+4JU15e4V5C90KDPYZZJt2+YK1vSBCT
alGpVUIaRFxk+C1gYnp5zeipVZWgTZCepLOhgdWxiqhmVmEuspfQNA2k1HFI/cFIByxlWTy7BJAE
L3IsVH2N4dlMk9O64BKY5aaWTX0OAPor1A2zSJdKCYUdkTxaWoPxvaHgsX8z4mnYhIOXo+R5zws5
t/gFUB/whqKqgDeXbzg0jSXRPV/Gxs9k/s/AQVCYGxu+GxAaXizoDmW0Pjd/gyu5bDkpS4uacu+k
9932vFaQomFAsPe3btOsvCNNFDQsAMKnOqL98mdddVkBs/L5Y5KW5SA58+lI6yOanbOLKIkpifV8
1KH3TfBcBf2Rx9zmAtgSCoIhfx/+zfsJ3zzBL5exO/L0rU0AVtmgxIFd/CQYk2DzNtZwzBq1XDYv
+nQX39jajqFlZhaTWQ1D/ye0gfwnKc+rQsKYIiXt1Od3owrVXEQ3AjTM089PbKuMrH6GKp1zONqa
yR4088SRam1j0GpyKUhRIx4AWOQD2WGGFOd7b0+nVr96vKWqpwLN8kJPl2jGJzYPdy4dKttGYh0n
ew/omZeHyrEeTDYkaWBViJWZ5nHwMFim01v4VlysCmr3rebPTSgVMbJJocYSwm+FHN7ZtR+pp6i5
57a27GAF81U5Yb/LcPlmR2z2oNMWLLxIjxmbBr0QO+BRPcJEu6T3dNVLKM0q/5VVmH2LRtZHjYfQ
8Pz9SkVC4hzOXnaS56l5819q6GMKxmGxfLD73uqPtEQIcK9G6gf1WozpC93sr/PY6zg0Gee1+AXg
4T8BPSjmgQTvBiIvSg1A1EPtcya76tUZgKIrFk+6GPfDc3UrPU/KbyFkLtI36RpoePSG6OXtx3qJ
ILkD37Q6dUKMVS9TS3v5qQbeZPiHhQdcUr2ygQVflDI4k1b17hCP5XdobCLDiCJJ9jXUs9z+DCRu
W3tybd0ennId1o8SxjWUepjBA3HYEXwEtbsT2cIUDfOoVejdxvemtoT+2DTOJ8UPzvSbCV2ovE3F
RBS7+6ncE7bBrQuW6u+do+KYo0qBB2ZOLIqYRurIKyZS2QebaP/RWolUUqgKsbpwQHhHie5WnDux
t6bnvjxkLxKgPndsV69DABMV17RtJbOtE2e7JpgGbSiwffJJfynakFi5LE0Yw5wyqP9fHLOK3x5a
Jpx+JdoBTzF24xtQCYwAT8GWdAN0yOJFkKj1DYkaothzcjLEjeh0G6l/pQTQkAh6PcYXxcvHZTUi
ixTVDzVkc8ZQA3dnR8rTVzQmdRxv7TXTD1ouZRPE4TwF4exqIB+X4gcCAzRhAJkahp+Md/JNMQQB
wBXM6S4IWdJX1GKPLqZ7p4hJARWtSgEXW7ZMouVvlkFMksj8s5YvJ1GTe5A3SafRqVEGhOGQ1UOg
J6Aw37wQkWQ7t5ojf3zTe6ULDaek0sk/inrCy07tX/H8l0TwpSf1HcYnBZqHIB/3OKz0GHVDiVqD
k+uecSEWokN5inEQraKfhYJx3fIYTw8xjkCA2HBw79U0t0PbAsmpIlgf5qnMhyeBzWtlOz5tP7dQ
JfSgO2LM6stOmV5JUUkO/0Yc0iuG9cv1uFL9Oj4TB0dI+4BWVQ7FtUxlFyoyWc7F3hXEb2VyInEg
jNa/+N1sNciTKpqAp5zbV0VLL6IoVs46Z6Cq4i3piSITKe4FpwNEviunELJjUa8MjMlIiKxItfco
iTdlveBue+S0NRMQXgendAKBXUGdAWpo7f4gNVS60yr4Gk6IrQBqXicX7MZuY3G0/8Z9uf1bCRgH
/mabHhw7uOfLg6e863lSFB5XJ+tQz4Yl7EVUKHsnRARyCycKUFMe6/uQgNrcfvRumK5tIbiOHOr8
1i+AFdAs1iMSFc81DJIsZMVgZMUGe8Fg8r3uY9XblGGweejRaBxTxCDQkMY/cOG5M6pZUzOvTe8P
JShoF+bsWlkZl62ASVifU/NhSNOkYEs3Pw9V4mtIbNunnJAXbTMKUBbqeXzYLZgWXYvDueUZa7b0
e8eS6TyRP+HHXH2jU5d1cTthv9cxsCou2bQQGyOdQu5Sj5+OhH45MNesoJsd7C/ZZIrTK09hJCSg
LidB5pPPxnftv4zWBOQ2mkASWuD+JsIg/Pz+/97cEBCZr8H22qjaO6MYQ0ogP2Wk0emTBNkSve7+
sFt4aRgPBJtN2WtPEiX6KJBpxcOppCFJwZYVMlTcOc9UDHE1jbuUwMBXC+72ayGyHm7vuiWGcv/1
2PJ96Y5vMcxeAZyadTYZxMdRG2TVLAnY8O5XuwBMPyGlvnIWysdK6Me1J1q2PI++lnRRET7UvXoo
3JqIhwcz3NivfE2DfX2jIyCoTVZL02yGSjJBFobQ2xEP9cS9dEIJjcA2bWdeiyXRnYK/fxVeZe1t
kdyrd7UCes8fWyTTLEoCNbtKmu1gN/jzcPDvmhexpWhziiTLimd5/0JcCayx0y4jQBs1xe2dLhEm
sXEFN1iEaaBXxTPRPQGFoJuc6can2tw/VosuRxrYsAVccgWTmMcUL3LK9pymM+OpYIUxcU43yT97
l3QidM4FAw+9kWdy7fHVMk9GprxdtbQK5QGPCZIYd391upVOy89z1iOqYHaJiYc9ldUnyh1cLKp6
PXLEWA/746LlTmIlo2tvpI72mOUeD2JNs41heljmYPBgKx44ZDBAHthSM5y5ii8XormZr1Xfl1Az
6+6NlggcQX2PKq2/dSbYkFLZmyFpfsDvWleJc28shkRGRLsXq7gLLDJ0Sq5Dfpn3s+6ErAFVc2xM
HMh13/BdV9xTmdaRqyIjKTB06+yO74L6b4SuPjZVd0rWo4Nu9oUnpHXPi2m3RDWQtpIDcI9YtbeI
PHQgovIMO6Kkxo6uxf+tDQCa+JPwpdFpOUwRqMcUXKQ0ZifYciIcfDwPHl5qoIR9QiS4Ri9nrLdq
Wn7e+kDyhg0/hvso1x5jC1KtCWxlt0dzxxMXgD9pAErT8CoHQJV8pzfXbjxgAyTkHbYZqImrcT+l
94y0FW3LXVHAPSWCC0iUHdq84/J0V5C/84KZBRzhxwy+FwhPwCLBmgb1l0yNZ2EsDc+Uz36FMSDU
0QqeJNyzmbSYKEJsQonEs3qYEH/saBU+RFQoBg+uBnzEMJ8QQKNQXEvhsQYrO7UHm8Xy/3oE7bdW
M8qS2XXrUGcdSLEF78Xgj5M+bgviKSSpgk0baayrP0AzFRFW2ZjIPrU6h4Fa3zEVUD0fd8itEanX
kBacvNAgt51IkjYNCyKuAfPPwtcYtDej4mBz6ae8Wjh52yRzikbJ55NgK7dIq6gQmusVWX6eRxRY
gjF/VMSmBnW01MakZn9Fw7SdlwC9gDRMGQ8CbriG1E+b2GJjdT4TxksZ9YyHnhVe6S8xAQa9ZWZe
Q4dmOmx7acJWufyWVv680C31kgnJcrwriP+m9DXkLQaVMwVWwqwhs7k49UA9S7/zuHeVgyR0w5PT
HQ/1dPtK6DLOpgfrr4hQB18wxb9nKYddrF8748J6Jl0R2o6Y59sNBCmY0kRCYMsFkuHbpXqGkLVd
GTbbul09MVOYnhnBqJw/1GyRBN8rj7LNh9khECi1Y39AtNyi4CaWAUfT+9hadXQfTvBdbzetLFI+
DjD4Sk+7Xxc9OOTqeLk67UfnG3/X0Pr7SHkpXYD/DOSBPu1YexJPN0Y2sTi3eThImt8UTBMJykkC
qwEs5qGYt0FISSm/9Dhu9kQ4IhXoLaxLFsuhzsyLZ6CuEFiBHNct/rj8R3uSeb1wo6lKYvTs+ACX
FeCwuRy1VYP5ExweXJzdOWdSQ4x+6dh0aO+r3VKYFym4TAKGfgA+IJkyp4NoLuOoo1Ud2ly1P4Na
JQtmcw6G0WSQjzT855k6UUu4Y3QZMnZjgaCQa1PU7s0bcaS629UWD6+eBMO6vxjYQS/475q5qN3u
/XMkAtdRUl8toE6wgKoZTj0WXf4arlSE2AIhxws1oyzd17GrF0cngka2UWrjS/uxdq+x2bHML+Th
ZI+9jVCOywsAYynvQgIOJUMNd0rrOocre9/NPtZRrdUQghHBfzuUJFTC53z6oWPkblgLjtL8kBsM
HepgCuo3Yb9XM42/D2xXR62AhKP6jxtOPcdHZ8sTr4adqwIO5a1WQLTckg825Shc+bVFvrP7pwbw
TiDImc6akPEvouqRsoSW+ltTvvz7HYdKB1Ygr37EPe6RcwDqIKAr4ALIHmk7dMXw8DvxDoj08MMM
yX7WkX5lOaS/0IsuTNZ9dpS2fELSU3GMjVhZuPCzyUWaRNmCl4QSQ76gf4kYsz5D7LvDznEva7wC
fHYqI/CK8vVWP0IRVNm4FT8XQ00nXdrjzf91VsIJ8QOnLMsqpYnX91OipessWijusEr7MQvofkPy
awVbBPgHJN1HzxP7YBAziMvfOLsX1Kd14/D587fy8Mj+VUw6pNUqv322ZTyvTaMuRMTKbHFqxuYE
9KJmO8MBj0vNm3g2/fpYYT/X7afZ1yamUvu2E/8Lh1buRGh+s5ByySsK49OnuxfcuefjyExbXYrL
7i4BzUtKQDzQ/3uTNZNj/Z+zF+VtIcpCW3L+wACrpFKNG6DlDuU0yNSlg8dDSOt+/y7fVorKn0aZ
iuzdJUz2TQUcCXL+6tLqXkYgDwAFqrYArbezRIfks1rZmU4Px3y9mr5N/jurxuR5PeK1lN6CvoUV
lH04NGs0USqZwAzYzLsxkJqmTVAxfR+NRMVsZBxpr5d1tHPn9Xhyz1xqMT0U3jgNxGtP/GiF3SiH
eOiFxMy6wXSF8+/cEI3KYJKysuasYGpiGzK59rYiZv8hftGruYZnjUhdGWzV16sJ7Z4nvY+Sb5q7
bR3RtRJJ3Went9AD/NdaKL8xY8Oc9dj0vfloj9+CbrrNXxI5c2IzC+gDxkKHXKM6VGLy+Y8Ta+KH
r1lfRVHCXHHzBgKraA+HW52f7CKH+EDVQKCnGtJCVSqZhU+yFVC1vQVfibqHAGkMtV5qS3qUlVxL
+3AjGXAqu+Npx3gCHcFbSIRFTwJDKcQo/KX+BL6kXeCKaWdQSTu6YeBeFBWo+UX5dMePlKqLzXkM
00aU2MWzGzZ7dfNwTZuYe1/DGbpgZGo8UZVR0i/PX7Lnru3akJnQHdpiu6V3gC/6vSPdIsdX5nT+
xPmvz1KoRO5kULjx6NT1xpSosW81PbB7S2CaBceT9++dKzWF06LTBSEsB4temeqvJX4ENlxkmv/Y
/sGRW/NcCx5bYtWJQ1mBorxWCTbFawynqq1BREfjBd8pjWEvPKSpfxXSJxxbNoetv6ROOahdZDvt
NhCX5Rmo86lOgCRpAm5osEp1U758+fMZnbDonU7DCXaxUxgTOYH8b/SpCOcFsucWkC+yzD6DWbBd
JqfhKr9pCT9ATxCYsDUDzZC4FS+JoA74P18hDFuK2ZJGXcUdzAmwq1QiJo7nAgrxGPfNbR68BZSk
NXm1YDMI+iOLoA5/EwqUaajKk3NdKCoWHpy3ye3hW1kufevrouBkHjlSanszv9ZrjnXEcl9sre9T
hcO4eXhBipwKb5+bqZzEOBvZ6bdKdsVOEiWSmHTvNze+HeQQTz1cHgjue9+0gUFXEfrCRdUum1T3
skSmd1eYmg/T6PJRzWtJnUNmwJmlgVieKdbEpn4qD0n7H0nk5Mlvqg8ASwZAMNcK1Oqcfs5eCQpR
zfvGcl4Lgj3A2jaH7enUfFpr3qwNJx9ruEZZzrsUpQ+/3jAvFsMO91AV7xUcUuQqCZB7j8Caf/+/
V4DzFX3XWV70RumXYE1QFp1fX+bwt7zsHpUX0HvSCP2ErTD5I0Yb8ZMeNtN6bmkKKKgvS1rWO1gW
IOi1IDUyBvPIMPLM3x2ipmL+CWBa3/f5eWmkCJwgBCbRNs+iF47wJKuBy9EC4MjKTJdcEVqoJdoG
BRSZtiqsd8t0a+roUyrSG3H/pKhdl9/k2gv09we8DYqZ7JjJEmmEdFItdrOLJEyNjSOEgek5xPkW
kZ/f2vkuJ/7dJnCchx2o+/RGARTNHJHOTOob4wuGGJlh8ZBEO+poem08aaBEdGpAFTCjJZsowEWN
iN/2carwkwms0+GcuSy3npPpB3SQrbYFvVhllJ+cLbuGCPvxRjPDEXV4rhw19v6DKItmnf8awrNc
CBJ9xtrFXVMIaJulxC3ldWcL9X0cI8De1fVoThWIG7vwcSbXUQEWj+T8Sp2THH10k5Pk+zB6vmtP
5/7ZvH3WTdLfguRqDH1JaDBs0NHydncDoFV8vtnABpM/J5KlNboJWPT+FGUoM8IscIazC+U+pVZz
8OkzDC/eo4CBsosKR+zxXXWbRtzR7izKUxf+QDvaBwLOOIXPwntQv+hVkba7U9T8xN+W50VVKvG9
SteBUQwJSrDP6E/K5rcwA6oZF30YTKIa3/8DCg5QsS4cNNrVSJFmD7jleGrvVEbs2oIRyxCZYbsK
IXlWZWm0JIvsvlKvIFlV16nWsyLHP9H2iV04Vw6snRWeSiFVV9/1kTgjT3hw3W9pri2Z3yVpGHc8
MzJsKwD9kpwJt7wLu4jifCf05AjxoWU4cvJqw5Ec4zdGchAe5jQQW8wdYJtjhhv3hATXO1ewZQ4x
JRB1DIgCoUO8tIGKdvTG+u5wbOeoC0Nn0yF2H78VoiO+lJVQTZnml4d4HlfwIYSAHTmoycpzeXnW
XgUzDzOTX0JV/DT5rE3EBfnS7cysDzilGEYCBBYI9ENHQK6v6pvywuyK/lVqNk8t/dNZxfXNg6gV
wqHV0PLxA6olQm3FiGAxa9faoHRzOu4dC6EW5Mnc8aE+9mX5vPswCe7pYBYblJNvEDj7OV89K+QD
Yp9MKnQxBazmdKQLB8y8sWs6pyf+89230t8YHi1Ubmp34ASOwZ0vBq/DStNgGCJm8lhKzJ8d9Ni7
4lAMeIVyvvGSHnuZhYBsqngkaaQ8ffC/X/YWhouGsekAcs5FMa8oCf2NkMoCIWmcETNvYWkwAD8f
szjHitcU+VwHi4eEIjwk6VU5KEHOmudMfbV4Gmgr2EbmPgX6NkYK3Ruu8v1H01BvG93doKPHQEWz
r0YtKPYziwIKc9KZ+2+onIoRMDxztywQEzJD36TLWEfuQklc9PQPZKsIB/7Ac6PoBM8zc003VctK
E/fWUjMcBlZaTm4brfie1GUwKBA7MFzgCO9w79P0wP9RP7vcjldb0zj87wtTJaKZsVM8R6u5Rot3
hH+QG+PeUbJuv5+vCOjEGPCXeg1xeuWMSSjrP8wFLQm/qlNq9q7S3C6lSIrGpBQdLBW6ib998QYN
xuFnRBHmtvbYdFkIu+X3B1K/mwn/KITQr/BOoZ4jctF/iBE8ZSm3Ugc9T67wgen9MLh6dsezmSSN
vgbLXgBC6eldTn+4WnFPiiAHA37OZ8Jhn/svlk6OymbHYb3Q3w/QHxj3tt3HE7u1lMrZRClxoBF9
HyUifttFe+QqvzL771tDtR4xf0wbfXyjGGkkNnXuSX0ZMdaOv6ZcNQoC+beqR30Rr7bm8Um0ePWP
V0bieQRrn0bk0GwLfj4A/iNRVQnU2YUruhj8PkFpIduSsPXlZKFo5uXId4Ybruyn53umxoMTHdv5
CQJEti7Gfg2eSihUyccTXpSrBFG7WsyoxlpZCQ3zdy8uKSHGBUQG/GO9ykVma/4+3gFjY6Nc9rVB
wHg4wATCjhUSMklGGdvQYmbnG2QPgFjaEE4UWzTY9G2pLWtT1uoYY2jiHnVVH8gi8OXt6ipQevLZ
rxqR5zENc2myhigc/YULt/ZP4Zx5jG+DbflGmvwVKcncIH3hbRI5xlrwaQGrRJ213MZe0FRHPCcH
bosZMwfRQCj9djYoYWffSfGcbSk8oM4Y/GqJ+7a4QNXXs9raEa55DFukZEdoxGlwsMQCMrKz8fpr
HNDi89B6jzHunzwg7/JmdCe4LGvgpzeh9iIJv2q0V8A3RdqiFsD733tJzaFeTlKHXEr+lbD/eGfE
Rh3Kkh1JlgxL9aZBiq+eEzhwhCkO7HBO4alRINAuijAhDgz5Q/+Gg0kFNueEt6cZJAPzzfJlRJa+
tKd2k1eS9Lbqnpz2Ybmm3hSmJpdqmu1u9RET9VJgN7Lieya1bOiNbjXgpWMoQUc2LVSY5MUHokw3
T+ys9JMATKe8d2E+BhzNMZXjqTj71FkelJvYEojr4KxMGA+Ma2IwKNPFBrSZfOMIhZw4KbkQwi2V
rN1XiYe9Q2IaUhjIcAO2B6dAKe/1Ug98mL9x5O/4Hwxq4C5NWLgZmy5J1MEQOeQICqGNyEss3+4m
1rYyvi+WL/LaMTb9pq0GeYiTf9VKsX7oQZW64v6rzJg21KZIkPGUp7uQ6LMRIecbfQfyUNkwoB51
X1BsX2Qo0v6ZZzxRocGbGYbWccxLH2ThCThnyV8dako26SCrl8P/3H/H2Nn5HUyajutmO4DoQTnm
jHW6vUqyyfYhRPKZ+7PZWSHI4laFMBBa5EBJBhpTr7LCzp0W4VqTxSrRX9W7GZN1akm05s25lyl9
KVX0Dj8K/r2eGbg/EJi2/70H8hDYjw/TafslvloUnihi3bJTbx4OBIDDEMIQ1R+Q9dzKujDbM4vk
xR5N+FkRsVHm6j1aTsROknC0N54wv5l4THZj4samHHjZUhOSprhVBKkqlNSTAF3BRxxrZRfR/ycZ
OoPtN5J0JFBWiuJ+4YKR/F0+afD8fQrdbzS9Mb6bNHKtfEegNc0+Ac4l/4YuGgLcZlpU7KVNZqKJ
9cycW+oURjC2O8HGDQANyGEC+klzJz6EaDBYzvxOCyutcJ+V1BZ1fyg1tR1mvI0w2fWI9jEQHMIM
bID3AQAiJfsOainwtkWIpfTr7Uwnc0gilTcuJmgO/ADhF6zQ28GzenkzuuUuBJW9n9c4zcRd6EbY
xwgyjkbq+7D1zma2UMcgbssgzRXHNfcbl28JjLG3twrqfMe2nXYYD6Hn8TAbR8SWrTGn/S5bsPYt
iuhX2ihwtrPxJcP/x0gg1c5O9a1jIOXrvrmfvpx9MU34nNfH044lXiz/AHfVUE/fzZXQMDok/Jpx
uD5PRYxVIS+CGDWT5N3kbmOgJbHa7lzFQhHC+3+/sOScR4Wj08SgVwaPjSzAoA0aBKXnQ7XTNkWU
LcFSnYvOSFvMmM4Lir8GdLN7uyip0RtJh03itUnej4xhYGBphztOzU5FFdSPE59yK2HWUCde/PRT
EclDlmZ3liGYEXp4FT1e6ZJlgBICIYHreH+ntrz3lwz1kprBHJU90/+jLYOXZyTWzsTbgEGtQW0Y
EoVnDKyHT2m7BETYLsIcwBCr1TLcDg+Zw4WKH1TeFMDr5N5kK5tyv8Sk5BVtYI+tn3/O7W1c3snC
UeXVKkr1zD3P2xJNV8OoqPXRqV04xPatsB3IIalHxYSmM6rEhWLMHJDf6a4TFAQ01smo5I7HSin6
ChcnvfooJALiqySymc5lZ4c6IWorIkPHNYhDSZpmQaW5zST44XuKpZiKMiWhHkRV9IBMwYFYH78p
6DY0M2cyVUuOyLaT4+Fa1R54BK8U1EKfWE4pfA5nTkjquPCT0ckjXCFsc+gUo4wOShed14ghMKzg
oCIMUAh2y7jMOE7YMJEdaAhS+yNzuBiJEVs8N5JwtVlVujErFDGfz7Q+A/vv5nzsMDiAxaXEFvl2
Ql1LZB2YbSEXU0E1GJGcUcSX37tdqBFui5QtT62rBouP0tCq6FbSX1GopNA8LLBCannHNO7mKHi+
JJnReh6No7Dru7Yf6GWJ/ZxGjbF9AVBPFmf2kMNEJtS8SdWN8Yd2+/jbj5M7rwR+rvhRC7nkA0MA
/xOuNYDJHZssYmC6mpg3aUA1n7qsjdez9cCBLOMBWBBf6EfMM3CP+3alWdaF/rw/R5/TEiBnI/S6
tYjtcEhCUnmAyuvajQL3ciB2CeHqFYf7EGwj5MiEEZ7M+MNYkLvv+9zPBqKDMuLuz/YiKjEC+0Ua
/yXxbEiA2kCcGCoNQoAijSMityrZ4zme39EDL6zzW4wARgh7uuWI1oMnkTBs31ZDNHkDuOByRdZV
vOYu1jWJs9tW/r9UuSsD+LzoPulkpRM2DteOclu+wcb/YzxVGc2YyGPX83Gp5vF11xbpnpVVDey9
CrcvjMYE7HhMWKxGFflXDNSX4m/JfI0D3Y5GKmlBCHc9UwmbnS0UU4lIEHvEvMSGqhbuWxNt/P8p
qUu92qkw8zhsDtiLDERtlrlQek+/8Kn3XP5kE99AzTAyTC2Z4ATNU5+dQK1OiykndGu/kynO/PhX
S9WqEEFBrkE+rD5q4gQ4O1LmBQLjSxOmXwjyX9X03l5C3D05NHg3Yi88xRP3SU59CeWCwxVRtxdN
jlwJ2nIweNVmmT0QZaLlshMTitetAbNabNnWMjkji7/fR6wBd/yRwO2ghD2++BsH+hXapwi/Lghl
r14edQR8uKwvxSCLqVzs+ur4MXc3m3aYELQjsSbrg6CD7FgGa7tuXAzGZD1jcMew4MjsqSlbpG13
OggCAI0jFS0IL1ckNV065Ft+YuA9xUCuANtvA7NIAnsv5izoidohSQmIxgJO3Tj5VeRItibo04fQ
lrSuHqwWSo7nW9j5gv4taJk46pPuKh5j65LRqP75Y87tR9Yr2pP/lKFqfH7Cx4zvwDVUQZOkdVlC
n2dUxVJCkxej/jh25g3JvNa0FJTLY9kCxlfsw2J1HN8rqDn8jsZOdSjbqL4C7BWSIAwjqS8HXggi
4u4stgxLDvXIqYQb3JDbPQz00Ysrtdeimf7Rn/gEpoH37ZfrMoLWe7BjxamSh2uHt/RypRz93CJh
Nm0p9ggE/kW9Vuh128zuJf84n+FznW41LNoEFV9pII/XghNNWxD5IcMVrRTCV4uZX2f7T+iVyvrJ
/AmhGvCJaTNvFYUnMkt+HDFpBGY0kBLmEDPyeLO6AXYe1Dv8I/157OXSgk0SB8sL6OOG7vofKRZV
mJyPfchbyDDLC+beAvGB1mPuY6bDKtyOmMe4JF/0g4j5a9l+/Ash9b/ICYuHm64XqYRRlbBCoTtL
aMnQt7QoFmgHkAiIaMwaZIQzPCe1UlQcmxjZiAljW1jRdmeWqkPvVd65ajz+RgWgsVVwKi87BoSl
KBgTmOg+UOJSXjmQWUQiwqyKx3Twmud3qs0yTdgSinM+gD/9KsD8iiubjyCAm5yxDo1P/ifuF8lm
0qX7RHyHoDw5QQl5hk0lO1egwweMr1o3Uxr1sDl5dpXBcL9AisnAl0pMMloKuryFz2LUkp0/5J/S
NSFbHHq4qKYk0KXxXEvYJC6bm83Z9FrYZ4/9K2yjs4CKSF+11jxY8dtjDyDsNNS9t720wgAxpA1Q
0QwFHi/vUS9uxn4oxGahb7Pz58sCEyqzUHsuOT5N2nBi4lsz+EkfFKeY4EJ2wm4uz7I7pAWwZudx
rzmN3VEGRNzt4LLRgTdq8N/IL5+KprIkk74HW3GNXe1UrAMshesWA2OQ34Y6iI3vNT2zh4LufbNe
mV6YXruEKFhkIfNDF8iRido7xHyfF+vo9f28kOXw9wjEKGwfXgDFAs9x8rjzyh35IGiluLRdaWiV
iwK3v0RyjGlqi4JylkkBNQj2FMy6FxIEN0FPez7BX2jldgWZKDtxcuE+Behq5T65grG/8TguKvzY
Gp7k4/4yC1zvIvpr2Dm7ePTCCuhnmFj3QjTbw/bNOs8gAq8KJVZMOMmDGA/soJ13qSMSfizJH92h
I8nEZx11AhfEMrbUTeZWq7mqr9UsdevHI4IAND+uJwZFDyluNDeoUF0KtGfZaTf6AjuUQGpOJbdi
/9mm/MBMTLLjhHrGE6BPoZjp5iUNucVYDIQHK4Evi71hWYsU2qXmHeauUrCbF5El1rujk+6JGtQX
6iqBoZcOVI52MA2X9DFXvUfZq84N9K1+OWhcwJpdCTd2pGE4FOHd1oIN00/3yHQN1mSPTpeyGhn7
CMKXsQzA0uJYIhdV3zvUReE9CLzXbU3lS/5T6ibOiqCYkGskLJI8+pJZV165tN5oEvh/CWyTMUhb
+1EI8sV3AnhyLPqxtJFebXQaAR7/TDfR65+klW1XexhwXH8FVd/9Ttie3s2AwIqPTiQxgtrSJfDe
00N55/St0cTSSUQDYDmRLQLJZs1zuvaohgbhCzQv7VBM7OR+q6E0DF435Fo1nnQHzMEd07SDzSMM
xGkjbwQKKIGkkhHpS2i5x4gI5slhNCxQ3XUsxaZqf1RLZ/YsT4iMgmrLDbl2Xa6eAz+YsnP8Qb6/
aT+JLh1Vti7F+knaQZyV9rJuNhs22vDH4JJ259DWhanzBxjR5QaHwUgV4YJNYAYM2sY9z15xPsAE
jXOU92Ljp1rm1f+rPK/2FfMIeSejIVISE8N9hk8UPURT6TGZSbHdgEAUxBgbL/Xk/Fm3k3G3xPCW
T+llFwf0/fJpxNxgQGPqsCtJ8vyHG3yvPfJLtdb1gh6NaDbMRjOGJ92IEKsUfq9iVZMKPfUG7RZg
7elXBI/3613Nv93WhkBirl9oxLL+BtUXKmCDHpmALunBNelL5KTMehq7lwv2qIqy5T5VhwMqmgiB
T6RgRiMZGvPiPswY/TIGv/5RQfDy2uDeaWB27uDMZLbWgz7wCAL0uBxYk6DSnIYECd85618nsAQ8
5CR6FJkZ8Ct6IYJAupZfk7e1nBDfUTU5KCMgH16mZttQo40H5Kf6EuXd2Tik5WRWPim3Ey02lPDQ
fqMqStscG52YCSFjljG3UojLicfGgV30P3gmr6n0kOJAQJFYYUysGTXwctsvVVVN3likMjcA17fF
FAqMTWel38mUzpyP0WqwRKHStEcwDgy54FuLgsEJXY0zwhCL6342jICEt+qZGGin0BQmf4ZnJGg/
+jwDdc7zRl2iiGSt0dCGEfIRA3rQAKPEd7/2DuI5MIEUDLvFHPuJ6G/Ga8QkhNfYDbLWnR1O6FOz
xq9OuryeNI2g4tqpwamSsOvq823QLfKf2wnrH14Sk1umcj/vCNy0n3CLHUN/4JMw3wcbYScP0n4U
wbMGN9VhSGCqk5bzOBmOBtjsIh4hi8U/dH7fpJbh/hbKhaEQl1rHw928KMVk33/wMLtDxhNM2sXJ
bFxwHUZ6NE5bLIjerwi4zYkmapN3LfqHzVr76PB+/mLLxeJpApIXsV/5jqR9T5sNlkESlYLk+xVX
HU9A12fsCgulXECZJ7m0WN1VRuy8nyWrt8tsUmwWHv2BDRggOG6rGlujQqWbEfOSWp/Papgg6Jst
xDALp4lfRpr/O8YO50/mD37cJ7amX8+NvRLp2u74IBzMJqYtCXFgpExQh5qFdqhcqIuwUgJ2KLir
iHXzYeNInC/0v+6kt13rkQ+CmK/Dpu/EzVhjx2KC7ZVNlRTzEcxCfRGw3ALJASmWJlOO16+ZH3IA
RkupL3yJmTKVAGlbbca/Uu2sTPMPsQ5ZWSoqq3c0OB/RPOJGUkAFOOQesYOpE8QUMFQ0AW4hMonw
IWfD1Bb526ec3nGoUKwY1rCHsJsuOJb9v6QF7e7skLB7hApPvNLgoYpyTriPxJD1Wz5gHs//e3ZK
zjjkdmSQQoHVbP+T3FBpggwA5GnrbwkVW5SJY6M5XJDid3nmohT15zIkE3AqZvKaiv/CLj+TKEsF
bCIXLX4IKPU2odzCiOYPYpP0nYFeM47M3FH4Fjo6iwjpdvhCiEKpvbZOsaEGK2slx1lubdOZmFat
V4ImlrhpR6Dnbsp8vZaXPectqGu6u6qcyosXY6WtwB/X9/+jFxC+Zr38pk2AChOfOw7LjuxcDkoo
kxaNSuy+W7oB4uZWspiZr5uwKIiEl/fFcbnXroJHq0DKlRpOQ10SIvPG2yX+cby0nqwlt6Awkh6Y
OoG0IYBY5p1AvlrLISHpzSQqlzmEEqwYBcO7tYW+qAlPE9gdYXEUk5zlS6/kK316/W65MVpIH5yz
PIR6pH3z2gRerQPkbam/mwTncIkC52+s4wbXI/QqHZbMEcw+Z9hzowvOB/4UYHQR1P2DyVxHS3N3
TuAdQXcPtDhHaCo+dkjmY4tr61PnzxMujaZxKZLYYcH1x2ddXXIDhOROfhNDb0KKqPua4dgT9flh
LtUCpxi347CuSdd5+nFezdEdlexKNDDSldU3pYzBFvfs2cIPyLvdbedXQ3E75f2y2jIW1I6sJfzQ
a6N2jraO6E6pFvPXqD6CVWZhNHfuCN5JiSighPKvxVCMYL4Ar5cejBkNhzaDdTojR/OF5uhyYNXj
+BfKEiUOz7KIp6XO+B/uBaK/DKyo1tI7IkoO55rMXhrdsEV77Yk7eLt+h0Rc9l5/THtcc3r2AZUo
W1IHgxwnnH6u9iflrILe1zQ3N1GQZTSohF/9ShYR5y47+1YOWw2+CX2Or2UbhJv9sjz4C7qst5HZ
4eVakgWZMJeFq1mVBfiB2CKyREZQJ0P0neEH9EdFjHy2CGZ6NvRNXWHnYgRDs4C3VrqdwvGSnU3+
ka83cUGow//Vd7tTAkATARmjRRp6RmCk5U7jG6ugtGnOwn0Eeaue541qogIgadV8m5YuMijp/Ejy
ZCZHcAkcZvM7fe9H2IN036La+ikW85WvHZj1IaNkN4skTaGcony6v73zcA+AGeALwod/K1a6BAC4
qN6/FE+AEUmfgZ/F42+0RscCVUtDVJ9ZI+w9Y0TkZlH8F0WKLd12EGXgeuTq7mJYfzlmB46SpksA
Bk95fy6QBCEqjwuuoHjEAMmS6LnGbzqYbJ8SQmTHf6oWI29lljQ8KsHBGCRJ2KCy9Wk+suIpmzc2
FhU0c7TwGc7Gk0kMPTUz+k7eTL7z92Vqa39mNNwhFnxGxHzQSdf05+OfChLcHFHDz1NmTAgxzL6y
b83tBzt3BeO4MsY9cnji0wWtlBuWHYkstmT8kOmXNfmVBfrVs2WwHhbvHi3KesTIY4PbZMOoai0d
BYW+gyml4Iikyy2sXqthvqEmO5208/fjQxu0WJkJG8hfD5BeiTKruVwnBtwWB9HRQFmp+nq8q6Hx
ljdVPTUOXoi0Oo9gePh/IesSkzbvMRLeszmOEgRz/BFRFTNhupsTiFB0PrAgWn3jqT5IuRTftyBV
gIzGxwj0MGH6+nxl8Gk2HvjcmmNBWZwVQwjzgx1X1nRunRtLKOvB2LUTIj8trYHgFwwVbMxkZg/T
V78MI2EM8XFf3Y4iF91VmCgBrDoF0ihzgLCrnOMzzjdN6wVzH0OXsWrvZg4X6fNiQLaAwXRmXjzZ
da6IlJWXQ9rESe7Tt1hpKED3xP6zSL7iDYq+bZqmZ3aQq4KN/gjrtc6mHZFdVV6FpMRI8dBILHzA
ymIelUcQYUm6xkphZaGQt8Q7XYB5UMZHoD0CwfDakmvT0fEKbQovuGvodRjvFcjcgG0SPlM/LHqk
Os8+tAZO9+0rEM7+Ws5zqSTBH6Lh5gItkWqz7bD65DTtyfqomQN5eCsc2IWiT2WKPRz+e36qxPds
BW1YLdAB92A9cnibHbxp4APbx1UGxAnS0+oju+gyq1xmTiSuHmTmclbTI2hB0J52g3r2Q792YY9g
b0HMyJz0gHqGGhNqBWpkeRqJaeIKeZASnFklG6VbFFPHV9uk3bS41udjPpQJGLoow0G4zZF9pzWY
uEph7YeE3O/Fj4r65N7w2Jzw2bFD2VkFDDk8Ixjz1rMoYeUfdw6FVRTJpFFXhkRxze/IkduF/HdX
ZtZJD4pSZEeBdwWk0q4suHZMQG2e3aFp3YqGdAKc1Nx0OffEmqxFWoGrNJUc7b/PYZLrZuB3Z78d
Doqriom4CCpO2ZLQQOSTJubHxLO7g/O8jH4AuKg5RgOy/pshcZqWsoF9XE/Mdzpy+iPLEjT40Q3p
vdk/7NK6QrSpdgZXwSwSJq1nQVhZ9fJjHY6KFm+ZneMu2wRAEGBCT5on8l5LkoW5O2J0Y9QTvuhV
vv1AwERk4tZs5gG44V/6L8/W6rWyZpeXaGZN9uqOAvZFE/RB4eLr3GTndrhZ8I/2+2X3S2Hh5taa
iA4YQe84oq76EPt/1SegJy2PkkbBNz63eBwyzs2H/UWo1UcQ0nyN309TxQjewOYWxm/M7zk1cNoP
Uu0cnO513xoX8QEHu7G6zUq2srxpn9keJt1uG5pAfSYji0TistLqYBkxxs43TYbzxbo/koyIy3t4
u8NQqLDP+9FZ5LetfZqjyLaklvrzuU3gW4taTP8Apqljk8clP7Keq9Z4NS9pdxMZOie458lkx/QJ
g0Mx/vpY6urc0iTdvgCkniVuZCJ3tSNo8J2jvBjjdoR11UwmrNImtz8Y5pfXv5Ue6KZUrXetPRwb
2N/fX9Xnbyy3x4LnH2AaNhCYQcriQ32R4k9hk4rY3tmf7PuxTmEGMuwb5pp1jCXzDsrUAdEP7Rf8
pfxm3OVd927dzKoaSCjS/0Ny68GoEF6wCnfaOWjy5vg7AmC173GwpZ+Fq94NL0mpndN+8Es4PVhx
ngFiwHZ/XK9Rc9cxI11ZeEm51hdjfmVaLu2u8XLdoCxXFNRgyRTjoNXUF6LipftUSm0MoNy3Iike
ToUllUu0vLW4qxmZCqBeoGk8iRbHeLhe/V+IDlneu9lruhF5C5g6BktE2UeW6rh1ksV6JEPMubcD
LuXYa0y8WpwvaTD5Fw6S811SGv4BbH+fjb+t4ACDixQ9ctvd/h7V+/JTXGifcS/kQzj9sVAo24CM
SOh+jI8mGG+RmQclXHVQbvroiX2kWRzIEjk0qfO9xd+zhpucvVUmOxstjaDK7LxO9nelvJZXC5I2
1ZXlSWK/KMZsGvTZNqAZq55yJa/STVPEXJ7DP9DWkJN+0geELBQ1o+vwIX6KBxts9vlVwpI7HU8I
IIukzM++HINlHUf2lHGZHN6Hvaiht15DHyV0hNDCKFV41MQ57M6YH4e/8BXYhvNzWS+LFY9hLeZJ
3U9F/n2vkDZwWgg5KLcDkEcMw+rGPey9UZKnSNmQFOoWWPnENjXeaKAsJGpOtNEP7oXwTiH2B4+g
ju1A41aXTRlQzfj99ahPUrgtUp6eTS3Bkf/762abJn0GKJsTf+1jTPtGxaSdKQsuGeeuqbtaHBy6
ur7jbXTlEjeALCrZ5BpQC73gwdR9b3Ktzc5Yj4Ckcs+LJW0NQojnYPqVqobPI2C0eLZTS8cH66p9
JfEQ+S0cImTvnLiJ3qG6u336i1Kx5buHIHRMbvehHeC1EJFk6seCPEJgYaxZ0VxQFA+yu2ItyAVD
c4j0barrteDU69tyOy277UkQSIzZmIpjFAqfuiuqjzyitZQdN4eiAmaPDT7w7RgJvnI9uc48Sg+A
YoVL5VQ0U3P00OPCeQzpbKJUga47yKEQliLgXNK8uQuFpEMndjyAz831h5Ep1ZauykAFmxTTEnZf
UYnXTEQHfO+EKlEzeiHu1JFLxZtqUUcZU2NBefvZ0l8an+6buQ526acayUVEI34pHp67/EgKkSuH
SVDVZXKRSRCZsQUI/czQaSntjc7zyBIRxI/9to1zax925wwE/xjNNz+SAE0QdBKfahPw5XS1Iu1O
9C6++42FmTQ/dnvcklryda7mD7LoLlDtuLEx4N69veMFDgbs2naNFD/C0+m7GQ0KG8oHN/QkALwD
SGIaO3dNyZKc7o9LhqdvYykAaupqe6YskKQ/zrtzYrnhoaEYBiPyzOwpzy0XWVGPBM2GuivDBLmD
QZ0qF8Z/WnYDS3/mWApnT3ib//xG/98lGc+AiBvmB9KC9f2jGSXSiSqNyyLsBaUKboPl/nXgUYrP
/27Tddqpqq3tg9uX8Em5tG2Vr+7S+vnD08QvZMmxPgFOZUKNcjiSM/Uht5HAYgsk5cDsPnCLjeDo
9lo8dAGsK278F8eT9Rujy/uCesMxmkNt25pZ+aqmBi9a/b+tq1y/TxRCAIM+goupMb7srEoHoWJP
IW+osIdRqoSeqzYAyxOXtbbEpmXv4bWpDAsFSvuxEuJy7aMc95NX70Ci/X0xEvIXxGhNvziI9H+s
55teNaCAYoG4uhoHVILtpL4JH8wAdE2GnAwMNBtHVb1nmmYCxXKQJdoeXpye4BRTZv0zdM8gTbmq
lzLw1+RE5YkIh55xYEbzxQLbPA+Xz/VJ14cBP7oz6hUj9G2jf8JDLRIpoDkKPpFTUEnD3eT6/axk
qNEsvFRwnGTQcQcvPryZ32f2X7nYGkV52GMBPbi3vJFLyeUS9IQ8Wmc3gSKX52lyt9gL0x1hh1Gu
YWNIeOIRPkEJnZEdJ8BXD7WhxCjiYY9Lg3HsoEH/zXTPH4/PIIqS2CoGYJADJZC+aQqI/qZtTv3T
wWAR/UhYCJNnPruSnNVuBY4BtIBoyKoXFFiGQ6qxvhj476bqHMvnjNFzDR/zb5ZLQxX4e5sLbWnC
9ZvYk0fp+WW3QqXaGoMeW8mWLIjGbCNnRAfFrg48M4UoPWOXqP8TruO2pT5gqSr8hkRsPl8AJDJJ
Z7x2oN4EzPixMAvazQwpAs62nNu+3AV1G2TxH1liqIgY2HrBp9yiBcVfVKUae/y0K10ydbfAeSSY
dr5TOgbEzCHla1DM5xlRKYL47/W5KoCzBHrSx1SWmQragch9tSLyznK9di0WO3u799qb1SD7MOE9
MVpnrPE17ywpVX3fle5fzA8FeD3KjI/lKJ7eMnauKfOqQauzlT7HzYPswP/0dTj6XyGMK5LnuDdb
a86sQwXloFvHTIJ29nfCjw28MMqamNJd+KxMIhcMmSARY0uGkmHfUkpj17rc764l/OSjM4aCthfP
ersJVH9z7ozi7+c3Rj/UMDBD9iQpr8IDlCp36BU515Tw+u+vY4+cv6D1E2bEBaegUbzWUlPmCh36
yos3II7Q8b0KTRCNl8kvR9pAdArDf6C6KfcKS+I/a0y79la33tz4EHMdjlMG9RA6Is6eLrUWhlbd
ps5P8N6iOZTIKi75GiOWrvhd6wsLtIVBBrjGd7y40Xnw0b2+YgSS+Ddz1iTtibmMoIZQguXsCqBZ
0wgc4No3IYWzFsJP1ySY1wDNiGmjEygf7PoT+XleuZaze5fzFzn2NWhX7QJm4zqBasoGmQ/Gu0x6
bTznZfaGvc5jGxfeSLJ/eamu/apjktl9353w0uj1cl8uhvl2Rer1xakihroc8PZ4rh+VR9KuZ7Q6
oGt3BplQx9hGev4KCMFXIl5gJJr+vnEBi6U7VHN85broqjq0DzUgy82VSGA81BSX/6eSiRu3V6ol
mJkZL05NDoqzvg83JP0BzqhmrzA1Pb+GsW2IHoFkD0gEzW2KaQz2HvpO+tMSGYG06BRf85Se8Ged
s1UqKpFEMAl8/nxKqfLLzD9fGyTxVmv66hVS0MvU7XcsD+a/p3lMo0G6g+KNVGvfMtb3AHVfhpu/
Rx0HiY/eD+l9qTBkj2bEM23x8eTfDZTTkkgZpdJnmOLqChC7JQOZlewOyp9AIi5jhHrsesf2cEl4
PhiuXgxzPegJiAbaFt/d+aMtnQW3ASTgxCLfdp4WnwJdmBCnbSEqXO1EAEysHpgflevK2Atqv/sV
npWwgkWXCKCG635vmc15RiKhJGa+uSXUu2gpMoF3XRSTb+FDOcnt2+Rbn/a3aTLxvas9ZapPlwhu
Kr0FtXmyLIcE7BIu+N5PJu6O/+fe2QIDIn8H2gYSsLvEFLuTIhdOsdGjYS9ryUcZTBgYktRw0+Dc
jRT06J3zw1Ew0yuHho4OzuyJZZAIe4fuGWQC6TZF57X6MX55fxVYOuYb2jkFJOrHV13jnlMv2SP7
BSAI9P1zH50J6f62rAWf8egf/FlesTm9B+KtUJN4HJmMXQMHzbP9miWzSJQXsfbwVDO7zFJ8h/On
vIxh8ZJU+dCO1qPbgaOz4fazDdxyd2IcoEZaEuYlNBmInBB8TMTwpv1SUSGJx3dr2wl3bW92o19C
0Jfz6s0O5qdSyT0BJpBwe+vvvPFx/J9WDNkmxgqt26nHb2dp2t0dAn0KT1RVEA0gilulnkeT/R66
WEJfRzmEAdJ1hEokaloInXa/zLl6OtCCL5ZMrhA/419/XpZNbL5Y1xVzJTl8zrfUBA9AjY03FySD
85l6SPqhIBDqao1NGvBlCp9XNIOm5n6fAATDLc4c2ChNsj5kOPy2xNxYdSRECNvwMXppgmzeP2e1
QVhhpsHZ0K8MoD7FyO35B74bQdkyHNjEu1zL+tnLht14LJZBShlOQOuvTGOlceKtNiWiT0v9A4zd
HjeNIv0LEFlNLBGEi7wSxXO1YiYIlpNqN0POMbU5Q4T/Z1aIteG8HwGKNZOvzClZVAuGWNmvFqJw
Q1tL8zWx44mK84kKahRqPZ4FYIGHAnXqUwM91qJoFMtL+QQzWPY0bRh583a8ioaWI0la2tER/RZS
4xycIZwq6holSnjd9HWuc8CFF+ChS+Z6jQKk2OfGJN+jZrv/Gr2uKx3zUe4mFipTVAxKIhAU79iQ
dIbDsByQdRlCU7OU5UzrkW2Ih7kViDI5TPtYgIkpGJFdFmJFBx112g87ymz+NDNUUILeOrKKvlXG
A7aWJ7Zg9G9jipmfJ4C2c3JmEl3NcdkfGLzTXS2LJzS41eu3dTyLvOMdA2CqN6zhLMuBfr7CczGQ
9YapxDOFyiwd4UBfEAewsiP7TmU48v72nlQnk+XS713VtyiVzqxjWPbx5+GcXPeXsB+oay5pUDU9
iqnsJBaieDLWHY7BSoTnsJl/hRZOVpgSl1r5N2kPjPGoSwq06fxOCvDCCz6QOVNxAPbAmcxyXBu7
C9T61x+TwzwFYg4HE5yIcN+6ASnbf7JCigMUBCQFn+ZL4iFkBMEmnhUXbsnoFAsVwYmHXKdpvQi2
rVEnyuWlGDFD02QfhZcgRWe9rV+jPfVAMomR1iKI+r2r3qe0xXLtu9tvwJiwKQs1ObfOPdniLDRZ
QkL+jhDBU2p5gsnhXTaTFAzmIQwGP3otoF/c2n50GQvkiqy00yVAuMtiHrQPkPJEgkazjOLWoFGI
+ZJEBRR5f6/X4cwTH50lGI3xku2ItjN8xU2eZOspUNStgFko75P/pRdxbX6zmlIihYbSz93nC4/s
cT/pBtYG1Vp78Y1wEpluqkVL3Vg0bKKxdXbGBHOCd6UzoDmbZkPvSCm4BqJGs0KZGL23PUA4JWzu
9m0JUbh2YV4McGrreRJnz30wNCEaD8aNOdhLCwh4s0B058lZ74ApufQEz/bY/HugobYZoEmy8BHt
rjXIdlDqdCMbjDu85vW6dOmpnizmwrl/i1Na8KmX/6QpWjEe71a16p3sLSg5d8LsIK7hI+xeJn8K
8PM3zfLDILJRXabujRW7xsQPcfsSQIlu3KArFHVBtMBHm3DDCT+RUuy1ilFdktxHSCH6PPkmd7ZL
vyVVu9dkNvvLnPCQXRmq+MrxZKn3g4L3dJdFuxD2WRP6SYlZllCQmHPEzPDVZkciK3yx13Qqbt7C
YpDpQN8HO4DzxH05nJVAslsSbQWOs5Mtk7vFZ8G3005UnGmy/TX5YaJ9/ogEi5lBW6U8L2D/5FpK
ai4MGem9NjcmtiG8CHePrHGhGotSKH4RfzbpxBpLdEwKwo6lsl4o1ETLwAwll7ny0HcVGwIbBDvZ
hPKUxRcJJEWzx4lPrsdJa5vrPnM7muVCF9zJ6BbF85OUU4tAs9FkoDGCSYVQAuteuCXl32ce/8Su
kHOEg0j8sF4NaUXtYCcXOciLfp/GAHLbjO+UBNPHpEArWfgKmlo2hbhOXKV4pWGsf6bOahW+/Gop
q7zFA6Kw3K2IvrBIO/TF4vDY3jDoVXb89W9SG6yKQcb9eTCEGofm7PjRt4vTN6jBR7h66IQAA5Nf
YdE03xx7PAf93pOYeLKEvTLX3m7it5e8xa4069I5Py9z4FohGmCKbYEyWMA1vaWy59zfOi8KgfGU
yEQDd35JS5DwJNnLJdXV0Pq4tFTXqvUYEMD6fCPowRyj4p45OyOwes6oTTFx/wfb/9iXhx9ZYule
CEqFFLtf4bN1n+2JfmaC1QNBlMdDIXvJSCEW0gVp5L/YER8fWIvGFqrZW536iciq9KNhKsdwTrU1
wc97rir6BgYqYiuNZ76UaV26LVfazxcBb1BsxjuRcHd1sKdHSW8ZnzBk1R2Tfc9wnilpfzB6icRW
stwqvzqwKhxdJXcna6LcK7hKl6REreQedMpz2UbXR3AyU51pyw7dpkc+U4F4vUVkOx0BYW2GyXoz
WK9vWKV3hbNTZ7aSg+FB9EFbRv9EkmnLP9rslcSTPr6KowWTELAylgEaTgd1HtNo1kPdQ3qxRfDC
LAQW/aHpdBzWjjthegrF9TPNucU8usRIBIxSy+CCSQRKdhIS4sq8jgbTqctZg2NXS6r2g9HkY/Of
rK6S/Ct8S0MHRguPcXRh+3GI/Mbkh1xHO95xLrhR/PkRwrV4P2kB0mx7NGYGjGWbqMJZhdcsviqt
dTBieNedlefEL17/Uh3EXmEPvLxKV4OYu/9nkec9vZwRqd0S0DwLoEaAnZ8fkMCc2VBoWZ8SdpXI
vlq+YTXdexJgjGIZA1y/xfM+8jqxastoX3EO0ZsWm7HhyqdhVr4symBh07Dgcj4b0Mww+ckOCJnC
RYwjz0X+dq7SX9KgReN4XG7NXiW/NR1RqGnoskCvuGu63fcl/nLVuBYzY0Y6YuNkok+aK8h6hulu
bIGDXXwVK4GIciiIlSIbH0+gnpzRBL9fXeC961pSm6AwQ/fYbkQSjjrlAO6KPxKpR8Y4LAXAvnFf
5Lno09C9EI70GWOqFQ5WmAsWV8WpbfLdVjuCDFybqMmY5XboPBYquiDL3+gfCSmYAI40lI50HwzL
E1ZSFLbAgAFZ4PiTdKKs+axxYTe4hUNzr0m4J65N44xKFt2ko3q3dmc4e5a8nWU6/hfbsWsDcE3y
wXkZpA2Wwz5I3GM9HWiVlaT86D+jmruY8oH+Vc1zZVb9zwgkVpF5IJNNs0CNu41T6YyEhXnxTuFs
tLGkHFw2RGuSB2GfD4QF/4cAtS6jxjKcZPrQd+qtmu3D3D/TaN7ZiZhxM/pQTlldYjHQGtH1jusO
Oy79xWu5rto+1CvBY+jWQaeuhUBidcsd2G3SiXfMs4CowG7jW9qyqHHPEzHdubdieMLP8e6qI+VI
0CGdiiCVMDjjxd34+BUIFND23wBbGD64Ji9L/n89iU3j7jXpQf/pien4K1HJloG3Vtu9IjsTtx6K
dCW1EYo2xxdMa/1gqLqaE5vEndomJTqbXwZrcoioNMkE0zuAoO5+cAHFY31nXRWdkuBddNode+5i
utZb/nLCfjo5j3j/+pgVfK3cphzJXEiRWGMgN+AHWnMAGeEHYus1x0Q3oIiAOYus3khC4sR5Uxgo
M/DMOXNgthHPuf6b3JWgvyLGhhrrkqkZd1B1wMjqb1DLQbneWr/7+RMn+Q+3CFX2hOjlGyJHk4qy
80HW+840KqhvFPOJGr20t3AJylHo7arWMbVAipyCdUY7ksGUxVp7TgtSCo9OYPGeWVvk81UGZh3v
g9xX2viBFmZ2oH810zMU/UbjV9HkJm6A/SVyt/6TtPZHWaXZjz2NjLQxdtzoSMvM4oNhikML07/P
VdUduxeDewQaCdlKqe4tid8g2fmtJmtI3GW+SNqnN8a5Yc+Gd0sHb4bX7qJpSdHbvbFxLgygV8LT
KHmQ3elJ/Wtum35tzWw/hq54UfdRCi12P5w3Sc9os16eP4MjgkGZ75io6mlV5FevCEqYNqAeaMoK
AQR5I87LqRfjpc18i2jVf2/ZZXS0DecRusP4bN2Fgiz1TgiDmlviS3qECw2IXQqibgau0qh0bEsi
jqjl+2O8ud2XdQDcW53ieuq81sTAat7TnOhFVD9ncsjiXsiPoo1MQ8VL0da+O/OPFjPiIAparyqY
l3rExZnAIS8dwsIPVfaZNY3j8GlZQ49y8sTL4O7yqdNgdNS6Gl3uMZ49px2BkUQrGDmWXu1zP+EJ
UzkCAmi2PbY7lJ9xBnDMAgqRzhGuy4+RbkDUE332r7nI+AUUWiCdqyRXf249LdnNpp2A6PHpiK7U
NN3AiQ40tPg+tU505SNftSAdMShcDkYXdtxHcDXDKaLvrJs6a1ANMCcCtNZmMh6D4Ha6kwpUf0Jq
R6o93dfgZnBdEIvX8xOJT3SIsbNBwPP1oXtfs8GCRKcC/57B4+ZQQObFILokVL5KhofHK4iFKUZq
9l65Cu7D/s9rDotGQrJb2XX8HnO9JFbjdg28JYZ+FsfDCwpuImlSxiExKYrLmhJImWcXUhiVzxL/
UcLpbJk7wQde/5bpkufJuZmjFadD7DEHgtSrY+ATuOAwxWWkX+UOlieU8pxI47sirZpDi6O7lH8R
pU6m3iC1hqVodak2fK5qfew777DUr6npLHIKEH8K5NfObr8nDUndEhRXFph4jNsz3lIuIW+xo8bZ
PG2aYUQtCNleVmq/sjq4L/aZryT2tBnnzb2w1NCTPKST9gcjp+sFqhNOkuPrFSKWycXtSZ4S5wgp
1i3kv60KtX8l+axlEWp58hsa+4WTqc1ynH8kwju7CcaQCvc65ddn/llTBLSRiVluPBacrqt/KEXb
7zLEJcWC7qZPWeIH0Kkdp+WAcxUX/+0aBXjk+UIIwmJdgjvc3+GHhreShOZkKHQ/jEdVJpRRUYId
UslXeoZS5t1D5h9NGlWu9RguIk4PxO+wtEedS210tZhjNuuzUG0MklzBRKAo0/MsLihMuR1gZf1r
zrr7oc8nI/r98nltfBJ+YcxW0y7Rem+dmfoUVZMOdzC96u6ka7L5mbWdBsaFqJui0wBrFQjJ9iA4
DZPNEbkFuWHZ0HY/+R7ZhSLg2eLqtSUYqUAB6mbPyhChNqpy1G35NjPP9xzTjqPrSC8rA2s58zSl
jrIgOjcBWlr1wfw1pUFlnC9zv5JUFBziUHLU+hrSfH504uLonQT/482YIRlmaJ6InPeHYGTuIl//
fTIIcIV16ifnDSZM3goDf+105ZYHYE5wt/+h0bscFrdniMM90+rX3Iz8uJrYSRqA5gKIWZ9thfdL
zYLFPd+Y2Dtm23GEa4LquOZp0x7/aYg3+Lzy4ziH8biPpHP3wu6IZALVk066aVvJ+Iz8TVhjLlSs
KaHOeftTGnCtYbHPtV1lLgba5n+95YSW519KlsSkBMMO+l850f8u2zjRM9V6H1LDoLEcyHm98KLy
JMzAfzrjwW6Cio9e6Nb2GruI9l0uP/qusAIt0op86BF+CccSei3zfW0krgJsCGqJH1umfrR1/3Zg
hgsp0NRRK6nhUu1g/PLompMSawAOP51Tr9C9GkB5ZvZAXec0H74+uV4R6GFqBYEU7+26KJgUezn5
L7bkODJ/jdRUVfmghceHC8xRI6gVrlCf5weLm0KYWrGgri26ALPiiQzXHl5uu7ejoyA497XZb3Hg
TXDJJAnsXPmNgQpQSo5cnohI+gREuhqrr3ld1i1DbEgx76ItpmxOCKCB7HKI/cvi4Eph6Fvm8QPe
QFHZ4XmhWSzwxRKekw5zWhdOzea4AVIK5toVZOyPBYyl81sQMCdC4cKs3ASitEUi+U8SzHX/Diy0
oyu7RXxRwnNAARUk0egpRPlzkulHfAnFUKN0VYvm8/pzEaNo4CVtONDoGfFrrciofqgIWY4A1OG0
cgFcdJAOkoDf6kkaBS3+XORomqqD8tM380VUDPvIY8EF/xfSCr03mvU+7xmTSylrUO8rZ3egYldP
WN4daaaflZ9iDiQNESGwQGEeow9OoWXbxd3iBvoHphJwCVgorHaI4xMSZ8uG6IFk8PG/LGW44PRK
3jq2h2s7TAq1v91cceo+h3KK++3OFb8N+Vw9ILX3cVg0QvoDuJEOadUtTfwgBeIE7JoYkvcvTiA4
X3JRPdbdZF0Wh0OIM8HXk9jo1tS9yqwoINsq6sb/elIx7WrEwMzGaGyShzn9nDqDvFen78gYEok4
LPqux3yTtP9GtF1+BnJWzJ5a4j49Szr/Ois6OqJ/XCz4XUMB6R4wjfHKO4ySpu2U2LRxslR8Hfwz
5t937IVrJ0VcsmE0Fge8TLSvnKUNNqK6GHUfkkMLROEnGMN4frbDUjvwEi5TG4oTCTBfLezk1m1b
JheETIMSxgK45KXlNtoWjvVgeBZDBYmZyzfpwZM56SowML7cGtGEzjfnW1kZ5GzBeZ7EfHg4LlVx
vzTBQIayb4ELEKR5KNaJ3NXWsPAoJJyJNeTc+e5NaLezg9Trx4jAUvjPEgjnAL/u48UfSQ7A0+mw
/X5KAReqNsBNXPmZR/RJs9x6fgotapooamcEfaUG79CBmHtlpXj/G/bwQqyY+sWyiHpI0iH6qf3x
Vp7mD2ynAGk+c1GGULx/bKbBKuXZwa6FUZ8QCQwHKblDL1tX+av9OK//JxzME5Kt75c1nUVDazmT
Ooj280cORCVDq+x1CZfceGmV7W0dP5RYMOb7/TIRVt9EQ1L8vSY6ouYP+NrMw91vuseRzHhKPtDs
gFBl2CMl67q+bOU9/pTL8JymNtJak9diG3XCQsehli4OO7OfUnRz4QBKyHSoVqgqiqPknD95YVXu
F7/jEsHfG+eOMINhpIKW8+nBUilQnE5VSxTBXoMFvLvyvoChrMLQBPQj/4WXSKto6bBmoEnWeejO
XEhFBnzh6Ndm4HTLytCQranvac376xd0rMGT7A3WZkUgYoup1HSnsDx/0M8iTKnBBhV7eH+Yuf7T
RUsEms8z12U59y6j1IesrUJ+7oN8ctK3PMOnEgCy2euBoyh+/QG9zlcwLNoBktXdJ7OijXCkeP58
kTTlftpIiBBbuQ0bWazMy8jVSTxIa7ovoUpas9tcCYHILz2oCZiHRsIlNM7sPhrXKQoDW6UBSR1P
62ctP2R9OmXEJ5md63ZgYUmanRITSWzAg3MZsV8y4+0BL1vg0KZADGh+QMOXmBch5rcE673j32yN
1tNoTcCxf14UDpjkbO+blBPPrqF3/DGzTzgOqF/hmPxVVOr1htcpo63MqLTuRdVxbUidOtvZnFR3
b0lB4V2XSi4Wn/hV+jvnVbR/Yhny8+AZ/HZf1TR8PrgZFyhKwu9nVlUpp5+3nfdBLUinTFTxpQro
VY5fgewl9Kx5z7z65sU4lW3VjcIIc1oOCAgYGJZ73yzmmaer90hS+a3e+0k1s8CLV8ZZ/Eo72vxa
wNZ1yP3wZVWkOLBIgxw+HRzADmao6sRHbnJjRvMqKg+ayJJDLLrPZTvVa6DY1zkkAUI0N9zhGB3E
bsQHuVZDM5De5eQyk8Bhc+5r/vJisPaU9tZ6dtdzXa1zMGhDugQI/5wnOk0gJJq9WVCrTeFyb/mx
SFlYCJ0uV509wHnlXYdfqII0Yuo/+0YSJ/CiQXX/PvACMoloh9LU6mxs70xvXCJV5xcGzhOdc8nj
G3SLZk+KTKRusR3vyJNrUvf43ReA14eylmMLWfS3lN3zto6JVnohm6XoK90GfcAn21UXayd5C1sx
ZmgOzkU+Lt2yE5LrJ1ZVWE7kTdCYvoAupujI+akKX4NR+cKXC4v68fdjcyE9+cpaAGo/Iho7Q8II
bY2O8vOsKfJXMtWyDFGbfxsUoO1FeghGI028MpsPM5rR/m+cNhGV5JMGuRpRJ4nzxUnFEwAyf6MC
7bL9MYdcYBifZQDv+jKCOFtUphqDVwgv/+0SegGVukFm+adZ4/Bfh9qZ4l8Nte7DsI785H46N9M6
U67d+n/FS3nC3UyrFs2reHqx23hmASa1ae1NFMXz5JuCjsuNE4RS8i6MVurwpjvy+3XLh8fMslp8
Afp8B3K2+oh6SNX+GEvVJmzAZfUSUUxz61bj2ks3TyIFuW6RpY+qDWIc7uOCIB+bk1W5CLyaXUda
axiQ6vT0FjVavbblLM2F4zdGozJuYbyPJJMIM0nyLxkqYSppavQEmkvGkxrzxJ5uejO5lhb3tw+2
PBbMOR3ubtYIha2XI3DsGsomBTuZcYvKQWpTXHHhjSopBgx4VYoH5pxP/aiyeRuQ6kXjeyH5lR0w
3Q9Sue4PJokoffyuegN6e33+uhEqDR0wB2Tq2SEWPO+Mquhh4ecSIC1DLec1JysSqqN3TRBuTvH9
z7n+oSD4ZSXQhZ1sMGPPVV3cVsjDau9eJ3vUBbQnNy/uJcus5KdSmlJVQRwdi9A/vskPjeXkaGEW
M8Cv8aD1NnaFQyi+8nyt48tSXBcBAC8ZSuRK8evGU4rRGbs5HQZmaL19CWV7G/bP1sKzx0PdSmiF
JFjoWH/gGalMzlTP9+aM2cUYjSjb3XGScMJH8fCS6P4n2FmMj51gaXtJWl3zuoQqr1GgozfmTmMx
pKNLcwrpgFvs1HnP2ex4hJ9BqasbqL6uYZopdAFNdq22vJajGs1n06bHu0fyDPyc1F7/RIkz3ffs
+e9Hdw+t3M205d3T4Bgvmbm9WyyWEoWibvyz3mcXADMFgieVg9WP7XvFxmUM/l/e6o6YR0gvHjgE
h/PHLTaTSvJZVgG3Wwm+HCVUzu90xea5R90288HVAlr9WIPYKVQEOapSr5zQKGtYVWUM+JORNf8a
V/NoP8rtIWK/ir/kkzpt1dDTV9suqnzMk0I85MsYVnTLrFuqrCG8b/2VyQ99w+tSy/177vyBqWkT
x3cGeFd8i8luPyR1TS/eDD6nNDXiZpUUf72Au+500Dw3bxNmScAgtTAymc7QLJ3Uuvl9NLr1jqBH
X8SdW6V1sGXA2zYgAWXBdM578HoBLVZGvqnx91yHyEQyvf26AoBwCls3sDn+6VY4O7pLeWFmR8c2
AMcPMKK2IC1rWOrTqoNpsqNuqel8KwC//LScLp41ymOY6VE3VsSNzXGgYGEiLj3P+YJrdoNPxwI9
hi/YX4k7+acsQFzMRr7yIQib9S0CsK7mkpPjgbYwKrhu540+ikh9TCs+QJNbwuQ5ieNNQEq4CTyz
pqj4WSsJTTKUAVyddN0CjRcn/9L2OTI5CxibKvs5YHVOYUYSlZP3UykzS1pA5Owr3/gB1Y2mlcqi
MAc0C55Er2mYhbJdy7irffZX/kZCGL+Eh3M2/en8sP37Rlm0Xu/3bbEyqmreSy6XtHcxQBCgjs5A
kiQIZ1GzAWl6/nwnr9nFW8hPcL8dIhw0tt+khHAOyuxUtRJNcpwGzRb5MB+IfwQNnmjoB4+dVAvZ
BHsWOqKsZD6ocgqBogtCVVXwOIIhhSIXSHd967MNjgNzPznqYQkuVF7KVPADN75+T1a+PTzrFo9v
KI5udreIbWLQOTaqopY8apfpb9O6fAIOqmgk+FxcQbPDfZQx3PtJZCHhkqez4AIGwnzR2m/uC/+y
CFhAHPHtoJm3xPhop0v7USofw04KrSNww/txeGTUen5FguvDAfbrv7CWld3bd4VRDTJfX7WanCgg
hqiCazE+PSjK8RF6cUzIE5k4tZc64EO/zbZrzPurt0Hb1OZVB/02buCZmyH92ncv7T+raB07P1f9
wwKu+qsmXYPytorScT6+NeDCeUokgQ82i4UsaNbF9b7aqUtJhoVbCD6luCnOUQAU50KOuEIV9cOq
DSHDqgP1O8+JyXtqdb//+Y2B/HxBVLnfzq9HFzqg5WNM4oCiyGYXdVb8KOnnv+HRZWQu+mnSCUZD
i7zf56l4Tz5p1dVtEkOJ/+BDkY4lXh4xE6rhSWsXmJqkDhCxHrjhLVcr+2uQw1h2Wuablo+7VaWN
bnkpPsudbRVfaZ0j/Yo5/If+sJDIYYHoZOjmcvhDtrB2K/HOFwwL7tANbmzX/xpSrNZUfjo8Q9cw
7Z6oxNg8/6c4hO1srzJ/3lDVA8A3pv0JiAZEGjKfOglyYpVJEvb/nL3+OH9eFhfAIYZoZ6KuLmjQ
8gyiFBd+Y6akNZVjdY+Rz4wx3Dzq4XnrWL6uL2JrTjni7oETgLHqDGTLGOTURkwuVfGIO5KusFRD
7v1001VUur1PXqDGZ7TMBsvbrv0slMpAeTAsW5EX37WzXyKqLeeCHWGysODhk5m2+ZA1phu+oMDj
0sMSi63i7unsg54E2JQJTT7w5MEkbhjzvP6DjUxkN9d1ZOQb3gYRGLmxc0e+Yxw5xa+lIKYbwtAm
SclgDEW3yb7vCDO8G0dXj5xBAmTN8X66AwXZUboGP2dy1/rirXbBnJxVDEYoGdKLW0LvYAdevV3l
j9lzoWO9X0qbW5Rg1ApihzJNELJMfzB4R5hq9XsHCrndfU8ZtUBdWWpBOrgVWRlncATuCdi4eYEH
1HUu8PUa76oDx9AdWwSQI74vh99DIAX29XK1+vsKgWAxZQyKQ0QfIMdZHNPPktk3OJKpmapyI8CJ
r7BHpzn+padGLgmqV7rD3VA+kZIeuOviIV3DLxuuIN4yWiN70EPJlznc1TfJNjYe+WmG4eJvcxm1
7NfZs4lLYMpomhnBeW/ZB7H/Pva8shfoZaqgTULwknUvMy2huXedCcP8NG3nILyAchqVqlE9zVqz
ZZySEhnifGOh5+KP6jMinDma3lM/l1WvPnRtOVL2dPMqGrfLA+v+1cllVaUUmhP2hs3PNHG0RPFg
aITNH+lFQFN71e1VluxDKNolBFM7RdJMRtVrGTzCkpavJZBEc5PJ2pbgF4l6S+rhB/OjPfWLjzcl
VGPcDyzkIrFM5braBs3HN+7FChOqlEM7B1pUQrUI2WpkJ6YkE1DkJYhwH8/xnbgVyg6hX+JGltRo
7p6krgwTTd6hJgt4t7WtqkAkMdE47TMZtwdY/B0dXl+tRYClMojTPxfu9t7JZxjdYBMmcpli9cTc
LOpUSPGqk2pJjLp/CNRReHdfg0XZbvDTKE0aMiPCAAMogYbOVFF+o3U7ShAbnuv5F2lwM3UM/Km0
VjIgI4cn5YnQtHRePUtfkT+Ize4lFB7Nx/9W4NfOZQMq+7M3vSPUCeMdI5tuUXC1zf5/xAwlwFzj
QKmfWNhnl3SaSMNAPJ2GMiIWM0LSJftcVl6O3xXrb/may3+k98DobQ+V/JC+tHkJAW9IjypfNXvU
zZLlT3NNiLGvPccP2YK4iOpe0wnHGAZ2P6KBBPC/Ui2BTxVq0ZhOT+JNvXbpPRNpElIq2DKEafOG
gTDJW4vXzD5veQUqefVk8IvID5krgSzHggRSsSOXlGNrKKXmuW0wclwMWnFBdkNt+fMUoQX9K3CX
IpZ2zocec9FUFeYScvaKixp7GdUnJGlbKY0z1C1wXSvVK+xNft2Mx4g583pI1q1oKUKI60wb5+Zk
4LTMwOPwNnAUoBRWoOqig8lbM3EfkWI9xhwagpLBZjGJaGNezBV191Zisfq09DA4HoR9R/NPWJup
y2W+5EmUfPUEsEzaZ3el727wxkH4LlKPaW1BhS9z/GjY5yCpeU6/cWgOks5R3Upt2y8c/x4brr70
2CDmX6I4D3EBX5PdCgq9cbqJoFhDUOMaV42ZLdyCbEF1hgKuSIBNA+XeVpWi6Jq7TiynBqVUcoYw
I95ECT7TKjyd0861QZxyKvck/f8MXtrzwqgvqCIrVYKBuQfL+adw9kJ+n3Z5sPDHEjK56nebVAZS
uMwxnFoQnEHhcBeJvOghd+ENE1YTQkE1706N4UclObnvlJ4mv0kCGHHfC5S3m7h/FfH3ASEwJgUl
bB1wIgmS+zhHk4VNbB3+nOnn4GWV/v68jhTsUhEtIvKWUw3xI0B4HZYFGYdjCW2TGiZH1mQHrb9d
SQVHAKCqD8obCGBOHjgh3j4B7M/0tMeJnWkGDfzk2j7MOZ7v+RY8JLYQ0RqItC3uFALG2xNqHTBV
l1x18CO8dUKNCKVIGH2nH99QevYVekuE7loRii9pMoUv+EEc3s613Edrek5guT4IC13+qjwXaIEC
TLN+X4YiGWHl+NVsjQrP4EL86I7Fs/dmKV6HyiCJp5kavVYQA1vYfNuZcRCwn2y1lE6KKYUiSw5Y
gVKKz+62Hm/DoBTadhYW0mJpMDaBlE76MdMdh1CdfMcVpxoTQVsfohUm8ryBx6G2yt3BCd68RvRl
g1VtaTUu2skHAaKigialtHhBfpvbjJse7lyqg3TTWGBXXVUdarpacaDhd3iTB2ihGof6P84LaP/L
GEVq7gShxLj8ZxCcp3fLBZqTX7LdZbouWoE8gYikm01mQldSQKR7OvSEmxQsOZAO9lEj7UwpbHTy
6Vy0xckRAQ/HZQvjmlXvmxl85fhrZz33/0oKtGsoEb+BTCZn7B3UnUnJuhwGr/15ZVqW/xtaMl9U
5t1qUo04yVGqUTuU+JJzUEWuRKzmiaMWoW3f0V01qwd51K+HMjiHY1dNHZU9SBuNiufGawkZSHwP
iUxOjNoz8vjcFlaDrO9dSzQ/jkQd2A1O/Ea1Vo1KrkhSwdsF+A6DOD6NPzqdoTx0tj7CTC69Qvi7
ce0ldevtpxdR3Ds/MqQBMDJhNO5X+lMGfOVd08mlj8Ht7ssphwJ1Sv0zuUXgeic3jAi3HFhkljaU
QsFXAH8ye8eIPE36x37aiAZ5zlQgu6iDI0EQDlhdL/XrG68YULLc4mFrP187fTPyJMymvJvMJZMM
vFDuGFstOWUyQ8YyK5iVOcohjNIa1JMLDDlYNCEzxmDuATQP0nYusWCgnL3k/EPkYqvwUMLaXgl5
rxAklrDq2CAr1/BV/Yq7LLg4CQnRor7oBgFa2BTD/Cgk9rUWHZU38MmwuQfvpdz/RdrEH0FjeycY
O1Zjoa47NaS42AFxNhMQU9SK4718Exz8RqVDprlBuelxQwWUOs9SCcit35xBlMHw+zTSsNQMM9+W
G8zba8quj4iPdrdmrE03XUU058Y0nHYOoTp+kSe6NPKD4pOb/S5xQ/X/lydPNpPN+byShs0nnhXJ
79MDwX1dk3no1W1Dagv7tNJcBs3Kqcj9vsDQ/3G1UIeCDdy7IZW33MdKHOPtcx83wf2d6ZWM0nhu
gSHLqkBO8y3qdNdyScfXY0R1ffsJy98VJ45hkel9Yibs0xbf0SRhJ0LOxIRt3bvM0sCyDHKXMWzh
YV3wbfQU8Muflv/n6CVEqKM3zo9cpvQZgYByesePiUNmk79Mf2iurptg6ptz6xpPMsWaYLpaKzHp
I28tvDT0ywCfa0/mON856QNjuyJCmtgH/1utOj4rWRUfIOL9Dt9mqlgNWTudB9zdjv20p9PevCS9
J/RkvthCB/T1VY/QL/A231R8C9kUE1clS7z0Db9ibYCjDRPSfzEahxWdplEXSeIaiczQBpFgWH50
rIehz92GBdIqUAbvXFZf17hjAjjgOVrmoLcKdyr1lv8hO5KES9zn7xSgopJQE7mBb/x3ZfAxZE3p
UOl3enAo3m9LM4kU3jAPP2ucPZePAXg/hW/DKmTOCFz0SU9gc9xqU9pVOioPsR/5yZdE5YSTckvs
0i5IQJK/EuPp+2OBQ9dY6M1OnbOKFou+ClcaQXWRJjR3lB2R0G9gMfDtPvM2T0xBathy7q0KVwr1
b9162UiS0ue0BrLzRzfwa0r4eKq4usSejMcB37ipDHWkNR253HULRAbnd/ass7AjQ+65AMCwGw1+
Pfn7jBXf84of8SgMABMSX1+pfDAIIGLuq2l3VFJqcpFJN7zUGcYKND5pDR7eiU6raBAOBICULiZE
80iePLi0YbOa5n2P0sFD1T9u5aEhLg7eL+ODHN5xj6cv6O7xrXC7m63GaAjCqo90VkK8y9RJ3Ynf
ChxjxyOFsgoWYLExDCylmTq7u4a+7W9tin5cFpIvV14SlPNh/vNVIFIf+CF6ICHP1Tt7EZQ5TtnS
5WKM1sI8AE4rWAqCp8/QLVWFXD+59HcPGzgajM+njDRS/yZ+m+GwsI9J7jghloAuN/RAzfE+Gtzg
+EFKq3KUxg0DJyFY94WrA0C1EqDop3LvehGlSpjMDANoPkJbaieFrAAtwm7zT7Nxl+7bSag+plU+
ZV+Ly6T5XUOvkjVhUIEAi5bQKztWAu1s8KxWsP0LQxGYTAh0BIWWoBAEn6Icndw99u6i7e8W4fe5
XtgrjPR1Fs1tfYRJDnL8YZLtcKoJt0pfQAslQJNOnqBw6oh6CPvcouq1JVHddSGG6LSekzGbHrQQ
jirFWpDd4MvDqdzcalQ+dAvOo0vbmFEABH8vTk8q1aDpPN/enNcFIxflJgjYFpK4PwnEgUyWRepw
Tm2oN8mtd8Y9KlV9pik6zGsf9e4V7Mq7gWhbs4xGeeBXiSY5M0IymlGT4XhhC/WCtaj/qZthaQAD
KVPcRANA80wfWUzLFqX2rUTD2YXfl/xTXgoQI8Aj+GcQPcwaHO6pZOhYvPNF98s0RtocAsOUGJc9
Cse3Qwx9dSmp9McctpIu2FHy4Ib3ZP8GX4u4Fv6zeeEV4xf6TdIoMeMTUvIt+2nQaAISbPIH2y7U
C1lhlxlqqMjlFh6xMBlmgY0fGKw8Yv6Fyj2sD8Rj4FgRWaLYc3SgRJAhSVxmYBtLwbfr8P4lbrgL
TjA/ZCOdBC6Mb57jOaSkVXl8eJqVE6AmqoBGJK4SFmbZdC0Jj8HALr9jmZXADgHbqgjcW/v5NYaT
1nw7jA+VDOJVyK8qBySceqvm2ahuRwiIETdazXRp0BXUbr9gSNg+1S6oybVDsok9Gnh1bUtK22AD
7Mo+vnX/uz+ziA8s9ZcKiChuFDtbeadClVlDjAUx58HKYBlaEFKmYripxC27fP93au8ptzGW1njK
dL56jgKhuTdrjniInVZMlsP0jTV8NCjHoTIGqwNC/vL7zNXlW6BHRda1yXhvq7UT8qPt2wgSNu0r
oipib8bLZAaA9U/9Ro1QDxVkR00GHwL9vaXGJkyK4OumQq41jWoL+nmllXwVePLMZpDc63gnnsyp
frIi6wWRb3CpjYUlWwCLCRdwnpJUh3srKEK1koij8FQ84OBz5K4sbppHe+Z7ABzpR9xhvgdMxiug
/kJ4D7uJSuiarBcHo5hWiynLGfYJ6WpYSC/q/1w0AtSPaueyg8ElyFDSKDjKd0/0zHU7Atfa7WvK
K6RcdWD/yLZiTtzjn6x0Y1r9zaOOj0b2MTzeDKneWtkLbWYy76Se8VQEdArIk52O+SPMxGd/xz9G
HbZ5vcZF25dznY8uyy9yh7OGGnkg4XZiSyim+2z4bTzyOwP4nNzkoT+oRRAmreDFuT91ZrJufpRT
5GsVWqUS5gwtYGnfGUSJGeMs4p/hrJZVH64voh0uQ0kbG5iD1smtLA50qfva0afGBKFJhmCAyDur
GheQDTsXdzjgn3MWfcWxKHBY2EukSL/67dxI59kLC41j710zR9VRDqGgjyQT5cKXyN9YLIa5Omdt
qYp52KD3J2IM+Csj1mLG2uqXTyrkHGpswnEfNUOyZAK8FIkshklvkjHWkqSA9QhCuEPLX6lVh118
L14A0k/PcFQGtksxiv1wzfeEs4NqePdlvs0t3Xs1EbM7MKAC3YON8MqNQIJDS2IIxg7rJdeKlP1h
QyYI3r/wtqmuIX/ZmjHoA90NDZoWAAq1JRUBodPuiFHxzH51CXNU/yXHeM9PaX11rDGmItLQIelj
9fL9hpbnDkxTz6guyjaEP39jZI22vzOduMnq4UkSl8Lx8mEDoxiRICjZGjDsde7LuLXTOep3VNtl
c7Oo1raFN6+fgCaqsqpUielk1tDABpJr2lw9SQyRsCVX+CmJq3KZ4bg32HsresGiofgWxoDiKBLK
oh4s0uSgIxWBm4P20FxyQb6vHjNb6eerDAnEBTr4bdKoe/490OrkdZT5VdMJFvju5E6SXgpWBfCI
vPkAbyTThA0D+p2EZ22Ll7STGTYnz0O+3LV7VTKpvrNbh/K2hkPptz+v2xyFzjis446BsA+TxmwS
swi0QxAwONPTdj5pPLlbD4c49gUk8g/iE99YAHW21SLhbEo7jkCt7Mv/9nWayWLpRW7rB9hBE9nj
gA8HawQyWKwp6qII12QvoJWb8sMBYJmnp8PVPzUyX8Hvp2VtnwEhoNNwLEBnzwCRG/3LslmWO538
nCQGzyK6UgRJ76KaqfoM3k0DHdhN/ElMH1NIHN7ti0U0k+FoeBz28Le5yXztsv7k3X2d6+/unad1
9JhPltAItDckeUvdlG0Angyf4vsyNVf7OiPiArHGL/k228aT1JwxNzt0shUXUOYYeCbcYR6BZeEW
aDWQdxUvdpBCLz3eMeYVCCoGxE1WXNsYYM3Z4cGl2qTtKJgc21gp1R0GlXEJxjAe1AGDUBhnMw1z
KsAIn7ej4b1LGvfuvXRkipvICV6M0UyK+HsEFFH3Pdq+Bsd2d5mMeDI/j5dt+iCqXmfbdq+5VZNL
FhE1crFZT4biq3n3lu+8lQzalR85uQTSuzSBpKJzPkBZAnLzc+R5R4LRdtZSn/oUopplW4lOu6Jd
8L8CyATVSMSNITm3E6BXMEUIbE8T2H8iRWivCNv0zXkIoAOLLFvPrhn+TI2AgKMtgwDz7pXJ8n37
DivZFjhfegwG68vx0g7rdQXy1X7zwVYzMMGrQ3RPS8g2ikINYIUV42hURroZt7TXmwyPHYMeyTcf
rPorgzU7RrWddA9TVBrrdGX3tBDFssD/5HxfutKQPxT1i4Ia43Jlnnu5gMSKkFgrz6TKXOSvRtwm
enXXhxJTXB14IWK/ls6sBmwFBkKTvNQYRe34BqCJ0I0rxgoGBlxbWCEW1nVQNVlwLFvnzH8ebFYj
aNMGS4eSRuBTbe5Hn/ICyPvCdVveNvkHFV8Ra+PYBD+K+3ilHlD51+X+hn70h1tzGPjb+f3aLSO5
scDaDJ+7FC8OamCPzahOfGUFoHgbUXPDRwJT/hBzMYyVCGF8RdObShR92ODAs41HHRYhGAOTur/H
tnnoWqMeJu7/SbsyVUkJX8Z3LvBduVbTAUzEGBUUAJvfdMGW4Z4Mnrxh6jnurdoBIYao2JodCOh9
qymqxPhpUT/ewk+xYbywaDS1vBEnyz0W2AIT5EL6ljB2xfrd0XnYhfDvaZbhliBvl14HFlVYMlZr
UXBIqKuxSrmkEkDpLVHDYgLxqFurBrm7ItHehLdhGH9ae+CV5P91aCJehvLTpOa28+FBrqPjajnV
4Se0AbDMcrIKetjUbt/XT8oErTla2+gpW3Ix2d87jsCnmsONs6SkqooQczlsIZyHXrQXTZZG+Iir
VSSh1VqgIgQoPT7S7JntegikyCbHk33Q8egW/4EIfO7j66g8oXW7XrvBSplV4KcMKalVUM9skMTP
Fm2VQpBW321YDSg8mGqd0MJL/HUSCXPj+ZQs1z1u4eOS9+F+jVrKSXlzkRv8IkzZuRVzp2LhKCon
O6muPN5NOVy9tvOy4hNLHdpYYNwkm01dbTJayPQ3/QM6VOX+ZU7wsUSi+FoBDn8bRJhtoVwpxI+p
YIzFTa4NsABiM0zda8LDepQT6fKQZlgYTg4C3YzYLdirQq2bMDWMKwzZxCm2jsBfnnsbp1pZoVfh
tMK0ZAOx5gn6RQGR8au2gtKLlHDNaOy0bBL0xpUeMWsaH/AZgtp7GTtsWdSBhjW8H52AU+zjQsLu
bWLILVTHEjyqvVF76bAKstOwvpipghUaAqUMS9HJXKZqm7PjimqX37aqU8ggK+Lv0MUGqMejJuX+
0SzSGC+8ep/NnBOJpXydT7uWe6tQz7sdHr6WOm+UvWehLg+vHASZ3bQp9Vp4aC2wAYG6i340qtdt
c7DF04pX9YI2uL1MvrsfCKd73p5aDRADsZo4Rc4PBb3QJSfq6ZqvAytmkxAQ3NSWF4D2mzIUM5GF
evWE3vEWPw8uHsJ513XVykKwMj++5i20hnVVJl9xwNDzySknFqaTJv7hqqj3/Aqr1eRJ77tLOdTA
0X4ov8E+WHfz0Rz5GVlmU0xY7yJr2qf/UIIJaLfGH83kmurWiSd8Oe5Ty7V2zApwViLtoP6tRWkh
3gYiuBOiolv+OAu9mTrtBeBF9BI3BWHn5wwiLVeMLGtS/vBY6yDt7vJ1GTO37irG4zcGBPx3m5Fo
ul6mxGaqtjXunN05JOaHbVXfgV5apMrd1meLBDL+0nFA0+zXgVyLs4M/f5jxZ5Mxz+VdJZddb/wx
boEQHbLvT3XhLL0Ozn6uFVkOSi2WzX95yPIT5bNv4HI6luTZK4NtaD/5fHDZ6RBdBMSUUP8EFGzL
hD5qSfvh+IAgIZuGWs0EG5HCRFbOYBLsifpaD3RvEQPUNhlgiTrWlCGCymET0rezgUDHjabRxhR2
o/ySyc5c/EnaFVKUKRWerIf/KEul3lR6Q0H4WCxaHFZZ0nQs4tFoiWAmxHnnrBxC6AdBFtLMuYU9
YNc1KkpI4fjuNemqfKGLkTo67NNnHXTN1XBtJz6Y87P7JDMcxpx7RQOhMUWH8kRbHycPyp+je/Oq
XKbX4cF6EzzdDeClPev4oaS86SyaGYTcJZ1FERwrV8tQsJNGiWV6RCAOl/lfNPmanCHUYn4rZIhn
WwuXGDPrG6fh9uqKNtD4EdTNS9nAsHNiTXnMsyDNU3SVZwyZvKy8h0cp7Vabb/ZvW8GpTQIu9wfR
tVQUj6Q2Nw2KTQLrWAZd9P8oqd4SMEQTaRwIpM0YkRXbOqG/Sc73W0ZIhNNyu3NMtVruKmoSIBhu
KjEfIF34RNdQBa74w5scytZKTyAWwwZTUCo4/+3cJxwucpBZzfGOBsYRqUUkwWAn6e0ajkjqh1xh
ixoUkz2CFFsGIb8KObW+0kFytQsn0Z6ANL8DWyLAkNjli6BYl48n8YHnvMDNHO8SecN5sTZv5FZC
jv9PXEbmkK12Qj6fdaXmCbavMLIgeAq5k4/p5KEYy0XIvQwWVFiAaEupnsXaH+Gj6LkUW8nh4KnO
A5T1H/uvh0QjSSKAyIEZ8C8A3gCgIU/Zps7z8Yee/kI17ULsqcl+P1r306Jn/lcZx9F9VzgM9mc/
9wm1SVgkNMuNsZmfyFVkMi9GoNCGSp8g4nj377SAtmjtNpKDW2/OrCphCJlmsaf+R0Pd/f1Sifr7
p2/EUe4YD1ZY/XYQIpy6nuXqytX5R+4tg82aAtzMYQkyBfiTmnW7WUMvg/e15h0j3aq/sG9RQovi
IRcF9s3hNGAn5Zxp+gkecvHsp1jAfpvtvVc8InY0enj9J2NuZSgSLyiQljG079SGnQZPy7Xl5Smc
PUyz7MHaQI9MIY0rN94qcPWGfmgZV4trmu7fBwm79FC7hhZXcoEOzCPT6DAi5oTi12T9lh9mhVhU
+ND1VS6RAQD6xjnxBJsECgJup0W8LBthi4n7glGcZ6wrx/Mr/wLmzIAjoIhwcTNas21VQLVuhOjt
6XZvjxW+4lBMCF3TXyJp7axL7vgIQz/EJ8JQBF3ZSlqLy4rz5dr8AjFqH06IUlbi4adlrQW82+iV
3HpeFe8XJwdF8jwy/qUMnV5EBmmDe4z7v9DNwapaYLnO9v85LKLtGM+xW3r5M/rYSmNd+DVDfboU
fDa678euxeTenOeeTF81o5sd/8AePkS5MKSgz0SdzYL1M/aA9+ZaJJOOyYwBd1HlXnkFTkxI5hvS
5k7HeuxXjFkmqHBMWSLxlZZD3NFbNlnmauhL34Y3nUJlhwmRidDzcP9nChsf9tWGzDMtO3BtxfHc
IE9j/Qk3dVlpjuYBuw9UBDuxNEd3MEDG0YGynHRZNlUDmpE+ig9G6JWCZixhEP2qzGZ1eX3OUh4F
1LD7Cyf8ii+nT0cBqKiC3P/hdeJi9E8MNsZlm5ZadF7Wso864/oV58usdBI6bApu2hyo3ZnpvVXw
h8AIZfZGYeoAc0eMEc2jp+ZIwBNH8hYeCOVQZiAVxH5n36KMv9BpEx9fXuxA9Z0LRKhmB6siiApL
FO82wsfVEl2rqEnkozGJra13zRWeMuS4YUrdbKD1vdHmTXVslkY+PYmpw3MjO2ZqMKUc2S9jQ+G8
1GcXEMTB+cTrx7Ep58Mx1DiIMA5hDZLAl7qaf7FjqdTACJrs3qqGgh0s01pKsG7PForWF/ZFHSvi
zrHqEtmeeVIba2mxO34x8d4zsgMtkzTj2zofN8UZBUOnCdMFTUxscrzu3FuzXnG0ae93hb+h4+e9
IxJk1bdqu8RI8Z7kYru3KUNmLksUvxE5JtsuF4/1dh+vJK9Zyg8mUYEI2r3n/WmaWY9wacVuRg0n
l9hoFadMUA40NuF92RQ8vfDhQsy2wy4+Ge0bS7EHezG3sfo08BdsdVVZRHtx5SJXyrK7Z0GpENwj
aYAJ+6zfF9XGc3GTAN41iaEZ+Iu865mdoBQruYtmJBjToU6y7TAKhfd8qBtoD4olVVgPXiab7BsD
wi0W2Dr3uGGEn4VnDhj9TOvAbShHyg7DNbVpsFlHhHc0F23VsqF98NptP29j4lxSgKW3KC6lJ4Tn
iUSCbCj9TgfzGSwIaSkU+/lGHblKa9vus5CdZ1eK1wNPJaHcNFnFRvudxFpYtod+kY1GoZ+6SnYd
G4G9B2JqlOh6EOHYCl87ldlYLCWqLMbSN4UNDuoQPplNn3vTh2o783c3n+tGPQPNOjCZNUkMhDBp
to1BLmrMcmnbIwcIYBA+KNQT22/WOddEQQSbtk+W7xpQT+lxy53LZ5OyykK2aGiyWeup/fo+oAXI
5rvJlPAOaihBtKnCQQKm9cShXKAkzXhyTtyYdrI3fxouUgxyGPKF8jIwpXV8ty47dJojFGPUAzpn
U4ZmVFiN3uUboACvyeQClXHeyJQEuGgxh+m7aByOGNNQ478cnQKHwm5HZfSrrf9lSSfUn3AWVVq+
D1SBFQLIKgHUb5eeqlJeCFB1l2PeykbUymqNAnUaAUWTt2Qwmxd+83WI0UXQ8uE8QRZHWimLHCa4
IGsmgYr+wRAf1A89UAAGpg+2egVOQ/ROmXMEmvR6S6RRYuXN5xra0BxaqB5CRRp5A8qm6lZb0xfR
hp70zNHne2MSWiH2aPnB6EgoWDikzPzZIqtcMFyNOMuORubVnQ+45wLuDo32cOjM9lpCp24E4Pbm
hKGqK2Ht34RwlohGgUdFoXgrJkAnl9D91SHsIlMWMEbdS4Ysx+eJKwifvnh7b0LJMBXDfMVQHpl+
qUPIZ/hTE+mj7a5BLorm4+nLt/1AnWjNOpqBZwq1iNEZTsmOzOHczJF5WRjWWdSbG6M5NjdSsCvY
MDhNQfMm+ke0f7P17pEGlc79D1499lG+oiZSRRHcfK4/cegHJbzwnlAlLygiirnGHCVwJI13TtN8
/WCfzEIqKOkapV4IXWDevoHsDGu09PxBI6GSHEGRmxz7e1+TyY8RE0+yY7XAHkhAPPxPEnHJflqO
qKOgpkIy6R3rWOyqBZw2no69vyymnzMga2/QrZ0W4AW+9GkkFmjY07kn3/KfmsUuf4DtIwRtJl06
RhRAGslih/DuXw7YGGg5wJcgyPTunGAw19L10G7XTCVfY31H5YhdVfEdxVtMrEzXa4qEUdIOiQZJ
Evi8YlAvDyDQdj0rd3nGksjS5RK3SAc0hn4t0He8YlYop2kgWHAbbO6a0FFEnq+koB9ta7INqnT+
4u7I5fEFrGU+xsjjh3mmUt7wvsIG0kQCJMHoNKa/XW/B0C4F5/1TZqlqqiJmkbhJzjYsjcvbImfH
C8P1v35ONUVbnCC3H2Qiy73vhDxQr1Pg2YHURsN1aPI2BEJHNfIiXx3DiBRP7rdrsVYt/9K+VMdO
FRlH/+gx/V0aWddpTtDZAb4TNqrVRRM4aDN6C1OH6vg7E3bY6e06aP+6VL14wXV32rrrwnDtWdRb
uitlSCEJtwevWrVEUljs1YvxV/9jc9/5Lf0SpOvVxLimAlm+uEl8R/py9Fn44vXUY1eKaOp/7jy0
T9IPef/5RdqptS/8D/hHXfgIcDE//mX8ce0OssPCOYbHliVdoR5ckxRBXRRSfIly0ppcJru1QR62
vMGfrFGx4fAm5Zwf4OLKiUvLfF7BK6UgqlsU8nQdpiRfKxaJ4D83afPi4R0ivEcZN/zy6DWQlVqS
1VMmAf6f+cPnwK3mXHBUr32OFnhDED2m22bFoUC90GTjXxJHuxsEpxDxgdzpgU0qxvo5I5/nFMji
z+89mijKWflVqQ1ZxJ4PRfkSv5PcbEaqbgM/Pw3Fr4gYAb5gJGpgLIuRVBYzZQKei+cX1EoewR3j
oqymlv5xRT7xDC7jdzEzZQHvnB/UbmQbFYvBcapRHDakKGUb8acsgJpGttbgRK2GXUAOxoALAbPg
YOzvYxit9o3SUqhBawTqlW36noyYyFy3kbu/Y7Do4U51neLIf/obJs/e5DhJPtU/FkFVFt6mVF9s
lH3eTejOxbvkLRaUF+nwJdRFZTI/iR2mHSQfXt9bXXRhyHE3BckE1D+ton7HckMzOJGoLc1OXZta
e6Bjja/L+9j/Jyyud0OAdjwCc9r6tc1HCQh/w+6SYPvq3AnJVoWeGT5g3uMxRbDdy6nxiIqg3wMZ
DGz2v3fBotGLCudXOFnzzBDx0qgtalqDGL5P/8LlYFnAwhFnIQ3DMw3gFXWCfNvIUB5jrCtyYh4g
z1cWvBEMoSZIsd6pme+OYHN6qfrw5qY4+cBxUXd/rVKWuHupmZRN53fNKhkE2Bf/r80vd4OK5sHq
D+DDhrWKFN+DC4Gs0EtGhi0RKiWcJZWHQELcv1m7DNWv8RGPjct1iz7WbLaLKSS2ok85l6zJV5tk
JL05K/IS7cJK3K0X573uBLyPgfn4cQ+HMnI44xjgS8tlk+ibTSdzhZdawJKK3z3c1N38P6YdmiFZ
cwAd373QQns07fCpfCWWvkzr3plFmuFcOrYXBqqVkYB94UylUoZsLlVwCm5jYS0i0QrOwjqnMLmu
S7vKvZMpSekIYw73nZN9RCsqVQQMTf7TxZbAZgU/8PE0LspjkGQQ/5SCrHDVCArmgaMqZtp+uqs7
mLBIQ2mP8CX86N7fVkQZviVF391AgTfpH8mX7tWU/lqloebjFpO1JV3zspqS9dqB4Y6MxEdwwOjW
ucFoCH475HjtOjyJ2VF8Tcy/dsrPnWGi/VGZuV4Pi2sk4q0MoF6kK/XCW2MQi5FnH5PXlK7Fgo0y
KSVVuuhVWkkmcJwJd/beQrqUEXoCRFEZQ+8i17/7nkaH1HxUSLM8u66cgyu5tp8vj/MmTYbF4o8K
YqaIFlR5ffiOKEm/LveA3pDksZqTzGUA+NGOOSY0u8Bk6W8Onj+n6bSunywKW1TNArtLsnYIH5Jt
e7z3SZ5yRwt9B9y1XR2WpXSNB1nSWsd7tCLZxHIQP6ZRMnXprI61xPe4f73e554Bfb+2NK3d3O+3
F/rKiU7e0E0HKv2w59bEsNcAHZUS0e441u5oPA65b1S5Hc8aRrXvDwqLn0Y5mRIcoB6XpnWe7N2Q
nXU50OOcaya000erZs5DntF0vTElUL0PgY7s/ly28DIWGarYddPxCDjjISk/dU23Wfmdut5Dhdga
BV2rt/rlEfVCN4cZYxPuyEPR1Fz77SD914OjceztjtOns2sSsgI8XpyCW+vs3EJheJdxNyzZAHfC
dMuo8mygi9jaR55WkUUp7k4UA1KObo23KUR15iWy6Z66Gwj+fU3K10yRxRrO9A38wEAyE+VqVuAM
mNSbOIKZ+pYJ0lV3/MPL8cCQ9s5vPm2naHLsSCeEW3hNERfQbZZcy4Nl5tlBwVzPmB+qDONquV3W
fiLRmDV5PiW6eM0fAXNuF0ofVTCKjXulXCdmELeMQGlo+wsX3sRhgJWkI5NIxvNUuX+uGqdlYJ6J
M1eCGiUdkiFfl5bGaOvg0sLp9EFmOCBnoxIY3NhqA9U0doestow9J1hnAakJckxb4M9DmGTGjk7u
DqppMSc1GXEQi1hQQ9r7/vJLNRcTPNB+be6UnczJ+0ydGPYMrSJD8n31L6ViGtehZr/g2Elf8HMO
76d9PYDK4oKvb0LupBNCSzaNyKH0M6kU70BjHBnCZvwSnVI9d/RiyeVMHYrh1EWW6Tf7ZLtfpXWl
3nruquSUx0ZpMmSuTY2r21XQhu9D4wYHZoXsgPL0Rfy+2WcbJxq14MmiXG2XKfhZhKSuloI75fCm
/Cr3OzT2xrOi+DqiO2/3CKFSD71LpcV1XNR3f5RJoz7arU3sMdLKXeD8zrsR26Lq407ElB2VAoH2
374Sar7SUZkAiMRmUYhN2xbStp4429fdHEhlxeZ7oJfr7SNxxCAN2bcwdhm/p+4svhIcx13ut6oy
qT3o6vvnVWcmZi1DAmI31WizdS42KyQM4tn9UYsJ26AOfoBd2I1FFwyZh9G9L7mOpnmozFR+jEUh
YZwdcp/aE5kRg66tshbQOqXy/PUlmrij9ZxPbkHmH84NCXvhSzYw7dREKFBl95hZHVjqWB5ifYsg
tWtcY/tQ04cSZ2xcs8ZTir1FwzL22Y60bGTa2opyhzr5gwsKlKM0GZP/dRu5QwFTewU3xhgorbrP
0OaJe9zzCaER3BQ5n4N6K6y3Uaj7MXHIAcqATHX7vcavFT8M4oS2+DeSwvwkh3ZqDeMpiXVcmd81
iEdgvHiaZDuKpkQnJ9cfsGgF88gZdj/qEJTJ6dl242Y9HZGrZjCe6fmzHYlMdVIjSqKiHwriXngN
HJNoHQFAZ7T3oL/NFLhAgjV34LbSXqVmp6328EXbOCMGwHZnXoCqaUM+us+l7u5+0WYWOW2Zbl7Z
nEn9ewXCMxCIxojkOxVIzoTLKLoirRY7Dnyu2N7bFumeQxBDGLc1bDaGxE8TDtywigv7h3mIQDu3
4sdJ4IJemyHGCQHvJJlcRwoim3NumXmzy9vZukg0P+hTvphEXBA7DsvRkJDKCw+q2y6cpyXmHNhT
Q96ixSvtDIQTTYaiEK7RjKpU4NDBRgW4cd6NiEAlnj+HspEG8klhPeiemjCi29SZ2sOUA4bs5QrJ
wk2ZngZH72Ml2sl5Pw9fa834Ldb7TKOmmK6eCW6qQoJmth/TgQ4SA/He/0rPFT6yky7XoApo+kKa
IthNTw0YW2S+7JWHdEeKBNqK7vXTXVtcIZrRPkwflfPO9LJghw2tNbvRfYEwbgDZr9pd4qwlqx+V
N8dfKoORpPOfim4e4vwxOklDBOgLb3JPWF0MATN7K10tJHYlKWrMj5dY2AeP10KNnah3a4qIaeER
uMjf+YZlXokQOrisKFJHPqEzk2yWcohyhvNh1tPArmo99HSLIYwsirzc1MqBahjm817ipi8zIDve
Uc5zjZmQtuuemMr33EcRmjskWSM+5CNV8zrIV7xftdxCLRFhyuKFvMFm16jvFPz3OfVO3PIBrAPt
51di86vxsIMZu7SmTJ0wnbk33aCBBky1ReZUY0OcfgjOBWnRAqOvxKKMicAn4i3MFAGAt49swsi/
vS9/2qApfHT1lexjjuopkYxOmxuak/m6gQ0f4ezbtvCcsP3leWJ9ROneZMqG3FLJRgQr/KPuPMa2
sI7DfO0S6b6mN9J0KrACxnWWJKskMCoEbbyc7smuS3BS+q2TitdmbEvrd3e0vl3B1TMPig9pGwdz
fQ19Nr3uCc5NEZtSCoL2dgkgM1RW3wrnsvJWfG9xrWgZqxvlRkfmU0G2Ntp9YgWXKjVJqySS3dy8
xnp3QSSLYEB/utPwmyEddiKmE9Z7VNo/MdlW7tCd58R3mIZYHsFvKDqJ748Knc53KbpQV4poLCpd
kb1kGPWJlnQlDZXzU9kIWsKPBGItZ7S/7KPtcE9Tjy++uUVgbJLHn19VeROHDR1Uz3J1T0/U/e66
EVPe4gcpAATfxr9unv9FpY34JDyYm1G5WLK5aw+WQOgV3LuQB+wCJ3mcRZVKNQrgwlJ4h50fmqBf
zeYiJ5m3SCb1/seqjqDnzdhSbM0rD+ueHuzMbh70x+2C+B2JhVIjnoQiYHY/n9dzr4BYNX0Qi7vt
NJiFHICzlwmvIKzF3ZOKSaDUO7G/kYK8pAhxqctpRPnBT3PlGCfhMfIMV3MlEY0Ay0+00dKKaOoY
xK/XufZXlRlqL7DEZSrOjlPd5E98PPVA5I6z6G1veU6HLVj/CQR4++f4XzXUy4g8lEH95Y43zZYe
fbN2YtKEwHXPMf+SYvElgjIvYmwpz/XVs5C259q9GxedyG63hJheRlNrKXfLM//C8lXCUL9Fwfo7
F+zoVzCZYbXNQJPu/13lrAwrbQNx1TJseZcqx+J7gyT1CfJqGY3KytBRkM4TQ2nC3s9lHcAeMrOz
hYAY76AcwnNEsLtdlOnFAldX4KRNTYFY9ctNRVQi20u7zL+oTM98ypR99c8buMclu23971FjuP6i
c2/UxsH90NdmNMTYOKCRzTOR+LtclUllnuKTTxrpdnSIEqmcUxU0LrNoi3yIhV1trzB2FASJxS43
29dHEPtiM8LszDBhcGTDDIzZY1UHqJ7NhpzDCHYjsTHcBZyYlsb0QKsRQn6sHHHj91bnVATKhk/7
1lG6sas+dqvHMOaA6x5U45+yCQm1giDNt9ip8XBE14VbMIbi5KFtTYOUR2aNGPjOdZH2rE7Rfu44
mPOaJFtduZ+CG23J3yygNF5hf/D/S0BR5he2qmhlgLhpeVx2AoiPNQfY+DVsdoqY+Dp1TbsJDdN/
C5QXRWFYE3d3/lAvbYXhF3pdao1vAHDBhOX7I9geDuIS7lKkkeGd5pRmKaAv4RNnmEdJFQzxCxuI
B7XGKoCZ6iNQdhJonle8R14kvTxLLNIaSDJbBxPPFImZn4L7YmNtCD7hsk1vy4He9RJeV0pCFL8M
v0G3gCunqH2CJHIykN1HICdGOsRsREOC9urET4TCtVDRDL6aVnjnS9yP3RMRT6PKGsisz7l/GDlM
rpqHED2jcpvpaSDOaNuGdge6OoJ3F3jRxShuTAOJb6gjQ0jvr4j319MFHvgDteFm9vj/OC5p/+vE
z4MhnNKpI6ec20UA8JwNpYRYMMUMlu3SFZKrFlupNcCothsabfqCoQwNzoyNNjpQB+YJIASXw+OI
qrzOP0GZI0ShKFKrODsb6vt3/4aEHUODqQeH0V5EFJ3jLzJTLJL9+gMl9bdOvhc8yI66GnRebwL+
kjiWtfRCKOX7AXrrnFj4PFoLNLcVjLXSCrclczj57n41If5EIVJwZ7BhgetzpmWw7BPPjHtoBODg
CLCXxysUM53VxcMkRoWkn+xmds6iHIUa8TNUVobdF1BGVkGp1NysXWaep3mxjOhZw6RIWW5kq4kB
ULZktgKYKzTro2bB0lWWdBtSA0jnpLnynIge2i21lnLWurD2KNg1if/FMSvRafnrRDn8o0c6cbvQ
bbZd3CaK+xlXNeeo2F2uQ+ApnPOmICiS4abiwjmebu2+bGsRCwPuCN5BdO6vQdML4PBb2dKEMMQt
f9ZqFG+dH5BlONdWnOysvICL/Nzk5xLAobqkaZmkRpfY4xUVLd9sr45OZEL/fAeYsUp7I0lIfNKS
8oPQIp+/fddelzFCxRiS+z8gh8rgxwCAcsqSoSeO3b9N909PuaSbca6A6wB4XSRrGVSbKOL8Dhsk
q45eWZC5i7Myi/4EmOznzP5E1GKx3FZ1S9xn3X31wVrrW7EqguKghfd84FaKfY32fJQ8zhJWXQJx
zUeRA2IfBe3D9bi1lJPHywOFYY26YDUE7GOUQwkIjid7hoek1eBOK1GmD3JRV6ssU+j8X5hoOIPy
VJsshVMkrBdcer7Z6jBlJfIgXGxGGJNDli1UevQj5edSUz8xj0dDfyXSxuJMwxGM0fDqjx/7zXPD
PeTCx/MFwP7b6pc5o2wFm2/LaLJBwr+1Y87sBl1f/LxCvb55Zpd7Kx6JyJeakL9YM3ZJtowhwELN
MJsARYZmRb5SyOcrLWWOLeqU8PgyLrGu0yakyCkskigICb+5hwkh5xeu1Vmvv0mcpdpejhtIFgWv
FncxjztPO2H+E0BKbWO1Rn5VX416qXBzj9jkM/wq0IAnSLmq25jZTbeI89GwsBKQ4Hw5opWAymlQ
Bb+r4jXX7UWMJ5wdRU1xGHBgTYZ1EmjIVCdqfYOYt/Gdb+tBZnGQjOcDLagu7mPG1rSocDMHGUJG
BoyQAEUc+9A620pv/6KN4iNY/qRsmJsZv2UfaQm3BqsLbk8E07ZOeFTcW+542djbIoAJTkgWHoG0
7MMysQFjCu69knDC4FZh42LWRrIUUlwpzyRNxhc2yoFjWXXiwQVg6R9DBIESx2YXgw1/ZAKNdaYe
CG2tOrOtTZI9ukcDln5vU3SWF1/WyzLK9qn4HrtGb3Yru1rr55CVEqhhI+XDPpvmyRKNfcraTIoD
8mKqSjhentHBTUB8wIxaQ6qQAbMNRBV6JnBNhvgshSCdysMsJjuLC5vg3YfOkS6PDACjXwUpjl5p
IUxe2ttHQy0JQs8ynQoiGe2UHpB7GdRrAsXr3/ceoNr2C1dg+XAmZw1xzVARaEsdpuNJbar00/QT
mpWOCWtvWqxlXEz+gXmqKxE3viFZ1KKd3Uw4LtPbpglkrLvfanXFWf/BnXAVE/AO2UCE9C1U7qvf
idveP+u2yLAThtEqY6f+9BvUDHxpYqPeqPoH42r636Q4vwT25P0QlM6pGArkkfCZrdt1I+seu6fd
4HWir+x+6qeHh4Tza+z1ZFQiGsVHoDr2xxdpXWQCjcpOx0F0X76Oa/YR1SlLwsT5WESUuYbq8JwL
gIiilVpxmOLK4kyIG3g8Drzmvng3uasY4M2M1C5NlWfq2FtL4XAskUPnTTHXnlZJxxRxnQkGrZJy
BRgmE1x6E+RRpNnBR9/KEA9AJmgDBjJ8QwWJiq4LVJ58SOzQK6bvUb6EXrPJ+V4sEWloTQnyyPmI
v5Wr6rCaWcG8NVyxrLOpC8pav7cT70UrvHA7NXgR0/OtXuuXj9uL0nwShgY07YwvH493xjaAe6Fz
1IQeg4LfMHfHqTc0/YNWlbLknd8X/7p1PFsYCTRIsbwZ7396pycKH9Ntl07SVWcgjgCZf9WazPcp
2LLAUl274C4/ryg9AhgdDQelj6fbDkF4P629gIh1D7Igt105r21W+NdnphawQoO+XiK5BjJdliRA
Dhof4bRZLQfE0jC4i6bCe/8HTgRrYX3tuuyJu+IRn64Sa5dnk6dIFqc1TNyiGBMowf9C7VHVlozk
NOXuzJ2awZGmkV6oUPAxG+LVR8iC2yCqzJHNUGmXXd3/Vu++PERY34YOaIboxPKlKM+TDhpt8LHh
ctPz+k4JKvhfwn772hkcpXDexv9S8fQZ00wj0fMKUuz9tQ78CvcxhRZgxnksNjkB/ZT4BS5XfRNY
rdFB9o5ndN6gmW8vWRFQgo16Yp5TiZMTFUThbpfsO1nyS8GfoSHUFn7E4YaeuCMkzEU5H2hjEduG
tfdks4CaVWu/Ion0Mo3f4KwYAjcojlo+CMXle5E8cT48kcqSZAwhEJZM+gjDWCEQGsceescEcmyA
Dx57XRwnoIby/45pxgncdH7fnEHGCAJEQ8FLKXg6ytKdU85mOGZ9I2eCsNnOdQGj+l4P3yihBw3H
NQGgSvT4K1znTOndEqMRlAGN7RKV2aB+n1DYO8c6lXJ8IM5u/qPEMcg/XMGQhTouE0s1Loh+WboM
e6+f+N4o9rGEYZm6nw5FQEJZ1xmrU28YtR22QR6yYwGv1Jcz4a/kPdpOpm9AEd1IRnC/1P0lyahF
TAV82KaevNtHL/uzU310yVoIt/2YL2ICahOFeerBKMpz1YUeHrDgOPu2z+wYjIhNXkfWlJOqWmY/
6hOSUVcdhqs2cV8Q5FJZHIvqHRDHjOnKjcN1VdXnqMtVRnnzvF5rZ+rH+JO455+duuWmTc36widp
8r+98o73ShqrsxBNUieZM6TyRhr3zGjuehdcM7ZqEn+4IUtNEntyigHM7ruT3IpfusOMc+dfzm8M
XUUGmK0ytsLfziPca8vVtlZ2B0B5TUi0J99Xjgi/TB+hmUBklqONf5/j1YJbpwjq3wI3Cn4FZFrr
ZmhrDTd/YNxPaFf7Lx7sw92pSZeagt4nb7eRqMy1CfMnxdck2Jkqtdx9OOnsYF5UykzPTt1YU7Gn
ZRT903QEhGccbvBrEe+rngBBiG5Da6A0vgD1s07XB2gCr1CxlyoML7e4rFll0FwANZnka3BuAEL6
o77QxmULVXmaS3IWKjY5MLV5IT9uFCOns5962yLJgauzZwm61HHEfpC/ctPxpozB57bHtVugycik
PA9sBb4nkSI2JZPUAe54Tm9Ixe1zboCIaVclXeaoN/Bgzs7/ROWno6bBvZiR98yaWhSidGJKEspl
AZTodvH9ZH1CTiJvsO5y1YRs3P4O+c09pgTd2Q+7MJmFXXjoXJNhdqtRrkaIV9/nAQf1PfPDdqMN
hk1V62NK7hVz5RjjLDhySwXxdVlDFzspg35xAdCr0VJz5MD6rx6yXWhuKrEjxpiE3IBq+2FqrjCJ
c2itCnVPWxW6JyCU/lMNoA5ihGCWrdDLdt3rDZepXuSBRYGSiShjeefn+kmPWqmbVwV1lt3cbn8/
rfIC4Kkz4XA+h7ns5kWrxofvs09JxVqovJntuPOs5ap9UDNOK/1fTAHL8GLBAO+BiFAxtaz5z+QG
+Mz/Rm/IH0ymZTKnI7OCsF3KZgR6IMW+D0ZKNrx6N3lZKRfoHihA4kQ++nJZAy6ryiiNihTmIOfL
+UggjVdf6u1KqMW0iKUvPXe2LpNdwL7Qd8Il5SKUPsvWZjRCKaoddRkLWm/w4R2esmP2+AL94RRG
r368ZBl3ZZ49AA1iulyRHKKKaloT0is6nGA7hjPTWlsSOH7GB9F3sT898wjHWmWgExGwc+5R6Gvz
hqctMSvxc9mNjA0rt0DT/NyhKTa1BHE9YReUyB9mc7RIIliGd51TJ242WC30NUeaqAB5SrTO14nV
tW/h8Uwvxch3+FpjUU8PpSruKpcJZdLCNWgOIOe9/TNrM/UK0yVpiO6EsPC5DFv4WRTO27TCTJki
uBisWuNdl9m5PTWskyBPfn0GBJlZu7B9vPk+ECNQTuHbxFuLEIzrIFQSOb5jdkjuJbiXYcx3RrEM
5a2mO+6wC9xviJMNmVYmJpoafMOodNG4DbQxZ/0jVSch6G9s1YppL/vqVRs1g8NQuqc6/sHokaDe
mzEsGnNOaWVX36e0sOyGEhDnKiOjS8cDpiVaFtyVmEUbxEfPxTISO2ozCdP5j2EviKumivU+kpkx
9XyLbPJkrGP6PuuK1WN+mPZzUT5KK6tCKQlKAgU+SQXIElxfPkxk6qWzTlz9bwuyc/bn8uEAyJog
ffqyJVatgh9CPqgIRthdKVPWLdKTVg4M9G1klfSsNk06LwqRPZOmMhkJsm+vudMMJTRFkRdFA21+
DC2tOegwB1vDcy8e3MjEGZkag5+i/+oKxLTyqB6Ti2w/zyb0oWINW2wvPhWPz7xW/3j5KtcS2npB
HHZ9SV1szX5w079QsYnQ3c273sxwt7eeMly3GdaWKm7a6nZ3jrBSvzTiHzC6S8ZHgSCseJg9mPWW
EGbmQr/TD/temrvqgISYpn7k5Vun7+YE+V2fdJOWQIdJIrvmrBHQJz0e5OPEnMleNYAlrTag6Tm2
5Rkh4VpVLuLOPKwWjswavdKEoxM3E5kzJTrpZnQYja4WdXfIy+Sz1JBaUDwP0hD1aBWzy7HOtRMi
GlfSKc25LJuNX4wpM98Wnk845LUaosywG4DJH5LBEVEb7skT/bkF+QJw5DffqkPfEed8hwNb7gUr
R9x1cFSyqaMkznhRxvbhiIoiUP/G3usrRXMUXDxzF/dHZXN2arztWw4rvee+8pLZW8xgtFdkuSqV
efjac7JxmJEOGLfYI/88mYd0vwjDF03lr6AxdtYNnQa0MGc4RDemb6SEYKOvvv71ukw9WwvMPsbG
8WMD4ajx/PHEGFiQ6SU4eXr0o2VR5Ww1dGj6OpscRdkv0jgXpWSbGiLghyEn4nMQf9WxO8Bq9SGu
4N61OGu+G9YA3PjoFwxqaMF7H5MkPPZuSfCFQZgjuLAeQX0dEX2z6EJz5zFxdY/4x0765x8OBTtq
QHsAxVwYNcH1esJelLbKHdTx4bPjYrZz368Gb87kdVLHMZ8RtaX+nH3z8begNka62SQ3cVdHAppT
IzVZQlPmajHkZG6Z1NhW3TxFNc6fLrRaBVW10LLLmnvuQfhwmkn2knAySrmYWk9sZTu5QnscMhhX
SuubVCiLYhkARJy3kIPh9Yl/zGytl979Tt1iSQarE43dnSnwUQnMFBwKLeNz9UmBp1BDpBF6iWs2
9LOnumm7V98v7kmzzWUawKvydwfpn3j3hOC2do00YZyf3tBM3RJ5UyltbEATsqwXFC2GgF2Q7xaR
JWTpnrWOj8Kz9n8+dXDAMOP99XzD8scveVYcg3esJLBJhnu9r/7pXwM5VXdpS/DAdJpXmbbVTz4L
mfkoEqHCWrPIoymwFGy3nT8/+W7JIWz2rnVPhSIBGTNX4z3oBxBiwcjGoS5Tx6/B+TxygCBT8W9/
UP5+PNwmQvliKvx1Y/hP6pbaQpo+qBCcOn5lPxRxvycK2lYqXd2mhP4qhOguIhKYFH1kFyosob/V
rHnbXn7PY4PFAEItugXsHpH1bJdYHbTLrON4tPtDpQYqyRa6mDWPxfc8KX27JSepvWrFDI+9vJj7
kVzbtIDmEHIICrBvbSHg9GfT/9neLK2xRb9ACvw6Cjt7zLfpxT3A0mNgBzZ3SRfkhbZcndBLBWPk
ldYX/+YkraJldzbeeFv1TA/Phb/qxoqM5yq7shHxOBqkvxIvjH/SIO0v6GTDFhtTgUsnnzdOY1Jk
wXnFb/iCRLB1cDN2aRgaKmgipziIC04jpEjpyM+m6skYwaUq4QpnG6D9F6SYJ0CVXFXwwm1wRWRH
a3olVFUlbCKXhVMNqtLuYuIahMVI/g73R90pBhU0VZqOslC0swlBj8kVZy0hMi4wucz5T2SWnucC
ohQ/fb4VrAxTjyE7DAMvbY52G0Ck/jXOwTqeGCwYv3cbC6qgfuyRfZFCIc0vvNUzdkBV0y1cZRXv
OKPEYjPRo9vqhuJwh7ncYRdaz462fb9kxoPixgjpo1SelCKrB1EvIVuCytyLy5jb8BUj43ghgkkU
rlLP2+1ts55q7UOc6xYAcNDVyv0TyZ7VDoZAKAs81KFCrz3WkAvjb7WOSTEkFsz0mILMw/6fjLBD
Dnz4N7Euf5v0n2Y3+XDbhfqlvjfypVDm+800kPpdZ0TMGGM2Ch6P1U6nJ4DwCjwmHdLK8H3TAZZu
9B4JHwL7iRdwwkk3GVWqLZ+xDibG6w2HkkDCfoyPMgpphkvQ70W4/4ovXNdaRYJVoxN4O0+W4nu/
caDHpyNLammO+SKOsEakR7qSm/AAr0R30n++abdmTTTME3XWV9M1JJlGEW/c56HnA0k4RoLLJq7m
zVrIrXgQk7QQ8CEZMUcLtfxDCut7/h52Pb5tgdHAPRMzhmiOHPyawZXHFKs/ebp8s6yJO8YGTKW3
OPNmQkNFAKeF0GWZJs3+N7ffeszDdso/u2+108qx/OV589OKimFpmHKBYc35pxuNyvzSpBQJ+ssB
Qwu3m/6Y3fqCvgoP9M04EOsSANi0iZCiLvFAQaoYSPDq1XsGJ/X5XJyePiYKdpatT9EbQgrh+fMp
s+6K+nG804UB8hJcLac4hbMMEP4S/x8A1L7B0z8/1UitUP8hEJXdywqNqVw42BWm9pwnMG+nn4DN
A0EZKkeNWLfaUz17Txd0taxfCDNn56WVIBUDCIvPlaMojZec4mViBFyjo173RZqGWrbfJNHhr9ec
S5eUhhKT7vfIIfg1WrjnX4XuE1UuVnCJH2vPB966KMMUesMEo2eAktJUOLBBxoBlUt8DVPH5uYT7
CKwvFuKZZfM5+/GZaM2fCLKZWQz1OvVtFRadHQhyBMvRFWLTTt0N1Ffh7H/oH+AYfRyWa4UwrXKo
GsJYfAIAd595cx2BGihsZbxPj6LwqIjFpQeBGIeYlepu5mTiHUDduhGNDrNXbig+xwh1FwMH55pd
TrlBGNo985K3CNcED3ZGz3ONDKWYTuyMmjFoUrm/5XjxdMRAGzXbEAxkH25OkqihaLm1HUoj2Uxg
0Cn6sFCrY8D8DNudPHYtu4VTFwLkTXi7Hn8/cbo4RMgoo5MtbjZS6cqf5dB5L6sUuzq64pASRxFz
3+bSSyHD61dhdlcStfk+Zve5hq8iFMWD/BEe+ktAMe7hb82nyTs+lJOMW/SSQxbjucZvIGuOqBQJ
p8poJ3iZqQaPJ5xLcPKTQWyYb6riUTTBeezOdmAR8ys4Rvn05+jHyTtZdtRatTDwsKBU4i4LBh81
enY+EttTtPaj0j+70cL2GxxntcMICwKrZvLxi2wzO6Hr6GjNiZ6A5dBCJsHV09VH78zDU+p8a5PX
ePpMPZx8tfNu+RTvKeevpH/edhEzw9IUF6cQ2MZM58faikBZ8qrPqjQoEZgIiYwARrvsiC5CjXs7
tZP7BoRYFdkUA8Cpu/cbB9sOMfL4/hb+tQznmIBvTz0Ew+G6QUNW8TFRJE6LFAlMwgx10tQArCpc
4Gx6bOV+KMTKObPspOeVgc0z3sfMNFh/P/YrBw2m7450H2jEZ6Nw0ZZY7DEL/cbFB3Qc/hnlHH0O
30nwCReN5Eh2PRn8LPV2Petkdop/z0tz7WwoTCSAmLpUnPzynq7mEgRIlug1BtmhO5iWkEZE7hvJ
3g3CryQ7y2fwE3XuftCFBIbd/gaFs1vBCe8UzWskxB9A5+HaJUVHlNMxE70f580g+KwE+PXNHpbH
NNm7Iv++uwsC8FPwYlOWzpzrRUwuZHPqdhtOQVNJZYZl2eYofj77mINodWlK3IwnmM/dBogoYF3Z
Aqtk5UQzj1HM57tt4yuf9Ulud2CQaUuRHp1MJ4WLsa/UlzkueSv+Ngb/WtN0ZBX19PYl5masz4/R
ceuT3N9RYBS+VuJubC4x+Vku7xY0CwbWk93jODqWZJZvyIxpwGvoK4b2vtY/ja0OthNXtkHrGS7+
JTgXOkFO2V7R7/GDKSCmPpW0RcQO0oYgEDTs1HH8Q7r8KvaKriSbnp+Mg9ORKoRvEnMqmTflJ+FN
r6lyk5gYAQAyjNgLcLrhXJEZVj/fcpY27Ab5KwApP/AhM5nOX5U+LPKOwn6FuLn6CVTSsP0S2xmv
k5kEfTlBk9GnNArQRNPZtzPZbtuqlDE03vrnK2uZjWo4eEh5r2FTraSoY9/yVoWNKTL5zj6HZ4dN
BRpIUbZCUqOIZuCGY4SJo+ihXOSLTJYNkcGAxzSV3NxYGPwIB/31ZO2Tumhp3JpGXBYfoaMKjqU9
kkJpv9qXvP+gIHAwgeyDToEkce24weOdY2K/m6u9z8vxp2379D/IqTLT/Gn6ygFWW+ySmi/GMyb1
lAkLL07EzE4P/uSe8VQF5NLIXMXWMfDnx7+gb0RTM33dSYSotgEQFFYKWc3rI5KJb6dy7W4JZy86
i0NZsf9O/iKZkJl1lDgmlvrmGX44KhFegQ3Ar/n1mapp3UVDb6NJAZ/dsPwrud5GwzyAnAImDgic
2JC3Si50msv1QrXfRsOYokVoD2gBpZMIBqcjltFQYe2Jde7Ckcz3B3DYQwfJsRrSXm+fVkCOyzGk
b0+1kTAbWU8EhUId0hsMa2tPHT+fG5fpHzOi0p9LCpjCTXAkhQuiWvdaED+r/0hWoAwZeiUbl04d
oPgwRh3YHxwBdqhJUh8zXhkP9cazH3smmVuU8Scw2I5l2FKunU/nJJxrPsGS3Q1HHUrbJlYV8W0S
dcYPgFUjIkkJTS5lhKta2WPoz0Qj6dhnK1S7qHmBW0Ht7CpVpmHScNv8MlWoQRuU++jgqcQerXxI
f7jmyBkefEbORt995Ed4+krgviLu6INTwbgT8D/x4SpIVB0yFd0Q0Z2teAZzJDngv+p3SlhG2XYH
WsJpBvaRGouq84pDxqnwFdJnalRKY38qnxaCPKzEqhoH4uqI7qrb2Yqi/VIrvcoNNwC8qpNWgGN8
qHypyTP3vhyC+0HOL9PiTngr81rh2JuLep4x2G4ZadmnfwjE2OpDfG/868pYEe7c5yg2HTcHidD3
s7MgYSuAVZEKbDU1h81KBTSj5muxqF+FJ9wJv0qvB1d55UWrjz/4cffZK/5ugOWFHZQxt3lt6ziM
2aZQL+/TD3XjRe98tmtqE79Y/ftuyv92INwV0/So7GMdGW5HbyBkSR6wY5xbrg1unihnXcGJXaga
MjzyWDNqpcTSuRKve0alq+hMVH5aRCmHvU8sSUhBJX4DkarOt3bpu5c5WL7u7BHpBs5Il3Wo33d6
YdUEexrsHdJcqdDS6gNdaEiTKPy7R0Np94ELvmXm9SyHcUQ8URJu5jSH4FeNKDUNstK/y3myGOYa
GqH+SBzMNTP/YnMB84AksquTlRfRkNH8JRrCdnUI8XdSn4Jk2CFGpCCQUqpIGYF6wIEeVLAgnv3A
mD5ngF3GNtksLHkkjakR49C3ikZzJ3U1vV8hop2n1bxJn8yWFl8dBfRphok/AMKrkKRLFVzTKikX
sWPbD90uvmzs8LGCTDpzmHalKPCqK5mVHNpVndWAPn5OQ0arnYkQWxgArY8i+U95NQhkHc/TP+aN
G/dxklZf07PVQ/TX8KFVAPKaa7dV+3KRL4gtgKrwajBtHXuP/8hCn6EPRdjtoIKCmX3WyzIRddDv
ka1uQwJyYujl1VSnMXgXwb3/djlR3lrMNmO8yuRixquGyABxBdjBaZMZZQ1ZcodCwAHAr6kyopQK
s1CjWc+hZTyJhHSd5hodrGy/R6uR5cuvQuPylCGebIqMmTutNNmlCE0tHOGV47FWEwZeqc6jxu9N
RuKAoxvsWfwoQ2P6X/ej3XV03aHUU801OYiWBVpV0QwaS9iXctKOrk3tvKxXaqsZL2S/Oi32D+3v
acSKSe/Hs2+ndllZaxP6lhsMR6x6nP49mFIOMOg72Kqx11f18oN41OtrTj3CNsq8zZkN6s7awcEr
iFNY9TSleON0UmDBmKJaPriXlhOUVTow8ZyAC2+H0zGvIvm49tyS7l4cmP+EOyXAcNkmki6sYPXU
3aO+2nWW82ySGMVtuiwsQ8+D/eVxS/ku4x1bW6Kshmien0dhY6aI8i2sHyylaBbIL77KoGb6x2tQ
n878g/lLH1Gw9SQ9dwFDkWxx95LfjusJ9hhEQXhdvTtRSWHPp4GooScwLHoUX0PfxbQQl73lP9ax
TkkNPnZFYKOZDviG/yPiv5wXLlaLrheBouduBE9N1H1ckcEYSkgwU46dH0sdjmnxaZ7NBtdADmsC
7JFesLoi6qe+LYFAfjfhERnBYoW6/WusN3JfZ65M+nWUK2zfNJoAcuX67f0kj0N8EZ8NAvubfeyo
hQ947Uvcy1KgfC3bHXdkIif5YjEC6bV3BL6UFB4T9UI5Fbbqdr6KMeEvbhz57s4jcqLQq4w98hYA
4Lm06ys7/kTPSHQ/uS2X/yJZPym3f6b9ifoe0EepZI3Rkn3Kq9L95rtfGK9pDoLnz50Eum5PhpJ0
fTBlW3gIkXQ5sVLpAENKQR0UH67gRioygbexORKRvztF7Z4M/+JwZXGzrW2X+3MdUc7KkM0Mn94C
tA5TFHzilOqpUwq9NpfrZ/+Oju3Wdg1ckhAwNyEcLIBCeAXiK7X1GUdQVkgVsOtg60F5gRyhKjsW
/h8sSh7saHg34L9OMBF7h8wJVlS9dViXBHtZSj8C85SwCA6pW1piS68JL02Rgvm7BoqL5TixFTm4
+SGc3tHFjiwopv5/PbWJKGtukwRPR4IRg/arKeVlAXDymjaf0ShhdRgTDiMDF7CQYvSQ9u5YMjB+
X0xClmhl5zvnnLDkokwIsmyxKJFx8RcXsXEWMP26e8cny8+C6xHDC72zkNY5ZNgb1PioEKURKmzK
9k8f6ys6lZEFsY4ESNJrsFkoRoo7fWFyPpVGN8pboYyaZUgZush84XFa7phhpTAjo8KRSgQn1Vf6
5iRHylhjE964mS/pvVN3tyLB9KGEtt9Nwk2/ASVaF3VaBsMBUG3SrfBIVGngo/4gd/AC+zkejtuF
U7D0xWTVum+yYWQSWBOQwo6t7WM6Kic8OwesXVUb7S+ApM1JmdSjVD01zC7La2dvsAlYlhxeT1N8
RgyzucUcRFEVbc8FR77JMDgA1DXCygkV8FFzhWpf6JWgH2Nh05mM8Tj1EUXSxF7Ar9u5I0vUC3jl
lsvU1zpO1nGB73MDpq6eUdGneAft4m4zlTEf0vkkLUGdEm0CLYu1rGXUpyvumbHOxdJb2iYoniBw
PwAXsOaSICZ0PLtjT6AjHhDial/BICy70TonUha2q5m7HUVYmhdyxSFZ1g+IVjwdedJ7Wxr7NUV2
q205gICTLWBgTrbfw7zwtbcV0bPDLc8LlDk2vn2XM6m4k59AxQj+nxa5NSy5XCHU0hwDshtHTB88
W7rTYezhGV37qlz1dXPj7OsSlsmdCGE3loU9L0EmB9RxnPMGB1ACWuj2JaMFiOwzuS+TIT9sy4au
kA1DOeSZbkat2xQSNNtGCmnBxB98D8ggM1Z90gAG/jtjNXrxwVxqEcERFBjYdeUXs0WiZM203jZk
C/NlBA+MTqtqpxPaVZAH3hcjtxWt/JfJZcEOq3fDmzOn7RYLQoDEbSZwqhoHwFpiPJj5gLZ8X4v/
6yGT+quONkkNIiIIu7MjdPQKeF/1VrFvNlWmrFmnVlbZv3teDSss8OwFLbkHjTZzHT3KGm/j/fAE
sbNp8fZTsClEV/zMAag33a8plC4SAxIIoaqcdCt3jg1gyo6D5bOj/wAIgbUKHTyR34XzYSJ8mlnO
mEbMRFlYomY/fz697GLWdbMJH9Sj7uRqEeZ9CZErx26wVdSQkaeG8G01CriFdcshOGgZyrYASTN3
ZNEz7QhrqdGggGubt6tE0z7B9CNaADjeJ4FjF6wL1ZhbxK2+oSmL/mBzMgHFDL0WsxegROYZk0dM
OoVz59MZIuOfmV9a9pJ6MayNsTYXFRiIqdHiOUL48iAuhW2yGYAz+j3ntQ6clXwn/eFk/f8hYGtG
ErDep16Lo31TnIlS4l8+mt/mx1GUsZl+/iP30Z+1Skw1m94z/F2wxxl/nCthqXeGYP6d7/sQ+Pwf
otAOismeV4KK9xlMYBtJj22XgVdSWfebhss7lCcpH3LwfndCuQLqo/Yt+ZUAUHLfh7rfLg8EZoeY
lhgTzl3oFuWNwL9uLA9sSi6gItWyrDuEhDcZdV88vSbVFXIlhOgU2LWqzPvy56A3+L+nF83dgVhU
ameiOg53kl0XWj+Rcx/mHoNN/iIZCktxLUmUcI0iOvLRbuzAdjrP4KrGCNlUAIioNJ9qFa6KjJtq
UZEbEGx6y0YCbpOpaDOJTRxc1SCRxH0DyEO5qVFKG1M01FNBiAOKiaXTZMO2GbqXsFPjzEbTJNdz
ZSVSn7zSo0k+smnR9OA/1uGTenFMghw+t8875IB7nvsFMKGWYVyuj3zMRv1vPfweWW9F33clTzsY
I5UU+PETeZPmTna01wT7dkLGHibBaXU6r7vHNXnJ3d6PeRt2INrZjjZ4Fok9rBZ/2v4Lk0hzjvsd
f1Tzb5Ge63mPHzdRTN+X6XWX+PevJzq69Ssp0dkXcin6fsHJNkt8/uj9vR/95P1BLuYt1DGSIetH
8G+wdYB7HGJwfCXIPHqj8DahJda2Effq5nhuFJMr1T2SHAQRXYXhW/uYPbrUyKTBt9wwks9Pb8Sf
/GS4rJSyLjqgptVfZAJFe7zrG69VYodq/Futalhla9ag3cdwSp7hzi47y2iKOFRV1ggLlPhBcFhk
z4uZtHH9+ZvJavncvahfgf7LYxAcR1iOG9A51Mzhk7qpfwJG+ZYLKWnFnLgiBcq5IQBkln6Rq+pw
waWj9lDhti2DbTQ+QGmhxNWESvNebW4DyvegUCY4rUoTFfQ2/QHilp55KGoSA2uMaScIR6rN06c/
Ya6rpt3khXYxBI6VPGaoFrjtuzd2yaB0VLjx1qPuAVk/6FQAqTpcQ9xEpEF5uIPBdbP8i9ISplsB
HxTFMBL2c8cV3hKyJuuZcZW7Ygh/AcXPVLbpmQDIdR0vMJKMtJ4iJbU5tTA2h6e86itB77D5Kb0U
pT4aif9HtoOhII50Lf1QZi6GsfPvesWupeo2GDLpA5LBp+ELpsNfuEsrbXsCegNs+rqHpKZSvC7I
FIJIWpFRuPNE9UwArEoyY8vWTiLyTx1f9Qp9yWraPtgskLZvQJVFxjt1ZIrZwI+i6iKZEWQOtSFc
qwccP0EtbSn27U9LLKZBI8Z+delHidpFhRRap939SnG7Grdm5uWY7vnWaRY/0Ok/NplPT7p/CPKF
3ZGNTIGhtr6vcm5vCDhTG2RqnTGJAUE4Rdbw4TGwtr0cy18ip4htAJ4QUYJALB5rEZZRtDvc8slp
MOTOwcUrz8DD3ASdrJ+stCuDKRuUA/ts+5LjmcGuqdbDhP1j++6j8p2t4momgIhSTNZGl/ekirPo
7e6KwD3LgZTRAdmltts02R13Y4K7nIO44n2R8IjBiLoZNzTzxPgVB2PxDDwKLTcN9LDuxJt56lfV
XdBBWpAzT9hWqw6hhoQWG9VowLQV1RhwHXhcvHCWbkXRYnLcKp3oh/5ovcJLoY0GAIZSi2ZTa04l
3i+98n2fDqRm4g9wSDoBUxrIYjGs2+OxZ3LxIM6CveUZbkiHOHrTLERSQGd6BLq8wlVjWQF4/yjA
B3ZafnsdB/bfl+JrrB2dnv5irFzZwaUMzi+2q8PJ0vNL9MqRu0UAbW/w6Iuhk4DSNxczqw3HWsuw
euQeDqVDplRCqyzRHuhf2XuvcU/zHh3UWH9USZR3FS4MLBmtw4KEO4ThrSRlm6rvJDGd7UnuX/TU
NYHZvt7eUjzOzZopxaNl5LwEpn2mIBNBsy5G7VVFCDgFlaGyMTHa5rdWuIqoKndQwy0KJwMC4mI2
f5zn3kI9HajE5Sam5+dSqdtfWnVuaoWl/NM+zyQKQrEW7aCCnwQn3fGG1PMXlHYCexyV6wqW11/r
Z1z9iIJ6eScNpXcWM9YxYMTq35MzHC/m4UfraXWZUCmT/Cza3v9F6sPgDpHUZFL89JiLkjIOUann
2auFSpg/pnNyZb5Sjn7LFzoEWEsUk13UIyympainbUcfhy6hz2JoRL9RMDwtZmJyNXGgukjl0Jk7
TaxNyX9XLx1atJ7To63I7Yeuj7OzJHmIbeBrk+GHRRiwbj4GzrTgIgsWG//3cbuQqyl4rS8VdNlm
emiaKxsR1BhFxdHbx1d1wSa8up9orP481iKJKK+Ih/pummGwG3nHgiAncDeddt9b8rcmqtzATc4E
+eJyJwAVEHbF/gp522e+k0lR8WMF7dfwQiXAgR9r3iXCA4CGWGuVF8fZemErAfYCAN0NJNG8OHaL
rx6ALjlO+n2GA/4inXKLRoP48vYZAe1tWQOOA7omAmOc99d5xsFujqRJL1qna3aAaqS+XseqxkCx
6PIusRdTJe0wXjWf3Lk2u6HGyWX67XZb4PaaNbrAz86+ZcSoJaabuIRie2kdTbTYnu2b8MWcFDzP
MChaOAC/ftoiO6inu2gEheyJO5pJMtiq8DkgfYgX+U1l94+eUS9Oy197DdU9gYGxNkYtRY2FnP0Z
EzBdDlfKXJHeJRz/SvJgEmTOuViOrd7UahuQr5aD+U1eoTtO1MuX7c7Dubv42sxZDf85B+801c1B
ft51jOBFUz6ZNLP8p6XZlM1STybEd7lYlq1hjnBdljSZktif49uxs56fn6TovOWA/CMhk3GWO2vn
ZEcH4bnWoaZ1uNb2F6xAWkiuIU5B0krvNu6EiOxiTQkB1z9JNcwG0B3DRhxDQd6npp1jwSk3Gp9i
vuX3/aa8ppLJaK0Hj2GWYhNfn2ftHY+pbuBhGi6HT1hadD1x8hFFGgPcpPHaxIDu/ZuB7TIQMTmv
SvFTkiXtjSRx5T8xQ4p0Zr2a3VLHNryLtFh/Mjat8QABt/CDniRVo5TezHJn/Vo51TmxpabzIzq6
FhgRNG7q4UoIXdRYWBNIzCQZRmC491aVBqU64qcMgCqvN3xpPmCkD8Rwuqjb9M8VUz/DDotlktbO
iEGM+NGZinyWt9dQzRcoBvsj9hXBQJbYOllUNVK+nkO/0gMbePjuVmMPk29YfcvYaTpgfy/lXIvi
Lu3YGn8Omix0kCsaJtLqBPZGKtucj0KYQYL+SnxQFGNmGl3wqdUuHVKV15MxTt/tsXV2irHbG8We
jMYIRLtDX9W6WZD8qo3B03dtjXl0mW5ZT6hOYUhXqH3sCY5jG/axXLF5FZfeTAaABsJhp52I9tiU
xKe9cMQup55DuZo3AEfyabZHzi7T++Voj2QwJdk953/dpbnVHaZMObvNrh/LKW0iQsp706P+yDS/
cKgNaBIhnxBR+VxfithTUPkN3H+1+7tTihwZj8iHj9LhVVzr+wunO16vH7LKOwDHOx7yaRJdOk39
tEKs7QWPdbkrUB22hGTGGYF3gACiEBDChE4+8EdyVO+n+SRrtT33tjvDeDZjMTvX+dTisdI0RvnO
sfgJNmBuBV/pvo7GKIobIJZpgbgB/zCTq9pqqoC1nqvW9sz8JBJYN/PnwqRwxxYzdyNCI9/kaCHz
OvNUjiaS09b8OZ8B3526GyhzSuimCuETcV4doHQkQig+QVmc2gRvW6b2koJ+r7bmhPi9Aikadahn
JqT/nN89t79WMOPJYrOO6RAFVwi3BFY3kaT+tDtPrd8le14kx8JHl+C+rGKJAw3Q1Szhiw1S82e1
i7zZ/LpmpwiUpaWbETdsfMH2viKlRJtdLgaAR5UAspH35As2LITlNVAhY0X8RgaE/YXjdhrEKrB6
yI6EippFdV4dbD1OMilQHfxDmAmeUx6q+wU1wCODeZG9x13P4UFSJFaCfctFHIsUSFosXFXtuL9G
VFn/30g70q8wN+T975MRMgsbk3aYxz3IiYJqomoiRqwv3l9ub+gCMYXnm6KJYH9mXoLF1Z5k1MfK
tFinsTHBvN7SJNj8hSr67QwoFdn9+8qbEUW6ye3fP0n3iNYWbz7XXXts7MouEKAWlSs2D3T/NX5B
n1mkuLsUUQpwjLKlI1Yb1+DTKNuzKi2V/3r1gWWtUuqpCaSV2luUZbZIvNQ6j+XkEB/w3WeQ2V52
UFwAE0U8DnGSMjZyQIpUDYg3V/4EGRyY9wGI/UucIeLiTxtydemB1EC16EkC8Fe0fUyESlY+GiAt
4uNBXMSNGpCfThW7x/d2JAZUovQYpKs2PajmVC0AeqDHebl45MKOecEkRiu2eO72WcgP8KLuGOu+
EC9ng2dQNG5p2PxoKxF2LvE0X0KKWli/uX2nv30Yqf6q7FcN2dEzBQeVZ3fJcl2VXXE4yrAVy6fO
D8/4v4VUBurVy4sJQIhsuq+WaQB13C6Tm5GzL5CZCg095NcoscmKLN8kMsUYMGyhoNhKVtTZpHhb
OqkJW8YTps6jKk79JZBUQ43mKbnDu47wC+sDLOO8gxDGTLuGwYxQgj8miefSFTp01z8fmrMZUnah
lcGh9cLiWApbLPmRdhPtLe17VWJuWM+d4QShH7GQncLzqFc1kKD6XvQM1yyxzZ8jULK2xf2r7EvN
2Tz//UbLA9hkV3MXiCA+MyXPm4V0RYdmGfMUxjsclLSKPfvJZfRmKCci6xsoHXoo7Av0mmjIJfpf
PLnIe9XSvNFr79MRocz+7+RZgsY50hu5K+ld7O2u8zwWY17u6a9DzYlHCA+kdnRsyXdgBRXAts1t
wDJqAt9Xy4oxG3FJwVB0/3f+be+xkAf3F91aPQbCWXpy2cRnzNdN50jW40zTH1h/pcqXgf0SuJGI
7t8O2bt6XHKeb/f+z3AFuDsZ1D0dHk/7g3kaJJk9EJrZZJ1V/pgKaNSZHmQuxmCozgmg9px1/BOW
Q5F7iomZEBq5Ug9GQpEkP8nw+BDwBXovIW2anHweDrw2HCyLonvabHelWKFuDScWzRE5sh0GASmc
b/NGPhSqY/jYbovbBo1fF1CJ/MqvHhskir0mmOLh3zgJrWaomMWLZFQYhu8tAOhY1ZfHxrYDbu2t
xT9eH1GFKfsicD32g6qnsUtik+n41gwVpC0eAOl1bD9Mxyi8B1MssPkTfG9WxZlR8RytkdBtN/Sf
ROsWFLNI9wV2nwkm4nkkgLHrrxLpbeAnTsKOA6DRCrHoz2yOTUL3x6zOVIG9NmULkv4BFNJxdr02
98YpjmdmKDkjYWbdfzqepgOLhX+vvxdR20qEtgScRbAb9YutOU2ZIicp/UI4vzCMjGapLEUCIAGb
lqfUU0SeJ4vZcLdYsP3Pc2e9v5u4X4WuluYoZiMT3d2DFKrAMt3hJF2pR8hV0RJWPmqNdOMHH5o/
uxdASbI8ezAtyoRxNH2QwKh8F/2ttChrwEbmNZDA0p2cPWLFeaSMl2FBxqn37YNab4tiKBJNkeaM
zG5ub1eQ4Vs2a43efLdTA4TKIfBGLrc/xW1o1rKbe+maKK/UuJeYlhMEOxqpjNHDFOnPTKlwc8Oq
rzAPns4hhhw5ODes7L4oLg04KOBpinwiMeF73+7lMnYgEzz9XQuDkwCxhu2j3jxtNivIAThdvF2f
Y0d4d3cgNXiuDlZi6yvNoI97W4Zq5owvNXDuFzj2Q1ZyW7IqSQ+3D36WnxAKFVkslUfwqR0EYmH9
cel03Z+R1RMts3N9N6N/hXFZQ2DgAuOnfBHxxF0lhrGiiNW01UEbSOTAi9vPgglkv5PD8VSnXy2k
fEmMEkjeUVk8AOBQiPgl83jyOAWEf0IDBAv/HB9raiR1fAm3G/gUpsosbwa2BTDDzjZAE71HEC6r
BujfHiVHrFHgvUecTu0Sy3ZI++h9V4VDf7oLit9zKsxsRQccbhmGyk8cSJPUy0FLbedRstE9hLQ8
b/ZEdKwXJKbtwcC6RLSMKpAkG4e1XXxhvPylXiVg1mPwP6jCUh0zskigtaDeDo92LZ0tqLF/+tqI
VFFrVbgESyjKnJIKiMBUDh+pBRQFniiEsYM010LWtzcmszPN4YL4JIqD4lf5IBSW0ZqdQmtlcT6T
HLYvl5g/TMgSKEimJFvSh/T3QcCO2oTG0BlaU8PWOm5o5lJjdKJQXAgdOpUt6RgAI50RselgIWiJ
owps7dfXv1CUc3gm2NVSKu8EFeyyl80vJdWgaCbHtrPXtP1sXLIv7BtQJa6t/Z+DEY/V6nhAdpnD
V0l7rbpZu2Mg8Oml8TTISibOTiWTEeLp3Mwq2W1/mVVk4KHDhegxM9RjFfAtwGR+i1I/Bm0gTxvA
Qb7oRdszi7fkgHyweRUyOVER/w6bqIAV8HAvmevSNS9N55WeOhPhLhO0C0Mih2vLaG3UwIs2tWkA
TYxYiFqOJ5tbhjpg/30eeGqr/pW50zl7NcamrSx5T76Or9xrk0/kDfTPiYtVwdIS3TZoFW/1tse/
N7aRGXBmfhF2HILMl4q2eME87cWps51EPTJXVntJWnct2ouONMlmec5GpQu6wfgPSeK01EolC5Bt
tJ4415V5O/2WzyxYxdKC7zB8OjCY6oEXBXevG5Yq9xPNf+JlVWi/ybtBmVH7cTrnLyp9xP2azmWX
7ws2DB+D95QFxVECPeM5XUee5xNZAvbCYLbqBBs3e4GmJKhAGWhag1ppPtH1MjwYw24YaOBw/Cnz
YydwtBuR2tvfuohcP2k4VloShj/yZXbonyIizvXyEBfmGaEeqTQgQKVNJtr2dta6QGGWIh7XO4KK
Owk9gPFpBMbemT1OGTjn+TJnLAd4EUScYXajuvrPf8y0gfeGQrNwGuSD2eWzi3jT/vbJGMgTEyNz
lABM8KjN8NZafApseLd9o5CBHJKfyO3otT5aBVVZgxgJ0Z+H6FWAIDu0O/pixb6PQOG8cH6YAxyn
nVz0Zt7FHJJ7GKiALHD04N4bz7ORoO2qVfcZJqMYKqIm7yuoD3wANY5STBvM2anIQDZQREamcTle
ESColuoTsKmdBTg2dpSktWIStOHbuRQsBR5LRlfktuoPY4cJF6BcusNSclb8nzZXQ3oE2HLlNkSU
SVwWfhHNwGVHvkJHxZ16NJkHIoEWkK68QVPIx5ZBbSfvOFdbcqNA2ICC9JNaaIjBJ2amRd/TH08C
GumzD6vNJHqSbEDdsoVkHQW/rG+qYXRrHzpaG6HfTCc0JDFUrw7qNYG+G+rDjoZR6up4pvcfa+Pu
F6qp44s6cF0rrpnVCN3SFijPcZSzT+AgWz1OdXpv/mlRtC+5eClf1fOPwNbDjKfL7B2C9lolpsk0
7t1zcwlztP7NPnJogg31XwgurE/Ot+sEPxUJ4Jq/SRa6tqn8RVS9G8Od99G08MKUGO2EZ2tYmPG+
vmjGyClOcvjr+hVDBa8cirAPOngp/IxrJskM+q7L3+3fdYYYqkucjCKtM5/+aLTZdsbKOIP7Pr5z
UgN+wxMQFsqGJ091N+/wiOAxAxci7reyeakmICv79HCyYbUPXZ07zuDxL/wGF2EKe99suQcZD7VW
C3dCzRLzIvReq9tW6lU5UTWPTGfUgvrOmvvc+x9fbFDxcHCloV9QBCOAOZZcEUQL6Zf5oMEgRvCi
hIeQgMcjyH/c8Ps2lj4Xr4JSCaXS9BSINUJnjkiIc37y1fY8JWjXuFj3Oo/6oyZXQQNEq96I2W3R
oTy6hElgMVJj0E+ykOPf+7aVzn6fnqrji0lFY9jwe3E5YI0vGT3Ahvsr41LO8SGfJ6sZ/MF/+WJI
Xrgz4gbRN2s6Ra3hJYcoqLn0EfATkPaeIt+JlYor9c6haAnVhUH4xzcmELAT/DZnnnGJhzP+iwOQ
P1Y+eKdmXcETWlJP3ehzVdBnJN0UEgS0MF709gFFGUgqnJQjT2e+Weh3mFWW7TsqG2XXsE6IbNLB
9s1ujtP2gKcB9dab/CTCFoSAu0mli5fktyVuna+hVq+DUM7hT5eFR0Kj+MeIR9BRyqJtbFIvBaaN
hhJOpprVUsEPa9iofmVQo/rSBtJAWtdjSu+qqpO4dYJvIK6B2Vt/zdWyAfg724ZigsYRD/28xNm8
1L86/ddoA6nR9TNlSLZKP0gFJiKK5bAMJ90lFAclSkT0bWGjGJZhEFXBqK34lI7BygHDosTiwrVW
+r07oeQmbsLTHUGBttDmcnpfocxlc9JQ8psGUkFIUwf18JhD9cLzVPT7dClVg9ZqWlpbMZQtw3fi
TwkhtCwjKyUgNzNKMgcz4KMK0MTYA9O4mcluOiUVtCxcel70SAUIAiFtpzvavd2Sgu7k7QTRP+J5
FlIeXweNC8VzJN7Jb631gRTu2Zs3UpfXaGt0KFyCHaLSm4eRPrYxpZfiKVYBCShkaVCded3Nh8GA
qFcIGlNHxB5r2bZRWfIQl9W40GiKrtJ9DXC75pyboBtuBmI8xj2i3Uqi/28POqEog46EuPQKmpve
guIPP6+NdGWmcDHLA9gWn88xpwQXfAMTr5Y53YSEXlo5jU5677o5GCSUpZDpHf0/60OFTodnIGvm
lGQt5Tc1xnA9SkAZC8d8Eei5Wfx4Ra3geI1Cy5yp6ls/Qmc5gTzZWqOoIUFCE6lghxeIaf6Xk8Wy
GxsBN2b/fWK4p49fw7ni4hZ19jSue8jk2t7lOvQ/4FobrZolm6A+obdTJrUVXGeYMxQvIJOGX56X
2WzEQDHTNeLOruu4KZQtiyxBBk5XDVybHuULEfsG6f/rbYbZOr9tjBegHUYSkwFfljM8ja3M91Lt
LB6uIbjcMWgn1fTGvEVBrH6COQ4Co5FfF5zksfmRhzWLpXrGvboVlJSZurhpqufdpEUmDfupCCUc
tIOMf5g4ohoZ/S1cV+BGg6gqfLCeFZ554zWZDYwhyyAB3beRYhquTtl9MH7b/Seo1zUVIx2DuLwZ
QI3x+tKzSG3iOMilkmZEuwOWfz41Ei7uO6PM16r3xE8wx5le8nYkvd+ronQa+HSIuJcIlFm8YorN
Qb813oT1yvO+GDDxY60maParS5rySpPtuhvQuBdTHmLzME3Lwx7lNWZnckwl7yuntij2Ex2gxrbY
9bf/0Dq3PBGMuzbLFbv6W7quNGUwWf38B61bIYb11oAWXcSQbBLfyGIuzMbGnEAs6bGoC6ic4W7W
ccLZdasXh/3IkzyFw+LQlrSOBmOJbSXsxmjWfOovBhEvNsSBYLYznbBxvOWZtVNyTZeI9ZYjYiF5
kmQn6fjTuKV0SZzo1aPKZtYZs3Y1ZUWsxTvVY+aHQY6K0kDNizgIpo/htpsxprADCZgsvnxdnA4V
qNrgFk8bpnW/tqvJ3aKEG3CVL/40SLtgrXDr3MsHX6opU+Q1mgsFJ9PHK5QVAtVrHhOVKae7thWJ
sd0+o/k0b/+cgkGtV2TSzx79ApVRaKB6+yNoeDEf0+zc6bHnTo8N8bk/Dj8mwvgumJIZc2R0Nsew
on9cZ14U/O+m49jbw1LZ7yNKC8Y1VvnuyYpZOxin30s1s4QQskE7Oc0ByaXiLCKeNGGlgqTDpTBa
MqWmk2IkxsBfSkQFwUUUI8ZRUsuLR/3gP2p9oDGL/6dcgN/b1h9rUBW/LvrKEeEOyyQFslC94Z3b
tZagzc3dHb+zVsurAJnixQ5G7S0Tl563icDfL6laatYmRpR3dDwy0fKnI3A9hYHyEwoiyQ99jiJK
HtGezabKfA8nBifAimbWHtW62Xmsz5bMl6IllkM+r33QO/RtXppW5oFChYCOuore5Vb1/yxtfb+f
KmLCgnJltlpCzq8dXKcuSZd+b6on918DImk2QcWbnBjvtJJ82dl/Q8IzkRe+oBlBf9c465m8lVr3
F9d5SKaOtGpyHTM89OH4qKKemcFGCPL2XZwA4o+LYhLgAXV5QTdEWCZWcJ9csrFCp8CoOe1UXNgH
bvJyT51DAcUqo3wr9d0LvW73pCygyiCWGSbjWQNN0EB77AXqJZCmWzPL9otnxo/19IDRDjUBTs+D
fmZlAFvzbiRDYOJkDTn92khUDToengNbYhfRYrY/pCrDVOzt1evsletvxqf2M5Ik2bkfEwS8bRGs
T+76ialNyMPfTytjZ3wPjFqaMLAn/GEJAeWTtLj3K12Cv/1KXAsNwo2UK52+wZr099HC2e5HxkHy
urEMkOTopbbmt49YmdM3XJh9Yf9bzv5tGV0PzPPJCTfgedQQ5MQeSIxUvaLHuzN7qJRDeU2Qluxe
07GXfrBix81VURI+KOPrRYRD7aAekcWPyZwU/9Xw0a2pOHyBhM0vcXIJ1O3nohBsgcyLJ93bDbWu
wZ7ArX4RFxNYRc6emJrP67EiV3iPtVDdfcxwghlm0/OrFRqNDOB0TsDaiwP/qQSXwdOFPTxaO2CA
EtMRMBavz26mV50DvgrwDCfMWCZFGd3GCrlg+d43CXv/FbwsRkhvtTUizKOH8Tesk/hVdzaHcQXK
1Xqcw/6MX9GCPdU5nWQ0dsR8vAYJjmoWvgkE0s6PeO1454vkN792gMvX4y0DkAjNYGAUELHZa64M
jSzu7dTgC6bmBo36mIWN2OHfmzEGZigT3bTzMCfLiGJ4G/NlisUbDxtBz2l14YVXn3IzFgl3Nbrv
0yyfrFXeB45NRRP3vje/hLjv4M6zybkNopY8d2a4wH06HEscaWlwXW07AjR8Ze4B2Rc/SyrbOaRR
GpaH1IAFTcUvPUZd03XGj2wy3mRryRpYotUgF25MS1OVbAsA9yj62n9jxNu9Dslr0ANE+GfU1VwA
s8MD+F1ZyumywJTYssncP3jOJxtxsyv0gz1MqsvNMDRpsXWTFprsyqlkCAo50ycKXcVxRremvYgU
cBlSgyIrWSsiAZz5mbhP1jf/RMR/GF84omZFictSo6i/9sgYC+DlzTvw7GqIlie3H4qGirkebMhE
miuYruW5JBBfjl1yIAU5CzVbcvwvILGZR3IXN0THkCqkEXsYsj8Gp6trgFMReAQ/bKNPIy8OL54o
aN5TNayqhnUlyPnFp0h8dBZ6u3f3cStb9EXQisCb/6ggTDV7W85qWlOInRPHcAclNpUB4lPrzsgp
oG6zvckOiKa6m5k45ylW780l81rAcNkQxuWW3OqKRET06KVl7hwdlHKfij1Fy211E86CxyWW2CjG
7/PsqeY0+uUm3LJ7mqS2jCKLLi7HeLhy3C3B/kbWbZuVXZvHEWO1bLRELhDUE/6cER2VlDuXzyIS
Drl3FVF5QN0UJCiuOV3KggoMdgSNWFTsdCc/U+jwGmZFVHe3tsGtPak7rvKERSc4X9DTlbRiHGLi
5XeBIa8c7LmkIyTTJiXYvyttAFMPpn5nSLp1KvcEICkvA5taLu+x7A8GmZ1VhfGuHn/RuLFZ4FyW
nGd/OhAHg0VPe8siaTVKg7oG5s4wrYhD02SNV1LTYqaA/34Fsf8rWkNe74BPYYlSNtadVpb0Jx3r
O0XqpBWldDvGYc/TK46NYSMR/5ouHEDUtXS7waQELJLO5PIqoPCWV01Tor0vbwAFvaqXuhJlQCFL
S9l/ohOkxejlU6SXfKV+lBF0kCEE3oUHv9TPYF7mHWTV1TquBFgNkuN7+XPTJ49LlManfswAAjHV
tcObSjUi9Cf4Btf4a/Kjf3Ku5kNmpQn1j6ldgIH/6WE1Pawd84LfyGnxGQ8xeKGTkHz+mS/zNlPV
R45oFHlP7QF6ySVjRxdgjBsu4drXq9VA+qJZH1HUjG7+CUzhZZzoZWenWkKjDGqDtysvPKdQFSSP
eV4rSkHAnX9wIyrBNKvC5QKWrEQYHSKB8P/9Yds/+bidD2TAWh4Tq/hEUZMV+y/NpHXa69zA2ZHH
TZcm3dA+CNlQT8FwdnqM+g0M3DoIpWDV8CefOGASVe752eWOFfuNIovXOGfvLo0QyqEuPgMlTZXu
RCPdZ+Z+GniyW2eaxzGqwtlQ4okmj1Qm1YMQF0NxdWSnjVnpfmgzZZ+74BT99292xPp8jmUwvXU9
LuydOKZL+gTEwWZaeBynlaMbea+9vVuPPMhj8sXxiqVV+XpNEw2Axs1BPXrR8wDyw6ObgBZmbnQB
VTG3KA/4s6cdHcpZZy8fxBQ18ehw/NZIhrelC8TPaKyCRBTbTSc8f3ma7dmcV23MYftyNVNkOZYS
E5yE9TMxQAJeXy0JvEqqD+1boPCuoC8Y6c8vXvCQ1quT3iztOn7C0XRmDF3zOFZzsw8IJOa40Ive
vaaPJ5KUvk33qF+VtS2yOxpyP2UFy9jDZC8BuGCYdFmvrSpZ7Hu6s7JUfJFkeUCLuT9ONead1jhk
Q/IrC0DfhI2eVMC728/8B4CI1Wugd9OIjczF6Rrtv0Xb6lyO9fik+uMq9psct++jVurCDSJrhcAG
tqcjQPGAwIq0xJond9o160NxBODfbjfy4Y8kKCPqKoDpeGkOvASQnVdOLKHdlWWPUPjS2w8MrfAX
nVnfwVN9xyC6JqbaamcYFBZ5nGDJOjjR/c+PJBUpo03f3txmRAplYikedYgleeipyvz253roKEL0
oY8aX46FLNSSnDYKZHyB2VVl7OstoTq+YrJqyPD5oIfvnx4CEXkfYrQRcNSb+qq0Z9CtRzC2eLHZ
6L1RcJSozVmtzc9468CyzvZDkhNaW+V6WHgy2j4WwNIB4ILUsNM//T9XptL6QirWWzUeWPK2nlkC
vi2qrY/0JXX7RnEPnNz4rOQ4Nj/4IMFJyPKiqLYlNBI+izBJul/6KbsSZKQloGvHOB8XnfzB9t3/
vkqJMZKv7D3LuZne+V+0iS5u3bevd10fQkXUFBBbPFI00vnWyIBeWiyoLwNaQKCHoSx1nWefBSXZ
bs9HTKC1Z9AoSX1INv+KgcTapcJguBIHjkz+X4LHbvzPwAnV4RIDRbeW8oXRPD9CkNq4s9PXlFIM
2B2BiR4IPcSSXaMMScxGPPywf2cClop2oTwm0S720dxKo2OwFUOS+tCuPGSDfU5e4kEzvQZabHbR
yBLJNNS9NmG3fPPai3BMGQLQOOr/gabkvlEUJlpsHYobIwbt+nVh6YuhR5IBLDDuiuGXYxCLqSlQ
+0Hejpfk4Jm0pjMZhvjZGOGzuPsaNs8DOg4yCRutNO7bTRKyEdfNZbqGA3GfLxD71b4DVA9JdVFy
tdZbUd8ZtnR8xEPnBU3fykhZRUnAO2DFmlWfQU2X9rvd3P+/LO9xgpS3ci5kt+CjkA+tjAI4TXjL
K7KjakydwcW2JF5o0Dmp4ldMWIBmo70JklQKQz+PRG1V5X9tOBwCwXGFqPERqTE9TklsJHKdq9IW
K4QmOsBec20eKWPtwaW91p2nTOKUgMKK43oNueiw6fPkeu2BYEMt31HNbP4BO1wNVaWoVuCU1HpZ
VdjHBvW3CDCqc01HdH9HUVgNdqa/r/V3RROrMkS8Svu/1Yrr/Pj0tFLBN55Qe8e1iPEm9OVYKtTB
DXQvO64Hxa023Me4kIrcXJrpEPRqTb2C4DiSBvV2TvSTeBynzb7LX6c0XdjDAzylZr8QcqgZ0D6l
IXpa3Qu7RDt/We4tpuiAC5FBaclK2R3H0/fvut0a8gDpP2us8S3mhm3p4lmcBieQyXQixQc+LaUG
bel62kvPNY9G8pMvbidy+cqPNFt3Fnq6ho9rPmaKDBpcZAkf1htj+7IlCnK2U11CZxoZa0IGRNXo
pX0wy9Yy6Bd1I9eo44VuKRbGpUB/kgnY/KijMSSXgg2HYRSD8SXMB4+B5p0kOEgz4NoYfA9cbxR0
gpaCkvsxIPDKT/rr39S+HxdJkmUX2CBLk4xOfT3+mP7jO7JnE8TUHA1CNHSA9vxo4wTOLaHe3m9K
t3worBlFr+TxcQbEsOAxtecGFqGpt4xmE0s9xCx33rSiD6DEKbk27PfIfK4U8mba8ADvqv1jlDo1
RjwkaOqgPzhi4MipYlDdILFLM5qM0xARqWOzedvqr4Bf9a5eZHFOVQPYg2rvIoZXQJFu+hS2oi26
tuo1bqsV0Ie86e8azVcmtZj3KJ7WSmQzJUqfhNThU80RGrJgJnTm1te2BaqfGjHwL7YEtgYpr27R
94BU+0SBSpQ9lPxR0VYD0P+nGmi2yrfpQTg8DN/ZkB0kXeVjKYIbKZJw4njqs1rmzXI5C/pdkJl9
YaDLc9k4Wd4tDWXjfLwKKuEry1X8/lrMp7eDdOJ6HaQ6PMsBK+dI2/3yh8Kldw9aYELhppGu079x
3ezSfM9u5LcUPWXBkC0fn243g/GYFThNTVQyLxZ1lmgI8/Z8Ah3no8cCmhYT9EVMHI4585ZSM1r5
lXQyNItU0TUC/zyFGfK3a4cBh5agAeLJCVlDKituoTnB9DTBwcY6DEA0fbBhslm3X1LvSw8dXIYK
BCeLe9K81xmqmLieopsdHUtpMre7qCAdqjEq4dRIY7H2Kw5dGojernyp+XU3vcOKeZPeBil9Cooz
94LPYsCpwwYfCGVSx/FDUBEScRxT7H9MnZ8j15VQqjbr1c31mSDIWRY0mL48Q6Znk03CWsoj76Pa
nWj6QRdyX5+8yDHqQ8doQ+K/P5UUy5jFrx8KO1OdikkC7EOumtxPkvkmLI+a52CMkwrLak5T1Lkj
Hpx9jkQIIf8FWF9r6n2wJfIeQvEjwnq0SJOaBHVC1yHdH4kdrDtCe90QUeG7UdO4IturrSM9fNW8
Gx0tiQXVBRR2RGUBw8TNfL/4kMbPQbAXB+hqml72TvjxfNXeiEuH/MPseaZizS5IJlCUFf2DGgFA
Cmhi81G7UPMkMPHFKbAjbAUCpdqY62INn2umyKZWcE2swG4NQN8+nZhyrRRopBZeI539g6cVP7eR
VcEApln/SfK5o/4lwUi1AvNHQjl74z++E8vvfy8MpJesmnGyNaDHVbFgC4XspRo2Mr1OuHApVC3n
PRMLxX9nptqlDgmy3srfYRyHAr3jDfDWz1pEJbzeKmXaGC3y5p/02cNCre0pJ1XRm3B7i4h+wVTi
29FykGutzNOLX+mYSFQMXQXJOjQZOlwM+V2Otmj7vrFEUaGOfm+AaQdy8qks/9JqXm1sb7UdSSBD
3fVLP+RR8KowZZujBkn4gRF01kJmOLCzdkJOKmilJMllRe6Pv9FmddWpYxvYfCdeTbLL7HtzJ8Zi
+CD6l7nUQOiax5WeHl+G6l6dg7GUrXdYqDnDOEf8fhFNspTdzAyZEvy5CzpvDBtJF4s6qLDXM85c
ww7EG5idc+Y/vWYfEAnNGqOZbPrbNFy0I2hpUikzoX6c1RehdLhZHNGIkPa8LlMSlmsIsE7+axIa
16k/ngazcdtzHrxGsb6BY33bRTi+JVvwNRrR446hEnREXQ4GmZDpjQKKSL6e9MpNFUEGsB1nCeH+
1X8mBnNOJsCoCl/nkglhIVS8pOOthlwj4/0iN/z+eTkx/Ncf5lPfqN5nxj/9YDcHDWZAv9OsEW9p
RwUpCODK3udEg/n44qXRz09gwUbYS3d68fGLJcVryHtD90K2yoi77l/ETnNNzWnYRAKVTx2M1TZ9
EfQofqeORys9VQRJU8PqHwANgJyMtrqpBbw1MGzTS0oRdtrC/3agS6JEU38/SXVFVQFIuy5naPKH
9HPy2WUfCOTIgV4vlRsEqAVCNoIymdU8DppFy+T12dLFO9tYZ9MNe0IUSfAmPZUBquaYLdH2vv8H
bizjAblQNz2YQaEHFWZNabyNE1Abh4SKajsiqtkNeO/AjEcamDQEaKuk6/2yPQmjkfgRJeRm3aS7
ID1DIrzxBajje1dZp86ajd5+SOuMs4o9ouSHraXOeTR+0Hfwq5JuZGw6oz1sEsd7QxQ8sczmAqob
GQLcOpdUTp2Cip8AsbXK4r3gcMUZ0r5V9zHqy//Jcq+ZbOs+JNSa4/qU8Tycn21mR4gbcN+YMDgL
rTKADc1AKAJQrJt58ImovaI7BYhY+1V/XpI2n/MCTv/RFK1flcNFUDf5+rwaZhPdlB/0EiEALXyE
TVg0V15ev7HJY6e8vMGwyuzssegZOuJOoWbvNhWe7N2XVJoWKtZtHDIDW/lLaBIr2GWE5B8+QkDt
sQQeM/QFoygvkrvIkbioURmhVed9LHMyp1djJy09xYgHJRs6zlqLSrO6NHqsj32D2Aw2UnuxcTyo
XZv3P1kEM23KEm0trUKAYxYaCwCAEGeG/Rj3TkAIP+LMMlVBPX1vLuXjabdunfZIKGEYfjSd/bo/
l8n63zDYCxP7axYWZwev0ozVsbKDL3Cp+fy4+uHwgTAZPffZZKx3EU6jx4eZEc7RqdUZbwKNZyG3
IpLvgu20pi9gUUsRM+Z4usWg1vTLHZ7J3sIK4gLRyTVD0Tb27gWx9FF4zMXDPmfY39S5e+FYiZLf
/EI8oTxK97Xt4TNQI9tp+uFaFk6FegB/5iEND5it0HMiLfI13mHOhlwd6LgPq6aLHQiWaVDbuhlA
Kg5l59icgjVVk7FQ/ZEoAl7daNjn71a303kQVJJ+5Atmpjm9uGuIQG5rDKFcsmeV2+uM/UHvDdcn
iFcDxs5M5bkhWLb4TfnjyZN0kieHrEpPwsy+foo7iXyxB62Y3Z0aCn9TwkkWoXS/H6ibgsvd3QJd
5R4/oHtymC2PQP3x1sq72WQRVzKGEnQ+gsxvDALDqnspXTUX2S556f6lE/AK9f8vl7/tOTwT/kP6
fVae9DbhwaZbTMv6ajdLZ0oJSDXf91CT7O2K9OkmUu5RWa8j2Pow3sVfj+/6T2ul/K4uohUjjftp
L9kYVgof9I7bdC2D5W0n1ynB3dzEeUvLmcBJHdDFx5+w9bC0wpsbJ8z2mHpwi64IxdVi9dqg5bvt
x8ZqaDuM3WOWgh3O0b8BurnN/7qGHrn90XFbhyurXlZrrDq3ffD3jdn6M22TTRQPWBnu0a6CR4dM
pybQz/WghNgiQ3ZTdr+Zj6iqz8j2T5uKnxsDr0xPW+b++Pdhrbi7wvx8bZovj1QGk9wC/y/hHiYR
6aU/+57jrYzUXdM6mvho2mSoFCIu9pjRa5xzxkEl9FeZ990FM+49ZAUXB7c9VVa49+AyqRv/SnQH
+Pa1QWFQoD7kL2A+iclf4wJNjEIKvk37EfkPeWLLBRKNdqlIXpF1Flc5kEYyaF4GYpfGkHBWhVJq
The0E7uRieUJZGnaLsg3PfHjo4HQKEuiS/RUtuJsCLclcnWNGDbJzdgaz90WyKVv3JtvPrDueSuV
UhRA4WhZ82LdyRWcyDCsYw3eB1ARRv5T8zl8nFjxakMCNjrQl58t3F3vN/OTmf2nY0hwkoOBniAp
4ojoRGu2jL8xTOcHSek4llBqdl/hXY5ekgMDwQePzSg4QlnV5JP8wV6I03IAX2TbL0qsLlzmHS1w
GAZ2wMVximHyxyXbS5u3fFITz073Oem4BeJ/OMLNho433I6pykSqoTC+CnP9gOUeejhkEqy9XgA8
spIZz6icoStWx/4UVgmk80psX5IhM9qL2cpGPxCRUGR/eU/aAVoPfF1et/hUW0wQSpkO7Vqve9nG
ydEVoX0c4VrhwGVWwr4pU/aO5/S6o6/5K0g9HRO2ZBTb+aYeb76ryPaRAo2dhD5U5NSUmlXlojrO
zTjbMBLd3KF5+0F1OmhFx2ePcU1h5XLUM/W5PSSxo+fL0HZhLNLE96RBBpgyskUQ8RoGnmKcg7eu
3TXcwJl0U3DSbjm9UyK2LxuDxRH02rPsy5ekZEM7o/7G/RtialNmwXgi+spW6MGds2G4X1PNs+5G
5tzedcauTi26DrV5CP3pqNjmXrOGKLXBm/22WUJBhVjkO5j7dp+SGWuKXZhzkXRMcPCR+6DLMoU3
kkUBHMDdRZS32q8nhCUceaXT4OLA4ULVZs7mkO7cJnUtjmvNC53QHjHZK3c/+eYzq2POXu9cz3l+
1hSeg5WkJ7vl2YBVoErsCeOR9UlAk7jOD79818XO8jj0qQsW7sMFYMTdup4BZjRhVlraimN9VqzA
zoFpn2cBl7LQ/DCnZY5hykvLMKo0GIWNBL7EucMCpbr3gfCrJal+0n3A+x2DGQGKXTIMOc1i7/dl
VkMEJ8Tnk7oMC5hMn/yh1928qQbhHWAARQQ8wguc18sikDZXdqZIMgtgfzLzeb1wMiCCKBTyVMXq
GQ3s9mgoLrtm059DaZNNndR05vxkHFpXWBgveAxt3cLCHYh7NqbGtQ+89HX6RJnTAKkvLfTVGWuG
F8XyCRDZTeDdR8thICQrO0Otr5YY9dO9e/AfmsMq5I75znAljQXpY1or4s1InuHQANDsZywU/Kgk
4h4rBENBxe1BcKyc1fRanLMe04CaY7vmyGM7/ktmixyZBecCU3fQhW0tga/4R0kNIVoyqodbbwCp
qnqM58uu3f9L0teHGG9toR9XZ9tVDJmOJjgoc7MRDO65c8bvyHZSawQmxrJbTkNQGoBz6hTEi5gE
f4ZbLWCslYUzPG0quBfamA7CdHjT7oYgN+SRMtaroWJ6qfmBZBdI6PMgfj1xV6yKFwkak++ZZHPs
KDXc9JPCz3oR7vfP3Tqucx0z2Qb/IqV8/LOEYetH8oUdc4NsljxPjPNa5AH59Js2uezPMTZQFyPd
44wpaZlf9v5F5lZH8gI8gwf04D3Pv9xFL2Uq7hVZ+DF2wc5ZT+BkCDrb7t3yTvmwUvNdfwtd9dIR
N/j0jswaEBrMnNlQ3+hel9oRF0vVydlrf+B8ef+ixrAznSsnHlQ3vrNLzwym/RD2eyfejVjnI+i/
+T1Z1S/VwhOnX4b+MPgOecTGyRax5FRtfPfrQsmTFQ26LfwECnAAwM4MF2oQzp2WifEH/TBOTw4s
dGoh+BQUIdf6flbnSD9lc/QuVzRc/Flf7aHWcWJt3pTs2zCV+X2Oy7JNEzagXqIWu2JtzgJrIxPI
9ir/n/OsTGP8GDD8QmbVJTaFRvGwDsOhHoy8GP4v9eHifTcqT7aBjaGjPRSBebKlqGyrZBefPEcB
Gp8zd+Icgo7NZRLe5M9/ApZ0NHEoePXgxKdAyjnxJnFVacXayHUUaKLpY5nczs9YdNTL9yCow8Uy
1jgByTr8YmyWnzC8UMr6xQT6M9qfJrG6/e2mJQhFsoGl5K794YE8x0apWWQcRKjSbgAaojFClKCv
YrBA04vD8+5VMMlIcA2WeIvppBVHxjiwU8J/bbbSpBvrPVXrddhVcL/lA5tFQT2UOY4WtKNSkHVP
8V6QKyOicVB4SyQqN1rWPrFR+n2T84hG31B0JNHIc0Z2DT7jMhyN4ksTWCybi5IkhmYR5fFOfPWK
UNagKW5JJ/bYqpz4Q9dXupB0wXUOuz+gLN+C0X3zYhZfzjSxLajCLYyRTJeCGEyO1PxvDS0/ofro
AqZEOLpWXEif8mF0XWMkipuzLNhIIRyBXj3zZCR11fWgA4BglRSj3LD4QzrUtBGiq3MKxU79YCNH
+pA5qHYnB5VeiMxTM2n2rJEJDV74Qr91nqpfH+FfPMATQXQjZvlTL5dRj0l3DaCV9b1fp5TpxXWx
hDN8ndxhS5I6jt9aPbjJsAJrnx05raXa9HxEdQdyoqfsCxmUujdTvnAoHJPbUxz7IqWsiwfYnzeq
Pb+Ua4SgOf9GvUPlXp88gXM9Q0DvlpnPkwjWYKEYQ2EuW4rOkV49r3kWpY3R1dnNYtb4oZBhbjwk
gQOCiXGkUhsLjeMa93eTJhW06GPaFEr39KS3HSpSJDb25GuhXTbqLMyGt7VDlXHhNQa0fHuPv4Qo
opmvF2BcOS7ylHD0r8TJpMvFdtnEflJQNB2NZijN6tKf4mHLqr46XlQXfAKzNfyWtheQ7NjnGx/6
umyZFtJ3LVNLD19uaNda+RN05VNQdYhDsO4IJeCvweCXXwJfxL+0gbrgteab89n1B4JFZDrGCwhF
4QZIQhF156SgOCgWx55ZXwIkXZuBxTfVRpxwrTHAajQfeJkr1r4VsJH8QKHDyuNwRn/w+lcZfSyH
viDzxxrkoyUGXGPeX6JW1ZDKuj9Q+sO1iFO3N+ryS1RdJ5WSjr67RGQfjHic/4z3PyLYiaXG1PsQ
s5OeqRD9KlLOqeppjQAwkwBz0Ko8jiyAtMh4UhRqz+7bfqm5DNS09WH1iUsA47+3U5oX6RD91ey1
AQTjWgLFBVkoQA/OzxiK7ZIDuH8xHnA7VsUpnkHghuMxbmyQg9x25atojqQByykRyCxTsvzPu6Sb
6wq85edEL7FknomQ6DJ/sL1CG/ejY3OvDHHKPe903q1YLX35gCpFFcKZsjlESVFed7bkhAC5ch96
Ht1Frlrvvs425z/hFeBUcO83mfU+x9XlBPm7powPit4LRhZXSn2HON5GlrHYiMQS4/QQeTk5Vu2q
c6euARfd6u8bMhckIrIqVH/8B+06VmiWODnqzzBaW4KoTRR87zes62wWn5EF3FCeRKgqmUPqkEQ+
LEOxtSpkYSUIld1q83VRl+CARgVTy3kHhrYuB0J5GhPzU8FOrgQIifQuAuEJE7eLeQ8OGNdJraAR
PCsdHEBknx9gINie05G3VQEL8gz/SQuAxPH0aagAarrDXKnu0R3TtkOZAyd7kntsy8Kuy3ciBC8l
MeZNLqGykWvOa34A71nvPYgd8KbWvqGo87tYfKewBF7B5swMF5bJsHolZ/8zELJLKoikn6nbTAIg
JaUI1IyeFC8oEYcq2lVGklK/SHz8giHEfDneQ1IEf1WiDE61C8z+sxcYc9dysHRtjUOmkjwMBYe4
++U4bNqmru8kC1XUIgBVhVbeSt5kiiHkytSzbwU5pQRNl2+D+O+4yZ6lFrInsinhWgLKVecnFkXU
TSR75Tf8juRbLoyjnwk++j18vOPkTF5Cd0jDbq7JifuH07jgbPlvN9OS0hHCGVZO0BRuk8/5spOU
Thyi7WqrQeluEnG+2uWjRb6hgwaFYDWSGqK15SIiBUozjHyEPaTz6eDqbffNB2Tm10hU0ETTNjRT
g7mPoYAX6zyM2xmp+k4jwEO2pFldq6SReFJYzk430y8Ux+QwGb4RsN5JP51hSaXWiGDa1uA204PG
6+YjXSkseC4q19HGAb3XWQt7UAr9vXvPO60aTYRAjGsWmQ8PvbNqR2kqZqpqEehaEz8Py1Aa4zIV
8cWmHU7by77Rzd/glxFu72GrRJaGzqv533boyRr0nJCkBhoPIlJ1Mb/tRs24pnph50jvo+qYoGkV
UpEKa0mN7RsDRxJQSmXQDUpvg21IBcLjQ/v/7CkTHDcpVZVM0qDYCWn+EcOJG3TlFlgKT5/8EVtJ
uM/QL5ZumpYn6EvDDyQbOe1YJgW41vgjG9lywi/T4LRRLQEpnUnMeC3rqvM27r/WM4YoWKRqpEjB
t1CJwttr7wL85OlS0fmgKRgu35rw2ccTI1pjRW25IxXEk7QOqA8Pm+EFbo+th9VF8fwL+4IntgSB
PSs2cs+uUhOJOrIBCdSJk3jtlg7LSn3aRRkitvxo499F6hOk13jUOARgd+K+Sj5Y9P5T2UqIWD20
WYMychrpPY5iirw2R+uTkZ67zARF42cQPiMzB/d2IrWGxH5yobgHxR5yk7yVni8C9h1uejDkFcwq
rZGM2vCkB732My37VbVi3vsqKD+UkWcJxWYcK4/PNAHDlyVmkOre2DAG8KDFIDXmabQKfkI1rFB0
A8+dYvX0ykwSnYYSmmpxg8I56pWmrlfj5YTPpZXy1QRrbaNZlQLd9YOJqY0GXV7Thfs5NtWuSJa9
YAcX1Plhlq5tbzPcFnuAHRrybNm7aRLSWIoLOLWgyWI9N9e12Svz5uT6HUohETEqko7k6ngyoQ0Z
wDOHDO2+6gRloU5HWh9uQM/F9H0PCK0OZGi8zWD4wzDkCmJFIBCEqpei2JBjTd9fvwocB0PmMs++
+smU68JlZ1QT1JDLBhIrdZa1GABj0uyOPaJyFPbA+fBSTyQd3goZBgOPu1sO3KUgJv8/eZZReDJn
r7p/DaRQmviDCqTUFYU5QX3bVZvOKc/6hV//rVabd1ofr9ULv1wijXcE2Ss0WgaUJp4rfKTmfAnS
Sk8dcg8QMypI8yt3gShzb+VE0+FGD7Ka6nddqfqGC8ZhaZDCg2wMK6xBIApnRgKuP2b2qqs7GStP
/Cfz3gABQBinWx2RDSbyD8GNMeWoChoo6angALB+QGiNfG/i5OAec/njEqCauO539uLN8AgM9e+Y
oOc6Wx+Mkt6d+oIm6FFdVIGxmVWu4hNguNfwpn+hVLjiuPxIY7reFdHsAo0k4f8PGYL4wDNW6Loo
0tzvgN5DiE06j0Lrb33q3KWmGeF1aayWV/k37ffd9hIjTR9PoiQAlnXz0Iu8WhyfO9YBN26sxPaR
97eZZlMLeT54sdaTE4kt7+9GVbg0GmYEZezYqPwBz+DIYs61MUtmxrMJOYrjRA5iKAdT0d7Il76S
PTlmHnnN0G/uILCZrzPrDw0Rf4L8yKA4qoaeNK5LfyJdlpdwqVA0EIEWh2lMotevYWEccrULq/Ez
b/ACX7cHPR6uWBTHAfxtTvMw7WNX81lVggw+bNBk5y9v7XGxsKe5AIlpXBdlKzNWztSZWs/o9oyn
nScBMa8cackAFbhUQnzKI/Nc9mvbnKRQFA1iFwXFz7aWdjkiShDibns+DTui09gtHnqJDDAMtN8D
v2RAIuEkuKodhUQ2l8tRLLejyjkGbFU3UdoVqP5UL6sm6wG4XTlCTYd3NQT1nE3zfauXIBRVfQEs
Mw3N2mDuUyFN5V8JgwBU2RKyh/xzGUsBbcNeM06MPdwr2+VGjYg86a4ImdJ2o47beDAahgkyBiqS
FkosN30iKcLJvsIvmUhI4DqD4VcWQfocxy1qxVpfYOofHPwDO1i2qTUNKjA3n5Hc0yKQaaiRgFNX
6zZ7ppDP9sfk7Pi6cFNQhC+tUx6wGYJcpl7o10+NTEti3iZBLxLCHDfLhDTaNa/c11G/4ptoE1NY
cTea6rM31r3xcPFu7t/pujfoDYhAJfjvDtFS5TjHUQL/X0L0kJZtQbVMLW7iKKzkk9PSs/1UOy4P
LqhTd7O/mytH+QdhnmefuOvOw4DSYcvGRtnDzIe90EUO/ta0hrtAjep5w4ZE7V+/VKNvISQgrzma
ZM5UgAq8HAbxI0BcUNrsNWtibX/pymhvbJSu6Ov6UQH7jqf2UDq5YtM4YAEFXRfJF2uamwixdLsq
SME838HDBHOwYl84AFx0OEz1CGUATOfzWsdQSA5pB18FW50dMInJ1b1lEQgBM2u/yVWXt4Dqvbv6
RtjtcOlFf7uMJp/C+hpc+lP48MuuQWMlXQggBxPrImAZJCYIbwlDjLCuh/MEXdX0OD4etWgh5N+C
6k6hPGabPWaPyAGaFv2XInpXhSGxxI3u9e+DO/kH5rEU3mlt6e7r0ofKG+Ys0RgP/ml3pZUC5eqK
zAHXxKBX4IN04MgDdj8OrTQolHxmiJlzPNrr9PMFPzukGP7+5jk2rmPw6x4//lQLHDd2D+NfJae4
pWcfaAWn4G8LLECtabFFVMtw9+i6xR1z7ZCb+JuWk1+V8Q10D6iqmC+NoKy48Da41uMVuO5FBzlk
z4zPu9yyepa9monrNLRelOLPSNqdV60WmV/XY0Vlsv485UcfgkMn8U6I6AVbK+4fATXL7dyMB+Hb
Aij06E5VYeV+Ru7Ojlai8w4hPe22iEBLbzpYh2BKDAlv8qeE1MJKUzAbEoehDwix3Z8Sij52A8VN
p1sbyxDvNmEZkVfZpvvuXM3ANKZhg+gj1hJ+TWVZMZyCOjEpCt6jJTzN82+7K6UR8n6DRaRBguLn
Fu2a9/eTZzfgcnbYtB3pCrM7ukXKbwOC3mbCqx1dvP1w7+ynkuErLb9erenfjjzlRIN5WX2y6mzS
unSmvRTB+3FE8407efzLgdTJnc6Owp2T8VnmUXqnHLt3wOG5iUyKUS/tqb6e6n1t/nYfD0DloAPg
qNC/rQtjH0w4/EskjH1XGKvoOTkxW6084ajH1hNrMT+ECC6mQBomyp9i+fq7oPPTPQW8dcyoFEuH
aTh3e7VkATcqMA605kHVz1FCrKJc9qnx9fCs1ifRPLH7BeTT37blhPdwZuoCSTS8WFhF0x/5kGcR
3pGxrjN4ZKjiIfq5pnLqnur71PkQP+ux+fBdEex7bFVTvcYs0PQohH+dwNIabQ2ucMDDmXdyKjrh
MGJmd9znpU8Sh/xBvY/KKBOxASNYQVAp77uOaNXr6rF1mpr20LxY6wKr/wKit2aJ+Z8IufPKYolr
Lv+x2eKjB7+2ZTbN0xzfJh3EUGMfCmRSnav27Ugk8SUVB1fNLMandHQkLf4CUcZqX4FFZvDPGOSC
BwrYhn+PXhT8UysTGjozuA0HLpUu+rBWcDQWmes3eljj/p/U2ovAWQyK8OSjPoha5cksvhuXM/fb
nXQdCpsbFazwLC53ZW0dV8VibMHcUC953gRAtCur7+NCqEJVY4S0YTcNy5fhW6FqTFKKNRWlH3ej
reomH7Z6ZLlIOCRIoXOnrqWqcmu6wV+2mI5PSzD2WoUBYfuqxwpJ3vVz1ovk/RI3MqrveqmCTWVC
vmp7+nzMf9sL4KpH60Mlj4t9btroP8lmSPoYJSHFMDbwGNe5Aydh3sd+/vPM9K15Z1uLS9PTiipD
LGcgIlGSSZ0ZHbGXRYuiuMmsY4/7K8RP5HTVAw8KLKKAgLIvniEnGfGQmo/4ExD28/glj/8NgrEC
2Ydl64KON6B3g9HYMKBdS/xBRrTejo85S9WEqcmYsIQmgShVNKYA2oTpimQ5t8diSYKfE0btKD/D
7opAodVaxlPxNgWos/aV30PvGhTwxpVEVZVHAmPLIrv81fWxwRNht5l8GkmJbL1vQh7Pw85Qk+xr
yzgvVI9ZZx9l7eX6jRz0vKeLx0Hue76C1TSlwdrOS+zZ/J6nqB+0zUZNz65ynqR2kD2mDy/Fm/TM
h+wfiF094XSdvAxPUTo9dcVIcVhx/PCRWpXx76xsXRhUnm1r8VXqO8t9SZCq2DiiF8L3rzuPsNCq
rslF6Qq60e5/cEaoMro6ycrKzwRmJfB0D/pRGCetF9SMURNM0J/mdHBHOKs0jb+GUp1lMWgToSnB
NveKKV8xJoncCsEQgPT6aDDFSmTm3PwZsWUbJRIDahz1IZVxPl/FyHIjgw9TkoFjEym9HVE5d3wj
YpMH+bPZDrirJGmawI5T3BYBS916IxqhyIGnArR349PbfwbxHtgkCdZSwySssVSF2ovmI16lskeT
8ApvWn8rWdaJfoR4/qDm6QV1jQlRaJ0OpyfovSUqalN3+i3v7mRzId0E2tMxW1k5ysloBn3x558a
68voq1VnU7/p9gvUZbqZfB7dvmH9DlpRLtTg1xKpm6ndApxbQDFVromyV/RcceH6+inUKsPxTsih
Tv3WuhjvOEJ90fqaHpiCxOmwyNRYVvJXtjX32e70r4L+xhZFIVtZmQfYMPB6gvwxMrEizM3pYi4g
QcLfxelW3mi5N6YQPiHM1mb5nyfx2Xl/JHLuxXXiC3Epy0PhnXoG25jj6hjlWTOlLRsHJvHM0m4J
QRx4FM9np780Jt6KtkUxb8L9o4cA3JIPjTJJR2MJeJubC1ucRlORJMvT10xUsIDl9+RDjAN8CZqU
B7EK2l1p2td8/PDFQXkXB2wFYnkYrQB8ZFS+MOWi2M+7Ai1BtCcgzFm844vfr939u+Ng5YbCA253
VfGSRz213tVl3nMeCPOA8kUxRE4YwZHFUtaNBZzuy9rkJymoHscBkx/FDLlIHeFZ+9VHXvrtePkZ
wS5ekm7/6h5da5XmDth7SC1KOHh1Ltas2ElDVKTaDZbfD4Xb4ZdpOcHT88t99ltf810K9sG7ce51
6JRsNBVD0ZZWXQBKo00TXmJVlvaJmsLp7y2mwCZKuSuuDzZPHz/ZS0oUB4h7c8r2vuIvgXriLaff
jj/moM37AoAhHdDpFv3s+PQH4OWMKrRs02DizbJ3VtcY5tchjYSoG1PlcTWSj6yGocJ3B6bcKqln
xFxK12H4hj4tnDMDJp8K0FR5tV8Ogze39V7fnolhhPwkyVTrDcMrU4yYruGBTWPonITAoeWt5YYP
tyrnL6ioudjEEW8sMJDFpBDKplKrBVJ0+Ubwq2in3ZygpXQZRDcgH4yetaOE4lB+bgstBTmsIfNz
W4/qwRUyQLGkaQ67GBQCYxrVQ0b55pGprEZfUPoJMBO2f7TcOKd3/I9CeHS99jUvzf8/6FtzTQsr
l4X/8fRzCf8sekdJV0yFqW7w3ikD2CzamsTSosv558SfkjZ2bizc2GY736ruodNxief5qqs5cnva
KiximILAMYswkWWVRGzMq/mFoipNng5FwvG+/75dd6YulZ+fSOiCI6GX65YzASFgQWBY02Vaknvt
5reNB2W4cR44ZGU5srXAySIrwkTrvI09IXj+t+0uQ18yU0AVGGLUam60WdGV2HK2NtgKQp+RZvhy
Ufsayc1ZG7CH1En+Ks3m5Pixd/G24Kg42MdL67NHwIZaaSphun3T5Wg6WSc9VevKEb+959e8CuLf
EuUa0m/EtNeKqQsjlqV4TSUx2VZOq5mVkC/E+y3SNOPYFUkE8MbwIgGdz++KrgGH3XsyiRRU/FW1
VE/PbSWduEnythXJCX4yvRWnTK3tvWWFTB5BIdHcV9IPjcZ/rg3lUJOg7L0BUA44Vn3tgh88GGVb
0K7+jrcSeiLNEVZsHoiJKfWFoRP1quioYmXJ2CPoriHy9r4VOzfyHwBDpuTPZPG1Fnd1XFeU/bXo
ZwU4BFijh+mhjbvO2ceLFVAzCA5BmxPLThTXAQvd2ZXvGxM8HWMwq8w/oAOfNImJryYhKeDRAlfM
NMIqJoDNevA3nlMkRHrKnXE9x6F2PpagLQG+IjpJkoxe04DQw0Ec51tPqt3nGdHb8McmTGNfgJvd
Yrt06BkjEOYvOHCELpHCR7D/D4tNKYsUe7VvS1oE/qqnTG0X43WgZtzI7AzoJzhu8Jhc8neoB10O
mojVuccl7zjJ5KzlzbFnvZQUctTOAJjdaNUIXZLRboTlas0He889hKotOQq3eE4DQRK+bghauKpI
hk7T4Ja/EHb0DiIgMaQF+3JOLZb0xMubPCjtfpi+7LC8NFSfV50y6Sg8fR+PMTbdhtIHr9ReHj8c
c4jrmFmUcgn0FF15o7rsTaogqTRlPErjCAjNFSOBIQzQfPuzNec1dV5XUqB0DVEY2XZUOJikEIqs
xHJk9oSYlGuExWTNI1UWJSLc1tsVnzoUmcJjf9m1E0abpAY9ZlYjuiD6zgbKULgQd3xnh/3sXzaY
+86GfuceypWlPjgzkzqqxdslIPbRDNhcsy9pjTJ7spOE+ZRIlvNcjNJEx2yx4ZcPGT7iUKO+dpI3
7BEYUOsl5JRrvvZEUZH+07R3bJCdP8TQUbwLFCsLaoalQ2ZJZJQAWjBWKRtUSFf73JIxsLZUwvyb
l+w0D7R+2t8fzEVLKToOTMDomhras317ggU+cNo5Zr0lhKuaHydIR40U8ywr2LkYep+CJx4afum7
uSPg84bBlk+lOTH80ce7OMdUlIaGP5k06vHJS/OtGuhd5tom+uizJvwt5wOK4N9gyyEgnSufOUcS
027aSdTt5DUrbdgHCcWNG4okhIOkPAb4p8s0+W+hnRoByfuSMxJIhHEgJmvohgYRm7J+Xsakgi2M
YaIpW/EtyxokZgwYewft2bOzPSdRgs9cEGH9pAKPjwSw3A3ZYATAb2XA+rCjdZEodWh1i8UUNzmI
oQl37kKnpeuS0N1DsQ7N8Pk6vkWnvTGPEBtEnpFr4Hd3gF3ip2F0IuQqLAFMSKFPGsFASydPnBU8
Fwgqtfm7EHnJuPFmGpURGpITFkomoc6Hc0BJ9yLE3x1XDojZogXx70IL9NTzhB+fX1L8/XziDunQ
Z+GKxKbizz3dalt/+DM/Fo4tj37mrsoBJkyVsheh9qucDmIqLlaBxXVyUx4NjVDcaSEoBSrmudem
5Rhmrsi7luB0XCY7YL+xZq3U2n6Sige9xltLLS8yIlAENIXXB/RH4H+lY4eO+4bKh7SVEjiUIzwC
VL6Fe8/7MuSsmygdldy6euJsB5vNIu+1MOQSqLZoUyEMDRk1l/0cz8jdhxXH16qFBInRnu1U/kk1
AScCw/ol7ZcZ3lUyDjH79IH1H7hQwv/z9I5tJsMTC0JXFkbGHDTfhBgfm1JBfCTRxZfaw/YtCVm7
iSPq1P0T5rX0k4ZFsbLyUwv8dlLMDdvftDWzSjxEb3nyp3GXSD7t5438JQnWyz91v2diN3be6i5T
4LqkiRl/IMVl7GINabKc3GhCu1VxtGCdfaKSebyPdpt69NwElSmjrTe/Np+2uVOpWh2XkZMyw0T6
20xgpoNVDt8ZS3E7Ds3WDiivqm3rrUH4l9xppxt3sEBjiBZYSQmFjRxuoljP6Xvxy18Q4rX63P6y
LKmXYikg803XZxltB9AYcxc/LHrrqsFkMG6bX08EVfFupsIiYXPopef8wuup8rVlORbN0zQztu8D
8WJkJcBCkUW7ezQbLhGMoFpdScYhMt2UkGWZDd5KtrPEM0+zOrGxPRY0crmgtU4FSo8emNulSXhR
Bv2IVFF2qbLescM3ULdWM45IWLtCsfnhhcpYsc3GVX1ePBJrrKpr4NEqOg05BUNLCc7SRSGqXCLs
2K11iEOm6snom6Xuxl1NyYW/xjBOGFOUxklJeN5WiQrzmxxdqdqafTT7BhYAuzsIbpwGLm9BbLDg
hvldaeBKGC8Q9rQIanW4lFT9zLqbaFdEUVl9JrJNPr8uvHkqMoN6fBy8DS62+/uW5opPlnEZ+L7A
97SI1yeOa1yOQDBYQ/zFX5Z8qUMj1NrKtq7B3Me7o2Fi0RZPtETL0sw5Rz4EnBbnazcIhGVYFK57
YSdCreeybYyfIUkIKW+doyP+l+JX8uaK0tuXeksUJh3t0gt7tj09ZygF3fVT0n5xP9XarLlllew4
aZfMsdr/opOujvbgEZGsoTBrCYGd6mqqAAro/97uptZMhyayPDdtabxn/OUC4Idfye4WYyvI+uJa
s5DMDWEZExk0doKnWLm1wpInQemUfJyNBevKUe8r00FQ4z3EwApYaRdkujgP4UM4Amm/LtNGN6W1
voYSUefpwjWJeuqeX2tGEJVx8zz2D10hbgHG0z7L2OtA5rb9B6kW7qun9F2uAAz53tjBw0+ZCTf4
uorDvmY1UmzMIJSV1CgfsgrqGzD6umxb1JJgC4p1LfK9lihIEsFWqUQfwCX0iA91PsH1nI99h5Nl
SS1hA4Gm2rrj2iCUK0FRVXoA3/BE/UB7iN1+ttgVV8L/2tUVdCXRG4UTxAQF4T0VLq29Z+ZESnQM
PdcgotYfRw7q08t4tesQuentv3Pykk4bJUsqMMWbVK69SlsaEQPJfrf0AT9skHdao+qH6cwYZYXZ
QWXTZpnj8XxlNj7wURaq3W/SaSnQ1wyL7W9qAjRxSZV6moxH14UbHK27wwHMw485dyB8SS7ZMugY
JereWFqgYSwml9SgtvxlisWXrfs74eXvF0QGE1B2+t3dN+g1aKNL6/fKeMmP/GUzauzykLVT7pnf
aZSiEC0aPZned54x5cilqhvNI4KWCP2buF4S5RnkRkeIQ6v1pBqBxmv72qMhSo7xoiCZSFyq0itH
J9e2D6RNlULNkMjXYkdW0YvIhBvL6GnZxO94tRIYzeBv5mPjacnddwLkJTNdxkHcfHrdOHInsc3+
3ZzJmC+ttW0fe7EnXDwAw6yMG/fSDZ67JhJ7uh1gBSgPhu5teaBr71+2cCX6NBJZdqVEh6rqVSjk
HQ49DKFjJUPD9n9VxpmzWUdrI4PUvGhw/QCddJs1smmIIVlQ1puZx1cCFrwc4SKotELd2cHK5hyK
8ujhFXoDyx6V/6iPGc5HcjxqkLhguJrYNop8nwlh5cgx3F3q3AoTYVrOZ2AM7I6KR4oRQXSPMuYZ
saIf//g41j3MMMRPRqZ2FVfkPTlCa2H4bgqXBE4rYIc5QWSsc19IwU5TGx2jdg/3utA5kIo2qOlO
ZpvZ1TWQXoxs4vknIicLSLSajA6cVDpyo5E2ITptKy563jnrvGw0In13n5TC1PqiPuzsst4EAbVy
o17a+srVfkruf9VnAk9OP4xCjreUljkhHDu05bdJ+EdVLu0bGb/rj3TiPMNKN/bCDlM3Bq4fsugO
e2aRav5GCknfFLa8vEn1FYBAGb/FTsGtflsaMSgO9QVR/9nMMD2MNO7crHzMjqoxb/sw8Q/GnqFm
vBFkFHcKpqJOSI+IS5gv6nyYbLhhHSAK43Z6H+XGjfLoAjxPphG6ALq4OX3cejKhK2njLTTakDyn
S3UJ9GsNK13sGaPVhFDfsluixxSfmyPlVyn1z3gnUwSODj8vwOrQydcR/UkSxmr0IMoCngouzWUJ
X9VMPML7n0W2X1sKceS4Sp/7CnYWWzjMCDpTaVjOlJ/SkieWiJ5pfyO18bRsQk5tuIJ12M8/aF2P
qgTmvHtM5aB0Dtv7ax6Xua489UmljM+fDJhMrg2OiItwQl0dsDV/Tfzl3F5B6z7t/FIX+LwKmoyc
hyOxKKCQTmhM5yfJf8nqaADsgWas3Ge5DHAeUB5HbSDozot/bU9yCetJE3UAaxT5YoU6tcmbVwyK
nY9aq6v5C7W/gadDCrGgpSnA33ojZtACgRAMIKFJInNhB4yKOYpsA/mCXCJCFqN9RyiZ8F7fhVYw
x2UbZhN+statOBm//MNJgVGSxAPDLatLke2r1CQvS0tN5CXftK0pGvdvGVyOjFR3GZ5wQSSe2BlD
XDn3ghNjwRn/2WSbpUe0ITORDcKSR5VLnrq/9xKgZOo+yk1bICkRuuupsPTr26CnlvwWg0CgB+Uh
TEbkutuQZEAwylYwDZYcaWyBksOBuC8eZzcLBxfuJqX71qZLbT8PrQ495wToV5b/6JiYvnnsBziQ
Pmpd3OR9uFiFti2FJzpcDMGKmaExLxSt9yLv/GRp4WANYHkuLCRCR1cf0kPRapbAVX1XVilqZitp
7+CyO9I9czhDGlph2KnUwQqpUAx4v4kiMLuJim76dKCkBKOBNvsd09GQM3nmVajU4EW609e0h+x+
QLyJAONxCzE7SN04rB2N3xfcI0jFesmT3hH8bJ193E5CL1RIXMHG0Zk8DgG1YCCUQd57Vv6mv7/y
aKH7RGQ28qeInNHYlXcj23zHeQyTnjFiXo4rWInB1B7YimWdl+vpQQTU/yZ0a5XZPvOGrI2mmKIG
hO7NkFryZm2PfFddN7btOJD3qq3RWTu/SxUTyfMmRVaD9UDTNoxft18cM56Q0Mec9qXzwY7GQXrj
Kin6PTIrmDr8FbmbzagrfSVbDEAEsgiQhXWVzQXKdJdDdFEGGrOEZ7uNxJloJqS6ASUUWkOl2tYW
lp9u1VGN2ZXBI8jo4g+JKwbfNk3+leMfZj+lj6wKIp3P9EHYmvi509AI0+hJ4ffB6tVYKohwRZUj
fgs1PxpPaBc4uWvBaAiFuEYXBH+C1pV+tz3DmWhXNjiW4MzEu7SmJ/NO8ew0MPjLdwXjcCxJ21IL
sKrQrmSfDZKPPLPT9N/yVPHhnrqkPWBM1f5YXDVRE3AuvOVKH9CTT6wNRNAirhn3iRMDCDJe7W54
+CypZaKS764gpq/BiYNY2w33fkjjNtS36gJhJCNQupMWKQa16/Ap9ysNdqG2AdOtquWluWujN7wA
bAviJt4jSqX6IjrNiE2K0WqmzWvpCkgNuVrSV5t7HUb4T6TG75yTR57zs3WwBBzooh40QgVHvCJF
8e1Ro/Fvql5QqmTbzDmnB6hPMkEFVVjuU89hIHcETiVFlcyc+Dd80uG8suGuqLQGQeYEMXQce+Rq
gIEPShA+Soxb9ssW0AXZ747YOpact+fxwLZAP3+vphpol8PtCR7W+dUjVbQM0oeNMtlTkr7Akxhd
HAoGrnlycVSvcTPqF8ECo3SPlpMWBch1DdzwrFN2T0nrt0Xph+JPbNeDRwOLLeDIgX2+QHfATlzH
W8hZi2yublTHriKX6q59k4oZI24Z7M6gioAIVmAn7/AheRop03PTHAYgInSrcVpicO15lxSOPfiG
f/afcnoiAIrJvvYA0bxSmhMe2LhZXToa3sdU9dR6d04Do1cNEE0gtvCOJiTLt0ezVGpD+7vtBXus
N8SM/t8+qIjU9SuC8SOi8iqI3RclPHnuLdG+o2mnktgpMCCwygFnP4uatP2UxKFH5Gx0vqPR3sa5
sfvODsztq0Tdkzvqi0kTTyXes8utYI6w9mmZeDFkYuRh8SkH87ll14MZ/c/Oa/423FSuRITd78Qm
vaItOTs+uiiYF7StNa3JV8vqlX6kvO9qhVHEB7pjqW7mhgTMdX2ezW9+0irDisMDJvkkvNxxSYaZ
o4BJZ0DI+deawj+IHAEdahzyS7/ocZu1/wsPm+j1rdFTlCV1QuDWyv/75GXRyJIyLFfjmdjtYrwa
CuRQYru47Ro8iVeuDfHDrIsx0+sfsRhZFg3m48r3CPq09trHPgaed9mOLPRgPTOYx3btOZx7aO/6
avpTbAmsJjbPHEY2Hz1Af6KCCUa3MyEQVAZUQjARc3FgoUW21nTwn8CPNEnRvkNrIKm3GPyRXFgG
llDLd43y839iF85j4m5HMm4DbhHPNPJWACza2xHrhahOsNzPqZja2ZlSP+q3dD5rxhrPUG8rg6J7
oJovhAyFtltpkmd1Bk5xEGpcb4oqDnd0N7bFcwjfiCCBzqs3S4fHySyowPtsBiVHd8MiVwVqPr7B
fx/DqFnO63FzN/BDcpY1/z3cm7OW6NEWxXDiLeQr9accPXdVtmpNh8ODKlMSpuSpcfK73F/uK+Rg
86NVP5ySjA0c7gxrobTAdTVsSMUY1OcoVu9sfMV96nH6OX3KpqXk9FZ426B2P6fn9/t21sMOdH16
OSI8KWb9gWeM1+xYNchQh9Qa1coCFpct1HQSMEbmvantvirBVbNPCq38YhhYyD2oSfCJVoraFLeG
J9AwH/21P/pz8tlBVuo5+Jmb3Yb2evNQKHqVe1V+L6j3F4a6DrlTONKbFYuMiBx0HvTOKJ6n+LDK
ssiYRuRsS2RRtzUvNSgJGeLuJST7piRzQbWFic1edaQJavh5m26CNU/ON3LtMVS0vX7jdguBurnG
wky5UcnsU96mfd7mDqcfp/v6UZpYPfr1RAxqCU+2/Vj1phRyLbl41E8PogtinwdGnLZDrcU1vcna
0iXo5yIitTikVvaiQ/gqHGNkl4PvrqEdhwv7SjTZKVqRkZWALKTd3RBaS0I/pv85YuMxnonZxj6w
UodsfeqUsa9wITH6C7fUhFEw4uTwJTL5nRi8E610KtXgc2+T4ZCgejwk6ZGR250jHdKJHvLbWBul
moxZjZ67CQr+bhprjGwwrMiY8gaGSiSdpNpCO9QMqVuQjlB5p5RqCh3XE2FpO6Cf/iMCGdJOf2Bm
lTWUytgUMOJ9TQnVJaoh0E9XFXjZoFKOOP+nFBiN47123CDHSwA3NdxW72Z/C6oNyVTb4++TH228
VjIqT7MLCD/77MbUr3vwnmAVWGawoPsyHgQi3m7/KGONOT+1E9AQBzOCwojIK6sy8cNnyt/KIA6Y
lCv3ojtkbpfFWJc6P6/ZWYirHXTjN6UjfpR2S5zJjlaY9ESCcHClSC9yttUFADT25MTVYsM22cq2
TMXjh4y0g0SFtfyy1R2ij8BWjHbHeNk8LVbb+vp541rIzgn3S1gw1mA+WDtjZ4GZfnI81IxdpyX2
KgGHFfw2Acp0NDBdFMPODljtZXFaLoaY/+mlekOre35D3ZvnZLx18I0vOgXvkr8252dRea/0Sjlu
imzUgGh7FFLKCEayuvXM2E7amLYtpEAhnR1D+t+T/6guU/GXKMN6H2SQ2MMxYRkRe9Y3yNQO+Lmi
sU3ZqaMircdKQ9QeoZqQoBnx1z5RIn+UvXuTTA2luwnqhBXKKvS8iwCRURoUSlZ/q2ifA/g/L52N
1NXRPpS4zukrd+FuP2uDQ74pG9+4vlZw+aMpEq0wwPI65pp2UB+Qmq5MjZVrEQ1GSUqn4Y/kO8pg
oXvXPb96LoEkJlbp+L/1J4mq+0zgCiqIJkySpewIpUZryYN0zTCfprB4gyh2y7brSLnIrGHL4ajg
OcCKS6m5g1Bj5VgCJ04oCrM3rO2iE7DyAH5CEULfYuF0iaraUKNmoyBoWKQbrBNmBaGAXlzW179B
O9bpyS2UoLkdSuT818ez6nToiqKhjI/kJS8D4eNVkj3ggGQd1p+WXh4nK4vdTKpSbw+gtz6JEUpi
OBaa+wyJErcbP45QdU3qi97ks46GPt/KfE2XmDotq75ZxUkAQKVTWUjDeTi35KvNvJED8d7+lfhT
w6Mn+d54h2HzNN0hOK8g8L7fbH4UPXbVuHax5GN4r2J38T7KdRTAh5iu58bK1AhqXVJ3jGSzZUqS
oBlqd69BUi5iOQu3iKABkY3+aUQ5scs5uUEEpR57m9Ok2Bpbs0yKW5rfNpvATOWL+KOgfzaPAtI1
RnmhDS8GiC2I0Rx1pZc+spp2dmdltkTcwVnndkEpDbRnG88oGlL1oCZcmkpoKZ9D96iDVcLuQIpc
7J4Q7ixBHmR7Tei/wyETNNwgEVLEJaPoJakyuF8h1TlMLV1biBZi/e6qPNeiLCi3XMHL0ehgrnFy
Cd0sXIWtgDbfDDmAtIzwdtkA7uiXYp7zifI5eroPtxMKYqq2bpngqIRL+FXyuZ/W1rY1IUH+JnZ/
Ze6E6t4SUjT6f6f+YVKeIJcq40l5JtnWBZ6LPtu1lAJJ2kD4YKBHEh0xqiVNnpwbI1SSVrrT1Sak
roffB5+vMvQc7L+B1Li6LT0EiKY43YSYEzk/HA1/Yx6eEP+lMCCYp4gr1ap+0pm5SIc6zm3H2WfW
IOqNuDJRHEwnX0CIxrTeMpfmlTdQ5XI6tRTM0em6IQlLpT0FDxU/kHipRzKuKJhuHUnxB6ZMV0oK
wPXPk/sGzbQC/6VXARvtVKmDS51bjZTVmzc3GVEYAbnn7SfmRm4yJSgOkL+YpYaTykww8NPXdnv5
WvbC2BjwqM8baRQI6OnERlBmAvoF4knvIMZ0qgnOqtD07AFzX6/mYr3MVNc6dOZHPtfIkC6n3mS3
0JrWw9LPZys6s5Y0yasFO0iwT8zLyvBgtR3MUs8s3Qu7mtQIimUjNkpcxIUz1ZynjPZcHNrp5Wyk
bXoZVp2BFeRQxfqeXLAm2vlb+0dq7XxsLwyj2X0VMsUufkUNxdDxEeW3+bC1jqUjxZFI5V99ZgLw
7juisAfH22/bcNhf6Yd7NZNBkZ/369DhTtFT7rOz2pfXzGAoxi8Cf/+F3taiYEp371ODQgT0ynfm
A2n1WsbhPtRytC4/4y0KrVlJaHLU/Wbgh82Q9kf/AILZjVvqRMBxKjHnepbZ74xtFmmOmT9Qwr9N
Yc10pcuHR5qVT7t5JSfe5Ms9Eh9imiyI49UiPVVwo2oaUSw/cPAgTgde1QmIDKFjIOjBPKYGNneI
Mc5iQd9eXQLdUw8ghOXVy3blfk0i8jkS4/deB/Onl0rFktDzcgNY3SjT3momAMyx1RAO95LVQrgC
b7gvt4oHwrzMgkBM55j1IwNeXt8XpI396BbmIiCs3CAVgDdldl/OkhuuSts3UfF/5ZrVf8VF7/Kl
sI+yyXXbUxLrDAoXJGYmc+R1NH9DPkVLRReCuXg54Na2yg0wyJqWZ6z2PDifC+edjyxLMP/hFmyo
kvTA3iNLdPrURJ68k9cBhnckuprUercM40OTyWK83zsIQDjL8KNE8j8WiHssay5MTbvxwCq5no5h
t/1C2vYwOsJ3c5F47jSTNzZeKd8U9RfNmL12Rb6lFFY4/hTJdTYrlUtGg8KQWJZ+wzismO6oGWPY
yrwrsBnsEusd+JbQKCsuZ37k09e1OTep40nMwMq160/FEqdslhxZUQcJ2Ju/oZOWXyEXbFe1Xxh5
i5TOf+hJxqJI71FVxr9h5pSjiuPtelwaiCX8xoUGBoD0ddnGMiJKUqtNpFttT7VdAK1rWfB0S47x
XEeM3raHoYrvK9hDMxlv0UVFA/XqF0e/YQrw2tV8V4eUCtdcc6zgr58wlITAcKMvasr3menenTNj
9bBqSBIODUflFt/UwPBbFSWp6DHin7VMnxNa+wqCXkGDZCYcPhj+dV/c8kisX7bznIk90cg3dhpH
z7P9V0YyBe0Vi+kQqgJ0wGRmdrV6SQd3ROe1kIuPf4up8u60Pm35Kk6FeIbPmUHeEG7fjg5tk3Nr
oV7shV3b47+XdellmHxn9UA75L/UHaDHSga092Q9hf71ku2OmXJ2TfOlRvzJGI43eiQHkcSQ+Miw
IOM2dqQ1GiNLTvqXCqGPrWBykTIZ/lwpGBcuD4OKwPZwFdjjlWPnPRPvRvi5PQIFuJjfm90pQ+MU
0aeIPAz/HSn+lFqkjsYwdWpq1yuvajgUOXOfAe+rD4RuDYSWRcZ2vTJU90HGmaFFa+Objv0aec4U
Me7rOQUG+zr0UyRPLEzOk1BleYBOiHfS5qbDCfjHBMqFGD9buQYQLg1xua/CiF2MeDU0/uA1VmKy
wzcNBr13v2MdbaLUx7TgCbO/GeUONZ2Yw3gmnl01h0zh1CzAc6DJB80tjffnSS6i2VdwP7lkwTcB
PYfNMswN9gko+sUrYbrmXpAxW1CNHZ9KHX7AtZmX/yC4NlGX/1jJjEXgxsVhh2Q0GHOg76A81v6z
CHsZhQMj29eYD0RsYkLG1PEVq6EUoUdrJp2v33mAFPT5mCCSCL+wdvNU40Mvl7GCYcowwAPLMGnm
7gMpB3WuZ03FyLAe3BnjLnj0JhVpy7+MBEpJSKGaiAoZZK6UpYp9lcXjGE8hRtRpKpT//vLZ+dLk
3xqIuI00K75Lu6DTacmNReRUqMCTAkOTJwyEorYxCb0Xd/OdhEBRt3H/jXvQaa2y1VulMKUu7cH4
x5dAs8Js5dDmqWrRcICvE7nTZPWktjSRBr7B3T6M+lYE93ecmRUwEkXFRxDDw494NK4su5kGLndN
b1MMtPyR8ObOnNaG3Jog4We5pG6WE2RjB+UEwljIPJYJGGo/ox+3vofGUlMylRvVv+EwCd18XeSK
nXC/TQDFKJOYQWSNhZEUcZdCPvBEYXFvjFf3erm1VbckqDQn9vNa9vMsPRC1qcj8TrOZtGRLJxpW
PJB7gmg+gbxCUp/ytfEJO/dNpVMhVULTN3VgTRp500eVv6n9DmcFLb78xZNyE0aMgdW5cGlgF5JJ
t3jnaFbUmenJd1PiSAJeu+0Zc3ZAk1r2AKjxkawqBu4miVdXl0ioko0peILk0G+Yn7Di7qs3GT7L
z7rUQny96rnPGhxO7ioF0vzxfYAtjVXrF70kndNvkdMCMdG1Vh5s5+JaCnB8N1xDZVijHKuD7FMU
hcqgDmaYYAVjZ572jcKt9v3E1z0uRR9FmFJSlY0nrli/sLvIRUoZunjhHIJQWVGqTHis3HvbCxh1
QAg1+v83uP0b2hHBxTqWh6lBF363dcWySlMVktE56AAtUKHllgvF5aJobmC56EE4zHfySRTFzpYn
nxrKp4n6VoDIOxK+RcLEmchlInQvE0kdT/osp7sevq7gyj2S8KNc0Qg591kBOAyqlrA2yFHTNOxz
ZO41V24vD4VT54ulzkqjUZNTQ4uRNntQ7WDFtGD+mXHeNw+14bsBUyv04rEXJoHyxUnBhBfXaGRo
+Ql8cKJ0zulE7na1G+MDK1AfjMv9k4BMY1yvNFHDxFS5966Rcra+TbdpCEc+UgpSSqU2Y39aCHEu
2/lhdKjxhLsr5JsuMZ3AfKo2fV16Q+HCni/LYNRrX6z2nRdXnk9TdLoATV0XRbl3pofKnMD2+ctH
nEdUP8Dw38MVFoMCT0M7O7FbZ2zX/bgzmLRu5OvODda9Y6GWGuskXvrbKyP5LpE4f7hREbH41vrb
ZVttO/cJG8j3UKf+gOzlF1cmv1G4BTFOJyAkktRVn/aOFi/75kOsMsCd2undeAD/hkCMKzUPV1uU
szxFIKlnSSJ29Q7ByxPOj7UGf8jL4pZCRv5xY+tQ2RsUfNoKNBx9DuMPdMN4T7FXD9DHzXvgHv47
UankulqYthb5JJaV+Cb8LZjCClrTwpdYgQFcvPf1u9e2BHy5ZgyIkxF91XTIN6FJGCTKgXjjv5dh
XOm+kREqJ42rDdowQtRhk24Y1JIdFqWPgBksw1NWNwZEK/Wczz0b/XWpwSOt8dMcEZUMyw755lNQ
gJvnEYr9qXjbABXV/KF1u4ACrLh1RhZsHlvOecH866gyNFEMhRP97j5WboV6aRG+/OToLGMhQg6O
FFrTia1YcyHxmpk/RLTI7TkM6sbd48KdqU9ICfYlfJmRDCq87/NIhBEAJW6LlASJO4pT6M1Vb3ke
2SoXz7kp3dhi3dLiVcU7sG6pxJh0WTduvAGP9UH/w1XOQsRpm5mz6/nRBTfNJJLB1xXB3gxj6Gji
KMhq8sD3gMz12xTRAs45SnYFFn2GvIqmOjCHL1Ikl22ZrNGN8wdJ/O8LWlnaOIvUVQ7L2XbEIcoi
qoQTqu9/8aoarWLHYMYlXRptXkTsX5Vr79FZ/4q9U5z58prH76fGypu/yAC5pHy0oqu69SgAod3c
0j3u0qdqD99r0EcjK46McZ1bwK4V8x9ssLHefnJkC0RavAu/qTp7IoKM3BQEEQCKpJ125zDQ0ezH
Xhjb06FnaCJTls+Pw8xLBgYPKEigks7CSbQzxgTW1x9JesUbxgVDegjkIX9D2+NQe6BUYFFAl6Fc
Ai8mq9gLPh2WEem0nLj1s+ZvlzsQL0VS81gfebDEnZnEwpN2LZYurWQaUrgI/bFbg3YxFgI85Jzj
7wjum67jB0CO5pg9vXIH+OD24OrjC8sw2H6KTTHOnWDp/is9zL79U1+SYVmS6UlGbA2AMjf74Lx1
jQVZ5oQ78vIfVAcXP5sW3rDj6Zj/zvmOaE69d623Fd5tnAODYDHIhn8I7Eh8afbnPkjIop2ONS4f
Jrx7RYIGQxpjnGj+lEyWVCewzaZ9p6HYJFoxCbqw5JXfgRydyouu06ki4qPQTmLWCLFUtdY/MiYI
BPYUFY8QeXHqdePG8ejFJxJEyFOXKI6pRJgld4XHHpAbSqaGB21+ZWjXRSWO1IjyQkty2Bh0Pnsf
XSmZvLGQsvP9tu+4IvXXr8GWMzJZr5dMDPNyU3A7R2Wyt1svG3ZRGBrBqQAPaf6oV8YYMsRav5JS
f0v/SeaKTN/InekFLy49tlFAwYfLqyv+2/n7+7bJpiqm5FnIaJeboc4vuv1cGBSlol7r8JWAJzBF
MmezYfSmFlemLMfeWZCAVKlcoerXiOMCN80zKKWYfOXkI/okiiq8NH/vIp7tkQkCKMOxzf8HdZpr
i3vrSqbmSILSEhA/cSYhGf/jSsYv7boI0PB7J/1Cxa7iytNjRKy4szRuuFPem6dKtWxDF+ht6X4D
2dDIAHPI1/P7mWvYw3MxqBwnhamyUPGGtP+GOS1LGTmQL/NJDmqBQeKjveFTnM62+ocLM0sTxyma
8t25czPyHeuoKZxjgp4UvtGSV0OfAYSACCVidICO3eSQ7LKx+VNBjuQfECcAPn6GbdCEynMgYd59
j3+xkEch+OGQai1oU0KO6oP5Eo67+6dqLknXRNHbYCXL3Ubc8LGQ8xJrT7jsC+WmfWQkKXYl1ZkY
s53gDpS4mXCgVhDFBc2myLDSOshACO3/cbdRnNZTGVANy7mCovDll1qTjZksVFQTkjVQUTJtJ51X
b0FrgJZ/xtl8jRD/oikY2jAu93HfRoWhNOkHgFa+u14+GqenVIIkU2Q6inArNZK1coxKoPdsfIyQ
ZShogow4cqjVYmypZCU8o63KqLPtl5bcXrbP9RQt0RfTf/zd+4GNL1+ElU9vyW3Wka6okvpg3gNw
6wmcBuM+JNijZApKj0whwBGVfyhwug5ytc5hXIbwpiiKigrf+UaXsSYcCXliYbiK6Q/TDp0MzxfW
5RlqIJi6Ky3B9Kl93ecgoHLWtlh2v5EE9+Zmxm94hut57OpWpELcaCoujC/6eFudolSNY2F+PnKk
t4VbBTe3TAD/jW8IC7+EGJyL7g7cixPIPNQFNFtCOg+nX0MOGoQLsbCZE2VSfCTYTVWpPXOa9KIJ
iznDeNb4obCX1mEf3F3MuAbaQn3yQtrxW4qOqzmRs1A5jVwbMMebPOHUYA2S1tw1p+WPpw49mkkc
ab5CRtvyDTOO7fywZIotg6Lpto93lkBNa6ECHcy91ulVxTP+opu9Ie0qwoiU6SDa632XbqJv3hAh
yo538tRS0bqOa4W8jMPf7NT4/wPcZ6X/972sGBlZx1NGv3VToBGtQBaceTZ5zRHLn0U8ca66CxdN
KYO/aNA1+LvcwdqkJqMTSYHMnUPSvqLYqTckSmb8K2dLqq5rek1rRJX/HGgiytUTBeEUMK/+Hzxt
Iz8miVSqFsUjy0wjRcQIU4LmP5GNB7pAVLe9AFxKJE2ObP1RDqszFRTP4tpmTGnNnQ17oHcWw/vC
hA3L+V7hkNL313q73Brz7VUpGEdaY1fyRVg2muNIGjGeRGCiEUX/V6qyhJMAwzbPL5jW3TdbKueQ
iviPxfcbvXBDoJwIPqHIsZIXC9q+CrcO/gsSgbgQXtex6Wja4y8O+SV8cwHnaxHZetFsczeN926i
ZB7oPv1UGSFk8p1257GhdcMGA9ANBBhnm8cr8oCXHdrWC/HVjoBJgoVyx7RSdVadoR2WcZSzUpUN
1LAkOqWKIVjIUfl9j6ANvj4IrpdvOnZJuMu34RnHhv2B0dT/OiC26lJc+eTs2GGKgFNCjXrO72PI
LHx6Nlz+xsRwHrexVm0gSRmYb0yROy25Gst8pAsQdczZVhC/ff6Z4BUNOmFQud5Spvzmf2r7uqmi
f1rOqq3PPWe8uoE6L8aChncJUxn5R6Ny7pxvW7Zc5z7V1C2TRNXXUvqmM7Sle3Gg2EHZcwGEdG6L
6CLw9RmQVY8o0ZxT0x4I27FvxtrhQSHIngu+49itXDKVfIFJAV7Pv2QGaAhHef5QmHKb9+8HpEuC
GELZAOipVQQtwHrueKreqtAoR8/K3JPBXf2ST/M8EKfQEl/WSI4ZazqWniqPEDhR+4FloluOd4EY
dw7Hh4T99mZcYtrKWtXbP00vMP3q8nGiGpXzAVxPMpU9idksaKG0HV70tpvXlnUq6XHGF35VX1aN
AjEUOVWLLBe8ngHqtAaAQ2twdmuFHbz0QCVBS2RcaiFYuEPuNO7xIuC4j5ZOtsP4Z7uMZigqnPIe
gZjdAX067uQjH6EHZHQ3S2Ci41+7y+IxplAECk/E9rsF3OZkIuJI5GTstD8tWG+DqTpi8sMKHu5D
G87da4j45xecjyZqSXq8qL5bfAvdBz6v+DY5sSScPkI2o6vySEfRNBWzCW0u5fWyxwsuLhDvGy5B
kWAk618k42DH1lIBLrZjn+1A2s4rh1r9KVVqr5P/wGY7RDoGFnDWC3St+WlFGuDA+E3Z4nqMUxYJ
UnRY/pMAy6nzFn3C+isww9JmOHmsUEEkEsPJNIy8Aiu89U5KCBZVHEdChcxS1VAcwJfBqshgVO68
S7Fwpxv1Ea4fGkfBLy+McatYDiPSYwJXi8+7V3girkt552CN2s0azvs6gz2vTfLpXy8wUevGQyu3
RizLGT/S38alQZOzaN+UmQleCJ3kNzmDoMf8lLAUnEUB+alR0aqOkEfIc2Ty7HzalaC/H5LsbhPD
cSh/45K0uvdTdCKTz8ylyW58urPq4Y8GJXyYvlW0ga/rgd+F+CLHx/mIoD5m9lMNYHKQplDP0KPu
GrcM6VCxwdXkPb1owjff+b/xEaAa+BS4XW86n2Fdu/7ObNrjeS6eR0Qh6GsBLyFtln8nSgso9zLH
J+yqBq+HZQphyLrXwRZrNkHultc+81X+ViBJVM2fkZ6wCgji76C7F7+NRTqzkDLRKOaMs/0z96b/
mScmLW9GpnMjifnQFI/OoMD7ATHrjh7pblwWz++FFfzlrs2d3ACsDIDpN7zK2du/lbodL4FcTooW
6n6f/EEwV3qcwt8OW99lWtTQB8MAFrL546t3QOmI7ukkMIiayjv5vDczcRDBCvoTbqVWl8NpcxRT
Lb1AM9yUxkyBS+cqJ2Rw1LGGXe4Lffd4JENTdpkmBaNAOBl4qsAKW/vGKMyhMo3XSU8NmAAvmPFJ
cwdQbxZK+lg3+jgr7rWLEiTAi1CGTYG/td6usFga7UVjsMw8Dl6+HqKeG18QRF5OOOZBrcAF+f6n
QYt1Uf3OA+iJSn/MHjUy9uh+8ttcl3FghTppCouj5Vf4xjVyhD3xkpAClghPTbMFm+B6aygf+w97
UV8Ck22N48e6wILyh/9OOi3EzhwKWv382CvzgK3sTN5EmO2T0TzgC6pjY4Rk3156gk3w7jQjTQ52
BEL6MDsKjYb96CLk55j8s2u6uCF4X17eAczypmC1WVo0o+kk1IwKkIr9F5E46IrUEr3/SjK6oTmy
qiPTMCo4C3VF3sk449kN7h4S8KXwgZRov8wqHeK9AosYfoRbNr5hkCjZUoFe/m58k0Ys+mKyBvMI
fEHK1fHX+Dv4b+Bk9t4dmqtuUcW+o0hM1iwJdVkZ4IC25e1bWW4wULlE7W2JXagY+A6tSpvLu0Lf
boytU+V+aVWSckOXG/sNYRhilEQyHZmr60c+OtfaOaGw1kHxb1mk2LJYNWHphKikxc0dru+57eXW
K6bkdAfEz9N9D7G+Pjrti8Rv4KojnMaa+iMKQ9RBi8Gc/x87wQJElbwDsvmd2v1YA1ArBQqwzWWG
Omqyj1lgeMPQA0NRB3xNiduEOvIabH+dPmb5Dq7rcssz2+VTbQl2TgqjEnW5uMKHyqvqj9/NNsni
flfFmd+cadOT5BQ2EgNkOCS1IVxZLNuydCE6F2RSCYqSD1DjaC/Cy6QWGsZ25vF/IfMNsiasCAmt
xe7ysAi8XOrHtQ0ckwXJqYhxRdqtq26hoEBirHNzG2MAw00v/OM+7urHbh1uzqFsFc7wfLY6PHWk
G67r2Yuix9kjG1/Ml4BeaElfMugYlnrcqna3ep4wbnmrxZcp7Z3djB+zKK5IwcSumk1yS/bEMtL6
59bUnJqXwZVFQQrTAL8nGcVPKAOp7kWUYSHDVc+/OL+zrJKTVUvaMvBeIcopMr2sk3udaObqqJCc
7DFgKDcsBA+d+spZMi27ZFEqbppPejH5LecQ1VWs2bpJ3ciJ4JCM7A/5foKMBRJQqFa5u+Oyy8bv
Mt3YcM/6vVc96cuex1PdRAxHNSpW8j+vWEWzR8DYjU8gW5qkpJ1DFZkXqGNAhXnIk2YHahLSSDuc
2BlAIMqWClNHLIGroNam445Bexxx5tezKXPkVARQMlIDk/BK7wTAWENND6CKhgl6e+7d/jA8dqOF
gnIMXG/ECwt9Nsmg0qpztVqcujNUbQ2bq5OToVlPDbRG4CvaCOFa5kNDNFl2iWhrby0F/SLvOzmt
jJe2MiUEuBl15p3bi3TibmNw/k4FanZm07HOmLyQY0mpFQxz6tfDk5q2fcjXMGBDRcuhJMHtiRrb
w18QSI8Sz6lVNr6O6XP+pRIJ/q7oCXHEU/JrC4f0jSgwLeqaa/RVPUq7xem6eb5Lta/0+fimLJKa
afwK0rxK8yaaWRffcWSbKpZmwRjVcivXairP2PUGd7xskZXBiBv6w7AGPWkCpog46pL1VauSV0ng
ms9NEH1htkLDaOdOy1Gj+R/ug+rLZhtllONEyQIPFIgnBHih0UlSHd8/gtkzpymeXbOX3ZRXlp9v
6uwVFs8gk4sGcMYJhzwp+SCFsbERnlMOoXtUxULBA/jY7PunOz9B8MAfA796bEBT3WYvMqHeeqmE
VYjl8HOLKWq0aTRw10kos17XR5CBKhqeUGwto6Dbka/c3Opm+ZacGNk/bGAflbT5S+7E2wevbQNZ
KfJVfS+0rNrcRWish2PdMLhJr+utiJc/x8KLKhvJ6EvIaesaDoY/qYE0zufCm08fRm2bDOJJWijJ
NMUaflhNSQJ1QlFyU7VR1iw7/W7uAoF4cPyY/RJb0EB7R1FRj20Z2Zj/b6XpeCoRtQdXD8BpSgnZ
6968uDzYEw5WZ0VQWjwJj5ISSG2KWTMoIrY1uIYAbI/WpGn7dp5EzH7DYvfmclM3wjJ7leRVoeS0
7uj/ioCSN7PccywwyzCnXKe3HzE/ic6zfDslPWjC58+5FWSHTNauspFIfjDebxT/4NXO0cqFoC3C
hceWRmBsp/mfypXG6ubtS0IfPnovP/Pmy2uQpbfzX1HCyxiTKjJnw0NuijaVBdhkyX5cpjFPXdQM
vx1yC3jIpxgCBMs8wAZ5z8zdK33O9D1ooMpmQcXwmcVJ4nfad6i6mo2r+jcOlVCMe1New/Mk6Drd
bBTkhRuSRi4qg5+6lTeZXeDtmRU+VZb4C3Lf4PpxRz85ShuSYBRv1s5UQlgy0j0ZgIBthEdlGz5/
OztCu3dLmb7BdFXRM5/t/wTtCx3vA2+dWG7m25Ua9ht4nNxl2yW1BOxwfUCdjvXTuDFE6rUgbc0r
Hcg0kr5xpN9SeTccEvXjiHTSmnKECo4MRqlm70PIwWlU2zeL78VfWiowKTpqZc5HMr+ZqBVFQQ+c
6Qea1jR66LVpiDd3L//OrZcjexS+CzokUFonu9za1Y8MH6k4kYTONY4eeBGdCEOQXsrQKNtQBI6W
0O34AW1yjV0rRfk3dVz5+mTgkTyPmWiePaJjDxLeKGzks14rJLju8crKNOqEXOrkw5xgZHGyWjXw
47QqL5RkWouZAlNxakTzVRmxA4o/e9bqdW9QDiu05krH3wYPsF0I4aTF3uBGpnwr1NdhyILXmZf+
LQuVBNE2GOhyg8YNyQHRhg6JUX/v7S5ZBZCXv8o+YDqI59CJhhroZWRbrwGvbDvgOwJyshzArTzE
f4MvpKfwDK/0jmYepem72cXw1WGq9SwE6V0FC7O+K+9NhAgYgo3FULwhY02xyBk8iPO/C4ByKvWm
M3yJLap3BUAhmQIyZFTdaaQoHNoD92kwXFdr6p2X5vJAv4K9cmdxvYrVbmaLodVEIeWhOJVoR5r+
s1WT/6jwYgTC3q+AhVLphLsb83LEKVuTJQx+RRVEYow96+Qq73FppZnQVUHGolSBqJcVhTL4noAd
PSLyPCBy2ISrxjn/DF+RXsHTPAb2d+59ci+639aAUyfvqcdevkMAG6/rnbTmS9V0RDdz1Pt88tbU
fiICC48KhJmTAytA0vp1FuTdtvXyjg5mREW9lnLpWB3DvFS5mnMOCE3COW9pmng5YBQ5TTzBR7KS
PWGhkJXwiBTlESdJQRIjhIcG+IyGn87z46lN4OKZBzixceCeEBI6AGKcAVyCgytI0gppYxH92mMN
DTBZeqfiSTzU+2gASF7ksxBzNtnFMzNf+07IxewuNFepBSSC2OK8UYFBz7mf3OeX+czPUaCacwou
4z92NYEj443VZrkFOQhPCyQjTkraXNOqXQTrFR5MrRQoS5M8mwUHu5KcegjQGzxLunkF8Ah0H3gx
MAMSMJfi/XOk5SzARYJ2ZgCnNiwmnDqMuHgd3G1EwVmALJYCmFRLap+G2nT7zzWoE+HndMGqockM
kSIJOaQF9lU7vU1tyrja0g4m6vNRCRF/Ol+wzDXmthriRV4Ia1/fkpv2xDn7p1liwfH3uUqawNgO
xf4JFED1L38jbx+xD3I8yZIH24K9cE+qpg3M26bFGD01EH+vkRnRZArcKvi2bes7bMlp52V9Ad77
coLmM+584UYDDos+DeBDYZqrJTQegGGSZTMUa+bR70/xKyX8HCu1fX2SH1+ifni8gjrMjboBBc9G
mHd+Ihea/mfqSbPuYqNLz1pEt6W09qL/WcaVHFOGcqjnAjz1M25k07r+utgxIZOGirr8lmMyvQRd
/WKc5JQfLaiTClLzNai1C3716sPyWbZ9Oc0OoAUkihfhvB/3h0QAhI6prfaiRcu17jQSSRrohdxM
r4Rr2B+AeZsFRMhsJB/pbc6HInONnTSGQ01PVGmU2kr6V2hG1veq+UfrqEZTR/E0Na8Kp06mb9Ps
RUmNuoWWI2pC51Ky1OmNe2uiIEIKWJ9dg4l+JN0Qc7VeU2OfTvV9HNtDeb8Fz+3Bj1kTH+h2owru
wWJsAqPmyE85YgkroddQlMJm/rw79BiU2GgGo7mQ6ClYQftHnO906JF7CGaN/RbelfYkDKN/6tUC
IgJd3dSW8te+hLQcYQ8DDPZNT9ROyZ37hzm2BbN8JCUFQGwFmsWLoRpd6uRFH8WFbRkj1QjUBl73
cOtnbraeOO/otYX2FqpivwgmzJDxghnuCBmj190c8urghsWpikkD+p2rDIZMQvQOvPZ00Kr3trRf
PzOA2PH2+pApvNgtUdZbWDyQPnmvukXArRVrOr2b2ee/MDaFZtQWs6QhkFa2YWieDe9DzY9umtXU
gDYW4FYuY2yf9Edg41fvRGK+f65WA2wdO6x62dtG1weK67TIkqbKy1fnDqUjLGsNJnWnpnQ7w9n0
aAuUjmgmWt6PvYTk873E26p5kp9q8BfNfl1I6dHYDDg88Xet9OwameqdbYEuzPLZkRGXLuO5zyvS
5qMNQ0wvY5Q4jTjn2BNbhQR7UIATBn/i2b+G2WQ3eCY3S4y62rGZBnYTh5h2uQa09/27OrUw7lSI
I0bWkP52rPLh5keWCqQU4ZvCflcoHUZouYM47zWfLKzqwtSpuPNi9isPycQNObWbdBRzeejyMqJ5
2LVGjxURcuSmRZFPrSmflByZ9ZT2eJn+g63injTmFNeJ9tBwBzNT2a646Us8QPXMRjHJGCSfDs5Z
c9xFxDd4m3und0NTMMH7Rr/fHR8+2vsDkfW4bsMG5M/f5aL6aaSacIggxi7bjiIcbVyc3dIMDXeO
ZLBTr1mSQ/n//mbKsVw5gqyKFn4bl9+jdsSckAzmPUckUsT51VJBeZmh6gdVzod8ai/n5FmmRzZn
4gXHEpN2KkBoxLrvPRJIdnV/hGNcAby9oUhD2ynmxpcrPC6amWxyAtSnTzaem4FlD7U6rdEJc6UL
/wsO3hzrkKURlofO9b1kzFsFx0rUL4dpBTLfXvqCz8wFDbVwxYjTykV1rLj4F6s9Rp76ut18oCRT
R1lul1feBdZjJU2Ux+tw/vnbscNW/zT8KviYW89llLZF9MK4DTdUjr4pWKXt4poti6gTWo5weFHh
c5W1jlvgPEghklpn3vVlSpXoXE9stWkM+9zykuHFjgw29RzfXfDkYBprubjymsWZwBmnBhwmu3mz
z0HdJP7bRtG+jTCGXNKSP5brKhQyLVEWhJ5Dsbl1Sp+ksruQuW7fP7dMhD2lkhftxZJk10ffdbmB
qK8P8PC3xKYek1PDjWIfiHax/Belinh0+6X9TZJDF8iq1SJHDS2Lfr8MTb6YU8PMiRkTVEd4WIV+
dMDRsztlxmoJ4SRNTpHfuk+sJtIXaBgDCdmhSMTtMF7dWgU0lFl2WDsqHe9JePgiy89lS+T03ME4
lcAyQ3TalmADJRcIa1hzO6SdVEyBvb2JcZyrJXI/ifX8ieXxSo4wsRhSmTzbB2o1310FInUAH2Pn
sJbIBDpHVjU6XwoPzvmaA+g5khG8CsGQVBETvx9qtf9qXj8K6W1XKaZT2J83xNPxFCuGoSpnTj0H
8ryw6GerJbCTf+wNdQtbuknWz20eh6+GIHoEE3SToiHK1vM6/8kMneF4hsK5N6wemoFr/feBgjGR
JxOxL7MZ/064XzPNHeGQSoZ7gFO4uWZT1Fq337CGT8ORGjghAR9RN4OJ5jNIImsA63ytvECVQMYZ
q8mbE0bioB1NqMit19fpPfVxKDHzINeBceijTurD5EYi/QfpHmUceggt10U95Gtq6IakbmDqOGjl
UIlB8n8wq3yoR6bsD8kHLn7N7rBDuBnYIWTk7WpRrWmp3TK37+sIeZ7PENIG04QXpb2nhuDlsNO9
OHU8m97DLJxWXOaXhYiLc5IN2mH+4SrF4bN6+HTHrSI1rLtQLEopqdYiJNRyOwFwwyVoL6XAqhw+
3y2qdqWN47RDqjrrnq5kBCEyZIOZror0JLQYGEufRuXrlmuuRei7FwzXDgreFyQSAlhsoP2M38WT
rqY7Ix4DBib1IsZhuNfZRl9EUGgii7Syj46hs0kAMr/gfNofgQW35PAXYRG3NmBx+ZXhs6QJSjIJ
6+7L9nCy4qRd+6xqyrXdeCGDXZBJzmRrlPNH2A+sboujNDzjHF3q/SCoiUA8RXTCwVX1Ef8Oyxip
I8S7D9mid/yd2l/NNl//1q2AOdgen2GwaLm5MqgTMjfYQXv0on8xTiSmgm8aL8ksvlaFFbbtFJVc
043rAOpreCgPiN7ve1WNOtxP7L+LFngWHgDU47RGhGE2hRmDMQDRP+jgrIVk4Utm+kYOinE5zF4G
WvJFfUrrAFbb7JQTQRuIvnSp2ZoHmsTLwePCIhjwmPa8Zg4GbknCuXyF7yYej4d+KKx2be/E+l3e
Aez8izDSO5NYVTYBeSot2UMrfw3OaoJewWk8jAlIjOtea6zd05jeaVf9sbEtmO19nxgBBYDSwEWs
lhayYbinuZOkKH7Qvf5OCkj7FZ7zbDYxrtrk1uBYf0wFumRMVbEZjAXEK4gZbVe7r1fHtp0sSHjD
ywBhE2qWIMzkmwvJWKzwwG+ZnvQ/VsQmLsaOXABoMab810VmVnSeckBZv/+YYIwIQQZuOaMajfff
39S1FxcFckapFbQZQdUCZR4x6sXtvgfK54Riubs7WhlAWbrzrszOAIT8NdEqIbW2DNHOYvdJlUZM
MHhjWoVmtjRcwZpjK/A/h2iJ2N8JZz3vMIBDrgNeFkToHGk3YJibXbV4XegIYNtZNLKnmRVlNnwF
WQzWffJ1QwY90Uhr5DBmcfatT6YfNCZKf9sEovNkhkzc+tYafWC8kvavH6H/XM9lbhuj5vkdH+y1
zR4yeMzZ9v+PCnuJp4i0Gt4YFhYuvLpiIAcPRuWLllBbmTAyeQTik/8eI2AJqt7/eoXAPqBvvpIk
X6c/vdw1Me0hyfcuUdYGvT77TGtLoXFn328OlYlC9YLZXbdMRZ0RfPXwthH8rAOO2RAWvgzw5Jbt
v3IoCUNh9KgovJZJfrqQME2zINimECZOxFBgiEbEQQyR66oCRdNlrITMMTwIzHUuAsmADRzbye5/
hE5sWhcAMaZCfB3zYXPGCTmFhf6gaOg7A/FOLFH0zTjIl7vjTijJaumifhFVa6ufS3xY3WaH3ck9
X/91G5Z+E61y+3ek8mHUzDmN+Q6/G8sw9AQ+OjvvJxyHmfgspPLKJkJ3C/TaYB4Sja9LPuJCOdWN
R7phHHp58TaqzxVKl9anmc0kokAdoZQhRj8NQGAtav3wGAqnu0njnTvnJMBECOnXJZqo8oNT4z6q
nHKsitEca078tDwPwTC9IFKUN/nuJv7wW/EKpffd/GEt8AY42Xi+k4Bbm+sftD84jOw4LYLtR6UR
G9Ldg7ZlTzGM2BdUDw+ladVORF5WsVUEbHjyRFTXIe/2SNK86jQaNdsCEK4AnUBUFQ4elTTVyDbC
eKYXNHTMxE8QJbizW2Worb8xDww2g1yEff7ZPCYbU0aVaO1sRpTfyiLFpG60oZeHFp5OnSffdSrn
HRtLotP2whE0nd/UHSkrDm3lHU+HLgKNeQdU36/phs5OhRVN7nUZNHNUO4COxv4jUbmFB6zrC8kL
mL+GpCKuH3qVIycvfFE290btMmDd/tTZZoDXhNTJ2q/Sc3UEkbFCKhHrB9qTps97eRBnkrKe/CVg
rk8AyegI16godtuUWQKH+z6rHaRWE2/0RY5FjzE67k/uVU0PP9PUhBOfhh294mdk5eF7k3K3XCJ9
pRsd3W/JRP4Iw5dmJ4ICRibCa09be0rPhut4I4LBMEStPnISDC+fPuLYSvV5NFdaeF1ChMag4tdP
jygIuKR9vX1ZkAaFLu2hZWPDnpIZpTmcxtYc/gzA7He/Fc/P3wkV3c1qwB+yYO76qXi1wgPd/Ikh
QXo9k5Sx0vmogD83kzD2JE97C+iAs2Hm6Vmc2yTBbbePTFDYiv9AXDzbrmuhjPs+f2MC+rtBx6D1
QTMh42ticsMyczIglo3d25Yzd+TmfFCukY8631eqMH1bG2mNLo2hHflRIdzleSUrpQm1YS4imixZ
2OMn7mQijNOxatI37kTcaGWaiklA4bO6hVs7F/KZgWajriKNRp0Efjg0uE3lLCx2Gp7C8uAqtxqr
3nzonMY16Tw6gBaDa2jo/5IbinLiInwPrgeP8K+ZhvAe7Cw0a+soWLpds2omr0VPouOaWfrCt8hT
SvWIuj4KJ8wTulgiSs+1Xq8Ax5rOKaOtTBo+tz3JA9XfOXIWz9bLH6KqK1iBIakA9FF3mDZ4Y2Oi
Q+4yP8J9nfTzLRBqPu/iKWZnzUBSRF1tdOaSZ1j3tzMzZvVTXYq5HPsUETqy9IZLAS83lPfIq5U6
xqubepAnyAnDc9afH5zuwZHqaEewBo4U3urBtLyYWZlTjDSzGFH/jeoQAAl+iWVkPaXbEc+IhJ2U
KfL7Ug2f0uTfvZrPG0PTybaMEhpzQQfoDaDRBPsDGbCblB2eJdqGJISyup3UeyRFT47sBpcOCgcq
6lBoFewqJiTEgAsy2cmkIHdSgvlGFkKNwrav6WQ5K+Tyiu43GfTSUEhtjuTM6RiXqV/p8tKNXU+n
uvClDj9HUWVkP/++CPlAcf0q6n6pWJt+Vm1tqrNgSDgD3eLkKh/rN9H50/nQLSisgVkuxZNhwQxH
cRqwPYQTFiF8sllKKiaVhxOOCJKJ8XeWYfNgr3NoaYTtwNFEZ4heQkg2M+VaU46oe2nkazb2HaLa
DjIVR10tLJsmbeoFTv8mFePCtTmRJ6bYW57y6p4G3G+Yt1VyDxaMgW7OwNIPzz5g4kQTyKW7P7+q
Mh72G0rEhBT67KqRTejlBGWF14eL0CkOF3wH0weivEw2Hj2qHZ3T9s7oobxf57BIQ947UpuYlt+w
qEF5Ml2ahZsG71yIlyFpT/Lg5r0if2Wru5GUaO6nAuULbsY+ySMQlPh7X6FsJzES0k5NtxeXb5XM
V2C9lEV0Y4OrmEMPR+mXNEDPoheqIwcIaMuXo0uOKy2HZ7AbkBIaEuYpgHx+b0T3GaqZM9L/2WxL
ZAagD0+Zn3IFanIoD1O1gnBqKk8U2pxNvj6bf5D+WO503BKVxEPwcwoVLnsDMIvwrsQQTOLMkCOo
HJ/qPUSVXPxkRnp64KK2WAoqRGFjnJOy6kww2wIMaY7zmvZqwP18ah7gIGQYTsL0PYEWKTbcxC3I
ysLpzSYSyC+yQpWRiOC5oS0fo95K5tLJ7Eu7tm8XTfiYsdjixe45tekF3acRhaKqHZaBLWbLvPxz
ivJnZ9KFzyXiGw8vtPWPvkn0eoIVz0iWMS061I5fm93tlk48SJpUWI9dqn3DzjpajvoWijNcyUc7
d4g0FuIpgalX43VYCyhbCOu1uN2QOfLH6uAaeXVBD+hmG6nbOcxXjc1lWhKks1JsLGIFbhoThvWT
SA0RcpQbx9hy5+bad5Pk3cM1Wc/xHAXMatwyjhAhEAIFiwRpBjMCU9IieGAT+tEpzUx3Cwyu91we
So6zxdtaRhjxt9MVo+VbtmyZD+coJghQJL+6aDku4s3/LXIrbeWpLwbld99drhsZCj0PhbUcIsWK
UWRueEErGE6XqF45yYTAnT5LgvFLXxg8nT6FytJbEKMTjTPxULLkISTR1pmAdddUKhudjvuaHlkL
1JPWmSwwJwnXmepFmXe3o8SVe9+be7Al7AuIR39y9iAj+d3ZX0QDUaU31gTdxn5Kg1M02B4n+LYI
GWwndhavb0Rp4oUufdtQKOf3dyWIqsuNQCFpUAJ3UFbS+aGdIrjF4Y4LZw7jX6z47V0TG9uGE248
9WIKa1B/IBlsE5nqDNQBXimnpbopR9sGAoiuwbmvJ9wg6x5rgvhPuE0Hl+iRYCWc4I2zWCrgzcWA
p3K/AYFgKnvvlLq0AQzcQuHNSN0FGdrhvmbnKJAKDtyjmG5ELryvY4wxBFKQmQejlpDBo4iijXW9
PUXdbX1X+lkbi/21snVpJMdQNin4LGBrd8cOUEDD3TtcI5wX0uOiBW7m1nE+1zrJ9aB7wukEvGHk
qf/oQRUQAgOT1X5CTxuvoP9V5ceMewU3I25XOOGYjAK6NseRGWyahfzD/s2TTnwzFIvtXcFlfOUN
Q+7KqdlPez3cE/AeqisQMPa5krr5hWodtgJfOk4iVtx+Gio0rnFA8gXubvsNjIBiEXJvbFbFNoL3
wMgnVrd/ylkHqaM3izS1W29Sv0IfHABaggnKUUTQGoQrdo3fLa1Im/n/RU/Sopo5IapjlnagOwn0
paEVUu8fgYHIPxJpT35pu6Fjap4m4LVIhnRhMMNOvdmyDKDgowszODDHalZc9lUxj6FtVYTFEMm5
09IIIEbbgAbZDZyVU0sU9Mpgqr3KiDOm6cKqJkwEy/ZqqpNqNH2btAmACexuIyK//Zwdyz9pnhdY
OsLUSu2tgHU5aVlYquBGc58U+fhRgl5Hhgg3S8GKlQu2dK/BieGEbFPIvG/KOeteSEn1VkbNXmD5
4IpeQVXhbl/Ulb/zT0WBQsFoi+CJMN6yBggPiDlbtI141vM4ouuMf93FPzuA7X8Ls9aEMJpldRRU
nVUC3wFXqXrVuG3uk6vwmW7vB9iEKeIHvU+UK4BFs1jT8ZLM+sb9DzivnEW2aqWWNKKldk/oWDoj
tLyXAL9lFuUcljSKHRIvSafMjvzjO8aSUl4EtQYjGsQoYWifOenAlpeD2meFKr49nSH0974dbRPb
PEZiEEkzAkZ/aY5bMvebmeRO3uozukcepil7B3hMyAL2M+q0dJouZlTmPq2glTS2CLvjd9E1H8xW
PyiJyZA2C3o1aeh3PKyuxNcLx80MNknbPBNEO+KthXKwmiUhjF/XxRiJb3CVr5IaRPmK3mAc3s9B
+IEW06+MAdsaC6GpV3sqjGK8vJBjwuChvMJp7OqhCY9RLPFVIRkRC9BKqZMm0iy6AD3asIa7L6eA
HNofNZ+pQOUZU1o26ditlvXh0np9U+YJtkND/OaW+is9r8DKvt72OxEvH6G4P45RiGPUQMXzMYHB
LbiIm5D56lkAFbRA+kTbRLSCcVnioZ+o0O+XpBXCPT4JeoOAoW/MfP3Ti1Kq8s/8ACFNfBQrLi17
ffAqbzGJuNK1KBTyiJCU7jj2DRn7WZCetndnJYzKdl1ro1Wj3K4UIlUp4XR0BMJbi7Ogvlb3GkP0
r56rr8sO6oO3ni23TjzcL8yTt9Mma9ZmfYQIYlx9sOERdGRML0Yvqq2GuovgqWgaTCWJwISCfl1T
HDxvJKl0Wkk/OewyoGxYqXKqRh3ia21pv5HCUZ2zx/Ymd1lEBVGl43n02g/nVe/cf2gX42Y9VNC3
PGpO2gMoPxbM1FCO0m5s3nN894TiHUG8MWPn/5Pjf/JheYA957ky7ToqE9YgL1Gml6xVPHmUxhyJ
vf33pmn90Kvnai6FbOCD9vclMs3Vog9DHjek6W0GI/xSCiKK5OTgBNU/G5IaKHHP6Z4Bp+VnnFVW
fHdjJaeKuUY/WeAHwbCXCLcrOQmmTezW4LUU9VzT8j8VPkl+kWF2poRrAUKXP1UO6ME38sFitO+l
x8oELAnQgzv6Oz1AID6wfh6JknAl4urlBrpc11ewFq72TLPskDST15Nw5wx3r6eaclM0FyGUq940
ZXDJ69eYAlrxIcEpYqBdcwSsgzEqSzp5+JqfkX1xB9Cmt2FLz9KGLYZEzXf9/MgrTiQmSFeLZ2Do
GNC0ol1V/BdCzKEeAtTGid/EY85vJrtln9mf4LXZ98ix+Yc1CHiUN+luUO8tlqTQkwa9q0QjppB/
toqoleKHLVHYYWGjmDyDcdGGdmbl5f9VEEjecfXyC2di0uYnVo2vkzv0fXcNyucJuYqnRdaSWOHH
SJA3ClH0s8y6ZhgMcsy5whH9aBUj0vlfzMwE5Le59L+rwZeQX2H5FXrLR9cVtCEhZOC5W+kA7txZ
l46h9NjL2d4+CeGuzt086iyowFgiYRtUMhj6Y4aTyPGGhiz6gjISfZNbP8zg8ia+zwkqiiKYoZ8Y
uCVOX248aQL3UV6//KXJzlmeswvA97AXrQSO4EgInhgHR2yEK+IWzjVN3OWKx+HImVF+9uRmU5rH
kar6pVSjyW7mZPbG7Eb/5EgJTKQqWMVl6JcWHvgCPKqE/jYKyO5mETe5UBlZe450ns/mMXoygEb5
AYoolmkXIhpOfoODEQdcWABxab5F+O2beAy/2dQrcuzncFKFr4V/DnkzBtLP0yiR6VpgZoJeo4AV
/TMXWrHImCCWW2+pOky1ovO5xA+pfcg7HnxN/yQRrrl3ETgPHGC3eaZdlOn2SlC8Dg/iItsktmRs
rErnhxRJZb5DN1kewC6QZWsv88Zz2GCAE0Kf36BUWqN6f4V1bsj5aakVkJ6rI89oVGpvWQ4/3KZF
Enau+1dcQTlq7GhFipzhUDtvgt4fj7qsh9J8V3mY2iJ5HTCkf8r5sqpNjOaP9a3jcNUirmwVhebd
ZQQ+6oRlNxpYW5mWgs7+1EAyl9IIr3Or6uerYkXYxAQnZF3RfvoqrSQQ18IQIiwuNiPootrZ8EBf
wdPIrUOgzPvLFBgcr+iM/5C0gmlTVPVz59dU1i0+qZ3KuVXLSQwsEJiN2K04G4crMYtyu/nYT/7r
2F+zFGLj58BIo+kXwpNbVyBaBjtLkJyLZGFGDRjXVEDY5hluC5dtQYzBgW2Hf2izpcZBAZ6LLWYc
EQkuYOeD5r4XdpSO6MM3YdvCrSDTsVPxDyUlDRstmsPKSd4AFXG8yCnyeIHtxJAkQCcZANl+iWYl
TObw2GF+haRG8PBksEEMNZ9nV5zzi4GDXAVK6NxI2RKjovNMBGP/yliltjvfzE8uoB04pF5jaUGl
ams5U7f1siVZj9iF4dXWc6YIbyeTKjRdLOSUedwSWtw3eMKSUbGkhGYemPvPO5c46BaFf5qHvDdA
VuV/biOSgAzWIeXVOnXGeFSGb4ZJi6GjDOOEIH/DhSIA7khlg1E+bxttbl3KVRzGK1GOe1uw4NKd
UJpL2ZBOPsi//4USQ3gosXueNRZqqNejDutWDqlEOHEkSYe3TDP4iA3HaRgAEXGian/24k3qbNBo
XUXSKoLS7e4wowvmFZJ3wPZrsLy9NKWF+8onD4Lo6cHSju6YDOVRoXPioK+aJjOdZGteoNXRTlBG
e1a95fCdFWtJLukMPUpd1gy0nX1pqm1za/DIIuSrfCRfHGBew5leHi+r5Eqpumd1r/931HiTLXrc
fTQ10al4/3wmPirH0s2U61UZ2lyml48+sHFQqNi7MwhVM95ZbR2U4vvruHW6smrETVIEAMVJ9rnV
qlId4yEf8pw+SwYR+rlEArJry1Akeaxy8A1rKxsJhnU4LK8o1Wc1lm5P6RzA/FbgzXkn3Uk2XjGo
eaNp9MPPLBGjCqURiOCc/n3kvh42yj1HwsgEkYtWmrLQK+O8jkrphG2lxHqwRB7rHs6crrUA0XNq
iD16ki3UR2F33EBSM/zR7PHspUZPuYXZxlxX2L3UxEzE4Ag7OdKSuyA0ilJKQiavidc4mcmi2cSV
h2FOc9joYd6QBsfqG4xpqPKif8FXVsiKYjMgBjuYtZjNfKCtopwu6qtPJWLoI0hxhUw9pRZto8FY
sty4Cii489qG9ZJ1TUH+cZMQlRWB3AqIYhxIt+swDj5exV0m6XhUpVwS8Bt5hXJcloE/1bFYIK1i
NHw/1JGTsfsW1fUO9qibfF5sJaFTaD2GizAEmVHpLlT7Ya1webMh9ZUKrRdPVX4OCHFAZwcc5rXL
MCfg3YZypM5pcuzdeuZjXBL0yr2gkvrAVSHbWHKfe5vWP3qSNRDmdB4iR37yFA6qaqgjxyNwhmST
9aIncKVrGzKdAnkGLhRblgXpWOchfUeV+ZiiEGAI2UpD/aPlaijVKaXfvuIJ/rwAAYT71J2JTI1V
YT5uKa5rNdUH1Ha3ENlE5Nw0jQKMZxj68WZ20z8HIIcsOhTQIhpaQtRQVfcoq2Kn99iBCFJAMv3/
HGCmPL07cbh0KPLnhPoLMbceqXpCmg6ypvPRjxu3f1vzv42faPDTr5RYtao3F13hbNa172UvCWl/
U2Vxm2+s19RJ7qZQYzO7LTBZDgJUUu0cKKRRmcxvqD8X3JRVxJcryc4HWOLN2OQZUPK3JF/bT4Sb
DthWee/wyrm980CeRvhFnxDfWZ2cSNWj6cKap2Ms43wLomEdml5TDVhcE67lIjfOcpOWxaBziTOv
lSOUF5FslB6vmQWLlrOol8Ub5G2oMgSiCpBpRIOD3j1MtZcdbY5nzmrBmEY6KIJl6zl0TJbebrBs
0r6wfWpm7moESyVEXQ+KYv6nncu5OulxlXSAdSGrXICe0HNo6Y97FuUAA4kW6S808vEicVCYMEBd
mbNo5NIki5J4mNuw6VXeTBul86G1C3FOdWCc6w6I0D+b8uyRvJkzPQB9utRcwthqEKQ2fDsCdr3C
i5/PrfHPbELWgBlWzsm5NEb89vwff0xJr41b73XjOPEaxP0cqdG1MlWJWw8/j0yJol45mBBO4Crz
JppX05sLjcbyIf1M1xWTAc8vtu84qb6B/y3XBUUmq4CvaxJyl5MNG7nDCvsn6c6EXItrjhmbH/hr
4uR+nXiIDnN6ECcAwwZaFlvg5GmwlCRua482v4t5dwrRDDPASbmwweOcyEb/3WMfCgCU39etnjjC
qOAIWEZtQGyDJgd4Pc7H5miUp63S53MROlBGdr6QybcqTwE2BAgvpFJp6jHHgNx8KCZilV0sSHiw
k0u8Gdvxf8pbbC7xTpZ2QN4PQxKIqXbKrqK/9UmBAGAWpaku+JoFGt8ZTSbljYWQH/F1YXt0C6oN
4U3QsnBg4AIP8IR005yVHrP3sfMk2MCE4+9uyTnI4myTNP/E+1shKtJqPhjliJRXuwlAZAigWiY6
XrKdTuWBRiGMCLVbBhljRdJRqe8uST+1RthkdVDUoZ2z2adUk9G8CIQAWxXGPlY/jFaaTiesJ88t
ijaIAPm1dwVCTVI3ZSfLkE4+h1VwJBGVGijpSYiz6tE6PlC7JEC57O3LqH566qcS5EMU4VSeKqRl
g6LnjlnVa79HyTKUyDiNW2kZrPduNrCd5i+xOJfURIub34NrsDRva2qRgh00qHOjrOp4H/lFQA2W
JLkgoT5ZWlqIicoSqro3cq/pEeyIlcNGBo9GpkWXnRtTizR3GR3SJiGXeLG0OPxi5BhGLQtrEsQl
in2i3aGjzEu7ZDYevLWnsgbXI5eCB93NiBo13PrttIih3jGE7wX/yDj7A2RukTovHWYMNDbujPpS
9J9qX5xAQYD5FLOmcuKxALEYjdg7VK8WGyfsO7t1lRYcMloMwqAehO/AtbgXOST0/zWTNl4Svpyl
jhhQdFx4jigY6PofMZR197peIpNdN0UsImpDbsMs8zBVRFk0orpX1EXQLDP7Uic9l9m0KdziWUPH
PdOQyven/zgrYt997MRjVB5bbiX8tGKmx8V5mfWeO95DxStUHLd827g1ED1FfRl1Ka9iUEvF6jWb
DTg/wGsGjbVRThtvGHalqcL87PkcnzKj5bx1TZJndf0jx4jnecweMYjVvkEPwtH06PwSDv3K24g7
q1i2Mjy5MNIXxzPgRQhY6/jE4aIFoM0H3CKfYLnjLH0r/1BSr0vjeOZCsY+USey3Kxj+CK0gSfkU
6adZKqxM2LzbEeL28WcN3ah9POkVMzJZcm82JzjzsY0eNLiPgZRk0hkaw+iZbmH9d7lBVVsPNK03
TSn7Aw44zpiUHBRGIEsccdiuuI2ar31sDOoQdFsNr4qCaiteFXIcp0p5jWhWWpRBxQKhXvcO3p9H
7RO5b9bTfwJEcwzRvbjUApy+fe48Ay9HB7J34qvFURenckVd7I37MfSV0NW9KRBlOb9Ipfu05DKQ
hygA2yRetgJkJV9yri/xrNPOWRazzW6LOABcc4mIxez9HbQ7TTJVCo+6iUmE5o/4eyv3TvvIDldl
UQ7LZUoDGsN3ASZt7vaTUK4cVj9i0yAqEpCwpkGI9b5Ueis4QhSLOtEAcAzaFc95oUZ4S9LXH/CR
5jdPJiFXWeoGPB304/FKCLg++tv2yhbD+6+4X7TlUhJ6rrltzS2ihZ+9M/KDi5L5gFSbjGtENFG9
6Tt/MYS37W9C7xdvZbMAh7Yh5NWaVdRZFdjduK7G9rfTv5jXhbmfud13QdvVv+qRPbD2VnF/RMhT
iUVgRSaMqkOO0sD8J4pkn/jwt8QZxBp7T6z/c12UqQ2IEcybvBwYEmVPSna4DHYFrd3+DwBFe4LM
T4RW1dKTG89j9j3x/z5u2VgFuccdFbolTx8wiuTagYNYS/kUvm7a3Si3DDbSDVKU/L9ParD86awJ
NlaCMjwyR24nnnD84WjdVWzR1euu1GLPEQX57BF8hujgwqJ0PsK5hsWIVBrDpZN32KvjL31Iqi+n
jVah9QxcvJyiUABuRfbTO28BvJD1auJgtP/CzI47j25umbjDKUIfSGl/JahWgb2kmYA3n4MAyGwQ
+KfC/rpVjPxweEwkKphxsK6DGw6jee/GnjfKX0syNy7W5MzJykbFVjVYg3ctdsfcisWUdoUW5sCB
8J6Iu7V09qJQ44dXCijqJ3vIJPOXq72iVxw98W0MuXGh2uZfuaNOf5Ro6LWwa2Sv+zQ0R277baPk
hm6w4XbjhTS6cVMNf5nG3EkADyOSAoVS8OrZJeNy3AvaTpdmvyVLwjYhHghXF8Ff15YdTGygDFAw
108EL2a/Qc/4re6UpjnkhL5XMpdBCuCFhGrKJdBlCdwwFfPvQ/iqTqMypfxBxuWmggm/EUfkU4ZX
CeabBfsPt7yRX0JgcnhTU1GccndsW71dR1tK0vgiSlMESfl5dXMTDoY437C8MXQ9SjQcNhLM7Geg
GuldeQ2+khieGv+ojz8CSO7eKbv7XO8oihTA1RM8saBvHGdnA7zddzioVmaPIrBZKnscRko8uYRA
l6nXx+DBcOwvB97td19l0UPfOdw3DsL+jponBy2x5au0P0g53hDifjudP5+YtH7dLaerEl/y7v14
rfFusuonQH1AE+ieAHDlB02uaSvwmgnOaJZrt/G7ZDMG/b8phBr4UKSupbwdIvcK9pBQZzdvizQe
mD+0mmrp98qBggm+U0yMmqBB5JYhfFbwgfpB7nrh6jHzitKVLEd1IC8AQHL5PflLN8lRLRW6utsc
Rw6SP1bz+ot9GMRzG3BD89jWkKsBK7QnX7iv16Ae1m4+amVVIBym16IiYQG3QwgCOBI8Qxsh9Jin
+4JVn3G5XIIcMjYHPDgjsci4BCSgUDgX/uhDDrPpmtRbVOxrzh00GiATP0SNeyrrR7G5cGmSiCC7
mpTE/gAlVcsSJshPqhaoNNvUSwrAiWUdfxsR42rW9uWv4YRPbMldgyjOTqmPT0mMKiRUzeKF1+sF
ao+PT8K/QWPsj2mjrQDsvjDSjjH3qRp8Lh6CU7XmityEjLZPsGZ6Mj8QK/J+A5Lq7QTobOQlyh6r
Prm/eGc+Q/meeCJar7tVdFO/3xHI/NvMlxGrQPNo3yDTL4jsouK7KJUqLhA3yH/XwQMQ+RypcoMs
wh0KjGyi95lEjcSGR6Jxgli65kdYI/oRNqG36sFDkM/WifrASgMTRJsvMXbR7iNGJTmHr07gh2Aq
tuuOU/PXVg9FOfdnnqTCD5uJxRCxDV/oLFRlXbr5Qth/6H4NzAb7XYRUNZRG4hcPyJ7EkRosV0ri
ok2yZmo+/6rhXM3ajGMziiGQY8lD8QKbOO2UfvuZt6L8SKta7TDX6dVxeELUBxDcKxWRWAnCaDmR
0UCJE5b4Jn19Y4LtaYrGRivXCqE0JkybLrwv4DmVJ6QMxGsI3dZebseNgWVO+E7yOdqX0ue5hZ0u
tlsruDr39pbpthicdJ3vEq/Gq8ZrDq1XUmv26p4MNVg6zsxK+8Tg1JcrqsuB6Pc266ynxDMhhH17
JsVuN29T7MIcQ1GanwEBpdDopcxndF5Fu2DP3FV4/Hb2R4wZQSK6+p5Sc9Gxu2wdS/o8Euohf/We
vx06zdhxk3ZMt0ES50UW2huXlnGr2L7aSQw1MZPuMzFfGShIuuuT5RUYJHe4nv9HvTdnc30silj6
SIIjSikn6IFWc1EVu/6pUGITyKfZK384CyVVBWnxXa8F4haeNub7ndtOiQ1sp7HJSbjb9TCZfeeV
6ok/gGcG24CfmY8oM0pZQmbJlE+nonOFVH5K5BlevNNLcL8ujZgqlxTuqVALFTlbsK28yPfR0EQb
X2qZ/xaXUReLj9mgGnfVMoRNZhAy6CRP5ucv4Ta/2Iu1szn2ZXVqT8xMw+4DaQFY3pVJd9WDYB4m
61K71PjXlqkZZe4fnMhEnjm8vb09pJBdWKZ+PD+2UTb97x+p696c87WAJMh0m61Jg5SwvvwQqRL7
nktWh4CF8Jtrzgr4F/ueQnt1kUBYqONilSHYofrN5DuOH+yI1XfZyPiZO5F11j+gvJPkVJN5vUE6
3q0g85nwMC+geLRCsx4DpVQpX2vsJfUNYxOmY5W/40Mn/VJMbIUUmxhjTNKlZzu3yPSeikCh9/vn
VqaYrvQO55m0S3CuVV91bLlTCBpDPbQw1rMrv8NspRGGcv8ZeivlVoOxydBnSCveYwG6T32ymD10
msV1gBcSSUSLYBMMWxuByTRpdQOmvS5fE+aUGt90quwjdnbDUOgW0a4mpX317sQ0rzmTLz5Sndeb
KegSdRjAHqreKNs/BvdUx3oV4oaqrcUkcZhq7e9hqoUSaPY+IsTsdlXccU3ro8gO4P7b+Fz0mwgJ
QxS09X1LAa7WO7TXvoS68Thgby7yROPA1kMYSddS3zLRWYhhA+Claa29gD4A25Kck5ZBSopcFAzg
Nm22NgvqQO/Tc9nn1fOn6t9nGRty2wxLtMHbtGr3bhnnJGQ2QHien7zCM/0R73n2NIgqo7jSoeBh
xs56MjJzI9O11yH0n+wt5tXYSBdzqCYwSjl9lfEKjJVmtYKUOTOfL39G1fhBEXW9gttT8UpKJQaD
MsrS5l5+M5fMUYaNAdZ0kFY9OcmlJ0g3+B3TLoUcXkTyAKhHDKozi9z04dFsIaqX9D5PpBzKFago
5SoFLQ2xY0sZ+oXk2OVIWTwto4nTJOK1CiWf5Z9LnH5yFz/B03keBvDFdZ/I2+fMlhi8gj62OHUG
s8pkmHFdZXJ1HGtLSmq4cwnw4GrDZKG51pmRKj9dnCUAlIN0guKX2aQ3AcKuUefPwPwhejg2ENPY
TvtxWL6sDBP/lUvrlL6Qx9UKABsTjjZvC+y2ctHBNM/ynR+ZPvQih/dz9hbUDLU2GAftlaC6kj6B
ZNMaWsyRa+5hPhm6cEvZNilu7tg0MYRGPRnfi3mkwwYAJOeiy4V+XfED/nmkLnkDmrxqL6ETaxR0
iBIGHuCO+YoQgW+qmSHdSa8uN4We02qltnrLBEIKfBt0agHulQTizNacQDFMjoHsAL8/SXQmlz1P
WGqAohVBd6XfHrHF9uHsl4hjfC1vniAQ6cnCCYsDEPeXdBKPgS6eMQS8pYD7BrZk5SjH7BU2NWHF
EjWLr7KAFPHySsLnyWvcdxeQ8MvxkfrN7ae0xE5cQo8IZI8ssDm0+yu2UGP0NVjdC+kUPdLXIAXR
g04/DoELTXQBNPMrf0ywb0cT9XcLnvKQ1TrAPqwojAe/glHOhZBfEBqIIpIw7oB3nGqSI2XHiBIk
V+c/aG+T7miviZn6RDetYJWE4smyicKf+NowbJwcEFC7hznmPmhEDg/Qya72gjXooOIwNuJ6fYYk
If/+0ct4FQ4yKcp64nYtOPWRxMloT47PHUAoKcEDy2qB9ULyIdTGea6r+xZXkzwcur8mwP2GKpho
wQt2aw9SAOHT/39gBNCQ+A4kGE7GHrDUMYaXx6nRUJL3xS5ZAUrs15h4ba1uQYiP4yrJ5q+YsFf+
y809PqWyV4dlf62do8tCpGLdMn5buJmwCxbrxYR+FZkILlSysR8RFBR1AqTnFy6KtIPPJmeCVt32
t3NzV5iuA5xh41uC8Qjzxrg7fJ0JIi+Zv+UmsDR7Hglw79MXsDY+o1KH6C9KXPP6knXdr/5QwQWh
yiy462DUk1f7R+3DLI90fdk5EKEYrfU/e+/itLswc8P+xunVrxyOU7qP3QhjY2H6zli7XdSX5Q8m
l8SSG7a+DCKvvAx0mnMSwQdf9zF1+Tqb0gzlCuuoyDkD2jE/v8KS1OjgmVeetgX+KUSyLOBRKOCp
Ykqnee/c4zwwRpfA30Evnq4Ao2LjzUmjVLGL+1NLbBRWfRv0tLzFcxntGzADtUne7PeUs/EtOzqq
CgGBgJwVBm/0SKIU7SoiJdW36S+lkCNSb6vIq+Z7VZZDGiDVQ3ZSFrbw6Il+HYpth+sr+6SAF9hd
b+Bgcp93GhMuTQU3+fCwlzRdv6vyNPchbp9Bdh1clf3rX1c4zX3WvLV6caVLbndb1zps3COIAA8z
fPpYChXbYmz0wzlf/kryQgMu+uvzjHNZXkuXpe5jeCtA6xnqymeaecHphLKRZFUZych6mwsipTJo
t9+MgFp57iyNpiqEq3h00zr+lUijmA4tWN3+KjVK1OuCHun1ENa5iQzWUe310qQ0Z4piuwwr+gVW
L53wmNQtMGIzVAkWU3qjIHBjNeJvWWdoE8olVY9+/LLmIzFCh+qBnSN4/Rr4dj7x8U4EmoAVTAYG
JlYU1J4q01L9cJDJG9PRRQ3rgREp+t0qGA8MhMImpcmE+QmfLtW0YhVwZ6B0aaOtEkUbwAHel82Y
sNZGBZj1Hv/all4gX+zbNF7R6kwBqeMhKbfXhXtU7ulU1sKT55kD2QgAjA0t4bDwAppV04mknxeN
YzB8Zubn1KQKawktuB940yYSF4MESg47rpeUYeuZ7J5ZDSC/gH8pqzjLdksyIrF4emPOlG9mnbal
qIb65nJ96emAgfjMRORsCQZ9LdIFpmIGlU4LwxXji/3ldD7OAWDfxWIejANyzu0mvD4RRViXErM3
VZQlXUZPk/DYNu4vJRXdjDJv8LkSpyfTn/zFYckUcW96O6FIkvFSqb6QzabpjFKfRXVoXQaXIpnn
Bt147tqgDCRwfKv9mLME2rbaCUfczksFJZ4JaCobSsq82m2/kHmkaFbhgP03kM9HnLZJrttEJoOO
wm95xGSM0McFbEMGuZvHeLYzpSiFBkVbGO2OW6i3NFAOY6MoGjqJe50DK2Brq1QbN/V33dt8qtwl
9jZbilBOj9o93bPKcfKmvLUjMYTAwCPv2/dBiYE7rL5Ou5WjAZ1bY/XPNt38oXF1kJ3nKjYSizP6
+7QcNgtI5N63we6+8jhRmIx/yahjhQXsasTs90R2TkMNYDRWLy4hk65zwYeBYaP84JB6qdXw4jaa
XDaXqckTX/vz32XrGrRo3wvTQnRGRNJV3orfpMXuJ1/5Hz0TR1gy23LIwbhkQwAZifYUEtMRD2Ar
gC+USQiNs4NRQMbxWBN2kj1E/QFx1NJK7gDylfqf+irVpeQ8Yr0GOkAGYPvqzCqdhbB0kFrSb8Ck
iimav8Wb5Qp4mZbyxrrB5wWjtUotW046lvPGO1ySbam5JfQ3FIaRQuT8PeMaftpcAVhHeZp6/2n5
8LegNnJh1eZhDFFEVbBrDAboLd5xSC+MSjigWOSTB/cY/+lYl/qqZ1t7eJkVNtQa0aDdjFzCTJ5/
MSY9J7OcrjSRASA/VbDA+nEcKyFS1QcyNL8BwiV8wF+mFCPuFyibbP6oDjnF6kuxIdPEq9RMmCI/
7CV+hla7xkKjhklEPVWHiE0KoUyA4g0TOUY3mMjccKjIFU82rXk9OUF223Hqytu29SJarnK3IFio
2Wjj7ZB+Wzc4+nCgzyFRk9obs3pwI6LD7RZ2DcrYXKYS5d4HWAaMCkrQf8bz5y9JB/OXA8LLurCb
0kXHOZfPMk7oyPxJjX2TILB3bw8+Kd9BcaXGyv/MAv/dCn7YjLqdIkfHw7GdubxZ5Eep4TM0AZL2
fsWt76FiRpIUN94ooaXJpZTkpytGSZedijfKB3bqYx87edv4O95aS6x49atVNJuvRjVusmnLVNYn
4jupholnXk8VAx5rEJJ2cqGNeI+N+vTBSE/vyQy1TeRCbndyxRHtZkmqr+/rmizALpAVE8iMDWfq
0Glg9SipfH8gU8fZGh4Z4fIc3tpi+olLNww5aT+RwzspDMdiGu8D+wd/9d56mNyHPBZ5G35t6XbH
J2L8zfpXAWVUwAUFRXfVvMnlIlc4O2GZx/BRsHJgUqqZccpBSvzDhmoYc6/ELncSbeOeu1SQ2g9X
eQQXZtOHDfvUsi2nLphpRkeTxEigeG6AcnwcNA9HDc7hBEJtkEhhV3qZbTF41iYSpnmDxabhzEQc
XJVo8XhdvuM7OyPmZFc/Yx2tVD1Z3OXjC9JFb1pOv0/b/K+Ye2/GGioDweInma7HgPnRfs9kCCbT
I0i+e3Jn1n+tpwjbV3kIJGkqSaG8jS2037UdImmKKewe0vg4s3p528UIhu96SVMcKn9mmvMFZEsF
pY6T6XQ+YIXQIbjTsMEMUJKkydP2rkw2t6MR5xFLv9XXOOy+Qah5jzkEKYH9YXlJn9QijTMi0qaX
RIqSyjdfZhrVBhSkiozSHa7Ddmqnb0TOJiz/nkLnyfCtszYbBrmWgBuOGGsfhAayjTxbpUrVfZ54
0waluJybfDJqhpY0y+HWpKRyOs1sGRgcQ/i2aLs1BOUI/EFfLzq7KoyaWEGp+sjGOljh5Get0DPN
JJ5WJotWrGJ0XN9NIvd5kdJPli4gmf6qmhuWJ1zF8NNc7CDFCsFAxwZVwgccQTfJwwpeZDY1hfOy
6SmFFemCkkCiCQ3VZN0bCaawhw7RRSvXPTFs7Z9dD/8vHoSXoIAvdAPgyvku77bjnBi3EQU/Z9Nh
OgOZ4C5qXvuSA0PPv+lVaXnBLcnb1a5S2j8ZeuxmiUf1NKyxO1npeiukGROjcmem7/IaNI3QDw7L
HJL82VZdb7i1PKA9Vu6++dPLVs+wZ+P33JHNFf3slsyuXPJy4JboLOE1TgNMSWsEbWwtvhkAUHi3
x6zNBrDFG6BvIwE0xE9iE8QC9BCcHtkz68RIwFURjTYcZ1jBb0scYbX8mJHbBPgChOL3jPcE93ac
XWnDk4RnfqSUuPGm1qxJgAapNMXBdMEbNeZR1UD76cftGOkP3ma5aFZNYrxRyKSkMtGLz5OhDZrf
y4cUpUcPNFZJQlTN8L+2rx9t1tG/AnY+XYAPWnu2fFGp9w/TplD6jYZHk4pEI31H1JH93VjtWitf
n63FCDgB9soG2zCXvseFA8FgdcXDwrBHvbYUB2T/YTbaK19MrtmLXSdqWuWzJvX8bpLitcnZ69cp
Kug81k0SiF2Kf57c77QQMa8jloWHQoTDR3K0IYOz5Ukwan2PGrmg6bpsG5qbmEpqZz0xcesuWcAO
bzxqHrzuQHy8IeS6w4DMaAqECzF/OsmmK9MhNpDdbQmiOGYV2fOlV0NnAojt0mGkBaBGv+8CXxjL
8mQSgj0EruwNHTQTrEc11qJDLGlDZCqFDdvkpziHzuRkiMxZQ+WtmGHnnS4MZl7qGMuZLdypG4YU
RivGnX4+yLTGwTZnG3ijGgxtB5sfwj4F7lk/qgBlO0IvLOK4M3rQknDJoSmvbqfbAAsn1Nxn8meG
Sf5Th08dsrNaCqnZ/4t+ht52TXA2mbcs6o/WJn32/hqieMl05uKbTWGpQBMWkagwaFX23oFnaruK
SCxMP0RBM6Ex1VdJc15HievypupbFWHolyYnz1G3EcEnd5OA8xQ+q3RTPDT8+hE9S16x0us8Fg0c
t5isSl+WC0IGQFDMhSSiJxZf37QG9umKAIO0QlOlaLtGEqdx1mcO8PrxodCPRqaosiX9DUpHiqSy
UAweemHL94OdJAkp/WV3zW7ezeI1nt5TQ6sumUFnS/WAvYmFuUdcbkpAJiL2MLYLCfpI9SFcPcoe
VE1cb5Wvd4oaTJLqZt7BRte49WDx4GpDbNlbjToNuDtvIeFdhLVsHkB+PNzKQSdmgWzfpnFsRrhD
kZL2AyW9SpPd/0H6pE86cq7RxqImRuO7RSyU5n8gfa9PY01KEDIYxs5C8wJX+0syRswI3XwwNuBW
IZnncBoa1pP+laBgvhdTHOgzwOAQa/UIYzKUcnfN9bvrWG7+l5moOJVqOcye0RrvZBMlTm4qJiP2
HqL6qrdlQUoCsqqGjfXocAEMnrcryFrzCExqC9FF8qXX6pQMhQ7oBIQ2DuZyVS8Qy/DtgHdJX4B7
UZ9WCVSdmLxP9e4cF0l50pVSlasibvRjo/PNKLSPNJWWSAYen5Z3Fm6gpGkLz52I/kVxvEHQtDxL
Cpf4OQvCEpxysEniQMYVvZzl+cFtogKkxp3UOngVFfTJlLPQBwIkPxzC4V7GDMDXqz2QttrHUMG/
7pVlPf3pFf+D3GjIlsVdlRNk4v2jkVxExYFKU0sQ/Yfryan2dofR8WZzUeztanxQWJOjoUBOSck4
4Z5ho+OS9KzZDcssgTyoYNzAbZDXDkId5+P5G4JPF2H3bQOlFHYfVUN5qMHJ2ssxTiZzRMTKYmEM
QWnoTLqalCgmYPkXXOjOCPdTIxplE5mzqfGz/IgdQnwkqREEwSmOO2y0/I5SnMPlIEVCuz5sdpU+
cByON4tkuoSvOLsM7wf60whg434RFkCdWRPAyIinVuNQ7ykhP2opYBaOWgPl9wAZSjXqpQZhNCiS
PAzlPWVRyzDQORfmx1iT1tDhbdpnDGErIPeA02I2jKlRw9a0wcVY4enPWMjcpnwFSWKHekxmJFeg
0IYtCbwv4thB2i41o/Dmw9U6qxWgCnJqcWqvPqxFRk6rjO//rjeLdP32LMQmUKWHdqfQX693dIBo
d7rjyGcg6mriavJ29QVH1Kbov6HFNyHbZ5BkosjARXBwE+H/2pRP4AV1q3Ft/AUrwmt3XkzODeax
xWIi0MjFfnekcayF+arKnyV6DOK4mr44RjQq3L4pGUSn5ntLtoA7hpA0hB4h59OOTvJWVldFhG7n
AC3m/j5NKNfvWBDXQTqHHJetJSzdQ2QO0SeZWqj03P44k2CwAV/J/0Dgk7q9UEOwE+NTGpQRm0mx
ftBY8CWtyXfujmVFrIMosIgBEP4UmePqcqwlP4zOWuwZJgEEg3vYGG/4Y7OfxyjF2Ac7MXOlSAnp
re557JSlGMnVA35eX9ZLuRNyE4a4cWXnJ3E9nh65bE/btlWMzH24WW2bv61R0nX14HXERksNIsBC
GUJXuGhXYBaGjH/VQMTv3feEbnstjm2HOfhziJceCbhMmsf5keAg8o8TSQDdIGAWy/WFZgp+NQZo
awlmpp2zKyG0odnjHY/NrwDxWiwZFxdjQ/XMOWDnNuo1Sn/qFEYZJNuyKCGe8AyjvcARKzrF+7yj
22j0QqaEPQOz+ud6XwP1tp3fkqLw6yJfEBNIDDlkJyVuC37S+t+gwK1o8KCoxa+6fqFfru/uMR5V
iAXfOAAt6YJ4xN5KFGvRbrOFG0nVLANsrDPfwTsAMfmwUItziGCnVnMwQl5cT+fCjPbVofInk7sI
9+DDk0ia2gAAcR6PxwqfS0sTThZAQJboMvxQiHLEyqruqjJp/Ji/4yu81blTKTCvaqlzFT7gv887
Razr5KYHbIH0JnafNumDMpBJpfkgkMAHUJ7IrtdTMmstT+ABFuI7OGMrMkNffoLnC523o9Jvf4Fu
gFUDoNrsuHaSs/m9UjCgmFhNPHXIV70qKSFGyqDbWJhZCanU3xn+mgWjtEW4upAiGaLQVL8BCxGO
clXQLEEk0QqaJ/F+eReIJNPA90HyT+GMKJxxuFHDTS7G4v0psi/HrRInTaH5g8XEuSMXQQpz4fU+
NTL8u6tj0sdJuDlRLu7HGcflfhXRXJMN3a/5oX9UAIvoyfNXwSniiFRpYWQMvxoOxZjOr5m5cfKX
7l8jqqQR5CwjEdW0LDLgrmlioaRyhPnKcU0yc5YDQcmtvo3M94zCBu7coRZYvJLUFXgktVfvrKdp
19siFdgEJKcAcm6MNmxvj0vZhj8sVCZnyOskYgDCPMhZcmEhfmFeh27MkQ0H+dcYU7QYEexvesks
71Ejt11xTD4s9iyhNhDqCX2ETpc5ckHlAtJYwnITI2XmhDDFSn2tw7jkQf8j87OWr3ahg4TR0xdf
fRbgJP+FxTBXE3cywmnf1PZP95aIRPYWbfOgviKfQdb9kf6BFr5w2agvPhPzG8w6ZKN/p0pFqCgJ
zHwdUtmILZIWwy4sMEdUotjCHvm/L3erhcomn6YrI7eWutDzGI7jeAjizsgcDfCtAREm/QaQdatv
jStK3WRz23b87zeumWUiI100gXidA/uMrItqLxmof2ztYmnuXwW/R95RI/vZzt3YBLjybt5p9D4B
ET7zJjlfZvBwaOnDrJKeKTHtIHcP6+0iVft5b4ECqkZzCztaRf6zAAbW4CDWMflkEOFlfcwNEoW/
dU76TLL83yYzE7RmxLuVqihRpoEsNvf0Qb2jwu1+o6Iw/A5dW1O0U32Df6f8kJBNExWN9TDCPH2O
bdWtJTl47CrT7ry6i8BXh3omPQApzz8ssil41GnAWXqMUieZwRoSaSP+inkgSPx82nW3VRWN1Vgd
dfWal0pkQ3lfE2iNSWX9opn9CJM74Id1V9VTKYniqP9v3ysjW7Zkc/PSV6q7DF23zqNKlOVYdZWy
hirpOjGqkUrWXffe70dd2RdZOE1bWP0zKw8H+dH10KUatLHUHZZFRj7/PrzFEzxLGXFzhxTtDY3t
lEo9DJx7x7vZ2xZ8r64uov/9fqft0rXecCFXqay92T1dGnl4KdzrWsJQ0gImWLouHdjQASpnjFQt
xxbjz8/AlTNc9ZpW0+Y8yepDjkxIj/t5lK/TYAjEn0V3qS689q6Qy4TgiaivC2erXxJG8Kj5omIH
0GSAFRcI7BQF9triFgeIeQuIR9Uj32sLQGOmsBsdmifbl2J6uCL+6+dfpwMTeqmqTtyECnpJTagz
GwT4EzopMipgsg4UckrU1vxVNo+jQsh/KZQb4rL5wRIHvUn8jpcO9AXf1zfZzmclDQ/oFw78sHlr
mhSkZkGJ6NGwAlaYJs2M2gRBlp0K+TuxBRkD/rxsMcTj//fBrM2FSPkYSX/aPTyzymmu/DvTTclJ
qlvidZBIy6khOmDN7EY5kwbbrhE6Mibbyv0oOWcSOl5KHDTtzIfkjlhRrPvXK00uVCzKrYQxmGk/
Vc9KYLAjalNjWUS36ZOXkOJ/i0E+1w1oauxkATOuxGIXtmRjonKOe0VQxVjsGOYWl/9mOC3ftTo/
6Gbtn1+wuFuD01jsBExttgN3pCIr7qxPEdvQEUYq6JOrb2Fq0sSIkQ+c7A5lyv0lifRG+Txx5tkz
CoPC+ozPdWqRzvkrqjqmIFXmwQszJSp+BkDSFgQe+oPjyIVZD5goUP+xrNB3SonmTfErl0IBaxga
rUSbzlxU6j4hnRTwMyvaTgxmo2kwAL9vmtJVwg3PC+Hmi5Bqmc7HH6VN+KV6Z1az4ICWCIcX5NRl
ClWeUt3/QRfgXuVoUWkGBgz+vAz4ZYK6P4H8CVd6HEiKSvGyscOmqMTkUmZro/V5t4yf7Q4nEOzD
4TGPySlwG60+zVMiw57y/XPjUmRXn3em9uluYA1nrxy0bPIH/hwNKClVL06Y/Y5cN9dhfbzsEl1i
VSe9KnySqtSpp3tEpMy5IXuUkIFgNxoXUwMpPjrcBp8IszFbpSYp3SUYjOV8GpigArKwQB/OM2V8
9EX4NO+CYrmfpe/67E6DaqzWonJZsDqeIixsfn4cmKX2CBoGG2X2yBrbpnVmcRkv3vkmCF4P1BSF
j/JU+p6HoibYYhgGYoXdaH0gIxU3YI/FujpfDRi82jGC6ju46Jm/aDJ8wKmY3AwG78KOj4NFH+y6
F5Z3+HjG4LoHmdS+0T8OEflwTdXhSXPwhxo5bsD8GrioKrzMRL++JN+QEm+UnzYxZ7qm2m+AiIy8
+8ODpDEdufooRLL4ZTAwGMfuEz7+kNd0fc7GgxdaK6LoaTJb4TwivsIsZgTgrO8E2S8Djve1EU58
B4G1dvHiW/2PZ1ZYuJsg07sehZro0RBkbbOVcBv5h8Q8aD51t55UuHKtqVOj28Nidf4hVoVD0rSQ
0om9NG66p5r+e451Hcb5VRkMlaKiFHSSEC+QCMWnyk9jdSe8IduOrOVlAPtfRTvX50OAel/+27qU
KVwhV5E5ojB3iJguPp4L4sPQX5SK3rv2CDOHL6GeFriUAS7VJpaj5eVNzF7okNMhhrvwgSnI8b/w
e3Q7jabPjz/Zg2E47Fi/4Z4clqmLSBhVZ6dPCetZ4Vmlvtc7th/0pSqbHKSdxjwQNciaxXIWwpmp
2+DxaC8kv77cJ91etOHGxDka/Vkjx5h1CcFvSYZ8s6TVpMcELMMEVjaUZG2QReZWH5SESbr+MtrY
JC8Za/UmsA66b5sZVH3HMNVno2RNw7kCrpYO0LMIA7AekyVUX/+odgDYfHI6FIU60X6MFfM/Rl0g
sCWrcCsQyoZELwm0cbNodyD/Ti7fmP1SCixaRYJLVsXlzKZT8m7COl1eDebEZ5OUbpNrUrC6FNmG
iZR8+XGE+WqoZg3V0LH2k6rDoyY5qgYIBFLfBv/bYdMWxuRl3jQ5QuJD6X/1ILRkIr+2CL5KCD01
gp4eyqYEMdXbWoZX/u4fjwBBQsnq0/4KjKfJGYPi41EnO+oesahYfyTh3h9jg8WY3vf65tYsLRCX
Q1sPrPcTicOj7mdhn574Nwh4obUbS8YnG0nnCQQsqq6JmW96Jn12UWdT91aUNQNSQvTueUo69R2X
taaiyljSIhvJKDyfNHpCoV+YPHzhMZsBo94B5qDY5Vvu8k2l9fKw0OcrOaP9/rfaVtR8uR2uX2Kt
mV/Oc9nS9ODzlNuKPzBDJydwV1W8FV14vWTg4UeUUuvm1dzInUrKuNIoHrqeBr6+0VLQWwzCmzYv
ZRhmvBIMp+0ozs3ruyEhhYPd4LQ6hGL5hgZenfOIPMMXCUdQ7+cLhhd6+11TREO2ZOQwGXqVQCBf
BHobO27dCI4iq4sP3nesfGp929J3lCEsSJJwBtsQ0ZxbT248IizvM23oais/o7ZgnjKMNkbEPord
pLwH/3mw7oG55Y8t7nyEgy9gAAEX/zuM6n0zB3VpFbgn4PIH5t9sEbBblqmgS4qRhB28SJT+mIqP
Jl7cM5Mqurt5MlawoPdAwa5cpjD9Y3a3vpKr8X10iAOK+x5WRr9LgPF47LluGeVPsyA2AX+x1n1/
0dV51ll2m6/yULMQBh653kTHiXFcHAyS5/mm6pL5MZYVuOEfBpadF12gGdW+eqhwOtxvNGo5uRty
VSppg4EMkZ/tFnU7orsyr5SGs4dDsNixOI5PXmq541hTU/F+oo+9JZAhUXmGev/6CADAcBJLx3yW
a8zD4AOacAr7Oqt0+GGLBT/2c1ndsLTn/gjfaUMN+GXCIhe8AWTOb6XXcBIMQGqgBknEppcmRHLl
T0aq1pZ75NCzI6m1CqPh70Ihh7M1ys82GCmDPjR+FtwvujTMPNc9OjW1Ql6Q7npOcMQpqlxzRg+N
ldArtdzmYuNxJuTAHeDxkhCFhNJeD/okqUBNbVpdHf8Y70Bf1PUiWTelal4pA4ghYyukb1Q2UHBT
Ix8zLszK0b0qGxnFGu9te6J+KF/mYU95Iae2jMvs/TVFfNXC0si1F8gu6ef8uA26whfx1xiIaoLc
I6c0RiuD3DwtYhYp7J0rIEEroO9os8kqCjORxcDDhS5lD74lYQAZeoA1C8vBvuF0DLuumuv4JnCc
VvJ267R7raPszd6mO/PrkhbPqMFKqj4h7UApAulKW5c8cRIqm2LnLFmWhJPlWqlDYonp4UkDhvB+
PNK0APSPSVLi8OuhhEIIIRGJlWnvin1C/cntQPW3wgp3VrKOp5obEQgkXIFYhMHeDAiYufM4fsHx
wImiTZIdSQdncL9sIgHMh02NFIVS9xGkmRDUa/23RWdDOMXzOUsDANH01AjCSmvkruk1+PuF+/Q6
qKdEO0wcgETrVqee/oKXNKfqRNMkXATNqppBUzKMISAP6j6qN16uKtWs8JacbfUX+UrvBSAUX0/z
bEVLwz1rYeTVOlB1erlqEX9JDbq53MWQg4TCBxVxOHS/Wn5QVR5mhyAcwkSdUtFM1wOb/b6ftFrD
R81ANM+Wikvu6laPUybtSRKv38B3X3C4YUC2w1Tdd/v0GXOzRCm48aUg1u1f7chaxS1Pwc5RLsHy
ewou5B6e8I6//hlVvaW6ZZ0uwk3qC828VJmnU5R3tVWAveygf2SIWN7386t+2hcQVT3tCnIOGY7v
UuhQ7QZ4gfN5H1WazaOVWKL7WLaNDd1bKTFwT3sWi+eMNW8Jk4nHWybKGGgKGUzMo9/32vao9lP/
ap75tdBVUogbvGFbBkh1xDSKF/9tI9cQf5hloCekNtIdMxvg99hQoWLENoyQtgw8g7zmL62HicZe
3gcuw9JL4kFHqqsOWMPJCQ60nmixK29gudIxjZcGSFPmngS81CR2ZzD4Tuc7l0qLhS/7JWKDlstd
9zV1o7+BpSIsqIHV0OT1yUivWr7o7MaVi8ESDSEqpqpviuxx4uy5/sq70zPnvqqD8XE3PFxt8osa
20QlLYorLLDyUeHgfp672gdCUsgMpZyPLW38O9SasFs2AOjUPL7W8cgdmZ2JNauQwdnsJpCBlbIK
5+KaGNZ2zkV+DQJbh4lvmC76/repDdnRefCiuuMJr8kQNf2liAUOW1DcZweH3M/qpJsxq3G8i7dh
1GoYKYjNeIlWuGiLW02NKyDMP2oDNHa5D/OXWZ/Uk2wgWk0J8ecq380/e/YuZ1lKMgkH+8DHccJP
Ei0+Mb3eKYCh+KnJEaw4ki6kZUwrcF9zj1+nlzFokGxAYCBryXwfyFe821UET6rRqwTLJFJrKg0/
oNKw/40/wL7Ap3wzerMnQT+ExoszAkeF7bWKDkMuuFlJxUNazvTlQO3IvKBfil496tPSsLqMiEbJ
P4S3mqOaKkfYh0ybWOKFyEbxKEfqhCPALgPZggY5NXxqkbHFSypnglza7W8ljfu/mtum/VNPjaLu
zSLGVYyjKOouMhtkDKqNwIDXliCIQDaaho9SvdxjgvYAWK0ujhgjldpevN0wgbSkAqmXtaIBR1+t
wsXI2nmSp/zIkL/tuZvyToa3Ct1azPEsJmR1YvkJ9P4B+FHXvIwgWcHoCIQc9iyXi2z2H7id1W7C
kNvHA2sTJQBcRGBs4BzUsiOzefPN25qgLpxijrdmsYuhDWP063XyjgFlumiaO2NLS59+LhQmplsU
iHsvxehzupbGP55T0EOHYJRyefV1J4avVHAdjimOkkAo8ESvWYe7+CcWgT2/VCeupFlxE/tUs0r8
98fC08V7/PeWoKlB5L1s49pHkXRy4/L59XcgM5bW3FIDuAaEtQAFOIFQM3Tf9xHI3Quio/OjxuRI
xbxhxYSSWWIw/SuVjEq7W2y7wxC3VLMtirs6fPsMRBP/bvvR8aj/lFtikqM2JR9h1CTuKINBCewu
SVedjv/WZ/INJsbEy/yVtmUpWydEblcFbjmd8n/Bx9NtCi3FG0fCXILQfzPfCa0TIj3V6/vOplr0
IMw8oVo62S7VYkXaEhPlmCxGKX3wi0Sp2kTDE97C5Jo8G//Qbk5jgz2o7N3r8AtfKkuy/sIf5LoK
9p96ng8+0jzSUxeL8g0V1DLvZiLgdDeJM3GDjHP6UdBl9pkwRpKydeqDownVmVtbdgkeUhpGqWMg
MkaAOVsn7RemquC4podw19SsxXnPRAvQ//bP/8Co/nSRzN1I40FlZO05paLHZ60Nqk3W2UwfWUOg
Hu4o4h7Idf9WWqcF0zlKEZfRiOLve7IS9qZlC8zxXFbPzkHT7nC5xZFkqF8ykGTGvDLsnaQCkSui
H0rHdkTH4OHNgFgXSrO2IUzs7SAwIS2Ta8BzPQz1lkRoJDwUIymPLCKYStxFhJgr8LooCCe14cys
SI/XS3g2+vc3ZI4R6I7YWYR8ztquc1CY9Sv5Uha7RvnMAUkeMnFMnUI3qTFQSlDE42qAW9XJKqKX
qFRWHaQAiiGPDDwTS8ZeZLFF7/MlHWDfxODj4g4wrD4YMa+T8Tj1d7bF6ult/5uCmw2YuWsBMCoy
muIomsXfdkgU0KpIqyFMjbxFVE8b+eEAhN39E6JlxapWqxcG+W2aDnIkUfabyWPwxlM+kFNW3CWV
38PWV9Utm7E3hTthOh5qvX3aUVZF8ofn3Bra4dCOK6bb0gizFyr5stg4v7tT+m1iL8vFJs+fHweO
9crtqeSRst2UTKEFrfNlB7XjEdZmTvd6cVPfR1Fti+Ya07KnWiO/cNXsHVjf2UMpGlwsrN4bu/XK
6rDSoBF1WkVoEuu4ElLXT6ztmZgAIbiq89fieVpNe7v5tXiTNU3S7B/ilseTCmOddmVWX3o61TFr
sFHCXQ7A/N9yzZxvZIijkRkyUu0nB/dPlCk/G6/YqcLqUB1HCxydw4OqdTmBfvIo4NHhfAwksxgu
8oj5IRZ18IjQ3dBYuE6XbZWieM22W+V9DuKCFAy9TGrhmJnVOj4/8fgIZ5Jj42V4Jl++Bmlkfqjt
PNScYkNiScsgJuF42AbKLSntSIDAV3Xtv4znTLJPa54HrKXzq2Qdh1kYKFzrGxoIgwbREqC0upyX
t29DVfD6l/afbzhKsCtp8QLmL4V5ZyPLA0Z2YA/uRMC1zPsM8fwZtUA8AetxlP6LuvpKHaw6/BrS
n26Ai7rRt/J/LNhp+OwXC8Mnhw1kErdqJGeehlnJKg8L4Mkq+m/WZYQz2DrdKZuivgo3gCIXRx3X
QmSVyj681/wqctBgv8lBPj0adfsCPVtW1CZrY9Oxee6RmDIuhw28l2yAKxnjp7V1JZztNk7/NBoU
EWrrTABxxMM2l9RnObM38JiD2VnGsA0z1xdoFXbnLQNcMF6uRt7NJlaxPT/BSHQ53jJrmcDrYAnk
yf5LotkZoZJWiyO7NoHnWN4qSue7xKeXwgc2qrN4Awllrlde4TO2aUliXR08475DMlu8eldJERVu
rr3KpHy69ATiL59f24qz3e29YwgUYryOzrAo1f9hNpHb/V0mzfSQRbAt3T1o5VqUFMMoOZ7gFhiP
a7TDQExJ2kIlLikSuvepwg0Q+U7Lo6XcuXvKJLueiuAz0N8i6WSY2vZlyR+ffMrZ8WviCMILEApB
gqDgUgUvZXH1aRBBBg48bhT3yCljyF3eCK4RcPI0cBwbOixwcbFJdloIhlNmls4JFiEKAzyZh59B
WS9uD6wdSKCa7UKCQyiajR06fIIpEtz61somSeumP2F9hGIoUzrh3n5tXW9Kh9pzIdSLaO2XUHOX
dnSfcgxCTSb++7R2A+fc7QvT/Ai+QTNEuTXtpvwKf+2OuWFrWqXxRj45F4EWQhJtQb9bq5+cua2v
EfEXgbXrUYUfCwtCg2sA+xvS1MQJRjDlQH63d9sbmnuo1UPN6v8Fv6kOFrnrIJDrWVGrzVMNjUiB
6zcwg+zB3Rs0wE8jdiN0ykRDY85QLHi83E7sw//rI/exdTI0RS+YB2eQzqWwrZCX7hi/ralU9pqV
QHWibiY/zg9m0ob42Ywpk+rsI+vTKOIxl+VrNC4Memtg0CAhi9QIMvnj9ClSaqmRdFmsIaFyQt0O
O+4Mh8UkBnnQ8Iz5ZrSLF5IDXsoo1616UqPGmQpQ40GyOS3RQDru5Lb2pYwsSUzyaHgLZclPja2O
xMKw0RRWL/BXdMOJ/bWf2HYf0hOvLjcp4CMAwB7HJqlgBGMIsTHamRtBHqc3c5wRv6whiUApEAul
21rMvJ1BuBFx/YkXPbQgkug7IHZlH5RQCAZAiwCbDL7ukGDOVpg8gDhYEcZL7UmBB+pOzLH3AAQ8
O8+WIyCbY00UFEXeLc602Am2krfh7CbZ12MonBaYkNwTTREVq7TRA1pyWeXS7P1fe1844x5hN7B/
LkawkhjgKZsd4IwVQBO/A6Z/Au0aa3S7YUMN6HwE0BsQ53HLaTteDRfOPJaW7lDhd5BeFoAxm02O
JRUuvedOGr9/S2lu8qxxe1rY7g8BaN/p2jrLA3ddfQtvFCOx9lRE8vJ7xT7HAo0fKyNAp3jkqWrU
Myf/EIF9P7uKX4sQGzMAd6McCYeUyxSZJ9DL1zPacsQlAyxfg7neDQksF2P1McmYh+uPa7hoWKSS
6azQBeeAlshVoXa64NGFtxAw2Nyf/EXajU99RxMlTEwvuAczG2WkpNYS30+X3ynx/W1M8MpY7Z/S
YQsYv1f6ayx2Ovi+Vpp2+zVP1ci05PJ2M481Dgk6CQ+lexwzBm62vKwIK6+K1gJEJZLCS2yhas9F
+EsWM3t78XqBaqTEZbVMI7QGhZ+hIX8s+T38d9RwARrYrX4HwnwS0wl0t7FMJ9okP+we6/5NuEYB
VD4PjumfOvprjmwF3H5AdTuMdNnEt0jZq9Wv7z3zQZJi/kgzvriBBioNWmh0BLSXv3oxgwxVif8j
yo2ZLdtnTodmOPs1E4GdwbYerNw1s51hOijBUvbjRi1/ZC5czfwK1IOEcqOAX+mQnhrsSno4RU3H
51gJhhlhB5nVETAh2m2H3wwphmb0rBQEDFRqGE93DT1yVKWLXLKxP9Nq9tcpYUboAXjXsi8zMeyz
GKH5trmo8duXvVWJmqQzo2qYm8wxg5kUCy/EwaxdwHSENcvMnKojLhzvGJ3IPEzYZCa9L3vhx/jh
9lCervMegpwaMKw3idsQw26YCb+Cq2Jb+scciWqeuuZk97GhHVR2Pne4BkoOwv0yZo2AMNBveJ6L
BTwYKf/vFborbAbkVaVL2XOzxGyh1EQqhkNuSlZFCOReeQ2ubzwZXt+cJS1yYF3AgimNanDRprOr
ucUXXZonFyvzzdv7EtEaC8kHFeKSJ/1ppxS4MwbhnSYiAEHO6rT9Q4hZFpFmSt1F5C30omf2wJ/m
9YNaLBilLuZEzm4Y7YfFWVKNbvjEIjT/2J6T6Nwb91qtUJz1SEEROvZ4lw+iSmn4eBcDz7CENelM
rDePoworKmHo6cCVD2tWuL4j6awAramy3LJqaW0PpvJ52H6gINx50IGYrgAaLTG217VK83H3AVn6
v0fdkFYQZ9kxekX412Ex3qVS5ojpXWa3FQt8Y+OcuJ8t+F+10afZBDfiHky1wOZg6GJFhmGJKqhx
MRh2tsLxyQT1TVirnQBwIkUYPMlJe+ZnNy0+qPQJDtbpAelmHrqDev4mLlLa6MAKtUxgTlTR+hsf
rgBzCLnmF8qU32lEVaZu0DxygquUhVm13OlqeqooJ3n4UdW9ZjcajZh5GiqVuZIB/r/euRsGQBOV
GHbqtcADceJaLX62/gQZ42RPGwUP1htgTp/pg/02qDtgPOXJl9PjZoU/CD//nPrFYsBWS5PpctIA
FJIcJUMD3NAZGTq3XzoZ1Lc6wozyBW+bgb87L06TJfPKLQPg2sapdCw40t4BNOZ1hgXnuugxFmW2
FS15moznRVI7abw5KPxT35UVDEVg8XDH0A+z+0p+ZCNrNl3MGJEo6+heKTxYGitnJDk1GI1JKBoY
66hhgt4nk7ffYwXh2dOBOPCrx55dZGRK/6ZjZrXWqLD2aWX3rp1Q74j05xkT6rk/pf2nOKz4gOQR
mLM+9xsUF9nOZF19kdQCovTEcHA8juOCaAKUs52YYKgd9Ifjt+FDohAiqlyrP2w7z8Je5lWjTCmk
pTDc+L9OOpVbHwlD5GF3FyRzmjfQmqqPxYgVFaeglYvULyNPy/XEiYGhCI8034R20ZlIPEwh8VSD
2iQY5o+8Fr9TG9/KZkpqvIZjYqcfrTdZw/1VvWwfdtEIoDbG6E+2esm9uzxbOzb3DWNTdWOTOGjA
fyhBqpQnObZ2gPBWPaRQYBp149yLKb6okIkjh2wFbyYrOqw1iN6WlKkOgxA4QH5Ezbs3OA21bs6U
SgebkJLfyeyDcPiW3YZU7/BCAnO/t0eVWNkJxt++LEVrVqgniLxr8mx2UpOHYa2piczV/rQZgrAI
Pgcvjmc7i8BQsWQ5NzsBLHS7HTwxo6IMW9pbNY+Ux0BCmoTbx0sa7KaVocC1etghZ2b/Zf1piI0Q
LBa67v1aVN+lv16dGAA46oYIjT1OkYahCQCbVuaPj7M6EYEzawqeiONMeZtN35vdqZIF2zny7vM3
nH52rPSTBxihyANd/Fdrcj+pr18FLfathV3IfKyYJWThqe5K67QfJe8oSg7cp5cON+VHyXk4gUP5
3a8jOb4Fn+iuVjb8w59N/MuQtF+QSLw4n6oxZJ+CuHoh23hM9gb7nWRSX6YI5iMK4rO97139D1hj
clJEk5CJ6t7LJrGLTimVpuYnm3xFM2gzhFBAHFEnZYWmHzR2O84Nvi+g9A9DI+BhQ/QLEHKfKoMH
g99oaTvrL28Lj2m1UuMhjSmJv/rZkltVLSG5aKN03QUXGuEuUGIPW4Qq3xdLqGP+EFx8S4Y8s1YM
HmCoG5d3wP+RIay7VF77u4rwfWQIVUv4PqfdJ5hmBJDi4a/ye+KrG2bBaiKVwniN6wmg48q7DN4n
QTbPLYI5q1L5MSr7ojL3L3kSkfWCscVn7EuybcF15PCYb5pFRqsjiriU9sNU/oFt/wIW5JNedE7V
0SxP6jtbQYFPxVz/oaPJpjP/PxhK29RF7j+gUzqQnf8TbVydEsR80QOFDl9pGrzXBstg0K5kr85G
VDR4OXIJ6BE44pnqUMW622lJo5L1yr87n2lKUD77v4tKyAik8DrxknM1VAigRSvIqBI8DsQkr+IB
qrhnY6if5McCB3ueBBuvb8wHcnykcuCwhiga4rEagTx0to8prO4IVWoVSbSnLOLIJPZpi6uBjCiA
DQJekX+lYOYpdRIfe6G/Js7i2I+blIKUGlS7ifB4rX9+cGuexAPVcAHypRNh+vIPl4sdO/oJyJcu
hUDmQavqN3WVEf3mLKkAqEsxcjj3bWXDA51xEvYGPCB25pSjePhLwQkOuDnoyAFu2CHw05FtQX7h
7BDVgGPLNIhuAajgFE6/fcGmzJB1gM117WtgeeYgTnghc3eM9s0PLLBNEoB+KyXKwr6gvN+DCc10
VUIERxQZY1F4bP+NjiX4sCehllbqZ/34XI1UGgO9T21flRvqwv7+TAzoseNLZUYQJkWh0J6pxU07
Cg4TzZsLVXmB9qUOaC6204zIaFSC2UJ3S9yINnx1JV/XnudgVCuB3YDUCbqY6jXzpICQ/YRYlOOo
8NlTeGrc4Z9z9/dxakSCAiAsw2bWSeWzKTmT6aECJy4LqJCKPUk/f0q+gW3eYKswBZdqrTkNW7bW
7Tp1zt8FGvX3qrJdeI+lfVlT+B8KgZx8Gz4yMbX0hZk0ItbVaPlvdKkrOuDTu9G924E7YVL/Hl28
/M5pc5K7m2d8JbydwW4jT+5zJZfxEOuN81oZIZN3zUbaUbtuXogy3sFJaH5ey8jWqmWlCRM+S4Sn
olRYrgIDf2Z3Zbb/ej/FwDz5AeU/eAFLaI0j5ot2f/M4HsFfzmGiEC+Ivp5XVGpZDf6hLbhYiGF0
4Y+aqM8RAFWfolCYe1InxoixYow6DkbceFREqtjwblQ1xiAC6QUPAvfp7SMpbyJTef55Hs/8mC35
7DiFlj+ICSrL5/BUN4mmgmguJc5YTy8pJYviD+1w1QWFet7IMXpGewrcdjbixLmGFAH+gFdGxGko
wDK7Kriz8ttGhj1bWsNbHv5FD4dLeeACmDrWUHRQeHn727P7OlQjV/nAR6R1Id99/R9YXhQmFSfO
4oqrayAp3Ir0EFM2LfKAdWoC1Objy4Ve08nOXoRX6kAtdbaLNOFPWTvJgqkOIkpxm8qtYqzfcBcB
ln92ZnJfgYKigpN4vSArI27haWJsB6IL273mMj58fvurUJE8wnKVFnf1xniLG/Iay43so91Wi+WQ
cPp3F2g/vVnRYu7FbGnXyuIUBhZAb6cAjrz0FEjFp98CxGsL6f6MZxpdBrOMgbP/gq94DrG602ex
vy4ZJFWgqjYD7BCyLMKzIiiCesT/1GmEqJCi4VDkiXe82gE91ER4Q6+1Qp8Fo4bmGb4Id1uTSrdg
zrhksaQOBjbgCDi0YaIOw7qjDphYR+pn7TNLCJYOrdPyEzh3H6oxSf7Lb1Dh2g271NiFc/cXrEEa
qNMJhWVzGR5LsE+3CdmCGVi8YS6L+ZUfyVoc7poZT4EepLI4Eaa4DNfUhI0DJ/dVTgkvnjziSNoa
zOUrImoD1EmdpXjbLaFCQZ73mET/qmx89lF800+sHkmHrInmp/ewK+cV1+SGGHCpaXPDBZI2UZRo
NcH/ChpygLIh6Od+q2z/QMJlU3DijeaOF3Ug6zqqXSeEu2HsstXvhBXMkvPZNLJpeuSyD7JbXMFr
sFqDJJdnZZQqdXDntvv7pOd/Tt8YppqlEBQyotVsRWaaLP9ZhItZNVf4klypc21UuUHp+AcwWiS1
8IK0QLdT0xiAvwr7IgQXsQR3GHzhS/e7dsgnpeRE5ulWYSLoRauoHXHNLU7xhNQ8T5BoJw17M3GT
ea6rKcMjywxgNE6hRSCmthDkkrIglSlMf6OLk+ACUJCBld6/Mijmp/PrmetDkDtRu73SRmFAm4mc
e1LlB9lQoZJ8O9wz1Vv26uTpFHhslf/uajYQojADxSO1nN0SdVfT0ideq6yvn1VnkivwJ9U1/Dhd
GARB/5h8XAlKeTf50NjR21CZ7L1leZ3YrlQ2fv/jmPy+yn4lpuCwJvJ8Krpz/p0Pzy9vifI4Zygc
kUw89l/yPg/fu/aJkyXvvG2ui1AD69oRtm2eqm1J2VvM63BYNVAf+yu2krGV4wyBPQ1MY0SRcayg
knXNB2isEdaifOXezOBU+eobgBJNfVEDcjLZpEWoXU6iKnqyekk7YPCuBTeN/jGDyijjf06srwri
GvUPE24XvVxFgtkTPEu6u56b9pViiQFqdn4FaRDo8qGp2muOg8jEod1VfFch5sDDvEeEfS7fgsjN
9XOcrBEPvWE2Swv3rbzuHkWYlW8WcqqCIuXYaT0z9FYBdtltht+Exj3T6kTXqhW+Ptkz6HLAX0rN
zhaSM8sS75y73S/qZ9me2tw8WIclt67BgO5Xk9MtkvKD7cP+UlItVrZM3ktQ2KRVz3vr2OEIIp6g
m4MtktZTXQFj/swC/UObKz8BOw1A7sZDb7rEqDMQIakQ0oE+A1gpiTsyhUAhSd+hA+EF61eIT3AI
OMVobLdB/7Tub03NhuzGW4iG+7ufLvbba/Z51iMyMkj4rW7tTU9zeq2x1E6NmTcQ/yxkXv1sYToV
FR30vNVqSbWWmJfgS4fiDzZ8FQpFa5ZObtBGCaMSV6YTEZRMvG6LjzyoL/SVxyfUFP5xj6Rd4YpQ
jqHX6dKLEvFpeAs0LzCiEQIBQgPYG4do8Ii8vc2t2zeK3ks+NCwMzSuSmnRLN9cabwSWIvhtAiL0
eudELx7bZbF1FF0zavYc3Ou6qWy9RdTPuMlHk4RcrF0Uj82/rYsTAks0d7d8ih3KFiNc1LXkJnK+
4W/ZY2kg3qXwmgRx4ybX/SdcwxzGswCO2u7M4Q+l0d6npYOJbLBp/RtL7vmueKoHnGVUA3o5cwtg
dhKfzsHb/Fev11rWeuUEMPuqAvzv8QGvePHAmpzuCQUYZyudaX1xWJ0aMbv+KqMpuluMBx1kJYDU
FtyQBBw6RAhfxOaqkikTis+2MneB+2l6Kz6GOCeNIM/QxlPB/pV6qVutsKng/Ru5TC753iwi5Fcx
EvINzsQzq+L2Vx6rfclRGLjUxnH0gofp2M8Q08ptaPsHNFeRAg8PTTbzpmn4N7dFdICKA3/BSBHS
zaYPbCdGWSDnwpyWGQa2ebVwelUOyStC3dVO1pBXW4R/3b/cmyFo14Y9jNteoRkZFnbStLLkp07t
e+621puPcVLWWG8uDSyKLoShfkGTEypl8X6uVBCGEpF1Z7DWhyLEVpmg6j1YA7g9Hv5mXibX5rSo
wWd6Z0Rf0JzAm+K+TLZNFIwHLze7yPcIXvW/DwIGZf7x2MB5+9SCARwLB1PAch5+60Na5D7j8xAL
okwJ0QY6g+T+7scFROW09sBBxvTjJnNluyr2iHOaWw/vAKNr4yY7EFTKS9TdNoylYxvGVFjODcaI
vEdm9hQ1KzB8c7GIg8HaKToW5K1VueCQjAAnHLi+7m+isoz0Yil/ohJf2uDm7V+Yusn2ggYDmpUY
Jjv4hundmYdO5lpIAdxzzNlF7LBiNadEuxB2ds6FTVXQQxWXTrsDqdD6ydtEtto1PApcMXS0JzKf
EE1Ep0yGynjf8P/WdcuS3Y18xOQpse2nkb4vRplBvONByNK5EYD94dGLqk+2TCSNZ/ys7ZpGSWXy
dVc3qq1me9Jn33SjxdMo5oz4eDTMxJJRGRHlpf5QhYhLFnJLZFQSsFqChKJDMFEHAxpcOM9YsHds
iUXI07r5HV1ZMn9HJC8eTFLb+1m65orxKo+F9INBu4NuWMZWxVFi1kN2eAhEkoxVG2cAfhqG2a4A
U+e96glf4ThNcc+IwYuOuyLLO97eLWl9w6LMKvKr5Lz1Z8Uj56Y0UIXyRZhT2Tt/JgcNPHnepk6y
beQTo7Z434bvmiZvWSzNDcNCWSZPoOVxhcs0jLllrQOpQekQNgJjl7nJcWCQNWXxZRGa+DLJweNK
tgz6xvJ0ITd6bhrJHalFcCby7f+A8M/C/RmaeQbhi9XiEvK49rLXLj5SvrgJ019WnstWZFAUN7XO
B5ABiMzmQ1P3BtZTOMXxtWKR4zXiH19oJtygHdG82QFRjQMivWufAISa5hyAuYluwtufZBq9HxIW
Ca4QE4JiW0Ef+CKEzQTc6OuedPMTcdYFCldbaJsIMg8vq3wLlPwZ6RkWRGibEENE2zFHH30O4vMu
uZ7KVsqtOj830SCw+JHQp2mh9jNSVM/t2C8j4E1MryKf5/r30Ie7KNYiq7Ua7xhG736fP4adcXMv
9r/EOnrEzl8mjBVLnMffkqjv4+KIOUlcSc3RzCYqzzY9jNxFGK6vWiaw9ROLthZPkf/JLORNybHs
Yjh1PvBq4f14Qze1lOC1eqMtI5zDshkImxmydC3XTt0NxnbjTjwZoEgdXyj1R71a36rWVUliwbdj
FfTj/keEYbwAxk4z88TVQqQ5RdMf400acMTdWIfEp/vhrxGd6ZWZUrhsOu1zuL48DIpSKHIbjPIe
MRAYUzHafmDJ5vvSUR7Ji/3OKncwNFEr6n7OtEfd0EzKRPMTISsxUB4NaxXeXHawPt8r0hI5FSo5
iCwMAoiA2Moi8sLi7mXiDq+CDdSP52+zQJgvgf5bpBQ7lzmToksFSg4/qjL21cfh+qQsi67cp9Ug
pNp66lhiXgM54Vd+WzgtMy3DUq66YhxJyUF7ocm6xGWsR0Z+SrYzXuvGdbiqLO8JgzuNo19JQA8l
GhEs38KbPbCeXK58mIi4KqZLDbsCqZGdKQPpNbaxwQooK72wtTUqBH4Xv0aa/j8ppd++HwEPtxj/
V9vvFSPBYOxSHXRXR06lYwJGzW1wDmTpkZyYTv1xOw/Buo9mdta69jlvlFIEoquHXyTEfEGzkVH7
qMCXjGBdUL+OaxBfEpv8xZwJ9CwhKYgEjfrcP3XAcMDXc/1SsShLUOkblfHixxm/ybZHNvgmIkyD
xJfISBvbCGiQohS6r9Mv6jQK+ultPTojw0EA1wue3GDHKpJ6amVFLC29eKrAS5d84wCanKYk+JL1
hJs3/KaDsckhEybLmSF+gxKvwyANR7Mz1CK81o3sSZVMkXq18IxN/Xnv0mmK/n1fbRVXQYSY7HlE
MhBYqsQTZxxorbu0jdU63rPcUaDoyCHyTszKwVRjvbvVv8sKzSXOroxfeW3IOhpOEIqyrFQ+Xxtm
UqoWRpzIKAci7V21QoMEp+6dqzK7w1LAG1LwjjJQqJOHnN6zrjgzVP1zyPaex2Up6Aj1e1M5NIF5
TRjBvQt5gWifc4WbY1TBHFFMIOWL+jk+LgbP/18AQx29041qgxhRLoLGlzdDEHUOWP4sT9xSAuPN
ISlQD100FvpBsbBVfklBOTWWzlbWNTnkJcJ7ZR+sazEj3Da3v7vMTuMujIy+A3LuhYYZHP/aRHQM
GxABOFTxoOu0GefjodgKdP2mYWCv+1mmETjrJqcPmNGLtFKR3LQV/JExBRKWzc5TItBg23+rpi21
Wca+noj/sSxPVIyamchpELcksj0T81t9vzQ+7E4l1HlYSv4Jt6+z9m75YB5dX3f8BOmeZnsO3S0a
mIVSWotcEo2+kwxlMt//JXqHtQaBTDyuERxz1DhwcyCac4dztwq0eyU05EHzFwCLvw/+6u5lJsfG
ho64/SgdNBvpzgvWXumgQy8mQ0DRsBVQReXft1UEkJqZu0KxQIuWmW7sAXijPhjJe2Jg6OeTDYhy
hjR8LfynaOpgFL55idSQBQ412pVdaRwnPdI4J52OLaItQHI4Bkux5zwUw25929E1S6Ql3z9o2c/p
I3dQFNQ/oRthVzKkO4VMpTaPZdOLZPDQX29uWsv4e1vO25xQO/liQlrE5JES+9gbgo+NFhAQyNbr
DZckWQy1Mbsr/FmX607M2cMtSoTRKQlO6RC1GwwcjfslOKNLdl6RpGFOgYQNi1+MZNkUlFvFvXG5
w3GRAxfnxysOXKzyyfA+85tEYhY1OPlDcblqb7IKqCCyvvT1o9ASlM8lKAO0D94jgCD86nuQpb6W
LOqCL6piTrUt59u/1y1C8AQe3PjJ6ODlAneb6P3aAi2B+jyyxtI8ozcmcweqtoCnhT4WrPqodWxR
lJx39YgRgIlMicovMFpbHJvaQ4YZfe3Tq7SqX1rb3isvm7k9MgAd6spAY0XrOjOMUb/4uOQxoCYH
C/+hNqgFsOfKFdLdMCH0aEyegb5hG3Tu2cCI4Z7LNIT6+VnU5uAFp5lA7+nt0f3t03hHEGeN9ojJ
0f5xnUszUM9g0lLPHu1WZ//4TR+PcJpLSRRjxVqkJF9x0kAoJyEPHVIRXDxz7UNBXF0jOXGSAZWB
5LyLX7OysKb1Ow0HU4oKxxkeeFmN2SW0b2xz1K33IlfwP8qVQvhWrisbCHxNsVFkyKcVP3W5Lr0T
8RWLivfK68QB3TGMKJ4IkPObFPgLBvpw3vwG2cJfqNHTjb25HoFC0biHwdnwu/rn9SdKPIWvIaAi
JNfR6BIiaXjtu9jnen+i1THDnq9Yu+BudHk9grBAbXvS8Vu8f9yz6B/lmJCPrAYDo2Zzt83UOYgE
E+MIYBsJKsyiZOTtugdsTG3h+jotej7opoEr/xFAoPoi1YiKaUmvuHO+ZJn9SSKYvV5NE0a8AtpC
G4xRXgdGCD+ZQG6M/rT24YngaQhaQTbEoH6oxlLwZgm1SnulzRyYRCIrjixIBTpIyMjAGGqZftXU
kCyj9cEKLQ4OZ4Xy+WgKPE8xi9pYk3qvdKLlRyEb0VFhz9SEKzqkryUewQTSJoEeE5XsySCp7bof
qNviqZrVZWzRjl5maP9JZPmHmzdzL70RWngWJer75Jd2ZtibdiSjTqrZ3qnp6GIeOU2xSUcniJtO
u2ZQIYI2ThpBXb6H/X+Qw9Sr2UGQGtJwWsDKYK4uE3+FqWVbEngklgv43wlJb+v2EU7n8fnv6i5Y
a4AdKKZrir/coPu5BF4+kemHQyq9NTVhYyZtaIvENp4G5Qp5LSWoOSAoiNkkVZoAc8fkx0qIGGMU
a4/xTt5hbmEPi0/pLfY/hZF7BMkXVEpwoTR7vZRxAnvF5vV3W+fUX/era0kn+uRe5TMhu7VerpD4
repsWDFylupPwhlKZ0NQFoDfkOXDcapgWWZwAwuGd5UF3WmDd1ZX2MTitcGKtk+95ebFd2vNpHXQ
MybaZ2MRLmb9qPB78NvcaaJU9JL54cuNDG1I3Y4y3ChdTFrmlIfJ02FoZegZo9B+xzl1QYa8xjHX
Nr7ZAFr+6yWKh9BtLr5ZTzFD3mshm53S5nUqObWQmf12RQvHbMHBtx5EAS1WAevluzduLo6gr+rf
TFsmFfWtfS6nwevIy/Wux72OwGVh5D+fXHjNaW8EGzwjI0HDpkJaVDooaK8wp1CqNMYaGApzORo0
JTqbvAYWeO0+v2sHhIFOPuaLqZ9BrPAS2kg36uQIYIYEJ5iSGWmSCax1IVFnkqfICmX1cQGdcja2
ZkDytbtuTg+PWNit38/441GEctzBnCkSuW52Fq3xrjw4cZLahSLkV/8Qfw7+S4NxLLdJI0t5smbi
xaDsL8YGFSxqUH1LEDsLBI4NHhkW7VCGv82b9KlL3yl8pmeUbsBJeuswvt6Vv7741amcv76uQ/Ma
wjsjM4qQnAly27+A4Gu5NOE7T39od92lRXcgKQAJuMfYV22POCQ5mOIHQO4+O7s1TlEqD7CWEX83
/6G3GZmWEoXWiEz5cBB1heWOOSYC3bmbOQ2Bn7iNL7NyZDCX6TFCK2Nku2iBWG5hTGUwNwbYA1A+
3U/eFOrdpuQzF3ku8pSUYU3+MA4n3Zhfoh0O+P4tU/C9WiCEM6LG39pkfKo1MztgOXCRPLkerM1k
Bg4s0wV+GZbuKFggdEcgYY89C1chOEFs1xyXRlk7VDnLJqkT6qjyB8tFHQlRrIO4Xw162EK/A01u
v3hkbU4qBP+0WloC55foVWhb54IBhA3PCkpokaXLMrgRmsAIDTmHakeIVkVPszGoLI3sXtrBp2KG
ppXrfkEnPEfV8C19Nk3k5XW5akDDg/+neluYh1IKIarqqHBd5CQen3tlihb3CTzsvaQlAXSFBxIi
Rdu/lPY6oVxh9wBieg1qc71ZCvLrgt7rDzyWkSMWIclZrBdFw+vFP0cIkXYm2dM92z3zm2rdYCXg
HIYlDmt9AJ94qKfE60xJpFWRCsIYpaAopvbqfKKTktMjX9yLsCaiPVRGue24fdkCeFrQ82E8T0SQ
B9PbhohzrHR+6aJbS2dbmcJg4YpUALlZYwGYjHRo03qVDXTBTjz5L+DC/TXckc5ZoMNShZ21WA3X
vQGfg0mmRLowQu26yWM86VqkHtoexdTDN0KYIewGXU/KYAJ0DZp0sK0X1Pz8fERi1MoBBdJLGkO5
1lJ0JibPbN5yfs3D9RaX/AC1DemRZjaFbmE5uG833cSgJuN6xdSmqG26ogZgWLfZUu9fEb35R1Kr
RmhoRjAkaQtWgYkGejiqr5z6Z6FTWbkFvaVik5Dnn6VWUpEQRRMy3I7DYQxe4t1aPLhx7fS8bx97
sNUvmOe8NwRdndTLvwjbyCtqtPpeB/X8U05SaQk8hnVA1Ogs9YERZGU/RXV+IpruSPMs658Hd4Az
PDPj6Wnh74Bwe4mpp5bLXNfWQ05FnskP5SR+DyWhvPVzTXdj8DvS9KgHTgJhKxGPfipl944f4C88
pYovF47bPsXBw4NBnYRaeqc0zHGWdS6j1npXEI/TmX9vxxxl0paU5TpLM2pekReky/edgcUf5ZIJ
6L2poguqxHdItCIwchNyUSAl/yAZBhGHXJozHxPvxlt4ODG9FYiulyyGgU2gePivXlO+hyjrWIJK
tpwudRh5Z2x62cNPaiOo9Tkmgu64donySv38LOw+MN0hdqBm+0DkbzvXOYBbk5bWUrBazWHgIu1k
6UXx+q7cqEZWUVjhjYXX6jOjxjlNEEubPClBBt5XatMtKfsstRmx33zEZ81VutWJCSMvUc+Vas4e
kuilau3a5zt7aWOHSiUlnVvFucM6rimH2h9PUVwCPIm9+UJBhqhl0hsvoAnhfwKju7b2Z/dgVAEq
FBdVV0S4lklRf39ol+QPHCCRxvRZ/LWXmP+ODRqNX4R2cU0DI6SVR8CZHs4ystwNuWKfK9yfRuC8
zqRRyJ9rNj4iPDNV9SWgwSvtlcR6U4yZzDRq+R5GjiOH6d9iX2F6EXLWzqWeSjv6TQl+tU5Qmwyw
TIwQyb1Ng3Xt5wYEA3nkHSO+x36PA2zE9ltTUbskH1mBSatjNBgKkyXeKWvkQxY7OFFZ1ROgPNpq
tlWGWuE6P6ebYN6AEvmCFgy/5Av8g9S2DZZ7uO+Mp1rWuep2kdOdk5h3rAQNKFJkhy0TbYCPmLxl
1yWtW3rg9YlQj0zd/x53PtHgR09FzrGnepuhQjp1VLkpGSXqzM8xRVkNr1Fn6HWpp7VEp5e+7OAy
iBuJNWGq5qFUT4WhN3t+wKy8MjLcQa8u7LroryXQA6yFh8vVRSDljmZNX/6nMJ9U1DYxKcZibL6S
YLMrV90VZZAoT5IlSGAXEJHI+Y6NRKBkZUnzSTefe2ExAfzCbAmhgJ0K2STvxmz5SL6XKjSOudq6
Mk3I47YRNzYsJwrTv9Gfu4VWzqYu5JrmQOfLToKS+wc7uHHvHCNaNGDlG+3YNGQf4Qf7oJoVhKHo
gpjmRaXDaVE64xM1XEupOa6nPTvY+5Rx1TaH+brQmGQbOy8BPiCU8Y8P3SxbCDZaYmRbxQ8YgsXN
Qs3YDAjwG7KpES/RX0oxp59JXXf9NIbgSsZ532NRFcyYfGcCmF+2/AXWFHxAITuVSroDnrW3kRa4
RY2aFQOz/bGBbHOinieMiNIAjA9r3leDUj0dXrcrAOQzqQSviRpVyuTMvGNHHNRDHUFAOL4FJI8O
dSmLLLd5gAYVbpCQtspt/zKvGzDpc38BTl2UcBHo4h9OPabBKOPj4hwrMcTMS4UIW36Q7kZxsuH4
Ip767FdeTIpzxQ3gISBgPAa+yx+Ycj9PC45BGxNGw4gUDJHfW0Zgq8/9mGyzLbz16MZIytAow0lt
Sokl4rYvauIILcDzVyq7RE4pPT9bJji6KgijVq9lxXKUqht0M61Eieclo5dYKPRjVI4zxqn2gmpn
Ux3FEDNDFtHygB+zRusN+6H0xO4w5eSw6Wv/buKaKw123O0GTrr+a/d28VxNUdTQPQknflLKMIo5
LXUV+5oPCcL5ybF6r6spXw0dTeLez4SV4Yu7Hwlb0femXh1E61Ab+ztcV7gMRUWSd2p03VR5rWbQ
mJXGDd0mtk1u0up0tw8GKIV/hti1Aqr9uEMQxBVdZKEk1YXiCV6+pD3j59zUJuHoV01NdxqOjcnJ
W09DzsC/Cp4Tgwurfc9wuof9LqU9c7MwtfNPElWIpMaKw8XlWZJwq/VFgv/ZTlsd1Iyygb2ezAr4
OqklBkhi40zv2itXSOGssareQEx2BP0ZBvB1yxzGIqHXZUx36XEYiPn1QnVX8+RfH9u6cgQEdkQJ
pBn7kKI4HNhPTOTqEJRasKmdThRiQa0xOam09rkQQggD4NIREn9ZJPgOeatHAD7bQzI/TKRkMwtn
Fnuf2xmMZdF4mCSPzLpVNE+mQSM+XDpNE142UD67G9WjUTvBg4h/GNKhTOUxKiP+3rCSJLfddz7y
ZahMYZLydJqjurEnAcoWvuPoEOGGFHcPTbXqPZnh6uh5bZH9+H8rDAyy5mnMTx8lb3JLMzLeA4PI
cYhbNdPhEwyCITGtJb6ac9DehjHMbnrgXPAALItb8yHR536dWb8XmotESXy09S+EbHGU68PHpfw6
LGwCl4R9WMhaCbO8oenzn1KOCu/ibxZjArGBJoiYulcqyv5s4SEPyroMRyn8PNiS2tjXfn2pb8Y0
9lrc9J1LyGc4puR8yvUR/XV0MEjOj4AsPMvdJNuyXOyZSX6HOlJo9d2UbiPRRRIB+sdDi/I2wuww
8W56z3mzguaGTaEAYJD7lDX2o6sPG+hVS1C0RrQENYId3gYMwkDOwY7qEu9+T94qKL6MWF+9HXA4
0CyZVpkMl+WWGtZvw3CSKVODtUcIfSC/xot6E4npDgs+wYJ283inWrk3WdR7PI+8z0feegUtq0iQ
uiL+OXivlCtc60+kK5o9WSncjAbfJ7IXb2J+c9VK9aaQrkDF2NwgsKSnnvgdxdHyBJkaaNWQv2tC
1qEszAx4cFgM5r+zA/azCjspJyfDL/Z3JqPnwYVXBZQ33v+rhmU2MQfgw2OsNGUrmQFX+gyyCXsJ
H3GJFgFfxtvz3TZEvtf6Et60Dn21p+m8bJnxnQgeTC2rfkWiqOInljwpNxnSdfhLALShgrL+TIBt
D/l7rNZPK861PW85E+XxCFcWbZDtv77ggLGBlwPG2ZAPVnIRuJmJJR8TerMsXNN8L02xcLPEUWZT
7pmQu4u358QwsOHGNpB8Ry9Uif/+lmufk708GqZYj30vGXF42+CKX6fGqrs873csvce6HHZqw+Vi
TanupDg22vy21Yy0eLPRE3q/EpeSdcYLP80k7Mawmq5a9j4onZXxuyYIP+wC6ag6f9tIAOBmkgR4
6kFDSKk0S2fhVkkMXOwtRqp0bBDtmhRQx5Wc9mSBVKVo1lAmzIx4srOHZvoBXpp4MdF7ctDbhz/L
kxKqzLTh3X6AmytpYA521kVtPnBp4yu6Z8rFs3BUsdwuY5rMBPnKWyUvqNxVIp2S62PvoACxJ6bL
NGTT02XSlF6oW1O3zII4csPnMZe8cJZLj+N6ffGhajyArQw9YYjOtCbD2AYX38wyiqLUk8A38pHz
wFga8wrNeqlNKkrVsqwZFpFuQ0gJ4jWsUZ1wqxg2KGTr7p55jvB32K+AgTW25ODTZfuSN1yT8sQ2
/O25WqrxzC0skbRxe9jBdmYs52I2qfk5qA6sQBS1JMX8qsSmHabMGzfLzRTEMcOO9JmaMc3f6DbH
Xa4r+k1qjHo9nIo5wcdR9scjfXvgl3tlTlLrH081nvve3YuBKLc9su3Awt2wJbPucyngUIiT4Y8f
d7tk1DucZHuZE3TcyzIK8kQvRA1fZPRceuMnsFsws0/87qxlAoNdSN90fBgAd3oOeSsLnK+jnuxy
isuQ16Ldj5hKujGsq4mpx9lDgAEinM420lMrHtB1q6ZInD5YUguFoe0NtKFxJzm5KYoI7y/ZSX+U
6NACzrt5dwgs9eFAC6GIP2DUN/16Us/I92um9Btd9zmUgK4kPYtsw7qeBnFziVBu/10mgUAeEQjV
4j9Qm+iO0dJP4x5Cyseswaqi3eyXL+Nuqwo9bvA2pY3coml1dmPjsv4NnoFKJM1CG9cIHVxVJmiR
phpXKrmgWnnWiTLl2dWp6AEd0shoNRgUIinl4hpDqUb4F5ZNp9gFvWn6TOuSSQEtEOPmR8i/7cve
AoA3+FienxwnXhZFAwskbDHJFlVTM+RzRpzDJlLnsuTS3dMYOe21fxPpJGjuOndl7MiPdu7Sx1UX
2wU7SAQ0/rFmw+3iTi+MjTNj1YyjK/sJS3lWRpC1RTL1o1HWR31JgbotzBoO58A0GrxM1Vm96Zaw
JxhR0yaPTLn8DNgady9pjMbaEF80mugD028zHynVSF8foTnh8vpFYkQ/9YmfYxWdRXpbPlZX841o
CtpSXctyeN/73CgmqFHNE+B2Ovo2NSL2hP9LwH0Qzh0z8dywc8MoIzbzd25wSYcQKuZl4QTbH/Pa
b9g/HPdKyqd5giJktq6b7MFfQgoOAB70N26Rvq3xSt2M69Y5yzBh8MKuP4m2KiIhQIPLzd3kUei5
4MsHmKOtnP7BOz0uXAoZe6cahLnq6OhVaNxX2HV+RyKT99kJbFIPzD8QuJQL/lgjloQ/peOgwSh+
eZswlWGp77it30EEqfrUHACU4a1HREJKH+kF0HoHahVN2PhRb8k73/75E+9/ORF/KEUKKYtwrWdR
2mtW/ToccyDXLD113y4+ITKM3GGollYWwyYoLSZX0AYUYGItsvpoLJmWOEkBr9BI0PF+BlMAaq3E
4Qr6cNY25SyNlDgFrvaPXM0LFPM5WDe9Q3foL1LEmdM0bGsIBaGeT8PjnwpryEC1T9RCnGycwysE
RCKuLFe2/BhmNQcSTm3qlTHplntww79arfT3PXkfiuRSAq0VhjMIPaXfQsUN9KqNTOE1HfCzof2o
Cf8uoci5ShbSfiGw3VAYz0I+nvep506JRLiIKw3DopxFwu/waitTWP5hZKpRE3G9PAJPFHlGLn+I
ulE58RhVA2xptAnJcO0A9H+ojewPydOWYV47YzVB8pvHsdehEsUY/Abc/EHMhRcGXNglc4pXQ+JF
s2a0tjrcPZ7rm6ED7G5u/qHKlVPQQ2RlPeACgp8I8dMjwX7YM3KgxmTKGJrj2MqI/IMGim8NNY0w
ayKhlkcC+BaSe6fV3ynxN8a/jyvu9lIcJ9/OdisNOHTMz+GhLQRAvjFNGgRqGQEUXZpxwXR7Ye9L
rFjKheKNif4pRNTsbG2y8aT3v6mmz+X0nsL6zfq5Xt02G3EMzHf/rOJT/Lp+IBof0Ot5Oa2BtTpy
gGn9iaLFbe1rA7Sd0uW3/TKdn6opdaHauyEzh5uq/IjhtEGA+9S2FvW3PdYDcx5/SOpWIDE4efj7
2U3LGmi8B5u2G/l3I+LcUu432XF1Q8+hqfd3oozEz1cX0gVnZiFiTHKEH0al5Glpw0hByPYH66Oq
As6CKkq24mP7CXc6nlFbsNOD9/JF/2zjm72NcemShzDnMVsAG+GvDAIhCHw0Fim3DFglFuA3XQJF
E+GY+6Hs7pPjZJN1R3iIM9H8lKPrXB9YAc+3Yi5w7MKxpYEHzzEiMf8zaPdho1lIodaEVuOFhqyw
6CyanvS9q0L1nLxhSAlsqBLEwnsgOEqKKOt+fsVX3hvLGIW+mY1/O0sAXOfnQIIS0H+9q3Wm8EB2
Udtmx3V/KlKqIJd9EJmu0g1HbXE4gI4s7QQVFKfsFxMxTDobGNluX7ty4UO3+8NUtbN49whCvvJD
70p+VfWE8H9wd0lOYdKQoqUsCPjdX6aeUeqIyzssp8+J7ZKKx1nUACv0L8dr9RkN0pT8jdGweWj5
su3ZuXsSmC27jCQyvfEWvn4T3YlwuMnoMdP3mYdIcX2quVXlDCBWa5niCyzQFSX9WXHa3Z/LJunJ
EsFgLJfp/6ccjS0md4yE27kuNXN886qR7ti2K9XRRY+Qavr6VyQSlUQNXaZWpLsioZEi9oYVQUsA
k8ULNi+5wfOnH7Ao37ZH2I8oXOn98rLZH7eFSXisP5nGtzAEjCoWD/lE0C9EyK7fLj2yVv7oPxqq
5HR5w8K6wiMWj5D01JNJAlvDtagoiCKroD2ZJkHYsUaX/JyOvcbz3WmY+ZAmwZGtUdhvyAx/JA7t
3V9sGET5apEklfNq0iIA1A0RHr/oJvmpILVuDjdrD/HSAp8On6CT3s0gpVuFUUsxVuBNC5eRD1A4
JJZ61iSBrZTqyMHAwLBZO3cbme1LLNpNpGHC4gESoXhfllASl8LP+3Y7yWLr7kSh4yXg5dUjughV
En3S7b2/WSA+Kj7pkzXtOqvJLz1vp/KtWWPYgSPNRZISD41XXr495wvJMLnQLK8OmzcY9IK2eS6b
M6Kl1YJLG08E7W5PCOsivSqCSXm783mzjokhMjzpL2iit8dBRUDSiM+ogJA83Dy2izkgW8k9FlsE
/7Gdwp41J4NU4IxEYbZlG7qggVV9PRWk5JBi6hMrcsjkIllb7kzYnGFglicKT9b7PcMYLRQqrpEB
VoMsL9A/AiHVlfCmXOsQbJFCTbQIue7cXx+SQxyUChkIwyFA8Bajl8qPt1+nhhurEFbU7KxKYKo+
Fvt8iLRa3nk8us2O9IBxtmib6H6ZPIUtSrnEKIh4Dtllxy7bUiqGgnVFl8GRchhkHvON9jzxaJxC
0WHv/9tM2u65z19vAGkZD4nVU0KTML7Permm0huNEO6nzoVu2XKRkrdDS1Y/b3y20LPqjShsUjS1
hvTJ7JT8kgq61r7cXykA82oI896NRDNJsXPneNIjsfIh4ZZrKJvd6ncSH0AYFxMrqUD13ywNXTpx
ukQxhVZDQDDuu/qarO74YvJI2qPLNaICf/Q9WCPPWvj2YYhiQ78/dTxX4xcbaZP/Fq6QT5/Fw/Pz
VmSv23AJRVkWgyeR+DKVnxdu2QUE/f40Yr8TLU/8gBSjBx9oEX+f5lnxSe+MNaND8GWaXDDhVzTo
N6CG4iIgNA74TMSpBL/mijTUcR+Hf6T99JaLb/TJpbKQvW7AwvnB2DAx4gtjlGjklmuAWgnbpqCR
FwvuB164gqCmI14q0PdzSOs/KCMp0QSe2b6cFGvy+XG4KT2ZXoCG/PlnRgkYUrVBWYJuX3ml9Ojb
VmNykaeYA8c4bb0cWVbvX/NVr6QlzLd5gsgjf/SekqGACI950Bt9wp+iBvMITZ1nMoW5Ei4034Hl
kC4IwD5MaTK75L4r8Q42CraR3CgGHG3TxZbOE9iaTkUvk7RAcb05Lm4XYhmRu9ii7eBRIkbdH5+h
/tPyL3ayShTjCYF9XtUlWGJGx81koy5gEzymSC46GbVeDOA/WPk2x4xjnnIMIEcX36s8sqyEu+WN
i4WVZsMRCAyns/EvmCysjFjnl+8avBW2exP81aWY3n3by42EaV10+0dFutJ2gMuY6E9QxSSzwXTk
KvpKqdsHSQ+6ZcuCitLvrUSeRyM19E9+lV8/UsiJrx11yAAYKBYteIjn+GEp3HlKo/FNT7heofzT
xCcjjK3YlIEF0LhaY5EVEaYgpjju+SGSRd3TWeJcnBgYULYXDgWCBB3620P8qWLNDgr8RQelSWQ7
I4cBpx9wTlDdt7NHo6Dpo+oJNkDjvrlx7xDb9D9QVQwnEbBw6Tn6sVINA26hcPlSX3aD3u+fvyoD
XK8JK9ALNTCb1U4tCGp0pZ8ZwO1Lgd0bS7+Ps1wXi38epqrga4o1H8RyhKxLYWzXS7xKfzNOFvR5
ppxDXH4b/Ol5w4eVwkOc2mOJl+/EWkSQguu5ZWShFNY/zwSz/2We/G0MxIDSDwDPIaavAsWQq/C4
RgVQjjZU+IIZlrX4vl/KANFuJW6F4iZow4LLZ9/GQvNJibgzVcAgFiPJxA1XxHRtmZjKZ7reKim+
fdKh5l+r3qnAqRlu/DLNd3gM2fAr5F51MF8gUrKVn32YvyYbhyEae0g+yMPox3NJvmdAqRZwVJeE
zTjG9FMRQGtPLoN5iK4sq94eVP4ZcDUgpX3CS2qE1erdxNEasHUNQBJvru3go1ijhtSfvaz+T9tD
lw4CqZNNW8CHY7ylyZaYE69gzSlqq1BEdGNrwPN23Mx62s4bNHYzFGxYrdK+O7WBVj83SnkbEShT
vhcSa9mduRlD4veZ0N5GEEwmC3etgy1YP7/ceMaELQzyA0nRe2b4ExEnntSj9FT42i8zxmjiXNrs
CrjlGrC2hy2yV+MZtIGlrwEM7aaOir1/nD2420dqDmp8Q+7wXqyxnUw8TKpt/YSEKLXH8QLNJ0Nt
ApoDKHV2uLPaej5/GdbM3N9GeQFJT7AR7VqKJzq/DU+REWmlxmeGBjMGIAxF2KdIr1iTzHrJy3Xx
o/GYeZv7oJLVKI2n096nO0DIrDclNi496UcfE2AnY2N2vlp7PNzAy0Sp4kc0OtAyGRsql5JNZzlx
IwUo0EBab0QLnvMpy2BNZE+P5eoITlrQfWO6I5Cyr0YgHOVXjJWlV7Tb40HjbxbbVSlcE77MuTxv
fwAxCtlv7OV0WUNifNBbJ4SCUzmLTI5zaYFlfwr4czfHf8yPAj+cIpoQ/io/sRTTqjt/PFBkfo3u
sXEqFUoafqO6rxp1EFD+NgjPOix4vqBlI73TyFOPpFTuaFpCBs1GXDPrDtJtHCnryGm41gx1NZUm
EF+dy0lfSVgXXQKrk3oTziCONKul6lJXlabWYNAbNZvCk6KUutXkd4N5e6QnVI6Fi3vs4N1s8bnH
MdNu9ktqlhNsu1/QvpnfmAewT+rMOttSgkfX33s0uBiW0GQo+4sfTWWYaQ37Ewk3JE1854T0q5n0
YWdrMDPwCX5svIXA/ibnrXBD4dX5G0rVdoID0h19KJn/Dlo7Va4ug3cotRL6C0vwH4MT4eZIaIU/
Q/Y8PIGtF7UDaEIbZ22DqG/nlnikPbeUumV3QlniKYVTO9SbYephlJS+mX3HNtg/EWFMg7xnBp01
7FY8UmnE2QZaV/0bz2EewhfwRl+7HDlZd7m+blA0IglQIKNzYcVCgkfFVEdKmyhJpPnSsd+1rE3y
aiRkUwRFPa0UWeoC07TUF7DX0Z/VQuv8SZrW+nWX5d0SNC1cjF1evjuqFFYLgsVvWbyfv9zswOPM
I3NWhrEpU66pwyq82xN9ejTPt5OnmVZB9inz/BHW55l+xVXeFnG8FJ9NyFzxh+xdFyvablAuqlo7
DOmOrFjSi8U++3aa0kldIAcwitpWGyNEv2YiZMapMAOjC0yUGedCd+I7FwykdaqGZJB1qtwWSctI
niURMrkqPvQfhzRSgVg7njMn80aVHizOGTxuYItIpu3MHXJAKFalWhXRcLEv/iv++ttrwOCKsKOW
VGl1BqXv9eQmxWW42ayfo+Qrp43YfJ4wX45Gq7PbOpc1ArZawxDKAelCANPu6NwPzcjiJePUKXcc
5g8QpyJJGftAT0Z61EI3zanNGr0hMgOdJbehOnFWqPi1v7n0fXUA/e9ynsNwqGA4VDcEgIPsHLNP
tsj560gWtHT9MOQLTjnrS9daotXkJ/oUQk/15IvCCE+VD2JNMyAtx29hEg5Dy2egObo+8YXw1N1+
Zwv662Ri3CO82g4rOp1xX6rUg8uaP4NapXXPDgFYZn0GduatnMS/rHzlh4954RXkPZGMppbfIAep
xVE5O1WojJtJ/M+VgmEBP2t2i2Yyd0O2DaDH0JUkowEbZdhnnSRnDu9LG+pyW1WT+X8Iojf/BTmI
mcT8sHk9Y9snNNPIqS/GvRYGRPZeTKqLqCWtJIRtxlesaX5QrHozf7YQk0KK6IHotwetd6zN/J61
cxXwthOgJOTivbfWXXYUJ9VbeZ09ZDs+M1kW0xW6uQiGaoL6zMibB8V7rjPqZm0SPBz/2Nqm3Ayk
a8v9GP3GKWdBvFLs+0UFgKEDSPn0w18+EIjtvT5t893Aya4o48WTsYgyCFaBVRB4Q53GeDi19e27
6FZ3oKAEnKwWly8Pbm1s47bGmHzS2Hj6bYYcRFsOTOVmNbMenJr1gI76/wek7lIX4/gC2N7M9INu
7T0lq/EL7ZFb1Tvy4RBMhlZddqBy0pU+8CpOQs6Dzou3/kXM80FA+uczkz9WRO+z3j70f6VjWE+z
RdD7ukIYho05LzrBJc0ZGDwscgafZuOUXwG4aRWs2zkaDT3BDEClQXLQyzoPIduthFaZ5ixbw+hq
8FwEPULVir4TkhGJgeGILZvFnJEIFEfs3icAjwyiNZCQXjflhD9DIP6YFsANWEYQJzj1+ut8ZNTP
P3Rhp+qcR5ZgLU3YF3EdcK1PbvfLiH+ve8oV+lZnvAj/EdUkdoyJziYLR/20GLZTYwwGJVDnG6tn
xXervJWEv0DtzqSgUGZfzQ1C18qNfGJUHGaI076tF091QWS15P/f0RzZxFW1tHXFi8+4N11iF3RW
QzGQAJnQEcvr9/BMDNsVHhfm2yRRr5xhy+sLs64GUil9CJWGz7RUfCKbwPM1R/AIMuFALXQ3jKMI
Si7ljiw1i/OmnujosCgp8eP8k3pJ+STLrv/O4vnRpSw1hkYzAkZE7b+Kflt9PV8XaS8fibfbESl/
Z13uHBubwTDCOTNe+DkhYEcJa32fTkPYwicxlu9ct9YBMAJ01qA08XxPaF1eKuW4nBVuzupvq26B
9RHfQDOmpYWGmWGba0wPtsbBgw25ipIT7LR04mqTz/7KCgokaEH/R9f/+c4igrqbk7v1Pjv1VufO
5BJS24WgG8elJmcv0F0zDBAYQHdJSsZCw/oHUdmXl77dVH67mNgmAzS8stDzo/1eq4Jw8nWCpwoH
/yPyC0+icWGTH9cTeCNTOnedsWgTCkSaAD1mc8nv2Fbr492tUYiXLTS4Z3vKhHMNICLVZpG2gDsP
Xye1Pwv0nE4b71bcLaPD0CIpXOvkHWS2otIxTIVi0+2uFzfuBRuYqOx/qhtwYfMS7dXCQpYN4t+n
iSHM/OPw/8/pkegIAv1OmSUSq+uXEL+kUYrK7bIg53+cTduLbbBWSP0tqYxP1AujeVz3qoZopKvI
Wplc7AHiXBtc/LtK7fQIZMqhbRr3e89iYw2MHspGjkOHRMPbaV9yICKCbaWWJN2jL39Z+dCsr2db
ak2DF5YbuZGDRZ9jy+QZvapvSSEq4a1GzB9qPIxcj/ts4yfJTI0VX2AXOhpqXFkw8Yy14BLzHPU7
dpVEUDz2UntFn6HzgqqoG/KvxaFBhpKhLZ0FL41gm6NTi9kNACcHoGG9gpNPIsdqzg4JTCbfMx0f
HdAJS8/PjnBmgInsrYyU09wvNYELOB97RthX4JngI+3yJwDAJHKDO/jGarqnNzRGuD/1aiebK8OM
dDz3NIDa2APKs2T98B4PEhbHbNCAIYbF+Pk7i37zgb2ofSlLkB4CgME22rGNvzgIfj//vkniZrCu
5JFKQAtw3eyCjGg+R1uyxB3Zso/9WvwEcwxuIoPkmqBl8AslyB3X6eRuFeKCfId2LLLXWk4YJT+r
hlYhkluwgoxFxz/wfa9bxMp6HVp8I21MHKO/mBF/iXKZGcLgfeu4CoHWSQi7EqQozbgnFMabSV96
gLtuPy4tRqszMv0VOmDVMq3BDFS29pVqwITwEN1b1gCbesKKkxS/NnVifzV4A05PazGQ9IxeqIJb
KDc/1MihprtMA74r//DVZMjG26v9qD0dKKA8qn0Uz+yO4feTL2z0ADLrrypEGxIc66HB+rq5e+Xh
enZ6x6yLOL+GpC5MabAn0IJDAEK5iSyLRNKb6fYS3uIXUJ1uuoQdJX3sguc2Ny1N4q0EM65Certr
F8DlnHE7WqOxwDijhGz3fD9szktireHXlfzBqfGOO0KOapoX74mu3Qm8CezYnyIX5fgTuCOJVlOc
v+QbNdgKLZGISBqNxsuPKcfYHjnRseSSXa1fiqgqSbEvvMbGZRN9Op8NC5Gr2heBWQ8SfLzwR4qC
62J6aDuL/ykfbdtyKFEbxMHgtGoahfIeKZv4T1Rbmlt3XtdXekud0PmSd6ncYKuODArMZoLcj6yd
1Z/JyIuVtNtFom0sGWEMDS70t/t3UVHYJ5S3ufPF0EYV+vkPBca3IEBChvBnluBzrMDDAweilU1z
1V1dOYqVv9LOy/kFGwCum3Z6ccN6ipUHAqp8c0MTyohk7heA+tzhwuUxzQeGZhLArICM8VMIwWI8
Na7h9V8FaSFS7AjzORBgBsDfJBJLI57EWPsikxxWyEREtpQ9PbmaZDPvoCFrlcjSvH0oyo4yU47b
jjIj2M9Qz+7Ef5ea1ikAu3xtQv2iimyBIy0QUJ87cMmmCFkZRAwUp6n1j6F784SK+v3VO5WxZ2xe
YukOXY67PzAP4eczGXrdgoq+yvFmNTureOW/qTQjtn4CwvSobN5SZlUWCzuVYf1lQ3hQuDOBn0VM
D5dgdjx4wRVintKIexSJ3wUsLsvxOUzlNVDgaY/xUDizzcsFYbK3/XGhUIlvW5bkviuvP+5fJSYz
u9KtYPwASWKv+zSBnlYVLgASIsXAgKw4v2UW97n6MnpZXrYVMm1U5EjWNNLP6vr9iSJeH59lm4lZ
knA+K2JO3bOhWfX5oLTGm6XNtTeLpfGZpURk+Ry6pLrQtHYjLsjTdJBqJQiJ0DL85mgh1GcQ0eob
Q9smH4yCOU/EKlOsYAmgbXXEd1vgcUZzOfbio3zGXMv23JJnC4Cp5i/kfXKgm07vzjfgZvsNFoe/
+7no1y/6p2XWJV9CorRcGaBG25NTM8MnOylEQUzIepvb23MIdmkp7sXwcJO2+BeoYLm1QwGXgeMO
UIC5heglOs1GKm0A+kb5cDc/M51XfmP8szGKidGrvX5PUsYEZTs8LSXyb53qjgyl6LE7NJn9ZLtl
mVFQiO4KDNG2/J1/ytlWdky8xwRKklVaDSMMUqiP3fFN0tnJx5v/5f15rcc4oVpJViq8HnD7laQI
2wTv98bNPmgJ7EwDMSC32nj3dL4/pT+0E0sXZkTHR2EIbUaUekB8ISH5QBDXjSui+KUtFGpB7RB3
jUQLdYtsPRXuUKjAq5Ztt5ZLm87/IapSS44ZVf0+P413DxeG7ShruxnkNo2LFTHvcS7bOeAJcufz
oYPcA6y/SP+Uxym01khCgy/iVZxom5ZqgcxvDIDLAioP2IyXUOaHmxtRcwKvMtwY24ODNU6MI9A0
nWVfruRgDJMMJQmCqojZ9COcV8TJi/zxIcdUC+GnRIYsybRI6oVxb0v4nTY02nFvqwlsGFNZgRGe
z0ENtdKmblMLprBSqso8M9+ojMM66sdv+SZtCebu89eFJ3yNDZGIDXZX5Xd+Mfg39YPCaTFDk6zO
l2WAh9GyFHnk1oC7xNhp7BmD57sh7aEV4wKFtdnA4IoVH7dFwzuOA1oJz6h+n58zLVKLOfc9vnsR
uX2yYkFkDt9bh09k6leZ7TMK8+bWQRkpnOpxHa9MOAurkWdi6WWdbJ+OS5NbdBGZUTzhyqLKDU8j
znHMlhoisJgOyoePziczOLAhMaT+Su/ANOnf+hHKfFVr4CeMry+DJeZAasfQSQwzFMFThtVIjwnO
JR61ndSK8deaxuDTv/LCvxX8pT8z1dR0GvMNE25R8qFcBqaH8ZMwYtBAOL9esKl4TeIZnwwgnjFM
OmWuDTA1C1DHJg3WExqzR8I135FZyF6GIrDYRZI5KZW992psnD+Q3brO6VcLfWKyTLSAqzgX9XB/
AODExn9XWw6DumqwFVSEyjt9PqWprB6yeKmTS3Dbr2amZYXqd6K0PA+YJ2SLinPfpSqhU/jKICX3
efaE/a7ScnIMQoD0Z98iJUlnSplbH49I+WFkYZeBOunEb1dziXRkarZtcHQ9L3j1T7lbrq6q5zgz
3vC1gM1yLIzb3p1afD+h+P4Tej72oWCQa1VtU/k14di7EBCeREOBshOVvlUnERpzAHu52xC31IW2
QmVT+oIKIaahvR7FTiTuS5WtNj5CX3XRAJ+MNY+XcHayw2Q2Xhv2GC297w5m5uFOZji9NTBSVWkB
RDih2SX+8rx1IaH8g6xrxcSsyTWQawSEipIYp7H3KwjqlmneGpF1err0I7SIZjAcl++mZPp+Vj1g
bZTmcv0qi502tHTHXiFVi1coRwO6NPbxE3XmsaTy8qpFti4LBgsjw1yjI1G8qRWUnOTaUSEMXdH5
jtA9389X5PjDT0+OKS3zOI9WtghJZg9rCJVLudx71e4Ss6Nzmof9Xp1cup3n9zvr7oJY8XarWGiA
ZVDo8CLCHTqC/AeWJWHM3g9E/8UfC1MvFI975diewLcSgHYpG0ThsgzfKjdkLkqUNCjSElpeqtji
AkonCHd3/se1/K7C1p7yJnQXFT6mRhPbKzBgnuNrT9McecS25TDHMCWxqYlxtaZ7xhTag5Pk4aJ5
TC6IGEDLDx3Ma6amlIDRt818J7n64YzQf7KXZ3C/Gj9EdkFsoD0bHmhwUAEWkSSkmJDPeUtfdu5m
2PEzTjbp9h2bBqZ6mslgsSt9k5c026lEttA+uv5ANqWwnO1/x8e+/nk1Fwt0Jnl2vwWewsAdiWt6
RUpbh4y2DkpHYRyvdYdqRlvuMopx965aVM7VBj0HpkMUhCWtwIKMz9CgOcauPXk48m/veumxIYDg
ZfqyupLt3OilZBhVr3xmcAi7srqTJEROfuE5/ADVpM64j+/eagf34xSjRCh6SrVNC2TngVTABBAm
sY4Qm5yTTwMaHJ5j7FDbutfOhPC+b6p5983UX2Hp4OhooXCY9eViH8RKK5NblS6DN/70E75SSlfv
bcGEqoTSU2+KJDzCrvQtirwVhucj7UXrGuGIxJcaH4ql4d2Gv1JBafrsuGqCv77DKsQk0btM0Hxz
jfQYdI91LTW8O5DSgqxZO5XhmDtMWO/Mnm5oM/0iITo6Fob6IpyQWznh3U+1KShY3Ak2tszMEHP2
mGfXjGV/5xc94eHcKCO6eaPDF28hq2TFnfhGEHi2DWVz9k86rxyb9PWoJXUkBEnWkzL/kukjCMiD
cRXHJ0cCOuYz9YhLX6U6quTyVIB6P9b/Dnt4qljY+PYHA9tQHcMRiPOE6pbfJjWsISbQKPvj4PTY
4OVyILvqmE5jsOVCA85tyw9HYcNFv05ojYZBikYJhyx1NycraTfsRLN2RUgUjARaQMFxd8ynQPdr
90dn9aF/cnhfGQNu0to3lOVEfeVDgNm6/irhQ1e2fEqArizC373fnY/jHPYfHUZ7vbGz9jpj/WQw
bdszVjXGEX3TnyYFnP/56yWZYb5TtvoS23TWZGl2Rd4A1e5xr8NIfAmXJSu11EFu1NIJrbsl8STm
dkVdGJ35d0K4oeMjczPGbDQTxkpi8wzelAILze7u2lY9ZQ9t4XnomjWQKlHyJsnOg1wza2cyE9uv
ccfBxXZrBRq4r8DMGMVb3VZh7IpHH0pnKaq/Ey+jAA0gWXJQJorO2/xiV7y4OR455AQ5aYX5C68Q
QIriqnamr7rDDj4HpsTZOW38iz5WN6UQRmibZ4+t7nG31NngHDG3pePdFi3EvJMRuM0ic4F70UFo
Aj2sFLGNCzkAtEYYVGq+/Il6xEqSYeEbRZe1JmZc3LVJXrnhU0YqCkyG+3ohIVy5o9UwqhrxrDKS
D1ufabH/ssjQbEXknqRf26s7wTbuUrjIon9vCwjBM+OwYy9DnmYJDNHGauYI/NJf8qAjY1UJocPz
rncrJp8Fkp16sjEe91sMFB6Iw0tEnG/kfiMHfaq0naw8KJypfVdUxhVsy5+O3Q/4iX7u6OAtVxgH
tbdf+Q/yOByYvQhqc5bPAmvNIX/FZeBbR5351V5/NAKsnwuQ1pS/PfRDn36mmHLbwtpG9jvDv2cu
f+1yKihLyPrnJ10HP6C5ZZf28vm1xviZFEXej0sJ0DrlGs81lYtwrF3oNMjRf/wTmoLYHMIfWv7B
ytv1HLJVy6U4s8iV+M+2v5XDMUJaPlcp4zcq7m4fUvTVv8Xoy37E0MRNnaHsFoibjxtr1XB2TXlT
aRIXUoA9t9w4AbOI83+rT2N8Hsr8249W3Yu6Xv2tXOKVaRR7H6p7ARxvhPMbcj5fwDwemcTiqR8j
1CGeTm94yrz6hEpddYUEFipF10T5zMsF+ZVILFjyB0bvHiQNInxBvrXcggJ0tvJHknemEd/apJyy
5HL8D4deEbG03JPdEIdD0eLiEwr10C/UVmfST2SFoMvv46pRg2zSEEJIhaqYKRwe9OKXtRNlyT5j
6eBA/oWhvgY7EEg4tEpwi718oYMgdOJUoW8tTH4Lh65HzG4df/acbHvW+8OAp8hhu13ksKxove/w
ShY6eU7NlHCnsos71SlDOKhx9jN788xGKmYSmWXr3DTFyhdFmIn4Tg0wcPmLNDxTkb8HAkI9QXWO
WUxWL1xMjdoqRV8Rmc9cVIvLoV2m0I6FosNlgnSixcN+k++ijKZ748/L2zZgC/UcjxqqlEwOE0mE
/+hg0g64Vae9mNEGyo4WKTf7XYSI/msb/0Yl69BHSbzjg9KBdyft7ZifZ12qyKDPJnViPMIU6jWa
92muQahP071S8DmJSLfh7sOxk+4ltuDlYVOg/6T66J+PGYpj9aS643xNnz8LI09hAahHxznN6KTf
yNHwUC4AVqtIyDyu9LjyWHgXxFkyaOOPA/joDf487SeGKZggMvdbxPVJyNGzvP1XJUpC3K6qKYWy
wLmwNJkdCJ+t4H3/dzDgHVImPjwDQfHUdAC+xpQVtnatBUhXoPR7nnYi5R+3neQr891uMs+x+CX/
nvvuV48jisdW9u4AeZGRmaxcmVroNEEjyNS5FByXp/aIMESVDNbtSn5tTkmB7PkOWGKJn5rsctNK
S2EH9ZdNBTaCkM2HHUXvOJcPYeeqmh7XctW1Fc6M5JlcRvghYqKDj7BZXTWet4Bk3HKHXOck08OZ
ATZH1rvn1jQ6mpsvl4xgdpm9bEDXfWzIF+BSsKlyqQvel1sknclJ7KTI/BEwLrsQYlWsnxwom867
hGmmeugV73r908/RrlTwyj0Q6lQmjt1YeMn273dKLRk5Q3PHEpFDyEgq1zqA8ymGVuAoWpn3hUg7
ZkP1PN6+19y7+YqDN3FBwbTaekwOUb93QhNg67mNxTKqZ1NRQT6iEyZQVenn0v13AJ7LwW9F03In
OTY2hqJjmo/5lSUGM4z7tQf9BSS7445myhSyvlEXSKLIO3ypTspUKbezBhamt9EhF6Mt/8QZK4m+
q2lStXqsUaiZGQlCFpocHGYPlByAwcuZUS5ZQaN4YfT13yWCV6/QwNZTMJoC+HboSaDqTIgLDwqv
JQzBdkF4SaLwZSQ4lDubgg+lSyucjTPnMLCV11CijMha3AAXh8byfuwRmAC+XQtT0kI+/qtuCj0d
1m4HIzscPhLSiexFX+hpmdDXUq9/Hw7hHTVW6zQJ5V+qtCYveBo1WjXnp/QA0O7WLQF6NpHYmD8S
nx+7IOrdX1CNdxPWhNLabtyakgGt3SLvjflTB0qyFMVjs4aviqi7m4SlbYetbPIOiXtGF7Hc5ZGL
QBC7Xzz1vKrKF2HVBIjIIqs+BXQgG9MBT0i+gKDnant76iy4ffxSylObZttgYjUFdQbFoRtnK+rS
rFHYKIhwghYUC98cKobzK4lL6iTaYLoz8wK7DL940GmgZaGNyp6zvWG2B0ZxItIAE9twLvKddN0v
T6CE8L8gx4wsgfsXKIDZTb/9K1Avg75xx/mKFEYtizoXADvlnDVcBdNPTZtjzYkO6ltG5WMDukX0
ixgKV0uqSNRoMhAddg11VTowpjA3Gx4LU1vMKZyCaPmK63VQdp1J2MgYS8i14WaiVM5rOm/msddA
pHAMoc6s9p/hQlFA2FAode5Mm2/O8dVWHg92S4cLPOxpg1USjzooWC8qNYmCf5gygnfWh72sxPgP
JWfKnYh31lLuBDuMsl+1g1fJNPEsNvkV43UndoYxowPZo1WNnjRa1HzXXJ8kzFf8JH3G8kIXfoks
VadUGRjUbn7/C37SLjA83wci4VOi5pTTdeM2SWmUjiKTsh5z/+b3uPBRZS/x0OC2uGE7RAOjUY7F
Y6TNEC+96ieXMU0g21PY5FtW5kka3xIp3dWmn6gumcDzBZTnbyrt2SJVvnz6JHPyvciqBVLygIhz
PlqED16D8aKOiw4IN36Wm9hgiavYuCPG80lfoGpPKM/e4XYDRahjxwDGlRsAaxJrO956z04TrjgS
nCNaKlyA/maKmH4PaxYJ0rKR5t7Eiru9s2IXviqmlPtbE1gsfOQt1TCCh40Ao7GWoGDR37e35ndV
D6MH7sUwgGxURXKY9eei436UX2VmeLH6Rlo7L3Z3W9G8FH+frVMv+b8BPoiuXSiuC+4f/PePUk6x
BDDqTEZB1V1oKjo0SEM8MaVjyA6YY7AUaAhZLoyX0SxlGobK3Q3Q1CHqixStjL146PodBQWCNfvz
cZXV6gPceX7M79tT0kDKWT4LBeueo8TtynKcrtwvqaLPjy7fIoL9vArB++Yazl2hnZxVsGjLrKWD
7wwz7VxOclfcMwhE0/GnuYpwezC7CE2+puphpv2kmJ6YkhFBPjSdF5rCHdEmI5S+w9EY4ME3sAnh
RzSDZwhYiVXj/SbO3axzySE7IEZEVfgLFuvl9/8uU07zU95ukylQ4w3P7ndqMUYZz4Grwq6Me0YA
9GI3JjmzNkK4xcgwAejapV8wCfRcXlVdZxrUcnD3w07w6oOZnsHZ1yPjRtuiPB/cg9EPaBXPYuAJ
CcXO7oIKWoVRSGA5S8MLiMBXkdTl3YZqLyyRj7CzATmjTWGKj+1GRrVCDQ75r9npnSXP5MkBjZZT
ueIfRJULec/VLzlgjbMmT9AJfEBWs1Ayi8yiDEB59Zeqr0DN9DlEbopjClW1ddnBHiVz1yAxsMFJ
9bE5G2P6N3whHGuiXoVjdL8YyQHx39qtlTzaD2wdvZ/w5jVPYj/cZRuBw5xNmO3IuwPDYnCGjE3t
TCKx4XGBvfNf8UsTlWQVFlSRp/55M/2J2Vqu2I1zptonsFNSbI8GFNl4erq6tB6rCwUsR2wyXF1N
Go/Yd+GvcA29xjj2XGFbOs6PWUjJlqDR0kaVu5C+TGSsE2VGVx859+i+5x7/KUAAdXxAhMET6mcE
N6383ssW8LBjYtdMp36w9plZktFw62Y3kQqMuwTX4DMuWlH54FzQPfEOODpmY7Ua3M3a1tEOXU4X
IghWKvxCvsPSY9mD2+CwtbvkIJUTc9M/Q3Pqqw4dZ/e/nuRgnuTZ56uyIp2WNNWuAfr3R8CPaM96
nNW2bADkJnBkblm0fPuDfEND34zifBKbUqzMvKjsJXvWk1nUGllgLlzH+dmqIeLTyLtxvq4JIeb3
FcFVCruwqeFfosFZYi0NUv248BpO6emGdE/QuD3rijviG+OfJMRTtXUA6FOYuele9LSE/5XlFGo6
bJGplGVtkhqjetvXRHiMhG5J7hDqclDIFE+U3LFPogVdczSVcONBlaLw7eKJjmRq77Ayod429OlI
8G4bmyiDR+PVhFsEfI/B4y+6SNOqB8XQEWLa0ijSFSXVpzFJL7Mr576w/HYh2j0+ZoPENbRFXA+j
GMGkIaeqwF4BgyRbrvOfg87S9ojNtpRcjTu1BinmrAHnWEDQpxEhCbWKVPudSSuL/D6F12Cw4hIc
H0rZ2Ae/tGmq1S+GGOgBtkWQr1/JXS7DVO5zbis4IhKXNh/h3It7WBr/iIghN6L9+5gX5hzzyf4I
QUClsrXz3ILaciXcXHof40VqgxAgedHmB7/1NjwzT/2+bJHYkgdK/IeHzua1irY+gkPAzCYrvNL8
gDqGn3IV/o2R2xWdGmbRIt9Mu4WBpW65ACF4GZvGOYzroTxVAiib9JkRIyYDjGlkq7BEUTbRQhlG
j2nAbbb502n50jyXaLcD2StJBIEaOkWZje/z1uxHhwz0vP2upeSM8fWOmWMvChuNcs+dTHbnJpgJ
PcMtD7FxquaRCpqbzLkG+6cnXMko2PRyTwzT2PELsZ901/Fbiq7E5PrwHEfPMud8stHROomXRxrZ
W0BvD7frh6W+Yk6usSBFLhEJ4BuXBYATjRPAYTsWdgPN2zgc2HwIxuVPcNTIa21AMQ45pXybEBpg
VW6wmqRZoasdTF8LDnO3VkpGY9PUs5JWn859G0OomFp+MUMZwP5n0oIjPSf4QjWfWL3Q0yNCbDvp
+E0X1mZY4YQSSp6+QKOMDnlLG2zg4tXsGfMU5OwogFhLGaTuacsk9Co6XA/D6Zb1mvn08s/HTDdn
VMYOm29eqded6+dNHHAyWMWLdvmKjESYrER0fNZbwM5RleUOV/kJVzlVRuLXSRoW9P+1W/6Lg3Eq
OZF6ks4brbKAxBUM8D6Jc3ATg6/yCPEZvH9h7yTsTJ0XsI085IDHePK5e3ubFFXHDRjdOXo0rTNQ
7PC2v47PISuPRhdc9xrfEdMEILv0H5HTUMsveM8/giSimNECTqkEUnUGlBAbeKqQEacKj7EXE8ZJ
BrEE8Xv6TY4pX6Gid3H1qnWkaAirdTWAuM5BaVqvx6I1KZW6VhsLnsw6p5gvMqSfk1dPS5g+h2KW
jE9CZ3ET+W8m8Rp1Uv0cH8pIsdOoUutSeLhcP/XtmpNxxYIpj0TqYr5dMmRVqhkZLOS8IAV04c1Z
Ltigy7CjWeSZehK5cYaAcnt3XvfgEoU3sPeWUeu/ZhWxnma0gQcsjTGZ85102F/NFQXRzj1+5Rsk
8qQ8E4dIp4umPSe3niVZnKW28aeq5CFwfrA+aIShYlfbx2rBD7pgzzWLXyoq9PCLJjUsdk1N7GX8
zPDuT7zuvhqvIhVRqNoGArM+kKAQV+alhMvyQEdfagRGsmzQ0R/9fFus8TGTsVAIJgH+eCLaO9nx
A3snGdWSyOl+Lx/4xGEV6E5l9kSETWNFOwsMA6Z47HMfYgwuxFBQaz6zaB70JLOdHEyTMMQ26kCE
FQzGm5GEdZDkOXnyvnHoDrWNEP4w0VXEMhAJ8IP3kfTWbBafuzY7U9KbE96cyUcBcCDQ/0Y566WW
AGKYaUb2pwCQ05qkIrTnnie4h00bvRZ7faloT3FvJ7AfLOQ7XR+j7Dmvqp/Sg0uL3k9b66hnc7Y7
2Jm42+Ge5JeJ622cCy6Tnouh66RLaiIc8ZbtRKzAIEJxqUsIIGk1BbaWCQ+fJFcjriX7uN6QOSnd
oYexct/nNP/gJjkbLYtnulsi+Z7z0JGncIzWp5/oUHVkjWBA+bh5t7ccfuftkU2iQgDts8/04vit
82PAAcozL1q81RX7rfzXS3Ux0ymMFWVqnN0JKbrWMgmap18W3udIY4NPMtoivP7ta7MDwOgcuQ3x
bjZ/mNLczpll0GUWpdPZ4Kk9dbM0XqXD7uixdABcFPTFv12hbQ+gvq8ZbfqCYGfbwbiuKRrRK1oH
F/+Y/UlNbxMw04Ki1FAWccXbcddbmcCc1Npl/jgtnIeo0CqW6OtgQvEatGtJ9Xj3BKsFjNwNi59C
4V34ClLDFx690NvkQgMV3rveO1cA7GH0cHubMoYxCrR2VyUa+lADBvKtpY0bYWrR4is0ZnCtOzZa
R+oGDPrHWGpNGTcuDYR8BiDKg1KkuNIrRaJ8knAER/HveGbn+hUUisn0jaKKT4UHCRyOi/40iWiq
CheDkMiELrEWGAZ9aig0EtBmhGnEYzS04ijEVBqJmzpLGfVjLaBBSRxRhqxFNaZrjgV7BGtvCLb4
iyGqbg3oKPzLB9ueDexnmwR56fT7jBt8xUi9PShWwf7WfE2OPVs/N+5lKrGAGbJZFbG8tl3Msybd
t2qD3KIgXCYq68SMGn6HTjUEbe2VT5jR1YItA+A8kzlxSNdFSDhSfsSG5YincMF8+pT144C+CU6R
c11JljXFhbsTGb1RER1qr60g6RJfJhHnxfNgKJpsMXLNbGnX933LVALwPrTsfCDmgFebB8V/P73Q
GMvnYpWgFRrAoQstBlOiAvnZ50tC/ZZUP6VbpTg4GNRJ+/OKsWwKfFZXhlO1ZoMXZ2wfLPNIfaB2
6rM1LxEFIC1Oz1oWqtbi8EHuGt7LljR5NTutyifIkITVmVTiW5kmZnWBWxFrQxgu7doWbydpjcSA
TDBg79yCKv/X1BtqTNG+dBjVjU0uBrOncPAHTufN2fGtT80t3mCpZ5GzsnmFlx/8KKhaaKN+p5en
sUXiBtLym3Orv985WSDXAHaMI/nGeuGbePmQUKd8rs21AU9Mp9iq36n+0ul7IV3/mEjpEUKGDooW
hz+jzH1h/PvnPGH3PaHfV4OKRsOr3h/VqNXq3yI78VyRrGOtAJ8zgNFUGYEoSm+QjgnQHutliKdm
G5+YBo7krgqGugDf300WVvOTfvS6N8son7/jELv1UJfHHTmGxqTVS+p9BmaMGz00/daJew/ataCz
8EDlfo+Ud2EDsKGwN+A8KUQnNKrvNowEfpmqIpBOx3eN8XC/sgzwsCkrzZMAyV5CrD9KlUhrTORE
g4vUTkAVBkqi54Hz8D81QVl55AYAWaIlfCXzG+xyRZise8OH26kV3FbeFfzsTSek+WJ9+zCvR3d0
8qK+wzvQSDfg3I35P/LsWoSQ3dduChLDB9XP+4zhi0bNmsDIiG5wq/je4aTLB5kvYFOj07bfcINK
5X7njA6yU0z6cjqu4tKsL0zp0zF7pbUgUPJgRHZqYr4VKwe8Vk+ixOPdMRKLJpuEiwRwbjzKzyjK
r34p0AqeYqJs/o9mL5pTgxflHbKb0NAc9tbBuUMENIhYaHHijN+oCdRSV6pKVnhK12UpA0BwRipI
R+Ufz9n0YfNLU7ukIW8tEvD5jyo4xR7ZnsRjXbk9reSQsighZrRUtD6REf7n8lfvfuhyP6N1Qc6x
RblNLMmJFnMUvltNInDH5zEVJHwl+7wBGRjQ6mYE88q/T5d+5O4LtwHL/eZkOruE0zksHdXdDFHm
n0resqgU79Oy/VDoZMdln0KP+XvAbAxf+COODdgXBcotwc2eOHi6efoBKC3//KHmAYWAvg8G5/J/
/uJ48xfWNk16ufCGzt15V8YaE6Dx6h3MGN5AKBaoWwnll3K3DE+TVDwbNb+qBg5wQ1R3s++l16A5
zjEhAF8pTfEWqR31EeYCA7mr53xFHe2bP3855wwJCM1116xqbT01RqKma3I4rMwSUtd77QHuNIq3
d8Kkb6IBi92O6fgIPXHOtc1xMwoESHGy5LxA3cpiqkTUwrkcT4BBZDP2ppTXEFUBpxB+YGYuHhf/
4+JXM/YNdPlh5tPiIbCEZXK+wRKyu6pelrFP4l0BrjnRXJhEyGT90sfXRA4lrQluThuXacuSimhP
+qc3Z/3mPUIpO4dpBssmsg6FsERBmzBps4mnffCpQrwTi6nqPBiNqsvRwuks0Kguz+tCaV38WUaF
fj2ybsretBSjKGVEb1wiWoVt+8+7Ugj1ECyPnuO7s028FkK2gEtVewmJ8TiS3PirnKXzp4kSKWj4
0Av5y9D2IfSMD160PQbgKW6zuQ6Ov/uEG2P6mTMyR11EuXxWs2YijIAsLuGBx/jUEtn3kvIPFQtT
gVm1wsXAdEcM3AC9jZOAlgBGU8/CNgC1G/TayrzRyhOrbwjj9yYYTTKkxekvMFdKoe+EUwZfeegd
s0ftg8+1JXH2D7XI/EJZCVExs6otjSE6iYUn5Qs8wFthRi5V9nActVznuVtHCHsuQvWitKCQx4SN
xLnsV4XN8MYpdfrIc4zH+vdLzKb2l/jgJIvT7O1PVRP2+1ecojVznb88LY/rAuRmd65sdMonnrYZ
664p4T1H/WU2gnzbd4WgcRrlcpTetYnCtIgjJbA46wVv8UgS+K2GgyQ4znPHuiy3/aAjs0qBSSac
SfLYFb6WgvRBuOv89vZbewoQ8FxXNgEtentbMZooAX2UPzmlDasK4yE0Z0hfEqK2TJQm1c71hevU
aMDB1TRdSgZshy26JPyqqZNWgUtdIVEUSdRqsnfzKv4vtpQUu4JU8Z4+DoDbc7A3XRZWYmRGZnKD
Ywdn7EDlV6MZO5mLMHD5U4PyEpm2vBZ1tue9pTCoLDrEhNP/fTQEOJMoVal5gbeNQhv4D+gPLpSY
1W2FpeDkCNH6rv22gLoQIq8pNMRfDeQ3lez1XntiYWySi3kxaMeeWewbrE1aPoVk3KbbOJPrOyry
8k3woNem+KXDs97a0Q6FECjn43MbKKeEQkf9pr5kBM9CGgVNdtnBHcELFGQHz1Hfu4X26eLusQDE
alE/oa6OpD670Xg2scby7oSRaS1sxKvQqHGxuTqjEtWGkAHEt9vdN8bgAegN9FkEiUvQD9NBCpgX
EzvcMx7H2UZPd4g9eAsYAFeS7bp/fmWjId58k15q3g6v3rikoXldSXKNXu0CM5owGesBHoMNyXlR
pgWhCYC5aB00VquBS+0xHZ8mTlzXlxI0cVpJKjlCflfqEzRABUc3P8PlKDdnpffiDKS4p4ipr3ET
Ypdi+fHPHvCw5cOYvZIn4veoVL9yHjtrORge2G5Qa+oqEc8lcjEHEwcgExaArEgrUylge7zNm++8
A+WO6ramGpi2UqObrOS2dtLDKntekcpoD0BLzSIC74vU1sjz7KEEBEmEjuOEVAzwY/ljzGAyitfP
Y2hLGUZ/BzwpZmXtwykF/VCs4I0L5Tm5Tv+lEi5QX3O/bJkTUd/Ul5wzm2FvHY00FOwA2TPUttll
uLkGE4nL12/6bf7Hh0j7bFwszp2vTIXFzFGRj6d//3UoqORrA3wl2MzxL/EZEK+2kU6dCbOvvnql
VIKOeJR4iMLk0kU4qvdy6RIX1ySVwxPGEdxYhhtlsdixQrQj0c8rUXiNCaUCp5eUf/8T3mbd84zR
vb2FYBlFWPY3650Nla7+eImoJyLkESGsAz3p5RRqR+vWTBfjmuWrHAa15uIPb6+gaBAu/s6VDytD
Vk00RVYupm/m1I+12fKJJhfbHEd/m/Za0og6GBMNtVgTGk90BG/BIysHyRdNzw8KyBa75pHSkMXx
MbWKq9cQ5l5CzpC7+7GatlKLH10yGMKvUNjo10eQCb/MLNSkBY29sHrg17WWnA8hSCtE0Cxuq4tr
Jpi3KStxE1YTc/4btiSWDk4iFP2welgP1Of8fM995oZAmFsTeukscLpSo0x0eTVdKNCL1NDzjqkf
ieepPie0BsBkNbWd/vwiAlzWsAW3Ok4Vpx/Nz+8GJJmK9QbWmkEnw6cxvPadEZFpNUBhAPDG4fk7
Bb+8RQ+NwuYFB409aa6vYaBn65Q2sBSUntkarzBRMg1KYXE9WW+VEW898Vj9zJZEdrbEXNsgJDae
pMTJG18r9ZvZebU+ne/lL+l8cSNoZA4kRu+PS911oPd1MZI6FN+eZtvpeZlt78Kd7SRoID9WRqLZ
uwNW4mjZSGePsrFa2m2FnjDKhcpmY488ysGq+/kCefkuOSchDu9OXfdwEkf2oDb2MRcCw4HU1WGg
3BaBcdw0MoQ4gdm3I7qpL/4t8TWRan6bBXcMaLS1RIdTXdwhOZZgt2s7E/R+Y32EBfEphUyn2nPB
KmRfZvVMGLTyS8xxbFjs3MwaTVj8U94TM4S/8n58oa3DbnAq/gXxVzMaC/uq2yC/UrSm26ukOPRY
vGiMmDNPycnEauiVB76Tu8PNiwOEy0TkLTIbiiGTkqHDdJ79fIcNz0hPj/MYyVcEUKB5GHoGTU63
YkdRXbyqJaRHzxRH6V90APJ6wWIH9Xytt5+mo5Ul+TAMvVpaVkByX8uOE3m28grLzeaJFD5PYZs0
AleyifF66DNooE602OK1Uh3nGOrjvTWBxSzqQsrf4+f6VGthDJlsFLV6SV7noIuUUDU0M7ICzUsv
EwNQ9909xY+TFgg+BmycKOckSpJAVv9l9NtlJgMdtankLwanMfyFcgP+32uNM8XQaj/aaW2MX4wK
zGs8Kohv04Q3tsTLXEIltSM0t5I4lb6qMI3trorjSWjRzg/zRJim2bbPOqRrXF4jM0w77CaOAF3u
7Rrq7tztXow22ATuftnUG37XrQF63hAiIJfw57TaI+4YU+j8z6bLNP3wBUcCtRb9JQ/cQKVt8Z5+
SvIzOhHZmV6DrP1xNRhI/ks5HLbviXVWQrxCGwkeHnd3/4dUfsSyWdcdmMH3OyPIiXvf9dDMoO1U
pchqh6jJRe8HEiJfe4n2UCEpPvgPnmqyH8Gv4YKYF9/zZWOkTVSL5jSuI0MvXPZSvNBX3YQ0cVcY
BsY/o/TmDNtpDZdUKNsvUNtcTa4W00Qih7VnU2WKHh/TfPgZXoPUYDU/Gk9qhvvPYGYkEdXymrPf
WkNnsKA2Gg1+xNhtaId5ndsOy5FYZxtRENBMsFsxOrA9IGoNQh2pOwFTGtmENy31DdABhqd8vrw+
1rdw/PypwRVLSMEFLcyFONPrOCQx32bUMLgxgLdsGS9tnR09ZhszNxzDOkaQxAYa/CL+DiwKLXcO
BJ9XLjniOBoz98V9omPgS09mxQoAocZf31mwukEINnFX9WSB3zYLR0kDGIowcysi4ICy/qT5mmxf
eqTu15Ekjk19cLoiKWPMmMnF/GqTHHTRskKb0NlRPlwHy1rJTVp6AiDEm5g7iPEy3wrPAikBxInp
3oxjeX7drC24oP0IC03+oTxTrHw2lpny0qrfPIRq4yKP13uo/b4kVw45+do9azHYTlzIRSrWXLTF
hxfL3o6rR3Iy2wGHt5clUsCsW9+hKM48uNIlf+u46cJyzcNO2izjZSLV0ca8iIfuuNPfJutvhG/M
gky+IIZWiGGdlHcAc217tDUmgeQ41ChwMXYcrVG6UpCSeeqZj1l/EGiP6F27/Z4RLQJjoyAl9HTV
dlQzXm+lEHPJDPyo6ZTpHy50RxN+CXGSHoQtq4Q6Nuh1q9c6FGgHDpNsKb+vFpNhPXRgrscWGCbl
xf8VdJBw2WnAH86aeefSpH+/7zwV1ShBqZ/tOS8k8L0+ZE4JtPrXEIsBRgSxoyCloeHW+/72j5Rs
N4IFpVlymKM/2jf+YwckWA3WPpE5r37c9bXEG2c9t50zbMqd3eH/5tAVX+YkpMOxbWaXWXBcPLlR
AHIl4ujg14qeKt4jDO+tfWQY2CCnIxyZ8mEFnPrkBSGfKFoO4JEvfTTAdaB7cWZJ+UbUHUqJr0Vy
DQBPcf9sVqEGwMBHZPFCsHD2LMBc/ST1DiCR9jkb7rEBWKzNCpiaz24bvc6e7ff8bhoRyRUlMvQN
e4SFZCum+y+u7LuxO6iNe0OlZlLeffywi3suFkxIhKGWQnvcKWKgBqu6BeMrvckDnrhuIrc37d30
hdht0PTszcC1It1HS2Vw8N471JxLwWqnOghTJXDa/z8k/7uxLLNyZ6qWypB8BMnrgH30MPA0McG/
W5E87RvZ+4+wylHlxKIs84KZc6M5TlAH0DQaUO3QiqRzg7E4qDFWceXt1itpqOgiwl9YmkWYGSW/
74PHsQjghjgTtPw0kGTypaj/Gz1yAUmUTVJIL6/4YGWenVXleZS7AaUkZt5/v7V37v+DU6VmNmZ3
mnCEqt/A6BgMu1joRItKtLuB0r9ytWKURM2ldekVDIFPBwHYkIFqQoTtdYu4AwfWDDnAiidhFcs3
Y1sWwCgiAdd0lTPQkaZWwPcalfJWFA8RzmK5eJOT2V2SGNqEzapE+xWZj3qR6c5CZubW3XfzMNIR
cKVz6pwsfqyz4z6jXs/2n9bjCLXBlxCstIfVfga6fA2nN8UDa51vrOISXtoQQL4dvybpCdPOzD3t
m1kTYpqhP5uYmfysjPmoCcikcwaJyrVi7oW5sQ04qDRuIBjlo24Nq21r+0wQDluSlWTu7V6y3Al0
mVbgkH3zzXWFQPtylzBB4q0Wq1QDkcJJq8yarx7wuoSwCXoVIjpCoRu/mI7bCfDBU8dD3qIsdwZf
FhMPUYhBcm68NseszDMj3po+A2VHeNhQBQDAXWZtDzUbANnERCjp+6X8y6ZzBh8r3xnU17dvzLr3
VrEVUeps8gvyGPGl2EDBZktW7D1aEooTPCZiGdcwRD7bjN3RhMiCTLgwUoNBT2gYNdxwYy7TUxu5
JkJq5yTkl+YzMtRtMBu507L/gkoWkLKxkeccJfL0PLgZPOGcPIe3skumHWbjZzLh70mNaShMUvuL
JWTBoZUG+grlWfDlmcxY2w+jswlHhdCgru60HI8ajDGpCG0XADhrtmpbinRCNYpP+A6n9i9JJISH
f7lf8W9yA3LFBV86yVyOFKjr+qJfUwN3I7hxPsw/jcSn/T9140CRd90LMwI1LBHpyOlMJlxeO2ZV
PRGrsIT/oq4Knf67FqmdO10tIh+nYM16y0h9/o5ybSmCqoDVQCphOXz1ZIp1tMXQVinJ7vokY08e
Hwpb7Y2n9+NsuuR3oQ8TXYjpiWSK7pIPtq5eATabFN22p7kajc2ketsIfQ7Agf5oNgUa2sRIyFJ7
baPMg14VS8NKn22Vpld3jNA0dI6vfeDsB8cwkRvgbE0jzP0LkWXYa2qxUesqSv35pzykYkweUkKX
G/Q/jzOyxHRHVfjtjSNQ6GqUTvhkAhglzJ/Yrhloyx2fzd2aC3+qamJwIjDjZ25zU3Mnm97Rylu9
m0Wq/hh1eliozIq9IG1x4GcZuLPmDm+ab3N1jFqcwX9H1cRxcYXDg+4KbNwm+MlpMMmrPOuqXLyi
so+tXGLzTU29cOl+bb769ZANZ2dhyX0W6276qsw42FwdeJjLA468aRFBPGhB8NqoxHwbH+wHfYrR
k8WtsREg0SIEg2hu8mkizTaxGO7A3fZO82bRas87ef4/TqA+iB40fjN+4kj5J+D9V9Y7gTZm3Rw7
X34r8dcwfJL7/0jbFQW6fdAk5fOLDrnxNJfk5PtCboFN7q6tE1zORRm2XztELznuB/Pr+j9LDSUJ
CcFOzeqSI+Ke+6RqXYTNJjl2YXkIsOEczmkDj39PCQzRny8D41h5digKwNbqKDcLltfw1G9NWR+p
3Bfi0CLGO5OqXMV4WjKKCT5NKcFq0T/4iJ6J7g6dPZBiorsZuXf1ziJjiSytgXb+T8C3fy2+16dt
B7evlfUB6Emv05wYggI/3f7FmL/Kr9kcV0Msmz+rI5MA90d39eKlSCSq1T8I7lgrWT5akIuUi+hJ
glcGtNXdU/TRdH7x63L9mjoy8ecvGBgibTir8JvGBlx+60Yd6aqsPDxO9qiaKSxTreazEin0RFpF
feiR8NJa+g+PIOZjhrlQbp8/uvty4Thc5R1EqcBv1rJ3OorYf9jIJV6OKmRVpRuFWVuOM6zKfMxk
VsuTuamVS+WEWW6rWnofc4GHjzRbG0v0ChK5kakzfTMmfs8FS9RlSK1smj0HS8JrsVKCJbtESeyt
+LjCEuJm1JRVwV9u3Uadjp1Rb0oD7zvW1ca7UcSUkQbjl6+0mnnd9rf10abj8yZL4vZsWz64NhaC
990uoJ1zzDaF0nKV926NgMRrZbNvJZZlxOcpNKhyV1sul/F8+smw7sM/AYWW0ds9Rdd5UpsXmzba
zF/HbUw9PCHDwuAa2pCx8+e5n9n0xyORwShtRvq68sFOQe/YRdWSM59gIwc+x+tsprT/dfPkuDua
0qOcYFn+C8Y7kkomUFbUBiESjFepK61/yMtApOFufxL9PzcdThdNp2/8U+DOV3VLXahPAqfY1RuD
szNOVAjtlZHrkifs+5vYNHeRrbhxjN88oOFruhdliGUzv5XdASmqRkA3EDYo614/7b4kvVadRJRI
XX2hhS0tJwhr2OB4VZI02HiSeewZ6b9eTQtMVtUDD25uJ1HPO/DNWBSPG4/Dh9BbKpVt0ngH7ChZ
LGyIMjJ7t0ACsVEOQm5e5Pk8dTaHQAusUBydIEvz7IZqTyvMijDBNFbxr51S5n6hlxSHre9FYBqW
ydX7PHSBD0sTJkb8Zuz5mqDTim+VAgAynyi9OA4t7FsaPf6D4x4Hl2GlKuyjhD1cW8cZ+lYyj4l/
Jdu10h6b0DjOWueesEqiF6n3PvODlLvgH8LEXNwgJxwHhi7Zk+oNSBVOO2AuD/5kGMVqldP9hzmH
TrXEjdNB3CqqOtgyWNjywtW/Kixw8oK3H1mPqrkRhrf0rh1ii1OS2JvtWZ95ygPjA5SQyyGwixld
72Y6K5JwK0N8ceOBDBDx8p0HoZVY8BwG1TylzA2tYOLVmFoCZgZND/WugMosq1zTIkqoz3MBRV6u
X0nrNApnKYtzZCTtjKytpKJIj0U30obcHJpxFs72CZb6Jo6neHfzh6iUuLli6cRyXTRlQsZtTXUY
7LbNYnCJ3C3m4VGoW6DJ8AhrWKbusJHuzSzbcEAbuQb62n+aO4RYqSwquCzOf0qU+YhopgbVZdwc
7blf/8fEjFmstMl4XV50G2sHJlBGw+OZcCgIMqm1PiEchbkSgnvnJlBcrUsty2tpzcNsiND49hqI
lMAob8+lIkRUnp8uMpE/Mitn3APqZ389sNJMmbPijRvlUzaIy4ncfd35lfYbKUD68V3/MFTAPeY+
yRRHj362iFJz4TvFzGsOAtMBBBigMSXUgU0bnl8eYk6jyO6dqAPxL4oKMIaBrvpmW9KWEsvIw0IB
S3R9NBLHJ/+OsucBPTrHEz8r6/I8KTs/+IL1HsR1GR71E4tk0Zf5WBJeXol91xsr5BUMJ4xs+Nx0
GSVSkYdqxpEWs4n5pNr8pQR4wH9KIlFiLugaIj7g0ydzTsC/MI1wBtTFxJgqKkSRMlcI3CFCh/6r
LxozCzGE15o5r8QMSrRQ5b9uDQjHkHWZX6+r/YStLzrs/aPp4DTn2UCAoWi5h3BFo1StVqzOZO24
Z1iEsC5B1iMRSUlMsZtgPOPoXedTrPizjbYoF15mXPFdQuoKLHtv8QkuNOrlFSpsXdJTxyTKkOcC
8cpXCXkTHEcV8E8TCBpnFfDNU+GWcCCOgDM1Wyu/n4C6s38K9tsuKEly7szYXhQOtfgWedFpn9Jt
lIEm1q6whQNkK+/DnuR/k2wB8ck9xtbnZ2lES6xDGeyPRPIPVFcy3CpfzvMnabImteWFKP+EfOQB
vEGIkBvirS1nupRDiD0SW5YV4/21sydvJnP8bB1rDFHqSzds3KtRClZUabnbB3c5ejZ2NXnvomZX
Xd5BPUb1jvNgbbRwF0TEhhpVgQYUKnXgL4Jva4yulfDUBXkVz8Sw+l3K3frbDEsVTP0kbrVEuSc7
cDt7huqaOeiKEgCuRRi3s56CKd7In++whAUTZQQzhRjHTsQEd4bG5kz0TQ5mx7goMTiDmNgumCJg
irDsZTaNfEaT9JRVEUYZFPeSiy5DOxCeTqr5ZN9uNk/2RzNP+L9dYvJ7Qwfe4vOWNt3nWkRVNM6w
NBWW7eUNE/J2hSQYIv8lh8YiKd9ixjCCv3VSROnmm5ZEcUCfA4NdiaAQe3swOzhSYggAfjjHACxp
XM4yPwlW2k5pVHZdhg0U4LswHKAPCiYdKcUMGYuVA6UY1pdBSOXci3S7YthLYmXlplwBMaWET1lP
B0aDg5Xmc2caAd83SHS7ZsvadOSWwo+IHvDJ8khFV5zKHBfnJtyI16tLHddUom90PD9Sx0ifJgT9
TQkxvNvbsnlrLbZuhYKKHeQTn86zM9Tsk+P63zPLO6lbdnkKgj9XuEBVqulTfJiYhdHbWuHeZvgG
+wVDa4RAa3Uj/rPtUfhnCCDRa8F2Yb4z9Udb/khL9n1GcLPRtUsz047LbMzCEfytbNazLwmsPLfR
yP7YeIkSU0XrW1dX+Xv5KSzZ1KMtVw4cd8yWuaE02Uh+E+cU3Gii9sSVDHaFd960TWNKjzcl7gL2
1zLQu0drX2rx55xUCbihWV/8RPPHay2PQOYqTsafwN25qCn81tnx6PriHikQDr4uaLfuieMjMkV7
B5wuxoi/KsbCTbahIEUFxFTW74LQ7zQaWTUzKuys0PrNOXfVAyZ9qlKOrrKGVJS8JHYxoVCHGJ8C
dCB8jaGi1/8st9WYvRB6ltoGGtOsE+5TMMcrFUMf9oGefg5m/tF/6unqPjiZsp4KM76cGyFZzNG9
F0uZYNuvwCxRutLzf+BW90ORynZ4qPSX+FJTgvh3dLETEbAyrfCYudpJZJ4A9r45rK1PpfHmYlWD
ZT1xm7pPRLuk9a0lM8pE9amAcYgdD5nX7IS0SzpuEd3f7fJJfFSlWGKalicmhJsZsigwaTeTFdYB
upnRa/3xz4FCvYbNp0RualEVhzmbozi4lu1iQ7x/EX45lt/D+PLVAIHBFwKrJ7IvKlVFfmLAv5i5
t0NE18LbcmtdfORyMn8GCF5ResNBdHofXdKJz3rZr9E7fPZJlXlDqnQtn/NMcgCZhqbt6mKjfOdJ
sQG+xSAugDctOoHEyBa30ftBQmChNonFMISYyfEKdVTCY+oLWNYrH1Y955zcPuUqWCKXqgxZcnZy
nn1oy5lYKkmj3+QX0re6Rl1Ply5FIQqvWfOzrckcal1geviboh6ky+4povYjfVOb2IavBkR3aVW+
tuERosc5vYRZQsUqqXKK9CNedM3MQiOSwr/LCPnpweindttnU1RAU9Yc6rsVkvm8hqWPqPwurvcW
3fTivhBf2fuJ3G8x9iRuYQQRDbe5bnOvlmAlDr9aJ6VTtjpgCkm0reY81MglA1N2kjiwODQQblSN
qMaobgV4ya4PAUw6r9MKWSBNilo+SbscCU422zfb7APAZHsIuA+cgCx+0g4aVihZbQUAzLuKt0Zd
r/BHolbRpORHZZq4nEpuZ0kMr6svqVKp/ufzCg4ivIwDdIUejRR1CjgGSZOmb2dPve3LPDWlprYh
x7dY7JHQdyQ2RKvtZF4tleZFtVvMzqhXGzv0yGH+aVNpDD3ebAiPgBJQWmMXM6KJ+qnzuhSRvyIs
nz8sDWLn3YDtR+w7yM2xne6q9CGVB6/kRQdDeqbQ7+DrVCOUknWA5dK+HII9ZevKfq7o3btZwzya
af5Z3Fw7XeZWV2Xn7A3OGLcGlYE65bfvt8Yg5WQRiOjmw2iXX69i0OfhscN2JUFqsYobjAzjyqI6
6HYNai+qVgSy54EjNf5RjulAKlB2EwwCXXPM/WS+ttlmNGVrf8FVC+/I3BWLkSuNxMIVaFAEaOth
XcXX8OOeHMMjh7hesatJiCnxjoH3o5xRuFZnus5H06J/SJrDmC5d48rkauoLslAE/ayzDw2qx5qM
ssHyZlB3V3AywHikKyDu/9VG1hfbsxH7rJxBsi+zFVo4tJxgpm0mOk9/THBrXn4/VV4wQ490qYc1
LBm1zMSGBZpCs8nhAgTFPbpV/HmteNLE5JhFdI269D4vPmBlnbscS2TJRa009jNEG9Eq0TJh3Sad
JSscedvTWWpCFy418a7rgI0sZ7rZqLIwXONl1/TZtIEPDaf8GbtATXiDH5/6a7NkEgEAwe+2uVyZ
pkxDXdrQLxurggUSGlQWrFQMMUG5EPwy48JQbQ5oScbP1eLUQ2cPbCtpcxAW+go4M9xegh6HCXaa
APuBcpyCDVi+XM8de3617W0CiBe4OsULhhAzxJ2tcqVss/RSw5NstbDI3Pd9vBDhBftzutfHjd6W
UJZ/bixsMy0zx4pz1dF53chPhcQCyPsDtYmjqrXfvWn465JWYJksxC7Zu/xgbl3g+0i3D/5CQ3pC
MXgKkddXveTosA6f9Dy8F8xgiqMkP+Z3huC6KQpg3Pk4zfIUE903PKs9lFagQ7Wdk6zhZKUi5GVQ
xwWWeR3iMhwav4HaJQx8FXQ91q1ipZWjD7lzL/GVeNXoF2RRtua0zzG8O7VdcIz8PCJH/65HhflF
01chxkre13PmHgvfVhHvoJ+FIx0IQ/wArFcSRKsERteqLYlmLj5lJM4yBCtX/y4JFSZKif8nyPBj
P+06NxvtN4zxwU01imm0BTnw2RP+PCBZGY5nwyOcTQsNQa092iRmKWZNRe7x0VLPGJh4B/AorPqK
29wUa3IgmSXynWh2YD5ajMKGb7ioHC0vlPzSRHUbao2AybTsFdaAml8PZ37NNHqNULzPtnMyHfjh
uFhJhoaze2t6uC94exahcPSVO8UuFWayAuBXdrtRJgI8wnhkoc8yumLgWGOJMKMphkAJ/HzRXYRY
N6ORcy0X5Ps6rubsNV3/cgayJIbIC3gRGYFAAh8Ty7mvXKIW5ZCzB11MHSAlPQg9wwGz/AMIIMNe
Ee0UfRJSsK+2xW2Gvmzfc0bIxNW6H9/dC+o3fOsELTy/5gDXzWDKvApi4pj25cLr8InyHcwv6AE0
5GEUi+Cy7OIz6kvM9xGZH4Mtc4Z2m0Elf1kllviy/Iqz5suEgf5+8Z0aczKW/LmZnFwbL3SiJFUZ
9Ri/BzAA6K/BkPkaUj5x2bgb1819Ns74x0KjvqqQBORCHlQMYTJraeSf2dzlzgjJZlJnr8LYlpje
/0dC6kR3NB/Ny8d36OlC0JwysnHM0KlWVdKNh/0UGb8vHJjngJK3KxrP6Ec0rhcBXOlaiCGP46hE
N8rqX6w1TGa/chO0X2/CNf5nFpXWi8Qvm+rZvdYN2LSnyubXa5xLkl9noscfNszwg/uAxtrlDw86
c0djZmDGFM0VVFVCcGabhTAUfH7hzjh7/H/sbZg1zcgtYhwx17cvuS+KUW4MWw5iJsRhLv09HmkR
HbwjsUPTXw3SMwZ2Fv3OoYp3pvhVnyzoUVw15PJCK0W4zjzcERcnyX0H6oijjTm0Y5kn9XE5s6hl
+pVWrRam+u5sEvZXi8Ehkr+3RhgjTRV8dCU8mwX9lEdlhCBuNZpUphDSf/Beq0Da+lxLusGd40TU
tFtJiIfAbVBdoWJLNbbVp8Gizxuv5KeJRhRWcXAGcSyuywmTBYuMtbX4DyLafbGrzo9v09gB+4fN
rFr1N8xjf1iWPU4U6fd2URStghy8QhiXP2nklMNx3YgN62QN1cTgClMqxt87TFsScbOWjS2TX4Mh
f2bKMg/kP+MWNRPXvz6mlIi8BgIJaG+0UW4iSkUVxKRwMp4DjwvgQCcirVEjLT5s2xfHInENkvAF
2namWU0Xw+F74Rt3qJD5qr/pAks3E99r7k0k2UufFo3ZMfMtm6/p1dNe3xd2F37bY2WvBe6LLNK5
RhMzuz7rBddUVuS4y2yI2Q/f1wQpM8FFGixiLOearKsRAJURqvwsczJCcuhW3k5UttFLtlFL59Vr
X8E2hqQSWMiV2uMryXQJe9+t+lSctmsPgYe8QBSghWFHkVZuqLKNKZ7AZ7kpXKeUEMsGyKLaZW4k
S63cfdgqfWzQ8WfMuvgIYjy25gR1Fwmt/amJngY045yZX01vwtXK1AVI4tPa7F3x/N1UUa7H7i8h
Q+HFYSQEpaWSHbbObPXfY0XG+7t5NUuRfxANxS5GzT4iDYEYDwo9hIC1+w8Q9FuVWvrNuelLQr+E
l7uMVlv9s+oCLt2F1wgH48uVRJC9F8GLPYRwNBVbALBVQcKCZpCwvBhttCiuyoyGYuZdPQcpMXCI
MNsZpHmEPbSF5wuFZ0ryVVlE5WWVbXMK4OhDte2wOEFBH4D18TbuQnWQhAjWgzxvOA/6JJz9YpaN
S9J53+JDuZkZiVbgbb7sOecob6TD1yBRT4X1Xtv676dJFS70PuZMbG96BkT5c5kr6g+/sOEFWwN5
Ral41Hx2N4+ng4f31wHzmBwTE1HllSFfhDtHNM3bIl62BQcxgylaJonOB2b1AaWo4aKKwCjCoRI6
TTso5jqhfwVLyhDwvsx8TI2ZaVPymhbdKRPXayTq7MTEZ7YOFgHzY1CHEO+ycxX9ByL+3Q6t2/Sy
I5wxdn7JKtI+ZsCrN5m1mcEjZCD1gQTdW1/nhBSR8SzfJJBZz6i2AHP3bNmlrJlNtC53gc7O72IQ
LeXGa7VFMXC0u9Rf4Rud6rDQLhCQ91tqnFSPfALtw38X2PKvvIXgLWtrWwT9IAEX9Z06rjCVRynJ
sy/hJLvXdTiRIcT2ItpB3gS+3bKbEiS5dBvlogo3C9p+LZLYzK6JU7MYVUvEtVueT92hXrI2oUVC
yE2LRClYOokFBJrK07MmkZ46QYKQrcybq1benGn81ntDUjDN0muRIQedUvz79JZNSXn6xoy0iU4f
oNOl0HKderGFy0wvTu3Sl/e+rT0irbiysD+toSPhYUbhGCPapEuTvZ/l9atjI9x4uNaMJ6W4U5fO
5b+9qEZUqW08IUtIyfilLVjBZl6ba+NgfDx5Sjx25n9gmPetYLXLEveQxZndOEpPXgrNrPBoRXSA
og6BWmjMFJwbplFqIJTtSz1PKB/eCy3iAqiIlzo8enJ71kpc9EMFdBPm/wF4/oAXaSYHY6v3/7v6
IxORKihN5WO8GZYR+FVBTo9bxuJb4DgQSHqqZ6rgt+2q4ME6nqQvDIQUdy0SjHXp58FZb7Dw4nFH
MlzyRlBZGtzg/Aqm0YMlAf4XszepTzN44FHCtYw7aaV7DaOIgPBkQClXqak9Ox64hWP18UBpk2v5
aZgQmlFjCLGj7ron+ZwrSlI7NobCkSDS7JD8MVyspdtVin5F/c83H+78Vlzjedjvzl/LEn/zJ8Cj
q0j61aRpaGHgQYrVMnKbB79yqqeBXNG4BZAYapUXgNlefdDYvQD7aaYIFNB160/KcMRmqj3fcEiE
GEXvatV5BXB2IoyVH4uL21ZQoiOAHkpF8onSZDsd+SEdlpcIuk4mZBGNd8cWIfQOBJbrSukMl4Je
ScUmzsfawGP2Xpk3w6ZEgpPuv6BPU3KIUtpWfyYTAjwoF7U4/+FsF+aiqxjOSfU3KnPYKAmYNsTC
7lU/jlHiwyWntq2HIVOEgAJsEh4sdlHmdhxgXTyUWvoPKBaVgZmeT8OXJR8gGMcCjcwxBtKcE02g
dSb67cGc4+TTpqjLtPdEO/9D6zj0YmNGLO2k6OrqAJh190C7Yv13R9QoSKHbiAHXHEPBbdzTvcfN
HGOG4Sc8cPCcAIrO68SXvjGk5o9e4BCh/ttFP/ESDP7cubthznBP+QcC2pGLXqClmW6XAFBmEKL7
5zxKj9LwquY3weoUYV7YKNJHy8UElYg20iHiHI6oSrk0lYcqgtUIjHM/VJhE/hpfdXE9DQnDguE6
OvTwnGiDjv+t+wvhOdefNQ+qbYHtUGNJj150EU1ivj0ewOt/kk1cXQwT3rPAiSdn7P3e3ylbkr3g
uIdVXDmmeA7+ShDvsTxTZo4WAziLiJeL/yoaAJZpGyPwbnklph+C6c1jV5+y5ayfBurlW0ai9O2+
jGfQH+eeaSpEgSahGScQR9wFh607l2ABg0JRdLWrcgHyHg2W7Rw3o5lkFlGcf83a3rlXABTu5J+i
yUlBGwjhOd0S+tnzlDiTQj5zSPOLJRHUvwnKBIabJR6S38+ixVZQutAJsYNOakgIbUbXGd20t6zw
lKQJl5UwsNMn//uDxKuzwJkVGl4NYx5ZVZA/yUI6YD+d9KbuCUixxkwbVz6V/59VhGQ66qIlsH8o
cpjZxWYTaxyBBHv6ZkXyYKCc9PRdLzv8BGHFS5eCDm0N9tBsWAV7p6lVfTpR308G1sekE4X7y69A
jGbEMZko/f7e8offKXuiabqwFD27EP2pJ4aj1wvHGMS+Su9KCcPB6uTwo0r5AVcD436P/C6D1vy7
Qfla8Aw3biF+HkTwQpF440Yj3zUvSanMjoo0sU2GlRv+gYGTrgStLh2YBuUrt8v3V40fjBuSovJY
YsFBcdrLcgjS3WBORBFy4KjP1gGi+i9yzqJUnrWx8IcF96bczFhknO5y5zV89AvVBkC/Osc57O3y
2k2bifMWUkpbr4kMTQq8v9G6iaohAlTLu/ZfJerxmf3kpLyAvAqOtzDDf7IHyeZML/x2U91etPj2
ywSLMAvrr2AWWnf1v9kX/UhiZM0OTI4BP17fQE0tlzfV3UoIeg465dhyrlQSA9n8/u80KZirGLsw
gNh3cI5u1qfEsWPS+WYMu2U6gaRxO6loF0zjz3Ju2ZTcc1BeV2P6F9kSR1h7HR6C1ZqiEg/JxOqq
dbQJ90l7xtmbd9eBCXGZBVmdWHfBFDtAE7YTdH4EcuS5iA9BxkZvgNHnleLu7eWvL1TfHS7rg6tw
se9XLn5SdLuSO8dIqgBMAiuQxwc9LvZQoQAxU5LOtzU7p+7N454OOwlGYuCROsu4xm8FtcFKlXmZ
HZaHG1HD8DCBL8tVc0+Wzjc32ElABTsD3LPPt4WGRbOtJ4m9WOb6ijWNkJCztValHKOyHM/EWeir
ZgLTRJm4Yxg52tAJOaxtRPd4TMYq2MqZvvWM4KhW8aOIkza23se6cHThQwF6EJ0RvS9kzSSpaCNg
7QBzeadiOW5Xsw3DYY7q7wvwUwHWZm7KTIj4mBKEugN7/u/QVBpoVxTUoNBkFp0mskcIgKfeQ6Y5
cfOzTH6A5O91Jf6v4Gr5hLiUqj/OHV7xAMvWks+/EdU4xU+CxfNKqu9Wa0iUP+GhsIvt3mA20JNt
IBTSySWdp1URodgpK+mBPeRDrzSJyO4z7as60ahm3mToTDvck6nx193R+GXvfu6rzWxCtKZDamZy
KTbxtZRR64igL+QM8Z2CbohNDwWQJr+SeoyrJBEobp0LColmCXhuu/QYir+tB6xsPdu5PEUSglqb
2EHgslhtiODFzqYknNcsxQp1nD6z9mb6nbuIUMSC22QL4UE1acwlgalX1UeIJPjEnmjZ9NsdCNVI
csvBfqOmOjDJdtwIlevAlGOiz46ntbcS+uP0Hs9EgeH3SbccV2tOoIVP66cSj68vJWGW7iKzawo7
iLW9qZVQw2bbXC358Nf9C1FwFccF+6Re4t6TxmqnmyW6R1+eguYfvdEVwnz0yfrCdi4UKGWR6VWd
KLFDrG1ARPhp2gK+Hw8sfASoAAF01m/jC9mFRLxMhmrPK0TLAdRKCE21DoAs7mGSLcqGJ4/w5CSr
UABn9tRz7gg25BCdp1IOwzuFR07KbZjQBF4I1ErvYg1mDMgLHez2Y7Y+f9gSMbtVuFX42LWu5Blo
ylKrBJ/wr6GUik1GK7oHthYz1OstVgzXuhyO2nFzi3v1/9aBMiwTNc/Cq0CdayhXqtxFzAtEQmkV
KGoyJzfRA+nRyz/Ow+YJVKIjZK476o8xNQoCEdTTikRX3SUMBcqsIiMRE0lTcPc0t35Bj5q5+cTY
9Whqnc+cA6BS/6eWgV6Akub0ExW8uAT77h3cI6W3Ddac2ktAI1ah9cEC7UK8w6tNa8013dF8pGvS
QPZfrA7mDRciJSNVDGXtvZVFAMvnQZI9DZCCelERRnyGqxHEWUZTmPOgRy8GPqKoEkJfyzfxqCMO
hOGxpeJmONWB6KYieUtEh8kLGVJ/iUXwhvBxq19M9oJtPy6eMAnkLMfSplT328pJLhtulp6leRKj
RQZSvNrcBJmGy9AQ1CKbneyyHBkx4bpMjodcoiuuj6UBvAZJ0PkNVd8ewED1idNbTfmfFbDzokcW
/L4Gp88zGzaZP5pc0YpBXxUCthN5ExcH/9AkO+WdbKUzHT1p2zVE+mVYfVTSW1LQUCL7iqiw2XDE
c5eFbkHh5JWXom/iQrAbXVgHFblvxc/T1u/5sXsvps0ASIb2fbEmGt2Mz5CqSpFCEI+6AeFY3ZbI
aiG5Xn3cIFwERq6wcWOU2v5HhDQeFxBLwB6uXhJ4YWaN088MIUHPzSCAqEcoSPxJgfXF62vHQEu+
C0aGCUtNfZq2LmRXHy+32psDpikCmReT8IOL+zHHglXH/s7MPKUAyj87WmZ+o0bQu/q4Zh7Btu68
19XKgIfTQOcYxyqRs6mWVElQz+2fFn8BIPE72moFhu2t5zTQGDvUuavWuO4bJziNc7mFW4uunIhu
2XdDKaZeN7ZU2lH91OtV1KZMw+fBVb7V6WDVsnPzk3pTRqyuDMBmXKFCnNXj/76x8ATGlHcPxfj1
KZmRCyUXf9eMC2nSgh4HxerHflrXuUYvyJtgkcUS0Xt0CL3fsBHyMRiWDl/iP8UoVZh/xTCZyJtT
mcBycTGtyUBVxvWzwMM3LR/IM5VIqqgvVNfxnfH3rH3aL/EmJV/f/ayhtB7pXfbRt6ZYLBBDY60c
pJYwg/ozoIeH3OOeyGK61Sezk7BaZyfaNw10KvV2Ax4Njjtem+B8fngR2i9qkFMXWAJNet84c9Qr
V9Jncs4LHHdoy6wnCzczW/i5BxLrz5PMmZvhmMPieHRGo23Is42Oh4fWncXemi7r4PyYwfxHV6qU
q93cov4w7vg4LKgwWdiztp/7MWhKvwy8r259GuzHaFRVaWE3FPlx+CAM7dtrNoLzXyp35LWcBHby
dIDoSvZ1mNSwVAg3j2h+djhwNhOaHP/v2ABPu6rvJXu1Lo6KCrToOtZvQgKVF1yLvMj8IZ0+X9Cw
RcW3MUb5BF5v9LuwVa6dDw0wHka4G5/K5zdSrvAd7l0ia3oDDQAge2Mah+kmXxFRbL8azI5SKIm2
bcGEQAeZheL0zsLUQze8mFL0ptGKwP84zsrE0DoxPBKbinexFo5NgTAQG4EEMA8KvFsHtd/lE4GB
coxU/Fzs+hOgtVqFZWeFwHwgi4p+QBQKOmgfn8KX0cTMzaZ3Y9LfjXTSYjghhb50yozV6cJez5Yn
d0sKtvCv83+9U0pkz7CM5taVFWB58zmiIzhXJKrWPLcZy+n1B0XKbGDhk4B8GvFEaOwFjtBFwBfK
LgG1XtZGx+LmsLbhzONGqatRKs9XvLeP9ulVIwGiYT78fsbWgnpuG+ISE1rGuC0pozLqzJEZsw5g
wIDsRr0yjXTP70T8N0QRYHfLx+7VAJneZBkoH2W60emfob3YV5EUchUGZHob6tsSk5STKXjOvZ8z
FZ/j5rXA1y1bnIaPRgXXLQwB8RxuqNjUYCpa1hMd9eoRYNHn0Z9SSsTampLqFG+4ydBmWfLIa/wR
8zfsXz+2FHeDGjPJLahVVquH6hssjlHFu01JoDLRT02tTSV1rQbATQiLQoilpWHz9AbJNosQ4fHd
Nn4Bq25Sm9mallI4O6Sg9dlu/uM88HDXyx3A1XUykvnOG0BOPnuXdQwjB/mhmsodWIMxq9r5Q2JR
e+Joe1tw3J6CPv5KgKNx/CxBhe1MintX0MdLyQ4XZviMDD4yWYxOrsefSI1/PC9clsvNVcfJ6j2U
E6IxSxGvf/T+qa2aqHG0CWjc/DYjxwoezwWFLZ/2v5v4RPZVo2DRBMUYk8H/z+FqfQoIBbm7vK5N
FAGqoM98vDG657rElIa/QwHDrcIkY7ZVntQwXRtJgUdtLpTFI8a4n91jbDeskzSBZyaoe98lG9t1
B2jFyIi1m/ninPJ+kHeBog8F4CSokX1816vdDe5RXA5glbrjvOujPFExN8gcGOLHx0Lwnp/tTHah
wJPWO+v8DiM2u0GKHRox3ChIOFZ8T7ISwlcvybleSWS0PQIGCLR8yzj09KLyzGtJVET9jRshxDfg
WRIU/2NTIkuv5ARrBYSZ7hXLfGIIFcGZK4eCjrIPlafoseVKnyyA0u/05UMWqdfkyrbJKZFB8zS1
jJUCFR8iif8gyCYfg+bY5g2SVWCqpMObNmIgmh4yBJwr4xOGiIBqNYnwzaApqMIF+UNCEqwNeWhS
/zFlYTgUS6o1ykAojXxf7CeGCu7FFh0QRsXtIjdkSTxPEWGeaymNHpTCBLwuDVsmn2QRvCpRXWsJ
bk/pCHDjPCDoG6BOSUj0UDb4Gn4O1NAcnT8QlsggGBGf+lL9cLnKsOIzfihbfOqwuy41nXdkSTCg
ZcldouyJpE4oV9l4aMoEPYYqPc5jJ7G5OxfU+460LBCXrcllMJ2ZG97kuQ8oelTRMCAWBFhIe7qX
FFnvYh3z9VBhfRc6MXpqYGYLCVINJhVfkfnw6bDm8EffYknGFSuzpR3EC/hLk8okIFAJLBzRyuAs
5XlnSA8+V6vS0whvv4/6VaIeO8fikk4RIPK61EsN6gRGh9Bjdf38CUVDdWJT15gQPx0DNY9uarto
d73AuH2A9vO7d0ouE9iFtkOuH/u+8vzuX/73EgPV8nxy3zozsZDKDkbqtpwbQRInSeZYxEsPHV54
ZT1dvci9/DzA/HbALZG0BeQbL0EBgz0wm+/iFrd/ipT92JOlN/wDwjrO8z2E74hQaHvw5Vnq9tCx
rMWNIzh6hddkyJVO5ww6s0WeENgZLz//iaZm9hKTzRU/r0AZVNJvP8Ilqo2gTnr3xRTZJfcYIEgC
NV5IKLFEE69zom/tnAwkwfGi/rCw0m+c5Budr9AZ3luHb6ydW47+L9xne0SuE2Umjk30FsUr+M5v
MfVVCRrom5Wi3gpGEJlEHNRp+5BVZVAMm14oAv8nAw1Qk7xsi+Xi+oGrj4V+9fbjs47XvsnHEDQV
mY13msp7sKhqtYNyz0bsJq2+aJbIaxbaCr3c9+mZX2PSLPSWgNbltt1cmQNvGAjkb6nMHqLS7YNx
/d9yjty/1zupy+PNd07oGI6JUTVIqWVzO5lywnLOSJZwUsjGxGWtvv/4NxekN+GQigGAKXchFdMT
dsvDdaZn2NsTsloYoJ74V/+PxbUjB66tuHc8ifQONdsizlGRG60mU+ctbHeHrCi4qN02WyO4g0ZH
NNu+TnOoBqQgliIsWgJ6aXqGAwaPpkTCe4zV3pyfLJ+ULrYHPuXbgMJvkLzkAdA17ssEgQXE1oSP
4pOWsMstWs0VYWzcIL2h4Obm/Vgqy1T7aGW/RquEC9jHD+kwgKJIvEj9buR91qvF5mkgRYfIm185
o2m1e8EUQeaiLQp2+gVQPg3pR6WYIXmlQh0tZsVQr60o97lQzyLpeDD9JmHAHCcQkAt4xWG77TFB
Gfr1fB7v5JFK+gBvu9DeV214JIkbcL65OBUiIEq79QQoGTH1/oFS61xNNnSCNhSFefcCIb0UqZ6u
6TYl2g5b99S1G1FaRQuElrz44u3kzSAw1oXbgfIMfzw1Fm4Qjsw/alxVaIiM8pyX4+1+x5tUjUTz
czqUN00YnpQQWZaoiy11IseHzgrY49utT+yNyJNFDeiUTgbQDPJHsjgSbE4pQdhQe4H50XRmuIC+
XTv2mIzWl+JAv5f7nzO7tr1M4I/VZLJME6WME/eBFXWIK8JUTUUMYwAB5fVjR7X9rmXSoOcETv7l
NpxqWQ3cOd77skePLqkt4/jivmYFI5EgWwz2Vk8e4lR7610yRf0ZMCMY4eILYDY0aJIzCUTqnSvD
ubmw1onyZT+5Qbc6yRMsucLUEkb0OvhTigUJybSWXAAfxQC5XTNf5GIykPU5mxRlvgNECmdopjUv
FxJTH043H9U19l4xlD9WaHWnhFv6jD56C9+4ZGgipJlCKKYK5fVRuRSvxK53fzMDlPBuDJpZoRKo
ugIWeWqPYrMbMeiQuo/tnt2MhHUTnOYP28uEb5koI30qtV5Z1l+MSmPIKOINxkdKs5VmWLMWNBcG
OD3Tsg3E6aNyREj24WmjdUDW2gwb5Z9Wv4z1UAch1lFbDQPW+Jz4c8rD74tzCTF/WGR+Fb8mD9bt
D5irK21FFACX3KmK53heja7AImgJfMIq9+C1dH0Pc0eXWEKuBIZhPs226EvKHgS5MSGoU3gdIJzh
p998KjnsynRCnMtZz2tQiuNfGmfxNuOeJhyykwt1CJmDqfFDIGBIT4nUJ8DpAwYJqoSHb/tnyqTk
JKznBd8axM1wVPovDKxkElgv3Dln4CpNtV+TFnE30Biy88qY9wgxPlyOPaWYChFTAU+A3lhzgaIm
pMmKbckwD4PmtPc8Q7uGXPQdq3IO3lermlZGfUc2Eyap6z7ElBeqYFxVwMrol9LEGUBu4HstME0u
7ugk549l/+FzgIEnUk5VbrgSpSVlsluNIC0L7FeglIlZHW3wbcTlAjhyLnA/CFkCCBrgY3S6zGK8
RJoWCRJzS6+gIr+CPjOkmgBcR4ubEc8AECztwTdu8JGHrbJaNEH19PgOGBYxyb9UzdNvh8C6P/jG
b8WGLjP7ZAsoZpqF7v0D4ggVt59IGteLV0e7lOkP/1cutG+heCCQSleFLqy0HjMoSl9Xl3YcyNqA
O2DmIcQqO8RYSpoh581xqM3XN6OoKd7obitdufO/UHnMAR6gObIgfSJDTmMIIvR2LMZK/cuXruCk
M4UKP+T3T6Y05UHNEvVCJ4Ir+BALWqBPNm1tdj23hTrvGHXD2WpwxYrTb3HbcxwVi7KOxzQC8Kap
8OWvuXfqA9R+ltVirYXf1LDjjUUVUzN4EuMWW/IhirTAixGXOUS8h5RyX/CtvkphXgxG2SeOhojs
AQfvRUQlfysW5ndw6YLa/t+Zi05vHhqz4fzJf8EWeFE6BVYcYzlOJc2xh1rZa8tA0OJgTReUlQ9x
A+cV5vdDu982WpwDFawBK7/J3VBkY6TZVh8hWDgCuvIGlv/aWCh32TbOv9GlcCcDmdcfUW990DpS
Cj27AUGZ/sVT/8rbLK8e8aMG41wpZzP8GCzM7faUbgmDhy/diA8KqXiCny0/kFa6HgYafFQHBix8
uzKOixNfhToQqe5XFFv3jRWL4QfMXdllXHGwJ65YAxPvfKnUFowfj/xSIzAnJMau5VFsW+Nl2L8t
VubcibfvEY25xj4+9YuQTMJr17PrnoX4FNZVWVXCdI5m0Q4+n0rpt0nic8lNg1eifYU/Q1h01aws
9stK5unKfWE/QNt3I4vME85HA+FosEIsw7lqT9z7hi8uPOj7ihVt47McXD3eQCT8y+rTtqBHY6J3
XnPG69YO7OcVTDTgAd/FQ+CeIBRsF0kuKR9oJ+MQlCRfk4ceYMKfdOct+J6Jved5F9r4/+2+I96Y
RxzSkheW8BWjmXWkkSa01TXTEFN+1c4EKYxhshbgV3nlw1R/XmOQVdHT83akJ8MKfm3T3Az+RbhG
VDPMjQ1yh0cvbvn0IWChBt2yvY5bv8ljZvlNZ8BJ9Q8T/MAP/0jwllezEv7xrPQHlkBt3s1m3wvU
iXXMZjucfTAj7SwCD5gS7l5UCNnDHxuiyc8Oz3drlCsfnqog685/GIpLrqMNs9s8f5F/RzP3/osc
0Xvd6pnFY96nvLumZ3k9VT240Ova2vV99Xk4uYkGZF1KFg/+8LF2NIEyqLkYOeJ3MIb1/C2TpwTo
QMWCHufBEOp2xwy6OlZ9N9Kp0Ch6csmXqG3ebIJp6bes7oJ77+4cNCXsXDIrJMmjuy940DgTpWaz
DCIEKaG5A9kBe5vBbcCrfLmM1H7SZ5k579xTYAo96rIloBUtpTCYNo+OCBZx30F36pZSIXf92fOw
rWAMTgPc53YkNV+xPFvvczHPccgxx42VSJYCO7ysGc1XJplOKqCbS3GQXc/Hnw2+VZSf2kHRCVSY
rja2rBmASVs4CK/WetxLFIPLt2KpA7vFg4a2dbqKHCov9RDIy9vAgdxjk0kvB02VhZHx36lTtJUf
qHeE8VkomZaofHAD0AeWGMCttGvLPFwaiNuFzIU7Hf9fTnlbsdN2fkmPJpwg+qg99JKfGVS3bfcu
OzSnBNdm0wpHXJluMrtp0EZuR+YLbi1thzkEpNHuHB6OFl81UGE5YYglwK5MrO5Wnympyrvsqn4a
LsWHxiVtPKtTg6sU1Ouir1+2ww/9qkkYOnhKGXqLmx/6rdfws8d1DnZvFJqVQd37JmzNH7jXswRe
OLw6rab4zmg+OEsLIEWKTVxngGltbIbuOcTY8jqghvMYIUE/li2WGme79oU//aVKZG9J7ZXIzWrH
ucF7SIZ2Hk8FnO2yuKcRNX7PoWxbA/nZCgv45Alj4RRfrpr8Th/sxwd0hJ4yf0Jdh5jaHjgEsDrx
UZM8Co9OsdeSjmI8pokcV/7kMlO0vpSJkaCRdzu7zeiJSwsL6+FM3PL2hcUHnyZLifCy+LN2zXeg
bT30Xwwbzp/b04Bj9b7QKBymC3cwByZXw6A8fEqEkGqgTz8ik5TwyE8dz+YILimS9GbF7zHZpVKw
MFvWBKt0rInC3h1609kHZ8/KFG3WYqS96PBCVns3dasd59LTvRSNcCPUU/XHt/PoyIIzszzuUoH+
v4pRvoDbhvwk5bG9DIP81PDf6g54IyzFcDVWO1Av9Zo7EYzHJznnTOI0WjrWXfmJuxZ3JrGG28mP
ymdFJTcNU2jKRS1svtiix4RBnS1M/XbDbj7za4aFVbjDGG0sxoJn5s1Cb2jVB0Onkb0SyI5hQNXq
JmIyNO8mb3bK4mscFA0JvwQE3hHHCtq4/EAIT5VnC+3FPfaoew+chAe+Q3rNCUdTSKd69oPbgLuG
VtlNtFXFDm7Ypzrh8faCzDKcnrYn9GzaBx/eyHOwrHHmwh9uZai5lDi9Q8dLt/SW57YCUvNBhxnu
essZdPOPFpGFYCkGGp3AcJDPlbB/y91X0BQ0ly9Ba+LNmW95FmwmzUS9XaGK0ODT3wgtTlAFIKBz
CClt56mIeP8PDJOS+JLPhp5jJn4ksoaHl+FwJUo7SqSY/EkHP4lL78HUY2m1EhgzVztOei5rEB4O
JVvJKKWRa4E4MKBqEkQPhZqDL61byC2NWceUNiYmsRGfhQ7y/7wa/laoOLbKOZbFoVmVDd8GHZyO
GCK93Yrh74pIQbaXxlFoYBveyaADGvqLBQ+FsOAB3l3ZYIvbgCcPwjZLdURH6g2jfnOUVO/jXJJM
gd3gAlKLcpCH/emgDYzZ/bT/t85WNXqsW+VdB8pTE89fIbznYAjHNECL5ZBprtVeHaWCNCprDvSQ
FM9TNGU/T2VxXUAIjjnubuGfCXphee8m7CRA0Zeq/DV23+b+QXJIMUT4cquv9zUEshf4JW6ZzWaj
VxG9BsxtupiJ9vt/EkE32N9IYTMrP7jEorQ/XRzfN/RngMOA1CceZKaQlHFleusa1gervWwih5LT
Ixm7Muw8flQe9kt6cpwtVGUNmejrVZkU7a0Mlzry4I2utp7T+amNAe4gu080EHW9+cC2MkIBuHap
7JydKV1tFpWkv48I4IK7dbVARS8pf/9l5hyY6ZjL1I0doGLSJnSfDmibQhv8um1iRrHoyBU5SdDj
VD4aPajG7ORaR9xhLJpeOSS2M0j/sf4DJin6pbbCEkY/a9wvceistbE9KLjjsnmnK5qfxVbFoEn7
2qMJwQbZh5j7Lkd/81/WM7K5G9FPOKCxHyqhJ5IfMQ9v3IN8Sm3wi/o3i1UNneH8BJWCPFMxnSU1
mQk+r2rTNlUzgzxC/p4oaLCCRE6vfDrnbvw35OvyMSAljVJkxzsbFiKzAQvS1cqpCG48oB7dLB+X
NJ5br+gEIla2Bolf5OAcNT0MGyuQ3zWUwYDZR2i0c9WJPCQkggOiF/dhh+PGWP6Db2cBYsrfbH8K
9hi4i9HB5IVy4qrVdj6Niz6WqNuARK4Fc4dIvvo5JegAXIXjhr9r87y6WFY5zu5cv4rkUnvmg5un
RuSQ3Etujr048bxWWzNw4dinK+dEVCm+5/6ko1FcBGlILvZFMUUnvRQnu3hqIRW/j95RAkJue3ch
JVzT1YQYjBtX8dwP+gx8Zow0SN72r2YPS4wPXVJEv0Lo4qK777h2WwbS5ol35vxu9e+wbU/vePi2
1UNj7DWkhzWKRRXOXT7AZkcLnG0Xnk1aSjcqlGN7OJlUl/fwQNezNSHWmPAz+yi1vaQklLNzxIe3
CD/OZaOl1Cxb/Gm74M+AHbplOyYOe627kHYgmP5xgtpk+btdWitSNPdkX4DBGoZQ0TV7gxAzaDUj
gvPnmt5EjAmMYCjsmjKFdKrA8GrnPtZ8cq/W0eB68/JdbBl4yOUGiQKv2JEW0aV0jid9Vk7j50CV
Ye+5IJTSVcaIAKMJ28X1Eif+c2+2x6PoYoRpLCe5yQfa7e6azz4pWkG9MQFrHWQ60Ct/3KPJcMEW
pAmuPLJkpaiyvBgKSKVK/jcvuHGpQsBVPjHDMDMi/1cYu4zbF5ZVP/uQZC552lQTRbch2Jf5EgGv
i5uM1nLU7Y6Idvmdc84sXv0aiX5vwv07FYVKa7wANmJ8kvE3sn3bls+VMkkVQIvII2hY06lv0mnX
b01Kz32459zMiGWIazFDSB47dEyjN3ZNwAUKu6sg39U1ieTIOi16QBoyh0T6pKOCAStRvSEttPA4
8oTKdjCRHs4x0h7dEueuw4ToqeDwrPOXV9oULuMh/URBJ36tRwNfpdHjBhcYtj0zUjnw0Ih/tzRE
jybrFur4MdJ8wIHeS2zgxbZlKdZt9+k5jxw8htQCbzhGlARloCoOChXVtAgn2/0ZQNpAdR7YAeWB
J9ZU4ogocJK8V/GZ6K4K+npVSPpoKnyRkTxn6vMc+XCXLIRJKNdx6suXD5AqGfS6GtAYd5L6FXh7
eD4+w0BrCK9LzuuPHDJsL8XkhenwndexNpI/RIz7b/eutrlNsb6EhywHWuLTS0I3rQ9ApGebUszE
F+LSPDc3vNIcw43MOoc6XnB+ynJiranxC88y9L43dTXC8rsOTrxZYnbsSTeG89hxBr5f7jjnZH8X
bIpp/QtvDj15RdPM8rAipZ+9RaYGWEElZHfpVt72nAUpbIlPdj33ajrW8Rke3//KMUkzCZBeFCFC
ayTyr//7WpY8Q/Paddx3bTdt7uB/KnDxX4WDkvscMb74F4d4hyLJmOQrTj/uWwY4P5XXNpKT0p0I
vsyFEAWJx8jUJGaDDM25ev/1izHLQIjRJcPetXbt4xImpLWpXXiY8X/QX3iOWfHR4Tf2Z3MSyOeX
/8y+SadvdVmcDfTbJIBbIz07QMvvQ8uvjxlA8f2r2MdymXpYokWxay1A20ZBIibng01eECIXMNep
AX2YKJwsRoWLsRtBN6+wxeo3k+/gNuGIekcoMVEIGMZbVyzcukYHve3ChYMu++D1GRt7wslc5t/L
rVmNOtTbyTwgTn4gAKD2XFHxMGX0fOWMRie74Dtvm0/j3TO3mZ/O57EZNtf/znyuhndS6lTnWRwH
26/4yTbxCunwOq62N0kzLrgiXqOFtEJtIAC0Eq/dBZqokYLI9ZpV1nlVDe1p2jRKo6MD+6RgblI4
h+BxepFz2RXNsJoBjwZrSsUZzsRJ46crLnXh46OEHW5plS2y30upryY367SWdOSv7GLDYcttgvc7
2/M3F2N/sPsommKsOo9mQOC1uGFNlvus11pYthhND2wgw4OKqV03oQCSWvk0xT5IGqPcJ/5cCAmw
Y2F8LKEKP25+oCf0OdtZTd+az8dlZWHpUmXchLmXgLe1S2HIr4VLcSgS3kk5oJMHtC3LsyfvoQxO
Vdgb92SQr/Ygi7bOderooiFnlQRpe6lGl34HbRSVnQAkjCJdxKOQuef5hdg/1f4Yy43txROLWvHk
z1altbeXCnHYtYAd+zaAdObwfYNgcFXumltpO5udOLg3QoNoSEn5bsOWKUkdlC3w2o+1VPy7PX2X
hytTMhu+GFCcG0osB/G+E434X23q4O9eOZK6wmOV5Xb6Ji0Gu1BixDuh+rzrvV0TqvYakUv+QaxJ
zuZOmZmhQOtwrTe3NpEc+1hdXG6ivNL9bpSVCZX22iP4f56BhjGzkdKl2G0KVUl4r/BThRuQ1yDq
heUpa3JOQJk7yUMJFykaQ3xRKewgrd0D2Zrg7FVgclQ+qQZSphMSz9HgZND0zdYDpKXK29BfBUZI
pqo/4iwKM9sikvlQGZpqZRUCqK+tgau9mbDGwBJbHXpcK8nX0by1xLlrDbyZ0xaFI9q+Xx9ZTOj4
FqL3M2qI/H9pgRpEOHbTJQV7uuNs/a/CsdPuTIY5R22JA23PIjIejoyRSuxqaUzN3ivO/eXzNI9z
1bOKv6mMwVppGDCXywI0vuIt7tffeiy4aXN41rSEY8XxEfwEUvz+wwIemxh5pBbCbiBUnPxPHRjm
kuPQWp0hWmEzdH237/JB0j9v+98lzBx8OhoPYxq1kVMcEZCC4WU/0kWq4q2fJKfV16iu3INFD7oe
nj9lN8K6MK0NPCydNg0fLpqXgJerXyjGEXv4F12QsAgywxzaUkR25DR+ondT5oHwkytYMo9tcjh+
xo58Z4jsl6M12HpJfdTSy2bIu5G3jcfM1Sy6zFTqZW9NJCEUxaQHu2VAFjEq+hOu8KNGS/l6wg/5
ja4KOv6o6IVUohg7oLeZssaiv/g1WnVmS4IhqFEqBRNdGXX/TIHlg4u82eJP8HvqR4X+VqVsOwMc
MmAngTcyYeAn5zSDwgag+9YeKgRXP7/3GGq81Qs9wUVOcl0Z3UzWv16JK5adTjAFq14Lv1vZlNAf
DgUnwYScDAFuXPKUs1o9MF4RSAxTnK+mWvAyoLc/ttZrBJVcQpJez3LRHWs9GTfy9IQlqS6EU4zP
9iQSDWL++jKS5227w8PX2+8SfORx43q/n1LUYj/NgnBWixPfFHUcDqjzdNh0Mw37dvnYxZ9ciQsL
6EdYZiyNb5VOOiz3ZxQbOFAwezP4Yt0vfi2koNlsFebkuRLum4jjzHrc0GajLpXOAqtslHsxOtFz
URs7uOgqs+U9oqn4Nt0VbHlENG+YvuF77z+IExoh8ziOV3x2u4xS7tElwLbXma+F+HqiMrdTgLW6
+F91vGGoyjseydNtjowztEf6OcmEf0lGU5LBTn8Zj2insVqnYK+CZx3xUTkEdduo595Y2X4Sye/b
ho+ArcJK9C+Dl10YFXDYPQeqoNKKqhEr463ngoKeFFrUC/YJKb+clJW+2mZJwfyR9LnOFy1Y8fOW
/yjnpXEBUC0uvfylc7WydUW2Jn36XkWlwEytyYhp3GyT2fDzXIc/Kc+12LeEI75y7ByI7eY5JXvj
A4PC+XawyLdHfEjlhEmt5bA1dSIzHDe02mG2TDmZilgvr8+m8fWxvnhntKKBfraJYb6uS65mS37T
vWa1/p3aYZ1hl9lwTsGvAtCbwwKqAWsrVSKLv5MaY6ZlJlxiM0ExbBmv7tB0s72LNxl0c/OeW9hV
VxIgVVUBKg5tLHEI/yjCtQER495uiKubHWi0tA+MmRsfUgRPU353F3ESPSlJCfrdaBfSmBJGwreX
Id3o4w3b4/qXX3lbaV65G+KiwzDhLE/YzPAnNvDke0JubWm86bjF4PCOTinuE2Pehbd8ZDNHa07x
o2tu+N4kElg1h0f4gcseUj007MKnllb67MRdMRSbwb1gHPPec+5klpu2Nwz69vEikR6dRwtuWShF
xQWMCMYwBBqkM0ovdmoic5d6GDCwdIL682tw6JbY6IoZZUCR/ZaaZfDbej2bTBY29fFsxZHX50D+
EGJAE39/c+cv9bwriwLcUtOPTzSUt3CyKg4nqn0e/JWfHyuWAoqseh4a+e9LWJNPqhAM8WUZgB4f
c85u6IbiuRivdo71F2dOJAd7TcQcdHUJq75mY6EOUKa8ulhh4/XHqcDIY5p+EDPB4gxPO7kO3yuc
Wi0yQbW+CeRL9s1Ht3L8Pdfo0140On2lhzLQTXZ3QDjQwwDPbaWugwBxbkeSPIzUjlXBLCH+/xsf
wEO+LzxAl0t54FFkMfhKvZ8GmuvJ48WSQV9ec1774GNYGZzZWNaEMWCaTw502EZ6XvBmbUtPBn3V
S62IodZOUd+p3L8AZl2NbYg2E0lYv1EAssoLLa7z02MQb6NPPVh0lbDIEQ03wV6o9nMJyRS0T7Ch
R6gEgSe+OZGusHGxgv7lZ361XXCrUFCwfcWLh6bt4EIaoQ2c+XazXoXLXxzV3nVKXbFQkhMovfNs
aEmmNz8h364q/uaE6bHsJGTrjvHA5JQyh3ULf1MMfmuOWuV5HIYpzdDEQxDPgMoyvoC1O1fmOpD7
naoaH4IH/aVlh9N1qJBFFe10Y+1874dfdzAEh2OklSA6tKzokvEMLEcGNRzOBZaMuleSHwBY9b8K
09z7KAI4UXlaDMyZYcmGe1zCKFUxDVCueYX3ws/QVlNeZBYcf2VU0xmhoq8KhNjTFInVfxeVNKK2
SKyHqgqdmt3yBZ3miJdgPh1yjrl0V18UM23BwGPNQHevMg7RCmIm2UKKv5XSsLDVm/2+WG6AxiDi
gzX9BOU5fygJRwvUBNTzPXCEq6cJWbGrFS11Uo3Xqs1pK9RdgTcHOeZNxY53Hrh5CVOVJNfCKCE4
DoOd2WmjEky3L6z5ooIPXadZIzTVvFNO8LaZUiAdgi/SXb2TLnR8NIPf1IUpNOMKDqpsjl265hCL
O8AgiJ7N5GCBvOvOGlOMSYSvbR7Iw0BxjGUGOoZfoadJ9Syjlg29kdGL73hCbjurE1cLyZKTlw3Y
ojrN9JiYDssWGGd+J8HnxOsfZ1vfyCmP61NSp6hxnVx5sm4dtzl7ranwb6tQBAgHdauNobGLrd4t
0KvVYGEmW4ZkB+n0ezEnw6dtzoEbKT3/+sV8vVDXLGJ7VbeeIc/qQfQUfUyiTCwrGJPay5HXLSAY
ElI+iNUYFoijfU3tmGW072xYFWYIepnIP5UNRTDalAvMBnHyT4/qQPAlzeq8h19FlKRHuAo1bJ8b
C45THCTD7qIded7j28v3Fk43qrEVEGElt/3YgIzppoutW1uIKqMsUyTal0BF7BFfY6CFDQTqOnUh
qZeduE+XYSE167ElQFOs4CL6zax5ZULyuP42wPL0x0+f2/v0VTgRnpScI0uDDZ7iLlzp4ltW8nYL
QyL9LoD78ZIkYiUEP0MwKe27ct95ae52qAAtESwyevCEhq1zjVbD4zVSeHD5j4H960ESwMn5bpcA
v2zPSpncfqpneN/yqJN0VkcP/Rt7PsX62tojeTZ5+rOHntmmlE27zZqKVwTDnHHjvNOhI2TpjtEp
43P7NTsOx+TUusaugAl/4hnQvAM8x5gkPp753Fdmjn0NRkHkLBXeUDluSUoVxo5iO6u4P81jCoDU
ygU14murFdMTt+CtRrTGwoTxMwsll1FO10T8kWJXXbYaSLw62G/ys8gFpkk7xicOlMpC89xT5sTa
+VkLUEhbCHIQ0JGCEdu8vC+D9WyAA+8kjZSJ4jHikcqSct6GYzWdu05xCBFLpbB12YDcsacz47BQ
wqMonLDrIYwl6sp/A6o/CCYUDNWExAylPGwNoNv3qvFIrep92jNY+KtdMIHNGtIa9YP1/62u4a4B
f9OUKlNQNRrl70f3Tgeml+4Y3eIlUNkRBp/C3QHz2BtpfN4Ac9Cls098IFmNpfJIz/kxS7TFaWds
QvvVkfJaUzWRuoYw4cwPTTbFOCfK2WwuGjny2Wo8KLBFmq25IYaSgkUboVuy0dJ2TsJa6rzl5+gq
OrMOr7taU6LC7sqafToyE3cnnclLIIkTPhLpa+/C2mVFDCz45av1BHK1r1+aOeVTZJc9YP1eMBid
oyUaQKIm5vc1MpJoHlYA1EUkp7lAdsqdZrEGSlzVbZjAVhh7daExtLYVl+Dm6XdHGZPiEx/uFb5a
ExCFwIEfILxCP0zGkKhPHEKz+V2UomrNmNZqF9fQImei5U8UKdZ6ApDIyDwwHptx4vfhx8KHz1D8
aKXvkTqgeV+ltEzuR1TY2R2cGtn+KYEFBdMIkGmVhnlwtTY0Y/CCmNsXprxTOM+tXiKGjzbzd7om
Z7tnt85CnJmeozLdxK9XVMOLM/+UoaV37JU71z3ek01MWRZyahnrkcK7/x3tGvjE58+5Na00/nyo
TniWz4lI2ZfFJ+8UFjKEYbP1JyQNGcl/M9UJSlDsk52xVWV1iYgLrhB4Tu6bsVMWeMMjhPyUth1Q
lwDg+7DoNs7W4e8y6S6RwIxlheBweSbmNDJQib/HDsBpgrJkpJyyh+pabEJYFdj9InKcLeMbwEsW
9aL3IUfwvln0QjkcXYFHzZkdww6/mAyNqhsh+YVT6/XsLf5/J1iJ+g7/GDwapp2RRmtCUohU0WF2
cbugxsDLfo4TSh1chy/ftTpltSvZ6deIlAh3boyMBcvc0sltPgdJBR+Jj9syn9QLC2GY4n3fZsr5
31jdLFppFkJObrNcjkrQoT3ItoXBGFSQ8kIEvXd4a4B4ytkS3pMfP+0OnjP0VAW8/iS6xPDGDr48
f6t2hzIQJw949GkbTPFyBZLmrljWmaw05HDVe+2Tpfc4G5q0q995TgVlOqtUgn/iqy68+8wxerFu
gsiXIpgBXMy5rY6DW8xjXMns1gKNaFJoaljMbc9OzwFd8H8WkJ4oX6DQ3yMqHHm2VfRbdjywNdKj
Xl65j7bPD/OYDgvKxeZ4LtdpNdosX13Fw6xLYBCtomSLWHMGoYiWYeU3b3vzt54OhvZ31r9XyFki
MCaE9HRARqboFeRJl4kmvForEmBSPH6b4j+37+jZMA+8K5xWF3Zcd+c1ckSK8KvOOufsMDY5WOTx
Bgey7pro51CKwuI2z+9OLNhshzmOPzpAW64qCrfaAm7u4hl9NamJ5blXS2S/HO6fYmYh8pOj+LdS
7C6t+d3Ns55qlK6xpY2knZzgAAgkTiQF2K4JFbuc0CU7dsZlCp4KyQT6BbB9lRpedLRCk+uEqve5
9JfKKCgOJoK8PEiojdMr4v+D2Z0PqZtf1Cmj0R0Ikp4+3HiVffzyRRAyuyOx6kevs12yLr4WGzVa
yo02KAtaMaoB1LBQ6MT5Gry5z0MRNQ+/9JvWSK1bwV5m0NivKIMRgroq+hLmlAw5VduwepdosW70
5/JBvVsbRz2AyP040/5egQvjo40QvT4BtMowUTJ1XDeVXfPxOqk+gOCFd4GRHB4tUPKha1cPIAKN
bdZUDePQMqLUkJcpTef8++Outiz5rz0V5PGIlS6VyANIiMYh5FFTCgdf+1ciEfBlrT0FwLyGFNgP
rr/dFDpWr+F20VAFebcVqgpsFJd8mtIXkFPKnHha8edYNBS2RZ6Tl1l+y49GDH9D4urLyCd/iT8g
gopjeD9/i9Y6HN9Ga36OWYS+3pi/bfwWUz+U+o4kYLnF2q0+MszBExZSjKwVNMqIT8GLJ05dg4im
2NpvEY+tzYWL2y0hPspeN9sPKBPJRsyYImPMpcn3cgMS2e7rrYwPgJUI+QdOuNWWxN43buaJZPl1
JQZrmVlOQUG6aP3d4GlgUcY8pnvuoCvV38osJeV0k0ySQHBwUCQGYR5ZN0jAa/pg+4Y+qe+igxi3
M599TYCToo7p1lTbNO0DevrlhpN1NDiTQP/LLx/o3PCmJ70qbt6AQ6olEqEOvCJjzHuzDrOpQQhK
VuCApoEgfswgzTJQILCcw8B0RCJDJerJVC8VIq+h8i2fzUv5NKR8sqAhLp6d0rUYFf02sviKdd+5
sZqbZJlxFqJ5wS9dcEf3hjRbPjhDfbygKYKFjDd0QtAPZS4I8CO46zvpUj5WDXIy4GvXhM0vdZZ0
VFpdiRMQOd6gx9Pn9pGVG2PfK61vJaSF6S7pOQF6dnE/wR4OouCspRIMX/xhhI0PtdUSF5xllXRx
BTPVdKN/Zvny+VwQbSVMY/2NN25D+7ZK+3hfyrjcJeX1ThVMQFz7icTbydt6p8UnYAj372Sq98hC
7zXJacTn3kIMmo1Hml6PXLSySa2krDL5t3hrk+Sc087mrNN3kRgaOTO1+ICuU04Z/JzjYJE8YmdP
lM799G81qc6qZHnHFP+6hjAzlMHCTfJSga+an8rEYUj2pjASNV23GeyzslyMiOm+3XAtuEy80sKr
cu9KP43pClkVAUuF4hka6Iy2uy6hPw38sGnIZdtDJfA1CY379Zx4CmbqjhKaQKQs3+Pfmv/qjL64
TWx5tYsWpb12qzIhH5xnbfh2vp4TpaFfPT9Z0hOY81N/obJqqAq9NiKimAAvORIqqVyfNIS/SPeu
xh3cZbbPHRFx+uKJDce4/jhTFJDGhxJMEAyVwRGjy2Jx07ktWFjULRoSnwiwojfQiTWlmA1vYQgh
ClSUqGwZ2+ODnAmpfkAVdsZgXlxVrVh4Zl4+NphzEERKH094yWHO4eo2n5BVNLtOkVU4ozkNSEsw
22ChQOfJM9UMb1KB0NmwPwP6uGtmzZVrkG4ZH7zL95IfZehybrQsWAUCVmqUZMnajvnXLR809hnN
WLZgyW5NXAqtnXPXYwMYo0M/JsnvpnU13YyUL8SnyvXawiCrlVmQU0NMkwebZu7mRvuEDdJqgYmS
zPIqIEO9B5toav52qmwSGpejZZAF9mlXsxwri2chMgXgZge7ZKvpNQdu5iIjJQbMYeUD4jnuqIfz
uKzkbERpmgck+FyFCEu0nYZH8msoobVbtb5LkfY0uMBd3RJigyZBMnlUI5Z+4AKPoratE9OtjFoN
3FRnxhARDXGY03Ll3jH3Y4REoSefl0pjUGiDPZSGeksSdGdSmkwhH27sb6+8x8ZaSDraIAbIY0UF
pEB0125b63f3xbjYBXa2lahKuJB5NnOdllcvKVhtT5MXPO/bW0AfA0tDvMF3ae2qTlkwoyczz+F2
IE+DFQQqyg4J++cyiuknNKLtU35yvgiT2FXlKMBM0+jCb9HBeBTrZ2y2ZrygzBpT42FAraQt/02g
rXISBD3tKTWODd7gBcrhrP7XD9tmKk6LDImYoS/NnAoRWlIZJ3eI25L7bC1wWeXmOisBH+jvCNJn
vA+rgB8XHxnYwDlVly1kuO3AHCHE5MpFJJUo7eIHkzcb/OGrTmss8x335hBT7mH7BjcLw4kOrvoM
v/tAjcZF4eQnYkkSmT3EcAoAsak6SoSJ37ZDYp1XQcM3MlLHdJScA0oJhVtXprdq5lA03aLqIsLo
D7M4uNewkH9YKZEqX9Iv8GEP/MEp36wDWj/O4sOs49eN4eYWjvkeheqwAbaCyxSZKqUWZIjUdMhh
x4U62ystdhCH6PFZJVjC+vO2X92z9s9LbnBz3TQzgqFoj+0V2a0Sn3anIzxnUTGbvDzSTobmNRF3
91TiyaNMEu5RQ2en9t4ue9RoRwJrIGsfRjsZ7QbeqhRrrQMSrJh6qR0V32ZZDGa1XrpPHthkkEnU
En4P1Yi4PmxSMbzbfam2ovQirswMw5t9jDVVn9/2rZiXmj+Vz9bspPJpl21Cg5mcPVqM/fq0ATwf
rjX2shATmzMP3RBq3zZ3t6cJuSRa+FxvaE2mG9cP/U8cKAoS0IR3v3Eddq6td/wX5vrM3uX2cXBc
5+J29HHHxL0NmtJbLGuO0kCRArrSIGO6MQOac3IoVFpy3fnZGB15z6aGyv65Iy/7QemORGxqZty6
9wSgjxP3yXTRu5XMwqh7aG8W3wog72vbywjvbVKEqpw2qhJgSd6KasJYIYUnPnPd+MsP8Z3jNBse
sjhK2hgqPmbnSyvERYQg4ixEW+/nqw95Uv97b5qQ7Nb64JMBydMTLBF6Ak1MHZM/zWKhq95t+8BL
WSxiOdfUNjkGxQt7x/YVWfaU6z60QueKP4bK/LObgBZg767VQMtgwiPqQUSiNBmoaNEBlC/3hhi8
B45sS/yJAktcQh8qyqDDIUWfkvCpllTqiCRgJG03H4P9reZH6MIaY2Q+N9uKhvx3emD8Mm9DIwWD
7xZEAfkeZGcig+dcjiAOfk7EiCQFMFnzZDOeSk1GDB24YqRdsLYJVDa4X4C0iTKb7Si6CqSl/goB
yhcAQPvA12K8GyJZSuBML7QK+C017mt8fbydg7U9Kv5Q9Un6IZG2s1as2vkFgY0MeMjURTJt8MHZ
kf+9LzXrCrfns47Iaw0MMlugDvQeUSbSHY7a/Yn2lvb59ryaURgxSjr38TyM6kX2PsuC2sytj6e0
OUoEUs386ERy2pRJa84hq8NzCshiA9240GVj2AX9g3IOMtXD/2u4K5+F2+RV/81eZbGqVcLNEkxL
AtUqcPfu7dPxfzK7l+UvNUUDEsrS4USTGE8IKwat84QMHERc8UOLAAhxNortlw7p4u1zRFpi7ket
G/r+N1VTf26JyuBwwW5QmxHVu1mK7FMcDywRJDreR9I0ZMV01KsYIABDbYcqiI4Z0NwlE7J4m5dA
GFwx87kz7H6vOMi0kUYiurVV13T5dT5Ab5NdBVSeSXCSrLFUpVLlH9FJrEGEf6Wd1JVtYrwv42XT
QxE0FzZse7S9AjZukgspvxMWgVc4GBPyrVCGjLrDB8Y3WmPOQUesrz+WJB3y2XAIfCpUmiVVWvAF
Nk055zqVoWLUVWmyjvdpraHbpOibBv1T1z2zpdfKCNPMEIrUrSR272jxozdvCxhQ3a8ArAD5ko3i
ZstwCD2R1M4W+tfx1wbR1/SUfNp5Sc/J7pVju4Kwldj47TjJiekHVHqXfMN2ulmmhnpRMMAXk3RU
o+ldGoqTkL9RvIeigY0elH132dYlG0ATmcoOMZY7EmA4L6qvzMxzn7F3jVs0ee+ny5iHFGmCmDsH
dukKICs+mKBFIV2crrYh40VYahfy2mgtsGW7CyAE02YLa41gtFi4lS+q7JlM5uYqGW5FW38CCyi+
aMFpEDzAIjD5v7kg38jiHEjnsmW1AZYTakehMZaNskp6JGLpGt7b+kmvJfKmeG7nFlLS+c44Ia6y
x83Ui6FH5k/eVNWjVpWZdHE6sLu5TvLfR4IvJb6cod2XNo9gsiedwYenx+XhfcigWnBemBHOCW/I
qt91nOumLYFXxk1S7mkh3K6zJxS4xA19ZgaTkhmFRy1EIL1y1m4zRhVO247rpUqteLe700d2f7vK
ZB8OqCdI4mPt9kGY4kjcx2ANzGQesO42ZdtLz38Ma3Qw4jk7j2Klu2XLoMCdvI7nQVsYGWk7fJ4n
RhgzZb/TwkLODLDj2K7gDsYepv7EfunluBG0NnE8hA15IzgbjMC6wCnmIc3EisCTY+aunkE3yuNs
adnjRz26LiZQy+GmebLIT9hEB6oai4IEl5he62rO5ONAKXswy5Ys/X2r849muqLXfwI+RmWS53t5
G4Cd3yJnaafI6BkigRBJ4KGmjooc0gmn1ks3DMqF5uniCxA66pukIuFRkKigOHXlqcNLepR0kCTD
r4NdN2aSKQbyK2S9UhFjOswHfTGkJB8EGQmPOFiDMXdbqJJmSv7vCaKs118kbKyPOmZomxYVNQ9j
nY5POv2tIpujF/ZmE3AM2pxtlkx5UmGcDjnd242MN8UIqicZghPOrxsnSRN/K+mFq1tLPc6ESH/i
IuoBOsBl/OTsTFj6qtsxqYakfIisnW84UcGn4yexxANH98gNPG1FcfbRm6OcT9RHS1aB8ikejvs8
5J+6FOBMTYvMYhwhXYlnLsuld1yGDAPduaB7kvf3Ra+gqrmNYr5QjzEpfBqUCMROInleH7qc1h/V
861qK2kIs0tH+xC4Jp+lkxoMLFyCH0ZoqUBvOTc0xKAbkSpLL6CpaD7pU9W/1M2LdZXUXqgdXGyl
DLa/uR0qfJMHXz5dF6fQjwL2iudtdgZnw3jHHU2ouI77kBK3TO743wNzsH36L1gHw/Xsi/D0y8BW
SERYsHq3oHOxgwap/aZiDQnSASf8jmgZ6Bh/IPZOnNSdT86Bemt3nQK6Ttt2DUGBOtxq9Vajy5or
c2VzLBhOBwkhbgIesRQa/l8erODgIakM3svW/5sjPMQq5DkgfaDt/svQxdHqoeCOwEA7H2DRiWi4
wlY57zN2G4z4AULeJnT9RReB2F2KwN/c33rPR1cO22Lqt2SBu8lXEcbp6IUcQjJRvIyMLFMYK7bN
i6TiBf63WtZQJFcrA7IIZ69/R2ANAHeDNlJke6NNxivCRgfV39vAEIy+Mkcz61ETMAphDU2q7kTC
xFtLB1o4NXircMgBydiFWHbO2HfczVaU0ch/No0WdgmS9o2UQPKqHM16VW0ffPCap6Lsf/MjXDIN
bff/zp0Q5m8979gxq9Lc04CTIlDQFWXiwu5G6vLLo1opsflPcauy2vv2uZefXCG0NEpAGJeicZUV
tFNHBx2ITqhQgnIMG1QnvQ9hm7daoouvC6dhseI+H6lash1PwU3/i7Nonc1eSCXa1QIF7LwcWsVA
Qm7TKTWY02fd2bpGtTeLK7mYcQJKaeIzulsxx1w9hsLfJCCwItSqTFpmN82rEOjvoUp/HN80jD51
y9y+e7cHl3EjypR612cgegxEGHyKvdjh6jLSlrKP1sJRGBAMFaeRM1BOdS/V9yaafxj3+SLK3A+F
dEMNaJw5QEODrYB7nJ/zJ1QpQDTX9EK0RubGF9cEZfq9kdhIAlsEUGToPI87S3ulSI3xWDFOyfY2
IZnDuV2gwHlA1i7vvNGvYt7VkdthOzwkjHERr87o7OcpsvBlbog3mWjOOHmpWY2AsyCIRsQOiysO
qx0jIeQcn1e0OxrNp7Ti22gN5w8ng53ff92GBt5rvtw0vDvLE6JGpJ+qYuHtvlRadDGJtT5MsXO+
NcKg/ZMDlR6KfTbHHG3xopXIHTfPKTOt8ld+lDy+9nTi9N+mfapgDOXC8SWtC9zLBYXK7dABVuLH
q5egGesC2UDNKFGbrdFCzh7EyLBatY30TH5rDRi/ETFEM9CbAULrxUWi6aktMi5zUONTWj9mm2Au
L5+PxQ/zMy6aQAVc61p1JJ39xxvZzHs4GN1/PCQtKqot97Kedr/XAdFQCFrACcSqVingS5bFimrJ
C750zjZu/Jm5rZ3GCT7GX/kiwhg+hYSw1H0BtNA9H4JgC/iazCyWEWUtmo31pRcrZ+ssThJWTSIZ
S2zDYN3nUmqw3XJG/SnNpFFZx4mNuJQvyYAPzSELQXteKR1IR+mUWJg6tHHEkP+cChuCNNV54A/q
6GT3/n9yisHLtcJWfheP6rCFNysl/wqex+m7A99uYBJIBnzhHk/+1pXByJvC3xV+a6wERv19Abfb
ZDeJL9zd5lY4SoUk9RA71mvOin5MA96fbdr7YFhU0SCsBIi3zQz6SBALzrmz2a9dEypg+W1Xrmbe
GZ5v3YaIecJnJeEjrfLCkV4XgbQ0MZIxnJkDjTcKH7wdJ4vcvrk4Gig2fO9QbuCWiB90Vg934271
BUDdOvYLWdxYE0r+v8SeeYXtob5zGDLG9XXs0fm6zOvavACZL5jXzt1n199BYSG61je1Ak4Av+io
p4yP+vRAmzosqkHSP8K1gUKErGWoeTmifySoOc6Sqgu4I59J0TFHQ0EZIefyU6b9rFkm4JOPgrA6
xbw79TVic3G+Cj5HcF1yrizJEFX5zPKbfnTKvCcUtO8E32MhPoErlLt05UJ7FYhqaZmHpTwTZ1Qt
m0MrJFzWPtN/b1+7LFAFSQTJv5zfrXuqFbEXCKo1bFQMqkS9X4jgm8NrudJFQM+vDEZi4DqeOYnY
9j4Df4nYPUl1b//xEywYvJ894FKcSLWIXXsHSaAPHskRalXQ6eJbrQilBsAnTjh5wW9nw6fu7lPT
w/uhdCKm53FMYYurkwzRO5gdWEkzdzMO7987HeRoLLx3+tw8yAgbQJa/2FEJPgro0ukRXLvr4a8z
WMGbN63/MZHJXggK0XZQLXo+DqH8oasTR3Ye5bNNagj9YHC1Lk4S3dFw1fTeSDKx6h+gFxIp3TaM
K3JT+cL0UIJ+AZhm5sxSTQPNVP977swpw4BmXQnQ2QtglnPjd7wn7j5egvJf+kgzqshsZ4sBoObi
cRM7fOB7ouVraBqenptvEWDkDsBQEmbNpeNQ7U8H75aEx5/hTku19qSPfvXT3v6zvLTWv26vNaf1
fSp9RBdMxe8WU3BUzfK2O6Q5uBc2Gspm8wN0uPUr33fj2yDb5ZpjqR/Z5uogndmGURZU2QXtBD39
eOnLHyM1TtIuJ42hlun9JusGInjf+EihBc9q+fcgSLbsYf5dATryQV+e0G8P75+TV0a24NAFVyXW
kDxdvyaFzwNw7/DbWBbfELE/6EeqYaCRfAo4nLDMc59gYfjop/B7xRLLF/tiZfn4rxf5fptgHssb
R+yzRuGEj9/9E5cTFN1/eNN5bVbgT5njgGs8canZtkd7leb8drYc5AkAp3KARYUjqAFnz+iWqBrM
Lurtz/9fiJtsrzhmohWEFrgmGXLVGZig0SMUlCAk+OkQlw2XjXdgPShBAmt/WzofJX3oXt6aDOTB
XBJZMhMR61qYzvAqHS4M2O7DQEC2XN+A2q9NBdAQbU8kdyW7UD6Dmp/XljdURI58Ztg3h6jHOAMK
w/uXyrWSuEc/2P9rC2FdQPNnR5WBuIc6Z9ZEYKOryop0X4xuHLz05mNvoomrF+oqaa7Y/dhrD+dF
iFwh9+1F2CKPG4ARX/sSPLA/PxlzFtQH0e5eK/mEe3wP72WqR3lb8tLoA15b4i+nhSWgKU7WdAr3
FlJH6usugXnJ+b1yY0BXUnuC8S8fkHy9qV2ZdArqt+TVVkcLZ3GJBiG78PxHsHf+plE+Kp8svjJs
rfeprdoATfllkml4Q6BDt164l3s/2sBNwAzaxuppneNy85ciGU0r3dEVjnhdzxHySDsszQTcLlC8
2BsJoDdr7HJaCtoG0e+zVayZUvJiEDZeklY9tNhZeRBQfWxJ7U/LBUDP05fynYVgV4tfZLghgYC0
B8+EPlgtU/cCSyq7p8GtpMv2Fu4ZbaCfFY2/OPKlecMiZZr++KazpW1FikoH1ilUrast/Ml0rSm9
lIBJCNdb8NWbz4eobGqrYc0rs5QKrtVaLW27qh/jyc6V7/gtAOnmltRMnwbPvgnQBjpUwHUWj/yD
ENIKPAT1JPPsQPGEXHtdybHDkfH7vfg8WN+l1uI8eZcksPgSebeSO1zFvhu969c5UELHc5ElMJL/
opdiR5cUXgxbMz/zG66/RIiJQdJ5BE89h33Y4PoAowz7EyRVlcrVe2uu2coieu4lIZ0XOWuqaDYE
ceFHF/RPvE+zn/+Ic584fi2B51hQn7aWK5TZ+0EdMlSFw1Pvb7EgpWu1UGYSNiOUCgpJQ6BXWPVm
6XuRHBXDPzg9xHDkQuZHm0Sn9p9w+GLIkRMRkw+2kV8Q05oeBLlWwLYJZF9r6oiX1SHLTYJzzR+/
rLbQmOa4Tt8vv6FjlY5drHumPyxSypI4cJT77LOe+Nm7v6JiO9xtSlcnXaeSrghCZC0JlWOHRSix
REKqPCokeKAHd/VIcJ7VkgzBb2UAfQ176iwN6nM0YQ5qMXadNLS6oXad9UXs2rkKQnzX2paDWhmB
C0U6RcoVGcAFNUf3la5saE3ITSeUDbpBhBI3eFhe3gtyw6ka/afstx2hyM6zvkl/MjnbYKpQUZBB
wDVfHwXuQNtPhBBSZWYoQLVExnkoDccL15/o6QwXv4RBAQr4GIQAsurNuNCmMr4ZuCC+6FN0bfhK
3b6u2IeuGBWy0pT2Y8ML4P4W0B87U0S7xqFnh2zTPmHaGS+eUCkth36vcBe4yrdZPt8pGOoT6yOZ
q6MMOO94W+RFadQdg/xP4bRTAvGmilRCLMqJ2GpFCDPK5/+ZLBPl7HeHFAPw4C93wnijKJw/+pkW
YUNaeViQvviKXerl8yhk5rGTrNZl/cRZ+/d7xlsPcuE0C9jvkxIBvem/JrYJy5XnfYsZJGoFSUgU
jiisGCCVDV1kI499UEh3OiB4zr0GrzmqAmwEMdROSr/7JItKy+zhILtZr+45DJnwNo6wL3fD1YLR
OnK4E98FhmXEZvtLprH0YFEChbK9yngdFC/Rm+7eTfQsfJzkuYVmMV2Fcx7iIp9lkelrKFeEbGMd
mZx8zRu1nQHwx2IkVlDk6xdRw0sIqU/hZmvRld88OfF2SsFmeoBW5yz3nwh9JyYYEQJBDzf0agS4
g3VeOuKznTIaymGejhyPCDqP1MCeWgm6ZNAUWfCJOTfnjbFVuUscPlwVEAdahwYLEX0mD+JXDI0W
2Zi95ykJOo1aby0u+jhI/Z4RRovKPvnCDBIK+xWXN0Zw+tJJ6I8EpPg0gxVIRDVOceZw3KMh5i5k
kaw2e+eFyX11ZFe+w0y+rCzC/d8zgmg25Pd5oAqLONCJzqK5MNkJ/lkGj+xfuMlTCZJ0qYgojSOr
nRXAGliF6/NgOcHEnYd7RFpxGsJdnylh9/qqHCihdiqNCYQlq74Y5jq6Rp8kYuWtNQDBv2i2a8gR
Xzn5wyEYk6FH5sVQ/eZDrXPmar/L+Btvym9VHW5c9idVLITD9zJG3Edx5CwDgv2ADoaMCc9ce6xm
pxkNaJHi7m8P5LnDjFNJzP8FI4GZsPfJGeTdq0RsNTxnjHq1xcnRHZzoccxBkfjuQCL9xGrM2QxM
VMVlZxQO5sUqkyEfjOLCkiLNihDMDvGupjDk93QNiK5q3OGuX8exIYabu+NnvOYOoJKqCqotJfPp
ZeR60+LcSKtFZvLX2WJwle/1f49jwKFtG77Iuj6fnG/4IOoUlSqwvqVzyqYKyLgDqfuRdpEvqKfi
+KrykHsU5MwpuNe4WO26BPW3jKE0dzxu7+BzK6bY7i7jj4Grt01ZCJCugAimpyIEVOCB0v0qExTy
/zaVJ2HDNVwxh3MRdGquvf9VGt+AWJ/u2WaEkpszXAXHs+sBOpJL1qtss4g6xCq0bqlc0rpNTQX+
+AAm0bmJPjDTYgBBNb0mfGNMO+h5BgxVVPCpiNyrK+X6hrmpeRXzi9hdeomH3nY1zNF89hokpp7i
xC96MbhZTEn8oW+np29vwCMSaTH3a/1LGX7FBdjV7OrXk83lB1RWs/kcUWRyw5XGFjgvWrr0afMQ
5HZIMSthVpc0XGs8o8/kM+WJ/e0SRF7dAqp8UDUBxCmuh4Heo0BHkDk7ITTU9oyVp184you0egiw
McxdjrdIEOKV2olKC+qR44cpAbH2mpqCjTtuPmA8ftAbz+4xm2lT7CJuB0NkPs6iNQmCS3hh8Btz
8NqjcywqYdh7ksneaG5y5Lxr8tol5RI7eDcf4zDvL8WgbbgFdkr6iS40M9X+8lYXnWXI9lNujmuB
YkGqdgnsXWxnW13i5MZAKhduwryZja1fNBgUSld2rrCvFvcX1sSP8L4VxcNS+ZsL1ZDAMI5VeNio
1ufarMyTtsZPtOZf5UYaz0R+JTRCL0/Uo1BuSPAu6UC3Jmc8tRrDnqGztjtIIrwrm7XHpgYq2Qqm
RHwrZZH6Gn4jdTksMKRhygVjoVT1I90DyVwtrty8Waq/Ju7+9CKfdu9ZEhSzFOIBv1y7Y6TX7hFP
CdkbnF3qjeRTroSxxxR9Yx/1c1d94fYA7BWRLW2d+RegxmP9vxXflm892c5VhpghSyCGME0gCCw5
t9yYTzct9GeAKKY6CX13jSw84K9H8FnmNa1Ttl4JP7GXSORLEybpWzlDfCN0o9X7NDPBtzhhr3nR
oig7vOAT+pqXubU3iTb4P4Pf8v0wxMfUn0UrkksJTANzxED6hjexFFCNcfF4l1Fxn52MZWVMrcri
y5AR3v+oCDETu57oveRQ9maVXeOYlAjjVP9uTOqzrHoaEy/pB/+XkQSWqhhiulWJt/EbdVjHU9OJ
FLlzisgqkCSmRykSQDpYIfwOiLdgqU0LBEBfLTWk2M0TNXiSObMM0QZntSCeR4Vf9fcyhVrflxxL
EmDgGZQspt+j+E2pE/Ni+mGsKr+M/WeTnPyq1SecdCuD5bZr/2Ffr4AS4FvCeYzFXfRc9JUHroWh
cS1U/+t+JosBURVCWLlkdraeB9aTxmzTJeD4965oaXJj5kSo/Gj6jrYYsliIfbRTh5Ct04/g9Eo4
p+sciZVXbs5qOUsYpY5BlReZdsgEXhrq3B1rf1k7SOoS0TbA5hEbTfxSExHngKEknC+qC9scefLv
H92Vqcd/QaXbT7C9RfrFyP4mvF6G8d2Z/9heMAl6uODyaSG5jLM9v8pHfEZtKp90PSRh1hZGnG9v
G9sO6e3GMKJ+fogdvUBgXczfT0VyGtDhiJnzlL6NGU/L1+qN9jKAyur2r7u1KDjQfjrTWCuZb/AS
Cl/zn5gPC7vPPkVJdkpjWi5wT/wu8IeHWZQizlgOTZmridClyWw0c7ex8kvRY1042jDjo106XW9Q
uX1lLKuSnQsECGFtAtvbZLBvwocntQ2pHcpwKOMcEYSeiF0ZjwnAozK8BF+12svVZ01jjelxN2Fu
eZk6g8gS15hBBgAo22SD887G8ozqk/ijWJOOyy843CojdwoaT/2GBI0kacbEt0V0D/gT1c5vgOUl
feO9+KsVlFHUIV40qkypC5KjBn+GggR2vjggsIr1xfjYmdMkCvYr97Udo8XI6foQD+BV48EHXR4O
fWwJB40bBYp296Qo6FxwKUjZ4sBZ7fF1TsxyfUGuVFHoheLeFi7i0yu8WIfJTAwK2NKAO+sXC+kz
QTO5lt08MpZe6p0gloXSlNyMnOpHD01nMQ6YZG4HNKp42P6lRp5Q8+CEZ85Ks7oFhBdtvegpKwBl
hB1tTkgemGdvnb4rGHkEPqHFxoRBXavrYdsIN0YHDIgtQgfTd20BiBdDfI8WGxnAEP+Ni9W5TfdW
Ls/rhqbxOpMobinJLS1vZWBaoUSyWq/rHgZycwwA6whZcPEkRRFnT04CIEnS09yrM08FM3qD4ERU
s/ybLpEc2ear+nq/BrHi/JGNyKEfIuFRZBHqdBoSpE9XAqUDRMF4Ne7X+5GcCLbg0KzHfn/6c0h2
GrP1Pj45mwzD32MUT7Pqoklle6WXPf1XkMfVfbwd6KNsXrEhZpaE1RC/0Coq/Un+VrDOgxTn1qEs
nhsE9kLs3S3eP3q/IgEpviDBOZiJdArbrUn7m6hDFU1MYxUVvkiHFHcC9VNVCQrKm0qPRRqiiVRr
P9Gidz/AmSkutTseSX+gidzauonvIX1jYZkfdtL6boZvAjTVwjam8pabb87rK8rHHlmSZrEIHVrh
Zux5biWL8owYLiExNLWsfXGcIVQQ8L1JGaQVIUbGqTZUZBAPFx8X/csasR9Z7UiaF0DwKBMVj8q/
6HKguoGhjA1P1PJwV2Dj3/v60/uDG0nwJxae1oV0n+aR+3JsOIbKo5HUXwytdRdmFDCvTWgyAUGC
f5df36tInKXRiKdvMDBZdTptZltMbYAgqlM24Zl2D4TqLKARlYzN0GVzYa6oMYb/QbzZ3tYjv359
PR3BuwylUVgSPd12uTvSMxEbuY1nATs/25Gj0Mh5r0PYibrIdI0isHG4qCIHCS0Tn6adN/d01XQ8
fOhKvxb4KJBiPmUdhRI3zYeb5DW0tXfGuVX+ceKNuBjGhbqZtF4ubg5HN6nsDYYHTNnRfsdmMCBF
9BI+q/tvxySXPyWIyIuS1lv2Z3JbJ6IqSSbN5+yT1qgRDZSNp2eBomo5s7neC6fJKpz+Ww6dH0wN
N3cNO4F3Mc8L+oZ5kDC15yA5RGTpFxQdm9sUONchFhDUmEXMsQos+6k3x19LEVpVAUT4Zo58KSf3
8jrXtYT1DLAsNE0MB0q7KrFcyQSxbRTxEgxfITNJV6ZPvf879llrUT8lh5hqiyG9JnWXMlGFJnKz
WadX+HSbvqe/guOshhedxo9uBU9pzLs/DSPg9JOJ6i8W4y2TMlF9+d4JtVS2nGBSc93anaoMMIML
MNSEDJwcFVQ489NgB0E83vR+D7pOY3xXcbnZ0CIqNGup3f4fMj9nx78o4HYhD1zzHNkoHXbb19NC
S2WYClwWQTQ85Y0bFa8dUI/2XfZJZ/eE6xa4M3hQOVSqBFbhWpcxSOtymHbVVpn4uTQkTMaOYTg3
++9HnjWQIKdduKZGRL9yFeUXvObdorNSI0Q0/9phW4sd15+u6vjkrVeOTTrIKIDn1Z1wiqtGlf9A
DaY0/hO0YKdeU81lI1uxYT357LKXSRbUzupmSyEPJBtc/sGhX7x8OwBd7z+01awM4VinnHxB7p6X
+T1KQ7782MTj7F8EraE+rZTYCgaAnuXDooLLbLY5ug4zhlbAnmZKAElqRvQPiyh4jbFtOivP+M/e
e96fX31z/OWuBjzs1Qjdi5X1MrNA4lvyNTcq/NxsGtVNsl+GXQVl3Q7C9ad8kTsInXqMxDNS1ntj
HG3cwAuEMK5R5lC6CWAF/mqijs6j0V6eMxBdXOlZeMu8oV3PeXa5T30+kJFl9xtk1VNn4IbNCEib
zbloAzw7N+4dOjO3GHa8vQM1qKfm8/W0z6TfQz0apQN99b00TiikkoH96+0LNJoe/rgpnp26N/+Y
fuzain9LxHo4wRmzloDC5+YlTOiWe8HA41hF3bbtN6sIhGZJoIFVDw4axgBKgF0hwn1EBO4Sw8QM
ku6FhZ33aP8iq/4vZjR3zrH11R12A9NXbgteO/Tgr2GKfF3d6gsXhlyQHXVWjCKR5XWMMKzxSuq4
P0tmMsubac19dge9MSN7BC1XsSmLoz6n7iIsOHe6TuoG1Qe3RdqcDufMZIlrYoRAVv/RTBfDPwVL
OjlfPzTvqJQ/5UxN3+0B9b3LqlVocGaq84jTx8/o/rWlZHycZJDAjdXhiyuUwlKRBlKiH+G3UKtR
pxExFjCdvglUxz+NVmjzdil8RhpXH/y0q4LOqeMHvyXTGvyL05idXRV+bviFvJJUShj5HI9eNIWv
iWOGTGrmYqjDXQkteXMAiFwYtqE6ncjfIiXsQCgtOO80mDT8Z1GtZhdFaNajvjN8tEa3VkI3q2dq
qJapNmjMOm3MLruVmOFmJ24wD9zY5E5aEdO5DfxaQoYAfsUKF4CpJWXGTNAZnoLmtsEAJAFEAOk+
BXzNUnhhvebt4uSEMnUt9ZzlsA7m40JcZRnEqAzKTmZcjjFxjIge6QQiDgZHx2jxifIOoLNUobqk
ElghwqHkhPH2g2LAI2P7yii3+lmEXGvctCohmMH5CEnnSr2gxMmgYKp9eP7NKbmMfZbrl0qX9Kgr
StqVkZMpBpRat4XoskQCW3U3WKZFGPyjWk9WVBT6AM3y56spBRBaVod/fSepXlDfBUJ7M7sFS8zH
mpmnxq5WyaEpwA14iJJuMn1BN/HbBIYQz77OuTKMr9ctIi3xR+Cvv+pQKq0IXkeTPiCFsqd3r6Sb
R3T7MM2NuBbAeTT6H0gshdJ5za8dAE9wO15qdOp3bqVWSMiwGlc/V7l35+MfKOC/dN52DMRmhGyT
DFE9Dh/xC+wvk7fH6lr4AKD9/0UGvclCIJKhpozTHd2qu2ul4Iix2mulRws8Dqpy8J2egqf0cilv
1ZpRujHgGlA4S84jXmw49BMPentoOvHZGeegD5Aoyh5+9DTxjK3VuzL3Ey360gcbmq0tVLwZLPkn
a4SblEhr/4MSuDvKTmGwdMh6JCbHcbApN/uaCaZdPanH+gUiMd6kLptcDx6gUN3WCDKC9LIfm4DO
3EBUmLy7tnJRjfiZvLPbaAI1Gutw5Am9Mzau5M/uw0wKBYCLm9xgbHngXmpaGSvkpxACol64MS3k
2MpyCaMRFa/daRCfTyB0pw15BJPWDBwLX6dOJnWUlMNDnm1VtXePwu2Ws6rXrJnM72xlbGJjJg0V
sBRP8pEASQ4/VbIHX0xPayIRE4OLIzhT1C8DgFR2qGoGVFSN+bMAMFNrt2eqF6Q6I+dfzI1CjVzS
14epGg9UImRlSHfpZrOzxpCegYBKuByK5O12tEintJ6rl87J8Tv2yfy9kkyx2KTmr4NcCemQZHqi
4ks62bTMA0m5ON5cws8bqsYvQ0ZGOeStgS8MWwxi/na++nJ1RFnSc2pDU6FsyDAuJPM60c6dqfu3
8zs+ya4kzOTqMAcEAhtOn6fhqfzUPE0yAd9iEvIG1I4TInHOSFXulfuLB9Xq8cwLMC7S/k/4X7R1
xlaqIKiLFeB853HLODevioPGL5MdLXnkDXslk+/QWr4WZUP6RkRehsEfyShM6ZcUJBoPyJfoo+cs
Gz8NQFWp8LG7jRLih7llNnE9Wfrd3uIMqSgTa1hpB5Zk7m6OYORfrjVt1tZcUW5ixhQhCjhgr+4s
+Ip1x5/Zens4y4QqBt7DFIEqNBQjo5+B+1dHHjjZMOeo6XtBXD8M2CfdvqT30+uSB1nXZAqESepT
mKXJFWUBqq6aVXg/il+JdFRmhbX6pwvFMMExea8OSOU90PTOPZcwjH3tiMX6cIkPN2EKxM6pRU0X
LmGQCNSmiAdRo7/k0RYF5xbWOmLNQfILbZu52P1tDEX6sk0pZYfEP8ZxsxH1biak10Gipype2isi
bpTAKDU/cAFuVHVlWAKbQbqU6mthNXwSSiDrylhSAXwW5tHLd6FQ6dstpUxI1TY54XGR/9C3vyDP
PcafrIsB+qPQ3uHR3UaXhE9yA/Kzrsv9VmfjNK7BjaUctJaMu8RVYdMiXG1Xql4WGKVcO6SNHI4t
ZzsDJNGIuReQf4mBDVigg6n7qANr6oYenENqO4gNxb1ZW6lU3cQ1Vi0mVCvFWLt7BASknCCqdz1u
1/kgLYpO0TSeXcXpdXM/dqmJH54pDFZ5ZZw6fGtc7FOqoYWLL+h4njGo+poxl9AFwOu7M/QGNOCg
RJaowLJg4herwtllqTY93UdAGRdtIZCMD+ciUi0Q3XBDApe/HhJ6jycqoae95Q8iTMQQ0OlkKp8V
jQcpmLFWu6zJAH/z792fshNVQNFJlnSXp4iYvM+uwN+oN5hA6whEd2Pg73Xwmv7+D28VzcoKkXtM
SfeWtbvCjeDmskk3Kr1Udn3ovw9LhFCKbv6Y2pHyMPra0/vCo9ixXfoxDTN8CwRTbVgQJREwVG8Y
dqc3I5BdZNnbKkYVC5hLyluKX+vgdlHIP98iJxmkeRkBVOhsIJDdq7Taha0GCxuy4xRfoA8LO1gb
kMWRUI3D4OWd4c4xsmYfeUPKr/bes7l3DB5BsPahu2eUSCQQpS9ic2AaABLdldD4suHFFdMToCf+
alxtlxdPiEqIzCiEeOVBEtvltuPAThRJcmu3AkMByQLy+WEQSh19d9EmWq9iqTcJZnbIYSNJzmCk
Rf5qDLpnrBH6n7HpF7AIspCHPVYzIKFQymTgjxImE4d82gW2D+KRVSlrTd/SuIqERDgv2jc0o/xF
5cEc2NPZW/x09/oXs5bmSiWoN2qjxs13h8ZzgorvPLHimohLAJuaLmlk/+5pbMZ5buHOxCcyhh8M
2WeQI6sZ2cc/GoRh8It+bsKNXa8nW8Te02CEEU+7hMdIGfexWYw9nWc2lB48puXHelv7uLc9LplE
txE+ZWsoOIvkXG0wP/j7TdBO5z1MMNNnAzDHb6jb15d1NTC6fhGrzneahShIiFhvXcKgucl7XxaP
ZEoOnVbiVBzjnzs3wtV/4Fzp52CmT8Xdj+A7Ciy40XxGoSPZ0Mno18HMCXSMurp2RpQx8GeGgZNw
/c2EYfT9iJaKJB/a5xaaIGLk2s2NOWXLx6zIs/pzhZiLD+ORB9wCve1GzEmN2QdlvpxpjSyawzQW
hNStXoPdMXbeP3XzjYpns6Mp33GjxGK0BQN1iLx3+hXhBEOZsJ8i5MPg0BfFiowC3KVUzOYSIHER
7GzL7WimIHFThgpJ5/IWTp2D+C7wEysMaMW9d+oBbvE3Pnt+lWTLSHAkT+Nu6ljyaHk8kVBBt3rE
zC5BCcLEV8MLWYXpUmYCg9S7lHSQALE/IIzFhu7iJPCWcdkLX6arkMU75nnvZydHJ5B3y5doh3DR
+4lvPwDcztQxaQ+C6Ft9ZOtseE+s8caHexsX+du51BywD16McuOkoy9uGEnHyDJSHFaGpy4TxN8p
5uUTtPStjWB8u5YnTyfNO7pVatM5m2VQcx7b89Dz0tev1bukqKisdFEoqcu+uRUsaVRdMFo0ygtX
cDVAGFJ4XW0P9HulF6E7IFDQAYL3E5VS295xoQkeCss0JypR/Z5rkxCXl5+cFA2U3w73JkugzbIl
kYuXDTeP01U/evO1Qxmia33I5YukTatxnckm39EB1KeOXDQexZtosNsBOrm1AkAjCAyxtHI2LHBK
nHibqijXKs1xGgSeJ8l5NGh3OfVbw0cOEUG/ELpJqZljaTf/ZgqmWYKEyaWzYB+4bAOKNVobX9Pb
DE/HZh8wb+mujX76jA8Y7eWZBIPosZYSQORGcGm8pDtGos94qbtAAuqva24fFQ0dsg40FUF+XqKt
nVn1p10+yMSAVuSw0rgb39NUPFLsOvXX0ZGv/zHcyf03omSJmGgap7+0ywQHfnsLMPPrtbi2IqQN
pWx+ZWdLqx52BYuExe3UphuMMe3a0DWBBq3vhHUTHGJDy8Lg5YDekh8JE89zC7n/2F0EGh+biIJR
CJJc0ReQDlI3T+Oe42T7O9gZpMTKDGVjRJa9eXAJxr13ohJ39MEXjWztNcVfsvMbKwvUCRSE6gq0
rJ91ZSqlrQRKjW/FrEqmcHHFXQhtNKCWkj0hMRkNVeBgl/vyITuLzvK3GRHJ0GiX4o0E4H7ozx1T
tPTocsxT+WCSOHeY1M+F+gb1+QFdeeipBCeCQDqUFzinaHDhAt0LkulWW8R5sVbqP2iPn9gbs75C
6s2wGCp/WM5fCyPFmK4kiPrPpUd7444ZqiYw5TubqvWf9Q9aNPfO6d7cN2dMUFh2feXEqMhxFndo
QGpBiXJkD/dJV/JgFn+UyBfykHJEXrUR99wws5Q8QljvzfT+2qdHJu0Zxx2c/vKL2DlD6RQ8goav
NuSmjHmmYOsuaLoWI+2bfKJecER09q9BhTfLhtEQ4x30nxbxbL0TH5Pye8JZTn+MG+tDaWK5Q5x8
foPQQsNDBndgaoctfu8iju89HAk7arLwytaWJhsrD266aUMAwtg3jeWd4TA7MdvJtCsShz76wcuj
j0aRNzKnygOwnL4iMn6vo64FhGQTwGmfQKAaiypIsyZspVILoUfKevSH+VUm1XFWp+jEvfLA/kma
XbZHlzJ/GQ+hoCHn546FAc/ZQjpSbIhpLaZ5j1YrMbiPtd5rnoYGciI2ft5kUCKrv95uciIn+hm9
gROVTiuCxsFKquyO8PUWX3mieN7wuVljU9eewdtnbRNSMkAyZ1rd92wYA6Gp0wee/vpFk0xWdgnr
bvKVo9IXkSq3jz8aOUs7+TmAJUIKWXu0BfwqMe5/SzhXnvRzncXhRhANC7R9e/dsX23yfYBGcs/O
CSWkfrijyHh0zmoWFEPKbhNSG7LsWYdPMuO2/z13X4djOlbGDMaYFuSNsrQcc63LbQGhIt9f4rPQ
9tSCNZZyb7MqKlGL8Q+E7bncTRCadTS2rKnqZ8KU4jddlDuUyQhS4YuyLZkS049TWaF3hmu49flt
fPA4VzMiHTtRf84JQMCxKmXAEVp3KB5WzzyG0SYXsLSf9EtTP4kx7P/LpbEhmUeKuxYFVzknujWW
wrj+iamkr0UZBhakJvETHGhZKvl5uTGBbOqC4bRyv0Dk1960Wrj1bWbM4fDM04T/SIKQNMBDhFUv
aYn3lA4DsWgK5fMyw1dGN7kDlW7hB2aS3Wwkelu0ZvVVLKfjdGbjQTVAMVWqojooPMAXbWww6WhL
oMH1bEMec2lnjHm24ppYtIxok/Ljj5LNhd3j9qud3DtSFC7okmTB4AvTVaLWWleMZ9+hhvqVVuyZ
QaoTWQjSJCNKSQ0SaBM3gz3qvY1Ze8py/fOwUFnnews97Wtetow9f7Z/E0IOiVNmsPBSNIZhe69w
p1OpQWmKq1Ilw5nZOcsMYrwuUibEfcNVyzQ23CEE6j4yp42F1qiwhsdjRxJl8uv1+Tg7/pMvF+Dj
k07EJxtEsSML66eZ6rA2YMl8j7f4thEU5ObsiZ9n7ujWwklaFdrrr/LMjDdTwgAJlgpvcy0VcQTh
PGykblaPs81CAsh2j6FjDwF88CkNXNi9Yj8nIMxrdq39mpw/oXIcEOXo0HBl1SuBJAD5zt3LkJdt
A4paHkJMhDZ9hVdBXKpunesO4gHn2yA37w/a9BzLqA5njfk94SMH+tOZbOnT784/hULHrTOgXqGJ
jPg2ys9079VXB8Hl/biGvwuNq50xvn/LmEljeBu5rTDqlAjVtUM0EdR0sW+elEi5jMNbhNkXn3Kp
tb6Kc/CfPTqiTblb2LY1WiXqWz/taGImoklpNbu3LfIkeS08LkCJsKahpPllDC6sEoFCNxnQofbv
HVRHd16RgkS7c7mcO2lgWDSMLV5mS2j7BLmzP4KZbdwB85mzV0SoE92qXxXnrBCD5QER3SnUr9Yt
z1SQoF6dy9y9JniwY+ndmA2KqMp/AsTqfEIszuQ/7HGes0jJHj/J0hK0xa25rzfUU47hoBH8+H2P
e2Npm0JAPxPdxsD76cQEiB6PDxeR1HL7TV8iJ64G/MRWdA30/N6Xa++eXtogmEvVIySo3btkiHfV
vhfOWAOSSUn+awzzmxhvVcX5pASbZL4mLl13KWnjmrS6LG52ImrRWBatF0Xi4Xr4WTiJ4bj0nHYH
Dg0ZJcI6mnHyESPrhTMd0VCIgSfy3slGdamobOPS/3AST4xTlcq2w5N2asKjx/mlX/1S5GhKgkJ+
tMFoclk86YiyV3nE98rdTnFCQUJ8a4rhPNZv+nqY5Qb15IZze6qdGW2Gpz8TIt4S0iuSRJGLL775
N43aloM1pPqOJ8GOlPQX354usphMJsxRzEuWho8/3osM5gjUrV2ta8mnL/nOu/EOR0PikeQQJ+SV
N3tlOgbMfi8YtbDWsuMF5ZIiX+FwVpHRg0fBKMkZvOzxTG/Td4EDOnSNNumnK2KT6db72Lvt0kZh
57hoJrkxEVOc8fIrLv5CYVXQ0qp4CTW3DP62qllv3lrkvcXVqulkKNaCZUoPbC8Ex9VmhvuuAguP
fEj5oD8P4hcfJlMpuq2tLW+/W42vmuRHVIpyjY+irwFH6Jt+t9GIq+mrq19wIpu8jv493oJrWwbg
ni+6y+8PW4Eg+6WlD9Gm50PW200jt9zMLS45YoQSVfy8WoCgvs5V1slcsyui1pFT0HANSDTxiOsm
iNJisi0xxt+0rHt56/SOOpi8OTT52FJOca6vOarBtZdZRA2tBgKCPRu62S3uOiDm8aZNC8R5MNzP
WcqKA/1JqksXo38R2RL//00PfpzIdmbtS7Q3UG26gcV/3Dug28Kjuqo22xhceVX1eP0pyebsD9qx
mLhHrNMm7ZEFp98+dlsow8FVffyLceacl2mo6uLrIOEA+MXollVrz4a9yO5pkylai1RKPrxTOGoe
eav6ZuEMst4Ye5iwP6qGsFwTAbugxmgcGraJQdxm8qpWTCHiUDdiv4nkvVJU9sxupIxkeADiedo4
xPE9/c2FytLMs6azbHseHHRK3vTdDQFA+EMJFRsNKSqryQRxqcgIs0WkHI4kBBL6Wsqclp6g+o4F
xa7+b6UMMUjk7rMruLuVuawy0XBPOF2wgDIzNAg9BHmusK3Qdhj9xSsEb0DyC6IPlIFO3d62PNJ9
2YOmxRDyyd+lY54LuxAXLgniv2D1f2CD7D432iy7jHa4t0LtuLqNVOQ6BDxqUN31DdiwKM8UDYTB
QasKCbwdpnzv+I6YdylWdR3AlECm9WoXNBYbiwnbscqYqf9uBUnqtPdo136jOJfX/rp7yPmjGCkv
xqOhUMwSJJ3WOh0Z+usq98PEuWHS4fS0UudKhD9/6Tf5e8lwPY4X4YKtmdKdgeKaw0V260UkKNRT
PLgz0ZkvKUJVKdNWOINr2JKU6EL/vwaaJ4UJre6ulrjUV49XL0U0EKFUAMdkhcIYDxd1dXu9eYCH
xLmYlnXMp3aXbdchzL7ctw9m1ACIYtfs4fKpT30BUqj9AvVOa3I+zm00gUrjfOPw/wjgicZ3/6uJ
mIx7eK2a0SQhDcSTtHMJJf23Eb+hWOw6e1kyjh2Tvymxuvq4lXiFxp1qfOgQrywSH1FZZmcEy2FG
tr731ceJhxf4iQXw1nBj5cSnZNZvyLFMNIRWSY62lR7orJyIThjn/Uuv8LiUOpGODs73VY+3K/ME
yZ24s06Hos7xu7e+ZDWmL8S3Kl0s4P7K0OUI5VOMG3inDG4DBky4acbmsBhaz1367kplWFCe04dQ
GJyjHQmkzBFAzQ4Pn3QMNI7SobMBaDKKS+SphzMoseqeuJvswSDopGFJkEY/VtZD8ONBW+OFdn8M
mq9LfrjZXPzHTx39w8eNyevFSwnYMMvsl3j/LWA7ZkR6Q3/C093lYaq12Jr7aJDt3gkxYVVJ56lK
pRHkpTMTkQ9pfn+j7TQVuuwluW53W3gXpnV4xKHOU8zBfzlduf55gKRBm5sU/+tl2wsz2R/ET+6b
GHMJ3iEV/aD1L/b/ld22jxsyd/psLwI0lKshca0s+30t/SyGOeApBFxIDIrAdx9WpHOJUsuAc7+U
gDnYLjZIWZYoUPkjN+e/GR+rUyb//xF0ssrlprVaPHtEAbLswLMXIuJl+lcdiI2OgqF1B9UW6woN
mkSlSRTpZ5A+UP4JUevJzt5FDA+5D4GEs37ii1bo6RWvQJ+9ukk6brSBaJmAA2LXv07nkmEkm/Dc
vR+IEnmNyEmIyiPwT6As4bZqzD0iEvVy1k3SIxUi+8d77AqFUDUqN1yrklkQ4WA4yq19IAvsj39F
MhIllFlMSLGH33EwFkUfWepDwGmcv2JUsWAdEUvWPruH4bpJAQsvgxvvbVrv0GBTGyP24ggoNbbF
YYqdRA36gfne3QTEtuNjpTWyteA7hBddZBXviIDHBEU0I3hcVLl2ZVWHYREeUEiP00yOJXoA7WyE
0j+zX/wcH42ZJkikANhJo1kjrn7sqncFlkp8kfGoBg4dyOVllciWj4V4mNGQJnGjYhnwRNfXgjbM
43mZzpMpj9Gg2XOzRhQnWaRzKVg4TWfo/WlSrpdWGejwAhPECJwYuMFZwps7N+xXabzDUw71memr
t9bCwuAAgcptieWtZzeh181SwLz5uiOqJZVufcIbfzsjsOJs5z4TjpjJPYY04g5Jv/+UQ4smjQaJ
vmBHXD8M7d1EQG5kRRGQYUbB3rTDtuMjluIBJq2231bkawMjjc/oHeBtcyBDY7gyvafNHT+uDEWs
dmm30qME5pAwogyhYShSYEffYZ4CAfncP3RdM52qjtZFJ2f8qvtAeLl+qsO2SsQ+OTv2gfn4cRu7
2onyYrSRRw+m5VNGYZi5/naKiNyzHWeiMddKN8On0UFRSNO/MkEkyL8kOxtFRBrjp+500+fw0gRd
fhP5YNIYsttFWgQMwNgbhPOpihBi0ILgxfKiPSeB2u1yXaM5X1FoTFDxEt5Ar9Pv6wllFCC4RT7E
kiS6qlmITyG2C3SNCTy9rsTQTwfyDzFfTjk1+LjEjMfn8k+iaKEeGuCb5eYkAC9f1QnBSUcj6kR+
YhsgF3Ene0iaPA0ZPSyelZ2lAISYa6hTZPOw1NJ3ZaRHT5tcvx3dg/xRTciit1/33FK7W6qTlkFP
mUVIi0Pv15h99J3X/jizkexQUg4CwLFexHa8T1Y3C2Sy6OtosLVPz1tlL1mnhyC3dWEfi4rY0d3r
504+OifJdZEXVL9FLsKWgRvJRgE8zksBxkPI1U6xkreB2gPdgA48ABT6SkdNA49hdgi7y89rDeqD
QGPURE2SzjslNvLfXGIT7lVXuisx6fzons7VhUzdp18mFQvmh5DVbqrOXpJV82/fUr7+QtJs1mIc
nk7leUc+RiMwJTGOy3MYprOMvFslardddXm10JcV/65nUz8edBwmf8wgOB4fz2Lcgfse5L5uuGqy
XrLU84znm09QikEQYcnpQ7YV5H/BzMehPxULsHnYeXDJA9vafiRvx6ZACydW1XPwGSVUwx3W6Ovw
c8e24jAxR5FZrqCO/XCh9B8U5jiNS4aOqoevlNsg20+fpjoa6m9+d/E05swTqjYJxX4YlAH5HT+k
x8lOCoTqTGgBlKbf5wyraR58XflEhBlHD6nInJLAnmTvRNNRNGcyrARCus+wZwfA64R8pZrz+Npc
b1bmT3u6TZ0ac2PfYySl3XSNFxRSX4Pi+AlL6kKiXtt62D8Qk04wHPTvY8ZiZQbva8rHRQCRB2WY
+mjdg+HwqRqCsypQ2OJ9+aAjFdju79F77rxsgIRYzEeIWIGQWO7uy0mC1MDL09yj0FKf4KUnW++n
W9us56IeTs4JigHKt6CQEMVCcd4G7yQb6D8XkPDCDwkFhyFbuDClE3oM26XBaiHwYv2/itnl1xD1
LDM5FqRsZbRVrrDYtTS/gXN5R6OZJSA9qB3cbCjj05yOLeu2hqnozcLS4AcJ6wHScEGULsWzGQFm
m/isXmcpgtPK02e7WEmmCXkj/IYC4tDeHVjTQ5/SH4SysyhcL+MMyzSMrzvGds/Vd7r4gTAz0HIR
7lUfsrQQMV47gDinKpDcXBpXe2ewvLc+yhV+7ZcjhHZC3M2S+BKmaRJBkX99amFW0T9jSHyPeRTF
QnjgzJicEJ0K5MBx0MwSnN0Kg4SZBKXYmpyYPTX/kPijRbxlpOd5Rne111jsP9vymeJcCAkgiKf9
d6oTzdYybWU/o4XV3tJwFF32aXTQXVwdqsn/Pnvbv2xczx58u/FuZS/gTHH3l6VY0xlHrOp2dkhx
Bac82jWjy/lmFKnVda3U2V5N7JaZ5Z3zxBzthIo91aLMqXd5ROCgueooVgpcd/C+Pl6rX6fuS6kN
aXjF+JErtvTq/YHHfRi8FWTlZznzy6rxg3irDCZp+uMrzvmEBKm6uo1odH51UPVczSwLCIdCDpxR
FmKkCJSy76BfE756Mtkv5Z/DbG/yx3FlAjLRzTgphuMC2L4uQ+kEXrt8elB1QNDR6Cwk06usC2Jj
HkngzzaYak8NGX1jwbdXFsO+LE2Wh81MmBsySMF8t6BvnrX1xauZ0Z1ijBxVgEcjZYrQpMkcP4Q0
dvIlUbaGLhxaRlTKU4a+ZlFhbnG/qlmr540E5gG1j9u8LkbwsEx9zXcEqmJvJb9MMQB1emE4Tlfj
kzfna8D3Vc1IUL21ZmQfdddJsXVB2NvtZpHC5kwDOpq5Hdmwdatbi/aCV6XDwJiGB2we24dyuW6O
57nfZ26jLu8J9di9HnnupUTVljo/Vam4Cyw1AU0Z9jhYVLceW5C7a/gA61ogeDP5XHreKZhksgZD
CXFmvOL1gdVJBvg4nnLWLXEbx6r9thQ/deJFl4BN782+tJSXgGxgdBkyWVJIXlGaotHD7TLGNzvM
5WkR+jLnGOPbB87lZFoZaCW3rzjngnzYu60uzD/JiQfntSpdAv3BawjetwMMiZfJ5twmOB3knUEF
CuPS+u47Oe0rb4TbT/YlQ3UcZv8puhYK/2ZYl1q8fZhK3EtN4Tg5c03arlO/pfg5qcDL5N5bS7tx
z3cpZgj33UcdXVZU+xBsT98W6WhM+OFTUINttYZRjfDQXa6g5mCEG3xBmKa3BTyPgKDgfPKhYWul
yL6yMB+JM2ZRt0o2KLQ+CNApG7/YKQJg4wtRLnoCsgrN2bjT8CNxDlS3QOMX+5uioiROjsnZ8v0r
gomA8qT3OhMeXxw8IxjRjsHpAxzwt1J3CN/6k1qC7ocOYFhQ7ZtShdVJSqruGvc9qKvhBsFLtpKd
FzhKpWceCIvatAy2DTbjHMhZO+VM2nTEzBu4w5qL95M92bWhHgXbhP0VDt2n6Wo3Xg+ZSGs9EyET
SeNVDJduhlPI+pKUM/osA9M1eAN3zxYB7tsAJhv5wtYo8QNzHOC4xvxli+3363Wvs+8477SIXWAN
dOKvAu/P68OS6yZhzWBT2pzaGbd051Yf1+o6yltpeM2Cjhzg6Prs1T/qNse7FTcnkU8mhAwNHMYk
arB1CmReYUHbkXrVZGYmQ/dssXkcxqKlMNghwPNdno8i8cTSBCMJp5vkbNoC7cDq2HD+AaNYWLtY
dzAMaZHs4zDeCUOCBVm3Ca2vyzEVnWgRwjB+djka2B2kRBo8PMON2YIMWD5j1c4R4DlbE18DzQ0e
OZ92MOma3kFqDPARlce/RUHUwd/3/mDb9zrNPhmcADAqgBPvTbdCV1hgV5EoPLogaskBt3YUfqyX
8blweLFUPs2ETy+JQllTvfkgpA76LzLgfwc3WojW+mGCNKu1lVFBJ2QXjmzZsHhAU8gF9saTMpkP
fa8J4kWr83XM9oc7LPr8DT78wFHKi7tu/3TqsJxcsLEbH1s1PtERjxIsord4e1piZ0GIE3SFikX9
IBfHm0SGVHcpNPhgOHGeMg6kJZ6KSjfH9whktZJheiRZo8rO6QyHE1y8aXBIRGc/uywJFekKBlj8
ehjuPqaZRY4yPz+mqHRNvI3rGRjrVKKQTxUFno1tVLjaH1J90qqm9JdO/h30mWeQDqUJYVFWTMz1
ebWjDw/I++bXp+z40HkKmq67s4677uTOM1Dyt0QEM2Jc7o/O0+KBHlQ0PB5Mkd6ISGVEZ6VXVDU5
vvmTNWWKQLfnf8HAtUGEns39iddjekSPMT87TzMmA+eBfTyWqSQmUxYz5D/VKOalsNBlDK7+3Nyv
i957ys0em4j49jyVDFHsjobbj7LG/oXGMKe+/Z94CdmRE3oO5tZq3cvuReKX6J3I/mDWfVbJtVUR
XyWpH4xc5fqPXJqez0QKDzNvph2OG+5/LuJiw4DeKr+stfjswWFPVpCp2e9eGhhcveV5xcaRWCMx
ra0JaGLLr6OKC1X8ZRqsTp0f2LoWL/W0duUw1ZxpaR8ruvpEjoH9MbTQuBaf82J8cngA5gbT5k4G
siAHBui/rPpYwHZvGzuWuezIpnjARWto5Vr+8hDWJ+aWc/G6pnDzDIZSN5ARjw7Z0Udby7+NuTpc
xneajUDelITSJGcWWyi/5zefJSiUdoiqqSH8Cbxkxgu5YGBGiOBaUz6i9gtnkVCwVTEsk1goHaR1
pxRNFfgjNgJibryII10l7Qam+x/z3AMMvkX/9St7jm7ecfBEKsVOVo8tP4VWnUZAmZwzI0QBN7k9
EdoJ4Uz8YtJoqKeBaF7Hp5eRFnxMGwjHAk8rgmmXC9EzGDw0VZHSCHfC9z4wjTmmu3Mgfe4Dha+b
KFb3HBVKbeBivOKQnkh+PXPnndz9cZ/4VGUrwCWYBrrbKaqsP7pYKEJdztx0+GROo2q2XQLkHGb0
sgQ09Xm5xNzXJAbXj+9BvdBrQEBOYYqWWCVKCm/3y3VbcA/qMriTAaSjcpqoM9pyX/o2QmOFIuIA
w54Y9k5TCWjaF+tnAckxynRqy3CbJuggtOO7cIv719PzLGW8OP9Qn1Df0qwK4Nv11mOEwz1LSQm1
DHdu0dNz74XY266WWECGSubSrNr07t3vJJ0iADOEaDcGCzZY5M+YOvPybecTXOOqD0iDdJkBAQqH
vjQreTmAHPANdFmecEXpN9kXKWF23Nqn4/rlVaQZtehjTfTq1The33KPHT3bJBjlfiYuSxQL8G+X
8jFIiDHuKJSVYhi0gdxo71iHDtvEE2iYC7pS4SzRZAGCPmfJBWtWZCeaa1X86KrDk47x1wevv50z
H4AoBtHpA56E+0KmbiuuEnVzC6bDiV4GR4JncJ+qbWn7GwrN/oC5KF40z6wQ6jJ24X1CQUiQkgJE
kmpDHfPTi1b8UgDdK5XdQB7CX0TndfdnZUmN74kYNT0jId3UhPK1BDqHEy7OBd+3dPmZtbFLypn+
6hN50XzmsGuP4OUx6Qgjx3vCtltXZjeljspA2RqIFphKQznbCVq+jCfsIduXscksSG602h/3kmf/
6l5AcB70HUE6t5Hi8x/NDEjDr7jDE+zi6HA9qKN9oX97o1a49MYlwmRqM3OjpSPF0m5kJo/h5FZe
bZOp8mFCO6L3sYavHp5OM4ty940vBKZXwxOEz7AMCOVmt6JYDUmqW+Dh00cCY4axmCwS1qph/VRE
knAr9tR/BALpIK4R7KXp1XSDn2bON8J9D1hPiwXJVGDYfapOlgtbY+DWgAxvBSX0tEkw6SsbOzzA
mzQJeK9ZErlAZcBUmO1Tv1F7bk8wxJxa/Djay0UamjPyo0EzlzbFV7D3pk28XzB53LXYskYsRxW4
qM4joGCGtUvXVWSjupBIubM8qCNkCU7O/4+C+o+TWUNoEJsSaG4I6ewppAtgqzc0xxk5e0xweiMp
9YD5lw9SR+hSGCdPno5mc7BShTZ0wR8auHP6E7sa44PZyqzQ4lQVMs2oLiY2/4sIT8P0HVpJTlZN
p7gUw8t3lNqDcq+K9mbX1I//M8csCDRNhBqmlzQOc/osoYTU6xdTy4WnGwKSkfNKydgPdmeNwKl8
8M4T0BWsXQgrYtsklZq14ZwoIReIuF2/Ff81C2Zr01++W9iuHmfCw+vz4BzZSDZPnP6q9p3H1ycD
4QgkY7YtqCK4DfF5uYt2Q+W/nylnLYYvW/ElvSJMsmoSaMt4wjDbr7IcPr7ql/h5xFF5daO8FwwD
AAG9ytpABb+mKcOZtHClNzs6yFBkmWpEqSQzjfvDlZmSxpxJYeiTZV052v7aZ33AhrP8gKwt0a1G
iCtq2v7J6kK9dV5PJWJ1lx0y2Oy9YDW+7Wov5sD7XWRvUGRJtjwG9TnfwFjsPhGjft4hxPPlz3+4
ZTuvFdchFynDOYu5R0KGlsezmtwVBT3PC8REGntcuOjHD1Ug++hvckNi5GHRJ8xIobFY7F4S4uSU
oTc6yxLbizMIoLeQYhtIrsqWbeW5yRinjRySjfaRt0fk2gqc6exH5W2g5RXXVAsBrMpPCQNrxk9N
RrcI7CXyHVnaT0/P1jJiKQBGcDH8yCZZHPjipyRQo7U69Ak0BQYKZofbH/qkanuipBVmebwFSvQ/
dA9nk99Fkks0mgKKpLoPwYKp08pYBLoaAnR0LZOmY67Sqyin500nUCqaRtfYvQ2mD6QLAEp7MWiM
IiwG0Ss/GiQw/rRBGGBDtfEFF2TiUxtjCJpi0sveNGsdpi9NuGa3NRhhORF6XqFEQiCPGvQ3pMiS
kTGglb8xEPz9AioahlAd3ecKcIecaCiB9hBCnSwbVg1wFTk5rTCQhaTS9yq4QrCi1VpPody8Hn1e
JglPlCfHw7E91RYe96jTRnPiqgw0hhUXT98W7yCNQGiKu84fBhLiqNU9CBdNS9UM+AHf0+T2j5Gs
egkqCq+WUlJr1fDPRhUfWpPjF6BJcQ09eU45Z6ZUIcAB8MmZg7J99pWCWcg/TQ79PKk//lbyCORK
O16/9s0PqdKiPnw1dAS731kKDtL7i936R5RZel2H5rtXXG7sGKzUA//PkUVSg02Dg4Vpu/Sp790Y
H43G6EYT3J54YgCjFmRhoEi9A8KHPHVq2CYPxgaG0x5EwnQ0nlD1l8ZBU397h9jVhYUoQintx1AL
CiIRmOKYZdbRZaUNR1esdGzEoWuBEntV1ESOirIEgYCAgsDb024+ZRpUIGRSgPvsjEJm9hVc7VbQ
6xH10/v1dHnqkjcTfBx/uchPaQnakU+Kr4kWumw5LKP1XziCP/tIkTqCp9f86Bd5qJH2wxWclQwX
LtdwfO5+wxM+dyrRPiQ3zOvSDwYUI6v886VXOyazHdN1lzPmN/CbycDXhO6ArDjfPedhMHIm/ZL9
j+MCs22mpwWNdWuyUDO3BUyN9aKFVtSO9kZz4JcJ5aTvkS4KQ4xg6o/ISdvrOXHRQJY+/F28fZ51
z1GRb7Gblm0q/VC+zTu+zN2p8Tk3KD3OiH6n2jrJunRr4CMumbiQU5gcnRz3rmRPp0Iqg/waYiwX
2X06gVcyxjgjzk3MRtkCBR6FudvqeWGxvfBOWPdaG9T8AND0rkl2HvF5HMHFp9UAz2yP5avk2b76
WhpvNhEkm4Dx31eHCezSfOMupAroGUqL6OCuhrG3d7vqlUR18e91aW3uyqic5aw0gCDTjgK0scRG
lJU8dxAUA+kxFB5HbJZpRGwGnmFsBUaaS/FkJxHNIonDEsksbQXzXhLfobIhV+fTRbms+gdWi5mV
FaOJ9UnfvGgbNR/y0Aahlp6IzB40gNILL7CmcbyC/qr0AUhemsW7KyaG/3pMqvQX9JeoYwI3YVM0
y2fNl1RQC+rd24/cyFYVrs9nsXpzUZ2L1pml3ie08lpUauNL/9QuEM3GsBZ8hZSf0BT7JECvd/7U
1Ll1ftaKSU90ebq6D2ibDUDOrrl2JF8tYuvXf6VOuQiRaeM2oOy8iZE1NExi5K/z/a6T8JNq/roO
j88DtNESLVB/byWXeMcu9+unrVUmay4O8A/9R2NSOMili3mP6Gx2StDGp4ffJZ++YGkoZf7cVkIa
9IunYCi0mholoUbZMIaKRnjNQs2B3xCiQbkVYmrbiTha7CF/5Tush8ArxWOTCOOMVFgbc+J9G/mZ
0+VVuu+ehNFVMy72qWAiCHWQJehbFUNVGTtIZfuQE/9RFyzzRHATW1txgWuaT5d9m4TPw/8l5PuJ
EQGGNUmJbIf+owWBy+YA4m6r4nDBpf5ksu5Wge0FXJZqkRHO6CpaQMox3rTRpggp9qXCH/eRDBOW
GHakpqgMtX7h9yTKEEw9pvO8Tg8/Kzy71WVASTNtxouK3P8Uyy4R6csgIsqJOmL4cepmtzkyvSaw
yeVlFIpdMAd6j+QNpTnkIVL+L9214eCvQbn2trN+V9F0YiGRG6+cYO4rYGM0DF8EJ4XLLF+rGHSi
3pJd4HTdXEmZTKOkYG40CJ1u97EexQO3ceX2Du7O5vyunGrbGEEmWF4CNPQSkocA4sGwxWTHOQXr
uI9RkxDrKf6dMHxADPGjUkSJJixABREr6Hot+3WiCzv2tAzGIPqbM9MIHYqZEbw4FT+09NaRebC2
t7/rkX9mxpXyHnYgvBbo6GRnTPQ+hCdYY66VMrFKmKaT5gLDbJcYv2Lzvl9IVIXeS00inntUiB7L
rJQkKsJoc8TBfxwWmKLMPINzCuLfNLURLVie58cmx+B6LmZVqwj5S8r670q6x6VU2yKTiPIXkNoO
jE6ow2s8egI71ZZRXiGfjRfAo1Jr0CMVpse/8W+iQGOnKTtRbeZJTpcIYtsAKLDdU3Q9vnX+z8mG
rgzSKRLosij7urv/nIP0MTfqSrqxCpjhSNbW5dDqrP2xxZ8HbdzUgKquvQOImitUx9ReJaMQTWw3
J/H+lKvTXXs7IHKC6cW5S5fZCpHpEUZC+DQQF0U+FuLdwOF0l/4RnkwO+cKGJ2xqUZQv/QKcsPxI
IYT6phpwSuBpl7InY9uizXagWZhZpv37mg+2FF2yvKH2GfXALVojTpT6XFR65nyAeTterdrvgRqu
TdnytcCgDB9oaIVyeE5yMp/t0F6Ov3eRBlRCYd32JDHmnZeuTvveoq2PlkRcpmySw8kMmJGj90kr
3oMs7yedFbdFIpbeHcl5aj7G8KJi66q2uZbplyh0QH2upGrt2FZhAqrq0M3lY9c8NQRfwLv+0Okj
buofRPoZ9PYZrpeaDJxZcJbKFBkwKYiScYE+mrhX7bGxLLwE6QhJeDiVrfKRV+PaRYC8tw+c0dxq
cMamkDhzCObGn5BtSrg67maxF+Fe5FaorrIc7kIwVhTmYdyeP2LIivIaltfXlZ4g4oDndmAsH8ji
+A9UVpXAYLpsaqG/V+c989Hwgv0S5TqoSc71gNvn7TgC8u70cTMYlfBv/r+pSv5l9f6zPX/1W1NS
Y40oJtS9WpFg/9DVBBMitbYD5Jyg6tlqOeQ4g6BChDYvbU5nd1pmuMSVXZDgDxBEEQSAwmO+AqVU
3Xar2UNqZnig5ifPE/6w7+SOqfh7NZepgKYt5sOlKmo7T2BM2XlgMKUXICGANRDq91VVXR2uvOod
ib9soM5FjXWgN0qzRD6bk6/8CGQf7/AG32kkUbyx+FSDtuOu5X3z9m4jEh3JIk8rSKo9naiGem9W
CUqEGUyOgdcBnPH0Ukdq/fWK8PoPhWAUZ3cLCh+tgOin977nBOCble6ZMQKHXtaqaRi+BPWDMbve
HD0u/Dtx3gRW/CnsbSSNzQ3ARLGpI5TbVkbuEw4N3f72l5/XKGe8HJdvWFZwtMDXX8IU5elUDBXa
Vq0PURC0h+GzQIaPZfxvb2L1i7d08Ui/eo8bZbLMgtSnwO/1vrG99eH4xlLvGnzsm7YKJ6tLIb1Q
WLYvRPs1WkmUyoiIN4dBn3iK0wnhIBTNDb3lAozV6F3pA8Q+coTsKGGT8K7NKdkLuWxran8aRAO5
ZUNCg5XT68h5fetkbAZqtKmMELZfK9Ody9KIaifM6zOc8+3jRn/ki4WCbw8XuL4F7xURg2R9tXmk
sbXpB6HpSByM31NWOj6eqBt6wJP4oMvTNiICLbp6KEiQOvCv3r/ObBIoOfBXDGNPGh4Mc4KYKE/I
wWcgxiDcuAMr3cINjokiQIGpbh48bzAcidZRDCkn9xSVc0fJGciCcJvueOcygIGtptD8dnZtUGCn
2YdTJ+a3ygfJl63VSTkOBCpJnTTT6wKUIFrTyHKwS3BAzrJWGtWm5koP3XzqVwSqzcvK9nt6yX8J
k0V25wnQd9ylE9qIwdARZNQmw14U4UHuzIC9IRxUyEJSVessaporFdl3u2zpiqL5oTiLqgLOvyON
8638DLWsvI2jzg1LVlpNKEro65QlE+/QdY7L+FqiavrEDPIJldjTVYFwvfgi5jJ24Bxtx66VhrK8
BH4NWvDXC5lQ3EQmkyOmK60Ahp2NE8I687ZUfk+SNTwpceH5A5CWNEaHV4LW5fgGFzxQEctOKU2p
udEuJT+ZG+dmAfiBjLGNSu48XGNp27YvLSQK/VDGRANCxl7b5e/KWO95uan6OjTpYVV4Zefe/W46
yTta697LYxyNn0izf31sclLJlIVlcYSo2HelxSZMUkXBzhlREaajN4LxjYDUmJvpSvAnTeK/KArw
kR+ymFSdIgWG0S0tALu2FCTD7eUX3Ukht4T6JZwZgZW1dk7a7Nml5FsY4p7Yg25xxVm7ed5uCCup
t713u7uQ/wfC7yxk6fILoTUhdOU12KGPM0A/gLwGHfh98d+zdFt6njbBr2vnE4/FvIjgiQnwrx/5
h4X2SczNKGn9kahQjH9Q6X7rd7OuJ5d78UX5QZl9mvENK+Oqdr7tx1FuvW1j3IftlLqNM0eMncDj
ZsfQs2Kwc5nKOwgerXGZpa6w2/8RLYuHLMh+jGlaLBm/ktzogjL1UsGD2FCvWsrHJIm0rtDflsYq
R0igVH2eia1vwCZmgAHCvI/hVyYKBrpt2T2ySOHu/qaq9y58ktrIQ4sDsmX2ly/wl5aOc8Em/+P1
0P2B9KUUX3rpJMmzBnV51DY8cdolzdkSx/YJSqo3zxPKhCwj3n6EVI/S38ieUz8lg3hw9TmYVUkY
FWoaxh5vy+F7NL/+TGfX3sRMHL7LNZJZ/0WInNwzagqYKFqTBecGYrDectRnP2Qzawk1OwNKSXj7
A1k0uzS2f1cpYIOMKyv7x6sUu9imq27kDuhKc9TPODDTGduunHQ5lgXu/+wgIuGbLuaE1/XUtlsI
ICnklcI9YLORCf5cqaJQnxx0/J0Kh4DhjDHvaluZwlPNZkCejhN8ZXnfPaxciobRB+nO3TFM5H7s
150qThc4TfxDUyXjqmHa4tpwSQAljFC3mAWpFzkGQAGk1kcbb3BJ3MMuMbc3OuNO9CitZonz3MPc
zCx92Yb9/61p4VtRSYRuLbM0Io6ut8iNaagIxZUsmnOlkz2PnByqb8zpFCD1pKP679+2daQh6WtO
GAVpFvSLyeQnsFX6NG+VfMcwE3Wsj/MX5IPekU5moSTDhUoILpPaPyq5KQLC6/7eZkzY+VnaLlGZ
PnGy5CVPPaAZXYiRe1eDxr7z3ecpb7HmEuuQTZiWxhrK5oNhTwqXiv7QXcN4obBi/Y0lhQu5Oelw
67tkPRh//ePzaDhuZJmFRofJgNvdzk9eb37X8jJRS2MR5uVUl24Puox3XdW5w8Mj9GDSMLSOVXEw
4EiFbxsx1oGwUC9yIdIUCVq1C+mHhS3vWs6lBe0bcmM1nAWqkt+qUACZzjxBlYuqTu9+9yzyfb3g
TbW5/n8BuMDZq/v6OItCx/7osYFVlFNLI5waZGauhrq1GfVRSQlQ5P+Tq0X3bBVvdYfy82e3+Ebk
g/zmKKWk958laiEpM2CfwxcZ4+JOI/KGgxgHwy0aXuHFEPre+ld8Uc7mDBHxa+ByCj45a0AYsfHz
dM6cX3L6QLrGgUBQpOXkJpq7sxE1xZU4sv3/XpGcXyvhd+AZuw7loaCZC3wJa0PUeAbfCWxBge00
HokjGaoxxWkXp57GOscKBxvPVqWcAfRq/VHhpngaPquEudxZtbZwId8xEfut8mAoRKKxwOKRIj/H
RPpyjMLhAnBFZ36KGGMPlZRvKZegO0qa5nWBlahTiA5HEEwaYOs2uO788EQNBEs86RqfFvpOw8UC
riLtXeV4X7rxVc32ZPdtNzodcxUo48JPEP22+ZPcL6w4k629ZWyHGKeFjvwIFuQgTl7cXIAM/G/j
fSoElBVKdG7Wo3HyVAMUGWpSISdzDqwIwvi06IV+17OhvB/euvDfhGFQ7wSlWyln4FLGfeOouuJ2
NNgnwpkFdESA7LMdZlVInxV0KQK0bVxuG4XFTRvkdy4EGc/putzGai7HhO7yvlZQQXN08Nt1rgIv
1qQrGMzFDksD+7pFEtHwJJbfteHCIm/jKIY0vGhYquMNGOf5b3c13cLKH5//M4YWlNCFpviialOz
rDvDAWnSNdaqyoaA4M6f6z4Pz6nAC3NzeTLRRipxoVKfsmfgAeTWWAjn9hE3DgV+0DLVOc5PXwqA
uTXUf4S3fnBErjUzJrn7jJ1kSPXlgpSwQ9xfV7lQewmADJ9hQ7HU4jG4RLqSoXJuiY+IkMXEkkBK
BfwA5w5did4KeukWOZ75KZYbKDgZ9JzLyo9NZ+hzVhLTrmlm8NI386QNTJ/FKSaROlhEX75ti2hb
qHlzZPNZ0E4yEBZWguA2QpvDWhjdMYfE7PIUsGmIkyhoNbdu4+MjAHShDWICqlPwQHJ6GyynIizX
dR4UU2RgFh4FQQ+gc9UfDjfIQaSO0Hb/+RGtOwt/ci2q9EdM8ajNpCUlU5lR9CEsfFAAkx1K8hbL
JRssDEKTRxG1+9INsLNdj8VkphLit3MuID2JPRT4NLIY+k0bZOZKqywT9DObA3GfXMASvXTVq0bW
1GIBUd52aE9yW0l5Ihyd8yGJf2Zo27Nu+H8wPeMP0Qgfe9ZwdFjYr9Jo6Q+Gj6X9Un9i2LZgYTCu
5dLvd6ffuAdmZ1W80Wq2azvi2T9tMpVmP6e9TxlPpjXWU64nw4u/n9hpBhReC34c/fcwMws94vz/
cyVXbQnCdn3ZRUWUOqDgwmX+NFI5+UMytcY0k1NxtUBHxMbOyg7iTFcLUPEiG5EARABKqd/77kr+
Bb1nIAGTnewx1CNLuR+fNQ+vAy/LaVCffJsKG+OPZZjKbqY1I4Go8oH1r/Eh1gdM5orBYNJyb6LL
SIiWfhf029hBlBXPqPSAbWFnIaevK0ZS9CP+qKJPl//j3UAigEyyUFTrkDGfFoA8j/3ADMVzlJTm
N6voSo4vw3bk/3vq6EORW9ZGtvmCSILJvMbosjTZ0Dtj5hPxsbQCxPPRQrLzg/YeatgGxI+0wrcZ
5onI/CRIm/84/EDJ4YGqhjwrmX2tnBlNhT81YcvC/ArrQqDtPxQsku4kttpqCkTWDVta5usodE1I
HbqjV73PEbls8wJlC5dRongma9LYMXy/+BbkbNdwNCwgO93ynkYIGMDVzLUJUExH/NF+dv9fcPAf
Av4+eqLZV4TnATjy7iaE97IexQwCxzglyRoOhVAuYMl0rGgutVcalhtLicj3JeQFopERndUi4YYT
e982ofK1BWJJgsiUKcmgfpE/1zqNVVzyZiefGl9hzWXm2oHnmQPx7vxOT+0zCPLBJGa7ZjYxdvnF
4F06xBgixWLDG9c2C1xEaab4Pbbe0coQzW/PADGUkbI9x4Eszlpj7qW/iQ05mFJe/RK+YBRKqulC
WuwgvlFiuPc/f18/3oUL5u8UFQ9IoQDg1FiaTDNUVlXGjQBg1sMT1hDnxa8w6radguuJAdbMQcSP
e2WBT+u3Kp7epRVG7vN/ODIbCB/06w+fVLphVupQw4wXIGtwYfJdJ5tMTD3EEoeg3SQWQCWdDqwN
B3mTA3+KF6qE48EACoKmRF+uuIXK4FZY8Rl2C4bcCoxeNQMi/BGRYYeZIYuehwSMeos/GbLF+F6t
cSYkp4PmIjPXDCo34PRmMkPiwp3dfa3o/sUHlmvYbs8tj4TZzhPNE/8CSVawy+yQPyJF1aKzK9M6
mqtt6caaVl1WoTMTIHX2pxmsZ3jHsrDo4JOhNWK7zRDCu0TUhHF4xOR738jvw3xv5uRttzlOS5uM
39yYYQFeNRVkAGlP16c4dYuPjFYrsL8EXNxtuRjxcyzf2ezp8PA0OqNbvn8zPZa4jSyRB/P4OVXr
JUnqSnC0IJnQeL0VdGh1FTpdFq5W6VNa60ncZh6oGg8DX8SL4n0eJ8JXyjKAish0cK7HdRF0toMT
W2CbSplcEMqsgTUGNt7pTFOWQIGULtiaPtflZnMu2bQFUfFA9Bjs0SiodJLHTRxhSLfJlvsrQmPW
x8SE/FuM8kccQ/1KZzTPmhjqT9HYBp87K1jHbM3HQRTd54p8KGxRczBpzpjf2WbliiZkbbCOdcID
jleJRP0NoKuu91lbBhFUqSVDu6+vp9uK/RwgJtPw3fj7+TlI2CMUaQV5jDSlLtP5ZcGdFwUbZHhv
eGsqynopY8VXJfUKtAx8xz3fUxriK73OGaERqR7n9rjg4hV2FWsv3mFmeKCucE9MGxeWwIoxxGpg
sPUQRc0sHvdfBW/ynTXYVr6TijCrGw2/X0NoxQio+V3+GCKVXVlqjMV0gicCr0Ufv42nlBOKdcC1
NTbG0aJpUA6LPoX/yC9HW9oWwWo4Z0crHRvVUU5uLs8sxMNsHKsFYZhR8BS4Lz+j1ZUAAwXuF4yt
6Q19UCZBl8d2XTe0evesedGdW2hJtG8bGi3amJ0Di0uPa1P91nV5fmmQWFrGqcJvh24Aqk4/TU58
CwvIluuOu3Q2MZVD6sHRjZ9t89DMZpL5Z4MOx0nZpqRCcaZ9NaKA+s3vSqkwBkpsrnoq2ulgetJT
yxkcTg6NJrLum5V6quIWi9l68WNCPkA/zPRuaOnZMKy1rOSdYmXoOuMrhHerZqtPerHSB2dEFZM1
+CjrGGvIVxhGULYobPNAAmvvYtt26K8WvS1fhJcmHGhoB3gGOs4xAHE51xxipxqQXixhYrCU1Tcy
uiBCd3AYdWadJYlq1gW6DK7q/t4iiGvQkgE0ICsoTdTV+OxaxOm3wagDL6431D0Gtm69RiiltTjq
CC8Bk5RkG+0x3eMA3H9TDkAHwdAlv8E9em09e7lEv77CGK2WCHFOwVP5IDf5mnvRJirJS65SdBc9
SOfYyc6jOQcy7ANn2ZopNfB/rcF+JaOTZo38SUUJvCUtLJQvwlicLYodoRVSgttV0KkajQh1mKuU
Wk1F4C5+1ONeOJUwcJguHdEzNqaAnFPDT/c8iNRux8RevYAhzvI5NEiuNMpZX3GrEtIFDiHUaV+0
tfmq+mgujwRDSnwe+txknGXe8RRGhybK1/+GwnD8fLi48+ogQdJeVWErWyfQ8U3t6ceGoHF4+6m+
+kWUAAhPmoBxdYLcHMShy/9yX6hBUBK4tyGmYIxGSiCByT/uJzQWZ/VQn+lnJPB3Huny8eHVTbvU
DRXyuu1ll+i7/EfoWR4vrSt9syhm59L2VykKrpwLUc46mG/yYLm8I/Ze4PcQM3zq4DEgJxzFEmqe
+LldjtrWznCHiu5+Y4P8flBpLCPtL2QXnSowQ/CKkvwvUdmKKi+W3XaHQTsZvQJo0ZI2tUSbKlxL
OsSzeYH7XZIDwQgaD2NOLESsLkTw6hMV68v01FIeWugRybHX5WYSbYrfI3DqxRlfXu+BY4Q5ZZL+
ddnwYXDi7bub4OXIdYYTPcEBy0NGSpsNofSPj8F8diGw4/GZB59859WYUmyeQz68lNg9A64t46Ca
l8uAXZgqZ1a580UxEbx7obeH5BSv3cXF6gDuFBaoUc+7qiO2NVIiPgtQ/LFsbZhlU0cIG7HFYWzp
yqV7QDqppnWcugRstS7+YvNrn/JQITJuzfqdc6D0BqmB/lmX8MbZDDJFNaca40YnhBg5swmH9X2X
dbr/frnyxjTpWif5tj1846suJYITM+9m79tgt8v7nFtk+kU1tsz8MdYmf5ILTjXHL5HzWHBFJ0l2
XemBvwV6gtN2/6l5zlS/tsiC4DMYHjFybwXpqqnNy8+nMrdvvAnaLUR1TyuRRXNIsphc8Rwrlte/
KGfCH9Nfu39y6QzelOI7I5XVd+p1IjUSRNBBs5IFykLU07FD3uRU4b6E4ltIcx9H39fvxbp/3Xfv
C+2Dv4dPy/8YKFGZ/NNr66VS/OEHhEl+ZzAqVfUKfIUi19/ZJJ/Xi98u8TczASp6JRM4algO8XYl
85GyU6eSwWsQxTM25bFdrz60WAmwXCO8CmRviLA12JWoITJ/3D6JHu4hS/0Ng28X98fmw5MCc0kW
MU8zQsQQ7xg9B0ER26X0rPLhHv1RqzxjqkJJz0anZY204bTDuhyn74DvMgL4FJnVtaTLxxwdztRR
8AG1jiZvX/BPIVVGhdbRiGsfAeVbZMWjWHCV2VEj23zZYoztXSD2I6SM7oTItYsjGcyj0dv2poKp
HESbkQrClikq0TVNJ9S0udufjJaGWggv4mxRSymF7aUFWTaddeUusZc9fgUMxolmKA8z1kLeNOTa
i2RyFwlRsyXOHXu/JD+Q7IEKy5CaM44DvXAz9YYGOToD/f5jLuwfR7hbWav05VehTtnxUa3PXuq3
gHwT1BO/zbndXoz8dpM9Le1nmbTtJQinAPhJM+GcGLJU2Iny8jLm02xLw615XmL1cLCS9nmgFr1v
6agQQEdWmb/gs3HnJudYnriwajuKRiLScVq5IuQwEc0W1s26Ly122RhDcaqj4opuRhNlnC36VE4a
Ffsf1/dG6AQ0XsSU5SnZWlaSyagz2nBVEEH0PSZxVNovH6Ox/k22tycZwRDtW5iNcoFtGgmL0lgG
3qE1XnFVS74uqYUg/rVkUCCT3iti4E5eOripSF3Kx7+xJnZ9PsLCWlpG07mBYlpn8CwyI4HKBHOS
4EcFzLF5u0whmoIpCLjZI/Xu+mvWWqWCRyvQLPzhichFM0/Q5NWHirKHTXmaalMlBDvNJjIo3oT7
CQq+g44SC5EwEqrzOJzijq/UYgTob7V8v8AOh2PGQmu3rRc3WxuNak48h1WU3SxGy+u+WXxziZSJ
rgHTHqI/HaN6nl1UR0O1l4/fZK9PrqLueiqxklNU+iC6K+gSEIAOXIVBsPUaTUWNayCOw/ORLppd
FL0T5O90cXmXKaJkzV4ZjljSlHIc7bdFydISrUPMWa1sxtNKIfjBN4sqgAJSwDjst8uP5o4dwYWg
edfwL4aRNVmj+J27VAq4kAAStga0C4n46GN0u8hMHf58e82n8L6tVTZSAonqzLZVENkmMxpH1Q3R
ooHJWwoXWPk4rWHV/ojMTHoZN4k9HwnUqVS2tWzKG/SYFpcIJc29xRDk5DGFaiT6XWZMr7f5Agbz
jTO6Ojf/vWt8X+FAr3PXtAFY0at8AXf2UGTnGHD6lTt6oZJUS6au2rsUcZKf48eenhktl6I1Uyhb
mcYF/JxgdUBLIdk48U3NBhI6fMY3b2Bp4FcrEvZFzwKf4ajVEqWaj8oi8UeO0Vy1UgVvEgpnRA70
P304bRkX2gcJHNRZALnX6fIzVVc8X1TM+w8DM9DK9409kvXujTr7tEtwBFEyhNT79Dq7/JdqRtiF
0jpeYkTtU3GWioo9Fd5nGQDzM5jOVHjlNJ71COlmpnjNJSKW2ie3XnsnEnhFubw7B+KPeQElyU30
S0FkMnbckraniTMh0eeVCwSM9+/zVe9E+gwyoWDcssEfk/QIN0LDgxm77fEStd/BMA/hi+2de8QG
i/P8+SuKnGQMKXoSTM+cjbYaAVdMeRY6B5xBFTT9rYJo5E+w5LrfWCzC8+jDhYr+50GfzvlSQck9
Jf3ik3wrNVKC//USzpkUUu4ALA6+M0f0Y6lDbVFUcz9E1Ik0p1aUCkHUlCcUwC4CY1zVfHZ74Q08
2eMRdSTgNTILN/K7g7PDfp/XIPLukLHFI4HXeoM682piJKKLLZgozyk+orDyiC3K/TrDnSOxwu0x
qoWFS7f1Rohz1te5ZBAw/o1Sm7Qf2o/BfVZ0qqJ4T8yGpL+NIi7ZPPkMQDvLK6c2yUYgHiWsEMZL
V0E3Z1rjbcZiWqYnNoy+mTBg90PnPcWkTeh89nrPIFwTBRr0BOnPzGNB22kdlggXPvmkh/H1OBbI
KZ6wiHIL4lTjDrPxZGzNdG7gfxXqgTDaywT/cLsFKoISnzoy04SQgyUPRdZzG59yzaEw8ZknfWVf
6HtOiELZeP6Tv4yWxgzv1l/UMxGGo3LevczNoVO8gbOU2N/fui+xUVmE7J/c5v2Z9ZXER3o00op7
Qro6ZqlpSQg6GIm4TwzB7Pw7T8w+sBzM6pFPAvV7O7ys64DnhaCu4aTodFF9k6LsylJhOhGmYe9H
ft+lAOxhNEd2yNvsG5J4X7YFPc2tgUDAcsKf9PNsmw5obcbxB6XRIryFX5rbTJ8NIMzxdsGQrmpl
7cxv5zVx3sWaf5VzzIyJrEG1h6aYDG2B1tKS1QshZ02MJJNuIqsmQ15ABhtw9abM/x/CzI+HaGRg
IS+coXtONlHHP8sc8W2DO17wiiJGG7JxpDQUKWOqFVkHpvykceR1F1aciQ05wne1PUkz++uHXX2r
/Ht+LV+HHtWUMcPkHy3uv1dlU7rd0Lc6CRxxpr13IVUnJRUSNo46eYqI8X3DsER8IuaT06bZmk3u
JULhwwXWTBhEu6pJM+EmoB1r6twxMvWn8a509xKoVQkV1vktzL3t5p95MR/IsT+ZNNt1eq5wlW1b
zP3NoWIYbkvw5EaQYvrHVDqeLxSZ/IQbTUgs+r62ESvnvRJmd6113MR3jMsWDGCYkecngZWD4vDQ
xYpsIwkfUbcbNddE7NQZ+z/GHaAtkaxJCktjVj54grBChUpPct81BnIMB5ro8TVuMgp60mLbzWAk
YtKhcxofLY8ITG/Ky+cClO41wmKrrND/8iOW6EYuopBCiOXJiJ9mKJAn38U0ZYkncAHUEg8katqI
wqUzTFgvCwyZWA23naaLLHRTGvxqXAxSdNL82hF/aHV39xq3OUC/Tg3dZPV67uXbJvUM3NFjljiI
FYBVoc0ZVYneX1ycHxekY40xvxbGmi/tjL8YmMug0aqIFmX+9spg/t9D2Gwd4F6lOSihz/kTDWt2
54K1Yh3VeSXY+mZpGrXNDbCYE6SWrxclkwY/LtPEcI0lLrBzhnNAc9LhHKVDTMKMRvbMbdxNGfsM
d1KECDNkvacrIrqvjzPX6Y6we+lPHsPeZ/b9MALDhaZvlYPl1HCs4kC1xY0+mFibUAgBVEA0tpfE
dYzp21vAKDoXCkSknHbhzt7BQcTFurNTIodIl+zNIGqS8AMGBQZl0hDpD5mfs527/FG9UD4Wsk52
UQwrAV9nGe0V2WUQiQPnpOFLQvmybTyNSuCh6AplOWBC/IQmDi/Y8XXVjJmTMklOufiYve1MGMlo
DdCtvYp4R0bQSMaa2VovkgDngDbgIOlYN4w0vGKvcFtXBy4A9bfiEwccCjsg06Dc7jp12jZkKwSe
p+WoYqma3CD+g7hqaqDyQM85mt8GRIi5FxHVJRvrAtb2Qnz6m+hF66Pm61UEfY1T+lT3UA8vWlLB
1pY2k+Uj0lZuz0ZlR3R/PCaxrChRDOo/ObwJvodCxaC+0blGL/q315GKxaxmuBi0NjSTVUAMigjZ
LdGg3SKnrp3Nz4elC7Hfg8P9/rJFmjwAKHvuRWjU6khnigEq6nUk1PWhRlwuJdiy/zoTUsiYp81l
zon+L26+8W3XEXwMHrvycETP56KWfkvstXF5EI4h6R0VDAVVoZuiQJnLWageWYuvFEiT/g8zukK6
POBmeKTeb75By8sPwkck2TFzrkNyDV752NDeu2sLVxviOgJiZ63f5HsI8LOC7nYEWt4SLmwlL5Qp
1cPtVXuJf6BHgpCuqIcj6gJmDhEve5bdvjK+jKCF7cEOH0b/dAmyfHhZ8k+JeB74yhHr16IloLG5
4VH/sWrSCH/RWJzO8FWJ8VQ0zUGIWC8UbGRZqZ2haiHWWFiw9tMUBAuT7ZfEWgZp6DzPiNieKYEt
o0vrNtWgTbdcsZwaVcU9w48BMx6auqHbrmQWzlsjUm6AfB6miKzi7IE5UYr6gE5b/K//WipOolki
Ycqq5hgc87YKBuSmgzAnDpX89ogoml5gVa/dpSe0hzMymKwV2HzleN7wWPEbMm3X81+UOfeS56k+
ou0fTymFZIQIsUXzvBo4v5IYmWP1KkMZkERBhiv+1byeE2qsRNPHQbDaw8sl/4/f6w9Wjji+oRAC
y/vk2X/7f/F38FCzpsSXJJYMpoF+vrQIr+1iOFrQYKPuwPsOYr2P2kPngbJSRJ+mmx2uIsjKi4t1
cMsvlbu+KsljQeR3kQrtmcNOmTceK1M6KxOfLis1hf2S4TKTQi1Ch0Z0Or65uSSfglqExZbCbeeU
S+Gb0TULA4y18i+TlFG0exFMhTVQi6tcFYa9JRgdXBBPQvxFEviUek+MD6hlmaB280I+lg6S9NeN
aMfKvU3WK8l2DT9P3fuLUlpqDnlAlv3I5R4sqvkHF+2wrMH6Z71+egdXLJY+l2OUjnbYqq4vIDdV
El89oWTh+zg9aXoxJZKca3iR/fgi/ZNuLgafRBDiIb4kIMK7+qo2DPJJKzbOJL+l+QHwURHP3PPH
4YH9YXd0ycg9VfEQ3flB12MC4MYaCL47OHpdJTOIofQa7MrCLqZg8+noeRDEBvLx1iBSEPTyUbQQ
/x571eqRrFqIJKEDu2YOGkzwsb2A2BemSfen5MwRu/AC4bKmJrD6e+CYueOrFmYAkhY1iFtGKtAf
e4NfIPJz2VZEVANvyHim992v6oG26LgEq43HL1bqEC0paV4T19RJgwAnxHU6cSUBUHcPWEYdvjcw
ZZGB7WNQiUdfJQIYGuoB8Shq/EVu25niR4MuMsM0CszfGJj1ZKG8+APa1NahsJLGW8Qwq3olrTjk
vtu6B4ySbylBU5K/9cxeZu7/wMdC/+/T0NBwnCYfmPfWJfZf2wWvjRbibk4wc+BjSPA0j5gWkEMn
SxLgHHdWQhNTW9VCSij/RhzN8gv0PXm1ueysVyiTxBP4ThnJBc74EfyvxN2r37DzaGSQOoTpX2Jv
l/jpbKLQaIoDUX1LHg/taTETtZ/kJlpQ4Bjypj7/g42gowdJPjTaaqF1nQvOOY0pI1TkPoqXpS/J
PSWPABjODqiVm4QusvtKRwMKsXhopQbo3AkMq10MIFJNBb3+r74regeyzhhs9ghdMdP1hKP/YrmE
Rs2QQT1Qm3MHgROhm8LfTS3bG9gh2maMLjLi9DjnOhRDxfvAaQ58k+JAE5O2tnwSUVnoIpcvEOom
Lms58yD2Jiacq7f9cVbdtr/vwt/2q41MwmFBLgT8nJc0SHBz+14tE5ujkUts7fONKBeKvhTWXyCk
NgjZ2bvMV3LQISuMdc3mRfTD1eorUKwoTQsfm2IS9KOARBG/Fhx0am1q/8GxyCfZKS8U8uouIu3x
I9juLepeOllnbJUaOPxQQhKxoiZKyAdINTun1GJ1X00ri673iXT3gQEV+Ylwe4hh4E7ygo7U2dcB
Ar+65sHGJB7MfVuHDW62KzDbqWGO1wRJB+ETIh3NS38QE+WScw8L3Ck0X6eLQq45LkMtgbJJ7VTK
4FGqtS2iJYydbvaUgDifJIwYNEvW1yBGfqlxzwo4rDpnNi6/D47uEzhFhTOE9g1PC6F2yZAbCNAT
8d4inxSrxrC7oOijvi/MXGMOltW0p5EP2Xk2im3ekYH0mjavJhn0JJH6kKAnzfm94+Ht+uBCFcPX
1Ew7jrAf/tOIxVdw6bZUFBhE/QQ/qCc1p4yKtj4LfkWZacrKqGPCYm1KdNj1nLN5M7ZxJkfRJyQ/
WXcChdftYCRTKWD3eV/Y5Qf31hL0khFYiKBQgI3oWlKO+WPZtXMPJKtGGYoaVPab4iLDA9+6W62t
qk9Qdc1lulnKgYBe4gldIhedz3dFd0UDIwBj2LPzzIGgwKeeLPndS/Nlv+vKMow+0gpIozCw55us
ZUVdObY1qRNl1TtQnXbFP9P9cgSqShZqBqEMbPytb35yimwX6vhPLUPRHnKn+q5+voJpANxTAYKc
nxE+X/JZV8sLeGYaHBOU2bYkagkvOMZUihQnZdP99kUpr8u3DsFcAoaqfSEzbOqfpEFGWfQfzesc
lgYzB48Plp9rMkY0eZvMsR63gv1ysD5rUE/6kdlusFo7QoIdmbEikjg5Z0bwIDCustVLIzncy5As
DMVexYAx/Ps/RaJnSCzWJUsSJwuH4IVokgZ+r1Aj+ewU1d7h4OPWF8yYUXicsaQZ53L1lHqNDOzO
Dar7CigeiXscFGKlEOiStLGvoDw9yoUc3R6mcl1ugbkcn4ElgG55g218vI/e6BE4Yw0UL5PlxXsv
OWuf7isRhnt8m4MxBm0jT8APNEhldI6zLjhHPBMtWdZz1967XlJCb9WOEJqYdbLyCaJumNAiJQby
cf3iDLquTagD1GtkU4TqJfPS1mZdY7poR4ip1t6PbQ/1j9a9wpqBYeQfm/axYAd/X4VMVmIlixdJ
nciuK8J1yYeqDJt0zySvmmookw/ZWvlAzbaCgwj9Vohc+RvuUCHmVz0Ma3OPl5RTboHVF8SLoXEt
OZYi99urkcdX8s/kz/fl/XwsjbKz/bym/9+Q9+QqyWL5txRlsO5oZzgwSOmgPWJGmmVTE2/+HHAv
/Ze7ENoom2L8BWNOZ+E5DGcUvJ83yre0dZaWbJbTp+K9zDvFCHkn+hzQS3zcgfvMKUaierGC35zg
I5aOfjwO6ONhMpdlrQWcamsYDKSRmvdcoxwAaoy+mll1JHQxQL7jkfT4lCOvFVKD5f/RayaXWQ5H
HmfYFzgoR3U1zKoh4Ru87I3MsZD+1OFsvCJvrH08O7+jknc2ylGF5EyzQp3rZrBe2EqrDF9Mp3Q5
i2Tj+x6Gbm9cKL3Zbv7LQ1wXiG7qpezP+m5QBc0PhCHbb/fX11JWY+eXOepjUycpZUtLKU0wVUxC
Ja2+lGjZINw+7Y88XnrpOZQkJj69cTgO+Lz97sAdpwJvFuUEih9nzsWRhOQzTV8qCJ5ni9pBJeVT
FmKgs9rXGbPWnxuORRqjH6184Ji6GWHC9zl7IAZHZltq8HnkFkLKglrJSH4axB8n800wWk+g2M5V
iDMkAk73DDmKSZEooh/KEFLTnaE4ElvjIbs9+R5Kk4q1tBa2r5N5WJT3gSYomhMEVfbD3wU7WR1E
WFIoD41nBt786bSWcRD20Y2DgRBHJynD8PcxGQZAj8U/p8A4JDAoibUpmtZqGldPGonF2icVkzuk
bh+4DRZV3GSqbQZZgFL7zL4woM5TzGPjqiJ33VBurWO9wz+3ziN7zHZqEGreH9O4zEf0Sy6OnN8S
EccqDLl61f765M6WnVEF8DwPDKpuTjNgmE7BVrOmtuPue4TCocCX5CtYfKwm+axKyKe/Q5s6A1pu
gDOG2lMpkaMxoduaIrtoxU12JolasWr8O4y51tHtChL+0Vc/WPsM7Cv1vPdRujrC5EbUTtfDwywr
2fABICPM74lZ9iYv78FTkuGd2v1dkYiFZLrfO0kIigUSo2oXExjg28aE1B+EF5e+NCUnu97mf0We
itAxEV8BAgDOrJpMzVKb1qou4GSiE/KhjP7i/YcZqm5pmmzE2AildSooIjv79pXy2OtMQJ7DYuca
t4fZHy/Sod5ACCrLXc55ZM1tbMAYJJzGLc4wMjI3K/NyZKlHcFNhXo/btWJ7IVAgaqMIO1N18Jg5
/WulA4m+I8EJgDnsvwXvnQXJDfxVlBS+LMiIBu5XcTkMj4J+x8i/GS6AVs42G1psv5crfceouVhQ
pg539efg3k9wBqZp0xFnQJYh4uPUNrkyOEDORcbiYYHw0R4GDrm2gdzWe/UpbUUltwLAmT1sYqsJ
XqitcowLAgBNS7TkTxItLS/A1Ri/3mUOGx5cEsc9xTPp7pfRRQpDkWJKH3QiQz15TUJRDTNaZ9Ti
DvJCkHDFFHx2Es3mOoEU5zi8nFReW4FEScuX0IIXPrebyqmJ98DVOJqeCwq1ZEyPEvO+0OBZDOZ5
p1zSSGw8teajqreQKOPXzcB73dSraS3a3JvZ4x+ppRkkkqUuHQCrF9t7kgghPvxBc5w9DS18qs0X
V+BWB9V+RgpvHmN4NsrDB/9FLUoDw7gSm9T7zH7BhiIe2W34i9/b3laGE/0OMqDHvDEiCZYvth20
JOezrigJj0MUf2j6WDZ8F+vYLw5h616ekjcq6XnN8QVkCZv4uBz6mFfiHJ08lg+Fc4ODAFEzxnSg
YDNazJP7X0hwlw1MIvT9NVmAmRTD8CMC4NDhXHfUaIcjv9MO3KNUf0jSAfcPTPLk+5IqidmGsxmi
QwKAPhOJbVaCba2/24AzmGHLpRpFQ4iNRDHk7rGuLskBfyC6acm+0/FcZLfXTKJG8UeCt1PqI9xR
+Vobb9dRYeBNuOHJZxo4O1ymrIQ8NhO27mYI5J3SFaTqgfWIT/8lU8DWqL7Nfk0Q26Jj+jJj/VR2
m+0StlUHbeEYbcfLqAcBVI+hUkUIWd6fWhpU9YCuoshaBSeML/MIV4IPivw/te777ap9tZZDhtQR
k5hisTloNmBYSObP9xkL5KRBKnXhM9fF/tq8SndNsXIOgUzOSxW8w/GboT+RULLmHIxUIoQ29OCP
122RLYK2nbJ6NRsd2vcOYbvnRmw1H/nbNvVHa78qDVlRb6kuL47+E9OJSbhDNafalWOZLVcAa+iQ
4VjLRWKo/DgHxq+ceIm6KlQFVz9NeJhx5/DCdZtDQ1ITXTCcDCQPW89c7bleUSdhifpxlCqqcy4X
PmAv5H8J9aUkUgjHrEVp0DQc6Eyd3nJeZlr6muqopCZu3y4/Jppo5qXuEBRf9MU87LHwBP8eF82w
/whw8pg9L+GZZgzj7TFPI3xcF0ucZ+d7Yl9pp/KR+O8WnfYqe5llmAZ6vVRNdgKSkwoe71HjFokj
BF9IPZMZM6kE12fkUxsD7crXsNcmgnzUNfjPAZc4NU79CUULQudzq5yZZczhv6+ULdeeHQmaWw5z
tF2udtL/hzYw+gCAX1oOgjX/r18PBnuN2gv10JjQ1by04VNpG3JWqXCC1Ln36e8AyqL3uqYtvonj
dn6kTJnN2eVKjreEtME1BhuPF4ynfBL14Ds/Lf1ky3q39kuJ20Vlvp+YanhqnX29SY/me3ty3efz
V4c1YFGrcJtiAzwg0602KyjMVEz4+3kINFp49D52QokMESpD3SQmTNf/usuMuFhdYL9u+o7pwnL1
Bnvav0Qlr8Tt/8XbxSwhKMobXiwR2WwrG5amYPu6uEQquQY6xQOl4IObVhypT+A7DYhgm82WYEs1
Oh557DjGR5lzlG8eTbhU/Sdd7iiz/IlsMaoY5EE/wX3Slblafm0C0jJ3UwGYTRaHZ9Lvg7m9XDPF
z9tpccnKS7UoTKYJG4/hfIgaZnhEIdaGAfyJOmB3vkgXUzbXLilYdXAAyK/bYFu9hRVXfYN8JB1J
zZdqHEHRzx+sfIgiwJ/BLRu05MsFkNULOOQoPaLrwUlV1Wq53j7fXA/xnQmvtW2Ga7ExQBDptM7V
0fJ7k+E1U7OgqfAjBeOAvcZGoV3mu8Qdy52wfXbSeC7wp1kS64EuQvY+q7eCs/H1z0iullS0eWUs
qGolDyHCrcsGavw5rGsj6rbJEzIm7qt/4wpcooh/chQg+F2rNCd/PtlLSlNaIYjJY7FI4Q8I2AaR
LidPyUAhCWNIwYRk2zbjwTNUHHimILSZOcjCVQnE8K3AL8Wt0Fe131aX7P73FaXvlqJsAux3vYte
L+KzefF4WIXdmLsSoYdnk95mmr6Wdb/yeIhVLtCvq6ELEOf69l+nwzt7A2T8CDmo10eR42TrCIBl
s7C/aWHdQ+XPoUgDVC4JXDdISXUnIwbMvt3TaB9ew65b67Vq+1t3mCC0esJtsstLEHOdnPBSgtQI
wOE0YsXB7qWZfIpfKxepSBAaQrYeWmWJVY4Vkj3DlpqcfnHlexFAgZ2+Hbim6IPWakZX+yIjKLhm
0crFkaJhxk5ToRudlUxczwoRzwagumgWQGtPLLtseSv7uhjBMv39sMMH4TjRHOg2NB9xZ3s0eux8
Fy7W+a2t/vPzTD0xCFagrJRP+3RPVrPhjW58VdaIrffnhvYWsbW+qU1yiVXoNLSRoJh9ViQLhd5C
NsZFfjtjhouuZBjjNEdz3Mu2k0evdwSfTxOCFdFQkS5G43d82nyYYSYMLxAUxixZrAWJynp5yve+
CRAec58QOOUI6tAXQcr0GiVA/g+Ruz7EEUxkIYfzAERcz7fN20pj/2rAJGRZqvD2HcsuuYozXY2G
MrWPtyNjPgJylUXvBgBRyghFuCXIGTumUbIdsR/Ie8uCA0/1tXot5M5dZTEQp/vx8sGX2u10t2QF
aZ0jV20u7DloQhREC0hdPLCXOg2DXEoLArLZZ0qxwzlfin/9UxQQGJ15yGvgsMxl4dj/ctPCPlBl
uf6mAmhKmDuSR4iHjEWsr/nW27NSGE7ORPRmRbe2M4vceCdFRqFWH76g9IRMAn5RzdSvg5s3S9fO
jmSaeNRpdlIzyhulcTLpZrLLtJoKRHI+o4xnNNUKiqPEiXWCMGi2QtcZtCdsHx5Od9CRi3I09XRf
sHLXpfvxHU2V4D9MQdF6nAVScEEM4ms8pKnGxyZ6DG10IS1p4aSZ69YMoHqweGITQgHRPvP10PD/
WK2ety4giGqoqsqNr48SnIvwCbRkh9hxXghhtkLh4DjlWWFsqTu9PIH2Q8EtjuAgZ0RG4UGwxpvy
DfPl59ALuezLJbDM39bzPOCPAVtBf20DKiEo9Gcd9FUxvfuVpznUxUkXPSf8SkPh5pVQqEMGGc7F
fxchDVENme+qD9mebDGJ3qN/4Jk02A/l0vc+3kNYxVqcdUlCnyoOHYxnPPiqkzdasa4KqXIWikSu
mWqypOiX2fyzEKs5+GvNlGUw+yP+2GnO2CUIRS3UA/kzGbWIC9Zz5tRH5SwHSGI7AaH9m9XQra+S
oLM7Q55VzoEfZnEWPGPzHzl420BjmTgwM0FlpFpFFHR5xf3FocGKrMi2/rEdiIC3rIN9/j1tJDke
HpCp09iVRKk6uxAupsSkRPMbDaaMPg4XmZlJYPJ7m7VHap92tr6X2LbCtwcZGRuOMeU6xb8C85p3
TMqlVHo+PvGtDS9AdVIVjIgaELq4vPau+YG9g8XkZU8l5l9mpbpbofGSKbJMdwoF7gE4Ac9JR+c3
IrRGC7/9PG3ItE2xpP67HyBjpItw3Da4geK30l29gpO5KDnUZTL7JqSEVipIsI5ZqF7hfM+Imm8y
TNov0f0ELl4+a0n8mOH8I8v+Oi1iGRyHT5xrJfhTIqPVFQXJiEn6CFAm09MllKuIpHZJqQu+LJNq
cTlol4HVS/+cy5Szkww9zHg4rLWyogVjy9Hh9Ki/tmNv3LtddAeRn0Q7pjYCD7vswR1H5GsKzU++
YGSmJRBjD6kUadmscNjsAubTlT6AN4BwBFbl2qTiBkxkwWlksWxlURsXd3ZYYS/CwESyRxQY3NkB
JcYHzJE2ZE0HgDd52n+4ZAjH0Ofh2B4k9FMS0b98FZX5aoxs1p95vb4pmA+M55oNJusVLjC0sZl+
ZRBkwZqzTwvaMmlANau6UkWYuPmx20P6ZQ2Md5davhaoRqPMXyUmKaHjzIze8eSAikwQ+AjcZF2c
SQSp3//PTqTMWnOKNN5X/t3lYjYn6sTYfaY0JllJdcztZjgolIlC1H0oDJTM7ycpHnB3Cl5fbrx9
Nf+nm7aI1Hn9awLFWoViItwiVWEsSvgG5JsaNrp4WIsJoxmT+yfpofmBe5RBgovkFgoqIz4OMUF8
R+vCpnrXdYVQCh7kPVuDL95fABUpPeYi04mx3Ntt5kbawrFTSJpYOLNEXmPErdB79kt5V/pP9oQT
Xv2LZf2/V3RkDf/RqlRSkiLMNOjhh2U+KDpiSRyUk3QKs93aFBo0uqsSnxlEDmCcB1RyF/teKgxJ
6D77r8Dv+9ayex6me2XOPHM2jEwL03VbZzhkk4/PIVzru+8WUD74Yvfe/L5z9ozdSghPhXiugkEN
A+3fLlJtg1DlFDt9KqcnWuOlRvK05NTR8q002R6Bpon0QvCNK/eaF8zBpn+4vFWIbqgto3I7E38Q
x8UjftEkumayP2KVA9X//wD8rPbWdn8IpEN0p7v8ywkp7o8fgm0A/VRgXXNzIzGcMhX5X9lnjoRx
bngdrHaj3UPYnMwgKlxMpxhp32BvIFyHZWh9Tphq60CzWxSW5X1fxvEy25AKED7ci6/PriC5UjEH
u3AoEQC56j2r6eGbhj79/uijIAHMPy9SCIogFDVTFhrMSmTW0bRKWygY9N65wIdu+64N7gdtqXso
bGQOrRKBlJxVWRSCVgzUJ8Z3hwPr/4UVrVZz5q3zATZnTlqPl/s52B6KKtRV2Ujm5gpwXYEQ8QSX
7PYdycgTD05D0tUFNHPthAzgGO/CBej6PKzYNYkWTMoiGU3ThkAc/M+Hzljx6hn8MA/tqtNPvcyP
MTQ0AAVHSyAcyU6P9rOkXN1DgZLieF8/wO/AriqdzQiKULfU9Bj7d9W58yqcTTqs3zdilDS7KyVc
q0HKE6XqwylxZWzw+/u8a9ITTg4a6SYhGynOZuFMircS9cQFj+0sJoCG1Ytqqb6QVWyrPILhl/XT
eav3LjAdIHkFeiVWRgHQ/qtxisYid4OPESlvJlDH59MQ1AQvxN+QRwBxYHffrk4qxvuCcGvU90oh
8DmZZI1PEJ8NzDvGHx4bqrOWKsTHOrAh03kI8AMYMuwvhBc9AiNNZ+0TO6AvNlqr2HgXAr2i8ViB
cw6O/OAollxpF4E8zhH4kYvyrArsMAer5uD7J0v071A1wAwN5asyfOMNsw9l+2RqhQ6UFfIjICfH
GjyDR2QHC5+ewjsnIzUqWQyyHNuk4qQ3FnA5xG1u20GaWSdBOa+zac/v4YdrrKJbR4ynlEB7b6Lu
4uW52tPFj4UAHOsess1zycnZU/nA1Sj3az5TLm/V8scEBHp6sM93Yaj4kWlIfTkUDKNnJc61gODR
mdmWzBJGQFpjAYLMkEqjeqKgrsL0Y2J5G34nd7x0cLeFSa3HgBD3hG2c21zHvTBIVZ7D1XecUGrZ
R4lKVdNL2+YCeji5aT04KqUEV+OPajSO4xyZSYAz5Vv5TOzTxII7ciM19ym0ABer6BZ4qUmdsaVB
3oSCnszF2KXOLXvRdD+pRfgfKX5hwVhCSTXCATSMQJtsBI9cOGgcc0QXaIEtlFwvMnOMRs9qan+o
tSIhlTRN1IOHRDbJyfirAcMhlO3qMi5j6vvYRYHba3AV61Jx0tQ4mpak7aTlEb/GKMvDu99nRxVq
wnAOtArgK5NdSwb/VTL/tC10Y/GJqYXQ+xcZmW9UXgvPbGKN10AOHBqHANOJfpaFkTPI0bocLNWL
8TBsdvMScszIifN7er0Jxflqsdsak6iUJCZVliBctfOtt0XRtTj+BmmxNEVWxO5ZkMz/k4UWfrh3
YZuWA7w9FQC5hcik4jSkrwLwjq8CzML6toKzQS0DKw8oH5DDUnepINdhyAPp+hXGVtTzIJ5RVTaO
xn+npYvr35Rxq+aN2tz/LEO/EmuSXNSITxciYTVxt7ExG/OyOykUr7EIugp6Qs4ajRPiiTir9qF5
OBeLr7tzOpULZ//ibUhunHqcJ6dIB71KfdnD6+zRfWbSzs5wyXjJ2kf5MUr5wvlJSmbQKwvcTN+z
Zkil1AEsfMOKvOglolC9adf94++NmITnpQHoqtMs8sjOZ4Qax1gMARywKPww52nKJl3xA5xNGHVb
PnaaBBiWU9qcVWOB/sYdYPqFx259zP1z0wJUoMt+i9EJAieFcuLS6ZPBJIxDT3Q1zQSjXNjbdqnD
pch7PdcsmY7GMLC0KSM3xmJaSejxpCL6NctApfA7AkePSI+hFgDXkTyG2002L9zJWF5rUdZJg6vt
p2B3tB22wAnKgWgJ8e3pBn6cW22/f1IXN7qbQt4Q8Bqcsi71t21TGlcOO8gm6yVkGaTZOsXL4krz
IsNxfbxFofmFEn2LTsnxu3fGdNWw7SNDaGnksODWImzHKaH9yCPFCLgxzO7Iq3oUBSyREz39ndWQ
qucmt64Ov870oOAuLSBEI34sM2rAM4pbMaU+pNhrWsKdKejXkaDlgpVgQ7JXV6aGJs79GH+vWAAp
ga+XZzGfTFdxIWgISTeNtvZznKD7yabYCyJ8W1HFYDNHDU0dD+7ib6EyNeZKElg1e4fj3/LHmmZV
lpWjbO6qFVWpXqeyFd17iDPdTsXXHtHWBunzG5zozxKM8Hvu36SwF92YOgB5Yq0AMQ87PdyzKRCD
/mfyDCTcUeUA9azNuC3cqDf4Lg8atlBg6SIT3hAa5X7MuX4cnaH+aYWxDs4y7fUn1lot2R4R+J4M
AJDsKH1kAssp0vE2/soYW6Mj/0G7x+WM1Ry/x8KSVUniIGhGfr6EnCkSMvTorMJa6INIkot5uYkP
oZPbNVYyVYiL30lbr+AVI/RiNga+NeKBf27EW64S76QdwfX7ViHTTD/QS8toem+p2+Wmwr3qfKCc
s39Mqk1xo1e44r0biSdxa4KuVZuiocyUiHtN+/ZGo6VeEIzX4rHTVAbdL3OkrrD6VIdyxGl/Id0P
ODCdqJjaKW/pTJB/H2SYMhcwZZA5xduoCZbuuVtx6gxZqp+cInkUnttx0qXWcUh4UKhcOTF3b+dL
JfQEQq9LN/L6LZUNDcKujM4ajySuUupflaxvpbUweeKwuI2D/DGEIpnsMndVNcOtKCzzFQ+H9MGA
7KYdRAi0q6Oz+8UMqkGer4v2nqQALZtV6sMDR8y4g45Y44uriby3nkpYRjAml3B60ijh/+uDG6OL
xbm+UZlfPNeBw9SM9f14sqqQj2PVfxPwnzHen0z+BySx0P43wMBb4ZUN349G0Tx2t7Z1xRcY4lXB
nPtbuQCLzBSmFtrOHQr5efc8dBm2EUrDba3/T3rvQdr7667oesyeyFxt9dfxFJUSfP4s1sezT980
xvlv0Vb/B3oCnzkOhnDr3mnyi71PVuHO9mM0OEXAUuIeVLqnRII7/A8Ij64UofkLbmxsJRNIHFf7
VYXrGNjp1hzPCJTQvWNm9K8IatuMLiBAhgWUbHYJa4RkHSXr92gde88IxGqkDTuwenYaqJBFQk19
I+7epeiaFjwXjniso7hJVjA4P3opSlUTe5r01qYIU8H7LCS6Nym9+Deus6zXgZ1R17Oh53aWJScr
fW9DffVVWLTiVN8degQr1dFKOYXCWnB5Ftn0BLKkkifGTrI69nQGmifVwKZ25tB5Cwd5WPXYDF4M
HiaKf/yuY1iXg2fYHwekmHX7q+0adlL13z/Arra6kI+7sSUn7L4ygBxCBdV2kpRBfEWNs3eBoIzL
8o71rz8s3aC9SmABqM865SJfME22l2mToLbsRUXmuWomQiGDKPqFuYwx5BgpgLNrGYbGe5IkdcfJ
S3MD/jJrny8EGuJai3phas5taIp9zUei5GOOZZN696gpkPqAm9HoBQDsa9AUEbr8SFR/c6y6CUbm
5lbIVd8g9KfTQE0sShhdFbe9d76YLmBpy04BXxpjura53WhlqPH/msvklj6o5v2IRrOupfO/uWuS
Fg/4byd+qTiNWymuQ3xD1Ealj/tgb3y7Vx9tgcKRm0HwXfAp9GiUbtgGK8WqTnAZjPlIVJWtNezD
jhQmFmLYnSRJWryfGvriLspChNbkkwlz9pCYnnh73nbjf8srhiVca87CXn0mJx7IeWM8D0zX1FRh
i7vSi4QEL71GdalnKjMuXAJFAd9zC1viUk7vs6r78CZejihXudaBXRtMqiPb7ECzrSe0CfhXQqgC
n6r4+88cddd4vXikyV/BFKrr4klU/2AOzrdy86xT/c2hfrtZOLKBFG+SLaO+Khxi8JLUQBPOr73G
e/YetfVZQN6dLQPGlIhM9emnnLC/6xBKW5St+zStb2AK8naA6flGBcMjfOymOiKKPiOo0Hja4Coo
r1jz3F+cajFGZn79pXz7HoqfyFpxZAvkOB85QtuxtsH+2Q1pwXN1JULyCMMBQ2x0ZWG0sHbo8QJC
GcDjW4jUp4w2nJuGIIRnzw1Sio5vjxlTm/7fGvLJIgVwgVbsew8IdtYNCpUc09LE8hHAPPdF2+ME
Zxa48YwmuFKBh0gBp6RO2yaehPK0CULMOR3H9PzZA80mfy685AAUajl8HPThStRqmuDHbcC+LICu
jUujG5betmq7l7LyG5sAc+mZa8mLQ0FQV49Il1oGp/i1CvHxreVb2ku2PpQqWJwAtX3iZ9oByfyh
r0/2b4aO+O9BhkgkEPbKTTnqqK8J+m3fNwZc2OGd+rJolUg68jSH0Hl8cOpOSkeyjRAaln0MFwBX
37p1cIIWnmg4iP0slPkKpA7Rh3tXx+5XjgxXQOxTTh8NKhAx6OBGbIAl3HX85e55bvGlokVmQMit
Wa5dHTJq5ushWiv7jXb+GepY/XooB1UD4IUBp8KUKeB99w2uZ3W3UnFlRRNC6jibA0tar9Uyh2cf
NizpfD9GUup/aoiGG5BIU4UoE3Mol5J2apZOcwvfiNwKcYSGFrSwGZCNxwcrOJOQaxbOwNy/RFVY
4aQHGTUPViCEmkWyNuT6ZwSnnFzQ3jn0fZxe70JspczMai6c7PSGaZro1FKeVHO32brSpdE+gFh4
DXfLK0uyqOsbQhILKRx1usu3HFbrqr99XZwyK3k0EJqFJMIYv5Fp2ZlWA21Wl7prlQdWsSgoDZvm
Djm42ldaX0iXvsi3Uu11YLvuJL/ECgPwyeTgDETwhWetnyK7iR9vR0y/D+OOYjD6mwP+uszaZA6s
CivBtdtLC613rMlMDlOxLR81dLBwCYTGg1ARWSYo5lJaqmlLdgxhhpu2BSCYCtSTz0AxKHJ71Www
NFSmcCcETVSrxNPypU+7L4o69j/jhlL62d8o2nLmXVvUVd0EhserI1XmShMh1gJl2CI7brkZ4Fao
3f8WXH1Teqdh8XdjSALxwFayjmsz6lmsrasAYNU2WW5YlgT6yg1CwFktycyXqE5gCWEXwr/13tHG
H98WbAJjjDC4CMygdZ+Bm1eMJ+joCNZl5PmFQvHBU9MLjawJJbmJTmC/b6PtfhvH61+7a83E9WXO
L2fae+AZO/+EWbjW4VbP4t9kHqBjfvsjvbvFZd5mLR345sFSvvVjHYsPsAcowRxnu2pOHuS2fG5R
n91hCJIdNbWea+KjA9EK5HftOvtmU5EACSLI2cJdEwcbShK+UJbhD87/IBsz/PpCNfAEJiVsQnr8
ASi1in9sm62N+r3bs2Lhg2I7dJsbYVl9xWg+XAKV/3KIQY0H7iYGMpsRlAxQOEm+mBSgYECNt17v
URSop/HoV1YeeVYWcfunxISDypx0JnEyrr4Zg3u9Hzp4lFe0Hj7yH5RIohgTzxFuepMc6h/4pnaj
l6c2LXp5hd0QIhRycyNRV6n7+/wEg0aG1UI1CT/Vc5XgxfHk8NsSb4yFjXm1UT4nOrbip8Sozos/
PiOf8j/PEACRlGStGfcTCKguL7tZ72Dpea7d9+brN1y0gBjuuOganPLb3oGKhDM1FnKLbeDV4vuJ
I78usYtVxEMszTZ20g6kKkkYa7Piqz2p0pyrb8Px6NCpj5WqS5tBKAtJGJ1/VbnNtv6CwvQaGk9z
XUbEDQjpiyrrH5pgZf5iiSJdy7WLa7PiK0APZu3oklgDC+BmMRWmAb9nyWt1S8V0hRZkIAfpmHVw
jdMVwePLVXntq2DDliCIW0wwagjcxXztAF2zIoZNe3kdPE/v8M8r9JQApU8Fqus/LHxw1xxym/H6
lFjtkUKddvl1x+8gurUPoa+9RNe2UJuCvJV2TwdrjqPNaQ52YvJsQ6B6G3CGGW6sPLN/FIubURbw
Ud++etKnvGuVWzFlQSr8eHBKim0Cca2U3XsBmFmcBvOK5BXotJIjnYTKCLcO5dYCt9p/4DbuEQl9
YIK/WOlDtJY7JiF6duKGNV4JaQ9jLKc3GVm5W9pkeY1Zgm72+qVTfV9R1kIP/vlSrChK7oduQ47n
jBctcnZviO6VFKLT4HsnofpNpk/OraKep+OnPtkWF2P0ip2RJyTsSZvcNkQQv0U4L+wf3KeOI3jy
xIhoQgytMTNjJSfD9Xi86e8o5mn4eOsSlsrCbtde1es57G941SgOktiPdtQa/BUylD4H/bjA6ykJ
QZnQJ30Rh5yxGk8IPDPvB95RC4gr325iqzIa/HFasKKY76/qm9j/nOqh9q6VSjKn08nBfm31jLKh
etiejAS44X+L3xq2SSFLzi1yW9amQZGTAFUkafbxn3xPWEna9qOx0mGgoB5KXAdjqzUjlq9wu5Y8
bAmu3orydAB6vEAAenlz3bT4J8twW5M+7ILbNlZieYl0XtisGUd6q6WmU/0GVHQas7XKFoy9GeRM
cH5pzOz/YYdYbziIdznyK6q38whaF+wzdfr5D+qKNa9M1NdASoksr4jevACXXK/4vhbgQ1NVls13
1dWb527uOJ0dY6qM+LJF1XJ7okZ10cDpmT8n99wJbX6SIoKHrCX1mOox4nn7jeJteT7xsdeFxkT1
jWS63q+LMlyBBdeW/jDWdNhlt1qqpiP270Uexbv2SugVFyMVTP4104Y9HqE+VhqqW5f7ge1/FI7G
pCsdRiA4JOsdmu+puyDpyQdLPNeg/21lRFnSp325LlGwLZtoYRW8aACNFvOa9J4rfhQdVNJuIMmZ
kkFCOjOdjLetb7fFa9n0LUyqJRNjLUFZA546SQ4UxH9Q4/I7ZnNQZVmwkIy+DLtF0ElVGZDIwICr
YYfi08+XysQh6keKvNUoiCUzTf9QNxyWo9H5TW6eWOJA0aqAgGgDOyYVO18Z8kzvU7U8dlMIXc+7
vH2trY15I8FQZlSR1RR5mGQEJMTPFTo1tbuVXbUyhkifT7UjTV/aNiNgiI+mfju0RqofmTIyJepR
lCfA7sxS+wGOZSOkzUVDU+udm8S6lJ57XytFHrWM98p69aM4dpffZ2zF98CuuI4kK2R6qTmN1dK+
RZgzUUdentvcsmyg8dnZwH5DztlHyB5XlpOFpp7gq/iGX26tQc49g9kTvSMCCPw1lUTjrju+i7px
7NeTaHw/kluw+uM5jMobkIWlnIEEiGGEQ3HdfcT1r+WcaNprcXyhqbalys/TuPrIqsBu1mLN8Qu3
4Nmpv+no7IsRZIkVg1hVgs2bmYHR93S62yGCt/eQcvk6Z9x0CMCrT9pi9vDvHBKvuq3u+ZVzfOL9
DkRSFLvRSyLa7RWedP+wBJeGlfYzKdcG39M7DPIjxMWNgT16RT5+qbhmw0VlFW+m6qSHRyBktSWU
wOa+8yYav2VqPQFDjMTJusZv5ViFzmFyydFkHGFw45vreuxL+YMO0dztHXg1zQdoWrwiMeIlyJJJ
MNiwXLMlQLkKgEKcIzDOPEvDIHqRaFb3SnWmXezw+BxlzFC9eguUiCmLrR7xTgbXzByOOqAlLUuq
mgzeo6wlkwkKyMTgise2k+uhZHo5jpUfiSSGCqCK3wKwQNmhsgi8HRMFNaCpAB+cMnAVm721RkXc
d+s26aHSTRrsi7t+HjAa35lHG53hCpHUFxEzZoIraARt7TfkcSLzIsHqin6/+ILob+T4A8OwYtSW
smMUMtx1nGeOv10CLuZWEGeInre9OE87TGxawjUU7rsyqoHVIUron7Tr8VdNj88EGUk26eAGEZCh
jxnye/QoOz+g8uQGFliQkLwXLxsOIxh7fgdBA0ac3322shcM4pMssshkitE1txN5Ioc8iYvV2a7k
qcK76wrmgbOz8iEywO+zO8fyv4Ff2phTw5a6NJWwS01tCr6JFY+/7wsSaOJiO5pVPY7Pb/fOlVEM
E7wOBTNHslst9+9VkwNA8aB+3Q4/7HhDlFXVp3cPi86AiwvRSh5iYW2vthQtH5KAg5bNPisFRKgQ
rTGi6uXJ1g9VaWD4E3JL7pJqsK2FaVg61hwtF7mrbJ1s7nlMoJEfUSYwKbwz59w9jcRUgJ1Z+8SV
8z3pRAtTWzaPbkzR02kEWgCicTTOpHLt3THGAwE89lvNkjq0235SAqPixkUiQgpKx+dQnE4pHj2C
oYw+nCSJiuzxAZMe4jRn3BZjpDNgFH2Hu5TZMhJMvrzzMeMKq++DfaBUxxwcfYSgfGGwtFViVIeP
U2uWVVOr8lY38Jyg3CXQULN3uAlXiNlMwKAleCKK9NjLo3e0z4Db2bh6e1y4QRzmrrS+YpROLf+r
T6iU0zGde63XJ8UYiGp5TGG1CPGq/fUMo2zMnWGUAL0jnGwWsTlynhfXgzlkAieXUw/WAJVEagI1
VBKIkzbjCDfMZ7X0p+TVIBLA6Uzi+IVC2AgFJ42a07q0JlJLbGu8FuMZrEYPW/poGYC8eCy800df
GLOflqCqb7dSdmK2upQzRKEIZiq8VlCOcaw/IGrzF35EpR7CWPP80VlYu6ZcSc3Jows1lU51s6Zu
V8rk1eGun1ea+IV5v6afjT2PnEbspdPgsWKgpnCi6AfcyVUPl4+F06eNaMg1Ed7nisIU0q3qsSoB
BjOiO7YMPo/5ggYkhkgGzy5zqjzC+MScc1aB1f8I7S+EbpPcZa7VwLANS1t9WhkEwGdqo5sHG1rd
6IYzHxhXwv6HjsI+upAcPC/jr94aGDcQwyiYYKoFARZgl4b5rzmnqHe/aQQMgwqE+IDtXn8wsRAv
tVrcbHqM8wdgviZ8JetGZSP35kTpoVvGsLm+2AIrZZYRbkwTUzscxqnBbv8dqOUOcp8to7uCYV6Y
ohUgzfDr+yInpE196sL23OuDA8OjxI6PZs5bPw4RyLNjVPisnu7YLJBcfw6tBXs2OzutlYbV0BQ/
i/OjeDLt0ntYmL6Eu6aETpV+U35rEfiw2cu7DA2uyQkezNnEU7vVa/gbFprnqs9ilAfo8HZvQ5nL
fflKN2Bmfl+ckFr5zKYRh4GVkabds4aA0Sf7hnkH9KCy7/GWkeUrLArBhmrT7CV4d5FBWdpZL+vQ
OAesqIiDTPX3plyvGX1qGc1NcYXOE7qIyd38VWXFyHxU/FLl5k60Pw6E8kjhfJsDfYX394pyVzU3
FM3oppeBgHSxeUbfhxUoM4k01A5hTKPrkDRqIUZQceeUZ+WsKxAwT2Q2mvVIF9slCmV2ev9/fmg5
EWtqcIv9Dc0D4OhNghFFWDbIFj1lNh34T6qVQI/kCeRyQal8Ls5TbKgVmtbhUslQ6x5ZAq3lnzrO
YJ6R+9Hbq7W9jD/F4YGLf2VpMxhgjOIuQMaRGDK2XYvffdRgmNJ8b/kG/LbevkrE94rqOqG8C5/1
Gai5H8fvpFlqh9bAcBU8J+GG1A8INI1OLqaubzhPPBBWoyB+y+V/TVNobtXZPH6hCJpR5swf5ijU
4pKCpbdsHoHbSe9kGBzSAd6fnLyRilFxirUefizmEcTDZeIhZSBmP2lRjh5CI7rXcaTdp78Q47Nw
KOiMxZjyunPQTJjnE7vaEVcRJhm4yP18g+73pT6t2Ed4xyIzbODYkRh/allRaHBR4Rk7Ft4cTKJz
jPQHr1gwR/nbaJgbXsI/F61t2eTUruShDxXUCyEzV7f211otkm8BLHNGmD7BukTjviB8ZI8FLmJ0
EG9oKqTOWOtPJzF04NVeCAK7ITDGX+mDK/6G88/73PnLQcVlyZ+Rf/EnjNV6GeMLeSItk3VFvsg/
7u/0jSTtJGKsnZH98CwLqYOhtoRUPGvRTuHmQbxaLvOffZesDUtGNXOVTtYzMJGJKSARab2qKvux
V4AI2DmGA61IFJDFso8Gc/ILrwRPb1HFq07VJQCW6qzXoCvTKVLDJoQbokW1ltF7FogErJHAn3be
xVYq2SzGk5EMHRVpbkS3o8hok03hgQsWDhzLPUh4BhFgyqs2z0Wd+1yQYsM9Tk2ICKyC05STmkna
Yfp05ZKhQluba+mpuP+aPaaVqDxDe38F1z0emB/DPDD9bzsn5BR27bMefkC0ZNWSL2gZE6irJC3s
VhaW79FBVqdBmygQZnNRGd0GRnLDmclngmwKEN6tkS99zzVWPhZ+8rXOdNWgzczftyLS7wTLeliG
NLW4BZXisKTmCuzxP0l9uEASmeL3Xi9+G+GxE+l7PcIJoOH1BuO9yKmuR4LksZN9sekLHP1WrTY8
cUd9Dm4FENyYNAoDogHI6dKQPY46BDLjrZB37qlDtSOGwCSpsJSM6GS6LTnS249Qu2ZHStfFFIGD
xmOF4tMoDsVGgpjAweZiwvpwcokgJYBFWZKKU8La5aNmIYpfF/g9QuRYQKiOSKYUNrjlnxwUjJ5q
/iEajlGkvcE89OD2Gcn37nDFuhgvoo/YLuxQs2pBZZ3pDlDdpEMNQCLicVShBlhVAcGEPu66Yp9l
ktNZX8zT/axkhvA7dd5IECYFa08o2dk3O9gLADHrfAuXg7i6Y2I4ZawoAAaCwQVBWbt0Odlv9MDg
0cqTJ1IW17p3nCbJg+qWqF0bzGZTofYrfUqpPOzWBoU3imQIVazt4f/DspfKURlj4OTDHeZHNBmM
H80IqJMrYGCYjJZUb9VE3i2Uar4c6OhvwAYnIt0+DEGX+86A67/fwZxspeAkLt1CgGBvRqhDwh9g
AS5dg7js+SVtG56MLEsby9izD+5gWgScQsCYoJB5qqXNA7kc8MMn7l3DjkW10USnvy9rCKE35NaB
1pBC7DlkZaes1YfTqnJcPMxk09YoC8Hr6iDRW7+TN/jLoeUFUm4M9F7wJd9jvDdhfVLbLNDL7w0q
S0JDQvwhthpQyet9rGRBvmgFgxrukWCKJj5GhRQ8c5Y4JJ6Uyf0S2OkBLo2cCHq4essA6quhVJKQ
TwcBMZmf8fiD1Ww7v1n/9DjFfbaT7e9qMBDr+o18mb9h/s6Q39nMIRcbOCcfWhXWlg6ZwpfFMQYa
/5x8kOoTIl0v5d03HMWYQPd1NpkJp1/EZ3XxggPXnOtfJN3Fjp4uj6016wzf3PVL+UH4yK7jf/yk
21R9CMchne/0HKcHEOhrTUxBVDmMPmrgSyMySJMABwZO7CeFBCbucEIXXUoDe9O0X47uoV1yj/ON
ISpiguSx8Joq39EFiOG3cE7A766axKSz92UAQINjIzGPMyM7979f1wZRLWrm6s2tqOASTDlhPPuH
FcCYAMTUMr8L0nijZI8A2VLQdT6VtH4PwJ5yXtdvKpwGKPgGUGOh7yx5v3Qor1PDHJCK6UjLUP4i
Tlfv9mnzQl9TXoqUktWGqQtUvT8nbcTJWHYjXZsvWQeuL2vrx429m9EhRHOfvi0EaR+zqTwYLrY5
Rqy944gcxob9LRF8jcnCU/058ljmGRtiwQt0idM16A8jnfLtc0goZGlPmPPrxQyNkDH/Qk3qJwwc
va7g6mBfk5XfBSE0F6e95D52odyH6tPsisgF/Z1DJBoSeOJuBkOGRv2iNH5kthiiiPxMCpzIihCO
zei/eqggP4M3FXwFyrGotA3z/SgVQ89DFDsQtNRPPMFzNeAXcknuA72L09MNwIYMpw3Vi9fOuoVL
0Lj6AkYMOnbQLJvjJebh1nIYf+D4bPwDmdIN+I7JFA89074ZUQpK7vLwqNRV1HGwijYdxZIcV51H
eGZR/eAZvtKC3+W4Y0mau1NB7sw52CFyo46yGnE01vTXazsUDP3jl4xB6Gb8a2vwj2PyA4vpEKfK
jsCii/ha8lB/IjUjZ598Wkvj44cb9D3GSCqVr/pzv4GGJ73VITAT5tsD5zfXjUqa9CZVfxdSc1of
AbknkqGkbzN47gP4ukPvddZwstdHyuXyLKTV3cpAwQHfuGZx+u2ZfpRUl9htw5pY+TsX9rgC8w27
Nx4h70KhS7iYTkkwbztfyd4uHHUvL71CvKoMPhAw5NmA8KtunkAvtCkTiYofxd92f3l1Vy2N/Zfz
vnF8JZ9818ps2pjBLsi8Ne4CkEe06e7B75+D/4AbwZTpyhF/qacyy3kYgkwdNnlGIyYHzShxJKSN
sZFfbGxAX73VHT8LTq6jx5j04W7cDF+e1F519t7X1JBhXn39AjG0x2BvYJqYDabgEyiv6cscmNwV
CYT0e3Wnqn78gUXoOJOpKuRiRZls/1vX2PcEMuFRJtqM4q0GR6FnG1kEaTfqJVx3bN6JRYRhYZRp
/0WEIchzFl+7CnDSrUs00PDZ3WyPf/YYrMDv1BOneBrR2qQ46CUALjoFhUg8cvpHYSrCvvq4Z4Rm
a1QcapqT1LxiZmSPoa8BxSfJ5Q0dKpRCJdWnwQ8iE4GTY+lb1Jr810LzCsxB2fKhAqZbxd6qjFG9
Tb59oQ4LXT7N/3Hwt4dn+WCmAUxVX/58mlsA5ZurlRjxtnAvsLNGuHNNaKb5GYy4cECvhKuFvksN
9cMQ6FQa+yvX7GxZvL52/gRACJGBIBtb9KjihaSTxmwr/W77UfWMB0k4Xn6sJwBKK/iWOw5GkbG3
ZEpYhaRJxwXHe+Ls6D9IwnaK33DeqwqWKQ0jroh3pcd9Xc5maPsIfAbSDCudGR5B3qjrXRiMCPmV
a5O5oKfX6olyJHnzN3kKrsMgmgstHDVQihlJmWMJQuDJ237XhN8ePomNmG5QpV+NepXrQf1GmLY1
GGJf3V/4BewngmXHVsrj/o0609DsDh/9aET4nGctBN+eSwz/JyaUJ9v9SgZSRCjtRzw6YQ4V3JMM
BIP87FkxI352Rk0ICUUsZJMtpkLtiJlq6i7xaJaCF1ONHVRw1phGs/WafvKw+2y6qH9Sa/4Lf0Hl
nDBXfAy4c64KXe37iAWBJ9P3fPKhjqayAB3n43l11YMpCBOZn9uCOWEfiksGI6Abf55BxivO7JTr
pbtp/YNSvWOv1uB8ZIFRFD7Tn0jHaoWei9tactmex8/8gFhQwjGbenFMH7tRoU7ulzIIo5CFc6E4
0jzd6zjaUqo41IdwJYthxG1TfAqXIqtnQo7YfLrcLV9ppdM8bN55c/me3azhAodXArgZamo56lNq
3yOPFmd1HpuObiAmTSv1XCjjLoJ5NqAvh6aHzWsjoDe43RW0mHzarndy0WVwe5E8Xm8TBk/h4HIM
ukZD/f/cNK9tWuZB0eQPFEl5G8i6YMylKUpJ7IpeSCaU7XyfS8VhzfXXyvEg1cMiWqEydoHOJA22
aBK6b3RuLrEJAqbBGb0JmOtbClZzFuA1ThmXft9oaQ4FVjlh8BwurUVTkQFDz+qkKBcDZvxZg/hB
m11ogoAZD0H1A6M9sSxHeKB0I2Sr0x6e1HRQNUDtIiRfeTjo7f8ShmUMDVza0jXZMo6HfD0eQW15
XtWOlheEywuzvWqWVlZ14FdBf+AIAR9fxsXas6oG90UfN5VvirJNRljXDC1jYNOr001wgF33uOef
euabVoBZS3PCd8l2Y9aqyG1/NhpRpwOpB54ZJLwWPztg7dOxtMWL43HyAZ3Q5PsrzXYF7YwbxCKi
kUiIujBKwIjtq/vY+TqeUcGKxj4TruZOrJ4pl46rEIEmfHwBY+bR2f/KEfxEW5TECSn8FX7c1Cxw
0i0UfKm7m0jDMP9gM7FnpQu9jrg86qJQRqkwK0Vo3KMLzrEQqZ5lyF03eaNJWB6yd3BaA61Df7yF
yeMKJOMkxaDkvK5I1FXja/BWcMLXJEDIrEipCLVfqmGsm4WE3lMmwXAj8QRqr8VJbLXI1eLem2gq
+KtU/XsxRPv0m6FHzKBA8Bi11uyNjyOY1ONShGT3Sy2I68WDuJZnKLiznHU4AvdM2BwkymvQg8uA
XOhA9rlJBqF3wZHiCjj/kxUj3A4zpaRPWNLjxK0hd2O0PitBU9OfIgbx+M7GuxkECSR3vgUOYL3B
+l2L8QyLSLCG2RMjolr4vsYWlZttkD2O+j9x1mMo3hnqr/eHA8puSs7cNJ/UhSpzsjDGYJeIhwEt
GZD9gO5T9K3B2l2v9ISuLt7g3p/aMUQV1jvzyIKOXUAJRRN4mrhzM5Mps0dY5BGQ5Jawuq2vFn7d
VxqfvL+0X5W3/3euWvOlI6zADT85nQL2RufBZPGhG077n7I+nC6XFUnlbN3qasr35q3zJXXDO1pD
oGcVyryjc+4pgyvV73mi9e1S1ZwelxgjcCrPxoNy2iD/xzqzmdSUs5oo/JYDmVlBm6pEq1YxI08f
JHyZaKoGx2CBtUXbcIAKsn/djgXwqbRysUX2Rdt7Qg/7CR6IMfLJKbu9JJoOcnFsD6G9iWEOlzgR
mYbOkANtpI4W+hnH2q913573C7i93Iu1awWKXDrGLMhWOcZl1NAts/p/J+Sps2Tdx38+pdU6hGAK
VE8uBjhYv/v9t+6UAsu3fIVYZ3x1sEewW8rR4Qs8kyD7RPo0HqtmkjmM1lNo3VtJzi0cJNelCXva
fG4An9KX7jtwqQEQof1PwJthrQlmc/POQoid690bx6kR32Q6md7IYbMvjFQ2RWI/B7eeNgIWH/sU
u8hxmHCOhswKy5nDWcSKjsq0NdiowG7PKIwu+v/Ufn81O7FcV4g53NF+71vr+JACWimkWpPc3uz9
BSzu6Rx4DYIMrZBazyOYG6SMk8OYMDBqzd7YgzWfZugqG8WSmxKcAMceawh0ZfOEhwwxyRLfy1PP
5YvcMV528gDoh9MKkSoL/KoLSH8NyQTbS8BYmhmFrLiRkD2VV2TxkVZOrsxRVfgnbv3u16+FEIgG
8tHCxAqr4IPC6vmGVa1nYWonzTp95pSRBxefHeJTaXTOcK8PHrdhwaKCnxVtisZcny53dZ2SeXq4
LvR1PyScBJibbDz5hBujmcBW1XRwCKVGOs2w2mC78wfbmG8JPwEC9HUrWoMFpv+o+IuFrJ8gO6rM
spRwXLuwqpd2NX2dg6/B6MDTFEE8OCQ+tHYImovRBerIZWxeU0dhyIr43nrel0tz6YrUz8g/xkTr
fLIpEYeoEUgU9AiQhwEsRgXYUGi0AIOKAYsIekYQdNW5GebVlkl5k7D2uuSPULoOdlCT4drBwmbf
EcE6lA/yG6xlEsATmBldmJ6EvFPjzcRPl3de9mFbDFr83zFSajzXbH2qxaMKLj5izfpSBGlkA5eJ
QddMGKaqL/AGVitoWtxDTTZocXBAhguR5kPEQUl0QTHUCLefpWUjqyW5Fm4pQhqYwqt0vpc7Tty7
akv4YuNWfmYbEB8EtT9SkXIR87aYJIEcxSmyi+5g4gQpcUvhM4f3O73TNz7rmKqSYypKrHP444zP
mgxX6GKg4Fr3jZ8M1UKlp/8BkE6pxSIvLuhUBsEdi9qa+DCWP7nb2zkC89ToIzFW2sL/4HKD7lZ8
0wtc+vVrYmFwQaDmksf36T2YY+4Fx3d1C3pEqzeAgqZHfwPzJAjLgDsDdmnWE/eRuMrEQ9/k/usI
K0o2qIiXq8Ao6U5L8kdNUBOd1qWZN1U9JspxyKQGHjVTxZjom3uHnOldzCkA9SNU1AJH/RBdlwBR
xzumm5WY5Xf+EOPXLxCX1ub85eaYk+bDJssyAG05ySfIdePj5sEEAhJ8UFE4jNH736+LDrei8eQy
8TsM7X9ZHnihSnjLzfvBa3zFKVt7cDn2G4BnYN4uOg5Fq++3ZAa/u5IF5yDhL6QG72UkGb54cc2H
b3MCasD9cM312SF0CbRrbhJQFFTKMBdvZlu26YkOEQFGErNhC7iHqtWHEDqnDvz1LHf4RcWPIRPj
TBWcIY/JgzkyoNlqDC0viFzaTMG3nRyzQxCVrg0+LSn5A3O+xMqddk4rVJ8FZGf5tC6ZTA8HNMKC
q2wqZU5vHFw7lSTxDO/e6/STxTnTazJgZ0DoS3tKJoT0RJBpvhTxjcOkL1E1OlX4eS6hpeZCpXqq
jY7OojfE8Gnw3cEBGAjkFeQzetZfD2bdAlSEnbMzwhNd/+kTbMVWNeh5SrGtzLQQfE3ti3bWGHVC
Na7Ty7DbLdPr6oVsw0sljVqwuQH7Yej7gWxdifZcOp3ld+h35P2JIw5rWVfwXh5eptEIPnHwF/zI
hboceX6epNk8W5veTsbUjl9Bl4FM5N7PsKOjzrwe4G7qSQxe9JWAIrgl7NFPFjws1gvNizIIRU3i
/6iNCZ1ttvU75V4v8i/kzy1fMPXHOq4EU0Up6dhl3BsjFsOBlidFLNxDWfZ5gTU1nJes85aAO0sm
VstIUkeedx0fjm6o7q7FkNpgkrtowqXvVY5LS9Z+ZD9hrKDFErng8OHveC/4yct7AG1cfeuURzpI
memALemGGJqeHjbXQiOoNRdtq9MIx0fDB5kkHpoiIR9Js+xFL9LrIiRE9ZYmrotBdy5Npoxps6Ms
3A2rIt4E2ZTJ02AhYKC2cY3wt3TDjr/MGa7+amgiMag1dIcfTF9N4LLTsnpuSZJJztiAUbNJ8a8i
xY8E2LST39NOxdYWRePis8e20xY3TWjLRk6QkluNwaS7vDolzn/P7mugBhtWWyxrH8APXMOxsNY0
Sj0y7EUi5mkLOI0zsWtjIFz1vZvPvcy+V8QixPLT93qwimz8PO5iPm56pz31UrVHxFYgH16K1lZz
pcZYa3dzaQb9nTtoCW63moPBoSOPM+aW7MM1UqIAuMJ3IqOBhVlw80duZB6zMQQek8YEBRvpllWg
4S/jSooSKev5y+OkucFZMB35y30sJMOaqEyDe0uCG0xnMZoQwuuTetDEpB7gPSmU1nM7Z24s2rpY
gvPPWqQdX/D0yAyHymMAApTy7dFQGVsXO1sNUJWWBwM+6119tcC+0qSF4ljIHD1hy/I7JI+ubmne
lB46KA2Hm+y27wBYrz4OygMSncvAGYYjL98NDWGY65H5XSPweJWWwhViHKwzQcTCgZEHAgVNxsPh
1dwRcr6cOcWkEvdaqaGz8BU6alS5QpLliUmtjL0cfBx0w9qPwWcxiwlOrP5XRG+FLMRibePXU7kG
/R6aBAQko6lJx4D1tIJiahHBrHcGW+yEt67YO413h8OXqO85SQtoNnlWlEyqFXhstilQh56hVRUZ
T1b5/3ldMKbA6xO8NWj/ntMetbeH1L+g5bVyMnZ6Frqf3RX04IJ+3y01SH4VfVBxorGW+cBAHdIS
/qbM1S4eZ7EHSmj2bi/mBKIzEstWpo+BdR04Se5CRp7L1r9+1wi3l/GYDWVYHml36Lp7hnmW/iy2
QwMPxRWB/I5mneQXLINPfLjW223PfmRmjMAaXYEi3UbWV3wc2fXA/q1tZgzQxL5MlnVkK+3rMq72
BA4tAJxUS0BfW1SwAMBf+iUQUHD3i59QHF/q7lBrlPzRgQfEhonSDM98anZ16BSnDnHAMIpVIV77
CZ01n6XhJqsYe8ivBMpin7/JDUFRv9GtOgivfmF7PS+I5oHjgVtLjQBwCA27CRSuttJiLEHQfu5f
65wKGUOnkBqi1wOvodmpFBuOgcR6Ho7GUDRt5fYAx8OMf+OoqEPAqLpiamlNiICMHgMXTdYcJZM6
f9l3okRdjg0s/0/NOAk55PDJqfPXA9nrwaiG+zO2uhyZBF26QPa5iTA4OcM3XG5Sawo9Z+OIYEib
/vvseOTjNOIpldvr8cOGiw/9v7MHVZGGPYGY+EAXCtEcL3OmzckfCIaczi741lvM95U1zCmpIVwK
8idIy1O1KliwYj+5u+o4wVHHNnwUKDeqLEkQyMN/Yx9WZjBZHGGMHJ5NyH25oEbxVe2AOIKnJlUl
axQPRdvtI7RqPDrsNq4aDZJoQYXAB25X11ZfzjWgTzUDbaOuz58ffUWk1DiFxZKIyBRN7O6/g0Yl
cns8WPMyfDZhpJcKqqLaq6isOBVGs0Uk72EdLSeyLX1xF7G9yxyHsB309SpIrdf3/Nr1H6TqIOyn
iZI9n12u9n9cwC6XyoaDTgFaoy+Ijbcwy3Kewo2HKCpQUKRntDhBykTwkuHjuHEf2lDlh3+DLf92
JNi9+qHWQ9Zjn+T9ivXqjFcMHebMU7Fb+G+tppJ1rzX4AjoRazsYuiwE10aytLkv3sB1EkcQFYBj
l44a8HNh+hVhY3urrO9DLBMZdszvGOoi3DeDK5CG/IiNpsKpzIq3Hq8JZhDs2HRne6l34PqNL4YX
Uke4F7Am6Ix6mkTENNxGaej8pwNF1a8XlbDUsr/MkW3SkvG6iN65qbhzQjWhyFuttjFNOl1ZUxfO
btshx9mZ80un4WUiU76zR7BB/JdaDNC1GihjHrsGETHGrFtvP5Av8JNsvlB9r2x5FmIU+GmXCbCE
IJXEzyaS42ec9ePqi4phbfsVjOCu1coIfdZi42zz4y3jtz1CIi9r1DqjD1uI6ejSeLJBXvTNow4D
yFGbgdXbCT7p0dpB8BstNXGynUrWBP9+PWRGbDQkFxvqc24waGWtmKpnY1Q3PvMBNEiHXhphL5LV
4yHrnmqUPnVynxusaDxsTLMu0NV66h48AEFwX3JnD0OcBvBP5+yP7zpt5Yn0vqytJhQYcWlyXKOM
EkkSTDdDI0qozg0HGu7350yNci13n9ASseoLDGf+KYe8BYhFaczVvzAEdJG/y5sUI0i7M4N+x6Cl
M+Bpd+4lU5/4xkyQb1oBcPjZZDU3GcDq+FVmnHtedCKG3o8X/uHKdxFECsD0UuioUoIhKosG/A9c
t+sWyKNnIatKpV3rMzbv6pCUq2ch65Wo0KieNrrpeLdiMO8OtOiwjti+uUQeVlGaR09VkAPFkRYK
eQiRzXE1U6XEqGKINhdNmFg/r38d0VSZdytAIZOENog0ivFQDt6QzQpcMuPKWSsp2nauyRWjnZIV
cOdGcPGAoDgJ+72rOPk3EdEPyDbwUmtG2J3uLvAAnx0hW0HgjRDVC2plq0mvOYzlRSB8TAEQ7N7Z
8GV4cA5MfH2D6A0ruBuSwzZ1Nw+/3fg/oFzTAbCnozI76yZyYnQqUK/WBrykNNOwFXSHQvMKrKEw
P1Kmfab+XKpcfbG3scLoCR5slbMRlWeE9z57tQ2rjEhQ0dVtsnU98uLZ0t2N7VybdC2mqxg/aAy0
0izS9+6cMQ5GJAC2L4zXGsftBSQVPWAdLusHzUxXvvN5flaA17LKBH4k0Geg3m/itSz4wyO+VGZO
QSoLz0VdHEjrjwxV35Ba3qQRIOv7QGibYXPQUKppiIJck3pj72h9+qkCWyj170rtOU3NOzyv9sXJ
Tc9kjaJruVBJPTyhZaCbucxD/5j86Tkbz6DpqGGJg4cl1sGNk3DFYFU6uIAh3kB3aAaIaoInlHOJ
ZYF5jrndmt+afznxj+73/asqTP24v2/btLGvvonbUXxZEVpGUPJVMDdmY14WdZ6cDVI23Kl2GFL6
EIVaMSxlyZ/x4YeG6IqqHLeYwc93d/vngbaAtS52jG88sN/ZCkPgP+xyjUHelbAkiGtpKbsjSaqj
To5CpKi8QQfanyfymkEW+TUCMiDXeQAeOp3MJvdxNPcr7uDRT25aL5NkwUqM4GnQr08O6AH5//BJ
SL2s9SkZwdK3tEi/khSgSQYd75GgtYWaLifryS7LeJkz5H+raWQJYQj6b5GidKdqul3QtgSowwb/
m7uBxO8eucFo8A+mXDxgEdINpN2geKT2hh34TJTnYZKYcVJpyU9+ggvu7z50D03SDob73MSz6qNT
sCi6lTaL7G9WmSEu4L/Cz8m/4G4Ij7g4mTz3DWkxt4z2SgOJlIqNDpE0BWxfkb6syTRlw7fxPbMA
tOygVhcudu6rzmAXyHAZny5ofvJ1CYyStUUIvh67qhaZt+hL4toLl3qWRdCOqDJ13ZJG+hHKmDh1
JC1kC+i9oK/gkx+q7OPABvfJTJ79yuz3diTrB8YIhdnROIifV2uCiAfeYcMt9iGiPlbn2xDQePcn
D1lHk7FemfVaePwnKpC1tXPUmXbJV8Fdb44NtiqZRGvTN4QJQ+avMwTwVWretVVjXdLpNE8QBqu4
g1LVZ4kvNn7o8REBM3OWF2/vZ7C1H8IOWm7Vnu7C+Lkfq1036Cor/lcpjg8o7GoWGep6CEi1tZq2
xMAiRJR8vqZs8gqUGcY0rW/Pc0/Rc2AGmVzFsljnMo1VngmfJGfR1XhjuONGUfXL9dy/bgFRXQHz
5semvNx5VIQ6sAIl0Wp85avnbLNV6sfa2gWXcumgkjQD3qIOFHYAwzCgg2njt2Al+WI1tpF3uc3t
i/Ws3KU8LWsfiur11OtNnzNeB9cH0iKKSrNh/cQ+BjSEg1nmQMPwJmKmQR8Eyr18gIznMdWugSui
8PEus+jzKWN1FQCCy6Ki1ppORVGa0LzcN0IQfKNJvdmAVsULUV/XOkYU2Tf/BrLB25l0O91DOm6u
wJwQLpO1GLpIp4tQz6Zr3vn1yUu6dyviuP/fLbIB7QbX20ijEcbZNp/xn1pRNfEC7jumPrCzEk//
QIYTj9l9rDar3Cr5XnS1+0u4xKt1vDXlgygMqBYnh1Tp7cup1pPtLizmgn0LUpytCgbRLo5yxmjY
EWUyx4pKbZCAJb/s9W+Wlo+CAainrcOvwF1jkpKbF+NMi9CV97c4+k8ndWnPgd5cvlDD74Zng+hb
nX9i97PuxPpYaezQ/fDMTZZyi/tPeTE1vUH7BCybG9mvnHHuz6xuJM0M+//FnJIufqfPNPhPKsFH
pu87HiAeOL5ZIgCcMqwJ7fsyCDaYXUdojFBWls45HcP5iC+/fNAdANtyIzrtavwoKw+qXNmAwLmj
5rYmRwXU+I/BmkMcHs6jIMmidvSjlZ4eR1VRjpKu89r4sLj7RW8NJ7roSPs3tm1J52owpiJkuJtb
sZOSG2Plk8QnmtFgft4R1PaIl6QciQRZAHYDCXLU1SmFEXNt74aY43aL2arm2AU32agRijvOr9tP
0ZQRXRHrEiCltsSG0C5Rq3OKJQVJrHjQy7g+C6u3vKoW8BwhnVzmBOL080Kwuucw2JTc1WS3jhGP
vj5fcQa3fqIjSe/lOF4vkOLNAu6syX90JLu2BCseXiJnQko4j7vy72eG81mBIlDIA2nFqBq8v5Bx
oWke9ZnlbXGwxpGXqy6Cl8kXPQnqEvg3+RgeYBy3WeP5xGQn7tJPhhy7RUvSUku92063BBo3pPHS
nODSS8pqMWMvoSEiANVUz+hy5KQ+z8XSnG8RzVxLbrgzNFmqxY08e0z4+BBxAgadctNRs26RyHsK
ssL+kO/zxexe6RwkJtO2kbxgvGw8zlQuTih8A4nn2WoFWypytTVONo0FlJdecdpJeaMpsUq2T9QB
bGIrieSJ5UW1xtTfgIpCraOCo6EgGXbxedeoJDLnNeZ1cxEXGtgB6rLCpJpqR0W8ijOE1BO0OjJd
PVUoPxyp0YF31K7ble+srOPQ/PpgftkIbGkFXTM93c1czW42m4zvEV3ho4bTzLzGUOVQXPLa/iKi
bjUstuFkavYop1WfwG0KJmwxuUVXkF4mhXgReh4Ub/jUQjr1TWWTt17KTSrGDaAJzlkkm4jAm/ao
lfCRXXukxwXMVUYB0usvNsxAP8Jf/sktAzZdubevTh/VDsgy481UhSabXHRMoVlL9tE/66c3UQNm
mVT2dL9PllT+/OddCYTtnjyMtfo2ORg3c9toJZ1tI/ov2grK4S2GWTJ5OXSJxn1lB5OswZgHjOea
ogUnDNnUrSQkgw20xxEO8fQ0IkNBKaRpMmR29zzLRLMn+gPS6rcZy096a6P5C04RzjnbnLrtVCWQ
YxYOwg/2jq4kmLnbFD3FMwGohHcXWrtYEo5MgM0SJqHZwl89sP44H9+fEuH9cJrHB2sQC6RaPPKu
ta3ZeMdh5VrzSqqACtoBJm12b18+PJHXkal3beqFQtlVGFCPaRlGDwvn117Nc/UrHGK20AIjT1+t
BDLl8ich3Nj8MrqxEv6P52vSZqSBbU0Du2JZS98BbbK4stVsKZkkVn0dM6+mztl5kW0mabcoWFt3
IC3slEcsBxL4qbpJZmFjujXn6aeCgletpAxoZhThDBtqHTuNJSdAhn2sLTcayMqoy4dwap4YcFUT
cLHZP5PfoEyozQHnT95Y3jezdfKDp81xULHnnOwQPez9eE/sjLjGJV8dRzmLPDCT0a/B6hhtjLS9
rAdKrjj3BI5ZsYolXNdTIe7HHYGMkTMRjBlSNbyLKzskVMAT0/g3q9nXtwWUNiFPpFLY8Bm/t+2m
vD67fqmyzUytIDs3PrZMz1Z5sSDjTkV6A40iPrOhuvRBonOZVAe1laAxEM2ZZZQ53IH5D/+bBc7f
occkZLnsiaqC2UJc5e3fuwUUKwxu1j7OTmXs8kM1Yych3P5PLuvj158uVHh9zenbIgnOu+Pr4tz6
0y7Eo2jMpK7YY72Xx7YKJ/94oSNvzbIctlBvpFbubTW4b8IsfHDhuNaK19hI2Ef7i1RXl63mNX44
XeTu1PQdja/JniUdcfM4Togf27K1TTuMD8/4VIUSPjQBKgzgpTgx7rmJln+5Fv10QgVidw2W+eCv
k6P8q6WiHh+jnzY9mJCEJO6qWWMFIXFn+xois6+sQCrwKPh9GHOxPRK457Vk9mEm/gY89PKf3wMv
ySalrwSgI6JCybB9MZA9Rs7yKwy4xJEd/h+LaCmUoppaBB8DA3khi5HF0gsQGHNsXugSgbk48k6A
ifMW2Frqc2H4QE4KJ1oa2w0qGeqI1OjA6wfh91ofee6DCp1LHMpISEjJw1/fJfwRxLAh36Che15k
/f43FAyaO3zkJJYS6dLIBwgprT8b22VYkUDUJBe6RWwz+wggDWfMGjpeqf1fL0QyJcLA5A0O5ws1
MXitkKPY0k4lXqXwz8+jC630DOoxepU0BzRzuHJSFtsLboKa4xvg+aW+uXkiuSjfHEhVd28BoEXx
oyf+7fF5bgdX8vW2yempUV7aPcbdgY/w0/onQo9BwozuqmFCWkECb2KttAv+Fe9EWV1thBt6LrAt
+RsifE8RgvOAelgkbjfBi1mbSQbOzfq7S/T9xSErPIU7gTrVh9wR0zC2Ut0kNZHdTGkGufmOIOxc
lAgp0cG5yoASJO82cdmrDdhXnSS5TyzoLVOV4rrppmarehtwEJmzNR57ooXt4U6SK8m2CSEQ9yZk
WFfds67vFjgvr3HZX5u3R5AwZnUCpNXUQcSCUbdLVqlP1O+8f206fvwDPpiVnTmG05D1VO2eIirh
tqzokBR50OIjYy+1JHByh0ed62Gj5C/57ylLxhorKnYLckdZrjqLzwMRN/EDrVQdDibEzb+KJoPE
8C/tTL3TNDUJVITevxOqKarKkCkVkET6eIkUZGKvAASaX9JMBap7y8961jdZUoFrvI7HoLPX4XTZ
jmJ0mlTRTnQDUCJVVbwd4SWhYgVfM+7dqhdISjLY1EogO4nrwDnqWFM2x+fjio0bOeBBiDWDL1Qx
fcsKPTn4pZ9eC8p6Sxyo4Nu5ratNjNpqmiV4ksbTXgqI7Ri2ChFobySgjvSgO0r2wi5BkzCK7oc4
DS0WHCVHml3dUs6Bk//MUmlNFQMay3xv09bPYDervTFOStMLJSiGkcSSwRo5uZALkSEb+IRY0RTi
8pK7WrYFA7xdau/OFNBURSJtov1oYK4yKeZEmQbM8/kcwoury6h7dP20lZPhe8zldN1uziNkg614
b/U4V5kzmF9mS4L7RHAvg/pSRZ/HrvHpr7ed1q/X0ms01YjokOjbnNhFURPs7jHzrF+YoCh94GhR
T19L/ApLd6vhO91YoCG8n4dhZKSaPHj+y2W/N6Hd3JxAJmGi/1tjXEuoV3jSGONgr264o3U7aXuU
YYhvd5+tbZ0KF/SDlOFld/SWfmIzukjvCOzxhoDXSNh1aLgUC0+mjmJqahzY8xki0BlNKdxcGuMk
OaioeCee4ape9kkcLwTPw63TUTwlxixWSLJIa2xOol8id8fkTQ4yX399URvwSqf+Db1yMU00+yyo
6VAMHoewhyueweZSX5lpKtFRphNz5n/b+H8a24JuPK5jnCzQrPS7ebNz2Ov3UunY8dLbLZ66+//2
1jSiauz4H7o6W9Is7mUYLtNy3kW7twR0ahh9FbA7J62TTMsBs707gGmcDW6ZCNHrH3L/RTn3Lcyb
UeWvMPZerd6/FVwk+yqy4VQQFLnRyp4HtD2cvAUprhFpuL/Qr1INzPEB40uit0LWSHCG2xtaCIhG
jdHsGSqiycktq2w8iC+1rCcVKON4W2BF+wCEnJ7MAVVBkLiiuJ/zcTutuE6i9V11dS/lJhN6mCLj
MYbU1ynK48pJzPWJeLMjfSVjCcsY9IBtZoe61Z6CQO00k4nqukH+WqrNU2vDE+Z1iKWACQ+p+QL8
41gO9RVt09T3xojfw6X5suvxcoLQewUjWKo+QW6zlYo3M74qT1yssu9tcs+hOEZx+CPGYy34Io1R
HoQJbCTmKFKYOYnkguLyNRxfVhi2205sZf+W76hjlR+lMz73mYVh2fIxMX7qeLqQUKSe9lgqzfiY
tlDfewslgLhrJxk6FR1kcdXvZXgYehZtvkdPCYSLU+IgDzPztFK9KesXzqezqsPQMGLksNkoCWVh
agqWJz6stnYsXYJcS3/HFwbNHHUGqeISoktaHvjH+5gy+tgyEDeA4G7mzxsTMteO+sT37nEzlXAv
YKUe43h09gripSbXImPqlcF2Ltj3WQbc+0ztiCdwdm4LfeW1+7cRGpt/yjcXCe04lQdK5dYYnFty
mjM5MJjDs6xhC3K1AKQEK/j8UIRKx02ooONKPKGe6LQowD1WGZq2qjRFaNQbzg9zsFVyno8fgpOs
xVhqq9iOnL+TjEB4cj8NwN6eVPiERqBLi53P6dxvIZ4dcFdVs/WtlNRqmYotLTWYd4loWYEjnU35
bAQJuJXygPARuiyOGJ+woap/979MF2ErHdldiqGtWISrtgfFR3toSR3VDymvTVCzar8IWAVv602W
qkUMHOJN7Wh3Z1wiiTiv3rzp2HJCBOqilWtZNu0EU6qc7iZlxijfmv4nN0zR7BCt8cBXPFUebGCo
rf/ThS68bZmFkFNV3bLnh0AaRTz8r6oray2m7ELEiYPa9ZT/lsGQy3CBz7zAfRJZSSSfAb5L+gGX
cBPKL4SPR2MEoswRmE8qJzqWJtYPRcuKKeMv5Pu2u1Qmm1f1hzclwDeocoB1hBIU/57cShE4+cuU
fPaYeVKUh9q3X1ZrtzMx2MsWSbFJ6xd01GSw2iiwx6YQDoZJDFCmtNJ8V7wpCmfp/lEPHdq1kLVS
XeazbVeUfvRznzJOAcnu2BHD25lkT0f+E3a1gFJLXGo9EZqqciQdtcT/Ir4JdE6Sdo7haLVwjSBI
hNCo1hRQLzFIM0u2SKw3mxn03I/gQEkNmU4z0mZYHxONXZTet7AoS5UncFawppYAMoShV9kY0l6M
beibsiqORLbsDVB02joM8cFbjZNzpk0Qav3Qb7oY7K4sBvvV1vbY1SIlUt8N/X5bE+95W4tnQUyu
sLUkumdlSiaHgnny/w93TtyoZLq39z6ZQb5+ciDE/5lE3x0OAVZKC4oSixJZIBErf+qcB72dCryR
2oC7wYP9SvIEOmdG/snnD9Lcib+1H82WAGl0pz0jRAcowzq5jnkc8MACVdKC14NEIXX2APeSyOnv
HKeySMK7MITYQhHWOX1ggj/xJ+Ao1X8xVgD+wRjKzF6s4dM4Rv9aT5ITtekIpnZiOdP3OQauKtAM
7+PR1yjtG04Jy3pmrzoa2KDjTwfv5ObnToyEAXrvKsEDk0tNhKAvOxS/TtCcRhZ7NaMb2ZFDIy4C
+0AiKNsf5Cmj4IC1C+PLDFnBTRKRfEF+ydWcrwWsG5hGbnVqrUVDSt3M5JlViHJJk9B7VWNXcRIk
xDcPbN6znlQgBW1CzX/6PrtSh7156SJitM0bw3RJMaSIF19n5FfDGCE1We1lY+XtrDJbQQXwJUSy
xEfZ4NvEyVTCEcnReMsNM+kIR1bI7XojUvoNxuKiLx/fok7ND8e13CVgX7KoqNlbze7ueB8lX8GE
pk35HIKht2BS0S6k1cL4GZLGuYP2oYyKaREGF3TPJ61W71R9JuyLy9xWLMlUt2wp1dDn5B3Bz0Fi
u7cLuAuPq9Ro7BShETJAdN++5ygafAoq8QfzCiMZx+sqroLF5q7IHtp0wMfRwRnEAA9h1Hx22pp6
OEcaMqU5YBgVe4NwUu9SgnpnNUcVp4iVS+qYTJMBn9FHRvHMVvrDEB9rkWg/0dIEfAuQRuRuGG4H
DQ5n9hjB3LS79yfmlc8kShW7krEpldNUq/45Ic9p+SggHrJEbq4oZn0YXeHPE+rRpXgpCRUpAVsq
2TprFutQxfS7b9Z2BDsEnR/hGy4Ogzi+j9iOKlIdGK94v1zoeWyRiACH0Exyzerydh/10M8hM/OZ
/lmpW/pMJ1IucEOf6dnEerLMwVn4zpFzHIn4GVruEr7DH3VNzQHLwKUe77CofnqeWANey85R3ClR
xrf4U/A3HCJhLQE1PgPDuE127KXy4nD35dJAbGej7rnWiXCfQFwxynqsIiwng2PdaGHWIubhKlNN
6gTpU0mubxtUGVi42Goe89md1hZayoxnv+iflsHz38i7ipzp8ORR18F6eegPieRkVVuU6ufvhXls
F2Tk+f4W8jF2sEH9Rm47Xg1k9N3vuv86LPWzYuljjuoPHIZ+U+by7h8Mb7MGyylQI3fxtdjXrDBr
V8qIgxEtlrZnd4PYojHnGZwL4BfQKw6YhNXAdt6qcXXzdQeleUuYVhkGd2WFKqDELyBOEa7q7R3h
e018qc3GG+pxdVBbXihORK3jJ19UuwVBc3n2H3pBimFa56DuK379JzUmTd/5PzogYOpt6uVc2P22
ByIToXU+rF9AJrQtP3I2pOpKQQ3/aL+E2K3K1/J1gu/7ltyidWnirhTkuv7ddlCaGxQ3Kiup8MeU
SJ/VVncazxougut/TEO3a9MEcmwNFKupPdwJHqBO2JLpwyu4WuwQpD6PS+lBFoqjhDgejsqAJpVy
PCzwBz/K26ikFewlwRHOm5Gb4YfnYpfoxbHzZG8OZcIcjEXuXST/xKuonDzV36dPuZi3r/uMyJOr
dnzE2QKKZjs8e5Ph1maOQ25nhMyXqzDEOYUESJmaD9QNonF6EuG4FwG0MQVdCgm8XNVTm2V6Ffuk
CmGdrtpcO3wkjYXQJvB/v/iZmzhB/pc11U9uOKRMjv+R33LQJMkaQuFac6tXjXifjQ05e1LgmLLW
ADFg0TnEYYgH1g/taiqrIyS+7JCzR6i0A6LN/63tjoSjuhOkjhBr58rbFwnknnxgGYExZrsb8+Xb
3u6Kk2/wvMGfID2sJ9PC3I+Npslqhyw/YopWP/F2PARCezr6pXNUt3FwC0cPgaYmjEk1XUIYwXzb
+PPU5ofGBtZjtHsfMypVpqcOo8Q6woM5tM+9uKY/RM6EE0twJ4hjL2YjRcTiv++SDQiQfWw2jupc
Fj/ysgWdc8bUu4yOFmPXBjCDSPZ2P6Bvi5/qVSQCE1QIhUNM+NxfCq2rRLpcfGsYD+huvZhXf5RA
XucFQwRJ8diUefCOXPWViZ5L/d44asxGGYryV8lQ6TTK81rjA/ntjcuY24lZCe2+BGoukL+S4tbD
aQfwyxVEuF96lW3VygAuLIpAAtNTihCPTHRMJysIdCM0Ug3zF7xQq99rhM+pw20KFSmm53oYAVZV
Sw6Ma8KuhPEEX5SMosNYsf1nhE4iq08xoGKo/Io6rrfoRc0RZdwtLFD6L8dm9EVyt+2IYiTz/dnB
Nczw60LlDjS/9HqbAEmxEvItBSYKJHNJMFK5Pic1TLmo3RXaB+XF9KfQRd336m2Y8nfxmGdFnFiH
LrcRxOew/2Vmxl8BTdD6GzxHy5PwC0m9uZ0MR1rfr3DzlTfJtFumVXMKJa9b1F8ZsYEbJIdvWd/w
1CN2sfvjpeAnRoRa2PVtS38wB9jqdhD0McATk/CK7lC2Dp+y8dsB8bAZm2wlM2o8t7zAzKauZRJ+
J1TcQYVT8AojMIFRcxIEu0hwiQurKQO5hj9kYB8XdV5Zn6r3R2D88zyGmZXunr7Zei02CufrS1IG
9YkYoN4s6NcfROtGocp5dISCrwJBctZjvFYJPUNtUQSCR6b93mSto+2kdn7kthYcCiiASNqlLtwZ
KPBwdLVNt9DDFMi1YEtzS/9fC5pZX7Qs0l0MWAWe3JftNq5NBIV68KKHTGbsZaASAhOztdjJqfme
sjTFUMv6v6Wj1CPfD3CdDwNmY662lfBHeVeiXl4GQp6qi+HfMuDXm0+nZ/rNK6VUrsH1qbrWM4i5
I7aJO9ypXs5X7gXZsrCrCjG7JT3LpGzNeYmAggky6NpCM5e45doe0MudZvlivzUYuhEWY1HCH3GH
sspFB2A+7pFEGqdgHqXP68hyXSOMItXGGB6CPc9FxelFXNu1VZhjOKOGQH+KmL9+tw86e2VAC0Gl
O5D6n+BMoolcsAJThxHxX5zh9JlwSSV2XOURZV/lf29LyeM+CvEZ1ikIVBxz3eE7sKKejMUP+F03
TrOhJj1KKSgiHeCP4HAdGtJdY0Ujy1kZt4yTA4lfU1S2lKY+4PQIsgVgKhNop935tC29r09w/Hq4
4YVoWLSw0wns3M2WJVi+DC+yPMbTY2diF0ZaZOb+qB01J/lnFHLPH7rL/xk1AmiYFBJcBh+gp8nn
ZGx1zt/+gIsF6/uvEl5+ax65UJw4Y6D8dcsDt5CPHfSAw3B/3NRNoYnOy5SceRY9EoIhXLkogsZu
gkNmgixFm/Cynvh7DK9Ff8rdzqvovIQJbf7j7iTH4Mu5gA4BJztYstLW2/xMCoLbTMWJ+Ao8g9p9
YDhF0T07dl+F3EpAPRxuiQ28IC1jlMuLDKe/yNmYtXnG28ipIivfSUNomHlkPgi9FWO3u4lF6IXN
HwAX3WTwSx1E8hAOJA1fu8V8O8YwDkoc7hHFFjtz6JLPgt8lUXbiMgEc2gYjtA49ILFS+0v9zibz
UBzAEphOQ3rJCUbzVGuX7ClHsymYVf3tkkygq3QmdXB3F3sv0krEtMxmX2hxU2D0hHlDnioFzOsm
LmH36VmNTs/+9hy4zyn6GFQh/q8FiSRziWh7xCr5Z63z4Scb89iQJJUvPCwtFSZfG5Nd9Vzh5PMu
KVYSzqqBEzSOl4qE/q1GIwGWGyLniDEGg//48DdLaAYklhFrs7us+VJP3fF++zrzXcL9d/J8f1zU
hm/LARMV1rzTdmMYnzXRTT2zTEDddgASRa1Vs6u0DWQ5vErtbbABr9P5+wSgAzLcbL67kPFUWnrc
ocUAdda8levV/FV9PJpESdTHVytQ2Nz32Mma8362cwjfEUkGUVG+GNrgO812pDWuI01m/VCZ+Gyp
FkxTuxXJhVDJhJiq5C/t9MncLSx3wbi9cpbosWAocHPtWwyb+QEQbRB/I2Vu1VqHlfe8dP4L4JGO
ehV9MOkg8GXCQz3n2vBbh+W9vj9Mgjkwc2BZjoBFkwYHsuPOHb1pYa+2o0xao+hjRoygezi5H7rg
oAxHZCpEs2o20xPNNUivT2vQ0TUC5foh8pC5lQQebu6caj+x1a9+hyFut6k7q80llLrgXN5oNiak
Mg1+BUkItgY4wtvYdHiLiAqa71aqMcNbeXTzrHpKtHM+ygasmBNNbpSEbUf4JwTz0HrxMhZnMM9k
3F9X+RGi6X1iYK4M5d5mYdsdZmp6iithhZtLPMv2ur8zaY8/rihUI9pvebz8a2SklwbVOoK3n2kC
Kew2WUWR047iFnikl2nwCX5KVX4mdxh4l52rUkkTqUqF4CF9NWq4XG8XyYswDFrMqNvs8fODLPEI
UHAIGR0TlXO/NbHUDZzDkFOF6fUKrDOReLgbhFudId+lJ/v0+p53lBR3FPniI7k5JbH4Eu3FGuyQ
vg3pg9QuBJ9/l7Gk8Qp5eo58VQ0EpT3T0Ov6ipZVuZjLpOJn/BMLC7Asw5svTDc4TSC1WCEnRZtV
fCHiYvzRAC1x+RrceIJApdy3GzC2mNpLZoMPe9kOQXz/UguoeViqxD+fXG+JhCr1RWgUCjlM3OQL
ngTluXAiw2w1/fabbLfm6rxqOMFxAjreJWCwO3KgxIYVIqSoBeIZX6JGKQ/JfBlxiCk4zXIIv4Kg
/1te8dezDyaVvjZ/w1hBdTp4Itm1Hri6UPtgQuziSLcO22woJyqfloq5i5Yxpe5Gg5eWjmeIvU4C
JvDEIKKS+YMqSDsPzothD5faGr5hqCloLxuI7xEUiWcAnQOGSxIWfZhZIMeO7icIr9YGIzm1RGK/
seBG6ou8zjslNQGmHQcf5JWNr55ytf+mZeAi7EAfLLN1t4a+lY+SmPcBzor9t1nX24kbcduXgTsz
03EbGr+KIW2HwWpc9VvONKtUOoPMTRr52L75L/mAIdCfIHWTebgwajW0xvLkN5i6TmGN6TiDE1fV
4uLznmz/vu31upW0bDkcXC84i+zn7XpUQJAThXEFaOrrprGUdNXMPJsmt3wCwcNJQoQXT5ZMoA/Z
vCnz2K+MzXdnjfcGhy5nUZQ8M83bWreecCVIFxkNsqCmAyu/aHEvHy+miOQhEPvMumxmYAdRfM7M
6JZYeFydtOWGHybkaXgZlpZxVB6C8/VyMDn4Bp7lWJhD/WmmIE7fLkwmbMaEOjAXJ8KmylXVbw8X
u8l4LitBo+P6vi48B2r/Mf+Yd9k+PtYFU0FmGb9qK4RCQeHht+aKBZpIEpWUbpXSDF6ahYlNxx8J
d6wx2cqdmLdFUFcFk1sinqHlGqKpkT6pBsQ0EWF0ojyo1zhFPp2nKgnKayz1hJP8VfCNlGpqqZuJ
rDVkTiJqtXG247mnLhEjZqPUcIe1Blnqd/Yo1EtpR1PI74W4iLGZUMlaXiG3xeh1ontSGmswwFZh
Ae6hvnj5FQER2xTwXbbVWFVO1x4xcD3GLXyS176Uk//QeFR/vlVUVYdcIFpFG9baVt5ek8TFdNOU
ZCVV/vtbVKVMFQSh97wfJL01y24y/YsPeFLPDSPujQ3/gmiuTXBJ7kXGonhYROtEMj6T/onu4Z3S
gihDITIPdZqAhnmiQGQnLn3A8XBeqivdcVLSlyQEFYy6m5P4GEktZUfqgJw8pFVKBxJtdhHoySEQ
MyALoQikuQqIIRdHZPn5pYwOuxXNovvKeZxqL1FB6St6bgu9vXUKI4E5j5BYzzpUkM48Ng+ikOcU
MxVHQFaTONP1r4WnC6Q96pAGH8c2FqmY/uJ5ajP2zYHfCOF/S0ruwWO5/W27FUJL2ApIQ0AaQMyt
CroErl4r8nlLsw4RUrus347UZcuYL0PsDGQrXDGzT4aQU1nE4LK3t7CnualpKUgUm9Jp2KguDa+d
NEucC4OB22aWTa0tGFEFqTHSxjsVHu5UX/HCdcTxk+RnclYmWqnDOqS6BbTf9B4uTVpMEITHuScS
j/RAJqpUxOKqoOBViFDFZdXnV5oKLSzbHN4K4OYw4RsUg/mOVPmsopFy0oHfkvuRA0rcIR/FkkpU
vvvc87opUvVJ5pGC04DkReieYWLVX/PzmeaWEv+36MIM+UKM4i3kZtkETKWJunJZD/q7PtttxDGM
yqPU7P7sqz2wgixGgYKxL2VC3hVbwH04gu/u1deKwDNn2YfgNf/DzYoF5j7VKGETCdtNf/AF/BTj
EVk/3nF8EghRGX50TQZTiQ7GmKXj+RujgkHqy8aq+PXmmyTNgMgboSp1oU6jA6G2SlhNJIoN1KhE
l6IiZttgYl//82+BdFuvLptkLkX+gWeQehQeNS4n/pOI+3PU5fhQ2S/gyRa4PL1Pi9+eec2c0nhN
Q73JUhR5uUpTJ8bI5SH+fRhFQcvxCocyzPM5ef2ILGTqSqNPVbMMLEaZOY1Nd11cdcxb91yueYBB
nLvccGFevRi8LWjFnhagXgFMKkbzTytDQwTg/PWWCWF8AlZyB5Bs2ZjGo2d+da+YPC/1jJMyV+SY
orBdQqJfF6PTRxwoMT3FzY5ASM/MA1qNBAc6bwnKx7oUSo5hdJhs6GxDxUQgPZwUG3gbSRtMpVrZ
0LEMWIP9zpM3N8CB41ZRVUa3yFPuGwLzGiP3FIjbaMFxV51BkCKLL6J+d05nyOoO9m8EgyxCZW7A
vi13N933blJd+e6+ujvSMKwR53gDVmlFavfA0SJyYsyMyD6KLJUupanSt1lk3V2bVsulbe8pBva+
ZJoF+lWiZIDeQod1ueAh37+4CQbepG4BnHbdYK6BILCEfhLEXjTBkauP6GN9oURgARamzksh5JqD
VJEdpCgMvt/uD70dwrhX2zDoRggcx/k4S4McHigZdDyeCa/8pUIw9ZOKpF0Idycf8DuHwq9FlA/N
edkxNeO3zr6NiKvy/oSBNcb7DTdru0NbDNufAYG8O6p0WPhsXMC68oCaZxYY10F7b0/++e5KFi29
OswIBrdQumxsuSsTEnxIP9CBldDHv0iRNTb/6wEGQFNYaRCTKQCh1k0nRLlKff8dm/7S7/F+N3Mf
OVmD4pWbB/vFkQSbE8RCl15qYAEC8I4qZFxxCHWjx/3GFC1Vfiocud5uu9aQcDMRwxipPIR0Gbws
eQ+ZHV1cJ5Wv8lD1wawsmU4W7vO1mKoRNOwvH9dnrK8G77HOfYcz6oN1jrgphQHNbw7gp08ecYlR
F/EWP/H56IvXExWV/0Jr+tDzvivKAlL+a348GaZ30kGsKXiKVPftSwfmAs9V/cRavdaOAndZTeZX
oWnNQQbz/LdaxTYc6OzH4R/FfnCMwXtSR3KxPIUedzArexq8q6GxvpZkECl2+N8I0cE9JnNMAwPW
WRNrEQqrpUsoiF9G81A9QhYc31PwLjCtrYz9yhmMD0q21jLqK9pATLH9MN+VuBick2iocF3uQc69
fFudYAdoPLodib6qbTkRwhM8b61EPSFSJtzHpbFrHymwXIH3hgHtVwZ476RFzNLs+FP3cgK916PD
KX/CzMh1zACK6yN8m/nl0JhWhZA1dGNQMj40+IlPDvWQhJTGJjd8LnX4t1RPRXvo4NjxGMkrPOPt
IavYjRBRCUakTNeXuMby71A84FEJrzLdnFY5bqVBSYUaCpGZu+XAQB3j1UNOEZhBBmZo+nVsKVdH
Hn5afafobgScyaOvHlM8zvkuhwf+qwPD55+eKpteFRPTkT/ZQyg1gJgoNTdHYvGDx5i6f2mu2Hm8
+4xJog06kqyv2ILRzQLFOwkOU54PwvTQge8kO3mqWlLqUH+4ueaPLdgexTt+7Vg/PfpwFuxP/Od2
BacIHB6DEXfd+oXFia/hgEETvncYb/F1lsUKJoACAUGN+IeK6v2sW4jXRn1gXQc2cMgt3zKFjKjn
7gTnIQN3iRJvP5ezU6bmyreMG/w2uY+Vvd3kwaYorCe9+3EYTnaHSW+XZuEDUPCCRv0rQ1wldi5G
QDO+vzlyIoX8ARPbhCyK54l3U+62jiAZm+OHiKpuGbnM+FEN6pCpaXxDNC5eZhppr2YYNCDPJc9J
WVudZIi7iyXkSMz+TsHuh5FpDn8EVZGVgUWHupT7v5DNPp07IajMyXNmnqaWAgjWcZ/ebKiSLfK3
e9MNeu3jNROnRG9+X8Mjl6lwOtTTPo7wnor7k9+ZnGvA0+t5gFl5/gCzyjV5CEFl7+VehyvAYiop
jJefHZSXBEY5Dfj5+7Kau4Twy2MHhSwq9EUFFruFlfnUPd35ySfZoGoUckgBFhjZgea9RDze+oQr
fWATrSOgxZ+RnSFYyUku9CaOw5rMCUURyjmQdUYxzYtnBSFg2+ItOiCZSgJPx8ebmFIS3rTKhCKz
YcOzLxWCkdNLjHguAZllBWkKHZkIMHmWN8HKHxP0MTBdtgagqhctEK7CFx/rpB5cZVBOqAccSUUc
hnleb1KIJAcNrjvWrOxqFdpcK53qXmEKfkftLyzdeNKbfhUN4SQmReA/QGaXAde3vPqf2dDoh36o
D000PXuMk8Ry14eADdjQUGsT2X67RQgj9r7+PXE6V42WcwJJk2wJeaELdl9iV6sg20Krd9/+LwAu
8MMtluPYeSdBMkEgrapQtV1GVIzPBtxqjH3pzfnjKgB8Psa65C517QBNIaZ76oM+I6oGdC+xp/Oc
VzMJCQXQb1jUjR0KQ6gc2U87h6pwBh24HZ7wujYO+FBnE0KK+G7XPeYXew0basw888uma45G5ibQ
Zc9HZsv1hepYQGGSvc7h2LcxcLuwe0A3Kfqi7VA+cMWdpSWpOVMoL5D/ZHm2dhPWG3/K0sFqhphK
2op7tYBNLbR/NILiX8u+gJYmSE4PQAsko1Q7vVeuUYcIBx8GjSPlKUKGRCEZKq+jp9SUdgUlUpjs
ckiVqpg2JRjlo5ANDWSRA/4MxCTkPI3sH5eT7VIHQMczs2XHdYkcft3OdIOkW+4RkntchB1o5ZaN
NsNYamjeCOLC+YDLrSrLGdVbHRTI5h7rWM434IluTXgG2dMwCQou1vo1HyZSW32q7DzEeMP+ZAtk
32RIk7zRMVVQAyUb8n2nm6SvIkDfS02qZFbmIL/6v3wnSBIslU24HjNp9ONyCEndskeNzUfht5Y7
IFb1r1HqGR6Z4jHvnB9LBbpPKzXE9EiCz4GhsA5ZYHcyljFMkbB+CDFHNA3doAbQdD/hK+OM39Uj
YSu4xmBHhPrCJPVTSPefod3C1wRXiIA1MZkBzIBD2ZBIx7pqi0YWyE0gbzsB1mgYPiW8F80RtGaz
uAFDtXrbqRdxCqdm/L/XN3etZU6RActdeEj1ZuiPtM0s5PurNRQUsATVyxiXcH5WxeCPElvjHRpl
M1ZXRknrK9HYycyer6L4utdH+NLxEqIhI5QqEIJS2eZ0t+JABHEghX9+aWCQRkoOmAN1pRlbU4f8
DJdZLmkVU65Os95XZpXV2tGKMSpoQmyCFHYgR98NOpegBYxpnUOmOb2/jwonINR4RGezu9LpNPt9
5mB/0hAoM9lQUdtsEfQcCtZcHH1CBOI1MltHOe8wpx1LBvATkzSuemjulHgkggsuERf8GGCY8Kp0
Rkzi/fVHi94/FizuFzIE7x/kXbtK/VZcobFY9z+5cO0MZCALLH7OTrAf4fOyk82bLT7OniINVgCT
ufvlOjizgcLvc7QO9DT/8GRKC6Cq6iYrKmkVFLr2ZwVQuwv8vguMBd61BeDSQyC6Jt9ofJO559Gu
A9/CAvi8fQSv/OkYjkrWCt290bGmzDzZ4qo1e+7oQ08BghuD1XDoFm4Tj6EHs3UVeoN9Kokckv83
DNdubIy9VjXjpJanQhMd4pxaGhMEE0ttNsMoh3b3jngUGYFhEUVc7VWgNYo1mBh0RvTLDKiyNvDl
O63PL7HLtlhs9sXRbN1MshbSP08l3IsQXm+wewg9nKM01elN4w3/hYC83l2jeqFmP59U7gS6Jhwy
j6zpPNKiSamzppemUTQGCe5wT2Ogpo9LlYSmcMlkhNCVQpT+IfQftDgCAcgOK7gVseZZOtklCRw9
909DPRsC0rGQYTTr0DNVKOYTM66rNK3UsIuRmFtxH8EvwWZZcfj1PPLyt8TpAyF3i98cAxezEAnq
ZrmMrxiSkEcj1VEsFSyuhVdYroXwIDSpfIOgECA+Grzraa64QqLxtxcpzfwrzBc+b4BqCDpEot3T
XY7x+1/vzZnvRV0nZ2d3hWjzNyk+zIktGrKXbOlZtPIhAeJ7ZP381nhiZFBk41mokCs4awI8fFtO
6aZ+CIsoaOzRV/KQqL+Amo1G1dMY5uJ2S6gBS3eGIDeQSislAsr9PGgzciJj5BuSzWtBhrqPSRSe
PQUShuJ1Javbq9BoiU3It4CIAQnhvcjo+rILHRQNYBodI0dYELTAI6e/aRCodzUWqYxBq9lR/KoN
IGjX7X03mLE33Zy3Dz+miZc8X5LIG4Lh9H/5Il56FLgvuPWISW+z0k6jpT76+MW/m+YB8z4Sw9G1
nxOODmq0BPI/b8CtIhdLZwUEIzO3qxgkHwdhFS+o67ox17X1kn+DGNRQmsQ/xWDAJ/fdWo7VZcI0
5oai+4V2qtHH60VtBQUKMCOmCMZ+xUgc/oPwblbrdxQ7vTGhukxd+5Jly9VTco/2ZXFRQELvL3FX
M5b4rRJozSxIRpWnWu9KKhZVm2Vl5/GsW295DykXiVfIFqHNq3ljul4wxNK6NUE7EgvoEB722GEC
PXpVGCreAYurHzaF1bMJlIXQXVPxSYY7+C6WVl1CBb9aHt3OEsv3as4cDQfz/FIrg6IncKK3MHpA
TaUDIM9pCA0rA0ykUUDOKtYGNDacgcs4tYCLu/ZbU1s6JMb/k6e/nzP8/GmHK3l2xmR9xGZQ7Ekk
SiypHHTwpsnTDxI5YuKzzowcSqoYexWSkKcHR3sUuhvuNRmSaM3eM2mANFF9syBVHfmvhUjXg5rj
RXMrHO2BWqb8eQpDV0Di+nQDo7bwpykZJQ+oj6TD3iqNsh+VphQ2lWUJ6Vhs/FPl/EYRaMg9DcpA
clcRclD6QP99SbT3AYgS8Fd3Bjl7LgSmdDIw3wE4kwJVT2lySbAixnSm2dMc9hIyNs7tZYEinzV8
CM3bnThdN+h97W9U+D1YP6v50HMgINBNLRHKLYX36NWP+EywM3Pmmq/ma8ET2ZM7pBa4SeiohEIE
WI0NW4FUDgCv97FYenDnTQmtPX96mS+8qHaAmxB4fS0mgj8An9GkmUcy09KgZD3Lc9PnNMRK4Tqp
UZvzliQtkswcgorkXaEPeuuhqQ5qEc+b75sK1Y6ACQhLiXEhlA7IwKUC0WgsnX9ZdKiRJW1zjqLD
yr7BHfWk5UP6qyUon56wRKSAfE8rVn9euvyIwE+8POlN7La4UONw1RzLCQbfuT1NmSge+gP2M778
BbkQS+Cr/AAQubVLT14RU/bNwVlX7+yvVe5e4BgobqAPgx8h8UnSMz74ZR3XCqeqc0qMq8UdULnh
bFlsio62CyyxsCqbybmUet30scUaRroZq3Z2+ZleUAfN5/+smTEZly57d4TI+EskMAsuaqJUk0vB
udV5QTeATP8N7kh8iy/2q9QMEg3G4Xd2EM1sCX/uNjuwsg+5fBqXnedv3Lpi2pGfekaOHzI14glh
206eYxCfZ0hgRem5HhIVN7HQinVLAyUcWxZ+QcupfhgQe/U1k7INyaa5x6gv7MeDyuN5CzrAJiur
4cyYIXRux755LqpvfgvkVma5lRcERXp9Xmi820J52qKrC672aukPfXD3oE3RzmX1cFMe/RrVXgoM
UQQByss50bZdwm1EjrPdiQfPK/sf1dSodoqGsWMJNEyTw8xZ3kz+U2Cs6MJt+EqjWxeMGFnEzoDc
FF3JkWPKnfOOLeP/JJaC0srLJ7idZwcJW4ZuqlpRcPh04nDZbsxhFQyDZGFh4/R54C20y+aG009h
fH3aJnTRkUFjEPHwwy5WeDXtTrZEvXzDx2Cvjz8Wd+nXEODQkK7z+6iQUKKoVPrAWwKahr2d/iXE
YNK60uupRcYK0XIRg7BeJFMdvH9Dqaz4Oe3UmJBRMlg+udgY6nQ1nogGu/FzBGLmRcU/ATphDrpq
cTeBFvpKoBgshhTXscgXt1KfEPCNJX446lhY1LM4pqlJqdEoZOfhoo4c72coIvQ5N/0GpLNHd5pd
a8puOLAT6FUHWdjcstcYADJ+rxc7f0UuECZ5+OF/a+GKSNvSOELuuyhw8n8iBq1dlKwxO4ucB47z
bzqCh9au0sGmUSijOMp4tjsxN5pUvtKiVBNZ+NWcYfjwXtOLGjNxI848LSSD32DqpYncZ30T1q2o
t82/L+BY+nJoYHQmV3+FN7eP9/pvVnF38kZ6x1fpVF6QfJ7op5nQzT3C7/x8eiE4OpkQxqSCicso
dQ6pm6yxPAr8NgeE9AcwKlEi60BwGhBhwYAMFq8CJhzIYIDlSckPgyqd0UNutrJ3scfdrJ+WyyGv
KvQgVaWD9nob1+h5BuMVghH4gp6NJ+Uh8swtM3Za547OCnF2Elong5ywzjdtQzN7Uii6rePLRRJk
j8nz8xrgiPGa7rGLXg1VnLbm+5dMW/vE0zHfy+l7J9J+dj5+jmQH13TD/iYGjcHA0h99UfeQBVsY
RbEcC+JYiY4sPGX6aUiQKrmNKkb1lYjGV9B5D+FrFXr6lxdewnw0cgMAitz00+ti2toF+Fn6khTA
A64F3066EBZJkGx1iDVlf+QEhF7B/bhaSfD+XRSJNFJxAVGwgWeHSztqXgB3Y7RSBJqS+YLB2GvD
7iMuOwRWtTGRRyaVlDLfqy0snmv6pUZrECdz27AJG25J/9GhOVtdbIgM5VR+py/GjpXLu0uS5v0N
1zXKs7tE6iflggY9PjS6gRy7vPEJoCQSstDLcWnRUWTB/4zEnWV/Nxt4NF1j+wY0Hmmk8cXMZUAA
L1QCqHz0khCDoRmDI3A4zacmo2LbKCi6brN+LIwsr+vgeQN0FWB+iNMCXVFqYNeNTQmGnB3T5Ytl
BlLe8k7d6oQ3/D205JnkTz5XT/zMCXblgMVm2oHcMuWWbLjU+7NbB2UBG6KBEGVczPldlvfhYNKp
pHmFP1m+iff0oWiG0waaKKpmlN4SfgluMP6S0J3sL30DwBKlXfJvO9uGGUDOKSBVXJ/9FRwV/mVZ
Fe9U5tqHctZQ23PsF+TmtRS2F0liieq7E9XXag/mWhmtLb05DvK1k36xOxTxaAQ/mOODqGy31oJw
uu5H7NWsb2Zy//KTK1VVihXJ3PkbyUfp9oxQ4GR113uVu0SF5G8LLBqtaNLrWgmHTAWKyp2dyNB/
RKRNydCEEYA/61VoIO9fA7Gi066ZFtS4T4zAgYyeGlPVWF7bE5e6XpQjKmOamP2bSh1tAJhYxhVf
kYJAPNaIsDgIlJ8d6AWaIQdTkpW4LyCosJeh8Mvps2oQyvhYCHw9MjmZo32tzFsJeT0IZTHuNE3W
ShmwhlkKtbVDTUziglji+5M2FAkD6ZXK1EI28ilY02o4M0X/jpfFTWq1FFaa1udYbF+0RxdbdaO4
ZUm7rZY2RdiaezxwBgfERKLT81AfFms6cslRbozBUEAlFxxmhEwDmLw3gNNfivJ9leKHCI7MrTxA
9WpN9ibJ6CnttNBAcqcwsVvMouOdxsXwQdR1V3ZD0+5kpz8mj+wUwNaU46T9M4p4MADJWLCCw1sX
aFXwHdyEu3GJ0a6ErpqxAYwDgbQ6EX1euNG1doKo8d/80MVU9c0XLjwbaHTuZmlZhJH8CzVHPzt8
5EGpZBYfKCxdvZ9l7V6KF6QWT6WMe+aDwUsdyMSFpxS4LoHIh2zcImEJ5EmbRe2HvGL5xd52LU3S
fAcRWxqL8VyKAr6ruhVobZfL97maj/qCZ2iD2pA5kk5CaVLa7pOuR062qyFJGWmbIvgySrTyDLMF
zsi1cDzdWv4JNlfeeIGbaAxwrk3FzI9fAT0zCT+nBvTLtAQbRc1Db8OrAjByh8Cn/MXkNQnB8UDB
RgLlrfLYoI8MlHwrLThHd3MfLk2cdF8g/rxl80YSWG9giD/YY3MvoAPNZDoipdRl6GTOLsRx7bvg
mrl84RG99Vw5HRBtmYTl8lVMw8O1pHsWUeAu/70eh9oM7+l8hieuhCUxnlVqBhGC24MV27ctpvIE
eKKibHSOzlhUwN0ZQdkR9KleX+9CAjT2y0rx7SGwHd+JOmweFuCtGjezl+RRif0ee6lee0iAxDUN
OWm4dYDkgGXXL92AF/h2Y1Qth+pUKASEeNcQj2+rBqGQ4/AfzGi8Xix3/vsGDAhAPMreeUBCpRel
e6OHTwvV0BDLIvSyrekPY23mc/SvBGhYcwmqUF/tcssIF2d0dvAB3duS+jGkiow2G27+B61kNJpE
fpeezr5P+Q3HeOaBr/DdVFoFfxGr9PHA5kovC95VZdr9zDsQTJ9llLZaC2uYvlrss4+OHyJPDbCv
yy/gc+ndNP2KxKzpXNAbuIAABs+6RW61Vb/ZoAKPeKkUWag5ami0VtIWD7ilC3iBAJtQpRJ+MH/a
rmuGp4N5vJW2yPb+tnpRc0oweUXrM/fzLjwBQvu+Dxj6vTsspi6TShudoKMrPKiJ3xVQUYi/N20s
AKAP8kGu1DabbX1BzxudtlJNrJN1Pg8aYBSlOGYOl0GC0jgC912pfeLp9gjnBpO7nPiE7wf5irjf
MPAf11m6jvhMVn1G9Uri41DHQVrWr9Lf9pCihLDwT++rlZm9NLMJ6Kp6rahWir4PJwgaXUK55+nI
Niv6i1V4kEziHFxrdmCjx84JJOg9aUZ1p4CVi8ohIP12IsBVk1TS2avPVE3Bs4u9IqVKUahk14bH
jtWTwiLjGdgWw3K1fSdxBWlu1m1hpJuT43yl0VJo9eCAm2qaLJ4/qbEaVExIckV8UvkC7cpuUMAm
dEWDjVj5aEzvKg3yFWj3sEng4KzavvZbG2oerHEGshX1u+D3aofSLV3kuOSpIzlTfHSGYuesxvmG
syvSikNEeh1LvmUcdDpEggqx+TZIFc8Y3LtoDJhFUsJGG6EecmnlOBxD3WQb4M/i0MsYEsA2/UEm
2W+c57q8lM89egQRbopnJyvr5E4Zx+/B+8LQ1IACOQVXGYwTCnjxjooiVkGcQ3w1h1IBe9YxzzGo
XZ3PmAWWkDaXRxlTkVKgOx9p0b22LNx0aauArGdZr6+tiHSfnDQlHYPHPi/tSoWPN6smMrMW+MHi
GaJIxqZKLKeUP2ic2YIet5gyIKfbBQ3p1eIA5ze+8ZyuyACIPkLNLx9l6ulfS5ZdJ5Gn+x0RPcoO
V5F03GCzf2RLd9CALMTTVervLMOlBGFqOUqDG76TCzEYg2DpR/ogS1MfZZZmbFrYy4MBkP4MrV2g
JqDVZmiAsfldG9w9cItY1yfKhddNKfuzEAIXhu5KZyrfCz8xPhL4jyJcvNnURPQGhgrL8Vc26rS5
rUlk14x4gik2zG9dbkCAXjsgy81we9Yx3kKzWCGvE2sImx+cYTOTRiMYzVkB0Hczpn7sEo57bVdW
jSRa0o+yaRqYN4/mEYjroiT1mpj0FeVTQjnsHAvCFu4vLl5JTkcf+ti3DlDsvtQc/5jl2HFucsSo
iIU50ENq677NJDcwM3MfESPliA5B8mJJ9QYXziK2mjDEmi4f8eDgG5Qxe1WVx936JCNoiDfB1rjx
JfXTtD7vV/QBfvkxX1p1w31ZYjOyW832/xbGRMoTv1U0cE392WJxJdyhh+I/4Mix+XExZu9j9Eg9
jYUJyQco8O04hp1cE10rSvqkOX4jX5H/1w8YGCQYGFa6kGXIA0aG3qNEAtOLYPwr+I9j+UZRDPwC
f+YEZ8dvvmXGGIVp0nmTJxx7n74F/NDFjVS/v0g9vSojPHbUiUUuAkFXZ6p/W3S7+9zVPjp2FuX8
ILi2Ww8T5hWPcTrZ4qphi9mfKmsaD4JnP6I5h5UmVQKPkkPyEndALcA5v+F/GFb8Kjb55VVSLQJe
G6Y+VgC/75rZIADIeyl3gFhYAmFIilGp/YFDNDGll406P5nvoEd6e8VRRvxAdY99fr8Vyrzi+DXh
JUdE+jQBZFYbcaCU7tqftRHYHvmDjy7tY1wswV9wbKXVSaHK69JB1Fq+CF9BRnplhO3PnQOw2EyV
oSCR4fnmwP5oPqnBdVzH4eJRqesYJCLXeqIbVshsjBCT7//Tv67s/jQ+DqPqVHxQ2+rVNnbZTN+Z
WCU8+FAtmH/ej0jNlxxJSe+cibUXRkNBL0B68Sy5qyTnN16bM96lNij3YwS+ojSYUcuXYZyKGSpi
cV8CLLNED2xyq4Mv7Lup6keNCuoIAQicZfwe7rpoC58stCj+oP3J8xKyh79htvoSAx/4Z+7y8UBb
Of2E2RYoaPff7vRemrF4C/0+75Cin58TbF5VpTToTK1x/XeXs88llVIAqVvOm6MOWO6ZPLBS+Ngk
qP9EoX5cUSydvR6G9gydRqYJjNUaNeB1a1kphjguB4t2XnMrv7efLiLkBkLZ7f5b/ZRJiV/nJzzg
nmgNqWl/x593hPBl6nRBmXZqDmPqgh2EEzmvLNCbX7aeaQ/P033uxFgZY8KkNrnujcWS3DzVBGO4
YjSMjYSfTWfrDBOjZHs//1y+fPCG9vKrec5p+92izxYEqVZANEVV+/ps7H+10vqtp0VFu//5YzHy
mi1YMdru3oItYoxf4S2rjK6kP8u6Ks7+t6jalCZqNi76MiAQNt+i2Ejt7k84etOFcYpuBCr4Q4Gw
3QN4Ap8f+d3yn3Te82dquHWYLNFeIK6ZxILnyXmMIXpk1EFxT3puSBAVT3AX33JtGfqFWTFv/YTf
fS9oSjAwJmmZNvENBCjfIDEJvong44WjucOPlrXwImLnKH9rWOJl4a/BM15N0FkfPfygNFUTE9gC
IV0MXKjzjow3F9xWIXNEHtFMoyLfH9yfBRfIQ0zt0vH+k4qb573Py5CPShIWhcm2vNPC32m9gPPw
7mZYT2VozHIs+3QHV9m290VG6tGpPfGAvfM6ngeBkg5c0y39jgku28oUCKMYg0F+hD3jovkP41fg
5WjjT5wC05QazvgVKCZunqG/K5MdRJP0G/8HSQ2wPFksS0QzvH/u5g4DDScT6LsD651UsEQnb7IM
ZZnrr/09NemLUJ9dTWPC98eQdOxZ01fppY8o+0mm4tGO3pWEAW1faELfk68CotGdclO6XJvqjo6R
K1fbciaUzXJ+B5kAM5rW/X/rh/YuOWIcSmf8SyBNIk/henVbzha3wqN+ugnjOldQX2rLXOOTwLVm
1BGSCViF7tCLym2aZpiFxR3TieQ2qFMuKvpddPwJMuWt9IRa6Spgkn2T4IBvrzt1P5HoKPI7PYHM
SjOndkRdZe2jKbtN389U93Sm8kxqcqQduGahxAENeucCms61I346F2CSBr/oHoWIamE6/7uNvCZR
eqM0xVCxfmyPdnhw3RFHVTuzRd2J43BUKKboso5xlCfvh6QXpyMh8qrph3tGWdkJo8mbVA4bU2Pp
oYuZnvypXbrhawR6KPfhIh/ZFshWcH4uLbVOyWjc4KZNDji4z22rOFr+waycE730mJJuNjZSbQdH
eVHymU6CyeHJKv8vm00kUslq0sCxQdV9hX76wGzSl8IUKhVAJ027AMDB1n3lz0CBi304qsgdrQyF
22pF1H9/AeaNApfdi87yZXUB6kj5sbEtaMU0ppDnMpyh6WiCHQXoma62qOu5GwaMJG3oinB75R+j
u1rIKm89BtDKvZps3aVfv6V1qxIJFlu3OvIOe/c3eBR8fOU5Rdx5c06Sx3xo/6987dX/ygUH2kJG
Du0smnDyRR/6SoMCW5FFRjRmz1jYh9i55WyDfH7Cys/DBj6ejC4e/e0dBCSKdhcQum7au19/UpBW
Uib23fkAzuuO3SUdVJhKY4Ip8WesgIWoqGOs9gHkxKIbE/Bk7YsgSmY/Ntu/X0IFKkoUN89vD2FL
tGTS4qrS8lLYcP/4qrIfLGjpbwm2nkAcJ5Heh5cXwRZBUwmtAzmZqWtcFL1yyCYJzX9HAdFvO8SO
6d1NebJe4ExG8FkuXTsMoqE8XXPXIZPqnCM5WZUPGESEuJ6VBBCUF5s1sSKz0rd9IP+PyfulFpOH
JR4nnZ99gMIHLyxioiM+k72/4PaFkN/yIALJUxI4pHQOwPJz3PHnoBFTzU/4Deho2nAVHrU/bNOK
AbcmQwFRkfd9kVabIgaYOtFIU8+fK8WxS3/cmWurg/aY5McURUFjBzU4UrhQdoXNWa6ISG80cJdM
V/eHuJNHPMWanemj6sKu0AC64ZBK6z7rKd2s/h4+cS1lKE/3vbvpBCwtcKZbjT2HCfSoCRK4wZV1
h0xA3x0BRCQ8APUQGvwxF5XEMIICP+AT2Q/UqxmBEL+AzeuamjaNMkb/Gys4oQqC0zb9bfdLyTKO
wQNDfPddNDp4LYIecIl2ECWRNe2G+wBVH83PyEwoFEAJEum9ciQHxXgvzVHdhn0+vJfMqdkUbjro
VVg8rqPWBhZJhR6CQzHUgZ4QaEgk7dE7H6wC/MDWC+oT48Rcww7puooX+PqTkcTmyLSujubr82V2
cegeJ/rQ0Ir1ye2TuN7JXGUH4bMbGFQSkWjFOOS5+MebIxOnYeUpOBvAxnnhecjKkfNUtrY/U64z
nrs0YkINeITl4BTCpqOL6s6ppDzR8pqM5U6VzlGHQkbt5mVOdGmsSrCmeRifta7w5AZBbCCFBRAQ
Dh7pWZWxQaKcf0mlGPRmpVJ2fTfLPbB9kl2NQyvB2ijIJwhkIRbHWdZqgTLtnERWyEphdHdx5vUG
NcSU8wdiQgb8USIIsAXezxrDWblF2hkRghlGD2e0OqvoYH8/6dZ4e5I3BcbjJv1SUjmx2wDdQx7q
31rZNe6GJtQt3OSE6LBDh/l6eiKnpP7QBlRL43/K2tPh+UztDInGqxbwqJckqnf0SdA5EomeYdfY
zdrSOt/B5dGawbwcr0JOyzxUc/0IRj4q37W+T1UuyZN+zbxFmsXcFtGsYp3j/LVCXY9XinkX0cD6
PhxCkdfrC2Mk2qI2pprjt117PM5UK36EONnHMwJmxIWE0Gnz/yOnn+28Iv2D5glzakpD9LOJW0Oh
LeQHZNIdHP+Wauomh2vH7U2H3bSzRQOXLv9+hp+NER5l+9fjiiOWUKKCAQuGndhlmwv8UsO5QeSc
y5jxZXQqBHOkvi8VOs9L5rVlm26cxEFCWZWDJ4O+UKmsdIQxFngNxheESnqYoFT8xq1qOTyInDSy
8rrZhM0WjvmIIJC88S0BWAWIltgzMRKyRlURz+MFpzZ8Z6ND7e56AU7PJy9QU/IDWyPI95E5gtI0
pSleafGHH/ZaP2AxS23UNPnvhCIMmEDcXFCG/cU3lwkID0uTVux1bcDCNBdAI/oRMk9LyoNY9AFB
AxB2RiqyI4Je0LkqXkc2ovpPEF6fl/7EAfZArluLxj1hnMm4wNGksq0S1lXYthWumkQewq9/v0Ma
YoPjnE8q/Fvc+63dOfqztd9GOxFF1k2uoPYj1Se6p3FDsRVPNidfviKKboDBYXGBzhkjFn5GbR5/
XRSFPXv02J4ucpRDW5jHGdQLtdSdt+/dhscvAuSznMAGQ5CygQX5l04xzljjCbhq1IowF/sqSiJH
B7HlVgn/UJRTM4A8Ody+YGv4LWj6c/fl+buaheis/vQOPT03KMxDZK3EzHJcFM72UDKZwvyNMuDh
adCpEgLZp/kPeptpfYARL9b7FxYLsHfDu79fZfsHUDyTvbhUDfLqg6bilayo71N9YWPYPq8yh77R
802HVGfkfCEHH4nJhYt0BOtVQ0NWrIY04nlRuxTDk7osolHjK5lCcjpAkcnG2jtweiMF/9DKvWpl
497p2Jt9++UUikA+crQR1+7PpPcH24gG9K1G2D7YBfjmyT/G2vbo9gdWXQWL3htu+IatZueAIBhv
ecpaGriPZK5xg5jyQxriHUVTTy4d3uRNq1y/1NHTXJScwHPWQqpr1KrGC/fvLiPHxvKFOgDYfR2t
8tFaN+rsojR0oFuZraPU6dg0+f9HPQESc+jftLaB7ToLzRrFIU2bt3LYvG4WbAERIoq19l0gcRC+
upT70yFfh7PsfrY42FNwHSpOJglEHXpzzySwJZRZn+zCl+pzmwh/9jdwXztxiscXMLFSGKpLS+10
nZXE0GxHvQJP9nkcjBmi+MGrWJiSgH67A12Y6dXKG7SHUiR/J7KGXLECEDWFqPoAdOSizBjo5iZB
vW6yfvR39Rc5htz6MCl+9psP0tmLqCjFl2hzadDRE7sMtlmpOIUV4YbApV0N3E8Zw+SK4g8GyY69
1ZBgjHvJM63pRpbpaM0TGz4otD5i4I+8NF0fKc/SK4rlhAoM1+wcCt2lMSf2w+SWmLUPDL76hRbH
z5ux0D5BPIWvrIj8u7FddxVsK3ddtfq4/mT35DwxH20EpOoBCKDVWcrLnsiIBRImFguXP93t8OMa
77C49+y1UdEBcUx7OTjUgxHV8M+nFzYId/vZPE1DdSWM1J4elAx+CJPFjPiyb1edt3UNf2VJDXBu
Xd6RKozEmAmyl8hSoUw9f/6XBbTgcbnJlroaLK9ygTPNkVuHN1R3uraJW1rjZf4vuh5+Qe3M6Gr3
Z0wQQpOLZ+it4m2+fn3J82Nt3m4DfcuFLLBWe54ACwY7DCEepPSI3xUDQxpRtrhb1pXRr7zFV4qB
8X5BmMnehxoz3wDuuFZ1zS6JPDmqyRdMyfLEAjM4ffy6zoE9r32glfSL32WWzz9R9I5lW5Db6Rjh
/7mTuGJF90kNkuHAlWjCgDkhYaLbPVO20+oB3lXQL56fWeDgTTfc5QLMfyBDVKEdueZq8FJ69NS3
n38rjXF19GtuQFE1cjf14joIroJrZJme71H4aufmdBO3WxWAovoaCn1vuyWpEuZbSMA62BAFt5F/
a9pzJuZ25hNF07VARG0COXxnfkgDYPcB5Qm6L0cIITdDe1xTAE1TkouD0Dh/COotA/An9jGIR8MR
fG0RTOMNQO8xg6FnKWEdtJk9AkbProcclFWGcm7eHUoOS1+v4395zjp9KUZ6SpokkKvX+s07I7lL
R+F+0FG5vH20v2+tuuxZNPqEwyxTebYNbouJsAqU/O6lP0NjOTbZSml92wTv611i81qZ15QYLUEm
NuqgiL0OrbIpnu1ncj5bYO50pPIZgLbzebiqXj+0b8TPgUTix5HOZaLrYEhKELizsoAneHzV1Fol
ivw8RWO1RIZRIzc+QYqnfy11dwmPHn/CLr3M6W3SvCDVFk17xMmuupduQyxi7oChm2vQxsVpvnHh
eefodYax6TPKftT32b+ZknFzptO55RCNIeKja30utrSc8aDxNdZJgmtX0NybkT+OjiXU014ufgAo
H+Nb5ox65A0rbYelAkIGhr6Ad9M73fC92HcvShsfAeZFTf/npZNLbQ7VXnrsAQqSXqQrOFH1zti0
P0MA9uy9UkYcMSdO9hZF3FGKM2EcVEzkojVD0icjryrLfQGI3slEmAi8ng7L5p0EqD3dafl+FeCf
W2PO2PApbNznm0kSvywX5BxA8wC2WnWBOrO/qRvDoZErD2jwTYg6K7BQVnMFks56NsEww7Mm73PZ
/w7iJ4Vuxk2Ua/ho2kN21dcgiNEUX4BOCn8TUF0ubymwJfo3nPEfv6+z+ymiC0y1sFYgVJV0h5Q4
LJ4nWPJDDO4lNHtnZnRGrioM8rzhOYknC+UrcSVfZgzpxWl1oG0NoDhdLrnsggwJIsCT4psivP/l
3HCUhIDgkVKH5LPDvZR8/pnaknUGHnwTi6Ccvhdjg/EgyfyaxXgrF8YpuSYdsmzAu9DGisFMXwgT
iN9sI7yc6Bp6Cr+UCci3twcGAG0apgcZooX2vEUfc+ktKaXmyhfLfFEV2dVswGzZdoxJJSRZsNNB
qp6cxxaAypKAGKao0+iRQOUjAMYPDjI/tI4hhqf1+dqEEgjAII1DS21GC+KIfcXl1FOmBp/GEW2f
EgMKo3PZNIF89Bs90WCIzT117e0QEeaqQNr29Yclxfz6nC8zyVZsU/3Jf0LqmhNZja+Uvk5WI2/V
CXes4MLbs6s/0GFoTFcPizxERDQLycVqduyN46otLwbDzpcJnll7XSvjzG2xbibXhyhPw28N9iFB
R582ZTHLkbRY476qa4t3P+qRgm2yPHseWVpp97ZMizmak/OvtV1aCc+kltNG6djlE9/45isPqKHu
eBM7rxvZ6E9iL5FSq8IDdfEgmMB+GoFHibG0vhnKBwWehGnf0BLguqKw/0vE0xVV69Jdbf240DrP
a1f+TUHnSjn6Lyx35hZuQF5Ou5qOZDsdJNENoeBSJqBsxEVzdj1OZ2Y0SBKfDJL8/JCa9FXpeQ/D
8QVF/F61s5k/r/5/kmNsuYW8EmP6gMeDjREJBH9z8Q3kv+XmobC1HCVs2Eoq/8/8KpXWdxEiMzVr
hGGi7nznhdLSPyOvpkkv9u/67OULlFzeesEAR3FT+BVrRS6vgniVh6fPMZ2s9MsFYD/2WhZu9HSI
MWILMRFsTLcAPA8IvW79gjYcJDKYQ50A4iQQ7bd/4lVZ5Vf7huruzkMY/HjEC9NVbxZleTEotANM
z4x6+KNPuup2hu7hqTrVIoWoWliNBM27bbEqLZqNZ7x6ntPGQtslspdpIQ8S+BFLuPsELPLu5zkG
eLmRxgEXpIcMnuckI37+ODQ6uz8Ny+piAcu1c5yfug+PS867qtCbrMJZZLf6dStavyP7DftqiYEJ
YTE4lkir0fb7xYgnTG3V0lVLLYK8x4zlvJYAu9CaO+MbKwpW7useNEJZXkuWFE6JLP/CuFOSkB7H
e5LqyB18eUtjJg17FsmAB5wFt0vVJPlDCW+Hm+MQPCNlpsWWKr4TfD9O2j7RSu7WR5DVKVLQJ06o
UA+GA1IbMbbq4pypSZXd8AgLUq9UKaJ91QOKLGgKA/6SHEUorJcXnibn/MNhTsA+o37cHoW+cLqv
goVgrU75rXly9t7V0r+PVnZk3czJ97pJR3b6kc/Tk+0lzH2d7G152xMo5XPhom4nb/qQ6ELt+rx6
dIjnYAvEaw+2bNkycN7oXZTGu7fYIjoUlM/GNDpbCqJqLBnW2gM9anK69ySymdUSrpahqNHDmGN7
I5T80CK0EQbVi/hk2BMTbMxyJB48W887Pc4yKzjCpP+j4sFJWsPZOgspeORayDx6R4ynxJI8nvp+
ufdXm/fBvG6CvteZwXrG8Mj0FlKHZhwGMSbLg5etx4Ijqnr1o1Y2d2dFGRPnxgUOE383knuYZOWk
MYlPem6MDCzTDOPKPYctkdk7vhu2LGKQfaXW5nfmVzghz/sKp84e5KFIK7ORJV0BkJWoUGWRf/N7
EMwZkNJt5BWIlxSxspsSQmg7Cch6H8bAV/VzeX542fj8NORhFd2fGYbBZ0Ssg3u4cRMIrCOtFgQP
6+elQZsmwf4LXk35gZh5vu4A+wppk5XTrIamwPhe5iwV8Wd9fMeRjkaajiqj/MaIN//2t9hqRGUc
o5z/ljUzCsMZ7ASXMjLw4gPZ5tJz838nYi4zgu8wx+azvxF/XxIWRpD3XNWdjoQTHS4r4NWFHX0Q
sb1GlePnuc4o23rwVBF9TWooeGgFB4/Me9zFb3L2yZTciVMwmQL33ssChhuxovuFaM0L7Dm3B/dm
4sqerN4fDgL4IhI4L2M92fLySIOXXT7USTR4GwUcp663vtTF6HieM/XWaZXsh9+fJK+fzFi7aWL5
ug70ChF8kadhTO/li+nsib8jb1PSa+0/wZj3Ldqi7dxhPPJ/gJWVSjmuvP5KviGTTtoOQnOWmOJ0
Rc287P/R1JSzR38+k+vgYXjxceF3mL5s3HuERe7AFcLW1MQ7UrVMJeook0VPqD+YgZiwSZWbxSCB
Mar1n9A8Rkur28slEPiE9gGY+z+dUQ4o5YEGNLGq/qy1tgTQXAf1jvGm28JGCtqG8L2TI+w5abSD
fRNrp05DdF+gLuMdtZHuNjv54Kd58H+NuvWZOibE0btXMZlrgB6DuTBOT8puV49JHmVS6XL7Kr17
0Q6HSIg8AFTAB12tvhWCZh9qsw9Esl1MuVDxf+LykumASc04Ty+BUojZv5Qa/Dfi9HBj/6rR9KjF
iO/FH6CXrmXjQ6dbt38opfRDD6m33OcFmDthMfKdAMB/fj1Qsbgms6B9Yh1T54CuKYOB20uRG1NT
l9lpta8X4QOBmfFIEhblBqTzZ7LSrTDmTHGtgsYN11T0yVKw5veMQ1h5G8OFnSbtbDqZbgSY94R+
8CxI6CFX9+sQSecXlt6Oq4N9afU5ovHUD/iEitzlQs7Wofo5oNDXzoByalUtpEOJabJthrbnjHbh
q0TmOZthSbT19+WrhUkmxbJmCw4VfsNG0mMZa5wOSAzcg1i9hAa6YJTJ/M5BDEpd783I6T/UfN8q
s+DTwReYWtTitDBxt+jnRzdbaJi7+e13ZWN9QY+fGxZ6TYH9S3aJ6+0y89caGAi252dR0hWS7my2
9TbLXdm7ysJ0vk4mWUTI4m1HXa8xTPhhIj/HISrNqgo8iPQX51ijO/kz1XaNWR7hW1F+NUEhaK2q
0HpBthl0Q4cbnUhaEZ0E+vfyucnhziJd0pgoRw5IqM0UBSutY7rFWRXyuu7Kao8ziXqSt/qszyeT
kJpqTBfxOR8s+ZUljXanffuyT1B1rJ/9Z5RmOInQpfqo6YGC/lsOWaS6aWFvfsr61oDPy2FPF02l
uefh+sfsgNafQteNA/Hn94bdAzhxocdf/J4xKwYN77J1q0cdNPf+TeEQDMRvXv2b+/+ifgK37xOY
C+hHUiiorvnPYtP7jWxmAbMBM59W0jVppEBY4K+akOvnCINSaM/eyDGipY3xjjx57ZgjfIvFpec2
kAeesrkHoA1VAMshoehFqkRjN+kAhL06LvVKNFM0Ia53vZexFa/TGtkXXxvjZ/DzaiS5z4DTcXBr
5l8la6hTQKBmlNxxcc3qFzZUCEU5sfvW1fzfw83Ts+Dj2BcKWAEJUUQrlk/681RFwvXCPBRNBSn8
Lmbz8AmUkqJpfgaKiW02VxnKPtszBRZf88Bq+E+1G+rLZIg8nZYF86jYTBQW5eGgAO8wnJvTUJ5c
yaG8yWPHcflhk8L5lkz0IsUL0BH8ia9SomIjf6EwV2+KBInqu+GNUr/fhpiVqi/iTLgY6S4xN2sJ
Ux9nmGuUZEUq56aDbwhzZZR4X2hhbD20v2svLPBnVYdx9GHUNRTTm0XXc6/UMwqXTWuY2WvGYqES
4hlIZKvcWZbhStAq+uQ0vGL90Qj2ttuiFmY6eUeEY8jHUWL1I/tynB+wNdWfi406Y9InwA8X4gzz
/s77LeXR2lTD7aXqRfLWwF7+ubunk3AM6FpumNOPkfoh5woYGaavsiz5rz+jJ/aDYLKkMjfMQMDa
xGEAS0gNiYWdtTY7D19kzjIl56Zn+yXX6MSQqr3qW0Ycz1ZSllDBl9ZzNl0G+y6U02vR2Xh2P220
v9hpGmUSSuTPXq6vT5CQTPO/cxNUWt8SUKhkan2JraYG4eTpjdVqeqFD1SIB81kNHCv0jgOMMr+B
dszx5LkZDojLMzNBxcBlwh+ejKvnoEHeuAJfxO5vMiJrHvpTmpfMCmQuVyTVBeEhkJjN9pZuLFFk
S5JFJ+V3PpeOHz8DZWLn/QVBDm0+9o12QHgov0Vza+WgP2G/3JbTmith65xZYrN6KwpdMq4x0v09
gfPT8I8OF3+7fk7aFbjC7kX9XWSOC7aDOQyN1FxZOSiiIG3+rOPzzhD02hJj0X7hkAwVaMnG8Ho4
DDi2+L6438ZScC20jfcmjFt9D5rvi3TF+99njU6rPrPOgaylBtcW7lE/IHnP992w2tD7bkRFUMGu
lmq9s+cCk3XIg6N749gMf6Js+SLhyrYpSi08UOBTWbIopvR0Whn8YfCUr0qvHF+NCymEhkT+GnFY
kyrL/HdJAH89WB3vxegUv/M7CVratBNXOyQAXsVnOrwJk+uPgxNM3JW6nHlD7aHnG/yptcDO6PVj
4H2RwdTZyDpPUbYwdNHuAQOEiWGMJIvvzD6FfCif6DIb0McXwYMCCu9zKBMbKSQNZOlwCLYx36jZ
Dv1Ru0UNw9nqsyFfDIQP2dFZxCsmFU55Yez0fFgs7d6b5eZ2tY9tYHaI3llp6xkNJ/91l6SAoAbD
akEq6nK2Ko1fdDUFLk80hlAWI6uWIvaZStQ7ZAvAgxypFad7JKPCLiSgpkm8nYSDbWjst9B0SgrL
2ApuWKoCRoPciM2lUMZ+Z7p6pWtwIBD3VfodRb9my86CAtd2cHU64YuGWs1JHHyjUR58roBQtQrd
BRn4I8TavIrbnUQeZq9LUgcxdygg4RgGu7b0+3inTwdWkX5HHqh9GUByYYOVGEG30MtIwhJShqT7
uT9akLLVeQp4JbKCpJ67nNuuWLXd2MtLwMcHMVVai7gNbt5gegUTCFseVxJ6wdsmq/S8CZ9mVtB0
KX+WTXgFxyR6/UMW9X3TRRXL3QN0IyHZQjHTB4V67r5+VFBA5r8G2Qe8Bi/vaTNaLY//VJJr5v7n
vMXLl4D9g5FOMTL4tY72GtcawuT9a/UGixZes2Zm4LPn22Um/1fzGjF7mYLzUmZyGiEBpUw8ktI7
ig95THdoP08up89jQ7t77lJCstEuQt0mSxIs8bH3/pU9hSg3TsEHVSsWt+Onqg9S5g9L6TT247zG
IJpb0aVrqhmBDrJbu6Onev7lryWY+P4MtEpvamhCvtgY3ffw6aOfVmYxE6Fsx6RWi3yZxOoyXeqw
WrI5eXXeoUTJi8t2aWI5/QTzEnGP7v9ZxT8FEf/dH94EQcO8/OgPdtThnw0NvhUbdzrFMIvmK2jX
N7iX/Nm+/8/h4AkznewZPkLHRa3oMzsBMMwKhFmP4xQDoCAFVRqvXEapOWzBpYfhxsJCEpXN3Phx
Zc3SJ5l9F2R3PGhHOCnw8Qy0bmlY4ULMYsHp/CFQIVFD8aG8ZYs/9rQl6id4K4y0wXIYLXhgY+hZ
ooV8wEyC45RAkD8O4+BjNH7jFpdnDNB5qK40YQp5WRpfjelO/HXc6XJHPDuOnh6OVpaJvfoE7MxD
yzJ6hCOYQvJDkpPoUaALrgqlq1tx5CW+pMeA+yq6SBfUGdKwMrGoQg+M1haFXpo6BpNwAJohy+Er
kRPw/YZFJ1UXKGL12kswoTj8OmuPx3waQONb54xkgMaqslBeeDyZI2VLAXaqS1TxWaRnO0gnwDJZ
MyOYQtUeiKgKR5DsK/PQvkWKIK1Q/FJHvK7AZKVSFdVsoV93zXA0+mcTHzmJybnteEqD0hRCsXAP
5hrW/y4ExS9mSOye9cG3hGhGNwaeRCXve6unb6Xh1KbZ1HwoBH+51zT6BUckUpvg28SH7zhppgae
7C4h7O+R/B6dCsKeR3Zlj1g9kI/pTY/WHAijppUc3j9yiX+EWnjzwcKEuL5sRB9WWlIPyfwWQwq1
OuHH0bEjyR0WDFlyHh5c58uqqpLzv2AwmnbodpBiVvFKjSuCS+0w0Weyd9esc/vjclkhyUEfvxsN
cuHMfGGfi6rHAK/x7x6DVY86Hd9+7RimcIeYK9wHCtfY5lMKhn2LYuJFSCQ1egnbVshSkhOXRSS6
O07G7ItxlzJ22jXEgdFzp+GiZqqk4EUwPCOCNIcIYSfXZXG3Aw6HJBaXJkrhhMUN08PH5+EJ08iN
PiwwRm3lOfapoq0lzfUhKlolXsziMwZGzef/2SLLt2oHY1WrvpRNYCivmL/gyKU4aszAh/1+byqU
7srS5KTXAEk0tC9IDjd+/ONYjUOPI7zcGJ+hR2k5/nOO89OafR5y6EJ4OV6aJG1/GAWBUBfARpEb
AlnHntQ/AhUxxXkmf3Y7INAHc9M6LTfveEELpLCiwCsovZwV27uH+hj14JfY5NJyX99ipq+PjegM
zTCpAdRNoiA68Ybrl2+QpwVfbFeo+cfezAaN9/MqJb2URHCQLuG6HyYFkcsskP8PHZGeO3H7KmlY
vhJSf1O81SNbLFNuoSWwQO4lb7kq+PmhmIXfITN97RsBxJrhXsLwrU7rHX5CL/QY9gVMhVUr1Jh6
EEyQbffOT3Na4CHQAvzRTfK1WMtp5BvKUyNFE2D4wMZlyEQQo07A11aMAh5JRRExkg/RMobDj7h9
RrXdQHbUlH9g/0tCEkzuikQ8D9gdJ0X0/xD+j6tzE3JZgRfRIeXBcBSGJO4Xycx8aQ0w6TR4xBIR
n05snfuc3cZVCbySNktFOsJrVq/nlqaxcplaAxbj4XhsdIY/qV9g8eTJGNV9bh+/VzsAmImPrqkP
3o+G2neoZMDZ8pkpYdmHZlcueeT7Ryj5BC4i+sSLDfJqN5rI4svTpbQr4sNEZL8CLRuRd1CGL+YF
bMcTpPsjk35i81PXUowsHaSuFEgVpftzilt2X2IfFQ71E4ZJ/B81JCVFkZkwcjaI2ZQXTPfrYYwE
bbKaU/Pce+s/Jkz0TVPK1FW5jeyZfIPzmq7dTOyQF2zoz5clcRp/vK/0b20oPDWQ/J5D1swfTbUq
2fFPy2iZr+/MfT4NUf8NCpvTb/7rK7YoYWt4rcu9b8LQtGUZ4EbqIuOB54krrHHqHEJirDGH6Q1A
PHy8qQFFIVD+uPkNP2ZpGS8ac2PXJAL2ANce6jcnMJkrGdiaXdDMQmsCoteZBNbtOLwr/WeND10F
It8YehD4k1YBayORIMiwKlEcsLC9GchHeCXOAb8w7QaWauJ9zKkTgkDNslLI0y66h4jd3yug5Hue
M0TyLJbiGR7YL0HvXXlVLoSBypyXGkwnWMS0eU4KYsAh7WLJf85+O8SPd0xqixZV6u1JZOWq+qvf
qZYAKe5tEo64tt0s58wdnyCLOXf39uP0LYlWAwjb38APk2eBCk5z1nARjIOjUXwEhWxxMzV8LNX9
aWz8jKarTPfPIUKp1L+6b15XjeKrIIOMVd02c7p1NYs1+OlRIBW5K+aC/DHPhSUlKQfVrlqyvVrU
GarlRa4YEpFHXsHQlIbmpi5utFZ5j4+HzAsdDwMIK3QhTkZot2kgBKdAALqJ7CCbvpbeVI6nKqGJ
f2T7WbnVqUwOLvMXFftXrveu3ooFubaKKhm7ZYiAX5g1RE5wfhhQptnA6a8IQ9aE1qr7+muSKytY
4F3CCiOAIqhe5B5YQL6HH0Sx0HFeI8VRdQ8SAPXWIyICKlJPBr/pwK+aj8o/4pFeiwfiRuVFnl5a
xQmOEBbAqKVAsmd7YAywGon98TsaoYZRVLxPfG11YB+SYqF1IRqfTFzyzOHSClAe6amIHWwojOlp
CCyXLugnPlBJYX0JRHXn3ZpRCSAnPt0O2OKi3HbXek2z3zQBtgIGLiaZ/gOzVm/mq9CMTKWLWroP
6ycGSMdVeCb9OFxc48xNrEABTWvXTer/LFprLxNx+ZTlmEYuRfgGIwgo7JlKh3/awy7X9j8clEQ6
G6kBlAHmkPyDfKaHDVLpmmDaD0mWxIDyeoqiPEn1SQd+aWmVg9ZPV2fcQQWHZJwQurjz9Ht4b/1K
1JJ0Fo6XFRvJT7B+snD0MBI0Ap+VXhZH92QJ6/t+r4My07zJ01W6TJ7++rYdAGfoo9LewxEUjSmp
pBLuBu3Q0FEp1l7dr4Qo+9fuq//0qiPX9skGBIZMe3vfIkEQTzEloK+jTQivQ1KbaHfnpI5cYg9q
DP0aa+h8/5+B3/t0itM5XeFMnifpCnzu+ICGnq8cLnfOOuJkGxVU4KMnuTIT2o9ja/WyMOkXlYG5
1jlL1d3dkwzpqa68/QmuO7SHztTQyB52tDA8OiixvqygPr1gRGiGHT/1GQLRaWNL++Vn8uW5L339
Hr8v+A6FKTjeGYAVPJAKqNYXKfy0TldFUWZ1n8wzDTSSz93P3+WpjfF9NJamc9t8a3ZMj+x4wPUb
dKSoq+0KsdNdPUpLvaRV9aPDFNJ+V1RfUOBmMUMPFS5uIK/eelaPQvAvu9tkxYip6V8HaIPLiThs
2kqeX1v4fpJSdY7P0va4ccmHceUosmgkMZtjOAjZI+xH9tvtUMuZuaqHn1RvIC8TZZS2fHtmCTi8
8WPBz+HVPMfyPRNao9p5fSHFHXC6ByWHj4Bn5TStcah3tiFUVq7lc9FsoWDgGbdtCUrQayyaH82Z
sBMemlgWBK6xoNpNvvA+lsUrlDVpW5oO6he0dmUk68xaj0bBBNFqIcWem89IWyl65fOfSxV74XAZ
LDp+aig26RQ2B9H2MnkiQt6sfi2O/kmpVBjegOynPGNgw83UuCn6w06simtnKXc6o9RvjjADdxOT
9CF7FJ3FopQvfhxBpVXSmUn/u6MPR0EOwU4LUdqWHcC1PBpTxQqdGXkoCr+rDWOTUG9JjL9hpoQD
12tImmmQ2HGie0Y6ulGLRDYngv4DIEqN9uKcGwoec1IZkxhBwFw8RL8ERMZ7VRenxEK+fa9JGVO7
2Viz5Lde6W8/u3Ieg2m4r0Kx8SPJBsvkZZ+YPkdFJNkMTM4pLa1+pm/TwCP4GFW1+dxQYhfSYVy5
G6SSaKkcJqWGEyG0rGAdxm/EmFY466C07H1eJZM5qur3saDWgw91tlKdVx68RFH3CbBD1hngp+49
y4dhqJWlDH/seOBu9IrfLDkg2AfFWXZoWT60mzRO0d1Xd4VMIlwRVtp3jFHymK/Ppqq0dxLDnRQz
XPnwUvsNgpOflFoqcuKsNFioUAa/OwSelYM228Ht7rugCf+SMxFaZVvei2d93kjDRPie4WVFCuaO
NOw5K8t9vgWz3oBaqWwAKx6aju1FztAH5Jv6hEb+lyp7F1x7utowXAsN6l+D/q0IG2UqN3433xEr
zX/lDM+ae4jGckOkiKpc6yHooT98yZHKNZhnti2HnR2jgSJwyRuIQ6ctW4q8VYYKuV2NBsyMBd8k
zafv6yL4c1jqx94IQRjz5UzqJABB0psIJyI5ZwGDQ5PryvU03EXnpCaeReNO0kcYiigo7ERVgl3y
MeBC1D/T/emZTe7ZLv3WIuW8XXScKhapjq4hsMASQVMgfEZmFw9nOITPzTTChqKu6wKLuvIUejM1
LIebjwydfp7MpbG5OdIdPJbKqm6cklAeFeLu9JIrot/A4SKQY/fo5T7SQb6Oy6CHC6SxkVfRCsH6
NhuK+0vLIXqqPicKMOuy/hGpSzEf20h2vQE9xQhs9c15P9vlfR9YyiJA5+em2+nzxSsqTz9JQA4h
gzjHSHXHud/ZPDhj2F4n+jTw04neFa4DgaBVLFU/j+XmeO9VefEtPF5rD4I4C+1xhdQSIdJ6O5L8
rWMlqz20nuDFA8b5x8AH0gY4KAYUO11W+NbdP14kSr6XpRKycYpmxYxm39Hh+jAltOLrXJvAOgu4
AqDWcVMSgNuMZjUeSR6YeMgE78GWNlQIaNeFlx92jIb0AqewM7px6u+9uw+E7NTUYJB17DzX5aez
xVoNitJqFieGRgLE4pau23rgJmvxFw5UrPlPlONLfzhm0X9q7pwOfRj2g3mzSsHMQJNA0dhpZZ2K
sJg3UjjYtup83+FbgiHIBxKhgAbf6G5MiR4a7k+sOM5GEhC+IXx+WPisvZf5IAeiWgdD3qUpSI+J
dsBGNrR6ydCG6ND/3heUuY9+v1yyeX/m0YZQTT9eOkikqI2vuv4s7aNssa0AHiii4lBV+Qbdby+e
ZXaI85jW8XXhxMrLUSqO1zcz4psPLHurXVuT/c5n4Vac1s6tt/N5wySmhDSNQFEo25HT09UvWntf
d7WH+jxq92I0XtOZWfmAQywQ3JyWFWhEcR9KVVI5yGJ53hrZoIUrm6kal1D3FZ+cjDbV3OlVyD9a
+q69eBH0Tbd06xJ9wMWsJTHcRkwbuivsyxk2zzZGqJB2Ij70sUVere9t7CFEjyCRrkej/zwvsIIe
sFVaX7E7CIYwCrCWFxe5KDR4Yd7RFc1ljFghMpqi5dMiwebikhCJo1E3JPDrAzLGZnoZcXS5DzKM
StdNIszomDgJ30nzhqQLpPs0bUznGpASjdIWBhkIzo4nP7eroosJ3+4vdrB8VvSYCix2NbfSO9MA
3JxdSBwvAqLZSxgJlNEn2wKGK2dYd2rlZ/jTY3Uz9fSlHSBMZK5XUh46IIk9ZZOzTbZPwgroIxpo
XVcw+WC5ZYiUN550Vd4i3ImPPBjtd8hivwN1RfXu8IWZXbb7RL3TEMbaEZOgA8vMtsvmiGd0UaXh
kYWq9EdbY2twGpqGH90pbVIhIq1uiBzGRT5dWAWjpC579LOWDuEhbROR6rrglznrkQyCL3W1jGLB
MN++9t/EY84DhQ/GI5/BAyLEJCEGJLxASHj5K13K3kYMzVsrwNz4FT9T6SpiMJn+awslzdxoTO/6
TX9WEBlhotffFf5NHsRMkEW2IWU66KAaXTMDVRnEqvNdx2Pk4ArUFp6041c/qpIO7R5LV6QwlVzY
zwY8+ZS+m6B4FLvTZLSmeElD1Fff00Bpnf9De7AAuiY6Ow6JKUXXaCpAYQmJygDvcEcRG181OM5N
lLUj0LZr3n9QyMn4FW69DCRX5nCGhK9fXnwGU+KdWwFAjvGYzAV+ZfdR7fLnOOD83NEyrXM4KoWm
uEwI1yaEjBNUjR6XkVbDeg+ghmmU8gKaWMOkpoZKl+8SZkNuk0R2H3OBH25UWaI2gUuDO1xwOXOx
rwYZVseSMr7ykssTboJjcjx666dmEYXt/PjT+2/xIcbbsmBBKUzOWF5wTaWnfCVtsoziPpmrXIOn
uDxRzAhI8s3EKp8yKXqkVtFLK9I2o+0xQThr+3L/HqmShkh8EP0gEsfiyLrqbszyeMPPwmXwgBC0
R1pD4+UnXNsq3RYQkekNlhT6nIcCNnwq6D8n3+w3AAbqdbHTmwOSS7qge2MY/ltRds9MRlyKGvij
IkyOAgaU7yJI3USTjtGjeSdlhmCECivFOKNB0+HbRic4/M/MKvxZrR6yWwzWsw+Tfg7La6TBw4cC
67TZ7kbmaBsnOXIPrSl+YpafinQlfGYZcKmomlTlWht2y0bIfnWHCL1+eBIsfU64g0nA+lnOH/ef
JlQZYQRzh+pCTA2OzS3ik3PxHknwYq7FShn3aj222rJUldewXQvahE8qy8n4gLlInZSlO9YCtZqO
ZXIMunpjLkQj5/2e5mp1SsCVXiH5hLg2t9yBttTh1THCCJvbRCVlp+v0dbE7tov8A6++gexBV9Rh
x5FPRAIuB1CYtxshD2TXbNMhCwJj57LHcmFZEHHv446SyndBw50vygcVsFt/qltd/Xug2fwIS0Co
3dxsGU6toqwgIp+d6cN3w/xUOhG+I7+jAUATC28gTKUxJpEBvO5e0ApfVpo/aQPAcou8NcdLkwS5
CJhO/Jsb82Eo3iSAJAVHcQtpIFqBL7wJDWu+KNBk12HWLdXb1ZjTQTNJd2+1UTF/7gJq/kn1w4kK
q2Sd2MEj5ThkNElOqPvnC63hRAZbMM233CQKfFI81fxIYog386TRs4+qcqYIWTshdYxkjHnN9oko
+ND7EFCT97Xoueg5PPQWooN/DAjjwHYr8jO3ELndk7bo59yRJrBuh+YMgvLS+3M85R2KzwZpdI1V
m7M+/ixqcR/UlrGKuw2uaUTOPJdC6inzRIU1rX/6MC0pfwMoGUxumnBUI0Z2Uxg8MYOyScnD/y7U
ei+ISkNK49zoCRJqcsa7cx2YKWc8qHBHpwPFrlmHIkMRYmNi5B/MnLvC3zmXeckswkhDA5aGaonZ
lbg/gvmmjYr6UlHAmLSk6cD2Lw6BrHbbh1YXDFiz6c4lmTw9qLKE1zNJzEAV10icNtD32BsPIZJs
3qT6md42/tUvzllXFEE7v0Q2dRXFZqxIbMQsumS1E3GJKKIXVTpR+53ypDd1E7NQjFUrKDDQYfYZ
+PD9kIC8ircwbohynMqVOITtjpjQMDD5QMYnRi5naQOwo+zrlxQnPC8CY8F+AsulwpUbbzwcKDHb
e82O2zofwuI89ws5WOPG1TFXvZwJtC+wiYzKNuCuvNhY+uwiGc70c8SRVYCE4XNy5rytyQ/sBfxk
vkCVryu3HAp8AfWUPsxdowJL3h71FcHJJrENKcp7KPzSoDC74AX1QCDmBsLm74ay3ZA8tyS1b2oe
hzaAN6FUzU9WkgCisAaoy22DoLHwcN66SdmBv2hfODhoNq8CkwcM2DUeY57DLsJyHP1hx9FjJ3PI
JyhCqV7DF4z9qLELXwTdy/EerYAS5Dr6oMvDXym4LUshjOO1QT1VAvDSbvu2h5EKACcAAZfLZ+Nz
vIvqVpalJU5b2ww3OMsPlK9ao68qy3C+fzWXh5fnJw2YPsnSIau99fcbFnn8UXRXYPXWyEdO/Jgl
ocfjQRU/XYMnk9QMf1hD2bw26j74YYKkM2jyLRw9JTzW3yWNxt47P+OhYk4BVUsBmYwNqOc0SSq4
MEMyk7aaFBLZVvYlWU+Al+PCVsYMhvLWgIoeEOSAredx7Vc6rMzDx2s/MC82IV8WmWvLBqYy5/AU
AvGYe9NsHbtJt8pgk4DkBKfw21gSuw39SiGpY1R3enx5wlh+YB5uD48SWzA+Tbdc8t5/ZiWvqEA8
hxwBINtX/g9A9zYj/PfWJhKL0T/8VjTZCdQhkXDg5s/pJ0Q2PcxvShkC9v65/756mEtGJ6PI0R/g
d6rytaQJZLA8i4QKb3rBIrUH2Wg5h3JlKBqmHzFXtTvgZ7j5ZCVKRS6lEqXAe1f+jzVr4E81tBA8
gxTZXSKuYXiLlNtx6qpoay0gFnd9QNbTmnGQKnCrY6VHW25OZRpr8GkqAifC8MX/OVJRREXJXsLb
1A1jmtaYW2KPhN6Q60B8l6Zv6GGZOWQeL2DuLYpXchXP657Oul6cTIrYoGnTa2OBnfgBWbM90Z5R
xvYfi+qyaGwCQ9rIdy1396oLio29SUx5FZkxsqFVzxy5wiD1CDdAa7hcZ7S2ZP1wEGE20uv+KCnk
Zb9Fk4dMGLflao0cJ89eUOyQWFc1rjfVxZNl6LPzn4xYohh9XYCZVViyELW5jb+C8aG3zjH/xlmF
ZTZBij4ioE8o0aPJmU95OBWI9+/3ospYiKCSFbe5vJZoU8epv7lWP4IdwWX2Bpq/c11vgERfa8wz
DzZiaLm6iPZ2OaAq8DAmj7JVriFc3Pa8Y99zMj3mfEkF4VICUHElEGVJrfGByyBB9tgPbG3stKXM
mH4fjWRunGEL+Qd/UaPhx/8E2xHknb8tqbZY10WWpleUgrQsz1jU+VreXjsalRpeZ2sejUqD+oT2
OOBVIjj9jCbKuK5fNbtDk0fQE4Ep1gPO27UDTzPKdpCOlEBEb0g9XlVZxWcWy1z9hHkg6rhYOla+
IrK/Uq6CtzGbWFidMQI8u97vhdoV16nBiRwyDCrA9uU7mWET22lG/1inOhG1Xj4CID1i1nac17+W
A+v77lBVFXZiWy1/4i9h8wgdayyt6f6O6AM2DiZLXoMJ6wLSsPZ5ZgyQbJgjiOmDmOZaz+Z6pucx
C9Mj7GvcrtLkPYKjCad3GnCA53ECBz1Ot/Pxpz7YyUu65U696Zdq7WxGbCf02N7x605QOUjVurPD
yNz+x3jB+7+Jq+i/xZXw9bCHQXUxDkMUMcJrXpQWODVgvXfdozXJfH4J5CjdrXARsPEBesBjYYe/
Ds3WvbthqO+CGQCttkdMyaXZlqB5Wdp/+v39OvVRmd/Nrc3KV3wkX2YUcavRzk1hzfitrP9OR5Dw
4d8Bjb/A5X37xgC82O3rvG7C1KyWhbTlcAqySTrz3LNJlJEkpc0iivwde0vHeJwOU1+8HO1vkxZI
/fbLWvWok1p8yFbNPQQmssbrzzhhp6ZMIzYKK8AvI4KK1pwEvbGcAcBrKFpvWeTQ9RIa57EgGQo6
1P0OV7diStdnXDuBxImJ4Vo1mlPZkiI0qxgnALl74gRFpDsLw3vk7k/uGBls/U+zPxPZXLQJnBJz
BOLCdmX+OAorgfigF+7Qj3Lt6oZCrMldVrQDT1xE84e8V25Vgp1PUXlOQXv95o3R5gf1Y9MqTZ67
IoUUu8U45PvMYVQKT7rItta0SBJ5498anySN8PBZwyXQHyF0KKwcgibb6iwdNJss7c3U2/173z5U
w90hSE95StExIY77Ne80L3tJcxUhgk1RBreMto0y3jvcJ8EFQslQzM5OwWXeea4tq9l6qGPSVeN+
GSeG/D4zQ5d0rod0Po2SiiH0N1g0IP8YNvPDwCeO2A2CmJUP1UoqXEgWpqmxf0NUEt//FLNjV6rj
ccoyadvHhMAYbAHMdnpIoEHZjpzZTD0jlgSYhiGB/AJ8blw0yiyyxcp9YC5guF0uyRZw3NIzMTqM
V0ToEUJNKVUluQbDW5EL6G/VhvgRqkeApoHluNP6mz6Bpne9Vs7pDGxZunTnX/Qt8MTMYb0ozWzX
PdmKpSmjV8Cpg6bZKZjEf+bB21vRQedGNI8D3cDhdpr9tMmnZyWGcdKdrGVtDGz6Fsq/u58Qla4E
yixGFyE/At29O/Mb8Riat8R1y3gFIn4ce8+nmlmj3qwPmhio+6qR0N83d64IXlnnjsQRX879ytTy
751Ms1ucId6f46MdFVdPz8RGbpWTtgdkOJbODTVWVp3C/kUwi0lSxjTRGlkdyrNtA8Zti3W2mpzw
L+7Iuv13g0ksJ/0TZRYauzIjMgjAa+Th2gCVnyKM2RNHXpkVUJVN0QsDVI921ZFtYCrJe4/WPOTA
Rz2/tktnhPrvll/7Uk4+i6zSke8iFaUNh1KANLbX12ktPjXF/6bKbkIbB371XA7Xw0PYEL0YIu94
z9v9WgAvBtu/3ozX/LtfYEW248yld03/1zSccGkekGMWdGmytcwDljeD/oEz+AjGDbjSAdxQ40kj
hxY7zGedz/qAdSPonOuvt/3AKS4zN7GI7flXk8Bpr01wDNnz3cqgVBKcCjfIgCzzG90SYlPQ57za
MnMmVelYtugvN8InqQLi1/wk/MzfTX6oVh3CL+WHx5LqCI19u1WGZp7Qn6R+V4y8nRo9k4CUredU
w0ec7LlYfvmIXihq7Z4sp3IPTtbRPY6JG7LXKI2Ft+mUS9wGh9LbR354ZOmS0SZwev3cHY25TwZ+
Pm+fPf2tTdDuT+ForKnznVfdDVjK/ve2pzWxKNs8qy4vWHBf6cZIPKO7aevqKE8m4W2iTyazVC6a
nwVO5Dm8A+bDVtfnaR0a8CZu00CHjCPWPokEXvWqkTHZS4ZpZZ9s1eFlS4mRmpR3pAsh3N9xxyzV
eH/P7/B5P/BZD42yCcbbrIlDT5o2VFDAZUGLm6YoQDU6+/p7puAUmNaC8IDrgbEeKHtkEVZdW8Rd
38WkUPXOnJkkvDPWKYaAcK4NyO5rqi3H6EfojMy+s6r/0qOct7ygImtJpn/TneOk4qQx0ssi9ARw
elpoGMa07DVEmYYGp30+Yl9Y/nh3f5HEbONPpviV6Empcb7PL0h1kniFbvxI1JGPgEno8SZN17FZ
zgfwPJ9d4MSxhfXRltvt7jOXNudcA3rUEgPDnJ9sWhWe7srk7kEcpkm6goeVWKywFa2cwODssCmn
Hkyc5h9uMmo6seCWkWYIUCsnqlxOAqN2ZbLxR0PK1nxsdW+ajhfqYn1vjXuwK+bS3n6vazjYZ67w
W5XIdhR7RzUmkKOhVGlSKTsFcfxFrVN03/wLXjzDEWrJJpBp4ST6KgHwKKGAtpQ/EIYyiElQRivf
CbFWpCRnBCH0h31FvXcxbCBrOd4SiL1Enbfi6sD5sFq+HYBt40uxlpOXUVoEGObDC7PT0Q3vDM0/
4e+K1ptARSAZuV1bgKTZ8X4Z7FBOAcbQ3kKbC7Skfb7vc1ZLn5c74wMJj2+5iBkv+0pFfQHH8Xkf
hXRI9meofTLsCNwubYlcPzqjS1na4ajakZZloAhAK+tqx/g4hRppwil39EH82oJ2406HrLHFVm83
kTXljplG5aZ+BfWh4pX//qoMLgjHglenqLXCecamECuoazlVaphkdLF6uflrgSL8e5WqAB0nQ3rQ
+ESjWXmRkHznyLrHyXyV02E/QdsIRxu7mW8bqSdd8FX2zsVWjDd4mIJNhCM1OQiaPisDbBIBwCCm
er/i50i1XtcxXH8lzOLT6b7eouq7XGvn7EnxVZtF8+sDOPxZr0TeAMsW6yijZwWoLhROgCEr8BfQ
mZYuJDtZISL/2pAeRrIICQ63JZ+8x2ULrSzDL6aPpGSYiH/h83BQ1htohBW224L5+tHKbUXCZzWB
93Q4Q/6qyZFrJdjynt7p2Pn83B6seOLd6KdNMFkhQwxaOz+ACDj27tgfTPSw8Z7fDWsvMyQXd9jI
o1XZQCQJ+x/Y4hrw9oinSGAD/Zit0L4fS6+asbYJ4bMiPSRO7NQ3Maay61Mqi30UcTk3689GKdRd
dVlVebjMjyTyJ2g2xDSCvU2XJYriTQWKGDI5HSz01Rw6s8CIubqq6GkL+MG/RMhPVa4RBJpZLKKB
ZNYnI8H9ryxk+TLczlROcEh2SiwVKpfAptDfF5mfVoKuJGUH3E4EJgYbTRSHpQRHGdqBGFpmzJtM
nZxiX+EaNhzKD+c+alTGVFu0Qt274EFLXB+eojnZMibG9upE5ntefdOfe9fKa+XK7iv1ZJUKBNhq
F/HwpdwfSjRvwGJ88fk2cb8BNTYWWe15GtK3UDcjxowFEojaXNDoE1Mg/wBPwEoE1KB0a/hERgf8
fDSzH+MZIZAI5W0Lh9lggzWqWoSoF7Y/d2uE6lXsW7jPb63/tNTUWgsUSka7K608j6FpyJZtfePN
Bop97azZahj9XtwRyE4sixAtb4Ws0KBCHZYe3Q+Uorg13vHUoY1SXFhaUPQjLUSlyltTuCHqYtBq
h3d75oLHL3F5s20J+PPJ91kN0bFIHrpeltUuNKXTWXesibRFLm0GBoRvTNXpG0BF5Y1QGtKW3CeK
8FScpH2c+w2k7PfBf1fj1ZiE5QcOQ/VkHG7U1Mxh8KGyu4iD+k8ukGfi7qHz5DJUy6faWe/sW+1O
tn2Ryw3uxaEHS6SQR8IDs2gkTmgLsn38YyZHY5PNWZkWt0QQbydSvwiUFrosBZEykUvPDa/TBd7q
jSOBp4WbpFCWfWBkUfYQdtwSUFgxm/rU0+9osRBd5mt0KBLtdVe0ooVOf9Q+RuTIPI/8ngXXdspC
6y/QM+KPxxFpu5VTP086T2eKLxZGEDFhZHiLNbjUDH4bK8xIdolYvAardYpifUIM0BgxkH8tCbHp
daAWIflk+dYiv+GnkSRAeeyVa6OaTUVZ78upau2a8/CU3stgut9u68qiuo2GT0uNxs8kZ8aCNzpx
aD9ld3ncwo31L6q8JK6BSHVzTXsou0Cnne+lDR2XAYZ4iDT5sGXRv1o3oyOMD9ysLKkgt+sr8F5y
4LBdN9lO9ZWS55Ahs5YKWQC/zUcyu9We/bMAYyWsqgH+hLDGIAMAuvxIT4mDLKWmKJu3hF2uKDi7
cpG12aTzi1FNouS2Gs4jn0U5LjQ6T4mNYTsqZs+nDmUCs7/00LqyYRxOFWYNAhCfT2jqDVWKPRlX
nI5t/dAAwG75rFkvaTA2fkfHYlc6w7dm2fXvcYZrv5FdMCPBrJJmMaXUEBjniKZ611VvkQhmfsj8
nc2Rqx/+dqLIfjzalKdCCN6AsEo3h0OjjH2OziXV914oZ2t0N184uTihrS2OIwAHgopT030rNWEc
WGPGOaFrFQ+SRsZRNrBOYfFRec49Z+e00vYHyqF5n66cw4cr164u0bmtVOOiDalMVVu4/UVCsbPC
fIVJ99jYlv30KPcvrVWfQ5skX+YztirtXaEG3mOL2dz+nHy5m9UQf50o7HzUPKbxTKkTGIArWYfF
m7rF7R1qSuGNINJT6hbVaNm4VPOWActO3QcBaZboXywpN6iNqfUtXEW6GlRfYlNCsxB3xYzpzGR0
UCFk2LwrXiRzDZg8x6OKdOKH1CXIwsq8F4N9xomb8Nr3QJ96k2Vz9i4spP2tA4c9phE3WGrqkYSR
r5pNh3CQIQqdL2aXrx3Aqoy3hBMtIwcY3E7IqsKJB6wgYJSNlxNAqCKEOc2jcQAx/Eu5aCx5M2Vx
cbuLdVoOA6qZ3WrX2nL4SsLBR1V+MEZlC+tn3GE2H1mjsUoP+PlwozZDE4Bj58VzvSEAoDS/FFDB
hAXC1VjB8T6sFfIegO9mRjJeVdjWJOt8OymBmfJCkpL7r2x07qRtMhvSQMPaV4yZzAg1ivUxCBqT
YYz5WjJry8VVKlnZuHph3NZdUA6KeN+VSx4XBN1ql9ZbZDRVVIro/GNVfWVVHlRZVSWkNm+YINo1
gtJqEwIGs8TOJt5YBHn3QfqBNklPV7WjBXIAOualffMOipoXV0/NNpvqyyc2KsEutwMC5ZbfaFAC
jmtjXcqzXZ71LJo/pctqqnp8CzauufmwB4iTAf6zV3MJ5bxjaZoas4b7MS/26nL6ZAeJEyxncJDs
ToJEIZsYM5B2Se8fjGa3KyPoPrkTYW2++NqzKS5JThJXs2RhXuGEqj0PlwdgUg4L5tb7D7tK2QpU
7jFN2wrlum3N3MKgbG7EuAAwIoLVw6kOUhjHW2z0yrxgncMMG/D9wwJ3/DaIuOxwENqovHHJ0hYy
vfagtMs//EWbSzzchNwwMdWt4+7kpLt8/1vWMNn5ZaEZs7HfJ2I3GOp2nRILc1QiWX5BqgHVYZ4i
V2Q69gUjez/Nv0ZK4Nm0mkkZFvA7NANgmKT/Ku23J7CIrFT+7euKX0FU7CsBNvBLtoeEcN8OFaZb
eZ4Bu5HkqdMEnb5V3OXXLl4bh4tgu2jl42ReZz23gaZtjF3hiG4KT6zVz7KXO/Cop79k27wmlnmS
1xTtAqvq7bicVpgjZdPj1/NCGCzC8H/fHr1KAVBeqbbZa7EVgu9duE1sP8A5fIulfQQBjGYG6chx
PnS2OEMkul8VJ5dqX45LFfJ4MLwnXOkXHJ24nNiuWnpWUMFqXNHRo98TpixuZR5pbO6S7DELAii/
SdJK8g+x/UyCE+gfNT8to6FdyGRl2zRz/Dd5UnDeX3RvAV/v47+wwSAlKPha512wGmeIcs/pJC+f
Yst7rKcgPfbUKTc2CL+w7pVuwOo/bJVhqeNogvSSuEBkf+ibs4mNn6yxUybVooMT9ySXMbPFizFy
8hHiqVJ6kM4ZCuShL5f03B3XwWwREaYj+unuedlw1WgA6gWfZAiauoS4ytXj6sVEMUAv/3V+21AF
xc/vzAf8Kme8J3M0/Bee5pA2U377TeeaDVmmw9P/NKxTG6fF49qBgPJ/PfZNzAzrWq3KuDkpG6ZW
ayDwxIgugQ2DKtNuO6uldQrIYPmbH5oHbQiDvXhv/YIHsGETeCmoAft6vfgZ1pDc+I0slU0/cgaJ
Xm4013kfC6j7BQJ+0Z05e1dGg/ieDvaapeIkj8p83qyi9CFzQSuPeHk4MFD4mERjjmb2XdTE/PDh
2+3JYpnmf5uNgLNYqS/0OJeR3Z7P5upfBnTy+2Fmftvdzd3zYBUkINxk8fRp0wfgv+C/ueZqAI0A
yugOn5ZofVEGVoeDWwDMsLd+/j7R36ZhFmcV2rlmlDX0ebxmhHIeBG1Q559kfsla9A9QFzkKoc3l
IGgOBE6oXpgjNxmBPk499AnHXd8UFU2mfJnlpo378UweUhAE9YHEOUr53Lnt5M3DbNTizkb6FdCk
NszhZFVnWMpV04uvyKnJCxS7zN8W2E/CmlpYjOBTTnMoYTMyyj+DZWSOVl4rl0SVsw3agd/nmlos
DROBp7qMVEIaEeNNkb29b9oFWzSsy5etZ08iJaNuq0k+IRrKXdCRdOnqenN29XpAlg4cLDM6GKC7
G4FmNqrE1zpDo+PecWqjYuwZW9iOt4keGbruoUYJ0N0QMx9CkfQd/v0GKInH9k8I621GnSLr+KOU
4Cq+6nlqk3K8Y6Vx38C8DvxMdGYF7yUX2i0ZRuHBXDtSPHx1/LjsEWEWH1sGvxmC/nz8XqdqoxMf
QsEKLqa6pDGHnxy6SPEJRIIGP/aK4jw/Fo1qqUve0PnxB2NNBofNMKzmsoMrRY7gq2/ijH5DDWXl
SKo8o3Az7tPo/hKkSYdl5JnbW+m/Mg191fESj2HaYZF1/wl7L2cQgtuG9uLs954uU1kmDmxUOBQl
2D+sXlnObZLRSH+wdpdSMeLYDkGpPnrjuwpfzhpg3rNM+7jvvyvokiyYZNz9Ypk5ZmpIxDaGMBb+
PW7H+WPwfy4WzjBla12P4rZyd0C+T23A7s9oHjX6YmvO6oSfNnjqir72Wd8KhmpcgE7fl0k0HIwo
/EzNsxpdmTeEA0IMF1tjsLbU2MFxhyOX1o6ltDygkPIQFXoBnStmVLC2K/0zG78nJ3k3M95u5mAo
wB8yRv7xTF5D8yWC13Y3EsEQd9A8PDIx47+m7ksLP3e+RzqqK435Qq+jNfyqS8AXN46MAW42f7Cg
PCHQqNtagD9sXLclrWCapPLT/jCGjegS0V8xCyfoJV3fvd31dGA7Fph04bgBnr6ono7zzbff495x
G97vKmroYuBxXCSFn+q4D0yl3yXpH+WlBmWMSFrw7+Wsmy7xVnOJrbYLXs3SKEmSWdHwlWsUGRNa
XN+Ex3zmlEq8zETcc3VRZt6XLJw2DMuXmj/6kzlVDSwryskZ/9eOPl8O+ir8a2lpzhd1Zv9eAFlq
3Y5Jtz4KyQXwjMmxGecMoN60a2ansB2uovwZDmMRSO5xiqNKm7OWKrNZFsJKe05/1sBVBtKNP5JY
qYQclSaBFElq8DfefqJYq7/V1vu2324DvL4yXW/aBqXT/eLT38ZGoNl8z1UFFykRWlO+ZpVn0iqT
28T49aLeZCgrN2Fkdv1dL9q+7M0sBEcSHMJKNTu39YBkwpw/ptYmWfr2FbMzhZ2TEweaodKN55q8
pTWWigC9b+zmSgc6NaB+MFuAUm98IjY8ocShWYEVdmoYD9QOofP/0TSSh073aBEwWNmCHzA5Mgfe
1hBiCn/p267uwOtMXuOmb9ZGc4/4SYGquwu+IjqbAcM17ICP/MOlRVbB767r3r9zBknZ5ONCfXvt
uYvFlbqLeEjmmkwPmNNMRomwCSrfv0+9i93nwaDieKb9TbXrroojVobcNpiUtK9l0CfX/WkhuuII
ETYpFu75UgZDhbht5Jvxe0cv5nZmv5jqqq9tAToqpjcprO4ZFGQtMvuax8v501CiSlChNiDTec1G
vKL2uQDdM3toS6o5ICUBMzmwIl9tLzOVP0C8RovHeMNW8hhtVITRvXz1EpEFs6JSKc01Fqpi/d9s
mLL3YnfMQVgfr7wL8AYdpEuGL+nuQxVY1ixiEbJ//mDw2Y9S8lAkia1wJwJvRBP4h6IoZnyi6ZFt
d5UudynEkxeDd12WqhbfqWtHMHToot5OP7vIYvzezAPUVf/cWM/Fc4vJrFpd2J0uEQI72yuJYKTi
W74SWVlBz7l94B+xzltQfb8bWrR1E0ebu7h32Z17VmLxRrGesK4UKPlRmuY9yeKLDizp7Y5I/fG1
PnPYE5d2w3hFQ6VJ9EFGD1WfqUmHcnMnjXt56LofLbg7XskNxtuncO5G/LGeVFdfDnQh7+3Ip3LN
afa+Cegq8iIgQG1AJLlMVDyBeqK69l7nJdTb+ydqEKMV1vHg2nNB7zGEyCx9u131Crfgb6pp5w/U
LiF7MGgEHNNgkG3zFXbF+lXN3cXFEKe6l1Dh8SxjQ1W7jtAqJzam1x+/moax6OZvn0kpb0tqCo+D
ZuP4IvV9ouvNlspjEAqh1AzkkNT4PDklPLq1lkvcgot1AjqtDqH3dxcwa2Sfx8WhTIBEHG/pkIF6
so0H4As1ljUBykj8bT6KYk1crTpVBzDH2XdUh70XX+ZO/Rx0++8a2J5HVqAFJb1HaABPwGWEkLwa
01NbxkdsK3Q0bqWc6tEVgLIJmf9PoWCt2OXOTrtchfeW8ZOEJO/IH1obnhsSsyyw25GIxrksx9s7
wq4cqKj6jZzzy1/f13DQphNX2LCo4A23n0YbY5LLIw/j1c+Nqa5N86/+hAFI6e/xx7RKQdLCJrpR
aSXwE41BciwZWYL0SznjmfHe2dGOJJ74nbNZfzpWFrM/Vo7e0o+98ES7vsJBdD640fHXRMqTDI1B
+zZwfHcc6vP+9ogRqaQ8wRtN/mxC+77HaGO4k/Rf7fZbc1QJtgF1qNrYd+WDA85tfaPFkQ4NqxNX
TefWJ3K29S0xry4Cq1RmFRstAR9GFki1dz2m9reqBY4FphkZqk3X+npXhiCp7sPSIJGwYN/pFeTa
tSARkjXbS1Y/qT/B+1DrAkLCvWr7XuXx30CGxBBzLK/a8YGKXUN6SKbPS9fsYMcWEHdg40RqaXcW
GP4+nSwVhsWeSYOdNwf8HZCd2KJ1iT9GNaZ0qZS+1l5ZDZ2kHY0nv5iJ4QqkXAXN4ptsy5CVeHg4
4vgQiveO9L86bFiGVy7JEVaXr7JR/ERpvEexd83xkbDd/e9vkjccsOyyGtjFTTYU6pe0B0WJ4Xbt
AYkPrf+BVcgYVTv4CrzUwqeQH9Gt0YaED/+L19DqMI8UrLhtboUVq77od5VOzTBQjmU2oZpi7YG7
JHNtMGe5WvNhxicDGwdWgiJp2zrHNrQTuLvzjfiTHL3GMBXTV3S7n2vHap1DLTpGhm/44bVwfknX
XRcYzSoK9Ww/iIr3iPQSpwbtXJODY2SlCUSW+7WxuwDb6TtGnqZH2mXsh3DCo8HMpXd+eYq9Ae4m
VuiXRGT8/kZNZ0YPbCmy5lc49fUiGp02O4D7JCT8mLPzOJG2y4/VIGVQSrlhCo1d5eM5K8X70Srd
huzT6W3YCEaFk6m43pcTlsLkAO2MdOMLzK9i8KNgTU53JS4USd4ApP9oVRNvPmcM4XSy6Ixuw5hy
WSDaJ0ivyJMK/yOQEOyxhWmERZsKxvJISC5Bm7IlxNrEy2+2Mm5S3UkSEtpqknHLf5FsHHgW8L2Y
au4WinOaSpQySL3W0iARUXM/L22UwU1nGleqrGIDvY4q6EPErLIVEQCZSo2+K9Y2TZaIuMnG0MhG
4pPvzC5I43xX+hBL45qT3NxIWoHwnP5uii9rU+9/L+Jd2z45Tp6+E7CP4XhqFRgbvL2YmKseLdGZ
Btqe+47AaOZGngPSkSYT8NBf3KLqBsW+Iu8qxqDW58zAEIKfyDU50QI3Drhy0jq/+dBCNygJq3Tv
rhAH15X+RpVY5LYNjUf8/6es4XM4GcwIyRsihIVZVaE5j2F6ZnRfplYaiUzk45b11O11exBRHNyB
HDuoZZNjPTkDB6ZP+O932GVEaF/0o0PNTYokcXvLdcXjaqFbtnbM5w5I1ntWUBrt4iJv5XhHWxE6
Tw4bAZft92ok6UP7VX5s6uf7yi7JlrUiyMkeQu7dDdto9C/IebpEGX/wgSxrqnrpyXpBmiq/0YfK
YX3DYser5M8J+UDfuwK2yys+6OkrAiQ8bzU0To1jxeb9QIRYd/fQ/TQxrMf5AdcAuAvug0tDxUSz
rdA37+T4y3Pw2tIgz+0RZeECtmzIkKZnguMETrrKbln8MfR/YMw/vTyN4+OALx1U6pVCSjyM6Aqz
GZProDtPUVMmxrTOZzSqmXGXh8COfvXxDEum4qHx/FgZjOeYw2swg/1kpW4keOAaavwBurol0MVw
ZYgx1WRdNuSSyZa23+x83FCLif36TzY1fAsV0Npf6AO37HzpbFcQllbWEaJ811nDcsvgCTaQIqey
iQZvvj2K7ZskcEkN8/1+5OFPOO16kQP4WMrdbAn5MSzjYIelhmLOpC1D0HIPwGdufiqGMoVyC5sn
EYAisKzI6KVMijKdekBaccOHGdxnKFKtzHQADc4CQINU9xZ+noavSMCJ/s9p/5+53CJ/BIOKC4ch
cPUUK5Ms/4Q0wvbwNY+k/4g9oe6kQaKJ1o74BSHN6SNls1z1AfHchuLvPt2qx3kvRiHX8RvKeCfq
XhN2jC5CSFGKcc/lgxRC+WQ1Lx1db9GIkbGdBoIDGAsqQwdY3CLfN0fERPu+i4+Q/GAeFeiV+FHU
A4ogtzTRFYbE5Y92o5LyJazTvYV6tnGIIVF/jhqtSgqiuZq+Iaz9JS/QK+Wf3TbgWrF8DRM3XhJb
H1rPK97hyE2gFI43Vby/qy65UvvY1gLgkWxXH8/+D+MvxQSXLsrJ/tDDNZkGnSUM/r8gYU//W219
EsT8gefoGwo3SqXkUgPZdRY+eyz7czS29KmB3DCenG+5Yk9hhIqtwBZHBZP3vfp5L7ZZ8wj4PU8y
UXmQxRy1QrpFpu+NE/PAWVq+wyl0nFpTKmZaMTJDXhcMrPm4oXpc+h6Qnjk6KgvRjRFr9o2Q4JkK
bAono4K69nFn0sYTfR6a12sdWHf2zW+LH47e5V9Jn/hXARw5+y5Tt48h2M61Dw34clqBoAqIkQfz
mAU2HxhOdsPDfNH/L3VdB5QVyHSJFHYdxkkcK7sD24q6lxg2yDklUb3mmZ+0kBL7sEP5axcGb9N0
ACjSWjKKYBEV+n6JgtCV5reaPSEEi11tYCFD9i0e8sasDITLkOsM3nfD76omLpD4tbFUOEDBHqs6
fRLM4bnRpbPQR3cGIHM3YXIJw7mv0m/khkMzSGuUBehL2Hurvf2MIoU4OIZG7rSAKFHzXxhdvKVv
2SKMElvi4HaW9KgX89jb+SCTMgz9dzU2zYdsI8Z8kP+a5AoxoGxXrqaCw08HKe9/lJ5Xo5NU+mTZ
VHbLIHA9eEOR7MT47Tt/JGxjBnNKq9DuXL0gp6j1w/aKCAoNlGccEG5XZG7zZAt9EexOguSCEcwG
237nW6xnAHxWicOiST9RoTvtkXMPt6sDentV9IsTCJ87GQWvUv3wPUaI3JnKOOOyRda+Q2hen4uY
bRJMgfBtMzKe7zhEM7rV+omgt4Q+xGtCaEeEiZKMEQXNIFaTPy/8kbpATOA6hVNChG/oM9ZR8Y7f
q+8WMUmyuffWVRJgsLNhXfgSr5jpM9npaZhoLycSX3ZytaNmDfek3BtgypC0qMovszThQncrAyBE
dYB11IIMBQfBazqM3O5Agxw6pLrewkePNcYZPlq0CbGltgxrN9yE/4M8daILdZr48YsE2k1Jw6lO
A6EiyCs2trsPaXVxbQ2fGC0c4R82zwtG4tJp+6CW61bmVmvH4AJVulf0k3CU5mIcRF7DVK7s4D2p
NOw7mF4+Tq/VA6QUpEt3bQXr1Y0l2MEnm/KCly8yiv7d6lNy5gpVY33GT879LxT88iVlZbVNE8Rv
MCa4/WNA6G0JL2GvWPaDsAmLSVWnbIMhGirqSjbK/MTlrDmTVaarQOrdXP0zrUfygUaYjo+khEAI
X7Muxzuy8R/035KtBkQa0jY2IUwtkCsaGIZkRhynQcULZ7HClvNFnx/ky+3hffkvDFXoTseqUaox
acHkcLnlbw0OEWaMclq5qFvhc8g5Ztb0vDI1p5mDOGDAzmYMLUZBTNLfOiHk7f/9sw//sZ7pYh4z
zmdatWWHXlJoQ63aC+ovNIJcQvQCF7McpSJ5kdCTwzMm54kwDt/HwI4OQ47SVMKb+oYQkI3na9cM
9efMEKuQrY1jlbBy00YiS1sx0pC+7JCv0wx6m45YpErWnD5rYdut31RTKwdXt2qSbaSZKblojy9P
mPKODbzVQsT59s2CZNTE4sPG7l/y8sRpViDZAhbGzP4RKVhhiq0lXp/VZcX/HPMnZRg+4iMQfczV
kHI+4arhPuK46oICDfJnIkZtRL0JDI21krVmDrkRfA9efljvm5xn5uPcWnFlhOk0o4Y1A4gQdkTY
mhyEYb22xDMIpPr0HS/lLrNdv+F9zYdsZ4JGmEH+p9LrCQ729zYNB+Ad0SdifiQvs4TeN2KlvvCR
XgGye/JJcmmiC9ownrF/xyY1QweeSSCl5aYpFIdTWN/Cvl5yp8a+8Iok4hsMyZjzmzuFCHoYHWUZ
/cN2EjeGJeSUO/PZwv6R7kqLQR12eXXLCXucDivcswsfgGtV+ODR3SmkORhJwVc3QOKmZMvl1Pvq
rLNt0pLFTPYQbGKqnIA+1ahGZLEpQXkWUhZjB8sqY1pxt9q2V3mJfd3WH8tk3YAfs1lJQQ5D6Bho
a2M/y6C/1vJfAyO9ICeLecjSg7R6WHprQeLuwGRblDGtOeU8+88pZPB6XCRwHjkA7i1tGtvpm9aG
0DbDghPcY2TLMuHeI85IQij0SaFyv4P9Gfe57jEVdm3wRRDGAlXLegoRlYrMyn3MNsPljVc2Sxd+
Zhtse4f/8kuN1uV/pdo0WJrs0CA+SB7H9GTOGRhgcozeHzz7GKp87jKKnjEbIPRnD5r9eFG5daKD
b4zJlN0tM7F/wa+mkTH5Sn1dhZuNshvhbWxo7WeyS9QIeEcXufdkuQwcgQk+PQ3oyhKpfG3c4l3P
ivIjz3gKJezDHC1QB9uhZ9xLzY6gSs+BQaRsWST5cXdK3KZLAYkhTUWswH4u9SdDyO+pCAYlrqtP
boTesyTVsw1V7zYIinvTCw51wDfQgVBuPmZ+qQ84g1EzwmC+Q7mXUFVAL4xNEnyW4h+vzqZ8jNRg
x4ITu02cRJs5xQbP3oP2i4G/IV7aOThQdc5O/LaxRGpPSEB9qk32uBh51IqkUg+Eiv0GbZj4ozNC
BSwB+USMuR+BUhqdxQRHtTKCdmIqsPCURLknS/l0eR3dB4reaMM6LNYgKnnlYxlTjxT2p/ZlPhjQ
foZLyAJVBNY+VYqkWFKZhqpKvgnQ0jWVflYQbHg7faUqmdEzpl1l8/9/eNuRTxYush7eJOcCx1f1
rmDippD6WGGPAiwVaG0k2DpsWfN2ygVCmBIerQX6+9++Ct6etxm29wtQmAh/Z7p5nL1l/RSNy+QK
w8M55HUzSzsR72hzxApzTrxRrCk08c8LRRHjZ0JfU1zqzSyHtIgxHgZd7Kd30FI7hEWAVbV+IqgM
3fz/+TeJUa2vO4GD8zs6GbNDsKjQxNtUSda1vS0Y/Wpc7vWJs0dPZlbAsuAAf2zIWxsN4EKv72xT
2OodIrGyrRaQH2Kcpqmr8Q6guABYVN5Bk4IMRIY2AASJZ1TsPz9q5+uWKOXMga4582G24TBeJ5pM
+/hNPLuVnam41PcJeOd8lLWUtvZxqR5qR1QA2W1PCjxQsWSpOTNOuhQHzMKSI1ROUsj5Vqo8Jcu0
u4rucwHCrmSQjZUtopnGcNTSoDhenugmfxwjNzZws4Mc5+W9Yc0nxrz1SyrkZ+7h4Yq6pLZ4J37B
uUo39feRjXwXmOxUimzOiHzXHA6it5prJujzVV31mjplrb1VAZ/7glk8LtekR63MDlqHb7Ts7VJJ
KpKGJte0l/VHVzhmix3q/i1GQCymKANiyQvV2bOuOclPAmKkXRgRDPee8oWBaK8sjNw+/DJifYZA
VyI4n1j0rHW1lVHFhKhORNNTKJFopKaVYCcyR9onuYbm5rQJxDRdPsLDVxCGRD1bIHp5vGQQduQn
zprr/BjZN2MJXX7E3l1S2VRcEMIVENMzUvsEL/NdTQdLN73tnPduJepz1obdZPK3kz3QYzyNEUl4
w+qKlPoNy2OGwoS9alx+iW70t8OgzZsh4Ce2nn/hEfjDipG87BxgH3LYF9sQp3e/UzQhrWcQ5cUj
HwH8cK9nkuYQFGiBvjFuwnLFKnhlPpWc41DSArtrKRqJ58ACVoYd9CwJeiDRWDMdFbbNyw3e3JQT
k/Mx40KLPrzev4pgyw8UpJFtG2LmBpSCC+kA8Vz4dE/X4IkpFIGztJfP1th2dsWPSKtidyvxcVkf
1THIJps96M4S/lIe85noKOy16cViaR78qS5cdxWAJ0DmttxS3G8jKq7Nn2GrxITAahlN0mP3xfPB
O7NVNFDbHUvRWNZE8u445U6S8+b9RZ0sUJvo6fN3G8y3Yn0AJAC7+uh5WmEnt8H+HEoHM4TtjQ2D
agJmtjHNXgUVu9tmHEGq+18GLcHOMpuKvpQzE3zy1JVh8qBfjcbGJqiIqsPYxGCq/gwSPIrxn/nv
zAoeDNR0o61y8nnC53YZCEnXTlc1kvSXU1jI8gHnTmkn4cKHwICVeNbeL5iT1/JjD8tfxb066Ko7
AyXJIvUNJE1iir+fj48sUKBu2IRS6dg6D9becTK/LgyCOMDO5XStEeInqIpSmmF0Int5W+TiiC9F
12PqBpkkRW6fBkyEDA4bRiKluF507rUIX64eqAX0iNQjvpFum9H0cL2NuEaQaSOnWpnQLkZkeipz
wgX1U2Svj+UsIGdV7C0ggT2z87SRlc8XflPnKR7QA4VqqA0pELMsKW/IoHL4O1xAX7OOctN+0XdK
Nl7/mjDI5q64uKDyKNK7m+UpqASskeAQC3rn88rdCdGBHiIw/qvIpRXv4pL90IiBuh0mzBJiocAO
N70FgcvEClvlmtVcUKJ5dbv/w8i9JWsOCD7/s+DwH18R+AfYw0LAUM7ZMouca+C+uBY5t1zDOvxE
lfyKQhqsVkNMx+7mKbMxXzTWYKbtgZwAyghOAfLKLZ16udEZEq0pIlPl+2ovRZdSMYD9DmQV4JXf
ig7nwnnVmoJHQiQRR8653byp+7jE0bsErjCvOEYeCEXnxLx4FQ5uSdkuG9pLpWwskvT4H2082xJM
gGVS6cnbR6Ii64Yg2vA+EkEqbacBnPAmiPFdBmH93ySAuyj9hitU2EX4SW21mBma4Rl1fXeaHzcv
91H18NgowEkZQucc26EBliPvNQfTqzIYmuRfKEiU2I3BG0KJmtYpHsyzH6aRuQcgXJdBX1d+x8L6
TzGV9YVKA1ugIC2YIa76exUrkFHN/D2onSQjvesCBp0PyyYeGgk+Fw+0ivFJPtiEKrc9JzG7ilUP
1OvU/ExhbifQxD4cIpBWYWp0etSmbXplhfaXttf+MiNsCSpO5hrPjSybz7+LsVztkkp4z8a0P0oi
0jtj6Ab6n2GITfmAcLsiEb9Z/1Px/Tc3ETcn31jBcljMtVQQe7PI8EWc7eH0lUfwbjVu2XZ/ciGM
HJC75L4g9ndp6VdCanU6qxz1VuTPr2w0ZMkqCNtAUlPJJ7R2kCRxjC17MVTj0mUbYzGFkQ2KUpdy
yhxs6vlZgHKrlc2Hc1EUEEFsqesZbXMFBn+5kURrvjtb/ys7meRk7tHv7Wyn5S8BL0ELrzA9Q/7p
qDQrZA/W/eW4pK4LrwyJzs/pyVIRK0a7CdTGMKCAohJQIq5Rz7e41BA6+LlGmlXxDshPB5v0b6T0
qMN2REfxukiHNw0q+D2y6v9BDQyjYn1jC5qMftGWVfZ4nF3GDFv8RZwiw9HdPAwIMwkglnRgrJV0
R+qDS79BN5L+PCB1xV972+J4Y7/sB7FoDlURNfnw/DZ+sdF5iXwoRRg4FslrZlqcavgcYEmSvILY
65ilcX44bQuYzOgpwGRjtkbDrH2S17UvmfgzuvyLjNHf2NRyqBG1ckaK1EgrClDVJ/1RJH6npUKw
V/XangeU+ezyoChgaO7ebYw6jKBfLWDSqsMEyqhs0Xq0WKRZCE/4/vVRvP5p44Vwt6OSj1+3gFvT
1xichmZc9yp9zBXB3OMwm7NjIRybM2Fg6TZkfkDjiRSJZM3XjBXG+DSQYn31HKI2kR403IsVWiOR
mvwlf0vdNWEZfIiY6o/W9wsBvQipYQY5IZNFcWBJFE9IFsb8QLsPQxCNk/IKTmuixCFBW4qH4GpE
RU0d7nncIMe8Nj9UVLRCRAui4ug7vgYGLyTivMtwRt70ancWYpjRiFZy41SMLz/i0W3fgwcTc0CK
Iw1QnOi/IE/lxyoVN5NmQlFNED87L/Rm71MDsSKUfqtQl0se6cFse1ic+Pjnd8GVRyPICsHELR4b
ChPeUcOu1OmUcTkJRkM/V9UuLX6msx+hpfT8kICYcHXx0KtzzU66fB9NcQwlQNZ7/ffvjaN7/git
1m+effwPLDuUAElq2Z8ZyyZF4u2t1s2FRI4bVGt3fxBFmpE4WcKfCvLAj8sYsjVNl1VB3e5kN5no
Q1FMFHY1yfvxkYDj7zvIqBtrWlQpQCRtMpzwfnLGgbFDOuBwZu/MwcOxKQzEvK+FBm5EE0MLg01O
jS93I/8bULUOYdQEaKCWncbXSxXzYbW0OnUx+uJ11FM29pFQTr7VKZ/cP8SRGR0OxgkTFnIiIPaR
tl2UNzASs198j7hfFV7gYEy2Fpg+Ju4Q1U/+DJ2X/yh30fr+85VVpXoAOvU4awXoIBKVRBNZKnHq
jsn5nQZonk9VcocIdmin7Twda3cddC8J2Frvx5/aqJGxwepKg+vhlpnLiluTLIsMwvqFCBCLzO4O
8meviTCeMxr+PLaEHBFbgMyXj4kmB3auj7BfXOAFqj9Zqcz6Mb9MGy1wGMVUaLcsDJOuGG57w4hc
5D08EZPahikqdl3Pc5egjWBsgfdhxTHbhRdFFAPfHihNIUyYsh1Kg5i62hFlUNmmruhlDofw2LdR
nEf06Ys1VPP/3hdLnCSRpcAo60YlLX2wCv2/Y+Hlc0Pps2CWj6pNumqPAP0Bl6gGwjmetminazJU
N9xkF1ddy8tNst0HXWbdsDrKRxmAGzq8jb0qwDwdQgAaJzUXc4IAVOVKGSv56f8irte9zrkejAEC
g2D3H1JH2WAtsymlcfLuHTk8/glWKKzbYvyDHk5ERlq/oOgXlSt+RnErwxDfDEcRgodxJPnkS1w1
0lKdjiNXaiYoMZVJK2CrsB49DSSBMWD41AuXZKI/NhwJK46HOJXVONIuOBIk8EaQZtZ+8Huf09xA
yJZKTahCOuOoWKnBIJzoLWuahCgbgl8deQTJjkQ+unkSjqXHkJ+ozRklRlC/ap36FOZ4+HbvvLcC
8zBTZq9RZ/YYhNmS2R37hK4en9T3wbqffNNIGjg0nZOaeLARqxuFrbkXDgMYlEdmYEVSuKvRItZe
+NCNl9sUypsRFxVXTB4nmZ8fOFmfRyPVJGW4BLh4JmnS2D0WfAX9ID1rwfWTEZ1v0V7pKb6m3GWZ
jQvTzl2Z07IxVKC8HtTxXelaF/kR3vvE5yaFj6M+vN0PyAR6rnTkAoHF51adOIyOKUB51/Kuf+7n
LmXFJSyAJwzwYymZoPLsXVJvypvvSxheB/s9RzCKS/tdzziABNsZmvbpGHSu7iWIU0bwj+F2bqig
SaJ2P8ndzT3Ek84o+xw9f8nR4Vc7MLJXAof6BvdQlILHABytPqyLaHiUdwQqwo7dOTajVwfIHKgn
kvpmIcQaQVmuX5PAysgB4bMfHV8P/6Pgoj7g5KeoQISU5igfLrvhCSqDIRauz5sgUJdok2tDEGJh
xQnrLikw6oG7d2YB9bHGXzAuB6emyRA4NdwPW5XqcMfmxQ/f/DtcqLbzr8PzrR6OYt9+zFkUl/Oc
s1gfq4rMdrg2kAPhH6YnVwkkO5AZ9Ly7EBDfvOYPZanf4lZTB063PRmUZDfjBM/smq9/pA4y4cS4
qgJmeb5RsvUx1mFf72wmzVO2t/4T4kODDM1VPQDXv2QhG/r5M8P8/3IE3FOKb51oDotj7l2/3k3A
vCSd6NW/qK1TH8d7qgZEummrQYXAZSFC/lkx1rYK3GfGCwmxYUriBgEYYCpq8ln3iAael/Fi51QK
TSUZ0Qmwb7C6GF8CwYGIsC9siLSQGFzr7C67QjafK2vcjr4MA8hU54/Hs6cMuNBKhRI75o18eHee
Q7Q4xN46xGX+xUlPzdhedkZ2KxZYkaRd0eU41S2NUSwkadLFmrF8jCD/tJXru700ghIKaEX4/YGt
KUhbSRobbcm3iONDYmqU4QAqlLKPydF62eQ+D+zLJW87rNs8v5KNmvBDCMYoUlBZfxekr7vux/35
iIkwAmaMBW4e4bdvRR596QKGi3VTs6AViBj/kX5BFMcf3OlU1xMct7mB6XiAQYP7v/iGlZUM5rVH
Q3BNU4WaTzpKfXZQDeqitC2qADJvmRXCdic2hw/q6EVCN3dy3N162GnucnN+EJ1pEIgj/CVvGHVP
rPwzkSHPVL+TNBN9S7+jBA5Fk/aGzXvpSuhlY84PIn3jilmMKHuOn59cQgrWm920tisU5/7Hudn2
M40DVsY8sHHyZLfASmtLKNeX4PD/vsw92ayKB8bTnAEjDJqZGXzvApgrG5qxrnavgP4OrQSmKYea
JFBONBbPHjDhojd6ZPihT1zmyqBxNWlpa11Bn0rwcg5Zr7SiIDLhPc+0CAUsVuKVyAiqP9reKzxk
3OeXqKPZyoIYqX8wxrr9L1ddTUu/GqxFbCSsX+hIwmWyzR8Ko8V3YMg42uUnW0YHrIbISKVdF7R+
UsyDy7q/gD4fJL8RU71K5J+D0/Kh+XJ2xAmZRklETtoYAZC2p40yiEcI0CkJk9NHZbkKuhZSIfdb
I1eR5A0i+9jgISzJy+ag2LYmN4Q9douejOVL/tDOQJVzxOFPzt6GlwAE/jiFIsCKS8xykqPddS6v
7WxaPM2m43GIgDe7KY1bcXEDUdDwpOpARZdgPkKwy6WWQ0o8aaPt1ZkOMt3aaq4EuL7VkOmJ3BQc
MYpQJrLvF5P8HEZOPfE8QpgWqZEwR2R2EJxIkNFjqTYje2YMT8xa9y/sfxiuk/gWMMxuJElCdIZY
PNUZHwHwCOEm0kMYMB3qLxEOGJeUcgFtELrsUPIUegMHQAle/r3y89xAVpgMeB2K4Ouz+yRepwJF
NfAzmS7KLMhieaYbHUL6ROFAEUeNoXxYNRipfkzZa5iVVcnZkn9CCtJ53f/nCAesrK8ZJxCfYPas
0sOPgshLyZ8Ktn2VImvEN2tM93OYalOuPCf/t/Ulx0dpG0f/9/s90MX9482ZvMx33bZ2ffGVeIXz
jI11SsNGDH5o5LKxH4fBDxE5kzvszmdNYIVbPiNqbzzw5m0lxA0/dOkKdIcpMr3ufUjMy0JzDlvR
8joMD5K8GMpObOmOngesiUwJIJBwo/KkcJQT1HpVpnkdxytIv2OLLMyKE/Jahh01MKHfdpDqpKZ/
nsWxM1fBjdZtfEwkUvoZo622gLb03rEuwhc4U5/e8j2/xuWRT9y1X/yn1xsFdlpnez9+Eq9l0x+K
qLeyGvBmthU+B01uVumuyuF4txc+Gu2T5JPSYe2p3BErhC8qmiUh9sUSZn6hVXfjhkbdOkmlZsjX
WZSdrf9tETXwF2OCfw0sZznhYmJXv3JhBTgnGnDNoFfYKBMq/gK5uqarZvk7LUHnjw/zEDQMzGVv
wRByUFmZzuBZ4OGOUlzrzl/pxOUVqVlSCBz9z9QpysT9zB4ZJCtGUf8EBAy7IBpGft0C1Qpx1BCr
KnZC0mJ/+iUB0zO4vC2A5KVcMPbKhefRkR7BKKBsdwQ9xRZdYx6sYSSEtie2O52uBF9n8JOUA1fp
kDBRRom7p9yiGNUf86PBwYULVRKVQ5u4Jv1JE9EXVYr0pd8Ose7PNYM+k0l5aEAtxf5s4lRGFM0X
qnYbDf+cFCHXOauAHQTHqgfTY8m6ywI1F267AFzER38Vj30qyL2gc7CS6oMFc/2C/gVq1ruaBJ0N
qRpofMmtP6e4uFWAgcbR+A3VWsVDSmsZ7EhWs+gs+mg3KNi731U0dljY/lPdyQ5l9FRcXyCn598z
Vf2qbluSK77tCvVw4gIBC0184I+avQWxtme9s5d10u9U/o6isNID5oLugM0gdxIugDXL+aWnpYuy
3g9GwWVmf9HRJblc3RixKPQP1uEhO5K+WdVhaafqzTXsv0C6VbJsir4rNb3MMWlxjjhjM4TaNp+v
Ov+hIqZDw6yUUNQAzGxdWpAEje4GgGvKgFtQfSCTYn1yCT0U/IMEjp7s0LmEx7VZw5cPOzbRHdca
qPwB/86engxrV1tkioNw3UotvBrsH1/lGxuRyF5ZaRtg4DYGliL9THEpWu/CSJeivbjNsTbfpO4M
NhggFmyuXI0m9WRZ8ANwL6vbmXnQPWrePTjfdfTIRtkZ4SyQUsAJ5zPiG04+V7TXyAOsxjcifD8X
mezh4opdbRq+W8eRViLyFdbEcckqGz0Jy6K4kHERXuWeoWdddbKJyY8/IZSBOiQwtizm0ymBnqC1
3lqyhGS0zJX3pB3U41S5iE4dZm1s8/CtbNskHiHQSIhGTRDjrzDTrQmk8QC7xW1n446sdQ1HQzv+
DkDEqZ7ca3d7WWfXYUNfPlVtsKQUSlkytbdyRvKPgaw2MeucCaquIAwXlhYaMamNE/azq55v6vUb
4w8Wo1tIVbRz2M7KxSK6wYoDN7O3N+Tge0/aX348BrYh4rSjxHGSsUYRVTq0tRcWJkUYQXloixPt
OWbIHfVYfthl2aJ2cCQUJYdcsug4plmVM5QgFPWgyKR/tXUsiIRXqs13oR+hPygQaCY4vl1he3Bx
iCig+Q9YzvvoDT5vK5uV+dAbiiVyLSmkI9sh4o0EqCFXTwlpXWjAmpmAYOqUq0rYgaToT/iupXKM
oAVc4UATp7mHfMiXwep5hGDkZXZVS+RANFptA8re7aqWIj51Xz5YHi+EJSq+gUBmx4jbpUQBqoIM
W5LrfqY7cZkXjS7jO/pWZhqf8KT2X/m2YLdpn35ZXx1kTwjlx9NkP2s+sOJ+MRbXI2HY22MoX0Iq
0ZtF8FcQ3pAinQYcxlJ6BJK5Eh19hK2e0HbkV2YVstwcwz7IoFOY8hG3t0Jpmi7mhPKMYrC6eo9a
lv+HtlspZo+c/O/WRSf8XPlX9XD70ie9zILqSg+44kJXaxBogzU7oixZ3uijLx846Uceyw2O6YCo
VJWX3IvR1MHnV7/58QW8Y4VZgDURa2W+kmPPfyWN7uQvF5ym/wwI0J2YZor7bTCmDeiudd0rb17u
tiBuLL7T+amLbgG4yJo9XQjQtHf3XvTSBloX4EtnUPhhQqDQV2kKkb75UjdtEcPjvCOd5tGBiqTp
8AbLgoxT+2eZCotgHxKDxH2gQtR2kM/gWUc47QHKVG9WGkP8KUgQ/SFlKpdGR4COVE5GNoKjbV4b
7sKVqNSC3E9UdagOZrx5fzH1ZoVL8wuYnpYCF/efs0l5XhmeMgma0UE2B7yLN6woUetvecnt0i9C
tVVKmjTr/Rrt10aqtdWR/0GCtAjOjdSyjDy7+76d3XFs6N17jRjRxbydnQzTO5eG25XowIPUn9D+
6v6areZcrl6odtfo8Uc57mFlFsKwhKtpYgR/s6DY53POwapiXWU9LCz4HN85b0ocNwe0gfmSIVJw
/t/M3m6VGLUMVC14YwNzRW0ZVCIfkuAUdP8YdckCHi3MhTqGXeHPt/ETr7tn9tdnWCOAZ7dok9bG
L23/gHch5tRwyHUBdVKCEWMCyhEZ4G+N2CyokSzmmBg9mWj81epkDt7icSUJjDNzd8pEOcqwZBGT
QUR5YIUgH4pxxImixd55Rn0nySwa+GNvMJpS6gWJD+TN5+NlaiCq3mdMCehfzo2KE41br2iN4rMw
p09YI/g+6PDe/qb0cLda64nXtr4x4/si/B4YywEjCCB327dDajZst2g08vu/hglbMl6YexY/9+4B
zYTDMUF3OREgSdlYF6OgvSbCUNWUiTP9CVtMM4UgZ0t5vuTnh1z/TSWy3mMPt1EE7zZmAvF1NYmm
RCg83tB5fcedHWY1eB8c0Y+4xQzUQekEicbu78PcJwHocB5h626QlYZTFZnDQvxxnbPWdkFMSxlu
/PqTvIM6OWfkfWbCOymDRVFpw+qRCtxdu0OiB1TVjyOaFfNTpQleDVrQFvs9+Qv1DVpbIRLk0S51
KpUv6qjyrsj5Ua+i/QtKtrNnV8DiJgS9/j/aF286g7WVuCNbMliAv8+H5L3W2quihbeK3r1qyTyH
dXEgRGkv9aL74c5qNqRSAJnJ4QH9obYPK1tkk/he5rldmoqxiTgMZ83lCSyrIL8sap5E6pBoaw5a
fACLa1Z0MucK8cYSpFQ/pXtRaIGqC4Zxq7xzULuKJBkMDpsvAUsIKnDA+i3VGC7XJU2nDxAdQX4z
9YR3VkfRqLkZWXb0FLGqGEy4I/njwyl9FthTscAb/Y9wCwxY+AzBwO4wdEvWiB5A67UXJRHrJoBK
Co3/kSaa0KoHTTvhAZK3o4XxC5Oq1idrANSC/2RpqvOIZCKaGjF3om8gvvjbmu59vVtBAje+Rkm9
9Wz5BbF+vm7UTPT23GF/HdF11c1zaGAAH1qyFUoaoMiKQwXx1wrfb/MOOmONPomxTMZqXAvrJ11Q
A89+aWCMtzgtpNP5nr7XqkzsIbABH48hbotGpeDejkbS7l0zgSAwhBILgAdfW+UQ1lhWJpk5JL6o
fGhsBCQnwvjHgweRDRrD6ZgVOpz6fXYMZUBYvpK0Q5ZdkQ1+p7bBeZync2E0kxNWOq8/UQIWb5ui
gXjfZtiYFXqiglvV6FAlyGmiUozm28SnOY7PtR0X/GwzGP5/8HvLaDKSOWH2NHm/j1YxNy+p6EPm
soCtKbz3yO2PY4naVEj24age8xyto7SFf9j6D7HDRtKabzWLUiYOCs9auSxkvgj6YJFoQrsgifkZ
zIFWOz+D2iqCk898nnupqyrOOEXrVjQi6k7QDHvSTExj8V3k+Zeu+oThFq1vlXaDK7auqbtutrjP
OodW7tNx0OPnKebsV0RUyF6kG2fBVUzutSu+VlMfH69n2Umt/TsmlY6NDlV16yTg/e5LkqxJ823T
uGvLpvEbvOjPBRsf1fS22jwBZbmHnAI7dBUA587RkGbNdhhYjYMs51ZvXlcVDqllBnSFanOA27oC
HoT/1skwDoAHMAcQQryqQ7hFYDg+ae61uauPExqTeWy68RdsOM4XpHizh+MXxySXa+nK8NrVcI4Q
+hUcNmQHWseWgtEU5m9nzuxkKjjh2Sf5RtYjKW1iAj9COXaCMS5U0xPJTff2/KZ9vcCExDe2Ib18
MQ3wDL6IxjzESGDIypSQzvW4DjkmzK3cWF0tbbf8LrTlwoNYnYDUqosbd0Q+9s/R+WSnfftJL6K/
qlNUA4ThH/bakKiqOXkW8k0oIgGkImx9FGXd21dU/CdJsX5iEu4ocOOWW93fEIBjB3O3+njWdVwe
EcgvYkH8TrCHOnpYWA+J3i9W3koDUPDdhHMzQAkEf+3ekYu8sxu3x65fh+0S9VBrBZgVdfWu2I2r
1CEY5zoD0dqXbmaBGfQZHi1KuXpAW8+7ti/OpNwglHwHXXe7ceULzVoTv+uxtaVJh+xkY4ZXtFvW
h96WKuinftWar++izUeyMfC+T1NAgoWyA3qNiK5FWOaqeN5UkdX9yAYZjnIfhxTZzG6uJPYoinHv
r6wpe35Fiu3moitLFHR5EpItyF3X1fGHQoRphgPTwCUSywKnC4zJB7cW/xzKWY7fYU5vaNAGtE2l
KOSME2vWkD6AJU83Cyoni3ymiQI43TeIa9zcGd2HNkOpBrKVrkP/ZfK55Z1thR3U0UnBePzafow+
gGkqOoZlkoLpm8HFbcHqa6ridy0Jc90o+SvazSyZHwOGTY1sKSYD/z5F7cw1qNS3Za0sK58v5dRo
oCJ+LOhfxLtQDbkZLlT9J/Y9BDvALuDvW2B0N0s4lZNrIaWEz4sOyDdVYL0b8rkd700sEG36wrqD
4A2W3GbkMYydhO0pooreqRyZZcWq3rR3OGXf5p7KpHwnpq3itNw9qX4kDpWJ5RovdJay4mndicPJ
QkZNhwUihBANHZ6A0Zee4W9dr3IfFpBclv+BrIqctB51I7dsoQiBmldzWImMG31EykTBrc1+DkN3
XnzQXvuSBi0KdrAXDWI69JLCBiLs3gjdRcLKf+XYPbmK+PaidNK/SxuMZc8GMB3GHMaV04GXhNBX
qciUAKA3YokVWBzo1Aj1PtbS1CjCMDHTrk16bJRT6eS7wxbCB34bAGj5pQ9whwLfwNXOBelaa7VI
Gcj823uSv58SvuCEIxwD9B84SQeq8U2bY4Zxwvtzyc39UjKGIv0Kp1LVaNibh0/Wv2bdqUphkbo0
sUHjGUSuG6DOP8QlZ1eNwOAkC/1ZiL+1NMn2Zhi1j4a/iHGtcxWAuEVjDLMhINp6TluXUyMnKiJy
67h2MJInhsErg44lOWyVgKy4LTX2+ctEb3PvE64shPcefYclTiQtm2QSYcY97IMQUBveqHYsiWtn
lUtqg8D3yxscRe1zSqrA7rrow4uxVUbZnweXil1Q805v2cL0IzD4bbYfSqv6mdJPEqe9t+I9G/oo
1eb/hhEtJJJbN4rr8A0DeHvDs26AU8kjDfyFwbfBXN+SQcjaVc2LtbpnZMFJtBpy5jy6SWjOndNh
6T2TmdJO106snheDWR5ABxxKn6JbxHya+f4fk5wA7MNdU6+P0Nk54HsvOl8QNRjS85VNy+F+Jk6r
lq4dm+EYg+QaUmfF0lWFqI99plklZQJ8pQn5COCD9926FUXysWgKp8V91gnm9+ExFM5oHVA74TXR
9NEEwSJNNIDD61hLzXQ9ma410WYEg56k3PdOZwF+oPQMhnkKQImzmoMNAJxd7cj2dnE++ru/WGoK
uvhhZgynAmeNFAHGNijkMyB9hkuthejoX9qnKwDsqlaVKXxrL9NdLVMFthx5G1aJiQ0fehXHTJWy
FsLZoMFfcFaQG+hQkv8c0lCzC8ojdu3RpOX85SktPJkiz07msdKCNcjTXu6UFEnKN91Q7OvwP70h
EuCD3qfFQJxjepQ5Tl7dOnhuLnR9yphGWlw4eCe4K3Q8IqFat3mclyHJpkEF5AkZ5F3LFoQHwIf2
qhifWaGIzzWyaBFYcJjdv6PsRvkmAmjVtNiajsfDfVNzrHpJGnvNdxbye4NDoc+VcPLjgnCCfYQf
uLWzRwkrChlOOyAKQJWSTyrqf432t6GlWsdnnf8O+56Lyux6IfMDMfzQbNP0J2JBy3p1XucgTvDV
C/tgO1VNN/1Xv7C1yhnPmesV1D6itUfb6MU83tkfX5eQU8HfpSdnNkU6hVSeO3om9AWa2hC1p7QC
F6yH+6FfYyaXMBatQqAwrCafptVbHY43y868aRFRitaiyK9Vruqi1SERsV2SQDY+2Y8eFLecOhLQ
4+m0E6B9kTIRZS7LETTlVpk5yE515pt10QhbOiczDrfJo0067O6Dc4i6YCI2eWRIncrWEe1nIEt5
HZUo0dknZoReMfLfiazJbAcsIk0nyu9A9hG33Ho5tPNQ2H1IMtBdKd9B/Ltm1OzkU6wrrgubzLU0
WJT56WwVo643WXO48Zz0qlM+jOz4bgu+oXa3jkYiGqH5tp3ZVwtV0/9FGEdeNBTKTzoec6H1RbQJ
DjZReY3RWeDoELBHgm44vGRU7oMBCVPT6CQNyzO6zorMNJdr3AW02OzwLAnSGKP17AamNOZrISI6
udc+ojzmklx+w/fpRcEO4+F5b+Cl4jycT2+ruR4FBEqP9LuogXT1f1vMp6Vhrz3V/nDzGZyIGAQp
N9/i3S7Z/66A1x3Ig2gy6jLcaeMDQrGGop3fOXv4LFxdoDTv8nkWj7TwCsvMmIf2UqwJPBhpF2I1
ck/3/ikimOL31wxYwZxBlyBOHQU9kB42iZhz8n+mUwaLmxtkS4pFF1PbEGjULV+SRfGrJsmI2BfW
zRpYqvYIwzFvO2NkJ53mmzFhQizQNb6qAbEYEDXrLetGi4fgbmePDmm3othGJdDDFsKxVah3/cBk
WxOJxB9hhUZJlCzzuwEf/LrXI1l1K+iKA2wS97wygnJhY1ybu3z+RtFhTYE7aHW1XbW5TPZbuRJ0
FYwTgLqUNdtEoMfAvNm1WkjbKUXa/y/r/JedjCQcSXDvufZ5qLEo1Lwrx5ThUuGVzXShDTrxQhlc
m7WAFc9dTL1Upxc3zxwQjVNC/GP7HSx78L77Ji/8idKiSzQgR11Eo0UF+/iQdE33yhTXvgdp/YzS
QpHApD2owEPZhqoD7ptXUUaKhXxGzhQluGyZRIgtU5p0I0gL5/00kB1/KL0ETmkk+XvVyjBgr9g3
Uk79xJuKOsumRqfkxceQQebFf0LkqYY9sOwnBEh9ehDNvKe5kutcvsWnzcHy1rTJ0oH2X+h6MP2j
0UuiIm3ZHrJoU63Lcgqh8pP7q8+BSGzhSZofvJJ7KWz7uejgEB4pe4ybJXaNSYVlqyDoz+QY4PLr
Vg/7RnyEC/qVV7+4xfma+Ok1iZZcxM4rEPTdqUopGBKH5fw6G06zrcShD0kvcqTZ+HWlNpRLCQb2
VbKt73cmiiej0orzvvtw+2F3ywErkI9hwpVT5Z4szQILtXGGEXWxUsgztmGEYe1DbE93oMbv13nO
buJIBQs2usfj7A0T0kbFWHKUzfkIUaYJW+D1Gray3ChojPMaKOZeKpB+Q+8kYprVXjE2Kf2E7KGx
8aELdPWueGFAmqJiNQ3+GC0mrnfxVPx7uzULqB6T6p5lVIX36GnhAQjUZdv43g6eshz4SiMtW9/H
YbgOaGeGVCfQeQpVRQg/IXScDBv6mugtwN8FBjrzHGkSHjyOhjASJ9p8jI4zBC0CcJmxfNcpkZQQ
vDDeifz9WLCVvugWDWHnUUiPW7qcsB9CoP6qPgapvDyMZtcrqyX2WkTuW/wtkuBryteIR4M85FXt
3zYVqCxs9lyaqnufqdzMq7YxHDcMDYtvb3I5S2sJs5V1QnHKaC2zuJtuJvnWOVIr9bMfUyAboHvT
0IaOLV5r6cLdiF+MYW1D+CRgBgmwl83N+seEm4/KDFYicKR2kbh4kzi3BcUKLsGZPzWQec990sf+
A7Y9NhgxK6xYP1lE3osBg/eXsWIY3h1Y36jiy2fm21yM1PL6thtq04FEu6XwtsBpKvVLrNby6ym2
NZgDuEC38SV24FjvVYgddQ4PMYNtjYoMPI8r5Zd1k6VdsIQJnLwLYteHQXOhmKZGgZQjO4qv0loQ
gdAOAKB2FZr54ZLDNeaQKqnpWjalANk3TtEVh250lkd6RpzKv8u+W21OP6vNfmEOfphu/PMrMzea
R0zqNFcH1iKweGA0MJw0wADs5uEYW/2gQfdX7dw6WDunBoWEMgRfeJpx1DZqKU+luFmLGvpFzF5e
48rpn8eeB2RIlC373kr4f0X60l3Rl8cJsBjFUHAH+0QDCz3N0BlpuGJbbfKld/GnjgXybKxJ4G47
S7IYGVOHhyeUnV3vGxAiYFv5k4cAtTcaMTLgNzK/4/y9xgG7AZ+ojOU/Wn7go7/VLSb9lw7rRdET
8nLF+TuC+JXw96ZxjRDGiiFQsZEmQmOCfAg/dFCfxZ1PkaKJM8zwIY95Ki3tA1Cd4YK5ZFvYcLka
5s75t8iJMZRr9ISOJbqhLWUmpXCpD+5ZdFSAsWKBHhhY8c7gjBGXr6FNL+w7Usq93rQbYRRmgVlY
Vw9MRsbOv3qyk5tl/RZHQXUmAAzTY61t6bfzLgT/noCXoWchXbjfBNN4GAPpdag4BeC6bEtRF9jS
RkBOXGEg2+IxS6NdFP0y111VcDRTi02CgS7vMz+o8eRQIY38T3Ow+H41dDhY/F2d5JIHv0cc+sUf
2eC204g+4LfCwNpgUBI9d+5zHlqbCy9CNMT5DKPw15qJl3H1Vp+NDfs5VrlYDhU2v0nMpgngeEPj
0wRfv2xoPLbINOmECiZrgssT9AMelq7OIFmwfCQDu0iFXCDqMu4MbqJxBDudC0A/+i2cj3U548Gk
kHb3Za5yFgnBjmIFUQUghAluN738fAY6szzrsmtqr8cE852cu1q3zsRN0qo5lB4Qf1OvpSPJkC8M
igX3GPZGTwydKlgqbJDkjxoU4QgO/bkAjfU/Et2zEibytrRtOeunpqlHPh1VHipK4yPI2G8JhRYa
64JaZpJIkdIi+hPpykmLNB5xSHHQZOrsaMwWbJe2FXh3bew3lGhqaEvSvb8Bjf3q/t1mMxWDj87V
QuhQJzFjeOatIvBokiRhoXsXrmT2HPK1M++NLd0WUBeGISfdfWwvw2mcSx8LqCYBC/ehRPYKwfN9
x4lputtGlMSCMrBpzTyGNXgQ6Rs1PPbh8dWlzGZc/jYtD2zVzc50f5ZmYA/t296ULURTwvWgN4gj
o8ZjVi8NtrC++QZtYoWrMOv/uVYSHzTB/2Ab9et0DH49aNxoV57bAlG3Bwnj5+kJIH7ni5HE2KjX
V5oadR0UT/dwyzasMd/qyad/pWnkfvIG1nIMyg7Dws8aO2ce0SB6ovw4jKQlxhYFJjiOWBbENq6d
BRTAkL2jmfcAT73Ycbajt5o9l2WQpFKy2AWAoVjwgDNbZc6Dgkw4c/eCqbiF5ZGrnAhlBzt+Ztdb
5Y/QJZEONgKs4Al3K+REOBIKTS9H6bOoztuAu2Fa+X/TFA0Q1XwzC4dkO5LJQABoH7cwfxeIgfmf
p0Hdb6ozMyhZP4qWUklZjTyPdjiHU+bdBi2osYGLh11cbAKVLv3Z30M+v5qRkGCmX387IOJRn2Dy
vit+c3LldA2eDTwiWrEaJ2/9SezOJ6lX+SY0Id88Lomg4OS8fA6Z/deflQc6yHm9z7G3nwfu5npX
ebD/W3p+RqYZ/VhtH/FZR/3Gfh8O3ueMNgmDlt9/QA7HOPOrqoxViqgZbwn1e4RwcM0jvCiXgC1e
rGB5c6nzZoql+nnBi9CaQlyIxIrr3SW6ZhST0oMB5FC8PMvMnKv7gT6fBfJS5r6+x+wG38BnWiPc
PD0zqA5Oi7q5xykPNNkMMHr+RhSrbLGEN+shORIYDqWEpswGssGCFYT+MIEdH/V0WG6s8duSx8uO
pUG2EFV8otHiDNT7N7V/V1EACIJpRKvNrLeu/zcCmgLEUJiLw92Ls3Xf23L2INSyMKkv4WB3en0Y
FDzWPws4zmeQC0RJzDhLavTdZicDHc+dFm6zLHDuhT/2WOAuLcDFV+dZx8DxLKwNG+NVcDyY6/Sr
W8dVCe+2Sy9/uGhXAhQvjinLENRNaoGMzGaAIcEfQJJfxUOZQ/zhXyu9uULpMptfhWZs91vYw6sD
y2CV8A9wlpU7crYWKv23LJ82l0vDT1oamKXIhSjrw25WWaajY4ffvXwzrx6UvbHkzqqEUSe9tc7z
/YArj4F5keMVK/M3vPes0YWth+4PG4bmgzUTceoBvgHygHfICG63jG5C3rxttYx0E8wkQi9t6fd7
vai6LugCM8pOvmRi5XUcU76PludHd3eLZlxdL2fgMwlkf1ywYXzAJTF4JY4r4M9aECivGINwLpg5
RtYVuAR6Ja9/ZiOpL9DiHe6oy2npK2uzWgrBN1RqTpDw2Nxuape+15E7PgDFvCgSbUtjKDGxR9Ru
kT0oRXuBJbUtNCl9YMoXEbX4vmtU9XqchVS3wYECE3j7+NaxMXSMD2Oa6NqIco4J72+CAE44KjY7
pnzvFQvwf5wTPmRqBwkF1z9IOIMmblYSilPEVphdAlC7dQGyRQa07l/kBtaH3fN5G49ioS/UgJTr
Sd8fC27xoy/NTD0aHrYb4pVF9vkBC6hlvZ8qo4uPRt2+GKjfjL5Z2ejJoiswM+J9BxFTSoljp1AR
9vf6ugONN3Qqsd3bvu0tZ1Ed7uWK/hAwSVzNm5kbDdIeTWBigRy6OOqcnpYJ+7d89n0twq6s5sMy
9d9+V1Gn2N4eA1rNCCpW0V3WTcCzsMz5wFfxT0SFwbRHBaDB5L6jbGamCq7o6XcE/ECW+v5rM+oI
j315OY62Kj0iMd6qPM4rEIbtPTXD+vUW61/6+Um65N/A3B2VYygoYivM8czIyiDokLJpmIFc2BQy
qw6XxDgfNfXIOLUyaGZEaQ1evngnDDlIp5qaRxD/AporEukseogXACQqD3T3GkePus0hJEbdpbP1
Vbx/TNi1aPoHGdHvLXign1yFrZ6EXKQs9NvqQNcO5ZD0AMHpmJoKciY8iOpVQZnfixRv4BMkXfei
B5xc1iRYmO0nQkgu1AJMUl0GmOS016OFOfFMtrJmFFk+R1n91vkgBCEx2wQtU5PwlkTyglA2rqKt
3DnOIvrKHzHchLSkgtkwUkpVrZOMdCOG2QQ94L94we4LzKUZLuNUyHdbBcMIF7TsRYxSCqX6CPkz
9TH2yHI5x8WGUfWKUYZf8rCHCa5oRVtFlbHjGGQ7AahCJWMGd9tayC1UihKZFKnN8zWMsdr2PLok
69jWcWpaxNnXdaDveIR/z7BaB9kvKgU/ZaDtIOKG4cpGxw3b8pJaBr1ipZoRMhb5sQ7bhLEH/pn6
VHu/3IlNsw3t2J2aDdstUPmkHz9VZl69jc25OKwqffNvOeFEz+fzLQ1RuhMz0l2OhcUY9hR2bQ3Q
3YNOqd5tVRHYjnizMkWwpHOwCFaOt3LnPBU+jGt1hIOb6eCeAgtfFi9GbsCfvAEToCHZPjuJ5HBR
w3CgcDuNay3SKw6sKuL58OdBcFh2j4rht4WBBuQ0CuPp+lJEMlS+UXz3ZJh1u+Fe+AbUnrgtgMBd
r+6bzXwP2tVnSEjmCccEi8+oqgfGjTlgdu1hPOLPVzPwkUA5yfxRm1pDQwMZUN+3pWE4+Zt08Vwc
U6Nt0R0G+9xYeKE8Rerst5+PlzAUXdJoX9aeb21dV/Vqi6z4GH5F8VdTQ+VNJZ1YDtRVhjWdWNth
NiOHJs2rDvyGAXSz5hWO/rWcR42Qedgp3OGv6UqKYcya4zUx2QiVzI4A8CmdQEUImyXLwmcGv7b+
ECeJKFYEAq6jzdHyT0NgH1AtzUBc5dXAKrXptx6OIHhfDPP2k4P8ifQBV9cRzbrdMBBOLwV/Tjf0
FXQ/K/eoo+H9lR2nT/mAkFBAAJzE1JzDU5k7Ie10x+t4ShC2rxwvf+mjzbRjF6yA/XU7+oMdaa+7
khqrOXnbV8p76DbnVGQ3GMPjaFq9kzs3mP79TTTmu4TCkclo3YBRQdaEz7JwJzXiRI77840kavCp
CIW6tP3cPfigGkKwhQJwpNodf+KCzEu0TYOsmEnnIg9K6roJnCnu7uG5MUI5xrGTdZUjqfEADsdc
vdcMqkdc/oG5Cx5AoWc7Dnfk77krHZqtc/swQucrKqpqZf1As8/ZMpbWW3Ejyf29C3F3k2NJAlo9
1txKoSmRsFDv/NWfavFIQKhR7Fq7PLaBbX1d1kQeMP5VKckCzEARq7oBLLE1PucSQEQqQj/XtN4s
ZxQjPlcJO3sNw/3uWR3ktd5tPGgYZYN30V6Ek2qNRbbK0JSDQthu/4Qqbntu/OY7JUMkTDlpg2do
ewQCRIjwfSgPD5wQ5O+nLmUt5gIm88kB7oHnEs42beOqfFA0XgrKlLjYI7a+tJNjzSeEjTBaBUtq
97k68Xc0fXAsunrwVznbb9ys54LY29zECTPV591dvH8KVWHfek3s9NSrLvID0wpGibc27koyB6ap
FGgPbz2PSbOXZ9WQlG8pufr1msArMZ8ZH46f1BMhcy3dNdYZMbcB3EQtS3T8k2VfP1L/i2yWl/7D
+M0G6et/m48zSvuJZtVK9QYULGgBZkSUoFP2U4+l/4j4Zc+u6xb0Ksbqen1WedBz5jx07bQZr225
RTO26XFT085pjL1OzahXRTYzL7IWscbEkogvmub5vVL65SrAwiNtu9PY2yYQBVgbwBZUM7740MuY
sLB2csS3ML+n3WoioGxSvGJTgnT9Or0jEkZQ9KuaukHATQfX+hovPBEaTP6Qxl4NMCRPt3WANgRO
RJuSAIJrpoyHp+9AIwZhxk8nIsyQ2HwPIbkGz9e1VVr/3JZfZq01X+XaPmnnuGWbvz8sscL5w2uk
dzxJOoc1f0MeoJarvFnnn5EXHwPVR1S/DRXfP/2ld9qW/gvVvvAxiZI8cseQ7oDh1opeuEggvfk4
ia1Yh835A4KazUaDj4jYtB9t8tow22zkT+t071QxjamnvW7I79M1+MXoQbio6dcLWgeF2HG6Zla3
SJenugGa46q8SrvCuRNxtQaWKTfuoRqJpNgCNT/QGNtZj9kUAR46J1be5YDEaP0kmP8bIVoAgvkN
CltaCfCL7NuJoZqmudBj6IbZnqpB0PlIxQ89K1iKWb6yoH9dXxPNXrhC8QaL/PE7nS64Iirrk+d0
HG9Lh/twOpfNjNPhBiKk+8yU15PkL6sXfC+KIE315XKHpbVUfLItnze1s4KQGgQXg/fWkdShW7MS
n+gZ5m/7BrWgupqCXoz1vs3fCCFx4Y5/mttjfPtDbddeIwH0eCUQd+iuc2/x2SdVgvj9MI/OERlQ
AtxaBHqe5xshyS1W7Cd1l5yMd04bR6XYwKfREZBRtXX+9sZxfK/dwWivpxd/gVxr2VCaEd8RGIZ5
t7VRDUpDDGD0kHHwrAjmiwSqktfxNb+p0zRltaqabZhd5e3MsjlnZpsfHmnqzp6sRp9ppFhMqNyl
KMYdsyWm3nTxLlQ4n16I5MVs3vEO6NUETbGw5y/Co1pARRQpMOTFglb2SWwMR45glBlabEPLHHjD
2+TcbDI9e7SSa/JyqiWpgMIzoL9fcPyoVQd4Wlc9ydmUUh4mSb2OkiUetA2uk0Zx0JPdPAVnyj+K
fXyVAHT1z089XTltdeN9YsC1C93UdLhC8Ft1xpjl/YZR02Uze6OxpE+06tX5EazTylGy0bHENcoj
9pwis1Glsj2r2eiNocfuIRViGs+MfFtGmJCl9Uypq4ixqVOpUOG+Kl9v8PnV6KHgB0JQjRkcLRaW
6WHhY056LqXN/gtAyqwoTmGDJVCKgrdKVctJxupzbHoWp7n5AW+IlzCb5DzVBhs4uj2bhk/rtPU5
x69RGvsy+vCNoivUreiWTj0v+JlF8ZR4Ms/qUQljqFHT/MXxFf0DIwI7eYX0ncXaiXmI2KbxtU/g
OaHkdOp5PB0XwPLLuE5W0OC1dEBsvO9EciLkVrLOjNcyDt/150ps0UUPFXkEU7XCfsBHuS2ltJY5
eCoLm6DJbwX8HuTCI2O4Q4tXg6352NWQHhwuMcaxTS7klQwZ1G9gQccJhQ2MeaTb31GpzhLUycZ/
hqXlOF+5lxyxBCbw88uakb+rmkRP4SclzYSTiZ5OCzdD3KccDwNFPna5r3w13phbfo3qx7VmovBK
xss4STdiZo8TLD2i5OGHXPFNVP0kpZhgA42kBMsqmRX3/W8MgZm1nTmPgsEPy3UJObNhaGy1R7li
gU3lB9gXppbRymbP/FTfD8Nqb0mwx552Pek/eX9FrWEYmX99Ex26wO5ZkSjo1647zaGvlxIDhjT2
OTW7yR2T47d85c91rfzlNd9LXtBva1Z4tYmseLHCZPkqekoom9JrTbepH32WKh+nnU3v/0iuk+1w
Zig0HG8LwiYUkyUmHLs12cQGOyGGsRQH8r+7uw8SNp+hrkCXMazJx3YJCkxI+uSGAe/Md8qTKrs2
Q0Kirq+6eN7Txu5cIt9cxDDti6wsxyWj05gBT0dhEZUOXanhB9dgyVraAxORBznnVAV7kGfeM9Wj
EQIb7zMMx7IJj2L/Gn4C2LD52BmcQ3vM4pHUscGAKyVi2z+0PvQKuGuV6qtxYIIhbFSC0hpLbfxF
YXtPonRs4q+3FcxF3FTXd7c5WXT7Rq3AOqkgBJ4bEvEQDBgJLLHJGFEy/M/hdH51UGlErbXoUIUG
Z464IEDGxVhBHRYLnl892V01SrGBsEfPjxlHsZ3fWcnEszcJPu+a3l3nOWuatJeSEuadqOvaBfjv
mJvjlUHWiySDVR0LwOiuRr4T+KBnfYd0Vy2s5Kxg6GhXv2CWIuObCUKsSpBFmM5wPyw8Ke5Qq0y0
EYY5iSn2Y88R+ZQjvAgSdHJxGK68PYGJunEDFkrkSGMcse1Dlxp76LKER0+Z/rpQFaQwokkrNnRL
m+A7YQYlpeT+wOTfZQdvQhp5ewdAddaVJtyO7MiTlWDSZaRZ2PctZEfwqAajtj5XWij6VWxJ9srn
B+WawvBdGvYfMccCC/90ViMDtOiKOSmZ5J5d7LpRSzd10/tM/id7Ta2YEfHAJ4WXEN5LFJ/nm5+X
Y/NWwE/ZkFZkOs+mM9/a+VVSV3gSld2UM6KC7bxBTGoug3pHzSXmQ5lAaBpGxjWmIHR4EoRsV9nG
6L8k1DEjLMXdzOy0IOytoowSZVSigzfTcDDY+/C4LPTngBK4VZrTkgO28/0O6X7LOxx6MljcrR/a
oOcR8NdslLr77EHKapsYWkuLD1kM2MmtU4aGvZ84Nd2IRGduF7u7yf/pqPp05EYQA7HoXaLkJ+dm
8D6wn4PsRYzoEn83mUnBLiMB64sn9MGUsX362cXO4cNEqVCvzRS/qKTKy2m7oMdQTMHWZE10CRN6
XFVahe06QjE+NdjMsuC1ha/zm/k7b+ECVq/TjLIjXgFpxh0xUPC9gCFWQmzlHh3V5W/qBC1Px9jc
jRwQYTTFKsdYhFxZfuG+ZRU/E+mPgrPx8xEGBXc+SpS2nkSpzejOXpASV3TnnjGF64QVQ67aX6ZQ
B4IDEifhD7+f89ElM16UPX9aFlkrD1fo5E6w600Ae9nrWU8uGwUXOKy206G2B5hUKBZLBEznG6Ny
BRFYHYi1bKA34C2NyfTdgJ+V69pu4By/rMKATUqX6ldrovqYUJh/Ere8AcDKGYoc0R8z9rDMi9hs
PX00ixLmwFk8dQBZJelwHDPZDyCJ2q9UO9x9HeEhwzQotr6jLizDy9PrQwzEy/OA5Onq04SiCMbd
ID+5jhDPnKIcGb9i3dRbHIKx2yAk2OV4pCtie2VasunBUrm1E1fbn0m9tFwjKmETJe1RKcwl9FLJ
gA4ndELo/ukn4fMuM05JFT71xHFwNWzfuOpWCDKQes7VC2uLlfnhVlNbh6Lf2mRtL2jpfuP+ISps
YR2STB9vvv972m8TeW+pbf2vH0/VSZsPOydS7VfMfxlcWznNPaFYRgU8OKelzLc6Y0um+PSxf78K
UHpFNAVfI1WVrRXEfjPyBxMdb1t49a48B0bbCU9aEy5fitPTGhe0jo8AQAT7uHLyXlISSk2fKStR
mP/R7zX8AZpLpG5lklj7LK0qQI6wsIz5vB+LVyi+JACO7MqY9ro5Lj0LjHWVxRH/iojpWxZ7La86
xB69cQ3JuP7lzUXEPcbFw+Gomg53e8PJOzjEvBM/8ZZfGQaOmv9CsA5xfzV+3WSVLGBbQnvnyF5G
c4rNkAT8P6z/fi8D7GLMWHOj5ixZhwIFqoqUiDJe9nnW6KqNB2s3IWAyGSeg0RHDIbVtrBacIWkV
ztbWFY49v0828vS5uAnGqn3+4hUJAOsi5hXHcij9wJcq5XI1YQGpXqDmgiiK5hLOWPbTVh22AZNU
4CnUGTyPSMbmPkf80d0D8Op+SmfN/71zENnNCV7/+nK/udrQYeFUsj8IG/zr528kXwUDchZdgHTq
PJ9F9pcduUYlT6h2hWJepEJxwCDZJdx4nJHOCX1fdhUzcBXYgk/DUlMbjwln2Nz8yPft8IdsZYg4
6iopbQgDb25mxrmjxfZRjzHNF6SOFPh3YO+jiJ4IqJpg5wj1GiWfWx/nYleCA9Q+YOD+70VOgfoA
zgAfM4TZV3Zb6bsahrzeZAMfs91p7YTJey13+0Z2vOH2Cf+pAow7ot3lbrNSFaEJypleyf5zJbxC
wcgpo9PObCBvehndV8ikARaMF6IgTYghsBvzO15imESECDWaq/9GQJJ1bD0HB65YZzzzU/0URC4n
M8zezAgM9hqG+/nzYPiVrH5wiRbVebx+u215UJ4kJFgZUhau8TK0rnu9DJVyh2pjZ1jz+g2Ro7EF
+lu8W+giouJ7fixL0/8THJMJhNTw7aknCjCVkOTjVj5/NjJx9mM+QEfpdt9qBI+DWZxN7x6x93ZT
meP5xI3qnO19TnuTqNZi9RAcBze9prek/3Kl1KjycB7+RFDf10Vz2rsC0iWoEB9bKaK0GjkySzO4
roR0ckFyGeOd3Gns2fUMEskzjT5Qd6Gy3vNBXjn/AUQ0McIgL1L8i3nIVH8IpovEveCgjhEav4Nr
b5AbWDnlnqncBXA8vcpE8ME3f4cGm4YLkposTSpi9jYr4NYoIlm6MyCON9JrRJJsM6xXxgJBVZmn
57cLYWHrAqcBkG4qAc+O3RCcSLZyGHAeQF3/MesaqOvDBSb9mPqinPN4stn79RXoqBm75lv6WPrp
diNZOqaTggdqnj0w9hz0O1acL8JMVzCTf8jF7Y1zP7L4FOxCPqEtZqDwX9nrexmNO0OK0IL6oO3l
ZUUpKgBPhpUJiqaaUoiqc5j13FQ7NxUbjpK5HCykA7XfDlH9LYoriuYlFI12sOkJRSxEq3X30Wn5
s/qUonkrU/xdLWThX3BtHaDtL4ALNHRJMAMr5QpyaE1eD7StG96EyosDoA524A/KCCORvNeT4tBj
ioPTM1X1T9uA7CGPXFbZ5xDxfVT89ORr5dEDAQmJ2/0SylMHqZn5W/ybc0yn+3vHc5/lTlf13MmO
T2M4cBMkYTOjAuc5t0k09UapXVB5TRjsT2yUj9cr2S2N6vBbNck9amvF1oi2UF8oljoAJII7cIq2
FgJ9h2c4D2wgySnWS/NPdB45PC0meUm+N/P//BD9jQmRj5R9z1e4FLFsE7dJ30ouc15ku0V5PIoR
ArMa10WHrmHBeEESyMcgLYgG2tegy5zJ48nMLDDGPWlm8FbAWUrB/iTmbOQ0CuTSuZAyS+m5sRjW
4tUnbr/yQbJwwroQiuTLCxXxDTStWafMgFhOkRuQYJXs7VFTNFzGveyi5wol/S7CMu9h1TeVde7Y
KEsiuyBBfxYuXpb37xvJyzwkxg3vt7ata6sniGLBsnGcIxDyahH9EMF4AAuizbjqlvYpI8VIbV3i
uzifPW9g6pV41CPGy1yH4r21G8bGdk2khtAu54GyfNHL7LSrVpCgzq4bCmziJT8yRGU4irRb8ggM
fWV1rNB8Nwh3CYur5/KcnkKeFrPAoxsqcte/FnuN+6OkoLBGGFbWZ7u5TOOQbT4irWI/GEOcN+yv
0S8ixlm/nMiQgCevTduNVcjNFApIUbTrqmmehcXNce1n5jaz4G7SI2fMAturZ1/jvRHmjiKwy0tU
1HhR5yTl9YuBDQUnURhsblDvy+aIEC0IqPGcBKF/lbkSGLMLqOz96pOivRc53Yowm/rJDxM4SrID
ExWA0ATYnGVwvz2tvawEQj/2lS+bQmjacBLj+vk1S2BF0sXjV/TX8qos/oNWuoGRTAHntQ0ViuSF
IdeWpp6vI5s1AsMwyWwH1Gtk72WCMYbRLtTPBR3cEobIUiANY0NbMC64whwPKx+WSxC1YDnZLP6H
aaI/N75S6+lYN2aDrKsvWfselg5M0lRSE1FLuLKUtnxD3NG62ZOboepd4hlf6+x5WfVNzQWRdzNq
F2QkCMnh47IFUuOUWeMf0Fw//yxlkQDPNIM5+7yaFdcqj+oW1CcugLdjWH7XraaqA9NEzdy9E3Mi
D7vLvjpmUTgxIiCONyQxpw+dCA5UcwdP/4+FLfK9TklJ+nDvQI6S/g+VIBIROEi46AEACDm610tX
wpUPuyIaP+e+0f/1I9Ojp/o48mYzCMApHniDj1Fy4DvQMVnjH062/ByTcNEtjUBrN53qm6qiF8Cg
rZgXi8UcktydnTWhW85mhJbVdKtY3yO/tEkPHXCF0qB9iUrFJTDqxsJ5GIh7hARu9ndHfr474jZl
D0Z25UPWLX0G/ySUZoGJD9OatjgzmwJRg/ITpfHov2Oka2hBdaH2hRr8MnWrDa8bpaJpMFdjXiOG
lWvaciMwfLs6p60tV32XY9beVlWQpC67U9Tmt06KrqkVj3B3NV2bi3J2IQt15for/rvdU7DbeT1C
JUy/qYmSO8TmBJcl6f/Hu8CgMslyPQgvlpdN5rmf/GL/7sHAFyRlGgp1S/CotwGMSedQiV0phj2H
pPwPfSn2oFmPjNsVhYGmY4/X6pjVQRir+rOLuFiZeb1lpVekLGhOclt3b3V5E7gbyr2bYlzJeELx
7jR3eZ5nq0t42q7oA3nOVXOL09m2wxDSeDToe350R3ohQGKMVbvO1vfERK8JeW7TOMulcfKKwxTI
6JOcrxgx+LNwcdJfmV6shAawkAlHYa/x162ofVqXiN4fDiFSvBcrOVz7NgdBYO780o5l+1JjMTrk
Y2SuVBg/oSjByQn13cAtZp9tYNd0WuKQCXDekjcsau4ZfuP8Jky/Nrvg0/g/c08OSKN1AE0J225O
qcAgec2LtCARrIPWYUWfKcC76AR27G4Rhhx77OnxWrIbR+7D9lSMuhppyjpmoEJ4oXUwQKnprl2G
P56OqYlQMWn15CZL47+XfTURigavXs0R94Me+XBfUZBh6zJwmZMK4KuFDbI0ynp74Y+DMQub1CFO
wugDCW3jPpr1qqPm3blnpmtFJoZgRNYPA2UUMpQoGbY7lwJYWAKbJWkagWe5qKHn+1hbFaHWUjb9
Qlj77e3CvOdQFYNw+P+hMQA9APveunxtM0qkfnXNv6wyBn3sCatACW9R9MvUERcLMfhkSF5SLrUe
5F85v9RQqjgh1hoMwXV6t6bc/6fB8TpC8qBLGLaDgRkWS5paM3qGvnfwYneMTUvlUinYeqXnSZRJ
XRly7GlRfWC9bMcmGoB3x1a7yAHY1L965wUSdsMSfwY6GHsJgITdEJwZJv+MzGuEkMsK+tO1GZGT
Uw/v/8ftGq2d+EfiBWIz90bmFIUUcvzkbye3pL1KIEn5/ofno/yNB2KwKcK5kR7KPgK9Jpe8tmwu
AsWZ433IrmOTmouiUWvWUXNNT0eEm0oRqYoDoZ6SZgZG9iXIRqR0IZO6dkkp7lqttPZ9VH0TISTR
JV97y1X1x0mFpVhG/B4sdviK9lctPSGRBeefrpD9smoR4wXPIqNnSQwuN3TLDNhPsWlCDrQdEgYb
jXfYzSslMZADt82ffwTiEQDGzLC6FJWcTssmt+jX9dJcw+yv56Tw9Nq4pKTSj7r/KTvj2yulH/L4
0WalM/p+odoHFU4XUsEpT+zEYGwiVuJ/BKLDFeHeoU8fvQgbeVyvcNy6m1EXmApEqvrCGa8T+kdk
vnhMlEcu+24bWh2d5h4u6pu7aPdL2qMJODmdNQal+pAErZe17xe7RfYCYai+xbIk4f4bp3WgyoeO
Ij2VupABL6y7GlVleaQ0Bcglugqo1sUt7zQDcme7V2O1pxYeD1VdaaZFXmKg/mJJUuHP91MByAOH
1gDh2CbEtmQIvmrx7QOiJtLdN2EsG1kPB3+8bD5RXrAhg+Bja5t1U+S+xviPpooJPxiBmGW9fRwT
eR5N3PK1yOxHeeIvWVRpZshiIzlQ7EIUIWVPGXjTK3VwVqmdUHLVVKH15+b7cTOO3qtRMhEVwgkt
TvBQ3vCM0p5hzwy/nMcs2aLDewAkt9FnDTX2Sp/f0FQJ5tv0Z0k3GsNY8CTq7IJsHCbrm0IWDcit
FNLdV2EkrFiPa1jjpPBxLvhBT8W6daj3SIhDSqH2z6cmhj8cQvlZsRsr6Qng/PECl+KspvhI292M
Tys4mV7iEl8ddMGm0Gr0cbcMpGjqHuzS9mse3jeVcy+ImD2f5Qibbjmo9I6XWAAXXOOMJwD1T91x
wrRSwX8uTTlub46Bu2yVI6J32qU1E0IhmMvldpnjmuHYQNRfFBvSAXkCpiujmb7GkrgWXavPAJ8p
1rkMCAy4RiIBtL0cO+wXu4ROd+ugfFkrZv7ciOk9aD/woq8jNdw1AT7zyFVOfcvElnCDnehZQZia
q6diXBTl/cDPoQ8/fpwA4IUysFzLnbRhv51rq8ntpyBLoK2JCcTvrqmkIzr7trZ9KD0S6QaihGav
AyVa731zroVTEjqVweuO8Vt6DFYNHLO1kTAEg67b2+bJ9Ub6cgU1vN+x7KUaXukbrO5F4E8oyZz6
E8hzv1B+wZPqsED6UwoifVKv/3/Qmszf0bVCh+fl4945mvytqF+MsvG0w3I3DQAhD0cz847BU0y9
PeE7cMclsyUcbvcdbinMdbAX4lJRa/cULfF5w9Ty2oABY2RWl1n3XV9Jdmlj+4/JrY4eq6Ad1Y6w
IUEmveTWMpj2p48m/lckMFpbgbGE4RW18F619VFuJdYw2no4EZEvceSy4FbugcoP9dglmkVmYwhL
VAuCU9DHLzbMmW4IIi9Ew0tMaKtHVniKcVwSssF6vd5zxz+rgM9LCsqLclxd5VdTFCHpLpYcbB5Q
eT4BPEhYa/tZaQLl/qe91lVuMOwa2y9dseZQRCrGFJC6ulpFU+aC2g0UjdLgWBF5m6DoZLV16DKF
8CZ5yQQg1ttDcjNRQnZhxUVBdZBq2lXF2yoB1Rp0lfQKh5ro8LSMqZAHOyMDeV7lSbzcMe8nMFpK
l2BNwJMIGlIJdMqPqn+55JONbLRFw1eh+BTQ8Rq9vM0GY0Ku8eYeWx4WWO0RLt4pwZSHJSUQK6PO
1NIiHRPod3HjuKKOnfK0lKP1QYTEhhgL1Qr5inENfZVCiapZtGnA1aKuSJOLlt/uq2PJmliytp64
1leWz1FkS3H5PfB2iwPS+Qivdc0Vh0tjqKabgrb9xbW/xlrGx2YGOSPmKXAmPPmSv6SyGYdEfkOn
CCwn3ZYoiXZ/jXvIr58qOy3mAps9AlAidvu+Hjf3JWK31xwsp3RACbayhNjFSXbRSqUJ0xwycinX
tRDjNSPgwwIrTN1H+Ds1G3gdd3ynTI75HvWR6A+cpeKA4Fr6AC7khJs29XJY0+Mb3R+s6cEG7SsU
/rW0cZdSR6e1mWwizEgZnS4hRSBDCNqtLaTFJAaDowGaxv2IUiMR78F7CFVG9co8oupDe5CH+Ycx
pGvwNJEf+LRAlxNXYspps1ObfblL9CxSpeMZLKEPbI25BfSNzVehS+Al4Q/WCzogMqmtD/IDRHAt
UaT6ROC/dDWbxensecDetlV4LImHA1QLu/x8nF+mr3eCagMrrM4UZMteqL4KXqr70POusvOuZCtn
bCztbwODl/q+DYQIkxCeNOVQyeQ4cOpyPmvAkDS6vx3ap7kBbUBKvOh+xeP0tIpnwR/ysENnUNsd
pyHPooNfMe6V9eHR66Fi2Q/zuh5ooELTFN289GhvhrMiVSBUVDnvaO4/XAQPqJQ7CF7/PJh0czFs
8AD6Eq6+TVVPDlA4bRajVf1ZpgOyuJfZc5W2NcMRU08rEES5vm8+A9vLNa5c9lR06Eo2j2M3H8+t
GX7TfttINpyAodbs5/TONwlXK2ChOvsTTLsaZ6U2rMmctQA9TADh3R3NzsXUc/duuAlHJ7hQ2DsM
THmLdfTDKplD/ZIfwPV6PglfeORfGgXyubhHrQGsLYP4PugmtSHcvpnodz2aYBiS92y3IRrgQ9o2
JCMOtn7fUJbzXArbolZELClF2bcwpEzNvG383Re7JRaSn+sx/4cG8sXuCm5YL9evRj3SNP0wuRMf
YbQDi+L7BNtnvV8Ct/Cgo/urUdHudsjPCnfXVhNST0qkzO4KPoQR4sMEmGQqX7H8MPVuzCxynH7O
NGBvDFmiRiYFj0PfAYkdoPlKKQdnI99Ylkteg63zk7lrvZiJxLb12URgePy+gObJhVUyhgI98Udr
COtzC5p4ABLdeza2JzP7gEGYxmX/y1RO2LUT1j+YW8SZO9pQkokXtNebhXhfe2w+DkHNkAUxbooD
NkKF2kfeWobCX+wYLejUleyaeaMagCIf0RzfgPiaHQ1Kn39XG2Ys5sotHWCs37vp9/fWiMb79/Eb
51QYwr+sdP4q0n1QxkYa9bQm7YiHXe4B6QB5l3ZhrxUdof+3tTDDHbJTZ3a4/kMS9xa+wzGSWQEB
FjP8hYo1Go9mUqeCrZ1Fo7N/dahAmL8nlkLnwA1FMyqwhNQNnG8K/whF+QTDvT+Ik/rKCjSvG9TN
NfRkY90gIblSds0/593v3GxJahEq4N3g5cRZCiYao3F7Qrg6Ahw3CeRuAR1g8tuSyrBFy7yOZ5VY
lCHui5e8jZvGqW6tlLDLNLWQgMkEXrMKe8Wzazrh2KVMRiAR92OHLiOgN3AApaa3FdEmYHLTfDYX
v5dLGReJ75AzCWfipX4ks8wtN6bFBvq9w4LBxSVeUNoPCGl3OuDtnBlaYkIpVo9/jtZlytjiWoPp
h28rR/jVqN3cDRD1ImadYlKbtxR2k1/1ICUmEAvyNSMJMDjGMjBDWqmHY+XboTdaf8/Ao/vETmGB
1SpDMPSe3OtQWTzm0gaY7seWZuvCBCNf3uky4ORlqsk8b6HUzyxMfqu2ofFC9zhtkLBoRN9nnJL1
LvNXGiwvKsvD50x78YkxdyGguGY3dGFWOcmj9e563vqQzou3RtsXg3qdLZ8MkZAMnkgFvY+m6pSJ
BtfjTu1K3BgnAdVY3lt2I/hPE8I3gLFv6N72XOtn4k7Z2VulCW1Yq7SatI+XAI/YmkESq6a4Bqls
eygMJcm/wBEFQoFAklv7VeCfL0OfMS51ACKQAiAYI7k1mnvKkb+IfEitE/wecNAUk8PSQpKQbvAd
4vizGbnaJx9eqctGCmborrKHWs/ZpMvHyaiveT1DokXGYpQZ/h4UKnpq4f9KPQluItt7PWsP/wd+
2BVO3HtYCZz5hTQC+2GwiXoSdMoaHh386+z81NS1btxEeD1qp26gnfiu08IFtC91Q6laJABNU2PP
7dx1NvNhcDlFksOdDa7ma388YZWBrtH/RDnaeB4Px4G8X3dN4+jAcaLX5guH24bCesrcFVmKGMB0
Kii8fX9WCrq998+WKKdh9EnfEFxtZRiPjqjcgV1qTnHlXEZXhM+uPBwks6ECx/2gumHn2bXr/wWo
N+CxHpxp2MZ9ZMl5DcUkHpA+BmMoDI9tqppmHlwAUNRk7cAZ6XPTF12qqrFLsj8FP9OJ9dnhATx0
3KJgu8OIt6zuo87vAn+jgao4yKVdIgoLNchoHo3xnOj0+09LzIqEl3BhmewmaV5kpVG6mJhKuPxn
7SlarOWkx/GdxlX7gZ0pTt2BuRvCzZ/4GZZb+dqgrKChtcfe41hKrbdNJmmFihG1+hwHkcrMH2p3
8OmrhxmTCmtGpI40wiUy59h5+7XTLZ11glBCCPJVLxb1yT85VH5/eqlduNgNVzKBsOq8GBDKAw3L
trJ38oSsWOmroUARKpipW/WDuqeEDb188ePqdC7G2ZEoQcG1XlXlSXGf1rCUMOeyYvhiguYNFQPW
BezFq1ACE2PjsVJkOk0FrhAa8wBF2WyAiF3JMw6amsMIUkQ+ZruxPObp0UzsxCS/IVmHbpVye7cd
c2CQEx3Xjwk3SsyxPjeBwd008op8jj0v7JqsRX8lcnUXur0PomKLsedKaJH9BNXJGQrlnFZ0kG+5
4+SAzths0ZQJKJD1gkgdxi1KUmtwJ7iJawJ4Lv6YJD9C05rzUiSR+YEo4P1+SkJOwto8QOFdT0/G
y1KOy67AixDo3y2BhIcgAY8DemfLMkCW5jQPLT6hem4hjx/PbKySKz4RKegfc4ClGjRXMdnwIAzv
kZ9MHzxreF+pwW0KEgACNFBEDv+wrCSNOrRXkqROASqb/Z25KD9S3ZqrwY9UPBoGLJRv3T9tzRGR
g/Pvla+E4MbQjOmMyB9afTRecVw450T9rs7WkXVLwhFwRGVTPfJJXjo0X2hCHVKPmTbH1zUjFIaz
RSx+Pg68nKryIU3z3M92C7Oe7GONowOwqC4r0zpiLls0lSXknS9vyym+ERzIozwOhkxH66RgduX7
WItn+ElFKTaUQhUAFbzfg1Kt1RVhqIbazx6XxhAH1OzjiHbRz7lJBwGxA/tHtYdxQiFuSs1gfRe3
KDLl1ny3t+7lZYslemivb536azlhMGf0jhh+SrEvgyo1RKK+mXCppKxfCWfVKR3AboVM8J7awaMX
AXpESfwcvoBbAPET2I+AirelHPZbAutXqxIy72bSgTUN2Cu7rNK9Po33gYMIBCbRDvfTknYwHOh5
ZDM4kz5Wyrg+ynyUE9EZ48cYA8aCqvRVhcIBQr18liPJkysC1FEASDJ2wtr7TVKZQCYSwHckBKbG
RuMoSBi/oKL5OM+j9wDmvFTfkDL9jv7/r/YEfpczjFfZRzX6YxPrff39MUAIr5SIuPKFjrVXD1Ub
uO1eIGknatUa0MepAzzkZEJVezThe8Kedaow0yYSKayVLPQEsFTSL/tUltvVHH5PEKyaCuKOybBE
bbqfoBbfulpFVGB16oQ/BIyJDjG29UKXmVZTjQXeFhsUb6y2aeQNJcCqCDphnYdyCgKhyRyesKdF
M64DNqKvStK0SsnvQ3kqlYnhOCXJZVlpnJhuVZFqpGajLcYOew/rZsrJpTnMKiB9Iz461w6MU99k
rQ1Ai6RqaucBcijPiE0OyOhGEMl4i/vlEWXc8QgL/QVUeIkcfTcT7dO6Q85T4InhU+1+AvlLz66/
Lyojr37avCQBECYKYQE76fAqN1RZ7Y4TyqgMUbsX5zuiiqsU+TgJAh0CeVWCwrUcSUW1qSyLcN/Z
sF2a+CPU5U+qYtfa3axDO5l4OCSns5BWKmLYgsg5nwQEo5wBxkQ8hw7AT5eh5YjFecoHfYlTCC91
nixPqY/FIxRfOcc1b7UZ4o+58lP2rO9wKT10VbhqqFFSRfF1acCSsUIGyqBG5ZFHd693i9KspgwZ
4lc8JS4A9HuSKQPgHXsI7CSWUjGrktusyFT8pCwjrzfLNCOMxKk5c3KzlKLOJJw/CZkXse3PdOKy
gEsPMAbRgyYANkfq8EijYlz+8MsNg26fchQg5rMcHPBaxqT+cpe/T6qwiSqVjIrjj+XwyT/K6kuG
zL8maEqIPqfcfXp3bzjN220Lx6iYoD7bRDg5eubmkraeVTB1TlCX2C9CDs9u6EwQcZtKdndL+qhO
O2I/2y+gBw/gvbe6mIyWi5tGxFbv6KbJTd9gcab++yVCmBo5CQM0wr2ZP1iasZW6u/q3O4snnMLW
mI0Jgc4XnTMV5mIXrUghucl/8eEkCzOjpM2JRPr2y96DbkEQLCIgi47um81YxBK5Z2cnHodPFomQ
1mxuKA11XhxOQhd4NV3td8c+bTjevFG46yWfWMFTHuO+8/+4P2hReIZLqEZLNdt9lXG0eLaPKkER
BQUzJ2StN0CildcM7q2Q5Vsmi926NZzwPZQR+cSwAsH0Qv58wWS9U68kaOT3zp4arwgUPjZXETvX
XcW+r/z5cEb6UIuedKifp4bPSuF6aXwwgSxbFNPuROgvdAXmG9C8QnspxjZWqSOZtB0Ha8sicCD2
pgpi7WGgKVx2T2IttZUPTpbg/DUziC2SsxbGYG+GZndINbkoUcXZxnJ9NXbnrtEmZRX9kviy5IEi
iRZqwoP0PMNswnkli2TW8fnNGZelAj2ePIpSffz1c11RtaF0ehCy0XhLmEwPQ9MlAn6sEQq6A1G0
zZ+WnKdFecNS6CV1eatTE2eW1WzXLjycwgCTP6haMdoNRteqKpmiqsPrewndxP89mN6qCjnX3HNL
x7BiPwmEaPG9Q09tqQKbJW4kNoNH/SFCPsy61JRz9dmgE5+2iVOY1ofiUiAk6uaKuD9s/RVHTWJv
yO7pHez5tDVHy644C9GWalp4QYnqsbDB2xxTc43e87q7hSHLfMfvixKV6wVEOguTT0E752fejxif
E6nLBtdE25EExweYZbfVwhypKF8gQy/L1cOk+5A6VbY3c8Y69wfuNMEAjEFE6ct1FbbDzq78KnG+
kgpEoJgY/Mq+Z9JtRSrWyFt/PrwnfLfy9n62WWtUAy4aRAmmTETs7rh7AbjynX/2yDA06/9ySN/Z
btlyLSS6QLqvSJDH3Q9mmGHP6OFJAXUP6JZeormcLnlHncIpDcI1rGDvP2tqR5DNozfssMTpNOYO
RAZZIzmnaJ/G7L3NTTk59hN7aAB1+WpRP6o6kd+F286ljZb+icsMsXhG9Y0Qda8BNTkpQ2Wtxzge
Ip5yUlpDUrhnG5s/moulUr3IcJB/GbCsxksYLqoeSFP6hLtIUO0Ync25F21Py9Z6cNqTnTMcQ4Vr
C0TLjWy8TXQkxJTmNSZJbu/FK17xflv5UbhrMcgQCBC4gl2XNHCo81iJ3xO1Cic4qUbuoCzprOJ2
xfQjIYu3i4a4dCZdiEDuh+wp6b1OWMfCVXKkcx3HwnqdR/wYQ6kus+xWOLrD61tBD+nwHh7AyjJO
B+WEPDZvQw65bNA5JLmG53tkPzjnFJSOh6l121eQNI8MWWnT5m3u6HNU6v7HgZcU6OciJy1nfITx
A/U2oTK2vEuslXaIdEYOKC7whho7c2ilqYSg1j5/nXfXusgDi4dArQXKJ7TnkDRs9mZYb8GgGG6K
73PAgYPurLp41A3J5aNDUOop7qFNOyCE6dkaF3F6XurkOhP5+LeW3uMY2rEOkQ2lqR4vQgGh/FHw
LwpiSOifGPXxJSCQKp+qGQBqqm4/LVspF50r3gWXeXNYGuGG3QbeR48BfMVZ6pyykq2H+yzuXzxL
J3E0qqketCtHvDurSQuHz7+pgSrZwY67Al31QMn3Ec8hJSmGgTyXhMbijDky4uKkTMxWt9VoNq1J
99W+8n+ijDvi5OxM4ziCCTZgmBFrvdkH/CgidyWH5PPnvSZpdSn4mNi3XttUDIJiuECWkh3Fz3q4
lrUJx7B8BuexRc84cv3F4H+wYLQ4gAA9hqKHCXK7/wtWdOfE0aPUYXaULUnq5WXfyX4lUWIkonxj
aF3AMZFwcuPHuXIJbbJTW+7KkeC62IjtnAP9RzLVHBdKJMC97ZvQpK04RHAgByM19W7AM8MtzNpy
fWSap+LGbTQac0iixNl2xGpt9J0R/9G5KklAafLWnewsa7WGtO44OomKP+KYYjbEoIWwjDTTaKPp
e3VAEwpOoBfCr3Q9+gGyktnFhXIxZK2PZoZUYcvasd02v67uxGy98Sbc0zSNi4NYYI9YhsS6fo1R
T/MHeqZsr6ke9QudJUeD0V24goVvtLRhEQJ3kWp1RYx4VNcXbC9U19wIT40A2LtIOHaAEoQAcH4f
vLrbPPO4b1xemOAvAW+Sb050MzROljuGj3T9ZbMY+DnfH9hY/hgWLHYQugPho5lsmWdefBgKF0tk
In0b5pTgPmswbYgKgQ8YipJHzruPMhJTNxUr6ScvyTOtWpd8NZhK4pcZ+J01Zt+HleMoiIHPf6ov
tTfDckA9MhiPSysxrmvb0BBlWeEGxkrbghzBBupyuBTTp9B2dK4eMPDFM9a22i+y3nzc4i91gzLK
u5bcJmqunuWEoDVrH19IYOCNeMVt25lOxwkDZirFL94bqH9psBRYffsvCV54EF61TQOo1TIbd1pP
agcaoq0kJwESDOEl94n//XIIV/co2+7ovzVcSApXYdhosyntY4NJlLshbg7z2W8ExPSg7vyjRHIr
vXqfVysbyEj+AWgwyRDzfJ6uhAn66Ejf3EqbmRISMkToyHYKdrpQh2BFSHykxnnPkhy6od5PphWS
s4w4PRunPusgauzc13nrIW5O+dY1D9EyxoxtWDAhRvAOnfxG06bFgyguuPKk+2GXB4Shmw/klIDh
0vJ/IPN9bgmgwSZACvC9h3tyzUVKhvLwSldtbSTaWHqmx/pyjB6RmBP+YVLB/S0aPBRxhpubfpb+
7DB43mGyBGVzHVsUlkHk57IhTOm5kneNdi+iEagsr6s5JGpeO/tNValzvNmOBhLJuI47Ct+KnLTG
wMdKxhiI6eJzGsjvTwezZm3PY6fXQKxYyfwATfVoWAh7kH1MrZ18sfdszeLc+JJ5HcK5R/EPsNye
gJa0v/u/8KjVUGj8kkSWUobIFgoxPSeWCPPaf7MD0nhzFymMzCeU5YyfcT7b2lv1bFuZ57asCQ4d
qJiJNy+zE/0OSTjPCoobjvtPn15c9NBFzaoe5qdt0UJiI1rkmflJK/gPCsfSn9Gmu6+ODBDsTFp6
eo2pUazhq7kAgZNHdpa6su7yHyZtniLi975C8BBNfet1QWUyNNtL7tj9CA12ERSsyr7BLzSyz/V/
ZNQ8pscURPFU3bBbQ0q+yt9C9qVrHLkRsVRDEx1UoZ1Yb7j4HqGatcmmp+Y97E2E5C/LMIdMFZBL
T1kFY+fpBIOjKmulG16xBpvKE32L5olV8cO4c4p+Qwl39Y6PBhYzTi7Xl3XH00lJpF1ouANgps5s
mcMAP9vB8DA8toAedVDuiJ1pvxXj8T6UoXJIrmOOWsgSBoRR21IX4hjjhVqKDk0ZfJhbGGbCx48Y
TH6M/aMJ1fj9ai1tk0GQ0kdGCXJc76frdxQeT22LGm2reRY7V1tqeE0i32Z9KnSiR8TzHBg+sjuo
jlpGkQX4QovT9tWqCJUNtkQwCqZS67SjhftoMJUXAFTSAAohU+Sw8wX0rv8n6srunMCUqjPv+bFq
wfhmQU/nCl355GV2A09fXoTM3sqAj+3zGW6k0mMa/SoMuKDKxpGyGnYeO1tiDARLZ5s/NCs6jG4C
ZS4HQ3BioPSPp6o3zwOoKTo0nGHOkhCPuIR/HArauA8U4knl+y0oD6E6w6WAIH2Qc7uRPxTTu9cZ
mAuzuFxsYoqMhZoci1E//folD6KVakglf0tdqbN99cR3w5PJ+n9NXe/9gTvmI9AzeX9HC0nTQPCv
PS+doOJfgcaXPDhs949l3y6y7Lrqes4H9g/3zxH6UuutPBMY9IoQeFGrf2bXYwODfgaXRfYZF6A2
hL+t043HwNTGhmmQ4addrOp0KrGrma87RVSSrulD/XP4fGyrdYqHCayLzeyEec5x99RgdilHzGh/
qAT3k6cHBS17GjzezUdz8c13LboAj/0GGVexE9cZ5gNlZxsQXLxlAjZhik4DPt4728ov3IbsE6WX
RFTUpeDFq2nUtsc4QBMLuZaVPKJqaux/F97QcXw0/iRAIvMKEG7XJ+K7ZaB1QDOkATZ9Z+Rz22r1
OV514T4BKWlFAIvQT4CCMWuU/tZVVKSl7hgdG4fxx9Rfe9hgVlam08sjAh1EKrYxllHK8PgzOrNf
AWYv2FmQsSew/+EUsnbTnUSn52cmc+K0SSo/Ucpo/ibJRvnj/fmSYpTCiOXQgK6b68Uv3xBfD29I
2Lq4DZsPRa5b96LdAzAtvjcU+jHuHHpOcVJXLaXmRmciQM4QuehOvESHlst6xketvCR2bLYyaik6
BcHwhRoftpnGnoz86cf8yZCGjlIP8b9XRfR40THdlC4+N44C7e5H7M3EtijmN3P7S0XTTMoycpjV
XS/mywyXwc+6rnZF8hHx0fsCxQMfQfMB6DfK64T2uz89pumWNrhrbaZmdjar0w4ApZYSxBfN2Y2s
RTkhuwUsU0AxksEeODba9GphDFoi55tMSU4iZVQ3ahJY9CTwSa0xtHG6dAuF+y0LXN7qXVzWJo6o
mbvcMmVTBm8R25GsLZIuqu3875HI4bUCC9jud9hN9jfaMcAXXdTukBAwbemLeHSyLZw6K/VDto9A
Y1iKrSpGkb+rA76zdVn/ImFwkcd5XBKk5cMYjeMRYHUbe3p1vy5ylgNNr20tN4hGlbP+vAFBGdk6
xJU30qJ/iEI1MSjZ96T2pQ4Jzi6V8Y0j4ruzngqYcxDFMBygqTb+c7qGfadlI7PHb3oOwn/biaMu
aK6F5yDVsfpBIlo2hrzZMTp3Vzu/rmr8g3InqBOnor4RTLgqEswuJGbG0VPE9+b1AN713C/TNPy+
K0W8j3gnqeGrZ6aOG23z0+1anU54N5R0uAlrMyAndSlOIj9S+NBzcsBOA/meds9O7g8mHfPrmb2Z
0KXATf26Isr1PG3uBcaOtpxL1DVd3ZuBNme5K0H4/u7iHNGfMGkSTEtmi2T+ye9JNk5HNWR7GDNw
98VX+hUFSEr4w4K+7HQ8ACYkth/qcz6sIlgVa+T06d/N+JJDPEGj1lx3nKcYXCl5E1M9Vh/fyVPQ
OeEMZCuocDuGHOhqwLkBTVc2Oxd7uB6KmCIoNEY6L82/diwn4xf+cDAyaarCHAZf5zQFcznmXNGQ
eHbt4QKrvOyMBINIrRP3Ac6na/gVPvDDv7OCArJta7SLzhyQ16dxRF+98bEwUXDcYOvp94rc/nks
KkHmWfrj4wNdz+9hKvIsS7/EVgxZRwcET5PdOEdyA3mgeaMBdGNJPbJM7F1j7mPSmJiF7DRwtbLy
mUo1p4iFOD+Jz3zDFpUiwHUOIdbwoLScH9sZvYQTujrX4g5iTuyc4D7BeJwq4KY3YHg9z3eiHmKf
VkIPRXHpdiOji6dCF0w1lSExxTMadMgiuPZ1brr8EF0fC+5yZI77y7eV6EA2en+8aXMp9XG6ywLo
69ZDYmhDChRktucOzQ+8pX09OfWbKOjre07FoKKx1/Plb21faHbi/WfxILxwDQn/DMXJZhst92YD
c0Caz91l933916LZ39rrf6itLoTwmGyR6sXJA7Ew7J6uFsE723Zn+QTJaIIzYc6rUdpZZGW+p+Sk
WeaIPw8zjWJ7lRzHrCST52WTp0KpgWE/lbav3R9bd40NTQqEsFGtKicAXmz419j6LzyrOpWZj1XH
Um65O0AyQxitmtlsYZxujAxCZsKLpPdmvP10yeeqEVCuMPRLMtVEMnGsyv7RIVtVk3ksx0pWa+xT
AiIZ/l1ryERa6pCf9RajxXPUbbdOmyP2hjplteAy0fsGuCE6cK86ROyu8AjxVdPTBevv6WU9yQeU
BGnsidSMfuPPaemtyqjKraz4b8TpfiLp1yMWDnaoSA1K5803Cztioj+xJhMnKvwQm5sCMrpxQ5/f
86S2A9+U6tHzq+OSgSSD3mSzwacx7nVir7ktZYpHt2XU8K1cOg1u12kx1O7Y0+R6jIR8VDssi5eW
Mo+9a9HwjuISlYk+zKgGsDAyEiV5umEEGGxsNj5xBuSfVLHVN8p2Za1xnymzr2NUIavuxlrbqd9A
BZgVCmbptkU86cv83QEctq4C9bDAJPqLPlub5evMosSplL6iD5jQxfgoAii14tYWpI1Xc16NYgwn
jhxCQHhBNRDsVbGXdV6S7AOo548GnYeVCS5py8x9nWtUnM3CBvKir9ViEJr7NlQRiOvk7/VqpVdf
sFfYbXn0SdX+mINaJmnfU+U1By2tx7P+E33U2IK9Ky4T8NeJotp/VA46g0uZy8hLV9FiSfaoc5qd
JPFBijYyEeaK3/+r3HEGE6YiNTyvLygbnD+rXjEJP0kK5edEpRoOeoGydqiz8v5ZL6dnyaRxXD+u
wtdrCb7Q4dHLX1Bh4z8t+/msgHP4qNk+3M4j/KKUeCzGn9f449cRRXstYtKGXQtSl+Uyfqv405Q4
gfKeQ1GxNEOG54qcfPqWzT9P0iT7smmvQctGycMYJEJru2/jMFnRe0tVg22iYTDmEHMiUAzhHHWb
FbaX9K2k8oH48OVfsyGXOf5PynhwS55E/vNGgtZ47yHPoHAp1XcUUjp47gsTAg46tCUIxueX5ipY
JiZCf97RQyut2/Jzd8oObWTp7r748DV11s1SXpvfbdEYq3NhgKAsfn83h67K9Lae8BlYwAnqv/px
dZiHwfuZq2fmfQkZAa2Gafec8JOyZ7cUSdsQz/H4l0NV1GfO9rF4y0ibNLwIpAAN3inXzunC4qVQ
oa1eMyAsbOpikcfgfNtJ886A4fKgzL1NGfUwOVCBvQCFMLjgrlNWIa8Jq+8JKJtPpUDhqGNPvidx
ENMNwHaxdc+NPvOesQBmBV9vjHENHc+4VA1V9RH9J60fHFN0vpktvDoUn2EZGt95ft2qB77m3B5E
Bul+sGGF7Kmi90xBpztyity2xZvoBPK5D+gWanxQK0qpPJXn2/xZKa9Kbw1t4nKrXmjUZRE5baRl
o73LxCaZLc9hyHkXtRzWQMRvnHEDefdUAmxcTENBQ8f8ewkVtVfBN0EFisZ/MXI6v92cE8gWu+lx
NH8lqrWrXfVP8fve0hq4/8rqH18hvmnN1KaxJtInc6kGMFqRbGmp2E66vz+KL1snsyZySbNrsj9V
aRJm5XK0tfr/WgHUqhvW7SDomeklfzyH1UtSUR72o4cKMfsfUp/JazZFYGcsOp9+8xr5dKJY41mW
YpMUi7OnwuDJmDReLgGgd3DDQmSt4nEJ2k5V8xGZOW7uTIeyY/aCV5k2BIT/lV1gHslp5FVSONiD
kXDrEPLg/1sQgUn8TsWzu+cLpixPKVsdsBmY2J7ofWYNllDEoVqqV5j990QulKzJhZZOHeAbNKIo
ZwxiJCioXL9V3Ee/M5Au1wOnMDoIFnYxbN/B5XhtW5X0Z+wkjSTyfZTRR2JnGLW9q6hdCjg0kKUO
sWhdiLhoaw0qHvcDECAA5/oOLjQut/X4Wl+6ton47f2u1pgPlFNqlp0YqkcIqUkxrjY84+69NHvs
Wf0/uA3RMiSjsBoJXlxJbOAKGZ+exovxyzEGQqgTb6vQG8zNvHPoRzwWstH0TYDdvmC9kGehUVX1
rH+Dm4d/d5fGZYvswHiFObnkv421easgsp7Q26nXuByhxG2iFP1lZAv9Dzq+3WtxCnzXOkrO+xsz
62pBxoW4eFMG/zhRuyRO8Hel1GwKJ/V+pM5TYxunAx3V71Ehi8BH7i/CuU1F/gAWFCx0o1266CJa
v5gKSzBjV+ClTLTqEcvT1bUeIhXDXcpDHch/uyPVopbDDvyBf40928lDbRiiTvAgKFkey7C7h3Zw
gHEeAYnfdCt13IR9iP0RlrHaOGGgC6d1GIBgassFuyLFlIrqgjn8iv9jFr5qq6hf5AMQrJqhBd6G
4Qtc3iyDDCIAQ5b+dwkzgMQJdhRho3MPGRTBkrmDLsXch10SSMKyq+ZPi8/6+3g7TE/yF0uNF5PO
+BlROOLYIZb4zx07EhFAazkYL/IR9WlQ+5v6PLeCPbNaZ0a9yq6D1VyYuYWREQL7zQK5e9yGgSm4
cdAwgRkRikmsTJlMFvtUKYpmj2w+U47+KVMuqX8IU6dSVf4wl4yoAQfkfTIxq7cNPA1Pq/uJPKai
p1oOYdSSE6S8ETHaVs3/d+/q2Yi1lu43y6MFBQQ5j4P1S0UlqSVpsWSR2+o7SaYNa19Ea+D31xVY
cD3uieQLB5S7A3J7VxpQtssyrgMluTllNPgNe4NKLJM0ZjyOa9wfJ7TXuC5juzjF83OdS6CCQfej
sesToB/TMFXL2OdT0HBhGTBugXzpFDe4im42+PcfM2HUIbUdzI3WXo3FtDbXQP9SWprFH3B8Ffof
FMNk9uNATYqs1v413z5njX7wNXbECd9o/xg9Sl00qcTSVxud5BeyfKydsAC+bOXkFVHfdOxFkvFC
iJldeY1eDSYnejwdtOA8LHqDlNT3+aOm1WYzpkVma8bShNTX1JsItkI3wk1pSAP3N7nRE5TZWcy/
AOweq7sIxaXOoTjgT/kXNgb/xpxCT6xER/gPlI9K1iIxiv7NJqwWW7P/GtaLmzNSgrOvDXvf+Ls6
RoZ7YvTaiAwpxNV9lE/cY7oCD+3RBG7qh1mYVexEmT3LjnbBIjUECLVVw5V7nOaGZAUrtJb6p8nb
3EdhvBlpF8dAtgo4lQRysrwv+l302BjgL93RNbLxE+ralKZcyhlsQNpesAhaEdxCMGcuqtMzt6f/
hij67mESwBnyJxQ8dEkZCa36K5RB1Q3XLSm9W+zIVcIqcuSZyK7qx5vVpey3e7asWu+yPKduLKlj
FIVexZdClPogK0iY7DmaCV+FhF6Fr4shafnIqCikEFdfSvh8H4HLVp6ZnxHZi7IKEuOjy1mueUXo
WvXTKmsmuTGu2DKx9wrGdkeFlBYGwMxVkR1fh2qSrayN/cYo0euGonqNMjT8L8WbErdqrxUXH64H
L1m90RAhYj16sLzKcY2beF/5xsOYN7SHO8B/XrDbj5GhHaNXEcHmWz0uWelHEIol1TSjYwXVxYcx
kz/cJSpKhlTKbiprgEVQNbNVIYunJ5+9mIoDrM9fUm6evHxy9yA5kcI9pAFApISBXgs7oNV1FRoh
F2eK2w9MWST/dqS90Kuw1x8cevU3BomKqOEavE+Mc/1odP70gLcJ9yT1vwumHQSG+ELjmhOhNcf+
50qEC2lBHfQalAZsqL8Uru5+/ymGyv819C2MqtwgrKR00dfK1Ci3p+4bvWloExh3HeOZpI9QztKq
sM9keM6GdHUEeZIXYV0qMTgPIrXtaGWmqf4uBhCiZ7Ko7ydgWCl5u436LxGP+JV9bx2jSTHXdr0q
WYZz2a+OA6yzrcp6LN/WxR7My3ljTicewapR1talwRkfoRtlxhcq0HdOMpG9900WCvQaGZLInB6u
KPREihgdyaNSjaGF1PGEIClsvpmlOLVzSjTgwWaoWBbdqsp2gEoRn2ekRPSZjisjUinHMLk9FSEO
58KNSitQqhRdipr928VdAjclFgVmkcPKnUBHoeH/X//1rqyE+LYx99iaahVbph5Dji4JI5IVrfB2
wLm6rQUDwje+wd009YHsAtcQA9HYVa1k8ivuDSrkOaQec3WorYw3lmbyUWCJnqeO2maWa2z16bc8
UQfb1fLTCuAlql0VnxCSz8CfhBI1PHovLDGQ5fN7NlLgsYowv1FVdRYLOxhCzFe0ZFQ0XwjTqIip
Pfy0pDWpSWdx+nA+RTUiWTTxGjgtEPabdmhUsNWkzQPiuCJxzMkqfuCOcpZRf3KEPE7UnB3ka9iR
MQnzruv3A9tbeMm73w+DvJsEKaFlcuqu1J49NzCGk/N1Ac4mLQu+qgtkoRtxCJPOryj5QTr4DK28
lIbU0Rg0+xUNp6rUKiY+mHBhvlMI/ZK80cYUGgyVyqE8fEZPGw0nLYOrrLXBvwMzj0Gpy98sgH+b
CLFCmjphJ2vyPa1FWH4dXewkUn29Ty91EqglTRpGCjCcFIV1J0Xq4GdmIv8GKd0BfPRbA3+/yK7X
iETw28Ya3ihNn1NfBwnM3t+mHicz1h71Gg6Oy19al6usdE5cDSOmXKppfstekiwYzwAG1/ly7/Nd
7jTetRQNtqpD4wMDlKj4ggVX3XwFrZbY8C4jri1FCXOp4kGHY3NRvRIQ/+vHHvlPBoVCxjAFVqY0
aiUvTWy32kBgpxWJ8HjrFfHtFQKq9iLh43pUGTqIu4KYdg0wVoKnMssXZe6bZQvCRSe8eng1GX7V
49uiCLsQ8a/pEgFw4iPd0o6bhdblXr5IFrLHxOpzKJYLRqvZKVdqK/EwMqeX6TznDBBnqNxYnH5I
e0gz/6JlEeIhHnthLu7Syzd2/s402nqTiku6fxquFx/1gYKDbJ0ymtOvt+gvrXzyeEtrsd8o9iVP
R+MvReNfMSrMFYbOLKqMG/5utV/9WVq/FP9Aq+p7OE+JpTzExaoZJzXRRONULTjO8hdHh7vQycCU
rUeUHdUnnF3Sw5m9MzTHiuu1Rn8x2WeYcEmwnOzL3cgFuL8APdaC6OiKyeex+d0r6Pq/uMZCGPBG
uKce05a5t6/ael2fZyodhHiYZqXXPBoPzsIKlMWpocfVvsvQcf/8MTeBswrUdcwCI5bHvHtcAWCH
A8hUKjiFfP4RIn+nhLGT51/o5T0KYK4ec9/xsjbKAqYtrkr9PTvaGJezrdOuZoldOSOJudbTajva
j+U5oXUeu++yvzoScR0A30nJYB8hVrd16pds8hN8IdXUqAW4/qXzVwH9b7eM7iEscy6M5hXMmZWi
q5hKLT+aZnV6caEVibtPK89/KfBNk1JzxYoatXNs9aJF5FjHylvXOXHnRYuk3AeJi19o6JE2hRyG
9a2GPfnoLBLUzFWW1n1XBuUntR+cvaJYIL/+S/eMInATcpVaXF/Phinrih+dLhllE206MThWfxOZ
0ZivREgtSzIfzm9/Ius5K/Pf3eGL78PF7hPCqR0e3YmaSBRdGSyAakSPD8c8s07KSV+OReCYzlhN
3gTKN4zsJ1zs+RPRZ8ZgvGST8tEzLSbQ4Q6Z6ddW8PpkbY/MVnrssGOkFKcgu1KJcCyF2OOL8sJB
j+hUPT/IEsmS/F5SWkBGm4xdgfjS+80rV2VVjoue9yZjRAI+EinT8SpI7pIcGVeyU3sEKuX2UuQ3
J8zB1kXBWJOZMKEQiLFn93Pnff8Ih4/+w9Hmn1HvQlJknYg27ERf2liDFkPbrixs5T4kXcADpjVt
48knezHVtymg2t8KBMdO4tJysZxYB163LqSrjGHT0yO0Xk6S3PByMYIxVB/MBe1x8c0S2UWg1BTY
MaqxL0SwZI9vrC+tltgdtMFY6iGkXBZLCUVVeycQ/iZjZ8bWFpS4mVXmI6Ntz/8eBkKUeDsYkg9m
1LyW6gFI3sEXdn17bMW7D+l5iwg+HDSu9Bg6O98MGH/3BQjpA8m+UPd0Acr9eR7ZGV2d6H2OvfZ7
H00zthGiX65Z7aSfy+ti8QanluLo9UFCR+ecJABTvpHw8EQDfSxbke5r06cZcUEhFnwtt/6G3gOj
jBiVK6gEScu7gEX5/m3pFs0TTIAtU9obuMcYcJl2fPHUcGVLJqttEYintVyb7Q71mIlKLOITNow1
QUpTyCVgAEHhkXAMwalBWGWXEHMxQxsTOHzPSgAb0zGD0DyBTEJy4yVkGSCbdivlj5QqvT9C9jCw
6UQ9dwuS19spI3J4KXmBgKT3i50KTW4lqkN0yTeWzkOWwO5VOnpYVK9dnKQs93UoymcJOeZYcq4v
Np2VA5+OmBJ54tGb3ghfKGp6xX8f+cJHE0TEn0Slte4FaLwQ19rrFVa6bwObohsykCy3khppk7Ou
j9PNTHrB+nnmpeOL93LPfznn/jLr049FjcO5V/hfbF+iMUIHE1oBUjTDGK/XDXmdjhA3RQOHZ30d
BdRisoKXE8rqhoQHobEMOXgRqA/MG3+KympUV1HfkKd8K5jpbIyrcAYo0PNh5zPPhYBDiQ1lpUXP
86lFnGSRYdtZKKCkrHCGtEoEJ/jOrs8NrqVQBuO6KTCUK6zC7n0A8UNsuNMGcUjyAeWaEkoJDN3B
LoTebc/LKE5ZsMYTo9I5AlrRUFGIteXAphQzSumyBeM8WenhYvpOAC07IFkpGXY7pS5qP2TT9gtw
LwjaEx5ip/N0LwAssoMA0DoclRBR111SJ33EimeW/EJ+KPIQoM3h9XTRB5GKuYFm4zl6BxTx6bz9
VubBhXdgkHaOii/5S7ygIS6/uxTkiJ+9nG4NRXmREmhXilPImkOk0ZdyPd7s5vgVINFDN54pvTFl
U9pAOCaw+wCMYGIwyLqK+be2MJPhLhkgDcsE1XWhS9D9WUQdnLIPuJVcWSQ7AURRLM+5XmJOwuzv
yqrW0isWRtcIsICCaDpWGLQ42KG9j+TA/Avy7sIuH/Ipj3PELuamm331nwJZTnDnXVNMjSzEz+Wf
0IFGrN+lFUaRVG10U4PQvNU4lIjjd8zP9BEQ9dTLNnyV/C6tdByvUpa1C6ts0Y9KJCIC/vvXNYE6
RGHp7NfQnuLZmLTYE0ZQp8qmTzhzTpTKsOwDrnb6Qn0WynC97BinxrjvToECTAr0m/w6AIkmQdaV
d4sgxn1bFadDCZZXm01tonwXFPCY69shvx/Ul3kuGJkW+py6pDQwk6fmUztmnXqHjXS+ihuKqSVz
cFoMeff9/JXXtBvevEYqeIEkC+8r0PSp3HjaOc0MYuOHz5X1/b7uStyW45KTcLxOnAVV/5CzPv7x
/AFDna9N8dqv5XFkxrYi0IvrwS2OOu4uysS9oheM2N6ZKIOuHC+NA/9aEHSUEi9FCK/HMj5KZSAg
Jwffb+zP3ibjOKOy4gxTJ9TYULmjp0Kqj9gXMag2yUfh+swtbcoIL6yzzQHvS5NOXi5PDo6uJi5V
JMrph6ylUMJPuuXqWjXGAAsyNusxR1tgCuc6XzpbsIocS47cLyzP0qYi97TM83AByHEMJLyYX80T
L7QgB3C6rqaO3HEig36MFMaPqm0Etecy9oWrBWzYddpnMxg8DiyBF3K5pEwiR7rEiLVe6iz/9IeP
Q3Mn5685LSbq1J5N8+YkQq6GA8Y6h0RMsOhtfRhMvelM5UlSH9T8OTXnMU9tFljxnR/HQdvx8JGS
7b0e7vkkGkOlO1fv7PTITv9unMCUHBQS9DyOg/3c2nuIYfHkLRvA005FOEKOQDDa1P7PaSIrr/Z3
43b4xqG2zrGx4fEseVAAt64yO1fIFpiUH3yoOcKY8PnTFwWoWmvy7KKBBUGp2lw0Qubx5WQAOkaq
rC4QV3R4byzIVLFyd0hILjJaefuuo66N/VLNcRK1HvgPPHYEW1+8CC7rM6icklMXTZWHPkaMQDDb
oTrRBpZA2cLPLt4bBsrbwx2OBdmewx+MjIAeiNvkJHlcebwvHTGcPBfVNAf2ZpSDE7HmKfjFtigm
yWPfwlmzO+6+n39luLbaHGx5ut4K0uBlM0kTNy+Pj+9B7Unn4JTau1VSL3rJpIJW5RgYt1edSdUa
0pjDF0DLlatBOOigaDqMXupTkjOYIUUslNHMusqOhitf04sByLXCnywDgyoQ81M4Amo2Tx5PYFh7
LHpsgU63O1wZjwroRQ0yhN8kzFjZac7/kj69OQ6m6fZEsZh3ChnNmOdTwG00fZfpg6EzyuyBVHO6
6ImsLSbsifVyAnJczBlE+bHOW8wnoeXfusTkR7CpszeWqQTdPnZHfZm9EiXEbmMlZ5ko7xCI4MJl
BMKVY02EMGqptGQKcwTBk6zmdAJYom/A1kVi1WNlB2LTOoc7w8mRjBbbv+6qVuQKX/GW7FmaLNGc
V356QJm7vg0ubFi/ny6EljcmIZf3C82uLkWLcN7HgP5j/uWzTM0DWNO4G2Dw16iPytGZYD4s3Vro
3yThYhj7o3r/etd4VPKUWY+kQfW9Y4TaiLPq3pIO6FELlzddyKHnm+9BGXB08Mur2n/lhFPyH7kU
J4/tOaR/Q9FzqV+zayuW8GTMxPX9pPgil69th+8oggLs0UsExthvIouSok9WoLI/FaMnxzCwb2oS
IhQeEiVdGJSxZNm0HcE2tr3lhy0z0Dl3JXY76aL289aigSKj7gPYQn1bzASg0i9n+qWKRZIOZbLg
vntFiVBtkjSAbT9cuVDpNEgyjopXcXAKBeZDFeelOlxECFep+XywUXqIPQTgr41zPLZHL+xQeUO1
M4YQYpqvAC60k7cb7A4OL+V84Czc2sgg0XThjNwJcon2wqm3czgjA16QMMQ6M7haP60cWDR3Y6QP
rNfMx0KUIzNm3OzZKIJn/UkdOBtUKnRIlK4GP+mSr1YnusToUwjp923vGOlESUwbdTEE8Qdgqu50
ZJpxApHqZk1IJIqyS5D24RQB24dv8s2g6GibR7lGqJBCySCAEhfEjLm3D5+4axF5cLNUzWhGEwid
rqKE0QiRPXLJQ/8i2SIy97qXIDfogpsBB6VViESkONnpUkjfFaK8HECko3pcCwjtu9NXdAAnrFzP
t5IKEkN/znBrlL450SOgh/C0hFtUeqPwrFe5+FXb1Tm7SxiPHWjG9AgSjkHLmxBT27bEiUBGtCs4
3CHVuYdWz4WuE1TZQ86NTLZD54xKSJKKY9DTWfmCFDWdjkZU5C2809Ruy03N653w/szyp0TGqnB2
S2DMAudLB5DgnNPUS55N7LugfsmuxFlyJ4lH8BtwVRwaiGSMPGQAGRnVtvLWiIn+tk0Nirv2vDDm
AloTRFdHIDj5/D3XQiL7DCb/UJ0s2n7FinVmmZPB/49DCao0bnuplD7NXuR34pdKk6ZC6ucIs03D
0SQxte55rhDNH5b1XYtZnotk8G0Andiq58LTR3pxWl1w+uSScHAby9G5rHr1hCSqfp2zlSRscYSZ
hxAJwIAtHPtMO29v6UtpFHYcoHls42/hAA0ij/uRbW8/FOCJle2wU6yCF9sc8u5xH/Ar9an9jrwU
r2UzDGpdRB+E93XVF3NqrKgWhEqmsmg20RdPhDQwBp5yiqi67QrTzKimpdm3AghzN01MY+ksJWAq
B9nXio96mgEzRak1bJcKM3tIcB0FOAJIPLGa3thVlTc5nKNazFUZp5BS3Uu8e4cZFvQQyrj8nnH7
cksy3aHX8aEFJa/L+l6uXOtXEONyURenfB25E7VtwqUdqj8z4B9MqZvfwXnH5o9oe7vcZM7JAavs
1ZzCarMN3I2RBpT25irmoGczXp1tj6A+qG/QXyR4Y7BNEEMQizRLFEQepcriMleIE7ezbDau5F7V
hQHzNOD21tqqf1D6XbQgjB1S9LJ22jfPeH7Eqh3qo+86CJUlkQxV9uzdB/nfXuqGkVih/6S/GxjV
BN6dGv/JfYoYZ86ue3/Bmw70BcNseIjIeIJN+6u5IIn80OcqVU7NNCMKYvmP3t0A52wepoXeaXYL
LEeqsJ2a5pnUALuXTPANFasWI4zq5RtCP0yDEKSozmxajlMLCYm8BX2jTnKS7JbuQIiobyfTcnuY
6klqo+2WoZElssTK0j9F4D4ck+xJXKsrYrkDiKhLyu/n/miiVHJ1d/fQP8TOoh5wfTqYUmRa388b
gdIvzrXGzO0AayAekQQo7DJDJ2Vn4g9vajDGDvo0JZw7Y1fcIvC0vev6+/BplAC8Z51fGfp44j/A
WRSROtgr1JERFPUyWH5BOSMDfVtoV5Rhxj7HeM/qn/9yvGdYk9v+neFYlvf7IWqPgAGBFpj2rCb3
q/HuZGD7b8bXRr1iDowPGEgDBZI7RrWBGra/oZ2b9KuZl/3Bwdl55WR/osMdXJBcA6hFJovdg5JX
Aw3aThZ10KGBoGLyn5/Sm1IE384MqWtK2z6AF+EM4SuXrszjrsqxxe20/waOealdeDV+tfsLv7Lg
hPPTMMrGuGUE/0yTAyOmVXdio6Da6gxKjto7DluAGaHiIXo9mqgKnSDQ9GbXbbcAVKYEWLedpTa6
WOANNdGnw7zuPrlHG8DPDb+z7CJY1PUPlYULAzyTMo5yMbmpqg6Kgf6Qi3ruAWJzHRy13jLqKpgb
oCEON0RyGCZ3JH5LK4t4ZQlLz40q8ouagD/URtpaqYtxi8LZdh0KZllbo7nJoY1R6CK4IbmluaGc
fD54H42x8m37aTcVwkFUHQVTpV0FfSvAOAY9f2TU8TJNDVW+VK68sIKEwVOXJ/SDw6jFnTL3I96m
rfBsXw53sEKri8PFHkqZ1T/xsD0B3VEvVng8Ift6VkoxZUNUQqLFGc7BcczzMpL2pRUAyZ6xmCgr
07LpURlLsw7XcA+3uzOAY2ZbK99NIPSai3H7elXFVjbMlroKPcjw/FF2DckQunU4kW0Sc0V90pWn
5GqQN8Jyx7yTHg1ZQb6Eouo5oKKnAp5MWg+wup0RH7Wx4Hj/XFSCXvlM+BjKFd1huD5lRvFsagEr
Yq+TM0QOyKqRYdcMxEq0gT21Fb5402/aDHbmaRVLgDjTwWaA5wlKLPzup2HLkM0CKhlPnVjsuVYK
ZL+yv5S+abnODU0QsCCE351oDQWbAQvgFxiPxzSKKBHROyj+2qnQMteQrjZcHBH+TKX2+9LZz8MD
+r+If+2IBCBNUNoPpcSMfQZSVT5MIxFFdcxhMsrStJNJ/5Y+nXqyuBzDeEBPprYhjzh6Nxj6/VT2
E95r5xuDRNYudG6LcEKtCj4Uc0Hr/uJfRGT5srrcKo4rh3Fw3Qtuf2ezL7bwgeF3stGwmLNnfzZN
6D+T4VqXU2j9KRW/mdPuIEatGTWV4bfd8Jnu3AI7yNVgIvoJ1Ca64UciQqLovuhCtdv5Xw/M8IT5
/pop2AbKcWxtN1FVk0Tbo027b1x+Q51TysEFK1MTQJqQxZeoGY75pe4NPw3rUyDr3gVxaIh3zdJT
uR9LD0DfZGNffVJdxNZniYe7Da3q8spsUGl/U60XN7H261bw2GA0QF62OS/K6eleQlUfmy8JiJmL
2hZaQB60I2kI9kduiWwtyS+OqcoQ3OhypflvEpH4NHTlyDB9liL8CV6UQqRs8FQdvEBEAAQHNvS8
Wd2QPvDJrGUZhYbtHmBLQvii9bv6N9fl6wqbXCy4gdg4FhPZAUINB4yhvwG/fX6As4Z/bbTglSqS
4uQKVRUTMssamR52isNKm/hsEwfCv1U8cLjn16lZpn2hAr7g+2nsHtul7jv4uUgXZ47p1habjrga
ZVt5N+d/Cxixq/oOx+N8gMIFvtB615u+FspygDHnDucGvyP8u2dTIfMV67qeLSZ97ukbw8TZosKf
90uIEX4NIMuC0naeR2ecTyZx+DIRgf2QGIfNbYVJfujD7NrOpaFlWQrzjXEciRSNeNG0LQjx+9CL
xwDveAm+f3OwHkQkAVjdOkM4rRC7Jj5B+0R8Zl1wABsZMIe4FBbQiUZiUdDm18RL6uEh+f9vIM9O
Q7R+xi3czDmQRPIp57B1yCsLutCfOyRjLHX/4RbeuxO7Yrdbqf0FI+ZP0SbmLg+hkVEHShsJfN2K
iUW1mE0UibNsosSy7/ALZREoqXaF/rM+1/p4JmmNaxX7H/X6xGuufEGm1RUbytWCYCvv3MDqFPt7
JTbvqsCQc/d5J4Nx+oZoptvXwnXb+SAEnNBVcxR/HDH1lZZ4c6O9RChN/yVM3/jf7sanMqjZS6mU
ajX1fPzNwzSznBfPwjEweCv4DkaLLMo2cxgL+7IkQIgwlu5M1A3XtH0tCoslEByvwHltCPPf5Mk6
J3X1UjzZxPJzebEoZe2EpMxNnz73LUDE+mceBADlEj/xwBe9y0rzVtMPfkHYFwMAtM1TS+lfwecP
+AzwO8vBl5GawMEFzPrF0ZBbr6L8tTN+/z6NW6qjdlEldqgaJYP5JnXXZ392/+aA3Gav0PPWOB0w
FaZU9+EAt50IhAuQASCnhOhRyC4/NqKkmx+MiskJlZQB8pHLYfuCeB/Baqi1NtE7PshY9OS+BLlN
+BFBReeVCVNbCRt8CSHCYgSZY84njGoxQotNvizrcGDsqWLibBvd8Uf3cbYGDA0nb4CwF9feO8Yo
PxPpvq0Jrm7hgyIKr7XaTBHRGbYI4MZq+C7XMRp/2AFNgzjV6g1FdtPvq8Llo/i3oc1LcIll2VE0
R8a7UelYAlXUUyavGlwl4y/OJZ1/o/qXvkCxG/vYYYfGJVlQgWxx5oHDPIRxOo5qgecnsyhkSRvP
OQiI+0HYlBT8GUG3G2Uprl1gJmw8MAtHtdQwp7uXdRLZG05TYjgYm/OAfC6whsaUZw9gY/yrgPW8
+8y6pyFOxx4K+AGv+IcgNWh28JR104ECi2SmXg575PC82V9NULnEiq+iXcJ+1wm6ECXD6da3G4rw
acsiOziLc7GRLDedPDIQ4k+K61jf7p87NRwQ3ESJUoa+dNYipxzHMWuW3F9/2LPUvhwHYuHbyP6z
f9kHFe6Re0N9nhVyzbVJ7+7GaWsmwDJJDEuCyGaQTFgqd5Ss0d10zUdydRNUdYoccAxy8IFi02Ev
tnlJAo01N1GY390sInnEYU5wpeNJtr+mYHqI4iNMfxRrBKQEijdpnRCBJwzdySOdnFKb8y7I9rgr
GvIJYpmSKQFMw4/rByXS9/GWZQRPEXLySNvceF+EWn6BeKDaLxThXY1zIlatPwwd73DHIaAEn7gN
mCfi/9psp3+Mh6roo49Eo9ETsNIUa6o28sIF0HK2TWdomcB2cNadgM6+7esdrVNrhHaeDORYx86n
xBJM2kyevtqyKzgmQ3TQJPQ0ULf9xx5MzrzTFSngPbqm8bgR8hpw8HSCCYX+Gmn6DJqbFHls6Euo
EAQU21MFznu+TU2XzAQAAd/zozDF+H9fFwyDFjOtfjCqEh06l+hlc9Kv+wk6X7yYiMGbmqCUGqmT
IYppgaWHeuBINMUoMHO86QC3P4+RBe3YOTYd0C9M3+iMoDDoULFFFuABr+x1qHKV2JxfOe0oPWPC
lEuEQFDZ/zs4J5sXOaMJFbDBR+b3qj8I748hMEqugvC3c72IlHS8SaD5vxUVSPB86kHg3nraL/a0
mCiw4usfUULuw/uKXncBSI+90czj42MPu5kgpmrVslUqgAHSm/97vfxGzG/BmYCMk53w1MJ+uFJV
gn47RQD5Egm4ZLzxSxt93pZCWvuk6LrJtdpQ0Wp27YsMSzeS83tabe6Gt93P//7fD+/KRmoh/TtX
cK/SV5voA+8BbhXh+KTJODiHE/d6DJnBaaKI+kbwTKgw6PTFuWYWhugPZeeJo1l/VZ5r6yF3Z8Oj
NDrIAPa8x5uaP9y2HdIFvxl0+HUtphY5LPFKtFieuoqlr0CIVx0ZoBc42h1Uv1LuhfOGYeJpIGPK
djC3LXRrCs5DviRzUccQjp+HluwXr3BcCGJfScZpy51clxn8phWb1qDoTgWB/d5L4i4/hIdwf9VS
pETD/bev0ZSsPGg2hMOpoqWXaua5nTvw7uT5QeE4D52snD7prdpmRUs634ORgzsB4QF6xLLLtTK0
VcdGXhC8NL+YKU8Pkm1W5k2f5btnUxk+D+pMVwIArDdK9hacRLyb0yUFwArMk47HN5g9FyvW9CVI
XFs0RZBCHmvQGTjlwAbwAg8w2nwUYcnxgt8UoVOey8n0hclKiGRvebBhvzC00WVGNGmsaq/9JhUQ
TWtMLPzpVsgxEf+fJCaHYoPriJNlSkh0XDUdmGGqIvbABggmUXDkGLWXedenBuMjyMPORgvT5RZr
8BZHkqcnFOzqJrISW+9cTIU/1aMmDMJa4RJ2zwTPDJgRzKqKyO5FT7A2RWR/3WPaz3OI1X1G5sFp
7Dv3pROx7LJWy4p/ImPZIItVVrf/T6uNSYIYiPzLnl3kn/U5bAAU+uIzDeNkjD/mJoEvmKSosrE3
Ok6fjys89j2koIGmxI9sawKdOy9erlcQkw7WvvadFoJYutGPj2639Z28HnuwMVVOQfF86K8BbFJ+
KRHBV9JhWmx2eGzDynLm+x6pUI0Fp7OCTjGJz083iVzQ6b0u+yk/lXC58juu5VW4jf9PuGT6Xy83
dZFaT72DJlnQGDuuphy3gX0Oup/bXdi7XeM30F+cxvPM8yzepQI4cJx6Rrgqp1iLCUy2wY1caZd0
HMJjTy0Tg1TqvQabMv0Jgeus0v77lhs+hFEyNm2c2TpA3Ckor8y9bnGhGp8NFsjU9996wiZ20iBP
ZM3xwi6yI7k7B87TYaLSPStPhqRcXfHSAQinreQxy62nNW3qu/xinPITQvUZYT2qJ9UPH+dWZJv5
9mGO1GLdf/oIVdoiu8vEvQ1DOh7QbhMLJ8QVopTiJWIch9ZYgYkka9TfVbT2Nf0EY+dMsR6ClPre
Sppwjmwh6S/INBR+gahmRILi9ZxckqrmXPt8JQB6Mw+BnH1wvIa2Sq1lhPWGSawpBh3LItyHdyfl
G0wsgnjF1Yc1Gjq4wfPse1Nw+nLhZm80cUUa4oq5a1dL9rM+zxw6aGW62UyYuVvzQ0IQc2CV8hNY
qB+io2vdnVgtX4+xn+pcP3o/m7Kw7URBhaSpKdFyy8ZRP5U9UgpPcYO9B5CDsLNrTfkMC6e1Ox8l
0vQKW0PZwntA1xY6BB1UUwNmi/UEYth9fBbo4DD7LWH4Rsn9uZXRMdvzlt1FS9ruhorkbNZkG2Q2
zkLQCxCzl2SOngl1qYgh6GC5V4iARFrIyFqRuXP4QXqVBWlVhUJjuXIubz/0CSLzEsJAu5dpWXRu
ucO0m/JkWl5nJWNYbyi6VgDXXTwilqCNxRxZrYKTz6NlpVrHy6V11xtS1nSeRZqQmxFVMj+utFz3
aP7is7UMMi8gbRyYaASAg+u21/BefoR2cvUYQ/iZQHhYd1/QVYHAbRqM+MXJixAQom96U5lXUKMS
ohESdIcU4R41/9ExH1paGlUl6xLcttax7PNWmLaBOrnLk9TmwaDxf77OD0yMplyVa88mOJWlGsMI
NCRIxPOWYccMGh34kFmh2QkMChaHxH3xf0PLUiAFqGucO7qUO0OO4uy5ZFe02rKh+B2dUnCF+nj1
h7HKiTRWlensjpsjnaGj8oXCceWSqnTOSxRepW3JRqApt1H7YwfJjz8aRxFrfmiAQdD4v4XONrWP
7Nj29wXZaGLsGsopl9pHAKSjv+wyNGIqSxY3E31SLIZUvJyk3Le5XK26TbAZqFc2e+K2YWRmOzt9
DP6Ga5a/zGVGAhxcWa8jd9KGMdIuplOlDN5kOB3ZNCkicMTjleFJ+g07oXSNP6fNrIKPZmw7hSkw
DNOTFx5pheb8MEFjoJqu+SLmR/ZwNa2FUp/6jU9ePMDKqSMbl5UWvB+HqYqX2XcnfVAR3K3sr61c
NtqCHwaYBBgtunXaQROyhfe+vSMlVW8U7DW9XawOCE3D17Wj0DUdOXU2DidHldMGEGd3XzHeiPGl
2p9edoXUUA8J6cOwYoBaLkRwtfQkFL/RTtQ2uHk4qvWq5jwKN1rxwcoETtNxbunVH/hADcLg/dp8
eJ/aVKy6kG5gXZQpdD44VuPh5jaLuXG9fimmR9rZU8yvSvecVqoJUbNaK4hAL79wGPbapJHES2oV
l3sNwTCEAatHdXoniSaNT53HyTT+sP15BnpF3V6ekYDriAO3ErENtZB1BDsLJC73LA3P/tptg6q6
GDntV11Qw1WzsI/w1GOwLHiGyTT0siEh3hRLSWBnv/j20K73in+1AF1mBmS+xTc/D+sBGRhIL4H+
fizyKAFBvaclRSWfgMZozqp0ZCTUllYrE+6c7WX8wVmWxLrEw04kAL+NGq7lt+a8h5fY1lrRmAq5
jIGbZxZCWuAEuI+7czoxP+G00EY/SDQrbaCtK6Bh0bW0LP5KCRlPlqLku88n3CeZz/TwgzRYTOlQ
Qeb4f2BTJC16sZYpXCjWcT6aXudVnwZHEASmiqxZTVqPHDjtRTRPB19iL5l6JeMbipP6SyJp9Y8r
onVlrBEqzwRVO6atuWrp10u+3dQUArOE5dT71vsAjsJR53N7eKzC4f2LQk/DrcAKElgxIal5AwnI
6ANSpYjvZ3yXM7xbelYTyuAfscZRq7weZkgXDm/Ff8YZLy9KcdZVH8esmCe+vP7daTzN/Jd5DFgh
rxJLNfZYgdcgFhBqHfUxZzkfL1W/807RN/QisQkDhUdfEUwF85qIHDMH33rSonEuVt8pTKwTZxoW
gPoT3pVDSotNmATF+2mOZmmG2jafW9Jz6gMLCJkb/B2p3nWIVZHROKy4HO/dhU75lgg5AihQz79X
ZfEcvqfkLHNh8Ms51Tw+/gMuV05yNS0iCTb8aDNqsxFiNrBulUZukpK+MG41yNamfCbB0VyQqB+7
MCJFVQu6mUf+9AxmX8BREUGAW5r2FDizZXxpR83U3DBUd1F8SYm9cQgxYhu3jzbduUXJgom+CEZH
/yZuvTp2erbTEXzcQB3saJMaHy2tp/PR7liYya3qtkH4q7//wBDvD3ameqZ3vH5D2mmEcCYd4F+b
kCC9HLLxyNU5bgd5vcwtkybZn/Wz/mDpyRaZONZ2mWxJPxu6fA8vtRqepPJ4537ED1lU63U5V6xt
wWaTkDjaeE/6bZTLXCtsf+E6uIfviiDqybJndlOMJlAP5zq0CSOoqUAnqw1ALt26CLUl12h7W0TC
viP6Ty1zzgELMqJ0lvd6TldgxsI3ZE98i298IHZH62o9FwWp06fGHepULZzICNCsdnUOKIMpVvV/
Zo0yEhqSgeEYOVfdu5mybDbC4t2sCq4gZ6QempkAAEqMMEn2EWBbEVFFdAI10cYM4RoGmrXgQ861
YwzIGbFOf2YusUuHSP7nlwrgLTihZZEk/kef5KTMBUBZPftCKq/gOWWJp2csksqwBCmfE25doSBE
xHMUh/NWYInO+CrnCtn+2Cs43jmXXc/a0zZ78sEWiyWE94kfaAi0MEepVBkZGh/4Xjrrmdv2qZyb
QG3HP/9stIPbCRwtrrqCANMg1dwgUeZRmb21VManv1PuuHFACCcDCNi77t0dMoCsrGEJGJ74XX6h
cmMT0+UpqkMOzgueJUtx32HMXyKuOfjvL6shkw8bQg9EmJyyqN8blQnatAC01L1UHrSehlGtmZES
MzFyo45VKY22fwrq+LB0htTrmZe5vD3RHSSruQ7OvhXG08r3m4pxztwIdIrQDR6jMXBgJtkQaw/5
st90M33pG5WxkEwW4gOul8w2DJcejccaHa220e2TiL1iKBgYGd8TYJwO3WIn/HLKRnB8DDN459zZ
UOBm34yppwYS22A4aFJpSGIfKQYeZ/hPEQSmTAb/haui7POfT8sD/zBMxptfl7DRqmYe6rqb4Khs
oSlwaw464yBdQFlEuYDmk+3g9U5nxYE+9gMcenJswKYtAVW/00A1eEya5lXWVPrIc7RkQbHjL2zW
8grurrRw6yl0XpDw8dkaCp9BXd+XwOVNwe5yfg2/Z2ner1tMqUlnuOM3r2XiKUtkF+uEsent8/PK
MW3DJ9amswG+D3Qx5R2BUUVkBLQ2uUvaaSM2e+cVChys2xI/+8hnTMZu16VQzEAF6ifDxN2jW6xm
DD19reajPdhi83H9fkaQv5+XroO+dkR2PTLllTy9z154/rx8YXP9kP45hkdwqcWmIVISHvSFZM6H
kXMFexgGHUfHBf3jYvNK5+JLLfjh28bW0Vg3elrXVd5IbO+HyRNSbQk0hijQ6SuTkOw5GAleO/Fv
cCykg4zleF2w5EPlDZb2cpRAjC3kKOX88Hd3Ki/ew4k+hZ+zp87t/BzC5Th5dKeuMqxAELCGGyix
gE6XrJ8z5mgI6qLLjzsn+CQasWLvuJDCd8C3OGdwSpub4NwXuB0eb4UkObLcARnLYZB2TqB2a/S2
ZAxU7RfJLyMF40HndiaoE1eg9RE2j4LJx6xRxUGB9DbZoyPPYITKrVHwu8QZJFqnAe1IlxsXm/sE
gxmxbg/q6JmVPgc1tgoa1P5Mv29ERn2sbJc0FWMS4BgeV/JgEyGb/Yd3xctxyhICpcK+T4V4Fbsa
axWCqeL1P+kirFjaMTxJh6fOC91oprCoiSaXPdWTCbDzHNaQA1t2vddhRXTKe0pFfUJ4zHSV874z
3fcLD0/X7PnohJ9J0lByF5ECZTrXXYcWodNAHeM8Le8SycZaXBGZPlaUjY8cX9D7HRD2HG43ehHJ
Kpyib7PK2/WZjnVfdg1G9co45WFZAgluvcxP382wKxbgVoFfNSyGHMZnmCYxQHyoXwBBO5uRTpab
2vuHDdxwaXIZslPBjdqZWQpnb13FTNX9YhAJktAMqEemMBBzCQYXN+nx4HNGhmh2UXZCfLQf8O5P
COcs9azq2UQuLRNJcwfu7m91Ip1dTCTNl+APhgSH16TKkmU8xa3OWW+Ujajn4otHAAxr47UlewKK
P5SqpmNBmRuRdkLiP+GafJOHwNfCeabMsciYmYkbMBZxgmAUDHS1rZ7LNa4KFHTl3gjwFtO8gpua
WAP+8fkU+l5jIZN7r+UZK50YF+u9WyV4W/U+iJPC5gG7SrkD2sixPGk8wVVd20aYHmqmdNMqBB/Q
I3QoMBP6OYVRLok+qkatjnV7RzBlbd7BLKMElyNlps/jEb4LYFYP2k8Uo1SCsoMewIRzBHeJ7joT
a0ikr4b2tpptuh6MLl/IKA5zbNRbGCMkQ5u5BQsz7dv+CZvMgyL2h0Ys64HRV1x3FVmyrS4Q/zY6
2/eFtPX3yLnERo/OAxG0JRRxgdhQVr8oDtHlNV2ELM0A6hsEI9ksZGN+ttsBvEoTwS4EEQlZJZOa
veRgAr5hJrwfna1yvaNm7wJIjOdgRxhLR8mYySNQNSENhqGQqPX+5vm3SrG9QtqwmpHH4B8q7RUS
Vsemc7CJl61SHGWwHPIShxCVI6FxMa+c1T2Ppvfy1U+35KBkWwWkPInekL0DsoTeukRAvdR0RcEa
wnUgpZO+dmS6mOgA9p9yHydEVN9PYeUFyb8mPqUbjNq/zl5mQ2rMQ3NyKJ7QbjWEtA0q4sSrf4O2
miw+5m+21iCsUqf/iNpr+vOYTJ2fyOcEBFqC5oEIGRYUPaqmn0pEbGhxfh5up4BLOPMXU9DB+7El
u5iWJOmz1it1/nA7dksAXwqiXkQE0efSFx0UHp8o1nGyL8mOiGmzrtCo9f6Vn40aPtDhX71I+eOx
nagGYcZ2F1e8mOMDagZI56uXSPcsASHZV0zRB1xY/bEMj/QNHRmNCMQ4F2t1sQJ+IzyePyCCO77P
8E0OgSvRdL8t4b7OEhzFd5h0P7Vtxu0eDDdWrrlnffS8+Q85tHJmS+nnnwVrsLYY5oSxrY8g0WQR
q4oWTTIMQ5+NK3x2f8jVcUm1ihx6VEtTKRl5N+kvbzP6sPqfrCOklli3X2qnivwLQ8p2Ug43u496
ecqXOC91f1mKoXJuRs5TESoeUEEEAjJ+oSWFNgw+MS0oZNekIcSD9cJDeSN0i7/xvnaXRhi38T6h
lovXd0q4jKtS1GfhfaYb9j5BQq2/MbkNfpILNIZMhRKB0Dm4OUXYnQ6IXawR2pSnxZWEYzoPtAhA
4e+ITIPb2Ua1Ft8pGrBT4I0BfnsstSF4CKKqMCSkzI15bdpzVVlsZ47Fcpx00uV/+AxLn3vhCRAD
p9R93luOoPMVkw7BNHa6lrh3dP8q2wVmZoYVYkYXN8P70eb5O9LK9X9f+OMFFMY2XedFhtwWtNMH
TBwWG8B47gXAocVqCndNd6V+fhhsQXyObLt70NTUYFPZAoVWo/OYa7KGWMymhRBvtmYyFMeCn7ie
3h3BHd5ciWLtpQMZOfqlYHDnHEKWYffqIZziQ1FwAlWqZ+sIjbRoIVyqGUSp+jolP2SUKlW6Pcqw
mq9y9lMara7SK9Wt9K3AOHJYkbYiHXRx4VmVDjYK+Uh54EmgMsshVb6B+reMHnwubKyzJBbxFKE7
y1ICW7+KvMgkGY7UXpG5pv/6ht+P7u4L3de7WnFr8bNLDNjka2uzVdrhSOxyhA12iGoComq/tioD
Cgw5cToMIjfFVsDSLzujve9s7zTQ47hHAO8eXaQy9mmpmMnQ7btR5s0xN9tuEI4ei/QVPZKokgbi
+iy91PshGbEhQkmNDmH8yVozx6fVVUOuDrEbSPmgATmAjSAR8Q6j3IfOg50vGq9DZt7zePTcTbxI
WpQliD1W5MRso5IrXVd5nYnBEhWFlhkcJ2QSoC+XPEQRQPxclyeo0JAYDD+dwFef8gdFuj55bSAM
zlFnDC5VuhYhIslLX1i9q2shz+aPUnaMdAy2bvgbKkkZE5WjCUbdcb73jrkEdmSHim2P9F0e13D/
VPgrDBKRUUxOtQ7RGqlpjHRShs9g13IdIfrQbNVLDeKodIh9IZCX6m1r0qa+jXDSo4tKAF9Hbsa+
rZmPQJDNH9Q3udyqrWPk/YZt4J5duSLzodpM4/yly2ulva5u2tayD0sVuboFZblUCiNzFW0sHw+B
qKO22qp15F/kS6P5vCGU+lprbVLffmdXAayejks9Vh6eVF/FrLEkctQVUK4lIBRVbuHI3gSrhNLh
TAprDOKJoCYgolaOh+m2xLKoBUYNKVctIS2yf1aqou9Ca30YXe/FjWU3EyAXvhzLkWMwYeBTAXvD
BzVYVd2xlT7fKfPiNYpIbtIz4rHgIK5/3/OqyqemTiMICRBYfwfuHJPlpYEmSrapbn/q+Vf7xKxo
qw3t2ctGA/QjmWyI9f8CSOpOXEdkf3JgVoRZQhoWsjG4jwvtow17FOoAWJIVGjnZ+APHHybGHSL3
2QSTNp0lRjD6YBjY/NlcOB4XaREaLyzrQfVXSjxFbIEEDJ+ds/tlj5J/OuuaodNqOffwWwZAuk2b
bYp85HTD+pXb6+3zp+SUWND8xsB0nje9PLlJEKxKEJEhwRNA2SG8fcfXcVKUCLJS3yNZsVZj5Eql
4KA1dgy/NLGPZzbEpRPpi3gRbkN5GDuClfUfuV7zYPCpPlgiQ1SF+Q0thrFwu7m4xvMYqqkKqEoL
R+RTH5dKjx/ccHofubNnZ2vOGiqNnkXka9XNZJ7ysX/Mmu+pgWC0FVmlxsA/9lZr/X5MgZRW0a3X
/QbJgYIcZntyEkWg6HhlPxbpuS54GukHQRk2INJNNGNrJdWwbf/ZZQSnp1h4zDGEa0nOtvDxBnFo
Mf+D+p/o09iDFy0O/ubGY8onA0HM28ZDDIYZ9yihWke9b88A7xppWSQTWHeh2nhuEHjnHhQK44aK
PLlybNHqwEcqByNOAch6aWjuRxt4zhUfDvLjjrsVbtc9bDKSo3ZLLJP/5b+obQFfp+dpa5YfjOs5
hnx5QzFmi9eB0YA8dHZ3pmqOo3fMPov9Of157whJzsn/b/ytNOHNuu7n/b5lNCaFqAPk4qCV/9RM
VTwYbJTW+lvgcO4dGQg1gPrL7SVTMRQeOgXq9OWx6iRA7J0swmPMz6JzAKc8NYfZOrdchr4gQVos
p8mtIerDRhqOwxOFn/K5fm7y+NplNlCTMv0Bz88T12mzv0fm2nU7iit3epxGxv1bk5lL7u2Zcp2X
OxcYp4hIlsv7mXbk+gF9mr7KJS/zlIHV+1JTBG3O+hZaTyOe96kj+LQ9af0qGr+Lh4iPIMtojHSI
gN+GegD2QxAla53ypgsyMc/YBm4hefDhMxWE2HSL7AB1ZEOHybINmBYhC9kMKzyPSQo2LJ+uesW5
5lWutticluE6BoyZ/1NHwS2SNS61T1EcmIUVPUdAyE91Dyj1N0MRjCY0aN8SDETH7aunuNdh01Is
hH/2xdePsYYyCI62LC/bzfOMgLAb1pzypziq5oLmg8g249aLcGb9R7LRSdQ8YeS6DNHsU0kg6GJo
r9RcpWtogPTVZxd2U03rYCyf1PnHr35KK1cx/KJDLsP9ktkMsSuSfn/H8bdSoYS6hqEFLOGGtIYI
Fby06T/XaBlrCCdfBvDec9i411az2P9UvboFJzl7i7JJuP0A5jBhMouex9xFQ7FGUalFqnktDcWG
nsG9tYadGkwCEg7/ojFmlVbHkqvth6yuzCz+P6bxkYcpKquLUSdGqmWutqZdwgFbQZ2ZysmHt7Tf
11bva5U4p7A5/9GOxJqrhTrcM+36NUSzR3znRtQF1ws7uGWMI+HmfpSEr5KphdU+QSv+BbwsXXtP
PATsZc7PDeGXMSssB6m9WLkErrXp0CPROnxoKZ/xB4fSRkbNrmrhU52JlfIdfftZ+v4MPKgEhoOE
oyCOOyJBdHw8rx4mW5b/QFt+2z5mBHU8G3+iBodRIpoMQ3+1eNhK9YeVdlzFSOJU/XYOEeS1CCmn
F5ptxMGy+g3X45lQLxLd9aTzaSIl6f9dmIsJEo6EwJ4cgqUG8DKd9NUNvcQScaMtSQ20gVJI2jHe
UW87vvh7GsWIRHBc6JrHZAAbr1uL51N41YGSn5ZXqCWhgKOFOxn+BMIZ3JUm3CyVE3P+16zgrvny
15lyaeYud/xjZ4YsODcShtxrvc5rmXNdxC4EfEGhQWdteCG4Sj6/PQCYeFIw9vQu0lSmbO7Fy5CX
eHpkWRNDZicLSRaXFlY9nbAjT3/9/Os/xGoV3NzN6tLBuym7zjPvNd/FEctnpULmLGIXpjMC/66k
km5bw7ELvA+vVmXtJO8T542RuT28Q8jJo4+ISieYjYQj0gI2s5uoQZLSexazTCjyBGbO++YVzeL4
K5WEXJPXtJKJ/mzez07y23B8zUmCy7d+XRwPLlvuV53dfLsl0iijwOoga1amTkU0iVdcyf/S30jz
8eYOIeSTV8EJMqedjfPI9xD9nj5kq2XNK1ShYNhxUYgAvmkWLsDLRUY9cPKtp0ukptVpMinqp/Qv
fI0mQ1IDfeLb4oFgSU/e53jXXxR0+7gW34UZkZ9LICP5FTzEZ+bf5C2oDxOgqmctpbSSieaefCQW
BzuHXuKrzklm5kWMOG8+XGXHHx/JenZQUmVZuuqt90cNJ5dDTsanAxoht4VwlT6Fcsleh88jgLC2
zeyVod8h+bEUWmDCyDTvbQAfdsLw+zHSSzLtDJfRnVJrUQSoq1p9zheG4wWAXQLPSQ9jPUBpO9Vr
VaKhGHIvszI4DHT/nK4ccDeXCVwpSkvUDd5GfrI7jiIgm1aJRr9BCi+7WTkKDdBqCeZ4JVCDFfm6
XmuiP6P6GLdU8pFGBOdGN0Uz72efH3FCk3mL23270StfaTB2ckY+v9OYyb315BZDRanYKG9q7t2p
DXf2amYLr759cNJnZ2+5ugd30Hrxv+mc30d0XRjaQ052pkjDObKo1mflYYkFYLCJjuPR9Fhkp7ID
ggB7wESCsj7c2c2EGH7ppLwtLgeEGmxnd9OFO6AEOD77wrXfWNGLQm7Ct/fIa6bfQIomN+5zMD60
XkBf+Ge62p92Mv7B+ZJuHSrQhke3876Jr+20+3L39gn+6L1zVjUOp2aDQIvAna9QhuVN4FDj7VvI
CziQM3/5+8zG5WyNzvktdOwxQLUgTdh4z6M2uuS14Xza8x2W8J8KeSvfD/pr6RGH0hnZnd2+QFWa
81ka/F0GrA7TtsiHn3x57/LSAS935MbPV2gE9xV75+gJiH3aRGwLN/UfATKc+QX9rWLDU2NWD9Nk
99M00OmWxcubJhhZnCNLnslD1+xDGK3HoTwTLaTPQ4gsPkwF9h+Z6AH/qOuj1gP3bcoEKXxNyhRV
gsgAtA5W6weg7aI/ipEw3aCvGWr1t7TfpRyj4wy8UbdTkrml4qXEll7gjp3A/z+tSZb31H8QgvBG
zJQWd+og6CIiMnX4yQk9V9Xcic+Ij/yoBi9lQW1EtpoSj8uDFyv1Lr0+TpbBN8zNCBc9vB3QYHEu
1/Eb+zGkMaTfg84d98INaTGVtYHfr/tDnn/BNsxH0BnDxHKJQBcy8v/MaZynX9XKVl/mkuv43NO3
vJOmxGa32kflLlYdGKxFCXCLx1t/068YiNfqFeFBTkEkGNNeoJjq1BcQUaDqAcgma2Mift0uwPvN
oL4iRazIpLke+3qu6otvn6EZcwnzPVnWXHcNB4fEy4rYfeHQnqKM5Z0yvIbJB/HNB7q11Fhcq0G7
j3tmame+T7jRwc1TvxJnOfdcRlh1kkyhWT8yE8cZj0YQlTNy8bIdKTaLjqfyRFkEm6Y5LspfpsHU
56mjbohq1n1pGSKi7lcdRkbkIpCt2XGKqllEEesosiitq1sBdnKMuG89FbB7slfsI1t0a//TmU7B
pfSoEzUsH2ujyNQ0kFRDb4Q/3Rewg+ontxbh73xefD0o/1ZzWmiaw+OF9ySO42AHWRfl1EQVXxOb
gHpUJbU/Q9svy72GVjvSTuFEWGWMQ5E8nIgboM7ouQGNDQexnPWnc0b2ueRozSj7arAUu0l+sbqM
dIpa6rRevoMXdGMN43w1lDnya2iRbYVp5+PHeKLqKPF4UqEVWCPLZzTja+4W1AIItm+D5Uxwe9n4
nag1+SBsyhK7t/Iz/4QRwLtzYhb50tGRcXFtfqDhg2RqYXlW14kstaKZEu8KNc9mIZGPsNTkhPD8
NwY3W204eoCUj5g6DjMGLe1/CFI2jajmL8LsZ9B+rRz4wCudE00DyZcCXZJvckw1SmKJtoNRSmDy
lkirrqjBQvMH04dSC9iHkIQoihTC2f1A29XzCSFUhpfXTa/93I5s/9TltbZ4KN6SsNmKKRKNAKP7
okeMxvFTOAN76mKf/DZRjTb29J+ocBF4wau5sZGy1SzNybfRBNq1pZ0vWRL3nN/ovBX9odxICYd0
g2PiimMFdCU6nRxcNAdOWy7bSVTFgO9g31dhrhi5eW6YX8mJaLIAb0Rki3/b0FBPAziwDqZAcwjv
WoM8W0ULWNNt4bRej7LjF0NzgjuHu1JP+bN6DJQPxvNIN2mChDClqlYLtpjborLbUIMEiaFNNuAg
LLZo7+zFxSJza9ssgNDGZZqHUg4bpViNQcgfhQnSVCdyRjcMoxJl+hIlrHto2spSwxunk5u0BM3m
MKRtMby/5tC+BBrmC81ZXdelV/H7fXu4OHADifuqG9LQAVs9ZXRI50Mi2hR5H5jZgkogw1Jy87RX
uS/ug9XrrrLms9tDhystqinKnf26HCWMfuQtnKzp7dieWYF/ELWeun6K9eGUQCLu/8Lb20lulxV1
YIU/uSRTGS69HTTnv/z6bRahRC7p9517RgnB9R9UDPl9gBdzHSL912YOWMTmk1d5bR2YY6c0tIKM
UEZrIBzp9OhlXf5v3ksrrdvva0f3cTZNjKKAfLbN4AkL9fpona6htQTexlHKersD/ODiehrIoLEU
lGeb6pCFOtBkcnP4jm4O6Qy8jNCbvogiO9EeMXoe2R/ZAzEJEz6gTmcQNLT2cuUql5O5xNr9n0H1
Hjd/Tv17ZO94DgYaW4SMAvVxiXT8QPOvVVqn38X/gPeXOhTeZxWUrNpMeBj+rPGOqugIKItMmSan
jGebUPcvdaw0AtP5jBvz/LDUZgTvMK44xU5JSAgSeWzwDBxW3ab14Csm+AB2xMLncDEzHK143fMv
Wz/4KThZ18ExfViSjfDhdt+ZwzDX4Kgftxl0NaFjGYyWswq/kf1p5moEfxzjVf9yHefRgkMq3BZS
yV2rSTLNam90XSMvdEnNf5aI1JPwjB4Umktpqn3EWYEP6mWIQ5tjACPz3d2cF7/gyd0oxYVtssmx
NmqRf2Ga/0QkSAUdHi5C+/KYXwED8DcPUlVuiH4MbzTZcu/bW0qeCqupBADXYWl5hZosj99qkFLB
9kHTh2d2FCQC3Ge/5QIWu2gd/+tIe327Fw1o+MPObDJHev8nyLvYr68Zzyw8B0LqP08uLyDxvoQd
bnUF/J5EkbzpmZRNG+nlDaOtlNY7Xj2u71WBh/StCDEqM/5qPatDyZ4KIl0t9A/TYiQZdGWPDcOb
fErKbYRZ4zhBxFKTJA4gYwpJW5Yfq+kHpr85HPfRcsHzeAQhhyj5jfyOsfQh92OzZqRHP9vCeCPo
5Tb2cIz7uf0nk3uGgG33GEPdauuqnj2UiFqsgpmyfxylZ8fXomFf5Mrp29Uv4pvbHDJzUB4F2VQ4
SfgUJrh4j35dJoZIr009RBZxF2bXZWH0W06HDVwXjvkDywc1ZhPAKlxdr2bPedMaW7vfFmzXlvHe
KGMIEaH4ty0rrtmaKJ2IAVIlshB+0gS2i4mEHZjXeKflbJIFf1CWo+wEp3SrcXU+6g2ZkKwcBSI+
ChLiL3g2Nr/vY779dkKUXHsaSnXmgoBkJmrvK3jCJSIIHvCjzuQtXy5xwaDMXGzjYeWv4b9VTZk9
HgiRSpDVLLffRshtz+Ea/NirjqlKTznOl+i7fCwXLeZbnDiyMY3OxFDaHkWOeD3Bai9dPBCM0e0v
HVwJwtJZaR8owZ8qC9MpGW20yGzz1dZiV8naGUtz8VYos2kFOKQWqLDRFce0qDf/jWd9mzrg5S4j
PRfPgY4ajRFUZZ+qN7F6mzP08B5U5Y8p9YH/9BSV0TgqVBIvlGGkCd4rdLYzwWo4c5UiQMo9CI9l
P+iWIKbw0NAiyfL7Cy8vpgw9I0WkeZ5Xz8ga8Zt1un18slna0Wlia+zJOs9O1BDfEyjgRXFAVNlN
OWqzoq4E6AWemTZyTwHdyNF/jA5+O3HyBRhRMkJSYatQy0y0lgxjgu4qgsRxRfrePkysFEx+xRqa
fMpkOLIyWq++FS4k5IW1M8clGlRnNglBxHwKJwZ8K9FhkQCkE0umT4zI1lCUo4+OKGz/790vnqvn
dxTQlGF4yL/WH0RgScGsAiaP4LXFkWpRdsUZ5AlV1W0hLB+VqnVwHy+mWe1nB5j6xVwDpC8OW0ro
klGpZy0zzv/+6XdSM5uAOf02E4lgeOQ90sclmKF787HGpBNjJ+jRg1eP6qp/5bRdzsTW23LGwIpJ
R467a4GHM3ArS4dS0aeNuqw3pHMkNJt1o9BMZe1BvmTEmt++zTK7UwOXCsHVG6djwFq6BXu3VfMW
+c0sLr7mNWMq7SYN9yZdNPfItsP6mSQ7fqeuJNAw3bLk/1Sq1DWz9qX3flq3/Q/6al34fV8lTFOa
6VHuW0PowrQPJg9ffPCFcrEjprdZZH4R+nyx4pWorTYwU6I1tHeyCiES74ndI3updXbEf6S18muI
SF4TEiIQ19GWZLJZtEBswx8rSyz68/hy0f2LYdUFnGreBuCdYYwmKtVlEAhUF1oPEcqfNB+gQWzg
w5kHUF430rVlIJnAjOoRUlLkyr0km+g5c5fOt1aHWlQyd+2LDSE9KRf0IO73jQb66VYVUVuzAo/j
rZZxDEdOSpWzDtHm/UftM54VZoOxuHxX3ah6vNK4KFeJfwKAfQiqNEKjcDXLrp+hglsaOuMBOmlU
ynsz+UzEcsT77nLFJAUSXa6ykoJkx5KrGrOzaYWXcK6R0kcJaGXWGETUZdeB8jCVf2XqflzOEtx6
gMWNqv0DEMK+T2ngUA+y1ypPM4MTh/7Nogvukn/iA2V41OEa19cktNfKLa9F6md8JNEFyz9pSvRV
+Z23FjfCCv+0IC9R8CZAGeYolrfhUplnYCU4UPXuYPIHMPs+lltV1vaEiCJo13SEUT/Ih2ydKH8S
llKTSCK9nZUW7VB/niOqbZ1XHguUK/lxALMubGAd3uSV0dm2yhW5nGW75vmLNGrz/sqY9wp9FyBC
h6w6sMGEb3qEXOhvIemJeP/3t4Ezay1xIh6hej++7HiEG5s9FpkRT7t8GHIswph6k/ToX714ejdX
qr0sKy0YGmnu+gvr/lHz8sjJLc6q27iM8cpVT92bfU1f9AtICXwKdB3YjqKaeqJIYAUkPxagam0X
+Ec93fY9JoADRF7WAAO9VAC2FVLGosU6Ce7yBWmM/RErdPdzj71d060R2SPYkpeQQxQKbmUOgnFK
7xiJBgx741aNp+S/3w1Mpd3JUbetM8L51QNE9rnulAGVnXBmeAkk4AjD3S25gAMwbGzsR7cY2DTr
hmyt+eT8cc6i7pSAvJ3ZntHfJHIWQHz2Frmw6rtgGqWaNhdnsinSUCFSS4vbsPzJAYhOcVQ5gD5t
uqHDU/B/Y78lLtHyWAiY9r/wI3Y8DWjMGeQcD0IstALhRWou5y23Dq5YfKukMBhE1h7/55AxcxsS
p3d/SmY64N/+Q6i+OgK5rQuh2ZAJBU9wgY99qwcXtA49+65SAxEHsZUNQcuSdpw9OD7m/EORK2Se
GJuAOeBjrJXE3R+Cwj3oYLzadjX6IXkN+7boqiXg0pN6nKtPvipCacc48Q9JWb9CRItK23gQtuEo
YV4pUXJVcHXNEZoWn0OP2mY489M1GMJBEvPOfNdUY0iTjMSXMbJ9ewWEPEc8OWsAEOpfg/kbw7Yn
fvIAk4aVtEXfJfrje4qy1fHVd6T2CWyFhepG6jU+rEvrnY1XW6XuAV+dUmUUTl73uU67kL0kzRzY
lTq6L/6tzaRfkfnoCGC8WXEdV8Gc8hhoYsJNgnpflcBVnmQpdGT7LKU94yd1B7JUUOkNBrEDk7Ma
S1rW6dhYKitbf7UT8FYzmXmruJtIFBNoclOujx/e5CZUTOzj1ypYmM7fG3on4SPWq4DFqy8VoBHx
3P17Ppjnr5AAzmh+XBYroVoLGfQvZWFcxxJbprS/iu2v7bl5cumsQ+Z+DriJlvbnYFY/3oLpQ7IJ
uH8QQTECnNfDXcBeBaLoiZ2mlna3KQPXjNehuDZfiNkXdO5FxLkS/Irjg0tf2ogkVrnssH4oV4cT
14vadsnagEFBHpfg8I+MtHAYYjBQ3aJPdGZr7js9fFH/Wpz24jELHhJpn2cL0SVnwkVeGxZXA14B
mVzggDAHHXcUxQeyZQQLLyAky+nMgwmyT39vQHs765F4ArfgTDVuKF3Burh8EPh0volijhQc8PzX
EyWF6/dHNsiiNMvbs+OJ1wLvrkDxIx2tMn9j1gs16KXZoEN9mH3IMG6tn9YXv+gbBISDX3bhaFRz
V8ZwvM3N1PLoQGdXmwntD8vnMiqovvp7MDn1JdBcd+/nM8YivWlO/yAB/yE9RPe0+3ma1ACNbHlq
egmtsinJN373q9gYhMT9dBoZrHEDtrlHU64SkB1GXkoVHZfcT+WSdPRsL5dAzuV0vHFCDRhW8EGu
h5LNYnLoZ1NhxbJdwu+35RxDm3QTe//m76gehX2EZgG0HmyCS4AZwjnmVgzyMQm/EOjePfrbr34M
bOYfn155FfXZMZduj2ghBI7+VJORNPnRsEmgWWTzOGk0tFUR6OiDNSFdmWWyprvKrFlhOKIxPeUp
bLhDhjR57yoXgYgZn2zr8leT86Fn5iwR4RwOoo3FpNs/5S2IDuiAWuQwdzMstN5FAKoH+lR7Uyn4
Hy0AnEW5CNRjLc4NvvmDY0xV1+4+6vC279VEn8MIg7yvLgwYNeYAw2zl19XwdvlSXh2xfSAyM6GH
v7vOal23L+bjakzZzWR8xrG37/HjhNicAfFhbBkcfoXrZ5qoewCXrOC0o6YlHlJOu7ypciAhhP90
xYboFKlpF063CEJyPuiWhA65ZJyBV/JIJB7vUgpJIVG7g4hfslDLBJYjflobSAb6PIkjlrnwu7jF
Tvx7259IiRebHkPVlnRdx4l82uCvtaM11vylvD2KtQWJFMo5qAc9wLJ9/gF98DWYRedcvAsttAhA
1rvDh44k/J5doA3YpBXNH1hnRv1SX9limjADUFDx6mBUNHBGkH3oXIQ7ZOsntYL2g9yIq9XEYhFC
xW0aAJXHHbK4yLuGVoJL9KFsVyeT5npTItukrfVsIPK5hKsXrZU8O+WJUkFQQlv57IFUoFbBiSiA
Azz7wKRM8rNtK8gFKEV0BHPOMGlbhM9efSGN/XMDHNAQRVQD/5tmdGQbjAhRnjWW6CtX1UC63pLG
JsLD+yRDxBEngV/ycqth0lL6ipiWH3OHdSwVNOgIu8UKtY/Y44qeH6Mkzy4OjvhQGpMBbV5ib6CW
j+1ekxaNZQ2CjF0yjCrYuyNbFjzNkTcJf7r8FLAhGLBCwslrmqWfuvkfMuwN3Lc47dHiZRut5XZh
WksbQnufoQxO3N0J5xDOPfbRB5GJlq38lFUXu0NWY9Gld+jpfo/Zv02kkDN8iYoGDs/gbtRcQaco
taCPOzpoanWddb3SdZEibvjxZrXmpxePiSq7FeIBYxD5TDDOBmbLipfBZG+hc+pNqhtZsxq8mMwt
jso2MHe9tw2koYchUPZviesfpy8gpbbUFcN2r444EwxnMvSysC0g9/CUbXNSfr6MxwYHMiDZHdZz
TI3HcOANWBRrQO1X2qctSfWt6ZEWUP7kP10BF3MRgXNVvZNn0huksDRbP4FGwvT5ra+qrGWU7HGc
mWmjyhGfOmJLzjkhJ2doSUaFKfXJrmouE9U+fbjQPbkK/UZKN+veuiD12fdaeGedggzXvEnW0MpB
Kr/9xA47Kgb+nZyWDfpEEDFEpMHsnGsZSIHAExjUMiYa/n6E8SslmWigXDFCFpcLAuouU+SrzYLj
sun3QXIIRZGMcMhXkVtQVJzdjkY5mXHZo0ojNe2pk9xgklDTN0tJQu4s+B7Q6s8l/aAQRGygLs7d
agKSX1L63PprP9FEW2c6EHe3JeaRr4lLncIPVQOgALmhf5RbN2CXuT5mzL6dmrGwOd7iO2vjXHSN
JcMOYk3uOWlPVhtc2iyc3FjlzaLz50uAa+Wz0G28k5ptdldr8IL1MA4HcFRnxlvUefzpQ1E4RTI/
tb3UCvJs45R4u1CqyKZnEVGq8AM5NU+soK4ie6A1Od9tzBfrIxlLM3qFaKSRcfZ3fa8XF+CHIe4L
d3fk9z5mxTDp6yKtJf3orv9GWCU4rW3/W/tLJPI68dAoS3jq2eAIRm41tV+sZ4x1/2qz1em9FMI7
Kfg0oF1jrE6jSEBShcwLKLLGEk7OHoQc9txxWkNXnb3tXaIyAIYSFEfL5lXuxwwjbmLivkWKu2CH
uaq5mvSaihCxIavxoX5p7BOp63DOB54o8c3c3vWPBjnvkeD7DtNHKL9nNf1T8t1HK0BWw4dVHtE3
akQp9y5OcyfMt7A8ONXKZns/0zf9m5YKsdtHPmu8BAcIP9JOJMJvIGUM+w7JBPnnXeN749YzTbcN
E12ks8/NpaIAG09Pkz+C/oZztFFTEkHzxWxygkezHxDJiquVvxkEnsPfIThETWinvyr5QUtPEmhk
Ko8DriyB9bTckUmRwzvKb1APCX9A5/Avom38+T6vCAEcbvPvsW0uRBBK7BfsOed31OetWk44If0s
a/SqQrL4hIZ9vYVo8wJQGpdGvWCCV29OUidnxhDAKQwIU+C2fVOImIOp1kQTF+F1/PGeLKiadNVv
3E+Zw88dZPlIKhtQQC0M010mSklSSoNt4b8ILI9uvteBpLyn6pRtHKArqA4XddI+uG+OARt8R8pN
5daI05xfQ+2GiNiSD9w+TJCAYqRxGHGGuG4hp9+te6VaSAgYVhbnYh0UOlSOTI/FXarUbZqd3051
Y5tubRDYjlF/2FLtovjD+GGgvsf1b8WJyiODcYqdfA2iOexLENWeIh0KOEnEOP9tLrEklz2e8hIE
EcaGwpQWiqNlkDI/sRXuBt62Zm2F6N/ES/s98U/qURd2TQ7eAZXu4T+UFuf634XB//9sZMKY1JlV
tN++7i1b7nSIu+9Y4njnGESTiSzsGSN6/Hpvfhv+TpdC3wPOMjdzpCGaWK/6JfT/gcvkE9czKrCb
MQAX04vZtXke9KDdGIGLzOqNnJzVajsYWzEdOU7uZOk+6Jbh6LUPT54PYYJ+wNaruetdOC4oHylL
HvxOhd8HAIGi0Pg4A1fNPqYlzEPW59lIBXUfRpexNqR6iZ5ZQcP6f5cJJC5ykLhqBf6lBeAdnWzw
gefolTkDQ1IE/2RIAewAx3IwMHMxrCaATWGX43ricFJVNEzlLn67I2nnsJlE0D2HLWHJPP2efdTr
LHul/5tMTnaSHNRKrTsZiBDvXrKL54c9HwvtCEfOATuRJD+feU+FLz/upae9AtOa7P0AzdSz6qCR
cEe2gVlZBVFGZDJvf50yXGBJ20TB3lhwutSQ6fTNVYmHPGJtq/St3qCAfm9GEWFY+/j6zq2HueN8
bxFvW++0l6/9d9e61I/3yaRR/HFc4tmB1y89kUFRO5+l4NJAOaRu6HUJ1s6UiLypuTpym9lB1Cyl
W0cWERl32ASQ3QI97Y4jRkELYtgiKK6VqnpGb2x3R9/Qr0oREifSaP1dVUc7y+MwUMwbm4W84SM/
+3wRMEky/dpD0WqS0TSfdSONxv6E4vDbFnWQSjgomQCxM0iTdS9uSjP6is+g+CEu8ARCnCtFrvVi
+xpVjUPCtiJ7Wb37viCLB9wLAG8Bij8ujAe2jnLL2nEAt/h/q4LbdiLS8LkYR8Nafy7cRo6iFGwv
ZKKkrZHQwSKtYSnBo978rLbHBhx0TZmcNhcRW3/iVVGtFICNj0oDFVzFjBPEAHv/iJs9uV35v7vf
SugbwRJp7/1y4eUUe27JorywRa4zrsuFrxl/vuz+lJGfWS2diqNFYBO6ffcGQ/tPRlkzm1OE3WEG
29gb5QH5FUQp/pAzAGLc2T1JZ3CfmUA1giB/rOHb+F+AE0CFBNkLmZgb6eNzcXLhEJFPQFP6Jg70
H9xFYALFfAI9bbKqfIp8G154Pd5D+4W0xBlASEfZRySpjGR03XCCmDckWGIjnYEEC9KXcd3G7GAv
zNtFO/0BgtU7o4H2PlkjizY7A4L8e5la3PzwSJzxsSzyWUzOiabCBbspUENqFimARRD/w54cOy8u
GUZAky/dtqyEljZkjouaZDEvQcE5vMAAqa4cFHTME0TnGj9cckTM+RSL6XtuZ4+/dmEaMNqabACQ
GYUfE2gyouyAArWfQxFGMz3OeeJD3Q3iN5yLG9m2DpiVVGHlFoXrpDkJ0Tw7KQuKb1BRcDTOA4kr
pbMBYOc4NSRtJYVwiN64p3iwEJ2SjDklbyTHX74YKJSS3HIixJBqfGe44wz1XVJmbMHAXWs+Nc7V
Qi4WRvD25qpSU/s498/8LxImY8yaAL/32xlv0S/1XCI3F7LN5p9w93xWUc23/zu+1knRn1JTvtjv
ISDwL4OvoZQzRE3QhMmgJXVtQTpUBXW7QJbeSXeV8oLDSCokFYVkaYyLEG0jZObqmImYOdfR7teN
k5JGbIVOe77yXVA1B8uRtvzSIO5OIUNGW03qk5AOMFFLYkF/DcPW9t0ig2eYFjF6D/Gpjbf6ztch
SWVssYMs0sCpme28nyTvfVDY5zfCU+nX7Z/mfuoI6nUL3M/Dmnd9cKZj9S9tNKM06NHCfgIyMkZ5
xQg4PNZ5PgRSos+rje402kVfwsFQTFx2bpkutp/OwEiq8NYueRJOXJ3kZseVb03FImxew660oePW
24n6ifvLdyPdo6z6gzc/FEwrs/Rp7RJp3OsA77z4qkiGQxg+ZHZKQ3P9PYimcRrUKQEhVTmHzwBn
F+P1yzD/rfAX776qtbee12J9TqY/AKJ1ICWGOM4HcyC6lqhObXhVTtHr/K5yLbTMe8IBNj9qkbXa
59gkjy0+Qqqwb69NzQ4rCf1/3Go/FawV8KQ34tRd4ynEM7MNWEbFutyZJsg9/98xNeoXOgxmOEOJ
J3g+UhOGSWEIAoGWKB10H3oX3vtflnGZNRmqpBHPRPJljIZiPJV17BnL6KYF4Gls1OOmQByjnehJ
a0vpLuEwG5IRvEeYyHk1oFwMBvk5xbTmL4BidVASmYMFltLmWCvKUn+gDqqXOtlRr+R08CNn+2Mz
s7oe8xBiFNewXq+Bru3MQnEiynl1xrq3IRk/3Baa/7YyhzxFxiZGvFJFNOXfpZolzxa7BO/R31Xw
VOw4hZ3T3xwUknpGmV02mIok0OtDKr/WwB3gve1ZyBhUbU5+T4nxtfHIi30vZAggZq0c/MM/OqfC
UURgRCcIdA8etiReINi8uABCpagl+Z2ala0TsIsFQ8DqyiCsvWLaqP53RxRXUfq9hyB61mpty9Zg
yMNpm1fmVD+GnoHqxnEiwOphnqpvQ7XXfKlyIoCn3yLYiYoxfYTi5Jt5ZxYW1vPANHxcDp1x+CbC
JR9xSvN9HvEKLDPn6hYJ1+THO88BuPYiZu6PqCcV3rwsihJX6s4V+CzH8E8fuEBuV7ypHIaiH6Wg
3Vg5vT/r+Nkwq+OhURSCFf9dj5nCr+J3ekKsjrSapsOSeqfNX9b2mAdRGMy+lGRaaXsHQGLvryBg
zKiB6tbc1cMNcc9WFTOQehc98UZvo/io10/3n0eiNXLQMzhJCc5/Az94sTBnENMFpu2TWVMCdvAW
GPZu5rj73gzaoGRGzfvaAUlUaX1idAA5CNaa17ji/iCfrgRpWebrPfMxyNmB+bdsDSG/e0ltJ5aJ
T5YHhyjjreV7NjT6N4EjhPlAzwbZtJEj7Qd+m50YoxqBSsVH4utR5kTw6Lcw2HXA2ObZ7dl4On6A
gxl4hoP0C4v0aCuKUpiO6p1a87rdfhEe0Qbp0o9tTdaFEsyI5zPQXlOEAO00mvK4V1r+9eOZdC1X
h6naxx2+gstTxDT6w1a/0H8dxmPq2JvghyDu2NNpgJ7y/FmHPDyL6EsjU18igtMkAPfZvcbe2qoD
OVNOgHKb7hzm41ERtxKtCopQhIiGiPMOKsmfoknp/2ehMX9bh0MDpj1aEm2fEOD38blj7f/LBorG
OttW22y9QiwHfKpG8FH9WhgvkwTgwGw8fw3n3bcQmQ4bj8vLfLZepRCy3NL6AsOI1v2oBAW3I4m7
0i1dGNaC0my6Uppa536YM3sjbBCENUT0hfeS1dOECURiF82MT9Zq3/wvg2fxiMGEQJZgSGCsYqYk
F5DbS7r6AeirDxAFQegZQr7LwEwiL3CNmIYGBugfUrP2lDl8SuajHeLHxKaLHGf112DwN3uiG3YS
h3VnGXrC4bS2p9yCk1KF2xiDjLebTyM2lww+aLXMQ0cQoCEvKjz694w8cXPLN8ftoRXDDFx5O4E4
vTHVXvUAKCVJW6Qiz0W8V74tOs/u4cOwoug4lmezpLa/jKe4UdZnydhgAkUPtxACrWfk5vfiPlSk
hgvXZuWL2ZVadE2BTvfNdH7fbzgvoRRQig2bxewuVrGpRkg1PQl3lcS+d0brv2kt3rHBtIzEvXVP
+Rwpdq8tfAjKSc+mP8wCF1wnl6iL68sh8TIZs4xEDY2N8s0+UU591hQrub2rdHG+JmbPUx6se539
tpntn+KrBRagnD0OpnvIrIJLGP1EgxhYuqXrapYGkafRHIRoy3ySfuG4eFmS9HpkVrmNCRomfJfk
vsqU+mBw2PeEh24CRdSU+wcK8xQD00n3c3p/f18W4NUHyQAwNgYdVYnjb0/drRjChqRmhBty3GAZ
pB8l+LfVgOZPD0UARYOOh7BhHjqrt2abK3Yvcx3FE5kYFXULDL8npKMHw9MGeKFMgHnfUaE6m+gV
wMY+udUFvkJJD1qwlEHbO8u7Y+otjTTXFNQYK4jXa0hrBqzfxO4VfpnGnrt54+xGKtHWMVEb6Y8t
nFgxh5KPXHFRUX6a+69uwzhKpBF2jCxyukR0K6N502mVU/PD8Lyu8smg8SWNW24FNlcx7Py1KX8e
AcLtfMNGoG1bnjApC8qwDAu4VZ1DoNqD1X3MuxPPmhZK8DXfxbrCZPy8MfjHSr/eiPIIbrN6J5pe
J5M8dtgrIoEt1zXKDIHbIzEfF+tl/WF2ZSEKGv2NlCdUkTgqW0vKqkG5Fx9xC/HSGjeXTv/lN8wc
7JpxccsJmNLAZ0WMZTW/eeLyQLNd9R7ds2gLgagaTjFnFUyuQu43HlRelecU9zmbt9anbpjrAmVn
K9BejA7FZ6VfpUolV2YeA+xoPaW7sE8O34/QaLJf7FVvszHKtOdAe+dqjSj3XwcjODq9pexVDtBP
kGg9Gs1Y+x7zAj0V4qqOhb4OM4o1SsiAOybehqvS6oCUJ7XTMilTS15a4bLYzG2wj/8TkIisHkSj
jCA/Uat+5aJ/Kc8eq+q8atmf0BV+9jEVdCEDIHIYtImudk6fuP+pXWQ3VjlZT4wAXzLPnJkbZTIZ
Ab3gRX/hhqkR4V3iZXyn0xA8Oinc9kmCKbM2i1MGdr6nnIp/q0q+oBXT90hig12XpJMiTh/NezAA
6I2mqPffdJmq9MpoEP33EFk+82GpiftIo/5n8pwTIcRw13TROxxDzAf4y8VkMo4JQxx+cVvdBV0e
jLj2Uh506lA1U5hOuwcHNBvHRqkn0Ok0EhyCi0ao8F+GzgC0MUzQQ9F62dwtUiU0+jYT2G0jwVTH
kJsSjt6PaOXoRpm2JkMyoyRksUPtUB3EMBG44KnRmtrbbWDQ5bM97IqbcXU+RKL8saohZcJBPSJp
MNHJiCnNFMD5oy7wT2Zv/XW5NaZLBjXp23PrP8n6FupKvCDYcPXimbesWR8L8ushtqoM5X0FK8ng
cQOM4VMyWdhZXugBwR7rkd11HxfU2rCiU4czq6x5+mHndYSHZYKhD90+i1THdaJ0qp1UfyGdTLYB
wwf2JUzh5DeDUx2TFiTTqfmqJrN83R1RSAZSRYJTymNZUBv6uz4o+drEGgsbZlMxXr3c1b0D9m9i
IYUvFDX9ZdQdD604hUih8zdWAJ7LUm6bd2UsdQrRTPp52OlZQSaGijiRzqtHgQVs4uetAMou1ou8
LBYOeCrAxQ7gwomDBR763Yl2f0TefyRDKIvq/u0YKMQ3zx+2UxvurFpgYAW7YaWUZ71MpXtaV30c
A2IylqV57GvHrLJAQzVXKEUOL4+2C/mYvKvNdnyIYgndPFuHNGmgPGg6bUXChw3ea7qVmU6LKHmz
OylAh6/WiWqlTIxjDd9CVrpIaLVYNbk98BEha55hWMwIx6Lfo+VBdR6m0X/CA4GWc6Iktc+5HGv7
3UZ8IrXXM28GfzxqVDRMTXXcC+uQiXDdiwH3VAeNbR27hYz0lHZ0uT9ueW86rk/bhmJQWErDdT9h
opQqDFSv9BVb2KmZCx9XsY7QxPpHG5tq4ut9hduj9TwDkXsANHNFZ6F1ngND3I35ihFQYdjnHNvL
Lio7Ma5tsqvMSXA4a0dNu/cmeScZs/9XUVqGsLFpPfGDzcxWUM4NgJ+vWkjtK0/WZnUl3sEaBek6
VcTHoPHMANgEzXiA1HgijwICZfUDkLGmWSeZfyONaUoq6Q4qYulY1AUMDylStpQ3DLDAhUoW1QXg
iV8hdpeLEuQqIwY56j1aU1zwoooLEG5olzU+s1rDTlVkSozNkdbk5dh7czAmzpGBnnw/M6df8Mxe
h1dSAEiCyT8t+ozHNK42zJSgOpgALAVfEvTy9BCVEdZbp4n8RXiLIignEKF+01NXjNFDJ37lDZqj
jyIDfsEoSA2fW0oChcPHMak6EE8ip7uYdphtimlDu78biEDKoPxnzbmrJZ3XrRjhjbvVbLzmeMfv
zzJ0iPY/gChUMpE/d45fGpanOj0cBczYDIwkydhe8aNmjirabNBfg5YhRVdxEHD164rIw30rsDlg
UDjyDX6FuJevmdHPmT+pVAnZOE2scy8llyubKOEmm+wwrHd6Vz2gNtNluZh4iASh0OWUNniX+WBJ
xTr9OvSkdzNZshKR7qAw6vmQkTxB/pp+btwnUs5HhO4aON4NJg+vSmhZr7n1Zbhg2j84sMAx9c0N
vK6CZqW/V+dnjoj6A9UdinAVVR6Q66V9zu066zUHXpGTSKl2e/iqarkge/zRzGbbS+IR8sc5f9nf
8xF+RsOhBwn8IqO8QxFgxzlwsmUUR3MyFKuTDc5gpcsjhSQSWvMtjGGcDNXnWw75JZ4+J6u42l/O
gyoO3kPrtoRC7uyIFUmp4wshO2ASDLdJ+2jaJ1seucaPWlwtciwao8+H/WDDCT07A9XcuKaR3yoY
jYUskuu3jgLBCeQOR2c3NA0kGro9Y59c2jR2DkN7uiDayzXIQFG+r95y8Eo2YouH+2G0wddKPDQP
Q9gPtqeBFeVTZuVLzxP2NjdfEMudoZA+hjfeUKhmBUrEzXMiAxNk7Edha4ifaq95ukl3SGgAWv6Z
eWaw/+MkR8pTQonCZ3DK2pts8qQ3CxwLNHZPvcLA2cbknartZhiVCKwxI2q9upJ6NZATWzhKXA+G
at5VfKKB90jTrTRvaaModZ7ULDHLoxW4GEM4nYpYOEkQizd+aN99ZqfObGJfwpGV9QENjE2+eVmm
x7ddirAJgHdaMg2nMNRsAo7ermpAzwJYvsD4ZTlLlz4DkaDdYXDRPys9021A2XM0hrergdJYddKN
2Evl1JW+tG2tSwYwCVlf6awL5zuqiRdByo1/ZqwYKM9v5RHBUCS4uG312JLixZG6Sy/8HsOaFXxE
u3RIgVbuBo9cNSsXtzdU97463er9RqUkpaJY7vNidRhrS1I2aYjVKJKErxDIwIgpufsIDJPOevcr
/8jh4e8CRCMH7Mx9eHN/1Avi9TPUCc4CHkJ/q4XtysgR16Kj83ll+ZhR4z7A+cGeb5L9JBVRZjqz
W/ulJVjHUU5mtWe1IbGEiV6dZBfEI+4rn8WRUYY44wisvFBGwJ4eJUoeZbobfiYyZTiLKTwIEifu
v5KLel9KLu/xJTvehW4XVGFXpTGfYCAfoNmyIpZ9iHxgPm4edAl9L7K593F79tlt/UOJBvBqyO06
EX/3F9yoElnTXoR4PzglzwJeeQl2PSpjLwFHyrBm5R0HKZHfXIUeCU/wVl6LrGEesiLoEQnRYuC2
h0+R6gcPR1hLhM8FIP0ukKjQM4eKNOfMZ1Ow4MaqbyyKEfg8TQsOqzaP97IkKo2fRtvwn/nBObhs
XK2ujkyEd3DQ0yy/W2uSuSOllVm4vfrzqesa+unVA0mVc++rlFTjhJq5QcEyneWwx5Tw29UbHPDY
zmfG3N0+h1RJUBkqyu2Oj56pyilwoLdYNnLXo5ECBWPWF9fvOF8npkcvhBEbCDPtY+xsMGmPzrK8
TbdZVaMO3lWBN55DmciHLi3igR7uXZyZEVqUI3PZtv8hGbKRjemZDgCObxw/WycfjpxHtK0qTV+w
5yjnaP6apDHoK6rU2+5GG61yYD8xuOq42DEVWo0/aN/b8N28mxJ0ywJI9kiGerXcnti1haX7dt5X
8I2JKsC4eC4QPqypI3wvN+e4wYCUZqDDrtnpWVeERneB+uy5CqlledDCrNU0KlPXgOdZIrymlHHa
XInoOj/4LYgScoY+vyvhh82SPeUO35eNBySdZtPM6RGvdbKc05f3QU7amSGf5z+DYPDI/beBJB+R
yMK05Snp7zEu10T7CbrRjdjByB0I8WlbbJduXidAbhnKnsjhQx1WzApvkEqU1aSN+PIY/qJSwpQZ
9+NupvNVkSATQsd3uhYGj0mwk7xQMuMi7HkcNuuiFPKVZ55vHXnwUanmN2xzF5k2FpDxafKdxIBs
hkG5HhQ+j6q4Qv+KTiCmDCP0xH5zqRYP3Wv/J+DbcaM3n8in1d2NPT8liXpS/xf4iHp+a/G5f48D
GWdSzX31f1o3fjwvPfUZJRnzlIvhiSGe2Dy1r5z1xushnxhTSK8Z6ktxIDb/9OAFvIG2Bsh+2pWf
ZCst9RaKO86pB01EGuznwy6BpNnhCW+KRH7V/HswJdUZyiySNizzxNETrZK87nq2LSuvLMfIPrxG
BE3+szZEMTb6aZuY/eLnueLt34ec+3OexrtKlBIBuy/43eiV6fHV7tef8JOTepfhevNXT+V63inu
KSru7NrMlN/Papy02jxq6ejMlBYKkfuY0Lahlebd7yidwN8SqQpsT6jQLIukEdkOjz2ypfPtwL3y
K5hNBSPxOZDZh0kqPmvi4t3X/5PF9drNzEro84a7p8Xva6fYNyXTjBUVQQfjZHwybfXhwHnEa0OZ
yaXTYaFvbqHz+PK51901tYxG2NE5FaaLUDWKW8+SNX04dIy+Ak+3mLh/1as43A3nKP/tMFuarT+O
pJwfq9BDKIZGtQKwoYliNoRAFbJaCDQcUCFYrjdzImggClLnpUE1CotloW5Ote0XCPLkK1DLSjd+
tuOLHylArmnyNi8njgdcvTZPNuO5tru2B8ws3F7CB34GNz5tbcbXXiN3BwjZamJMC/b+QjFCFgqb
/Y0DcWmj+i69CfcKxPCvyOMEjrO61u8UoFHo+tROZJZd5LDEKRHwdoL2VfZTqQEBNN58tGZunWSh
DoEKHO3+ZyHb/VLWn9Ua4+7+hX9Y7xbkb7ianmwv+Ltx/d9RlMEXeCQu5FZWhloOiUnuVjpDltBd
EIRxkp51jDfPOgqUZbj7d1ij8t6WZNX6CtFccKYmGI83EIt+daDV7D22oWd1tfT+3XeHedJAUgdZ
gadILZtg2hvuTYH5EDhnNsvvZKToit2B54D+HoCmspfZabbPXoq2qDrZ7T52lv4aoo/0SE3tnNxz
FdsxO3YajRxY2cYQ01mTQYc2age0LhvDwyTxeYJLOXJWq2mHqcP0GLv+SGkwZ4BLY9e00tGsEDnz
oXWSnTvm/xUfaMQKhDwxyNb8zbWAMVxdpvE7RtXHNWq+RnYEG7v2NqUMpVKurNarWCWLIQVY9CHd
cHEte35kzZEg/b1+tAy6W20Tebk+7W4UipNJUqjdaFQOlDvQs//k2drGqi2CnhDv408NgbYpehtn
O2VwZqg9yxe8Rl7msTxVJ+G7ktJTtGERuoY5BW+eHSpp6f0IHvjW3lPWx0uxlNXrqmf0Y47yfGOk
sz9YXowZMg7iHMUGxgUtWizcfp5f/CSpDOBr7a4NQXM1bDzNnqOHtGoujrTxZT7b+0JuCymESB1/
2EXzNLVlzX50iIowKdd8OKdcIGwjR3LioYocjhAkjFzpmhsv8d+DIbgp5J9LHsNZeEdeuY40oW8r
bJ1KXQ/9u7FysKxloi5rHcq57EEtEdtztE7FMqqz/TuH2tZSleCCFVnVCEKCSc6gLWslD4Oy86on
PaVWhzSsmMLwb4AwfsrM6iCqezJPid9DNTSIKClN45lvbYooDfUyTTaT8qi5hQmS5cV/v9Gegs72
LecB+y/KMxadxjbbNH6efNbuyVM28WQhVIQ0Lcn1C6SUAP79zLtBdWkEAV19b5HjAxWPkdH93sxH
+RKmxRa7Ku47Wror4C4Xqdwz773IMcMOFwK38QtFtDaRgUsauid9nv9UrGhmO9Zskks29eqe2s9v
cYt2HITpBAPB13E3FICttuZHBywy6KczCcTutSKl2/qWu+LHVD1m9jTz6kBcX2VJ7vMdMol2y5Bo
yOpzmg04vPHEwMaB1yFISwjfJ5+OTPr+6QpLgYz9ycrZwgKhmMhVJtECeRg2V7tGDLbePdUlWFdb
gj4r069f8QP659zGENH7sML5znFAqct0+5ZLAboEOjLz+5kAjyCAgc1Jc/mPhUlexa6LZxZKa2yK
87BAE7YIsL41ENEVumRM3V2UXj/Tw+lTUjL031hF4zUQcb0HRzVYEJujEGav+8XD7B/WdZHdca/L
3vAb9nwTC9qsBBCCy4a7R6wPWug84pg4p/CvA2UFQ0ArR5EdH31/yH2dCE6nmtPH82+Ejp/e90C/
TR7aN3C6ErAidVkllcMjOdZEaBUK1xBJcI/k0lXD29QFJHDQH4Bv29JM7edBHzPUPNfsVmGsMhti
wvgdyCegsk+52o3MT8AnP++Ns/L9OcYfuiYaQ8tbT3reTqO+LEWRCmpo1NSKkNykUBFOm3EYI3Iv
6Uowme68Gt0DxhNd8yQLPJF18fLNLY8WtDCfsPXb6zpKL+49+724T2RqyrB1pwjkTNNrrbO3JMqv
Pe0iGsLbgR/Qmn+xuzRHc5VPZisRdEKg7xnv7eIGFoahqOVwheipjiGb0DCjopY5q84nwvqwb4GO
cpWpnsuKz0STuVHvXu6cSbb70nPUqKeSuDwpGZA24mOlVMUWpY3JK2zSowrlayTgvFHMHlN7MltH
bDx0HFBORXhBritl52O5YQNgC0+ed6L+COm7ZeRfmQ/pgkHNXr3FjTF2WP55Z8Jetu1ACUXqVQru
KcakQPbt1RyM7MgHs0SvcbxlbeKKCrHMPJaWuP/MD4LYeuy4fzM8zy0v780RR+0yuLMUrr5Q74Fq
PjR82CiLJS/cR+Sg5xto5DS+O7gVj/Zz2olFSGiuuTRbeYu7WN+sUGen2s5VVvvPaYwTDbWN/Lny
W56NnANlwgd2M7qfK8l8Ul7VdsN2+rJkq64v4yqhGSGyY2wfdFnbJQLKgS1xTY5lD9AdJTj/oTMK
l8A/RBijNlRWi7LYmu261c+4pv6PVvwOW0HlCucUqPBoG066FENRQheC9JD023wnvhf0vCwA8kuK
80xAPWmhbZraDx9OD08ZImEWN5FLQzZ4HGz5CYg7Xai/9SeqbhGknSvlQRv3KnBkCdPChAfUZDjl
T2ptcuEhWYDK6GxmUKI3L5ensSxWuRCCOPvHXf2VopR3BooGhQ27UZR/K/6k1JEcljrXDPT3EC90
ECBDU6j5blq8n8c9LnGe+NMtcULMuT7RUTdntBkGU1zThvIlaMQvEvI+b3jcTTi3xAs+/aQ70t6W
fOmiT3XXHLV7GUedziqdeJQ9Xqjz8DTa/R09xU0PahL6OWFofMcEVuIEDjfPqykTqwBL4KbOKAdJ
gLvZ8LNy/hWBglz+rj4jbrkUVn2S9QlF3SrEXLNmVE/QnE2xgLG/Fgzq1MLlko2BZZWljDYELPO8
NHwkKYoRLik3MOXZ9ph2l4vcUjzbwlR+WgN9DLP3mZifHOkupjWGrY+ieMoopsBJvMyGSYHTWPtn
YrLEZxmaRjK4gT6eWCc2koX4rEuYFAFYUT3avNEhj+e8IDpCkmoqwLLqdMPDH3wplTJcaxUWOU8n
53w0Pn9xcE0jGOKJZWz2LjHlGta99qomlpD4yd6XLB0xGZtroiOeRu2as8386GuJpKD7UcOMeDHN
n7I2345u7G9UFwYvfR5EJEiEh5mGnG+L2AVgQ/8yRYphwoxRIYOpeZaZiMUzOMgi5O/xXFOycI3x
bHVZrNV1PU74xMB/8XXqd7Ws/vqYxgbuN939anb8FK3ofASE/IhZfPpYxJzlS0QENEgXd9/OreGq
IkByw/JIxiLfLZ3ifuC150w+L6OL3Try3q8jQNU9PQzJbfrDmRU/76AUw5cfkyfiTLNpAReIQCVE
EGhay7x+DZF9ZsEaJuN834fBHS+2IE9ND2J0Jau69IDxsPsgk66MnkTRbSTcLv4dhfPKA+EERy3i
nJ3EJV/19ZR8ULmROEWBhwaydVqZ2Dn/2VadPc6n2ElEeOe3039AcJfRTHLPmhicCxbRsBnsd6qi
+ie3WSgWLB0KrlvoFy8P/n6U0lNGuygVUBFtmbimbyxps/FuCv61DpqnPE6k2ab6fNXq6oEgQJf1
7JkQpoNGdcU6nvuVkznX14JVe1t2KTuIXxEnzwpPQ5mU4mYb2rJR/ZVN4A74NvaFjEd65BxbiQK0
nDkFS0jgo68sFDZ6EGoaktm/jElMpMa5xelqQsVqW/7I1hb9AM/LFUpzT5H9aSwxAeA6yEUSp9Yz
ETDu/Oj1hOr/BFkjb6a98mrovC+9ls/hBTvvULE9HJA1GmZRINc8ozpeMkBvPbhqBjg5CwnC8Vd4
4p6n7/L+sR/Ud7X5NOfOIZQisuZdnY6N7GuZMoP5SLzXKIGwBlmPjXj8o028W63IMV9HDcxy2j0H
3lDel6EbzhHQCRI5aqc3pbHQxG6PsHRYyAbGIuanxmPIWd+Jo3m5E3S5akyZIPddLXP5AcKsG5cx
KN9FGaL4ivryCRxHU+NUZn1VHjbRdm0pvPsOATQBtv88rqdffOXiDJ/5SAXoXpTBhhT8nMgiN43t
ix6wkobaM4+iAtu1XFxWKztrRiLipnLTx8mj6dIppQAPiCbtPF6WYrKSDpfbj/5Uc0weT9yBMciO
x02vuc4QCdxp7tTmzwFfKG6cTrCtLOewl5NmFWv4osTehKo055Dl9YBrE0E2NurYdBGM6e6CsdCa
dtLPkfJ64fj2tG6DEqXVTrhYRDjz9MuvR89C+FsYZDI4liD0gbPUkTBCELH4+AfjEkq0sbmuCF8M
iVCH/cbi6I6F6os1L1jvtQExPrhIcDgIZK90Dw3YqdNcoU+KxvjchVL2bFg6Yi6bKyiSVxJwKtaJ
BNARB36YAjVSK4o4KaLuvnUnjdxcB6UjCCcuUiIgHT4amPYWuknpOnX9iu9qz1MxvuYNpOxrkhju
e1YepkMZm4N0cZJkwipNY29JoEUbrwPViFHXm1BAiELPeQzIulRS6nF0j9/5m612EfxNmz9C1uJ8
Kshp1S4T+WK2PwUmtZdPKLF+vpkmjFOTsAN8r62oT7gdhf6MsjERn/ViF1tETSSFgtMKEVV9Krn5
+60cWhihdHMUG5kjyE0pJlAVWFC8EcZGbzDvMJdKJkY1lKoV+NN24DBNCQ0WSgfgv/xIQG/l463A
N7aEhZIRaNPz+duXCfuTwl+/vj4qNBGfJQr/htoh1qyE7xORTqyTVz7/lgCyuNP3os+e2giH+DKr
859HAgjggI1Z4VQOtry0DEmktv+VYComHAOsMMrtBzmSPPYtzD5O5uTpfN7tgWWs+rbV/dZ280/M
I/5xA0bGKWS8ndgwDhDKrFwRzz6/tdOjdLm3f4/gtkQXEmYlVvmiBkHgj+3uxbZCHwyxMsMCBN3C
AfTlmSr6LeQDrYtqcijjxOOtUqSFRs/DLY8bvClQPy4q0UOF46B0Jn4iuIt0VKqq65/JThGzxs+p
6GOw3Iyt2/yGFoPneHP8w/TF7z/v05v+ebHUbj8RWK9FTGQzzA3h8+vm9N9rEASFj3t0zE0e6WGR
mp6zB/AD4CqvR8axAOFUmNsjuyOfExBMwtHOTRYJtiEqbA/78i3WPjtYqhhL8DR8zNSRuTPZ6hAO
mjS6d/ka+1CTI7sK5FIp+iwGqEkwOjwfahVLIHlcvzvUNVmxwos3U2BMsMijd6wcIBqzZcmHqJxY
WzjFdR9W85K2Tv7JdkYreZ9Yam8jRZANGx4NkllFZ5VWVZmpfjayK8E5g2lSmgEtF8zLK8lIpYEq
6OvwgvorB3zQnOzu79b0V3fPpX7g8GjS5RwTFAFeKmmRgFsEYjHksjUex9PAgx/ZJ3/hJ0oGBIXB
TKb/DaawRbw/wUtDt0YqfEAu9y2t1Vz4krpZVXXTBjSz6CU3kTXAzIYTXHVK+nHVPGQh1nCV7xn1
Rp8TDPqGpm/BKTptl4gphFs7kVJXAJLBNLemFGo8WS4iFPMHeauDhloCqXSXqbCsuGa3VW/15GWs
mx9ZUn97uBK8Q6bfKrLG0GpnVEcHbqjKYgTLdj56Gg3mAeObJBqjGvYlDYJ78bMAu/XIZX0zzDPd
qOxIHr9LubpUFSTJprjjyCWlm1QEr4chSU6xjJlNujtzgmr8Yqp0QEHDGHZyZsoRZ1IZd37fPlAc
ayGA4/hAByL6D+xAptPsVcHaTeXl6AqGIOWqO1OlPJSrEgyJGnOdnIUlJMTTXWmpndANwywK8QSl
nrKoBfP1b4aPOHtRskOZqGYQafwRtBUU6j4Go3dutYy74FoB6mHLTn4c4y+yqvAv/bxtBQZkIIZO
h1+nWF7pf85XgMZhHY0gSxyUa0jhc9ExMz60dHyN0nOP+Cew6kMbdGv81ycVJSWcsJ0LSTprt0fN
Xsw0SJiBIM74Iyp+4ct9u0Glzysa/WtRNfDEhA5ckAhLDpVC4ZkaMsIANtsWSO53ZqXDVyQnjUH7
TZ4/MUjP/Ejg2HZcfwtLPHrziGOU5K0pOgArcOG4+i6Q9/m6j5UgNctElQtuV8/hS2R2ZgIQZ9W8
KLPFB3KdsDgjEqrIX/fTgtDRY+LbG0p9DXkPUFtC3BgNm742Bbft7fSIvmEj+V8ihc9k7cNvql9v
pEmpvMTpN2GTX//bp7lAmMne4eQxiCt8Y1A5AMxWBdisbLzjHI8rW9fpt0NxAtjjlA6FbknoGCYi
8HdVmCwZQLz8ozJi/mAa/0Ld0G5lqCKSCQ6gt4owl1tV9OvG1yDC7/plEmyWrlZKTimVFanD3mFC
MHuegbSY3erMI0NySFT2tr3YVZfniBeAZXMbQTpHdjnIzxiKNyyLG4ZvC6njJ1l56KbmU68EjGKp
HcuESkmZjN4S12IuateQ1pkTy5Tz168tXQzwF8KTEz4IKlRzuEIcKgzd0B4C118fy28zl58NERpP
HLaC6xoORqwko878fxVAiS9m+UvA3xsTNlu3HZjdF2u6KeGHW/8WyqIvECPMJOie5xxmlZqB9+3/
vj/3O77mOYvZE1xOn8eFvEbzcYLHSHbWMkdNycqOPJp2iDDKTd5AP0OYEYmuqIupjjB7sS4IJeoI
Jh6zhRQTVxU6cZ33KN4RrEhPu8oVec33UFKdPYy2MNGgDFhERli26rd/54D2QQsUY1A7aCrU52Sp
GmtZ4RTjTjlYa9nWAsnRAu/xbrg2zxup11BShsg4P+G3q74xGB8evLGx1YJNjBTqq3iF/kfoGUZJ
9ZAsLrbNh7sJjLkrbJpoDGP8L/XVz3GSnq4AmsaW77LnisFOKMCKIQ5fVS0wEbtWy5K9Cs4RS5+s
U95WF/WipNP/EHOXCdp8X2/ZBCla6HSjO9dUDEciwwMrVZtm72JrHWTs8m4BaFcx0Fjv11rxxtjg
mWajJILnvlR7AjlqC0GMSGpFVjgfWVTUk1FDbs/CMym8CTPMEEcU+6DZ5cTeTCeP4P9DyHz/DwT/
fDZMEeO3P13HVCqWBfn5lyK0wMv8usWc0OEXQ8RnkolI8YPDK5d8oyu8A25SRabSInTyfpckMDPH
jLvqShuNP38ooEX/AyM6OwJlzWPKa7yDmKhDYE5dt5SeXIg3u38NdyE213MlbtMg6LG9XrLkBoUA
vk1MPT7fTS/WmgHUvO9/8sIO8JmemC/OSQqzkLLksZWHCO4dNMwqJqw3R7zLRcace1yx3zU+B1/+
E758H4aA134tuy1n+9cO7nsWBLNpmMRQleCq8JVbZNtB4GPY9OYU8XT1oE5A0CfjyKXAjHlcYn3E
848zB236Le6/JQDkly/63GIbip2FYatMXCSUPpgyLOne8lMNKxQorE+unNqxu4lrszLuDT4wD6tP
zamkzkhWe0B7nRrIsWKl8NWsCb/58KQa3QXRRsY10nEebOzdRNlae0wqQ+00EN7tJkzKi04u5qk2
hV+ukIx1OU4x3UeXsYRGEWB7N5CpXbP8XM5UtmH6iC7lX1DTYdXETyhh/gCrAInswiV4Mu4NwwvU
nSo7pS2BBVsm/Bac5OP4wI3A0nv9PsHgpKoMcqO3nNcyRfEusg4XQm/qffU/ICtGwoDKXtxu/951
Jscolv2B2BkJzmMs8WgQxBHKI+vjrzNQEQDfEQNc5M9Sci5XdtKX9ACdnC6g269TnFFJourTX+cR
xbPkCHEBOL3fZXzFBL3mT0ApvuFKothxjhf2jVkTDcz54KvD6rCiKUBQDislYB6RXTiaIIqhWrMI
7nK0VzRbxfWCFwx5dSFNaWaVnqiNfoP8FL6io3C+gr1sDogQCdwjT32xldTu8uMBCzplR/py676G
JLizfNFb0SQu4E5VWB58fBYobc/h9d+lyuT0CrFWXzHo3tDlx7TX+oLS7QFhfSHpWgqfsn1s7Zmv
2dfMCLn2Kag95joxOH7K20vZS6fkYCzaVoKxazxxPxQo21QxoTQd0k/LPNvSmMJ8o3CgJAaQxZiS
U72X5pbrYcogQxxy8JWGMfqgWPsoJONte0aNPJNxn9OXn8mdo7d8OI/uCbjWabOdNWwTU1MrUeCZ
Humn4ACZIhxkEKgmbwKxZWiwrPzyfBZlTxA5bDUqJ8Ys4VEpvpEjvMUsW3V4DO+eQhfH4FttkTpX
FmBSmGtIGtN5SmX+NRdyDxX4GrkG7RfXWmt4bDOzJo69kwBKZD8kH7+hznn72uMktePw0Rprs3p9
JWk006VmF+JiV5xEl8dTwCm5tQldY89Bikv8Fan+ryj6HhQh1482pRyE0BfO4fwHRD+XdmkwOmVx
3UAgqc2DD/sL6JkH9+gbo1ZvaBwzJW0r5CloQcdwasReh4q+WmgzvKXrTQ0I8GCc+XY7CjddgAGc
w7uLfZZItPguonKI8z48WT8i0J5p3H5OLLfuVZz1pn0Hg8zDLDyC/eBg3G/g8kQ6vjLzAnyyl7aI
lFuxd+Br3amMTtAktFQNQeMa/iWLlKrbmziqUsTw/clrGrg5lR5DpmjkjtDCsnUadbYenbkbAAE8
DQSmwmBoMblxCcnvVIa5Qq4ktSgsGdNtf7kbi05ZiCCcyoO0G7FB1SDrndbyq6T3cpXYNkAyO9oV
uQRCYtYmDMwpQXsOwf56h6hyR+KWqWLIK3svW0O6TG/Iqvmt/qa6xgM0Fl76IkOswExkqvgjFpFo
72vu5R3F7DoG1+5L8hQYMgWBlHyLZj5QLiBngvpMHjmnk4YVLpOg12ciWMVNcX7UhWOl2igWUkFk
VHJq6pQLKgRGeszjsjjPo9CkFz5uvZkEw0a5BvhR/z42WR67lV5HsQ0r4MVWkzkg2NfXqiNUi0nF
QHEkWnFkoG8p5UtgBNZ3tRpdA45yulVaxPAIn42kYu00rOHtdZqlwYQVNsi43cA7GjfP4MiyQxzd
Gas12w9gFPro9msg2prc98VapAeabYs9caIm24FEVi2YvCys94om187USc+mLzDBzOZ1b/MizWWD
0QVceGHDMZLgEih8939PU2MdMJqo5YtVvkiSOeHnkLc0g0OXkDOo11kWkaa9o88NrExRZkW6rWxf
fV89SGHhVt74VNwxB0N7e9W/4K6YPI1xUWqnqm3Ky8u/980BL04+9p7QgG4OJGn58PPuwWP2nUTZ
zImKgp2RipCHj1hwYHuMdNH/NgGF5xVqkXp9LysI8UCNPD8g8aAu5/C056850OpcSJ+YUAb2p07n
roPqRWDbX9pkmuODDCpPdCY/uQBbx2iT4L9qRoQLi/BAFC2yZDc6kIOuWItCyaoFGQYA9psvdxG4
DUthirSz8bAsgCQ971IImZyhbMS0Y+53JOeG8TQXIVUOhN++mFBUjt5k8z3AhNAy1JjhYpFklcxp
/bjKwdf7FC/10RCDFhqr6DeSnw3glglJb2q57pyg1Z+9IgE5eEOLrq8UUKXPnLtkKAwoYXaDzYOZ
OC5S4V6BH0D1oqAPyH8X5DekJZTUluxG1EydRPPPKLMPinXfTlnag+dXxaOyVYKQMXRNV2UbwR5o
f0tzO11L9oq0qpLmH+6STuMU4aI4qms9+PKocd3cEPl0LMtFdGV2ErmGwKO+QeGeo4ThCzImqUzN
VRHTAsU2mZ5hwJ8Arf7bwjJfBZwc7dFyiH7KIKjsQYaKeWHBO48jf63HdSK4sr1sGndAgDOC265v
1OFdlgE0E8f7jZkffLRWEDyEpMUmhwH4qW4HJKQR/9dru44zEgoQHNZZ0Z8i6SfXIjCzuHkFPEsZ
QqmqRk8q803IZKSG9Bb1G1vbwhMtnL83wi+lQE9j/DS9c+SPSaSY7tNWIr69z0+W8iEBgEKjyLhy
tVQVp/7ksBub+DwVlphTmgHN1WTngPRv5BNrhEzRG5JoUYloQQ82WGCR7VhRRXHydCuzBbxaDjbK
FBlXuR98RRWgmv1Mb61Nlup+l4fsjBwK4SznZ4XViW+2SsaYwDZ8EzMQnEDeIMWES8CvtHU7j/4T
QtY/TIklZ74iXh3JH+J3LxvnzkDrZM72zPxJiky8/+YyoEUX45rrS9XvwI125wP5knR8crzjbePT
umGVLJDM55/LCF+Vx4QWqbYGzwTe/UBVcGDo3WHdt+i/sH3leSfZNBucqXHMoTygDfmJebRMphur
02dD8e6wIAYvOBEiJRfA9KM9uoPmQWVzJ5b83xUJKly9B0c9V7zilTcFqp9isXDtAYnwZlaaevPy
fXzEv6gerDibznphUA4xZeQArP/w20HB6A8o7rTjIMn05kBz5MRD/hNoUO2rTslyn2W+rQ+0ODzR
DRG1F1j7SddtEan5gqQFcCGsXYC3LoZtwnbsIR+rrX5u4q3fPKB7lGj7cJ/eakomgz9bmbsaqdBA
5nWnsC8J9vBt3zXecg4657BAZbLTlXa/JQgHsx30NTFXHVa4MVpCGayZq2q1wibtnmQZsJEN8Rbc
7HD6lBjI+u1SgG1NQYY6hjEAdKzRqydOPN3rqrLSmabwLtQSiQIUd6fj+jp9cvP5a0QhVWS04fCt
8Lqb8k0Ik16e5LOY5RSILHPCDU89+bi4QQ5m2cwxazI+EjfHYvQW7IObbdebmAYJf/Id1IJui8v8
QDBENyVFou4T+vewfM5MpDPLKLLOLPRaYMN0d0Y/X3yF7hqLe/XmKB5YNVUa8UZBTtomLrvLKdMZ
Xol9n2vRx3jcGts6xR6ZBXjLD5He0ND3xwMAvLjIZbQ6Or0w8FmVZfyOztCpMMTeYtVtQOR4OX6c
iZ0dJ/D65AZ4jEqoou1Nbd4XHNxItugTNn74trGuHqBGTfmkFNCkCo9kgs8xkKwzzBouq5XVG0sP
GZJ8t7iw0uKLm6FU42N+YoAgjci+tkyV31Ony+xE/ABe9cs+qC6JXrXe86G0yRgb0AAyIuF2qpbF
d7Rm/XP6/WvkoFAoDvEG9+QAeIhfQAgPJZMrOhDjPQj6ZylcCyBkNSUKBAusenEprwOiPDQ4ZXtg
vL1XGvzNICp3WZ6d0pw5k29JYhg6E1RRKderbU1S+1k2B1bsEN2tMKEtSLsFUWx/21pq4MvX1ROW
dhloKpOqdaUudKyqxbO4uPXxPfB674ttcfDAhnEU2ADnqXuu6QO4QHbX6bqYInBFJbcE6nFdCCcN
MHmCFjgE28+EackCsbTlFB6CpsW1zMwgb8rZJjX4INU9nNeVZxxOslsgWFG6SAYrhRy29mPXVpFR
BtohFzj4KCAVjIddY42xJVBteRbvSYsEGliPm/4AzHJ+alzG3XnozoV12Qa9KgnLfA1fEotgHvQB
eGtMYyWB4D5cVSYzipBd1laa178oSqU5bi7xeOIuVofy/a3TEPdYus1tEj47hSXXE1RaQeV4yxs+
ilv6hq1G/gpAuPLAHCXL+SuxsxQZNzG4AvsJJ0AwjcDBm3hEFrELytVCdsbvpHTKf84jlfn2kh5z
p55JMDZPvW+A+hQ5AkTAI0u+3N1fLBil4AuPx2nbAexs5FdUWktWjVHi0O0EAsrU361W/vc3kLXU
lLdl56baKU3SORQrFR3Ym9/a85Uhz6Y02Bjdzdsz+cHUQnGIahkKil1BFb7n60/j8vKsH9mbHu0s
3i6Szgh6RG8XSVAVNeqYd5sw9TT4b52OQ1QE+4lCc1kPvE/ndmby2mb5nKwmt0X80Ww1ENkeLqaK
fqn7MxYmLqfnDQjN5/8YCqf0gnkj399AY8EaYi14XPltRKQUM0H7xFxZCqE+LPS2RC8bDShq478Q
QqOSJul7sBvPpd0pGTY1JUPK7kY/x1E66nur8K3aWu+eoVSk3VNK8DDQSd0d1s8nWkrpRjd2kNdx
lsxs7AuALz3lKUOoBy754HoCWNHkCka01P4yK062KImnGczwoE5s8gKlqm3V0FY1FBiBvIdQRyNt
/1URhH0zXhcIAgxpw40kBQKR+kpaHNsQJznbSdjWz1eAbHt/F4HKjffSKkqQd7kn2tE29QSLzzf/
M6WLuPzbYuGMtBpKfZi+1OYrxC+0tz2TXfL8c1JIquSIF/iLDqPB5aulB1uvJ8T15JQVLLS6VafH
ATKJZd6gg3aFhESvJZYtCrjJU0YVqJ12IAD0peRxWxeRb+PDOnlSaepQ1kQCxN8J6QDQmm35yPge
4IgoVlIJE62lGGBejTqvWg5gLO0MnOV8O7d25uWqg5qOMqBfQIKV0ngwGlsFbe3bZMh0aJs6YL1Y
oBB4vWy9Y4P/ijtQyhE8zZy41aCO70d7R5Rbzv4FJMEgn3Q/7f+TPy3Rx73Jgnbj8moWR3I+UUMj
C1m2U1rCKTlAgzD9ctudgRwMehIva2c4hNrY8GujiBibScYPdIylXB8pPivEhVqD2O50oqZRP2G+
KOCAXkKRHgX0hDnVwj1nWWc3+LoNHpVNa36E3sDRHZbHhhh1vuMJUTfCGeKnSJnYCB+cm5KyuXcT
exHyVRviIYO2UJxy+VTqDjzzwwnoFvYyXPRQL633dZ1Ok6Mn7/CZruxJJ/r6QDxIW06DSDaf0SKI
SWwdFy0e+NGRsQGaEeue4nssqC+eW4BPbRWQQdJ6pd8xinvR7SuXz3JjltAFKFNL2X4EdLQiBA3s
EyczatN8IajNB4iqfxZBKCL4FO9lNFqEfZBW4QGIPdF/6UJKNIRA8y0FGFZGTozFnWaV46qCG4l3
vfb3Ba2uamGuQysEuKOpZhyXjJ139LV/r19c3g8VpKM+YDJjd8LuuCW18mmWw8v/hAvmbLdjXNkG
N2RqRo2htS5N8oqIIjPW5OW/L3nBkVtAd1fr4HelcHrPBlqdnwMLGbl6kFpW0d1noqy1J/GJq8TH
5HdhmQFFbRap5HKBayss8VlpU3LfBeN9QhlZmbjYF6BpbhI6o73SnlZxcZGjueGEjzJP258xZyzf
Df1VcbfzBgjTUay4rRAwcSdhSFyJ4s14YVSD6kKICVGC74ZC+ZgfqA2ovGimeb9H+yPJRblTjFV2
lp7PV7jgM71prQJc7pVff38oZT2ql07YiUEMDVZ98AcikvtXw959Z2FlSehln5KhJFk9GpFAzkLY
iS6TwP39BNCeKl6dOnyq7PxLu0aAdYn8rrtq/CJ1rXU6VcgI3nEaCwgwWb/aMNzTCmszy0X9Lqgq
cg3PCcC9aAEgqVISMhOPw8+Wr7Q/MdsHRh+WIaorDZccpxUfUFaZE8y9eRitVfS92pIJZE8/SBXg
U4aR8oVz5Ok6uMzB55U778B9O4UzGTwhqhOnVzf+yjHH3Nvcqf4to0OI5ZInJDVPxwuLiDK+JHIM
b8u5BqDhIrW6E0fYh7sGBH2+8/mbj1ZM6tZ+BlVyS6jZLpSgi5xdAbk+ISv3jXWCfATSsns0IMPI
aVDxx1RSBqCYbU6vCV97HBM6hVQyIaF0oZvcAVNiC/RUpTfGeEkjor4aS87yFT34WZDgCjDrQyxr
cBcetyWH4ifLbxg+CyphAcgkmC9Tj8p38E7qHs08JElkx67karJ4EZc7K9g/tmiM41cCRXCDu9UK
gpzk5V38yZNsg8lXGP0GZsDX/DGVqe+ED8bBfrMmy35XlfIoJM7ZyLQKXIg0/j26vn0mQpSGQ4Xt
GcMs6L4z9JMF++eXyk0WMNu37BpEbDqlX4jYit1vu0k5itIRyMYhYxMeQNedsYelhr/2jF0dCzWH
bzxEf+H7+mEqd0XE6jTXGdCq6RiT06V9Pe5AH+Oz5+QDroBgR1DtdtuFY0FNK2RTfZPbqH/G2XZc
TUcp6yNwoJzlcMmkMX1TY7/ddYfIuahWRooiN205nd9z46v11IYLZW0UWwnds116zcQvA1T/tJ2D
JLGrtnuYEU33taYHDfBHMMu4uNnZrgcRveRajZtNVcHWgmUf3C/weB8T9Ui7cgf3h6uSVYoUbp8A
fgge+UXmCYN1zfVwQRLo0yjHhaUJAisHsnIUTfKbi8FJiFoRhv5K8LKfhJzabxc5vqjKBfxCTcMW
k/yXC64yxLmh2tQEBBA7e5h4ODBgAJqg6uaTX11vKxGiigKQvszM7CJBkxqjcMDRB9sHY8Nx4Acw
k2MaFkA6HwLE4ixxSDj20njNYLYgXPldG5TYqg8ARbRqzJRIJT47wegWb+zRTGR7Sb7Byv+VS0V/
G3+yyWc/0lggEFW/wlau3rTCumXRN3KQ9lgT4ntdXgXR/P+wHoRaoytnWcGW4j5fE5e9BgmOGaMD
9wwadwRDMm7tQ8B4qi4CFQiCciXNWxSppDsi8DfPCcQo0E3qS1PQRiQecpjHHYpseXP+vIDfRu4L
66K3rMXc7LoLF0g7vDxXVSwuWedlqZKR6MlllRzqEHuwRdrakrmViboECd86oHAabqqPjm8+zPPB
5FdiljXvOR4+vPnEPy+1SffeAonAsuEa+UFpkL8ZVAPoeiWq0zDI3O8OxS69WdW3rYDtS5KQh3hW
Tge75UXB0oXRmk1+yEnmMI72QeIeRrspWWF702V/hcGNt5fGM/Ru6WwfpiZHTWV9ttnv56qY5AkB
Zu90cW+uWFpq3QjqaRncECVc+c3SulE8FXLXhmivDoOHQLRSXgbO2jdQ9tNPhU9Ol1KKodvk+lod
oB3bImKX2ulZxJg3DtV90UkcGoia4w3EDceNqSdYQojqJiazb/snjb96RTBjgaVV7VNQZTjd9f9z
j+qOED4kBDlWQyfNtEEGGKVORNMfiktHQTpKeqoFZ2UNxO8kvPBZBmQiqDjeqk+4z6huOZKukcVb
EHbJWsmijcpQZ0FgTkR884cozZhlbo2TXxh0MYLrw+nrx+OviPIjVP3YhkWOHhnDWRBDT6Ve166R
+VM4fUoLw6jC1CcM9XR1DH+guL5jZqq9gkfNoIgFOO07m8JNReV28S025AzjP1vo8y61T1YU11KJ
A2IS71XY6wZlVClD5sAa14aqCwpCk4rPTgxnItt5zXO+p9czobDb0WjSMXqz9gjsd1QlbA2nzhJs
RFky8IFopYW7NT8XZD4G7R8K+gVmUbwK+DnyhUVHdCWN7fNV2Eol4jslGnrycn1B1dk+deVuI0SS
BuoL3w+1j3rwRkS8k2AFj2mczewnJUtSBMGlfFC35AylP7illOaAMfXellt/dTcrOQAst+T16mX4
qh/imUmdV5ZaENdhHA+G3vUvC7p6hi0Z7HpC5Nc19bJTgqKsepd/B+tbmNMnrB0RbqXIX/I8t/5Z
BoYAFOURVGOwM0ItnGwY+eex4k3kf0cPPifZ82sHyrtWFdvp58mz6ciYL9N0gXZsGsilK/znUgVj
iiKTxk5bcxUqiJe+bV7KauIu0J8rqrfVDH/agiULJvOtfEzQubQNFb5mRskzbAy6WtD9/z1RLwm5
6jNGehyfxhSkWOCkfAGkx6gfHd+LMfUm8GP3199g0wO2UviMyardF4gCuO7A5KHq661lpFTVHuKt
b0bFAP1RqmJKWr/Cc+NNhGcNN5EeEWg9l7YfJjrOqGt9bdzGPg1zxN4s426KDQ+lwE34MeEQJb95
O1XbNyUlFMFYtoZzWmES6+ShBChmd1G71VtmaqgDPAsQtZDrAvAAb5A57MWlt88uCznFudaTpR3y
XNV0I0g00VnFHD9RAoqugdNTyjg2JugE31ubiKiWyBnX2lb4CGRglyKD3SaPyn0MkEuoqmGzXFMD
FJ/+ZfzRmXq6oZxDfurNaFlV6OxenMyF9ah4whP/ne+rNKbRYhKQGUSXRtIewW27N3gnU+wJMU3I
OCH3WwtZEoJV8vzQMKt8yGFLMK8g99uLYJYGAH3gwVe+m7reFtwA+SzSjJ9HzvtXHcAOrjE+NBT0
3saJSwtHTJ20+aJvgsqM8S0LIEDHhgd+KY/Kh+JSgryAXCXihzJImJ3WtTcE2qUXAgOOu6KM74j6
VOg8hJM4scuu+xr6D/slC0RuZQevRAdGydm1Sc+zen8qs71S/uHzvkTJjcYO9dxqYDgvWcWLoFWI
q8zdypQhO5T5KT1JLCx10E8X4zcZ5w431TnXMiQ02dLKY8urd8pTv5bd09kSC8dHXG0a073T9oMx
HokMvHKFxloQfDf3NAuslSlRnqA/qpVYAksvjnKQzhVC5WffQhfy54CWgbXek0m7g6uZLzVlBIeT
/KrK2VEhnJj65Yt8V8sAzQw/SjAme/eHgJ6MlByoInrijfBvVXhFh3l2L1BnA4Fm0kzdmnPMyJkj
T8uHyIjL4AjoSgMGJzH/luJwG2oKSW+mZqZSR/nHZevKatyxtvicAKrdtHaFY0hPoc7vGQfdn70G
OGMXysqcG0SHJFxkfEUdCEAhWh6YO8pTZHwnMqWjDRzkkp2oVR7yL32JD2AWVDNociKSnZ9whXeH
NtsToCY7H265i3TBu+n8j4KxpjX2r35kunnEVxGLrf5UolTTgZtaQltcbRxE9M4n2FUVFog1lRup
h+38vc7KsbI/mQL+1lDPz4NH7wy1Fxe0gjmvWgCzb4Y5DSEaZq761BCQCbaOysMZxUbVmqsy8/NM
rCJJeqJIH2MVdd/TSZu21T88olNHWenolGYYod+cWuh3IZJi3y5FnxQJDSvwsx2xv5RfArX3HnSf
hEc4ykK1IhUM2LUQjJreiq0t5Y2INodrm++JcMIasgGiThM83tQPyFY5w34iHy9xTJtOidtrMyBo
mLdWWaMflR43UE9LSTDirR8X5WyCbV9H6zwywC9MSoTZZzPOMwUPTvRC2NnCQlOSVl5PIbhcPm2v
6vh/edmLiVAXURmyDyoSvyVqcxGJM3Wp/IFHC1kAWy3qXG42GdlPh/TtqQvPDUnG+m8+wmzOSH5I
rDNu7HkTb/Eu3iQIVviUr1JKh0h8nboBzjvR2SuWIghqfsyY3a/s4PQD1IRTcEfOfVsUz2vxQAnp
JjEdtsh7AS4w79yIYGqKogfCNB9ZsL7vpLGaCFh4RvxFSjXmZnXX7KQvmFPRcSS3zNhStoZxbI+D
rVtzkQFeOSkRxrQiDijtovCRpae4aEsznFkm+HCONSfC5vMAc/6bYCIv9ylGOLXZOyUF3+dNhjYi
5160YBRqW49wtYLW4Eq+/+tL3EsU6861Z/0lX5Hh+y6yHNhRmXdcLhKfbE6itBrrKhEpg6ll6uYH
7YHcbvt1/4hU8z05FU+Moy0Ki9pbP8G0IgKdw04hWguYAoo7hpK2WdtxGJGH6/Th7zN5nkpfpgfv
qKX2bcOAyIEmNE37vEvFcrGU9HlJ6EAhgJ96yOta54Id1eL07vlULn/cWxz+6souVD2XMr2Vz0w4
Jctf50nSlW3SHC9nawUvP2nHqohloJDkUe6hggGnd0LCBeUAvs5Wa0xLFphPdjwCVVbfD0sYFqvW
HNGTyaFzT4PtR2499hs3Ivy+Mq4//ZHOMEcr1s9p8j5Qmc/RNyM9AX1gj7aBjH377feK3MtD7DP2
wsgi/Poe+RAGvWC0FCs3VpsSJ9DwALsz6Yp/7whDygp5tgfSDlftcmXVv3xsHnSHQOqvV78XBM+d
jXJN9DwQr4KKpLyuJXRHsEw9EXyMTLUQhdmkQuJYTyuHc1DFk0Aa1jNlmyKMkBvB91TjeFH0EhNn
DKrV4pvJQbK2sv4TIF0+KPSz6bkagOPSg3eXqAsUjt6fIaofD2NkBxcsiASSr8FXSChoVteq4C3Y
DBsMnhGWrbQ7/rxuWFzJyJP22hF+pm3j7PByXa5ucgeQO6/ldCBiCJX7qalRKgOr/Pb88lZ9tPUg
6bODX53ACouYCbJ6uA6ZwbJQSn/yDQyMMmBcZM/wQBiYLSEoL+G9vUIzsdncM3Z6NKQZ3BZLMkCc
Z5da/HdZcQN9ZxIZBfbcgyHaZQ46TKdy+tQ5HXwWL4qF08LJSth5WcBQb+gprWFDuYk4TYy44mjB
PxPTp7Ggl6do50OIvAMCZhYwBut8OCDbxLh+Wv7NfxdyzSoVb96hvdvPG2MH4HRGnYC5DrDyS7Y5
Toqh56rliN4cMFvAZHbhtzjv6mboW6f9KZ1H72K3dVn3gAN5VZKIY4gUAUbV60qnG2/hawAkcv8i
qSXDT1rzJBCNE4h08sW8yXptm2XSj6Tt17F13eaZVgmogdryZfg+EkXEnlf/9LodRtmwGQcgBkAV
A+rKRHiXnNxe43ToqjppFO8biWIOEpAj0j2bI9gSYlbLrDrOQfiHVGL1o0b0Zi9Ig+/4qj5taDJL
VNIyoD87Y4GzRRq/IWOYkHWNon2/bcO0STTKvQWB0TXf6I7XWzNL2lbnM5EMylNhG3UiUIk/12z8
pSrrI7t4B/6UPxY/0rDj5OaQjn1TyEHIO1tlBkRWojissahhtmoJmX430SO2JJBYMI9pq1yVEcW4
n3xarwCnNPkjmRxsMnk6cZ8o7ZXjFt6HO/aebm1ocg2ATNlz47kQ4KALFmcyQ+JA33o064rBTwEQ
5m4RZrLn1Ttat1vD7XqfLkq4FHyp4W+w781cOqbSo1iKNxT75XaNn25K1Tk+bCdrsRWewS6pDSp7
5Xg6lnAkE1U8s6NO1AUsJcgCzuduNSZC9DdyEtgaTqzxW7cFvtRFGAm5vbbpQVWJKiu2ckBilpeZ
Q08LeAssh0Pypjj+8VjZTgYhRFG4a7mgqA3jnC6AG79RhwUp8BYUFfA1h+cKd5Y0N2IikJP7flUb
1+EyKnF0BYGWAPcHF+hgORJY/kWcFaEKyZaIeixyF4GC3oCZsorbWjRDuHc/zbPNOLkYPlUAeWEY
qfRzg8D0l0p76oh8M9FEOK3OVnv2yhY+OB2oRLlk9UD5Hr80poLOuOteYEiohEYjVBE8ZYVJ2/08
MtoUHe5LJnrwXh112sTry5Y1uG0lVBSHu3dNWMETQjfnwXdLL0j+hNhCndTy8SG4gVG6ahnbeqo9
bIQd7KQL2OIq5yWZ5fCX6mVgYDo8gp5YGepwKmHIkecCGc6WruOTABz1MXQRX0dQf+10Iz44WKbM
o7qC0wyQPzMH+Shqanv1E9Z4/UUdHKfbuGzYnSaTMTzZugNRjTz/h08qk82fTPNi6zhOPQWnDQyD
vQaPthSdrdDwegbjCjg7M5ViEf8LE3XuqW6coOHs8vD86XirX0qSKMZzoANmtUEGycqGwAuX8GDD
ISGTRKFASmyT4DpevKXomgHMKYPPOTJTK6tnF0tij3+SEKEwYlCSPzYFHJ8aWP1Yi0MU0CB3uk4o
uVE4VUWcccmnYBDyDMmekj/8hAbEUEW+IcjlF3vM6BHDyG5bfYIEvp1qghK9JyeMQifhnip7mjdB
CWwvLs1fSNB1Yligtye/VV/Vs7WxdRT8GxOrYg8gNoNBbcZwZ0kYSsXAL5AKO+lLWCO0LuKpChMx
eUQdXMUOBFwit6tYqBEvFIHgDyV3K05nXGkvN7DStl73ebMH+9KKK+ofSrEPZ4HHp1li5RWya6U3
MbHsVLHYIevm9PvtByMpUKiJbKIxqImkHyS+Rx2hj81jlnLefkTjpsWJMpSL4yO8G+lt5jSQGPe7
hAbpXO8BePZOneBI1PlOe9BGoMgOG290kv4Ib0/n1blixJqzzyS0ihL8Qe21Fe+mHcVPgCSP9p7K
2yjAsUi1+v/IXcetjc8TG9pEjeh3gOg0tjtgCacttqLp/LdKOJV3rq8SjPCi5c7xLPR6umMKoZIj
DFLnsWE4byA3etVvhDZ02hiqGLwIvHNRMUS41+1vtL/CoIL6XXLGQoEKyijDPBn7qYYj+nGpRgnq
tzT9bnCm5+Q/c22t9IvcGS5fYi5frTmflEtBkMfGMsZBeVayFdY108b7D6FLS8M1fzpF43G+6Nab
VGCVFt8PT0pxak6eUiXx0tQhso1rXje9jS0eer8fCkju7ry20wRBeFreIp2uIZhxia2wS4CZuC82
rfrdWivEwk5LtJzZdJZB6sYEDTdqJtkUXzLR9qv7Ukz0hoCvYzk84mUPZmO7cGx2KBrurayr4I5z
k9wfgRp9u0VkJSGXoMvrzusueiDhc8awoE2GxGNexpZNTt99Uh0uswlntZ10MxYZ0WgvqRJxebvQ
kAfKACWpevW9FuFdgjazZlcSjPXx5x/NOpFvgIfPWKRasSs29x1+TVAF/AfdtHsAdHgznxccsCR7
Qhad/Ubi2G/gWtn/pay1nhWs7K12sggHsUFFMZOBSd8nfxUC6Jz/oK5vIhc2bgETVV+lwSO9wwdI
ABXCTJJgz2sDL19TwsXdP6Zgj12bm0vJqHhKSoGCQPA2cv3hVqLY6TpDAruBh0NPt4ZNTdxJR2Wj
GOqVesajvb6tWY/E040jGo1r3v5JTDTCWM1RKUrn9G/Dr5gQVxC+dpID3tJaIMu56nxd5CScXYgV
5tZWuSeIiWNdAA82bhp8Q/qxI8aABJ5J4DCvZoq1u9jLix1tnL7n4gVtXdqNymnbwMN7fh/9Dzc3
zyyis1uIeKxCgy0Da0iXxbuzTxDtvtRfuFFpXy7xy7IYm6dvXr2eaSnu+TD60MxWKLxjs9YOkTKc
Rc/JLIyeuG5ObMh8uTm7fK7Ijtzk2zga63sSjSUNYxy3G0VPpCsdFLkEzBnjS2QENPCetH0phuNW
M/Jaeg38dgTWCy/aMTXPzIeo1tggzEzAXu7SNlltduSgiX/NOmNT4ukWK7FWUsWeRHDBrX+bWNCs
ujFBcVtoLz7XPuGvqcoN4RyK1Hs0riA4EgVa0Aj9KsxW8rJBLdNf/Hg4ncHMaEiK3G+ELLay9mqR
wOUBnQlRahTCZxFcPNMEjkSoPVzxbjluyEkn8yecDMnT5oOGvFwB3XNGfOqdXuyyYYTE3aYXTJgw
zZ6ooKpiv61QBCRA2gF/rZxXf5ntpXxM5UcQK/19mZsSolOhEbXDu6mmpi2VBeYeARwjqh+NvZh2
GFYIv4rmda+PRyLQFsZXe+wDph8A7uNr/feJnnjyYPH095OqHuMGMX0vCx4FuiA5FmPFNd+W9SMQ
UgkqLxIMRfgiRmy21K1vT+vjvD5TvgfsNjjtlEqOZUkKy69gsvBX3LSwbNauKZqBARvFsAA1c6PE
3B9ku2AgAD1XHMV01qarR8zH2yPAtdLkaML637mqqbYe1GoCHsoUMJJYl2kgzpSXBCB9FBnzER+m
b+RNnK5EnuJetWGuRBvTxxnhnjcoiuuY9AWZ1OiMUR+O/bO8TZ5njcVFNvIlS3BkXiTcIUY2yaf+
A4iRPoow3AFjTyIZFge9boVT/AbcfB6AthPDnZyTZ+VSu95HLdir3DpGyCf48xmbfxmRTepomQwN
jKOCQ7ckC7LGaA1NFTMISDq4IQbpA2hPD0boLfYMqB46WCMCJ2qlj/Z8cflqfIOH9MPkYMJ5quk3
ydjCX/KCNGuv9zpJWUfBA4gxLBLXDOSW+s5sD/9bb++pDf3yOFGhKiiKL9Rq6tqexgDNnVQckgt7
0ECM9aJ4h8s5U0D7qHfaakvzhpeM7NU2OOoT0a7Wg6LAVpajlyPUjY9eZYMsunjxuhF8x+zmoQhC
V2SxbHIU56mcoS9YcaYansttOl+8BAMdQ8XLRfdIP6wK6tr912bSGAqfcWNvSsPQJKBeGvjmRSzk
bP2FQ463cVSVcNG3EODpo5U2MgxlORGc0QLl6iBqYyq7ZkRrGLVYcstTyVoSdkDIdXCL5NfGLdFs
trAY9H1OQe9rH4My6l/S6c9IMm64Gh+n9LUWZ3sXBFU6C5jdufHYT0/u9deHFkJbO9aGXLfIkni2
IZfuzLO2eMDgXAUt7pzOshm4eKBKaRdluX0kv5q1/Gg6DMkBN3Z33ZTW4OdAq4mlt/Lks7SH/StP
NhPq/Z3ZO77V8ALBiw0/BniL0w60XHn1wol2dsc/n6ZADdY4a2Yw46vqicwcuMjbfkfIU6EiR5Et
XtvVi8gHmEfKV+0S1vHX/JA7Yw3UkcaXCECWWs6DDaLFJ5DE+BPYXv+nmzxez0TthsQEEsAQUcJt
ONHJ+Y0LVq4Bc2X3WXMFT8q+Zmw3iqcp7r9ixY1ggCus8Nlx3Eqs50JAAIKZFpCQj/feSy5FQmx8
XB07PQnatbLa9XPQz1IP24q58a1pu8uUpBSQqXB0R1jPVLLTtoLMyU5IZL1j5ck0W6k9dmIWyi1J
SofYfxXhKtmFClbDxkGCmB7kC7ZzLb5N781uWSzuibGBBLzX64h8AtEr0pX0kYbFrNZZaoLuyYYn
JmIVVCQSEBaE9fHpN2wHLu4rHa8bVenKkUGzbFCdf2YPlZEqJB6iJ7kMNCWb/6cK+rPJGvQ+n5Mc
esn8eRr44GX62YLkYKRIoHqxXSooa6NCxaz5+yvZPfETSMlcpOapoOyyVoEGlH7uzhk1p8x3QNxv
bnr3lL7DtGKaattMRqvarFfKdNGyVqtLm3JWlpfb0yrXF/FctlOrfPG6A1y5TA0CIpxmg7QhNhJe
w5sLa2BzeyIg9icGiU/+nu0ff7m9k/MXGiQihIj9CTtNvDBGtHYgRQ/7ITU5rn+U+Hax4OB+Sqwu
b80A0EZNpCF34QDq1UHfAwUxxzd3mg2+fETTniQPLbywYpnTvO1JrX+C0EdgbCmw1CECo6BcH17w
jxjwpJPp7idnuOXyEdXKzX7jbHOsm1Lo7+BKfCmA9J1qdorNPXRpww651dzW87rLbFefrYqTpn7G
sGv21ra+aR1rlcides26JNlZtUd6ZXnUTb6E7UBemb69S5Vg4VUSxtlBGnnR0NpJUX9Jr6rO7GRy
eLxarhF5hYZYQte05z5GOEJxWvGt3uD/3B+7N/4nI77L5NnNxTYo4xpNDzT8RJdx59f1l0t3Xo9u
1jknWwoY28A5T1GU7oFDDDLZqh88HZ2S8A7UQNgR/cZA5EKOQPeElNRSKXOF/PlgUtknAec9dzJs
NlH8CJv9WNx35qghe74Esp1kxFass7dziXcQ+xZr17jc/uHtWBvWJfjXdaYd49lKPT8EOzyPuCnG
hjq/IHms15ApuB473lSDjKGVgDt5NhPIWEKELiyEqieXQtc3WLe3Lkrc/4S/a7GM7TEaIbrTgKH7
Uirg26v4BPDxiQxXLGysvNB/yyxTpdtuIC6qj/rEAc4hA3EVaQKXb+25iGmT8yyY9601qESBzoha
1nwuRemb/PS4oH2wd+H2W4NlNwme1nhKA7j/RmioT9XiIuiwt8HQ1SMveCQUY5CB0r2voaBqyZKn
ugPq1R8SwY4M6urxtD3IPbBRm1ki81xBxPsBrOvHVX7ApDBq1heTTvT8JigUbYw606clEzHvqzLJ
oySV6HSmsfA6nvMR4gs2K57M9GIAZvLJrB5Tx8qgdqDSEus4hlEQoo6l3sy43n2TiKH8lSsualDn
SqeZnveo0fib7O+DdgBkLjVdjZtTZlkAJdokeNArYC+w4rl2bf2Mn3Odl7t0/vnDZu0i0wqIDvQW
QdGZVTieovJhkCvBs/17FsO7DmMgyrSKG0lLHnzLz7tGrPyDYtETY7OYsq5MInUGCeLTBSGeS/B3
gl/vwyYZEDonTFNbjEYnPLk4NgXT6a6lvhdbv4xuCEzEqdgHlV5kBd6OaL6c707cQ/apU8LBG5U+
/BYSjx/lT1K+3ZaUiROz6Wa7xXPx4gJ7NLrJKmbnf4oBH49qP0Q/gC5kxy8NfBzYqfEatOs30cG8
iesOJoEA1ctnjjBY6oxN14zksrxzIfrLsaZEktz/lT8kEtXwv1WomsS1Z+ccna7UC9FMiNhUgCYZ
EDAt3n7FJbgbE8m7GhOSwqXtNTSyLSDjgNg6fjy6JMRjFG/vkJjJ173kPCsyr4Akej3Wxt9hNOkr
F2CRc7ZDicHEZOQQk9VhpuKJWX8kB392EWeZt5KRtPiXAAUUQ4Hsx88KbWyRt5oG7bJ+AdIY9pkn
ffOD2cqKpbL/vUP1dLLhIURZ/cGHWtTxU/n3NLcoS0YLV6TBFDmYBMSxYP57ZitmY1E9JPVj+QfA
SapLxpKos3MgEuoHFKo8OCH3t2Wo+KZR+qIEpeSODEkxx+ht1Y6gBgRnvixW3dLVApJjmh9XKmA6
A52OCFDGrxEVVDfs0e2KpWGdWAm4VpEjhl2KihsFiPug0j479jqozk1942tAU1YWE1RuCon/AZxi
okaW8/H0KS8cxKYOHMF5bH7yu9Q/i0hPWTQ8L8qahjXJTK8kLwzZBFAYemijbW8pwqGFp9YqTXRZ
NIiBcLpxlGP2BvH8fhDt48OHoJdMcrcjG1OtIWkq02OgDPu/KUsYG6M8RVUAZgcqm0o7SRt/tjKm
E6WdalblPEVnMkfl9WPNMBMUe6Rq8ami3pni7NKj56dTkuwsIZUt0NEEfzFfPr/11FXj4UI+KbZG
T/5K7Oprm/4AY4/XV3hnjBz6urIupBE2qwTFNv1VTWXiZMfc5F58hNd+Nv8Xlf7ax+YWEcKJSzkk
tckgp/riUgoKgdrp9qlT3BZu7a6fwQWmO/RRh0MNSUxVzlqWFeJbgnNp4v8ON2jLAr4EdSQKCUlj
O/d5yTpZUW5AXYhy0Hb8589oKCsuTCjX6qdNFaNH0YsBHmfyV5AQgBha24QPAokIQtdCwSGEpu2w
A1O8JCcjU7106hv1w4Y5WL2Ewti6zos/rrS4400DKK5xxLLJSFBAntBdM+m26lkdPc3QcxQBwSnX
KZqOcjH/cZlYUTl97Z/uWGSSvS9cI59+nyHBq+2Ea8gV8QUVeoPRoprqBa7PK819nxlwnT2rEqs7
DEnPKDYyZxqjCHJ93Efds0VuS1m8UKLGifIwupjpPVaXNMvEcwi380taH54dvJquVlFIPel0ncyE
aqhndylFNALLLzmrx4lh/zyVsK5oZUrTpLyXh80gnyRG0oEspubjwGKC+StfZQy5bloUvEAG4TTK
qjvPN2S2CHAOmhXsuHWIBVJAmK3RJtwU+QZgAa+M/LM46GiXdskhn6eELye+pIBHWAOjY9M5IPGR
dnV6DcoueAS5s9p7WE8m2lPJJmrDpmC9t8iW04+mFFr2+EZ0HrG8hh0MYLRsdkVE4CU85XLV+8ua
swpe0oCNVZTiLEPq+qcK42l1t1ZyLDFMWDJjPRZzY6vHAGZfY8A1IlPHtAwLSyVaWygQZoKay6Wu
lqKfZ0HgOwL5n9Ry4uZxOqmemibbqwIf9F4WeCOwB+Ypx4SIk/5Xlzld0jzZsI7XfsdkuP3DIvYT
GQZNpnhP1w7t+Br1jFtS/KugR/N6NSBiygI2M1g20H9wkPBbvAScwYQQ33J7eGCOfuZ6SAWy67Sa
NTwcCzuMbBN9eXRKsARABQW9Fr1dh5aZuGz2rXsfE3VATcN0DKk+KyyQK9twJwCnkZcx5yjQeK9r
m8wibvTegq10FaOmwZ+HyKeYbyqfyg40gNh5zQH85MYqlpo7NgKwSbrTrj+1yfy9hh4DS/aVP5BF
ethMeubdDRISFcQnAv/GUKpwXcvtEZ41H65c10elg8QG2s0FkjyTBGxkUk+iggNJQqC1pVBcL3mw
srhPhUlplqZcvIcJU6kerZagG7KZ7mVahoNYMDv7vukHn/23HYo/4cYpGqwtZnnv/fyvttu7zU7w
/2Y1kGmW/5b/mEDSIkGouJOzpFNHuv4cW8ZfF7PVWYbQoAA3AqI/+EqEimc+KqhFb9Y6FB8HQycU
i8/oT9PtxAmnyhV09wz8NdsYbf4emOXC6TeDTXSy8gaf6MMGxH2VJR+aiYt2nOFTe6yJDaUO//0O
mcsqwCX6GFPNuE7YJ0D5dCnpcdhE9E1ncNxRBFyEnKVGE7MB9RLqEuD2J5OEcbhTXGjUSQTcMpmX
SUd1ynFcC+NJj9klgAAxs5OlUoBEojW41x4jnqloeDqUAK1u1xFzsCTd88nsASAJr8u6xyq4aEi0
Loiv7mBKMAkTtRN1zlsGi0M1UgoZqXLPU04dLOo5Mua8JUS8c4msdfp1HPnGyRFy3cpYvoJy7Jai
WSyEcXhvk6/LtLepwMGGC/y94s8WFs+SPjScy2y4O2htZCtbsCEulN+aAu+tU+/qGbZbZyCaNT+F
DtPYeSaMmqRcH9bE85eutb90EIVEGvnIgUmQdRlHjVOwelDMbLYEjMV9zvqV3xfM2za74JqmJLDt
5VtPP6vMvkPIT1phoIn18HgcVRrRDTMWogIV7JB0ZZAxqKX2FhfF0YRq7zPEDBi3zxqvfdeGnLva
tCTFE7lHJKEh5CTJFpU+Ji4t96IrWbfXCxhLIaTtmFlamvtPmrEYllZY4+NS0GAc+3whWPrXDoq1
TH2wJP2ZLONjdxBU3wFpa31dHKkhW1HeUR1cjvzP2Dpw/ayj7OkwCtPERvjFkxxCVpHwsKvU8Bm4
9LTMuFwyoRrwRN+MktLGjnz5AemN0oGdRyyCo8BAulCUbOiqQPFZCmkrNoLKERgcDwhW0upc+XTR
GZ/y8ME7YwxMHEKwmoZu1X6M8L44Xcc7V6JgqlyHh6Iex1tYLxSoM2TVoskraxzgMFkNmkaYoqjw
aMFJ2T9Z6f3O5aGQ1g2DCrJCwusMx23ABSVUCgoL/DdsfCctuH27/5aX4ldIIYVjmGwXxulo1hFy
1CqnODJSZf54N9UmPref8UyYKt1GAdAI5RzZbS268TmiVUitku5utGrNmlSYXqrjakEbXEi8go+I
9rrLBXLKSWbrYCQATNqzPOV+2c5/jGlWjyUs+9YAvX1C2QtJGu+Aiao/wI/pqp2ATaVqhfZc4tKE
FGX2Y41YfO6dfcRb6dH87waOI/VIMW/OkCTpEZ8zCaGkKWPAOYaJsPBb5DNlF8EHIOujSDCu7dsb
IXk0ZQTGijlPWpTukYg7M5bmb7012A240g5wekNw3PUvmJ03bn9clwD+4Z/bAlT7cQg2dxa6I1O9
dW2YKxqKoV2B3eP4MYJwBzDyuM3r4EYtdIbo6hox3oeWUV4ogrYVhv91U6dlhMakqZimWlYVeCOw
oRth/PMXhzS++Si12hX+yJhiJC/HT5IBmipJ9MArCb1L0H4Jfd2helyM+vmYRHpLk2mPdvzWn6Jm
HWL6VHf3+uRRvHH8dSeZx3dgowYJZiQ0OXoYpjh46Yl+4ol+RV/wLEcpr3PXCHHE97BiOMCDDwtM
ao7eT+jP2T0sJRYWFxKdqf1UZerzo0xXRyGO4XrI7l7a4kYvxklIwwsQBQUSRAzeFrBhPulGnFPr
50sdmKDqqikrQJ2PoIugKmMTaenrVzyf7c/CmDVScdeT1dWOw9Lw1+rLYt8i5BbdNKeDQU3GXeCs
1zonu0DDUX7yg9i7UISokBzz9bw0zWnb8XU7DJx+Ec/ofm5990Zhl8ygKpqN74Ic2df1tKzk4nsG
c01Nsphd5Hvpa83UZg4ZrJEptJ6fzd/1wtv+Yq637zdS7cQVriOBINgpEqJbBdx8vKjFFOVXoO/g
YelNtiW6d0sM1YDDDAtceQA72Hcte+ezMxle30W8CsljYs3glKgOo8M7C7dKeWiV9vpry0dk9Vf1
CN4CuaFouMEj3Ho1dbHm1JSGmKue1oDxukdBaGgQ5BFOeM06At9lBDbeRbVYIfJfEnBywLUrseLZ
H66fO1fQ3RRacujF5mhfD0LHY+xP/vCVY27F+H5YfGRFJJvFdm68vbWBWfQ7se68P8dvCSUEIV1G
olzs/wHkqO/PUHj1X1AAzsDiIRKu/M34YDD5arwdk60EWCOsYmKJ5DVjC1GDNRZZ7xf3KV1YPG8G
v7aGHAl6WqXf6aqJc0pobvmX4rOHcajvfdJ0bQeH7+NttzGTZBWIRaKuHio/3AnkTE2Sprrq4n6P
64AIsMsh1ttld2Z7yflcHhI2CWg2YuU9obYjbGSL7FcmEEkLnTtECB9XsAes3bIjShxe8qvsYQDx
vhiIhPnT+yAjmfrXUTgtTrj4t/uu3Qi5e3O/LI8EfB4YagAm2gkDWqgX8+W2BTmPY5q+fy1tEYIB
kMR8v2ta3ZGXkY2SZFcb903mNaPopkgc3nCZIS2s4/rTDGmxeQxldrUI1lqIcVKWHn6TCbPtPd7o
tQ61JPSWFcAsLHrxFUzf6KLb5Ons3VdA/tU2XWR9BkjGOyonMfyAd4I6JB05GKjgaafAtrjR3Q/V
BNHlc88V2yEQG+BSgF++OhZG7gnQBvhuNdnACPklWA2VI4AMgd2U6d02XAcg5jeEyhKs1+HQyyRY
e/RNu/5ns9Vejc1DrI+tVBdJb4X7MezVewh1lRRc9yIbDyoOVvFVu9NFyf1Ze9li3tWc7AQxv6n/
d3boxD/HadewTPxvoKvk/27/qUEwrYSZPDRXQHlLJaf82CEuCzcuLoLeyXt16kmMCQH8PE7hRrHr
o5p+IwfmcqbBWM2BGqX4FpvkeUneQp8SwIdBK5KuKIDFe7Cc9sDrW3DoLT7v2Be165IAZCoN/eWK
sKVQwHEo0IG4+YIxciiwbjXyd+8tR+NQIyfLa7k/beh6382qIl7bquRA3L8ILhBp4mm2Mhz3Cslu
yqOvTDbULcl4SoeQJx4IBfazs3ps0c7vzs11Nn0D1UrRwSJguvX+ZEdziTfuUKCgnjQsiiv0sL0z
6uVh5mBMoyHL4xPhVxt82TMvrvpUsLLnxTTXtTzEkm7Wr2at+NlUTpEhORpy9Id/XeTO8apGoI/L
TCKJ5I6w1CDe9/tPL4aGGHctHQWWXhG7rBckFSwqT0696PAT/ibLaNG5IGvPnRbaGg9f7yInpKMi
xv9cJYgMEtKFpJ8CP0S5W8hqUQW6Nf26OGX6HENo/70fSM2pctRCwAptKPQNBFHoRTCT2eEYo1sC
mCj3Pv8hsN9J4gHHaVb9NrkLPV/eJ1Ic0Qw00ZE3Jn4hN2f1ZY29SPegevD4m3ScS24Rga5m2Cc8
/jvsR5quthIQVwUUFQL5m9vdZ5BuZTVDU1xl/+jZpgL9Or4qZDNmZbPBV3c69wrHR3zE89tgDaCh
PRI6ihWklahtRh6XgSjiBtkNmD+ryVgSniQHj+Br8LXC7d+4p/fjjq/jRP7RtFtXIU8hvirVy/BP
lyAmTAr+lI5+v1p+huCl4AiJ138HtwHZkbzPCEwhM5hevgHU6+XH1lf8kWAj4j3nkVw0A6bkeQIU
5WpLpFU5zXW6RySoOKEiWe2UK2LKlTBmAdFaULbw8F4WjPxWUO9lpfflEYLCucudEg64L5huRVNs
zcQnxDbuqJGH3w6/xJReBk9A0ou4dxgYRXNh/CHWVYwucBcHtYa/T7YbImhyPzCo+X8cBHmt6BFy
cJiJSkwdRAPShQL8gvs0iUWzSDFEq0utM9q+4Foj/VebxlCYk0ZI3B98lG8RZbFuQPW8/scdf1Aj
mC1lk87fr/MoGtiSpwdjnfA2KASjsk87XZ02Hlmkuh7XrFlq4+45JsNgRNHg13DQxYt7Dx/ZTEZ4
jx5mSj5s2uX+CHbdzYqagnn3aKC1X1+ni7aKPiyI7Z6BVzfiNorExOL2Bxkuznfrv9ULCNSfN1tT
R4Jvir+ZNcH85MjRa13L/uFeW1BZkiQWdqW0GgHpHUXiKr6i+y0jaCON9esq/CUJzMFQC0nrSQ0N
zqq4DzWue14ClSdAu1eEM1DOgQBzkNXBr7K+c17MPBRlD1EE2X6fJ8huFZ2/sEtPUVW7IGiERfEN
Wq35sv5KP5o/8Es/L5qIJW2tXIsrtYsqbNuq8NaLUGYDNY+YLaPeNKdqFdRS+dDN032ITIh0vdIe
1D6/mSmXJAEJiW09assUhp8nJg4fzr3pxVIB1WRHvK6NWsUQIpypKHJzCY/oXy+mXfhnorvOe1n3
p7y/S7pbVYLwGqyRniyPkKlApQQBAvhhv6Df5erYjph462eAuTYtNQ+/7Exe2/5/dpdKBcdzl3N1
miMT3RJnBh2ydq7XVpGDoyTK2PSI3MT181lljBBoFU9ci61vOJZkmSuV1dvzpEyOi5m2JEmorr6J
wmb9q830bd6mHEosftTVHH0VYTf0rP0aZrt0jqWU/bPY2E+ZzABoWhU7i/IW61WI8ztjYh+h/5s1
4JLFJo0vBaXw7ZXLIeQ5FdolZE1hUy++uUho7v8AelQ27SiPWTyD8i5xS86wnBStJ3JnuBDpK9Lk
O2j5e3AV3RJx6JbPTUi0Qvv9VguGVSmYNda09DZ3mrGoX25Akl22r4x5hQnZ6fU0T3Pvgbv40mq2
lpE7AYCBPYfoS2JWKn3eGG1FpEuurnubkbfxnpjn8Xw03hh5GZMYST12Z39xa4TaN/Pk57B0rsnk
LtRWO834vW9Vy18PYJl3JvIUHrxbsqXKaKl9HQ+8+qfEYJz71fRie4GIgKGw0K6tXLlDi7ad65Es
74c6LZ5zt+8oFafcPhskq/q4OH6k9dzh9abYQMBsfIS1Pb080LXg1qjf4JbAcxVpeiSDP2CwIBaA
Yl1lEVOvZ2/hGTCjFq4oUowlClCZaBplpSwgiIBtoHY77VmFBqxsrzs5g6NtKSEVpIkBSt8Aoza/
z6WgUxhFt4zRvD28YO4yo6ZbO4z7m4SCrYaDqxqvQaMQfDq0dxSqV1y/mfht4KckOv+vAF2eAHmd
L4jeXtJifFQF98ymNybw5E3BFsufB4awZayeUVfFBMzJ5Yfc1GXaS722HRNSOO2zUkJDhossyT/j
WUiaW+qJOvNw5Uii+lJf5Y82GqavvtQEme/a2CTBOPDezVijbVMEl/pClWWxSHtSBZR9LkSPd1pk
4v6gQ499HwSvCdQPSrk1wmstRI8QnDIs/krAuX6seKMjqXxlHX62AHphkotzcUqZBagAPvqHMKtT
xL7gZUXhDqkOXgjr/VH83amx59oDEBpL6fsFFIeBuFY1HQ4mgsBhmXQFSG27BG61vsXs/ecCk1it
23ZPtsCymxQ9V1ZYWw/B5yuM8ZgOaMExcFP2zg+0LhDTp/sruSewPHhs+shkIJuw7bmUiMgVTlqZ
k5AzbnmXCx3TJCaPQckIk8h2TJxpD9XEvEBDdcMPNa98rNYQu88zIE2QO5NMY4G86Of9er8hUAoS
buPXTOI9Z33X3C1BxDVAkZESlSQx3bvpnuMFmqr7RQnN0Of1OuAQ0b6OuOe2DtGgwY2IRXZe+WpJ
/uEdLHm7HL7Syb7N88LzRdgDqce4740gPiuOlvZf8OU6hQPPQlbuPsXZk+cEkS8DeoWxbgi3K2Qz
oIoY2fRR0cQgpsMg/WwvfdIJZ8euG9ZGVVMb9pD3ks5S7tV1L9ROjCsEOaWEXxoiXSiO1fERpZqn
jEg9JavO7l7X0WapzMoH56dQqjPe/G4kL5J8vRj9g5JlsA2CN2LKxiww/pG2CzKmHW6jXIKE98MV
r9ysgnxLz4X6L5tznO4FyOMbjpUhabs2a4F/suEqePtT3w5S2YwaZ51s0meehVupbXp+JzRUUHjI
Ncxt52OshxyRpb5Nj7BTLhpmt6OTK+Tl1trHNitl2EQpuJVPkrukQl6w19lkcVwlTBOzSMkTQQRg
17pDPVanH48hn4lMxW6z1tA4UJU9nyhXzvXKwnmX1iI9PwemsCQ+gsVIcWiJV5m+cxfhMtdh53FA
pn4Er6Lu+0GTAZ+QMjdNpxiTsmF3S9NKgRyjdzqp+8HoCgEkS5VMo0P07XAUoPVky4ffgXuAgNJ2
4Qx2xYdByd81TZjVkrtKi4AfdAQBEp5mQpB39XxHqnAc0WspuabcMfTaSI69THZuzcQNikJRfF7o
cNK+TRMeTsEklLeBsSFUfaBw999k4Te2NbGzf8j4r0JRyJBTum/yQxPWGKmTMuTue2t/45Z8IMAd
/amdU6QUCtyb3VGUodZDvz4ZyNZ+KybYuC4b/nCZpLFrJ418RDKxma0TjocG+wkNXMiM3QOvL1id
qNmgb0TzxIVj0CGbQiry4b3UbkhhSXpcaavJHn+RQVGbCvdwfHKdZMXSrHOpeW7ORZyp8s2ainnQ
9Vtc+guCk9FMIvauxB9Su0UExOS/+n4mwI+gPWc7sCUTjNkD/GaW/HQIV9/pnYFZRYUqfe43oH/C
o2v4RQ7Il0kvmPJCC9ElfUus5iJszVskwsMwaQaoM1n3OeKE36+QvxC/e/Z1iXeduoBI4Qpzeh49
hgOgnFSjTyHBgou7veeIrB5RADVFBRay2Zgs8TUVviTjgtm+qZh/VqZzpTX46tsCklTaKMZvm4dm
njlsATcn7wEzzT9KPxZqZer0nltQiM+8DxWhrhykz0vEZBqb3XrGVqUIq21b59n5pBF0l4DDCAF2
09f3jc6vlwM/1Gi2gwdrp6ahLvnQJShWVin0RE3PqfgVY/drtBJ3gwMNc6kJiQmCWoeooBgzAR2r
GQrUkZTkjiwzpH+3LFXGiW3b3eUPh8uT+A3oU4tKFlRDwDcYAL/YjUIv5a6i0k6sjRNsVto0vZ1j
1D8WtTup+z4vVGhmvsGKzb1NNujBPVt2UPvuLw/OuubxU8Xv1jKX9CA0xZwkpRmBmr4lWC6uANIR
wmdNlzUHscbG4b9Hcwtg6feyaiyUy02DGbOx/lCyFoacvor/I4TUTarYVuWXlsGhP3Gw9ocLmAX9
PkvfBjRWpQJZEoJFnhdTbY6geQlmniKfbghYgFG6+6fxkv2DW/JYvBLxlNtPz/4V9LtvGRGC+WdN
m0BX8giSi2nkoa1Kd6sBCm7BSmU+/1ODt9cacnxkVfLTgLKZqd356TBGJ14FTbRDXnQ6xamWKnMD
jSwAXi3jJR06F4/W53qh5QUyiGeVW8sxu5gXliBZM5gR2MSYREQ+uwygEzBQ46A6Av2ixAEBOKvF
BXpqN/0OEr0M137ZxhtESMJWGgyTXHsrn1YXyW6cuSPHYWb3ZE0WIOSQXNwhoIgiK1ir5cRSJ59b
FbEEBuFdjE0cVqlOqFsIiueiH10qgSwMUE9sESEsOykVfvB5qUA3vz7hEHDmrqI738ehPiiMpvky
jrb76KJv+JmF3B/WOTvw28wWUDXIwgSLlk2fWO5/QwyT5gRfAmyBCawduwdprOIMnBD6AHOR+hDe
PVfSfiD/5ZfktiT1P80HqdXtgCe6CitssNIcb0aFcrnFlzN+GXU4VUF/D33yQwiP4lJP/U/IvY7C
8j7qqxrL8592yv2bvNyulnhK3Zxdi+Li/kPttOkvX9eEQPVj4pRO9CTFqG568Jbsv5CSRl3LN0oy
+4dFbLYF2mtAJ/5MVPeNmd96SB16lqmcdu760G2X8EfDPhIxfFqKozlS8XA5PkRXi4Xgy8e8Ym3y
9IsazngYGR+k82EMWgMXveqtyAwvCZWhZxDZakfyaJbYbwoytiUgrNg9iarrEQgsLcdlxCM5BG9X
H2Kt1q6CBj38hm6NkQkSeOeRmhK7UdM9EOdFjrDGu2kimW/Qio1Dlwa8+bXCmLo/ziUNBhw7/TGd
0vIG7oyDZ7KphEjoF0v6fKa5NXleG4kv5N0gQEmDJPDujY32STKvQ/wep/NhqQ6/Qhpa6iPN+jEN
Z+YMIFxSwILcvr7yIvMgEWWEhF8y5xGUrJWTEwOkQO+YlApLQz5ayMRBJPtACeMRaFsL+Py4eGMC
imv9UircbIRhZzVcoiUPAsJr4LRxNawoGugWx2GlPugboG36VpK0l8v3lNHUzml7kM6UUElB2xmg
7exz42fd43hd+YjFzj2/4DE0I50yUBcPYrlRZQjjVHWLbBoJKYaMFwt8XMkMxj0rWwvlFc4Yv4j2
oDswsPM1U18+hNdOTFa4ai9aTs/WPX7b1lHiTyWwQcGqp2/FsPm4R4LdVjYfqx5diMGckjY6bHwL
m6cCqSXDOWdpIbcMpbK1YhKLUcE5ebkS/5IpgSQ4ZKYxU4MjNk4ZDEYP+VszgYfl0ygsEIouwXO5
GS49A+pers2VbsEpI/NHJj2Scl1zIzmOajDlOVcGhRLQU16czK6ojjyPQoIVh+uK9GVdkXxIjujC
pTn4DtzrUNgW8cm80pb5H4Vl1gGYVxA4nqiaD3+zHyN1+98Nj1jT1bCVNszUKptv/HHOyGw0zTBy
edW7CqGezqKCyPc0+FCy2LqU79fJzLo14yBeUs8fDY2vL1pWw8DpChyQwvRWTPvrYDVPmHCgB7un
r2vEs4iMS6eb0atper3eDX5c+3zV4Wj498J+JAgQbJdECjO57iRyzIiGhuEsurUE7lIg8gpWYI3e
dLbLvfh6m5WljVQnRZWcHuVpBJMRtd3nuxz/bysyMqADzEmGWL5ztWb8CMDB9M8stkXhf3pe6L34
l57brNuzVQMY/bvH+79eO/5v5apC5454rBLjpYOwEdsBd4VnzbX6wvk+v2SdbQIrEL8oEVSfSa+1
/gJEB4gIgTBX4JgYONEcHbAO8Xhoddk3rek28q3o8KPKPbe3ur5cipL7nlewAbUTh8zyGvc2bmd/
02AFkNfoLg9hAlcut6hHvLcluNgyGTn0jvsz7tDnCZy5aJIm6l35i9uukczqCx8V8zOSgdtfGUyv
Ca6N0h/D5Du7EdBXIJWbOaak0EZTyoHqFy8x+eho37dscNKDsH7nMBSNEVCo4RtAyHjFPKgtyTQR
NGns2JHmXTbZRmNtRuJM54zrnafmyT2Yc9rrjH3gE1URwizoSeRu9yrYDHQYdMyl0shKpFwk5Q1k
Aq9nwWyE6A91xd7WssycAibaV5ucMG/wWJBba5gQ8LQt14q7ciIfORh9KNvOyDQk9eLEo3FdyqyF
rZn51tkiNAQJEGyX5x3G8sO5f32oYn2j6v6pzRO2VrZtfCMqchaXHdo7HpP5ikeWVZXLYgXrks7A
9p/FoLHcAS59S/Gvh0hMPqbMfkm5/WAcIlyCavT96ZxLUjvWz9U7pAl2QkWteA0Xuly3VDkdpLgs
qntrJeoS432wOXEEnFHEqGFL4tgnyDj8qDA0eJ8rLgSD51/hEvAs3L3YL9Upu/1eGJWw9RiYE3bj
nsWkPM4yiGezQNLp9FIKt/+nckTKd7bc4+l1OsmU3n4qfUiAXIuaaFyRA6XCznnUGKkOhXsFdgUP
RIgM2IDNo+ZfqXE1aqmlPjK0SnnqoLHNFAxk24iMl4ID8lN425gHOCg5y6ASgxMnEYY/wVuR+uo/
pxELF+tO9G9DAVnH3DZyQWd38cPdQxVLC2U9aCmy2PGeqxoaYotVQljRHr9ZyI1vuI4MC+rvpO55
GBeeZISsweLRxVRuov9IKsyiEtU3zoP6m1AL4d/J2ElqZgSPLP7CPzy67hFC56rWf2RTZksMrnE4
2hIdSQM/faQIUmbo9QP1PP4rxwlypwupHWa/nRxLAxMdlqQdn7O95QBHTC3IfDT4xlxGyp8brUoU
Oz4qxA3BHtcCpjLQfU9aTG14QFr1mZ9GbkhyLKQ37A7qa29zAvAzle6WmmCpfv9WxzyV2JOvFpFE
mAR6TWEdstziYjaltua7XfdBJAAvCTPo/Tcr+SC2VIaV6/NsniLT4HKr1tnGPRpnr8jtcvg3cxHd
gA/hM/ozy3qfVXlSNH4nNL4UZDy2IFky9rfaDzK/5XmLrf0Ni+gdu7vZBXPpo1ym76DWUkushzBE
uBLjJI+vxxv8eQbR5xFGQ4d/+vzmcb645RRtfjfgI0qfusqPRE+wND2NPMTjL7qa/Ikbi8ugVYw9
wW7FI8aXNlEVaXA7AKCh0Ypowvlpw6Zq7lfpB5H17DO4j/2KhAnH1gAmf4+Snoa8klpU2nfUY9jN
qgwJL10tl1+DQ4nvHBLzOZYIPFtLVXSDv9SlJAWYw4FxUZriDFgn93eLmc6XZmDnhxG5k6PE98BB
djAhtVJ04cZhVeBZ/iN7AgClOGzC6sMbWT5Gkdv9anCnoQdL+NeX/vrPYKKBRVe0nspRTIgwwJkz
PctDlLRvNkzEIK2xCpcFreJxb8RDDF/QHZ0TbdaQcDgl01qevReRVivjkRLbhkNU7gIhfceT+C87
fI6mH/OhuvsQRFwwhv+wEdeRQA2MoUhVQczHBzDKdors8xKC+wBZ6pIZ+Bu+b10I+Iqu7Z4mP8GC
Dz2FgQZnfAPWmFo7rMt5nmrCiWVgPiZPTVxzMDLmWzEoEBnVWOJTXyV79qbao06kRH7gx7usbde9
jR4tcnZ6ff2k/zYRb5f+BLSndisp12A5ubJdntREz55oynb26rpYrym89g1D1nzmuRqocIyCPWDy
sRaLsSpDPxLpnDNn/rbU/xXN+7SQZQMMDdRcNftfctfP2iFE0Al2DiWyZ0ZWQeXH5zE8axNa0XwQ
TGIjMoysKer0RIob9Txs10GcFGRCHDxurBsdV2TmhB1pU2RECTX7X+auwiepiHktGPWmaJvniESv
iyCIkqfTH8DsDQoQ/bqby51NZy/umnI9bkoBN0ETt9CWUUNYiSyndZgqLWc504rUJD4wbbJhNMe4
HcpP/lPpJuRigS3Vvia7OPRZC1Wh3qQ0lgc77h8Q+1IUvWEPkevev8jaW/sfQ9FDQXAtrLt0nSvK
nx9g0S/yZ3GxF7RwZk2cVSDTdHlCW72YR1AIUNVRNiuUj9L8fwp05qzU06aSEead155OnBydQDwb
6xDUWureNkZj8gqmth7eiPVOHPcVVJenKMGyJa0cXDw+WWWjS457Epy5bmRmBpaKZXYkYvSwc/7c
VAZq0itVsc8n9ohK8fyMmkdd5b/8Ctb7R10swkjk9b4x46WvD2M5Gri62v88GbrSim381UXpe4ZE
8JkNfb9ZKca4GeBJH8cWqmu9y8pNxA7OIHBOAe1VaaICMKqKgKiEVINXtxJL9yYUwl8n/SnZrTpj
t8XY10bodutHdysRppTls4KGHLHRj6CDFqHMBDT+2kSPPgkfmFxM2d+jty+2zx9K5InJF9LrAXDf
4d/AUN0MLfwaZThpfItBPzXVqCkrM54wdWdXBC5JVMfHa/IrbVGq5bqiBnMS4ocVMozVzsEIB+ml
LivAQTboYodDnOlvSQlgqpPBOd45hsysaT6zy+Yn56vHKTQWRcV6Ow+syK4EZFnET77P+DfcaDbv
d47gfg7p14xOMobhtsg7YcJsXrm1j8Sh4VY9f/3tech/RXr987mSN3n6FLRwkFqkoV126J/1XF9Z
WvPNWjMW5Q7M4axOsfbj87o3AvBay72UEFJsD2sdXQNa5qbxI0MR/6DJQKDZRYYJ9CfLrodNZDxP
A0Kjeycmc94tpHYxsJwQmw4EKMYn6ezH7SXXfL0lWsPVgTtLik7sEASx0wm3zZUn1Bqk7yBIBogz
Va4mWc0wCAZCrckxcGTXUbNZrLTFvBSDDzOgQnSJzYUAb1jZi5wKteivWIK69xFP/OD0imqM4wqV
oHum/BI0Ki/9vFL5tV51fk4VLwSS1yqFDS21P9Pz0FnjH9Cl2rSGGpK14o0+WhrbHBehqLRFI5e8
Jx+GL1MSlZe2WuoqQB2E0j0GocRN6yMfwd37vZeoG45lEyw2MdvjQwHvDp6lj3pds+eGBOtDRwRt
gjGD12Ce4zOrl0W2+kN2YilEhILcAT/JcX+SwV5fskwQnYYnOZ90BMWKsbesrhNT3g4PpJwI3iYU
4bM4iupBV4706NwliXPcc2RdKTRkTcieRPsTwKoJUPYlDHfiiCYzh6EVq0DBFAUhRF/EGmHzUI1H
aZVBpAOlsZ9A5HMVgVg2CRluFk/7Z8fzSl66+pKhtITeHQosVtpbiuo17Vpmnu8QHwkVabA0tjsa
3gPOgsJuJM19WA3F4GyLG1kkzihCoG4GLZYBbIsCgIo9CVX15NsTq7+qSJHNX6Znh1p9vZoRS5UK
PKQ2N2Iw6nLfbMIG5WwYoRZ64TcL+fkysT+YNw4zo0aEIiYS5ttcVGbpXBNfBNY8qF+egVVExFYy
aiJiyXiNxtL0jMuFZ8WEE/DUqum1dxSGO6hhYQUOldm4vf0XuSmMcwQysT5RdTImvUkTETsqFsWE
V4+X1dv/rAdo9OlSYc0sfa1/Uj0gytcFw4tcsOEGaCbrYSLl4kCBHSR0w5JP2JccOqs08Sx5Yqw7
lUeUEAuhj4r2iO54gOILl7tfOyJl3r1BzKEOpTlbBwFa/ilUDfABO5LXGYIoHK8YLRl3SL6pudHC
+ofIVDMhKt9r7Y3JXoZCBi4yOzJievZ73cFpPyotspGNy/F6PNEX5O4B0vPu8G8bFDJyNtT1mjYF
MmOtZDHAo57mWWMD9PZ4M/nvtwCpkAiXOPCG8ZZpGHlN2p5p0UTzdRneE4WlE85Dc98Llr/34FM0
sZz5NHxhi59s99IIKH9LK9lsySv7sJnEZT7Eo9l34TWNf7HtpT3uP627i6J2joUsjHAXeDQcKUK8
6cTtQTShSVf/bUYToQcOSDvzO8za15IwyWF+hj9AoajqwGV6ft3CplrXgtlNfq+SPYSbBfUNQGJh
XEqzQmL709XLvM++DQyB3p9NIdUgPmAe/S9Push5Tap9UwoJTL6X5TZeCXZPu3u59f8srr0uQHaZ
rUqv2TBofdL8SkQ65Mc58khJPQw3qDBI8M5sESF2wKWoQWAZ3nutLS8EtA/dWdMuAtn5l4ZomHFt
KrMQPGeobBYB5EhL9SFKCDG+wXSAl492civ/u8wnq3fGcpPaYDiuoWfvDp4wHNbtQA0sZdgakpfI
pA35n1iq28ED0nTgeykZlinnkEFRodGVOEZaVJyua3NBwD5HRXiMJYJCLolwDOYBpOqlWzjQCul3
3LWyyNADqxST3E4pywg6q5Kv7GQM62idgu4FM6HZkUVaM6UcmzI5p9zjD5Jdw6aWpDWwJeQahYGo
L0dCQkHQdaAGec+f2t2pFmT9/1W1rBZPFXTYM/qX4QKxkd/wbVpTsx7XaQBqkxuOe1nUiL3oX5L3
eFrNveRBhMLenS2ZLdXt9ucsmgmaaK8ilu35dh0u7Jp2hc5mLZXCN5gZ3KZosf5QXqRiSzbbw0L/
gn64oimP47MQ+hiNqT6rDH+EwlNHIvf3riwA5jyWxuL4pdWJ0wrW1kUmr/FV5HSpHeC1C6ZbxuKh
tykbBrT6HU/f13/AUqJ4TkzZagtSL8whJ3u2soHcevk6rD+kQ0LQW8mvBI2H4e9AumPB1sLE/a6N
+tVXzuofOstEktydrbpEJ6kZwWUP74rgmRj/kKxvT3sSYs578jT4EshzG2zWR7CQVZBP7Kl6sdPH
egOr1ElZiSMbase/mwMk23s+PxoihVhxBkaRqwRUGQaVcFSeYwG4tJVA3urlGH0K86NQVlcm7veb
UT4KEGXRhlOiOsBgN/GM/GIiCfDsH/ssEOP72aV5clV4k1yxsUBlbDr+bp4lnd+9x9V7ZCX0odNg
6maXi/LqOsC+MxVf4t7zwb4bNg9/TNpEQaRcIb3QC11Fs8B2/jDaDjEWqGJu/Nxsf6U412R8PDKt
F7r1nv2psUZCADF27IetotOvEy4O96zFn3EHLN3BzxRwKMMNythBD3mtP5HeuZsmfpGWi3VOQ48H
F1DCI69V0vp9UDXCbyC2i/GB9gKrLHQGyhGZF6IL6913JNM5SObkeUpO0KtiUSyOvfMAE6gDdgf2
6otqsdTpe3ExnZtNG92xjanYC2owTa9TEN31Z+T4VTrwD1YmwkEFJrVKQNFo5cEdA4EvC/of6Mp3
24BLBIg9Cyi+Pgjp/ttfzAuiz+eJPg7uQYMUdeJt4ojW50ggtWPHnRr4ffDCe07HQNWtk2QP1SHT
03mLDHCv3xyVdkiDbcJdBPM58rMP2Wi51BJFa//otTgXFlUNh+iRLKtZccAHT6DpULxuO6cUM2d0
qacuCmbwOICFpU7e57Ni5k2I7Rsd1Nbg7XLxTTCisFO8WIVP+PDJvvHeyfEGcUCrdFBcHwpM1XAJ
M6agJV4h02j29owuLJ9D9DtXAKhiP7cWeE37TUknSMNvlTx9qbWDXeK/vzTvCgziu1bKSq6g7mpe
L3oDEdZk5E5KnVcAUWHHO/o0LMg9+TaAwlzslvbSaDg9ass6naswJqHRDG9CZZC06I+1MmLw5Ss8
OUWJfLNJFpliE+Gu1exfJvvpe3k3rDnp2LHFRUu04y75vYXJIVhtCABblcGG1jTKwR8NK0OM/qCW
vdx9hj2whrdWzTXXabS0dQ84dAJxVatBet6+2/65Z4Orz0JsysNoBFjZw9dnZzzkkhqanqqVvShR
2jbgEY484QVUWWbwZ77WcPdnvJZ6HGabO5q4y9kECW9juasIjDeHzlnlumKd7ZMk+c1lHI1jPmrj
BT0Uv1RbNjBtWriGgM9G+PvG3/nYrVJuVmGL8CVwD6m77OphPoFV0jTIMr6bL733BM+I1LmpqEKS
P8B6zOvoWXGVoz28PZRRSQParJquY491eTzWy9jQh3pRRzDRr0P5qj3hdzdX4evtRgLUte/gEP48
PLfzKFMGjMSgEkIEptJ4112O56S9Es0JyvgB7VU547jx8Of87EXhdz3EzTtu6AnY4MNoe658vI6h
ip/58g1QKzGIO0JQFcNO/2M1orWvuTHKtCCBUOwLdzQi9SjKq72gW7+IRStMjQIUYao44VEKOcfS
Wh0/j+b+KDTrxAxxQUDH3W9r49eyTX0f6cwTqskI8mgW8cYIqqXcISsVF2TKFCEOA54IP5D+sDCx
8BdCHoDQqzaH/4itTZjRdD6V4oFSy863R4CXzI/rqSMDWJ1M5xWAGVlcrkQGFhgVQqviiHs4A60y
tisFKWIJFizHQ+5T8Fo4NYEUT0Z+SFJeYsh3ByQ9p3bJRWZbj0Dy9ebk8Visl5tOAyK8as2l7Wfv
Rw/M1lHfArBVApzpUfEsD3wRy4NFLT1vTRr4CW+To3PZrDw5k73TiK26UrLUaPY2uNeGDJl2fGD/
kBvxt7H1eHRx4tcdRAjaseNVAqbLJfvD+Y92WqRldcXM4WhqKPCJp/9U7EI6yyfPKCs9Xg3Al5KQ
dz0NTVNHjEg9/q3lwXUP0xuaHRpuRqeSMwWcrFtVRrjFfXiw8kEVAgzxsx0KjkLl2w0PKtx2djgL
y6CrZUmaeBBt4m1Zx/ll+S3Fv93ZtwHozdbgZnluDhFXV5wXFghQvPeiSD02yiWXj1JYwNJx0eGK
30pbizwzfjjA8mFKxHNDwMty/v+cKblUOLmRSLkFpQKG2vzoAD9TAUtqS7S5KfBY0QBrIB8SKYOA
akWNB4K6yDfZcOuyBuFDs8o43VN1TQKb2eTyJqxuSYlk+mCkCUmEIwkYWR+JjR8oDZhUbEbL/dHX
WckF3g4HcySyStbxtMY+EUxpGLbq7ZkmmsPH1SD219mvMQWA7EX5VMBEqTKOsNv51QSbKlBev1eh
lsl1PInGfhTNsKYswR/PMC4AL4Zlsyr70OHcctTNLj3sRsB0ivCJlffJVOoUBbVeGEhkAc7WdQoP
jRfUB5s3CT933AoXUiyfddU7f/rN/NcTH+4+SEZBJh2/4b3krpBd+zJPGNtcaqBB1dV2YkeEECf/
YppOTBKexY8xXXbdmBI8nu/BSqyXnlqKR3n0e4IXFx0YF+sqJ0WMNBWm9BfyUQYBjrzzIjtHo9Uo
Y1PAf20rw+Zn6KDIzc8N/7AR/+XinmhOqYYHA70u3z+uAZ788mBP9UTeUoAHDQ3dXtz3i2pAPC4y
aKd+ggNdRp8fM0UkJ33q9JaidrjLiiI5QkzLfiQgxMuerpsWKiWZAoFUGKWSqW045JGOPza2/t+z
04qG5rqpOKt30M33PQARtnuU5NsIREuQiLdb4nF4Agfkg+MaqXZrh9iKLMJPu4Gjj9FSUDYKVgXd
lV+L9jWZhzTk2jxs3tBU1ROvgeCZ+TBFnRLoFgcZGH3qta9LYinKF/MTE7TzmSc2jZDP0Kftact4
KdxCKNTC2w0V3C0b3ic8XroY3PQEUwoEawKGXlyJlIu7qAMqoPP0olmjbZNPdfj9TUjxXg92V/HI
zFh0gnqSQ0imTTW1m26Yvsib36ec0JIYMl/6wUIgXuyfiG+82ljbcuyDB3lYXGM8IAywKBgpF2hF
KUHQ+fxEXKwrkWtDctQPQCCD1ONJmUFLB0szP9973b23QuqrdeoCtJj0J1p+TQDSZ3y/u3rkLnm+
zDD9ojikWysSBbC8M4oETIdWkKhdF2OhkwelX8lsbe7HOmx5dTqg3tqvI3iZKQI85hfDg1eIQc9r
XxuwNU6ASHJEJfo38aEecWe8UsaPtn0gbNRJwf+f1l/I2L0UPdIRiGEvUXqJ+SRomuwJcZTluteS
zqZ+CwtceqXBfo1JD2M8DxLQMK2Fxeyeq1SDnMmtoqoNp/pWpOX3VhNX270Lm+C9cJxbfLJRPPSu
meMnYf5plkOe8UMcs03rVYIZh6UMUKDYs9k7B1HeFWbukvaz9A63F2+tMqFdNir36ZFrcs7b8OU4
qWm8cn1OdJRcH0sRMCwXOY8CGqXUGLWBlb5zDKb9YmzVddwKMPe49N03yRPltYT5ia0hqEiDZFAU
SVD0llpCEMUV9GXesKKp1w4dhHGNoAHI5hTO/VwbWdHFHMq0gvlf0kE9Cqp7ldO+Wj8UphRVeZox
aF/UzrG3UeYA/VGfypcmq5yurjrUqeAz/EAD5j9ZVwEOsirvhtwhny0NGkiK5bFjH+Qow0ATxxim
FFrDde7JzEHnN4oJ4WnD0JRMzeqX8+N3BQmtw9sCkvIBlAMRht9taEzv/6/P0f4OgD4hsId1lRxe
r/9Leta78y3IAKEsf5ARMKqce8nJC83zkjMtzHeBYwsRPc5Z1fe6ai1HZqiq9y88qi6daKepz8eX
92p8DBk0EuyOlwg7Mz/FWIR/7jwlugjqlR3y+IyEMVfNDFaUbSOshq/FkloZcJhIZ9XLNA0WHjY1
qEg2qhz1N6uCUWWEvGPE13kS+ABxzigQyW/NBrXIyj2vf8bhKB5M91+xn30f77O8QC2bUI8x9E51
NIhY//LddVeadKp0Zsyhpl5XSpLbapRh5Jl0YNh1ZNnFYYKyivzvEXUPP9nls200HumgQ9sGgUUz
XfKqUo7OlayFRuXDhg4pg8KPB7tCeKHSUpfw5nkUr4g/axF80fOXnjgpej/yp+gFd34xdmjf05mx
HGIwqxVa+MMYGFaisovc2pxE3cF/PuHyVGHSn6ICEhyJD0mNn8mhHW/bT5rStDPKdWPZVPkA424E
F7szrWUEQUsRAMrkD7QdJDzA9q7r+G8aeFtvSy6zMOBv5JeT5mPQDgetUYxAGjuGD6GjyfZ2SMc2
o0AAEs2xu0yBhJP7eXLe0PYTpSQdZzhNyJ3elAYNaZOdFR67Lztck6L/5DeRjyfnb8+HqcvLO596
W39RqQT5lRHfyHbTtBmColasIUFCmWNZwVq93caIKcXbeGo8gXA/OqSyWpw61mvqlLFGK3EOMOhs
ePWk5eHhVyN9LHx7svXjh3f6vP01yQsit1p5/Y5y28c4VEOWrwPB8pEWm4iFDgIOwk91t5mZtxTY
vl92mbKzjTA2GmmRMA3Yrzgyc+3E6qzc6dUrdY2YDEJxfF/r/Gw5bN18mk6uQAKTJBcs4wj7J3iR
AMcBCmIWcIVT77rB5ub8QaOvuzY2BbJ9rCEut6x6T8WaT1EgNhKIZDXe8k2oZ7c2SZ8/qfvdPKmZ
sMaqlsUCLzrtdYISc6n9Yb0JVuhELHWNm9xL9sdJIzys3xh5Rl6LbeRlZ7QrfI+crnJr3wKRdxGR
DjCWzk5P2rn9Lvaie3dU4EiAGg3suQPJnTVOT7cXvj8aMiZR6JjL/0crlKxAQLnn8EBMUbWXZ2w3
TvqkF9QxauSEJdZlGTWizAolAcg8CztsBX4LX/RjCM0+YiJGShHTrDj37DtCSphCHbz3nizhj5U9
kmrw3dtQB1Y1OWYPeenBqFkZT8OmAfMlaL9MpqjGgL5VbEQMRPYo6ZPWtgqPfO2NZrhrWWLWGcuf
JWvHje8wvfup8d0Til/QgKX4P1LQXQeYy1bnlPJVOZtZgjoxGTTwqOITwi74YCUJHTgpgPRKwuAE
GiK0f7afYOFBy+EOH6mfOiExJnaSTjdwxkr/mBwg/n0xTwS22UJb7q1/3gB1RjiVgqrMG12LzVCS
DRaaIo+GxojEYrmSI2iFDCnhepaHZSD7wj/o5K6s+9wTSxAYS7uqO+O5hZlThblmZT2r9qHkAG4T
7JkMLpXzTvs2Ul7bWmlQKZM3ifNf60kCLX3xVq2crvMLaBS3l+OoJp61baT8qEMFlc9BlREjKuDZ
pKWLtRkF1Z8lkP6romjEE7kYDXcQAEJlz8oFhOZ505TZdEazMc+s0Hzyb4eh9lb9r3u9ieHTiLMf
DjyrEhU8tYxn2aFOLPcjoPj4EkP/2L5bitXqEj/LLQNPXl1VxydNAh5OnKhJd3fnbJVX0CCgUA7W
6aXXenwxFKDz1GBVnSvNuE9OswEBKtuW90c43dbruCgQcmQ9umFSp/vbklWaxWbE5l1LUfMxXT4r
HdxZAddT5oj8ZxgSf2P0iLLIFaaF/b9mHlujYU3iIZd1K2h+p5+Da/a4+4X+ZgXMREOTEY5EZfEJ
ahEaq/iJEDoOb/ypN9vXmDJJVY6Z/r1aTGWPA2quAj2W2V8sjFblo7A1deguuPzGXxQlGiYmdoem
FVvQfU0qHx37o4mqg9HwrMP8uTdu6HPgVOm8uNDMRvCpfZxSFSWM9XbVAHhaAhP4ttBPRfUhrXlL
IyTdCTmyRP9qyiYsycs23S/dKauH2WkMBtcbO/roeo2m/SvmIaLEdbx1bzgnHB1ZShlZz0f7wCNK
qPjo6cjjM8g86mHkNI93E03cYqz98E1KnYFmoXBvSpT+MAkFrtYWzagrymNfYVOtVlgRCE0Ous/P
W+cwgCVVM4VtbkGfrVBc4ixE8EMP9VIkXwWtkpurpZC49QGMivsgc2MbtUWpSo2LHfzLP2ycu/BF
UFWGRTxZPDgdKYaR/yZhNAQXNblFj1isQXZBafajN80mc/B/PzBXZVYwSLRaNJd36nAsOu/nV/z2
3eFFKPTEmJ54dmBLhmoFffndhd5Q8pFl8gohTukr1ifs3glwvswk69NUz1tFkcpwOlw7it4pkOza
M9L335yks9s6IHkkfg2HvYcQeyB/9xStY7Nn2EJRmlcwx8utGfWVc/weKNTT6lCd6n6hOgisNfa8
SYYbGhhFR77VQKViFDUANSE2a4CMFbYJPZMH7mXu7CxmT90rZA7wAFEOqUIlWrWNYG+G65fblWef
8c2bEdRDK0ds95sBGMG+grG0tFu7suhNpDNItzdz94MmWpaHw7+WStkQ7vu+85/KnYgCZsEOiGRb
8OqWrJnclTslJc75FO2vzeyuGnhTs/vUjQMZRSlDbIn6KXX2FxYCKTLRi/pzVnuNCyUksSN4SHqG
F1V0kfu6HO94Ja216rQmZXcIcGXEdAffLbcLLXKniaH3DVz2To1k66BLbpWWUik4Ni3aAtLa7aRb
sHUTUTArqgbawizYIMaLGQ8f824ZSsJqTitwoNWiAU7/26y/rlq2i5EENN0u1N7hnYgualm1YWnx
Nog2WuvdosSAWMa4dY+qr69WitdMeYWTZcUAS/5vC7KvxQzu2B28vNU06hG9ZOUXrsCpgF9mxldN
N5w5s732Wpsw0FrQeCDzq2TRDqfGNE34Tm/bT9gqA9bZZp+DjG1z3kCbyDbNDGhZffwuNDx32MRN
dbToA29Oo7k1tyilW8k0xkbjJxJc+/6z06JU8JeEIS8Ftwk1yBT1VOOzbK5nroSls/BZVlQgn3K8
FJ8QjiG5rsHpY7oWLO0NFEmMOz5ECEQLeGfEQDdjiyWAdReqN8nqUTqhqnDnEH+0+0sla/Rypa3A
US40iAeUz9OMX7Rnh+QINf4t18dSoBVNfo8w6fhXaqlJZznvxc4tU48C06M44opEOz9Poc8Drox7
oih6NI/mw8tx31V63Adwtj9aF7fpdZ6snVBp4TaW2gATxSuOjjC5F/PDuDfbXzBDG4dXgODlwnhP
sBjyUuo2qCMwmAzbWTNLkJshFddurihiNPgI5eWDMgSBGN8SVm1rXZBCwEgvrLCOwF5mYfxYQmTj
FkJDC+Q2+2QnQ3qJ+c62egQFrjM12Xpv41yLeyeKx1YfN8ZU2iKFpktWHv2zZuUyaPG1RN5tfJnQ
ML814J9VoHyiI+30c2EblI8SG2c1OZ+VhYoMew5eF6SJ+rH4A7SWv2V0LgLeNyF9ccIewoRJLPNX
4gGUCXCB7E5JSMxUPrHLE+Dd4mKSH/xvAlg02QhfrE70hRkwhWjY+i0nKMIyvCpkNg3LYwgNWZm3
i7a00YZ4zEBsIvNW5QllkWGPEiuWtcLds1tOvjGZTkp4ifEJX/HdfLTSJx5vkQZZBg9UaL+sWvDt
FlzEqVcaSXSCBfXUQAXhiyLIXxC99sVyCFxZO52RTbD+gan2MkAiqA8ml+2mcJnK/8pqJIeVNh4r
dNppETLIG7RybR1x3u98Jlt6ibVLAbDEYiMs3NEzWxEmEPamt9mszyA2HVIYqIs3JrD3B/g5tMOk
vTRgfqEAkdR8cK4/UX828dbK8dSxiFScXKMfxWccbcj1+G7fhQL1MZl3tyudszSCDe0fdOdME0zD
2dVOkvTS8JKcebxFffgoe/PVJtjNghKMN3YVPyw7I2nJrh1ysbEd6cPzn0zS6JmJcGwAdfLv5CHq
tQS/HtHEKYkVpQFOrvDNvxe9FDrlmhwV/C4H4CgXDLo9Up+Agir4+C7GIzl9UIgdDd3QeUieoWmr
Phti8Lc96e3UtcNx+uGlIdylANbWhVThRI+ivBu9x2OXFf58Gpc2zHjmV4s1QsgANi6RQaW6IdMf
l8Fo+tlkDfuGdtmUoEosxrwr3iBJETO6bru87cJhTyPj8GiP91eSBsG6nVQFQnvsc7EmuBg/DGiZ
YkZ7sF1K8Cp8YzKtAJMu7pb+FNEdfXe7cXmIJFXikQOcH6yFNmNDE1MK62X0PS1VpR847FHD/cBH
cQvBq0nuE4J8+6EfYrAHipKr6R2GXfQl6imvfS/twS/eOOYee1zmT2c7y/nhYitv0Ju2yKM6O3hf
mIBfymI+FYGPVeU4AfMcBsLTYOV58z2sp3B4jDQEGElHFauBpRSrhULT5yeOHyZhrqjLN+mqUwZ4
LWol4O0bjq+odhQHv5/dkn3GXWp0/yjf7rHn54tl/XXwxHTR18+cHuM0Rd6cgi/dB15cdvWhP/75
Zf0A8FwXE4Jwl7kP/6hP7UTjSCZAaeXdyvamNyoWPAUUEd7oFo+jKnDNqDWFt6gS5CxlpNdiP8vk
RF66Mj2Sxv5+/bqYmsw7bMGyndqRhALUctygXhKDwwaGYpIcNodAHv8Lhq5BcRi+JCQeNAmUpmJx
nmDWpLkzaA6Ol4zjVqNuLjUS3s4kFiyu05wZSqdmVLjqqOwFwxBNzjyKA9ggT0qQmEAhC6NcB+BS
riv7othA3FUNya+u9C60Nmf4w2UsE8ebPyNX9i8CpFz41KLQ/vHDhvBSWOGUenOnq2QdivHp2EKY
gVufO3OrfhW1jAnncPlGgkKoMrDfUknDM83E6jhyihb/DP2sjxTfPm7n19gdTaKPoSk7l0PHOW16
/MvO6ds57bFZ28xUueSgMYrWOHkruxe9Lbwm4LSCD46zYlnaCs5VjfTSjlhECL03IVRFB9a0jGib
gMZfZhCSXg2bRDY47JMaIhl6fj//8HLGzGw/lE/acBb1sB/yxjXDULOAyHlcp1umSmbLBMKwOk08
dK2fzoNtrCBEYvKfJBWSJ070CUMMr7s/CKAw7mVpiTujyIb2g+PSCIMhyyeKhyqiT8XWfIZaGzXT
kIAWPalNBjpkyLIshHchRmSvY/NJIGWD5oqQJKWUEFEAVk98mFAmE/2hhCUDNgUUKzBeP0XDsjLL
OUFziWl8dIyNtV7tZe+OC8TdtgH/q0r7dJOFKoolp5pmZC2PpVp5KBI56krHA/O6xUCqhSd9N8QK
h5OkhnNoBdWlNPFCqtuIc4h3MOW0shJ8IYQUk97SVAh51R11NHqHuCtiWcBYnuQfWDHrlPDJgUrN
girG9WEuab6rnojYaEKCxTrhr5uFYyygz2uLtFUHaBPu75b3DMPqn3Pjaa5EgHpG3dEsPCUrY4yP
e9wQWwv+nK1YASC8A/liR0xQBXENfz8HVo/ShTL6DsBuyXNO4AQtJuann6pUatHvz8xDtQwAiDxx
BIXg22S6Jncm93TL7MoFYPFbI6dH+84jQdzKT2aAbD4+tzmBITFY7jq7pZ15uS//dyrzL/ITlzLq
v+GRuyeYv2U4v3O5aBdgB4zxrfOuXfZ1nG2GhWa06u5sc8OMVddaLYbiFDOkObk1GxYd7COmXSef
HmU/0TC5k5AF2joBGEt7TM7mWCfud94Tl/j1ZO/2hgyqMqKc2xk2slSSnCaXJ2UuBEoYTzS8L0V6
fOH/bbXPvUJEfsXrrbK9ZwZnlKiMYgMaWGTg5aKb4e02ub7fkaffmbGWo36Bs3rNagIw/01Y4AjD
AKvXU6q1OvjbtudppdbRXPOieXOYMltJncMIN9Pa9NssvgTAL40ZdA9QfO9m+w8qLUAZR7BoK1M4
1aOChujSjZmhsR/fSIrXLAq/NSAEdDXYuaxgn7GM8Rs7C/loMhiqSbDihroHp1HhyswI3viYtg/a
MXqbNZMdQryFHD8xrDkKPXDqcrv0I6VRx4fM2odOVZthYuGJa7QQ6wdg+2xLzUV6QgkbFbmkn3JW
sTGfHakfI0N1Nn3yLS/O9WTQR2jcXJEhOEewMBv8S0kq/+rTLUssC7igwn33b4pnF4X73tnOFiXC
ek9MWUN7he9vSRy47B05Xj5rUX697W1Z/IHwsuNptKk+/uP5Cg6NavMWiUMWejph+5dGYxlEnk9w
Ef1zo54UkFOei9Ee3mMkw6NtPIQaE+eBn7eajYQStFjYXXCvWQ1yDVkH1Y37iRm5aMgQzpvNoV0P
bqJj8mx4uIsM19KZe4t8gtS0+iAa6imQDJvVBYfI/KDI8X0gna/FQZXgZab9c+ha48piaiO4Bal/
7aJd17Cavej1QH5yQpQ37TEa4+2EmiodxVsv6qy3wV8lWhkNzJpCxhOzsrwqJJkb4xaTWvVUBfIm
mbsZ4kD78lIxjU/g5tJZ2W40ZY5b16lzQqLPZx9sqUZJ3BtolHKqM2CixAX9B+Avm1M7PEtnQbGb
7UxbAWRw07GTXtvT6TFiHUHyl2tN7+sPP1kYQzQx1VvVYARpuZPyP0upllnusHXPzGpV/nKF587g
2kTSY+p9KlFU8S+5eF+6HcY8cB8Xa5eJP7/lKz3/urafGWviKsYXJZogGLEImIm1prL8IcQq/suH
IpbqBkKvmNpPjcQ6osflpuZ3wKK2QBaVPioMxfhA/gFh60FOLV7ukTF7+s+JpbyDROjgDrTJxyXP
wDfUN1OdkACJB0o8hC6GqLpR0ev/PI6Ur998AQ94sXmBuWfd0enNEFccmqQMyJBoALS6qAuvrlb4
N44tipyHxWZ3nRuaxlFOaj32sZZXvTXk9P9gOmD0/stjYela6XvPE/U53BfIJ0XcRpG+Dt0oO1ID
t2uwO2T3cErrxrM17xNM/U7eOaSayxxJQPtQQZmCq6zBMDa4dsSWdB6XyAa6XW+EWdGAGbm8CDZb
mEI4S41oS4wVBFy5x6AK3c0ALvegLoO+E0r7s3epgqLsG+LueVgR7kK4i1n/GcMwphtSbjLGMtr4
WWfdKw/i1DU8iE4VGID6P2B0UOydPZu9nPfNR70V4eWfaKTTxAE2B6btJ955mphH8HFM6ycvByf0
Gz6KmDH7EBsLxsZtcxBaLTpg4CEk/a9kmxSm1HrLr9xthgO57HIn8vw1B49Mdx93hJV4gkcQ1Rk1
qu88BI0OQFDPA2fONfY7W60PSW2PljizeIc6MFZZPh4Q3HE4TgaeoOZHTZjodXgVmEan9k50Z9rT
PHx/Q/yxPqpPuZVpqolnTak8FnlKgZ8Jvj8H/DMQEK9yMQBQAOL5GlA8VudORxMi6FFdIhoCFc0C
dB6SFvbFiMnflu7Dx0jpxcWTUJmBoacCWvqH0d6l09GHwegJtjJwekvN02sHCSqtMbswAJHb5MpT
yI0F7Kc0RNQN7wFqlBhRhiCY0cXpDSvGzX4HtjyxYYVf7phC2IEETNW0Bz3xO793bLv6GB8NXIu8
rPIzWYZSAqsdxepBBrLcS53XsrC9u9oZx2w8dQgVguhQtJ93huiYRRpOy6JCIuyQapAqLQgsgbe8
mJMHAjAqKQSg45ZGwl/oFTGWH6AmwajAK7gGJoCumzJDKxXnN0pMgb9aLkk+xknjJLgJ6VTmLWXp
lTFw+rO7PC3oYCBz4DKkbyBYmNBdY5h8V3jn9IcWaHoOHnmv0NkjInwP1U274RJMYP3C/B9XTC+9
Evb3ZB/s2vxCko1O+BwZle1ZzDNVMMAVd8Jrwj7bhOqw5hTn5uF1iS4Ww4ACt6ZKCRoLxQmZWJgC
27IgrA0g5yCNiQGqDZE+uC2ruCQuzahw2IoxDDqGCIWKSrWoQxX2qcxBCHV2sRS6Yz7gww8dNr/b
QgGfrvUUemhq0cUeLhMQydvy+CLHW6+fyEo68t/ckERIHLLi985ohp/B7wjafPtYdvmI8+5mj4ke
kaB3D7ppdhZwYCEeI9Obq7EeyLqPT8COqn790uG4q576mYftnSs26eNBypahwmwCrp4OUXTn4f0T
5guvbitvN49SJhmOFFEOGaxtmX2Zrj7Scd8iU7hm85UOxe/5UgNX7T6403F1dfjJmI7qb2pYOjB9
oC0B6RG7x5FmAuFKx8fWypIwH0xJDwnq6LixPs5xQLvnrasmAt40NzMUhxL9si9SEK5ghdIu3oog
Oq4ZwtrxvNwshMaPM6lt94n1yhxT+T42Htcauy+83Pn/pUB/o9BUAeGb01H5/TmoXudAFIe/D4hC
uh8EBHJwWJ/tbuWXS4JhJ0trYRGapRumYUs3eFjEVRBD3npdV7zBB21ahvFKSZABHt1uhYYbg39O
RNGFBQvrrNcfn+ShBdsT3w1DF7WEX2aQ+mZD+10hq+K82pmRiZ8qkNsfH37/3Mo3RlLaMaKJfX2K
f7sjAEVfz/do/jtYh69roh40ol4FTQNI1D3xookJlxs1OKwrXh2IAvnCDi4jQ2CqeA8CKr9kNULN
FN14DAAJLhtwR4cBLcYRdRQVOSMD4xcYbCVvJa9YFQS3CdfhX25zCHVrpL9oOMobuR+lNtlS/6th
JXRJwKc6rkDPVovJtcTCSs+A9cccDnS1RFEUmrEZt+moSGm+5R/ovR18Kp9xSZJZuACU6kqqlktq
cX/TSc/hVlDpGkla3gWHnXZN2dbyur4bpRN48dnU7mhc5bKbB3g+ckol36N6bcgPsyKO2q8nVxcL
QVQ6DHLWhxa4ONf3lEOde5IXROFXqHt9rNtzfFDb0xO72kYKm71ghrbOQyjMmQIgn2qi1D0x6Zxg
WCDmSWGx4u1IXhx6pJc0OMvhx2QKWEQ9BiiQUJdOymTlqW/iosO5Z/5PtSMhf4dIozs+2fnyrPF6
LsRzlUP6uIzpdMwbYIsqnyeFg8wI9kpYyr4+m1wyUUxYpXDENKCrlK0IygbM7QKdEK5wtX9t+NGk
py4Qkq5O7bWZiRIKAIh4dUsB6MP+Pyn+ntRQU3DizMKcoGppuX/x6xW23+Duu31R50NQQItY3VFS
kOMHjzqh8002E17ly3ee26bJuuSV8SfEBGt28LQCje7kaKccwWY3vXiQmtKd4GQYPa2wpiCKF47j
8dTxmHvSkr+3Kv3F21hdV5cL6lhx1Si7YwT50SzUBmX+DBBkWts3W5YbzLihKd4Z/qT9RUF7ybWZ
Pbik9KWNz2Cjpnn3WplDaWzsvGlojkbII5/Xc275LmB6cw+fZnmZoo3lUXeM63Qq4IXF83crKzXA
rJtfUoPuBF6GxvYiPI8X3K2qJNx/M4HsWfKtPf80+A6fk8EDwNc2Y4/2qPF+56LqrVWjyoNYzcCr
93huFKg/ormb2iib7fYk654PvpK4i2NZohPls9bpFLsXlFsC9mOJp/QKTqYMtsTffKqrLicdQbq6
3Z8owP048gbSMA80qt7VxokB3la2HDEA++3W9mHsRx001tQrooQ7+sbj6aLebr5dvVwXemutntAd
hAXBOkjJ/ylf8GyyioxpRG+6aEZqaoYikGPsR1klGri0bHdNYBPkHoy20TvHc/7/+78u9vpeiR93
BbYD25x7mv+/hp/Zw+ij0FvgstfIe6NjEOefjZ+uOt0EPsE+krpEP0i+1Zr3wPpjfFGm9v67Gfer
lERyyBoSwGXReJdUB+hWx2dUoJ5ITipsrB3J/WP2aBr2ktM1CEGomm8s+o1BBzef+rsnbeXNCN3c
4Gs9/cw+T4Jo+TxcInHWg19j/+RHwAXq12yMkS6xFMmsh7yEEo+HzwSMrYiYhbkfGn7Shr62wnYs
ZSWbCsNG58FTgLbyCypbw0PVij/4nxDija2tIVMASp0OJehtxIHL40KGGNJWMo32l19n1ho46yq9
XIctcbxqYhiEuQ/QXKnBdTeNIEMaMLXaFqQ2V4pUzLAvFOhXHGYzVSuolbIKgf+AR5cJ36zzet/q
lA0GzcuwXQIEvB0MoI9pa02UxeGqhK77uwR0qV2FzqQ2C5X28l5ThwmFgZPm/rZm8mE8S4eBLc8U
esrkaDTWwJVuHoT8Ms7sizJLIDQIIfFaQR+MhAhMDH4XliFtngjcDrJhtP75CHxYrLINt4lhYIAP
ruODIcP92DgTfAtrVTFRCS8rnX5O97P4kQmF9VYxUKErdb1jF+KVDhtGH6KayuN/X73QpObZzbJL
MsSVqd5rAnxQuwTN0Qm2w1teYYrzNGFlpWDyqdmldRvIu5ZIPVv+Xh126lmufxT7TIduSs8gfyUc
3ywkYzlE0eK23J0o3pB3TkPAJNRCMCa3ktp8KWGgICGBKhPll8SKuBYRuYMQuetz4jdeVI1V9/ws
vCk6zT11ZWalSe8ag1peS63KV6JdiuxWVADAPNzdeGnfiwyl9oh915QwvI9Xiom7S+xzIyM5szbh
kfW7+/gwqqgv1DVCGQ/FJ6Ds4eWzCCGehc5RWSaEbv6o+kziqYf6k8km3g9K+HswV210ybVeoRX/
hiFMeBgfqUOJJO30BKvJN8nCv+uD5CL7XgaDj5ALbEomRt9c7WF3KDYhCVkJ/QpOChMljfUkUwe3
zG9X9SIZrWr03HhEUMQmMeMFg05Nki+QoguhywPGBk2QgOeqsPiaOE8Wupx+2cVhevFz+F+g9BSC
nNVKUiP/k9HgUQ/00i0fanqg7yMHhHyTLyGRvGXQuaPtaKTpsA/YTL+ZllzgEFYtPGxEmCFt0+KY
UNPmHS+lCC9Yd9bUAm7s+pIahen8Qk7kQhEQyh1NfXptEyUj5KGTUoszQ2tuH9HU1+81Tygmkkrr
Ipe2nuIk4vkqSVbNPzvH6iZwangEho07XeTJzwa4LFtIgye2YPLc1h4iPSopBsw72T0t/A8zS6Sk
OUWW+GmJZwWVwu/4EzjAFgnPY6bu1uBSguVAUrQh0d30fNo8mkAA2p40R2mOoiw5YyiThdF1Kox7
q1VKkpkBlJQmP1ZM+x0csAvWzEnyW6fR4ZFPtDFW14yqa9nIKXGNJ7KOb/6SM65EFBUwUc+5rcUh
U6xu6GJgDDwjDLZvjMBGH/1ixoR+TDEl0htSQtt1Byrfz+XvnDmJM+1vqkxib6EHTydrfxZkwN5D
Sr74AGX1+ts5VOtDHGN2cQrS2GiZyVPfLamQdw5zQOQ6C5vB7A/krGCuGQFXxfoXuS7F88e0TJGV
k17/B0+iKreI03zSLeUzQrHNjYDNaGjU7xGhfPwV5PjYaCS5Ym1ONnxP0JRpAPnTAyGU1kGYZp/w
5fpB140dnPO80Zh0ND4TPec89mYYfCfpgFRDuELi4I5r8j+rqtbrsipiKuZMCtP4Kyj2PILBX1/0
T6mPL0YkkcGLHYWKnM3zt2lKyE3xzXfzVblK4pRvyizeR6yEYjSzwjwS127mxcdRwyQEtUCRY606
vk2cdI+C/cMRA6bcVGjlblJcabZbyBFYQ9VEHgSgREEc6heXJO5bJGH8j61VjuJaj/spiQo5LtUt
7oLDHONa3CB85GCFnoDr8X/BvZgqX/jXbVdXWcO2X0nbi4VYffoPv0XsyXiwOQ54GiWkdl3mPw7H
zR/B4XMGVObfQT3N2ovu1Olh2lTQXCvfM1KzjXrrkI526r+2m4G+FEfD1QAgx2ZxWrCEwNdXpt9m
XQixX50vvfnB9uONVsBRp4DZ00MrrTdzDlmxhEltDOFp2+W8zbNMFg3UqetPtpRHr3KGVkMHkmYe
KLR0lmrXr7KqES69xkgeHBTMpkQLxi4dJHKWxxlSaDCT6lR3nC8BlcPgPHmCBkeE3o4GkLBDgYmr
lpuapu+P61p9wh8JW3JJG4IuX89LUEj3nnRwLZaIAet2iiW88IfEm15ppyTYvMRInVsmrNOaoZ/K
kGMIJa8QFXSWyCXiV8UwxRbsdOXUFJLvbTRHnYPbYp2eF+wmEmJT93uM+hk1OUXvf+AvAjYO/Hxz
3KaF/SB6gfEsuwqXwimcxjGW574vTEOsFI5sFK06JA3cEnBxFRfFLNWMhxfHTOYgDsC+9Av9nvRi
tvayDJdhxUn8gJRtq25Ts9eMGSjaeEs5FQKClhQ1W58NgzeqpYlbpblb6uSL0hRXOI84ik3aWGh5
tZmjo8PFujcDR5hXAc0TmfCweGUrcmZhqEzxNpKL20dsDheI2nvum9ipifpbzV2zIECz2VnxRVYD
SYi/pPh0acVSpuRk6XWR85FaQ5Gdu+BhXrXSbX7KVV25W5gPZCOMA23C1hfdIRaSHH72UE+CyC5H
ep5izSmWBJQY1PgzSZAadWWkUCaARceuwCdT6UaY6Vau8Ljgb+lpAuJVXeyM22fggfOPdAz4l+Ys
qDu/PzyYGplOtXaNR1h1OLp3Y8zusTyOkp3UFnx4W/lanl8DoLlKwb2Y6Z40oTcEoPlALeRSecvV
PBwN54PpDxVOv4GhV7mfGfROHn2vpKd0aCD2XHUrW2VVXWCW+87+Vc/17tUfwtbdYun/KXZ5Y7zA
PMLTtcsqfvrnRhllpRT0fYev4ySHxHkDKwTfCF+4Z5OgglSAQH7aRxvnHn320t7AeCHsARdCnLrm
Y6oivOzVaVo1N09Na/B+uAhgGMwpiyNjDYARu16ueFNvUxGG5KrnvIlYJLLJq726XAOV37geYOYf
MwlWoWVR8VAMqKoubVU9o8qvesa4zi1xtkVvF2VjnjFcC0++wCTGL5ANIbAtT9d6eqtVjYUtQRh6
yRpro0OCQDMCYjSLyLazNst9mpT9CZXv7dqnYvZP5ya5qRYE/3zTU4rq7DZ1Ff6JwTHxFVBel83f
RMr+tALYI826K5K9j8OdE4mo/o52KK/Q9VIklicksOZXirgaM1/paOxru+FI00LXGQVkzUpllcgi
huxgjceDelhekcPj0LPjPR1la/qh+GuJEK3yfK+//YJsTMtW1+BRx8jegbTlwAK74igKwVbhqpNT
tS7ZaXGM1QaMooRqVydXt+V/Tjn1fYtCfmsxAAt0IpqcdXmLnnuKZdWe2zq7maOIzE5UNLUAtrft
OhH/FqlIyoXfianrShAi8BJ/Y69Ws55hugHM9/9tHgRf4q/IB9x+0XrJGgzcpaCTOfloZTXp7JEz
nCYqNynNUbburerJm6YVm1Wg5n5QXcYm7V5MZYwjobuqC74OPsDD89vcvnAdhrJBZUfZR9P657uO
p6fq5XNh5FSGq0DnGsE8AJCUGn/sPF0juF47mvDROqH3QUcnbDE70QsHc/LwZGe7oux0Hl8SypD6
TLoazwgl7IC9SZ0A7to+nYvzl/5S9yUtxNVjhY7EZdbSQfeSKvt6Vy2RueQnUcmbhentVT1Dv5S8
q4o213mlrjy2F5FxiHlkFiFvUv7c+BgGOsqyJgq6iClJe5rnUVq/78ObvIJbfujLQWyxAmXjwW80
4lPd7Tj0B7/UD/R9dcy5baIxcqDEKh+ZPj+JzTpM82woIFcEQKcDzRlvwXR4ByIyh7eiNkx+p7A4
N4PTHP/ke9clKosVkLDRjyJEWbQ01yR8FSgFCMfhHPO2M4HG44nYwOaT5RYF8QqpuPtaNorY3IG1
w33AohpZdOp5mA+k8bWF7qJadYfMZ9UetT1FK2WA5+q4x3qDK6t0qVpx6G4+zFTATXy6+SCAJUKz
Te+PkklrPPlFpaLymSY5dpDoElnH+Ak7roERn+PS+CsacWVmVv+ndesWxHe5KFqKYVK80VkqNV5T
ftWalK3QzOh0pN3qGPuPEtvH4Oi+sDlw8DJJJ8PsM8K6Qa8N1ne2Sv7OehbRVwlDc71AamBMUzFO
DZiE8qol2gVM//YarCTGg+hXtJ9KOTCxZVkc71T3gw3r/buAdT273d3YpDM8pUB69QMjhQDaBLvi
QzRiDG8Pxl935HYF7POATZvfmQ1ol/mrE2VBM+k1SiKuodLJQvpZIu7OdcGWNTHfWpnfzuJ2CsFv
elJrWhdNXfkUi1po030wWF0m2aLqTt70soPH+1q2hym0/bsiCtcctu3TVno1JSKr2quRIi4F+d6d
O/sfuRw/ckfcJe/OUj4E/W5jiNeMC+oKVq9t3AA+3bjwP6l2fXF5pC1AmGZITlLXbpjcV21MfXoY
T9sY7YwW1K+4L3c/f6cZOu4xf9g2cn34kgRrG6mTbbuCMfzcPoTcwrxuhVVnQEDCRu2LJTcW6ITP
Tonm9uRrAOwf4sABqvoDFzLA3yqkUNsFSRBXvSBRT5tiYyHloaIA8XE1AhlPqOwmwsf562Ilvrgk
M/A6bd9jsld2ymqydHovhTfskuoP8+OqyU5583hf1ItEY8xjFitRxbN8rQx4JS9LNrWlTc4K9Y91
FIopRBf8MLucItxNK5Gq9e1f3ibjp+h0vkHRoo0V3iYnN7VZz8uCvTxd1acRXnNv9YJ+JHVkCXUz
nh79ityAjLJJJCJ5R9rQAfgP1SOfjiFQ0TbMMR0m8QpvAQkP8NMQABDIIQ6VK3c0DRVBj8nwI6Bf
aStgdaUChz3UFMH2sqp+tLckkh5FpSVZBos0+gG11d1wzDVPjhuv4Fxw63F022NJItfuLZDQ6m7y
TFmINPXXtnso18uy13cCUme2lTcfKNVehSQwkoUjiNNpEoaku7aYw0hL0S56kyE7rJ70kLCc8PbM
44Ly8w6OnWx6Qrp4dg64VRIL+0DVyxGt4PEoEQi2alL/GjfoNEAr3jy+fcjtzxjGsbQqhIhoG4qu
ZQ5qbF06H91yOpWiPwpE9lppZB+H1NafzZuZ++A7h+XdgJy1w/VEi6nqf8VYwR1kOHsE2e/hkjlp
rotGaAoHdX1mQWPor63QsAEvaHJFx2eZbb8mp7hVb3U2xZz8IgnZppT3/yv7klrcSKlP4VlVJSZh
QspS7rOdLCgpfUH8Ow4wmxmEMabLR5uANpGC2VPXYIqAPSMHcUqJN3lWT5dYFX7nuJPAEYiHu/FM
Q1/L2EXGcYy53Q1s/RBpQOM09z6eW4GtplsaM+2n+x55tC04w1eLWnkr+QqvhYh3fxaVr9R7EXxb
D4ZFg1G7mtd7FOW3LVe9F1CFoiWN8G7cs5k5o6qvf+KCQkZQ3TxrChlsM6AxvETBb9Ky4k6tiqZA
7JUkHg6YIpUtkyg2GcfnckZOe5EA+BkaWckkXDR2v5E6xeAdhS/jN5R/tJSqDZ8uylvMKJmQxV5k
xTZ6YkBkS9LIcbJE4YpuI991DCpMkeGRtsJeOPSfA2LmxgRKxRVKXRLHB8cypSYzP0U1T2W57Om3
aHmACgq/OF4jiYSU1ngGjCmj1Eram3m1jrz1XKGTHbgVrA2YaxD/azpG9VfHrbxXtk55TBZYjr4b
JKX+KyODxd9dM2oj4L3mAaLOQHYhn5KXZ4TXozr/CIoSDeEOtryq39SC31HX2BHaJr7/xzcYzPrx
tnNrVi/b58hayUCmUhnrsNRnsJIPmCKDHaoRdQgfIqlWFl3JavMxwKGvWhe2lqd3C7RKIpdVaA05
xjAldBg04790DMcg9D85ezhDKqMrbNHhzSfGfpXacG29b0H6AFmWKhCa+5C+mSYECO//VuD9x+v0
M0Zpbtm+E+RHjwx8/FhS6zKuSsaX+bNno6V6ttd/01jYYoh8doofpEVLl9+n4/8gqhlpdLUsDfzS
sjpKAkOBaGkq/RpwwfTSjEypN402Ng2+9w3TAX2ZZU7Hk2MS9Q19FMC5s3jhGNwJE+/pbVCdFxf2
OcpYj0ZufiNba2P2L49rwNb2vO48JtSBFTD2Renr/N1UHOVgkWgqN0U7QiWojayYknew3tG6WNZo
hnbeYbiVixw092zIcjmD6Bj73lMAg2Uxyj3rAO4GppnFxw7sFVQjHXkuA/sULoqaomsMF11Yk2zr
xkYd1DEBAkCLbB3GLK16iUvrd95FXI+CnslT1kz92gxheYdWslR2GaRoPB8FJxbyMvOCsl+VC5xe
xN8xRS/u2dZjYamPoqnmBuytreRNf7F9Gy2q9lKWzFYZR40nUujLRQxnr9VZ6xSBJcsRvty41hCb
UjzZOVWxDEIGf7ejxCJ9PmuSDClzS4CxOOkfaT+ChxyH+2tw/m90y8FDEXQp+r03ems4vlIsXGtb
fZLwhgvizfeCtrO4BQQzWAzQQJWPKkvX3Y2kQEeSqcZ8hb8gTRf2dzY9X7rCbjhaDvJC9fCeA2S+
1LcadTgZOTM2FtSuS9WpJFS84sUWUITirZAXB+yfuoX0jEk9sTgrgrW8y6GH1g3priXmBjLZZXeb
gp7Hqua5NMkIMW55DzP6m7MJi2hh8nTvEzg6tF7oXsTp8tKIYCKj2g2I1vSLf8M5BKEdp/6gvrxp
vUp8nmYWC8eihKnuQcSvd/5sg8VCQm/BgoP4d0p87VnSssNIzDCjTu6mHNM+owIOU2EIUzP4MoIJ
pwfQp1rW4kUWw/YCfAL58KhI1wwKr3fWiMxpOXgJ/XTACMMhCJ+FRDB4Z8heNBWb/obZig6/k5TX
dcGtsEzbUEe9j9mE3jC3NVT4EHj98SBq0N2J30TyyOQP3s1bFqBwjqG95n0RZLM+moeB7zA3Yaci
ZVMMfFUyOcd1Gm6FPlxhckSLxl/Vt89ZUM58FDRxJOroIVvkHn9xmuqs8q0QeRsmJNC3BBe2lING
p33qfO64sa0bvmw6um21HqiLLTERE/Pydns0pTxMEks33d3sonn2b6AjUTp54yhCpXkFwEPeRdGx
fda2ggCw6+GA5rKUUTUfv7g5HyQpprE1kTbIsOgAeTVB0XPHZNusPQ+zX/dfUt7rM1wS55EA7nmt
EcQol8m3BZx6fY3ZibcptC0HXOXaBmTKVN9vP19M4VWPhdgqNuVk4jex9NwmSSx1pJwJaCBXP/ws
vXwXVk2vhB/1RF7voMqPdBLO3ulQ46GerIJ8ZcwEEwM+uPqHjxYcTPhrzXLZFA7M7VNeW5A3paHT
TqrM5vIpQNOvr4oIN+ys7jB5NbFhY4jbHF/7Lf3ZVLj3rLDkYa4O5hpzPYznbXUuoAO+/JWkTtos
TlOb/lc5yKrItLVkDgZKQiyt5SWXxZetjfd+EqYvuXkLhiDtz0W3YHRvP8Se7ofA/rzencCvTpCe
nuRbg3w1IwWqel+dAeVbnZBU9IjXVda4v4ckzmZp6RxUfDyumyuhFTTzFHUCOcqLf6yYBccDk2wQ
HCJPNpKeVPQAFLPQbS3I6FRmssUAShMKlTjC8B1DY04kIfZtZ2mwjylRQgHMRrjmWm36SulT5A0t
5HATYFncObCtrFCPwv7r5kEnx9Z28i3PGChWEODzSSDj46MXY25joTJefuEVVWUwsCj8RkL8NHtO
ynd1wo/vUNrgdBiANifxB3iG/QKrx0JBC3g3dmMFE+jzNae1VdPdJ8LMXnsaC4FuO119vi37uuxj
RNa5heVupZq4xARrhVfL/NqmgJk5tqR36eqvgYjz0WddF7NlxW62trXMEk/kA8KKcKcjtk6/ONix
TyR1zvUV09axzTFPXGVCvjdtHuYZ2fPhJ1xQjea8ycH95pEmV6eeJnvuYTHNBKvKhoH4h7rCBQvN
vbZ9sRBuKvpiWju5QygG1dKVX2tOHQ2EAltfSlG8laEgKQhhNJ/o6AV/lO3l5pP5sJNNCcN+ojey
NXKXi7/63Bya9f/zcLzsa94EIB8VO+qpeQUwOxO05LW6v+lSE2QkLTMO1r/p27yXUE2UC8smJi2A
EuNYXnbkUZNKlrhm3LhJOyOAplcYHNn1rV0UgaiFhdN1NLKjEnCUwBDmiQ+oa/0cOpeIf/qvIKOM
x7Vh1TREQjqCyZ6ZK0ngYc5YFVGnUe6G8ktK/mk2W9UGMLGriYFbtZfRE+8aS0RjAQmarwgjANZj
80ZqqmT4yaheuWI/P4HGT4na19KXk3h0umHaxxEQhtnK9IVJw1TFNU8v9uzOud3pxD/PxQ2k+Ubm
Ub+D0/brE2ggg+G+zyp2/o7ZKt7bWGoqK24GTtcDSU08EZELoVwHeAgJzJxi6Yw6hSnMcg2fRapB
/QICc8tQrfT0HV1gB1XDvqwR+fXqweBnF7SzBCspWKSvZu7eCKlcesk0eGesl97RE33oOi/jZd/7
rmYXfo15KqQESAoN4KaQTzK8fpL1O0eFY7hpor19CBoVxf0fF5xPdDscMNSRhiqBOPChN1PZ3O1i
SeIAL/hx/AudVZcvoM4a+/V52Q0ducbqjVFHgcwUUl9PDVxNuut8wa7+OP72nT4oFbZfdpW6rrMK
tEUBhnKD3L/1yqS8PnUoRbVziOIauDBE62t/vHdCXlCHg5ALbiu9p8KHzzXogRWdErnNNukai/3c
6XVXw004bojpYuJ1SwVY2owKHZ49Yg+pg3YbQYw4tf/RiNqOS2bZ0SYUquosjEP/5tEvGcwriHMf
z5zdSCoFQIsu2lj5jHdsV9b6GdwYMLb/RAg9QMgsY+Z9thyfQXE7JmBhbYVQZBhpeemDBO6h/7aS
1nT44ejuXqutIu+o95wSGuQ+2AdEWmcfwTTBa3P+e9+Ce89uUxc4xfn62w8oYigDDvgkApaKO8gq
wk2Ysz91Z2Re4y2f1fb7yc84un41HE8xunSr8aqClXieIlMEM0M2f3JXyer8a+zb2I89vw0OrjbW
S8z25S1UsUlZ/f4vM6GiBMuAvWvzyqkEuTQFh6hlogcqzRWLMhKHmka4g8pzbPPCnsOK1B8kAC2V
LhV1uo83DZAVclDLjJn+PWNFVeJylxxN8JfV52uc0CktZrCCHpIlp4T4hLDJd/yNJPH2SKCHg+Gu
/a4ycIFTlkhwuYePKzPhJKxhxUUJ7DAgZd/2//bKQ9HdczPMsiMcW4nDoP48FLU66m3zgcNHzLxB
sohWIYKEHdQgJMYCc7z1pN5w9RcrU5MPaXCmPqXS3LmVbkCnJyrcilA0ddYkQb/75Jo73VifNsmi
ffQRrSrLij/PB5E2M9LyNkQibTn4tIKg1zRFubSVNTfOybK8+U6rQkyAQ9YdUSqgg/GCCtaY4dU5
q+j5TOADJ+d58reO8F+PuKM1RpZw1k2DfEybioAUd/19ZkllRg8vXQYdDTNh+eyGx06G1ribnwJS
nO0Ysbf697n6t2W7pLTE2ri952dMyWqR57DOoyrxG/m8Jwh3il3+SluYGFApO3aGYAIMrifO1H+g
HEkMtiHWk8WsRiWEqInAxfLtmi+KlHctY0Q+lEOEWuFH54EpPIxBjRj4MEJPiMciPxLkwKgRiKEG
ZsD7jPBdkc6y+G5g5571WI4n0iy64WXsZH8fQDL/killvzvFmdzrVOeKjq3ORhHcBr0gLnzhScAs
8y0+2c6fWHPxTy/kTVSIv6uE4sBrd2n8YXOsEgiNo33QvQkTE65IPf7OixXhXGUakxfuoKuuJHX0
eujhcRV/NuoSmVV8ggt/qJ+gkYeNm6ZWj2tbgHlfmDqgW9YKw/urMKZ/J7zY9wtN1iGo41o+t/kz
uSHtaIp5plGorzo7DoghGCqA++JeWHFfYdINoPwCJ6lPj9jhlF87LXNd81/aOn4EnF+uR91JpjH7
LNeJ81BolMAkfiu5eHuBkRmH6m7uUdlRjwsNudsVrDA9+Gs0eUFCzUYxAOMAWl2iwmxI/K1I7dW0
cn67ACN8QdLvp/Id02JcnF+tpf6GbZMz+1ElGK88XwNwK4+nxnU25mbGQnwooovB4XDN6xmNjf75
MhRWIuTJPFt4YLux1VU3UXujnrTUoT3FE3lCA4mcgGFwxysQ3N2RyJELDVoLX+nep6ssVWYr719f
Uf1jkL0ag0dFRiKJATiAU4Ev7BA5/QhM3O60NaZ+7jMJqSELIZlU8+eL7AVUqUWPEuHwCGuBWvKD
myqxR63xsGQ5Q8bqkcnKS94SYJAp82X8BAKie+7VX7F+u8i1b4WOiSnU2+1QrXXYkDrRV5KD0/Q/
ofbBocMZPpt0sXNNEdD7XwG/XUDbJSz4c52Q2OKb1P94Kx3THj8ezG7FmXp7wJ57hbXM7W5UuvPS
MHRaF2SvXERk3tjNp8ssqYJB5DZdO+vAHXN3YTJjrtGokRBIplx95I/a+ovKEfzrhrtDzhxnNUgf
odA8Rbz3J5p5CLqbKfXxX/gTO6cknplI+ogBFgvw6fuWfLnciYvKUVf0o1uypFCGDdboMSnZEMbk
h96hIVLKLP8zR7xncW3goRbEzCOKa+wFqeMsAASy8k9RYD9n7Byh1KasrSlkyHSUe5zelYHi65uq
hW3uy3gasswZJjR1sXAhlVHzi4zJHxIsGbHH5QFDRMy+tTpfADB2PxfbmsuGax/cNaAeimRB0usc
ocpXBiR94Wk+ivmrffkO0BDsr0vLGWArzGsujb9lgX1+fg0WghmVTCwp0Rn++wOv4wBGA7ur2nDo
kN4tj1ozfgPWl2uFfpE9uSzJ/6KH645xEIUtCuTfDmE/E7Sm9I61xoIJ9IVHQQ/37Qgw67y8jNRJ
BpR5UWNtaWeKaSsaKmYj7Zz/Xoj8oYxrFpQjce3GRzF0kMEDarDMQvDaaw6m1jTqGbOu1TiR9Dwi
j7sn/rNUSMd6jEZItl/sK5RY3AZRLDAkw/RZwFFyLwBP9E213D1+WkaZHIuDUmxNAJ4BRoh1lqc8
5cMsg4tTSQO+Wt8qKsHso2YbmwZe9rP4WPsXTQZvwASs/A5Cvjq5Qa4fm09ajEuKyKppibQG7PIb
0+G7cDFjOVnWo5lekLW44eyns6PehdZHo7UKtSWPQ3j8ic6hdYC2qk5km3KX1dGXtZPvuqhKDQhG
juWfgkeRM3eZ6x5hmY3tvh3cmusOym/o8R3Y/Kh53W1KVD+SyuWAmYIsYVIkbfWFidykLZFwDBbS
+YIMzWQU0TQ4RSC8NV1N8NrxZKaEkcCk6Tb10eMs7B7kw0INPOOmeSAQ0ad0f89oyPEYSjF6r31K
MgomyYAJIok3XFeUnkToGQ33bnXMdzXFYKgPWDGTTldK8cVBJSd7YinxeyggEdmHGMufOGDbNlR7
pPyLHytklwx3We6PxqzlkMceV56cvON27jfaC6BwFPIRDHfnMkkKBurF8LMOTkKiuWLQZ1GfmgG+
9JKXD2jjHfOmuOIvlZ2jqO+YXtwcRtznaxQnLrK/UZv36UxqfER/Wap+Y1lEfgyiIixG08X5ZIdn
dixupK2tpHKmX9paWiIGU1vlBMxfSUxLpx0V6ZHOe2qsXWUovSCU8uLq0nvfpGJLZhAHxMyo2ogl
2SwIGxfRip7x3fwnV3LeV2+Wu63rsG3Ln0Qnxd858qw6SZD7x+V/UjB71iKFEAtNahPmHiTbdsxc
lWs59JU07dPKDZIuZgWxwFC2/ZmXhpgYkPgMiIlEg97BrfkazV6YWESJLeDZ08c1jJNKBieT+1g4
xZoAbiM7ipNE7k+WEZRvgVc98h3EA4A1kqlrh1EkgjJEaLsc99hMU2QQhM4M7md+nI7YxJrPqvBf
FnlvoXMLPwAYEdbX+09VNaq563/iuXhsoeJy3wWiCvR1PdhYbQNSzjQB7jXuStF+Rs9qEAhkqX4y
+G3PkBqZNKr9Z03R6/tlGPuW3adH93GNSeC/9hUH7rWktZpmaKmYyBTl+yw0YuNanTp52bSzIjQQ
2OVPdKjNvWl4BXYsOPSXXa3otV+0zeQ4Pn6Cw9zcKHw21TIsWfkrv/jWqoaLeF9kA8Qcde5essIL
kT0gsPOieSugwUoyHh39+WDKa9sZFaxQDrzdehklK4rFBuyQxosI15xgqH/sqwmYLdKX9FxpmQZi
9A1EIeKQAt0h8I52rkJKSklphfhwjIxcTO6sZ2OWPG0D5StzwKr3Mqb9F5/9RQ7SjAsudpQh80RP
09OZra0rxkKazA6gYT+K3Y/kkPlX7y/L2QB9AwIGZmcwMgzHxNt4L5RJ0ApdoLCE2XsnDo/dimF8
PiHfoZGo9ltK+pp2zQwOn6Q6oroc1KR4+Ci+O6439WKcAxpyf4kyz9cvXJ2HpIpz2iOABUbFln+Y
5L5Q6r0bTh1qecYgTrL9uUIXbay6QlYNKuAkH8vZiydV1Zv/qZ0+aQc3Sa0SqnRv6NjfvNhxdySy
/tSRHNadRG/cM+8/LR/k6C/LZ7t+fctE2ndt0PMR3vQrFHwnRbMBnip5/uh/ugh7SqDGwRE/NT2y
3qnZqhOTAKHaf2JaYoPseE/0wImbpgLdGlUIBfGAccYEbnjzShYGZvAT0fgNXAgCwVgVvXy0HoUc
lXbJn0hBQKE2K1qZsOg0bY3PH/69ZB/tBGQuZ8TnW5NPYXMriYYjEUcaE5JjUBh5+MA2kY45ED0j
23JWZnUVvyIq60ZW2yISo+LORLnPG7ClCe76hqKE4cFy8+/ZG8YDLJg1oIVeYVOguqsUZ1nSGeNv
B0Ujgu1DX81Um4g4o6a7Ue1xeKLlDr4HYrdUuXosJozKrWt1kxZ8SwR8lqZ9yfMPKyVZ5K6fhkSl
p+KreEveqSza9ec8NUoQow3WL00z0PC7hhoki2mrbj4Ed6XaQLkowTKvq4yQni9rZA0hduV1+LLT
gxfrEexWV6F1z5bdeP2ClaUMb8pstihQf4F3uBYail22pO7mss22aVufzAX13P+PzNPdjqQA78R1
vN+hOskBkO7JDz9jtQwblLFkDqVdsl5niqIt/buvKBY0BBf29g4p4BChFPct9hnBOLMWW8Ly9W0O
IjcJ94yOuzvKyGWLzIqfWau/p5amUGaOsy7sz1GSyyRWzAbM90TfRxgWeRe+Borh9SWBn/AH2UIo
7h9oKnzXByuC59NeNaNhQbwB+/kgmRBWbFUGfEKUp4OiLkb03pXQtLeK6yBOUr2HeXeoO+b9WhDz
38mjZUdYrQJ3CUm4tAk2/Mj2qYazVettPOpwS7VzFNB+njJZgLOIgg3YOlc1BH7f2V9r8BXgKCNz
ZXxQUAIVwdrEQksuwo0gkWPZI+5UapR5ReS9o5UxvKFe8j/Ks33JXGcaNVxMJKYG46nMhWKqfE0A
PUxiClCv6KJ3OGgNaQX8moZFCHlkGVG3pPglDJoKd9/lusdDE9mHWn5+xLYSivc2BWknIIQ4GGgb
0//e2Esqm5xUBgMaXo93S5QatL7VF3VhM7iCT2KR85n7pJLG+kmplXfbxOwbcXGjnWwyy2w/LJP2
oXR0MqNVjKa0CrmqhHsxX09oL/Fzrnrt/8y4HPHmE7VPFCXo7eJs7RGOZqTO1w/FRr/PbKnduYuc
AuYrD2jTHouybvm9PXf/DrVBVouzUg2gX538R+s55ChzdBMlY9kyF6gbJHJlj+EVNcsOWwA3f9t2
aGPSN2r+160fmlvt4e1Dam6Ygak2A8bLdt5iEDUNikEKeweg8BD9YipmTGu1Q38t+iQgnxHK+UxT
ZZkxPKPtypOCjWi48vXDP0RqCz+v6bSgxk4yPSEdcAZ6KoC38ibxklxUjcIk9UkTKEBT0J5ZqVU4
ik88SW15EV9hq+795IFf3cTo5aGWmG4KdZOwAoVaIApjBKRnppAfbyZqtxTBr8lcwNwTUF9lckdW
0rOqKgxVO/OM1rELLMqwh6ufHmY7zrR655Z6JkF+UysKtKct8DFiDqJRSk8wsYhRPCrBTn2MwM9Z
CCCmwOyIm0WnfZ0du+YM/7h5B+R8l3ZCF+4UETiZq2Sbcjz1IjZkel/1lvIYIQpmd0HtDpXyPT1S
byEBSmwgrVovupf+/FVXh3ncp6/1qy91kangMxlV8GYNutMDW8jHwWQdqMntSQ0MZiuolul0Lwap
4+MJUV8wBodG+FA8eRF6JkoWXU2gZ1rZ1SKPYxYSq89lDVo6JIYO6RBb/kTp3UE6iduIpSZ1x37C
dZAq9OnPqlt+CycRZtUyVOg9gilsbLPZerox3sJ/TJUyQ4cYN8cgjosfRE1PZlP2guOkAv5ZXtr+
0A+EDeY/PYhzhehZMLu2ioUIHRGYyQGVozsX5us5Rn0msWwpnDNIr7W9dUL9nnC8FXWhn1iruyRR
PIpBISsHpfWhblBfhFZFr529cOQpB6kXy4g3BRKQDRjxhopKQ21uQutiQQ+py4tMGh8Sl+tQAIlm
8TGPtO8diN9P1X2KddeLNYzLI1q8sNEaaNA0lWkB9MfXw1LVxEyw0iF6L7dwoHrEZMkQFaE3YsuI
8QvpMTztbH35QX2IK4hrwi+EGqUxNvRn4glrQJAOaHagw+K2/cw5tNXncRNPs3vbUvIoh8iaJNM4
fYAAyJaJ72eK1deUZSoKqtCSnFAanlW0xVP6BnQd/RLGXdlEf4nMe61JCBQNMpuCPRWuT1LWvKuB
5myRAYP0EFoCq5/f60/i5O9w2iz0qUyOOY7padL/YbJ9DSp+2yNVCuOlt8TvQJL5JqIIbTrbv5pf
MsuuVvGofUw9BVNLxmO/6gToLMDVJ6UE5gGyavfIOKYms0ubq/iIpbzajnZXXuXyvW0cpRkVxnSF
s7Fo/a6yeC5amDcOzUG5HojLY8JUDLTSSlFnPDVzvQh4jBrrQWZQTyqsbEBDHIzZVgcCTLkMOcBh
MFMo3WeFBrf5cipQIpupWsgURfWZBZyCW4OnMEhJawlgBvH1ai4FGceMPu4QMm9DMRA7/LEi8hbk
e2fJBwg51SOMLAL58ayB+0XMHlMQJc+EenPb3M/GjjTnB4eFD2CAkmQPoNyXliId3vP8ANl7axVe
vse1mK9hdcPdZIuUGDf1vav9nFyDF95DsWcxrkhxG7hUOnVljpy1POgc6AfRPiSsHvxPTJeXIu6o
GDa4eaUcp+krnUvowSza1XjDC/Ygj41aQ1OCH4BPCZP+4+6y3B63FtI248uUXi4cP6CfVkyAFpaS
A3Y1dwj1xi4c2ih8nl1Aqbb9o5i2CJKDq84wBtd9JLNKCWHdEHe2Cv3+nwpU4mqw8eJaiSjEOLL4
n7i2KitJJUGYYyOKByuvZJLmKWdkz+5aO1uK6kQooNKBuWP6TsZDirkJko8nRZGnVoGGMfAf40Q5
F9jCH3Gd2UC9y8ayt5yWZetVKfECCYK6IngzZ2TTQZ4rgM+u6u8wCJnpDossJpCs6vnka3gytM8D
2edoRDXWUnbRJCP1jbzJoc3wbsd6ytr8Hrn/b+OjfvEl/rYPlyG4UPtZqlx2Oq68EM9KU8XuMfkF
4WgUhlc5kJMgHkPwY2SUZNmu/a15koQKjrKqpYBdIwkP2h2EGY7lKkXULMO+q/MXE7yyUD4oZleq
4D2sQtUzghAqXe/tvaL79f8cxmYULcqplm5vGocHMuqlMtyDr2xJGf040IYHhUi0pQynm0NnnOtz
kkvTmJCAUMQZBcqr2Ewx/iHedssK1cuvMxuYJyFarAUQHh0YRrVfYD6M68JoF+wO9O9Ksy1LcJAj
vt8kQZOHWBB6OuQ9GtwijjVi+FKcemTqmBryIuEzkOG7wy27Q+RFjxsP/GZZYm3vsJwniFIalPv6
jGBUb9fct0oi2+qRvwJMmJ0LkCBG4Ci7oiA4mFKq1WdCDhpKTr2GmuZGpVqEq30QsEtJAGhOq7N1
e1ZfWT/vIYhtFfE2MHesjdzRPzlg9HqUb0HyglcfpT/0NiP3ySqRm6NGxl0euBMAM4vYdytsiZ6/
qpaGlutWWVAwT4IY7ttskIXsD2B65S6A+xUSRMs1/h+AalQscHd6EmOnNZ97sJTq1QXHLzJ6P183
n+tHvzqsKOK1M6G6hErov7SZlqbHZcg3oYF7OMBEqRMAwVWSwwsDuPkSokWk3raD7dg9XJB2mqt6
onyUB13kvf6ohIKQ1m4znTiFUVbNk1wYfZsWCqO8prMt5j8DbHOfIvL+Ryt5H1wTXtHPV4x/mn9L
QrFEkwJ3yCEdnCW8A7rz7gFLyHhfjrIfCrseWwB+dagHsCTK2aEPeDZybZnTVoWdEOdq07zDbbK+
j5rrFobeGpGpoEhXuX3deY3eyGjI3e2coovY1SSjRfsIEc66B3xCBOZoe4vPtMIFciLhr/Y75DgQ
tDt5OsmkgLC27y1Cta4h6y3ilW0vQ96Y9G2F4KuiZ1q1QG1B0y4ER+zHUPgxw5910Javh0iD020l
RIipIq5RaVUrNTiR4lsFLZ8czpHWg2Eq+x04wh6lJJqs3wZxe2+tf5cMGEPTRf6nuo9jDMqsNP28
Eqvgpd1zQDptm3atO7rL/BtvrN4ZeOHquQJE8K13f/gtgQedAuyqFVYfxJ1Weuc5BFNHrNgoKcIc
m3qpG3g52mMPQ01XwCvLDjUnttJE5JDZj/y1Ig2lXyGwU+l717+HftqrXKKyd04iVgOd80A5KVvO
/0a0vXiE3PDM+943kqAy1UbA+i8XJmnMhG4iO2neUadjjo1mpg5ynhhIDpDwd7FLE6Uuw+mOYJWH
QNu0iT50ePEt3KEm0k5V2ctuBnYcaZ7tXhUw1UMHPLSjcaNfGpbGm4MgIBc3B+1xEBQHdyrwXmil
CtIbluE9CQfMl07iyC7Ps2vsKk6jhy9Y4BZpfTzxIsOoYzLPGDgFtQPUnRwOsDCA0UI5S35B61HU
uY/qyc12wngvNwC4qQatSY7zwu5EUczl3+rFKAN7F5CAvieDC1aHUU1KYWQ0XOgPU98+rnrzXMzl
uqNOrPhhR3qgYN0t3R+tiAFBa1eZqHEHeyX+CBl5HtBOV0crXklcO720alABjyRNgHDAgC0vnfoo
wkPulecIC34aM/H7umnJfyF84jR+YuLZR5oRt05DDiu1Ls430vc8cuPjSS73jE9UHH1eupfB6bxP
LGwbX4nhz/gA67EechVCMeViZYaWXb0fHwijv83r+2wwzTZCgr3/ng4bp+7/V778QTxvDCPqAgSI
1Oudc5dWF6b7t8JqMKt4487K3N8laRFM5P3+A+lXkSJJpanXTf3cREKkfTuprOo+4CxFHbB8fgT5
w0eT5GhR9zzAO+UGo12nDWddq18XunoJhBz7OAlE70UP93v0HKHUy5YV0dS6JUE0/oeS67Dlu0Lv
/JIeEoKvW4zN9kG4fe+8RLBloXlfYRHcEK35It1tpNBB5O8xgUVBtJxiFmniOZWfoiCnHi1qq2K6
gBnujyjBuwXFx9xSxMBaFiu56jk5MkFEfLM76QD++970r/GGHEB8DGaCjxBqNLHG0+XUc4++gLnm
myc9/NqXlx+JKwR0HRMachH5bPXj54xSGlBimaGsD8x5X7IvGEZAlGTzcF6CJzTVdMKrtjoawnZ+
49rqi9qblEpI6cfB9k3MhEdo8D4P69Ds6Jpt5EUP4GZDYPh9cg+nPn2uylkbFfcn/EsrQcVslXik
RegidE6o1WQ/rMuAu45MDfPtDCGVpdfWE+ti1uK4oVyr9WhseyakcDh2juJWRv487cXc4VaYEnaS
RioBfI8cS94OC4FHGEQZkSpd584wiu+MtdhWsFqNLwgsaZ0FHcaqiE/bd6ZzbI9VwqTUAALCPcGB
eJrf4nHvxCMHFFJmfd14zEE6NTHok5nd3S6kBlsH+HwrVMiVLiBdR/y1uWfzyFWfIpM7uqpQ60rX
FKu86O6bwID3nc/H+asDEuzL2Ay1M4/Dl/e6yoRSCF6u6f8oGXUYiPE4Qbx8zJ+nuhiZb10p8CwU
O0LicopZ+wR/P1PKEw5YhXyE00R6uPr8sN8ZO85hqlo9l8wnDTqde4eOAy5JJ3pq3ydZm8oSMDtY
JZQmqlOU+Ac0Roby14HwNbKkBNacn9javiitz+4fdAwKrIcgIP5pijV625iGpxCO8PopXCEzaO4W
sKjBqXhE0FZF54V/HsIkCIex2QFRJicz9i8yRAVsyeDaH/1aScUUE9VqOLNphtAXCQfxxybgV0Le
5Hxm7K+aVJRIOJq8peur/InkyIoS2R043dNmdK9+OFPI3ESEHLgFMl9lxkZnncRNaWPZTN7w4WlG
OiHOk2LGNyZXZVQcHQhcuAEPxAIlTdNXOrAu0vHA5Uc/a0lG+AI1VOdEbZcunj4QRypOA0u5ioLf
R7MYxJ2l7dlZ//zQitrTz6vVQTYOiK6y6DToKWJ0FLlR/goHmY1MBCoGAIRbNUdVJMdhh/LB0GC1
1cGo9IG8CmMVDFWFm2HwiBaUQ9Ieo0i2R9HNcsQlDouzDnMpfUO5EORvPnXNb/hoIA+F5V+ZXucs
IekXgd3nn3LKKjQDao2uBhUnK/jxHKCgmRlKdwUIRafmHHrtIiIZ7MSVJhCpBIndaxE2X4Fksp4o
QSD1FnPYK4Igt/UdNGackSiPZzsEEZA2e2khhdSulzv9W2R65Knh3AmJZooPYcjBKowK9xSi5Pt0
xS/YvjIn3F+YKkqPYT7jEalSXMFavsACT9bxm2E3x41HbtNk7B7A8rD3inHeqJhABZzWzi62gIs+
fnQC8iwb5ZQjsJo/66Iuf/bXpmBqZAZJee5Cf3GoqTsxpmN6pvYQSN/KMJM9QL9T5K0af/QR3MAR
Sb8mcVZmzEiXCyIqmuIbh7MspNB0UDOu+MFB7yryy3ivibYPuRS6vnA0sb74RWd4ZZl4qgJnQvW8
d5+5O+6ovGM6QeT6aIABx1f04xYvupsD6xKcHyFo2g5sQSajRi0pURAj3zL+5tQQ8Qub5HQ3Rt8R
QZnCT87uqXJ8fRk7xyfdJrHjtEVx5kRieyeEKIbtgwM9j8PoEe63QC74JReXn0r/A01eBr86UcHy
K8bePDFRdmsZVlB1cNyRtIA3/JCZhk/S346YXLzI2VtvIHghdv0uLaAsOYJAMrKFDx2QBVt1SNvW
ASt5wtjMUa2jNT8LA72d2QcFyTKU7BcJAm5EcpivmbkXYXM1nBD9jwlQ20j2HwsyVOfl99MSVq4k
bVuELoYVk98Z+jXG75Clcjv2vtQk0w31cf5GP1Hvce5tL+PP6sBwhKXsk2c4mVL25GiQEeBJKH+T
/PyoPcJBGJfJNJH3E5nzmDV9WxHIBAsEqT/lSSIDl4996T7GUyvzGBGA96mnXHuyzMfkOgcr2Bje
G0ark5raBHNYT83SmfHseizrjpK35FLelR6OC9ZmlEow7Ms+EtKZ/DSDwBNt+AMrq0cwqdhwOKwK
Damr6LZpUAj/wjg9OLjSg/pkG6m+tbs6Dn5PwB2zUrfX2fD1241ISBCru+4eDEzaf3NhYNY/5xX5
VCh6GQMpnW1wBfIrv1tcsRv6yoaRJUgZLF1uoCHgRg5SiBzqXIl3JHXmwzoS1SyatStKwXVunh8r
TOts5YQ7ColCtG1sU2IDy5CErKAKtydt4GCmyN1Ac9nrU+oTFaSzGCf+0T3fDt4s77+lomxUQNhg
AXJnBsh6SafK5/CTMtory7KDMrFLvZJyJMJrJvc8Ftw4lXcrrtAWgOj3pJTgXpmhjMDUnT69XD2X
HUlOZ2pQI2r/PLTiEdILhZJHfStKyNgCknVX9Fskda0t4dwVZ5qVqjoGqesPATbPm1bKl/TeesTJ
xd2S9dZ+sonZjAkZO370ND1Mu9+csb0XAnCJegkWC3suomAyQyHl3q86YpPTJOInCGezsNoVZD7D
OM3rkNnPqLnoHMTZbuWbZcVMs9PaQLOvhXUJB6HMWA/FSprBmK06DdKRJS2xQYztFcCW/S/MYKub
v7BNp0ul6Lzc7MdTelhAILlpOg2JqcV3UNX4m7iXPvJuLU+OPuaKBGqxNaVU84EQ1VeH/5E05I4y
pb5pHVXlAFt0Ov9nSdgWvPEtVRVVGs7qoLaB5WQMoBsn5zSDPwZtewPYb7VgxOhdX39rQQihnajH
zguiv3ROwLjgsEfRGzo9ds+QxLwttihn2rzxuQUsPMwGVEM4trfVa+4dmkB9Go88ykWroUgdBtDZ
JmameByWK0tFPgjQr52xDDnZXeNeBoos5qljqS2wvBVUFTTc1dHSHzSVQBsJFRxs0KT3IdK3OjWC
8grHuYvML7lyZHlz0wmVE4yepVvw7J+yQwfB3RQnVd0xCSTSXTga/p48+y7s848ezV3RphfWvDkc
aEWs0df4FHbyszLwfUODXP3+DhGMQGvlEdPvua9eNj9AxfXamfGUoBrdhsEYSiZXkx1I9J5wwWMM
h9TVUqD3DaHpyaSQfoLKl5cjQ8wYdGxexx6rb55EC61Fz4IeWsU/DxVPGrWF8LLrrNtAtHh6eYiS
+hb5gGZl2hXt9apN/7HqEcN78aB8T651eB6vUxVVI+kjZxVfIFRYtUgrKNeqlNmYGTLfN06AO/0g
xFitNENO1XG50JrWCX4ZYTFL4ZUIHTkK4Nm7AuuY16a4HmeeOC0xw80TRK3ck4oRSGEvdK92tFN3
Rj91j8jHQuq1j9317J1+tLyZ+N2avf/ZKcbvN20lN/VD+fElCwT8Zdirt936qb0fEM+648iXp3Zm
1xgwPVBWLrnMEQODkkshUNypguth/LB5NaJbF9GiVMuMUPvSu7i/aMb0C+5PKGLH9VY7otSCpau6
h1lsmnAEDuWYPcvI7oOu5IwGibL5nx/NXPkh4xlzYCMGr2IsFraVjkCQCo9JkPcNGXngrV02Q0ss
d7dnulRIdzIbn+xmpPofowlZpNCYZ0T87FuPDHsX3ycNDn0e4YuaF4GTkS9BkjszhnCqQoLaJepG
cf2HHn80kbOCtR4YnayENz9SP9EpHIymdOY7Z2V4BkUjGfqyuXS7TLxUfFQEer1pPfBx3dwvNNS+
yXkUo0fmAPrNlykK9WzJ6zY02+97qOLkR3KM1ZGX8lGOv9D4/9GnOFJqyJuLSp8HuKsod3EdbkAi
AxB4//DFt7ohm5eZ8O1lpnzlA/fB9K0j5f/F/SVoBp4Y9W7tIE9yhrD40XJukYgMHA1gPfCKmJQ+
8OOTx0WvGBRHQo04ukk/b1JP09sOOORAQP21ftFfPgufTWoKUgR2pg4clR1EXHT+/PpIFzFmmq3B
BGeqO4DmyUXzwTy8VjlbsEJXi2/yhRshXaRQZSQRa3F2DqzyiM+DlXpNBRXn2Xb2A2qaXD2UMkmV
ehvAPHgGyJyqzDYyLMm77s12cnpKEkrbY4iD71i5ptsnMmd+Sldc0FRNsLRw8JAX6YAflnX5FBI+
fAMPp2aAzca8og6GyaExyXIfT9v5EFD6BokfcxS8mKMWbhuL5E9bfCkL/b53WGn1kRo9kULNBnvQ
l8zXMbK0jTCBjbHrZYTdAprbEF/YRgFK0WT6nVf7VOEbAWfaehNNdVx0plkWhJwDEzZDcYnU9EAf
UcsE4qUQ7Aoh56wfdbgdjBUAEmVhedKjz/ERrv/ZbR+trh7rV6A34fv5pUncY6gpD9r+IdiNtTGT
SOo28Juyu6TQqQV4Hg22YY1vpfdKkxregF5FdXsW0NXGl1BF2WKLdmKUdXY5DWopATrPvLRoEe7d
EvpRzkfkeTIhRGJuAwf2vgQ+gdslMvG90GDiC31cZZUrL8W00mQS4idJA3WvAfjlAmaZnYr5vh1d
0PbyKJQ2CPbMYrHX8QcdSjfLKjS0I47Xrcvp7/HDE7ucrHALf0ThxrnvTjtFMHQbuKm8FEbYWxp8
abpRI5cZnaPbVF3oL5FU9uIQTdqflhx46eFC+IwU/OqRnZhQ/sRco1v47z9fEyPHrDuu7DtRS42J
zYR5rm2m//ndtab3kipr9ORJmTikBohUQ4RaASkvKXXMpDPdgmmU4IpX4e/aoHuvNe5F56ZYVs19
icnqo5Rgfp+yt5kInSZOBt38zlJhAT7taCOaWt4ySPFOuVKrRUVgOf9K1myaxyA032HQrWRsb7Or
SWRPu6nXSGffrM1WeMyquLemtHJO51LCQU+9dbb8HJWGcaapMKC60aQNenZK78CRmmqq856HmRx5
Sz3TYe2yv1Zmbt4PlxHgTATNvkCzy183/g+0MQ8ecoyQcoY0VLCmbLzLvfXDK5/LBjHYvqqANYxQ
tdrm1GwRsUYCtGxPdodynCmDnj+x8PTjiKInOJlY9jUXtCb55tas8TUn3QaVEil8bSio52ksA748
kyOB2GWFRaePDRF9C2T76NwliqTiWYSGiOgCsNSosxZI+7TnqhB8QQU8UheMi3gdU4bTtJdPXIWi
PAS9gvvh+3hh3NkCcLJPMu4G0EF8MFDW+F6BX40WgMrCcPsnB3c69lpQ1i9w2t6K98hqzWfZuvLv
t57hy+50fDqVitrj4nQmKW/dEktT7pj4IamL8kVmsngpTLBuClCGtQavjWoAJeLARSA/ZU51RheY
5K2+cg62XGEGdXl7n06mUSaK9w3B6EbJ4tt7lq87b7Wvg8weAmldkpKGK61uJEggbefxlrwMD60H
NNWyql7OAy4gWcdGjLg+Jo2nydmURMMHF5WhCsZla7yvCka3iKF9aU3dxyadVyaL1F9eL53vMk+t
/dpd5JatSqotHoc8Ru8+MSZVQ9KuZqpGH7Z2rnn8vOFyOlRdusoHCS8BkA0RDHYbc6dTz3WDhDZq
sooSb7cG7kkIMQ9cbqj1t4ZuB0jSqJ0kdrzo4AM1kvfCa2kLkb3Ga59whOXYApIjQAG9PdkmSSin
GG+sxYfKT7nztzdLz/h7Y57kFqhbcVjLohnnVqY2vfuvwM3hR3gbZIHKtLYcqjMkrnu6Uz9zcvwE
gOjMt4Q2GiVGQoExX8whWyWBYjdeXXL0ApUzr9lo0f9ALWTv7l/Cg4HxUgSUspqtuRVKAOlvh6A1
+gxQqLLa/dDygB+qGpDzM8P3fMmbAo9X+2FkWeC0BlTyqYKZJunvNfPdmUGtrU9P6lHPc4AA6joh
mXlhCLeWYfKHAgxD5kZAAEMRv8AKeqRrJzaZm+8bzL1cjfgio3h6e7WJ+zF5QnCv+Gh0ih1z3maO
VpiUMzLhdmb0u8AfupLLmYivR/kiFwN2vNCK6/U3VL9D/yaLFLnEyCuTUo6RjGWn3Jha06Q/jzEQ
x7j/IOI1l1uZGqOUje0FwQKLFlQjNrU8bUiAFCKfmEUSfiujOU6zNVCjicAgTbACdctIYPvvjSEQ
WI1zR0eVJ8AhEIdn1n4MTB3Iu7V50fUfAKTJOQOgkreDED52sR9uXqA39t2remkWfI99uYAXKxku
8KcvppbJcu6XvAo1O4egOQ6trQ8WcUuIHrJiFdAfOSwr4bH/U2z6gRs8zaQuJbbMr/WlGGA3aA+D
hOKuNR4u0Nt/5dRy+PRj9PxXUc5CncsXXynP5RkdAI4jhamn/B0HLHCXEaYgzun7r1Z+7wNoutwm
F7cC/TdzlQKOPSELxkiurQkZr7xMFiJg+3QGYcYhlchOnCnM51ODa+d2LJ2k62rcSSS0czyxbzul
oh5hVSdk4cR4bDMG18jN/MIOwd7s14dOQuiQd910RQq6DJ9IJhijg6br4TqOk2pfdP1Gzh3ZiWBP
hBPmulKVTxyop8VWLXoMm8JkydHotaJxuW9/cHuil7tbHr7iK9aawd4YQL41aYf4xkjC5oJOgkZl
/h8X8743UbhwHyR/fGUM3ezMJfB0rE89MrU3fK9yfJfnSzu22HYxjnMeZepuuyEMVjViEXJO/9y6
3hBD9GWZE1kIKjbM61SWW40Hk9g0IGKVoRY8eWwjCMuONZYvPtUV+T2nFg1TndT038lysLwPBy/+
AXZ0rog0QNkcvgF2ygl2BWdxqxhz63eSFd44ryYCV8Zh+90s1bXHff5ixVYEO08WjDGNljFX5BdG
Bnfygk8xdi8Rg09S1Hi+zM4HhdMPANjh5GeArDyLLZjubU7K7dj5QBuZkK4iegbSQpbme5/o1BDH
BLhLSbQzlcVBI+LKqCv9RAUm+N8UHq5IjlV09JZas2j0gORZH+AwUmvdXyUx+1LJtyLcGHN8zGqI
POCtAV3f1WjghlA6cJYrKiY4FRACd0+Cs/0piMPWV1SCHpx9eIB2zAF/h6jkO6bDpUhC+dnxWNVq
5mmHST6Qk//St2Kx8uY7xyPdjiqu52u/6aVeb4I8OL0Gy0WlVZWCWivPDq+Cfwi5EuUfDjehkFse
ljnCMr9RlvFVfOO6Df3/iW1M8yGt3v4oY7So9buxiCTVAhZDpSSSdm1d7VPle8OY5bTypMd+YzZP
L++qHS+6jcNzg+bM3rS53jHK7VLxpdpbUvdVz8gl6KLl8/YBX6B1iPE6Y7cGHGBBD/T6Phmk71bE
ikK3hL6mKWYeaCTXriXpfJAtMJPNptn9kOJQPvYXLPMhqaInG0mmM9L5yBV4r3omVfZBI5ByWgjd
QYODRhgX98zkdZMAlq0IElRIn9lvPoBwU4rnZLs8WtS049gxZ7i6aCUV9vUdKK2K0Fn5iAnByjeV
GIqKiP+QbXfTapZjtrLw8lJrHVjz4Lt8E4Qqrdd8UyQTtVpRWXLnEuFK+ev9a4T5r8thX2PJEwEX
1OH08OEifxeoDbEmwx2ksg2Db4T2EApoCGotAHfaXJMlCIPZWaSi/EHQvknqCqtk57suAkPCQ7WN
uUZuK74l9ca/B8xkERY8bDgklVcOdRfm6tqGkR3iwROZUuOkK/LGBIB4nJ1C1xeZq9LYZPxGDv+P
vI5ji1nchPEx0DbrqF5ij0/saq4e6O7deG0cUygKl+Z1WGV9M+RR6j4zsLBewsAV4+fa95OY40CC
z/AbuUTh6KTAWvhPmRWjlOMTkgojtMOjt6RywpOuKwG9jJfOiXBLJQmqMyf38W74X3CqYZHFy9Ab
4YEsc8N1R1AxL25H1Z+E5tjlOtA7a4gShXwq390w0gMS07WVI10h3MuBuhrxvWuldbAUpDQeqpkx
IgMRhhOyJXQrDUeuBkq/b1ntjK5wISPHOcMqgdzaVO0TA0gLln5jmy3Jko8ztSGvS/ECQxuyDG7n
c8psixvz1DB6BIBcmdbBoSQwbbqNmTME5y3KQwoN/ZlOO5rmULHRc2XbNRY6V+2zHW44eKf6Utwm
AJkwst0qGo7ic/obVWyxOvAR/0gG3U5Q68x3eG29lquGVEBlHVmrBx90OFGmCoSP5vcZrBuw+kUR
wNzLC4v6IvaSuby5ZBdvubFdnkddIz9KNPxez9u7xfMNXC7SQAP4r2QIaF46fJROYg53iMZ4fSEY
+uJKpCV1da0uML5MqTMnWnAqjEgOQNBXq05731y3GgwEO7dHih2Er/VE1Xe1d+FFwGIBsMTg0Cvo
ZQBm65Ic9Pn2yc5SvoEAIKbipWZMTNlfMQPCvYjk+y67izMHaHx1eDZx2DrSdksnIBc1Z+kd/MFg
mnjxquq3142XRuFndCFIJnVv3sgTAUzINdA7mUQknyn7rrdxcYQWyFC2eGM+5TQlMGX1g4NEAWoD
F9tuUBxrd/BMBvwQyKnU++hOhSyPgNihoZec1Jg60uhL59kXPbI8F5jQZVULPs9VykuE1tVIxjd7
KhlwPCEcdNwlNwvykTktcjVUlo30/IUl8KgJPBBdCq/SUZB7dHo6UeMzTHbeq3d9bIJcmwLmI6QM
rasSUxCHKPqXGOzo2asaEAUmXLFF2j9YZAvDlesVkFMjukwa+aH8cBXHUzabjSDyVFgeyTlsR8gk
fABVXgq1qrQGM+Vj5oeRPUtPtsaNxGBSrxlIgnxq9uo3lwtK23q/qDyhBle/lY1SSLdex5D9gd8s
h3VcxbLG2Nh4QXkZOh0rIXssk4d4WI27x39vlQmZcRKbI1T38XWyOedHvc7h3C3cFVs2A0sNftOL
d924Nw1dBoNxU1m7hRQdmkJ/7Guhhvu+WiJnAqQ+ZBDsqUsw0/XGyDR2duO33afU5J7yYMeJkhGs
V8vy5ddge7MrT+mvJybu4fAUhbLuwuvXWJrGsQuCfHLgLyK+E7WzU1ERlmOxdi3XeYhoBZb98UC8
MnY0B6qIWXUAAeU7w38LBG2ksZuA5k/dS3faivO2O6WeZdw9HByvvjeUnMiGh99LQyAUpvsO9/I4
KRP4Hx9TAsKWPLGjuv823OyP7ngV8eK4IMD+4dSssbLIZfX/ecXRVlrgmgCs2bZNTRCO6mUxVP9O
aC4edPIwF+5cshprXxVlIpTmw8av4jIpEpwwlMKE1GfSq0IUjFb8Ch6TWVwd3mnpZ29NtaVnj+pq
co2p2yysqhv7REPESIoxigkn6+qDvRRK6+TOm1Kl7NyzZYC2KAvjZLqe82MnkJre7jChotXD9nWA
HoVP1QueiuiRLF62f/NDLYeL5YPQqVpy+4/fwSyhWGH5o1qlXAIyrFZp+h6UXs0Y7QN/Viqg2UWV
lVnPAFjf0D6y7ftfCkSryl+O0zjm54/MCY+OHy6ZvX84b4IHOuojlJC2DFMZBQ9oDQxzMuNPRsNB
jDvKnxuzK2jN7PXl7NvnrUtlb8HFfDtdcUmNTCSAQSZ84rBHnotDP381VYXdc9Pyt1ATNUZyB369
h+gVpO/ouW32RsUweUbfqF6DTfrtchyzQJDTHpHUvXVmjtAyi/KTJfoHjK07eR5Oc3svx/by2WYP
FIcAnCIg01Vk1v5BjZ/IObutlBkVxhI8crYVn3fTig6sUxWvKOHHpRZfD8Y8XErdhrh5ls6YBvUL
J3VUZ69aW6t3+52zKBp7CcZWaS53qeGOauWIDdHTmBEbkITQIekjLTru6yBCiBNd+s83je+402g+
lwG5VEjPgOiW7af6/pFbKBkjKGLL2rk7lLVDOET40J5WrAAOA3C5qYkAjZ6JMHRIfDx8BsHzoux4
IX4bWD3PZHeuKxe0MNC0pRwcnT2x3+4n7sOlYAqa6eWXdxoUNuEUNJWV6SsoDwC2aqW+VoN4YRn0
H96NX7PvwA+OMGhNSfmJqisdDADT2/2MmdOYQf6lRkeZMLfNViSZi0rtcGzykLNjda6WZdwx/I8G
2pTjcIB5Vnsgh1d+P9ounIqSyv6T3ubAbaXy2h9cABaPsfhZbONPe3ENwHqmaZ6wFhsC7vaf/CBH
lQymgwBtSBVe06CE/E6IUdWv4ZM+0cjusJYsxx8C0XApWL0XP2S7DLyV2iBULGl/yUCTCkRILrNG
ZApv4fxGIFA9UY6FKsNXYcVFvR6f1GAb8x7HrUCIJxw/82+YkzC2pwv7JaVK3AnyQ9x+fgcHdoIS
1DPmJcAWa2mnhkBH0C+HboDCU8Kb0R01FSzX/SusK5Hvbs3uoE8RX2PCzXy6zZiT95e71kSo0cNO
AMnMdCxebSyKpUfkGnHfELopwYlKdg9ff8iwuFrXhosq/qvuyy3eMzMMy74nY+mrM3svt2IuRvc6
T0eFEbnKBNaLqEGS5LYVyzN8qFW6HU2E8T473lMUcch484uA/BRacKanuFHmmC5jYv1eU3IFw93A
57t16fUUpdjh4IERrMuLPnMn/bUZbs926MYPjckklSFgygjql5mgu4kzuLHX485Fqop6F89sn/NI
PNTWx4UI7rA3GRMDOZ4Aa4ZMksuQa5VoIiM7Tj4o0R5GRywvftq1A8dmNaRarTtd2ljmQIR4yuXu
m3bxtzlSLAtIVKoe19hntfCOK409h0CtjpIRheL+2GXxR9UpyOhgVXX4ft6GzEUtT+XePB9Tv0jb
etvOjfelHEP7dlaPwTjZeP8XsY92IjFKMQ3My0/oJQNfI4aS9CCfOaUi4VrFtOeqAunBRCepCsgA
THhkyqaMeivKI0Zv5/Tc1dbwaNkreDnxlIOUQsL7SNswy9wsODiJ5JWpU/03fv7PXAEo/E/fjuhq
NrX9x9QGUjXzDZgp7rbaz3xKLm21ZsoVySTDH4bYQLpXaPsxcN6r4865y70xHenIZGaM5OKOBxOp
uW05woMMEL6Yoe3+KfMPzxOtorJ4RSjWpHrtBmCgSFfQ/FbkYXvsY1kQobb28FqppfD8cu3m80Av
EDR2pmTKhcP3mEY6JXhnGvcdj2e83vUJIZHf96ZjjLPGcyAyOWbFQDicUZH+TK7nZOHYa9pRQIO9
BZJ9l7O2BwXX+2K/R/8hMzFwytg/7mjJqiPpXjCS+XzSeuAx/ZYeUFxWfynTe0uHPXaZk0Q8iqvU
ZbUNKyNZ//B6qLYl/lqdLDDbpa/hQIc5nY9v40wbmvJdWqmQ+Zi94jc0v9eOGgLt6VK8KsDqiH0F
0nndRkM9HiqohEzC22CXxZAEDks/er441pKkPMeGxX+mG0QJl1smia/3+qgHtM0SzzXaMbi5+vEz
dwjwxUKddM7WJ1uY4rLStKwIus6Bb0sr8ehv1E6mnhp5ekQOLxaAjY0o7456rHE5BQFan/s4oVmf
nMBg/ZkxgFJKR99Fi0XInXMn835jX6VbysK3E4XHE2s/NrlYg/yT9qc2T1SACAFRC3NE4gMc1faM
LserL40hYnIFSTcoTtWY/ZGiMbiNV5r8Se7XDrCGWPGpx2I8atrB2P+mE6lT9RtwbSeP7+CwUEPc
n80cIUV+j7fZ43t20f6OPxiQ6kojasvrit8FzspTdHSMNbAC/L4y7LYBqUQs9Sn9DKgnScOMveso
5gRlq6drVvBQbPt4EbYsW0EiOi7jXpI1nfmXcU+Z+eC90AoLDeksDTCW+iZuvG+IahA2bahZdMiP
K3J7VtGqLK9PkF8UXMdgJ0lGdeMqT9a/hezl4G/2auTd+k/Wm80/lTQftiMS8l8l/A5LH3UWpwJt
JlOtkU4yLYVbUBn9f5yzLS+sV42qWlrgKm5XB9cutuSYniDKZrV7ZtKavxCF1noTly1YBLQ9JmUh
Zp11WpA0pNpCDLVCFpNO+K7FUv5VHXVdyhBF+AET0bNEuXd7tqmUk69SFbIQjLQu7yn9TcC9+gfl
icSNTggWI1DXJgv+aYqkjZh//hbtf6jCapjPrrdXwI37G9yQcI3UbSEL6HUX3vjmuVbjfg9TrbjY
0GBel5ep0f6JvvfvjKoLYXyClNB2R5mByDpXLul7wIUmaIqUpCz3G1rVN2ZU9zjguFa7qQ6iW2qH
US0JVR3BlXf3/N234d86QGC1e0VaRe78wymEQRFWGmc07vo17Vr3kPTxP6OJZ//gChhvaGWuACEV
WocJqxSKYZvDgbctuRDZB66K7gQ/gVUJNyOb4sjiruBaDr6b9GF0yfjlPcmxSEmDIIhJw2f18Db3
U1UuB3co6LwEpLGX18PUgjghWE3j8n7FPbW2wtx8KRizXWpGCjGLO84eJylNun96irLoBZkURSJH
LNXULYjcYxk5Z8Xi2qj9dIVd8prQuor7JS1oHmUrRTY3R1jVLYqmMEwmL9eYvd6J7r/7QLaAasDa
+mv34osjEC+8PJpiB5iV1+LRgtYuicK7JfGjBNGzkT1c9pugxw0+v2dYFjT2TtMkbCZjJfNEaDzJ
KZIaxCqZDuVAfyGhYwlmneNntDuIQcC6thJQwvB2JHzrWxFVl90zesjqJPMoUdl06oXRc8FoCV2o
qBccYtGEtfA766wNb00hINFxvs4tY1GurssA+wu63riGmEvVPwVIidkYjuktkaOgMUUU/fFHvAm/
F6zjnPgy0+2ULxAtyNP5cnEkiCl8sUDV023+liTgOkTCtvyrQojojRDp5jH2Ee/TXsz96Fd/UW5T
KpSyAATF5K1iZR5gnJAru3BA2awl9T34HZ6+3M49SFsLsP/C30YvN3bBBHuBh46dw9PIUHCcHahY
TKeyECNn8kbTtjV28g08eP8bTaWmrOMQWuslIgXZOxa3mxG7NikhQ1U37r4mPCOXuE8YfnTOHom5
F5FxCn7mB7ZTh4vN6Pd9FuUTp3H1WDGjYuHXGOK8eGQybgOS9JiEDIl6cuu+kOuIJs8gVNjUtCAV
lw6U/CRyu4OCt24GJQlxwF9TgDtvyKbtEunidYFCjBodLGeomAly2yxysOsLM7Ho3STykVXDLp3J
DqsDJV8z0fzCJLUGirm/tsZuXt1ur/VR3zNCXh30PPUUAsRKAgEmn/2HRde77IGws84QmJlpj26D
92gNp0BVjZXb3KaS+KkdPpI0DDJm7Yq9KoMqDKEw77TJsSytobcCw5QZC1BqCpqJDmsfppz+1dp1
sH4oIhVFdLCKOIzrH2h2EB02U0jIUHsi39aMg+BUJD2ZLn2nk3+Ep0sgeyBPFO5RGzbb0cy+civB
jQ3uSYjNxBOJLZ7XN9AwCJaeSwr5zhFZYuRhs+eaAPUrPqoL10/IKGKeVUiPz6yinkfAC83G+/lV
VTytLsydf2yNH4fGb+dzYld7lgv72qXjli5exxY2A7RYCoczr0+1xMydXUZTR/CxhRr2BPQR9iat
B1YI97f09Z9GRmZ3numEZUU/ywjlJWVcZDIZ0mXer0BsJO0AHEfew1wm4dbtnJ/77O/6RKmSsv6S
MLpG+S6SuSwpYgJniCVzHm+T8pPypYokLjEUwrYVM8+IIimT2Hs8lGsGqtlfjGPULPIQ5kYnk/8T
jXpYABg4NI6Lknbpqvzevq6TE1MOnAQJ/rL99projmjdb+ipdXr4LHzsR3y86TQpiBEhv8XSE2RN
58zq+TCcD+eAaz/9SbMPM2Me30ONF0UdgFX+ix5hAPUX+u0vBFqkJn2MDLJETsPoYtbUwHlfdeBs
q6CtsUXkrhCB03c9078/2pjVJBYnKthAv3/ZOSDO7pGxj3YE2/QgqtUXv/3yCL/4MPmZYkuHNoSI
qpe6r+OIqm/00Eub+SjPq4vIPFB0HhhcOU1l6CxEWY9jI67asQBVEvo8MA06kHy5Kwg3vlCcct4e
qxGOcpYM0HsVHhGx5UFVMynoAt10KO8TpWrfl+y5sQwlKhICuSxBxOLiaeOmvEc07uj2Dp41rH75
jHy8H8yn653HJARy5nzqj3Lhu3Qur/PBFknA6+dymb5Ym/uoYC/qQrzTPz4v2tIAsEpJgQs8Xgoa
Q3JP74sBy41VK+NQJxhwxLpQiteRsAt6L+OKJdx+edKhgdffDunxuS7i0MqjiqeDVDmC/lbxk3HL
BIAAWfGWSMEhR6fIVwCHXGPsIibn5/hInzl3NAWAK26Ias9BJoRP0dsD5vdVrnY+Z3I6iGF1jxPj
Pn2IX6QIAOfJ09pFFi2XH+89aSBwONcnqmnTb/j7tS3JJdJ3Sqzpof0sLpoELJc648eC02PSJRXN
pefRUB9zM3XX98pyEGjfF4oQjmweYPBtVn3b2NkC2btg+E8FYSXidq801MSBzTuGXiJML9Q8VUUn
8hWisdJP2iHQA4GiCSmR+p9/9ByVr6ggGzRX8lmJO2CX1cTJ9P0XGaLGrAInG1ENrdTma8fvK0oD
jy5u78a5jNK8obWwUNsHe/MIjsAM6htGfxGe8U+pSim+V2LlzcqPKll9zMdu42pFPdyxV+Ap+kbi
6y9lRKDg+JMdfm4VxVRPZoLCNgubbNA/RuplFuTjgYnTldo5nRdoWeHTJzRvyLsZ5aXZWnAql8m6
sCvMl5zEqUHx3j/kfMhHF3VeN6i+dm0MaHmaLTjCJkO64t/SLXINqJ52nIA9bkdg40SMQFjEvZYU
o1GRJXhmIWaqEWadglz4VElh0ilMjZ0tQkoj0NB7ozMocdQA7V3fnm8bLizmgW2ah3WI+8IHGHhN
G4xPoLRXI7Aj7muRJN/LhsuydYAna+sC6mQpEv8bgIOhvHLUKB1WOqPnD2C28XyYgM9kpzlJJNHE
+y0hsbIZf22k4J4C8OmAuWNDJXfwyw0f6oMoJv0tr8mZD+Gb3bwcDqqG9W+/J/xeObvLb5y3nv9f
t1CXwfQgeDiNz7GL7LUxytc//h6bdB9GvnbGp3uYALwESkh1uDXGXquOnhQ0kaRi9USk/eGgw62a
1KLPiwq70TEZVK+1cnIfTdDFRv1pREHdgCcjZ285Wtavu37SkH4hMtyLGltHORj4G60J3LgTgZC0
QEdQ+JQRtBJtqqcDdE6Rpz7UG0RLSMpSNjtFoHH5BB+ZJp0uboE+kBfNmmhDPbryapw6kAiuBMpn
7dVLAx98Euy0+dK3yesZaC2+GxiKvrk1ucaxRDpAE5QwKz71x14n5+FgR67df8mkRaAHk8ut1RS3
Fc0k9Yi22iM9HKGnlM4C24NKQA2IbyXvYjl0R2bPT05CWmntymSHkKOGWDRxELoG64fYrmp2JCy3
v3bYElsREFVIA/irT/DwBjVndsrj3RRSJrfiEeoJwkPVao7LPMyv+I9b3ZETcBdPrZrpWfK8Z82O
cmBs5f9j4liww/AQRrvuernMv240AwNDikDnM5GAu+/gW/hcX2oa3Na9iHzYVcWv/Pk9hkqaZ6ts
XaOUzH+UD/Tg4d7N+NGrs64QeYzmUPF6LEDLZaof0eGJhKvqKDEnGYbtLGQSOWfKONM80ALbSbkg
d7jropjyGv+xDsF/rOe4UhDHLkvRhF9dlaQoCxjLAFxBlkEz5QptRxFQlz8gZ4uUfu+mVXfKf3B9
Ylv1vWTCHujsFbl+L7vFhmPc24zo43CJU22amTHvKQI7nuU8YG08mT/vU8tNoeJVSLhVVII4vaMF
Yxy0aJPzD5LXmqaXrmaj1jYlEJOEyJvgBVUFxKf/K/33IZ4MFyKYF+kT4fieLWJAidk1Sqp0dtnL
PePcyjFqwfyAbxxAL/4X3FmjDfhMICI/uzU25mJ1VAl9efP0dekrxkdDrBLhIhRD1nAG/g2FSSne
Uh/4WljWJ0uHzuRh4vNtVAfdDXUtOGetHdkSQQO1+3bRX9HJIGuZDJvqyAo00s1Fq0FncEIfP3kI
/AS5nWub1NOnIk5iN0/h9yiZHJt5jHMxfDT8rBxkerZ5aV5K5z8xKoAwMAFdeFciRFliy7NIli3P
/UOCeH0vW4IPBqr6/QqraAg79GqeySVpZe3S3/bOWXykkOrQfdzrDkPe14RTnMZoCBeUBfM+9M4Z
PEH3y+tiC19rNZkIi50nV1nt2Br++l+uQlEqlBSBi3aXSXMDiOpF3snJncXLFQQq5WaSGzQ+jEB4
BsP5Au4e1myhwEQxE5Tik8DwDHkcvWnC0YLdMG50lK+7hMms9ogDSfm9zbgc9Xx/amfDlosNt7tE
G50o/kRc86kILFZPu/QnmpOFUiOmOGi40zbtKCtO1Xrw/7Dsks2qYoz+Tk4OQnWWAJ6xf1F2FWgi
Pvvpd/39lzhE1tm6VIgBlMOSHr/BWHi+uasqJdzfPZTlCOFZoBQtMx8sySnXpQzAcv+9lcVIQabQ
ryUwLGFBsdydJXCg4Y7RJhHQnrSsjkLbrbbleFDnxiDvnDzO8ZcdznH8MqXGs9V2icvI8axD67U4
jYgfhu8QvaCI2emVoiDGALPwQve5vAuyoksEyPbFvMwriCx22w/Dlv+aPIkDmk7xCytDXfx+Pcnx
AG+KgsSiLvm88ylkCW+yI4EzRDxI3pAJjV60ii2rCYvhfH/MnPP9MKOF5tb5qHMwtAI2cICENNS+
qyHMirUnCfBGh36urySs89eh27FGdQcD73S7QuuU0ugpQvmw9WCUwQG9VdaM/n1D0WH1rsM+L/8y
dEX5jhiPvd2cPdUP0AyG6lcuX6MbxqgBjmywGihGLKqwZPY78JqNdfjZSsvbgcBuZBI7Pldi+5RR
G3Nh/4drY41moxQ3lYOVHfkdL0Ukco+mSp5NUTvR7s+JAnzRqsOfwJLPdCPZBxOA/njlphn15mMK
cvS/e7igFX684xTjwF4PQQ7fCINJ9fUCojszgzdbUptm45JBzQAn1azNph0NwdCwQ+yUTvYRJxN5
YPHrhFocprMAVguGLY2tBERbBELzNuATgfWQ7LfXq4AnH+pZV2oEMiSorvzwM7B+Bam49n5I84ZP
RpKxg8GZ/+j3E4aZq6W3Aof+fOjXRV/8Je4Nf6xzQ2QefVaVVOKy7Oof2uWBiuH5uSCC7bnDmpDo
IdI+8I+x4Xqn0RKM3Sbp5BvoKNyC3r9DbKVzm2pkaUfZtpq8BrEZczcGYYmUsR7jpInbAkJdLp1G
mAWtretEBYxXsQGh3FHtyC45L8j2SlhNPac1lf5XdlTECrJA7uzkl96WmG2nFyZYPFMdq1YslOJx
FvrzcANJZxjfz/oAjt3Afn//zI54NH8942Zh8fIcfNrPlbAsgdfZg0Liq0rIdnmkIQzVW0KO7uAR
n+W54oZ1zLOajHpttN0hrWPCdrVpn1LszVt8lLE9q6Mm0BKYQIcK57hza5Vr9EXCjo8w28pWrXxj
/x7H6WDgxPpzKzu6F8m2yA4wgw6AnbFu4r2vbEm2MeWGiraKcNNBcf3n119hbCOgvPhNOH7jNt5c
cWUr4k+e8jeHbXsJ4rPznoQuHITY6xh8ILvxM3zHSunHHd660GLwCNJjsN5qLyH2oRBrifiWcxwm
dqMmiVdYZ5csZ2dy0XQFlBdQDaTeA5q2q1ZdKvXyDomkljixOMpZmY1C6qmV+Q0s8PoeLVS/90sq
NI6uf9M56uFvFbnr0VEaMhJ+blocd0JzBZAufZ4UOssb68P22Qs2D7kAGCBDyK9Qgn7cQ4vsNJ2v
H1DYS6h+L11giY7+we2L/pWIv/T75IVe2KDILfAyKKx/FUeHWb8w47iht+6lMQU2UlryLsWN1wav
DG5U2aeTEdq/2hTk1oxJKl5s6kr6avyQYMFMzOraOt1yQ9ONjhA553xFSxWqiVdjv3LY4zXW2VJW
rI1Gs2n7jTHbksCshXwSXFXIjcFkZx+tTEEH5LZBhgXyE1JPWbGF4aWj1tPZtbC1wTCTcIuiIhsO
uWamF6NO7XymIfqzR6XSWjF0AbwuQcyqa6uq+fdq4awinW9ojDErO1ZrQdqxZ++NJM9NNLh5Oniy
IovNOZVo3naz+2FUx7xLJAet18fAqR2RZeNrqVCkosxyWjLqYMOC1R9VR2jeCCk8dTBne+qsp8/+
ni6eppn7qyBs+O5SUrvig3rOQS1A8KFn6KJaleotf9jv+PrBlMp3juNYZOwV7ghnl1AElR9nnDx+
C8FvndckPuNX7mrp8CN1FCOCrH92fWzzINDNOG8VftUSYLyTTIBzf8SPri3NG78AOaL3GLvlfs9X
Mr/2mvYNl9B97HimBsFD5YhqpjEQVCHdRj44ZTC9ec2miIss5J8AsBdhsdML6kq5J43bKYsykLaH
gH4TVRJCKRzz11iIgOzUohwvkf/B6IFDxV8qeYEDYxGia5G1U6y7fMm6h4gBjkYx0tw7TcwkV7NA
JmUxO8i5UxDif1Fzk00DhDKx2hA974QtIJEea+nKHWYaisQ7AzRhNdSjpNZVnXynO48sHnCGaRPE
5MGeUQiNWOynzw8V/o51/3/0beCgrLLKGVeqrSBKx74NY6xj9F/cinvk80+257DAipr3P1n1ZmyI
jFfNzvtEMrZH5YyLYLaNFZmFbGRZD9DxDPlKsGKszrkgWWeXyLX5MeXyFkG11mZGrPCoizckuYHa
f2l2KiIj1MuY0edOqbQX+KGFd0whwbBjhcYAd34mZ53PC5AX/a9h0rC3tB8K94cAHmtBHLUJnxxE
fhhY9Z+VrgNoIFLbqH+wcGaWKXImdtZxz3+6DPcF46xRHbq1bbCDl2PxOzJKhJuxNuB1/l4kJpvs
VLeDW3Vu7si1UHrZjq9mWHq9ZM5XURDFGbo0BUmxee3kD8N8OuXltwc8F9xBAWGiqZ157JkLIJmu
St47ih3/gNCFsGSLNNOAlvWytRe/dqfsFPUpHkvB2D43bLgjGjSu0zKO1CkTwQLl0wr9bgM+O6mj
yKWgbzp7REHLiXNe4eI9IF8pO6b/TddmOJ6KJOl23lU7BQw1YUWq7vPGZ1eRhzyhRxqlLlMrycKt
2AirIPnYqTBkgol2RX2gaM/JBTGQT39b4fA/tdTSmndg8QMrD0pKcsC2uRnqWA3sOBfo3XtvJq5w
Ej2UJ/CGCYO9Q40L5oPqjbCZQ+CkSnBlhji8bvGiidlCRadOTZAhducUQc0VXzgn6aAA9EK7Iqah
Dai8W7+8QMxszZ5BRjAe2E3GAVJlu2gpaoUUtu+ql95vVlGg0f1LG0iHKSidM9dP+bHUZhDu6VOD
4B8WEC1RkO/iCjhz996Ej+CnGTukn5uxBDvaDXWtkJ0hyIfhKrrb4SPF3A43MkpRjg+N0xNTZzbY
dN6JvCelvSoeVnKXq9ws3H8Kj3B+sqVAYJkx1sIWsq0+QyeQgxBA0dkd0ENZxjrKVNILO9/AtE6K
QDi+zkCHc4Zv43Q9WQiIvFUsU6ykE3fgh9Oh2QUT8sIbxrubkBqA72o7D3ZSRcxzjys0rPoyN0Kx
R4MWDwguV9HaWTDD19DSP02fIvgfKsEuMX34xGQvF22yXh8IuMf/XSnTTVoqDEJvTsCf6EyC0BOt
p+9J+AIsS+1ASLyUs5Hu6c2W1Dtu9+37QC4HuKInY7qReTMVFTFLLBF2EwK54WrYjMC8lkQyGFkI
AmaB5osd9Ip6WTFPLCe6riO9r+xBLF2znn1L1uToQOT9cklOhkkwM1NL4qqfsY9c/LnXLqrIy/G2
Jvyml3+pAbfsBRlx27fN7CIuoMCIN3eeZ70UnQxpRgpoPvDl2qMwUXENGoVfgOT9XauBePkiKgJ7
EEXyoGSWvuZNuNIh3CwBQxusXVJ5Hs70CjAWhOVjiXSf40PryJZryn6dC8beNcnguEAZzdkm7aU/
FDhdPi8l5SnQDpa7sz5okdftsG3OteP99FF7oEViv4WOZ84uUU+lXumBTf+wd3br8oEL/ePn+42N
khXYHAuODFe+JFPxI5uQcujcwOQVyg67wnPL0qkQvKFqYKmQfOFez4G0n9WnuadqXvhfOBXhNa+x
74bIYslsj8vskRxHs3tZ4oVR5ORvwzUz4pTAlIMiOMn2l6m0hmhK6xbOAKDsmsWsfe9oMOH0OC0+
Q0nG78Fo5opW0XzIMZThfcI9KxcWqVbYNQqpLfQONjL8gEuT4tvJU+2b+jGk1AoygoMm+1yb3FMs
fdiiI69f9gumytK2cO2fgrm9sxZXR34ngzz43LZbb+SldTSZwVDaJlR9pwlPUEvnuU5s7uhGqF3H
a1DaePZflQmVMNRE5L0D5+fZ1oswvdPtprhLpUcDIZ3exkLCFTLHOB1tTwva+uPhHde7+ZYEzzHQ
ceFW3dOPsUXcK/y4VzmDKF9kG0XVj8Vnf/dSrxQ4oJNTsHQhLEx4j8/6dABHhzxgcIO/CPqGbiw9
jNUDBitTbEGI8qx8hOchHXKLfpFkoHKiXLtoZu/wQSKUi7YT3XshA5hCoA4OIaaBHrrzOXBahpDr
YBE3PtB7vCguaMGQydGPNaIDta8LuEdlGyDQjyPqQgiJu6mnlIjAIFZ4UyacrXgNWjA/m3CHmO9e
/MFZ8Rnilingwhb9gnSKxEvBMg9nGfqCj0CO6ZW54RXbzDJjYjot3umQQaP9RkJYFBR1EAaX9wBa
gpRxXvL2W3vAiv3veB7hiFdqJB+UQMAiEzOUvaIClIJ2o4jGk9ZfrRxCdbwxuuMfoQa6dEzT+XKA
uSpqGRglpxo94zbZQHyuHCyvYFcNWYnk34zk9gAx5wFoxZgqIq2dzqfohcUz/ek/dLrwPEBltjg4
4cgHI8cI13vCIYegky6YNci7ua8tH4xSsLJlWaMOp9sO6LZgxjPdvxChXGlB9xsDZuiaUiQMxRf5
PtH/Gst0Pya9WqGpOe7MLmTnTN6laIviHzneqd0QqA2L/RWVFjWTYRHmdFOw/Fk2MvMYORSLiBRi
G3lRywYNAlSuwfZTsOA7mOLg3+oxLrqtep7nYpmmZCHNVc1lUHj/8Aff3KB1oYPBx7GoaoAuwYLi
AfTFjaEaSP+q9DM3dnKBQB8clKKbX2qW9Hk/uqczoKYuCcIlNJl493O5QXZ9rSJSNVE1odoOum23
TQTJ2md6Vla5DCv/QGfqIJbwNmu/In9KWcKLO28dKdC43/yp3IwjnyFdNlSqax8C02rwB9IH9h5m
kmeGW2JUTtLpPi90BU5VWAM7+7oQV9acgshTyyCzdOHv2yLD+H79w/QgvLyLPI8kTEdJt85Q8pW2
O6/69AMeqS4Kv8q8MY4T9Qe3qfZUOsNjSdUF6uCjEGJ7Nv3Oe9sTfsTvURisRVAEtgpIiDlb5kFv
C183CHq1FJmsBlTg5gzxF1yHtuP6QwyMp93wI8ckYz9nM37lMxfT0//YXbrTNmCCk5GKcO+B5WNp
krL/Z1xaIyaUF05SVk6ShOiesGVrGV22sjNFO64n1hOtPV/Yv8M1YYzi/xjjXJdDY5f582bGDu3n
CyN5/1y4714TPzdpV+oDOFsYLD56AzIjflQg0oV0XeK6F1FCP9G+NDiNkGn41e6KmCRUE3ckIB18
RsxI0ifrqDiEahDZYl8oOmFIdDDj7X9Eo7LFWYrZg+ydLjre6BJxvEQCwJSxeUaSViSryMilKYDI
3zU3YXdwtAT5f1HJtsDkQ9ArpjxmWYbFWK/i6yPidlzS2xWXamncpfP7c/HLVThG/GS0HJpPAm57
XTC5MErS2zwtymUayrzMrccZvxHaJKrwiFKgSXrsk33coeaSjDvpWQ/AJtVOnidwHjoibXb2SNCW
mQEm9fvqXqZyIYEC2X/TdDApFvA2NhfNvemfa+Jwzs7n0hNdHTA5aFEa/dHJprmVR/ptmFX4m4OU
cvkiyNQOVNnyuYQf67nMntAWFLA/XlLfY3qsjWzVtdzGurFGXA2Gj+HegOEUNL05P+o4JAe7lqsX
QlqtAj0m4mLzWDjTWksz2bXKkcvwyg3gcKD/tasinhHhnux5rqQW0LpN1xMQ1jFGRWs4e7o321X2
qYrtDaa0St0QofyYkvUsUjvP3JiDL4hLHJoTrFs4vD3T8r+raqF4TN5kqK4mPUDI0yXzfWqYjh8t
jVU6ubrpYs2KqW2aD3IfrBU8xztgZ5mLGEoEGt98q3zsQpX4wpU2C3IIBk1fokfp0DHSgT6oKZEf
OuQwOsHVoH+0K2KmmaZ2wKKJv5FOrxFNn1EB/RCkDxjPuutpMGX+r8zLwQI3t44LHNlMJdfkcHOX
Gq6HubDsAezsya5KV7KICp8Cr7j7LveDuicP634cgcSPd1+pzgVyKeC5FQ4THGZMWAC53Ww2oNQ4
XVVkb++XBMxFQh5rKCkgOGhT+4mvUx9zhiDurj5Gtkx8NhnOg6WQMhqw4lDOSijTvC2Px2FFabFs
b5MF/OdhsXs9LWPjsQ7TJqPAe2hg23X5e9PPsqwt9G40iRSQZ+32ryrA6YzDvYW/rg+ewMfIEIaO
LDZQSpPj3ELuo/3iqRPNBTZ06jX+nbH5T2Z9soOfcfknK3ZXCsFLVQSA+Ml5fenvGShuqGd7S1uh
pJTSGRL/2VUqEtfyaGkZm5LfipVrP7R0i8aRFJx+RPF/12i1lmhej8pGoBLDFwinlrb1xbPh60XV
m2Mubrna42ZdcBteSAJuF2e6WcwY9s/fFUibAg36v/mfPNwjaW9xDpK+i57xBpcQLgXh38IIifAP
O3AVpD3Vdd6ioH93uUQgiRQmDHnTsN/hkxuoZ+lCFPGpMdkD7Pg2ImZWaoTvPzC535gLIaP0pzHK
/Kx7MlNltR39petvclyc8D8DgYasCaMnTGijB7kzPst6oRuGrs+8d0bBrWpA6FTWHitjToccNQhK
phwpnSvzim4ipJb0PxlaJdmQNxAgdhOKcxjOLeqf/WMQ2xwLpZJ1re3dmgJxOxEhqysJqXtNVu4B
do7DyAzaLIZL/AUFPyRT6wNYGFrMHPQ389mElRqvmrULh697DmTJmouiot9rw9m13T26cQv/FJOJ
uAIF5Qo5C1iBVDO0dJZ0j6c8yZl9Zu9JU2CExePQhkIVFG2ySV4YFj2GLu+QIrRZtyJ4V/TChoWg
mr41FalFRMLaB33NacnW+UojrTk+aX0fUr08EvdD2bEp9TewUqx+FTG0H3KccCRpq/lEAt2JmVRi
j+m2mliqq8iakZ2fnFTxiDY3Hk4/I//ZErNT3Ktrw2oxisXRJ52lq0MMEGtzWwprcyJHjnglwgD9
upp6BOkO9xPmgdybNJY9TAc+qgnKD7IJpiVAgIL+18tLOeYHbFijKJbmf1mw5mAulOOZQw1twguM
MOeb74Tv+eeT34yCNnvugaGJ0Q8TC69aXH+QLlaYMwswCA0RzAL/XXmQRSuykcWolCg8IEAiNW4L
unBhzSzRyTWo8sG0opYoRtQXh5AozHYJMLx4qFJ1FQLcaefFauN1xRDUhApbEiefrSYhZVmiOcYV
Rm2LS1+0J8ItMeKLYcVLyIR41wqO4sa3lmMr9otP3lMW4IkJYaC/WxwRsY924CQXds4UOvZhXxPT
xKCoyyh9OOx1GX3wXo80U7hXFyWDzFD2nUkbvuEQHI8xch8O9JGM9QnBqKIrjQqUb7c5IpFGLdgv
czdr231kEPOi0+xJB0TKmPMtOEIMYDu4CHNhoGx+XBScL7Xk8JlTmriHk8TC1fzAvydvAobf6yqY
ACgf0i9LYt9lDUHbYzSbMNQag2OyQ6ZNvZ1OcEqeYeRnZyIVSyRFNxkwMuTWjovyLI5Cx+Lw8DsZ
oO/MGKctNqyMYU0DrsNrIZ45uExNS8WBpwjMtoLNr1z449KtLeaJeeOvdlekzK2igNRwpVfGZpnO
qwoA2pweNu7xEUAWG8NXzXItqeKPff+mlsQGgbtj82zFQLcogTRVH2lu/lhniz2eVU9MltdskgXE
ZIMDyYxyKXvqD9FfZ3EEVnAcg7JtJCjmOgQbEPq+vE4X9KJjmDrrG1i2Q5+VEp23eFKYS8+bWrXl
eSAZPAcaHyoH68LupAtbHvIyv7A/lhJ7MXCMB890puADllkp7moLXSJRlEguZ30dty8U4WzoTFiF
hOa9FMw/ZBhyLdncBovcNwjdYkR+4e0vCzxphz3EiJKviAXse/QHFkageyToz7tCNWCsv+4RhV5S
YPpZYWPwJi8lOUPBXw3jn0hp+BhMcgCaUTSnUTjk8vy2z3ETTxaoYQBgIDzoP1bY0AmqLYi6+QR/
CB+Rsj+iCG6X/Kg+UYlM1XjUFuOlKeRHtqmJvuqOEv97PR2kIXH9SLR2OJTVcSPoAeMgLc3i+t3s
3zhZi5m/ETkF5QwS51Pn9gJ8xAlFlZllpqniio+PAY0C4kuv2ZFHn8MifOy4W2GXdHiRdtyCAnHY
2msFbkDnje9lM7buG1GEHyXXMEs4vuDd0zRED5Qcj243CB5jcIx+VRS0WgSOte70GmWdvlPNZDfc
I/qiBdFqTnqzOdTQazOdF8Q1jnhytgieJ3/VE7/Wj7TnTB9/T+RX3t3bJZ2rnMP0rGF+ha3f7Z0V
+nVRxzwUSLdxK4A2QaW5v+TMJ4M0uEYghiPKqXhzmYJ8gynhj1J7FFURQ6wIDNaYiW29a2Maf+p8
OCEXKZ/dx72qhN7GXDd1MXJOU5qwKYnurAFItr2Mzzh1LJCDlwEI+i7UOv+Qj/H6EuElEauRVUlU
xv0Vk8F14JxIzYp7ghrXU87S8mS3Eewd9zagMHWTVRpuTM4/5xGQDlE8dlWhyr1qcMIPbRGUnkkc
aIVKNARDnj4cZOPJ4NFMbqIsJWkPWjvtmBVd5cQe2fNtM80spjFFwALZ1RDA/ayf8mrGuuFwhJ95
wlX+bQIXHVj+41c9KSscEoT026vsmgoXSnYoAC21sD9QHEMEenziwf+IZobP+f0EB27Ewll+d4nn
rKOWr/5cJOHKOe9uMzhzrbSW2V+iw2MSf76lNLtYamTCr6cFIz+E9ig9jfPMRQ1QhmSwcbeZw+Tr
472dngq5QNtv8fx2E7VvIEhVLLHWvng+0HoE2IpjaFhNQmw42KgbOkjT8tJ7YNaSLV4DW12r2fNt
oD3gV2465gP+0KwkT62iPgBSrd8U3oUbjJyXgnQigNb/7WSsALDA4oAeuBBvW2UOSL9A1AtskI2m
w9K5ZNN+rbLUvjemlEoMJGYYGOyQOxhPEZqUXPjoEgtLDWUv9X8irEpD7M9wGBoyvVwB85MiwS/D
DMxV9db3gLcnxChR7ThABwVEs7afLyST+W7JtSy93gph7IY7BKOmSM0gzU68W0rA+VfHklx5/aEi
mP27qR6ra/uk2YSDxFGl6Uq+cM9p/arpGpY03vqLvWLpMGHtI4tPqNqSKDZKLY3LXO4cG8iYqAHg
63AdO0ssRcd7cbGmN8gKi+nkxpdanwyMNfQEkHFwxTE4NIAJlP6KhOiQJr1AEvtoL1C5wd7BrWf0
StbY4YxvlcNs+Gv3ajxLjwb4qStXwD4GwCOqNJ2hG19Kv0WyzOUdITW4ingxA/ISovrTWIMOE3wd
wb231wja7GX4LvCizcRvg5YXe5Z/7Uogz9Ne2DGNnig2xJZYJwfvAuRzcKbRv5hLjSCcEYCa++1V
L/xxXFeb7WaPKzydUKDPjoX7emF/fuZFAPhg+mjmpcrFo4mn06GcF6hoGMPlFEMp9maXH34K+JXS
GInUBj6AGuZqMAirLIR4CT2GOQ+U7b+ChyzLax/PA0k/nDBIHF0S/xtePREfHUej16KG8HoitBih
XmPFFfhr7RY6EpXnrLV58coAz1q9SBKPgk7efPWo6wmS4jUd48Huka4IxjQJhyHTl9O+iB2NT2dq
0r15Y62oJQ4jRY6EhgBS6suYSwn/LTH8v0qLPSWGrgDF9fwuEtpUmovdllszK/bsruauZ9KZzw/z
SIOILwCmkb/YeQZDwZjJfctDgB00yg8a+KVRbtopnnx0SsgFpYDIaBOS11gAj0cKYqJCuiCN7jz7
lSz7QNsIa1e10e9n3i6XkFui6HeDuOVI3PubwerJY0sdvCI6ywegkIuFbowXTB4qXxQrf8zzHDhh
hu2qcQaVs1TO8ixLmJrDDnXsWbVVMCaWNALazZtuPwInOyew2KBh7TB5pHxcodg/jBh5i1rqeSzp
o3gDoY5nA+ejeQ+Iaaniw9XhjGVX8Vudfv4aPnNGuhvpGpqct6Bc0hj+33MMnNS3Y0ZO0ThIWc+y
f1Kyl4majNj7BHWfzqZ6VL/2IjFFe/533B6vaJ5ZnrpxUF3TYlN1cJiPmZFrXwthbRo+KMSYRy4h
9Ex8Tphz/lVGIVC7YtGG0DGLEG44QjVdvTiVu2CrDNmBJABwiPIuYeO6pXHmIZ1FK54tgD8OFXSc
MOnKXFooAuqFqyjoIJ9AqBF1q7MWGT3kNFscpiZcHBKcCZeMaE97TqlBnH1TqHfkhpvk6iuByFhy
8EjqLHmYzTzQ6i/42vG1prNrSTTj/kkDeX8LNmH85JrosDlqoSzr9fjMEnlmOCgfJdpLZnRw/3ho
YfXOmUpDrC1k5j1J123QD18j2SmXDzBqPzxKUjce7dONw+hejzBsdJw8PYDBpXVb4c/UtIpuJuIA
avd+ub31L89heynno6ZdBa8ypOa0J66/QOYxkoZ+S3qoIc2c+cnSsaz2zrimC+qFOb37bxpC4z0t
jYhJyOQlp2QrrzPXVBVoYi2skvYwBSFNGk328Uuy34cwlw4dixqKN3KsE0pySV+gZM14yh20Y/c0
2wueaJ77s3diQ4eyG2g6inamFFF3x3DSxzlxohaZNwV3Eq5Yo60fiNa3Ngbz0nD/fbI4pVtHi9yU
bNbDiJIrisxTE78kpCySgmvvUzV3/b8397PN3mro3Z+ilUkyC2tnWUkilSEyrXV4Ro6skXUXjO7C
Kr/KRgBwq3DBnYKI52GH1pmKqMX+4o5gWrVmccj/+eDRjdr39XMsYRGRC9m3dDLlLIVLZ1ip46bu
s5FyESUMk53qdvtNOzlZ6bb2b65aG2PENl1lxHmYDmp5Vi8AN5OWOHI4Dg/VqDZl3RJUy/UHmEmp
vXnmOiFcn28Urk0+xumg/ISTfNPFcfktrQyd9hDNUyxQBEwwV6quFlntfhJ8i8z7ay40f+QfKx/7
v9pfEy/WKotkCfEYUjW/oHdWRdGawDKjj6EudPY7SuAli/l9/pxRGsKxr+E/rKpIyogH7Qn+OtsC
UDf/SUNKNNMIabPtf9faDo/Ip0LFg4t1yN3iof9adBcEVRO+iP+WDyT6nDHrLUFiAnJok4ny9U65
FpaBEdbqQaVeYDbyxzGu9KKljUZTBY63rv/qIECZmrgEZ6YR3aGCAs3Gj+pp6pqTWnVovTZyItnu
oQR8gkRpPNTs/RIxTPSDqLVapoZtqaM/CbznZrW+UugDIV+7ehSROSXEs15Vkf5BvM22V1Rk2AnL
3abFxz9I+kfHnVlxZQckh9iB/Z/eTrCShdVUUiGrPrbqfeD3KGivqXG5gOsFiFn1sKRB2kJkpjkA
IQPs3JnIakUEwQsZZ3rWpTiXNmamQFr09ZEf401iJzp5y1rmASGI2kVD43/vnIfZFs6OMh3JWnPa
Tsd3HhGR4ssg6GaL3oLb2KWqpDlYgAm2oCzZCVdynRYBcA5E2jH7CQS2qU5xTdkj3NqJUcbZAECb
dDlz+G+LvUCw3dTOs8z+kQ1rUb0xV4oYMoMDHIiH8ynmADzBH6SQwjGs7hZULHVp3005xbmw9xzV
nmwRya0RWrxa+sQh48UD0Oen7rlGakwFgpAlTjZK8jMP+InxgfTQm64rvoxPbQcqSV4a/a8QFsk+
sf/z/+TmOVgjVghruEHjv/qANVK1GTCG3XJE0t6lhOjcjubuSwhUE1CgOZXZuSwZC3hm4zVr+oQq
InU4W5RZnlfzrQ3YiROpve3mi52kGcAB/hPLmnsiiL/k0VCA3TAV/g9Ge8gtY+JbNU65oBf4OzQI
/NrZ7z4cAGGOG6iglb6+wsKvfquZCH4Zc7N+NBTUIZEU4/w6Xv/OXQwOKB9s1rpEYvwp4c67/8jO
ZZkjCSCJTfX20lFOzOpQ31fKW1Pv5Q0Ix9GuONDDnGmkzBnJcG+iZIIPB7bPIVwM3yDT+3CuD7iY
LjXdeZXUFWUkP97MkSN41WrY/38Dayd6C7fLU4LTSStaw+T6qCq2d4vOOkv9sTUoGE5BKzUS9a0i
IxwbV4xV3RE34nxVTmx4YjhjM03Mgak+Z2kvn3AUNi1+8c5y/hCEvgoMMTFu5psup/0zkbJTMk7S
k3QMv1xeDZFIX1oPvXDngrDyoY8ESvH8uomIc6AF3WjxtBmeqh2Z23XIpaUT0uiwGKFbvOKVCUYl
aRTwNgFc0E7HGybWQS6LU4KhxfWUbsZbUMmubQlQHgJMiyOdXXfleFinyhO22l/S0KO8B86eXwfT
0Q8VLcWlPTVHuVZ8Bib3kuKgaZiYkluTceJ9+lJP+A/CIaXUnvyyQgZxtV5/kSd6kF1oYhjmuxt0
nj9AhMtNPKrm4y2YAXBk282eWCz6fBe4JAgz+yPkMvvCVJ73vn319VdD0Qv9dCCQrdO7F+VX80oJ
VsjWCqVs7Yakso/RHiINTxQyV0hH50x2Vx8mK24ejurYf+vnfHabJDbQeONp7jNRDgHUK2I5gwid
EA7gh8P6cF1kjZURwWJ/RlEWdld41bWV8pyCIqmI7eaeb2OYKYeDRjt7qffKJHli7uixHckk8y6U
G65LZVuTeeZw0jQ01XzJ5pVdA5ihkDCzUJ9cRlKZs9GK9aKO0eX1Ndx3ldCTITaBleWgLCY96Jlt
UUEPvvn018otn4aRaOtgJRXIrxFZjp5m839tdAeGiExkrZ4yB/iHInleenOqnoVGAV8loFhgulB0
2dFJfnmCgJ3pm+lWp5uqo59Q1uA04LiL61OWgIR6FveVu7JS12jZI4Ag0iqrRuEWQiVI5XU4toXP
ReQS7CAuXmra/7XeDWwFJLrI8ZC0sb+I4oi5Su+tTBavVB5M9isOGvOetVjWrs6ibWwcZf9DufKu
GUlBcrYkxX8ebOvL+nPN4FC5N1o5apSlijwifd7si/JboiHbTEu+gn12g3IQTO++dSJRTTnWyABB
PQ997Ubw9tLH7tk4pSlc3Npj1x47TFZrwHeJK9B46gaqmGSWL2/jZmoQS/PRwgBnptMM9rcsLGep
xsV9Gq06jBnive2vl3EfQIgU9EQ+1T7tVknblUwIdhEhycK6iDpy0/GZ6oN3BhpLpgVKV6mna9L0
tqhCh/x3XZ/cfWWutcebediE0Q9LYw0wAV4mMaWb7pYmYU7kZQjBwlixDck1y9pFhPBMVxtPNSNI
dtRD3MuVihWUKxNT2G7/X+Mu+JRQMCAoYyunyW2MMmBPT/Y27jABT5849txdDW+HtFXY+qCh0hii
lJXF7vWqe9A/jPZ7YKTgF5JYfNq/o0kZadzFWH76EOQYCkx3S9Y+3t/DQcQiZpazGJUjldi6TR5f
CT2Jg/jqyKVNzJ7N6JoptSsJJEzDQBsWywPUVEiaf7wqTZ4O3cXCBFGA+ky4Sp0uJPi2jYcY5cX9
FSpdEPU9ktJap12i4lGuVk5J+30xXKDGD4pqFZMFynq4LMrUhDoonOy5bb18y6XxrEDEx1GEkIqd
OHtKarBhgBCl+Ayv/HjmmraLizGBTywNyYZuQTGExrViLxWfJCTW9wpOnnp2lUUXn1dttDU0rJLx
2gwdHv4lcqjGF8C9y8XMVAuiiVAi+iHaqrrrRIwj4sdxnqrOJB7ElDcgsAFguAXU4haYKELReCRu
cWhhKEJTOTnH4TMwWajnv+NqRkT+AePu4L9rmy4iRhVEJ2Ox3Z/EWYaLr2i2W3Y1rW5iRXjSC0MY
AsWqf5l0iO764RpMkMwiwaME5xal0eqV0X02+b0hRvKqbdcC9u69p+TG6Qhg97arSTtel2iUJVf3
kKKgxWp8PIXJzJR8oZikBdYSROOjSg3EV+veJFvrLFJ2JIhQXatlxyu7Mjz7nxflin4HbAq90oJZ
0iKZTWqmmLcBlxurK2dihSnILC7o+9KrDXvdg1XaEYKNSMrFrOFQE72TbFbzk527wZ2okn17/fJQ
z7pq8WMqp872laUO0RcLa+bnuid6VKlufUxdWr0YhvdDyA7OgcZYYqWbO587MesQS99Dy3Ew9IiG
odD9jjd9R9aMSGmAQbaXlU6cWWX2XRT1XeVmLY22OPw8assqkskRm/EdK13jk7vYOFUpZoueDdzo
4R2UpuIFN7ga2QYuKxZ8gSPe0DULCWGKTTeUL8st4A/vN/15Fp0Q42/WlkFEZQDUIaki/2OoFpPS
M1YrmPSeRNWC8apn0G0BHYG+JgJAHg+eC+rZu4RqDY1JgYmJgKhJEUVuvGoEbAUqlUlJM52Vdd7K
qefSWgRax7cGVfDkYfg4ew4WlLsbhj2Ve++hi3A6RsU9aHg72TMx6NZOVE/4XEYtUHc6nKKgieUp
PUc/30U9PHYWg1ExI9gdGYL+YVMSOHrUYmQvTsFrW1cFFta3skksezbK4JLGpbKbm1ECA3QAFnWK
fZvpLCPvuC5WIzWW4FCenfaWsm2IJN1vh7W1PipNe12oSDLlHDBPdUfUQAd2/41/8moOCSA5sP/G
kGx13swwajATXFLqBlNCOUMOS09PYgs2vtwUUB6kWh3yAk90rMkvwkB0wJtc91hQgM+pOqNSkUVX
u6fMRFb8gjRtt6dyPU+hqKNwCly9A0d3HlcV4/xO/yRmzsb3KAWhxOXtH1jqlxmiaBkGMZ7l64Bz
kvZcnqMN8itI2dcqr2pJ0xtnUIUtjzOAZQCkjDS5GRsk6hJdjvGecx8+Yk7gO+m82nEoa1g9i253
1BZKnYnl98s8F34JDg5JiGtIVCtH/ZZqehcXwmYRw1KmqQBNJ5ruM4rIO5ZxLGsZf/hkyQrlGnZK
qo0udxrw4lXSHP2dTH+Hj/iasJ9ilHC3PmjUhEtz/Hvxav55+pSSUnxRCGU++ut6DtB6gkBtw5WD
UcKIFVLvs9yKLbKC97h3ET9fM3bdGcT8CwPIxHVXDTnJ0Q9nFtpUEKYmw7m98mW84HJ7mM6ryvCA
2xqOHEevaVsFp8Kf6MIX5UEP0fljpajN48RWMXTeW7mOK9ReFjd8AShPhO/wZ6OuJHDKIwm045Bm
qcbIXEDh6F4Tf2pcrB9OARO5ofGaiWY9wHIF0zoHWz6WEUh8KiPXGgmHUFVpk3578Jim9/tA1IXb
8Duhz5Y/Qtsd8CJM0eI/ix2Fxo62N/IwORUyfPUNp6zEHaxli59aHI76YxW+RjnXxiqfQlNUOPOV
oSJb7/7BELFe1SBees+fokqC/ifHOGfDpeYx8z2sTWqNP6oiCoh5+z+eIH2lGUEEpE/0Wnt8neJW
2peFz9F9FPrJekEVEUkmsS1kmGpAQ2PUqqgO1SuCRtAlUzU8TzwxZVqdg1qEOctnSmdLQc7qX3rY
CtWLjU9o2Vt/U7kfhESBN8Q+AqQ6Y1ksFp4KthE+kM1kUvwW4AyQk1c7xHvN1Dnnol0GzjS4kIB1
6SY4SjysKw2swEcIVCSP7fEV0vFgf3FEBnIwbInYaWu5qN1wVulbgeJbwbg/WmKgYzDbc/811Stv
2zsPuCXG3Rek1p7Ydg+4Tbp1FJGR+4WFplN3t7qeVSp4/pOdAyW1BIpVsGuF0FvXsoeaR4sJZvtn
VNBiuuz5xjeAmoYYIcpy+yH4OjIPfz6Gq8L07Ti3D4cCioIn4zQfWRJzqrUxG7+CubKwsPJtd+GI
I8KAiLMykLU7i+ahxNJB2kB1cieB3TsSvzCQUZ2jqDLeI826xuwXyAkTDFisyb6sqxh2UHrptiuq
9Ci7+m4xRBqz0YbR8YtVCtQTN3dVWCxWaBL4O9jtQWDD5JOcYyCobkc9ZLtg0PyGjE+FokcUb/qZ
JF77T8Ry4/4uQbhetlj/2i1hdDMirsSkriGxITvXOOfZAPxGzayWLPZidpP7yXrwMj5UnAr102TS
P0YZX/xUZST5KCmuG25Yogm6FeT1fJHwOtOm0YNnwm8Lkdx71DXtqSomFyFV46kK4RKgmON546Hs
i/AnkqyrBlBV5QJRjaq2IxYlJV0zHuwDZ+oKEWLT3j8c8HW62o8Y1utyQJv1k8Jid/0LF2iKb+z2
xD/d1M+F/vNNFgawZGWccfijlIQ0Tevhzi0r8iJxIb5X6kKpDhR6NsOCsSdyIzE7Agjj+uH2p2SR
JC0gYHME13w4le468NSJG7Rxdpm4QaBQ6wLjeRR5fFVxY/gHGI5Il7LPhTKo6OgUpSbh+yvUXTW9
Av3F6VNBBKdoBqzIvFTDaKJZIG6I9Gd8KwSfykyJzYDLHkVdf/qHNEmUbZ8fYNb1kZLfU23+Zzik
5JB4Yj0fTDkGUsi0+DOEaOXaW5wX09fdxdba5qy8R43a/nYdGv3xyM4BOa4tF0IvkA2KY7fpbFkS
kIPGvzsdl8jeMbyDawMV2YZzaDN/rtKGsN6fFJ9FCI50sMnjhZX0R32wRV73ijeWnVS6qzvTRYv1
I+ZA5u9P7scpPRkuMWh8NCasNh6+4A7KDytGVE1lzuma1CXZfe1K5FHwagF1zHzAmDz42QTpvk1I
ulrVjdQ8Npm60pHsABMNruwZrvYnI7HEkceouORQdngwJT2bDml5b1iEijYnj5gHZvrv/tydI4ik
NsdDTuzk+b1d1eJSfp5l73V5qXPWSNByzshV8dm47Pt3sMGocGvI5rZs0F/RjOFqc+hC8c+dx/CQ
siDMZfcziBy+oo1JsoHvcVXjXYGH2Wu1rmUwMTyEgMQtwCOUfWqUZRPBB5E2f581xtjVrXgSOxUe
ClDn1MWhGJiO2GYcqd/fPmf+BKDeYZdx3LfUXPtPqOzWuPktDWt0EldtbHZKa51iWQWkfKE0Ty+Q
afuxt7azR8imS2ZWi1+qetZmeBJE+H+M/IrfMe+GWSE3oKk6dm/aS03TDVYB2TMffftKXRhiQhMf
9WNxqzQmR3aItvfbkHljsxpBU+yxVXZEXkrdXyS6cHdOh8u2oGPOqQt/hHEDKxvDX5Wjfd2div3C
9+U7AE6aHizN+pwkW4HpC/1CnhaBRnI27SlRV3eqH/hxyfGN3PvQJnS/3lfiuHV5ByJuGUNlYJGa
CfSeEzIZp/C3MA99bzMQErbSl00ujyRscLZls9l08csA9Fnu3DQT4Wgc96tqbIeZL6Wkx5nJLZS9
5czRXIGgKAqTfGaMr75Vqqgr3ZrFxPfSf7/YSTGsPhDMSWZKKS1vlvEUAc+WKAtzvIo5FNH55uLC
cqxzrimPYIkmUS9xc2m8OdX3NC3WE+nzXZ+rY73e65c6fVKUuRxJDH4+mPdlQ6IoP903SXIWJdzG
Obl0+BGId8knVYmPK8Nf6cdngWmt0abbmQqW6zpXdUgC63PblJ1AqFivMdiP/NfcqyEHylBwJDJB
4iJrBbJ6MnaaKgxPQxDFVtHVrHtSykp4pL8OuFL8ye/Zc9nWyRZiTiaBEGxQOKzhYSdU+8429f+i
LWHxOKDKKudGzvMt8qFix9Y9FAKqxKi4RjjNavawMlZbYKThDayLQe/QAKIQHu20jSvoCnJ19JdZ
bEsal/jDCD3p8jB5axtbmgbaJCBt+QPfBEsTpGUSU/SE+ITNVdiEL+lxIJ9iUgfc4eiPiz74jKuh
n3F7eCFYKsDZFVCbSgkrg0f2aI+Oz9pqvcv4LElaDHce4as8tjL9zEv+NcEavtNUD4RfWk6JO1mO
euNTe9hAOuh3+ldiI5WPwGnzrZOQY7B3CeFWGIvwGlqiVjXZ/Zi2MEoz51GixNFVF62DXeYaZEPa
ZANS5uqVX6lg3kse9JBw2Kq4Gm43/TzyY5f0QpZZasT5lpg3LzERr8PUHnUNNVx6VILwTK/xc+0/
wOb4Poycz0ni2hZVybA2ZVhKbZFklGP71y8mNoFFZ/YwopCCTajpPuQGffPiAQ2iLHTl2SWMOrYT
az4c0uttHNT1RJCPncSVBzkFyF5N46XOAk4TT+ww7YH+ByoXDO8dWWJHAc42Khy4qdj2xZyqoZ2x
4nFXF+Xm5vxOTWtOmJ1pm2ug8oi+BlxWkm95/dhXad+8RhwRyss0Nzd7+Kt7srkNPVIWHIt+Zrlt
I13s6PjJEIK9T7Yw4e34Yv+Q/7eA5mLFoex3VFPqqdtOG+/Ek4LOXJ6tUeLq07eoo7by+r6JikGc
wVfT57mreePE+Rmy0C+LWXWcPf1nkQ8Qmy8+Ljp4X0U56epzeDBpgH6VCfEl/b3NzuRt/SdkfrKU
f/9K9U/XniQ2BMYIHXdQH17GAWFhyq5SmrgueFRVgcfPza0kovdVNzr9xRbNlOoofDH2sLGaDBq1
ZacQiOSMFoR/Uu3zmhZBT6MrjZVN7zUT61XZ9exgNq07VI0ePVLUkD6SXf2zWZ5niHn/jVEZ9ddb
B3hcMjejWwRBg3TAZsJUm4LqYGLZAuKCJ2ouOxU8ZlsK30QdtqL9wEfZF9uAcNfs1VBTkFmbzAr6
vBZ+QNHx2MVKWRPYrBx3ol5O2ZqJUUmKDLTmbBksqdCRMSR+bIS5c1oJiSub5DqvUl5WjaLQ1Jx8
JBco2vO2MyMq9Q1Fp+BQbZ2S2ZMdA8hHG94jWFXYgra479uJPE2Ra4ABW+vTVRBVOEQQ1MSsmRRB
U9QC+LNli2MCAlHqAnVIexrM2VnpeR68L2yqBxAS2AvOHxSyi0UGIJnNwgcUDa2XQ5uvKIN2Xbh7
KpRrFdIrWF/zZzKFam3d0jVdt/CnJ6mkGxMHmp16ebrCjmny3ZTmMWGHeEeob+8uOuvlNGNeLFsW
Rv1FBITSyRRogY3Mbj0Cxhu7juoyVk2VoXIhVjs0hCl+FICXx23HttjzDzXfKkpATYbL4IhE0Dqn
H5GLTw5Vs5cK8WUqGmnDh8YpMhxeGoPGsDnH63uApiaOPulW/Q7JzAMLMHztMt4B2aRHNef1IWo7
e6AN9+iaFRqdXpBm1G3Fh0CnutQSPeBtzpBDaxxXkJL6aqgJ7lUS6maDzC3Q/3axiQgdVpiDR4Mr
czOobLGjHKRdd78DkpXxAjKEjDdNWjywG1ABLE/3CNwQtXE3ges4mXnRAsP5wbAfdjmr0/sqsgab
6Aa7nIz8zAzNJza3fRCPqLtlMVTS2c8KyUtGsm6zaO85gXmTDkL9Q5euXHGboUE0/1TZoHuP7Jk2
qbgc3juhiRHT1LrNkx/sjM7gYl7MTj/UWi9vo4pBeSK+thDzZh8yO7B3Q6aIgfWwiRJb79wXpZnH
mKfnW/T2H0wD3nIXbFKptmgxxxXgykJ6h3Vh1OvhbtaLcftULNCOZ6F6bCIXIlHs94YP/gr9wUAC
1Tbl6pTKCT5faZr3EVN/R3XOCB/F/WpjXuUy5hK8VKL6P2VkwURZPPyX95RsUUg0pgGeS9mQ65P4
cTQ1cPDJ+nkYivpPlucIjcKxHB5QqcvqG29XD0eazjeQuN25WEer5GkFjFq9UBL4L6kyMDook3kY
mPFJD4VBy9N8LUkbvUZ+S4Nf9qlKw/GRCIsHTxs9LoMAeeQefeBWMIAiOpxh56ttNlKMcsO70AZU
u+XmLdztc6NH42tG+zHs52HgnkKMkVxeljdgzvtzLZNfowvggSLotHfP+YXyAYJiMWfhGKfHW+op
AMDKSH2/Q7ZyP4+RzaWBG6DX10ApJETDQc3fXnhxlCsRqPWfxyupEEGWJC43TXx26RDohvPw21Jz
zRL9PAKKatiMMtMD4oDwerIrOVr5X9eO8ouc9qAW460FI47pXEED6bU3LcJb44RxTS4GH7nLC4MQ
/851MAOazzfF58TDHS3l/DE+a8tVFALtgW2LlEjE3QzxxXgD5V/aVzE4YqSVCKCgW/sssXWaNfNZ
8Wj3yOCYcrAVkckX3SemFv+gQz7WXhkuFXiryK4KPmk2F+wLaGLg9ls8EpVJSQiS3fTJMlR+ltbd
RaNLq6pLgZJttFqh9vozbQ297P1inogWh/uYIpScbjim0np/gjhdwtHAfOzySbg9wx1yHb7k1VxH
3MXbixgLuD5i05kGNir89vsQZSlmtph6VmB/CXqtMSE9eQh+PPfi1A9rTIk74v1/9ygYgxzKY/eH
fAoS9YagXlLzmkWsNl4D2pgC0xRc2cHdHTFlICqXDcVQxsURd1zjjfppZU/xGk1ufAHeS349VoWS
Z/kPawEzSs1Fzt4KN2CO8JnXTw7X/cC6jXAQouuL5x3M4Cp8atdvSE4S2Lx90KPI5jnFT60WOLqt
k75/9KW0qEIT4U0K7chnEnnwdcNgweTUoxZuO+Dp6YsbcblgIAUZgZMiSKiRGqIDve/v5mefMNsy
Ucw5q4PeAL0/AzIRu8kA28SPgN5DU4Vx4x8lUK+gwzMEGBMAnpAFZnyIxKyIbUUm2E32sEY+qQAW
PpnMVQUpRnisDWYHeZC73/Gb2EZLJ+8hnd85TGoNLyd2a8YZMZs1G7Mq+rfgWPflPqV6Jq0IdNqy
mJGpugSaTPNOajc4O7FbM8M0Jd7LjzuqUxA027vDmVgbXt3xf2KAMdFIP6HJQ3VGhhhc9R9WhJr1
1laNUKUBj3iM9UlvUjiXsPqMJlfJQMyD83REuZz0gC7DQWDObtRyuVxC0eJhNx1eE9SgjJ5949Id
iiX2Y1NOvwTmInhCxGAOBIU1m9/UxhSdabvU0Jd45YtvHLvsbKH7AY6OrvA+G9wHkDWjE1leFozF
p4iV+tOqd/eiCjRA4jF1H54s9m+0vOkBC1TtbfHSerlS3HnIu9tBw58UlZswC5F28VsyOAwR/awA
kmoJ1PojRH0FglM22S6/083WZCqOyE8m3BTBeEeiJm3HTy/yFixrKRrvSBA9Fa1a9wIgndvfDo7C
Y499Bo5aiM2wx3vacDBfVxoLc7a17LMWS/lWbQ7nLJF9SGc4WaMxQ9EA7oMiLqJIWV2xD12chotG
PPZeEJmzwIos1NTLi40Vl4hR5mOyHWf8uG5CiMXONhX/6VsuYh41m/ecEFiAQhYs5BcE1H0rQ+cv
hmY9dXDm0tmFxGUl12f8VJYm3aTR2x55tOqZdmWhnHLBwGzv61BREj6SOl2i+thQnFQwfyPKYmSz
wqSYHJkMcdFbO+C7erTO8Ox3Hav+ca9XnMcQeYwp1Eanwe4FNcTpHpSkzRMg5QXJksCi7i+3IxfB
gIMrImohecIDAnUziC23wwO6YlLLcFUdylqx3dMfIZ1TJEyfhFv7BpSSmEr0jXrwvi39ATFUEEjZ
E6hQylbQP+ONDD18vpYLTCGDfizqwCmCQLVT+j/n9Z4j+XoDLdpdCvaTvs6RLHyzCCco7EBhZJPi
C4PBrVftl3wvDWhT786/pLOq/GXRue8zpEatoXql91E+8tAfJWW85zaBHb4oKank3aGVD/4ZjtSN
yS9NOoAvpRwVYiDBi9IiPuzpGTwpRWD6YsWZqEiuQs+zkFzAwNgT47Bccyl1/85u0+4llWgPdCc2
Pbspb86RIhcgekkythruv1MxF+IcO0CSdfKNF9koYldH/v7zUIDwbHb0U20BePLp1m3V0qE6F49e
1l4dRNT2yNhAffxNhQNZ3yqTLppuEirx7gAaUESEWnTghedCdQbT+vnSmb+dQB2mRoUuvjr3ELHN
qG7hvpyq23N02oK97JkQ98NT3HUjSstl3dAegMDKsiOQ+cL4ZJCLnvAckloKRjHPYL6vE4Svj0pX
oUQjnxqYiOmgcd+1AafSkgbjMlHJlVBoRLinTg2rOEzfOh7n/mMeRf7Z49L6TR/8EhkqfA3F+u2Y
i5uU/1EWOECvnUz6NRoC+pBNJplMLd3T0A0RkjzPxPlZFacDQ7ckBmtY43Lh3PFYAKW5Ki9bTYWr
bazY5pPgHEyWam0kvg+zwqvJJRQh4F24xnazfdf3and67OUn8qyrGwPChD3i6deQzitW7yWeTMFF
UX7NwENMoU7rhG6aFItxXWv41jzPOhT6O+wOsgYvr2Go2+7QbhXB1I/kWJR3l39Nt45LCmciYsbT
Kp+yHnlLN/eiZsjVS/GmAhHhr9nFYJ8RITbn8JyGdI26UvQWyGtt6j8S0ng+pc/yLpFcpi422pwl
XNE/Ct59S8c8GU7uFWyeA7sp3aXk53EI2WTGjEjq4JSo1YFxkoz43bEyf8SAUOkqSZ2l/ALIjYlQ
0GLzDw6wB4vhScMAfKclduuaFwC1oWCN7SdvO4Cxm+mnSA99nL7YhHUT7nMty/T/bt/SApckmqx6
jVZaFQJeNgclmZ0XNvTfg6ZT/ofNFj5X1Aujrl2CW/Fs0Oo37VEmVre1EMM2G+dqgAzPt8Jr77LA
lB1kzbSp7EbTf2pekiCr6AMrjz/cQLEBKybslgFupNdyP9ympJahgs7383Qs6hvIdPnpfObIDiBW
Yu+YLp3oBU9JpZNmZ8W6iqowxnhyN2yY59x8GeGDymKm43NjENFxujxcEfxODW+74bCQB6SvTnYs
o/5sDDwbS1Ulmii+ynbr/Yk4jNF7Ey0eFaEG3FhO3jxOjmgFwHKsoCw3H06bwXQCgg0vXl282J46
DiKUUsznG28nun5IAlX96nB+agWGX1oKIRoezJl1h0zx9SKTlkRE3tQgzAnQjcGqBnG/4du7KtMy
/zvmUwrOYlCMJGPMOUpFl0SpZ6KDWpuVXbGjbDowWNu7X64MI0NLixlAcgcHa1eDnS4ksi1R5WxX
g1s5MfHk5tJHjdeBlToUPb5fRzPl/s5uJwM0iHKit4tcv/rfq759BSo0zfsh0rzSimwJN0lmEKMF
mlG9lIUEMFXwg3UAGHyQYjdmmJkQjK9dtIjL89xagBvbzNnIk/VVpdXT+WhPG1SqwYX4fSylDizl
z4xItIrEBtwqYSCnqlzPSKkh6cHnyTcUoWgOv7EguxooLBvr7upsp1UEIXSoMXWs2uPGe0VHQOWj
TQlhO0nm+Y4NtuVzxaeZS1W2dTrOgfLiBh691GSg/hdbr89yZjbbLtAZ1N1IwZMU8RN1xP47cfYl
4PakMzXswWr+fd5ImVwRkREQsL7nteB5K0zXO5Ac0BzwxEGKAWhtwq1qokI0ov2Cx20R5MR2MANE
zrzCxaCdL64EyYCxqhORi9EN3NJxEN0XAMlE1DXfSnoqeJbBHHK1jF6mo4rwLe1kouZsT8BWg0lN
6HKtwzPg+HF9nX09YiixwLsHmwWt0WakJQVeyChzvLBhakOXaVZX4mj8TChpXvAURuscHr0kZ5md
OL1quXfHjNx1CMkEHXKDQgQQigSk+rbzVdWWJd2YD6pVIzOwPL0C1QPjysnI0QiGFG9tUCdB4J4J
OGaNnaaBO28aQYSNekXca+f2QDuR1i+Jyq9rf9cjIeIlDfu9cn08iAq/XCy9A4O31i3KLDqe+hL7
eS57W/znek1DkjDjezH8+kHf8ua4PC7vHXd1M31cn6yb7xk/9mAUefJri/AY9A2WnYliAoJp/sdg
Q8C9BSTKw/ZHXspv4ar6FzbwSmBJgwnORDIhbdR1V1Dh2h5NxMrILKL/3vOyJtg1Sreb4G73tqIS
HI2U9tpDuiP9DVCyss97ZKTTc6ddfyGKjZIc24TOSmRlj0xHy95c9qz7WtHoq33VW4xA/MvlRDZB
1BH8/WaIGGtzjfMFdBP1IbYd5qqpMWwpLvGadxQZDEK+RN40puUO1t1nQK/g1RQjyacPnxDEOvs/
4qbFlWscnxp9XG5MRVlpfnJgBACmTuzflpHKsz53fuiqTtyO5v9iUwNWxMkqCMfqM8AWd5wHQLDa
FZJva9qfFHeJSphwEO23tr3pKYLdOtLWpRCgyifM3vlr//svXME4vkqbVdF5MVY5NjiC9ID0YNG7
U3ZnRy0AKvHyvyM7Rjo60OTa4z27Klr78lWBZD3J2q7AQDqLzUjbXsg+ugb6LK6PmPoMRmBYedFd
hQRHzBS0Szyddno78CvfpTP1xwxcTG2Tr1n78DfYLSH4vQ/yq2skUiVyG5wngUv99hgelvdQnPKF
xkKeHVRbaoVi+WK8PWAojTt7Br7UaNERmJIBs6vCrLGHntdvlBhd+bhoAyYS/newq0kscos1upfC
B9GNWIUvsYVjrJZsB2wxA6NlN2Y4a1wwQVvONjYRyxkhrkPCLkSPVfnZ9U02U/p/nVEWkBCjifb0
ifxOHkHJhJaLO0PX1+uXFXEnuHnUoQrwsd2FudxJ2pIr7Pnlu8c4jdcER4vTMRW6LvmS4nthD6PS
OM3/E81oChdiah7OrDVz3OXzuP1Ha05f66ZADfbH+pJV/CMR9c37Gza3oJ3kYHPvX9DG5KVl2P8F
WsVdtH+xKQQBwpVaF8Ffs4bc3f6JJSqi8gTqoDqtqRp4FhK+a84sJfNcZoipFc7Du+8cvgk59eyM
ATKcjWCGN3FU0egqOSltiOcFnLn0d8zJEW8olRTt9qW1vQk8Cd15iib94fYv2JxW4MkCAyzO4kdE
W/flr/yXzRZgUAbGlWNzs76m5sDURP8TB3M7PdYDQgSYYyZqQJ7uxGEShawwRVDvzgZGF2L3BPlq
VXt7io6eSNTsRQefAx73BUqqKrz+H/vgV2y2TgYI6hRhTtgYTwwV0wKY0KiaS0UmCrkot51YymHj
JaPXyPGf9DRGLU/tqK/6bND48ROtim1uMiIKVKOWoVwd3CTjUaT70jTg2fpMT08xLDk8ODaY3P9I
yHWwxr4tRTlXRBm1/wNoryCmG9uWJ8XSH1o+Imi3+pSkvISLv3u3ZrauEnAGsoFfdC7iMAEzwBWc
n7kmf/460ZH4USmzkNnyFbbREvzMaRLbYLnVFX4WgPSYJ1Exl0Yx109pl/I+eEgGRpvHXAaX/YEJ
ikBuGYzWQHNHrxK/zcajapQeM7W5j3ThP0DO0IvmvsA6SAiHQqNX8lR68mfJzDN59IgYcmWLJhQk
TOPRz0eyETQx9KjnVnL/X1ju30din0gi3+xvoYz4q36kkzWgKy6g/s5p5nwcTovO8MD56nzKt7Nl
i/mOVrpYqwvSkoTpYlqI9vvDjIawR4PIoL2KMayF3a/gVc5K5aTdIAWcjM5lVKWUungarPpoj0x7
EEZMgsRUaYeaSuF5ZO7FWpPIO9ra/xAmha22l9JcaMAjuUM+ewYb/CK74KdvociAsKFb9c3KSL34
JFGv7kZ6lxQa5PXbmmT/W3Kf3Gh1pbM1F/uCdsBYGYdre2lOecbYgC8lcRCVtLJXQCQkRGnFigVU
9T6lq+MDFZ4FzsH+bhmOZ2i9rU4l4PY28fh4LCK5vpp/IEGa+s7UWWkVTUQDP1PFDD3RlbKuCVdb
ORRvVqXH/HiZYiSTP5jJB09TRuP3oZR4ld6L3BZImaqhnRV56E5C+GDj2R9B65avlRGGokR/A2bt
EMEJersJ5X6087SCo5vM5wi7BFv+RvDbQv1yVY9KY0EocjATHqjRFLKKeUYFbEearY8Z3M4KC+7J
hd+WV8/vohDgSnRP93K1qqTb8cZoi6EylolRDO0YN3BT365RDo9E3aiE2qNFmsRpU1m2oihXBBUE
UC2ehIgs4jvSeavTckyLumU0PyrabUjPw9n1qbqIi9CCqxxDjSYMmPGsBeeMdraotrZ5UdaALOmX
V4lm6KL+FWO/RCTEUcEBatUj0LRhsIJCWiVUlwLy7ppAwiOrBOFoxpNMu/LgzPz+Q2imlPTSCy+c
nPvQqJhIq5uI7gBPRJVy5X/LBhUS6hhDBGRXY0p55lOPAbaEV6M04fi/ApI66V/BbTobU5oNoMLG
BujS3LQwNc7ESKqNFXFm9X49iMrOw1MzwOGTmFZLO2UWZHwWF8B4gOaN2hRdpcDHZc/02JgXsO6v
PvCyzNZIV6HPkZfA+JejVRdJjejz2RdzAGLe/jhrGI0eyCAw71370vCGCFpV1KJXL6Ee1TewPNFU
DNezL5qzkyeKntRDHDdyDHtkUpTPvU3FNw+ZiGBwSScpY5cL+qGpHjiqj6gQBqN2O3FcqWUnHHs9
+2hDJAZ+WUDn2G+KhsO3wIkHPSSgMtTzmyPP9lSAUbeyRRmuqF+dsB6veN+ongIyZDkPUpyYpeRH
tpcqTFH5MQysnkVdBhVqgLhs0ozkaupkpw3/chcDdQk/Aq3bwVqEw+ewNXD70x5oUXJdp9KeAm6o
N4uv3tXjbVtg34ojQnFIJm4Mz7FA/gWfYeJyqod3dTcbqf0vKKJq+vMcpyE3DBnb61zfKUFW1kYV
I4DX9S9CaNP9jIEcZ8aga533KR+wZdBx/14U2vSl23bD98aZTrP5j8qsX/kD3ojgzmJPwzBkCBXX
r0ZcctVun3mvz7D/OIvh0Wa0Jr9lghDO3RC8mBobejmsdwlk2DlDYLgwS/DCEtGkmwwSGjGtyxg2
2JIt9kqgwcTJvTHY2xVRI2w3gHVglbCzgY0H9ZNIhAHgAL7nWu/Byz6k7dP9Ldu7pYp80VMfXX6I
OFJQ3XqZ0NJtKBWsgJR1HME/1zR7Mrd8be5MxtIb7RSt/OpepS6OvBE8pU0XwKOFsth9oY3Drgjs
95BM6R3hrQO56u1neltyMt91jVX18K1AByy8nJFb3ULB2znF7BCvjT93WsYZR8aypdg9xIaPuzgG
+hiwO6Y4rV56r/749L+n+l2vZiOh1Q1j4pG/g+8cxLvDS7RqBffyIqrzJAAJuw3jNok8amQ9lgnH
oJoi83RCMOWEOefhntwb7hs0XkiOOfXEv9Nka7MsPgoZKMXEfmZ+K/iq0W2X8ryE3ZApBgRYP21H
i5pkLxyYACgqdrHmJv20Em/H9oNS0pVheX6ikQRuNc/0aR5g/0OoDmh7sArCj5NSy00tjyiPAYbq
hyFL3lNf0Mf/v2xIFdRcEkcIRTMkqzt4cJeEiiGJ+QAb8vDY5WDrzVDy7yLhAtXnHz2QJBL5ZDWu
tSpfSMBrR5BCr8cFyTGcCl3SLy7LAtNkAQFmGanGMRYY7GhGH9doK2w7XRDgojcVAdJraxE9FIWx
NTDtaoEp7s5bSRCoJm/FCyeWMowYswYNEHnq86/Tx86Ser8rz74caSJf4ExaIMftstFoUVigta/I
6ULjdrQbeFL3kevJoSrMU2c4G+EZ8vCNWh7FaIAFoQVs8yhNdCtaA+LehDipGZZ+AnfMmK7MvVtG
zKGVqswKAaxhdUUV5vH9kYYB0GD70vnGHxOnufoJdN1RdhNC4BFdkecImBvetzQ+ofMfmowa1RsX
DMwdzdKnCgoupcH94xhCejLHIbeQaynWqlbjTFQUbzDbgLBoIaULQCwuahRxKoPi8/BpPCaSxIqf
Gr6iQzY2B1iwH4CIyzQs0cKe2H19u9Ojm6JTjtZbcVVdk6bAUhdF6+ej9UyYx5uNxyoNA0O0D68P
Hd+ogX5qr8Az0h1gX3mCTWIzjugvH3VB+1/Wb5UFRoa8GWgzkdLj5xNBRHEwuaPMtnLTbjhnZqE1
Kzz8vEr28xalrAg9SGM+P7aYcCQMgUT/vomugY7qOBuJR6LHlvxAhNA/IXZXK420gjFJRNywxyYx
2WYTa+YAOvvJyNhPVgZfV/2ZMfL/XRzcsZPk6dlz8/Hq+rLOVEXnlErqskZFpNdfBsdx+o3vXoWb
36gvFVaz2JtJjQimbv8KgkA5h4osSZwWhGc/4wCqUqdFY26FhvR9BS13/3C9HFCY2e73QjKyFn2H
1p3pWx3J9Wq9c/sDZRuU6wjLNu0YZH4akpA1HonydiW+pYBFwcfpW8iJdo0coWyuNJbr/+i8AzLc
j92yQJERglyckr991g8UThSkNyUlbi2Kbsg3rl2lvas3cXBCIIzr8nETvq3Ql3r4R2oLJ8Kjhi3S
CRyYP1mksS/HQquJ2lxNKnMe62XCwvcusVThwJ1ju7aeXtjzKOslL6A7u8c6L6lI3mHhIEZebRkD
E2WInxKHnaC84m6pc2PIASzSdkpUBZPS4XXH/ujSSJXZ8VJtPJzPxHySuh6maiVY/t8MtTZzJxdH
dQIUFwa7F8w4y9tZTGkoSVI0IfQUSk4Y+WeB4wRUBqnEA834A5g1rxnJMrgBJJkuMlsQN0s1LXZZ
wDdD0wKQc65ZhQQ2wmiVpP32Uf7UHjzy5XgGA/3BdfLuywkLbi2YDPfNHD0yl7IrNBx/b/T+jiKh
13VZmoS3rtajxCVpahWJmsGin/ojmUHKxD6wdBPb3t2ExflDBr6gvN0FRzKZpvKmu6EjH9pIdzYP
CcaiEdj1KvU2ZiqXqN/N+j1jG81epE8hayFrdG5qKwLNoHFwH/S4L502aZ1d+PnymeJPz3NpIvZX
6EFbPiqxv2ofSXnF1CoVC05/rYryHyX8PnIa5CFgUjujkK01GGGbGzPsYN2aoe5hoeg7fFROwaMO
0JtC7IclqwYK2LEiWGNZjBQCs0fzrN2hR0hIthS2KCoGhsKfRDaG76GSEa1nmJhikUxmKSco2gQl
yga+XQWlA9OCFa7bg7P2NPyWP9K6kqmp09utzHKhKfHfc5r8VmfbJXr8Gz+nrnDYyOSlLh7Cu9nS
yla4bMXVJB056UK13idyuwHBaLzotxoap3oxicjRDgAKCd7ssvuW+7FSb/jDv/jfHsFe5/9B6QVp
yupqmOd0gv7QvIffl9JzgWNnKI1Ym+31KTEpIc4tCe1yrDFz79W2URXNl3nRcHHuBi/gzTDuHqI0
m0+/7JBKd+FC4o8pOkdImcSAoZHsdFk5gyNTeMvGN/GMtXifv2YJoh2dys1GK39jeYBOSb8VtgRG
TTnDQ1KlJtmSk1NoexS2QdUgC2vwf/fmka8d4T0Rdyml+/Bo8CIhA+mEpp6HR3Wl9AAnFhrEOnnv
532RrocUblC8dWE599CrK8XyMnocNopVOVcuoWU5gSKzENHjKIfhjVpAKpazz/8hiaYKR3d138z7
ZppOqJpaIOGrZkP8nBUiVTn4TiESFKpZHElv29TUmH6IcxWprBiFmSVMwErzj8B+4qjuOfFpnt1A
ImdfCLik3Va+BiI3r3rf3t5fwADEAfOn9fJhYI5VqnalKmaLxUcPahffP/wdMYmHR6DMZti4EGGU
xl9R0/mSZ9II3bU9jTq4CE4sWu2BCjRAFwi+Nj/teX95YBiPB4eTkdvaiccH6TE/4URl3gRHiEGf
boor5jQhJ+ROXtmx41n998j2lfVS9ijFB4v9T1TjmrtZCKK34Y9JGMhPgo5Nj4u9ppYsSQZ7cQZt
n6iz6uwfNXhguQlej2SZ8WbYEHmSOm2wumPk9do07Q8c97P7gedDmZJFbccIEuXkd2KC+DhvxUkE
P0oUdtHzNFJbuNJ1EFUHfQMgkoMP3c0GL4EnpqfGSl0z+OsWTbANOlQqUFfIYrVu6TUrqb+LKelc
BUysP/5c6It9iFYI/DnyUglxvpu3dmm0OX7M3tzbtaXV3lf/hz5IPtvxhW+1ONudzcuS/tALzTQD
DZurF24+rSYsg5VLNpeMhF3CHJofGVHAe3ubAH01UWUz7nGBhvkx4kD+/cju6NMwzSIRLamQanyu
hcngrC3Ug9POfMGcsoo4FETRT/nUOzkXXFEAPNO9lAzaiRsdK3eTxTzE2hC2GdVy1V63MazU/fis
opg0hVf02yjy7W9c/+T64lm2lQ/4rXO5bzlgB8nGEcL84B/XtAqTqkK3Zirp+LtLeOeE5Zm+5Y3e
gJaEQsu+jwq4+hrS7ACVVkZEOqgB9rmD0X2KbwkMw3F11V+GoRO3RKMRILFMYOmwttCKiJbzMRIY
CF1yf8PHZIwKGoKV+lnVn46YvnIOqM1Vf1d3BIZvcbF8YeMcZH7dvpqyQhFMFz50Q2WN5uNvVUtK
gtxAblr5Edc5jfKr2XMInr9NzaKHRY5ciLuSIqvde4K31kencmmB3hoNQN6zsJQWJQd6+cMQwciy
5G+hIL2cvC4MV3oo5lI5axmr2PcaoLKneNoSOjjCDvRF5gaicjggYuyr5ohUKTyQXsDck+DVLNO/
nNIaWFmSJZbcbXq7uMD6xHoTBgzjlPWj4Hu4dVgi00gxCU5WepPS/pxQXynf2SU5JHSFuvMivB/u
swIfOQHqo7nDJ/kI9cQSl89TunfMNtXl0HRrNuaNf0gGTbCu3/it7P6ub+ffvyS/6ju4yG19VB9l
owkwhk+wvBBtqP8FFU6AplvI2qDqXLMlqQlOWX4do8jgqeJReW7/vbYTrWd2L7yhnhbKkFWlRxcR
0ZIaf48AGupOaAJMhZEv4G58lrd2gQk7FUobs+GiZ1Goed70w9nYUrlqpNPrvIzMiyuHWt7B4zNO
QWHQxUYf3XaBkweQot3w0SdUcfRgpKHWH2AW47udxccoyiGSl/e4HYEh+ZJE8RzinVwUsnBAqjL/
BxKVFfy4WLsh1y77OUAxlFPCwdnNlHs15iyl3XiS8Z5fs0xmrSZQRG2+uP+2IMBJNQJSN0ZSoY5U
0+zq2VqDwB+WYf2tr7sldrYYX8eOpdDxPNuK3DbE905RfcQf1AJA6X1tBJpcCqahNLRLFBBCbZZt
0ZY12Pc8ESeZ+IKf+pgLYmX9sliqlJqCoRC1bRffz4j55TynYMveMFaOZT8ZNIFxsHNBL511Frnd
s1kEdnfCnkKagDgVjM0ibwf/RWd7UR+FB3ZeotYjROAeVokdF6l/28cOMcWR4Wq2nx+e+v3LLMx5
uFskL4yatuIenYRgdeeHE2HoP7p0mIhovs1KYZs9LOOvozjm1tRGA9anUddlOFZoCF1Dl8e5zzrx
0LUvfLhXlIgbrrGjV6HTqBwYPcSLkVabHojA2i1ETnIU+W/xAvPZznT7euSN0lCJ6PFYLpxd++sV
gz0WPZ414QTlOLFM0KZ7oWYSECnKEEV43e6Nkc2kNTJDZRJSSLbo9om3yuoCTDVgwgpfUFopXqjt
bKJ9t1pjZ58Uy5qZrXEh4/zeGy8UVH09Iiipvv11zatAKbIRkAxawhTSXpQP+2G77xYv0CuhSEpd
9eZEY65E3H7P3LNj6V2Y4q9fSEECbul1rdcROAIId9ka1HLSwGuTqMbi6rlwDqy3JJOFS+lhIefG
WK9lkH0dV2f82VbWZB1qR4fyRF5wTrWDGEQj6jpZxbrSNw+0eVjQHnFqRdUuMiYJBONo6aEktYps
UtumZBSYN1ox0lziiTWqf+mDSw2sBRUoL4TZvGH1dUO6vi7alPFAz66Ur1kkRxX10wEJXd/RwcTN
YGtUt424Dyxzguuxim5AbReYi0vaywdFUGSxOyN0grK0CBNX90gXtS2wZ3yFS5gtUNLH4x1cXYw0
PpwBj9hTmuZ4C7WruamGSS9d3OWPR96dnpE22qM/JjTMh6DVmYQkF8GCV4SyQ8UZGGMLetTCN5MF
rE7AgQWNgtPUnxwb/BaTEgTFCG6kaeoZ7u7h4vQ+Th/gV6lZ75JES/zYkNtmnJoSSjmfrTBy1xcI
kRI/FQ6nsoSCHJi9/GAyqtbBF+6IIytLhNa5mI5pi8fxLs+prjF3xZfOyJBQlknTC60jduRw8Qp1
SJtZ5+Y9msrAyJFKzt/Ps5YiYSTfWy+12/PZGR9BNqt/ZDu8z4KOSDiF3/GvspMYPxzPDzl+HjmC
3pKw/NOXM+87uiMTRZPmx6cb1heIZ8OdOm76bKoEseIsXUJhWlHnUcvGNRmOlhwB7VGG76/OzIdJ
j2ujvGnV7di4jJP7XJJzfsoL/b46VRPGMKTOOMotJKq3Dvk1flnIhVEM9rP3je78DVSPlswPaThT
gRVqb9M0fWYsNSW64QR2q9/bdSoflI8vyzOMnmVsohQ+Vz4AnUXUguG5k2WcUEHycyEyjUw/RMAt
G2Cw70f8ATnOXAObN0uLOK2KOA/wFoK7hyqlw/WigessG8gUgqT6IQ3tNDY4cA5QdK1RiSDORo9K
lOyfaIEy6csZPRpsuv0m8qlYW7Db5t2UPsS1ULFnFQoRSeXS3K1RIzjCdagJgYbeXbSlNUcLUwT/
yoGdL3G9AX3rpowJyhwKFVrENiTvgqc10vGHtza1i8Vs+n3q9I8y4Vy7O0mNyDJbZZ5PdsoQlAxp
mazxtlbqXrwPV7FmpdAkQIO5AGNN1Swrj6NNp89laUKlieOsrLLNnMvv8ZF8kaqTCSGU61jK5jas
iWuK9PLVh5CAyjJS1P9xb0dN3T13OyjwppED7DKQ5OvzfAjVjvSTzNQpgxkZdlLmVl9m+SIBtCWg
w6S5BFAQM8V6VWfLpYVekPU7JK8i0iGDj2NmJHq0rix4TC7ClSPrWiASZQMt6+1k58ApuOxbWy3T
CKWliLd3CBAJ2JSHTIk+V/F93RAb0PmgMEUqXEfFWGH3e08Q3jKgRIzMsoiB3GbO7teD+t0DnUmH
Qi5ya/spfnTnn3IlIhQAOwld6sJRLY9Kn1gUfTu10L5pENoNaM9Bb5Y+dbGAJv86vEb3NO/GwBIL
FvQCCTGexpAzvdjcA4OgTDnsHsGZCeEcsY/niV6q/MM4FKHVjv9i3BrOp2TxC2nlajnQ3B2iqBaX
eb65sU1OAfnFygTczWoWwI7Ckyk5H0QFnc4Knn0hidWOr49tCRdDBKNhM998Ip3I5FQTRVXr/OA2
5WMatfRjGQkNmqTyjJ5jaKslsAzYowIgBGdUJV+jov2jg30fDjTEshpbMcOJtRXz0sVNlwsUzB/c
5AoKWMhoW8A3dWqxe5UkTVWOc93z6/sV7SuRkSo++wZAvh9qfCKERTfBHzJNfHMRbn3SIsLpw+vv
F3To9NkWrGkqRB9F0ZLnOZ2YyRhOE8vlhGjBYBNxSmvjxhLE36YIP5dqlUYWQ6IVWLTwjr+Kp92M
rf8FVXt1e6/Viy9Y30oPISOfKj8HG6XX+frcn0738uhG/7aBJUqI/5uLyhnjsF8XLFdyPCvFiJU6
9cOJ50nb/J1KqVIRzv2QxAAneNAKG0X3qR1gGr1Nbtb6YEgDnp0pHlnPx9j7emRVNKX9KP9HxxHR
L85dGPv94afijTleUdcZFmfCQoY11hJXEkJ1iZlBC2h8tpN29LIdCZTrPCE9PH0okiQWruhcMHm+
Yh8uXHTTrk/VffZ+TxEDivjkuYgQMAfbqFn5xkJKt1vOnGH+USDMV0T2VsJunndx09TBRMfuBDaK
T5I50B3zEalj7EAPTLTBKvN+/SpZn5p+xux2/Dkk3JWcC+NxitjmjBiF48cD/XSop/NBmVC7Sccv
TCzpqQ3v/K5Qx2a66C0oDgXXACq4SbniTPcrd62l2QAyRFB6pXOS4xNAJDhNzGe4ZVZ3kOGaJBEl
wjl7u4U4Rqrpwj3dKOc5Jyuo4Am0usaSkQ7Q3Tr9JygBMcUgp4pvd9aOw4dGxh5N3/oCvQKS3rJN
QgB99qA0Gfgd1EC9BFJY55H1IxfCGZEGYNb4U7fs+W+baqjRnC3QnW4txzZ5Q10muZfAkYqGArpp
Hebakd55maazXkE7LMRyGoIOq+S+ebddlFRB0sj6swKsr44ttcS8Bt147/F3YK1ZxTUrZEWEFn+a
nuFtjavNdApRfb3Lop8x0MxxuvIc+cNgbDZj8cVffFnkwQO8M8ua4pzD5ZrQXG3fh37ow69CvZfo
Se+O7do5DruqhhNKMvh858gnzsQrH6xa6zT0SA33Z1N8bG2Zdql24FBGG2Q/g6Gswn5cs848qkKs
MLRlNrnjU5UFb8cCdpzJnS7L98f/ZcWeQnLb44hDiQwOTf1rVZvZN4E74oAdQU4q8bmeS+gUNK7n
lFKGbcVtwMWT9bnVhutIEQrnwMXQRq8Wss9JzVz52qeDAPJEMMLhisa95CtzHbAmknVTJBUB7U3P
4J+VCAudx56y9AGw+A6Yf4/8Tk4sPZho45W1O74gzH1uxllDwA1ozoDNk1OVdSQ8OmFJJBzRhrCn
TYhTPx57LeG1wHdaIyuapHgwgjgWZjm0oVDvJalPMH2eLo5OClGX6Gh/4LPwYAeC4RD7LcZKP9AI
eGfBWPaC01G04ekPlR8p4za0x1lXUcZ+MirNCEh439kXXDHWJViTkBN92BBAs1I8X5NuJWEOb7yg
LSzlq+sXtxSQTHSkHba41quWullFCIcfsJMuCD3Xq+rXdvskpNS7NT0z1d0aczx3OE1UGQLMx2no
9V20j2Emr/ZDGwUEXcnWajg4XObnJNnv9MZ23lpVxsyNT3yUdxIv5qjMrnrVxaEvTvhe67uQOP11
mfn1F7PsEKZByppVWsQrz4nlmkaibyy3oigpomqaYtbXVJrxEsJGrOP9P7HExvJ8GtPJxQwhJYYA
6VmqO5BQbu18S9Q2vBRqWt6byH7PjzYwqYGKcztwwowCirmK4nwyCMPPMNfhhxz2MhSjgXmEeRIo
6U6W1HxOBStoNIHiWouo12tNKuWhbt0185c3ZjAcU/DgqS8YSu+oBR1GoBTDRSP+zvay4kmtSAir
7rZfIZBoin1f8VK9+FQ59FrQNjv6liKVxSh0aZvl3xBMYeMXyvwN8ULZlHfbnzSsh927iEaRnQFe
aa036MaF63P2MmOSQ2JpKopoj9vbkfhK+rUUVfsjrmosS2HGh6sNdrAhtbz6/sDKPWdBiNfmlpWr
KzZWMRRflYPG/3/bNgEgVfqG+FcJLT8NC1vKo7Pv7y5WvS8fnAaop9QXTEVG0mPxmetNdeNaU0yQ
iL5RhQP4ERYN7vxhBeEqZJ3/mm4C3Lm05mexSSuFGo9bMbSEgyL2F5Ij/rbCyT06k/liri/+TsFC
aTqjYO6NmaEgGmXAVIDWnITaLNAyw92AAc5bVHe65uW3rVhIcriuO4emspt9X+TFtLR5MAs6CE62
JHgIW4zZd8jv23GsGA4GgMNSlPKuDiElYjeDHsToo5Gs7B7dl3Ud7Lua0LIN6sL+aMLnU225c165
I7P9p19qEsmRtRYLavcEIOnvLzHzj5dndTqOtOlgRT1zgJGX3m7jyp0pH0haR4wadS9jvs6uYJFT
EigmU0oXmYe0wolqb6jBWTsKOsT4cr3bb+H0pJBZr6pA7JGlEIgJeAVpcMwW+GZUVTii9B5pgDKQ
y7k1MG/R05cetmkXE3PpSsjmxYdExWlAJQWaaklmJIjsUOQmMXHH6Zgs8CzRBp1cwIXaB0aG+R5R
eyHoFQVLgDdPk081mvjMVfrLhJI7In7A+uuKvFcMyTQdKF15FU++bIIOOevtN22o50e2uMjJhtEn
lbpVHdVrwNV81nNJDYW/WaGKHv+amSx/BgbahIoJJoyPxl1qraC4EPBptmMU3FBwayU016C9TOti
yhq1JXThScAVVQTbDllDnGOWdiIleZbNvvI38mU1LNc/xBDDQWL9zeDGOWeU+c8Ymck6wDpZkFnm
GQ0STFIaVQc/8+woWbzE7htNgo+Ne3mYT0WCXrifI6bVYRaufx9oA1uGQB3TasHHA/kpwzaHnbYN
OSRv3uuuohxLA3XH6Vta0xL5VpjRxsqXk55lFHQ7vpBqZaMJyRSU4nBGgKs7Luoy3hkQH/v9/uh1
4i9LALfc33w99nrZ66YBZS3bztF8CVgIwJ1eeElV8f0YYQTs3KDRD3X9dAkuzw8IJUMgl2R8zY/u
xFTy8Uk333b6kQP7ifKhRQO9MslgyfYYznTzWfDZt2GAZBJOZ5IIwkPymxtbH0z3/Y2ckMZn2MOF
NezHdF+IoNv/ZrfnMpcFuxf5W4M+eAMafIE632FzV6dhuDBOeQX0DuRzMrZmWpvx4ZlIsY+gcBJL
raNtqJdp6a3iSZaMgOEvgjskjItB+bTw1AGQCrg+8EeVUjulaFPDOZUECPKOjFE68+CEU0NukfQ5
xRAccdUnSWT1iLwJqJOEGxXsWQTBzYeeEF7219Mi32YaXsQHfoJ1VTmfQdvndpYXVQbj5TM7WJfi
mbRr0Jx/KGkyZDmnJlHnfwrPU6uykelalCsXcvHt7OOgTVh8fSJzgK8AWI06X4zUmVSbOD9JoL5j
ZHhnjjWac+KvucdekwlO9XuzQhBElJFRPeQgVKSu0GiohNkcXgtUytAX7J84fW2VZUQ+7ZyX/whg
0Z5v9aplQc/GehUppW9Qgxmvo+m8bZolIFyPJF8kskyMEG4Hgo/2HgC67/41hfGTR3jrWqAGBbVa
6Lp8hzQ50rlxm72+2qoK+oC2U+RJyLo0gMTL6UeVS/ohwbIdl4rYvi7lq6kTQUUYl8hRu4ZiTtl9
4CQ1UrSxG8sVK09mniPJOKCQtwgHNg4w79pYePyj9iPvb5fv6L6+Dt05kq6M4ttgIrm3UA1SIq3j
LqJ1Qs6PSUjRzo+JvJtf+3SXrNv3vwLqIeiRQwm1kIJaN1zomru5o5k90Z7iBBFIc0yRkDPzZAzP
9D00coQCP23UTNlKm5o9qAUNmvYG8dGCNlFLIpIVkDBTvEDFrnPVoXWxFfF+VSGwpQuxL+JzOlxS
cNBXjhJ+sL+2SZLcP2+xcNL8XSm6t2UdV8GznZyPruiD9xzCCpwJI12ND1G+r3EwssSF+tESN2Nh
cgKYJoB+0oYOdZl58mF04z579VjcizrcUG4D7R5lHhvFgQKIohnmFZbuwjqEWrGMCdG+yaMNzbJq
/Qh1OkEA3wTMbpJp6TDoUP1DGotiVxCsK1LvmJgKzMRZTu3O0paA0Jhds9yqrlcWvwY4+zQ8boOS
+Mb/YD/z+5HlVSlNvIHgPGBSfSqE7zyqaOXG0bcgFAGmi8PcBJso7yvHfkIwgan1K4GYOCclBVqV
dWrjxblHGohzszIS3bgFc5XuvKNYxqe7m0VTGDqEX/A8CcHbzP2+GA+Q5AAcybFx1t/XOchHHV9s
pFIt35DjQhyEMiqkI140V8HkcxyBfXmxxqaGeShrl7Lqc0Vlv60TwvnTxSe51SM3QIMKhqMFRi/T
DwTAV6ei5yXJmPKGQ/0bTSaTDQoiTnFT4OtP2SMCmsGvGUeN5HdTzDayMFFphvzKYq4R92cpB2DF
krTg0BlD3xvYDkJMaLB8JKOHnf13rQXU/z8rCwI6Uyyh4AQbkFHh/i6glWd/ESYTzw8nHr+DWVDT
XuYKmjxtzJnA4lE9RQqQt6RnYZLmco6EzY10a6mKa46Qa4n6G1wUbVgobOn6CHalNiXh4uPqvbQt
oMPMcGNC4kRKqfs89YnjT0QUj/Yta/YjmN6euK8F16tTlX+7SvDGQ0GeLx2JQ7gW8orhK1/7Yc7P
Mc1s1JvOM9okcN/yDAMyRoTXrKuyMR9crJNPGNSPwOn9w4+wlocxEvauWmWUIB83BKSE5bTZm699
lISmU+uNDaxQtHglM+kqygyNCTSKHMI7ZhNz0Tu2f0FJQN4lhPjhHJpPhU0G52en5q5wW5UKZ+qA
5xyWENrdXi0QJBSIcgztE6inT3fRmw6AW4wCiUvhY1YAnXdodvWuIVTQc6hO1rkTkhb/CEm1nK4A
/rzBHzKmm9iTWF54aRbS9oKC+2psqiKGKZ1XZF6y39XQtFW6qvcs9Y7CrASfWDTv4V2LCLUjI9aP
QhhPn29baLjLeWmpEQqYYsnTsvfZ2I64qYJjlTlL1iX9ZiFY2BOuIijuN4smZNittTX0ltz86PXi
JXRnmuZ2MiVy30LYmEw9x8t60n5DMXDh7qRKDKVPYGS+mN9pStHaPhketRqvYhdO0+x4q1MpaTP9
wsA+NFcODi0QVqQkDWShuCeTZLtLODGk62pqknWLwEWn3ko6yBQDtjZvMA9As6+QpFGrTPx3oIeB
XAV3ht4ombMDH8TX6XFHFq+pM3pwicrr7pKfDAwWtWDiYQmtm8Mp++dYuQxCtsQcbsjnKrPdz7qm
6KeqkqBlwDEkh6JoRT4NvBqmM/A4f4KEQ7JMEnM9F6nHKuSSlxcxkxRyTe54LXpSIoeVY1HLjCmg
j2RWT9jSKTOqQHW9/RsczNPQtEZu1XkmLlzy7F9Xm2FNNMTBlZglRYuYBs//BWNUp4gz/MaubDWX
nYh1wR9658wZc+cNCIATsellM2GNEYeOKiGNpXUdlBPN2BdLtCe9gTu7GSleb6lPBLo6SXa5AoT2
OOKVwuE7tiMLgkv2KLyjlUaRoKi0XzYEp5ScSiPYa3O/H1ROrcjN+YrkqmvcSlyk+zVO3DSBFYMY
+HUriv5AOCLKabYlaSij6GKmimzyJrYctu8qRXa0wYc6wi8IblhBM2HmzxYtB2gi4HRiS5K2si/a
XBzCMsvJlNQ5yyuy9TN+7B9DUYhcBjyohOc/oA4Dd0Ji/XLqwowYtUkvsuYnIQpQerAAN69tavfC
KaLv1Xca9ZG6xVZcgL0plAEY20rO7eicaQiXdKnfYRyyyvMW1WRVTA2XF79/jFEn8ePAp0EDb0XW
d/X8lZeWw2tyCjWOCHqRRtrtcdV6iAZurR2KdgMO/3C6yfgA6pyfJbrr5/oK9ejInWQqyePl+ZcS
gf0wvnysz3jCn6NBtq9LClkiMsNkB4G+EYXepkKxDw0vplCQzObdMaWA2R8npX8akLVIK27j1c1l
zsqYbBoGWd7FyaJXaMYq3QQJJ/kwIhfbQ8wyCgMwZxhVeQMxpBLVyotAbUN9p0/c5qJZLHK2AtUq
eOGX/1gYElk/ZKaVECHOrHhDBIRZ7IOJseTmn/NgOdQoeK/1aGagmJ+FUuMMH/uM8k3fnMubotG0
Ryco9AS2QR/V4SI0LeuHCUH6YIK0LvkTIdhfjfSvDKu3YqO2yYPMKDfjySe40TYkirRT5IVu/8pI
NpZMe8CVuhCJ0tm7QgQa0FK90Gd176H4jeKbeg2yLJah5vvDe+xW6/8VQoKn9AfYUlO/WQqPiA+F
Tt+uxhR3URAZ3eZZgHNQYuJFq4pzM+pPGtjIL0qH7o2yHWo5iBUfo7tujC45K68xHZFoM26HeWs9
gAyWYTv/RVYCX38ozQ/C2SwdLfYCOGVpVHTEWu2+pI0Karxp9L919xhIRJEAM1V8jcUn08YcXuR7
IMF51bIB+VWFZoJ4HmYtwMgpZ7lh1HegS+95YZmn2feIi1A9+X1WicDBDxxi5ofxkB+YzRaJ3GqO
bfCNIvBxcbPX90ZLQLCU+8YiaJEmj06b4mre72ZNjKH+aaY9F9p1K3tni9pAl/mlDwjIdTlBUH1N
365OEKmQ18UJQtytASRhAzUr/+yv/ZmmP9fUI6Tl47qW74xyOS8fH2R9KKuqhMPx0d71Z/fXxxpA
/m4p739/2BVWUk00O1d9BktArvcfyFfYg9jyMtwtbuyIm8bJyRdF92g06+weLsUjC5s+HeDRX7uX
s+c6NEpWyrHMf2lbXPCxJH9aDbAQONkpBrGKtFqGwhIWrf4pA78Kb7u3fXFVMqoWo51FX9PxoRRM
gnjQ+rM3v2bbBWEXqZW23zYd2knTDo61bUbSBWvlpQid0f4JjvQtgqgWCPbC4iY5ENEuGTpHPqgj
pRk9WA1Y0x0BCFtpMQqQBUZT4SpzdZtdxE7XQjBXy/3mqy7x9AYJlJ5vdGvrP2Yoedq69yW1JizR
Bv6W3hda76TQzt9eOOBrq6GL72ZXj8axdWIKgHYY9ES1oqOVFqEpjhgejv7xuz9ySXTaSePoUndA
RH/D0bANBy0D2+xMbzFhi3hH+nyoGWQU5io/fXOUZ92x6nT/63lPBvMwj53g2tQmw6C6/1NY70uE
kZDizq62jOjATsDsc8IhihG78dB8fGX3gQUuLL91/fD9DEArMV60xe+Dx7wW++TJrWGFCvP1hoOU
f/vktju9DcpR7Ofm+F2U7Ew1P9/mgXLGNW3HuLw3/WlTeJECilIMQw/iXefwowXcYPPRfZKe1gHr
yNA7yXmZNf6h88WeNmL/BBUhRFWHaiHMjLCKrzBQd8cpDw8vFmQlfxZNQBt1kV5rWa8Ggg+3GQQ6
qBvm+NBE65GPMgFlUlST8a6eZETgWgMm6dMgJ3mzLwvXutlsct13dxoAYLvfT0nPWZpM+rXUjnF8
WfkbpFL0HbxgOS6MaSH9GpVncnfDndl2oPlaBcXlVWKA3EifVXh31CN4PwG9R0TbRa8K/0lLn46E
7eOrN+f6ZaEgk9mWdZ1qEH3IvkSjQOgPFCMygI08EZ6NhSztnZYyroIPLmIdspEksbjFj7gC0Xdw
Sw3/5+yX59g9TESCXUruEXOXKWY+fD0JWJ2x28njnu53zhMcNE84pxnfVxcWwzafHvyzQBwIFPJB
ZMbFLQbypGk7b1NXyvMGd/JZvU8s8a/0H/fLHC7cW9QtjRr5tGpcYzcQGQtxzFdpTOLQ08Zyy11B
tshwpn8uBEULtSncfAT/ccvR5bB8eAG9mt3nD+vdh4esyXEdlZghWtZVgGiQrAcW1rwRegx+zYlI
j2eCNtgPPcSIZBdq0Tq0sX7FuSwRxPe9wG2YL/edTifBvCgDqWerG/TCdGlldpHYaw3IbsVujV2C
Y1h2WQZ0bKXCCNpZ3dJJxn346QGHMxzaq1esCm2WrrRY7n7m0EwaGmoL0wIHpKxmTlIs2SBrrvVC
TBayd/lnJDlEbzYbRbNTKPAUbvQdWH3YvY5tgMEWFcNwaCFhGmE54IFJA3qqPyhD1xWJnrkC+iXy
FcqZ4xlyAon/5ujOlT/M802R7kmEmwn7czBUc2Wk/BKyK7n9i0xDddlFQtwt+f5b1PRDZZKL2s72
N0xRdZsNK5NXv59eMUpRHmVNEpdlO0Ee/FECXX2iJrYeNhJHUVQDgY5cIcirHu1Mrz1Dop81cSLu
kAVqQuc7LHVZe/EMYqihTQlDhTqhMz32FOfkVfPOWtRJiAnf8LoZJt0Sy3dm1F/HkhJMqsKagrBq
+ejaTpOJo1KzddeOM+bUhqBObb+Ulr2MCkHXw7JAUwe0k72n9S/KmeNrpbN/jO+jsFCIXCUQAkev
CeCTQd9brk9iuibfBZTwxkeA1zC/0UklHWy/V6iBu8DH/2FVRpcxnA/sS5xmXT36Wt9BkIUFiPfY
BNP+Ns+svynEPxI5Cejk7ZLrZ4A3unDWsgjamX0h2/lS0NJWDkUVb4TH27JDKJXmjMTfNd3bqfK2
LmKnR1EfyxSeS4QnC5u01XMLadI570ymdzm44tIqvp5MTjJzRrJk+X6L2z/5uiU9V8rl8TzPi73A
pnTH3WGHmOjlmgWXGzyCLgnj4cRI2XGvGBPK1yAnO5j2xcXHcsaZAoo1u0AnZMgh4FPjKaX8r1V6
JQ1QmONoTePy2flvplb9Z4K9XJXU5GLytxJiF+5vPUgnLrLni0SMyAAHPOBUVSOaU9trC29VDhh+
RTz5//+UWrYB7fk8s1GMOEFHSCr56u3yketnEBRbim2v983GdjG8TNaKHNc8FeYEWSv8AFMmKXXT
u9hK/8z+Aorppua11xtxwjKLxwkjRuSaNsAoPH0x2YgnfJnw1om2yvTEL4VSGuqEw/yCZjzrYOfD
360ev5L/P5kPilRmrd1rtg5MlglJ3VNI1S/yjg4jBKJz11Z6kNh7cIm01NyYLpeRua48FsSFSSwT
pEg1kdE63a5M7r978PJcNy7ZOuzB9gTr4kwLDqCdRnIHQZFlJ/OcPzeLCYd7C/SiuINWuXpNR8O6
5BZbeV0ayQI/UyO5wgve+p3UFR0MUGn+osiGTTqcQJ22Gn0liDWpRY8DglM2b4CNwg0tK1WxdMEb
WOxiLKaeJ23Ra02+NvCyMlY0y98Twhijq//Pb0hLEOEzhw8WCs4qWE0XjrpOrZ9s0gbx8pVdEKXa
IabhQmuatYvw8VSEr4P6BKNCRWrQwEkg1U139pXbp0vom6Bck7yHCW7lp/L76xZbQ0EK745EZGV8
QiZF4+jaFEmGaVzlCt6jZUqVFC4ISBhbgG5iizvP8yN9JsciYXjrDrIeV2qG/DnqW5ff9lRtTdkW
KOd2kEbMhCVmAoIWg1fei5e8t1yV/OXxgtYitszN7rHEZd+niuv5RW1sQT22pMnfhpl7KZphiGwX
CJ4KB+jm9ELoEc6S0x7iRievvZ2mPVN2fIvor03KiwQTpAM0FYZ7J8WNnjFKczP8qoR3xBsvQ8Dm
adL6mMOPjwTKe0ZIf+/qdCN7TUdhePtyiEWfugZa2dlNfG300cknLpva5sBy7OxowJvEP+5BWz5N
W8WMNBISmJdORocxJPkjnyXyHV/0zwzdXTWUZlnRBIZYBAAIM47GJly4IZXiqM2+LvZFsyVcBQhk
s1kMaEFaeCqZwmlq0pQCCICqhuM1JfjUKKQaRd/lLPuJtTZPszRlrDnAMiaLasduL71elzJ+2n8Q
yiJ2bTtFiOQ8Q67Tj9PouQqzGpY14dyYFd6N5/bTNihA4ooXBJbzuJ85vB9dmbOEmfiXEHVPzeI5
6rCYgQ4Q1wGfzC3YZrkLsPRxh022ilLHn/iQhnR5xLxArHo+7IZW7u+r2KeNgRC7tXjFVmNqj7oJ
ypb4JgNTdtuZ9aZ2dhnAo7+uwvmgrltF0rb7Z0djS15sxacFSS8xPLU8GM4KHEX8Rp5k/KRvF/op
HAjw5bCn5e5iR29/dJhVkUlxIeCVLFXvs/Bvn048+MRhrtDbk+J/43N+GgMBFzBJwosCaSnsjBY8
arLzQ2FkvNl8bY73HN4oKE+FyTfqThDAy85sDtACDbjfeAH0hjSB5aD8LP1B1BATNvIe9n5NlOX2
uiumK/CQ5j6aPEqkN1rRxPIGOFz/hCtN1TiQML2QYGLWNb4Ezq49F598jSK79uTuigKENTD2hHIv
ZmnIEikPnzKvlUkQNu4uVYNJxiuAtmTSIvTtijFRGdyVGiBl9+wOUj/LXsT+BaNDKeSlhNDNVTcF
EBSgJ8/KZqyocWfHQH4KIpV5bef7KpBgxYhunHOcAe3LgzOU02S/8EKzIzV7O8iaYSeG09Ks4C4m
DtAd9H/QfXRMWFt2oZi1pwKi6f7f2WrZ93pE6kvuVCTMatADc0mvGjqWO/yRAAsUntHTH5Kp+umA
APAPedBVErdxhE1GhQhB46VY3WIofRaL5SlpuZ91HxHlYVk9uaJr4El0y+6LKyifr/b+Jl8wlVZ9
YDhtgtFZO6Zkx867TgMhSFkmtWmDP5cqoJLxHs0BAgm7ZFFNUXkVgy9heoUC1rIeN4Ze5EgY46vF
Sbg7CxDKcodw4g2Nsr9fz/U77QC5JAgVIv/AODbIt94h54kUXwtkxAGbX5eekIGx7Br2tQkm89lg
CTQzDqVzTsv3VE1bl/QdVM+Hf1fNiDpXdb5Xly6BHB63WrTZ4TcmON8YEt2/fXqELr00XjndGBpS
/4SlAsHgeOZkCEF4B/K8G80hX/2hoCj4u3DnvpvCXpOCaCGD0cP3IlYho7EFLjCmCPiEXzhDcjfJ
v8VpVORxLg+CWcHM4HRefYoBUTfsdvWTf65YZ9ORO6d5y/R5ZxIXR3xJSCXQVX+USbo4mLOLosfx
FvYdid570lCaxtmpaJczHL+Htdf8L25qxgGH1VG7vnJcHcPa2o/WwreVU7FsuNNh8MmVlvw6Fz/G
kLic3Da8iunPz2eqGwene2D30Z8/RUWWY9MYtzEEkLYZMJSNCFPco3PFanOrRPoKHXErCK4s/DCr
pPMG5kHUbUBzxAd3dViKTNpydr2nREQhVdxaohs+/moDJILZ4vgZJ5T8SwZWdMRxv59YlRfEHMpD
tzFWY2qd3MbKjbqrT60+otN8gnSaFsqt2jUsWxkzyWGrsp8+vK3JD+C3yQOuBdDusTS5JTnMLssi
6EbnRj5yqVAoSNpChEASA5UuRv58saeI5A5WeL7b4L5VxbOyfXziFNufmzyaJX+MdtiUJ2KMJo7S
9/ChJS3fwTeoie9chkzrsCh7Dmp9M9uNAF1HCpVgoPf04rMmO4aSvhePW2V8WjHG58fEBkEdQrTe
5aZ4d3BszvztUJP+qDwGLgdjnMfugRmXdQej0QZb0mQSDf9P7Uw/x/1AXLjfGVeHcOBLTD9E6czr
oM9wMtPYXJ8wNcpAuA35QBbfEAG9EraYtTs8LrWT836EV5S45aQy13M5XICKHD2unauzyGh779Hq
ZrqwG3xmEAwiQ1uhMe8Ft7S5YUit/CIlC9+zIKgIneXK9VEC0lxJGh/Bx4js7VYs0OxUJq1OV1jm
Yf96zwygmk6amXrU0d/Di0v5sl4gwwOHtdSGRPbZSmYY8r0ac29624By+uNsbd+JYxuv1vUkycOt
SprRJE4t+CMGjeji8zjIgJ3s0LnXRm4oky3Vqb+hZyMw97hc7pTFQYds5XUfyJt/EGd2BxyjMlUz
nSKxeEEF12MIo2hvQg7HF2XTpXJpjLTdNqQEov42T/B8un75PoW/pJRQKOzqlwSWXKAELwQKrpdH
3n4+DONCuccpitSQ1ojr6u2Ao28+UFE9BIou2TYjdzLmwmiL8rHS/GYXhrbDA23Nij6zhlVpsPzP
IcPsXUbVHDD6QwRtqav3A/z68qgcsGy5rxXEwyyfPdbHkRGIJ4KJAjt/nkJvJpoY0qjXXcMF1ezr
Yd/ux+wyB81T4b2zT2Q2BOV/NitdL15ACvzgudpTV39/JV7eNiTHnfCKJ6imyx4Mle4shl+OP/cA
Z08NxJS/QtyHSrnVwy8KhKroYM31/hMHLXxFE9REU+uOeqZYq764Rx/zOqheqiXOLSmOxG6ujXmX
oa3FfCxSVcBDYg75us85uSANnHh/ep12k7Vk2PpOM/PeaxMUccpTIBBqZUGAh7FHlEFF8YdvnXMf
FobUhE8NTj6U8VNnyXTnDsAEKlkFX3NGORSKRLtWUB0AH9ZXPv6qHch/bwiqTvme6Q5TxfaWr9wr
CTRuAHN32HLsTAfM6AMf+iWYsKL6gGbulbBKvYc5FlFhyD4xHY2H9RVEjuvmF8oq4SsBf/PLD0wF
ouq3N21CkPAzDmIyrwmRggfGBbEZ1JHGTnOVnEwET9Vn+m36DGypQTv0eiF9FZ1AJkIxXDEEjUYz
9SbDtFajei56iqMmtATYlls5f+SkpwX0KET9o5hqSoh+fk2WBXYv/arCa5T4Y+X3crR5OsWFp9iN
HuDOtWHceFWF6xBM3oixtLsIBHJtLRYPDShNxJ51UGfqiDsIcVkk0GCTyQUG2kBSIX5iA0aJE+Vn
UIDiROUfmZ/0dQyqFNUzS2cD0a8cgbMxn0ylzWAwtYmqLlHB4D2JJtJ0whzkZzrwJxA0uI1Sw5To
cwPcwe7CZ5+IVl0ngvfkN8JYm8XE6+cr9qmgPgJp9extyqb83hAQvOtbvFl5cPGDgpRyS4aai2n5
sJ37My79pBV+OjrHTu2VIzbzI1zt8pHbTZt2rQwjerCq843AVQC2nOvnqu5c/i6DAfRYdQyCXy/m
v+fNS4gvu6e5gU3BXN3du/zjjiqQJRrD9gVgHt3R8HswJri4Q2sRHMOq5awiAUP6UpFUJ355gbnE
r23E0wMUm372lo/2KMjbo6W2m/WX7YQ7t5WXUJVn3X9dSbuCgMzB7hDNb9Up6nWZT3L4Xes1rIyt
HzOowpJg5TuJiyK9XLqEPEpLmT3lOfU6wC+OZ5xHNDn3FMzGs09ofINu6Nue9uZ4IjLMVYXHHQlQ
S6Gab6w0XfjTVeHrlbIpPv4kddJuhGwTrpFf9LwhFeVQ88MXBteCUzWrrHfr/MUtiiDbURUdhQOu
ZFDIthNErBzHvM82KLiQxr+X8MwOfY1RNV3VeITGUIx883+v5ixa9v7GiSZCMv5+H6HKejablIEQ
6AfTv+zC/43JpyjbtyF3QSj2DU7l/XzPJ+oKNPlB7Fpt9pniYCrmQpwx9BNb70dnP/H2JdZLrdPK
aUhaoE6RLK9vpOzg7t9d5MGl5YWlzsampvnDp4MvkP025VImaWC1AwYJLVmnlGgVJLwk1yF3xRdw
TvM0IHasdz4qxPDXBojW5pY8G0O1B/p5B9cOjJbn9TvfoCgYLr8xwHFPWpuHSNN+Yp5o147IrojH
VZIZdliIuSRU+ukMrFCcrUHq7SztvD+tiaeIgu8WGU49wU1YbuazoEkj7rI4Fh7nCMW7ozV4ar4P
wN7AmCVxGCVMyUbRKXar9ei0wf0Bs34EtVXE8HAun0QblDeT9PlM8SweqwZJGwOFebFO5VgiSXOa
Yt4zgpF37AzKRnn6qXxizQ5lsCm4IO74g06Klc5VslEdhi7LZ6QponALnUdHFChouj35FMY1sWV1
TAIYpsRG5GQx0tuFxHUYYo9hCTCMvWig1AwBu+gqaXiuGAkc3rzrtidIrDQJhMVS1Y+R+Fzk5kyg
/ol2Dykxj5+MF+FPlwMBBx9lWTk50NmxJgOZDCm+pLNat0hTED81+DpiYAhiwOq8rGeMkvEDSc8a
ebmrAyQg/b0lRfT0+6EiPa/SdSD/PCzpgk0mAEMG30clsH7wZWF4iXtGq+jr3qVpJ8vsHnQlCNLS
GtOm5Bq5doSYkhXOtSb7jy0wypY1mfT2MOqiC6S2Unxv0pSnve9Z2hhbVyARgXCHqxhMnb95lo4P
16hzJhQHv0baNZ+eEYbfv6/cCV8VRpIgMhsSecgAr33ct0NTgY6J8VRcv0y9ySaVmWdJHWRvOVs7
CYCqv/y/gzIw35CSiuG7LnuKQCw60ds6XSwpe50jBbCgu034ALQVnj5hHFDy8GfP60X7XCaWgN7C
zFLX1ewIr6r/hERCAiWKWeq03kFONfoFbsWfelPFJcnedlDOAMLRVF4DJtgNeH+kv/aDGd+VgNny
Zoy6Pvo5rZJJLlyaKg+VHM6PTGMU0hZumBWPD75t2QujZBKemO1LIPTtCNTd+pWmxAHrU2zGz9ZD
dShQhNToSBLO+snAkp57AYjNtAFhjmSekpW6PUNqkXJvxhNKW6lOSStcVBhjLZADjQHuWacnOAkk
puxsFtfbt4a2zPtdDXQ65m0CKG6EEgUk+K4EP0g/CgyTWEmD3sxmBcYOmSlyIY7IV2MmnoqrCqAH
0zRDF2+80TMu/BvAtKbkVkz0QfY/Pb7/Jw705Ojmo9ztXYSDng06whgw+1g39wr4+6t6+oGef54i
zB/jQAjh31g4jkjbJmwL+UamwlM03PjUm999Hi8SmpwEuqx7TdX/qFFeWQzVBrmTHYazuNhzIB6h
icamnnpfQpJ2FqgY7ItcBH8r+Sp1aFPVe3enI+9YOJMDwYxweqTi2W+RUOZxhqQ+wfa8KEbV24cs
KbAd3KRQd4PNOPjq13AbR1uU+UC1UPB1+KOrqyXkLEppT2DcuzZuzrd138fGxjn3t2w2THjmYILt
DYQgun9VrvE8ROBSaEs7IWoBHAkBO5Y0d1ZLdAct9KaGI3kBGYe7MR4KxzDJ0ab6yAwJUWAmJwm+
QlrgdRfjXD4HHqyv1yz8hwyaNVrREb5h3lDGDFSCALIWGOhMg+mIwjMF/PcYz38aNx8gkoW2Fje8
+/IsT1PTckR/qwCPfOx/i4BfEEtgrrUbMWkzZwu7x+Eeyuw0b0y7J2BI/C2SCAkO436ZnvbLvpfV
dQMHowgMXhPgVNUWpiGiRXnTbYSAxzReAR3ooZtduHXJk+ntmT9zQS04ODm0ab6EasRCY06pEQJS
exogCaTJdLMgF2gmwoWMb60qdgrmWRDHjXkmRBPemNBUhoZ/I4gJifzQhNNBrpXXBzeNE+B8YiJ9
FpN3XLwIyjArgjiarSCw9A5FgiZJEMYccDYQPC68M0+HkndRXZB5GwNydmRl+TwydBjekjBNn1cJ
Ip+UMnueSp6OHOxP5QSKtnrUXVjtLwjMXvpKd0jgp3QTvSDRz0MOaeyAuw5yjLOItl6Y2MsHPg3I
gC9VQxa3O7h7dOuNTQmdI9dt2p0ewgjl2xLGmYt4uoT4L07joJOhJVQ1QCU4FwIPTGbt0ZHnv8Wb
0OeQ80rNVVgYcXZrwzmiGwzGATj+4AGdHGLc/HqFL2q3SbEur1o+BR4LGm2C166BlTv90HpfaxXZ
TmGx/DT7+/7UKRj4mvSa4DxxDO3YGa5G+zrFkqok4XSw9LLpsAOMm1aBS9KA5pXOShAeGIlekv3f
MMUztT0X7VyxhmI5N2XNrhkEpj6PlkvdImA8liyR8QV/ZsvB6oUu5wnTa5TRkzzzx84XGIJClVg7
RqS5MxIr+AxMPvOWzA0zQpDy2C3mlMamhrcFzX0IpoI8ucb0K68FN78zL7OFV/xCjcF4nL5+7qGY
nsl4wYntJ+M8FOo0ea5k53tD216sokxB3WNOCKC38KAp8PPomZS8Oz6J3ckNKw2jvsIKuoNzBWXO
SoNv+B3nLSjrwsOo8tT7pnNza+EPUnk8Zo1gJ4tpKR+QdM/1a5Q+HgNvwfdzJaEx+r//K8AB55Yh
mobzbFNAwOTXwJLF3cEzzLEd+a9rrUE+Yl++7ZPI5Q/RgfdKdQRMPuz6yn5kzjh5YKmL7pnm2GH2
TjgIWKz8p2/EzZAIwL7Vv0DPkUOrN6Kvgw90gF21eknR2hiWy/BWltmwPSIqN2PWGLIaWM3RuFou
ziSyJg09LNa6euJBIaahlJlLkcbNdyqMyXGL9OFqcABNpthqUp9p/U30qzOqoL+o4PS59xkIrThX
0NrJY3WL9sc6o1JwYnFSO5AthFwhVb/Fj6Q3fG4s7Iso3W6PHM57CcqpCosHvhtnPxDMiPaec3dP
LnFWSTnpQIhlD9+OV2MZFRUEiEfS1oORXAhs0jAxdqZcwhqpN0ZpXj32XrWBbPcIE8/8rFKzS+aH
8Laekcm0k9U4n2d3xSyc7lRH8A1Lk3twG31TAzm8DZdTblffG3bY4g7/5DPkITnRiVGlNAdTjDuf
39RVE0QFaccY42P3NezqWpX6jZ6PVLTMz54r9f1IgzosfJva0Dr45cuLwOu5tZ1woObNoWshRrbn
Q1YM6i8pDR/9cRsPxw1pfeUL7T3YltZMznuoZoslvSGPUfss9zlp/1ZAH29aDFvLaYoDeZWOHkXt
Iu8qha0inhzQrFdn2qxO7So1AbZdIY3Qo+7gRk+7opxTBICS76zSB63bJ8vS02f6LAOJtkF0IukD
u4Rpf+tC9hq4FaHV84L7QjAvwMd3rTET1/5Da9ihJqNziNcal2zWwK0NncZ9+LY+moPoOTuRlMys
YD8LaLcL/sXPfQSAR1/AoDB8oDyID4AljxnHnRlPyMAkCwK8wYuVq3KKXO6v0QwYLArOmqmSXJAI
LA62QoDnIk1eMqu2IFv03e803zdVGMol4AF6fT2gBvi/1YoOP24bW8OR4N4FsRn6oJzl9hIedlOy
vUZ3CKGWIBt/+cFG748tKkUtmY2D/wTz5qU08/B+s417t/UtdhSeWSk5RqM9kUX8uVO4s20snWGr
zwJaGaARHfF77iDA+kOyHsqWG9f2vnKNBAki3tBHYz2/U/YpNV9tXmp5FTMpnhgYpM5EOUEOhY5u
iFB+W3RR7pYgoSc4940kY8PXmub9X05mrCWdYTMp+Deb+FF0T3VjKWbUnOry1cz1gsZ3r7fSOjDc
5Lfhpfi2xuZ/EX9YQGzwMtByJqiBTzZOUG1+eU72zDm83LbDRqmD/XOzZy5kmntkpuMHfkDORf5o
Ubxcla0KnUz+s7rDPAHuL6qaipLCr8nFYz8a/OhYEUGmj4sWK/ZPyoPrHD8vdGnEIile3BGD4/f1
VwTfD2OL5cJyqf73qPYxbHLXdD5rYbX9X4i3GWZWQYv6fsKid7XJ3bufMVaVfUJ3NA/AZd3h3u7I
NBAVcisjUXLGCrcNnwfAeHDXay0ZLh4HXtbRcBlKLYyIWgc6lucI3HRKSFEEUyY5ObPGljIsCE+E
YLd3PFSo/9aD8adpPSWxkN2JebyNCx3m+Sb9R0XCWPQjKxqRAMHxFFTA0ufW6uPKqsqwU5kXarcU
/1EmdlR/Td8iibzWXig/vg1knV7AfLLajQYgDFJ6TDbqu3IfXIS78BYuUWt06MJw2Yq01obhdiZ5
gg1VmtXr/7WfRjeIslNHQCgrnc6Pwm+TVrT+LyxY4L9OvHDPBQdyfvL5FkMbMQIY+kcIi4Jm0bMn
Fg5VlCbx8GCVy0xNf+CGirV7MKmoPUEctoK4G+TuhB6JqFbdosvLvrFRI9ACZWUDEp8PQHpXicSw
wkMJclKxTQGUpF3agUuhae2Whi1Sm3dEEFugO4/dzbjCn3Gd8BQk9l7HgXIm6s058shl6WdzJddO
bhQnRLCit8Q8r/yjfwNFuV7elqSwypVanx5a8ZsL9oXfndwhZb8uv93ZwbPz6p5nIUvr9l7HiXoi
x5HWl9oxC57+3rjRxv3LqNaNjh9DdbLZP7JD2ILJOrG36NzIGGlckPzrCIAbUd8FmLDK02/dRf2Z
rWMKViMgdBwDu4tzZrM2DZeGQTgWGJKpOkNPmtM/oJx9piKxybhmaNaU70Hv+ETZDRIhjj/gRIcN
iySQ0XVFd2XiVehnvKxfp6ykOX/p/D6kBfHQ4tEKsExkzdG5fvo7ZHC7JIzm0ixSBoJIfr2Qvimh
ghAzoGpoY8hj3T0WxcaLD3dk0T2iWFfMmTBxFZAaOmzBlfPYD0FBckyANaP+whuCzlbE7Nstb0NT
JTXdnbC0xIA6xG/040e53MYc4bE/rCvY7x2xL/l0yZji3bOIiRimCjhom2P0GXcQgmNSjasr3FVq
ebE9Dopz8U/MWVH8IRr+adfuCTu9myqLt8tF5MI3xV4bVHPDiUHydm4A9C6awx1lw0vahmIfp4pq
3M2aw3F6MkWqP5KeXhrBQtTZXZ/RN82favU2HZbGMszSs3Bx9cRZJ+/e2SSnkf/f3qquY2gGaxiT
lFdEq0J3z+CV7reVNykSARF5bLmFtabWtUTO+N0kbYkX+OajaOiCqbybVuvvapkzdXO6mJAil1Ld
ZbDHPy0L+ZUEUHEGxEPNhYZrfek3kysq3AzcBdMdoPeWEa5Nf6HyvAsgzfZ25X98fUsJS+h8o2Ya
xww93AVa4PNvLvSBFBnWG3Gwwomr4MGFdjH8g+EGZ/7FCOq5fkI7yOY8CPJv6dk3SEM43haYs94j
bzQvgKbvRl3c9l2CDHOcIW/1/K5lCs4pC6JjI0Rgf7Di171xWtxewjSm0sb9JT3WGCLjy+Xa8K96
WBVd4WyV6y5JNyhAHG5QbR76J3/Jf4EDeMn3U8+N/evl9Cyko42dOTR7WCP+zScfRHlckhaBexzP
o9FLZsxsC71dj35p2U0OVhaumoUmos9X5/BX9ol1Hzg10akZQBwUVhawXUqgo8uj8juW/7JsSJGx
1koTW2vTcPlq7IUgqS0OXJEw2jI9CNcXJD9UDGe7WECtcLPmzsZIXScViITB90gpW3cV1Saf1dMd
8oRNbFJHo27Zk3ukICv5IfpCcdYQz8BvSsVTb8ay16TkCiXMBeY4E9jEvksR+gjVD5sMORTVG2xn
zIiPkkjVbY2yg9tw60NdzoE5pX1ZYEeBunfsma9LOYHtWyJosmoqnIPO903U9HhjS9UnXETOCHLE
r6Kr8Ja15YrtjWmkEyHaH2zmTefpgPrHeOw1N/rJlJ7WMLrmUKD6vDDz4EDTcyySJUQC1F2O7ych
XKbC+FG5+bkeacMJXAoMMiJyM2r45FAqO+/C+HchX/pW27KQb3WZjXv6/uMlj0GzAYyyegxhp0HB
PDlEETIYgcOe1nXO5LcCQcKMReY9pzuX1rHRNUT7shejtx8Y4p+li2gXkD/IiUlKBikRcETWGrFq
/qA486dWDI/4AgPb7Yl5Ju/gX7MDBjIi0k/+xQ4zzbT5pO5OG7msKhjsqe5cT0gsv749fvKVJIZt
dIGBy1s9B97ljKV0faKo1qz0Ll1JwWe7pL/GSNgSB3iTSb/VvaYSNnuiwqPdQSS7BI801/iOhOgq
85j5oSqy2KHPbga+9Pf6G5sgnUVZlK2EDR5qfmZTP00SDJyjFNx01XkM95bZM3W3X4F/ySGvIlJG
dxcAgxK+G3+iuWU9zLsH9xWJ7IPd3gGtvbZu81CT/P+UojAnFdSsHUOh5X5GEntXGl8MEMCzyeDR
r5EngbesPGbNM1dz2NLZ9R4HZNGRZgnNY/gm0kt0ak4MTRWinthd3E78xDboW8b0iGYcxqPuZHeS
M2p/JRfc5igNYEne2MH+pdom2dMKWN7wHK/+RJb30RXXApAymCU/4awCOSyQF3bBj/49rfeSh6NT
6S7uMu5Lmz+HiZeU0ub12Uj+yxZKRgQj80Q7VPTE8iZERxU4/BApffQ6H1sQPrrozCr8LmIuoTBR
RLE17wdZ1ZaPfhyh/bqxG2EEAeszP+HRYh3nJ2tr0nLIQ/l8Bb+/r4TyisMmPdP6IRVorsA+FA9z
CPXyz39hkgduPGw/TQKjhqD2zT2KCI8WDaBbYPTEbLxsuqJaTK5UdujyF/i1vUEMEmdvR6SAw1/V
0Itlj+Mp6lT4+fQgPQLpy8dYbFc5UnC7VD4hOWa7xpNOFq1wR3ErcluXF/7bS/1zLSPkjHF3pjsM
TH//N32or66wfR5bz4G0wZecNQW3opu3rDswoDPLvsiRGCyq49rJbUPlwSVsg21lJ9lFIFSqBc0q
kZsNyJxqPtCzH5IC8fRgQWJ43Fu2W6VRm+7bn0c2eT/5DCbfbhtfddqrbwp/9Y4AvVndzZvv4rIx
A0HZNfbuk7qVcGBbKXPt6OCoB43QoLae1C/DDxiubq+aPukVSkWHVGNeIx47zQvhfYXpBByvcHJX
NT07Pq+rGvgkXksOI7GYlQusmeTfXtj4f39aPPv0dkH9NNSNN2S4OBvicU6sa1y/oWlXYNANEOwl
gI2UwJNjPUEjYYxng92tNy9hKdk87RcsFxNpMif9djyQ5uoM/Cx8bx5lN+/KvTh3FKoIh0wJZYBr
WvM0krxoLsE2EH/aa4/fcUa1Ckq7val7zZ9HJp/sqEH9EZ0JSBBTiLj83303A3kcOWkJAwxr6rbD
PZNr0qaeEn012OW/Skv/2oVJWhhxGUhi34XwNm2dKLaD+taJ9TgXR+Suw6xvO2FnVd3UzEg6HBAT
f/OzK+e/yM3+wpc1NfRq1DYOi3m05o7ekwE/M3Y70RYkOvWJ9MoiVoyGTTEXiRsbewfoJ4VJ9wPL
VVBdtOOpCR6QXyBUtB7By0CNq3ANYwdRkVxlhYzp977q45NCrrsvrEOM3aiHsdkKixnyE+lkYkof
A6Mjm4MYw4/Fe0PE0jXuv0oTY67uK5ctSygC0hE6KQCfgEi31jeJ1FSIs+oDexm7iLLbwd2AxAkp
tpNDWFhf6JG9dV627FSMFlVlWf5JjPzEad1RDqiGAvkPGHMcFc+UFQp0wR/V7+huSbQkxQRWtqzO
x2lTvuvuSYbkJC1FQd8ZpyVXPTckX0kMT3nHluEHVK32rcP9p+i0X9RxGzHy6Yq5I0CqjFEJxzHq
6gotSWrCcM1/db/2GHWf2NC57yL9Si4FbD2LICOVEmhTsds51ENdSvUfgCkOsInCehMtBOERXY/4
4edvo/M7WeGSOe7huP/pJKPJHmW9NpyRZgVwbIxkkGw8umGntkqK6+rZI4xWo2V37U0tLfH+RdBt
KLBBv8YB8I7G17NkAOV5CM/pqhsCr8wvmfHQ+nMLRVev4Tr3vlDD6eaC2mxULLHo6rwC5n2VvWmW
ppm2QkxOsFIAFBMIqL5fc6KJXF7ZXll0geEO9r8v95DF+vRUk6Z16mPbOi90sJLByE7ZuPSYnCj7
Ks6tuVABwgZQku2sPixhdsEOLS6mC7ygK2XbfM2lKhiikcuMKSAdgkF8n6KOUDBZz4ORTYcaHZRl
yGAYMgg5PV8iMe3t/KDENvusuCucP+z/9cd3Z+VWP4kC157g0CmP8zkixWzYIwVYnEVtuidPBcEv
/d1e149BaPXJ307Ca15XZpAxCc5rE1SrcdAUxyr8c51W0x7pHtejBiixjPn7+AAbj/nea9FE2wxd
XuVqPsWbJzxVor6ZlY701eOpLizQ9PjrZn6hCV+vlXvXe0/E+uWLdauHVtgHwA3i00i2oWOp2JuG
C4/z6zqNe4e22JljXdFVN858FEHlE8HT6hlfFJqfXyJr6V3JAemqMxdW+AvJUe+dJ1esuBu9xQQg
P9BYxnkJQxguQ9R5BBu5+7bsAJxa3BDVrxknqUQ3TMtLfmUDGHj0fC3vSlWh6MpguKLNBG1lOO1b
N9t2ptS5MhdzxEnKx6ObPNdMdbNY28QwnWNKUEnamNr0+VSNzqy3Xw+1E8PoBRvAM/3b/DwjU8cR
6lWLCSYL50jl48AwsJomDYI3IkfLCl6pyRKBHITAVZXYx1Sg7zAeV0iUK7RLt4f35rO68ZGBKKp1
cb3CiXMMLy6NPhSGbfQkYLhEPcSLRzzCymoCi4pfhTVJlU20vEQnFute34pg+JEBE2sST/sOnAlH
DT4csmMHAjw0qH6rUedr3420puEzhWqWa8W/Omgpbi1OH48Ghk2kxHW8KV/XuCEI98oJIf2OkBaL
P4LjDiKzGJCz5sXepi+O+y/WDyGJdMwb6HULr588QuAAHG7sSDnXszdYXhscG7B7gfJTXwy1RTyb
9CPdHjLfzRmlGPegNe/xDCvXXYOqhXYpTdUUdx4EJ/WLiIe4s3DPY6Toi4APUaC1+4kSBe5RVPJ/
6VXFOcg7pRaewu/B7zesbZ+E/wMFxpCYp3tBiV7R/1sFM/749Or4kcdQdzk0ZAuKiEFtlsw0pasi
l3zdNvULsEukuhxiRW46Tt8/1vIviX29ewFv4OkUb8Z0zLMmKcmLvpN6SDTgRLL0xWAODnxU/JAI
lIDs9rrBehgEHGYtGnTPWuHM25wKrJsPj/3bb4vbr8SHQ2ZjgMIOjZ6L5E8mjxK+tMW3pcBeM012
8tkQN7bdDyT5PzuIcSEwHCMuCHijkhmf+mwkMfcjvf6oZ6a4VXrqkJ56wZoHSqJrxkPhbYEY/dD/
sCEzriq9hrnKVfQyG5iRU/rkZtmJ9/TLHHu1AUjdVbRLXOV4EnoKmdJ8UOGb8Vth+z2pJhCktBQ2
yPe8lBuJVBl3R5yEX4ICsVXG2O3wYS1iF8piO9rWgRqle9RNhIFbrAYT3CNW07B+jQk8KDH16M5Y
a8Vl0q4hSAmbWoFuS0wxtjd/tlYIn+gtjmaCfd0fH+lgnCXQurg6/SWEagdkWKzEooOJi98G+axA
dTQi7fnSNNb2G8zUoAW4C/pt2w5JPMAfxbyRkOWqzPqv81tYbLOJQYyHQdg8AdqPIvaUuAgOjX8R
WaczUeSgv/K2tPQK8dgYfv5Mk6AJhqQ47EyI8T+m6rcfDrYraO7qL9L6c87IAjVV840zI/PITFVH
zu6EQCMKGUaziDs9woigH0BiZOkcpxpO7GbmImm6wIKmcSTeGXlzGVP81Jx+Ezuhfi14hUnmJZ8a
2mQ5KIVVsZLGdBnJBN4ebU3ZZWfl2iRY0oe2R5ZAY6iKGR+C7s+6qF1tDVz5+kwfTxJN0HZR73BJ
UupgQzx1kh64nqswAOZQQSk3Xb2xuOdLVV9mqWmhY+WjLLr0qRuWOtuKfJhLhRtI0n7p8ivkpey9
j8oQy8c6uXlEzL59ZiRaU6784+Ak0Wv9cSkdE5S1IMcMMci+7gzPgw2Z+wALXHZC/xXPkckqdtfH
H2H2uMtfhaS1oG6mrZx2R5JKqUZpL/LojXW8vN713P44k2b566xvcOvAUetEZjSzBtCx9plZ8UaN
THmJMPUzNjgu4fleo7hbfDaEFEN12xtxHc1bAHiAbuLrZ9i1bcUD/60v4iCsP9dXwhqy7auJ+dli
Ovm8FD452chYIUtcVleWcU/FRbmWqJ9rU3haylRZrbj3mFr2xhWvRLsZz30UDBCO5jDfyC8cjWwe
nMRzdFbhAWAuWt4FB0B2i/LYaEGqIkTac82y1tvhgKlOJYv0PFNaoTBVPrDLgtxmLbUI98bOqGvv
L5TT5SDscgS4YxW5dmWIR5vx5+vbrDVDLsIXNigH7jHp1Oaa1r1wfijswaFLLmZxAUl9CrHQ5QhA
apsJ1WsV8hYF2ZQIhikftPG2J6b7iUn7CJP75hrrra8CNzkCLxfpA+QA3QqNMB07FM2Ur/3CLYXt
6Yuhob57oxN2L8UgJKazch8RTOlfwBWXmv8SNkqd6aTj1zhP7pU4UFhMrUjU0fzlv5u25DYNBBb6
0yPFb2/a7Ns6/LLBsIZx79kbN7SjnQB/tbKc+13Rj3GUEhVx1Kmm1CC9RsIRtU8h15Tb9Oyx8ILW
VkryHVKozqbFAondSkNBCKAPgFManp/RsRjSNwA7o+IH3oVE/gCpGkziUJTDvQ5nh8GcZf4yFmEd
J0DjLHgn8vPhhs3wsOpWocRYUG1EG12bg1RhfJu5nJBluf9Cnngn4Z8DNZzfZ2guFnI86l5af9Dn
99yoBDQJWEo5afg6WFjygMU4Ih5Vk3YWYTUn4nN5q0gGbxWdFaUUiQ18tyjdbJ0WFKfQ2W232oF0
erse+eBJ/OcEvl+RobcSvfv7Xf24dqAdnGfLtEw5uSYacFaRGEqi8GTZcmrwoaGLGLB0ZSVrj5ZQ
AjFKYtnc/J5JjzeQJh0yZfJrQK+2nx+z5A8B2Bxo/QW9IyvWnBxSsjLYX+KN2vKgTwM7VSgQCdp9
k5aMFU0Sg8UIp/NdnKgVT+d16TF+pTUyt8/I1WFzSQJc6nKrSwjA5Bis3fikr9+MDwXTYOPnT4bI
CWVZrgsbleLaqnbSwhSzULikCjEO3GDsqFaSI9vleFRSPs8WLz8ehB/5+3AjvCzjIF0jA4+HDSva
bU5RQ23ItXq/R4JUcshAi9crnUt7nImR+9vdlhwrMxR4YLKYtBGF/iF0cc53+rQpOt++c6XY3VkI
L1FzAAOD/fQWJySyMTc6VbkdD8XSAQvkKGqqRCv4d8Qq9+bMJOkRqnZQV873MBKaaIxzLVn/jsF8
jjf4BtncdaSiWJuVxZv8gerwwqteQiKcajzuvkfid1lptq5f+oQGHdtH5hfeUvyokog72qz3ZBU7
Gn0mRnTWSIWq1+0rzb23QDqlzZ9mHiRUcKLX/EwLMV04ZdpyQ3/4Vr9/1/8m8ijarIEdxAaKwnss
XsIeyJtKVjrJjRnsUAlpXlZJF7F38Jp49/T7lEp7BJoD9Knk/eIPAa4mRiDd9ZrZk1k/3aUad5Sv
DaAh6hIKlMO0y6/quUZ/IcpvEy044ZenbXyQfeO3BiPcrQCPm1R0WNcVkIJTLrEQ/AxuoXtwZSr3
/iH/6SLgFeBF6Dbq+tbpW1Iqx29GtQiFNS3XOzjMfL57BlcTmYpxbkDC7k7mwM4h7TPocap7ckEV
yh1CGXtgGZxbv1mQqvlxbrvU/QLQlQCPUQGxfCLfddn5jdKQkpfkjY8OJ10HO/mq00HRPjLK3GG0
yToeIkKLS0vUiWZcAjf482yiq/0e3qCaWVEex7S5js3OjPXqd3blL78DbAqJLJlZc2M+EiRx8dJJ
jFxompvMGli7irN1YAYBwAITozVG+iZTd3p+Nk8K7NB49lHKgt9uyq7oiD+ds4Dm3t5sM4xftK3O
s8ysZC/Q5Pd7ZZEAowB5D2WhHF7OTX5p6Wox2iL6OXmt+Fac7U4uhJqgrkBjGJBhEGaotuCxbrDO
bqdX4zCR7Cga/2xzTHe30cicJ+i/kyzWXgliAvWsN4Q05PUR6X/tBEsgA+3NC8siXDTUqbjZDnIt
4ietD3XGHLnDF+Qk+5Nuv+fsXGIJBEDCWg0X3YX4p0k5HA1rojlqSM2xjFLnOHaBk0Z1B3ENisE8
bAD/EecTRnjSMCopsohqUbiyiT5bQ4hMKCVXyzh+uD/BjBqE2zKXRajF2Wx3Lm2qO3w4KpLuOUPi
NxJjp8g/ePdFnHAoCI1kNfOZWq+tc8JeYw/Hp5ZlSPibQpbw0A4D0iU5zpKx4HPXUwxsVZYHyFTY
uOmSHR6r7DjUoD7f5rbQyhzmqWYOUmYH/Ux3HSRHUQmB/XvzWbxRW0F2zMZ8Ta7TXTpA805w84eD
gftAe1b2EXMvkyYVn672qjcITsOdAya6Qxct8WtCas0nqfjnCKaL+yPMkjaGZegQL+5t1tlkEae5
qPTzCmJiozpA0vaFb/RsNfcTbEw4FfaEQeQEv1DXaptc8VPYiwGc6Hd671EoyR0mrpg3y5okyzo3
6T6iO/4xisGjXFuy3ptKST0t0XDioOYlGn5xVTFAfCcmgp9dvX52Nd9o2WThJpqEnBNlphWrMpXe
Ha8AOyrFh9q0rEtL/NNCwZfyRx8jrMyoAET1KzmTsTjamVhuYExKLiEjMApWTMxaBTtM3X7kwQtn
aJ0wm66RYEv2S3OdeFHcyHrk5KEa+wfR03PigKL6ZYfYDBugYi3O7ymqW3YtGMrPrDr9fVY12MhY
jiS3Fd7FmnbYoET0VpHT9poGtI3rUtd0Rz71xx8XKzWYFsA4wGVtkcAOhvKq2+fbvkIwGsuiHVu/
3b16LUhWj8CU0jKhgHLaU+ou5iJ+1o1JwILr8k/ZqgER6VMl0HnFHf6Mz0U92eKV5PnrnIE0Ogtd
MmXWTrTR4aFaUOdWUPKSrv2mKxkLs6lCkqoQueVsvxoQkhNJoltskwANwFNgOqertA6pGehvme5A
sOqQTZ5SknOsAkvZ5SIYDqXTX8+xnsokduJU2WAkne3SUJAETzn5BOrAxCU+kwh2dS6PfzdFFMWt
29wyrkIO6BoyIKhagPOER4/jHZu+99ezwl9RMMRKmr8grluiZr/r5AoUkdm31z9qvK3S0mYwJeXl
jJ5zyNRBLRiPQ3US1bCzv245ogBz07exekYWeIROXDGB0ph4mxdRzh1Oy+Oo7zN7KsLic+RUpH2i
eFrUDU+4LLEJKAhe4t40a7N5tz+T37R6OXWnvFu1KRbGdT1mB9XdRXr8RB2pyIXPbZ/O8E2+Jsm8
0qibWAxpRSnwfUs2ySczSGcZmECQL55EHBV1TJAcuH0KY0+g2zmTO3SA9hyFowjiLtT4WjP/tmb2
mO/mPTrwe2Pkpo+SodwPWE3XlwtUqzDQG1kwp82bbhZ+eT7WWjMDKqS9wpslNUw+QAg+pwcPbCR4
F+sPvj/jgRruwAAo5QSTTL6avNAB2n+Z9qZqUdi4WPlLC4d1s/sNFNsC37T1qyIhIhirxvEt51Xb
PvucWdUdYVqYYmCQTF4DA4vZE8G1YboySKm4HhcQqM9O2BvUAYAbyBm5JiOqap+pCap6hddA4gKr
u6OVLFyLNX9KvXGdejG1ao+u4M5++aoaYtHuaD3ICxNdwj15Nia2xr95pUhsSDiWTWSqTlPizaPE
qZ6hMXZiggCw4tVzRfhUT5qlK0ZtlxPn+oflRV5EjRINj1OFCYMvineIkzC5lCF+/xrwE2TTRQKg
wPeCW/2a5b9KQFVwkIPjJBsui7gAaWFR6wmKxPmi5A1z4HTk0VSSu9/6G5uYIYtUxfHoQGnm3JAl
u2GNpmG0+iGkfp9+rcoDszrs93azqyQ+bl27X1H/2tRUM/70jPdFYMlDcWr13KGXZj/OQGWltMy6
+IM5ArMBxJAuSYCpU0jACSh29m2BddYy+NyvuIf3A3o5VXKx2enKv9j/sdxLTG+o6CuhE9jK+u5q
mq1Ac0EK6opVvjgRsJAOuwf3M/5tNuTyCzZHlosUi4R7kM5pWQh4i17gC96twntLaXE3hHB3ieC7
oA1DLswsGeu32OAAeTj+B5g1TFs5Hi//1XnwPEXImFFi+IMIrfiGTtGPT4hiQ3w1NkPLMb92DFRo
KGqYNmq0dtzI7Bmzt4/L0aYaib57ZyqPJT32JxdY3oMpm+WpVeK/MaShOMeC6Xomvd7ELH7bHt0v
xxfA198jfaosyD9Jh7tYiOiqsIhQZXQ/2Xw6U6Ymod8OYDKDQAQWqhk8t0lMcQblosCSCVpAJSNQ
7/6F6kYjIZaG8vk24vorNvfy/0cbzZHnGD8h6tQQsB2jv9sJui2WoC9ihC3zxkwD8r00Iw0mtlbV
NJq2WCaPL+MHT165LJloSnsEouiej+GtCW6orNHUpbDvxyx6TWqf11OkG75ma9PLl1iQS50tV8XB
/C8oDJKZ8q111w+rRc5eV1NCah1+SbM/8gP+sZnHoaD26By/a5Ps/IH7RpHUX3Rzr4ThbIg3tayf
VvU1xfkr2KWJNuQK3pzgedRBqxnZ+uUWVBm5Aj03K7k3FUTKXVGyPrfywLaKalHo+gKXG946UlO4
UUr942v2k/y2hC1iF3M1x0DI443uY94Ai2PBmygg7WB/wnA9ixXW29FnQalOmtvja3dJXNvS8N2V
qYjhI6frY0IWoL/C1H+ozKj0i1XEWrbYNcSZ34VfmoLyL5Rbs7YKB+Q0Y28fwKxt9M+FecFuDt5M
V3O0o1obBL2GQqOqKuZo0mNsEl25p4jXpiwBSylcwfOno0qBK+znqSPObioVq0qTWhCsaB3lzEDK
VGUXSobBC0jaaya7pEM3+3rLXeCfHGLOCTe2FntfVOTCVeOjxyX31uTNcWCTATW44RLN5DjP1x0I
Lj9Gzk4t3ZwbEzXGWszxEd9vFmLlwrkOtZ5SQoyEku1lwEWsSZTCMbT3Sz1dgn8Ty3CeVkFx9HKl
/qO3W1l9Hjcr7PGIIjq98XDt1fb4Q+/ME/XIWkxnvFUBNM80PksYieBX7jeoXRG5atF1XI57Sxyo
GyOTIbeMHidYJJkNhkeR3uKKXbI0W4MqQaRS1W8cOlAwZ+YJiBIfQynEGu/0iMfqdYrKvpcUAaim
ZP38G57YQ3y3ZHPv4EY/Rz2pTdE8iMjabG8GuBMuoElogk6AkC/Qt8VOxfA97WdoiUCHq5WCO25O
2JyRc+OFxUtJ2DaconKl3z+cu58Ou/veda6aaq149eVUn6LM9A9f7GeN9NmdT3tQEoEctaRpmdDt
/Q7oY3rLxlRh2HMng9egNuKVLm2dj13gokZKDuXoak5dK+mmDdCws7Y+1SK+xuuBeFQagFKdnZ1I
y3wbw6I5MglQoZOgMpgJMZ5lyZpxSETR63126RfC3l+BWoV0MXGSx9g+mlY6R3Qcr66WgCeYKVT5
NGU5FR7i4vFP9XFtycX6ptGZhmjkfeBoTuuax3r6OI1yVbECHTVZWYDgMBdKMWsuKtmPUgeCZXTF
xMfI6lhTUNd4C9b8jLvpGSczm4pxU4OfzQNlpxFsvYeNFr6Q5KmnPI4GoXMSJIUcXLV/l8Mj2rgX
VQVxiC5CqFz4Hwfflxz8SLueA1rjBU3/tBUd8mAAdQJGFHsSePpmJayBPfwQ21XSvFDigPQ/a7hq
oiTfkfiZ93b3RtErjpmIX8eOR8YjjZiD6tryvpokogUJc3aTLxcl6gKgCUxPTEMUidbvKijuh/fn
ac5xp45WyqH3G/heXdKwOAj4VE9q25JbnA+b0CYyLL6s4Y3guiSuXQYoEpvdYV4hANqHvvnssZzL
wuCt/di0jR/RCijP+Q6xH2TRQQqayCTMzT9jgKmfTfcF0TNSgaFmJ/gLGZgD4uvjFdwe8XdfDv36
ohhNP0gMTzliYVzEcSpNBODV1ooemFf4V4MFMtX86UZPUQqopHpaRT/uK0v1mZCZZoGred+DE7+p
Wd/ROagzkRpqRLJ1uN+JikfAPFAh8MJxhc3PeRhvKBN9gdNDePO1C5e675wdpvKduL+VvsSCjJmF
38JPxJpZ4cUpEbUM0Ydee4D7Iln/QNvB/6rfoKm72yVGNITYGuocMABiG45M3d6aLdEiqjjWGf0t
8/0d30Ux3ecEAJ/KExuep0p81Fkw6yw4FlZTbwpQNqmVb0BjZCyvGuls5P6yMK2YQirI2seZ8FXT
0PHLpbfYixCmkrcF8JPrmP2Lz1Cn8Oj/EgUsJ422fncVRAuBsxUcmhTrc3ck9qle/enkFPWgJu3R
twNDphcCg4tewHhbbl2njvRzzKDRB5L0wjUY6onjsO/3dTRE+I0baZm7ZmhpU3761IipvgW/BikQ
wyG55+lE+1y5yXm2tTM/lQxhAyITQ5ZcSEBPgsnvXZNowbre4htfD59BT2vm99GqmZnCdEpjTB7f
vBza8lpgSXa33q+WictwPzEiJqOLdPrNndivKvpUxbJjA2d/xeNa6U8xJy4L9Rc1c0uvwskTFNnq
YkD9HBOh7WsnuXGlNWpj3z51xGr5Fm6F2puLax8SKI50JVu5I2UPoxQTaX/Utc/OwxlZBBfmc30f
pXPzWSSiRO0kJAd1AmEeUjcbYtA65CA6zY01ODboRH9NWZNGyYtTDJCBG6WUmRcFqS0B53CYWy1m
7cxhpepMYnAs5hqrD8KHVjQkoRq1zpy/TGa2GZltH/cGy1AVc1NTAJWVgf3kfigf0rDrVkpe/eLh
dHRukFaa4sU6rdJsZfv0nFMKvXLNzSdwI5rH6xkCjam3Bpd2yYhn+ttKYMAfVpeVBgMniqWhAhgJ
uhrXNSaMo001A/I9T7BRLMzic2HNIdXb5J/P70YZNTDqG9WVAAdtLOdRv48lvjkuqT/i5L7uLBGn
4Y2HMVRXRTgD5omWGH41D5fX8aC6/7dyStJbReYR+wdESAKTMEfFPBK9RtsXqBjN9R9ge0tsKOU1
Sx66l1XJb4V1kzVH6H2BScBLeVEd9dOOds4zyH3xY2M1omWOqV3y3fKxprGVGYJ0F2IJlIQi/mVf
uEIiDq9zyJH8KnRw9i1B9wTQ8wl2InLNBYCcLESpElM3ABhtVIEPMHcb0/MCcTJlTwLRvwTqxUzl
iOU3ew72DzCMAcASwnjE19T+BmlMk5a21EkiXB31hPGuCreeS+ODYNkRyJKI8P4yjbejwWNugZzb
WX4JS2EsEoeJNAfhA8IiyZuqbK+wUfKnKxC5vQ8+Xop1DN0D868RjsGpatdB2nYxkf7aPRryHd5q
kU925DBmuczecpx/Ak3Rg/Bi7FvmYqfUqibu7LerZAnzvwQfU2eMVIbX5/cyLmOcc0PzTV9eGmiS
L3In50zmlIlkddbZjuMG65V81IynS9/URJY0exv3m6EATJFx2EYOiLNNs29sV9bfEU7q8zRuIm7h
qrY3Y3vHpbFu8z6v1zwiGOvKVyC8dZEWP0kkiTVo9e+uCY/R90m1beW3mxf/o9FeG0kyzpUV+tsr
RkUb2lLGMYPZTQPBEYzxF77hu4xSM9Vu5HRf3Ii6bOlu5nDi2jnA58ELc3fi8f8TQKwYlm/fYSsS
HdZ1qTqgozY6Xctx2y6vncyHuFIJsDPbte+3cWRP0hhPBrI86ywkFs48wh18Np7n0HyqeEPk4K1a
6DC9I5U8yo6MmCo6CBRmjdj0bRZ6D7/R/vHLSORJfKQf+A1ae51a8t03yLbHLnywvMcBuuq1fJso
lAOQXSaJoZmk242zBoxu6yWva09UmIrkmk0V+LQm7HxZhsCDKIdoTPsKL9iw+wryC+w64IrGg0WI
AFR1RjJPSopJxEo/LMQQzaXyAKGLWWm+aklwuWg8SBWVF6zF2HPq6HqqGFdPdD8m5yojUoOMy8wn
jcAIZC08oBIb2ZTWSLeyiG89r9ZuinGnCxbQUDz2Jaf6f3Zk+Ce25r560nQ04Scz2MKJMBRcofy6
bZ8UIMkQ9XazYcK/3hMq7mG0239Usy3A6cV5B2+BnXtMAWxwCxC40xTkKTkmZ7NwU9eucsEV/uhh
4hNsnU+DX3WgKPmaEpJBgHY0ZdhsN0F7Qn652Fps365x/PCoo8eAU2e2xBCJYT1BoirCBx5myxXY
zUZeg+Y7Gd5UchpJ8RGcN5yt9YNxmpYonYTc0G09d3U0XpNVgZQZqVZaTuQLjIbQP3TpJwtjkQFi
hfW3t/1XZwpmffEw+2+yY9brA1mnVBAGR+JPAZU6MIMQ5padDNDPWW7r043GIZ1Hfglcy1i+35hj
+Li5lsMan0tFYHmlfAoDD6R3gFwsGOUwZrvKuxMnlNxhHTm+ywQivfIYDQAcsrKl5kiNSyJROsf8
6CU1/EuO81w1CMuEssaeWymHjvbm/i5G2VohJo9Vip7fAIbuYGOB7RHM4ddy7fI9TF/wMe8hX6o4
FkNekZo36BceVMGhFSX9hTsaHeI8MyHRJuyBeoPyDKI8flAtxGFKzYu7/FqVNDMq4D+Y2DQkc0U5
jNpcvTJrmLKtRRhQNo9TvE4kYSstO8HraYRzzhm5OnKaj0Kp8b69Zm9LEynH3BxxhWUyVvA4209b
ireQ39EDgHTWiV2vTwdYkN+Kn3kV1FqutvwqxZPfKbPR8h0GkGhkCWyeJaGfC0Y0F5Wko2UEX/q5
1tphkRSjZQVXGhRqUpnPWy6gnWDY+VlicVNjJYyt9c4ben9ZDccQw9A8hwL+M53aurSjl/hShtOt
j1dmuMGIh/0qLqmWGTf5zSiTKysClyTJsEgt/c/CU9oHjefG3uAyJv3ZlM++LnFZUBgG+1c2Lyaa
SC1lpQu+UCZc8bUcXFmetkfQeTqqTM3OEAiHqnC8ivT6PPZp9gcrZBxocw9gMnOGRiNI/ttBDzRa
xhGBT/YnOPuEkWLw1r20tqL4AJP8HfqdkzMW4wWduY8+AFMoI2eEtWcRKzjeFfoCEYytoaNBy0Dg
KbcEZMCa900DMbq/6UMIg4nNoGoSdVu8QBqdWv6LF51dFDb+7E/icZzCDgmiGeZp5frGXlV98e9p
Lg+lZYcL1EfnSai6sUiCJuyJyUcOp0BHP+DTMwlgYQa6O3JttVKfpS7lEz28nTHhj8/aCDqhj+RT
ezy9x45ZNsfJI7kz7iicOTPqZQ1XsekPYzcoo04PJaK1CXjp8KszlCZD5blnbz5WnNfDi2sxqi56
KDJw/9AAh0n1EfPf+Lg+QICcmn/95wiUuNEfZngxhb4jkDE2No9TUtcA0Er5fMfzzOblEPsiD/fa
mS/Ug7fXKyp6QxCDHdGDbtnz2glZLXHjNFDggqHPJVwjtUvATnxxakJrWN6kid8Y4iA0q2vmefEL
WSv7xSruiW2KGD0fQhMPFYlHed34I+YaBKl9F/0zsbYbDRAo7vyfA3dKtMxHIPHoFIeWSxUw05qr
J/oE8QJO4lVeY/xlx6eS4PdlykCEUZk1b0FHu4Scoov8zVwnEKIShfzCW78xZsnCO4+/7Kxb9WcC
gK4B3iZio/e+d7pDVvek1TUSRPoHVXz5lMInIuA6Ro/2lpcNmjYz0kvjBL2mKjcfzumOKQm9sVMH
OXIrqZU3nKq4VJq2XubBO9XsR08C93k6IhEIVP0+CfxqlxtPpK2gHoJUgfGXFsDqNLOd9gVVHbtu
b19XQXFaUIev9PmNvFxsbMHIr2Cl3C/jozA17vbttuJDuRijYwVuYTgJ7fqPuurAovS78VnWYKsO
tnfLxLuNcN3qQHEr7GHCmpO+KYgp6+gZOcsCVcqYJ4cIq+5EmrY9W/zSg5RSe+v1Xk9+htYW/SwF
BY8QkcWSY52Fzw0ebCsS9p0QuR43U3NTuC12V3h4paWF6rkjFweksdYHY+pnMRaqCrO0xno4X8IN
bvs7wQ513jX7bHmofuVSvQRdiBzzhp0c1ylWfdRCqhcib8ainKMfyyZObtS9AN5cVFKqxiIuvAJ7
iMKXg0Ee+99qaSonJwcuBoVJjRbSdE00BMi2HU4zuUPyW+LU4I0wxcEJoBqhOeDNT+hItUDWTVRE
gk21Sr9eJ062Nl04XFupph4uO2Not7untz3gbcWMqLPVW9dOVeEYjEK+iDhNDo9zptB2XnADYvvi
K+mn7ioI5H4MLzpRVkzBlvQPLdRXKHeyqCigTuQhRIsCsEhVcREF7P4XkT3IQ+z9WZgn5m2dYBrk
3zOPoBP4TtgStZnHFp5Te3KuNRwO20JOsn5Bx8SnVSnoIqbdrzo3pJ9Qk5A8MFPfmVHVZPxrttQC
i7jExMbPVgk18RBP9hgwU5pHGGwrZnhUL35tOYEG1W9kkAnSeLYiGT1SuiEEHZen9K8Y5NNvLPOj
7f2tvQEjF56zJQ8g7CSvbb6aaKll10xzlHYkZNuvNf1cxL9BFTRHw0sIWA3PxrFnZZunWtwfAA+A
VjjIkW5fc/ZuTlm3CgMpPpN/F9wXT009kzLMYCjCgRQLygeDLISEZk2rHEKhtJoJ2cpQFiq/tyaI
h2+Enr/GU4kfvjDWAnOJqdXPJ2OtpDJt1pNat4tif2qBzwIX8GTZc6RiCAIrj5WDzpvLNSsLa/2o
ou67oLHV2JWQA4KvI1Mvd1rfxbRVGOsfbAyq7W1sF2aTJvaJ/rxOGBdAB4CQN1Iqi/vgX+HUm53+
Iqg8efWCS5cOY4mLbvr1yzZMMi9rw35+gERAbQU4XRoq267mRq4VsNt3YjkoZ4hrq/JcCJx11O0p
Fv0CIEDWMggXWfqCvBoFSFUTfcWOHouZZk2QvFzhtju2VRqENKJNMWR2CB/ECNXpxk3ZNtd0WKZL
8rFDrW5l6ZuBrdD+NWwxil2o+9+expYabGiToNDYUHH/BAowFFxBXPlpFOPMiouBifBnLGMmcdM3
TWEoQABkacqn6oHpXramhHYAGWhPeKvb9IJLRGK3AXZeh1xyd3hKdIa/F8IdCbaBfS8nBNA1avYl
vo5Eg6elfR3Yrk5k7oUKoOOpR+STO/tFucqOm9G85TEHFammXuLM7FFNm6DWhzpIVnXpvSPVLeWR
dT2a6psvtLbE6vj2hWtMC1tWoKkdrNxC9MkbkdrV7HqI/rQsWkmiPlCUzjscsavr/69S3DNvCvZh
4QmeADLK6vrjVWz2rMN9IbaRDfCTqBdIlzURxHd49sjT2VpVCL6heBc/lCaaxtZ7CV0iWrKqC/hL
EYUkdSwtdOt7dlobDGCXBOIRni3Dfl8wPqzht3ADZmM2G4htTs352Jtr6cIprp8Ghvu05xvwbBNh
PkESTvffI1CykFNjgzuEEm/ieG2lW8IhIkV91MroLSsWDoz8i768atxqYw+nCePMaLRsPyJD2Q3S
df9DRiFdxoW9luAJhLTCpgPqv0ZQl4YST/RsIOmw2jwNSvqcQr26ve22pWwCz40/0YvL2f2CqNne
3ezTy4/KYx0wy1pu0nQf7bkcBmmxVjEXLsIefyywLgRnVf744HJoSKqEBree1IVZjeRAMGXOZVlZ
n6EMjUKD6Cxh+pQ5drsMxXS6Xs0M6pO5cQjOX/bXO06p51cgMZpJWS9snkFKKy9ddwx6zQP1QO8u
ivyi91lwTkUZ6Ngt1b7BpLiOrpyPtALlYd84YqomyLEwp7kIlVeFuTvul04isyEvnFrbmlEzLVoi
MbqydoNDiv8UBqaWjKbzae4J3dTrVnm66iq5g7ojWkJ3krYObCDjAR2HqatT0fZc7xuWVeQc/Aos
qDpyiW6G9fZDDElVGxWzcla4JnJSP9D90lf86gSjJ6lQK7s1TcjKoaEWNd7NBapUmIIjwUqwo6TL
o/pAhlc5Cio7h5rT16Jlui4saLUaOKUHhEvwdUw+qfQYmrzHmk8pUsu+mLWXQyiqWSjnXhKP3Gxb
IG4/h7GCNqqlAbCr+60ynapgNu7PISK9OvmqvpXle5euBmjJ9DodcSc1gB3UZJ6HrqyzFyvzHTGq
riEHEHsF3uLNNYnT4kRwUv2Mq5fE0SQOWD0kgXiRju0i4W3KVIe7xveiOCN0nnh3TEf8r5/Klf3L
1XQHe+GiSORMr6EwfIL+X6+rzbGjTdWEnRGqKHpNrLIMbTwN4lgSgqo0cQQq2kB9aWT2BYME5bDc
XeGDjwPASjg5XdrtRX6t+6ttmgFPzcjbkhLhdo3TCJUV3farFtrCcV8joG1bCYWEbRntWNrJfEkJ
MZ8MILzQT9cebCxK6lQWzBQEkF3a3UBKWLQxx7TYrzN/7vSB1gxyjb0LJw0WlEjalfZho1jOSYes
7Z2Crwa+3aelJbiWVUcfi8cyUfK1HbF0LrvoF+5Vq8hB1nNEqXrU6GXKflSDVyaWPm+5UksnnKNe
+5zTNyDQkIeohuE5BaXotcZa+knDI3VpHN6Jdv7t1izQXx9yyDN6Uqtmaftvl0lmDsTBBOFOEaMq
z+wjjRJN617MIE6I/rGMv1BgZeJvtjVuGSCXg2bNrs4P9bnIcC0uf/n+12Jga5LryMJMVS3yvX/u
1/1mc5XbPaoyTEvtDrdrH28Ibrrh/uMi1NKWbRAFCNLWT6oseqh0zsUs/IYOreK/qz72K0s7ugwd
TiSud7dsEiuej0JNNLeDgzRMuUr+MWZC8Wf/iz3kytemXzlBAeSa7tN5dyvVZhPJZ8yDCvmNFIYp
Loa11p5GlkKDT5TaeL3SRMEg0I9/HyQgMblOnOXnZ+5ecWHcc1Kf+F8U8GQiZaG6O3yibt0FiDLG
tpBeVhcaeanbPCQ7gwWunPc1mYOQbpNCZBkJ+YTSbD/gJx+qUR/mlj6iI4BpzF9MD+XlI1hdlT9t
eflHGhtkAzsIzs2nyWqoEgxqqyCGFYvLoezyZhe7ftov2pWvB2SkJ3rEJFKrMKDzzhp3ZgLAt94K
mtVxGB9OF9LiRMFDaWn3e5ibEK7SlV5LK+bFvhn1nR4qUOFtwPygsg4CHvAee7ahftO1cDnQlLpC
wq2NoI4dJeSHzSA50Mkt8EWGTm35B18E7MXg1DWbva7dwtze4cDDqhqF8vGuyUD5N/tGHe15jh/z
sxSjP3jfKhn6RmJ0LTz6M1+WRJb7SFqcgAuOz6J9cVTWtEyKNaGnJ3p7/G4316s48nZI/7CGa5Le
xIUNTx7QDVSMt4somR1Wf/l7HebHz9jfACNZ2ejBPGVlgL3VETwBrga8imiO5XFUyMvGUJrgh3Tr
1cncXcE6Y+vMXJjtjJi4ug0FeeGkWwpW8xIMHy2wAtbck7FbXjoyeLubKF8KPlJSbOk2DbNmC1u1
/9jvYTz3DzomuCvk+k+7ElqFrzyGR9wMNetbHB44S66iN9HT/THDDGd5jSMVcNDjOJrhFBX0yKeS
sTBw1cdRn9izyRHs2sKXPECsu0Sk/O8EtyBYLKVnaw6+TfzA3oco2wbGK3lrBo913LwFl3yCxAt+
3PHsD4zuDvBk1bEQ+uqx5L68QMdbyF1j6VrdYVJuMsD/Mh28Gst6sRoPFyGmFKgp6ohum1EmXIeM
smc69UDOQPPjzaFUMwmQ/o57iiBDPEOmmkG7+NAQKUqbPmbFiWuM62FLCyhtMLd/vkfP61plYmtg
lHHROcFqVcG33rlNVyz9yGpII+r5nqdL/Y2JEspjLEpoe8Wh8r2leQRIOztld3779NX1M4yS8CVa
GxF1jmeWz2HwesMZT6bR5HTklbHCnGa066oyUGNeOjAA9BGPZj9vyCBMhrFtrQa/j68q4DZmV+7Y
vbKpnWzxXV8HTs1CqnX5ryylL/aiBoX78R2PdgqktgolhdmxerWBh8Tkd0E3cBC/ZGTjPJlROFaw
e9f2XLwhRsHmo8Wi61lLF3/5abWqsS/ZU3x/nb0aUmJ6uNTCpFhwic8uixQzdT4xqldBU76LWt2w
fq6lKwb1+lS+fdtUFqpkbJ0GV36uAXOQ+5jCnD24/iQ7sFZ3sH5J3m+uZXyT76nrqaXx/Uma4nL2
cxUIxUEH9isE97Co3g2R4TVXKZngqun/pj4X74QnMa5LAtTvH5GYqsWeiQc5LNlWrtPSgJ4RPopw
Nst1RsM66AAgbiz9+mhkQKynq+8gVvmHzLRd/F3NZktntnnCLD4j0F6MD1Ta9qXadE6RJPQMFBh9
As9CQ5vqt84o/SNtzC0l5qwVPEs8+7iZUnSlYCBSrDBKSu0USuTMBCcF2tD+1meQOx6kNMIekDrS
eOXZApm8KHTzFHGGJUWlK23KCnoCB+HEh5cK/AKFOZ8WAjSRd9qtgOfnXku1iutZQLxZPf+ivL0G
68xfhLV5BhLYmA64zT5skc+xO4EX7Acb5MKcnU7jvtIDaS3vGhjpq9zqyQTSq4sepWy0Hd4cBkLS
/HnqWtXWuM37kQAYWce1VvCyS9j4EcZ8kSsxZrv188PSGGbTyA2HD6zWcQsybtjK2ncgX78TDvhP
5j7F4OhqG+QphQnxbDcqNpS6p5Zb/tWSoa8VdQ0WczwbZY4R9hov1euyC/+lDPHs2NMlTzK2fLEC
12o+BUd1mbQiHqgRXAebUpHhHKC8pBnEVLcZmiYmvIOyrMFHULEB8FqiDrV1cD7T/PUyfwkbA9KE
W0mz8kEavNv7CkVc0EOaZmvnJWqXFpM5qxGFOdPagZYVtq8FA1n1cqdJfbNm2Kl6PY3gKaKYFmel
bmaJfNfSA6UCWi/9psNJHbZvWG2cYSLaSCMWxSnqcNemLQ2lpTSDoHK6HLVvlLPkcacl6/LTaGfa
XArnU4nS6aoSLzt8JfmVwAXItz+op64B9b6Ovee5za8zRsGQSjFfud2XDEfXja4VCjmUEQycxa1U
zYxURPsARhAWP7JwRsOZzvisE2bkFMs9M1sZk7yQVuICPRQiCUGjYZOg4uluUx/RINAQULOSBXQA
ditpZZpj+rOHVSkbyTMi1/fnlOgqjF1+ifkMad72uCCn9AOJ2BNb1xC9OyggbAwjYQenoQ3psWQL
lgH4ZjEtet6b5S7GL06V6iwLjWST9F9/3vPNuCFwM/FV+uiBXoE/Lus7jDUTvIsiQHPjLYB34gFY
gUI4+tsEE/U2i8XjU+4tE/1aUhvfLAYI1tLRZVIatOqX2SPaidENaiWifY+BLo2Ctnl2uUiYEu6P
e5gayWCdWAF06v/7yISwoLXrKspPgDuLb3wmWbiND7JTcxZBBcvDPoVjcB/9rYlG+KEM9x0fpRhM
60zhTY/53cUxzVFBeDRRvfDt14ZTW27U/lP2KYM2GGCjelrbQrZilsnfHCNv6Be3V9RGrfWkpyPe
KUf4OpL+ouJpjBARujGOCeKvS8rU8dR0+yRx+4N1U5pgGL26ugFB4D+5ZGoM2jm/KBc+QzIZdZq6
N0PJOsK6QAtT6AfEt35DZj7rK6ATeGC0Sg4x2zrPlNZsm77m1I6hW95eHve5W0IYqbDiXbOviE1H
5qj9cWW1vhqUyU9EHfCEFe3H1bKkYuEkWQ/AycLw2nWhBiRRhB7kvei8nSJE+mP4VgReSrC56lgA
+liH8AkLzR0BRB7CYGFl50K8YT8ZTg93PsL1Rkm7Jm8TxxMLUI/RgmvNmgJNt4fXAzm1Tg+gpXtb
ltFvpWffnkO60p8tJkfnKNN6gCrTyJYOp4CB1WSBmz6rXsVbCnPPJdHBmWQdbiaWM5g+UbpQUhAT
9WGfulOkED1hCpFD/g3GgBppLOY2DEIJZsXoDdXPfGcy3O3zO7gfW6xg+Uf4iXSBciEMrAOVjdh6
Ahd7JQjnvGEmNKChDPKRDAGIX3GujfNqpZ3bd5C4ZZiwj3lSWtcp6k8sRrXZfphUMhVr0z6ChGDi
7WyMcUY+jQl6AmxkYdCdbHjyU0k4Uq4rffKJ+KakanE4j0fZNvd8721cbJz/AAIxICVJbRztmSr+
C1qC7VMOdIJjliVKcig+IN4I03mLAU59zG9ApCTm9msdyi/JuqWGsHGt2wIRxMeKZ6LZpAg7Idqm
ZrFFgMijKHBJNLz/48R3Mi7vAWa2KXV/U5mVDrAu/Y5EWwUu/KvKlXM+EgfHaeBH3A0XsCmIIoY9
IS/k89QMagGOLNKAQTHv42WlQMKn3P8UTmen6PdEok4/eG6OhDi7RnJulH43ywUWSL5svkEvyLRF
SvlyYjmNbtljM3/uFeU3/0K4c3hjNr6Tv6S7Cu2pnSz9jnyn1pr8tHJOZpKeJsdvtwlpxxQ7lHB+
hzlTs8TO3glJtghXl1P8tV5ir06zQE25qmNbGQS0WS5cMGA4wpbzvi0lq4PRlz3rNKoHFhXygT/c
X4M/0B7+kAd39rUTYaKAzHIsQo0M47KCL6G8An/feVWFG8I51b5lhI6mu/ZdTDxobGEsQjUqj8VZ
b9JQgGrPiFnk/CruHNarBTE0IFg5DOAoIsk5vZavmkT0IMupwoefEPvH1jDzGcKhZ3tjUgUsCLox
R3t3U7xDQTCMqAtYKkWplYXNU4rPnjcaT+ROr3H/nDAne1cv9JY1bzDNrDTFrZvsFTLBeuG7viTB
Xycl52u0RLDfnR6ECbmDzKc9T0CYd4SYBZMvMBMZXt1Hw0oCNEYiLxj9UUAu3WHsdeaLUyxMG9qO
pIMP0c5x39UoTMY3eRlJwT0lDcTwKdmjGjCVg/djcIogRsHXRn4WT+t0jCSmMbEzU6kjntx5PpR1
CLTohsP3vJWieo5hAr1J4HIE+M7/I+2c7okuxd1/E5OldodTB3FgSmf3fE8aoqGnOEtqgsRVyPyH
LlIcPNA2IPzOPvVD7TKgHQBzEfqbDczWO6dDhWxt1lVv5s17ZHo30J4+OhEsJiVtTqXgJVo8dzqV
gTIpnZcchZO76GIUvRfuKvI8MRi0q0gCdQf3i06UBoUeZIXRP/QFMMLNH14mxtNW4qmLryk51Hyi
iRkNB4rH/BC3vEgh/1keThEda66rS6UID8QenqG4+yq2KUMvNYRS/dZnW/UjnVzQm3wnilRgVLH5
lfpji4A/zS6/4TCavFN6QM0sQA0+cKK0yqdqxXImM3Lj4uFxdLo5QQW/qtCHI8ByYbfKi4IF5Odc
tuNV63/d5+utP8EgmYTg7AV5ILRUCGCHuYrNLxmUzYPdN+lr0pg30T31QyLxvIhRme1ikplxa5PJ
Hq4Ibw7YNmQZC18gOt1LablIuFlAAg4IBbYj50LcQmj2mMg7IxgrTexokROSXMUjM/0sMd0OoGcm
LisYqYSYzoRLHqoLVeVp+HPvmufR4PXoBkXyC9MKf32MRQCe0/bZuhiNuG6FAuKXcT0ib9Z8jOSo
gwV9OqXpAXW+Pk6PKQ/fXcPS+g6IJ1xoJfpbI5eqXbQoxSjr1l3oHVMOfgnzuEJyzbZ++PYrcAzR
EcU+/5F2FTqgMGSNmipi0Gu4hraF0C98QW6q4QI8cv54+SuJSdjM2wMXRParuIzmAoByBO22qYus
vOpPPYbiK+1FEaZL8JTGDBoYD3h1+NYVhqmdhPiSj12Br1TGvmnak1HGiIKcNFuTYIBST4m8mGcr
bVhnolmQIwgVNV5WuDirMqKbp0TTrZvM+HSuCa5wKCiSQIZuxmrxzcQWsF08WSELOZUGGs6mxmTx
vsbqZA/XMYl8stHW75LP8cPwaY+2LBFiNNFrFXmNozrzayrxkiYUvMNpxtl+g48SHbJ8OAF4JY/F
lpK/bqCQo5Aiu5yRtVdqCPU+9qcsQF92t1r3OVwHe9M9oo403QR9uo2YEJtCBMKrRY1ue8yZn/b3
evPlAJRjg/ESHCe8IhZnUeQlsNXqWzdqIuv6LzOWLIGJLq8YHvWIFMNmFQ8plSadkKdJ0AYx+u9u
43sNU8e7vtGlMylMLluwiqWi+KgDNb20jhUbUIFryo8X3kpsmu2wwv0NX77Y8Hcsrx6WwKWUXANs
nUaxFpSKXQs0b6M6TGd44cTzA4AQs6omZlMxxyMm2iesin7iCbrVDQcEuIOOkNrXMzOAfAaYwPFL
XA++QA+BFg4Fb3hs73eFFY+cnQdZqFxK4sJa4EkLNPEn61nl9zucIE1/W0uiFs0IovvmXeUQaeRh
VTxev2vZgFq3bvBiOqvxGdPrV2jllJpDLa58CB7CviP9yFeLAsvXSHut3gDZof/rWXLfK2K4fGXZ
rTQzQhcWfMUEHXRAJRqe0AbyN1FYXRTGKc6+xeb3MMosU32g8LXh+ZxBv/J5hBQVM5ne2ofu3bbM
eXBwu+Q23keOJJFRfd+Exy+LEMJGLvQW4VIIcojz/uPlmx7vLD8VIAPwVx9Eg/pAtY98L9WfXr3X
uF1uhCcTa0EU6/XCg8svNObWqwvcJbr1Nd6TimmSbmvOJrVtkjiQfONqhgH18D/uj80d/bb/ph4m
ik6TRFGJqFS7YkOWCSaqVTJEidPpPWb2G42UMOsI386xJ0uwb4oqKANpHsi2m6/5q7aH43B43xAo
OwCEdoOjymlMQURsAmmZXUqVjwSOMHNMkqsmuB29y7f3LcNlmaX5pIvAtNYwjTECvuxzVAGYRyC1
05BygZ2+opS+zxLMv04ZQz3LO7FEPI72VYDa1/mT/x8j1oBplWqju2taq6B14OnWIYlPZZHj3HAM
+VTT/2gTen/WmWbOUSGJzDOJl0c0qZuxBNnyuYeFEWAhgeVbOXsd82vIQMbd8Y24QGHOgTHFaq9g
62Awz220At9JlIWqozkSczXUgbon7DMRXNC7/tuDJ7IOiQ4wA1znMzuPRBYpLOWvKaMGPxl6t4jA
gplR2yJNVxX95arg/Wx17I6seCWVvYMw/GbAhHrtbsLG2dHLcFqfS4S87qsnDiQ9S1thPoIkLT4+
7jx2nb6CiJXbomc8soYnRzF3+T9FEhMfHBfwM48MbxLm5NVkibPdkoh5AHFHXdqzo7+MuLKyu4Ta
ITQqPENMx26x3bPCO6BDUhNxKvVthrNqYXazIQyUMB1rx/uuHCaP6a5qzVF0X9c/mZm2dBdSz8Do
pm74/luDLEBQkOl/j/fVhzrA/N8VjR2WKNHBZdDqD6rYfWM+cH2gu1oVstKJun5whpzy5dSF/caD
UGfwx5yDA/efrbuapHnqycxxWnW5gWq2pNOcH/CPLiYTzQfHQD+A02xCCkSCtolSaDwBDoq4E3xq
2kIgPZPADmJNN36uu7a+jNkJSuRCFcpy1uIoeGNXRqxPEEIo7ZaTovN3vmli/FGPOwQMHboMbldO
BJF+9PwhkKOPpWQFhaIqJ/DznOO/mQwew27QeYvHhL0JNFAb3iZuNCqv+lviwbVQoZHdcNmiiqSO
alJ6IsGf/5hFPgYIGhz9ZeFS2bXVY+dfV8kABeL0MZK+q7BshBT485jtiomoDoe9RMhXdGVydWw9
+95021rKU02XgBXbDyJYoqIfsNRi9Zh0q7K22Y0nKdmVUcL+uxT0z7nLUehxSgNfqMd2/fWcA49P
VyGBIDPzZFSMeP4M9sk0v9lgjE18gylRhAA85mpSworkIIgxQxyHw5wns9YR5xUmGOC+9bpcIbaL
9jEv5J1CEeMaZkvzVswE5bhDzpwbmvhXznQEmqhxBxVbhyYNxI8/7OUT5M3/6LxOK9jlC44KzVza
4GJfOj0CCaxwvtPjunF9Hh04B/JSTfbHLeoKUFbJba7mwRXJdVUe2CJaisfU+ZskgXRMhDzUAGZS
XU5xeyty+7U/kp8cIc1nk64F3daisc6T/f6UMlO9028ux0TEz3BeRWuVEjWnU4nJLSlAprsYpJvP
BQBZRfom6PVTRaU6d5mTc2kiqkqkdmrwh5DeJ4hlo/znQkwWMPXxJiWMzoC2ui2X6HuI8A3gylrs
NmM1+vgFHwO2PpptElIOyOD70W5mGQBdnMfF65CKkZDODnJEM4IDyMMPdClv2Em4EFKH/zO0ksyH
yvOlxML5B2YAY9Av7NdSS2C7Vtu45kIw40UuQtICga86CWjC5lW1rK3FzF8QweyixqdG/CAajJub
DvdaKCjwTFbAP7+oHUajAgOIy8p2ZXqCg2iqqljz6qNihdcgkczq+LFQJjbvt3wwZj5Cb9eQcoFz
D3TfVkOBawydi1jrLKaecuzZLf5/GLTZE3/1qfbu/++XT7lH+VqNKqcgqVRlcaUjmICAIxTl6MDv
gayHm43h7p0dZJmyT/+hiNTbGXrGC6xS/TuTn3yiMUBg1LZksPOW7hjff7rmOtq/116NSfWCBl+r
IlcbSodusKaePi7GQ0HQC6hOUfbMnQHOBiG+Wktv8uAkuynCCSaUVCKokra9+D/iI2KyO8OhikBI
x7QIPlGVBQqx0+Cow4K78H+OyN1TaSO5wgBPvXT7r3KjMyloxuzz7pV0ga3RsEQ5Qo+aKYgtyxSL
tsYa4KMrmGP6aFLWm+WlQN+5t2xij95XSc9AbqgCpvXHTMOHaIpqMxiRhI0O40Gq7ot80n5c2hmt
2Pxmv899fI68u2Wm0CPbL4BdZYfe090NAfAxgdUB18xKZsQaxZV+KVSo8/nKMh1yyB9vlNrjGA+C
jM4p02bBUHTJI9nRvqo8SgXSUm8m99dSCMbP/+uqjLW31Uyv59yeVaZ/QFOU7WGTazFU3ggCh1tV
dw22GBXgdDwgCTQ9M9vYGq7tdP9z7uMv206kzzLeopIkEm+VokJRNpzHmEuiManFovp6zGiFLZNv
2tUhUn9WRbdqZiY66AD7BndS1IO+p6KX7AzB7I/yd4KeyXVMxJXMjvNpdPH6W84cl6ZiBzlbUubw
M3cegusD8EUUQDhbo9DvMSDATWIW9nsvqYFkoODjWJe/s+4P5eieik3PTPdbYKwToiMAjGZZMZ30
0RrnD545KXQG1BaJtNx1gBY6EH+/z+EzzcuPIWEIHL5L8feQjonT14MGHLbEy6sNPCatyLFRhP6S
klm7K+bvbS7olWlWXIdiGiCuWr7KwdP0kkLAs2HghxzZoYUuIo5CmBLTccOunurcOULnIO5UkhU5
FK8w5aylvbMAe7iCZZ0l0+wCcf9LcN1fa/NAiKtpgY8jMuppfA1p8cY0uc0X83FCxjJgwvyDzSXJ
z8LmjfGXhKgvnoSd3eS06Iogn349QI0qmVEfSIenEpx/7tt1HwiBz9YdmxLyUyMe1gbOi+46w061
r7265OfrT7z2oXR/fNpGsx6wWFBJI5Uj8yvL9VbnxyL+RWY0i1WnyfEdmh1TTiMKFvPcnwxPsRXy
WOry/vksUl9kfzj8nD4VyDRMORITozoL3/vUBBeCLugp0UmYpEumKrvummmFX7Yh31Sv7Ux7hhhz
TyVmN91zyfcBWYyZnjwEwCX9pSqLSCSh/cJ/p/vD6NQOSjr/8JpHohzCea0xofk15x67fEudSIu7
/pr5JMoqysnndHcbJmE9IM1AHowJkzrF+z6JzRqz0QS954G6rC4Xl0bClk2VMA0JhNookILL2/XF
bcLj+L8xG04aRgaPNOQsK4nq2ZUhaH187airmOSovrgCDEada9E81WPeh0YW4OQca2m5zwguld3r
ixnLmE82vPK0+ycxZfVYzWnRNBPqlVAgfLJZ88mYyRKNB4/SmLXR3pKmKfJPRyImZuAm98KyI2+l
cgkwhgIzy7xPjUTEh7T7BNUGwM5Qk/7K6sq7wtsyHkVv5cY2ZQju7FmYg4m7SI+GWBiotrZL9Fr0
XNhfZgUY1cXZGWx+J+IAWBq+e4rYHBs8kP066I45ruUbgS9qe/z0r3UpOVykKaclf2MWMPrP0SrD
lpmC5U4q5QMVJbSu0uyv8BFEfHSXfkcUdpsQyRbUa/JQO6aubDJx/gkkcFzc2Bez9kB+CJL7JiX/
LbyRT67L4WUhoXbn70Oskr8wEpNUmPT9Z7H7SnlCTlIPcO1u9Cz8GytIqJAMk3Y9oQVhswGCt4I+
oohbEGGvz+2UCRDI62R6U018ONdE2c9Qenwss9wsbl39T5IZQcIJNcaMS811oXAsd8b5aCn4Befq
zczv9/srLGIhHJfrpOGsrsLHJg2uIczDf3768KF8vn/owrUxmHkueWDjtMwLgDC3lSlMP8JWhXxR
0u923fezARWzm24RC32qmuAezZ/Mp3lPS/fCDcSZvoHCHeGWsYDQ7pzYEdjSTmee6SIN8nh365tD
QF193pBNmI51j2FtKEBIMz5RmkK6qVMPT6Q9bTvvWJ2hUur8v11325OojaX7tYwQaiqOUvVBlkrM
Yh0SWnw9rBvMkC9oRWRSa6SVDUDizCA/khoF5dLyEP+lu35Lraoo3lVBbqjKMaRJG5GHg7nJvTWC
MRsf3EAwuGdMUNjfjPs3pYPhRc12fNZQRwdZQZUlUSPCQom649TtYCCzk+ZUJLygCKomTzbhYzSg
9KAMaAdo77qEem7osnX0/8ysrSpY8W1PsLbgQr4LgVZ72zfKNVfyg46Up9yYvCUIWg3TAtX1Kbo3
+MQ6WPm0nsVK1TsrnEYylQ5mHnESbeL1e3YewfITAvvYUqsHra1PiwYMjr6WUmUECodviDNw4yYJ
hk6Eq9cwmfe+GOSaie4qv7Vx4Jj2SZ/NR3IYSUYVA2i1wrW0z8zRzRj06SKJm/qUl4LUqrLRIg5j
8dEj/wSxZ5ChniNweHwiOTwhTcGUjgx5p8NtMdC2gZDa0VNt3DM8wSKbI/SZKlWLO4q/y0PZCc8M
YjcmtzN4AEKKe90qrFt3XjWw5TS7rwgWIe8otJcF/YIuKYtwPvfiPg/SCcAnd6q/u1pk1Az3/8dD
d9GT+yJZk/rryqZgN1CPFdvElB9KNaGDBFmxmVTVn0F7WAPLOdjxUv2XsbS/SBnKhfeJOd7f1zjA
Y8sZkiWIEDkhe6pmqV6zth5Di2WtWe+ziPygjTpJHPvm31YE0Ko8/VRYoOJb6iK1p0d9wlBveTH2
I9mcXL/rPlhP4O2FPSqBSUUQlG3U9DnK/h/zl1k/03njY7ULEEr0Wir3BFp1NmUd1TdUvhrFUR7T
ahQEMi1pgBDnJYV0Z51I7lB8c7wmCyAGoFac9cnsgUtLhc2u9sflWF/OOCwfiJhc+kgARoh8/+/r
xTzrP8N4v2DXiRvWgGCkjqwUhVI3PjWswVFH2W3aictzE3VheiOwKGWKlABvn3E7hiZYqQZSGT2H
/VfssARK4nNhPF/I0tLScCQ+zQhYytcX3oOP2Nz8M/xrJPIVm03solBikNIJoplm/dYkNTMxNI+Y
GsXdmX6tcDe44wmGcmIV3Qg5xZvqhMxeuWn3lhSxK8l/p8B12UyfjsveTLoJ/dNJJl+FzujMeDrr
RFNpvPIKUOTRPStVwkN1ExVC2PhEPmUe3L/JxYPmJpft+c2cJEWVARasTj2Od3lIFFTIkUegFpJi
n4qSYDVpuOxoxoHiU7Qa61ceRbE7RarSl36iqaV5d98jGdOmNoB/WfIBLX34PvNcJEQdC8SX9CVN
NltwwiB8qcfJgOB51sFUzOkqSlvKvCvMbajn9DxqmVWLCmoyBz2Z/vMlcj8LOqGmdZfsCrusu/mz
13CYiVQEW168m9v2JE7SgnAsNH20R6b17bbSYMvJ2DmtXjebhM8J/kceJsi6Or3aa6Ur6nQwFbig
fu2wKUkn3MuhCry1zJNBpxV2/Bv9g7l0ue5GEpg+gatXhm23tGxWm18yDUvx4ye2RwoqoWlnLckk
tjD3kTu+Mdm4sCVSz4LLnDERbhrGzEY62r2Jqlkzpg3hG6h+H04+CccJ4oKDgp1YORbNTYwHNIAr
p1dxz+fIvYy06jr+byFgi2YyWBsafglCXdSxUgtW7w7KeB+WozQScud+M7sbdi5FulsmQrW7apwu
UASXfF1YebPPxG5bXSUrE7YhnYpSZrZk3+uYzViLSc+xvtd7pRVIqgCjuaWD6eCUyink7350v2Ju
nP/F921m7s0WJgc2vmjSjeepSHZDg5FVcEWpQgLDBMrQk77zVjrC73ONkuTs2mq8/Ir8Sqo5s5DQ
9hXYEXdem3QDlRJ9wvHoaanHxdZ7A56HShL+Qdw003xxIhmFTAhomt4+gesrWlM9WDq3jZlcFUbE
CFt7S4Pbk3azfkeqRP2bz5Sxno5s9S31HIX1YU155tOHxBcPBnFpKEAbR3XQWy2xQzRQ8tarY/x2
nG3TUbnDsYXFK6iXqP6UjFL7Z+j4sxZtHckseniZfxkP3gk0bf+tAHavEkIEYhPcDlxfMamPNY6s
unHqCoO4AvFl9LFPTIqZABllYTlbSOEmW7BihsmY7fUBcVqk99OY7FU73juCljt05ypPwheCeKxq
lUQyxBwHk3rd62STMYsaurbXpIkm7ZIc5ePwp3C7MBYFDJQKRyjud76WuqOiRabGD0LND1pex8mA
A3KKKap6SuPxep9velL2GZ1j67e0+ct2541YZkym1QKHfZg+HwoDH/S/fb/A3IDWw3g6dIKmgIK1
/drocs+RyiRsnOPahXkE6qa1Ymj2vhFequIWwTq08urBcnYFAcvdEGstFX9h9r1M8rBxfaGXulbg
XRMwgGUh8b+kDVCiFUVf0DRklL9H7PNJL96EeZOrkEstOuzid5XichZFI7V5c3r3oQhWJhlSdOPl
A2XTMx9UdV3Vj8zpk7qeBIdjR146kFEyv0/zPn5hSmkkH0BPTYcjei9u8X6bl+s2rtKEq+m3xN7k
0yredBcdQw9ycV0CYrcB6uctHRa4VMMT5ExF55nGws2SB+tLAkPHUv1NC6P2zqXqFrEJLLiGjTvF
fyBVEY+U2Mblt1NthuQR4bHP+OHD4SZ2Zats9pLhJCLg9xttZdaThwQqin0/y6GMMcHbX4/tHVum
8ilPXYhdRxKu4u3o5SRu1tuLmvTfRSnU/jjXINEQ1Pqjr9ee4ta/Gm6zJIsQ1DiL3krtpQWwWoEP
M1WM/ndm/H/ItD5+LROSGVlJwlkwqKtVPsbZRcEx+s36t1RKZditwBE3uBbgqmi0N4PJSWLxLTPf
jHaUdzo6aHJS/m/I2kiE1BMrL6mTJ0anDaC7xGyRw85AmduWmD8D9whtZTG3+9tggy2AZlDDGtIl
RXicgZlAb6bgTW0pJABXqp1UNmiJkP3TR6GlDJSQCaLn4ZkG4yEHkDtdfXscNaX7aUYBMStt7LR/
tV4ZZvMz/PSBWE4jKrugPt1iBrqYyFMSLHlbTOR1YguOUqbNEIjAMF7NIbXCVQt7ElIE24pJsGXe
oCcf7Ry5zNvq0MemgPC/nhMIRhQYt6y8ZDXSPNIjIM7k4asMXdPcE+2pgDg26n/rHxurdwec10WC
Us/gZyyFgekfmkNE3iLfUv1WGiGrHqu2mhz0NMxicG0z5VTy5ShqWN5sDfFdkwvAHwJGe6zTFJF7
25IzAQx3TsLisRKSYmiSGW4dDaDCqUuUYedEZcVEg/3hIeLl4KMqhuWbU5Yi9ckttbetYK2L9lol
PAkyRowzsCXaKXUfV+NCFA4k1YbWp+9uGrE13bG4pszGoM1LCfbELgi0zhmJErj6wVSHpcCKHUc0
0R7rNSTyi6dwrsSzBcGNyMsu8XCXKNwO9+EiSAh+SvX3A5bSJo+EDOGcaAkM/v2gAkxw5HsNtQ8f
rPJJSecPMkYXl9yPzG/s6a7LHZa0HLunjp/gr6Mq187Xu23teUB79RurVhmO50xdgZkDub8dOUJ8
P1oQu/zkY7aewVy1YaBtI3JIGPzYK6wGUCPHUPujL2BsoaLZyzwjM2U5PRtC0mkQzknS/ie4JmqT
0la4ELMq5kJvM5yjN0T9tG7pMq+5Jla0Hl+Bj8Y5rzIy0qvfqkk6JqgYC3qgfsXdgKOxW/8xsXSy
GRtv+8bs7BrB3WUBqShZV7O69MKAgv82gddRiqeGw8/1Eyq8SyhhquTco6p9lgF+n6v1KGLXUAxg
DsM2KvqkD254dfqLKNvTFxTwYboELlMfpQwiK58rLVnQqD0e8PddBBz1E8EnR1M7Xema+w7NMI3k
/OKNz5llPI4bvaKJN7o26DrG/IZBkyw2gy9g8AbcFIg58GNo/iOav/+d5xhHwwHYPboR4cd574dM
AfINIA4g/3+X+hkRS9sbJHaluSK2K0SoE0b9rKxZr1YfkB8VXGDbSCiZ5NWjX3ilJU5fHz+Befqy
ZqzJt31pif+BlyIPpDQjGH9YUzJlgEubeRSryeushQk+OkC5kAEkdYuLfPorCSoccZEURkIIgITE
9DYK0QQwgIwSJnR4HjlsZUituTiCDdQA+nxFE2Ezf03G0jMtHhJyKWlHqIccBpFW+wVsv28wKkId
1b/MjIOmkpcXzCd5ncolr2BcmXC57S77QKqWgW8N0/WRu4/VgcObyP809d10s794Iuv0qEhWuYW4
ucKppa9+7VRNlQWOvjTdQfQqGz0tb7eumg/KcvsAzyrKe5V3KNeIEWWGyHVg8Qh45bhO7IDuUb9B
ihvFL9y9gbhvnx9Bp/5OJVRkTmaCEnGulnDcqMglCJpec/E63nff2t91bBdJULf6KvNrGRxXQveQ
kUEwTpgyM15D0YJwzU5milCz1in0jHSG+CanqjwblIIt9szKdFqPSKD/AAHfw4lUHDTdjATgS7j0
lp5XDD17OIDjMAI9YJQ4kTFxqHmXAhqV/BARuOuaGuCXfkcZ9tKG8wrtrpAqPu68sYI27DfkubWu
qB6/RiugXcuv+QwRX8Un9eV+jz0o5/0uqUOrFXYeJnyzwl+uPEgFjY9+INdDxkoS6QZlPSd3vInY
mHA3VitPkWvrgzH70QOAncZlZMpzCGBoyWUY1n4LEqWmtsi3fymlN1rwY3R6+MpDnUc2oiZSbZ9U
XHLztULfPqSI6uYgwyYHiTWtk8RlH6q0qRkZRpITqcGo2vkAuwlzi5XXOT/Ob0pww/Pa4hUHoqRA
mCwTajdlvAQMisUWQy92oJBPJtg9md3PuoiixcvuBumRPaL7D9gmsvm5C8T2Rep8ndEb48hCW5lZ
dzBEIdnLwMkUlfvEkE7XR/N6QiFvnHFFhgBAI6NfYfCnnymPz4n3idqAHpeNueVRLL/BzHZ7e8W4
1MG2uhEpoYhSeYoHyxY/vf35DGOyMs8DQAiBQQreH/Eg2rJjh2UKgM5C/94MWQ8VdYN6S8RGitgo
p+F4rPdzk2hT/ENU4azQT8uXdr4VjWt/HKM2xxVqb+vLO7SK0pK9YstYmt8RX9IMgF05E2tgxJH5
HkeCwqJ3xDFeLdba9sq623SwXn/mJ6UOG7fnEhXoqlcsU9qpks8hX0r0YWavsoUjPZKOF+uU1DI1
5FfczRmbjBle0vq9ldnfg0WD4B52jPlqn1yUSkU9U3SXG6+1BClR2eSMV9UWHl+rR5M7nDCPayr5
gdWTSMdbWIrgt1yNgouNH4ebGEJLdcKkOTNZD45UpBZKc4lkbjShVxtyYIMiInhGX0lCVMh1xaRW
AafRK08LiJq55tOIiHnxnshrRLb+P2a26z5t/tni1rf1uHWjQa2QBnRsu/KbGISMBUbRcuchntHe
GiFfGaoYwRcGjHAHQCgIusUaxZsOtX5hTmh/Bx0KLJqBVp0wfeTAy4YJOc+E18xUwL+1x54x5FRC
VDis2AyfYHMSidqCcxgGH7OtX2EX6Gk9NZ/FcJzCQhN+L9Wo8K60/Knidz6j5lv0Yqp/sheU6LIW
ZY6mEhdwFwgsnIf1L+UahgCTXDgxUQyVYYFoMJJ64Po2DTfCyet4sc69zV+y9hQnZ5wpQefM1trZ
YlxflLkcr4c+J4L0O4BtZl87MvQaG2HQlrtMUed5tWS3oiE170pSQNFVZaxGIf7HSbgEXe+cDOPj
lqZ5XUvSQG2Q4x3UiIdAlld5lqzZH4/TOShz5WGFr75GyRLNMGVmGpBoo0SL2yaT6q5dBVG7I8Qw
ARVQYoJ+7n0QiH7QnUdwEthWunu34KykPk0PJ07RwsXh6ZdrVd+ftuOfGLR/aKZ6WSHmx5yo9uGm
4jM3Owqd6ziXHiN4t5fvs0t9JT36prEBnDQuFvAhdB5dF3FLq61bR4UzqB9Oy6Nqn8FhwtZ4wBqa
CcfRP6+dJpaYhIw6GUo8hFmSl2xNfouCB+R5k669ZdjWlJ0sBc6wu2PzYhSb5G3R0FVIaqlrMuqC
uqI9Ha1V2ITqUWfFOcGlrV/G4NuLmfEXepHQdG6CBEHeLM+gJ9lrde/i6md1YxAZZIKDKzIP/1mA
vZq2JvwhDPTMhpriVqz+Vr5Z3jZnhIMGWZk1XAXMd+K97xtvcyrUTu3ndVGWSnlZVybVx0k+1uk0
OMukn08/gb1B0ILIa0gS5RIKpoInctZ6d81xXrJPL89wENMLECWn8Fx6UoHstDPUUfOhXsPaqz81
tu4Gf8Xc4/tftGxED8uf5k0WR/4hwqhXrKwrgQc0+QMmwAlsWArnZhpiSaHa8/+XFxyEwIZ9zJqf
elI3/NAsDGtTmTW6OV2Qp3PJDR3n2yFyqu8YJPR9LZjXmqUhTnJt0sot7tkPq87f+v1F7z2bzzok
xYuD9UdP56MHhCbDE3lHl4FJh10qmvcAbh5U4yKR1GY0NZ+inwBstnKyC4322ZMWYODWSPff2aFc
39HHtJqNAARUvLdrjTBhzv+YdsZbSq6NNe6RUc2S2DKjFkIi1FlauMCNgUpWBbF1qAgoBgHc2r08
ETpGAttQ9n0N0VT3Yf2MMn3jkRaas0FCv7Z6W00jvOdq/eAoFlejIvGsW1ga1+U2eCgDYrNm8UVR
us5IkPVdcJXY+L2LSbDf3DAuC6qLuz8fapKcaoMgr9IcYuQw2nUOTWxED9hf9UZ25iuiJ8+uoTvJ
HvUP6uL9Qw6NdYGhUxbJlAUxR9xcicCtfMqWqq5M/b0B95t+4EsTqick297trDzBbyEKqIOdt4dI
QrvWqUcExr3q2DGmg3N4k0Em753DAtjgWVcMQQxSknjjEY4G5InyGspWddsxDT8tgIWxlVBtKPUG
l0XjlnHboAolauK66JQ+sMVoH+DXWPXA6mA3JSGKFccxV2TS4XQx77BIYP7eDxa7RPLmHUye0cDj
Cx0xheHILkTDDvuQUypT5IWKOCf6tE+uvGtRQ3PeyHXdJbS0X6r+vdHps2HlbkgPrF7kI0eu9iqk
9/oDDUIzwrUVJyQ6E50gJq6KdfE2DmFT2f6fe9QrRnIWy7IlsBNBzgcQ+dc784TYGWJdbNuLkVlD
6QOHUlbi9nvn0MFpJ/R94N3Mhw2A2sDf1qIINEyiswmNVi1Kl4Z5qU1FWrBCLFoY9eAeLKvYMxBY
d+qbaZsBJoK4OodSCa9j5Ji0wE6tkblk+pNNeugHgDpcWSSoW3rrC5gbzt0MdZvjsfBpcnvVs6rL
A1AaRpGvpDuZ2xgPrZJPp53zu/s8vYFA7AaudM2fA6smL6aeOa/sFt0Z9CR8tSbtrUnFv836ANoS
JXjNKi4etVvKcnZ1a7b0VSQee2o0Re4/y7ovTFhtEyoejcrVA9fon2peH7ZPpixYRmdbptNeWk1S
XZqyhpCmkLuaEonvROsfhyiPJspYc4DIf+84TdiUJKfC8c5kEp0uHbL9HkN1Vz1LtzP9ge+TKwdL
Cpm47Bx5NfDuuZAgqbNB/ficzWIu7HkG5PGVky4o7Bz5V6oBPJBxJT+yEnp2UOVr2sUrQDxTrOxg
cQRvLrJcboLrIP2l2hv0vfttCIkRYnsVCRbIgCBTuL3NCAON5NDffFPOesZxFWqFDu9e68LYul9k
QQWqKPnGjX3vWBEgbFpqh0/bcdOaUR+joDCvOXFNo4xUJw3Q85F/OVdDQHXAJuaoA4LOtnuZzCmf
b1UZgcmwCHn5Mk46xJqZJbnUTszkf2z0iuzz0zxI8d62+qGg7r0//UrPZW4ArRCGksv6QgYq3OfZ
tJcmDJodvJ/ViqlW9Zl3Bdz5JnIj8F7P8x8UqWV5+0XgDtw5Bu0xAvs/sAp5d6+8b9MEfOu9M0Ao
7UnKfhIYbVmrKp6EPkG/Z7f1+O7Rh05lO8QaVqASJs8mACXgiWPz57zPl/qo+7NQa/TN5ruvB6gu
MF0mYv96xH5+bgMwKFgHENB3SQF7x95F+CbTWo+xQmd7UmWKCk7sekL/FP0zuBg3y5fN70jMYzr6
yJUby3+mbYIvDoihBs774N+CCubP/9eCDOQcstpy5waD5E5YxR0NM3l29i8Vo0ajxI0ooBCRGO/c
cxMjIsY1dsUCGDKmg2EQ6+GRFu9WI+ySTyyr5/GYCLFbphEQqbyU+IULDtCz0BhE+C7oDO8jX2kw
Q/igdqK6pBFQqqENgEq8/MQ+tLfB8qv1v6z6STS6qceR99asoLDKOuNKZFv83nJ1wGYD/VTYG3FL
vzIZc7WalymiZDbOVoE2tqHYQ5XlWjNQASkhCFOtyCSMklAJo9ZjQODGrroNO3FaDCVaqYcxxsXl
lF05DQEyKDt8U+j6pTgL4qoW7sY7CI1RPhM8yHbTYTB9EYHNfs8eTNAyZxk0G7G6LX4VXAWm5fS/
VUvohdjpO1Aw9Ils96RIqGkLl7mNfIMYfX9y507OWkByjCsd6nNiI4JsSA5kY83JOXUcHIzuz73i
1zT/K28E6Cgv5+vMWOUdI3I2jlljq4Gby6h474WQEdwYlW1c1ocmYUJlK1B/svQC2b1gQ5tgpABA
kGUCx8iA748F3IfV54Xb51kojzG+tNILFbDZcOKz8dlV5tghdI/v0D1gzVIC3I0ZGj03KJCpeKyn
rSNS1/cIY8EZt/d9H8ZFen0huX7M4qHTRZfyFWJgejoMmZlN45jOGsMj73ftcerLhxzjz/a6uigJ
ap8kFcvzI077hxWj5sh1fXtZv9Ls1AT71bFO6ydGxn1e1b/cusBWgi7/G0nH9otjIw2U9JS0Bbtv
tUg/1egGXZQzNOaBocQZV/tWbyI8I+MsTUG14uS9mPy3jxByA3vMDv8Pder6ePDamwNxqFJkQ4fw
c5ZLeEXFXdKhDqbom33F00btoSjGK/Jv1pnri6B5ov5wKTTfObgZP3imDlEBxU0ZYzR2PP+kM/ue
fBimOH+Xj0fNy+CxyOH9jtyY+S31pTa2SKTANRFwxj4bskfjaBo19qRLb1FzXCsNwolRqUOYA42Q
gXDtTJ1Lskt14rLEbflYiBpmPgE1dpjdTN4DJy0Ke3ie8SBz0SIO8bX15/d0Po5Fo7VsyjhF+5cH
dxxGQHT8xdlhybSMab+765zEVHW+lUC5AEEsWWV7FjDJBupXRRtnwYtGwAwukrkqRHVrrsyqL7O4
Jn3L51J9H36tuxz/upq+MLF0NgYL64CvLgkUiwgdEa7pwORPCE1iNm+0sOkIPETSERr4i8UjwpN8
1ruFbEmu8x9Shqp80WByGC2svvZ+NYup95tucBfHHAEJMdJmPDcZCV7aZZgCBZx/9/TIVrbp17rO
9F0xz+z+blZySdWshg3xdVaolO9K19j1a/d1QnO0BHIQYc96nSQ4xM9VI3xPKKHfUMP/Bzcbgu/T
ua8Amq7KQmUAJMCuXwvJC9HayByUYeHZoULRo3uGtUyOen7HAxrdghJ/h7Gg+p7j6QdymG0g8hgz
xitVSIU6OTQv/S3Hs4Md9PtCHaq2LkQn3kGlOxuBMNeSL3Gh+stnDFZgApDS+CUhj0jZNyNcNBHr
GOOBXqbjXxjsB2ts+QCBqcvvjOXHGGDYG0tSqCwyA4aipZGvp+EIJmIi7MPA4fgKJLc0ZXAe2N6j
VVSP6KhWPknK77avPir6aELWNj/RoJCS4sVhR9cQpiLN+ELTpmLJm4n1Ta5Kiu6HvVpNJXban5bE
0C8a1BakqyULKl9keWa2xYBTEbH7MSSBL7BD0L8EhoZOIfJ/D37GgaCR8qkgFI7S8O+ptmmVioqZ
DgaYHhFIl5maM/sNd0RJsoznUI6/XWQ0InF9dUFaeFpAejYdlLWSrdFfw/rwBPVW35cDj9daQ6kU
5xtPOAYCtaI+LUJ0bFtwNCyQkR294MV1jxKcSaozSFgzV6zHAs601DqM1Hdhvt0bLUfBhcw5H/Oe
SsQpLZqVlTCTPHEau50ZFM4hwQyp2XFJ+lWxwNljaNB/zSpa887tDBrt1aVhCHUh9zxM97n6QhCG
GsmBhQRydX+P6NzFt0NtcsDpeXlUIgeh3t6fBHB+O+zNGFsbMxkXt1NByf4mnsmtbp5S9axIa/Nz
Tp6TMNT86i71X16BSiWnaQ0ecOb7YHH3PHTROIGUQ/UECqJsSXr7QiSNyRjT0bXBby5yg2dNnMEv
IcY+Z9zyBNGN+sr7pSIHz5HqPU7esEhFMkgYGbFPrQQci5wmvQ4r4pNDhAR0BMJvhFy8Y+oefWHA
SiuzU5fN03Di3HEK+u+T7ygOLLOgHOTsQE9CTlT1Q/aGHJXRVTQI3YD7zTiWVevW5S8qaDmsT6gT
nTnScYS6UJTfmFEV2xNgcngqVU49UoIh/poDvFV2JQTX76GYmg8b0XXaKozOrCkXSw0qgKrnJA0h
pOeR1YsfRmgKUEMapDsxOrRS7sO/QMy8BpgG1KaQJIc8MZUNUbFipDqJQCN+773dT+fjJwxHCh0s
8NHDoZ1JxeBfj1wfgHW5oE9roCc/o95DTWnyPnzjP2Q6jy/UoHgfuveVhnZ3KGOa5kCNoK/XM5Wd
i2IBoxvEzMAuG824e/m923fon/Img3bwNYENMU2Nj5X6DfCaYKFOGqRcybm2am/qfEhnKSX0G7uo
Kz6X+Y3OvLQIeMXclu1qGiYRSt016rsZqoWGY/C3LFWC+U7o7Te0M3iyyfqiwn1B5lJ4OzTcB8Pn
IjNJ1pG9z0VvBpKnj3NnrxW9VXtHFa43zxpjKxX3j/QU50v5sktNxqCTfFm2ESFAIHewzx+jpRx5
C1KEQPlj9o1STVEZBG9rVGin9hlrv8Hjf/yDkUrPTByZRi39mvLaB5ing5T1RM0yDMsnItPqC9k+
y4DzuXpaSO88HK9bEbrO3g5kYmeYFZaPUQohp+NRQBH21rtpFr1bsmkNnSuqvV9V2iHVTmzHKtFl
KNWhd9XkQZEowTIQva9JMhCGVRNE0yEXoo3A8PJ8lClmVQ7pOh66oA9HnY+WC4A6VrKGJOt7dowD
LmORRd6wwvT8wPO9in73tM0JeTY0//jje4Tzf6HRf/wCJezGBAzW84tcBCbLoAiN445IWgRL/C08
+Wp7HiZBGRy5NwnHQ6faF6SohAEJlsF09qQqscH4nUnsG/RsGikaJBLHkMRgPwCgIAXIVQzn1DpE
5soBCCUhMItR9x0aq2xG63N++OCefq+Do8A9FBqITbtwTEpVD28Z7+GICg7OqEMq0OlGZt0K1bzt
Xx+kqsSCT1R9vIZxtr1hxsuI8Od8SggqeObK5le22EU9hzjopz0C8lYm5OvBhlwkmvW0RY10RY9o
Go2yjJsGIThnvtQut7R1UrYFeYoDAMcVz7AOESDSVjPN5TudhTdAw0e1E1UF/Nh+5LbdHE56e4CN
r2YzpxPdFzO3VVR1qfXoilFVbJIzoZ2P4IaHScC0FEtY62XgFeOiW7efr9FBQ8N4djgMphU1tEUU
EJjaiMi87Y7atxNRLbbIwY0IzlpKFSHDvslpsgmYMvdjD2bo+AJL6B38KzRcEqHLiUMsi0iYWkp9
5NjyhrOCsMt7n/AvCWDGn1fVal1hdyR7a+tVMdHBVIyrUXJ0/egJUUr9vvVhHWUFelBLU9x5+44f
ZQH2eeBwzw67s6/zl2F2dM9cHlDIanHhdz4cgX+8DrB/ahjmCqXcxNKOB3kuub6HbqDINJKJTifh
cINqGQdzHKXyy9DJftGQmeWdyFSEffsUefjxrFDUHllbK85nKEo0V/Lt31DAb1J5YuMJCSEJlBA7
m8ZAoOg7Q8Qzb1ol97fkytiBqby5wOUgVpHwvjJSGOlgbAbZInh0ey8w5jcD9ZDPMf4sLe1fU3fj
BD9D661P4tIBNia1DwXcyXNbCJTgbtmKvoGp8cG33DenY9DP6pnynH1n4YFhG63F73FeXaUGDl1Y
uLNL1aoecqI+5WdgNSFN1dClVbR+Qo4XWoT8RuoMBHCq0CkKPc1NqY0DKpa/hvZN+jli6I1EJeBE
4DWfaf1WnqQXLjVA5NisUxnx0eWP/p7WJvdhJq54B8SMCNj13YeE4gNUrP07q4QC5lUT6I9w4/aF
thh80qsYurFE1ne22LXaNbjWFkXFYTUqteY43k4Ncsn2QXbrL2YRzOYfm4HKYdkOBt/sDI7M0Orj
PbuHNM6PLNrUoj+0hl9O8pokMbiM9aY7/y9wg+kc9K1hY5NJZxczTB4qhJYsr9Tt7vX3ZsVeX1P2
V8T3w3fjG4lHgUJ+qQ1lB354NGbgdc4tloa08f/E2ppmt/pRPvvjnHRqmNbrE/5irNUz6QZb6szi
oU2MZ05tYygnsCTLbFxMwavUdwiy+GwKfC9/t/eN+SyvrLAovGT7iwhf9z0/PYxx4j6HUeSOrLjH
10oT32eMZcmkeysLyPPlOauY9Lyv4Ppr6cBNs1PA66YNA5dA8ZAvynXxliqEfMzQp0pwtQI63TUp
JUj6czHY/+iQhOPKvnrlRExlaQRqfZ7lf8meuOBdiOcko5SKNoyVAqV8dj+TfZJRSHTqoxmduZI7
0M02HuZcUeUoxKWbeEkVWZikyUVtk1+ijR2qT6r+bx8lqKBaXeiLiVx4stDzJUMAIdJXk+V9Y3H3
R0fMMkemLZU+A1//fQKW0nrNsHyd0sgqPiN4CP+ZDZWHKiiKsag6t0mf0nVv/8BXW5ZqVr301phx
+64bUdrThRFSXvpd5MT9s/hItjkqyVVf+0c9LhEaY+TlNVR7StoC3tgX9L211BMQylxa80ch1ljA
6XCTKSO6XkRgoZmKkoSu8AhK2/vMxbuEmQVk/8AR2bjowMKmarht+r5lt1kO1HZ317W+/fEBoelu
3aM02+V1NSq1kX4cADqfm48DH9HHy2XgGqO6ssBdNfhc34C5my+JTKiUENJDk3zAMGSfx2OSlMih
hhuiXpmUC8+srJ57Wip/pQnW8X3wiedO+f+7o3ctF7738oTLQI7CXCx5WR8J0HPUWa1xB6cFdZ+L
VF5iROmhBNdgP1hiyZN8O2VRLGcjaX6411VEx0SHsb7c6Vqp3J8/I5AYMHp9D9ZgQdZ2V9VbLS5u
pRIWh2tCxAzyzM3eQlhlXYodaUiCUQSduzCgptAwWpHQ2LVoWD912meOAEugcg4es2yZ97Po5WuF
utapWzttD9a4garH0MWapRxrpjXF3WsHqnqcUdLCp7gUd/dSHYHIJBJ9zHl0UgzPMspF22shfiWh
9eStsF9ugtmOU2+5lW/a8IRjQmfkavRqwZzbjXt6Qf6CKMc5K6JKGc+ZFLXq5nuBFfO3mnjdg8BX
LuZzaXSgy+SXDMX0UMK3Meany2kVd8zo4OZ09mV2iZUbkG0CP4vfonIPw7NEig+IwVUgSEQU5edU
4y0t8Qo14GXDda7kcqNi4puEMaYD70uusrSdMN05++nwd/I5DLXDJchebOBEsq0PF1kLxP4busOV
Xq/kB/zoJIs799dIeNnd2VBbBKjLMh+giAf8owK0X9OMO+BASlrYWCR1q+FHz0kr8lpvHNIIfDk5
qunjuhIQGmsyob+rOavyNBOCexleS40pO+XPlko6GFU53OSyrZ/24GfTauXojsB0zORZDCSf+dtP
q4rTUh6/m2z7TpNBCbrZkML1ffueDS2BhYPLsykssg6iNLJfI6iOx6mavh1KmWKhwXRnwBU2Qg06
Z206GrRBhvoBX79/Fb+wol8RClcePoCyH2cvhGg9ebMbGzwCUT/+WrKyiEVtpOu6vGoTUcu8gr3W
BplqYb/URZk5un4TSiZ/OUGo9urhLo1FDiEQcBcxGeLCT84PM711oqhbtrOXkBY9H7k6Pbk5iThO
26Bizct17LLJ5TBj1MQJSPJSFBTZPyixWIC/Vv20uE4FRqF6+Dsm9TNliOpL87XILRaFcTjPoqeA
X7zfhBP6BFlosECJANVYqel1g1dyfFsJg8h5jbTxW4MAiP/VURMQtpQKTmJuKPEo0K4+0ZJggHTb
pdZ1PqUrBRprII4p/HQzXZTm8fMuffQhpQmnqhNaYQNacin2JTUbZl98G70+3XcJngx7EH7oSKYL
6UtExVDMylKITwiXTFsJD3mmmfCYPLtY7HuMomWcN4tvIHLOt3J5wbUp2JlM6F72VVHkexPdA3X8
ANQsfzPBFIIyixjVWbJG14k7g5K2HCsWhTS+USU858sTX1K1RmPQrZUYEnLGuYrkoISUm6NsF1dp
sxbV7DuXQSgp7TULcc8iQEGVkUj8ubvJHCdGXpWFEDzASUwsgJLJqvR9wBkyUyuGTE8C98za/eO2
mL3ofRyv9sYpKMeV1Q0csdTFj8UhQu8k0YNTwDaa3fkIuUqJWjoUtgE4HkygahiwqHulxkgepLd/
ulkTEZGcFs6Q2Y/KgI4JQ6RawDEjE9l/NvsQ6r2wlldctd+wwmJEsvZoPxiMl94gFYRlQXd4lq75
2y7CZ8Rh6H/Lv9/x+yyudHAts2BqkOWtPEUV+Xl1qi4kej47mOYO7GV0Z2+mGZDK7+a5ds3JCpa1
jttv6+kQq9LONszOeTdeT2QKBiReVGampiupcqPeV8pq43vkmx4lFvuc7o+BxyHUHgAs7QdoVAe9
js3Q+8s6nIMgHPpvSt50udqACLUA+FebCDi7uej4dtBVwATIWaeNmHzPpXwL+mxWJxw8h6PVF+m0
8A/kGdmao01xlK5K0W825SlTzGhqub++wUxN0ZHgu2G+0zg0mJwPIZWLNahPyumrxQX0cN0ha1QA
apKtda1a9zZHU06s3M9tyoNjAbyL22jLTISG8uvFIwiAP8T3ESP7yM5CpxVcUUwsrtWN6fFNe3LC
ZJqc6gXmF9AwCBjFQAEKvoFZv5C91HnORo1o003HATUPENG48mEl5Hix9hMCODYG6HI8UZs6sqoV
X7JByo4YH7XOsySobXmX1NufiLUz3ZMG3/d5A8bBrI6pSGqGbBlsB2dwcje0duRq2I2AThmvPYca
CJ3YFkJKm8YUX0QC6G/vBlFkHHMZ+Usg+7spsllppCNeywyYnLXXQ8I6qgyDLnugvEKndWUksTZU
mGm9GLh7eGrKdp4c6QIFBAnUCiFLgIhvU7WLBdFnaXeYU1MTkuptN/r8u0BGb6uPqfXm7dZjxQ68
rifyvXlOBrwTY8CWtD6vhsK2IX05yTP+buTi2ZSKynjRIORVAGvg47pPL44uogzT/+bjB/3A3yqw
4qefwlHCuilTxqvLZZW5a9+mZ4F/fLG6t/nRa0/AzdMxowKq5BmGHEWyWzXbKcftEbNnsrLF+TaQ
9QnvXkKq98HQeRI+T4qgrJMXClIXHZQ31bgOqEjXkD97DKnpjo1+4fieAKLO3Nqutx6Jx4oi79Og
G/EgUC0Os2rBpL79uqiUYHdeDxmuy+s7/7djvmvPgPbSg5LLLiMBI3cPhXFGpAuPUUeYqfqkQtUQ
lj6zKDdCM6zxoX8/hD3x+QpcyS9qAZV70epiD1tQA7cWEjCuGUAc4wlXzqAzmkSs9kM2rpjLY6Dj
klrt0tzAV8gP28YGxsyBHZrF/dA2dADE6o6ndHcDg8VII4gikvOej0oxKeVOXK8F1fvU4tudB8Eb
15KGlAdFz0BNkJuMBdMl4S7Ia+Xv6XFqb+pN/aB5PPYgwg3446cX15W6kxnaMexn70XRo0z6p2H2
f/oafYdmlRlZtlfqpwRqm5pXhhlLzLgUNwZqIAAknpG0hPn/x0e6OiGM7Bhe2b47qsrV2yFVy5WZ
5CvUahyIL2LZRMGQWwwLbtGd1nob1dYqJ80kDa2uZJbSlxVp1zfDY0FSLVY0TPVzicGzXc1mApmr
rYsWj1mGOD60oJ19LD+azpWTqPRdCFub1Pb4AbZpzuS1yLkx/8wrB3/m6w5a+5j/j4TjWAFszhOj
M7kzleA60QnLTw+cs5awNhAQ2CrlYdNI5zbDFkPkH6KTudaifkUsRtudWSmBKezyarYYhI9eDKFM
FbD72ri9B8PG3PP8A+sAEOGE1rrEr9xOiXkjNreHaVy1UwY2wmfxoDvU/ejVeGPNY1aLk4YTnoVo
Gcxho+fkiCVnXVbW/JCFsPTgqE92CeJBWRbOLUf+j/eRKW6WwIQwICzebPEGd5XnfA8yU5dLvcRi
RA6C4LOOAs6jdjzJOyd6iUdWuLHbApn8dr4pJGpszI4Z+Ubx5Yq4Co8lcvV82rClg6gCUi+HJel8
EBICdmmdBq22IML3DseqCcT6g635jvC03lEezznxLhlwtYa+yLvRJT3ZXN3uFu0zZqbn6h3RBp8r
gS+CnAHqwuXjBL48qC0buTtotUtIARoZQv4T2eiq+EWDkSWM8itkROdCCR5Nsnhf0ImllLK/Hkkv
++Xc0L0FU35dnIYSEuYgBlh7TlRhDzp2Eo2jyfSyHu+n+7AvqTIBeJKBDyXTl+o2SCcEwC93bs7A
MJW4w6/VA8gnZWSTRboXhQgjVJcRW41+PdLFYXY93gWffrWowTpuw3RrZusLk/WMFiOZG/IW9LcX
G+h8ycuWqbNAS8M0+c316185qf1wHjrqSrlZVE2QRNFupoyH/DVhowEFLss34uf57t7xbnuS1DUw
nSopTswXCG1mVLlfBNsw9/pSHHNJtmb2qVOafgV3jwguSGJ1cYN7HjGXIIAtdDkfiJ6LDxHyt0Vu
C69PQ3S6AnReM+QpBHNX3/Ho5J5sGC90ikmHymJ6CwMMmynAIoom7ZFgylkiEIVlHcue/RRzU+qL
FEMuLQMWBIpNYH+Vb4NlCwPX2mJrfLsyueMNuqFtuP5nFnWBBgGNxu9jMzMoG1Bg3amgnA0Cv6fp
bxgrZZchd46bpwFDpd0/2/KhHTIQwKSoz3O31zbQaieJJ5apI91l3KINKscnK+0+8a/cxeSIygUW
smzVNxu55HmzUn74oGwsRVG3iQay+9J1EmFA5BcEa2cZDMiQ87c0vF9TwCa/cwvY/93tlx2lcUfo
LMJf8V4CjZNbjUXOW93hVLv7Grxna96xsQ0yKYgbfUJzMPv0GKgFI904ZSSckbiJpftIxVUtS45b
nl66MVKisffLIMYWwAGUp9ndRQJOtTyImxfcAKDPfptFk5N9q5jjIjXthxl8cDYShu+2w6oFY+JI
qrr+6CrB205BaSb2Q45e4Rn6voVboO+sE27Fu2dgClzR8JxytlmFM7cQlSLu6bXXf9lv/z6hr6OA
/Qv56T9fBwIv6gl9ScSyhZmbzWUxcZ3REgimjEdh4gBq9NrS5L5MWjc9UnQLge8rY4qjNGN5Q1IL
BogpJGHpPMjrwDRTkfRIQ0DmXEK63YBNDxDCbD7FGTZELJHfvZqGhLLaTOYt15EXjjMIwC9xDzHI
vl3IWugwfG69JbtYSV2NZ7uK0w7YlsPhaJuBJYwm3VCGoV3bOBD2a83VIQpNdsCierAQMa4xIm3h
ZgZb5U2x+wzG1T6pA2dhc1UjWN9qTxeGL/nJSz9SMihMdLlIvBOMidaeD8o58qhUBqVyP+w3AEbP
QvkFawEJbgoWQm1x4BR1IADE3XFzsBzfB0Xx0waJ3knu6ZHcGVeproVmHVf39zttOY2tUl6PABY3
Si6CaiF7/iwPFEPOs9l9MnysNDnn1xTJhory/oMyZZdpkOwNNI4E1mQdd3FY9lMpaOGCL06m4RVj
bHd5sps8RaiMpk4DDZX4NZQqcLCk/W2EsTDAqvSf195w0oX0PRbww8mCauWmigsnN/82+1fSWIof
aXWSkobNaC7+G8wBx8Wzb6708TTa+rstGazbD8+f1RtjRs3lO56sZZF9ks2U5SQtXUz4zIkokd6F
pdzVMi2T5IIF1sj9JSr94jVS7ASuuL0jBF5v/2EYTd1z5zqcKpcbH9wybWBjbLxUaQc77YjQqsCU
qgoPO40tWvhQHBkZ9aF/bhm011+PUV8vfRBI+lRIQa56b3ZGakc4NOt7qnt/wufFnpqVX28IyZZK
l+SIRZ+W/x0mJL04SMQ2q38325BCjfNkUlvMFKcKvLodlZS2he0pLOt6G+7nY+ICI3pnWBbpb83n
e3gVwN8BU/vr+5Q9RgZuBMl2YvnATQzXbksYX1Pw6SL7enb6IHt1BXX5EUVtrGg1eDO6JFUuFSLU
hGObGdr/bWXHCUw9ux2QihRFOQ2BXFPHpCQp9vP3/hykZbTQaOepAE5EdJMamNuKW3tXm6zWrPKk
/QOTK0PVBLWJH3QTf4ROuxN6T4xKyPUUQy81/Su/5jRRZfASejla1sPM/CvZENmTCw8g3YNVf6qQ
fZpLa3vbcdLOs80Lr0Ua9KKXJ3vWLBNEPFxeIiX2CRTksEjd11tXmdF8tLMu/YeC98J6TeGyBUQY
lumeRaM5kTVUt3B2RWLW2Vq0hXituKANurJVTj3UYHgJ86CLPaDBf6lLfXQtd1J8wCAxHTORwQc1
PgkzZp6GfXH2BPL0lroGm0mTXe6Dvyp+fHAWmazRC3FWONWjBWZCB+oUSrsK6ACPvMRTHMEudp0K
0PWoozxeucNIr4rRCFb081b38rYeVVta8ghRoFE9reihXE4rs98hEOPpFGpUJNtPoVUj/wkniXjw
PP8XQ3XwheL1ul9vcnBr58NiaKDGUTymfN7HcNckzatP2mWYZnqXiLUkU+DLvUdHE9oN4QuKSIIV
5ZuKU7jkn1KmjUfrOB4UPEGvwbkTNC61EmANk7Ib+A0I9UeNrFvw06gFpSICqncm8VBg69eqsAjc
fUfoPkXcMeIXJu+ecnABfhifx/O4AnkwU4kLMOwE/XEA8QJyj1VQzNlX5e8uPDVRz3ahbYXYXYfJ
rbxsbCPuNs+yAhE5KcnM/j/MZTLpRoXcBd8kipTWoPtYBQ0fMX4oqz4hquxdJLROcjFnaPcJUJkd
Jh/9lwysNtTcP5I6nJDKmmqmL0XuTywNGe0e6U3FoFXokvtcnynLFziLxM4areYvsaPWLdM/81jd
wRAhyVlnO3M6p3OK9fu9KB/+GdGq3Z8tB45KZOdpl1JI2pwiqTwyFe1+D0+kCwHpGn/QLYweaDuH
S7jc+0cIQCjk2DP1LDLI+TaYO+ihQSI9LL1OHUXf5G77UxhU+iI8XhgYkVvKqsYGilcH3Knh85rK
xbOU5C3rdx2/X0D14iXjcK8KJhUrGEPIXIbfINf2Dd73qn9LsRyUYRFya1iuSJITzujMNVetgfsX
/zaIGC1Myutn74ZyYdXipXO098NvslMJ1oaqvWDR4W6qISMqfVPZgYsLdrLRE81bH9UrtIV3spWz
NF7t4x1cMA+aMi8plp9eKlcmQa3WGPxCICITyVGSs0uqBLN9nfoAMUQeM5CWEnEZhUuSrOo7/D93
QOGpf4jmBJ4ZHIZ9moMVD6G/Y7HxZt+N7BZ496zNYj7lAFtcaidyELqpLFR1BS5Mz6ZmLHNRSBAq
K18m8g4seJjxOloZxfVNgmLgH3wbtsV1GaminCP1GLm5E1ClQv5LTbWIlOnmTi8bG/ZkD9Slve29
+94imXYIlzv6m49XCOXh8pTIXykYx3uYshbynJ0i6vNmqxMx8nup3M90v9OXf/6Z6LFvU+kLhZtW
dFoOvl7ogWK3jle+EbVmPEMgN9zLDRaqU6Z/0prbp4y/BdpZtIBIHlmV9b8tXPV6e8j8glG31TTB
3HIEu3GJssb5g8/QsCDUujzzWkPyDZ3VjIlT5gM1EQ3fndgS+F8uZdFipsgCYJbB8tV4aU4suDqS
4pnQ8iKnkbZFQ/UIBxM4hsd+9r14tXmd8VUDcp3Yuyx+yGxwG1HkNKfJLC4l0dEqO2Wmv7k7sy7I
feXRlALmDwFOYxtI2pJnXmM1UL2Fjj0UBLDLygHd2HqFWuwvpxAco4RJI6fa/iPA2xPoGW0ZgDtb
zpeb8JXIS68AfXJ22Wq9QG1tfTPSRKtmnDNVvbtk4zsEO550rpDtRXC0ZIA48OqUnHnsPm5TYhEs
6mnT4bfwp7kVeCryDmjwXrQdObTSF+H5RAxYdCavXkxTpFdpzc1mcBjbwRu3iQymbsxKPhTHeU6b
kEaysHs3tbzA88pLtzDZAYZenjUpQFiVR6OHM1FJe6Nkxj4a96wnU7nqp4QQsN57k1vCZPqLrqLo
9l7pHpuvtukA3PRt698cDb5bfm9ngPehYY/Qfc5uanpYSW+FsfgFhWOf31olLnyYLh7npUEKtgUu
Ki6T/IhtVRD7fTt2CJbXbAyfzARB+L2vglZ+llKb05AjabU/FtR1DWOEoaNjwr0a14/qd2qP3i4q
7gPXX5msLeRfiFdWSp0sOO/ImnwPijDXTADdk4o2/xeF4gs+ipSHuioglMcs66a98fnPCbu/01wH
gLpUqWNFt3U3NzLCvCqtHOphEGRwvIuPqp/7rD2Ne3GP0EA5K7d6UeouIh7b8REkiQy1Hme6WA9L
EaHNnfn/NcmbAu+KG4sHWU38JYq1PcBs+zaJA/4ECvM7VgYSvDOjL9aDxlYci9+xOUJm8hKkoTfe
9sKJTFWuOQsf9vIhq3ulRBfcymaYwPDhvRccAnQUgCIgfJidL/zz8Pz3XvGUox10WGJQGYvTvtag
rT39gIqrlrvHZvDBsbZ2WGe3xO4BVIFwEbtnzvnLjwp2sKjgG4RL+iuaGNxGnXtm3+j1lTNHi4w7
XAPdYWYoNS9s+i0BZiY9z660l3ZAScwkYE5JNN8W9rDDysceAVE9gkipiCPXqkHh3gcatO8n9aoO
kROjZ0YjjZu3h8QfQ5GXU0spUpDn928Vsj+SejFj05PjYa/6Wfi/9qHj31WwFoYmPI6vRgVxrHgp
+HnLU2075vY1RxDBCMzXtax3sP/eQQjQJvX/SlRTicbRpza9I1xK2uSThym3gKrC/G4daOq0jF8M
o18RFKrDisn0oNPjrYc5Pa2oyf+258KeapQUUyTxEm79hkD+GI/wQn6tgVKqCMkvxGGsaeT5t1mL
Uz0uONW/Y6eJDrRKMTSLBq1GZodYzZt6AhAE3qlERDsUbQY4y1FvswFcGBJwl99L7K0sBfBXDpjl
/KePZIZgJDHPoOfZKldnG0/svqdr9m/HxSVWFnRpskpKenCTgftI0SwSgkxxejbzy+G+vdznAleX
t+bnuq8ak8t3yTN/jm3LLQTbEZ/3cKNpLE3RgitvhpdUcIVQsKMymY8hqXMdL4kzVqhGO010xGpH
KfG/UjaUE94HcMjAok8l4ve5bDiIeMqS+X2aYuQFuWu6J8cBQPWitKSupan7TYZUujxMoLPhEk+3
5Uh0gLmP3JdoIMi94AZsqhCmnRTYT3RSJZqX9XiHiFXwH1rOhDcQrCnRodrwKncDoloWz2qFHaBQ
FsymUaiX9Rs3vhjERN/ifLZmHlda4FmxKPa7m+K2f2IffiZx5tSe/jnk7nGGJy51Vsq2y6Buahne
C8TyVXanA3qToB7CSCxDvPEVBDki+4MgIWPw0bEv4utRAfBu5Gp5LbzEek+Uxj4lAZiZQY9a2Rx8
ouhGrCi8rj9110V2ch63I5fmDmoczp8bD+ywY/y/B/UgOXCzRVbhEDLBYSD2D5NUWZ2ZPZ1mxw1Q
U1UZtRUpK/CGk4Cs57Byl1eIjes26Um7LbjUulsJ40KHMj4bqvR3cTVf0+flYaQPuNs8ZJZcXaLc
UxJflQ1a1NXPNduTk+95YYiEhCrgcc1zPbruNyWHot5NCDJ8PIrRe0GLnAU9c9sn17ex5oWoRlF9
aM3ygYEa8Y+e5bUZ7CeofgTfYCCGYQnmvoah+eE75GjpzpwY9DITJyEIsDh852hiMkOEwpbBctrS
llZ/2XqhU5m8XfdPaVn9R6jgmY4+8cguS5bEIfHPdqKfOpea4dyj8dVbuwSZJr4wl5LukWQ9ijGv
H5rDQ/kzOdig9SpLOmYbA/ErdCyAwsYA2UXFnNApwK7ZWJvWl7oFFWfAq5+70rV8CE/LxOTX2YQR
KsXyPV9xwHYTX36k877Sefq51e8EPCV5fxkMxaM1oWbfOFe7cO2Owsl8eHLEH9FfxWI9ULQmT9A1
EhYrA+APh8P69GW2McuLOMnG1dxL3nQtHMRjww/EnMN/XUXmkBxMI/Z4veSCvUaJcIrnMjGepNeQ
WTFtfgGLTBmP6SHR5U/wajKZR1eAH4SfMHqeVgijaYWjo57J1d3rVKVwlxoLpyRXoF145Sr6a0sE
m0jYQbDQkCG3T7X/3CIY6RGRpz5zLhIqH5Vzj2J6Em78ZbsSmr3s1n6486qDANHjO2tSV4vUEdf5
Jrb9ye6Bca9380uKyC+3Pir0tC/w8OxMwXdkQfi+75+/rt8exp+PvaPH0UP6gNcci2y3AD9k4Wh7
eYGhoSnWcpAQkgrxyVyPgOyT28CGbJGOPzDDGViYbi4BC7OLDAm0BN/RFLt5EGMJBzofmxNBjHTx
KzeMt8rm3k+VdaE+bQLj9QP/E1PPh1CvUmeYFT6Idjpj0ewg0DJXM+SqSmgyYjh/xSuyvlR/YvGN
NaQdaP/+VeASvQMilqAtRa5vdNgqjxNWMVRQzebnRs9PebU/+QvQis8VJyjKepN6GlV2saHayFZv
DJRsosXeegV7Loh6RdQ/7g04pXCjWrPdSkM6dPlaIaan6vxtqZAz8AxyvUW0gMsprxnF0ATXpm/H
3aeQBwEn1+o2mUQw98zUrtb/U+wW3aAxPg0GlYiEdiNnrThi6cvvuU7+iZwAZP9C+O7BGye88DwL
+KPY/h4dmnLfggabGrSznTeg1wiXbccVS4xYdDFCKWSxNbc4+4DBhHDnecH7pm8CMFDolhU4N2ll
KqFy4jXRkwf8cH3XyO1+v1xG9I0N2CrtYAZiYa3O7q+RAxN8djgV9mIjmi/U2jLb1AsbYyfyZIuC
nW/UCUMRhko1VIjZK0iDFaQBnqnzdbK6/gDFlvZ8loB8O2JhCCGW3xRIYrkVEwIW0g2ECOLvU9NA
3dC8dykvKu+6WNJoE8BaiIVjERFcMBAOPpqNgqoF4pMsAL5OOS7bAJJSz3822JPyFnl8C0RppDh5
ZKFA9RIvsimVBpb6dSaEsr9chKktcsiyKb7G9r5wf3Hk/3C4NUDQRrWrBJiUrWmAhHPRKliLM9/Y
F57csdLMW/72oDs2s4SjZbXy6S5CNGQjC326wYM2cTURTRNKaVzyIV9UO8+qgt8ynicUOmxJyCUv
j2xjoIzuQpNK8AtcCQgRApR4kyHj8fj/xpPLl/z6a6Ana9crTGlkEgbXCnyjArq6LxTcM0dpoWik
whuV2Q1Z/gISDsvnU3r6+VztxN5XZOaDGCA69OgCiukD1baqs2Xm3m9j24FP2FH/0O339wOcmp+d
aCz2p66kcyytDDmAQ/d5R+GmYoTVBBA0p9DdumLP1dP6LviBVeqmIQ9RwMEUrrr3aB6+h4Lx+b/D
gC2gzFhAiBlgEA9Dr34OBADHX7pD8vLXMqrT7Z5VT8lA4pxbFTmYK9iRuEeSEuMZiJPSosrAnZI+
MfI68GD19ewqJZ7jgwrg+sTvO4jxA4YZLvlM8xXUQopO3zYeMmdNZO8qWchLXU+iIBwlGTu4ukJp
EwqK18pYkfBE92D5pYK2fDyYljFBK/TQP7mUg8jrqKXJdjWZ95eo8lT/Sqp/aFe08JFc/r0XosTR
CQ3LdBEuPrb8EG9XzLs0XZDqQo3/gJDf3H/wSNyg83dqxoee+RnkVVbBzi3KvD9N1YXbFmm2V1jI
Gr2ZcZET/uJ81+ojoc6sa5JdPAM6uIzt++GDo+dH+zl4PFXWPDq3GyWuXyzEztLux0Xtg/pJs9PC
tE0Kz8Fw+NoZTt6EpvzHYTL/prerliwaHi440bXv5M3YACkBY7VXV5MxXpYlv9DIfFsYK2ju/HER
OxAKlFzrPz2nf9Kz0RYZy8q3vUakcgrLYePcWn2D6m59hH8fBRvSS/S4Jda2RuWJkKSGmq7ZuJFg
a8BMbkV3STIQiftAsdOdvyfcXMW3NbAQi8LzQwGkov36BhcpEai7t6ZsER7a4ZMBJHqLMZw6k5qD
At5F2CbW8uBNMUMnX2HK4kn6jWfEOzOcaMk8iBvT8ISqJvtS3AvfYpATHzturRnL3pIJ+eceMQiw
5nKhIIcsidLkthI5fL6PZ3m7xJmHuDQYtF+mHnpJWgcfD0ozFLa6lgSpmXMAk3i/vYTEfxlC7N66
S1FIz0U2SYa7NL7sRX7nWDzHI+pK/c0qg7lNXFDgwqZ4GkbAIDsqH1KQfTfy5kKJk72Qutqgd3K+
5UKKeMEIQcqpxaiyNgVoC4PvP2TCFOq51Oh3OosV2e+f5NbWRh8akf8EonlGCNi8gHjvcrWlzqEn
Oatx2zu/fSDcWEOcXQW0G67xhE8j1N7tMt++2ht8pKQwT7anJOaWEFHaHrxAbfcp3cE7rU/qLFkd
tPBlt2UR6JnuP18KdNVk1pNSKreGY8FwC7NjOunRL08gUBg85PNMxymE8wLBT34Vesn0C7S4fbj+
4aW6a+sdjP/x8Tlr4lhF/7uipopqFEvMKnP9k/RwZchTyk50VDFSjTDoChPuu0s1MhFzQc4/gZhf
ga3fCUtnUBBmfPO9w8ldHqaoyqOuKblCsKhm9Iv6F3lFl05It0tnMOFHPpm9HzcRW2eoiwVCDTOH
c1NHqLQ9W3P0EGwR8+XVMyWiPnaOT9ASkItnyihR+TxFVufWPX1wcxhbY4J2b13Av955BOcRf/ub
yF9msy6H2FI8MFa0/Rt4anzF4MEnlSVwrL7hry6+buAPI5R29X69teFVNeT6H/NQOArVJGgxFAt7
JkA83b0lUbv8U734mJ1iQSlZuuPnY/JYDemy19XlUX9wXHga4af0iheUA5Wbysoxvc+3ov/XWKYd
Cns67+0vd6Ct0vBr9AmTy5m2fDwSOrM7fW/JubPRSDRzQ+LgFac2dzvH//N8NEFIqecewRNOPmMH
SBjAV//zTEBPlZ41w57gJlGSXWh4dwMbC1CqPUmdip60xorDsBRgoB4MN8I/x9VQL0tnQrBPIxBe
Hkqz9FS89IoQa+G5VP2c7SWa6pYDzHdsNqgj8eAm+87u9V4SgzLU5G3m/9kxvCey3mUrEtEdjZev
BbebKV8Tjc+zZ6zDFXZNnC7DLAK63sBtIwkzeHQ2CSFZu6ePHM1sLUbLGUCIHOrPHSJJV4VRGpTq
/SKGcEz/i+Z9wyxPA6W1nqnm27daQaD/x+y+PPLVTZnZqhktovw5fNXrqOf8eFhRlzxTchMdxqym
x5RWCEheMhqTi1nOi4NG4zI6CjHmb5aiBmkAEuNo4avuEEIoyLKFH95ZEcaqZWOeVfWYWYCJZ4AO
VACaHjxufgG37z2oEzVkM6i2XUGbS0AJKTvZEnqTS1GuRTrQFZE5LoRhDK0gqCqAlYurqI+djyPZ
5MmqSykv+y8wD+qX/49oVzDMLsX9DmOh9GeEk6gSyWHLUblT5Y4Adxrwl9GTvbITNY+im7pCJTcx
w66GoHwfaBFItUVVw+QpVPPwUnpTQcVwKR7/mfZRWFxvrRmMHgxIYbA/pyJ+yrL9oMwlCva0fMvp
YTOUr9MDjk5jfApKfXGkWSwkZrsXFMcVx0DpXWCrBUrZ+CWAybmWxuHlXY5xiAqIOZkxsJ7/Gjrg
EXI+JaQ/Ti5BYxAcxY9H8TmpfRPuVKr/1GTcpIihBCFytxqMW6zbAbwtK6qRVRZYvksiY2vicZWh
4hIFYZ16vW8vrKADHQEa0nUDMUAyzlS/dP57oJhedZFDDPU2dTmfXeW4tG4OnTkNeKgSz1acbu3l
PTcbwDRbA2W2CQW4JeJsjY9r/K1SJzAcBjOsH6PyGxLuDlr7n/GcCTvZ/4kkmNgYyVgaUCJhc8Rv
/Ao1nS61qgIGVFt9IWB2HfGdLx3SE/Q7dh+cHzOjWsErQETdgZWO4gfIUjNB7i7ONqb4K38fnmzc
yF0tUOJZHLNSenXXAnW0KuOvMfO6CO6gMNSfXi1PMQ2/cL+n8GuU5CGeqJUHELftx5pSLu6Y0nu/
KL3BqNKm0VUxXMbtyaeBWU1nuNoxm1QJJLShuochZD5tVgQRVnyjTxVr5MsKi8+E2rmMB8HUS9CH
VBCcergg1C09pU0tkVnfglL+2ykhamhSL2Qwpdh9ObG1rFqILoSJhHWmSWL2Is54AMeEaUGQkAKh
6DcOqMcpYsIMx295WzOxDvBhUkvfZFx9DpUuo0QUVR0z+c+DHx+QL/c1K1JlzboANXU69qmmPsc6
HbhHpP60/lfE09/k/UFoajPwUYDI+GMeELXjcb7q9oJnc1kOwZjKhshhOepDfOkkm8old3j23yPQ
uKgqMM8iUUs0rxopKWrMUHehqxTe9hDIGpdltuXdF1j+OhnX29w6e/48lbB8q8WAjttZzNiQz/bB
3rG4cYjLiCaxtGp5wQWxVzcw7A7D0zgtp7d80v+sexJg1fV5JTK0o0qKAroYzW1S4q4dN0xu3cNX
771xRt20TNyZ7uLv/WllywZhGYd4Oz0O+YnyR104QAQGv3rTy178lkEDBoQ6e7c/TqWZX/Ya6gY9
DabDK/bmOY040CSnO8z/NA1sDiT9lozlMo6Jb5RiPEaBNKOgHdY2VIDQJp1TnbQ7LJNSLbF+ciDT
MqiJifH0OLFTv/zbjBKQ379BSa8HSU1gb3yO0r/cqmwCeXv8NRf9VWUXvVh98L23wpYzTZS7/gGv
lum8s5nQiul+2DzEJTccY6EBsB2SnNqMBpRBgq83hxLvVLB2T+Txe0keBHLJyJUz76zxz8pERd2c
wiAMgQ8HZWuiKqlGym63cz7JpDtTqZoqW2kVJPkq9YgOSZJxGhJ9sHga7foi3iCEWWrv8dQL0V9m
SIGeGPxcHZB+IWdTjXNXM/HwhP5b0mpTjtkoRB51IN4Dci0zw124X9ff3tUL8PpBs2ftyaE7f4CD
Y6t9XGTctFptcRoXmOcuza4tiiZpxTWlnnas6fDL1UJsMixMeBhheLw3MZtk3W+cVc7zcs6x0b07
88nkVlP/zyEL97/6uzZz7ZzeABnQgBj2m48Ms6ehD95ehZgDUB5efU+Zlkf+VuSjn/WgMLbx0A4d
jsIZOeXYBSrsJt2aXsZzRwq/SB9cTKS64CwfwpW+Ih6Je8K4mr6sCCKKLwixyz9UFt6MUDQhSU+V
HoXvKvnYjoqN6HNBnbftAHBpz1z4/Os5zP7Vl1Tn4ooggFyKUjcNReOnSC5Yb781OvqXVaKyFO6p
DxmwF6oxyDdATyLxVk5pIfoZHISnzKxuwmRffwFp08tg42W71fdC/yvaoBXkVUQdarGoc7z4t94+
YZ664DKa8v+twob38XtukMPJeZnfqnRHiuSaSHrPwqu7MxmhTo4BRpKyl/Krnm8dB4iUZZ1d5o+W
NgHxub3Hr8vy89TDXluhkbwIgQWveTr5qyxjQirg7xUSpB7nbQPMr6jwugPuHjlGiK0/UEBuBfHp
EQqsCVZcuyjAHdIUNtmpOw5sVFu3LKliBvfkVAp17Om6ppXwF9UKYtZuIU9k6PtVUxv3jQp20b12
1mGBl9yybM/qrDr/nY+hAvZI5fTpB2vtfmvWprAFMuIWqBGaXU8eUV/uneWVgGRktjTyZcgAyHY/
WdXBPuTu0JetSSUg5LvJNXa52Z/jD70TmNKN2CPY7kVMs+KuuaN3iwwAXi1ctMMsjLodcNEM2wBz
eJhLS/4mLcXYSi8Hz9aQfB3M2q444Vz9E7+ip7AVh22POdxKrTV2n8lf8PUV85FznK6pKNU5x6Cl
hiAew4lioPvvh3Hkr7DWKVa9oFBQd6hkgsOYjeBAyZMgu2siPaU419Z0wEMywNb6mNcfYDlpkxvq
8zSJNBZopqecf5DK+44zn3/EADyNktyKkdvlVMOdPoFirHObCWwAUOc0DU69X53N3LYwGltfa/7J
af5uCnA6EvA0xBDTQVdTJ+AoP5GitaMMUy6/RVUHN9l40run4PB0TzW0azypXcAIkpU8Mu4lVZc3
GZDJ0kQzmKfRkoHp4xFDWNACNyVfeBrtmav1X5OxOC4Yh1m/ooBprOeZljm9FzifM6tyLZRRJq4M
C5iHHqT8vp5wHHqA51SFvcC/nULxqGf8IWOUF/cwcQfMxl8Ta2b4NbMRaJOxb+16sRtYUJTOzGum
iXQwkexH9hriZ4tZ2l3gXHpJrUf028ZCNMU0EPskR+kMfTVvC6dDyDVw0F+DuoY3SSh+XLYLHeLR
KXsGrZoiTPpNogl1Kw6XryNvX6CunstewXWrDKgjx1kdkF+AzQCRXcQVE6fFef6wTqHtFg7Qan8w
PXcicaHA4dsA3AxbD5OjN+PMUzyIfKf+qSkelMBWhrClEGsefdIaVna/HXc5Rt6RJvPtXp7O4HnN
DMoeJvd790vfkhhu34JJ2fnr/xS4BGFRz1tqRX7KL+SwRHoVHBPJVKTVe4wXeI6RZnf9YW1vDSX8
S9WL34m8dSjX9K4jega0i//H6EgeHVDuP8qV2Lp+HbJRFMWueoDRcSvyGfGRyZ2rSzbzIRjEd0JA
kfZkb5O4weZogXHbNPsu5Q67RoxANcQM5u3Rs2BjRuxxe0sfD8jXM9fBrAldlmdyLzpxNX/Y8oXx
bkuv9fpW4xa27igkq8vNgLzlzCpAedl8PVaxw4TBImmR0c804EdHd/sP+0gObeWIQ4rHIwy5s6tl
/TqLAi2VolS3aUFvxUK+zAp9CtBWF8ILQYaRX3KNrBDmH7YG8iVgluHrl8Kp0olJPjKVDfWFTIld
Vx0hJj1BFjhQHVLsp6YAWLoPx0z1KyERU9gLWN+ncxXtvOEM2v1x5aY/U/9bjJap/JOKqDl5AtHe
UVUjbZkfRB9dpMXVg/E9Sd04d8pXCKjsOaJ7N9ybhyMerWvUdxSwgIbPMYPJeXhskANh/LXoHv1q
9q+ZOXQoFwHTQc8H9cn5QM7HJWssyFVqiEzose0HGl9sZrS01N5aJkQA8B614ouHEKA3l+k8nRYK
VHCycVCwB17X1hmD6fXNlxJj9tdtJnB1Jd3sJoq6Gp+OCBtTyNT9y6m0B3ArxJpDMOc5cMgxUwIy
imwPKNDtpg23lrCBR+Ee4vzN8OTQPERNMLqazt1vCskQC9akkDRChKcOvw+OTFRhqzOIS1SjHSXB
aO8j7SYyAf040INMbF9pMqeBhIA/Q79id1ejKKdkT+VoYkJfGEe2hVGgEMBu7Q7lM/SFDypNrA5s
7EkfURoRbKKfaXnZ2470oiUsSJm27hT3QamrqFLKCjTVaMBs1XKojBd5Bi+anSyyw4F6Bh8Fij+g
amGivUfFEDOsb71vY0p508guVVbpvSfZNolv8WS+03tJmMSVDi8ek1lYtojlSexsElvKsp4Psqd/
6z3tHBCfm05d8YT09h+qZqdup3c5fhVf00IhFUs/JLhJHC3zpBJEosoZn91K3LwEGp7YNxJcajzF
nblTGkSR8Ax8snpvDNNyU6jhVmifCj+Ke7V2QCb2AB/N9J3OI3d0V8GxgPU6xFXD/tLHTQ742JpN
UUbpG8SSqtdli4XrkMy6SNDvwcM+LrL+bGhp+FKD8ULBdgBKlSd2i8wDMTCe0FKRKEVSbmgbgGL1
OkbhptKoMBwOzQ2MBAwCF+TtdpyLECMITXyiVQDXPpQioL1hYPx2F5bXIYpiBSC2XyCBZsHhhqS2
QEVCIFmiAGQ/JpoSeBdiDM05a8CiXlZLzL1O17o7L+8NTnxMbeZuBBjqasK73oKUKvwumGW4/xL+
6DKwgIfxcIjNuBDwFdigUwMyR3BR24A98F4kZTSbwzqam77cCNuekkv48H/xIscuaga3Gi7oPfpO
n3PBuPacIDfgBdxvsoejSJLi2yhs6Oqdl6Qalip06frDuMF6fl30OhecGcQdhPzSP3npkKOcGlrP
XaoYoDngUqQ2++UdhLWLzRyj0ISGF+2M4dXeBtIN7OTbDZ5/XtMA/2LL5ByKW93123IXGrAgsPGY
IR068m/EfJ4/AvvUepFCgNbF0utGasXf+JaEX2RNt5BVZlTNr6eeZklmUiPfBvlGzfWOGy+kJhUg
5lugNFNlbjpGYoYtTlZ6vgsgv5Ie23aDs3UoaXqBO/gsHeAblXkgDpqm5ESDI9wCJHNNilchvrJy
vPihzFWgeIlvp0//6wcnbyEnJZu3f8TsP2tDLZtB7IfrBiPWPJq9SxpBAPlgdvHjfneH91k7yY1i
Um58AOK/dLCQHW5B83tJBVIs7WlCBazRgqWfqkf0czkSFLAT08Al3wAOzI/MBUYr62nFuvZXO1wN
5KcaeeCZi1Bn/hTBzZMzzJcmJYRpAys+MUvmt+GaAdl3xqdlnpeiuvpUBkuUeBOOMNYPhMTqLYcG
pERhvSG/+81/vx+xNclkwmPGPAdI+W7UfbuAnnQ+bXdX04dqQBGUtDBcgD/0kpz5p/EietwNeNHO
nJX0oDKNrqIZ1s0EbwxST6YR+V4k3thJ2/83HqS3GFY31VR+jJmK2pVperaJjhjSciTYI9Tt0+e2
CYtrqFLPLxs1a7/aEz5ZTy30IlxK0hN/mzrmKCYxirTkgwia9B9YMTJ+XJaDkqxmvnoOzi0f3lE9
xkhmdts793SX8iwxJ0eq+JZQpXMeu5K/uZEyNUzE4CnN9hHLOhDXIm9Wl34hIn4QIuE+0xcC8+xB
EZ7JUMl7n2bgWrmkFjKAFG8Kk2bD3zEiNEjKsMGViBUR5DUe2OiVvvGwTsnomA5MhfVldeB3twHw
Dsu4VUzaBZ8DBlYEC9ZWdszYneCE1bP0VGvM2FGWZftrvbMQRuQUeUxoccnYA2PEgcZMrIo2tO+J
Sf0irXAQeNCrMwZSsMrQrPtGLe9KMn1FD3H4tb47ON1MlA4xrw/ftC+B3bxYjjBWqASjJL8B8c26
CvSDL6AjN4DjoYjqnvH3yoZdFdn7f65VuvZwUtJCs18tRhr8InGkne114gn/4NogYyFFlT85epIx
WCs5VAly2GvDWaqxcoAf9taKr81yKNBqDvq0srXwEOdtuQvs+umrNmuuMKAYXMg4wmsYURvLztFs
rogbC7qUOMeMGwQSYNcWOfDDlwqdl2eNa8QmGXJhiTUDRN/pkPv5vXxydKmTTVUTvgnkHDsWhL51
J0cl/ghdFaxBb1UX04f1TEuUFiOMSCNB44UAEcjsj7a5iWwH8refv09uXwPFt2tIUJ8yRxWBDcax
8gKek2dYnmQbXUEp6P/yfz/iaTP4nxMxMYMK24sNH/7m2Byef42sthr9atnYS6Je7VByS4xtvypP
sXxorJJd/exZIJ/Lo6XAS24JmSYhCBh2630hCbTiJK1h6fjXxdRPh4dPTd+5tyGjjCXOo5qSNAc5
Hrb1J7jjWjw/NZeFVJhkRmONcIUEYkQCbUVzu9ZI3g4hgcj99dzmbSJsisfSc9J8SsFTg7iDttv6
C09XNKoHmj6NkGsXUaM7I9WuwA5bqrO+wIeRectTJNwvQdU9pjwJF5iIw9c+Mxm1UildSsvEPcLI
KYnZjbxLH9sNB/QVV2XiCO3AX1ZRzG3ioPuijKhVJYUNyZM5cQSCXK6PP3pgUdHlpiOSZDMg1YHO
lRCCUjVfzcUdPwUCB9QSFnhwW57NoBe+U716dXBVa0dsiZx8E3eernzZAy2WN84p7Q2rF/5DAGmd
lntVIrnWUKY/mg+3yJxD5Q0+oyWYZhTiECKYS09i2my2NhCBFYemrlyfC0xy/FAXs13W+tMAr2c1
DxkIEW4TIHka59ywrNk2WakHbcGtbftqlznkDSYGmVMdAljAswdZg7vzoKeWC2P/j87Iupz9U0Ap
iPuI4c3Kwdve21RZACtfGrFayylReYs3TGl8+hqyrN6X7QbAa+HubJIZbK/liptw3QEHQdRszEEe
TDGMvjTCzmP9z68YuqsuG2AR+JwWa79zNUmgI4KRhSypHiW20OzTZ4bv24ByWbPvSVhKNMQLi1F4
DAchTg+X8qUBzmEqoDO8Sj5uKtJCuicg+JV76ro5eWbvCfz9fFJo2FSmilsozEDwfbIbNJhj+CGa
HhhEf0ZekDrIc8odRmPqFvBI50296P6OBjftGK/PnrE2w1Xu9lgRi9bio8saWL5+L62TnEHVAkGJ
ACrgSc3CHrubzru4INyWWfjORZJqTsZGGZ3z2vGDp+eCE+s/HHaX0kHcBkZg9bwzEZWRpxX2GDd9
X/B+D9VPPx6Q+GGmksfDkSViLENt3NlnOAb97jplMsDKEZfNVmu7UgDWBQiU1N1rATy0Q6pYcdYa
WChsakL77N32qsrtIRU3BaJV678zRWinXCq3wKKiA5Nwzm2g8tVUwGd7jOEaLCXV8o0hpQDMX6R8
W5HMloNLRMO4UnY+GhJNMBxbuE1zEOZgYAk5kgFdqEaqHBo85yk5y4yznNKwepsQxZcbub8hVeiw
J9Y+Da+p+ujz8yYEQl7+5g32bVHlih+LNBr7eodUuRlXmu08Ezx8GNV62aJtTs7Awi52cmmiWTJS
9f23c1+Lbm277hheKNWbShDWvZJbA2w2Bis+416IzTmLSwESJT6sXwAi8AvPo2zrRYmfXJJYQz+Z
dNWrT86X6CBV9ANxTdyjTc1FnXnywl2KCdx994SKxJfMHLDGfYiZnKDfm8vRKNyJ5ne7mZCGWScr
6FzSZwLIAXR3dH6cJODxE1gfmiFXzWlrQVVhJ3GQY3g8GijzZsy7OigSNeYt1Y0DHZ7+dLkcCdNS
CuXoQLMn0H6KBAMs7fjNl1CZSnjz+FtE8V3vC7YSpn8b2ZI4VXSsZLUK9Ss1kogL8gISYTsK/Ori
MpTjAG6oZ87T8HPKiyeSj3S7yODKI3jZwiZSt3zdHHbUvWYLEmhtf/mi0ZsB+4mvCnX/jj0PBwL6
uafj1REYtWvpVDOsRpJVztff6TyZ6Uj5dxJz4Nj17mZisVfCcnBVaV0JRri0p6ZR9ygTit2jTqP5
J96cycVX3vr9XXrQJroUiMZI2lfRLWP7mg+Z7r8xYa4aYTrL6Vz8k3uZ/IfbhZosodvzXGTNFId5
QkIG9B7Vv/2wZsvRDqlCLdiF3X4EOj06pUf6xBoUg/R55GGutxwBj+f+YsCsK6qnjgGA0+G67/UT
4qNWABWgsof/ftILyKbX8FmTCcUV4ArVIGdJ67+hRmUd1shcrt+1jfm+ZCeW7JldXHrWMkDqomQu
6ZABLKGx03vWnvuVu/VPq9wU+hQdT+rtp2SBHGhZd5BC0XBYmMh2syiJ2dYDgtcf1cWSeSVciD/R
vaYB7ro8BB+Rd/Nc+3FLx1n0z1JC+hiooC4YymZ4mrWCkrBpU99UQlrEl7a7yW8woLXAHC1ZIlvZ
bjKrgk0iewbKS2rdNL4D0LT2eJ0/STILUWNdPQiAf29seMKL2rwJjz3suvl5FhxlmAaiBrJxNwXI
9NfwcLNW2qsR3O1P2eacVU9rakSN9zqWyZIIu51QQHokAPF24+QcpJCyUkBw84SVNXgSaGc+A3el
MnfsKEZEJ48guvDNy/VLYHdJVBGwwn+TClR14k/y4SZj03Ox8NQbpfcSy0NdxgdQGKZvvbPhZ7ai
HWeBALeR6f0FedRoQGxdwxlktd4S2zW+Dzbc9Dl4u9mk9yNxvYEuZcj4xwPd1UPmtD88NrYpuDjJ
m+7QGctlwRanxV3uutwzloMNjC971syzaPYdLQo1BXGUtIHPhJGqXEDTkVsR/ylKm93QduOxgzsF
aDHkIRqT3XPfPVMIBroz28EvN18aJxtgramwkqAN2WueFE6iF/h9QCi2uV2bQBgwMbj7bkpml6Sm
5wHoRLJEVK///6lPXTK/QpcjQkK8xDDFOXlgNXvtR4hfGIJ2Q+CYgjanVKRjiF/Syx6EWsuNfILh
APM0byIb8bnFw86KX1R3yOhc4w9v7jQ8mJklLOay5u7YXhgkJInRnBoSr7XZNjwv0xk3iJkxBimD
XW6RNyFClqb9UPsSLbYwJloqopYAuMXsGDZbmwd/Y4M5WIO60flE5ILR6fbxhARTAT3yzq11Y068
WeCJIW3PLfNbKMFH8T3gcuwKEDzkrrq1VjMR6g+3YTjsevFQd4VvPsz1B4wWseqd1BySh7DS3yzE
EFby9qw255L86NGOhEuG8wK7VXEeb8rAA3pj05+96D6UwyV9UvBeY8IvKPMu8kdDsc6dVkOunB5c
f6Lk4B4yMLlY5WyK27g+QOCwfVnadp2AGSVnuRttvOD7CnWNUwuypqf+YPxeae2yNTlpv0tVTdmX
0V3Ip8tek6HWNOU0wb3msbjb/DunfvBTWEpbzAFReBfqUQCnBXtmzPdmvNfZrPh9lOoSpxFzvr9L
1epPFvnFmY2CQQI3vuIPPPLi3RNZwgfb0Dkp5MvLge/kc2zFa4YUR/nTBloh4VzPiBl2M5ckgnYM
JaNY5Yexd0A5b2ahoCPE4ilADPca//4nZdIauKlYnaVGDi59QA8S439/68++5+4Oy65cHOw4kfZP
MH+DKFpUXqbemvr57F6RCsXfWQXKcuB9SHD4Bj5N3mClm4xoDwjt9Ab79QI1xqggi87wZA+KJXdK
/CrgSaL+4FsapFieqEsy+7VUsT2zvzR/LDDpGQMF+a7efQ74wQiAlS1O0oxeb+HnD3/jc4r01YS2
mJR5+ZstVGEAghC8zy27dQUgsAxasLtV35bnZdtEfWrAPBxxOMIPPRRDlea9pAf42CsfBdWrIIcF
JWgyV9ZSCr+Rq6gRptRBAPc8tZmt3NgmYCY1Owz5Mp6dAd5HLcahhvc+VFGzm7eBACP2zuIKrAOJ
gL9Ya5oC430S3ea6qLvwbNtyyVi7f9fxjdWQETvZNkwr0evEu82Ep8kvWdOr/mUcLIOCOx20c6fP
KwdOIuQBZvTdcevZseI8IwcunBTaulIFXfJ86sI8+mfI6iLN6EgGhty/Lz18SAhwrTqjYqu+jGLY
sW0XV5RwdA1c4cXyS2Btz5nHb99xll+mSWWSv+8NyBcXMuF7P7ssoYVWb2NKIaeGjLgmVmAIAhNS
qOpej4S62KuK5Af1UoBSx6eyu4SYw/aGaIr+W9amoI3t5uPQy+aZp4ZPIePOYGa3Jjz0xpHbXuQj
Nww+fa4JM3bHbwq8GwPqa5ivLawbFLZsGPCbcMYk4Y+pdTcLva362U3I8te9Z3KxKLeAmMupXBbB
2X34Dnq/xzG9NJL7vBWMfgTYqs29Jhj7CIldAynlfPd3JLJuJf8FQYc47k1d3GHqr/sz4Q4nFUKd
yih6GX8muhH9TuvA0bxfUtEUxJJdPkO8uvoq3DSv+fMIEYZlBMEiklnZdSfsKfU2GtGgP4YRWA0W
7Vm/tZrCYD+jkkaQMhhX8eKZ/W62jI79FRZHZV5v1w8eU/YloAM0ezOJDjpC8YgWItwPst2FPVXj
zqLzFiwd42Ip1P58P3b2SnJI6kwIKyQqX4tZYtlrQpGRUQHc+oAD8wwd3FA8yW4YPes/lyGt3Ajs
0RO1yB1pmPDsxwqr8hS4o0nZfACh52GI0P/Sm9dLAgk7CiTCzSJ5mfS3mQA5ndGtk7e1vF2fEoWt
e18H31eIn6HGFAICw7IV/EUtniiK65Nz/HszeQFzRMZn+837uG23lpFc/MgE2o+ov1bnd0DS/nwl
GnfAg2UP37zIzZ2od7IrWS8KFyhhWG4IJbhGhbABOdHeNASKCjS0sDHG9MTAq2BNIJNyp+Tptf2A
zWGalNVjRh+kDE2t4wqg2rEtpMYJtCn6ai90vSbV2J126WfRRXhsOZBDKxxpRxEPawexs45dX/u4
l3LGf41T73jwfrEqPhKBUS7hDpzb8huzlssbQK7onuhYrKZG0G6CbHSzF+S1qINP1KmA5CICxGv9
b3dnxKnyJj4MaTu4YM6tGBUig/CDnj4VmBOlw/e+YrBdPlHLs0tT1lkNslhWQKtaehDdXRBobVSf
alxb7HdN/6t6AJs42vjI0FAnTv3i0+zAv/jK28l7qu8ij5lESAf/bsVijjqCeEF7vBW/3z1OyxSH
FgO0t4qfMZ7KuLvuKdqoPALvfc8oQOAjR28qo9b0u6ZthgUR+r/lUIFSBTG0sI7dCBh2WgzTIFGw
ElNT3OvGv1uF0Qt8Uzz2YVmjb0x8OpLf30Si2SFtNKi5JC2wku2nqRBnhVKzz7mE/Et1IX8JyuGh
8SNrimrS4VnHLNiYsayXSBlsl35naNdjvI5oyNkJO6b3mFXpj1VpPR3gHwZ5kXwMzj8pQhlkfU8w
bPDb45xqld+e+r/t2VUR+emO2DcgppPiurXLAEN3ZU3NLOo4TopqhpiajguTHfdTgQZCJPrDjy3A
d5tz0p490Eq37uuxmDKJVGrKv+aLWhPnbW5yOrZ5y+P4cuV7le+ao3F2HfFXQUKffFCNalM4D+AX
Y84f+obAM20zGchwtBTcy5GcmRuS1VrSKbQ/N341tl4CHXba2OJiPl4GNZnwWpIse04+0JtGRbg0
Bs/Tu2ApRIqTEgAgCOQJuHU/arjQWrL3Ae0D5kPpmv3ojYhay6fNyF644XitoLPss/JuScFch7jd
q1Lw0ZfqiRJNG0BGS9OihA1aY6t0nlsq/25TYG+uuyk/KPk3JKS3ordu8rtVbEDtnZam+jnf+5LC
MvbIEbT00IZYYI/CNAZYQYGxR/FVw3n+6dUdUf/2xFVKMrtMF3kaXESH96TqCscS7wPzY4Ae9DSs
7Y7r9Ra5VTUdtFRc1hl+x/ebmb6ZtpzhGKBPxtDh26YJG3e1xb8feP/SUAdIJkBzfewYVQcvMXIM
Z10Gr30C24Mw1mGMdx38Q58ZAkdZvSMm3VkGTCUz5G+yGh4LKzMZ93qwNaNI/qw+UCal5tz5GDLZ
EC0BgBnYDm5Y1gMdma0moBlK+t4ia9CxcYryMyj49DD7Hz6jU9C3trU1TVVxqV5OSxurNpJO2T7Q
9zDWqEQuQDyNFUfxS4txiFquaTD6BQjZK2Nm0ZP3llpwYwvr6ObHHjG05xHyfcnnIMBCYfDE7Lx5
43zzJTwS8kKQdKcwxtuIzJEmKosTXrswOVqV0WHvnTLtdNXC5Pg+qXIa5BPT57VjUBirAzbkb+pj
P68AxW0kx3DARPKN3z21DZMS5jc/9YjBysyJR05+zQnUzguIuwV7avDcmFuqjvlUABGmE3K7u+y4
NCXCaSgFsCjcS4UhTZjzwWwDOZS+k9IyNFjXwUzpF9xAloYMTRSJjIGh1txm1SHbCNRtwUg/MFw3
gQItns3dkqAp513yqi2E6JXZFftzEkHCxlWTvmn6/a/J+7W8jxzIJecBc+KzL8Te1CfnPr8SINB/
DF6FrAVVLLyGagKxbABgijRkVcvjEO3WcIwt3sl1GRslEBt7dsiaHwoFbb2mGQ3OyilnRLPRb/Ih
8TEbKS6EeMCeS7hR58gOWJW4Z/46HXlkS2t0thlz40e7mZyjV+c5BPSIFULmL0O+neK5WfzLtD6a
9//E3Tbixwu/QdsJRoiUYaUH3bmWtriNy9evIPG0rgUmy1/vPAgjUBJXjFJ5rgQeMLFq+ZoICgS1
pbMDLBg18Q6OT3ErJiS8/toB2n7Hz/am3mtPzBIKIVONpz1AoLGbr1Ju1R0vR2XKC1/8ijXDums/
lsXdCsLQsSrtTnOo+E/33M271dPBFJlaoTbEtChKUUDWpD4HfELmNjrE0Ir15PrsazerfnfK938P
JliGslJnG6koDRQQirYrv/RUXSkWGc3xXqVroKAlQgY4FW7c9EPDZDViGJcp6cfT5DXFInHk+TXB
QWPCYFZIORvA8bYSgCnlOYc5JzD/X+QhAD2qOI7Vpmdpy0xZzsDiFEWPhYtX8q6wMRoWiqqDDp7u
9AhbphU2HrUrVLMvkRI1JkM0UjrUIHDXvUo1rayEVtBQa024s7z+tCAUulaT0FjSLtmJVct+U4/n
dVNzAuyZfei9p2nsrLbPBDuukjGyzu8CqtyEPgxbWSHtyVjwMqWhIVDVPs7BGdl1txWnfHxe8+/R
pTOIs2L4Ra7k1RnpExClJ3EcyoFSV6mCHsdmkddABtFFioMoPJ7rC2kk9oY8Zeic8LjnYBs17jyP
9li6dnrola8cF5RLo5eyPANe1yLU+eQDCrmbhOddxBHn8/7jYmeVC5qEj9MCLeECKYoqVZLCz+K+
wq8DfMCgaCggJA0pAA3lg8rPbtqXyCaZPt2CYPo8J1R1esAWfrGqlRfsCa5X9Y0Pbc37h1pqlYxO
5IdUtkhXiUdDVMi0FtQPhO20Ko87Wf0kJEh28JrPLi+OefEv3ZfKjfXaoOvJ2qlDH6xZ+qK7VpVu
BYFy9qwU2vpgHp+w02A+SquN5Bg0Z5kdlUnabC+JghFpviM4VL1KYkrdUvNqPqprorJW60QWdfWw
j+0IIKF9jAgG2QeqDjiutQNqDtKm/ZVm4ukdpmeKTENd3Pfi/pjFgAwKAJ1pU2IuqxGHRE1/nTro
T9abtyeWs6g0xQKSlBO7EqmZH1RSsqibgKBP9m1ERgvSsOinalQtu6XGgwxVvqVG8O3syb4NhLVD
60O61TJ3g0+CpM0cfF5K3THznvI7nxGILBsSuRuqpWqEeLBX8+DN6xtj32zJY9Ug/Jf/AttPIPxs
ZVK2LsvQLwWfzIHuEsQIlmEBRW6WWHrIKiRkvWaWrpB9RirzvZD4MpSG5/uVw+zfYrr5hjqWbCdK
PPXPtOAdOL5hqRgJlV3z2h03QosWOFKdEGYCNzztfSlTJB1BjPRIymsBtgQkQwLeNpRrDI23tJmF
LO48bgXP1S9ZPa97DLeABRCuoed0M9WNJ4yvgM+PZLPc04Quz+AMQNSl0Ix/r/hVv9q0WqeB2fBr
Pj7FmiaURGsJCY50PlIjQRbhRsWXYbDNQNjM6NKxw0BfVkbsH0d9pAUBD40FeNBRtiOvU4aGXg8L
xyiiP1i79FgywJqJHKhM6RGaLm2nChqD7g5LNarAhjCkrpTI1Go9a4Yeam0JPdpSZ95YHRo2ldwf
cnDYeseYdWCzz2u967ZQud3+FzNGU57v+FIs9sW0TgNT2sGdWnyJzPZMz5pxyPCC/T+znPLZ1erK
9KCkmAjWbYugIqbparftM0l6uQjc6F5GeKRYaLvmkrSlWkPXx6lPav9SU0pLm+eGsolDBCiL7SZo
cdX05LAi0TYYVgqKCVuMo3KA+LP9efeIX03zHSHOElscAf31kq6/sJwtz+iESm6+lII3oMqolCXq
BDEPJ3EICWOOu+f2otJvy1+tZwx9MRWk7BZ4TjHMKy1Y+MF3Z/zTevijtak5rvs3mTUxH2Qn/FgG
Avav4Zpg3tLreHcP6WEZxGQxiYgsD+JKfACu5qNb5vve18WWcUKac02h2lE+9AM/VIucIFUok6S9
exhM5o6ygGMvnt/dFoZ/pgVlJ5RyH32ixh8gn9vVMt67Ek6ViYfZI++0KoTIyh5WAV8KujFXCOx+
SsyXvBmoeFfsbzRrJCLvoTRUEAqf5lQby0pBBf66r6tGV2JPIpZ7xMfEHHYYAeCh889ZaC7LigGB
ifHZdvBjZmrrXYUAiud0cmLlm3fJlVX9kD5+A/127uVJVhH2oxMB9M8P+zbG13v94j8ZZpXO57m+
PE5oLYt+ifI2C66salOECdSLk4kgIZdVLcl2TkIJPrwUnoqyiJRkzvWCWKAIuXQHbgPlqHHda3jy
21po+oG+GAndCGD+ne/HGnJ7QefMOJBDSMTWGN3Hm3ruPXG1sMc0e2Qtwii8AMRZ6zpBpd2FpVIH
zQ8msrdiHF2GYmqqu1km72PXbdVtBNMj7flpySYOtxyVBBCA20bUPsrgr/0/0AOrTl3eZcnGWrX0
REGlSdsOy+OiX4FbA93+vbuJCXB7Ou2tag+bj0/Xws438Of37fAAd1T6cg3DEcqaKZIZRO4DXjeq
pPPiU44NTuaQDOyvka1BW+pgiDXzqoWyjFS2C5mdZee1K2xPOckVJZidvE3PipsCeM5+/ZmVvIhB
ZA2nb9pZ9EbYvOnUCKOD02iE7/ewc5trz4RMVAXUTGNLYbAZR1qzmPVSELHqgHJH8GFRsYBiiEY/
PWlSBNmsZC4d7qdEpVvTeqB9NoJpjtpk5zdNzfZWfrotEgTbwkKpxwp48I0RSHJjIHCbROMIQIc/
PCPUqEke6kXSFa+gg1AcWV0XnjBHLNA38SCEa3LK/t6EYoM1ywZ6VFGj5gnZgIB3jivoQY4AlDlx
pTZNi2hsSHQ3aeBWnGKSZ3oX/vFeLqFwyXCLLKZsWG1QZ2K65Q94/TOm2+5FChJC1dTx4FjLVJDV
TFmfLnAkFOIf5+2XbfFQo1v+jyn5YXSBZbAq7gOfEQN214tPMQPhg/HZ7oT7c+VHySLtZmAMzcZG
Tt/nDVJL7+9/1aUIZSbVGd+lozQgGQHJFvxv6OEI0fpgjGayjXKTgySmEqGD7zYkgs2NduRSHkpd
/sp6tWS2Gj857L2X5x2Hl9oX2ShCUdLjbwEHW2Uw9GW92ZYi76Ju+JikanwD5ei59xSIUaTuhU5z
zMkFTAqdB8MKuQg/uikU0IfaUqO6ClhY0AkM0nQ2Vdrj+/2l0Pk7jQV27OOaeejYXekIQX90bPpH
WYlEMIHajheqFM2UcMcc/N+nVCLN4zxxd3kMTWd/my6yBxx10DjEy+QcBhq0iehbInqr312deYql
nrzYAWDQEFsL9BT2xjCltPpg/8tw58YYIkaDoqXJilIxjHc4xvEC0SeJJf9p75ihySEVG7RHrcRW
Xe6g/v5DLzGfv06BGHBH8YPhZfp/bf97Qq+jrznTMISGplY9z3S98JnxdExRzQOdaGa97oeaTBbR
NHxQe8WDR5LiFyqtEFndzfGW3sJXosp89z24JesYcljeVKvUTE9US5vfwThUNJHyFymxi2KIPVF/
89K1u255+RatlbCxQ55PHGDJngCZJOpiPz+at3b/CEIpHEO4ISgbaxfmMDaztc79urA6WfHYZ30u
xN6DLUEV7mdWE7rAnw576W79arGS8rgare8UEBkDy+Z8SU36IBMwkOMrSvd5RmJAyB5FNioA5jzw
RCHEwtDypPg1NWnLeH3NMHYznTOwIQp5KmMJssQjqJvIa14Wx/8f3IBzM+rC8fvup4DUMZx32T0E
WvqMn/dyhgj95C7rt/KHAjNxzgoGxyqo/UxpLzlP1pluy9/voCOIXED5/WqrAolBvcihfgOcbMXq
vWWwCLSb/+xWCU8p82qZyWiD0d4RVXE6i4N6+zQNE7f2pl5qYME6mKd7Nz147pCXgDdbySAHTshd
Al2CS7kcsfM+wGnpwZ4lwThmTRlO9uBjvcOlkljfcPDOqLRFCWy8NRjp5/TDGKg6E/pCVZR0Msua
m5hQmp/Kx4P+iaWkekkDpYuZzklmtPfUa6fZjQfsOk1QVM5wiciCKRuFTncQ62xnKj5ycMAg/z6I
nVSoYt7BZnjvuFVaO3lengnnyTZhQcdhl8+MeANgR4+abLAfO6esD9/5OCcv1WivXujr6fMnIuqS
fxeiwUc+e97fQySw+u+frzfPD34gJaAZjMB4ZkBXXY0niR6qIMR96DfQF4UvhauRbfhrdpp8wlMV
YUmaRAas+Eo6QHhgxPk2ubH491+of3qRQz1mk8SRCvTcafaxFT8xp6r0HFkNTxFS1yhSFOc9grpq
I3QDEkjDB9zoTq99GA/go8aUUQ4M7GwdAOZfCjj/7s5G93SVS3lqdGFJKFdr0PjaDfyLPeRtca7M
dJ56tOn7mDKlbs+MUU2DzRI1d3WxDTwaqCyPAeyfFMsv9JyU1Ajpm1ZQX1PUdgTp6gDGjeXMH1SV
cCf89OvyxukQSeULwf66e26c7o7IHfEAHZ6T9dN9hbqghQFzi018Xna/NLWDFO4YdbCgqIddgHNt
tX/SWI9cv8151IjPd32qRFUNS8To0vd2WyX6z5VP6qm3uR8XZJvoc4APxP71HReIuBaOQaJKaFsO
ISWdXY2QRicZEl8GIZ0ZXNbUQiKklaZ0UW8IVd0o0jhde3iXlWqmG+ZbokXaRjldRkwYVWBjJeAa
rwQz/Omk0JAiKm/tmF0EGfOkgbKYZH/jehu8/cZWc1icrRmemiJrfHnpTp8IBqWvYZh/PCkK6EFP
km4dZZLUwhaT8fr/aZejsX89XypTj8RkqXjbNK+fbNVKXl9pxcTohuV5dWNnWJWPGFpPMSXgK6Qn
lPWcHdxnxG8CL+Xlus6XevSsj788aVpIuiHFJlT6IrA/ZZ2OOAEqMq6qol0co4wE++y2ADJGW/Z8
KoqlvEA+6F0s7dwGXS/UU8hwBmnXVKO7lVNLmnDM4sg1pKXrzIr7hZK5wCG7dZWDwx3y7U03/scY
npeC6io433AbYQ+LIfviG2EO5ByHZvRyOVZL+KnULuwo7Q8xn7e2A4Hq/quzromiVSsjjdbEdmVP
OFqvMxRhrKCtyxuQbxJTD/32/lqfhpTmIPodEdF01dZelhgoC8NPpY0+RXGkFi9KRqFBGGmPXUQ0
H4MpOrA6F2BQKfKFOL9UlH+eQ+12y8puaJcwiFWqH4l7Pq/zNlt2EmzDxb3cwkarcw/tOvopVgXc
2GYiA/8b/vgRa1f2TbiYP1yDhJo/RjzUdR4Xm3SfHL/W1cQ0rvnt/Ben9JRgyRvMuzdcrd1loFzi
7yZQZc0vSUFC8Gfbur/AIw74+5jIKSiJnbuHH6Jws2JTzi3Q+Au6TsGXelpAKT1u09nW8/u1T3vs
8k9RD3T+RW6Oub/19gi/VsdKA/fErVS4yNPWyXKF3XOyRtxpg7cJMcGLQSyfeDywOsKtncq5zkn5
GJWMmyv3uUMViwqmAuMP7XtxuDzJNi5R9q5v9jV7IQw5gIyA5JWmgZDjxh9+sELM+h49CtneNgjY
GlV3+t5wcwDtFiB2L5Q+YXAeS7xNwnv+l9vc2oJRV1EkyDGJgFhr5Uy3s7RHZ4IRoveUJ5smrJG7
XuHacvDRIHZ4zpOy9zMHYb5E2/CNklT69412/b+vYcpQcWeKLL54XSk9cIbhNyhJJMTsskolVQ2h
IhERwmZg9fijbPWk/vZoSs3X2bVuwnexsmQ5uZalEDlJRioNzsCFa93EzURTC0QArGqijXtZHu2c
jhXT/u2ZOjOgFIrlnHGM1P8j+TJigKww33Otl7uilqm8DjjiRhX8QjPt0IWwnUTWXJKNwLF7CxgZ
hGPgTv7iGPZHcZW/aGGs6/A52TggAfymOJXaKSBrflXoEvHrFlusptWuj7UnaIHyPKjwrcIG0uXI
4CRrHxGX2ziNTXG4xzlIyC7E8FRDVGP1tEly+RVuOfZqoOJCWkQRdggbvicymmaPpzeIlp9w+fsZ
m4C7gk8NizBV1iHk2y3uEHHADUJexxAi3gK4ZPd0aH31DjOW0ZYFvmjEwKkdAyZhE+LDoLZ/ZN7Y
ft3i3sV4WEQ8u7zl7CvMlvcLXP5rKWVi4Rqfjikz8wmlDUGzxfUD/jUml4HRqDj6SVJZ9NaCoId9
CA151HdKr54g6ogYOARZp0LlRZCztTCPwcWi/n2KqgUbt7rkJ2Qv8rSYrXKRLUECFs1CLPW8o/KL
Jo8m/7+uHJMyzusq8LoiquZGxLTEN9wxj6j6Zx6I8uvSgFFX2+pV/oHrA9qSrcmhJZKm5W1motJ1
7Hi30qUIVHHNKvSIYQFNITyI2xewDWH4PKzdDXlEuvhtMu2NEioRI3wzhoADQ7tRzDWafVBRXP3q
Jgq1EbGcL7m/97ppvwuSFNb6qiHjpBzKrPTeSKTYH6iCdJU70nyChC9RwzfU+a2k0tjifZ0QvWvj
1wEv99+gBKVYTSXcIzVqb+Y8ATCbz6ZrWSJZIW4u171QsRhuhJGUQcFua5gbx6frYKU+EgoRAKSE
G1xZaldv1W/QuDyy/YrfY+MdIztJz7UIcJQL3cavfXLKOITWDsnoI8kIeIWspxuY9bEeQkCHpm8w
DFOiQljrhgOxcbKjDxj/GVy3AdiGtUH6Zoqzw4xx/PQ8zcEuRuaW73mKmNY0OVa9tfryuCT3ZKyr
nYZjHhpXEUJqOZOLLOIFFxU+14Ft1JuCEfZJwMXlNl4RJF4Q1rm2UJ8YTZxMdloPcca9TaRZS5Pu
Ou3tecRIF/+fymjRGvhC3VQth4K4JO11TY8xKVx1omV/dzIP2ccLXSjPgZXZtI3n4KlPv5ovwTgE
yxQnxnsSnwqkc39um+4gQV1W2A7FnH9suucxg5KpJZ0/BMLxSPBpWw9d5ClRvvqfbCHVAl02QL8y
vxiop2s/W4umGF5ndDsrUAe5PV9oxUfAcvXWd9fyoL75IArF5Urs/e50dh7T2yW2CbL6AYUnFM0e
GiqKuBvjP7EnC59Wt7mw6CaUKGTomiuOgJcxfOW4ADsxyQ5tv4o92wmPdPGz1oObfWsW2VlnN0XR
eAe/5eZEPJO4V8jm9qdjQvFzh+LVBF5Q9c90OCfozewACx9blhfyGCvIzMeYLX1C0F8Gw4BPZCRf
xgb6fvKpXJcHc6xjHzX6OHaoX2BfgbMsZ8Vsqmp0CyoNMmxlFBALEKXiyKP/FrUs1dYC8w+Vh2vI
aiwuul5eIE/iio/Aq0/JjNMV8ua57z6aS5XAVUr2rI/i6Ti7fPxky0WISWd4jsO7cmEvt+mWEVf4
iYHmgquJtgTQcXqXuBYDxJ0te8noUKXr5hFodIGSc/OXxVnmjpY93onnMeyI5+J9+GlQtertiH0+
SEQfmS3JwbsNgLLEtxLqWTEaP+sOWDCYdny3u34N1nxAzueSQRZd+RYAUOOnsY/yvq7R3hqeA1/k
MeRxnQtzprnCSZrx6FY14QfUhGQBFUB8sk1mEyLqkVdEg1jW7FtakhxBWQ0nzrIHO1p5lYFFbhtY
4fKAeFEA++U7WuziKGMFQcTUwMUUyXfNU6/uCsAsVBNRpQruUtVrgF0YzhclqTi0YJal854LvduF
Cdd7imYKujwfr3+d3JkB0EsqI5gDzsp+DCGb4Io85a6XNZ7VNChXyu3Gdtk9nqN+TQwrtFISzDqL
G1jkwRYrM/IpmER0HMcu1L6uiWUO0CVXaPII3GxaytalimNkM+r6lZ8v+4IPWa7J/fmbFV63/TML
C+vT8Yt2r7g0te7N8tgVVdc2+UH6856UQZaEFnKjeRWl2jfgPQyGFhk8GV1tAm+ac/pXtWBgSsAE
AFFCO1//V7NGrehSwGTqQcDlZ8+oi8jdmR+iX1YPxTT0nBjALWfcQ7Druk1slUtIgUBqzxzAEOPK
eq0b9AuGGAGL3J2PzrrmLM3WZB8X+FzJfoKoNtAaZ5tHY+qe3xEPxu1srhJdEJMgQZZC0LDae9Du
KvrX7om2V2OK7Q/9yy2Mc+6jAEACEhmVpV9JgBPhJiLku4ykSmN5KrOhU7P4aj/orNdkhWprVl9G
IrN+nmmHeQJtiGPSHswRrxFeaVtSQfB0kX/IrvZL+sMDQfQcJDEgz9uxPQfGUrPSwPpMHJrG4NPO
17ewcCyo2KHHnG/Klk7UcCW+nCrlCwLKmbAXfk2GxXltNsClRQG3idrtBb4xF4Dw+ulXgKmfOt5C
3CP+eZXa3NgtQRkNgcctvuDCSO4Y7raRmB0fKdE5SO7RZ4foMkPaei7L3+xvO8O7nrtMFV7+QqWv
PxG42M4xZRpY0A+FdNqylRyZe+J0Y0+RCnYcbVrwtmg624v+eHMzPV1zFOrnA6lYIDivQNVJSgYX
nJkaRHS2D96vSf54bEr0dxT6g7klHq3Mktv8XBzVpB23wR2k/hpXSsllRcLVWjiTVhEgpQQkEd+4
gbR/mnOuqT0W27bAEljAzNePiT4/7dICgsjn+Cge/TEDZcCdOQHw3ONfPLZFO1smvWF7PGkTty7P
xR2951r30KdPyG/nSvgsattB1BRXzbJp6moOS2jkNSACVp2h/KVGN0J4IJftdccfQ41ZxSColYPs
mz1vzIeEwKpIXSWiOoZMlI41h68oxkJm/X69x7o908y8p/NlwWtFGm4/im0w1kCoJwVJufnUoZau
csVj08w+sV4bAHdJcUFlAynVnVUPc9Z+9piBvOvapVrukYWOgDI8K7GQ6dqDIkXUvN+HCD0A5mnr
ole3rXLIuW6MoBjsh3cSk/huxXc+73LdKtiuGbZcwKjuh08+OO2m9NLZNOHfHdCVhyAK+0a6OfKg
IiD3ssK1Mc8o2mzTo00A/tNbA91uPgowgjWrJx5TCEdppiJ1lQhhLRHcqdjZ3hewxWyVGI5MD8lH
U6qmHeWenQDVOXcnQZchdxV1c9ogM2SFPeh+tU9RlVyK1rgFCLhFBuWROa5RareiCSFR7/zfnAmN
LRE1/ke7vw6n1peFzjogFxoOICSETu70j/jLSuAfGL2h2iVFGEBrzLca0DI+VwGCMNrnpHTsqBPp
bnywyOdXMdhg8w1mkginbYJx7WKLTfKCYJMfu6LiJuEcYUTI4cmdNJH/e1PEjJ7h43pFLkAKJvgM
gnSTQm/qTEkT5kvHCuM6aPNJcZ/zutUIpm5o96Oe6PsC7TOc2Kdzk9bJb+srs8O5oVEF/WBF+FgL
jl5VKRv3ak1Q+ilkhzHatzWRQ8vVrqS3nsKRItfF7eTSTYH8MJXNAoLwrlo5Me2ZTAWDFuhpxE5x
Y7+yQvwGNNPULtVuDQYn8ASBwHXhaDX74oeeEriFK9KeM7ulSfnyMiHTHrtjGNnq+GpbjzNrDAga
DSRjR3ifgaY+M7RRvG8FZbyt2VbC59m56SXgujsTkkyHxMRpBCgb6b84eUJ7Wa6HOEACMHMfxfPH
DBminoQVkeG4D8Bc99DIMmlSNW4Q6xW5pJRnnn97bjcvcrc1gGEKekqfHHegWw76u1k1ViXetbEY
cd5ldk3GstNV5wGzXRQH6FDHSmVudypChXG+j28ruYHRDKD+x238ZrePeYF7IdXkWYIsDPZSaTh8
N3h9z054vEdzQPycOE0vxzNqZDt1rCYztHwmlynuViBb/yq9lp+hY9vwrmgWjdaLmVhvXlYUoxY9
xG7VxQ5pGHYD+PuZtH5YkmLv6qQb3pJ3XG6WmUsiauoWYcVOUsb1K4chAYd/WhAezyu6q39eUkva
mhid83jaxz4JWpyfl5MDGcC9cZkuKe7LehC38Y009fTwiPSZZQLTgb4FUxARV16/TEZRp5i+Mx49
CT2kvqE84YrYeIAvxholit3P6bcgA1Fyfo+Nrnb4MVUIzqBZuHrUsNclZeHWB5dJD2b4ym6AmX2O
IhWXiAxb8XKTEi8mV+Xl+iZT5qMqPb6rHByC0L7uE1hoG+4FCownYlrFy0EUCZ3f02epPijFS/e9
JvaEygzUm8pgyM6nLrWtYuIEqA31Tr02ZRfrPpebx6L3IQs2ERUOh6tHRM8HKDDeXnAkwbpqLYQ4
UcEvtoEFwAZjcOse8TudzQTYvkj8TP8d7tYdFYk4+JQs3vq57CIwc0fUf80H1Fd8Un414Ws9vfSK
8w8cMvuFSbHbHehsOFFaoL3W0+lYhPA4jjhZF/5t1ltWXyd1k7hIH+0ddHnSPz0Ut54NOr1m49pI
OKTAAv/XW0K8zQFSwxhaF+Wlohh8fo6OajItv3X+txKNYc3A+V9Pm5e/SMGKoAtDf2HBXH8GwnBu
lRlF44ozUnob9eOt/87ux7bRTCkLKLPrw5XUXGok+z3tJr//b3O1uqTtEJx0PaNK4RhY/38HfiV2
YPity/SoW/V4D4ukxZW4Vd4DXmFS9fxnE7YOgFkBOnV0aBIn4GiUihm1BWgR39I2qucWp5Fp+ZW6
O/YNrlvegaDon7ooYRnVeZyCG4dX6qYFiCzwc174jugmDuiijx8u0NKtBmkDsY8sMFULx4dkKn5q
9iV8eW7wHqWuX3s3V7bQm9w1rlQr8VNhVFba0IC1C7Lh2d61pK5jQo6yflNrE+FNX0aWUL2gtdTn
co8RbY1j1z3kIa4APk1nbc6/Xa4PsKN+mVSjQJjAoKwDt7ywwdGAx5WvDhLPvLdNFq/+zv3Xg9+4
kW9kuPdU5BcgRlDKedO2shvM8EUGJsQ3c+9ozZSWqDq/GxTzJdCrVEm0SZMN57qhAD/Yv1mdUxvr
vFYn91Q1kjX7JHEuAljviY1rxN0UbFDubGgBe4Iy6ttcQpik3Bdf+IpTacD0aLYpOvfk3aTy0vUw
HzY+Kf37JbqvzJwK5VsSwWW9BKYMUmDQ1P4XGGLRQ4MVTQry+drCPAqsW1s2W/GvYB1GD3FsYhVG
TwNimbGPd8u79Jw7afR5l/P8iwoz0JTpmN7zV/HVrMW1oLhcQQMckqvSudJ5d1W2M3YO98sVB0Dl
oZsbyMQS98ssGpYkYqckTapeNPoztwSO5V/SZLl7ykWLw6NdBJ5nnU2QH6ipmtm1IQJQFchFDw1v
wM128JeyZsYRe2+edPm7F7x+p/yl1RgzK5RZ93Bq4xeeLpG5KhiH9FhUdWHD+nkEK4CWvm858c1R
KbLP/AzrD4X4FEUYgCYCIVqfPW2XByLYGn0nzRQlTIbwUm+02wWmR1ISYMSdIgLm3XHGMoP0EyJs
ZG6R/PyOs+2FWTuEhZTQpSzVT2c+ONQ4ocNsFjVYI7f6sKwgCxFhasa/cATnmHRR96GxuMssoisg
ThqJjQmYkhFKfrIDC+euMflwn58cKmMJnmXqwsgXuuEfTBrUdn462gBToCEzu4WZzPzJtRbMaM2O
YMf7xjsKZONEpKaU3utiG54srzhhrG6t9xfeO5Zt0BWZ+hBOs1oJ+ljL7bX/8m8jZZaLpQeLOwoC
KaV9dxz/DYIA2jlyOTAuvYlHGGBEVBoCU7xOEuMR9QcvHxk5c4JV7CTDksLbzh0yKW4426Mp2dvk
C+2PVNx4nEK0feB8808ue3lP0Dz/9ZM8qREwMeznFdtKVa+2u4u/qEBvlPgPtTloAGk16yqGXT2J
jQPsjDj7GNOnrTZWODDaupLznhJql2/mPmsLTPmsEwhgMJnK9xMUTyBU9qjxrNeIA84i7NiGSSI4
LU7HH8Lnsal4n8g0amvtc3B8KHu4JxQy5sn6jOBe/g7jVVhIvIFVjFsU8lOxI6vu8z8AyAQRJfcx
9gK9A2NchKgooT70j8A9FepqtffKusbWSbJiZGrDeewgbHyqsHANUnDIWBqNm9rbbo/2D7ZQSjx3
pYqhEaUcFba5f7g+wjQNoaS2YrIMuKYo1rWerJ7WhUoog7n31juMUeNSROjYLrtJD/CAfGIN1u2u
mgByTL5rJlijr8T9AvP1KcB+sUvZgqKTs0zsUUvBbppCebyz3zLXBFfKMPLN66aijw+zzQ8e6bJ1
gej3Z5gK9tieWc1sJSnQyglQeNW8wDUPoIcZNeiAOGqYypp1qEn/dpCBkDcZcujFBnERVXSijXEq
whaOHulrKt0dE4bdPtcnZeawmbX6WqXwLrjdDoQu4XAt435TPcdRH0Q0TRa5wHDNfnWLHdh79ii9
76IkB3xNHvkNEBRHzt7zcGIRrSe6m8JQE86g5kHs2x0yFjYvk8Rr67NM3jbVOgYVYVQu9Ai/cL/h
f7fycDtFWbxVgUJnZIgkNsUseg5vu87qeLbYMpR5Dka7i4jXj+2+5/JEdU45CVo1k1BGqBbID2y3
fdRIt4G8g7C8nZ23EBMjbI9QzwTkrF8glvHId6EKiVpN8Ugs51RglyjCWQzyhx29HD2vwyPlPa4O
Z3EkbxJnPftQkU+yBpabwZtzLjn0zhOmdxE0bCXCIkCTvdJhKp0LS7Ne50zxGzBGF9f6pZuYyS2/
hA4u7KeOfrCHB5O0H/YsBHpmpUgK6OOwCBwfcxGLefBhL171GRs0bSEwAogtzc0b/p6prKz0xIuV
a3M8QN57K9ekYGACKn6kuX1m2z8hG+VuCWtse26Ds0+YZ8kUS7L5eaFtDJcju6qFh1r+oXG3RxK1
tQMG0bBRIlaVQPXOy+CsCb0E2R8alFPbO0PtoC/a/6PohJ39tfQN/b4GBj3gNOCaJVgm+8aiDzPg
4LI1x8nG/5bIS3Ni5lQf0RyQpVtDfWJipESGeNubgl0G/QNxCchY9sh13JlBgJF2w3LpNKSuWSRa
O5wyf8F598yYuH0L2XEJkZXCM/I/AvrIXmMCFv0mRz3xobL6IdNZ+G1S2evseLUEqOeb/F4zoUGY
vO4dreu03ytgu29Ar1tjTIkq5cQTCr0Sr4YofeOvL0zHsXzPdJUNuF+CGFIg8UtZo+GoVmfH0EKm
cs9K2Pp4U9sbHp4TXdxsUZEEgQKy/BodwPUAQGcjO04f6tNfj7pa22PYpZ6oNzzHq7G4Z5u3PoXx
zbA6ZDH2ZgrG01/trnsGbl2RvB56kVoacaX4xNX1b4cth71Vgw26l9C+ytmGr/zsFSgJCUDvhQq6
xwyW6LMA3P5FTwaNT3lVC16BvQ/6sxjDy+19SBGyQfZHGka2beD29wqEGvHg15mXkgAU+q90F0JV
txixiWDj0FTiiCIoGbXAKhy/XjE2EKycDEnNShRY5WveZowQtYICjVUEdbChMiubCWolOOrofaeO
Pt6sxN6PqE1JfhsLtvCRgTprYp5KReBNqG8+A583nzUHS8Su2p/2Y88ShlGMDPcP4dC0ID5OnqRc
Xczp4YTLwwJmvzzm9UxBbm8GRcqVa7FJ+PZhvdEhaRyCR4jrc7mgzOov1M8jPCiOtHqWlO6YjDSN
COACN07P+VSmqviC9GB3TUOEUrEENDtMlQ5aIc71v1lcDwiFx93lNjNtfxqyZnY4QB2LAkL6c9Z3
iwO4PdYMW8mDzUPH15P7/dd4iYj/1zszBHTuKir29mRJOLDUC5gJ698xj3Jfs9kjxVl4qn3mFUJr
RMQXb1ZEGQFQ68c5afNA5FrCUGoWqtBEnyGK/xcNKQUPTlKGFRiIRz+WkEgmxBzB2RGX6byUGWxm
LAUNcEBed3dNf6BJifcPpmEAL+ujfNYCz1T2qvH01ysm5lFnzjRam7P0jh8kCwaDjDN3FAQ/dHKP
kQ5XhCDSrEHyfXi+Vj+g8u8z5zLA3yt0qGFucsdRJm7Z14lwtw/UGYxjrANO94Bja6Tn45Udof3j
Hvq8dRYzuOSor94ycU8AiqzENHOhas4UNsjKCKP7/aSu/lNxt4bW/U/RQfja/r78DFrKM2xSpaQs
WtfY6rTqbkcHC1of15O9N8gDzKANv2zep7/kRR9Ovmq1k05DpQ9p5k1KtGjXr+OxjNPoaIJOfTMW
ksYtMRRrWbKVbDpjcPNwazJQepURpM0/pRmMw6K66aDzcaGC94AG5v+krB90OJL15zWbbNaZivun
oKJ1YZLv+6tfVSRNnnBVWP2j7kXOXQdgReOpXuOE2K2BK9EVCN18LQZzU98o2Vca7oMiWd/firPm
iMbCSNabrHoTka6F1tnPXRDJnt7QrfPFZiWYaTjcNEbt2jo5HicSzhecQ8GBhrvR06LhvIgt2nLC
g1TMXzYUIATxl5rEmrLnzGY3RW2bK9CRCebYsPGM4+3wX8K/I1HHDGlhvVCTG9ISmY4jpbM9iblV
4GAni1E47u855nupNx364IHWMLwNXrmwVV1CTfUMwszbuALuQq2QYoC/dmb7kSrC1CrKQeHJSM1f
qHRIRP0SbBsEmR3kakANF5UG4Z9uTV4x6anwvCW3YAG7Fk0oDtpOOvgvaY0mmIcqMNAI4uPZNmfl
ETWO1DqlQ8g1meucJFmUYkf3I4k3jRV2Nk3UMI1qO3sS6fQ7LMt0HB6focZSda7sQhKcRGbk4sXu
BC2lHHW+jAQD3LfR1aF7OGqpMnAbZb/fHZvM0C7uU4ZvyHT/ftJIDB9kqzJH+MCtz1U5JQVXFtc6
QHtUccjchhv5BzjvS2KGaE2ob3lvx6O4bLqrVM7Xg191cBrXf4ND9q8ZdiGmQfvE7+qaSAqN/Jcn
aW2uvRSQYOFgEko8WmaEh7WEAMJD29l5wvW+LP+SnWZR4bRa6n5BPOUVYkoTWD7k5Akc+wAzVsKK
7NqqYfCZ498VtpNCDqprfSFQOwAic152LteSStUdIKhzI4httZMAA0JV8EefSA4G3+e7M7faADqw
XJe4jlcpOg4hF478wPBE4YPy+yrpFg1LCPLsZXHWQb7yDvjC1y0asH8TGHw59cQVZZ8Z1Ik7TWhf
RbAkHg/NuF5lWWZzXTN77xOL39+oK3Y8xRsBjHXvo7Y4LQUlsn+03mSn05tzzDTiToKGdPlVWYnf
yPodzDbVG1udzkD4Uht2YcBN8iWUZeCSNdlKzskzgQy6cbDhGwDxaG634GXiVJtJHQIeUXDv5EmN
MHKEdPvVziHqGlLd2D1F55lDINkOLirGfJJnov9CMOUcBRSu+6a15/9xVgSQxVoLD5zDjn2Ln9D/
lH0PuNk0Qkp5VQAMcG4X7wE9USw9I/46wh2GxqIPj3gLJ4NGNbBMf7c3NHtiJjFD0Bi8QwuKAdNg
x4Yv7i+CRHo1+rOxenadiEhUM4VQMzI0BHrHVMazC7ZZ8Y+rjvPkVMRE/T4dk6sj0fqzel8q3Xuc
t7gOzBrDZjfyiu1At59iuH4nl12S0L7or9IiHfejNxRGj6d4JcTd4gQKGO4yOXyu0NK/xfwhO3cg
5daxHxzTP2JykcwwqNoGf6dimUQuqMRldjzoAOYSaOOWTQgZb0toj9VZLxwdVQpelpfnLaoSH4fD
JEZ38v0AYI9nFlOwxMshpaThUDwlwM8YC2H0EsPKColUIO04QnsAXqY8ZWNr/2l26HOYag2vPDbt
Hu9P3bDZnjWBHfwOe5vIOguYyDcFqHC1T0SvTRgDEkW95ClbGBMSepiNcRZXxbzfSP3YRCJUjHOK
zYjUMKAp9Bx2Cw43KS4ltIFuhRqB0dKxVY+oIMP0o3ibwG9vGM13P0Gw/qhgh/zodkP9Z19OlEdf
fmJwhY6BCVXAzHpKIbbL4j16cXRUt3seEj3ISyU6SpscHiIYWF5SjarOhQdGo8jgChBzm0Unk4R9
UPFdC31G324wylMyCokTwrsu1tAXwVeoXCsXJVxF3v5Dx8Mx8UKQaE21h0mPg9ZdQ8Pxxf+6Es6L
8OZDerb19+C/A/P0XeXA0pUS8czGREG3KmIMn4qvAniNx4n7n3t+lYcCXDHDcDQG5xZWxQqi/4Ju
QYHErp7+R5BaGI3BcjWw4juZ6a5NhhxLb0a03vk8KUUUyIyfEXHnGK27oerNWFJZSaN4DZsdb7Ob
MqVHyDLS3HBWJCbUxZ8NL9gQbAbJxZw2bYjVOHHmtcAC8+IAXWGSlVQacC43VD7T7G00vYEkpIlP
mYvUIrSQdPsg2icIQog+tDdhg6X/ikK5uVNWvLrt1Ou8IT6o9skNvycT5jZGwfdZkWasJX6I2rkO
OG4b+mBqEDFGtEj+vZSXAG3xWRxGUtNvQGRI3b9rL2URDU/USr+BkJgKsYknCzGLJ7kPReWD1LSO
Jo16Vu/uw/HDxjFfVPBW0neykNe5Xm41XT4UpKzNGHdtzW54yYn1mClsXFWGavuzhFE05pzlzdp2
vfXJUYGRSkyLerZyoTkf+raNbg1b8j71G5er1r1OfDxJMZLjlVHV4teMT/H61VEnhPk50kaQ2pUN
4UNetViTNGzv4jYwYSpCmR0DzUVaqL9UrEJVDmbe7Mvw4wVozm4sej3mGbaFVIh+QVhAXW3q7xzr
v4PW4NZ9XWQj1Hhp6Y38OCa4xmHNjiHxWxRymB5xF/m9fzRq41Lf+7pBFEkSa/TBL+fwwtvR0ZgF
ccqfY3T0cuS8yRIu+cfuFZcGJg65czsJmVLT+Do27DX1Vmk8QfInBJXCpwHjunTYWzbWclyZORtf
G2xUDXlXwjT4duD2jLRx5IbMprlWNnRe1bkrj05icF0vfEF0QSA7qeZP5E2o+Z7Stb9X387Miluv
cHY8TOAlBgJTnotTTfVd1HhgTCVJiTHFPDR491r7LniDBX5BBl2Az4hfK3c8HKWEpiFuyMjEDh+r
I2gDqp8iJhOT2owYojbn/CA0LlzLgSpkwJFNE/TrUxfGDkQhx/w/6+6KlExisaes7u5Iq1W8iMYh
4dQMEFGm19AoXm7txg8jK7QKyV72c0Sjc0BjxQ+erWacffa0gDaauZtym0cK1A4Z1YplSSKxaA1Q
EApWrtPqLlTpquGnG6Bv92IW7QVV0ZW5qJtCbMan/76Y+f1jHHxHMbWqeS79J7ZKiqRpd1qSyk7H
bHAMZtKk5b1mFqSmKkUz2YPERry/GadF9/l61/wqow/Uq4ezugDU389JxKgPBlMPJa9YuqpTbWvE
eLJgRdAyEo0SvsSD87VSTCIh2vOeweL9DSg0pmkIujZxRTTz2yZYXbW0fkCJx03C3t4UsBy89um+
KdXMVZwjfqZHeBFijEsfOdrAI4xfJapEF3/pld8oUcZbiCvo//jwPHW8NJ5fyDWJWO6Kiu+MtA6V
BVr7RFbsgO1jALnOPXI2So5HTd8HrMEoUcH+8kvgl+IUMuKYKAwyjunj/Gt2lKUsCj92QmRwMHPz
30SyQeAKcU0XvOpgVd4XcHBj1Shb0AB0Hk7CxErXt0w4+Geh3/Lm0JFjM7dISBbgY6FB4AV8L72b
KiXlwR/Lv3ve5rFww9engVGl/2q0tNG2lgdao4dQtRfq5l/YNyLtBOpVGdco3co5cRZ3ePyTp0qL
g179XY8cQ2V4lUx1eGPlsKOsE4vIEICNOIVCEZJ46fKgtFJeml9W4Iz+zRAcEtamlrInAeNVYwxm
7ejlheGK1BWgH+TQNB0PRT8zTfT5ItvymGPoJcPbC2HAuydubwH3EDS6Yl4tRSs3q+dVnsfXjvcs
Y9i/VoTTJuxVLoBvSCwke6zfwCth2lSnJu2vnhZIqx7lDuC567ig51MY7GlK2b7VKoOta8HVSCJ/
7pZ34rPpGbO0eiQCAQBJhamvMZOU8sLccijhg0gv00E85qyA3cZppOlTBPTrD70Nvo2tbi5FR4fR
qnV8kXgUSKgE5u2K8rXML6ieyyez/+IBK+ohCZ4F5jnNusQxAVmM22ApIzHkfzEQkvT8ul08ZOkf
naZFWdJt9O7Ib1aD7Gc61qlZvyBvCnC1iQvwjPR3BhkUBZLvnYqX8ZLLeme5O1XzrsKRq7ch+yNW
cu6+RUVveN9G1UXlm8K5vB0jyrdWUU4d5dKDBDh/rHrGltebj69kWK14aaR2D5cHm2cG911wNoMu
nblVELPelJqYJnxnAZNz6Qmbiw9WhY6gM3+jMTDCPShbItUX+1dNFX/CJqT3Wy864wWA3G115Pu0
1xwggjSqLUe8phA0TUFW5DahmRAP+iJIo+agBS2cMBOtQGnWPETjt9vKCf7ya2fa6tbiyslpwJtt
zlYxJhD8jro8iyhpFqDrJvQ590KH9Ep8jxUq0/tNc0MXjB6SibyjpM32cgAcfnj1Iew7kXxD9pcS
u+5ORF7b2iIyeFxi9Daz10BYGCa/ev+S+/msVKWxOefiQww/eFPO54Ed5h6OewOc3jbAtpoMZtp2
K+Dugt2LtlR5zILeNpRcyTPhlOxGFTiQAQWgXQWUEWdF/t+za7jHqQUAjlIkxcCcQgOt8kS8O0Gm
Q5g2qRXHuH1WH31a03pxdvJGjx33WGMz9sriJ0ceOGgRW0f+MV74U8IbZOUGkIHegifxeNvviF5Q
9U/C02ID37CWtW6qQTnx5zjcL+uOQbr3+Y0OzTdgyxPEYQG/4v81REsD4DsoESAOr/AjLHIpHB5c
aOZFDvPtKjjYnFO0VgOnLyvhFatZIn6d3dUHTGDU+iYPpuXJae9z29JGZAp0XazJQF9mDEhGqIS8
cVp/zkIqIRM2weZ3LSKvjfUEpYohemxOkhmkoPu5BPcIpSAdeW+SyG28AWDyq086ij5Ic9Sj7kDr
8ol3S3a61Wvnusr5IPn8RI3d9KVcunj4/FthdXqQspJvTBGe/YMukEE9/ztQaXcFchXzMhUIEzFt
GlaIEun9gF09JdPhGk71VCQ/pIT64hpoclFgwLCRJTG7F+EIb+qqgTKf8kWXNMoWznoC1VudppFa
bbWtaVs2boixh5Cj2YNQ4Z9AQzJwZYsjKGUb+PB4hcY5SSP515vTfzG4hfYPDwFDPcrt//bxgYMk
nvx6s1T4IArk6VTZ21HfBvaxo+JxasAELXwqMTl5IAJ6c1jUXaRWNAVP8XwAtDSH5S+5lerfHswg
D0wUJTiXts1Atvj8O5UUSmRnIVsprTSWqSGPXf8ON1XgpUKvjI7mA3UIuDpROyvj2UNPWG8vfinO
+SzLqmm3w3CHCz1hrI0Es2WKGLiMb+XFCT3r5Q2NdhJjKKxVvKkq25En35vqncHRDATeUG6aSVMe
AeMdKA1VBnoIqm2fqlBf3zX/T87YudO0/ifeSRtEbqgv7bCWacFJ/8vDN9d5MiW/PlwloM4veS0+
2dPOtocaj3HzQaPs0ua2kyTKP2IDym/JZrdt572CuJErzxXmIjm2AysvMH906grvxWADoNeU81f6
lKeWh2bFgMkVP2cAf7JEUdAHZoSxmBBaDkq3rhETNdXCYfHC94Zijfa4rTe3OCIATu5rjgaJ2NkS
hThbdFWRjFDI/OVpk1rrr4ZqzuhNgZFRoWvyCvG5lp5paM7OloZebhFo3sPsGhL+pthWVB41OotP
Wbj4UKKTBrRqo/b+pVja4xOa8+LU7yFHgz5I4NFvzvxcEbQoMywWOUakmJ8coo3QzdxZsuHRzqiF
Fl803U4MmB+w8ULaUQ+3pOTyL7PkilquqUCJrhFZ1SfU1iu5ozbZjHWU0dF9H7fT4wRcL6McDPWL
SM/LqUqPo91JQmk6Gdqjj+xMlPbU6SaELoIGjiTIPOCmHrxwRgqwiGXWsntTTXuc+lhLN0Trgqdj
7DmLKFm11luF1pXWvXnPO6AL273rUTqyI4SM4KAVxcH6jdptmc4c2kXgSXow0BdmA8F8i9zjowEf
LNS0MwohBDEtNjG+ZTvl7nzLGI7HwA8Q+rR6b5PYrsyBitZCJjre1VMVAdlNI8ZfHyhKSqlTafRk
CuLbTYrNnYPaPP4JJi4L3bpgJX3gbb03q8/4csKounXUkA4cPviNIsLE3yj2tndsX5yd4LCL072R
aLrUkgShXxyGFf3NgzMh2U290G11weTLZQqHLU3/zT676R4tOUpWd3GnM7roc9qv4Doj/COuMsRy
jj92s6f2wngf7inVEsJAOBIX7YU9f2g3DXEe/eaNOBoPTpzVzeJ1g0vl680BQ1tD9imx5nBvND+G
YIP6mO382chdow7N6npIIKq5bTNsbc03ctqnDjfg2aMNnxFqwB/ne3WN6BjPI5wfPT3ALvkwXT5+
H4GI2POXb9tKzOhZNy8LwhpkRtSvOpUGuFklXHpgtZbP7tD8uXM1Wg4EpruDlRlUYGsJ9lkL9w0D
CBzz6EMTaJyXRgIEl0q5y6lKCI0zDtQhrf78dISBzMgZdLe3nxJXvpHsNw1in+TwDZin+gI0hjBD
wRtIw8+6MjRkbWZlLlFZD8OTymrFrZtgFdOH5Ml6hkJP1heB+ymUvLHotlKQwZUzD3y6p3w12a2+
YVj67UHQKZhXe6SznHuew4cwk3LiBQVfAFnVt/4JX4KCJ7BUBlN/RlokG6Lks5ygWyX+F9W2z7ga
x96QW2Iof5qbpScPcfY4xO/GljgIQhRSwgFuWFnawCxPTZ4eg5+emaCV6WvhTwbVpasBM9FzXHUO
OHV0cCtcnK8i9wbcI+fdfsLqqa0/0MXZoUYTySGhsD+tWLPdV74Eqiog0hOpCbnT61kbHXA6kQVp
1PaBQKFmS6Irj/67UTmN23mz2KP70MqUbc8FhcIhfcbB3bD0pQzo/hNAasvwhBukXVvf3hYv9I1F
k+X+km10ixZp49zwBMsAQTxH4+8YQ9oWjMjBAFXD55wZZ2+cXNTGWPkeS8SYikKmrevEvkfQBgU0
UVCIk7sHrXzJE8hWOyIotWgBMYspZe2DByilJWlSCI44vf84IMpCp3uhQOPcNFgE0Hof+N24/Mg1
nVNbDNZR4HcgIWPsNqATCnJqpHXhrsBLaLepex7rU2jrtazomssj1GZ/m+ulG70Fu4qh6FQZ7cjO
8lOniyHir+ICFF1TiDJg+X3z/slRH1k8//eomMspil9rD8Pb8AhgeMWmCKocv4EPI7BoJh34PR0/
dhizsLx+V2kBQBxsRamnXJT2ODrZdvQQGauHNUcjucpJUy4jN4Rv7KM9X73oF376o71Ai9a0fplS
aM1oTBDdJUtnFySwzq6WE4CJh207Cz4xd6sRVs0S3HgRYhh19u8uQGyuR0BwpQ1mEt+Qo6AuHbZ7
q+569ztQF5GOPtISYxQvhQxUt4VDnLZz90HwJyaO2TsrHizjYlqjZ9f9v7txuWA/L0KDhJOpiDBL
T5WwYkkh+5YJ07758ZecleH+EmF7wnbHNZpLGWB50D1uD3CvFDxxz5VYsVZx9OPQLKe7yhrc/faN
XP6zLeaWhIVdP13t2Y7Cakn/m2uH40+WAcnSe5gjwyo5OsgjJwD4Kerw8hyeg0zcW0hw4qeVA1xp
AUgNZrD2Fb8jRR1UkqYIV0GKf/umYlxwwbP9zQVwAx9RzrGTa5UDKV2IVRf7gMktbHDtdya7xqTb
kbioyTeSgukg4UVAWVTw2gg3bRiqf3b56rM6EkvAaSrSTUJTqKGTR9gT4MpsKFlfjIHmuXMN8Xso
sC7Z0mEbR1YDlPhVRLIpMxOPBoazCNCGrFFuFTt4XAKwQbCmVs3Awjqc6gmatoYelcboPY/dx+G6
+miEpmFJRjpml6hW0IGCUpVZxKPaNiVYuparYW47mQvU1loo7PNFzLv9YLDo0ar3AOm8fF14wf9t
52PG2er+iKq9hZAmM9dGQXd3j/lJlAnnn8bhnBqgszGvfl2lmN16yG+WXxVbGlwuqsVp+BJ1ShTr
mbMtcDtfQ8e84y2/5klhTo2zkNyTUnK5L1DPwEoJ9YVZDgycIc6gSc1MRh/2vmE4CkR9pZ4aQkPm
Qw3qYQocK/XyXaoyRXd87shgj/l+DeihTK3d1VXf1Zjr71L5xMF3wLb7WphWXiptv8fba6ffCPHp
Hry8qwmkgIOOJ+kJ4+lKq6HetvWGk5raJFnhMqoD1JGl8hs4iXX9baSaFM9Ko9IKNSfCz/JzFfC8
YjXmgpeTZB17YJiZeYGqvRmVvZtVQYLuWU1284LcNagQZmFEoWe3Hwe3f5fCjt0pV4ii5wLPW3Zw
tP3CIqZWY1BErAub4zGXL4oQCtx322jkeFlhObMvzXi6AhBYQJ0kRC7wDcvzXOG2T3ZNA84lSjTX
b6NuOHkXXUMZy59Cynzo9cqHidrx1GVZJDf9GNAGwSaBX95v8qUaZoLkRqVBVw2uuE1olUByQ/1B
KTA3ptKzUQFkB7RXnqVu0roAoy8FruJmHsuHr0L2mP2uZ46bw/ESnEdBMGGyOsqUH0ljqsOofZrp
lYtKq2D5tv4pnTcFmkhhE1MTiDDpfEJVC7C6XIpznE54UYTCj6IKIU3PQc/xY/eQshlU7rArKnoN
g3owiCQjQBclWGzdCi6/Hu1Cpw53oGxRZFInG89JH9hRoYhIufD6O29jbwHLUUrNuc/eqnW/jRQB
oSpGQS2tbBJQ8voCLWDc7TXXeVoaRPVmwg9L/rJ3XWGH8Z8dXkVk9fuh/sFNoJTWkIrLD/bzVJN7
2Caap8WvM+LSucHKCVkvvE9PHHlwRa1LxzVYkcriMNXjdonUhHL83Kny2wge92nXQIBaUmT2Puu0
bG1Kc3QMCJcscGCQET8nNXllBn3FP0ivLLKRvRIOOLoAzx+CXxg936uCaAwIDBP5ecRfLe+EU+3e
4TEYA6E99sboF9B1QmT8Oevs1ujugQbTr1fcOeRKNtHVXmKYPyaGUVwyJDaW++OmxXCRKQ2LRsn9
ZF/+8nciRqg2XdY+0Ms9Q3t8fr/ctycZKszQBtIT2ugWjYdDxHjZ87sKbYgqCN2nRzMIum1kRWHy
DKeWFYeFjuFENhREkKWqi/VSMfHaTS6yK+EmtTCXw+eaLFyLJEkopkoGZmMjzGcZlvALxCUaW1U2
Dk3ku+Q9ErACm7M5KpmKDAsEQ//OaZb/3YQ0Y8lNlV7lBYVY3gaITcn7Kmg51tq0IXtYNYt22Dn2
6cO3x/hCxhwTKdFG1648Ayij64DayrMhWKz06hb5QdDK7/pp2gKuv43KfMObPFIBvkul0msJcaOs
7FwX0Sdq1MCN0zyOTMF4LAIw0bWHT7zM8ZD9GolOEovxEtOJiSy1H9TGIS61I87ET1bvrkDaRGcq
mSGrW5NrUzdMe9HzvYRqLPBjvbVUWBI8jcPpb2ttUNfvwEPvFzQtghyHt3RRLBYQ1OgflS/lb6WJ
JB9UtMRZ/Ugm0eFsNKdPIWObVXtwQPx8CjtrnDRDw02lxyEUUOGIAyUf8luVBI5qudrZrTT/SwQk
yY/ov3OYBEmtn4+P0qhz9MKmm9SMX6SBquZFAsOFN9T2/A+Zw4J0U2kTQbyj0xZZ6Gpkmj0dEiDR
JmsOS68BmhZ8+y32ZLwMcQu7pkhIvo6AXFmTF5bWXQIZURWzGTBWO9Oq+FujVk2Xv+sqVZjk+EEU
KPHCkZ5Rg4J4DfxDFJ89aqQWQFdpWs1rSQW11ryi4/olohG+ljBiER/2heZlQVZx+4mxvAUanDHf
IKT9f1v6YLWLykecZQaKfhMJuIXulYi2EMDiCXJevTSSORx2EvZyyCWcUABV5lzoorHSmjMmKKDL
26K5lGZv7nxZdfsazZduiXKPsiUdfLhF0uENwMmk0ii9pRnjjUYd//hTokdZfzF/oxJkMbLRb0fu
jtrOSJNgkUtOKIqI7FHSZnfTGBw4Je2yCrwQGN5Tw8hUUvWj3mQrpySo6AwWKautgMwHuUDJJCiv
ZSYxTYBVnfwFuy9uW+2sFaJ86uelVoyO9L2ume5cmNmPjw2P5Gv2iFnNxQ2WbiLkF7ZUBechIV92
56ZENOww7sxs9BNwBPTqkDA+U9rGhUqdCp+dB+4iQ0nWOSbfrfnimlCWUlGmk0/qmbIvgO5Io0Xb
X4BaGnXfyaZ0GfphHnq3H5iYhA4zblD+w9bXB9OGOEKba67eKSNxPQEo1iHLTeH+t5OwjqWC3Fev
LXshus7u0KDmAQME5lAS/jEsXxwKmumn9I6hfoz4vI4b5bs+50UlUn0n6PV83461yiMsBrDBnBrs
8F8rcIlQjPcmQAeP/oW9bxixV6gDYXd2Lf4y+cjWk9ZQ5QqcSimSydZI06JCgaMTna07aMkfMeKg
I81yyLs0oDWsIeCvDK2u3Px5Q+K236unz1oTi9ghTuAuegmcUQrZQA67gx5gE1OhO9nrkZX6DlLM
J08ixfqQtc+Z/4K1kJ7Vgm5Q8TXDNEpSf+QRwGWEhO3ehikxMQU0Ds6nunjALXvsKNjAK3lRc2Tr
zIurg+BTXz2woET0P4MAJnZJXySJM/xIdUShI4wMKGJ9FOqbmZ3J8j0cPHveLaOJzU+JMsTV5mkM
UTjjHNKHCUYMninXtF+Ci9SpkaaUzJiQyqqtGGIPw8QGJO/uFxcRbhPDqMD8ThLWiuZi4WBIDv+Q
y9fHd0niprRJwMOYGa8j27eOY1kur+mP8IR8QhH3obEyqwW2BPgTLMeDhadIAPpAhkHhOPZcEkHF
YtQ0I/Oo+fNe85U4zzn7P0C/910Uf7UnSqO52KthqSpfyer7vF3I4vVe5NNbz2zfYRTczqjO2k2q
nnUCVIFyNIR+hRWxA9XlT1QrJWgQs2W6b5vaxCsA7WxhgIcfTEP29uv1F6CQFfXCrVIovdwnmVI/
FO+fHdUHwlYhXED1RWJ0ZXxn8zc1/YPdJsgfezCmxN4txVCqrs2wLb/WalvB+sXL+Y7N0QD/PeXH
hMExdv8R0tIxqsVHeJ6tJduMg/qhhBucivvYyGOO3cay0KmWpx8gfeIqOTw22vd4e9/kWykiVwfW
5H6S+VV8zTrA5UIsaohkcWFtTmSwUxBW1fTbRaDNtKNc1mLl/7MspswMSLsskjmvmLqQdMYYf5Ku
BSjv4qGZ5lrWwrXSZ3O1JLNogpm7FP7PXmcDpNGqrOd3XjXSoUhFyLEpTKnrhsGRnuY5C/74pKfA
6Z7YLVl1VYymzCwXqqwsznNdgilry6RyiftFWgeRelzndk/ad6y+1xRpc0UeX0hlUwH9Zx3OxuQo
CRevNoU9IgBp9c0MEGR0vBYwWODvSuk1L3GYMk39AJoecPr9rrno8rREGf6z5jW91puGcQhtAKY/
9iEiq8ViNXu2zccbxAiDyUB1iq9cY3nlqmPBwj3BbzIwfNS4JPO/W7FJuorK1yITjW1pa8tEUL/E
P/Pe26Y1igR9vCyKWkq3Bun3aY4nMsge/ieoI6cdD4ynWiVBCnWkSxRDI6pS9jbeFfP3/NuCISsn
T7h9jeXbFxz/rEqexoIkxDPDXaHQ0itsHPJR1KmTVTDA+MwbpcKVOsGg6un/dsuSMEAFVScwK+pP
NRi+5u2b8Yw84YlLGQXg4A7n4v4l43VIUGQpUU/tz3lO5ruPfrPqN0OV1isYHOduId3JHRmf2GTn
ZVbWhM4KWRRbQDOtX3tZTqN+IPjrOVVbt1QRa5t5imV2/zcoSzpf/MS4OSnbE8d8FXOjtWgEUHeq
HIglcpq19+we7UiQ3/xhIyZqFTHoQAx5J/WvBkJbGDF2CyiXxG8iKH47qAmz5t/BxfbAyy9NKXby
ivbu7fVm155sdZqId8RQaGQ5fomHgGpWnxCuvdkKgg2PQcar6Vpo2BErtlWKkmq3gS9xkXzqujut
mahkrq+8iwGsNZepS/tpGRla2npVkz1w1rKp8xrNhhdh0C+nt2NnU1vqYHcbbJ8gFGRfQ1nLT1pi
TPj9XlEkdRuIhIn40hi539hLg6zaRqC8sBCVb+Q69rfICfA+nAkD364mBJGWb4LQTxLAVUYLtoi9
F9j/YPHHXH3GUQLUaJx+Yq5kYgoq6uc+Xzn/Iv+y7xNXN92oqTOc5RTw0yiokigQvUqdrvb5EfKO
U958Dr9oTCqjm9KkhGxMLN+DCnNJO2tUSmHTntcep64InRcMtQOVHhKpiFhL3nTj3U1SXvbQt1If
H0Om/qSiuztQ4B8tpV5H5Je8Y2HRU7VUjRa/AfGPoM4o8EAEiUzz96Wgk1vqrryHLtHkuG9y2+6K
NkidYpqh04pNRbBv65V+wjtZX/I5wEPydUYAJxb4SAjkWw1MDwyuZu+FQvChoayqnXBN2ugJ7SoC
VXSH8MgazNHEFX991ciKktBZS/99Ehy84QPciDM7mNm6W8wRAntV2AbZXh134XhSlpfV0hKmFJz0
aaezgrDdtIUly9E5QpjiX28HQtfzXq1EWDcK/nJ+PbwoLtnODvE/jZrrr6T82w7chIYAEIK23IxT
BbCVrZnSceUvjPGwm+htW6UjxXFmvObO0kzcyvihJuR7F12jM7u7z8LHspnC1xWTSuU+cNC/H9Vr
boof5m2hgETkaF3Bo3o6XY9FhU1RM9HTz6QYC/ODX6bRLTPhtjvt9eX78VWsc3IStZnkTblsfKfU
wDHk+E464Pe9ypwhsizIzC6YFSSuVzxXyxafGR241E/zz3XU7w+A1syaswWlA4gAYPbtBCdcp27V
b80+A+kdsMW7jUU4ZZXqR/OewSF6PFqxXbN/Ts/nM7M9ko62UqPGYzROlaFgCJOdAXATf63Rb80K
AxL6FwwTfr8r3tpHRtQ8u7Gtbdppml66f4n0bGebXXQK3PlTPefJJmdvMX2xN/086p+WhkUXVNNH
mKI9Gsh8IyzKvQRQrbgm+3pOZaqRCnZsZ3R2Td2A1zEn0qEt3hNpC95a7a5KKYuKBBTFVtngfj66
k7JoF9aHZgMnVvW2biYzNsnNeKWvJVcXJDTiemwBKGjsge4YGhMrtB6JQMo2ot9zTfiYgdPkqJkS
hvwe2DtvpbOOluUOLMIKcOWfmI3nWrLyuNF6joAWER65G0Pa7pZha+8Nok47XQUWjYz56KmGH3SA
EVxuHXDbqvtigW9wFZwJOzZ/ou0/Ve76wEZ4CzDBQjr2lRWI+4R5jUCqS8vvXEQURo2FzaB1S3Jb
DjYgRturyJe3r4M8EBGmk+N1CLhXmnqktRi6eefQNQZUELOT0v2ZdF3ZPi09XO9KdZQebjvyb05r
fVsW5AvKOK2pHXf0RFXeZzPIyTbNmAPGVxqYE8qvlGNGl/W3QzRigedupeB/aBIiYfXxO9oEwn0L
d21B/y7VZmkx2gnDiGjFNQaoUaRzwNUDcK9PmdTU4FPa6Ycx3pfPK3NiHGTcRmyVgDn8IeP1aFow
/BnfMmOHhI4VSdvkKA7yqDqMgSSzlrYuMc+FAfsYfnWKKe5IT/k3slACffBhcEysqlJci8K1rceO
ZEEN/+A73jOOJ2AePsvB5P1xuFGA8ksFAsNVhR6xAM56issvRuWjOvox0iJLwTGvvWbZpO1RuhMB
8usTnScUdzUVitLdT+J2I1U3sHp/6uu2qsSBWMTzKCNikMK0th0ieJ+RO9hSCQE+SMyJtQJth9dR
J4RpgmUPnl1Yp9c9h76reW0qTgSU0KsUZMc2By8KwTBklNb2CVcNXEHdZBAx32/NwR3IlDVLUDQR
By2gdKcNlZ4Yph0zjrA+2ZjxA4j6bBZjiJjiVv3VZFLJ4GeObvJsz/i+mOQfAGt6sAdp3oQufiqC
9Xb01LFrOxvs0zHlvTOose9Am6qEr9dREk5wkIesImz2SQI8YsBL0FntQKvQ76nEXZPb6vwHBT75
6eBvruNxH2QFjrwNd4WGSuyiPSJ7YmzJU6NDX9nwT8LtraWtt+94u0o9SIY/k2TZu8yQEzvWRzKH
Zka/HUjNjm7oqAhaKuFya0LHCGJk5Q7YJ2rtGfIipo56/N5qQLZ2Ndf2OMyO8+jz4YNGnt0vmJr0
AzoTGHbyrtCKmEkmxHWR3jZZgndLxCD4yW+uXpf2k+Xq7pn4JL3H6zRxDKb+eFwkd9Vex8k6NrSm
DJfLMZC1TR3IRvpivTkFUpD4S51bfLIxknkOBFesAu/M4SBVmGH/AcT+tZYSdbZEKJlIxIVC8CPa
yf/O0FwqoZd7o1dr6/UH7zYUBXeBt/Z20xh8gMGp0TebE3Cm6N/GSsilNsp3TYfkE/a60IogLOLS
b+lWM2OH7wcv30zc6UJCRaY9BjmtRhxQupccFGiwbAGtVJXq0/BY8o8KKKthErfCy0hoOx8LDD3P
49n3SkjIhjkVdsBtlKQraly8XbRIJG06c/SVOQalRVAxsFf6o730yJ2vglId9kTSyq2dZtDs5bB5
axq/Hx4X63IHv6nRrK2D32142CDl1P0tUEBHLbFsedp6nCSHzvPEhYKibGR68xYLKbAZQ15t1CR9
0zbhsr6FpeglW/Z8gqhzMtR8Ce2jg1UTX6IPWWr3pd5nT0PqKChE4B8as2Rs/KXGqqgTDs5jbpvn
r6HBYo5SHuFE1zQLej5S4NWM9TQNqAE0ZwYsFOI+1S9+OUsAsunr75cHlJpx6wCXBXCXEK0JFM1L
QlsR8WS6brVD4SiPBhUR8E3pKwY/Sb9ICcZjX/+6pwfAHBpwoCGF/SdeVx4ie5vjoElM434P7u7P
5BAH9UIHXPDDZ/oQrjbNHNV9jBo9bU4ZXEXpUtLIv+WtG3nosrlUQbT1zRPKnFTS2kzN2KtFYrxm
eE0dJxpyPJodz1elcTY0FNwdVK6cmlvN3JjlEBVkfOkQ2zKR2U1AL7hgAv3eV3UyLk4Svivg+gIE
sPOJe1p3cHcuGAMzSVoUy4+efCAX3/yyFSO3ygdMekSxsSV1I5vnDfM65xQqIJpnluyzKslkJfCq
DTGjOXI2JPCDqjw1oAycQQeBmfSC/jtUR3N4Qz9pzRKwdqPBFXi6zRUR+BZViUK0ieamKaQ+iPaM
PV/42XjcJASIESZxAtd3owFBGc3L7cHE8YhOAaPKKRxmScSivB8eostsEFM9c1e836twBlPo1Qxd
hgWbcumqBB2HUYBuzX+wzA3VAvs531FWd1Ajyx//imtNljQU41fBdyDA80qUSw8UTLveWcEDneYW
oEFP73+2ykMvAOhJZxsqm7kytxG65/sQHRfglD4jhUgvl/rhfNGMA1xOfhsVkjYIRAcoNyxxoI3T
bg9H6IEqocFmGG03s7ayJlH1rn0u2bTXa9thkuz1MAyf7uJnqcgjQgxVKGR+PvxWTJaOS0iumi3X
pHxzzx5MsioJ42/lSQRxgRfC6FQKqXgEa2MqE4c4EMCtNTmWhlyzaP18wWs4mulRdbV1yQfZFB5T
0Gf2iXwSieN2/GvM8LQIqPFDLuHbyRnXCMYgiFd63Gp1AmUhcyw0BXJJJWgiZ9aN9gWIEviZ7/dV
iVxOJ8ztdthlYlQZQ3VzRRY1NbEZLjWIDUpnxEm8PreI8A4qZz5KzOIUfEYw4FGTzYfy1xiwGgpF
WHG4RRnrIwjMDELGK4hNiCJ7JpcSjovX7tFzkxC3OnkspI0VLsPdpqhXYdpZb/uTDGimjUlX0bGv
l9+y8fmBRKPumqVDI5J6MCQRL5/yl4a0yGz7/c2zFy9TMMnzlt76q8pRv5uhfFzAjnTTXvvR84nU
7IRCV/Nx41dkquifdoKDnBApCGbIeOrdjCRiDDhWK0bRUcKc9gwXiCqLnh0KHsPfvZVLr0aTt2tG
f/ml9G/kSsyok9srdWugVZbjTz8Mt+kCCa1BVMwsZjLmxMViLFzSb4T9nfDwWLxm16ZWmCaxNvi/
WzGg3dYCAC58gZSQMFiHI95S4h3Qjr2thSI6x3SqSMzcfDcmnjx7G+v/BSB/q8Ydeyv2ODPZD8if
GdR/Fylr2QQg6aSVLoeT3S26bUm6++0/z3I9t13TWHHSr1ArdlnUaVxRbf1mu5TzPiBTH5VGJAs8
vjvm6g3Ip06O8RR1NYXEZ2wS/+0NgNWHn8x/OqNoHT8Dgw3m/eoqAjMy8w7/NP602yblUKCTqat0
0EwjxLYfu8NAklPn3GZ4MF/uuncxOSGvu0lBwUku2K9EASTFbsF/Z8ge46JChYyhZAAX3pTW8GvZ
E++wyVF2Jx7Ag66mUQZzgtrQNNxXZD1LQsXXjrmZKeU839SVKQ57hSqrfEK+kVLgcxwUqGebvrze
2Snz+YA7OHjtngcxBQZKsQWuNV3C81XPQATzTfYx6mEzsdibe0C/Zb52+P04aKx8M9HW/AFs8u6u
2zCN4TPcbiRZGHbfg9LAmdrqY1u5I0n9iWhg7qarzqRgeLI6FNurClO8Wo3Y7HwrZ6X4l64ZS8Vi
cc+y6myhAsOND4vWPDQJl37BdweaernYb26X6caovT3Ig5ppcR5aiUN1PYtAGZL/EG1Mwg5KXDSN
6tq3UnI4K//PD7m5AKL/nghue5nQYj8bkQ97vnmt8dtrabvRZ3+ohzAZ3QJewY640U+R1407C5hR
mJIC2CBELJlT97Jhehpu1p1Ai+XfjHlPWiQiiNsAoY86HEpJU6I5fDHD2cBB31OdLfPEbwBnCDQF
Wcb15cJDetXd/ivxzvpxOLeZV4Ev/ySOsCRs6ZqT0EU8VOFXfHIgBQq4F2+y1gaUWMm8gA4nsLYk
2voVqZrKfP9MndwSBD05SXz/XrkZWd9B7NI62EaXApbTrORZtdNDir0fzFqv8ArDHcayqqkTQ/G2
9q6e7/kQXx5crbRmMXGhDImqrViwXeJE5Ogcdc3ybd6ixymI1Q2PTkNd2UlmOPJI1eJ178qQr/z5
K+OMDr9SqU7XUKIrSnRd5bKQ5cjs9nUOEB0BRbR1pr0R1DVrmtGJggXxUzkXxewn9CIhATV+yRLF
oggybeoSK5qUngwYagm/XXBpRKJpUeAmPTVbc998EvQssWm4sQOHK9+aeZVo0hOTwOX911fBtbnM
AKyfL2xi7cpLSdwsrrizg2GYXs+bHFyRfVaunfGnwYrVS9wcyhR134vBJqzigNrnzZCPpkk4tgOd
y5btFVQ47KqzdPiNRNbNGm0Xw+P315TyVbaM2JlHjJkI0bUG3/WF1GHmTv1ZpLkuEr+jvogeLSWy
hWGFNkuaDsQPiJ7ds6JTS+wmqTvU++ICtuEb9nVYeWr61LCGFiKs2PmSXepGWx9T3RGorLpFdvBO
xzZS41s02CYQplczFsmHOhKCbCHidE9IG1fTGAd2F71GFJPW/XdggWEyNfi8C70CJuCpREigBj7r
1V8Pgw3CHLVKUyBlm8aoYSHOZJmOxFscxdkvVLkcrq3+juSO0pJUgEOT1MGS/tzTEyYoe+eI384N
gAaoZGF/aMt02Kp6pM52+6SyyuZG5MiOCD1vsE1+x24LPm73xdSIL2byBcLjvB0QHRwQp1aRvqUz
h1kDhDjeV6iEFVdUwB7UOR7PIoa48QUnLaR58bKo1AVbz0wS+VjoHJP8mkP0OmOq2zkWUUmrWMfC
2mw2DSgbn7Dzz91dWQI5lUaAS1vrBgc61Vmyu//eeNogBlBL9aXmTiY2+vqN9sAwoIDAjxhpv01x
cMi9CHqWISfwejbF29207vLj0tU/C7FkbhWtqpgqeoaTqpo8sIqfHjzA7c4jr3zLd+TspCqrJCKa
LFr7QXlH1+djoUjiQw9GSMJ0UE0zSyvjBrqwX/FnhO1WFOVrXdseeqxCZVLTE8u5vajBHtQYLowN
MxTEHkcDy1vOqDF+jhrN1YfJw8iCvDbtLsy5A6twFEwI1XydO3MalPTiRYOCQjWeN21pw52+7Jim
TYkoJVFV8yv2CRjcnTbOOO3gZwT2lGjrfMmiPCRNM6iyH8wpfxu9c5diQC/WKdO6kKo/6aMWKRVy
XGtVk8B35cWFXUB+agfHPJI8B4Q5kLPaeEYYEFa8ZRAiGVNxHbjCjC26TcO00g86wYre9DbPFlXW
VUGHhhohW4RBe4fvK+I+h2/wzpbzSuHM+3X1qMx8GXUA1a0jgzlY6G3YGt6dYnT57cV/Y91fJ9pB
ry7GoIQ/ooVw4Mr0GxSosNzxT+TrA5uTYeyFecSVpnTxVJJ3462dI13twNdOns+7PfFKsUBwdVFW
0wfb/nRsAU2++sW1sIaKBP3w3vVRah+ag+s7ED+6YyMavmPV7jE1BANTPr0aa5kbvH+4g8mxLngg
+j0XPeU7HhtSIgnN9PsHCDnviEl9BtKk3olMhDKoTrPipaS5DI1Aw36wKNwyddlOPUcM0CuZ3R4r
h8v7Zg24FYf2a7g4FmEmfFoy+g2PzvswoNRxxV4tIFq+6/FaSNyymkXBNr5IC6q3ssZTIDv9BtTA
//tyyGHLCYCu5vgXQ/gwxX1EPqslrhkgJz6Ygrv4nOlMDbU52otLgzaG4YJwVks+33JxLvXP5ecp
TTKIAlnfpKQSqS1yVy0JTAvD2pmpiyq2nxCSGv11cEp7fawYJecMyvWNsWFopJNLOeMpLWkVjltS
3HkquTUQ3FV2hFpyfBycnVo6KRH0fdaSfl0zatA1HwSNDIF0urojvLHT+mXQRreL/ZUt+lwjZ4os
BCIw9//pvJCLRruaJQdc0zT2HIuJgfu9F58Ocoex8AqUrtYBs3w9AHcSoae0Cjkbobpa0XdHV8ap
DyFfndxQtGWc1jFcNvMMAaeX+D1/4QFM/M6KnCdoGQ/191Gq+ZdakxRWVy+SOvoZ3MA4Teo4xEZR
m1rj8+G6kf2dlO8l7K3osCn7yXSOTj9DOQD7olBl1kIJJ7XRWWUEm4JKcd99//xfNFlX+SiLwg5U
vCjHaqraahsVw8phYeSrkq31cR1++RTbEF2HQkFocqVpV0Qox+mZ4EMPcxLKHNBu6MqaT7J9D0/Z
UH3X3Uxk/DGaZ9MSkuoFgrSYI3msq+vK2HDIhtM7x/vO0Y9FN4EFhuxkCCaELtnlJ/9U/61vizHQ
dDg5xTVo/SqiRSc6/xbvFT4ywiQPkZnVhyz6FV4HexqtpoelvrkJwSoIdupg4r8tqOtkIzvzv3LQ
7vsMpWAfLA6FJPw7S30YjPgtiXqlhmsiaOwpwMBe5YWali0uf5leCNytjkcvaGQpvwoXKqgsx56g
Bpn7EoShS3JM9k3Yg9n8FQZHswhhJdy2GWkr7Mf4hv9dNgUygHUqCcHEagRMcn3nu/0faokwDvUg
JmTvYDoakE0LTHh9PM3vK0ywIZtICrATFeW0qoJQH7ShFJS1ZgfO9kAu//vHtH6AB+m9fXqmJFhS
D7HQlXSkw1ab2ieDW4HAY9BRg1bGeAORlEz2IcfBc24IsF6Bm/IJsW8LQ2A/d8bdS6v5k5JFibS8
86DGoTaZ2HUWE/mk3nOIllXcTVRqXUUezeh9CPDFSnev4gNOONSgkhMa8Sgm/xhbpCBnERa2RhKI
fNqAvlazeFPmp3yKQTuVJf3vhPSc3RJUKHqLHOIg4jj7w6spXUaythE7OfJgHMjtNmSawnyVO5KC
BCMl2pYJWQm+pp0VptU8gsAGNwAH19QBaQgCe8Zt6RgJaykUfnKa+Sfm0LMJmVfK3CS9C5PhT9xC
GLiuFIBz2QX5ROpfN0XipDgnZ8kEGnLfopx7cp4qLtdFZhLMmyZC/WB5N1rqdIL1zmDLEOYOvZRU
IhVd5EPZv4VePA7HfQbghQPJmC87g1i31ruJfDIaDIY7wnjKV22C+pwZ4CFCarwwfQiTV/KQ2oLE
VogzdkbnumO8TLTdjqEbfUSbmiFx5oVJPzeq08zjKF5+ZL24UeAl2xnw31vsKYZ25tKFkUzz9gDw
Q41kXX/OpVnLrtVgbCqG5vruyJLe9zdu9MKGiCy4TCe62cdFesMQbttWy5vE4rbc0jXg8WW+BE0+
eFmSmAOcUlaPgBgRfK7Vu44ff+tlcPkc74QC8VOHOJKXpShcOEfjpR/nPO0tJjkbvxNJLaJRIFgN
NA9lBwIgmnbCYzWY+AmbhuhnrHGUkZf9q0J01Vp1VnWX/DnxgK8gP7heASH0+Y6YcBaGk+pCJ2IY
DSCRL2kK+sjAzNe9+ITaMuYY5UiZU9RhIbIQR2zDvDjd4AIlGOGWh0dDBLeVnU3NuYE8DtbIvNNj
kbm5xgOohO/V4OjsUI/OKl0StghdO2BFLXPhObj6SjEBor97D/jIwDj1qnOBNSm/wzAOvuYXfIdv
9foF/cNNVKvZY1L/p+9vizZYte8boYkbYEjMLLzQEiHvkUiggFOWQrsgugLT1Na3Im1xK1iuF0Re
bq311zus1/x8QMyXIqAvuzLmGuFpAnCo+VOuH6513t2nvV0kUEWOjXKx2BGJjp7pOWC1ZOeAFX+8
+6ta5Z6cRjqTXDdrO6FEOuZWqhMLbkOMhH+Dme8RzacPUWC8ec+hHNwqiGnsN78EdPLD0E5o9fKp
RqQxkQReO3a89C1ijtMNzWhQTbEM56h0hnjhSN4CxzZcWV3tEZEXNiaKZDMweiDKQA/qXDV0rRKK
3+I72qhBBFGkvmTC/Qcx7+mPO6NJtOON33YW9FHv+oaeXIpYAnYReCDEu4M3NJ33nfPkr3VDi3RP
a5bQne5N/QzDm2pmQOapl5UCt0YuvuQw7NmS6utA+Gfu1TZ8Si7ivueqXriF47i2VbQTWxf7RhEu
BM7gjW/dsPzg9N4cXkLtI9NbVnW01SiS79daF4lb3M0nfSpY2vtGYY34jOMzqqIDeMhfZu8pXo0h
IRpf05DVCxtTGQ2epEk+ki4Tkg5jZ0HeOwWuVa+H2itJZMqeteVvmuKsW5iu6C3kIOgEri7SCl5h
s0GI53IOjZ5QBoKU6O0abHWshi1YTo+8dk631XYY71jfZjz41SxhrLHzaiEfrA6dKKkqNYCp9AjD
pMWQdaNnU/UiGDJGa3T0FrxiAfXid0n4motcihc/1ZuP6/yPu4tvo8Vzi9Q640iJJHuk1PHI+akt
nQ+0wpphtcJYAKSHM3UEsd0BcyzJM6kDxS9/EgomESZxZCvEZfEct+fBSAJEYaXPhFHYRO5b++Af
dx1O2AMMlkLfeZtvGp+dzEkYrYpOVo1vilSgWEy1jTA2v2sVGsFMFMNGOh3H3wUedEMz1OWGEMIp
Gkw30N61wvWPaomcQhR4FyRZGY/PfVQcfIpytXchQ05SNELbYVnJJ6sJDGP76Q0dzs0FchMK2gZ/
3lchY/wKMYR772qex8sACZfuJHiKLBILY+zyo8BnmgaGGrz1aK62rEKuAc0DfQi36QVTD84V285G
wAFs3WyxJ3dJZel57YmIho3HRItOdBiTyjvAokYfhyUeM3por4G35VRls8K517Qsbnh98tW5desz
FUjldOsGxFpVE58f5/EjI7YJDdFUAgT95yiWUJp5XUO7YdEp00XwdfmAWeLUw2bIy73emVkv+P/7
bCb6GfMXqCzVgN2G2GJKNfSvGW827BQci9FYGFNP3GB4XpiKacgrDzfxUiID1eDplkAhjN3KuTNn
rjgI1wDjmJcBn2f52wQZqKw6INwBfsIFZYvCWqP7av89KhDvSTu1T06acgnCMd8c28INhTIlmvL2
MIRmDIzaou1NHnFaBsvFks3WQ5OW/QnS73ksZuTsILo4a+V4d0f5cdC6E5IUbTOOUXAp3AKGlfYR
JZ+8V3t8v5VSTN9yixiA2y/8j8/Lhj1A/7/riKPCBKorQ5L892xJCwx8aReC+hxXKDvsi+1hJtk3
/g/p3hi1qAj4mBAkGnxybh4ERCGv8PW+ffwEmIhgURZGCHGhsMhmGXwGP924uwrBlrruDLLisc+t
4o7IOiM6D793XcK++p8gVtO4tLpsyF6W0TWT/bcg5NsNFGeshXMEQjDmC9GdS1AoZT2Kzo8s8Jj6
2MN2gM1tVtzyMguuE7eww3n/DJuiAe5yZjYAK36nn+qpu2UmPEGHbhmjCT2PC+VNRYaqrKPZQequ
ITdr27IMzhxYi0qk1JUiS/dXujSK9eePhECLAXG8mJyqHWtkTAMmDkAJM+UYAM/WG/rXzmc2ISC/
UGYE720LLj0gG4w2KxI58mXYb+qUG8bLin0I5JbiZtIf6kggnrB0zoe6a4Ww0L2HA8Pi73ne11Cv
o3RAWjFv1KIUS/Ya+F/7Xs08jlR9GkPbT6L1f5p56VSCVC2ZAC4Ot1kXdQQ/LLoMipx8TfyoL/tf
YpS8yY7vM5zeyCbwMpt19fKdzB5N9YqnwaHKDDDc9d2W/NvxSkhLnLHcTdtcv6VPiS31s2538tIh
XlbeHlcL1pqZZcAis+dvr/d65Zgne7vwx17s4bGnvf57JQ7P4HpXMjtA7ez21d84+dNrGQ7sCdci
uQ3ShCiFSJgvMigoQ+neGlvmiiBjrKVEuuN26+dN12xXahXKWyjJkECHbzJAyjAJKYe+1jwRu7G/
fmz0kj3Gqtw29ucSnnmCwhBeunwVzLQuEurNbDgfMRLmzs58Evv3JFqGudeWvlWTN55QUHG1tID6
0t5WC/0Uyg4EVBsaGEOZK97sn6VRlMhy1KOn6ADXnqHYLiaPl026+Fmol/X8MmlPVAymj+t1O9G7
V4u9d/x2Ksl3odz2T+Py9fYwK4soAG3DpSwCb5AR2VhAa077gavixKr9/eaZUgGL4J20Jfkh53Er
vlQ4MlLkwP/vIQR1eXv3aRbxBWC1akTPl7Vvf/Xx+2k6RUwKtUm2O9TK8K9vrkqf0RDG/Ac0Omev
uV/70OdyMhxLUOJVwXxTS4ZZnWmzUvz3K02WW4vMNX1Di8W1VZmq28ZfAVHZsDLYSzf4FrBehT7h
1Pkdm42Dr2ze+t2RshSOVhnA0Id1uz0o8wuj+LVc5f0jR/A7lKuKOf+4lyZqBiemS7AFAproDEqL
xCASpE+wMd2rIxR85UMElHgCv7q/X87VuxavT39YltfqHv4VeU7tTO4cgJXoNoqE3+eyLHu6g3d7
g6QQ9EPosnF/nflmd6HIUDtYS5IJM9RSh/wseNnqlreAX2gd27FKHSA6JantYo7ZIRTeRfVEimee
cKpGIDC4IYZnV/YOGZFwb8TnjRX6R4Wp12YBjlmiZjxtrNaHOnnCW3FGjBx+d/HD9+0sjoysXKeI
71b4OnDFVnJyB0O0ttlzORp4UnhYkHmclcWggSvHrnMwLW1nV9toafOy1BUuaNuTOztCDwXOcjuS
2HQeUd0z0Cq29bJJbCTbb7yYfnatmo/gHXftGD+2jBa551ItxN0mlrNjSMCRfy8fIVBq992oVy1W
UZddLz2AgtLw/ytLQlA3N25N9yQvHzi6m2CtniEU9r0MVlsSVn89ARfmEYUaRrvqTxmSaxvNI0WV
EPzNhGxExamLsQMI2hKoYlbc8Wk9a9wKXDY1h51YAKyjbBY+aM8ZNXrVojhAgJ4FILm2f1mC6bLN
DnaI4gRZoYkUu4orOA38wOaoPD1gCMWXlRzU82xa6SS+G6QvNwubsgAOV2vQbTAVTdtU9fCL5hNI
Hl5oRGXz7ZjzYK2luSD0SwCTNG73GGNQ0tSezP/cA4kLZlonG79ydPqrK3/rRYJAWSaOTbZYL3uk
rVceVqdzamibEhl4rJDmTe7I29qjrEd7UO20r7zNwPc40I5zPVFHFROGhbVAjHoE1b4qyXr91bCn
qRdh1XO3FlMNVDVQiFKJMvm7xq9I4v4dzy6uWarXoFYBlG2S45DnTFr+3Hfiw162MUOYe4qaxl8v
uzUAJC59kJZBQvXvNK7Apy64xuEXL6Ntkj6wugvF3MdzclMPEtOTvHEMGxZ2NsLqcqK1m8y9Pv2v
i5+IjmYsNtFxzTTAUth0ArmgmyrXY+1t6OHOsa8+pMDwwptFHYoPmUjBk/O9nHjTO6mSArsPqMnu
z9nRklL49uNyEIRPq6odnXEcUIXGJU20y9d69N2ROcCb/sCCFfVTj9x299jDCHQBLOC7yXn5Ufe3
hvlYmWKAJxyy/m1PBI2jWz9sddvz35UFxSvB1igbKx3J30h4L8yJRWFTLbbViwd6CQOvbg5D/zQo
Hp6ynVNpSROJX2aG3xgb7xv8he0Bk1IJF5cWB4jr9QBmSJ3if1VNSRGM+JdKcoQ6ynRIv5dcbhPy
2ES7wwPj5DcUiNmM/pL/egF8Kv3npGXoN/ogNFKSUI2d4+LH/bWzfGe48BtWuXiq9ZsCe2rlmXMB
Q9UxQK0nwaslBUPHntunKrjJIL/OlASjQTA2e63YuK9QCe4Tt7Q8szIlw2RnnVJF3VUFYxr41dQq
smjOe7UxjRwbUEccbQNMj3aqnp8ynmqiy/QHKsOte0z3cjExgGJNGSzezb3YA9/NCNCaS4MsRzK8
vChTKmMjjSO/iIF5vF1TRtxa/pa+i8Kd33XHQ82Z67cErA1I7c6OT1M8fPzYf4AX4AFxk28+AaJW
jHLvj/IRYXrC6f/r80h9xOoOiKy2fSEhus7qsXGQl7yWQ29DwLkULkROFSenK/WftgYLoxKTrcFS
Kv4pWAEQCBt4omlmuKf2dTUkgvQ+eJsghPeIuFwTQuvc06Z9Zw7GRMBM0oU/v1brb4J3mzUBD+Ga
PB9+JVE5HSg2Dd5kHlupQGuP1t/ETCG3n8NrZlU++koIOddyZknY0MG5jZ9BJTepDmofvthWrS5H
tTZZ2pWlDeUzuQEHCK0ivzvGpZlEbmJ0hKlDs+npc9DjBpY71QKr6ziqzEMRbmJ1X/t6QPabs+P4
u2GniaxSzRnlfFgLiwJiQRcC+KPmlWcBx3DThsSbASRfn4p6Pmano2FRc4TKjuCYzyF4srHAWgzt
IyvBw9DUqqhL+B80Wrirh0ioQ2pAN+VNXg2xdBx7ZjFJqoTV8dDeRBV5HXPnzUZV06Jj57Hr0YUV
UKcpySVU8uqbldqvUEb86M7LKbaboSI/uB4cIWOO2ALnoaj+eybbQsraiZi9H9NQ5Xozts89yupj
K7WCrfTkSSa7E0sBxyDVUwtENC8h+0zs+CsJpvxKySAJ9FFbMqwTDoJ2Wyl8YCUkceKrHCIK+zyM
7UkLxh6qJ1W8T15kCDSAmEMcjl11my80VdHSv7UTbOfb1Jy3MYg2G8I/XiF+7HejCUBe1l99xZdx
Q/7kwXwZzqGQGGVNmH/vcelQBuCdo5RoK1qCia8a3/8UGsLD5XFza4SslqOT/SD6gMw1rdM8PIGo
m2FRGeuaDJqC8uNhfg/5pOMRB6BHSIsA0WggBmH1OuurGdvGLWBwb2y0z+uQWHD3uqwqb2hr3MWP
8UouampoT1kVzCm9fD+k2t08DsSt1uajnqQPgy5IySTWrOEgBD8AAtKDc7qaXK0I8QLrHK1nea3Y
xo0mQaOj7AJKg+TXHT7I8JjCasg+rtWViMM80YecJzu52MRv7cqaNL6stcVS4fQNV7cKRX7bQY8U
m04iut/R0R5AKbKnqWcfcS9PAllpiv9b7YctNrtwks5DdBkoEd8cZ15tRWns/nISgdc0CNx1DP34
vw+WTA1h7I7pvW6SOQHmxH9v7ifaV6zjiF81c9I0DwKx8bk5ZHXF3cER+q33+Vpg81DxE73KBH8C
DSCeSnYJ2WPgq048kcdZiigyfAupMGWJfWKAmHK46gFtJNZxKf8XJtaktLGER3TPpORW9s+TczKm
AK2gR3FxhgxphxslDSgWa36JYcWfIo3MbmwS8mQUNQDnwzy8fJ8/DwXfbik5PDnS3D9EBDn/e9io
N7zxJOtohi4N99sPurxp6b7uRb1ZybRg2pj8cr0xuMhms4buUQop1llwiAycRbWvlbdJFbjgaENi
BY+0ODbMoVELsvAbBbh283tBY6U6Xg8lpQ58FJOoRAi+xqbOvfFgcqNQR4NsbbINqWwY1z1V+iin
iRK4NL6Me3icbBD2yxB92o8Y/6wZNRkUCg/4QJdBSCI8pQZje519PsUuMYN/JgKmW7gH4gNUcz/k
ZwsWTQEBBHq7LOimBZG22+jchqfmAPMDjwLRyUnGlhZ4A5gbTGxKd5OCP/q7biTOoH75upemTqbf
HCAxrZC5lXwd1YNQAlQg84wsDjLrCqXGLsJHHfC0YJdN7WZ2ePkIIvgKMFtmc69hzmugU9H3BPhF
yJTp2RA3VQQK7qxyWYOSX20nUpQL/J9fUfRgh/pmkkH8PS4a1YpqV0i1TkcE0T0EWuz9zME2McOM
umlQ8MFDv05d9h8lx79fSGl+JXcfm12UYhPd09eg91fJZSL4f08ZuP6k76eYkHDsZr/Y0Uy71MJr
gVSmLKKRm2alHIOE/o/vf+u8EWpuO0KacllThDi/QHxZNPjeIIdNZGmsht8w8TjvvLdZC7MA14dA
HqydNWtfmqzWZp6Xr3myLEp+1cnVgZQd4LYRqwf86r4hrNA8/suzOvj8kK4uMWL2/WGxOPHsRzFQ
XO1bkdHq6A7BzTXWr54IGoGJmnByvAJnMkacq05I9ahQVWLdIm3wIZtrZTgi6t8lDRgpyEO9ucJl
wtKTPXnsYS74RHuF9JoNQ0fATK15XH7ePE017XjswxXnBZA/BxzrvcGyPQ+EjysRJg6OpKZJlOFv
/Drh6/3sHaexa/6S/C/5HLN+d+Roa+TOcoCUaxT0HaTe/5h8qtLoF9DV3X/6oQmZBdPCJVqURmDT
fP/q4hLcoX6u3EgYjmMeGVBEP0HpOsbipTqNubnYIxuS/Ed/uPY7kOQFT6CYDFeRnxVs5UIPWTwQ
ECuXHd7ouSwQGCfdYgJI5OOyr70tq//HfFftpSI+3RWqI2ssILNA1C2pOE6iysctyGhDlCPKUgPt
QaYi7dvKgCcgHajHZmpicdsrlhDphd81f5mviinB/mcP88on4cfEIWD4OS6bDCF3XQ07lL7llHX1
csjkekMd7OygU6s9SmWUt6JS5SPyLowQr4PVxFjh2+PCcmtTel8SZvP4WVsOAEEo9BebmJdsD4hG
VXH5Ewe1ZAtZ3ySudlqBfuEZz9iWC++OjaJnaVxHn6zsb+C3/psiWmd8Gycou9wIhMAmtGYhSxqd
BkCBnJTS0oG0SozKFO9/CAin+4OvqPuZXXWLHBUMIRgkmkp8uZDR1VneEyn5SGuYxMLoplHcGxNZ
GWZqYqk01IH+Hf9cclFSqnlLJn1A5EMw099nFh1V60r7YKw8CZ+0d4Iw98mq7oZOEqgMNNRh270g
8L4uHwqssHoHt/dKcrcL39/o0kxwB4qYaOzA0JC8R4ZpIeho7H7zWWn8BbwE++jTNvGb0EOncSGJ
wihZ+YSlPWeArmU82w4v8YyeQgwvI5a+e1baJjZibf8IYPAaO3BTQDmO+hcPfnMh8PljDevtOvlM
XlYmM1Sb6iKyL5QNUc1a1Ps0WYart8MNYrkQ8zLAuA2nYnsiWzrWIKbhJQFBVa0W4+B2pAnv0kyq
MDhoy1+fV3MsTNRk3SM536bPU8v3ZAUDHnr3o8/UY2xggoetK7GBINzw9VPrfEBSLvhd29SOxu4v
oMvNZIT4cqol8vumTQcRibDGoT2A7qAtSDp3xndpCa1rxhZr3VJuYdUbo0L7JRkNCfArSagT0Eaz
U500Qz42Qr6gD4o9KRMTdiIdoxa3hi74YtnKiG/YxCJttP3PE6fsZcTVyrsJv3EooO2Dkq/VaVyI
j86bAQzIW3soCNoxnZO189QcLXV5qjUGXqD1LhPCKUPoFCmFH8KvFFVtmM8khEfAKYBtlSdORBWo
uY0zq1SqL255yIc6wRXlf4hZxmxS0LwuF6bvp5qpPAktlC1yiqIwIE6tZl9ZCG2LDgVihEheErR+
2Wr2qeLqZcL7teyagKSqicpoFr6ggLkMzqVVcQveRzm+gqzebJ8+NT2s9pynU74EQAMx3kWanUuk
6vSkvl1MFitIhOhhtmqTKUW/3BAcLslIGyetHBNQe6VMPP8AlJ0x9QbqcCJ1dH6+yvgXFT9GafHI
Opetr/S3EQp2Uj7RZvd5otgFmZkmnN1r/69k4T8FzZ5A6BQfVwuq38ig3VHFnNyMqcFk0ZXgMYJR
dsEYTmIFj2Ky5XPJ9OLQDwveyEhmYOgcKGmj1Kxfl/RQKneyXhSs15g8Z3lgvF5d2PS4qe5w5+I5
jejejV5yhSPw7OHggOSiR82S7kA3F84p331YTk2x32s5prfC0x5NYOab1C8oK7f2aoefb7w83odw
DnG6l3mZ/TAxplTosD1TlPSdpy//IO637TLW/vKQsfDb5t77szndIcCNJ8C7MpF957p6yS6HfDfZ
31tjZVGaIJMyUuGhaoVkr5nKgBcw2cbI1RN8TZYikmpvrFVm9QhZlNpLshIi2V805NnM2L/uc7JA
k8h9++owoUZ4Kwkz1FniW2CiUq5ykYvwtkPvGNQEcJDs/q2wtOu5lvAX95NFVuLLydo3LQkxYvBE
za7IgCzvm05fmkQfbqlDEYabV0Sx43cULrG6bbxKNKygGLMS5z1o2NijsYIP5laagoUvyiz6B2QK
woYTaSzB5sTIwoADq3nJMFtt8qbo5FfftQZGg4kBCWrqFpvbzM6z+J4OxJSoF75zQrYbm2E4Mha/
dhthFjW8z87j6rVop8vqvLZrrm0losa8cDUBtMxJPlOghVcgRWrogFWjtunz1I0BKPTdfNZSamQu
MMxruPBK36fQG2E/rR9QhzTOm/svUAf7i21UC/Mq4U8AJT9IdJ88NiEYZIGOI41sXMPUY1MwNYLc
xWhhzWB2UQEHoKSJ6FjEQvjhLn9QKF1a5FeNjpOT1lKnsR7RILIBvSKeilCZlB4UG4WoyMAPBnUW
bbtTrw7DJdfyPr2nDyPDRuZ239sHymwyfDHBsKBI9UV1M3zIH+l8+NAw6F5ybGrZlbvgPdH2TlYV
SLcPo5IZPNpbBKitfqD88VVKTn8oqChk8eMY/tohfr9TFz4vuMP0KSrzxmsAo07BUTlLvbB5I5M8
me4NCKAjQ7BBc7veR7ya9j1KXYONt/rXyc6KMjmBsVblJNCeKXVkMH6VnogAk4vrMy7v5Qkt6Sjs
tWQ1A1kDdKHxkuqS/xoYu0GUXQ4+jO4VQUDC67sdTIdAEdaLvv0QK2HweAF5753Dga6xAGXkBOx1
LGfKTGmu3AyGvY4sJCMjQW6KUQMOPom9hfrS44/3BiyBI8wqXtJtFYrtIUYQqGrXIAgWGYqEXdgS
Wcw8UlEtxCe41WYqlAXZyw1oG986TFweRBVwxY+FE2u4aY4zQYcv722OSoGvyMXcU4xnPpXZ0cLN
Yw1/pnHTbdTKGi5Ys6g1wU7WmOcoqaS7Yxtfvp0jtwrwCSrljNQHdjk4XHt1pe8/QB2zaCurcvev
R+7JKu/5d3sDyxr58MfRwHJig8dBEdIznvKBofNZ3Qkb1tuZ5wE/bOzIt2S+seUqgB0LYCwHx7NH
KqcGGfipNEpxxK4pGJ6HMc3BNJNHt+NxqXM+OxjHoHDCQ8aHIXHCrS3yXNWtr3DAzks7VKbvy8k1
Om9Tg8hvgcHvSnzR6Cjgsek+kKEeuxIydzqPzNuBBm0Ta2rwHPgSSfCiLcU3GcM0w0u2G2ssPgeu
KAHGfAKYU5RfiK6PXlV2YHglBDQKYvwTLuKmxMCMU3Q/9gkv/+ogLQaHamJG8xhV4hIL9+KaEO4c
x6yU5DlloNTa9aRXFOrLG7BfVuQLvVsCjbvC8YA+Wu0TOXV1zrL+RnkXGBqmBoaXLqoArEm8sIQS
w63BhKob3fxxu2nIBWX8vmo2ihSBIBVusZ864QYk9nsjZ7v/rJBMZcG8nMktmaz/T9PuOl6vjus+
3G4Mr54ku8H5dluvQuCFhR+Ip/4I1uTIIGzY9Vt3hZ6D4RCfRJLtLNQyaE7WKb0nPEOzmqJqh5mq
YPeuGEbMW9H5SrweGSnzDsaENIwOsfCjGD19FeiFI5hkFJYuVNCovZI/2suqOT4EIiuVmfxTE1W9
cmkdBULhfEf1SKePGmdCJ8o5FPDOrQoGLeFPpva2Wd6Qe784ysnaLPZpQPjY2wi7SNCi7EgikdhN
GE042ucRFG5NeWiHwiJK3yXSbKoAjeof98XHbF5JV+2zTI9FZCp5MFI/uuCZGbGsNLgz8wKz1OV4
mYGcp89uwt1hunmIOOjFIyIVx/XiAPVTZn48etuRirEP5Y+reOC9zPmmNviucyTHrxZAxX+i6sEn
2DfrN6sOjFzcObWfNP6clxL1eKpTGQ7gL7AI2I3L7SG15g1vfPgeR3NaxHOu9uv1hZO03ZlXbxyh
8F3/vBDwms/9J3dujnpMuvtEtARB0KH0tG3uXdxhlGPiCIGTjUMn2uyHL+B/EJGSvMvs7BidA+gb
JMsBCw8s4fV5wcEn+qXetVAGlqeYMY5CyCDBTu5g/SnR2T1rLaKgBLbcRO818p9YvHo0ONN0Rx4t
AcMDepu1jDsoMBs0IkqX+Oj8jBYd54cX6nDz2O25IiquYkroZsYbm6lyUQ6hQwz5Al38D5tF1CgB
9t3DhmIqlxXPU48H9hOfY0NzGAI/Py6oqx03hiXYz4QZG2DmRi36AizKoOkhqI6CMVKPYbHo9UVl
swOij3lOWxL7sknZ6IEOhoieiiiPbHoM4RBmuIfjxLY2AjIe2uG+WgLGUUTyiTevkGt7D3VjNhY8
06e58i2b6kWz1DATO140KAzxC0wrJ5xPGLulbxK/WrFjYZTpr7iHul5591IzmVj2J+hYscsPSoMQ
WBNjzKH/+T0tBPHg1yBNzkOKzgMNzGODN4Hs2kkvPY5CsDneryjKSgzNCN+l+CM6Q8FLOlkfv5qX
3Kp8ojuqBqKGYpsOJ248t9pjHKe60wL4oLp/tnWG/P9n7A9VeFG2gZSdNSMLkAd4Gx4pE3x27pCj
hhO6l0fZJhW2rnRrXUrIvZuEqAeBSQIcJ6QiGD76RIaBmhU/RY3pUn1Iev6RbQtXN0sWhqzpYv3D
fwLxpLhlQpi27lhM8S37JEnxlzUx2A64bUMA4MCafOYazPjBIOyXr6yNZ2peppC3cCJY4zenD0Hb
oC9QE0s3wUNdBJ+LemKbigPRpoEx27MVmUpo6Z7WDmeH40huoTmyUSqPRY9dWSIjKOpXLy7oaZ8R
PdhcfctbUxrYxjUvictmWtx5Qxj2n6lHrNxzY52zXHw/ZbqU1Vyfz0tTJ7tDYwztzkOofgtXCM6x
I0i8+L0RoCUCGk2sqQZ5PR4wc9884XwJz23FxDYWkZkVjFNxOlZsnUZ8OWP7E+ZhwWljlFeBSrqh
d7Kvi+2hnnJlOiNyC6m6h8ip3MGplkLelhna+x3TFXcMC44aU0oh5cmp8W2Dw1wLjuPfe+FdqMNm
P7KlGP2M9/3hDbJqRf8XdMpoCBM3HFKqcl/HSW1U/VF8qj6HNyiA2bG4yBwQKJhv6OovzlmZ+HTN
PNVtMVPLMlBVtWB1Rt9oVcutl1H8sp+MCCdUruuiAZJIwTfIqwyrBdcGnDc1IATtSy6AJWxyHjhI
VUI1D4YrBHEKzairvSkid2sVcKA3FmzPaPJjXQMnO9zTvI9VWyNK9LgJInr6+WDIlaMYtE2flnWB
632cwn3uyeRd32jcA+i34F1e6XXqbV7lrm3+nZgs0ixHR952sAuCMkGEW8T5p5jqtMkpkj1+l0IW
9ELk20ESxJeUnA8Lpu7UuhjHJHDL4B3w7rWNsbs69NXHl6fwOplQHvSJ4y9lxXf4mZK+oSknIxJW
R4g2uYGOonQX+HGjbbO+Eus6mPY31tOSRi8JaYVyJpvqLeRCJpV3TrHr6NMEuZ2vzeZMfP7Vpoul
O+4PHbL4fc6g98by/9plPr3A+AVtGKVMvtBvgZKPaavlxz8jP9lQHTdJYIsuzrAuoJB/32QbtC+R
GbA/EoqBGpnMcu/4CxIHE6wRh7IeMoYrBjg7YJKlKt4EJrVBLqjTpvfjt0yoZ13x5KLtURIUBAWw
KnSOGpXDjSjMwGKkAEPskEzK4l7qkxerM0OyosgkWl96zPwyDncNKSveu7MJCoJ5yZhbGDSZNdzc
+ST9mBLpyi0t7vc4pcrpFGq32/gKXDIq6MXTYieUZnRwrqAexK5JzKQFxIs+RY2qmjnOZb27H7tD
AwoTebowmOIAlTJ5oKEaF9Ueb6Q7/4Z3ffTxidr9RKu58XRWsHUSioWHwQIjQPvXA+ZMrZEpzbGa
7TQv+NkMSYGORPmIOQha4QB/O8VWMEbRwcAEbjRYI08DPbnJgKy/t/luGWf7kvHf7uOP9foaPN7s
I/VCE4p/XJr/RcF4VIcfIxP2HPW5TL/O0QzfWnxQLqN1tF6P8wIKN3DBwws9NT88Pj5Hn157jbio
iy7lnfsbxdqO9Nn2zNXPOwKSG5GHRzFfcTKHp3oAVZ59u9PH8yncJpZ5f9byTxrj8w+yq/asrmqZ
vqn3l23lZ0IgYyr4WiSkJM/WzpGkBzbR7eB4hWNlOaEZN82iwdwg3kc+9ZA4mvxGQzWofVpJk9EL
jLsIqm8+YjQAImnkzTr1Z9p+wde5UA++axYd+XQ2Pn1q6LUJNCWoN7XdItU+y+9BJ6Z+RDLIIhGe
X9LJ0FKGCgzKjfhvGm1sbrlP8jYYpG/LOZu0L904nJ6HXfBJt9Irg13s3GRBSVx/9IAHWVzj4gr+
TByp584Os69jA150wDRJ9n3vLlnw2SEBN3ka0l73RhYu5IEVDxtTyyUnQtBVnEeo7gDbXzfmJVQp
TwXOXpu4B2AMIFhugpau5sXPrPT2ce4YNWlKFuJ+TTdowjlzPszVDOnqPzorBvc2oEhh2lqPMjI8
VnQivMRPvaRu9evZU+IyAtFlg8vjzxIYF7Dx/kJZL2vG8htKg+7R6LHLvB4FJO8Bqs5FJ9mrQLCU
IPGxUVzGhwdPXQfGKS4LKJyOO3QV4GvC1oEsx/zvTg5OAgS053QuNb0GXv8IbCo99qlo6zERsXdO
RnW19lqP/MBq0hfBPtMWZun2tLYNnHHQajNR6tXXyNhGN6MnHzW9qV+YRV72aQjLyZI6J8KrZr4h
6bjqK4/zVt/fgwmiP3Ea2y7mAmcDElm/Rfyu0S3oJKkuMbQb4QNXgSEf0XExVsBsYRI+HktLRsa6
tFN3wCXblg3MKnEMUhUtollzBPsN1I3g7pHsy+/21PUujJ56yL5pTx+vjapFDjA1XBFyn9iJAwp+
BCIXXrGshG1LYEqyyvbqC4Js1xfVVVPneKTRZvwV3sb3gVBvxY/aCY6Rf2oUKIeU8b5YbmME21P8
L8YmvHxinyAjG/AczBpINr2FKH+4VX86AaJjoQeQsXl3V8eiylVfzZEssyJX1ekqTl5rytSgziG7
m4+CnpK+7TWbZHfa4RpJOdx2YPBit0sYmX/eHtcRo/XrAZQzyB7Jz3cWBqKROE6cUnEqVLJyBPop
oeMZRIQGVupA8VYnd7LHvzlBxWnGMvOlUro3/yuMYywWL/dR0cLtWaAW7aYnR3cT6ORpjtB6yX1y
iPhzhgAoeNmFzAgW5PgmbFaqhoWfzF7UpMrEj2A7Fl5OGoe6AxPf1TF72gOsrtidqrJwzj9uCAgE
0pQhNaJWBZQ4Qyc3+Un2ScrQnyp668X72r0AxvNodDjYM+xXebRuKU8sdO3PwLHjtjyGRqaC61eB
/KiUSEWqv2FW8udUyfF3pidMkFOGoYTra1IXKK+OuMQRAe2whQzQV1ggQJm0VAn8hSyOh6RJjSgF
rs31o4AyWNokPl7GPNXRXKIaL0Qv9jdNfvPtKKEpmLGznGghwsZ93ehBG3lPEKEgrp026cU4KcsT
G2Ot2VAxtFMZsvmr3/Whch2sFAOaWU1/Atpv/PdLC3UZRcPdfdLBjvJxEug+2lc7hOdw6rLQek+9
HlONBY/c/rwFX+Bo5k/AzzdAgEAI+w4WRqq1f+xNQY04vTlxiH6HLvVrBaFzKKmoZtBvU+gjHO8j
SCjTIDcfy4HAP3tGAPSS7Sk+6HB0rMrPxNrwlZEp+nlImg3dfVjp1vqMzTXElrKp1DRL5hFHQEmX
9HeyF6wWykKBkW1hHj1QSXkv6CvYZ04RwgGSRSYKmP1kj9AcaYGzp1/AFlSAqqRV9b/gJ0FsDDdl
KU4DJIxn7OyTiYXl1jXMkVWxzcf0x5urfKXrr/eetY+VoIjRU+FQc9B/y4P+gpw7cVVtQMWKyZi+
8LqNkr1I0Wp/uXHUfEcmoUOveL6GROLgxiADJYspWbGCL6kdOW9AfSl+fMzG87YUMzalyydOvZIP
KwAppIccgpx5eBXUCsbZyWAxAsemeCtCsGgepR31ZuPwa/yPqOoarKWFTQdtCXKahcvoq5Wkhnji
QlLVcA1X6+gR8mq2+En3rmiqoP6W2eP4v49d6yGrWj0t0S3ORPGZ38ZGdi2FvfYUXog/4P8i/LGm
KnX7cFqoRs5fVm0wTQX/fj8RPPl38HwG9t8t0zEAjMQUnAu3lPO830RRjLZsPMCkdhHEqCkxpCtx
hsuRhxQHknG9ba74vfKc/EhzYE7q4OEK/XsWyrluWADoAy9PZ19tl5IN1aNIwbva1/SlkEMlUZ6f
2iNLuM30lCvB+dM2d1++I/yYdgpCjvN2BfQ4LT+ld2TRc8RO6GjQdS6TgXRkr/n+ajdFTMCykdKj
uY58N3/lYMh0UdKMC8vys+AY7M3WbpHuob8F6RCzCGZgNdy1+0grBTN3oz+keqYbNR1nXs7mPNN7
FlNf0zj7Y+fiBGn+qfxV5qJhHRAP/udU9pM036x5ynDbCVKyeMA11o7MTbjuSpcT56rYdJHkvXMG
nS3yss0RubNQK1M+/C/XXstxqcedRVv16Ae+mLjoNA/RBjWC5h17XB2KgJ6Xpd23/HvOFqv/fX88
zuFiXthdYTGG0wefqel/bhGjBexKddmifQGvp+8yhY+sjlmUWKxEite7/yPkyKyvqDC5aGigb0d4
vyk4ARd4zyv8XIvUXc1wMwAIu05eocy1CmpjTi0v9D9+BKmKa0CoplOILXE59PXHE7syGpQ0HPxz
E+m42wxySeDUDxfLTODWipBQF40xL3avFyJ+OV622GEIP8GoeH2G0f0AUG71qoEhwQXOsCYA+kIM
YlWqLR2UT9LTyXldA+C5tjWz8myd8tdPcCHbRAgyBlwc+nv82n1spty6+XnQoiJ7zWkX9JwloF/q
c60mPJCtXs1C2VQ3qLWsIVeocyYEUxT+06EdypNp2S6UY8/owAE1nrFkoeC/MkLv3xlLL6umMzDB
nYRJcguFEHq8iK2bzjNbYAjgcThBHrHZn/Z1J/PsxiXNxtSFygsn7qDvkRJVNeSa4fFPQ86lgUT8
rFDRPGlT5GCPapDiPHA55KN3wCMpRAbQ4NpeCOsO89baYGAiytm/MohXixP37r/31IuWv3pTCTla
6QGd6tolZgpVEbQTJYzMqclbz/DIQDela9HSrQWEhIi7txGSakVdtZbhI6WmQyiZdB74KEmSIwIz
6dsNKMQh/B/bVCqNmptUiuKxH4Lh6m9gGXccRj9TmoYhGepUxYGp80T9LubJD45HvUAKloqnlmrr
arc1VzhNql+AvM++YzdpRNQ79JQaUQeOZWETgpt9SFqpU4q+xLDScYwNRB+QKvCGimY4m79WGBSk
hWGd1yg8qOc91Lz2YJK3asx+uSgX9lP1BumE8sW8a/qq0LnD1fRMdoYE2AXGVS8gLRR7Q6YAXfqF
H1PCKD+rAff7W7w0WZ+akcoHunZLJl72ugEL9N2FVDfyV0NL/ESnGLx//rSPYzPobT6+cdkwkvX7
LerFDlIrKp3B/5UIUQynrdn7URfyEqPSXKQqAuBmG2VgL0KAigrmBEDLfURc2o61pW9Y4d7jTyym
g+eCSE6aLeoV2UEIhNp/m19O2YHbPJqYe2nafhr0CcNlRsVfAxI/YK1ZhInpbKIMZcINrQmpWA+O
ctUcx5A0gjhfPGMhz7KjfiaA5YgNhXGq/VUrlXGvTahHTjUhv2VoSAQqdtXQ/TS4whwFJwP/Brb6
C3bCe7FvCslORm2zPAUjrlF7soX8V7Dkz3jijvb0TNmvXso9nSyCAJleYJDUtT+tBxi7kmp/J6Ij
1T8B9qO3nh0mhxMhrvAgRE7Rk0MKKOY5+yH57sY6m3ErGkHBg6aeV5oFqOXCPO6Pp3n7BvmlaNt0
kNIMIGS9daOq7r/fHRDabcz3fGoykxUYjaW8DeFalPcj2WOZV7HVCt993SWCP2CuTZqa0vjeJpq7
8wjnRNJrMuozqRM/r9si5urxvEzOh1gabkqgtaqd2SVmBDspQbnMQEFZbe4zUjVnJEavYXxjVZky
Nezm1jUVqKrGMYzimwewsghQXZ3+IH0AhrXnRLon1mJW2PGV8MkdIyQxxoLAjaquKKxP403rSb4W
s/274ivntWDItz5wq7xiRi0JFu/9DGlr9KxmaQFeUB3WI+PsZzLToUkCfLcIBFr4nw7P/wlgkkD2
6uQhko/skM9TmeMiAGikdDdopRzMEDyBYw/N9peIPLO9WnZf+bEpZWUZ+xi1WEVmRak3wvT67/oO
VBh8+PyHytWODFv0Za0fpTURmj0uVAynzGjF15EjAOB5E0pz/kPjV40ZzPNQ+Qpz3fSmEAm/SYi4
foVOpYyUGPEeyo1ERJj35vC9m98hRFJcpvib3B5wDclQXekRenJ98kLJoHXN2FMX61ix98dZ0+Bu
+11i4zZ6Fyog5D5pq5bHxDamC2208ybYMf8epehytLewgCcr+Ra4jeGaMsRUiyJ0d4SmzT5vPDJL
VE0PoCAbZ+uLOZ02qtc2EmILJ1VTqoSHyYwpG5IUiUv2Wp7vu2xkpuADDkub9UrOHajY+TOqlksy
RWSPN//LvArz3B/bCL3zBi9D11WwSFJOOOKbBMDodB8sV/GwGvyLfbezdV3IrUb/E69DS7vkJjN/
BeuO+iDfkG6v8VSNMsVvFmz/96JA3BUXRD1aQyu3NgKtY8u/NM3Xx7IEFzFVrbiWz3d6tOxzAENX
YpdrlW4RwuqrLj6d07uLvm6VqoCraLDXMGGZH4aOL2YnOqNsXltax3roOsKrFO4HaUkihyyHdzKf
VMjCuDEBMsmM2vdToW8Qg2oFIXnUJ86xKeY+IdSVNRCmdiFp8B2schIogfBBI8DwNFL1qGSFWELt
ZcTbjn+HHQnMGQH79/J+Z/h7xyaDrkIMrjldQoI+tz8BbOwKLh22k1WZv2PWMyKhpL6G+uDEjod4
0iAffuq3J4I+mN/nBDuCMXS6v+1MNHPP6Z4eVsk+nDoMkozatKNbT5F/123VLL4Ap3/tPJkpKluW
n7g/DlhVInbqFvSQ+L7GQTzOdemZ/VD5n+GysM6Xy0YPG12S7thC5c2eTdC9MelkLr8Qr98PRzCB
bkARu/aOxoV6bgfOzm+ynQ8PmVxOiKFvYp7vScbFZb6SvTpMqvbQhsfYSPVLYcQ4JI/6COGOwoc0
pNo22Y6FH8eyZPUeNB/nT/i/RQndQkkXgXw9PqRhIRjRZG9JraCcnYM6lthgyq7gEDC+n7Gv9bkG
Lcr20z27d3/aWT3YdTzLahhvuFDt0ySV8ED8ds55azXOzR07a5XhDdCpFVBv1GKJd61q1S7tDSqe
Nnn491eSnYlK+4ltXxtwBbbLcFShrSeMvMiPqnydyG+urLtw2yLICDKfRwKfp6sFKIk/GQuLiPag
9pBojDQ9Zg2BSSfHaPZ3EWQZNiKxiz+aqm8iZtM2gMWgpL4h4zpEiDJ9qvDOsTBKqsQEJO2pa2Mo
Z2tb+rQAquZOBL0yhNRwUf7e6KqfNbshtgt0YNrlDq9V2m2/TPVsBzQ1S06MZZKLX55yt1PdmWko
ZWAv+85A5VH3yc0Yf0JtNsgksKme8BHO9p4dFKfopP7ct4cmRZ6fbbksWS4KIx5+3oCnTHJrG66w
NwDyGpcAisScwOvwfjT+l3ikKGlT4XN06ubIqWgZ7z9eNy/4ryZ7KkGXEYkZxLD2rDGt10nblsYE
ngzQaTQ48t5PkrZqkVUd59mqG+UAewjxDUneRA+HJCHnk/A9cCq/QWM5XFFk/Nj5Mgk+LMCydcoe
4OMdEy3pWyxtQ506gRMWXkHhF+PszlDfV7rSUod4x/1AuBxPFQyCJ3XU1/tXHUQ9cBw6PF2dd3dG
ZFWaI+2YTRthV9trL2LFLsd+E/G2rYnUXGuU+VefHLGQj5+UjztDOJp17qvQduedtMQ2n4e4yJNF
Krr2uY3osdi0h2PETSxZSJNZKFdQA6dd8L0jVCMuztkYDZziwVtacyfje+6G1fJp4yJe8/hKUNTo
IweUhpi1z2ja0KKybaVTDaJCIFqR7PEZOoBB3uKTBwDz2oAoH9BpmTIvq9kUhLZhxkIsR5QnDrzQ
5Vi3XHVuLodnc9UmnJl2qTqtL+TU8/AG1l2qrrN9iK8xzeBsJgrzqCz08qeYuBdrJAqiLwJTREUO
5+Pm63/U8HV902vQQ1zApYI0Inoz3rbsa+NCLVup8jCuace0I5D89aDkPKWl4ZoptBWHdSZVqU6z
2Anuc7IfgQxbaIrpQqVZMfDEbllLP9XnpuBF+4q3UYIyOyTS1B4k5zTCeojoWqfvOdkFfBlAHn9t
SV1aOUUVn+HlYOrYhJda9uRMkUEskU96IzjG6/nbSzPCJjbOdDo+HaMexWaMgOMLoRKSVrHjbLgk
nSgj0ApZzLIHNRJOTxAMPYEbyqlkiO/vr8gGOqPM3CH/O3TBpH159H3xa2tw88Y78oN3EHaq2xVH
/qmNuDN7t2SYmbF/n1RWbhBvMCU0IrkLWjKBpHU7cRcYUfjpbUeEXraKt9tk02JOU1gM9qk1G43u
77XW8k9gNHEObdTp4c6GqGZqLCK0J/E2bTu4+njDRhfxTPsuNIv/lPUguFdhKj2iJeNDcwts4nVd
Ouxlq9W/qvfdBVW7W5VHRTc8sdyXBIhu46p0hR0rqlIROBrom/N5/41Y/6Xg9OoScxLCt1edJXUR
UwcrQOVqg9Xhfi3zezIDnPixYYGeU1wiAclVDR3CzVsmInyzAeXqJpHOF/5zptDYPy0ZQuldZUd9
qf/tbQ5q7byaemk2NBZRg9VHKM4fyNudndYSN+f3U+lkQvcObNMNeQRHM29lTeTzyZEn2nFdVNJU
opgW4fsopowhOoOjvlvnSXdBSOPqvRdlBDqa+/l+Lv2QKlNMLgbZ/D3tId48VVBPEho5V1qfbG1T
/jdrMWYW1+eFFcJJ33okrusYS8/vvxP5Ejsx0mjoEc+xjrygrqVtDhQBzQ5WUT7qCCqfh5m6gWrO
G0vVUuhOI+rlA+PyScxJosTpw5as54ZzaZUfpo3He6CG+q4u20tDSLQSUiqY1q8OARXN6+e8q7/Z
QEhwKd3aBdS7oLGbBuahjK7A3HjX9z759mjmKwLCsKFmSk72vs/dZHXAqvO7CFnXn+L2CchVlRMT
y+9nO8F5OKgRT+t3GH28RY1fJcchedGKBg41i1LeDDibl5iJ7nU2BlWsfRVp7RL3UEJjGkSR9gPm
ac35dRAyCKVFtnWzsEkURq+yuGIS34pdUEfZqVck/KfvfIVA3xUyUXV/eDSQtbmkAKcAo9GIJ04k
fH20kDkdVXoZYqbPiVVJNJFp6GB4qgdZjhl639By50XEC/pnKawl6MJvT3f0l05H5toiAC7gjsK2
qBnxHrvrHtQggSyMNzZw6wHI/9T+dSkqsFBOwtg8unlMaTY9FYeJO3wBEi24ubzWqMRCOEBdo/LG
lKD3qW8w4S4Wpdkq4KY0fBnays6g0qo6YlB0kCovxt/lXsqHrY9kH7MbXENIUWzq9a0cuzOA/gsk
zuAdBOmaJmjGMiIQijukUmulB8HJoHQXS1CIiwMupQDXbyikyU62K6DG4p4NEf1G9w55inCtSLCe
e6UiuMpvgbJQFLQv4utLVNtMR/oUiRKLO8p6h/nQIAodCKYm5hC1ZTV9enTF9v1qY9yD/tz7f9aP
KoucpZqdlHj43ps0lM9w+aIpn47ykZiGrMagNccYC6nJ3+gWmZ8WKi3fv7Cx/aVT5Dn24peBC9kh
x9RHU9bhQdjgQwdioen10r5vXYGd2RSdOrSKn5M/TV6osxUENTmGzobIRk5P0d+h95UlSzrIvUk/
7oVT4rypyzoAuP9OS9oXu99ACOEfZugrU0H4i+RjDxDGapl+eFleOmqTrz/DBLBVKZ5peFnGY0zQ
MZ/9UJ38/Nsdc8NABWY7hZV8EUQdsP5e1aWabe3F6xjHn3bIpwpc1V11sj6beEq0W2R9rUvSPmZJ
i2PdWrq31zznzA71NkDrSNs34g3hmz0dhphHm1y5xDxHPotSSMD6b8T0TmMrXzons+hhwTzaK1jA
xmnzET2NuvrGbjCk1+E9CHXmMn4vNaaK8FLDIsNjLcJS583NUzuoEAjalTaCN8q7IcQp9JkC22rz
Z1IqYUQNL+YmliquxN23M29uo6qbC8XdwcRH75J43opkUgY+XKaARNSByeo1L0yk2G2v65jSZGG7
FunI9aKWcS7Cu6rMZxHvPk69+2hUIkVfcWnSqG5xSXTM5tsloGtgCeA+odYW09AQQVLbL2pvhVzn
mx3aevB3gptclcvODkiGn2NG7OsUSjjawglBIz0VTJwcngcib2c5p95doYpmDskCKhfoMP5iwnBn
mPgfV+aJ8BJFMP9rBpcJ2jnk/Wm/xiqtM7XwVP2UPii7iI62vuf8V9pc13PFjfmFt/IDDvxedVNs
fEQeoUvXv2iuUxhnXX1kbVkoU1blm8TG3CJZKTipny0XH/2vqWC70ZxF2Srqkr/8MMsYJdLhh8ms
VwnV4jFRXfrMMaWaJJp51MlyIzQ86LyCVKu/djDMx8q8+OWKSdfhCfeW85uPuY4W9ptbV028JhU0
H88Ib9+UGiSJG5fp6zPlyd97Zor5RE6T3b0N9482Bos38mbZi7jhkhE9Gkmwe/C/L9k0WN8mcMdG
ks84enxpay6DdtLDysqHS6n8cb5WhHNIECDJFUnPV8VrQco0GRYmXsuicHOOueLWJ9enhQAooqbs
Y0dfmY94OlRpUqK8+f9xaIu0FoCOKucb37F2WH49gwxsn6fLssZ8wklHM1G4p/MsUj7I2n+FIF6T
pBZs3UOq9aL+0K4sAI7PzAt2mVf7fZHaIh0ZtvIkj0ImuPOBCUrJ8rrb5qYgneVze1yuJyj0r0cn
zOKz1osT/CQUnif82SqCmuh5duGuuZcw28s9xKYhi7xHYKWUbDBFNopLe6o0iyTg0tAnRdT/M6Of
FQJIOeBq620a1dt6L8dQ9R5iesGBueS3Fw+w+yqyxfdo5q8mxv/ySmPiiSXQGg01yC9KbMJ6RWJ6
KcQCD9BdXYB534QUGKWGcAXoQKHXra8wNCVF6uUFZM7u2R7PLJycl94B5eq4wUr2px5cX0Z9g/DE
cZTc+4zJNCH6oWajc9RlyfPZpL4ivp+GhouKGxmtCqiLHDNAHq72yNSeFdBTnHygC+N8YayP+n8+
vP55jf1kIhQxXNRB7F8c+ido+x4bFvvIwFVHRj35ACXOGA8YWjX7b/AyVxI/uLAFc/EPLchVaQxo
5Qsn9c/gxhvzmlKPDeCITQkkYY8nSWhqMJS6EcyVHSCEBVg5CQs5VY7x/gD+EH+OOHWfwqhIbIRG
XCYEYpra5UfXgkiF4CKNjoaNxuA4X0hvVsRiomQp0eAydsk84AU0cqYtCFeyGXBg0GhNXfJ7YLAf
Wyau35xXwf+ye1AG2Fc9w+u3X+IBeAMoaplj1qAh7OQQgK4vwYM4Cfios0BFbZcX+i9+WemXs69w
I8bHqh6CM2dpGrTbPzgHIsT0EAlFzVxFFhrUf4kyIWzZmMriqnErKiBgMx3Bg9JnWSIKMYdgJJPQ
EkSZia7x+3+Nl5xmwyTYfOwMbVEK/93XFacIKPSOqRYTJ3NWvab0JebrGaIu/76y5chsADxdcPyg
wmk6Bae16ejk+HHr8tBd82DPdCScCPv3ySzUQhprcq3h3of62alHL8TSQ7aNR6ywfeQ7OOzTiv6h
NCMA+6y4ELoRiIetCy0FEZBjamSIFVfkKjJEHnNlb9x9PJGeqPAdgDC4ksKu2+kKVnyq+sIpnedP
lw6bMMFJEh2gozcwsEHynpioyftdMWhzxIuXnnevL/KUbvGN/FdB3QtnYhJ1PnqKqhhVx1Q1Y779
z4P5hrox92ja0D5WRkDAyEa5ZsWlskoqtS5RjZWX3L595hvHoAB6QjfBc+w21bB7UibTvWN9Xxoo
h/RObd7X7ThLke6MEPUsPc0JBOdhi0DGuPlaQ30LuG5ovFx80Gws14+eSrc5M1aUV6ITWULMN9j0
MGOTWZBm5iXPpUuA2LRjmzsbK0aCxhZaIV9NopCgBWe/hRr2IEeLIL9mSVRPAA+SqOSqe/rn87X5
45a1tRegUYWDXlf2CgJ/zHu4wID/Q98hNqClRNEiVIDn8be7uVxETIdiEOudgGwOxx4h90xl3TXd
jzboA9KPMmSa/JabeaBZLJP2iA82bjsTZIwvJ978QZ7kr8Gh/C5DYliyrUnGbr+imBak3XOCga/7
ukVU1ydX+8WhtQW5CGg5PXrrBHgaIDDJbGIBvcKrBqkdvtFC0C3H5VZqJpOmXoIDHQAc1QfM1ZrB
+L+NxUVGPuLhGQMTEeVlRmssa2NPJtkt+gfk71XfdidLXCoYHzmmoT7yJFsw63vmjU7H/0Af5PhJ
qm+Z4BPYQ/s5fdFfiaqbUJIAa7njGMNxXlwFRU/OBqOwl1H6F5HSBjtvmG98tKBwnV1E1Niz4IIS
CUhaKOAzOqi+uPZEqv25DYPYj636cTOn8upZbdjMDza4aPmQ5b0tnluCQbW8kzgq5cQNcZvzhhQX
kzGZM+1qRglwh9jYXPyo3uJIEn9F0zGtxrtW/v4riYUpA6eto0P0yrUKugvlA3ItkoIvCVZMzhra
ZanWZvA3Do/wZe/Hz1cVtitu1mgOyhtNFsrvbkuL8ton6Imf3XDu+3R13+MmFuytWDdn42az+B8N
klm5V77qrHJJc7fQnNJE5Jn1SsZmGrqAlJegYyCY1kIXXXE4J2tvUC4BKw6oLEmKPas2GS23Q3H4
l9E1t+ZM8KwjMFbQMxAy2+5jmWu/tH3u8lCEph04KZvoGWWXY0Cpzyq0EAAH7zHP7HGz4PRx21Y1
G2qvESfSknnwvR3gg3SdNWA2hAaXgsAqj4iQtNHwKRAGWdI5K+4j0+zN90Hl72ynBlZwBNFzxfEh
zswhx4lNoREcuyKjzaWL1PKb+0aRe9e2a3F5RiDzgLRrWaaXaMliHR/GD3TtHHwXqUGvbOJO0Nd1
CJznhZZiknLyb0O2OVqgMGGdMZf862H+BWFdOZrPROA9Kdwfd9d2Oyo+F2g28iDgrk9GY3RuBlET
I0AOf4DrcliBNRccMwlcWoPjlukC16BQM7YsI8/NS7rxpbtCYAjGWuXmuNzexb135kmf/jCMD+Pv
YnrFIrTC/+vTVv3JJN4JN2/1dZjbMHn4DOfsVKYwTMGOvFcBSzjsKxOGXNj+lTqZBdoxSvBsjK5r
oLDhOFDQQAXlH5evPl13+TpdPb2f3qJmngtxq7CukPy7j/AMP0MSLiAI8AKhSk34Jq7xEK/fxwqa
mRKt0iXFwMY+6HYHKZ5o7npST8Aqeo2OGPwE1LHhhrMYq6ii4yXuqXefOf1ybCEBsT7X7B9VjZBS
mWHlaP2PxYe+BQYf8hZM/5MGdZQ692RYeiSMrqQeIjRdM8lSp8Z542FPyJ44yklp6AYAnKOMENON
OZO4g0Aul4EE+lpoWcKPQv3PzhMhRW9b5Z9//x7G+39SN2lmJgkI5FDe0xDuMJ/yp9vSQQg4uSke
x8ufucwntbxKNQgl92B6Xg2/GNwWEqZS4Yzaw98GKFEeOrz90SA2q9tOLNvDExU/H4Nz3wTUL3WO
1JY9Q+HI8G7m+M42AvbofnOu5j++hahu6oI4dhVghTzPdUSlHV0m2fZ2P33M1dIZvnnWRHTNXSF4
2j8gAxvfZtvWTDOG41D8XGMornfo+K0DXlajxsWI2JISy3B1asdVJ8OBahrwfp+bgKmQZ6H3dz9F
oBgCYhjt8Y/XNqR6FGp39szYDrAYwWVK1YQLstfnCqxU9kyN3b99+f3nT+I2NN2kZJ/dr7O9NIhW
W+2/pMEtTYrrsC3SbbyaZUG/kdaAvCI1Fb4/k6jNxR6zZStOC6N9bGmHILvLyA7sz2wPWRHb5Iyl
GIfbVnAuepANym4jKP31PTU9pPGSFQGJP3IARHwh4iGZlF4OQfXiRa9dFUQxn4glGUPmsVWF4ckM
dy/ZtC0v8DGz5Sxv7hR+a3KSNsvzfi94XxPi0cAGmh1MVknjSmFgeei4prHWXsRiGrTpn7LsXqF0
2KeqNOwhGqmPhYQOyYQzDf9beQq2mOoatc8dT95oVDWdyN2JP3bTjIRnv91WFagnPlL/TKeYam91
HuNEF96hiGz0vwvscrxsnnOkgyBzHBnh/JkqQiEVdLfufpTSAcNkmo+9KDJahwTR4uaDRPIQOktx
ykHSkL3VRk5C0+U7OfkvvLJ/BcVi19i0Ru+ZN9UR8gg/Opiqv1pSvdMq9zOPgB+V/Pl+GnVlyi7T
CtTDyuDCAa5vGhjxTBDKJuti1b5mJWK2kdRCcHPO9Knt+OYWRzL3yt8zfQ/u9s6zRgzUPMZBnFYq
HeLRt1y8jHcDULQgXDSohvl+V0+vAr6IZmUOTpJiDWtQ3BayRdMyTVmvGXrDlNyVf/calIHWZUSI
Y8YaXUop0gqxa8394exh1mXqUcAa3MyLD6RLCEjE0QtyNRq0jrDYnwyi8IJdMenmp/6FLwswfbnN
SXFayo4mzLUJWDSzjppPRkP/KkJZdUqqYDrbUzYmxE4VTLFTF78JYimpAClSaAuHao4EJx4AJeQr
3wVwZWI1sZqo20WRCCZhT/gxRL2zYldFeaLtikJxipjtM6CS/g36ihBnRVl+Ixj0DFbA25m02OQb
ITYYkBSeXku96J3AFtG2zckyl3gasrOeBiWVg1KQBOWdUPHkxngfMbCUT3nZcPANi41IgdxrzJtY
iGtUJIiuDiEnWvGZFkSdcuPK3MpKD5NA6SEU6WKFSiUP48TXoF6716Z+pl2KY6pQvdxszXIirrSn
mnrb6krKzI3fPdITXnS30o8cQtmdpb1YRr4Hyown+S86gvQQtOV0HsGyiHoenoT2wG/gNes2q/dF
GM4nXT2g5QuBZ24fcig2apvy/NFAAmVrTktvmln83Gs2eM43l949Sb323rNRlRejefN9YgylUFdi
L+X1zD4pmDWa+P87z5LG3MQVrw50OIb+uFqcXhc4YuYBrAo8w/+aA5lEb2ngJ2RXTLsy7OBg/KNx
DIvoH6PaI6voN/IIKYlh+juNZgrNA/GID+1bd/wi/fUZ1Jx3a8Px0ovKoEy/frL4O1ND9vLf4UCv
y8BKcEotobH2T2UXwZs9wg9bCCE8HrJjiBrxaKEXX2lBJ1lHTdtcfQYV1sTLVX8w4eXDZiA2uQL3
QzZsdhY5g2Q3e+uihORHCdBse0orojeFHSXiITqsH5NuQ94yPQk/3HUJBoS19FdaM9LEqyloPhdH
9K1VevfPStyrqTTcVX1QHiZNf4DxQijSAhcHEW/OvXmm4mqvzrX2uuCv5tTdyqNetwO/8yq9Tfun
VHL8qk+BIJRxgsGpornP6xsw7ZAvwLw716TbkJ8xUXhLdjw/ksdhQ9MxxUeWB/ozQGwMNlaBdPSR
AUPUPCpQa3kONJejjlfWUa8qx1/xRfJjBz7saeBhI+3leRpopfZ+hs9j91m5mFUNOgdUeFat8PG/
BeYVOvjU1de8RUF0GCsM5hK4VHkq3Gs0tEAa5UTvBWBm1EEseO8Alb5AYZ46LOLFf//uoJkhFCZ5
cwU0iwECLlM2ki2gNm0az4mY71JPraIsMGuyHuDIsy0QrsVBaInwwUvLAUsY1ijtINPGQ2OPDhHu
BUa1OFrexrvLiaW4IY2Q7d5z1GrS7Wz4Y8NZIuuwl4q81pQ35fUeVN1FTYJn2NMwTmaqigcx03bz
KTtvz1q5JSi8EXsaPjhqc/MJ5HraJBP0RkRkc4c8gWVVahn0HMBt+6BnqmWbKh3npIKmlxiDnlFx
B3hlmLC8Pt+pQwf4FCO5FC9Ty2muBTzamgtEG4E3flFW3aMnQtYeqeWCtCBdDpxObWOO+DwrEAFx
AxXdtTEHIY+mb4ZxjhUoeXhaNOSaMq2HZPUCDf5W6NWMkRyZv1s/KXBG0MtIrQvKvv0gTX99xqes
pjaMRoCwvV6lRLvf5g7K9Fgyu5FPnB4TDPKzx6YqbGQdrDxGZFdjf+381nteVPqS9A61dQVJ/70b
OTATq8d6gnIZTJSHZNZyA/p6smdIDMkmxVlwt5jhd/WDGUMUXS5FG0ultJ4f64lHjqNNUz6l3Lt9
cRbogVk9TQl+NOjCY38a+kAIuXy70LMj6pY9jxgRvZjIsLU9kTI0TFmDMF4AdSna7vlS+DIcSQsE
T9T3mL+QGUwHx5g4zf8DBT0wnX92Hm4LCCYEm8VpBIkf8LSHGSTUw+h2kGRsiPX5QC6v41g/K5SR
2+DcX2OE5lRlzplvjXIrdvdxTTGCJbWxqYXwZ5ZpdCdjAoLUvbWZYZyDs74rEG1RHI+iq0dZeB6i
SW6YYDCRi8ijbsznQPMXqbCneHop7m7N12HLUIGl3HENbZpk6Xlvutg/jLqyl5ea5ySzjkL/p3TB
TpLSBhZGtDGzZsg8ZkeWdmvyKEMDrQaOir5SGi6wZj1gOMteQarBWGsQI7bZVhB9eLoDY2v0vMI5
v1MqtoQmDos0tkm5TI8BSo2tG6OE/B97mHjLE0iLd1Cjcq7yaIsQbyscj1TXyxurhkNZGwFKSql4
RC/kS7FFav7ihx9vlALCibnc40sGopcQbokTmRBUqYiu36mggmlhlnFDVJJR8Cr858Z5Ao+Qlbo/
7ACevMVz0OzeSGl4x/470FdK2MzgqMVfwoEfpQX9QzHmG7bEM5FbjsRUgk9d8koTS0YAQbt+cUUH
2qPeEvs/3Ru6j/Oa5W+GXwzGOUJCk5F8VGWQGcQlGl6MXIQovSZjSncdVgJE7E8/VoSXyMXqzm7E
v/S3cZw+eWs9PQR93QRYVOc+0LfQ7TvMVcAe0J/2fUsX9oMcc8WfPogrx8I9tnyRgydtM5Z5FoqD
YumHE9vHwGW3W5FE9P4FuRKMO9iPgg0jH5pF+71HZj5wAhB1LFFBDaB2r6rp7mII6MoLHXucrJ6T
71MdqyTMiOuEZbOekT0CNP+K91zw00r+ju4Z+RsxX0OJLFoRgwaTlv/Jpiu+MhYiwSw/NV9FmbXS
iM59sxl13HSZ0hnGVABQOJ0qneQOPpn3d4/GWN5fu2FsIUFCfJ/YHuyxB6ofE8XgWKItxOCU4a0Y
y/pMP8n8P6rPvJNh0I4iDrY2HrwUBCHgqbc9v3qZT6sJySwb9+MQFqEXkghh90T0uBrBgWwZAdBH
78llNcp+eC+ICPR8VDWMHlzBwgFqy+ye+TpzWgCYk7DW94CbLhyGFwwX3uHDjkIpJFXWQQM8VUUo
70yuxdk23KHxSQxh5/9F7KbtihVZNXM8+R0o78RWU49PwMiCFTp0o4uotknlxMiN/IT7sujKDhLq
keZ5Fwb6dws+IPvbZNvBC2Iw4/XUJfZ4w5hM95kVPs8VHEbnyC0mh1sEeeOosnn840xAc6e/MnxW
vxRvzqX8I3dlNab2HJQ9XOUu6AmxYA0T44Siudy5cQH7KbMiaOCz9eZZzLMjmcmlCMiW/cCaeUND
qCEMYefChY7MjjzgSUpl3le1Y2y86nmLFglMtXLIFDJgmY1mOa2WIlNnc51GkmiC2oCKeaqSs9tn
zRJYxy2KmV4eXdLv7UNVvpHeaP+Lki//tcC3k3SC0NTnSigkmSy4/cizwhD1IfHEkQh6p8k9eReL
nT8KH8nvr+yrc0Uci9Px9jKixRRrm0tz/Xnyz8nJ1ChqNsPIhXIEuMPkJKOZs1s0C4xcNDSGYUqk
p+MjErg5MxZn7dnsVJBdmf0u4MZ5tPkcwgwHS7xj1bB1FDmmAjOlM2+dYfHfPpB4zxjSvaGGKOWM
ezNIetneJ36b0NcRxKll4j6k3B2i6bRDOgXfg8hkwIDZxQA2ZSJm4rpH+I7IYH7mUQhfVv2JuV8q
DUzOfSW+2AC5hLrJapGlt7wwMngBEyXyqeERvpPcm3ZpGHqRd12B2amrk67h9odLz4/bt7JN5/4r
CHF/UDCtSpogC5iA/tJZxTzzgW62qOfmDuQ/wK19r1c+JU3wJT10I1nqG7icoT/yEiZPHbbYDPyo
OeYra3P+/efiJLXgZuhSbpPm2h2mTe7JcvDq0rhA/IBPuVJ+vY0J8pqlxY2v2ZabnMyt3bFlPG/b
bEm4vLfs/NFIekHY9it8IQVNAUI6LS1ZxUA6UHrAt8oDbL9uVwJhz94c+Ysi0rJUwovjMlZdyKrf
mgh3Vt+msLMDsR+GmsO1A4d7Il+L6WgYrfRC7i1mB0ZqP1NTbRLcuqQSnZzMI7LNjS7drrv+v8Wy
lb5c2cf02KxIX5SeJwANIP9z2hKHynOT9cT4z36tL83ps3wgyyNt/htk7gxQjiGIaLsIoZx2bJyv
N/siE7zNDVOOw0GZj9FfJPQad62IG2B9/600cwxTVERjd594W4YZ2bjjnhydUgZXNsmdUtzn/sqg
dW402qnz8qxHIlO0ITiDvPGGkNISesCiIrNuCJ1O6cUEsv/f8ACxJVjm7Mtcz234pfUGwiQHgh+P
JCiDMtgnzr6qwV+o+X1010z+HgVJMj5d0QV5jyF//IWh4AoWQRuBsbUi96v0IM04Sj7dC6Nm5cav
bVpGsoNsrvUvRt0tXgVmeywsNihwWPQp02XwlSsIAQeBqTb730OwId6vTfWSnMQ5JythLTOy3pPh
jZfUNZKdeduwtFrdGYaJkQBArVbhJhXQtT70PoFglD6zaB/cB5xJidhCGoIrnQKbNXuiP2/gBg7M
Y8w1KJxpc755bvc/6MpZ//n+0LoSW5WB1y8WNn78MChiBIMuJmmaKgPO5yvcESt20yMmJlW5ddWG
8DxYcs6rKTFThzTmLN5x4vfZfnfZmRfwOD20YFYZNRaKdr0Sxve7jJ12IIzhU159HPP7ds9KGVqJ
NMrawHangsO5oPOWremh1KfFFZBaPp5hucdCDjXnj/10UvITC5qzfNXOjhb8MSeu5idhudTgqSB/
hyeuThk0sFvL0JA9eE/gnUQg77bGs/+fHHT3WANY2fkU4BCxf2mUoa0UNu/30pd7C/uEcM5rSUTc
Zt8AxnUs8arMNB0R+rBMlRIohb/CkD7KDrUZm3hnJwZHDz68Lw83LrBdKvvM2rtL4tefa0qhH31z
oj0rSbCXmyy8FkvMjHvZz9ob7ZrXtS1jFQSqAioEasHPhM6LOevvPNxRkLj8rOxZ3no9xdUpaayZ
MczH4a2eWYDz7QnLRAl41RGdteJoS8YAbJBxIbJJ9fmqOhN8nAE8g8pMmrowDHiSuUWy/lKomO8k
0GjkfnaDvDMg0eCH7TojaarBN5ylUZ/8+QuwcWjEvcUWN4aCpWy0xa80xp0nYur/ENdUOt8YqQDV
TqFH5EzGA9MOITOH0+gnFDrk9JNajsfaqkRk/+LXTLGTD4gd4rhjlifX2bww617Q07/je8lYjbGA
myZ1qJWz2vDGOS6/peXZp5wFjEHr63HCyR6LeLvBWl+omG4pF0+h7qp63FMXPEP5VaUcy2+okRKG
xF8hhsKFft4BNUqWcFGeMqNaDg0IeoL/epz4iDemeDxhvX9fG3dV9UdMniw2LYnoISlakeAlRsk/
LeN0eR3WGNI8vdvQ2TojVqzC7zqHLFs/cwro2jwGInq3s0bOhf1NXHHhlZKHiO1OHuVSa+W9QMPI
0gbcBqX0frTU8r9XesBy5Asaj9Ed5h0fvIE6sr/dCkndL3AqUubu2wR4F7d//wKhYfin8cvnvROg
Zmif6R7t9/zTCnKbKyZEyYbonIyyO+iY7tI03vDPHPjobhzouOd/yessAvzSac1JK8cDHxvJl5e7
riqID2l3pX5JQ7hD54jCJqjOarpxgvEbgVtSgSgFsIGLSnMhmrYsEs40lx7RW8nGLuH9d/NxCGlx
Uirb7acRgcOFyrs9WI8K076kyFezUkyWrXzwGEtA8wAEOdsB1OEqrcYW49oXGZuk+IMlko7LPv31
I/iGO7teSrWosiQzGb0L4thzaMq1Ywd7vtKMmiFSiGrnMRpCZzTWz19N/RGSb3/VQoNdspXjZ1Tl
SsRZWu4pLpjDCZOaAIHSjWXXiYL9Tkh0mF1t2fGZivX64apGmf7tu1MfYToRJKnTOFRVEBct8lZG
EpzRyJtfPyKrZxDWI04qAAjp8/0s3LmpeSwznJjX6Zzk2Apf+Z599qp5WtaYBbiH9Pa59RGR+Ite
H+mC7rogPHw0QvWkTIr+N6JgTXkclbeOWB8BSy7H/AgpnLDYZRujHrMgYL2IC3AKN7sFfVVaRYRr
EJnbEsYBFN+azy2DTxHQxmWe69FmkDq5qV3lfoHWBm5KV8H+5EQ5BtSJMTNHVTJb9aSp9GGfeCP4
wwd6mjNQ6XbRlIcmOuMcLcqVTHBa4ZNrkpnlggFfd+ZS025xaChxb/E7o2vrGaDjVTMmYo5yzWFQ
BUrHH6/2fF3wPcOxaSSqzdNOzl7Wy8q6ZyLgR6i5m9DZjG9pxeI2I/ONs3+a46nh87nsnXEoA4HP
zjwJb3JZXbcMB7NyGx9HkUusz4ZTmGfnGVrFe2iATzDhHvS6nzFcMmFjzzOAYVQbQCNYQO/1Anpr
DkzQfXYzwA1vKkLM7tJxZMLcjL+hRAvPh+n0vydB2TvG/PqPDF2Rwj1pBYb70s3OYQ1EHD+WHoLN
RlMLrQ4SF3lP6NmB0kXkp1x44wwgnzEhnQ0ahtS4glC3nVArugkZSHVruL0K3C2FO0XmPiIYdbCh
2p2XTvoUde7LVe98WauxOWj2s56sjssV2cIKk2Fl6sr5DCI8Pz+WNC5sDM1fiQ70bgP8ex/FMD1+
VsdpaOGyhWmi7tbMiSATyhwgXPN+4IIgetFEWhei/s/zaAY3/WqREncfRva07TNxK4OaoBvxHLbr
vl59/rUf67hN2Gi6EozjUzwhMSm12SJc1frhcqexyqplTUDvGLfw0ipjRs18tF5jCThRpG2wFsth
MP0xbf2oVyBzYjNSqT2k299ErkMKEexbtnzKVcOKf4SwAZQIJvpa2XipiRzpVk4mgrqaRIhKAhU6
KU6IFku8ymFDfIOSyqAtTWsXmk96udxi/DQMZG5pE7nAQ6vwajXex3eu3rLkDiBcRC4LOTGjJosz
uavIXJa6KPMVzx1ne10yrhreXGx+WHElnROUv/PwpD0/PQDwinhjdvOHQt2A0JQ6duxLomOYwnL4
X5b80o2LADidu6JFDUsPtkSoPvkdokTPzygd4TTbck1y6SryTZlFVZrXzS8va2e6HxFZmvDKBxat
QOA/tmJytkUqNtUraH27PuFDavJDWS7cNUTE6ILT3iO72JwzKV02369We/ZNBBrw4eiJbmUQ4VoS
lAs4ijPqtM9AG1120MTzfpgeuIPJSdyV5B2evLt5lgx73kFlZup+FDsH5xZGo07GcW2MFQcb9Znl
RjEKUOn6k7P7UBFo4LOiM1+NfmfuV4ATkn6OSOfx9GLZl2CZcWncJi/OVBNMyGcYAZjKQEMxUUb+
J29xNzpFm+7Pj3DPuer2DroSQ0qZqPGnTjczBgZpuDFiGoL914tF/lzK532NVqUgaP0lOPMpSmj3
BW8ST8In/OAaN6DTokaqOMvBfoF3Kh5bmH7XxcmBXMo9xVfSwxiW5h7JEZHsJR4IZSNIeN/N2tF/
g5gjFkVbVcUl+f9ezODrqHactUw8VEBQ254DZ0V4CcGy7Irx+0GzvLV7b4FKc/gKZexfydsrLwwg
yOlmmaJNdDh9hZ2hHHmbUB7KNfTFfYpHun2dWS6eYrH1SxJJa+uq5ETrQiQ3cD9h1pzs0HyB6VUD
VZqPqnp7upcqRukRLyXwpDsIF/hpPjeFzcmYCByJPd+bAVmJw7Oe9Vo3kIG71+WirqOBQXP3S/v8
Wlv2qQOIXNwuHQmSdEynWeLTW9zh9liYp1DQdZJMRjM39/eorF9k4Qsc6vqcZ6lGIk6wbNCAn2Wj
AbB0Hyk7+Ka/AG+FcG0F9T0nKjKwDJcBmNd/0phEAgXohxs7BqCHgU0lq1qrFqrv9SyX5ayu7Bwe
otYRbbJa1YZRD0+LkjPGt2hJEdR816OrA7FQE637cONOl76ogCOEAm1hfmFrycCwMPs3jEoKtBRB
ugeG005F2qxMojtWS+qOxibtA6rijBhn5AEvH2qijDp4s6+KpTc11dPx0T2kBG+LT4gmpZ0WRk7Y
wEdanJdyMW9YrRM/kGpRYi+UDdt6kxT2tzrhtzlkAOOwKBLk+NRju/yOV6EEh/FqJMDLEoaP3aeG
ayHcaE7j2oT23+LR6l8L7KxuvKSM8kRLBNldFDq3IPXpXrDQrQBAiH/0GZbXlq+2S0PM+BQqShft
jUPuEmwc1wCU3oB0uT8aewtdAg3/NOaRN2e9jioKlap0QB4jOzElVGRu4rXUWnTpM8M/PWnC+w4W
GfsAH+uPkUP11Urv2gILXqRUWEtcrTHNGtG71rnI/Os6mHXphdPGW9Ad4ignWSWUO26MPLatpPjS
A5iFaLNofmwikPwV+sEXAN9uUx73CoocxArXlPkQRbW1YZPvYEIsMLFwaZ7Gt+CvNo5ejL5As97D
58nWonuwbSeIF4A5ikCidz7NhuKOhgA8zKYo3lEkaeBo7IzJhzXpfl1gW/g8rbXRHp/zqjadH72a
+0e1VI46GAE3HEFDdTEDS4PJza2wT48Nt1iuaMZGXLp+TsVRpVK5N73oaxKQzAWm/75PvqQFN1DK
U1BZFbfKrSQhmGNePzLJ55PrbgLGNGoOHf+bLi9F4pg0oTkoTc8tSr9tR+4aC0fvDSlwFH0CS+he
usMnGnQVREaC8ymoSKXqlu+EqhM7PqjE94ok22K77nhVYw4ehpZftg2NL1/5SAGGCWpkjewBs0DP
wBUCF+fCN3jwxlSxxnGLIDEr/ThckLcwsZS9zD3nFbgWWIIlrITpDBy8tL//dr4ZIg141WCvm+fh
qogIK9tnV0APZcWg64fe9OHygC2qa2ZkzLg0bROjJNXzo8V+Iv+/IBMinThQBjmWGGgFsDwbIYXz
aMljc5A6IWqVL/kK/0byIc8x2icqGfvU0NDFO9/UgO4ujWjIlKdyt4S/NY+Ot1U5gMLJSKxAeabk
O6TXkN7SjOfDMqbQOQUW9KzLRwAK5YaCDg0sOik6t4VZgKdtqSJFMvZrewDqiveY+7Suj/XPq2sa
drFcERcRhbEJ0HPMuKQUPzWz2eEPDC2grxRf0t0YtIt9WIMwGfeELlys5vETonbitsXkeHWBAHEZ
JoHvoX+5LtCQb6Sgwrd1ZG8THHCZVnLXmaUAHyEO9+yirVwycteO/TG1qONGDRCPULtQrMnJp6oy
K/F60eSRWw59vemWjNLcE09TJBqIrRLq49QC/ut1GaUCRcwrdqUp8+voynM5L1p5H4Ff3XGXG3Kl
6as9mYHnzXlhKrWTv9T04NAhLVVx/5f1UymCrggwbwIghz/kJxCML4aewC1S0BAW6pE/UOfZZKH8
BIiCv8XX2zVh0/fH6wXDPnVAP0LjM/Z7qa1mZk9wO33QBmLVMBkqx5qGfYpy5qKd33gOsqe8E07t
yvOb+Q2PARw9TnKj049Vfv+OlBgKpWDoG8yKliQx6dgXc4hS/18hipwjj+2oMPrN4fzKpkDyzq/b
jp2pweOR6Vl91twyIcJ+XT5s2NkCiRVUf51MkCIZktXW2pnMpZ2nU1c30ISlsZvvq9e3vtH874CT
sM7QVOPN1sSjldHqfaqb95Je4hOQl0weCLryV88K7IxRnyojy18ITmBc0cQJxCLLee2bEJAFqJ8w
pzpZpqVGyYPOmvfIIEvjG3NZgKkyjmo3T68uD+U9rcTxL/gWHtlWntb5/9SbT6KB/LpapW7B2pXF
fT/u7KzBKIs1ILjzrMNG1kOJV+P9f3KyUO+ebJSFkh/fnzK8jBBaE7FyVZhRcHxb4l58WgW3V7f5
21HPUwD3/J8GkUkEr+RgsS6oi3UAO1x2VhXQkhs37S/ONUPxPSqzF3Kk5K/97rKUqvnhC1BEMW0k
v2cuoswgUbHkceFzh1Hjkqqj5kwMSeoc7B03IH62MFSk2ElWhQsnthXKgtH8pzRKytSjlQitWCUp
Rans9HM9otPLdmQ8VvLcRUy48K5x23RaIDM6qDf0rn3inaaHH1xVyfSYbKHPGoYyh3VB5twIate/
5p/mtF3iXMovl4b3PdIARPZgJ7vBHgz/G3huFasfHEHgVFY5zg+q9b7EQwRuGFm0827AzxBE+UUZ
h9UVMq1v5MRp0dZHscse0d5ey5A3D98IK+Qe1fhbtAkVHSlHKVOIM9NZ8WtQNnJLkp/5OTSvjun6
h8FQpX36EWPKIgNC2vsYzCnkDl3XdVoYIDe0NvYDIkX8mJCwIJRGpXXWogH3K9yyWWeSeF6oEmmw
UKHE533YAFDjQuasMP1/hdLJKkye4UGp6lUhj8P1n8crXCARU1HXfd1TQvLmFY4Jly4b+YtkNogV
h8Dy7AhbJNVtokx0DelZSWb54zVSVXHQfRexzjMpBRFIG2Uv6XbIqqq5FgBs0syB3wbtyTv8n8gb
dAZXrUJHk24CzS0UuFZdXsC0rrFjq4SfHWJY3AiLr2R8xb4lZHLIueDMxaFgCuWNDdH5B/xKSjpW
gl9kxPGkxvoI2J/JJFACqo+FlrfTrG6XRp2R7K2WB4klX7+U7i509J9YUd/nn0x0M4cQT8x0n+Gf
7IaPDrEP1VBCBchGUjp5CjcmhU29caVxivr1pAwU1GV7kz3kEpJ/ltPLKaMn0mm1QWet3W1VslR2
nUl2ORhzE8sAQW9TXKk+aEN7w0n+BJ4P60sqUYRw7nkaAmL/uUsnCfKZJ1kUwh6RlCRssGRAMOht
NBeqeJHf8kQIR8yt3AA04oqXdqGndKn9icqBeu8aLWPLfUVXDEi0RnwmiiLGcPZsVF8+CSk693l0
LKizrWpQWAEzOmSnhbPQjMOUkcRsiJrcK6lRTuihYsKy3dADMt8qGtGEkUJnoQYclLUSfl7ON3pd
fz67T58QlSNzDpZrbpDXoE96OEpD9DK9RWICBlQgCsY7g8PZa7kYfMihL5BKFD6b9t0t4lz8jhyu
PRJSVazEz6oMqNt8ejbvKLA/uPfULl8dULaoSG5u2sC/tHRzYDrQxtfK/aCcLErPFJJLsif5KJ6l
dIoCK0ffZZG7ouGOhw2ZRXKmHa9E5BnxPy0cfsk9uorHSUNIPPxA54vETNQSV/oDPkn8CaifHvxz
KXEKYqzHq6NZQmuSKVUlptNT3RIYHc0SLkUle+++ZhQ+lsX9VwtCvwQD91+6EgUM1/GAZEYR7AUM
igpRVagiXERx7zGSF0ZzP557NeuEi5aU9EH6iWojaFNz5pXXXnhVgEpX6yJ1V7Dj6tArJ6CYBjIG
c/rrW6orib0BV837tn2SEhkHTwW27XLH0UhlwAPMvNr/6EDNXl+L4NpgS3Zx7JSmXXKXO01VXKG0
okHsfjm2RuTCS7TY7RjJYXB+HMxVL+RkZDV0gmbpZv4tMk3hpgWBiySfQ8jsJYdzSilxHCYdOSkt
XtmuOh+YR4JB1b+4R9NixCgpOo+gh/5B60nkDSWupMY80cWsUNkkNu+Px0E829gsdFZp1H27GJ0m
dCvhshN9Ycu6pk47TDbu34xUrO3/glsjo+9dp1Z408eoV41BoX7D7AR9jdBbh5BVtUD04OLev3Uj
tGnQG473r2pJXXExhiW5yUIDmFc6UDSIJ8pJtPrLHvW/+ZE6WT/IPjLPlv0ac3yhj9+OCm0Q5SFf
mmC5+0uj/i9BoMCQMzluwdCfjgCU4hWMRV6liIO75Q3qM9nmpZnpNRMYZ/SXfn1MqlTeTyVu0Y+7
NO5vdEaZNuWZGvpKEdABhLXck3VnzjDxnIP1+DZCPi9u/kUP3BBGjyVLBksaYraqt+DIgD0HlMzG
qzNpaCYN2AJ96Jlvr5PCHw1k6AvnL8ta07dZdyM4vFLzz/y/sm3ug9hafMvOMMnGk4R9iP7Jxqhm
Y4BNzivs6WcjNObc+DPW66rMWDpS0/JYggCvMzpsaNzM/N1ic6t9C7ZwioqALgwiRPmSCoQDapdM
Lv3XAcrxSrev7rMAFo2TjrLJPl8bPOfb8Ca0jSNY/TKaOakW1i8cpajKxCarrBCeiaJZYlr6hMaZ
Fqvtms8pG4BHyc3qXvW2jBsXZ3IUqPf0dlCvoxraGf0oZOswhWJSaSG7c939APS9l1nOsM0Xp8ww
We1zbhATl1vC78GsU3SQWzXlOiBplucDxSuzlRJnZkwTMIq78bqengQgcqA6zydRLHuqfsUS0d21
GeyGwAo4ZAmYOzmLeFNNiAg0CDfNa1Cb8zC4EbmJMoyfDK2pa1/CuHTeMCiUpWzq4LSqEOXcDgpt
5p8TiUsMsYlbU48d27yR93pCm10tINIcANN9f6sVpnbBMqwmeONbf3Y5hlzXWTjEhv5P3K+erGPt
jMIZgLtbScqZ0F9TcLDONnNWZQGnopYWMu9oYPAjIJy6NYLPO8V+SBXf95S+7A/6VuWkZUDI4krP
33uYVRt4P2H+7zJIPa8aMo5YUEc7SifMFvmJcuIXz25nxud4d9uv51eyQJqrL/HoqL7x8mAZwLQr
Oh0W8wprXSQ230TSt6Hx5zqVmHIWCcYrelPkcBIL5bMPf0ZgShZisw58UDuY332hrkGAfXRe00/y
tCwPXiBUUlKSFsOCLGOPM0+wgwleutK/iyP6clniHR+uX7e8zK35wGCq7BgG5qqQ7ZAlzYyao/iZ
cwrf3Au4VNX9jRby6aOgXcTbGt9sM0NQ5ny3+K6XsrI/eUultPpq5ujeheZpKfOQEysDjw8fNdzH
46zk8J9+eJHu1nXcHf8RyQdO1CHmw/4440tVl3noo+5UUi2M76vsKFFLzTCpKZisFM4TvytwoO3F
u1Jdt/yWIrn6oahP8uSwefT2zRaNTSA+VqQu/zJU4ehg+0sYLXFvCT1JhS4ejj+BwftwovGam5zh
HgylZXLxjg+nWePT2dio+ZlOnC1/q2AtiTaeJOy8w7/GPL8cSZ1sypaBEUriam8szNjkHjurkC1J
RZ4t+9/sBfq7F6CL666qyZNv69ipL3VygxVh0xJKQMFZnGVJOMM7x/X1Wfu9p6Z0bN9RAux7KQ5o
YKtWE19debu607BfBXKz4RRBFdZx8qr0krnmJsPKveTFIPtTFDap64oxNu8TVqUFTA0hx/hcMxrW
9J3XLmxbj0cvDGcEeIzcI4wgGjq2ZgzbdvTNmoe5jHlSvF6xobnomjkwE+EQkGjabI3kOaOgkp1I
VGeCJnlOzMWyMrulWqoWkPyFoxfAtrYBiy+nY1CSv5xZAy/HbVjko82VCktkMZGUC+gc/j1PVl9S
5j3FRMaWKWbN6NlnRCx4FQACZLCIfA2pODI2dYulsrAJN8z6MtX9U4X/OVTEQZ1yGP+ZLSyfF9By
qqMU/Q50Y8mS7fBgq2piOzX07vU+iCpVwPKEse2EEVjJlKwZZ2GEeNkbzuqLK1/0L+u+4RKh402Q
bmVujBFC4PIopYmr97444NH0fgk0Gou4VgeF2D7yLj1Sf6eUv7wKwO3ZdPAJA7yXmpsvR+dTosrB
e+MXrwegG9hdCfI1VTjgtLCr+/dh9H84cu30yuO86xNy+JU6zpYCqtLD1wXfrA5rSH4oU8W/a9Tm
vntLb9qNszJLXGGiSxTv5TCWBvRvsbdhWBT8ItbKFi1/T+lggQA7thThhDJ3MewRwz+GKOWtHWrU
rTRwtKj8a5hJjwoKiG3NNmIbuq89XuvI5jKyl1yvIzelIBNSn/RWcEMFl11aDhAPWkQ1R1SJ8OgS
CIGIriZIu0ZIGhVS+hYDxLY/7SSSI9hiICOAkMjlPeGKMA5ek+tamWUP4su67/B5qaRfwClCTbMW
Ze8L3ne/ONd4edPo0HGzIbUYswuLFSfT/zaNAuVvtThEiVRqB1KkDYB4fGAjBGFPzwGC0NQKcjRh
so1Iku4SMVEgvkNaUL/XSvtllgKF1I/7rjjt1ytFKRzk4kDn5YXAkcesxWhNPdkPLliBrrOdLb/0
t1FhD5KIewODjzsszsdK/UJv8QGs81hR7kMlC++xjH5vbeO506N/k0hcSQ8hxPFq2A5pzyRPW8WL
S5zHDia5yF6huVMJUXDYT01naS3aKZsTi5CaaenMrMl97l0eSyOyPSKx3xyDNEfgc3UT3Ee3uPTT
d2xOHkfqMIjbXVYhFsUEtAHCIGA6xTTkx+Zah8ioTOQJNNBVh12VD0NPgZOGhE9ySohaO6Xkm5U1
bu0tFS/P1jVP+bXLvr9FayZ4L5nGwzDk2Vc7pPoNceJStV09LvLYg65p4Bk49h7PhHVJtd/b9sQN
hG7in6C4QeZWaVWybDX3p2QF5wuGvZXVb2A3dvGqOL6cmPxOzE3FSj8Hy66mGh1AM0KSr7R+6+Tb
e4sq3EwEJEof6vXWGD3u5LvtbYH9sYfOJyKqR00mawzoTClTbUj1CK4dZHw1+k53AL5z3DrySpiu
X7lWBOnIUXFWPaGOJ3ZKmgz37lrOLIqGKmpa4hkAce3Sd/0Lyq5+odsVjXV2KC1dbvBlMiUVmZp7
z1kNdsA5h9lGIhRySkpFrihtcIn13PZdlp+A5rrlna1eAzQ3Ijvqm+q1YUPfqEVLTXQYPq6mC614
Mw28I6BGZkdMrtL2bfu3VaYeC8Do118u8fNg2spjdZKxxD81cv8Jm5n0BmVoUEsq45XALxtbz7j1
wWl3ad++tY2QRspX9u1fHSnFBqYJ6PECZbd2t4HO43TKrW7KiIp6di6hZxs7Ig8hM6SWZRGg9qOZ
LfE235CkpKrP1VvQDGb+TvyH2l+lDHVernJQPt6BzbNIasqMNlAF0ADt4lRyTeGHE03gV1mLxudy
4moCtyWjyTmpBeE1wL0AywwALzwlV9Zu/ZXiXDbGwhv5LGOjSvt92KmB/4DwAeIa5u8ODZUw+Kzl
eOEPNW1MhZXNcGJ09dpWjZFO/E2Mjq6FXijUqzTdan35gF3DBp2qE3AiEJFJyuzbQPFNE/yykvcC
Uskgq9L/5jHp29osVX8NZa10fBhbPRTatdT9UNRgAfvV35jkUPvbjsXT4KtT0rmo0wXfTw/7/G4G
TL34nz2lO4Qv4/gketdCZ83CpmEyCDmPEFRNlX/AkNvt5adP/sFHo8GDhNkFROdPKdkkMYt0gUQI
YQs1yuK/eIvOH9WKWrVnui95kdktj2/cpB8MgJQXXK92D98Yjql2vwnRI6yjoFUPrflA/oipJ5hQ
HnRlwdg+37O36LAd2b9kqBMnX/b2ZfSupq+U/iRSfvxXpt+hcPXA18CX/1/49zlu3BArexEJDejf
onQNIXnIo7aNZcFw8DQG5oID2xJ58gjSOyEp6gPXIgahmPDmDIcDBvRoFbutQkbHxNRp4+0aUw1+
Yc2MqyoChbeNKr64NWAIB2Na9R3zxHd0zk840SZ5nXacSwOhnPuLKX4c7AiOwU3cWIDyCTYtxZiX
GOXy+ov67Q08LrGAI9pXGmi2/P4Obqx+u6de8+QsIjIHGQwjQJmD81/IzLIP3rkrRaSsfFtXb6qF
1mGgB1K/9/GtEH/bLgK54IpdgL0+Wt8o9rPTVAiHVkocL6ULCmCJyMCh1BHWNYgLhxZqk1v8rZ+D
9U04pUhWEUu9o5r6Sxb9kLFyCflKdWioD4UsJzg9RAup/gz7yavrH8JaaLCMwf7W3QCOH5UlfPvS
g86EuahY40CJfGPaKxshVX4z4cu+G+lFkOPdfP6tkWNIPU9D20uqIHN2BKM1q4Gs93xiCHmHJk6B
hTHKjW2mGlI7nxCgOlKzNhDzzXQMFj1yB6gim3hn2LgWR6fskzRdls+QrfixiiBaXfGD1qA47zX2
y0nwoLw7c4DWSbEYVXyiz2WwNuraxQEZkVfNJmwhINUQoDgX4X6qjj0nxJ7VgbHQx9SYiw2SgrsL
UK/VYNfspdTL+MqF9Dmgre94McV5mZSM22akYDwGGfyr11phECCmQY1r/Zq+GcdzNN9hXoE+btbx
arA37B5/7z1ykH9UStstThZmcNhzTJ4VN0O53kL2dIqjA7R+nndv6P25Wp9tvJDxYvv4NP5ANPbz
oBaqp5gY00QAJJDnPzoLJootXhplEHafeFV3hirg2CVc/eR+wr49xyJAKNMTfPbj/f2oo3sRMDUu
pk+daxBbMq6wEnwSk4oKMf1GWM6uMokGpsQZnOEhpeBZXvt3iae1esAUL/L7LzABnT7b512NxNAK
4d2QAxPGx4vRTtnea5ATP7oGgpT/tb/7HHeiLZdXeTmcMaHoSaIoXtlkJjXOtRmQo0l53u5RBtCo
IvkI2y1CSrN2OiZJcWgTLa7RvuoRKRg9PvAIn8t/2ea9sVuUbcnE1CwvnZOQ6KUSSJ+d/ZZjIQGH
0r+SWQjx47lB4q/AS7qUS8lPz9mqTTvSLiuCqnay6vRpAoCTcP09AdDiOlXhYq2QcUes+Bc0zd6+
A1cMQJYzInqu+ycTWTibIhkL5NQc9O7VkLxTnFapUKPYWCbkLGnwam8xcwrUKtNKlh2NKLPQ29m0
J6XeyBQLBslXnAx39hLSCZ+rG4Ixmngjj2lnt26oRVi2pb4k31sFEX2ktj3QGTFeMDLmBS2vVbvN
9NywEb3LDje2yf4dhUAV5FaUW0HbOCsM1XOaFAY2jeHtlDulwShBDHtHkL8bhUbue8noDdGKeSAJ
5XTqnqVJmSt/btcgcZDPyFi8hU/IOXPijv9GabHLcFgry+IGih4ORYeEHi8k99JoT2RcHTrH7Gav
RE1FxJn62ehEBFOKK31rMrY2DGMk8Q6NJmtq8p06Cpa7FhjWbASY0494Pf7p9xVYiMlIUjYJ3qW9
6M1G5/0yVR18zImJLIYFJCaj4v7JT86owfGqq01lb088kbNoQHFSTp/rkY3tZCDD1XlzYt4dDKGb
KnEpVg1xHm39y/Btbeo0aOtSFQT0LEIxgMdRWHpek2Z6qQwpQLG+xbfi9GmLrKGPB3sP8HmTwM0l
ucVribgRU1IJD3ccdyoPZvWLvNipYFahxAbo9bPifDr5B6R/FkrftuvEyhvLEao6ZOwIL0CeZZmz
oj1CTBJhnY35n6Dj6YxVq6tpJbPBHvPqSjr+Ox+QR0oZ3YoeXmqP4SSANZumPt8rz2WlHgIvEwgs
pJdN4zPSs394jm2ryybG+IVJEJ3WFfM6fYTTsV3hOYku33S1VfW+uTB+OjONrdJs8BtaeEr/3TOc
jKXOA+nfJkLcWHb4SaJtmqzfxTM6MOtzJWq4nx6heJVuvOWO4cb7xym0Gd10UogWlql9Dm3q2xsx
DNnmJ2QvaoiG3Zwb3ZWzMksRMvw074xNIfCSB/RXbNgBm0nXYbxhQUIho/L209uFs2F8GG1Q5PeX
gkRHlxqtREdU5UAIirVx4MxuEdV6uNxK8ZKFzeOc60Xv6mxIbevyIN/MDsGRHNcsw4PNcrYxscVJ
RZmWr3VqcXshYEdQVI0MZAkQiCFWE46VYf9cVgaN98NPMDYQLNjgSDM0XK7muPniw5GxkkXYEClk
c+GG4LRlqZb1ddXWJg20K8tEkycrid9PK9SS3hkWKZ7b+FtwzBkAIyzrtOXqhhkIINOtuerh/U8o
9uApuQ7OQAzuhEyFRaimg97yEAcnYqIoJi52ADJakSoCMlzKoelrICbOta3Lt1SrEyAgW3PjD9zF
OMEnfSlqhP2wDNT4g3Ivou9P8/fzNv0uH0BnBqvgWkKgUOCtoG300iEq96iCIKPgg7OKa0PW18Gl
qe6Pgzq964gYfZKqAsIeC18jtBXWZAXUS4DtXPc8UzqNacWrReoKqFmQoYwhxJ6cj5ZjS7mgxZA4
mamvghE42nTr4u54IWIjvBfcaaK7bsUFdu8hrO5NAjMlzlduI997yhl4yYFF1B8H1XCEBuuktXuQ
QFKiAc0FLXU4ldYoUDQpLKmSNKoOYsSniRGiIX7o/FHpLiHJ5ipwkGN0/CERzmYRfSdoPCGjyDWs
HYZmdixOu3YAd5Y2ZHJTpCJVxD/xh7ibuWaRf1iXTcoP6eE2W18UvjVJbaHWUDXF/B5KyfM1WCG7
lbephJ5AZdK/cuVAVpql396mJMpwtJtWnk2rKt8LrjKLMlouj/KHD/STw+hCdqJfOGzt8qAKWPB4
tyko7tnQSJq8oiLePB7OKLiXym8h9PPPNY15wXA8yvDMlaHhenkalM5pD4CrRDVdu6/YppFeAQXw
aBSD9+IuUZo8ug0cDQJCXIsHIKrbutGXacWOeKm9W9+T7M60l4PJmupv0o0LmocIPjdNOvVyGQUI
krM06xGzaqXdiuTpSIua4mYG/lsW4CI0ycZ1jx2JkNSchVTP6+8HJ+ZV7CDJXVT6RsBJCkXcWf5V
YjRks8glQ3AHjYP6ljOxG963PufG08yP+OWQCG2e4QROvq9e+4kiXCraYEOR7+r9rpCru6rGUTwk
bx1k5No7iCVADMC2njysoMDat0HJm/sn6tnkvhpr7W1L5MP8HtCM1VueutrmRROQPsOvXlfh9ozh
2z+z9mD03cd3QW7/f+8dNla7r5g599DxrXNshtWqpsbRdQ2HUM0oFptiojifR2nQut+y0rfRJDVs
hvz++r8XW+n17BPnOrl7euxE39eFrr9TFO2uPrbh+62Obs59GAMnrUkpP8SlLxMTi69grQ5S+sHA
wGkMr5Q5BWtrjew7LsHoHFBpxQMzxqIdquBBUP4v0PsSxLtT7hUORS6C6a/dswHGOoZmvxzrAWOh
IB13YKDiFht/xTjzTXDca1GA89mRsACJzw09lCOGxyeZl+VzggP47R6wC0smV0q9ixn1GS1GqMM1
suqUDZxI7qygqIVDpcpyfB1XlUWHlACkLmZsRw+3yRVP3WyoCkdMpC4RQCP5O4crK/3Wt4TfH7mO
AhjfrpfMis3qiBt0NmgCaMp2jwK3gx0bgW05JWusmc6V4aPKIH+0kJkiI/pRM0oySG2ajtwjSyJd
8utF8/x5RWeoNg2uQG3x2i6I1U9sbhBcHAMGmzImXK99wgoS+C/PuFPBJ8lWb3sVgSrTHp8lK6ei
/9XiINJPgwK5LCpHZ2DEPrpy7pFi8goOZS1YQ/dv1vjjNA0mDgm3xaK36ghr+cAL0iY25bVwbDAj
bJVtCzui9ZDlLM+7O9BqslG64enxUrcSOtS7q8Cn5iuLi6UNlF3QhLPPLeDqtoOZPMaOAD/N3r69
PiDWT951eV2i8NDSfcpZBUotaQjJiNIh6fknGJ/6GmVn0MAwx9ptcCrt8oQ3/IfRZdkJ30teirXV
3a6ZkFaN0yrEv/MFmenoGyWufNEvwOGu8TC2QpGiARpmrTCLtU7SQxVAdH2BDO9ysqSMo0eidfdk
oM+7E0MBIVMxgcItyoXgo4Bw7rxMP7UVRApNF8QkL1kzEiuqgUnPamD3g7qo5+Zqi8+ZUzlA2jtG
LhnysMcOh4SbaUdakLKlH359KeqYi2GGXsblF0GJWMKoHSbZR+VHtzUQUbAynwvfZnDHrBiUJBcb
Z2jkc7fhCrYSNSzABBw/+09CTn1lxLH1d+ivvNdxFIjWFm+cNfUVNE6lpQFNwS7s/3xK8flfwcms
iA3kyrw1oR2pU+DPRHVTrjMZglL9nW7l1wCbURkhxGTl/43gmzlgOU0fY24IS6haIe1Ou4AqD7Br
tB/X0TBxtBn84OXi0fRzEhcRmybIbdMokEo+wln/CIj2A6Q6lvZ6DtPRSJV6N/78Jq8FihEWJljt
qEnu23iTyNBDFld44iqK3hPz5tPbHwUVkcL2riNodL8fZ4KjbjlNcFFvjoHvuFX1CTr+XJLgY3qF
X6UnLbOsc535OmlKAdHHrOspP4sibSMtVmiYxsEZAtsmdRSo9fnzVQTCeA35FKAN5vCKM8Glg3UF
fJj2//gxKLO4aJ/3AlSM8xVpEv46jARMS8FFirrCN6TKU6d9aibQrEKYmolFP//H9V1/eVS9M02x
OZXf7Io3WBDZvPVXWxKUqF9B4lzT97RHYRiwKHZDbDsgiWe3Fc9NLPzNQhreVCXXjnzcmAHQKcMr
suTJXDUSmq5I7k4P4b/Q9m2UKiz8rHsjIfu0SWiuUfwXrRxqm3PYxoteHc+eSUYnwcXkPIAInIxF
zPH+Ne39hiBDmC91GAiC5SMIzwaeCjmpX5dGNV6EAlq9yoRERl8jWQ/9E7AZPOTw92PJd4WzItXm
iudYTmCcuaIQkU69meJQhWfme4AGkQSW/+YGr2TixaeVC/k3DH0EMNccKNzZf4ud1Dgm+aqceGIv
Zu6FBq08Y2BR68CDkXKGmJUkK4NCYtIQoMd6p9fO0zpt7ma6kWf1k8JTXEcc6bp5dBJLQikEOnvJ
ZMWcaGT+9rKAM/omHut9KqmARNAMbOJFdDFynQ6RKnoCQeb25B9JTXKnl8/8HmWsqha6MbLkp0vc
trxVc7GFnLUtBGcapPmSb0ztJinbH+okz8klDy3EG6g0XHo7vYRFQWLSsJbUzKQFdysql7Ncnn1j
prstYIS7uLXmYdUH56EYG0VbC9m1a+/i6GhLNLusgeMWJfSUy9oEoGgvuzhlmoV9CJ42noYlzFgV
FvuXzp54DNNKCUY9C7T0R/aj1RZuibK+6LRqEIBV8FHwlf7msY7SGCRn67OC5zTJQQmZL33QF2Iu
mOTgMGPAy/KYwiJW2aclW/u/PNT6pEfqufg1bmiDLQYhOnAAeW/FMwHcRTzwgxsINLFqi3//D5uZ
6metTQoaiS8jbqjkcH98RBKowBJC5dMonX8gHFUm8wU9G2c0kcnBbBgWmbQwDle5L1eTIhMokmt0
T8zXYF62O2JH8RYbkvLOBHVLHaD1A8cUXox9X0zIT0V/tty/px3LJbqHab/DfJRwyGOjdpmHbsup
leOJriquUu5aHQN/zONlYtTwlBtNdwSlgGOthOztsl2lpIRKPDWHm9lFwZmq3L0JnUtSnxLommeS
0g+SAxwbGUL892Brzvatf1haQE+GkMVO8HKgdt3qsJIWH+ghAwyWeDpYdyPmGczRH35IUeo6F0/6
joZNDuN7DY02vI7LcQDw9cPzLq2u2ozeq8nqCvqBtSeRQM/5c8aVYoxfQAY1K8QdA6mzMR9eJ2Kx
uz7/pupZFJXZsLFcSo4k0gifyCgXCjRzAV7qmr5RBfNp+9uwRw7XHZn0UtLuQmFAlHf/Z/l4HqoS
r0gHS9L3IPOxuy/BXgbD8IeUqLQvR3Ial0jQPI1rqQV/PAY6B42dDKbZRkxqQ31sIX9KPmKxC1IL
5KjKhy+M6eKOPS+7lyGLGifr7dicFdNSyKGtmlZplieU2Q5G1htbOgnkmIw5DHHFqLivPpVX7VhM
u7/66m/3u7qAiJfQf/qcWyAarUp+9xP3PiBPjtf4HfThaTBlujYckJf9G0GS/GQed3YLDknXuVQV
6ztkwp9NbsnLKwzZayT2idlCPEWXShw3FJh1bUdxLXAhGjYHq0wXQgBhjSa3/Zb7n6M5cNaZLahR
C3Q+N/+SOkJFBffqDFVRapOS3pE6X35Fd7INnxOFV5oijscnVlvWnRX4jJxPHNx0kkgpfIAa5SDg
D2BKYxgZV8G1W152BAWKOlIMcSQOFTJb106rp8zWBnR6MK13hvS+mo+b+VCiI/ihG8i+3kHo1RCR
nmaosoo8+mhsPLkztUEL7HDx1sc8FTF/6dNHhjHb6zJnXTpdzBjU7RwpBJg98yySH+ILK3UhiRzN
JOlF4HyL3Rumen7e/JXpcQWdr8xL+zLGLjjbffLUV16STCkudohrPszr55/aC9xm2TOS77Y0Lg9L
GWn2BAwJq9u0SZFIjZoGn3yEH7ClaTxMkm0HuFgcosKtIwdtqHMJkFtqmoW1B8+oRXTS5AYsr1sx
RrX1DDMwTrW9p1LBAAJynK1Tr3BjBlVVXhFrn2ndkA1wi1w7t6yyGfBhuSvDH5Oxb5rHEPiWWRYp
2XW6YGzTL3DMUvs81rehWVAKKm6Xszw1NvFXXSVsPLIlBrNyuc3yw/GZXR/hrLtPt9bRWZjp90D0
Dyr16p5PfWmqwJf409vWVkQ/ZBDIslnF1uSOfZF0yNSU02H6eYJI4kGorC6BUL0KxqWxKHhf9v6o
Vwp87liqqJToHv6+GHr5TG0iWbURclovEp0lkQ/fVd17i6jx/cmH5f8RKZEai+Zeth2EI7wnlGpJ
5VdlLHjjhTeb6NaQJkKvZB2UDxXxrearkmAF9w0bhD8xc86BTOG3Bxuw49tE+oVZwUYJdGq5JTnD
ovjGEezo8L4hKa54BzTFXTu4ObJ0f3P9owxCNy/pq6dNqxgVJm9yjvG16VkDOKaXq0gCjcTdgWah
qcBOhnH6Rwzgr+bkYFUV3GPA3VsEAScwf6hq66Hg51bNvFEwP8B5/aHHjm8W9Y6rYzS12SFuQy68
334hLQu7WKMMYPIqSDLbWjjbgWOeLzkfgW8N14xShQ2KbNNHagyd9ZfAzphpSVQluwqR4V2MAwZ5
GEvmOLdQKGcQzWDAuTNnSwHjO1SA6E6dTyHNjHB5ghVvMEKkt0hzDQPWjM9HxF6HZizp+H2BHfjD
1iz1WWQU4xi8FJCFIFG16BYEnetG71lQZ9pYNjbs8IjlA6RHjGAwR5FyCTCl3V1b7fwPY4s/ehF4
d2x0kMKPAlq4hRpV+D9OrDpIm39HcYq5/98DQoWW7NHOOHEw3slMGoxlWf9CdySWPyPdo8gy5BP9
mgb7WP4dwOEVc5ywgcNMHy5KeffCuoLoMcMaM1p4Z6il/xYseGS/rHZZSeYsiuydMBSy+a8YDNFH
MSx1dvMJlE7UdCPWV5JBT6ew25cLJnDsdC6qMN+OQQKzce9R1SajaPZCaUoNfc/lXFksvFVeL+UU
NO2CGbUXSKnDucEh9Pvtik5WhoJkMgt9L02arvzT8Fzcwmjmz1Om40hmWL2bHbAJKUJc+9kUB46X
Vpr1MFgHyznUL8J56DA4oZjxJdFfKrW7M9ZTSJa9DhALUY4L1wt0ESJLUEoRF+g6/ERM2FSQHxdh
/guuvw0c8Xw6sRSDOBGyULsZsRX6zlYRTBzaiCDwwjIUr8cL+L4HS04aewak9Lfvn5zrKdgWGVkw
n3W68w7jS47kDVJKqb7ABQJk8vBU+J0YlZ6IVsB1LGd7NtI+IloRSOZ5rR1mhoqa9PD5Yk6VYOeF
KWoof/jyhpDJl8q1ulRDOpSU8Id+iV/xVGmo0FFCkFgoWinJXkaGppAWDveYAWQtzEkoyuWnF/YC
536bvAryI+FWDxJOQR6U2oywNMU9mRSVVOyXFFcSJt1E9+kEeurYde2jUp+xqbMW8QF+0fO4/BaF
e/uIT1kzB0kywbNVdc0qH71h66NEo6Pkxj6GqCbcIt5fzPOBNtZgPmj8/oE5dxDqKWoYPbBNve7S
4Fnp4uOv9o5Zn8LL/SDugKn7OlgNrQ9pJMtwSI4JP4Rep1KnAK0+ftl68whyP24Ji7BS8Axbz0N6
ZirufMdOkvk10H2iclrH7xTixwGYzec3Ki0w0mUAgFJ2LHwO3CpfWI0YBGqbaC4sCJ6dLEMfQ38Q
qO/lSRHbhLDyF7Mwt5L+O0ni+sX2YQsUNi4YO6ocFpxGzloHXP0mqCadb7Tlg1kJWPySYUDE4Q6+
fsDxKPSe5IWY6x5OpabDIqWmfE2KK5takozrlL6eKfLC1sxA9GQG9wp1uZiXJiah05vsazlOYyM8
ocn6dLgKVkbe5JMaPCihDRNuj1y2We/5WBKyDKRqSn77GhnEN4hvhBbuASsnVo/pCuCV/DS75MdZ
wSo/8vkLKfMjYQ2bXt15uvBIuZSfqDXWtOmgHbclzPwSwPGQAUuuoAbyo3UL2IlewH1FS+FYmMih
mvQ+Kn9dLimbFClbpc446NqlWHjMKvq4bg1/V3PfZ6sJbQr2QN+K8ACtz081a4+CJkDmSEeA7Hz0
FbyuuNpu2jvBIUe0eGaOopX66c+x9bH+FiOPPXUcArC/h4FpHeWiRAcBZ4rDGLdcOOLRe4HEz7jZ
/VffFaSAF1n8ZLmlxtOy+0aWeVA03KqabzCVnRhc4MISJHmNICyGRBbHZ/hnU8XxmPxZASbSZlFB
sNpLczu5J6wQ4Mxcf4lc/+RXhSpSBCTVk2GSfjJzOKl5ZTv4grqjH3tAd3jgocP5CtiZ2iGVTBE+
sby4/7lERBAsj3H2YtRCfe+03Om9Hmq/coxZFY5HKGC/VQjFqRxYXopRdtw4fU9P0A7YTDuF4SlG
cejA6jWxEGQHJKSFSPfe5vN0t4+Dt/MXp0Jg/jPbdJ6t4InD1d5OGxlbcPAYrCUtJSXxgMzm1FpL
jKh3m6T56fbJVf7UJ7Tv+pYA6Npu7XFSRc/AMwTsFgGPM4NeuyZPTzUaSFXPpZwgVhKSb/fi+Qzu
g41TXYTkfmNc55YqS6w8FxyKrPNuHq7N2OyE5/YL4vEYM+t6b2Zm43KXo9C7wCc7XeKxXZpgBFup
8oyVORxqEh27K6JgStmSslog3NTIPY/Q8danGNBU8X0ZULCoxNlUk8kit3obTrL9NZwRAwluxx6z
ejINldRyriuw6xs/zGNJs+5UNSQwOEb6R4Ouo6ss8fGf0cdPRRcD9DmU303XLbpBGEv2TJIP/4Ct
18J9dV7gZq6giGWHxsx1N92MUXDEiD49BTD2KJ2kqZqcss8facUfGKSsKLJ/pyt+xsVIbieEPnPA
SXqFAvYFp9675FU5M8XSyKyo8dupznuKdQ9ypDor2mhBJ56gS7b86jSHC+NCqwiVZbL2Hzu3irJ8
7hlUkJWzVi6LVC/MF/F3/60upv2sr+GZzAlWdXedRaNQdbGx5G2NS88FczH25lUD6Jy5bwwiHSfz
VKoDQ781P6vs/Xzqiammht7WLVcZmpZqaolMK2AuxsDjFLZZnXGzcVOOZVBo2jf2Z+pwGk0mJhb/
UFtHTVtCg1mQxcJUUtlQYUfk+soTYrF9/0qbj+ihk7hc9nDrAvGaVh5bj3Tbpu5AKkMoH+PmGs5q
CxOt+ALK+4LsSLaXTTZ0Yc2z3lMpkUH/1LVxb3FHZm+1NU3O3/zL429NUOOa59uyCiFB0BEmy0mq
jalKApsqyoXRXeSA0lYIdHff3phVU2pF/c2wvsBZ1yboCoMtDe/3aI/xHO8s3TbohDbjYXg19s49
iETHX3PHWYiol3HHbEkprs7tNv8+5WsoXf/QxwbWCFNrHVfgVdftonvaCBQgHPc8kcRtdKDNdd86
D7PeGTd0cJvzXV8zfJ/bIsB0/Ic+ldwWIHX2CdZ394rJbBccDH6+2WHlZuVx7F/AF+9eHATW9a0K
2MN6UXe1Uf7ToNF7vqUiSKPlB+K6J9uwCqJHNqO1kWbst1bHVv21LJz7PhONPzehbgXXNuHrvff8
MoLpiAHXK8bwUURF/NP7aBW0ate1/DK1wm5kK8ZqSrqPF+0FvJX8d97wlaQ4F+sWTJSvcemUEjpZ
W936ayJ6oMYbhSwPda61ALYU4k6yMqNCNB3aQ8E150Cl9M9moKmWbpUmixW1mzs8JtS4t3doAwCQ
QbZnIrwZJiG1rxUVxx5VCKb8//YLLZbUNvxAS2fpRkQfEDJAU9s1B3gZQumXXGZ0ITRj+bsPWMKl
8Z9lS5PEcBk5YdNRjF45IPtfFkmwU9NkixT5utEd66QoKDRh9ELydwl75aNPbKSRdeox+ImjCEj/
UabP9wzuqM5dMMyaJfp7/aaSPWzXMrU4DFMBncMD6c9OqBSJrtP6KDb8PUV9BnFdnoUIVyshSTAm
mJnkubMzwTbC/hUngKDPj3CVBLF0+EUFDKX8fhRQ9lOqRw928Jvr2A/GWqbjZ/l5UKW4WKJlwa38
3TxwDvTYE47FDB9wD0uwCVlxkvZCpwIWrk/JnhGoB9JH8FO/ojRP1VHa65WLUWLJASxERkhWlTBn
ChPJjZPwTXZNIV21pC7avZGlQ2VdNfWQkhoQEbQzcJaRGBQK/JjS9hZXMs5t+r8kHRb9hhFu4rT0
CrTlBb+cA/iwmQFmm5i6vf+/GX7BkrMO/nvrKTsULwQ7GbHXcp2ZI70+svrN2OQKpenOKecE1IKw
M9Pl/1Rrgm+e9YE3FOO7VnJe0pp32l5Md09DhsRPRQ28MHwhoQ0luo1NIuvuPMTaGS9Ws/HDo4AA
lBRZ5tGL3RoGz08YdNYurX1OnsEpyuaYKHA+RVUg/tQytrpFez8yfS+hb47/t3438pgVt/YUP2jj
qVYwtUFAvq5Wpo5Y6C7A0QQ0K4eObcVK9QGww25QOQrUylj13j1ZPb7U8p849XCQYCs7jfyG9ygP
l6sKS4vTX19xkD/05SKWRSAT7jLwn8BAC8FsgqDXPF9yoo2otSdWlH/8dnKEbjwrGxHX2QdwE9Rh
tasmN5AGROqdsf4zbNj1n72IeTtGioOS4qGVWxaGYJYiuw0u4XFwfMtPY0hTa9lOODB37TnMgjpo
1YZji3w4nL2ZVnwXF3TJ5SW9OUOvTCWyqDsEXa7Sh8PJiR9cizA3wkAGkzwMVX63SKoWOrl1+Epp
nBfe7/6TZnT9pMGQgc5M6pCmN+DxyBF5hoiLvrLxRPwSy0jFq2PhiwIYj3y/uCzM/VOlBCmG8oOM
SSRSA2HSGLjUZs6lFHTvcR//u0ZqqIyp8EWj5sGI1Dccjkj+gRfCTdZaD1Q1oz+3sCOhbzxWV9gb
52x1e5+bUIsbQ9QNACAAIjilWE4LsBoeqFT/BOcT1MQCZOQtXqbqnzNLijN3GbudJbu9+qWEPUNU
3jnchH2/kwKQ74OgbI+UHiuZWsHQo5wpJdcVwyPxWTV0zk2mkYbnqoclst55sNx+tFQrsL/kJgJe
rPkKWsncHBEnNUcSnhdJGVTk6zbcuXeI+0uoagnTknaAG2OcsaDixSLCTitTfwnVfvoVLx34OGB4
EBszmCXhhmOBedjPwLpvg4Z3b3LGhjOl2b2GZhTYcJoJlSliYYh4IEZemdflgCrVqDzJXBGqzygw
0gLuox2rd5UMQ427LXmWs7h8RFge6kbyiC+9xJptqHFqfkCC+Zs/gRywtgXyNa12zX4ax/HeU3a9
WAulrZW6PytJyJLzAQsU1sH+3NHavzX7dalDdb4r8W3u+y3Z+NqkvFGBCBqkElxsOoK1E7W4O8ud
7xr9HFDQcu7oUEOUcgspgwHuLWRjcc6KbV8lVOjl3KXj0pUx3IHzLFISfwLFtRvsb3/vWN4YK38y
V2g4SQiMYhmiLNb4TkhrADRw+uXVgZpIgjhj3kKYJYImg9WvcX4m2VpgO+7qYD//4ZrFYG5n7n7x
Lp0VO7tLYyVQIVYinCNDvLB4a65fyWbV5jdYvTX6D9S9HfgXJELedt6rzsJxvUbyYTMdeaT8VPFt
U3+KxIvaAa/qQ6TChP/pWvkRUg2OuRc85Aa+NcwCgmH3SOPnIARe7eNyWgshvDcim4c5K+wIsxIp
XKGph6blKSeFXuyhMy0gi84CNOwiusR8jQi9JUP4uj/oqRvuWLANqaV1aJDbLuG5Y00iYAQaH4Nr
iZ722eG/83CSW4QbXWutksHz0N8Uv4ZF6Or4Fv/wNAvczIyowchlxWGTLH2bg6irLlmYT3ZZTEpi
PS2gsfov4UMAFA/kqXxXfLcZYvfIZjJR4IeJv7EmQ7XkavCLj0hl4Rvohp5PAvfXHxI+A38J8x03
ghp1ksNqvHhGJ6oTNxKb0wblWoAZ4U/dgcNa0y9r+t9ujjhqf+AjXpKcxtbUQWzCntklzm8MSL99
uAIFa1EEZrJc/2vAcH25zlobL4tvctnnb4BJ1sD9T+cViUGvvv5+X+fkxhT6VGGpxOm1kKmB1uYN
XOKUiwLqKphMekRIfXoI6Yb4MhpJdD0v0tifQ1AwIX+OETWNS1veK0Tbw7GKvR5CeW9Z3VilgCLc
Qwzm0vwKrOQADPCM4VWOatnq8SjfH+qYx0r3IV7yK49moRp89Hu23nJh1za8EPqTXp3kFDR1D5TX
z3AFkb1eq2Ctw+99Ww7X4e7Oxn3hLD9puZTBLWN4ZqjWxyJrgz1i08QXtqeawVCLhVqZOZ1KeQ8T
mLzKxqpz+wFm1kxHAkstbgb/YPmZz2yWVZQn9IpmyszTwyHTlYZM96hjYxfcb1R7H0ZfGRKccSvd
FrE7NBZRp9fwob8GOTQkX48E906klOay6ibENMU/CLXdxnbgbSPWpJTMyPaHjqHRyMYV6abGSGVm
QwXb7pG23xdTYKI08zh9TU82It43pyEKBg2Wlbo15nSTwHbSvT0WLEgdWBQLekI/natNWh5ysur6
Qj07uHglLziGQZ4iSu/WerHh4JQHhreKlFmU6W7hu2z69WtKhs8+y2kUnU+z6t+PhT2CRrFDl7dX
GVTOHPwG16+C3e3B45tQlcGIBYBR17gMJzlEq4ys/5ynUsJerUKkjXPbPQxu2b7b3c/enUWkArlL
vjhO2hyejnA8vjc4kkTk0C6W/D32za64OJ8vl6L6Y96xvYIBAMb2xSWr+6AtcNgbPhDz8ePTYTk4
alwGD936EHaWbSGXnMYzKl0iZDeyIqDk52QZsMPZA9lNdoqHzOA9QkQjMtZCL87CDN2TE8bhtUvA
e8Fj9YCBUugoCzPFN8JbqdkfWOkM11Ppr3m3AO5Ay/mh3QBqiu5tYMx1EEh99vNFBQf1s0K0ohZ3
mvgD/3LLFMYrHloR5wsPSjNYX2Zb8Qu/grPpWkW4DyXPPge0qG+IIfmjMGuMBA53LRfgvASQyTTj
A1Xf4kIvsH39XQif1aR43509AQXupc8tkKNo6zX0ZoA5ZXv5FEZUU4pBXDObxChkOhYbyIMWdGfN
RPYoQlessAOccwY4WWZ4qqCTXltCITJlhfaPRIipXxEhkCPMmPpiPp5N59/TNHVOsNLRtCcQI0lo
EBqrhAKNFPYEk6XXIUu5IxFDvYS2bnhER6HXi3Noj6YMR7NWFL21RJR8WaLr0risZkzrE701j/BH
d+LJjdCNdrDmPghvsEk3WFRBuyRpue+s3LPjdpXdisqa8aOXbBCTlKu4CEeGdTc2fEylqvyz9Tjg
strJYXImmnjCWbB5yICxsXLgIWFqoLmPSZ6CVBw577mMZy/RsvTjTWPE2qEA5EL84kczPx7QRm93
bx7AniQ4qVxgAX/RPZEJVqxkJm2iqeK8/AdjmHlsRNuMakN3Njj7z/rSlI1iMRKVT8IJJXB67u5J
rA3mROmzAvsIwypqpA3NpGkCgWhNeOrwJORPXc3Hhv1nD9o5pyBJo7tX/0GUcCi8LCLifzbAL1/t
fH8Exk0Ust1ELrU9O77vLZjO7igUGpAWKUUhChin2OylaNtZIdsZ9c9CAI5fdkf2f0uY4XUtNWi2
y3Je4h+ZMqanNgvSk68LcBrnBByAf3h9GCKfO7DoICmPcxr5abQ92wy+4Tcp/9PTfZorLOnxfCAo
B1rXC6CnOeZpJdKg/7TgxjW+R1g9Qc1/W6R73c0Pm/R2cCnMJX2ie0EVX1hRwxSmYSBWSCr1okB+
l9Zq6pmmM1rkN4/ICocdsGXmDp0mn7ZeeGcaP4wKEh8zMpylFJhN06BjdcORU6VjV72xQ8Q3aYEE
QDNuL7gGfuYuDl/2dGvh1g1IbsEpWSdFlsCrNgLIOvkgshVUK2KXQaIifj0QOPyC80Dx9yXI0wYq
cDodAx7LMDyWWL0T1i/jHMOB8us22lUrgQmZ4KvMMIaZg5lZVkI21PmlDnAy7leu3mlz1Rx1HyQh
1o1qG0+AGEVOzTXiF1YQ2E2H2zsMAXR3eBKlYnIsCi6cJfo9acO0vZd/SPaxwG8ci5GCs2ywfNJN
fwSCAa+9AtCbfa0vnusuaB87d410oQLuSXcipJH/pRlW4nUMcLygNXK9WVPnjKJ3o5Br43sBdAaZ
7kN29eymebI+jAdptfLpaVpKQypAcMGvgzJZvBnpOBmvmqfhenY9Xj33EsuQ8tDK/P2ou1JbXxVr
/D1/W+nUQfYhgB7CYtXixpCcDM9Vn9AWjS+h98bRx3mwFA/9VbTQfpPjALlgXMzi7+Voa/sIWsoF
G0u1ZeCNvVPtTvXibqjFizarDKYaD5ILSQ4dz6RRoooWKfKw+UG6zKIxsvLuva1DK2M1ESPQLYv2
iYuT7zzZ2UgHgbmp6QdGOqZefBoh5g4EuHydxHNbUYxKCDZ/iWCNQv4vX77k28zmnFUYOGV5LN0o
OuhruZagK6ekkYUXZtXs9yyEbQaHh0unYMKqui/6aXqb6InyCKlyPuAxQOMCwPCKIy772r/V03GV
LgULQkLjWY3lS07l2qUoU6SsO9tEu7kv25cKpiNrmHkligK8aYowmzKanzsKBivYlv3K/wDZfe8R
NftoXmG38B2uuvbNM2PE3xDo+wEFCyf+Y07A9mp68fvZMvvGz78UlyfiGXGDQvoDzCJubB2pLTLH
29WCTyMpJJ2GEp0CAh12D4oM1WoN9Losti9dfiFTccRHDLxWvk3X0r/aD7Yiv3cT4MHtKKdBv8JG
Mtw/69Yc/u1E6fB+RV6SPISvMPjf5vdQQKZ+T0sla82zGfkK8aPEdxV/m9+BwFKTZBMj52vKylHU
IhGjLWvg5k7iygT8nENTp09QYjwWonjnSweKudRMjG4o2BNk+GCY4/zH0YC403B1L0i7WiXJZBqR
IUWgYa54+E4iswTdvrPbPY7mS5PetGhjSgfErSleLd+WuZteD7AuAYLmR361KqmLXN+/GneHG1OX
1YCKcAoLY1E5Eou2NIKX9ozkNV0/pq1foPnofHRGAY2Kfp/800OfVpsuJh2YBgZJ96sQ/V5A7CQZ
GaS8SpJT7jvjsrULgAfT3hLlWq+GagL0z/JaS5G7AUhftdv3HTTX9nJt8kJa/LqxvZHhHpdOC5wf
ZjAnw9/0KaEJGIrCFGq+6chEYapsRSbkc7f80vGtYNldDAh7k/U+SVgxFT9+FcUFhURB9L3egGDO
e4c/dU7XVEpSZymDEN5Z8+J+ix9bCxUA3a0yMOfCaYa1sZSKuiFK94DMAmOkIuGlo2WUHLWsXxEw
yQD9R+E+YzqBSLo2o0cqG7KrxSqfowwc3HsKaFTpqK07Us//KZRs+KfF08p8G6KWaDXQR3aEtrKY
WA9OerfmEX24MY5+vq9xgK2idGfZPlvDDoqFPvpGastVWqQKA1nQIfTiO+ni/y3vtDf71WIVmMvF
chW1lBX3uV+dcTEwjroJHVHhhWI7WHEU/qby5pWODlesro+zEWqm6zPyd2F5QCMKkQ3SjArc5TOV
1KZVVGMp/LBuoY5EB2gavzbHjAb5MvW+1iEnbbNiPd574l5EMs2u/sqXsMXns2aRpPrDlmZd33Tn
YM1rcNHciqQNWMvXrEjBjWjV9H6kzJJepkqnxDQW4++0d+gLVcTT5szONpMocMHhLfiuR02bFIHx
WPky2b3xf9lZeRJDcIBEVuZP1SG+xGgituTC9Rji9fgVq25iLQXlqNToA9BBR7ks0HNc0fH5xSSR
604yV+tx3v7NBMhDE+dnUD5+F4xu1yR8jz9fV4+xoZXTmzYwEs7Alow+enWoRcoMM/J57Ismf+rF
o02rhNzyc/lSFWgII7dcbG5MUFyNPgAULE3PeSgtfs9K9jAlw3B270RESB1PB4u2m0+6RBTBIpp5
wJKn54fNvX3cKUwb2V84RTc3SqT2zbjAwtB77cQTsvt6Q+lz+nQXxEXh4/1aIq/1wSzeTNWzEUeD
G907oxbewTCCaXQp1sFfQLI5bXZazjLqq3TIyxR/w9xKXYxwnTaBPNn5sEN+EN5SkB74F+AJj6hi
WnPeCwx48WQJuNgh8Q8mjUfYrmQccJjX98L2EfEfBOVIzv/ohLkPeKy5v9no5mpg4GQbF43OSLep
r8wVez2C3lkV7PA1LcFOOsFVzkDKmaE6QVJaqJdKXPHTt/IksdvLj+X5UJ98f5TuMhCqJ7duLvO9
ql6ux0zPFdKzG520aqqsW8rs4xAfr+3tERVARq5jhHaoOREI7T9cGLznPY9suONv+uC+WAsPMYr0
fl4c3JdQowlHWlcIAMhDvXlyIZLC7DBbxCBG+Fa1BHTxAsyH+6IJUWnQsHlL6ogC1KkQD3XQBDl+
uf8Xc+4mw6HR0JByJ0ZBlF2APeQBSwG4pG8gUyik4B5GjQK8Zcz1ckzwiMOigdY9a62u+tyR9M4t
QIQWrGQrhOrgFIOrl0G+L9+EFVOwW/3KIyeMYee/ZOdhnhmPZujieTSrtR2a5ZcSvgJWuA7L4LDL
glWBQ1f4BiDpI0E4iPCH4/74B1MX/TeAsCpT7lpyy20GtZ72Gtjdz74fGhb6UWgym4Olnungd274
IizsVkuAyYW5Cf15yCh6LCdT/tvTvTm8MeHAQEMpHnSOmXAlF/Z/EOdFxNecEex3em0nMHb3MWd6
Vl5GVv8yCGMVUf3Qbe4fNuH/RKwnyoNRTxRm1OgrRRfJ0LBmqDMhSCwkmaJyiAVaYzAUtBz4VwZk
u4xzLnII0E6PmJut8qWkX2cMdR+FDpAxaDIIboc2oCtrLvBsdG1hYkaL6cD6ObXUr0E/f9sfXzKq
AbBJAmtc5bz6gYYassH9DlH17+5Nzko499EUYHLqu3zSMlhy+pv5vwV7C/vmdBvuYC4SZkpGRgEl
nmY9Y8LfD6diNBTwpnujckpBrWTaTxkMK6My0HrM9T0A16EGbW2tntQ+5UzFpAsm0VdsiNRlHbfB
uDeYX76TiVjxSToj6U81bdlJZ/FyFzYvKIkELTM4k5rrEf/Yi7qxIe2v9A/PaNBCH1DMpZZydS08
Hgo6Wxydwmb+oVlPzCozdNvc0pTicvFsbXPYK2TAlvg07nNS/KnxJHpCcKxICjUvP5TJnzODOYSP
/kzhrD2UBsj4zLqtCoyDl58l3WVjwz8Hg8mTp4Vmf6IqvM9S/Ib13NmdlCXVgWZSiQ7um6kZxMmH
SfpcFBjoIgHtw1J+l1r4sapCNk65s9BUMz4RrbyhMMALMMXGJTLhv7B9fQedJYG6LCuxArxkb7yp
4sOkdwEMe+Uwc6S1c1cvp7G+07O2yZiMF8pebYYOA5OKLycVBGTNque5zhk3lQm4hFyiMK/hLBoo
pBH/66LVkP1NxrFvA2w7UBEJr55R5ngVhi/kQKuFCg405GUnUJedhp8c8H6oz1vtiI8f85Nr2HLf
N2l+/HvGkNECqOmPD2chwDoEviW36W6oST9U05GmViqbE4ot5VdpQCbRxPtf5Z7BkwbKjvj2wzBT
0k+NW443shURb8ZxlE8LDkcMi7EVsPr7ayOyYDFhCPs2Ja2LXO7h3ucsHvx70AjTdL4UAp6CJgJh
wFO1O0ZGQUhuybiGz3uRLp4gzYPIKmPGmMmhJ2Hlu9dlWYG0KEau2WA5n163OeI9V4WuTN9YxB+R
QKIhXQS+VNTbMHroKCGNH3mvJ8F4vbA6qzCxT871Fvmr23LWqw2ZMq4Mn/C3TlYad4xKxHzO0mr1
CQ4IxzhrhMg+BIEbuByeFMpX2c8w830jtO5Yh7pn7OZZ1GBweIz5yX3KFTMYM34D4ovNSC9uwC+Y
JEFMU2wSh7PX2MOjpED7sdUUva7AcVsHiykjG2goq4LQ9nTIvwmg4w9L+eIbm3l4lH5forIEFqWe
C1EqtJTn5nKAfpxL4mLc4F9jXXh2gQLQ2oNiY2TwVzgqhXViS4+VZ2wHEaSphezGH+tzyXdPNNkH
zyQs0l1XWsA/M1s20XEK+ILzlygwPV6WBA6QY9n7rkJsY74MwW2GcvxwqrwDh/ucF9DbT6QTwZwR
aVKinwLEW+OtjnXJKoBt2cIlXxiUzURX9ErvIi5L9w99mn8FgKJEzxXuCqhSQPtuqNul41iWKjFm
xncqITz7sc9CaTKQYzHO/hZmHfIf2H1UhLrR9GRhg6GCZrww9YtVpUukTN4y4PcgmdbYUiWLx6xd
olNPgvDUoeGNFx94f6czFQjXajlvZUMghioSD2bKmrnmPTkvCt1Seeuzzl7L5Mh6p3KtszvqIeKl
pD21gqq1DxpXqo9fui+9nhNBwb2fN+UQ9RA0XRw6ppxnXk3XS8oB8GZPDRiMPRhUyGMe9lIeZPgp
OIAf59MwoTlA05J04xumDs51P3wro9PgTIr4ExTRM3ADA46wc6GXeDyv8oG/+kvozb/ieRGSnsFv
e5DKO3gL6O3qQdRxpZkSf8bOrbKr4rl+Jg3NE7838hXxp/YAbnOksn2YAr35/RPAZQrPuPqutpuk
UnetdL9eMiyGjxVmV3htZ5+W6zJH0JPOpFJN/0H3V7+Hyx3T7/eKYfr8d4A6/NXRILHHV9J2+mnh
soLnc8ojKxZJPlegmETzaWSK8dvCJLeYc0GVYi1wAAAtPCXP59Arh2OCaFBk/7Y0HaG+N/zdP76m
kEnfEPD1ZNe6O1m8ZOJp/kdU8Kiury8vYP2f3+DkPQ2UCler3gY7Qt03GwH3qbCcREtjQPaYdjHt
l01ni+mSDJkp/eQSDGeGZ9sPKnI5dAEIjHKemSnZUAvEDfftPs+K+aRJsPsLjnrjEncCU4zPL3aR
qinNVdEit/y9te+TvuD97uAE1DnRrVDyQsku9UTTd9QjShRwHdrN/fzlSvthMnXTWBVQvBQl71J4
IqUtyyXWbJl0FLrId2vIlqeF4PFnexyGtORm/fcqUEP19/Qft996v9V/mxk4Vee/Kus1vF+CbqsK
XWIRjXrlHAgawuPKY1BLzxK/vSeZCoY5FldR5R+Fn1RfNMoiCD+ldo0CnCslLnL7S2t4OAZQvQsY
7W13NuLeQjwfrugBe02kmDOkmqx5IWy6NaW097E2/fXI/TTOWDqtIwSMEANACpWN5h/zeBaec8NY
4Fh8bpVB9MfykY0lX0i79s90rBWaURW4gPxK4XGBMDmKEe8k9KuTTQ1MKe8pdCJm3Rxj9oqBnIDh
f7pQY4iLWVPVLXb2vCqORSGZjcl9tJLTMgMEJEAbFYaCT86ZcXAVukN0B+JslZOYyse5lQmO6cm+
8z+d2uTOwCDLhS4mbqejOSILlV6g0RToc95Gz5+W6ODH2eDNlJSeE3qjosFc/QDkHhFH6vv1d3FK
R5vzmf8i1JovLKfJL5SGTgOCqI0q+fDVKS8Ku9dZ1a8+m+/d2BHGyf5D1RB9BjPXKImuSm+aJ+1C
wofZI8XUHPuDaiRVvnJeL6VsGbjIAz6hSINIu3eUk+hKNPaBAz6riyotPER10aZeAQTbyiuiveae
nosZPkyBr0XbC+upD4FIdjVuNOozdvl5vRp1cozpqg6C504qW5qQ/04aRj1kLiUy9DrFZKQpuiEu
4ZDLgKJq7fMIlVXRxgUr7MQQ3/LT81lnDybBQ04CCQM8qDKbI06fYxLsjSW6RGggP6/gKiY6iOSB
2bbQVPO3oeokXwMcibJhL4MHfDN3nW+hhes2gfZeo4I+5n3XTakdrTJw7GYj24ds3XHloWkfOS+e
9IzGhe8EunKv5chJ13EjYJzuP/LOhplVbN4Kde5O2EO7N3wD/x6TvSO7RHJdmBl/TSVO5JAEDfpr
+5RMyji4QKk7SCimwRTVYD4iT0xo3XmuktAUh+atTcpCId9D4LwgjhkKBaprA0wZvzq+lnPSAUTJ
EnkBP4SlGf7tv3K5DMIt/H2IIXtWFEW2b5lLRTFMbkeHmPd0jZonxLTTcfkI+MsLttZz2HZm/3Xs
YA0GbzoZJ3WtybEiaasVGZ5bMT5siyu1Kevd+upe9ran/DursG7bWSPtyk5lWLtzyJKlGdk8M9FG
Iw5YI2LQHwYogRfEBYTrjJRB1khW23OX4BDaM+v3JQRB2K4wm7Uyv3saBY9Tgqo+StfqN6OqLlJ6
AgYmCxT/Z7GW7YOEJBXnx7XYIsO3NixCvv7kDn587dlp2v1M4HFystt2kmcFLOJLYsIYfyhwh7nz
CByc4kBiytE3OpZzmPvpQIUaO8EIa6g7eSmo2t58oDynvJOhJ0SX6S+ua6ky9k9J+lMPgna6FPHi
726kggxTPsHSFULm8mFja8e4v6PkdMeLXLeutgy738xHz5ceS4wgUrNrvRL7wbKI44NOUGIBF3NI
sbJ+bOCtTksHqxJF8JX3/G328rhbNmDGIiWFfXS+eTIRB03C9g1ed9cnamOXDPje6aV728vCZWUF
xYlEg4QXBW2rq96OPpt6jiid4Plz5nHQjjXYq92zTtA+9tZi8yzO7Gh+zbJzal5OyjLupLBL22ku
xvpL0ilNUJ7lOWUihOKd9BHZDgJU4QabPw6pbTaewwUB0BboincJczZAgAIMATv70aec1qnY+Ms8
oaqh1+bTxiAGPzOfY9ZE/HpGk6avUEzj9gg4moe4M+Cym9izxAKMMDW5874ANCqUZtLK6+7A+aV3
FhEHoY2r/UHYfyoF1a+9smxJK+vkKheRyfplI20WRkBoMbPQKAkF03Te8fzoCyU/voejsFTf6tqv
FiRCD+M+zbOP1mAOd7pGYl4cq96LPpYUGf6ecTm5ctB8CgC4Yu6XNy7c6UBnrE85hrDoRPPS5ker
d0P2HZlgIXOm/BFaMDw8gUP0qkSmMomvkMpF9faumiJtrNidxwhKcSRTkEa0iHBNkj9U90wepMpp
wun5DxIJ2xgvCkBWsoLy9on3uPH2yTjoDo9MMdh3B664N9O/yZ0uTn46ODQq77VvQfFVgzw/lyVe
dimTb5SMIFO3ZeFcKgPgxNodoQameDtg+8Ye6TPF53V4eyOZed8Yt7kVuzfFTaTX4ToorVoqG++Y
xjQkyWC5GMSzcXRJIKaI6ycyNrpkqR9QjA0bVu6jvRSkwZgTdwh++E0y2r47kly3aWOPn0FMiPGx
/YJpJbL4ePZ/VaBUMgOlEwOg6odF5exgiWsNPHH+Bdz5RE9YZxklS1ZIKAEyECkw5xGp3C2Awjp2
Km70+QKUj34tdGvfBQ2qIpAIBr4hhkrP14F135op6K07IuoEhmr7eDuLG1XIS7a0SYUQXnSbHuAa
4V7LyrI3vruU2kBYtjGxAYKsL/9mn1oB3sLdC/yym1LK8siGQDKjSzNJXK4QXJhvWofafj4c7iuh
ZJvIkYkkku/4ZBSiMKxQxrQ1CmoGYYWfQOl/oSGSYAbAQP1k32nmaP22l626W8DTlQ11M3KaYWoF
/qb6lGu41r/L9/sIdDEGOnIneong+tXI+NDkxW85aNa/fWphCYc8U0Rn/FmEauq/ai1u3g1WNDkL
B59LgE79sFoOamJppJH16sLTYRplCMDCaM6SyHgg9rTavcGB+H3woHtAuV4KKpEf4a5+dpmCBQna
RkuY5uvLE+7PmlF9xUL5D0TPuVMSKClMsikx8+eA59AaJeWo+qbw5UM/nHqj4ac5UrAPG80rP2Lv
9CO1J2jEUxUAet28fNydzzQ9YuGDklECoGy8/oGjUY70Fuy2IrEBi5K2+m3EcAmhoIocJoJP0X+z
yqZ2OwvNtd3KdXErVXSaT5M45BtEATFo7j2k7maIz4hxjhFCFewiWFQQmtOZ+oyEJ4NtD0Rxoys6
35Aroh1fmpt9CoKnYMeSUImOmVyshaWQRuS0eFGNxUHKiS3xipu59Rc5FXS4FoQa6LpeGlIxERbU
G2NJCnNL6JOVXPoQITn3dkYmx5zqeGW8mwlVYPvn34UPa12n8rg2PXN8aAFL1eeta4omuE7PRXeH
EBZ6hh9Jleuau2Z/S7Buv03hJMblbr+/Dzu+rv1XA/c2lVq03znrSAH6ojrtb6xXXse3iREqLEkW
TKJlQk7st11jLktlhp1NlLAkEQ/z46TP/c/LDHBflybwbuf5POhM+NknswWznfZBf2s75S7fXWBL
/EKEd4em9tnj7Ew23SWKoebdLhPvXqueQIxjD3DPjHdzH4h40hmz9yOJhTQNRVL5u9XmGVLlG7E2
rEhGZN5BakPems7iICyLo91ztDwzOig48boyd3nZmaSvRHT2EuhgTHvQ/Cpd974WmK4Ot1CcGT9t
HU2L95fqYxfhkH37uoN/qXqvefXunEGZZbRpaBufVcxsEL95O1nkDkQjzTXXIuke0zDAXGoAcio1
5Ej3otrhrsmgk3CrjqYHXYqsjZ0iB24W7uM3/gk/R8YE5LEDB1QIjwmXFts1i4r1LtTKIAdIn03K
irdUkcklxCeS3sXjhg6nflsWNY0mhGNKHDDSug/7hop6Ra7W9PAHswAWnNh11NvHbbdAyewFNS95
nsUO8p1ACXOPLuepGLR0/GscuzIeAHhrjvrT7zNiGGfQvq+ptTVRHeK6XDHe5givOf4umkwAcyPH
N++wdGqff4K4XjG4c1kOhbw80buMeAsIjbSJ3TrEcZxgraKzupi230nhW98io7UCanzfJFURULKL
MPgGtR7+PPOEQQN7wyNzQP9ersJzvY0rtyJvGEkl0Egfx7jae9N+HepPnZgfp6YnZ633cc1FpRY0
OYLTmBOgdUQ/zlFVY19y4Nb9QVXxEqtaL0WTK7yIEMj05QXpRSJR/8jpfKxkHiZmPWNYNo1c4Juh
vLIjCDGWLzFX3xdhfNpRleWlZx+JilETdBAGQMvE78nGCbN6CcfUaU3/eZsw2zhPqSNOn1xf1EU0
yJ5+aHxUPdn3a1S5MhaZatiXqZE3dxdiGLGCx0buhow/PfrvKrWxmD5XSF4+2qJuAKOeYVZGHL+2
0vyKA2OyUcELIeqDRNFgTspxWsNs0C/19ClFbDYOj0UNTfcRmrhAYgDBzFMkWvqVrdZCVeD+1mrc
5YDNEn/Q7pQfkilu3ZxdXZA/whFbBBNAnwrvmu4PAfE4MG6Qdc8imvAOzZGcsh7QTIXijJQ+Vzqp
597Fs+4yw1yhUWeNqwHbE8w1SrLwKoq9XcZq+/G2YexQ9Y3UDpaQEIBByDLJttIgAg6G6UZCGUcp
6WaKa059xP17SCP/ye/WiZTqaeIse9HRwk2jeUqHP+caAoqsk5fq4X/8IgFtI8mjhw0QwG5yAbMQ
q2sEXs6Xdbq1RicTEnXIF3TUqKwOVZX2/js5hDWC5pLWS7bYx5scHCeSwHDPJckmj6S/+z9iAuxp
IjB9ZJ9Nx5Sd6VGX6TS+Rmkahc76TIwXz4ZXXHLXW6zNFInfooQX4oHEylZsXT028mImDjPcoOnW
fkov087m20JdW4U4IAfEIF1cd9X+vyxg3uty/7dsoQJa3zU7aYMN4jpcsIB1EqJtNH7Feu6f0MRg
2rme7IknVPRbp1R+GjxeDGXtK7xWk6lSfrSf5R9+SKlutSU/0VwghjR6Qfr2aY2U9psCxKlAad2E
2NYv9kLrbgXGc0U6j5d0lU5wgjWPpmqDNEUBIA6EYQFrg9IpLl7olcBjnMHzzo83KtBpCa+/TPjL
uUelBHGle7je1n6YOgbJdt1pZGfvCyNOzoq/t45J4CjAC4G/gzank/K+n/StyV7sDAFnSnlGWNBh
ZtHVI9Q+QGGyYJljGctZBC5hDfujTVlZxyhskviUFY/MlkjsKEkLGFR8OKQwTqdaLi0HTsL+BvUi
gxSjw6zKetpkoRVbpz2bW4nKlpqdWObDBrAPAQ56z499Jgg0MQfx5M0cHJxHN/8NFS2olC17ouve
FxsKdpr5jhRnKWT2SqFON7Dg9/GJ4d50s7i2eDWEN7GwS7YoKJ5szKGhgzVBzE3Q+7BV9Q4MlPj0
hx0pm7ohqs6rRTl/z98cbvU2RKsgbJ7nXXDqlY6H1OxLheuR4JcAT6RgzJ5nsWarFaf9gfeZN0Q6
A5zaYSzLLvltLxMwl9JyJRWEkzLjW4PN73SUBKGG8F/WIJ7Bc4VSsGZ2yZfjcWm/7sMT7+Qj/WPO
xUZCo2h9DFUqKMi8zeD+QHo1TvECz/bUQ0YkXzAaRk8X1Kl9b5YdCeQX66xW1SJgqluXIeNsk6TT
OqaKIIQUHAPqGcjnpYBf1owlThwbtIXaha8FlgXa15CC95x1ooTsgw7q6SbSM3nQrH7AyXs5qv7T
iYl2TKnhdq6VUvYKi0/4mu008LqdK+RH37923AOS7y+n6HfPHvVUYIdcLtvwz9fqRFXOL6iwkvZk
2wANvnerBrUMQr7vYMI+1TckL7me4en3WbrHkVulFqyZdIvTpzyqTXE05h617S2Hwk2XEo1maKAV
/JCuBjmsDWUg2acvpkb8GYTgT99qATWPzUPwvKdqSznQtARwcTT4ApG1/MjMLCyIgnNZo6k5LKdk
WNsBze0xNc76ffaiEqBb++pkC9CM4hofGULSR3SGF7wcHkhrRyldjlY4n1ri4KU1+ZfSe1+c1nht
eV56KRkcXEhbVhhco5k5SKtXjmNb4udKgVdtF3GywQJun9MKfg0/MAFeLQtbAXgkYJSboBRwL7de
sWTU3G7REHutht0eikB4Ajmwf5K8qaPhJ3jTO8oL3Joki01mkkAzWKTq0Wk8qnZu8kk3BZTTAZlR
7YM1QqdsuqyT8ofKIUHRTqDIhociHIWOp06VMiUOoJ4pwizFncHW+yFcAKZ6rhURCpd0hSvK0dNo
kw60UO5uyG8LAes66H7WrJ2f+qFcJkwUrT0y8JRIGl2fboEzj20iBoXlJwaEguSpSOj7oiviRYaK
zS4+N1Hj7Fy8o0rPxt60ZyPgZesDMV3MG9fr0PLqE2VXyXn9ejzxcRxR6EdgiDscUj1lxLiAbZAV
PLLEVZRShnkWcCHZU9/xXmHjrhIZvbzt9SD41qaVpjKAo8AsRY3DkGWmEFQ7bIRZOjMAjwLUMG9G
gOkMQxGHwyVMPXJfokTnPsqcFHzUCUwIo4O+lqr8SeMRW5ZljEQ9jlqgTnEwcZemNQv5sA/U+3Rl
777tqOnFfDSiCJTrXOWX2UfX+rd3QEVl/4dPZ/PtQRINyZfSLI2GqR5W67SY7Lwen5HDGcqNquiU
AfLGKcbQ83k+47pxecWOJToRqVF0nv6sdy3QDUnp05ziW09zr21WXQsls81BADMhSYgAECBjAcgM
i5T4Y4vzyFNmSznJtRsYSYtbhLyb4rQ8urO5VmXQfo6MqSKSxuMEv5EmNKmPfyD8o4N2t9Zn3JIg
4M4H412LclQXgg3gjtqalG0YbU7eLtI6BJn4YdIQOWQitr9eqtqRf7WZCE/h63Q5vMkP48t9uEiS
+YA3uA55DC1r6ADk8hntvbwuVf1z398C9EchW9Ege2jwfO42QYcolrf6uXAQd2EHFAUSL3qMnyab
qrSaqILJOTHkLdeBZsCW0na6bBjx24iOJv2ZDiP+xwRwvpEhWXFgr7yp6bxWl1l7zl5sCpp2Iiqm
z9Yx2YDy8Vxx2wt9sPzu1RSjx7wHL+EHbeqVXUIwy9LeIFIL8fdSnHTJGrTnydr3HJl/E66reaow
uCJxV2Cg+xQBj88cnYthmjsIjTG1AbB7+dLxvejLnHNavAheY7epSXYVoL0pyT0D7uklF8H2LRTw
p2wlKrdVYe5mB4tTI06cikzCu0Wj8+uKppLuV9vRmE9w278ZX+SzG8wTz2TepUicRdkc2iZE54Ps
xFN2Dq9/uoQTxHmMdx5fIVQ5MrWqpoG1me230XthwCcLgMe0czcZZzjE/s7w4W24u7507wl78UBI
jTgKp4PrX5s4lXATKSbsLdg2Q0S5W2czrN+BQ8ChW60f5O/3IuRvuJD6k9mFpcms9ectbzO669+u
d2m+LUDOgH1lNaGvevqSSLewf/Bi1zaJ0aR53EZViZqaupq0awa9HBMDIZrZTKGqbTneYmBF9LS1
8f6Q1bQOWWcxC07jQUlrdJPVn6UchAVOizs/HTc2CBhSvY3SLPVTbakQFWsAmhNwz4lpVPbT/h7K
l/BKVDRYoJQd7wX53FCM8fRyLRRlF/3AuE5BE0RvIciaq1Czga1X4ChV+UIepMvbqi+9692m9aPq
CERWDX/2JznY6gwWO9cPC3iF5tKzUpxGgygeDF8jewRyjrm6PA2FqrOkrNQayOxoguoGc+eVZJ9r
yLUb/0bjQ5UTpwQbywy3PfX4kCQszVgDaS82uBWbBWzmyTWmfr6ryGca//+EbZgvh47bDRD1P5nu
adfEUm8qqjl76hNt3GpCcjY5/Cw6cTE7cqUvCp/ocKLl6pWCYIasXqv3ZI6jC8xVdXvqucFpDfBs
udMsjxQOqEzjDzZRHDkLbcqaJ+v4oaRMgMR0U3wBH3Is5GivYyhSo3fXkbN2xgJlFQSv6MjBwD1Y
iWJA9ZJPkSFAJvWrO/pAMFOyazvncwyR4ripUDuPJH0n0r1jqrrYykIZsDtNOQroh7VJ5l6lY7Y7
9jDNFdEU8ZQrQYTsHqtyeJu7zZVP9N3+VSl9hYOXDQpe54NJkuTYAE14j8Q78sD6jXqbofWRM2Vf
MCGJIfka5Okk5oyk0xGEHuD+92/X6jxjueFSTGS13sK87Pl3JltNJ3TJzKmmABfItGaA86vbgwDT
6x1Kt9TcEJIkB8e/27qh9yRkq+p714aYKMpat/DY+4weL4+3BZtVteeXlwIIecr3EH/32bTXKCbf
7UhAFePbbmNgW/7WaIrkJrEJQ7LDOrqgBQEsf6YdHi4JILFH1wWHPZ7iytUggXfZiPJGVHfPEx4S
FJkvscyl3fRJXHePaozPXZibm3CL+jDtQfmoay9P34TEpuW0Ozwo1R8dHWLfCA/7jqXm6ppUpz7T
+B5RSxmfyuk8r0uApmFw65AuLV8Q59MYLhPRX7xjs0WEWIdg13EYA43IBZJG/gNUszM7s92cmHcY
IOKTzd60N3wZxJMfhIOVWJMt8+k50nQa47BKXrSXUi9kA9CiKEMD25uvbxMQjoZFCK6+6Rpf/L5X
H0jd4NKPSnbmLLGacM9G9w3XX8NoMzDJzncgoOIE9UrR7Enb2S1PqD4A3/No62sBLk0d1Vf8lggT
QDydyKluygfnhHLulvmrPS9H56dGH5CRg4sP1xgQjyfvIS0r9/88FgeH+bYUtykCAb5017XDRVPg
JDsVvjDeYi1cRHVYm0tmQeKWR5+CX4aSUJVYw8HHuBEdMAONCsjAy5inTi381R2HJv0iXh8oJ4Ma
f63+mjnSippZpHS2db0ECjUKV76QAdyyTxzCctm++rXpsmX8g4TS8wOJbq09+Q5+nZg6XfHiVFH5
iQkH8ewwRGKMq73szXpEBy3rIQndHfck+U2WPQ5TY74w0fiAi5NcQW+Rah2yL16DwgKPJ0CI9Gr3
KS7Hn41LHkS1LcEfnaMA+sP5fvADoaMvUSuPAGvbfjtu5+XNJsPgr5qTZkx/uXMNmCi9A8Mme4wd
O9gm9Tc3ZVScevO+Kf2CICpS9hh2flImTXW5DLVQJMtZ5iWh6OFOoBsuGL9nNPKQK649xKe51aSA
Pf9qbiLpg0dpetq6/aEcoFzzI0DCfr5KEPYhyG4nEZ/4DRrKElhxvXhCgjj99dXBPShCpt1ksSV9
qLK8c97Ntrz+4MMrC+xe4zMNL4+y+CUfr5WBkcGN/xchWU8j7Z1J4yczjq0WtuYBFBr/DWjqhDJM
SfUZNnEOLOjTunJ3TYv09SjY1XAs3rgnEAj2Hi7Up3oGEfT+V4QFRUT//pRicEjp6bH+aPvgy7VY
xyI0UzEPI2BLuk8drkVSo/V9LGvYc2cZPTpBbLlp0B5d0ImntoKpQWEs1g33lRx7ohV2Jw7NV8aT
/d4j/Ma9+uB4F6xOwLkSyJudLhzdVSa6b5m3gvz0UXGgjhJXHr4WTahqOdBqZQjP/ILIDOn3kam3
vYmB/YRRZmgM95FsR22ixthQM+Ugr3N2DxX+kw+BEu3+4mgjmCympi1DFg+wHwWvoa2wC6qkPe8c
vFiH+vJeFMAmHP77h3czOkC0tErc6iCcAm3qNDMhQAYVd8v+A2FOHXk4pWeN3mz67olTWAUe3Mgc
HK3+nDdkmhk2aHi5+ZIHElaPZTQ24rNVxuzrjik9cOh4YRw9yYlhF+DjJHxunSlJ9N2LCQRulXQA
7iWlo/dTDHpxlcQ8jgipR6nR47qKj75jVZ2bmoWa5KbKioMCXcABjTotqms89z0doKulnVuKfosC
KEdAFSOmpp6wM4fPkKPe+7tbr1de5+65B40Rl90KWn//XPELL1RrZnmxpeGy6SBOr5jU57ylbDNc
K7pidboMkJZTQtwpgoR/kS3WA0GKkgA0hUlov2whq6vjrn/ILGKpVV60v7QeHpaWItAFp4mVdtTY
79uY9jVy+uob9aFQmKYI6PG0bGjQt+IlNQv8YpoyzEf1n0mSKv2upx8ah0hCg7a5KyJ8RXUWFns/
iad2UpiM7uHc84JnrA6AJmOoXkWpGOaW43L5Dl4Fml1bn/U7sHtECtZna70CsN3attBkiG5nVsxZ
BQHh7P6/eGHlfpchkfC7vL4pyGUjPq2zFBj1GdApCjOoOM3SKPbrUnUYcwIqIqHhKpR01Dl9oRic
AeqgsaAgSQnIQNReUuPbhXThDc7FCeX3PuWhf2ZOc2XHbB5/n5oHna67p2pILRLqz6R0T8TPfBDq
EveQ++qojvxXiMwXQag11U7b41z0SpHHyr26dM1DeUmzA0odmfdRKMD5oKrz976jm2rntVuuoTc8
LPGMjhtnfY30x8l2HKfmGDuqSsbCkyr4oXAEleMuij82q7dcz9zdYTwZSqRaecg1Wwb59UxEoYnP
ftLKfVaPyaUggUJyM8D7DUGOgDNUCuiXaIkMs3jiYcznAu8fjV6tsLVtUS6eGOH5wDBOU8dqKmbu
idKMlLMm7lgG9nO4JoTwCN7t29RRHdKkjtWfenXuEtRB2PxTPZTUZ6zs5lF9X0G8vsev0MMkPD0+
fI0nogJadtWJfr1JiHycIh9iaQr3Z10wr4eyGuHfekk0epDWyTS6pnp4untKsgfzx1XVg3GYpKZQ
oGT6ioFFK8YNQ5d6E+Upo3CKINm+An17fY+l/Ootx6l2XziJE7eGsbkkvDiP41NS5Hpx3FYzNGOY
uHnARp6SvIU/UnKblZoXRtAYNuBmVb4HhAhpDIPgwAzTavvLhHTnBoVxSRJ8gDvd3FQ3Vohj2GhS
hWiDJFbgjxCruB9Eq5DyHkxM2BmpVqzk0urjchn3aNXqA3Dfaj3FvHB05COx5JIA2NC5DjfAbv5F
jxOT8EHtyJU3UQbmzEPAqovfuoXDz5nfh775wDQkpJBCuYEx/7BgrqUvrIjZDRMc9oEB1rqBbksV
hjg9ouc+WF/CDDeuOVcPSBB4FpaCz+CTC4FyA40PUsivPpSqyVYmyCh6IODUXB3S8dPPviG78JV1
1SkFMvE0ilYQtVFXRtay8CSLZ1B1cgaln0ljN+s6bkfqdJQ7ygXdLJaPHvaLUcaEO+mIccJXiBNe
C0C6BMcRP0WNw6FJwN4Yur6Y9nhPelp5M4A/fhb96eEyTfy2CWRLgJfONCYS+4HbKGYvzmF4sh4e
/EDpIPkBpDIFgswsdOwSIoK88p7n328VCHuHqAA32hDppYYWyuFL2dRHN8eO34CzVF+/QYWk7k1G
Yf8UK1H+W1Adkxp6G96x/bvuaPopwvaquNDbeRpzlnAl/u/TxOkzxBMzLKbMaJdXolLbctK8s1a0
IQ79iJfnSZw/CQkcXwFbTTQurx8pG3tQZdf2IUSdK+s8jvAW+BOtSekJxSXkMUNID6d3v03f0bcJ
cRqICStMatZhdv1Ja8KDybTdUQs+NUuqlUS6JuU5gywZJwBt+VWd0ipF4ljw5aMGwghQDAJJB3iI
8nAjnrxj7I5rCFLXXLcyDntB/vUaEFvgpNVJhGqXCzayNOgKFP/kFl7hg8UvqxaUzYF3XxUu4g3X
6FGAsXbA0Rrh/i+DaLJnWYX/iJbdSAKGBbdd47K5luJxh0Jrlj4zrBe0fSZSDf00hg22vJpjXhra
FZ43PD/cMljAqCRZ0h53ZSd/Koh+T4kPBi5gFK7hSRl72tsdywBTicUr5HYNFpq9NmnKaQJWLnxd
/BLqL1ARKVVjhYgPhSz4AFA6/YDRYpBEJMVDGQD11skXvPbuf7YQpyR+g05pbPMEcTqc4cKkF9ak
vvhv+/dpZrQ1nvnB/DpPAa7pcf1pSnlXiC+fLX4trW7MYIhStuCxnDBhAR5V/7bgQWviDANHVGip
jIPUlTv7Zf45K8Z3narRAcTKqW25FqvqSPPBMSqotrrKGNho4q1if0v3mLw35ze0wQMtIY/kty14
BsQqt5OF/mEWAefGZvs5NOvzfAALN747PbgtMJoOv+xx5yjMWBiM+OTjkB2u3fjPC7K4EdWGqyXb
3ePnx7yVx6ErtdntSJfRM02yEtPKiRyQhmIRsHj761RG3R0YwArPi9FlHKeCh7Mr6vzmWbb0mjhv
41v9QhD3OjoUgwWIImgdoh5PjUbpGgWgkkAJLLa1FxG5sZPW9HE8sJ0ZCeg4Lix9CDyYJzyX70yo
GdUjWh9WH3vUmMGd6U7PPLPFEgVXPxUmS2iVKxnWy2+rfO+m3EQfiTlFatj4msGCIF+A9YbSNw2k
wIHAYUsjSkBa7AE81GRBQ9rq/AFjorcbv9Bs7kwDAtPRCGzvrsdFQav9ZvRnoliDGGcbgJCNmw2J
C67Poma2XINWYZeJv+M6JSOjDcXvT0TI7H3YUu9iGoYoh5a6xAXp1wNvaXqTqztjQBDhDAsA4d67
3tBhL41/hyzd+gZx1aRVcZpeX9Nqq8z0RihGOapAtHOL6R4z+HXgfZMxTg05MgdswcvoKmKqONd5
2BIs6ADDRy1AT2hZnMLTjsVJT4YtUYPLVUGCawwOQTyaSBRCEp5UST/y0cQzSf7cuuIRzzOnd4t+
/0GROGbwyWss+qXL9WIu9ZDl0j4UCoFVzDgkRN7PdCyxhY3MA5d47kavdxx7gH3dv56PZXF37Ibd
cq0g7mEsRUnT03OlTjPrXeN4GAi+NZEWg+NU+aQJDqKHYLAZFBVVNUNVTTNaQclajPN7oZG6SvJa
8F7paK3ACIXC7r49lZz+/qvrkn/EbAep+EIdoavW9b841RhG1Q6ZkumC1cWAFmHeaCcC6bfq1njo
ZWkbJo7WQTBPRcfEoaexstXUGQfu8NUlbMRdVx4n7AxEW3CY1qfZfNjCL2JzrZfybvbo41m2NbPd
symr1oFhOJrFPGp2u0kNNY+XtVG57mIm14kJclCuI5T7xuiAESHiqHyUlTA9qlWmRwhZpXUOELU2
yFlnMWdfuHtw31h0uNPMbYqmzWAWYKHgLe59/oRewalxKrNzt+GAYGmn2Gvjq1bVIpaRNITqlKZB
dnV7UWb0/wMs0f0QkaRklYTRVVWQenU1v5NU1Ccao7PjtkxWr0qI0JfLoj+xp1i/4dtiYlcCTlCE
atG5pmKS70Ct+T+2TyJr0+r6D/G4yORP/iUxTudyRbFLs8EqLwQMVkygedXj1mBhqrzEW4B+3fLI
DFYv+Kq0gJ6btHn0nBH273CH6msFujvvUDCAxyI9FBKeKgl3JEwEp0ZEcl7lwO/hLnyhvt6G9hXO
XzCCgte2zH95bV8PliFYmlsO3soqxCKew4MxLI12FESrvglEgNPQ/Mii+36oHxlwuS4fJFkgnb57
/qZF/9wTFOS6/Hx6BItPM25TdylGQnIAaa8CF2vkNp9xTfxkZDPLZhG7RolHoPdLo7HU7zRMEQEM
k+o4mzkwHhC/iN47rWV9RUeNfTxLqARyRUxbLapyDGA4e14kXgWgyb+16E+qWxwKdZfGTDFmzKpd
BFGgwUd9wwAa6gH/BysUlFXxr9dcnRIgHGv630g3IDj9a/TZfluC1s0h4L5PjyMXYYWlbNrsfReA
NBKdY4IpLFhS+evRXW4RQEpr6XHR1N+9BHFW7gNitz74dkR6YwDQd+XRDcYvc9DyS3IeTxMsNbcn
LQC/aSPZzv4m9QvdfWjraEoc1mGeezpa+EWKpNNqfEGw0wxXqNFyXnLYrw0jPj3DgKl/FWET0vmO
ZFwEXMm7h3fqYXoY1X9rKGV6g2z6wy1ld67AvnC8HsrweCR+8XFXu1JMseyMDxfJcpbFI2HTGNhI
S1/KxqK/Age9cspmxIKFvo+jCWsdKd1M0yI037DD1q/4s/yULhKN+Wnjvxxvp2gHFBa2eW2NA70W
zPWIbPkwee3vltRK3JzrLTuWwdLtGRqFPcHSUdjAwGiC0E8/Vc0J5XmSPZUlEZ9xweRDIgzCfjZS
GQV9ASBHsaJW8xCynCgVSf1NiTcCBZ8Lktmhbek01iKnQ2o93HnU8I5lUrFS0t2abr0Cpuq/BNzf
jXIsRSpXdp5c0XCI5+SJK2YrBOOeXYknviYnIvs9YYc5AcABEqnAdm5JbUw64Elkgs0HpnirrQE5
gMUiziAH7RUirtNo88QCfculLFz+EFCTGo5IFuq1Rb6rw3HzN1rHhOFW/kE4AHe09jNnW4CpwK5b
H/9EFQHvVAGG/iNSLajmg4vkGwXS+628F/80dczOgngpAT+WCKkqLFYe1R2E+r9Dde7mO7xSp+VQ
gDEkhTIDFW7nlomZ5XWx38s8C+isPuBRPzVWXy63DyDICYVRP6no2kfwy++3m0jEJBhMz5rBczXd
yN+3JnhwWXZDMjDu0Wq1l2PS+LirkzBDmVRMYlCjRftlkXW0UyGkz15Mwly4yLmVtN0F8xVoky4D
g23dGUFhYGjwcJrAXQFlV6EI5N/z+z2YfEiNNS+JbuAi3crsTxa8w5wwDx5gxcWTdHTyEGq5mQpH
ejkRZCoxvTPJLAxiJ7HDTUuOP46zDK1PF01X1nBoaaBC9iCN4pjD1V1qWGIE1v/gl/ILwsH3m26b
IZlCC8iKTCNfScDrJeyuJmkli43GWMSVBCFXVhUJwRf0j+UdJyFFl0F2fNgnOqaybB6GbW59covR
puApnij8Ti7QZddKbIaR0SwvnbPGP8M6FqSywjXxP6CzF+RTneVyWGIjMRCy7gEkOqfTvDtbIdN0
rjAwUNrkvV1Ee+ZPoJlvyOsSpOcmwxtTAxvAMZ7PM/3QtRYsBvzc1xuqg9sixUWizdEzJF+K2eog
rrtPsMAS3LHKq0xhXqw6uu5MH/QO3tLKwoLFDIADVBM0p2WzBuGj5J72vPRJMQta9X5rzyNTcAb1
K7CaTpbYcQqhIRhBRXQeW7qgs7d/Yv72lJgC9c4i/XN3vMEa7BGK8wmZk/dAkofTpdfJM3RExgpo
VcHNwBS/3/eJpjqO1X4C3pnvxMJBFI5Sd/vOsS5TZQSxQEkoYO7RExUzNoJPZBz5dogtb0TgvRCq
pgYjU9YVuUNp70lkY7P2WOzt3eeJj0F8GCMrR9ZaybPjAOz3cCYTvYKo1UTbN61VTUG/iyLKjNFd
LV5/Gf/+pBM95DfZf6sWSVWDOoWxvXk3MuF39goyh/CikAlWHATboO+F+Jtjw9gOmJ3CqjohgFMO
19iyTt45hRYaQv+QlakCuhPGQqH/+fJgwVUux+jZv8hOGYolbHGmbvDG5kOiWjYxnxR84ooNPPyF
gNWzYQ1ZJCLyrj8mzJmQrr7PqRdTdPZl3H1k6VdYHdQtz7B0valzz05e/TzdOjvm3CpZSIFArmoY
B17NuZymfE7+t+feIupZyEHjENLBe0Z5eL7FnHWNa6A2Mz2gNl/t/xTCZ+3pUVMTz5OW3X5Y1Zvz
Z6ehHPcKjJN4RjXNcUQk7FXuYNw+urLjpljMJJU/00YPnx0ABNnAj5a40pxT6pyu6gaHTCy18f7p
dy1LCKLleA7eGVTCYZYZc5vDx4W8NtWeQkBuJgBEZqyoQlku75N7Xhc5ezWGQspQLSfPjXMvbnRt
2V1LDmc1kZgXREgBGhW6m6yqsOXgrBQmMgdaBA2tuVpFdTH9pehjfs8RQA/ihZbLCClxDL9v/o01
eLa6oW2gr0conbmiG52Qs6vyqzUrg1Riv73nUwSUNkkCs9bdOPEt8t2KN7vDzzMrKtXiEVZ/XfLQ
r0+SGZlXd6PLPViAdZCwhUEIVT6/Phqe1c/BUIV+ga5YDGfQLmYYdZ3dj58ZSAgfqd0N+RaEPrBU
ThqO2Mxo+kjNFaqihub/srpfwmKHwRV0mMo1XHmWeXgVpAbQnQVzFMiWOwG2OMzX0h+lyvmSMR9/
KdtIVFidKCCbEckTdkKsqpWS8m4CCRgXeFUKZC/mX6Zv9ZlJPdkrNXIi1z+LrnI7zZy7EdMh4Dqj
MtQwMw4a0EbP7EucBUfhVWdmNxrFlKfOqge3shRV66RpFU2Kgmi4H2+/GYq88RtJudUpbVQnI5of
kXlbTy9eWbxNZwuw88w/CnDHUTQ2TtYSJoNv2Zd1yzUQhvdbz2aT4RH8qAOQttOlbYh23fuD9+eG
YCREQ35m3nya4w3Z1RX/qjStDotqd+fCGbdZ/MIr87iNFZrWjuzzuD9/3MP1eimSWURK094IS0Be
Sce3h8hrz9i3wX8CAfyAgILGhNd7Dwed6/ANAdOSuYX2G4tmjrDEcr7LaXdRU+8oBDkit7DK8IvN
v2pskMwtuNBmUWGgOgvvBz1g0F+IiifMEX+cB9cqPKaU8PZ42IvxAEpnSLmiQWzvUsyGbCaIz2cC
GiF4B/xPDbyetbmdzIyBOOqc4bEWVAxYBRmFeTPTg41shtvnh7WEmoYteyvbKG0vPskmqPPmy9R2
hWyZckF607pd8vHyCjhdB7vlEonEAXaD+pSZXsZlUPJgXV5MavF1wFW4nhRcDpubx4pe8wmdklE+
TH8Wr7VR8WcaFynOG8/IBT0Kze+XZ4wE53wPdboZK2jdYLWbo23YDle2Hlk7qqBbFaIiWLuTB8oi
ehj/OxEyAMn1GLiXXCEipJcGawpioG96IJBPoGQB0dQekvolnvaoxkvVRErtd1X0umbe6ea37O0q
dnwbWPI+aPBZflgI733zHvWwrog2ukvpVwLVs0WsaoyDGlJ+MGUnB6uaQNQ42d1UkJ28Y8sTUJCc
sB325+6YnkreCXxXQWGuVvsz5ORi+09XUrE6iGZsv1Sm59bN1TjzRGH3veKrsvioj7+T7Asz3BgD
GlyqumiIBwAA/NRqbvfxjzzSuQuzLTd2qCRjrNiD4qJjkclKBVTqpMeLlMw8NIp52oAVkFG6x7e/
z0duqH3+5aP9u/yQB9aOIY5WlqWQFW29U3HkDrcLnU+sJn/294yQrubXAXI5anyZOUVMxG9UHdFx
1YzeZ2uocRONEBlwgiaSGJ7MJ0ZRdq1gWI5ULCVwPsCbbUpezQlu9nAvR/SiPc+YPfejlj4BBXiB
aQscI4XiVRSGI9EbH8KSYZNudQIdyIfD4LGqGwtrc/n37G3UEecWz4dU3xU55qQW/icYA2qtnj9/
YHPaif8UAjTeA2Q+pnBvaPRpWPs8qXl7sEFB0OPEWNIqrQMYXSFSB7U3msFHo1dUH7Rlmpsc46SU
rCGvqiFtn14RqaxMEcBdMMfs2IJA5lw4wqLNIiLPM6zZIhhRIdty8+AbHI7gjZ8ECOcTXwcrc2+i
0+oc6yRcJiCGuhSBN3QaHHThKneDT77S1wucwXF8WpZWnSu/OF0Sm6RSpQjfVIh2uAhgzUBxfjAh
pj6m6YMSMLRwyaYbcdSQhvUVnstwsTp7wDGysA8R80eesv1qHBT+u+jUax4s2aX8ljYk+LIWyv7H
KePuGPOgnqBmq8xW5S7jb4EtEzdRffaPL8PknbVMzYhFUx8J1jsxty1hj7oR0r4404kvMTT5NiTW
8L4xDW3dut0BNE2ASsMhf29oC+wD09R304maaWz4ipSyVh3icYgMw8dFtQv7iNFqd7tXo3Umhbjx
1uaa8rpX1DYPiBgg4MtLkF2bn8uvkx1LdQsDqr0Yn9QVltAk/UchT0M+3+O2eh0O4E6+l7S8zs+c
IWen7ZJ0QehMuQN1cq0DDHRKA4fc7ITeeI4Qwj7becvmj4IhnC/AXBOa4zopXjPd85YGdS9qGtMa
8hURnPx32ZSrs8ffIqzUiRQMCBBcUikpsRpRdDoZ0SbHth15+WhgES42kK2SoLyK8Jc+zwJsq7+y
lmlu6QmAijnYWtQRbFZUW76DOUe/GWMlceB21fjIJnjDjSDekNcFrMp/K3QQTYmVkN7gcJai2Id/
17j2Mx27gN9ct7+4XfqnTBEx+JqCoyHC6zis/yr9plNV/sbi2rmZM2Eghiech0h1JolOCOmOIDPI
7B8VNYz3g/Dr/dJbso5OMaO3UWja/az5fgB/YKc6m5Cs4QgKRFxXQhPpFKckSJwlEvScinlhbOxF
d7aZzhmKOGA/TVgp96kI1EfWesEdPtcCdXMB42QZdO+v/SmaU/olNAhcQm3cMTFGDjuWereFsdpW
wz9YZByNAde2SVmrOB68iz6GIIt7FesTjqjjJgVH9M43gz8S24Lk8kFwCwHFZXBcmvRmqD9K6bUx
kc0mUkAaD6KQdCVtenZmpVj/Wfrh7RHX1DUWYqk/Sz+OjiaeL5/YIJErYxrVPYvDcVmPNrP/qYjz
cINvNxfgEfktRS+L7J6HXcBc4p+E5JiS7CvutRe30hyy9zoXPLEFWaSmKODHtF8REVJeJ1xShDY+
ZtPXN2LB1m42ashuYTprQ//E2XyADnYszjhW0qXdt5th9G05SH+YtazpBn4PU94t2CXYQbdNvpzA
NPpqMqSViySrOkHF2eJUd6rJhFYSq1kiF20pIvTSPyXmP8HLG5nOsXj3cdVTDkHMH17PQ/kcnVjB
eV4GlP0AQwvayXwtkAmGMZ0/fHISm8h8mhmPo2HHW3r3/sbLcYaSATlNdJmet4URM3nGelMzcM/5
ktUhSEEGtZRW8t6Q3C/XoXZl7u4gODG6uMpqMcli7fXN7Qa2Vlhwqqb0xh0rV8Lg2Y7z8/Iub7NU
4nILU3T9jefR7t7l8jH4SW7wNVSJl/4JiketlkzRwEAN0+mk+vn/WAvJPohFjuKt0DACRo+/l/tj
v3/JWFVGizuecpOewoP6kLAlf/H2JMOd97CkxnBgWc19qpYM28/nJEkQBQ36ScyyBgYtLh64Yjvf
ovCvL2+sna5q1iGLs2op2Ks+9zeyPBSkrQ7t3dc2t7vhW2/zADSiiWVEJvq6PjXhVJn1uS3bp/Jk
kBdcCOYoaCgYXB/VTWV/2l9n9GWspIyQR2zv5zLTeuawTekTj8iB5/CiT8TEmuvgEjdiasCTk9yp
bzqBAnICoJLTK/jrVU4kmXk285Njp9YFCPAoSOw2h8lLpdBZVGv06QzjkETPhPFLoJ+b1loERP3w
9qmK5iAaOhxOUQg5BjKyudLnlDyNAi2jv6E89So1CvcwFhRBW6y5fS/s6ietJ5Ulrd4Wd4Fo2QEq
EJCBDHfHomuaKjHXslQhWAPq1lNtQzcGUDxnRBwC36QUOxbVROy+16K8sCRx/+paNApUB5zCxQ+/
kEm/P+wPKw9Sb7A/9kQy1GBzTnRynXzomzu7eaR5CAXWQ+cLqfzCj0rqjX76h4gsu6c/11+Z8+yP
0jlLB1Yfut2TVnrNo5uXXhB8Z8lPvYZxPClZ1lAFUgciZEH8hUCVMalhV9cv+LBMoOoC0ZfK5h5j
HTe44K+gdBBvpmO/9FYm091WuIkbtuy8JWMNBAjfurWiH/dEmdtBN6rU8T4jZWNDZq7cBeP1yK0C
KW0Tr7zJch05W9z7tM5s6OhL9ut/fkaUEvSw69kjEWXO1iBjeFW4ileCWfaJHFC0sxfOp5qtzCuk
ZNREvtdrjeWe6Qs8xCyg7cZlptjEe8FM2CRt2ZH/uxfGbkhcB249agQmw0rMWPc2c6m/7pNHRFO3
fXh33RNyqermJUBsB0daEipcxdL3FMEsaGquDqKUy651+W6L3vzOwp4xdLzMc1BiIf0/Q4DHPwoW
fub78QAPgNLW+KdC3xO7iqlw2fC86HUkOGmsmkrjPm4VB/FmPFsGDB+NybkPXaJ2anyjGzCJ+YxD
gES7WVekScfBFIe/xwKj08wKFnjs6g18JvFX8ILrlQiARC35XGrgogQvZ2ZYSOM3lFLlCMxqm0a+
U7pbkywkwHHzBg1T/umpLGyYvWtTxm697uDLUFQRfOq39sc85todglbt0uGtzv654bFbxHTgqIvQ
ndjfs2796DkE35o86nJgM6Ap+OGhp4IlnrsZJ0zGG8dBSw/jNoLjEU0houYh9YqtjQjPm5OIyylW
spsmi/McqRGDR1PJn3kPRMM0xAr2atJR7sw26ciFs5e8Pq+0gn/qFVd0TLrZRTOapEuLYV+Kg6mQ
IqJq5stZ/Y3h+uhVz0AA11/KqtUE1nGVljU0VpiuyaVXer4KStNAd37Q9PdZ9d0DFn1tlCzbzcam
BStDtjkugUUhKw9NxK7WeAC2suLq2uVZcJhUv6Ek02FeO8bMnvPMPsQRb3qpdUMCCp96wjSNyp58
Fo1dT4ejr83016RSx1hPu5PoPDEClKb7QJoOzSICMZwp8sMl/DEPbzWwmlA66xPgIepF3rgFaPHT
8ouFrVRLcW8rWb6g+P2XvDscvfQc/kVHsp29OiOL4eF3M6BcCMiQsQcYrTEkLKzfWljJfRgCYLKV
mT2Yk6QxTytcgQXCHjwVVk1WA5vo5473ZGrTbZTu0VXWRN0sxqV0uuZCvZZKLoZQd2H5u9AOZvum
mokyiHs1vy3cQUR3TajZsJLALLFyoVY/arX04exyEZtGawU20XaBgtT3FYNphkWK4B4Cag5HxuBz
o8+Kg5fDbaiCbKpIDGR/RFVGP4CWdKrW1InqZ3Bn5U32V1+1Sp8aHvc0skbGu1UrDcdwTN5nrFOa
qRuRjTFrUFcP238SDqYTmq0bxsT4uzkQWUTvheb/jhu9qfJOL/uJbxh+iXnBhwNOX+ZWgJy49HEN
86GPB58kdSg435VzdLhjnzNUB/XfLyCJluBljwFTZdhCzhcLJcbBNxYXwS/Y76SRmdKpoCsaD6Jj
jQjUaTZwhlHhXQkVOEMtrJOkD8X60u9na8t2jWYtFDF8KUy/MSQ5B9wpoYJWuYZGx7GGOclF3txj
Q7RNlkc1vBc+karfkg8aYcDHwYQlY4oGG5Pae3vXQavz+OrmjrJllQTqQ9Jvo/+hBUnCBjq83RST
uR7nayYmqA7pz7+4iBXHn7F0Y9MXViVTeIbM07egYXMm4fKv+f71hiu1LQmIhbcCDXlhe93jqyzJ
oxG1zT/OVQo7b8F1Q48R8rNEMpt/2h0uCrw+lXDxVTT4q/AIaeYVWufRIc90QvpjUYElmtDDt9AV
7/yIkXOrRnKQ8m6vo5wIGNmq78VMYNq2HQxyRYBjtzrf1YUAX8VgqiTyA2uS/TenFNB04Jcn9miW
NiZw+wlCdjtnQljjOjxJ6xemF9ygMvth/bKU2MuY07MxWtN6qA+xnD3lIX9tXtU1GH4hrzdpDK9H
XnCuEHwDhLzDEQzZKH6nv1cTQxa9fjC71qk5SbaeCANPgi/AbWAqwUmkarab59ruA21dlhvs5os+
DRt5f6fFpgvD975Tja7PhXyV8OzDa5UJL8+5ZdS5C9VCRs6I7QdOTzM4X0avbDxa0UO71dCMR6Ha
ifDPLuon9H/aMiUw0rS1eAEAPFHCOLN0yRGaMV/NSOwGpac6kwmNBej21i0xQLtNE6O8ud865/Nt
oEmbtRskyfmwIdTtHQO/BhftTo1qLssErvAcHtRhrFcZMDQ5HDIg6wkL2wclkVP/GhfQb4EbJMew
eTUUJQh/YO61YcNcFn9jWZHIHtfcT/TKGInbaSoRbuBiZqK/qPQx69ejKV+4s57r2o6D5JqXNC9U
zUgi/u1kysUMD+3xy5/fW3jDZ1hyrMpyf5fBxG2jccQxwbW1XlTtHyinrQwazSQ2ARVYz2qUixIE
82DWh6HSOzwiuMyp9R76kvcrc+ZK3bv6kSBm9hRSZxH7jE2Ll+lwopFhfjjeJnCkvO83RMsGw9Js
nCjxJHPfkGHeD+V9MszQJ+zkBmFEjk5DloI55mzl1U4advlZq+8Mo8dj+lhdC4CPkYy4R9fZyQzL
AAOb1+3tspekgVilLb1GLv6FcF86+nZD3WJEMgyLIjxbtK52TcsFgd+CmT3cxW7+qgwVxFivYim0
FdQ7T0xES86Lj8c9v3bhnciDDyZDpUszxmNZb4Y+wV5FYs5abTIDFc9vdP1CMi9LH74NkqWcOGnM
w7SpNpDJSvOba2pKS9m/3yhnsnfFXHATLVze6p+KCzOydyESfDnF9TilOuWOVPkpQEE16QZeN6FX
uz9BaPMm0w7eWSVYaveGF9JVU8pTgtao4VG8ASXffdolqrflfiJK0r5MG7/32MfA9zJ/LA0t/V6A
lo+cJKHIM19ejg6wuJEsKZ9fYfopcMF65/VPpq4/Qflrrfz2TYrqTN98rZIePcS0tyNTj1KQEGqh
xyTnXzMu/s208wYEg54jHANSOodWOcvo0vVwuYXhRU8AWNj/+MU9f7iuiNwIUL3C2MqZlEL2HE++
V7asTtxqTfgYsb5pZN3YmpAPOIoIcgmGbj5S7A8DBgKDyS7xkuTwcC6c7pGzWO693yNI9TJZ3Cf5
j3utNzkQlcTkLu9lJbt9yUzFcfE6LtooulEg+enZ5gRuFBVdCvPoRWRt1+wfMTycmo8Sw1eyPhK8
5CmCIOLQN27se+IAul3c3C/DK6+w2jfs6BNKV4VpFQ1eHpW1CItbBXC2eQQZ8tgA6L4x4sak6onp
gWsqVpboGVy1Se66/SP+LkvxnqaOmTuVURRXJn1bKahMAm78F0rm87EprV0vcFTfY9NawjH5Ea5T
yrXpiyQO2hJw9bKYR5acqro4p57id/kGbBiislsFFRvMyocfZiIsvTUyVol1Art1r2mUpEfmQBuv
90QadGG1EoBSlvUcC2ajUkZsB5Ra8a/qMB4bWhFMdQBMQBQE7h0AhnVYOgY4exASXhMBx5pWmvIb
5VKfzsy/SYWT+z5rN1OuyoioA8AvDeZzmKY5nF1nWQyKUz2m1Bhs6hZEAMedMNMfLHbdua8Llzjv
244P9CCYCvxjRA7G7zDECHcHjndHMjXdz64PaTsAK+ie3hRIGSYKmrEm5SHSpEFIaDCrBL83hVEp
QmsKJP95aqqtZePPh3Q88UGk4P69dU5ajiMPFZnpKq2GAvKFVYevkXZlI5eeL0Tk/8tew3hcOq6w
55+5F+D3A0a07H3TUBzGO5t+EUOYqI60lVkVCO9A1meQ7FZieOTJPy+YakHrRJ5zX2w50wlFRdUA
ITHQXMtCQT4AoWXwb+CmWQhnXd9i8hpaWkWMV5J4nBtN2Qnc9c347qWhM1m2quhy7vQuDOJ+KtLO
CzpH0z4nnHZltPlOvz5TYffFr+N1ODb07OumrJOQ/nFAjSp10twK9Cn8ARc5Wie9ZsNglESiRKPe
8aT0WPeiddLDGL6HGvCfhWjPYaNDXzcvNh9kEI7Z/OFEtN3OwY0TvNZBQ9if+zQ6W7h/p7C7v8Vt
9tlppLOQoZV/qbbfm3RK7YKvDDIZIGvdnTiMU65coJo5ruYOIEBR7pYyR7x90WzwJEo+8Iui0ldh
pQYPAuvFNJy+K4vbk4YZ8J8ynbawuflQmymKmNGIz9lVfvzhr7fbCu0ileVYTJoes7bl9NPAOh0s
2ZOucaae+wkgCTVR4hNkrDyHZ4VF7T6nln972Akn8DObVSfXFny3NoA0tpY8xAQRabcLXeQLmZ78
LUreNobViyIYwaGLJ2IsKWuW+cxLbbz233qUaytoRu9Z3D0JR9EUzWYT1GogDFioW1CfnQGNps11
WF5B6KEuP6/fqnIjIS7Xfhsnc3Iyg01YWrhvTRZ+fcG1xqxdK0+H0VhONGK9GCKlhmJuKASGEf1B
iaKTOA+FRPusPYxtwyZeUE28UjJwcAbYrcaF8G5x/voSsxErE3tMhzBm/T3GAjQkEDRldlJvhhrR
4Y2LC4YaXTZapnoEqiccQbBu1ghnKawqLyUS5Xv/MLL9oL9uBFHWUSO9cB5pAM+9EiQNYMfwubSS
JbcdQnD+lE1fJ6YSGNb8SXbb8zRxDzcNM25zj6Qt5OTLLiw2W3daox3b+tKzukz0HzqKp50W7+Oz
aHjWQ5OYk3KMzaDlLBzOLtw25sCFE3p3mfzGhiRtddzz03WfiZm4BdpDinJrUhd9OaPhg0XvLoYR
AafPbqjjar7oFWR9xbmvtfAWqOvhOm8NOczgvVViTaid869jz+yKr8HD38fPItAYKjxUJsdvVqhh
3JakcFTsdXoDOvEGVal79hecQFwJi9O199l7RswxnTy9t2CpnpZOaFAsdxp8ZtSUP5Qw8vBRTrqa
qeAeZWWcRxMyukrGYHODTcKYn0kf+dMeZn12OvJ49K3NCoAHPzaIRV9B4o5ZwyWK26IFZgh6tw+C
ObZUrHRMtbXXMGfO/62ClrB7JWO5aXIcczVZqk/IpR/R7u9R6/OJUQ0yvz9nVer59IasiiFF7hK7
RF2OLFuNQpvHBXxB9eqS0tPyB/Ctvyxbj0j9OrN18KcyZhlK7OHJtJic+RRskjODjx9TZsuYCHxs
XSqRt2yVF6QvP3fEnPhORLr9qNjcEAPDmyWwhK+j3q+yRjYzMUoWAGJTNxViU5QHtWbYAmEbl85h
0qhAlAjewxwNwAV++mRA8szv5VLXA2B4CtDw+cjlxoShYNcW8xh6pHhDvsjiShdLzCquvyCppVeL
3CTlzm9WR/2e6v/qIk5BUKmsk1HrZsIUgHv/wcn058ODesRkDOVMjim0Ph9QJG3fNG4xdy5RFHE4
iOdpYrZv+CMXDJKQrT52nvcpLkWBB7sI/K5rR652qUdWHLvJZNfZ/2TnD+rRAcLX044t2qttm6dp
8jdod6B9wS/dNA/pzkngfdxk6xe75sf+7SFh/yLuQCrDkoToO+4KRgW/vdP/sGUbtfYeBGjUjbEL
5qiIy8r8NRKmxZdSfvTK+JlviDP+mdSpeVN5miN3TO9SAonjG5SEyKgvIo3fuftlQHB0RJiyKoyJ
4ENk30rpzpQs47go5Ou1QHI/8t9psql7wk8rNkjVwEoGTKhTxW60cdpugEtsC14TnznAn1y9MrB9
Mj3biDt6utAOfS7sC/yPBND2Py/Q9BHfxBE2XBTVD5B6k7nm/ET0k2AzeZCSnLLZ0RAggXblYA9W
hJYwCg+hWhAswHQesGfP80xNq8ZWc7pR9Kz14Ux1R25ckV7cp3Wnz0dYI7V4UZDgDpjYzGzlb9/v
hk6FhZj1HyOY3x3q0obG8blizUNV93rmzhmsBaSw0l/OOU4BClinfC/Z1lsNinYitqnosb1n4GT+
dPdlLfM3fy/r5Pvmys8e0R8yTfRoHAgGq0zjfk6mcpu0GeZx4bM2Ztrb0uDuQG75FmxwGhqg8tNV
/p8oiccwm0vZKyavlzAY5JVq1zwWWC2Y9n9g+7zW0n83Yhbm0f+ekvc1P0rxLtmhkp6Bq22ON559
KVmtlDtw+Pj1XrQxdHvKoL/HbWqViv3O9J3IdHQpjq111WsZx7sGslceZTsbg7m1EHIPF86pWKLd
VjqAk6Q4B2sPBqKVTu/CJjK+RUGNn5xRIvbwhk2NU/bRRSMl04W6PJzhRr9kNoHFd6S9d/0Gxjn0
grMsy5lZvFky7HHpEbQRhrhIHWNl2nqSyIivW+CSv5qh6hRFat+KDlEQa4vsQHtgngJO2XKbLCo8
z/M0zG3a2hen2JlDkBo9nVCzu9GZpXzOnQtwakOvI2D8HCtJLM0M2MV0jQt4q1U5z8kquqYD+h9I
a9+Pmwlg+DMVI4UwGpBJsadTD2KNG+oPhHKJywUHChmSVDWgFEfPwhpozZWZkcLJZJ1BibEwhDnF
8KtmO1dAQAlZCOblHwSTcfu0GHpFpEPfzW5pxSa/FZUjJCwlrHGoJlzrnThR2PJIZ5gTgG2CraxF
L+Ni4brL8F9o1t8K3dwl80h6B97ezMgPZnEycpxYQyzpJnFJe17Kp8ksNsBul0a7M7ALi8pTdngi
KQhNq6kLkAdw8hhfUOX65TV64GYVgbiey2skV4fR0JQQTWy3NIHCRlxtQbhItk45GKQN21D9uZer
44Br3To9JrK0cJdgX5tYBYl7lcg/xV8NWD2M9JF2onN/FPHZobw8rsNjEpnK5J766WLvyw5u5gL0
6ivmwLDOMtTPUArzTAczY5NAbGv5lAQ+5sMWx/xQbJSVAcsfF8pcZiFPbAg6ZxgIXdbvCUufuxKF
1XgsYcM5QLo7y115FwU8eJGzHrEZbn0S86TbClgi4G8x88rrLkE/M6h7nsRZ9ndg8r9qdqm5e07M
fUsF0KRdIOegkiD/j36+U2uVJlo9FDZ5OVq6dRvfqH0tzqOrC2cnzWT5u0UUyQSQLypXoBEACfbg
R5236WnbSXROlNJcoSiqzmGAzUjQ0hGZ2Qly+t8cUt7XWd9vltilKWh0HfFVXE+Haczmht8aWd5k
ZJk9GANrsQuE1ynoiDyXXKmHCQwwuFHC9K2VK19RbsGu/LoXz0qc3Ko95v3ja16t67Ai/42tdLNP
v45+ClVGMq32V2f1yiFXiqMnNIKXmYGq+Qyk5hN3wC0bqOkzC00gLtm5P5xmZMq/JT8N61EutTip
4rcm7kKwoj3MqCan0X9bGfOQFaAQyuGxNdcMOUmF++pV8np2tRPZmJ0pQPNpZ7y/L/sd8JkRUXyb
Ag5caQil83pq8H6MLGhdKmFcA63StH74+dKGLnatJKaQCzJjS1Vk8BRl6wRTinrq02FG/bO0VqJO
Mny+X4Yd+wG3sxi3LXP1aZ+IWquda12hP3iEwFzL1iLrbkbw6fUfv2S68lVSHgYn3McYNVN++WqI
7ezBxgU/uS3VE6qD9YVpuuXGFwTYCE6+RAx8+/OandwdRD3rVegUmFPIShW8jibQvU2JHkHKilpG
SCn4A1aoKP7dQmtOyGui1OpRAGViXopTiUriLHoTIPIT+nYzuFQySFSgXcQQ2qqFI3FjPmpA1mTa
F9G1k/7xjaulAvQ6s6QT+SbpNWH7s9HQrDSKkXnrOOY/nrtE0E7GKM3+VeQgq7osuQ6Fo0bjZmIU
fedbhfg8z0snEqftT6s9spmbkpyx/Tfo/QGNQfW0rpUPY2NLmNHxPlliVNcZfn/6JB5nHoLZfo8y
sby421Y29KsSNVQcbzAlXxVpd8EUYHOlW86zLwcDHeOzha3XeA7VA1y42yEfSoZv05ooM1/PESYg
WJYWY2wymOpHpvXkozCojSSZulXrxDhI8M0qy6grs3cbgmpTHkYlAQuG3a6tOo91unGuEJGzOSkw
t+WzroAY1Kolb9rOF+YecYoHYgMVn48et3ptXwv/Le657/HVOtV9Hayk78sOqmCaN0azoS3nyETi
QZaI1XQvTY7zOPDl+xPJg9W9droH3g5h2LxOD/lF+34AZfZ114jd+upG7Ne9vr2yPqK6wlwyhm/O
LQU3QnmZDxzjCVhYVs/jemQzZrQ5mpInsOiwJR/8sj5tGac2WduDquWPSOVvg9I+pVnaCHwpsnrN
79XPkTDccA8AJCtMeGBLFXP436ALsqWBm2eJMQFtS9Eq9PMS7iIRC1eKXNuc9rZD6xZuuARKApnF
8JTnKFCnv0h1jeSHN7FXtFAVAlJyrQjWvlepp2n8VxVuKOPaw+nb/4aJACTZhVlIs+86fuDH39zk
XHsaZuZgR4eLGUFL9DhhCOH+GRUDjOi8KwiBVgFhINl6qCCyiGwus9F57Dnfw4cRZq0ml+cwGhj5
sugbwGmMbwSZ/S/JRQVTSXZ7UclxsEK7++3j5kwnvNZ+sUUSCZQ9Ogb+DtD6jC8ZY5sHwdcHY69c
TFa8IFqEfJEjN8pUDSATKgq8RltA3bC81l1lAd3EJTrhX5Sm0blPextIDN7HgtH+dANZVd8VksfH
MfjtI6YRr/mYuGSPOmGZ8eanFLxsQ8rkTnAur2/h+OINZunjdBEF1YYsvqhp831Cy60B1TX5/kAB
mZXtnGLNgxNtu1CBX5CCb7VrCAgCAovmk+NXVLVH0gVS9OXQMRENn+4J5rpmMn4Z0rQO3nxOqKfr
dAQsmohvEIEtyxUQvFcDqSlIwgqdNzjWILskgkaIxML8K6rTcEPqNJwvT+zNxuN+wuieq3Yr6W4J
zuEjywJmvhWjD+elxp2Ft3GYLJqKEeE+QkQQyxpJLoDD1VreM7B/XA2jxquJku8+J42RUQT1iLMo
w0wVzMjWrbnJATQObBeXMrekvYLPu1rFKDBcCJjrzCm5BThPEtqx+YnhNfWVqwPvr8DQpOILKsLg
xfjRXxZjP4MK4fl9mEBcUTeoUXbwTKFlFg9H0PLugfZ8X14uBpZrnOjLbQFLQ4Go2PLwzcqhuO+a
GrDS2c0OZcOTR2iz7R/WHuNwNF716oRx+FAXw04OVqxeWYan54NQ5lFK43CzZEGfODB8FxLdOGGc
MvF/XcJfy6jip31uQ6yh4tc7wJXksmZJqAoTGT4SFrAYYZC2AyTcRgDu69LPMMRmz4zis4mq1jkG
d1DBEO8qHBlJEFawEHt0Y/Z9SIFE/CiHFhUktcVibgrO5fTm1Kp7f//n37CBqjHwsqLcy6JSzDpd
AYTSliBy3LJjDhK8/LOICorqXam5kBapICwcMKzNaKTiIaCnKyG2qJPx1F2Bgxx7MB7cErfHgsej
jTE23J3v9JVarU/n7NwNokqFIRNd3FnNeNpD0ABzLgB8y/6NiWjtXPpZzfQJl1uzEAY/RrKCtDhq
9KAGyrDr7wUlSif0xsFHDXS1ScnkektHB+8L5b5rOKgorAHU3wG8vfbvxZ+COjdRTeD5Xrz1Yj5U
XKcrCpDiM9I/047PEoMcvvlKzx2ulN1DqmCQyLZCkQljeehPRlZsRgF0WPLfR3E3QLFx6kUTNAfo
IGIufE1Y5gYHUcBCfZiEZg83YHy7sIHGyfpvU+hYS9cP9cq5+haT0/krejS83xEu8vFOnmtWK3Bn
/cxSIOtkEOpvFooloQsGxa11U32Ryy/wZfnfOJPuUVbmYGSr6TdkGkwIisXBNSytkfj3xtuONayq
7jcLORa7Sw7ybHXRKblKJw/x9UKqhLV0FWop1KVw2MDdK5kYekgRKcgC9HrP/E9S2hu44mjwoTJB
pussgiSQdnOWZquK6nkb2MaVOPPiPmzfPzpfGEIw4Iwr3Fg1Pq9kSdSgMS1r8jhqzq9Uvj7YFNTt
fW+Yvha9DRMCmJF2BZwAlrPzgxAeeHX+1jmasLTKT/YtQM2riEs8TeHxzFE+pVezHvK7XTG1REv2
EofIj05XkgP+xXGxG68f2WXxkoWKwvXo4X4JQqn00ea5AOmIm5H1D/eGEAZtXiEoDR8sl0hgxrTf
q7Y6lETTQhclx1rrhXB096b/8WlVMy0aOR4W26AFspz3rxi5Ot+WOATcjgOUzDF31n9sPyJyej65
e1i6HmBSFedqqa1ZcWNfsWPiBHOY+SIBdrhxbgd1ZYF1eKY4++7Pw0RwOQaGd56tpLLOgExPmnaX
SteXETqpICrY1xpl0v9TKw2Ud/GRcCWtTeqZ0qFXhng+VKST0ZcmfcKlG+3QbuJ3z/XFYGdL8f2f
zK9QfI2nqSlS4AycfFx/F2GWDvk30xKSShnHleBPjh+9ppQyRx/PfMbiLA4EgjbTqcM7b2OxG9rt
B0ZUrLmXySlEJ4Y4BCxcAI66T2Fz3CD3NUI9vCsILME9Pw4i1foQxOPojAYF+zxcRnkpUtyoZdPq
c6X9/7Na/ba5NYgQvSs0NeKLAhew7G/UurS6BdEhHdj5yk11q1xzfMbAUMK6F2YofbTHABhTVvBj
Aj4WrbXWAgQspom24n/aSBB3skbRa2MuddEm2n3bpqkazyMJR0mc6qM+3zExhiuCyvsTouDvrn34
xadXT1VqLEmoWPsVEknfj4ClZm9ekdiYupD+Sp0Ow+S3vc7a3My1WfKkhn7LgKrZTJaJpLzw57RA
KZLaiPJmPuDZtDIbibzvKq71JOKxWHfWyBeN9lOCv4OLq/hPjI578odwepWpUtViM4W4MJuyA9/1
42g6G69wEbQVo0KL224bsZOmGH/IojOj00LSE3WK5NOnjEOZ25iSULEoEOFbZf4v+Utg8+VI+OP9
qEAHonITZBCQb5IqGPyeN3CydfX5KgpBbw0C1A1gM1cC/GXaYF5Vbn9u3+WxTE5aZvYeifqaLcvF
cKYbIt1nbydNie6e3AYD79OgWSm8aqnBBZLw1j6R9OP1YWpgckwOvtKY68aaLhGbq1JdNqC1ovYw
flWvIqEdkj1CRcDUX4oPZu/1qjFGh/mAMwxIv7eDrYVU2ASR5IHmXsyEBeBKMm0YvoxOLTI3CVXD
BSj1r8vpZ3j/XT8p3chvaRbSzhJyye1J5YnAcF+fRGGPPpHKeDU3MxafubCKEg9gIUKfnICwcDaN
56tH3UAI99rdQ6M8iySW4iIDfLasP89bywXHA5kGGG8hvn6suJx41HGtl03XxXPGJ6zEyAAlAsHX
1XgEgG3UEkCVHOxC6lEJTr1VQaNa4v78fpMWaJ5JaI/NjHjyVHd0no7+aPMaseD/WzMTzrNCojUc
7g4x/t+XtvMF0bj91mEbI4HBDTFxRdLyNhf1/L3mE+kxyeDrFo+NohTR/57e7nPoEoFkH16Jrk5a
fBkumHSB6lCsovNMlQXVmb72vkLHchwvmjt8avfgHvhEV+eJ3wWlc3hQ7hYCP8/ZvOnoofSFbHIU
rI8pWD22coO5UIEd92PIqGF5hRAAY11DQOB2NzjnDX7+iaepcAwMIJ9YiJ2XJ+a41yEOTNsNhs2v
m8d7k9cP9ZYUvfGJgGoCihWGDZqTl9raXVohsHC2Du/SJ1X4oiOrfYJOYaz5wKHzzeJGclXvXyjd
ooQsWN75gMF55THiDvFh8Lv7bvD3SwOovr1rpHBnXzebmaUl/9iX39sKgvCpM+AbnVdTiVfhVLxo
DMl4vKj6u+qEZI53DO297mIWtuhlKWe+z+MkWQiyVZEgz7BpSF0WCYWzUbEL/6JVug3GLCkhwRPc
lm0gqFU8/hacd6S51Mve6Cm8x97+Q9gWBMuK42CWSfx/bTlAdK8R/tiRIT0o98hCbRbX52DFQTqh
Txgh/wXJY556ExwxuW+cmt0wEmgZTWwZfp/cn5ZhTdnHHyL2VRkqt0dEPC1CriknxORE11mptH89
cPTKCwcXcpfUqVItbaIKf0db+vl5BuRX+/xhfoCDkJtOZUHpGb6KT/6FZX6BnE2cWkqewhNThu47
UuPWe4lki7f60RolFo03XPdubEHZITUQk6nXHjJbv5hQGbyTBBy+dNv7p4pMSUsu0aMMhXPo9Di1
KwZmtxkBJxH0WNQsOXYet/enFq7g/stwRliScN9FI23q/x+cTPfKlioE/1g00TWM1yfGlZvY3bLS
3v8N8oIKE0STgAHDQcbMuW5kTADWocMa+0CJFCsaWVqn9ZZugvZ8H0Fp737E3TowFL9GfygmoFTF
LRj20JPqHHqNCr50M4naHPIDJ8sXVq2bmJcOex68zloNLRazF963fkXYV1tPQXTpFqzr18xykWXd
Ljv3DRd8Be39YiVS6WDUt8k00Ceib8QshT9FaPZ+iJjT43MKcpk/lbXRo/DPWLabZ946fbcUW1Nw
mGPokCxExME3I7WV6VvMzFBGaJs1RvbnpBzdIUk1jmeNvQ+oQgAGHcHiNI1topp6oVoi7Nf5hj3V
HS2/YzE+W/hC/Bv+cGM0e+2hOQdzJ0PZcOCVRerj++Oomr+kCn49PCHi0kGLmmnfNdJ2uZuGF5Ac
CHpd/NnPmyR2kXl/7iVD72qAQzK9RJXVYmojR5Zg8PQ5wc4N07nmUU5jqQxXREVmlFuvxI4sS1Kb
kMzwoGMhdwlBYQVMb/XYS1uFYkHexWhnOe2dV27uupFLCXSScIKICwJsajqT+rvag6qG93CD3z/7
LXqjYEbNpskYJpd20TuXZZt/FDXLwqVcrPzNcQhehSA+qGgAIAHHsX5uJ5JTPyf3Gk0A4YF7Xz9T
V3bFP+FYLllA7JXRp7/wK6MnqmtkQiDynbGzfNApnIvjxPDq+12iFIlANQ7nG3n0lLVVvw6b5CqR
3c7d/A5U1fjeqGSjTgc+LPogLKwTWwcUOs2aUas1rXUNBHkXj6J3b2Ylk9xqyKjYhAUFTILi+BXt
ijnnmea8qGWnG/gfXd/4308j5VBdrLO6+yAJsCNujm++0cNSJpjBd+cnMOwkG3lyIzk6LeVwDDSj
HA//iivcVJBx9v1/N2lG3cnFyjFaIVFOGHooKmqtd+gQJasrrFxWpOMlj7MaENUaDZZ9vlA4st5p
bmfS9FyGoz/FiYdz2BCNTu85DZft5MI0VcrmBDXaynieuC945poy5SXimwiaff81jGWAGge4HOQg
HAC+zmNXrKR+fod4s8mfwusi5Hy8fyMHvMEbmuiwD71xhN/SA7pyZz2C4SwBcUNZkFw0UefCf+o9
IffqLFp30eln75DKxxnVuHZ4MKwKYdx9IPYkXPY96LZus4SqAu+IJjyykLffBDuT/O+FEQVydexN
AEBo8lIOf/8ctuOo/+rWXvfhRZCzlL36vG0sk9tEfKypVmz8rAAKCxeUScRGnKZW4BWJ8mnCtpx/
cQB4+mnaL1PjQGPhaWrrk8i/l5Gu0utkfdq2A0gTKryGzyehPu9JPFAEyF75ZxMiRQ4wJ7l26OF7
uNxncaFzNe0LMOFD0n31AUJw0VFPDzDadVLsVFxhKt5Y3G5Menx10CALV+QWP8p/o6n8khGcUpe/
/lfefgpieDegy0mOA38UAFI9ggDGiZdjGMF0n+9oclGnsw9hGohvxCaN0fi1JN5wuY3He9mxQtMe
lhHcvuT4ZmSkweJvOYrsE8wCXpRjW4pqxwCS04TBvLlJ+Jkpn9NUI016PRbaW/GinucUJww1e8qO
fG0hxMEayY/aw3cID/Q4jmJKBMSUpOuXdb7/1oUwYnWbejp2uOsXw3EOImzYMr/XJ4OL0GikyoXU
dF/cA61NLiqUDrtCBPNDJ+AD4SmBVr0mzJIjZc6PRJC/G7/OobkdPsDtc//60hmntctzV0HeZ3wk
WEUZweGieRY32+dBqsQ65HGMyfUj4GGw7CAystWUlouCLskkqOv1yMbLWtQoqPKHnaGHn2d7767E
rEBethM5yci5krBTqKb7EIkW+XG0vM76p7b+xTuQUyFZ20vNQJ22/0jw+8RfU0irUX3sBEmaBY/e
YkVrv8xm06WqgB6Fd1fjZoEfWueiRmDeoSFoEnH88z0IvwAVTXRjXKcmJOZ/2IE0ncg2sOy/VWz+
pHltIlqgGdN+E04NazJilOAe27Mo/BIQGOwGg34YQ1zNDSCBKSrDCXwTNxwps98jUetNshA40+1g
LA84xup7cJoqZ4Gpt4gnaySiR7R3DHwIiGj772dJ9YqqROCZhZbIAw60ZnXoAXSJyagoqaNESbaT
lz0Y2dsV4B6uZDK9ZX5tfpHx0IScMun1znIemTnDG1MBKazylOj0syaJ3awON09oi+VkvVKGRbIS
U1atXKDxs8Y3xpO5YsnCmzsjf0uvk5V2S0e6iGCfZ+bWlNFoZ+M9ckEpTZA9C34iWRHlfs6GXA/b
W4n5QVuTNe0mgivXO9HM6Rcka1Qp1zDkf/K8tk5uHy6lTf56QrEw4AE2N/MibExeyKyx/8wt/jKP
iyjEK+s1X7pRmZ+U0PtTOK6a2+uymmygZlyCm9YzjRNYa7T0gZubcCleqcDPWLombBLXZPqrEPA/
f7WT4Lrhy85pEtoTn0B338BLuQnYNqsROaLiSDijbxF0X3S3aVik6JoFJJn3fJ+GK+S3miHgOEYJ
KxkJZmk1hvjNB6DdpinFY77X+G2C/A5SmCUEcNVjicJ580+DvTLbHT+DDY6odag43kh4wGGXCRcq
V9XlEE4CF5GH+9NdrB3WsA2O3h+xHOgAvkZEQWw6Q5FgmGXKRR4myI+STu6wK90gff9PYZLfInSd
jqcMZ846xjGuJV57xqJ8NFoid+g1koWKX7h2WeHeVcWoYv//UEm+1aGgBQgnfikDcVimoiwRCJz0
JlCO1puHCf78B8FbG8L9D5L2bnhxERbWQj+MIQ1H+FiWhQxz4XJB+k/qVWBZ0tyQCCpDFz2YGU5i
egV0dJvyJJyBjoUXzT4xN5BnmGrDEMM52H+7YasHZvWXipaTbUJcgTZ0cIJ6mwV3vZRFt0J1Fjri
8ijStaqVDyPldh3eQwNz/1vV3GQ2TVlr6ertMdXmx8x0q3Ib7sQL7xdBnL+0dy687nDFfUs/B3O8
VbJoeWGg0Xppw76u8WfjqD/gAu/vuaEZqYuCrCrB1ti3nD5BPz463paimGI7mE94jGMZMutzl7gl
10KCFqqo2ebaBICat8NVYZXJMO0++E237PZEemn/C2qJe1ybNODA4IU07zMUJTItPlDmYmipp+H0
KoeLwgHQVAHipBVK8MGnbDGXS/QgtFYOaCkabGcD3H0jjDHjvoKx1LXa63rasb1bkois94kxkZfx
PiBg3ODM4qv8i+n/v4mOZlFVgfntuQLy7t0+ozOTJMKkiLjWKFWLxpE+8FU7hEqtDyy4dOcafTiM
DYaVxBETahfUC7sXZWPfDTGFM0uXZnixt13ffyjQgjpbuxd5ufgDE/YLVRZVE5xJodVKjSP3y9Ho
iwYMzZQNJ/BuayDpFhrkNfoOcAvn97rgsI2Ph7uggEQiKE5rlFJ3zDuNsJffhyiuSqtwVpImYYT2
WXsrZ1NMYzm2jweLXi9CSdKmiHLzE8gkzGZyCIj8Pcp5JiPBDeohrc7eGAi0ifdnQ/xTCWJNNtF9
hhCGMg4PdUrh9c+swbgFzUBoat2Azty7WRmE/dxLuyn1K/q8kVd5NsxkaNRYtZxfhKWvXHASBr8z
DbRhEyJ11ZATTst2D/mTccOxg6DXDjnUodUHfbtXDDX1mpqn+IPyf3Iy4DbTPuyq5RO8gdocLdkI
uMg3edyiUA5YKMm0MjfqK5y4BuwuJOf+fxUyHUYi3/6RcYJAailhTIZZ663rLypA4LhOynWFFDY9
bjMYnqSUCpOxkkN/MabUKxv0SMZE5UP8Nf6FxbTJgKbYLGLvtzYk1Nfh5QpMrTfbwg8ZoHMd7IfD
D4QOQHWz2XwiS7eDgEJOl1g+AdUJf5DWBzJsuzIWMyqzU7mE8CDdghWa6dSLLONozUir01HlY4kx
UrCidG0HtBbb++DxaU8niK+0bB3YoTiY8qAIdplIb07J66zCpMYcrPdpswVEzI+IYBLExBSxaAey
8TCquXZ0U/eoFAea5HEdHnWe+St4eiki38dSgZ1xnzFkac+iBAT6hiI3lu594hwUj307laLKOvb1
dybnnNKeB0Jm4e3iMLg9pmNgm9+Nu2Iz/NlxRSqH/MOoG2p7zJbDo/jO+uPrxrq7eqUrycug0ru+
f0PMJM3MuucauBRtKyzLQU+A/nVBnsU1NsafDeO9sErozInF3MGknm0pUnJrdmKztAflnXXpOJcU
SfBICgq/ovvBlU4I3Lt8Aeq3Uz8DMpb/8Z9j1CLwVp9nYUVEwevBzWYiR30TrWpT2qqS4535AGAy
PIroebovY4Ju3Ac4nmN+2tgkkW0v4I5+STmDYuPvjurWCAhxgGbAXocMi4VTf/ZIcmtxmJj0FXfn
G/XR3yQJeL4EaTbl0Dm2ZoN+i0nD5oVeDi3QMecrrySjd1f40ePrTrXtkJYzkO5HYRckswWssspE
gEQxRtQbj34nYRSYI1XY92V2AY5AuRIvEHd/bNSEe2j1phDVKfv5KuIoOD7tknmxGxXGeMA7slR1
Yyi1xSHN3HzY8XlOvPgusUzbbgUr0yswDOJ/Q5vM59WbaMuEZWasM+4vp5uMJPxcoYNT8D08BBZR
/yv+8NAncV6kfrdvoV8q+VdCEHKeoGfYHZv4iXTP7jVHC7LJb+OEUgRooaAdeNhbNg/jUJ52cA+R
paOeZjLs1ataW0m7IR1BMhvzZGPURISnjn6uuAWE5sXbvzzw/yntpt1faw73RDQrvlwM8EUA1jUJ
9Qyze9rlBriU973qAlUD9fIFuIKAUi6e3SYNfb7k5n7yiueTUUJAqyExbYyM2PBzzOU5nuIQKn8S
ztKEpcEcenuCzkTqeq/ZIRxDP/F8G7wpypq1AIWxfoTL5GiIVnP062J9/4RcHxdszr0CDmuJPIcB
2kHuamyDNK6/5Vur9d+BOUd09dQI0TkwHM1ysBNPeJ8repKlZLrO88nA+roNMZQ5y6VcXAcPHTGY
wTrE3p7sWBT3U9rR9gEMZsycEmYFT5FzAO9wb1mUJovyDUFXrtR7SsEKyRUY5VZHr7YMwdBdQP12
v/Y30+LZm5n/TaxSq7iv9X6WUVOY7VcqBzTmgwSnH4zlpkKB9TJoj9iQlKsgU3zjiuCVYrlDombM
i2hp3HLk4dvM4BL5NMJpbCFKG9e6zPU6t0asu0USEE5REeqzPXieE3lZzOzd0btIsXQoZbcYiiHL
xaCzLr5LqjBS3yNYlLHl6DlGwDxxsDfoJjS77UM1iHBA5tDxvqhoz6GinHQkNB41LpXgQUq+2aKh
YW5i9vC0iKLav0H7gu42kDoTsIIuYojqtbLZdukEdZeK9GWD0sTNV0CfyfN3DVDH7watJSHsohu4
h7RTmYzpdgFfwbjJMdIiCedXr8RaNc/9rJZYG3xE5O+MzCrjTAlZArgBimbjZiDnvXNR636x6Hhb
61h1f6gnGGrxRLY91d4Sa7kwdozrI8AxmYNMZfOz78zGPYOdUxPfhiWaKHvduYCLZa6F2iT1o6gy
yoNUpt6dfSXoajyQPYglOeGCIc3AmtCfcIXbqXGwE57jr44Pn7ELE/YlQYig8CTYZAC66NKIrffk
brgZL0DGivvWCUSiMsViDWKWiV/5xKrU9RR+ruR0gjD1DsN8pH7G9pfxpgsWGAHsb5bKLqJmhSip
Wn2XIchvv8BjzovrhyodZ3Cck3nVyrnKizJZFBO8uSoJZQ0Mk5/eE0xwexqEr74BN7O/ufNqEdHR
fajvbn9DJHt6urTjEuW04cEIpMPKWJNILN/6u3dayMaq+t5sfzcrl1pVhrvFS9C5TjwkMEM9zGcW
+C4cRdkqAnkcXfTcIbozX6LPfkgV3fixC4U9cN4J/ecX+g7CO8CzCRf2zxoG21sb/t4e5bz8ZKji
COBnrHhWvtLd1h7GTHjk7ObxYMgjp8zGu//RHsB2RVpINASxgrc2vDxXytbDgKv0HZzQuB3LTnjt
khrDzZWOIArA026qk53cfhcBd4zzKmcKOrgzlsR1ORFutrbg1F44dXbwFfcanUgJN6rWKjWyY/tn
nKXKCoSWWqKJ/nQDE9Lpx56jl7sw/Cr9s3t67/mO54PnXJSFtPVUeSSSlYkNpMCXZnxpNt01Qs1x
HTdgdym/b+Z1flc1zSsTHuYnoZ+e7pLeW5rsl2WAphywwqGO4pyCnf4KX1fN+vPdfirtAIPo5gms
i9jzW+5WFQS1HvY4u5lz5jqV2irkoHWBDY+QGeJ6cO68DTCgTqMHYqunTph7Z8raTNbEIQJnij7V
58mfmxTqv/7cmV1FTVnWX6bKczYPbRV5UtLkT4ULM0NJAvR42nPWXan1vSjteRC6qKDOL3E3bAvX
FkYwPpf5oaRWQMFevxZ/+JF0DdTNuA3z4CDTnDkJPiZTv5iqolpY4YFxnMnWnzLVQbX6ElJQZIu2
daWlrMygDts7GKPBmyHst4ikGs5N4fjO/XXKzpeukKAIH3AjrQnJPideE7F5M8iEk21ArxSNqXcU
jfCNy3ps9MxHd/h3tfhAjUCzY0pdZcc/s4fvrxlEds3kRuhiQCfbKBV3KR3y2I1ftHoPIg4A0HO1
s21zmrUDBUNBf/LcuduPqZXBdaOzxFzETre2eyI8OADsAvwq+B672lkgBHIZ6QzaihrgfLUbqHCe
6Cc/xCffROYpjEXrimPvZhJ9jmrqWREhGmegWSfehadVsQEwhm2N9nsfgIChUZNywM+Vxjew/+jB
H6ep+KXakmloxIXyKV7v+I23Zha0uWFqZBXFPvyWFObooRL2hJkRj5NsrGUlLekh5HZFhT/Bw+oG
pdx9wIHlCNKkcy5EA6uxQveLDfaQ5o2aJExYvj4QKMascGQxij+9POVerNi0D0ETsMqBDXAlyhsL
GeZqhIy/2FHrMLtMVCVYBl/BZbuIL7RWulCRGBY7l20jeqC16bx0tthxoldhBDEqFJcOMsyyJHc6
m/jsKe0kmoHMxT7MCkgb+8gFP2GnsbfYwh+TzEAgQna8Q/6iXoGziTih9gEAE4yMlqIFAAZhlhcj
f7QWtcB/eQae27Uz8pnRMddqgecv0+nJkCkQq6K4CkQ+15V0XvCe0NcxHi89rc+vY9npT44o3p5y
RGzlbVZffHERX5B7S5KfCeENMdj5pHKQNZzNFGNKwwGAxsCMmBHFm5fCfggCioIQSn8TYorr1aun
U9X5Vgy8A5EvTMyvo5h6G70Cg21i2anVyXqsl+iuGoEG2PBOb9khN/s/fOYzTCxBL/e273jZ2TE0
anSv12OE4ifaAOtxCsLHyefb0YIhSvtdgPBe4oCLVfk7RoCeeWInlb0IoK2eTOUHuehzFPD+/vMc
/B4wiwgrUAIdadaXdk3f8Lep80Yv39KoHGCeOziiJSrWJJ6DYKPwXMMGbO9eBR7ed8UFM1yFdKYH
RC8GST7XhJBNhzQAB0BtPoPcQC/5uTSusaUw1cXLRKOx9umcsVTIXmAKJAf3mZdSLywgW3unwnP8
6atwxP3OJMEeYnnQXogQqRmTTtbmcuYrhUDb49OlPErF+RprYNinFVcjVdBqKVe9hoI/KKaafh82
VUukmB09RLUTmyT79MJ+vFn9spDHbb4Strx54fbn413AyDy0hpK14fvMQsYzJEkQv0OPVA7lZZmM
AxXddh6kyDYAL660SvLKhymQ50sjyzV6Kj4ibQiBd/BoqKorQi7DhKQp0jAaTdCvkhe6XRS4vvN3
9Jbtnr8MykGH7937blwJsaTH4fWzF1VRMRhY5vcB8CZBOF8oBMSNurKpqVhNKYXPPChWgGcCKqYR
UZme+RGMmTTro8ImkCR6vBzsnWOg2Uy8iU/t6Jo/yQO/WqwTa+1AubiyXVhKRx3vuto0nSnn8IQD
SrTgWJzFkXZlJdvd5N42M1o6E/eZzcRj6ZJM0C8jmbT7SplVtUKEoplngOd2r+Z3k4zmELa5mDBJ
YOEzSyQiynwWHcUrXt4LpfoCUoFZyRFaOhqMe14AoGPglYGQKN4EIwbmBXGgycKNYO2w1p5c6pX+
3fKQ5I6Z6xhYlcl+FRn1TgKEPgmz5uzMlVKfz/CHyzw/8OXcwRXdspQ2kMyKVeNAj9sGGNmZTw/+
0Gg4rk7uoIQ4h7D+e1iQEJjLQycDETlaQWmziBpfqO1CyFEsO2NbVClLVuJRGZSNRo3OK8O0IkkP
OtTUuHerM/YL2xtQJaks+0+NjYOgHq6XT5SAqpofmGIzA42T5htE7PyJlCYyPXc77C2vNvNKOp6/
1Ep3IKJ/Q9vsTEUE1FDN/49BLmjLsHJWBxFIuaBMCmmYOJzd1KBs1Go1JSrad6Qxon9gzE5RLpMC
YKWtnW19m4y8axJ7Be2wCM7yzSNsH6ffq6e5aaKBKEWhxMEa4NhvWMjfIHYazjNGmwIAVnlXUvnG
LV1PDjyOBoAJd/OJmUv975NFfg0QEmUga72KWeZKpjk4g+4vvCEZKcKLKRSGdUNX9EOPNGxeTxCQ
qqNpYu+iS8OKRPNtNovRxkyDiJZItxCus0ZemTIAETHwGikUnJUfkGcvIK8M68C2BZ08dAgbBsQc
K07bJDt6OLYr0VZDEcDHHN6+I4tPPSPNupTL/ean7QwnB7ixVDvS+0pNfW4j0/io19sl7FrlwHUV
uz1Lp0ddl5hAlveKObXNgkh1PUzeHJNiv93OJuDIR+4OTH0JcBRU7cnGfog+hPFNR4UOrNSK8l1T
VmVn1P04fOQViTOKEkkS3dx264aExPWbvsndKOPznssoN8AaKdROkEUXssF3afpnK3V1Fl/3r4dd
fzZHpCYXT9RlpMy6k50f0OCQLUTK3ccjNX/ke8rK5CRIRR8VdEzoiJ8YvuBvmS0ji1jXPHolnWhf
GrO4PT2P0unNVnGbxMcOm5hy9up4HNupAjhrVr5GafOwXa+HhoudNR/ACkpoMUI7OcW95A2jqIm4
yVtyCtrgOOzyQfNd10F1a2lpj29FRr8Wmiw61YKkYeuDbZMFSjUItvMyTRZZZp6I/bddtAJ4Ko9g
XFN47OU1uM8zogl1xYhu8qTjqwQtVNBcQKnxx9DZnyTcDkL7nRsrq7MByB3ygOKAZpluc4zahSNX
UsIEa8/e0gn9NN1Y6jg4I/JiVvfAot/PTb+kqEfo+KqMyUmOmBskSIQ6evz64eSrieFfvGYlTJZf
ULSM85/193KaKjcydaqKS/7xOWRLhRc90YwaOYp4cx/DNO1fFU4whEnh28hOyd0DgEJEZ1aZ3egb
fxyyEedo2x4V0+4akdd6sdB+DpbieVxwA30Jxpkk4/vAKwHCcqqn7mTBdm4zashByY/TvmN1FCnS
g+rCRAn9OP4DxUBVQAIy3TdpXY3ZKTXjYw0Mwclur9FOKnbC13iOxOhdSligXUQg5Z+lvtevPq14
BR7CHcLsdRBzN9MSXk9yk7nCvfL3+i14HQJW1O9+uoV/XPa+XQoRcaq8FA208oSPrTtmue1Ial7v
MdSn2IiBTt1pLO4512KD4lgboJfes7QRtYU27jS1F4rR4btj09/GOvZ6GFt67/y247JWYx5MubAC
8vHn2qnZMJ38yNkG70Wj9b8tV48x8VupeiYFnP70mBFzDxVa+QvbzebtLahfmaJQUL1e0kQpHWr0
aV2bKbWysRx9NFrw62J2vRE/Zw+HVjxTDKRk0XdVtuo8+JUhySXgXY/VrygBHieqa4p2aonHXGeS
SyKkdzI09I6o2fqJJ+3zz0fK5vrS/brrCcWiPX1jsj3VYs87WcDtna1AvBXaP7eTDTDJMeaHN/UU
/sZdGz521ZQ3JH1tECSZKLRGA0OOv6fBqBKzM9i01yx6TavAQ3QNKhF+lUvb9D1Wvl/eCUuHLM2O
j1UtPGKQAwOR/ihCO4BNddwxjn0MzJPdn00TLQ8PXqGegcFk+ixH5XMQ/uRrufqQCnCN2S1jAXyf
jQvs813gFoMi+ONgT6C5ayLDgE8SyRhDwSV41NU1w/+zMAIdFCUDn2tAQk/p4CfV8ehXs/RQx7gc
oCSqnldFRSF/dAYkcUNLWjcm/sWOL5fC7Aoh43Xk2cn76MsukbexvyoF5w72qQl4ssTzkoE88c8L
7YinPUhKtIo8B+JSir0WKTOh7mqhaM/fDWiJv3CSbD/kbpa+5vXnekRzwbxynaHlsp23+5kIdLa3
YsYXy9kp3i1UaayYW0+CFt4t6P7H61IC4J8UPo2Bmy2+KumTuTFV5oTCZ9lsSpVjk7irWVqYQt4v
ZpoBG+6g62ZaS29af0cqE2FrDDwqUeTKJNcW0eixUI411PKJjLZdhSmw2ECG6LMMnXeuVj+UKoKl
0eZ1PxGjAq7TiNxCzY6b9bJjXPMyvugF+Onv3nQtqJASq5OvavSyQcnB7d4ZddfLLxWshvHrBXDz
Q9V2y5HUbEQYqX8iIcfbHkI5pDyEN3LbJBUEMaTiE99Hg8H6nrgAwRnDmqY40e++UYznSXG+pHzx
C7CGFAMOvkCyRR0sVLwHhfJlf7UK6q7FpUwmgesMW72/yoov+BU/w8/xtEkNLdo5SddiTSRgfKVH
yykS73rImeyOTZNkKrkq6diirCnFPi9xZqaaPFhep0jn29bwRdZNHd8FsXeJ9oIFT/a4oh62j9GG
qTf6bweKs9Sfu8gEv1StlsRPR+WHSVcvsI1XwY2dCStxM3AS0S6ieRfe2rrX2gN37/8bvz+dW1PW
p4Er65ZqMczqf+pnpbSwDRoPozFxccRhNvGdj1qi0Rj+mF7Ewt2G0NUy905ingV+mW554E9PP07R
hDz2ijvP2ZjnSfa6IgoIwurwzDsBtkUobBbEOKJhH6VNExqbbfGQjRb04IcC3FmaAay02C8OKD/1
aOilAWTtFm4tO3RCyGKMDerZVdzEzWrEkpkazgYVIxb6Xr6nQjG0fuzCQE7lGnEFWsM1OedVq1FI
4mkUu0NCMSUnx7QepCPMk5FwX/m5sP0C5nsj+4j/qejmelrpddhXx5CjOuR2QQzhP70q3bEN59hn
O8Qfpr/1XZl5StxfIuu2G6ZxtWL3JhZ2sP424V75QpU4vPAYnFQL9CThPp17NJW0+J9nCff4EIQr
WN5+F/4ozNPL6iUMSCtErBYrR75XEbaB8u4JtXKoFI0nf6kU8NP6mXOrau0XN91kkzjSYXEQwXnW
lG+0D47SaQcaIAsqxMWiYRF2eqTOaEaM5HHgONdSG2jLAn03nyZBALQsrYeJa3MMdbvREr5de0gG
KTDQPuAe+rWlGoXXoME5hO6dj5dGb9Ac56RXfV33rq2LXfFIAOnzYYuY7pUdTAjun9D/1MVLE41/
/X+L9mxBNaeTcGUubDorR7V/qcP+doZjqEiCgManEe+reASW1h2n0ZExMLZqmQSbYgCKdKNI1w6Q
KEz3X6GSfz6L3KxxAKmjD44xWAVUR6v5y1XlrE+9kckdUwcOJA0Kz8bbyqLkobDCajH4umg+L85+
NZohaFcZxXIxYYq2ACavvfAztUKu3HIwnKb14blpwDnKPjjqC0qmYNgMFvlFg/PzXxy03ZdvIbFM
9ByytiI2cQfEr/sSuIebITSUgqiTOvWp1O7JZTAI2js/bj4yhJnsruGKqvV20UwmBXfb4+3RNBwh
Z+qnGhEiVjMx/0/Gu0sQKheG7ZELFBz5uK8OLmdlQU4lJQGhoEED+v61JyShr/s6dA02u0xKfvk9
gAlyb4+Y/Vr3hvkNt5oLI+TMWlZFymdX6P15vpMCZR0aSrDFYkZpy7LUFN7uvO5LvssNvDtQ6sh8
RChpaxKCznR/QLu3JGR8VleAJ9Xvy1EPqRZdu+XcfH+HjqZ+sKRpFi+46bMcCkoWpPvkfjkEvizS
DutV9Nk0mPqLIt8iI6y2iWmMMHraelLbbvHA3nEhCRuRNBxTrKG/paCNWb5apsg+4ESJMOKMfnYL
hAZWLEDrvckZqvDKQ4s2KdmfMROyvtEAmE2NHsaqPJYZnw9Td4CafbMhtcRMdFS44abeeGC9Ncpo
OiN0JuzCID+Ajtpb/QrX56TNsmU0C1O4w99HRkjJ5d3bOQ7yFlZ78Y3cH7HMax1AqWwSAO9cxd01
yXAdaElhQJOAzqRSiyEVfdXnfQrT7iMJ7U2Sk9LkwnBCgPTf0wsFfCDUA5Xs0DMfGHCKEOYC70nf
TjHQ98+JUE7K8hiiAAwX1y0vVDXBc/un/ln+QG/JY9cxmcdCeLZ4sW2oMx/mSj9eBBh8NopCYrU+
JJBlOSgcCeRl5st4mPNnNA1RowK8Hf+WdCDlmj1wFK7fJB5CKnXp6Rlpfxwd/8+GUj8z2Y59nBEW
fY/GxwF9i1sJ4ufPxHrlmv/V6+C9OnewzJrFgaOdl10OmRHDjuuiNs8Q9cnlXvGumOPXWmk3WwLT
hbHrqWvv5PUJBbECosS9HGXYdTE6OGQrH/e3bbimu5gc1rs7tS3eWi7DdGyREcp11RZFwSVbk0vD
mCTABLfo3oaaRmbsptAUHXogPvr1VMhkofptWOfNJXCV183Mh/52wc0itRVr/7Z7hv6jnFlPQPga
N7xHwbBP3ox322xZbfkQjPuFxXo+EXNESTJ4Bkm5IEaxS37JYwuzoBTBbNJKj82AT9QNoV+013lL
J7jSKVShVyAAvqPcYb8i2Sk27ARPvhvqGVtSONizDK6+JqbaWUmQLJHJfFuJ7p/nJ5Yn7tmV//me
Viktmr1KyeZQrRS+qSiLRTytWqPRLHDG0eJ7vSa0uIoGhnz/sP7AV+j4owRB86KGG7reZOqdO21t
fgkYygBWiAO+875XyM/GxCku3Y0OBzuJAn+YqWyitnxRrEsRrJS3hS44DV7Lh5IjMVg9Drl4ZxeO
AslH8386bVrOZ3pgE3vlBCjxDqZGHhOPHL/qHlsNa7vq1Q7ohn09HKkaP7VcgU+iWeuQ9NrIiY2T
a5Q79+/CdPOAotqPFMKL4O4insaS863CkjogQBWHCoGIwIQOE7de8ECD1QRF1SOPSba/iOwwL+v/
Ad8hukxP48iJbPD967JmOQS8Ac9jTufEbRfl4jkc2AhyePaZVnqsjON64MqPfMZaANfBw+iB+4Vj
kHNl7/CnVRQ2ECGFzfuzTrECi1PVr7keOKOoKtwcm1iLsWV5yrJRnBjvDtLthtwbFA2ffb8dOuIj
sNic/+4kfyVt546vq3Se13QsdUNHPL6U4TkCeP60r1hVHrNu5j7I7Ib3UXTo11XesBBboXqLsFAD
ThGDCnft6RwKTNwk/nEKLmER5iPm5zE/d0alPBV+UMauGLKfUB7m0BP/895muA4BKWNKXE5St9Qu
Wt7CqapzfNOqqm7yel4qPYxC0n720XzW85Y7Adiy9aNiB5XImvgIdvxkfL7DLAu0XW6FYF+K3QgT
DdxxkG7qfZMKpVkk/fJZjvZevncC8wLQ4y5J9u004d3Rl2llgaSR6q8WlNcVVdK0KRjfOFmEYA3D
yoRswNBp4dVMLZcHybCAEOsZGG5xSl87NfpqwTjwbu7jW1DGbjGaaLvXLiaqZ2Kie34G2pcZS1tn
HOlyXk4I0C7YTccdMij7nXfcG9GBsEoY1YRRyZABCMteh2T+M/oXdsNTkCZ9ehoj1vNxnmsHVCNC
aoHKyWsWzlGQr1Rd6dkmoVODLMNkPR+AZ5gPK8paSCFF0cc+IvOZ/V0SOhzAdi0XNgJGXmjHUubH
3Rx+kWbBV5NenXoY2qRA0YSbeb63JyrjQqOgAOyoOoN2oB/0agCToI1RNDteK/zU7O2wjfKB9Kny
TGSNqvraeQ9TGTTHWlvro353GWq8pt0A/ObC4bJiAN2vuhyOVhc6N09etFAfFwDz6iqgOcsrAxce
VfMp9/gGRY8MQfDgIwQ2kKIID3Imwyi4ozH/SwxmWkW9g+FQY2EGKx6UE3TuleGwslWNHa6gisEy
s33GoC+7xSpdsXCmZsyAY06nhnssy0wJaruG0TNHALB6W8oNgaZDrtIgh1yhAhSRuzZHJ0wwKiaJ
NKTiYCaZg5xfS9y8MOm+wuqEER8ub1IxRy6A7ATXba1dIJ7HSwQJiXubUXLSYyYltgnANh6xOaSf
7RRuoewtC3kOCxVCjYbnHu9iwznjjsUniQiZ6muux5zbdT2om/FBxQI/8x7CKEKIuAupz8v9S7Uy
4gQ92Sb7pnmKfsBpZc8thb0+DZSE640rc9yjs69NDvBx3lV2/8RAAsvmNSVfN2oP2Ul1cTiEq5HT
PSNK3VMh8y6CWlFS5rNKJpwUd6NO95LNN4/FbG54rYP4CRv/VHrw57+BqHxDBYrwhynz0vExWhI1
nqkz6MsBo51eAGGm4mCpDQpTsZ1qG1OAS//PA7DDEY+TELitC4kIQgkNL77mGrvQVxVjvM8J8lBh
lK8XwtzWaNSc6Vr6yDDC+5R7zwqP6eZKshfRbbABJq64FACIbvqxlsW5wkmKR3+BhWqDFLxesdBl
8tBDAb6R9XDCekAWqtO/1pQsE039nLa/TlrC8L7KlSOD5GUzICGC7lj/NLsAxjk35lk3Qm7PaMVy
Gj19F4JlPZsAQz7p7j7TTlJkc50DlAIbhHHY0QMR3SG2jTWVjsZhvnZEq+Gqy/1sKRLeDR+jPAYY
0UrOvuDWKs2eatkOqemDsIb9LSxHMDEnAww5GwblxETyUKe58lTWjI/gCF25fQy78JDVizYZKML+
TOYay4w055Scee2bsqpYC7APXsf4UPtuz76EpYQ+FIwodvcw/3nWlJtC/j8+zkmTrJH4+EklgI1B
QtD6CWssRb/d4ZsJgpAhvJvnn9IYM/rg6lqcJYw/o293a6AC3zyzFXoUKfA05XIWp4H4FG6SrJjW
hCEMTyqCgKSQfgz8ZuWBLS7+Zm6jXyj1UDtEvJcHvaO1aySfDfDMBjhLrPG0h5uOZBo9y20kKsxa
Afa1GC55nxUVvGgI0L0vEj28UbUDdlSNWgfNcUVo4flGvgGFeEpPkUA5lQYaW92xqtX7ETtJdI9P
pqJ3FGXCXpSaV20GijuqmtJe5tLJmAfwgwqqTHViMq9ZGqOoZh+ZcYSSH8DValKZJEjA5oZxSi3r
lFLbQ/8tjxvALlDeqgGFUVD6wp7aueL95TvN8avKbinUa51WaL76tdpxps7syjMpiN4+i+ybs60Z
ocv9ASbITDfPrn0wbwtjJX2q3k/W8X3BZajS45R/h9XL9kvpI/hrdRBwh4nLey3glxDnVLG0IxT3
S1dys0Y0G+ovYt1uKCp5vF4aYm5jd8JQltP9Bhc0b64cMJiybc7YYjxyBMyZKvaWXOP7z/dCJ7j7
+kNDHYDi7e+LoNDQD/Mf3N68l4gvbOn6z2YXxqMVufllNeqHhjQXlTEDO5rVXod1LS36hAHHDrd6
yaxJ2wSbfP+p18J4zlac7tsZJxmM/t6JoGxEtuT2+8MXuCwPPhnVDxyOnNB5Bz1K0iCcfW6G1vqq
CavXteqt3BInx9il/AXgoXI6Fte7skCxYQ2P1aEmN01dcZG8MP1uK6JO8V6O4G1AP0t6SbyNIGKU
youA9yJW5o7FXBSKI+rS5Ui1qTy67dwSpE3ZSLVTbKIDUq2LxOxsaZs9kQ+gZ/GBhRkyX40c6ZnM
H5G1OjEP1m8FUB2CVBQy+JQrAIreZmnX4UqDPJQkhyMVZdOOZTZG3RhgySr2At7o0/u48QJSTesx
U9iGnTI5E4SFx7026G5KunD2anX9Dsj8VvlrtjptDCHL+N6SMskbwJH6ZVmCpTLAFcx3PNHWJMKT
GudPek4zXZO/7cma/uyGySa3TvPB2rTbxHi3TI3M86txDZx+/eYl/6208Q1EUHLyTwQwq9JwJBlR
SDyfJ65Gw0CNaq6/L1yksxScL1tpiqSy0NU2wk/eRQ6zWMHMPCQ/Uc8TjjumZ58DeDyhM9Oo9DPY
7GfV5HEa6qXB3ks5X8myVpnxhuOgo3nZ0OZE49vd2fRU3aQZYr9/P/Y4cE1WjPxSrLMNB3LMNc5O
NM97n/iXRewwpP5yWeafnEtmxUU3MdzQNvBO55/sZqHsxQTz2KsbOhAgjZ8dsLZHKfl9aCAvC9XP
FcGoxVAvEBvkwt31gAdyuJxlrt2IQOzaC5UJ1VMHSyTqnOmPAMil2AQhbE6SU7rmwmxhxsRT/pzD
ROZu9vCV9OC3kmOrakpmcMuD5P+Klvxa9BeWZBXeNlV/2xyjuMEe3vFS8JlhjwO69gY/GprjNyjs
AqeEan+ZIxnUWUzXB63VMHt4iBbmaVbae0njKzYH1l94MzjkGzJsgD+CwyRJmBziMVb2SNZDWEfK
phRIebTlD7sQ3Cfs723VdtMHQgbWhnYA4OO5hBn/CLdcBqWTbvIBfOGGFu5cmwBGejuj2aIUmR5a
qyfTev1ASdcSWLhpSH06Vb234u6kX9riPAcLUoXBQox7qdSqr6NRaoT1U2V1jizCrrrmprA2OInq
tlxILP/FBcu2cZMkTd96H8lFsXNjZaRtfcdVXg4Or/X+PFO8eLdySCcCd9Util28HSADDLaC5aeJ
jROiexU+KSDYFBxMXJw9qtLY0FMExKraAnqtmHFIJhUmbOzneIdBBua4q7xweW6x1qW7TRi6X4iq
Z94YdeU0BYdzBRsxo6tUHQyoUBfUcZXQ2fZ+qyCKlTfEfdBQs0h32+dt1mppkOAOXgMphuPDHL8m
bdxWz0ljLEO979u8huuDxAHOa6obCgwCGCcV50h8zgIx75B9xT44JKSzhbsZvu1tiWKHvcqgyMeN
BNKhYCawZEHcw4vzclEg2GWhhYc7CSnK571e65P/S7Yyf8F5ecQHp5Qoi+lZknXZ3GML7m4bYbxJ
0YwQCH6DcAR4+m2bamu+Xe6IgBrN/O0K9EwKL5y4rTUhUqHIjiwtJZW41n6hZPGbtv+sIXUKWZ2U
bcvZwAVVBhiJc4vL4Ok+hfDzqOQNYpdKeISWex4KD2XmkKAzy4qR+/wp0/PfkTFrozQiIXJIx+Gg
gysqhebb7oBwf/lSDLrZVT5C+IiDUZWg7drrjOgIsjavD6RkQLmfu4L5lgoX6jKksrjNJ015gtHi
RLJJyY+xsML3n4JqzAJmAsI27YEH9TeHIo4aDdEOmYUlF3S4DbsJjwbju2diQV2MwugbNqvSVW6f
vgFrBNehHZXW+3xz+L1Z9GJjvQ4kBcLmMxDc6UtcJswkYPUtkVJ+iQhA4laKbZwfAZybHqMX/JLY
s2dukRzhocqySS1bRriwMApqEOonPwu64xt6Tm6hIS1ATm3gKFdHMzKbZakNlWLY2VZlLYqPTe7v
ubvQrEsYW19T1Bne4MR3X201s0rQjVAZfKM0VTubBxK2bqxpfqpvmhm26g6EK8ZXXlNDag4kvi55
8u/Ps2Mf0tYburq7MOiJUJSGSCkuLJQHTRjzBRAB2MGlOEhmIQWc0fsJ/UiSAUYYjB6iuPeAc0pk
LNuZiwl7ajIL7oSg3dS8HzYEYLXBk5U+nThSpxu1W4TJlacVu/febRUOz9izRpcz7l3Djo+nzA/G
lArG4LMrQlnTkQCj3HdcJuj09Eva6KlEY0v0WnFz1X9f0jT/xSNdT3T+IyNaMUC2eQt4uNQFTUMt
pw6PPeihQR6rcX0U5fVZQDM9+zxk2x8FtVAg/yYAa/jg3D5Rjwa39t0LFKYTPa72OHLLshPo6KTS
5HBYb/dVJqkhCsMOYXoTSvLvCUpkA2sevBJiS+aXgEZLkUlE49RkEnUjzf4A+eRIUMKatlyA/wJ1
jJotQ7U97r3Hb6wbi7IH5B2/GNET75+DH2V/dVskyPB+0CuZloYs1Nmh1Qf6rXgAukL+1Pzp33IL
uLLLStAEWV4oybDJAldJuDLNbvynFZxyqNbPfWlIRromseYlHToZOB8lRD8hvZKmdh/+Yfyfbl6q
sdpK1S4TbB3NuP3wZc6YQlohsmwx0VGqGOXz1fLx48Xxcf8RkQ+gmUBv9SlkjO4bi4x1Wi/ysbS+
vWBF6b4Ev2vACzvwp8Xw/bJggMEWu/33eXQu/bTsHc88syzdu2sTbHV01/Bue7Phj9UmXSncYl8w
5btgYMVv62EiNjv7Q5LwiW/ZdFLrnLkuQUbu4SKw1H3T2yKjPY74cQsrKgvNBA+LtA0a4LFEGNQm
H7xSTjrbo9YzV/yfsdnipouP7PQxH8gKqfQ2tTU0lO0tMDKlqpoWH+ccUXpLhe2u/thRwHSuMdKR
nsss+YsiqwdpPOtcZeyH4Y621FNdkNf+uPZNmtBSjOEwGDdvedM2JsLiCi+TsU07BSajBkOaGy32
A7/M5tjxH2kggj8WtMUccDVGd9CkuEWb3aph9e39Z2ylDLrZEj/yTqmTALGqwYwu0gcXG1SOUSTW
aC5P5DbEOD+1ChIxtcDOpyhnhPAQn4hqglcGzpYNT3tj65xvAFxyQ9wXg/HyhasPYXXCRGmLJOHh
1aV99oLmRyT646sVKLMuaLmQBOCiapWU/nY3GCbqJiNKtycLAugHjyq/LQuduHMJgvi9lP/pW+kJ
zpTJ0dOnh/Nkhte4LAgyR/wUs8OK3+AXr4TDAJCDFchJzVskTiNWj/1hP/2BHG1PU+dbesYGezUv
x20QxRDbheUqc0x6Uy2i8rpjpQzIsHPx3+YZhJbLhtdvYBRVIRmtsYfIpnvKl1sgsYy4DTjcl9eq
Z84G1YdCIy+NR2/U2qHaczuAxrjU2mHRMGNPeWi4dcpGGiZAsKdCvzlKme7Ixxo5hz2RF67xo5jz
3ibZj8LDlxR2W+YHOQe6Vbi46/goqJIKuf3x3XHrSRBE9wDKZMnmnlkAl1dpSeaJ7naaSbvzWfzK
mADSMEvsWbkjL2CcWDR/1ZUMkQvcXHvHdW+1w0y1KH+cMthqFWkODOoeGBIt34g/n1AcMCOCHgKC
01+QMdj5MoBm6FbvOx9cyvFBiPYPZCsedKKMmDC1Fih7KxdQ0boCCefGF0cuaSdzJbTJtgy0urfx
KyW3HxT5iXohysJSpPSkCyw9BaCJh7dp+laKuwF5jbIFUgXAxtWP5bf8KGT+ks0MW5OPMDQTprkx
GosvaoJT5/McQ9wyZvIFrwsKuQERnD1OKK9jEdsC+VZZ2BAPJ/ePv5MVYT/ycHKfjCQSYlwWj8s4
/GuVgCG/lcPE2hJO9oU5lTMXFoszQpY1sRM+GaAT2sAouhH/wjR9DC0WVqGSqcZ3MElw0NkSKDs+
0UrMijfx65gdoKjczF0V7+CSGUWqrqifK4zqmmmiNjyz1cB1YsUF4dZDRJssoOPDj5TLP+LYOtY/
3jcoyQh6t2knZ/Yrqf1NZ4KiC5qXT/iz4HbEi9sg3M8D0pkgPP3rzwSQf+25ayhowJm6d+vqadKS
XcozGNAPxOd2FSH9ymTb6w8IYWxfCq5f/pD7rQhbT1pNy3mcDmuzaQW7tdsoTvcUKz5oy61Ioql+
Pju4RGEP4SDVnPACAFE+hmnDZs53nlmXiwImsGH6HuBbNgtWupetkvKo2LtNE2x+lWxuTlRYHYtt
YTnTFyRcQNNQpdM56UvOyvKb/rEbsBE5ugPFjepIspt3mjq9qrC2A9SgymaUAnOrKRutaEQ/H5iV
7Iy9Z8EputHpijGUK6ScOmNyrNvQptD4UJSoa7dUmxlGT4smp1LpBqfaNJuBvb2Mr7zaKGFMJFQN
fGmWaLiOh3UqjTN0Cp6a/Upmx1YMIC+ToEPGi/TpqlcavAcXzYXlFr5HWhQVgN9FAje7WuX5RNfl
cfr1gVUZIhrCl4fgZtVfOgk+FcSZ3cVG7tvQsKpwQ2niKJsM2GDf5nKqpFIYhFk9k+uYCziJXr9B
FG7RRewiMnUCzCVBE1zytRKDS7DzBvACK8NfDQ8FSGjA/WtG1TRafhe6pp6NyKnFpyQudNKOwt/L
+3HZCQ7QHFr4yg49AJEDcvRwTNQAVcA66B0D5Xu4YQ9MzniICoeAmbGWe9lWMt1WFHnHgr/JLhew
xHZ4sFULn1CrusZd3IrmUdHmRZQ3Vrlh6Mu97dboIlczw/xt/pyiBm6c5VUvRG/xtpnaJ/S2hlNl
iPfrDuA2YrN/vdhnn9GRoQrBLDezYQINgfNGTJZY2dHA8CDKodanDzlB18/NHhDcG1jc+Eh6LckL
/lN661WLy0OfZxISzw8wDeVwGGhwvQcf1U1tbkLEcamUl1WQaZCfpxzwbkdNAKok3HDak/lNgnGX
sdq3Q+kuCc0TLb/zuZq++xEItPv6mTXg2T102L2upPGTxAE4VgQN907zDC17+5gsW69xeKfUGSx+
JRDaSyTFxoaA2yOwNO6HETaWPiopBS/BpveptYhH4zq6UxNaO7bGQYrkg52sdZgfCauZTMtzRmva
Tw6itfRlOzTgV4kn/rk8WDz1ohqudoVz2Nx13lnvKAv58uI2+Qd16mz7gSwxbGXpdQQ5lcAX5w7L
Psb5lpxbMHBG2FqgLB8zJryrthwuOUtOQJFxK3OOu6nxG2uYnTvmH5DfUj5UZTVq2vzQtSE1QJZQ
p0LwNeAWyfgotLSvE6N9lXu9OfQA+nwbiMYrHrQ26G43PCWd8vVTwqcMSPSULTx07LSMD8SokmaE
ceKDF/D8gFEcdhTFChkez6279scm3OorinUK6NYP25nyevCqDnQaqcE8GoGc7omeJveoPLKtUuLo
eleJO78ZzuPCQieJlDoJYX45/VLv4HGHpn2YokViFjmfOMyYNevpoUvYtI3WvBswp+ccKGuTlOnO
5Df0eG1AK3DbBggTss4YWeyM3Y8JJGVOIxae1ocYyjNqRLSSxHi00CEoiXu9bDyE4u1F5CCpLMe+
Cp7ddIgZjLmtT7tyhpZHrl3m545R5RepDxXIyl8Fa49jNlaPvQSt3KWwCDazH477rTUU2eWLxnLW
djn9ytuyvbkx0RcaukVCymwKg+03EHUOpEcyiAqaV0w+fblDBTtTDWnpTjvum+M7ydP5PqOrQ8Mo
0KKpop3QhY+I+GdDQrvaFAZItqPBWbCCTvo8Edhnx1vbw++hZCWsdrlLEgfT2T18/IPhPRr6sB6z
zBveJun9oaFWFupwj/GETDTSwjcwSyt3Rm7CCqwiWaqGZP54Wo9gpEYPMNCumcYfv7YfefAoG5Dc
Yt5PIntMYctCSy0dTCQD5DRhLIa0TFppOwrc1DPSeZhKDkGBf/AGUATsLRKrGEpJIk23KdWxpxO4
SWv7Up4IYX9ph8EDm5pMmvUkkI14XEoM+o4SK/9uxHl062qqg8DUCrOlSGZa/bttYFhZ19a3GXH1
BJ3jL5rNi0zVZqiTonbDFcoCQkQklzp3UmgMwCjvyqDXZB2gDf1VaSwJCQee6kar0NnF4mmdGMO1
gOOrx8cTe/qSBTqmo2s5i8Mop6zfpdmmkuYphzKPmmW8Ceey+EmqnkkKxFpLO7nQFi9wc0ImVkda
MR1XJKv6Su/sgh9xAziwBleNncCori4HB8bBiuuMy5v7nhKCuCL28ers/X1DAaEbARPZ+DA3ojDk
XpsQkpFAtR94abWKSENfAdeqz6ZTXmfeGR57jgBO6k/yM6Gf0JaPCoGWFv5cTenm7Q+UNQ3M+j8K
P0qn/QVOX8dqAj06C16KGzAvHQ1Wvubko8fKocgsITOKgMribTs7uXo48VC+5VE6y41sXZJ415pZ
eN+0RDR1gsFI+ciKDiM5PM0wMjcfrNzWDVWuk+LMEWelFOqOM22OMpfxPOjlDX9RmLBaVZLgy5TB
AHsG7YX5iJeAB9TKrC6SA3US1Xxmpodc4khMikTyfWOYjZqgFwiL7ARnGZHFZHi6j9pF7ZAKlf9Z
RRUMjxmDz6DJMEQTK4mavuxdcrigJ0dJVdt6sYIqNsF4TEut/m+nz4P+g7I5PYV7QFj8SbY5DeCg
q6Ys/ZdPE8JF//FE6nCNCNry8iGS6kahXHIcMehhW49QqNa9KM8mJuU8ScVO3xuMAlIwWJdz+l21
AseogUPaIElClHHGQIeVT386JkK/OjVP2JdJB/wzGXRWrHUuxvmGTDFr6/qMQls5ovRMmMoQZkJ0
TtgXjCpsRF3f96jngrK+F8tY8xnp/jLyO791w8pn61425P7fZpPhz2orujKMMNFVQeOhb4OnhsbB
F+k3abl8juk2c/IVCVxYBK2wY+FkWpUbq1474lFZ3Hjx85tk69IKMIWUmD2SamW4jQgzaGzsPOlH
wkQOSf2TfXhJay21x60959SwPPwqHHyLc2lzSio+IBoBXpxHItMsuOuMHDSw65Hb/qvFY7US/4Fo
KSyRAqSvv4qH/8OZhkNhUaK3VFJrfKeiuLckByenMYGqs43wroKjF6xVasxdu2zlZ5t/aao3mfOk
D31Y+WmOE9F3pjwIY15d5093SdEHNY0BXer0E3iZYMT25yfpEaMK8dzcnVklFWg5DegC64OKC/XG
Q2tei9lraLnmHGeDFvh+hZ9aUsgHrFlLvw8HF/qMk6srSbJ6YMWY/QmwhRYDjMniuQ2tT8akipd4
R3NTbTO9jzlnmksziyy165KnRWM836Cfj7IwthivvVK3bIHMH86lfuiQcGWXvQGh6dsOxL+OVdPr
lGRXwg/xFt8t39n4EVcYaYqaMUCEow2ZugbYM9wpuc4ShOQ3Z3kZDuAoYbz8QiZ4y8gzovCNIDJb
JpezrUMmfWlbxg+X6ShvA7lQ4tP0flZk/1tPYGUIoWxZfoFTtrGMjmZspD1/RVyPLxC0noCo0rWh
591/qjlebpY4t92CIcYQAW6nd6IQsDc2ApK/r650vaeEAso/ZNN39M1hpCNzY/IVptxQ41ISE9DL
auoDJXF4RT02WTcVJ9db+Z5QkVaGEU9cX21KLsQRr5EUg9AXxMFH7BBiD6/77UtAHfhGMgRwE/dz
90uCUmTkDQahbqhx4fAChKaUaHSusbLD4u6yEIkMWw30/wkFnNBC21Ld+QB1OgaBfnjMj22XXvDX
HM8wkM1JnXWHL8N74wxVDhoen9pHxuBb14VXiz18qUMlGrTLz9fEuESilXWgx0uqZoqIsg5nLD2G
3JcWvA4pKniNNqz9+aVVruQfIg2yr56OWNsvM4x195LqknbwsS2Ai9D6g/JuGWkKCqsekU1XksKN
IJ+bCplqdOjkzMwVqOba9otcS75v0PHkZ0f/aV1YR7t04uYJ+OTmD4BJn/L64SxvEZ/6U1IGMwmB
NiTBXLyTAjyljexh2a4z4K3CI+2GLOy88YVSFTnjFZNDJjlzPEx/ankEMOASazsoxC0w+CqVqzfb
GCgLcuonVyMH72PWc2Ae3VFUhJhZeR1lPZ1bipSE2i3INwv51KoG7LR1Vnd9eKKYl08nqXC5/Fus
RgFZxEeB3mdAW2+hQ8EqAQ1D5URx+M5jQ69/ar9V8vs0WCO8YNn615LsPrvsK11diJ6TYJuCGzVD
Y7GivQ0cz7r2mGJImQrffV/zvWz6KU0kA3YLnvRGStNllUj9MykRG9Q/rp/p9jn9MdesocL4Fa7b
UTMLFWGGNkR6STHgiHi4WGN1swh/sq5WijahiD8bnHLadBg23j/KpklrcCF6gcGvLY9+UiC0GtQ4
NYVvOoR+OIw4ri2s72j/GXdX3d61DrrP3oYNlXZRPKEc1/mTNGtTtMoV6At4+rH8agrbrvIc4Thm
5jB7Gdk7dMHluov3lxpjXoYvnvZdV89vZSA59waafnJ48sN0Sv1N+HhR+P7dsfnw51jxQqijCyyi
27rSFEHtGbbDUAA8WLoSbWbgW2WzDYc5DpFHo3q0MQpACVJLNtQUIZcY1eewXUUK/dsJWk5WuqxY
SYWprDlU9SMTn34P72VnSyBF9it4Fm8iIeqsyHlfutcwdpzb/9zLmtYpA7HouxhVKsWmyj9ZSIvW
9E4iM83tmJRZBOeupASLnWmHiFZfOaR91HfjvmKrgk/+wDmS+zEhKGo1bKVjDuoYDueEGmvcAhFp
Gs1wf4iPAByvzv2RaWC0Qt3qTk7i9sXsRfjuHBMXyYG7FtcKQ0B9J5rSStvrWLGlB2XI0ZLpfgXF
EK0GLZI9rbRuyOBzLMRb0BCd4qd41CwJvkaABiJluuvhjSwH9NH3oVHomZ+nPQADkB46ZEdqLKnA
1aquAW2fB9MO2aO4SO68tKxIExnvCdi50mnOChT0oBWY1ybz81Uz6k3l9UUiovFYyDGQIgEl1E8e
EKYjPa0DGvBihcEJhfmlZoGbuC2TSpp82diTsWHejln3bEQ6WsTi2GmoHkb5LSwlp+NCB4E7HBde
fN64LTkGjmZP43/ZhEmplbA/uBGfqvlnIBOkdbnu/Van0SuVK6Vl+Plea4ss36wqjulqQ/6mGVNl
X8af3NIdGpypZad6X5IBKVcy2s2H9JjOBBE1ODwDHIPXBHq1BJ2kaMCee50yU0ORigytPdh7nUZx
xHpW3EMET376wilh2dGkPHg6w1V+Q0hJOa7ys/seT/o5RhhP03Poni86oI8HCO2gK1+DaX6SbBMr
L54mypPuczIPqoeJDuFDjTCSng7pTmn5LKR718s/EPGIDcmR7LaWYut5RW3A0CVgfA2JHLqBA3xD
mBkKXtaaJVS7fbPOzykD49yEwptdzH758uX/jqhQzBelAR2cp9b0kcVDFfk1mfYuqROP0BHC11VW
W2uJfn5r/JDzJfFvkioX1oAv1n0/zuF0HXazeyvZg3fe7ufvRjhS2s05zd6uaQRCJM+wp1jgmTi0
TY5dqUp1FIBHKj4ECNBmOjpJe/GJ1pia/u0lEXE+wwh/cmglvgNDKYMPAwzHooBUFcZBT4U2SCNy
wfpdgD1lcQ8dm50XeAbkGwaqxrQJgnnccJGMWDzAQN1ujbZ5BcQgSfKqZFcan7NQgu7yC0SWAsK8
YXoqeI6EYRPtRj52Fkf6OuISeTvqn4f44Kzfo8VTsPBT9bwVpyZunLXuWkf3FnXMuAxiNQykI8Uv
izGCR4TMghFMtwpvUfGMkqcK4k9ZP2GzDY/G0O3rp80zir1kAu8bk0Bh70LbSlTve9W4xFmfH2UB
bkeBg8JtZCiw6mZYpaNjMS6QVLLaQZPRg8UuZnMqMSgiakKI/7Znlqh+F1v8kj+Hvda58PF3cOv0
WcLHOUz519Ru/mhpJiqxYJIOkfO+ijSEupNX0mxvLsAdgsaU8SM2JgqEOwKKda7IoOXHzKzuGeXC
pcWEm2mTYV7XD0DRW7l3CjvjQsT/OEtdmTc+09biWXXjyLh8FB1alNdCTVegnWndH3Q7tmptMA+C
r7QoOmrNaXElZ1H/RwBEFCN1ArWNzqujdwM6JAqZDJABOTUbNI2KRfd+b88t5GI8SnhPL5CtEKcP
kEWNUkzvLoZ8s/Md/SeaMXx6ovt0ZCiN1ufoBoO8RvBOrCpqTMCHKBGj5/4VbmrFfAacWQTqUUiN
smePTQtiI1CyvHltNDu3sU3F2PrOppboIl6AC0b0JqDYVGTW9+M8QfPKY4dEJ1gfZ8zV1sGKZ82B
WcBLvbobmcNCzL0VU3wfN5o9LJliYft8Nb4/7hC1C7RT6ZFvg3dAYFUaXjUkuDHPW817u7c2Ruf2
+oLiR4LVXSHhk32ttLZ59RzuCChG1jZvzKhtnyAzUGnXid431I18Sds2sCa2QhH+Z5VDrBOH7Vdj
Ww7gZkGyvsEbeIu7d7Jfp4bS4q+miz8l5aBaEScBcWLNCznMkkA/gMUT0daHc/c/POFPDLaq+ETz
EChDfrBRvBNAVBZST9k85NJxbDCd0Be7oE3p8OS5iRVUkA+84IkJcDie8lEINe9QfR8g8KhoWZbz
oD5xpIYJa37WeN3AJtQrTE/8bu7x7Deons1Q7ytH0Vwr3Nj2xxFBd920m+HpvKGz9v/MlX6K14Zx
EvkoUskgbdUbE5Atnb7M1ZIeQQ1ab/JMymSxUb1HTLlRcdkoph46osSec6luY8v5pqiHBoQwhXNC
tUGpOS3k9uaVUWtRFMEtjdz6O6xpO9ovZQNU2MsTLGq5VxW/FM1cA836b9t5a40fnlYmnLnDw6Cr
sgW8uza4roQGn+MCd7DEqLJkkWXiZwgjicZJeqKGoqCxdYAOXu03btkK7pW/4TFcy0sDf+4qoNAx
nWJST8lCeH7uH6tJoAaSq2j/p2D6dQcrPZXFcYkDMmn6Er8iV0aLe2uspSQ3vx3rRLEBwRdUmuU/
EVLCGzzGq6U4PcG+Kv3OV4g8YGp3lE9Gzu6V7BfV2A5oH4jNW5MmRIHlS1H/ugZWwGhUl031VCuP
L3eQRGPAfz9v0Dlr+tHsxpiOIuolW0CtmIHC1bLU7bMLsThI1n4N3eSMhjVo9dAWgy6al7ugmbgJ
Ntbl0IM1qnE7EHA4U6YV5r8oKu8Gne+NGshJKxzdt4lHY7xrTOqwRYnx95ajePwS2uDUEKKJUE3z
VWjNMFax2yCRqka1EfapZ7PVHncQE3v2vjyNbbJpxW/l65+PFeOSuix1vQceW8514NYXf+XWoVLx
gEc48dS/GS16+kl16eSnbXINb3hp4Mm4VKUHEphLTdr65pQlbdEP8aLBhiM5VTNTV8yN6CYoTcib
rneLqCUPiaT/p75rV5o7bHFl4O2lzj2TeofNtiNVKopCvAwrAmSJbq+CI3/FEYCiZzsipdvSFpvU
BxQXQzDGlhClRbVodc+DgTAskaqUUHOak9XYNEuvdgvq5XYNhBYUJMpvYl7/ctQDs9MDZRfhDR2K
9BOYXGjxEp6A4V6NZyIGM0m8uA+SZlTG5Qsw+B+qwTwhUWhmOnNRg0iy3Nq5zt0C40tZKDogMyEZ
vVXQ8EdKJ9dDk1DlziK+lKvQUUi/7hwBCmU85TlONxM8E046EVWQeb+j0jUYM35rtfp9lDqf18Jf
dnh4MFrZ6FGwxsfj4bFKcH+vwJpmR50E3AMl5lwrhU3QCbkeSY7s8LxsadJwz9kvJgEp7/iGO2Xq
eq/aHWfmLsEPvfJ2htO4nRCHMjWxb0Z4nrBAlgzsazAqUK1dnON4eFBuMJR0Jq+BwmewpNKB85LA
zOTRTRowuhQ68AsVfGnKSosYlUgr17mazRY1Sy3qf6iDqC68CnW7uoDIGT64j8ta14FaMiQOGDDq
cAPoDiQzkp2hyuKenbeZ7fTHPXjs3FvXfvlHsSBPiXa8G+24sVGdiGe86SoC5fFDNOnUkuPhwZKL
a3vEVXj5/eXU1FfzHowlpArLM7tSNztKvpIJM+h4w9PZBO4G2ondjxDlQjFuZ5oOOVyH2x92CThT
Gy0CnEUl+4cLwBCtLwez0eAha6PLXGkqDNBzLkHV1GFYnlW8VhEqIYivL2CG+oOtvHWsqMJXPF1S
Gi4Ff9PvdA3ORB85DEv9WfZi8IuKLgPB3q+vpK6PP1X+6lS8QDRfT2gtTgiXnxoFsQjB/vj4xGaD
pVyL2ZU5plEoam5X7VJAYf4z6saR7RatFFk03TVF6povWCmfcpMcccMRoRjLFPOqkrJ/yR4tGrRX
gg678+LQDXiQObJZOcPniqKjgB//ScWf1K8RCrsNuGQhAsigVUkF9KKGGBQkSndWmuFPv1fVu1i1
Z4VK++Z4r0Sz1Be88gwhXOQpSnEsgEBtb5f/e1wnl0ff2ZnnwazrlbNxeNbNlgcOLk5lJodWk6cG
3xKXBGYCumamsgLHG9oVZ44NiYPrtIq0dJkDQgvwFIi25Yo39lWAWf4aLV+bVsqQRIRqm6+9JSYL
64iKamrzinAKFANnImLxLh99jtG6bXvpI2b/8p4N4bG7leWRjD9TTVthuVnFpqsgyxnLflamOtwZ
pZy5eE9y1wuNPfr1o/m0rTxjgHlRo8aSuLWwXYNnJh9/b93pkiJn7CSVGcJj45meqcqFUDY2bhlP
uLM/r9n+Af4y0Za77PAw8l9Umd3gcbWycFFcJcd7QWSt9K2Wrtz8MSzW2cCdLEfZvAhJptnuibI/
cwU+6ZpkWSJG5N9RIUnDoOML8j9Iczw9zzSlHiBiYBMlwFUv5XEUVbpJvW47u3J4ttPaOkF9LXSI
ds8AfE9ryJVO10vjm7ltr9eeMwZabRHguGj56Troa9Xg/A08axuJ3riRydlvzNtqJ51clGX6Vb4v
5W9qIoDNdYQpwwkfI2MXEukB1Cm00LVVJZ61Q9U3RlYlv2sEx/ZXXhVjLd7jsIHNDWQA7x9XIn0m
FYcUlncFYcvJVJSHsnxdFn2yFCWuPXLuYqV9mQOp2rSxuqUQLKuLmkXhc7w8jKxlHzLVJwhXnKtA
nK/hOKOkiA68dVb3eGzW9ngOCeWHkAti3nmk2ixC0sZn8ejGgnt+5Smv7QXyrerdHCoU3T3u2CTd
c+IIOfa9fKXwGF/sl8U0wnO+eoO+OKXmOKGQgMdteRPvCt54856+MbrT+1HvcSkFYIqS47cTEkGh
S9BkeXd2QHys3C4lDQVaKFoDq0H3U/IYX5ehHuBVWH0xh820a9YZEK8CfKJ4Qbj5F7KbORVNsJ/d
7k7wrIkY5mNw+LMa0VzYHBh1TfMZB8RXF4t3t6i4F8dDeyUN1Up/YJs7rKh/oQW77eaXX8FRUb5u
9+fuZf3eNYwN+WuNlIXd3dvJIDTpVo8lG2rs/zmGRy7v2pn7k8UVILqDex7h0gYDNPQAW75JJRQz
6LDdEjxfMV1vaogCQd6dXZBOb9+LSwVdVpHJv87Gpid/SVSbHOuRZjyXNwQ8c6we2PwExwNDRsT6
9nHkwF4mtQRs/fJKt1p6FHa+QFIFdznQYRPnf3VsIcX3/iv9DsE9Kb0VLmqS/F9OzbCireh/r2Jg
1vEM60E88sDiE758xd9u6TLKj9u4IxlCTNexeQIMNDNr9VmqmSmPGnAth3fUXv9psafvK+dHuPjd
n/Vu8VpzDPCqHyyol0L0CnayRHdF/fhhC7X7/8af5kpzwsovVl1C4fOXwMlpFAjJjajRcAywUs3X
4XCcgExzs3wpE1bsdyC+Z+ynCFeo9RCYUkHhL+PgWlCvOiVKLiRR26c+PIaUp2M26oqzUtIDmiZE
g7cxlW4qREZ+G5s4kPSSjjAOfpMlF2oFvB3WERxELIiJOCJmTozblItbkZE5wTHvFk6PXPbUYRxh
JG3SD9cL1kqdnMtff8ih+LUvAMTcH86FGvL9VCwA5bFq0WbfQd8/eqEFNweCHbvnScXDTtPePIaB
+qJ90PGFDR7qbdWoXjLjLZlZTNmh/l/QBNgvopPzaWJso4rt9f5HSZ+oR2+pS7OVwsqXUV0mbM9/
3eQgbRc+8pSQPoyrn/xGiJtJvIxecixA7nfxT7Uk1AKFX5IaMYaQIB0irWwxJ1Jio6eTKsMv+Adb
aJhnksi+poUJZcwm5yyccfNQOhFlaxw2dg+uhv6yK9Q/tUJDzn2FSp7WoY164rYSCoG6/YIjPSwM
JKxE9EhoYPmhKxVESzI1eHDliFnrGvGlRyNxME024WhiHJDuK4dMWXun6AjDtsWymbpMMDz3iT3Z
Qx+KNO0wDIvJ2TE8DWJLQCRcqW5OFPS4FYCoUSxwbV4+5eTpnq9nQfTUJWmQ8flk/es/AsI0D8Rh
/n/WBzkvqRGqzXYkDW8lU8fj2nKEuKaLBXeHS2sP/f3MWKgz3xVGPB+3TCoIGaUw/pIxM0MndTx1
o5WTmwcuq5+HE+UDQ736DZ9Ou62LRwJcSp7aH3L2DmTBMBoRQFsfmqFCg6ZQTWHcEryEQy55MoDW
15ErdNXDJ1fYTf5ElO3xIYytvmlgxisEHoHnGTigrnUECc5jyY6e16+LquvXK/J9sXvAKYRJ74lM
v3hmZnlkydVuNQ82bNTywlLKOrdUyyGArtn8Em8BZZmmkxwnkiz8JtC4lr5VCppV3P6GSgm/PENr
XgcrHNVDipo7//l8EEV1HrGiB2FYn6vSefWXjst/e+lbqo4l6hqnZO3D0VkUXYLvqP3rIX7C6v6G
D4jddVi8RHcrQC2B3xydJE6EJOOru6XrebmvrzrodOAkFNCnieCaYN/w7YvH/i9E26qyZv7/vdtd
MbgFOhuopq595DOXPRBsMRhys5NqK2e8wVZc0hb3krCLmHLauFf2bR76fzQ1xlMmVVYvGKk6juDt
MfEsI8Sy87FSi9q4xK6cV9LxZb6pLXhm7p1/hpQC5qP7vjzT6eoYfTZo4OhWyx/HgUVr8ZLoyfij
sRj5hjS/PattA8JqlPUAK03969KTzTAmL5NxqYcH9C8+NT7Cf5GDfO+VqDRIVA3rXk8G85V+a3QT
P27pA5VP7tkZQasmnp6Mmo6VWJ2FWYtrtd7ma7MBQGr6zV1X3P0gkMca1D0sy8JGjPaLBEaIxxYm
g9C3tM6Lg3BYAurS3N1qn4JkE8Q1Mmyqq/mWKSKa3agSaGZR7j9NxsU84gXubj7RKVWnzT1sW2Dt
voXDFvOwz6e+sQNLG5Gm8BmQEe/Jhak3QERojFHNE8344n7v4dprEyR3R3Ilh0OuB+LUsSRVvcn+
TSwuUEc9brbAXIhjO3j4G/0CrSbcJChvKSk4UeaBgXxI+SfcYnc12LFKMoMdf7ua3lQo51d1P3lK
T/QFXtXUV4suBqXaxt7hEz0DxL7GriPszccBRkTumDKeWk261uiFhZrxpCX0QxDAPS2rMLpqIcQL
ioECREZ1g8Tb7c8LQfUyRDOQ7krSezdHNKTfKB9XTe1V5BE2m3ACVbokNqjYseC9omt3vUpnYd2R
BvlGnInKmPKykxT5i5jItS+aOMV2al2ia4PILXa1BYgKmg+c/uyZ3+how4LuizUvCToSBZPQwb67
BemlY4YK2pzMeaocuRCa2hq+UspsPA1Bsw2vbZHPA5t5VFjrHiJwcgJCAUqnNDM4QJ0/EQHtZkIY
xKkjst5d4EvZ0um1hpQoDDiCJGKybciOsMQDd8IxlBazB5w69ZR5mBx43IK4qQy8c8+96g49JGgg
vAP6kIHVawX6qVpELxpiOp3z7iy1GGSyCc5trlCV2RZQvuVs74hp7qArNW46P8bGnBfrVFPE2Ti0
Zw0uA/PhvV5RLgCPPG05EykvHjote5+BfBUCWbE+w4mpKCGUsoUX8T2E7K+kMXUxn0z2mJWlNMno
mZYJyqkXZ4NeKu7DLkEyMXafU3lIQFXhWeErWPHAqvseVzbQL/DVMHzQ8qKROZqgdl1mr7c6M8+O
cald3FXYzTTONuDvcRXXCTFCDqgJkJBqBVOKYXR7FE3uddToFG4Dh7xzwRHwbGtPGVkJkl7o0l/f
xrqbN5OQd61XXAro1tYrrwquSV78t5zZd3Kq2TZnBOnKLMZTKjf6VT9+R9IRTmwTbCHMbjhiT6z3
N5jt2ddFcQqY8xFqjT7BIobjNp5p2py3PxH4JZNAPDGKhxScAq4Qeh1WEK4aO6AQQC6aASoG+77w
Krr+2zP+pyGt9aO7wm7UU0Sl7uBNmlRJkIeJ2CtvVbMGFbojL6COrzF1B41YL6ZB6+xgJG8hIj/i
Vz8ZSeRCdY9f4jxJip6YQgLQB58RRI+RNJNOc3dtZV3ufSAHUPye028TJlMzKOoKRQtsEdhzmEJG
zY6y749kznOkmP+0+xnrKB7iZLZxAPfGiQHua62k9ZowOXR3Z09RjOEdNX+Bjnuk057F6m3ig1iJ
NszFMfAwrKK8kklUGCGdJRCrI+/mMesAuIElZJ2a9DOdZ8WSlOsdqK/kSOmV6a8pSq3W2hQkb9Le
sZTbS9RDXHBZeACqr5KNg8NIn9yCjcj8Wr4xQYsCoMpIOzZZXPgNWpX3p6Hl+gk2u4RocFFP5L8+
Bot7sHtTTw629pdwPJqeOop58jb4/wEwICZeAh4GWXtCNngqSIQ8M6cANz8EoPqZntwNkymWRXcn
c2zDPaq8AyXd6pUFCDYgcCJzQcEILcLDdbcnuJcWOAASk8Y4Y3Y/q4qqZrATOLIvDRGsB6itaOj3
m0rvAEx0mQ+S/yBzHZ+OwlxaY3LXuULgeL4KFDivYpQCwvt2iYV11x8eN23CYpfbkiltCYjNIcng
CDqmbtZrCaDi0gUiDCXEL5q5Cpd3vj//Ph6JbZ0pupHbs3lZamQjydPauiUPF9MNDuvmjlvgfaRf
MsccEs23qreg9Q0rf5N8iLKuJwbn0x9EUT9DNIf5lIDpy5hCgBqPMxxPwUJ99y9BcV8fL9rlEocn
ufR+8mmY72q5fRxaFZ1yzLTW1vEgPkq+0gmaLM9GBhDLkY42KAyBjMCGE7v5Lqh0RdYVmPY6QFse
DowRDCrVe9UFl8H0wpCalMBCFDHcCzu9B+ZsZFUyLQSDgx1r0nPxLwVZd5brxvbM+v8SNl2FKZ+d
V49YCph6Q/u7JqtqUZGh0j9Y2QgD/53wVkNd8PlGidUdDc0wSUQTKLQhwRBYxz2C1cDRuybDVgx9
eIoUl46Jf818KmPyC2su7ns3lrzCIOACGzr00yREbgr9ASd+xfsWodHb2ucWrB6GrVUCIp4frTeE
8VPMuMiH0b1SIEgt1T956gdJ7qRlA/ikoK05AO2KWtKfIWlO/m0oTkGq/99lk6mdt11YZUqkG2Oq
YFfRE1LI6b8f4N2l5prxFzHVuuhfWiSfUw5Vr/AjCQChYAM70Q/7i6tq9GKfYSoJclu/rkcTo/Ha
Sm5jmtmkpdjxDffSeYWEHlZxr80KVioyVBv68SGzhjJO3pv00Z2quEEaDGYSERVL5eR/ju/CdzhX
RLzsClozhMHOGYyCqcYK2KWEu8noLv+lPeLtuDBYBhX49JrmAnRy37V/LiDGTmEMyuV1fA+Q+sTh
tAxSup/tNJ1Kho9os8BDrRRQlQcZjhIyZFJj0yXnLqkUxRfjv5Wl6hzD3/t9k+JXN12UiEAa42PH
R/loEQEjMUJ1hMN83oeC6PnA7RdrDjb9WTwPWPDCbAM9P0TQslzX1bVRtCwGDWGIdZFSHFz6JCrI
44lWgMvASZaDt3LR8MzQkwyLuxQeZg8qmYZpIzG8me3jT72ZmJPKjSQsoHIYKNvrcchaxpMjkUTa
lTyHFxG7pa43UipGIvwRklaH3bdDgcmPj4nl3WcG1jV5bRfsg8hATJrb5lxCXTArb9Z2m4vg55yc
hGqB7f5PiYZ8126keJawPDQvBeP5haA36gmCf7pQOmDXPv9uLaCjRT7AQyKkjylU/IPVSxjVG0FG
v0foMB1y8z3bs9mfu5J1ZrJhi/vHz7mb4E1RBuupvX1FQqF98aSYeOUJ+DKwqd3bHyQN2Tb1O5C/
TRTxdFk7thkuQ9OLbqfYT+VAblqdsiaRrqhXTpmpgTqvxsw5GWMxyOsnfhBG/NzL69HG2tm8UHPX
/5tBPorBVW2BC0x/WUGKLSsMGW754dwc+caVDsL37WgXtt7JxI4znxw3qACe0kX2Zg/FjTuifn72
9G9NYB8zq5WhDNGLGoW5J4Lc9xZgqZrjKLq0BGMDIJVxENumcp/oK3qC9HOW6sGm+I55v/fhIpsG
cP4vT4zqknyxvEkNYgqpd4L/IoLSpKC41KJPNxIvebk4QvfuEAy2vtCPH5G+3tBk1Sa3KQHeP2tQ
2AyVsBeojAmbDSS5vN5TY+XXz/A2t4zPSCCTRhdvx4hvKS9mXMy0Ak1BZacMYhBrgDltJRtkX2YQ
RIrqE+H9qgNEcGb7rxN6AJ/EQxRSREUGG8Zbvp+oKu5o1WBJqzPnuJehqGIjvFjxPaJ0qopyRVsZ
PtBRCCFA+PBNhzir1ix6RrZIfm9lF1lPMGbLnf9vxktYI/quQxUYC2i+zLNHgGtoKL5UDAHnNfUy
Zvtnq9kHXieslXZicx1Wic/jSxBCj2PDJb73Db3WZ8LLixERNr2SJOS7yiYXtNL3op+jTOzSFowz
VZhRYClILz3jJIVlkyf0ewjl3shYl15nm93Za2YGust0zO62q84JluSprIJ9N6BnamMoYnRRbYYK
4owiTHsdp8XTcMBYCMJfx3jR2lrU+xnDZDg/d2tPpsshctX0MSDUX2+OWoU+2qU6Z8ot2221fClV
q5PAK0LP4UQqsLvARiKsaM4HntxT9tMV4gy1SBAMH7rHKGRZJD4iK++xx1It/7OPt2FJ7slNxQf5
awuZJWIbXtaE0VKWZg6V0m2nwBQ6JOH3q4w227p4SQAh8CxQ51OW+wwssRroRHLQlAhO/MoDfZnv
rF5siDdSkwZOU52VeHYxHfaC/aePnrRIPzEqmsaNEkWFmElF+oyCrTjsuEfZznBm/E+Vepv/hrjh
dRr8z59opvfz9vvB4Z6Rg1vBdXIY11eGWrBU+KtHzYO+JJSEm9u4gcmKAsC+8JTy7KndyYJcIHoY
YCuICIbcv0JjFvLAs6V1d87hmqHOv32Enx0ws/XfRuJEzXLGkooeQjbOJaSSyLKGMCMu0hdCmJ/L
XghnaRybX1qS/5joaOKYEB3oCrREklkp8lOt4ZkN0uDIumgu6YgMzb4ztrswSilLt4MlnhOU3Cdz
Z83SfKr7kmk5vhxi2L7GKzHHmwGxxN3w8rUXlz7G6DOI7oYVUixvHGsSPmbGBIJNRSw0mrCpUsmm
XEDc+NgVqTlf/p29RplvIF4K/2t+0Rt9RSweFkrrAZWVNm5WeD/fzrjDg/EE+YAO7+gbo+mOtbbe
L5hPsSwh9IEZjunLs88rMBWPy/OLSQHdUSnRR6+tBy0SrcTpiPOBKyN/ILRwyYw4Rcqg/AWkJjwb
oyajkezmR+pghD7cNSyhu00yrsbPaNDjpSDAQ9zrTa0IBDpCNhcLePpW+OjXfPJBPV3WExiHU4YG
WkEM9Kvfqh+ZrQS1znzT+L10W44R9xoi/GyM+GcT4P0YGd6m56lcGo3FLsQtlepgmc+IOeLrtWgo
6GOxZH8Qan+KU2m9wQ0UVVjDCXoxcm78Ha423hGmk8KeBlfILalqOM3xfQM4WpCE5uzMxqYURbRD
VHcaVkmZGUoIPactfjl+bYZyGnk4irkoL9EbdwI8cocFTDftOyhA8pKrZdUDM3aErF9048dkw2W8
S2oJr+eEt1eqECidPBueTkkbFZ2vOfytNrX4tJPn5MmTZyNxi1HXzxWD/Pk7ym+LTmcAdVAunfdT
mPUj7AhFolsw+3NALmQmT51QkLsvSAGKwMPClqzo1+1eCswKPyQOJ2WK3QqAbEg8TBLTheH48kF6
CIUYILV2biAKbzNq0+fdthgrJ26JbzNUucpEyfvVWwoas4ZKHfb8dJXCZPoK96QqY8OYXfltBAPR
YvOewd/XYhU18iFFuIeQFkwSw3aDadUwpI8tsD+NbTdhJONkfQ4NY/vpaz/OhmcUxfdZA4N0KtjW
eV9mgi1LVF2lIzZc+kb6teW26JvOzlVoWOgiAA7XSqcG5IHHF0YisE+5c6ySUB00mSdSOyXLMnzP
FdEPbjvolLRZ+UUGMQF1LdKtJ22no7EoXrfycs8hM/jAzcxFwXVn1n8c4B0BXiDl/ufOaqlX4l0p
FYAI3ljtEDZPXL0WvcS8wZPKdTG67gTdtgFCFD9SZkmi1rmy49ejSiv3b22Bj8rDRIN+r1S2BuP/
svoaqqSEwTPEl0zo2aZQkWDjj0qEhVP+zS0zLd++mmZ0k6aCfp85jH+3YnIYsu+hz6E1fTbrKo8m
zubKP8jjkNU8JTlwF/4rvyk3y51dmiZxGW1hVuCNE5LAcYMclGsby6Se0QIQRr9KiX8RXUI7FUjD
lPr6JRSwEn8uvCt/0k8hvh4NEVPFg2huUfWkGOYjIOdYNgZ+1usXNF3eL9D3exteYCsuOJ1Xpdzj
IoZ8OzK6ZmhWlTb706hY6PwqfO+lOPEqXAvEblHIJVQypsaewwH1Ldr83+0cbAOOAHCaxJvqUEAz
6fkBpRAVKs9bPlaV3/X/JgI8197yv3RpTa06+fLB71DB5zHnfig+JfN88TX+D9jYO4pnlQ5g/9A0
5/cBkY/cgm616UyQKgE+x4cptOpYeQgJ8PreHR/486qgJkswaM5re5KxTzgnQ9vB7Z1vlmb3h0Kd
HXYd0HrxtK5XVGsdiiKKlCR8tc4+u0/KXkRl/1qbOtM9d8FcHs5/+8zxQgOqaDxAELNeQIAnSb0b
UAqKTwvsXqsrkOb+fsBxV1ac3wnlhGyHJ1HL3zN/DKVOSVikORiWEIr5BUda4ZgeadZu65kOkZac
OIQx7nr2EXtLWKd9s/l8W0KWacR/aJ3ND+nr58py1o0ADRRWdVCkhp40eS6ar1CP+3+HEF4pSBP/
S3RLaSk5KWATLTHtVWTp30mo/t5xvDJX7finn7p9C27c8ECfEW6YmTZp+zlUQ8an+66jhrNWYqRY
6XgXv1H1Iq7L4iDy/krOz3mwIgs5aQ6KBLXgeSbmraa/2MePfabzs5tEIM6M6LBJeahkKAvdzl/o
8ZugMfojLCoj9AQ8ZqfakfSL67Q4uxGVqYXB34bULyELc7tpoE+IWwxAfvWckDlat1ZSHjvErOZ3
wgetuO84rHXlCmSTHEBeMJY/OQPMEmuSq5kFC0StmGFxo+xAlK3VgNhDEbyomxRnxck7BFErrGBQ
ui/fUleqOmE29+6Mj22IL1qCgMe27f8Fyh2zGoA+nmrSQZTOs7n2RY8phZi7+n61G09fm7qRIC8q
5JIluEKZvFuWg359/DRlRBIrGap+eWTDjS5FSwNO/yvtqcEXGZH4AiGgWBqEiYurUFfOHOV368SP
UEUUzDpF5Uen985b2rUCpJR3olyMUeER/agb0IL9SrKMigkoydFkKOUiL4XlgQnOrCUaSr8schQV
HbYSBJl0m3AYHnlSC0+lCWvPR+uiXDDQzUI5Scixbj4yxKZXSIB3q59Mh5Pq698m5ENXx48PkCwn
Zd91X5lsve3YFqfHC1cWgCN8Oyz+tOsEVjIxUMyPy0ODeSMRX45jiioGaEde4zbsCqXPqflacLJD
zt8Wn/egi+FWHJatSh+JWPjcIvgj/1ZfhjLpBAGGzNZBMcIfCH40tw5WX2KK1pS6if4z/M2O+j3b
40NIUudbQ+pie8KYS+eXmBOVijBubvZtbPpswnV+CYD2fKcVXIQO+RucB2s9Z4lGQ2kEHIq55rlO
34KA2utFEVpu/AQTrbDhOTIbirTsSi/5mWMbdkvIDOayl5+YCeKLvQsiUh9D1MUOh62w7rSQLBZu
Ch6dGzgGZHfDcTqy8mbBjFgShPnQLOscFq6ZT4KzmcrbTSO9sttb1WhoG0JKxNi436s8bM6HipgZ
6qG0ST2MVS4tL1n2UzoaUbeVGQUvdkEznOq6HcmzrwyP8xsrgjYtyyLLyePAtgsItXqgy0DvUXbc
eou4mScE38MINNkVLwIZUmhb2vb0F6/ZKuK5ou3tVfMyjzs62Lu9Gl5uPybpdV5sChMrIxene8Ej
n7uE42O51QVUOkSqCdhAvjNYD+79lS5ARuKkH8XSy/RXnYdFIGxTiz6HM2uHhJMbzDkNDF5Y3oI3
N3q/7tqYZ6hKrYugTod2fjMO/MNpLTM3p5V6SSOQCH2O8wPJbZGDYwAdgtlorOI0MT0FTCbhsJLb
ThZA9Te7ECVnaf4RAPZyLwprx3B6T+tEFEc58zlsJ6TccT5ug4RmRgZtx7cb2wbIMRqlciqSFipN
cHk3QI05SD37Jj9K2MDmvnvGNWhhBYDt94R7kj2rbsPz8ynWWV9BWXji+2m77JQVLuuDnnhJkOmz
xffY/8tldP/N9I23QZ45VsPdQSvUqUU3Q8frPTm1oCqWm6Bhl+DfJh5D7umvjG/M5ags5GXKvhKt
Y7E/jTfpdDw2ZIou7/4cFyFRtTrfp3k+NY0JWZpCsSQeG1aSaF7xVZtpWq6uAKIn/KPAs4fbqUO6
AilfsW3ZcHK27KOeEvmKi5PTLxm0j0luMxAWvyPeLrt08C7G9k5uF4zHF/eeBWckjAwu1LQGdIfq
+imSN/PUUVTlsf8Ph3PuOSiSKD0teKa9ykuJX5DekN7n52Fl8VMESRJG+PomV1vz7HsmZlaNQ8qg
xs9VpdQRclBGEyDPWGJLdTgO2HpCWTFwwsA8WRrT0rOOJFLhe4KfKpjAqf8OoM5z+fC0MjcQWp2H
bBjvO+lbKUH2emEbvrOrH76XMo2/JSol2RvgFOdfdduNz4kO9P6nphpsovaL5g/aKAdoFZCLposz
PI0/kaF84+033s/WUHO6W2VqqexG8E+oKcQnYMVQTFswTgZa6Wu1mV+s9+RVPwGZWUZ7wQqd8e9N
2xgbVkfpMiHMVAvtz2b9FLewHnFX9Kjgx7rb289NTdWraEYGmUmz2Tgzl4b/R9G7oLWanHBilUGq
LqDrdbEm1cBF1MgKw1L/LaMo6P3O4MEZGMZfbv+vOSZClJ1Pr9SUTmjncAuJgL98Zr+0cxXwXBag
44eyT8G6OhL8VjzH37dz/CNjg5b8WzxxflReaLOYT5nM+RVcfF0oWelMKvs8gruB0pJSj7pR6MhG
vfyVuMaeyR1LDQu7YIbVkglHhEoazWiJP+ZhGPw8v+oE2uVCax47OAAEJK1x2vBPKjUr14TbfcFA
y2nAqjeZ5ZRMw4rCSiE6FdN9GNYFckPePfwI8Z45MZFF7VX6DBg2qlbMRsqNjflq2wOhv3OYJ4L1
hWLSczV//+dtcmrufDxRXShLpP3avDIj3gAKY3XR2iWF4JDZ4UAVDl8awDDs9QH4QPLafab9VWge
bxC3P9h15UrLZWWCIH82kay+rgMvKJ0MjmzMHBR91L713s3C0p0kOEGiVG/uC5oaRyTGuels0iOW
+2OCOkB2l5FPGkxuV4gUzd00eROK5aLzp72s43vkMbP6XkQbX+GLF1XYAXVmxIsxke6uTI7BJ+D5
BsAeH9iYA929AtT5JcLXa5b9P4F+oPNp7iJW91WbFbvuIxr+CxX4mBDVu+5cy5kaBd1fyMMDwYHQ
mINs7Ovlkpx3/kOk0bmm1nh3A882TWZ4LJRDoRoKIc/3pRTPCBJDBO2ghgMQY8Mo9walEEmTEQSL
wsSoMgBDUSDY2pnqyXLyLSAYY5KXmSIKLyNCqx6yS837hoMPvfQ49D/0lLHli+o5x/Ftsqd898Eq
E7xRsT/84t01AFRiQQW5j5aZ+Of7fsfFFDwVU2MC5wgEvDKAmvXlMHnm4HXNcyNd90yom3keMfmF
A6l5oqlNTiMRsFPfIzYV3yeM8f+HJvQzY0UA6KuJDq3kYI1RHqLxT4+XLSLFs35cMP3Sf54w0lCw
DwYtlhw3QnTCOAzRgixzyGwLEltIenGxr64yj6TZER33WsofGLY+aj5P9etyetqnDwKqlfU0A1vm
EjFRkpd3NPKYEq344N2EvgPx2zyL0tes8JXU/nLKoO5HrcV4kK0ey60F6tgfNIDvcja04r0BJf+y
KI7h4/QIMzDJBD5Bv4TubS06KXt1XOvMmeqS25pRLHET+LWWfkJxTk3vJLmULwQEKggxo+fjMBwp
q9eMZuoVHCdEYCaOyacLtBzFEppmMygU+JCLpvbXNaj8grO+xpGmNzSr3mE3WldduY+GK/Fkha1y
7SGSBdcychMlqaN3tEeEi3F2orOU7FJax2v3/QOahgrUG/246sdg6RzSbBgDuMUYLr9aBS+YR0s1
GbmSP+JxQvdDbycFiPoloC8gW3EqxA/Icj0GoA3VZVzccS7DDuH6cH5gmIADB4IzGzpt7UTY7Idx
AZsDNlcgUmAoyu7gA3vYIPvDD/1WPnwRl1hueziRaV9MtBAQSUeE+U1N0DQKRS4RfQ/zZGEsKt6u
WqpKMzn3BHYbew+tCioeNWr0KmdLoPbR3WsqcSbpXKj/QAMW8YNZEInyUcehIv04JHACGlfH4pJZ
0n39d0hgv6gHaNPyRF6orUzqoUz4ZRVW/Pl+Glec0JJqwK7dsNn46qiarhqeNStwn/hQWetppOlS
vhAKMHsgHGfwVQUCA4MRHRPLgovOn6wMQnIgOl9hBorCLdtYe4MKOY4fu4HufcB436HCyTVV8Bth
aEt1/n+NsyR997jmwPABes3wb4LTC/knwf5M62CDsem9FI6N89yLW4O/V+FHoI7IXoCTHEFjQHeS
/Ga84IddcUxHk4TSD5L6wu4nMyuuRzpw1i/pvMKB0ZRBS6VpiuUqpIBrFoby6Gt28+yW5BbJkQjc
mvZUHrzSTTbXFTOS/gOE9kPiPPBnj3oPPWvN+stylvpCt77rE9+tVgNhTTym9eTSkWzU4RCHPl/V
s+njZEOIavX4NE4whqA7lYdQT3XolkNfy2SX05EFJgooajzo72a4p0yxSV1l6ByP/qPX5QKm8cMO
sRCBIYZPM+9InpRWNQTXOUnOfH9FB1tcXMcuc+5iguu84ujholADgbc/wl++cvNv9olieun7Y2/J
E/zDQNVz5huMhCH56yD7p1dFoeRjzZ1Ord0j2ViF2x3biAqJ7vhq6o73iRPR7J9x9RX1W03bb3su
hhL2qTr2QkJANUMEn422oSy+lom7T0eJMyLt1HnPGH0UA67NE0WWGfV9/s1OqQlAkgiJhXMW89FG
eT3t10eTETOiOwRypKZgJmpMAmgbo8f7/uwzWvUNvLYV3ogRH9NqWLnRDseTkoHQXTw7MdYcove2
gNm/PTD5NhinNSXjRPng3/Uqbs1kj7Vo7iN0vPHtZrfVed3qpEwfCXGzsLskJFQ3uTPuYAWFAhem
26CWmjkbCMWGSletpG2bzl1zvZA0kZZwgw0l3IiFJqXTnetHqwWC0wszngfkYXEN5he+kO/cQAIV
3/BW8fg2D00iXMS5SSXbmoJ6P2RKgB7uMvOolPVA70NUDXcRLh831Aqup+pE2me/47headn4OeiQ
UH+qp3CQubGoL57vXZ7PDa3bjE14CQNGbWuoMMeNNvwEE7PnVMUQp6jsR+ydeofkOFbOcjnAjN/L
EnWLaZbNdGi26KLbWzwPTFV9Jj1nAod6REltI6dnAkxCtTHHbBjk0T/x8HWm1g/+yvfxnMkz+Ls1
KNkW6Q6k5/gwu9ehRMIgqzQMFpP0JzHS8av061bJQeOIyVdZFXcW4owkalOgSSZLCy8ZrgUjSOKn
2O7UpOZv3HhxQcGr5XUzO/oDSeB+/SY60ITnoJZHxPhueNKWBNjwMJmUWo6yatPHby6TIETkPcBj
MDSL5WRJh+kOwCQhtAwo36D/s0C4GNT2Mt7hvdSIucm2iW/JjnJeCk9vJTVIrfX8TycoGWjaxW4I
lOpoqy5Evqb48cUooMZvHlUGDlF19JZFf3umH8hb/EXRsr/lhPU0qWRmsPJMNQ0Tqnh+O+2VVCnV
Q/qIWsoF/rzoX/BQKGJEYNcdyTuGiq/cb4FpkM2XwR64FWx5pkrm2h2WHoa50A0haoO2jSKjpQOL
JS+N+g5Kt7YMBU6Nfi+87TuJr7yNYzBtW9Z+odaR2WTYMMx3u7pKYj3k0vb5Sq2qG5sMmHoGI4bY
XApsL+9uPjS+uCo5VQ69TKJAIMZJQbKORw/azMlHtm/p5nt2+krh4y90fT4NDwIuGrd48NRz517g
C1s2lzto5MR5tZZHVEn67U6Gyy6NEpEhfC7XjN9j7ctE3v0Qqc2xG/vPGx3BMdEcBI1/0OshIrIG
65L9YXKf+4DTjTPZ2A61343HuGts0O4Z0r16QbFCikFrJIFSsxBUK00mj3zYA2pVg0Fma1PzJkPG
sQBMS78x4y0IvGojliaYFWUuJNm2kKM32XMQ6q/jDu37haBUD/jsfUN2kywf20SNnXNNcV7HWwu1
5Iw/uIdL6XQc3e7paoUOKFLgsN166X/W0vnaUIIKvvDHrj2cQU7dFXfk2Fx5NEBxsLu6utABAUwV
r4zDVm7YP0FfKV3YgQAXoX3/UfknePrL9+y89UY87k0i3DcZWxEYkWu9xp8IXYP2g9dHTKM5VkJg
LDocM+9h1ReAt8ySJ8ghzZgK8wQ0e+KGTuahRkdk7aR2kFwk/o1nlq2wIhHcYcs+IpfgZ31pa0/Y
TAYlhOsjAKVnTd7fVd3uZJCMcN2VrSuYg2nx8jFsPp0xrolkTjzuL8QuOG2va+7PeyplpKuOk+wX
HjsCfW5m1iYptGcLLtw/93AWIw+0fUj8hZ0zBJaWb5MiqfSamX1Xm0BcFFfz1uOcyDI581esIUiT
mgxy3d3oQuNbf2n1wHr8A3c/LVcU02NV0YA2A6sMm1/R1Ml+QWTg2mryVzVIYFkC7x/yBqJmwRQs
0QAndWRNBWXbk7lpVWAcPWjNM9nxD0GTGGeesJ5XTLJvrQnaYOWqcOjHhSf9NLganOrTU6hRo4Qg
JCncrXtqby9YFzEzxATQblIVrq2SoThLtxSdgEV8do+GAUDmNtWo8cTTB22Msc75iz3xaf7C/ch4
eRygBTX5DdR6FeUBSAr3/Mr+NddLdc0a/gFYKQQDBCnPaCg8lNviIpHF9Ov7QbUa0IXl/3eJ+gCJ
vUh9IivMgrgEwBHdOjXxtGQqm1i3tKL9SryDsRiQ+GUkpPQ/M91tgHFWROefolujZRzLrEMKJxsr
X+vD46ijki+oGO+cXRYkY0qrE0c5Id4b4I8YNdzjBbZ4oDc7XNrKvq6FV7SMMOXBRCNvxGJsSQlO
PCAWPSscJhYynH+qsDp+lovBxxzdCwKGQupkaAdi8oqwliOtSiDDuQ0T4xhXikhlOeHoGBx0MQ8C
FYMrmJe788ugygo+g2ttY1DvvEWt2wQx4feU2I7uDFoEP098Rc/okMKwdRi9c9xHSFBXRqjh1rgI
1Q+Gxx6jtLxdaT1COoETOwKb5tMwjEmfxWNoCceTiOUvvR27LfzYYgdBzetvl22tbsFxnquxb3rb
Tq/ZMYVSDOzE3P3S6sEG64zbAV05B1G+luJEaotDdlVBH8gVvqaIBJVmq6nHP9SqiftXEOnpX+h2
1Pe35Wwz/SfgXa47v/oPmEtWQ667frr19jxEAc+Es9B76yNuV7uPkoiSeX1FZLMm/Zp35reknyM/
ixSjUEB4aWRB+LP+QK/dJ+lOzCFpE4vMwMdzDzGcYpy0rQ+ytO3U4lKrXkJxjtLNTYBU8CWPWwta
Kf81ykmdQ1slwxzK42sMJH28Rdjmkon3UdQ8BNB6LSlVhKTqy2xFQAsdSV5PUFbwU8h53AHj09wf
W/RKmXfbznzHtfR2aUyseEL9ap2YXtObEbb4DH2PRK1fwvD7b+OCwLa2QbUliiwtVgVFsdW5SE1M
JqlTgtULBXEzZ948XgM4K5/MPd36y5iUNt+b4JLZRht8nVeiqLr/bYCqwRiESlqQfINqosVUzZKo
kBCN2x3qW4dnNENfN08wO9a7zN18/9rlgCciYvDkiRB3anoWfErpoTVzXty/g6Hq4QFx7zbmiHog
+7VU3PxrA3bt1MkQPjf6dJzl1KMQ182K4aN5nfkIzqoriUt+KE4OWzhvz2cOyM3/jx+8xfvfe+TC
xtYTKpikrUgYwF6poAN7KBKIqcBLGoS7xuEDwbYQu6KI1byiiFeVw578lU0Hx1dIxqxdA406IhY5
fY30gxfzJtPMVSfarDWVRaJ6yBseB0fDOotXxF3zrysCZHDpcWyh7fw7eRFeyOnao/E98MMcL9aS
TeQLfbqt2t4li8KPCJ1vHNDm7zBdtgEtmgmp1vufiu5Dkgt/Y+T8g0gZQjnc2fXu7L6j8065lNpZ
5eWvy1PgWQiMgbPD1VdLlCuRRiSwJkdKE6+I/kAr4o8aHGkiyitTHdFybjix8sxL2RA0nyWgVt+a
XrrYRCmvx6/QiYBjQ6MygqlNIEnJkboruyXtD8j2kP1b7gCDVk5T0Fm8K5XxiYY4zlyBcUe71pel
+yIGAd/8G6JWAORZ8rzshxgF41291T5Ti0ri8CMQZ2ybvvm97W83x/ZebKE6QhjJ08azprQEpvpd
5CNnC117KicIo1qheHbGzS02uOTEuLLM0Rz1vWMuTJ0FnAuv3baaf7UUSJCDr7josWOkmaRn82PR
e5JOUuEJcWR5XkRUTe+FdCu3LdcjcCK/2LWt0XiBr1MXIRwxjw3PQgq9yUmaElwnxbomQEhft91t
vZwQ/XNhyz0ttIjzMdRR1ztkglwNS83s+D+zlwlaEQLXzfyf1zhBdlAJHizcMxqNv5ONX4pmsqC9
0NSMRJm9YSWjcjHQ+9kwd0de5AtsehTG3YeUanR67ibLrODdMcFinVntTFmkUzErtgnGapiRcl77
g5OtrrB9jccZIjOX0QTWq1BAJrX/wAgj1Z9S+FzxukTTX62rAUNbvhvBuAQscIaSaKLXPvWJPtBU
8mdvOlPjWbaX/teBa5MiGb6+U0TELNVwNt+4jLnGzs+L9HvmtWeCyuobE4vQLNwPySsTR5AMB+Uj
gE/yzOS2qD2/q+G3jAwnwKYSF0YJGyhuEfjfdd8CScVeooypp3nc0lK4C2eh8rY8Wqg7XE/QtTdk
DaegRQQtcIdP+t0Vyr1YTVKaB8Ri/gsftwG29Ivvv9HPwB3YxKe+3x8ddxBo+OjA7IbCUdsjUkH2
ZdEGW5YBFPSLiZn45N0NrFuDztlYM5JmJdo3wJzVQdG9fAFQbZLIcMEF1Emm3qZ6XB9NElsrGl0b
pzyb0UFnG2TrVeRv1QplhSEvEPAyiuMEuuz7VfFr7emFKWLg7yp8A1Mh1Fg1uujpA9nFh4f3xPFS
7Xk9k99LEc3UEgPEygVWkB+nDAY6rWd/4OpX/2ChLQ8C3Ed2BhGtGnPmuCLlswsG7G0TSVoytpBe
8bvjrLqZee0buVHdlzR1vwo0CdqYFOmsfVlMUWL3k0mX1XFy+2lamZXui4SlR+QgXSrjpg+PNclU
TN3+dmZ7NB9gaBOjTCcTLwMO4I2az6jQscy+tWg2Xq+qXQdSEhcmEStCTEQcIutLjfCnSls9jpxy
HC1OM9bVXysJRkuZpO4CKUT538CbkXHosDcthwNznqEPjy8ETpOs1ftBFDibAHLFCp1YBNItfIAt
bRz/h2NUXFY6MZX8J32uXbJaxGJFcIicl0K3jxUGNN/aqwrQMxvv8muXS+SXfHfP+4qHyMVoCczO
fhmOeYQ6IVIPpLEllyERFuvOuYV8+AWAZXHAJuPkeSEhVIcX/z002zUi8uboEfSq0RqCosModXc5
zo4IpQe31M5s3AFeLA2GnBDZuQtX3d7qePN9QBIxhi1FL15N80umkP47jXgIIju7D1Qmv/L67uBq
fAgK+t9cgPLuI9zBou/s5LNFwQ76HGqCz7m6WwsjN6dp/kTp4NvITyDUjrQsV6rZzqLUGPYxHFpF
wTDcVQskBQjzFNt9+wG79CPCU25Me0pLeOj1XEcPI5xIplH94EUCkuk+/Q7Z5HfXZUD4g6xntkOz
6/kIIrLd/8YVtNgEKyxnqNdteUL5fLzmIxMloLIYChU2q9yQ7WN7/XW9yvyjXH75GGAuzBywFQIl
v9AW2cUUSIcLUeVrF8rvBMI+3bN52LZ0JIf0vOVzvW4bcPM69Uj5k1b6VEaZLXQd+0sTxgGSnhJp
IX2IxKadwjLccHiM9TH1ugEVHzu2FKPqLeRha719sMnr0h0wQSbDvsBuyVmWjh5AF8pO0JJiGyPM
rbpMUUYRs2t1cZ0p6H9OJ1xVUnzB7hY5EYNrjO0neM074204YO1YCxiM/81KFCjoV4TbHCWKWvPh
aGfLViRRL+xasBx1Xcrx2nc0UK3Tj8ucBFOAkCICLaKvmkgzIY6TFxR8BWp4CyA6GUjTsWNgICR3
Ybya4PxArLBHY1EIG1f2etlBkcXAEkYGyNwTCASlnIaqLoraGkfejqKU+Jbiq6rYXT5wjr4sKvOu
qh/cqT/du9e3TT1pFipReAtloahO6fVRMKv62e75/tuI8/JiLfyldXTN6+VHRoRWTpn/j4e5TqM/
mvMf8ic2agvpSRm+S17kWyJCb52Kw1SwXiGhvbm6Lex65BcLuOOErGTqruIjq+CcuNS5K2Aci8Di
XJU5hrL23vBPYqYVHrkgReB1AXtRb7HpOmTxh5GRuxB7jax9laWyFoH+0iklwFFojOAVj9qMl5jP
P17tXJWtpJXgYHMJMQTq+fwDsWd5lpOiGDjPxpYb8NWLJy0XWPXlX5iB7/ru6p68gJHG/s6naSg4
4aZKSTd6Fa2qTJeT1CmK9Sco2wvpw2tWgX8ytRDwSuxJtYV8+0j0eDgZmjsdoGQBOgM7JPkI50/P
psMS26iImcYCGw0qNHlnVIMP54S47xHDN28tB4cijW5n4cVjQhD1tc5xuj8GGWu5hyabWvS1QAlU
7SlNNgqFEFFxMtbY1Z9jQs0Tzz7dfqiZqGqDyCF7oIz2ScNWvqbOjBAn1lY3X3Ihrnj9NJ0y3JbH
bp3OYEXEaGL8gClZn73R/mUShGFboJ9v40H90XoLgGykfzTr3kGDTPqox+Dp05qxm15mbOjIkLMi
d5RZ4uPsTRbB9iMnJiC+Ni1CGCXKr6nqw/hCWxwUwY6btcDxt6yEi3ylP5q2DRHKl9WySYnl9ecL
EwHy7SxZ+MiN540DAv7mMnYl5weEFjXlJuUZmzy1a9OE9dspoKh7+chjKNl6oZSpezBud2fxUC+n
ltV7y2tZIaDNT1a0wbbLG3epo9mIpBjtxR8hBZKOB+ZTvov05O0COi2kAAFCztoWBty0Nuk6Y8MI
x7zP7FVrIot9PC9u7bZUIj4XDxn2swMntATuiKE3bW4YkCFxbqMkyJlKm9536dGt079Os2sxzxBA
vCI6DaWb3nHuaXohBJeiPnSdOO0a2qsH1sXvDyhJSYB8Fk58M9LE//DZU9ZcmAfPc0JcnYOkpW7b
6SPHxpmsU9JfjNDhxh6uw1oejmQq57d16SLYTENqbJq6QiM0n8vslo9mBACSE8JN56UlgaX/m01C
qKLrT8nM8O+yRBzZGu1UyPAcCRffnIjf18bq2/sH2Nz0GXsJLJii8B9eSsm059uTuktcYcKrmMFa
F2wKyFR7kZ2Z2O/56+7ci/E/R8pi/n+74o4PNDwtdCpzgA5N37uYyJT8e+hnFVWI1RWtCrhMuMrS
308gpIJbpjuWZVQVvCPgHRj/cJiQfdTIIPzO5JrirZhHnqb6DFiiCktl19hoVchmjlIaohTFdGE+
qKZrjFhPC2ZBxPBOLyoIIM4q+0jItjEJLUhOGcn5f4r5vZVfereaj3+b8bLjOYqYm+en6MmOAeL4
293xlwKC5rCNwM9cq6yftuPFczyGiFr2/DcOmWgKV77ww51LQKb1OTuX8HH/2MIX+wEq2UV+IF8j
+IL9zLvdojazxBvzXDHNL2uHIwWsm/HW0bnY48th40niLj/7Ij8Mj2KgHKcPB1M24ZA0DYg4vrNE
EJqp5U40x+DujIvhLSm9GFs9ebM9UpIlj+kQ1PiZFp7B/weH3sUVzf8zXuvYdngrTY6vyLUv7Vpu
Rt7RE+w+ExS7Bp1NFnMBDZ2eqCbH7ywm4VVdrUV8Pty4lruPymhGH0OFh+9bnE2j4CyXRRPy7VCz
E7AS5NMqsZEW6fhSn87e3hpDC4D/EkAObN1Rt5l9qIxFuhr8m/Yhzu/5FtVkZdF+fFi72HXO24aI
mKPI2VPHWs4Jwn99E3wo3a6+S7kXtxKhjxwEqxq9oB6O2dWWOKW2j8k4xcmtN4bR/E2moWDvwRub
MfZOOe1IzwU3vtJVAobtZiIRMhEPObAkFWsuWuJmRBhHK3SApixt0WwV6J6E0kvakvQXgwbnosVH
ZIMykwN0P8VMz8gJHfkFx7mVryJpGq5geT+IDAwfK54FGGZPIR0/NYHDwkZ3Q2M+xInLh0fiVI9K
drNLZhUHj1598F42M57Jx/i3NH0qWZL6WQsPoDw8yITlDGxc4e4yWgIhPPnN9LJYCjo9/fKGHhLa
RPOccEg6zwsJsdhblM1OXa2yFeNrJEkbNcsjuz2Pw8aIYYahf7DAd6G1+4RRGPX3l54IVNRLcPg9
9LsEFFJxqBQIJIsIyxjwu8rEjE8raStc2Zfi7p5ieq5LAbSx20OOCYWSWQFBByKQTCv95uHmX/BV
28JZDfwJfpbZ3vA4ecvMEA5rLH/FOzAk+/xpbimcRF91HvOfoq97aqbTFQtMvPWxoKgNTcv2nyFs
yRRTx0umdznPDo/mEiaMqAW8AIOUok1xHuPO8oBqht3AdofUoIwtoNT4pSyvGhYQuUcaZoFXC2yG
9KL2Ix9oJgBnfhgZOW00IB0Yy5CvdEiI3tkGoOKX4B0wKoiNd+5ciCQqbij9cXVh8bwAty5Fr5/G
vN/GLy0iJ2qYZMLzi+CdcaVgv9X0f09WQCfYv4c4Gobw0YPMAHCWnnD/ZPZ+JQUH3u6uqIVD4dar
fXDYkM9zpSicEaDh5svEe3QmFGEW16GA4RD2b3o5gFBiM+jJy/zp/UCRJJMLY7aUrBPgWge5BTi4
DA7LkkGIPIAustHBXv44t9dvmbysVz7ZYgnZuR/gtanQdV1/NI0JGAYCzD0Ma6lkVLQWDiPVmMgJ
B8kG+6pTpHgZCo++GEpo5OzZf3V60e9hi+v4ln0VS5xpHPBSk8xU+NMCJi0byPTQPNxzO/XXvxHn
+k/3XVbO9sPBb9Z4yUjY3VQ6rVDF//iu3GQP6Ooo3NNhxEo3eivhAo9LrxvbqRfNXE1Pc9pWqkVI
y9OYSu7lxWBeGRYeDKXFO2i71/oiFFHWSOcYtU811kA8cAqjkgcHp2Bax8IcWNb+4Rjs8f89gKJf
vUQj2PweDQRei+Tl99jEHn+wNs2J6yJ/3DBz8deJlJ//peNTWDtgLknMql7oswyfUTsI8dwe6bmL
kkxrOZh3W9NxcJ+SXaeA7H7bMtJBMFuk90QwcD66iKaHsZ5RoXmTlQxLb1I3yTOxajqKyJHBuxKd
Gh0uEarvE56wyr1s4NdYHgnwLv9qu1B3mK+rXX6kBojpoWNs4BmCYNQIve0hZwUxTXEcz//ocec6
9t1MamBRzILxqvfwvA8hGAPXHvDanZS6bNDsjO5EJiDCWUwV1dQabXPFvPO4Bz+R0itePHkRFhrQ
cD+W2EhzOTbd9MbGybkRvHEUG9aO8dvOHkIKmWMAZhnITN2lznJPiF2bIuVZvxSWOTRn0Ts5iAcD
estTr/O1UOHtmeSQ2agzqjzCoSAGaJ4etNySi/eJpjVW5SCU4TCabTHn5TTrOD8VKG/5sXK2nGaY
sWjBUxmH3gmOuy0Jly2W1vtUUmHf/jEupgFhhs/6phQ9hF6ROEz1W4uot3y1jNaYcV7RZYiwXvad
rqaUXx9P8jUrOZxs76I5imPM3GuhhybcGVJ+fqsdxeamd2TtgMUzstwRYFlTfQfYFaOAr06WJkvz
3oaWnmTNQGjTqs2yHj0uzwyDuKN+e0DsAysIq6PIKdq2BTrcI0teMRV16XRSBNaM7k3HWBtBUxG2
K+jpcPD/SnEqDuPST9+i1PFncJbrdA9Z3NtraNQ6Kg/5gwdfrlPe2EwFVrHwnILIGdg/tDkAQVBL
CIqPEquohSWYonxY9rk1+a00QjeA2Gmv2Zj6mOVTvEzXpgLvsW3+eZcFUSK//IADkixkB3g6f7gL
graah94jKMCMJfMGFy69wP33lc5Z2z/cvKPfj+k241doGh8moiCbJEGJMNN6W5AHpFuhS1Z3N5Lh
nTC70SOJaDt0Uft9+4p7i+NoF9ClZLXVF1Xk27vNlLKB+5X2lt8EF52Er3kZuIc7qFPVLZYQUEnq
1RDE1XI4V+RQQX5AZ2a+Jqej0tWscCesqSa6n9AMoqzFHd+FD4IYnFvSyuxo5VGf9GfqQsGDcnTz
CYyOLdJnEMZ0LgSTN2KIgkCDxJ9kQkZgvmhlyVe0AFlA2zDp8kOS4d+RmavKxpfA1++YSEeQPhDa
nI/hbbcj6x0lfRC6T132BOo+o971NTgtTN6iOUjry5K8hhY7LNaWZlnOzGET5qanV1OoMxQ4UDFc
2uoF9dADVlqMtIjo2l6/G7ZKnosDnPz9NdNPGIoZCN6Ht9uuPh4hcHM6JIt2iasue9zyckqf54CT
H/+MKPqqK+6Wsmslb/CidmfNnwy89OfVU1ArYM7evuQt/Jt96MM+CwdKrwraj1AeNvyvhzj+mXkn
EHwsPoOGI7dipmCYIPj+u1HRBJII5RSGIFtQz4SyaVPBWzXcnSnoKxJUsA18iZHUf2PHyPTgdvFJ
fioAX2n4hQPmdb9bJVN2X9EZ8srE+Gy15+F7fny7vi0tA6deh95v6ROoM6cdyVn+f7vh2BWfTm1T
K+X7VlDrT+Bou/eqY+OIMwQ8cn8fa0pw9mjXpxvSVj8BNIGhD4fj5A6Nicf3zsgdD3KL1dBzo1xi
TCU6+fyWJFz6oT4qOPo5lKner/ljZnVVW3NVdyIcBsRo5fi950s++lt4lz1BknAVgmvcaIkNdVHq
oflVmX1YqDKgeqGy5noE7uJ84xRfZl++ka8cIEy/wTY2y8fyJsV/gZTS6+gzrW+KPX9hi6EXCUY4
HPiY7lxOnMIa+wq/sqcW0Ruei85eYQIcaU83BnNfPsGSvJdr5C7UokQDYydAqU/Luq0PvrA9pJe8
DNMujZsNqdRThflanft+MMmZl+U1tsoV7dimq5uBHM1aWlKeR3qGYmaIio6Nla/NmesKhMwhDemx
ZaNpJ3EeJU1bNBYT19nYc0Z0r6Cr7v3rb+f5YveG6JVHFhGn21qYupdGJzb7zeXFgRj1QTi/00Jg
k9PcUw0Jb3O65VnKzEbkUOvy2rLE4z6qhoH2QRBOQhRGrOzwt2F+6IOOwh3gHeAmtaPP1VJZVn4G
5ZnK3dN90r0JtrEvntaVyZly9sBoGZCFEj2xD4ocPHqZdXUbd+NZX7QKuRq2tWuFYuPdkXgeSNPR
5Rf+pl57Du7ZVjvCixIvWW1BlNEk0AXTLUIgSj6mk+zlMmydsWKfaAjwMqPqs4OnoMHgvThIR8zt
glyu24mdkFuOgoql3rS0B+ZyY2+7UkHY2FTCW+mmI8SJrvD8xHHhk1OuI6Psizi6sbANOq2m3s64
3wQ54FIxDO1nRI730PRj2NlHGUduj5+lCB9uqAU10QV2mEm/eam6wFYMs97brgzMppC+J18cpKDM
mwKFh97h8UUqeX9MUJYlaFc15aGMaSpSyKqjuSv6qclafKzgPPRWZziy57kU6ige8gb/pyYZmO5l
3t35Z53Dq/uuEwUwGjoGQoxeJoKeRt0SqgLIgMsbNtnkBxvzHrEcHiSUf4EIJXBUyfv5N9/1/ZRN
jVrUiaNZg150Td7eh4j5GskY+7arWIVmK0VacH3gGtsLwMfU0MqmAeKZEMoTLXCzbLomxCFDv1Hh
wevefm+0nm04mzGIeV8CkITZmrlHDaqTQ8bcXLu4bklciRmw/uptKPvNfZmFN/EqeScb/f86W2Wy
gm8n+pe4O3ffzPjrSXhyxnZ38dTrEwEQf5p4pQMdf//kAg062kr8Q+R27y8OTyJnNGXthGUurkDf
wJFr7Wufhbm89KfDjQcBbjcRFmJHoG2vpCGZSc2HcQQf+v+9JSjTOQ6hT9y0ql6s9E9/Up/kDUNu
FELIOyCycDcXYFAWR3PaghfZqAFovKaDQWf7N8Ncl+jDYzIho2CE/D++L7rW+nXzBV55Kj+2S0aH
XGA6BzI0rXe/YQCpn7X84ESmb/JA6UY7hE9Dl69chKiG7FfXyBJ5igNhnIgHhjevct1kaytyolFi
ok6f/K03sF5kE7U3I1+lMv98hmE3wEjM3HLFD5k32s4Eb4UG03e0mpZI1IZP3kr0+SMcYche7EYn
4orALA+M9YYCV59ytOotkEI0MgGgY6fOE8oRkTrO2b/xkOvQThc+kOVxQ5D9Z6NFLhVFJjA0Tq+G
5EI+CZTDVZAVQaokYcSEQZ4JIPNAv+gawYiE3LivA8RBQWJHf2dziahVvdeLvnVwa6w0hoJSFFmp
PkJxZfGzVtDnweFkJWsFx68J1Nf5pA48aZXEjdslZVS8i+1cAl/4zPnZgdWvUgMtu1H7oVNGB5qL
2hYOMMWiVBT/0V5vcM9wU7mfGER6mO71Ehj9+afQ8Z/VhX1I3TeJnjEExonVWyoS80AQNLeNw3bY
pdDJ/Wzf9xLU5/RLGG2Lr9fJBCamr558iopB1V/MOXNsqwe+p2Zf9BWT1Dl80lT0bL4HxZE45da0
xb/TE4uJZustW5lz+fMGNWDdud99+phPiYKzuDkraP9W4fE+Dm8pXbLfzFVBxmA3xoD3NnK7i3bW
7GiFTfn+JM1PnjxtuKxGCnLtu5lJ9InAn6P4lO2OiZ+QdRfTN83BuV25mx+UXXEnNn3/PkeEsXzO
oQePQSWn6/nct9j2a/9Fg/vKlzBmuQEzCPK1aCE2EI47okKJxzMjUOs4N0dHut0vlNIHrpdUZaBt
xxKhM0kkIRwIbBfFJSf/kvMtqvsCy79B06kSco1Ivo3433dP5gPZl8kZ0esFLKFu/ggzpYrCsmHY
tjBN7kY1xY6/vGyNH98Hxzbnkt5CeT6O9G0nt8QB5kj7HCRCx4vNg/CpaemJnmsoBbTT+bf/MspM
wW5N4aH1XuLKV5eaGPVp5XiCDU8mxWj7fxlClUiyQPYC+P2EHp70olVxuK9GafPAzUp/mvZaf/vt
Ep0tMz8MOCt7F7gr01POeH2viogmuEZ9083T0z0NOvd2Ic9agjCMv2aTaHzIyfG85NucKv7beTTn
7/WoA2IllaPbRQijsFYB6zvv3NKwhGTCyP1N7wOIsGcxzkh5i2EMhDU26WA1KazGHg9qUjz8IKqa
G10Q663/hcB5ojMYZZdz4pUfgr7JuiPKYQtY56ScAB8WcO+ODZzfPKSaU44s6JS7hTe7ECAYh+Oc
/1Bl6T2fpawzqq8f0hqsIknVF8swpLJqP5oY8Rf3C1mjkvNvspfIh8BZd0EFYe6oeia06UwtuQw6
C5JRq4GCkw+MtDggMHmNsIFEruIMQg7EOO+Fkx38bQKDWJvzCH1beaiaTI4Z1vj12bUOL/WO+ugP
fAp0IVwUC+lbez2kd8UNc4g+seCMBxCQ7lIx9Igl/tKMRL41W2PFMvLu9+VlSKoj2KqZ17eJoH7/
pJ845UF1GXCxPhsHssozeoCdVeZKB9MJy64h+cai8b37YF1EXVMWoHrBjt/9vdDRytZnlj1q1Zh2
kLx9uvrOhIESZdZkvBGq+A7/Iu3vdd6NeI/qtnqP7dTvwGg9+llAThIF3msowofczpgR9Ic2qH9R
n+5nGt/Xw/cOXXo48IOXO7ThFJK+8j6r5woHfSGhWseaabQgmj8LYsVdXfUFIp1DY+rfOByGT5fl
VAJrupgHX2JUMx4pPFZgmPQK8tOg8oBcL7EGE2Z/GVEV98ODCGONV73DZ81WLP7pL3S+Z2TLHdRa
prO+WXrdy86+hSJiAU2yjV+7KZOWTk+ZsT2yIUpZ2aaM7D1soIR4NQuu+Ww6Vq8fbH1tdJdPDPMh
BC8FO/KGGhpvpazz6dwmjOJumIbaUtsOT4MjBeHv0zZ//3Qm6IuCS6QQgOXLMQo72UsjoGwyf7l7
5ULOVS2+Y3s43GxfkaZRQwXuY/OpRKZtfQYvME2g+kbNm3ZDgUfZdyWTAR4s5sBSmK8W7Dxu3tdN
LvQeccr+EywsJUxK3Mn94c1QnMhSqrC8NaUjDqaBQzwkpYmxTLmmehMGbBXUQO7myB7GUlQFybFg
n0fo9rAN20DvfB9AvNY0K2fDGpFh/5nYSkhsFwVve6eaHSSd/S4YCof1694M4JUaaekxL1vwsefO
T5/Iy9s25iWV4PlrjoSpKoZuDWm0MbFIztHR7H9M7NOPSYFKdr4b7pt3K5NRP5SaWdaSQ0iUhs0y
14jYARKElc70loo1P1QVVEoO14jHwkqqNcTsdPoumhU/DmWxnDB1V9cHMauzQPyoWaJ7iNqY88ZO
fkUnZdLhwNtItOfGkYBom6zVlRkqWNzyx3mVG/4kBE/eNfyqEXObineX8x6pikES8m7DtY1BEv1W
P/9HF0Ob8vFG/bo4Nd51xPc4f2pf0REdEIc+EJrYDl6BtFke4WmzjYSAO0PcpBVOrnY+Jtq2TQ6t
6GnmYCaE7TlWxfozLkBrGVCxqFIqR95jLPknZ/yxLI5eW4C5fuV0n1nx1RqrmtYw7WG0b8LJP5el
EhSaBql94eLtSBG/HyPU2u5YnOWf8Kl1U61wYv1d4CJvGEiuZmw6NjsllCfodn+YWfmEwwBUwQRi
jfOmGkBt1DctLndUMJavDR+Hi4Vl4Nke+zG+3kSj919TT/nWfpu55ePT7+hg10BPpd90mjOJX9dQ
nf0upTd5u+pO2cU3f61fU/xG/+dNgTGB6B1p1iGTmDsubGqipMvcMw61xaVQYOAqAB6eLFJ4MLiU
Y9OXCkX4liqpMu+gO7ttlsarylbJpnv0WqhL1C/JkH70f8BiRnWpf6pwo570R21cowU+TIdhgl4T
lBOuy1hVs4qWKedDwLughpYzZMiTswwfaYiwtiKmgF7G8hU33WtK9x/nsgk+AwTHPeq/U3pH6+hB
QZnQnQ7eusknQiX8BLcKvJHYn3PBGG4guHxFxFskIpw/CLufqEaSMt6DLQfg/eKrC48swOidtSBb
kuhqIIgKj2u5JrUJrFbugKxD/OeI/Fh82LN4DgaR0io1MJ9MIUhs4u7Ol3KfPGK17RvKpsbvjR8O
O4yCeLcsn+P1xO4J844ytrNCK3UMFt8aHku8hYn1lsyaWmAsrvCJPT4aZQfjEzLhPp92fChGZJZo
NFeerPI3TZFWZEf1FCxMh124k+E9lwP2NDTRdo/7CQKtunQWKKG2+4NlaIAJH8eOnbsizAcOS7Xe
f1yr7MAiG9/S2dtFcKhE58GC7YFAaPNHunFP+1E4CsGF5LEbTbc3Gc273YcN4zYYfvqJCKgXH+qa
umUwVx4OXSEyK+tHPufNI5mkggW2nSpXw25R1iS/NkTfM0Sgl4g64TWK88oICtYsCF0w5tLU52pB
XX6m+Xb4IpbtqkZ5RJhHhiFIzeYvjNVeswTTFrOZZFoWSTeXtLWhfWo1l/6BG668+xW0iQO+w1yr
IUBFuXONnCz0rLx9lT93PPU/ezLxo5THxLuYk9tKkcpU1/9DS6w/Hw35SrCIDCVY2MTMYodT27ne
udbdltUsv+6bhSbVkv3onlLkGElqykha7jLPakhA1yfR2fkU/Nsubr8Vufmq+EYoZfeQMomDo2FJ
e4wa+GU7VT2euzFtGYJzkAW2gW4LDuYzkQniBJmVEpG59ZCa6u+L+ziBj6V3xW2T6e+2trwKeQWj
cvDdXICLef/GYGoZWwI9PiU6p8C0K/mB3RDd6hiosEv1UVD/TFrFfWNaockFJmnMXal7/BsYQ/Ve
1Kj8TubAxC5G1UYU6rPffHCug11wBFUiJKnKG1Gu1nWOR6HlVnkGQRxbkJdju96+kgCUQGiwn+2z
YIkVNhjR9NJVUUxG8Ta20bMsXjzqmTtex8/yBqCcdNFHlHcC+LaLZzptyWNR+5S0QGDc+rQk2fCO
MfMrN7hVdheRER1DndOI29owtXOAVOraqpe0gbVJGFwQXBURMnCJSf0GbyMsNgFUmVSoimv832me
Edl7DEh33NHfpiyg4+93Dzgw3VtiMnClJFe2adD+gP1LrqZOwItTUIXJ6pnAQHx766H3F2eU4bYJ
637aGv/szCxKk3go3LQehLKFndlNrOny/uZuHFK9vXH01O7UcDLvGfQW2UB/SWSOkAzSbSfqMCFS
MtQokMTDoY4OJjEONlFJPMsVO2OSc9XcPqC5lVHvlsEcVOToWgFsY4NSzG07Hn17If0qs7cdAj7I
kxVsS/XhWpoPEazodHTdJ4jlvFEM7qfGhuTU9plKlEtEbZIQ6iCvlOUabQI+xzDfFggGg5nApuFn
eFi69vy2Kq02OLGyqmnwm/LOxyCWiUPjrAzq5Dc0VKytCcFcLm4FJJibdq/1hTOFPZADY7fUXZ7z
rnr1qzvM5yhXEUN0Aj1p2C4zDsTEW1d2tyHrZ5KMMm9nkDAuMuku8PdfkSm9Bz0+itNfzZ8430Yt
CBQ0QFSOuIbTm64i6phDKFisGe3YKXtIBIcW+U2W4manMoGenjqxOvITj1JeglZGXUnuUuEAeYgW
/qZHIDoKZXyHzUV5LU01Ux3wv/uG4mN0NBD/MFJQbSjv5aqzXL9x4DpWS4ytbFg/PKlYlKoqXX7q
MUhOYTgAy2C7kB4dVUg37zH2IftoqbYWqOcgXevSEN5F6fzHbi3vFNuFPvgLAliS/cORfztlDQBJ
77QDcrHhzjOAVVP2KaNAI2c341/+LGMy/fbYyYdAgEc11QRMMvOvHK9MW+FPTg8tE9pL3pWtMmsg
4Szdce/SyQVPherMeVNV7uhZDsaWwGKmUw0RCc894XsjdFRf+ycQlnYN6My8f5HpKH49U2zoAlFb
W6sROKRCYcZVttuO0BlmuXGVbKtsmOcspuiy+9QYjpcsvk7+DA36+WMezgIDMfykxVjglOCMFksK
Qr7qanbHzjgystUx3w7DHZ/F+cTHRf+tYDM2+cxZPCPSYDb1VNIvXEul8yhI5TWwXUa5SiOQORzG
uznVGCAOSQkWhi/ZG/LoOqKEmeIr9PF+BoKLyg85IPY9QZqEoSQ+yzj+JpsOIeTek2w/xR7CGB5R
lmOiMSzVIOE0J+oOoz/c5OkLcBrrLoNcIweEN7V8oikhLS0XHMSyeLdequQl1vWUepLg44GJc/9L
T7CQHUNXGVw5k919ytbFsLoeaxs2qmdFo2NCHT40FSTgx/sSVcEDK7HX07wiO8auUFaD876ZqysZ
7TADsQSo9mjPukmtcWl/067NfnvaPuKnn+YT/zVgBXyxrxNn38hiLuuXTt2EisvRxUbC511C4fbD
Z5tS9MrDUeu/q77BgjvV3XdGBMVP4biAN6DfpKb6V7KSfkHCrkeF7dQjk/TuOtSkn8O1P58R2m2w
fVvgpfIv9BUIGVw45Hy3ZbnFmhin4Aea0g4zTq6U1VTOfr0IiLYx18iHTzKxagfBKZmB/JEhb8t7
fXCPO0tGPg4P/YVb1SzQ6hoErlMGwFGeEpn/D4Ow3G9wsel6vY2LoONudAxb0xmc7uAuejLWnH5j
j8rohSBMQcqcxgfbG5Yx+UiEAMsNMX3+yOv33B8Xg7+DbR65VwTzjafeUpT8kjdBo/0mEvJ69LVa
419JrPD7TpbIfPeG9Uyw4Qf3sHXbf1ES66OG/ussCWeljaXmO5SdWbNKEGZoPQwaGZWEHC0eZHi9
lGef+wHp7DVgPUUnd75DKLNiRme/gQrN2jXI+lbOxg9RMxIvK1wm2/3YFShEDoEkyGLzKQLXbHp/
5LQ7uT+bG9abbhWTKyIP8Q7wZ9TKuHrQlFw+OTPD2xS8umVMPznkP0sJjH7esoKaEm6nwDwEd/4Q
hwVmycACdVruMQ/7453SIvy0aoOzIzRZzUdKgLrcbKg2KutPwGuDDHQcEP5maeCd7GLTmMaHTYjd
w1dW8HUN1e56b93JrlWteDSS4Vu6VoHH2wqLbr6nB1txnzCv7vcVMFGoywvGd4mW7QBd1dl7dPJq
ZFbG6YSZLP9yzbSdQCPror9dIXE9jBvtcQGTzw82dEMqXfaNQFKbnNHdPy8r5fPKKqAStGGa+MjA
/uD43EGlUNZLq8PzuXhAh3yamK2Qg8mpwJc3Izb6RF0lL+qT+MdBchkXeOgpVA9F3OqvoCFpBDmj
9vDzlfFp7cS1nhkL6M6r8XGfzBnYqYpRqIXWhsDrDX7FWEGsyoIRxx6bz6ejyOyByXEgoIAqpzZ6
6ehTVewAPmrkzZ2DvhdLnifNIuaagbQ17is9FvjSkMnAZKfscHyIon1WPl//la+J4De+2z4W+Z3E
MqhP7aCi72Kt6BRxQ6oFafpNmIT5jq5KX3A8UqMCIYZkoJn9eKueM0jsXbukszF6RM1vRIyqkoM0
hbSQdzQoACLXBM/a9nfS2BWsQlinNedU0/Qf7c8LSOP/yU+3Ao6ZP6DDEe0o75v/NDzK3e9GzwKb
sNO9MgRbbrOsmnJ6DHoa3s1K4zQPRWazaRJKzzea9C2ajW6+hBSpx8+I9FeKwpMn/sfUPbDtXaja
7Cpo84SNm9MicCqBujZG9eI7UcpXCJWZLd9rznvklZYMAw7ycFxBRKknPh1Ey9H1nk5encU+zY1K
TwH+E1X0QQAiW8D0iMRnXzsMjvfZMrHyJ6+oOv5a3RD6kDdywRmlvDvAF9VuLkKJAAlp5wPxH76s
qmjWj0wMDNMW4en/Uq4UES8BrCi+uIoQO+VhdjG5p9aYCwkSp7dZfYIlAPG4Cgv7gkvek2+6HI6J
aN8Sd4WtRP/Hs8HBfbi7natXMmxerojS/zB1rdjqTkxFE3GKcsF1ezmWWqKC8qD+uyVJUy0O9NU3
fNGqGHPJWfok30mdY8MzUiPuhJZ/A6Rlz3Ir8d0WMb5gNr1fAkyBtIvU1VthX3tegeNEuvG3YkSo
jq5ybdoc/Ue6/6Buc0zMCbRBiK54Wwe4YCmUm5PVX/YDvqvhysBG2mGyG0ZNbFuwBLHhuPJ6ekQ/
CeSiwciIi+t73t+aIX7ghjBmjBSeFoNpHCSYsbjQ1bv2ea+Q37AW4jU3jUZlPzLX/IoA5Sg70Lv3
QqcyymGftl4nANWM+7JPMgvFmAMOvSXwdgMv7wUYtS8A6frvp1mwkk5jSV8arVmdebWpQebYWCi8
qce7CbRU5oHDlpcLYhFT0SHYXPIDH0vxA1uFWmIw+8y2jTiTjhQIqwz3Qb5uG3lxxcbZ9OgXDsZR
EDrcROuYCiRVx5xNOjudaa50an2GLDer2iUX+Q0SGpeS9KDkqDdPlF30asLc8GSmBUWVPrjQYcVg
bQf95EyfbG3aVrh8vB7UyThoAJjtdtOXQtpEajwfCfCohu15AvdiE7P9z43tlILkmrK48/3Z3+tA
5MIzHsCFXqo6C1dxq0MshKOAr7ZXEd8fy0nWwPkfkBEuQGRnG6KcD+ewXqUYHhGI/2FNKoBVj5ui
n9US7JXM6WVrGKwAXHk/5HKdp46SBHA/cO34RmOJ6Jub7Cxi8aBvKFCqrSQFDQRP3fEGaY0mfHTQ
mGT9w81Eru2lEbB7ldXkNmN+P5sDDaQUn2U+jkTxYxhhYRBJqV94YYcKnpKRTG3bFwDUsQgHbLP+
L7EszgXJ4gHGhp672RY7+fAe9AQpbPiLV/qONhUUBKuYEnuSxBnKO6Pf4mFa+G/UjACHk0+ZRDTM
s1beXsBS2VBE5KY0P3ZXaEhYNPHgNtVasTwG4iN90u+BZumk4/jTiymG3n28pjKV/IYHdD5gw2O0
TjwcHHRzwjTwiGbX1RB32656uZDDRMc8TjPPZokrnKIfe9u6o9xtFoufjQIh5bEiOP3rlVjlGhPw
xDml0hA2z2NHzpwhhVmDAKBWF8lUBSXBLCrTbByIDcS6tXSd62zjQVBVrm1ijf3wKG/IE34vZjD1
0fBc6WCF0Rci9Rfx7bp3Xn8hBKjMg1/TgzA1k9UgYc4ORQSNd/RvtWK1rir0fuc85YuKHxeeMgeQ
sUifu5B5seXwJWOdZl+BplLnVgWLEg0GkbrbZmJcaP+tg8e5fsA8Sp4dQFUZSGRL2DtIRoQHH8Ln
RkxTyNngKdP4oPRF7VMEOSNzHRf6NidglSW9O6nhd/jtnTNSaaOtG4o7spEoI60hkhRiLqdNk5jU
BXDGAD6bVBsbHoqvUXmuyP0PoO432oxIq8zaRv/grx8+V8rK6bw+o++7N6QtocZQU6Yvtqj6rKhk
miTrJ8B/kyYQglxQrFPrppUjTbowusEGb2965Ogopr4C3LhkY7WgmGj4UymDKFIEz6WFxwtRt1DX
Vg1mZ+8OK46vShMV/GdQxNvaJ7xfGqNH2S9TVMx4cvcrrKuiLwiTnL/ZeIEAEMt2SIecJjyfmLPC
zMJUkWub8D45d2oVMh1LXbbzA7MA0bj+J249QfL4W1OdJjtR9Po0Vf3kZHFsHW3j1hF3/4MT/aSW
DrKMQOx4s9EpBoAA2vVqdFS9AO5bcB6lx5V+hGysvkY94F7fvtT2WdsfOOrgBXRlXvoYKyPllxtr
mKvUjBEULx9gbdqw1gQV75Mzzc/YMNUBTHcgmEvI7msEkt75P6T4h4W/GMY5qqdMW+zVcOwrqi/V
MA6AlR0uV33/4GYtnHHQ5jHyGRySV3xnVgf1QZfvgotW9iYRtstCU/lZWXUhVhBTt8fcpPNWlQva
VA753d2PbnuzkAFy9kMMvYahA4U2aZEOR+d+KF6i9y+g0aFzvQeNgXGlwK/X/plLUlrhoHAaEJTh
eAfH5fYlbd2EAGYPap7CwXL7WPhK0GKW8xW28Czf0FFB+XOptfl1JIcBWSIOLAyVAU1xFo3ZpEQK
u0jpKpHF+PTok3FI6+puuuI3swRu9cM1KrjJeAhT37fAT3VQH8eWyswbDp+XDaHaDz6x1sI5DT+e
mpE/bpVvkXSXc9UEIVvdKdaH+JjkzktazQsFsugZwtmf/TED5OkY/goYeljdVqjSA5ujsaqeRqXE
Q86hT0FL4WIb/garZw73KboXKavVuN1NLoWEIeoK/GKUIsUFLBPhUkXXj8tdkfQPy69QqByerk3j
Bhvmz4BsZOIuoARHLHF4zUJ5SEXNtoV9u8a0qcCa+0AU4OLMnZ77D26LGew4m0TW5T0dXYBftZ34
FeNZMeswzf8tLDEBWJ7JfVe4uflSwdBAXuGNdrCzXnXg/PhHU7RtO0uhOYT19UaTPv10PIvY/ch/
YaAs8iHHhJ7LCZQmQzcA4HSHfn/soM+61Bm8n8q5loLj6+9aXWjSIAbxF3x77bV8sdLFgKUSV7Op
L34ricDsse8F8bOGGmPqFzVBONYz10Odh2mHzujs3NF0/9UD1m23+7EsVHr9IDZMWo6IJD0bv4a1
sioXmKUmlUFKSN5VBr44PdLL+5kE8yYGUF2hbDwN9ovnkMgzGltdkpPvxde63/BbpArgLALkJZmP
jDXc2nhBa5X0JG8zb8PuSuueLKCfXeSgKnNo7eTHLjlxqunlHhdIV3IvLqQE4oitUk2MEtJuXcdY
KCszKkm/jZq9KHYMlyGRKfO3wBlNy+gfjYI7ADG9kHxPlgDQgRbNiFKCGhFju04CxVUuDFfxj87W
9juuTCDDyaVlXs1SGNzeMAWrs0MuMX3CPbqyMdZSnqt0lJMlakQ7jCZwMz8mG1+0dmdw7CwOBg9j
G8lhUYJwwGscwxRxRcrqlkCwLBpBrm6xeHAlqYmOncx3d+++tVX5ml9kX/vzpPcRhDS0jeftefDY
54k/xB3VdPyOKeNHOCRMH3VWufjR3YuOT0AHsRZ01Zt6dhZ/qWRnpiU0mdk24heZP0N1gasIMGQx
8tw0DxIZo057xGG0bPM37HoCowHOq+giTAS73Qg1JGRl553GssluCBXlxAQ8T9qnwpLQJ4b0HwHJ
Sfoy+Km05VTJPBcBQzzlkQYupy1BMfNwStmlF7FZfK+hPBUFOPpTOL8AQSzrr2TQLRiphP5VICrD
KrfbICckzYOpL/uFE/X7RUJxNcQ9SsbpazuIyCFWYeWRFkR3EKRq/CDwnCCjpARin4YADf+T7vry
cznN3+hSiLOEmSh1kM0XTXYiWvk8VmOzjFAY8PD0xfCAI4OaqCtKJiwsxPcUaxkpGF7+LEG84sAl
Uj3WX3iZLXO5nuB/iQ+HmLJt0MmYbtmawXgGL7vbmRnuUnQCMH1VqJp2ynAUszJUdtXD7XW0i1Hp
k/w0suVnWROpZQV2DAFdRPIbrw6J6j3vdcCUd+MbQQ2VHfrmBAmzIVpwE1U0Y0uDm1zoCSiAd+95
7DgyyfByDCADAwFI/Ma7yEPYKaPKmsfJphDUUYPpSdiFCYXQcyFfYLShOjhgr8p1BWP2ewh5jaZj
r1avnnw/LXecT0FN63RSosFrKDs1m//LHPe7AjPrtqBYhScMvvgJwCjfqUKkUT3jewdlPxxPISEV
kPOPmlrXxSISw6+xLQ/kuB4l40T2qC67CF5sT0OXyIZiiuopRcR6BcZv/NhBWracR4ZkKbPvq3MR
FTmmxMW6Md3Wwl5s0vzSTjJoo014oNazLVaVHEpa9Jqj5GUIMJFuktg3NiAKV+T6GKEo9O/0yAc3
GF3c2rjiV7qwBXqA3vUHWH5dncLId8AopIinhOtoI/8HaxqZQQhRquXdhDyznYCbZ7acBKYw7dX4
NagvU/hNKQggCY1MrCet7sIxDNq0A6IdDVm10MmYqkRQHkfAjge/dS6WGVe96zaoZZaH7B5byfoV
59m6boOkmqfMU97YaYwHsBCuMkeWJdcDTM++wuFesPKI0GwdWZbNjlUgk6u3EBeACV+OmwgPmvZK
8rUBhaeOO/+ly7Ri7r+2xvziI8ESj+30MnP+yVtFs2heBnPglTzQB4N//ziCmnKGz3J5kR1KMcss
MWz7kNO5ISUM+kn80KaCTtR0PBD4mVHbG4ZvKvne4KU+SQBLU55OC4g3bM+DQvVHVBI0MXhzv+KU
KJ2lpc0GGHOLG3RYvfBzvUlpFItT78HycIVpYtFuRdhna8c05gc5qk/XTZw52eFExHgKVxZw4nrf
NKOuu+nwbhek76k+x2YHxwUtDtDKhtO2ak/PzWR7Hpdrsp1N/ZhCK2LlJYjdUdSn24SkQ8QXGHht
O4jLGmZgaDHjiI+2PnqPeoUlvzruwCReQouyNIU6cpvPL85uX7QnGg88u3YF6cexrwHZVgpUed16
sAa6nLvrZ9SzfWxiSaeUrQX+8qFVHp2s4YqpqIOq9MwtUpox5dN+2LWEkelX/rHjAOp97c3Pt4xN
Q6cMiwBrgbWtw875WSsEuIVecIwTCeBjHy/ErFL/ttDMGgPer1PVD7ti8YvhCgi6fIKwHn2zSJnA
gMSaita04d07gTTL+504vEvaTD48fpA7zOEmRJ4tgp3FncQNYayZwK6RbDwBEY9eOUiOYv2ea5cG
E/E3ghBahgdUWb7n1i3W6HjeIt2bpy3ACTrsIiPxci+K46rVhuPpwoHgDRJ1BKPWqGJC8IgoZ1KG
ucNk6ZfhPPxUqEbSWprfDkpPeJWGXvN0ePkaEhKZYliciB9jdLVBxbFDi5RX9gFU8yeJm8GdnRZz
n2OGN5MU5wY9BP7YFglF1gpTero/LY3PaF5nuMEFfKmVD6EEj0IsvFaZxo4k2OR8e796ohK8SENu
4q9Jy0KuQ3aK+xCT8f64LjHVzTtK/8KS9L2d6WCJ7dS+Btz2bDrLjxqHWqP+r5x0kkJZa5pCIJvw
se5nh9bYDXc97DNDn/yVZoxb9e08tIeRoOTvonpY8xvxtHztCKTcWLOormouXz881JF2KtMzf7Bx
04B9r0WoADK5v/ooNblmfpHXqNEWKx1pEfnen+Eb/6m2G/hzzgSgbCo6zYusAhhWEjirINZuwreR
GA1cmvLG9SMujiWUsTomITIqhwRqakh9ewSnCwfAkzaEVy0qt5TeoR8ifdBLFIsNKjdxOyDDz8lV
dgvcwoqOKeRM0+igVkoepDcm/y0TSdQBWJFHqiWnwGmMLhtFtDykJdKIHTpBQ6dxz5a36SIi98Mx
zL7+Xg/TPYYVyfl/3z819X/vFpDl3ejcRh3cZ8ocSW4sxfwiK5+j9t1bYljvHOJBE1Ky1wvuCTXI
zchWFlGIW4mkOlGnbYte5J4eR3vzu/RC3lFj+UlDqvTguVTlUI6HQlc5WIPCdwXaBhyJHUMTATo0
Px7TOYbZ/r+1JcLOwXRAORfsPgI5hxOMzRHK8nouLAt1uxAHyVXZtTCs4T99qJd8uEagh1RqTV4d
p4TNdMgxdi9foFRRZ4rNauW7CV0D9sK1TAwB+EuQklkR4J5451lQf/2JYWvUY1ypRxuPLHvZEljn
8b/7AW9SR0zard8YT5Cs3lWcrtplchPZs0jzJFUwm4MzMisV+fwtZQdN7HdJK5756F5Fq5ozNH48
3PMH51CXqzlYkOt718saTXlTPK4WFApGRm1nAX6KdviMvn9JHppFtkMAIkpgc0tvgk1bGHebZKrG
GZb/HqajwYiARYy+RnJzzhuRMdImvPqrcd14ZHSyCs6p+WAdFRcG4iDMWKNRH4jfqpt8mWzYFncF
HE77WU2NQ/6gW1HRS9ac3TuKR5NRFmxFNebVFQsghxqEMk6RBjs9rG9/J89mWwY7UABCDd45lu5a
qwodXY7MCuilcaQgisC7Vi7cMd01zcv5RKkVivVhMoJ0+3A0is9q5UpbUzUs/eY5WDEFc+9DS1CK
c43y7ZnLJXImD6qkQOVqIXaBJHpiHhNFEW0IKbElPSxyxzxJaKeCLxoW6WXMFPvDwvPtWSPrG2KK
1D8fxorBlZG7aywMuYTlxg4ZeyA2cYEabGpJh8O/OunvguNBNl654itfZVsbhe2Y/s8hQMMWVcSK
sJT96RCdVt2LXSSJqVnLeUorEseIaFZNeSMYGENolaA57WXQDBVthaKMP+SX/lRCs5wTNXOD6lRs
OIWnlZkRQ6v+hdMPYVJCiDYNA1be30A1EkrXRdTRKb4jnC6NM1GqDQJm3UXFqBhilRTEcBwwDmeq
8TA+XQ6FddCwqHq7mxjIN2G2YPmLbMOx/uimYaYoegCsU834kUivD0BrwWRMIerYFikKK/kgcJPs
fkgaukn93VlAhx3z9ylHH6Zq6o+hDc3use1Ggf48Xj3OGCUburbHMVsyU/KneZNnxZw9zUigjgud
jM2pHxyqfbnB9UrS8tlY7+8fZ29MfiqCOcuUBNutoQ1bdqVMWGu7dlu8Efh4VHh7KfrUNxgCcmt1
SMkxKAoswWL/v4Tz9dl5K1c6yNj+17FqhDu6vuOlRNunTpeB5nBs/td0uajOD0E672VWs6Zu0P1B
WW0zWU8KTCXLufbxpZpo+1xJZEuIhjk4TVHqJPXqSakkPD5oqO687q/ZyC0WRdDyQYuiV1h7ipSl
g60HcjuA6CxslS1JOwFSE8fWeFhl2gDW68HXkRrjMN/NcZre8ETixfb9TgyvkCMHqrakCOir183e
/XTRenQMiEzref+mq/1PWvLtMIzLA2RJ3txEfYsogHAzKshBMq95LHpEwtGkCiP6fw+sVe9Kc5/K
N++NxEP9ZQd4fnkqS/T/b0IeDBmXwV2pueOKBValYuYXb6kZAy4TBp32iTCpjGiR9cQDGH+EQfqV
X2tPKb+erFIxPxJXW6H51FRvl7Gzh9dtnUIM2Ep4kk4ZAXGthGkk+OzMeyxPwF8f+W93Zp41/NbS
iVolpo9qFLlqoijjPbK7Bc2K0II9v9wjkvSyviSKIPQbf9cNGtE7bSJ26yniSEuvSIc6+9XJ478N
SfHcD0HrUBAmdDy65FB9iTzy4jTDfwaHBEGN04RLgfFawY+WKwqXi1sCXhVfKRu7Z5EGxIv/aWtq
JSn5BzHlgriGjrxDIoMiAJWyW/l94xVHrRO4e6J8xEMCBlgmRtxporO4TOrCRUI9ETuRL9CL43dq
duoWl0Df8KQwfkaxU5jVXIZhWzwLyHm6V8otjr3Fxw691JksauDgMOpltx6xtdNX6DizfClwOtbL
iHzE9ng3DKY2lGJJsPUdg7PDp5zAQsiuURUkDKGNdUZO7Zvtmzd/3h22Ziy2AKr2/IC6Po/qmvwM
BgIHz4md7OK3HqN+Q4ai25eh56IdKvoWR2mXHK6399iXShWZRpfwkiRz1HhvvyHs7qcu7YHkt/MM
uZQ4aIcqV7BeWUZM7niWmJICuChOkDBGMNc2IbqPlG+FhTRhQT2X2I0pypn9MD2xydfNDv3yYHlC
GPfbo5vOzle5OXyF0prXxQG/wfYWI9spMVdQsn+ED1Lg++de3OySAsiUSjiddB9Iwfo9gcdwRyA9
0b549VV9aKsV3hwOs93SEf0CKOpWuPzLt7DcHHzbK3y9anb2YrxTEq8HI3xQPivh1uCtNQ26R0a2
EnRgez2R5DuXbXypRzb3hUeRb0SII2gI6DE2A2yVTRL32KeV9OwWDzNDm4wV8AecznAmpuBJunpN
bqrappYlCpNSeFC+2cEeAY140Ag9OE2LsQ7dK3x4gOfv6iqPkFgKMqRWLoJ8Rk/O3LOV5hvdrHP6
KepWLfHzi41qonZGCCyk4ZbgRUnGSsrJG1pBrrEfZU51ZmoUVvoCcxs1DdwH46QI1dLXGvGAa8Nl
KYUKHlnFKzj+o8xUlOOqIPkA3uhoX3q7I9V4BZttymJe6Af6qpnx88V36D8QydH1tnSGckt9OgRb
90N6Zhn+00/aKbilquTLy0NwVsRxWPwvi1tRn4Z6slOGF4PTya8lIE14sHuEFsIbK3m9/qzoAR3g
mnY3XbXex8PK2JoOLFYfqrll7CiHWxGrHzxQ6vOcx6bDxnsUP8yPdmt08KECDaIwkz4qNTGeEeK/
fUQ9dgzD96ZLn2uE6OL0hvYhq/xQXKSaUCQEnXuDSEVTuA8q5lZ3uWVy9NvJW9tkG1yEvhat2FBs
sT4hzKFpx4UWEsluhjni4JKBWJxa6STORFHPU+Ycmnc41jklc4vrQjwdwNHTvq0e0ZLobPiX71Lk
KqFyZgtWHREk0VJdXgSzG8HStFOBL7aomAWuEnG+iM/HDkVqza3sLz/7MilNKOVgf8lk17xo9hVc
i7+Xbk5uDjB0TWxRXIhsl9DoPaPOsC9RmajauE0veS135qinPJJg4ogJ7bN1GJfP0B/YTpn3b//R
LZgNTDj5l/nXTOlfc1K5sSAX7rWVM9ykD2Jj7U47+M7rYH2zSsX/55Ri1ZCSguG60UQClv+WWBU7
alW/vyh6aBDWDPXwgoyAhhHdApYRzKgEmZA84FKNgdKisOqMMjiUPRLjZA5HvihFG2mzPbka0juW
iiAAxfHJwqv5Up53wGP6bxiymJlJkr0IiWaAVxJJGdYeYcZN76VlnM+COb4Z/KeFBai4OgiGgDTt
AyCaVddWlRHXuAaYkpoScBtIYUHOL1T0rHrrEwcFdByJH4yG1s3ky3pJOtlYFC48XghQjquOKlC6
n840mOT/ySHrnvpIMNNGwSH5V3/mZkShzntbbJxQW3jVg7AWXXlG+iJmaFZn2j9wfmguJJEenVMn
bTRIt2EdM1xRKTp9naiG2IeVVyiWmGTXCO4OMLsG7eA9kRKpW2lQuLvfcUFCfyhiHtqdDCSx5IgK
Zkft+Q0RLezT8bgR5/AYJpU3pjKOt2/tDGdTV4j0OnjTh5ZQFs6kVhcXEh0SicpEUSr/Y3wGWZI+
wCYT+E3j900iBy/ANbHKHySNp/5Z2RVIZjTsOuSeeoGieH39e1y1DoPx5qWdbPzD+fU1QlbE1HaQ
OiLiBd0ku8M6yurZdd/FXoNkDRotoOcaO3RDiie9adbyE3cgxgTrrk81eEPEAlp+9QvKT/SUOyAJ
AG3+sXnlTvOQRPsgznrVrGfTd2TLqeFjVfHVF/OfCoBmtzQkq/hujh/nySvVXTU3LnbMxUEd1xU3
UKz9JMzhSOavPzqyagstuYVwmfqgFBnmMHp60fE1IoemfsIMjNO2TCmDoFkhOQLh0RHpLIvmPED7
G0XPK6O6mnHrzJnxo25rXGGtb6x+1WHRGziirkbdGiwFo+uKFSVJyEjQBV+LYOzLMCRXFjmgB80x
RkLx8q54YSo02JQYVAcORu1y95ekyNoELCveta3FN9jZ0GCSBx9JnNHfzpvVzfBKvNSjhwQiqPwV
kvBV/qFQtGYWE513hwScdmZplSyEcNVIQO9KpS9GybZgDmmqv98AQ6qGkC7EA/6DNpx/vcNs+tuX
XdR8EOqLBAnrptl7ajJ4Yc1VXuQPrRnN2ppdzLWH/LtqNZ3zOeTVlRNTF1UXVHudzaTspdd6bEY3
gzGlLR/wgDuigsW4LygtBlyk/RyzlHgF9jsTMK3EkRp2SgYluJJjZqhkp/lASt5m0sc/yInCOW+E
OeO6nxjpPuRMwB+Rrsv90ZpPc28q5ezy7iDFDSG4PCj8y6pLdi/PxdwmjRSXjLmpoB446m4NmCbj
UDtlh1WBFHgCklvLFoE6h0HBmiX8u368veMvsFOP5KAiIuRDNkWUf6CvXEPzoov1TNJgy13Fu+JE
2gDkk+UKv5kI888V6Elm5SvzAQAaO25EaPCknreQkAAZjiEEbiQnJA65SDb9PKn9ZFIryp8tRpSX
bGYm0W/ynaXIv8QFEb/gI1OU4My08H3NlGgx4agU2zXDpFk52T9JU3Qo2xBvb69a28FUWL8txjEe
TBbezMzvYEzwXc8QlGL4T/Q3LvXlybS6ZooDnYobT3gKR1bNCM8OsnAWhbvw6iTGWKxTf7J8xkiC
AdkPxXPqTqTKZo4IJ11s+FyEnHjAFAGR76bOlDRpPw4L/ZdgRNJG95+f4LjUamqoJgBnH7eDIUK2
gxJVmhz6RCcYUh4OTQknVal19jvGsv7UnS3oaPUKrfGf2iF+pNGgOlUdiWToKAcFyl/sFsn9c3kX
wsX63MJZqX9TM1SiIwmrDTyc9FFl7gmA626/Ff9hdxG0EWYbZyPqWbaUxQL7ADwNEl65i5igH0RR
tkQ/Rqrg21++DJVbLQXBceCWHxSsUTpgGcsiZJUwvKWbyyEWAH1iDVXhP/LaF+pHnqefMGhPw1zh
D1hIXvut4Yq9ceC15+15zaQ4snJF1G6UE4DTgsrQzMWpBfcf9g49l9qbO7dtd0wzrVcyyYoXq8IY
OJiqognrEGkiIIaH+hpWfNc4JYBgzqjNt/6rAE9xkczsshJpUlb3hjAk+zuLE6lU3wIeYtX0Nfn2
Eq+gHi4SdXbErb4ap7odOMuowvD9yKhALV4ulQ3nH7S4/sqsLskKV/90Ty1RQ3YFz7gDqDey1LTe
jgAsHmoXbrMPqFQ5JpD+NfWlOYBLy66k6X9VBEOCq268pYQimzxowBFG1urYkwanyD+KmLmgWnvS
93fl46HBVrAHGfrlaqWxP/hwrG+HXsypyEmkaUgisP2gOuz/qSdmuNBQ6k9ePyrPTcVGvRjIr7QB
BiSwZSjD6ThtBEoLFwmDYSsTv501Q7BZqI2qhHt0iJI1AQc+8YIMtJIWLJj6lRJhZWoyIFgh6rpU
nPYBk/7QkE0lIJuCVsollqi0Lqd7yfcubPUieOGt44J153dGt7h78jgXXsfQb/hMdGt3GaiWIib3
PRHLioslOYbQGDPQ1I068PGfDErGPlfH4rkbE0lNm4L3DpmYUv49dgLSU4sna2gAiYnwC90dDx0c
1gh1rP1p5nH3/C6e1WlkOKx3jG0vTEtQy/XMVp2IhgeQY9tfNbTdB24u/PDk9wTP0rz05Gp5R2at
fyUpL5sGhheUZGRJcaZsiyupWvLiycZbPEoH93VRiF8mT8D6HGw3PlTgL3ePheh3+zgikuZBVu5Z
Y1Np63Mys62xOwrLQaqvDS829GFVjREUqFCHEs0WPIdTH2BcduKOc8j+Fytfd2syE07nPju51S0t
MeyoU1virI8nq6gOfsMtyPUqgJLQXmidYFp78Oe15RMc6WAxlfOScGOyTuCas7liCiOxemdI3Y7k
wTfrbAPvgsth671zaBE0tZb1lhyXrNINGLJmLUMM/JrD94uY22lFR/7SfJyrH6YDEsn/aR/RZwU8
sWWJAMwYOwkNQ0SD7kuHCBAfmkY2t9Lp0G/pYOpcmnxIEjdieDoa75OgL5dgRIwsz8HhCN3z2Zk3
SFKYnXnfk1RxcZJLjdLDf2bg5o2Q3zoxoWfmtnB3T1BZocPXlzflhTBPZn9sWxQV38TE2aaHLQUc
pxiLGi+EMqcYQdG5+GMIsgCipwKAv4PvdJo53/ChPTMjs+NSv8WXARFU+m5zz37BB0ZVKHi79e0V
DB3mtXU41REqR6rIJT30+ViqjmuVioqN1fmp2zVtZgvVqm2ElSjaEeR2sn+Zcm5KhnIdqHCds2QL
p3o3dANWrWJ1vWGFX7R4o7F3f7Buk/CCDzf2j6emowhYvV5L0S96tOmAGpTzwPB1Q6w1FzWfoxiE
swYegBH119i6V/GKBGsJSvJ7f+a0WWYurIdJNFzGqUJCGwWi8IvdH/8m/rgqJNm9aq4utTpRmgSo
ByYIuOlMXKhG50tZKnylU1Fg7NddTohMkLVxxsHksq+EHPZxgMy7DXMXQT7jOh3QBJloWWx7zK6S
xpwglfZj30CqsDsg/lR7R72u7u5W7dmClmCLhbNHTGj0dMmIUL9NBQWXxcNGn++s+grP43q+a8d7
uPVoL7uSfsG14U/iJW2OI+S9tLeSnua/4Bb3iOgT0j//uSVOr+6QshgRzqpsaWxI8vWMvNFPc8KF
qY9bMNGHX4JZhAmWF5AVIUQrOCD/Bl5yOML5WPlHUkuF5Du6pmIlBptOBdiAHan6NXGDnsMMpFAm
pe7EitsK0uBm+rpjKcvnV+b1NapILYMjeXgRsmqboDp9Ze2llLrvye8htxJ365uY17P8/wdlR6MQ
812uUAIw9kkAR6l7leUEM4mFm9tbg91Vu8Dk0YJhGAKDNzgCGuRpOHtT4ekChz0SBp5maRdv4DUF
sEJ8WRv+Cud/oLx8F4H+ag8AViFozW75CZ3YfrBfqa2/s9Dbhp7pPgYE9cSVybBXU5MZB1lG7FbE
SJOFgn0gXit3gW0E/vNBR4OC4aD9t/mOxUZw5ikcgKHRatQUOqgcMWdknRhmpoRkTzB1OrIOQi2E
+7wDdwIpSSjLeRf1sm/mKfe7ureHY2zRC1eJVbMCrCqlerNLyAOphZ3INSbfdQLb2Kmf90QJQhkK
vhCNv/nAnRytSdx3e9pLVo93HvRgetz3a7KcGNlKprGUIAkt2B8QFA7N5EyVtFcvh8zLk+RLF5NU
0PyzOU5BQYOhvivKVXOKJ44eMVWOHzyVvqVxrUWe1QCa2cJWcFlSQ8yPAniZtg1mSAK2eqfuL9Z+
NXDz9cPCTXa7OtqogfmG7LklynUy4/hB42rsbh7FufRCqgX2CwBEwy56B5VZAzIxJdmbY7YLgO3w
7fj+N4loL0rRCZhL66pJQiS47ELVzbDwL/RJEgZpn/N/ao2bcLogf0z2+KlJY/wiz0/e/qzxLWqi
OxUc2QQmwhSuV8ZjkAzDUTn3FInshI2GYQesioF6Fj5BioNSSPE6Fv3m+NRnQcC6ZkuSWIujYuL4
3H/j17gshaXZkNObcOlmuARHIOj5PGTr7rp8pD+6RbhCsmvMW+EE/p4UiGXbjC6i71Oi+gpU+SKh
kgakg9ImuoHfi2UBrFj8jng3alJvJet1Kewk/Y9b/oYwbHp6dEmWkyAmvYcMLiSSaDUcTs2OpNnL
Tdw2JVJVBFjpDrU11fQtljZDxr364LVJPO1H7hsjR04AlS5BolLiJ2PFdn4eofwmW15uJ1Kv5h0y
QggnuEMEBclWoqkVS8BKnh3ynCPML4du38iRr5nu7e+pxR03R4BAJdh0qRbgLL2AAk49z7ajBwHy
ghrh9brTdJhQYsnRY/GWASCs9sAwYYP/WfTX/NrEGygGfP6dYJEjWobdoaVsyfYFVmrSQdyJcA+A
4tVBAzyVJaSTdYSSDVMcKKtp4Ln6IumM6qMz6gmUneJJVvJRoMvgf8fyuPiNQMnWFcwwglHDauAc
70m0KC38klsHiXNgmJ0BRz0fgUEQLRiQg84iisph/aOvZcJ/UfyH72T5imSCwkv943apflwnJFHA
LKQyzsyeA8pZLwVOnzB+Je96wfzbyLfLtjFdRN2A7K+y67lL7+YZWuP5L8fmVmHRNdIeMJ1z86vZ
GejCz6wI0qM6dMV72dP7km3gPmDpBAsM3txO3yP2t0zDiO9tRFHwpDCoixTJo8iqzbgNfOWuJNDi
YVYNs/Tqan7lxwSdtr/dJ4m7FpMNJ0ROIj8EcnWeFyl6EzW37NfNikcjqgxgv2E65yqSFfmdqQzH
Jb+YjU5eUU2Hx8+dvmTBxenZoWnE8ty0AsOhyX1YlKx7VP2AudVUAODsF/tNR+bRGPOsqQmI6Qot
4ylH7hw+ZqjpEaQGHkLKMxQY4XbFCv6YKLNghu8rBn2NJ6AgOk6Ih152nHU7hFb6NMfkKIr+xj2q
rw4wCTD4pDltVtIKgohRiBvMph+LknIGM6wBeK+lBX1Azz9fm+D7gN4rkEZHraqR5eWJ9sWHV3hF
UctbMPcKzM61zEWn0BLeKSRbBBonqVY9jJX/0DHvlPQqhSFEahHA1DC82L0MGG7SS7b0eC9aTkXw
oZRu14QMeRN6Y/kxY8tmKmN59Kslv/8jEGT3gyoAPOWrakK1dpyr3SI3V5Ze0KLBRMvcU5avuH7j
VX1R+Ip71krLkplY3kM3zwOVJZBjGexOvd5bG6zr7Imxr27LCRvOjjSb6xwFkZw4KcIZpluqv7zF
D0cOOpqrRLbTyGjHP+l7xVBBb6McSxy2GouLmV6o+fXy75Xsr8BcRcK4ueFk8q7ewTZJ7oKX/239
UuhDwjWIPxf4I8cdLLsgRfPpMDAID1vB2GeIa2Xu8zOPF8LF4ER3yuybhKUKjwa9ljsKQIF3QGtY
0XbhKVrgr8UIT387B4MGao9ogj7olx5SrljZOG53Y1MxD04ZirL7gu8PYK4rvkFhgNshgSYtOppr
CZcSTJvtT1FS64zb46Wej2c9OldMILf5G6CQG93vaEEVxVr3rUpQWPQaL+us3ZMWFMHMxcJvcFtT
96x4VOd13dFUJzWcxIqPMMm/vTgwmILs6rvomBn1/IjvB6GECKwrhT0JVB+WqOmWXtLu0mOCzE9V
EstyYy0erefZ2PhhHKZ1Q8N0WRNNWhZKxsqpr5+mKy3v3SEqd+NdoovEN8n2pzk8++T7ibNjHGAv
F+vccCGEWkhbVBpehgWRKk/bbJXd4f9EvFBBdIEXkCWSzfY+3ahaFoT4TMcNhbyJWBYzttYoI+8m
Y6ZV1giAhpBS3/gAxYfyMWBHowaro5XwnuP9jc6QMeIc3u+fwiRPfE8dbZHK+yvZB8qoBYUAesR+
+o749uvaheNOHvt2ats7uAh9ldRMJPWmI6KB9Kd063cSIHylNQSool7nySJbDBjMXsOwDK1wqeAY
mAJNTJ+oIO8Er27iQxXwFoWigT6/0C8BK+YwN2rD4F5ljPDKWmeV4IRJHyWncKmkxvWmFH50Jcei
aNijn2e6Lg2EuqV+kAfWPelaZu5nIsRDhFgpuK61ZObvPvzwE/cadcDqr4jqv3W6TaVc75T41XcV
1Hkb1lxCyTbKixP0Ecga8gair9j30LIi7HnexR00dv+I94RZ8e7p4dH51Qog+W758bome2wMvXVl
1d0PC2E8CGS0mqIkD4PDwTIYUqGjgUDPzNqxIsxqoM4f2Zdq/oOM5OlcLq7zpsQI//HQL1uFHTz7
P2WtDqzOTmfd6FUDrUvwUPwmNb1F62+PemV3sGnwtz9NkcvFcVdA6yh5NDLKsGgwTE+SaNVaEJU5
mcnuA6r+/iWsMrjy1iS03TrdNgPSVDg5KBAWiPx/ZdNKfobWBCvcKiT3DWRV2IMi1h8+ivxyGz0Z
YNM1thZJ/Tg88wcW54/0nZ7JwLtaYJRAJmzZ9F14HLlBtVGGLE67GnigCSv3katKEweg3VtVh7gM
B1tmm/ir4bAqvJO4/2Z+IQQQEyA1wViDeQUAwX6yvEEgBdKIY5+hMYmY4tn9Mz7OzK+LNQEdDlpm
3sm2J3ZH/Pzg1rEeEcJRFDcsmy0r3L7/E3w6svP889wwEVjM2h0Gs/Uxod6FkJmB/XasHHA1iO10
ZOQt1kY4UYDxw71M+bJiwMfLk0vDT02RdZGZl/MYtJfqQPJZ3hNhtRZhEm1oKD9KwewbzAa1ZkXA
pVJIyfLOszv5Tmys30X5zBqaRXBue08ll8WJskl6217MpRZV4n+EfbxNpjVlSLZC9WauUE1buF7W
x4E5LkiX+WQwIrXSzHhxL3v3J1/fDiz2ZUvTfY+HMYBmipQ+R47hlyFLoxytFKnDIu8GpMZ1qULN
pSGD/Ydu8E1Wuoo6KQCG6pRotgRuh//pu0vl3j2aHeMUNvIh3awlLv06MTuCrHgHD+M5GcCWcaml
pFLhdNShroC10MwOp5PyVHZAQvQlN66chS59wsJpIwOWerE265/Oey0ZTLGC1Rns5tnZdvm/aEh+
hw80eX4M2O6C4DpmHBnU86e4wks1pdVccPbHD6Y8KHTbONOlK2vDcR+AfZJunntHeWyXf4RGIOiA
mdQ3YfrvrJxES1+ZdMxDyX2r8MzL6lUQ0x6kguz3Q4GIwAwTvdqPEWcPKsDDI2b5BV3ZctoOG17v
70pFTu5McTUIF7f2DiP8OwIn96P19rGSrjCSCDfOeXTC/16Tkx0DyMmW7QcZ2PM9ZlQ/CVTFl/1m
d/c8pQtyimxPnd1EJW5d2wmB0uIt0VBeCtFiXGGFoWVxj3XQMgjaRX9FfK3kK8fURjiyYNJ0aaKW
4ta9qIIGr4tfpxO6NKrx5E2IWXR81G4XPZZw9nLC4gQ40wUNt61Ww3DCitGy2lLT8emXkjBmx/aP
pnwU9n6SVs0BxCI6tbsxw98EXR5EAS+oCc6pAU2g+8lyRYvOQxdNG/udyGMXMrT5OzjIPxDFIrM6
jWZbPQWy5Q3Z1Jx2E5tCD4Rm8uja7KFB8VNmZ1Xyf7Fd9+88+ncaYFnBMxh0UYJw7N8i4jjwUEvT
+SIbezZ6ktbQo/vC0wH10PL6f0Pgdpee5wxg/l6SkRkL0SSM8aHvPUBabvPNU0VJvLOQweqW8N/N
9Co/nV3czan4lQ/gvPXPfvIu2aPfVZBaQz1JfpJbXYuVC+KEgqqyvZVjTbNlKse/fObUz9qHWgsR
JKBdsnn0NtXMOdZgblO4AsG0kJ9D44Y8MdEzr/WvlJuvXWlbmGuwOSny8X606unw/QSTlBHV6kOA
hvXdmUdD5YLYY62Uv1w3d7+6D+cQ4Rn0m7n+qmXjylBE+nX06/i3YsHJyIVs/U9aZc1Jld470EIJ
Xi4OQfHWWLW+UuG9FeP2pK7aWD7SwLDpB9t41MgoeAopnAB5R3lfpAkJC/OQjrNfKAd1aGXkAVH/
cyySn5ekpc8eUfwnEQmt/hwfpQo9ypCwK6qv6INcVxuQscMGCuQAqQfktVs+uLOnrQRjq2pEqe56
b0hAbM9GGzFiyypvm4H4/KlG0WR8tklpdxRIVeBSv95uMqgv7wLhbO3AkM/iMXgsj2OF61t7GiEi
a4CBM5d11jqKBOxw/FEuXZDO868/3sN5v9RBb6VNBLu7bG0+CT8J/Trie6InD4JKQk1WCV4x85dU
XV8lXEkqNZ2/045E2hk71WGJeGitDKy9ptkuEe+qc0qkfVFLeTPCuTWqkC3BW1IX5kAQ5q97uk1y
QPtDDbGJx4CeObT9FvcyA/gCqjnmhM+0Fycty6ygIBbXYSucmr0mQ+pFD1ECJHc8Pvfnjg24XyMR
1/0U6mgz/+0knWcwvWdP1f8Kln/6HGntyfAS5luohAXvExrD36BpzUu5kb8bYF3qpQzBSGcMkdqr
/zVnT03yYZwQdoUTaU4t9SAwEjqMCFJBnhRJH3J179Z3zBgLTV4tPUSiZkiXxbhWo1WU6uIWqiqd
MDaN8t1EaYooJYb7F+uK6YV2FH5AxjfWlY4L91HjvqnIKWX/nGYgXLKd5j8xInCbjBjdRwu6AZZk
kG21/umYvqYzmQGSSghGAVMaWas6ZvvPAujNB2Pxvt0FkZ6idxz+QHB9AyX9JKGqW/vOCfFDihPs
89XQ9v7hleGF7KsUvpZwR8amTTcPrqXyIWz9y8B6s/VDLbs4wopWgqW7Csc6nUqBp0/yFDFRN3Kb
M8baa8cfKbecVHa9iqRJPJ3mw301NatrLfwg5idc9bVrF5yUNJBeA8+ZumKYMEMeWMJgyN6Lc4Vp
G9PUg+vO1TOo/mH0uy5CpKGs6MiXBbDFuaftcVKoaIvuSLUJgX4Lo5hFHQLkVKKidIC36S8SovOK
x74WXsAc1vTi9aWQfUSjB3YT/q2ATIPmkJ73n3NBK6MfkogLnZJhusp2QUsGrq/PTMFt1AVcEsO8
9Z/B40J5xkAZ23+Nk4Iojd3JahZcMEHr3br5obHqr6uTNN/FmPlt51YUWW/5EedSwoEPeo71xkSN
cYbYUM9z+5AeVRSFvVridMVFLzcDA/5LmsQ2Upy4EoiH32bW3J34kiX7Kcy2VWMvXoV3h4dcDKcT
aj/0UJVyb9CU0C4HS/gV4521cFL7fml6Xs/LnmYjjW6RlItIRnKos8YFbuyNVI1tEMj7CbF0Y2tl
tID5xqPcDliF34AjY4AN/DsK8Zp/zlrruqdBuFZY6hIeiWlzz+SpdnU+xnDtFJD+DFbF9NCyGAyW
VgcKmMIT1Wzq8D+OjRHAnWdLl8Miu2D+F9Tu7O53I8EkKf/d+1nYSSNHFabQgPXMBMfTmuRMTw9a
b5yJbctMeYULu0KDI99NLKT3vryODVw7KC/OzqEi/ZmEFOo4g8UqNrzSJ2T1oye2psso7QzaAFyJ
K6MQSs+mFXeN63y8/59u0es/UawgRiMDzQwsCWqdhWWMx96z1+Ondvy6aXO7o4dSOlNsHwVtwKx5
cMKNuWfe16oeSn/DwP6OACPNW3PgVXDMJoIctwVEGLfo0BCmx+CFdtx0uyU9EsomzhtbgDc+5IvT
R+4D4RewAScmk5NAHA5Bdnu5KYk6ZINNYKlkVBz8QmIPTDINq6W62D7ohybtneVBllGZs4LQ+/GJ
6w7DdPiSY+xhHB7AQqpVD+7PW9fmFPV+raoGJF6mfSrAqmVgI0Yrr2Bw5VfDShaMq4A8g0JGl4NC
C8BWfBXOuQCitR622hZXx+eyMk+N8oVqUUmEvcxoCBiXw9D2un2aClT94fTWy1j/DhLY2zYfMp47
lbksaScOVZGaSr4QEwfwbtuGG8SR1rmHh5+r0wlc0AulN8AcQe0JyL6kljou6wAhb4jUNlr7SEpX
1mYkmh6HopLWrSTDrqB93n9SIqlVPO5cGt4tRy2FPEPs9MXPgmSOwrgGyT3VTdK6/IUAlNq0/HGA
6s+vJDTdNt+7CIja4s5of0k8qGWgh+qMTa12FR3Y+BXPMCtN1RXJKZhrN6z1qTC/SRA7cbdySV1e
2JZzjX/sXKNK4SVWihOBrq5xkCnFDzazCR8kmzECKIt/Cy5qxCVGshygaTOj4M7TwqxfjeThXEQ+
fzZ+H0iXaMKNpHNJurB3ZbKDIzyhD0BP49TwWVcjznMSFLiudUmWdGnfW5EDHDu8dN3/+neO7zpU
RFVhTuXd3RBSSop1gf1Ziwd67t7RtiYg3GFfAHXoa2KsDg8xH9ZTuBfgRTbHYRyPdjVO/Zp+PwBt
W1bBLDoogZgN8JmAO36DDH2pH6a3xWdvGJvLJyJfsXRmos4Vuk8c5M+/G39n/lMuDEZ+FYNME4Zb
g7brXnCcld47EV2VdNe4h/sk8m7AVbcHvzYPOckPLQpf7/Bof3WCx06rFmhtl7NFadjefWwunR2N
j6KM81Y5zVvr0ObR5WOCNBxpRcpSJCvSVDy2eyTCetDA17g6Rh8ABBiJe5tEo6VquCrKXM4evAKz
zT4JdhbHUe5hBczInMmKNc/a7zTzt+xybdokz1hCxl7SjjqiNZTWvJRP8DUuMqp1kR78HybuRUrR
y0aPsoFlQI9xv7652Oh8qlurVBXtSEv9U16O6Zilkh4gvV84DeSM1ggjGh/ibEvwDbivB1sjcFIx
br9iykQzNCjFFxlL2vICXDFL1y1IugmzZWp2ZA8Hrg7kXc/VutAfSc+5n7cmHIY/usfGsFkK3eVr
Yk473rwI8wn/OZhj8uXwXajlh7Nx5wymfT6dGpOWsh7aK9RYGWeHqscy1FMx6SFL2OrWNPJqPrCe
PO1YurvOYm7K7N6W+aepl/rbo8EGm3ge50GTGYs1w9oy7ZKJFPplMALkb4nJPyzkhfpYa8EdvRVX
BfzarukGwXdLVIAWkvIxeZHHAU8JqttsXwOtqUNSRb0ZCc3FJ7v50GyjnZ2Ie2T6hx1JAn8OR2Ls
b6DUihdQDLXzyhwm9sGqZUiCnxcYYoyW5wreM7olTr8ZfInyToRjv2QF7OSA7rNv6yLIZYl5xPOp
IiI5Fos7KLJ5d0Vq66vrObgEhpJyTiZOZ3Lxyu8FesCMCwPi3Ieh6MmisnoUCBJjH8GU79IE8iFd
xOnDk/zCtJhCVZuFx4KE3Sw52i7gzpEXSRe06MS+G+qW89U9sQdBqSX98hIh3mw5rlnY2hnvcziC
L/Hwlt5X2nwTBD4zHOnG0e1u1RLy8aIuCo56FEJzNbKVg/5aYghrDrQRng6hrb4+Xq08oZMonq+8
PtXt4HZj4hTAxZyl7vYDT4wp+BRMGUhaRgYRwuI1LcZ2DPDU0+ckHmyN/ypFMpAb+VSZ8Wctmh9W
nF7/59iQC0sINgSaqixqXDYHBHBbs/3DcYjuUx43a/CcWRILkFDumzZvE/yK012iXKHkCO+H8w3V
7A9vAwuo2tgwrajKdfzDyA5YKIyYlhJDscfbMMSArBqChDWct2Sk6veIy0dWQvqq41gJz9982HnU
GY0/voTb4hjJlIkZyUzWqq1cHmBYwc/U8+1/VaEbOp0a2nCzo3sAUtVwFyVsxOFsE8hJm3OC6xJm
Yhqjp8IbbrlhQVjyjRuci9BGp1sOJM9fF+wVNmtHByoORJDYh9RjgUAzDt9y4YRLFEl3j0NCbhpa
5x0rW87MoVHLMUaOYmJ241PK9F9yf9/XwRi4XQfKX0bohinvXk1d+m3ohWG1Y7kEJZ57ngehmpLA
MgvcfCCfO0mFyzNDUrel1lKR+PrrObHVpaqXRdiNWTK2wvSLNd2Db56mRDavWPVjxwkOTqy0WbSf
2zeiIUvqhEGcZr/4cAyAPol7SEJN22WjH3qggIz373fu2RByjLhrRcN5OXfSIeWZJqGhSLmybNDJ
zNryHblMSmJZ1i8pFjdMffO844XryYPotONeuqWA9wvaiom/0S4o4EN+56CkXdiXU/dNfLJJd7GO
FfiK96jnkOOS5IzgP8hzzDAPLHfeN2tlQ/ZSwX7VCdPKEi2bqzYXbZpeVe363g/rcI8zdd9YoCpW
UFsx/ukAiAK0/8qY1SNWqaH+FjHqZWmoCRerF3hdUmNk4WpJKYqrDhiRsWB0mn5mkOjw8iw8ySxT
+fKWU6SQSd/mOMC2ozb1Q/+Jg8wi3twN4flbNG16aSNLl8TcqPLoZj3OkDwtdhCg38/OV5n4dPJM
6vAmlxTVmCnUCJPYtr2x0eYGBojg+hkaOmFdRMZmgzhu07sA141WPjmObDSunSp9xLiENZ4xq0UZ
gEciWod1LvS2LZVSdw9Vc7lx5cT12a3yPn99QDicyNqQZZXWYNcmEneDBRFH8Gx1yf2H+z4V+X9E
oNu8FKSKRSPAXZjjp9zB0XEliY7V7dZZfXVQFfJff+He33RPMW51xU6dmdtQMlJoKlqvIEhUcPm7
wy6UcYn1GWaFcWj2zeu1IdCHYeNHTsbQDx18pOTUZ+gZRyQdiaK6BqgK2jFKAvvbZKfnh8Olosk5
rN85bo4CEK2noAFMGIgIYMu5XcuvcdQt5xJYIOMnqitBoUEoR7NjA0PItf9k1Z2F4WQFmvrGhXef
XnM3tzXHmlBQ8yc78JB6bVdDzSSzqOCKuTu4Z8mVumspBqMZwHtnBXQbinZkuza11oW5VovqOFhG
hN4znygLYt1bl71IMmzFnUyViGkM+L0UOy8ZKLhOa3kTlNHV4dP/5mvRfbMidFbk4mvjHfEgAycV
QJiH8OaCc6FfWv4ZyX1LMunttbLFGz93by/tsBSSBqUE4iSefxwC8kucxLjUj4wk/OEo12OAMLG8
P2ggrZ1XZbKgGJayxi4v5fewX0XV5/DVYKTiWjIfSrMfcoAdOl+NbwBqHjbh4wLFeKcaNdbiafoQ
iQCA0fsIfcroySvsGQg1z1vfB8VA9rFgmFxlWvLsDOqWlb6Ut3y8U14ajvmeF6GXSmiuy+JfcEVE
3P4mWGi5WtcCFaoNXqcrYtXhVqhRqPzaTS1iY6NKNvK7oolbQX17fuTvs4G9/vjunJDHd/g9wMfN
7JRk+gT0m1H3hds7uiH2Ek7dooyrM4Wj8jTBV15siEMbvrMupI/AsdxlqHeH3gEkTDAFU/ObQl5p
ElhD/UgJCOzAIgj0t6mymR9Tr/f9RBkeeABO4Tr/oYm05b7TC5+ZRWnfNaXNFhJcMM9MHCDiq1XH
MJSm1amVfT4dc0hF/IeEt5VAGyMNVpJd9xxkzk0QlboTJCVRnLjVeY8ofD4SI4bav0s0MD/goBGc
dbY5AEfXhIsBmmJBQIAdLvmFFFmnEBcc8F4yoIOXsSVuAjj2ZwJFmZeQkTaUMuOhpOlfI+IF+86X
T7vsyRnaMl7DiPn4BkL7wcPhuYH/pHzFoT+nVvjs+9fWbMGL70Ij2UVucdl1b3BfB+4AQ0dUbHCo
E6AwHizGV+dOB22tpKYcSTEKSlvWhPyL0SaWLtdrKig9du+tFMXYCRdEVq6sy5p4Enayi8AdjO2a
q3Y0W66onb0FRJarx3w/AMc1Ev7CcBNpsc+vg/5cTA+PM2PJ+5a0LTpcJBVIbiy/fJN3VnEQr572
BhecI+5j2M6RW4xZbyLQ3BKKamB91ORpx7SmOiXfqDZLC1A1wCif985BIJjIuW32ZpeiVDc4sMS/
CpsqTGdX68JSJVJb+Is2MTY3d2GYpcZ1v9dt8+Hsyl7BQuVKdzBA43wyMVnGuVm4CfjwSeUbpi1o
vbNRR5i+0KW4DWYKlS+eg2NE70+oNIKNYFcbawWs8vrn80OkZLl8MJEF5KUfwJWTmjz7vrCooLJi
l7XnEg+LGqaTNoE2ERLjmJyTeokI1EGGE1bO3YCyugBsKlBC3fzraq/MYkfxOdeOBbXxgweLNhdp
lH6mayTTW9zp48e8tXMaayV2twOquGSBG+opsroKUEH3WsEBNM5GUMwxazRsegnd78oEBAJ5FpGj
S6gkCz6L/qbcSkC9GshIFN4dpyYYXNQGUuPn92WPlOU043LOD6C6d9IkgJZOezFcnNP4uJiJA2Jm
3zZilX3Ws3ndCdncu6rZ109HSK1YByZMioApNQj1O1/TB1tg8LUa++IYXRWk94WV5fQDR6XW927I
1nXq8U71PPHD/RvMIVa1Djsmmjr80X6lnoU5t8uXBbd3DoGa/Mv8SA9cQNsuj5Jb7rP0xend03EH
9vJ8HL6HUXmuNuF5333PocAoNOr/p/wgkukmY2j5tsDwlOg5+0vrFO776j61Sqicc6nZOvNQQSUv
l187u/n9NUwON3pEBqC3V04RH9lkN9YPt4WDbNqeaiAvwh6OXuLYfqKb2InFYuBAXr9JDS7c5sZo
7MMtTP/VJPtsnKOrT9dg4mXwa82jxk7LFogjybBGlElbUkH/obZHfHXNnSG+stw5f/ZefWICFZ0m
fiZcnigiEZKsGFcs5Rgini/G4ah4Zq2tXNY/8SxEGcL7Q0mstEoxrwcX2oSwLa7iEs9IvuptwZZB
ck7Ii7gMkz9R0+f8jS2mrdENa6mar7r6Hw/ju4P++ohsSehp3VL7G8gGSGHtPNEmk0fJIqv6j09Q
XeumsgPV10flLF5aoe0oCzBJOIgLdVPfvmEOz9NQ31zL6b5FQUogROzT69ICJ8VbV7v0RV1WrZyi
u+o507Et9XzEOJPPwSLg7eBHqal+gA/7IalNjgrhoW/WZ3dHHyeL1vAratryLSwgEZCqiGAMP9Xd
j2KGagDFmdoIHj4K3D9TKqbGHNV0Rn1pajQ5smd8z+5HYIDKg7+9G8JOOi5Pbx03rF6TT+FseNqb
gHRsY95ljHCcsYqgcd/nm+G9p46X485ZXrh9AKAbOHFUblrnz5Rdw3ptfC3XXnFuYMA9MYsStzrL
bKw6PcBNAODnB/8DrcPq8AVSPLptxmtePHyFFznXQ3lrw58p5aFhaiYSB8YwNZa7sCY1vnqyTrzt
0XOmPz/R8cT0MU5BcSsyJ4uxYNmrrwN0mXDe+ZsGrFA+6KqD40ao21Qgd1z0cwTPCdIVF9R04M/I
hg5aZVeA2b+8rWVAbT0FYRtBNfVmrw/Jcbn2AwpnGhrLAn5+0RE6pXEOMUc8CNnaMHaHriM3tVzs
2d9pG7tpEuH8/CKjmx5oUyw99cH1S6Zsp9Dcou49VZNdeYxSriD1AF020/YkQGUKxIuXHR6n4As7
M0RVXqWrpI/j2DJY+vEI+iO5+xGvLa6Iymfd5E19aOOrl8d1sZ2NvZmEchYtk0/tiDegUj0meV8W
JwHfAy4j6zt45uhFgVCFVkQvJywsS7XfH4VVCS9grJ3sB/m5kfm2ayC1AP5Gpq1FDkI2MtJgJaxh
h0gFVnxo72bR9/QRJMzw15tJgvo/60gWI238itxYsJ/Xonn6CAUzqBP7FuhG5fES3z/gY6C7q5cs
Ht12G2z58IqsE+BYKq/d6xzRw8aUzI4LvvXiVJ2O9nNHYjtdQtdFHo9K/buTgV/Wk3kyKAiZJ8CF
P9bKL3eeQxdoq96CnqlVmdAulzgWFnkCGfXKshIJlmcosTubxxlT4qJ7bFGzLGjK/1V7QGoZTCdW
w0sW64Y2UW2PAJrrSJUQJzAtdnyQa5m9s2hi0BpsCsXPikOFVifV2aNp9e4bbm+wgDcWvKHbusvM
g7C2l6jVjQVHoNOWruPMBixIeFPylu/eyOChQGw7GNXlw8iewlkDCOqVmBmKY6kwMD/UqLQNDaQX
V2TF++FHSvFI4Z0bMoG5aOaHIPTeIMXf+QXwko9Ie3hA5ObjPtHa08HaKdNYLHCNg1pP2V1otb/C
kB2LM7x9E8DyhhILBIygNRYgyxkZJyu/rwFru7LrBZ7OLrRGxXtjuOo0Sr+oHzFxEZBD6+m2f62d
G2hClZ1JLl4419j2h9WwwRJ0LLu43PnCcmXRBBKF8mBNEjlOcDujMmjJyaEWMz5fe/m6U8gDpmqG
JzZ6V8lF9m6byjAXK1sOMa4O5gkrhDG8X5gJysVP168vWz+UWocuCH2F7lJJo67sFC8sUFNIAVwv
OyxCklhvjjwdQ1Cvt8Q90bOYepfanzxznZfi7C2R1kpLCwNDVjacQMFnsbx2wBDzuRlPkWJW49Gq
XnphSyKBzszXgc/aF59RghErX0J3eJSQP0e4rth8Baolt9YefWiHtNkDJ3mU7JTfm6yzfykYzf5r
2lDH1qGmgGRciENN3XyjOXarUxBS7WQ8t2Gq5W/JeGLghaD+kTPSIbKAwJe3FAkywvcQE8OP/neT
EipZdMhzrcxBr67+m+m0VgH4lMKMKe+9Tk8yz5uXrDQgtJOOl4UV0k4PNfVxGGB0Mroa9QVTNwZD
COo9fvK7VCaCX/1abfKaqZ8bK3/NhM9arXxglR4YrEjWhu6SAAV9J7My3CGhDuiTyqZJd7WQES8y
7KQu8J4xkyBslIhr2Svtq8+d577epp8cz8mOlfR1Ur+A1l+hMUeB8/2wYxIMq58LxSnFN8/eGv/V
OlyoKgswH7Scaz3lHkKxXYKWD/uUr2WzY48AQlPdPlFbZnzWoI1Va3/ih1BqRoGz6LxruV16NUS7
YTiJMAK0u0kedgd9S+MEtqOeZEiJSrZs8DipYcPSWETYpMjF4oGapTBzJQ2LM6PJxxOabqikPBcG
oaLL1/VkeQma/ldBJlG8jAl0gRYng5ycDoVkSt7JnZJCuR7jvVeYMWZ9xpwTXz/f/7Kh6mLS3Jg/
3hV6bXYmnRw88DekUDS5WdP4iwks9sD7sUYqxKbtjb8HppxH6EkeKsjL8/5zAkujH9TiCUIWdhH9
O3yC6IrPTXDAJMfwhCeCXm4gvY0XE/1Dsmnmn0Q/RLHA2blT5idSqgOjO7uqQOAdnNLDnGpo9oIt
9dJEcHunj4f7LtnfP7D4fqyPhtkTsKeuApirQFrXPra/DLrYiTdcFtrcWnAlKYEQL7gQ+bk5hnk2
CtXkFEc3umg0SN4EnLYTvNxZ+F9VXiX1SqAp5YcWYYg1nM865AcsQMuay+excXlFH96HyL5/HNwa
68CyU5uCrzNO8UiPZ103QLc/ICMjaNM5D7jsv9xAKkk8gcDpVNqsM5KJiWeCcdzcZQ/vtvUlA7Zr
bCB30nd6JJXSKu25DKx+kd5zC1/ns5PPA1cYhrF74jouhHP9CGdqRb2mRhoaTl72BlRTuz7dBtAk
08DE8eBCEJwzZ+Tkafs3hO2ySGeFg7SD8kVChrA7hMijt7xAlEoQ6lhyaHWdVzWaJHw/buAvXBwC
+HLuUE/8vWei9FPSNYYIAzFYF0ccfTCJsl4pIHe6crxxcX1nYm2uVEC2HcbGQ+ZH5nHywjnJhgmU
xuPlRcs95Po1TPUJn4BRN0o1z+Zb0tRzhggDPB9kgongUVQnhMeg3tGuPtCqxACwmG+aYpIykfyG
oryDjF3LZiB/hVrFCGC8Dxmz+1zXYGRnMKFneCwZhPDk7Bt/Jjuj0dQuOCSXhD1EwCGkFKdphl+S
M/B4aVnZ2MEk9hpulYzJGQ8Y8TPMeJTJp9IbpRvulg8IQg1KccC1V/6brZnzr0XrA4u8CgpMej2v
cMO8BnBUGzo0XLjFzgcwbnk5kbifK/L1RCH+cJFZWCiU5pbokUXqICypCbXtRtatZb4U/g+Dm2mJ
Q3dBEtR969PCYllpodVJBdrUbsILWrE1+pOJEIyMBTTI2RXZdGoBAhRleGuCIrKLvqYlIuxRmrfO
Z8/HwuHXoUL86lOp54JMreiN78GSi3vN0mNQ2Piih3n35XUiaAbNYw3JLFrTuTcT03KyeXvIV1CX
dM2iYYZDTmsF+ct13Cg9BqladnlNVHmdP7MPDPE/251OY4awEHA/zddlzbnUW7IXH5Yu9tKJR3Gi
GdX2FJ/Kr+Y8+wMFTs3+f6Ay5zRy7yRttNiRZYEx0zQl8f5FLqSKNggNOi8E5hD9y7R8TcBSCEHN
H6UKrGTuWTyK7JvQBBnrOU1zSHGHmjg/rhsEF2JlqRUaUh6m96yHSlainLLY6ZVq4ygC2svLQeM5
BFRKzvvTXYX7xkhyfcxI1bvb2JyljUGh0MAvwSMF2CPe5uMmr8hKm1Q+9u1SwfUZ63y1yc2tHVWF
lDPob7lVCN/5uiVa4Xt2Ontn/l623uHR2LH7n95cV2r5+p+yGWlx8Fc98Y8TSAY0IHbZ1WXk+GWR
1kLTWaS8cR0ftNO8oJ5XabbD3w3VqKY+PkeB1W6XUy+0w4fHT0TmfqxQlDME3Tuz2YNy+b5YfmDB
/S2V2cLqA+VIF/Eqn+u4kL8zyMQ2iwyatw9VmwUYsRsYGUDDD6ldyIxO/oMLZ2mlz8AoP3vEvBLk
LjxMocbq+nLhm3bhjwFsIPkbZFpwMQCz4LG5XSa4a8HdP/OJlguXRa9RzROsrqJXhdKp6M3rBUOg
C33UDZGFcqIPlvg1lYGN9SJzrqi/snNDJNnBhMzhiybkiUJ9q7nC4nS7FR9tHrVBblA4n7NGCvM5
tbPz9xs8eOr3+cdEeBTKgfzf9mk0qKq1eAQ3ewhZD3+KajU/wfyM1Z9wesiwKhMy+220eIlOH8pe
S71AbOuJCSOZLAdXqIHPQtGrE16LanPTNnvNph8yOMN2gt1timxbARU8Yj7Kc0CkJUvWMT0adtlV
uBlswGpSJxsojLYhAHO5Hx+PbV+lQzPgR7y/aYuHm80I16UIvyDLM61X3GF2ZHxEC8m+5Dd7jt3v
gtBsMxR5ROuo9MDoHloDkc0R7+ZOQbgPb3Y9aMFjG8/j5funLPyKZzlNDOr9SH0dIRH15GQa68h/
bg0j0mfC2+XJ2Pni4kofkJOobJWCTBWz5cOI9NuogsMvPN9DcN990TGvz3UD1UKAfWoPYrcAylhg
a8U/7K8I2OEyDF22YS1N1BZOW/SOK9lHxOnzlXAzyZ3HvFReQNGbtJ8BCBCcOTbnI+paTlS7WGFg
R32Z0pocJuGxQRi6pizIXjO9y9jQCNie7A6VfHyOPzJDFPfXxM6kyrOjnKXv/O3s7T1GKZ1OnUgQ
YslaOy+5dIv11MxC+RqHQogJp8BRS1lMx6Ce2YDQ53Tx1pRGOgZeez4yEyu5ei5AsLUOD0xje8Fl
Gx5Y0hSq6qAJ4y6Nhf9+HC5AS4ARuzUdKdgArfa1+5NRWl9spSz98R5DNH1mkZKZaGLgP18F8w4f
6FoPFGgarj/WsB4UY+kwG8b2s7b148OMYb62YBQMH+4Ml/7W+m1S40HbQcdZofzse0nriKZMhQkC
tx38SgiryWECjezUdnxFbwkRAqOZNbirgpwZpi5Em0t3D2k+HEnYVaX+PcWCS/8/jfXv7U2XYUqn
TB8qosD3N1UcdyutnnFOGZ7O23Q2J002bqLr6VC0xs0cOHBm6Sr5GngVNnQGD51DREcnI3/pUanh
PDlwXQNwLPNA/aO9tCKOxFpqKDqUKRnlu2V70mtl+SaqOxRCErijnGZyCpnxIrpUZsB/1r9zXDG3
wobQ7ANKQXSi5KntaucPQfxbeZ73VcMeuLG3p7bbJ8fQqndAD3DkF073ivy18vyLzG2u0TmiPabM
nhMans1XDEyZeKuZf9n/LGzHDDFQAFICOGEJpGAmPQNNdnDAJMr+Lq51nsJIqUHnun6jFyElql3N
0kwastvmlRSA8f92/zoXAqoHtNgMsL3R3H2PBvobItQgDjrWFqZVcsfSIYgaTW5eTL0eqC1g6uUT
iaBGUzvH+tGhEDgTcanNqk+6/1rxCUhuFps8Bq234pgWoYqWoqvKqjgmP4nS5qauGBtJcBi0LRg6
UfqMSstLZQ0DVqAhfjDxhrtalok69sEG8C6qhqs0gtkcHCAxq3pd6ZlNgKaBbQrO/5/O1MybLXwH
ZvSNJlep/XWpJl3kQ9gXUAiHXK0e7/He603nxWHvhR42w7WVtNSJq0wYWzX9mpXXfR5vQQT4xEMT
D6W5KsVLhqg4o8+DpJnYk5UNI+qUgobudxAUvkZzlnM4rCp92yT7dYfDqvQ1GdgITaT8yM6QsJPP
Bv8pM1iTDI598tasES1nhphUd81dQxWVAgSpVsqF67Mv+fZHgkaSgGYflcld7dw5BA+NcsEDcimg
6iD+2kqks05RAq8BFAXmW0kZTC0Mej1vlVfJVNnBXk80TwoWEzWZdT3V8Df/yqYjOQbCcRwB/MUq
mzBbJn/TwcTNnnQYjmACFCsksFg6ojIwGU2NcdQaetBPkUZKP/jqoDNQ2HRr0rj778fmsT8Mgt1M
7gM6tRpQRneFOYt4ME4neHAPq6UidRN8mHjXP/l7t+grEjtC5SB2pnKrc0diGxB85ZJmGWZMewA4
/OVP5VUpQuuIj2EPALLLfhTLL8b3I7uKrMbN5bPnxvL9DP6mEUWGvLwvmzYF2z1pn0D1Z6a0eCBx
48+CkP3/D7rZITrVWzkf/xIxPujCFvkLv6qTDAyS8QV8UvsBnQc0/qKnqibCD2a/mD1PltREbob7
dnA4n6kE5lZ1KXqodoRmN9VTGA6ML5XbuVnoOYq2xKXDkXQVewZ8GncM4TFIw8zZr+d8IlxsaRgp
t5+MnvKC3ANoN25IE8tjW4nAluEcuazHSe6WNR04+rjGPrIDymMYpZUF18nXmL2wLZRf8geypAw5
5krTz2I7P5A52Dzvq1UfE7U0aDmAx/1YzSU7aJeKFl4YG87FQBcjXvqWz75QRv2Ly1yqAT2w56J5
VdJQwEm9MXDDyJzh0A3GrOCAIcKS+Cur/Q96224r3qGfHwv9uz7gB4ZtA0JFO7r+7N1F+bB3GU8u
Z2H8/SJg/4qAXlr2yisZPLWxBMjsRCufydAPqJ8O0I3rsvFG+xIjacp2EZ54ZRCLe/1iAELecQlt
CvY7QdPvWoZRg2f8oWJ1aQicjTryzj7idfnDyII3XGgbkLe/MDm+ikjJxE3ym/Tp3RYwoIDzhnce
aGgsuc76FGN93wZx24Z7e3qreE8zns/yxQwNe3QQlBaEXoOPg7/1AObj6tn7quHuW/yZv+rh9ymj
ivIuavAB75tpF4oVk2xxxKr4nOSMBDJvLnQg5qDKqMe/5trwhCQlJyb7Hum9TPfmqRIjyRDFqqkC
/ysOv9O0SBupsOmN/goDOcw6K2lb/EzPD6hSYfhDoEb6G1ecAFVzwe0EwvGBUB8yHPdmcVMZ/n6Y
mtlQJ6ISO94n8le9/YE6fY2XxzwIHq7JXSC0DmZRqRV6E8ZcfyNVByNebyn/CW8zPWjC+rE3e6ww
dyg/V+bIezBGUI1ah+rSHnl2CDFMRWdbrL5LtWLkYQfPCoVMdEJjv5YyTD+S4kyKNgiC5N7EoH3L
jHnW5N1YGXbJ04MIWLu7NAistgW69pgaOdVTrgK62OTOlpJ3WroGfb+TomDKe3oMsqODMVuKXH7K
J01a4Vaf4a+XZ4q90DY9igw1+UI82BAuUKwORCa8aqcD50W8nbfny4FsLAw5wrNRmrRlRtdwwyK9
P+/eqgWSHfczO+Rc9SGvu86WkufjQUu7pcdK1qJff+XEf5FbghsbF6xNlHhg04qtohghpHH25Lgg
pVJZXJgA9DtJib5Oo0+tuJGxxKDDewaJe4AcPhkzIkYscNr64V/bAoTtIVFx+iUbQlt0/ZuQZKkj
JdXP/w09BN79RubdJ/8LSgZOMw/5OqWPowLsJcz2Cr9LnzHtrFGxJvFuN98QqwmIn1p0Nr1HqSbH
CkFBEwuAt7dgwvx7v3OcMyUwOdlNRi2HDA/abNGI6HoA0Z2jnSHTbwHhtQToa3Fy/utbOyY8X3Mz
8C/E4eUYDvz75spGymzLBzYZZoJqWd99WcYEFWeOuLQ88RLNOSuGfjD/MtsntqlDfzpU52rmK0R9
/Jl+L62I2PcxMLybXcfv9zbFNKUk3TYPSJaY+1DAUl0Ghr3TubxiktBcgwl00jKpPG8z+PUNl/hW
7chDJL5dnHV6fiPO9LtyhcPGOYqUfwMVcBKo8Aaonf+J3IIKfAhVPSzD/an70XHhcm++XHiOoluP
J2Q5mgExt3tb6pdjZzoOv8aDheOojsnwXUvnnsGursLSNF7JBnmWmKQ++iJqMDgkSwTEmut7yXnX
+D/fywveq37NSS+eXilUo+oLHQ/CkoWz0ByhKpIRcRWyTUG+sEEQTXWlp1aMfp0rLTof41KRovPp
D50iY+4snNUOCyx1OmwJLm/c3dXffRabnbtNxVRA/3wepUeu5G25OK6Jsbb0HLYIpMvdqP84g4kP
h9Z7oSTw+vtv6TKhYgJ8vWXBsBGrEdw3cGUbPRosyjA0OgR//R/oxhRoppi8l3Jme+rChuZFN50a
ht2xsyX0+3j+e19nAZVBTgaPq1WRL20lq9OvXenIueOHvl8TWZL9uXyFLcCghdT021DhhsUfedmZ
urDZkSBRqrD2rpQzdFyl6qRJStNkR5PEhb5iNlSTcLBuE1om+R2gibt0bdbNPzjJHRojQInw3j/R
kcaQehdL3iOJJEeyaCGy1AdFLn9FQPJu00qLpN1VMMXtvr/Sr/j5FZBpklyrbi6Q4ueaqM4Rkj+d
klod4CLRcAhb7D+77n+lASDAqe/RZA72Za6IlK4P4qbl8ndpm7ltox7sK21fTCPQMScM6Ra2adv8
08Ri+UWPIiJjCoKQN1bUByFkD5YpV8ft5pwji7oGIMPn8Ruk9tzGYC3nrr8X1rYBbodY8P0pNHcp
DJp7Ge8gQjLcfrr35L4VxewN7+D2eOmho2Pl+lMrowqAls34lly31dc9k7a4wT4RAmAQ2pR0mg8P
pwvBrZ8YZOeFKRsT6CzND6QXz1MH4XrxdumCN7WcXVxj5/we14GH7EgcQ+XWE+U0/b6sDaRVlpq+
Z6/kWbH4sORrBm/q6qLS745YyiAlxQkj0t/aKcYn7SsuooVkYodR18ukKZR8XQuNSinFrIIeLpqY
0qryrFZMOEC98Rb1sbRZxvTDlq9DHQ8VgoGd3DTDaQml3n0S80u96tUZUfkU+iF8h6T4k+giMBLl
/SsrttI0rZdNHWQlIilSvDt9SJn2M1B1MRSYL27DcRtJHwfTcqfu+5iCnzKuqOVhT4+Fu3cIcOff
9Bj2MFR0fohoweLtSCAff4u2ydUyVFmNFbhBvP84Yi7YQyZPd+yfW2HH652NRnbu0zO1iyECfIvp
ZlHMhDQAWPdH5CevV8AAgtlhiWaORpeIXYhLZ6DXLMS0203hTOmNgdkL7xHto8UuOvkAuwdwt+40
AIEH/2jWOI9abTjhKzpQ1dm0J6JGn0TFZiGU2MqEWNEaSx/almmCOt2hEPZ1Iuc5h0j1E/Tqfakn
iohNkm3pD3+B8S76ZpyOU4AvhotLhTywaTndog8eyPxEUUXWnCbjZbZGupgJCf+0m9Yl6BkPi2ak
8WOrnRP96Js3ZY6cGsJDy2mPYZ5BfIKzG5BnsSfVzZvELBUhibWm7QIhHVXx8ma0b7DSbZ1K9s20
thG/T1AHFtNnodE8dNnQuSMXbHUVgKix9D+MMNqjQxUGMsAq7485w1QgXAslaHvBMkAAyTaCsvzI
hKfA7aAOJ/cG5WPYr9SdVyEqIHhA5lVpjL/K22q9bVdO33WG3VvCWkmkYKGDFKQCIKTTTyU/SwXw
U91+jtjMTEE5rfw3yJb/N9mEplFmhhoOj9Y4ixlTpM/Mwf6PamDeaMvj3pUsOuVbvXoA3mL3SRAL
e1+2+EnN4C807w5xpSHLqyOVs5gNmgxzP60VBkd010LVnynzml6HOX7dfp06cYDpluQqcwhxEke1
LeKm2kPKlEHFX9ut1L8u2C1+BL64i7/Zk8vhHlYZgX5kuXEdV9UsGyI0sZoJdF1PRjL0aoY3Bnr/
nQOkKVSIK8jeIFX4H4ghOEegdP8gbP23DFRBdxP+XAlvykezj2dV8MpEqq4fZhxExHqm0VbwoiFi
+O1mGDrxfGXUuPaJNzj3SqyAe5bwlWuKKGfRE/T902dxX7W8q8vek+wBFh+aOwx6qFlUZp2kOWXX
wj2Kh0iJy8FQiXUl7QubHZvHVZ6nSEFpZUgmlbTMLXwrTrfx7teuSwXCrBFX12bLMu9efKAnOeIH
0H0Hh8LJyFzJdHenjTQncw4b4Nr03sJXInf+iociRfCcgN9ha0HODcQPz4gKLtxZBQ4AZeWt3mTo
Wf509SHwdeWa04KxXDa0+ko9NaEQsSsUZEx8+LB2Jnmj6IJu36qJ5jg8lLM6LARlFMZDAZGgR2U6
aVnlNxJUKiw/XI6BjuKGDPbZcOVWEckaCFBTWi0ClP1VK7MyqBKXK5k3ADZsHpmQd9QFZMj+5Lrp
rlZdFRzlW3QpAPQpwAimBVE4AMViDLeZkqyKAfrSFutemP8HGDFEjkKpDEiJHvBJkj7EGSY6AMkX
923IVQRU2+pHXPhjZHjrPlUdllTubN52HJwZPx1SK+mSGiN6dif7DcFTdNW9prnjkG8JISDAx+3l
ZlxI3Y7adpelUPF48PG5XpXMR/mBH8Rg8FsxSujYibjHB0+yj54Xf3ZLcEAoMBeaYBb1WNDbzaGg
Yz00s6CMyzH54ItgekEIxFyhgQN//ZAbS058zLu9gXaL1n0yAPp1Ow8O3Tsx2estDAgv7wXQkbIX
QPzx3rJ7okj+hA2mdVr1TI66CrsqvogAzYJsVRFRA3FAqyMx2eRMvumN+Gfp8spToXy4tDZbNpNd
kmeKAgg4TsfvL5M6Rwcak9fc2VhnnHohJFkt9tFL6l+c7m62QC4D815K1HC6w4w5yJ9j/8PZPbSb
ZliomDkEFXaPPzyoRz5/9YLnYhA9x9khpaKFV2yJZkv5xx+7hrJO4AQ+q5wcnGOJ/04hey6PRDKD
jBDcDnwleyBztr7hTQcBOjuHkrpcbs6pxGCwDRy7U0iCgwBG3Mpn3UQsuL+SghlwHbiG3yBKqSj+
iRDRo6MHla3O/+vGr0nq0iofr+r7l98LOVogUHQhkaPqd3ImxjMxZWqXZaTxecCXRW6R9mdKHn/W
um09TCR5nRPCU6weBteCERSoCeLtR7YlBc5a/74eNRNbXosH0mYvdwhkArDVvUo45CB6FpOypDyv
NLmvDbGjVOyITj/RqrJrpJgqDlSn15bwh2Knb88Jhj0rtFyCR6l+Tl65X6vbqIJ1oz+k0twofoWU
2TPDiHBUb184AeuQqx3yz90QQjnS7ktMLX3lr4V5nWiW/FBaD/D9Imvj8ZIl/RU2XsUvxER/150h
VX92DWhj54mfN2MWZexES+h5aiHVkJFGOoI0mVX3DSUjgey5g6Xw2KAqNCJi4JIIqoAzhmmrUQ5V
4j2TDrL9DDNVoo7L+6UtHtIypPUl3GT6i5TZCOHzM7eIzkQU8khcTHXChSmwEgydyGQyjyY5N6Kn
B/S4NtCAp355rN+BPFyv7c4QUMuzLkok01KGbkqeMDi92T4LyeE9KR8fMQNn4Dx2mo5iq6IGG8oW
4P+gocRVGb5pBcUZP5nTUr/4r5oJEBdO8NgPMmTYf1+dMBe8RrZyqiC/NLWWLq+hTM5G1tk/oExc
wCfEClaxgPkExm0ZklCwWU7S5K1u4Nr1IGSqCTsDN6CM61LdbSMRe9Ul4QUS2RtLFTXqVg1PYKQA
vFQpDrDlzMfYGsWsFBmZlgoabF6jJKhefxxb6+mJNQJvZKuq+8Bww0eBRhZIh4hXhdYSOB8mz0m9
G6Ve04hqLIooEFPoxWz2Z6KGsZZXxqYUXUQuUBwfb5pnvtQzefOzJir7bj/wW9cbjYLCd9gdDeCU
GCpGa2j/DczuaAN4q8jibPDoCzjiVjLKOzqzdH19LJnD+BVNFxKDK20Q2xYvmZtDK3vuQVtfw5XX
/tyrduBWD74Ge3wAd6GVVciHgF+N8BfhjSAn3N/GPN8VAkw1RRvUe8WtODhPNedLA+lxX8ORZP82
0/eW1/CW88wPzkNwgQBiMQ8U3mo8abbHo+EJfsTLcfJr/SL49F8VHpiA05XWOATAa4QduxXMQLs+
EhM0FOFg8cBbbZZEp81723kwMHJVU159TwdscbGGwlgUARJ9A5jeX7O6542G2i/ot5Z3k8wBCM4v
AR+VG1lXgoIHJCfJK02V80EHgsIzYQ8zSMWm2DJrBx2wkyOXqVZ5va+19W6IvQ5fP4YtuQSHxdIg
3Xf6k+vaOyhp62lp2rRM0PW4dpDu20n6s3mxv4WWnPx0XoAYGJEKU082f+R8rE75fqFFiw/xoxYg
mxFC3/U95KsRwFghrXC3ohMPJzY+CKtyz5m5e3ZkGh0i+OPi0nOFslYwNhuLytcMiGVUJQARDJ8Z
WwzObHA5DfO7fdfJHLeljly8WXIiZ5Yv5PJpiTE3Mn79HCP+OKiAnmzwR27VHTXiU0p3vKzsFpSg
gS1mLMeh2fwM98jKB1xAS4g5XOfdaar8uX6F5CUucOtX25kIYaFaZF3m+PBByr2m1ZWAGK/E5oQQ
2/+HZrz7BLyGEv+tMZRIpitlNDW0jIjYGqkMpyiNVf2VO8Hu0/+BWZG7CjeR70+wqSbd3W5CrDDR
d2SyTES8is1eUGs+Qi8ai6a7S3nkSHNGwkqTuA6HZOoSCnhyniAJkSumenpiawIq2Lu3aSexU/MK
+kksTiSHHiglRW8c6+01LAqhOHsiXu9NUU4RSG8i1C2MkRECpSneCyqURIk1DLDccXO8BbXh/UkC
ReamssUZe9J4eFOTwgHo9lpycK5MYAYsJmn6zzCEOu/BMOCLsPPsXJ+YCclneBKwtEdVuNxA8u+y
4nOQbvAyZIyQ06CDvlMYSjXVj1lR0xQYEBXuy6qJRyRN1X1FxppNXZJ2I/p8v3dQhXOkzIEeoshp
4JJRLEgNGj20yFDvrsqjMLIIL5p6cBC61wecnd37/gT+JBZ+rIlpeCIQrufnh46JtMLZb0zlFA2P
vyVvsz8Ot03aPqXRNJR9GBekpBc5MapvnpIfM27UqPsfW8Kz5ubK58zqB41M6zNoaFP/ygIC5Amt
O8cetgCXKB5r5y7O2U1shl161adFSva0X15Ww9Rk4t9yS4QitQpUi2k1cfN84AAtt7Ygiwb1YXB2
XPkwjzLY93opk8dSzLu6+YIQEu5q811t9TxOPmUvBhXPQgmAYmdLOvM/1Aj00sgOXeP7ua4InxH7
r40r/fJntbLgCFMo0zFs2S2/W83gqVcS6qSKZBq+9FICvZ66XVQzmzPzrG3xIG9d5EwcH/3JsvVH
IkH5TjozM6jK2WQMpN21D0aHaeI1G9krn6CTsi7EoZJmVlxlp7CukF8X507jsK3+BWAnRVEz84fr
1MNe1+XSjIxwRakRkyNyLUFOqy/Dj32Rvb1FT+LiMQWVlF03EDRAGX02q0QUd2wIG0MjhoRS1ieb
awXvzQS7MPHsxyxAGPv1Y3CQQdDyL7mO5Ujy19VTRyHsaUhOWbkPLaNqkJyrlQx8uMhfTVJIMh6K
2zJ3airFsBrQUKeraMjgTwwYB3y0+Wgw3gFcSJ74XVtTavKxrS836MsOvdHlveULNXfmMCygv0j1
CBTeDo1L3hnaO3sRV5wnRfYuQrgcwZJV0mfgYDHp6Hv0AAgcu0sJ2BC3MVArKrVAOCkdTyfQG/wm
HEw7TpryD1DIGr4V6qlH4RMkgTWRdsAg9yQrc3ZM6qzHNM7+JC1/6yi7vVl2MfqBEiNjIjz+wcJL
lEXuiIlGN/0b1De3wdP/osK0WInJvZFpDGAXeBn1NpJ3KUYKvOn6LobJC9mW/UPDGImqIivhoRFu
fOOaIXw62ARAY/zbRSNU8cgrUMscC7ziEYuz3AQ4plx/saqc1bY7dxbu+CCvlW46rACAaNWLxmKP
50mTkffNFy0d1ONepPFcGtgtqprtDic+dB35ghe8Xp9utWr/g5WdfX+fMRpbAnfYFI+ggaEQOyIV
wG/GZ1A7MHE0/lGd9AlCudXvMqhgpJKm4O7v/KS3M4MTIiuxYiRnOAVc8bMx2pg7gn39gX6XfAvR
UWXz84J/3M0nqPm0DYWFyi30O8+HcocShK2aGuI+uFeAQWNVw4roPnRIrXGFi4mcl54YLR2on9mf
XWc2trehcHvGaNI6AyQ+007CeAL6/L7ZJhGOY+5LBLBl07vCOOynsT/78xEMRfoy11xyNTQAvxfx
uqyuirdRtehb+/x6j1JKt/4UGEilcJ10q+4oVE9FXn4V0wkRZF73kdjaqKL8J4hhYJYBQ4M3C+uO
vtdYBnNMPDPMSytqk6DUVYJyKCxJQOC2ZYPb45ppw8+gzN7S19We5mdVKBEtgZIuv2lTl5OORXgn
i8BR7KUJhdyk2hZTwDHnD4Yc2baAcZ47X/LqQVQl/moKXEdjB0Tg02X0KHOXmSVzwFMo0V+5WnNp
NQq5OWNkgkH5gkXbp61Y8Po6QXFummw8yJS+mcqB855ZYJsZ8JTxC+jXgBWisRwLq0itkJiHrPQS
ASdYzQ8NGh/x3gQ8S6qFWQWE3MaG+6KNaRTsXr8zGs6EsCG7giK14/PVGwOdjRfiILAvDhbee77s
48XSbPpfTuOr3gtItafKUxzBulJ1Lf7mSXsf8c4vjyf1teK2iJjacTzdsMLfH63XU5mNxzFyVJ58
WoZfRCXZJcXwpDoYmukZ28fnw1EhW3tXVEaCQvM8qPHw/Bn5WDDZCjtQIgQ0JyVl9YMR61NuTly5
qb+bK/Qmm6mWHejJ9UT8s5Fj+PpfxhbrluFN6nfpuBjmzPAvdg3K1XgKsdkXtXc7JkM8SKYXQCUt
SESLU+BvMJkYWKoxdOpIV8dVqMdqfDCFjtxByaMhnqH2VwIScWHJ3VfEBKRLaMeFCK9ir0aVcFIv
LMQMUCcrAfuLTFIQbR7bokkAq2XCwF04rEG7bRUIig6Qbh+q7nSQS1MYo+QmvDiCuBXV4WtE+PV4
IMsiKRAut/Qw+ZU0p7F6skvUYISYY7Fgtb94p4ClHaSq7SjHOA13wrLwlvF0WVr9x+m4eygURyyl
ZguGHUE8OoDw7KWsh23Y61/0kWhj/XQDCRNDaNobDozqE/pWirVK0i8S9KP/gbpNW3uEvA8fccMD
/TbtYL5FMr0WgJ/VHRYllwbHXZT0ZRoNhNDHZ1BrP5Oe4WbIubbkpl9mZ+f1C6/2I+2Zj+lcWhUD
4+EkdxpCz+wvYauk09IiEZ/Hc0tD9vA6VcX3bUmYI2xGg4F7klM4loId67o8CUF90SZNahotWgsx
iiFTV/yDJCWcokBDq20wW0E3cSPbpKD37NiR6DwbWkN2lK+fhJSDig8cKArk6grxVXHXkcUHpvVj
CVau9Z2HUcQFFdr0vrw2qDD1A2oEs2P9/dQTvbXIG9QeSSYlQ7p2ugCNBrZ8fPkis70BePqrV5LD
ZR+nwWIBYYNQ/23znI4htcI6ln7V4RbS5pjRKwqkdX749ETVbAGN7bvERHgiviVQCTIF3cgVAnjM
c1f5f7jCNkCXLA76W8FLW9LIUN7PGi2ewsw3HmNwLkONOda2DoPseE9sVY4SBe/a2TGm7L6Tg0/7
VOp2zljullk9UlWV13znsIkDZiKEWliQZHnAwziP1LKaxzTe2FcWWn4T4zBiCe5p2fNmDwOLRvGP
/s3jPAMVXZM5bot2/zND2lgIHOuvScpiIv66e3i6ANUfWon6McQLxY8wfw0r/+Sllx2L0GZf0/QI
hczwyT6sE5NQpnSqei292H5IZNkoU300tTVh20qrnGF7B1AEgQz86dQSmE6Q7Q2nrLuOU+gMy98g
mDkrMKVpGCTWaqU+zbRJUidlWmt4hGTfWdmxC0vrKpllbhkxlebz1g+dT92bfwg6yeL17luYaZVY
cVJUD5zdpAaadDoCYJXzon+UpAD7k7/+AVGT8oU23W54+k9JofYKkFDjl3kzUk34sfswW6Mh86kW
FCFGpflrHlnSS4mptQfqc6PhLeCSr2TmvsN9ij+PWyvXjOC0/uVAV+luqgzPl7mHnYge8Bim05bS
Q5O+RssU0cuXPqmWer4O2ogBVbxb/u+UpQV9jf2tdWQFQ9as5/OQ6wDHaNjBGTT6tmIWLzGiljeF
XRlaAUgB5ffr1MgJv3b7G8Rl++7YEC5bWxqZ3tpxXlJPAVLbHgGuvfIyeUnpfycFfuheGo2GgbFK
h/MgPv2gdo158QG0byDZT2uUo76iMICEqTm7i/no1xwh/J0BYoPAKk5ZSIQS1SF0ofQcQ9Uk2fsT
17oA4Juj2RMny2dVat4eeopovg6kjHiHQGxam8Hv7Nqe3qe1n3l363KcPTpqZn0RtiFBxKVOSgAW
CMT1Ncm2CZUOVAAwvwkRej5aUrtZPwUxhpJk3MouFBLlaE/7b72+Zz09WNfXa6D6VTkUyoaxY1X0
w5MeQNo4xfprEy3Ku75/pYwRGwGnMeVU6zkUYfBXEbnRbwdanev8P5/HZbVAQ55Ee9AxEtaw4+pD
eMpdz/NjPSvDluQYrfgE7DiVABlRAUayp33gQhC7WfJ2z0TLwdZYazLudx0q/sNlQQIa12qK+QDG
PB8SQEd55kvDiSVofdNucGXVavtf1c5M+2Gr49nCbsNeq1gATrF1gadctBR2SkVBtyQiptqPOfnC
wXMN5t0b9mqUEifhzO/xSs8wqexByyYZacDpPo635u5d1sFntUYj7NPKb2Wi9yI0JtLuejHCA0QU
fCiTYeRlzmyR/CyXw2ga5erSKW6DbGgVgzZG5WEiMv/a1iz2ucjhfosAFmE+uktNYH5fXGy94w81
3/AwvffR2DbCvrrwfEytsOACfr5fhAm0+Dx6lFi28sZ/n5O8nKlLtt5txD6zTZWvgH6B5zBfa9qY
JQOH/XbKMswhWk/zr0yX3iTujPKomwj7nSbs5pWl3gHrm/0oY2FosiPT44qI+U49HBj/R9OAhfeR
alvuETx6ActliZJ21m5ROgRmouCxOj8/bKGU0uDLYccA4q12PnjiqtWvu7ArQLCDjFBUFd9Cei9p
u2RZr9F0f8XXOJ2PjCfJeU5Ig3MrIa/uCYxeGoleFg4lmFap6NMTitrQQMKeGFrdd+4+XHgnF/No
ORz7VeWvlZui0I+nSxt4gOQxXFnNOPUWhjygILo90BaZPDvoqNyfW9kqN+DBm5RYKIuKno1z+cD0
u27v0xyTeWAAj8BPBioFhWYp3PfAiFSQbUuM5ndoSQOO1YrB7r6yzczHxuRg79HYKTg5mgibaxkv
A11NsMDy2LhGCUX8bJXOt9F38Il+OwkQYuJ1kYcxMdPKI2sndjwTFz/RhlXHbkbSUoDpm/nktHqL
ekfYZu67bWURpNKkw7rr/2Dv4cPj1roDT3bPVN+/Ky7kxdb+mUXwADfXnE7K/e8O9BfrKRvPnIUq
vRe27euJHfP6A9+IiXzTMGVm+iLTIrNthuMD4WR35cyn9G7rkWoGLjEPgaeFBhSzgvwNeEsrAkl9
/UURvpc1304Y/3pkw+GThz2d3fgDQInr+3qIYokaIfr0btJ4QsNcklaozAlo19+FkwBT1DQ300FV
XHyvmLOl9UYi5IwnbV4AHyq/Xh93hbyLJ++FAIWVc7ZZW8yOA2WlvYS3Ab6c9b8ypSUEjXwmG0uk
/HsajRiy/IDLz2fBR5cnKsqzkoLTICj65sBzuaxjgGC4D+aHxWYB/0HHxBAm3hER+sStYwKbr+OU
bhQ26KBXizUImP4ozX61KOgegY5JkGVThbNeQsupFpcDbWtZfFVntq/bBtTtvuMtxqX3A9wgLBcd
BVQSEYvMg2/0t8KyL+F0YuH4ugme0olj+JvNT6eLxKM+YmpvdIH7trMvml3gIie59q5TIjJ1TuAQ
/6FzgcaShD+nJvjRHPNNO8qI3yb04Jlc7qXLhlxPVGr4R10+6jVBqd5QbyUrsJoaVvhG9byVZmJS
G35WVxUjWpHRNCzHjhZG1GnQLngulS1NItNo2zy2VRA09Q7O4I2/2v6m7YF604f9zGEkmhKbH9AO
M+S3qWsf2P9wkMyKz1+5wt/A19kIlZNQ3tTzbtlm+FGBYLbV73xOIrhCU6kemmro70DPywQq50NY
F6zh0xaorqXHNkVGBEIjf8z5VtdPUibTgA9uIAxSChGf8tQIjL/EuJKVp9689PrkVeFAAx4EouoZ
FtAsRpahfJvRWmyF1AMQpb5veItscW66YdxSfkhoWwmphqn/O8VNou7S2zHPfcaFNT4+3LReld4Z
FDnW6HbrGfjtA8mWDX3s+IjEEA0MaqZPaYTY4niqCaGhpJzF4dWEZxqhtP+9I3S6JDgZkLWr3u2B
NEqTlPs8/Zjach2h4KtE+K1fT5fAMjiOuHRVAr46mmNyuitbkB3o91peVipHzEWv68KDM7hMJHoO
Kf//hVXCEPneTim8W6E3jMKd8a8KhooXFPgUbfNqT4zfp/btYPepA37D9GzTUWMwwOAOBVGiDIlL
PnJoZ69jxTEZuUqnpmcRMPHE8TXeEt1JJoc+5Istkk89Ok7w9j9gJFZ2rlVrVmxeNM19Prtt9jlx
M5YjlIICkl+Yfh0DOwSr1uhNQzO56JMEWQynNa/1k5iG0BzlQtkTGWSgcXnPB97MDh10rtcn3gWl
7RtbS+7xjKOFPlqGj8VEbFVuhmBzLnKKZfZx6x0iW9Ydq7lDHELfDkokqBP85zZ1hcLh5F97nnyt
oczS7D6V0SzYW50vcaR5YbFIlNVzYcBzelO3BKNblgE3EvNddVmesIh3ebkVFsbjmePJulPKxMEh
jtRVzKzXHb7M8VDVz4rT+YQ8RGfevHpBCS6eFzhwbgyA4Kumdl0jhMVuUFYHispgfWKLj1ZTk1iQ
RRwVoF7o02uF70sGw5BtZEqiFQwiWDSP0gvyU9QWCdoUrBG2u/6gTGw5lO8WT+5Dg+g+fok6ss2r
2Ba1nPtqSAWysPZJBIcRL7EKMVBsPyNG3DXQ1l8gEbhZkklKGTThzf5RLY/6dX3qQX0HAgEIARxA
Yq/LOw/67OKKrvrt4M3ojwj5rvaK6B5Dvo78+M2JsyRCS5tEIxzxj5D5z32v7VZojM9GNojMSJhF
wMKnw7DEpRxMZHmkWFy3iyxQFKBuPw2rhb2VxIVRvYlslx0nE3KI45hYhV+y245KBrMgZSpNSbLL
Rs6umjfTZERfl0fVqi24VEZmpJ4pk8nz/ylgpAYxh96tRELiKfudmEZRf4SVuJpPfHY3VfXcKNZw
20OidSsD10oEWfqhSVryX5trug4TrMqUBwrHmMXav4Qxfnh6ryXwEh4TldrbjPL+3eQ5F7yRJMfe
wyuAuZ3qBv4MTn/HKjpBWx9wd+flrOhPdiWVCCpBqXLMv/Itkm7KNtL8WQAgk7pxUNE1tUYA5tlN
2+gDS1rRq6KSBi1XLHacfy05bXDCZ9gaxsug+MMxBk2xaouj7rGbPhzUNJzwfBeQRkKkhAT9U/hr
YTeG+dvmdbslC/av268FBoTe5J+qP1678UK8L6syBLeSthwgNf9i0XegH/Fa8B/P82UYgVoW6np6
eBDlCOdSoKjWcfiy6hXYXMtnDp0/w2PKiT97LLpJsN8PqOPMEUswBWQOJbPh5fYhcKZH272jj0oL
2gQAJ91Ipi+I6Wdjd5uJZGPP2TgcFlCTEMjp79orni8I5NeVJ1Kwcq5mwB6M5bbDyp7X2+pM84x+
ph6zq340J8gY/8KKz4t6QWQfiyDqkNpDG0M0ahwPoPIkiGxJhE3ZyK/VbuIUbOUDKLA9bYnnFbPz
c/f5Ki4UxsYBTJYlfOzxtHU4a2o1AI+uUjEnspY9pkOCoWRpriRF9BTyotTbXwPeV0Q+LM1R94nw
6MVX/yIrFEUmEl663b/lxi38tQEuOIFjXa0E6TPQdFiNTLZ3G7swCoOuQ4NWqG2Hfxt5FIVwDszh
jKDS8X9fnWAr9gGKhrfjPEKZTutsDQdR3xm2Negk6qgH38hR5S7VBVjAicA196OV0k0dkiIqJc4D
4Up0r7FxsKmk1LJiohv1dQU2NrML7h0QqDfqqvwxUVhOYs6UBFp1XC5wQxxIa2VvKeqMBDGbjJQT
lW+3f1TZzp5pmOFxVr25j6ZQFo4GHGiItMMFMMar7UrmXgmfYHIz8hn8/mQsgppuDn6IEX6qjqAm
I8iQNrfTimIA0Gd5GO28ULOXRmScVr60VRRgBj2Pkj7JbbMoanKQ6pwVYcO6D6T/O/nFwFp68vi/
fAtzpJt7SHMzVPfVfLpVHKSQEp5yP0KKg5ep/oghQdmwRvgV0DKSVDefFrNmP0J67uXpezlZzkdJ
dhtDUN7YqRbbQKQnx00PKpJii3t7G8dCUFZ+nfZMef4TE+EPiVJB7hfEETHkdWZQHDctnXMDWFMB
dCcd4jVfr5iF5wKfMBcbKX0GOKOYoi1VUmJIElexMzy7hSE0ENormVb56mxZcNvYOutd/5AXOdGw
PpMOl3vZ5hLzJ1Saxn2iKXUI5uNJz4geFCJYv3PfQV5vAz+gWvG+2NAxT/T1EDW7KUAzcMbq9mHT
B98xvwkzeFRtPi1N8uWG8nCWjuJF35+rPEI6trIigfAkBbNDEpNn6t0BOOvJfVjTtdd6y2ysRRrM
wyVOwmcPLS8U4h+oJHIu4DSfPfj9QebenQIqx/x78fnPSKzMqyynKRcEivzC31Q+AxnLPlr46zUA
+H59AI0+jmOjG77o8srD4WHDgq1saRoX2D4L2z+QjIlyeM58NpTeHI2CODDDShR4dLpfB82FGRp1
kO8GHHuhGwl09uZ0mYu46k/1/bHN2l6Gry+JuXT7sTZcEufN3W57NEB3cfCAKyZfeCJyonr2NB+L
SjJyv5Vle5y0pMXYF4o3sOWYzEWJAmAFZcerV2Go6wp1NB6BJlHfhzmxDkvlsmu86GYsGjDV4aYS
KzYfbyRVN8Sg66iPTEpau87H8odsReh6ivKB0iKhFksSY+K7NRfV9kCqaJ6XOFhsT8kpGr+lm/zt
+JzjwyJi4aPkPu2iUbUTLvWMhpfMViNpGHxTN4a/co3GpPoZOT0ApueI9rBZQBNYF3l9smYt26ro
tL+1ViGKSGUSg7OumyZe4VsSdyUF3Unk3fkaYM6Dj0Gd1vw2+b/FtE2z2odd9jpM1GwPETPNRX68
LMyxrSllNLX1gaMI7XkCOecaIEkYwa/wecDTHX45BVYyDnYe6iL7kfagb0h0kMOMPZ3ICuxJkU/i
Bc+X2XdRc9PPgd3l7riQ2nkpYYUD+E1wN8NcHu6NUmEASchJYPgb+tAe0e3QmATp5vWVv4Bjmxna
iebBse1JW5jnAtjXZCLcLKCWzZ3CUOTlVdsT9jFKSmqEJ0d71184+jbk/nMHsAZ0NKdS9xe5hK10
vDm4sdTj7IiEK5IqNCHX4w78aXZwIysVHxIgu2Z8aMH1lljjxdLSZF6P/cfOtU/S1cUK9DHXw5gW
Xh/2C955JkzkqwG5TkzAu37jwQ1J59n/rPcz+T7ieJZnCOYcEjxuo7gFuczP8+oJQH1YbwyEKCR3
x2z7RDgT42b54q4+vZ8fu67LLBnARGmFcKO2r/Bkg2Zy7udp0Tz5mT2x80WG5sDYqhPulthtNTju
XJyLHxabzcy9rVa8qTFOAA7GtCiKhIKXwthEtKgKA//ZdjjLcuUfZP/ui6EyG8ImL17BDV8KyCjU
Zdtr6PWxkJE/3AXbsGAFJrKm91Hov1RB/SbNKlKg0veayzA1X0Sv1/C3lLrUOKg7MI0RgRjiF10o
cLKsJ74Oe6kTvdhoHOyNLwSDbFBsw4Hnl/KMzMLNssRl1udYAH55mTfCXeXvh7Ay8jMWicjZ/7p3
orROx1mAXIh7Y8z1a77BDZL825v5pelzyDIMgspSg2pcgUjC5W6rW+pNj9QsLac3O2gIUD4uJ+j3
4ibqpRdtcV2RBuOrcy1lQiOq1PMy4vDeSC4n9RQ0M0G4fU6fDERw1RGGRc5uAcUuesKkB2Vx8i5w
ahQ6YtJYCHiTRz5tVj+mJimb5N1l+k7Y3N/q/40wb7X2GJuum2suZI8ZSMYtDD/9LMNoMZ3DrcT7
blAGBs76t1WYJjGrqsVbIMOe5MFFNSmiN4hAjpJXlZaXmgC8tHTjZ4ps4VtK+qI+hsD6m9z6QKy/
t+Q0M3p7I6l7utzhUpnT9iQAWDe4jCIQwWKi4zCjdjNvhzvO+B+9qhBivUQ7E49fobszfLIXvIdi
KUwXJyyWEMYmQ25GWTl15h45TmXN02V4GQP2iKZ1fGBFCa7dPGtA4TUqV0NLSvMqgej4lo6gbfJy
rmWvfwyqAveirirC8fJXD5Wj0Yz9xYzeG5eGjk24MkGV7NxJYqcpYyFDYK7+eMu1NpouZqZYpYud
2uwyd/ped3oK6mmwPaENh2nlA5wwtWdcG5cqXCyNxOuONyKjek8vy3LAfuO4D2g8+/0XfUJ1v9+l
GsEBE2FdjhTzb/KwaZPJWZp4yMlDeUJOnj3Zs9urSYUWF93bU+xic0QlqpUXuwbjmOtmHmotqgSF
fkuC5/31l1AiyVunhLkfedGJhCW2wWcw2U3cW8J6NzNOhvbKDwb6iljJVf6SUxbOhSAmaXah3f9s
sSIYIfKbY6bV8dSI7KJk11urR+/wRqgxQzWWtycK5/8mfuyv4afNL9ZVb0pZ/26NNX+3zPBS4OJy
V6N0ta94aNloFwhU42vCiAoT1aqU6EzHgeDKLEcflqPqvACZWSoJTglULyJ4fbiEOifdzPcfsTSH
CMuGXfwShCPT2jASbxsohhiOVA2Vs+39EzHMHiKkHYgT3gRDWtQXr0rwG8hHwa9qhcLnXOJPDTc/
Gk2FZhW13iBVsEIXIzELgNArMxblC/0M4uWToePqfrDCzwjoKl1D5Y7L/YAaj/yvRg3DlV9c5lm2
BgfGpt+6hB7l96wSYOF+Tug4Dhj4LfipqmuKMfTqKlALsyc5tX3E0MAIAAVmSa3M/GeHCwDG2aBa
ZF+ujO5gItgnjkoQxfOxFbuwNECqcTmdtb8JqUw5ngPNLD4VNNZNJXKP0UyaSvkBUdmH5VS3ZvGP
ExRz2pWQPF58B6u6dQhZ0zrvCmjYrhN4vVqjMo5vQCOUTin2AcBUcBfBKOT3AEz4lA683CE0gPWN
m+rHe+ASSDEBbenipNqnNX0ULSL/cZCKTmq7OORr5E5U4YhnffJDchCmFwpbL88NmDbEpKvgCxx+
+mnMcRrf3aprCTM/PDG6IP6rw2ewe5oe6xR2Ex5a/ks+eGgJOe7zgDAJ3gaqlpfdCtElynLin4/j
p5tDd/EEL8LaN0FPjtm7VRUKnArDBzrMlvuqje5aONT0Y9U2iw7/wRKA845oJ1jQuVQ60qjsXIH8
WD2bphpeRZGPlgKCCvkmde8ovL3WJ6JB5gzf27Z0bwdMGmPBMzDGZgq9j0Bd8JqiWcB5jWpX4Vmv
TVHv7qmhmGn3DYqLE9JXTMzZiApPi3AJokmco+86KrXKY9O/qHW0ugXfhBNwDb4hGOuF5b+kaJo3
rMorq7b3QRDK//pFyFA4lqm+62ReAYbGwJiOp3/6zpUCVRkF1bxKYzmmDJwqIL9JwL+fjLngCzFN
HP6kbIuAYSRcKpRU3iSFO1abIiWAGQPxoLTCrAxD2q48EzcqRrESCrdl4bJZdvwZ2taC9b2VctqR
6tTS3r40i2MHFmZKcAul5/BUg5zlGlP1TmKYfA5dTSI7ZFLkxMJT9FzBzuTOaHMh9O1n/X1epCQq
ek5jmZrK+mEjlEIPfwF9OMCoyoaJ1HMjT++ItvWDdYZ7KtWUL+afk+FvkEQUkXil8DanVXETSbAL
1NzCVv4JiQ8Hxbv77q6HHz8NpoauWATL9Lm/2QHDpcJI/w4s0cZ5lRgqVyScWjBDgbfwJneCn8ei
pHtjoAE7O+zYm5OmDOZUrKJwYKnAbdvM1zcLl8C8ZNSbXUE+STJT1byTBEQZo/XnJmJtECTQ4d2j
g+98af7wXlzep2iG/pvXbTmU9lTj849Tbu1OX7Pqz5uFbO2MO0/dWr8PWwOraH/0n27OMvThFoXz
8y98Zd4abqSXOd5gKu8Q43hdGAHDP3bu5QcvMBmEY+L6rsoJjH35NZAl8rvqTKJf/sA7ReNF/vyO
G/3URkmmsgsbDHIzT47V1J3nKhm7FogZKwh+/Y4rZhCFD2bNORgwhbft9CXqEWUz7EPu3ScG2umk
9r3c64jz7ApN+mFzyvpe1EOMb4GeMqBe/WJ4AgV6Nz395LZuXBM3mjuGA3birfK3ChhFFbe0Klha
wAZTKvN1wNJUO2sHRqw4DxMRKmigwemDPuf6Y40fB9FDhWoICBZz21wNM79r7APH3WWZQujNjdKN
pDlN46M91ONSkBR522MZq62jpua8oFDxNjmU55KKUSusqamjNOukuSHziOYP3O5E8jXLxKtzvj6G
JNx9s8kfyo8ZHM/yTW0s9bZ8B9H9vDHxWzFdSZ1r2UtCC/n1eDUfV89ZH8u+efYDDqOd27X8lpy3
9DcvO3W+cedmoOg3tEnXkJ8Tk3hl3FaalUHk8jCeKT451FlO+oha01yUtWqXa+BGpep4GCSJl5wH
yiSZr+h/D0SELIlFs3xPhQcQWyw06AOrJiH1Oiw3rrXWmhWWFcTqsBpB7aoIEq1d/WFLqJH9uSnj
2uV8sXSnmkEncfW9l9QpgtUArIws47NaLnuRiL3BKCdh1+6eZJXasRDLyLqZh2dGh0dg2SlGhRlg
mif9sn5Hhp8KLfzTBbHahAY4MCV2cXCKhSi+qaIVJzCi5fiHK87uGHrqQaLyjYKzCvwjg87yJiB8
2SyiUcMEq4e0jdxz4JbT4pWtLMo4YBTTtRnNhXFVr1Ro70LvMen7kBhQmhQ0unGGBreDigxzOmel
g+TDxUbHrNzs0c8zey7w5Mwd5lTb09sIaI8waVEtXdRSnJ/1EI6azuSxN6VFNA9d6gobg1Om2aCO
QMSmBJ4xy3dMU2ANxkhQgmbrInlGeilkwU5tNgKWJM5S+NkHCaJfNELWLUIk/4cLr1lt8IWWftpn
pL+V4FWvRSp8gC/XfqYMeV1ctE/GAymT7U1QcRWeJJWldarjnWKlFe3heidh4NjdedThGzQ9O4Au
AqOrhd5FFrRSR+29mYaqS6NaUd0GllpShxZhVHsFe98foqmouEX4uOb/1nSjGG+sSuEObILzOcVp
GPRikH1Llhft92ECNVzHgVS5yZ/VpilNBNWmXw5psKixAV1epssfjMFhMM6EYjUsAr7B/aehQuEo
RWIZJn3TtBolBuU9LeOozicRIn1uKX0ZeCRp8uAayD1No+5O9kOUT/5ZIQ349ZboLXKLAFl8cM0p
3fo8rApxRLoeXxIbsO2sHUTxnOee7kX6vEnJElrcBRo/Pz+z36Z+5TMKtDsb4OJOEAgpmucfZVeq
opiPzVI9esUJntoeRUo8Xh1ISnXpP2lZjb5Hm1r5YIJVhCMmcwYxrju/Ko95e5Alia24N67AxbiN
yRe/YmWhnUamlUgUeDkEodUAbetHfW6QBWo9Wlht2ilXf6pQVJUUw+rycHuEIhf5FgZcRrgHR4TK
qww3c/KLkwF1T/U5zr2zeI/0SsD7/kWSfRuAZF17b4Wvusq8YxtTxrdTxsfGsdb7WqphfujxnYxg
hPt2+2ugtuIPVgcI9c8dlE+TfEBWG8qwFzrPmIQmdKZSYM/69V6HLx3jNcA3KFHCgZjPC2tfauKl
3BwSezFzPfnKf8sd0NBc204hKF+cG4oszbnAqYwVeT2bZhQ6zVHOLeLHaieqrv6rUbHsGCZyXp0U
3tGYp0ZI/DKMCynF6jqdYvFiZLCNqss4OV7trkZQk3Ia1xPfL15IfexlvqNGyHVL9tVjPBiMXdNw
hAriXjrGj1yGGvyEi90PmoLNzuN66BBDHcznsLaMSBtJz7XtV9YIcllPE/0vJIfkY+TS+jS51XzH
Jp7E5q/cWkLwZOFUnxw//xkwP28SH9I1OxbXfqhMX7vJrEJ+Hzo671VE2UM0svHTWTAWfffqWgdC
Xs8Xt6kgXR13EWskGcgcz7X8m9VtAqrAdcRSWgf7H14VUWUMV6PWUgUGO0S6vPgeN4OLv18UerU2
DBcK8qFw6JIYI17o36o5pcQw+cNe3UEbALMqhZmyD1l02tI9WG3LiioHD3nNzOZo2jZyLoKgmrhQ
Ig9Lzvg8K9fYwWruUuHVkqkGMoCNBvPMWHr0D19q1pxsh+uiHmYKOnDAuOnsgaJaOT3lEHncXCD8
HEJhS0L2ycJDx71K0ajiJzHXielkil/8S1EXfm4c/Xg0PyahbCmWuVLnA1ZU5bZXqB3KJsEeAV8q
vn1jdTRawIadI5E/5/iruzvxo1v132c86pJ4lYrIPAZuzLqqTwcNFmQPc7L8+RC6MAce1xNBhG3y
/p52nwIYQmzoDmnm4WzGVxIDjVanDvhXqfIhI8dmK5JXjIi8Wctcc91amTpCAT2sotR/R3/a/JFY
QCuczp+mGDuidUix1lcdfC+Nu51I8Dx91r50YeQqEA/ZRpVXhe/jRtD157aTyjVJoMwvLmu8Na5H
M0N7Ex2geEdJg3dIaCcJv/n+0i4Erh3yGK4/mqh9TbRWd7Gd64ZGCD/VwDonMUNS2A6LTUTEg119
R3LTsMF7jHImOsLGLzLju56xXbZHhV5r2n8j+UnE6D2Kzm0e+lQ6IWaVZ1sZR3waQbiEButiEUly
kKqUYLiIdPWK51EQ1g3/LUYu06J497bKCly2xJuwFqeD8RQhSCYSoYC2Es6xQkeDbuVyhGju1mCJ
pmjeYdT0cu3+GkxEmbt1AB2rIV2A+EYBykBXJuNwqc2VXfoxznOZ3F4szB3Z7Q1AM846AO/I/LuO
vMBWFqTor5JQD37s5L3gM5QevOqIppbg3usWyenGGw66Uw+EuGxhZbk0Orm6NdoWid/3XVoK7Tbv
73jUmOepz2Ro/n9oJn1gpskyqKDjorlM/ppdGyzWmNWi/VfLSEPJaCq2XhG8yYRX4qK4dD4CZe/O
U8hDeRJ1V8V91N7PqH1yuZmPlpuOCu40bW7ct1klI+1W+luGbZbxw6tiE4yxjQqkvAsuGh980J5p
n3aEuBw+1Ws5ulyQv5jH5rEZjj/8/cDXASAKMWt3hZUiBaUH7cA3HQdYbgkGtyBgarTMInoApAKJ
ceU3kpN/IgIof+EGTr10x4r031E4fZUuvmyzGD2DpbdV4dnaCDV2nXwA454rWO4pz397hc3+tb1W
L/FZamZvJJSmx4/LniqBCjrTZsnu6vDOL76aDWa6nTmrsxV2Vq6ZYC3ALn5EpyGshINWmZ0Am9HR
epTSmunot3+ywdxiyMOVD5L4tVkQXbkLayCwkVUeFd7eRaf68D8lOKtQK786W29xaoNC2CHtJQVl
ohVSOh6DPLfxYVFOSN7KzQJ9q2Azm0fTA12AEd6QzMtb386szkqjs2mpJvgmFUxsm6snArMWnyjS
7dFh1PvH8qpgjHpR1c96Q/jKd6/uMKevMDkhV9Xksg1lU9KMJUftcmYCB8OAb6z0I6Fv1D0KWDCx
7X9eUOMh0nPb6xIFiXoBRjimZG48iF2LRFdv+yr6zY+LYRtrF+yw8O5Ln6pm+pNQFNBktQZpqnuQ
H7WUmYCShuO1XwlnMn+rEwHu3RrMzBHT0/mUfnkIOx0pBWy9DECPEITCnVS2v0hH7XShk1YeyOwo
7vSolqWPDgmCyM51QByqtDDd08o2mFl67rqXwCki7BSP7wAaRPanZ8DcWdRK8At0vVE4YyLnscbb
qhaVQYTKHc1u3EWqbXO/6QDK4kBv94IfS8MO0WHpyvzFrjhntoohVigLxc1tacRcNuh+o4GiOurp
TpIQWVS4GqnIwtGimxqiTryChkCk04hCVirYPCMi2Q9t/PVgNaZwJaPWkWEBm9IrSZZPlopEoY5U
6pN/UHFMVLQ2SSEYSAMJaE/RVdDrsOVr7u6qcggKVwarjbpTOug1oDwcwWsDMqRaRCUefEIBSLj2
XegZXlUpyIv4B01QYxAXQ9pBzYlDoLYIz92wg97PGY/6j/DUlcPYYKuH6kxP+uQ/j9ot9McRpSkq
cobfSlpCfur7QdpsZL+SnXlTFz1tT8wkMmYbC3SgyRw+GPA85rvefH5xPuqF866r0cJkcKqFS5GM
p2IbTREaiQjqkS9IqFYYAg4CS7hr6liggvYBW8U3ijyqHRATm6JsvJZ0Oe4Vy7bWVLPoWsJCLGbT
B2N/7XxeKsvA5fOr+PHXIqnEbCU/ULEZLuyAmRhn5e8IEnjdjO/avCeSy7QGoeLjt7weNE+X0IBj
xgNiKaIyjqTe+Sz4xiYZlhtDhVvsmkXx68U+QbsujVEXJmzb7q4RTxW48110Lwdq4IdefII63lwR
KDPUHtRSO9Zpug2tT4CYworUJCwHlrmx8QTjoDAEKcILV3D/ybAhuqVJAiI3LQ1Rvax5sCPLBqHZ
bmRhXRHrMJT0XHCuOvJU/3OwM9ylcyQ3VAkqgRmDbsmABamy6XJGXD/5suuqW5YH9bAookP1HJkW
d8vOypIliQlVa47w4repupkdYEKIKsKroNUyUV079iB3Rb9SwiQ9jND7SE2Z2ww5rk200JuM9s0H
yeRQT4eKwvWWCnLIJw5RMMzkHF+J0l/+mNWbTILHGxUrKODldZtJSFH0KQ9Nlwmpo0PiHZsRViTg
GFtvp6TWfZzV5b2bIGrrpWpkhR04goWoOgFgTdIGI4XLIaLaZq5re28Zp3SdwfRpZMeaxVbb/Fli
K5pDlytZiHQbi9IWPLodcibkoJzIkX5qx0+80dzM0H+pgNtSGH1QiJYl3tcYkVnzZ+7Fz8JCVPSJ
1WChKG3RQml5yXkgkxVKo3eQQPWcoenmeCj8zlWPjWc/cduRGaGa2FehHnzHUMmJ+wvv68rP/7BE
Gb1vl5/hNeJFJO4bpAQWojmqKq2stIt7gtO5jABhxQfubTil45h5a6oDsl0a3gv9m+e1Sd2J7jcI
r9Em+fz+ezpl+qhrZefBmlvHxsR0yf0AVzQGwuZpraBADibgdTKxek04yNdLKuaMy3hiTcSNiKM2
qzJN7e49aC8K083mq9J1FsrB8S8VJyWHIBoi9uw1TEtghodyYVDFiizRCst58iKj7d+edmtWzq5A
eJxeHkeVyO+R6BaPoPP5m+uEET5gJBbNhLNNitHAjBTVyWjwT/QAl8weTKF4IOcgBRPOYAkHYmz+
5sK5pKbSMW0HoAvqjCtaNJcEhcUsro/mGPRmH9tH3eN1oAzwhvpNwnNAKB4KpF5htaGvoEVR8m5G
C8E7/mJgIA0ruC1vS/mF29zSlFV6PVZHCi74Ht5HJZmjYWjqgwBbfTW8VmZ+NKCe6TDginTSNVw5
m8Q11L73KPtxB8Gpulwh/46Y7M3sJw11zE9aTESg9au1NxKMubzsZnQoiyJ+gQHkS5PzFlKIAkmZ
3DQolf7P+ETEoTWVGQchA3MZezVKuCL7bpCC/WM5qz7wxzP8SwJPGwxaqI88k6yKW0BgyVksEwGR
YpfJxX6D6rzSYwM8eULVEIvc0gir247F1xySG4yHfogOclqCGyXrjiLIHovo11gjiKLPmMtResUJ
1txJEN6S0Hq92ADqCIs1NuGIMMZ2i+rod84b+n4vEZpNKSPDZjPNEx1n2QNKUS999nlVreRxP4X4
3jIBFnnWiFEGUWJ/7Kp6pgg0EWbmq9x2ah6bPp8Kp/0KXqFc8slLsNZ0ykW2KapL8n7wYrT9I2Sf
KitOJUNxJv9k4WUcX7fdr+v4JBksWGEoSF6cXqIRlUx1MSDRHb4rU3fbQ7NXNNA4yk5u+FpmQJZw
u27chEQ7VFqnAkxYbiRTvv5rmJbCD4TLPyjlNdcvrUj/5Qh6OB2X53SYe/78Heb0uQ/3DvOcUrIz
Ww2rNDdydZYuzRDY9aBnk2rWCJ2f0vb73/BZsaDC3qkQeH5DJCHKOmC8tKajdKa1MC8fTNpWI5PR
eIzKO/h3xfQ7pQg9R30T/aMAiiePEJwYZGkyEYre5rz2BEcbzhp09e2BXQQ82h94n3K98kc6jf6g
PNFREVBDYWkyUuUH0qHzw70dNo9XFLB7a9fJG6R1p8viOkNrqb+/YNVtWE1yO4WDuelr4Weugfa9
LGDcUzDPLVCg3L4ohGeCuqApYw+eseZ9gV596v2pw2tEiJPmpr5ilpDa5gHdAQs49pK8Lznlxzob
YuqKpJXcKmeOEjt6rOPasuvb756Lrw9KZNvNRDgFg5J2eeqnaib/U7yvZ9CaOUDokdwz+fOC6321
tokZTOYQ/xMud/96JlIfBN3qS+lAsfPp9rvbsOHrHhrLdIsVxO/tqQiVS+pUm9d2jyKa+t/77xn7
umvaPwmhPY6YXCET2vT9x7tFiPEU+PemDSarNL2QgLAtz04Aocb9DmRVX6pQOKNh+GDTACu8BAWd
tKko0LZZvnPEbvU5VSE0ssQ6kt5Z82nHV2NdVYOgnVG9yJMNyPzCCZ9ZBI8COCEu6SCuMYI1xDr9
mrYpq2QtNOn8G7v/vX4UbVz72kw7FZ6Fz505G3fVliBmvwploqJSfWkY5+S0zYpRtny4ckFCEvJn
AcnIkJSmmtFiEgVY/kLKnzyMExXtosxCHXOjw/TXQu0O0HrL9bagaetRuqkjHpf4qhLGfw6ysCBU
yPZGt7Fxh2ca0ebFYFwnxPEqIkHBfVm4DE56A5CP5FYHVGCDTiLj0B4WOrWzY+rXRlgxa+rY2+Aw
w6/CK9GJt4GDFcBCI7WpRBmrEbYYCWo31CfeirY9kDrjfvtesHHrYvBYwA316fqd7GkPEShYeAHG
rWZqB6/s/0zml0ImewXFw178C+EFI4/DuZYRiftMGwC/Oa1d2Q++t1WENtxFBYeZUX3mC79Q/0fl
HGQl/DCKChsBmO8d7lGMqxVFMjD2VblQIwgPNXtj5vKa5GfT/23CyJr6p9dGFIJCxzU1Wothy/Ma
pQrS50JAY1xzeZt9O1Rw0Fjuc4sgfexmeP1gQdwqqufjGN1mkekX+DXRI6wnXZMQQXzFtrpwR7UC
Hkbsi3NXQh413N7eMaUNAKqA8FcGHwabNCHv6T4mo/UtxBPCsw1Nk7WfkEtXTsVh93l8ZYr+/SCF
lCW7Pfnib4AkHWEsY1Sr8TtmUaw9r9QoJOHTCEy5VIUmUlJLb8rBXg5USbyX7gY5finmcWC/0Qku
nOtOZrApWW7WgiRsc9xiE0Zhs0oB9/48sYDfGomVm/eMft40N0byCg7Qlqsz9ZeghLEVDvdzyb3D
i5ggQ2PubXFBWCGMGA6/PF8OIyJbv2Gqhy/qwdHcydgTAmk+XQrsD1Vlc8Z/lmeaQMe9AQNDf2do
G/kg1GiQda15RkSPYq2OGh6k4wmRxIOqWBaXWJeUotNm9KurVwHa5anQ/2M2mFvtM+6XomYBVBX/
X9/yd2S9wWTHWCaq/3o78/ZdsPUy07kr1X/icrFAVqg1mRpcQF8ui9SX9aEG0eh5uBTXQtVlzh1r
eeH8ByuxEQNaSRjilA2A6or7TWSDvGFVnTgainIMW+sCylm3NAietK0KI3pfzEAxPM4EF7r4PFy5
8JfeoasrY8QKjsWwUfiLIO8maY76iwisEd8sqK3NcCrXwAkEqaj1iNvngDxovJvKp8bD3SWUaApt
6dclpJF9gsN4OsUSRMFO6zTes3YnU7jqUNrsYMwCddHlI5+TF1RdZhIAdvRoOGNSo/CuSvBuY5iY
MbEvcOLj04vPvv8upowzlAYvSRRRDVciSHVZ7K7ynvDT0PSXnzF1H1i+dOPqM9fyPtDU4tRChG8V
/fyjHoI7ld8hWtiBBhaYyeoNcEOkJP4QaexCfzqwW3+AmPma42QmoQ61Vwo5970/p71SpnyXKaWs
io85WqtNV9uzI2nLPftRtqa0ehIug0NMr6UKv65GJ+UIfXg38c/vGm2eRNXxW9wkqdCEYFWHEd4H
0ZzaqBHWSxDrbZt6Hs9UqyZaSg8sHA28gea/Ja6lhOv3QSslhATTy0dEG8Kt+Ar+rF9rE5VW/uvE
0pvyXWG381sO7pNKGxASw25TWy22rR9qutP2uHkM6a1rxCq0mwvBb0P22GA7HihzGYNoxMTQX3CR
U898Xzy+ZfyrCwYKJ1nBi1ak44M9Iw36I7rYgLXJ4B0v54954bQrNEg/XQgVlwUQVXI+uLxQeFHa
R65aR5YIJAYX8Tc6fVX1+08SlFhnHVfk79GVqpKchC5TAvVNw9/+dGhWiiUxkfcYCHxxPktFN0Zw
62eyBuBRFeth1TW59cegLmsn4KPvOXjdilR5+dTiZPqNm6SvjVDiTFfhY9xLCc7rO9tAyZAPK2r6
PvFT+qr/M9AkEwVTffgSzVXhQssIqALFXm2wX6jY/B+Czh0dB7Mg1n3p6i8UHMzX27FKkQQvM8pJ
pGRNbM2+kULx/1tvIYQBknmVKFmr+/nDWOT90wIRkvsci9lfOGrTkmkhYUbqfBMUyehCVVb+RyaZ
or21fKemSBOo1KlZ5buOCQP03WbkRKlx8kxT6UzEf4dwvC72lRqPUn8mmcp39nURzikg3brumxiZ
iPZOUbSzUJifDqctckvxaQ6k9Pj3f8JrQH6KBwRuZAko6ykmj00A4AaQAFyKiiIDF2r/XOAyADNm
/HTTUNOimJT97ICGcHkBnbU6A6VXhpKoXEBCAKNiUff8l9kMRjqOvmmgz5Lspt5z7MlHinIj32tJ
1U/4MZ4ir43mow0p+E5KBvl5p7nKInhe3EjdPAuhwAARaWcCoFdxgSx9A0tIm9GlFCIjHIIWgyRq
3T0bsQbWzfeDXRkvQoOSkVBqopASc11f/rqqNE7akQ0eTmzTb8T093o1hbOpwVsasHjI7FPicjo/
7iJFgwILMLl7dveFP1KfG2b2ur/PXwEV9Si/I1jHzoONUrGpGknEMjaEu8PZcVtmaMTQ1u9GEzLW
c12vpWELw1nGsIu0pxm3wKBqhb/Tcuh1joYAiiOlGLdg8EplHPhKxRacmftGIJdnu+j4M5GLiRW9
bfA6Ub+mnYTKuIBhzYpznnKPsFuzGuvfmuLNMP7Hr4PJw2D2TjXk7NiU/2SgbCJPYO1jJe3CzUHR
rnipGnQ4yjQnraJxSF4OsBw16cXO+FqsL+AUkVacCoavmAXB4tw4cGlsEWNMoYohndhYjZn7zf9x
1XQ4nYThkdBWo49/VdGvOe5Q+vVmahJpFDStAMNORHkd5bZ4obEm5n8eqNMMZUgC4kHfbqtvVHCK
uchSdMqk3ZCnbqittpYwPsUgZWzM+MGqPQIWjiJ6sAlnX3zN3heRuEf+UgvzCsQWIMfDVawOCxEM
JCzrOgjGcKcnpf66iOWGFPigR9Ly5xRazYmvzg16FaYL/LYnocBvqCuu0feiF7U1s04XNHP6k0qx
0A6iR7mRL2TAzMWcMURMCC5SBae5IOmP9OuGF8XKNsxaMawU0/j28xlzs5LR+3Gstej5rpIFDkbT
158zJFPCThtt6MJZi/EjZ5j0aDkGjBBXOYWvohz8P1HE/MXya3cAzp0WpaokwLNWcqimPbrPhfhT
Vp9hMSUuq0db0bbcXez7Yghpo/L1hrMAlcoI5FZvdEQADNzkLpJo01u5XN9IAGTkWmlUJHTX1JhS
fCEeBw+RUC9HXMFPHWXAiIITvE5uj1PjVi2FKIHQoVqlvqsUikzi6zXDzIaf8An8mgSKO83z9A8T
KPYXVfC+nGef0a0sflWASZFD3JgcE57wylIQc8LCSW0bkBxCYFOlRVVlZHLKcOyq7uOeciAmwRAx
hnKDyyIJRol62ZlYhmO9pkngAvy82ur7zM8XKP5r+AzskXrXIBtE8NHhQx+33P9QJSLBfES37mlq
5kuAWoACK53txQS+d8gHScjA0oosBcwsSaZR9s8vYbnPwXB2JQVsUS7BCd3P4S4HkcV1jOVT/e1H
U89N7f2LfbB6+7Vu41mogQpmqJSOemtymtdeZ5A9eYwEGUjqiAncBSjmgeYQoO7tqsyIknHug4yD
Xednhn3/+KSTWHWhqo7h4cHpYv5ZAZVJ47KiAEmM/FCJJn6xpbLhPRkqUjMqpzz7S0LFItFNY6Cg
5TJ19um/9uebxpNpnF3wB7kj2dLyjKKZvhzQVH584v0WknS+i1YEzzqZLdEr6bXyCVhQXWIVEC/a
1jO3RHgVUijvrXqR96LLtTF11Uoa83FKNMUH9eC0vtRwvARmiNQJxV+BXB2pGg2eV4H1w70BfsPp
L056TbNjGIi+tELhvrY/zxNVvi/0Sk2fcN7VMuKvH5zEtZCNS11U2xgMQaAPfzALrh+WREvFuo2/
EYp1i+FvlsFPtoFaactzJ0fNzQbsXJecge1U3MaujbfT6HDNpenxmfn9hbVRq7+zYPRcs6t3T9sI
bFRLoGdTNGW0fxdrPHBrZiSH5HrmKr74JaasUKeowY68kRFx/tKbKhhaEZED1LhMhF4l0UNx1UOW
F2q5jXHo2zhBgb8gj2a3Bz/oHVd8Z+NPs4x4L0jOZSLq0ouo5dDloL7+DgrHcwFuFnG3Nr17qr7K
6eE2ins4/eCaxIOQC8lxkfN0jsXKMt+kg/OJ7XyANjROLqTgMdZZZITTkm7tGZ7YSUL+NiIm57q+
1SMYuk2UrIduxQ04o6tCcPoEoihE86BFJ2GnvgMF7qt3dk947hMUIbvDNPd1wUYSpr+uFQv8q3Fp
aeB9lDzL1qc9UXqrMMU+ix2WzHgZ5q5Dd49p95qgpZ7wd0IxNa3hEWR6Gzq11swk91AqmRwQbaOS
3bKWdIFXJyxdkTdtJ6WZF2sICobjKY9xpyr7Sx/wqgdEEY0naqP1k7k3QbsV5AhjyIr0xxrNZk8Y
XMfOT+Dy5wrkUQArhSBr+9hB2+RYFdefzurqEEoU+QD9nqmoJ1ZnlcFfpOpExKMBwqfidxpQXhZT
PaDdHxte7gftRQiDKExeouzS3oP3OGgxk5d3Z3JbnkYx9aYz3mpHJP6IF6Tm/ik4+XFzfmJ/+OOq
OngepWKKEii1mj3fj8ZJfqhv0cOtyp/vQgPWJ3Pk1/UXI0JKVtGKWMQYfcyqRW/fBOm3+BrrBbHQ
sk8zRK0ustHhgnJ3NUP7/KFmUtKlB2aIwXSMCeJJmrNzGqLWnQ7xiDg6/L0sw5aj8HggH6BxDiRg
lMFi5yOKVB6zQx+5TY7XohrbFgv0StVa5yzMbj1YmrQWGruYqyzcDqyKfqkrvFjkxoWysmfIfj9q
Qo+3yKQD5D3i9a/3v+rvD/EWpalmHAtotdWBeMAR2WurDPXvNHhRetPSi1ZM44zbShNcwTRYm6t8
43Gfi1ooQimX/Ma2JR8VIBnGdIN88cnESnwBwP3bvptmFUD9ZzG6sQsdirTTADb1VAHMErEgdmmT
FFrHzJs/YCEqvUJbnZSyh2ULtwa7OhlIXWqVmcPYPIqC7TAX/hHtrlqeWWf24WwswYmyovSmQwGC
SGID+bIDwkbT/GsEQu5Lq+q0Q7nub52dMApzZg4s5w47y+o2Ier6tUkX5t5TloRIGTSn9woGJT4f
wL0bVhwtiQ7sDYqH+gD6uzj85AmvtFo6fGSV4/G4S81EnAtFzaQIaZN0vvQnoQteoU5YMBeqP6oa
RCV/PGn+LsaNzmdGPPZX0P2cntWxL6CNuZ5vk8TnQpXNIBvaIRKDB7NBQJh7O53+QL2tI5C2bIN1
Xhi9voIeNbiYKdSEZ5PMcmM8gtCNG/husJuNzFTZ3qkCWpBExR9IozLK/YLjaTP/e/U+A2MEatTU
TVY56A/umZNDzY08kFFMCTcGgmbMU7UB+LnhPYLbBwk10TLfOIdCPwc6p/ogd92k95x1xMat1iCc
ZzUnghP/xhOXNKhx4XuEsn7gs8x+DBE16de1oh+V0qLDOC400IhCl33kiYqGiNjC/oRVMlyaQq08
kU4y5DJnX+HkJrwhtGSZcHIZkbTxaLITqmeuUjrfIMYrBRCxM66eiDAFlUiAG4AvXD4NP8CqGwU3
+pfp2CIzpVqtjzUjj1wDemxRKkPgMamQFziE+oTKlj1MSb1TDGax+ThriWJxpY5R1nadG7wr/7hZ
WxMDYOOysCZGopmwByXAVUnnB2W8shyPc+HN7MwQwKMg6W1U+9KO9J8Xb7RS7vD2jPSvQ/iKV6eY
yYcmWEY6bd0rWeFWQDmQ8hBvVZAQdw/naW87ZE14Jxj8FYPSC/t1HSBqRFzA/ZNlNF0Jn+hRV8Z9
EpAPuE0M/aV+T3yGba65adnA9caMk5qGaI6ycPmcR8bpgSQr79yyi18myNHrf0S3mZfBZCqfJYVX
rOfbqD1iBB0QR564Hyst0yrbl91XnNFL3+QYbgyTouqEgJLJ/n0GE8b5UutxhSYfgBofDwb/TtwA
odylhFSNxmuqPOJOqLiolqb4a71CsbVvrh72irDzknG2nmBwXt6MItgiFKcYsbohSV8ufn96IRBQ
HjYdctsibACaVWNAov2fDdHHfb7RJuPDE8ZIMES9lNUQpMBfFYejQoKrSB5M+rDfjmmieC4TBhrx
fyEFHJoexnPF52V8Pccdh7uzIJgYeaufvjJ3UzilK7Bvbv7MbprCTkhQijrsTXQOCVzfuN6ce0UP
2v4aILRt3OAjXVDy/Y1C5Iw1F1v2TjVFeyAzYwbVvd9gD7T6jq1a1OCRF9/UYIGpVrGl+imeRTBK
DvHT7ncZRk4taphWGDhzkKwb/2mAbpHFz+hU9I9Nm0s0C+1b1jq5rHT6HE6EdLHLMXYtpJIS5gl+
e+Cba4D5vsDy7Q0oiHfpLDDoBsSgN51hoHEgxcWhAh0+jYOKkOJxXaFtG/UCoShzQA/EgiOh4C1N
YdwNi9GkWAu25IJe6EVYQtt2geC6uobkvrF97kzQzJ4I91Psir7DA7rz4fBrV6de+wYO00qqun2v
gN0FHjLgheEv0MwfQHG3Q3oQiRb/FR7BEIyTJ5o0EHEadPul81QEjbM0c4K/j81nZdbd8wXDsan/
g46kN19wnn4XEnI+wEv2Cv4TQH8fukIK9KQxsR8otUxzcxf/xPzy13zxm8tvcuR6SLS9CDFBt7+D
ZOxAhwmNQADIQnNQrxHUTkOhjldzcIUsbs2u0XZJ0GfurSFuX3a7vqmkEkQsmUEko2zit/UFLg6z
iM5/UpExVHiQWX+sx7Ee5ksOUb8gblc0bVPHLbfSPKfaehK5Eo2mYQGB97wEfDMo0EC6b+VosV9m
/DSsGakxDFsdu2gOHY2Zf4E1DfTK1awCY9uMqyJAepOWZzAWnELN/n8SfYH7PzyoOOPyIMhUhkkA
3rnvc1c2lJZkjrQDYgpy9/3/XiLdQNBtq85b3c4X6K80JBAfVh0oZNkr9cIZUD82Z00s6Oy3Qs6D
gRArXFEuMuFV39kGyhxI2xZOyo0Nv4HSm7psB64CIUCGR3NSG1maNe6wRcZRPgOlzY/D+A0HP0ur
xSigAfxhQw/FAAMniQijP4ckajnzwpy6f84yl1+IGEj4Rct8x6yR0VoXei6MwMR4xAuVI4iF4VBZ
mTH399XhWiqD9HTXZ0EkZ8S9MNPIU80nIJq5d+llSK8QowuktpIuQ8LnDDX8kr6ksfT8PGN4R+Be
CjH4JcQWnVn6+Q82gUWjyqSTWbvPV8+eR7eJE26dDGIaWcsnT6sxf0vUBgtgTI2KaJqIi8u3FXvz
V3YON7IfUWMKbJThclpklCdfdOZjNK4s7pjDc3Zkbfp4BBaTYG0ac4UWprNqrOLb7KLNxYm421jY
cCMd0Czcc7RDLjMRSnpSKFmIQzc+YWr6g2q5/JbCK2troC9CGsfi0M2BaNnyxJTdnNXy8DB+UT3W
ecO1br6xSN2gt2Hzayt7chZprzO81zxG1EQcplKyCAOhbDR0uig/Idg4b079yVIs3GtOwn2qAtv8
b0vZa/GadmWOui9fl7KY62fvt8kW6sTO1s6pQi2IVTau7ARSO0ixQ8xe8F0XobQ0WnysMcDhMzU8
U169nOUDiwZMxTrJkc4oNi+rxfu3LV122M3KjLB9eAuVQ/KqGAIrfbRevE9UhtLQVSACSAcvMHrv
6CMceG7PgZwuC/3ykb41uXSLKScS34zULtmJyXP4ZWVolaomsU7fAPvbQnxE2s5ZRWPr8K/1MwGl
fC2xG/PHkxBn2X7Vhpg+LoWTz1Q95Ieel/wGhQFVdukEpX/ipHuQV7uYL4WB+7DSph1FPwQ95j3A
E+gbIxJJmUIuX9Z5Xd7OqliFfZyGG0S+fbutntM557M6IqzUaRW4WPF1Ap/7t1nObq6mTJU1OuWA
xfFsJnIITVM+QV4/yQ+FSKjZROfe62FaAcyfJyi+ieKiafiR2EHjFWf9u5awb3u4TZhd1Xg6Mwog
Iqu49TDahQhZaI2XChZmDCH0p+OQkeiPa6x+lgsZ5g+FXQpgajEMk1oE2oxX02kMJOpHgZbPL/9R
Ap0cjM3G9DwYBQO+ovrpW7nS2dTYTfJZ8zCOq2QsUdxKIpuyKpSVhU7cDB21dcyRHToplyF+owU6
VSN5C8ypglhmxKd66GJzQ9j5IBLjZONEVGQ1PUt+U2CCw4ASsMdv5Gl3Mt26+cR1Q6wHSHCvRBMN
vikENGPiJrjIkNvObhztoeaPDEmY+yfdqfWjuskzCfMDlvIZizCD4TNGMmoMdTrXYmELrQAnOb1U
j8Ign7PJBdme3dR1wjb4TBoVv4E9RkSNHttoaBb4G4OklRs4wGX3x59Yx4jiU+iE2mJicXlUCYJJ
5KCNJNJcFTLWI03jdGx5Uie5mInhBugRsZwl4iGA+X/jkGZ0hHm5d3i6nNkyqU3GSnjVfX8pvMBN
bgMh56lIKrZhBvIdL/vQ2BYgxw1J4OXqrcMpq6S41/Uzav0x+oYH1umqg63OLrhI3qCdrR3hIg6D
LIsqt8aOzcoajG5aqMxNK1MHrI9FE/nrFGX4TEPlEPkV7vFdTsyFyvd7Vwafq1Eq19l3/UknGAwT
tPOYjFUwyDDNv4hQ9+ak1nmw8ZNymSak6HDTJ71fQIyB/eWhQkX2ickwrGXxjSqDMu7c6f1D+LxA
V+vGJ5jvgIj2fJAJzKDPZjMZsIN+ITP+RlEH2yY1CuGQG6dScQ0OgwGtLnJd9sR/DV23YABM7Cwg
JttnfQ45fiK5e3dh73wxSF7Dex0427fOJoWyysHAZMKo98rdRPx9wwLHb6cxfgDLoQ7hEf/WJD1o
0kmEXlf41/nRAyx+EeoYreyWki3oko9KkkUf1cF34T4G/vUIzr0olFPrrPwzveQUQWGebhdXFts1
/mQs4B6N17O35c8DqQh8Qsj30nve4h7avVN+jvj2jtMFw1+vVoG9IQAvCnMz8K0NMSh6QQNLZnpO
I2iWVdfn4B6fA1MSB7dN919ljp2uKLI5e7Vj1/h9Lai5UvRh5HLPmxeKVg7oDItR5Tw9Pi6DXcxY
lNCEREPTp2OIUbMYL/Jk/klWK/TB4k65dm/gu6akoAwsz98BNlIteY5nLzk574/e25H/hbqoY/pZ
rNZizLCWV9UMQkpbleOS3yc9ZOPkNBVZ9HYcqwpWHhQHWL1hIya6eZ+0ABMnZ4dK64byBzDKRVcS
BctKiaaKfQE9oNAkgKXPXkIZTE0YcBApNOZAf3QbpEjBocSNtqHc2FJbCXf3Jp1Q35dHXd0TuSjS
1qv5NO1ouJUvekY744IooVVx577IyuTdF4jkbmcBsX2o736h0uccuwmWVBWxSLE7bPWZd0J9s2Sh
BFDhU1+BvMBGX+UE2d3qifFi1uY/0ISx4wOdrOXUQcnT+xXkIqueswVWu3rvTt0seUXJikcLxBUy
YZOPyhGgf5CFZ3TJgHt/3EXZy6YE9dOMDgUH4EZrfzApHhqq4HQUPsRtmDJ+gKhLlEAvVktLf8iO
gVCDdEXKuzCtRhpdVCn6DUBjP0FYQwtr4Eq5v9XqI5yVyB5m7HMAHrtu7UyZY7gWUPDBKE1Jn+6F
izasi5ycUMAY+8ublqCkq91+Uw+P4C0KbUj4bOV+yUI8+dw73Ku4eahEb58V2m7kyc+a2xLfB/2o
E5S44clS6NYGGIDYhJQKb4Mzc/GN+f+o1zxn3uouX2yVWQ/iko6TvGA5oGWH+wVlvuNdtMT5BodZ
3Ei2T+RtHJlDwWg9s6GotcoyPHu7poUK8lVp5L7NrMqDFvfO5eRTiWnZ/6TynfQcTkidsp6bZXdB
sdo4jSEXcSSjDQ2K1NLtW2r/FZ4TK+hWRGyMoNpGdWnnaPFNJTXHXz/qcUSMr25xv4UoAwNK5M9g
NiJzr85kajoj7nfmob53l2D0q3FEq6PKt3gU8zKyriKpHjEjxdAtSPEyJnc5JWuTwqtTFIhzrYEr
qVzFPaNnJZzitfLkljJl16bBszJAR+T5NVXp0Duhn59aTtLfQxANCk8XDwnnnE6jRKJwcE0QGgtR
hIw6wedqOcaUFLpeSfFNKSL0hY4WpC+EcpnHjjaHFbjOMuvvXm2X/NQ40vbvDNqDx6ALLQAhY3vR
+BoF9LhwdNITJAJIVwcIKmnXMusK5yQxzrHJG6hDOSJyzdR4IA8dFpN/jRFbHNKq5Lo8gdrqkal8
ZssWI3Kxmt9fv/CLTPEU6DRQWzhjQddwvBZPEP942AHKaq67KAnVvO9U9M+MX+BByxYN3V63MNBw
37zEf12fKbTpX9OyTRZh8SIl0WjfWcv7DsRoRu6p/t5V0QgfOZNagFED+m24+xubjmouFt5+ZQFv
WpxKj2LiRIYTZ0IOMNcEUoOZxpCf3BQhL4/LGeMjgx7LC1O7cYQF1I1ZIsZQSEenFaWCPc+12ipN
ohe8S9J0+5oLRXoocD3weFma50yNcYsEAVcF3xMnQfVE0E/NTv57QskK8ky7B/jQxYHFphe9KWFt
oF04HzDCjLMVFj2d9nA5r2YmlRtsMYQZsOE4WSqmw/VFoxqEWyQfyYRSKbGX2ARA5YtUOA9H3h2g
JCJBD0goU66gBm7gYsG+fKZ1d0MDDQeK0LluS/FtvSlkjadK62ZvMJeFnX37CCxZ9ENuBcruCuHn
ijNbnt69c/dgmas8xV04nPa/L9p9Hk3E2vzBrgNWah5+RpiKwe+fx4mNt170knbQjDu6+4n2oZXn
54ZTct8ZHmjJSFKdpHHzUVE6V8Ao+xOv0wuwVZYcxLmhlKm9t4CjH1Ku4Y3YWqGc6fuZtM6oWJ7g
GH96wBmDMME0YjSQcJdxDI/8r1c2qRaU62pQMILGn5o7sXd1lJ4kDaF+5PA9GctD8h9hfybt0PRu
P/2MQk68bGvD/ftSyF5/eKFUcQireeerStBzZlE+WrEaLwLcmST1Nm4Q+Nd2t9/6FIw2VmrI8RZs
pp93Q5/pDoujsjv5BzYH+yKN41asMW5V6CInMwLO0OUxJInV//W9C62P3lcjOqThbtVlP+GtPfPM
uchUilAuj0mM7kht6LJoIlhxtv3MDo/tcCNbMPrlCochUwvCbx77Ut9Wr0/p1Xj78wsGtpRkMG0d
RH/ScgwnLqtCH8Pm4QkXw0Ft8TJOhlv88cNeiv8lT/t4ba1H7zwUWC8UmIUKFwIUme1gnyYirRlJ
dWPw6XxZjT3K4sItXY8hhX7M9Hf85wgXRrnjLW9VpgndlQWankFV0Kr9hJ5t0ZjFfBhx44gPqN4j
kM1Kn+Cx/HqlBQwfnje+RxCHngMb+cJcfJwCdGJcaHVVgAnTrV7t5MDRnPzcggkbC7UOfQK+pqLx
1opwc5knDmGgcuJLLZ40GWykFBjk6DCDMd85gQdf+PWMcLzlkXvQ+2DwfQRnXFKtCWkv0c2MbvMJ
aRT2z+0AEyxGHmANueIsYa7gpI/CPdkilIX0rvut+Mvl5yedPtqWyGzLNT9lmuiZF7X5fC5BlSwl
tI40fzQJz5ZJTzdx82vEVDB2T2Q7PFCg1MPyAZIRtFgRBtAR3DlrtuzMQO9kjsSAz+pQMNP1dzh9
XMqqi1bPBly5I+tZuor363rGToFftnjdIdqo3D5ELTP+LEM04i5hrtEHoqLSWY3lazuUpM1yegrZ
Q+q3x8OZnuP8nbtzH74+KrkAiLldpdu10H/1AoSjeFjHvyCvmFHr1u93jLZb3vN9E0r6oBs6uGAC
Mg2RD6iy7dzQQjqKmsSrySsa3H4zz2cwJE9r+4Ymgm6gkppBnIScNj4+wrlRHmhsGLwU4fIqWm77
Suqm0i/UIEzC4Cv7gjNgDPPUf/BrG6m11/EYuOoEGpVam4RP5DfBhNS0CLytjahgk9XVm50dv/Fm
Brbgt/r4rNRVxeT1wlV9buS/9FxvfTZJqXTSgQF/JRlQYtY1p3sFG3Z4C8gpxnulNmXSjMThYoq0
z5xGM321yihhEXzSlN28Z745Ug3uFF+OvhcVqHNMmSrhwSxV8KCVZ5E5QUaVz/2tme2X2SAHvDpO
EmhhZ1FOCjaXOj8iW6lsp7JyFflgE4AcxHNg+TfvrwDW0aQgIjd7XThIdO8d2pNWWJi82GmssRPd
MoO2O34Gx/aIAUnmQ+SL7dkghIlw5V4HwU3H8L0AHsjff7T2U1RJvJ2iXA8LvBC37cIGWeHYgQti
FK4s23BmJP6qHus+VTxHi0Cg2IBlv4TdAL1CRIUzF1SuLrhx/TqQvrniy0Ep0ffM0pEBygry7POd
CZpBdMLlxaiZ+Fs+GxJ547d985A1VSaACILEOdRKiXDbNy/OgwciHNibDwKdNkG2YqPFZxiA0niH
BPVnfuIi/Ciw167goVIcAkcZiJYzIJmRTzw1NKIL1bkdVoViG57XHbM2aYV2H7XWRqkUdMpBsS1Q
V4U2EXEEpE9ZQq1sGmZCTb2i36UQBVp88SE8NlrU0CISS6o2kB6v2Ru2pbGKyHe6mOarv6AAZGbm
3MXR9UiF3I7KwcWMIk4SGvVFpBRBzMNbIFcevK1a+YM9kh7lZtiq451hr+yPXSVURyCFEx7/dlBE
WSevDTlTkb0Po26O+XzGYWjzJi7hOBAXu8M7vMY7pfEjOhBcglCDLNC/cHV++Lt9AtD2XUICLDaE
cHNnYeMZ3ViU3ADcug4+htxA2xm8oQJgYpg3qxcBu4c06v+aK5/WxLiCQy77/ExGs3NEx9E25FK/
hLnYmDrGggvxwoox3RsUjkdlQLaKBFKyHZgQjBP+mwwNQ78h7+lvBkmtapmFPZeNGqx5ckZEOJD3
GWQrXPZ6SmZL2HfQvCL4uK/h2J7+4JdTX33UemOVAkcw6oyfVT339ThQGiBLV/Rg7iOTIFrbJ1AB
UvY98wM3cAf5tjijfeUc543ctBrBuCYr6nlwdN5D5xhPtBra3doeLcXBn/GHyrF9MbrPmoYyBULO
OIzeopMz9KsjXguJidwV82GhKNqE7dtIzlcT1KV2X+xbJD3M7ZYzPHZrUH8rMIaPKGxPcAAKf3pR
HCK/ap96UqmTlKPIZXUnZGoGgGyuE+oFcXUKWrzVt7HQmQ2aTKSXB4nXol9CoVaGczvEKL+OmjB8
0cPsnOFfghMj9vOOuTSFPOWCKMzjl5GnlAsfEmOzxDrCbzklIyQuL52huKEpPzedrWXjD1Ku245v
+Yy/qT8XbeoQZzJckddb4cFsaQnMg3YK9PWtRxtuqDqpDAZ2qx7eNeK9ddRaFmf8VoeektyLmGm/
r5i7ZK9mVzbr8CqJEFxOUysWXMxPaNzAB732Hz37XJ4WVw3X80sSFaq1TaxOvUFeELHfG+QVRZg0
xuhqBIDEXuvVDSyvMBxXASZ9GBLkPuJAtD5hH8YjrcoVmDyL9map6hlVKLs1k3B6+d5Jig6CmTe8
+KSEtgUejXaV/rfX6ZRUse+1s9FVgaPCzDgekHh0p2ob/GlGZqPIGVL+33q8E15o0nfwRh52eoKW
PNJBs1DktLZ4mnJr6b9GMeOJNRyGqoZZCsgu1mCZI4BnVm36e5DddZn2SsyRbNN/1l+MXYM1TYLi
1KzOXRsUtJSJ7jV8ewLsacZfVRFpcHrpNZzdFG47Sf3Tot8mleLzhfiUvSOMaIy7e+ROP2NdTo0O
fpXKmUs0AtnNQDvpz9KnZVZWidnhWJfv9qwP2s/O+YaxhcoZDqpPsnXQ46DfV62ufNClL6yP+oRs
KUt/TbJzXdA8So/RdUS7/Gz+mPQGw5kojuQXrnitL/vzVGhoBs2tIONfEs4hMbPUIqNX8mH3fVGU
T8ft+17t30/Fmaou5MtwtzaVRZOURLjAs4uKbsllyaCGt+yBECs+/Lew+QrtbH+MRzfnhA71RDvM
tNA4jZIqZDKQIlv4NfulxKzz1cCpjEUa/PDOwL3fDUa/++2eE4ASBRMuRv9zE+KWqxeb+louQx+T
o1BgODqvFMxGqFUxMmD12afGCBI6zS4IKuz8+KvuGZ+hB5QE/IL6by/ixhyZzXgk2YdrSq5BjVdH
Wlith643QRFKuvYn2Vk1IAicen0Yt3gcCGnNxVsVrRnxzKH0hLd8cIMdbTRprq1Ip4ufzcHDkmTs
NwAdjqsfgO6g4gYxnL7uzXWVu16QB+jqHT+qYdCv4pGFy44UO/3p4NE8bax9mwNX8gJ5DMhmRGcI
5fPHarrqkuQqCkNrbxl4e/3hfxR/CjUAWTrC2vRAWknFUxuA4wselEK9xCvzpCZIEWR6WImPrcKW
m7iyYt0x8spC8MyLpVsdrcxzJmDTTPgItQ4/jHM9D3TfnpNV0brQ2NJaAiwbooT2C4y9XnZCPpZN
QJKRF/OFj4Ib2BsdwrEDkqpwXWlyOYNvySLzBw/+IDL678NQ2FJz+nXncqED1oHD8enECCpj//3N
YrTgsJ7Iz2Tk0elDVN3xk2if2WJjmkGZdnxzgLOcJYG40BI2mO1JioiKtp4FRqJl/CgSNSQY5akK
AcSkHu/CU28Sz0Xk3heQ6RjzhIcjZNEREluYgbPnWHPBWu5bjZYHBWAoVaXh8Ky/GGCietRBYjgQ
L2/u/op2HS0RT0lGL4NSftc7YdLpR1I+mcQJA7zJWmqz+XJx7q0Lk8KxV0nKceAIZ83FKBoZm7Xk
xvRwuVbc0gtqkhEEjqQ3uU/O9LjD6zWZKolywfx3/noh3S64Of180XfOt6L+rB6iWDx0ysRnU/t1
4/4vsddPLzxawozw+WHkGh4q1JA5rCJopqyhpqQMJFq6EnDPs9A5MfMs88MWus6uEJSLXJ0rwX8U
D3X9gk7cVTkmh7e6hO6fl9ty+fgCoAASjKDmAkphhizRWUlE12ZUP2bBbnbSy5gUoiqmt50uGkrW
/dFUH0CevwlLH/rcmxqmv05CCVBEgQdYcAq6AOae0IuG9zRHnM4HWdRGhAFGIqm64NmnxtebF8xI
/QMT3FnEsEO+cgroqhzzrHo2hhARbVj5RwAWkSlXzFd/mCaafAxYTEdDB/6UmBPPkY0B28dWQY6q
RUyHlYoeHdEh9BPRsS+VG76+ieeAdkBGJXvj4XCyqZ9V20bii6tkEuI/fsRnMOS2OMAb1xnZGgw6
Um26x6DFypx9H0PzxgOrG+uAskdaX8cxJCnZok0SPkdI7f3xNq/MCUihUUxvIY5W0Z/QXT2w1/MH
ZEUsBu4BvTUM/vqOra7dOaT0oKryVJhQ6OfJYusJVmndRfr4s1AXE0DE6tjA8YeuRLny3hw5w28+
hJJ4A16EuaHaD5MgAOFDRJikqfRZTEmjpSadx/CPSquCEZAxZhwXnpZsIs1i/6tNSyRF+AfGuB70
izF4/oxtJidxt6GTNMJ0LQa2bO4KxG8gUYm0uz0UeoTehl5niuK9gVeX+KsXWIe7WB+Gd53pIDJY
5L04adM+hUrc9K1MbENYKkuUm6J+x7OML5ZHM1ON26fU8hhQSm1CzYgMzSsY+FSv2/xQUUxLBaeB
R/52AJkS8Umnx0/tbmkVZIceAwG3Z+yZXPfAXsgcyYTrneyhIY5rXZ1syBy/XpRSvn3s9/q79r+v
OldU6dCcZdVh+M6XxOFIgWNENUs7QVUZPl7xMXrIoY/Z9QqwpsdbzwI43wAXOJZahTC49zflc/rD
XNcI2GjH58/H4aIda7dUZX6OqpkSYD03ajJBJPnOgXIVQzEOWHcZs4uvY/rGH2ZyF8cHBQ12COma
igVVDUzJvWgYO2IIdnqupJxvgZbLYm/X6w/4rpMRCkO8BWrNwfPZBWv2LI4ByLwas6wemeVs/v93
gaW7NfjNmutpMiNZZisubZXIkJDZkqGVlq1SaOw85mZdSp+csFOmmQcaRA2dlqWDKns4LxOUEMUq
ph9vIZtJmGmiBw24TSrdO912QR+yyQPTS69YmCTwBVDv6Bkag3uBBnNuLgCdzz0eXN/5aVtMMwKd
WjE7EJNYl+ePraGsKi6PaiuRa3Osi///1puQO7Jx26QNR7LoKb1U5ObTZw3zfeha4/3GA9hZwnuA
bZAKsJLnX50Zj7fKQwhr8N6LVOw32KIVMo7RGvGERaFD+8o1nGixTCVwVdmp5RKR6d7ya+RRCD98
yc2H1O8Q5E0GT86qRoxpNNlP1jvFlQTS2XOLhdNK/8mRpC0fLU70MLWrs487KFxTNByRl5nzoh0K
RbFHix0b65Ut2U+6LDO1+bl1N5QlyuWylqfkCFWFGn84BVhwNewR3pqZUrkCZ8ISgWoEfJ0KX70Y
JwtQSYRnDnQKO1Om5AnunBY3nc7p+gxJFRzmgt9l9QTCLj+/hNU/UD+IW/5DI0ORcgpjTFkjt9H7
JkH/zo3Ij4eGU17DkvH28sgKC6skyC7iQXejxsULAnSs0PWyJjtHHpe/s0Gv4B2Wc8Q23hbJNvkF
FDmg0Yvy6HVu3FuO+927Yi29n0wQdw/Z2c+6YRhy3kKCA31CiF/W6rf5RWwOkO8r9aEL7QRqeIkO
ZaQHMgrQSoGjL2zf5lopqZ1yV8LehPZNaO6dFsTm/FPKBMfvkLULtrBUi2MIhD/TPBrl/TBjynrJ
g8+DWaYY9PvgyswPQVr4O9Xbrir256+foloptXoaqktgBKQxbi9d5Ot1uqcQC4jUnD2Xht+1DljV
G7uvJyGfZdaPJVElOkO3UG7O6Qn6C32/anojY2a54W1cOppqeI/h3t1Oah43EGQxr0qxdEutRaIU
57uzXbotFYdBDiUOpI4qKXjNf/GBzPZz3HQ+l2HnXPTGM1TQQwr3QDMOEifQ4HfYLnAHn3xmQbw6
eq89KhI6XK9FMTLnzDV1fVgw1wHni7vSQ2+vqeEawE2YmaUUjumq+OzObO1A8DKO5BJ1aSav1FDy
Iu1BkBPeAHTpU5jm+k40XOqygDWbI/2Vfnij/BNGtmBzl522bxGJp2cv+sWZvW76w1R1twzHcY9r
tgjYwpOJ3VEwOrlwZb5glRTEO2VYv9wc8Png6UQua6FFVqVguV9TOvVIXk0YLIBlqxmYBT2c7v4L
IJx8lSoWx0ombtt5IjiaHL195gFBD2l2DGeF1qMR+Vyg60BhH52f8jfh48U2chpgGcaRin6n4ImL
Qsx/ESWojH1D2OOQJPkwXk9F22gQarP1zgl8AkM8IiPboiGwACRhlbK1x+wM7YPUP6MaIUJ5lham
mlrtCb8vA1vzhtQMAyWxDYkc8UdZrfAqwDftbTRNQo60h0v1szo5o76c5pjJYyhIOfqc0kyogXAC
DGIs568fJU1UnRx5M7R5YYYGZPtSFOmY2QaihxZ9NHy5FjKntZZP0y305uaeZxFcsUJGoqVpPf8H
LCUm672lFtuaJV6bFD3+MiZPBWq/bYxOvDbmbvmNMZdvOlb+wmRfUjFCxXyx5GZd/3Q61YHbMLal
6tTBgfGchezGlMrobWiLRw5WkzbZ7VDfVisz9u8ENz0/SoHVsQyTAcAdz7LIMeHl/xfTrbZifhx4
jpz82TbGNuflrsE8JpBP62THRM1HJDU2/Y+D5F3nrGpbHnkSoM2A6gcm7SU6UbYbLpWRpbxElDd9
xKFWkDnmrbJnmQTu/5+cpOIzhK+yzRy+AOLaVeg2JyrL8ZflAMaB/lbKwa7u2/tD5QkzFfTs30BD
V6DBOVFGMdcQQvIJtdgnrVn13Uv7/yYXTAjgtKaLjS4LVCrv9x0a9/8Yp4XkQkn1SlIdvAE0XSHb
7yo+sQ6pUZHx+0R/Y3X5PU4Sj2Jz71T2Kzdu2LM3fdkddeMfp5rFVfIK5lOrgUPAK1HL50pKkC9E
gU5bWGzPKrDva1pSHA5afx9gzSPSv6gpmR/tEcw+LLYCRM+q9pGCAMzjwPDI/8Fld+f1Qvhd2QKD
r+t/1sSS/S37tYyKpBQHpTCvrhPBw1O9IH+N/amGgyrbiLzdB37xpKiC9xGXcSzruDCsIs6/LBe1
lgo5OCvZ0bKOPD55k47XCEXAbEEsnn80D6sD4XdcNk4J1dTSQ13pOdobZ/1CqzIDKXxsiH3nsR9I
GVbDlA+IIsaEbYl81NfZoFx9EeukDmRniPcDdsIKMbZAp/si6iT0a06BGrPfSfPMDXIaI4vgeCeu
hj7adxbG4nQ+3FSwIfDrutKgs1G8ejiE/ihprs7oFFJ1XqNdotK/0gyMP1JDJ2G+EsJ69T5Wghe4
Paxs8CNMcLMT4IPlXhFeDJKSFtykhu3Pupaj/AoiAEg5posRIZblnymfS87zh2rMwk39V+19wuCw
9mabR0GQxRKkabk8fZ2sWAwQU7gTOkncTcJMluK8u/sB/xr9qbAasTqdHsuKSSa60HZA003AC0AK
feLhW97Aqw5+kwMlIz3TQHb4wvdHPAEp6GiVDbME92dLQTQqAVFnBv4TOlZnyOGdSn0KveswAtiw
SmL5CEM7JjyYhVxLuISein5xMbSu72N3RWxeHlAMAAgJrLZKVd00VLgRtATaR1ZZRatLxmyDVVdX
tV1rx+zx0wYtc1J5xsKuZj6SQEGxH/T2XP6lNwQy1d4ckSys/p9iAMXUkhuKX12Pn5vZr5esCxOf
Agi2dfttVg22/sKWBFJuBHKmhIVsqBnaD+BJ7nbjFIePpmRrbex+VZ9s0dUlyjk7EY0dVsUxxZg9
yPReSnOgJQJCukpmAPU8r47KXaRZAKX8jpedYlwWibEGD1Pfac6+KaS+tWBhtsVbTfqevwGH/mh9
FDemswnS3vNWBigjtc8hjrzU26doJZYrglKkwtBbNDuKQwG+5aQNjF7haq/qL/rdfitASnFYSbAz
5a3tpzXM+EZifNHIyTAngjfnvOLcY/WnDKf5J/BTdG344tx26gBYdimJexFHzbN68ttWcsG3VmVM
tXHvWytcKoVxCsQoEMxE7InBFXGLp19bJNJFeVbl6ZSEvbWiEn/hfJjyG88baiuCAK1F1CX/eD8U
XPtim4bA8l5oJpm5v9YvHHpNvKtrx3lt2Cx2ADpYhhM6K/uUnbvpSzfcoUGy2NQ/ZpdypmPtRIu1
1WVfHOdlrFr3O3tFSQ0+o8p+pwoyA5pUyHjOzvTZTNokquFS8jitO1GfQLqf1128oxZTXKFvunOD
NjCgEeEuSQ7YZLaR6iePBCAvmyo6V0VouaswRjHx7tzRb/YpVxApXpz9KzM0VfXDUGt1Ep+nVDJQ
7Zrmp1MIFMJqjFu3bx3zyt76LgXYh/76ckurI84pS+mxonujhGs0MCg8XMGwAgO3uW9Oq7C+NxKr
WE9RDw5p/62tSBy7DWCS+bYwQ0fg39tKn/5garQaRY5mzP5bmt8+tjKDv7fKKUli5JYccUcgOHDg
PaaWQBGFsBvX13uRWUGhhRiUVv1aLl7/x4XdEhOftwCAGIQDSvHIa5egtUnJVkDmQrOMTog9uhGj
ZIrnteD+sWcQrzogJ23LqBfk5+4kreQTdZ1Y9gqgzBlNMzX9R+eG9vNjWsX79vt/C+Telsx01P3l
f10+YITzG0YkRMGFq9sLtdo6WqXoaGao3wDAM/N0vfaYw88M7VZibLLwyheWhVGbj/DLMvUCSoh7
5wp/HACKmqW+RMzYXQtnIXTPWtBE7WtK/AtFt4BnOFQFOtvElM7+LebnVu/05EZwIRtP9Cxew1Wl
mGX6C7U7EvC5EjP+6dnYQqrWCfafS/OCBxgpLM7yiSqHVbCJ88wYVgV0PPGxGYMGEtvLOP0AsKD6
SxeLj/9oRSyB1FexQy/hHVpcb6mR7fV4HoFJ6wy2804pg6uSRW6/qY9Kb3osvU/jQlTFqADT28F0
yzuEaCQ8Z3Mk5lU0YWZjgWYLHh71uIYtPQ8Ah5kjKQZM3/cgHu7mtnt7MsuNZanDqoMIorBJyzN4
kHfVzOmZHAu4+WjFI/Jr8T4KKtBqfGM1XJ+aQHiiyU/vXBgRExgvt8tK5Hw9qhTB87JKQKcorFhB
zQQr1lV/NdmdzCyePYh3ZRuXh2UTYPPkzgMZQea0CniHbxgju0JHxZJx9Aku4vA41F28wdNzSw3S
UXBV+ejVacZaxoKE/ZeubjB0p/AqyjamUssX9+e2W98v7mqR6JZqio1FxWKjH7OJF7tO8kS48urJ
6Ool2ezudmoAzuPc3u2mWctcxWmRgUuO66GlFmbWECcnu2IlhkA+NxLBiQH11aI7UMpbpV3PlDIK
LscZRkch0nrHPGP7+nGu1CKX4iDbO/Q3EJWeVEF9OMhDeut2l6L4y1o0FkFtAu4AbDZysqXkP6xm
R2EcwbiY5wd6hpllmeqxiZiLYndZhVIQsVpkZSXKnqP9vFklxhQgEzgA7wBkzy9sS5GLlkUt4XaO
G+kpi45aD/+kaUJfqa9wjyPrQBqiBmxz0ZGwEztiz3J8e3d/V48G9AIucBDvdRlbBi7AODFFw/pr
ChHVwb4R03hWNMvhLb5alFRtzyA5SBXoiFeRZvmgeu4ilsQ9tTDAm6bmxRzn01yytdRDGwYz36Ue
V1oWQLxrBy6/p1qcea8D6+sUr4AbcdYLFAiRLSxE/0/LmGCRR15Gg4fItkYFNZ645PHoQc/gSP+P
mIssiufDJh+j2AiB8gmcgy5NEFrS/yJZXNIjXaDpDxnno4W4CpXDlC4lH2YlVuM/zEZ0/7BDIov5
druPO3fBB8h7NNYDXepHyWnxB1xmXuf9Jf9m67QwZj9lL33fBWR6jjvbfvmcxQ0dIt6PjMIC2BPP
PYq9VxHvV2r6DWuHNrIF67HSKp2Wkuy/b0pjFH80mB5A8L8XmESLrJz9rznuNSaktdBglsofOF5g
7qMGp34/hxnwf7ySlL8J2UfJwnoGcGOvPpq1UBMyLISmi3IHewcp7dHyeIBfRi+wbuvBZoq11XNi
TwFjtmpynDqwb/venuesPOb6VydVVkMyZR+Q3N4FeF3O3zPqUiySLoeQwycRtx6ywKKB7VsU3rq8
wbLvfuSO7MkNrv69QNi1ynAVY9VOYFGAQD7jelgJ94usDkehX4AvOmqvhVfZjx2rpPc2OKKejM4Y
lsV8drP2pbgT9GGzQrwsJVg4ASLBVWSnnjhaqFCNOP+nRJdYjt9+OXujzBipC0KYryRTAQLzC/fq
3/jI9wdxhva0Fj1vTOJkceiIdZibGQPQPLAgIVbupkMgZqINnZhwxIk8kl+lz+GHfyx2fmm9cQ/q
STPCR5tBE9ipNbDKYmI4Iz5PHF0TxD1hLmuyJwVcNMtsoorXnp/ozCpiiK95sWxXsqSJeYs+b2YL
ZWaxY2A2nkO+bTxWzv2WFluGqummaAsxyYapMIvD4k+J7re+6ZtiKokvP7gBk0X2NASwv7689JU0
enYV7C1iyGHSC/9Vx5ebA8m2SAjeOvcvZCWstXAZ1+P1X0V6ZIqm5Qa+F6op4ksaa7GDJ8E8n1vi
egGY3rO+P2rd4IVwWlVBpqRQ46Jvj+9UKano6OwTh4MH/z5j846fapCExoEq0vVCKkBfqOsPJS1Q
gs69eBic3JkFZD0n6ZTLgG6kBMLBh50FBenpxtjznq+VKqTdY2xJWQme8UN4PoQvGdrJkGOLMHJk
HYLLY3yUBUaQBsACmfydDZ8hCn1eHCyeuTakyGCnnP0f08X/lk9Y0u6RYKONfq7OzktVeXHxUCJK
xGsXttJLaJpcCK4O7EDnB3C/yyLqCWvc1kN00SQUKwcbL0Nry6xV8z495qgfxEJeZNXXqlqBOmbU
2lICriBmZW3dzR0mrdJYnKbOyMcC9HcsrjzxbktFmmB3fiLFiB6+wrVRfQH9pJaOrRNYLlaY6tKC
bturdl7axy/61Of4kbvT86RnAoxElsq0aARyNTStewfse4xm83jV51YKDZQP5Hb1KgxDNdtErLIZ
+hiCktf4CY9fygXXtr5jpG3XzEWDR1Kk33sA7ftdueTn8165jKhOr/sZdMT7pDHP0skWLiIciC2t
XGVdOu9DVVqxCOKpMQkrKitE6K68AsAt3rZn3anmjOEmDHDkZfT4CWtthNC4dGnQkHRVJGiUuKBE
UUNQ+uGa2S0pNcONC+PaLROEiXBvnBsTN51QrEQ38U9zE0iILJdAYXb0abFDGlfoHs9OO0uC9bYd
vw76kGILWPwylzZQdU1aN4lkA3LDvl/HpJ5Nhb5CwZQQ13hVYaJMIyhhuzUKIuD9eokQcNik8BY4
rEByPsw3Zdhf8xz648flR5YiPz0e+cxip0Z0wcgSxf39h648i9iwajhdeHf8S2oocm+iCeUnt3QV
lGUocdeNwKDRF4mJNwSC6s6SWw0pfR/QxsXIBpwkU5LdrE8rAp4R8y9fu4K8RxAzk845tNGAO7sK
4xugkZ4H5UusgZtntUsBHtmXWa2VjNFoFKpHf346CvcpH9IqK8WGXlFuQaG0R58bduBtqQ35CCjw
PH6Fq0iGD/z3/8UjNtlqnTehomFBKpSxSVzB1rPmjHGlgv+YU74jExNEuo8rVQ/jx4w54Yv/QOYL
hMuBo+aQjU3TBWzKqRawHWTnmPaVvXdz/OWltbXMYmCS35sj5ELCBbOgP8F/+bZwayucRAWTEbVD
DS9f61Fihsz/kLs7yFslCLfO66cZCuJJY2A0DxubJ1W/nlpGOmMHjpBAb3NWIjXbhMV9xPiUxPad
fDDgW6dEnAAH16hP3ZG5la0juSXrHKyD/rA8A1LX759HQTzGULVCpOO5Hu+vzwscy6QF2TKML8/f
/VHaY4u/qlK9mARE6Z+cYH1LNM2kx8eO0iwsrRC5n43nym1odUXvB1aIlg+X0p+8TSjeVVkneecd
achK1CAeHwGbQ60an+Liak6ib4Bb0GSn18i//w+Div0OVCvCqHla++sl93XtHhrWcLNKkiXQdtqS
bVSaw6HYEnas/IfznsgfO9WtLck0EQaUhC9qgMyJ1IB/m7c4rpsAhQ+mo+EB17CEbzguP3FNXDrK
mdz2cibokXY0EzJo3QOEgb9lgK8K+6e6eUC64/Uf+SRLyQeLFnhY7WW4iOy6Qgk7I/EDl5RmvSxz
R3MrQErtCBFqgA/Iz5LzKS07jybrXIZ9FE9M8akh9JK++mTKI3j/YDmp6daREcUN+3DRym6TCKsK
Wxz+fg0NMxalzlWKdEJYPcMHkrqcmlBzvlIicnKEv6A0V9K+VAkchVEYWMN9r32rABCKcfHgyF1W
9C3r5mP3LWX68rB4zRYGEVX6cgCs70AVKNx+v3xil5Qae/rGYmj+CEI5YVBdndJYf5GEVDo/MRF3
frUBHPSsT34QYHNh7RE93ky4sFbYToVX0pvrtgAevvLHeK/tLFrxNioeAZ2rEx9ze9fpgQdjH782
O/Kc5Go7M8xDReLHY/dgaBRnawE+qMJmRVksH1RVwq0MV9h75yGYMrNsomAeFcq8ifhlSIVV7h/7
HsMNypLw6K5TNjXxNK0lEDMEp3QxmcpeN7CqiZW7dicsfua30DF8+DDwai/RozDXWGLfLU7R8TTr
hDxKEcHhDu6+8IHLYV3ngReu+jgjVK8jHo+1B0UEUDzVxUg/Pg8rGauLuNTBk/3eyIx4LCEm/yRG
9drXxKVChZc/UY0+mv3fZehLVHdFgr2ayzDa7xGVlyGdrr6g5GlYgovbDlUeMly27XgEEdUekfKR
jr9JAz6qlvRUdOVNAxDaUjESjc2xdrpW1a0TuLwHatSS+VbOIbxoFo8ByGxP56qxipYQIhK6skmh
4/zaLl65ejk/HRYwQ7N8tKdvlUDXfVlziTisPAFQ8bgLG7ie9hUmh1z+6Kk3a5yj/I2twdK38ZEN
9sLekVLsr81Ka8HLmPykD4Ji5nq8U2ARDbZex5TTQLbVwkMc+chNkIuLngTNzMOcUswzpNrpDpr/
ixeFfxzPI/L2hLJFSoZP5VrzaRgT6qy/8GwZQ6u+jlj2MUdl/hsNjXgno4mLs7y0A3iAacbOvk7W
JmMPlWbBj864W1MYl3BCK+mPCRQIx0mYI2Hts8ojdjyyaOv/jqP4PNgejsmFPvyjWzTJLtrUh7SC
2lgGWhkWOI6T7ea52fqxy0fDV4FTyaNmbXH7KJ8j10yo34eRgoOoLD1++Vut9O0jMlpgqJv7bybT
9gWm8tPcsvJJdBWgMZzl2oI1eMhTfk1mIDum+iUcOCKKFQVLE+EWRhaYuWcAtecnS/jBQarjwWSe
Ah8vETHgbvV4bAvGLOjr4r1xy/jqdeJXnX33rfVyXK3k99oW7rBy4tXGkZQ24eHnEkWLzYP1nfxy
oL58ypJ09ENuAFRwTAj67sKV0Fw9K+yVHy6b2leASy3rIz+OXudLwiaLfUIT0S5v8Js+takgUQOm
QNsj7sRDoKpaV5O/prMrx7iGliwP9yEu7Brk9WUSG1/pM/atLP8O1Exu9sI98suhuerBJB5McIpN
kUHY262W/wLV6C4/ZUGZZ6092oJCdqfFWd48marKR34yPme/QdeTkRlz9mONhtxAt6akF7KJChlX
FX5hQ4b2ojopbwuNl4tUxwf/KW6shEdsFTOztZ6aiN54s0AIffd2Bog3n+zUuY9WPuQ9WDDiUrqD
n0S+et/W5m6FGtz5FI2H9k5M2kJ+yx39c2cAjQmQ8vVDsHkem1mp2N1O+XVFhuVRTbmXIUxSLu6P
wjqiiRldYVqpRHilrRSOtD0L4q18AFgRUSbb8pyRskpzH/32p4AdQsNUxCz4DjNrkrQWwNrlY6+q
qkBjVQAxEu+2ppAjhqcCOhnKxW5qZs/3pAR6mp5mobcYmLVKP0z1WD4e9XppokTQjC+FU0F1curQ
5QMaFsoD3vzhU/WropxXDOYZSQTjbGP87TKXGdDGJGwtCtuAmpZOepuM8GJbmQh6oPVbMb57w2lF
JCWe3EoDQuOvvvM/F6iyqTkQqLvM5CoZGrR+7HTya90WHGorPWdGL8wubqq6GyaNSjXJfXBd7JbL
9oeqrM/OngowlvbC2CNo8i8RKqiYg3n9UTQOCkk8hElwssV6ZGMaBc+TAPLeUujwRq8h0N99I4tR
SHp7LutliWVPyPOCOH6s5z5s/Otq/dXnqbOJ73ACoHV8vjydLkITTaYvdNR8LzZwf4USGNxoO+Pc
mMrRa19JeDS2x2wLVm8e+CUqUogXffPJgxMA7aG3mOMFUfXmp8CWP9RMcyK5zE4W95Ae30r+UkiM
muO7v6jTB3guyNZwixnUnwG5vAlaIK0nhzU5d/Mq9cDd0vfWlR/rxVD/YprhuJT0NSuDrsdndsPS
YG0UGzKks23NMD3pFnEMQAtg3fvtn0ZGA8Lj2UAxWJppo789DjcD6qTyRYourrBlWaRUWwzf61Gk
qtNJ5RZv4a3q48GP+LQOSA8uDOVsBpLPnb1lw+MYFRC52M5vSOAJji/1A/kwf50RSN+nF9qKYjMH
FbTp4wrHcIwAxGTMLujcInABkWS8wBdoNFK8t75FUBbpQKoGsMbaqsdSmhcJqHesmyKALBJsGN1x
WHTtikoAjSVRtHNh+2LFkxtm5Qv3JyYfAn6fEAgs/aaRck/Y0Mydma402+Zqsp/QHfVgOSwF5Z/V
6DUC/MpXtsbRNqfUkr75f/nwQJcfrvWW71A6aebB/Ps7KopRVRd3Yx8XgDhMRS510M7E7Cr6s5eJ
W2fBLEm+YeMqaQtHXuAjwiMzv9bcyjcUpv7DLzcJj5RODcKrZYhfY83/gAhw38lPQHKS3tjmvJp1
RAD2pKvcrfHArqG35U3ndcTJ/SgJl5NaazIXyA2SpEcW5kfXkdE0dfuRuiqG2bdY53P0QbnNTVWA
DTIpW2a6ZZ6aXM1GWiZ/1RqTBd5F/JgZNsqmiZ32diBpvZweeGGTqrscxYZSvY9jGJIYByvtBh8O
d2lbQIXn2HSBtIDH3Uv/wBmgeJU6tcfUScYVbPUExYKHBG4KWkissF3U2FWeHG0asuHzZY8fzQ8O
n4HmjSXB+XCL4O7L+BVH2WnivJfc/sR2v3ZWXXUmfyMnoF1BqUkIqoNPpkOf22PwBnIxfd4nFp1C
CuGynMa89zpo8o/KwTek20eb73oWZ4w9gbE7Z4qXsA+nSK+6gTSixR2wxedb/k6L8gHOqXn3uhWX
bcJcHChx0ycE8GMy44lZVGOK869x6Hw+6odes9HukimOHJVUshLe5PZ40M7t9+Q6kBPdsHMbiPad
vNsiJvbaGzyXpVpJN9s5u52gzZfoxSsVI5dqi7F8E+vunMpjyNzy41c3RqkV8D3yibH64bkSVvth
rU0roSZWI90dbNIBSX89nBTR6w/bj/MWrqTkZv425aSmt8ufqTWplSVFYp+q6VKBGA4odUvclAdY
FxpSkAs73h0lF7gcogwPnV0bmpjhD9KP4G56h/GToYL5vpxDT+ovVnaLJapkTt7tl+uN5L8tMq2E
IdNYrpTYklWz+ig1tuUmQjwlFR1DR8rhR4XXT1WB1P8EYyFFBjxkKCHYCHxepLhbk4EHRDXheTOx
Btekoc2+XSsc1H863RSFMC6+h9NoqG4Bi/30Y7P3gcTzJRfwKZ35Q3y9uEP/LWQKr3AEv2Ss+vTb
+eYDWUrDyV4wjoSY8xZMv0I7oQvf2mtVh+qeoOQonU5NUfWLflgMr/vT+nlsbIqiIvwygaInyzDx
AZ8T/4MHYxMnhHI6P01CFKdeLC+J7bWFlm7koY+wV4RD7u8TvQo4Yiq2fNznPiFIS2PtFAQXkfXD
wAfVzwrJLd6iG3/Oi/J7lTRoTwOH9j23HH6QEq6hrR6YLJ4dr67bOWWlYlrw9T4YungLtEQTmKFS
4zovk6SQSc4m3Z8EWXUkm1FjR85+xE2YIQKFQVkI7shnL9xKSQBoL0/mymp/1ogosrNucnDTsSn/
tCeu6nlAWSlciGjdaf/1VjpsGFStonu8Vi6CTX+9YBm4cB0g7Nd71wawZLoN0DSK+zWug5a1O6Tt
LdWYFc7sCrqVNFS+3gduA0SENAMyKFPL+9NoatcCZjktgQh7nwOcdKJ2dOIzFdybv1rRYipQYaOJ
bBMoOm89IT206TjwNWAQCo7ULa8nJjWUipXR924jAad5v2Ne9ade7eeT+MVvUbuqsZNcM4isLYwM
HMFzEoR4ymFWqADeoufAYhkTHGdvR4qz3cxqNoSako0Nik93NR7bHWtOPFA7ZA8RV0IUX2i/D66s
GxO2DTez4CHB4Dz7WuQm7UTPPFIZiquzVOZKz2aCzSnBX7gUGI4xdnqiZdeurac0YZLi6a5JZiez
ChI1dkVNIq5rTcEJyUujm4My0i059orpSXrXGQHHr2Xovu7TC4U3Nae9HEAud+jtBiBc2L0DVfJa
v9XC91ZfKKdv93Q61xmMvrTpo8ClFM3s6WA0nm0dbVlK1I2Z0xJ9Cf0eOWfN22+rMA1DB4ZG7QAp
Tx0HhfcsPJdV09Oiv6hdeu9cKaKjLPCWv370QU/9GGacyxFTtaReatDxLA/6IdwxyK/fRqTd3FHF
fUJx+cKFb6wqA5MLzwMmMdnxifXtiH5XdAWb61I7rQXvebxmrXPeHR29SqUK1PpjxhBMRvvZyjlp
lPo2bT4ZqACFK7D4pmoG5kwCv5MCL0YFgv+7QG+pm58zNK7lxhH5hVqw1G0AtloHPXlNjWHYWQnk
c9VYfIZQh/KyRtU6TFkcift3+eLdnrvkcLVCBvE9gQI6yNAIZAMIZBr2vWm/gvDny5fyEeosp9OX
ax+zGFK9pfgPkzl9CtTto+VVybHSe+hYkaqglXsVJjkj5N7y9t+KVgY0uoRd0RlSE2YhCAnsfkKH
VGrf8qu1noAgJF3z47KAjOtZVT2K49t8VIBEEBgQzV2+y9cALyr9ztVWdCuY/bqYWkvSIOkxbKEt
0fjddx9xvZbMNUZWZfK9cC4UAdq+3j2MT+PLfuNLcsIdlGOFcjIDcCSE1Fd2BuXKvPSK2J+nZWzB
p7KbFC4KMe1c7FWPrLJ+n6WMoXS48G+oL3M9uuK5PMjmHswlSs//kxgF76htGX/CFT4ZvLcjogcs
LeX7c1NzLx1Unyv3C37ii5316RwKyXdcsaUj8RbE4uSCVlVVW0aCBPCU45vNi28Luz1PXY3Ap2Fv
YBsppyFhnah54SqzLBo0ggzQd+xGy8M+KdIqRg/RQ/ScpZkzKJoMhZMXVDhOIQ85aOWHpqjnn3qe
rtGEuG3rCYjDur/0BNoCgIuqgOiozc+708G/vbkxG5QLwJkcC8aCxB0/4C607Ox+6oNrrIdhy8FY
YI2QL71wdyD/7WnarKXZkoDBSQ7ZpOY33JevofeKPrDR+025uxTOxQMgjqZQMw0SuB40YASVQd6a
rIpTMU3yuUQm7/A9XbBNMKTcSR8uz8FHVjGEF4tmH8ncEZQfOvsAxT5CPiiVhKlMYsQpVOSuXPWP
arKTBaNCHxnD5vVKt8AVheJ4dnZS2+GOa4bGUovXdHEyQTzJVqPYYrWVcF8JZhEfZTryRr/QNR+p
oUJHyaBY09AtWSdXBYF0r/U95ZCMOIYFZrVn+SbO429za0pxAouM6Qn9QiMHAgjG4o/f6DgcQgfu
/n/YCX0FjiQvduIA7aB2+0au6tqOcq07eaoFVIOMLlPw8sMRfVgFmfeLXSZhVmkwnGlAw+H+heCC
JCx6jRnRCnN82DF6bxUy1EWIEcuCgs3DeDE3AeRb+LshBNE86js1X51gvpSb+eXaCBoWZTLhIYXK
UewJHAhnzbQAM+oYp6lYzcJQvAG8JLrdsZZ9p/JUTGJ7wMmNOBqkCdWqcGNHODaIF8LC1Bgx+6/3
/LqBVMq15EqFwjp33Swlgn5Mrc4gV/P4pGg4rLHpFyV0HGJGknOUXGE3QM4j4X4Rm8K9uboehh8p
Ap2PtGJujn2R5cX9wDZqC5kneBKb9C1XNja7OX/rGWt1cu3xDGAPRZ0G3mwDQCZEpWfF6U/yR6Zz
cS4jEji7OpQsbmmkJKX+zIpI1rq6r2RxZD3si/XcDB+x5vp+aUGS1ldf4chURx7WAatidIoB4gis
F1vB5wg9HwyEky9heyA80NZh+X4jfQIt68pgshwtx9T4GGDlgeirFQ6xt00cdTxo9tBjVtRCrAO8
TfnzFilD0+GEogSmYEZ6ADIRBZ6BABQdOrJ1X14q1kYeC+YwwGYRQXi1K/eLUclvAFJsjB6DXaLv
ApgSP0+0dYVTIuVS85xwq1BG/biq2JzwXlgzZiAHuVN/ADtHhJ9FtWD/sXurxp0JhQYRWyAG7vzH
66uoAIwWU+8CUXCkZA/3tW+PE+66O6YDo4xDS/rDA4en4w3BwncMfnjjjqc8GWetmTGisNwa3STA
ji2wzTLpjAsPBhebXtFwX+uA8WGKOq+XCBaBmloFYVC+8NU+3qzgiDpGK7+2DzyY88pll3qXhczW
P0XcGTyvEkx7xGRk0K9Acq9LsFg4i2Ihpgm3lljRpqzVAexBm9SVfiE+8jet27MtI4IoWYk59Sdg
FqqOrTpFAksmoR4mzncxMC4srNPxRJWG4waWDfntFRE69etv+KO47w0hhG5026yLpcaojUEWo8jW
KMtg3E1MjAKYsiJnvw0fTfdNvexl48dNAyRLSkYnZce+jR8vi4cwAajvP+NxliU0BFhRNcQ3wMy+
Jr2eIx+P9feOqI3K9SEZ6PzJSBwhOrgeyXiH0PUoUZWyeaEFG7yiPgq0Vs0T3OGtK/ExLoeGs8t8
95FgYFLfjyFFRnNSWsErEDKD9fDtKy4SjWsI3m89JYLVnrQNushld6YXq7410KzhnDJeDIWaHT8r
Huel89TT7Fstek8hSgJnz9tDICX7EjICTtra+hvLgdd6mhCEQSB5LXCv7dfdpmc6a05We1996c5X
g+mbWU/JMAnvxNhXUMg1S/3hy1u125YpZvIyjX5mPsA9G61njXn7wf/l8ANe/vf4jxC+3kE2B6sB
quqmybF8T3W9FoNGpvSGXEzfbRKEl8zXVnu6/G2C2+AjRtpBm4kf6a+SPNjOahse3x7WrEq2Dbih
uLAw4oo0eRUp3e3rwBXxO5qYsNWep6DURE0KAQjfpVoFuh1D/tHNB3iCpOW/af/vdhJozbCcyWWZ
64bIscusGB2ehKR9QJ3IO7T+ZNv2fxqXQz2/0U178DzxZDs1XVapQQLv/ptF1PQMNjLS0G5kMZ56
benrxqwiwao459+k8V3w9yYa/Dh+YnMUd/gywLXbNzEcqUJL8I9MaVwNf8fi+rCnYTSrxLR2pkNp
aCkomWnZ21zJHACgeOCJS3t0/ltZx7R7hAST65qjfZ+Tp2g0j8hVq3sGZGADh8sXO4xKi4OubKAK
KehWocNbGATcPUMl6zjFLD258Casl8LGzbjugQKZ7CKMqJ7EhFu6IZ6Vh4BVUonn2zpEeyeA8NEX
lG3lgFT7nI8KMcg5BsIF2Mj41BwqYKJrD4L0Zt+lqA9VOo8mlggYoOgUL3CbxKBf+O693FZ/gtdn
fg3XeG3OTr8F0wms06OsiDbRyneUcoCi1YVXhcpd+0M137A3Sc4j341OYpLuB03coMOn2XfU1oQc
jczNFJawea0FcIb1OGFuKW6+YbE0MORaiAsF9KbEQ94/b9vjiPhx0m4jb60/hg57nXJBXW4NEU/7
tnn7Jqb5aoeFVb02Pf1qknqGWStXlXwGyglnL6P0H+8vuMiz3qvoE2MkivYXrBrKC7+9OUriutZ8
16G9TlIi0jXP4zFyGIii9+C2L7hiIJh4vKTikcR2RyFxGS4779gU9LRw0W3MGEoJ47PEcaZjaHS8
TlOSEG/msuEHDQ19DRjHZTSjlbVPd/c1YqNMogGyQRb8mj6xmMKw/miwPobUDz9WhAu+iNNan0MQ
Zaw9AIPNdK5tR0arU/JqzCYRMcfoIu6zW6uHtX6BgKKhnwRwrbziwiapfJ7k9ixLDYQSSCUiP/1b
vfXEagoeM/JKH+eBpLb3amdHwWBUFhJtFWot3JgPtNRP+BKpXBciAOXioxPyH6KQgRQrdMY3BjhW
zcC3mPAzJVRDNOmV5u4FSUG/DOikVOV9BxieH/SocNEX5rVtr+znXgRHnzstPXs44PG0Gs4kBJOG
qYghQepnpZQ5lDJv/GWZZd6gw29ObNYAtaHCQwlvGz3jI6sCQqMqfqPO6mwXwGpGp+vQuAbD+yCT
Uwmh6p3tWiMwF3l7iiwWgWhntV8LWMvNWQuzZWuPsqnZzM+SvYzzfXDib6rlc69Wqjj1/WTmOHnF
X8aRt5Gfhz5pyHH3gxVO4/XNqcSnUoLAgtlPe12WwB0vK1VJE9CF2Hgaq3Mqt6QvR3fzHdYeRItp
WFtexYizwbwLNG5urHheRhT5nY2MgUiU/0k/M89IThoP6ZKCpIxuVFK1i88bfC7HRoeSUo7+SyOk
hziAEB1IX/9SZ0HPcsYjJlyceG81ziLQYdKOi5D7B+MvRiTIpd7BbwPVA/H4xvEEYxoJsKgZzJYE
N3ZxhH8TVSlUU0rdNc2aPn4sdoRoqJLzh0vH/V7tq+miH4Aes3C0IIHSJrnXtyZHs0hb08VFph61
EyPLx0Il0n8MHcAQqlWytxk/aUIsLFuQ1ckUCP2ifSu6UIkFnz0LyfkTYmy4SUV/ry+nube20NkC
NVoLb986e8Ot6yS925heqdctNxPGXispFsnmtOT2Is6VnFLvbMhcqa8Q80/VNPJec37yx4UkXEZU
CNWOWV3wgjOUC1jigZ3gaY89ffmAA7KO2AgNWlLKdsnxzjc5UEn3Ddi1WqXhVw6wT60aEA0uRLRe
jvmiIedL3TtdYfprBJ+yrEr2SdPMP10Dlz5/v7CpjaDElKMlDpFuUsII1FvtO+WpQfdDZ7llOWTv
UTj+4IiF+qgdNfWY040ILx7QkVBLIJa6gtdSRlhFWU5vUyUXZ9ITsot0Po+NsTqo9CquwoVDXPFK
vXVBriR6shADgbIBXl/XTJBC1ezF2YxzWgDed6UeJmUumMagR9qECNYTueNasJt9e8Ma+85ogaXw
11nU2wcG/t9Oj7ImIiFmwE6Qbh8dr79aes4G5abTL4X61tL8mSf99mETeF5so4eZCWaxdq6dN9Wa
/4z4FxnxAMj36Jwkbojahp1I51dpKeHFU4i3u5mIyHJC121hWZzCWSX6RP4+SwJ5UdJS3XvvFVyi
Zvjfq+RF1BARtCnOWAIrphyZtBwXS3rTmBh/raaX+NipyJT5M4eNkJq1V5WWkjDe16ukeYZ+h9aW
hFFjBQxzNSei8heQ7K/QJadLuQgN4ixXZ8Na+tMRqB8cokzCeR9OnSK4LMAAIF5pUEma8dDpnCSL
9Ibdd8TIsBRYx59pFhIxHRdoeR3Ek3GW3FWBFrUnDThaIS/n/+f42Lxi+cIaXvPvxda05N9LQ3Em
1B7U1gHhJPzMnwejV6hcQsZJJ/U5XngNv/mj5v8dJrRPQjfI3NmilISQpiMP/WbfZSPnZJXxF2QH
84AxLLJwGNh8uoW+d6dQ432cOTYgSTbXtYrP9H+Y4l70ZENBj91BYu8gGQvFOfDh9etEmNRDusm1
sos/z42h8vAN18lvHrMCVh1A4BOcJKrnYbHWzJ3Ux0CT2dp8koisTj9JMF3jhU684sVsObhKgC6Z
ag3zNyuvcrs7ubRLkDhkJhQg0ya7S7axTgES+tKC8tAepqK68Z49YrqXwZ/JCOhSCXEOr++c+Fze
u7vl1kWV3zpbaH9i7ZA8jogqD5JzmdYcefumsHc/ph/jU3l3vLPsQVraHnQ1fu3JRd/Xg7TcHSE5
QEv0ac27ESwa+F4BScMkfHgV46OGjfjkmNBAK0CDDUSKTQCP4yuUVUXeISqkEkEMOnkKyDBanxSG
3mT6uGIHOxdF+6qOKyaF91s2zKI/axsiXGlE8TN1y0sYcBKfVDPmLcfxWfze6492IFvJ1BPCKHyv
VPwBd6XjUlHuGKu07TJIWaSw+3bCgsSugY0NNcSi5jol89KN0qJH8aNrRe3AQVnvES+zLo1Rlpgr
gF3RM6lswtMKbj650+syUWR4tkPZUI3/dyh5DVP3b3asV/JBxdvF9DEFjhiauvagP2sjAcxgqZgY
f0EMsK9BunxWnTctUu6qwNP1nXWhJdNT29KcsBK0+l2Wl6Qih8TSW516yusWYcXVLzHXvLTUEIrS
ckm7tzwnBQkUzInwUPKeuJmW+Sn9Wgm0mMsnBrYvg3qtsjhEhLI7XV4lipcSbWUZChMeOkR9wbEH
/jRfq88gYZ8KFTD+R+WYEVpJG6uu73hNIf8X+TMx/JNCfsJmtC7R/dw0cgtC/LZkxNUQJuykXohL
9VZoNA/rlwlq+Tr9TUEwRg/41+0vXoFmhnxqgS18Wiz7hTyMfZ7Kw80nTT9E+PcocNuJTz+GOW0M
h2aP4s7lInnhjdppp1vb00omAatX6MNveDrzlfz1Z1GQRhknd3k5c1fZZXrXOky9v3e/EGv+c9ZG
E4AlIlpIU2YRFuuep37qBTTx1Iqun8s4TP8NMD1gR1bSxPW1ErBpvY4cF0VXVoNdwJENWCELZb8M
YM+NAlLCTFTjheql12mDO5VUy31Se9iVCEeGUz7ijLCd8NB5Aetr8dl4l5yu/+QnOqNVl5pjeXX0
A8fq0AF8gyfASbHCG0gLJB+EzSgGx/OFpLuqEj5eQR7FQ7fB1mcFKaccqviwLRveH6WbXP6UdTpv
1Lv2m0/LEFQ89UtlA8bF76NIj6Mq3xiWKdbxccgk5fdIrVt0D2WkJaKw9Ax1CYzNNEC7ZggsGXta
SqqnMKgPPMXkq0OuIYhw48jJRzpGOHKaUJTD5BiQwRVxNTvP2HccEA/YCUjziTX4GS8Oqo3XnMzc
v1vZbd+uNpw8e3HstszLKnRxTMU0D0T0rYMjWcf710dkccNLcYcJcdP7Md1M5y6lfkR3v5oqtGy6
cAQF3TzV6ZvFLc+1EdDsumHJcR9skg/JoIzBVlUhZ+9E20C/fkg6lxNJap7whU0HoEzOCPrKNYJT
BSJJZd4eWqIrwuVdUjAGPD68kBYY3ylNnJ2o90GQwG//35NSgVU7MrYDsaIL1MrecrEIAoLqll/C
BgU4Rl2r0r4qnnKmTjo/pCka5saXpP9w7ujnAUsGA+mA7TKgRecZmNUSLlfbauPYXH3Qr1xotFyy
oX2a4NKxZQVH/kXYkydfJ+j6yV5pvYabeG1PzO9nYXGU94c/5iQJI76zEra5aZn4z5S4XAh24987
82UBXvIF+WrelGbF1Vpk2f0ElYoo/eZ9wWYovry4AVfnwFF42Dg8Vpz74/l432Yw1Zfj2z+/AJC1
LNNLJ37KcrOLFypQEp0TG7ePUEvxQsmlz7104MDcb5CPOguexlFq3+sPseaaoYbzacdyvvYFa0i6
qkfbCCMcVAM/B+12txQa0HZ3S+iMy0vZ/MhjFD4yJQ7R9/WfD0GD0iBcGP8CaHJyL7eO1KGvGzJQ
5S/TJuEgs2H/dpaDzYAbdAU/7EsxdmsjAjWUIC33RhXny5YpBCB+U4uTSxBppmHmeBE3/y486i65
AU8hH8NrA7hrHt32Ah3fwDIx/BGRtYMxjHC9V/nrLx7xZ4plwpmYvqSwQOpzGQXbk9/RpAHZSjMR
LO1r5ICc9ReGyzGFD4UKxc4ekXDOcP5MLh17inB39UJ7MvKUPg88OoUWC6c2fAQ0kEcqrdcNP3DA
l1IxbnLCbXX2H1i8qKATJ9R/4HmcT2/i7RkD1F6ftKxB4fMMF/j6/wMqU299j5tloQ/foPswldok
4/kF1GCIiGM4dsUJfYEYxeYsQPcejRQVFGIrAQ6mBvlJKAHRa5lpyFUB3bDj1h8FYLBpkaOsSGTe
TbJ2eqlYfm7g276SsxV4l7v3dvyfM321lbdm1MT2lp0GAo7RvMDYl60Ibo4jhlxLXP6XVRzo1M52
ahN3pIBFA+6VovlJAtfypGxkxFXnP32adWw2G/aGxUveMR9aBZETmTRF6eDfIMj/563bssWW6LMc
uT9sS94dE/SfKAansyoaRzdLgvP/QkAZLqiodmYxykbD/RzoN0/4iTImxxlnCPnFgSQoEb9RmSVy
4Do0I6FRmeAFVQODns/0PaZJey2CStp3/1XO5S0MogcWX+25oIGJZpT2hwYVONu7cjz+VBa7h7jo
9t2Jein2Pa6Qjmy+US4wXosEl1IyH1BFWPl2VaVGviQ1NYvnt3Rh1KYfAK8SWnnlpDf3VYnfjsZI
SqmbsmL+WG3Ssrdd6hWPxb4UfBpFWhOc7WRcZudAJO+HB9JI1/p+aFmKhzwXEjrokjCzvWNGOxfq
HgQ2zJEjWAywwbvyf6nrYxKOX3cGqT8K7jA77Cj7bdYpVbPOzf0Dzp5WAd3AP2TcytGykz3E4Cmb
Z+hRHfycPJws2dYOJsF9v9P8C7EOp2Lf2aKOer1bU+vMJTBiJChLRyTEa1QUYDO8CvDIPxPk9Le6
BghqCSUXPVy4JdWYz/HQXfTdJCNx37yi/rs1R4NWgStqlHM3hA4YsvXgEI+3pN39XoWysydFM/UY
QmU2FHISBLVSVRzTUr2PSynoOgI3UU7ffzO6jqiwjW0S/iADKejfsYE3QX6hrp353ffGXhxhsODL
s80pWoOtlLMqdBzf3NMhZHQb6LPbdGLWQ2LXv6OIifWZZzwGuzRhR/+hDPiTdBLjN6TjhvgdAVca
s5TWQ0qRkWMGbCf1USUU+B1jeypRJnOW0fq6Gvkie2nG6kBpqRaCatzJsqsp/T3Rx3Q2Cfjl8sw6
mt526Ho+bSzwMDRcZXcdqBBDTMVpyRzsxvGdsLyKXSO+3NfReL/0eQMtR2UZg8F3OA26P/IuWq1u
fKeTWQtXWP/xGPjqitFiHxpT9g8lpICAxBKyPAyi8R1t1M84zbmrOmQGel/03/Zsme3Jdb/2vwcu
wm5BSp2Hz0Oq6Tp8NX9a6k/1Jo1Awfdg9cFFkotCl4jvceuWh3sfmsL/46kUQNPRDySt6W5kSs2e
Qk9Tz2WjvyBsOskkf7oMVZFWdU3BvhbtVyQilHsinAA7oCmsQLmARHhUq2/6pRV2lhu5y9id1ALd
X045doTjINsd0bslgxms+g+AttcdIb4X4FFVL1vBcZxEP+q7i7vJ8X1o9NGJeXOYJ/idD1LCa/nX
RxD3xt5/8k8S4qjc2W65e9VXHbxRlAcYBn4DtSrm1wtyOOFZqdR5Hsk7EVjwZ7M0EWjdeufA8UFW
i/t16xnIoJDluO1v/sM+tRMgQAMN1D21Gu3NRo/XGMnvjlRtXfyZ4H3EVaSmR3zxtjLUVSkmTmR9
lumc2CRqMXuhZF1ytvNz0d4nRHfYbYheExqZomCAcbW6L1b4T4F4f6E2w3BDosg0b6nBLVzqd4Bu
jkh1nk5oF5CEOgVTTq9X/7b8suzYCAaUEtZG3J/kFTpJ4aP0NIUXaA0Y82uCRWEj+LgkiQ/vzooc
AdMSBbbZ020f0ErfK39e/vJOhq1FngMflZYUWkFa0KIwUiotgRmR0sF7miarnJwQ1Z43OWDiU41c
KSpRoVoC6G6GVhWurYXAuZMFpKi+3r7GxTxoS7xvSjQ9EZblfX40PmM8/1mBPL3JmefWdYeVZb/L
47NThfBeeh1f+/BMF7dnYz+1d+cPO1bbCyEP/wgvWOMop7RQJ4ixLkhm6VEnaikCc/rl19fAuuzd
YPz2tHnAiV7qYMKpF5r67+LXmwDolTvcsD/1eXWmbL/XSpj8whQBwEcRLvLVq7U4r1gbBmzutZHW
ksg9z421kIbMq8cgVaCHUzA4+p4POJ437ET5+BiHHLDB4toS2KxTic/URj6EXx557OBQD8WJxEI/
Txt9p4ntc88vTJv8XfOCTKOVYiZjoH2NiZukOrlBGMU2sctIgLxALOXieRIWh57HKNXupgiXIdzM
kM74chVoWNOEnocCktxPgHIxVQMgXEK2zw+4Pv2lU417TVIjkODSgbUqn5H5Zx61h9+T9Vf/r0fB
qRSkjVj4ZShGMB91wGrMCPcnTtYsETgs8hHFGSE39rxhnPBCsJGUcuFwGVgMFb8x2iC602kBG9Hz
SIBANKviixAbyWfmX0yhjyNf5ifbTIaP3PSDEIWbvU8FtsIGEIhiOIyAuqNoU5MwF3ZaK+gJGTEb
MPs+fWmwSW8KEy32h43Tcz6SglBUVAE1HfzGkROULbMR8CXPNuS5v95qCQDtWaM52D2QOuKZqTdB
dMaMGhmirbiSD11TQ6svPEC/60NbmjXzZPBqek9PtMH4ny3Y5m/bHNTeSh72j3Uf1J5bIo0n4O1m
ULk2l0ouBum9t5fnn9rTDOwVZ1FheVyTpMx0gV1NxGAK1Evaq0lOADEvT9Pjn7O7xD9Z1PzkPYnV
stTSkdT7nXrEdM/6KSFkGgLOWTiYLplfr0EHdi663ERubyVhnrtugo0LVlpmr/AcjacpdQ6mTKcn
9ycjAbqhAodjvVtMeuQx2yDalpdZ4cAFyCpvAvQSuJNjZeeYjuhBz5VTHSw17sRqJbi/bHzlvNB1
sjEVZutgqsHH3bB/x0OfvAs8neIdht3YEV64WFovqCQLGEXCZuAQU3AVbF/h6zMi9hSCRRPJu5sp
H8XoOEAdqQJU8wNdCwiVJ6HgdB4g5oMqlg3iH4JqIXZ76nUPxRIj0xEsOgUUxF1le6WNcj0xnApB
CzxnZBTFmaimARhD3TGnjYT8fz2x1/L89axwCUP09QnQXqMHvGqb3i+dJHQDX6W7dKK4z/bCMSNq
jD+pBs3Q1UsiI+ArG/rGFTSNWfdi06XN0x7uRBEymoPyozyhMVb5Mcs8ok3zyKr/Xbs3DpMdUNLp
NiWDKJNYZsMIFrmXyqiXPi5Qhk0rN0Vt98Z7jdMhAxqtHQxPRQW0lP+t7nGjBUvw+cEhj/dZ9ZxY
2XKPSI4LW8v7xVTOuourEIOQOEzwmCmZSbw8Q1mHg8QWEUUOiwHfHKC+ZDENKwU7+0Huo2pxHsBs
ENnUnA7TV73n4PzHohKkGC12k823L/NhBl4wvAjOcNSazsUyQsvfRXvkOQemHm81aRF+jQddHvvF
gVWy4hkJCGh+OYCAjR0uWQueGOgXOoMchVDXRTQel/okp6vOuQAtwrB/bmTdQe1EF5LCPZOcIkpb
eWMlinljyx2lA/22Tn6ahGGfqSm/GQRTjBm5jC4K8qfbloSE99vVlGMYfRX3gtvUbCa0/4UCjnoM
pE6N7vgyZqIJiNBn03frrfaZPnKdx0sqABGWZwwg1z17z3ms4CI5mF87LoAXNrBlEhWoLdUwZMqM
jLolRUZQAv0kP60F14ed5upNr9m9YhUdkB3AysxYPljzeRhVJCLkV9OKzt4R5ynlUDp6z3ysFRWQ
8Zm9CL0zpUxAR2oDTURubi2wBtkcSCG09W/KqLv8O0QrcfHkNVEbOKGrQUtltI2DHmJa5Jat+nhP
5LN4eMGXvW5YSBYkTLokjxVM1fjlVEqRM6yonsugz64ZdPePkZC4J0hhy22UIqbcsKX41evYwzOv
KGrubGSO+oYN1fank+o0ZcWOtEQdUcie1T9vSqD0lBrZK0dIzTO7yQcbb1b9TqxFCGJVV1Gyfzs0
KurVlXzxFNglJ6l2pGjH+tI1kh4lbt9ksXPU4C0DDpdg4/EbQU7oZWnwZi7CU12HMUuwVmGfiNYm
6IgbHRmrHsSwnrDUIGJ6MedMJHqFh/Tt7NTOa1e3FiVu0BNAN7eZquF5t+62T+pPRZiic/5QGGpW
xPZjSi7veD88xIpYSV8VTJQ7ZbHTmDuk975zBo84AsZN1z69GrVebteAZBQ3Z3WDs08gO21OusL4
Jv/r4yVv8Kqt2JVP8M2tVqhRcf34dvZpHQu8FoUp9PEOecbxzNA4XfukhSXtprcWTOkbsoULlF40
YmIVM9vp9We2UrmL+TN/7ZRU818OQ2Li2QlC3M0NxuxqLSA+uVUoq2wxqv4CGad1VNtdr5r88r5b
GWyNjYeIlHYJiQSK2CxVsN1DRj5i8jR9WMDBBJOePmBZn8GFw7R9ZOdYdWj9cnN2bay2mEnjFUZI
QsLWzkICvjqeocEMPu3zwNtnuN4kZ9tBkm20CVwoZ24Q5F7PRXrd8q7QEQ69Y5xkBRMIGNozzpxy
IczIuUcQFb1yLGgJEOt0W1Hcc8FbfXe2vzg4kLle2ApIBvtmAQhD7Wfl402689u6gEG02Nnw3NrI
F2PcQB8GhgfuLWuxg7HG50hfjbJ0q1bdi9sEaG6WwZvwwZSNFSOCAZZQBA4+PcS/jb09sfNaqFw6
5SgW1chLVvqreNoZjlk7EqzHjnamCaOS8Iuk0yvw6E4PhjVEg4rdfjKOsvplJNhsIWYq75exld98
ZGdOns6Q9WNXfNirPpUT7tbrRrKnd8aE+ldYGjPjm+I7pLLayURYNmNrCksJf/LVTuTHYlDH/S5m
IOCPO3dItxxKtN6JEQDNzSErtjsnIVffm4MpaXmhiTyX4QMcegur8XHXC5vuhGiXXJlbtm7njKP3
K9UsdRqQI5LnFP5vSWB6RF764MrliayLZSRMVmtDe0CsbNiSFnN62Dc4cpUN/OWK0/UAWyA3ydp0
aa6C984c0doLPaPLiSu+IyKD08VU9o71GXyH+ZjQcOYBX6Depm4pEvpVRtJ7+5caoDaUFgxt8fvE
Xuwv62vIJLD25KaCisQZqVWi3ebM4cZeMzUrQiWI5wSLiXbaQ8glnHMwxvQS06v4itoi6GrA/INF
pIN+wERRbi17fZqm/ebn2ay/lBBLts4TFeCT7u34EzdhnOFFXg+eFUHjnlVmD45NXLTjt/PQdhYY
k30BwlQHygFHcOQkrpjrFfXs8FmdLJ/oZogNaek6C+kMX5Ee14NSv278xj+9vB1mNBk+Ed70ZNMe
P1FmWSZkZpmiEieZkkG9VNNNWh1+i0qUe2kQKW2Phrx/BeDqSGCwzvFnCAGbLzYKIbzVpYqqdVOZ
Tc64dATdWX+eDKc3uKA8u3WtIC6yx8MK/rI6haLTNuDQsIo7LhIZmdDMWaTQyQe/0RqQUlboLufL
HI9FtL5hJP13CUF2KbIiNdRLXIX1MgzmpXT20+kfl8FocV0PhEMYuToiQcgUJQCUR67E/yBNb7QC
alR1of3O8tSmOhZVnJVvIyVWCM5y8OouYmqlVoUvhTPD2TkHQm+zSuxnF0MWvVwEfg1qC9lOT0pg
SCqK8h+0VL7tLm0E4E+Ba1qmQDOrmUNaJY5vUPmlXt2ikYfBFuMwEQJxc8AxbkXSJ61g0+lJolw3
KhSYi0OfPMSOm6086vfxIaKfMZDJv+J9Le3bv8le00Q4oEaE3NhyBOHmzBU5VbN+b0dJswsJ7xxq
Jbi4LbdKm7XKhOJeP7l179G080Pn882rLIYNxpC2sj2hUbf7hMVER9xL+3/7k7qwdoKbofmt0CKX
/EM5X//7P2IlJcqph2TgfnROr3O8lAb0ezKhsMyEdGst98gntETt3GUkMPlhcM12cKHgsQVd3+3G
rYY1aedLeEDP1Em2kpM9roieWg/CBfb9sq9bNMNw6l1OyIVCVmJxsJYQwTZm4yrZ1C/Nj8D7x0Ha
9mcSd/yZlsp64OZeBWd0HEn0F0dSiYYp/57KDWhKmX9gFXFuRDM+Y98tQHMVbr3m+xvracvvSVJM
RE2nfP2xg4IO0GarJynY+lXG0/ijQtBkX/aj9HlmZ45HtvV4rKQrv+JHlZb8jOimezOXgOYcwMu4
3UOuxV5vlqiUc0Sp7gZ2h1SeEAZnYwfMlnaSnUfcMI51FEk1iIbn7AStpIe/HDHeNKPULdP9uvJi
dTgO0+gsN7AOoYEgVXPGZo9AHe7O5UvdpdwWDQAYQdu39zB/hkTMKayf0MmqmnuCP9Ch9LI9sNvc
CcxWqOwmQBkQM2UDvmS0o3ym/kJkbBMXSUSp1ElFXcj0S8nHfMX+WVOK5VjiRILorqiQzTeOwbqM
4p524LoU/hBA39xpI5aiTVEtYfZzOcwJgTJMXKuCpjAWrwTBOnh9irNWVJRpmi9ONv63fzhhuBl7
BjC2J6TXt5tj3oRUM2vezaqAt8PbUtMbxhG0ANY+9HUcSMD+wGjykKTVQOvNtI2n3py0+r7HePBG
xJvNQrG2AgVWOHk9Amkpyf7vGozlpvmfzQdlwxGEuAeodYLGoOoa8MlgKVYvsWwt7L5rjZWqOuEE
Wt9AOVS/PoslHbGHisH25eAlEN4PKO6b0zqTa+TgjYGVSlwVkikVFfFMp4+VVzIawuiQs3hhzwF4
zyQoavzmtnJyWlEEUeeM293qNCPNS668rC1HjR9P7Z/ot+VpGV466MVi1EPK+fGkeQuGMS0D0HGZ
jWhpgEP1AQCmCPn4Y3j0WXybqH0w4gYdyIhMEfqs8juQBh+rm1m0Kgw2a2S/KxKAZ3opKTa0j7Az
Y0cBfUpWZ6ErT/+cY5t7lSqTPL3L8HD4Lr6o1mCpN4Z8zhmnWH6raA8uDyBZhShO7n8P4Ui2zF1i
oVN5XlosDFRO2mZxMhyi4ckfpvnRStOGm653fE3b0a2omypSVI9IBZEBtgXx37DVu33efaiUsPKC
AWiQHn78gcKeDevijZdUFYbzwTYPFWn4rpPJmk4VmTlo5zvuRsiyNGXEwdCaqljwQrTCkttBwr3C
ugE/9YQ3AxsAS6z52kdS0FUuVae8u0e15OXxi8/A8he7EEjfHKDfjuX2U0OJCQuW7R82o5pekHjl
HkolEgYDiqwfJlIuAdzdvevZaih8JEnNV4wPib6tgaz4OkU+I8211P/4vhZfYhkXy0IgQBXyWntc
FmJ7AOq5KYew6Of/ffvJWh18WhaG1WtifRStqGIZja18bL9WiXY+CsHu7InUYP0xBRfaQoDkkKDR
6QilaR4uJQ90L4szhMkClHRrkMmLh+iU9vtg5T0o60jQZH1qKcVnY4e08MLU+liGmre5iSiURph8
r2nGrAOH7773VGzXn3miK6symSy8LeoAv75bIuIpW7KNAqB8sE0HEa0Jy+R8va7ki7Y+MdLDTsLW
5xUOhVLSz8D4g8lHzBMacs8w2jnNp47HVeZPa4GdJ0AIw/Sj5pNXIWHtxqjKc0sllasCFH/S1Epr
7FpbRxNGJd3nM8yDxTUdd2XF8faLgUE9z2tttgtQrbBOrpuZ8JnR5FV2ZVv8Z0c0pF/oJYbxVBpI
0tYyY8GXmhClkwkWlqX32jTbzBXdiMAZ/lZXfFlXxztsswur5LhL6hSvSOGhJfsnrM/x+cfTIpE4
qGvI1Vx5grIOV14vfUtH5hUBlTXc8RCieD+VDryk+mQD8UNRj8hkJzWMzgK7KE1CSBIIG0JOGEKa
O02ygyhsJZCTP7RPVycPW6rnOIwMmdvrB70jhsIVgElcLrjw2RJ75xqCqZ52cJ3Ot2yIGn4z8IiB
5HugnlriSsD6szl3H+wQQO+qy4jD6VDFtZO4hckI9EOsGZQ/HMuqgQATJnT+qi158HTAH0A06LTf
dLVBE1GwcPZ4NPlJJuxXGrEaANQVzj5a/wrdb9VyXxT2hLl/AmUfx8kaY97PP+32J+3PB5EUgABj
ObDMUpgGYD/8FDsoG6iJ5EwEM9SAsBNYvMmvuVS88EXUQWXoXltSl/X8fr6bb7RaLghF350Al51L
PzWy/TijX20DGn8/L7yO6mRaKfpTyx4impyLJCnmGZL/VsB1Sz7mPcDmzfq5ChV/l2lqwrFXaFC1
TK3JizHSGs0TuoPZlr6tdwPwB1Dkv8/5Tas85O+moReH6L06V3E+JSRM96pUsmscQDOB79EfdMYU
/KOLNRqzJBy3biWI5IWv2iDV6TlK5QFQFLs0wo1lfEoVimnLB8O9GH8lK5zgdTLt1PH8cSD+MHLd
VNxtAuKmZA4vhPkRijPryDZ/Cozc+ewxpBIxjQb6IFqwnhI9lc8Taqfw7V5/1vidhVVHs/dTHXRl
5tmTwLXkbflfuDTkjbF7Qh0dCQABmBpXfim2K1BY3EklX5QA+SmF8o+yFGgaJyPs83qKDGuU7pPO
ObbeORhBCqkUAj08EZ1Tv3UfKL/c1zlyYqbHMm99gtRhBG4nfK1GtzIn/cASFIZ/YlRVdbdSz6Fy
9686JpIEBMAqhndikhX51/rSDcu8JCtpfJD6Ps918JHFP7it2xZQeltuZCL6Ljjw/Q6GQgUrk1Ee
JF/UZbrrcTPN9yFRogUGOAQYZq7f5XDpkcL+WB9sbJm+DnWxTQqTAopULeoicsXLiYxqPFu+4FrE
ZP3riLACyDPrUX9Iv4zX9v9LtOwXq1/mlTieszCqJQ9pRqcxk3VmjUr5CDl2s78JoFg9M+jkILF7
PCMlyYxqr2noEG5q4tCOR9bCkvqoquYnNMFlBwI3RStfoKIQ2aJ0ClmQKQcC6FvDzIWktmOQjpPb
+N1OWUMhy4nE2QBt9IL9e3T9irCW7S1zzLZERdtPri6yRH3+pfCSTLib+St305dBC1C7iZ1b+QSk
6k78ho/sTqC5JrrjpAM+Rq56JLnCnGalNzJcuhi0lh8xypc8c7eec7/0e1wnWSXff+yhd5GOQ75T
y2i4uMnMrQwJb2T+aDeiERlXvBGcoN1q6tbuF53DJ4Hf6hRqrP5hzkjeqH1BufrrA7JicPQQNjkN
5EYxkDHAuvfflg9pwe3jgqCPeR7Z1fAUZi8lIqxiASMtyI9lYpEykh+X3wizMbJmQhkdzYnFDTCI
Tq9oGaJK+VO8GwBEFqTIpO7sn1XbfdIi3E0jamMulA/kErVJhaEACR0xHIApqoL6cyczBUbFixaz
7jiFvVY11TZEwV+sG4hqaOz32hzpAZ65KKHwexaHq7oQ2TPIIaPIfyuVLpBmcMPN+4pSreh3p9Ty
d3MeoKZrEWgkHnooZZ60kJMZ14woOdCebMFjLzK+8yzK6QwbJDagY7t6CnWFIoCKfHLVwqwWNDOP
BFoEGh9NtdDF2EexKJlvcRLYJTzHozUji8RBdSYg7ZIGNz53LXaF86QbhjXUehtFi2Pxtpp96SD4
YkFKxcRXoC+rMrbB1TSMD1tmp7H3oPYdQdHt9Pn70YRKeCmJtqG6Hom6tss72WifIf/Tp5TuWlCg
W9zJCyeXNs5rqbczENYW2/uei65W8SRayXhQ72OdoWof3iS5UIGrFcldpi4RGsYzNItyPakYHLvG
AJYx4xArRJTRD7JeObwmMTS0ztwqfZdKrquQ9x4AtZNajgNDOXZuUJFYcGHqu6lqPukHQvaBwURs
8T3iwtlthKbwyC2Cu0eR3J92dvwThR3Jm3BCz2EiipUuwvvXXY0ZZtBSoAmE0h1C/bBhjq8voRGZ
lVV+aVEZG2Mt3EQr9B3snQiz2eUfrYvw/EUq+Vh+aRkwtyeXZ4xs/jwLIPd9Nb1F9mU2+/ce0OF/
uJkiY6p02qatJFAxf5Bysms9V79a5mCwf2qxSbXt4tKMqkS7Xe3MPMfn1ngzz5fQsgRj9jR6D0R7
ih76CCYNq1NE64J8k6C4LTe7rgM2o3X0s2qlSkXfvhlXOkb/xMglUMRDJ70owAUlrxRmNlc2POki
dCGqDac7TNueyFcy8ErAZm7xeWmhU8m8bIEe82bkENH+A3RdVmfRzEtqz+pHuqKx7nvS13ii9yoo
LgxofVpqKFGz+Zl06pXUym/CvHVU5Vd1D+7NqHdzLrLR3uVwy9BHMQuOOq0g7W4BXgyMPH6kCZq3
WxjCI9ZjGFrzcNOXzSbh78guzazIzFQFwXsad1E/uAFXchm06lPcM0Z2hfVlhZ5EZSKFS2LZham0
a5ffQ4uqaX7Q4C1ouvNq2OO9nlzwX6ze3CjxFkvsFZb9I5P0dtu+wdx5DpAzgEEM7I3Aq/mJmObk
LNNScHcEx2eZAmQv/7veQvcSjko4Ru62wR4h9KIKhaHFzdPxA3o01gzPmKVGKbiTyLaMRUH5Csim
rIzzhsR2nuF3yDGX5CNv6zJ+/UkY+C/BwCRslpL72C8CwhccmvUmzwVlHIWaUb2da1RYbk+dA+qk
4uxBC6G+BFLrK1KWEOKYQRSCLwWQLFCT7SGQJjkg4pDI0KmCRSAlsVCZBm+Ij1XboHOwvjdmYmsA
SEXjzfBfypu+0qe21yxOXuDnDz6spFwiOThP/T80aw2qIRMvOma0Jisfvgvy7hDffvqNdTmypVSp
5HytGPCte3CN6LxQokR0+WCAd5VFZqjf7MprCx9Wsq4jwt9OqJySstmx10KkmG9+xCMQffZUxScp
JQRDhZ203qDmU8iLRxYrKD9iUmem7mthQvjhj7eJWriNWznbKgTd+KeoRyYMcpS9qEpGmQqm0Li1
Sitm9oXDUXWWOdblwsxKraDUVl2N17cFrRLlvZxZeFh9xMC975g9/1oIa4wzmBlGRC1aUkHr0JIS
Rwhvfeydbxd5Df4D7U1H+M0klk9cDvPEE9nSgQGQRRYTmYwvK54dKlra9EApQPLtR2ixzUIunbwx
Imlo4yLiAwPEfuq34Yg+ncyIggJ+kxzvksVRcpdu8mcZRc+O0h74YpSoacdmiNwioHlC88prAPpI
RMLZ/9K1HUsYkGIX6BfbGkPC+QZ3pCs5eU53pmDDw9kpFiilM9j4Lo5boPeEU55EprMWD85jvwiV
9XaZ88OHkAtZgcR51dOZkEhlbr60nVDLQLB2ZiDcdn9nJ2DfSeb05TPZKcjjz3QINgDJla9IzHJv
3WFhYXNykRIEzYAn0qCw+fj4VjxnAqKs9r8kZmdDN4TqUQ6snxupuatwo1R0XawSH2MapyksI79b
9Tw70EYypnkUeaQuFyADoCJZYsqYSVPwo0GWE7VYPcAH4JIuSmT2jJ2cV2st5OSe6B44J75B9RyC
SXsTNp1nBtuhpwqWVtI1ozk8oq8pBDgbCy4sQpCN4BeHCniR21TpaOV0QLuQUToHn5mRqDCpqmxQ
5uHeQLOVlll0K69PA7esH2rHF8y0PjIuio7/BZg0HgwMDRlDzXD5xawjmqKI1oEbfv5VQrgTTl1M
z9febdRZYW7rIZHf8O3ZlQsHA7uw9FO5EoxHHOy4A43BXEmGTJsZgB9kFHjpPChEt8yqYeheY9iZ
GkwCurWE989O2kvgpMJPLZ4ESV8/RcmOjPcVySxq8G7Vw71yci6DpXuk8SPzyQwkWCK3r0MxPUPo
adP4WRZuJ/ce8qyQgY39uqoJjAUIQx32k8A6W5yg0eMTlUG83RZFdy/ek3amjPvtkKuz5GKeix05
3eFGNfs1iCY9y+52CtJzVfxNAob+bqvxQG3iFJIYEATqxmuwOkEzhJv9x0efMXyYrlg0T7+H3PJB
qcHzsMQxQECskuodMSE67Y4N9F57CwqglmFgxT2zC6L+HObwhMjNXQARMVX0NuGHKcVjAt7G42Lt
oqvT6opqaZx1+XdqZ/+AajbgJ6Pk/qqZjz5jdZjTmXvGUCnVqhnj1jWSDMir7PduznkcQw17qr3x
9PdKSmWf6Oq4NllaayBPvP29IjK2wFtA5IEW11QNRDUxcz1/50RNnhdUYaIxyrScwLcE2LonYf1r
Jb0EPe5o15FSVEveKhkcEV5tJ7i9dK/Z/cpVhsd/9cjf/Wxb3eVpZCYbON1GtjNLtMCGQOdM2O5A
CV3NY9Ptldr51VByNeC7Qz77WX64vQgsh98ivWuG75lCqkt/OxIkTyUkWFxBAuj4EMTtSK8I/Jjj
Y3LEFwXeDVUxsaJyk9d3whQPpKywqpy8Q3lDDpuR911p9QFoWsMDdsI6z7YczWZCx8Sr6JHMn5gv
Ycjqv+1mpWvt9/Ro+x+8kNx+tQjK+kDkgB+vZheksmZ/rJazrjwtKAvzQHnz6vfEZSKV4R1lyaQw
KzJwpOlLWg8jSxV5LnrFJy/jhnhgNw6KgbvsKoNCm5S7/TgUB3QhWn/txBBlH1j0pawO69g1BOvu
EvyMNTbzqU57EINWKp8Uw7mEirAub3LEOr/ypngXBKfKKFV+xqyz31Tx7zFJrrxYTkmT88qg6xcP
SoxMqs+jvuiML9T0cY7oEzDhQPb5lJny6IWckcLdckng4aZk2bkh2pbGQMDFUONWAqgD2ASns47u
vfFvEictRSz3xyPezE6XtmprhvSYwNieNS+I6oXZUsyshSu6kkIH9o207SeV4DbZl0hQ/vRmtFjO
HJRUOk0i7o+PkWN6sv4/6p8pXCdG5Zv2RH4HGGv0xGkjOe6tf7CbqESNt+eyVwZLS9Ro8leBRTwX
h2PgRSVbh1ivMWmDoplHizLWWL48wGKD7PkIy60TxikHSoli/3dHPqa38KYgY8BvTVWO5UWE4zgE
e3cDRFpm/MMAePT6RKHPDUs2VYzg1l019Cm8uOzTjAABG+B1K+FyTBwuGK1WS2VRupcYLuCwfMKE
6OD2OL51qHN946TDzD3U3XzGp5bvw1yjoyukBMJIatsmjxvE9ETV8BjxLkF5dJNO946tMDcYclpi
2bQN8gCvS0fuAbFVDQuOXpSAXrjcSiUBrcTYX0RviBj2TT293JkwSfErLOKj+QFCJMB2a3qA6Zk2
0WJd6AJeWtJADmjG8iIgbDoFsAZLsXZyxkaF+xS2UcL+DjKp8ku0uGEIR2KQoeUKCc01+BZf082Z
komcPDhnnLdrpGyESCEfCFYMe1V6RvhlAxktp+Bvbw4mDcBOepnzPKyTh14ttsOVgUtSbhwUMzud
XT/W9KG16Z6n5D31FaWt3KvDGUcMlRI9ik1Gya5OmLYtivdXZX8oeIjeZ61/suhcL1DZouqiIOLq
V2rt57oVLfMTPfVqlxW7utkVs2hfrU0HK9y1Hm9QRAgybCq46X3eXFJrZmbUaDShjYjeiUhfbpjg
uoUQFKHjQW5R8u+CxJiWtAsk2wMI4ivVddRW083Hd235y0v2QrPuMI1SuNUQ0TpIfw58pTaHWsLa
jkPwA3TFplQzDQc2MeolXxDtHDR66pzVTmw6xQTEb0XM8LNd6i4V68ufDQ4/QJxiVaq2+32PW/nT
xkWhOeSwsOi+ezJxmBqwr6nKjqNwZhL5SexvtDTjz+4NofEmj7kfjxYhrqFCm1Jco+C1R536C3jK
mxcHvwic3CXI8SzqutDGI2WIhSVn8iMJiaKd7FVEBSTh/AU64nsxPRfJWrMhVe9MvLn39XTBeAFj
+JFq5ffHbk560ntgziMMF0jyXUVgoXCNh9LFY4Zce97MMsO8+oq0xCAN8hXQsLVGMteSPhuQX4zd
5TI6APEElqMOr6zbOkZTUteBLRuVF09htjBkenkZPJ3cKb61YMK0iGhY0/Gg4xgTLcWouMcJN2l5
trRh7V2lb3DkbexUID1AevAronT9O6bSLK6xTHzWRF6+tyAEHDyD0XmyNH/NoSUaOLAz7Xo5wMKh
f0Iiz7Vsa71Tv7o1F7IML8JVhrlPlicYdlet+PRowBlUg+FdmYasp9wAKb/o6tE5rCgqToxK91Rx
ew9P3XrZG2QvOoOtCCbs4NZJ4FMOlD4BHzpdavH8NFd+NUvcS4/5rOsHOYvecoaL28KkAZS+p7SO
qV/nlJ6zbHPUx7+4Q4Kd72AVIbuCIrhVT88MhY3NP4jmjkAqaOzVStHmXWoxFpSGure+bHPK15Z2
0WLfA+RxQraaasOnCtPDTHyGN7rig0JJ9feiGY8dI1OW4hfLwTFFQFalSxrmjsVtcgEaFnIopVvh
9ARk1RdZXF0VauPWxsP3ZHYtOTON1KCblulaS1JrE+DRAjLYdGUOc5S03K0s/s9jNfy2pYWZhu6/
P1+5wMaEYNa5VAybeIRU0045z1bxJJXwi7Nd0bkM957HBiYWbWQTK0HSfRxbNbuwWlZosLVrDTYi
q7dcTxmDsrdHub4yrj8S+Byku3UeNtMYzOLBMOwhiFjeFrW5IQ7gxoO5zqzzQ7W5ybdietZqON0B
Pnj4XbKbZBtIhZe1NeUWev8j/aYLiWXwYReF0HoUzbDG5PtbFmUJJIMfIZ5NpBBOGSyIyuXzPHbJ
hqxdDQ2RVs4BbuEB37r7QBce8yGOIlzoRNOEu3AGP1yN0fB+rKKbMD7VsdGMQfGDQUlVuzOucCqz
/ghtGMzv3+ivfJXjseY/fDxyVcFffMZG2f+y1HSfJee2b+rSa6bh8U49uGUOUoC4wP3XdP1VUYhs
CWA79z1T4kPkbIkBixaQLrry7Vin5f4XEXafl/tICIJR1jz7HKVucTqlMMYsJXk/1oY7h9JELhOv
nmgIqcAnhX67diSX5PP1WoLcRgYDh1OslpjbIP1W3/1cO0SjcMR/HuHSsg4NH5eSMNybsizmHyWr
E8+OcJCBaaNgqKa3MefEAulJBJZoaRU+1GMBWueINHDG/cVKzUvANyGR/WH4yK4ARNF0GyPXpyWP
PuAdWUfDre4bfRF/BfWe+Vk/N56CsND4v2QvFagAc01wRJLNDu4kIkXHdJx8IV5w7Bw/A7aiRfpu
TJKcKm4S9leNO41UCWWkrpYBjC+Ws8hYqVAVu3W6e0hNOoqY9pPa2CWv3j+k81rkDGkKD1RPXKRk
zRgJiTqP5vO/l20MRHHdJERj0Z1RUw41iZGa7QPg8b4s/2tLaAsl9Q1eB0N2Wwd8YLnnmbOiLarv
8DUixhC8wwki5zSXbgI7SEJX0ZPPaJSYERKgqwgOr4flypfMgRCaw3mxe9308J0MG8gUH9O8B1FL
43Gv0nvvEu7b4r1WmuirgmRzCD7mIaPNl95ZAHmDOtnMYWvYWNt8qCHeSyMbiEhd9vXJiuxBYvyP
n3fk020XoToR/P3gNSwcfNQWE/9ciY7ftKbWhya0awtA8WDpSW+HHEvLIHbDXEndd+P5YWke9wf5
muskhqKkGrdnSEREN6Dk3AdQErR+VO5+bEhxiR6DxmzPkYSv/QbHIfDCD1U0hEwpbnIZuL8QtQUx
n3cHO9zItXTxUGohsb6PKE2bGi7sDHjRpIj2nkDZGtDLqYEqztnpkTQcnnc9nU4xDFwipok3aDRy
1NTEL5Q66TWIA/UuTw5ZTnzDy95eY/CcmB5gBZj0mWoLmzP9KU28/cuClV/194jPBKlbgnOOx+0Q
kYB92bR1WDNHg/87+APi8O9DZgGp8LkpwKi9Jd6Fp0EnjNr+k9dNQD5XqpZA4b58W0iGqFYRb9Ln
Y7KMLoCreH51LBMAGCZ6CzB1Ln847XTNxnUfCkvCXNKftbYJVho+6vC0W6jXqTfT17o7yUXsn7Id
HJ6B3dObUB8tkfDcVe363vwkCI9HIzvnChnoGB2Rq8Ass7gy/oSJFiXZvobME5bKavRgR4uiqXff
w0Y1XuZOop72/VR2MG73MiLH2NKhkocrbfjD836OEWeXhAeSxq/Vrwibq4NJQrV0NEQjGLPaN0+J
kQwDh91PRow+L/TusDOO4DZiYfJA5loptf0TZNQrJ5k7LPBnslJWG4V+K9MWbRmYoRYgv2aQ2qk3
KqIhfe9ppQfTYMaE0IUHj9xPuvMp/Q+Q1SS7aUbP2J64eURKBquhoymqz/RyB9iMNdMwhiroKXmK
zYh3qFhJ9sHcou7hi9Hrn1KSmCKVEYdaueOScmLCZKjT9/af67mOqbPvD12YuA599V6F5GOhkIQE
uHc2kKGUq+NcRY1qQAJ/ncOM4D2Q6AYU0gnF8rPblBx89JpM75DwmscB7tBHoPXC0FQR0oNRNoCF
ky6pYIdAs1vxUFl+9zAZvJ+HCLR1LHyrdyywIsbjV3fR/n+FYYR6xYY6buBWcF7LY1HssBZCaaNO
qrddjObbK+wVl+EzIfViL+bW99j1d0/IamjwoSbN2tIO/TSkZ8K6pzdi/1bxw/XomTInScg44xg6
TlPcoYmhyXWuDyDxewoUi2KeHEFN27Mc3+v3AFayvcHQDHUTCe81MrBGmOa1an5lk/T024bc/p3Q
cgAALS0bg3AJCUHnCYJzoIp4qqeyBLdyT/eva1O6afAHDkeDyVARbiRDeZylti1AEChuFeKUNk/4
st2hZ/ybnN+PNwslbGV0jyB4baGEXJnbdqdncd11owtHO4XeQ5dYH2qYvRXTuNfUtBqelIhwL8zO
uBuEFKa42GOtHVQQNUSW1MdM1wKm7UxYyu28M2M6+wmHnBk7hyW28iu+bcJgBK5PutL5utQLnYDs
ntnqKMmqZ4pXhiyXa6rWXA3aKUqiDwloxv+Nz5Vla4VAfkQXTM6CE+f42WQVY3UcYo4ms9WVmX30
hezp8Xdqd1hRTX+RJmDoENONjSmVIpv6fwmyDuEQNGeP1DHRPtcyif8x1VooITbC1BtUgRWk/oPy
szEBcrZOIB4sHOq7xIChgt20qCrm308/SxLdE4SWbpWxw9CuwvSkw+9vPmBGJm6QehWvROhCFZPo
tAJAnWsPoWEXD1fQWXDQgsYfpFdStcbbAuvwFWbrNZsL6kfbkBvd9DmoJPQtRyWIBEWn7tKj4D+p
E2Q17KSgW3GIyZJm8C642+EXe+erW1DzdIVoqpI+cQzzIyw4YUQ8Vqfrt8/UF9WT8wgp26ptnzKE
zimRm6RIuYMvwTRafJB4LPnVCoiMfkDO2D1QRQwyC2o0DjoThxWbjCvvVCG2XxtIEz2KAX43mIzV
iCXaJXL/aIxvo/A0/Lu8bCN72naxaw1kM6vEn0e6V6B5RrrJaFgRHGfFzCba5dY5PiWm/zvtviGE
PLrvMrdt6qzMa9OaR8kbCQoSbEGZWdY51AG4YpSM9B22I/SChvzPVgDcgG2XkAJd4B4aQ8bxglTI
2QZA7M3Bj9a7CczQRSfy/gNjMbjgeBshMCaQcSLhxPkkWuXV0Kij35NoCPv2AFzfaoDhtPrwnxrQ
0nm2lgqtOHXsYL7qHa1nppuAIwgz7zRv5A0I4r9gny8zw3tLTiAR8vT7YXyMXSKwjddvJBlCnDhS
XQyD/CMHYA90hbQBIhZvZ/llIcdyT2ty2Cuil1Jcya50OEBTYAVh9okZplZ76C448nqBV1HGwO9S
+WZzVS0kh+9IjkDUHWGMwhkAaoGLy4N2gXg1GlINgUhgT0uCMbOZPJrEAY62ps9aq0YKhu4fBqzv
+I4mSVMElSxZh8eVnx53njw6Owyw8rksKisFVi40XaTfvOGV7j5gWEkFFgDnhNe0x+/H/wCE3Ua0
fc3gMZPc8bnkZVgVVH8wYHrsY+RXZUxCtolSpi0X19DLCR+X8HF09AUtApCNuhfkCuWOocKIVOKX
7LYvePEnsqJYBk9633UsusoZU6yGpXdlW4a8Zuk6bpqxvnXOI4JVLffFqrBRsMop2i7aJY31W1DU
j3OaNmFXk1bG1MRYtRO+MHmdTqkjhsyZ6IzHNXvSGYWrpDahr2u2KZtgWyf5NBvSW4AzGkbgIIC7
CkekDQmLS3Y7wdbBbBDC1+Nzyo8zzW/ID41fnOfJsyBWaIQLy73XyPQ47atzmjvAthOGqVU5X5LV
CB3hOtuog7ay6OIVcvRuwt1yPHbIdac+u7o2efj2wSi3w/0ZNBU4GQAEA8tD+K0Ea1KCfeJepTR6
G1ggmXNWF7IQ+cQ/efSGaYvbJchIm7TtN1/UuZaoYLpACsAWi79MqDwBADxtLkAHndAnjfiHesP5
xvc/6skphtKVZTcyktDAjPEPHT+haY1GfpdWzkav6YbNmsiejGbGblHXf0bgcX+pQomtgAjdOb9J
iGZGZ0DxPNuiFEpW4JipHyGwDOPMnhKDLVByAbr3m7BhTrBDfhRcKPU/4Nr0Db1Z5p6CGsBDSBjB
rLbhvXWsBsrtkggZGjG0VCmrKJ+kkQT+F/EEMFXCca7KylMm9QgL6rN7VgxIfRS8kmL/v5tYsvXO
XiZzkG5vzbS0F99s26UXqUcLJ9MBVwj9QzyUL3o521y+q2h233EMX1q066CgoEMS/Y6gfDoSDbGe
wJUPGQh7yXU68/k9/XkS+RLJXoN83VtK8dnwLWFBlNKgQfbqT1G+pFN1gHQ8pX5cN3GbwhJgPLEx
37otRTut4m4eAIQ8K2JVRSE+oUPHoCJRc4M7EvV63J1P689+m641gIR6aUqLXW/ng0VkixC4S9/2
G9DaDnxDTtdwkS2nXGvKyK29CS8xFiniTL7J9KEsqwcXkqVdLF/bnasbC78aJZsd570z8dct+0eA
hx8QSJqIZn9ercLCrRVBMTZfwMPp/1Eq8zvxB8IQctvFwicAllNDWHEIe2ILmPCDAFWp3t+2ZyG1
2vuprS57KUi0LuCvQ1ySdeyVAN5e4Lztn94JS+cQDk8LtaCB3Y8gboi3jgXwRjUNzyQC7+vlPVUv
eybOXxC3IiQpa8JejrL29HsCNrQpyNC+zk8gONWc0sOijj3MtaJPFnqNlqHQAHkX/4HlPnPd2Ayx
D6PGkGulB592/sn81WgoM1AU0RGhNkRFWqnvC+sCcRx6T0VbhN+kPA2ByA9iBdQL7mHZrc1jZytu
lrMWdpXyXHnyVYbs/ZN5BivYDMidyPz1lR5adC3X1n4YcTSdl1cRCOvqcEMwndP7lbx1NhoR3j9B
dRE2e8wBnVZZsTCr/2LMNOiK4OFEdxuUQ7puPcHN2teP+fCNhkUf0YYudTl7w7/Y5vR63VDE8GXW
nriRhKYpwZR1yeaJVr4Bu9JCyXCvFRrEyAGQcuGNxzwFuX0/gwb1aPT/uTxi55sFfMBZMYGW8KO5
6GSBkBRU35H7x2/BRIkQ+4zgLsoAsILnGsc71eotcd6Nl0zLK74xUlAxiKHMvgv8+cmPTmiEFjLg
pYQSvchTAV0pG/KC71y17BbJ+Huaea4L/a9IupKQ9xEiI27qWdQR/ZfOmr5Seiym9wdKMlitQ4rg
exxOKQ8PiWyc2D+I5D3eBrU1d/acew2XfBPO0NhV8iXcWLunM1eWuficUNj4lR3x41jXMTnSgZWz
T3mMKNrBG9c74+N/sB6UG/vHBnw6ikE5Puwfd1b1a4ubM0P7QDM8M91bGY5/Gs7g65DrpKM4c1oG
/Z7L9b3ZYmNuNn08O5a+6Vu166VX+Z/4eYflV502bubT/xIpnGBekWdlEiVFyZViaoyVOSg22d98
0tES4AAZ4zpid3kl1VOI6Hne9FiFiuei9v6oWf6sxLmir4NaBzs0ieF1akxsy9p5kibcmSBz4wlp
i9JCqd2qig3bmwZEKpUbjBL1FVBnJU543VgAPwUdZYpnyNeq25aTVaDP2dNkSdEl8iC+DnUi5lV1
Q4eqQQRmRO4Zm/eFKHxwcKDbRMRRA67poOFmQqaauP3cwgS6KZtlJ/rujyVqk91V5Q4s11lZh8+f
E/vGuymSgFOpKtL4bm3t7MB2GHhE2WYdSvE7epx2PsCtdpemjSrBmbVB9S0I5E0P2vczsq7olOn+
P39Cq35VCo94fwYdVrQZ2eQ3z/OGAS7ao0GQtYagm8z6Bgece4i3lvJailNfIm2CWAK08Fl3Wj2b
gNPFEaQsKmpYRhdinKkOfF55LaSNIAEby6OChoH/UfV05NeA9i6TSK3FbnHDAbkaGrOFh92HX803
juFQ+x5Aw667wkPmnYb8aafw9+s9pORxFk7o1QuFxfmKTFqZyY1txBSnA+YXcnRusR+5ORPdhvcf
W96ewsuh/oANm9xU7mj1mpCqpr6Puy5bitclMLJ9USO4BSvQHjKytXOeDRI0TahmkviuN+HbAeAa
AGyJS4HnO+eYJ4UCBmaI0sot/s3AHSiO1tzfmyWeYX8onNVsckEZJ4B6/Tk6RxXZB7+dpOIOs2Lc
5kD8+fTHRnkQx0wp2zRANWCbdHjx+oZBAQaxgxTBuz4MsO17ovi0bain8REagI/91CA6J3PXSqwG
H4EDtVB5bxccklj11XA8D6yH3eGCtpDSYA9pJuEAuh1kCtR/jmWML04WZKQ9JXGcqwjOPHMBEUBk
h8nIwLGbEOmMq1qpT8lf4ztsUt0UXvkV3tBrQbMpp/k5IXj5jJ8y4FhlMj+OcyvLLo63yY5Z5P6Z
BD538kYXgVRnv0MzO3Eqcm9RWPEPQ6R9s6gYAF7N5LuxCqOub9n1rs9yhxGUd4OjVOfnyX8Yv1kO
D7KpixgPF/lChuCu11cFcllHBAb5JbHFNJuN2OUbjiS9M/Tx8fypomsnElPtI9gaoaIMe3goZP8s
UP6dp7sFFgttj/kYz10i/Sw6ASoVwDXK1OKRsYI1PjlzuFenK+ZLNlrZhFVC6tHNZcjdGbNFsOp5
0lWXwMxAptW76gtS1r14KfZOjp3D0aJ8JGRHzlGm/tiHbv+fe2iOcAlfXxK4MbFUSTadv+mSjmj0
OEHIyH0cY0lnCXwSvnkmG3SFh+ZuKOdNhs2ju1IsCmzSB2D8O/S9i2Wx5j0E/ioXxLVG1qsEa9g+
1rNOPajGS3yaVCTmhJ+b0ltn9kiBO+9PtouTg418MRcZ+tWSTXFQCZyPLcgIqPt3qM5VHMqgYKdG
4VKLwGXfbkINI3vqavUf8nEuotJX8OdEB46LJvaLAk42mrkZ2DBP+Kft6Y5v32e00ioo3mNZVcIL
QA//S9x9VEtHpMVZiCprHTinK2hk4voHGpqbdsws5MqM/0DwVQJu85+D9lGOCxU8UXxc54hDm0SI
3f7eqQC59ONNkUcqJYB37BiPEwg1jl/W840yIu5bx92nT8fzA9KHmYG6JfHSq2MUmWy3z69Si9zM
gK53Lb+YIKtT4+BVk7OCOmsPJC5o2YcgW9DPHAsbG8eNjxnwc4RGiOfJT14mgV8UrmCwpl8WcePl
D7RF3R8T53PpRebDb0qWAos6eEF9gifjs+sOJGIG2OS8TDR4dyMo2Wxr291QQJXorfB80mJiCZ6a
rC94ZwXDMWseB3ulJkmgLOW7aCaFQOImeZR9tgFmV16FY125BEx5RA9QLcOkLXbPbNan2EMnKrJ+
ova6XJnCeKJTyzUMZC3jWGZU9KUWvfvDrVWbJe6uKPC9ZoB3Dg+kvKbg9KxRP+XUv7TONJJ9CaHh
ONu6WZjgWqRgonzs7EGBe7/hlIAu8aQfvW7qQdAIDHsEXQjK6ORX7V/Fy5Mf0+khGpq/Exu9e+FV
DF66pCRl7/8Ehs4y5jqWzWm1kuVo5/oAsFDK0col0VQyc1/l7c4SSwMLL8PC6UGoc22n2DQG2y/p
/tOLa4FdtRXDUrnA9227KYYipscTKT/ffm5fCSCn+R1srgYFPBehFDXp67iK9yqH7wlpVhkEPO7Y
ap6CNevfeCXvGY9hdqAaHRWr/QgxbSYXz7l/KiqflaW09TSxymyfCFprjbiaNUuenbnjiyBi+o/6
m2v/z656d8pYRDAZL8eBS1p4SNu4xRYip6R/1Wgp1K7MIgNlD2YWZo6fCNQ4NuagXJEh83Mp6hO6
F86XIN1xoTrWOjQuK2dG+QA7DNEjosJ1Olmhfuc1KJ6joGMnp96vkQOL5UWt8/SAG8wRWhU8rFrm
5+JW6Q0fmK6BDOzKouIpZ6YoWNeU3GWIBp3zYgSqe0ixQrzDOWTWMHf6UrWTz82E5YnB+tTgkhU2
DiZKjNZX0NsBWpJEa6pZxX8b1sizBgbN4Wm0b6BHJErLU5LwF7pADh1htzIzgVrujfkQPkr7KIdw
XF4KHbCjgK6/pNb+caF8Bc+Y7fPDdw1Yral88hSr8otRX0rhjaNmqhcpSsRb1YpxTYXs4ijIIA45
nB1BGk8xxL694LsxxiAE493HY7dyHlh3DJGYY2HDQQ5pp1n8hH45eyaOJBj3uCzzM9I6VAE8PuY5
j0tUX9EnrXBxkE9KwUzGa/ZTPW2bc+HqULpTd/9k610RljZ9VnWd/qUMEErcU+f6OrAyXXhrxZVu
AwzaILM+xSyATFOGG1+9v++k5292N3oe3r/70W76MXz4y+2rkrNLAszKZTNwvlPTqfAQ1a5+IdkH
TgK+yx0r5n/rwgFIisKpwchv2v9GGFFuhHHJELqV3CvIpLNqbgDbxiZflY0Wq01bxip1cxaX5dJt
gMtO0QAtAPMPByslYIxYLOFqdOhexm08WpQvFSR+TLLe2MwpcFRxqI3u7bdrlNtxGZgpWqNmUrN0
uOeIGIfOhNscfP94vZCcrVdl8LZTxQ9B2Uy2kTr47OTr+7oXyv77PI9QqPzOxvAbLy86d5ViVWNE
fdDVAY3dtvA1lMpfzXNoieBCaK8ETzG/Wt5n7VFPrXhIKxtO1lbf7dT9Tz+QEP8Wqki8dHTsJ1+W
UVnHEP+6xPrLVBnXia0ek2BNBYX/gtecU4aBC02vRkQ6lIZOguHyqoXOvULrIEV+9X8HKyHIdx7x
a3Jo4yUmDwOoJpxOAohGa8ZPFwPrnvUMWpuJXquYcK4UmcG7LRTB1GUA7yVGfUWi9vHGWTudSUnQ
V+5CgFuNScS7GFcIsodIIgMWFxUR0av+TtlSxKzXOYxTf/IWJTcMfhzak+u2Uo9XAzWQlfw7Kl+z
77PcZjP7ht1W6MuaWTjiV87lcS2O5nfmc6wwpbjpL+W+dmOYqRKqvewK9b94sLXb6zAwCjKYk3hu
6KzmgDEKnekmPTEPaPStTIimA+HpQkmVKBxl8FQ/tnpQUq9F3QlVNHyT4N8OwGifsCRCI8AeIL7x
mF2MJzMIxk+pthdKJQTkYcCpKauAlTh/8y4stwmBUlYAQ7Lk+N52NTXVuir43KR2xaJVKI/svaao
sFb5j++GKCfzNNK17uVrEJK9wKYdr7Ni3L6lQbR/WywqjYyPBgjT7mmFXCVxm3+QPoes4D7OG0Ih
OKviA0ws2X2Fe3Rq/qbeClcvLHd130Hf5mJty15mk3svaJaNWAmv5IOCxnoyCAeHGLsXZcHKENjd
0zzzc4me+NapDCfKqm44/6hYHS03ykNdLzXYgO6gwDoWGXVPkcMGz/t/YmHnvqN/i/CwW+pUdbi2
cReAQHIgLmkOYOF3k6xmKdR/ueh8gbRm9QpwPPxpNX+uZwf50wvm/elPCRkjwB1SltY1IOxFWTLP
Qud51qk+7vTpvsRD5Qwf+xtbVYFm3IPBlYxGBXlUdfcXSuaadR+s6uiih6vcDQXU1H2JxzMER4uL
dccY4Nkuavb44itF/rN5BXr4r4PDGSY3rzNC3gXNick1mzMZ1qbBpiAytseKVXAoW8tkr6wRWaKk
xwaRt9PgRYlLWVJyZDL/dNy153EvH8M7YcObMrdNMcZ1vqRroo0f866q2FTRQR8e/8lpKQRQGd83
IeRFnszfAlphy4dbVo45Lr3uDUQvqlsOP8NMS++5H6uK3mE8gphUHrh162QbePKVh9GQk0G0YFY6
Io/599hIH2sufX2UvNqWZ1Ggp2Wqj/dOsznKLmC0CjRxola8vhnu6H/6MBeSFaetxPNROmzKyLfe
RJ/NqxHl/pAgtGl4zjyC/NJcxtvgUeBYxWYNqo0vWtLbwuea+B7lbPxYurqLHun3lCKlkPxC+Oaq
PcJ5eWXQUjZqc8n2ZhZd9uL8bPfvjzyG6HX7Y5bNtvPkiEs90Li1jX7YVFloHXsH69of7dNSjayu
aBb7WFdMk57KMAh9a6Xp8sT2J8dKweubmfD32z9iw3guMEbKQgzYxs5Hb89SYZw39HkPxloUUWzc
GWlzqYgOMqOPmFNNGPb0AVrGn7fy+GB5oK/WcgkB/407ic5J8ECiDndmsIOfDlxppjcX9VhYsgXi
wkXeEu424+EYEjBk8964t6rvUyuQjC94m5EGgBzvva2fWAF8gofGzDU+QTeefFoQKRae7/+jfMaZ
hwMZPhBQvczqAyfNX5iqkLNthEjJntk8DW1XROGW2BVLnYODrHGn/z1lih/yrHDnTL8ZSL/Mcwzd
cWVIboGXBKPE4knTJ/c7jttHxR5wvxSfByou5LG2SlRuBKT/XTD+LWwrmCCaf6ZD8MDskQpRseHX
zO90IcbnzXfiX09yroQw4E+zctgEIXJQDLhv2c8Kc40Pms9m3pZXiGHXwvVU293zoSr8+hjL/L9X
UTgmjGgUkVrnM573HPvfsklEe0piNcGPfQ6FmxjsNLdG3TiimpEQfaN2WBeXPUAN/U8zaJZ/WuhO
6Xouz68iFFO7aUyNdpXUUUiYdJiZ+8yZQBF4I2WPLJZyI+TTRDwsv20p/Dv+ohckMh4//i7U8e3k
MJhTA4734TcvM4v/yJ0X4zPo0UurS9/YIki/rT2Bjpa6bKfer+qAfL9WGFZPiLhEAoICJLNagie8
JMJHKmI39Yz99Jy3FqYPOqP6HYPQxGVquySaFIunikES1ZGeq1i3+udFoepUKN2KY+fiHKQBRzRk
LGWxY0ZLvt4v1A85Rbbd6i/RdokOWJ7TeawCkZOtzRiACYeSOG3A/mIBCOGDWPBBknKQqO0/foCy
dp+NoL5sCPalBa5yd1tEXo4S+DFA/3bD6NokQxDQ5NZAKzSxKbmSnE7DplqY3Wkux3iNnTRfFc+z
/TfZk4wJpmWlI+zwU+hM+HktJlHinwHFrpiS8y7eOxxrXnrjtyHRy6oHuY4uI/x7uB4lmvkYmAcU
/obDGd84J9xHQ21m5nZXyNQOqDj8qrTfsk6rxXRAxSP/Ucqa58iOsDJ7tleFDAxrQ3nAtnzD0u4D
YGoIpDwKSQmQErNbaP0dxa5AETHjU7no5vWCusxkoPKniHDB5tmUmtZTWysbmq6iAgDuBo74XF9f
ggnQAgFIs89Aa5Gvj0FCHvSsGe8/ozUwyNATFg9mqu/CHduv6UFQYgEcavevws2qLcqVqmyhcAZB
oEMopO2V/Y2hgaxe8kwDGbrug7CO/Iorzk0V4xX+S6ZloCkNqBkAsKEyyPAbY1ZnunFfAV6grQYS
c3GwrFWERwQKAeH7hi/7QbVEoqRVEkRlDeNlhYZgboagN590Y8sxFZsSyAQCFiLJ8gm5mkUJ8qeZ
onDLy4Y1V3gQu2a605BoWqDSx63JdFg7sQJ1UtLTk6SlTEWqjUamqyOl/rFTow/VsXcmX96Gs2Wa
FiJbsHazVL/U4CdST3iljGH+3zNhLSW2qgvw7+dP3et+PmOalpXtCcsumkF8auz/gMQ868PdIgjH
7VU6mVLk1YskDuC4+Z3qWmcUkGlO3vLfZ4SU+O2ddQmO+aCfZWMpulr6G9dgGTIbmEv71Y0ytr5S
MgVzOeHdmwnfhhQHJXArf5a0m4bXv5EY2R6fN5fT6Zj3UMbAEkzd1w73k3xQheR19oTTFrFsXlXQ
NxjI2sgFMsBXoxJmsFknJWGY6n3FmUG8H6sfQ/TLJwHatyfBxpnb/Ew+TaMUl+tg8UZmp292hhtm
WQbRh5XJDJ3wrU9VcrXC+E1/M2unPxblUVImXeYbRn0iuIu7y79muAyJoi/kmR2+GpnyUNEdN0AL
yHf4oC8LpmwSt4euMjBvn7qMiOsjrbML2Vw2K0lFsBqsXeiS3u/KAgkIXaVn/x+hBVTACtuBO680
KLuUvMfZPJUhh4d+Szw8zpDmtigegNgKVdCUoYGOirH+iUGk/xcPyah4nSjQkW/odkEiURGMdZMT
eQ6dAHRhYmBbHUHpA1m+PCW87DevSbPtZY1pr0iVAEESsMPJVuvvaUr/+5omP14DQwFJTa65sF9H
AMgIA1c3kNBSErp/JyBk1uXsS8tgeMdW4fNgjrRLKSjZ1HDtfSLPQoLVrI0dtsL9Zas5/ani9VfQ
Biil+0An5uShu/6engR7za8Ut18IyRAwg8cK89mqcROiGTWdxGZAbztpR4xGf1ygAvMVZUPu4XXw
Mf3OzQ5C2gfgn/meHKkk5CPcgjuxdB73gJcwLmEQ3aIs0bXLU5vyDVDUmZ2zvrjs151pcrf9MZOl
QViqL6GHgOc6j+CBjARdgLowfCVXY9MZFP3tbkkQOVhNQETcrEK5JlAhg1R9D//yEhxpl/CRc6yb
nJr7GUK2PvIZqQy9bOhOTf+Wmo8Inns7vmb6T2k2cHEWZwm30rU3s3eU/UGM4HObqT0/+ycIkr7O
Ny88MncSNyP5kcYqLEmfu+Nsh1gdDXNVykm4jnVvhL+yHwkNiQ+AEHQcpDjhGmgIYgpxkxwwaHON
3mJ6MWQfGic5zbbks0vDvmMRdY2CiHuCu2Kyp1dc1VjrwgdXWjGCukTEGov5IypmngFzwwRwYlEv
4MUl+cwTzdwTqAjin7KDnaDzrQhNB0oo8u1ab9d+ITZo8Sl5KovdAVmmw8+oRAr3fbj+Vzkcx3P8
f/tINHGtxqZCKBb2fNLddRKPyrBAegDizFgdwzx8euy9viV+HkSK0R8IwUUROAsQliNAzfnemlpq
ijowaetTlMe7HTNXgQWrOYBO1Mk/cs1kJvcPYZkhlK8y5+YG2hsJToaKg5nCL5GYRzqzF0R14jJJ
m1sIYzaXwGJ/F36FMzJ8oACcneBOKpI7iSwmbhF2F5o0bp540e8shJpLagLK+kcZD+HV1TxJyORO
AAYkJp6APmfyxaIrvUMwr2sxbJ0P+FID9L/YBITm4FhrJ/NZ5ZfwNMR5KGVvAFAlPxryTEGGTOoQ
zYFWhTcRyrgkcXY6XVO7IKl4Q333Jznf9nsuxKw4Ba3zefEq0M6X5/H2GkFmgGbgDUTZ6hi9nIPv
1aRmUHc4GIQyu7U6JuTbOF+gZ1HJfmoOFh/BhQi+AxT3fwoJ+xTYIciEaGvSIMNLFgek9u4rSz+e
4rpVPPBSmLQwW4JuKDOgDYdU/wa2g1dmwJZ6wP7kBguE7LZExesp/EaT2fYUvToZNh+6TuLiCKiI
Y0LBKxHf7LHgt/8NxY8tqvEXXYS81LXG/9zwwsEvRnij0dw/SzP8+Ll3XRsKNbdpc9XuyY2EWekM
7lrAbAIkjaaXOj/D62Gz9473wOmB0X4n18/tv8GpJb4eI1HTBMrf6CdIwo7KSRt77nZgJ8dx0F66
xNlQ/rtbAExVvj25VgmVWu4ezdLgD/tkeuMRZWA7lbo5TkBvGnVHW/sl3kODsPFwOvBKhG/lJK94
6VrMo4pkM9Z3JuVkHR95OMg1eKJjXTcmzoLpkIrxgIUYJ58WBYZ7K30jUWnipg5gCf2W56jD53fW
d8YwGDDQ6qSacjR0e+uRKOMD1GYpqt5jFmz8fUgSmD20KSQ0LuKUkvsEQTX3upFvu7LjhLicSEdn
Exh/RbUu8h/4ZbnNlTTeGKIdAt8+ynhcRrPESwhuw6l5eacB6pj8EkJTHepsn2PiFGA4tDz7PPu7
sPpFqQaCIPirarG/Gmj0DfLJCE7Tp3GqQjhPGQ/rxh6j+Hngmegy1HQJnmoV8FJbb2589diYUfEn
0Vn+8oyB1RA9LiTBTxX+s2H0+H1yXzYB1DRR6cmiZn9rpP1gFkKsKtLE1Sh2vfh7Tjb9PvbhRE7L
mtYwegwh0poI5qsrnT5nOiXqsuvUMaDCdzQekUzsD+80MFvPnl0epEnA4s/myxEy9yE+aprwFPqW
Ko9WqOSkL55taqIqCIThBLlaUQWSm1sX13wIhr1G0Xq9Qr+5ItnQewrW9Sq4qZ8z2NQDUryQUUPt
FZJMMSuNkYPTH+6YUJr5US/0jXm5Rc709t+mU96me1k55lXTUMrW+eOu54sFNP2nqJGakgsTMspk
YF2j09tuiqmXYJY1poPqle6mgW2EOm0qIavOO8c5z3nWz6zq+I7vmhb1MMOgReobgyZIi3RaHb6i
SEwz8qq2X8mjxmBFZtZBCYrLSMM4nAbI1BGSiAeeXBNcDEfYWy0Lk/NBnW3hn8paMTy36HuOjbmK
DAOF0OgTkoLQUndyM4m63DnA6bwrjYd+KgCQCyonWg4o2RzKZdJAJ36a/ojXtQahOuzdBtXO2pOR
Siw/vfoa04aKirNHrDbH+7YrEYqJZgZX0DDsrGV+WxRkvXh67sS6HPUmExG20f0U3e+4CzVgxnWa
BpFjKOb3H8lRtnKCeXZ68Qyt5S8l5uFbxRM/F3WDCmNWjVVRWRyy1dkQOzxbP+fC/b14aALmDpQ6
A/n4HQXeNuV+MsGrw3Aly/DfwvQYorm1vPuQOMbyO8htAMAx9mqOG4ksEPpty+yXZas+Oqg9fxga
h9cm/PYK3EAL2A3pYROnD/k3wtMnqSSp5h1ly56+N+MWKG2nKhvuUmt0ucVDpW/2k6t+sRF0ovT3
3ya0z5bPeiIrBvRnCDWEofHOD+DGEceC7mvCpkRFpJhTST5e0Ty84M3nVBGv/ZwBlg/GCBC6W/uV
p7Fv5KfZNs9GFtDw1JGIlzzwRs/PY/Ro+Z/F7ISI/xnbRMPHOzlJTbi368Y3MjaGYPe8QucbCx4D
yITPiVBKx8MpSZY1Q7tGQ7Ctnn+Ma3Pj4iaXeJqgw4H/bz+E/064ubNwyTajFjZYmfekb+MY8gTA
SuDryx4Q0m7Zfm4S7MXq0wEWl6OpPsMzfdEXO6vplYz8zHHT8AWAECMF4iZLKnC6uYS+rE9hkFZh
RsK7GD+phhNOmvLqUoL+uMG7s9ZOAtOrzblGWTE+/Tl2b91AS0XspKtmpv1pF2cSBc7MKQsK4AAU
P1CeZbUJ3ogJ/apDMdTWtOD1Dg/oU/D4GdgyQuEsGeNCyLQN5XZ0nk+2VpgaUv7TBiWDn6yCHAiB
wjovTuUM5eNpnixw6mBV846py2pgB3AbQIuLF9Oofp85E/+8/N1DPdcrADPYpMGaVcUBd1ZgPf9W
RrZp74L898DrXtOUGALJuRsD33utpe5/ws0ukO4ST9CazB3GxJEvFoVT5uZfgtdCcRS3t9g+kz0w
qIlr4ld8rcqJ1U0/BMRP5Z3hpiNymFqnE92qHiuCrokdrxT/fm7W5gy+diKqmjWpTpmwkfJx4nGE
hNK9smDEWSdwfIPOyJ5J7PfAE2fRbD5ceBUoCDTixGsAvvXXwmWO/UrbpsGsM1lCTnJr4RAY3n15
K7h//rcrtQQlhWNljm+zMcLoQ3J3NojaLe+KGoDtB7qC+U2Jq3wy+cUqEmVv/qtQ8LJHjBcRmgIL
puVhVG7UC2bMEUB9g2gjeZN8TxylE2fPuf5WX4XeWMfLm9FZvMMuODpchCHPMRYR1WH5skEp/D7N
WNS5Cc5s+lqGmhFtSdCYRj4e39uatlKXq37CUAaVXmwwXCwIHBaq7/GQOFdcWyXrK/DcpbNt0yYD
IP8dLfvKLl9d8hui++nfg2OfabXsbmnkxmetCJDIaHZ2uW4QvJXiD1cSWYzTE+1xFH6CwJwMt3Nc
qxtoOp68ofnf8XB+eU/4u7r5MgAWRLRLAcrAcAvQiHb71xkOn+4DRn+M6OXwKh4Br1wzdYk80gdu
PR4u8u0cdGLzuplGaAdhkMvVC48wegEl5pk+OWe2AAg2KcMdbDd2LosxE89IEAZs+XiqX7YGNNzK
ABFBPAFhwKHw9PQXxgGdmDY3WNCJas2rWBdpVS/TRTWABSFgy3quQIuBPnXgDH4bn1AdPaSEEtiI
/2TML6P/HxfXJ3mOct94iTdCg3z9z0RRtMz2CfQoXShr36PxuTTN8f41HRqUkMoU7ZNYY0jXdWRS
721Nud8Xg8kuKh/oyRETuX/aNN1i0e0iiFmojOEHqiTjy6LV2lFDxn75bysC8WMdgbDKDR5QviW4
Zg2bhBDtmzwXdMJTQOhikQzSovAAds+H5qLgl2mR6Raey1QMGoiNe1rbFd25vlFuwI8yWcnHN/uW
uAngTRNnyOimMp/TUEWycOuUMYsiOdSWeeI7Ai0OyPrCYt2PlsnBkK6kJWm6v9spX2KllLV3DNvH
iImr7OK+tA6TEF2tkm/AP/JLV8OX7e9C1xHXmvjWikiy7Tl6H3gkUOwJhJyO+9+uo8a8tebWIwsY
IOQyHH/AzbLryC6uV7M81NrI1kL4PK/X2gnUIQW+Re7duWBm1w0NDbHn3vOCUIWEfcTR8YP4JWSv
r9mnzu5g+kX7AHpulqSSvmEhVl5kMNMWN5mH/D5qrvhuZEgfkr9NvvgsbgKHP7aczp76qjjZs7q0
F+CaTc1SmKaFJvnnygBIcgmQr1J1t1rgP3t9e1QdScfztr/U4QAHBrD5NPZeDPWdqKRXS68LaPzw
vAXhmfGfp5PeuZwvRR5m+M/KMSp5Ndwv2Xt2pawP6htdLAKmGnQVzbNOY4GIBLCVPIk4TOJeR/Lg
CuFB3jBFNhDC1kWIUupDhUmgYOMNSd/iV+gGROimAdZwJiDPZSiJmkR04kJAGTxbgGB5WBbY3fEY
vbuaVOkxZiddnqi/fHdL4xS9APOaTqzwif/WfVqF5JkXXVqRNISpe6/DWyK4kZyJ12TqWa1YBQOa
Ca3UeMkNBrpIaPU6BXq5Px+33gw1cVgeVLMDnx1fTozOUdx+grQ55JIQHIs8btWZgHjStRUfpWRP
kSKiXZh4jBuZQX+vecuTHTxMezzqs3OJTPvzAjh86qmjKsImYpLYdE7W5X+KJ2Cfvt2LyvYXXgbr
xuuSYd9+X7XrNdNRdrhCBNUf2uJmuB5eE6nS2YK7i1JubJONTJtwOAjmlE6dw3J9UPQf/F1AHsSd
5v1I4dq1MnKxT3GJkTfGqs3vgrNsO8S6yG8EX2AREXCU+HVMmszzd/OXak5HiGvyKmaJdIK3EXcV
z1By/QTwln45m+lyeKAcwpYW/myf69qohNwc8jaAI/pGmNcykakf7yRBd/krl1HnT47NFpmUeITy
VNBF+NTF4EmeH5XRnDGdeSbAB95us7W4e12trY6Pfq3DTYhXxY2ic2lSCJtyQA+1IIRWW/Idr+ay
f5wpo5VmVVikK4rut4oecDgFMXKvq0dNzqJbvQ33RF6lflNdBRuLhXwijt1Wxra+6xgRHg9SAOF8
pLHXW1uizxZXJ4rvQ2qHDDpAFPaDhKliNHHFj1wr/H48VkKRn8E//kCJ3+qGWr4TFw2SPPD58ORB
4EtFGDBIfGZxoDiZ8LaWo8b5bHnl16r37LL7YNw9muETRR2oWcxAo50rzoSRift2TGM7+AyI0szz
SE/kiOx51rLscv8pNm6QOAz0ZivJTM4ZlUfFNuofjZMNGHbdyWSPR63JuDeKny8j1BswT/Mn8B4+
+i6N+EkEr3PnvECWnysAiuRbfwOCTBww3T4eNkXovIxo+Ss+s9/FszuhvBZIpb7zUKAUi4xrkZ9Y
Xlv7lzpeSmCbbmmzmhIowFx9PbL/5im40l4b1CJtpphdrdEbP9nn+KWvz1BZyTW4Ru1oD0IE1n3/
Ptw33gaOaqIKiJ+VdxzPOUBDVth/iCzwlEGs+0Fh3iu7FqWJ36badnNc2m63wBpEgVmI1Gd05L18
Q8J+Gvtqond6DU9gkFQP+yZqcVFbH0SfYY5EOfOnDeafIhxdiU8m18lSoqlZW3laCtF4bo12Tnzw
+ijD0o8z4HBNMkMz9VcArbsJ9RCeC9b6x5HPcZPpI1ExCEx+Hl+VZYzPl3fQ8+W5YYDHFH+bBAB8
vaXH66E9wN/msf9jftFNjaas/Nd8WBkfXnaHdjAZcOCnntqrQiKMq1gBSCsOcxTmGyog2vTH1Esn
w9i9khLURtHu2gy49gL3JIiG1ymV6jpMQfa0n+vA4kT6XVM7kLTXFjufRo/CouNUXm625KfTY2/l
6RIl3JR1xgXYiB78VK6WK3nRhJZn21dojtNWb/eZJyuctbkh1lKZXF1Y6l4L5j0eIggizVdXJ3Au
TZkuiNmGf079R9txed/9biRcehA0PxpLXYMBsIKeNZqXDBKB2l5mtf7CDFYOr7UpHVINVDsZV4H7
+4zarIub/iL+uP7NezC4MPffp7TQES2HAkTRTaszGnRNbqt0CDg77WU3zHlP/EUWUlhSbhM/GBCJ
iBWtqpDWE4f2EdOG9cvLmrNTNGTD/4ZD/5zQAh/qBmJpJLO9opWlyNFs9CD5c/ojAyh8pLM/5GM2
593TjGa33MY1Af07CkfBUsoDhBtzNVGWuGpkShxw1Tqd0YT3qwETuNNqvlA4g3Ufh3RpUnsCHTXh
edo71sycE6bK+xzBDO+A0VwrIxG56J9Pt0d/gbHGARjebB3LG8sW8ohA1T8tHDbdC6VMuPetc1rL
qYfNUwsv2UMh4mvOpgjnzyc/hPIlolapiuC5NE/wrt8irG+uEk1tH7eaXIs99740NL2RA+HmEKoO
RcRLXDpySk3jQwSU/B3XWgw6EIdsdQKO6Is68yyYAvxVJIK08Eh8wdAG9OmrOHoladizW2AGaUJL
NDIufhc4Wl8iCenG9xEqi9Eowf+rmbL0GzCVgiNwMMbwI4laFZNgI0p5W42fG6FGx95np0AdMUyr
NAsXKM7xnoX7gFaVARIdbqhcJauiE8nBp2AWYbqIB6AXLUv9/RO/36M70RdvCu+PQqHYM42z793e
dcyvgNDP+hrrKLwIrtW3gdQDqg1WxiVsoHMvW03D4gMuUuJT57IlHiEx0X24n1BUu5L09ZEZrKo0
5BjpX4kwazlhSLjZiycGWfrbqIJlGmnN9r8b7fSBqFMwuOWEGuCyIUQvOKgcaD/q/UKnXQi1Ucpi
DH0/NewiwnpRryorCC8Ul9o5qr+meZchQwJPBKWVmBCWktqkDFDgJ7yjDtCHZ2Bo5qzMVvqo6XfZ
4eMuHID15ZZO/Lx8qxxxF/XJIg1SIMXoYw8B2SFIrvsneaZfYR7wnmOoducQGeKBl2WNp87AUqyL
Tv7yO/bLWhfsbIqwl+b5M1Z+cSQRYtZPchuuDP0oMGEdi834sjF8OAKFQLkCuvEPfCcEY4wGfy7M
Ku0EQETy8qhjjNrQF3I5K8qxOSXXQA8/SYG4Px1A2GGBIZeYy6PzKGX66Je0mQgWC9S6mwkawEco
hwd/p9sOwsgiSi1t/lsvgh2fZD5VnCYJ4YWY/42KRV1GmgLvuLA0Bl4RhfIJX0u7PpzlPl32GTER
LPhSA0DriyLPJwI0kUWuKXxh2M4oI+hu1vnjm4cpxm4FZFn+9QO6wOilU1bdMXZryT3DdHwjxfzG
bHtfBYarTVNQuW5I0E5xK2gc39CcN0eP4TXAOCMy0xr+0dgdk1E3nb+TuesI1lHQr6rfFmdXQe7D
+ZXl26ZA5FAg9GrKXHcZhGnP+pLHtmwhDQDjc2qu50s7vW4X9VAaJgeVAQsFyWt6+REg5ifArd6m
DHYjlAk9fuO4Mox1BARK08xFngceUa4gNEL7HPYmx2aYrgwWwyODN9k58tSKJBze/dlHK9qv5d9T
tYlTUumVLQRjtBdkahxOlDpR7cKx0ZxbGhls0GB0gZp10hRCSroUBZmcT6tr/zyMkHlyAtFmd2/t
NdiKfVRtgFaSlpIuQAnX7WckSf6q3R91Sachadqe0hFUT7YTHZd5raep2ryLN7uX6SnhOi4YRhO1
PVu5GvdCuF0lxdJSfzGZTS0BNeBf3jIgBRAMNXDLiUKcQMTxzE64rBo9s8iluOvNP06MLceCky1P
Mk2nFmOjQJL/c+84+/inW44xiFODErBzCIYSK8i9oCONLWhE3Ljtn5BM3ClXeTQ77CsRaA0fhq6P
+umBGqDRP/Uc+0IQN9fUp5eyGaAER2Kb1XKU3nqvbEjFib1SHdpy3nBAKgYNXzBIADME5AyFeH9/
DEwTmZR6CpSaXlm+LejNPvaXMWjss/UURVx0q6xOGahAXNj0BGrRPZY1ARV+C7XtqGrUfBH7JOo4
yFs99MbS/XAHK3q2zggqYAJ2gRRKw4mS9RDWV5+BLDjWSd6lMn7xcw4GNm+sSzItXzLcUoI3PY85
WuwYu96Z4Mio7v0bz74uVTcBTPuajhBPBzx++gLY3PP+VwACvcRG0o8KO8utXWkAi3bKbI6rewbh
KCR25tzx8JUi6JNBYfo8I1rs5fiHBGyFVtksedJYxUj2rwd1Yqy0CUV8yhF9asAxtu8wqbEWvxvt
D/v2sinSUEq+9ly4eFbq5/Vt95McnPTcJGNw/A3RQDa9+OMbaffBLUUIAVR9hY2a6AeBL1IeumYq
y9m2SCqMJBsbtXXc5cw9jakLK6XUrlI4YAohEmNxIok3WB/I0ORhqVMvdNU5CCs13GVB1AsrxWI0
rg9s6PPlf5NuUo7wP8g8l5b6FsqFdESHxmlKf2nqNSr2/YeJL7yjujxUXFCAx9eyG1n9wxrPBToq
v9hhV147rMuvLo/v8+Za5H59fDs8eR7oB960YA933uGO0EYbfOBk8Ws6nIfaFR2YbwwGJcuOjM2R
ySBjJsmKBBbYnwKDc2jpczRI5RHYq6J5kRbzEea5Q04/jX5bNKWqFNR6mJMTyGcgZ1T13sVZ3N7A
fPInyir3I1x9sMCBcwRVLNSUwSgVXcJ2JEPWGig2PWDWpMjXBeNFz4/CPNufqF0X3G+b3mNHYdM/
99VNvntgsEh+QYdQ/0BaMLeNh7QsPLQEfh8DNgLqknAxWY2FFI28AOUbMkt79RcMNWdJ081onhK1
dy/JwOoXDOL1uLcTFWyK2BE0HnXuMrk+BPiKYDIpRU6Ah+PEw9bd+EMaEnY0na5LB64h0DoYXaDd
zbhjWPKwMJt5Cvq/jBBvChmb1pv1kw1/oobDKPTvkStIBNpn12Jhy5MhQYOLflVf+gh/sVP4d3Xp
uf6oTjhwlUYRCPbsHln2zyoNzyXvnA885sJabOx52ruQbW+RtgdBHQccl7MAHS6C2riSgpRNG5qW
pRyj+u7Iofk08DW2TGvzpRVm4rex4fA2Pw3+BGWVL8huPJfyfqJ4cZViJX6lxTFhrkBBrrHh/XmB
oez+u6ohiimVlfgJHRvrb3kiQ3GFf/ZfxPcln3Fla/3Aj69da7+TSkydMkWrQ8XkujhAHuswBwav
6u/k93nJbtiXLfWRRkT4RqJ5Q+4hSbdn8aKL14AWc9ZmQxe8KbzDKOddriJSPmgTzaNd2B28B5HF
scNGPjGnATveQ//ZLQO76sg4gVnVMa01uAYwWBnk/OyJc+O49igtGaTXb2Qgn+/vX97GRwMG+5CW
oD1pFpy4K+6rISAC9EUIki5IdVCrzSqi70fHQf/HoIaVNMjeOvJlEoQzZaw2J2Tr+EPLTcPtfA4V
CB6PLYctLmaobtHXjq4UC7MxUo9pTjqVY9P5C5FVgtsnqUS6En9klCwgDj24TebxotLVITWKHl+z
IeAYWePhyahl12loB4SE1pKXIGo2UGgWE38lfB+CQp1XLopXm1hJiQwTiZ9iwLpFFgzcwrLZCPf5
B2auVhdoDnDlaAlCB95xAm4HtrkfCprJrStDq8MiBzTN5N9fZCfd/nN1xk8M96rHVIRwilFK5aa3
i1qQvuL9UlTzzOT0hveI9LkwTfjhixC9UsWEBxS5CgMhQsuJfe7lKqJGS7RyH1ZaH3s2/pfyE/Qj
tyLyS5dfVqDnJNIuZPTokGbLLUXwOVj6TU8HJa01zRhRBJAKgEgQs4UBN0VsSADhGjMiRUBKaHhZ
OBxFw8XOTeckG1pbP0IPjeoOxBQMeX2I8oL+i9tLqbVoQv+P7dmo8b519C37zQ/hj/p4aFJZcU8b
yYpUudebG/A0u0ff9Yt+hVmZ21PlLTC1YQQwV+JhrqQnIrRdEWpPT7eqlyzZLm7ubKhJptrxGL8/
Wc7NjG8V4L8PlftebSsjHbk/hKZAQR6QoN7qd8zhCEafFs30QtYWxS9hnRSv+TzKGV4RtSgMHGcn
UsQZcBZ1HgK/nrFaV7EW9LEhP87i/ZAsl3WPQ9TVrB6e2Kwa/GOMwsEDq49AON+ONwRov9V52H5C
xWxo9W6K3uyFY5GRKDo644xTGExK1ZAYuUpkigaFw+3949md+3gx6L6fKS5m6KtyXo3gjvJuWg1E
EioRllHFn8eNz6R7UvQ9m3uLb3MjgTMKIKaxt9qwcdiNMwKq4W7ZH6KVphxckMf/DPoqfXJCZBT1
qyToXVbjB5NHJIt4MlZTtEHxzCmJMmZcgBNi3U5dW6D2TNsPvRJx4LqKPOFuQjZldRgW2qA0AWlh
OskmvK51aZfEaR40xP177iSCfEY6D/wFXG+Bp70BZo7TBciz4JXJveYSbOTe41iTDjyJA6nllPQJ
y4xgQrgb9J81jSgqG9EnWQLIL9bes+PwNdwJ/5EYIRedG29ipvzARYxv0aY+8QRVeDpVrvIvRGgh
whJzU3t34zniXI9CK7nGdB8Iz/uUvyO3JmQNa4+lDVrE1U+IhneVZe/3y6A0WPkGCjoffTn4Eea7
YYr51R9q0tvy7G05JIRC1bdPuO+Ou6h2uaJzYZP9z4EhrPrC/2MmKU+oCvX2tXnB1IEjDtxoDZvd
ylSQWluHRM5iuGjSniYFxDElhxhFTtHnr9HXci3M406in2ozqP40RYoNiGk0Y5uIjaRe0kqcLUkY
S1DqLH+nckNl40EXQOb+MiBgaVu56iESEoZ797kCdVvF6vba0Bnb37DUd+jQVpGD9tJHQGEPm3RO
QbqNdeMKzTY1XSfh6V27nSFLJ8JeTzWirkPNFEdrVioQStO+Zdx7qMw0iNRV29JSogXV3+yCqs7K
SLhw9Oh3ll3W8ktsuMxLbXubbl2Lo7LPiyJw52uUW/mKuIWP3tFfDWJ1j8F1WIMPAdyZP1JlibaV
seZSAe6deFT6I4LOwE6L6ExwqI3gHga4AB2WEVb8lHUBj3lwMO6Q4m9KU1KWAfMcpA2TRfPpD2fK
jdo8Mndv+Ypp7NoReK3F5hrVWC7ry1gtj2MQO2g/SciHrEHmTjfhLCEMlVhfde0QJeepCiL2stI5
so6Jd8zE02/2jcQjw1NZ7GyhfbPDTHlQG0w9VlJ0UE2u6MfMwPp/M3hQfqfAc9BlMGlbhF8Ivwe4
D0Rcprx7bdcFQtuovaO9mk0mwl3TIwxxz+ro7ZclTir35YeIibY36Cx7ndRMkEqZGrjDO+Cq7sPK
h6b3sKA62cAOntyqf6N80UuNKKyrOjcmz89glDCi9l9BwlC2+ObWwLWMk8WU1JUNqIwDLsyyYKsN
unviAZMkHr+UfpNxnfe5yufmLPoK2CaxkC+jAzzcUmBnUrQSwgg0Ql3HFvac/G+92aNxF1JtYfU5
+VPIb2gaSxFfG4RR7dS0slED1VVYevYBWfDudAfUznvoZrRTLkxloYRBDYwEbUw2SFAok453HCme
ZgcXjwB95QMD22DIrL4/NihZA0JfYYfWBDsmHWEGZo4ETWhgeJ2mcWROFcKAULL1ResG7fV7VUqW
QQJ+k8/AHUqiagv3Z2dzMTueK4d7NsgoeE38swTT8UYmSNDp/EQ61ghgLHICF6f6uivDSh0anuOO
NuEH77/QTSg+pDw9B42JVP07xq9iJmPLbSNNoyBONCQru1p93wDsS7mFF5dwNAu0YUrntzaZyftA
peZfBERXQRaMQQUtOFaFrBkDj2ZzGRmZl44BjEgpc58koMCjKgP0Vgh/FYsvOl7sPvzJ0dJUztwV
1s3Xi01Ok2brJvKx3wukvotWGvyc2ryZIKTDFcuPKo8caYDv7MSquErU28lCFRIivMBRBr2zvDtR
hpwmRNd3Y+ZJXoSPzRCF7Mgwz851WMX127pdMrLHJPJ4PF/6Qdkw0jdYAFsGI1ho5l1+LUGhnj7t
ZiZBHReOu/itHxWDWNbIUuVa4Xtd8ieAvwu6/oW8d0AziTUSyusIJswkad1pX7ReGOh8hzMwCdh4
LbxI8Ez6ZWT6JhQfFCvFPUITCyaPbokN9XjGv3C1/ULt6UAN+72F9qHkKjqwsyliobPtmvha3KD+
7Vtrj0+bi5iezucb0pq5pP8y2A/aNsrxiyDNfY+WNh32quy9ro1q7SOhMjVoTpR6o0FT1sBtQ9LE
oX26s5DLzPYQsFb9oSk5wQNgh7lrRwiIXLP0JPchKoyQ5mp2+dwuxZVsNtEHh3YB7DVgcCfSMLwG
ijgoTJ7Ta80viBo8Tkn4FYDCEiOtGkTfe2WJEH91+/tpusfniXFPbf5+BlpKyTMxwklQ/DvzwSSQ
AEopEbkA6EuQkGOHdTwwL3XduJSAPvN7TnIl0gxWDA1epbwLLwKT0Gq2WvefTU3wdwBs7J4kNWP/
zqA89x6E2K/R57Y9huhpUGoO096kHT6efB9nu+5ORMCuPKTox+LbODQPqMK6XS9ii8zOS+jyYy9C
VhBS7Q7p63SANXdX5u7kjS09KOpu8H9rVHb8/8jmvhUv+k497Larh0hdnGtP3uLOYUqh6cEAGJ50
NY46cHqkJq7gMUVRdnUw9KMDLH2o7LNZ+B3kq6JiNEaM8GmIJKxNULbosCcxRQSgXjClcrRJOyL5
HvHzzP4TewpG2g7qd2L2iP4QlDHKy/1knGHjM9bQj+naHgTxQr/j1KQZder1q7LVgKIZxrBiZFug
cKFtBlAtPf3khYETmkqnjFWijQ9/Dx253Odhz3DywRC3rASIV5iOD+XgdPnPLiIFNHLT1BMcGkjA
K7JK7bucZQVVtEz8S1pZZkPgGK7fd0QcBLd++44gpAtcK9as12vfcrSPsZouukWbTKEZWDVAjAIC
wvmaDjLh6sVN+oAepFpF8CthkQ255DxGnjvtKQK0tlrzOANDITOde0nrhd/CUt7K9qGu+utc5vI7
Uw1IyGeWyEuLJB9cO4mbAdy5xWE+rcw+FnCrjrJ2x0JTQEc7tBjLTzrTvPKPm0Bxh1SLtU/ILKI7
EnmHwE0Jg64HwlgVmpTuXW4HzYLOrMGbEaeX9p0/Ba5paDIKPitrOlwaVSgcGRxfgSzrNxyKFiTu
Qb5FrliphBdQPSeNEkfWxfJT8u8OuRJNGylBW1rE5pWsAZVSV+OI4iZves/wk8BzxTMQJg0UrEmn
5aNw3gU4JzCWL00SjHyg/nMOScewiyi5WgQGbtG6rNyNY1H4TA979G31E0rmqJvQIRRCTk+/PiYU
bZ46Dr8I0p0iTUKAQGyNXqPrFvwoAneJ3MLYN1X12bzfMelo2wF1zYFxSCtqLi6W8TXpj1zfdEoG
DUmzD1WPbUyP+sMecbYssoEaWV7U5mX/aJkx+mdQTtL/XNYt/fD3Ud6QcwSxT9EZu/BDRTrdfXq5
em2NsrOrm/fWBTgN0tpD5OYn6XyTpa6UHrEOR1Pz4fKZa7CIkyYAanCG1KDyZiszTrxIl31Olt23
p69tk0omVCP5JXB/jStZsyxp1w798CMULv7LUrUaj7efHLnO4D5PyDOzqitJdTPOuGvwetwQdnVC
QCuQxlfiOBnN3F8E0yMTKXXuf7/wgAdItmAy3AlMcBpnBQ97TU3GClRYL7Hm7wcN1HiR8MEM8h1b
GmpLjc6w8nWrE3L9n27lz/XZHOFqdN5+4qpbEme63FehRftdgbZYNWjbWyz+uniHGZ0yqEyhGV+e
6hxgzvt87SdJ2l6uDAPl+GFxOkY/3DoVXZxNXA0AN+soPFFH/wsTSzENUQv1Ibtfos+MmXKYc26y
n/WVun4dLPtdWmKhVecoe/gTBHiVOpMvIpAbz33XmooM/ewGLRyubBmhA7Wn3SPJG0htYP2QSIvl
cF7oD9Y2M3+RshTcIW3JubG2gTzy6/WlFRnGOAcihj9+CJV0R/cVb0kBLWiHxrIDelB5lXUCCjXE
nJarjGwQFjoJkQshhKJ2c0ZsSO1bhoXmDR6P3xCCxV4P3tPnHOlkLML+JD6p2kz4BY4UM02D2N19
SFiw3CrdYYdeqho6vWdgfYbUT3xzOdKgiam+3ASrBHUNVEiqnCApa4IiC3Nw/qFOKcJuIZQ35fcx
CBv4Y0O1wfbD4SN0fRCiakVPKebtG7lJEWM3NcAwOXfhFzYzCqq9RnL+CpLQQH8pagfJGg1H9SzV
JvtcWiAypTbMe4FIQeaGI5c/dDf0f9x/9DZV19hVmN0KIObKxBVtqirdTXJDqu/ONk8OWDgb8HqW
rwiWYEdNUmhpUWuN7nygFJLCHi/BDzoSEvti+692uk5ajJeWSYdoAxU2DEp3UN0KaOaPD0ajJHSQ
iNDeFpcJxTvt3WiO8SEoZc5KymN1vzQlfeohJxmXrHZODrkYg4eWABhFJfuUhptuXM61z5wq7NqH
p0wuOh2u+4KvDrjbIwkNmWi1naY84LZrQ52Kzy29DUrBzA5ub3pIxEn0OR+8Sk4X75T54cxFk7OD
+IsUZboZvJACWUUqI061UJz9yQddE+u4wYKngyWXVA/LLHK5R4gsFADN8i1gSnjciW5dJMOe665j
q4LTmwlfrMQDoFdqUe33EnRJ7fV41IDzfSXQKuZWRn1HphsYvJEsWodVinDnECvPgfi5lHP/RexN
SEk6f2iHxupuFsX/ar0WRLvKiJhyxVwb9an1J7f2r0bhJSq23Mm6wMQ6ALb1P2PzLDy/koM6p91h
mjH05Od2ND2hd90jh4EYhPqlN6EENsiJBKBzHJwTaJicgG6nct/BUeEHFl00BtRsUf3IdUguHc7y
ZEEIrsIRq8heKveNBxNssmo/7r97EQ1QAX6YxvNSp4J18U37Vqv78wjySo/Aghrc+8PuPJdwoXFg
5hsZpsfyRHZZTNP3PU9O0QqYWNQFNNKZUiBuUXgbTRwCocvcx3apEuZo9A+ilWaEoi6NwXJNyq4L
+DwyTfLrq38AsX1wHmNEwTpiFLugE2UyoW+MnGzqxwavwgnMdmAk2iC3sjSkYokwDHYBtzxZvF+1
FkE9bSk+OvjK0vETXwAXkeY/VUmYODDTWQqXyPuaZhM2sjZXUjET2FFqoXFRC9OcX1psxlUh+Swr
kyeWMzOwMj2Di9kcgZJyIMyOXrRvfcJO4MUknapKzYUGLkjIpASUaTCr/JtxiJ+CfPV4UjDZaVBW
8tFjYpuTwYCdCjym0cCSZWqugVtLvfcIjZm3DGanPIjPnb3/KMtmWAU1gJcsXYSxgObtXi3Eqh0u
auLIkebTFqlK/MmnxeyAK5z0No+8MDUCOs074XZPh4Md8e2O50boFiDoBbDKgrourjFcQgmTG+xn
pABisOjJ3hjMXKKMfougizuTP1bv6yCp63vxGRI9aMBuzceta1b+m6TnY1jwqgQ+T4CJHWKEBUG3
5Yu5kZU3C3W8k8q0bxV65VVYCoG8x5TBZbCQJo/vRtoF6DlrH8xQ7rZif0BsNjkN6OT9SJ44huWz
UWapr3DvzBV3roBROcxfF72rXuzy6jbkgn5KChRLnJAI9ZrB+nuUTQLn+T4aP459Jdd6yL09TGXN
20StZBsK6Xqfa8ztTipxVk9ogLjmJ7FDD8FrWWfXqxtHpPr0rbNfFeXHjkBo3BubSnCienAVNXlE
8rF+O9oZNc7a1pvh7QWM0NPcdGbi+XwjobFwEm+NWi1nozCauGmrImy/uuNKrAAJVzM1RExCg6wX
8uWvCpSyagKr/zYwENB/AKjvIY8BMFBmlIHrxPVilzmj4bArNlJbbvAidqpqIw4c9e4TtlV+0wJV
dHzhDu0jWNtlilfL5ExcERYRqNCxgzF3cY+DhSz+2+yJv+EQwWNfAYLZro/p92yxGJ8iG0PRhpiS
2XEF2y3EMR1BoSkh3SIszHB5A0upBetu5M85Pto4xLS6MyWBWSIxyXc94yQtXPIoGEfis2Fwe4h5
XBHEjEszeQF7ZPbqz72xMiyca373RK/QXQzF6IPgm2IY5jSBphZtvoNLftBEVMWU+7ukmRuNwtxP
eBEjGYmeRvmJNP0cTHU6R5CbmBvBaP5y53YFFyyweszSzbYvXmpnludvuOvr/iHvEtSvCu+xb3wc
umjaDCCtGp027+Zyagsx+qnHhF4QmKEKs4MmAZHCYX+n7rCQ7ahzwXULv4P7O6XfKC21SGOyqang
vqBsclAEvnZolqpTtDaVu1kW5QU9N4s8O+Ewfpe/Kjjr4FeXvkUaftTZkGc/225B/f+sn9xJnCpJ
oaHxv+7zoL7Ef3s2fH+4ZfczSgxsTkxvH4SIUOiXRnx5B/ZBuBEGtWgNQaBTGodt2q1BRm8EO7NF
kIUDxLOh3TGtPHsG/7rU/kdn+jrDpsQXdFNERrZ7Nak+TOHckLsRca7SKEVaZcRs4BrNjE6FoQUx
M2X/BdlfQR3XItF/1r5+z93mZd10AQtWAI3Wm1EZSvb0zh1mwyd6UIkObC2TrxiXEwlOC54z0PjK
o3dzchZIBOejNN0gFhJHiTthVpCsGaw9H9ydWOVvTli8T6z6c9pk2bYJY8LUEq7XcxzdK9wXoqPF
pk0uqV45IBgF2uYb3JkKyixKx07Jt20xAJpQVCFyF2n5XXeRvniHT8gNq4/8ruEjvwLDOoLHMK9A
pNucZPVWWz21QIOXjJ6vtlplXDH+5AFV3CEVeIG0brmIQdIZzBszYbo5eWGhlKMiYXYwihAiWMtv
5U8x1MJhfUj2m3FWJKmHL7kgSTlGSo2pNzepapIsZ/nReliCu+ZZXdFR+uYkkb9bYXpSE/ArjGOB
KGHxbLzYNt2pW43OO9L6+EnJkj61cINjaeeL3bfjXKJtpgpjStFvK54X95N9rFePpGMh5rybzEkp
LrJuBLrYxJ70qO2egphHN8hJb0aK3yoWjWpwFKLdY0SD10fxyzLH43oFP+kLGql+Mqcn9vH7cFDE
Qnv84mJSblJd2VjpbYOwYnfW5et9xyoeVJnNKhCogbymsSXodZP/v5t8/Nrm7gdoUcjzpUKDb0yc
jXSXsFZF4NKGam9+H9GNEtuwclh3sGgDeUdI6TlTUZNFsrRpgfSHvSe0cEAHqGQ7/PsqQxcafxVh
7YgNrqheKpAx5lXJQKxVimeEM9akDl/XJ8PCfHCtAD9BKuBd7fow8F1WSSNU9jbUGSFpktuY7XtZ
VtfR/wYsLYdIlU+k7NouRSDMkB8CRKSLoi7pz72uVMTvlEfRSc6e9YaUvDljj8OyudIgBvc61SAI
TuhFcn7GdsuV5XqICa0Q79gFgkAHOb1OCGJwqeN0g68iGz+8PHUwRtpidZp4UcOlWO+fLBbhfXkq
Zp0h4ywyMVVWbCnHxNqYIZXVc5DPH38kSgFmeqyt27+8adF9lK61ctSTL3N/4UVAN0nMDqgByJ3h
wYVSyJMcaO90K5XZg+YORAS6KDczw36n+eRvVpPxZggoB6Eep0kwXFlZsqoImYRP5H2XQsOiuIm5
udh80hd0irqQNEy5rs6L/PuQRd/93mTUP8tCICYqxJfn9j0YulrJhX2Hw6EUlEHqn9R6PSxbZWk6
lxQwYNwxbe43OBE9QIWGPUnWGSvvtHZd8CSmapgaIC6np3hNVaknhWBO7YIEWq6Arq1ttKXFcKmC
7kdfoDpfxIVE9yGPWWFa9jWgHMwZ+LVKObT+jXsJiLeiOl3u9VOQe9adnzGKynhO4TsM7WubwXki
bKYjpyku5iwRQCJKetp4WE6qxjcCZaN94VtYbfx1lkPHO+E1UL6XfxZyr9bGuCL308aWtsE65ooD
tDC6Q9CnJXZ4ln0TqOg9Q2vcPF20Jj+vJQ4xOKMcN7I0cazvLTLErH/J7VY7YFTZ/tCupyeTbyk+
++DWCQyqfNwJulh7TORdeSVkZ4saN/9V973arRV8djkWIDzTH+cK4CYshTczUN7tKBI14/jOWRX7
qLQoS+u2T/+6n522WD2pDrFxNG7hWAe4A0ksauk0EQcgaWzhra5hK3IhHZDyRsDsgN6HwtU1ak8I
L3BlQ1xzHOHD1VbrOHkck+nt5lbtVmQh8tgkLJrG6z+yMcjySrZAjAHcwGRpKLlzVg3BXFeDedNd
zZO+jQH+rHHMROQf8GKZfenR+cu3APterLX2rq1m0vfRRedhGSLJHfPXJ/aHUUbir7i6IVTkYJQ3
nwF269MsawbVgEiX1aPQJSYdWDIm0BSUkLM8LmH8j7Mw0HhfeqgwLLKWDpFQ004gZgvt/fO8H8om
vxY0yCMAqtxxcSyACbGmUCdsN76L/P1HNm6PPMe/4G3cmYoVf8pT3cFr48f+BbRlSkgXbZfq4USN
Z2rSpKzDAKlZmgN5MB/Effg2Mu91ox0E8tJzVCwjiYKx9jgsRFODZ/2Dft7ifYBsfuH+mhiY0mzl
mo8ELnRRa8bKDF7QxH5Cjl6F6Amugo5/fjIt5H2GCmNXghyel7q/AmUHjxAXKDpUBVs3PgTdVxWH
j/uyfSU074xaT01hOOUOjNfqPT+tGXgAiN18ppfK4D+mF5SBWAQr2Pwl+N8U7QESbbuqxQgHnNQg
A/nhSERHhk0v4EDBmXrG24QIok0A+MbzRzpOGHsWkDIrtEzt9WmyGPnAL5sIU25C+v/jurTaoM7g
hasTwDpZLhk1FG6QoOFp8w1muIIySFjYItz9+JHp9HCaxq8l+WApouKbFlEHR3GFh35A5TpE38Rm
dvO6vjVUKrapdhNtW4h8N5mfRV6ZyBcYj8fJaAE9MWv2vhDJopLhVtqII0D4IfWrta2uQbTcSa2E
WV58YWmWL9viOdH/yzXK4BHxjoJZgYnw4wUU3VEYINM01qTA+8BjXvudFlFDwFqnxLSlsslIhoK1
gAEsRAqyBpo1r7V/tzgOa05sm/Abe47O8BrvkEPyVplM9uao6Q2C1lfKdOvJ4mSmEhdXkeWX/umA
Ycrdgd3CwTRQDuA/EzvhMmwzROntnIlQDQc7halKwIpoLksdLxbENPZ+p/IdQS+W0BOlaMAsBjKK
bt/hvSPGLXhub4KyJ9SPtQJNd+F3JV1mUsnhOClfrlVw6P9xRW67USON0ytxmOmgG68NAn5pEVxk
qjTqnU8Ch2ujIl2i0QwGIHI5mWdIroP/+3Qb1I6zPk7unVN6cHP/5G7O+GInSvLBp0QG7pBhCrob
ZDLUC157IbKEeVcnrGLGM7uL3i17fQDuVluTHyi/UZvOvAR3BHZRawq3BZCvdlxrbDOqGK6g8twQ
r3Y2HkQ3Kt843xuE9GW4WJTCmPM9f+DmCfN0ciTwc3FyFl/LMkB1Ggb564N7hsBNIPxYScl3bvaz
CxQeDF9QFckUdN7Z23ohO9EBnFF6kf2f+oUHbglbeQc2hCi6m6l71o7YH2VvAnMVe4SUjEwlTNwR
LIvon33eFdYMXFv0YUc2/uO7sAW1faxlMdjGRj8B3+E5aVZVVT2iISR8H3bKSxzQVKh9wN1G5oEp
QqLcNmhifur3z3suY+bRJ5oUe2i01TJZXVJCtlphVxl7C92oqZp90v0+1yhhufg0wlXpqwmM5xRI
gnQcRx9kAvOLCkVXEo/sZhI9dL6ln6ty1TrrCXzgxLouY7JsI2I0q7ehzdMpEANK0ENSGbrsZZil
obgycWJoFhwISTJ3BIII6fDEhI1q9OX053wUI3rOmMRuZyU6SwM7QjWQteX3Ys3Fek+TbPUPxS4t
X9Etib0ngwf/b4Fg7syz6s6QtRjXGy7pp7eAAygBw7qGK1UReJ9kY+50eKsHhPRq7ZZo1JlMc7kw
7Kp82X8NaMlSDyfIK/ClGeK5Vbbjm8KRj9spsa3XLRKGiz6cJtcPcTzVwOJt1Qn5162spxf6WM0r
0++i4H7pVwz6rvIZ73zWLXHPzJ8NVxeIzE+6dhuPf5q2+/VCFRx4QPveg+aSNX/f9Lq65rEbK3PF
nfbvzv/mwRx/bgs/JVBebuS2xIsQnUcYC8ivdj5KQe69t20Ql3X45m5ijBxGDP0ctk9djANUZqZz
9AMBLL4nIdxKJSvXQ7UApr2KGY7MMNanAzwqlSWZJTC/hQIqLligubSY6NXNDh1VHfiHA/OCm848
imRGOfZAaIeioRbdDuKDwXDvTIQc5aWb5AX+nXP2eWUSqWt99ODDea6gsBdfxfo2aemmjv69qe+/
om0VuWKD2FKrYcN/GL+2ukgKO21MM747NWi41dLK4LpF1o5A7bl0Td7hWD9h6o9ng97yx2D8EiU9
Wyk0lfCYv1/jhD7cw4IWS79iogxXPNDjEdFSVL/qFIxXxPSUqodMffLWXBYTIHSUTfNWW6LWrtBz
vD3ahDBhEOb3s9Em+e0RvPIc6X3/cyOPiiiDft+3MbtDLV9bDAAqmDrihoQmRdYi+CNT9L/hNW/C
cAaihs/11b7gzO9nLkNJIYoqq3s7Mb7MKp5X2AALy482KOCutaoJcha30uO0F4017eJYJT5Ipijc
pU7hCMi/f4F6thwYK5cbh6rF/yzJG3wqwEW7ESiiD5F9JoMa1JLUxEtQYNOsDI5J6L7aBIKXJJcZ
Xih9g9I0zzhYC51HrS87N57BlUEVE88sW2pW/mPEd2SrGmAY92BblwDfWbDnBrCqxcmVgYBa7X3X
4C6dcYN4FCkCSbBLv4OlvUPo4SYhXxH5J/2KgYxg2xe8efSFvAYXc3RQSC6u0MTugR7QSjkJzuSM
bsKpc8cQDrPfx4WooT4lly50ExXW5pgEWuIAWNWP9Q/1LupA7FMkg4CDXoVcAqRihxDepV7zPGJT
IJpaO76Sevx/no/ivCKb7U+P0P/jK/BfUBs9WpLBftv7bSnDsYkRgxrnOtGEDKUajDoq6ZHTPfHl
6COxkdFqF8Vo8ZElwvQevzSbk1A0E5nhIc50AW2Bp8cQtPdxy94AstlWxq1KR8l9j6RB/1P5ox+0
cRaha+ne9bRIkAHl4OtP46KcXutFbK3EAGMrNphAf9rng6+jvwT4DDAMG2n/pKkh1Ck7dz/F0Y/U
6U9HnTLTI0tAQ66uX0RvOqeR0gYEnGTqZHB721+6imQ83Y8JwFFn5H1jjIGdy6GvocdahWkea8GP
HEg3r98bfr2bxDgQpMkOfZKjvR0MPGRYCE4krvGwm6dyyl4qGcygwXtXyTwI92cib3AHL9PGHs1H
VBd4irIc4yhnel49iwVOdNPUw1rqUaV9qwQt32gF2ch9IfIziAXQwJPWrO0MLIAWjh4/p7gSDAiQ
xcImA2pVeLG9xKlR102EMUD3c8SKauFPwKfF8ZiC9TcZ/XDxGqpJs9KsYgl604fFMDiWTvjf7AF3
f2WRoQGDWwO9gvYNXFtK2Pqte7jTwSPK9E6v5TOckuQVm07uSFZ04ZTYYWwBLXnCLq/5jT0T7nkQ
Wia9zu5QAom7gNHyMqkK5ukjBBVjeJZ/ewUBuSFje1s0R2apizuByz1elloSQgtt306Hya6PSJjH
JxzBurHJKMxxUt4rhYkrZTS1JAx/7kGBQ1RmvUKfH42Eg02FXn4LNeFMuUswYr5uIirjIDTKeDuu
ByKmwx2WzaK2UFSOqfFvoELY1DQcgMxgcGMLZjJWfCmxEuEJSmzFHIAQDrIsnekTKAGKRE4cLw1J
U1RUs0awY5xP7urI32jb8clPcNi6IaGYYTSllVh7EIn/rfddoaPrknBKd86mShKFhIWOzsBZNXHg
Q6/hQz7hoexD9IPs1bS6pnBliW2xyStVTAQRJ8FpVLW6wjjKoDzw0R7rqaEWOYh/RLgm9i14bnnC
9PfnxBGnettKoG6fKsviO+Z1TcRvG+fYLUkb/4HCNGUoind5OhwhxZDUADoOZg8/XgGKXFf3J710
IyqhQnM9tAk9Y6KbXhprhE/oIBZwQxgOLsuCDkbydCdSW6mlvrDTCjOHV4CxIw2Dgcc8Inzf0dAW
5zabfterAsfrsWd429eG2wjgE5Eyo0BGWL5t4ozkJXWrpsyZt5xcRGGFMczKEU0PRDgg2zyqVxpN
BJmn4NcDaDoRLWjbtFwty3qZX09kdYzmg2CGbainIdoXh+plc+nVQB3tdSuZZ1mkChQCkMEm3Qxj
6rIdYu43ulZ35RRYCpK8igTDvQE9xUykW5I2bbl6QwqoctK6HrYfb4S2mp/ieG8fRSDvCnT8V4/v
2x1yVkYDRGiWGhvObsdezcNb9sXrNKzS3twpzuL1fqGM+TaRppFoBOatEJl5dg36EqWg5Wn3dCai
Uptxdym5ZokMh0RQ06ZxR2etd83KDk9TYwZBVJS26Bp3XT14pf/OzyMvouEYiE+Shv7Je49CF+Vj
wkW/k8wwNcHDfRFGqdin8OzD9fF2ARTKk5VItUsrjuKFS7/cvxAThwauVQss4JDYVFoqi+sK0kFP
nNfMYBZeyQKyLHXbTCLPGjxLaNh9n8TqJH4cTjnSN7iUaSHT7DrotRW5WWfV9hTlFd/ThMic42gw
/JXSq3Op0nFvoIrBBQx3cKnf6W6eMAZGy8HgdxSEE3KDbR024wxPqSaU3gFveO9xmO63UAzph/8w
xyh5p0GV/G6nRNdzgB2e+rf9MMI9uAxEO2Wy/7+J/xkKA4oPyRbBjHkcMS9GK9rIdRMKt4GYNlbY
U9U+tnoumMP2JKUAw2fDoRYYm7n9WAGRhruoJiUfTDq49Y6+TaOAs4u6/IZyfJJGNsKrJNW8fHYC
aSYjC1s57nn6acLsPN4i+4AOP0wh0iO1j+6vr4lft03gZDSM1JL6p1R1nxr/6XsbH831uF4bamEs
6iqn/KiiIoMfOoxtcdNRt9rfQxwGwga9QNwaCOVFWpD/J/kD6WyhuFJTFk8bih8rHCBPyKrBUiFX
CBXeBAjMFCMLD6zbElkJ/OA3HbgJksMIuqxzX3ei+/Xct9aTLwWRdzGcjaasqUcezZKhIjQPGKy3
I670DyZDgwgANgh6ZQ1SHlWVWMKM2fClaDhJ2jEx2mS8UwKHVQQ/FTii34mKiW1XFaAyhRhNWwcs
Y8UUNDQ1f0UjLetOEqT7ugX/ab0sTYWib0PHJA9Idt8Aj/NYiftJ7WtXkVB/mYWQCKB8pFoSC6/O
B49I1jhTzOmKRBBnyUfbgkRvI51PZogdrPZy1RCjcUDQUEx50oHElvfi+IJOTAYjIP/uJ6rqzA75
QjY+bnZ2a+/eFdwA5yTIMQuGV0ndqnDN99ifgV8Dsw92vlJQ7+ZeTgv9opSLOHTln2nacAjyKaRL
Q4qxV8wzzW06fJKyR37hUqKqBLA5ab33hVobsC6VOPeBJPaQ8Z/un4ZkwoK/b5jIWNc793G0A+JH
VD9GF4EYoiYSaYD5eqaaTq2D0B+reSMGRUQ0XiQoz3nyLaa5E1Krv/FulSl/6c91X4wOlMjM0s/7
Z8AMfHE49UaWUj1FpAEvFNlSj1LmBGu09rkyEW4oMxRBKCAaoIVI/bK5pjsc4jj1Flo9YZjrl0Lm
wg9LeYWrYWiV+VNJRSv169MSDYgW9gXalQPVG8CSv+tLQBPqsZ8hGYqj9AQL1HhJhRHdG/0eO1bm
DjwZ7l8DysjZBI5MpORNq4CFSGt+Hb1tLsEbxZOjMuqCH6ocUghFWrdRTAeEHuQCMM6HSF/I9ncC
r2A40Nc8mrb3wsd2zdRp99QZf8kzoM7kUkFCAwlNM6K1NokCyMkcb+pzlakxp8dYGoFUR9yweSZ7
mtAB7mz5ORcrbyWFQhrnQnxWBkGCrlYXmizN9AVOotqW9ydJb0i9sZGSp0lpUyvqEsw+VPaBzXc1
x/PZNILhkzXpbdaxDxvpiXIzgfsr9W3U2Mw7/UgX9bIdh1KwLLby9gKqF86H3iXP0JdNuagh9bPE
SvFWcYX5C+qeoBR4ARCjmYPUmNMbXHhIyRi6UkyQQ8Bv1AP6Kbuz6cHRyza0j922Q53OmBhPR9M6
2W+G+5pXlkZRWGWdNPJElDHl//jK8nbHn7LhWb2BtrjMBalMhNZaGUE6waUDatwN3ErLBdEch+LM
HXXJF1ZS18lGHdp7vLcBu4w6H6i3fYR5RQD6SVGkjN/mvrHcuVSik/bArACvSKZ3Z07W9XUSv8LU
QwZKsIM8L2Xn5UDl/+572tkYH3tOsqgQTQerpxYs96PpS4CIIaojJP9FcWAsZnvDHw03cqw/qGgo
Rh2xUJi9W3OXKVYZRbsIwKidtNsBZUnhCpKfTyShBb/IVDKmJglBL1f5stnruVlFJcHtH6/rBTG6
lQCht410/t/u4Hsj3GIJhK6jZjTvKkjkxYIywpby8qlj+yiHOQ4Y3oYGsSOOVnxTzfZGGAGlC+pt
xcvgCSAn0Up1pOm3BcALunSnj55UtMgzvBdFCDwn3WGrJ2tW4hnDIlf+gGln7S2vOvfxXHez2dK9
mfzA0hvow8PsQH11LqR4bSpxzqhqG0LaCJVeAh/RSt+jDU6Vij/qnn2VfYqFoXoymB/8FlrOMhWh
aAD+ZMRNZcweNNOumG9z6Kq6kYVnIVVJ/fjJ2rvDzUq13RVf3+1ta82pS3MW0DShYnM3F4QkMqEw
Z061pqYyrcPNmgVWG/WTuaNxfWSCKGyIcAT0FJ9mGNruOixMsNFQcYTz5G5qg2SnL/hLULeztlWn
zGySEayqmJ1vRIYCC4kuoPbSQgp8jZWhtduRC68cxKPE2WCecrl/A2L54b+cq3SswC884oDIWGkm
X/akiiyvIqyqFvPNOY6ek/gX5oSOMdmU4BKO5CtnZ3nUdyB7vSoWbiJZ0oIr4wjo77Fa0J3JVR4x
1dovKece8UgZV6XUSxH3R7EpdPGCrdVW3uTr8Q7lDH7xwUs1hfokBIhVO2G8yhUA2g4DbxQZUlVd
l9whT5xx/W8s2rtvsx9bDfvpKnqL1yMYYqBmVWuAKmfmq17ytzNPc3D2QlvcT6xtpiXOPwPPywgL
rdfqKjCnn8SmCRtAP/K+RzjPN+WPS12dcUIwgd15lUuq6AMQKXfxb2+KtqAzHocSWPG6o9LrUIb0
IqJYrWUZi0YBzSNab2wSKeTtqV1bibAM0KJguDaViWcXtq+CWXjHUpgliKEb6lg5/TAgK8FNoQfw
fZc/waD3biybtjxqfkf8085l+P3euKDUkpRjv1e4dr47kn2F1CdqfbnyRS2qWQlWZE1AbHD0GKQb
wL1ypgWzMWvLOFTqyGpcUPE+nMObgVgOWOu9Tf/qMHX+HgUhptz0CgEF7bLJCeHA9/sZhpKi3K1v
lWvx4gVsZiuDPmHyo8poFqnN0wEoIL+BXi0nkueMSkrB4uRgQ9Xp0xKv4Q5uLKbZII53ESyLjL0y
Nw0EpTQRbeWDx+tPjjivQ+VfqCteiMfa4+b5m1hwnAPpWnVZUxEKGOicdZpTaerQjcsMzYMrAAea
4IsZ/cRTdjVznpcyVH0s4F5JjFqOjmiU2//mck0oZnV8gUfqRrORJ7lGzVLnJcR2OEAswsebuPfq
L46aH0oh6Kip+28N2rwIE48E244RBQjwTezlDLJIRxAG37Y4lK4Tqjv3iIvcdQMQa2zjYQQZKby3
T+by7iVpb7EBc0S1BXol+PMgIPRdAQJsCeeCDx6DS4Qcum88S/H/HaEqcgSzwKjeYs5W13nrSbKc
Ztn/vpFpNwhaqKA/gylpVeeVkRa62D5CtuHPRBO/UHkiY+bwGEPSuyr/AwfVUQV9EauRdoA6CdzR
rPGaoga5P6uKlNPkwUxOfQjMCkiN1bB2GBmvCbofqNcStkbh5miFmwLphu8Ab05g57MoX7Yunagt
PyqKtO4P2TXyFhQgSBjYReSMZiOtgIkmD6/LhTTRBR7jLgK078vher7mjBxipvCeuvVe1xMP4HsT
7WTidM0bxRIyKBbdIRMezx8wzTlvCfprJGEKJbOF2medTL8R88pFTTU+aWldVDKkyHesdGnW6/Cj
UNinVW/IprZkyAwRKFJhzV0Go9TkceFxVFish411dD3IpGK3AX0TwY8jRuXSJXBYD6yn5va650u8
l3ZtxCgzFKn6UK80otCh9MR1U7Yvz1P3OOUCIiNM+vr4DIXbS1GknF5OhKMAL4nwrb4gT+o29bW+
Py5+7qZuyIKAfuNecIUB/4sQxtPfCgUlIhj1y8obd8DWFQ8nRNKS3X94QqUkwlq75PyvaE0H6IfW
5Yvh3hEQ0yGHsU5PEmgB2VIZ1HvEmTJTVnn/8/TVvyiE9T8GWqneMFRvYdPhNQXUh1IPjGiU3e6B
hLmMV5l7N55D03w1vZu/SvhzXunn1q5FFivmzdpVc0w+Xwm4iT8VqnKtiV9rChAQEWYZ/1FTZnWr
lIK9hh+yBLnjIRxlcrBx28O+9tR/yV1iuZc3vJtrv/JuTF5EP/vW7NKcSWbv7+DdPcR4OeBDGMAs
idk52PuZdqo1T6zF3FfplXMG5oJffEYzt1h3aVp2n0ZZiLC/roUEVu76Byg5AGw4NTJZrt5Gs3z5
t+RKD42uXRKL6IWuQXsLY4Zrg3yoYxnfT/IzZZlAUXDfulqUX6qfva2ETAVAHYwTsTZFDFHotxuy
HdsxyviHxLlxXBs5RN9eE383ZCXS/6WR97kvOzPyPynm0jSSWGF2FHJiRYYzLY+d6/UpMk4ymoH0
/9Q/3RhffI2+u+2HqiFaM7muTSCFh7oFhQv5zWeO2Ud2ITWexFmmCeS6m2rMY0r2z0ANI3WuzlPc
yMzk6qVod9jTXUGTZiSNgT4j6zIrnFYEFMFmtXUX+wEuRKAaLcSu2tm/woqQE1Qu2RqoRVjpqSiZ
WI112Z6bBXR70oI6r71+rNoymwQRlntlhKhB4VQcGVxcCoqLKc1Y2ohqHjDhRJULl1Ftps7/CodF
7tncPttsf9tLWavo1Zq0Ea4yt1KWfM+dq0HGHDEqBoJqWDC5vA8bIgiK5qrcw8H4cIpVGcez/846
79vUxdviCQM/SUvBfAGItS+5f4iw70ZgZRVg+Hzqfz0eLa5uGnqtqUuDuUxm5FcOzt+GgH5XqjlT
9oJhXzXbPjdk9FO+pbJFWQcDwVZrEBlUTqskwLyF/HCKyrzSSz+5vDfTPYsJjRBW3nkFkj+6HnKm
A048cnDris7FSCJR32XFsgg1BGWoV18pDWYZeEq5IrijQB6Yec8wNwl7lrsWuiUTNlN+rmkgBsrH
uDXgDifwY7Shm8mWfUwgvZIIFz4wFPH4ybob8dpyM6F208E/iFyPThStd8+niibUtL3F3+2dA8IX
DWH+ONBSg1uXbxB08SdWpY0eb6UveBJPEQIIffg9MHM9uSip5w9+/CntqrR7gfhAvaqunwQ679IM
0wLcb4AnU3Gt6MchIRmPUMUbwEvH0/MLmmYnC9QZTbdgGFgHW7awtDHGm8YYrSteHfV6XrnfqxN9
hx9Anqhifj5fXIcgrH+d/WMQvyofCFlbUHTdmxcQ5G2c1+w2SAeuJBmU8y6UcMtNGra0ZrNsCWyx
eGCMI6+jS5ZxHquD1rThNCrE0QWzlCsNrlyxYuEEGe44jTKqgyZg9Dg2KqN83d8+45UBP/1bDWM4
Mm1gMXvWVgJm6c6cMVkMAGlCTMfxJMZODUtKbuYzV4IAOG0VljofgPxBKLGw/3h8PASSI5qPLR4A
FjS0ra4pwCc4OFGPEbJyj0uBbp3nlQFIAkYRZ7/cPHiDqAMP3YU/oZXt5kqFkeT40hULIGqUBiUb
6QHQdNkWgRNj/tiCFBbhiZgV/aBS9cia+cCdSpCNgT/0WNGEHKzq/4XVdxwW4gBQnvFUwxQXn2ZX
GyJY56p7prehS/RwE9H3mHcgx8lf5f1Lb5hQnste03cJSGRpvR/POMrrn7JxSLvqfz3Lbt/pnylt
CTX1rrFuiRqsBGH7dQFN/O64KQj8DBhiGOvfLpFbwT5itEAWHsTEcmHGCMsecOhXZgx+w2y3KUYo
LU5JiDXX+gzPt8F8lwmcJBaGNd1mEVTI7XWmB1/E0hJPUD1mG1K420fnVXiLDpB9KMwRkRx0xLxs
TT0ov+XNhJhykofWeVIMhCxn7A/Awg2VZQ4P8LvnU8ZXGkjSEQjYl+gTZ2htbYHpk6EA1ubi7DrL
JAzYk4QU/kb9ISWcWso9J0Q+jRg/IDmcksvfTMEQxsnA1c23sfsFD8hsrHnmbfNHsGRHzl/ddq2w
YtMfbWqwIxTX4ZybKWP2keY/8VI19/5jF+YbKV7FTnxm69oFICcQdhKYG4uw6WgfmZP1k6JQ3crB
bTvZIFpQg6NLT8FfZkLNbGBadzkmNy8arLRkqurJJ9MPqsDCmEnfcBpz/eowJk+k5A+0JS6V0Vy0
YW0oROaSvpJiYdU2ei+HeZhWw4WjadHlSkm+z1a3pRTWI1i8V2Y60p6ONwOBIScAdVA0BiR1PJHC
yJl3Yh06uRtMCzJLeirQAV05xKFSTjRsRpNwGl+vmokXq22yepnuSLtHBYz5h6BeCG8wEAwTf3qt
t4sshuPKAzNMIAg0b7sgFKcosoRGU8zDSt69Deh4Wj9az7FEiqMoP+HH4CnJ9FK46bGLmDiJYsdx
d/byUR5oXeREluwHA2tsPRwCTmmI7QsR+mJdi6CPKUlLfZ3+rKJLPjDRTTSdU2zUc+LsdOtbs3/A
9TDB4rXZm8QTkUIKb1DoquqJAWXk6+018KljRMqZ7NVs01Q+ISSodl/nMTcJxue5W5FOLbWi7pqY
y7bl6eiKbIrK4OVBTlPgO9J6gsP1uO+c4twyFErhRKbwVXJVpuM+fQQb4rHg5T/3Y8t0O1boOTtQ
Drpq+CnqkocQFkbcn+auPAnl7VMGxitCygqALA5KW1eEpEu6PgLunwC/wBxY1H3d7SacjseJspm/
IPSmlraZVhLC+ZRNluoCI9WrzzHvqOUMZn0HZblifmTnpgyEZywCxWbpUMfUsy9uhZECVZcrTlzx
ndDZpPWcGaSoXdXPgje9c8BHK2fQh7nrM0uHVukK2Bv4W7Z6g3CSjN+gyBoMO2HE2+8Yz0/2wrsM
ajrNVs0CW/BBEGfO4ny4pQwzwMKElBfkD/yjbuRqV48CDve+JSwJVEQ+ocnkZxE0bC2BcWAzQy2d
12NI/clHacSDKJZ89sab5gFje7wZavNR9ox85fyP+KApMIncU44HVrdu6Hiduwi26hQ3ODGcQGGe
Dcynr0D9g1JYJjsDw9ZeJP0P6QGeUIwgKFGCR8Kl9Tkb2oyPd0zV5Opg1J3z37E3kvnfN8yMdOSX
UZuw14FLRYF98PegjbqVd7PN/80ZB6LyQ5J7CB/WdmRStX6CXXf3/SqsKTBaVQumWwPKXterYrKu
0GmeVHgDWUQFEPBXXhD1F/gToIt8m1ErkZYuyP1PEX/LwCMyfB86VBSQDTfIvReuO7xTtfx67kA8
1AJAx1gcPnBDEaWiMD0NrHkHz8ycXsirnL7FqsaqlUhgLAAzm+XvGAOnmMP5GHv+7OKJuYgNpoDT
i+BSEakIM6sZXm4YqlPPl39o/axaJfXaQhvI7parpCzSP9eeHp/lu8GXEYUPb1I2CianQUN+db2T
QR5RdiUMis1fJbleFZonD/rxbsG4k8p8PxNb8OIxwz9jPWvyG6ztcn06/ykKA4/5lFL222tMcsXt
3nn73xXfvIgutG1uE3yDRru+/iUZ0hBRhAJQhZp/OAiNvtttOgt3eC81Ex54q1jhPC6C+SX7Mjfp
418jorpzBfBCDRQp/7QwPvvgdAgScUYAinbBS9AoNdikoCbEqz35odJu5HptVDEb9d4KJTRk//vn
+cJKbOdz+W8cFxzYoOZvxYnjhg9QrPRgpFku+Fl6aDDUticG8wz9DjWXnE0T2Oz/j5RCzZ9LkEe0
tBq7U1swRoW1wEndRGn5SuAvE1vfzmN01oxbMWJbRUuEa0J7YF9U0W3hbDBObqcqvOrXsKRAQR+C
02ceSmYZr7Hv4KDzjRy6MZCrvDf3dmO8tpVXethffp4TiPPgAIQzFL7kePyxC9RFSJVvLNzxnoqg
fG1XOMXz3War23ieM8NXFKyarUjpiKbsAFCIxdVMzhgIA0nVmdvCxsC3hTGyhyPT05LYEnJxP6/6
GO/QnE0AT2GYmYQAJiDun0I5sIZMm4L7MGVIhUejc4n5WdQkpcxrly2XM3Q9gjmZ7PPecxMQ9rNI
8GhmAf/PoRpMZuOs5QSbVGwQN3CUqZvJihL8y5ImRE9VOF3URSo6J/OQSyM48m8SNLU9OgLTiKuA
+ki4KvjBLNqAcvkkHxTxwHcsoTsX6TaCNTfzmm9R8IE/LTrBXK1Uo7kexnK2bFP+h+rmAlx6KH8u
/cPgnY7EdGe/MfBsS0dMVHxuZFtmjP15Z9ef6gzFxUEV276cJu4rK8GkgdUsIXoPVLlDaiz8C6SU
2aik/EQarB17qUogrbiszDWTGOj092yCiH2Iofi7Go5fW/KjlV3C4njnJY10C+X6i+DJIIuR3WQh
wnA/CEvJlpDUOMd+uCxDxrRPVT+Zrn05Wl4aWzENqwbAY4a4he89LZR5v84ShrQfHy6+CqHerEgp
VSuI0yt1Cj1280yf33aNrxEiOUMFGaN8DNPuPTYSTcyYkOe/fX9LkKWWEd8oHQt7ciKWACihq5K2
9v9eb7fmU/gRjlKpUPicWhqYyo1S6lsLMd13cTlSkMxUZ0ZzusF5QM+4/GPGpMBE1X3NjvmgamHk
5UxKN/UnW7sG1Aj1O7vgiWnqaFMNw37d9u6kPrjByAQIZrUTqVI+X9dJj5wiqin5U/80pIITWwdO
2iSljzgJIan0YwybipbxKWCDsiyjsSk9wyDwCAXXB0mGHO5rmfbyyS2Y1HZinWm8/DXTgWS7cET7
TaRdPUvcnf6IPB/PmQULe0uoAxNktzl3jEivebJ/UWzzgdj2ELTmkgeIxVK9MxZguJwyu0JF/FUm
YDpq/hhqV29ux9cNMM0s+9955gALSOT4/fzPdsXYHVhFukO/B+T1VjIhDMalFWMPILhjB9GviCPJ
LY9NLa750/Cv3YX54atNBjcl9LkEHQ2AKr38WnYMNbV6YbwtYu0r0hlXngI5C4/54rZ9zjNgtmia
iVcJ1L5wBSpHeAfzHPCUqxpq/jrB7MSon3jbPiFikGVMICNKwN5fyjXXvCeHcY16JZrTxiMancVV
a/G9z9NPt7XJoAp6r6oCfDnaeTO8CzGSLeDMI+CNrGpyhLB0teVNLbfdP4G1tTSi1ZACJnPrtIi9
ocSCVzzn+cys4NSnk0QfsxXRc15+CdOxKmJL6+z+CEFxcmXuYTPrMJ55nN/IvPdyTZqs18zsvoxu
yEEmGcqV6+QgImdrkEP7GvNQP3GjPQ8ruVPBFc6DOSbZ37WbdloCn87DFF7fkKGDM9oUwl4+Bpiv
321Bqg31mqJZcpZLPPlkWRforQx3CXE/22RVrVRqs8bxwplDuG3BoHw3b9HfD0IAumvZ9Ydnzh4a
pR6Xa+P0v3y8uNWdrItuL7HE8TAZ/5oSOULVlQzoc8IAq3hF2BxqcgDKCJUvyQQbhwrBZPOKd05X
ZjEc3joki4GS3KI7+Gb+j6OYTSEGIRd7+xn86EQPOcCF8Nc695urKo4b1BzW4hGMWFW77mQHTgu+
/1BuEdVCAq+BG3C5VtBWGyg/4oPGGArKYqWB3aAmPkhn/VVvSSbEFQv8zLiB2LimKdd7Q0izb39B
Hm4zkKoItOZtBgTcLMnmIfpR03bacxhOX/ToAZVR3+OLsSK1rB3CN6tL+mmlSav+yNUG+vwffAYZ
Lsl2vwrxnLGsqll71oJp9t+qYdCywBzWGQ4eGesBXQoenQnnbYQlh2SYDhijubIrkfpd/Q5kSSMz
9/4FMBlwyjFX9mTfyC5Dx30KDZyfKIqyIU9ep6R8lTTfUymd6Fo0ZxPkUL5XMMadpUDIX6BHB17i
+8l8D5MjBaRMzuw+vo7NutrzP3v4DY8XEUV2d7lHQfccBoRUX9Hd8icKepjktaOLsMoMd1QuMjnb
a/OBShG30CjX1riP7FYYXCA5LA9i7PgALkAuyweotxYuHSjnTC3hVM97kT5Zq61+3IBDCQ0oGDA3
Sz9UsEcUa/Zuksan78Hdur+JPyEcvKM3LzKYa5ldFrjQXQQqf46UdRahxxA0vE19PZYWUJ7EL5Co
DWpfr6pFfaSEAVNEMZwYVwlVgr+GC/HyxS3w872Nq+vuswOpoFBEQU7Q9QJ33/ElJd0stZarm14j
KTwa4lfld8TpM5DI7a70Ij+zGvWAijsHw2xP9+07+JKRzti8xh8w+Pyuj1jBY8xIF2eX68CPganb
OBoH5Y1DmOSPPcck5aA+wfln+EV0v2dgOo8DFzcnGxDlKOHq1ix7ecQXipwlnfGAg2SxjU5m9ndd
ZqDtGrYnWrYOizMHe0Har33S4D2T8GRWozWl6RZuuCViPvXU1JMdcAY8OMHl06WfV4D/cnFt26lM
sarDsTc731TrvmInz14MFwRyLgZcpYmJ9Nc6Y6PLTTGGUt+pOFcl2ks+Wh/N3sUNFyHutHLkPl1S
/VuQGW0aMR+aYeCKhmozyRV20cfi2qf/1PQsZO6qKto2/0D4t8CM0+iE0vEXw4IzU2gK/igI1mHE
A2HJMU1Cbj8JmhmRR1xF5s7WdcQkOvBMNrtdD6tReMbCdi7+C31vff4LFfaTurwEYxsoYGHfuImh
+57vyAtzCrbj0+mZhV8KFWFEKZvAtXmiVoTlfOZu7VKIyReCRuFGhMiR4uRn1XFk3Ck16c++QYPU
tGa+bfVq7+R4mQbW+TNmV66OgwxzvHAycxS9+FhvmFEDNJ/us9jdAdW11tOGykavrlApPkhTyjX8
kY0CP/FzB8V5HiqvAIPKWC7rO5RCKfbuuP2lz9RsGwQncRE2n59w18I6JW1/+HPWWswkZC4l673U
GPHfPkAeejJmG+PA1fThmW9tjjApaRmr5Yzmup1EFID+1VuU5CAVg79WVCkKNVJA5gFWdYvlKFB/
YgDB0+LLXATnuHxS4njdeftq81+AcPDi5zE/BIQVmyzCpQrFisEUzdpiUei4JeZfAJjQsBDDC8Hl
LdMvB7xhq/6HLfhD99qBAyynIWcQggQobLBQhfZ6J9+CQ/RbotFL0AyRQIzKGimeajjW6pAPnKuf
8ikbKQUL5A1lq3HXz73xX9TmGK1dsL9x5FXea2RFBySV5VNTSbyodwUE37Erq1Cqin2G+25bOrM6
M3nsem2wxsQEFPZPWEJsUnF5g4VQ+AsGj0XnBxuLZLIvPDXtRjgC5Ni7WplvmficvlVRJaA5kaef
hvK3o22wI9F8KIYTsyY0jjhAUkrqsYs7bMnICfgEHtaROXfYkSBREfKXyue9buOzDoCuIWKAXQA/
mofUMeRcvNtfMSPpp4BEc4dwFCqTPhPA05JEj/tFPM+GloLrqH/MWEiJRHMk7AkzekYzWm20FJpv
BUeqWfUdFRsxP55FlPEriXdTaCNBCXAwK1Sm16YBBeD3FHFQdRDm+tU0u5uaQ3/fzaUAsimdQTY3
m3oD4QXPVaJndtSKMMiFovi+x+QLbkaRejZfSHZdRabLYtHcfAnzJgcVKm+R2bOwFj4NK2Zu0MYl
bK+xF8OSfkeUWi6FF8YaazH/oml0vDW7HbUmQ57DOsRQC+aFuuMtOOXGNhF2pR1GNAD/divTgZiJ
jcW1FSGymVxENcZ8599/i4R3Yi0hK+4T9wAVgMc7VvMU5aaVQgcOoHlkf3tTqnHudiNDGHYQOh8O
VMZyM1BwY7/Fua2yGhwl/d5eXePgrfCOReyK7wgGwM9fPZeskA+RYJJph0oqB+ifv0StKlPEnhx/
GsiAHz6vTtean9WQDuQpiCIYUbkv6GlEYNT6XNzYiPjtZjwO8SwnWdIM+iVNSAW7RJahli77mw0z
/023d9556pL0780O1OtrOHP6GRqHa4zyypH5Uhmh362gU5ILxd389jW/8VVXSsAdNfBmlBqioE5k
KgVYvItv015R6G3L0w01t1RPZHmgZegs6ETzuDcojoMZkwSXtpnqLme0GUxcO300eVpLdNZIqQOy
9/xcgp9H8N72a642G2sv8TEaOiuHMAy26v6/JoaC8fQMESh44daRnGfPi3C0MOxJqY29IgYMCTVV
bKjjnfBGG4Tzl4VRIQecv158Wq5TJ+8R46vh/xJqEv5szDgD4sYpG9/1myHZFTierMCLimjTOnie
IdXKGc1NdsTuDw/BSLWxhGwONYywTk1eslPk9C6R3ASl0dy2pwFX46R1Z+HlwPFd+CpWhHYnd6UH
CGkJ5BNAhgkbP+etojXOmNmz21aZJoaIKRd26wLW4o3/6+UJDcJ/jUVBCT7Rf8dj7wahb0Xytk10
/Jblo522VSgmnzx6f9qQyxZUjAE+Ut75lQ5J5ggZkcHR32fEYFpryYioTsEL0elSj46xN1xxsuP+
5E6q8LWr2hqfuUkkQgeavT/sZImDXPS56OAaJQAMi4zhbFXfgiqDkOCG66L+HgC/4kX+uTJK9nn4
MHsmcW50mRRiyzA6LcIsL5FrffevemMmRR9NhFwTG3ye+1akm/WjJDlK98y5ciFr+7WRaVhWBKn8
gQ/0HZVimi2ees4wKHRpq+gHIkhTESKvIWQUYkXQnKr/cMe1iBs7gQwlADVs+1idzdCxXztZjzfP
FJOcax3K+jsmXizqicRrRMqRLREStxGCs1aZXtz2bevCz6siMc1+GNmY4JwFU9Ae6xL1aJjNaOW1
1cdKDK0oV/OJ8LmGqLfhg59iZld8hPg9dPAUIOiXzJVnUkGJL/c21Saf5jnIs7pfi7icGzVnMB22
C9XcLupnFYQTnJ/K6keeViWheEPqi3mKreCc1niKH/+JI7tvZxJaLlN2SA1GIL/o+90+7RcjesRT
gLCEt5m51mLRDihpZyOkWhzgP6R7xKWtj3D1IEJ6x8dZkC8jv1fDCZQATVNG/mrhZOJJGTNU+2H+
iOTNafBcjXmcKk0Z+gzm5Ov3f550ux8LONwuE0MfXdnXuA5oVEkUGpdVKfJT4zSdSe9bvto7nwLQ
FQxgoVIQgB6044q0nj6Hb5xJXc3rESH04m3+o5t79cwwW4mRVOzwHQrEmcIZkb/R+1d2nL3DLphU
IKOh0euijcKWOLrOTdOv4LpUj1AXsvLDR9OK/lC+Me6D7m5BoGjpXtnrKbek53j/ydxayAHYJYtT
zbJgchDA0jgw+fWhYncQXukRfEbAr/hr6clrD9pGFr9NMpecSCNAnJ8fq8cE+Mojt0IzkWBK7zoz
46YObzdJxEHveHVh6iSD1A3mQBYrwkRnxbPpjB9hH7VZLnS8hqadKM13KHVXtRCAWeICIGTP6NPt
FSc5JkB4IQPXPqPcJfj7he6KivRvOFG54ZX+N7nF7sCRuNJYU6YlxeBBNuuCRGLf4KVSpDyRbdZ5
CASwEWgegEPtvJNR2n/MyQ9IcCd//KndBB+n1OHqXs896RSYGrQATBBzoNWbi1/vrgHACHBiCk6L
J7i6DOU1KuWjenjxEhonX2/sg0eUyp/A7dKgzr5VR50Xaeo4oD1Exlt+1gDsoXtpsn5bNr1NWnsy
qDzQM+vZgBJB3H1BtSb/HrwxJv/zoSjgHa0hSUHwLZmbryECAF8aBfbXC2mP+kUet9eC/E1eSoCb
DZ9XrfXLqAsMw5TKUXgJzSluVPftYfJjp9GQmUc20CO/ZKWJDHbUkFPaYJt/aL+Jc/prNVXzXDCb
YHE4mlrJ5O5XKe7n2V/Xq9ARri/cJ/s6puMjQ2aiewxmAC9ocHZYea0FyGUjPvINkUB0KkiJjAmY
o7oRt/Oi+k8BzGMTpraJvYJdxTGkrXFE8o4J+tO0IvigeH48srkVOBej3uIM7l3r/mjb8vD+iMQw
ZgcXC48xQ0uxVd2XbL+vZOlPU1FH37rCq/cjI0iwGPsLcFDsbrpsmLRLkUQgbnBB8hGH0TL39kFM
FsVDeuftMDXTY+G+6jQ+2pyZ0NKmOZp5bsYkM1AG0roJCrPp3u34xrFExrSlPqTEqwpztUpaIAXo
Rym17pUoY6iCdj/EZ6t5BqySEXlGlSewUpiannz7nGYG/mlNKoAD6HoHY8Hf1mPDO4oVrrOWA9Y1
gk84XZIq5SxgDCyXeGcNUYyN+LjRNPGB9A8nUwfi4oKYeg7c3eFcurNoOTq+3/gOrvHT2ag1PDwT
HslN1BVhbIVyewcu8pz2JKyu+dZAPMaGGlzTC1e1UjMtaB+NKSykaLhwd0rS5aJ05Sgl/sncCI0Z
he0fT+Tt7if+9phASQ2hmX0HgiwF7cFrx232mJa/eP97O7JXbD2zJ4NWUVa5QekFqeFQapPcRpFg
BFPbJYjU/sxqjJSRA2Lhr0I3VRhniBmyC9dRNtYz67nsfLuIG/3RVlNBQVmd09NWb/zePcezxmRV
o1FnFtjY/7m8kQL8jFyWanprnFDPkxsjOFqDViaTZOc9Ksg39lF4Qz4ak8ozhIIkLRou/WHKv6DY
FM+LnFRz9vFfSvm7Oov3CmHfT/s0vSkrBIBe/TZkIZXcIXH7xibvPCARrAUqUzGB6rmMIvpdki6d
YksULzz57EmsGiOKDNPymCoFcXjGxYnlpoUU8gBEfpysd8iuKv9xjI+3TNkwacRnGmcigDXef36g
n0e5am6FMW+4f/9hsbqU58JqvEmu+++ybUmrAXQxMP881DFmj7BSaj7FxlIpyfUMWN4JrUS1ZqpC
cBlcCcewyC+XGmRa/jSCYnKpQEvm4bBKF/OqJOxBd9QnqGzLUw/88bOG3SIWffd7QlbZWVND9MQO
XumAcdmjwAsK6FGIbc5dwdpEjnGO0yhUri2BUR3RpL6Anyao/BrPngi4mDSiFS9QEiUXmvwRgtiT
c4bQo9ZLD33z/Ru431z2kTGksK6lz6i8rZ5pNCnDI0lxZSomxTLA6X8zytcM4utpHSoPgXQ5Ayyh
I5XO849TQXD9ki0QRb90UQM0/xTlmYQPveuMcbUxMnvxGasdqsOKFUU7kY7h/nI4h9nGxm/x9sL0
VTtFlspcuJOBOlaME4fuY/JIMgZtEXcrhFejtMkRJauyFl/igOnj0JoiooCjVmdXyVCl9RsgTcNm
SvyzOlfC1Bn25XzMrhGg+KqnMJwmvNnFBKyPvTPjyG4j68evYMa9dC1gvg2DopB32DrROeEPB+gM
0CO95x+ywcaDVi6WqN/bqWDxrp5RTl5/oJwmao/vpclGlY5ZqGON9o17i7CgEWYgO+nJQnmTp6V1
zTJQ3sV5natcIjYRkvImp3yFkPxfKfIzHeDcRYr/ZcFxr88FR4pzSH340R+bDCSEAEmRDuS9CZ/V
gvzqq8awcJV3AypGXTBIy7bdekL/1TaEuLUNWzkCguM9DGvka2JrQ3DD8LKqXn/t9l86TPL7a7y1
ypctL8ySHk93+zzNTJw6ZyfAca/iYrPZI4dloYUyGGgvrgCKdSWefk8fxuq/GGY8s8rT9R+VcXKN
WxyduNIyGVRh+SyMeK7iwn6gv0rwFPG0YtmqPTlVSpRi6N8kryqyyuIJlOIJDyNuugcsE/mhzTJB
lZAuo3arouT7jZASnuWu1aLMp400tzrRJ/eyHPnL/rx1Fr5PkdhWh9BkEBA0O1ATz3GxJtIjgVnR
OEFa7DcNBZ6m+QC3ia8QUFWEUAjsyt7/iLmR/uAaozEQ/IAHEQo5QwDr+wY5fw5mRTptwBaBRh/b
h1m70vvpahDg6NK6wrHNW1kAvF0U9BtKgDV0kA7ktpPCj4D6Bzv/jI8RMs7D8+27DaLxzkrs4+6Y
UsY/8xeMyn88TM4H/LLr5G4josF8lC2taICo9GjTFIIAR9Cdl3qMz7I1xrNqxQpP5dsG5w9nv2pR
akDhaF/wgyMylqVgmNZseyQwOKyvYb5sojnx316xUVAlTJgO8TV4j00n3B2YuP5jU+6ig+mWfGRF
DOERGWFpF74C/wlVwsEkUnhxU9q4x3CLwja7u7lisvrbKzwYZDoQpq1Ph6bekjyqpGZOY3gRBc0D
r4rUzg+Ld9PrI5ZBYcyLOpbCYq6AJL9gKEB+irrOyB7yYDhB+09wh9ORt1RigV9sRD4fahfh5tpK
as1CHjpGaH63hQSEM9jhaKDRbh3kzG1C8z0ax92A4NfvAUqb/oZjfJ2vUYDW7Bu4O4G9k0eotsji
KnCQ4T+OEArwCwEZ8Aqc3XqPeE1SKmi/CkgWnhzK4Fi6I3N2mL+kUGYJoYk0Hv8ijw7NuRx/xzy3
sGp3AgI6FRpTLbgVHyQr6WOcoOOxBJdHlUJpbiJtp/BqN5JxCi7MJeWjKsfszmroSr6Cg6+MZWqd
iIg2Vhg6cQOLCcZ1ZWoj6NQQDNQJKtx7iqKgvLqq8kzo0KkH4k3KHeAhwVwqFM6RGdkswzzSJ1t3
dUfeVyXvVC9hbPCvvkZ1oGeMcs/ArZEre6OyPveJSAyw7s0miGwEogoC3maybENdt2khna0caXNx
GvvlYql+ahpWLqdH5Pdfy8t21Zm7ziTE0I5/trx4ZjSI6beCgbkDinroRLwlVjfY3378yG1AYpK7
yfvBnZfN18mK4V4Q+Rjan0ia2tc/L70kl2kDziLIltuPD2+HPvLD5+hAmovOpBbqsInMqL/DPuCp
Wqpyq54Bujl/xq5ljjkI/yMSQAiTtSPb0C1tFlFE1+IKbGRkfVBOH1r77Z8I8n05WL47IymXv4CQ
mlzP1hL9qkBecE9+aYqtkPFPe9hWAIAtfNWV66FT1iginWD1ANTaDWv6iqt3iAIII8Egf822qjGf
dvOtHDO90BEyIXg6V4/5zPJbyx6AT25hhHT1dhWbEwgqG7YPs7IGrSL2JmOPxgsHBu3G6zjLHFCj
rfAn4V4IiK0jp31xpWLGuZpT04yFyhNU+QUGVErENkHdZRdgwOXyQ9muMgICNHRtV+proT0g/Dy8
cYuDcgUkHdqqzW9kzTUjajE5XQr2j8g9ROvL30pB2FHaUVCeLRgMq1uxVq2vW/7W9+KGhKJUyM82
DeWorvy6VGc1NHvT1GwGXZumZHWsrXOuZuLA4UnzsM4TCeeHHSPlrQCmmHQmEYvsuJFWQrMdxFtA
KYjQkYycMj9oGUHTj/aIBEfIUaXBiQMeGSH5LHF6NwwiMtmpfVcrD/NrmWINBpjv7iJ4OxCbc9Vm
BhUqPD96ZTR5OA6rJsQMOK1VHT1yxoqzPOU09eWUuIrC74zTFsvVN554Vk18aawCZQplYV3vthZM
svL1k6Gey8Q5N5FZKfpCphqHd+iGXWuwDM37iBavvdBnOCaenCJMrjYcGMUE2jTYc//lvim3SQM1
n1box27+RHUo3JQf+rCy+ku5SanDNV+bLtpXHHqyzS05xrePQDsUobm8P0gJYx5hP2FmkSwtyPEv
I05OgX2sTm6d0IzCuc+ukm15cTx1G9oE+2UypJVEnu3axCnk8DOF9IhOzIwTPV0+2zgwU/Y1sx2W
Flz1bvGqTcG0Y7bMY61Bxqg89AnPj5faNpsfOPdPUmV/hcKmnWz8Ivq9FO04BFnr5hwKqekg6q2V
3bzgxkVqT0cKYe/fkKDKZoP5TpTS5uba56WlWuDzaDc0GBI+aCLI8rsZjMXmh+SJ9TxvtfVQBt5l
84nzrViMjwDfdnDGNZwE8urzcBItBpaWqvHL7QYbiXM9JAGQiHIPtJhXIUiWjqW0Ppl6wWb1OEgD
EM4B3y0wXXsnWEllWlSRky2T1IuQybE/4sL7Ki3nGONAUwhIewDID5rW0KvoHOrlRhgc9aK+vP56
cMuEPNDEoXH9Opr47t3H8BZXi6683yCscwkNWGat7pbmMtrfKfDQCd9/7xYVqgUmkJAShAVv1Nsc
xej2gXIE231FV2ajtQWNSWxOqWnPEykS9aUmAJ5fTRkf24Ui1bTnb6whAP5PJugVvKgpbRaPC+qk
BMWmS/PxqpP87MZiY00eNoFPOivHN381SwZlOoMYKb4g/h3bxT82Fokd1/cSBFOxBBoJxIcEniqZ
MeIxJEu0YZV2sFmMPf4PEX3SF+yn+na3pcQV1YZMux0HCm1M5xPITct8Aaz5XTmPnWDGkbhVrbM3
aBtRGHkMSipOgIVm38N3QddPRmkKhNTOnhatGQaeP0RyPUn7dTaBsqcYwPCELSzCiT8DKxjEMh/B
mtHWs3bEL6O+oxhFQR4/NjHEpYzrtORsZe/Ou3H0i9veap6UqDceCAcsM8zn/WgCSEC7rGvMMXYp
v17sBOaX+T8LbaP22pqg4JuXK7NcaGp73b/aOQvLe228NgUhFDlAr5lvJr3F4vAwOPoUzVPwUCMz
DrU3yArbXXOXZ6PttF7vnCg5jTKSuKbge1ycUSVDf4faQ752gyh3ovG6MHVqPaOtWsb7S+UbHP2e
83fm9HRXnCu9c7yjnZmDn8WEVwQT0Lhy/U3uMBamkKywkPJS74fqMHmZecfbTYbUyZnGf8+xUm7y
iDdWTFNMCQ4T6Q5xUy6vg1DuCiNa1DQo2vmueB8EBZJ6DhoFXJHSxcI+4R7Ixqj2Frhwq9tzPRGs
sF+2YX5z6ljPftWm9kpuaM6/YTgZNiACqIkQdHShZXkuyqOCNa93adYfmq/5cjU8pDK3cXKbGp2O
CW7H7Fn+Jywg+iM86xgS43EXQd6XIck3vN+rXzAr08FxHF7sjKdWOtDC/+G72Sa5eUuz7bBvNrQg
PHM1a1FkNRGRBGpuyo0gKG3kwWh3wAv44dcH7frwYovbDIvCchJ/AeGTRvwYsHJj1M7zxFCy5LKK
jlZ1ZDif/mCxxD6/BB2UGVxHwel1Ng/RcF7G5YDKG4UR8m5aqzeYszhkPyBkZLKZNV6EQWZMfpvS
2gfdkZJM3WX5OE3c3phlvWc5xlCJ3XL5/ueiVzK9bM78IlIdhj9Gx1994sstCy0WqPwQPKvKSlYf
+DWeDUeaEQ+6E8JsQO0Q3kChA/D/hUksWZfjybl5Z6bjDjZbxXAbMjsyCM3nA7B9ZlcE8OIQd3Go
tpgrThcZ1AcCMuYNIatzLuxbFWdI3g+PREfO4m1Gvv7GPPKb/4McUBWTQOPaqU4ESNAq47a1DIdq
37Xn1ct19aammIPvc3S4HicWE092hY1nsy08uZeZ7+B4dMWIeZ4VnEmy+wvu+6RX+5+42fldMbOs
UjJUOpxWI5SPdF3Tq3Y0EbiZ2bx88Gu2ByVOJDdSrX9lTWXoSASB2l4Q1bSoGbg26fzm8KM9NVj1
K9CrMGy8Ml5eeC2RUeTI8sORVdiHKwcWCPKYkqF8QG24NhauVyHsG8TMMxI01Ah57P0Zi4o/+AcR
mQslwXGWedxcPHjayxPSbNuWnUkYm5b7F61vpPyerD0eChaDLipWx6D3OD/i3A5y+mC8tGxvXI9W
DZfoYRvI3BlyepRIjFae2OvMkIPmx2FIZ2uMUgflC6Lw+FHBNfkFRyuvkspV+Qso5kOgahyyYFY9
ysCBFHwMsZWZ9jrBOKek09gPCjTuhP2HLWW0h3i2PlsfcrfJSpR5LaV9NttaYVk5moYmelRUbwXD
cXtx42dSRg9Rk8mOlI/jvllGwls305wSKFmDKabe9YyKP10iFjBl8SVo6SHmP5ycw+s8q6MGoFsC
ANv+TH+xq6XAKEHKMFCYFkbaHWR7KMUFUh4WJNF0moPwYYlGnvt8yzEkIgXSB2+DwJxg3GgI0tAr
iANM56cEgk9D/hbdSDYz2rhiD0OkNmtgNYT/ZWWIoO0LZ9KsDc78jN1+JQYayGAfFO0T3u8Dwjz8
YNNsQ+y+6YaLW9yujOsHI/KNKSdgUkzn/m1MFvd5T1Q4A8wd5ysb94ayJf5yzb5RwhJmj82sXbSf
UygiQW7GhFhLVZlXFZowf5p7Q6AWTyJZVm5LbbEMRHhJLF+EtB+GSgkI0bM+kyO4cJ8s+pl/cmGg
ZUxQduSZdMKKfoRBv2UEBMJk6SzeUG8BfDMD2p6tXl9lg9C0TqMDAvBqgBra6KLOKRWeRD2g4jEx
q0tSAqqcmTorkQoFjuxomvh0QeqHD+NzCzk+UkMTDn2gQ/C12uA5kngiVU7kxa2nbd4iYdCJ/MzQ
lfxLWBuncquuiPYjrc7l/U2tk8xvab0B1Nip/rw5CWagjZksO2S2DjaVXRoNn75ySIRcWCnk4Kka
f4yytTng4lrDTR6Oc3jfu9XpA93poc2AwYUfAEwO1jkz/JEyle53FdWIvreeiWUQBNHIjA4elU1+
8h6bbMGj5Jq7Mo7TgQr3qrHIkLOr4zna7M6QA4uW1GUrUwphrzlUQeo0OWLrMcE+9CDnUM+wMeVG
cXDtTD2TmT5NsxCHkqQwmLsbgU8eB+sgHVHFYx0B3A+Qj8MlxdcCY2g98ydmIRsKJt03tmhrLqOm
xO52Qmct48QsuWs9GH9syZKk+v8bjXbN4XnsUqgPTGKwsgyltv6JaZseOcYgJ5scog1JehcUGO9i
GZRHjjHbvrVoAWNL0pVTpXl6D5CzD2xVo6jvLXJ10cdW4ns0AT5dS0+N8tXdZz0uvbK+eFF1g1nr
guPdWpTgPDIyBqfv0ogjrUhyYW2M8Ounj1TGW0d4V+Bl2mV6eQBWHn9k8za2e2NwQlp/J4ZVwt7u
Kof2b5fkry7gE1fYJV2DohwxaS36ajYAtGBuY3d+T0v6aFie4Se0sYLamy92s8HcMxL/x1/JHmu6
og2u2J8r0KTQ4GeiGPOK3G7X35ipYQ9h9RZ3U/pRdXMcoGbZcqtqrej0R6EqtRJ1rtirrSuG0AE/
hbv2CqyI9g4BOastspn1UBSjE5wyi76laONefDTgImo+NQzcV2XL5f+TlKl5OrzBwzQgjEGCDTT4
lbrpuWab7cy1Rkxg/cDWzLIx6b/gqIjD+0QRq/5s4cVcZ/IhbXTTahedBrT+ZvABWAMQAO1/xnIx
faZBVdrL7n/7PZAj2ZQUZ6TTS0c1h2ECSYzHIj073/nECKBVqZsb7k6m9Knncr5HqaPcykOjP2F3
0Hcb3keVg6k+VlnXMGsf6JqzHno6jEA5lckBpLuoQ349/ryArH8vD4e3Z/wYbJ/CoZjwxl4RgqmG
3Uk8VDsnLgkkqOkc3XkXjeatEwjV8dhilZqVfrPG8tJR6E8gYeVeji2FT3MeB9hd8vLqX1tY33TK
Xem0rElJJkxstqEZ/74kMIVOR4IrOOXNUEaTcJt6Z2HEoJU+kAhoYjDl4PYyAv6zpcur1FH1vxRw
bhRZgOJKpOzsa4Rv19xfbXsJHFR1wWCDSzKajKAolnW0+nLlBmBDsCEdyDmMSGX4revzDmq0exP9
k7Pd+dsKPyCQUA4YyI6PwuNeYj9WGyeytaluId3uTrGXLYOB3xx0PywLqSjUXN7+vQsnoTG6Acab
7rkoWNfbG3t09e1Xm7XT05UG/xboKg5oqnY98bMP/JL/QcnYdP8BFa1Hby78H7aEHZ9SseGGLsXF
/Cn5QcKVi8WRfste9RyANGVhpvSm3vProcbJXXu5Fq5WsjLP2b7fkeQ+ekUA4cwh+LhvyVjjzspV
XO1SKitxJy4Habh812IozEBCKuXBMBvZ/2LFL3gviOCwauZ1dGEexiUWsrFJ3uhLMAYV1dE0X8qD
Tq9uOPKGMDfVUUAJU1bbTbqCmOVyV7PPoN2RqNpa/W61WMGljA91Nu4QtMNKZvmrs33d2PrM+9op
ZmwM7oa7vNugK2oFQ21SNZUMjA2fEJ6qSrOV2koqlJjsRXKQVKL/yh9hM9MMxd5ljLGsspArzoRJ
S2GTi5k8YRvo7E1hHmNto4ShGNgqZiWiG7UCyy2LOfLfpAmIvZ0liNvc9IyJNKuTBA64obPZEWUl
+3G7UlIxKwpKcpNVIbVPcriTqxNZrMfGIQcxfOy1cpBVjfR/4qHDrz7t4xhdrmdSZWs0ACl1Ip66
Prhysses0oKpql+aCQx6x4f5GRBwZbv0TYivgHcSH7wKFhvq6wBZG5TvHV+wMAoIGrWrCaiELPsF
sa19f4nmOkaPj3KDwBtAp6OzMfE4g+ZYSgm9dcoT0wwZRZxWC0DyVOMu5ScQHAk70Dxw26VMG38l
yxKlKnBqJV4azxZ0D9MLtcDzE/+s6E4B6lF+oLHZspXNWIbxW6B9/WX3MO/vC0vPgcaIsXUi4xxi
0xiimYDagJ4ui5FhN2Jfnu/+fmSqJkHKeuZTB824/fSPm1puJ8CGcdm62pgJiqH1qLxjRW0aMCbd
d00H4YgPO8txaqGUUP5Q7mtGoAQzMv9jicHdDp0ydjaYGewy9JGaEXwKCOpNioknHXS1uW9eZ7JK
eW5os+QSvpSPhyiXfwjVhZo5TdDHYOyc/4eZRxHJ+HsffWF1Ni6QRkE5WVlwj/PzdPNLsxi7vfTl
EguuMKwU2D7LPXLKVQojsOOG+WJ91wokJQQ1vWpGcnzzYAhzFT4OgA8vcujK35RmgZQuVOZEcULb
YS8Mx/caft6Vc2Ts2ISYsq2qcZxNobDtlkCIhcfv9foQUHd/eewIlsZu2GKi5XqWWNeKbBKbiyQf
Y5lj+La/rXQfJ6nfRyyyEwfTokBtd6NvePVxT7DM6ROGRyex+WTu1qgjTPz7WTG8AjjiMMOP46VE
VTZeNggNViNGq3jRutstHaUKbtWR/eZHLUkvFmg7NDSH4UpGz8uK2mohJaIWhFEGr16eyQciZfLl
5EpsLR2KKJHenh37BfxtanImTO1EJFLl9oX1uhh2FHNjWj/Nq1n1qDVZW9sddWIoYPvZO24jWvNi
nrzzzjzpME+cR24RuHATYV/4pXB+hvv4zxW1rfmNVqvhnLnws6OHvgvLTQ/UHh18mIiP6VHbRbIw
yWAUxACcvO2T3UBHBXOJ3pp/g496Q+m4xCxymNJLTlFfRHYNOQBhCCDz58+EObaN/nnzZy7xVUYT
1hwWbdPPJvM5zfAxoGI7MZPggjHiiRmJm7u83a4btSWuBD6oCjJku1b66zlVZBm87v+ELye1+M82
LvOz6TpFbcnh+qT7q1wMk7gTGmXTM4trlVOXS5MlS7nFBiFgF+kqSM+DDR3wQjLVEBUcfnsHcMWP
Ef5HX5x9eYqtYf5mufdz6nbrwh4HctkNvKdZEenp0amQ+Rul5skwXYQabMQizodHiU48mWQRRnY5
TTynNVuOsrxGayh4OhINPJufIJKjy2XuQWGQcxlbJdnMvH6K0LUA8MAWBO0gp0TsL6aJBy2UC+A0
rZQbXE7uywdvLU5JejYTaDWcG+i3226vBapghOdMHYmX8YZxgQPSsQkl9GjOHnW97pU2LOA3Pe5T
zUGgJWmJRiIQutwXqyl+oDK9TQbJMKYki4d4XYh5hL6p1vdtQzaHHzuYXJcBeHe9Kcol8ILooNjM
0Ou1hviP5TlE1q/zqYCmGbmeeeyIhv07l9yCDEwqpQYbg5gWjK/+X84q6oyOgUftXXa47LW5gdNJ
S8j0up73+kfDfei5LM3o6pny8u6xYnWF93YSZB1lDYnO8Vc4PGoZgBuESwe62EGWrEU2Whm+QzFs
ThSIh4v91a6v/JAc+Ve4R9ulNk00J5spMKb6BSlemDd7l3UQaynFlyyEcdNmRChIAMSpYyjgAvMr
Gmh481ixiCrF/Ngqz0zK8hkPnIPNG1KaNEq/w0r+KlGeYp7m9IjIKYLtFFHU2eQ61UeW2rqLknFI
HYMbHWScCs/TdXn8iZQmj1Cbh59fIeN7ERm/vqJffQhPbr/ImXnb3hbvCQR5NEMcO1OWzA7sqZfy
tXWp64jJV9Fz4e5wEFmqu+ow8LCgJ0kgJQ+jCN/JDhbsr+9NL03lOBVlwNORFjJNcRlgGCA9f09d
kVK4wCinSSRbEihnJ8iowHZJrUcCGyfWTyrYLc8jZbKb1N3JCZZ1g53T2A6FXR6Sv13mKJ6DfqKm
H7jP2FsxmQ8WlamPM+cRE6dhn8Yoaw5iJN8ymX3soamvLoxosZUuntdA2oOmHYp5qgkjO37aq6r1
Uk/mVcuHXmXp0E1heJPMfNQoFbkaZmkzItPFRZFJ6KGfqRNBeXJaxUbU/fAN3SJw8MShZ8qB4Gwe
qo7iqbfeGsvEtmZ3uY1QgivlPK9+VSZnmKRUGl/yPduXcBk0YDfEsuhD2lo3ZO8HfxglF87Qs6lz
ptx62JRgCSu2P4Fxe4AcowByPLL/xcS64PNdtJvLNdEjXIrPIXtfQu9KwAPUu4fOdNTRXV5vjDFv
1fw1MmPD3o/+ahcapxllYCbBKX760yIW4HT1CJghKGFY6NrwFsoVP5X7epJIcwFBLQkPVrMXEkR8
Mi5bOK8b3FGncBrNhFFnKkOyVxbHVOYbT/nBA6HZq5h28rA5i1+ASG6szek0ijqqum7VFo00M6X1
/Uq+3ptNES3A0LQsHJzZEs7jZbeYHSyzy0RRLTvTr6osoLSec8ElmYRRPIoTXQWds2cHd/p+xBcW
YMTAjfljjJ5Xrh+Ly5q+figV3kaivYgBqRnwCRO9l14N2ueSG0TinS0fdmFlwvKfxcDqpraIbLbF
VxApAVb3BPU4LKHZgeJhBZexHL3NfOI1Zi5doTqBv5SGdGe4ydJf8GcWifrFHTUjuHUYNiF2VmRd
ueMkVb8fywvkzj86VuA4bBSA+wyqFPQ66EOiZGwl6p/Dzhl7SW5M7gr04KCOQEGQkSNfRg4s3D5E
6jB9/+/7H+dtJe9Bct7be2dMNLa4kIvFN6pdBqOo7PgPO+hsqlfzJXCq7Pkx73vvu1GgiABqNyXT
Li9KTrYchjX7awyQVa0KBVvUIPuLDFjHlZN+BNmWxnFzgUmFkPhNmresrz1EKkCl3Sjve7umFVBq
sxTY4GZIkdwCa8BUE4XHSmc1UFReVUER32By5GNRz5fYUsSiS7nozRECwadAUvbUTL8D9toc5F4V
Eyy8hLv7Kf9XVCZf4TROB1NybcbbBcR8qBgOfTyVxzVGOMwyzUue97hCsELifvDSUPBBQpxNrbrY
y3DQo3w4BuqSg/28iA9XkWIVBRGhMIDdsRH2ZuvKR3lffaUfAC3pygqv996NxzB5qqVuqp4WngkX
K51e2gu1z8AO6dL/nwGllJUf9CosnsW9rQ1DWr5E4ZefykPURqUeruftHIY+/jX2nj277gclj65S
WSiFsXb/0jmQ4U6Bkd1QF3vcqYZjD4HMPfdWm7njGPtkrJy4YMbVrt3R1+2zzIQb1HI613pHqm2p
5iHaZxyLHtq/eMn7rTm0P/f8dzIMywV9Zoa8fOi31ivwBzdOyEuigSPZ1cF2eZrnI2g3tlMan68Y
yLEtD26Dv7X3uMUQx5pFaut0fO/4IvliaVPZZ0j9s3KWZJPm0RgMV1JM8C3Rf0QVrWUFoTxX28V3
6y97fjeWOn/gADVUwLViOafufRhj9oDDuXCNJ+hIlfxf5/40XuedSmGYVdmqhJvW3xjFzlxgk4zs
vq/8FX/yTAbgPKfk+0WgVCVUZmREs+mM0ykC0TP6MZGSkLveScVemcH99uQiqAClThe9P7UiYn8E
LiWHMMzaz8bPJAs1+25RxTClP+toBJOMYgInBveXZnFC1aalQ/wIskK+ONdelyEVZj2V3HtXBwJK
Jdzchq6mcHRuPHVfnsGEnCYjntN5H3AsUvDshLHi5VQa7m9/B8x+wYmCj1KA4hU71c7SzdWHAoLt
0Chjx+vsx0EZfdGc9PuXB52RTuJI5o8Jlg9eoocdMTTnEc8XTigRrwAFNHXAA9buhx27nz69f7W6
E6mrQfYUhu68eFunOETfilQl8bleMcLPbMmSMlKimgCxhPhZ4sHRckHeHs6/c9I0ya29FPMqyxL0
UI8SYG5dt7uS/XcoUQHcS2DRrtZUYrPVeszXIu00z4X4UfCNIhi4L+uPz4KYOIrWLIqNQJcMMhFk
9lmoi//KppSSndaRVGYvcnmEn4Fs6RyAXTuaaklvgGzrG5W8Ri3PzFgAHeL8aYf53wwWWUvfeMlj
X/u2AZXYDfs22laYmKf/k/6wHb43HNNZNb56v6E2OnIt/w67BdsgOSFqIZBmPIoQjqsRb6votfEC
Kxk889H6QPUag9ArB/v+DTtJxOFOGfl3HtJP1d6RekTJfrcYX4SoTMhdr6+ztfSWJ2YQ5Fkn/Lx7
zt/kPshI0rcdjo/74jTFdcKVAUauTC29McQ7fP+XJJGfL0ldrUb2kXZ+QXikyGm1VyvBssblC/m5
HjQlT1xhEH31KufHp88mRz5kfYR7hyzyClw6MzM9qyT9x5GoTdEkmRmrIGxJ579+ukYXaxNijHHK
Rx2x3ravmJNSkLAXOflQwkadiqeEHVNy04NMwH/7FK/67E2tKceGm/aACpwVev5dapwbcYIo3O7X
PBFkzn5UZtgwNn+pRhN6ZUkbNNYcBAMPHg2TW1LVjUL3fJXNJT56nE/WdsLd10qDyyEgpxbBpbE5
Q79PmKp3cE5eu4XlD3Kdxe9vT63SFAptfvapoEyIli/GuKgQWM/u8ALTsHJiIrbUj0wBDbSF4klx
I0N0+AlvLfUMN7NGEuwy96OHscSk0h6DgbvH6zLguRCqmiHXofBZDjCPs6PZFUOW822Ul/MeGCqk
oXwzjEsQH7m384mp5pb+xs3DYk41Xq0uckjuDVVrqTHHFkmjn5/XfXh8pHY6lu4+PTGUSa3CWYP1
H2JGr9be7gZiMJecAPCGImwUKlnSdTcnFTPBw3lOp7qHecyeBAWQ/wl05YZ0aDE+TqCVEIyU+Hi+
Q4JteEAihop2NBLZMAXYtsJqKCb4PPjW2UlE0cXHLcSBvxhQA1D01+jpyeuAvkS7f9vXAlI6JZKL
dIQ/zSnNg1e9YIa29dSEuYwC45FUBgYIgYdXVGCMGrdvU5uV9U1mhAedmBlSfDGf+UIIP/+xxkLV
kYeKLlFidS+u4IZfXbQbvYtX4+Kcs2yu5gCxc65X/kJOjyTXKKpXFPWT/8O3Iwdv6fGKqz7zHq8T
1wynzK5G4wFcKJ6P7INFi9ceiby+GyvsqQi3eslz6gI1qt99wI1EorxuAAk3ipLt5QDw5X/1VICk
x4kXn6xf8Fh36+7t5UGVBMHl58TWNlDBs1CzbjMpsPiwCslznx6iUN+9LNJ3jQsVVlcU2Fz2bAYL
YNCZ/O2qHqlyJfwzK5RgcGCiyp5B6YvpUMqoM3XzxBymhHemIQK1NW9aVuHf74HinuUXHANmG//T
f/ES1c0OKnCdUPQ7i6fvFfEp03+q052Msu8tE4wdORSvkGEytuf4LPMJIAuyrLUIFPY0O+5xXuZ5
W3QUuXgIoNpTtqoVNY25leK0RpPvGkjOEod3QZh5F4Z6gPv90pvhlWfLTD6OJ0Xdt5sCgf6Bc8zE
yBsT14R7sy5cKC+TxqFSRwm7GOxycbN3gqurySvZ8tGjETr4AJQBzQyU6u4SOX48gqjSa/hjhGxp
gUKJCU77Id34v8U9mPZQGz8Y21tmWky1EsAFHGRhfeK7H1t5y5du+cYFJHmnNN3ydrD/eoujhHJm
2Y1DSV8AodSQKkZj0slCq0wskY5c5sZhK6kKul2oJF9784mH4LW3MosQEJby3Cikr+VKzD2BSxQM
KUUAqJVGfwdNyAnkbF2L6ODJUmqtUzrfS3xiah8GhyuO3U6mCVDE08/SgGMa1IOgu7vNrbdIuKo9
5/T14gNbDzBBddnRkKadem7Nz+0kn8J4KcAXTPhnio69Z/tU2hvjUACsCrxgWs6yG7sw0UtmuOOr
tJwF/bEYV4njA4r6XyYQ540Hp8xtCodS16XbjmjwsDmvaiBshMO19ZfhJTvjPqwYp1Nm+moRAzNA
aRGLzulN7mpUE3xOY7kTctigrFga3/RCnR86QIc1Y0PiaO1QPzDOxb2wD4yeraEifsk+33J7dUIf
7q1ewgw1qO5GO/Ea46f19Tbc736kzxi/qZPoGz8ZAcokh9SSK6PqzOp35POp/iIJ2ZcFWz/RIIpX
4ZmOWOb3z+QhBsrredFcafTJ5CrpKyGcxj1EaPTH3jKtrq4CNujDuwQiwtf7BAb0v260q8QrDaWV
QUpta8cA4xZpdNqZNyGLQ9v/F7i7I0/yJCX/5YUWL/gIDQTlmJy2V4hoYvlh764EfNgRHp5ibci5
Pu3+n8UKKujx3/cSajhE4rndNqdqUgrnx6Jf19dU9KbD3sjKYXcFk/dbYAhkCLru0wsSfQsXo5fb
77hYEGBUPn0HsYs+MeK2BNU/ZfEaHLULd+wMevonTq8PJVPNuqJdyPKRuOFnN+kavVGADvkKJ4aG
Kbu35Zb6ctykscNLIScI6liNmXUo52RtSaqY9THWpIdlH90YeaMwgd3ejXgKETCw6o5/sskx8oxb
ntx6Srig6nj4MYaWIS76JTx1+6ZHq1sbHUyI2nHH0bUE68rLIw1WBa4zdM6pPIqL8R4ajJw0urCE
jz3rGXzozb6gECZ/FDF+zlTOpXpJAuRjSLNUXdxU4LO9D61bsG7BlBt5+YfTs1LsvFrK5Mznn3dz
soSMAweEYbOhLNWiJtmQhet1VVX+KBBDf1AziudH5JjXcBeoCHGi8usJ5KtxJWnWdEF3cpZKpAEu
IJZl36aBRQSZPqersAxAdusD1CFiOD62ohWc4T56aiHlW94SRErf8C3tYtL6ndtPGFqdl+rpQ9Po
eomi91pS021VhcxH3hVT/iAh4/31oiGbEEGN2Jm94byznM3SnqoN4RM0dE0dOQWu0+JgJF4aJNEH
MLO/LUPuH5sk6vRsGG15NHixjZtPQCzXgWvwJfUfCwXGhWZNvWkHfSzY8JAoYwZhbzaJstQdj6M9
kLV2+R7b8Zi3V7b/Qb+a4g0BjKlZD3ijcdELhkm7hb8SXuv2L3tQaRfxSJnyjNhRTkfedyHtueH1
GSQg4o0wFc2T/OPggEUEgahRZxzjv+j3eii18lJOmtjnbKgnKfQxZX1o/6SGJCJ05mgBMDlXzYiR
CwfpIqTfmIfmBAtooQBniguL+QFT/24UjNjXfsRv8XUqhxUCjXO2QdNXlsvQhVZlMb9upV7XjYnL
MDTJL9ECip0b5o4Lndm8CVPabW7uc2ID3HJ4LRaorFJXTOFbx2zxcT2ALYi23RqHFZnPFfXwZ9a5
a0xhUAyB+ClpLhimBMsilyUOkZnqJ47pX+AGRBjwhEKFHivLx6bA+eTJYUOf3o5YIDKoiDeJUVTI
NQQerHmxDkzPeIg4LKV5Os7BgmhF3KhNKLlJubCL3CyEGsE/E96OyHr2HHiR93B5Rxe10fgVobPw
jnTQ/BEC7GL0U64P6GSd9CSLqnmZssJ98ti/RK1WiXkFN5B9Ca9U5NmtyHpIxoJYi7eTk/LRtRTM
w+ibR2ewMYaMvftZppYC/tRrueN79ywUJTsSaUyiAuX7am1cIk2H3fX2+t9dTbx/cj45cLznYOP1
dFgjhkst1vlIxIVFfMvRAlFdJG+8qKtAve0ybKYinMqGJ5c8kwWgR44DwtqJQr2VjUS+IRH9ogXM
Pb26fPDFz6D6S322zLgH9BEEOP28H2dnnCXn+npH0itoJVTmQCVMX+/tGQBzvW2UDw1ExzhBQs6B
LQn2az+zirvRwTgCqyB/K5jh58ZN8k4ivn3dxSxO96xlkhhCceQHj3We6lKMo7Nn9FDfY3qevu+5
kje2jRainx9MAWumnBukvIEOpxt/lH1Mo3PYhk6b/3xyTkJq0mp7HsqAZAu3oGtJxOTCdeyAVsiS
dynQHxBV0gg5mayHKCO2JZBDfRUOeXNxUFWhKH0063z5PfM2hj8HUbhyNxwpFzaUXN6T3DXDjzFk
xrNiEHAZY3MUfOabjpcw9/NXtWdRd7zIJO1QdgSQ+i0UFPkgDjaH3OQHdxLlKGXbGjftZD0ejq56
LWmGgrUy6Fw+fof8VSfII5YjaP2uW02JPFKJBJSs/3j+cOTqcVskqmRek3sbmhwSRMNa7k/Zmuzi
Lg5AefJ4Z/TafnYlbIoum13MTzrDczZzO07OpwC+f9zVRdZUVaKaa50l6+RunlHBei+phhpdSe7j
uqT8a2V95dAm5jg1xaEYHr4DCcyhXvyh1LHjPjXv7q3N9QtG4fS+pnRzoNuK5MMB4Qbc7umwKnab
1JHK7ajLam6f48+EYJjVMABCh3TskDAeMFCw/d3vfxmjHa/fbBr9VNjyXeXP2e/Q1S+G1Yq9qEfQ
Cw+r1nCyqIALvnaFsju3mA0sTvqxb0hmhR/kohxDsb7qtFaeQaDo1onjiHWXAbX5fbTtvuLLRLxs
GjlYPuBx6sFIwAMt1bgBU19v86/gYKqfKk9dyZ08QzK50RXv7CbUltg1vQOQxE0DpBlHyOkxV6zk
kWed+gLYwuU2SMzfet/Du51TH3ps65mHlzJnDIo2wvUk5+/P8Qp/8VUOsefWDPhvcEkm2BtSIM4u
xdR7OGSSYhlu2d26wtcFN3mPcvB+5wlmeQPmluQn5TnYvzTe1UalaRNmiIiyewh35sNxjZZEOe5w
5bDEqsFn/vmp1QGbFklZOf365ZbQPhA+rlKkiI3U7DaEIN57dqpxFKZESfqbGcbNeA6Doiyi3GBb
6oQhpGgV+818R1BZbB6QcY+BIrCQZKl94q93tkDL9JA8RMulbJ2fLTv/hTPfYy+umrXb51e4jETM
/2gXTCpTyg0AHs3+ZwEdJS+25YsP7kF4Cv3uJ3ml7JUHMZPLKnDUPpq0YAERiAXCN5cb499CZgqT
t1wJ3CGBmyOwP4t6oQzGPFjN4ybeJnu29LzcssoHZy93iorP4zbdWmUwyDxCn2mnJYJ0s13YRjp9
Z1WaLBQdik7Z6nBUOpEKs2XS0WYBUBEGaasrzH0ykXzgwrxFld+bMOsKgLia7PLHmBZMN88mkIxj
Nh1cmZzb2lh2XTHgxTFhrILdp+ccH8WtbxuPF8sos4KPg33RZppTk1+AJ4EmTSkmq0Wa717/MrU0
zwgdn0s9Fy+QUI3qKwch2Eb2SUZUdgCN3R2MkXPkTOTEi5UTBzXjBs9BMiIEr8tdlZ02ift4plYN
vEAEkpQFVokw84JX35PckaAmp74spzODqc/lh2Rf55wdaKpV0veU0F/ErtBaskzBNBtEMGhpraPz
5KSBGaTrVufYqTkONiv/gXEfXQI4fwakGorkikzQUeBVV3cZ0ATdyxeCGNXaDUO7r50VD+gQ1Vih
i8iLehPoVDUsj2bhfs6n84QH5aON3q487qCY8OlgMhidho+KI79WVfPwnRk1jtmh9NYD3uFnyOfT
lhZbQNZSRvvNk47Jga3+1KM15ipm6N7e/YChEWxjb9alzMXCSacDzCLbKnzclaT9lxVaE/vHPgIv
7Z76UuBAY3GVb1UWSMIIQlELgk1q3qpj3Qd2tNbYiZimzYlsFy4OILqq4zqtt01+DAetyzMYD0TF
2fjWgenQ2GX1QPv/1YKvtoucskp051HK6UZfYYOMR4TIJKsdkEfCXnRUlRI7Z4fhZz2fBg4VW9UJ
m6OPuJd1M/j/W5Pa8tuhl5i0K7wzDVZ+kTeA2idiAXg1Qhd1f+tMQcOyTRk396AxqczKhmDHe92r
fqKyzpKMnx0bw/lsQ5njEe/wEeyobmfBgJv7/8g1VtbNtZwDV9bfRWUEPrhMI4Oaqaye7N86K5H6
uFM7VKVWal003WFnOftaZRiQwCbDVmaJmoZP3IO6iTOlKKCc2wom4GCMed3jTPPxySleb2pWNLCw
tc7XMs0D7/VluPUiF3UMtuAkfwV2KZwfBfOt2Hw7Ed8VCL/rsJEdwg54Ahr5Qb0fD3g22HyFNush
S1VAM+Qy8skYbUEhSgXvvYpuXfS1iMFU1v30s6s5b1T2aARqYB94/58tf1wHDy1LIHD4PCsVp6Cc
VUlBkoksibPPpSZv1bBJHTpZ9ao69KZ+8cFvjSh8UcAvhF7E498hRLBP7nENhKw4xw9JmE0+3vNU
B2QgMDcCqfA3LOwm8KbPotMQaE9PUek0wANzPCBN2fuYfPnJmq1C83K7WMe1DhyGyRo4z1WKSQAr
myPm33PovabrJHTH+WDzy6NtZ3xse4n16Dj6p82P3WwZsjHFEm1W7XRz08Dj5jYIAFISV7tweG4v
TSEOklmFvKvlleWidr6Nga1GV4pnTA3AIFu6M5np7p8qXqupfLRlVWkLUtpdChLfvjhPE5i2SJy3
7opoy1+yplLtb1b5sEod3PnOQzCOD53oaUjBe3qkFXlY98ejla2UeocCnvuiyXkmmy75tsTwJYqG
rrvxCLJfds3pXjivDng2jHHTTQPjA3d1DmGj70o/52Hi8A1FY/AoXDNmST1j/WbJWvlpH8IQnSL8
3E8UrREg4GdK/5pCseg7rka1ou0NVIePcnktbgCQ99d0IZ8hBcrlIrUZG/V9vXyQDamK2EfCSpfv
Z0CRzAqt0GE78zXwMICc9gVauQAQil3vPuWojsjLFQOQzjo1eyqL5LPUBrVVSGTnZxtEKIOMaf0P
jo7xHsrVVbHSqm96GQmhK3Km7BQsN5/K2Js9h5E/5Yu4I9lWwIvZKy+2OStRZf27/fmxmksY53wi
xfR32xsfmD0TSauw1avhT++bTNhvHP0WWia6VnyXSpyr0oPX6odNCPsiWlIxN8Eu/z++z2NkX5i8
Qr0nsrHqsQF+U5jgCGmHieoXecw1P1tCp9pJQIIN86MA1UDuOkl1uwQMkUiOBd59jmtE88JPQZpa
VsoPyLBD7FSZdJcSTsGCUfoEzMnJ0iqHOwOfWb9FaDKpjd0119tRJz/KnfjwzWo55YgaMs3UjdB+
ezvW6vQ23N0PUdUOKzO6WS7F1s5S+amT5z860JZDs/nRb8eTYDXBqRrFQ0ZLOElTrbwSSLyADZgR
9tmxPTVyNi+96A8TdrIm4Yqvzi0WUSYnrxviJzSZMuzkBkq7OmYi8WBIqGFtfkq1b7QwuvAP6k1k
9c1uWIhfjTYIDEx/Iqe7syi/p3beisbtjt0XEdrfTEuj8MA5+aWodRR/ZymbzD9fQcqbSm8gFMzA
sNzc0fI423Wuw9nwUDZGNXAnyLch/XX99+M9iNsQjg+nKbrfEN84n5kvxkb/72K/wLCD3yM4NgKe
+tDRr2VC7k5SeoriCeuLhg2DG44sJ7jaBGjU/Bj9va8/N1BZ26EMjLjuCLSThPxRKME3oGIIhQ1B
qE3e7qRA68GXUqHNYJisl7iGBtAgArQXYMstm84hVnXIEHIAC1S/G9c8gGDdJTg2jhSnblqQZ7Fw
AQM0p1dsu/lxKoTVIRUTsvOvE+x0w4lV0HzwwRRldsrLt1jZvTyZOmOqupXT/cFLhtHyCBhgsnqq
ox1Vwe/9wA3kVNzFdP6fL1Xm+9GGk8o3JkS7oaf9Rs7DNDHRdJjqpucGeer0d6ReCypz+a1AcDO2
oOADwLCwlaBY7EE/eqZsWRziv8DXbc9XGaDUXwEah9gZ2yYfQuFMeoeo9Tk1EohZEY6NhSXkfznP
emHg5pQic2H2ueyunuzZ6iS0gWn+h5bYGEkVU9KghzE2CudRDo4xnmCjSregRQadwb34v8tAPmGn
SxR4vsaWXHIrA6PSTrXdv8JQyKr8U5yUgZAE3m889r+rWcWylEBqa9IJGzSSo1DVwYOG76XLmSVn
wswNelD29JeKujw0Ji7eXVLOJwsHZLFztgRWgIxPCeW/duoScyEWoeVohr1snvQ5XdiSR8WEyYPQ
tWTroVfofq4uTdKEDFhIhOVhqzIXWJ6cIEQc5GcgVIhLWsD7mhcfk174NjymRThOgV2F5CN56ZQ3
w5LpaCAsde7B3HjQbyFMwKz732+eLMHmB7QKUFXPwwF8RO1IVBg/68q5DIs/IMFIqaDDZgGGnZO2
+p6DB6dckXIgyLNDxQ6SrszqyJVnuu8OLcw3Ael1U26dfZtanEk/ERvVLmaZvWd1sUZLt3sB98jk
mMh2el9e2PrVB/7ngi35td0MBHtrjteI6rvfy7Sjw0e3vbrUbKWhW8rcZdzaJA7hKj8qindn5T87
a2zPMop1OhDAVuDuc+APi4n1OPnU8ENorr/YKgJi0tU5Y4gpE2B146XQtQaE01p8s98FjrRfkOXe
c+V10/MhXLTy044Qcgf79Dih6N3uqQMuHpJB8gt/sq8GjtU/+1lJ+S6zE4jUx7jfne4T3leYD+em
oeV64Dh8K8oSV8aUmAdl58awiIdfYRL5D+oOJ2wVt17EZSdvyUdOl4wM1FhArqUJUfX3orhUJjle
8Z2S93lfGMOouFNxK8fB7wx1dHTS+wsaLWFz2V1+Gq1KdauTvUdg/4Vw0la2uupDw0BdCexmk74w
wWgIsSRbRW3aidMll2l94QF1rLGL/57XJiUhaYiu+JlQoJ8carHil4hdTtyKVinXNJkv835Qy8xd
vncedoratKwQheMQCzaDnVlRT+bfsDeE1gK2ZSEZli6VlCERqo02w4WECE8EHqzZaQr63Cj1yduH
ysEJmJulvLXA1e0zc2QfS+1NmmL0fjQbhdcGrTxbx0Zgn0+CAInSGK00lFiNG+I6zlp3h+3ekz6p
LNmad+IT7POwva1wtaQyFBFjd5zFcB6SRGNOgIFD5t6Calo351QtC+AfGmUGgyFCKHQJ34E4BxaZ
jOZbeD+OI6MHbei9QV+8pN26bRiC6Ekv3T3Tk2FuGfWNEO+dVgJCWBDMNoZGtXLO/g+VkCOSLK3n
Gdc1JSQuCKKfFM/sgHjOgxmVoOr3zGYKSfpsUClY4+HSch/i3hJfQtUncG4qEdQgbcRULcA5uYWf
QsK3D5BEzujw+YLSDrmYyJLmdY0fIqKyzH2ahEvq826f+jRbS68rwOz5xQeASqsBRrGRVbJGzEfb
mf+ynjUb1VtjbaSWb5PLRijaJgYBxirXd7zDEUXkktGwgl6dluOmueomPd2e/6pFm+OhlKMAIIqd
Iqtb2XpnOLToetcoS/qXhgcokgmfBjP77qcqFpQreAlD821xtzjbjIItOSvFFjZfRieopuP8U5Wr
7WfUJpqaLiIPCnCNjgOmkGZWHO10vpPOLVoBRh1ou/VMaSV9koCj3Xgh15RIFFtXlpFmx1bWFdbg
0BYxGWCOOLjYYGt9Fk3WK6SWN9uVfye7fB7m2+VE4vxGzqFc0Z9gUruHfu7cxFwZ/fGmG3+pubhd
b2TWqbRSeihAKG3vs/8LCCGUFdlOIHWUsCicwrblM60zn9at62pHL2sQk/akHwV9g/lun0xrNz43
jymjGFdpkyij4gvpX3F7Mj+OTtlg773B7OZ2v3+D9v828KRNPdkMY1ycicUmCBDgSjqAhx7MyCgC
L5HJv2I13BvplxtRAjnay1vCKK+d6Qlhq2Nkx7FQ2D7TXZS8cLCvnnh0rYTH1U38anu470sUULfm
DLyzf4zBV5EJ6SSLylVpYdSd6tnwk58Gd9oFaXVe8iV5w2ZUtqALC6WViey8OYMxt80eAc1HS0R0
iR4MrjsN5ctN7t02dd06wm6rplDKb/WSN0xrOpLSFv8VwCsxg2Dwo3vbx2mxLdQllrlIM7S4NY8o
MoP1gHYELCtOvc8uK3UazrkpM0GbuIcW1boMRu7r0NsEwK7W6fx5aL4kam4F2sacR/qQIslI2fxQ
ZZPyNmSxzrmVqXNBBHnB4VG2E093+F0CMtkkIwMGUhyc3VHPMIvhldPEk5gij8w7oriyH2zXlwaD
Gv9raVpg6oeLm5EyjYEL9Eo+gAK9esWACbbaNz0uBCq+OMe5qCnmyENLjpe7sKxHIh5UBVGKI9Pz
CyrpR2NxRvgCnhbzPwM8q3bkX8G9xvUICNrD3FHrkiBSxxR0zNwsHoLyj9JOQOIedpxOsMfGSeMb
Pw/hGLbsKPYZ14dLU/9J3xcbphXZ7ZUEBsDid6hlNWLhHs3tJOAY/vNij/0n5d6cADoN4PvvqkXY
T4O37JXcFC9eQTwkKOwK2jCzeEZp75djZqSBIIsD/vuhYrlFL9lwANh7+3RUGIfBEpk9NyhFnovU
O7TOc1IPxYfGuTAIcjndS85v5cb2bEDrrf5mFG/aXgMzane5W3ZePGr+WzF7v1vel8QFDabN/Spd
GzysGXePTSo7rdLu8/fBvT2DmxvPQMdPAXwUg2pskiXm0aNrON42ohbo6+Hip5lKiDvm78GvI/ys
BpwZAApz/2R+xZOQYk+wfZH1ROU7AYd7o0Kpk7A6wwVhKYfX0SY5GflyrLG6nzO2ckf71SkITwS+
XB8DvQ0gH2PgiD2nhPLZmmR0gRZZCB6cL/o1fzkUyfV27uZ50Iq4dEkQTqbEpjdfTf9OHcrnlNKF
+Ax1Si0lXTSfMb7VQkqjJBA3say8qT6tP8Xgj7FoFzKZwgkb0zS9js93pYBryiKZ/zG+kWBr+zfZ
vGNMJk154TN/v548eiE0dn1euMElzF3GqH4wo/++9HKqLiRfKc+VuOdNDag3kKZPwig1BuebFotg
Q7rpjmClMzEd/3NdPc01v+R91RBlNnNH3hkF5XJOPqJgaqZag80tCUkAh8Uxaqf8LsaUiKaeQdvt
Igr+AT/iK7I7Dbx4T6u/rFdhIFJpVrhOlr1DmzlHXVjaYshFAYYcsUKULHBEiRIoQHgWOE4JxttZ
n6L7noOzs4Hu6ElyA/84zR2+8gTFeyGZ5rQ6k5yXBeg7zdPx/30cNywVjWwCFCzJD5rWqfcTmekV
fpAFY8+7SJyS2Uw36NoHw4GhrG0O3p3nlLqUdXWb+mMSzvej9wpvylmmtyY/3q5yAQs4edXHmHZC
rdStLjvHdDCr+OqzgHpawjJdfHlItwk9tQaZp8iVIIUsSTdBV6uZkppQ4+HDPZ64rWXIKfW+0nKN
sLY9dnVQpJGx8iIUBYAVcoUQAgP5LeZB/w3m1Cl55RJn0dvyhH0KeBBJNSuYd52Xq7j/wLEBhU5V
+FV9Yy/5TJrrkJLYC+gNU2GZxepebXzxo77PNAMVsZXor0wqgLRw9MRse5D4UMNpBSIjknDoClEc
KxbLbomLoEc7Hi9O9Mv9kmwqUaisq71hvGHay/GvMkpkUbfKbVjJtLWFR6ah6Gyu++r6N9jFISgt
aECVvzOhyX4DV3ENFhSi/KU9c1POeubKeIiJiVP8ZZbUzCiLgErbnq/o6gAchh55y1lTmmxB/0DL
V84dgN2cEwJqI9AMSSM/zZz/bY1F4+cxSRpFQzDg0TJ77N0JgDNscZbr4imCS8inNTz05cxe8THf
tv4F//XFTLYOZaHPhdp6e9hKr71BK1taNAPVr6VTLyVo6nnx50U78OHcSlh/M+44GvP0QUod7h9x
wyXsJLd9Ml3HkJSdB9xUB65RfuwWODISfD8+o+UGXFbCny8ZzBt8xadvQ1lckVwVDi5y5dnxUt/u
nrpk+wXmawaoL8y+08LIshb4+n6/yU/2qtGmu46vg4eFxWPvVqtfw6Le/gTQhHKtslY9PoiwyEqu
fuuq3YXK2fsK19f4sH814lCELLQ5oC3QItGkdtj3g5Mbl/AZiEUFcSi8pf+pOO0e63UZdhi0UfsV
UUkL7ZYEQGTbPZMo2aQpCv+LXDPVBdmQ4zI9YreEUfFNsyHwokuJvdYLW8FBV9/Rd5qugRwdjuvk
4JeZ3mn45UVBdsEEkvHf4hPeuFoeExquF+U7NCPja7ndvz4zZo7triEkFpYY5Kp4YNGg9Pm0oL0A
ET+TXKrEMCR8s9eCIpVuZaZvLq5r1xgsubaQ0iOt8Oz0CVsCuIsUwlQKR2O9C5nvsQ+j14JqoxGz
zsHNpENHbBZr6SLNfOKkn6lN3EXzJ0eEahc94oGVI0eWY7O+GjmiT9ago5XaMGZw2ocwEHh3m+RW
+bPAY3k4HzRQWaShGaovzh8sAuEajTfjShPuyFnMkfyZmSb+xstn18e9+aQJfczzRhIR1gJyQRJp
2XuN4tS/PLaoSP3pyUHvSVigqPC+up0FAHnxoOSvWNJ/eyw/FozBYaoM92NO+D+ZHKOklJtBgUBz
VE5gYXqdyuzcumBcLFU3xVyNhOHgTNlt3l4PFP/i4JEjErnivHkwoILFGdVx1rAzsLGADIi71Ctm
OU8tYiDvQxLIkdjJCUj9LfJeAgfNF9DiMtXjCJjjDuQj1eMHTA3478mCvnF9Mw0XDJFwUN1L6mlv
BQjaay+2cxcjFjyt+2SY05noENrhwitnvTTm51HRUQ3sbej5aAfYyl4FOpJstPqtgHDCK2Dq+5QG
XiqQPJPdfeqOojWtu1hCCaCxUHPwgFDeTViIjlYPphe9K8wS4Zt1SkNq6LGSGsYyHhN0VOLzpt+U
2I7fbzVDsGFBUSeEYZxVzLvid5A247jxr/M/WaVx+TPYOQZP5e7PAywUUoqbiXfYnXl+kcqRMQMb
Fr4Up6LtUSGQd+Tx7jYujbCiXdMxElFE2f1kgj6PJV94p7IAvp4r94oi/bu71oM5J16b4PpHQaev
8o7v/VEaJD3WbDsfy3KtMkN4FQwEFKmSF3e7qo7EbI1y3RXpucBRgY4hXoFW1NWZuviWnUal1IXL
5z3pOYq9Fdqye9ceW+NmBq7FhN67s2xaWiYD1tyF3wRBJRxdyzhS/bHLDvChD6kxIm0SKg1Dy8kU
OvD55WRcir0FoslMYyKsSYdFOO78+rCyNsFCTQHdDR+2l9TfJ3pyzG/auvZWYmbm57kZ2uKvu4uM
xWxt5bfWyeWpOv0TpT3hBTMbH7tC6adJKa2VH/u8Lrv6cImCRjn1Zk+Kors0xMFOZFwBXYbnd/eE
1Q2lUl7CminNqp7sseItSlKx6EdOAZSOG7WqQpLStW4WsqpnbeVjGsgeSPJZTRqlv59jQW78V8YM
niERkK33vddwU/3m/UYZmE2Gg9kqL3va37JpRcaEmEYYLYGz4XfLdByIfGBqkbZyi5Fw8Wpq8sTG
JOCQRyaTrJueOaIlU9UM3xpnCtW6GJWVWXDmjlNPcqMOSB+8CYl0zlwEzNji+OqfMySR+vziSu4m
BqETAZU6+lvH3gLWXb1OZWAWlenS+3ezfrIyefN2eqaWRQ0A0ChnapNoNPvBcKHMAb+fKoC4Ljmb
K0fLNNi9/7T7W2jtdo/2wrh66wuXF1pan1eJFMi+Iwxib2VdbrU7K3V+7h69zGlzmYUpHr6EZZ3K
CGmsU7h2fUbJS/1bol/ifz6/B13Fc8JB/4z3BPfwACqF4q7FSvhmtqMHpDyd2EIFZsJqbdBoj2wt
VAeKh+RAHFnLwiUEmn5JB0tKNilkzNPvg9VTu98lfl9GSyFMzv7Oj6beISGyyw2PdByR5WKB8yeW
0NhbjpPexeP7oEEkLAxFtZejF/GPqkDSzp7o8p1opZmnuQD5qjOgc7Lg2eZOtxCE+eVHu1lS0lMw
f/bhoLp0PZErGWOafaDc0I3NzFImOEFDEBrmj3M3fv9q8SQqZn2I6sRxDfRh+QLwZTYrTTcR7od8
j0Hml2rXXRIrCSEP7ZKacx5bqnYu1/6Y9erRJ2TGye7b+yFCLEzeurF3sT+9cahlgLziHdJ1dKqZ
8GroguAvPD8tXANLJIIFlxifaVe0QxzZNjgcxPibyNLs9VkSHx/Ucsc4oa1JnQDT7gjia6Z5Gy9P
Ks8j5YfYCKCs8grm8i73LKBi5rE2cuZIwQPGGQiZfXTy/VtTpZvTye2nVXQRQ8AXlsCToF1Pbqjd
wn7gZuRutNkyFSVxT3xsG19L4muDvqJbtn41Yb87UPs5YMVUHgCBRq4ODu65/kzacomE5Y9Q5Qh6
PprJjFucmLGfDfllo3mXASTMVloe8okeLKAMAUrKItKGB44SuDcjBI1v7i0gN/j443WfCHffLVjp
4RsMvbBeG9h4NTfG7PINoVWIFuIgCpnrHfZem+cxkXQK4wxp4nRrXBkiHrHAeSh0zDEN9pQ5rk5D
WolOezsuhCOGROgm+JFMq8D6gFIXniKbQpRrq4IIBP/hIRNQuTbLn0ymH7WHKODrxGpzacebBQ0e
BzWxpQDhBghGI93IG12AGkXdwBrKJufp8Z+osL49AkguYA2lWuwNxbOyzifA8k36Hs+05WQ52Dn1
MYMcYCj/xDurJc+2Y6QowBAC4VWzZTkFlEt9+ye9m2+jNu8nB8CEac6kOVyLRMXDRsXnird9MPTG
qGNOMjWgjVsMRsMTpYbK3+k/FGdeGCVVsUQsFhUV6gBRObKriXaabuHrIx0tRvMwTiR2vCi9j49f
AaxDf45jGNaG4PGGY3kEIqbQOwQwUswuuJ/tAFGouUjwXJLZIUtLxm3byAQCJnkpNwjVjM8l+lpq
uv+uWRb5mFo/zv4oWoLwgcBqNsfiZqqqO5ewGh6zCV8uiAafN302WJsXPAXMBEmixu2B86o/AX06
0OjN0xHwNaIk6VjH0j8sd55mHOztxY6QWENye/S1WHrVG2aj2EkSNd69ScTRMEoyRKOad9Ep097D
qmzhUJo/vUF7mUbrqYYmMF4S6Oqun/nxTENsQVEKa6JfIgOiA5HthAhYvKGNgTnIF/7TDI3HxOoM
lMdczyQX5PGop1WLpwzZr/VTBMwQ3FnWqKTByF04KYBbCzCBtRCzraf9P/ULYm0lAXLXpBV2rlZy
7Y5+HHLq3u48FqBgEfVjHfuMNBNwtFHRGj7f4FLIeJT/+VHBRhM9fcSyCkaC2JOs8bRQZxxV5o68
Ygfgi+jd7ZXgVmCfpcZDovghpGmTTBo87rUIaG72rAuGlNzvJSNhTzCcq0w1BpROjAM+QRSCBgQG
7e9RQS8CujyH6oigi1YpBnXOBfGmAQ5+ae1qUG7Q5WO+Nrg8uLVjqVqiDZWemjfna5L2i7iOLXLw
OmPVESL79i6Mwqk7tl9yxnRbQZ6m8fylx8dIMmWyC64W2emGuS1++S7HPnupwCxaOnpNLMz2NGhm
NJnvAprtz5sxQuZMmEMm8Z8XXHOXmYM5wGHjdeq9nNLGPDc1vu76u8bOwVG0iKu6g17Bn6dSUACn
b1UhUzJi7cN48jqY38AbMPxxKxX83YAgBq10C4cDTKZJZ9SWbtRZRui2usDr5qVXU4C+ZxcOUDAp
v4T/vkMH+oytONZi6hUjZhpHu2kKMS5kw5FOCmecr+Rxbtt7DdBwPpsJHOyV83dxpfl6qxV6U0Uc
l8ToX/mynAqmJMdeiGn4TCIOZhp1lMlQTpFLx8MfEFdZdLvCU62uFhN5ppfmLAW7LE93M5dQcrO1
e38kOnfiKbXafJuz4xJ9K1Zo9mr3k6MAMx0Yqn9gyuGLEUrdrLydcqPUfUIY2X1bLsLULYQvAzSS
g4Ri/9900qce7VTl8ekvz7NQHn8HPVnUB3ihQlFv6equ/65Ipk1P1OsbTtV7AFSnJlqRSaRS+Rd+
+52a5gqW2XugEjIIp8yXTIkLEf/oMMz8E2nQr3DfkJD8e1pO6NCG5mE3xRTmlPHj8JtE6lejcU9T
fJDX1wR9PFjdPjcrg7P5xcRPBowpYSm16BYJNrynXHV/BdhPCkWxEo74zRWLvA67Uab3B1EigGk5
SU7mfZ6P7ZpFvIsWrAQ78zYP+0aLdNPQzCN7+g9wi8v75lfcVtu5EBAmkMdjCZQATA+WTh19sUKG
j/bFt1IPxJfcRUdtmxw8Mk+QX0P7Yz/L1Cs/eEaUXoqp+lZWMrjUOUpbh5BPDqpLlDbaPIorsCOm
R1mXDSLGyqmDBSlKBbX/JJS/3oRhkUPUcptT3rBTN4rwwoyMClCyLkm1nvYrzdBJaCZnJR7tPQnO
oosQqwvoMrAbeSueVyC928qOcjT6fm18AH/MUwxuGv5dO3sn6XcNBu7+RRFsrply2DdgQq5aQr4X
h7mhjr6Fk5L9DM+hToL+R/nPX634c8ZDlUZeYSOrqZaLq/9zkKynD4mriOCNu2QIiC9+yyPFb/Dz
H+bNd6k2td4GamZuuQufzJ2Sqz02j0bX97YwatL3x/YqRWREhGj/3IFb4HbdkdYqbJ7XgqirxoN9
qCZh8dS1klxvrsxwW9jOZ5DyjvmlPzmosetG6mLNW2t9hgzrQzFThfHfu0eY9GqdOq280HkfGw1j
XL09ynTQHnZ6z28jhr6+pyMGnIalI5K+fCrbXCsuzo2BqfT4P+Vlmo9Blp4kvCBTBn9rlbr0Wsy6
WP91loRs9JSx6geiLcnTZg8Is11AfTUEG0+sNG4snX0d8hjcB5Q3bqs7ni18KIrjMe2bK9S43WEE
JCsfE0HRk/ozBDnekajSeOD8mxu5U+gN2OvTcMs2yW7YAxMOosuOwRXBftHq+AS26VwLzkIgF21i
n1LhI1gTEMJG27g+sdKE3cJgO6Uprlstdb8P7+OeDUiRE7xsG5fUvLIxt6evE56292LtaXZ80qOk
4E0QBZSizc6arw3Sj/cjs5L3XYdCbS0eK6cOcVLZ/+/aCYwt4LTtTyMT1gR0Etn2IZBvIyElsuqZ
tvHO8FGRCF4CzQyTaw47un9VL2OeQtZWFKfwdiOurnvAoN35SA4ASbWT5Qbh+ZMvGk84k+pG5lfo
kJOIFTKB7p2hI+35b5YOiTNaMsIAUvaeNv1RaBFUiup2QuZEi9wtTuf1Vun0Sgpm3J1KpaiFXlHW
FC0M51qpnmbkBR6dC2YzmDO5TnndPIHOxXBR+wCuRiGCGubprIbEDCCl3BJcHb4HysqICh28f7ay
rwhmCVyZ3WWRDq5+0P3dQfBIM7yYjeWh49OCVuH+eICv65i5okVVcLdwg+mbDEdpBTr1IcD8gqp7
hknMFR0PqQMcXmY9RvnjVXYMxm/b6GGFlOUwajWrbnC70RBn4xY262ZWlu97FNOrnMr+u2pzkuR8
EcBYxnQDV42/J36FKrLIRjTMWXiptvaDozHctwAVjRkjYWkNi9fNS3m7VYvliBfU0jIyemW3SnZE
OPDte75eyjeDadm45ANNw4Ro6439bG3T+mEF5YnaKxMQOtpEV3iHqSgqb9NsgMB+65cMlnSr5bxK
+h5m8NG0P7PQ87Fh6mI2F19H5N7LPv6nr7wOsfqtn17VIhbPkL5uNw96JKu+dQo31prpUN4UycEC
/6WwhStUAEuZ/0WeFhNlKBkFQfKV7gfYCdepfC7acq4FEoH9bSpngIQgsNrSsm4+w7gnCJLZM263
7snZIce8KcUIdefGrY4/fns4zJTunMjlFbQkwARHFUNRcoC/+6iIXtMUIrPN0y55hUU7NrHl/czv
mhpXXQlL+rxrj0WrnLEId3/YQVpZc+bsfJs7Kz2eZUV6kVF+H0xO+6dKv5kl1RsrBakryOgqmqPC
lmTsMMGzYNsKd+5LoRCFYYiSe8tyeGjbwfV5fKvvNVCzIGb2c3hl5N4OoTxKnIukwOyYFJELqh7v
pl5if0ICI1Gn6h3d9DpDwISb7RZE35qzzPu2RC1DlkfDRhlFtaPbuA6j0Eht1g+doY+uuVsYrybi
dzFmthM5NrKr9McSR378WjcecY9qVzf2V4E0N/xxHQ6oNJdsGM6QnT3iu+UGGvLtf8Xo9Oy/A4sB
Ct/vvMGFKdwlxq+qYO/F/XOiYF8hlYqpeBHmhvVGOZ595QFxmt3LvqzCdCrfnEmWk6umkTGeZVhN
yOZpkHz5I8nRzldwc1Gsryk0XjuKnN/kGZWcgSYP7A9smteRyQwL/BtbkYPa/sMZrTDY4o1vkQGA
7WcztNiSyXOPnGzrAlp/yYdvCS7+JmySJCyPz2le1yKVslOpxyeVQZuVoQB55yedWUKBdIZQXbxJ
+uA2fgku35GQ4QHvpzslWAJaTSqY0QDCxuMt2ZeOeDMsgUEFlfWXoSClK/a+ByMCgix0fFgiAg0N
HSUOi5BK3HVTiVxkhiiYIBOjfyfRkmga5J6e0kTrYNacDUagkZUGkUL5mRhAbM+Gth8Wg6sqwLxZ
OFWJFwfMwuQqLcFMyWhuUzCgKAufqt3EfK1rF4+E185Ys5AEiqhLVrxNNZIIlL05J1KBFD6FmRhX
l5aokA5J9xmkJmhzDwR/BWhL6V/o1bMIuyoy0eW9YhuOwTyL553Rs4DmZjMDlzici8HMWBvccxEy
gw28aKgt/dkovUrD46sGX/oGKxJ+Zqk+NNrzyClFdJ3vTHbAwxScyhH035VdJE4HAuMA+QIIl4cK
gluw89mHtfX0u27i1Zwn4tuSGkd7XOdze19W+nuwjYdbSPO1j0mSUh22IcYoDPmXSOdMHnlseGXi
tAnIoAmvSaO7ERgCUb7hrVQmj/1959uZwStcBps7ACJn5H7ce1thS00Ku526sY0tSUw25vd2FEJQ
bAGY08HgLwC3yx6a8t+t7FcUg9laoUzfyEBMm6VMqXvrXTnKg/ohVojrNsJhKPpdlp+q1jTXtY0M
Rgw5t6i83UkgSx5/5GAgemb048fHrfW7gD9El/QqiYXuL/wcOGwGYNS5ByFVnAuUg2owzb0rpPBz
PTX5BOUVp6/hf8aYHX3aWM4jPj1SxM1sg6V3g/H8114F8PQJXKN7Hczh6GY+5Z2xSjJj6VkKm92i
105HKx0yOwXzXOYidgrpGEW1Wq6gE3y174vTKBkS38n3YLD0yuzgVmgH/VhPZ9pAsJgoqcSBQMBn
mvan93F5q2SqIFOIXIAiWI9iZYeNkPKUk5N8hj5JuWbVvKJf+nF1m9Fj3yZuBp+kDVIh0kA1zyuJ
TxUZQKKSfkWHe2a2rE0WKaoACY+1+Y5FxJVIvFlSFwGJq63rAXzbrMZOm4WzmCTLxRilgRklENtT
8B9VdoAehKtO4JQVry5eA8mzKWO+RePPWKMZ+Xv2Ax8Crq2S66gqLlAXqA+T6NtJlXkMHZRLUews
wub+D+itoGPQjup854hGhoEnEmpLVuYMqVLeJKBcnxTRFVqPWvbC2PnLAS8yE2eabuxMDmp+ZLaL
hkr78m5LGi3TXQjvks1/qEasq1F+q8VtXyZuYF3PXFSio6VALagdBZsQe/XPpVgfHw10OEveXG26
8qLiK/BW+0zPrWw2g2Q1hr6+qUonn0fgOz54IgBO6N+x3wSafDK7Azzm0N8xHMr1u4jAwVL4YsX8
8Mw3aRaKFBs06IOZOqlQ8/KtDpdI/3LbD7KI36Oz3r1rwF3V9x6+T66XovMT3v9qC/h3+a7bNrYm
BgMrWmNaov5VFh3KkwCAUnvHAOSNHfQmHx6d3g8wOpfg04rcKpGqeTJwn2chcjl8utikHfqfvtKp
F0+qvRgvQ5/WiaOnNEu4Bj2aiI8EwMQeIt7UB99F4X/E6ItlXE9LPc73533hZcHOtmHz8ApdyAyE
nAbDfOcfhwBxRTbnXzEQrC0ias2v1EPv8uoh2/6jlLoshLmSWUpZ60X332W+38BMccmUQYPaHaWk
cFpftIY1h2hXPL8hib220ZCUKto/b/RsHYVK7AcbpfPDlPpPrnpr+tcJ/wSUXT7a5/vbJJhTvSUn
Bi+Db+i8pqif/dOjbZ5mw9vgDMkDSIAA3jSWBLIdLGreAG7MOV+aeTFsoQ7NAIdouFDv3ssQBSG+
T1zQkXExAmKQN2Q+gpDSR0bxhvdIk32iDUhuXSQis5fiH40lKoYxbLY8uTpGg1CGGcpQ0dHyFEV5
utYCXSIKI6LS4Nmb6M//YP7YGlBhAC3w5qGc43xfs6Z5+tbHTv2vJyu6IwZK3ic5q32rTRQnqiAm
ouv9Or5G3sF1Wn6Ed/J5g/KE0Y/oSbFvfyEz9OMVWe333KxJ3pnFLGvVi38CRPbJruhBr5oyhGzK
3F/xyU9HMLFA/qI3FikfkQ6SFjqZ34jsrsF9ML2wdGplpovbV1Qnt2yfdpBtdosoXJeilXb1FV1r
r3+QCsGljjdgE4PGNsG2urtHdlJj0bIqALzbnQJHJaXC2PmTHiVIzzKB6g5DB3a+O+5w/aQZeMew
tyOZ5kb/X3v6itZCP/g9ohP61irevekHhmDc92kQ44YeDRGihp4cg24iZ0PjLmpnavoBP7062ljL
2WTQaF1CTqa1hJmt1kNgnIqujyju4DI7knLs44IudbCfYP9m3KrkaLemS+wIlfvwdVBbo53J03+1
Fbv93ndzaP8VsFtuHKlA+o83lpMF4Hf4l8E5NsuAHlxFDf+DhHOpCCPjnegacIBkjMZvGu8VUIlm
ADugaLRgA98Dmd7ARkKFuFwttVsrLi+VmmkjWK0zBzk52bDX+cwba5vxqAWVys+0kbghywiZmNhO
0DAxapkzLkWLhzsw8eE0hxQizunu1AinlHBpn1z5LWWK9MobX+Hj7K6VYRVWutb9YsPwIxaSfV8I
l+hNHgdacluq6T8jRI+3hDqsGbTwZ0sxfJJa9RBtTneq+dZ/ouICeVRqzd/3eOSdt50n6FLgtx1Z
QdBNgeK8beWJKXgs4OYc/4wJOGZsZQjNUPRucs/Mc0sBZLZtHPEg/pDPmFK7VYkRJaMkGG3fknfO
RMxQFIAoqirTRzyFyyQPtLBw/JYCSnIyj/t/CjYjEExgi1mwsh+isB+BKuElk7A00ON/MuEa5pmH
y6Qeuzq546UPT77J6vwEFdbDnqeZfVkTFfeCLIEqRDCRMg7Q+hm2HHYsdbDj/LtH29Tv3suNUyYP
EOMMz/F3E+ON1+TA6tofmlRLpZRH69UTo7shbPWvD8AdlI4PVgWtw/bjW4YNM1SuHj8yThmfMY+I
PscXMtA5B98O6n563aYKfogjsTmSVNLxvOyOpXxU42TAX67sSnAoPbBCoY4e2BOgtZVxc1pAKcNu
IU9oprkXOianjTCc9ZBMloEdJxPHyWX3+kE11y4zI8nt7iRLuIshlSJbjXBqitJ43H8CW1OXEs1O
L/XVrwIDfx9FG04m8OvMOg2jlTURK607J87FzwjWYtG6+uSHBl97j821KcyndJknQgfadjWd9DrZ
u77zpOwnRQoLm5PjgKtWLvqPAAuIT7UdR6SLS2lrgUPk35cq7KCpNBStnjVU4jyrVnDFbH/5UGNu
2z4lL6WxBUQ9o0pglmcXR/eFdshbBoGGjEl1Jtsg/D2TqCsD6jBjoKhbz0iI8M6xnYlrUMk1q3pj
zJ3E8FQRr6/g46KGNsl7qdXZRJlu7cYAGdlsoubZhZ2Oa5aQ0WQzHtJTW7kM5nnTmvMXOHZ6yt9P
Hh7EhIADRAbZNFsAevXzYa1RkQ/lMF2tfQZn85wQUljBVOu8cCp4c8aTNuJrxv6AJJ+Cob/+10Y8
dLAJH/7G7O8FDqpod2chgBTfg22K4DZorBFyEjiJie+QnZKBI+uYgS6qg//HCd4YyoycLv19j1RC
vwntImfbrLHP0SY2wnfsp3hyyJhLGze+dFE3KLDTo+D4PAEe3kKnhxQTAxtgUz4dVGVI3YOTqthh
JRbwlJgO/jxu00/nbr8pxrXxmqQ1lpenW3Ahy1sshps/Hpt6qgExPvW75qP8GM/Pv5GLxmb6g/n5
oIvGL5GeIW3Z/cksISb+zxXyWO8sPDC2UUN/z+5khB8w5UPFZAijn7iOA7Jv0IXdsh/ZH4fXCOK0
5KabrpK1X4Am9CW440Wq/HrEzG3UUgW33dDl4xelj/NXz3Q1nxjzr+b4BpRIfvOnDLO1p4z6zAlv
/GEM7V3cCNhAcnC9iKgwNRZ+WG6ve4EN19UT7QsvSg6wZyQfFrXBBFrYnEVyuNOuAR5BsNfGKheA
uMFWiIgNYtTZUtbD68/Mr61fLO6r3pe9j/StY9t/WqiEVhnvVdpvPgyBEDPVhq+dVuUqGCK3Uqx+
98ODOXL0/dXu5FvWWElghAUkefC1Cjw8+O2hQtWvvFb5u4wv/1mafS73tOm6h5nxPKJTB26KM3mN
MWTBenYCqzRiUN7d2o8GLkmcpQVDBCdK7j/TGlQu6+ufPCpLbH+wEvEGDzbtTroBy3/kG6qoUUwg
j/x+BcrdcqBXUC5FY+2fHWiC744owBYpWRD6jwXKas6qn6rV8M+0DmueIisFOjv78wWikSZpQi2f
0WrSP1xwJFpZkYnYi81QDzCA5tt3LC8hzz1b+FIpMZFTCJRPkYlR9Zx+OE+5RypIYtyB02VvcuyU
dAd1GkHi72g6gwvTntnvcTLGwegiqkDlGtxCXKPr455W9k9s6Cgyo3olo/mHKU/1KYBpjg4eCZ6f
kgyGEAzMLZez33RpFvhwFnnvCC0ZsIE9x2YZSrH2/QeO/8WsQ23/qWhAo2gfZy/kAwhDwg3FCkqS
c64PARMPjwJWQ7znoPUJJukY8JmRMkV5C4foY0IBRL4bJBOwyF+CZvvtPG+KRvYnHxXA6m8TfAKS
DZPsMNpak7QERjbD+kxUSLq71HXgftBvxJQH3UXMV3aDNt9aDLzFah2Go54UVE5YndHM1h8q0GmO
eK2/DRhOeSuiJKg227HUIdLDctA2eu7dzNoVbeQw1bw9TOVoqZFv4MB/enWqDNzIovga8txQK9eV
aI8GCzRSbdQzsqST0leOA5S8pk3eMrK80YbMG+JxOjH2KUzQt65fNyoht+X06fiU5PsfWEhY9/nG
abGmM7yUg31PuOSJH91TQkygI9tJk6GMEFPur/u5nKtnW/QgaIy/I4FvDWWh+hjY0Cki7GA4dOd7
uH1NkH/WZVh6OMnYVf6SLszaJbWpln98DkrgzI1wjd2RSh44UxDYRbxL9Rj1IjnJtXzbu41iXyPK
ptcmRmGcbkttLxCvrs2ABAOBOGrnOdEM7KgdzLrrD9V3k0HiKsAqaondnUygV3f6cM4/KemgoMuW
mhqBEUIsNvo5/bqCxZQVoAwRo3w/kr9BUZXdiJnjVes4qpCx9nl8Mp+6b4VSb8JAZt5zjDQtSaj9
Sl6aQSkOwmswl2VKI3Yv8bsGGHvhJnzmhpM9ErDanS9ZZc4zjPo2Kcl8Z3UtPOtmNyBxoN2VWsNP
E7pndH+nHwvdQkmndYAjgvoJkcP52sFS158xdVyUefdACpI74QtUhHkcjuvzQFEala5lU0jwLwOD
1UywoYsrdVeIeu9tEvlgyU13lxnQukTQoaRuljd2IQjAG8o0R6AOhwFc8SnADrnQ+oTd3/Isk6TA
hOeiDU1xhmhSlv1p/S87T47sX5rOweiAw134KjxBUOF+7vyz7w82H9JbxXxcNX0LtVndeLCMuWkR
fpXYwt6O8E1VxTuDuIAca10a/KjYizhcMFHsg0vRcwAm2BPJP2jGb92E4WeKvH5Bdh7dpcDPZdKo
+bnftBLQco68PJCdjGxz4gakr+vms8J+Q6P/zDoyEX09ZK4ejIvMrxmenzJfbpafcRc7HEs7loxq
w5TD8bSJ7TCyziBkjv5wFZCZbGNDd7eJ2BYU08fdfdoG7kwOHy6T+ck75qbBz6DSowa15NH0EldN
XkIcv4Kl7dx4LTbgut61eFDQEWitqpgXAMQKTXBXds4K3wXGltQDROYaFXjtSM0fNWDBhfRXA4b0
hgA0Dh785kzIzHGn3QKcaAX2dRoSyZel3T1LzgkXESCRwbIAWjDONWoMvsI1HF5IGe6E4owFkdPa
qjsi2Mo0Op5qRl1++UkgT3pO4TULKztpmP9zzdjebwfZJPYXlvWLgRPbp+Hiv3L880TccOda1C4H
VN2GdHKNRPUIb9eX9epZ/Wb82Mv8XObS2VN7AmARDLb0sr9yCMO/abM1Sk+vRdMimaZeJUMita9A
avvrhNCi36CBzO+JoICQgQK9JAOj7TdOOtAYNx7NLFuV6IQgn01J2pnT5CgZKuNpnQ6xxZ5p9m/g
He2xMWla9Jq2405i5azUIEQUp7Ck7VBIRzZY9gO2loTX+8gvGxp36y7ZSbkOxdeuOMPJSBUPMBy8
k+U4yfOr6ajXLLGuOiVhlYSCs5mjtiSyXNfWIL1WOQ7BdAeqv5rgUuViLQKxPiQXhXSCSUPqmvwM
HMF8j3G7RkQSYvdDGRA5M06QlGpeT10prQgpVFzg2KKqpK9gCHWGAcJLGs4NPjFBac599DuaL6Sx
TKtRw1x1OQgnmGBQ8AwdfNYK+Em2QojsUevHkPERfS/TvkLIZ8utxwNb2GVTYmmSqDpGazLDxjKk
J7VngeNsDrrRJPkraCMe6bnFjfto47/WfwK+ThvGLb2in7/K1pBd1tCbcAYQxA13ze2eExyQesyH
TVZFb2er1p3oM9H/lSCILupuwboR04T32ZgwcVZSJ7m3S040mCSp3mpHWXDNXmtlIEAWnnyk468c
omcUWqSQ6ssWZ/WL7ghELnZ3YRnuJXDBoU2iK2ppvLYen+aFaO13tQJ4vjAIBW4TfprU7pJU4xst
wj5ZaIDemI9V8n2iYSdnRnfiO0BEqibL1LAVi2qUmOvkU4eDCap2CZOFtQ6DCMexOh2Sonx1FOjn
c6NIJKzYMCmYt4P8DNbQXpzGxI2+H2YWDpRxdJ0n693Ztpr9AINJ2ua72ZT8GhjzulLP0IXNiw0t
KWfJLWW2pPWjDrdGAVYfqoyrb8NI58RpQGBjFu2V0tzponDJ8qtQqSQ2g1INtINgYKsauHCYbo/j
tTaj0cn0h9yHOFlHUDdWktsnZ8fkOzuO7wi+XJvSkIB1ellIvtEpX+8jThJGzEO6rhcxW9L4xTgy
t0k2ul34kS9ZO6GRp6VDQE8v5HeuUlvJmsFoKhnBEIcP+SXAQBcjSUC0OtvGaRijcgmlzFshPnVV
0haJn5SWh7Q9KQgb/WTKmSdr1SRCoZzE541h07M0joL8cRoyAff2QYJC4yR0yak71vRytrGE7G1K
HXjvGLReB1b7Sd5iWm8Z8I3dHjUa47tLk0McSzBWZLsw4xvHNOWL0UHz8DpK/FOyNwuX3juNJ8e4
OqkMRh1AFxntrKpPecXmGFIdUzH45eOfZYLzzUYY5iMEeQctM/4/Il1wMeQtaSYx/vtQea855p7Y
BtfaqVTn9twD+Is/pHuPXcd8sT/D7Z7x2G+9fEpwVhL75otdtRwMeyZUQE2s/85kV0x+UnBZ7M1f
KzG599lCo9n4FNQESzSeLPWOt/NvcmUDPcdvkvnbMqSOJhDpioABA4ad5iCVABAJ2GodsA4u08p9
Plz7wsF8h/70Klg+hCZHSXUTzbBEAQtDdfsLypPcrQ3IbGEQPRjxNLrCnXDvYVIHPnimuAVOLx56
e4/AxP/yUxC10SAdr66L8mprSroUwpHzyXFNOC8vpke5uLsSyZSTkq3g5vs5t/MRPrGqNhJm9eLv
jliivrU9Nx+9bYOh6e7YzO6H4Q66VXvtekkH6RkAajWXz5R3X1G8SjuZ0zDtvOLjkpoj61CEPEt0
MYBFzLenvWVvLUh5AUHn55lXlh/TrLG3nJDnSiISCVDr00xCfg8b6GIXg0Q7nU1InFvIOwLk0VKg
t+AN7GEWYDw27SeSFfb9wFrFCdMtWdWmrwtC8Hnw6/sPvC7r+hqi3QNl1A2F1vcgLBhj1bj23lxs
WBsezANPue+oEu7yrQGuH1YK6SPGoZw7GD++4/+nPAZYKr5STrQYmosJgOtd32RYtHyopmvdG7/x
1l+j8ezoeBnXkIp615JlUPX1qUuDEYgtITUbgH9LElfAQIoIBctgiskSv+mkBwMAPZxzxh82Ci7X
90VoMzwSdKB/fr9CcKmdkZF/cLmNDSe+KQshlTAtu/iGLgb+BUYDZSWE7aj0cDsLQyIivQdHx6c5
GeFN7w9saJJZkNPZW/fA8qUQeBml1Te7HuNtjRt49aoR0HnazZHW4fWRzEa+PFeMHGnOcYXMmB5w
huGsAY+0eqzubwPGDltCt3bP9DaO4cI/BFyrRmvojsaTKNtTA2O0YQDGQ0YWwiIB7zimE8c0+VAn
ChTU7ChiNuidogiuopcKch1NCf2o7PVsp1sp4rNiLtm1dKnPLrxqD3iZ+aEXC1GRsp02JtG3S3a6
TkfDSowao2BR2m3dYtkDbJa6IwcsAHa+WTOpEkO28UNvcHgl8yY2lFIiosSctLunYRP5na9XAQHb
tLn3TUspt7T3uyHNsShMMjoj3aM+FKCvjl8Ts6JGWhpEf+e5Eu7KSVNogSZxJvKCuUb8lU+KrP1r
FloENVoyRzhMCNxC23mG4qOGY/id4nGs36nDTuZK7lGSTtzSQLpnxIGzj0ISRppSkYHJoxtZsfGS
Y7GQTKI/QVX8dOaPuGCDpjb1Mpba9cU0ZJUHHCxMRL0b8w47zcFXbu6aqw7Ckrg5uA+4pyIy9uXj
Q2stcdbAfx8OvvAEYmOD+LVCtkurMXTMXhgLtwBzmh3vBShkEw8qxTYM9mp6hN+O14VVa9a5i1eE
o/aPf0q1l/zTFJp9LC25pQ5oKaH8LA+G/XeO6kkTJzlNwKaPCkWQgqs31iGQeISW8adgD4P4oxFU
Uzp2S5oysSypjUxtRkw7qk7KbpztbhYg+tCJ8Eu2LWWmkPFJxEL4WrR70nPjIzTEcfZiteUh3ncs
Vmu2jkdhW1DYDKyhY+k41jPU3gtvm9qOeB7nXgGY+kmC1JqLgbol45P4NK9e7Eqz2DPduzYRi24g
7vrff4vuv+fGHn/oWYityFK1/P/twMRgPz4bP1sZdS9N6Oke9Hc4Z+Oy/JYpQtQapHb8EClTIR8v
TdV+kQNQWXi6VdpWOXYhSMZrCDkUlhl1el8UCuJBFKEP7Aqy177jJddUOPnLnS+5HiOkGm6Px1eE
PW+1NRuHe6LrOQwJNU0yWyjUJSSXs6zaHPzXUJ9eCLkYsK5XIQlj4sBccsGJgmWLKyYnGzqpfbqr
EpRlFeY3TYNNb3iWHpAnmKotdOoLZGSiBJNvwLv5QeEdpSwFUDOV1UYyvloiOGHR+h4SD/PmhVkv
KDDT+6LGrsvbwKISGi6utjfEQZKICNuDcjdvtlLNn/2jAtGbjZcWqOI/qwTN5p4TtQY+lWKVjhlP
MBIoNB0NXfhQGWaVeAo/J55qRB1AT7DNkzRWbCc8QF7SiA29ctpSG14SJnIPxJPsFy1pilVYoXJ9
79jiRQCtrKfo7s/6OUE5NH2cmUvZLqNW5vQs3HzDS2dH+rTAuiUSc48mw16Eeax8OETQA9UwQhfn
KemhOMMQmFUt5WBGkuDGZYn5UVgOL5R2inqcejUjQOpdiOhH3eNJ8uoWEctlRg2aS88hTnVoUYyH
Vojf4PhoXJ2zxnNPN855UgndY7OPoUKZtUGBbLYBjP9EWhIyZ057K7p0wEu04tMCwsxJgAkqlPWL
3t5eRw3fiRdvudF425+9IA4ij0jI3SOTLVqY9BmiTSZ15HGUgefaB7W3ojhmr9n2m+8M3bglG3rb
tMxqXwbAAxVJblrCcRYXcZDZcuuJtxeDyEQEMrb7phtEVaEk5DTzo2m2lvwgXIi7pZiWiiH7Flw7
qdJ3fJs822RVVflpDPSX+BAzKexy4ZOQ9MmU8Gex+Qle4E25EYWFH/N9yB7AzjCKkU99rJtCQVrl
UVZ9U+/ZVcV6snOCuBuCQv1s0u3Jywie1YyMki43QVEP+KSbCGJk8sLjZZiQh6hfq7e4KWiZ36pB
ZxUIq9bVdTQL+Zt1bRGJwIi9NZpHZZGLj2Ik5/l2shU6G7i3Tlmqk+BZW6a2zZt3aQUmyKVU1heS
hWHZFN5anfUH3ZbVAUkOdlUM3z2eVPazdIBz6yR1XsE1+VDQ+MJfeKdenHbngq56mHrWx/84qg6v
DxatGhy1GmhvBgs1p6K0/Bxu6AoI25GAgDYzC7zqnGaiX1tYidDqIdzCfd4zytjhqdc9bF1w0flA
qerTIvGELdmAV23Tp0Djwa9XZ/70353Gj7zBljLLvyTOswu5Et547b+zUr2OrmeuPMgcvNuj2CMD
ig+ML0wPk9fMelvdWbw4TpHR8472g2MybNloGdbTz8qPL7T7uFMcETzCGb6owfWyUjkggi+GHZ0F
QrxKurmlcZCgqhZF+5egG4JbTHj8ISBm7P6fBu51OsS2l/bpMLmIUfiWffmNnGVAIkT/aZW4YNBG
hVuUjzuwMLOkYTV0Rhy4B9z6e0YZrl9bwHodTZFkXiMVvgSMI1MZYRMdimfExie7oHU5IyTZwlkd
RHK4xFOsYM9oEBv7D3enY/HPk7rQyTl+PQyUDjf0pms0JUyeJONdjo2D3v8vlAwlj7IVZj29X4M7
QN3pHHzzC1UeWQY21oJA13gMG9mlm5t2RNaJBXoJhIinD/ebeuR3X+UkIpi4Kng3QY6ajoJ0lYKJ
vKv02sFd2yCSyFcIZv1goRtpJoWZEaRi2gIa5IRROJGPWoaTPXN+2jiV7ipOC3syORmnXuI2xsp+
rInKGZ3VfxXXomgu8WfqEwP8eGx6yGzM6iwJDKMK//L7rewK6cQBJxN/Wj06konHCCP7dWQjD2nA
P8JoQPnkoJQbTyqbYT7IWExkkoS0WlWiRV5uCQY2rqdp6eY/y4Ue3q3byrKXZvQ9QO4PFkChmple
RyQBO0geo99FAIKoIzaskEfqY6NTvS30AuEmNwDwplbXeqvANj2KaZGGclKFDhQw6H/+AYaGVYjm
tFC0dZBoEKoq6D1F4E+/Zz9fwHgMAmfWhtHgzwl8L50PDKACOqJEogOyzB9bsrL4bYxwRHY+Z5NF
XSpHCz8wdOwraWjfv6Cow0x4BcZpdWXnPVtBveLgaNvCu4mEB7hSD3+jYKsNgj9CMklynTTuEo4J
vWi9geLDwPdMiUIHXL3OXVRB4grlXcfKjgSJsu0t1c0fbAm0SWLCeI5S+jVOWvCqx08LWNbZHqiS
fPe3XHUg2bIG/x72Xu/4kl9gZqW+XmuPhWL2vESZkWh9q2SBeiRlIJ0IPyJ7U7vec8WjjkBGh2Sk
9kPW5UVn40X5g9ec7dusKmEUCaTNBGf4/keyOSasAcIbmWnTWv9+NKDN1x0BdyTNJFf6ym1ZmM1I
OsSgKWpaGOMPEd/rmWq0dxeYXV0qgpx9QNrR/Q+XdFPh3E0f7p/MeiqRbaHy4whYPmR0OzblgxQa
9XU2WZvGGwh1NQZyimUnr5bv4aIT9OtDFt1bjvUOCItyDvx+YT4nawFSgMYzwi5hpWhav2DoFTnk
kiaXA1CW0PnwTOkWuUJQXznXgm9giZW885vq/efKsDd6ZU5a2UN4RP+mc6H39MRoLZ4zQRLhbXrO
TC5Dh+aXjlJwkb3jqCjQ1gmpLo8y+PmU1A2qrx3b6Zusgwxya8NlsZfVObhFzlOo/gZg2D0ZI5hG
CwOAfwcXc7mdfZG4osT3OhJla2ENlilr2IGIu2nZV5huoTfxxjv7+9c+n2/xg7L4kUU6M5awVqIX
SUlHGInnoJa1tFINRlHpJoktcmpF0AKmq70XYSpE0h3RaIiuAmhyUwAujsvLuIrzZuPLCZu8lVSh
bBT/HSUC8fs24HictaYMlcVa0xjHYAESyLaa8p4NNGp39CHhp1oP42pH9M/z5JTelvPIEeu9S816
dKJRT/3qPlumTSmftOni8VaUZleXC7NJByVMvi4zDJpDCbQOCodGPuOqAEcYS57Z1BhHz90PT2co
8nAomF0eEOK7gGfmn6wt65a5AdZMosZ2bF0uClgx9Q8DhCHqmz63iM47SQowbDJ4dhTB8JWYbOFo
5l2Lsp3YwiFKp9TAViijTW7FQhaeHQGohS4TtagBhLIQXcy06YIfd+dtb3e8rhEihKh1ww+WSC9p
Q57BpMMjYRSOKQAOLNj1szmd6YMSSF1oYP8FmK9IP0ro6/QnHhWdkBjhIMklf9GogcdHNg514XvM
XuBaNfTOGy82mu0jZxY8YVEMwmYvAzdjPpqz4neccwtlyIuZALS9vj0bwYNDk5wsqgMZpl5Dg6JO
vFVCBGJ1xyz0/N0BGyUA+etpqzINbgxkHg7MhKmjn/XPEFquYzcIzfHkc8/viYxNKEXjLL0P7Mlr
4/J5EIKu3XRTQyZ43qiVSKFwOONSWTcQyg2Nagk5/tNZEn02wpr71KDjpLrcfDGvRgniyGMW1Abc
7Ci2PAnPqjyRrHsWP0q5m4ljslgjdR8e9vOzs2CjJ0ZaQIRbDqoQo/iEOrU8Ab5/0lhgmTLJ84Og
nmmqy3KFHtkgc2EASaRoZzDg8SRtPFC5d8bhvPMYkBCn/R5zlhr4M2bnwcrswVUTKB1rCbkz7NTp
7gNL/KDDUuSt9KRtOX++Umzeg1OS42/ynu/mblxpsNp+eEAVeWfOllg+MgGclUHJi3MVqTv5Cnel
Uy8eb9UIG/cdQ91h6FcnueCO/XZ0md8y/dTrCCb1aKQx3OUIp2r2a0GCc4QjxY06ZuyTnFHj65x2
H9UIG0Zq6PGyV7RZu6Bbkj6zM1BNoaX8RZ5ZkcWA4sWV/Ov8xNmxIwR04BE5t7loB971nrpqVuoA
DELvOiU6x3Cxm1Waptea6+KBj01+7lXaRKf5di1aqPINCu4gV9Kbw3CA1XCln93yBSM9xbYKrZ5Y
tKbFMEvHUlLqS4jq8MC/vHcrsJ87dhcwtVwrDmBiFe2XCLyzxEstNO1dyb+shHuy4XZM8gtVxlUz
ckVY7FY38PaND2AocyIsBX5ryhVrUlg2/zdsDSuXWQX/q6GdJvYnVPMRNJ1Z52wFGbZruzf6Nqdq
R/fWHmgi4HKgmQuVqyWCF3MbauFB9Y6jV/KxD4aww4/oC5Lc/fVRPmpgcz/yGvPXW51W90QiP8dU
D6UUBOyXlp1oVgC2SH53MKdVHWmR8/Uut77duxVm8tMElN5FMnE3qhmafwKRWxaG8YO42UKPFec5
K6eAyNChL2qkQsT1+XrS0846JA2BN4mjSIUKj8UwV2E68tqiueJItYmHnmTkfBwXa2BAMrLpkCDm
gHd7DSOs1hNgFjQqLicYWR5nHShp1xj+4rdg6LqPyf4mqTdm4IoGoTwU/+DySvAUEHfghdmmFeCz
/IThW8Tfdao51hPwHRwGJesN4Lb2BhigmBdzsEVzrGh/l58Iu37yD3hSgeWKElYqlfIZ9FbpSpuG
PZbx3BVrGFUfZvsS8CIzMJhuQjEt9Wxr90tzYy3KixBHCW3jMpbk9ROxBxz8hwI5OO7dq3Eebmil
FiusB5SCxlYBV49khyUwKZM7NpJLXcCra0+FpYlILsNxdYJcOgGTp6scvl8/FS8JDZ5qNIwx6Uvh
bjg9FDFPjnYURBtRTQH5CIg1JIZHV+eo8B0cTa8KKJKP+v/lTT6EdqCfw6Vo2v8vDyfDJsz0oYN/
/B5E8RoexfScCl/GEUVmaeh216UWUh3ryn8GdVQBjnVdfbBA6G7yM2VO5wh5Zt08BtdHlJuf/lNv
8IQsXHZDA70vSnJ8cm6zUvqLGSEDJJp+/rIpz2oIVBntXpbXBmaPvfVSZ2jmVQm9DkCHA+3WI4da
b23rpG2lmomla9JPsVIMS9PXddznjXXAlZh1dqOgIg2iqU8M7AIPxJpx13Tlsb/cCIcZP5vyLODk
w+WN0tVyge+pQ3HXVpE8EsMdzusPp47tfciroofB+WM/j/cyBVkYU/0jbfYBounEohYk+Yus1pfB
okURk9BWyXCtqbfEsudtdKpsUKDGLeI6Y2zALS8oRFpfk3pql8IcNmUucjtaaPA7OGVDVaWLtZG7
V2Bw4A086zPpgAa0US2zR+/C+wJvDTd3PJzUEF/suxmpiZcMrcOPQIhpQH1h631uMoHyClR5JyqJ
7JXT3QwYzurYhaIwbDqrFcDzOG1gC5NzkHOixepyHEc4l3SthIwE7uC4jjy2dtSoOSTqefW3ljCF
r7YllKjNsVLmSVEF+jJqWFkiLlD0L34i0Nx6Zv17l8NpE5UYCIsvf0Gdu2SaQS+JX+UhuFfT7XA1
/WpZVbV+I0l4IrATT+kd/QHSH3QM1J5DJlw5OyVzLf7OcqZBv8ZfeJjox/JPm+xa00eXjhoBF7yu
re8O+2OnT+8LRXlh+qDU4uGCedhO3mZ8Onm7bWtIrEBZBocoi+wSIOGmXkPoBIU66uo94hj+2vk1
jhNXWNWjqskYMw7npr+iwbB7Di1o0FOm9FZTnmd1SFOvPyJD0QeRbJaA/+N+awvvamhYldYZ4oST
NBdvT/SKfNHUeghenABLYYrr+0wooWW1qT2M5y8i/6QfGA26t+X19tmVl7ig/2fzpNRHbYIMsLH5
/Cm2xWBvZqWS8OxKFwaNdWTYxCnSrgKkifU06HV7TgsASNWepinnw4faRIOfrkYQiSns8gD74sUo
J35A8Us+VJkSxtHVEKxM/81rKay40f3A+MCCYKYph/r8oDxwjBUxcDPBTbsHYP3LmU6ASOhSp9aB
XFGRAUhQS68P5vP5ih1z6GIPjpxUso4aey4vW7kz7z9+G2E3Id2bD/1K+s9TM7VKgpb0FY7hIPf1
ELiUXiJfyGA0Mu1y+qioy9NAEOpQDAW1J1gtYPnlPaBF5yjQRK7Yz76bNHhKDVhcGdAVfJ3Fe2ej
0Jx9QdQgEhdcFdxL/F1t/ntznhyGqLhdCblo7a1xlC4V0yC5b8uWO0JN9KczPPyir/sK8GhzTxsq
T4UcvQLAgiZFVig+FiMfrcDAuSUsObNiFZjuyvpqN+dErm5yZ9Xpn93P4+46zMvV6blH8SMCoQWG
TmtiIgaIspZz7KoB5JlQe4ir0m0UVJESDb8NJgyICgc1hUhBOcsVRhjLZOtTePFyhtKrexExfZHD
5/hwI+KhhIILZaDJPIZKfRLUjlkq75WaR3YkClNTaD6XKij3WmI4SY5oiWX/pMsJXb42rM/SxTMA
kaYS8bLp93P3jLn7xyR2ssFeAvrLzrGJSvw/dBsPQiO7FMqQCURB1zc7V5yeUnpOUyW9pD/m1cqx
J+KksNEb4TPK0ccdtGk1hOy/WhqF1EqkShNYkNMqnOrxp+sei9GuCfu7y1sbviZHgBRZTZl2sHLT
iP6QCjgz+H7torISztr4ZHUshkVLrn4zabVCL1Rz1xu/1uYwhpXTCeRY03sLPd4Rnl4AnLaJlIP9
8caexLForYtWp6S9G03GrcoHm1ha91IPoPeix78DADXihzr75A1d8SPkM+o625X+QkX4BwPcR7z+
X2Ep6aWCK6B/9WdyP9av2QcwR79RjKNIme8YyBKCUkyNzj2T1BaK46iYk4aufKDTKhFwU0wJnhOC
DF6qBgTEa6QWhBTp1XYeyTifDE3Rwu0GherIshdy0DGD1+JWZaR0eXWyukkjr8n5Ruhd7HbrhUGZ
ItL+ZG6KrTIZewNWhsX1Sej5sfTphtJ1a2LnoNDU0C+2wCRnGbkbQbFnNSCSMoimLLNy2z5MMjCL
RPGR4eRILSKd7fzlI9MC6049Yt0PYgayy8axHxQNpOSQET6/hBldloP37T1eJ+jfdZpPmA9cFgAR
MUNR2/AxBA8zdDl+RCb7nSj2L6PnHA2YAHsPMGUl2RpUDu/bGXmDR1D1yVV5hjZ3dd4Iv0pCxU2N
/+1V2i23UOBy0tTTpptWiHuRCimBHoh/mIBV/Gd3jkTStHoY6Bldzaals10U1vN+JlX2coyEP0Rv
3ixczpmia9Rw+pqBkfXgrIOJ4QhQ35VCcnb7FpSSYGh4vbZ+aBcErTKx3DjC1DVnIgswHA7paVgZ
cL1RN5aPyGxZDVywx3rZHT8mEXS4WsyN2sn+/Fuj9NyhKk02riDAcNMT0PQVY+WaOqfrVFELt5gG
YujXW0vAgtOMjTbgJ6Gn7HO2yBRaMrOCNUwM8iLLOAJx1NO1k3RfHjiojNkdxldOe2OO3yDYBwcQ
G8ynihXGcUydDUlSoQCprj3yOk1FuMxXXDQKG+Hi4YceHrJzH7rq1CuwJ00z56go5qE63QftkoRF
P0D0BZe99mmuCph77nATOqEOPpeQkEsdalpAa2WPor3Sw31RjnZfaIpg5FWiDqrmFEDW5FNqzlhz
fPzKBQRVzTm5j8Iozt3lPPg5682CInUpPUsNSHsU4pb3r+G3nuaGCALeSoURwbeUsr8iEkzuDjL/
eqXZ4zG0qPXz0tUKWRkgYcjZwfUSvgZWoUlZHnkQgKi3xoUmvzGe2PjB0cxjBJ6WS0W7TTXU8U/v
i9c+4CeTuCY3OKmZi32WpG49+NFEddFEP0ai98RJeROe7WDuSi5CzQYd71cjytc5ryQ9qFDRSLDS
MGO/EiL4p4it+aP8NJWMYp7qRovOOoL4ytYo6xL6JG8yzwKLVn/W29BXUiVuEJze5wT7/TcjHSpG
VmG7WpA06wRDvRYbjXQYoEXmqBGCzmNDMvOccqoj6SIoCpWwzwNilcf3UhWJKvJr42I8t3gBlH4e
2uOGtiY+cfL6qTuQ/igs3DcS9xVrph2TRHbnoqh01dNkBOPVFk2fiMBGaKN9wSV7SxSIkn5lhqOL
XM3w6TH+lfLkht4+B0bhHxY6tBdQZxdYBXnH2/88OYgKX/XgR/z5M4nczu24IvvvopmHLc+OnEsj
XxywbU/D5eTnePzhfme1I6GgAH9FHkQGrQjQ8a0uV4//Py4JLRg/8Tbnep7q/yslb3B/BNrUdpOC
U0qfyetfxJtr7q6RtI93bK3x0KGQlsC4+pw+YjrTPtWaNyS7VnGTa/dNfWLAIzz89cijvHJA8blI
amrqMc0J0lkL5DO6tEf4ZuRJswiJNkUKL0K7TBfMynrIp8cNFvG0i1Y4Fh81gxzdxYgcNlUxr7zN
wbvLW5s7aTQ/VDhMb7aocbq15sadDG6WDXGCiB2rcX88OneCgf0mRWo6qx/SItFmJDmPfAbgStlh
skzngnO5Xgh0W6/uNTNBnJuxawc7KeElj89VrjanUm6xuQh/xVjUmiOKFBDr7lBu+PKrBxpgUJg5
oo1krSbh5D/z26vBbBB4X420xr+yd5BEynlQBbONsnHe4lVsC158sHlEIVfNvrh0FLtif26j+u5C
csa9kFxF0fjZkzUiOd+VjnOFtYDkyIgfdkUKMUhEQ7+GHBIrH4CF/YRbXXII2Gy4mA0GJzQF7ysi
hMWR5L8eQFWVqum+5PeYnIvXvN/mCpfwUgdVtQoS9PTnQYP6fF+QquCDkVzVHofRoEMQgRoN8PsD
Yn/w3lc/GwCo/cOeQDiEFLHJCYzkPoJbFpeCyPhs02YZNleg+fkVE6mo4Oh1s7fwyahwS2JfUajT
NFOsKRXoH9GdsEiN5+uPbJUWG5GCTpbi8+G2BVYHHxncihFA9BfnD+Kl2lvvFqPtNENiHNk+x/LD
e0hAEcmCOMLZS95LJ7S6aWMmUORGvjq2f8yNW/zK86VULSDz262C0pqJFdndGpXSqtPMcgYeEPx/
nACvaKd+eINWEO1kW60aiGfih59a5CgLw5tmidysc4aNe7a1ghg1aJNwDzCG7f2Wa33QmmTiAUbE
fe3GutwHwDFFtAYc07KvKWQETZa9S4byXybvGNgE7OGSVmIsG6CHDTkoW0Py2KWLHbKnZBaxLaLO
STuzqgUqhtytLZYeW7caoJm9tWaEhtyac3GyPzqhcxuFKY1sLMidqrOIElPoT1kK+4zSDbR/hoYV
u5hSIcNzPaxta8NORAZvvVnl3/bxJY5h/lKxmzSvB+Zq4AOvoouTjAMpZINha7ABlKWbljGFlOOo
HRYYPYdneB2WP6unPm4YPj7FDSLoznU8BxYvn6kKcNmJOK76jKewiv1AMf7pNX44f2dBV38XTsEr
xJTlD9Kjf1uxfvYeRJR5qIkmhPuekMgajg3nwU7I9uEFqpaHri/Em2mOHckrbLoNvtvfhSIfbIEQ
DiK3OgX8FNT8AqSYUXNYpSL8X+cwiv2XPr2NpvlFSvf8KZR/H3uz/3fQP9AClSx8ey4UtfP5gh6E
Iojkvj0hXrsPbRdj/fqhxTmrRj5zE6uPdYLA9UDWVvzcmndvdfyxttP79igTBxYe+MTkMzDIM6P1
SGXgxl8mGi+crljWn8wUC6WeUW6DXaMz0+zFr9X/61WiRAOzuiDgm8kgMsFLuTezpawEb0yTUI42
oWZZPf8ONCmUyhTg0Am8+7XnaLS8QoBdHpbQ2UrAwO3zMCwtkhHRD2HJtoNbvYGvKZeLwXg4y0BC
SVQCsUT+mbtYaLf2xVNHXWEqpucdX6cFV5aUq8KRDXdgn47pnfFRKnU6KxRh2XEVA+oKMxX9z+s9
F15NDpwv4hutw2CnKGZCQyNLWB5+gRTYlOMavhQ+EBWQ96UbGQ/DbBU0udesiMSocu6+y48tqe0E
6RmExrAGStTeWwLxSywyOPf5qVVagZqih6/sy045Du7cyemEkyw8SNYUZlTZ0JrBWYDICTCBNB1O
FQklXpP1BSuOa2FmzkQEDPmHBmeYezu9N9J7yD/Lww0oQqHBF0uaa5Zi0qjILZgOaF5YaVuRboWf
bzgGoxzLvsMc/SAIm9vsuKDKuKbPMVqFDhfzHt6nnnXlAtVDXVAhnSciiV95ZAfeEfLrEMNsYnKj
Q30nx7WIX0b/pPA36J/Z6yowNm9SOMqEfxtrc+1BHjOkDVmwmrd94zQEl2cM74HeFxd1SRHYEgfX
nyf5t6YNcR3oB561I4eOkqek8ciuUxHR0bi01IztiwPoDpgWkEpUqpLDyu4g8k37DQG1oAYajxqA
mTkAPl4ry7kQWUuRxYGUsQt6bzZiDWi3Xddxcbg/ly86itqYkBvtKu9XI4NLYTMJLBQvwmjKAa2C
JxS2hYx9mQubWH6a5hR9vM1qY8CvFHXKI8/B4oyuCVyQ15B2niumnuhqlo3rT2Vq7nbJkOafzF6w
H363bkNekFipAaD82eNy0i96Q014/ABl248ZACVLVhpqx5ETVpMggutbW9GhXys1XMLp5JryqW7B
2t0acrZIeA861bgU6J8HUyA2mPq4PHiWuxg0z5GJCpXQUHhMdw+/G4TSmU989Phhr56uvnfbGuE7
HyDOuBDcSOAABCYTqxJnZApJtepst3b62qjXnRKiyAXB7zKgnB8BYWEL18Kz7siU8i2zv6cKJO8B
zEDA95ruL53nmnPtJTC7hoRnnsFa+gIJ7emmhH++LBQoeFsEkNqeF+6yl1xO75wX8XclZR3xsrwB
aN61TC5tsfdmdMKuaGIK0oSr0SyY1lhC7t89eI0iay/+vnesnMEIhMDImmcDW24zEyfiQYK5Ulh4
s2cWX1rSubf96HUhnpt0D4tAEY3cKHNlHplRKAghUxG5u/MSvXHkzTiRCIQiI7ELnJcfAfjLU8oU
T9/W/yWpLMFwS9f6pv29l0chE+124l3+Xao6JFYjQK+4kJkYfkniPEXM2FnMAlND0h+ckmOZrGnU
y4xTJi9WOTySRL9Q0yz4s9JVPMFpFV2XHaEZT/24geRmd2AHrHWrsZFC+qFimUvK++OmexOlFH5M
J11j7iBDOCf8Cbq5eG7rM/ZZ1CHmj+jOYVlcNdMoKlSQp4pUR74/svpcSbsdxOtojGlnmc4jN3mt
5wULp8YwagnFRQoZwi6CBkvbDj6abSHUgnU2aiM20Yf59RnQPOmGW9+ix0FySkAezEAGSSkryGYL
8Ed6cd28BVRyRm9uVeHTWDyKR0TIcvCpsJu1yvd3aw9AZXHJxSzDG09YykuUnsWCo5hQoyIw+j68
iEf9SxOvZL48l6lCDWXW3TIezi54mAaBC6UXey5qEqrALItfLvlkBgmfSq1dIIoFaRGAC24//04I
2UOTdO4AoctIV2fIe3+jG5S5mJh3EF0zH41c5yrj1i6crN45jbpehJFLejTQqm4tFFtb1Qezs1mL
pUfDs3F89wnxEGDiGETra3ULi+X9IhtkcBPsGmzUtxHLJp5nenSnrJQwuzG8lWyYwsG01VC6GHe5
PkyTWPJ2GVAdBjVY8WpIe0gjLuZRwmoAVQo6gQuG/l8ICQ9jCl9x9eGkBTGl+BukhrCRhOGjOWCz
XrNvFlbOwMLzp9Z0DqPkUMfRPWOsQhxyefDQnkyNbX9Xcbou0URxAW13jWwpidxxgxaUQddy8Nq2
edq8WUYB6WyI4avX2xDlm53CDso+eAIlUrAQo+Q+lMApDLfBl8rt/FN5SwRxC3V1AXpZDO9HvPdC
YIDt+vYjLych1kfj7lzna65VKhjRR9hS85OFnYgxZCW+oM60VVkNDFxFstABzd0wbqGnCI+k3UFf
X6IuzkCPMbZAihDh21EHeidkI1OxX9D7oAw1ZLkbva8Nkmk8FRMy/lwn+Nc4pPhbrREg2S/qharG
btH+7W7aZ6j/cThEO++on7ZWQyY2Y1NDuQjmsdthgN0BT5+QnFZyn6vnxUaBUDm6K98GM0lotumV
3AUgf6QQc3QhdWFaWHDuj0VU+6JSxis8me57X6eXzRZPhTqwhq7g+EStM0yoh165N0wUgBtd6EEh
n4v/k6RKMP7Zbbhy/yAuWRkiREOtnZFuo0BBYVimHrqgETE1yoOAIOxsXW1Vy9tRY5K4e6borEv1
prGUvLw9VQMDARgyoZhW0JBnNcFCp5YENB/jRqvAOhpv2gwYaPjpWmXHSA9HNBj9z4MiF0fbTviz
/HIPH7VXvSwL/Tb385ZVMLLLZPDC/mOb3j3RNDluYcehaVh04bx8PkC+ahqsPcSK46DaXFVhUQ7D
ZwLk3jWMIbRes1toC96ZN9Xe80xLTkswpsa+coLS2+OPGRyXCgCmXM2YgrrWDzo7Ek4u/fR5Tz1z
WHXzI8x2RwLoo+kAFrRB4Ey8/VDfpwgQpFZgBdk8OfLSit4Q24Y1BpTDziJAxmR315zO8CHEeZP0
3BXSiX6IDmGynOOyDrWRaAuF3Xhat7pId6i0UGrc63IuI7uGdyhI3BB7C6Qa4QcamiqH3G7WHXG2
jCWlnnubdBmJXXxeF9/lAR8//qPfmO6vgZZ6tZCMDEfUf7OpRoxHi1UV7q/qSAUJK9PCQzl5r2qf
O5tMMzBnzVeTme6WSozqshkHbHNjxL6u7YL5EclwXxuVe/3bFTGWlZm6G48p27qXghaFEhyEzSwt
ulyyJEXE5RJ/LFCjo/9eH6zFW/u3LlVNmVtoK1nSZ728S3xGtsA2wFODiIdZKDGMWYPEEZgI99uc
EUVU+BpOZvM9PLb0LL3nmE+t5H2imAtYK2UKIbuTqQuMHfuvRLDhNr8C4+UFPhtzC/uX+fiUcR8J
hT7x2Y7L40QP/BcDH81vxpuN2AAPaGqfwTTsDCiJebN+6NbUMSbVfz4ytNpHEmxUFwAfJsfvucs7
WgS+AxVOOdWoAkjsk4hkUvD1UUNJn9Ewqyi47yZDXo83pci0rs/t/ohyfyEFTUqki+qdjbdWBxFW
LFB84EEisL+/CJBUdoPg704TXhQbgoWFauF4PNibXsWeKpWaPX4+3WgBcxilMXPjYPa1UcsTVMcx
KBqiBgKtX2tB7Zvhzg4bNAdDzxTGd5sKedCeDEYvL+AQZr2DlbKOEs6cDVD6/gGcRszSwovf0h1c
vGckisJ8LZUEQ6uHvmxticdNr4/qX+5EKZdMYERKWnV/HVG3JPHUij0bNtLNVpyMqey0Slpo53wr
zY19iQz7FdggrIC+jDDl3maF16xmf+AB9xWbt7LZWTsKOjQ8FDpjcwuGQ8GImdYhRgLUy4kwmTC4
rJQ6tAH+uRQK9UfA3vBUGG4gkZ1DRNa/rNf3ZUoM6Hed8zrNep07LvUjW7hgmiSkThe7hXHbdgrk
oZ4FIrNmGCb2wK0dmNNF3DYg7F0z4odjdFDsHMHkcRDo/hMlUHi54qbciBsH0ZUQdLEKtLtNJXio
0s2MGGR70BlWMiujQZ5JXvWtXenhAJmd/CBBTyKf6JV6ALUwfPQqtPgCAZyjnmSt4m2+g6e+WHEf
LiHLBwKP3wm5GGUQxJF5s0gba4jEfo3yO5DYo6uu5F+Lp4oHltTazWd1pKlAg0joGUfHJgrfdOg9
7Jd6CynpYqI5XLxZgFT1FkSWt7OFKpqHhf5alPX2V3qCspmYA6coxpQgeAV9+4MFZgqcP4EUzN3N
0F3E8ITtROxu0nVqNpp4O5KO+8p8gAsVbCMpTjflpZhj6+Oh+Sr/ym4HemoVDWE1EHY75GzCVNG5
smG7YvwlCdDe5Bw0QntHc38R4GrZ4wMuH30OM+9I0Pfuucj95okUFLi0SDz+bvS98X94GLT3CiKW
JBxJp+SUFyN1f85/RtJIoFNKF60jWRBsm6ki5nDvZE/LF0hIQWluktmfJdQxhK2iU3o25FA/NRxO
8gxY1S7fJzURyiWGSSPY/iQXLFiX3P/i7gnZ4P7uPL68dQRvIPUAhyUTnPG38oR0uUPaFOmJzTvN
Cbqhk4xCvAnbGX/5SkKu+5S6IvypCOahz/h70jcmlto9fS3rV6Hosecnc+f5jxKXxXGMrhZ7UwAX
Q+hU0n3HkPV54U7wf/xNe290DLDhcZcsm4kES0NBG87gDgI5gnUvL+pmdSalCkerTshbsNa4LDb1
3YKsCYm9xqJDUSSq9qzww6bw3u/smkq9T8vqgxo54SrzDaPDkinXrYnQKWXmpZAqlrhj+M9YFYBZ
1QchrIlQDTHkUYvBE0iEKzEVxQ3HrxoC8t3TzzRJ4nMS2BJFOwd0RUCr7F/o7q3W08FQZXNfnWUn
SnxyUkPos2okJnskftpP1nNz4M379APaEROfJDPVHd8j83vWJ+Mzdhih0fPAxLVTOXnbIFHvNz+5
xL0++1IWZKGeXBY3uwxJ9pFS1giUxLuxEY1JB5b6qFl34zK58w8hDGrjQoGmZyjl8Kv2Ym9HPTSR
SxNstqO8+caxZCRjUBqpZadJ2/Qqz0a+xf4da2V+P8OqxjBOh/fKGWVfdIIxQqj3wV7Yx5i2utw9
bQP8OAdw272ecGkd4NebI8F9fNnNVr8NAjNWsn95HYa8J97saZy/aWl6MD3xH/nuq1iT/ZcQnQg7
zXuvJdubK+1uW1Qy5FwEdE5/IdPU3+nGiNpFNEzDQJjGnJz9iEN0M56WiKQoYP3LKqTm+xsT/tXS
EuJDBf0X9NmnYuu3K5xLrLw8wUsHiKCk3jNF1A7tAHaLHcjuZaV7Tcqsr6HvmAf87S3cJTQeYTtI
51nSqowJaSLGDRXcVpm86RYC2+Q0mw5ECMx+6oZWiS99jmR/sHpDvYw6a/8yDPhIC9vmwL6dItg1
OxSi0M58c8qTG6b0UM8J5PfhspKGqxcGaiOzPtMkBix/qJyEAWf0s8UmXfzUmds0jN+hTKOx+svA
GjQW3bea1IY/+fduwSzkgyNsM+dq91nfO8tmnWaocWjxlthGCsFo80K2suzlv6egBY/O8icechCT
LeQbPP4QJzTvkfzb3aBpzphX3hmbhrPe59HA5LG395uXpzU4WCwC5fG6X3nJ1vSi+D+MpCxuM2N5
fkZVnQhhZYDoGpQVm9hyEExMSZGEkWNPvNif5ytIcO22X7kMcRZawc+COlh8GJ2xH5V71G7Fw8pY
vdF18jRl0lD8iiVYYPXokzNLN/pOo2IUgRQa/LvUmrWtezY3VcJYLuGYDfPgEDxDT1B9l5cNqA/j
1jZhp9A/mWloGE6Veg03wxyfmVTcH43n3uudSWEhXrmnkIOgfhIbP7ATIfBOLLaJLc8TtGamrrnH
mHvFtAOJPNtRdwg3OisP3lkKBRcMkqAUyDuAJoRt66vWb43cafNr8JXyyAuZiqWeL4K1zrtwfgae
/j12VybFGPyGOBxntmPzcumxqsgIMXNvpcEP9EbzvTbQuK1EdFz4yK7v9UrPKDbcV5S1PRL6GfBB
nwetm4Q9UCanmrBNyWJRnxX03sVAEDXE81oHR80jB9qvqFPUeziGYuBXxJx3GgP2A01i+pEzkiny
9xDWsxZwlcookTrp1Puv+Ajm/EME5Hat9JRagJKGyroJKFBT454cbaj8avCCyovi/ubn0k9RJI6Y
LJOUg9YZN02F6ot6HUezGDC9DwXA2G1eWkiQEP0fr34sKzVayvE71uA4LOksXIJ44ZzELB2+goRg
FTx0K4gWVHJPXvNV6BVE9ND0XlbfyK60OTFfVf0OrifxVUBYsJJa5/psHVh20vMgK85WP7MoQ6km
YflTOZzZlcSzorSxQqDLhp5gpeqBsMPPOR4bnZpQdT5GznARJbwrzSgyU2uVzPS0IsvqWW76x1cT
0dPInT1lNZzoBtMxhLnr9dznaVXmLR/dDhfK+BQP924r1ldBv2qULv7uh29AG7+STashsvFFrDf0
8yxqovYBosG532/olar1cj358Vie0/phhrpdV0Kq6wl4Io8nkZ4Q/0SzoXAyde7z9MDzE8UB5fna
HBPNGWWKxfa5NAD2iR/8mA1+MYrweXASS9DcIW4K7LTk/8j5DAX5h0kPWefhUOqJcj8lYbNh8TjB
ZWZbkKpvan3aFMoB0QUG4TnBi2IkRbi004FpjXDBpHRJq+0FLems9XgVLivpkIgvhvVx1FGvGl3m
YWxf+MahJ4q5QEq3b1snZmNh/UxP82XCZy14T/ZbUmSHqK5L2eApgu/d1TMVdLAo17GQo6GctlMp
D0OOzk0bAQ3RcE+2lAkqq/d53klsm7cccUqq8SlHL2TDJFfT5O79NPnTL22qx9AJ1vyu0CAMIKFI
YmUDWLQvdERoyRfCxG2vBdIq9RwFsr3mSsX091mA3Sz+yNXjPSjupc0TFAsHFyHeezhkH5dSGx/S
wTIgZR7gQOE+3Y6GHOnAO9N0IuZ42M7/X9CddOrAWNdhkthlL+dFGaxO6AzOr4Zs7ozbqFXjNpz+
5WgFlbKypB5YYnEo1s3IKDBB9asK9i74Wj/1EIZ9gZC5s7pwgmDDnpnyh3UhxqOrt+XTd9vT0qI1
1GTV8LjdcedagZH2gPLseJwzmPLYZE5CTbg/R+gUShyAn1SQRemlMEKQVtsLO37g67BT7QZpNgIB
A94+8b6dqWCJi0d4PVlcpgHtdPQcxVM2kmC3UObA4s1r5Ljg4nOvd+6inO8yulWk3wtPlyXo3G45
SUVVC5DiCZSQIL0p1cSBlczoEl+fmDiu6yO/Q6Qlmhah5PRUTTPLj69IkLIQItHwbduO+TmF7ZqI
CkHDwiPomfkAmEi4SShvL1Y1X45Z/o5+GCKcB0z1aQA8rdqRI5DoObHnNGbT+z/bsG440zZFIeiV
h2I/e9nXet6uFYrp8ILPhNUslmpGl+jK8gcpdHzkZItbbPLeQrHdwsgSpxAUj9Sv9O1LPJ8hsi57
GSuRvqHdqSQXqZlizQFV64k/zViVjBgflSdecb13swBuZ9X5ZLWD03m06OW9ZOqwb6VwvoC3OsHX
3l7a0SvlvF0rApJyXzaNqUUzoRLiiU5PQUaBHgRx0SDCA4IBiAykHRPx4sR5PI80u2j4vUSYG5tr
ae5NpWEulu9kl4l6PdjBs9TIF6dOHiHlcG1ibNA1FWbwkPPHXLxn68fXzL+HYGHDA/Rt/BjMvBj2
/lCqrRBmqyemnldPQuVQkBht0wPuROVpti3ZuCIeYVqyJMGVEBOVO20AIVal6HW8o48w3jF0m5jF
+YJG4I5+CA8ckYhzhnJFLUcmEZE8Q0jpGMv8fcHn1A+dbkMCrN0OXLii1EDEPtjVIiXoMToHcv4E
gvGauuPwgh9Sm14X0AM8yrq/mYfLxapsLc29d1mIvxlJW9Yi6NDP+kFuDGJKtZmbcc0FhWol8oIc
GCvJxsgEcoK7p3KyWRM/joKEMY0CJdMuZm2m9FbUvUa74cEO1BxLEwa1hEcmqTyUM1cRO3R4KcVa
V3uI//btcHGlq3KOmdOyn2d1ApaxHKMTYK1gePP071B0A42iR0ka9bemSgVnMtcW1E5n3fzvkAzt
U5nAJovdPN1FHdJ5EkeHoiVzSGe3gkBcznHiHykTNuscBt4+wPLLMk1z56kf4kEIrynYuho+ZlXG
bimxIHnaolSlIjem5KLKVCXUqc1rLIJAaN8JTfwpZXecICLSjOMm0q0/8uRiajn6i7qkBsYgn7yV
d6X6hyvOnkj+ItvEADPKCrOI56u3QUy73t3pugt0EylZ6jtY9gebTmqham9li9uu81X5GOKZH2qi
KCVdl5brlcvOHJ7X4+oT8QFAsc0vTLwjBVrR8yAF5n7FWCQSDDDv+FSDWiUpnyWMD9J8eC8UdtEN
VElGqgTnyoLHRVbTwMGZOgUjRZ0EsH775weBtCaqt7++Vjsyo5DR39obgNdu+r+f9Z7I21KfpSFb
bXwWpwUoRaxgdxQpTLWo5rSiP6qj2DLVAVyZzS+dvhKlW40nC2MI49qbTNr1QQpOhV+uR0r8Xdd2
bxBMWj+9lTIvKMbEpUf81REqTyGpu4nrtWyv/1Y2IMoWcNOFOSYw9CWM71mTxjUcwyExX1rrvMPN
pfJWv7i609fCt+/s8zKY1379V+v67jlN8XCmj+RNHtuQPt3t6nhJPID8xH3iiwWpB6oNIFvQ6ILz
oA3YD/V3OER8xoIGc1LscVhqB78Sh3PpoY1GGKSypMpes5EHTh19ZYQ6hJSTDZvp7CKUaPD2Kl1H
8bcEdoAX2rQQ9Qa410C4DEFTcQY/XplpqjA0vL5n78kZyA+2equhOb/bPannwVxO9hXSZLZK8cB0
vEcyg36FrBDTfa9+XxzL1GOMA3V6kLCMtRNVtlM7yZNZyOwMYPh2ep1+Ss6aOyiqVyKt+w8Gk+/j
MZYxZq7xUNififLf3xLMa3wDrShpYyNCJlC3ypF+A6WMV6YnoSoe8/BOrxyjh15Kd43c/HJjL2vm
yKU2Fwp6x5Dieu0ZQvwuS1BtBmn3K928McokzM0pG2LvQRCpcU3XgEA11X3tgEspzVI5mBKd5dxh
x2/EKTpJppEKXenG4+9TUZoSOpr66HD1btHnipQyxxxpXo/L30ICgZ9xg8B9kz6BzfLofB5G1lnu
L/gfNY4TZUHAYzcg82QIwdFGVRwLrPp+Wvrc4zCXkhdSlK1JYIy+cxqbSVbyS1hcrnq7hEkxPtcl
woGmGkJOxZE1FgQOvbSA+nx+AwiHK+QU+aFA7MYWFeGh15M5wIvjKQ3gSVIm6udaaV6n+MHIJcLT
uEiPkEJAM/fJ7IiXdKL0HgEPlZ0HBLz/rw3+AuV5fohOqUbzNmvMay+dX8NvhipTJY03A+oBUIx1
640HULcDme+NV6n7mubbnKLZdt/COGESU+MgkKJ+aFBOXX14pPzk5griRQnDWiKvUF/SUgDPEu9x
iDcJuAb7b35KX45NcbbOJ32mAIM9lqQh5ovtuOyf5A3OT3vvxS4/n8o2i7X5jWD+gEmWLtCX/EDL
SL4FuWc4T2CaNBZqTEvFZecxAXIWG/ZAJgGelDggYDE8c0EbBQU9QA20vzjNkzpH+lG1Ztvj69c6
8O9jEbL+E5RQ/YanyNGcFfRAH+FO4UCgAqvPlArl1WS8VE5O9VGtN4kQQCvzHXaV2lj/SoTSnQcd
w+pAo4ns8yh9yllMT4xswhiBFv2kNAsN4yfIS4tvr54sP6VQsJ0LU1NaQtz+Onzhrea4p9I4hdg2
bPEemUEHmSI805+srbRe+hhav9A89B5sOEE/BgciO2eqlPVhhSDUxkuA8ZfnW5cR+xH1OlgH11/9
znjTffWrudNIbv37ZC9w0/0VEt2yAXipw+If66LND3GvL3EyPWlesCCP29p5R66iFRDrKPTgqYC6
t2Rb/r4nORwd+SfmR/iNJeOFewjiN9AfjO4n2Ue1ffyCjrIAV9Cg+t6Xeh285MZaBsqNN4fK62uY
wL9ujmjelssLfCdx0DjloMTswADgwP0tPVQC++3ZNyTbVMXhjYN4Kubp7PVjePl+eMtxLUxqND6e
yOw1I/PEH/yGlmD+vggkjwTDFhR4CkF/hmBZUn2DrnCa2pJrJCBogSKC8B9xzAU46lex4tgohBYQ
vDNcxlgCr4hCrKyKFkFr9zY0DvCcvFHHCOjVsA+2UCkRCj5HYrABDcrBaSXyYaWYP9/Ztgw78ETs
IGLX2DFwJym1yET1yPZVwU16qP9dHThcHJsLxeTsLuC55CNMluKRpbmFAwYIPYBJU2hs13VThmL+
5hNjUXBznQsHfbrdcfTzBVOj2oAX/RibfYjKjmBumFHYVYHUyZyryhY/0BVkPL6UTHaQhYZMHz8R
YJxHOgsplcb1I/w9ifCR6muV106LWgZfm9fpVFpzKPnsPaP51srAB8pY6VOOJ3FyZ3OMOinJ7bM/
1rOR5DxaWgtvs6hSc4oa0lOL4/rNOOa1xLHwBZKzpGzscSBxedeRMHgBhAgnllTmDenLK9FGpZyr
Lb4J671jxuoFZ36niaxFvnvQuI/55gy4LlrYY/rcotpfbPEP3PQ0uKQU6daS1jgly/1+FiF9Kiia
mTvdveqyeR/lUpC0ypyb/NkGxpFYOzY1C75Cd5b0ALpjH+WRjbny4Go0HoLOswSmCnPB9HJwzkZG
104WtFo9R8FpgzA89GLhSFgsa6xN7hZxtW2+xjCUny7YxbhbwT/A//IzF3wXo52XF7iUEU9j5nZv
drRBK7zr9HsaMBIt+3rCkU3axsEQGtTF2EvdrDKKOjndr7guxWTaGtoppiO6oNUE/FLxnWuzcVy3
PQZTZ1HCNBccbCTa+Yuc1bf8huIJ9Bw+j2CkJ9ibARH5DMq407hJtwxpteMD2IEAitufk7RcyYk1
2O8fOdbpHIXGl0/cfnDyC2MpAo08vWMjmSsL6mnni+XSEme/UV1D3FsiR+fRlSLczKO1yTPH8HXz
omzH9CHtx4vhS4gwajnIqiSBrG7g+m/SgXzmyd77zEfGuA7w1y0vmNca0L7b6lDrg7l6cMEs+pbc
TkG4//1MAFoSYdww4Yr2i9DYrt1gtffINKodTwDFV/Stxr3BcFy5wiR65vwFcIb3TdKUTGCL6IXM
5di5R4Dys+uV1l9B3YQMcA0caG4kZjWB9u6pC51AisR+MmQ7ZivV72Ur5gxLAjEmbt4MIvEBoYgu
N6Fj4Afs2oOgUeaS5Trspt+7dIB7gXYaBosl/1HTCRd0zJT3tdwmSRq7hX5IJAfvBdiYyIYTBUG/
6JMFWU2EMkFNr2oF10TEHBDg4aJp+uPXM2ZettVVallbWOZKW5v0DthQChO990FQ7Y1dPTtjUumf
PnpC9JMLtTmFYz2hHrHxS5MUyiBNphFlJ0yfzelPk4K0HBZmkpG1+Ch9sRkVe8ICrqVrj5VMCaKN
uY58nVL7Qpb3ELPTqYHt5FUL9ULjeWjXaO8C2kBNebBJP0LC5FcsjzY/k1pZ7AYoC9KwkBB14ETF
o1AmMwdkI9Flj4me3rZ9YdJfE68KXZxapbh/Pg09q8BN5ozl0yq/TyIm04IoRetOIhN/9kiNjObb
vVFIB0Yi3VqZzmrJV9h12JTp0zuQES0SDgTH6+Bqh76ksYKFKLneUaadYq0SLeJCxiJJXs/e79Fm
i48QBp5ubAosdG81zzCNY9FOT6UBJosjJ1qXwdYOzMvrFzYiwPePXXstkydIre1PgbgVtE+ST3BH
y0OeE0eZYLoIf+v8qrHvMFkkwpoTxC7qL81Axhb9yLoqd59FzdEyyotTBvV+4184mR5axJ2wKZ5n
Z51SB5Ggt6uECUEnzaFGiyvqku19zMxlQhLNwu/EvbQmukXigRkz2Le5dhF5FdYARnS2E8T0XNzF
n8nEUi+2ngdzuxOCxHkOULqEhclho7zHUg5W66w+t3P5BlyjB0XEYptgbTz8EZGPECQTGce2T40n
U0r9OWwhel7ehP7Nk9Epzl5hCFqv+y+y2C+xgfX+wdOMWHPtOtjq0ro1VlOPKKgeRGdhCAK7ZL2Z
qp4N1LGhwc81kTdSsq/G3t4jlstsfEETFuaflQ9dDGF10zvv3tOKivhl71H1DPaDl0ASaph9kPtD
4sE/7JfGxVlzw2Cr34HyAePcAZ/OWbKBBYgnJni6E+Xh+Hj2HFhFfrsLowsEvLxLi+BQObsibw6A
16kroH7zN4xR3Caw4iCt/Vq5q3n9wYWpVf0D7aXivoAB6FIIUnfo11CiB5lFrOdUTZ9O9G81kBQG
J+hVyPjOwQnR+uMGgk469v3LiiuA+vOH1G/USvJyM27oiZJNqyOQWm1PwmhEgFk4iH1dlQ6evaID
kFhqr3W9k9kjBQHmP4N5us1sBYwPyBxT25GfCnjkvLrY8ugg/4ktgZeER0lw0CBXkcKwiA02EyW0
PLzkR36dazRTZ9Rvz5mbcmSMgv6I747rrDoadrRwrnaooayM5anyzjSM2HKqhfCuYhcjlz7bRxOB
/7R5StWAR5pMYJ2xrSOH6+kypTbSgdXKVnTvP4bQUZ9HwwJNCM9xhvVdd1w8YJtUCxojNT6rudMQ
tyaua5edQ5y2mq+hYyel8veJVprh4fYrHXMH/+LjaxEFPRpqr6YMFB/arAPFUIhgt46vyyPt5GG/
3Ifqbl69/zxvebAsBVE7DjL1naMPht1WPTcznHKRgLnJi6X8NVz/zP3YinmVMvd9DKJEIO6OY2gM
GHRVH7KTIr0o6HeZs05zkgZ2W2SuoS9Dwg3qf3alZQg2ZV1uLcsvu7LAAIU1cKAMctbZPCDWshKs
wjVVSNafx96eO0t61mhjTyx8HNYQerca2LxUrdhRJE7t794CE6WDbf9r7Q9lsB4yMrAfZh1jo0+w
3eQa+WU/fj/Y9K1k/qATamGpgXAVhbmhNPJNDkwDOBn3joCDcZ8f6U3YrdmGtmO7GxH+qJEszsH+
00mONYNjef0xnUtEe6WfsQwDcP4LCAx7//nGeByEpmVeSRyej7P95/fD/S9CeAZ+cVN1/x+yR4NH
2i4fbceJN59pdiBCezG8NsomoO2CrD9R9z0/AKWanRqghG4CkxmmgV9vbUybsXh4e9ftLMA8lK76
TyePhINLAVW5c4WlABi49mLdQ5dU8m5oVE6p+bi4eCKN85r/oHcjnjX+Z/elklOFi0XBOKvLFMNl
L1qkNFB9wnYFL3gXcg88V+YUzcDwhwDqJc80DAbpw4UyKKEJDnQtuhJr3mytSTpR6QXdjRxNlEd+
4EeRKYJg6lTWFC63JIKJayi00LJQhprOqQbynnmREvurK0eOfTNozcUr8qAeZ6vWIqXFTFRkNGIU
YmDjX1CFD8aHXz08pZsP3qI/SIYopKo9xBo3bPNwpGFSAE+aGmjwduSEVh4FK++6cNAvt71ibTyp
Ei8QPFCEhgqaKBO5OwofcIXoHglb4zXXePh/nhAErggYag1SCNgVXpf7y1kpB24FSA6v4PsDCaUU
iZvpIaTakNzrCQJqLzzD2CN0t3jE6HBWEvzKIfKphzbi10r8VM6L77d4LAPb0vxIPlrL1iMTtZeU
kN5UdNzRthyeBvYNpqAhqxc6p4z+JNbTtJZiWqBlJlGZTjxk+9zxZADShe6xU2T7YAH/+MU7BUWH
9e4VDmAZYyFdZy4Bx6rDbH0WHCxsSS0Sdgc7N4GUxx9hHGikd95dRHQ2dqioVnaVRcsxHexip6IN
/0/21de+K9wLA38k7WBwcMen1uXZvsSA3Cd2vXLyp/a3cvWIpGQZAuY4CKyraRJMsiDRDL/3EMiI
dv4AsAdP80FZSXKQOd3DMEnMXNtxejoPRtVOKUE6G2fpWU9LLLRABR7tLgsiGBAvtahJUsU7ttCy
E296ijyYRQmXBXfvZCZiTQdpgVpH1272FwsmYTw2Y1C/1eZLtFH6n4XmU8UsIYK6iQj0ojpNXpNe
JDiE477cAqgZOozW/6n61iIrPE06t0V+tdHTdkTwiyF6JhScP5/QpLaAY63YZ/I2z7F1it1lNIxm
yGNSGCxHgG2hY6K1sj4bVlppKT6D2LLpF6vEvy0NeNWn0tzDw772J3cEWk6Qfvl8EB3gtQDWwyDh
1TXdkNPO9OwOYdFUOgYHBRzc3aiqghhR7+NtJv78j/foYLHEAVHuDxJ0CdOt/LPqluWt42U1koEP
uJq8OV4gBej1lu0XAv0tBhHF9Rp8JxxBOguYGcqFVJ9ayRyNUXfBnZSF9mCCy22Y3pDI2QlZVk8N
hguU1D9De6IUrnWUb3oS8tTQIi3o1r+2CZ5uNEp1XPetorW7I29fZNwLQHTEo/lmgpsxH81S1wRw
IhybaTONThVpQOu7M6qVE/HfkYeoOnhQqxozNGZlOZTX9Q5DdtW+e7cxpdcF7Ejh7LWocmGqhUJr
GeqoI/Ye5Wf0Kj8OQjsEi35xVs+SFD3RYEqt/oJk7lxarbFZb5tsoW4jceN12d2wLGIPPNCQo7dQ
PQa+jgY/I3cZZqhK9Sq/7PelG419hBf2woMJVcCtwikAts91uiQNZihQG2KQyyqvTNUZYEs2ALM9
gex6es9YXqi9yJisPbnVsyFoPvtoj9yp5yQbPSZQYhK+Nhah1SoSY74yk2vntyqsEWee5RiKRgAj
x3mm3WAQeOMx5ZOUI6bijay09/ZDth2p7PRPsraD6rZfEX7C0O2MfqAj6pITo1f8ypq2NJYVsa86
XCfcLC+d8gdmTQxovUZ1BSy3dTUf6PrV9IgR1d7PwhQ+NLjHX+HSNJUTgnlwB+FNtQs9urn27CKw
D4qN3tdFoUm6lr1XQYgmXYLuEHBbmBrDT7Hvv9kuiMYguIzUCqMdYML5sNhiy6hzsFmt8PX2JrPl
pu9LiPBtRCCfG3Msgqopxg7+WqW1rI80LqSJzIMMZAxhCwkn82AwIobRFsjE4wgEMX/B1y/TKiCc
VS914oheL+Vg5Md1INxOY6MZwZjixAqJzeCX5PzYE2VdENoLetcTHwcOVUYAI2rIJChCNPFa/ime
RvejUS+GmFQ/3JO1syNXv0ydtR6BzIVX0WUK1AHy1rCKN6CLIc50FYl+1cjzlvR2XLVHRciehwqr
4tP2bkl8I4rsukfBpzoTinzBJ7tIKaT/oMHL0hBb4GbGvR58aW7i7QVTCJs9G6s1OA7SfjRO4OOh
vbkXUE3vjwSr4FTG7MMZAZrtQ2mibeWW+PzFlAV/Ew1r83M96UKOZ/adgGktybWQKE2qiJplJxwx
H+HKrSnPxuVmsq5Zq4h2RwHMz0C5tE5Kfm3pNwo5+lH76Xg0NkrxmKfC6IPs2pDBIiVXeGcvtWDk
ypHAeOaAzoCLS5R2pRkvLNmknvSXGaLlU1rDQR+maIY+m0t8HkxwEK9LA731iEdDdJn6FR60eKgD
uQ+wds3XivWRmu45SWK0Asi62GFWyPSn00PMqO5RMYYalX8kHbRVTRzxQZJUERcVTR9lr3OtEYRA
XZ6N8NBeUzS/baglZGORFDbSfoqrnoWpol++w/9upn7ceTWNl9P3cN1v0xmrFs5B1+3T7w1IRfWN
X4Bz3lWh0ijI7foyPELvK+Fn+6Id3SwL3QzmfZW7gZYtH1yUugqEQ66rFjA2dGSq3Txlx5X1jxBV
fmhL+3Dm2KRfc4lyGjuMP6SlRyPt7Xp9N6oPj0ZYfLgoY4Z0EBWBNv6FVGvwy6TALUr2zgkQ9K+f
/LgGalRFEG2ZKG+QS+MbQpX2Ec6ESpsWqtkeksxpjTngKsWAF3JMfn9ICbZTl/ADQGq42X1+dvLH
CGDZ07K9HdB7tclz9dvc9uVFLPdyzc1ur/V9pyx2y34MLyml6jtyTeJXcSFnWZ4Y82CGJUKfdu5w
t+yUz7gwfSXbBMR2fglOsHKtPDwyeDnN1yjw+WOBYppiPnVzsbveEiD1ohRxjT2zxraoB6qZaaam
ocO9nEKApDeYcgLYHj/fYe2+SHXDq7a4FEOIyc3snKjLg7o0UK0+PYSien06uUIrxMN5pjlmV6eP
q8bbhyfuWeydUv1+28fqKnCZlruBwbDRDCdiGBDKJBfjnPfWhbfH1LbuuJGdBTeuUhJgV9ypn6UE
x/D2O6g+o5gwjjH25tnCJpB4Iz3S0grhTykQchJ0JJPXhExjhbmmCMO3aVrtGP7E5mmw7fnHt+Qr
nyfX8zjrsdJmjbK9sUbCb7aerVxABFxb5wx6PQ/23EJ+DVVLcaB5/ZGydVeakSdf7dP3r1wbwN0O
QwgwZhQtYuKIrTTMOXCZj+XLS/tR9Xx/NDuqHfGI2ppJvi/b6o/MeI/OWmvzpFuC3PDRwjUholYk
19QxO+aXba6/qZnF1yKTo+wqcWs27L+XwA94Rxl5IcPSZvqOOuHJEHEKpuCpC7xqJ8RjdbGSc+52
UwTN4zeZKcliP19eMjJbDLS01upuahHo9fXGg631mdJIWup7LBQ2Ps0p0e75kXUc4hm5mgaKz2x3
qRye/41+b473jpWWINrijxl9F7JhUk3pv126GBOTzbRjKqdi3EmlOwJwMPxvDRU4lsiCogye/uaS
/0XdkYmZyHgCoGzBExhj9muzezDUsD9Ug1MD6FeP7BUFDBhDO3q/+jCnEKldKGtTTAZyONJMjUyk
gV/uUzwsUC2Rofed9WT9vaLmP89uWlTASnFqsODgHfTMegrmmBV3v5KMJIwCE1SUv+U4Cf33IFwV
UxbUetUCf6DPB7V5xG7xRKPIY4dtEgTl8Ut7d936TKH6D7cI+ZyceXfvJAmqqfCo142is6BqxuQP
PwZ12Ausr68zteWuNcBkXgL+Rrb0tXcOYsBmvO3k5XVUGPynEdPPY6zxfm/sQbV9+8+LF/T+ut7H
Pr/fRm5ZQSXm7kwLPul2jsUPriAhBXXrmwh/bGnB6qDUdY1oly69D6gLJ50JrdcSyho4Uc2lXiDj
w3Da31dIShTapgYiA8i/SKX0bz2S2lnsurK7zmzio8pqOuhABX84L+Qoa283FyryRt9tr6gyp2HW
bKm0gjoD/cm0xBWulUZIfmg2HcOwVyyB1dclDwjDfUieMLka6K2rIeXC3y0slyvhf57PCHnUZWIz
LwJrP1j1S8QM9OpDNhGZTreC8yvn5pdRP3ztpY2WlRwjoYYR8dIdX8NliZSqk0BiDGu+GUcqMJnX
tF/ZL54N1B0Qh0nYDEnG7Qo1KQTaqE7RRh2l6H0Pj94Ibt/5x6qdbXkOpidGlhZziuymlJ03R85/
7lQZZAhJvwseoskh6+qoFxLAmvsCU2X1hApSnBYyxzGIEj2l0tyIlBFQZFByKnvWKueIxxXK2ypT
AlvkEuNEMTzobS7Pwq0C1hixEL6YasJZF8Yew/vgPorr3c1t6SjQmNrJDSwbnzHnjdLt2i/nmILz
zsJo0/Egl94GcucUj0nxGd6MuS7YNGSmvkzcnrXfzW2HSK1K08O77NRv+cSzB19gupKno4ZlqICb
Du3seJvAOZN1vYxncgPnqTl7W4CDvBxBO7jvJITv4cJFfwBKEl0uo2HPIR56/+Jh1e7EUREZEi/4
tKIKiPjWxlXLoD2is8Ut/CNJHHu99UU7afNQaA3ymm3/1i0rVOuFbpZpllMcuFGDZzg2vP3+GlfU
29yx5vQX0eqPmqAPRcQA/pbJRiC0Bjn2RJj2ZCVXTvUNYdsl8XuyHxhnSQurPyyerG0C8V9GIs8u
qPbqJraKursw7YVywYJjM798t2UpI/sstALCQcGDD4tsmSVcnNjwluPqipqEtdB/LuawNoOWv3gZ
95tR0PVey/mgXv0sBtlQVupYfD+ZsAcgGff/TBe6E4wVZg7drOXQFX+cg2t4ncTXaR3Jf1PMr9Wd
G47ftHGBw4XQWqtivV2REkJ2BWPol/uqMG2A8wtUbGMqVub5SjIOVAwj1xKCGREl+/q3KXo7lZ9i
Q/uyTcShJqObz+/rHa4hEwvHEs+BNcN+d/+ZU7dkv2aa8+T1mJKTEDQXaccACx1a+dtKdIKAEn/m
Hh/nDlY+yDmJ4sIDI5sqvRQLUbJnJpNWLBbRV6BVTk4I/sy7cyLAg1vN6EP7q/+SO2hrPyCG8+Qq
Jfks5g8LafQSl5EdBxwxmzcm9E3MlNF4kCI455HJXbMFrpcWc2l6Itm4H7FrA/XhRJTu4V8uVuPW
43xZsMANjS+liSCeQK2E7yyNvZeGPnXrrmSCAA/2ahOUXi2bhxLtD8OFnYBknSO14PQrn3nGFOT6
w8otiO4v4/afwjolE2vf1pRrGTplQ5RL6RpKY2XMumvBcjL/H+YSM8mChvgTnQePEV4ZXqAOZHF4
Dg9GBm9laLC5iwO0e9LWlVialJEQ8Onv4IWBvGZTl9rmpWZXBqZNamLwwCBJkwgEDAyQG7lU1uON
z99wSImf6X3Ix/3YiwDuikTdeDCM+hRLuinG4yucj0zvozTpgwxVCrqvCTWFwDv7g0Sm/inFJ0FY
GeeblRHb46S6AN3VSUQjwNDGZVgpCY5ScAwG9lzUGpynloCI86cDd+eiwWsuCf+lZjotOGI2eOlS
CwnqkLVhrSqC9JQqASgjDIvFVso4MNA7NoDGtp8meG1RSRzByFnIgZeDBwxsKYQpLCurqzMb/2Am
bi0hi2Tc10XIvfDNVvaCiJdN6aJvDXu80jBK1a+YKFjNgYxtisRQJ6M/h7NTbM3B8EvkDHofAgOi
IS6ky93JT0qZvVNx3cmfEINS+YrZKkJHQ0GeYXhQKxVniKNnsfXzLOWQvrECL9+7Y5JcqZy/nN/X
yKPFqMI6wPlMFazsfDsomOzXaWRfoTaUuoe+LRrN8YFJ2lzdyMvGA728baxsTdCjqKrBB8hd26TF
1bfhdZDJ8VRW0kyGxSnVb1rAJFkJfgOXaS0u9UDsXCd+9+59SF10yp4hH5/GjoYRt8ijO1MCOW+R
mtYZke4gxwuKyvAUOaUo8TFibDCBMpvRkPAvxBos7i9R+A/3uJW9GrY3fcf+MWAHoLhk4YA1t1uJ
k+WKgYLUOnB0XSYuZyTPbCLlFZj12JgV3TK8lSarI2NdhMnto4b5SkB0r4sv2lJP8n3ui8TLlbtw
mv2QuQpHD0YbsN/DQn3M/X5XfocvgXEGtArIq7TTyj5NBo52VaD78KyKlMP+fLtVWCewSd3CmrNl
W7EzTCjQ0qOS3MznhkEcjKHCDGO+zRGflke+yClajhV/AdMDBkAX8Mtowuq+7avYP6R5nwUsyhqq
VSXUu13bP/LhxAQODeKOCscB+Uit9+RRVheMa6xBSGx1nV7rrZTdJGCFyC78G4ALstzwhVn73y19
UyerdDM2HcsoRJGeGH5vYUWEtNs5EzaGX0VJMA2g17NQ8taQd3TM8WkYnRLNeJQXgunysNAs28tP
zr0qnxMFu/DvRg/XVFl2fOr315TjlZNjjN8VhSjn0eLMjc3MsAhspEZGws9n/JRp78UdscTdODEh
cftRXPYxemIvjXpbsGEdGPQSf5PM8/U2H7BSwDYkaPXdTCKwMPsO3yt+tSn+S+eJQr4HeGG+MTwV
3swo/S/AbvSVyUzvxQrrlcvLEriu2Y6VdiZiAYfWDxTkZRxsoE0LKazT+hP62njSpPmG02KdLUiJ
qX6Xn08MR3KomiKQabjkq0OGyW+O5C/TqRyH/U3TMnpetWWQHu2KhE6DhDFGWqkVLXyIULZISYho
TtqT/wdmyLdjvCWsvHvTc436Q3mDDsstCpm3MvqdXpyYefZ1Pu1JLhLt8q1XM4HSkEI+UxIti2Jp
6D3MmGBmDdqAekDsMIhk0UWMuq1hnewC7avtKVD1zuaFyHs6kMca6Z9t84zNfDhQ+EV6WAYULjz0
4Lm+eRUvbMGgwwK3fgORZS+fjAxLZLz+AQ92ROS1WVrxy5iMPRHCFPvDVbsasGv1pM5RxhjG3c6D
FOttIuzpJf2m1qDCmgNUDEH+fFedehu+PAgEktsVy+LVTPfcZUB8+U3g1PktypJ47OEZQNTYBz28
HwJWg5wQgyjkCfIfiNlj1r6WFmQ5r0+HLgIVv+JEk+l7q1d1aIJNDpbCN3qH20cuwBIVMJq+JvNm
9wrpvBSFicVokOTLfxHmx/qaMsTyxCH2QQujFcjCZam6K84RdafFBNaT28yjvFsrBbSmSzVZdhpy
rC0jHW6ZNFCpEtQY4mk0locXDEd2xfxem3PPuvU/l661eE4ns/ZlV1JdTjgR0wQSdI3fK2f40dpe
RiLof0sIDy/XYiNbgZx6JLnulDWqMM58yuEfha7k8wgkkL0Cvm0yvrkhIxusJ5GtpQE9767Q3Fxx
xxW+CHWQ6GpFABChMH9F3VgZymzHUZkJJv+zty+c4DZGcTwj/WSGO9spuUYnJMI2j3dt790Gjg/S
hIRYATbq8Y3TrRxHakAb/HCmHiTSGDFtMQ1gSs2qLEe9/xgjLUEERiXg5zZuqHR13DBpJEpxoFx2
sZCX9poEbkii4ISaxZXjwdnR0gGEAnSjj8p5MyIgdgC3AG8f/DvI2qqMAhEY4ErZShMXKJttBjIR
K0jwWR0O7AfbdJnkCLEhQ8L+BvYw5cU4uISMrB0LoD6q5JMzmQ3VMYTMX2LvVoY+IfAlUPDjY8HW
RvidyW5qpp7ezzbfPfiyMJMHEsfMZKXLVHsJVPIxvETUi6gUi0qbLA/djzkP3T63BNTvbOe+kE4/
YT+8b1dT7PlF+5lYZxS3f+zWTwan1vx8TSOulPbH0S+9cwRcNYaGUVTFryHkCqXinVmkAQw1n9OB
C1A6zLbhZAcnEsFsP4gWqgkOQ1k2akQdmzEl+eatoGhM4dkyWO4g3IulQw11Z0C1k48ITwDrD9ql
lwI4DldcB5ltc+FbaQqcKqbg51naAuzbCmk0i6JzNXXWUM62BlK80zREa1pSulk7lwZ25Khkc4A4
sqJ0yUEGiTXTTYI20CmdoW4x+e3laCccgQCtYWAMMjRwApcdnr7Z3GK7UDM6fGNAC4DIG4BAlF9V
CQRCkZYSe7qfA45odJFScOx2I/hcR5KZWS9ejv09bbSDgCCOnuJuDzM9D0XbNtpzeNwWFRU0hgXj
EriF7N75qNVyTqE/whfgzuJzHhhFR8AUwKPMsvsbA9t8KaA0WUnz1ugpmQoLxvqEBxQC4+wPKf9I
L9/JhOpTIfbzyM9r2zZzQ8SXNbPMXqdgjlvTraFe4jTWwx37NZmzclXp3jCZvVaolgdO8a8dvu87
uPtumcnhQFkFkeRpoDdipeQTKKxrsGJjfoxu3Do/kTLRiXOGc3TFkFG9xp5FT/Opy0KeZLSX1Ipi
6RTfQQ3QkV8HfOqakX6QKpCWXp+zTrsdgJswXRPh4Fn94tFvdBtrJ3iq/eyowY9pKCN35kCMyW6q
glNQs6y7QENxTTr1qZjIrOuPhQy1yrqj5bzt63iXcREHMsZcR4yMi/0FW0erAs042idbrZLZCdpL
ibgQwMuv2XuytUhz2iS5UHDzrpZI5sZ+GxYXWvuNqF9i+SpNVi6LAzhOZS+uAuq46QnFnBkvo3Bi
4Mimx/Nv/j4kPUC6UEx0rjC0XSqqM08XIZ+Z1bLld0S1qjrh2eOWKmawk8XzqnfWB/xlin4/XiG6
w4gwZYVAlV8mtVybBDZOSJPtmHtbQBYzHDg2Mx113ayUhGuh//6HNjynKD+BOhx1XKkEqBYdjDIK
f3pengmcqIvdyGDhKNKYWLph235/Uq3eYcwxIxDwYezli/2tUQjQ+WkTwQwdQXvRTYtfcZR9SwHw
ual7gTQP5yb5cQGPYza+Zs5HqTLhSyWpLOtMDeO14NdYgOb6T2IvPLsK/hE8UovwVUWHM3/u8E8D
rrbvohmebHuR0MdJV4yfgVXcso1nttpjL24w50wfvYq9l/foDn3s93BKu8N40UbZBkgx6P1LI6f8
vIY4OKjRwtB4sStnJB56xi6B4Quz70hUQy5jDplkdVxDB1IRO43syejqcyIAlLRmUxsC3j2RdjJC
MqvRTYJkOQKKoX6Wc+yxPFk+pmS/8Tj2FdSJeGRFOL8jr2rZ3j9JrvOlCJV2k8/mWrRG1Co2IL5o
eJY20obXVnXoUouKtls867Nk/VfP2pLoY6v8w7yS0gT04Xfo4RfS3EAppiO+X+4LmKTBsBenR2U6
Ho0VZz26VS9soPl3nY/ulPJyMWjzaoZNOe88+JYJXw6YaPT8Lba5e9EWizKIDJkufS3VvV5ELMRm
HmOOJVsy75TsUVipBBVTGcxyeRaVye96ZS0uUvRlRYIuIWbzhdE+MxBsLnAwERLh9YtNRqyLZsN3
uJIIkWUEgL3dLx72wX5Q4hkpmNlBQeUfz49ZHjHR4GeGZY2nUG/z5s7gGgbnLm+4rdyB6lnnIcah
0GHPgz8kIPo5vnxSiK/lLCOi28xZZYORfKtPDsqXXObpQ+ZBR+qwyYPGf88s5Sr+2vvs7AevOUbO
LeUy8Cn0bNnv8TJ99m1vOqIYYipbN43QwzWDRHOEj5wlyP7bQVEryuvefHy8LobxSWW9Rs18SU9Y
s7VrSBzXojgkxhkjKcrI2wd9whcrXshIxHYeU+OYtVL1CAvexMDyW+u9pKc012XIM+1DhRee34+4
aaWzcaolP6SoDZjXTr7r2iBXGnyMK/gRY0RBEvY/q1lqdFtSW06oEaJD+0XgBH8VTN0/18GCMLVe
2cjMuGhwd3qwG0n43Koi5AWURbnkznoOiemVUAr+m7+VjbUXwPsHNvoa/ma85j3RL5TIxT6nHXi4
aLvbMRAHFEvABvX9gYah/D6Jbk60Wcix/a+4vuKLrtrIC/ZgT+9Si1aNX1j0BY/7Xjdv0XczG5us
nz6ncsNYCMCWaTqM03FiHfEZ5zVYB4xlIq9+ZcVjJ++JwptHOek199k+DAKrnony24Q3gU6T3ep4
ybNnpXXkmRwOzqozVm1cQP8DfvZuN9v3uMcifefghGQ7ADNuVYkb8yyAlIQoO+HnrkXhxR0HQTym
KpGTgLVKSOePYKtQYF3EFStNqaJAb5ZbTfuljaPPeGwtT3ZIeAWjHymeEOgLlnG8famSaHwCMl3n
JTiQJ8qK3Cs+Esw2EtQrbFhYiFf1l2GseX9pSZ7o/woO5G2BMPwL+XJLG8oIhKxxNP5rx5x4xHhb
l8R5FOOVExR+ZA7qoAAcXXAeKPr9cEztrdVirl8DP2Da8sGhipBjghOVpNxJ0gAkb1dspanjz39r
hGMoGhMigxyaWnAPvHoURHcTWaPuOxafAYk365gK88kcwtqWWcX9FpxbNA5Knvp9yMyvmrA6Twpy
AL1UjUIu303DlvyMujfTmAWjuinA/GkLVL2VSYlLTmw3N2Q7qvdI5VevEmglYIs4FqTLmp5VRbC5
sBJm9B41R8NgXH8+GyhNxmlzRE0K5bM3udlf3h35XbeQfy+Yy3mb96IfWiGPk5dcx5qHvI3GIGq0
txUG9aHuznkADKvw8nT55ceBhBXEs/milNzyrVNU311g6nC0Vy/lnIIpPXQgTvE9Sl1DUK3S27+a
cNtwohJew9Eb4Jn7QVselYMl4rgtOBrrGqywbUOgXddQO9s04fwcTBKQXoF6MtYE28w7p9rApbNa
9DRXTgVcXZplWb7Dnw8nth7+igZl6znP5s/D1HeV4xLBuEUl89521ueZa8UIbe1jW+elUL8iwpdE
AAe1C9VMnlCDrVW4n2aAv4gqWAYDoK0dn3XAJKtk+7ABSCXl4ur747ru/g/BPiwNDelAja4WJOmj
AMc5vnra/rKTG7sldPAwKP1of+OOczXAivYVrotu7JTjjAoxyboTL95+vujetpg9XwzuL/K83HjV
A8nOoysCWKAC7mhLYo7F2bWvcPr17mUPlvg9mJD51Kzxr2Qrg0dDJyCzRwQF2ox3ZFth4w5BXM+G
R1DHD4rxj0enb8FqOG7Jgmon4RK+05bETxnCUSqABlfmZyd1Ev2ZGXb2jeUQ+U/ZKxX2QPsNVq0z
EmrFeiIT+0oyRYuN0GvLL3lcGUNT/oC8ZX2xVjA9dBRkqB8nzH/G7dpR4FJkjqTpA7tPRm9ib6SZ
YoxwHns6nvg8Lmey3a/sSqnlOM7lHWx/Al+ZG5n16R9prgIe1ak6FW7BB1V107QEqVZwW61OGnU3
Y21LqVy12mSdrRAFvLAMuW1QDEgtF2d7uMtuDyftBMnRr+ya5Nx6TVpGtnttVGmZIQLTcoAQ8eye
xZYhS+WsLmBXERYNRAEHP5F6dODGvdEVhHnBrfjsE4S3AOpexwAstj1xtdSwqkO9YjJhLM2xnwt5
ydwaRmO8sMPXb2ClQXAtuok7JLXmPPkgviXDsRayAkn/PkY0AfkP1IyPf7xNeHzFSvFL17hSMAHR
4Eq3AoYYNXXFESfMb1LA4Z0Xcc9py2RwiVSlMBsJ1nE5HByW9UEhVUw8uXhenYWvY5ei68TByoEv
xEmlQUmj5OL4yEc2sFqbCU+gETDFlr896DRhd8BFku/xdq4jMOOBOTZUDeAEmPgc4pI/si86S0hs
b52n/AabZB8Qne6iL1QZIyCWemwiB3JCXhpJoMvlcFDdtchJgDQTnXFdvI8DXrbXWlHOv+kue/o4
PmK6GZ7sqggt24tJN5JMkIpmFHk3Soa93T8oNNJE0hSHL7Q9g1j+lasBJZ3RcxenzKjuGjFaatNb
lRJBD8C+72Z2wQS7J+pACRj261SCGy7QyG0uyJkeoveBdEncklTl2EbJh3Jw7XjP8RbXwVz7jXzX
PfTHMuVIIKdbj+2OSSRdf+sjeSh7C6OdQVtzVbr5+2T3F5ZdOgahNFABZEGWQyEDxnm4tt9A9iyq
EvwpCAHAlWGY3zU2vmCVXWYwIF4G21PMcA6UG2XeOYBbn4ZwUyAiYz4uv5U5qK3lTxJDgbvbB3UR
yVf+114UOFIJXO9Pzoj8/wJT+8BS2QfEC2YzFojKZn51cLD06GwRKsjI+8ob81xcIPtypS738YQ5
qrQvGGNmDcy3ctlYc/805V931rPck8z5B1cZxMXiHHZvTyg0j+Ry0XOVc9H5gAnf78XxkA+FB/p5
5eAA27eA6jClKHwkV5uaBJfzs6G5a20W0rw02w8xuOv70PTSHtljCPN1PKnymJTDEgS7eYAB+RDG
Hgpnte6I+WWx/3YvjEhbH9N1xnUPOEJT2VrcZ+1hQGaNbVijueeykMfERtkLBvB26T3fhucSyzLf
cJnuyA4XnlWSHsi4CrYcmhNjzUPDOo727z6kHDWW5i6M9+TY2RhIkNA/CHCh6+SC2o7MH4GbGNrD
qXHaXoSz8eIXMMs5MI8ifqVloMUTJKJ6RGh6LszNnxGEgx2cjV8FzLEQffGQew1kryn1nRCxqFAB
rKfGMi9j7Sm43e3E/kXVSDKvDvjPSoItL0tzwkg0ASkL6KVSxAVwrjJ88IEHWzkLYdkrT+U1E1sx
0/Ehj9uhwDEjRQw1pafCeFZvtFRHBUXlIDDCeTWdP4qE7MR7LbsmRuVw6rILDl+TfxBdttoPDprQ
RD430oXG12bepn5kuEZEm0gYoEeDj0Z7GphClner0e1G8yRNJvHZ/Yu4FUWc731Wafb2+WJUSgjj
bWOEWeZzk5IQx6RnXv3H05hKlYxTHwv07Vdt6fLSkBPTfevXQdTWn+zY2Wuo/IM68/wlBVJExJ4J
5L27WlY9qPKJHVuQFsMqHe5MYkQJ5HLlHhoCULbbs7M0lJHa9fBjfx1MRlrzEQqdi4z4OqEkeK1l
/7g78gaNtkRGDSWBIHFI1UdDC2du8fgy0VIKYlf0eSyPBZVLH+66R8h0pk0iMYLcmmOaeMdC9fUk
lnPHwaxgiDTTc0S8HGzeObfofgUPusOFrMLTScpX2ni2Sj/zHd0nhXDtLLcvUXYRoiTqid1HCQR0
jS3ThHQiY3pbKSmVPSngBO62fyRXj+2gVwsoUNQZ0P8Lg5fPUGGiUdRBcQEOKqJtXI4D3b+sSCy3
e9WaK8LyhhZM1tfP4uio7HjcAQgTzG18LrkBCLiNqC6xdbc7lZZAd8wybd+nG78zDBWjC1vrSFcy
Rf7b822Dng3JiM+fZFdQWBsETlH0kWfnPc8Ldz07bJ16vCR7CqRTvTglZjg0jQHLJPqMgD03iedz
atq+8Ea0C4R5oka7WF1TRm5joGHIxzeY3C9q0BNFWxqY2tKKU3N8vk1BTfrzipQqCkS7FvkR1+3i
7giVVCPyDjpeybUY51sXgigU4bZw/s6RRAb8mvVNbnY94qqh1QlYjizZIIzgcCil8O3ZCaN6kVhU
TzpsRoIjyuXdi0WrzneG7A73jW1XEAVqOOv7snqsNg5i/jSeX87tRgQNfTXXaG+YuRkgscnOjxf/
qvaH21lX9uE1ghU+kDhg+//aWZOu4enjEEYxPKcIBeML9aBNHiUoS6JiBsgp8SnGORKGgeTyxuF1
ZSkYv379DK/Rk8JcMYbdg3rxc9gyNLVmMiuz2Ry4+HzBEn4ZaFv3y4R96pMq7lA73liPbAxfm8Vo
+waHW6Qw1LDgwPRXmXle7G+r5TtAwrcZGMoM7RulfWgDRGjpfkDxb+RVLl3Own0Tja9S3EVoks0E
y6hByv7nuPk1FNOzLFArfcIehDcA3R2DAItBE+IdyWXwqmvgtR9iOsGy7tYXY4X/Cw9eBQSykHMx
EbAB9wv9d+6jl9IqGCDLFbiRuR8w/PjFOwMTv98Sn4SKVVrzj5+2hdF9DWrwvLGyM4DZR3tCymyT
/pB7rluOd6HGCz1brQ0PfaBV2HVSC3bYCRtz0Zabm0pApH9LF7Xx0eMEhZ6CG8oDg3yooGpTuhxX
5zQibnA5v+8cSyOVDpsIFg4S4INIF3Q4x8kgank0e5MLMgRkRmQCQdrxhN0JdyP/OgNGRHPxUOpm
7nL7X6h4VDNFdNK3vT5/efHwnMAnPcu/gGj1q7wEoVQTTgBcc4HhsJh72+M5j/tmdT5GhfTW3gDF
LwdY95Apvt/ZG3UWQz2/QYNru053PDW4v0f2albFk5VUN3UMhnbxsuXV03wefRjie7n+ZAAFSR+0
1MMdr6JgIHVG+crWVeu4GDRxE6By97gU78caA/hzFuclUAvgGBLFQzn210dkAZFRUWURTloec5VT
Otv0Iyy0y1PyLev8xhCzhiYDB5CG/NL9VQ8RnDKRW05T100HUTakyG3X4VE/LQqfwRutyrQWHVdU
pFEkZhMForTfR2FVXL2+ofmoE5N0TnvLWVo4r75O/vwj4WcTo/Ox7NW3R1EGz6I5yR5g1K7EzxB2
9AzlkHBayDSYgQY+VXlbnqcrUyqmaZ+BDyPRjzKAlF5ZSME3Q3gPFO/iUODPQArA2FDB9OWpAw3Z
ZiutTHASYFKQCEd3BARLLIyUL8MLAQxD6bSydnJaEngz2Yljin32B3GU/ho3KGmxzKkH/faJixfe
k9J3XVmnxf6h0+90vfR7nQxJcXFCdH3FeLnc8K+dv0m+6net+c9m6hNoJ3ty0wBUKEp0bY3GdGEw
BRK0TFn3GdCJkum8BCOSMY4kcIU7/SYrQbMKrfnbwdmk4+J+wJnVhIznk3R3LySkekyTWS/gx2Ls
zFbFHj0BvI7iqetqKYatIkCUtl3XgMG0wmsbwoH2qfsX7mTD0cj+g5oHD3MsUG31GBpVtrAjraM9
yCl5+nR0eZEon0MqPCwiQX8RBO9fDinOojstygXVLDSQKP100zVRoaDrVs6vTnaJ2Beicbvcle7k
BtW+FHUFR9Y+SJpczOaiZoadB93n+dTjVuWdGI2dfwp/DvZJf76BSDTUco6xwLpNdsKUmBugQPAI
zdiYN5P9l7pgVgU9kn5bRd+Jz+aOZjeamUMeBbE/y7IcjLXDSnsIvFVWS7piVhPJtYJYN3NdtyRq
PTIyEXlWFs2tZ+pqbETkN819rHqDvNEWHpJuvz1m9l8wvSD/Oy/tBAng3kzviPmHOZASDIImnSGi
J+KgNslWMbePP1PMaw3ek0Y2o+esNzdVSXE3vXVHkeo2q+kkvlI72+mUcRb20Y3MGZ/vGRyEymIT
obGIsuRl4Fw80bb9DRWziNNShF2aQgUaXSboABJlePX/iVHCrE+wk1cTIeVRYfpQE9vIt5QPHlp6
XiK90tLBZa4auu67fNzBVSP8eEtOhJg16K+rEYcXRTjgHH5GDFr2HRxgULCLAC6TfNplQK8l+LGC
PEHArhb2MU7cNhQCnqfSZtVSDUF/1AuFdC4UUqeQAu5hUfMJLJJuqo4k6I77hBy+wDzKMr/wn+Oo
br3WQrkOg9s42G1x3MAhwg8P0qUZKtu9LwIKf5IQSvNBxy1MPQ5Bm/jUY3Zxx3JuYoy/Tw6WZ2vL
X9i+0xwmwA8ItvgeyqpCQ7gmL/ihxvc/8zEYEnczNfs/GT8VaZAaUz0VvGLcyuUlSM2Wc/mhDcBZ
fvsa5X1ecjuxJlM2I2FPtsLh4OiF9with23c6gBadXYczfqwlfJ2AtRkw742ibWjZWgS0lfMWqfz
NqMzrkdCxgsiIvlhXGkAljI8WO79ISTiPqL5vCBWJvOOaC/spnxvtUbXBX83Gij+6xman6iAXG1o
CpY701shiASVW+DKq2K3rlPVrAIkAF9glDpMuK/YhrcvyWTajoqt6jUbJGh6r1DXnOe6ugUQ3s+t
DBGxNPXMwGCpX2noeMMldxmolIQI0U8g8+u37SZsWPpPh1zil8y/kg6uXHnKXvUms7wSKZrV9dOs
iMw1i7/AyDe+jyCDOkpHeXZL8fmfCZEwr/vPEr03plUeeCGAgi4Pmi19+9UNCqDF3650kKRuWfys
AdGPqiQyQoqmJuOyrKyUy6eZAFG0ooSouaeizhnC+ljS759RWsBo/6cNrA47VkFfjiZ8+2P3FO/c
sf4e0HPBlFexC7e99uh0Hi62fkLX03gwdkeCgjNbfIHFYLu4AOOWyP8ogeph9G+Mnp7kDOK3XxrK
W9x7rTl+yGpp67yBa1d3a3FiWab2ViH4xfaInLi0fole3unH7wKn4gu3KezbzpFE9z7WU/J1Dnte
Z5krUj1x29YpW0N4Mm+VJUAOriCFmwNi5jm3tD6FryYOXsyb/XRTd1oXWJzUpipimXZ8/PXoomjP
iFhf9yN3qGkT9tD/zc5iyjNDwIGT9Ica1aIdOXty365xFRu+k2fLm8u6ImMxIfztj242ErWTTgJp
OVJIMHOCWckHdgXseZiQWh7X+zlyQeDD0Na8gAIAnXOL4xBD/XxzhbWhFBTgAbfi69u3MXgKQaGm
U6pDdbqA/QKdAyGwgVSMxKnW4NFaZ9/uW5Df+fWy+sqCUqE4yCr9lEFyCR7+VmeLfQbk3VlfXqzT
Zm/tpHuHQjns7xSStw8sKWy0Ctubhm4Lf+y/qNYh7JgIs+x+k5C19Un0k8BWh7m6kvS7uhM1Hc8c
fdGMgZZnI3ypUn9wCPs9BMHy3Wxe6cFpJ9oGN63BjVcSmG8USs7OppJgxNiyTuhZDb7v3UVkJjIE
fF3UDY9tCAclF1EnOVX3TfqZ8NuDLrtSRJsrCAVVFV8TmcJByLJ/qDNkI4er2d/tvkmlkmoXmsv+
he3yOShTBJviiU0uyBzRg14qXYcmeyuTqwQxlHaanCVeJUSK4bGH8wyRc0U6ph9hOW7Kl+PAFJ95
u7T9Wx2vBR1CXuVecZM3nyEJAkOfbg6dsuCKn7B2dy1oyEBZ2Ka+7nabHMkg3PAUAWMgQWjLEXeN
c750axaZo6SvIGPKABxLZ12o6uUXT27YJqOZCqqPCYJCkx1BAmwmx7Oj5AcPPrji8wl2yGDgaTET
eBySverm+P4I3O9f/ebjDqkbLwqiycU5PqDWZVLqzbdxuuWwonEvFodGAiacMiMB0TH86EOrMPMC
F5PAxxDabXGm73JL1LnvM4nINjBhdymulKWA2DZLAUTtL49/WgJdCW2VZRvXy3RsNeeSxdH6hLSo
OBQfZcZujxIRBZok5EN/pZBSM8knpcSBm8J3CR7DvutFIsEFDM4Robdxel3e6ZkZFI8iLA9r0KWW
x3YYm2odIVORFtbuW9XAMe1Qn4TqjXV9aKOhOwa3jEyg/Ayj4o6oIIgqs5q9HfVvh+Z+EOX7DbbR
sgNDLBoOg8unWYQPnCjUckFbnDp02ySlpmIorKEVRI/tXknli3MS8vbe+tbFE5UPyT9fd3fcxdeM
AeC/PrEx+dVhllbF6gdKhTPV81/LTnntkuu6/hH3bdpjGY+iXGp0QgwdSYoMKonJnkKJqZv3x4Wm
1ILmDF0GEauhhAlZPT/Glr76DJh0+k0wWD/vaIIBcVE0Q4q9SiB5RQu5FSphn5StVzc1uvLvu9Q/
cufTbkr3Osv9p2/dku5RMweT3KX83jgMaXDpi8DK6Lm6segCPDyonA2843JhIh5uDg+7Enotz5vt
sOeOUSj3wWfi0lJSIUWNGwmwmbJY6/TSq4eO9Z6pgTyo9ytdVO9SjVJEmxqOvxFptZ06iryjTD5d
ZkmxAcyD4QskLY00bsp2lcHcGBj79E5iNHTue/rreGDyXHyY/+ivaPk/KAMNEcpM78DS1AEMrnUk
RXIeAoBjxQdyYxQXGNoHTY4kGGgWq86pLyv1gsfzpQ5h98kHzbMiC2/jTVIw9MD7QyAALHO3NnGr
36D6q0DofesHzRkxhudSfpLNtU9CaxnWMywUslwXPaCgsRHcX3w2yPzuKGQf81I8kOcpui8O91nS
QM1O+gI2LiUD95hM6T6vrHhyzrCMSZUtfeMBMFLqWei6YDUDR1hu0DJmAxf29jKvvqXVsxJH4S4a
XwuybgLFIJtCbmK/o3tk+XGvbTb2AW/kfwOMkpaxA2dcvj8Z4UTQ1V/SaJpObMNQewG/iIgk/2e+
MCleEuwcWWu9koEE068Krqyx3Rm8iebIm/MlneI3fsgLCUijk496PqXd5490zuXdzXPdfy9QYCuN
Xd4rE7lu4cM20/idweDfksNSb4+Io1SDMFgAMyfGOdzfUqsJRIKl4jReNLpF+DM++022Csq3FQbz
kNZy7ipaVF2S5q4qoR98waQXu/9kGS0AJKDOuhuunTiZfchgBKtZh4x5pdgysCY4Esx3Yrq6Q6Hi
ZVsEm7sJrmcMRpmfOEUNgZb9+moScpS5GNk12nvTXD0MWLtVSo1Hu96I4nqRuP1Sg9TKEP4VSs/R
jZ61NyOGUNNpbyA60Lzm+K3kKCDFZyibbBGUJsAXyw330J5n5+z5QL/1o6Gvx8iW6Dy+i6UeeGe4
Yp3CkuIOSVxiNCkRxNvyPPmkGhk3Hvy9jlUe1eJmm0RFmU2/ZIqDHUcDzgsLtWZqa5dxSQs7Lr5I
we+JrL4ZZpo+Zm/S8/QHVh9WSnlUqHcfR+IfHV+OmecCKLGmiIXey/Ga1zyu7RpMnuOQ22MwFMnG
keRmWYQjSyXLnwwACkvSKyBj2R/SXRtvMFTx3mkWEHLxv0JowMB8oDRScni5GWiZiT7KUFxuxVhw
dPpqabhpBIS3P9IlV0+Hwdn+u5XzASINs+zQwlrI+wdXN5yqEf0AQPuwfEk+jL8beLEVzYEz1a4n
Gl8y7x5COjNRaKoGf2rOK+2xzJYQ3fOnewLCuoiAmP//3He5Y7E5cEpSG234n4Uu0N0GwpmbJEEg
fBu8DKPrOW71+gzkeJVS9K9gRtcpn6vN8kZMx5A79/qIyj6fT5aNqmpZwnSN3s/4dfuxgwoXoLUS
dKoYuP/co/CgIDhRkk7fpJHyD3chYBAZ4VuPeNI5yJ2ApH/J8Nylk1v8H9geKPyhQBOOZWols+IC
/5KZo8sguYhRRxNbJK5Pt5/6WPMbkG7giOmkf0aaInW7DZ2ASVHtlvJ2xYXCe2iBq8vs31M0ks+T
HjAuGYfkPt/RbOakKEpIpZZKunkygW/2y2pHpxG04oA8fGnvsdD82L4sWRyG3k6Vj1S9ZmuxdAj5
geHYlp4K/+P5Tu9nEjRifEa2sdENyS9rDcRwebxY7Iqo+8/dWuq1RHsFdAaqS3qdKZDXT62kynQe
GEuVfiEyokJo95jzC0hPfCprvq68iv3XQ9jRU3vVh+/pzHP2dld9Mb8WmyWzm/3FONIn2AzjiIW9
snHMwsbTeLDahRmEZ2BMLtNCVrXuM/uxlGwa8Ih08hhkVZZdLGjKYMjoGn6Jgq9pnXekJjqGnolX
4wzr5S3JPIqcE6nfHxKGPz7uhBtdjjnKXBZW6Y/z11WmIj6zUOShXhJJencxQDXW2WFdw1q9qq0T
hKhoethFQ9OF5Whv1Da2x4AoJfr4cUBIjPGNMwY7EbFX6DGKUv23g1taxH7izCirLpLsIwrTGJyE
4TnW2sgDt1wuNGnZxm3D+Cg3PxaAO3dJtblZmleWs3bdqW+7I/IY9CteOzig+f3GFaRbUkiG93vM
S5i2QAGCQY/dhqWRns2NvTt/85GP4ls1pTXMEWdBXP8+dU+26nhx2EGqk3bXhxS3igJeIDDpoXPe
gyviESWKmUVvBB9mzqlbT7JRAV6I/QzkAjBCE+dXc1D+RrOL1CRASyU+l4j6pDc7U5YAPuN7TR7Q
z9n8gd9Y6aiqLrCCZFMkBjoY4j2jggyVm1507M3Nv/BeeXqtKPiHCyQ8GLE7D9Tf/8T1Edrv+PX1
zt+/lu047246kuBsD6ynmbWAZEMR6Kz0c9eiiwRWgG3bHOPMB4dR+d9I6s3p56FYwkkLZj+RDqin
ARA+p7d4MRpg5icAYnHuyitiAsVQygsaoMJNigOb2eXEM/aDcbmhGC8ZtPjZDy6JZt2YFb1WfcUl
F8+8r4OGYN5Gp3Vb6AZvfoEsVyKBZzNQAeL66BvgjktK0PAcJ1hBc0E5jWzkwzrv2n4tVfudYytC
YH9pedTR5XknLGfbsB/GqpsUUKt3wzrK7fH+Tz96XVD6m6D/gdZXxN99Wt2OJRtipvuh+ZwebEMt
j1nP9aul6veraIh6qG2s2DIWNUU98IzwOqWPO8JYKifhEThf8jAPVSmIONpGrR4DEUVzynN25yP0
qCFifroNxgAQIPEP0ivdm+zuqBlhxOAuA8BoFZt8naqV6t1JMBC3t4dEntKt1gm3Mm/T+Z+EakD6
bpkkOjHOnAI21oN7rSlVOPJyoViQn7XJpuwIeLfhry6NdH3mLVnypXEMRbMCxRbkSu7BQWR5LaU9
mfSFC2C6pJHSCh7Tgsu/jQYzd/3IXBBJqrfg9tiwR0SD7BTY+4z7eihZy77EP/es7gmakug79hFD
WD9zWaBB85pYzbth8uZjnJqinBVbU/XCZgn4eN/Fkcdt/u/QLRR7x2HQF0dk/97/8G21q0988/Ip
ud2bAXPL+97QXHpJRTkARMHJjHc4Th+LuHrRpz2+W388VbES58FcrXWM3ajtfc9cvQMSNKkTsn/L
mA1/iqrzkwOFYkSsNJIQD5OVsupzU/Ibm/iUt3ENnTMLsqc3EicvWkIMFYmj2c6H/lxyZFvutZNC
fh6GeFEFN6zFz3RLWbGROPOyMEreYuPpxNyHB4kSIfQdWTb3qofMA7l0oh1EH8aC0O3ZBwlvY7vd
OOwTf+3IdoQGPAK3OTTUjU+WCDu33EJNHcOzfSs2+9f+3ZKYF7KVh4Crh6nINVmj8LoD9f6k0vwP
t8maRpQE3ir8AGQg+F1u2JBgquTY8RCMXGVcr6xM3OUyGFxnx6jp3y3C/hOyzKEYhdrkkaq1Ulw6
RP7gmHB4KiRNfF+GUECptFiJwf1cz7ztickpwIVfnM8ECHqMLfR25nVY89BPa8EDyeMsKvN5eNGm
otucXo9xKL09L1N9nTDblUjpi6odRkd4ERC3MQhwEO6d4s8x9TvqPKe8n/egBIl3raPxWWrumUih
PY8kvRYVdJmHxl4JzPZm4pDbO5To9liJfE4NoKDS/g4SZwPd0v4YhtUuyQKjFrurMU/FGjpJ1TmM
Yk2gkvE5up9GWqOzzNH9Xmids2dMTSKo0qBg3CWDCryuz0Xso4rtioo0kMhr/IanZrnKrARkhQqQ
UOZAyrzS1hESywfHuT7x3wSbRS1XTk8uD92KUwZFqYS6eJfq8J5L1Fq9uQwpXTwZBmb8Nhqoiire
InEbn28kyBaqJYfinYa7uH+vScTqCn7a45Ba96oDkLzWA6osRgadOwymZqLJsZd//X/Hmg2cz/xt
Y8AGJeoE9yY1zRq5THCFao2/Y4q3LbdD32fAKTy4odScxJbSIHnZ+mZsOWt6MQNnP2LZ48QV0gcd
fsPn8xQiU735keeMM3zXLWEihl4/1WqVpIDhUOf9x163V1jq2bpQiFVy+9PO8QkqGKsTKbacn+6y
LLS3LhgKQ02FM+GAlAvPCJj34r9uCwV/U8B4/hw5PzYNlrx6z6KdBaFY3jMzl3RRzM7f3ldjjHB2
c3VUHMVn2+4WJBJoO4gjrpKPTGGMa8KQb/R4CAl7w516+chHLDewmNkHdiEcU5PLUarOLaT8VJ3H
BJERx7/6e+mm+e0iSrhzUr1zBpCzxvbS719v33pakEnFtjeH/eaaD5iHuRPWYINCuaVT5vvZ9zvu
zaMYVtPPDO86pmWpGd3ysdYXvrJyjwUdEUQQT5wWgBYy8HIuZIJOAMzbPNb2EdtlYg/Onfukckhu
GR4RUCyCKYDL5Z/PcIFk7CuStoHJZTDZBr+XZIqZzqghzUgG+65mvHRZ6e3Th1CaZE07RU7dKFLH
M4O0MCODv1IHzm1zxigmRYZcas9DACBPbDqzOZg1khfYmGQzuB16DNbfVvQdDH2OcrRvUR2qoH4H
bpzduYo6eshIop992Jok9umQe6ufQlnwao4tLQKQ2Bi0roaoRDu5tn0OGIpadApWcTiVeWXfrHYb
A6QFusk+Wu5UQjIVRWRGxVHVMNtxLA5aF5lcThzcrMT6aaThFqjusLWkKHPfHc90FYIvWKqXhfJj
PA64JBGXNupNCd9mEZZwzfIcuOZPYObLm/dsyFEB1HAqvRtmck9jl3hnwzVnfV4wRRT/RYZZ+0qn
tHfkP/CuRJSUidTG1LbbXUiz9T2fwvhZmCbVT+KpTJi/KOAtPu424hayeN+DhXVGLtD4eHE6yRYW
K8BcWlyuFzpEHV7lkD08L8ExKr3LVMcRV+XZeZUuwJTZzxCH99RHJL8zVdKFooU0xtfi4KdHTBCJ
uoWHtDuRFaYINc3i60Poqt/6CitU5WqQ83YcniRG5R9bxeaqLvUtWmFAf54lgA8MrF9jROsF/5vO
HfjnMZC66Lk8VCnTUVa5VDJ9DhFZ0iqN2pBSj2jmqjc/Yr1GIIoTGislS8JXtgoyy57Gj3n7xl5U
fC/8OhpIgcMhF3WQ9GfyqHzx+rJJoe66TaLPUqt35A1DruVglg9r5N7eYH8unPkUdJADgOKHTbxJ
s3BKClQkTJLDUh1XzMr04Y7ZKO1GXKEJjyO0qL8Ji4ayFJI7MbKbDCJVWknBBoOI7tSvrfNVXSkW
Xb4HosH3qlHeWtIj6Bgw2u9dH4w6PkTsi/cXHElBx2P+RLTEm5lcUyveOiFMyL8DapEjudLbhFhL
zV9tY1MMW1UWWj7ZHJv8xvrM/tFfvYAEmHFmE1pXDyK7Grjf/B10MaMzL+ENNGR+rsASVE7QlPwb
+5H6C8I7aNKbIL22DRF2WBgAtWWeHaQEVgyuYyrzWO8fMNWIQFKVYGjmAUYJu1wgQpQImF2L35rm
6QInCu39eErQ+qmxrg1vGc356bo6ShV8NIk5hKCrDpvpMykmdf+GfQx1S3qqCbAUdxeaR0ktnCVi
Gis2ZkzXdDy+a9DDNqNfCgCj+pR72yBPjKwR3uUmmYo3XN6x7QQlY8pTx+hy+taJ8m6rHGJ7+okK
9C9WWqPpUe/o7EiQgekNvzdvszxjop/9Frv+fl5iatu7rxTqHlcQkqG6fiiyrv/IdcRuZ+qcXfA+
J+MrAPolLr9PYaleWMmgJyDNC9L9OVIxW4jvgzu5wjhUkXxKQJBjSgPKyFhbNZxQ5YW9MZcm9n4G
JomGDnVvQ3S7acvpmUojPjQbZ0E4h6aA4Y9RgDWc8UzSscOKl+7GJwS+bOec9HnqgKoZMLPswXK4
pamoXILx5T7koCdmxqCGYVKzmolA2+td8lzwpVF4cIga1/OxBAkvrHf44EFZqPS0T9qncu+stcIB
V4RizcH3ek9CAFJ6NQzNEDJvL0QMEIk+jNMT2hWtBTxRVYHh08JphUegIRy15XZ3d/W4f6haVe9y
nsM3mnNT5kjUh2Uj700TTBClfVvdhy5JMgHoSfY9OizJ/Du2ijtmLp4/c1IpqWyzXJd2sG2QMRvb
MYp1WEG1lQQhn8ljdlEmqNJR2I8+mWsuaqvkRvbY83TFSNTSdbEqlNAgMoMJawo3i3W/HUr3/6Le
GFPAVj4noAYVkPcy/12fgTPhuKoLt7N5RC0ny/PMZdLouJEdszDeAuH/3nqJh53rX0E0dXB663W7
V5wlylCkYogtHj25Hvrzuaf//wwIqVlxPqqLjdu/J96xOI72BZFKNpx9PbAXm6SMXH4n7mmxUTUt
81ymRuxenFYafubcN/hUD0IYz8GD4ij/SU2nWY7Me1ReOPQKKs5zkM+KWTmJQ0uSFN6rIRnKy8MI
uFT7A2tFaRmbzwdfI7MFMgthO/BLsgtoi9q2EoMA9aotHFZ9K283ffEFK9nFSfXqNULbhi/ZghQx
DhbTOVdLXnPV7W3KqUiJbSqynIHHDy9lWOVIWPL5qRDLyrFn4E7v0kFMUDBf7PHofURstlvFNpTx
0I82RtR+RRu7iVE1NqZ1SB3fQu2QUZ4OfUUHP6mEYO5P2V//LomIFEb+6mTswTBn21pvrPfgEQ1+
/pKjaxc6cgeNHFjtf4cbyLbDXDF+8VSwK1ZvhkjRulf0pBFP2opKg/SWChe1pWC2xBn9fA6M00CK
jM1+9cfszoHVJzHc4LFxpF3gLVIlaaDrN0vyzAqdNDV1fpPeD+vVbhnlINGoraXfA3+lTkCEdPA4
VeAhmFW6gEmfKTlN3iPMBK3jRF1QbAKwVlOL7/TD89ADtpomakrH5Kbcl8O3UbX+GSzgc6Za6bGE
aLQNOZuiCaf+8iUIk1hFAaTJn0CyT5im+MgZK+PHWe4YsdSDLKTZZty22qXfG5Puzi+vMESOoCf9
SrGSpSCEpF73dzk1VFkeMxtynsi2VFJoX4saM8RTiJpzQmc00TxJbi29HXrC9VAxSN6NJciYyzvj
zp2d3U6co6gIhfsvSvHFCEVr/JUx3/Gk1keQco0c3Ut8XZUrFUZ1EGEiPvafpVHKQCrxIwp9BfNx
/B7ugqbzLZyicDVClm3FyFpeyxWK6ZaVpBSs0KQYTMJJZN7PwqpdL27sjSpAlwf7PaghvY1AtBPV
c4718s11Y4dCzbx0PZ3LR8+I9wBE4Q+5XCZ0UPO9G/X3d292cPNA278nLcgXiUqqefBodFUW4Vvy
mzLt0IXIuXk12WXJxygscTnRdSSl/vp0l2KBe3WOhtPS2qp5OMfquH1795sAhThqBdvvgvg/KfnT
6u5OoQiQqOI7RpKBkvCbo6J3eEb33aXLI0aIK4OopYBWxAUqr1HKREmv1mEchHQTIns/3EMHNC6L
/iw+FI3rzVeJG7uk+r6irTAYXIm9daHWhmqXnsqens4lVBXwK1I+9IwwWmIgLzfYbzWrwZWTLEHp
LpaHCgxYN+oHtcadaa7NNL5J4GuCw+cvl/EBiPwIu8plzO8FUpX24bIUdyiU/IcP4uTsX2ZB7cxz
2pT8Tsmigv0lh1NatI2+7K3vlxNnwxGCdZos9jPHpFMOES7UTN/ARbXPo0YdocoOYjxhFm9H+e7f
Z0KFPDOsnALDEuLwe4iqZ606wGe5kmjyY5h18Jkt/IcrM0eQunE+3eSuWKF1GugSb8oWV7egV3YL
hwRxuZE6J3G9OjsfzL9tdl6/148FWloSiWkDok51AwVS/WjKLoL+JZ5PECHLmMdrZRSvPiemGzHU
iXTJ1qZ98aEy8xARTi1F7aOwOyxiQCzR8zp/MDeidO0ChfTuC1Naa/o50qthZJBDhn7XXjWPQWMj
gd8XbiMyuYvFSsVf7rh80nV/mlL5efzU0LOlcZ740+ew3pHgfEuFk7rnM/jUxNexcY7ZJu1gETH2
JJlErsQwVgtKaeyUVE0bRHTb6tQfMja2wkL+8/zBbNowrBJRPLEHntNTSrqCxL61aiWsY01DoD3j
EeyndaOIXacDLotat3tFBuSQiv0alWeWH41Z0SW86N4j3BFAYW7St+/456RMInfEJiG6d1HEATsa
ELVaKMB/dmVeBlwNCLg+fmEy5PTsc9DYJ6RIiDDtrCIAMa08lOiD/ndWZurBEkL2Ca0K6G7bSXV6
ceez/JbwZQWp/eIYQwzZq37fPv5gJmMGQl1wxtxi7hL0gCXC41+fJ2hfeTisiujzxcHOc1CuriJM
4dvHkK4DrQ8a2deTePxEETMWz1dlpmcCo9Howg7PIPGOnNN++KWr1l90u+k45lf3/L9iZZI507Kt
zD1+7VltUrMmI7Epj5j2PR2Q2IQ7+u5IhCHP3i1P4QM/jpk9PWXbWXufBE4xzSv5YZnUY8nG7qso
XtI1UqQZvMFr8VwcF1WIZ8Vb6WdXWKeiQ1kpYdK+GaKiAvksvPJvYnqL4Ldf8eGiTNwgeMOjLMTZ
TJt7uHhYm8P2VGc9xGY9pS0ny2evrAcYY/sols7Tg37r8GB+tdMwv0cRkiU6wvQhk9qzY5BdJ2VS
GB7kZUj/KmyeNy//sy8qqZbsdhgJSQvFz9hKsz2wmN0uEValgvems/YnhyiaAm46Ol1maFKdHpUr
iJiU6IpSBhzAP+sI9CGsFOxWrGVZOyN2O+BAfZ3dAVN/nfftJkzDLyoPYJXk4sDgKbZ9/ghp62oJ
v7jBgkjqMQVKkyxjmcOxGCWUkhbi8GyB9YOBSjjJd9Ejf1jMlyPdBKO9S0uEmxzaQksjfJegFgbf
oO9Qf5e3Cy10ewHq+f7Szcvvz7VMVy8IiH0mBM8JyKE6h27emKg+y7BYSA98soQ/YUv8prhSiLab
4xEuLk2LHxy8Jmg5ANhSE5jeR1wVVf8tFbQxzMvG/zI12AAFnzswn4dXbZl3E7qskvQuCtnBv1Hb
vwotWmUQ7HB/WaWKM7bh6ZgOWBWq54Ca9ayQ2xis2HDSVj04ex/ihvwVAVgTeqZr9E2+4Ubk4F1r
cQj+9ZtEMOesKNsdTAoQB4BalMuwoTDcVw//98QqTbHTPj/vPmcZrLuSKWoq/weiQYoKHKQh/1iv
xoxZxlK4kTNqV4VAPpz97+HnGqxvZDhiS++Zd5l1SruFh/SMmmXKlUxY+p80N26L0w6SkySR6M9M
E5TOn4hZkaHHBTGsQU6kUdvsEo90Dg99MWRFgtXt0IJK05usljvFps+iWZ70Bp186/z656yOJfTV
0SHTw6y3RSHtWbK+4mRWmbvTiHWt/dgLtEtP1dZC0UN5hz7klF53lTBP5p8wh0wvawQWHXTGzg2c
V0l5xc2xhKb1jVIkKvfSWi5ovmkPLKYQDGWckGp2kHGD6pOEbeJ6S3zs3osTBVjTsaDAkl+bI0r1
z96EIT+HCCvyT8grIFAKLTNFFAbkdsn0X8dnWT6TObpmexxKVjlm0I4FCDjDWOopm/dGqZexKwci
/qyhLMWxUIlB3K+xuhaZAQX5vLi97/88WgD8OztGBu/JdigaxTWIC0KPksym7Of1if+/uZsZ84mn
5W9VmwA43b7Td2n+TTWPGRDh/steJUFV+VD6TUkZ9bm/zhiYHpeky5vqnLbFuPUNqonw4d0Y3J5f
q/a3Z7e17xRO21O2zIOJHdo2EmQx0sY0r7akB/fp1bsddxecJDYnm6MsZwp1YZSiiYw6okkbMPVV
A6TUMMOZq+KU/P4S8K6GNajcpnnl85rHxYAOsfd2NOOpssSnrqQLth1MJDTqt03WcQNPlIPlV1Ag
IkancCzU67Ho38LJL4qXWfzfAq5RXpVbfUfwv2qfB6Wi7os5wZIuYaMGd+wvMbps+o3AE8yimmC/
UBgtg8gpGW53jspvFQzWYM6Po/Xdyi5ScW6Mq5DiQKfoo8FX+4KnAD+dornRd7P0+6ftGrUWjDjH
67sIntWjyZ7nF6JiOJgeAW/Cqwtqk8q7p8me80w89K4cSEUySTKm1RBDqRK0kdlnfMNUOq1VYohM
n8pajHDw04AzLVFmuTiTs6HQBv9ibKSxEqssG8JJjL/0+4vtobeja85300kHCo5w09RrF3HvJ/9f
i61XUryfyI3YUUuPk4VLJrdjMNEMDHuOvr3dBM8Kz3CG0sIytb+eBVsGK8/CVLXqUwWYWR/ay9Jx
Z15Fh4m4oNKtIL4rwo+DoBDK5dm03spWlq+HnV1KXOtEZDQiqmUd9KHOEJrCbPbqDSkoUpeq7722
Mp78ALyglHcRzI487Z+YKW8Ulzy10K6r9u7d459KNgEEqUfeTLdfXFgR8EmjoQy+oX1Y9+reAs8p
7mC2FNp9bG7OugwTJeVGPTMZo9OKKihJCSGqLgNTfTWjbdFXAXjaVGKie8IOHXf2zJL3AAIuIHjt
anBk2Kafi5A3CPNDXhOKdvXTpNmvt8UtdG+Bcf3sX2N2qgm96Ufa2++42NXb9zrCb5x2pmcIQdwF
oLnvu2UbGDvheRiSQgKh575tMjxInr0O+Rx/82nD+bUwII+AH0/vQVwlGad92ngKCqn53AnXPE9E
UiMbmdGuRfHNXdBTC2GD6Umr2OODWFc0K8g9DNbZtde43fovMPaecRk19Q9tjf4t59b/qxaFkYT9
YUyfqlkW0l16wvsajGA23qpktcJLfFB9jmK/5jKj+JiYFKhPyA493iIXA7/ydPKE2IjIYnfblhdW
BX7HPuZ6D3aPZtw7HSTtZZVBecF3CdhIVEL/Tr1c7/omtmozSN+ijPzavWX0nlm6jCcW+8lwQLzQ
8618k/ihpgg8aM98R2FHIUJDsaYe4S8xNyeSThtp02FZNnjWUYHZ/i+7hqVvnzbsayHFsqtWah53
6kCfwTXp6X67ZK8W/mQI6rDBhHeHvDa1cJUm3HcMi22TanXJQISzYsT7hWWHi+TEzaItilLEEztm
3CdN42b1nGDSqODgV26cq7v8LkNY4MgzG1ljQxxrsOk+LhpsDOwiQQqnrxwXFX/kC25QN/4wrpaK
Xg3QodydKyaJwPaT0DIU1j3cNt6aYCq3B/8e8iHJC65JckU/Hake4nzn0v2c8ZZWEksP0Dhb8y+v
6q1y3DnoiMOk1Xy+aV/j3Tlove9b7PEyyTXkm2BArJOnm9TmJzxzsewQyIaqvtlaaHjWEzGIpP50
kSquvqVQnkwUO4TIUKGvP9uITTsB0MAVL0M7HnU8lRCQgX899lQykCREfzBrR7gVvWXxIKMf1tft
UyaotCJjfMXcWze7UhZYA27fMJhGxgbWFh6FlYgynF8DSywTmbTxjj3GgkyLTfRpbkVUpixJNoan
HEd5EHK/llOIpJEbuNIXiS/aEnAdZbzdSRBYYNvIvRSlNXSNpqCRnof6s68qzEmKboTkkSpD/9Sg
sodma9pXxNOROGrM752BJ46HvPY6xeyTM1OPi+2pExl7mAijZgVAsTxF+TmHibu3es5QmgUMcOIC
ItBNs/PNzIT+2T4TnvGHxOqW5hFd5US/aUE7NiuWgwRlM6+qLMRsgxcQA6W9aZbTfsSU9AcuckPE
JggNS4wKgHU+wQir5Ttl7xHfkk6GQcFO+KLRD5BrKyqiQ4zpxUbJB55LZ56MXdGdwFW6UzXYoiZZ
ltKQ2LjqZfrTyEGgtErWBLBFrRtpNIZaSyBqH1/wokOBT2j7M79TCJbmc2HBDvVqsUjt6RKjyIqs
ya3dwUBUnz1dG1jtj3xgSEu9An32lrvTOf3SiLiHoVtGI8IDT30I73GWCB7KWprAwmOL26/81bna
k1b7rHgq25Ku/buEN9VsS8JkNr8mLMc5m4v3LNb6CqI3emCeml46UBDikW/4Dt484Y/x5VVp812C
BAeLrGvEcGOdunJnTtkOQPprmN9bB0uyewKxlNnma2kHShqOjEwyFCz5X50QJ4xg9JIRKBWfAlsa
3yDPTC9RMeOS4f+GtvVUhx0+8T54z6HGu32pNoT+GHGjQ535BNYY1YJrO4qH14RoWlnGCW284kr9
Z+80+8tAozO9t0n5+sUa9CAoljWAqcC+ulPGbv5iddHgzHLAbUs0ci3Kx3WcSL63qmg9MeqZkaUI
qeSuOkmzWcgpepzKklDQQWxpKrHE7MSFYWYFY54rsQV/uGXQd93wKODqRDcIO7nTNJvnMBc97xum
z7YepVie9zZ4O6AGgIv4V/X9HUFQAB/3uqrygv+iCf7qpSli/+rKWqe2A7FRmnh06yqcgRFUKE8Y
Jr0gMmkFZMUhvaNLyXvesVJM6pJGmY1ELGOCA7QhsdilTHsQrmmZzZBd5Us2WaJ/R/5aR3bO4ZP/
jR11OUHjucmI/Qr9BPLy9qyedQmVT8Y82nJZqqtCk09ULSBseCCA4D7lQ0cEcHkqw46MuabUeFf9
V+r/ZLLsqpRJ2C3pK5sZX8VWiS9nryP2EicrMK5eFC11Ggi9ElK/DDeTcJO+Vyqv+PMsAcazVDyc
Tuoi6GucLtkGFLB614rHYqOINpPYQSCcPf6zSu38WIUCXGJ+sGF/1BbBCfY5/GCdFMtFmv0R5Ajl
MowqVWhIQEFpA2Jk2xzLSAgxtmYugSguXO+qg5PIuJRZrr1nRWWgC97cQMno0ylwdNxrVy76pUE5
Asop49eyvHGFZp2SsMeJ3hxXA6DMwF3+73rMbeZcF7FMEOLzWqOLVaRaRopsYyiiRe5k9p93pA/2
PYS0YJQS0cR0YOPOAZ75XrqmbYpDiebvP2R2PxwGq7MuzAh+JStTHrEJSkC66f4Ne6ZRAe7yFqcK
hPd5hy7KyHf05PYMS1iTYTDTkU/nrUGu6xMtcW2RcMToyaUiKiVZKLHomcQrmSAcc9tp++VTvHy5
7+4C0Zs+Sk94z3jCdJIJag6EptZdIrt0GNz1DKQHhKibr7vpvK4DHPDSQ6yWHsXyitdl8R3hch97
Go+lMm5uFXmRFjQnj39yOEvS7D60O6OQhw8odWgnQNW171WtPd5WTIV398zvPnDGyxCZnBQUmBOC
LKfX2vjWE6F+ydkppC5mE3WLMg8R+NfnsWM1GcRqUpVjU45wpr0c/sykhausp8lprhoD2PG5qpOt
sSkhiwyxxHbsQmGyvxXmn2jbcOhMvNk497lB7hfEzJjMA2WvbBxRvkTDphcRj6z79DZad/1jMz76
6d1pfqUeQy/yo6cztcgasnJR4xE9VAjCOUpqlaFWNb0nFQOPCCvq1jwzI4ACos0QeEM2chaXGCQJ
ZhkIjU4BGrZ4e4/G/NBTdkkTb1aQJQRqxXpaGIMMFt7nzoBqrkopEUhncLtXIS2kmgorJ22md/vg
k645CQznFCd7dZZ/wAU2jn40yJPi4piUTyRO5qV1KEDYbs2HZ8W1kdp1B9H+8rH9TzJyeki2iGrO
7naI06ujpvbtFsNk1uL0rE+h+vqrJZ4RhfaYEW/2Gx/jl8rWnGVKRn6HLxwH7e5t0btQg9TVLubT
7TQ6Z8CSERDkmNdgG0D/7wsyPjajz/3mrra8zetTKCt+lDzsc7ALwJOYXu4MfHMr45KU0Ga2lF2F
jTDz6ZcnVbLXgCAEtLZh6AFfPep3zs0wixC36Pto4LyjxtR8yJfs+dpQVDJZbg45ChzPFZWy2TBs
2e9yzuSswGGKRZJo/A3qBBWFLpBd/dIKh5eYrF9jTX5diuU0j8K+YoHZ4xNmS3AuVMkq0qmKUL+k
anio3hxjKSXF7ST0R9968NYqOHb5+xQkKhEfGIgtj72ri6UtJtnJhr+qehButYoS7G/W6VD8XvpN
cffO57D5BsH2jG/54HE99kqXmPMEzghXWdYqBBpsH+0y/vWCh9xIdLk5VoTcFpltDo4Enm5Ep4vn
PwsIssTQ5Sq7EsG+waw6zsMddE5yj9Sneiqu0lD6wEJIwLU6MSDksWkUZZvf3IOK54bVOeFFsmCV
ERrfrSnRffDKIxxLPKCIPaKFSUN9C70H2c3PjJoUrsGzBLTm1fMCWWwG4vtT8MSB1IolzIkOCR78
Hiaa0jWUuRZ3C9XLl+XD7YRkyhDmZJKmT5TSTp2h5FggD+WHMhsq78z+Ld57DGiAbifaYSu8BPjZ
ENgfdx4EZuBWI0QRHhpSCWtFnxKWIbhbXIFISfuT1iqYQjgp88T+2GwUrhg8CmEb29mxzeZx612e
UttUlZpheqp5lkoj6G+m1aAKLOaoxZHODri9+ZyMdhQ41BKwqJtcvyx44RfZQctLmPLoKUhWtPbO
bX8ujzDmTP+8e8a/3JOJW3IYlfXPtKfGn65Vtoa1mjmB9krAUb1o/KF4Sb6cXJhokVt3sjqWsu+P
nm2pPRG+hG81dVfZ92rPDIlNQZggib4Apk998gpiYM7RT5tAN7zxaZz30A4MUnOILbUIq82NcYRA
O//pBUK6W9weAh/+Y0lPIr6Kz6cwBWYdCRmNbJhqibE0/zTpl+tiLydMP2UfCe6mAbype/nLYcnt
dJTe8zIsMXzPer2uU6+i+G4pIOfuh3PKW7TbPbOkc0W3dX67BU/XL9MoOFJ1NBdRKCZnH+fAgei4
IBMKPWrgigzPRLGiyS0vE6sIC+kREDcsMoGWAinDcGYYKX203fNp0z3CR0Wej/QhBrDUzfOPFz3n
XMJh+EyQ9F2eWIp17KYXnFcTW5cOCjzaHjfMVMJqMYHyyynWc6MzSBzRCr0YB+marMwqTyWFcs/R
IwWPkmZPdQVCIdCs6xlbd0cYc3H/BcW/griT1AAoCvbmeUjpM1CPOLHl/j3v267Voh7ED4W355vT
WE1ZAnYwjGkmaLZghl0G8qMIMrfCwjo0RfCERZpIkmGwZ+4EePAPRMsscfIBnP7y/cdjwFLpQGZV
yzqj3Lff9CiiLOQ9HCZxwXrjeKvdnu+l536I98RL8Z1ogYkZ4qsZnZueJsqjVNGpfcW03V+mn5lG
zOtqOwU4JMcLgALUoy8AGlvVRm5omXG3zlCNZmopsmLgBAFLBpFk2pGDTJQJ0NLNaSN5LH2cd4iz
QGFTgh4K1IJ+bWQzvDEygAL02UjbUqhg6JyMDvztWOehuJzWtRHljvthl7fdM6kDaZXrfLk12wg/
7AykiiOocnIimcJuqn0ygxzmZQuhy98DJkPfz+3T/8i+Rvt0QdxQgpslGcxR+XGZ9z1opHtViQLW
NqpW7L3xW91NVJyr141BccZ/XG+6sEFY+GQ1ymHcvqSQZ74ww/IPj+WQZBzNvBPQl8T1m1SxHRd8
wX0GyiV7uP0YhJ08gxqQ7ytU/Y7YV4xjzi1SMUayEPzYSVzzAUM8Cj2TIW1krr7AIu0+mzWsDOny
2i/oe3GGr0j83oZ2u/gzjwwR0bVFj90nEPrKlxqaucWUtrqGep69PDv06/AN5ymz5VGaxQDDRFuf
sLf5K89UA/xoKzcYzCWxuvlMbDCYSapAaHU3Q0cyzRmdVFQRBZ3opcxGiGy+1R9f94fd+ZsuKslU
QFklTFmftuOFX4EDqjfkBUdFMEzg6pdEBbgRXKXZQ9X3ZzpxP5zZ4yNyXJzFgbwda2QH89/lNne4
GD65ANRqIYZ/3jjoNXVmVpvual0SU5qMbS8n6naKSx72uw4iu6CKBD/5o0lsLBXUV7hpyWiFRpq+
G1YJArdePupivpaK8gE3uTu8gcJZUWHinQH2r5zxNxPYilQnLBFRnlqJM3N7913v9zXmD/ezCD9Z
66111/65p7A0hZKGei7I6l2h8Malf80vg1N8CbZXPwon11Eqr12VwtAADvtSSSMZYH0LHl7RZuY5
pqnvaUC0lKhy+RSyHrrqxQagv57QbdzLnHQ0wRsvPatM3r9XzDkHeAVar+t5i/9kVgIXaM0jUicm
H/0ndYFx9ghhr1T1bdP13G5/x0p7F/B/3XmQI1wGR+fi7rbQnzfNLB4MdH/zsjVAnJopU25za81t
Bn9hpu9HmadkSh8USX00npOUafKWcZENNUST/X0l6LNNkdMJwPwwjiSTwqISPrwynBZzXN1S3OIF
q/zjV2FfyIEvvpWUKGa2fC5X+JQg614EhZnoUtNKHDxGGMd7VL8bPoz1CxQtEd5HYpNo1KhlTorZ
FO7g61ZfpdWbIR2CzkThvWg3fXEWfBT+ztx0Z3soACZugU7ZGpapPIueM1fin//SrP5pbv4uOESy
gOJ65WOKV9teawGs5FYnagluLWSGEzLg5//5JgIvMhv2eGPk/Xri44J7qsZVmeNUHlVSkMTFYvTb
MT1Gwj4hWEWBM2mAItzNtxjyHvS5v2NJP4gzhxvNOeSkmDE+it73DO4BjV/3ZomG0XD8vjvuflra
1ma506UaXU0XTcpNiEC6CJuHdwIgotGvPbA9Z5qj5qAGt8zgMkqFcxOndHCa2qp5kTFHcryV4Hjb
WNwLCTjBckVtzPhecQNQG6u/z6nRl186UpZm8bSuLrSKxz8oraWwlZ4Yw0/VO7/2tqicpRcg9lO3
4DWQot/h729MrKN/j2PKojOrZ6rpHHBN2XBKU26xSuFMBdnldSxkfcdk4hfxk5kpSKMZrr0e4sPs
ZpQcALeNFW1rP70k8C91063kQPuB2NOBoG8z37jaJ6Qa29T4yqBcd7s+g+rUiA2V7pP4c4jkeZQl
CpE+oW+BO1PFfLb3BGCwajRz7W3sEBi3N0LB4o+tIJi51IeZQF5lxcILN1CkbsQjO3FGStGYg69t
luCJ6gkQ6JC+3WQr2QZLGbITpk8FSfGes9l0Y+/BYItik05Xn3OlK65u1W5IYOzWMw/bKtrsvzUt
aCYubcz5QtXO2/phN4ck8APhSHAD59H+Q34Ik3zS7fzvT+1fMbqeomU1ivvm8bh5SSadL1fK/B0V
F9JD6i4fyyhXXSjvh4DI/+UOornhRWNZL9k2DARyre1YNNgo461DSQJROTcpshQuaRnF2cz9T292
XgW2PEvj0lPHn4rIoZa/1NslsN1ct4J4EeQDSlBBJ2EHGzTonFWUhRG1PnC2TFYqfP+966zFLJDw
a25sDmReZIXPSXV+1ZxoF+VvmvzEf7mq1bVLMWvVzkPwQWVdsn3Okp7uMGLlbI/5cC7lUgYN7HeB
rZaA/8hOOKUNplM/VTzL7sQCbTa8eDDFbOMCFYnP6yCsMBtQqxvFosS/DgXSkgwUjsQ9FtCETU8z
8CVd0j0C0DkEajjzrwsk4N94l4vRnnKVZgIu1OId7vmahRLKnyaGH6Q8KBGpUDbpO8k2JryLSUz1
eV7qncWahAoR+e07Uo4MyAJtiOvQoWIAWVqfdYHjqO/WhbsSUi1NXWowb0+QqXwy0GfzsW5Ill2i
JsGhqE7I+YnUn/AJrt2qbOp4c9VgN6kgXINgWLsWla0OCjy7K/vl2WA5aTkLIMYNjht4p1EwBWiI
NzZf14+gZItKRiHzGn09s2YALSZ30RJPWWmsqBJdd2nUsGwUHC2NntLiq6HiOfBZ4Qb8yRgYezM0
DbMYLPP2ZncY0VCbDyD6na9ludfAqLWMZS38NINEvH6QM9K84RkPAb8MutEyU/A4UUmC+GmHr+6B
xoMnUslRFL+JmC+JbRKlsSoC3bfyilAFhGevjgfVy5SnXOCt2ufRlwKWRm/3LIt1kWW7Q85/fape
C/m5T54ORSwW3Sd9wrf0DsEDZ336U5M7LrJz3Xf7g15FB+jF42LJQjaWah4bLUE9DZXmeY8NT2H9
7BVoqYx7rX0BPfajUzmc47FvEb+ZiMVS+9l2vHV3aiADqOaG9TPvOnSNLn8KAt1xBkiVTkPBwv0K
ir4ZMQGzAA+TkjZ4wPHukOrASPpp6YqeuyHORG9H+tAMq6lwYheLeMnvs5sgGqSpX68urJAs/1qB
MJ25RtNLENrwpKkqsCh/2eknWehp2Ia8O3NrpgTi5LDmarV0XS95LpUQItPrvIBGFSKuGXNAcUws
Nn9iVE+3RORiMs2ikninRpatg1b0PPCH/+XvGd1yNVL5eAvTs+Q9cYiV1xIZYzS9fs/ceql0DFj8
CFhp9n/wygOZVfLtHAbU7hsSRZKwadXNsp58t0mN/han0ew64+zAknT/nZVLgR+KEicTuXo2VEmw
5F38ip6ZJIOS7ozC1SdlGFJ3ZozIRF2c473ZakY4fTJel/kWYbehcyhRQRB8tTTAVDKEZ1SeYK24
0wBlM1X+b0K1UcfBdkcF7DXEOR4wWJGTboIauUPxxJMaP/YfDfhLjO63Owo4t8qbiaKHWKLU0kec
FhSuM2VVGW2xmLPSz/97CTxYnLMihdnjsAKhuCfNxsT64noNa3ZpE7aclp6dEHl40QC8ymQDdLLS
16H+NPKc3wev5GBaK/k0SAigt/O3WsMX/jWHfnaduDOAJevVqs+5s84oBOlmNhTLbqz8onfSlJZh
RrzOEYwI9Vy58KJ31xtShcCzT2dErMg323+BlKUmOO3/hEHbMoBzSz3S69eJUIGxLgao29L91b5a
/R9SCkBVZNdLDBI5utsXkuYnI0uBf+YZee+yT9KwTUqgGi41RtwDfNxp6Ixch+zaDCv+Mp+bdMZG
M+ESwXKB7jWyv3klxMg0rRsVDgDPSCz5LqwkT/OgY1lkvDusDle0d3PBynZt41qMPHhjHg3HErXb
gjx73X6uLGoSYS5ath3tfxG/BY/JvqQi7MVagwiVNwa+7vZ7TgP126V9CNGbcaG9ijahDXj8pkmA
Nqx1mimxEoCy5Z4aUh5MUer/02eCA5Yuo/22e8es+AbLzINzG9IwbcSCWNIQKbemz2CiGQXbenGb
UBZ7Ggql+crLvpy6SewdDnR/Pw9zY+2Y8SpYx7+4/lk8bFaVriv5pbcmlJ9gAwdpjip6a+Ptwy3x
wHG9Z+VMEE0eC+uHfHFHltjDbxbD/ohn6gr8gwnMSp6Z1v2ywNcwBOD8AEOm4HLiFQp/oEtT1JOu
kUjPnyFwUqUS3dTj8kJxTbQqLSgOMT0lxaxVwjBWWVVrX7RVfHC0RtN0BHCFoVxDUQ02MesIvUnk
YLeACewUps0XGtxupYBX2EqBj53/OAwGwFdX2IiF4RF6sHzLpfFTW5bLEUMR5nJZoD1SMhYOPIyR
Hqk/VmZzednDs+TQPD2hKsa44jtP8IpRnRiQsZeuxm6T0iRpIs1RrpOc3tAzc9HX7oBT/6ezVv4u
dTijkVCRbDQ6xGAY20aSxFrpPiTJTlbVhOLaX3PH1/sbLkRNXICq54iztu9wCpR2yZw6woUypWzX
BjWHgpULLuFviqGUsWdTh239h8/41qm5aQLAc0sXOIx6VnyxmrWmGX4jij9ya3gMexThR8NaosNH
y82R1YqXt4SkXpkUeaVFN26pp8ioiiDjxwn1i950huSOnQln1cy9OG6BhbLp6bvxnG6Q5JZwDJxO
iUNwa3gdUc/BtkzuMg+PbGxIDog1biAunZoTietOzzEK25DGhchPjYBsSQaIvbA0iKW4kJCrRGTR
3/b8HJcalPHlEAFchAULTtTLNANTbqVPPPc5oC+qXqvS8Gpir8DWBug7u6OVeBb9bvn9oxpGgFiW
lYM2zBiRmby8LS0hBkay+1gDhA+Z8WCuVRgYWoZBOuksaEQdgmVkO+oiWOcVGS84R6vLn+CgFMjA
1EvkDq3CSEhW/DPqVnNhmA4u+9bjcTon1ia/BFkUjg96laC/b6aTqPeWeNCOQZ3Ury0JaLPkSvhM
hZwxAwTvNAsFD9Q2FTbylCELp4wNzvlCNJMp9Y5HlCpMld0P5Slo9dsKfAKMc3UFsCn31SFOE+V1
rrdGtBcwXp7bzOVKe6taE8rlQb9C7m//ImQONff9kAjblWwm06dLfCn6jP5BUNMBNzRrOmEj8tLi
z+uqYsu2j4Thr4qB06qufnYhvWF5FYSn8j8+vVrSOm7skrkkyTR4wWehqklAT5Hutns9fSJUvBr9
FOBuwD8ir1K3uWMF2/zzR3tIISleUj1ek2bMfmvN9kq6FsXEboUttdezI8TGJZuZ6mvTcHSO18Na
ze33PvZFkf92Z8P86GLSiujEYWF3Iv30hobCgrWqrixpVcgR7Eb4EbIwmrZir4a8oBighzyh9uAS
v8tvrTtdnnsixa2rB05EyZGFpbBbqmFH3OzOX6UAozUVDpxGdp17b0aQ1PSRtmoP/l/U5KkA0gyi
KqFy+7+sqTlQqMLOsdd44D6pQEj3T6+S7E7DVj+bY4nds9p1KnxD6RjGI0xfyyV5kcDnxL8poMQc
fHL6pQ01AGUMyxKsl+g1QUzhpwegkCZyePadxNdvvXKr2Y7j4tALT4TO5k/gPBBMZId3BBl29vMU
4Mcp9rvlSb855/rpDHZ3sOtUpgaNbhGeRAg4mfsctm816byZOOrDzVLp76Xq9vWCNO+kK3hBbd75
ogQhXz5NPuC0cgSQKrRplrLo9QBAA+nwN1xCIDq814ybIQaEYl1RK5ChToZHjQ8FXMmBBd41aLTm
wJNzccLp6qrYU6U0BiWbxr3VOx1BIt4iHGuAJg+YxCCZTYqJUiKjJSM2sEdxA9bFKSdR1f8K3aYd
Aj5jqoEGgyKTEkmRF8hT1Oo5z36/JmJhEB2qgFVRYlkG9EKc1AU7wnO1thF7Q7d/19lT2xuKPC5M
mWRlceRbLsthIGUlSI0dOz5xVHaCa/0ApVcRTdFuhM+WbGz001llLrRLnnTKNrZB23cJRK3jtbRm
yxXzfgDgfwcJves+jKMysYmEdfQjNdNmnWLzFFs7PpxM9TxiIX5nC4uwrDHVZ+YBajN9GyeXNkK/
K6KXtkl71vkTUQMRW1Fp3RNW1jhTUzJVfuJUbPXISt/8IyWAJzmf3eZnrUilhicHDlyoWfqxSb8X
juNHLVZGkA1PeKJ+DJTnGjYAgaoX5vDPaYctMRYgwtH9gWJRPMtbukpH4fnGDXfvii+wuE3B6+7w
b1lS60GuE93W0KwVUeS52pEWTOPjZ6dpKQKJj21eOtEkhSaVPRw9Nt/VbhavdeU4oEBtGJgi/FvT
PwEdbM1eyEg2hmF12yZxGxNg1UNHi77xFpRU1kryU3sA9xW6MvY0IoUYVfvisVEx7RhOEZ7qP6Yp
IRq9/tyscLhj8tcOIDE8SlIittL7WV0vilpjko5ZXYo0QN7I7PqF1An3CA2S4529uLQCtZkb298S
hr513fBsbwopVUOA9z0BWP0A88pQ21PkwuROpMFhujoSgQqj3ephGhUGCUDqJW67XdHxIVTDMTCA
TvJZx1rR+ETF83trp+HgLmT1OOZUmP/AObXrlnR/1YuQfdpjEceFypQp+irlcgMYJpelfdmzVLGq
Uir5ZvW+9zFHe1Q/e4IErCHWqmGXhis8lVqXT3co8QMaYzD8a7deAGxX8fAgiTgfrelDLyU2tLcP
eIBotFUf3A05sWjpQt8sTsf7+qfmknS5D5gg7tL9GMSLe5a1NhgYLimp/mVCfpRAQw0xuIROYOZM
fNARrvHC0FrEe1OYARq3kcScipB9wtXAe9y8PBejoWwKqR19vb7fYlGOeB6jGT6jBfvtgMEq+sTj
Glf5ljX7CjDnok70UlYAgkD9RX5lFVmq3LGk0AM1dZ4KIsluvT4V2ynqKjhc3vd7WMN91Yn03Xbo
Jmj39o7ktDZEl6TTKV/F1SP1ncIMANKHGDhJzvIYTeVoG/S/Hd42lWKgTRNLe/QDVlYdPAktVaKA
B+6gc7gYN+9DFP5KzZdMwimqEQjY5LK9P+h0y5DgcrF/PpnEKnG+jhGnUwdYQHju+JVKCLuBg8sH
ysehazoiZ8DwC7rM+RZ1EGn+iTu1A1h90G6B88ltHqoy6oPTHayjnwPHVd11cFLc3Q/x4gfllkjc
BKVLXEKu+mOkMB8ptAY/AZSTJItRl8m/dljUJg/jLkMY8XAooYxisyarTP2iFIdzJuqkLZN4WV2x
poJzY0uzb6lVNqKCLJ7nxUl3BVPRdRXBs2uTYz6rTR6Gh+ChCcNVfT0JMDEkq+KKWOROWt3rYXig
phh3JGqbRGo4c9KnWIK4wClhEKt9PJOPAIIv0DPAVa7IXna6kk/5MgYAfkk8fTJNdwR95Dx2HM4C
ecvqWxdmg7C/B9V6pgigI6o6Kcf69ClWtq56pJj2/s5LEvSnFRaoYLDfjuz4GoWBURXJsaetMxzw
QBnrbD9wa4JUxrV4wwEpoHRSuPKSkKH/t/2151k6FNND6gjtDSZDxwsQ6bL3XFECk6sHl63bhZWE
Yw1dSvXvZFwWyHNZatI4NXSiSz9OGf7YDiOYvDqSnd3EOaNq/s9w34wsEDtT7nKjYG1Onruph/YN
/1sjkEpbwLh5PFPrSau6UxWx/5MSp1YO3zNduvhFtg0ZKTgGHxjE4RaM5KOdfNlcBaQO9JU6isqK
shBev1xdzyt+qoNre2a7EtMXS/RJcQBlcBk8hDnrhJ1DL3wRqCdGJdPhreEwmlKd5gktfv68gJ37
H/wGkjIOJt+EDnXGwo0DJ4VO4QMFUTgVx5mn8vigY/CWyhzdzPQyepL/Df7sLJWQC9CZ2CSiJsfF
9IsqVzDYozvLLnSFjAaxTHqOu7ivdsoDCc6GP/SPukCo48DB69O6RvjvwqJBcHUwIaiZ9oS9ilGy
aZ2meRsTJ942ifoGzEta82Q63mQ/fGf5voiWMiMKvBtjgtN/aR6Cfiub1YqcDPcATdzYLItpWqX1
Y9ALhjYM5bUg7Eo4kSqr1gOKCT1ucYbFVZrAnyi5IFNUGnd1sNTFrlnAvcMZWXvBcLNi6ZpLkmpd
x055xBnKcYjkr1D9FvoT5vPy3UTmmqwSbIIgOEpDAGU+YrTOzDhEMfwAhNoPgfvMmf1MP2t+M1+1
cyQm2+BIbjjf6/d/R728PSDUdQP6Gk5V8y+SGD/jFW3PNhum00Z7brxQSrTiWQwrXq3vDhRJt5Gg
kj4YfKdwnOAC+XZcP1zqlibiPr4LvSd/ZaCmS1wjvxPNFMgmHqO2jmuPZhZmRD45OTNAhGse56Z5
ztEWeg8kw7MUOhwh4qrKniPkaWQLPXIR0HcIq6jIoIKOKDWl3hlIJ7ySxz55N1bKlvRPKfiVz0D4
YAmo+9we5B3iThummM4aPnB3kO9C5qvfPf3nRAnw+1jdPXykhtPRCxoQ1CnVj+EfldOSQhjjdblp
+XKoSVuQLK1kOtqmPT2OfMKguewT/Sr3VBvBqjXYdomAgyb+eAWeABdSTJo1HUnTKBQkPGk1b0qt
r0phif2uUTA8mUtJDvmdN0SG1fhDtYbHpv+cYKTDYHAqVdC30fII750XxMMl6NhdSH+FAaNuPpXB
KRbyQ3Jiy7dMmBcDVkkD05WRKzb8PAJOJwXF4JI09+ybHHIRBJA1RjTPIjhApRXBgzmrFr/HiO7k
RvVkZRpOv5NBoVNqXn4z/EHfUJQueuBHT2dllJ2xiPrHnKn7b80wzqbrnYLQqZLVppN7pgA4Nz8n
oN+/AhrfWzzADwSraxIYcpWgSHR16MQvZGQdM6NOdquLPl1rkqbjG1uisG82/r8M1a8WMSzcZWaO
E1mrTGLS+i274OF6WiU5Q3Io1S3HI6rSF6mmGa0yFhQoZd7Y/6hx6H1TdJKjxZgI2k0pZxtLdZuR
uk2RzbClpr00NIzHA5bdO9eIlwRLW2nNqEMu4j7sQeUooBduD2Hu8eeCEix+8mQ20BitISOIc/O5
8VTja+w5zQPqHs0TomyQI5/2qYuHeRyQOzkNPEE4vAECFjj6ij9w8zu+gZzWMiyyhEG7U+q3oTvc
jpmIUSNkWYnDEkq14jsCAEBorMNInoVla61wUpY+Z1moOz3pl8h5CUNiHag6LFB8/dfwTy7S+PE+
ls+VKVDjp2PEFjebY1ngHjmzFAvARQQppDU515k1We8h5DNmHvW4UhTacPpZv5oybj1J3Pwf71Gf
85iyQ7PFtox/Qr2R3Bmhlf6Su4E+Lzu7jE+SkKS4QESVuMZy1H8h5vYVw/8kLbA31Ic1dtBoXHpw
C7yJ1CP7tKO2gb/qXLUyZoxgsmWhVfoURPyRFpvpGrqYbiASeZloOfPRMwop8TWvijJufO5I7BSH
3IZJsGW+6u9Kf/E7degDcnjXplM/7PpoUiaZ9ZtUcwP4pL4L71T966HsnUPM+P22OICm0Vo9vfvf
5T/mWNXLFQ7eYHi2VVvV77MzTgssbDXi9+f0swo/zsljWAT2rnEb00DWdr7KNg01UPLTUHnmcNrv
LmBAKqPexR2deYNeQMMadJZodnxjsU0HZlc81m04WofZyvGEa0QSiRi1K9aiDTo6drAHxq2uKhfo
qQXoAJZHZaTr9wfV0gitX4Ufbd0y91bzXddZnk9OcOUEFH52B5R1iNhYpBw99sDl7FGoAhtyyL0t
ZWPMoD3aD1kvXf8hKCMnYAc2bzlD2tMOuhXsTtHo3XRymgJFw0tqufKKS7p4L/Y2+YCWla5WWV0c
vBGbz2NDi8pjCZ5LvwlioVR1+HJw3pHu0Unxp5MA0Y+gD96Q2zqEYrIOLAOpIYR3cAPy8Abeeo9b
tBl5gh8iM69Im95k5sQlgP73JjUhqGGgkfbAfXdE+GaCVuwe+SjPizoGVUxUdu6UDkYzxyT07wM3
iL3tq+Tx2GSDTIDleM1w7ZpmKI9Srgci8bekNSHs2xzCIhE2c3EvoCGjS5PAtC5ZBEQf67yCTZl6
NvB2fXRoODpMWYBAax0bsyy/8dTrbiMgrURESFNmuPkczatl5TAlelWb1CES/t2xwJGvrJimdh3F
rcSECINqnrFlGpEmzy6j98MsQwxLav3alvPxiOAhOaKVl93tHfngRqqExOtzyeTgHOxD6Eiz9RMg
fIoO+1KntIu8LkbirxZ1LKA1rgmJ0rfhSeCv/484TCz07TgFAHIu0whQO/de7YDhU7gMs17e455R
Mppy0nwH7rf0u2+U3nn1QKm9K9X40VrfH6B6QxkZrJhnVc1GR71bhp3F45mrjee+tWDLJi/CXLtn
XCxGj7vEYKZ3/8UQTz/Svc2f+/IPwo3SEUKp4PX4IBLgsVxrjqG/58p3ZeWmL1KRIe4LIJ9zLxmJ
GSbIMPTx/f+nWqacFqhRpMC/dvqdlFFWKpVqFYPpcCmCevHE5lXU24p0XN8Gc/qRr6Bpj4NBvdTz
+pxoYa1CnW+xvsUSUzZ26Eq0YlLtH6HEuIeBgxjB9S+oMrJ5+mh04Dl4CgpvS4jxmpTPJUSZXais
LfgjuMw5mRICFh+tkrl+tdv9622srMglZNTvR+dfZ/ReVjMZPbuEZbeXF3ir+lMCzOlxpp0IXPUI
gVa0WukwhIs7Jb3YtjkI4ZNJPxl2TExzIGEMHtB1si9Bmk1trXXkaI8uf+bWjynXYZfNd64I07F5
rrqDsR62VdfpdJjtEAhULiDJeFIp3M3590LUe2eX63fWYsyISNA5fER3+VSvqqLz5OEAQU53KSWi
I4cubT+q8pDCL32UYZk6AvwK40Jcf60/YKnbRmDTpOe4eh93t3d35M2CO7xnuTj8EMIIXEx2ZNHs
o4t0i3D32Ip2oG+SPy4KyIQWPiwGalb7UaBthNxdmyR3F0ee9JUtYU71xM1jL6uaALHW1FRyIfCT
Ki+lNbkQJYKz3jdm/lHeTwRTE5Vl+JWTMJnrx6K3syXUZ46AV5e2dMVaqx300kX5VdFyB4vrpYIs
BRsDx6/24x0YXhsb37b87Q01ovzlbfpQpJ4q34QlE9WiVdPG0iI5AodKxlyepwWukEjg3b/SFu85
8aE46sMT8kg4c1bvHAP1JjF5mI7m23vbT7+6RLF7o80OaN4dN2joKtVNDwnxxwZfW4cEaEcPvUNd
6L0dol1YGp45uf+mMTO2jUlAUjkHrnB+rAP16js5R7uRy68osk/uW8BniGDBIugxM9PoZ8ya/TN6
It4EW4+fpxOensA20sxW6Gp2ckzQwFCfgAhFiC7Iv2BmqJ5qosb70ygDtonj4ciY2y/WIosAWanD
jglUoh05oRAzavmVtTT9DQjxn8SC1RTom94j0a9YMSm+nAJGVLZYyS/s9Us58ycXuCA0Rvpn+j8k
pJdmm6pymQiXm7ievrX1/0e//0rpTOfTHIXKCah5ADibFTqbseIDEblsZ1EKNa2VfjzQM038S+tu
3p2PbG0ccr4CsRzxwKtvPEi/Ub6DF/NOJmEhbSdMnqhuVO0CXoDjwI7icO91bl9bX9zF1MLgLN5S
wLbK5fCTJ0vHvzvVtLNZ3Jka4Yt4zd2S0toAvk4gEkbALTeU6+uAI0q+PIfeZQl4KMwzQAB/o5i7
QS3CSy4IJqteXS5c5zu3TGgYR4CebKzmeQ6L1oXTQ5ZfGysIO0bbjdb7V1SXWzvR1NNeUGgnSKDH
eyM3tIoqKPMOkRNt4C982qpc9VVxfgoQ4Wqlvq37EPoCgTZ0FpsVOTQ2R4pqqB/c05IVLNSLCBih
oDatDk426Pl4d1OtdO0iWtCc5tmDvVdQeUae9J1yu/uk8tyRLTX86EXJnky9LosqduJ+qmryXIwY
DnEaEUfx5BE5l4uYHaM4qoGxME1IUBwRAJZbVm0LuNKkF5W0U76Q/8Ny0vEIYaG98ppMsKCrA10j
yCK8c0Ob5SqVNOJNq+Lk4xy5QygV+qn4Ios8Wor4r/PiREzb9tVpJqMKyUhr48PCJ0HbMesYt1P8
/ilWkQ+JEdKsN9BKXRLXMWfJbsldpmuwFxXuVKu51ee7wiTsfj2c8AKy4IVRkek1TtmuTwWx26L/
jYWeU7WI65Z0jsLCJ46/fzINCqXjhbkKs/swFCuyg5haesD3jlKZyph/xvtrOvs//oT1uYSaSECV
2q9ynh959MTI5EMszntdB3ItcsqBDukd9KRXHI2mv+v//bt9lZdfN5Yz7ii4Lm01qtIWk1qtedmV
ziZd9tATAs1UrHqZAMLfHBoFB9wRtZ+g/Z4maJn9A6JuFuACiA1OOtuuHPVNLFY7l1dw4JS0La7r
zQkYew3GSSsqNqjMO7HrC80PBYS4stXr7FV1+WC86wpgDWBl7cOzdRvOczFTWJPMi4koM1dewHW/
7QaCNegOulSU0xVAq9Ev43lHTXIIM+rbtJ8Or9dO1U2yV0mMtse/oB+UrHfH9TZ+d5caboHc/4dO
65hdttjLN3ZffARvdGXFyyc/JAhoxLreYO1SpG3MJzYd8FuttYwJgNSEH+gik33no+baO1a4seLV
fM5wGfY6PnS9zLWRVG6tu8rlqqsxPBRubcwUs0E8R7VSxujJyh9kUrcsZANf7txurz/QCOvbE/It
RZMdAvdBiMbOZeSKpMxxOMQpGghMRYmCJusy+LG6gwNq3YJzGgmnmHnKVVPdj3BTS6kjsv+HbgYI
Y5dFAQu4P95p5iDILOjz5lhpEiEN1ljErC6trPdqafswHnavsTcaO06jBqoMXU4VVZ/MkxCDVJau
+yiEUJt/4JFP7W5zlQq3SvpyprsHikAwfhYYPu1BUZWiio6/ictYofxrDwts9qfiE2aFs5vpj/Wq
O7vBr7bi67aBsTSLARR0jU9B2c9WhIXAJTKh/UaMAUOF7RG/ddD33AS0vD57M+hu6rksZ7R5d7Ai
BDef4JD4/K9IxSWcbpEveWhFuNJFhWP3hvGwWa5h3Bzwx61oQ8CwRMAUbW8/TCFcz54XWHOFevQL
BSmQxjEUFuU4urNpYU0lhXnr+YNwuEhd2u7t8DHCe90VXHai16f7Uu/cbhqaGqbr9+Bdk7o9y/0x
YclgSoQM1ZVFqBKqVKJwbdzlfaTUnMwb0WOR5Qkuof00iA/zyeLi7bJh96/3Kht1sWlvqA8sCMm8
lQpdKt3UjTGLcZCzrW5SjAiCH9XAQYBVQ7bRGnwttka7bwdAkw/YYM7joVc7hLS0rmpATnW2AfHV
us8pZw9+AlcC5QkRWFJ4kQyTUFusjZnyivx85zPug/xf1fX3VoeXdZniB36zW3zLFj5bLO5j98a2
FxFUzzyOUK0tBSNZmPdz8a2qmimLlD8YP1JjKPTncq4vrtQ1rCsTLWa6sAXXmEQBoQUzLHqY/Zsx
qs07iild2roHTtzooHW7lzLtOR01+IRZ0l2wf3tNL9aGUQEve8hJSzCfxB9kurH6+3sIp+OmRSOO
F6/oM9+4B6pMhyKPz1YuzBg4ax5mfrnSl1l2DeINuoUETzx3/l8fSZngaRwuVGFpjr45tOr4nUCZ
XTyimOar8tvQAo+E7SI9XCARD4VLkKbaA4ePzCyV5YvMuWhqkj9yzdTbZWHMvNsSxiv2oYHfByTp
CnDWYJuRdeDonWHjnzRyGV8SJ6O70Mp107hoaw2rXzQo7vIFCrl2q5KbxeX8N2Vw4UXZRKQ2ehzJ
H9JoU81kBAEs6lIeNT96HwOkw2aBX4wb4UFXebW5LNKBdoo8TyPtCIUVtcO2I7uQ9vdu920KlO3s
luIVactbMb1+mSiSVMaXMB0rYQtmXzNnKh7C+uzpJCfJ7SqNzktxJC8fr+1UY/TOwZIxMv/gh4VV
/aKx8LlltMCskK2Dz0CkLb92pqua1CIKwIL4zL/cNJk19gxXCqlx7Ez1yY0PXV3uxhCxswQx/VGk
bNDmQKmxf98GZmqEcMvIQRJ9cLNmilu6q2xh1zvoJpnCurEi5W6OmscMkbHd+nJu29jURnNqs5z5
/9t8rplEXtCSP7/GN8VKSiyfFylelrzHu5DDERhMXYPOdOboWt2TJ9SFEFCthU9toaehlDqQ7Iu5
eUOgMSoCrEwfInoH3d3krzg7ZQKw4obTqlfmCWNgeVkEASXYwfgf+Av5+HaQ6HOzYJwq7A2VTQKo
kiZ6/EADZjo1j8BrxhVsfZPWEbT5F7CgxPw+IHoyAhzxU5t5ncPzVE03L7oifo0l47y+mnTzz2vF
O2PndrOtPBz+Kv+z1bBD+CfV2m0WLJC6Chhu5lZ5I5GxXAv+YZdVcFc6u0JUYaBVl9yGJf7+1+yH
2Lx1b/gKhBGSEblXxUmDwjD2VrVlFYNMlpy90ku1epY2MwGXk4pb4R7IRbwvn8QBnUZieVzz8KGN
ma6MIjuCoy86LKeHUjpLh9qlhGVb8gQSmF1+Di+iYMLzVx7+YheFmavuXYUjSlr94Lng1fYI//qV
PO371nm3u0innnQnEeifK28bSzr2G1vYsgM/x++HcrPWq8WnnUcwDBj8QtPLxglgl7bEXxbQJhvl
dI71baUQ5RLPZyPba/LXapV2AGuUby82btUJJ79Wfld9CulEhN+HhaOxA2GQ/OHpUM0GFSz/D86p
9Bsqv0+aDDgn57zQz5P26bdFbWEtByG5D2/rxeQ7/N6htoN0NO/iyNBUZG5/k+HE5n4e0dkn6UHR
iK+GsHwYY2uItHO7OIDW0WbhkTbG8R1vhvilwHN2CSZHJRAJfgwWNGEc/Tnf7tksHbNADl8PT/V8
q0Xs/EbA0dwEv29dP1qXErjFsgRU0ZGzdgOllhcOTO4ez3S69N9qnNLl5WSklLXcDMj83mDDXwQS
YGXEJNlu/JBC+aKMQtvwVGjqf0zg9uT9sqMN84WaGGfoXrZLblOFZAjBOajvJhqABFGEZBbzQTKD
2Hb2GGv8k4zIP7TPbfiUExli5fK0TpmIRSObAHxrPuFX7EDR/EXaxnmzRH8BYQ9zn1g69DW1q/1x
edxJjJcTQrzgiyhSnNPrcEYrL0Je639ijUDrDDJSSf2nyFIQqGzJZ55DZPU3NiCJlBhbNG/IZ8B4
vmhr1a3S2kiKWdOANudWkiQ8bQqIpCI7dqBqVg9qdGGjQi/xtjMX7qcFmJblAzyHEbbs2VZVNuxM
Ifu8u4MH/2cQhrSc8OzWvSqgm00EWL+NbBMHruhaMOjRZgXXcjq3gS600jOogFKI3Pr3B3/0jECf
MbRErtX9LWf3hJH/HehYqZBVrledN5bXpTL6Mv04ZsadAtRC4IxM0LY5YFnO1eyFliLm5xrijjqQ
F1Ln/B6MMZWP4GkTDPibKuC88GW0TNwWslenbFsqNoTnWva5gx7ScU//NcnXoxcwkmy5JAVLPLeK
XVW4h2y+WN6fZY8FU3ciFz7W6PrJHHnu9qpOGeQnhDf2MHh3IhG6fnCCvy2tTMmWUAiunrNYj1bB
SVNfA4YK5aJ2soMBms3qBiZPNG2uAG8kzhs9VjMK1nIbrlH+UWBjOyhoECSpamziBB5OYCj7M682
EDvhDBR09rofc5+3PMOprME1YM+DYUJNdRATP3sdxwXg5IVjbxn6a31iF1XtC/F+YDLAou93APd3
q53Hn7QvMdgxz2cXtzIxO4fViD0+ZxtvwydlWAcf3lNQuYtaU8BMDCdK4LvATGdEIr/XaVLY+O+a
jVq0+92+jWud7jWBP3DCgUbvKN0oGk96PI9BJ8w6dAZT7wCriPH9/nZ+XDPSm/NGX4mg22nNNRPk
OrlQ+8PNElZtUk1icJGMrwCllF6IBKhTnL4brsmJaL42DmQWVKi9FAlS8uOcudjcmqfdz77FC7fb
E5mjQ52PgKCm8AHF0PEBbi1hytArUerkhD1ephrCOr2KTX1nTtGpGuhOkkeVXx+xqiQfp75l168a
p3kp4Q+BMsuy61oTGTokiCeykEsy6FaVReEiulKE+8iUEnzbcCJgUn1R9AMo/7DenBscamDTOzgD
PBZLNzkiU29FpAKaEDeHZTC49B9dro6Oa/IvK8kmHqs2VgmqloaUX3lN1ylChxesMMOvE+wWfS/W
QH7Hj0rESoSBLoTu7SMNuf/+f41WlPQ2DRqWNVauu37nXGlIRa9vt9n8o0yung+Tn8qE7n5KqO9k
eVFqih+9cjB2FrP7+uCmaGSeBCIOOjl2FYBQuugVxtyi0Bmikq8yZ76l2HumTjUCE0Odr1bKlxDG
3utuY+nZwdMdegoCz7+ljq5VLda6j4jr/0AGIx0gtBnj2Uzuy7wSHdqFcbTD8v8Bi5M5c7Z+3GDK
3LLS5SXddpqmgrpL4EXbFW87nLf9cjYaZRfGX7zqyBnMO94tSurRiaJzfH2bj+1qPbces6kyNRt0
5k0OBFCuWjTjb7E2rz2r75nqRDtqnyzt9fdQsJjHY3BiyplScT2hhzConTekGy6RXXyFvnA8t80H
CyTZ4wU5mRNsV9K01RpdJSKYKIDm8dH1R7gkKjfx9/chliewCRclRpR/UGHvdGRSMPmy3oBYlg4N
ZLcEQIxt3cOlQgtN981HibuO2PiXxpPVOXPLkKNSgrEi1Xz5NK8gSgldLEX9WOcydz4ZWOUkRx1Q
/zH9td6pbCmqInGSPKGJObQqAr/g5kOnWjse5E5APjfEzjz5+WVKONGawzwUq0sf0mNyTyFY+rPX
sjrYCVLQ7e23vOMBNHekmfY/UVsDgajEixZrrGG0IjHbvv9w3AYeptDmfG4z9cC+RKY57itsEG9a
FCLxPNU2fYCIPT9LLQyfbQdiTmQmANICGot/J44i7rYTHEX0k4Y1fKWX9mqNBvzRxb8ox2t4enY2
iiLu9lb4B1rAEpeUbbdPRkE3wzQbEOn/cQLyLhdCspHy3ey246tDsOWA3dLuf2MfYhFDptrHMcek
E5K/7xWEXRNoxzLM337Iqo7vIj+07FGqXeTsWWruLjDohxHRYMI1QwQ2riZWNVpObrdTzPfHhNqQ
u5zCKjsDvekYPKf5r7eb+f6wurjImfrnN7s0q4KfHuB4SatPIGWLVQCOeH5b/GK7A4poqx2Lsc/j
GgwCyuAmP/g/en2kZIxzAJPTYxAVHBROgejCk2lMfwlEhjh1KZbjsmNML60rDzWyER1RsWbtYbjQ
vOublN2AtGRpXgkfaT/PSI3Bta/oeVg+uqAVrTU5NlfuFZScmFKzZZQJuloYtvm29/lK86MXsldp
fcb1ibCT7n8chhbfpttjJKiHykHnEX2SLigAL3n6G3fFNoTdNTQ5ynMOY6ESG5yoGf1pN8mG6Ssu
9ZvkbUnuOX8NTnUuy5+NyNC5ujbe/LD6jbmmw+TNhZ0pE1X6SXK55oslwOV7zNnZinHioRIADrZc
CvbKomDEq1K4Cd4fnYuSgvwEUA4r+eCooSSOARJIxtQ9krhzbLEghHCpaeBVpw++JCYV6vzTCX2I
L1iqCrCe/EPjUAl62osyGRPDdHmU154ackAGkrjrSa5Lud0ZDit400N6tlemTVaTW5f8LYI2pnFe
lOixoCOzZl9XiaWQ1QGmyjaFqXt2Lp32ohvTmSSuf0Z9teHd49oKzTkYS3vD2Bp8FJGphBjQR7qD
z+FGmgXEVON3XM5k8n1P3o60wvTQyQPEu/cToGh/e1vumVE+x27aP35oV6DM+lHn26Jmx9F0OQs2
GLJgDtO1Q4uhzCfSoSe2UuQGt0ZT5Djn6G6DdIAIwX1odAaAUrZsXHpmjyj7xubopZgfR1zntvGX
K82ne/yva+1wpcYkGow7AK4cEo6Doot2d9FBD0fojh77RFsRxjFFeVzoOcjImFUJ4CdQ5G4vUWGx
p2AT2UDmqnquiEKASWIaLqOiDBzDMyxe09ZpRl6caq93vIQ7axlRYu+KsROgH5rvhvsnK6qhq4Tx
RWZggme3FxE8utky/kvEolDP+dKRQCFkJ2sRtSipEE5Tcuw8ipA2q90zywGUAC2rZ6t5YzG76BgY
Lhw2nFxdJAKgfoPeLGOrj+K6Cdw0OrceDCsNpLN4K+KH+EZ0uGAwvbDReFlgiFEKCGsrT7wtveRi
roeFuiPRFVvO4uKkuwKkdDWH3IExJbfkjkDCJw5hNG1txeDm+5NgdCmekDP8bcqgagWhPA+MODdA
pKnpBtsPLK/LnK4LdVuF5sqn4Eb39tRH/p98K2H5SbQsy3x9vif9vhcHKVn68DZO4ja7TNd96peG
s/Kfanr50vAUOVEOn8cZY7hfKplb0go3NTtuyvz8OEzl3Z5rAGCAIrOw1Nm3qMBMtM5QvAVbuRaI
sxFDV91Qqj3/gp5KOuJgDPtNBDDjacyJTBx5kmkxsJPEpmadPP2yGWJEhkY6Jnh1MWNzSf1egyu6
1WKKwW04Wwqf1mEJvlo0F/jtrvlA75V5mxMe+AYR+onG5MQF3TELDYZjvF2zxykDx2y0B7cqyW/T
qdUUmEgizjPu018toJIRa9yFNztD8wDnWYioxx3aRZNlpcytPhQd2ZHUMhS/M7kHrO6f51rBg1en
al5gMMz6t+PCBEOtxr2Dyv5UQJDpfhPsUGCSh9TlR0ptccvmLvbyoJVmY3q5o375VN6YCYp5EG6K
aeK/5AWn9meJyjwfEkE+s5s6SRgoTGweHpgxfbGnHwvYdqGjumBVT7Bqz5jZ3YDlB3aSwbZuFToT
JMJ0n1B955ws3jFQMLjTjJIVwBXb/4nKVSPO6v/fY3KHNIU4jYrxFot8Leb+mM4skP/inaylQRdf
OD0n1COp/CpwHewO3MseDdDolxUKXAoRADJaba7pKZMSxPa6q86cyHL/qo2jj7fPGxmx5TKuXKck
TSlkOLo7eq2EUcXwQ9E7A2CH9OsDBGytwJ7pN+2h2sYIov+Y+oee9NdQFm36D5Gd3sP12aUOOoxx
46I0HnrFpw0nJjQ5YB6ImriwKaJur95huYBHwEBgxED1WDe4AyEIu/Dm2wEn+tiuMglBL/SKskHx
LhtIuraPHsPX7iwk2+hRaW1RBGAcA9UgjGtnVMqLqbyWhlL0m7Y+FfoxNzpApOY0q+10hXFbajcJ
wXTXYMAsEVS7afYAaZ7VMCqmJdcW8LP/hxyK9ecS1va3YD5SYr04aLaewjsA36/5ch52w2NSkyDm
KVKwriNaXgHt94mHTfxNljIpRHqKkI3pnT2+NrvC/Me5iCKVSlrUk7+Spd2/MFPr24KO6uHcIdEP
RV4rTPbYU6/3Dg0TVrYOBI9LUKfOh+FKBO69pTJ8tLv30hTV8iTEevrRpT/mmU2nMPXMZyrpyU1k
grr1LcygFb9LeKGVt9slSgDWb20QBWyXAbiPWDkSCz6+ykNwjxe7W9/0a7g5Lu55V7n0ukvyo+JP
n1VWpzecCf2p7gZb6D4Gt8Ed9nmwp92KHSsVp1qrCwU/a6DIzx0NKUDPHv8Xcav0NzIgRczzLA/5
JWhqhhjgTVhHMV19oWtWgr+9RV9JxR8RZOlSxFGTJU40a4KrIO7yRs+bxW6iNR8Uxg/J81MWPefO
s+RV9pTe3VAsnqOQUh7h5/dwWL6wTF1NyIae3sAlNbCXK1Px2dUD0S+qwDKKZeOj3P4Q7GaWJLfU
BWtuTJWIses97rVhP6UZdPgYNfQzM6J11WYAMk8qvFmt/lzNAL6+NMyvUYqjS8tqR3P7j+gN+AcK
MFTzJY+QuNRYc/Kv/zOa0GoIqG6pp8hb7TkyGXdk9dBDzLbcXMslPNPDC3S11SdQ3h2wnlLVP2b1
1Xh/LO6yTQO3J83810ILqRsOHGGEiD9/QqtybydaDeduQvukUVKZJu+sBFkrIyREfpQFeARLL17u
SJqIEcAcR3jMnWWUaMZudZ4Y50EtN9zR/he1ff3fk2+4mt3XmX9S7bXwI7Q+y1Al69mSe4IV8w4R
Dae7zw7b/UvR5c0DHEH+zJMiSPzsoYAeYhr7WfUO0TNAk7Tczm2uQkFQTu9/6a6ieRn/0oycAYdS
TMMZXMhoNenuAl3MrsZpduE7lA7z1iRhwo6F/M9qgNFeA6GtMO3LH/njFJzNZraCqLVlA/jNZKS7
P1T2rfiZhn/pKcO2+47DVNl6Q9Oh3hH1HrLSMLiBxedmBTx3g5ITpJw+WP3B0uGnun+AMPLZe8Da
rG78Oe8sszSFTzcxruZlsOcoLaevo7+5fR0z0QYU8tMQyywvdq9kSgd+UGvQzgYg5SsNgX07Kyyp
aIIJ5+IHYRplee5KpehiK0/DaWvHmys2Jt7CQ+aEsZ2i1UHZ7HZEkSDV1Rv6VRdkphV4vHCwQfJR
74RUgxQKjmpkrpMjSYAt+dxYZ20S1y+BkWyw1/ehMKvuvjkmT2hihIQ2vHM5CHkVGOYVjud++zGR
/KoAj/TC1NOfyHFqp4Z+FkEfO2GN/dNjQ1/a95xpMg9ISS3wsP9rOIINYLDYMcwXxO5boVjN/YOI
1wuVv4XEsIaIJfp8xD+N83Sfub5wdk5BGNLxBx+My0DkMFTwWkYmgFk7bk9g/JiO6fKFpSnOa3yF
Tly9uyloUHiPbwtkwcx2yV11aFzQu/+tWKq+kxDx+aXADqC9SQiHY104FTbIm6tPJ661OYZa5Fqw
ajL8VsxQWrdKuZ8FQNHuUihKnb8elIxVudbm6SuQtXQoUN+AOfLE8YbiZSWPpZSpaFmVHKI9aeq3
SLHshAq6Mx1/OSP4ctUAnvq31wtgwjNQF0SnXrj5of7ehP31XIPlJ/6AByXXC45EsS2tzSTG3+M4
c6Z2aMcyu1h/Qt+WdLCytW6nPMPM3NLftZp9WfiTiAPxQk+IZgLhbJCe3fiuIs+oGfzB9W1GILDD
HltjLfQR2RdU3kYsO1U3Z2gbVxwdmXOO8itp17bQuN3Lnvo0oMfpgLlSs1Qe14pO/1NnIy2goaDj
HV+XuxbfGQHtp210IpWSXTAnHCLDizBzDQxRcWPbmoNmFJA26AEVA+R8PvQ0TnJ4X4U9EEZkHlPJ
3K8LRwJ0AMNQ8bK53VMJ9nx8qdmqkzF1FpNfegqwu58nMby/yn2QEV/p8+6dzPKPxEaZ7Zt7OoFT
2NIUD9m3jqGdIiRC5LneaYarxOoVitnDDVBwF7PuHIG28lEV7GGmoCLLMcEIca/ID8U29tOIJjtg
5Rr2y47L0ufpaTDVtOHl0IkRBRo7jXbVbqGHlwZZth+v+RGABbjbvYUW7dzK/GoAdSAf3AMtm4th
uIqgtJv46g536we0TeyhihEIGzBTQlB3ENDJYbI6NiDRUHGuHtHEksmeNCrkuBsz1Z6RfxfVNPug
y5BYMHIC7mHaJkmzXIRnCF1GZp17qWMPRX/Bhm7IedLEa2PBp/kmYuRJj9AzeM6Xjk5nybSFelR8
ZevLNnVidD3GA99TRKh2dC9VgvtBXfPpPbeEynBhT4lrQMbZWV0HFNeb+epohmOXQTiIyO7kubap
cNjXJFv5NBL6gkuzF6kT89Ez8bFNF4ru4HQIaCX35rFo+cDRfOIWruVchoKG/2zxPeHBN39ZvgGA
z3Hz1EcjDMDbHVz7IaZ/CC9KmYUphvk5Wyp2XzibiqtSmjb/LTClqFVp7w+eVmgxsp4xJ+Tg4XdB
UmJNebCkd4B/5TqR4SE/ImrpLN3bQbU67OxyJwSTh8r7D9T0L+Ap8eoQ6rj/jUfQA2IiFzJP5vGz
nj8NDAXcRoQFFKgGIT0jBMziNonVt0i29Ts0TnLZofRhknU/MI0MXW2Ij39Ru7JOg5yReLnK4u+g
+dkslYo/OZa+5MRKUVEuXoc0qgvlidKFiKiiUia8ViQ73BMwy7G3BrNGCs96yPJqO5YqZRlwTcz5
2kWCmQ9SSaof5KGOIl3HJycxC+FHYfHjmuVWXnARsjMhsu7a4AD31icQTjdrTjCNJYJpLXsTflYs
Su10uptX+lVGVL4azg4Qd6KlumhHtTAZFwSn585vZFi6e2eB7dyuOS9G6VOEcNRnlmgoZq9I/9n+
5K30GYePEuOJQyQhEa2jrDY39BbELX/et5p3nTeQbSQp5Pcc1B0oCjMDgxgYP+/JRS4p1Alt3yv3
Zod4Un5BEgslOBCGQ3awFUkvR0YIpOCrsDbcNp9vjNklMCi9jy50vhJPEwOgjefs2s9xnyB9n9KX
tPDcLloq/CBdcX0DW4JFFHbKnKv1TDyCF3J/5qE6zQxrVp8pyUA/GLQAjTmjTOsNIPriN68zYPpV
ABF3xCIGkih7R0gg173UjPQGG5V3edY/HGt4oaFNlwABID+AMl/c2hArpkeUlDBX7NbaxGPSCvg9
+nwEyN5ITJFBKx8tLU1yV7eLRYxhcascGCDLQGREYoU9fqgejjoJF2/dd0Zpdj2NtDU5MvWZGHqs
uG5EEJaJak+ywPGZeK5vs1T9v+pwGRuku0HJWml4v7d5PPVfFFEU5KMFzYV7JlbQCNsaIXP/EaFQ
9lvAIMohDZ8RqDHh3oTP4Ga8tZkLf4NC6A0nYphDHWEBTAgkkq0cdhH1wms2PPitTTPPXufRJqwD
d7Jlu03Ng8KkBwzx46ZMFGgr5WLCsylWvEI09RC5MipZwItL+gliQUopEpVON46N8wueOiVX9FF4
jcd1Zi/EbeFyGfa8O3MgD6JpJTjec8D7MN6tt87bfOBkUjvFXxK7x9VuA9msZ8bWLsarQKFkBMQK
5l2Ms1LNzze/TSaib026AFH9fT15bpvCvcswsM/9rbszzBvA4ICreDwGTagohwhIIfONCfiGrZz2
djVYNZvt6/jptxrKeq0ZNe6G1w0iqmC5Oyk8iw802fzcQzOIQOqJqMgvV9akDm3SczyqunqKYAvS
jV0+6CW4lw/ISM97dRbpXNFy1gpNqVyeBKvqQUsrgaJJfsybCWis/+bW9lZVR+4AJnRiqFWXYIw5
fAdAwXWYzlQNHns+aoCtZXLF/NY+aRAFc3gBBHpvuqDDQoG+YHz50FFGoIsupReyaGif01p0xFRt
HrNZ26Pe5FVxZoHLAjqOjQZvT/YR/4UuBen8LxkoLDvaKSfgtpeEa5iPJqGnUNyLohuTrTRQJgLT
1ZOZSL3AV6GmtGN7qOwEJqxPmYUaspESu2It5O5pJZmbMULhRfFb8lL4N4YARHY2z+cJpJJVinj4
DLDkJK4TPLUFtRoB3nvoEf+p+4NJfUFdEu/axVBImJ0Z69yxQJrfeDmVbLyu9PfjWa4Qbk+ToSc1
Y15hvRW/c2pGmWvremzVKHhW/oJttWiQgZJqXEzv2TB9rtYDRb6mXI4c5YfBK0uYyCTACg7QyNGm
f6P7GvAdiOF5vSUZmBcDhvsXm4D8xDLyN55DW+Kv1YH3xdfm5q7mzwnVqqQiFs6C8/kSZ1Be7ZWg
5ot5fX1kBWpMYoysg4/6A4jcrdNDfrNlV1Wl3LNjqm2mQnpdBIUFi1YzGxjIxrqfaHQpUxm1c5o9
uB5Lj1N38yuDGCdSgDJLDsTeFRuLhjL2atywf2xKLiMTGX4TgSdFCXiUc43oidS008+YljOJOjfp
RsBVJBPxEiiUl44Ih+Bcteplnm3ylDHbqfauiPbMM17n6kByAjWEuiPv+62uYEJI+0lrIDE4yDho
91xfVskup4bWPnKntS+cdoAWlxmXKLJbEDiAa9+M+ypyuitNNTgKVy0RX9+p07KQkc73jD7ABgWs
VMISP8F99Cd/cRCPYq+HzT5mQr+SHzWjdfFuN8tDlJW2hxekKK44YdcIUsgsV8/zz0W0e2cUZSUF
Bxwrcxly3mJDt91oXgpD+YQJAUWIj+uKFXftmNn7EZuViZjz6J1oGhzPP0qbt8eM5mZX5hSzgXkx
mqWf2zs2BvTMk1UseTdwwJB2bVGZxbKcOXCytaPrK9isuCVpLLxKeS2GjJHZnWDytTWpztB+xhZZ
IRnZ6ruOBTa2e5tyOeR7mpTem81Am2XXHZ91fR9y29aeOQ9fIeEmSLnmOjDDaWLZAb1nxMpkTPd+
C9wHs1DL3tSSOcdxUf9u7O6zCbc2C7z7ET6C4iL12y8cz6dNfUQ5hsYSp93s8lLaO8ESUVuC2Tsf
ENMTBexiZoxz6dN7jIi71mpiijkxRR4D1RDBvdS4R1pKZLknt8EhQJ+ctC8bHARNlpg52PxYCh9O
CgpJw4MUM3iLA6HQS27CZ1ysCTXPtAM12gazsF75VdoK0jwBNh1p0QLcPlINdDOrTKXD4iJiJwFq
gNwVLAlVdtyXk2PkyThnir0jgSZGSdAb5SeulidKWOLbT4HG02WiMOtUiTeoczlTe3lGf4QAG6Nw
3loM434ltaQB1U2lO8X16BKrgJx9lBpCZbdtSKYGnhYayVXvS/iOfH0OXKo2wmu44GkiWDklCvPX
YXsjQYItbEYBjgt5EmTiz3U+t/1xSPW4LK641LIJjeWvUmoAAOFwoIKX/2UjgvYLgCDrRi0zW2n+
9s+y5ppe1H8pFHhogCYh8+5u3QpWGM/UZ2o00y/quqy6TQ/dBnqadIl5k63W4FzfTLjl25juBa9F
8lyNnAM1TfQ0EYVyaGzyhdtrwjocNgXBH5QAv0DdeF4UAU/BmcsM/sugQ+0ylXD6eEb3ZCrUlr8/
oXPN5qqmEqFm/y7iu1ol700hKYt1RcGKYPOKNu+idOPNta2PDeF4kl2QIetkz/aHtZFxlZapuapQ
muZuZKdnBvVhMEI48f73a5CUdWT1WAtIVtZM6WUy2qiFZG9eAfHSvVEWNPFOcsa0g4569HLo4bFh
k7jvYYkEGueg3avvO6A8Dv2+buQXEAlNJkkvgtilj8fSMgNNjF/ijaaj5xu95tBSvl/hC26vUyxe
xBcgjbA39mCwnBAxH4dfAxrLRQ4zFKFd3oPvRJkmKJNtJKdVDpXkpYRjITKOC0FxfPIs4pIqrJEf
sK+QoyRSvoIgf405QwQLbLiVJHGAJ/9YkvR8AjR99duLurSXyHVRSG+ZLT/WugmBtNNK+T/mB95g
I+Xt5Qoaa6PG13i0iZ22OTZxWU4HzzaY3Q+mV2FVCx5gsp+hddys/yLJDOYIcbtlFo8747zqMLan
Njw+D7Tp60dz6Hs59Z9cTYD9Mg1E82pgGA9ge40qOZkvgRmykJqxLS7y+hBl/dfdIRjUxL7CdCSt
8AudCUZNpKSUCSGb1/3+ZWTeITUwLIxXlensbfX/RVwHwpD0lij+s+HvZnIqM46FTqyf09QGtwQq
PKrMiCKTWB7tVZuzsVtnDDhy+2Q5KS0oVec9xvI6rrr3g0pZ8sjCMF4tg5et9STMqVZUwdC+B99d
Uc8PvevYDEF3Qh086yJXG0fp1USEdThgzG0Lk8nwMIX5hCb/ULUoHjetAxYUP06uwKVP2DSyEgEs
cYhZuK9GXPLjZWryfM34HnZeQqocOah65jdHGLcFKMZ7zOMywG58eSmLDa0LF7QWK/BdevtN0EHo
HAA/ken47iF2OC2KKoxmjRV/2FqhDGzgDlyA80xEuGN3lnEC7RWbCm6tIu6MmZQBhi2ZrBQYgxo2
Ac0v+2BMr3RmJ1TPV+1EzKoBHZygjI65jRC0PZZn+H04qx+YnXSl5UeZFiFZrOFR6zrdN3ogeWtN
GXOSsSqhRAcRd6BhmFlKt53PxLvImiwu2c+l/DUyA5A4OnU8FAdhPUzzuJQZQPzB9Mkpgz7+NLAC
IOahRXGDbSDSac54HdEKxs4RCeuEpvRi9J9Yu4VnSZ+A/rwQkc9Yz0pL01y7NSi/AkOf7Jg782jZ
NzvWI8I4QHDqdb2/jYFD//9l9d6pM/vTF0aI5dkiitXVNvyL400UQKrOGHW/jSxZIqHyysRMpH6j
kht7wUKma8Qr3oeCKggTr4xivr3a823H0XEED1zRyg/XhP+fQCkdLLueynBtPcllTFYc58c47zwh
mjQ6NxMBB5++Is7TJEYAAPTFjCJ/l/E5898Wl2INIPk5bcA/Q1Pk+S/8l1ZZ6rRxG/mAZhdm0k4f
n8Qm30nFuAwdgf1kpjhXxdeNrwC0b+LeJ/USrttmVZ7RpqXZN0+hr8UkaY5/oyM/htE9VBIqP96f
i4N6trbTqpm8b8HS6Qhqmq/8UJbp3dl2qqYo+vPceNcflurR/b9TLKISCHlkoJ90P4mCvrFOlA5T
nnWLTXioWUCo5TqNtRx1MwNQ2bwjrqy7ax4UT87FE7Hx+bMKmD1cF/BL+P+VCADSoc+R1W2TQ9k0
GlwbJtqjDnRs/O8ULlOtwTyo36HUt1HENx85Dfd2D+8ggbo7yt3FwtksNyo1c8jZAfDFAMfmbrmq
Hgs9hUoScO5u8R4f39qp+pOuxQgHqfVoqS5LC70W6o0SCjXFKzK/tM7hTFi/dR54ECs6ncqpORck
ll9UuT2hNwNwxnyFdNxmjcPpK6KdsUqlCSvM3AuwTt7PQO6qnVZvRDle7Rg4PPCnBHSShu8cEveN
Mqd0525Qzbcglc4PKF8OrrMB2G1VJE78Q9kuWzloL+tr0h7sO58JpOqVDGCnc5uC7zGWEfvAe/dh
n8V1pmFyqOgQlMmNToa/3iU4gIwLS1cC/36TZ4vrObnlPoi/yh75ZiL6uEpnTHzxqsBoHB3O0lMM
yzQaY7d6ionhH+HwGQv3cuKXuPKwt8ffM1ZZ9VcD5J8EyXr9Fo7vJVCx+u3WiWy3q/sxy9o+yamM
cMbDiiHjkHpVfyneDfY9Bmf0Gh6MZ7eZBz2eU80tkJcAj5k1VppQfVtPYB8fhzm5t+zPGrTNGTOw
1fQrwjImi2Tal2ZbykHsOkQi8a8m24EEWiEo/70b2ePJvjPTN8UlkF+DsQlVb+Il4DWGtM1y8gbT
YGtI70OhXlKBpyw9evqepcCAUOuo4f40/PBEYow+2Jo5qnac6JWP2wVDXf+QFmHdakjTbua7iuYm
fm1XKrZxJXVZeXU2XO/WfcJ++cdaF1r9f9C1YksmSM3HupUyHHbB2ULj8F7eXrGBmTMi9oTbP65Z
gOmBHJU4VYKLqfTwAJFJLPJTr5ogTmwr6FduVVeatIe4c3+U6m7BQYf/HFyo+PdEoPKp9CAl5XRm
f65WEYeEhj/9ELsnQispc3UlETQGizLNdi9Gu/vRDOlgWVOqnmxcgxEgPaiqbIBycP4klLkxsivG
7SZiGLSLRakn65JoTaJfXutPoNf3lhCN4oqD7vc1clt8KoVlxq7KI2sA+ovQg2fQUM3L5Zo05rPb
XVGDZMW7ADdmUyKqZdiccW0DtUpRsEzYvau1d7VoQDDNrWSRXi7z5+UYzJ0UQdZmEHlkOixPeCfn
KmaMPWrxXxCKxVjHB4Zsr4c/xM5ZBzbLwR6hLEOU6ceQqQ33oe7gPN2SQvYOs2uicmsk2yM8xbgz
Or0GC10q5KIRczkOR9cRLveLMmQs0M540C1C/Rs/tAnNWkpPSMpb+e/yFkVWaC4Qz8dq1M8txTCi
Pe+RLWcdSVQhvxfyKgM878eHcJF6vqCa7uQ2shEaVt0zdj6X6o4x+OfTYkI/RX03c+gGSSX0FT0W
tHnogO3gUP10eGE308Wyt0t65LZQRffWB4dMNGYJJ8yC00EdIOy/yGBw0jVVdthYFYgtKTKe1PWd
ba4Udb88bCQvNO7IcNSAXqPo6tN596nX4xcII5xMc3dpSERG8bldlMo/bYgfprEu1m1dKzSnK7dr
LAiecuXzL8Ga5tXSVJN+04XDkbRrNtx+yuu9vqxhMeP/YuvThnHiTq39/Y1cV2EtkNETUxQkuZG2
XrNCWbbh4zabkXDrjbksGEZzNM7rhJo0aEWZJmllZXBiT0g+Hly6P3ig9rW3zwkTFGQfn83b/BUf
P6pQ4GAJgCtixoCs8IXV65Z85w2Qo+Rg/BnAPUwZo0qIh4HbPJBAll4u4h6WrhYvyUIOpHnGu8r7
ELW2mgUR9VP2x/AcJEEiFJYsCrJPr+Sdmub+NFxDqNwGsVTQrwufKyMDaFcP4WR88y/sbEtvrQo8
HvYTr+DulEPMVnJVZmzGt9tFqK0s6oUivwL7TEayraO3Wq8BpaQgMcjwGEyvqoEkOTJi1V1qiMc9
sbxQSz9Z+y/WO5Bvv1YuRXYN/TWvVEK38FzCuDLpuMLvJPHWVAZig3Xhtztb3I70QR9LvLTjk3Gl
bjRo/a+tBeQdAwbrL/hd2J8hruqO/OqHfm1QkQInFsLrRwm8HyXh9gRvgkkkSh5ZIknJnfxQAA0w
ZJXEfPN7jSWxwWvdY/+6/aMPgSxJ82Yp+lRSMZXlSjmnMPdp8DMjYn8FKtYdlgF4yi7ZBa3M0Q4G
lAlgNQToZRlZYI7C43bb71MMnK7vkOfHw0+k44JpZeTektuzd6pW93FnHI3LZMYTrsoq+okjRwhV
uy+ecoW021bolCSTbflVk73D92JWbSbOlzArb0M7/5FlCObVtzPb3/9eWcmYDIPPwhwUheyJrtf9
YPUVwGfAMSI+fu+zG23Q5hOxVvVw0Yd2SV3rTD93kn+AwUfwfOuo3D6XOUU6VpUH4uRGtJRJwvvG
7Z8vRMG/GbBL4Kb1hc8HKQn39H//JeK0NUna+cJx8jXpuHqEzeL7S732Lup1kaWQX/q5QfYDbhrE
hnWtQHaQhvUczQ8CmDZw6KvyKbSKTqfwf1JT+KiF/oEEkZ7W7MRMmO5bSBqPEsJmY4KAZ+T+5Sp7
4pRMXCzeKgArKRbL+81pCMQ7F13JIWR9+nkuTqWVbYr1YiKxbFlOnjsBFkqr8bT++USRl+Cf9Oi0
jF4Y4ndZGvgiQ8vXeQ2ozMkhpRnBkeat82w1F83FmUhyOkHjhevbCfUAgs8W+hOoULd4JNi/edl5
CmC68rNhapYK5fLWaK6eO+k8JQVtruBV0NTIuXoKS/LjGaLdnbtCeL8rRVSuIL79YvglNTGXrEnl
Ezh/sZTbq0mtSuiwtNt+rCh2YLQWZ60J9HyDca1cvQUu5ezAD9NOubzMx7ERhuudXi4GOqJcGq3p
Srle4lPXG8iMFvVIT27VAg9re/Jv6SAD7SMHRnC0m5lL+pIdFEL3tiyLS7wIs1kiOISYYz+c8lfY
A37EXSj8Xl7+vu4qjUEvxykuuyu6h+VToG+DtjQl1h2t6X4WkSvgQXamSJyaIETpWAoCnOlX+d9E
sTP/ZSV1CkgSjCh/9ERaSMx9R+5GBGD0Pd7SMtWA3IECFtjBKaENp7YT4+O6It42VNe7iJ9c9wfE
hNPI2TWNl3kwDKjw/o4NlPk3DbVMFnIm0xf/3YNrLfVLx4TCddIqWC9QWgSyhRA9l3UcEzMxpGBS
GgN53TMdvv1OnxU+VHTRh6spQpbxiRchtItO8Ln6/RfeU8Y9R1RuhgL5TwCRQONK27Hrevmc0kF9
Uxpgs71w6eNSGUmdm30M/ludIQA/tnOtgBaX2TbCbcRap1s8jwO7cEchp6wfQtjQHcOzKvwNQbHW
xTxa5kDe+FEgnrT/UwBUHFJt6cXOhZ1rD9qQxDqUw4u9gYX0nRNBi8m8WnE1Ku8R7t/R+DmoQGui
sHjS+XD2DLmzA1ePr3CQ88REqvOcnQEKg2ZMBlZuYI0LtcSK9Hoowf34tyHukaK//+hz6g2n+nE4
60wL/jdH90Zv2qtj7Rs8r8c8chR0zVVoRG+99Pyi7XTnZ/lQQ3Wgdi/dnbxNe2svEVr1yrMWgE4G
F1F4LsAUsXx65AIMf0vZBN1/aHi1Ka/rkLWVjxjglDuMCjdH5Qf1Ej8SjvyfY20DotwvcYACNbeq
fKP4c7rssQnEDWWAbAJjSIsKMDbbeZRUpGZFYDT4vSPd+Gb62K4XnJMJoK3tQ9/tWRYtnYuTun2F
M1Jv3nG4dZ7TGesUm7Wg8stUyu7yrfxGaWuRcRkS9oNVSS7XIBVdjZcDaAbkSjFDeKhwl3KiffH2
3SIWjAJaAPRSHpO4dRbLw36XMQgrALAO9Kb1wEIdhQJZIYYsrHetEihR6Ltbfq7UEB/iUeahul/F
OZzY5g4p7fBC9l8ZWjfcItqtlNR5OxxnsMIqiHSd3GhJHDSpCTzWnqgNR6XGtzv97mYcngYHxYD/
V9SYkGDMyItvCJNouRHgT5Fngw5wbWZ+dsTbwYo0wSlDjWBDkIuSjNeUvls5MPNmyoLS+7Gr6bFV
73iGp49BUAPorbnUhhfO5Fh7kF2AMsmWbqRB3Uq+snh9wM6OZedzlVqkGxTtXhwUzuCXDl4IYRQh
q9RdA+rklLvRiY2L0KyDFEAPQHOGtKMmLpHJmgnrvU5IfgCPzbXWRBa7oBgHe0fC1fhmIZI0xWjO
nAblonh9YAvV/JdS2shnpluxp5cC6e58Y5VbINFoMtnxEOdfFMU7Svq2jbfnIMJUcwbPUXgxpfqj
KOXo82EpFxtoJjCjmtKllyosiHyTp+9sLGinWhy9yYJ8emBtDFf85MzStuTKzST/dxqyMXRxfG8g
7WvWY2YvQic0cKrEVRiNElwvZzhhs5Jifjh4luTYa4e5OEe10crup1BfcMZ45Icuaj/syJJrap9h
vdVMNptsrWVGwyhvCBalVwjzo2Y0Fz0a9kMDv3nVyXQy8kiiQZrdKxtkUEyMcVDpILzbKazsgOvp
SUDSVkulNJnWhpuuC3AvdedWSysguyP/ji8sQyJqTfSMv5Gg8sWmo2hQtaf8x0ICnpiQsqfelGY6
5DsYWSi2HU8gWiUBIhxibWqEAl3swZVtLwKWycMeGxQciK7oVZJF01Ev8JguaufMsH0SCr8sWayq
CBESZjNOefeIdwkVpMZjOmtl+rUnbgdoFbjGE67aI0p4AxSsypzcDa3uScUtXUDfWA3+jFYiZNjr
w2CcgPFg+p8wKmGVH9iAcMk94InwUPX7SX2TqikRhPqohn9WSjPeiPt6G9vWicYYcayb3yRJOQdF
WztF5fEKWdHdxTxWo/BY5ASE3DNcjn62D9J3WThn0Fb3gIkwM5ZkgLWhDUxxoNlGIfslTEIy3aFR
CNQKV9b7L2zsCCG1OAJHKW3st6uEzL5KafX2CWmn94mM0Itjz89ITVUhIJ9CAdZlgPsYoVH+DdiC
ZSp5f1y66EzkOD2MioJfwWj1k+5OWwWy6owsIII69DZVJ6Jjro/8g5yH8F5ErSto2ScSxlc7Y/Kg
kdRfobFYssMfeIzsYSr9GxLtynlf1K97XbF2xl9gKmuCxiwpthsVBebcOnVTYhn5fn+nZDanoJio
35CmjpbcB0EjOlW3fLWQpj9ff4TTi7Np02dWySbMn2Rt7TmCRntDqRwie/2L90GqE0IKws+pQ5Rp
xkG5JAwnyVdxAcJOf1Jz1sjbepONFlj5aUdiVHyHTUaU7B+3eoslVQPWL3w/K+3WzXtDXME9ObO0
cL4oPgH5sWlZSxho70mIcsxqsN8vWXBbht3XYWZg9qXo5MHkttXZtSMB47QDPKk0zHy2Wg6nAkKl
fJ961BZuv88loVH8Sxs5XHWdIraOk9GqSPl3sWkTsnRF86aDll//bI6U68PKC+9PmMHnQ3Xj3v+e
7VJsC9siESR7B3kmRsOBVYiXzi7A7AFSKbvIzsLekjM3TyQ4bI2sAfaWWGTUEKILLZolq1Src909
B8gJdQNgfHoOrmTTH+tlfsy6dlh4qenm0C5B3j9Vd8TCMLnftpRO8F/gZlKJj5v/N9U0wC2USI0G
Rg5EE7xGBExqBUaJed8/4UVnlXNpFKRSK2FFY+HF9sa3PKwcxAa8ByEuvElIF4V8Xg8bu0XJz85l
3s5dvWjLjL4tBX/So3MVDjWCKJ1K1yHdWM29KrCe5WAYnbndLUqZmH1IHWP/0zijjkhC5bPJVV3M
DynoqkkX/u34HKrV75md20d1j6VdGgf0xOcteKefbN5Hkc9pLAGhiBrbxNmNIwuOgdFRI2JAMAA+
Vq6Iraxl8wK7Tn59WdH9UgF4FaiIW0ghHyvsuUHMFWajxAIiOCgVYH+9thUW2mfq1/2FlDgp7Cwu
+YEngt+tcRX+dYAw9PsOrPV0/5/60mQpIGHBSXRbhHLHUaabRHQFBfF5zOJLplrpCu6NqN0ilyaf
GMBLe8cyOfdr/j0f6P/tHwZwuOFM8fhcXiw7WfTfOQd5I2uyrK2KJWi3X+sUCWvHOKMcxOXasowZ
HcH4CmSLQpJtmiPcAHB8DBEnyTIKGO4o8QA0Px7Kc9pN9tvXpZce9MuLA6rQRsUO0vmBisgdKcK1
oIPE0u5MA28xTvV0PR+oggwnR38QVn+y04EfOUOaW7QhtB7CdLbbN2C3dC/B8Tyl47IAMDtwPiWI
9yWq7lrqKcxQvGst2XDU337HyNGOWTA0cR9vJto8PIxgHH8SAGWI/tYl/UvixsyzNi0IOGlgFEIx
XIOL2SrDlkRGwtxcZlosfWM1BimyFSNx1N2B/C9bikJFAmPz36BLBcRWufCxqV3pQfI//bjqAHvG
O+fa5kEC276Q4c7kbUuzmYgN03uY2ic1a3qM2J7+UGB7Bo4tSYEK9mwPqiHfOvqEr9KZMzH3xKk2
5svu7fz8SdV0cjFH1C/8/WA4BfP1og/lBxDTEPxPZsaTzhNJEkDF7IFjOcS21PiUw5W4WV4PGyd9
9OHFntjvPq53JZ355CIKFuyzYrqDVKzwAg6oyx9jBi4zPVy+WuermWrRMUCWZ7msKQK8fCcgO67Q
3kzJDu3SnyECM+Gn41Cd6umBblH4o75hlLdN9cvq7tgirUJZYfoN6OJSw1r7JeyYDFxjkeCV+6tJ
a9t3JF/DbOpdVYPSlCmDDE7JqU//yZJHeHtdXpYW1bvG8khEmgUBzKtmReDq+/C06fylbNVhQVe4
e+HXuaOC5oMnjHdEjPwySL4Iicfoe8y2FcmShATJbwHYP5JHVB/2EW4NOvaWJO7AINgtq18pHUwR
fkCvRJKnsIyC1XjQcOkYurSmL8Py/gZ2nljejlnE+6Qa8UhGvEY0vGMqLk2wfABbMHtBQ7wzKnpN
sEW6jp9GGVnwOa1gzJTuHE8CD+2V/CJm/TlmfjNXSOolpm/pJbBj7GMJdL0pZWtnLstgI8mxiV1N
VspZPeouHpe9GLJ0DHKWUQIT/3GR+d4fy4BHR0jOw6C8g6KIqq/ybOONGSwhZ3BY/yIRBGI5mjAB
d5KF6h2N1F5Ask+Oplxf3NX4k6Df0Fa/UhgzeixRlwvL9ik1yMPjsRJm29zR2MoxuBNVXvcoHTxk
e6K9851oJ+R8D30wzcPpBAPZph0GdMSRXCAqTo3sJYnMjIUVbQLMTY+qePSCqMbyeVn5eldeePHt
hj3sZF52I2j453K/iS8vXR1GpTMDL4xi9qXXQl4D6f0rjbYiDgmib1Js7XSYj8525R8V4RsT9w8O
sO4NnF01CRsHVsR9qC4AI5Yq2TsuZlTGYEwgyM1Ecn7EDz1FAugzH43t8BGMibmd34vE/o25UumP
OkXKoXDilx9uVmwYrX4bGaUIGqqSL/vdatr9QiGs29pZtR7gIbYtg+kRwJA0pqnuAM8UqiO8Gf2q
uT/PU2WQ3BZH0RqOjdDpPnsNMrCawCL4zgG6m2XjsF8sTmQ6kpWx8XUTGTPyJRsPS2jo6Q/Rf7c6
/TZ4xs8csf+cohoRC9R7fwalH+9d9q6BkXbGSdo3BP16kCBe20mFf4pTkdR1mu/xFuo9vehzqFU+
bntarxS8ZXgHN7/D7QC4YFjNo0nZFcm2jw/LXgZBE+l3bY7+R0DlDFTnvDjh/nSaolNGQ+p5HWyL
7Vy0agw68xxS1MHdxTLGi/fzi4PzJAsc5ebyWJD7QHWNlQAbddc43XS/lXeF5bNkYNbwBvCrb9HV
i902efPx6sPiiKZrMhthqg1P/zJOoxCZafA7E/KdpWOGTDpYS/tQdJlzq4i19ayULATCH/K4cPNf
F6GG46N3uQOHUE/Nyb2q/7eDKwzam5j0UxsArLDqKvRUlgv9fwIP872cOVVhiT5rkygl/Bh0nL8O
P/G5wBmG4B0jHUQwC9CTbkHxdBki2nBFEqsv7GU/msN5z53lZdkBms2FXIA4iO4/ofi/LHscawue
adeg7v7Tocd2DvaPjvhb7jr6HhdkR02HS1zStRar37oVGjKewhtdmZabU/rlJmloI6THf/DdKj9A
g/oKsb1oUWxOAg/kD6Xsl8BSKLWkwoBBvs9pW2Ei4FAdcBKeDuA/EkHq4Zk1pxGz8pg8ky2KVk28
W2WdiSshFFGtRVGkcNZq/CmIvsVCqbcGF7Q/LzkDteiOkX7IYiGu+/PM7JBQZBOO4JCMEjXuLIcQ
400d0sX7oEhgthY/KbHt19qSiZz6dmvjrtMgOGih4oyuavTKnrkSm8njiDrOrUPiAaojXMb5iZaF
155NqQx6U8/pyGFyPdzD6FqVd9ZFGgibbAXN0nxO8joSL9L6S4SPI6nRj9eDq8zXJ61BqQjySDU9
7DD5dima+eOOud32qg3/9dQa8ywiqrfxeGq7guf/ebE/1ptsnKw0fp89bWLvPTVbkOQfSnzpWbxG
aOkJ+fAG9z+hYdP6rvjlp41mESG4CquotEVmvbMs3NKlMprlwHbzpCDXpiLvU6KCh/kKic4Ar7nZ
1leOfcxmMFzQ0aHsVXK8MbSA/mmg2lkxtt3HV/siEnD9RMIFkVnn2iUENG0OXDKwWzQvSLK0RuSu
hzJD54JgQctewos+vdwsAKx3oqYkSbpMQEK425eXnwQhIlmXrXRUfkRgCf5hRd1TeBv8Bu3A1G17
bc2Wk730nOU5BpBnQXn7KZEW/65vSq5L8zlrsoc6DW1fkm4Bzz+GpCh1Ups99ly2cQ1j5LgVoUBC
2hY9hmIDhxlE+kcnNmDsgPRd/DQ/GjvZh1ayFaKSzo+ltbHV3aP7zkSMpBbfoYN5IbmaYSsfBqp7
OVo1rFysystTyH7TdhAn97gm7fdbJwz6AdE9/KxTJink4BJcWFckm6VmBui3OCTL538hD0Vn36q+
yOQMooNqogxHYp8Hgv1t1RYGGYCnWG4uz/yB4k/xkGAV19MWl983ozaU+Qe+QztNyZjhdrpL0OCc
i470H2QEP3WyUnhhLpjWhNWwa/5QvZpU0EtmVFnqj7pJ12S9GdoaUf340E6HtPBP+sB8TyXXcP1l
ELoN3c3i6uBHNiy4kQAnoRS3mXRhnDvy0iJ9ovnYOiCVUzL/MusrahaFEOX+VcsVWaHgos4voC5g
PVLZLyV8kwGW50h7fWmp/CkQHvGCRhxJ9WSYsaJpTRMwRcFPW3XIfXC9rql2+zQFxlSn6LPsKOoP
JQJmUh1JaJ6+M+CHkcvg7L7r6yMfthHvFWvueKh2wjR3YAEG+SbQGmVNe958x0e1G4bG5MbpK4Q0
jinznAsUpgwTKsxZryHBGWUjgBYgWO9LlxJMfIO61nYTZBwoB1cvphi/UUlyjwymnZkBKNihBaBu
/JFy5Ru99/U2Ep8+takWGaHEDnMvA3S6kf1cLO4ABdcre+nMcYoFJqwGBV8bh4uLKfEQKN9zEsnw
uGa9mBt7jr6/gDB2neIPQksVO3jkaRWs2lwK3blRj+eYqis5UBCno+oLKf2n/Ekj3kldEW9GeNXq
HGHmLEUnYGzm0fv8k9Z4AZ4EQwJVjBx0h1U+sxiXe7QuAMnarr7a8wzXfyC/YaZicwIp43zYcYNE
q5nkAst/64/e5A3StCLbV+l73Rtl8LMmTtIV4wEv0qMEQFqsnrnRY79M1EQzUpLW8h9WQrhy6hKe
YVebZPlkP04FNSPcisCXsrabcf4HjLv5uMmgzClb1N+iBLvuBeFD4QERhUPPjJ/Fv4LzwX0hhBsC
CpNTIDMwXTSzpK63ZexklVD5Fk7aKOtSJMCLRsR40PMFk7kQt8vvIbvEdfHFEOLmZ39PYEOTD5ui
OZSj1BDSRQi4RkLJSCUIZQCChRKvBhx7TOvfqXGotofIVZDI44bK4kpQASJ4HQc9I+/5Q9rSjCLw
mmJSLE5xcm9GJXwZ7YYBGntZYdIJULUSJrmp7hDLWEuaND4T2Xa5v++2THGlBPFzAx85EMO2tfJ7
qGu9MFThFDTZjXxQIS/mcOKtIM74sf4ErbyOTok+tmTPDOCRse8BuqXTQ3MqGk5gKNC/Auo2lDvF
VvmBubBLlMAooNReugz94nAlkwu9Cs+edG8jk5xANUOIKvi+b6jg22gg0kwhATkJH+a7XMJvvYV/
m+tcfQdh3yGRgqJAsyo7t+qg8FWIbmmO6uw+vyCH1qFuAC1jRHe+CtS9eH8H2Bi6wkJo6isKSYbc
sHJl/POjkyH3sn5sHbyLsxqaQ7LconR5UWi2Ts6MwORvsKbUEFo98BPXneaVZhV8DuTE2wpvB609
kIlsKkIr+EwbGSWL7ouoM9IbIb6W0+7B/sZ6HnPpnnXPN4u1G5+5ru9vaKl5YvTorC+dunP92JCf
n9TMh2JPnz6Pn/Gu/CZjneXWemh5vcgqWv3bxEhboQkDO4PZomWIE8QmF9Z3dPjZ+NnrcZnSpRgN
c/bsHGFGo0phEmZ8mNFMbpvbRk49YMrBZPT+JUzNjJFkoUgQ8m5Cba3V/tIXFLAmD0oBL2g7an96
QBx1bdMG2AfUoPsccmT8yRVmWwTb3jgH7RjymCTi8DS1HjOB7Eq/6IQOh7ZRWijeEk3890G/T5QR
xyNNM8lXNhrCt4I0b+jHIIY+xtrW6JBSRXp41/QyGGCX2H6y1JZxRO76rEam7yEGjM3miKxQH5st
jqowMHinyPuwLY6depMVm2VFml0UtcHniIB+1ddGLvlLmdTl0HfE/I32o4JMkq1wVDclz2p58qay
bPk9oyTC6tzFzgS9qr7MtBvYIC63/ZbCm//Mvd4pmc4uTyGYLJw4JzBASQViKa1uV0bZGneXlLL0
7h0RTRXR+EqEAh6ub0+FOcz5iuETuObXdd9WJChqJHQNO42L6SB/Dd3mb4hboc/imXBOrRIDhkSa
v56fNSZpnIGJBkDgrLU01GOBYxs1R/oIcpl/Piur+RVRONK6/J1u7Up5NgoajmOsvOgdq1ClLaDd
aZTALrKoeMM90tmKvOerB+u21oK9oK5ZLjmIScisIqooyGlH6u6tkdBnfPy8m540vShQSCfrHAnE
U6d/9stPvo7syoe2Ob2lV6kRCbZ7wWrEazsONvfUZdRQrKBpkk80qGTbvTV+2/tZT1PPp7biDv4q
cj0GIJyGvrTykfVlelrj99EYL7/ash64mmqg2KU8H30oUixREYClJpJByYl5I12QEYLWXrKQ9QtD
6HgS47eqY5V73HP43Psg7UrEjB0QBdijVUwzuDQJSKBgupHqujb6czhPQAOpoa9IWakrmwcsBN5K
vRzFF9OdmM3Jo2CywEqq+c2yuOor/tUsM5vpVg7FfVVFa2mcKFfARAJIZIksze86GqzG0XxxUvcX
xzwIAC30DKseJNTJoY6VcAm3zud4W/4VLnu55D+HpyZRw1fPq4tneHn4klD/Pke0zl+xjQ4dpDbQ
ho7GZvyWNtZV/FR0C1GlftprhyEoD8dgEmO9T0acEy6I6lwNQspJMM/Y2PhLJ42ndx13PCLXzNUQ
uDzh+pVGLypyri36fxdRH+U1fljMdtMzT9l9YM3iqFqXg37zzKLjH8S/T53ctrWU/OE8UqlxaBDl
0VqXyecPUfK0azaKTOsVy+Z+KNXxSY0ci6q2rko/2bvy3gO1muEKuHSTZ0lhHLYIJiD4oD36AB3G
9HSEl+FzSZ/EgAwja2JvemkzUB/w4SOY847e+8Yoi+86Kb89TCCb4SuiL3hLnpNvB+yiFrUOArob
Ut95bvoGm18h6kd5YPbd8SQCK21qFJxTRD+5+VX1QC//OKnFgvEW2BNgx6K1JpSF7YpEABUNoVcb
npY9xxM01LnsK31DUWw2Nx51iMCKYNQe8WIHHJhmtjUpUyJUFerw3RwJryhGwKdX+C9iGxMzELQf
ZxdSLwCZ5yrpFKz+tLFlB0ZYlKJ26F6UG+1exkvIKQnGgj/kKfvSCjmOBzDc/DIv/zzsWRW0RA7Y
pX4S02iYk1sOkXIUr3d/LHlOnXJggn1BXKkKUh3g2UVormC+JaYbABVDP/FntpAzkdjsGpUUm0h2
IfYxeb/J57UolnSxjMyxXgm04pnr4bP6yI6d6B462Il30CmL1NMkef2PnOQsogImN+jsbRxLYv0a
qxpZcgLS/77EZ4JnPurnKtn9BFdr50cDe57T6CDbhQfP6NFQc4iVjVs7bYe2bDaZp2/YklSU6D2y
nFViJFolYDYgCXitrP5RFbU5kxOS85zNAmZnFldw9ffhgPEC8UMb+anKtS8xmegkYi+wWAbGnjJX
dtlL0xa9jsOQrKUegKMquXRR3kY5gsXJd4oeKVSJHT0huzDOqdtzYe5SaixNaBcQn1cVNkB7AFJt
pJNI8Kv/XhIbCHKWeV+l7N5p6E9Dx4hUbZkaALEvJusrqllQ2WCV0sXagSNzPqpFPU7NmvFp3bAV
JdeOXjT6pSrblbW2slBtHjCxsOfGvQs+MC6RXUDQjNBqSQnwVLxpCZraQMXs0tHvPhux5ruqb7Fu
McgQ1cbyn5a1N4JH7q/ZbjU0E+Mpqk6R4W8Om1BFF7pnntkA9JWTtCIPWPvY3mKov5mUEVoiuStG
Pc+D0n9/SWyo9bjyd2v9a3mur70XbxtJWFIXO61u9ZByLV9J1NRKPJT4lgMzwDRRx6eVMMNxel/b
GqbbBf3QmBhSoiJdnomNZeifWUYBB9f4/oMQMkE9Y+7TJE7hmmEDwPxPNBXe9vlRQiRTlFn7CG49
BP5G7mih5OUYOKEUikejFmR0kn01Wv923epXdbVB2NbUFXMcIWViacU1yJYRRhfM9ZzklHRWPNQw
jg8KYn/nHPhNc1nUB3MfIj0TkzTdVZBzE8/AtkCyJWT5C7g3y0F73YLyjnGkWMTJ0YpKudWrle2B
eBTouZwdMbg73gDs0TdXmwvcFgqer06nbdjHdz20PUjmHGQLYhZFD9fWqzTBr1LrLZMgcPJYj4HL
Ojgehxg1W5bPkHgI0aKjI1ZCHBOxk9hMNbZCf51B4wlc5e29CuSImlx+VhjJOUuhKRaHyVkJtd6y
P9hrbWXyeGSCGZLKXgi5P2ewosCILRrLYsHPk/iAKIoI76+65APNdsZfOZEcO5LvBM3MNJ/lxzKK
ed8huZkWDJ+O9FfhoO+CQy8kAAshz/cH/fouaIzWO1UvhcHiyZWnsW1YUY62GJ8SsLa9DuCGA6nD
5/wV59w3eRoGmxjNUEzAevO4LCieVlx1WsfQ2yNJ4nXKw9VcWL6U5tKavVvaWCzyrPxxMHuF3+zr
irT2Fwhg8GngZIj1mUXhbtuJFyqEf85IR1Mjje1q02grw0g9cjyKGpDjwirWwDyoMJx4EHSXeQ8j
Nc1Oc7IeSoC8QY/E0d//8/u6aumLYC4CvsDSW4hVTSkFJMcnW6ZpTBzHmEgzg6Ep4SHo2d+0VG7u
UZKGzKrvMidWlAAP0Ygejdp5zvdUSx+E7H2AK9UixUX34u0oduUIj8j5/dn0k4LubywGO69gGJfa
XYllq1WoO4fYfzisA/nkEyffArhuHIGXXz0suqj4wJ+6nTMpKnGApSS5U1iT1W+3Zz9LZNBbkcRg
XF3U9kRWZkO3jlu35S5+iZ+aCP50X9u/r+jEVGJHQFvxYe3tePREA4gMtpf6/ZWOyxefzPryypz+
Jaso0SCnUS0pJoH7ku/y9rGGqyUk/I4cFN9lb1ZWm496/VI7VTimZuTxLMJgpTSB6IIUHNlbdQ+y
M91ib3cfUBr21Go+z9JW+kipIyD+et293m58un9qxBFAk9hGlBFwDRnLIO5Dbubi0AOe8zZeKQgU
4gJVoF8CfTczx8wFAvYajLpdk24KfKXxrmIbOfJhnH2CpI0DYyynx/GuVxN+yAb1cX2lQnAr2yWt
ig3zXSYIYQeM0HeBzAS1ZcQysNsqOBmVgShonJEsxym6JOAJdEWPUQHVi5qNElPfRrzmJlrSdiF0
N9xmMxk6Ia2YW44ccQa+sphz8VSFrBf/2Ol2nMoMiFjdI2NhbjGZxMA1Kc1O5Ky0ZHrqNjJq0cK6
COHkMSWPETEJGfzxnH/gedP6C2a3XmCojJTSMrGZVqveUJvi0VgPZMrd0bwHXa71wBgPN6JSjqD0
7slBKClzRc2c1+708ovUIQjEU5fGoD6JVakwMd+FE/IPpCoxOhabtd56UJ7jCenQx7E3qsg5iOyh
lm8+/xh2xDIwHge8xWdh2GYHo7hkkHITddozi7EcxCKGJAwWvBh8OzpPhA2qnisimDkgAhyNDfsU
5yNrVRVtsQrfgMDCD0oTL8S7p2gbBLMi61vCN4K8wgT+dO/Cu0PiumG2V19s3aeDLA5Baxlv6QRg
oaVizZYoYFG3ZJiHL0wVCB4LJxHU2eL1r2glfbtnUnEZZoemdivfrk2g/R7AvbQweH/EbfPs2g5k
35mJH+Oc38PMSqsERiP/QMNsYfH/NfEGpRhHnCAsOWjTWcTUISeEY+VlglgSGFuXvxiwYMWYENzN
cVhjmcr182ZRGf6M1rgqTJzStR6jAKMnATQdG1swKZs8hfJyQwuhV7gd15X8KPzv+K22tJRMQbBz
fX5PbbkIOOQBnjszySITTiO2sIbdttObOpfr6r+QYyWdwHHY5nBgrFiMDuxcokXrCYlis8XlKfcD
uI0O+naW+aETIaWgP7wX5V/Hrn6cW3qlHau38Xue1b0n+D9YCOBqzgOCvIMfuyJKrg+l+z+HyCmP
jf2mXpNxO7izHPisRlSx3rH/nhXOy38/P4cOXaet44m9u2zP4i4KGvOf79gq95f8K/lzf38vZ7RG
sS/NUu1YEEcKznXwCzanvmdL2gzK3tdMd7k+sgA7yIIYgP1oJs+xdg02KVipNh53+/LX3xB4vUMd
QCwJVKj4XriE29MQeHM3CJTq94WJc/PfL7PdUi3rGXfUsqG89kvWy3oTzAR9j8PYBfxDRroeuSbM
aYxl+mOLn4apTPHrszJkFnF0oXcPw+gtTzHExyURc88Lm2iOeOPiES75CGKgKlEqkaBdb2dx1cpg
jJLkME8qDdNQpbmunTcBkHVkPfbxujCoEHHtskfMYAfpAsY//E75pY9rQ1rzSCLVrYLMljxruwh/
UPP/C+SsEAUvR82YRz+mFU9QaYHawZvVE1GU1x3oyGQ7YjTFVbvGrEK3YWSFCMuqFmLWOGZ3IonF
yQtc2/nkWU8MjSn+ZlQMPgBQQOO2Cv2B3MqweIdB2JuSmvPuQ/i6wj2ffZwIkLk+0ALl6lDwik3d
OcKt3DcNXTY4PadA0v5Wj6Xgk6UU7HGlaEImvCC3smC/FF2yfsmj+IXkQipaF8hSnwMYEZRVNpHV
CVVEoMVxa1C5OTmVNBRdnzB+pUL9PTNiiqUvxec2IF6rmG0wagRGl1eC9DpuadsZTrO09Whj02sW
jN5r4E9Z7WNagEgXnkSK2t+1Rk91OPgmxP7/J3R7xjtrNmGXWYjG5eaIn68tKkPKYQ3TH7iEYby5
lnBjmPSmw7lhBF6Rtew7uDyAxYPqoglEq/PwtpB8PXTvJWbnhBBSfTxXKSrgsBHRhfXluhSgTFgr
dDWxARjL6UmZTstjGJfMJHRJ7DlQIaP9X8TyS/qYQsAoNmIIu2RKDObSJ6ZD2m0Zch4ZlV1n/+WR
pNKBVMEsHaeRbdOneszp8lFfyC4ZKj69CF7YJ8Kj4zJ7+RPSK095jPRR5puPmT5aE2bN383PHbsL
Xh3SUkaEtVY1DJ3Vnyn7wMdzDZf3k0kT5Scv1Pyi5p54UpNSfz6eB55hWW9YmoKVe1wzxA8TimUS
nVwCLb17hCIWDwXskZFFD/d13UcZXRROQXd6QI94DEqNMld6vD+6iaAVgppq72AJ9BQIItjeij2G
mjZmCrrTI2XPZY9dl1RW0RSKv+89GGHwCZRyag7yd27LoNj7ebaGQ3f25KmwQ1SdASrVw7HK3m6t
QRtOMM0PN/tzdXoAa0CARc0ou+GOVr7qAR6emkVRbDRetfuIZnSQSf3UoDJjgDsr/sUctkOEDuwL
yG23CcZ/0t/dE9SImYBS3LvKPMsGeYtWHuMGMxnQundijJ/FRa577S3KnzX5JgRRKlc834gzAPVj
/o9zSyC7XV9oCn5Mh+MCbIIwu6gQMv9OArLPfCxA1aD6R43J8iGPMFWvAvqntSFJEusS4VWeZLsO
Cn5ng1HQpXuSwfT9TptPL48WRl+S+Ly8/1Q8nVD/m23nVzmq8h9TEVqOK6HyagGpICo3ZIE9Gpae
hd18D15ji5gCTJvkGmHQo5vQbxnXgBnUHN8/L570sVreVBKftHo80JrxAOF+yfXEiY0WLscmPj6M
fr47Enkk7L2ECIbmh3MycG6mSNIkjdGtBvZ9Yj/6yFNSLRPXhbvv0HCHwgUAudMLtRTJ0rz1QSLc
d7kSmTsnjPxh3FoWN7Ef9Uaf35/IBUCI1u64XfETHb+sDkzX5yvQMZ9lZUxcDpdCObSijDSNfoxI
dEb/b1eBnks0VkM7rp5UdrtnKqJJwcKLKAgmq8kUFHinl6OYG/zLySl4T4muefNc5QsGWZVAkCl/
3XXfOklG4FDDyv0G3wlRUdkGEV648342Kb2Xl+lFOdIElSIaaFDyLI/DFr3Ntm6qx7mOWQayLhZW
6dW05xbhSCgOa6TRm581UBZsDUvzqNMXQ4NrglSnvN4UWoUbIDQrJA8eX5kDp4KrumkNSq9pjfsr
jYmx85ZUv8JD7+DaxC12pCGBz0KfebAViuGTllMsDBQ4FD+fuxOPJjybszYrihG1qXCyCCyFqCLq
Dclrt5q1ji/Q3ecg7yleTC9JGpBrBTa5k5fdWqlPQWO+a2SmhPFpfUzGseJd2PrYoEjOJzc/JxGV
unLEwnzSWqjEXrP+o3yzDasnqKTF6ARUqWIQc2PbCLa9ox4oyBR4vFYorn4udlxI0Tu627dDG2dE
+GrhkD2Z3hav54vL6B28UUrGcluws0b1nDE4ygqWTkXBtt193080jztqz7yn3d5TtYRZgP7aZM+Q
gVSmrLgzFkVuEnN9t8jfe/uylAdOt9fIQCHieOep/z2ZoFJlZgPhSflNqUfsowdPIvw/5ZddJ4OV
irRHQRjxasby44+PGONETtMMNtxh/uUePJGTlMUqe5CvyFXZBR9u3Kck4eMMJQAKRBfxsYp3JgcW
MpQoFYLQSddB/CwyoA69yhgH6nUSE+OjBxZEFUM0fBMPzosvBv896D9TCUW22vAYwOeaJR+1/Zsy
vsq8sGlmqOYH2+AHpUwUdLWWRpF4m4C2pUKYSFywzWCpZbr5rjVS7SRysJZcSkCTkwJuDsc5YT/a
z8ZUa8Crd+Yh+GJ7LacLOOrHKq+iigR+vludP49ld100YC7eh7EmboGghFnckM6Rd5PLdp61UrrD
lsqwCNUUvoB/IJYZ0neH8wk5jb15yNyT8bf9it9ulwWoX7DuaqkEIST1cAVY2lV5Klx/RYyns6dt
TS6tD7MMcnL+1M36QYViSGbiCJlGTMzBIVDARMri3MVaMVuRWiG13oZ+oYd5s7zv1aeVNZ8pawB7
my9ubOEk3bk99vbnfpGFDRdI3+ovlO5eB27qfmk736sOaCiEjd6XqR8Uf7x3SV2kXoUr+4Iosel7
0YW3gUJyuSkiZyDItuLle5WdL+oAgILkFar6MZoV4Bk9BsROHC3eBLF3Nbreshk9ghZ0jYIqtLKx
90VpuvAHJKA4itTd3r1YlNgBlY2qieag3IRmSNJOiNXh2fV+Dgp00LTlv00+LLNNO3Udx9WZWXqr
ZAfagLQAfBQ1rCMr6G5p9Li7BecizpNjODFRahZwMcTzMLRaplzYTc/YSUOPR2ruEkbre3gK/sM0
/NHwyWJWiMqUtojYmB5aefABebiYYOSIq4fdCu6VHX87N0ng8oH7WkcH8WTyoz+bUznSkYdMzwqg
AYxYnG0pL0sN2l4JSJlLpzyuv49aqJXCsFHvhCn+dN8UNHPhUdkBq9surRIK4YFy2B1bFsUwshJd
BY2lhFmATZrmC0kGDUuLS6JSvMw0rTv3va283eCRFGPPJdtQlR+tmmfU2sS/Lg2fVxR9rELpcBbA
gPsvWNvUNaVQzkB5io4Ma7UxQhAsyQgAR8793urjujB6YPgzgjlx00Gk/iIHIi1CwIZtY28rJEPK
/Pox2Tr324d64z9nCBqjRfgiYHOZzM07zcNyJF3WU07nxP91gJZp+f0/MfuC69ylXwQr0u1YK6lE
rBiMrnNSQwpSPOtUVC4PQ/TprRLwjlYs8hwIH94ogJdujjFZXMArBnha3y+/8cztwbxq/bCMwxIt
WcerCFj2hzDWVF5xkco5DqKiN8RQ0vuYoB48kGZvTyFmIZexRHpQZLGLiEXTOjVOJLjBm1nodh9L
swsw62k/jTOqXbMMrXcsmghgd2jGZJOsGhGj5xSiLEHbc1waO6rwrwztFIpJu4fG4fIckJFHZDjb
SGpHQ1BrUplYusHKZy07h1s4plf7ITaOV4mWMEDnLQkkyIAxSzXwUFvsyGDRp7XTWTj4R8x2wBnM
/H1IMz6S5azvKZrwD9H9s9+L0+M/gA/j3zSZC5uDapHTq/nhnJyi7xXi6vBe7ITiZJC18ijfS9Mt
LsBehGE4wXa/9C+Jatklw6Qqyl2enpjmnJ4hry0eAyrEL4ejetUSqpRb4yKB3BWDx/+zFy5tb6Sc
tIIUdOG7PzfRqAu3UN37fnY/M1pBek1oy7FVAw5CROm8err+DkHPcAXsxtFLT5wpcCeCfHn0nSNn
Jnv3K/2lYAazS07rHCktHn2POME1j+f/BSXTyhZV9BzkwD8Nhh0OnyVy6ZL9MMmdxIreHifQuj57
KMCj/Bt3Sfn19XwknG1bQ4IZr0N7E3JAiXSLNa1cfJrqSyn7gsbcb+gzbBar06/FAN3AZT29ap4Q
xecGXlxBaShEMCtyOSy5fghBuRWwj5TZwwAoSwL+iVCiVfbU43GkvENn1Ao4HxqW/z6YBYPvaoAN
6xhtyxphB0dM10jfmWaPtM1qd76PrzOHeCioxTuONA8a4l4AQ7ZdalvPQogF5RAqc9K6ZPkO6OrI
perzh7J2jOiHccFVGX+YyG/HDEzjrQeRH5jeJiQh63XKy7owrRWXiibz4s9Zo0oH6Oho/Q2baKvd
9Z/a+V5ewiizNtQTan9zNOx2TKE4ImJxsVnCp9EaNJcHoNYdv5K9rgyqIBhvNj7Mxm1xDskFdhrM
VJcm05/ZfHRvq8qinfWULPzDQ7hyyBBKbMybNJq3JsCOpr4YAyUJWdK+PdcLC79Bl/i8ScT7y94M
wLePddgndBC47sNalk3RKjDIUQXDfMLajcOM9xpK4b/dIFjM5Qpl8UiJg03kLowid86+Rwrq/P5q
VNFOWl96rXTUnAkOfuaJeB4Djz4+4B57SlYv0fSMIfc5gccOxJalAWTfCBH1CRi02U3ZULxLofOt
lKh3hn0PLzP0+nbdZbvmlAxlNSN2dmbLcw9tWzSvQvZ7Rw7lp4f1MRQNG9iMKe+MiUSEjfIosToj
n98iPMRWo7kL2UwhRFR42TcvpPuVkQyrUAfGOTPM1dtWGpASHDQVlsDPTZnbEmvmUxdGfB3IFtiL
yu/6MilbjGDlXR0inRD4Bbb7N8stP4WvglA4+pOR3uRz00BTZjX/nWLAmjCE04WfMTcDiFICEv/j
dnvJXYI7TzQMv1N7baxiLVdiS5J7vM1CCYGxSaTsloFRXltFXvSeWdW/xRuFX4x0w0XHnTx7imY+
SR4UgeK1nsTfMhcLi/Ciwt8jw0Hb4EOCH86QmSdUJZZ1L8UvDLyI/UfYtcQBV8TNGJuQnhPbExiV
8+wjgELJjqbEIXA63jTtyn7bn3UihPt0wiu3m7oQBDyW8CwHBbILpeBf0KHLhBdxeXalPKuKAJm2
i34aRsmfTK9P+3PlINULIORUhtk9NG2fllx3fRrqhKSM4bvwFQZORFztNvAu1FeI9Fe8rNrsLlw3
X4t0mcdfMyV/AgEuPI+mj0gkZqcbhJjKmc+pq0at6HviECWwwyEsfXeOihhG3zxdrdxtK8Grzf0h
fz13eqnczGMuIOl6+O8oHQvzadXwlTtd+GjfzcMkVOWRhjNF5d3Jp0CK2okblyZJlNil4bhlJ7yN
Pn5OR8+UFaVNCuxABWzBR+BE6EOMxGygGMhEvmVk7S7XoGbDgtFZqEG9Ps1IvnOc9iONOj+Njb5O
bjByu4vQ1SMzkq2ILqFVZcmuBXLzLTHWMDaR017KBFBleXMkrOlrsq4ZXLWDMFQ1MpDr4VxBf5n9
fa7p4ZHJ4pyN+uXWh/iCQih7I24Ii+xSKCSFdAFJdmr5vrNTqD9Cxr934VZD/PuhhBmN4YG30vfZ
aocGLDmvbh+lFIsBGM8tU+raQfCwD7A0l7DAqB9gT+cksPV8dF2XD71KdSNQd8XQ24kNCTiG7KQC
5zKFKopQqMdj+ee/9yoqb3j7lBpL87gf+5ws6kzh6VOBmHUFTlaZOobhJu72RbV0PfEtXJ+oi/Df
H8bqmunfxM5qWyMMNfYAhdJL7mSqFxzSNOhLKYwfNeiOaTvEZhhcgVnsVvyWI6cng6b441OpzklS
hILWrNz/R4/RUQMmowAxOZtV5FKzfIXSkC0CKmGNyupruysM6F+d92KEzJznOPicwpH1FvF8DcbQ
v4Z3tv7vor2udBeB9keJlsNhYWxC2Thbe4xlL5eUD+T4EXY5ae0tU8Bv0RhT5DrsQGd/ibFUnvS3
QCRDQucy5fi2J0TS1lg698sC08V8edWHlzQuzHznIxytUwPrLqmNGxAweafRsmXW6y0dOSQkDfTl
t4WkACoadfFFkjqNG4S9D6GSl2WO6c1q3AutlNJPwUt5pGk/rpvB1uDnJ2XHQ3KOfDBXYWTNGwCJ
TLrMDYUptO5xtuVgA4RzeiLyqmqVzYVVdOjMQo20z9z+FHn3wW/F+NpV51Iru3J9l3xFM+kF6qcU
8H0ZE75yePcou799SAlqJDRJhXVsGrlpm+vaV+C9aJIaxrJvpIaYIsHAhnvirE72z2XPz7DFzBSU
e8RlOLX4dXmN0+j1Tr590CbnfTcL/0UFDcpjyVHfpsZf2JhORWcT+f7yFFk0ywFZVI5UsMJlRBDG
ZkKBP9Ss3ilmtA1yhw6W5m8BVg79LMIWPXD99ZFWAP7Ypas0MDSDLYQhj5EHm9eyFocLFflpDvjQ
zLh87riAKtdJEQOmw3TsAEc2T4lv3emJFw8iH0qwk3pI6C1NBmzlt3W2N7ezypjv21xeSHxnvD7i
FPyKu5Kk+CXg/nC9KtZt0pYSaLmm6Ka/d04WmDBYBnGTTD6b/VtGwaSrZPbwlYdq+qRKvaYLNH1h
0MscZqiHiAnc9YiI80jWUTCyR8bYUCEm3ZwYw/b+cCL3W4fZbusSlsJuISMz9ekhP0kctIPE18Sh
K2CioTQGv6uJW8y9L4g40I8meU2zRsdXmVZIfXLRTrIoYQgaAikmxZbCXj+61z8LnJ+uAeRMNB2I
nhAR/4ge103+yLN+/ZUGUHm/3tbqUWTQ3bE8MlDXfZayJvUW47f5pHrUqYRtnEYkPotNfTIbDaIM
Wjet61WTW/fFUQhDSVnSc+Cis0ra0Pfts3PuCgYmIP0/LCIL3P36n5gPYGImhq5QOBMxaWAfJcNL
lXi4Blvw9GQ/m6M+wxVEb5dMVnKQEPbVS1yg2N1K5zK+7UjLMAyxGN17csd5JxB8NNxxsW58/G1e
HnfvLo9ZOdybDsv3oRBGz0rsLKasfVONNJBY63LrLGTJnsrSngG7uaUaYvrRfREdIXUQ3JolBqSy
AVVl4T0bdI90ks27WaNOKOH2pHnsY/SxZ7QL0W0tib/FhoVIYc5juG6dsncy5RTfYNrV5oeClnbT
60otSJEiGcs02Z5rZZmcoWM+HxAjVcWYGbKRrSmlGDe09Negg3d4/I0j0vyRb3h9Big1xBUVu9mX
iH6xMXd+UQRZD/GJBrEUtbK+fHTx+5D3nP0WiG7PnSvI/rflqcMTvc5sSLnntDeTlqq250ib0POy
PFrb8ge0ToF06GnOy6fnRtdZdswH4WtKujSRxkDIMX+M+ktgdoWS7SN8e9jGigbsSzHyXV+TGh8j
RFmqmBLQTfbSzqoSE07iZ6BXONuslHKoz910uAM69DtM51iMjO7cVgezIihNKlRfDx/aGXsmuyAO
U0rULb2bqxGfNgYkznFXqJQQEstzb/JW2eM/94drGNnQmjdZYz+y3Gve7wXP/uXfYtpOcSn1Dg3a
30tZW5Ds97xPhRnXtYfBrKwgfuYNpg5XmQSpf0L/LFFV72mWLHnwLZVY6m0vyIfh3XhH4oF9yFiG
OT9zWXcHaMApSx8YsgVmhYm9in0WkgLi2GS/WtCe+64gHpXWiM106YgEHsnK1cR++idVHnSlEhec
KK8+a664FjK5J3SbM24Tq0mXyjTboO9AdXXvLrC4coaev6e/P+GHFbL1ffOhBfJRg+pnMSre+R7z
uGGEeHwfTqEqkF6xukPN0L2vY1njwOBvRZ3fk0d2KzeXoKjjToCz2M5eiW966J+38P7ZUWGKDsT+
dEMZjRDqFZBl09aaSE2bIA0zGgwFJETlBH6CVF23OaWNHyhqOVGAfM8iaEYzbyHR6RAr8eU3pMiD
TmYRe3mSzrBnaux3FMedzJWSLrN2sULKtDj2QyJgtRFRsihhQqrHKHZo/yyG09GOtDYHpeOZBhHJ
eM5QWi37A0979sTOdA69tHLAYDQqUZrttqjHtL8rR/+rjVzQMm9qRryGvxcD6cI+xavu/3PXlTv2
3ZeQa6EjMF8se8fjXzV/F3ow4fHxvPW+hviyxp7qKvX414dbGyAIrMJd/YPllL3iBf302g/PZGMO
f7JsYNflt9JKPztcFuN/IXjQN+/kjfSDp6wByo+xKUHdPzn8VvtpW0uiyiUWENVge76Vud13FOdC
w4FXcpyjUNw0U4ucVB6OkxdLvjE5ONbvnTSnaIMdXle/nvC9qYAjIhyDDJiqkSq2lAGYp+jglZtL
VhcmyrCcVV+Tdx5P4sbv8svNUrHvxvq2mvUKwpLpFbjc8u0gCbbfOYgPmX4Evwmg1fhMxm2u1QCX
BgKsNY4K6fVSX+dbNzvJXHE+WrpsEaE7rF+DJ5DqE/H2bC/NPAXqzLAXHN4p2ovQeSw7qIT8r1vC
dzF8cFN6cCe0qlCSSv9WIhYSZaI629VKBlD/s9MwMN/rtAWbGP8NC+DAqHA+zhIMgRVPxBVoGWV4
b1gkB+xP6OzKQIaVxCj2xfTB9hiwytzLsCK9RCfDtYbyThASegLZJSTBvOUpg6m64x5Orm3Au/Ch
ffoGpNobq5WQztCD/nc11jYqpuqB/uded9RrMEZ3MTEfGJnsMzvRj0ju8xchN3vBTrY3/eAiblsH
2EwOA77WROqCRa48NfdgRVfqF10ZSSg9nZuyWUW9ohouAQOjbWmFEM+0tOwM+ZXoydTam81hvgcm
6l823vv2a8+s1yFJScP8h7PxkQix3Zd0ADZcbzNgWz8H5bmfdV3FCg45kUUsV2+WYT3FQfjWUWQy
GpAzLEkpsBwftEXNVeQCeEy/mmtbORR8z3KI1favFEHSYmd5xnbT76v9kMcxaQA+y4IDzKXXYs8b
kT/sgDvgOY37kS2hkc/jKuS5Rdf5cYQfCXA6j1CniDoY/c/HA1YowW+fbP1VjG3L6E64zQ0Jcf/q
sLf18vYpuP81hGmPEIUQngVIT6PI9vafAXCCbWyb+0xzu2+lEi5P6zjH3nxpufD5NeGqPBjCWYZ+
jQpVBx80+2yLe76+7Hr+986ogLo3XZyaPXDjP7HMm6DadqR4J4MaCNu5PwRNGDTx8dkAi8ymYOGa
ZG7UxQSMh2KH53WNsw9hl2uvkmS1co4RwDRyHqbuc0xvmsTPShBgVer2Qf2+ABQJNUjwVOZ8z7oN
C1fsdnI9dtLQPQb0kK79ChsVTEOZ9RBvIE/ek8VC3RZVi7OZ4T96/QwAvpv73I6ihrvFXGTqUcsY
yVqMA3Ke0qf6Eb9hA20K8u9+sy0OI1Qh+SbyUm2QIwjaD4vf6cSy6IczFYPB49TTOHeGWQGgF6GO
E1DF3gpI5rFitHTLfv7nLklSuqLTxsi0LRNIQ0sVrdtEL26iIQII9L4QmBiK6xCXi1u8OFhs/MOY
PQxVxVbjYDtrB94Blon6HYdh/8dla+zO5xUlTE4T5YVlcAICAB2n02BhlScn6wdwgvZYCb0RHUjT
yEVg3vBUG7eXXImWQiRQV3kbzpUvI/1lVlcZfWW3tyG6X6vdm6BavBD0kY/3Xajp0aR8rcqzi8yV
LMV/C54caBFvgwVgBkbIq08Xh4aWI/ayXzs1r/z/3LI+TPIKp+p6zns7gn1Mt/YI0XQj8mlLzgTa
leSyDfutBB7jipEDusEEG66IT/2tgREBxy0ZBzvf3xXv7ZFSJLJJLBj93nFof8CAmb+8AWvumOat
BRYFkmT7Qq9zV1DohqMdwRxHiA0ru3mi5N06p40KC/GMsCtii6kYVI1X2/Lx0VRM5ulxrECHosGw
fQNoAST0N4mFRo4mX28KaZQpiLlFzBnhnzZZO/eZ30dRlOrnPiQUBfkwTtXf3KeaulJUdRgh0Cm5
AtDjQX0H23iGyI5dX/IIIy2BYC8f3dg16O62dz0NMNxLXcMJnJ5FXk7YRjYROwNXliK7i5CiCWo5
K0crgJ1QftdSTa+9oqGrskcSasjRXuOjk3+4mYLTzCvaok0WYPf76gkruIftmL1Mhf/k+rOzK8tQ
ej7atxYAv2uBJU+xXqLW+EN3LpHJU40Y7bTnf294smAxFEYpekFr1bG80InBLoMqIdKRyc/tf5jK
LhotyG/x9w/4A4WOImYBJzhJQsJSfkFKCQRevaESOs9NEiAynUUk3phhsDHt9v6LN5+1JHuKToS/
Rka+7Sm63FqNjOlXb8ZJ5Bzk8EHY7VrTo2h/mebishjSEW2eRMKIL2o6QfPg7SnDtT+MhXmjVZVA
QMn1J7o0PITi+LzkVYYTiF5WKsEs7HsN1UqoIyZBZVu3I7U/NOSPFnwAlqH4+9KAiR/0Dw8ybDoo
ysWg0T4WS0s9N/8+dnz50c7tk8dPlLTNzCjKkjj8nCwmrRNSXg44xPNk/Sf0be1kYD7vb/eq9+yq
yhvKZAo53Hl7fnVygMWfcR2oGld4Z6FGJRIhvnKvSTCw7Mg+WNRAS4lKIdk/v1OWmC1IJea31QNm
Hm9zoZ6IpllpTo+fHdKtMuENE+xfb1isBtmiqwBLKMwli4P/2cOUdmdznV42xa6/XupbA/6PEN/U
nkt0rSAJlO2QvsSl9sYjtmjfJmstpOTRA0hfL9YBhJzafHgPcxvFieJ50s+omDVM0gslsaDoNzXz
Zjh/Z1OY3371YcnssD0N//1CGCIJD+iLGPTJgABefoPoO822GEAEccUi5c+wSf7DXZJu+z619bZd
5+mB0x1wEeh11jCVW2kvl+eWYrP0NYwt+bh4PlT0ZUkxOTgn5b6slbkuf7NYvgczNsE16ZoFR8F3
dlDJpHIipRaECRis8Pl26Yo98XQXmEo/MgjfRo/oHxfgFRle+77Z7OHZuR3NNgkjoTyWSd0OgPCw
Wsfq4L5OPfQBIGRtCeYXfvFKUUbY2tuc4ado0+cRIrfdC2VCvpD4V03Mjw46IgdZZj7LekN5C85e
k2j9/+nLwPX/misTEZ9XLtOEUManyF2a83GVGma3gCNbqNkQynhu1kcdACBCSqQKTh05bROYWNb7
sLUeJ9jMHN0vxh505srTQhfjf6ywb1HIldEwjRZJZlYFJPPD5d9ljdReSFIvSW9X46bcBBh8YiKS
DDr6ldpOXoBDZR5rv7QI1WdlaftRMUkGe5Osoj4qaJvCtsF8B1B/ofq2avNn1EJKxojBgd0GJkFj
RcbDuJpDG+lL/nsqJv0j089F6z2U7Q/kU2AzHhI6oqHhx6S+A2opmrgdWRtcGKKFB7s4lS+Xg+mw
yX0JkqmUXkd8gXobT5A61GxxyAudyipjCCVcT5LNEervuuUM2Zh7t58hW1QRxhJWGbJOmhJhb2C8
ZZwBdZkM1fIwnW5Zc4ptMiLBGnqCuAs1WGVaFuBCKW/IXBggcEytFqsI6TxfSmtSNwv2yVzDzXuV
q3MjkISRDU/EAJl54920Av0YKO+eVurWJVzAE40+2OVxTPm1h/HjvGQFf0/uTZYEvFvOBstwnoRW
bYiJMnMXPHln9pgmQQBfdo7l1tXYFKflXfcl2PYr+e9/Vd7wgw7p4zvXAHW6Tr3oEJzxaMh0XrVk
hyqhFC3s+SdKUIn24/aSJ0ZVzvvh97+J6XnUYjSpNePcr/7OYxCjk+SB9+gOwlbZTz2+b4+QJLV3
fuy2OpWgjoruFuAxuvFJ0j/6thuM4Z4TpwfPeupzEl6E+jDTZH1VkGq4ZMiQ2cpOj4K2iRLAMcZA
GMODRsAOX9BCL4B+qMHXxhcV+st1I+GcgrgV4nLhWFpy6aBtHf3+Cs3ARNfHmHI8X3Woc1468N2b
2SSYzKPUvtInqd7eSTsoDZCjqL6i5mZd0I1znIiwHd82QrruyNDTvK0eu0CfcwYArahK5/ocaxq0
kfCqVmJ79UcHKdbBYqeny+vVp4CveqO42TCNjBw+bLg4ENzlmQkSWJkuREjT9fSTVmIzqUgN/xC7
hS0fER4EqqP5uSolaKX8utDrPFtU5nLFCy8Rg7qWqrOD6xrqDwSHJjtXGpITZQCGYvjjXKGVlRpt
9GuIUKhe9FoMzU4Qlg4hrTX7gHfl2xVbdBYmI9GGkexRYwXTIN1Gf9iPOCdKfVz8NUpsfI8MerFN
UV//jVBxF8CTp0bgO+D0xHuEJQM00FNeGCBspwoj8szCTs3ZmPeP1Ovc4eKLqvalzXJUsK9ku/oN
o/WDtyqiPG5joet6GNj41miYH404AUjeeGjD7dH2wFlzolvokHp/pU4k/3zTbeW+YmO9UdmRH5+D
u9Hf8IhB7UNgR26NHKGD1W0DuWdzZYgNqd2FW4cPuqHJ/9YTLd5+iqSQ6ZsM3vgUGxgLCwIvm/xX
Pdt3XlmolocWZuC0bysbyT9vGmKBJgfMkVrEE9JMBoM3UKehQRFhMCJxn4CNnaZ10cqwKfy/dhjt
YnBQ2Fd7OMk73r4xTG1hbh5qxLSRF+cBXZpdiEAnrW8caI0qEXOvOG03nfhq9zzrI3e6wdW3P2Q0
CRXVvk/9FhwswLpFDkc1zBdKL+LIRTtAvSP3bKsre0wzkw2fGEQXAkRUfgaTwtMlm0e4l6g7Ukw9
4Js3JRZkbIK3LSlrAwtrM9WDKnARek/OobGvk/HtrClfpIOCjrOD4ic41OuJwp19d7rm6PVA8IeQ
K/T/38NoWAJ3RdVcKUS4aBf2FekH3WT0TfNWLhxeunTyig4fIbPxw+2qf+9x43XxZbvP0XJWyg/u
S21VYDyCbzhFyG2AQuxNCDzAknFTB7QNZx5fmmNmipIyTE3WxaurcykJdrB/LwUhVaGYHwbFkHCD
QZdTWV2XUPm3crHXK/G/YcgYtQ44OmpiwKGbcj+MWA9Qs4r6eiZ0K6GKKPGx6fmZEi9XkNSsNUx0
Ga8w6osHoSteUWMY4IIVY9/IiyqJc82uXHW5ZraKYJ1ME6F+W7KwIladFQUpfkcIbWB60KK9fB9W
31lf10wzyh1UvAiid3IKLiZtb/PynKCDvrVr1/X81IZimluSgC0nYld2AMf0kjCPjGA0Xbpnd3kh
mvzoEDUxZ4MCHEAN4/jaGrGIfzZVZw0n0sOHoS281xq9+pLh5uJLn3C9QqkHSekB2A2hKMrdoH8f
hQ5GROYsihVje+kpiMF9gqdNyaI8TGc9d1fLDSf4C3IXWSxfPsqOG94K1qYjR3A690o1NTUaTyf5
DN6Fkt9ViA/w9aPek5x0/jAP3FatBou3Htbz9kMVzbqh/4VLh2jWohY9weSWXvGtSt2cDYlOQPbv
QhlU13T5RR3sEMM6mCLhYURdvjLNLevhF5TwKJsDpAtu7HR0bK1Utq5RklRHau5oy+JYr+nQ3MyG
X+s4plyUxO5SFz1k0WRUFGDp7MTh8FghMeqOL0GfLuOFNc8D1czcyDBmjfolCBxkbCM7KIin/ffo
2os3yrEleDC0Qc91Q4dWNs5PVK36T4KEZ1PTICCwU0ols1tGtrTJd+jT/I1/U07T4/FMPv7OEedR
8gDvABKvLfCQwvx0G2upOSIrTO58Iw9TPC0MOitmDhzApmU2lRVqf6T7YiGrf7mujxCFmgEnYGRS
AgcVPKH2TU5BsI647Yl34n1I8mWdQbZQeEOmKiWymyuij0TeyQEvabXpj1us7hO5RFmm0O76Bdz9
hiYOOR4miZ85E9ZzhSMzS8v07kyOnYSEBulZooclKxJyClKcSGI+M6R7CrfstnV1C+h+DdRlWSwZ
lZUC/tRkioXJ3RUJMR+wamrnpIaXQ2oY80BC5CbIRlQWyZjlUtVtrqG9Qf47ptbSnQVCnegWdv7L
E1Jkf9a0KWsTH/kY3cOpJFfadQ20ChnYHRAZ91VuQVw8aVrPv31Tf49GtKHaSjgGU2dYS2kifvfx
3stIVsTvV+P9+84bWXnPU1AuzBv2gd/YMgS9RWqXrGJyH172VsxGX9SaVMmRz/w6Hh2qPEKwSsev
YR27VMnPPc5VKJXA5opDSTuEI2Zycpm0NYgYyCGMlAQ36Zl6Dv9nvUlj+ZK2drIgAl6LnwzgBW6W
VQH2GAgi6O/A6XOM4zZP4RchNdZcHCwLMFFLTBrDu3/4g3ThVxabodDarzKZFZs92o33eS2bP5PT
WjK7KvuW9VBmcKhCdyl+nN2JslpNAI6y3TB+605wzOaFezzjpMnFxTluP5L4W79PIWRALhRKINn/
JAEZ4jU4NfEHywyOUoAEF63xUB6/jxZfNaibH6Ji5nJWpEOXdwWVVMqP2vgZu6t40gnHTeP4aOI+
hBWRZp/wkj0eWfqmYhcazUxTkjszGlxkbJZ9pUKwMRHMFcx02Qm83/g2LNZHXIyBO4k/YK4Wswzo
wzYGiJuctBgu4xAaHIigvQEUIgT5cV1qrF4edozFfh4qQehR13oqgaagcNifAegyZwyXL/ed1dtQ
QDxXsMSMofSKfwXJDcYIa+Db4T4L40o/XLjSZwp8xtHO7uyw5dhq8FQuzTc2ZqUMOJ0ASuQp1EEG
L8PPBktoP2Hw2+HJpHIhauwZ8s64WdjPdjX0Px2aQoN1BpECRRZ17Be8HBjgCcHYEjTQB4rXmNPm
5OAYtYGqcsYmPOkaxhEpPN9qFaTyhuDx/4ya8lNrYXCyFevFe60xUrTiTzkjmot34QqHnvckibE6
m9OvS/V5GO5q8ExCAP5qjVD5Vxqiq37iwpe5Qhl/UzBkTNVySn/A1jWhSm9jBm3BKcDSwrTKyW7H
dTlyDAbMv6TlVV3/Ru7vT0h9iyoKr+m60SdIK6KfXyWy/Eh9Dg9lZGC272hOCT6EbCiBwjCV2sFJ
L8bOMbijFo8quJgVwQliQQY1NwkiP+VvcK2Ns4Gm3SLxMNf8YXVixrXYJIjSdjpDd0IBu/GBTVN+
livXdSaqCOYkgLfTO3GMshBIVOy1IG261KPDQXYN1lxnyLzvDmx6rgulk8FvWmxOuhLIOEJGzFeq
/DpLXT5NYJr4fdl1zAaAOw33/AZm+r1vP9Sq4uRDd+N8Gp8DOTlu/rX8nVBs65U1AQB4kUmTxBkg
px3J4DnSdiJbQVt347PXhgVTSj+IIJ7/ErNgIM8nHUrqUd1qX/Z3J7h/Ddu7xQ9PZ2Qag9ek84Lp
ZZEbYbvIDIXp+ML/ypJ2p22iWYzqVe5dJONvsKZ7eCkyZc0vQdZyh44C4fkXzAmon/msjk75/EC6
JdHvNZoT8VWb2NXpUVAMat3D9VyguU5DYqsVHZzlRJ7IDy+jL2fUSACYP0/oKJqGJcBzj3InEApV
QA6A40Z4Fy6V0zvxlZ612XHFRBDDWWje9DV3C2DUQA/NP3w6SfMgWN4MtxTVNJgGeej+wRiWtfh9
kzYrjDdc32QNSURYUxtR2uozskfC4MOaNHRaa6NIJxt5bGSqL00NzcqCDU4z/gdm5E5VfzeT9SH6
jN4yfxCyRb/VxeW7BecCjbFuUqvOYJ1/Kv1GWZRusgj+YoDRg56HASXasAjdC7Pj2hR6bikHQeSs
zzsOq6OAuh/Btq9uHNBm622ZOMvP1khFs/RQ+qzWR4ps5QxTt+iPEXZtdIokQ8VIAblbxQctICyw
wQz8eMYlhKlWnfpmh8in3DDIGG7Pf/dIbGKeD1x1VrFgy1eASQtAFiUFlF+G9NukrbtuWdpVXMrl
KCcsHiT2oi8+1C8MCCuHYHly6gw5Wq7t/FRUbekKTnIA6a7K4PpoVcb58KeaF69PKwPP5WdAl/1B
syvlY8h96SkpdsB4P77qM3a7+imGvC/6uYPYg03/haMFu8EccwuvLQDGmgTNPHS5AknbyiFucoiK
FrL/765muIvmr3FCVvO6BoORm5Jin888R8SAZBmdVzkz9sH7bUQCzGQaodrnp2vkFO0nUci9o89T
ZFbGNZzlU7oc7k+fi/76yCL2NHzMr+bTZpyI0jd9R4v5DqC7sPgb8mMEy0FVDoTAfiDuvkp8VYCB
Bd6j2Bm4bRDBTxhD8FLBbug5pjrBESFGsCEjKO4F6hUxOEwoRU0kPL8n7c40/BrzPhk6oPLjuIdW
HNoXWIsMA5i7ux5R7T15CLnMHFDa106Qa4fPSRWYgiQc5paLIM2qd6ltSX2NH82R0rx483nGf8X6
EIv5S1uah3LekQQH5KEEVZLv4CXADKHLkd9sGS5bWpxsHEjb1LvEOKV6x7X+eWQfQ7pGFin3Ujvn
xJ7+X6g3hRSn5hMKxHXwtb6GJ/9BCM5RmFf2aUh4htQKjZc+/99gkcWKWUO1PMcm0ld8MDLzwyqT
FJdg7ZZ9+w9Rqhmpx5NthAs6OceSV4mLyZPqZTz+TvkQyeEprRggkMJHkrkDQzBWyhlauHu78If0
Uqdv/QzmpF0S1yxxF3d9WFjMGCez08pm3vklk4tqRLms1ad+MLkdS+JOhYfut2iY4PNxTXG6kC6c
96BNDnqAkw8ltbbu60+JkUp6Pwzb4Ex3F8JF5g//btdRp+SFOk0uhIDG3kOD2aGkqFsdVpp3ce2v
xwwZ/MvgkYYwbkUeaA2pz6W8HB6S8kWTu9yaUi7eDsysmOKE8uRE7otLG5DFAMmVCfT/FlHpTdNj
8FRN2aPPWeIPLdXK0XTUInxW7zdjGLhWCWTfzQ5fI16FQ0VPkhwSmTWzd/VhHkDABGp5TEW0jIB9
ZGXsezx4s018f47mx1rsx6Ana10i/CIfAfaDMdMhiDiMEqsU15fFUzgbm1VWPAnpjtkiV+FbnSi9
8bu+L5DRdapiVv/h2iDd10tRK/41LdkNeIrCk2sqTYU5czCj6ghXEzNv58O6ktIxRWULYjvKmTFH
I9mxfCAyNsZF3BtxU8lzePlJeaincrpSSu5m0yIrFHin52W5JdRhgQQrX4YHMfmnyrVA7IObE1eg
nfPxV7EKn3pJG1oYmN5ObtNhyzzzsSF7o9TgmSd7Zmu3pseYiW+2b2Dsi68MIBQVcL9KJourIqNy
gpA40/o/lqr+cZcGn8ZYDzivlkpTwAqNqy94WdEP/iaOKUW1IK6PXbOSW8o+Wk2X7fa5K81xjTAc
NLjbPbeQzfy1HgWR42zepFiTEnz//gUnrAfeYMpGH1stqKNwreYPgWJvXz8teo5BBlQqv6ebAOQ/
BQVhUoUBA8tOe0MmkmWlgve3qy56VLgqzhkQ6lq/9VSD/b7yTPjXynKYc64wZItT4ixdw6X/VEpT
VIxKNb2svE33S/OXwWDXXfsv1a26gwLXZ5AdoUVyQRQPC1tStRSAE2odMHZkYyyPlkF5Z4i1BykY
k8/gt3lpDL4rUxVAMQikPsttuTS/vK/4kCsCfL6vKYh4k56MxLz+o9qmR60pNSlD8GYBH4V0eUHb
1q1m7SkN6NO1GleWbDAk6hLP1P6galXlKjQu+8CTfomks7Pwds6Mm/VTq5UvBL4ViJddH1v7cmF4
LStEhGkM1dWDdqb0gzcCMr5vw3Kqfyrl4jCFDPcvB3/GG9f1EqiSUwahLMwwSBG/7wi2lsht1KyA
1TPcIS5rqLilIZK1RRlr0qmmcWGjbjlSFWmlDLzWmSKOwyTWUtgXbAYGpLmpYxH0u9IdEj3m6xXN
6dSua6iMKLA6E52HdolwTCxvsVPFIQ7lp24Urj1SI/4ciqHdcIaor8e9IK1Q6f+O2Qp9ONGLCgzY
ZWSVL0cviL3ab2Qz1bvJlbyFSQHl+f2+w9v5t0dAFL5VJ+U+fpRfiFm256pDtFrui7HgQJolP5Yj
W2BpG9Ek3Sn1mOiDPizK8A5XW9pAoc5H0IbU0PGnHIGKN/nhbocZLNjtZvB9K/uI7xM9b2pn5UuM
kX81igSqV8RQmmiEb5taXtLFKierohC5Zyx5aQBz4V7aK+qYhomZoozc2zTQT8I6AFhQT6l9LU5R
IJsCSYTnodkVLjeYBpQ77EWXcFPrb2+6u6Sa8+YWCFgle/Vme5qnbVF3YzdTWrDCaki1EL86zah/
cYdW2bPGBq3id0nhqvAXF0049WPyqtdwsi3qlACVJZtDS582l4OVekfDTQAA9YrNnIRPZafdDBa4
LlyqdlaVEBrzqtlp49OiDlN1U83tvp70NEae8y1xIU9NbbuzpnudECFFiGuXztv71ufmN4ThMjDR
+fedbyvuehowedAT//zDSb60FPDfZouhfGQPPNmTQu2P8W1mVaRUj28zp10PKXgJrY0PJxLBmuzW
1AA4q+2DSakfZKPc3Q+y0JAhB208+133rUeRLv5wpia+ld/FOzW/R9WUN4E5FKoh+YFQ5IBfiqBK
SlgzULCvvhkelJNMgcgm1BAuFzHbJb8MYJYU6eLUO2A35NMs7j5986COkN5WKm/qa3sWEzywFT4R
ZUZEbMRtsUlTqQcZ8ABbcDdPZK8MxVeksbonEDSosHY30xC3VremIVaUOpu0hqdQwoybWCYoiXre
aeCaRbTOTmI4namkGWdou76AECXLf810/3I/Z9FEpaGxK66l9vnBaKVnmbFoeKGqb877cO7NHgxU
sHWdgkkIW+6Mnhdc7La+LSBgoyxO0wa0Z9w9sbivI2pQU8p1qZgWHeq5aurtHhT/5nWstd3FaF4Z
e4GZAPhUD45R+jmnConX5VOdYq/oezjTexyLxF3NabWv9FSryTEmg7PunY5g5xqmEQdGRh2BYtGZ
CVRG/zw+jKdFf0vfKtvqPcA3B8GTqY+4ZvLlhtAudV0D1HqGbTqlNdwgE7JFSwib33eKNpqnhEka
T9/bQoonABlJk2ZhiI5eRrEOZuJs0b6oX2n445MUszS0Vl/EtCnKWU7cofu9ucZX45QJprKtV7r6
Uwun+MA3/8rqgw2V7Cxaq7luQTiNiMwlWgURFdw+SBgc747/M6FvrLJO4EGioAIiBxi58HWoC+4d
Q47BH6dXPzQAeJoKdllb/7WjDFhFQu+9UbWprLID1WkYa7J9NwkyacA3t5tGOtYC1kRS5HNTHk8e
oN0ptZwMFBQSxuDgn3e+A7WWKCl4+DV+J0Hh3rZumZ45asPxPaT4XZVWuW1KJ9VYGL3KR87+6I6F
/UcuZPiINsBbxBJTKsTIfL7xCluMa1sricDPyI6Ou9GxvVNTHK2WrGz7j9kL2rr1xUSkWhXDTFS4
LZ6TcKQzLM9qzSGVeKhBlTOF59QATKFQDhMJLMQSpPQXSSSxAgkxZmIdKgZfx9u/JNAuaObUT4/3
4m8pRD2YFrTkxRlGGbfoJFk0PvNmtkTrrVTItBAKbnuMyUlrLAEwvYqhhO19jlehqpp4XnRxyefL
5zeFux/xRmCUZy8998GrFSSIufvhWgIHnkJRFGJwBinDxY08GIj7y8S80DnLqT3bymbzLGwPtZPQ
0pfhWKw2KaYVW/Z8fncSZ9oX0s+4+t4ngKHxVJ/+RHct0E5bDAJGc0vexeqiirQr5UaavYAfa5oQ
ctMIBd7Fa6wfwlnOzY9BYIUyH+BQ0LmVpelXvaR+IQAk3icL7hxxPEtnLoRtM0yEWRPPV3apXqM2
WiMqN3kdsm6K41YyMAEuphXtTp/QWyDyg+FHm/lGd2Z3JU9YsD5V2dyBnSGR4u0+mcKb2pbvqkxG
HkXLFAG6SbPXO8ZeJRuU2hDbCsRT99mmQ4qfB2jKzxAwZOJgqvF+6EeYdVnlE6EV3oq+P9SUwpw9
GmgLcQTVftS78dLYisst12BPwaZ4PAdOh6wOkQC4cqANJaQOgMdSQJA0PrUdmc7CpVui75b9hDCb
UNMVZO5eKpms0ChO13PemlkUA2sBZLqFnIxZKaH2ooBhaxvtVzq6jbuxjlkesGNVi7/U7hLd7Rzg
40DAl8NnUSg9NdgPW6OiNFi3eCNcTYck7JVHMVvAb/ZlGMGpMa0QnWJFj6ABoaxy2KcpOO1VvVmk
wx69VRXkADp6uvOWhNj01n6v9LpnCqycdhjbds3H2vUjc4CTStz1zmPKRg+2avysyiqq3dEFkyJJ
hCG1dlwImVSUkbahziynX38PmVJ3NC8JY4HZSHWjfup/KNEWs2hogIlsfy+Nh0AA4nqGsxPU30Ms
V+OUIAthmi8uRIlnx6k+x8IL/bossIqV4XbmekHbVHAeEWHppHaLVgtr0+PJzxU2E7jp2LdjVQdh
F09AJOrG1lNAoZVKMXPwpahYjhZf0FwGgDF2HaIYdbeuGRsevoscPbzTM96dabY8v2QdcpE9scm2
t7q6eMArXEa0jsscn/V/7ZErJk7hOIW9T6Samd0YBaCiiS1PzuG9AnCmYXjS3BUJO4hCC5U9wOuU
4oabFGdSMrc47RmtgPmN3F9oIi8C8Wn6V8zzvp4LC91NCdgfg6brsyhq8KQV1GmTSY50UnpctJyA
IR90zCFcY4aMH+9VzVKZFHYN1hmgW++PVmWEAlnC+NcyaPPGInvWs41YBvtk+JVTO4dqqQchrRbq
zsfZj8LbJ+bEIJwkOdRnvrwJCq8T3XNwcnnlLxdxLMW5Wc9c0yvuLO9BBL0PmTeyUvk9nh8BDaF0
r/fKcssL09xLWKEuidbMr1w8bk6TTY+1J/VaYT4tBMQmNPLcvV3giy3MUukWg5e/BHoV5SnKVBTN
gzOFHFQpKvZ3UicBx5xRPMN3KuQdUAa9Skf3a5ySRvTQS71DdcpBU0D0ac1ng6NSJIG2BQYjEEzF
UjM1ILViiLmGjcZDtHpcJsClD5fANmyBEM0be+hTVOl7HdXICzPlopryeMPZHoTvdC49UUIJlcgM
LuOaktbRHHvLe7+z87ZNSSfNCUSNVrgP8kugkZlf4wtiODp27s5Ze0Ay71ZY2R6dhc6i574Jk1Rg
M8oZDGS3ISrmhaCbXquGXtaPISiAZdnoZA2FO8Dkxh1yiBSdLTkjyrSFIHp2z0JmvDfYdPNtWlz7
dDVthDVDZhdJ8VuK/nLWkXUhmizXZP8DAAoiDttsqSo2XgaBd5w4kBGT8wJhMVx3CHotfIa84U6t
vyQZSIZ75jJmfjDJoQvv0CiL46XBS1oYK4Z4RJvZXEQbzF7tTvJ6G0dwKKc1kknYyyRmUukKNwdI
M7XbF3Xj6exxpLiQQJXtl4Bu9H9NjAqB29khWbuKbc9uKFzNLQBBF9n50NjqLJq9fFn+NyQFdiXj
Pevicw5GhAEY1r6sA/nuMOLumWs1KAVRFJ7McdAVPK8CMb+Um/E6Pv0fpUFOwlexXG2x+m0Xi2xo
EBqwNU0U2aP6QtaZu76si1AV/UDGs7zaIBWPLxFo13wcNK+KIZvFa3lye+t72dTuLwNBzKqQeZ6F
BIpWxz2/DXZkEh5Q2J5cPuxc3r7ugoHnjSmiIJXBT9JRLi+Ur63tKAxMDH7fJekdGqY5aREcZ6Mv
yiC5Vom3JtwhTgboDSR3fM3gM2DLS2HSNWdul20nPg/igyvNgnVTt2PeMeopFKUTCvWzMcGQqEpu
brQtCEE7RKwd+QKvjNHo+cZXanqw39v1V9x/amA15Ct23MXsRYuHYhOi0p4mLVdc2Xsw3e0kvhwv
kJdvisMaiTxnIkPklDzU8VkeMR70Z/qUW7vgLW4s0ntNtE80F37C4BgT2SB/BfIYYdsyWTqCx/K7
0FzbtsQHySAb8Ptnbydeb6L+4M1Z1vcyZPsqOkZg1wQdwVan8ZUULxpvTRNoKfQArFjnjLUu5Jjt
h74IETKoln6vwdFwro25RmhBVrEm3zQTMZ6UshIft0lZiYuM3lO8Oms/Xx3Xe7C8xL2opbw/05uc
eoc+lAHSkA7AeAk6mw7PilDACfVBefnwZVslrAoVxm1mJCyKldwo/Grb3stn+jFplKPcL1S8yihT
V2kFPpZpJw3MgWvdRsTUAXuwuxx9b8pc38sBJJOq1OC4J3BSb9AeDiUcwnSLicjUO6zzatwrQnU7
c09FFF/nZOmuwuhKXLXaqdPmkVx1w4X+6rHtwK8rp/Tc7pHzlX40PvmvQzu82R+Zxmg8rMIae9gw
Z2DrCiusdgSSupjNGN4qgu167dN+voZPfQxr1GOcYXBFlxt+X430KwSfyOKvoOYRheDLqxNSfRgg
D6ZI03ioqst6+sIxx46Uz832S6qjGGbmc6EZW2k3ywiHCTMhYvsOymGRZcieUVqwdaEeYe2A8ANN
5S96cbmUeJ9RfAh6OAD8lD8gt+gmPfxQk5Dx5fSgmmsPVeit4akx5jsOOTuesj9xvyLipAoUzTZj
5lMuPrn39+YjD5H7A7flGKJztv4yZxq/+BNNuuNWcvwgJS//AFcYjtyFmYABQFMF/x9j2ZTtp3bl
AL2JgYIlynzzhD2VTlrynlKrGODSwkOaKkT88Tm07jwqC8RHqX7quB60l7pFDHKxjQLKShwZ2NeV
A6wIOFxA/gW4UKGFH7D1OhPXn07yYTHSEhcED5XStbTx9HH0iTN81YmhMrYd7saCCbavVvI30G8w
5vSrdd9EZMDdglX532ZEjGvPU62ySnBPVtnRN+JM56K/d5sNgPruYRZtb59Nz8JklFI8cdlSDXpa
YhDi5TrHy8JKmScfZAH8BPNH+iknYNobmA/ttDchijPyUImNiFeU/+83EFFJpvPVa3v72fWI4y/d
Bq8MOVt6LulI0LML6rBL/fSPda6+rcRS2chocbXjTaJTQe/3lAPhIv9v4EmDItE6knXFjA8XZycw
NZo9pjkBSUMP6Au0d2W3qbHRJMHcCZvBu8NsQX1mJ4mtfGSsR6RbGWXeEBJpMvlHYb7iNWUhhRV7
t2Q47UPXbN4Pmy4N83Vr4le8EJe2CUA130reQG8/yhGjcOIPMmPCkJ/qQD+WRIbyZS8SDpfkkiAk
+SYqABTaRz35gkBtxhLPI6Serr02UD4TbqXYZo+N8+I0OHiRYQGB8gPbzh+8lRk0QhzNtYUDsOaE
P7VK61H3BoRmc8A3RN629orNm0nYlkx7upptH1QEWXQ+Vp5f6SrWVlel8A7kVHvbA8WGXB/eA/cu
EEg4JILrZm4FjyFmdq8b+btQmMeeZAmwkn/UakesgLvxPbrxwiEM2wlatCmD9jNtJlyQ4+N0unQX
M8QNVTN0nBvHeqDUfZZVBKbkANnSnEFhhHcCDcUtqitt5NhktrWO/9C6AsfTvIIjfPZo/cIhYOi1
X9OZhqLELyEtVJsxC+EHXAaZ+oBQMMW8WnXViYO9fWaOofeB/DLvm2yI+bHFiVQzRVtBecDWKubJ
Tjq/6gty9KEAiLRhQi9MS/R44UhfXTMQloPJeaCb2qPbNU8PLWORz36h14AD9SVvXOuLT3eakRI0
gvIiZpbaRnJVJLQnf3zPNUp+FtByKshZ84qQXeh8W0nMYN5VMDwAvyyuXXw6i0KD5qwoXHY33mbj
q+WwLuVnP96eAhKqYZjp13Il0eNOzRchxj0VtWW8Wtq4bdDhkfoxCTrsgL2vSO5eECmKH8mquvPr
X8PI57mdkEy8geB/HH9CoNmajDEkv8u/28Uim256XrYmsVexOv1XNJrEIHwwOBb2gDKv1z48tnLQ
3CSdSHBVd7Rq9SkYFhM8U3ANaTKlepXv7BUqzMfQFqQN50qbrThQxLNYOgBdONjh9cCzFvyZtvqx
du9CVRrZ1NKxfkWcYzKLaqFoKA67HXK0YbVz9rzo1qVALden+fxcI0vTVPiVtm/AHlUiVBddgMJn
SGQgY5R9ppCyPy2OrNCgmvnsxopzgmY0Et8cA02ZwwYaehVcC5ux5emP/1nUaMUMAHJ0g5UwSUQA
g26p9IYC0b32N1uSHjjamhrQ6D1Den/b42cOMzIHasVvvTfPeOYnV7RbcDajEPhHPLl/06K/5K1n
475eNE6ynXrdjiuBLnMg9BHGCA/7eXl4H4qdNrIiVwVmhL1czpPyC+lyJ7vpdxBpcgnnkSjHyjMr
pJYPF9SX9lmDUE7izQf9wjZ4kTgw/Rf6UKK/tvbGsRnq9vo2/gtxkE2mP70JziJNrrXuUis8nI0E
FSGZQTA1qaxSU+0crKNEl8PXzYJ+gR/DaTexYyOCJGlj9NW32lVlqQY0YewIIJAuNO4UAADQtlCV
jHNcSLpaYvytISQaLWcZX5i5fd28bfzO2jNcq0Cgu44vtgWC+bBgjJPycdyTu62ajihD78bRjSpy
BhYezOpEMRgBg6mrPggcyDSZPX2mJiluSdyvrMQRvpCgOarZ9ecVK8Umy4ZgUP8ct6e+wqbCPFk5
67uUeAlpW7Ov9tMuNRi3OFpKZBCWhNLYH3EIsy53KiBeZCUdTAiM3RRfcTlkQY0aUvdyzNp0fY56
w50bjIdflGAoXwydAzidbKdNj0qUxzVlVo1W5dAUa1lG9z1+yhlArmsqF058G6laKceSPzHHMhc0
FBpzuqLo6ius8txqD6KR+84DRLefS5i2xrUGMNvNKAW9HaU1b5+PI876KGxff2UEXo1sKpaAsNJq
DNwiPzHqNWtKlxo1wE8N9BTAyUJXquC0P0Curey8WCbXR9tKvCC44KpAX9WJ/pcDJIRL0kECUUzF
eGDU8bzd8so4HWibL0/dFrvl0rgBASfy5gsJfhXSM546QSn57iNRWpgrDAwHAFBMezJ9jbMZO/FE
D/zecuxvAi4nwd6YSI7BOD4O04pVrJZ+FbZF+WrhsXiCEZY1hdJuAPqV4nsG2RHQKVc8IZUlhYfv
r8/zVhiqoUUFV0/a1P2JYs1U4qOzs7aZevpkqK0zWnjC2hGNx34MIHoIauQtkIr0PtLkpsDbMFB8
aNnQF4eona/YVVw/H3MVCoLJdDFq9jcS7tUnTfvzA+27KEljj86gqdAg34jpo0alZevgL4JGGczk
awqYKvrkVJOOx983zCzMXhZCAcb6bGLh6Tal+KxfO8wLuiTDLXqlxjPFVXdS3ye+fBKXPovjt/i7
xLP//w1dNzlTbH9oR0t0bCIS7NZHDCl/rEmYid33bH3+zY67yTyTPGUerFtjQM35gJk4yk6nKbRb
NP2LGDFugt9XiMDJ29biDXEPCyX2pcKc8wzPe0TsKp6iaw87xmKll/GnX1IgeZiq5AYvLThPqmXG
tODsgWx73psBD9VMJcX3E8dqoyuIVzwH1QH+tiA3FNNRA0LWn3FXZdG0CHFT74QDupIFmePqzpaA
9WAHRlhuKS9U17JAgiiVH5vDlteKKDO7ccsrzsvFm+0Fq2UY3DL8yrgyKZhyknNR7EM8k7v+IAcW
s2c0T6Y8Eb6FQOnxRBZAYjyGhGicKpEI9pF6+M3xWZSlAw2w7re9aYy3LFyIW2NrE+Hzkaks0dS/
rAjTr1tjHYs441J4F3c9zSr523+TAnUJpHyaBI8Mc7FnkX2A9PUUxhapmILGpevFQJI4j4zpAEBr
61jizFIiL5zgF26WBf4aiHrXerapU+SCTL5y4I4Sfxco1GbxdyjtEE13XOmwyYq7m2paejW7GJWQ
uzU14PwAT4gV1EFgY0KOaAUgbEGmwbybOFrrMtmpo5NlzA8D+2byXz+G2l573HsbRvKEkfKR8NDs
ce2gKBbvJB+tlG+oPrxdhgZfLAuq1KAD9PNjsyIlycAxnG1AC5kSb0aJea8gbNP4gGIlVmspHsOQ
Lrrw9zlOCf3weHfOKxxoOYa5DvvlUy/mmfydeOEHLybvb7UIp+8YmoZ9dYyQ+sjJNqHQSOyrxTc5
1+oOd+7U1rGeIjp6tJSgB/5j7nW0W9SNgPUrSDdQ8sxCe8/AcC7ytKJAnYaMlB8rnqne6U96yn/i
eTtSMFzYiUTZUJk3HkZRny6SkZgJt+ZSzVV09aAG+eVLBmnpnnESDiBJS952vo/TYKVuH6Ylct3W
hlyqq2pHYgYe7RDT67skH8hbDTX+uWkgOZaO/TYw9Xr8gbf8i7tKWXi1AS8sIiSarKuIpBGr2hp0
reqE+PM8gNI2S+opWJ5P7cHpBtMZXt7PiY/QwsSPK2NV0aJZat+tqCK+8YGTaJNiWo9Pgc4V2WdS
ZIg8rPiTIY4AA7cSEdf8U+7W080Qn+CX1HjYLNbuBtiBgQCbojm8Kw2/vR7Bzs9MGBjfabVAY29t
hgxZDCinwsaIeW5jSTEHD/b7l1Zdshmmbba8i8AUYwtCeKWBhkBvtpCwlI929Hz6+WiOmzbhnUBo
SzoQnTbuGZFUjaTGfL9IriqXcns2cetmxtIVr2Dq3vfpa/ZC2iwuWzFaty6Rslh7ddC+wWzYTw4r
4mPzkLIrwu6Z4BEb/92CjKHlMTKtfTgRd0A9gR864lb9mcgz3ljW4l+ndkzWmzvgasxzaH3dDCTz
juss39hPB0qbP5u9y1UKukItgOZECXM/9f8rlrYSYqM8oZjyYlAN0J3jVnu6pIiP4NWpobpOvXf2
B973laDcmAVhxpYLKK2D6Q4OjKLNTWZ+c0RNztzZAcR2ejyKJe2nSDgqQtFtzompFvioTB1UQNJh
OFu5ekFiqLFmAipA5Y1bmRyBceWMv2nzjh2KaoCnqw631cCXbjj0ZtxkH8SCaG+JYXnkHjh14WtA
APu4jPYkiThrEBYSe7PlbUTNxV3YfrNdhKf1kEl5DWmygcqj7tr+kDXpXMLJ60P4zsVBoalnouGV
WQoRo2s9zj+ZhjMhMCGIVanB46edx2/fzeaGFkCf4M2h412fC3HT4PczA7sMaoTXRRLiGQiPnqPm
Ur8QNhNfp63VCfWpH2WLcIfYsrmUI92ZOWM/f/p4APM9cEHr/fJwraC5r9urBmbzt83w+CyK8yz0
9VOm3qSOCChfMrNGmAWCq+CN+jSiFykzivflquQSHfWsLvAqegUpfavJvLZUaDouomz3jmljqrmL
/h8oHOiI0x41Bj1dttSevnm3ROr7bgXJrLExuAA4THBvoIppfyret8Rn+pTz+vdUWXuiBGaJn1J1
OZ1mEJdiCigZUwi2C3vltD8iXfSC4Z+D2SvK9FZt90/oaybJNKaFOErowPpjGuFXdPI8h9lukb92
OM/yKfyw0TGy87aGR6X5p0GvnWh87cpxCVce2I1J9yCf7lR1OQhIA+0OYww/ERoPoERRFzYuELp7
Q13J+QVosYTUdmB7ud1LQvJfS0R1BWLYX1fjg7uBqPgFknreBFJLqid61xJcTmypn9fYekY2phbf
QnA7hK80cVN4G3gB/CXPPszR+f7wSNkHASc5QVyF3ysyzWoKdoOJi2AMlVnU78EEpKc6BiLW/bEC
2KidXNhWnpUdPdlUe5R85omiyk0m/NZ3DkyzB0ge2qjpsD8xLaVb8jtq1vh6RSo+rofqx/HS8HQ5
jEK42FOB8GkDBr+FAClYekeJF6jUISmG2/8Uezl0r2mdd/6ezEidqNQa6e7Z0peacGjSkQwCvAl9
e7X97/hJAuQMSPJLjpDnn6GOwJchTF8NFjnFIfKDb1Pe/8hvyj6CIfxRqWjhKEntZr2hN/eko5S2
lsbHswhNClgyFe0mUVtlV2pa//ye7+gzRb9IhQYqwOBso6V9/x5dnPWmPmZScmrTnFDJ4h9m0Jhx
LWLSgqNMDkaE+iNQHkoVP5POhGzzL6SUG/e8BDZi11gZ+mVqYdmgBy+tcVX6haY1ChnPFMx8hbA+
qMpi9yhmkksiEVy3iXmHLdAcEF7J31VfExutvsevuc5qh48WXes1gdC9ACrvqY24Uf/WjiWeVlLV
e/ULNC6ZnajKqIhzoRGDjTYE9DWOx+SI/lMrLMRLGFRR8zymRQZKOkYgihmawev4dDgV6wCXNvmL
jGGD9r81rc5hdjdMiTASe9QvE+l8ziOidevIKRa7LXhgg9mUQ+6v+k9d12boxofPGxRPsNcPc/OJ
iOV0fNq1DtWI1DDDAeIh92WiTue1evy7y3+C2hcP9uj3DfLC1jkcfRhwWzbwDNKSV5bpZo3Ei+ob
5fKX68A9Z15SW/Cu8Sazcn7BMAXvsXOmzys4GiU/JjjVCRKNmWPAvBtFynuxus46LpkhI+GdSUVk
NyHQfOPEaHAYUImeHfwRgOG1UnwEj9FmGuq6DeO0Yei48sJ6D0Cta6FVIJEvSBXbYgL982QRaGMN
EGIa1AKDe9d0nuvO9WGmMhwpW3B3WDfQs3WZexaoXDKdsbfP26mfozjDxlLtnvk+o8CjMOKcVgoj
tH7ub8FpHasA5OpzFXtI8LDvViHZklOMSkTm1HCsI8Lrll0UtzgHPvcp1vpny834xYzcUMVfXakW
iIknUx7nafi6BzyePfv3JOWT9c1oXjKl5M+FyI5QMTMPZCz+FKVpmWiUtnH7abZsVkYofllTKuso
DeD4e0FhPcJ0bvv8lYTITfT+Pt7i6i7Ak/dNr9iRAtbv7dPDGycguGkmwPr9bD3Kx80fNBvKYxjR
OOen9oyzOOaQuNtewismjE2sVKOnP/vSk3Hsp6gEgYX2sLfyE/YDPds/luQ4mJVE2IyhTqCShdwm
I5ukGkufeSTcH0Oa8NHyqKaZOSSigd/Q5mQ79tklBzjONXaWzp5crOBNWfz8MbCK29I5+ra3hmMQ
27eO+k8DEAoYKDXoDhIsQmtF6E31Fs0r/3k76EHC0de4htjeA/TyOK7+ELz3FNNak9ehjEWz9aWj
8t2czvyie1lLluC6D8ZxCCu3yEP89agbTHrHSIOcANtbTYp3UlgqSA4NnRV8asXU6Wdbe1NK3hWR
va+ZVsO3YN/TxkX1W8YEcR7N7j/VtIV+jW21bKUq1vMylJNbdNe0Yel8aLkCU+yNVZ9MmV43U3jV
gr3wdvfuqI9dkG22JI+74T7btXy5t20dq8hOEJQBERHxAkxa2pZ9QUAsxsj8mVyaBMjUmmP30XzT
V9emId+Tq08F0R2u/t9YTBRoWvQTzpkCJTDxvHpzEIKwYNYH43qCDjM9YpjPLGO7SYiopCH9B/w1
ODy4yB+rlnUQeRXAN/aQO0C5ZT2i/rCFTNnKBzvcN3sl05mSCywWdeBx5sRMefuX7q5RFx0fwwXu
ZiXtN3EvYo+VIrjnQQ1OIU/CzIfilGJFu9VYgrY5L9X7aZ5DCa6QMwZunLXZ9sTHe1CWRnfXU6pj
wxyMIcrJ9ZYrXriFMvKD3rQ/1m9YMKAwVewU/0wG1hNJdBjfoHGNVxgME0gQ8bAYuQCKNYOwB1jD
zREzJ8Z3H0FQy6Dz185xB92Rn0QVrbXqX8E9YaD5gPifoBAATcbTBlgMVw7KTLD8BpnhY51FR7Xy
3kC3kf8qr348LXL/5YdfjDegZbv52A2koj6m3ODanl4G/37kpZnJbDS0EuZEY/y5tiz/9w4YjTDV
/AKYQd3WTI8+QUxg31AZ5Zo/60WJvILlcUwXsOOgAYoyKRJmZGPAHugmIqblGvd7WVBwnAPyr/hP
T7ZcRRQYRG5fiIr0uz+YgTqfEQMQc9jUqklqJgvFDid6KPBTHH0vwpViv3/AyyQxMwSjgIiJoLcJ
5k1hA4/+0reem9rb8MLTypuepDCEUddM2WAMjJ9Wyg+tf8LSZrbX4QWLyKQ7elsQFh5DGtuYQ7Xv
TYnW35PKJ+6YiqYWjQflL2D29cb8KDhOlftlxm1x3jistsCMvVF09OzLoNxh8vub0KiUV2T+I+y0
UaGXFyDLblFflCOMO+jydHYuTowhhNh+GFqR5Sy0JvUbfK7SKkM2VTAoPWnPKB20XUSYYuOnIRKH
G77pxxTJcQncxERt4Xev6jDQvz1/gayPEL4FCFWRkdNozDBIMdKUFHm7nttJkpRE3vmG+dNnKgUs
//RYfv3lXfuVbn5P9lQAtfNNT+mrnQXBu6FmiCeee6ggLLBHFw7yTJEbvvVkUmAluGFnNWcJHBu+
SuNO9C/Hqm2Sel1S7y+dy5HxBcz8IXAs9udZJTVK2gUg0PGUouVQ++/FxtKZEdzwWxubo962yXRA
G1iILYRV54h4P08rhWCdQM5ngi2CSdbkZ7icUS7WnI42KiCxjVNKyoMb+jGdoYvKmFRsBgacA3Ge
9TjpVUl7WHs5rZOP/DpOOkAf08KQZPMaQLNb5Nd59QbxfaQ8wwGcb9lekFJEHgH2yS77bfGlTvhw
q5fKJ6VmlW+oJCv5knoEamuHqYxqS043tIEKLtSzP1p0JIMrGIn+3iTFEkski1yL+AXt0cVfqfwm
rgAaSuzn1xzoSEc3AENd2Tn6B35sjHNAX/iV9v/2iBnDu0KGEBDtiDHwKfddH7KF33bNE7fcTPiV
DVT9z3WAUAH3tQTBPLzUgXwSLHfT5G2JJZjYjbncnz3lrBm0MbHEuZjsgMe4WNu7as0eCdjg35xl
RaO7h6OkE3vIEycT7cC54QlYgdhLDzNJBpIbvNzjlqA5TW5a+lGvRTjSVxnqxnksY+ARbgeZhT2V
MIzlyC3yEwNP/mBqp9Ks1t+t/Otq0QLkE7sB9DS4CtzAXTxTqsOyFdXJq9TgpxsFifspFaI6/fFn
7DlPcEtQ1wf8uvohF3c9Pnt3D+ooFakMeScmn6gUKhJnMnZTTUl6s+nKXkMZgVcDqrT7AeofiTqI
hwM9LUAZ0HI1HJWZHUl+0d2j0G5hwf3pXmoV7HBh8QYuphMEFDQf+/XWCUP0SXBi+FK7odsdTdvU
ynhglBrMGxYb6LAuulSW2Wxe/Nnc6yxzlSVF/8ClXOjrMgNNHfOWo4cYeA+fono+4fbVaDlR+c2k
47XoXc8yL+bYQBqPLklnMsUUCpWnyZvboWtofaRTI2eWJEHPUzdUWXhSrtW5qMxYQAYi8jcBAVmY
H8NS+JLN4fpY04JgIWZ4uv3Wg6g8oKmrFWPlvafRIByoHpGhY8JW2nbwjlg61JVVhjoqZIHRDm1U
fgKm3+kwcTnNqYqVQTbRjfHQR7nlVqIC0x4DgfClKe7XqsdY1nckUTfCfc5IiQqytLCWrCZ4F3dY
EJJCu8nXZCTC+OwYUJUkWECam7cdBAo1K+jBQ7AkMm+vgNHqjqZDiURcLVVJGXF77KGxNK0TAg5s
pXS4tzhOkvyS5lcjfRzAWRTpbQl8hACgc+7AShPnaoycvxyu/vhM1lr+gKvnyMIA06wN1jK9Hxyq
WxgVgqDlrL6ULybssFiDIg+Vd/OFqDJu+W4QXNyRK3QwNhUG2QFZdX18aS2e0/TXIcJQoSBZ+J11
2C2K3rDPMH+xc9yBr3NIijxKd/xTfyZfnR4I5DXl7teXFXEwT3i7/1MAtfjuweh8VfgCrbNRN+Ti
DkGN6oyn69leooSI5/9bwhre3b5Kq9IqbNj7GlnvaPO4WeIIsRqZz86AI/gNqPt+ZMMABePPC77w
tkrvO1tGHUTSVBKrHTvzZujUH8ZJ32b7rlLYMeqiNgcsJOHZP4OFIWmKSE6v5f7XrVeCtl7N+USH
2FxCh0UHnLkcKmVTimOJAGzNem52dCxpUUEU/tRG6DED97szEK2xrAs2DUj4Uivm2td5R1kqKIEb
ETRY1pYHgjW18C75BXV6sWk1C1pcxadEAfc4OPmBkV2PT0zOoJDZma0TWn+bacWiPlZ+/mLmjBku
3Z+vT8DTJfPwYn3JsYlU+uzsG3uk6WXhSHMjezf88OsyLcsJO7kEvxCOruKH3CRKUgH9A0b7XXdH
vk0dm1lrnJUdMG/XleC0w4+xwnhhgyKZmhfrQjSx8FOP5cIv+oWoohTDzeEptgUpQyNqfZBS5IS8
8FRjPyIJejTcQcFHHknRjiRMntBrkfxM43pxOliWEMChqRFaEKCitRxDesA8xizhFqQwQBOcRP4N
XC0My3ssN6iwWCS8cGgt3D72Cda5ibD5g7Ieo0ncIBafhvd9HXNFoUGKcmYWZMCgDmbWqLW/l7WX
0UArBeNdNZfkZxHDh6vvtPT4UZ3+sPznw5tFY5lwQxHSsMGACgjwMJCorm7ZgUXWKEbroFGzls5y
JMq62q8lie5H0ew0bKCiGWkcNb3vZaHbNG9dVhuANvZNB0TlWHmGuCsJyK9nwSuDuUR3G05lpV2b
gByFffsiYP9De8dgWaBvCozYsrgjvC2dNvrvwA4cAOGM755achj1PiOqVo7G7EuqF5BqZ35ZUhn3
Rgvgzlk3MCuF5bxXbyZgjK1rWRYW7J62zyE59RMeX98nmRX8FvsfTCCxgu6naeXcBbwXtRDPVpYK
doz5spwL0Z1VNqHCowzJMcEXjlcKE/RllYUatHSjFRQ3JbJwo/w6CL7Y1b6x7t4kZGQwjV1rt4Ef
HMNBaJCQHHi7jJxWhC04rkq/sETgeWx8JKdlPhhKq5VgKrGTgsBSL0NEc2KI03ISR1l47uCl0qvP
OoQPvJVsVxFHynuSuP8llr5QDPVRLnVGMV9Haf5AB0NxtrOuAfjgk8g5GCqHE9i4D0tjMgk1kQYX
hnYgh69UBX0KZXmE3tMeeYzBKhF4bx+yX6Ov+MYpN3TiWFJBp5hFwcOiB0pSbYmz4rbiM6Y82C6k
2MLuN8CWD7hB4Kq6TBIugP29VbzrK6Uxxc4fw6R/DcRaIziYbOFxls4Yb+p++RQ0uvc/2W4vLJRr
n5CXgpYl5STwRpGvqt2j5kY2ruD5ReK/U8itjjwzfpvVvD8hfEwZYLbPx8s+i/yvpG4y2vC8EP2S
jzX5Hj8Cbk02e6i7jLDCvO3JuLzNkBrS5QiO5tsWHWvD5jS0KCuUAbGioO1n6RS636yslMCw5us3
6BtL879s5bbJyOYIGF74IkAtw6DJZu09UqM62254lVTK+VDYniBuf2W9zaNafIZEG6nQzNNHJR+1
pcIypEq4e8CGgzXm5GbhPE+jnKU/0KmIyF7swS2Qg70Qd3D4WooHHZn6z7LU8m11dMv8vL8AXGJv
zI//Ro/AqC3ht+4AgXGVw6Voja7v6BT4z1xOUacM4ex1jII2USP7KcTZGkWOyfQ7Cy0genQW/n2J
RjP++n0Y0fPII9nYzw4AqhmmMDw+EfOl0ERWwdj3WDWhYZ9UA5mPlfWFefzjJNRyeo+RUqyPNDpt
fQ8pVA0barKpi+fh6cngBfAgrCAIkltzXAhtprbFs6LxRBBfT0W/EICeSBqyQ4x/mUckhD3F5nIg
9SEZlQG1ai6r/vwkJRJyfzVI3XpdELzmPqH85Po+3wzoB7NxDiSQ/9FqYLLGIYCB6Rgkyvs/VyZ3
4eQZkbQpcc5qlcVpxxGt92y/acS5JqyrYjIR3CzihMrW5/ZPTd+ucci/XrGx4WxNHQrOE21ER46v
w5TWULNuVi2UoxqkX5MKKdfi9kB8+rpzHSGUY/1NXWhQ8EMPd7lD4QnPEoT7IhT1IVFzFvK4pHq7
6coApbyRbKyLg42NHSf07/zByyAhzh/4IFkXThi7D2Wm6hnK5PHo8SFBSN9MJfLGwEIKyldJLibg
EkkqkXX1uDZJhi7WyGpM7t+Puxoc9oNiOv/aRO/WAYkf02/Q8mQH2iQNQhQL7Fj1kwtDCaCkrk8A
pTyiLaDNhOin5McD+K0KBFRtMxEcW/gYENLO06+YVmEJ2YSardkepLEPjtTrDN+ZqxjFDHL7KbdO
NEkF/6ym7zZkMY1KyaFVO17bclo7CyEZFtKgt67mUNrLeeqVHw4iCwkphM2ua3PX51RM97zhyH2g
e3SBJD34PT6WrgRvz//Jio2S3r35AgGBtX8gfbZuSgxa4bdCRz6i05WlT2cdMjOeTKMwNGdqvRNm
q1U5Kc4BuvAFW7IBDHDtyFP1ueHS+KvlRQREflDKz5hgPXZ81yT1V+2++pF9gbjKj90gMv5CXltn
Yi6xlLJN07PVd1OMn/PDoIKfl7v8cegJzSO8HFHMMeE8NS0RhHoPIK922ODudrD/lay0uio313tP
BXULPTUwHY6ZwJLYuRtG6stY1Jm17SLVc7KcZRxeAOqMXpX9RmOiH8uvkxeAAwCLO5vpTAwrBoVs
gS2Jge6PGLCX0hFeJJXgnoStrjtgvjmETxWVnluC5P7/hlL5PjVYU6OSG42zl1AZypa7c9AubAUj
GNKHL/3W7Qvph7zV3w85L1zYY56MzumV92mqD2f7EMGj+YWSWxse0rkQmuhDG6ByZZ0tNcAwy8rt
j3r5v1E2tqUXXZ0R8P2RA9efPlz94g1za25recBRTujXhNuT16Qq1gJShegIDYJfEuW/d2mqBzr4
4yfX+hUWa+DM/WVncS6pU1gsb6fGxPZnUDZMcDxaKEZd6JRapmvNRNabhtx4/UTLhzmb4OG0+KoZ
a78+y9x9LGJ/IiutKexJjiutD/aF3CVsUTy8X11QqobuDVq6Xb3fwp5Do2ckiQuporOI9+FdmwDs
NoSq3biA5tkilG1ISxZrBb+QY8YH4U2s1Rp6tiZebEgzdUesPieVYRVT3IHFPi0TqWA9jX56bU+y
fVf7ixWfBwmj+5kGaMfr+6/NEpv2CSEGL2mTIMUQeP5JP7KT50bxJCBWHc0g9DVq8BZteLKpcRn2
059HTzqkxQqtGgR6Sk7OrlD689YHozsEhv4iPfUULU72jNQyb0i4PryvVE75s9fzty9hfL/Qk3jf
hSRPN1RFJPO6UocW4MNxMcc/SiSrOSOjODH+4w6irFiIlUO/D/QEdE2d5jeBgzlqUXPbeq5G0Xdt
1ZS8z+4JQEseeK/LV7fQXkW68oBGa30dLoq20aTKPMx4JmQB8QlhvK29jE8qMyjVSHewfjW++6ps
gD20m1N4+tuj710etK9WKW6o6TvYhLtk0o0qURQ1/yTxqsZffwrNtIaHnLeYe7RqAxM9MMPUkI9K
4ijEGQUaWeXNs+/4/MDB8oBYJyiNBxWmwYRqT2xVyerQiWFpKrh1RENyloh87mdN2CcDalACo1B1
ygbGuSm4cEEVDVJc6/1Or4uLK1WB+x+9cH16jvsjwlZ+pd2IEiVRG55XMPuHE07ggyVwSsTLhuQx
JkU9Xc5xSdY2UrKdl+aDHj3myy2mo2Tl+fYzuScawa28ggSqslDAWsKBfGGs5/CxQSrvIcBF2wnN
wc9CIwVCgL3EoHpjYQQB04HU0WIPxzbBY9BrZtySgTM8gjWymyIz0//gW8Pu+2QnuUP1aTO7hye4
b7GrjF0No56N3uOPYfeV9U4mVNonzR4NDDrn2PYLQiWhxemxRsptb5pUuF9LnqBeqP79KZ14Ghby
m2E2QWvIkf11/v9p/M3nzHiseTNEPW+dhhI98uxY0tnNMF4Uiw7h4I7HsQiV6/A42x7Uu9BO0uqA
K88tQFJF3iZ6+fumoSQQgJbuykCtGTBu3LXG+ohZ9FJORkKnDsw1pcpOVu9TRRQQi2u4KPIQrQ4v
sONuqlU0mhPzglE6mrtEe2trEUZ94/vjl2jBBmUpYTzq0mfdUIgnspf3254/6BwJakZIuErCBVLN
TlTtgBqTlmiCp0mVjGfBmeHt8nE+aB0p71JKqG5bHqQYlDDGTfhO81sQYoQ0F7lkl0jg7rGSVEdC
t29ykdMRjQY8TM2siECJprsJDA4MYJNMDZvg9+cOV2kLe06YReWjyCXob9tCc4uumW1g8/1VcsTk
8uqa5wIpyx/5zcAfa73uC2eSwkrAH67+l6x8BvyujO5ST8CXFWG6oy/y6nH5VkYj/vHjbVSfhOwa
3o/CewdxzAwizKBiUZ3j2TvLM7OYD732uxlmb7yeAbvggD47a/ZIi2D5+C1RaNLJ24LvezKz8GPz
FNPM2s9ds6AhO9H5aSBbr/t7YgEn3gW9FVlw7goXjXQfmorg9x4F++rgJvEXQTjeDNmJUlUslNvh
JBD73MK6rac4/ICbtM2L3kxcJr+88r5oxJIfGwWjP+ffdjSpcHaoqqzJWZ+La3jkldmW9bZm3y/h
zfD/pLeXepQQskCzKHuM02u0loqcwSTGzLocHe5Ma0z4FH3L4pPYywZZeQkGzPveuIUiewcHXoBM
Ql4h14rSRpfU6PZwLpIa3qvC4okKb9sqsbsVdaVU96DRuxl18YVdEvtrVWTjP/bvMM/KRIAO/buM
c5/byjv8ivLg1SGgD5A8fa+y4h2tyzqs6Ec8wywJCJ0iW7y7eV81rINam6a39X+R2CTxoKL0DVIa
EJdRKmeJEyuc44ziE/1Ezp4No6hYWB3DgTptyHLCj6MdvUXrQ5oVLsCKTbpi/ksvc8BS6J5stB0n
AySUCItw4e/ppgVCHO/9OGKIbMPU7jx0XzeP46fxR5DuaDbOFXunHvkN+3FzuZU2FPExmwe7YMGy
9gUNRSaL3/ThCosSDy0z1JEKF8w/cf8xeSJvAoemXnl2GVcrXMS/QDYblQxgLzp2XZ10gLLIm4vZ
Jkl8ZQciycRGrKIbCUQan4Xz38MaApNDdzYbt/KuA5QzWKwCcDaklD2Um/EYanz3n9yctm2J4m9E
h9p2+t9M/pmLXOfFkd+gLKnhm3hFGXq4K4R4jb1rZ2W5+mo0guAz3bYTcGd9PqU4M2h8eZ5E/GhW
6EvayxyAllHqTFjZ2MGDsUPFLW0jdDnz+dYAEVRrq6x6B25AR8tFF5CZWXz8vDDxg2qSVCMHeiZk
NWmmAPo/2sHCWRx+bfqVbE5Wq1zWqchCoyyHYzjKGt8+CHMvql1X/eLm2F1xaGHEH4qwVhpTnm/V
9ORdGRI5JHToOLnf6zB/UvTIb62Trh0LpY6JOWC2wa7Jq8kAsmLvhCNxyu/3d05+4OUVkIbd0yk1
cDK1d/vkGfzqDYhVUhWSsTGMcPsNqkJGx1dzRRc91pzCg4OSRbZKY6a+DsyWyQG3pYDJgAXfKK+Q
B84CHHLd/qLo/BtAGpmopd9EqGZi0rnW8qeXe+IwZyP6BnT8ov1SlICZ3n8uNOeB5xIQkXnraDi8
vsHOoF2eRgWWahUMe61/wnNebp5mJ+RsjWFnYSvyNF5htQKb/94l0Bd00L8WwHoUj96lOK19Y8ui
lYyn2YC37gV8CR7jpT6gKm6ToiMU+Jb7jPWH4RCH8zPiEQMq0JEbPQchKl23l6XJs7DmC4pht78E
gbwvI2dnVDkW8pL9iyNUHCM4bFKvI/ipHnaWCQMWyhM4ua/sUiQxxbVkb1TXICzHFCEKhBXZE/S+
AQfHKgFZ0IYMTl+CgfhiTho1tnrufAr+BPr82hyulHMU+zFiylA2suxD2+kEluo2EAGIKWU3Mzxw
qU+jEG52eneukFXjQWjQAnHBqzyNvRTM6YCERSOZtjPz/i1Ez6QLmyPtE1CWcUsimGXk6EnOLhdg
KE+fhsCFvhLAJwXw1bD/CkIJa5g+4V+/Ye2FmgZhPTDXz8EdavTk3NSQodChvbN2op7NoolRrr6d
ot1vJlX0ewfpAu7Zdjsz1VcOjCkN1zm+QGIlatSTAvM3lfsG18elTV7Jg+kmZx8pNtM/5GzZgt2F
jywO1ubaWQ1POxPGcPA77J+JVMDz1JLqV4L7YkOhoKw7Yz2k+7KHCfjouDQOgxNnkNm4bWjGFkXe
D9/35Pwdc8/JJcHA/n7oK7vGJnfkqrQFTi+sEjHnmreLYOHVhAtF2aNIk5v1HEOfvZGNZj3EY/qv
JshHCpDUjj1H6tqPQbo80U4O3E2/rtLkgtzATYj7w8M9ori9/DfRRx5ayTRuoTajYquDFNaXJz8w
uwnFypqk9iQJPrHirmEAaw7UHxsAPiCPqz7yYiMOxryaCJxTb/yGNM2B5naQRAA379ChBW++k8uS
Ch+VnjbuElyW06To8D2qxAN/GS3qDzf4JLvKAFSuHXfcVZCwpaPtoZOU3AUuStDu0DkGhrYA8hGD
IaxGJgHB0e4lIriEjbxdsNS/dBTxi9wcJ8lImwfpR385EEvlnDjEbq81QJH1cM5z+o7vtTm4LVQG
h6SqTFCQNo62ZTETy8DMOEQ8oi5Azc46cszh2LGPwBMS0BX7dWNiviaDTsuLAxMXuyzI5K35E0yb
Opye87UPUVuzgjhGmORhkPebyVwrMv5u7l6bAYwZA/AebKcXClK/kUtwr8/hiqvO/guCvzHxaa4A
N33Zz978uy0Nz8lV6WVtSgIBuKgdqwmmPSddmGKjGMDnUkHkdyhaqwfgJDvQQn/Lb06KEfSn34j2
Dj8XDq1BaOkZQlvPXePI1xyb3jtd2HIfyoknv4Cx+rT39UTwErxDJwNXsq4e6QFCl6AKTn7ro5/t
8Hk9v+bui+OVrxxkho3QYzZowfvOFXOWerKUz7eeXxoT1TW7aNUTfHo5kE5/thf0BFr32Kz/BJCE
7LGelwfKe44s9NKwcvngcckJ1WHdFsZFQR9E300CRBfb46XKxwyYaaF3Mch6WU59vAujJ1HmKj8t
KcIQtLvFQKF0BleR0RCDwQAI264kcUWS1/VGsK477Kp5CLYoIh1ZWnHhiGbBqAFmfk54SZg6crxn
0ld1+/0TW3R04JBwkaeWuinU/MBOCnJUYYpdo/FFDRk4nOnYLZDunvAhuDooHogUBpFQvKwAm7FT
mlWl6F3UsOMVeh92+jumN98IY1ei6nKNUEWhVx7XnPoFr7xCOuq4b4zkY5TGQO19dtzaZOsfbyXY
eSE3FmEy68b/bHshT5ibRIcYv0TxnPyII1cOaATyl+fwBxWK8mIaxJExlQ0WGX2lCUVaf0ASUDCH
DCCaPgDZX0/wuCBe271NjcQtdRlvnOJEfEI4/Boy7hCfI7kdWt8d25Rbas9gCn7UZAtNkIzgK1SV
B0nzVuVaSqKPrS++cxlv3fDpoAAcwAKbhg/cSBiarcLBFGNtwTZTMh6iR4WpXCah/+Pk46gvZAWc
0xN49JyZ0rLMI/g6p0UMsx/cLFweJ/iylOqGP67MbmunxEQfRmkILw1QfJI923hBipvij72YTJDO
E1ynGglhEg0mP6Y+hOLEKajKSCcULM4mMT8hhSDOVndeoN7SCETCi8Av+Gr3HsLvDdyIE2XhRHLr
6JvJfRqPnojiEtazoIinfDPj+uVDtsX8AuXrADGbdSF2VsNM5oClNQI6HK+ZSaDjDKy4T6ClSKQ4
InsZZx8SOPQaS+rz4rdd+IL4H5+FU9dz2dkYJ75rx8i6RpHT80yF8Edqd8i1Hmz+OfLPylKKGKXU
K8XM3Ajz/sRguw9dqIYsmE5knLif+nR8NOtX+n+yXklSiMyTsW+UNWHKovDFliqD9bU8PpVKlNnE
V80bGatruY8V8ZKeZ2pWg2XvbrXaDOTcYIxWuS4GLdRbnc8/caCEfQuWxS5lPczCmZ/JsXUld3Ze
TeOI4DjW2dRp2i3Fc2Ip0wF68WPStu8v9DbtxtuwZUAbMlTiS7sdsDqUmruSMM5P1JWbYg3BiVl3
lVJSbnoApxTuDvDCgpx/oFrD2DCIs/sAj8jKPEiHq5PYacRlfX4039fqJEhe1elE7N07mlQjX+QT
+D2FdywoPuAzNY5hWHYIFi2yh2a3etDmmnC6iH3LGAImmaTe6IbFFT2xqlpRlYHaVA8QWXZSOqFS
eXoFdNjvepPpf4L7Iqzdvde5Z/q+bRtSfjNn5XZa8eNtXQr0dKkRTJedjndnNJBb/AuZO0IynxO7
Sr4us/gB+DkVC2/MWp0dYJ59A++mMal/mDDMm7Splxo8sSdcpus2lZxYkDJYoTA+MxuFh6ssK31S
QaKuRHJKD4I4wsgRHj2iIDWLhfr4rcVUZ0VXvKKO8pHmdubhm5u6j3f8ZpTfk8ZxjhmGKiWBD9UY
ghG36ORpGoM3/uFQrm1QP1xw6SbK7Bbu3357BY+FGMFuKHChCUF5d+w9FewKR4Wx0JCjXdcEyS5n
pvuKREMRuBLTp4pgp7erZu6nO62KwNb0/QukVqL8+yNnX7yN+meMmrnOmjsjuoebf5k3hf3BMAAm
4OK09hUE2p9lr84XlOMtmXA4u1UiP04eT554c9kKVJAvHSWXxGTlfbjmOxqVe7PNAWaV2yzV3Cfg
tXjevfZCOadlx2/41bkRN7J5yNeCNMdC6pK+OL/CpoPvwRANbhGDe2gqvQex0XCvrdGa+CL3z94F
z7ZumPyuBpRSS6CUmpmtlvzXjRZSPr6nA/w+F9ddAVsDq9RKk0foCiK4m2TNY/zrM9vIe6Dv6Sbj
tIpah1FL9YEqqcqzSQ3mdgN/tHoHZTDuYdfHvg/T0wUgR8chbi3KMisDSdgoR1HwVhi+dVdroxDx
ah4aHZQvmZ25Zo76pBaCKykAUmaFiCBcGCbib/RKiDuZ2uQ+jtByX+0HnOPZgozMkg8J4PzwR5nC
p7mtAuZ0lljktXWFLmdHqmZCm/M9iwnSansDgKQLFzK+LVYk/NBhU+RohM3OFAx+JuVQ5Mo6MO9R
ToXvDKUYUzHYZ/3XF7DrV58FRcSq9rJsuMEZP+Pagpg5VdPGeadaH+7pj6hrhI/5UmdKPLntJmAE
SXOWlrWvr7LrjdhoPEXAe7taoDtQizRJrOCHlbUrsJpuF8HjCutxEij0I0712zjTwyGCYnkGmPOa
IEhkltqjOTmWQ0sWJ9E+BRtOL7oLHK626mq48tNb9OVqx/q0HKMBYioStWMrASDiGfydPEyXUVa6
96nCr0wH99ANtPu95niLdtTzAa6cPpOs/mcNztjrTKpDbAmyDV56PCWKJD/c9rHnxukMAdW1abEa
eyG2RTAmg2DB5/mUf6pDIA8YTbtKhOCEm3sFwzi9P8n1OgJP/x7Tmdfib9xX1b3u/WWOx/qOaIQg
piMNpQFP+nibYePQ+NNT27IbQzgA/wuUPa9KbdE7IQvZkrC0WRMka2lKdxD5Vy515e+FKgsr75Tg
3PpAmK93l07MThPh670I9KMrGuMdimCHaCIVepIvQ0sUoqmXtmNixc37C2y+EJsM4xSyrE6WDKp4
iTttlVNblYR1YVAxBeCkNAqF5Eo1ROPhyq7/K2rCgG+OA1U10fo10By7UF0bEgAU3cbez2y9njMi
r4zESs2FkJ+CLxTEy3dhr0pTjMS2ADmzCuKdZTgLhHNg3JgbKaRE+TjajJcdE5TgQl/1zlRZD8hf
2uAcvUBUuFc+cM6NB3OQsLPW5Cjac69yW1ko7MIE/iJUxBHegZu+TVHoKOAtWhKY0M7ydNp/yYby
QFcZQNxFZ537/8yXuQliG3Ch2gqD1uKZeBXeMbNdXLPdtRY1CYh1trvl5WvS6PLfpROsMawrfzvQ
RdrK9KPTmfZnCV/sTL+yd/idEozdjcmjdVAJsybfaimXyoIxUVbf0yFexJP0HHZ+gIl278T7VCBp
Sxf9JvA/h8dOH29/UzcUBHD0wbnS2fuf9dyfqGuvi5s9PhGGDA3zPbsdacgd+DblJAPvIV8KnB5I
DxQprBSQWfi5WJ2sbww53ddm3F6FCmktx2iXBP7AXaX2Bgt6zbpXGV9k5vaQfBPweObimQNXF9v0
LfU2ztIGxJO6juEzX5wJkunjU9MfcsgkXatsod+O6sqsYFMkJqOu5sUN1BvgZAY6ABXTxX5N3OIg
0ze/5cvLJBj16ytt8o+QJfsuguX7N3NdTV82fPGp/0sMAL89+eZ9o/YuEIueUlDkWJATLf8jsoct
+KYO67lZRU7RI9PK26tlpmpdUsn3/z78oBxW+69OvJRS5ep55m8dw1mYa+qMPiGhGnjDCAVg3Vsp
y+WzvYZSuSjAH7Va83IM2ItsF1p40YL7cJ7VFeenIjvvGwGeozSh+gpBdihS34TbPnZPO8M4mGSi
OlOWpokRFKHYaVYjorbYWZkYcmRT3xsctRZbWEG2ihxINil3qRBPVeQnlxdJJTEQBRY5MITDnE9L
YDjjTgl+DBy7A56UdhDChJgZZl54TMxLNjvDxx1LWZghLjXaCLgTPtP2TnnSfaxXnjRD0SO/5Zu5
dYXLjZB4ls7yhjYGXCV4ao+7lRyBjV0DcRmR6dnu6Id1j+jrQ4Cxr5bwsAOCzWU8Cp2GjZNjz7/M
h8FPF9+HIJCHsdU9urCaIWBC7pnzf/voT1U1SBN4+jLI7JZwJ9AP7/Le/nVlvibO05+dRSjSVJKK
EU3kzsClSmntYFsRR/wKqh8CE1MLj0aAXQ1YvkgzJylnBZsxU/n6pg2beIFtMnaBthuxCe0KfcpY
+e0ZUhsCRauVymWhPsKnRuNX2dMCZv4f65t6mIQ+iIN5R2+KBlZU6TSfIagyWkhkh/6vhiYvot8N
4vaIPttV1AK7c8rghqVaM80srreO5vyoGjeE0WdFI7s9m5l8dUs5m9DkhoBBVMmioHV0lCXfaGod
nhXr4Hf9xDNNbDQS/ItAwXbAii+bcyzrdbvYYTWpkPElfl5E8N7OX1fK1bCR8pvIdgUFwFS8eDcJ
5NuzpFk+retaVi7am4AU2GDIrCoMIGYTgwO3Fld/zmc9mZ+iYkOzNNdV+OUeQpUZjMJD8O9FvM2P
bzhFXBYtizDehkYqU21FnbEJpfZiQ8OIi0BJ+K9FnCP93hNsjDH4kKHluKgGMMsE4j8CU1cvEoga
JbrGRM31pVIc/HRNN/E+8oKj7Przy0DVqmD0O+LCDwLfClUTs1qlDkwW0/0oz4QHLEHn7vMDkQsd
RjZ/Xa2dQr/NBTNzu9zOWKIh1I6ZLeWaz5DcwD5JqQRwrBDVOKLVsSlPx4W8LjG0NIpEDVpLusgX
V9V6/Xv4ZiyMkHOeaVAxO5A913V3zWJ5wF/vHlp2IZb8UI/kjxcx5o+7U9sglaYO0LusZvCYCVeh
gzSscPAzEtP5YglyRgovwQv49YMo+4A6oHeBY6YUCcuJDMTezRJM8GQqyT16Xuwr7A6AvwpHP9oW
Z4f+5jgAWXIuxij+vO8bEloj5RKkx6UvUNcS5T1MOB8KDYltZllXjrDwd46f6KcnLgp/X+q+NwYX
LgnV7X6ZdQVSZ9MThkI6yy+8pqJrQnrqrJZXm+m+P5uy/RbocmuVdgfupSpciZ5vvOtvtmdUaU1r
cC7M/HU+KwFdQMAZgGnakfAYRzvcWIcdNhN/q254i7z7Td3MVOkfCqGaXc52d9QWjf8eKya1g01R
8jz193tj1TrHu2QCrkoEX5rwQt5p0ImXt45nKQpBzYXBUqw6aIDX+bJ3p/Xk0FEDfEUEnlcyC/tP
xewFrGtONxcV0iHYDs2ifcrGGgi6Lyw+YQNU+V7fLgjJ2bYXJgzIAez2AggY8e29REtHBvTuhg/8
FwROQ7nVMZrMQso0RJsFHXRAMRVGAaCFVOeIkw2HWYSgYslxfoXMQqvHOX5PF1BC8VaNqYbInP+P
j46YOWJryuW+eRZLsNlLZBQKVvrosHPvbiTi7NRPIK8ZOAx/Vd08U5x21/BX0Y2AdltyP6j1o5ui
xG+LOmGi1HwK3EEStuZ63iLV4zy0aZ6Mi+bP5CVbMx0kpxNT0NVrHhWhXZwX5HwcPzyc8s3QB6j4
mPCxsbuAUXkStA7oo5D8aQybcvAd2bAEO0/GRTkiikm/d9WxZvuC9TQ5EnaGdOd3rAsa2lAvOhup
alTRVh+CQA6fBeHqjw3GZTA8Zz+nDKVibOM2YVAric6+rRUUrxkbLQ1iWZ7V3qj+8ZljGKYGeuxo
aM/lB7gr2re0VgTZ4Fqt5NrRtxk28DFPzj/J0ehwsZVZHMDYz87GiBEbH0tFPGhKdmUP1mmdQRNM
OA/cMRqody188rRJD1USPbn/LbHCeNE2rFzS8IW5FQoGh5iu0KnxDIWe7R0vgZrFKNl5pp80PtrL
Aw8D8GuYlYFSkSXY7uq+OgVItAXqkBSosHpOGQ4OBL5rbdWqVzkOxIuUdfDv/FiSRiq7ysIoqcWj
v99cY/I4qCuWmjcQVpULioTMS2E+mGgvtvXHJk42VKd9tSgJy4VrjhryOg9tLfavS4CKKf/eW9fA
3I7BfWSgDrLPPE7Qbm3CxrRdiIOVLqxGgUkfxrrLun3gC1D6cM109Jc1XaMuAFRWN+u4iNUeM/fr
A1F2sBDjE8tnExQgHOkMVLq4RtYQy0KDBZuHz0gbMg/ArzjeqYYVK11wnwv0Pd1/O8RY/fOehIEW
BrKYIGiL9mSouWBtHhCHCdA4hkvpDR9m3pPAiOWq5emNnfYsBdL/lv3icm69nZodqcDfVCjm5Imo
OsLuAVaHLpibxMg3bSH2oAJJXNoKojy2e4CCfQ2rxrEAOwtpSmKc2oDbpeijIk8KRdXoKHrH2QbK
Y03bLJwpWzbN6uTTFg3uLCTaJ3/9FWzx7RhreX92/OuWuyb1soGJLVb2e6GrF26exufGxkevfijY
B/abjq9XFI/JW3cokdNGHzrOJRAXuM+CsGJQTv4GCUDe1cjNCZ3NOcusEjv424RJIajHye83eNpB
jHXzqRxI2zl01HS/GD4zhueItbJxxl3qrLJL5e0wBQC/hbmhO9ODsx/YpBN5kwP9N3CS6hBtG5jB
ZcQNQmTqMQtFosvrfbtA2PNTJArplq3L+QGwBR4Q4Q1Sw0GcPn2WPq5PYpdAgzLfdKo3vK7cwrZJ
k6yxAsoAgbWLAV4UQG8tze/M4UyqFykk/dI69cOO4TkFuu04t0OLZi0NISVw5rmXxdcp03ucpCue
zkdxencwEXGm8gk9tz1VdokjlpEew4NwWZYwKzbGkw98NBu8+l6XG1XojijDBW25LW76N2RiTwiD
BmNzQLOvZ3X8GN7Lyur/8C0kjPGjdxkf0WQPJVy3RluWFw36/tDSj2I9rEmjmFFxHV9PbtR4eXYV
qMLKa/8XMUeFnTGla8CcS9iq94jKKRrOTSC1Byzf1qFiND0YKjRbNNNWJaVDWopZOorJLO1QmP3r
BrSujEEjy0PKXnaxLRFsJPw/4Zy9/z0vqzOvZ6ferzowGSspCrbEub6n1C3fJJXxyRYYrYnSBfFV
u28gN2oQfl8ovU7tYOLOPa3E+iM4pY6M0HzK87nS5pAXPMadKu1op85TnTJ0mgwDyr+ZFx12AT0a
XgMW26UhwHxF9xbiO137ec3f1Vrvmvesv4TdNjNk3nN9gi9jq+RSPFBvKeW6wsr6BxgU3QGAHLgL
6Q7c7Lm6TSJE93uR2pMMLXi2HNP7gnEnpXLe97VpX82ocdz3YSbgy6tNg3fnu+ZqvyHaNMF4sf+L
7TQ/udW42+bPZzTMcl1HcEzjlXhOMAvLQqvQMgO2NBa9Zu1BeZ0VgR3jxZ0ztjyT+S/Ac/MWLA0t
kXuL6xb1GlCegdQtdnTem8dGPJmKrJd7/1K8+ZKoxxcrSwvmmxBB8HGx4zriPEcs2PyMyUDbfh8x
Og0bsp3AV+4kEayZ8RylfEOo1/KiVWHzywcpHMF+MF4iskHSHNsTqg5nEmQ1bCjWxxMjShEsAQLI
3YUAAYFaCXDBw17bDLTkyuTdPxYQF/GEG5uGC6QByKoYudnx0e8dVBVtmj9zJ1jlORYzttEt6PPF
tPOe3lDcHOkwcf91lZiOaLCi6OVhaKmMYVi2erKhcYLviekwRdqsKTUrRjSeplJ/flsMvkku9vaa
rAJo35MwYAF3twRl9pRkX8F2/NAyKexOAwmou4EXzY3czJFkcuKPR8RiwegDhdEjVRV+A7gdBz2F
oEWTrZ98NkRZIKw3eWBwMJO0YPoVg0EPkyv5bOmH1Uw2NKmqUwwppol0emk8Ugpe9JrNfWTWNpAj
bP3uaUVF1TM311m63n/hL+a8syoMHH+zWwscy86mkz3jJ94C4yqY8i22XoT6+s0XULH5xCH+Wg2j
YnJ1MFMZwDle/LGlvb3C1KNB+iKOZ59JqjWU1VAFJQYh8flGwwOByULY0z9jvPEwmcenyLXWSRZx
vcL/3aIuhd5Uixki6I6B6vSvwjqvJZMfxXYqLPsN+ZNcTFx3gCS9iQSinTstV8Kg17b+XveRsy2z
XZtQGzs8QO+TFhNdpxEDB8Gxb5jsge+huNeEcmU/MANh1l1NGMDYHbkiOfAwqB94cqSeCpLI0lnN
s8EH2C6le1DFZZqY+T6n0siHqrC5gnxoV9O5Y3AuOklSjyZh8f8BZDSZuTm4MZlQzgNoA++0AKRI
UvmmJPcCFZWgJ22hfcl1ATQZneJ4Bv8b6qb+lYxABXx7rL0hvJ2l8mKfyuDpE1vqpN/SBSJjySQf
SumhJQNkRPlbAJyqGKKBsVDxyMTIy+AmBZaAwi0YxVmMz4QyuUOJZmafy9OuHA8+U9NWQzc+7Qi7
/re8Gc85yXoKGNktj05jNR0HUvW83sDZPj1SpOxLvucvpEOWy7+lEODdD5huloMVJU7zWBPx7qJ8
bZaqQrAp/bkZk5Ffu4FXPPaq0gSHzpegTjDdDYK3+jAHRUGdrLwSsyQS/Skw4LM46U/fqbaLecbv
EiwEDGuJxmLKFnaHk8xA2ywQ5Ru64kjYogUFiJel0LpkkDT3jzi04KTtFq9ZzhmjeB4nJK1Bk2lw
sVQwTuFrM5pNMAXaORiHQpnFvkraV1lpngHSpn4r0tBOZWc4Fg9SkmcTmBpGlVAOgACPaiF/P6Z0
OU+pN0rGNtscJ9lAWba+rArBpv/sIqpC03/pNekipibsWKUvfvAo2re8IrnITPRIotM8R8JARKO4
U0xzA+XBsWaWqVDDkHkJR3cqppwe+YDAT/Wu0dx0nRN8e4t/rEsPfd6eThZXDWFi5LTgiIedPyP0
uoBVINzhmvdwG6nhFKdazng7exhtYUynattZmCu7xGtV1IMyZBit9Qwxr1zQmjvIwtQUJXnrfSA8
Fw+Krnc3MboR+2Uano1/ZZyX+f6Bt/PLGfQL8AFvdKgDSEmkB8ZZvzlTiYDrC+WqX4VCguug416c
HA9pdceYhJG2Wz0SOc+OHxMocEmf8bmCEgR10jxYHhGJfTIcrLVMtGrLohsLYeW7qovCmRK3kuKp
aHihkZVauzKY0m+Aj5xMIOVXs/SayaLNS0UnHfYNI8hOBCT8FAj3bhpRGzWu4RRC79IvAehpzFVX
pnJv6MtZNw7pT3PRoGtqc9fdAzd1jpyfWRRI9I0Kk8RKkfHrGRGsJzQjYAo0rf2WnvrIP0vh6K8f
cTntKdDI1sTUj6SShvE7bw2lHj7aLQsIRDgT+u2NderT+P6AIJzUEutrEju+XiJRoEnMsYxKiOcB
SaomFoiVP3NEcz1OP+FbQzvTa2jDQBEF7DgIvRTL90jVGqfJCmsr0ah/bcSloijYqtgPzHZJhYL8
gLxFvYcIK2f3fzAZtM8MItFAjfUNRU9k7MLEg0Z85UWxt+OsBALgGrG+Jl80UQSWxfNioyj2D4lm
sUfojALq9L0c6D9j6KelFEKdjCEkbBHI5gIV62KuuVi/4hDUqc629jV9za+4BDMrsa2tXcvrLuHW
nHMcLxYwXuUhVvT5hCvnz8lrAL9TPze2Em6+6E4BseVp/1qP0eghQoQf4/gUobVOGsuDaHoXBBON
kAAbjoZewWY4yOtlcAT5+QiyovWzXdxpEI8RfEE94c2s7hWDYiDwB2haDHomG4JKqeKEf1EYVait
OAQlzwPPYvCk1edzSajNbqyu0ARfq1Hz5xMUizmpZUpqG/Hz9njTaADqGWpX42QXBOrhzWQiv7V7
lPUlchDTczL6Y2eidT5KdCHNCE23ep2cenymXaPkBF3L0XnwpHNyvRbS+2qHCN0V6PxyQxPtbkv8
/RhWe6ed7sCjyM3ZXeSUx7yBFFSuxjWpX+hxUTeX6BPAvK3XaQF3Jyz59RDoXxBVjL8ey/+6kuY/
JA7k1xTfR/VwQGcnOiPgYgLWTq115qz75eo80gBAeNtMgFQhJB9fei4Kw/SuOj2TUm+nRhGnRbAK
BvTrvP6Ljl+cCVt5K5nrFcziP6PQaM1WRy4uJMqFEx7nNfDqO2rsjdAhOrCWIKN+gRuWWdQCgGsE
kXInGEIQmkMdxR75SORAW5akjXgcjUDwL3iwpQGCMEWkb5+5AvmRflmwBcz7K+wmRJcyg7s20AlU
CqybSNxITOWb8ZsY9j+xsUt8MD5Pr71XqmQCOe8xzy+9lvnOH6S6z2CSQhR8LpHCF9DdTws16nkF
t6Fs4FaTrL/U1bRNExzKrmGqJcQGdL1dTuneuEdbJnDCWl8tjMXnqn3h0Q42T6lMILKBbDJ0fAyb
1kKt6rEA3yY9rs9+ZIprMND3bklxBm9230kdcUqy/M+HwiwG9UVmWWVHVLlN1RUL32CECyNYmcdR
5a/B7G6a3Ue2s4CcKFqk/l1A4ID2lfFWtZZC78O0V4/8KINzMP5jNepTr0xmujzqoT9q30ThpN/C
dzsmT3fh2vu73ujtRBlUzGfjHHndF0mdOLBAFrrI/sTfGK0/XhSpk0vrrEfuv2jKbwNu0U4fk7tO
OofKAvWPac4yp5rqcnlx/F+yqxvXXy0dZImKvqRQRgsfLEdNnxBGiuUc5R7KCVYALCcNiPq8oWu7
eu1LDd8Vztc4o1EzNdQ+qs0W3RVFuNoZgmRxL7ogKQNz+H85MTuB97thOmPXvFe8YG+3c/UhrX06
bPVYHtXi3qPF8Zp2D2zMR7a2u6me7cGTEwzMtkOvarOu0j7RUEZlS3VFuBQX5ZCC2gQeT5tEHK4V
XLF48VInAeheAsvfyyLUZE6ja8/jnxC3i0bIqLRQYb26+uTh7MC6FcHY+W47mUlBQUnzfI6uv7Mi
+jVQb515J1nVly5RiVjdNcidYFGHhIJ2v1rfIGz5hUBJ9KdA0zgNusqO1iun9Fq67D2+F3aiNhVe
Djna6OZs+ttR16bYcYIqfvfbbOvl8A4j9z9kpiaZA8OHAD7q0NSw0Bf2R+s5WXWM0H5HP+g6bguF
EA70p34doUQ1rm3Q2ooaU3eXqJCYbLgE5SQ8DzsLPNiWHJWOVoYWY4qdc30TMDy+zw5G4/+A1hDH
sdCIRovbz2KqpOksnqjHkyxNzV6xQKUaDvlo6w2ItmDeXES3WwKDnZOalfd6T7rQXl7ltl2wdp/f
dNDsNlVMXF5Y0ZrtNhTuj5U8IFtc3EpGvF6N0vyZ1deRlC6iSE3a8m0/Hkuwixuet8RbZvmXrao1
iV8/w4iFaIVZxHTHJ7ZtHvh2PV/OlONF9hfwAvGs3SsWsh8hquo3HY1R427rujVWZ7iyPXJJcQE2
IagZlPk4aBtAUFyeN4tkKPHlK58D6DlSKnToPz5cadSkUQy017ik+Bc5y1rnpufvvwlzpIM6dsHE
s2eR4ypFatMfaJbo1xkWdwyOJxwooHg5fO/JbpEsSZ5goYk9KTWcRXIwy57PTLf9y8AfZVzJMsxw
MqtbZXcSPGJ3oX/216Fi57v+/8yGSFBtFPyOO8TCDy3QZ0fCiJxoJtDktbgpnhmlop+6taQpizr1
oBN+z1O5Bvty5/H6e/jNTM32IBC3jTB4o0whkmG6iOLy8LnxlPi1+rJky+4FIe7qh3z8zYSybWTo
DfczNkHLeVqAkY4Le9qo01wx0QDeOWuOi7uXfbgzpNHgycjBnK7X0e/F6bJkAbjS7Fe0grZsBjzg
Ccs+Oxp1KbEWS7F+VHJdMRQH+ZLK7RcMXSyNDUGKb3Mh/C6FHcy085pmT3/xiYMiuW2pJK6z7DhE
pXUZTpPiktJUgXU5KHxfntYCTY7ImOh/QVozM/x5n/wSXWf/8gKzalPNnmGh+Vj+CldnEzL+6WBx
9+FEMXXGuhgjpMSwjogxBhJEGVo3r6EhDOMn0WrzugTovxgJIx/2zmRRH8t/eQ60BtuX2zZPSOtu
3ZO4TcqRIXGGlT8QC18nIA/mGjLzpdAP1CA0f4f6Znc+3J0N4laEz/vB6pxQ5WKpT6/Y8rTDXg7n
LxBP2BOEKZUpbi0rG/F4RLCqHVZ2VMpZLaeJtruFnqX4dkoxzKGGNHBbIzJpArXXdMac3eb6LBqG
Ddnezmf6mgj9HczNNAJIo2LHQgU6WwhY5mGqGj4sNWX8dLPc36Jh+MVzawDm5zZFWx4IsHvKj0sV
+gpZ629WlKtxXWb6sLzUqtUZkJHLvzxHF7NBzTnh7iwDph6Zd2fZoymB/Kk3Nluoukq5TJPohVoU
LGJAHVJRqcOZYxMuUXlcGn8j44unrfjhI3TeT75SHe9wDzQbf39i/HhQmC6bmAtuRQkJ3D10iVg6
aVOs/ApnhqkMv52hNK2F0Kcj0kTpJbdAyW9fS3NSUJ/6l9oNL5Q9m4+GDUFrLGFWhoOioFbpjRpl
VRH1a2h0gzfy3TtW06smbCcaVT2Tp2EuMI2+XlIju1Dw23GDm8fn0dajamVlnC4MFUfeG/r1Zptb
fB/tD/6e+JP6b/qqLziM+QVR0LDnD6sV572U47iZHsaZKCwvmJMu0iejMinpWPUPMG4esRHVLxI1
FdXbffuC1X9TtMJtgph0McPp6TRb9u4mggF+llKAeJqp1idmYr7wWbdyQcCZeV7aM7pGNUgX9nim
SrwwyMr9x/dLABTsgvAbVAN+ZSvaQsSSv0cecXug4U0tj1dYm4RtpWy76F28YGmYJUN+KBIIrWtB
lMuDkDYJmx5BQn9gCdeadp56cHQS0mYvlFsyAz8v/mw8Xra2NrEdstIPE+BpWYu2HVflmYltlZWy
uV0wUxfGRbtBqoQe0vRU0Xk08C/olUdam3lg24V5eKfoMJ/3hciiJAKipoC8GnWm/9lxPBoTv8BL
XPhTyVKflwuv6BXDyx8JU1zei4f3tkKAsQzSbQFeqAvtSt9+atQ3oEFa/s1kxlwDC0ndb5d3HtiF
Soq6MY75j7FdnifRNMmOvhpg1biA8jbmrOCVG0qriUqYoQc3nTUnBk3BGdEkNx+/K801zzxq/OMS
J3rBI5qEw8Tru7nVoyx8c9xBW3B5xX8S4Ys5qSsJNCDHq8fIq9E8H3Txv4DhYptNzKfEujhE4yeB
MhmagAIZEUn/7/F5F/doA9PKURrZkPasgQx8eGagjncYiFGaa6RTWM581Y+63bp/wFf87dtwrtiP
sCzsiTHBzsiP+3zHSeLHv172w2UntyrwY5/mm4uKNMOTM8sRMnUFKiengSr+KTxo1HxB10YzIpWZ
tCuD8djgaVDYf5WejL1PzpBp+fvPE5gvZn6fEuD5ztYs/rez5i8c4zSFO54yKEfgV8sV+9BsVld3
vFOUlGZvc28Z7hfwAuaj8VCGakzxVHyRQT089LvYHfHvY+IZAzHrb+QMwjI2unqykSrwi4qmxgFr
raZ2yP7NLlxTSjjp5i2NMb08P1ogRvxupHPSFFRjNkPki73l4D3Jw7gLCWd4a/r6GbRuUYhzuWzS
wDuloVUSnQIs0pOIx9EscZ4mwhWuZo/26E4Fyo/anzNweFU4FZ6vXSEbkIAjBmSgovT/OrrIU/Es
A0m+Sun1yPQALsc1WZSQGJn2tgb2nG4S2IJCD3gbc9pFMZdDEEKVMzYxUPHMrtfajnsFyTOmjdpC
kBZSYMp4hwkTJdSqV35/ynMP6GIFOT0uLXHyZCfkS8YoABFmug9KTYtvIzdjKP11bFiT4QyNmQ+d
jQ/wCglGg17bT/605Aw+t0VTwjZfnrQwh9hPjd2id/gOHRl+S0H8t3ruDcz6ktnavX120wNv0CCz
3BmmEqgOfTUAOuJe7c/cCZK61PHEazMFrJdfdFfcEOXVvHv4LiLmZpDrlYEAkCSUOFcd1/iKGU+E
znH9bWArFvX5IoyM6ve6f2OA3yhpnK2NNPmIQLkss7lp+3DzCKR2EqahFc6K8y9j0Z00enOblpr0
czxtSXq3Kk/pHbH5sZ7rM5z+vM6u1e64LjDf3/UGSXo5PlXxOIH0EsEka5lwT+3FP+NN7M02oVJO
v1RA9zHlKWE1pMfCm0MxeE3rWGO+1DfTnhM4jwbYb1o7SxYg3ImQm8/Wf6qyfPKJLyVo+dFzPfq+
fNleR/FAGHIs06FU9vpfdi4Do7auHuCzqVT5ZAPqnHZNnb9rU/ikS4fyDV64CpU/uLrgHSo/JECr
9z9+uRMYXoiNt5dxc0Z9DGSKVRWIGtGoNNpsENJHu5L2ppzndWNiIQuEtMQcvzDCTzQ2cf/N/ayD
tLN4FnuITAIeGpmHptOvAJpeF1g3t1TOhtZkM5XwW5R5iIlDR1iOAJN81lMc9Y7cWIXQBgMsXY6y
g3vPnRcf3oST6wRD218s14igXTzZKsDmxjIi0WNbcORuwI0vrjbSERP8W31Xv+SAm9I+kT5Fb2kH
+Amu3LagicgVmYGbD8tJsCeJ11E/f5UGw4r7mL3IbOSVhvtOd32PQyBhaLU3DCZphmcZgnYL9c9W
5ZJWVnmPzFKp7p7V9Sg3cxRuqVlCOK1DCR9/8W0kqEF10dzutupvmRvXNuLvDUKlaZ8AYDClk5Y3
1yun05wvknAXmKZbYMhHVpRp18KpIgdwCUEASCVZMQgMe253JuR9sWLCmq8ICoDpSqbGOKfOorJp
GjPqFl2gizhU51Ds5L62f7RAf0m4XHz00ItgfJZZ56UEbp2zdm4YsWw+/ZsiG9z94p0KanrAqZNp
AYAN2QL30Z1XTrGp+7Pjncy8XzeBmkkbyknbzIv8in4kTaezDPH24eS6mXS/Go/hTkE0vVrsg1mk
1UuLVbAkjImsdj4oGEETjwZfvwP0P7/XouY/mPLADQQ1Vv83dgUmvnCCgfnp2upmKSW5et7flUOn
vv6MO1i7bd6WPk3/fOfOkFUcjMr4J95j0WZcgIehZ4Y0GaY8gezWsSYJtkdfhbdK/PH7xXuxxHGI
kAWF8UqvPs4DHvP1xBtxmCPRJDtyyHywc00QQggZmSzfYB4VfQKOT5lQx5UYOLrkqYZon2zrP+gt
eyaH1Ujc8WHzFLTvgCuPBNzTkpSNI4fw7e0Yo6De/aHFg9GLRtdHqJsfpk0XuzyaO8QO0Xjju+z1
AxPH1Qckesaf/a3U6ATlOS5Yy22YjR4TU13aZiKqkBGGpCv4GwK0KyETlK6zFX/mi+apjOt0BqCM
DvBUUu+LJVbhWtx/XmJrzwQ0h8e5x2qJeEKwIZG/2VEYNdkdLODh57xb4MWyhR1BzU/wBWTXezP2
mAsE7SXgUUGGH5EP2l3H6fP7HWNenlDuHfb0K8JOr7YNebOcUNlaKBeavI1L94Zx6gg+S+Cop9AT
jfK0mQIzHAnOsN6XT+ZluVDJTRp4bXU8PS+wwASignv9QdUj/cQINxkqCXSDHOCiJ2UsdGngliqA
QfHztoRK0vxEINQbW6xwrjUuCAhKsiuGhnd8esnfV9WSRo2eEomCc84ONh5+LI14VuAQylyke/mr
ucaUPX0/x9y4Gz3B+Od2lj8m4apR7jkzCoe8OPlrv4hGTjUeAytEvquelfFZhnF2pwj/EXnphFY5
9oMd50+OY5XcuxtcN5f2WtHs6T+SNdIEM9sL2/wy2MBQTZfPo57B7Q7JnPucIDX74ZQyGhSI1eC1
c7QKWe7g5Vu5/kopWuROSRX59lD0cW33SpuV8n/F3dH+nCThuaivhJvpx8ekUsShBnWmDfJ4w0Rf
batFHUF+ughEPdeahIcojilKYF8p8urBjm0xt3jB0h7ssJhepVAdhB6iFPmuyENMQiv8N4pOX/l4
ShXaPXSaumUV7kowgyxwoNaur2Lrj5nJD2rKL6i0tnrC37tpuTIlOFxzzktCAR4Xi7WHu2HCFOUW
v5acZqUkNLFOLqw6nzQagVol3KQ7+VLKQL5lneL4rP27vveC3BipfMfMRX3dXl1ReW6ZinVP/7hP
KuW/OjHQz/vOFHvdANpFu3W+wPoquw89pUOXID1SfsKvkv9wfzob0zfECGg54OwmFQ221q8CTkKf
xZ/xeRtC+8eRu7rI9wpFB3Q2e22a5lAD0LUk4y18B5XgsqC44lhidznSq7QlU/gWykksO8O/YfEI
gTqdgKf/4v2CdmN2k4G2fx/w39J80tkzpjgkGn6zMJM8EPE64nSAaFtl5r43fULfiv0ug7GSdzsm
dU7j0KcwO32joBnyvKvZncZc7JG3lJ7vcUDuJnUDg1Qa8UbQFcnHih44FvIDGuuu/8rvk3kYjkwO
+hEUNB7KYPlcoZciXjqY17631OMXJD4814/haOGPM7UFztHw0i21qhSUqRLeGUsSa42narRgbB12
EbMVDPep1dYMV8oEUaAiUYVpnJbrdrnpOkug2JwGrAum2hPwdY0PpMgdZebGOhJMEvDDCLgXZvVQ
M3XaaRuW5/B6KAGTSDtxuldP0Xh69R4fSX5JHuaEq6ijIY2iOkEEYvxBMfNT97pkIkZnafimY6rA
H+vEHllWZjmnjqmU9zYK4giyof09mxNOB/5oyl31pt4xp4/fbgIaMvLAjX2/gwRNbOI+XJvspVeR
oAomtf9RtRppRpc/ozsEbzE25pZxm8p9hPohy01lqgDGj0zeorbwPhA2gzdd8M/n2IRAReU0dW5Y
IhNQkkASGEZEV8nZa2e8lxkQDdZbGvzpsyERG4S/shOK1nGRxJidjfSwc6O9JgTfFo+tsnwETCfb
vNKWPcPKV2HOqJ/cKucSab6Wopzhi37jB1ORPqzb/mAZQlnwPPHGb8snt673y1bLOHNJgF3Jc4NB
GEUiAndfwtNdF44w327PGCrZ47C0y1FTu4WXbtgcDPmpsrW9Y2V7pC34v+VErIc2SXQXO+4I48au
z0TZ54jHX4El1u/lCxdbjH8mQDOipZUKeGCy0Ktqmn0QdZQ61Md84jT0/j5hBvthUvdwmxY7RNUN
/+yof+fgbasygS6xczUX83LXvR2VZwh8I6fcbRsjmleiQqhDH3jF0PjwX4LsXYJv0JTGIHQ/fjnk
T9LbsVmKvkfmMt9NwMjsU98ZE2sMPxb9ReNuxPvGU15v662gKc/UkxgFqUMz5/iKVTdNG5ak4Xte
07RrExY5I6Xit6mgdZkYuy3CEdbayLb5FdQpVz+rAFiBBXr2/rhsXavTULpTSCnW5UeaIm15fYHt
oY3oPQiEAwBsNiVN/T3sHm9cv5dVhTSMzsy+ZatQxeylN8G+BS8RL8YOzFzxd5CE9M8lHv6F60/+
PtlWZxnh5TNLUDqrftGyf5szw/DE/VtRtyJYOC5YYaD+m4ZCCeBxek1br/Y2QnLtvCUF6vaL96P/
fjRiwUaizS3BrRGikcXK+oYSaUwjMeuNwMWjjoMvLgeX+MdYrNEFexReX+hH4e1jp4LLSiFVfqhE
siShAkgZLjZv7n6pZBqAxkg1hW7iiQYp7VVkQdgvQYdU/gA/al5FfJMzhsnEYiz9pwmbeGZZlmBs
nLsuXIvhgseWZEbgPt3UazSh/GXiFJeCuAdSaCobqTCaISpPySSJBSFpQZBEHpswhRQCK7y7y9Z5
zbGsmXKCAjdxjUHsyIHZu3xCIdoZ7GLoZIMWmoAQ9q42rAYSVhf1QPj6sxUKjsSvBBvrZuUPN776
7EtK/OSu6V52urEg4qSXwOOo8UGKQ9njqJDjgTr5u6F5KiO2ghqyW65Be65lrNiwZhqDnCUXuRK6
MBoXfk7S7I1dH+ynjuWrzvhWDW7JoDLsub/qc3+se5NALonTaeWi275x18FxHbkUWpcLRRCCWXq1
Dh6uiYaVeWDkgy78aMfXQUWG1Rij3QbbNAOru5QmfSU6rFr0aCQU1I9xI5T+IzUiUilrtPZAiSW/
jB2+x3DWGfz8h0E5GY/3TOqyrRRJ7SREvBYgfvPv+v+kKiZs/QgXhPUr3dcNc34oMTsIqC3m88e0
qmPDUGH08a4j1Mu30HPtoyauAmh33s1PTgg8KyXfkyiHMnPCC4zf8CdcnRYteW1QQ0wCuQGaPdYz
eSnfADNIH2lxIDUsm8UQ1bq3RYOF/54nc0Dng7uE8D/Bu3cghtNOiHqQOW4Qkh9CAynAgc9x7L1M
UJC1qLNLlGK+yFzA3vhxLTq5SJjJbOoDKJK7GfY6ZGCYYWU4sdA3Y9V5s/BN+WcnlmLRCG4fGlZG
StiVdyIZGw9xo+YtMv7dma2ecFFj8wBqkr2eloXDqsXnSO5ujF0cpU+NoV2sI3uW2wu9hJntoXnZ
B+W/KvX2aO1s9LpQPHg3cPxUZkFTN+ugB5mmtC4uPBK7PAtFtrFKcGIUihlswBD06IlDDLiwitGz
eTd67EHY0IrRx8DEWV0RuweYEUM2vcUlkNJB1rT67mnJdpZRxZrSs18AH4SmaUWlvdcx8OtR3wTK
v8CrQ5kEOi2NgmlHHiZn8Eeeo2yNyr91atLdJptlMOKAcZH0lmIoUlqZjQHiWAaCGLpT3CAN3NdR
zgD7bFu/9nLXNzd8db2PpMt60mwb0e1go6VKg8Sc1STgnWao68mIJ4/eW0JWe7/7FAO+n0p651N1
GG/HFnFGBmvoEkYN54zIvfG62b819lplt1UQR1VxBI63a0YrbYOveorYAoI8Wteo4Swoc8L5EDg+
6/PVbwVFy6cjuqyUPK/bYgW3WZ/K9Q9imf64rZG7Z6rN5BaGRRYy6K4EGQIQixh2MLHknkqiOgZi
ME08pr4COrops89Wsn09fxqv7MFs5jjaKMso4aarr1bAGJMUXYVDTd7G1Xr9q3b/5d2pMmRrFYpS
KZVucKqyZ2u1QIjZ4dYFK5eQHeji6v2kLhDBXalxRW7YsUTGn4+XdA/Pk4EPg15mlk+QoWkvI5ld
Fgk4dFdm4xb8m13l7MGVOJW8PPoO3AoGPjRUEMz+28/aEPk5nC6VfVoHfaOv3QPuD1MOth7O295E
hNCzbdYrrwNEhH/H/mZeLsUsNTJWKATJuHpKv2IELrGkrhs7uq6BgM0AaAb8dq20jjz4Lq96s01Q
Q7mpowtSkfiXTiy7bwv8NzLoQ5yVBsXZ7i+vN89AdSCgmQ4xtzARHw5r0AKZDrUAAV1y5X4u1kNG
S7qlSxw+A5GSMtzd2mST9DI9Qoe+p4fuRrBPXuoQinU9dvhKbb4xZ7TdD5AHig8dTKmi0/4aIOGa
9G3zuaH2/hdy7sfxQLZEgLEW01TKs+U/QdGDz4Fqv8WaDPeNJlw2nDzUJDP5qOnGD3g+1UNq4m2i
/YKxb48ILcW4vdLGAGEqS96IFSjPvCtTtsf4PihMQE1Y81aKub345yiL/wjI7RkbrNx6A8zTmESX
s+Bp810LFNb1/RvYUCy882WcmuIT+PeFYUb6aq1XQt9w3WDMiu5KR1Na8vNOSQiiD3eWpnMt6KhN
wPc/gWjrtR/H/FRc3S6YmSkMrA+92WaqqfYoDIFgFKmND2SY7FKmtEzyWYZLzPQs0H43aZEkFJhJ
8pKX3yY9AqHicHDNQ1T2pXFw1MajUFskE/A661cp1yyqVRce9UeZ/t5i2u4ypWyx3XyQGdTkkXui
2QMTjY6EChAqOffpJVb7543mCbXhjlwt/7fdX7+ufzj5+emq/OaO6ek2FjsqHYVmHbkDsugbG3rP
LRo8oG7TBoXHg5mjHXsNGZE3cEaXyhaQJRyizJTps5O5vlSGgM0vEVgqEIrH2WYnWBM5RKv9ec9F
m67wVDeCddwuCu0B515RkW2BqeuwY3e7YC3sd2PDFOox0aepYLVUeGQ/ho870UfWFYPRYceh6gmb
FwONJyeD0/nriKMjNI5Updx2BgubxUqh+jufk72T3T0e8u4P6OjbMMmG00bykLhPzunh3tTm/++G
z3JfjRW6PNi2iwtsVgd13SyefaGVKHQQDwjsOEqzWHhk4qdW06DDsK7sNBe5CHV4ObokcDtQEick
SCaYcla4svLnG3x1C/UUjxrjVTPnz4+6ZK31/yBG6S7S1xJaGZurCzTffkM1mjt3JsDOPhKGkywJ
ElFkr7GidAlBP2CcxxHKbj+foB3YzyTwoQ0bZfmXNoPGAH4VAePHlSk4e28HawOjDWtD12hNR4oT
iuH4Ush9pzPrKt/W+3MwkoWvKHtKzfrNidOdS19A0F3TLdo5FM2SFcEqfMGTUJt5WXPice5itBuV
bdQ37bXTUSY2qRkgzdINaUFmh3ZWyHxPFDLnz8g2/D4g3lqqpMdmGFqh5tWHnR/T51Hsudjw6lgZ
b99vHQKI38o9j4Zjz1vUMWrVeMbuzbOjiB1umua1UojHK+zxxlWrtdOYQOz/uA5zSlTc+dGQAEkQ
Rr+kMy+td8FdLkKfWrzMoC6u2al6DBS00mNv1bkoqVPIV57jAVvfh1WAcM6hjaSeQIYSpSLt+Gm+
IVvNnWegJRGO4aij3/Tg3b1RrBqdAWF16BgddzInl/MD1XPNxSKm6oGzRNsNLHT6taed4EKSwUTT
EQdVgLcVwPbVzKwflp+JcCOcp20hjcMDvxP4IdlKpc8PzeJxR599HwAS3cl6JJRXOzbtTv3W+26H
+5h4GucEelsAPp2Yhm8Fss2LomjN3TrfC+mZFaQO2CqR4GLj+OOpMT9ud2RdYmv5hhkkMRX3LZGL
KFchFtfnjn7Bame0pp+KDgC/yTq1HWesTX+1DjdGatw+lVn3Qxc5KMrffbmFjqBHXntCLzeqkoAU
bEqPMrJ6ki/iKvDLjvCitlAmeZ5jNNrjQ5qQG1VezGQnOQL4aOoL23x0d1cDY3jFLS6uf1ZEbBhu
rxws6dt5LB7OWLu0AHkVu2BMsynjHJ2sZ34Qn/QDv/+LI+Be6rEgk6MnyYMELjtc76DPNG3X3yod
W4zf/JI6eyQkY+hpFD5Oz95DUt3SV+ronXdGD5byKqA95JwyUXphcIuybR2JEqutTcb6s8nyHOwU
FINZ8MIgSMiAuEBoPQBKY6EjMsImJKmAdrMUm+JzLVA22lfhdABwDnrmXjQIb9t3fcGNmkwrC0qV
uM0fPpB/E7h104vziA8v0S6VTdFpcXNeUPayNvWLnv+bZFMc467E/EdKYzGIscxG7y7l4QIwuBPX
JrnJbrY8BjCu5CheAH7QYxn1FyFQU1mAOMMMadRjIezcEaK5hgMkvVRHii0OpgXDBzyQiwdppQuk
DJsopw4a8Oju+9noE04Iv1RLDdRkEzBVZZrz2hacrvhSAohas7vGXfbMKWgOOi00VdbY1Li2NfI6
rOPQbLjXqnScGx9y4PjBCh6/hKE5yl3xg8xAdtAU9iML7dP/xIX4l82c2h9EjLeSlbp6PCJk3d/0
Pe2VOR8V9LaW+XwRNCx4b9GoqRVPapNT3xHQVDao0vs/0B1EHihqE+FuZph8UEh7i36/m+knghmD
H8NyN/FuPdc3NUnUmGgsuVRNObx5lTWXNxNsaVEX6xubLUbk643uMdLoHpGSy8oNGhAMbo36mBWP
YmBwoCwnSdQ3pVyZSAX4S4IpE1ma1d1ZLFi0mz5BuXSI08SXp6iSGAzos9oKP6k6R78AlH7+kl/Z
Uk5rta44oTzvWgGOoLfxBfLlv7socV5F01AkPSqIOU2jI7VhMhftSCqAXJ34mqbhoVdavZIz5NTJ
rrN3wNUVWbr7iyuya50Ps5FmEr6i9FM72eMoeCcs8yIGCtMKJaeZGxCyWmTTan1Vs0bwXn/vznQZ
kCj7S2XvJ9OlNNWoAPLN8RJ9nRMS5QovldoDJHfJYhmUWti8q7AuWf1GjAPMmKaU+tQpUQvNr/Fx
MCjdJ+UNlmIzTT1rr8NxZpQmMliKH9ygJtXv40vtUni29Jtm6MiCwHpy3WjFnZxf0+aE3MxO2Tqn
8+gQ+D41NQCTtmETMRJA994d6RkqEpVLS7Q3p63fGqGOjp1+G726lyBS5KdUkSQ/NtVIGZlzBOzc
3ramiE856SwDCcHEOsESaxyrcHfvY13OktfZTqBob9kaG0PVNhcERI5G5lTFKxJQYC8vrHcKJQbi
GdcaxYco4FcAuegD3JGSiYvauOTgnn/zEZ0S+iwnKPjt57oqALNzL7tJ5KP9dLL4+vL4ous1L/Py
qvOqAvGoI9zm2x02Vsg/+SYzhmFvbSSp0NLsM4XtjlQOAlzhF9MkR+9w/EHwmUwUz2K3uV+4oKOO
YcZXa4gVSJITaJIxYrsMfAbwVuwxFz/rNcVkd1SaJFc8wR2RfuR8RjYocIFBFJe4v+N2zTiTPdsF
bkOyuBreDFyXyOuGjfPuHEXs0Ee3wn8geMxijoxX71shB0zjr0JtwHl1gdQ/GrlVea5xWM/WiJ8G
bAd7gB3xQRXLkwYgEtqR/hHPsB9cNBlYRZJRV1PP+WICQQ0PT1bJUqfr8J/7MRTKKle83jxwyYKp
Iw4DQezEePk2DQiev1hhwVfZsK9HcE/TrBd18ZnQuOFcFeNITiKSTR0JuB99bOO9mkJ7Z2ISDk+V
MW9xB3tW+gipenciLZKJcQ8fKeLPryCD8lbjTZppkiEJXKoqKmFsCIXWrINxD9mE/pian5CHWQ2C
IbBGmRE6Xtf798J9sAGmygKlVtuGTsQUkIzsid82WKTLBGFfL28E60mLc07Wca2M0Y+OJ+wzUE5G
As4jOzZmADhWn8hr1rCi1PqVieNL3gUT7Mw5QwKvcHw/GLhku3iXYW0DgPDiVx3XXk+GhEW+JT67
/Kjc4GSGYMI1zdRpCTnR621/vHOuwfcAFnon+4mhx3R9qHMs5QI9kplFIBnCBbAnd0vPmMbo6BbQ
g2DVM15cM4BqlRZVvNxI7GXdDjtZuOs6CMUjrzAy5PprG2v+6u5bdPigQb8XCg3J3t9TTjrv979m
lwtfwiweiSpSmV3wtA6GhZD5RJv24X/t6V6varEgyvDVNs56FgaFiGeIFiRPxtC08Ss10M1ykrga
TUzABuSWv5geE94rrIfCgIZPefD0oSqlqK8cw790hUqKynVPK8n/8uziVcWEcRbGwB6wwXiNZaau
F//C1eijwjncCeUEqOygiUx/2rNXhowzRXDbuBHliwkeslhDhkpCLZrHKOR1dXXN5D/2opBNi7zY
zHsLrSkqnEvyeQ40lrPTOMOhX+64gZOGWMvR0rtxT4Z3sTQgqKZ/DbhIWK07mh6m4atU0VRgFAEi
D/eMBgXfp2mqexjmZegKfDnfY0y34F92TNCZ30NgeN0MmN5/kYXyoocH7VX4vSb4NPMxpX3eGqtX
EKXzW2Npl05R0XlTvFqGY0tVhhZYcu6w9gWxykPn2e5KTvEVC4SsfEy6zZLnf/bksVz2vmn4/TOp
5Lu4lm6mUv1AetnSW0FMAdbuwCQkNNeksx80XxMraB+ULmLhSR/goQiTzhfkvKgSXv3te9BChFLZ
fvrL6IjDiYL41jt5rbbJsAlECnOZ1wps8eWSe01j9/268/vWwpdken1FxeToTx49P9VMRSwB2IN8
ujPxe6nn2goOTXqQbY9lMvKQXuqXaoWyTym0cF56xjI3Ds/X8Ra0didps2nbOxUWo60jJiehCBSH
nk9fxFxcM91/0arbw7SlsmcSn3s4jowZx+oTFsLPBPL8wOdURXjFLg1vmeEbVazabpWdLEHETAgM
xEHDPxZgkkzqGtHGY/JRE1i6o8XzDNUgJfP0Ma/eHoxcHNt6oZ+TIsNtNsnYiLFzMZHyWuPpB+Mj
MCb8izz9h1wFqW6eSEjgC2jL/9cQXSXvGMkT2WY38BDMTBucx6bHbXoVW5Krc55YaD/nSo4+gk5k
KwdI4ONhDfpvE4hx77Iit6pBCA4O+k6OKvvO96Tp4AmIZukTATtUWBjS6ewsQWbTAptGi7iZe6FN
f3hR7L9EyPQPik4NEe+41B7c2i79wxvwqdFok6z3aVyuVZ8u250Jlyy7UQPZvFIpJoF7fYaSvm80
SpxdKcsUpgZbmdNxDsLU9nyqhe4toE4ucJg4P9ziWue4fjwiyelHT+ssYvy/KSCTnk59izKGccDr
YpgPmc8E/5/Y3yWosTi1bia7OV1B/dEJUf/JQhYKQ/t7R+aS//qvke5iFoLJKMNExuusotrYPwk8
fmlbQNfomQrUJ04fiRimVkDjMMnPZLPhaZC8d/YVb9ACpZ1Houf5jlQv2k12/8iXaJd/xdZaJTZG
pjVGwUxvw6WsdlQczd5FJX6sof85MjbRunS8zOAC+o3Koy4ZJD/pvjqfgJivW5zlcgAsRlq/9fzF
JfHYgBp52gvP9MENAU6HEYTEA7fruG+ES+1TIkQv/9UPJhwsvno5N/iHzJutLXG1cZuTrliNUJP7
GvNIDCT05G74hbGEQziS4H6MICUoFhwLdIVfFGFB78qIKUhXWbvQ74ybbYj6RbQZdar528ajKQ2C
Ejeja8fhlnlKhBVRwetZ6yJUgqzwFeH1pX4v37yrSSjXw0xmLP1CuKegBgI3HZY1UTq4P3YWJ+tE
8CqvMW71vpjbebIRg9Pt+zKE1A14FtWUOYH/q2R+s8V55AmKppLMey0lUjhmTnaxQ6HrQI5zEaCS
cNs1LW5WYnFQ0v/jXnri3C6iYn6b2w6D5RHrv3orqKTTxQGkhzb55o/mnI1j4ru6t2M2nl7ysOek
yuuXiwo7w/Bdp+2YOyFnDFFJYDUFcGf4tLsB5EeV5Hj7+lQv6wb9pzsn4rW7drBBh/QJnLBiBxg8
iaErWkj83VRguMIfFKk8JJGqndTA8elB1P2Dj7eFatARvALAl+4WlGYzJDcORITvYl6MAQVSR2Rb
zFRRDLpxSlGiPXSppIz/YGgNJowagCjGd92thSP7IrkSh1ptswfiqyxfW3W0l5AMen0c4NCirBFp
pZw8Zbce6rGJsOPyunsfUGJmFcPCB9M4bmxjyetd/iWptsGG5EwilBiUEjRWXf1yXsbhqlUf1LdF
1Olj7PeeZFOlui8eKJD2w7C+Z58J5q0RBX34aqeNxjuR7E2XImEdVQXR1vdb/qcZ0LkUDCAi6nKv
HnXadAHf1A0+HUD3e6AubIIlsLqO3d4BqPfVe3nUSyaq54Uf+RXZ7FX0ZH1dXsItIKojJmGA6k4N
0XjFg9bvkHx2ZiaH+iN49g/yyXvjQIbviFzkV0a8ud+kf5mTdRfcBPgJRb1bIUMQDD+obebYBnJd
yhJdM0N4vt4uJLRQwJ2zkJ9iVFn6PNGdzqQWTJpRUz84UoF06D0v1d/ioGcc2MwBrZ44D1FRD2cr
unb9uvzQAoZsge/DMU53gAapAvNjVy5Rd+SqeLxsOlpo14RqFtABV0YyGkEVLXqQklBaBd4jjjOr
Lv058mKVsznFmycKPCK+8dauxQVZnIK+NdziYv4z2IvRfZQgO5bDzHQd8Kkgbz/N+XEliqj1vzJS
A/HTpll681cRzMkKTLMzNilbM/9EzsBL2B3k4aU+cncb96VF0Q9V00PLyBnTM0LcQXc0o0bfrCdC
8eKp7wRfSWmtjgEHbPKnPbZBiuxZnthgfPmz2X3IInsuxtp3+NKY1Tg8gOZmNRU6435SkU0Gpflv
yvpPZq/KYZjH6QMIhwf8/R0U8ae/bVMy0dLiGpdsoupFNveQSgI1J5oM/8c13nrvRTm0XTVS/wit
kKSekQ8ZAJuc3vsmaPAkd9ku08QS11Vfe6GUXnYgqqprNQDyOWELlRHg9VvdzESe92mGeBkINLAx
Qj3KF4cP6UeJsSxq/3TDm2+yv8IHaOAjf02XtcgLnAG56+TtnMBjCuUT1hzv5+l6GntX2OXdmzi+
Wz5nqdRyTmmAP/6TmgdfJPfFgNTMVfaRyx/52beOR9XpVVnTKbFGdPmCWso2tRZY430ZxJDK6Jjw
6s63bx0xoZZ7DEP212vpfdPLO9bRPpNGV/kTzS9gqs0LVPRQgd8Gzjr8MGsjtzgLwK2o8gG/tF00
+hgRiPuKWl6JAtiP9eQlAOuCnr2RGM9aYfV1cPGTO/HYkoeUIg4FPCsKaA6JpAZ/1hx5AGB3Gx+P
zRet0lS9HT/oaIcGxh2nhE1WqT5zvnbdJg47wfpfkqM3V+lSPAtqCMmJT9XZZyuGE3QVdxP3JUcX
xn5zNpxXTKlA2uV+5Y2IfltddiPd2coYWE7WmUy8etWnj0FKvA6hSpcFH03+QjdJLRyuqSclt1+E
6TgZH3g/jehHEJQqRcQhHtvC0a5k+LEWm8ppNhRjuto+SVjRyVDnyiLHU9zYhhbYrLCgpc4G5yrI
2FSivd4la/n7ZtJ2X9KMQDfw2OKjXyGenXcdKhHbH2tHAgUX5ptnh1lxFFGvw4qGGxpd1qCtLgFf
Ce4TWwJ7raq/GgXotqiIceb6D1nX7XuwnPpMHDoSlcfsKhTvzL/RXdC6toLCQnauNxdGGXE9rwtV
gYn3UCGtvRkmf01nCUIOq0v+WIyqMjfgupKsK10fIAkAFF6OHX+tSYY6YsCRuDA/mgfe32WI+FeY
P6vKflB8VFEsQXJAahqlMA0o6LWh33WtH/yV216+23DY/obYXlrrkfPGNW8hfWir+uDg5+Sn6oKX
ciz0pv+Z6cCiFtS3wGZLMMr7Yv2rxV0qU2mWyJ1Zk6MREo3ARJ77cxQacMBPAgBQmINJn10wCmsm
XMJItqOaLocj613elXAnlZZLB9Oc8H9kFsbkbAQT3iHGTAJGEFPv6+MR1hFItk5upIFgELywsmsK
+GdCeQW2Dmd3hTFOk7buj+PhJXzB3NCIzthy74vjNpXireTBNNkMPi31qU/bEyA9KNBq0LZVcXvh
G//jiVS9dTPibGR4kMCNsmQJSEynHt70KN7xPhZzTkJIkCcjk2l4eqvDS4NVpPOBSUBSqm+W+Trd
BmP/GmMisdVQ+KKIgUbR6mYPRfmTMfumzAoUAFk7w1romGHt4n+jSxnnyd1NoDUOrxCaMbmda7Bn
QmaMTbOnVX2NZzOf4rdYm7BToh8VxHdo88iijkJJKdUQxYTvaK+CAer7Z/wZd8sOxvVkedLw3loF
13e3vcBl2b+RHSHU/j7KblU73s90EjWVAzLkotI5wQuw/tlQaZ1y2iutFjsrfE0ezeTO2B+1/eLz
g86Um7Nllz7GPDD+zNHi8E5vByGVCO9aJ3HQv6nyelQ9tG9W7hIW6A033mjHuQ1ooOoC5PuK91Ru
dZAYbZC1AxcIpb7qIH3GIWm6KOtXvbuSGAuG08iTcIx/+K+ZkMONzkuM6CwGWVD9qXAU2NHvnGMD
wOYonml2q8T9Y3lnDLUHLdcLEKl3YTMXaJLwdtO4EU0MKU9XePu47c14s99GwQZrx0uihD03NYO6
x69bHNcEwWOhiWjRZQgw7Lp1Sxtt66h5Mx+p1SBZmkhj/bE7XrGk8Pw9bGbX51tnUc7ztXheGtBZ
HHn6i39KbxasWztwZY7Ktk7m9NFvpECjGf6jGtmPHx+lKgN1ucJDMv5ft2Jz+Ur7tG2kdV12P/eQ
ZPQHQwaWgGDhapeHSpx4td3CcFbbBpV6pGAw3fXRF10zbSm34NjHm+nFnwFFus7R5SzkaaenGM7n
s9eS77j1eOwUD3SbmopiVxTZJAlmwgD0wDpKzhsuVPNY+k7ZkY+3qN/PfNozmN/lDTbtp4k98mmW
eWS5dlS1qA60XOY80kQo+ZJLz2ub9JnoShE35hCdOMEI/qi+HkJ8b2DS62So+jI1uh5oyLnhY6Fa
WCiDZ+OqDTLhm/A4eZOZpkg7z3Mkuwweeo3djmEIG+nk/rpXvyC/byIwPSLvbIUCpMLLmc2oug/b
55/LMahtOdAhVMJbNFyFvSTjgslxu7Pt9ATtMCsQfLdCLhcId1x0Z45vGnwdXrwSjM7Y6z4RD06q
PkI9oAUdXAbSHjc23H5kkj0awkJvWR8Xm7USoSgIaF82iWrOyxbOywlzoBflVUnXPFzFlQDdL43P
juwUMmb6qJeYcdSQkduKlFijGjrSe2i5I6abO7aQIuw566Q4ZJgRAchZ8CfAPDTPTQDwYnCjbYvQ
HEFYHfz98v1OfP0z4E/daBWFCs6rk2+bmeNehAvaf3jWm0kRXhpfceTlVmADlD5pzpcLpFLXyeel
s/ypxrATdzzQAVvVrXsX7HicLFbhvdr4tpXWmL6Sz8BXxjU1SQBfbfVjp2AtCfU5zlfB6qcAcnBj
M0+x+DR8qqj4UICKW5c/D/zlsJsWJG+TTdmTOnKRbeiD/jina7cXbCyM59VBbY8AjShXCbiSEHcC
EAczZo3ug/e92k744X9lQ+aHNh14Gam3hKynWIXOpDhjEoe23VM6k2haopDNRC8eF0ChPs/0jKT3
S64KPDadLS59FDZRcEz9JcsnyBgY6cm5cIoRhQR8kCaMDrplUpkQDLj3ddgrGetelUlnE6gUo5T+
KTDNlMcEdUVB8F2hCwvoGc0dZ9T+7QhCKCf4DpIdrzzvcosiLzMYJ/sTNPI/F//gHZwn+mFLZhqe
ZMODzcoPqmKN1kbJU6Fvf1stFFwAg9F6rP96ztcARWxabJhz6+MNo1cRsauZkgBL0FgCvNUTNksg
L2ihbj3MoW20QrySg6nigxPDQmlDoCX1C5QPAoazk4tOH+c9oOcQhBqYc34Oj6TYO/vNNbDnqHv7
90XEOE/cduiBaaEGS/2RrHpb5lFEG4C/8OUZE/+RWZX7Gy6QU8DePokQmKYeg3WtbgLxff+uE6P9
tJnvatP+FZjgQnx3RNFLw6QWHRQwVOFt5gVJCGD36Hg6hQPBwhI3ce7RDZnO/SH9XRsa4Fba5vVb
1DBBR+iOJPfB/KVLYF71dJ1qKXLcvSwmog+OuIPLVkHxDi3sdU7/VyIP3Bv2unDbTsWWod5+XJhq
3T84Ho4TAT01GaQmm9S2cZbdMbgxSKqJ4r7AhFC+phnpQfZVlIuvxlPgw7LBVls6DofWtZebDh9w
HbvSLmpMOt29cAPyYqo70MaF25rpt8YOixG5FrcR8bEg8nrGZ8hB+huXax0RZxDG4m6HWOPf1zZF
NplSQ2olHfFJT1+HJb0KftcVG8zMu+cA5uuWWCRJaEz6aOEeWe32vL6zQ8w27W7TGjqD2cTbOtgh
5Zx3TNPEgy6gVXPObJCimr5gptaVZqlo60qeOXi1mqdhYZTS8FdQIAdtzqgGmfpDKPK42ZpOF+37
PB1OAw7ZYlMj1Rx5SZP+m3qe9gzCdReqf2kQT0DUwDxkAaZJ6xYBvqwkyl5IcNMFqIkuGpfBUBqi
lalcsZFMFbv9fPCBiWH1L9H7rHn5gnYV6iPXi+ud5uimDkpd40MgIB57Y+aD6IimjIGzbch7l3lx
c73Isx5g8P3BSuZEkPUrWjCvAxOcb5JUkAPx03zzZoBnCR/ZLn7AAR4LYw9PAoRZwMWHTS7Kllj+
mZdWfIv0JwgHbTMZdTg6VV21wHiRZDtec8puqIlH+0eQCF4Ik/7hFx88OUJEjZLXUzMiCCwLeaUd
8delis6HtX1O4nLW+S+I+cBbXHvcgpjZ03O/g3MtOPvTVCIZd7lTODmxmloVbJIDJlvsxnhjYL56
2fWzmoZ63rgVev8KPKO3Dd9Y11LNWlWOcNGZ2eIfQE1Gh/xJx9uWPWMr96OkmQmyUo2HQSnxlcPO
8iafCA+RAzNh73gBxKM0hUxqOGyohU5wl1zkOR0MLDruaxYPjRytZRWYBBIyry6HXpHmi9lDwRzw
/9wfZ2sr+O4K7QAoP80cDUqAYKXfHimILiHqk1+fzRscoERofis+x9nHtHCxJx2pnTd/G2jmpJrl
IDXInnvvvawrQEjCue1B4NJOUFe4Xfte0XrGK3tJw/HWHQ/pAnlkUoG9trmjj5V9YojtQzx0A8gu
suepiq4wAJKLHMxhNC8XstTlFdLdrRhWOIr26txNXCZH5NaUZSe+C22mtP3dryelXI2/jq4uGCU+
7gWUycPSfIf4oLdXbFFOlr2rL4HclXwQ7+4NIVpGB1E9ATPH7qqRenBiw3OG09Eppw/FaR30Dfcm
f7qAzKZ7nHaOFZOtdQIygu6doCgNS7lAtCu2aJ18TQYGdS5297w64MIVBITCEB2ko472Ad8rfM4P
ENoqFMnZcrieba1omD9uSb2+yN4DDRDUrLdyzXBfnr2WL1WJZDVbr6+epq9KIJsu3yOzj++4MdNs
NlcraQpY3P+OW4Uqp3BGKtwaAcJVd9M0D2U+uBcomSqNzhbMFdEf1mQ3CsFsCyB7d1IEpQPLX647
rPE5mrxcoUtAIoGQ5Thj+P3U8ZP+B9iaQvdgPjenUdgjBknVGT4apaLnshyH8bhSafrLF43goaZe
HpKd8hIskoZVrADMY6rcCFU91ho3iB0e/votSKfdjI3tA34rPaPestm44YsyRjpr++Cshjv6tpTi
9JHsgCGV8R3UuwDolOp3m1UKiEAPDLk6bIrk9PuPFdZR07Opd48DkTOrRcxLjBJvWz3ab58O/Eb4
rZ8bTAX5HhgKKsaGAEvsEwDMRpP34QHsDA5cbTxrS7LJRjVS3dn7mkb6XT9PymdkjHQeM/kR+wF0
+nI/Krt5CUHkkEhRk+s2FAVbRjg6Yucv9M6DS+NawD/VWmswrRRTe0jUAow7+3Cg7bzWF+GIXG4R
vL6VkPrz+FA5nAblrfm9Gj8Fi+6693ZsrIV7E7EoAhuqP+dc7JwwscMuWbHyr3t01sZpEcaRnQZt
eghVoI76/gw+zzGLvCtsiUlgtHIXceOA6lyYtLvjYM10srn/1BpT4WTjGEMCSS/zPx4b/Jo58qHv
Cj9PXTSJcyC/n4fyTYi3f6I888m5WL8Fo3jkw+31LpQl5bvfeHvNgvtlheGfHCzLRef9Hav3O21d
dADsXN3t/Qw8GyEL/FYqiVEd3G3e2jTbRz8GxVVAOys5B5PayNu+WGvmmhPE7Hgb9DzmdT0Panag
dkMmYYhmyza67mq2cAsyQ+GrEc19T6TvDRO/dLiO8gOchXyZtuWEjJWrI0Eut3DgorMb6lE7jnrS
Tt7C2AmnVpBFvwFNGHvSAmzcGjY2yIP3AW6mYyBWG9K9nPZiDKeqdtlYagZeSlmIKqLGSJW5xOIg
ar/jFND7hNihkvhvtc5juTkbJv8HOpcAWnjmbN7n7uYi5uFZrwDnV6XQHQAe3JTpc4ionLy2ZkkX
xD64hP8Gq+mJfc6epqLWC8P9xpZNOwhoXRE4vsPQFRjYRtDC6qTl5MY+qEttR6kAXYadwzZ6YR26
B8TDcLeIrzZTSBh//kO/feYh81TSeuqjiq5tORE/z19S3McK2fEHjoBDzFagPYCTkdt+r+Rtbrxs
QEyH50+ZZ3rmqoK8e7c9HbuCr0ivEILEcCV1ZzCR5x/7Qd5UlQ6thgV6Li87pv8ag1re1p+LVPyd
AtosvAhqoePJhbS18Y5+mA7HBxwvcDWOkPP0PcH9Hp+9x2gYXOoPZqb5d4aEOFnswUXP2AByaKrg
396wQ/CcKZ5ldMo7I+sXekLjftxpTJpuNPUfY6hesHKp+l5AKUTmWNo4NBXWw0qIfMNqLTZnkGIF
V6SZEst1Wqzu5zx35nKj5OGUH0E0OLsypTCzPzj6HrPGEFmKOG2BMhWnhDCeEqt/J15mUJeOmHyw
UTIBlAWPSFxqqPkpUnz9pF/N0h1ZhLeX0MJprxw5RAhgM/C+9GW8RGJnj8++0OvE7W71sNbZ4vv5
kUtAvhi8y3N6mO50u43NZB7lKFmllgeUjvSpS7+DE0qGispSLS6SxpjHUkkVvJvo74n3Kfn+p6Pg
GXNv30h5q9O1c2tQoAYPaGZzUOXE9YYgk4VSvJsMpu8u1qmHR+jG/Gq8/emX02BOpol1DpQLTT+z
l86LbbOspP01OxdZWNxPodsEmUobMWzGKc3iUgdE1WWzk0D3vz9UOQwgVlePKhdlQ6mhIUrjl1aZ
5AIF0gnL41KGTjGqGuOWpQxLfZer6c62djJV/QQxfEgaYquHC+x2G2fHfuspQqNy5Vh8VRAKAK/u
IWtVogiLpKePLHzPmEqnX3nTj32jJaIvWtFcj2Q0UFY6nkI3HMV0herwYHDJ+EcWCmDWgWz2uzTJ
wwlVwzuIqrHCKf+G20O7GpoG+WnrLqJGDqyiD8B4pKAeG01yn9ct3o851PRJbQiHahevd9DIze/C
QzCt+uXnNWfliEn+uxnj2aDML/7BnZiGnSosiGNiyZtFwsBxkAqtbH89wKHB7Cr8lhhjegWNyDnn
6RLOOA56yrFlcaxTI5pmF4XcrabcKy05pYWvTdx/ttX+iO4utHAnmuFfN+0+VLuT79+FodAhhRo2
BBW3bF5efj64UKsCZh13ti9pgPZFpO8IGvrRT6LKqqCTGvtgHtWkwsEyiWgCg8xjalVoAkKLhoJp
Bdjx6mMGnIMjHHJfUsAKHFkpFDWA1mVbj1L3N45rdZnYqTAz4wLvie5hI82ccf1Dp6iegXeVb1Eh
TO6oyt4nnHg2gsAh6oRyC9JU+oe7OtAewMTeKk6BFdUAtn9rdJXCXwHFBAJ5GhJE/rBE8MGMDhKp
9gWs2/snu4xTNXYpxbbB4DJHTfuDCpKntk09IwbfhghltC3DrAvoE6NQ2w9W29wTNmBXZhSK+t42
xvMDtgIin7l0UyLNf0zJM6sgh0oW/jUrP3RoVTVfuOjkOaH2ecFq/HGw/hWA7pATAUcQ8lzkgEvS
dA1kAE6Ha4+pfeniAgFB0cZ0/66dEflaF1H+aYVal6b5IGtvdigDXNFJS5p99jjDas+wg29BePah
JN0xXm3dtx0Wrog3kh7iDtPpFvEt9MkN/KeGT/lMnnrQR0P1Kn0NAU2CGeCs/ZQ6LNh74tGONiBz
zXmCWiYoz1v5znt/ninFNHAspfo4ONvKkhtOfhJixjfBogACuHDCRHNum7gTI02EUrSi32RwmW+F
Hytu/6v69T3/G63yFxaGmlgxbxQOeCKvX3pD829YIT1btNFdAzzWsO+TWce46zLKTDDbpet1oINo
svPgRZTm7gevFpXlpx948YcNMEupZD+TMiVIm1V8LNdNwb68Rq158aKQzz+oGJltgsH646wBZ4ZQ
QEXAlhDLE0ukiDlYeHFN3eW0Oe12bp3XgoTyExlpTalpJstjUdsjeYr0V5zhdAi4tuQJxbAtunH0
d0d8pkVKm+yObu1aBvd95qHq39CqjDzkGfzJWr6taOooSjLFL+DNT90cW2aJczt79a40cfsFCT+F
kCoxfFJEcBpLI0CIt6UKcj9+bECJzse1XMm+EBofizA18fa/GdZ11/Yr/zXhsHmreUIOJFwGHJ9e
BtkgH7EorUw/aHLeSTlo+oqzWn8IqsmIQLTgpX874Fde9ourqA0n2PyBYazxWjdqZp5h/EWm2Bd2
WqavBJLbMvZCMWWsFp1kHpPZ4GydyagMVnGUJ3YmA91fMchOe+tYoAYxmk11icXVrnXY53xCNCzi
f+8jtGizcyI4kbdTUWnMZpz7/iW/FfCiUpmuaitMZBt924LzcIPqIeQiojcgHtqipW87qqvudzWI
M0ZMd9TS93jdbHSYzS59ZnAyQbPx24Rd85f7jWcYV+HPh1C8kEGKa4o+hiShRGMEdPt/GUFTtbNT
+r4Bx2ljLnW9eIYWYOjonHIKlwi8EuqUY1Qm1UwlRLC0w10tvaPOU0zcd9Lw0vwi0MUuMbcgIKTp
MYQceVZvo9DPPK97Z5f/u2dQtuG1CZXydPq0zStQ25X7r69KATvxqlZWl5d/Fpa217AEZxjCqokp
2bDD9u5JoIndiM0dvvPIzVaoPklK2N4+35zbfK/hvPHwo1AQwFRZsisIlwrgrmDsmUzLfNrvEw1g
QFZS4fifpcmrFgCU66boyPHe6BKvyUPI7XpWBumOa6ivZU9HlnS87folunSCC1KsyPM30ZQCMasW
cIoOCUS+cq1mmarEoY2Lw6YjZA+TpyN66mSuPnhJavzqN58QMpMdh4+FtJW4qcXe/Db71+vObPHE
QhOhr4B8+s187EKEBuQhtzBfJavYS8p0bk1vTaUp/7DNp9Iu4yWkn6QahILE8AHVt0mjQ7dSCZTT
GsAyWA5WDFOezmoFMdxpvipHBaTq+PxOsqH4Q1XXgdcFav+xIRXTZ2aaGb5ymow5Vi4aiW/3Whyy
l9qgPgJl7vEgfJwBkkbOGdJjfdpjGm1fNukMPyQpq8MVtmdWGzD3wC4AsXdBnkiBr6Ub7QTydES2
XJMnIjf0izDK5aIp7dQOlG+rKJmbbv1K7VRDydEPZ686n7G6zROP2UGQTb2IGqCwuFniXQU81+S0
6xcO2C+kKHaRCM35eHpp5qoyRPrtFqr6r/+qlj1VUOMqAHGOp8BqyEGfC9Dc2AB4aCRymhMcqD3F
M5hF/bN98ipSB3KBzzm8KAfpG1KoF9l0EZ4vfEwXFkd6vxxNb9pXhBb4YpqThs7yQ0TG9tFJ6kxz
EtFIYHdDD0vVYxAsG56U2r8T/M/6bKiSJNg6LegdMYhrHtwVmujSH9NJAeeJ8q9gaThCuM4qLnAF
SXT+cvVZPw3+pQPq5TVACTUDPSyw5dS3CpSBklLxuz1iiOJ+xng4dGDnYkazg6jDApnQ0GlcZ+G0
kRM//n/K3GDs3ZXrpF65HKjl6mRNTBnzaZkfhofC/bHGieUQvT+0X46R8cHkqdlS5hPSMP8DfiL/
Z9i8HyiIAUHF7mLMsrQHEHBTS/GP/EGVS9Ap77IU47Z5/ARm8n4JOwGbedOK9b6ZvRx2SJLWAxj6
E5jarGuiQLn/DcxL7PioEbEHXcnjrrkzB2912Q5wVD6oIM4Uc5NIyDSt64mUNcUwuif2bvumFVBC
11swYXTw1Vmm6ostcpxKlmSx38ekMrsBZnPANGzEfXm0KEJUMxMAR9rmHVXOipqORD7CDmecHNg4
mIoRHanSKiOvsbAxLQSx7nWsPIGfhyCEqGEbQ8T2sUMSFHTEhFDa8dItNgYSnBFWs6sXq8xNWpuI
hyRDi/x5Z3V9QBxTy74w/f9iBobevt5TBnXMFtrLD/CbhGiFN9el6e5toahJGTl3JaQQDqLPevx/
Uf72uK4nwIY6GBg+28BFAGT+jJ3toBTJVqQAC5q5QYAdlxntDrpbrlJTZs8QsUYtuT8etq0zUZVw
Z9O8X4tsFmIEKI87oHqZG3H1ZLvUKxkuJVg7P5WPV/i/xVRndvZ3t93ZU5xkBLeXI9WhBJkAGP21
DuBIdCiWkv+5WM1bPTc0avr7rpyTMEWac1dfvcFNQkmi6ROl1urWOraUYUExds1tze8PLQV707i+
fAbC4Hf/j1y1BrnsdwGi6biO2u4bJj9CbgmbsWnwJ1c3/qfXUIedgMzqcLzyFxKhIKZ+gWpR6UX7
yDa2vow4gO7jL9yoYfT94Yg2l5SZpNH/EslIS8Y6OUOnQcaWpR04WRCtAVxlPTU5kLWoa45nHvPc
eaDXdi8rPoC30IvDvBBfz68xw41/HdM8KZPY81ETOeG2ploUXBmeB+/BLs2IObT60NN/Aweaw1U4
3WuaO1xAg9dNyyEUxUkiL62j2fz4Vw7/xVolevIYkvsWi8Xa1hx+j1ImmWTGenMBYijarI0/CA/k
m124hbcSETpDQzj0rYG7ihES35JF0swlQ1WK0xEbE/WuiRWkcLVio4jRY4qnEYJ/L3XB9Ka4kHic
STdjD3dW+HOzbG4tASn3PqAJZPFHx5H+ngkNVOf1DEDHJkiiktvRzmz9d6pNaju8SGCx1bwGCuMC
W86/txYyzZqD+4EkyiGccxJwvnKrBfIP96uEF8Y3oKA13th0lxv0GdPfP5CsTSGDuPiEp/AyZx/U
Aey4agSaINDKm1VTd+WW90ks8ot7FH5T2h0c99AGh+vjf5i0lgUWBS5agAuRpWDULUTzcFPRTXYe
AcS0RylVmqGrgYavqKilBvkBHOlew5WRvcLePxdx+JKwXI1A6JS/z3qlmRWiXRuDiRQyyjFtoHE0
jcP6g4+5l8gSDTZNTUkQ2IMPk5MfHECP5oF/9UVuV0YrUoOZVg7pAYcxwHAbr3BqFaF1sX4Smxwk
Lqd0CNNhJoViWR5+GI1iIpucm0inQ8jYi/dEQB5uruwbRGB0NIqcTh7vhzsjAT065eaC9WSqWmCP
IB2hEHxYns/igbWAJfupj5ml+7KszLlqJB39XHrm2i19ETF+4vDR1Tns/DOhsws3cX/to3mbWKfg
nFzk8MJefOR1wZ5J1u77wrY4QOeTvYAbRX/KZjtkXkZiIJOE5Jb5nL8licq3YTkqJ892lm77Bee8
3rhvmnAOAcLSJCM+LPlD1eHetM+tYPaz5CWJo52ziJr1J4YdYgCVzkZ1oeRbdzl7XX54HINBmnJR
IKB++XKyETylRv8FtxlckHnS5K31wlLpsDi6KmLdACa2qQlFyplENMyC4MHdsOQa5BN31W+92b6N
Q+dGqcithJIc76qiEfG1WfhvXyLFCk51HhHlU+OfBwd3Jth02R3Wniy/o2WU3wfK3Qwa1Ua+Y9Jj
4UgcCQoqdREPVMvgqX71IKog4PXAaxtH7DJ0eNx3lotikl8/gyQPKAWpNSRAOUQbRqO0kuXY8BSK
2HysTBLqzXM+/GerXIOpCGb2Wk8RoDyqo7OzNTmmcJfLpxn73PFjiuX8R203ZtzTIRYIBKxr459l
wuztk11kg/ypvkDP2YY2+ExhduH+eS4vTemmbPkcfq7S/y1iK+Ycq9LwJzf9wYRcsKXdQkNfVxsq
XNo03i3G0G+GQwPKRmV5XPsrCESQBRCikh6Asf96+O/arq75C+/c4+sDV2KxL4LmF+noh9+H/EEQ
E1tMKpob7bwUC+mRlKIQ+PrLGNVZha32mdfcp73zyReSDr5qkIjvUQ4X7kuFVP3lXASaVvrh00pi
q+jgMp7VoX31wIVkGgsDHDcblXSg3DFhiMfDCOipn7Y85fADDVCau/HY+x8UwIPLDA5owmda4/Lk
Dwl2pDo2dwJjEu/+DO+v109xRSr/aPtop2UTF044l4WdkRGQvfnI3BYWW62tAqStoJ3k7EAgY0gs
+MySf5kpimcRgFm/hcOiElV0HHLL96MVBtrsJrXUxkGHj/5WcUDcF5q5mQiOY/emxXvebIzSucUz
7Qb4OQGCpid0L5MAIAWz601xoVJcLmErHYMX+cdlIwabYEKXilZ4paMLYMspov1Vqitosmc6Jg0l
fLZHQRz/gGvRUvNvlDXAp9Esm9LLTlZYdPEzhuw5vRdEGhci6zN+5sJpq7xMV+IHn/iPDWh9VI4y
McTOMU53loThYo4DTmbRcvZGkDcMJxNzMhLbLyXVV2DP/Xv4F2LlWBqKDc4XjT+4WJOsHrn1eHaP
h08JyZmoBlH7vp51+tZf+ihR9KEiPwA+/Ntty/MyoR7M3dTyTPOaR8n7MGhWzotV73mE2MJmnwuo
vqcpA6kJN3raCD1PSCjGPdLEqxKWUQ2efCNr6/scZ9CYOhNzgrrQPKrT6MflTb5cndkOG5J4Q73h
usFuZS7fqx9o3XLX4OJRndM2zLTp/bYZO+wJoZ9hSDzBi4ce8n0Dv9YRLfV85eH4FhlANEnici6r
leuaUtqm0inF9e7Ql9dG5vzD+ikXMnz8ZmOVtW5bG53f1zO70Yjk4jrfPOlX3uQJOsrZpB3Rl904
UFRlABtueda6bCojxy5Sav0CLHXT/26eHK6/lB+mi4ikyTtLVmFjJ1E3E5J9zfRFA1mz469Xl8XF
bkDPHgw2hTwynmlMrBQaMHsXYqIAhtlPqcd1dpC5rvJe3QRyXNS6u1zh8p3NQK3r/p2sJNwiBPqV
QpSKJNqfCJpL/yoIbcGJhUL9OGqhDr+VIaCNlDDkX//P0LaeMxLJQdYJq5G9N7DFHzeon0VShpWm
1vNX0EktAfqKqwzj7Cw4hEl9S6nRPyBRKhR1JmO5LtZ3kdOo6d0JpnBYx+hfFQKDgjE1/rpAMJgS
FsiSaNuLDTu4Gc9sjpF8yVNO42LiQ6k+0cOkPEy0TdWP/vufmr8hd9cJ4VxGV2sflRlFsZobl1xP
c0CBkKo/W3IIHbZdkWhwNSYSF0nL+yF5o+AGR9va5fTPOie5WESJ8rd6WmODFNM7wYjgHKYZzIqG
L7ypayfqTZkoheVjiz7zo2pKBxx6/mSCBRCnrR09r8Ipy1wieGwlk5nL6RJyD5LyfqxMoPRF82Q5
8L46babZG3MhGdVmyIl40Sb9tJVEbM2/cCFjW1w6RuIFhdimGPpwLk9zG+qCSK2166ldD3hPA2v4
/AXTJtL76FP+vkkP/L+dUY75UShSI1aBFaIstjCBX/9ekG3IKxzKJ+2CSM58pqLnDWdeZF3krcv+
NSyoMOQ958zntunUODT9zsOIQwilKDHWbEmVipVisbJEohzXUnk08f1a46aaCWXvt1M6VN0TB+Yn
cyNdlXmSJZaieDxu3+rUyWUBA9OHy2tPpIGu9NBl9CaHszrWVUSSWnPKsnSx3ai7y89GFB/OPfWv
xS3OGyjXsGFHgAkXbflpA7eMpCiRcVWL67v2neauTKapTvcth5hzA13RQ/RG1oKd1t90NjdeVesE
aEz3j7vrdGD8Yw0pt7tS69SifP5ydv6ZqLZen2nJeT6ZQZX5tyqqyspj1oIZr5niv1BB0cHxaVHQ
+pGv16+u+2aQ9AsnCxW38+3DIHy1bARIULM8OaGyNhchhKMyeAA9OImq2lFysVUy01G5ejmGO5M9
jS8jzR48r84CK0wPMh05UHWI/bgDDI89+y5NNkx38T/ZDM7aFuSQwUFMtLSft6zLWNEBLrt+hi39
bo2cAnbkXSPsIKrHMAz3H10mr+OnVLoEhJhvU78vuUa+k7ps0N8xbKjvHbaaDfLPC2uBRcKED9pf
tqNFNrhFzya0dH2yAmQ7wLklokSBh+C8maBt+6k6yEwYHggQ5x2k9D6R9zul8cI9W2nDdNeT0r9n
HhB68tihS8H+FQvYjDF3/Q/POyCS55+SUdidfv8Uj55JRtXNHIhwaT67WHK+RIGPdjNe6uV3K+Wx
emxBKX8itf8fgGJu09/6ZuXUz8z4eDOGLfCFMFm+FAfI/fKwpVfQKj9D/aAmWa+YGMMq5m1DmbCR
txhlo47hfBv74fmYawNaSsXiDd7Qt1OIcLWHohhg9X9llN47OvWV3yZcOUAU8oFFF8OmKvd3AL6i
JxY3cIlbRD1LFweyAyCSpFSoDZRYkbZw2qqVBSDy4go+4OKOvTcDDyCZoVkdiA2GJcAM21iCDeS2
IRhLYaM9ILEy7LSI1gN/nzgRdcGLXYW3olwwUfQ4wqcxhT1/fC+XJJKNYaUHL5qAnsca6S+BYvaf
abJBDctvWG21SMiw/r/FU9ctSUESYFC8k+tg9PcYKqkKxqiqKGrIY+BMJxlGb1tVJvwZ2jqIPE7r
s9zeyFJEgyNTPf7xki4pV8fuzR7mWrXnJWs9aTWQMfkBtqxI/ZMgfu7HVfF6kzmSkJQYmnXBTYxY
Emg9oh5l66fba0FHjlvvD3jpQcLEwC/j036XD8K3ZsSl35zkbHRExPmauIZItbO92n0NMQGVII56
2j1CWA3LVj7KWsSyk4e6NLk3aPyJvqe9fkim7vUl23T2lepQUWOSPm7Xeg5t2UGfvJDtfMbQ37S8
x2jEk47Wv7QewZ9L6M0RTRpzAV6SpUSVH2A+5Mu206z5dt84BhubxkNr1/uhETcgK3xOOmdcIyT4
nm1rWVXGSeo3+zy9/YMKtcM1tomIW9f730NB/tyvTu45VqZ/N93xL2hX/GK4RnBVZ605RC/16aIk
R9VvfzL10c837SWgl5DqCX0q+H9qgbZyCklNhiLkYJlodqbuyCpNcRvSDfXUGIvsY+ohT5GZqTfc
20nU/hOJIe+AfWHFVMLDXZCPm4YO4PKQZrzKtaR4OjWdN5eyK7BB/SgxL1Zmi1vK3mKblQyvkzUH
LBgeRquMa9ZrOAOpZEl3B9Bk5VuoQPUwDPgLwOavI2xpPgDQnQw7FjjgCntU9SWcGrHK/q58yfwD
iQ5MSmjpCnhgE3ne6wmOsRjTqT1aSQ71nDw2rFxwGh3AFe4Fcy7bzMza9QcJSxM3IIJDfckeJ6Gd
Wf+GTlBqxCHzvaALNSvwX/Mb4MJfwu403kEc213lOfC4dbXq8C4FcHWKDhba5emimpwW2FbZZrC6
Tr1nexcbmSLiTv/GBz9U/SXMJVSpikGIMcAxDzf44pWyWQCnzBqim0AyHd0D854OP2d5yOtQnqtm
JaqtylqKIq+IBahxcLDdQGcT5pkn5FrXgIWgIBqr3Mwl0rC0QKnsPMGKsOF5102zrisu22P17YXC
QOEAr7Xj7P3bepdWXW8ordA6+9PpIpnZqocLl/p20oykdl6PomRb0nk/k8sIXLfilXUvxvmwDDti
429AArgqvvIh+QqiDxw0LVtDmnlB63PReGdGzH6mDIZ3/3L1EwgsTTZYyrurNuowkn+VY1Hj25+v
6FQya4rDXxP83W2kd7cPJNZwg4zHRBFNuQwRlxxhb1GRQ/GS2sGoEA/s8C0ZgTO92ETSCXfXwFRv
uNeuqUcY+4tASDlm03xki7l2K4GeNx5TavH4DN8sWNMSEacMl5bGQC7qIj7PdYCF4j5e1BWIH3RO
7uL0hLe684Kj5HKjDSxD7vEaUGhSOGXLPIJBGjDlQVCX6Bq5UJsxyqoIWXt9wnyZ0Y4Cc4edJDFq
o7Vj5ZHC/OMpNNRZQa1tBZnwVIVizR/AVD1SDncE0mzcUbEoRQdhPiuOQn3btNeqVmF7NVCCW3ul
eom5ykcFSSP/fdZjLRB0mCcGsW6kpJNqjIPtDyMQXMu/V13dvpAs3WOFHBaazkmHwKCoxxWsgqIV
jBIcncZ6EINGH3F34qggcEOHQiLAc1Hvj0jXAZ3AQcBWoK3OqiaVQ7qOdnP4P4pN3HVzoOHM8iFT
QVZ7uYrkoDnC9JMq+w0q5rmlkrT5z1lqzHOUkrIDOt3X5k5pR8JvoXMcjPnrV3g8iXCGB1C5wpC4
iR05yfDP/GuFGNqYBhbIJfwUtt1fX94UrMLdoTT42x5TCt93TEhxhTtlm40fKwhqlG2west4wmP3
Wkwj2tLbQVknDq+i6bT8Oh1RCCQ3EaszcDiKEkSmORFDorITfsLKJ9m8aokBxRKsi31G5540EtfZ
6wxFI3gNLQC6tQQYP2pYgfDK7yx9jop3y9EqljFTWlX2ArXcPYYlXGw2hB+nOxROaiSNpbpjfKB4
a+Iy6O2bJlNbnwl2XahpFlyCs92dZshvMBPKLT2ukfGopVGJgtTTIFNIwC2EDS08Uvxjt1/NTj/Y
8eeFAkacZjcxPPOOykQetR4VdY3sY0gYKh8pjMqwIW49+ULSwC9RCvcW4ljgbCuTV6KQvpF8hUP9
PStdm6eZww5029UpXHdyfeRI/HQUIpv060oj2FaJLDLc8fr9QhOFByhFnVGvSlIinZAfEoi0rxv5
Uc9l41q6VQv2mavQYmzVuUGwPyZ6IALREBjD9Q8V6SvE5Zc2rW8uW48JASdo6d3JMaQGwu5quHNw
g2/dyfrh/KWKocj183MzYQdRD0ERTGm1mz7QXzfZ9R4GFxLMerggb8c93vQ8dtPjGgXVNgqAr8AW
djqaz8dMLCOq6kHbQT1AcoK36xBSftTG2y+UV7i6DZR4mwZtQY4fQ9cBiH2oUAokhp4/qdajokNE
ipzNSIoBoc52JCc4BNIsgQ95UyJcbNVXi6u5YWgJAVtCmh9uhRMAebAscjZgtdx+Bx5coRv6kOGH
3aaiU30Yu1aPc+pHc5IGMhiilku9hhQZutn4wjceiTsAA+YiiLczZSj/g6j2JlQtZ8v57I8a2GGu
DOd2YRRrxnH2ppUZbc9J4mLuXGlSEe+BUs08gUGfczCP5wYhWjFTR3AWEscKHmWnA5i4Fpz+ftdR
XaLN9b28rjUaMspjnCoU+Bf+nIvHHitjCXvVPO90HPFSpSQHbNjQDClm7Y/WBkHGd0wWidfNdzBc
OMNCTGHQCnYR+PpHtsJoD+oN562RiOp2ExIPUp7dQxK1X0bGxypl0jUJoAuUhPB0vHfJpZfqn3rv
xGatmwhyd0wAy/8p0Pa0iFmjC+gIqzrkK8XXsKBblkQ+usS+TO1+g69+vwVuXHmHGn/v7IGGf3o6
A6+wUEC2u9OXdlTGeokOi9RPsR14PGEo87oGV9sSxkM+6Nuq0YsFtLvU6VQNjELkaF3ltpp0jPAB
SNXPRCFGL2IWQGCUxHogCCrcPT7MrihffGTCQ2zqyuf7Nozqt5sCQALGkQaQabsOZ4Vnfw+29dWy
hVTUuQV9TTTXU9vUVpHtqLy99C/d++Ama+7Xkd+/LeXuFoz9SvsxwTzj+rMNOmqGn5ZKBLQ3hd+3
j3bzhj/ay3kbKXGPMGx3uR3rUIdIfD0JgzHPOw27LJdrZM5zZ2hX06IJgmUPZNxkpDMX2AQ7pm5M
3SkS5DJz/nKXQD6oe0URYPf41m6GWRyYewyrEztnqCD/LxlqOxDJcUe8eEGQYUqzTPwyWwRIxRmT
rpYSzjYePGD44zO4XOK/zEaYeV17N2xzcSAIOWU8+aqZlLeKJT96mTMUHjfPyJDwvxWxmllhXLNz
ksk1yHpEd82UmZYc0W2OtdYrkNDadBeb3EIVDzqQGVNRDzToQMmDD+Rl7n1VFUACpy9cIfDKL+wZ
Ec0D45KR3YlyMY9S8rLwYxKp36YCANaTEEhynJmcCsVa/WfsNDFxH0iIilX48BTp9nuFBMBLq1qq
VlHPjBoLFQHUIEFhVIY+VTwr8xjzx0dhR36I/NfjPta4S/WIM7vSFF57XcYwm8BDEGNcYjzHPRzp
O+q4KNLBix+xyNKcm5Qlmw8F0Z93s1vmc910csSJdeHSzm6fOAQdQmecgaRq3uU7tazssfn1h0F6
rAQIhhDy+9wBXwjc9F4ZEob4/+KJDMBo813I+o9miRGTzW2QH2/o8R/pR4PpDnJKABKRhWEt2BoP
eklCjXan2M/02A9nM34x5bOmHaroDhsKbbOSFQfhm0kLOEelD+47JDs9m4+gAyA1Jo3kxQ1fiRHA
JxT8X6wjdZ2gmMtiOvrHomQg30uiA99Bxux8b6CjBPug3+VI3WhbOEbdjfoLXRdszd9rboAT9wBz
Cs8uH0qOrHXIaSSDZg2p9cV2bhd/Q34yOjcu7C4Xf91mAWbhvazHcUPaCZk4FUUApnQEkD0bdBO/
RevJbQs24SYISjHmWVAfad/rr3ZWnWqNPCUUGwpKm5bAuKWayKOi2J0A6WR5jkktjtJIrwObUERv
zquQAEfPinh6VdZn/gVnbPeF5JdUZNe+pWVgvNdKUj7P5SH1j+2/bY1db/hF2BbDrmwIhJH54mq/
DsET59rYl/LIw1YxSNkbqS/+6TY0vXcQWTowd8VrLzFnbZGB/JZh/hfqn0tS3ZKYpRzirr/GX9Qb
BD3mddiTgoYk4m7DyZJttzHuzkoYJIKgEdGVX6DaxrKEoPR28Md6BPcOv0EK/0Ajs1qJMP5BWv/7
Q9Pfn3jNoFVRkxriljnKqyadSer+STGiuXyO2E5GxuePbisM/hE2bjnaUoUkZXIaWiCaqh3vNspi
dXnsbStdNmYXxrVtYMmUljSmo/RAyGfEl60VCQZlvhtBWJjioALpZ/zblQOzMNLdYQKPcNWSZQE5
Cp/Z2np11usqGMLYodWcroUw0uW5HlOdfmq0+nr0uneR2gQtzklfKbVHujZ9mvh5O/yYoydtigzi
Em85Pnau2kNtvnqOVdjZdPUUn/Rk6gCjvjMFGWDYxRViOdn/IuAnUqeGxE7iNBHIVTZqJVdUNj7d
EqE3xegyINLO9AcG014B9bD5L3/YTvQ/6X2sU1PdF6WUD0CLs5B3SMb0NGj2PhNxx/elxtUQCioP
EsxtnMNruNVz5GoeLC92/fk0hKJIOMyqCSYm7R7n+LjYN8MCa7cBiAzh5YjnGypm6QKE8SxyCWb/
Vh75RSmdCaqfDVW90XOgeSt17H8lupzKXzzemjt5l1yhKCi7Ig1O6bnKEaOJ+34ogWao65vmQD3+
Y6mJDg/GNfPtIi1YxMgbgMOCdXAbi4MkL3IdDkcu5LBm+XVhH0r7iDDwaXSGfPuMO5SBjiX67fHF
AxksUuRZtiFs5EmcFbYU6PisOlFQW6KdhtpOfXxzmlQCuHuxSMIQmUgpZ6wysdvia3eDdWs55Gnm
C3Mx/7QEhNvrCn11zPk+QjWb+EY+HQf5RUdGeAXzJdZUlIu2O8rYoGcFGYL9M17M68J4X0sGomG0
dje0DMUT2uuhgL2QA2w3qvxCAbES8+uHm4rRyBMnvR4Go1Ta/hnswIXhRfNzL3iDX5myEKL+obHp
R4DUFxQdFd6p8aa+uNpwq1P7k7JdY9Y9ssy5y80T0X1i4ByD10g1aaQAv2fT+IUfv/ziDlC+VN2A
+eVky5CiKXjFANUJmTCLhdlaZuI3MPE69XlZ2v5BWAQvzlr5TnEVXi/K2KQlpHylO3L0s+xTmW6h
RmVhUrNcKiT67Av0H+Y1C1x0ElgmF6jighu+5nF1EG2CUxhlPQF3QB/YLflc/fsHU1NUfheuvOCl
Bmx1XOfoLiZaFo+iKQ9AULyEgP0rEEGzKcyO8wCJnQuKfz8qDtpwYx+cXelE8FioGDgbp2GF3BCl
50tRCWMmEXEf8ShEVPJza79dYZbGaBs6Z40CxzRRgt4kF5JZgmdoLJA7cSZHSUapRAYh7Ww6BzGc
UT7m6L4ijVDaHPsJX75eEjlzxIOY9T6PBrsoIzZNmq6jDK/IcosSstXCpBD9I9q5qdAOq7VKGfhw
1Rulck+oHbsfeczOFxF2CdZ8504nR1UEWRU2Us6dn/hw//X8NEwO4zpaBxKC2oCzszdZWy8CVyA7
G/ndos4GY/TISKvW2oJIuViWCj4rAbBpXjvpQMNRMs53J3HxtaerTUv7wz2nIrqVgW2DufzFQG85
uQZ2PN7OGTv35lLMg+85a7MihROKs0O+C+o+ZGOFrwIlyRXPUck0ZGlimLvwZxppOKbqRUMMyEK4
MKAAUTqcp30ggnrVgtOqXwfVaWiklM6D233PjtMfWE/9oLeq/Lmp+zGufUOHgOXu1Gy3U1iEQypK
sq6yTkwRLW/7rAQ9CvaSKJDaW6fSAjz9KqKEng3h7huOy5daktFBGVNfGgdrCgus4+6dIR4MtcD6
ZU6oSeAmlWxPlVprn53GxynJpDCDc4JTT89udbuDf0FMknsisyZglYN6bui7eKCMna/owy4DWh+/
/xkCcAzQhY16keTCRK0VnXVVsZUvVWJGHRIYEfAKcJqqZMQR3SWqCvTlYdtkN3aA61kFma5eJNI3
Jwiv0KyMo+1xsqj7tC4PTXZkVzXWSnsEBzk49kWLRIOXuiTMnEgbWhO9rhrHnsgxByR196Pa0Cf6
CQIyuoIbPPSCCZf6bZU6bE/gaWPHQssKWlqhIHbX/WQlAp1lhiKqWLLW8bKLOxWLeH0GMjhmUbLJ
y5/kmRgi3HO/n+KXmo2ut6OGyTHHKkTjtGfIYMiZnVYlaU/BKMEo28kfQl6zcoahqedTSXTFFnx8
hVCJ7Emfm82Dn3zdwlgnBc7rYab2y+pLQV5p6Lc3aXC4NSsuxCQbbQfFxgjj3OCNmhmkNHRGVtAZ
//ookMmfQbr+fzgQmZ8rLDpp7OzYo3zjtHJPVVuT06X8yrsAqBANEWIQy4gaIIECUQo+tzFp14EH
mVgVw2vv5LHfRVbxVJXY19C7CB82oGa/cmtjXA26cppuwkKHWjwlivjT7yMOxtdCyC1W5IQ7fT79
9WZzfnnYna/+oTWrNzJeM41D+dS9FnBqKunf9iCSSruqIoVZ1C49z/VhehX0s8Au0mFlasJx0+fy
AB/0PEAU0bFO1eXfQOUNJH5zo3FSuEadzlM/IB4eplCTZijc4CdzCrIXGSQQgJ/SZ9xaC2Angqs+
3X8W1KwKAM1/ukE9KC447lAbZe3IGQ6VtzUSAaZebRYBS0ZZIczRR0o1z1faCp6uZaTn9t3+9cqF
wYdV9/CiP+DVKOMYRc5o3Y7l9iFXGfJXZiOv/HuAa+t8EhgKyx2FdwF424OFT75AmvhX7r5PJcSo
hq6VE75c2cSN5SI5UcNY0e5uBXU3UBfRjA599wDDJYENSoxkUcn1IoapM0wGzwULduQ4jMyjSx+X
LOL89kjbLJutqOSR8Syia2RonDAYYv+Ohm7yB+kmro9FphY2E0xoakVLNRjgCXIkznyoaBslbfad
hVryop8Gn5evk/f1yySX2trYPSxQg/j2BGySDHQdhcGedXjqxSZ8rSMX1/EHhSy7j6F+6K2GjU3q
LXEVm1JieXBApx5w+Qr3KhgTgQ20dc00GFDFiceWbvlET9MV3lsDocD3y1g8B9i4oxfhFDD2hWaJ
JyBE8RsQXD8wAKYfSu33xBi302Bt5eLl+x1/oiy0qDjiwdvoyP/FXmVFDV/pjNDhmjwXVgLYKF6t
aH52dvR1ncbpR9u5E7+a2TQb1TbR9T8Vm9mMQaobpKAbnWLPJFCE200c0C2thrVCITq/zyflpkHu
2RFqdwLFRhMl5DeRZgCdi2m3iNjbS439jMAkVJe3OleyP9f88E/QVaPYUZqVnwFr9EbXCtYd1YCv
+bwk6OgyeYuODADfnv9lSo/Wg4tRWd94UACCcCErRnMbat4mIXdK2qyxL//ai3mX25OpJNPAAASV
YUSALE2iMnxwzOvf2HItvp/VQ2lG0JtNtpBlYb6G33RgmX/1j+a1yS/yh50OuMkucvYrEDQzEBLX
RxXuW1GP1XSTL7YhsUEJPM1WGsrDV7p8IDcGIW3xaAoq7IFBBRi3ZhXfeujJ6IqDVP70++zyhBU1
QvOtzKwBYTWCL77f6h1EZcJFG7kzWvVr3rY6CImNbzZums25y3vDkd2x7V+aKrGoqhuY+/fz2OBY
nYlgP3jLIw8tBPlhCDv40OnPAkQpMTVRa21vgJm3DhEvXZMNrNNus3IpOTre0FI9E9enhNcDMwyD
G5Uvli+TWvvlKAU1gIysXq+mUS4TjoDyjfCK5ANF8aQY7ZgyXaU5xqgYmi/rqKWPjxwjBbOXDvqG
x4DaF/uYowBFrINHLG6uzgZXfMEpHKu/H2RILqfBS2T2Du8ccLUooVHuYMBoJKEPwZATkop+hItC
eFMCVEaDAdcZYZ7pThCC2MXa9Wt/dW+APWWH8DN04WK3AEVLZ15pvOqV3bOgbkCQscoqQn6WA1Wi
b3lYUmKbozxSK7X7rA79teTWvlR1DRYVGcXSdVAJVnamsaO1noeHoFdV+cbtCtzs8tfa0opFGfAb
VjeYUicC/172ECBaEqAHEGsmI+7BUTeyKdmoJ5HiKY4b1Jp19msvpecM2Pai+vX7lygcPS8ed4WB
q4D205rDCqkSotRv/pPagol6xGjnCDMlNCRo1u0gjQlM+2nTWjeBXlVhfL1H/0spIbnflI9zrQGR
uUQLvJ/AGQK153x6G7yTdOnqLkyX4h0qX5dngDtNeK15rwdcPbnIDl9aW7kTPRbfWdNtEvHXgVGo
AlVpNAGk+7MNHfLnSKQ4e9lWwDW6VqFtpzyiu5kU7SO2YPeCADEIZPnK/YUDA7MmF91Kr/VepALd
tg/uImJA+dxiyeLipVa0hWogFZ/HNaH/ZQ4REHn65zb4j72iBV3bgDs6tld0L9IksGGU7JXYZlxV
Yabwz/STXRLBn9AMYiw+IlRXOjMBjQFvYTheXOAhkvkMiNrQ+pTuK8fZpBaVGWm5PvduCgUcVDZN
9/ujWO+oltiXDv67a78/LlpWZY4aGwZt5/38s9OXOW+ymUO3O1Obpj6zvlsLTy9YtGk/BqKoQrpU
kAzY3aVIk2hSpjlPbll22uygtGGZ+jlJXwb5T3752WWDfDpiJ2+Id935j4LzNM27vE1ynjqchZ7r
pJwMAX1JHARrsauaLmMXKAC0NxevRiY5ZW1PHd8IkTXBDW1GnwiF/8JnZlM2X50Ne3sGsEbODdQl
NV90O7a+aTakUI9JRk1HeJ9t1iMK0zurIZQG8J0VGjZeMEhNVj0UR1Dz8saeGSqQiZdDIUFbugOn
SNOzOhr8YHa0urY4d/C8WaRolYqQz8yyGSRvor6Mv/N3VDeOVDyQ1NTqnU+B1eldSdmpspCo9s15
f+sxolnY7palgL/KRbBhgM7PScWVwz/Gfoq8q2isZO+7aCDSFJGwfURbj/5bH5XXHtLeva2PD/wU
xQV1fsPC++WSJCtgAOinckfOpBbvbJjCal5nIFIJoPb2sJGLaE01qcjcMTznvU7vGqrrL1jCqpbf
s91VT57wlb6oDiWIEJDCSTTzoaBnwcAodNiVXDOgCk7gQDPbvd7+Z4nYHBaJUNjjnsU0/lNmD6mc
fb2QvI8bx01VxQGvM8/aP1T3nmgoe8CZ0qKB3Vq/B1qFJhqTrmWLycncwwdOjamhfP+7i2EuuxNG
nG34C8DhUglr4E1D9wezvN7uyjcvgiY6a+fk1EYARnna007Vq2HO4XdR+LDn9j9kSRo/LgjCyOa1
sqgYmF4PrCP/6jLh2AokMKsCMxqphn17hvvFhjA1xDKHbvhXs/D5LzTNAXtTvLVujcVOU8ciL2ZL
SHXiZdjwiFp//NMYoZNyyo9BmB+jHzeDwGuYAcVdu/M8rF3KY+pD0+Y6dr+sQINrHSuOOCnIRusK
iV+VSDhY0mi+gH9e/bhuOHeLqmG2YEtFVnVdKlKvyhvssqbQHXgBFb0u6Hdes9ctZApYazQgh/UO
8DEygGKiZllQXB5STK7Ea/se/IJsY35HbCH2ctmNplCjrgYw5Q21yGobZtVNBeQe9biO5vMElX7H
kH+1to60OE1ZAsUCOs6+jdJZ9ufSzccvxB6Xr4jjtkld1ZJLc6S5JSOEItw/+3H3aTL/X+gwradg
e7Qbat/CKUtbqTEnF5fASxxa4ajO0AoRjpzS3nD1O2vUQwskjqoT6aD6R0mUIqfcaEcVvyAlElOC
cL3FMYyhgMU6be1FY2OX6VQTf23WpqETOTK+BXjfHzedQ4VHe4aBURxtNcUNpeudCQhm9ubEX87b
eQwC8zpl9ab/xrFIY2CSR0C+7j//uVYWGXUnrIP/ErSEIuNkOg5HM91V3nFUogPZO2laMDdWG9ue
g06whTY7qnAMeAZwH4kUD64nwmvlBjbqdqH0nPuDl77v+Ya0H4ShD2C3+K/kf1PfLZItiLspv7K4
8UPpw7XOaS1eGI+9WISiVqjS9CzDpTl9QE+CSRphv8I5if4C+JwlP05XvtlxzIiPu44XqYACB8IL
YN7yQGf+r99K8Djwi5GT2+65DLwCHWoJgIXun/JN5HDQkGs8nJ1XI81BZ/PprB7qFdeGvazUI73Z
Fc4+x4OirC1zWuuRUHLXjIvGCTrd192ZRGzrNixzJPt/+pS+A6yBsAm0QaTzTiRCSSuxIx3h1rQV
Fi0Uf795234ro2F3qUvy1WFPRkPNTngxUuQUyj4djuxsF9uD0HzXf/2PyUckWEBkMuhgwiqk5ffa
Vo5Rvu2acudF3MH0Fp3w+/EPR3wan+Xc4ZjSf/Hw1eGf3bd5s9ao0juPcm9MonWtNEpODNKEQuRi
Pu/h/W1AaZrnPEGiCvA+fmVASg5mLBIL0lR8TfvojJm5ZXhOXEs35JlC/jw/33qckSOap9TGoAV/
MdOPMgFBP7MSDU19HB2bKbvjUQsOgCu2LcUIqd0Cat3uair7nmPdezGQY5vQyzG4UU6XKUyLqMz7
IQepBvJGUXisLHAfKzxL+8PQpVc5UMRMCp+0bHFAP2xalxDnDF1JpGeHjK3sJJpcc2zY97A8XpuO
VZweYzUDUvf6O0L8IAWG4xSYY6JKU11LbnkC5PjarjerCokJ4fSgyWuFsUJ343vA5sSAgmbsjqln
h3LFyT/cxOLr5YaEtbDoEj9/+rGHf27RsydVrl/S1IE81xlqats42wqsl33KDkVMPfpKyRcjv8Bt
knEiT53w4Ro/UzO2cbjKxXGBNjDKTW9v9yzvYMqVBBzQ9FMqY96t8vO77mnJDtmcU0XnBBe6wBhE
BftKdoPps9m1NB5+UBkfoDLWlQ7vFmHedTcVfFLE8Zk/k4ipUkvH2G5OegvY2qoyQnMRIzlVb65o
iblQvLrwDllX8vBllb5rdxEbreXhR/sTwAHHBonrxoYOOqYeL+UGKGCsuNWBciODybAxagZ/heH1
Q/qboZScS3FmnXTOeshg/D5zlyQuhwMDcZDQQc7bMw7YLNsqCegyWfLDpQ37R0FvQb8mCXG8cH4R
u6i4GRJOd33ax/AHK87ziU6x+/6Sa5AGIie6CLjkdoA5kf09AHgEWUTd5J7L7dETwcr8Yj4jy5ye
Fh9IqhuKCimkFNMPIImjTGvmMPu4vCGu+zc54HP8y8XzNygoQLBwCzteo/Fkch0sHRAaO4GehGkM
u3sXqSdz0DTGJM+iYo8SPv5UWtk9t3RFJw49xn+tEJv0ujhbs11MxtLUTFgVY17osUO183rKIVCb
9KsE4LvPpRQjemGZHmlNvH4JVyrrFv26L3iIFNAB+0aWNPfoG2x8CBrWgjzH9VEYwV78vdRxEfUJ
DTHjlt59/FUFknKQjQRKdVvWvH+UvLRVA7YAFmnHFVzCBv1Ifz03LfgphYcywDudw7GYIn0k5dIf
13f6GkkEPMRcyfYY7RpHd4VNqT3kEd1qf7h2pClSR8BORujBqBawVus6fQyqV9CdW9L/r+ZwgQA0
3/eMnIGU7bZIqST62smU+Yr/TiID0QF08ltN+EG/kBYI7lDyWJ69T5eYclqinkSD5Y/Wk6kkwNkE
3GUqokELY1OxqsNlJQmFfou0CXwML3OHlKDfBFGqs3EMK1tKNiaCb4AXuApKu3v/X+aH/GkjGo1T
+BUM17z6esxkwODTwWTkKk4PZI9shpnZVcLmV+tCqLukOKIRr1FlwjRM8sKmMIPV+whTdOEPASPs
5TwLOWTIyRuwQkXoLxAnE4Ez0ISRuMYkyudx/o4AdnFyqaETv5oOqLUaTr9Zi4RN8xDwE7grHrnN
zD/X9u8p5opr2spjRAqdwkHYixy4gJt+O/h17q3SrUyqGUln3itSWl6Z/LndhjIpcoQJ2rNUgfrh
J/ayrAeuFLZvAWWOCt2VfY6Zv2KLvTB65zTFSzX2cqPgxPWoRpSHrU17bnZdbRghOWNDPHTFTwQH
hCLCOKzZUvJtdP243WfeXzs5IfIvy8zyexx9DT0q9COaEp+fD0/7cRFvadWPlL/qetfz88z9+BXz
ZLClv0CSDc0EXxYIVnVVQBc55tfmW5CSJck3MHrvV+Uym/PYVK2gd/puM+HsT/dutWHxEl2DmYi3
DJQ6kuUieqXRw84Wozc/8Yyrq1eLOLLh+ocbS3ZuOBfkZDctOLvVm43EvP5ay5+52QiyF0y+dRBy
P//vfbw2eHy7TqnIFtCliPJXyl0k5vW5caXQiI2+IhqDjrzmykFVcfaT08NUU9gvXePZ7+ZzRv1C
1bUW9CUOQU6S5y9Rtrxim8+ERRNrnVafRsn6N6GnYkD2UQZpYBLySpzqMDHqeC9B5CWUV9KvTiYq
7pRKiT2Qt9LdPwysSSo2Xa/hPiIkQN3OC2ZRp4LqHSQl44qLDVOoWM9Z0fgKWP1s7RxnPzAGoWdz
6MpukZERjYAbwGKBqCM02mB5lQYrRrIdqQXVcSNI3yYN9KqTrKStUYtYLlifA2D4PhREsZ7AtZ1r
DYIkDIYuCYRuHWohU6R8erdszArILdy3QqvuKO4OxWiPTJqJPUFvvT5EmJxNRFxic3ww16Za37gF
sxNzUy1zkIDFstgZ7C+VBtoNHo/5OTMPMwIBKsE1VMLljnm3nj4xYrK2Y71UVI4ZRIyqe7ibYaxs
CNJBwWrbqpc4g3IrhYT0gnLN8ScMvvzXbZ9OHLCY1V7No4d7dp5BA1oFL2C/zetyO+ICLmaRI51l
ejlFte+itTIHWdBt2+INjm0HXplB1DBRa8nPrKXwVps/a3AL0AfdU+NRmo+zOv0XN4Lz5z3UzJon
zLdVhOWSdLWc/FKtZblOlnkHKO8ftrc0mra7p94nLs7tSViQBY7jWz5rwZbOcjETUOsfSqH2OmN+
+ehJX/TKOMEBp3ZNbiPuOnqY9cm3/bvhy1in33LrXZRRtAiJ5Y1M5p+Rjiexj1xHRut0cXzV4hoR
qo2L7pmvzw10SOWfnZ5MV4JovwgBwS7m4zP2R0S+YAlCbwCNWHTwedB9JqW3ShHHzv3C7SFry4K4
e1p0I7emOEn1Be4NDT2JcOt8Umstkr84Lr9aFOpU94B5m+wLohvb/iqbqPYpzO+L721SDWLGFd1y
c662fiwc6G11zLqn3Sm974QjAHSRANnIGITYBMjz54sXyVnBQQQowE3pPpJpGV6D2+9LBPI95pKG
7pXm76QVsLeUSLNQ+fgbURMwJKaxpmjOh5+3spbDMgoW6cDZePdY6roGynllaGuP9Wy1ANNN5H35
xV9Kgvq/uLMltS+b6K3pKl0PJTlC9h3Fsf6mWkkeI9E5CdCmfBQkoOhpNKL5OsYE/NPjOzJic5RS
jf+YHOo4jWuvCBxY+Mkg8d8Vqv/D63RVBxCvc3ptXYwGfyfwDtBmbCaZDxofW8X8C2828hgHz0cY
DNJM8BSrgp5+Sho5+v0pNcFg4I0sINJq4QNExWpxieOEhteznFOYLjMIW1g5wzI1N7L3YURX+DwM
gWvVoT+o8j/9Xg8X+FArHJm+sK3FeBNAgBSOFyFVIiO3bIact8XV0TxfeLJ5qTZfOxLZnETP527g
fin2NN1VGtNgOYTvqrjtW+1HYkg8R6faox/8H8hP0hAdwxxWxO0lYlOsZbk2d+VNtl02jbS6KyBM
wKNI6F64DPeJu6HRd5UVQHRzJytWXmdm0KI+CAX6OrIYJBhSY+9I9f0XM54p59Ncjnuj8ZfcZhCk
kvVOyW/o0WXL7gn/0yiIM388UUB2YPPoUkbwVrc21Osp/EYdy8OzCEnFV3CEFUTInuk273uljIY3
h+GvtGZofC3n9srvx12TYXahDguurB0XOU8ZjjFSHG5NIp3b6JSfN1SXd0k1i9AqRVTzT9uuARaK
CmVHp+AsuXN/XnB+kkKQRwZUzBaCz9fm0BSQ5khmy1TYpvl0FU9rJ8hYgCIsrxaVUv6rBg3u/ubH
nn8tZfX4ygWAhJJSI+mosHGOlU0f5Ea7a3+rlYRAf4D+MH4na4p9RckUFDDFCWTHJYDCSx3WVfNg
nSGbP+9/xVL29aFHMmCFcTj8X84wxGrMcFIP8afailVTEWpu8QiTrgwaPGpZXE/yaNjPzGswd3rq
WNxQZAl5CxqioNYseCJR3o/XAaBgKs29SetaIKOQuvzLwHylyWzKcdU+YnuIaurMCDTts1OsE+y+
Ox2Gp8y5oRSTc8mi68FADt9H5NHDwcR8IJg7+3uAD12sz1lSqVH0uXsgI/K6qnTEUwxu2eM3k2V+
jIANVGPbF7uhqrmLExl+JazrMYm7+PgysHIkDslUSESYmLOec8MGGFWdrT1d90vcZ3/KgSrPs5CA
CA71TGZ/jHakf4qFY6p/4zF56QP13ujDIG5j42Yvr0KZjLrJErTh7CNt/hLDQJU8YndzzqVBLEFn
XHGRkCgR899nGykAIN4XlKO5YuuDrEC8C/K946bTxRQDQChUi9BvJ5/MwfbsKw4NnIrQWTKTAay0
hu/zjLCLg/DIBMijdJWJk/OndvEXH1qrq+6OsRSU1xNEnwa4oMhEBklWIAZ2osrhc0xseN/LMaQM
rwuyKgQKxn9/1gEeF/2Q6QLbLH/V2ZK2fjCwUID0cFOnK/dASSpZPKd/3fYZWcXx2GQhm1wqFWdN
t/4gNV1FjMw+h9uqB2fKAjl45QU+jZJTiVSBftHjqyY/lu/Xri2pD/oiOSi9NeQKlgmEg5LCf038
5lljBqHEOOFuwTTVwP0iEgeW4dCEfQsScK9KRkmPUUnPPHmZxNrvLs0UEi10nSt05rxdj5opEAoa
oMF+tjmF87e8H725XXDRyUt7Wk0tTyQG4MH+pag/uiZUkdwOc9LjU7dRPjfYnLmOFmSzVSGjeoi9
L1PtSM9sWGnOJS60aEkYb7R/884c3ZopTcVvxt1TrtFYtvPk+x9dGLitjRg25YkIJeK0tMF6t+xc
hWmDZ6MIXSv/t2Lg+bekzxIMthBMge1siEh0avauthkOvVhAGn+4OKzpEmCDGHBkLb8gDQaVj1kC
nfzAz8GhNGopB/J3xQOjIn3DaAUDImtN3mhfwd8EFACrnVzTWe/dpFAbkBy6uT+aEy8Tf6s6jF3c
W0tKrFrJ5l2/mZLSIiqvnjqqTZcNxbmK2+Amsq0ba/bo2206kfoiUDIU/9UgsxYGofcPKyJNPRtk
KpG8B9gdxQo6hyISp3DNJK7xZNfTP6CoK63KSsWARbrCuDYq6QEqdI+R0rJpKOGVqAPvhU3sOmor
eTtpID+MXKMu+otJxVt8y8RIQ7qpAEjVRyyyLDO5E52+obaClj9Y15qdezxFxEqaaCHpCZt58lxz
OVBdYyqOVZbW0dHHjX6M1UlRL4cikNF4ryI2dXH/E61RuphNAd7UY5+KT79Lq24zgUAjRkXtL51W
VflHTXYquXeS+GWeac9YvmJco5ADGMt+2yubymV1f5xGt1caCjcLcwfD0YGI6e3ev9QoGxj6L2dr
NUWh3VsILrg6wO566Qdf6N7G27nqGgeFz+vTJHXR8RaBlOr35s7HO5vGD6fKbXXLQl7eaFsidpbf
cZUGypdWNBDSpeLYX3ImRtx8lAUn++l+VZB/Z9ZkivN8oYWxajAWCNe8TAyC0nrgVSkR+pmM0eZG
kKGa0c6u6mIQDNML5mLD4CJG53a2XHSNZWXIYBCRemdZE4YZogAHg11b8zajbZhR0JDVxRQy9rDO
Xq3LDFhmsWXbPTNp/s6lT6yQpwRBLpf5hYuxP36of2xoWfUO58n3/lQXNnHrFP5pgdwccM8wONjG
zxM4rQkOuerOO+DzxOQT0llhCYBBIAHxw1/Smc8WQhNT3mvuthvJNw+y7/oe1Fty9Ov8Ua4GfWCm
61OcktrMnQe+RslHmxyOrrUpuWnzMsyYf0FCB6d8BmnWFIlwf07yqSYosOQD35rlYEZ8fYOyyTcj
+3mkxfSOau8bjbEtOEUb0q1DAAt0kkJtGODD+QvBwOW8uFeTzDyOie9WCMqP2EsFhHGsOMxMISTp
1IEyL5ZRTaW5cwZiar5zP/z2xbEOMBO4wyuSLSTzvMprV/qmijLVdf0JAR6Ygamwt12opDweATjK
DC1JrVyj1Ml7+cKt/Xn+mgz7qTM49PRMTriSzKDjCAJMpLDoI1mHhCZUGRZIhMFEEwsyniAx+qKS
mxTxqmraCi55vl23KKUbuvwGFUyTvcspXhQiexHUwZjXJWwifkAcl3ZymOvv38wZOiOld4wBGxD/
q5oNsqyCFk8qGeE++0iNdliJmqT3aUKN21iVrcY08a6ablAzRSXwXE/CekxANIUXyBr7XfwtUcue
o9LzbEBpSDlcVoC1q3yQp4Pl32QIWzAq4OS3RCR/4WHtD4oNHYkUg2qL1JG1jxZ25MKNQwRDErXT
jy1tx+9N7xC1YlSQl/Q18ZkRD8oDaGcbshnDkiNI2+wrY3dfgw1ZLSjR1nKhj1gUs8a7ga2AN0yx
auXjCjtOd3iQJSRZL2HEepgXh0CF/H1o0NN9QZkpdjVHtQ4VOrV0GscEkgoZPq+TnDVqudbmrwGD
Yny/J/RhwuIg8dRGl1CjoWRugkaJEiNKCGWklx7/ySjTXwFZoiPqa88AaFa2lXDrt0hWJ28NA7ec
hsXyq6Ju0l3wMEWJKU13jXXVRVesS0cDE9M27DNec3wJUuPzUbmdXsB0DXNovohK4MGgwBTKmp4B
dGOnfkwVNRK4SRtpUhBOcykUrD/mVrx7x1QZ1pN89iCiMgec5UF+0Qz66w1WiJVJX2njxarMni6h
XpYOTfZQ4DQolHxU6fukAFbUN5P+K8yiNW0GmwKa5q1h+6NPVeapRFm9wUHz3mJ5xMTyuWtlJlky
wZhPrQuZluEnFL+Ug4L0QEnCuYxQM7TfQyG9shSlZY8+2F9S9JRzw/a372rXdDG0QrWImlvqPhK2
xk5sD0fGtvtc8eQ94u5P3SGjq2XEOvcDbwbLtWzAIz8OlHvsBR79VPIaU4px0ckNfeVrRHhTtepJ
j1wm5mPiNGIiAeEBOYPJGrTh/fW6sUwJDZ37HDI3eiR0OPbAvF8orxRzIBuBDEQEd6rgC7l443P8
xNKzqf+RxucZ+Sg/7GzcuO4FG5vKgBgj8ttE1hOPyJqISvNpVUxoSY7LCCmcJpqmLKH26Tgen+/b
hQLQ1/4ZlZjO/UyHg20z6Jc4/lKjjg5Z8oENouyVfiG6+zYi1YvW8iFmnVPgPTjSBNZje9SBYiXH
ezXIt5NBc5BrhLDaU7UNgsKcC8B1EWqvpfNbRY+2kafII0j83s5+xb4Y+FwnfowUVLnsRDPwRPVH
2paffXeeHjPY43ZrJzBJbjZBGQSJNCCSqnhMdYPbvmAR2jAAXA1tg3Eo+/SWvpKH0NzDLrktQ/pw
znCgGAyPgUFxndaLuZsNK2mN2lq7hXFYfeuNB03kb+7vEly2kHVu/k6GwBUdYDAfVyAR7/IsxdUC
1T8gTV3QP+N1VkUfp1vwO5BqKc5yLHCf7jZSiVHXjJQ7xrHBCyLDJjIu7nbky6fWYcy5qSlwIVpG
pJnkfWAh1t9P1coOgkvsmZbH91IgIeSRj9cnUZJWIoYJUv4zUMpmTo9niFFLN1p3yu3a5DvOMeXl
ZFfy2mwqySdzhW4utg5XndnRQXLqEutD/YE30WFoDUJyCJvGaGH3IRJISMOslLmav4mgak9JTW9F
MlFjUPNdvb32Ljo5Ta1ZcXtcKo5mcjAB4QyuDInCmEsXiGt11KT354/qWDiE9SJHFJEm7RvzEGhi
71TKvvJDf1IsmDk3o5HAIRUqNk47HDAm/45QDG3L6rzpmsrlcfGlCx+phF3IC97nuud6w0x2+m6V
DDeZiAkY+czAIAC9IQJpKutgzs02Mpfg6UnRR+aWPzbNGaYLyassBk4vkJsyTmn8QhjiE8/ZVtm4
ijAPYl0gKgR9mcik9S0WgB27DTG2nQuognfT0Ws7d15+EV+mplL7sU9gUbkIM2wsfsW0/AsI6/dM
KSuEQaAVb3TdFitQcSPQa2dfknXL9FiQQmfbBLJhjKz6uMlI/gq0xfH61d44HED+waa6vHmkV0s2
kIH2Sd9T+OrUzVccz4TIwnSGb/eNXlN9DOlCqxWg7oWBeOJk752v0PCZJLQ7EgIlPOduLDZuXB1W
rsO0bjCQmJT9R9oGfZsFfmyAieOFyP2UKq3vO9PiVdtV0fhFz/oj9vbr+qHwryTZKesEyTdhzmGm
r3gjEkz0Ko7GLnbXDLNFLBIurbY6l1YT3zDyftw9k4MH2AlzQnm0HZdROK57cd5458jsZlKa0rsO
GsYtlhB5wOi4ztIjYQEh/agqaI8kqYSHnERKoBtfgWPkx7o+FVvSYOjCJreOLL8P341Ox0rSXyD2
5u5jv/6DGJ9A/hlMQHu9i4rruYH7bKmKPaf4LUQNjlhq2D9U4HJP++qqDOaIp4U+fbbLUftU3ePA
HLW2mW1/BgkLA1LIT6J3gY56vW5H2yu5m5xf+IZScn4kmvi41GYneoFjMLOSK6ZjfiNAQEedjbcl
N1RweQGo5fr8+jPWQeolUVYCc96n9tISleFRfPZ7dRfVzhjG/HM+LrvXXTOraLjOPUVHuESTNWx1
NgKGWQQ2iYTwuLyXxOzRCTnPyrWqC3B2cYLIs1hMuyCEeUXPbBEm9+qu6miecc3MXQBvi8+4FnVu
9SnynrqgXK5Q5oO7gM1mnUnc3ZmVpLItl/pPyOxv/NhAQ8TkQQDNQhZjhPZXlO/yJhDA8WM4jGpz
U78hLJrdEf6f7IKVaXtZzQRtRDpf0u5/8Bo7frS2WpPlKUWvR7j4PNy3JSVcgrOE/QV14hA248V5
+cHMRtzmSOxguGMH5cvDshASsX0fC3ImkKgdrAHsWcud5JpGed5aM/aQg1SZvt2Q6h8cDRjFKSKB
2HfnE25hwppWqBLkuWpjwN7ELW4LcnO4D2Wt6rDSmF11oFhcOoRxiAs85zwu4kTlgw7u4mMKmor3
kvJWyRN6bjLPnNQ1lEhcnXNgUvlCdEfEycYnYEhQhft+GZszn1sRVNGzKvjUEZHV6xBFD4uQTPFu
voGq7nzy/e53cbh9Yf5+9hWYDhzal4eh2/g7TSrzufgI1euY+ludnAJiVfOaNlySRVu9mMn2CquL
NEjaoB+Vq0uop/1+f2ClMF4ZHhXuuF4UJCrosp17SX1VRlsOsOoc6+h5OuP15Uc6CJ1fNxgy/mQb
pgZZRGsCo8L+BWUtZFd70MwAfh5habRtPZ6tjPavvA7zHj/esMklT65JfKKK7mzStdpOCAj8ad3+
2Jnq+487/4MZJYI31gevLiDAwJiy6gHJkyzOQDRjhC6Zdpnrr7EALfB3LjPWEuZ2QByJegEMRx5/
QMPunsq7xQy+8sIQz8Nqbjh+mj6FjCA5lghZsqKtUP60e/SQIH94iYWdbFAVXFQ+BgbPCU1Opken
B7KxFvVvxhuasIxeQmy+vom6QSQHdqRUcEx/RLx8MJccfIGT4WgVS9CkLUbLlLAWGJWXvOuqWKx2
1xHl1AvqdZIhm8Jx7QiIApYJj7Rkp8UEcEt2Z9+ALN0X7jm+TRMCU+gjIbxezDKXWvdpj/oS6Uxb
GjeahLgbq7mXvS7njVlQolLAEa3bj1GDb0mueNIAI+Casm2otQjCs4yzgaWSB+0lAMtXj+C7v3eo
3uVn44kRNJTkzGgA5JRN/IdoWRKIq0pyHai/pPOattVZS88DfCsgkHpWt/Tw8eeLcpT15nKwwt3q
/rZiIZFD1LHFxzekZI2eNLuQSNUT97RP4N3jiRZBVkubU1emzceewOxr65F4aJ7JWHHuK9mtgeLL
9nNcPf95WfpF0B6bgXl4iDSFpvbvFbhVal/cc0h+spBobRv18YOyeAp4CyIbBRIpfAmu/HMMcKcm
wEs9bhsqqUl6l6Tg2a29QFFXRTs1MSR3yb9xi1rVaV7GSVRJTDHaaN7R1kxgxutFekm6vTvGh2cE
bGr9wlZjhevNG2VSCbzR4Z/gdI27HbCUFHjU52nqbbGruWlGYNEOFdmmzIHMqoTS8o5iHNqVBtJ1
wQgGlG5WKj8CDF0Z/emolhNIvXRAW2tjE9998rVwRKy50ZWqBepnNfTMRyukWQIeotHHnYRTM0Zb
jAzmdRcF3N/01OMV1u2TNq05KC/fO1D77RYo8G9vy1/VhN08Ul7xRqZ3ARLwJIuddEvp0FACkk31
6kn3sEycajXIPVhsZXFD5yU0hNGjhebM7ikW8YxivoIQcGoeD9YnrsBdcmlZXTK5uzX/Ns9zXVKk
VpuTy41mz13AYxTNhAqpa6pRphNV3Dx/Mz/9G5OBDJAHSG1WR82BawraMF8QzaUBO5TlkQM4VHHj
ftSloMqpLADHcq4HuF8mxIX+liHH2RfK7Q1+7YnBQtN7SCM3IGEviIAWKaJsl0FDwZTnhrEuQ1k9
CPvKPGKauSm9s/mMbibgYr2Vdq48eu0fW33ygXm7JJ0F/85+p/dF8DtD2Yo4R4q0jHGSfkTbIXmc
L2/1ybCdUMyfUTJdclwrFj8itNio5tPwVKD6xxESevTIMo/VHgqeqAx9uzodXT2uDW8SlfZ3rOw4
0H7kh5uDjKmR+qyFrtSJYwbUct6x4sC25iWS0RN+e1ZMPfT84z/bn7PD0ykvMsFc/FE/riGU6OK2
pZoRXZJGDkOwBVUaD8bw0mEm8RPvR7ysPXlAK67aZL0HVlMxn9Ca8j4Fh84tLWSRU5djEI0ypsKi
1hBf5CvWvgr6HtzvFCA9nkc98inlTFw31WRdcpcajrNljpIayaNeFAbYkxLMZQlsV90luBSH8xNM
62DDeq1w1N5QiIqxAVgEl4UAslMZLsLHjNGoZ9NdLRHpFcJSjhKom4xTyi30s83a74xpszyFvloS
4q/rkl0BGnbnKfx6ll6vZK2q2FXkEJH4jolNf4v9VJr7E/fBxC8tiQ80Bn+CnWRaPWET9DQJMQym
pcPHb2u60eHmcLZgCVKTfbdmpD1/tIUUROl6dwakbbKz1Xs/nG9QSXEhF6n+KdX8pRiYRYnMAHBf
5wv9ffi7+p8cn1fyJxA1ZLdiWl4NWk7dYzM4bdm2KE6MUHxO0HZBBfc8lfmcU+Xzqv7dw1YRc+fA
EnRRoZFw4Jzxy8EIDXHjnnF6d+zeNPVpoBQx7xpVF/h5EN67nnEQg2TdE4jaI9jWTlHJ0r2jevKd
fzcyM0ssLSKn74u/zs9fBbmMP74qcEahfGxRcrmEmskKgVNn2KMo9llQ5xQIkErzJ4fjTFpSoAnU
JIo97Dza8tZ0GuK8+0m9BwMDYgTc0AT7LzEoj9KGypqiw99AsmacdQqscC1jI+TZFsvdDZScYO1d
AM+sGELd58JFgBdeG238rbz7/fstUr35cej5nl362zvlwwjopG2DgFksXV75oDRCVJ57Gpk8EAsx
eNE2pZN/sCWg7LJrgg+Si7gVEQAL0alxCm//w0iEd9/6wJYSyZEU64hwdMLh/6WrueaUKIqgB6Zo
TbLLsD7LaUmTMGLiXely74fOuHZAjBLYRW66wmrn3AR5z+mXy+6m7RxrUvjMIZBojUvv3nWwDaOP
IWeIl+G2MhIr43zk5Ohg+IG5AbfedNFwMvKOQZmaukJmKlzfni7XG4xRwhIrNJv6byN2GnyxRcKc
ZPW6V9WMnbqsJJ24PnfjpRLo82YF6eMG006dtVtT9GDObPTjmLjJsPkHB7Vl8O5I07XNi8lnp5aa
f9f4qmItYdrMVCiEcanPqInjM59DOTbeJfXZ4HvidXdeKWkSKKrCyJNrdE50LBD65mw0H0obWt6C
hy67HKFGmS9OEqdsmzo7QsiJk8PLgb+JQa/boAMYEHlsMnF9Mwaq0ERGPJdcSofyFDoAA3JcK7BR
qad55VyrFFxmQnfTH2EXW7DaSOnsVE4teOIqBUsU3J4Rl34VQpcvKCfhiuqmoo49ZvrXXKb9a+B+
ZacnkEdLt8bDvuSvSEJbkXalR/ONyhaZfjD60tELe1+Jyne0fmuB5r3rBxNDiD1EVk9TM8DeGsZj
adGQuK8hjAKZIDygiYfMJLORvgZ265fS27BR3o4Q7zkYZEScmMGRmsbjeWmXNuoL3ujKXk4daAjF
9MwbzN4xLxX5hi6MBF5wHI+8sg0Z9wuKiLbFQbVoWbfONJstLeFWLhlQJyLt/XIIP/zqKHpZ2tEC
MmrHkWYTzoudGt38ucYLs0VKNgUZrFM9dOLcR7tbrgndmioet/j1Jec2se5Lyhd2m8hraw+gAs2p
1WCep6mFz3Sp850E5FFepAxQFfXEHDxW0uq4OLdZtHdoUwEPCNPHsl3k7b639rUE7MSbqGgAAT/7
nh1VVzIqD/V7VnK+jly6iz2u2qTzxaRXYBxzUv6N7Vvr0zCFguXK2kMPPZN8qDCk1WlnoCaBvCR4
jrMOy1uwxA8KQIOpEBDx1PkOO4Pl89WGtaZPARShjEWTVCmeorQVQ9D0buUAu6rLIR275XXk+PBn
nuPoWMew+lFUMY5Ls9I+orMFro2ShUSPzPQhn8CRRWNPZ0HLAxZVt/V/OGY056UVIRiTf1Ns3HOJ
T16B7Q+mTtFlwKrRrEUTLke6h59SzeoYo4SkiXrUzeW8MosGfZSewpLX802Hv4B/Y5+CVsaNNOPU
DvtV76pX7uQJ4biUUY3l4f8C4IKkkqw5Nvstol5a3WjA3yAyr56Efyd4GlMPxD6LEOn93js6RgOh
4rABVys4Wtc8o+aGUaTbgQgNUO8MH37iySIjGG0STL58vmY9Lf7eQnImsz/mq+o6OW+noNO9dKKS
cfoX8FE0PzbO+apgrvFE+1pEwLwSHzB1JWyphOJQM/TA6LeatOgf9OZzVSE6qtjLer2hHdSEIG0/
jpZMVVcjg8vpgh4z0PrncPlb9+Xbd6zc+x2EE4MqSUoxbL2g+qGXgT1CchWb92pPhfufQP1jiTxT
D/evHOBOvTOrDgXtEvvcUxQLCQph2egwCOORniyVvQSW402biXShQ3SHe3VO8lkLtm6TXcSc+X50
MUsvn7O8QN2dEYHc0Vn99IcZ5h3YOWfHV0gkxYcrhLbzpxLDbJsvzGcztFymp57RPjph8Uob0goX
/ocDz3HeRA/wmyxoL/Od0Ly+4F+hugKD/66pUTlfnork5NF1SoyDuEZmwPmpBfhSKeMXhfkkkX3O
qCVMlCLcOjyJa7nccbQqX6kGqFxu/FYTOCImHMSfdqTaNthWA+FUqypb9lu1Q9A2Q4oM2bEeAtie
4etI1MFRgYDUlUyvORIVrAlLvZtIIUaAROC9kDfAqlGPwH31x/qp6FEY0KlWMya8H6Jg20c22CYn
+nyAQRLQhrrjR7ATTx/mASn4EOqf74qXafC/ib3q17upCpOuEJO3hmerXJaxaTIAteo2taPpVnwg
t87aF3+PMJDVEnkbO1sX0DOiX4q0202pkNiElxXHelW2hJ5Zm3lIVDmmc5L4dbomsy7wBjj2X8eg
552ZsO58K55mxrdlLb+WqLwlZbAnOV0ejI/B3+osbcftW3M/bR0Z766qRp6Ic1uM3e+3iOSfB0Yi
bpOgb1wySDC6BqsekYsn5dHQCGwqlmCwMZXgxNMlTL+ytr5sAqFLWIx8No9CzobhnNtrAR9brrE/
RZGMNCURWvytPJu0P3PBBs8wLvoh///tZ4JW5LrIu1iI8lemWvdyJ27I4vAnrS1Gp+H63gmOayHh
vp22LBkbMRZA6e9FiE/yh0sSVOqS+TsqUPYIXwg1ypJEV+7W0K0g+mrlmxLXHJW0o278d8C4qBDP
oEyWua4GLe3MEa86vXhV810EtcMm0/LefFSryVBFWLMpBJ68Sp3bV2Su+mcMG5Yxg+e8gBkjDoZ4
IT6GrMQCwiW27yNfEYVDXTUpIimZzAifAvAo/jDt9W0jwh7QiSc7iJ78TOi5COcLqZ+5ecmdRwg2
UcmZO9whPl/adO3jq8a8ROunqvk5QTGdZI9DB+g26OQ7EqXkYOuiTI7g2sLpreSMHynN64dzXbZy
pZqgs2i57cyBtuHu/GRIScdRvVWd2fnpkS3spAzyPu0PazzeCxqi+FX6QFp1jCDOTga1vbAY/JcD
oFhlxVBw9Qpm1JrCoeQWZF8EQOPz2zQVVOGVayxAmP2V3NZfRTCGX0uTFTPj7EeEPzf2IRBItCzJ
ozqNkV4zh2Q5VQnpYbaIrgAGZLWtvfrPmoMRnzipSPvGc41jxqe2BlHuOX9GHhDcn1meyEEtWnx4
fyAh6jzUmFt5y8OezJpgLqVtHNSfcj/7vqcJqJA+m0kMXxyls9BHP+UFQl55eg2N3bDrYNPegK/Y
w8cUq9a8r6NkHDBLdc22wB3IVYfCL81YI8OD5dLzp05SntezYLa4vyP3FLx/vXlzh8qQ/6coFgj6
aykP0xk+SdNeE5+AwBcbtFjbPpOfUYodcWDs9JNqu3OJKXoocfM0TP7sbNuIFmzi82MYAas4hxS3
TRM3Se3rJCydCF4koQmyAvASnhchrkm9rOAKTQu0fWvjfReeNuchgtgVG1z5eHpilyjgmAcvSYSa
lbQfpNg/VckGFzU3lYvU1ktnLxWxASiIpVyZXvmyIyCMLawgc8KX7ueSenddO/1Hm5vR9d15uwpO
/OMPi+H5tAxO6SIl/UMuz1xBU5QDl2paOhKcItwImZkfjy61RQJN1FADdI2NKLuhzD3OPQQd4Afz
bGb4sk14dc5BxLWLKKwDR9jefjKrIIdWu9UB9z5IEmwvDy2OFtxFypYV6/MUXQa18EBuXP0+Iq8k
hOi0TTtwV/2vpa4ee9vEgDUHTpSnpcMnJLPGgkQCBjVR2uJpQoNoXODgvRVSrKZbPfIWt80oweNw
MRojx73uJrdZCWxxIRzMoFwfwEO9itHObz4fgtI4ziIY2hiHK2xWOg6m4zltR28OMXVVSMY2XnNM
/XV1buu3EwMnR67FQGromazwU9Nwx1zRKdniKa2NViENbrauJEuzGaTTgDG59JYTDGlX0h70uK0P
BsnG2+lgmvsy00IKStIKxGyswCbsRznWjmC2x7t1We8La8fPO1onWWSXGd+EZxQLWqQBnNxGMpCB
MykhYTjnN7vMub0/6PCKW3jTKQIvNrgvggOcmrx648xJ6UjOahPBJ6t8WgnjTXZ1c+VKis0c3SR3
6nx6tEQqaBCKILVNVqtEY3/SXco/XVxL751EPjsGeE+P6d2+q2xdnOfzahtr5IT2qDpFc2FpuvmI
yAjDD77ec34qt7OA1UDVe9TpNYzj7DgMCw3zDxJ9U+eUbdkt+LpUJpTix6x+UITSSO1emtRfCUMl
3n01K0gMSc2chP8uI5gWVWF7EaPU5Uk9+wTQ14IDpFodwCZTP0a/KfaIT0zoWygScCzpjE9O6hjP
Bgi0pmXFLBuoDTkIxTpZIKPSJBUMWMoSig6KlXvAruZ7+QwrqcSv5NV1Y0nyxK56aeKJbpxWto9Z
O2V9ceXDGwheEgun/IZm82QRzYf6d/Nu6D7G9SdshI21yDlpYYc0cMQ7STu12oaT+ZQG/SpmTg2W
b/5D4FuuRNvpGK1BpaFLM1F7C3f7+lNxMq/dv2+b0l9mXMespJ0ANh0S25o2ehikXYPgGMeO+goQ
GhENgo4zX0bLXJEXycMnZOo7FucssWpTnE84MnX3yQaeB4jvJmhRZVp22GrxpF/9zb2bRRUNneGD
Hm2g8rBsoz/hs6f8b/STLR8zIZJ46Ly55Uu9vdnNs3AMr0LcpZYjG74mzn1OAfWYeihPB7U6kbP4
f9PcWM1Rid6tH0/LulqS5nRa7t97k2cKt7blYgOOWHQ19yihcbMuuzwNkn2Jt3ppGm3Tfx7LK0dO
5ESUOkY2/G7mjqy6s1lZIsdWqJE8yPfdpCrQoXFDybIoBIkd86fWF8eCrhLAWG5EwUXUcLKwfUOm
clgQZ4emb8yIywb4m0AjnrLx380I+IXN+AYK+50Z6kr8iUFmrqHV6cWbs8VP/KnY5c//PEEuBM9l
PkX4iPGR1U3n5SpCdryawtFcHA6wAkRwHu2HuC6rnIzkRC/NdNWVofC5NBzNpo5KDBtVKwj0loqK
faTkDLyTL8iMocRATmqXoWulQ8UNmI10NUiiLVeGtbR4EzeVQ4GG027d46mrhWrDfb9+HPHuFDi0
ewHkzlwyVW7rop/fFkg7EgIZbTpO2+Sn0pLJECaDYJCDieeTqaBodbS0XCCYGxsq2qyUDHoagR8U
GRlahLBlePG/LN0KooDKeM2+BzX5VpFB2DkN9s5X0Flcj3TM/GO/SkiHauLlRcep5vGFT1S/MC40
K3DqvF3D4PCU5KM5Bv8b4uFwAxa2FTPXhFsvd6sfTLXkinLd/wHu043HrhSDGvw4MQkEl9Y5eaFA
eLJE7zaDHKwSyoXjjDGeg7MHkqVEZDYzEueifw3NbPeKCSuCy5foEm8oCra+UqVKkAoyCAhZv62N
EMDNXMofJJSPv3KlTcR+9lqrFLSpq3CxvkngR76AzYhhiXTPFpFnbrFLZIExcvBCX63pb4tifX+G
zc5RRIH3yR/QQ3TMNf+x4l/ZE70mfQ6r6y5MqBVQilOfL4SxwXAO+cQ3EzOOcC6v2SUI8uNjrTGn
q/gugdBstZxHQfKkPtgRf4HRpslTwPcBXlzXTmsm3fUTLp0nTnpr+dBV7mfMvXOGiSN4LshNCpxx
XxWpvaFYRhRDu4yu1VL7PCWEdYJ+T7fpiO8Nvz85G2wE+8ZodjFJyKiA5aoVfjRtfjIMxTmp8QhL
vlI+ySClxE1nVobPYc862BKLqDsehUdXAax7Lyc25Ky3XFcjAaJPZ44n5xfkqOtlLtySegsJOtQk
86xanPxRCcnsdlF1M2UG+QSRtzX2MM8+R0QQM7a5kNOsfVs5rou+ni05B9u6HlV4pZJbwaGOhg24
i3cBPruEAMXlU55SA2x4HML3K+dIM0fb0rcYBa9N5qzXIfeLnBUSGrob0DBsDQoixbOdxpg9N79j
itaS4IrXZMRlu3qW/q1YXkQZD8mXE36OEE31oerLWyZV0EsS4C6q8F1cIKc0eg31eo2T4udE1d3a
GR3hq6//FPeloevcnsUWFFJMc6TZxx1cTTMHwaVjxawrBwTLeXmv9+GrtnRsY4mqciQ99FYse3CD
vSm1fp3b+AJjZlFCZ4tPZyDgZ4Vg6PzUowNpWGaA2vvrEHKA3pgfEdEM42OB0PNi0AUx0hZ9NGcM
erDdMcW434ylLemYVzglPw2Q/KNNk59yKdxfvgs0LERhMzAZZa7ytwSiQrAAyMOijpVWemo67aeu
Ikwdwzm8QKYCubf5aWEIiMzfuuUeMxSvMcmaNkQI2tKyHNXjkIoIGmwtdkiCDjzprI8qF3RvkugE
7TJ9GG3aRypzTx5M3M3BRCYamoFI7YoDEhRdW1nW3bgLcv40N+iXvTaofmgnHb/wP213sckUlu1E
oT5hSnnMCau9EAQIkEPWqRH7SLMwWWMxoy/V78Jz5u0+mcnAuZZNB1ZLChspUxODjSrf2+bYnC2T
JeXFB9jGbsz+x1EUE/nIe6N6jT81961vyoHcu8F4q2dDTkvUo6eZlOB2T1JonCQKsy0JyrkTn+9Q
mPBLOIYefwM+3GlgVL88wgRcRw1oqPYO/uHTNM11/05Sy0DQqb/+y2RFdc61OBTaqIy9A0T+zVsg
B6Fs8uxTzjMNiLb5ftaauwnTwdl7iWeaDZCzObC6PB1koXNta83JQkHls2OrrrNtrR+xgyhz40+T
/qnhgiRQOq4SOYFnHFWjcsqKvLojlglrN2AfReD3CtnM2GjNVmskiCK/ScdkC4PhXqc55g5rQBsA
LByHVyxZ4bOa+PCHqdaIb9ddZ6qZ1mVFVXENSdSC00a7Fyu2Bz/U3qsLaleDcvaBLKepVD8VUxLL
H3K0cOvgd0KpjbXDy1mDTB9NbzqwB8xjpjxxy6g95usbkisKzSbI2JII2Qm1l7fv9nnwFizYsNx8
o4EuS2MZElNWj3o8y6eiQCSMKDo3xt5s0eRSPKFbpFITaj88n7Eym4byueM1ESXJBPD2AJpjJIJW
noTgyWXoECkHi/fo1yFsX15yDhTw/6oRbXXy48LHg8RgWn5qYwHYYsY2snnh37tqrh7D/eSs8DPi
acLx5Y9nOFynmEQG9aarNdGzDaFiLDdR7za2FbNChtW1GnprGXm07Oynt3Oe5e71RGOGuijf69HF
e+pS4JJ+fyFAROvSOIIE1Kl7JipbkUKbkwR/0u6SrK2L5ci2MuZtS4/raLRvJiJ+nwtn/bmlcqg7
qECVtFrqhjPO7Io6vDtyivNZnRR/GpYWfm2SGshzw6ySII9mdXS6TqwVbq5GvUR+uCP98GrB0h1p
u0+68qcIDO1y/fjciXEBcVEP9FKRmPzc9u3TGkfpNvj3ZrgTNCzzuoB10GbZWrKSAsYx2OGUCCV9
r4srQRVJr8owp7rmz+HzdFVU8mL2GBpzgk0og9yMwkxS9DwOed0grRuP8JKrEX3LhmsdP9IY41mf
JdvolTs8mL6N4GuTtVuiQJXWnrn/0jJ3X5DEVEpdzSs2sylT7KpdSz2D2LM6HxcOjZXOokF0eKGW
F/Wb1I64EHQ0AKxk1QsI0YYTX409lEaQ/Q7CN/WHiKSUxHecD5sJWE4rmkvdOu/SddANn2ZmYIVl
UreitFeCmEAGz8g5mmAnEpR/9zoOwMEWepG/iuBRqEcGjUNhFIvppSQBYJFNKWG65DGE8BPuq6Ro
fxs99UFVdae/whBzVXqS2GUwvyTlLHP3QTDKlhgWKOmfjYiCSxAwY/8zh4O2JvfsWRbk1AmFgLNT
Y8AA1+n9FrHQEq7pfrEwJvF6W6zaWsnhY7l+D37dG9YfBMBGguT8IoWZqYmDFjCkYR8vscQl5qXm
1MXLeS1lR3Sq9fuZlNoqOJsoSJ5+AAzNkCFsgXBCc6k5LXk7usxvJiLuQYaoJsnllNUjQeB0WApD
wUImBEZycMvz7JHKNjvGMtXyQUEa6HPrNeYrpa7UFzl9B7qXfjEBVFySjSYc7jv+faOGZit7Yegs
NKKbgvqkzz+kDq07dOuTNObN2lkhnnV+wkGI/n9xh/OYV7foCp9kWRjAwoSdeNGiNOFGrxuirTod
cqDdz/omHhQsEODU61d7YVOUAmKb3jjyfXG8Fv/VA4OWI41ilrwsucJdwcHQp6hpgHB5hLL49CWs
R6vCQFHiLMasImKQ1I2+jrE3p8kZG3rPhIFT+VwtUYrsw2epdzZawPGVzC8F4Nsd47/2iGemf/a6
jurl2EvQ6cmxiQijJ9kYc1y5/J0y9SaAHZPYRii4RzJWol4itagan2Tt4jOdXuimuSQ2tanizG6J
Cl2OCIhJA5VP+SDBkn1IqcVOtiMUVjyX7tVQJTRHoMkvVVeSZ+ZkIRKFY1AQRaBp7ZwhqhgAzo11
JMIRGr/TpDjKYJHeRkuQelLmPMGoEQRUP3pApP8C7pvAtes8fdkW9o2VAoezd+0h2HIkk5N4ofDA
zYwFgxavYmATZB1Yvr4N+80CKZcm7LPcOIXc2xho2OrE6lZL4rsOJjKKd1q1UaAuQLEiSGfOIuAW
+KNMoBfNlX09ZUgnYpmv+U79djqfhR3C4Yhqwt20bXfGM8lZizXkMJP98TRIxXoNOwCCjXlntQ5Y
Wx97ghPiblX9k3Y5y3zXINvOQmDuNVUYK5vT0pAAS9vyfrhHdeeg4tgg8umIajmyutLCywUD0VeP
/eC5/XnjZjRDANi5a7xA0hYuPAOWve3fvsZFsOCkmtqBiz1nAZM3Bs5hd7I2PKfHFpXKP4QAUWSr
0mcjhTlmWVqpbxk2NIgGtRX+rdu4uC8j7hlhPbji8Is5wQdAgxloY6j3F4TlxueTirantRkY9Nfa
ntaUxGnsrQQW5kFJLOb8x4nRjx9Iy6e1b7i6OaWMdTzqXHXTPBmAGd5lBdXNMfNobWguA/g6MOCf
fvCNbReuyN1wAuxYHqzdX3Eu59Dh9v3IVNPazNceOP1Udbn4ZUBBxyhlMK2OkXxnUTCPPuPjgnQl
6478Xozocgl+w2D5+YqGHmBd/Qj+Kj3BLHsHtsOyng3R6+B6cYEP++XRmlYtfH7Y9PgB7LJArhEE
lLKDhBvk8bDtoz8nDSaDdXa1HGwE7LhhppMo0UKxfP20KszbmIT0MmbKguW5hwdCK6W63+LSNPUG
w12X+uzDGpiV0rZ+GDg0EcKqARsPnutq7iucgfnium6E5o9FwG91YZZE8r+FwSl3CBcLMFO/uoAw
8ZeASJWidhUG4/f+uU6vqV4Pa9rai/1UjDJ7UJ6ZeYUStX/7DSfp4Yw8XOY/Lk1i7sKU6O5B4Igi
XEVD3Y0tFx5AtsLtwZd0QcPcnvGCaQNPR7rDMw8v+PKTSCDNbLQCZbfS0fyjxSNATTZE3NRWklCh
nIznUD1p4FBeSQD8VeZ63w81cI+djcI7qVeWaQYQVEs+DrEC10TG0Ctdu+bpPBCeEUbjjVK8SokC
4aNL1RcQ8BD1pw6kxOHyMheBXX1qW5UM0xOms/BFgeMBHxNyPZIi91ePxUKnUNYwy+zUIO8mt1oB
10IEwUcLcRTA0zOePLRJmGTEJMKf20SC2mYJjW6lIoc3ufx8PEY/Z4HVs+TL72cQxiZmBoeSBaK+
ZbY3vFYlg3QweYF1aopWnboFn8wAowSmvC0H6OS0W2K5Sb6yMwLosXsUOyyAS9/JehTk6NZdCNO9
rRXygR0YKDDx3DeC7KVC2LlWb49l+qs0IwTcHmpctJPvEMzUduqmbxbVsCxv0mu/SEqhN5W1KOh8
gK2dVyUbigc9fLBlqU5cLeEwMg49Vpf0A7LHyhUdzNQpwHJM0qJFd8McaahQsyvJY3z6uDOOyLTb
36rJmYVpCLqiTLHI7iNCstJLdRF+Xkwtbwe8Gemf4c6LbpzkYR9PFP/8PuPYT8Eju1lehZ+8QG2h
vRfBKHfmyGbFSwhpoye49mye+bsIHhNbza56Mv4y/WJpy9oVdFL3glgwVgj+bLyzKAxmFOe2vCdr
YLlWtAxgeMrH0bMAJc6TxsYO5CquKCqManPsL9iMxtsUFlC8UBDpXB3fwJ6M/SCkTnHkr4wRXICq
AAD0B4OmdECJfBUQJHSFKUNmXmWsZ3V6Pol4qGf69SkJhca0I1raBuqrDDE6bS+NXd74rrRahnkE
TyVLd4sVpnPZEPMPKKQOh/FW9UH96ieubpiI4lOGU2+11/SEgLPCTPvAJJ1VFWb8rJS55AwV/Z6E
YmnvI9X4XiIyKHB70u7ZuMR89/RhLUIXJEQzvejggY/qQ2aqVmUnrOXKlhf0Pr1GeffhWLCh6Gaa
tRl9wzsOy2pbT7llNNNq5DuvIO+fS7h1nDyUNmufvXwjErcX9Mqff2jVXfLOLYtlhKLsPs3T7yv5
zSDFkzbOUsvfldktRz7EZWP/W4esz9iEXAlN3wtRCJit5QNiyM6oBlrfRKjXUdoif97SxLBwSuoC
p97dRtCvAkfBKwU69gga88MJ1Y74DKYrZGlPUtSHig4sifx6u6z0wPyi95ZWs/x4JAGzFebOs7SO
VdnpGd0yVxGarATPv8+Izh9New/ypsh6kVetit5AnUfuwi7pYXCc4RkKwpEIznJBMumfmD8kPTVx
aVXW+0jPsucUriCGXNlEQv+P5G7pcf5WpZJkAD656qn3dVPjikhnQ5EOTs/1V3B0kgVjK5LDzXzm
w14VeGs1izGK9yphErTCzWnO4W/xFsHGZg9ouUhdUaUJAlvKgixyg6XMdWtf4wThC1zLQkxyWyQa
VibhT9NMuS/UVb0jY5TAA0uY/haYx5dWVeQNdlfxkBIYzSmMxkFhdR/Xkb0riYd1ksglNqB0T+a6
88S4KKIqNjX1o0/oipXBpQ4HfmRVUUPa6RF1pDxN+q29SfByHZbMWwCQXtR2I+jgv+E3wZw3ylKU
GjIBrNkH6pRhB+cIN4MFmHp2pOl9Tn4SYTs0zd216ITv4DyYkIT5k+Ni3qGWpUCPYTZaUphG4Fp+
6zOvntU8IPhXql5sUjIhAIGYphVdQXG6EOrOQ5L35pjt5jV21xRcHPuN9UfFyjAzutgOa2qRCnN4
x1du5Wa4Ow/BUceFEn1wUDRNySln8wV2Nq3GJxdzcTKV/ei5R14aXYTM6N12eCz4b19fx9V02EXb
gQn1Aexg9F+3VYG8i8SXKVDiXXHRdHytEb2IzMTv0utzqTwkxMmTGJFmQTbV56w8Nvdt6eRhSQgH
TUJGIqI96hSRwAxUmKv0bEh3tE79NZzDYWE+O5xGUpLt94Sjxu5331N5Jzw+dBEOCt495j33MQSu
6syFWxtxpqiQvo9QdvlFp4fCEzAAFknWxnUt9elFh8d7OJnOAkWPLgkCAGNFpkSoNChFvrFfc3Hb
dJmEtJH0W14s9WGkIEE0F7alirpOjbjn9QkT+z4v+O26df7UDGTh23MO46K4q6iijbFk0eONq0Tu
nA6Dmxu0kKOw94c66QOHpJXWK/4a7IMN7hXzKQMdH8USJuGAtsfTzzLtwwQXchKAiX9OJjQdOtl9
0VNA3atdf92Z8N5E6Sax8+c3KI6sF3Mp6evCsikB+CQozukyGGGuiq8rhZ8EJguEdpSf2vSrRtyG
ijhUtxnGLI3pz1hp5PnRYQBM4iR1xo3sSjTNAwUUqkvM8gxHtkd+jvDSlOwb0k2UT3pDmYTkyeGf
LkBCWDBOTixb9t9lWda0QQeEg8C0D9YtAptlmNlhPtBJWeuO7KN6177TusyGjtpn76F52vcfx6/9
vcb+/EGnRGIVfChbwbhNroiYKWMBb0E6wCPSRL2hPpeEXfK9+yMlXynLWjIkRy/5NsMmbv6IE8V8
uCxTci0JhCbxVPin8kPvACCaxJzaFCRajNMb7zZvEENqN3D0yYRG4+xa71HVyQq5Qp43Ui2Mcx3W
KQZrP6CnZY2VAoA9y1GQuqKM1z93q1FbG4oQeyM2BEfJeEofQtd2TKCjBb8uBRoP05fKUhfVBBNs
WFslQcbquzfWsfBU2Qqqwo5Yt2O76CseKRb1PyHgy0J1fpnzjoa0UKf77JApdWkMzDZj7W8YBpHn
3dhP/7s8HAZdlWwTv1O3B55utHwO8qPozFckF3/pw5U79wWUUAPLcqk9HN2aFZMBpKPYEbd+kYDe
iW18O8lfoSIBYyop+cdR1QP8GhwLrxf7MZ8kFWQ0rrLALSHEOEzGrCcD58exd5w3TZY3zL4Mu3gH
kUReiB3N9131mmSmF1EsDsSFHJ1ylZyfYVJeOXf0RFgr8trrWG50M3l7SOEyVQGBSTmmFLd/lSGD
4cdZNcbSg9GsjteZb8+yjPYs5+a0tCeAiKEcMZVIr+9rk2ijX+PajjSJDxuj/Gr7xMjova0VIPUu
oBsTJ1z/kJ1oXgW3V0esrBrH2R6IbyeBi3bxSKtNOWEdLumJiwgExgsf+Mhj4Kvx4aqKWpbN/Z1u
9BxC1RH7Ws2nidOKp+kHIbfQctjW1zdkFWxE7OUdEdUL7MNRZsCOxRVx9QOd92koI684QuNfq8RY
ZwJXHIelXuS5DIQ+1Vi02cArrHfbanbo3wEg0tFTWvWySF/t3vMnRgTwX3iMSMULW/la9w3ec+l8
qTDowc9hsOkje8QFixIHM2QQl/25s63Jhfu7pjkqw4fw11xjNVlP8IPyWpGcxfPwnpgVbkkplTcu
QlMOdiHmz11WHhkx2TzgNnHvK3txkPfE/LK/06Ap7ypCHG5IVmxWY9IZ72u9WR7z7WtXMkHLHGzl
2D1Ec9Jcaq4EPZqW98vIFOrW9lWxeCOziG3cFkJlqluI4RXl03KGbYsdwt7WFiQi6AvWrG12UqQI
PAz2C6iAB7XQ3b183OEVh3jIed9uhCBkA8m42xN5cE5ZvrrBVa9q1X6TeWKW5ulPDKbUbJwqTKnl
AbAjXcjuNBWljbnhmqPf7uzEDY7RKtNZtycLAi6lsOCV7j/QX+aEOTs1XfAYM/lixPgFkwXI3RVB
apJBgYDB/OpKCyFPi3i5t7dl7Sa4l0Sm25OKK+Fp5WCtwDhJXAudunnerFv1socmqFlkgY1FB7ME
L9pG8aaiRzkqMiSC9bvUPRCfcXQZhLhgb2IkUZ3TRPq51L/ArXam5dfjMFm2Js0mPBYm7k6FKVc9
loG5PTGV5YTHoLYIgQRNtoXiJ3phK55dzeu6r08jY8JbR66X2I0wcE2VyIorEKOqnTIfq3iOTZhC
FGqxhfum0umuYdmqEgJZllmAwmc2swzDemnIxDV8sDUbooZrPIB6BgTRjxrn5BqyRQozxAreJ3tm
F3NZGhscHRzFAqPUry20ZRQNHFfHTCiWNh3tMuJ7osFk2Zk5pNr+zHSpxaCO9O8D9RMCGq4aJ2df
57gAr5KF0JL2s+juiuWEcoKkDcPhsMGHP2qaPSFHvUnY9OgPhuotr0ZVcYXknekThs1UB1wf1vSV
7kzXKv4k+5jnC34kbR658tzbATp2PhJ6YtlHXOgI4ot6qeOXOl/9FlYgIbcpEFtUN336I1TIvt0z
IxXdAyFSyl1CEP8Lwb7i+f7Qli1r5P/AcKfrFMBg4YSRD4Zt0UpVQTYD8xgl338AQu8R6kdtTeU7
wP9cyr2obDU1ag8SAjY2hk0mAyrferd2iL1ZrMqFgdL1mqM2OO+hYC9F4V/Lju9N6OIbqiZXY+AY
FrcIYPsNi1A7+u2Rji7ERpoQ5MYELVF6SJI1KBkFddrAFWlB1mzCMiKPzuL7yUrwazDglvBCf31Y
uYhuEaDzl6P/BQPHxoVTIqORV9W5dZW+831bCzBB8rR00nYD8AK3u7EoB/63MOVbesVQ5qqPskR1
4NJYL8uKynme8UtAHpB3tTaR/1UDRrnANEizoxhoAN/3DQ5ZeAbDvjtQN6GbGNRBbbUlkBp8oQlk
TUvTe5ZjKqrisBnpa7/Pnj3VVKVn4C8NIy0tq7n1+9nk6/LUzB6C6h8P00uTJUIUqMUAwJJmszZQ
vIPeJev4d+WDFRwwIbfNcZCJMgsJq0UD83mYFwRZWU+MHsi5BLzyhn3Wf4pNLtka8nrS9nOp5jbl
M6zkyDXc4WXd+QpbAe6yPbqbL5kLYnIbfCUJlUJP9OOThcTN8UOsERGUWuvKvNig20riRONhFrkg
ibJyMNhaLFKCMeuZ87ePIJ8fPVrlKZudzjasx/k9Mue9TbybCoyjBxmAymHj66G0g9eYhuHqsPtJ
QPKkw5kjQumIhxpskVIm6uomopctaEqaHOBFRoH2TV1fS6gy0kUN9oRKfEZifivYYTrLZtRIy023
J7tMv16OoxEIZzPFFMYzb2giDbH2z2Qkvo3DtgrQCcG9zTbJOfk4cmNdaukGjxZVA471IYrCTeAj
twFV6G382rM58M9EEFpDVeFcy+YURw3R2OsvGM8Ytl9JUa/YYtLH1q8zxkO3dibzBiWdViiFkU8H
tkDffocgu4FRGYlUVequoO08XKwqgvfJD7BqRRvGZShPSfZQUluwzslIxCIe+jbzoFxjp0t4eCCL
GUOLBu/2VVnuuflY5J9LTCdLh0srt85sKm4pis5zggY0qJUqy0BykwAP4an48SzxjbVxYBPGzDW8
qpAOi8EwyagdnYi/kvuDvtkeCTmJRzYSPsu6xfzDncwEbkDsrdytYqNGj2+nOXPzhdljm2Kif718
u+M/6XfJ4YANB2dz01gxjBxnNBLaOzVIfYGlsS8fACj/6txlv3MDZUzZODKXcFB8vH76RxegFbpS
fD7/OeSnJOhhAvCNlJTpsBPnXoO99K0slMOVJA6dK3rNk9QD8EfIqABTuHzZsDeJiST6H6/12MSq
6vZ4tjTyZASM6Hl7pQQ6maJ1YbeCHP6b/n4ZHXtJMAiH4OnthqRo61pkG8x8ZGUVn8l4fTwPGul2
YaFdydfTRkupGecJZib6Tgj605wWxIifit3PPUwuuXBThZ35XspipTtv/c/YMDg9wGdySihMD6Q3
QQwYRHt+zdMdTJRWgqOIOBgYbTiq7JZfhnpC6hIDX5PzJQtIDPlt+alImNhX9oTVxZBas64GfJ7C
UmVuMXvNAFpBRdowQB99jaHB8b5MIDa425uEUj6UpR+wiZo1MMa5hyIiQoIdEVPytIvjwp7y5A0I
KlKgejoCgY2+NtfNtIn0GkE+r9tqBVsdGqhPBAebcBlaKRDSyBpJxM1zdBJHKGb1OON4zKHmuLNf
QtyGktDPTUwXRSqQIrHm62DFg3w++U3oA7G45SK0itXEsRkfxZPINpoQr2KUQD8dc4pt06AlJNGN
sGGcfOLAT5nTDefVpP11zIOFiORL6CX2BEVAAISCjcqhps3p6fTMpbmVhvHl/2cajwGOP9jDtRCb
brXAr2KRD4MK9UkIQOVLJ1d+5thEwmHvtfvu9bkDq2SUjwspjDlhTjN2uQSZTJrYvQoqlzQz14dR
EjEeo3zzmDNFCwwSV9nNoTcbHXunP0j00Tfa47ApJ4qlPMKw2NMqiRlC37MW3RlvolelJAEVLHPn
bhDcVlTBBsckXRFzAKAJFuRtS64ZrKM3Ot2TOsGboqutRXb9MjHcwCB9RWe6lnzTx1fMTf90y6ji
581hCkeOM5GagZjQCO3cdzLRvni1LY3A7h0AA5jKx/xC+HWM4DpnIpchk0ctX6NyooosDwnaFhZ+
Mv8ZvUeALqSKEt4C7ucB0IM5n36/P6gByO7lmSCLmY8n5x033Z2YZ6nNl24xAVLllvJyxsKJlI2j
gQ1CHhIsQ9Q+SPYUsJl3YBdRlY6EadolaTc1UkYfbLO/pBavbMZ2ke7OKxd+tyiWMToIH5Hcttac
gtnzbsJ3cF8vy/2GsqwExQK0cIVK97aZnAr3MNCGm5DFhASCnsMAEXC5n9KlwyqIMOC3OFe49d1x
mZx4FM1oMbFQyLE69omTucY0++H11TPaO6XHOtTiGYuwxUJ/Lhk17ZpCqMfksgMEbEysF8qo71DM
YRceW9VTBllMj8lBvSnrhhzascWmhVroK55lB1bTUf5kzltFE/wvhiM7nA1PHceRifoDVh0GMUgj
GK2NfWvyLLE6HFed3AhbQDqBoZKhFtt7w/pA4NcVpa6zxfkkRKD5FkoqfMa553jXTUE04qAnFrj2
/8sCs5koUfeM28HZxRpmuBH+plhzSGo4otwoGXrdDYM86Am3M//TJsdO4Ugxfm5C1MjE/bznQaed
XRmBWPLt+kM+o5sXRplCE6kUB0UW1QGzo9cCMrK3qF6ixPN9FkWJvdtoQBM1vFCN78KI6mW97aKg
iWoSZ14PTykbyoVa84aLou3OeL7dqZlYHCwzY2N8aEcIk6NcqGJfUtSr7wNQ53CYKK9h/fyiiU0p
Smo7YgaRb7cxKwQyvSWwWQxxummzNEexXnMeId0GhN3UqNmRcrMtoHu0IKdIfaCk2Y1IdTUDSfOe
vIENKHHhs2ah7HDwp8/rlsz0Sc0kUbH0ukkgBgE6fjRYsVr90wxTx8D/F8tsQ9sXuh7NR9xs1FsX
h9S5Sz5vu5jox+SKpfPcwhDHnN6gfjykcmH6PenXowk7wK0JJvfs80N5/Uxg1dBcuQk4y16StZjP
fKhO8YFKHZqyB4uOBuOVDgdEQZX1eC+BCygoyonRa9XYqDJJMO3spH5nQ8nvj1A83epGtLgHNYQ3
Xjn6ikgHdxAmD0qLAmQ2+G5IahjdI4SVegs3Z00qZDP4jY8QbJKKKFnnhNJDUyJgJl4eD903F6NB
sulk/TD1OA3Jyoan1cbveDFxu7r5FgRNckl3nbsuSmWoM2qnXfPNkPtKTIJ9NVfoeO0VloD8SR+t
0zcHpLp8pmSoCbkbOtifQeL1SpvjKYfkwhz0c8RMFV9jue3IqkArwOcV88/yi0up0Wb78ufDY3vD
5hG/bM9Az43MDbCjYGsVLqRoCLOFK0zWqoYW0gQrz1eJyFvg8M5yyaNAwc6ChdYrm9YwZv558pz6
nPekypqCGqdwDJMJ+NxFAsllq8KYVOd1n2lIQ4u+QtjmYKlW++IYjp6r4wqRlQIkgadiCFvHlk+T
3eO79WVaEigZ2cBDRYQpWZhfE8AeJrhrog83c69L+VqwMRd3JAPAyGS/9ja7eY3lSPCK6aubnD7O
375QZol/SAjNtV4VzJx/QvbGf3JEs39R+G0W4e9iOIM05w0ltQIbVstbOVd4UaC5qmheD0xa0zt7
fuHNhO6tJ1UKpxkVSgEKZTlUoveohR+1LfRABJFkLo6TVHLEi6r4+1yLhWPWjFEFCy46P4OWFjWs
BxzijNv9dsdLDx3zYE0OCVeYHwAU7ftftW7s1F8/gblSHfnV3uWIhfg+HEOZEoSaESvMbxlZ0jNb
+W/zLCJPXCaweydQgzxkitdvIHZHza+rFJxncEqHVEBiJQeycmlG96/YrITb+obLfjNmXZ3r4v99
BPSen3GuhL8qaev78UEgbipJB2zcAI2ixDxIcPz9aWiCINfjjUhHrV2VNcjkJW1BumZBebMzxFra
XDkYU3wklDuB5yf1aNlg2CRg1Wlk39QQKWfqzByb5YESyhPitE0J+JfCC4VCdFOles/a6efQgMxf
pPR8kYglf522wKE2qYjOTVeIyb1Goun/ybInUS4E8QzhSM5dOVpptDyU3IYTy4UCiEWhKsYDhz40
nWXLT1xTXhPnA2l/7p5sMQ+vFX6Dfi0yBAZef+TmqkBiJiPBcnrVS6t6rYhlmZzknWqw4aHOHaHu
BDGV4k1HXobeOoevH7fQDCUC1QGSjIi+b6gkjU9HS/3gpJWbutZ9ux0N1uyo6oDphyFM9CPVzIeK
0gPOZKHcrfmahE8BBO+kkyEPPk+7o4hbvKtAi5s97wJ+/6Ny4C4eGLW86n40b++3DoOygvg8OnDY
nt+o22i4U41+R/eJxT6cI92q5IOm/bqNaY+BkHJZPcezr/K1L+/Zw4Kgro/hVCRnnQGAP7PO1izj
ev/GnOihxbmnNlAS6a0X4IaaqmlwmqifNMBDpeZBqtasqiPSY0Oow02E002KYKM/YYcADzPjkKye
jp5my8fZeWy7u0VTF+Ske4EgBs0KDmQP3X20YI6N7Cv11glgKVutT/B2XCF4vPFCizEgDkaP+s3g
+EcfPoPoVP7H5KKM8+sFMtrixfNiGSOlaIcvHOLHBENNr5vtmBtPRVK6Y+SiLF8pos/dL8ygc14z
ZG/2lTvN043e7qos8pGnZy1ORqGupGpnoJzj6YWz6GOlSS4Ozsjgfrb4K7XVwcSBAgoWttxXuOse
ZPrUr0XMN44h9/dMIDhVkfIOHKB7jpFNK/EVIjvPr6G1oQ73WbuBjm+MWl9zJXVM0N4qMicZuFfV
dbWaclCPlaB45VXKxhg/4kFN4F7SsPsdTDMkh3a6mI4NtiQcJlaULcFeJlj2NMuM1OlJj85jOpW+
wfr5PxTXDDU+zIa3m1AyEeESIx9Ql7xN5b4fT+MOZ1CD9ScEy/fqwb/K0zaLwk3CiUkXchqOkugz
SO/6WNQAVzc9xAs1tdM75Ywqcgd2J7qQYYXLLYglBeRDz8cQYMrlkuuGkxSSnUSiSfOXMWw66krZ
r1CETRpUdNXV6kHS4qOWGN+6yhOVPHE9RI7p9NUOxZi5aEK2q8B6R1YYaZYWnua12vXBf/G0gtbe
8Z8a63xi9V9sv+0JNgZjqhBRSFSswLTGbyUACndJT1uG4M9+Z0cyODOW+AZXwe17bvBi75gxqHgD
QQ6sydSsvgbt4v4Dl9EQvIy4GezrSoKTyh9ThD8dDXl0Ief6EvaPi6woosXd40JPcDS+Z4fRFyec
nc5pCY+8wxvHycipU4lDueHEnIOCOlYZ4Ilk+YWcYjDR6eDRzmUhAbOd2Svenvt7KrhQcDgXXZve
joUZsEp2PWBVeQxxM/Rya3vHXhFWirqccbgJ6WkS5KTsICR4qFNt9BHu45S1n0fjK+b2NS0DCh6Y
sb4rtdUVkbDwnfQPpZ1gpDwIP5IOg8jI5Go/xuBcfzfyIiFmbRysfMJZy8k0uW6mFt3GJSL5/jpj
nVP8BMVPrHuC85RdrShXgEoP/tvB4TsLx2wmqR9S2JVOyfz7ww7Wj5GFKVZ6B4c6vqfCv0AbT7mI
0sOlsrUQAGFGzviQ1Q/07DySiYJhfTU1d2WfyAmBV+OP6GvPcVNJD+ay+3UH9ajOT0tSfRNoudrH
0O8bJ+Vws1/R6rLub77VPmSLKjLO8Ucfd37EEHAiUVcmfAbuPk5GQSBEfiLlSmFq2x4LTIoCNO/V
gGF1ZriFQ6hJT+DDjAPb4tf5GWUA2dTMmNL3qpVzdvn4iXZeaMNYqHI2Kslub2dKf/o2EjM4+zee
7jx99mhRYC5nuRjcWSzPhaoeMmooyiBa8d5r1Wq2f0O94sIqQy/YHdlt93veHyNCAkNwS9pbhgBN
w8m6Ra9SbjNyiOFbsLudp8P0hUWJsjOXcFRdiMURIFfMlJJJ25TAK0B/HER514VpZUDWRhi42hWV
bElthoYFJbAYjVYFV+WGJcu48oJ4Bj3SmAgONbp9QPIE1EjX3+nZa1IF2i1zZrOnCnZrNVtH+7Cw
uB7xZxhP9NeGJeGVA15tjHqpeggGL3JoBULNHncx4PfyG1CcLrLqIRWS5sAyVT3k+gXGsb7AJa74
5tP3XSIeu8o3bxFa6jtT4U1YIL8GKwNPk9jolyXs89WyIb7Pr27puTDRRRKhOIN99Fli9ob4BMXr
57rm6ueYRBM+0BevXClkjso/5nNsCyRIEpF87Lx8oQfG+ta8C71bE793qcHZ6c9kHfezDD69Bz/L
HrggzgFUT5eZz2dqJgxHDzYMXJxYNh+Tn1Csbt927eq8np9mguXoEDodgnWb7eBXod86vRM6XnoQ
6UQEhDYDytGN27O23/3ne7/7f1FL1L8ET+P6cms1Ei5EbZ7sO9bE25o8PFW7ibr6yULG5tggBnqz
JKqnO1vqWuiyK83FVQEFC//JMqhFoQDAgRd5Ypjheo0W9ymyXXVMMlDJDXd5Y59wPsl/JrdNCAey
NI6Vjb6zb47EDS7GoLLwraTDV1FBw7b6+eGdKFgnF3RNozaPNiAYemfmu/+3dzrD4MRojJbbJwmn
I+833npiDz0ed2WB8INJZGPnGDlXIaP1yU25ZhPoD3phdUvjFuTZUy+pgbzxy4ut2L9/4ApgvZen
cUjODeWb7SLDPiRtHaTjEsqOkrhFNoyWjX/2qebeY2z+oh5+Wc1oFnOU5DWHROhNJNW46To6zzXw
t53E1t1gJICqOb2081ShiiKCbYUxhdTPyD4ns3sAQZcTqPXBZWmo4UO3qv14sR0BFTEAO93nU0g7
aRnMisw567pKP1dUZGkxbCk9nHOvVCdZ2QU2droWZrOWYMnshrk5cigtRQ3uDCrXKhRozVvddkLU
Rn71+/OLs6RAnV0XicIFa2K5OxMUKEAx/8EgdlBZophFTU+hVsuUjPQLPu1UAGDsmjccOgYsI7o8
GT2x0xqsve1sBOfBmjuCp/4bmK05Uwc/c1DGQ3LhOzy0fI3AbDJAkutCjsE7M0XxkgwV0DaZIhm4
uzXjNA88W370MoDMGghKVJ8LhWIN2PHQvoq40CbWq1vajS/N/FwNuk+u2dG4wfAZGN4hKguyJ0rT
z98qUCr5KXbEUfkmz17SETd7ETvbpmbnNXSwQzPpBU+TmYMc/xE3dJly0YBMKuNrurI3gLplpVYx
lfinadKMkY13ia+9Z3jfs/gAji1Wn1ziYPLtaTZLTMuRB/W7sTvbW+PxhMC7s2pbT4RhRiiMDyyj
zY45V0FUMRTBEAFBixu8bnuQBc6oosBD+nSbmtgNMbRUilnDeGS8U1z/m4CdZNUxsxVIe4BLd6bh
21Ja1oTzBCRtukKSJKtxMy41UCTnMcMeEuZdczI7tQ2JQwmLHCcysiI3anWN5eS6kaDXOLg/aAvJ
jFtBZA9jxstAnt1DoHieLc6TgIe2PPoNOt3Gip/KlnecyYWCfsMJ5NiaQBpn05mif/k5gA4Wrldz
o2uAxo495ffmV/DMDWpYTq2/mkOpiEiskcRsASYu5LQb0PEaaEG1JS/wtZB2XzW0TcDohZ0htW7u
9+C8VkNGawFyusBWHBM8HrAd1V3cENkm0kGvB6UbONyp2+R7EpNCRoustEQ9/2mFm6/ZEGqwyXvh
fc6K54+4FzZNP7PnOcgx3IhPX3z1Vm+WV7+vhIC/zyVJ+VjQYhY16VMAFwWS8rgkLUlUFF3oSeoZ
VhU7p9xW/E7QkUms1DB5PhCUMyBOQXd8EA/or1YASjlJhWvmxaCAj2wt+wFAI+BvVdGNE6VAXEzr
MCZSVUkYdsgYAll133QIocCtNKgpawlbgHCBUDELhGxEpqxE7n0ZPa9sMd/ptCDG8VsjzUPt23iD
PbAYX/fFJQrMlmpnM12fPS9i5t1qGw6eqYD0Dm31frHX55VFhaYNFBnFiHqqEj8p/rMpg5SpC5oe
kTetO5LXfoIO2DeoWgzitIY9p96IbGlaRzOKzPt3ZJ15cHIfto3H4qVcEckogES76JOCaeuNkC3v
Bk3ptMv4Bq770F86bCT2ee4GNN1CJ/QlP/1IvxXMZ6RWuevuzr2l09xgFBWhP0pdQRGY7rSgoAZV
jrVOxua59ky/TTn7lwSuyQdHuZSZtCnSkzOrIXV42+zvXrigtKu7HBX1Qeu296MPfAJtSL0eHNs9
U7hRSUjrxPCkZfBGH5PL9sqgNHifzo2V0S0cQ9Edk0GYEYC3Iw0OEl8klPRLIANXjrKMy2F7KRjb
M5ydFD+w7QCCVVqKX0peBnI1ZCpLMXQ6ggNUCNWDlDOk4L/KMRkyDALInD2LaOj+rMhjDlPPF5+1
uRVRzs7RHUuyidg5eK5r38U5y8mcb3SyHNs/Rrk21OROLNor1iGrFwSg39Lh5l3fETFb/8dgoTpF
pKQH1qJ2KO+BEyu3ev0vDefHuaZLV0rUD1xosMqzxxAvDGAFrmTF+AVs9GESlMSB1bIidIx7wM6W
XVKb3YvcDCtiHP5vX7onlEOkuwvddQLGb5R9w6lTJ6SjExQaKSxlmMXF1DopP1CabZIvb3YdtOOI
a7PmO3+OlZliYSB3LDhvtD8T5w5yWfRDmiNzS4JS/dMdciZK9cSYX1AMXHa5G4cVk6LPw9RoGo2L
RSeNH2T2FX7MWWBRK+TRbND5nPP3ePW2anqFe4OlHXIQ7i4lZo4EWZbY0fupGFr/kmfuDSQVL3D/
iLWtPsL4hjp4zLTQhJuP/6UxMsAaA49eqwDhmL8RnlAP9EInkw798yOSHx08iJS0w7yPIYCTBB1L
1Fd1jznRzEqETgU1v/x6KtEIFLhmW4L5OEeAGg0XGmhPBqB5uwW//PXphfSnFTIHcenBgdH3BqFf
D/cB73oE+x0XmR6X6Y3c1NrfdDiS8LhDlfy66luhvSi14fnqUEnf9dJFEhMOhMzp9A+YbEA616/6
Hf3dwJlxI7uULU82t5jPL39ybDkuNwmnI/c0GHLctsaJl+auLDYeoH4l3w+RIapQWWFZCX8WaYUU
7+bsmZTJ6cLTdc1G+mcjn+Hq/bM6ttb+/WN/41hyGvPxm+vY3O837NCCoa4louimqefdGyipFETX
J89oBpKDrxpZLnyJ42zL8W4YTNq0No7BJVPoZmINtDXnJT6KLm75Xu3WODf6lGmHYhyakLaVJo5x
N1qiP1DsUSLfen3SrZoDLVSfTGpeOaHFZMjli5xYJqENkU2cInqM5348LOSkvxvF8tRJYJo7NSmv
jc7wQ3nfz9md9QhdnR9kUehhdj3tLLLcPbQZBSymhpzz3MKF8V5NCNH+gJSD6hKoOwosEsLVuM2Z
CKAkj1hiK4fsPfE1l2DQ9GrWt1eVYZm80eusJ+ODsSCgPGBOThqU+9U/oL7okMsP4M21CMjqVtQi
nO9VEwNxd9dCu8osQEl2O19K7FkmLZdEzNTbyHXlwWQYRfc7q3OSxsq65C0Uc3eD8Ab/zPhsV7jo
CKwJecuOjgQ3CwDFTRXuxiJ6OlMM6DNF/+VpG9nvcVYoIdMI6b/GDhzhau86mAP6GOOBWbe/HLS0
RHRQhKZo3SOefrCr6JuKC837JWnkze8fQFsFKYa9Sy4523sqk7JdyuXRJcqa7M9nPe+Z9wZ88vY3
skU7/Gn7L9XDa9t3WQP+2rsdAGP/nNRJkrKzBYpCXGcPFqsHSKecT2WYA7KUYjm5oYLyffy63zJs
U4FVTI3yIBxS3q6P/3nMCSxbIZIxMjdOhFUZSsLd0LoLB5s4wXGhaa+7p1DO+vy52nAb6PmF0wVF
zUq99j7gcbXoOue06slC9lkXXTSkbVMoHz/5kN88DhOY62LW5Ga5KBxlRvPPBv9hu7+7Xsp/vcUp
MgeOHdCOTEdyIcxq3DFZguC7TkM9jAVelBVQrRfUNx5i4ofz91qnbUhmGQXsbuLpRS1LJBw6fFxK
TBpGHrxkqLIz8SV8ZgsGKF+VsyOSmonAwdbTiZI1t4NXbEVjuvV+6gYYYmCTnQdr17992E5u4KtL
HKUCUGTGtYbHbWFWH3SYCvp0cgpdND8xuAi6heMTnaUk+RNkYOwpN1hWSU3KmM/NIhwDFop1cFE1
bg0QFLNmSGqE6Q2/m/9KWJS+/91SuIlMcDqS4RdyomFqDFQRyBslMx75OBNYE3wU2zW8tGXDztrE
rFO82I2GS2YUGZpncNAfQ35jNqGWXUUAyZeBBISPWI2q+9ghZrEMfUiE+OPyOCHdIqhc25poRSYx
B7VEv1pkxpTl7+ZbUQzvJCAFP6U4bqfVeFQ1YNl3smluj6zQpp2Ng8P13LrDX1m2Tm5x/RV1pOjl
aAY7Ccl6RNgSg0udNeu/DdnlX8r+O0IpvQMqg1MWYlxD8FwsnTE1wrMaFK6PQEdzA5rKa1cxv+4V
zPGote1aeLA8HLBHclLdYs4Mi84/YoB1HYhWh/wcb5VLgGDhJ8BhRHlonlxjn2FjFkqYrH4FSpPV
/M7IHKoyEta4Qyp3T40rNnhJlEo7Z8xOUhiK+QbNbE/ZvRIrOZLxubdua/D1sQ5whEXY5OVgNX2I
Serdwl5E2R2XHiadObJIkXJlg6NKuGLrEs9GIWA7W7pppAygDK+VU/HhrATnYNSlfI1ONeWCAzLj
u4pUVC3SaYyok3h//OMWuk0XgaGorgghA+1JdhcC8I15rTHRQkvW0ec4P825tMwI8ZbBinIhwmb1
ipHnDyxHErnqvAUvARcDgy53vM9AqG7zvZQsQzNBPOezolKEnHLhOMevku/cZv21aH1NLZgShRne
WcCBVBXm1AgWuIEq/VwPvJ1dqENM95MfQEDc7L5QhirK1Y+QCZZH6T4S4XIWTWWv9HFLe3T8nVLQ
cbSZ1D2x4iiviDkGqbfXChNwDBsYm9FpRJ0LVHpeyfY3SMAMTTI+baRQsBexuCqCx9F7O6IAZd4i
SrtcisBIEZYuS5Ad3fzXW7XLwupLL98ozqa5S/gzGYFc7jvFkQe2BhwL0Q84OWNTSZNATos3TAvz
yVg4VRFT8NOavAMuVwfYwrpAMvdEabN8gigp7eBXoJjdmUWh+W+7rOcAbFGQn45qain23KcAyyGq
sPYdpSjIiYORRbTWPmB2dHrFPJ7eFuN0pfHRUJj9fQHsHvk0Ya+/EHVV0OYhXvZK6HTnCEQNaIV2
LeoHBZpGe5Td1kQlsoGqIC3Lw15CO/2Uf1+/zhp4Fep++KHAOBtLL5z+THLJNRaV/lkkRG0YXGBF
s+6KTScYlWBMuDGeyhWM1kmF68XDJhgrlPvOVDOey4wURcHbVNv1NZSJDKktzefrqToZsZaNhC6j
7XlLj6EWi8OykvXl2kszeOxViJ5uB0EoyX/PwtJnxGx2jf5MXCQwENX009XSmb+ULdAADJzrbR5C
0sO95VMNFGP1USViVNYdPK80pRH8YYufcCA4Hkt5Kk6itKYSh2qTkc7o4aEgqrCgBAi0z7zOJZSo
qfeXSEI/wO4QO/GW0UyAVRt+KXhti6bwUgVmYDQswDj2X6gu5Z36WHiEmvbuj8pCLO2LR9j4/2Qm
qbKMsMDH6rohx0DXu7Q8PaOXGrOfM3CJtjxJPYzNct3UAxcsdekgxrzoGKhLPU29o9x35ehc5q9V
ZJYz+YgXrtceL+UTnVM/iT7Wk6IvDRkoxp1qLFPP5+aHFs1Otl5ZHuhHm06eGJIy84PmPQe3z2M2
XquIC5KF5jci41CzQJ8lNCb6rEgNklDGFoQkzso0zGBW745xxVUixRVMjh0QZbx0VOshu2nEo9fb
Jx8ViBaLq2iF8azVaYZmLnmX+EMJOGC1BcovtZb7e8zK2Cq1tRsNWSArFeaXjwDryQMto7aUS2zW
GHYq/FiDKBAa4lLaed0efybxXT/DseAgtGcYMIcSgDO3vklXlUdpgnuNQ8s3FYAOyE8e6i8J3kVJ
9QXVrx3GzT88m/8a4U6r8bN1NUgjtwlEbMxkAQHoNihnkWJclu7QH9Qx10phpHurz3WxwAzsB/Q5
x1yIY9daL0i15DFo98oQEXoEcESm8NjfWbDC4ZZZNajUG3UTj8VrkyhZJFq8bhchkD0E/nf18JvZ
97q+YGs6jp6EMCFj5w9/RUm/dhA/+SKaRiH6xkHnVpFP2Y9UKXOMGNeuUIyeFaAQrc6Pf92Acyq3
LuQEZwIjoCDSycJcECOQVXg1Ds+tSbh+oiXU+PSnCcfw04yXTZ25DRIvSzqIu/jnjPYV5Idne2qF
8rB7ffKuljboivMTUlzEj6QLn2xdw9YivY6NdzjHk6LA+pTCn+ZH2hyhRTGvNDR1otoYaN7LpFi4
tmilz7DjhABif6LPSAefRbQ+Xnq7BMJbvcnkhsANqZMMRfUTl2TcFki/kydEOVMs4ijP920pxlhV
aqO+gfo2LVBVQPhS94nOq+Qd3vJVzARTvpUdlRgWuAfYay20G/2272Vsm7IJrowIzpMgqGmV1j8n
OmUaY56aSAUtrRQq29pPZOEoD4YsTi2FqAp2eomM0kI7YKh6Y6Eeh85Pe+XOmYoUS2S7Qq47wRRX
qEIhRRmNmKXHhiUEzHn65j+H+QuVPQ47smFEDS1Za6YGWeZExVZjyfw1+xaXZEu9EjBn88bBwmk7
WEZWD9rZwNPU9W9YBEAMsqutyYekVJZIba1GamU3YbJLFAEjrEZmEIbngbEGqoKUnhfhlmBsn8um
58XDl0QCdNMPHhGmwUkNJ0zaPki77nhYh6N01STt6dWnyu6uguStaR6yq0Wq3BrVictWsFB4dZn4
iPIiEbTSqNwnde4xeCQEQFCZYnbzYGBVRVEOjXGBrANyzHyneyCQGFvY8GvGWgbxnZVATg2LxexN
zmjlDUmciaWkcC5YfXilj6spRRU7fqGwxc+Sm0CcmTTKHHWADi1ehfn4d7qAh5fm8XXktNDsZoMh
pjqTryQdgGemOtmZQgPpevxPggdasZpsuESENOO2zIJjhrfjrersnlltBJ7pwMTd3tzVO9r4lhYd
EXjdDUNH1hfYXe78sqwRFb8NhZHzIT5FEv7LJ4lI9G64QD9nR4GK/lA23y/c8EvwipO33Gmh+BSv
FkTfGUn8agseQ5UGxyLDAJog3L+dcEvyktHWum9rRoDxqCWzzyCtP/UNovz+iAJ74C29GQKjYqKw
e5VF0pyaQEK6Xbx6PKb+RnM582wBVVzdxVAkBGipBomxPDPt7/fwaEhzJ5Hk17qbr49TLwhgy36S
v5z3gZRHIgGCXyKpnu5MxZnovMYXGt2cPuZBxkuM4gPChVZxLWfNy4SseGYgNfIGpxatUARjGGt0
rSvpn8OV39hvwbjEH0M1j89yV307KenOAXmiJfC4GjT7GHf+B8ZIl6YwtCVpTuBL6o/NXI92Q9Jl
oqdkORu9rZ1Epkcj0D62fcqFao3FzFJjqvt/vZtU8kkWfAvUJS+mOSjqdTz3/l3ZACtgmamkkH5Q
eS8G7k7eTG05hfTHlpW3Gq+e5WnjnCU6OyIOc926NakBffBy5lnaZ53FSK5W8KLUQsNKdGmUdj+v
3jju6wZ5XnG7LzKa680PiNHhAA3Pu5l/lUk+3tJEblavWTpFxtzmxUmEeeu6LQbnUBrJwjrf6dcR
0NOmr+Ky8H1qTvrDO6Qxh421nLvV3CfltNJ6pDqHGa28aOeNbsOqyUPAI9CLpIrhl8DiBzLHoCEG
puvMKaP77XOW0JSL1m0DSWQblGhXk8jazZe+rJ2TYCQAcsG/OzrtplVzozjN/w3v9siyhGcRylmW
CLyH+a/VUtBRBxLRs+VY5ML5T0FxbwBjyc1FY2BgVowJK3DP1qkgE3R3j6kTHzvB6OqiRSLXkqXJ
M5+nI7jADWLAPuPcNIquTmxnLSeUbsOkj868qjmPPGgpqx6f39Zji55yT6MS0/Su6VQQt+GDBe2C
Oo10I9t3LeO4jQb1k1CD8bAwOTMYSzsswiQhd71KrJahp6HjeHeOhVrVwIovihZpHeUKtKPg68fE
vSqnyJ1IBaElMxoUK7nM9skDZ35sLBrGsq7ozfMTjEteR31yZryw8TRd4y6Wo/PX4tNdBPPzOhEl
0+Amipu3DkoRggBeh5ZeDiOnosszrwAS8fq3jiTLrnkxa63CAB1TNlcqBNg8Aq6aDpbvVK6mcHeH
8HPRcsc1fswArIksZbaLH4Bhst6IrzTXAOWgeeyE2te2iKkKpzTGtmfjxltrH23iHc3lo26bAcx3
tao7VWZqOV0OTW0rxUPd0ch6exDkZ5S+TyJOp29vBxvKkqBDVVLVc1A83qs2YGv5SfUMaXyp5uWB
7ll4UIBkOqFEWAh1YJIsbti3uLj6yfbaprdvsHTSkhdlEuXx+rJSVwlMpwQzXd0b8nMIvWU3D4nn
dDY26uIFL/mD2gh40+FIZoG20kr+TNSVlSXhGnxkZ2MALvQ2tyqART/VP/v0AmWfyPFzRZYyK/cd
5htKO6jzhfbzHSn6Q1LZZsTQae1HTmML7iMNEOj/nkqkeLayLefGLQO/zHqnL1PasUKIFNTi1L9e
3YMzTuRcK+ZITHjPYIQnN5BteYF1Jws9QBcR+1ljgj8HniKBPcNsiBm4tvxFDs4D4Viidsdn36q3
YjqWkIzv+vJ7kpJTp82xCf5F90YqQq8WS7+7dvKt9R7cRRv53hTyIelGtdWfjjD0gQawUkkG5Hg6
mTytV2KxFNCnG/EGDPDCgnLWNCvLmuWuhUHCjpY3T46A3EGhjhk6N/dGeS+uvgVkVXZ0TNACK6BZ
9NuaL5lr68ihg12PXHw+ja29GyTOXC2DrYwMvNSduLSLI5UYWE3AuXDLlWqAfK26PGsNDukhv/N+
DINhcPtgrrebCPG4Ll+Fpem+mbqF3FkVf9IhJ//fmzZq2sRmlDbbo/F6JCMmvr0Mxt765FC28T4t
q4aXlZ5YgO/IibB+BIc//OfJQjkPkb/GxEiPRalm2jZZy7+JuS3bDCKWH+1u3VHCaElQPBzrDhKn
vvtoJW2yooTzp2JFkm2uFEqyhgZUqQYIqLsh4gRh9QahzwlBqmP3Rjn4CDwClj5kaD9TRs3CXE8c
p4TSem2BHNVZ7AXx0rVhvNwgkE55wAufG0/8DrTW+bXjy3oCktNnlJ3lR/bbh08Fhum88/+2bwFv
M/N/jFaWmk48rqKvsbU4yHpCInjSRwvdLuRTa29wfZ0Pr+q9kcrRuGPF+NV1IzDjzff/rumhIdfx
J4Ld3mXkeS2UgZeOHSaN8yLJZJXu81RfI3swcVKLKPUbYD9YYerUvybN56GTrZ1CffW1F9xMw+6x
nG+nKBnyppGKy6MyKxKHl92bRYnepuSnqCBIqAQ8FP1bVUXAkHkkxrUL/YULylSqNrSfMnAC83IC
NaYye55XvlY3JpPb22oB3aa6By3ONFUHliBt6DYGdmwaegQRYsgXmDFbD7se7VSYbknXQ+03nYUi
egnzkm1FfAVH8KZaAMafloVb32u558NCA8N11IShAO6Piw9YOeOw+SeQCVNVRb+hAiZS07eXXDNQ
alLtmOo7I0faEl9REdPHK5Evvh5w/RIN4G6MYoIPtbhJbmm0dHTz7/c97OZKHPnXGYQJVFYsf3/S
TrwgdhmZmdmbHDB683jmfCvnu5W8am4iukQt9SnuLoeqMM3/BaG41yYgnOCBaX/PaJC2W0JdZD3w
67PdJvDB+TdtYaNAW7SIt8bTB4Te4N4wUdsPpNs+jwRbXOS3hLfo+kbRI3+8S0BKgsmYdFdgrHcp
Mx+fFuXs092xYCGc6eYVNizHIKrwFvOYxjMIKV3ZY/sSn3VSQAqv+FI9H1ZpiUet6PjwsgEo+1ZS
QWraTqKfBQA/5jxnbk1E4B7lViPM4d+yJMJdAwP05DtVifCTjhP9Kfe3t8yXM2qTRoAm3mqrUnf0
Lfg/UJhXMEbRsKhpLXhdnSREm2DtXCTTakIgpEwMHaZ7dpJXhpzqlMcuzbDaNBXyqaEVG2aabT6j
PPe1lyOOYaRi3MB+0AiDAewlAC3ogFFnarSJhMinG4b9zXh4cSyDGXJ3SVJommUGa1uuN1mLIlhc
ff9fSGy8m94YTsMr3N8MPwH/UBP9Jea7VPwsOL8Our6Ul3ta93oPEutLLxF+SGswmQlIVi2TMTZQ
xMBSbiRThM6edz/ywo9K2LTreYa7uxdx+Uv5iB/pKcaHShD+BxzfQOHCDl39nleKUKPxj0uVc+I+
KAR7AV8HtOr6axV4gQTKbMNEC7pB7QoQ3QW2muobVGFVvNHqyDyMmSol12/9WoW4k0fxFoOqRGD8
t2QK35FwrKZmBon0nFV/uXQxtzUZ1g/OmliqnsZV+DzaryiAGH0JkryRNHT29DlacXR4UioEXNVW
1alVw/ewUWLAIbaIq2PRlGWW50AObH6Gvfo2oYt1P/+a0yuSl82FnDepJURk9VVP2FeW557tybIX
xEIrlgBD5p1dSX7yKT8bJvXVUrMqSq1Y/stDGra+IjVnc6056xlo16GDWdvliDxX1E2/JoGJk2/s
7bZzDBqvAmveTbHRHtx2ab/Sw3TeYVNRpWQcJl1ujLal+t0obF6ueOzACYu0y8tXyX3n7OHDvGqU
JB8/QTDrqWJfDqSUjF5DHdU+nPKtMr2XGtJeOW35e3/+rOSckCF2QHGxYVQ8JJb9/vDKFqDDtJOX
o7CwY1tlGpSbMyjh1uWKJfAPzqqITyGmEg65GFIODEU5Q267GxOMTAot1TVpyosDkqoCPd52xoMA
Clt3l0Yym2tTU8+AfhI8cf2oMZM+hCi9lHqA62UvhMCfVlZPp9p9+ELn+SAy4GQ2ic10v0iSBS48
Bw6gxFCuXW16IQ8KuFJpW/c0WNtQBdHXZi0p5VKKz7YJZHbs1to/PUSXw1Z2nv/TPB8UWAHT0yZy
TOO5VAofGHdxsdyfvt6ssGSGR0ObUIkND5BYgwrrjFxh2tOS8H9kepMFelzVhU3LCqhShuei2Z8b
B1Z7jgeUmUUzSVYwniirQpGS/lGqFRAMAL/aRHF8WgrI04VTUZJQ4ASwR+VNVekYvrj462aoR59G
ty1Bg3Ar2i0O0HoVafRltmwE6QuFoqBokB3t8vRNrpMkJTOyL+tXL1KuEeZf6Q+JkdZzMCRu8Oa7
pBt0mq46a3KiU06qVlS8SRyLQJ0ti4YPRErsPz+1tvv1UJZeEjM6XNxfUo5CjUskV6wwH/pRvnNj
pUzb71dJy7jhTHGkO6OA87ACiW1O98Ui4qNMf3Z5hF5inE2+A2yr5tLk7pbhFyxTyoxm9b77O0cG
fp5VI/SNDdag9/GoV7YS+FjyqlsHDFEeDjGWktzIN7JGIa8UOG971nVIsbJWSS7iYVDT5ghzaSd+
bpGUzRAMZ/hvO3ZyLDvpteAQ90yYc3XFAds6cIph4701Y+ZicAObU3hk0qGPu0/gBzUG7DGI6BLh
oVBohYOnz9mUJYPTZPM/C8ARjZM1ZENgW6I9WAbAr0oqzGFAy55aMjE3QlWS83UGPc69MfqCqpX6
RpW550it3QKPEgUd0n0uX4Z6NvR/6Anku+s4HXfo2MYfRn01fYOTqrLzvVezsRta3c9xWFJ8o/c9
VVPXo9f28uQwCL/3OKoOLJsuRn5sy6k5l+bUiH3Fe0V6srGBYBxYZZu1oxnNiJahKf1xmJ5tn7Wv
M7HLukO3pJmVcL93k/JF8DluWyCZ8zB2BYeWe6MzXPR/CRbONm0IY0tUXiFfbZQ2l0imbJ+x901l
WHwcgtJXZy/XdjjkDHzHcTEmFLFAFybUUyp22GWqGYUBwEQGJjiabNvRvyi6I091NmZe3ZSbHt4+
vAfdwnlu19HO+qMG9bBrxpOgcI92zaNuP4JBfXUVy/TFnP5v+vtXIazODb2HBBDwIl5O3Gb9BBJo
oBvRKjGF/7bLez84UG97Fvdo0xtivNPVmPjeI+rSFSRo2J3Bhljw4Ho8siVIYWRHuVlmlkVx/y+M
tbnH153ptsMeHeCrfIANezfoBXKc2taBTKme1dx8wQ9wwv2OXDg9mVIZNjsaUkkA0IoKm0HD0pxt
kOCocAm/kS6hfVBB6JPsZutFHzZ7To1rWaMRnQelBEojADxA4htlWKpEmJaHros5BsKaAa0ByTCp
9tJshFkKyWVPE9V1HwASWbNDzeEDdPB7jyaDEDqvWyj9hCQssZDSDvpR0Sv0H5vIvZqgDZkBvksi
eQMumvapLnQdjSXqb2Q6Mkk7utj23hLQ2NmONBDnZ/RvkZsdHidTaiwP9OmdGPPxv9VdXDnelPFz
xExGfK9XFrA12b+Efiy2A6++LB85U/csgqmMBN4ywsJdbMW8vYlwKYlSp5rNW0vMV671oqopZFRX
GXc5Y9jJ02ceaHmo7WqRkpKOATy2V6ruoeO4NbWm+T4GA1renYtMHUNRO9QDHA+/rjWl9vH/wJxT
/HslE4b75539vTct8eQL6V+1bquC5Mh+AQp+4RDIMj90oKW4pMCNv0t55BzypPhFNV3tkjj2sWg4
wDas70mYYCll+78R1BuazDAa9eenn+U8Nx6+SZqo2A0TXHKn2JuVqjSxeEd0LD3Y4Zb1SiRDWz88
bBk2uDiAeEw2qMiKwBmmOWkYf92tf11nKgjwL4t15IPhcx3tjPPZhtNw+WnMIyJwNs6qv48t3sYn
kvCf0cLVxiHdiSyGSCpjhb4nupmlfpUUBO+s4j3FkUU22sDOGQoxzHWliJgYze5L5/J2PSI/m1hB
eviz0uI1FbjgNEbiw1sg6Mk+5QMs4up/Al1vLFMjujjTMqm//ekLhQVAxFcKH5EUcX0SchyzLWVy
xk+dAKNl/pQWbzo1LS8zP53K+hdMLBER4I2tBcIdR5f7WP2O/Gyzl/6PdZ8el8warwq4cwyh4VpO
AEK5KmLm4y4DZkCPsPa1wux+yzRGzyQWll/MN1F9aCWdtxBABgDL0aIrObDm/kTsotLL7jfWGSjl
s0y6C6HZPedDe9/rMdErhL3LYEW5wRl5GufNOM4x0h3KOuXisc8OHVclapAcN5DqW2nZEb53xrN3
PE0SY5y69rdtOoZZKw79VO7JghDyf44RXtIZrUFwAYfZXu1b6vAvGIYhOjiISm/tduWqCtDLim7G
7ogohwx+Dhcp9uryP/pXr0rR2SdvdkpjUMBjX8GgmY8qBjYOIROaTvUqreLyR2WBEXbxmUYbcGQs
nHYs1MPDR0pwxvwqwz+ORMaQjFi6TRI6qu6I1zSyrE0Bq1bJKhtopwnvz9t3vQmPS+W+OGfW2zqV
NUoiY0lRjB36jAZ/l5NgpnvWuRcZfJtA/BmSxR2TYG3EAOQ6wn9ha4CCg1F6L5J0K9Hm3kpweVLL
8I2viIJ/wELYPnUUDC0FvhFVDE3Gw1xZiNllP4puDE1wjN8cdsu24wjihhVzxWAZfddIlpeDZuao
qYKU/tp/vdvraCh8MB/SCBFzV5XXTHaCz7vT6t/q9g8d/aOSgqattDvrkxc+X8j77EOKYw7nEQUL
MHa03KuQVsmD0UDHV/GemCnIUkpnbNnKzYkREGTY/rm0H5la7/SzPqlMHbAICAwyZV7IYVRjOumD
MO2G/yzopbB6rh5gIABFdzp5VOBinNwlJC1C9IO1ubOy6nljGJa7Fyis6grt2FaL/S+k08jsbyOj
AY6yLt3o9wwMaRYgYanAjdwaiT61krDpYCWlP4fOXOgD5voMx5V/hFx8MNYnEhLLpgUBGsUuCopr
kk3ZIOu0cVNPZVofncZW+wYBGv+Bga2R1wprZR+gWjt9SkYx1LDFR48gFUf+FuZ4xVDYl92Sxb9l
I5Ev7/rPhOouYGFEpwvP0rBbimwSFhVURAzAfX8Zr92GZbSXXCBzgCv/kUjanvVjYRZrX7/+6yRi
LbiYUDa6xTfzBP6W4BZ/J6vy/p5P+HNHqq6IdXrS+7jwykwgF8m6fNIn2ocpX0fJbkaPxAejVpB2
IyDowrglgRsxJAapdzn+OVvEESfRppAcb38QgHdUndG28G689gx9lEgUcojqgZQ4VWN+OW2Gfhnf
vsx4A8OYUrYyaqCrnDCpre6GMXTcxIzZHsQn1NwO/+4sNWK1+kYPZ09bzzuqYlnxeJ9cYao+likh
mqQeSIu0xr+a9FcfiAz7tiD6VAPrfdoEHspfoqbZp/gncGUs4GF003pklhFFjFpalPTPChIfrVgl
Rc7XFbpNda7hCIOUQCakuABsN6gOw0Mz+9itbE5Bvohj9dtMO5SVBjTG1kthIvgmrZdEObmdxu1f
hlpAMPSZcPsckh8xV4hus4+SYe4twVXKuyyglCKcxWl8MfBr/UUmLJx6qV2B+obps5mDJ487uoTB
TBqBEIl8VGmXsHBDvIBOGytgQLHVfaZ5hNkQzlGkD2bXbjj3euA5fXL7X7vG0PB3+lV9k4FamLxr
zIPHwHwFGxqiXbP98rI5bbWzQomPYtAgEFwhX30cmtzFTtTXHp4IqtPqVcY2yHmZBbboFDFgyPc/
6TgAFvqhbduqPPvLwtZU6Ixny2qJIf1KpO3Zy9Y5eou7PuWvBIYYdvtOyeUf9prdbd4YuYxjC/bN
44w6KH5OZhVw5IrRpfpLcoXd7UZ/jwoSR0/1VP2a8Vwo9ra5HAd1fVc/goHPml5LEpqFGRe5s32U
cvWkrYUfRlsxJl/TqfZnnbk2AlxrwM6rPjxZ815IViySq9hZW2PhTSEm75X/vLPGqaCymaUB9dbU
LUPg5qFltNsmp4HWx4NTka79e4LAiv5rMhpBD0uKsMLDF2mj87qpyaGL8G9Htqh+vFSPuX4UidIg
oeCefGsSJpWuHhNGRg/A3LHyC6x1FK732QsbEMdI6S324/VGxaRSZj7NBqRJLn9h9OqGNyYLPTJD
in0Brr/xshcqibNk8eE3poPLjJN4Iz4PTLDGzXq63yj9fiWIDrf2wbioMsVaBpRKRVbY+mc/0cOj
HxnJHiGGqI4CR3srDQEmITTu+1I9f53Zje+8lAj9FZF+rdmLm/njSsf8HC/392IpnjaPH7JYONnS
25wNBVwtBolZjlHI3sJ0vciYbIkt6mZP36GwA0PFNaYGGFjnkvmX4FTZYraFBY+ougMceIq229q3
PQIHuttxH2/f1LIdhwBCOPeKVtF+Fvq/P7uGS8cTW/4rYOWTEMCb/PO3PcJ+ohEb/Vf1EzfShdot
uaqclHj+HSbEoT/ZNSxfW9YGN7xOYNv3q3eRKpa9Xp8LQn322eTTitvcoXq4MTK4AaOODmodADwh
e7Umhg5QHQM2Yc/RRxFmZ3JDgRKQt7QcwVeu/+iRa71gWwM1xJsxFH4oqmX1JR+SlklM9V16fYba
/qpp3dN0Ohw4gtlTRzTHsFSrK+RjI7ozbZuO2kSd2Xp1QYLLjhwhZdKb1adxCkH6hqANIJHitoSX
AHQ2+LpYenRsfzkuWkiQu5fCGOsBw3glIhtHLuR9IXhQyfEErUjnzxkq9CJMEkGYehi9f0/fOreV
a5GaPHEi0piF7t9rMHBPcR1NP2eqSr5c/R0unH88IIDs+ZwYbn94DBghJIUPIownEuDhsbcEAZ5u
ZT1iZ070LwFc7tupig/37BGqW8gWlTpYar8xtIFcY3XhQCPZUDU1Y1Zgwsl0u9H9OOlbFdOlBL4b
3lsPEQrZaZaghq3AXYV8ivyM7NtoNNfLXmYq35oz6KawLm4cjaAX1yEL2T41/6hMo42/IAZeguKl
3dO0EnvKdkp8YlNRYpZbwFWpiSdIlxiFptvysIn5F3w1YA5W+UIxzONYADXDWqBXY5X8ZwYpiF6G
PD7F8ympiVpQEXd7K0hftO2GglpEY7SOEBfHrRsic1J5DniW5oSMordBStu/9m1D2qBG8JKkRI2K
xloLS3M/sUFfwbICRFTTo4l2pzB5Z7Qp3MimLOdKCPbaKM6Zh2loF8spe4pmczSELXRS10Aw8OGv
gSpyufRZK6woW5L6OSgo9tbFexnXNvvw4Y5EaNBrF/uhj6+HTFxyLf3A9IKSVJH8E7265p98hJr2
pACkzqJebci9+ms5idVp28n7huSshTkC+P3EqMq0STa4wsFPcVcSt00BUFFImUImDGkBM20J+tl8
8YAeJ4fOjDz6DBUGVbUGg6R+xwqY7LChf1Fthrc5uhsSh8TEJkq0XuGV7sdseZIUaClCLntt0aep
bT7TauGh97QJEh9vIOT7u98jp0R7qP/ZnPxq5i4BrFtCKCEFTd3PRstIUw56dVBTdoRMEOPvNBBQ
bkENrsbaQJZLUSj8DriESLjziGSy8bYo/VcmXmOfpxnCqEXPEqcls2JVmHQNZklHzphVDppppfXj
GIRJfFLQ7NhwnOWCGFlUVaUFunudjudpXv+CVeDClYt6TVG3AT88L60f9Qod5Vakz9H2wBrreoKw
QDpTal03i5+J9LYqesM8l43Z+TnMpYOaG2vYaTdnk/j71GWK+n0LERr8bci4hO1TecB8EDk5w8fR
jGVlqfL2XiMFiDr6mNqd4q5d0Vh/3K94xU8WLKuGYprnzeNguvwq+pQ98FUdVx2iHI3TK/Gt4OWx
g2PJAOTz0xKivpCI4dRsr2FQO2Fja4ibin9FM6ESCpFMMXhJn5l8+T9ntq22BgxXfLQ/w6egON26
RCIVJRw1q7EBBi/96/vk8ijtZ4mykZWlR28Ez+3csKNOj3/nW7rlzQg8doqGpch9uhUOOc8EcCYa
D2ke6CpitQNI9O3fIbnxOrEhVOkbAYfqVkx2ZonBcB8S8QAhVSwOeZskcLe5E1hIhsD+FzwSSymL
syHYAgnZkpftTi7H/tJJb6CkO9trRkgNLUCR2WTs6NrCOLzXG7Cm07Pk6vTO9ZV9YQyfvWV/FgSR
8P7lY4QY6WP2CdvrRmX+iIgDaHeyU5YpHx2ScjFX1Q0DOKn+9tICQMaXonw8YR+l4RWWrGfs2KzL
V9EL8yZK6OdsDgzwfteFJYKAIOn1rI6Cn0rw4jo5snTY98rPHOTLgEBDx3gltywCIIByCOHthqkT
G1eL3NGqLkdHURzChTgTCYNWrHdfki3osSeT0jZCsPsiSAWW46L4W2sdATxfprcv33d+5fuRqsSP
5+cHY3VsoA7MRQVOM+Y5OXotQDdWpFIEQkxGuDl0xV1wYWBS+mXXy6KG0H+R8xXw/Tk7SqBgI/ts
KNNaGcEpqkdm4ZlBSLvERojc0o8eE+bkCpeOWFHO1V41BlXoDgC86cJwI6LqoGFQQ7Neb/cP317K
PgVGufP2d14kVkP/YWdeD/CJCngr5Ez9Y/fpkXXG1fYG02Jpe0DuHdnmqFIuGGayq7IB7vUgB7Wc
PXpD7VIvJyuFdplXIJKlEPj3aoER5RKYjqoW8Mxgessg4wBtK4FsfdrIUIZoiVTxxI32pns137HQ
aLdwIC57yU94RxVprzAyRX4PXntUhs3hP2mx5zP66WgGOB5MF0KFmtF4ioucuAZhaClx1796tgkv
zctXFiEcRhDeKVCQVXL9KVJgcbz9SNKTNv234bBzexfjSkX15EzirmKVYYODB67NV0kUGjWEl2hV
vMbyokB8T+/Q5emDWlZ+T8Go4nlwWx1lRofWwp8y4GjH3dKb70oLweKP4N5O9U6HLG2eL451RpTy
UWEe7j3ba4Pgv0R+R/Bc4rRIkg5V+McoVkZGl+/LAnwYU35smxCHzb9XYVt31TtmDaFptk++1YhX
rHOPja53rj3JpFLrnMhsZOSz9MolzoFAImonNXgkfRj/hoC1A/g0EXOsIJmxrYBxGBXEsUj3frzw
TnzJNsR1IkzGA+af/IWk6FLXvmNcZuj+ekV6aEBGc7EQwPL5SEF5M2ANuRxAcBCQVbpOxBYZcnub
0Z4XitJfCMeOuBTG+5vEdP+slgGEn1fGM4AzVLf5W6xV/0tNfb1/PMLaMTXluJTqhU2AdOWCzGzI
j/d3eQ6cId3nvQAIaatQqfO1ZfyAXXkM2mo6seOLRRlU4yhIZEkNHYgT9pXPpdO7yRHUXwagLACI
MGXMEykWCiXWwgjucKwCa9RF7u6JSxIoslrqZusNKRG2fEtfjJVpvre1PeCY4xuWeBGB6cr6g0G5
d52KKVZblo9Wg2hZ5V779XdFffuuS2vBpXFQSWCUuKHYSv7b0PxgPhU1jL7f7pooSizoFKuxOpub
qs7zVwSVTUiwlnc4FHIQztbMn88v1v9YjeL54Rq+ZXc4iqzyZsaUIIN4eRleTAlyiiuQX+ueUjx7
s7a5NZL9hQPtyien0D4IoICFwh9jzKqwLEs0YUotw4e19p7KEM0UsHMWsVL6eHFgYAKtA5UYsQzY
75ZNExFHi4zF2VU731sFaWeZyztVkCfhC/FHtDwrO+5lAycCtNJwfOWsY6hX7brgm4hc0wN2QLhX
n0LQu14KoXbPkEhig3l+XRSr2l2dKXF2WjrrdCRBTuRg8TS2Q11+HaQ2oTWRDM4XvDVtsn0VLPU3
s46O9c21dTnwc9vpFkjIiVN2e26Vy5Un09PzwkykjyrxCDxcjmCReJFBE0o0GhcRAjcGr5lgCVu4
MkVYfTKxZcnLQELSz2N/jVMWlIRf1KIVemiCnLCKYRXZDCVOw/rktjNSTt1YMkXHYVTyBY+FUlkG
ED5t3y9O4TxW/aiIj46nPEInG0cX9lWh8DMTLRhOiXING7fHckziUPTTmdyHypRwEIN/O3PweKRo
GhiskxPzkVHVOo3y2RUhQMforpDcqadNi72gY3U2+srjDhRO3AaOMeMdGnqPWQAlwMqGa2V22f7x
p6ec72V+Fh0u7+U1qX68nkvzmlZUCX8lGikjM7gj2EalyH0OisMpC2EFEBSjT4QTZBZdl6DMpurn
WSSxZp6edDi37Nx7GBgZ5W6B3fWjC5MckAri/mgahh1ain4bQxzmSpfWtTlZSO0MCWOuuNdnu7Rl
Cm6TOv7f5y2gz7wxQZzZIwSOxfXIxxGNY7ivBnS800bQ6XgnCzQcUfVa6wBOY/KElQcO14gn6Ffv
oNXFvJF8t3IcvjftTdFvExC6xR6CC01bWdZ8LOH7fG6wCmNMUYT5oqNM5ge/uQyS+g/RkEL7bjMu
Z0TuNbC1FNKMJeRN8M6CyFI4JACSXyBqkK5AeY1pqL3EquqRTorSaFBrqY+OMs9nhI8QaL3UaUnB
bWx0e4S9JFwwFTVg3HdGtgLpHVy/9o8DvFHpnSN5Vz70k2WmirJabU6Atg9AAKPWamww8e2KBdlO
9QC5NcR4PlZE8DxWkoYQBRQa4ebqaxckWExBJ+6MgjveJ2X75ZimRKOZ5UU+/xo/Jjl0vFCbTMVy
PIonxHObGP75be/QzYu2LPcaglcVJd6DdnsFRdcAMnkISHSsjXSpBu32YLza+yeDwn4E2/uZZMfK
cQZvNNtwaF1tRzAw3F0WuU88gR2s4oT9k4fvWHe9SIcCVY4mk8EUck7JPrcnoyXT3Wb3YyMwcWN/
UttwBu7FQyzAlJHDUfeNXQwAiHeHSqR/8PlDVLATTnM08fooH4ppLMreMh5VKpIN5sPjuN3+WWfN
TDFIuI9ihY82ZgDNrPlgmDfgpKzkSDYYfqjxWhOUtMmHUT4Ni31m8pbFDK8+3Gt+8PM4R2npERMJ
lM1mkLF8GWkDocwqEK5J3KV/bycqAmOHt5Cw8s2hyCGTnHuhToLy5XszXwsTx1YsWRROeOO6SNKy
IyBbgG0+CfBuHvJwxYFW87ZcXp5JkzDYafUMhFU12lgKX3Q/iKRHO3njhAeL87B1Qu+xCAfbxTWN
IK/lBJigJfSWil5hxrWwyUvNteDecXhInyOW9ih2Agcnh/cDfrQxXGZF364winG80IRxWxFj4TjF
3YWSwC7BYvDD/c7msfpGBLRX3xpjbNsKGiDBx14WED/KCoj9inWXz4HS3rlmmDeKXLFOzcUwp74m
YBvFwIa1joIxH0DkG9m7s9ui/O5afvD9O79H/qw294jnC/k5q+19PT+KQ4T8iz4QIfhPEX4ZYe2O
dIEeXhpwi4G2GuDlLKq+uX4mdvRw5QQ6Byf4VcLSQQdyBBYBpfZSOViyuOZBoytAIxB5wneVkkZM
VvQse9gSpMPuU4kClIVBxY3JBvB+jkZZySlTJBsBu6n2V9j9kkJwSi6G9Yyx+RuqfF0cBDMhqoCU
QWTAyzcNzSozLP4k6DCdQOVFuV9QS/culhJ77qzhuKYVmMMqHCPfYUz/jpoLueOg9LMFBUlK4gVX
+sE8XhmxeXLyn+qMQUMvwBp7Ep50bBUsoxbS6e8xvHvKbxVIoEqjOtpkj5srXmt6MS26Law8vJoo
4Bx0Op+MVOFNBMNxw2c9GI27lS0noFnX/JAkVSNvv0z+4nRe44S6238Skh6ETEKEZ0kDPaiia92g
cr2zPls9NB76W9QVaJuV0f2rL+JD8hTm0WX8BBatQHU2oUaGKWjgMoDlms19zEhqxnJqzYe8ZtLZ
rwgFLBgBNOVEn36BUfBPQQl8cADHr69rBMPu4IsvgOGqEUDlePVOou+1DPAk5/0lMwCdR8qP2Szu
MSiqNdh1h44mcA0tuWJpTTw5KsRuHyOg+toEN7xabI0ohF5niWpxehdg0HuG4Ft8/9E7UZWvMpcN
IBGLNpgL5Cv2IMPr8eRYq5yw5tBex41OdXyrbfH0MVHN/n/1JeNjmmwlu8zqMwfzlu8mwYTdTbTh
so8db83jwTSPif08aWgAZhbSEyibWm5riQw4N2139yzSGrj7+W1sYRWHKsb1icZYtqJ/yDjHGhHE
ustApjSiy45qpXVM2iG2xkHL8EnUCZzQUBK65wRyRfIuqBIeh2zJjUkkEIG0WL0+K9+njjWz9xqL
UCbzdVS+ugbPUp2Y7O87/hspRIiI8L+aGof6YZbL0sfSMHvPTaI/HrCGGhSW6nxXOxQI7sMsJEIw
Ht0s9q9/beBLNEZDNGtQ4VJxxBcyF0I96oJIGhwtkcQ/qjjOZbRWgPJlMlXFFwvf5mokGSv2fN1h
opsVaNFMzuCC/AVE2jJfOFGE0w1rZTdpAescNGk28IW4gD3g4sw9JlZovgUef2qnjPOYm1Y7btrn
bCcV4s+TZqeYOH0HYEsECiXXzC+oEiIfj5/q95hsmO68xjqszpvR8ObbWXpogIP7SioPfWTCGwbY
Y2TYNCe3YYFIC90CnLTouv+ifPDspI4+Snrxn7YGuGG8kLxdsYYlI/Yu8owDvyceXcYWhGEyg5O7
Hsa3AjwDY3oWA/tpxouPq64pTS/jOhbDFLY1rqur47an97sST8cJVZIo7XGRrnZHtk1+mpjBcM9A
DNWB8IJ3/0jqGUU/h/hlu3weDVmC+r16Zz+MXSOJ7tlz1+JamWXioTeIo3XwEcn723BFEpaCgLZo
Z+r6VLubNXQdGZ1KsmSkXW/Hk+gNYFTYhlKMRT52S2nd1RRwnSObhJzY00cvfCgoXGPAcWWjw2SO
hsDyo5Y0G9RapmPGhWwYxfFsYoeo6VvDUDytUGSJDcAMnDhU3pIEBQrkU3AlENJA/s7snJqta4Mo
G0mPIn9bBlFouIu9bzQU04JE6A8pkOJfjf9w45jVfOUL/GiAnF4xRd9a/Zm5mNJIw+sjQ/CZGzYH
RZ5mCkK0v14vog/Y4fUqF6emKY9L/2mJpR+d5UN9WwcHpeEmkktl0+EqaX9sO0R4AJunXawcBrRn
AT/m5xkh7I1EMqknbgKoOoKmUr3y6PaUKhP8QgD/6W45IZkqVkGJmZHLB1/c9jXbC6A172TL/Sb4
PhTSSKn3jCUryomIuuqEkHVH56yJCBuMOfx88rdXiZGpP5De6xCag0IXBijv3q5a0NVsFU2uirxI
lADiUiQoLTvTOxa3JQzVyOvHHx2tDcloTH/GM3+tC9k/0QewzJM4p+stjai4r17JOhs1SyVYJf+9
ExYiHbOEo8Qf+knI4peBiscTcNXxrcYNfu0GsH0Vslua0rk6n9H+zmWyl6T81LULiLWJDH69UFSh
wOMzcc7uIZqdbUsKCA7V5GOX+egQZpeINgXDlxwVri2ZV6DtIxK0nojmdfXwu0LhDhIZFthTIItn
cwaqplW5XNpApD4jQKrj4fK2pN8zspDRdhSjQix8MNXLqbEPQ7f3ScgFH+SJ9e1bEWm92Y/rlB/8
2uIrTlIQTiLXp5zHO+Apa/gXF7Wf74AhK6XtjfFQeGIyXnMN34Tmm2opcFiuj+HwsGsde5fMSmcg
8047aMTp8T60Suyz4AqiEI/KCMaFwn0XejzWyHp2fNAR1eslQ1yBYsCF5NNINYtlWjc2Dp4xEKEG
J2f+4ImdXte1jf3t4zVjB/cUfhOfXM2SyAsq4vxIu7NgIqMHen055x+olIFUjNoEcfgCR8qVWdA2
/2zlpXLA+6yB/g6jqCeNQFXNXl788IUtqmrvDwI4Uu1DH/9dMquXpGA/plsrpFj8rRFom7ueO1px
Qkck3sSqvPipTc2ejeC6lQBzm9ieLvAEEszkwRePQ6cZzoFBjFJBC/VTE2zwC16Iyto5R+G4AOTN
jO21l+AGvv/lFfdDooVo7T19a7f6Wwn5909g29OEBlr+paGux/uqIFWrwvWTPb2Gxvh6mVPJ/PqK
BJFbQoERs8EY5KatVjqq79jXEM3E2jCKIegbD67vuWmn2G9LaxThSMZInE1uACSJK1eI6pqTgztC
2Kv2s/xL0z6lXG15XCX0vqssZKCf83OGGpmAzq2OfS04vT2NiwEyyR76L0YeJwbqwX42w10EZ9Vl
zyQBY784zRkwemW1mxSM9GSE0fNPXJb/evM8k6yylX5vN9k2GF9phmYlPqxFj1j67GeosRPWPYAP
xL9jqxbIhqc1NYo1sYxpx+g8PudnNZFgv1Xaj4FpkQRd8v1kOo5+J2zEcSuv5a/4CA4o2llDXsdh
7QUCZ7z4lHF6e/kWLTuCHTpuPhdaybzMW9g73ks1+XFpMuvnv6uhv6/fa9mQRajWZ8wNAWirmWq5
izYfDNwVVw9FBXi1hOakAURbP18ITHpohhz5A8+aznXdik7VNMM4tDOvPlgIWLuPtovym7llZE9L
fiokWpdOxp2Dhc/KqLQJ6xyKqLiCHulWorU8tlOkSrKddqYr7DUcLt0p/yxym0jEBDqUH+19UA8H
xB3psnxu3qbuypnGCjydYD1m7l9/ngzMW6tuCWSaKm6OZd8K07xu04yU4D2dxHFLq279HQIb/7Ya
BDi8/7Kh5DzNXHiHmcTeVARz0kDf6PVn7x29qch13KGNghiwnx6N4HHb92LSpYCfV+3dlMTRGpXv
EyyHyGDR3Zx2P+h7EmbEV+yKmCQufuSOzQyXCw670aa//glaIZN1XZ3C/yU8mEU6sWT8OaWuTxnR
//ptdaB1FQFoJWWOblZysWdaulFrfaq9scjqmIVE6O7bZyUULp9lGRsHtRISaqp/v7AAdFYAIYAM
BqZQBzTOdRTndRmqz/6xN41OheKu3hDG+AvXk3rCxIl5+9dy97e2DrGJ/9eLU8dKMiurhuy0TrWy
ZAbZiyiQ3meOf7luDbuy7MqhIe3221l58nioCnOFVpcKbKP0ucZE6K4LO8ZbVJIYlEAhjKuH8Nej
1OeGI+0NTB1F5yi4n8a6v21wP+Y80+5josat6Klq18/xGt/kUhdwVBrjiyFqvVSe15FxWkotA30L
VznZPBao2se43b2mUhIdZVU8d7EilPyvJt5Go1TR+CuefEzqRXD2jt11TTe3YTJZCgZrYFzxfsuj
MO216huxfvUh54FqsoTGzyULOMEl0Sum9ndpgxACSMjdYv34f1q6pgg1P+tigwIwa8kK1mgbzDpA
4vngmc3kQXm97mxcb3vNmFG6Zx2qPde3+vqt781JVwY4OBG+pVMpQZiCX4WV7aMgpdXSk9m5Ov2Y
Kex3oWBNwSMQT+ee+ilWOzrZqrqhZlownNbzNxUK++FWcTu/VDKfiejWcge3Hu7n5RGmKcKPg6qn
dcp0QqInBZmFy8HXpUIEqWRb7hkBKcvEdRTu4b+1bDLttiUbEmcw955OEAZjBBWkKirBpvfMMXTv
06CE6hEnyyERJwhl+cNbBLWq+XrZY3Gln50xCNPbNieI5/eSCb5LoSwaIAnxzXfsVQtauZKuWpcH
YbOhzK1EPaJYixIj93eUE5uPfThmv7hCv7ftNlLf08vl7wYYQtScj+Ji++0Rj4E2KWg5pK0kfZTg
kFr1UfGZlpEJH5bYiLPSJc6j/t2JepXACIZRQDSgNZU5siGHzfQ+t0KpbdkAOoZrE9w6d8iLlpQU
wRVpUSyR9P2trvNBd0gA21WNKXSrcS5K8UqQqFzAMq+OkGCr4vlmQr43fBp/4y7GhNzc/gjJiYL0
p0K2iVWKhA87kteuMXABBQgR+2CKJlXDJjvsnnmxNvApsndxeym/PCT0K2svdTxUqXe3kdzBTqIB
Q2BZAK8SXJd5sOfE2ufNun5zvWBAleamu3E3HX3baYD/s+od1xsiAc60kY523kyxExi1fRob3Ccy
kxRyHDoQsWZehGcVbSplj+oU/nYwIom/0oo8Mo5qigZ0mQbP7FJ4xLtAAMaF6gdbOG5aZq7zR+QA
gE9G6RKqLoKf8CPXdRXAYsa6g02PKptb1JC1JAqO1ct9gbStufAwU9KdfpJY/zrIrGU5dQQWY7ml
Pbwfs0+Ab/brSI42iGQ2Lbel5W0nLXZJsG7lAhQCzyIRWYpray41vZ7JQ1n0qN3PCZ2ai2U9nBeE
QkmfB/BjmbIYo09riBQLacWZDge+gSP7qmq6Vvv6jLYaxKdy9lxyo5aON4EeZ+c36Q5a1qg0goaA
NjJydwmwZxiBHE3X1YoHEXMUo0qPqbcz+oy76cLnvz3ptUeJX6PiJL6Tod349z/sZz4sQkzEpkZz
QLm7F9q84l+6wB+jaiArfsNoNidH+Dt7MltQgvie5I0xz2OhPfdmGRmCyP1mkCcFrPoBGtdtDEl/
C8cuH9/+Thl1sUH3eNWX0Mmcu1L8F2zKf3q+psXcL85PxRWmEYo2S8lq2XgMzaj/9p4vgYQkiMqd
U7aLVYy0+bJ0iz1Fo9nDFPSDKppvF8xZYCvmwA5i3udQsWwfigPm3pUZL8ijPVobKlI67POsyGe1
rOpGggaMJ++gJlQ6lTAxpjxvGRc1X5B0yanQfyXb5Hq+c6NNta46RpgGFj6LDjEWzy1/nx2Lj8LA
7bL349Jyc6lPWgeOhZs3epK6iyNFw1niyCFrp3ujswGuIrnqfS90n83290FsJkF/Bspa4ICc5iPN
43lUDSVH+BjnsqTX4MjyrZ1rNUlDc4MM0v8WZ4OJboMArbYBlgxO0Go27G1AR4Kj/EL0zpceUnPL
fMnSdVEf7mQn01V9Du06Nvv7rOx+qq8zNaqZSsAuInLCi//NJ5WVOwk9iVl/gnNEqofwFYU6IUjF
yskCzgFBWgNXBFsiZORX+0/CV5Z1pZzJXGLiVxTdLcoJPMvoz7+qH6GhiI9svMUH8Vw7aCuDCGdM
B0daxfkthP4O2BE3JpdfyihQmuXCsv6a0zzXmQ4PVwQYIv7hSoYWkuMA/1yqASmufEN7GD+mkpRW
w2D3NXm1pIS2qvCbfcldynZErOt6ixbR9ckbgGqc/NuW4O0OiKgFKhibzyZYNScE4Dfn3M+oSStA
DGaXUWPxrFbJO1/AP72kNJrtzIUti+XDr4NfGc12UWt5mU4Cci6McAqfXEk3Zl6Jk2cdgMWM6DWF
FpOoN1ghyk9A2HS0P5LU54q1Q60AYDYBqZFRSloRjoCIp+XB3cdoGMSk/f6Su516dGgQ8UsnXqN1
01gKxSX488kSRPpz78jklgIjkviE3jhMEwac7PLnoej4t/zZP+lJWv3XyWzt/cMRNk0ZtiQBruI5
q+FYkKJVQVy0BMAM5wKm4PKZiaFJYMme/I/3tEVWBZm6bfKITGuMU4PruzW8VQRgW9V/7PoVTISh
rC1gzoVGYbdawdgT+yOFbJsvDRiwne8gLh7WhUoFliwQvZt1za2PzS4klVf1tYCVq24ZhFAOtuTk
8uDJcV3Y1Xh9UyeS8S4qXa6r6JuJv5nxR1CoAYMzZYFWKRWzZyd3FHzMI2ZrZSHBKUtoKmedvLoq
FHIuAC4RpZ+eEz9RKEtgljugIGp4jF/4e2UaBcTxQhWO2EVaAuhUuL/fB1ywuEZn48djSLNBcFCU
icqnKq2o4NJxi+vS6xxtIA/QMOA5S/dCbSMcI2E7WpPGC5kHli90pH6QKcP2p+4x7Ge6D4XsPynY
uCVCdMcWZx99Z+Df716vYHCwLiMUje1NmWDA+GN1t/tQYBOdsixj8Vo2dX419cj6802Uy3RCvgMV
yll7bjZogMRsMeWxEAi7U4sUrnLvOnPOgMSP7Urm1lk7ijW0CPHUunefA4hjTD801BQHQUYNom9N
hS0QMFx2XcxzMbih9V35WizRvTzs7tKZURRHh3122gwfJ4U8/cFKm8ZYxwj0g+Q8twzVfp6rthzY
Q+DskdSOc1VYSU9E9iustbXFVjCCECL83rdfMGzOquCykdu/cH4o6Kc8r2uuu/52R0MfhH8JZoKi
Nq1JhVtZ5dYOoFqIS2C2OtFad5tkGWs8Mh3G6rliZrrwv144BRcP0jIRKrvynyGnib2IWnrUu/uH
JyidCSEI2ubjShobeVNNPxcJ4ixgAhAiVT4bx40/K7zhfs1lLVhL3/p4yjAlXyjtoovfGdeDmc85
lV3OoI8KJOVsEJjx9eQhydb77mjm/iPzQNq3+AImQIgea4PRphC9DXZ/kZcRzibDVGwe/KtQEvHb
xmkZbjv/tYB04NR5m+w87DgwFCzLWoUdo9ofRx0q0QzA1Y6BgonIWNp5Y7JPvrvDkByeyI2u7dSB
QnQaFFjEudq67tHm2CXd01LbwynZAuusknAdkLAnwoRq0pY8RDpBRqs8Sp1/8zHoBH504QRjgYp3
lweZslIMvJpn206axKyq0ki8Lp44GJZB/rAGb/b6bb9QqHs2/HpxQ7m3ZOdphHFxI5bLcGaCtwZR
lxbfwMaym7dkPZZ4YpW8brCrIoBqBhZDhxKO2x4dc3tJ1DkRlm6rXJlxY9LuK4z5K5d+XvBGhlcN
cQkqPXv4o1Bjf4kBOupOhQRQ4+cXFA6kyM1A9mSPbLBjsg5fVFvA3pIw6QnrJjACF/sIJYMKrjC7
iRSiYl/MNqZZeghDvejxNWYjRxxngMIJE3ypxsZIgnhTdAj9OsxUnhUrk3jhHQfoZunZCdfbljLS
wJhVLgQ9tfpE8fYERbLYxTq4Rgq6RSEmCKGId7x4c+l+DbWMjx7C4ku5k0va11colxDundAFOYcD
7h/jkGv5Mqy9Sf/13BRzThqVB/CEHYdIVd01GZrWwW4fMX2y/MKhoizvBqJtoglgbBNlZvq0oFBV
dPuoL5Sy9c/s17EBXNZKw4+DGzvXcid3zlLXR2mThPxmq6P8vRs1YgRN8r+vaUXrdOpNa1x6N/T+
C4nG6xJ3+LDd1DiiBOX3IiN8TsNp9gbpHnsmawlYfFVm2PsZe8LggabTMQRb6Q6CH0oLWI8Y+VDc
WJndR1+zSyb1rTnkzMVloShg8345RDMlCmRu5ATlyOUPtlCbo/8LCUHttVK2lqYDhEErnN5YMklN
zb4wbbOR863kl6WgFcuVfzCRpkxxbxmO1BUqTKiW23QmNwt42rnC2eVetHhodHgXHVMIa2bVIPmk
DbKgRICLWSP7aTZXS6yjSwLbXXoGYbdGwAkh+SJS6Nv69YHHz9R7HGOVrgCgA4roY2RsqquUTgpi
2j4ah6xL8Yk2lvOpAoMKmiCwdyF+UcQ0bjiVSBkGB43DfzVIkODbCAnYHWEwCNMXyc/aiHXdSJP6
Pp4qprjDpDvNeX7eXzGF02M5lcVeamI4iC5wD87o1no5it7YUb3mFuxX04k/oqsx58+kIrIjlZG8
rbKkvBXg4w7piinOf+/bGL2KXIt6P5IaIFL15jCKNTjM5PzTKDOtiZ/IOdeY+pWpVF1bA/cW+3J2
iOyH+jsdil2Orz1DQB0bvUmnkv+Yra7AoXw+whhtIMT9bVbyl/VvgziNYNalrfRBIHbcb+dUptIo
+Ph8Da3XWvEoAMDSvhRvAvyLhg0YDH/OPYuwWHuWKy6O/BFp2/Ekknctxy21pc0sSNKf7s3RcWPk
4aua6oZQxxFGQDRoj1JYHaruC/MbrTLh6hvRdty3xX75dznDIObJUH6v/lbvLZRH2/tlSoY8m+wU
TfpF9vDr11UwcWG5CBqMnRHYpFn5LYk2ulNT9K26Kg/e9B9HZZt/XobJwOZI/BTf81DldgwU4mAh
s+DEjbWQAolbcHrbbsK/ssaAYcZISGMnAFOd27gx992qaoY2A9c6ShcJo4g+behf9nbIvLeMZ01x
OUeAWvJFHAs+6PUe2uzSykTQIH/9cnzCWow9LlEWvNCu30nntZkHksC6YwLTTo6tLyO6qhUdFqKh
38ebb4GQ11LPKMPEVJR862LL6mD/LyscfirhviJLqlaCw1zVh7sWfrE+uXHc1Tz3dWccLFfOo3zu
FM4Hvl+DF5pd9L8F3ymJ4AKYA9xPjxGc+Os15Y7OGMlqRQKHrbwiCSyCXDf0mxh3VwGJggN6DYCZ
v7xlKEg+UR51hhLk3jm6gTzDECLtX+cDcUdzf9tY+SZzSK0q25LSrFHJpoCbH7jTvJLjV8maiJka
Byv4kfDZ4RXMUvwl9eyXQ1+wX/35Tfmve5uRbaFkyTepBDrP0Hu7WcT5Pou/7qugsqUguBBIILGt
Srs6Dy2PT8BW5U1N7WW6efNglcPP/tWp7HVRe1qFZoZf9jb4YrdGEn6Akue2kc0RtD3nooJ0vPaJ
wg+AmCXf+QBwVXkKTuFYmwIyKfHJh6CbBW7oojiIHkMh1KDdsSIzaS4KHbRVWhrnkd3WJK76wakT
G56+5cv2QRSnljVve58ZfIY6sUWehVV0s8KOQ55dgpoJlMQCR0twvDTcMhmwZqJdAihz5hEBYecM
edyshCu0OzxakTt7foV6ax6/CmEp1XBuJE6LFp6+M0VObt7owTWYSRcGwBd2SED8hrJXnuMX/7oy
7NJAR54j79wDOqjcr8v6kMYrh2rd7BXTFEKvHbXVS+cWIV37ubWcLAtfKxnDNKzMw2DPqwiqLChy
6hY5b9OcrbhZ2OKcfYUyTYXdAZjCppjYrMt5EPo+UINlsa1KgOM0XbZT+nIInPRPewIeYwyqXRhk
F4EUZ1ejbVf/JFnzpxI0k98flxG6nk2HLT8gYnSBhQM9R1Mkc2QUoeG0L1LaY/jDqZ4i7QKGAVAp
JB2zZS3tjUBe86vAf/C4bwLV2miGs0k4LCdk1om5/1vZal+b8dHUpH7eML+ZcpoZDT8BcrxnMKDj
/s8XpGljvtprjPwY6CN4vdjIggbNXNBYx335hXLn5HZ1iesCGdiF4g1xCaQFhUUxQRBEFwxkeGtD
dicHY0eRAgbP2viOIHyRMIOz5aqbjNb9MKn6tUnlUDdbcu3FtxBoRCARAXoklrTFgph/SOt6C24k
LLktyc4JpZiwDeTuhRSfbBwPzj2kKUzjeSsfhzT5iv1IueQAk3Nutbarhp9AGsTItKeZf28cZnIW
IScFUgFA7VhY8MHCw2B8+m/FsXe58y7L5ZCn4vaUjFCjKDA9oeYY0rhGZULB4inXuB2L4yOFxs8q
k3pKsCZqh6TwvCoz/xbFfuP1ZtDVL53vGFUFmJUs0ntgVeiErbDzCo44jmu3Mq1uOEZnPxkxzSMj
ihH2Nfq1CCH+zinlSgeZxgCDph8eHGVdOLrsQEXdQLetzlK51SLp75i9rvsITup59m/7iw4x+42F
WmGjJ/tPd/lExPixCFTSKv+73mbRlw7vVJpjF5fw2L7WviGbYMg20oV9FCSbna5BiopNDQm9xFbg
PkQqQyZo2XFsdYpBAwjc683fi3WVKEC+OTCdrlj8OWG359Y828Ix5ppEc6FizO3TGthEn7JgorBu
XfBUz+YT7crZanTQ1tyEWN0Du0re8OJcVKjAZ2347tBj1YVlITVb4/mtIP1/mLGoP0wnN320PJn9
ndT3X6+/f9tVOzmFCVtffk7jEH60gFGcWN+cBnNDM5PKW2RQbPFNSt2YaOodcimXcrfT8bAcGlXk
Ds+/W8RHLTmhXmtKGFpbVm91eO1wUn56RU9gl4BDpnqVGxRtrKdunTd2Hot1WTjUYsnHucya783z
uEwY8JpNkU/vUflD6Vp0ogoN9Oqvtz/1etwhr8ZqaJG89ytQahmv/Sr0tSPOMbdoluELVoIgrGxn
wNAJNNaOgj74+XS0+/i94PD8gb4uPs3bo9ZZprU1fB0MTX5HSTCYF3PuP4FaY+tibccuX1z1VENt
DYCXe6mI0IE+JIQxB9E9nIep0qfNNQYGSOlccR4j41crdXfuyLY9ooGsseB7KD14c3bBbvGjXhiV
+4DPl3dWA473SWz5/Kx4FeJeXhCnVeOfkPoPSxF/gvp09+YiMd68HBN2sv94Ddw9rR0a8O6P5HXr
HeDXKXRp6LG7qLnkL2cptRyJ8MQAag7c/KTNtGd6YxX392r5MSLeOTkwmMNHeY2FeNu9DScqZaBB
nU0nYCLVzqPaoBOucHnKaDPDYz/Wi8TdsSqiahXhq/nOD105uVOi41qjiA1oFqrPK4svrlcOOJ5Z
z+jH34woc6nsP5d2XdzoVUO9ZZJQkx4tl92bP+xk7hkDIO4hb9Ih20z1PbBuZr7HK2/R2aXq2Tju
p1TY7WcYXXh8itLvXbD30W8ZyHmSIxEz/VH2/uxn/e1xPqAELOQP1O2TVQ6jm7oxKp1MqpOb5a1I
jsMKm2bu+e/H8rH5EzUZtXkb7aHbBzBL2C4dFKBiBqX3b4jpEAhfRa3wCyGJ2qpJEN/r1uJ3i2No
HChBHtRx9rx3mymhRYS4CRLh9kUo3RxGeoNCmh0M8qo20f9HvxOmQ/PCwX/go9FiBqs1KLGHnr0z
UfaHXC0H0V4PA2HCDFfqcqU/azz/5DErDNHKC2zADNQX07G4I0s83u/t/BYHhNci4TegHaQMeob+
tEYYYSgLpC5iELTek1s07lc7xZJuRHwAvfZAPoHrZ8cdD/qTBeLqcEDix9DLyU+4TLdZUzAJnaRK
UVhue7oGNuBccCqHV8SJUdCd8X9VT/9UpIQDo6FHyYnDr1rth2cXzKju5s7wvnpXnEdUdC8O5c1V
k9KX53Epr+P82kLfvqqtqGchIyI0lSenwz6o2GHyToLgIF2rmG0QVFQrHcB3kufyoY+IElqLeqXJ
LOniqkeRViE1sQ0ozGPgJQAv2S7kWb0JlzhtLqpMx7kKXkJ+BjkVUNn/rZZFW0lJ3KTqTi+cytMx
B+GZ8LIErfK5bLQ7yYUGlk2g/AomdvxEqbH2zwVUPzBwhyrBbAIOx2xhz19iCue6eXatAm/oRGjC
+nQuk11FJZMlHWvXdGxBNjBO6GRbLz0/fk/DJj/NKlBQlJx1/FQrExTGQfNsZvKcJr6pdzInxsbX
/QQz9y8W/5vIEgbnimzA4KzW/Vx6RlGwPASWLFiaEr+0s0RLUZHidgrCGNhlsw3xGacW8qypEShN
roZPar0RfvHnDNTB614Nx8LvjhEcq3PlyI0u2ARARFqWug5IRjLtcVtTLaDanrIlzvTmqZBhj9Bn
XD+CFnzU80Wl2Jc0yuuQ6kKc/LPf9eyD5Z3etaPr3q87ny4ZTSXe20CVIocPWo7HJ1EV+rsJTKat
H25VHHyImeVPtrrPHwDKEyHZNGpS8yaVtZd7XUIKMOzxnPrR12Qtv/I8KjkV8Fn47Z3o8NHb9Zdg
++K1aptsobhKUzpQ4IRzu1ceq7wUb44m1ZzIeu+0JoCk1S27/AA34L3b228B2EfygVVtJcc5FaMn
8Bi3qz92CwXlJBGyGUi8s1DMisbNliDpr8FIlG1kIXlxH2YA0BGiQCSmjTT7OPVLR9jycb+Tt38i
Arr2IuwWCDX6hS4Va8GseJpoHTdHBXzOJzXuzvdtr/0pwZ3PozgBw9TToUG9rmkyscmLnKaFpR2V
sdC8GI179/WBI76xrvzWGigZDO0401huD5ENs9DHoAKpw32qJRXz/0pombYkiMSDZHYjnK16rkHB
Msc4lqCeh74abCyBtVtc6C/VT64emz1W7Ns3owP8JpEqoRHR+TjwLS3Y/5bebScBLF8SxtZ7o3d/
6vgrs2TaMBnUFGRMbhKWX9Iqdr37hQ6pMpo6zKjJEPHl0PjH1U2w6H0v/21U3uTXtpeaR0XR8fM/
BgzdjETH2Fc76K5Z/AFw1ilJS6a45o/dRA44IQsSmmR2si8TWqiBhty8LGRKwuvWPZKkb/POL+Fd
yPWs3akxmWxYzF9NEaiir7uk641u8t+cc9W/AWKFpxetbVXOMsLYplDf1/ZjyR0YocKwLZn4VaEQ
d3TL06jcRvbhV8+QASVtWOpRqc6Wl8uJ0iCunVX09P/Fb2+zU7m2XYb3wq6fj6So3ssjucTNQBHf
eMGW/W7pV+x0Y5zZLXat8h50j9pqen1r+CtT2cCYPJngOetZL+rACRmGUB6utia2pU0MgDiOhlKj
qLFzdBuWo0u1YhyHsSdTMTaoSl62tWcwNEvRn8YKmLCM8supW2D0W+sifhKYbLoRIuVzqINQ/GAp
NKxXDystJxRFHU70HONLa1k/I436OTdqzoRClXX4U7/8wfbTTwLp1RmnekUbiiNFZOjyb+DxFe0v
soO7/JwcO/RO8Qql4C9uFWs+X5j1upgQjZvKM8mR/kSGEUR+7KfbRMN+SdUXqblek6y8u/x3d1Ik
HEIX3nn6f7HnenWmD4XcjVm+fe3jR9svTKBXtTbNfJ418lZ2GLPBLsVHptRRn1/QWRePnRrRHV9c
/45dqUU9sPivE/k5vUp1+CYoOstSbXZkxqM5jRcGkG0NBN7xfjsPCHlUF3cMq8ub8RiujFn1yJ1K
X78La0NgKOXOZQmkphXACKaVJZ1M0uI/1c4vtPKpQFuzL1uo2fkXbf5TltaZtpC/bz5l4HqtSTP5
dCb8Gri/lj6nQLc4x/cd5f1QPV/Vfwa8FRhD8MkwYN/8yZf8+55MpOjSbi0Q61IbrC62i7aevas9
tD/D1d8J2mTWGsrnhnL5JQZ5cGaYJbfqU/EfkmP+jUYa6jAbHf65JLOb9cp+TATF3JySjl5e/dF4
KtDP4HARTqct+22Ss37zYcLhjWCCIANxtqVaFw7rcQ7yguGGqeIvvJlmRnja8rlBa80JKuLH+e7F
5iptdWtNGBzN5YD6JXQxeVZqXT43VJ78N4780Sl6GSTAhwNZFsHYN9bf5PHv+wuZ1RHBO1Iq7C4O
RviL3tmPZCraEidGDnmYvLMso1/CY1lC4VcOGRUkVJShG2MddUod83713jtBVdl0WwH8p1xM/gM+
WM+FEjsGZAilb95oeuKbnUR4aFe7LC2G8wnxjVfpDqs6Zf2k1Tr6j4UyMNY4kyVzg902A5GtgxcF
FcefjVax9y1+13xfLHF1KA0fIN2GIe4HP77cOt9govRTReM39+U2FsDREAjywFqMNHCjff5rXu+H
lDKKgiT+jSMg2oOBMXGNzBmsKokagXzI2Tq/u2j4iFitBFRP1cziBVlGw2OsJ0LbE2/szB0gabV/
M6cnZjdSkX86aiJcPK3daHZv6FBZwJggD5a70qQ6eFWFJF5Wu6W33Ub6oJEpEeepwsO0ao4ToWsq
XYwumVFqldZR/rBWiiLtTo7VOh/5QaYx/9VT9PD9l1P0b7PNK0MI18ajPn3zAvXhM5toxb/DYjqA
Ja5arhzMpbzjhVXLHPg/erZ42JRPMwMzX7H9JPGzSpDiuCk4wu6ZZSU32tNyeYuaVk2hzn8CQsiJ
b0vMTW3DsKIJDfWEj7vPT8XYzvhEALRm1ZKV6xZnMZ6ScbNiha34WFAdB6OM6lHLFU7ysy1PpZ4Z
t7dLwAs0l8lkpwKLmQjdnZ2a1bqKCon7QsIqDO/ApDm+RZmWTlfn6FdWGODfRLzzC3q+vqc1rTvi
imGHmlikuLJzaEjhRjS3Ay5B+Gpu4UNGZiVpln04xBhOviCII+AnvoMI3K7CWpMRK4qUlLi7JJmi
kC/f6+oTlXI6rMesu11IIaRaL8rKKgTjgbHHqKsI4Glq4dvEy3MjOKLjbElgCojfIHZeP3zZ3kmH
Dm/UHiW3E3Pg44lpdmzhsiWcvOxY74+DY4+8hJIc343+aMVbKz3HEagobyWu8Ak2Lyc0IOL/w+iX
DV0p69ztBzoREadlfuElcxU8DzK5PyslHHCB52CxsYyBexHXE0I2z8RtzzJLMs07bPGZBinMMtTE
RAntZo5koCiiokDqGktw3bZJJB9hfmHpgPRIeuLM4Ph0zWDesVYJeIqqhToAwJSyfZg9sc2t79cE
kZLPc581fjE2yS+xUb1YuIDr7uRxm9rmZmDdBygIBgnLmjzkF/ckgRJeUGmvBxCl0O4XHIyGhI7/
OsQWX3XEBUUWG8zo3u+EVwYOs5waL4insm34StLapldm4i8JaZrC/FMztRiUdduatPLQ5hLWEPnc
Qp1TMlT6P3m1zixKpjnFWU4kAQjhAo4HZI9gJ9IRWg4lvoHDF56Ijma10281w1l00yI+DBaHBr3O
C7B1RlW3xqKCObC4uH2jqvU8+oDZh5dFELIYgPeRCSx58SdLDIp+H6uU4M0Hcq96lGpjfwxvi27I
EL9T8yClqovP7MAUwCY4Wn+lobLjl9LlKQyh8HyVStH3uHIKcT//9sPHAJQKO8kZs6OrUF0h2jMj
9upODES0565UebTMGNaWqfmV1fh1jyAf7DjKL1QAWXVrfPL+lFVl23TNb07Hqm67napxM3lv7Mv/
mqx/olM+U+a3AoHQc9r39POX821KtRpdp75o5y1mgL0HtOwAs8kRYbt1CTqON4bKMxnQr6VZcEt5
dzdOWqC95XVFpjw/i8uHMnAOee3zaTprZTkeHoAFsSvBaUSy+d0FyKSy/RKWDhbOwCGvrX5Ufyqt
c5MEs6FETo6bhOBFvgVzTJgGTW3RrXWOrXuO4yscL2HNLXi95PvtmG19aRS8TBdYJSj1zWJb+kVN
xvP3qyaLCi40J3RuPlMBAHeb5t7mRVxxuNn7/sYLbiFvvDfktxdn5bi98LdYjs/o0ypXYckFBLxV
bMf22Tjjr+3f1CFU1Br3tpQ0atzIA9ySd1fe7Q7PEm54NCQfmJL5FELiphpL750cqfeTwgMSDcZn
ZY32aaziVJLPy5DpCN0W5Qb5DxhBAd5UmbM1lkP38ebt4EXlJ2KSA7PIwi0dLtB5vFaTqERsfzJz
uBVaoL226ZlvtE9Dte8Fy2Y+OktpQsEFh9XAfL/h7axOBGLtbWAXVcB1UaLGAP1kU+LRIYt+tDfI
YC5aMLbnZFh/nqNwAIbBxW6M5dDLvTQ0Jz22NBnzgWsUoTvLxkccKQEDef2poq4q3sVQcFxPGNoD
qsUqTGQjp12bPtFWy8Nl4ItacXnTjGalW9VrXuR40zPqomGl2UDy6PPIyjYKWVxzicRrBfsD6QkM
DZLjutGNcU2HsqgMU13/ylsDziB6dtFbqWhnWQ8xsSo1vveoN74LqK4iehduAj13rDHy9e41L+EL
JgWOYWVU5XkMHdoNKhr2AJZy3f4LNojsty4SZkvaaFMFmnXMkIF+Z+yPU2zA9PgQnwXAdJbz/Awg
c3nlapGJ40+FMyMvJvtY5Aax4JYB1gewnmXX3m7rlFx1XExrZl3cWQ1kSWDqz6US/YvcqsHZPIwH
ifatQPBaJCG/p6OFHUDYdJ9XdyRDXe5rLuVQcQGcrafwVG8crp0USQJsVuJTu8TVJrTegByzZAWA
wgs9aMeiU9a7SLePQFI+o49gJYvVtOxA+Ai3fjcA5848zdgerHRTVkyAKJYOF1emdcVF+a0bnxP1
HSH/MlfmvhdwuDuUGbvSi47+ou+jvy9yAVdkpm0esRW1Lrj5w25Xk192yqYc774PJDX5lYXJxr3Q
SEs00lROwqPryVvTrG1phCCEzkGsrWpBcqmGy3WQW1/E5e1UkDYVvntQ78TS6Km0WTjg/aOpRSEV
ER0VKiRHMdTXbARwk0FkZToOjhsGK5SX3AyRJg3kDvsRs2MsMZianIy+M+XvbRHfdGxf8C56r+5E
GVqlhvn/bwW0lgDpg8HZzO2NcSd+qFH9tUD3/ce8fIEys3zPKsnjysSJZj5qPEPq0VACIJfO8ao8
nArJcjmg9qSwOa98pO4kiXpea/2BhVArV57nRg+Cn/qKOqx3bM/iaFXqY2tpJpkYkMS5TZdxp7pF
KI2wUKqJyjK/xTDqmJhPnFLs8rW6SFTZKx08C7sixZvbqgk2rUtUuBsHCYM3xwT8Zfirs5kPJrxg
45CIcWdvYllKQfrdd7DOKjdqXgi5D8OkzNtphTvhpqNRBsjMhxUL7Mh8jK6tAnX33pl0KuFZVHzK
eULOZBlfjYb0DG9dvGwCqvPHY5Mjm42Bai+JO/URcOWtrcXn/M8NGPoH07nPP2Wgl+xUcd5lGiFh
bF28aX/MgvYvdHU8dlO4xofSJgeXEben5aQfToqGtIkL7SE/ec6u30ZW3DIxttdTUWrbc/0DfVD/
JICLYHFmJgjoNBjWkgrgqcbZf9kjOaSLaUOTa+HTcVszRzkj59xKccUV5m8l0EZPa4bE+0q5Csm9
omu/HG1AXieqrhIlCThldbzrMpbwDPD5IPlF5TgSf/EvhZuLMrN+lDJxPFPoPCFoq7cZdYw8jy/W
O7OHpdN43VXOg2BM/nMC9W3EgWTtsvhDoapDyOgqqUMqJP+wQCcWSyvX1Zcq5PmcGNWCmPMC+o+F
G8TLZVZAxjE8UrdqWmi3tzb9vdOOqu7VAdDtkgaxKCpxUN0ANKwWp6hFskSoxfZQH7zlXEVDHz0x
TQfUpHSUTjLx+/XnCCpWn9cEt2dsE4GZL0AHt2eA3shzdU8HD0Kt7Sax7BMOEBf9191YotBA+hm5
iUd5j6iiPkGYdQFm78zbi/w2TxNg1d0xYA5GSbHIfI00YSoqBKRzCdZ4z3NEQaPWLcJFsZcltq9T
V9VYC48+HoNr6B3CdiPiwk4Q/n2xuY0UAzP92zOuddvFWk5Psd03N6ihuWwtux/XbpbP+brdD2gZ
UvrouxRrpQkGiOGPWnA28CUzcvTjEf+u1NmVEBh1aglsD+uEDdrsSIIZ+yVFHgwApJI5BJmNZphz
KgTFKA4709ypqaE+Bxgu71ttKjlezOd24WQNEJRaWlWuM7rxp9FXOGXVcwPGEC3YyW/sKRFljr2F
+UXljeSKBj3WVijvuEq04gPzR7+0WR46vOAT+Su6VT3U6Cgr+ozbMy/X2842uRDlZQLbFH98G1PH
d6+jlg6zLMPR1S33ubED02ubhbF5jgC9gnkCrXhKY7KXSdmFJ19RvOXlRHVW3zaJ9PqpzPbpMFze
JTQqH93GQXL6V0ZlCRa+CyfshLrOlZ9Cq7EMMNjB1If0KuxhkiBi8H5+IBVniDWxiL+raoGUoK+7
VSB06Zi7j83v6xO6O2mDMq7HsDRD4kpXEbqK5LHsaDFlJBUGWaf6/cW3ovlcnqtBRem7TWjxq/ZA
ZYLcHUUhF2m52fkYrV/H8N4T4Cm0KW3GcMhaqOA/gpEvhsy+GjybxLONVsGnnGgtuXaV/YJSFhjM
i/YYHsqvEvxEkFQnLXAyt3Onp0brF7dbHqLySZCblSIT/beagPT5h9ZpOQv8qrftRgpbvzofara1
flntONyM9tDAacXV4usZA9bITv6Sm4wXQT0HqSwDy1PrrYCGbwUSub3SANMgIw/zSmI5QVKrgbsW
x97UviEYvJJ4FJDXCo9urg7CJzoFIVI49+BAyftv1Xv+GVZTVbR2zlJ2SZCqBFTkFwDuFy5hqbkl
YAti2VfCUaM2L+wEqmv+T+ef7JqJtRIw88pygYv1gLpGgaQXGumyE4A139k3wXc1gET6Thc33nDH
XVYuoheSImmLSNVXy0//IjlVxLoKgdMtLM8rNCqLq+btovfgxSkJFLTTSkUdGqOHZwsrwlXcqFDh
5PXCPPPcFQsEykOrw9z6t7mxdGGAVeTiNaMiMj3ep5Z7LuUa6Qcr6cZVXH/zeNHe+7aN+OJMHo9R
X21AwlJS6xcqNpJq0ndES/hfx2V9ZG2QswXuUbBaXPxR0eUp+Ruvvmanv71aRj1gQvjYLADzVWuG
SuB94KWWUe6erSu+1MiLqbv8hUUk3PGpSjCtQJz5CfTIeySm0jq7ENbdUDMv5sjcBlhAn53SBQpi
ZCiLBTtqQ96Q7Di1YclBlTFiv0/691nDletQX5QdJQ2TWZVyRlAaqgsy3FB6KCbhfw2/LCok+tUy
VZzFHLxgS64jvcR4szoJvucmVfXM/ijWD0anmOH19VCTR8iCcDwHpxzrTQY1JQbfhOOzyB9T8KQx
5Oa83hQ8wHFgz2dFtfeCWbXsDjBhY/5vawko+S1yelm0HXeNQ+ACNyoV5D64gW4Nr7hcoiQXOXuv
gDR0B+B5egmaSLaEihTH2V8xBqm6tyXAA5vqiI4jb5XuGFCasWCuvVTR5aNgRFQqbQHCU/OWdVRo
66TYiWn9heygPLXhTvyWaw2vYVy17BKM6gLFkPKnXXwNfnNozVRDFr3x251PV+KUgvHBBKzY++uP
R6q6q1tymexf6VPXR4Z81g5SnQjVN+IjE8agZugIQFNyqrDizrJpB1aWeBA1Ir0zg1q79xBGJOh7
0etY9aN0wFlXR0T0t6cT8ebgzOstE+mbPRZf9zI82UkD26Z+roZY47uej9eOBnfDXaQzdKNceMPM
6uTZO9Y+KnSoh7T/Hf4cNFXybqsWZyyGQLvsNOsa/t9Gzf+MWwsrybSJb5e/OgHJPWkcQ1OXjQKx
P8brDT6NyOBn85K4r6nIlqoAqC/avr6jzwZt7z0JBNwfUTjQv/2CDRgAKvVXTe7LxvUX6lAQnpXp
aqkeiFL9pDampzlIcvG2AcagdiW6COtNPb46F7yn1FNfCB4cABYps6lBJb3s1KspcJZlNnNyaMJ2
nyaCUjBrg39BeoM0ECPFZsRZgjEipvb9tFDVXXJHFT5zj6U7aFxmIJPDVvyhBhMExKgwFM81IfVZ
53CyLx0u66Ax1Am8fx1E6H1iBIKCXbS078ZAXIjjK8aQ/NFui7GHTOC5ZXG/EHHIm7asmlp6B3yw
Ssf2GWIBd3yscjvPPDtq1IYSsaS1LnzqqXrArjwlxF4EdOSoCn/0BYU3hV8/SZKXcok6TlTNjO+x
n/cLgH2URbO0pWUPbUkGe3PRAxIki0t3hKW0TFRNv/JYtSkNo5I62p3TYkutsbANJ8T/UqzmweMr
eJ6iSEZSG1FsOunp7Xm0Y24hJ5R7LGbP13QGmfT0YnVY0Yv79a5pauYQQgQIDgFXWxbArsFkGA1O
/KF8qf30M0i5AoVLn/CnrhP8ojux8zy1SLeJid+mJIbnxQbuN+bUq+oF/Bsj6ZDaBwOZ61veUDzx
1tk5nhjTLQeNKWF6DHhISz9uF8rRzCXlr8gvGiUtS84poFLqTG0hecsW3vxjA1KVGoPALzag8uvu
PWOELyhF0Zxbpc5RqZgwyvdACrtz9Fw1yLOmnStiy2i6F9jH2YKZSh4gNSJJt1Wti9lkMIk3js4P
XqXvQecwHqTiYvPqNNf/3CMRQMXJBdSTMtGBVZfMeMWeLDruZWWfMa5JXrr/M8gYHjb/4OLWMG9X
pLPGU9Ige4SOfdWo6Nh3VnA5IeHc1wMYFnfUhZwOgC7P0KqpSmf5YciOJO35DNWB/hFE1EwuK1Iu
YTCHi0gBJDLYk7Azo/XwY709GFz9WDX7R63eHScE3ou1GbVyxt88TbjoQb4/lrj0b1zkPS/SXne3
6vjU5JMObqVInbrhNqBD7laJHbsWqJIa2cqD4qfcKSwERJ+CtCMAU27UWjImnMEO2YOgpGwfqZG6
JBg/dncWU2dT4I/81ge/yOIyuoQGxZ7cpiTX0dHuNvw8/Cimf6KbtvWB4DnZ38uACdRuIYwb/4ZQ
wHjPmCiGY5sPQPkQuNoJm6QkXmjQ+MeOQfu020mxCQcjNyhuE4WoSBpLbmA93x6TQ4zgTXFi3cOR
zzZhNyAaWESAP0oA0PXnShwS/kS4Usp21uiy+n7omptUcDjP0spVdHTngh9NXgAEO0AG93gyiSd2
TkOLkC6iMLCCYfGVsSFqUBYYeZloxM18qAmgEw/uubNBSPRNSNZQEj3BDSgdEX5tYG5A8MpD+wLn
fLYvlFSZUAV/sk0AkxLmqaoXayKJ2jvQi/Vm/Y1KBhnzcNQbB2Zf3qQPQj4P/s2ryacj7ubImERl
TFfzO4wf81kGeY4V8VgFSf0IZOUjtVmMxI80KhPvSF/szZS/7nmT8t5zXs+gc4h/CyRPGiXflNJ9
ZbQP9QN+Wf+VbOl1xb1kWxvDfDkxjqkh9B/OtQi7hcWdWgupU82LCHJzX+sEQRncGCGuDLgIJppc
f9kp3TuM9Fvn4IxPYE1LYvmifnOz/PzpeROLkSoMU8dgLgfSF6fWz1zmnzpki/ScnEFtYqCql8CG
aGJ2wJM7ID3Snw1C1Jn2Mj+yZContlaqfBfPhR7FfQglXKcu0hOqG7nPhqIP4n6eCeIpFqQ6G1pz
kEujhw3lSF+BnM5YieZAvcmo+CzX/YTj+SrDBHmEVWdJM5nACvJTFnOVlfgsxr8pMxsWtGyzbe4N
6VuOTy/SZFHc5gBxf+EePpFVXC27n4TBJFHxjBjkeFqIZW8xADMJWM3g4TzPpGE0KHshIf5gts9w
pZbiYiEvOeysU2TP45PaspkZHSuKRl4LI22kFf9cvNXBxHcL06glaL/m6j8tryHwhQxxPId6UFPQ
FsVKzuvpeN1WRnbSoDFngWyE7ZLSnVWEwCJv5GerCcjVCiJ7gPJ8nG7gwU7ri/Rxrhv+o++aKY80
7W6aV3wrXIu6SxxtGCOOlX56TRYA7+aZPGxOMUsCK4MYXsUqWC8p7OkbGMBbKb18omJUXTgeiyFl
dJ6Iv2sFz+1AbIKeOEybFCu4S+18xmOg53CeH2zWnnDYHlaenctf+M4ohb2cpIg0PRa/G1wmUa06
sbe6Qc1TwD5QJEiIe0VYRKyaUvn2ot9Ypy00lOMoUiA3p9f0S5qBM5Yjd/keNFMuE4BWm3JMA/Xw
lLTCuls54UcUzn2XrVPiYdoOfJHJH92nOJxYqP1t6a0AlLYKdWeBmOJw0u5VoPAaEphc34vIKV5H
cY3vWna8ge2nwYODjZyrBoItpAt8vxfcd4f/lgVjLLyOyvyawseIMr0pq2s2ZvAPJrA4sA53fiMu
Qo1Um3qO6iWfZeOONdVnLyLvSNkUFSieWA1DxkJEZ6uI0KxSHxzUwOQKZXIZzOqC9jlIimqPg1oy
lS3f7WjTm0hEgqLou9xAOX0BFGrcXjQtFgaokp3909f00C/cmZelp+K0FYM+eYeWvb6pseCUS/zO
leddVbEb7AbiHvcZAK3qXQudZo3gHpKjQX2rvA2aVG4OuIYuqHVG4cDTPJ7hLz2L01u6w96nByCE
haRvOLP1caFcsyCDIHxrRswCKXWBP+kbmSm3XfUh4ouKiBvjXA4pOItRvqRZQtz+raf0IN+LgceP
0+j60ml7z0Yo+mN/FjNif8ByentEdEkZhpwcTxJ9qVescyVl6ng7JGyw0TqKgrifx2ZhmcelGxfr
phArwvfdHxYnn56/qMFCbbAWZtFVX5HQ+DQ/lV/JSUP2kFOgOQJ0+e/cGyvvczAzuJx0UVPLB4CY
JxOwFmooi9Y0jNGO4J0KmTI9cG//8lECOcizdFKCnEt5Bwdbp2B3mTiwgfLKQ8FovPSy8xHnDn1K
1+YRo4CwvsJot5uqfZS2nI99CcBFjLz2pMYSL8p1GnfzjdTdOeeiGIebI6Q23szB/S31OORHToxt
eT9KiEGx7x+FEHrHoFV5aYXqdvkzbSYV+XU5D/BvGFanDOC+V9sfVEl53sMaFjuMCOQcH1TaQM5m
dit2k+5wo5vcN/O+382YJt0S4HLYCR/TdApNVv0WXOOZ7Q4vPaFvwb2a+C9TBHQHy2NF0+wkSc6Z
At2Fec3daHqVq2I3TnuMqwlkFqXR65idvubovNKCBrbOwVBcKBS523p4DYky70okpCM6TcR1oioG
rgOGBKVYGY+0ljS2RBxmPKV9QdD2yqYCyOUm6mzP89mR2J+5/1YrcXElyYiPToJXnkAmvB+wgTGo
bagbbs41ZkeFZpyqmC28w8B62TKp7hjgY1n4GBn7yrCXJzV1ftTBAoGJj019ExiO504UEQmote2H
Ey7Z4is58jGMy03A+4EglJTG7MMIHxVVpcEfMebP6gKGqchzAOQsCvxr6YkMHrwH4+PF2PdTxRsV
gWNTz7uwDGSmcx09HKBUNuW+iasULv6kx6vw9j4iC449C/cFj3ptzcuHAcW2VLciaJBMe/AoqpZ8
Hkg2C7jqRSoi/Q8JBGQpQ8XNmdtcl3Cq1Zo3UOomsAhy/lO+skCWkq9IJZe4rRSKhuuEUnobcFw8
0qm0FXKNnOts2cvdZd/9SMl3nMjvvobXiLotWeeadVdLNIgNH3PK/wVcPD7Cdq98g5G3ecl7LCXP
mVktp0mx+7PQuCEp35kI1wQJTmCCXJVxKHJa9xzDj6lFx3qqBDnme5LFD+rzjAPBQTE5gZDOv1eW
jM4sW/pLI4leOfuRe4LuRbktZUBrAZC2AOFRatETH57ITkc1+DobqUESuoCfrZGFqpVVrnHE9aHZ
2B9usghIvpQxwoRNPtx2HVixaLcEaUNuQG28NpQmDYMA5CpsFbGGzSQUv8PYfWW1Y5HPm33QVGdf
rYO9OSbHmlNG+vo8ARRevYpzlOPvii7aWbvdIgbSqquEUvOJR1Ftrl6MujOh//8byRGUuryLT/ie
eDY0dzFEb3XN8ssnkO51a1dJV7TkWrfdLgmLEG56jjDWc/vUr8lgGeK3nELeCaXbk0qCnj2LeZlq
9gYoRwdOzd+Tw+dKbpyZRJetEAIaV5OlM0EjA2jgops/8Jh81zrnyZXVc171HYFl27BWuczGquSi
wZg3zRM9I0HCfm/7FEvAoFvi7b1JbfV1AWh2DlD/V2p9hlUfFK/bkWn54bfK7lOu3WFF7ualB06F
SrJwWtZlKOaL1liSrdMkB4u9u6k3SDj5rslneoEn/D6BxIDAboTareALgvgiRQO/NwnvB47g5wHz
4xMXBJ+0eH4opNki+L3Os8GqdEU7L+e0Oi1OFKoD26/wN8kQ9XATcwm4zHSsqPYQaKesyqPf3A4n
eauM9W/uHUpn65UpTq1/qUsLhX5VoH+86TktzTXn4Vibok81vO4MqVpkoKNlK+efPPNkvnJ4WJxp
wBTcFwCTQ3652PLeXhokl+dJfku52hHqDALFgcrkDdFv+DFqPJP4y3tapVWDaQ7V4FngKDU4dINy
2Cu3H8Ml08uaMxawXktz008TzuDFG7Ba5n16UIj4azArB9LT/BibUs6NLrpyzQNmr+QxHkEOFbPj
89d98d0+nuFrZo5omDitgNJEOxHmcRHJv1r7jQdcgV29JzJ7hh2w70Pzu9CrxafQ03EXGF+eOQdt
15rMUV1VPj/w8Yb42jZCDYkdlG2qtDAMxjnO+Y8pfNZrP2trZO1ahU+jZam+oTZKWj3vGav8//Tt
yBu10VksZ5NoHKxgWCFAh1PRpnUFVOy2x+wEjY9te8j6OLNeRAB59LUDGQnI/8NRrkC5krqnNyV+
P6QlURek5FMtzY8w6PGpzfcfyOwC0atQEZjEEmYcJJkQUTz3hCqcNU0VvMXHCGZAF5u036VJfyBj
qnlCEv60gM/7cnVQDSrGyU9ocq/8pGt9TWX7YFBvjGR5BlnMrUu5s7UNvUVxN1eey6t+lhjtK21z
cpCzJgxiX2vOGmx9K/EDjI6XnimBe77XoRKrVM2MGceuwJ4T3IKZqDXzY88Wmp29kGH3+gJONU81
zI02NgYdWQ5hThlIIUzH4IxGI0+ROGHZ0yFjEaISXNVK/N4FctvzN7+yI9D+xofIoqHvZ01yx7Ym
IEzMPxKC51jke16YCqFpXq2F6Y5GEEndXbtA2HRidxj8Evw4IUge0ogmRbBO/GLE/rKWjOM8IfZX
zegQ4UmlPXd6Ckdjy4MOxpeXT55JV+E8qQgBq9d+ggSyVrdlQ3BNtEtYvxDzZcZicm2nI4o1DPPv
MSqdQDiBbZJJnaVSabJ5NsZEWGfHCik/C0ZiG7TwCHitkRD2ZxtkktVBNAtG1o1ltc974QFRY4dA
5xw8K0xNZGgk9Cxt3K6om6XTWpeLE7MqriwQORwCpCw5eqi8zLp98YWDc4sp8DCoPoIsnunRHGui
/tpX7k0R2VFqeJBYClOJ8SvYEPHLzR2Ev4qGKPGcdWwMamxdcmMz3buoLdTIaxobXEyqXjmMCpgV
JkVOtdaX/sE3WWb9a7tk0G54XNO4zJGNSUhVvwp7Jc1VDvb680silHapsLEb5OuQY5dqH+AT5z0H
ysidf/FLdRnsF1SDkSG+nbc/pKoI4R6nj6HC3McKWHXgHTixeCZ6+FfMWM36TIO5zJsW621jAlFQ
g0bCX0b3lXvG+cEXKCJKzrEk2ed+tIlTY8FhamShZMi/P3Ztq+Qy0aak1F6w32dm3hFGchg0il3W
N4cpPGSAFkpxS4z7akhSTklmbtgHstax+5IBnEZSIKBWqjM7dIgophzW3DMi9B3psslJ6e7dYj6F
4sXpSJoTKb141ciaAlWE5dCeSBx4AugOajVDGo8joH0XlvluaLjQnOhZ9ntmaNlXxFV1HIkKsJpE
E7WARKVS+J6hsgzSHE2fQH7IW1/EIMcBuov2m4ESxellnvrjUEGrZ93rnf2zX0GQs8hf6TQ5uz3l
qnKs4ddD21RIa+ViDBG3hxLePdg7zm+bLMfXS21r/4crQVjZiLXGGTW0vDDdxeDdn9TRXSlOG5cY
OXu8b22nuZM4MtVvcAz2+dUVSMtjxATTUJXlArKeQRYGlRa9wNCRkwo/vt1dw7Th9JnDrt1vItgM
8MqSqAUS2aUy/4Htk9UW0BwgyMMkEsxKmVfcpQclWpuWrercjSMiKtYNNYk0qXryq6H90rEZSIZG
Vv0yXiVAZtXIxwgdWMOn8E76NG5QzzesL6ynyTlXJd/858xliONhywx5CJIXl+SxO10qRObWZ2eq
P/+RHKCSqFjCaGMNPjJBD0EtZarKJoOvKarWxtssHaE8AxTL3tNScVwhAIpaHS11MouMrd8QxQT6
xglCu5mg7sSvH/1Jd8yC3zuw6cbYLXtGy53P/5QDJ/chSWnlh/G0nxNcDik/tUkzUzMZy1meweAw
KX/nzPYHvSrj3mH9f8kz+JnNU5wV2aiYx7JQOSQmeaubBKEPIzbotPdwGkYduJK3WBv8aot0Pk/T
00+khNc3YZ16qoADlc2YpW3hUUBYc+krRgks2y38a0xh8F1gqlanqBv4m+kpLBVB9EVudbvhlIp0
/x7sAjDur57yxrlHG0RVvCvVrA6DQ5mfVQ2GH3e/pjUC6/LuQG0VTsmBMKFDvnsrK8IYgbt671aN
yNc9QYS53ajBuMDuxNqwJaj+CwC9k8v+Cr+015ZX4LbQPG7qv4cE0HIAImiwAnFMchggunkeYs1c
fPnnQ7MwCTreE4s1ZPBSxyhXwo2dBGFyrX8AeNxEIARwzAYqM4LEh0+dcdhXhTzG3lT4Pp+Fn59I
TjrPLDKiPiki//Cldguo5YrYbbLKtjgvfHCRKrluV7hn7j5mUUrJb34Kyv5u3stfx6AorucUU9bu
l4LEnLO/pRfk44ZEiDdY1lb8TRd4h6RL2V/i22smL4Rq7zD6YeaqQQ8pA96I898mehmKhMjdZlf9
Bq3BmXCMxA6SzujoGPKrmUugp/RIbDUIJTbPW9i+jRgMZwIhyFyT66MFIh31y56RGsZr1qpgvNRY
Ystj1i0Y0NLmlehmUDFihzFqbvasTiOg6FCkg59TcfaExbUxIWZv6bie3cI8I3EuNF5pgrcxIwMd
gCGmQMehgyVbqi3q9aUkfUUXMd2fOIbXzlRVcbVjvts3ey0xvqMnwwxh52Xv6ZFjdouQPVSWIiCq
Fdx+1UjigP3HBr7L4NjMiqCnfMpJ6yJ5GinFnz0QgIOOjK44mZWGgOJJTHjRbWcK+3R1RCAR1JXp
sJ2LmEx+jOehi43n2MO9YOREJYwt+lx2P7/juT7lYp6zzMyfN+Hc3RUMuquPJBOaa6FHKwPdM7O0
W7jfnyaEb183HrjrXBNZXkKagVQEGCa/N6BfOn7PkF7kEMBvYGlDiZX+SzcK02oSibOwZAxEX+KF
ihdNSiAn0e1pUwNIlBu+KEmE3A9odhq1pxtq3Egeklqt9elY9hCEoGBa8ZPeANdwBBO8mGorsbuc
3ExxV8ErZVYVwGnnjdN7J1XigPDy9n8FPMLgvT/XXed7WQHxERZRmMHkRO/Tx0udiDX6YTvBT+vO
k5PHL27ANH2Oz51uhcq2EUjhLu2b4ozKHR6/4hQEhcGDsdJwUI+wic6Pw9pKHQPqo5Ml8ebw+o14
lgLZev33jLjXKEjRYDim8ykgokVtLuCouFTiH+rdIRaenRTNz3GCrMy/XVlrU2y+pawk4u0EPqgG
xFl2/AfCyLnj5nwpW9LxzYiZ6QxyC27ebyl+k109Ktp/dfERQRwcP8bzfgeGt57S2Wu5fsxipuUF
TBbN/BRBQilnwQQOjx4732ooT2AdnZA5z54MAUZKynfwOR86jOOdUgRgsqIg7MFZDAF/L/3bwJhF
IfN2nDxZXWY9DJaXsGnyCe+Uxsv+/Z8IhU4zzi93cch4mv3N4ko6oiArkGPLWT0PXHi9Tty7SZ7I
NXQ5YpntdV7LtILULRlDLwVunt+RLNRPU4fOOV8XmRGFjsYTOXBQLO2f0KM6wzN3ac+6Hnu4RzAy
ScU2EJzJ2HIO5kYn2LWKB0YO9w2/NLIM8A9abMfnCHukUxZD1OMiIG2s6oEzOiNurUWJUdKfGbUC
kPd+fGlcL8akEjoA43xxnsBj3JQvkTPxZuJ8fRQjJnw0h2bFY4AbIoiHSNDVNBEfYDYJ1Gu75bEb
rMBjPTg9crqo5rBpSX3Cj4b8d7cydBaEsJ6P03MtdN6Xw6tkix9jB7trRVQ4mhJTUN8GwBMDgiJJ
mFRWKsGFY/Cd+mjLAepKTbitWRsdXftY3NFkUBhdHw83F469B5LiHYKFxsi92BtlGOdqeo6Y8CsR
iO4KRqBM6o0apEyFCxc9xuxWM+9UWq2vV9Prmj5OHjJxG/rvj21/rmSe4HmO7uBwHrA53smcQpU/
JhU+WnuosZ5OzWr5xOq5+CcMHAcS1Dssp96MhHF6NkNACF2+qshbWlWVo+pxZuU8Sng1PT/Fadeu
97hhzFUQ7arHmaAaP1d00/PBcZqrHY4MGhCzEVFnkZCepTrvF5MLyjT8WAXDHWupS46ijGAHIavc
czzf8qyl6gBVSqcTEgneC2iKOfWG4XkbbnQnOv4kVOMkRCjUykyqQ7y7WYjXZOR6c93FLxYQKBHq
2siGDYNrr4S6YRWwrQqfXajrNt2riRbQ3tgADqA7nfUvd4MXBEi8OZPsrXKwKMzouAOrCjNsLZFf
1uUXt60vYFX+/+oSXfxBXSFOEgQJo6dp60yc7FxTR8ZJ/0Hu+Q84YYIAEU2n5gn7BT8k687oqm5I
uVyW+Pmsi9U5PkBJwyPauYa2lW7HRjUv/np4gvDh+/hZeMrElSFzJpdo/zmQoVPiiTv0UgKijlPp
5oSUgft8Fjjirq4rQrAGrs100QjqAaoU6LH3yRS16VC0nzB9tpCHui9vqAhsz4lNOUdOyomldTBS
DTEIKjgyKy/ThYVkZTGnwR+tyNnEgGcw1tumK5JLAPTdRu9BMxly99QPuwQvEnXsrcJg/YkPfXWh
oY+LRL50+Z/G0urJv4AfaXEDKy1E4TYT4mzFvh7z4+bFSFm4LYtfe0kaUXo5Jk4XYMX+JPQCDGbf
W7Ge4jewuDODaUmluPlvQdjaslnaXxai4Hla07GbbbYLaQsDmTqB60l0nz8cqgcwXa7ohbuJVfyw
JQMOoFoOm+xNgcmBWRPvkBVpKBTy+o+GypQfFmdvipgpyNSBSgUk0ipansKWlcJ0JK9VkObvHHTq
52JUzH+j91T/xmNeu6U7JKD320nUuqcnAWWKzEDIvLFHUPvgFXUpNg5VuIt5eKTS2Yz45RFL1jAz
atzCGpEAlTxIdEcf0QSuFZalxhQnoelmiDF1V7GrRvzcKAD23RH0Fadi7EQj3sqsedEdom0Kc+zZ
Y6UJjff67YFpGpL+wHZ3843/dg89OpszQ00d3rB7dKWWI80rLD7RoKqCdRLPWhVsN8EcOyAr5Gud
dteQNBlI+gCok3JzWt4K+PATd7JSNDmT7LqduEer8sfFne6hW/KGonNg+AWQUcp2XJwafUhSCKdT
Z+eLsz9oWodH7wG11caApWv92rQBJxKYCg1LDLh9hvWLdr9EnYog14JIUUpYuoCmOWrJ799JaQjH
nGWoSORPVYdh3i8BT8Jq/qSsl3RvVINy6SRLOD/UsgGRoZn0VQo4D+knSvBjIPVd7vUeectU4bBz
IErOF2U1LbA1fsdpsm9I3PyESv5HdSv6xQOGvqJNB2+Om1tYMzMnwVr3N7FmEqfm+Wx8nN71XkLH
rl+DDW1LtYNDVfkcGJ3yOmrL2Vyf33Re/DhQJmT0FtNij+1L9hx0otWWJfnPPUUwKL8z/+gZ3Eq/
BdPxKnkX81fkK725jg+1/7XiG67Y748q1D0JzreUXMxpFYta4VQ9YxRJWWWiXZzKiG+0BGedjBqH
pvD/Thb5eAls8azpvkVcNvcCwOm7xPjxEcBY6n1uaxwfMqS3n5U3rjXV1OtB7Qus2ka3l1Fu/Q14
AHea6yLuNPIlgHNw8rTsZUxwRNgE3sfZB4oG73TSuj4C6lCirhczEHZYVLNgGblwmE37OB6mlXS0
ZoPtNafMdmIsC2aUL4WXaYTh+OaetcS/seTGSit8T3Lz+xt4eN75FTDeGEC4Acrtf+RzpBYDHnH2
sHnNAQTqlDmdjmN0IDfTz9BLJvU6TgJsf1clYcTEo1Y/gyguFCqQ/+x0+mwBeE1HFQy//v4NJJtj
qK03yf1qNgdRnh//FRTjuQDjji0zjk28WMEGhs6iEYqqXgdVuEIFOjA1/U88/f9LAva0nAm6Z2o3
xfFy8aCbh4FUOcLW1/dVctFz+TxImkmECHfBVvWUARIDtrcf9eFqm+Pz0r3cO/6BBbUrJplhYVOL
h41UoBxGncICFJ3LWn8UZr+9JX2Yu4oXfm7d+I3p6ud+dIjlXWd039dml/t4m5Va/vAMCH41k7pQ
5VZ13YFJ7yDV4BUzfv5B9KxLLDDVyYOGEbeJeJ+OjSbHihJnusAgugZ7mjo4ulkOzvrSM+7m+gIT
3mItK/YdX2xzw4vKJoHn7RlFG0rsWpqX5x4ycplY7TjPwTVgHfkdlgE3xn7DKzDrnGaGoalLpmGc
lPAmkg2l/iyxLOqq8MrvcrVV1I+tm3FVh78WJZQ3IiiRnTB/hUfCERH5SblNeIdGxF+FXXfINYCq
p5dBfwgO8zH+mPhU+lu/PUiKI753A3B4HxZ7vSFeJe+poJBzBHYUc/cod8bknihshEV7bdXpVf6A
565qsKw6DD87hGLdmMRD+UEy7DeBowheZ7/WBFHTkOYoAbAehHzGyXOnRTH+zvDZdblyLxphF1xL
UsSx6IEEHA3q5h+QbU6vp3+zIo1IHbrWFdqWKSnoj2mmcYpXRtpHhmnGYQJKK09KN/Vm+zgmtIa3
YzGybfTYoeVokraW69Z7J9WyjNbZaUUrvDZ414ATYl2ZzF1eNuOhnUsNWZqNt6TxwPxvmqTLiDaz
qmfnlMVjgBNslyXTjPtTyPFdSvEf34A3IQEq/LNkcemk+JEfBmrHfkbvBgh/B/NChYJCTMWxcfA5
09S/61s0oLuQfZzZhYR95M4zvWfRnruRSUuKU5a3YfOrW9ycYJr3aoMlfk9BQs2mBl0wWjPL5wV8
F2zI9G/NBB0qHCx/15hLtCK1fV2R1v39YSeoi5h0dSItMpDso+r6+aUGndsytI8IzBwFRqBiK7cc
5obsjA/v0sWn0qbigLbIToMWccLhD6uqv6Sa12Cjmr0WfsLv7jkuRFzp/+jwI//L3iY/dt944N6A
ytLEj0Vu0lTL8c+Cu4NGfNhHOspRhf5RucB1X/Y2jmfWGpecuPoi6Dd4bQu0CIoYtmdG1ZiQ9Yn2
EW8GiOwq9GpALwcorOs3pRqVyAKI67tgYcWuCuRPO97cstpLO2DDlSUOTI9f1pOEEErfA2zFOL8U
ayXADKDtAj6sua9ybvCqzQot7/ILk0mZ963RaB71kwMOoKL/jLZCvyOY0vOhY707ay8PTeUVMesJ
uE0PLMTYDyxWb5f1lMSPhiunIaSYELwGRnkLkeKnuteSLwhZiCzCX1DAlE0XrJQrLEcJu99FZ3tu
pYQeW9FkvdZ+nCY/8iQ8QAU/gEHFrD6jRPgCNcgW37HKIIz7qQ8ZsQ3t70Ry8jWiKIdHqDcJeU5q
06rWFEVPo1UV19gJs5kzRFHuR89Rft+i0p6RJugNt66UWFA0tnHktel/AaQTIEDNdCixZ+v33PTN
zEMq1bCRMJUm/RienckgjT15ArI5Rm8FA4/8J08sNUhPZrWXnKIAmSCEaski8Wi/LL9Y+4zaCYUF
i5Gz/Gb/3K3Xuh05EJvmYaVebexv2dHqUKWkesHJXOIK30QpO0ff/0+1e/ZvQ2OQsAZpxboEkbm2
IxeBOJvRLU9/2UfNCXQjkvZKYAkunYvnYNS3f+0PY1QdYVW4GpXczkZKsFF/tc2J84ZiiyoOU2zP
p3quMXHwvICTe2ZX9fwFo5s3z59X4M2Q82EuQF1Y6B92bT/4QakmRW8j/920bnml4DI8gy2IsFgu
9HvHcgw6u9u1yyCd/p/MisSUIhK4FeIogOQrN6+EWYTWt5saIbFbOC+4XNUYjDlW7QFNS+EPLWjf
6j29fUS+PbKQhX1PC/Ql+F2hCW8W8v4gfYqfjqsrl6b3g7xblBmgqlW5MtgbXCg9Sp1aKJz7+3jY
g32+aLFwraGP90pajjPllCPSLWen/Vb+uviYU9FVQvQaQwMOp3MQ0RajiPGta5ZhakTxoRzf0EgY
RprUnaiLntpW0SQdPUXI61WP6ELRR9XG/4zufu5zpRryOaa7rC6Dc661K9eqIf/fm36Sof6modO+
Js/gIx4nxRTn5zF6fUmSL8l7vLv/GQiY+x0o7W9lBQ+pMMWEVDrrlzMxd1sZElAoCCOnqBTqg19v
wIjvhyAeJ0A9TjWN2EccldGeEhkSkv17cwbbMuyqqlSBC6vgi1QQ4Xk0SdfTUSNAvutkyVYrWA+P
/U5Wk6qvkZAMoYJuiU+prjJrizF+WFdGL7aX0/0LtkgCckfs62YOBOqtYxg0/iN28T4TWamn4EUP
WmVzqDkCqWoO9uXHyqG4Vv9FxVi0YExvkgKCCOb8JSpfRIDeaE5TVHo03vSmoDdXlkwuI8MPAl2M
qpcsHkWR0GLRMNusBf7ewRslmZGxYQAxd0rRqGNq5PVHXGnydJtHQMhyBqKdIS1QiB6CqhxGMicO
HMTMbrfAryMboORYac2lWsbo71PNGXZZZ4aCUvtkNnPT0C4bPOxwm6JcYkpsiLlFQB2qXNo0qp9k
PthJtewN4uGMuBZZgUGY2B+PXTDACDT06fFWdS2dbS8Mmqp2yKkzzFqQreGWeEgnbeih5dEU8YyB
4DSmgkWEdTeeH7mOhmpepXUI5F9mK6DhAKTPssVMYrWeXH2Oe9yM8RLz+vayly9qsSHD8dW2+MN5
JDyfAW3HfqR2pUBQjdGmi+DN2d0J76V7UMPPEXccABhhw40+dTvobBPPhTqMW1k1n5d/+JwGG3P7
r44pcOcN+7X6WK8cV8dIMSUhsn8ViLSYLG+gDttkY+gn931+TCWwwH7h9iTPKoeoYBLBLXrn+01Y
jJOcOgdCTQWzzZvYGEEgU62bCNxTthuQ5Uut8wsYV4K67cAC1sk6sFfIx0lIhvIilJD6S/QufFHw
mo66blyDCh75m3cIuJ/ynfNMvs5/RW0hNgU23vXTzYR3Qbw1AVxsIcVlO3ym8EheR7a7uFfGwEa9
2ckg3x0i+cx3g7jVpOk1J3QIYKbrx95ayWt5ABz6Vo4oL+J7sZLegKcpyQsBapl0vaiZH4p1Hwio
N6WIF4M5gIKVg544oPUFBaYTnOOSfxpc2Xuw9LsyzloDEKFbyY/Gd8+NJRJq0zvx1APsp3pEm5sc
H0IBVU8LXKgteRfaN1xQjg23h+x53u8X3FmAvkwZljMONuCNPMsi9YR9Or+knUKtTuM5HaRymAZa
bhuwREiJkkRu5mPKbS/7H5vFTDQhkD9Fn45JklqUa/kx+CcH7D1ni+qpmLYHVG2rix+mPqQ576lf
zDUeXrhONzcpZLorAeCks5oGxcnIX+nNV6zhH92vurADuZXAfgRfJ2fDA1HsahgejSYVSKeX3iIC
1hIry3b5CKQHOe5JMJXyh5Gl1tZsBvy7spLPD8Y79WiAkZlx/6T8y42Br7YCc9/ShAopxwSwnlIt
hcdKmCSG8k0gi1T8JRI6VfFKkpln//EtLFX3uDZx9JPtPW2oHephjMa74O+vyK9fD/sV19JlRZhy
7bNBf+8Yhixifl3ndl41k8lbbcIp4vWUA0P5phIrRCSbIxlhvRIAILx1P6xXVuinm6ngb3gTWuZw
4FUSQ7TYtW/TpFPPXhAhFx6dUjgCT/oG90y5beEkluFF1M/EKoHM6LtPxZd7k1Erz8Us0ZsflbYR
dCwZV+2DhIARmf2mtalO8QPswYrBh0qmJ82+G/wAc91h1JIFVaiBlNihx7Nwe/oUeFpAeh7I84yQ
UZYmdEGd4URz/OXX0sxG3eYWiP96KytWgHirxnXUOeew/OXppJNm/t91EQ6QPz7yt2RPe1jsFUSY
BoB2Pzysly4Ch0mLxb+yipk7OFELNdH1GEBWJ+wXpfCfxW6absEoy8Zp1eyf5rqLoq+sF545oegs
9DeqWAyl1M/iUetWEFd2RlCM2xLSpVKByviNlwwsiD/jfTJ/YXGjmz9LqHI+dYnNCX8mU1HanJ+p
K9BIGU1so2dWmM7FGpA4C+Iv6joJka1/YrKGbKcEHrCsq7E1SWSZ5IeIqPMX+91tG4vd8Tiiy0zJ
n5D8bbOKQxbsweCVIzRBZoNMr2rhjqXjkr1pzb+Kkb7Dxub9zFJ7bk5kikKer+0xXk40yh1WKKIz
coVOnzUeS5/WJ/92pB5oWYaEZySFdXiaKJ0at2IdnnjSEKAS7j3WhMIPtBWDETqTfyhPVffv4sS7
rMjFOpAo57iTph+NoxpCO6uyxwqExu7B7wcBCmPq2a5CIQJQK/cu3m1ocJGHbbPd41SGIorNTzTw
a6V3GVdjm+af/4D+Nt0FSesy334GsCcUEqe9cDhMaibO0fG8Hy4q0MX+ALbXBtzWCrUQcDcLw7Uj
jDfUlP4QDNKJmNrERrS4YkydDmwSlwuUyqKgE7e9EFKJdSh3sMXinJpEZHdMMXnqpFxG/ZE2oCdQ
mEq2kiBCTmWSF30vcFTXCkXcIpqOlJ/Heimkym52Dop9q8MAzmdpz4ic8FFjh/A3CwOyY9IN/wfP
30jJnxnNwGgz7+V6Ijsx/hbDm+yx/F6fYINKE40e3BzQbP+HqHEOW8pfeIOsJKumRcvUinqdgxmh
HPfyEVI+wW52Csk7ls+fMr/J+T0baX3YmKO+FTeiqxwVcEzH2RiJ41HrvHl2nTMBy8XVJyONhgLh
AGLkMTjaNHLpbWQBmxCYlsK8BCICvHiZCNPg89F9hIXuMPeuRIAxcjv6kcEcjLhNS6yGnsfjiugJ
ubnhIxlGxTkRUgczOfTXufo2jHfkoeWQs5dTaemjDFseGV4zVVX9YCDsaTPNt6hD2Ei/4qcLsbFS
5bnMfbn8ofFCcNvYVIO0x2XX3dEBcVPqVjN3jwb9FSnzZ+b7Us6l6d1rIu6dosg5FuMPYkBxp27O
6I+desGESK4kD2V1Z7//cxkejmGniO2ZnEya30J7P/SOjxb2PQeKqmQ3SWoI3mqZNlAItMZ9htyL
W6CBeiq+Fp3U1u71njXLz4uJc1LdF5IQ8YEN+4ICjgR/VeSF8243M9Bpsw7F4VCwxjS4UDpxRqYd
AB+kz0+JUlVFj6XKMOB4JOdLwMf71jUM5mxWVXlyjkZ8uwbsuo8EgVncUWl87mNh68zfyo1vUTkh
olGxmw2MF1vK1W1ddNqIKHpcZg5cAU7Ihg3kKzxY18fh5r75w88W0wfVvH7TUGww6KB2Y2hsAwt7
2UDtF5y15sdosP5nbBmLNaVo9dDthfTMU1T67joL+Lq+BO9q5Jeyb0XyOdx+mTip9LFwwgfeSPEr
UaHXUb14QRtrHtc+6KP9EecTaVuj+qcGsmh3++kkwPMRvQY9wU95RfFWbnjtWqfpN4qqLlosCb5J
sD4Tr+GoaIGkjafJiCffuf4iaBhWPEbK1ScZlOtNWk5e7Nc3S5JdJ4bT4Eeld0gn4F7N4ns/MnsH
XGKP2olpPfCJY5AzqBfsHaTUK7QrkDpDRyWy3kt/GDAJj8lgy4Qrbxeh+Mr0Qez0l5mPlGKtJNXf
XJiPl+C2uTB2K/zvtWYG2rV8hXC0/HRJtPTWLyZE6o+1mcvhWZsUtfbtRhZes8iFLBrSDEBw6+oC
TNZ07w29o4kPhiwRUlf7rwHCwkd9oAt+ksaLG2Z5hTCV27AaS15yUUg+1UkFYEKsd2kiNoBqBUqm
AbIG3vXQ0Y35c8RsoMNIMrtGee6jGhBg9rguDbiTi2DHL7AbeUAvbcT27naooXzHX5GgziWFZfq0
wtEheiCRPzzf+cILvMLEbekhy8O0/0BU0+VacRwLa69sA9Lbs18JR7fv+d9H+73rsbiPAZyNqwhM
rFqllIZLHANqcCpBCWmLvY3q/O1VWjswiHLJeX0IwimQAiPWrrMXuinmNWJYhCMv6HxBYp23dhdI
a1cfliW89sYIdb5nncHN7hNaEPTKK7F1NkgawPhQFODnJpxEVWVGfU7nOnVKTQF/MXLykU67tAzb
iF5pX4L5dA/QTowlnIA0VtpfFsmn5uHJV2+Sp8B7B3caVqjyJCGJTII+CV59fJyItu5w1v5SXlS4
knwV/aq5cKzXyCjQ34GIkvekfDt4h4MkbNax6AY1t+TtzPnlpxTA8m0F4ddzMX9Q1qf8eRGqTX8c
PDX1JoOwNBNdLH9ZGzumRL91OSJ1APtVYjTTk7VTm4Y6O0mFes8LcxUXIcgtqcLEbw4MfBHMGsvG
lr3Sg4Pz2HvFyuMOTvbMD/aPgAL2xTJacRNdIKJOIv+DPcJfvUuvue8GVANR58Fad84GVlTVssxv
6QWzn3egy0bm5Xb74BJWl699TZ0XU0Jqq6bHl1ExeQCC96v45bzArg6NKu344q8bUiU4SN6WYIa7
glbWgXLgiqxvL1LlgBS2F87+z2D0F/QIXWls/GpQJoukbX1Og0t9eAkSfHdkEFBGi9yc2Ucd0s/8
aTWICsi7nCx40fQN+Pcp6+7uFcYHaBav2gxkp8mwpu62nhBxo7Zjg+ng7uVs1w9d/+2Yw8xUqxro
XC0eR+vVW4woI9Xr34Ik0/svvl+lhhLdVvP6QfDJWwo6FHIGa6Ar9jIC4eucRzv6Tgzxze+vJ2HK
ouCuS3GWoBwpkhTKOMvqbMFwca2m08Uffx8gbcSgXk5fiwm+vCA3hDORwMEdPq0w37BkfNn43Qhs
eF9TFKKl08j+yrK3tAfvHicLZ6k3pz8aeqCciMW5P2T2A6J6/WtSqvX+Y6rJ+kqN6K3TKSPtbXfy
1oaBxEF1EMlmgc78xel9/jWlYIeOxtCMhpacGZmOpjRsH3IWMZevtzhgsYRtC6Psi7kplq2dp8Yu
GVhjqBeMkIICpHmIpzM4/Sp4h/kjI28undytE5O9Suq9IZ9c1a/5rcHsumiBFA8iB7Axxi1v74rM
rOUBc0Mz91IQZdKUAs7s8iN4xQqyPuBYPWruRkqJJgcwVIFGNaoGGzw4AycsjbSHED0fZUp/BKX1
vtmW1Rw9NYdaUlZRu/LqBE6BO4xcftSzoFqUGEtGx9XOpXAXOl+FRy6FY7UZQT0tZ+bSBwhyCrZL
RaIEMOknogqGfct4SjgM9N74Wr8rStTbmyX3eMX5UAv4W/YZ9J1NKgAfN3EGRQ42el1azUjEGmLk
h8/Tr+XaWxREQ2feY1KyFO1ygkmiEPb371218j7eLd4669XoE2sXXrwFsP64fr9alqKBaPha1VJx
2lPjzXjNYumsxyvFM1ipjtIDnbHKKRM7Tg445JHrNlx0CmNTu+yokK11woOxdbru6k5fT/NCSHc0
fJjBweS6sWLY0X68Wr5Xh7E8jktm2K+Kdt2GF2zaLUsuuM4n+87jzyzNNc0mi2Uzztgw9M57kKJk
9RSpz97tjd11Ags/6empyfQbMLM0cLBJh3+TrwcJK6gY2WGozDx22lU4s4R2nmEFUUcBokxAtPi8
NGwRakLv4TaladVk1rG5jImu7bR4Qokk5xdnLoY2NHy3/wdzMH+gBuLJ10lPVDbG+03okN0DKuON
ONHGw7FcbCggHJAmHo+Vlq4mHaVCpabTaCLfv2g8VPp8pFPGqiQkst2HHPe/LmwKvISPjjnCRfd7
y3Bv58IjjpChR5jShhoYz2+m78MZsrxrMlpobDt6v3sL/wzi/ZMyErblwRlDQhbZcYjFevGVvA1v
m0m38egZGDUP6A1pxmaAJw4v6GFmN8SymvV0Ozl7zsFVrbUmKi/E/UQmTzE0l9oP1Ucmr2nvwWat
d5rA6CMJIDd09sArMUNN6mZDgitZZgtat+T6ZPcw7JqW3V0ITZjJz/3On0EOikOZSq3+KiKAAkTr
DclFIznoDyGNSk/f/6SYaV7r52wvL+nZlY7SXOMrkQgBLsydbQhHT9EzpbHnWyYXTL6MoOgdaTCI
n27r1ZhjcA9Dhgh2laGRPPRLkH79M4WHgnvaa3FWVI7B9Aoymr8/KxK8yCiWj7nh0f6F7FETOeX5
okOVh5V3HtCVWefDsm7lR/f4dJEw6lJjjcXEHTSfDmsI0v8hCjV7dHlVxwIhvFLRgiU4VYVktG97
BjocCTNqHRFJhGDzSO96pZ1jYld6jprDLN84XYSB4AFVIhjFB/sJVP32VWAINF8EZn9mARNiLWIz
vX7l9QGXQWOIFBP8ZfQd3GbiJ6sAzJn0Djt9zLRfEO41ioP2lb4b+GSuMrzw1Y+ovs9shYsNIf9C
T6GHnFU7/0EDx6HtzCPpG3CRtvgmOVsdJ7pUc5GYXNj7Vc1OQaOE78S8s1BUBspRmPf7IMNjdkWG
AKWsHK+bhJyIWN6gXInxalCIqm7cGRMou3+ZjyrccI+0scAlDFMSlMGLSOa9YidQsBVucHOsRYkX
P0vOx8DgMnYK4xuZTfxZLR8nekhl1ee7xaaW4zKnA6thKtjRlfRFmNXFFCqgV52BgpCCPWWXNKVc
fKBSp3makr0wMAd6Dlb/6T8oAXxblq4b8Hg4cgaV0roM2ZR4xAtCJx09Pdnfgv8LpqAIr4Jehimb
XHwbcMjyNwv/VYdCNrLg4E/aGXfQRF/ojX4qi0s6NfE+/7Q30OZTLhGGXCOoP8DfGoGMHQ9DCh9b
LYTtO5oeB2CwD/WR9ViGwe+eYHU4OtpqPWn6/o49LTjwJ5nZpJitrR6PaXKQLDKQrrLE1fmXYJPX
0T2e+axWGC3Yz1ujcHCjzK9Qyn0ND5bt2L5m+Gp2yEsk0/lHf2orgJtAtret3MTUAqNpWskDA0Vc
4W61YhegteRD0fOxR3Mx+9QcpwEWCvU6fDCE1Pvym0JjXKxIMvzak/srx4pHG/kActuEkrkoj4ds
lbfp4HM04MWZ9T3acUmIQ7emO9cqlezh7RoXoOSPkNRhb2h5Vu2XnIxvIlIuBk3hq/6LaRK+gb3d
WegqIXVsyJn14BITBcto0mdEqLx1RNAVDkJj4GFgLj+t6ysBoKIJlXy+gM/9PyXfBSe5dbSdAtIl
fRxW3n7N+px1LTBYMJSGTHgHI/R+mq9OjJjat8ChWJ5P+Jut6ktsW6A+2RQ41nOUWkKp2JNiC/su
OcX05BIKBidK+pUP3bcwdYsykywniLCZjFBneN934REH9JX90D+2QhgAWWdDN8tzGXlsbUyE6YJ+
v6lOo2wI0APTlmDcTtM4unwPToEC/1wMNx8F3yvv4FeneHhWtA8PVFDpAaXHy/xs7u5W/rc3OWAv
IKJGVXUP44wYZIWlmFRM9fY1z8BQj5h5fFmlbKJmJkFoZ4qDDGwKj1uB2ZXXE69TzX2rQG0ok6mc
3zlhdTHthSnMKAyCNr210QatsMAq4U+IiHoC1mYs2hxrAHxU24HTUaqfE2zmICYDnTuSPGdgO4I2
ou9k1vC2cQOup2ENsR4DbXmifdfZFRx4AxtKXj6QA34iLXfbrBZdQYVJ8iOfS1DdK6L8d08o11Nz
GqbDmVgnHPKVtK8Tj46NnbpPXLZJ8HAwLELbjQvwmwD9MLt4c5JKZNdtS34Ap42ibZrSB6eutiZU
20b2B2nTJvSqkrt+yMcqZe0n4BPiN/rZN+ux6YFRDnUz8KvSsM6xM58zyl5cR6cA71q5ueE3EtpO
h7aFRmkpXNHq51p2m5pVL2h1TjaAocNRuQOz+o70mlNIviHrbjJg6RfeeIWbS4H/65oCuQwg0NFM
3iTyfdDIFZk7oIuh/P0cBQEZHVzlGAM4D+ch4ODwZ02XkhZMc4EX5Ve3OwLasjro0TZAtTMiWZNY
hJsqx038fV3wYarbeqqEn2VLBfCHPpTHjs3zqBSHjLjWB1q9IgC9UwJ2Ar6/iVArt5htPR9jF0u6
qBQlwNrCOIMqne9+bBkckpGiZyzdWzmlX/bu45fU4Em20BFgC2SUmtp4ooFnUM9HcaNIFeqxHeUp
FZFIsxVJurn6pBuTyQl1rz1d80Wmy+Tx1Y9kV5+GbHBnLw7i23gvjDG+I4IbE0UAHb1w/wprWmt9
lXF8WdzqYfn8yAlvCUQcmwoXGfgr1zTO2/UF9uOGNdqOPD+KvXpP9uN5FpPiqf/mxs+VJQrmEEgQ
7y6RAVPDHtk0MA9xx2RlD0hwyEUHj0o+ibeMUbSjkJUKSAo+7IQ77XsY8lGhjt2oI+CHzwX6/dJU
xnVqoItWCZmMdtULf+GG6rLES06W3qKotpk17l+/hg5V4yt1fv511CgK0Nk/vn2u7wXHI7giz5Am
e7equTcsEhNxX3ueaiufrzFmf2biDdprcV/uYBLCVnSQivxmAWIjd21J8dBOr4eTPzUnGyagllQT
RHGMHb7/OLc+kTsARuxizCN4Qafh4k2KKA0fjsmXiYe8yRVJg0dcCXAyeyh6N7U1XhEe5sCd00uM
DSU4YK3IesBa4OSvGMn0tGZaFOGaUR7w4g2Z+r432gJhSrsLpIYpZE0TZW08NeKl/+aMSPwTvcY5
fHD+8DGskdfT1+acr7Mg3BkYBKVBR+pAvndLQ52kct1LFTbZbiucOpw6r8zmpOIOEiwhsFB3PNGE
JG36w4pg0ibVY1mTVrBd+fm5t4WWha5gSd9jFLjagKVwTJOGap+uAnh5jbnaq/itIXQBdeWw5k7Y
2+3BhvgWTeG8OhZiu/CxlriaSazoJl2A7CrN3G5zIlbPDKYBIVdWajmj8WuhoN/kfEWBUr27XDK/
5uitRsX53R2ueOnhIzbugPPx95Ogeqsu3jMmgKpjBkH6x0bJWXJzk6eA0efo97GS3J2KXHe4j/UM
iZT1sq5Ve0WHKZ1PJdpz3+WeIeYQ9v0nK7SrbQITrsHtgdJkqAMntZhAGWtyYPo09yKlEATbT5PE
WVm4TGQzKVD4KcFqDiJIuqrgLog8I1XNejiJD4YIOZkgEp8d0cKsCc/kHHx1qW1yfHORiN2o1SM9
G1T1dl58NbZIy99DujD00hjNt3WWq1xodpiAz6NXezKh54tPRAJfOPHD49R0YG8xBt5zOjp3UD55
cSMET+77tQsPcZxwWVdG15jsDXcjYV17e1tbzaLGYrlGYLL+hr9MW+aix1O1ntXjeJx5TtwNJ5Bv
p9v4+m4ejOf56ueV5uwdxIH69pQ1jyDo8oKzSbMuL71VZ5RWmuh7OlmhlLs/dLF4swOFSPzDOBZR
3IU6anmTppcM2rFfNy3SU5a5StpEhchYOzs2ppQiFm8PQmmYbxZ5y/cKSow4L4qziRB4nCTcObLP
yCk7h4BnnkhAKJfgKHwr4nWb91j86Nwzn+gF3Zjy1mE/V5JG/AkOvVwPNQrk3qle3E7upwvVQ0ZC
Xu1R6R0ToJrMOpcgiUg/ob8ISESnyGBheENfH76mjpSwAuZ4XuviEOwMTDa6WZR3RkI1jXYLDquK
wR8HTgXFHcNlE7PppP1+q2fQt7TEYx2d0SdTndj0Fn7/9bnHFjEvYakt9O8u/1/Wa8p+6QRgX0C+
/kP49ed2cZ0P7G2TU8LCbp8cclPsgMkZWgjOxb/tNbqaAlxHDbLiQ4hFawiVWPA8S95dgyymW+JJ
8A7Zq2upFE4olfFjgyQT6lb2A2bYZHo81tzMgpE89/s2/GngyAiXrhf7z2xYJIyqgTV897Ovn6Nt
xRVaSb/haN035rWUba8t0vcseQmVR4+C9p7Qioc41USlqlClS+v8NTUxvExpoiaffKtCkcZjZ/bt
eAWAFb2XklR4docIIUyoWm/dRiGJ+ObU5VWsPL3sbmWbPjo8bRay5ht9eHEmEVjrxFZRD1AWj1z8
DV07Ezz3jkjgoit6GP7lvMKK4ObYsMFj1FdAjql+WOt3/9Gj0pjf3BOaFyMOj2LQQCryPFtzUZ6L
Rzg8zyhFrMJF5PXmNCxszyBnpY+gu3xbANvj6DabZ1Iz9GaCwMmM3zrsQTG3pqAbMLlP0e7Pbpqr
wvEVKx7TLlaO8hDKazPaRRs6VGlcdGMR2E9hyoqdu7RGVYye+Q9BkCPmrtYyJnG52IoF8PzFrn9S
NDjEbbc8h1vBHS6qrXrsBgtsG2OAcNeUqlmzyzWjp2vKZ3gDzDGbNNX+h1PaxQAgKVt3QPiJuSLh
Budlos9kcGMOuj9yMJGi2yJth9rNtcEyxPFextj0f+dp4h9YrCGvswWmpBoOfQXmaiT2r+yzQfdu
E36T9t5vl4dJU372wttczYtpI2LEPaCcSttNyGCktoY3zdDP3IzGsp4E/T1vWRyr07Zj5H5+RsPz
LafPZ8UqSCtEju84D8hQUuqNS/QMGmKUctm8UhwFL628Y9CbzvgKjPB9CTIUBgvkcyJSMu0ohc+i
qttv6+oUPdJ/+46PmsW/1YL+a6jazW1JzcBo6cYdKsMKvVtOGzDbfAxl3OIDhTkUvnZgrqS6UzOV
lqXRC3d8gemhFw63vLs4QlVvmsiaQMKcd+93kr44yjDx4PQmXfFIj+IZ+hE2DvIfIHREodjvs/Vi
pY4tOBPV5vvrR4ZaG3S6iV126uooHIpOwksgLNNhd7L9xBB2XnGW/EsHkWqW9jxu92JsR2peyrW8
Hck/Nc9k85zgJM8lcq53IYALgxShzvrU3tiGJp7rOCYNLGWA6XRsTulrPKLXJSS3CFhcASE+LKA7
lQQCWRrbW9yEW6VCtg4a5oinchtcuf9WNLB4Uu6Rbu6lR6s7n+ZoIf5XPZiJcz/rAXIlqQ5Gd9tn
ZmTK4XRbvzU+tjacLLO250U8RnQeEoVLO7ELKOKTrJhj0XsA6KAEapYFIN9R5msdmwTLj9JU4frZ
yYQQgzHzzZTE2dyzyH+CCVuhUKGa3xY1U+8zr9QzUbmsrr8Q2TXft9Q4QZxoKfH5oC9Wpgd1M6sj
JxUf3FD7nhcJXTYO139DMgcdYxNAmfpxEG/59n2F4Tys9B3usaLcl82e84rts2TE9wxVZzqRkjTk
Tfnt4FIOvV6V4hhSgFzCO1pph6D73EQgvKVWqH1daFQy9cvzQ3SdbDHHONV356wObSEifoYdks/u
NPz+tTlyT6sToieOOwGeAtNiOpYU6Vc+AjjUIBmUP3zKB5Yqrv+/nyg2l/D21J0C53TTjWAcWojY
2ip0xbqibvaOHxBqPJ+6Upuo6FOjkjgxVxS75fcoeP3KkuKiiYuT3ajdriUtkwyy1t2C/TDgz5ho
PalKFv5Mfs3HrnBGwBKe++Z1BUtXWxzsC01A9bvrs2eTu/9VT//VMjMEwshkUy503WqZ8HNIC0yL
R9KiYuWH9b5Z3pRZ+5wdFJJvWx3+d+LKcsuu5Qz7j0VyC35qxbpkF28vFqbvj4uFNINGASiMpP/N
Lah+ITsm08/kpeeRTCMNLeHyLpFJrzfU94iUXQrH0BVQZf7b8vtb3L0xOOc5TJfyKoF9fQaWU7PV
IlEZgfXNDH0u1SgpoaVROaQU/2d2A5THob3kothOMHW8MwfbbErUV88eiSbeZjMG7nrzype2/s0H
+7+1Yp2mTIfMoOKQh1rTMeiOBFJ4vCOdFcuuwPXfPLjHm4uFry4pRlSIdp8owPG0QRS1Ctc//y1n
7GL9JzWqLw+ocT3T3AyS4DbqQAel5/dn5iUDgNln0nB5OwjudwHcuDqdSUoIqKqgP5GDK+FEtku6
Tfw79ufcKvHF31Q9zsJKgB5wCBr730dfkIwsDeTMMVdjB17zDIr8Fo4Wk7n/RQyHbbmGlHsSeYoF
8eDKr4ZEHQhLnt6jiRrK7tqRLZxidAn+0HR5WLterXuItOldhUUrLqrMixWoOdutiba191BsZntx
SQljlxgabXLk+N75PiNHoPFWkuzzxuHFk8YMljaC66PKW2WPF5SUIBEFiVTbSzdVMHgJTqqTsGfj
kbW3zvchussuMLQ9ej8SaB5OoqH9wxn1Lz9s58YwtdEgERoPv0GVT+/SO/B+lvWj0G1qE82QjvPv
d1+ThqaL6dPUpJSWn4eZgIhwlr+gz2X1GoJ+r2N1exiVYZ4SxiIUNapa8ylTCOy6fnE+Zhn0J6VG
hgn3XOfOXOlwsqa7j5zwIcue2CSqwvsY/gsBvLSemWudVU/Q4qQNIZX1XDf8FfUfdvcq4l1gWu3u
JUV4QzCAvrOt4whfw4WasKiq+xk7fWkhNODHxmlq+IhP4pGJQIe1gr6CD7AxJ5Sk/33yqEnmU6pd
SnhRt4z4hYfbsaoN2cTLlFkZAYMdjBCUuOtg5duYB6arhVrRsv0fe2OB7SSQIY4iz80z6wMybn54
IV3qypVDaXkwWlg++pmWZGr3BR3KolXMwSYKI1k2n8MZ0dwyOXZe066jaa9WfeZB4BGFMkUF2u6S
XGxY9lJgLt2o8HuH9wzymIKsAzXH8oAStKEWucZ8lYdDadesFgsujn162yTrOBybzyeqt0mATh+g
4Vup3+U3CuxTGC2KMgrggf+FkOcUyKYb193lpuni94bnQS99KhjudkQvTBDNR0aVeTwp35Zlo1kj
EKg0PEh3tM7aylYb1vvCOQiLHzHFRpDmtbYNFGI2aBaEQ4vMko2s6XwcFhPi/Tc+aATVVbtuC/rV
dSQUuwLGC8+pEL3yNyf4TNq+pk7eIu07uMCbfBEC9zXSPp3SMkBU3zz3ghjq/5q4Z3O8mwiCCD5m
XBdVRp/XBxYPdNkREnP1nhWgJ/gkz/5qhNpZODSFqvHnWOpUfdJHv/FtO+iHdeKHzEMFJNB7NKEj
2TvSD63yH3ilph/Dv1JPXOv8d/GCTFUtFzv6d5zIC3K/VQW8IuKQsdNDFxk755gdn0lHtpqQVMN+
R1C4yA2EL8hXmK9ZQ0RzbxlsvKFhK/hhTyXzmzwp1au9PdlL/AIH7Ugw0GBNczVwWtoLDhCM3szD
Z6JX03RJumUEHj1kx1q9ZKlU/ZQMaNUeYvOjrgJ+bKOppq2c+vz58NwwmLKhXjmrgjodEt+JcZ5b
vYk0mx3IzYYqUXeKhcS792nUQzrW+rDYhHAHjM1jrQt1QTf07WtisY+GSLQzng4Tr7nREC5UUN6V
02CP5n+g01CxdnREyyGjBzD4sFwFXrWaXJmJhcthH7EJt2/qi0BIsQkEFL0e+rp82mFC/LXmnY1+
kWIMbVPAofvi++TbIN07IFrmNwC6hks3yidwJaQqulo7VH1weF4WPrRmsAKADGKZUnA52QkWJOhB
VR7uzSVvcLR816F7I17E9nC6PVX7R/LjbrK0dXgVhlV29tTA0PxysN4mm+p9GdVhsnggbxHQD6AY
6NrgKy9fj7mA14pjwK0Sf7KWmO2hG4cO3VdBAyZJctLleuRCHycNIKHO5R1liAER5XLb/8izzj4q
awQTSeVUCywUkXIkw+LIBRmSOAYFHB+tep5Z8HgBVV1ZM2NuURlrI4sJLfgEsXuGTXDgHqXi9qln
20ruqrN4PT+OjkAf5swvZEe/gsJBIFcgqs+lEYqdjdE0JSBT5UM1GPaBrzxHyLxVW0rj22NErNCg
a6ORQnsx4J48NaJ094e9kN/nfGPxkNpfUHLp5FGDe3/JCCBY6r0MNif9Y+F043vLAkcql9A9Dgi3
kkJ5sgy4LIyXTOY2kmYT1pLtw7mi/N4sXUub9kGmIgd/90OR2gqaD5d1os/kED2TrU7pbpD3CZa9
1tN86vToNsqM2hodaM1dMlhiy4SL65xhGNj0UHbGPM5RiwHw9GNQyVcxp3P+l4Y60DJmMRfIE6PQ
O6zZ4g/yM8pCWLOPCVWHQZnnwY/sPQ07kmIObdNw7vtorruX+ndMUJTVmoLy1IgAN+REeqt6aYLt
GuatRXi2JVTgrtijctZ+mKZ27F/UkttxaXlHjNqEDo/i+VZypHtAOTNhxK6K+gWYRr42Wo+yP/uZ
Caa9VuSszEEHYj70MTt0yKl5Do1Y3DQyxBqfcsItpP5iupINr4zwLBfcANnuEEXezNMmFGbakd3U
kgpQSOjgEeroznhsQOHRKCVowxfgTvi4uHE0gSo+FT3NCgAGr+m1CZSCw96CwpERRCXNDU6Ax3L7
g3Wos0S7v7j3ZG7ZsYkdqeYGwZvdeEBuQJQnuN7ZkkreOWQFgsjt1be7nGm4XvfzL4RT+ByYiMXj
4CHK/bGag/5XeHR53A0bN8t9CEeNlQlxOU7EBTtr/woNK2r2hjfH7B24hk92rRFV3E0vAFeYeLdh
zV4llo+shUFtjm2u35r2J65B0SwoRiG0LQDaM3KS6f6qyZSS+erGKgTsEIk9YOtJVU+e8sc0NlIX
FfGkMl5zMTGFnXROLz8h/nytMNClC4//DJto377CvrEGizNoS8ZNYVvZ30bs2gxCjRQ5+krp3qG/
8wycnfcLaAJUoc/ZrLOBYWCLdWuJa4D+OxRhAfktTp1E1+ZAl6P7JjV9jIKrnH2UHS+PvWkgOv0R
f1kHfI5E6tsnI+nxMJq6j56/r+E0uuygTwmQ16cVOfPlIfPbRIX9a6kKdXdUBhBNT2l8UNCUEH8Z
kgtOBxXo7MxzXAAMzLNdIoajC4dQRgxMcvnKmE5U67IIerXBlJXPVHNZcmgtDnx0/DRcMkeJ2Hsj
4og+vCCD0TzEcX+XxKefHp4Lg2GPS9SExYExmAq7ctkAPLFK2+0D3Ny3M0lybgxxEqII5EJqAgvz
bp5LZCQ4YgB8G3QV7z4nyT5vm7GASVJNWmsoRGDMbokaWL68ptaxQASvOsn0EttQMnA/1yR3Dm0Y
BUoTl77x3dTHQyI0072KZKZ4+VtZq9vv0ufvtCyxjuTIqRYLIOmn+GX+MRnrpL2HEsxq3OaLHj5i
d4yy5x7ZkFhIXkrBXVmDoDMyIOwz1LsbgmucH8Xu621HL1V4F7/n1lVHX1PGlWm0uHPFl2edlWn5
neTseXI5ABfl09vSBc94jYMs9nK9erh+5QIVQ4Gf+YZ19F6MIDEE9raC/IbcXSZHY6FEXXKzWeR9
+P8SrNrx60sOvbTW1sZMCH1c8PDZuIbejCcBHQ+P8F3pyd5e9KoFcdupQ2BUKWdLZwShgoUfRPp5
QHaw+XRaA8elvGx4TEqm17jCJO3ppiwgPnUGmJXQlZkgKWv0r53SONnXyXA9i3gFV0Fku5JiIgM5
H2xdZ6UmA9e8LPSgnU1jEwOwzRcpUb/5Edt2nnxquRfrXSKpua7YaIs04xwAGm4P9afQ7flnKcJm
4ktDQmUTCGqEl2cYRpUZdyr/DkdQfQIXxUH1y4VOc0IoD2zuPacuDmIIl6mTtQ8ZXTKsbEPA7rvT
+nTDTbcFj4xmFP9hLJF/6e/CH+GZLuB9L2uPTkwNINeqYKv+seGOIJb5aN+42WPhZvLZVV4PvqY8
/racNHjtphnD0gVllJ/8ocF79Yrf/zo96HPssMnYRykSSBPyDPa9XiTuZ6cWikd3e1/lK7XOGllG
SvWBdLOO6HFvvx50U5f3PfLLceGY4opduGxJhWuHE7oZXWqus9kYkCR+jwqVVHW1XKzQi3Z0EMty
/FUG9mBeeiKGS5Bd2aWPU8xJbSv2JL/qOwNV/9gp3oZbPYqiu/xh8UJnnrTr/yvsACwDVr0UcY4i
EVHtVGYnQj6aerFT6mOiI/rRJIoDRuNB6GU9yYsYgfHlEEV/vOJiGNGicD88TJfzyUofBfYQeegL
g5PBPxcOcBYlU7lqTG5WsFRcd15aNWGlerzYD5x1s23sZ+GIrBfkOYmm3SZmpFxJDRZotJ2U9GtN
iwZXKpI+h/zvecBufOMwpBxwTN0TH5Uc25W+Y1+kgStYpyboajZ2AwSyoG3XgR7siXdHC852evI7
SK5DE0YSsNCRtJd3RWbbLP50rtJIuR5QVxswaGSjQ8xd3GmAl+N0mPG6W18DO1KeCD6V4AgF3XBw
8pS0vOQ1ZAop8Ub6cV9+A+3/fuS/9mzuACH035zpBhUr9tOryDNu90ZSVh1iSIeUZ1BlSYMKFlGf
jW98YhzgHE2yTFIcLQwejbtlP3W8BviZoBhpwzd+vwPIvKyZ/VDUWVaLlQDLS24ZbFAI7R8UxutM
EV+NK+OGyPpvAag+X5TadAWmo87BOFdv3PXPDxe0emzJb/OXaW3OTGginrH6WcYOFnbJB8TbUQN1
n3EPZhecALSWivlYazjceSzUDV3ieWGRRarNFVCTu+Pt34UiJkWr3f3g5/j/tcTVYdV8PODZYETh
0VM3hAoZL1sg2DdEzJ0zLQZ4sPLxIIdhqgMdZ5wuFVDnk147Rmq4/H9AeZTZrKr6tV0BkQBmg7uj
8EsCPp6OKcdhZPL7yMOaIXZ77Sm71Epf53lpOaVVC8IXOYhrEG0ENAc+nR1Nt3X16tLH7rePeFGo
d/UiuoYQ8z1NEmVvxyhqL+JutcQbpBRezwNNtCkMCI4a03ZyMz0mItK6NPGYCAaw3N155A04Wiyl
LFkkv3qxK0zZOqKYC3FNO2QTJLuuqthENfBxby4thmLygmbIo23NgNcJRc8jU3gJoED8eOFRPWjm
pDh0spId2G9jnsCfikJE1FAshCxLabmDEQAoWH90yKZ5+31Y5tktek7kRqODqpeObXj8RLHLkWVS
UNVNahc6v1oC8swlmVklqNUUF1DxzM39CViGnYcrMsFT2J8va/zpFwHCmECuvD6ppIBHngK3eHRA
56x0G/rs21COXl9zBuvz6FhyzvXw+ye0GHDp7s7DUURj6vUy2Fof9t4ylUDYr1GL2nVvPbUh23v1
AkBvn8D0wcWnFcvsttZ4oYtAD4zZGGWwRejlEPLWMxwzWGfoCvzmvVAj2I6w70s+E9AQdxHDdPvf
f4ECbhghDjeeIYGjULltpSktE8uxO8EJz+qp+JhyjYn5ZpS1GxHE1pPuMTp9Rjck7wqAC56deCrz
MSV3eMUIbBLd1OQgvMdRvX6xlBE2lqLMIX9IADw9zGmPManHAVt6xxKnK4mpInula3XhoW+B3/Nx
7IaADDNg3NbTCif5bTTgafzX7eOj36O7WPQluuoXNJtFnxH2CxlWU8zhbFHpAtEM96B0MLiIbxzc
2clfoxkL3VBUmg4tkf3kfbnadWENEzDaidFfxgxlRfj2TQT8dTpZy3MeuUOo39Ufvx9XlFukHgba
TgaWm5RGizWc/1VvLvQnZaxrvzW2AMKXrQUVsRWkYNxk6X/NgIG6QhqZk2yGHuAhWbKOkGyPqJP1
WTMpzJlz8QoJ7hvzxHnumP7TO0527gJq9pvZ3CUx8RtYsVSIhG9NN5Dx9Te5EmQbFNu4bc+FehrJ
XWJD7hWlCXXOYoyBGemdhe4VU1jicmaCq+UXWvS07+WzdZdN2qyNk+E3xrh9vK+mdV/oAp6I7vJx
LwEZ+i68Dkx8lRgEEB5or773BJbbtjOc+gkm/JTfApU5MeTGtmi7z3HxX9JfOQF900jF2Z8GPs9c
A6VSb+krjq+1SzUH6rj9UXNVql9g2VyEOSdtQ3BZKiwdpOhDojyqzc3mcWsrUyZw8nR3Ozu0pBgn
WDbPkwlTOBwDHn0uB082Mo3t9IIz485n0GQg0Ye20XW8dysnnOTgdEsR2MJSQdWX5ZXyDAJNwS3A
lN1lY6C8v6xMtCxVbRBWKMvyadD3woicT/wa2qpRJy7ndBq3ywSRGP5whEOgnnf/ue94Yb/dAO5Y
SrUD/c5ngpH8ai7xt04Bdwi7bQPLCba5EvJPBQIaaXPozwrsIM5v3IzIq87YbQir3M+UoChq2Gy3
fVBAWgOsFeE6rYLYRHBAk0sFfOg8mJzTFJ4Nz0B0T9IIzY8Tc4PqmtrVZB6mmfbu19HgoiktRJHe
lPHVrXwfufQwVRbbNdw2WqQ8CT+5Ij+Tp6/kzguKxEMxFAg/W+i0sX721e0kqjk7RDzLDobel0MQ
9VBEJwuJrQl4CRtc3mxYMcIu7gnIsN1IX2GkYMqriqL9bncWy3ff/mzOpi0EaFH2D/1arzCOuH8e
CpfYenpEAxbTjn2sjLtdTITUxuPVolPxpMcHAWAnCypR27PgOwgHSS+6yz2AyU2SqxPWRqh2bIod
8Q18u3ruw+UMKT8+tPYfwbq5VeUluTV7J5LnY/xw4nodpi4Pbji89AQjZyyJ5qJRKrqpQJTsTeO4
7lx1hXHB/iTE7eWt7MeJcWpaBVsgFeHZJk2oCwYuYWu08btGE2lQupPL7SQkO5srPDoHKLIDrrHG
Hx8oi3S5QsfDArugnqfL+N9hW/SbQtUjhBM9bu/U9T8oaPfhzNiSB8HojwIP1BTgri9/0gWdlXdT
SRklv1KHvE361j3ywE2Pd89KrFCB3k7otpA2OXu04W+XLKAdJ/0FOrVjjkpsdnHyQJAhoFVGB6d+
NXqrcpx98pCv2u+oqSxnkRazZMRqadoxXcQPzB3Q1VtD9UwzIOXGYtgUK9/+mciWpgoD+4X/DnFM
oKABfHEF/JLCMINiY1a3MuTopqItMoUD2hXHAq0pb34/KGz1IBazL5obAKjj4TKpwLScF4gL5QXy
TO+VmH3pVwp0LLY8RpYbGCTc7M6X2m+4Y3o9RygRCOe8LBtFeIdthIzl5AhmQYDuC4RNBspjRtji
dIBnaHEYI02F5/oqdulGv+Sm4z6bGilCdlaZDtv1c+VC1R7qk7IjBZz6lJsNDd2OjhHgKqCHnNdA
u5953DZY0fzsm/YIGeACEV26XQtPSirJ92MbRykzrDf+0x/pL1gaqfhM2Rkx6S619toSAL3EqSBm
5xAt42cdTrbuYywRbQvSU3pXUkv4chLcUzi6eegubn99Qxf/uuYSE3I/n55Hjmtd7Ce3YFGg6LAl
OmXoRxTuoICUCpTOPWBmm5TIfE+02KmoF9ky0R4TaZbeYMs8bpmTsgPEKna0gHFQpQ4LlsSleYnP
RJe7aBHWnCjalslXH5rIMHr66SXmh5rRfz+C+DXDv0hz+r/oT9g42jzLd3NkeY9rhq8Mm6Nj8HTP
Yfy1+1PckbfU6gzjHrDplgyh3IRINkk383IN5kh3CGt+QG8KyR+IKMy5vyHouXltE51C4aZww9ax
fc+lbQI6+4ZZRHaKRQUWZY+pOerxS0z0MpuCXszqpo9ysYy73wBz9sjRW5K4dgXWDFSZTjwZq8ZW
C9FbJONHOY/QsDZAWBZc0EgwRMJI5Pm9+odR6eJU+GH9Z6nH/LzZLyJYbMki42x0VCCt2ah0IGfD
oXBimk2V1RSgCB14pQ65tjnpNmMOB/YO8R5Qdk30JVCg3cFJuaT+7vLaDKJw+fS85R7ZYpQsJvyj
PFqzJs02//ZdJy7nm29VkJkINEiIz3D2JEuq33g5Wx7RuI1E0qPFbsuRVWwtfxsEz+gNoAUHmfRR
897ehjmwgpS/jhqZo5E2apQqpLNLjgD/F1U3ktEISs40hpOpqDMT7FqvUi21PalR9+87lFEhKGpg
I27k0YjJkCrfaf4GAahRQThGhsOYXhGC/oSCEuw/ZInoIiQ+VruIePDELPIr4FAAdurTPh17O8C6
smc95B8qupI1fbH/qXJeQsrRLEOZ8moQ4ob7Kjrbmvk/DkpkP7SHA8/DTHjsdH7y11jieRYolg+0
unRXonvopsHj2zPw8Hm59pYTeUdzfVWO1HdkmcnmSPTfLuimUeAq20THz63VjPfxfxGrt0vWwP4j
ZCT3R594T5uJPAmk3AZFS96Pw1K4lWbft063K79EGTgIkjuv+HYXQS9xwAJDTcy6YPSo2oItVv5G
eXvbolIubpCaUpEEspcobmADIdmslRYBs0Snu9gSGwEPK8QZMQO2PxT7taTN+5ywQpd3WOTpymeX
R1hsh0TZZ74KPPb85u+3PjLnYP3Yqwa5fKXCFqEkx8XRuKXPuk4l3bK60v3LdR9e2nTqKzr1h6D1
o5SzRLWYCR5NXkV/ODaVNwWXfghO1ZrCr7OFOivBcEc5mtP+/2cLfn0t3fne3qKQyNtk38X4p8Zw
SQdKAP7oBNyOWBsTfkJ/7FgN3viz16n4UngpqNTODLameGhhzByfDZ8TpZ2+Dbc2Hd2HmWEWDZjS
A9GPnGy8DwzWapnmLy9XSXfHQ4jL/8UMEdnOf2E2U3DLM5ZU4hZB3U+KgBk+U/KcfwMzwdA0mnnv
dHg13751Gp8ysJCMO4QHXukhh71ZL3e/TALjeL9DKq6lnt9bLwho2KDvU5s3Jupxx75MWRDjqd+Y
nW02ATPi20yIe5zqvDsXi+vluntkVStcxac1vNuiqRuSi57ZukXghkVAPE7hVdQ6QhucUaktIE5O
xg9PbHAOhD94158UINttHj0UTYf3YpwnlFRn2/LIZvaflQT1blKa6mdZEHd789POtGRXOMMZpejQ
uJykcTorWb5J0socgYcDQaxJLzfvcWnQOsc6KmBE3fCdrShS6uFi/7l/eCE2RaKa9sEZVl2OE/M0
erEZrSB0ohoJHqeEM9LqxhvIHYFAWu9KNAj2OOBmTYT9nAvjhqZmYU4KQlruPjkLNBhJuvMOIwat
cnP+E59mLo7BzRI+278eq28SawoFrQQi1xXeLINVrWG1v+SlmTrdOnm3/c8omVN5MJJMbyOhX9YL
oGIPABwO0e4zoXrNsIKKHp/lWXSm4kacy1OkAHzu38+/COppv2m50l44IRRJdtc/RzFWN8qzVDkL
O4f3q3ZsHi0F/VhXseXYYBFVZFa3L17s3/yRxH7uJ+NAFsUpN+x9uybyrwq14nKfXBvj0JzkHI01
wo9uAGtHJ9Mi1bvU77yn02oDeksrPKk6te0pRK9xCpDjHVWxPAgv8/g+ZOm2C1qWqAq5Xbv5BzYM
A2naxr/kBVMmPvGc9JaQ3E9lBoMxfa+NhrpNo2jjWe7kjPIX51AwvmdkxvkOinG8h53DEvB2thwx
dEDTL6RtW000CvpgODn7wK3Q6PxpBQiYloQqR3awIky+tGocTvNjMkqhN3WVSx6Kf5HP10DUb8EQ
zrQulHzK+/fySwys1VlL+tDPNmF/gHcG0f2USqNcmhwM1WXn4YHU15lvoEMLgMLLeU//oYwQzJq7
9EvtDhAfU0CI3wAjBHoDCfCGG0w0YQVl3E0qQztu/fBdjqxKr+Aqc8zyaIi5SLaXQzFmvo4WnoIX
9LEDDHTLuK7JTvdsPABfcdtQkT4PwLu7sKs2vPriT04XdDtxcZ6Ev4UeQSpzqa1Pf5tgmqjy27wg
YSdcP0Ycp4t7W7I+7woCeQI4irjFi5yrSybHbpu5H2YqVJ66iZbPpNjM5I89zQNLX/JQihsqLvRB
9lqHFA3A+eson+YhQeljjH/CiTdxsSn9kotZFj7Xi69pSe48H/uOOu3NoyNEl2kpTYseC2wBuYng
7c9BdRHvj+jcPB8fLR8NGNoXY7I8QeIhBGhPoWQ14/qQAD4qmiEaeCjLhtvNE7nPTm6UZxrfPnLy
qnFR05lSQ3H+ohKc6Shbk2jLMtqcR6MwQVM6pW8KnOfNujQcCwoUCNkqfXiTDa8Mg/TAN5QycKHE
HAfVJ1vhTdb3CIWb8elaIURJbEfam3hdFVX2+nsN5VI1r/vmcbQZUnNcLRri+7p3EaOpioT7oVQL
P4GzHI682w1Q8Q/ekEA+Uors53UbVqJ9HiiDZZs8HFxhccNkihxJkhoKrXqUeKJUSyF43T1O00/z
HvKvV82iYMzjKkOh69/qCg9JJ/fs2hnJIvPM88HneypKsLehCCeqPv5GQ5VToNl7piGOp6WiMRrN
e5s0hRTgLMyMgS9LsEG6JHmlBBS+1iAlVLbYSt/WKDK0B/a0Q1HwqayCTTmQD215j/FuUo8SH0R7
yNrcttR7wezwgPDD1mOPYM0r8Og2Vxyi22MeoivY+66ecvizK2kBsgD+/Iudj1/5GWE/o/csngG5
3vKx2eU3sQ+B6yKcRewojuhhhzaDyZjMAvUTxuhvAoEtkrH95BWIImZFeFg3H+n6VPzL3pjNYUqv
gCIvod3SpLHcO+SNhQdGQhOJVqqtMw/JoDE6gm/GIJtv3BBKR3tihyJH8pd5RIEhoxbKa+ZhnJIJ
NkqitV3j+OhD2v3u7Yvf621076Tx/gR1nLBIyelO/ldnNQuAu8ME9QKuuVJ53YjFLKFJY5ORobZM
u3uu3luWrlUUoLT6YuWyoErqnZVTNN4AfGIpzuie6myaXlhlMS0LCGle/zUBcZsBpm2npp0pDuIu
7h3tcTv0q4mXx7m4FEeNrWqR/CUwdi4tEkSWGnPXHrGfOx4l3lSkwdxVYMqOEdqZblQxd0eWfL3Z
DXbvGbuEhMBC9gjMKE9dVbp6j5Va9bfDNX56oHxwHfxtuQuYBwBdzT7HLaiyJGksGQi+qEvu7LhV
/RbTYZelmfKCZ2NLD8C60NU4xGoDgZbr+Ie6gZnEXi1g0ChRKcN/MmFFkyTDwY4NpvKWK/cz81Vi
YLCEpBrkA94gd9fdRseFqDVSyRlMv1YqWXQENcU5HnGzBl5OJnRPPH1+DBqqgncGJgwrv98CHebN
jmIFn6pAIXCWPFuHHA25hjEvvtAUqiukGxC+ivVI1iyCFDT+ZHNCwrXdvfnjwxVWRIpoIWz6ErAr
2GaAsh4IDwz8fHdXDXAyyL3n1VuREPcdOAKKGpMZg+7XOvUmWySvGQwaG6FmUUbm5x9J99uiN+7c
gqxRCPHiLPlsVB04qvB2+1AKErQUpGBXZT3EXb2h6KX87jIuoMucpxu5s92Q3NwdDWf50VLcXgwC
sCAk7Fr7DkEGoVl3oQeUZmrFUnrFM5P82XfC+8TuGvUVAnzkMuY1G7mhkRlbTIWGgEhN4lD5d6w6
pN43XT/7Aa+P9if6JDSiLstO7lmipmGzT+5oOBPsbzJD2oK92Vz5mGrcx2whL2boGoyA9nEhznWV
8aKd5Z8U6VOACYa6m2z1nCzFJ2dCbxvJvJMmqlAS5L/rJFIX8cDm0ufYmlFUnamzmNDhGffMp0n4
2lDA2rKC+FbUojtzIwheh7DQxv7x2o4GFlqnNe0MxYtk+7WIik4IJquQ1nOFzuCcjWcN1aRAt7EP
G4aVx68O4T8q/keLGvtUZFvCMFzoAoweBatXZSK37PeB6sVFq9CnXSO/Ey4QVkWzo5mWZI7aVdLm
viuiw6YA3vzZ1sAsSHoccbGHmcvp5e5Nk7fLvjBf1WPYa/Npaj6SsA6fsBF24he1WPGiEJGdncvQ
aU2HSBKJ44FGKQ0uCZFh3l+H/aMKPR7BY0BkYz0c56LrE3FOpNv7QYCpiCOoT54wd6/G2L/aI/dB
8OA9yjxg5LvhyfqHCEHFFhNqJSfREmlOPjKL3TYYp51WHjZY+swigi73yfblbnY92TnJuPYjMBxX
aHdH8IpGuQzNibTKZypzcsg39FmeFHnA13Ew0H6n9D9b2EqbhDaeDibs5w1PVlWwcePaJPSeTBhg
eILTIKQ81YX0gMoeV6nuAopOKeQ9KQ5HhBN0ynQ6JY4WJreg+atF5QMIrK244uzhtZqVaFO5/Yzt
Jh08KZ3Lqhr9a2SVLcdSkR9rnAvjApwFIjvuHesP6kr5ASLCJvz/fZrhsTGJ1FwS8nUN2h4yp+ad
jxO/M5hWn/wB+SHuxK7fepukfYsQ+PG87QdQAerWph8mfPz0yNWHkz0AjZJvhEE2EEOxlRNTlU1X
WOEhb7blc9Gxj3KZt+FhmF+hBU7YK0RhynljovFKcpQJe1Be1w4La8LQuYemmO/8yyfJNZtga2Mb
aswWfbaycPB9kNHqOQZ1mzb56R+gRrVG23BsBeoyg0V7Xg0aLCyEP038p05QgR+TxYjBWhFf1TX3
jJ6Kn1vtOLOTeod/z9pHt4raMR7gsw3w8r50CJbYga/dTT4BzrqIso2o5gWCC3J7UazG+R8Bdagg
TIMR27Cr1Aq+WVD5fK4s5THlZICmDS1T5kfQK3JIkpUoAcokCjCeSQO7wJfjnYxTj+RvsWlk8ROr
SDqLnjz6vfm3VGMUPlROaUMGJF9vsoqaQ9MnmuvjHf00vXmFnhccIKkbCAQoWAo9UAvKoOPWwzDF
2RA1fjD5SXnEyaYjAZYEpWrRmWgL2PaEW22mzMUCAil0o9CwOqBKiXFCyumc7nPhb2dUZ0eUa8qm
RbEyXiU+pTea/lKx4B+bczNz+/xJnlIkuPDGn7ZB+MOilP1GCbhJh+JhwyNHxMwcAZcMVLDYYsQa
YCjzbLyaV7IWVBLdVHZjz42TA5pX5l5HHuSC6B2opk+B5bhTJsns0flcZvMoWai5rSxJZrRT/A+J
jaOEBPten4Ibv/CBBBO6Q9rn7UTL2hAjKbK7lH01YTnFIld1WYtk/r4nZrzQga/jNYRgyeOy5yew
sk84VQDpEsjIP3JdNkJKrYkhJINCsq8DsmaQ6Jy8I60hd1JYEB6Qnc+XpuI+H0uTunwOWIX0PF5d
neuorL7rnROU6aEWpg6yXyZu0gnjyu9nwAEDgxosVxindMYHgNDVFIDRqjy5USEPklGFhLVXDh/S
ssWrd0JuBgF0nh6h1xXW+pbzBcKahRSOcIyHs/ZzfjtP5uuA/1Pyoeo00Fg5lFRoApzBKZiwOsl1
dzp0VO+WzZ4xXGkagQqvTHdw7U+27Uo3ndjKZYpsZq2vJlxSdgkbYPXiO2Zsj2ePtphLmmG9X/lz
tUlzu4QPBkJYEHoiu/EnK3c0ADgqFOR9vaWcdzKfTTQBocqNEVG9f9VsslG8dgwsOLlts8bygg+R
13bLneIQd1K+zLHcP8zeD1WSp11wBa943lXmfKM7EOOXDULh93xkVtZT/bPF980ORcfggbeo94jU
Ys7uCHQCl08S96my/+AWVRyhULyBH24sHcX6uNGh4UG/DwMg3mdbY6xY6wDnT3+DIMkX+RCSd65h
Tu0lq+soKsFKDZ9dS3nouL8xK1rXt2bdQ3ancyqcNXIhFT2BT96dPi3xjVmWWLkxFEe5IePaqUaD
KZ3AgdEFGbxeCUJFhU/HmjeujPBVd31JRDXjAhazmvvyVLDwcYSEPOIApKDmta/j3hSgfAUMrpJi
5CNEGEq9nVAB4Wk1Nx50I2H6506ptU/FRaHTLNuR3727mAgycdYYEq8pI9aHGZ28V3lT7yPYuihG
yIhl/FS+kFS26SUnepxkrOEgA+z16fFSgwwkrPUPRoyT8LST4xbhXGYBqScYcZOybXbbuXP/kqsT
OgnawFj3/NAXSNmGThO8hFm7OxkSmRokBWYSLTvi5oXgAksvu/DnrgWAPqjSmnBnWnbA8PfITFHc
z4YPGeF+j9dNdHUFMZL+ZfCsuIYRqcLx9eb7+TAQ1K7nRS+3MD+moh6HvegiLTR2gyj3xy62WCFM
agU3OdtM2SUe4ZIKea/TOx1fwiBY4JbejxOq+h5iTQZlEPd58gc1+0HSROD2sLKkcivAvwmjKJ5Y
7Tbk8a+wIXqywi30vv6QNxX4dfcyeBJ8LfFBRsv8c4K0QLo5DuV6Ajk/e5JroBPGeMZy5qpuLbkR
x9DtyE+JJ1YbgNO0/DHVtwCXRCYJUJq3PcUvD/KX7t55WvlCB/XEkNFFCGUud/sPgjuggXXESh1G
Hm4yxYVJHTrOrJv4yLn8z1JL7SIhwErYRWgQPsQJBW5Mxt+1oDJIOnTQYN3cuXD+iAN0VWqKLq8I
xq/d+F6YX4Q0u2vOy+GU+Xq5SwkpG/EhSaL4IIFVKJlaPte6WzBD3cQToCtxLi1llZwVTDViwaOQ
kv9OPnLYI6LKlpbviG3RkumUZLtkjSKJ5Cb9By/Uu6DiebfTJTUe8hQ50nNG0KTTYOM/NEO5qTM0
p1cw33ckmTKjhnIsgZKLhhVBXabNyDtJ9VOp00ZxTyiXdmD7i7wXhqM43MO0uTFvusFWTDfOZ58N
nupXQ5TQGin6DYGR/DZ3cf1lzph8O5BK75EB5ff6Vu+paCZZ69FjatnLVeNqLWYiZEDrp4hQj4pu
mBrD01dXt7xPWXeYVCnHK6atKVHExu1PDjmO2v76gPOZLmKJsSF1kcBjNYRwjGZ0ArHwWila0ZDd
mEpHIpyGgI23R2mIPLBha5IfEpOwcKGUhYWp7MBES2Q8Rzr40hT6+36QVy5B7FA5fN4tuIjASCNX
785GNkBeNGnQF1OaGOnVYaw5XSM0DgRsMHVxKH6lFz0DisqFpf+ub6BJ4STYCbjNupTmLvGg9yRA
2fEbLurfFuT7VT3/Yn6ZgcNigdiAkNAo46Ltziapw7AJ4HJOJ/iO4JbtGS5ZGjILfQ3k21213dg0
ZiiVcihOjV/J9wsOBOVSFopyclH1RmF2FfNj7JWt47OvwPq8fNSOTd6GVzSorvdzJmXPpCnSkG69
HH6vNGnH8BpeDQElPMKoglJRw6KrXBiLVrJxRRBaMJq9yaiCn86QV2Um+gezAfIigdY20cKmHX95
DqCvhJ0SXQ3oruUO4LsKWJIGuxbKHrl05ihMCh1ABl0BbqsUi0ZUsJqDWSiLKrxt12Htn8mS2g+N
AbinxJAUhiTmML3f+GvGMALjM5WxYmiy212VH4+Y7nQyeh1uRwFQi2OopNYJ51Kf44TNsORzOTWe
w/R1SzrS1Bb3y2n6fVEGifDR5Kw5CBHSJnjI7qNV4Ut7ICWesNc71AChnKKXUkmBT3LXUhOsIonI
o3H0ixKnKxxpYrNUkb+m72o1eXeoG06IfX/ttUsmqz98UTIWyxUnUQ1AO2cyY84KgYldLfH76vy4
1LxtMkpWeHq2Pu+D47/rkn0Ot9eo7NyN1TmnED93n2YC848VqoB5F+ppIFA75yWq4T4VTDCDmsx0
/g2cM+Y69arWEsxSlOe8z4lks4S0IvvayqZkM8spsHZGb9wu68AmcXl/ESojxsQu2jRjj50uyNGS
8xHjl/MhRrMOcTtA92zaNH0B4y4MN0b6w93QSindb2kTsfsAPFB7LiSpT+iqdYYg7ZSNO2xcGtGc
OZxGHASr7SRfMHY8w7aXHsfG2ZyrVtagGUZdywhKBDtuRUT6yDTSJMGaPSqc8RViVt6jLBtUG7zl
nhYVdZfmOYGJuSqVInZIftGKXIY33HLx3rMKSldn7+RWd8xBpWsoyZThZuz76auVMLROQYmvc2EH
MzC5SpQ84RLfYlMBvNO5ggxazobItGryUvbrJbr8iiIpFiT78a0DjozxA4KyyD2mQrfEo3m/zeG3
WBcKVV/kG/+TAr/H/DFAjvkNDvivnYHoPqk0MXkH5iOosOXMWgIr9hPecgVN1oC9kIjszIAdpyl2
98FT2P4eb7MybiaOrCaLuFzbNYwXvme/RICa+liE8WDo2pfwJQVft+p4Us1zPojl8LOkXicK9NsI
fwyGqzs4QRxo1v5sdDQYkpGoeXxaUWabacZyuSilfZ/AKJ8FymVYc94nrQwqCcAmxlQf4b7iNGmt
PyecdUatiZ3/QWhq+ThOxIlNioYydjJ06ksn2nI1HOeM1UMejjcF7MqADevHTsm0yn2Ed0K+uPNZ
ZWSXJSCD3QSDPyBQIqV498V/VpykPhlskpAVbt7KMSbQ8znSiyRjaug+rZ8b1i6pMzCZgEZzst3h
5faa+1MzA1STgR1tfbkDQZs8nK4/wtnxA+dbp+sVi4RZc950CnyNOStVahNp/+wd6SuhS8Ct0i9F
oeazzagPriykLveDGyBxruq9J3WRV7Vv3iKwTIvc+n4D9VDb31ASrHtztFuuk6KdAqTopruQPZoT
byEPxQ/Y8K6jOm65eqqewsXm0F7R+Hc0so3nJKSv/hSbyu3X3nbxMZM39Xgj0yZBDDX0h/HcYf28
ujmKLdqBBapqEH4V9sItUrPXrAvAsbnQegsfFhVYTQGrTpVHhh5JC85IMGqjT3gjRvWXdpUJCc6+
BFBhdd73C++RyJpFYrHceIekZlTSoQGGFxEw4G+k8MhU2eMISnqPIrGP79E8xrsFPQxpZ+nQ184y
+Acp12V71ziVIufyRNg4pfd62P6Ff8+/4ZFwyW7G84+g1fN0ZbzVVYB630+EoNolQQnUi2wBHfFg
Yn70U+NXWt0lHVoTbNIbgm2GfD52ldLM0P6zxkvuA1g+JgzbeX7qPmCB5QGMqrlYFRbhIgLwPaFV
9a2+0rwjidLoZ4BrGhpRX1CUTbE+OBx2SUSpJSIvkhCUytlTYsWqY8nS4z1PQN/+IlOPSkhzpDB2
LgrN5PG5R5pZZGErxo1uzs/s1xRbuTWOxCIZszjgP6gR2zjDYHARFaeJGTxtt7eH3U3Ss84fNaBB
APHwymmg5xJe+kDqend69e2NGxL8KBNwoNeoMgR+81Aldsb6BsTj8jDdZhLsKuX7eSxbvKdJGiyo
P6t5+JDX4vKqQdGYuJYNc5jd2AiOA/EtLz0dNbgoCJhM2RSVCZzCI+qtyRNazcPzgY782Wo5Ys5N
KV8lv7sABg/E7r5H9SnGJ6utXza0EUFhV5T5PiZfER0JyjCyUOQECcQrUWuF178E56bi4sIMp8uz
XpFokufsBoxs86/6A8E9FCtjSzJ+/NcR/cFfgv9WOSLTs52a0HtQeM96ugybjyJn4vcO+2Sykr4T
JhnTFonSx/kvG6EphXOgH2AaIHPVT8QqnDbwvbQJRnrz65nJaUHPtq3SDdFVtbNCsnB3kF9/dC23
oumWHGrGgQjpvO0q3h44LTYHpIhcqMANBZdVFKi2vZk7kAIpuNtZf0jelbqUg3IF1jFW8g3L9ztH
rCjrRuh9GTIqfTldL/0HiORQyJPkCZbYnTvXC/ywlQpUh8mZ1ZIcaEBseITG6nlGsirzOuYM2nz+
0iJVy3jKFN90z3p8zXwO5gY8LtL1XmgsmA4/R+wgogXyoby7SsMQ4XOTVEVR7hf7RPXZQYSstgXr
uQCFhiv/S29+u3kHpKQkUW1keqJ39aIsamJSTMKsErbm7HA1e6omuhzj8OhkmPmNZaKM814q9Fml
wpXkQwEhz+nvLPp/QNarmcfFWUrZa6qeVJe795LbdA7HCOBVEIhDG0+jURjAZazI7k9Vijo/7JsW
vQRGSrxBLZ5z6BCj2knbyLMKCBRKNsy6cMIxnk38Q7YbbQS7jj5Ub0bcoaWz87yTvEY6ZLBywzqo
vwBGXMqL7yMMLipan/u693+JAXQ/c8sWx7H2mKBlEP2cWv4ANox5Wdgc9UOX02gQGxDlelxCRj5q
aAaSRRgdZaJheJPSidwRntJVfN9KHzO6WmnV0WQUO01qBVfWDOs9URNzdjE7iLdxIAf4LaUlw/z9
gvl4xGNdq6huIhciHrfnThwdYEKpt/lFJ7Dz7rbvVGR2I2SEM/KI2WYljTYIj/yPLzBoIqUOO1LC
IhJGdfUz9YHZDWpgAj5nJNXYila3kC0fTle2Fe+iUJnKwuVYS7IiA7A4H99pTxv1y/w7cTPpWvAR
PxRRsrpfdjTXd1JsQUuW1LEaM9Wkxtbs+aYRz9zDIMgo8mzRPq1+k5Ylo8PJ+wGE2s2hPGwLoXXo
w2ynD4gobD7fnleyx25yyGmC5ri3+elQLoSlr6xgr0xItaUntNXlul0uh26EtHrU/FAk1QEGID+Z
rOBaVMEhJjqPKWbseBZz4tZQ2QZXmtZJU9BRt1hsLuuOkRQ4n20wgmCi9sJxSO6wS3OMIHswaJDK
3aEHV2Lnw3Do+jHxyG5qDaKxfzRTLniMWaGMz8gbPLOQTkK4y9QCKe506DNNiV7jzMNsGehf2SPZ
YvodCp477k4FJwprAtLP3Zejbnjc7mx5hfGBBCiadze5aic2ImAn4Uwnc4L1mcoTLqFWgT5E3z8H
6T+2glf/jjIZ3fI+/R8tOb2zPHO2tYratwCbIDNat+mszQHSM1MYd0RNdf5ypDUjlZIF3NazuQTV
SrGEp5jUpeoYG3tygAOMkM1tv+aGWdLGgqxD1KMd4qwwsqMkVzuTrvLgsHWVSGZhSRnH9LYTKwRN
lturacel7rrSkJVvvFjb5nDYydS0QKNFyIPr4JSOoyj7YfXbyaPaPArmTblBEOcXiRlJCFyvp7OV
ix4ufnbiuFlfgKcOA4aWthwvcTsiAc1OuheaUHACs/lFWfRJ5YtmEHCgwI9nfI90fs3rujGk7gte
v5xGI7RB7W+MBV7F3jyr/Vl4XBzqJ85vKeNP/q/QUpazTi0YUO5s+Gvp8wmqnaaFWg0pZj8DC9sC
Bp4daF/zOfSDmSiCUWWNdH7CuI0bSR1lNOVSURi6EQsAQnDaq6kbz/vRQp4pUtOazufN3MQGpGdv
Ip8S0i5CMY3LT3ZjQaEw95FJkn1R7BQV5ChR1RQ+86NAprN+Ps3cMG1SriDjtpN5eU46CbXw2HI9
QjgWKdmQTweSTaHqxYuj1FEE+ivxRqDr5j2fw9lZqFXZWUpN5z/jEVMj1kY35Ko35C9iAoVsGejs
cScZEAZ6czYjwsWGTxoiKyzh0yinpIaUfg6iAWJRC9UHx9eq/86qjFsREzj49ai4HCsX4WlZskQA
2+bRy/wc5TScj9d1QyQ4UAycXtEeuGqF6IbfxEseYCPxmuCE1dLmwZgO9R2xbN0YZIBbQknhxdPt
rA1Bs8o/fgxY25RAal4vvU0Wfv36w/HT9BhVn6W5+x8ywpaLAigU4uVVP1xtXSiM65JveGCnBQtF
6Vo9rbwygvFSbY7npObAYByI6smSRV69gXR1Xepf3v1iqpjNawzn3qJ84khgCKA5tG2os+LJgq/E
4XtkNy4XZf2L8g+0Fq/FQg9k1UUV6OF7VM0v8F/5dxARIDtxUANPZhby1A8wcrJKk0pgQ2ni8trT
hRzQbHTBeJRoPHIJZrfr5Dtsu3Iq/O1sc7Mrz3HaO1SjrBqvRPx+nSzoTr+6YwWULgtExlxCx7YI
Yd4p0LmipBd+ipcDPl4A6W6dRpimpJp/yvYm5ipv3m8+wgdO7J28yG4oa315MH5+Z/T7bZfO2m5n
Q3WH8G9NIKvWWnQuI8FwVHBDP3MNK029LqOmVg6KZVY4255fBdB8cTa53HorHp60VtAY4RzfNJuR
NJAa+ZjjA9lZbJP1jZ8LPhY8TR8K+1g3JVct6gV352bFGOkypMN2Gsy776jIJeGxvWCPu+UnCofj
k1Z23TxTIlQcWap6mq8Ar9x9vDPKWhaUP/hQF2inLGeq+IwWjFxdzxdRoEDvi5St5HrHHo8H9h64
jNG2/tPtKcTDKzmMcRQsJERzU12esxwJkEcZu93Wlt6HHPY5zjrxx5ZwU230fuIC5IgJ1JdYcuPs
yWoUjWUtxVZ2hq7fNUOpqGO2QPY8qGK9U+teyA+pP2LkxmsEt7C8+WxEmMuhM4ErFkwn4G38lv/D
mA1qKe1AF5LN/anGudM9Hs/K8vylHUgOHuUYdd5MZt/jVcUYx2dmCysJNYMAWw/+V0K3ieCJ6OYk
nBtKAOmZAJ00A1PA9p9qSBuqr8GOgk2WInuoCdkLtZl4Hk/E4qo4oIyApRGs88H8Kmyf6vXmKYf0
TzTZZgMws+PluKDx/ZUohbJOUfchDZ9rrkMI+ikzHNBlcaLomdvLgeLSrfb/xyFXJ3U7YtJgbwqB
DV8kEfshtXCo3O94zl6UgkyK6J/+MMYm10qqXmg9CtizKQp9fCikVp4kkt5bPbkuDGSuNWDK8Qql
x0gR09230N727C6Z4oS22Q5bitdGLXRcfGyV30OA4OM4PRgwTUKeWISNrx/O0UsBWyrN/svlXsZx
PQn6Ws4gcy+6fsKdNHhH50TZ5ZMuTdkceKC9PesYOMxzgB/RI9F78DP55v2zqDHf7QMY3PWP3w0W
a2YV7urvqYR2t3ExfQTf4nUEBtzYmSqIEF5h+DNZ7VcBKMeRUcq7a6Yf+zsGwb10skYMKSA4A2Io
VB1vk1SwlCW+HViEn4kP4eQi7ZHR/HDEp3Ydb0D2Ng3Xe/Sloc5pxKsMrrSSru/IB1ux/B9Uvjk/
d6ct5TJ21jqPu1RnfGpm7ss6BTOuerRiNHrER+U8pW4NNULt/wuS/ip+EnCwAHHZjYb9ngyiat24
0LX7ygeqkilHSHp1pZk54X5CoCXeeDJhFW6MThORYsWWvbeANv2jZg3iBlSj9NkD23xLDmcvaz69
EJqp9h6cIvmwe3qFTh9q2egMFlMcjpJMwKUQGRTahHuID6z6bhf78UIzY/l5FDWfrCDTKRYY+I4N
blQHsODYKrYKM3jpQWI8EB61TKp0E5ulo8NvaRAL6qry6FwM9ZMOLTwKCPf/XBGlJLqUdhmq008W
O4/3IUM3zo35pdIVvq3KcwdmEBti6Np6sCceWJLgkCOftBOBnXiGAPY9eJI5TL4PI4QenCRRPUYV
JNMMiK0YZDLhhQVucpwxbNKh8uof7g3S+kCGZElS7XjC52dy+iSjhOLcPmFEE1v/el09VKiWUY3D
xXWKckOLvrOiTzYaQ81drLm6YDwD4VIf2QvRCwMZIA91peGFyhKmkEnWogB55eFqh4wUwZTV85+g
TQI52T57u4B7l+Z2fiKCDaKjsN/2JC3mOx9xpWWNhQO/sJhGb6HiI7iqCbeE8mn1TwnbwbkdgeST
E6Ah2V7SSgH4siU3JtJNgKlizQq8jtLWJ/SmTTArdhYevOUdcD12MzKhKJVT8tE7PV3SuAJmsG9b
ldVJ6HeAvCptTn3/ziNWiZe1NVmSabBPk09CwT86QSW35nyVVZFDLBEbww2nMQIQveV+l1rmWYjn
Uy9ZGA/OTFCoL3LkzAjwjfVRfVQgqYgKSXKsMdcnR7VNL2anbvcwbuu/y8yXeexufnh3BWiQ278z
aVwM56HViT5ehp9mqwsKxqeVWrNyaCR3Qotq8KOYrXJN3AgCb7utCy8OZDIansy43kAXeIZAtw+U
JEwiqwBxgmOt2KikI60i7VzfozsgiZGb48XVQ6ZiIVovdzmemZgGXOje8XnaD9eUcNPD1DdyqLCV
gxENFS+nNT8rvAgXr8xuJl5cVrnnjzmwiZIVUl7EoK5agrhLuaf0NjRiW+XvkazTNbAAD9FmV5fy
PVK3d7oJ7IWZK9QqGKbL+vT7iL+W8M7fc54j/jnA8uKaoVv6onk3WT7krQRWhhKKLnap4Vk/V2Ug
Vvyp9PoDuaD40BHIoZXjkMx2BMyHtr3w4Z++w26IEhePb0WZVIoJT9gwXD6Ehxp4of44VYl3m/2j
p9y255KQbnK0ZtRxTFMGEoT7foWMrES36HAKcgdWGhTJk9vZIU92g+iW2gpmA9nBgZXGYKfde9HZ
lHdMZTJ9CWGINRLmHegteriBU800G7HZ27gHbxOE0Mhz6SbM2ZryonpVWhLAn92R3jyeWuotQY56
FGvGvWRA0UtHyduk20SJDGh4ZEhkEeMplZHN+sf3RWvhr5uEbLoUSlJOH1oy5fBgB2ccSfiSMg7b
GrHBeqwd77+stZ5sjey19v4bDue211EocivvOMClPLqC6iB2thu8MVLRy/uRSd1iDlDwUZ5f7J3r
Hx8rgJs6cA5aFB3+pvbjt86TxN7aEaDuSMAU+Fv6ekCejORhjpUd8TsybsaoZd87RUaWB17Frbqb
Q/25b7CD27JaRijHxNZDRKfc221dV9xtk/DQsp1E5S8he6cwVhZE21Bjqcwu+M5Hk74uM9Rw7G1v
D7Jgufl1+JIQjpEIvLzn3kNLziPhCtdqSN2M8ih7glE9x/UoatjtT+X/fwgkYHEerJfdKYqbVGKY
q7yW6T47ncOD4gq7b2z0PT2yZmv/Lj3VsIvuDK6iCrDH7+R9Co06TDqiYf02JTFArjMz5gZKis78
ADGtBmBaT+taBFJndfs795HRhII8qN62XT5ANHtYqo2vVVX/F/l4X4WAjCZxqPi3+yGeIcgVLzuR
XwxOs1vYZhjFi+Ejy42hKxeroZC/uxrXrZZL+0Ju4Vv6231riT04lBc2W+C169FM+Ilj67rQR8CJ
81Sio9R4zJt2xuqxDEX6+f5crNYmf6di1LCB9DRYqSZtb/sFNOfpqvt4HkK0MSo8ZJIVdUcGrn1q
E11gTqEyv1gm+3x+ck6C3kARjvrJOV1AHbxsDnbgBOkwdFBl3V1eokQ4xs1e2k5jSSbHhygoXBzH
0+PepaMCo+TRhiGbAUAVO6ph3FCYuVBmYdYdmw72GMrLjrFquSo8tjWOV3c8E+FYyUawoqCaGvmq
EiuhcQKKX36DAStweWLpPSo7u3p3Cd594HNCn0kPjwgpjXO2KH51Conzztd9vFuicXPRcjamP/Qu
m/DnwxguPb4znO1iixdi6r3SI0CrKWmI+z/IY3UgmaDIoNfl1hNLTW3/mOQpY+mrti9hwoh5DRMI
F9z2FZG9QqWVsY0q7dQRm9eXyILK6y5/A0XDV/f5ox8WH6VKW/BjUzv+m7J2euUizpyW3vnCifDk
zAsir+sbVrrbqQISxpS5MJGthvNjCQrs0HsdzsSjry9JY39kC4viqy7NB0p2gwhelbfQsecbyIIJ
dUXn2EQAb6hcrGx4yOSEtEDFnh54+F3bo1ekmknDW959NtNauz1a2XTPangCKIAGFix3OIflZGyr
k6mGE2+kLQf0MxLxju8bv/zGrCAsmpT3wqY80uRkwMi2IgQzsZrtFbkkFGXsdz/AuPnDdHDvYlyG
gfUR8bkOAEAZl4F/shhlBv5nJX8gtE5/X0eCIiGixrd9jojDVCqH0CMruiKSZx15ZpiNncuuVqfs
zVcmeG8DWXwObPDNVRDkFOnUjCy0lMWzmrnmPws/qdFyX/xSKg4D8Gsr+gageIT3iOUHxQMG/90d
cKb6l0QB5VtSIhvMNs/BGzpAkMSHLNKEKzb+duwb2n15XL/reHYDaRNWpIJCJhWCT74Dr63jayFS
wmOevpQdP9B+sbOaDRx1I7LT6Z9vUjxGpU86ZM3x9qr13JC6O+/sqdkRqgEo1dUM4H09g7QrDeDp
YV811u855gwd7X2kpl2NUxGrwq3XTBp42OMovQK+OMcG3RpA7KYp2p7eeeNXnBXSICgCWulVyIjw
sVSYW0HHym36olzVdOKVW3PxDM1dlRWqaVkL/ttqCEQuJLSD/aawjMHePCHgbfiPxhWTH4tuLju3
Pbp0r57S9ZKCo2WKx+r1bkjmDR7kAu9dHvuDDfc/EJt7Kopj15xd28uz62+nnOWMqIOf2hcz5uxQ
CrqqNhPDg4OV1T7FOtG1Nnt2KLb7WmphNXIP4ctg4ilu3SmjdgIAhyQLf+mhsSlm8xtSuYSqwVjX
toV21DB8NfoHX/3z+L4NC1y0vPw39Yo7lJJMS6jZyNkcA8ULxN0ekwf5CGM7LIsXUxNO4aL8q6X8
mha3Gwa74sZPkaDMizwmm7EPdtRd2NqL20lTICow9YEGv7qWpQlieN3xNB3ngac+1kuwQZy1RhuR
4tx8ee4C4XFgUe1QWnreeWWPJ6XDDctNy0MkqDZi92eB3JNDOVHD5saPV/FfL5w/cirR4i2G03zF
QE3XK04Vms09BlI60ELo4i3jSpdRsmBQJgbRWrp5iEu/1/ZR2fJC2sngxQgFJfmLYY600fNJsCXw
ReDMULOw9lOldlHnaiodq/RBS8m91G0Lh8oOCi+y42v6Otz85RfZOrkvEcPeLb1Ir3hoh83YTFcN
1DWgMYEBc/We3TXqAlLSc0vv5FCSQ8jg4vBflcCDz8Yv2jg0t8R6ZrKOVu1d10k2KkcJeUqgaCDT
FpNNd/9r+c2GrF7Dt1ig5tw6lqW/KUIB4DMjsTH3whaL+/l2LVmnjwYcU9bHsCYQRH9Iel/yQK2A
JaJlNZJFyFr4iSaMwQP921YqM4lnTJJfvCKcaF/5hDA3T2CpbnGouXrYZLGYCgeQbO3/s3QgIboT
pMs2rYWZk9QG1TOVP+qD7IyUW6aYWKCHRnuyzEwpu8KfVFpPf7rdHZrnOoplWIbooBnbTKqR3tOq
G3vvJr9B5jW3kS8C60kuyeJoJCRNzPBRPtn0xKX3T5fwBTHv7qDRkzugbZhIAMeoHwOQUHLA2/Ve
OBEmsiHMbj35kFy6EBGV+qDNr9rD4fJQVLfoqzIJVTYxuOyg56BNZ/imLbvX9oXfat7FBCn/GOAe
d4sp6bfQy+EmP5z/Wjl2Yqze6w7XviE98BIHssR5VItM40pxckCm4oEIlKoN+bVKghupvP5/dsmR
C5fpRDoPN+BjvKMBDntWQPlTTOyLj4M3s0veEEMnNxxiNpGGYx0eKCH2xG4Ys+X2Y5zAh93T4NY5
5Kz+t8glnW2Hy3xxXt/4qeu5/fCivmyPpt6CVdxNcAMLGgbqRHMsv6pEsKypj6r28qHVFRSoSaZM
cUN3SUbEs3HrnkWzSsGV6GARFjsMRqJQ9T6qt9i42SDKr1J0YOpJU8EIVEOBldf7PpNsgzc8po+t
tUZ5HLrpwOM1A7XFmyZoOZpiG2385DI56IdbBZjQDivpQ+Prz11wi+8yifSeW4P9ngLTN1ubohvN
Qs10VCxV9xZ/ArAOHXAOuRU7xo+QksyUDpqi0Tend8rq8nZ2O01rUpTlLUum/+DcOp9uS4chUrYs
VVZfuyw+xVSRKalDX2UVY+eOgFWQ8jWtJwapNWLFp6iAHojwZH4LOBc2XWzrtZAfBxjan6QCBMTM
WIZ/M/zt0Ls9aP4Ur7UNb9mS24s19zUoxce0T9z7CKoxs3wQneIp06Oum0NftrwokceX/uoMlHcB
oeVPfqe8+tOTbPViDGGCh+uh3ysEW5Q+1wTyFhU+C4DWHVut0bBci5IhJ6hlUJztPVfQuYaBN/aT
XZm8L2y1qiD4eLmNr4/A8rKe9a2D45rwRuV0zubHkVQlSYz6rko/KcZgXAReTXoHefmO0BLSw66z
9JPPgPVZhEmiNsYrB2puOVQ2TtR42G6M8AlXTGDuZe1rEgeFIhksLk8m8p1ub4Hv+TSPWkisittw
STYoiL4s7V0LPSvSoRPwarBC/BAjqrZBtm0QP7Yd/k4TPb0nNo8/vygccOacGKKogSwIVE0fABd9
6+5X5zoaqOFA5kNdyM3X0Jb42x3Zlp+wByERI3nwNCDTOwBcUADCQfWF7Xfqcd/tvxBa/5PV5co0
sm/z3lynTuGgDVNhh8Scy0RZO3mK8sXl2BiPejvPg6Y0/crXL/Zy+dhqHzlBNax4/beHIyFUQwYf
ftkoT0oAiLrNllkDti0NROxonI/oh6JdddrlBbix/WJmCHin6e6B8uqI07UaN66DC54ccfVaFSXa
bGrjxXGR8Pb3lRTC4w+0X3ULR+UPvB1FZJShDw9bi4HIB2P37J8KILe0i2fe5IWcZKd8jSP+OGis
QIHHpQynxDNq3t9D6E6iO260bFS2FeCImhwg9Sjm3ixBpeASmv3efWT/5zN4MS2qfUek0AAaEhok
8VLqHL/Wxdaxoa2N3+Snxq4ZevOXiYrqMKEPXXOYcNpcPhEvgO5cKlCFa2FhQKPa8waT0HlwNwih
3vgn0tFXmDEWal/vdCIZjUW5q0fULwMzKHyf7Rexp5OMNTU4DHLeiJfGup56WKU3ctWRxXk4pHU+
wvBtb+Bwte/yqsTdg+BbCRVl7EeJDJOcD/+YZxDt4WVTDE35Me+2SOHkDvfdjZC3soVzybQNKO71
caKHB3pHOCpMBSXvkwPiQxvgNfPYA56QjvORe26H1DYds/R+6GB8EnitQcaNyf+TmA0bI5aUVU/u
XFb4b2LZ4Zh1SqWaLZ/DQMBtDUz/4MJd0yc+DU/r83y00sQoM1xwwy5omBofqW3z0j/srlCpoF5f
Z28lnUALB0yJEq3gWy15ZWyuRfxgRHczKRAHKZ+sMX4JskH08hIkMJpzHQEXhoqV77zaCAxtzs8E
WnlGSIQ+z9PNFeYqP2IkXI2wp2p7iqS/TyNSnsFUy2oc3zYWKHc1IGR6sxpPT8Fz97Gh01qrprJE
xvKWrSg5bY9oCI/Grrv/nCNgRjvM5L2MSwNcQ4oxr3zeo/M7b+qlX19mzVfiAxCedAob0gvaS6FT
3BX+4zT0MWckhMRNDSRb85+j2XOeAk1RSHZnTBalwF7fgEM82t3FJ1Y00zRVn93qn2tASVaOGk+E
97YJ8Ok16Qvuz3Rml7KQdD6rIx/rboPq0NyzCHi2AKLux9aoC37ZZLNsbAtJGwGxHdCJ8mwzLlZo
WgZ0AlcMeQitRQNO8tAVBAi0i5CC+ulJtG9vnEDrenxp3eDL7IS5RIcmNYITwzmw+dW42dFLzE2H
sn24jl8kGUN6DrVhjADM7G+x5vjD95aY6tlx4KylZ5Yuh/kYxcX0AftjMBsNcT/wtLxu2B7+ocRj
5HLlZikm2nImZy7d1r5y8cu08xEQ8GVT07nLL0fDRmcvqdMSiJTC3Xg3cAzQU0OqWHdovZoHASd3
2DsB0Vo5otJJ6kLrivvap8hEUH+4K11s/D2bYQDeNVTdeiWWTkQhxB9mQ9yxJmw0PY0y4m/tFvJ8
knRzUpK5EPk2og2nirK+O8KknfglILEMkurf0ZtqZs9QXlPHCTFSBRgTho9nYD6f8MgX3pO7xMtd
SWZwrWv6mwOfgBbkCjKHd02h4ZMWsTTAi8g11wfcbTQIYmJNG9hq/lS/nLKgtLWc/mTY/pfB3sGX
Kx+IazgNs4LDTpzkwSPDdGuZYAvvKiaeCDg7i7Ia0HIpaMdy2C7KhPvhsWIXz9jKYgfP42DZ//7K
un9F1J27y6rtPq3sGBXAwSyLD9qHg/2yLlbxHqv81Fa0RWkG7/NSRMBaDcl1yfBLuiALozHGPeb8
61q/bJfhoVgmkGjJei5we05xgf4V1LaodHmHhwPTn+VvSA0ik+FfxSjJI/dvL14EIK4GlDnEjqhZ
SfPxtX8xqrxkHfGlgNzOLtCOmNWCzxcSV3stad6dqcn9mzW4RjmrNFzmBYZpgV/p+ezeFGLx8UJJ
v1RFr+MdL19bSTUcLhT2WNFNqihM/bhEqvvYQ3oA+6OgSqVgECybiaFJvSwvxE7Gk8UHYVxWfnNb
MZhxPc9uJyGRklTo/xd8AroCH1NsYrziMqR7dL31+vtjvSsTq0w1LRrptnu7roL4I08WgFwUI1Ex
WwldBo/0n9SOsV8mYlVGcQCwnvzKaj4ughCS42VBTL5Ye37uJABVpNe76AS9qvpcIzLdpAQmfRsG
G0QuSjry7SDR2SZ1e48YR9NV2kYzBV7P4Ump4tm587+bGLQRQJkgpMTyn2BrIrP2IEbn35cpbJTJ
3wN2ExVtUwz4idgHhCll/taI+VSUYO9oD1yyFRc/8sGhN9voGWYiBns8/Oddhx17kqkZZVTE8cy1
7AfDhS0ovfEkNG/6yvwbz7zsYX5l6b/u5s10dgK5L5phTWbUTpzD9+nVddI/gCBXz2NcQ86Ut6uJ
mhdgsp6CPDDYflv+H+2B6rO4jjNbSmAoLUHjGnKZ5CfuM+Jrkr6QJtKDtj/KTl9BU2X/v06Yj965
JabxDfBIgm+AJokHCZ6O7oTMt8SHib387ArvunPvEv8KDw5KG6mhN+KPOmkGt5vqNLfsbhh/Kd1a
uTEyGpLhXox7/oGC+idY+rJ9NOdSs0aU1wau0SSUCDZSHsa1zrMBqXivyaKEiW6VcmWvO1fSGvOT
8H+JrmTwRpl/WufrNWCSm48/jS7tDIgcVk5e6sWtCdRADucAUL+432bY0soWFb/VlwWhHaIzVGiZ
6nDvIY539DB81CmLkAYNRmA8aJ3OHzS+E3mQvPWP73Y2tjiMcy1YOSqoKxVBR6d8vqpnOcRbb9SS
Q1ttE/TbdIjD5fZye3G4tyl2rz3LYU1q6CkrkkZHVChGvzMXrQ6nyIgOW0gV+SM07Ubv+Gw5yHT6
nCKJuyq0HCtB91cd6DED+N/d1AlHnvBiaCgpTUW1S6Y705lHt+h1H8wfceLtiWrny+Wmi2hCiDmm
65nLiX7Cv/g5to8szPazSSGgRAt6Pr3HSmCKGhCL20hn9K5HGTbIhahw7WVCTLE9Fgr4KkcwcVzm
Hlp9ArNRFzZEYJy99q0UkvEEA4zWWBE+V1PMLJiY3nfastJtaPA/dNGlqSjliS1LgEvNVHDpA+mB
nWnmgBmNnB/nWxr19EV7estmNans+b5kdEiBF0L58NcSKHzcDxePuDSngSZ3cKrKZmUn93TI/zvT
GxCwn2/vfWFYfg70tGSZYflozZKazyJkI4icaGg7AB3lH0zX1vClf981SRzD88nX+LCq0WixJHqy
s8FGsExLwhFemRWpEQps3XSPxqhrXw84C9VblRtmia684b2/Nob4iksKZPHms2bOlU+uPyhUuh9X
AZRCPRen+8FyawPytvWX4yU3+oMSFg1wgQ++pEI9g5vJuadE3bXwE3N0T3o1ikDnePsL1Px+l2wU
rHs/5Chj0XunIcxBvYFgssEDZVFOBIbuarWsf2vREDfBe3thyuzmOFSG6mE2dZcQIqjuz06rynSH
0x0NBNfUkOafGzpGwBgyiCQQMg4r6Mf2HDej+WTA01ehY+C6xgBlkMh7e0zrDqncL0j0NQ8Da+Fq
glbdbm1Ii/A6VFPAFxIZTE4Oft2bUJCCPUz72b401SxOxRNtT2mqEzMMEthoaSzl8ig/uOAfrP+z
l9P4XkPO2vSONqwZJLOSZWY+MN18aVq5q36exiSKOjyE1rSEnFeoQ2FOoZfrugywZKR7RAWraga5
qDDRNf/m6pq+AfKutkv4ngoWDr/FOyw28+OhpA4ERVeUlmF98qXXZHejWGs91Ts20mHdWhA4uiG0
E6yfYjTrZfgM7L1zlc7G2SuqwR6ZI1vgHl4bDV/uT/UlpZxJqa1iavLV6o99cRDJ8xwuWhCpPpcG
3IA/TKjZxH5kh5UJNPNas1M/t7T1FFq+sdt/NRNaJ630SCmEVjztVykaXLA0MNUsh8lsTkm5ZuLs
Vr+jmTKqRKsZd9zSLOZ3t5bSKcXjKNDnHoLbNojCHkpapD3/zMNTUqpLsiL+4Wv0x++VrPvk6sfj
bzXXHqapiq4qhHTcdmQ+kFD2QUtynkor6p+R7QaUaEB8sYgsR1uHPe1p3RFzX5j+SOdTfzkJrW4J
gE//UEvXs2TfT3flKMlo6cIGuwri48Vr/yslFp0WnPP7doIIKThIZTaIt2w+WxK+TQt+s8IARKc9
mhy+DDhp8IPQikSfeKwGmnruNbgkfaXETYLWaoluPVF+24PTri4RHKVCVKFyK83SZRIuiqUBm6RP
qqCShXPcE8oLbA19N7AEAtV629wxXsyYh6JjGPOkZ5QC1VLOD085CwklnIo7/rjLz60yJiUOGfaf
gwCdmW8OheLPsmCA5/PPiHYGwWT3Ghj4zn0VgtRTqE4uNtHNBWktgS3x+W/05xhg3nKCqaUlFFhq
shuIUPckGpTJScWHo15IpaOsCYcc6UrGFcNcMCTLivB9tlwo089b8fVWlChubf9wrivPJYgbAOKX
t63+IFYYsvIkj03i4bprJOmQpxXlICcrjE4o1jJxl9F1TZvNHhU1SNA0ZDI9xpWEoAMBIWHJvAKS
cvNZXijXN4rfava0Gpg/L0nTt1ZBuUSCgHfhrY1HFsZ1gu10CG2i02XYFsQuWz+ceswCCat+D/xN
K6s4T0fdDbo8MJE4MBffXh7XkL/IARetrQnofOvc3LbQDjf7xBMbiz2yUwpYzEd0Mv6pXO2Z+xQ3
Q0lVmkDYhdiP3qhbnYp25RGHMhxqF/2ylzYp2m2GMvgEpVVWWS5naOyUdYE0ulDKTdJklb3nQFTG
sSeUKSgNtHDfV1hO44ENmaJF+4F/m4lOxaTGyrb6jkON4EoSZBLXaQwwV7pjvCghuyJbh71y/Vlc
FX3L3ZDdgF/L24SIfquJmD40K+KaW6FI1X3KaLmE8tt6uChjceEwCaHV45VkrDklUHs4ogv4iUnX
rlEp0lsH23elXufWMO9P3sfUIQCmHW8WozsmfyzfqeTmZWw3rvmpAK+rA3ckaBSXIfdiPeLU0pcK
mnfYjW93+4bBEshVYHo0EB0PbM+zeKWHFoQnSBBB8GVijTx8nANKEp2gkydDfwnm2vRN5zMf5un5
ht3wXsBYAQ4a9h+az18hnwYDdFkNLsiwb4KoI1YRXk3YB5did/WM32iQ1KDjpsAoJybTqsML5B1X
FW067RCgXXlnFhZWLEO3i/ONKfUG/SUx86BghojrB4OnM4CizP3P19E4Ivcnqecjd9hwdNScTvfC
Q4/rgxaTfYva+dxdOxTezIi5nIeimPaMW9D090ac5hQn1/eu+noGV6FKpc70g5+mQJqJqRnUunZL
nBcgthZNzosWieRcpAccJLCWzMzE9Nd1BGTFK2nDnCPv62DiqQ+7sq9gynE7agzpXQVzdONMy6sO
vAMmxhDMwSaQY0mJV8WhDO7h5F951vSjyslFcKLsv5aqCsN4BJC8L3fLttEpEraIGePvQqcjP94R
z3vpBlGpUIJTywOz6sTNPNzDcylKsUU9uY0IUwxRFUtO2InE7AgUYltCJjJ4nJvkOnxdCy/EVECn
/BZn3igkHVCLKWiaT9Q0+V9DZA5ChxPSv3lV2W1EQmOfYS/6eXDn3skk8h3EryJ0+V09/u+6aopr
vrljR/NDzUejDQETfUPjtB7lR0VDrTi0AO/W7/ssjURbmVv+sM5uE17hWp5tacmp5cZW04WAuniv
HQ5tkH1/JY7Jfbrjp8B0PmAzi5HyPGLou3D6FJ/hp+E04EgKE94jStkxrJlb0/2AWM69Ai8HB3nN
eTyAjVpHxsWFwDn+UHd+c5kHHQJv67zCt2khJ2oVQRuZ/qdB5Ee+WrAvEngvz+qDbxK+LwtOMuAz
v9ocMH707h146WHfTJnJQNfXm7AehBhsAVerVE2SNaHbHV9YypzCO+rbCpvMTdP40Z6MGv1qrFcj
5CxQXMPqEmZeCxwRKIk2TZlc9zb9LpV0bj3KZIXPEDTwx4evKx1fbfGv+FFAB6nvISudPJaVgDdP
ImRVZRkbW4QAygQsA3Z/Qo/gbFOr+Sn0qy8KuOtKotdZITHglUP5PMR1co7k+igdE3MUrFvvMPXW
LZFYvXyJY/vuKfrF2hUe5KgQLWsmJ0Otx64SXN/+cVNm/ZWwUIKjIJgMdR8RspGavdshMeEuppbQ
2Rgb3bj4gGNPAAnIjqGmnETux98YPU/8idoJ10zuVnZ51yqR6zHWDd4VssJjrtbLKtBloe9OHLbB
5RiuRhd+fPZjeyr4EyLst0SrRRPRFwYJAkd8oALLd6GeR5idteYzN/Sx+Cp7lS97sZucKGhOfyxF
6PXqd0W/vy5rfftnkYXuH0pUFctSRqwwydj6LLR2MyAiPIV1lJYZAs9cn/ucNpddVqjnknSHSjUL
VMUoanC9ToRqsGUGViCm7PbLFBe920vneCBEGe72BLgd1koR8gUIP9k4VdAuuirnyasC2mCkEoay
eysPVlveaGetAGThYOActOUEGj+JdxQBh6C6d+jKqfPFxl3o3x+52L9GyimoKW56l5Trafuyi5Cy
Coi1xPPMSPUH9acnh5+DMy+RbHxY3BMQ+WMk3lk7R/trYCkIaB9M9Os0zpEJAR1TAPD/fIz5ruUx
uTwl3YgFfaO6rz47Y/EBVuTT46n8NCzHdQNZcA2eNL8EauhOqMXVv7brcYE1wYZrItGRM5I3Qywc
d7DGTF7urGG330KPLeegAiXrbdfO64+OpblfqgibKYTHwE9VLoBk7k7sK1Ax+F0MVzMyCKL/yPdd
qhzU5/dgNS5XT129cAbZdp3lKzyyuElZbmNx1Ev/VSkUnbK9lBGB1yf1eTXJ9fGfcMvf9+QFObKD
673GptK/tTXXFjFh8uJKs8mdJrJ4liyDrYwlanslS6ZtjKw4X487o4U1B+lDjvN7MzHhir3gBPUx
yg4YLWdWHlz6rYeibsgz/AX4PZ3rjec0p9x0BbPimF5I7cemcRwRgsPczqLpdRTw9AFrAdWxaXes
EUq4ZRYKr0zCV244TiMtf+zi/Qwx7o/X0zS5NRCfgSxQU3aSYvs2ZoBJ/7GgmThDVrhjhyivdNpS
ox/PLtFv6/YfhitubQgZNB5hoZpbr/fj3MFmwJPQ8WobNog2KwDmH3olEAqUqye4HPj8uCri/Ytn
idb1X4n90dfh2DePFJDTZrANb63bmXd6ZP6XMxXunG8f51x2Wxpuz2UrLzODHNta9BIyECb4ajGd
iXxpljGBoBZwO5gEO+3XBD08kBZpk/yHd4oeV/SPPYZlPtLJjRKY+8iXz3TvaXHLDArE84cJtUja
9guCehLUPuOWRmglwly35BKBO55TbyQuHOXSxkc2wEjv6Jmwhs5mX+TCjfJC4RykXUcaWCU5Zuci
iL2f/BCstCygBzqfH0wy3Enj5t4PwDTZ5GYJHDP868VmhwOvJ+E5Yv7HAbzx/ogc3wdAbQSW7Vth
g9VdP1E/06FH9fJjyBXAah4y6aDrOGYrJ2ezSwF3B3lnj6SQK/Hqj7Y4cbQ6YeiaCafdlA8AHlR6
6WDIefI/Ch9SQxByaz1N44PIXAzWTDUJDs0TbSn8Rtc9UetCkQsZeiEyoSl1s8DtbAUQ9BWl83Mz
f8mFrZvUXVh3lP//u11Fxe+3C1G0TfvDZJIKhRque/G1QabFFt2G+30ICGxS/rJjqlZ2medXhbGW
tbhbt+Wpgxturtndff2XcCBEQlmQUlleHruT/vl5ZQp6mFD8OPCNdVxOshaDF8sF9m13qvZ+V4wd
f01WeI+UqrGxCDuNnWYt1M/2OOUKwBzzq/HAWKdhM8kbWF/TCPZwuzDUy/Z7fvTUsEFVFazN4RGP
BbVyOrSJor0BFVJdT+WPIphskx37WPlWtLfHVScmIzwJAvINU19V70Bw+dl8ysUQbGvsQgHJYYEb
xYPO2B58kVKgvi8g+XC+378xJENDYChGb7YW9Jr5sEdYk4BkQsNYKweml5D2090zZC1tYBM1EHio
ze6KpILSKoopRp1CoJa7uueho6rDLVgCOmpwjfsQceUWSyvwdXI6qyLmNHDd3XsKcX+oTot3Ft3k
A/cUQEFeTMDtgXlmKxEWTxl7+ppw8pa4+BMnVyXIy/PwT/+eiSY2+KIc2pWTrniDok2MVgRcNf2l
n82iMPBZo+lTRdj3e2Hoff0y6Wjd+etkGxklgmGEaxdw7/hfyHKRk4yWGUEIDXFKz9fd6jWR0SvX
V4u69wpTLbj/dR9vKEvZxJxnEFSF+4jv9Z417S2jGd0p8Yqd9ZnCxe8k41nNf7jtyYlHTvfY2Y5c
gBp82aH/7k3QqcZj6NthJrfnsvLp7G6JRi8gjTMVXboQ8Z/z0GMEPaRY2kHdljUGBLOgtVyIVQ79
Ld7Dhk25oLyTwLV0aqL3r5Ac2oOZBMRjkyZQSCjnP2edsvJ5UM5g7xN0csAe6lTSLjP87uXHF2mU
PiB8yaWcKJjTaLSs31WIHS7G/rhEOuPkhZMFZ1ElGpFHfTad02c0xqOw8meHP3LNPrtRTGUiB4F6
iztAbwDpFMgnI0p3E61011Tj0yhoxq05VHfxVX2AdJiNrHjKwALRRHhqIWdmiaeivnv2c3oEWC61
82CKQdSsHcsTKR7z5xNWRJUSq8KCDLxkMheqn+QNcyle3if0dlXwlcidOQHfFJxaPLmm7skqL89L
HjfQe8DDZaxc4Ub1xJgwKePA1SwPNxyvP3ibfOzQTGIF0d+RANT4iOtREGbDUBpJMr29VETm9ibH
SIlqaMfy7nFx7jCYhHBAyGEBzAe7WFGqAVejGihbK3RuEsq9vSTC3Uy0b4RKRa91/bsdddeKbt3i
M0Zq7GxYD1oSDmSfihWBsE1c4P8PwdwjJnQW5ZC6+BkxAoBcp/madiJ6KcOCuya7jiaqgfo6A+Xy
a/DnHjSygXBCGsn09Cr47YEfUPEG8kgSYebEFRPytys1nfhHbTVJOLlXZrS3h091dpLmqsOmnzia
hoWXKE1FwIlHaXR7Q/489YrZBY6RuPiNjGarzTSrtEjVfw6WRoqTUz0k3wq0i/WW/+kX8EHS7WUR
qLqfY9TSqtmsTMo2h7FMKEUcGDpvnEMGEiwJHSJ/P7IkPHmu9trfd27pXn26B24JCnOF9F3s4wUs
e3VRbfivFptPAbfO9jYEIMbUe+XNvjvhGw1S18CdkwghxHV5J5qK9JLKpZhtgc1yDwo75pUvHwdr
IcuICtQXdhUS0b0S0A4MARV5iKhdSA/vzYc6+4eTJwt2rUXtdxSnAF+e/+93OKMw7RDrvsEEsjVW
QKT8mwlrYwH16tiB2qmK2FEbj1ld45XFYowo2M4rUvSnLteP37+zF46u3p1FqynkylGsr2fZBEes
C+oePEk3n6BKEVcuNaue+mT0FO6nnwWzkAEGKJNbo3YQMK83ofDoBPS8oQC2wpgDHdNZYJIIawUr
+I/wXF/p4ezyrKBgU56/8z+gqXW3hm1/O5DiicmYDzKID+X68sek5QpykHCmGcBe6YsZj/8rcI7e
+8IF3cIPC+54w/wjY6S7dwbGBZoKD5OHZ3GobA6Ba7/KdJmqbcjbOsTulquesTDaV9MPiulrlpIO
hM8Pjfi0ORS507xdqkevFt5pRmTtM+w/Vmhzh32Cz+5RRhWNl4McDNIV0H6PSu1QFH/vgn62AFg1
MYNzE81N85eyEKx/+H0WEXDMsvbqAnxRKvm8oyi4yt5A/uJ+OyzkibJHghRuwLmrZw+FnAXn0OF2
pXzoOOcFUHq4/ZYcQYG+K5Ls24PEFGQufB0J7t6lrYivHtayVA93qdWCZs6wITzWy+MNa2NhNWUC
oK/3L5E7eotqUKR+tDMuK45gr9z5wZWXjx2n/qOxLp4SPebn6rvGLhRzySh2Pqky1dRZEQnY33T9
83eIqAfb6RpDqBnDFf+yLMg5ni1vYQngrpy7///1a0LBV2f5gB/z502j5E2D9PZyRtH8qOSq4TjB
K4iAz3Qp/tXjrsd/V1Bv71oVPsR/zQyTPZgDuUoGbQTr+Wei/md33oVmSJ2BCQHhTTIm0HO4eJeq
wzN7nJVw0L8Ebm7FJyBHNjJQQeT4Ob1Jrs1DPOuwdFVgrQEaQe7oWx2e4AHE4viT9NkgKaH+y0i6
etquUG3KYoE9jxiO3o2XokEV6GtHmotT/rwqTEeBulJTKkTCe9ocS4A8oQ2BfO3C8sCgz/Exgi+J
Mnhagw1m/gHLBLZ0DMTLSp900jsQ1cF4D82vYcUQV0QVmiFQBRj7gOm+v6LJCDdCpnQHdud0CrqB
fqBrpD6I02OjmaS2NLrpSOImb61PALYjKHevAgbKELzdzbqzW/tmGWT4LvNtNh5V3a6SkIZP8fTA
y4OFygn59PowQtKYwieUM+DDaBsCGuVZRNazZ0DIvpZYCSdvJm3u5W4KJqhm7IduXpQ9Wru8ZaLF
KOf2haCN2Ry495xbz5koWL9cxMEFU4W0uPWhdmyHSHIt5Jc/FsGTDdmvYaOziPqUWjPOLQhiOCNu
HAqS9/H14KkeqOy2C7hUs5gQ0dEvKKDrdrRFByHbuS2/p6pAS46P7wWOTztKU6GoaPVVqIFQR9cU
o2ABBgFIkzvrdbXWRBrnmuWbvaByHbIg7Dp+I2fu5IEwK3w/s1I3SZutxPvl+kB2th51O4AIe8xv
9P77ENGSdIGFJ0dcsBZEsemAj6wc8xheia5KFHwU8n9XkTU8nkmzpQ7RJpjjsY7F4vSKYzJLPbRA
XjPiXz4llJ9FH7EwWYGgZ8o93EhAMGPFU8pUskndHNmx6tS/61YrLbW5c9vBrhP11GkXVE3P564k
2dzDupRisZFPjSuUwX9jJnQdu/KCMI48BSLyVAesSY43gBHHsocwEAjB7HqyYw97b/oO3hrm6ZBG
hNbTC2geiPvlcnPVULPTlkMX+uXEClJ/hU92oI/C4YAjYcOcIta6J/bj2dh7HLEoNtxDF98OkVKk
X280Nk+oACV5ueMuxSY0ChCrGFv0BoA4/+c9Bvt/7CT+VcxEQH1ukHifdi5cGNsYbsWtFxWjA5uE
2sJkNyLT7utlT76hQj25AhSEMoA03GxApEo1LxIsQZwdfT1ksYfASqCUbO2hKWZe8jlBqsxYrfd+
BzF9ZmmAtwhcQSDZ+nAWjF2k8v1pUoKVwBpkFIX2MiAlA8xbRssy8ddIdoImd2T00oT34Uy4r5bg
9f5Y6siZXD6T96pknI8W4qeaYPFMiddYraahtjptMJO/cKbC6piFbaAmoqJxNYdUoBWphzwt7WRQ
MCyOrthCmHHz1iFR4/lnzMbLibOsXnHu1rjQSm/NRZJFuyJf6fL3ah2E1NLV1UgUKBNJUCdxP16c
Ww5MbDzeEVJrSX4yTb3TmT5YM2XVWdUKjD9WucGY/63XcKBLQhG9IPqQ68MyKwtefh4Wcz++aubs
ktpbYYtMN4ZGBf4K2ddD8bhuWRFvr30PqzngW4ylSUYHzIGOlo0mQag+MyXFP1B9ZwsZ3GfoblRZ
GA31f3VDpIjTrw8nvJPQSVcOh3Y9/kI5nEoc1Vt38UcMcn/EsZnhAmPAqdF7AFxATkqBi1qFlfkA
IeTffejlSO8vEw4rq5RdSz+QHoEIlUt7qJudqwTBc+sBR9j03eMgOJVVXQRs8YweZH6E7gvT6Dzd
xl8o1LCALgWarzBgUD28AtogX8EUgPs8KMY371GZaLmaFrB3lPriCFyDg0RAINU51pkCBuifUmbk
LH0U7nKptPRPj6bO8s1MR2HQmRXCLNbzdyC+cXGwKElLFMOmK2fKeGG0rKbHwpegHPf7vP/x5xPc
lk0oBQeTNxJxwsHp1/nVot7h7HEASDRxds/1XptAwVhx/VWSmH7XL5W5AMW+tfcrYEk6OKgSJ68I
NoY62ZGFNSVDxGnR7wsaPxAb9b0q/hHfct5z6OODgOEcnP5MzKcG9S41RKmsIwzRMAUzwWkhL2F9
ybmuUd8KiEw2JvME2mTUeE4nyliiq4XnxAUQWNbG8uTshWSakbOyobpe4+YV7v1+P18OS6qD/3uG
OYKlNW7CupwyIZjMf3bVVS4EW84fdIkTXFhs4i9th2PyMEw7z6TQMCQunEwgiQPeViUgotoCrSCb
riY7FeDVURdln6jXwXaGAaavA7TeR4dg41NFn38daUDxv1kburbg3aveqmlUZFfTE8p9WgUYz9yH
jLFP2RTrMT88uv45cBPxJAM6GJlbBKKroeGb5W1V+hdh4yz8hLs0xgKUOSBddPjLLRawhmheQYOk
6nh6cfHhcTZCGA0NWHdJ0+DKamymY4mo6AlsFq96lM4yKKGXQkAl8pGtSG5cCMw8anCBqj5WwVcP
VRy30uplCMN9FYtbvQapIMdV875R1jvyWu6YEz5N388ks8w/kDmr/bM/EGz4qiWVO+uuwFtHucIG
q2SnWnPIPvbK0Kukkb9zC/FgFagUDVeDx4/EAVLh5qw2tho45noJSwLCh0YmBBqWzGB5yWWhc+sj
AHY3RZ7qtzeE28iV7/BZD9nMMRcxwSEjwpDD4GTgFJr6ST+Acp7ZrZqi2hb1grhvOKYmzl6sclGn
OApKXTBtELJ5koucu3NIgTHWV7EbdwTfgWcbf6HQXzJxY6VJtKGHjm9c+48MkK0bBDNWRZlRVmSz
fF0BeMsZKV3txfdBdnzpolMX+Wq9T3kGTSV5CEUAL6KR3gye4jKIbNZcxoBAOKzKvgNpn6XSyy70
99QeL42Tu3MnObO1SA2y3aL056yMj6XbRiJ7TlruLhfQ9ZCx/EFo0kwIU6cTg9rObWvPY2xDQdtK
1nbg8chIgrpnao7D/NaQzjsy9PyCmkAA2TbRQ/vHNxdHxv7Tjit6XFh6iEilsnuUFXugqkGDeq40
FUaM9BInSS1gigN7XQhfTjOosA+SL9msO09C8+/PBaGxG1kEH2JL4LdvkAtQgEMvFaTAvASuSHpy
dr/W7wFmMWxrFOi7/hvQKN/VHb/HWeAgJw2yuQZlQu1o8Bd7QuI8ZqM+cQxddDXugMZcZx/ixEET
9a+49sC8WUTj2v9J/SQkEy0ufkYN8bWKDNnMixt/eLdwnjqD2LVtMbD8VbxwDPvm7F4TP8lHRKaX
vVCGo+3fQofBlCF3QLp3kXQZnJxZCiA1sPRwDo1ODeko5JeQalCnM4eX7JLyyycWZ/MilS9/40cs
TaJpnVdGKdBe76z0YK/qh8bk3SP6yqp3j77BAMSkbiybPU0cxAEUzEYcXe5W9BF2QtMNZrQrBbbU
zpTv3opaSe0o3TYMff5CMkzg2nchonCTwkmOBn8/eKq1IfDfTa8JF8Zm8EDZI5RVlKf5orKtgDab
rQlQ2fazshlNRe3igpS8xoTGilwL5bsN2InSNwu518/LxbNpIuO14d5SWgb9TG1y9lAG2R/qC5WP
0eLm+EfGORsFZMVgx8KPI5HrwRKn2Kqqgc6X++JKbDKbWPGMJYaP2euiPt5NAkqGA5jSuBTWKsZ+
LCDZVs0skHHDcJhi/xclXG3CNg+b/ubq/B3/b75O5jQBFC26E8AR586WHRE5XqjQfoybHvkHJyzz
ia198CG19o6ezOPpfLTrEYzMSqjruwd0Ig+duK2KNAlbgGV5o3CBYWgZ/GkRe6ASAGnbJPQ4LYAa
w0ZESyR4u6KYcbEIEL4URSl47HIk+BJojwpFmdqBAo3ceGmQdMPfKUkMoYFzlPLWJkXSU39IjLzu
lK+/385ltrP3QWQMRGFwGs8KmiUrkDQkuAfOgkV64THJNwjmCm1sfmY6X9NGnGevIjZb0n39IiRq
9l+aKGATOAk6Nv3xW3bpUaUAPG/O5R0ra8yWmeOACqifUe+eK0qZ+J/gMQznCT+Ce+L8YvlMln8o
LhKqEOJUa13wpWbtqLvYNWCaioyGyg4Nw17S9cwrQOwjhTBBOwBLYOuVJgUc0p0zsv46c90Qfqvq
1kYIbWpnICaVDVPDVmSOv6nYDV4aqBDbWl+zc3XFmOe1JwgsCsbacklS5ao4nJQSgy1fdm9nz8zt
4t2J7R4ottHEWwdwiR5g++K9g2iNTVAZtAc7FpkjvowFVfbf2qCS+QlraWHOMGAplE6HfSkMItwD
W1tcKsXJq4ZuDw4BsTQMcIV8VBW3aUC3mRKHKEtb08Qry1YzmfVQaDszSy1W/JIL5ikFOWDDkfFJ
5ovbFqHVPW1YTWbcbVjF/AiQmpczdoEcIAhaO3tY+WF3TicSLCVlJ1s8AlzO8KwUT/47Cg6Um2bn
I8rqi8YEJ8ouu+Bs7TtoFCsEUiYLHGzZcUeoAfPEgvCDFi04FMejH5zhNszJw0Tp6BqpZ7H8wP6O
vP0ApWI/YUxbsmeolm+k8tJUEz5ZsloN0Jgwk+TA/KKesoku09DmjE7+kYrWCj+r858u2UeaLJxq
2NSx1r+pvP/XPnC6VmUuM3E88KCq2nrNgyN2u+KPCY22rmNlQck0hHPzv3+I3/O0UU97jpkhvEpM
W8yUx8nESfX0DpO12H70jK/kqPFhNUlXIKkW412ARc4ZVRHUGdfxA/axvfJjGh17fC4rYl+qQ+QH
Ik1IIDtySCfumR/jaQkPCStsgZx/hmjUUOrBv6A8tFXpLhO5kV6KSXCfnOiBR+IKo1f9ykJl68og
zwrRGDpCa3qdDSNz7bb/w4Y2wW8pKimKML2nu3Bclr5rhR2Yx8n+wj3tClu1Sx0323Hdtw9lvp+R
6PfHMtm0P1wKwXqUnxwc9tiSoiLk5Dgjlh7uXIZQZ9UshXg6oaUugCILEsQhBKNM111Bl9WEVyne
UusIDFwVL45Lvd3XspecRIXc8XK5tKKcpx66dJt4zhVWDiZJBvJnDF8YLvNZNWB5GAa6B/cpSpH3
b08owE2iFf24MiJynLsbPp0uRXHd1RGTLs74ag/ceEPOh/YzZUr3ibkCVm1JNU4CPrlaPCi+LWQ1
o/98Phj4qWxHTp3PDH60+MMPzcb2MUi7K5g0MllNoYzEUjJNwVjU4+4PzWn+7dtrCnDVNsiHCii3
BYtzSpeKgX2fdwvwv5+6Jrv8XpiDupYyL127rGYSUjzaQsYuWe+dNFAYmXoaixLcXiE89b5aoTrl
sb0HiGtSihaw5EwqqlmnKT+3B+nRAqi1exPaykHSHOuJxbHjMSMgMlZLEh5iLiacChweBA7eZrZI
V4gbJHAonftiQ2V431crSr1lBryl5icnW42AuiReDvZHMaPS4jw4WLCleVn8fY85dGvpeGvl+UC4
+rfvjUpm5OXbiHPEtW2C7KJPhfrnxwxu210sACOxAkPBBn5b051KRBfiKgZHKfAixhHdzV24cEzj
V+qMbnNQMXUSSboiujkviW9QMt+s5AqemiVTA5h7riC+wRnCU5lYZVMwIaUw0Ru0kOhQZTa3uNjP
j4tdmkIoZooEf5CEWV51rJ6wf+ICkEhCOxKisOKT+JDrRG2B/yS8Zdr/Oogz17ICcOsfD4Anm5Mj
oH0BOPG29vjF15LFkHODPh6OqF4m/AiRwSPhoY5cNkvFVWxz+fWBmD8ep8NXZ2irJ34IkaN+bAcC
1+f61cT4w9EjJbX0PKmRlbzNG6SY6zBMEucwBhlBT12c2/BUq2odfU4CYK/esLdXac6hlnr5U5Fz
zO471Ubvs6FmghYti2XlU+djsCnwFDvIcGuwOkFYzWiMH4N4EAoITd961IApEOr9ihQVT27IDrqM
jCRca0U5Q9pXw8/8V0Vdb/Nk3EwUc6FuA54RLJ9KG4E2Nel9FvioGUGS+6OxZn5ljwRKu8QuKqEZ
6hCJvblM/dMscvNE6BEyK8M68OyDyYCzILzII7UfheFjxUxMi/byVLcKhSO24i3MuVanfXnkSYKE
RWiQiuk3I8RDIcaR+XmOHSdp8kvWl6pTfhDMNbX+3GoZKKzM9HElPjygTNnaT2eqP2PJw4g1+qtP
xrK+9p350bGgOdTby6/kxOqA+dAKJf3zUqOMDUipPKG4DOYKTHBYUXvJ4hptzIvZc6JHj4Pop8f5
GaWyOJTckofY7fS8w5lYLRtobEcUgxYjsdm5tOyuVNPMCSNNU8eXrsY+QE26njffP/kfhh8VAbAM
MKmZNT3JywkznaLnpggj43CRtVKvPuHA/JiroEBiX2bginq7ydnV9EUmz+dgotA2p7AsJTX4leXW
0iY52XZ11TYVbooYdA+moi9EfnFWzVqKeLmzM+9wjqcD+/RLkYuCr5A2XAlUHm1mGhVi/pK95IsI
kavinu+WDUPVST4oIB8neJnioRzjBEWfD7Uou/FVz65cqetGc8t652TJEYXk8jzr1Niw/cd7KxBu
t2/C9TClOraxUr/+jvsw+T5nm8RDonSfSRlD4Yo5Rq1A/PpnMlSERR0FUbTWy4QewV45sQNjIMvT
ZPZuCYLp42rkSXwPyRndtukdnzExErnIPiScmGHjD5/7eDTCigAMaYIMXWx/Qftb/4JsKUgUuoG4
ekbKda+GqYfvylUEmPosd5gLwSaF/idn2WBYC/WRkx3YRVsdGchCg3hg4Tw4AcGiEnvK85wvJLUQ
q/aSHf9Q/yGvVQv9clP23XXwv1Ir715i8w+XtrzypENLAEeZnUecihWXSeeVCaVqHvRySkhfOcoX
dFqnOSTrFgPyRK9WBmigeNV/8kkLIKQBt6wjvCsYY8EOEcSiQz24QDK93a+67D+zLNm3NT8AFRmj
ruG7gbyBGb7GQS0KFfw26CCGkdCnMavcCWc9m24N0+YMGTr9lhZAjmyjLnbMSDV1P3sqjfLTw47F
JBWjPwZhP9frDzjOY3TiMEt1P1AEJQeZ69UkIQbOpGbPUcBdYORaEwGKowlIgJ27nnAoRtfsOUtf
78EXta7L/WaCRBISdA8QrUvKTGcU3CFl/emmL5RlkCrIFBYOaA9kU0gYN91+dLx8fSwtRMK2psnh
jgAxd/qUC2fwXz8FdohIb9fC2S1SYWXFrBRye3qJW/WuxzP3jfNIvoS7Sfwbrv2NAjCHWvfxQzwm
XbEHbcnDDo9QC3gsj2MkH/OmeBhTDCtSd9wpqoFQn31qPT8FV0fRMYyBBCkBQ3TF7GOiX2AEMbTR
VnOTMwQFm3aiasnUMag+nTx3a5j4qsDGYylMeROf4bh0o/Gp3o2CWcOFUCb+9cXNf+otN9HyZQEt
RN4vGU5seorLIxsNAzAeMX1zYRgiqrK5L4JIq7bspE5Y7LsOG0sbCgMG/N5z65EPKCrzFDUuWiT7
O5E+F3l3rTZO1u72gHhy+FtpCTsfqfFd1OvCXU5wGiZbCtotSx9M5tVVZ4hcSyjOa3LPf1qMcRJ9
4+5inlf57VZTZuA+lVyCD7LY5lwaUziWIa3r9l0ru97nzP5fPCu5KeejSzAK0XM4yO+Lb97Itj3l
m79CE0ePuqozoBRbJWtinvC3NZ2zObVpR/JWEW7QQhRjjFH0X9SoD/nUCuHObF+zbxJdYOmqmzcb
9yDTipnp4mlaAJBO2IMt3OxVsJKvdDpX2Flk58MWHTX+L3KyxgPRxt5sRebqUjmYKfDd/pCl9kGj
EhussU9HM0A8xhKuRnKGPuw18CJDlUmNeKQ8jTIdpGG5IxuSONrw7jdc2phoBp2RPNuobBWgLl6i
JJXju8Z4eGg8siTx1XGSIorpKZ4tOPrgqaqbj1t6zN1kLvtTXVI65bxH+n8xozyNFdlyzy9FwkYH
q5xCm7XIA8puI7HjEA4yvCmeMsf0fIUc6TsjD3bQnIncmSH9vcxIehdZiTsypcsGE79iMS+GGSto
B1lH00Ma5sz4TBF4dvUKK7rynmlf9BqVbR505EzSpOMTY99Xa0xzzhJAZYJXyrwCmsqPzED2XioH
ZOMmj4DV6p1HgWQqBQvsJYfBNfsSq7yCOY4SKiXV5d3cVeRnyHygdbyoIbawgPBSQLXbcBhrx+7U
c4KL972lfUTKPmO264+kjuumIORUR+HQaGq7hyyogo0h2sVz+Sppolz6i4rHsUnZpeShVAJhxSnj
iDcsuUZbwt+umUZj4oH/wwnPgRUY8P3ZALFgb//pok1ghkphdEo/UDHoYwAP0yjAPU9FGpWTrm1t
5DkpCyxdXY/wg6WEtN+mqkaGetG9IzaKdocM//QlMQZHyN9yJl8vpsGE0m9H+ErQPUHF5PrBSUz6
HR67lZnHEztinQZ00iRS7OmmXnpk/P8JGVsHPlBlMdUAi6PdSkfHpB5gNj/hwTZP1fqyfVO2nukZ
K2lq5aj3Q5rVZeBOP1z2FxdGaYWHxESQFyTF6qDGGZgQ43EnM3kIgn+IR3tqxx32QQl4yZRT18pQ
l5HESdTPI432gGcdNT9qdAJcRQ81VauuwFWBALxuOx8SjQ2axbf+D9sV8Xs1Y3dHkBBKdTLvEMY1
6JT6PSScXhLYoxh8eSOFBhbXFiIIdVuyOcGHVWHMfvr5e+fuKGuth3YtBy73hDYudONKAXQO8rfU
s72gWyVNCWht9xG7JDdM3m4kYWXCvbButdF2QoeLmZqosbnQid6tXTqcaCcnMXQpmipmZJGMcMOE
rMeTv6j0t85iJXiL/LcFwAP50hYqRb7CetgeUyA18402SeF+tNVOCAksouy9LVVCaahZDhUNrWKn
blevtSRhXB6j0uIqiwGmu7xJSvVEr58uyMFlIKV78PG4VmUx+PB3FMIW7pSHWTJKn/VGCei53Lpq
hgGj561XmSw+4QXMYvhcn1Mm0VwIMrUr40KTVWuCtDRTEzK06h8uvrGN9F4g5y1mMQhmtFGTlohV
cmphzFtomlVTr++/gmQrtlLucTdU6AIVE3ErWahJGrS9K7N7a6g5hn1uE9l+tsJGWCL3yM45iVYd
iEMG3im30oDdnh/NQxken561DnxJSY+yLUxGotb+02ZNecOG/qL+yAAiWDUxbrdOLOzB+k/ZAIN3
FKGGmQFOEh3fYXXHXECZjOukFyvgxe+G4qhkqylAsPmGga2j6ROBiQkzkiUM2+vAOAlxI1DqioY+
nmet54w/Bp3B7rog5bMLuAn80njpmTlP7oIHX/xUiQ6Ftff1CWkx1PGJchwmXB48XN99TP3cgf4H
cRjrQ4suXchq3lDKJAIUti+nWlO6NupJuSkeJ11TRpNr/cvN8FL15IuyvIMYKOSGkeIiNo0DaSGq
1QJ8ZLaeC23WB2OegPup/svE7j/HccQVgVD8MiEos+LluxwqYEKKDRAulIJv0dgLb0r50ox/3y8m
CkPL1qpSpmBMxz8AaMVD1xAyuLFGw3qtCOS16WdBUKzJdQNgwVTf8LE2Ofa2Ipiuh15tESEn1TKA
9tV6KcGe/G1VCIljhiHCAcVDFij9kuhTqhZ/g7SXzjZgykYFow1OMlpU2VDNL1f4kC61zBerCECZ
YghzC+5MEGAHGIgdZw7m7WwjHOnBop6OyQDFEJrZvdL6tydDIn1TB0MQwj26N5geQ8zGJnNnql4S
/+/3hHKIJVG4h6jk10x1Xt/IIBBbGL0ErRuTn2GEAsWo5U/g0/ZrVgZVlDyA/GZQdPBUe0NeeAQs
7hDStg+9y29fzq9zVAwRk8hwizvT6p5kHZQTC5JBcFRbnZZgAq9AXZqPCQ+zosqAT0xBjCr0naMh
6VU4Or0AEAc8oRQJHiJ/zSD12WxnwfzaTtyHzESGU4thU/eE9JdZeB0+B0b5GeHgJxu2qlvp09bV
mj7fkDReIwgx48FpWwXE//5+P3PfHAdiMMh9IowqwrheQi2scx8htvEZWahwkq/xfacXsUknFdBE
UitJobaac3mrLSLie4DQKLnP8wd2tmoH7fvPRsr+Jf/7+phJfgDDo5ujUslYOLqPxAsZm1y75woh
QShs9e5bjwJUbT9Q7yZb60iS6xnWFtfgYfJ41BVYtEg1iiw8D8eEOixk7SP0mWdDGrgjOQep+3Rk
A7fIgD0DXACZrMxIqM1EObogBorzS/rb93/C00lBQHygA2Qt7ngcGt/FyUcEQ/wnJTn+4HOvXr7t
U8e7eizqETTDcBfpWseiV54gSFsSTJMdp4tGrBP9jkaM5u8eVMbWygGzjNNxN2sOJOSJK+DwyTRk
NVFjhxBK4cv9geQlRJJQHm9jIfD+b6HIWHUzPNP16OpZg71Cu5+E06QFUiBX6WgeAhD+RTIUdBIK
jjYyeBshLjVHNPwnIoUZ13mp03tEfOu/s7ryXQYHzfoVyuecVysMTxo8N2ATQKDY5Mzzi/K/fBUM
YUFwh0/pGPFETLnqpJmTeu8plSRn0BlDbgkJ0A7lXwR1ReqfBVKQ6UO0pDfUCbHEeESL8lqR7KJ1
UM2o2GYvtK8hMIFnJQv4HnN1Vwx2SR0FQQ/7qwYEvJ8KqW3MmebTN7Kd1tr7n9aX8sthtXqtK+qN
0+1vRQzQXN78OoZJ3wfmBIdKxUeCR+W8/79a/r8JNFSYhGTelNaHcB+cDd5notqgi7o5j8fFklUM
/w/vfPh8sB0y87sI6jWxWpPwa+NjxszoH99TsLRHGpkpXrUNpe3/vMIFGlbp07PbAlZthtYC+2Sz
sqtkwdURvcn6K3coHAnhq5D2b/AcUH+XPUrbJgOn8W2lgAbDLwR2UFlBnBln8NiridQ9obtSF2u0
r7h/qeqrYuwK7N7Eusvm29LC3Y7Qxmsnr5/L8OIN0lt87D4B/LcZ3vG+u1GsJCOc074A0KgFUNFu
Pl2x90eNw5zq51KFN4Sf4nxkQ1clurWwh30o09MEZGbf+gnEbGHzjWcDyW4Gn14vssljBg2QDMvR
Qgvdi8xYCHANqPPoL5MU5hnFkzpimdBd4cq4f542CFzWCOwG3hoR6mLd4ttHP7dXwFrUhaEitse+
6yz5r3UAe/3XCF7uW7fvvJGrsoVRVZmL0r9nkOobpWzIJDiBtpD17PTQ7vje7zoUyVCBvIuE4J8g
xK5fDKCWfXiXdYLvFVK57D6njLaGKinSG1BfVrFsQ6UNxq0ufJ/25IBFhg/tcLSelgzz64cmfz4T
i6v6DW6AL2+iyJipuQk/5B2jElYG+23YwFmalzLpm4Bufe2J38UsSM1hXVCAq6jnqWR+j8Ii3mas
NsjoLA84pJuNFvxwhZ6HuC6xZ2s9pE0BVeEwCqU8cSis5BxzJYEkeuiMYgQrnvMzGYu1shza5x7k
3fTs2/ZD5fEHbVkdiNO1R/+SXapa6cpPV4M8y2UXwous+b5uuFBqo4qLXtVTYtHyGCUSA9MtDPWD
qKHSFvnQlAiwQj1JAE+M9PCEdTGaeAebnM+Eq63crnPUX4IMKLAKknoFmCMMclsSx5b8NqerLYrO
vltND2YnTKlBDqXQdXvdYEj2Nm32Q/4cApCyXaKiF7KDsidZdqqAwZL2hed2hb4iZJlJELks/4j+
XspbwDL3tAbBsDcKvqm44SiEaqOBuNJWxb+iK0XTU0IocafXmEG6n4VEirJPM0GFSNNV/8pFPY0J
Rug3sWhOK2EaaSKZEzSI5ebG0Sf/N29PU08lMvyeS4/fka5fsARfBcTRiqVjiXKdGCmDuUxVobAW
7St8GIBfkM7Sp2ddxNrAF62dMN2AZ0A9Ua2GjscIfhGFGova1bbpsNizv+t2s2VAgZ1j9GJWhIQL
IKJ+RqWd6dKTOzO5mxCrYKx/Fm8f3wPhhmJJDkRVq2Ai2Pmz+2/hCKZSlzt8J9a+c7PTTefkLft1
temL2cYEcymj6Ht48lfEGiFBV1LWyITM9ZpQBIBOQ57kLw8oprd/ernx1ATZ0B/RVVks8Z8ih5bh
/NAjXW/iGXF3mTPCMfGFCkGC6+vI6UnSHm0F8XglEu3zUqJ00asUZI48kMnpOQBrTjP+urJR0lAF
sG1cNM8gjtTjYzER3Y2+INwaYPRg4h/Lz2427hhxzbFEFztFFVEuB5yhxGUn/1RRsuU6ndZ/rwYw
0xcI9w8N6idPv0Ha3Yz2SAKcw4jXbFcEpKQhOvyqwyx5ffsPpVJZ4W2UQkDO2Qb1lvq1hQGb0DEF
+t3V1tD8cQxNCD1uOvZwbFvA1R190FpwWQ1q7Xv6Jh2csgxdsCN8Km6n7g8Zu9cg2BU9M7lbjirl
Ju76aPJF6WpE1VPjsPKJYKFt6LxBud7f76Ic5BFlWQ5uik2G4R+9fNSzcw3Oo+46Q2o9Hgol0YyE
PVmFRUVnY+1ROmnSKqTvyoSsqXZXh1x3GedDMvw+KI9AD8xAK2QAWxW62FpCFLHIhZtFK90pxAJm
HvR/lLHPTIPn5aaA0UDfKlRUdp+4HDJ24IyGwcUK0e07fx+sJ6x3A5qz907wgREtoAItcEhV/ceN
6ux2Rhk0cjKf0KxDuQ8L+xkvGAzob25KbEhpEqKg0lokoXsUBA8vYpwa67pG/xuDu5CV/s9/xBLh
nF1tIdLpFJYY6nghJkxzXfBMvjf+Z8cp02GsatvwPK9BtfKt48LdJYmvjU+QX+zF1pB8fQs8/4xY
UT8c1H4f4l9z1V8ZQY+CWTjG5S2RFI0itzGIrQv3u9eFx9g9Rf0FwAkBjzgK0hQhTHUU8+QW+ANd
V6KO0V7rEMfzEhtE2SKNdhsGyZ3LUw0StSor5rpPZ+g3ABZ8tvBaemD90y80OCkIGYuS/urHXf8f
+hKi5HcqwOv4cIVvSHlbsuyVk12UyvzJITqUTzeWWhdMXSgX2IxIwQR1XI5mFVtTYtcNVAH3vqQ7
zYRn9ue9Cj/eXYCNj55Ui7maFtZnQt3BO7WsQ1cnWct5Svl7RN8+e//F9uRLNpHfe8FkjfPLTc4Q
IVoIlnaBNUGRu43sgP69EOB2XSGI31/65DZuucHYOACh536mWm7LzmK137Kuzvv8xra9WXJftzI5
LZt2oKJUG984h3zlxACPDGBkmjqP38thaXiR1ov9mr9E6cOdeZTk3gFA67lgGwgH5vU5EhSHuZN/
CPd3YiXDWpPLVlGPFHg/4OP6CgsYMUkrrEIiQOWxTHzVgNjCh9J6NHhcPWBK61A3bXW/mKxUsE0c
7AO0SW3Nr3KZ70xYeDx/uy/3WtDz3ZPfzCLIkU4TsxYKOqmDAR/1nJ53Q3J7lJp9alaNCrQa9nAz
xFUnbRJH7zMNmX08vU+ndO1GuV5QIjhWVD83uH6T33Gfr5gZwT1JMagKCNtXPkmCH1kB46dnqjvr
HYLbRgRYAwcRUOk3/3bPbHSIWcVbuUR+W31RLgINDsaxYhP4XchDx14iFYHzuQ1z4Ti+1BEE7QwJ
UfgDVj6FoJamdFXKLt19YPLo5KV5TpjgvnP9qBD90f5a1TuzFo82psvVFm2PNdhhEmxd1121qhf/
gTN6QIk9TUMsdyh48xsxzdEgvrsJ4ek6wm+k4vZuhwWESpIBYBCA/hlDNSS9wmgMZmTWioob76OV
zoNk1Od9rPz6dWTwmifnLcCfRfu/uXz0xN3jzG7OXQ3qEJkaQK+1t1+d5+L96hdjPO7jwZOeMAyQ
QY56vv0OQstLtHM5KcbCSRCVq7Bu27YVc+wcoIvEUU8yvSA7sG1IYp9lnNGaFLkr9sAlffOHv3Q9
0zCTEVPdXR+feqZYYWHEAZMYstZQrkJiVADEMgm1sCthSHiLwPqMp4utyPPAfDRhrLWzNf6B7CJP
yY83cDk6K2zucFsVc4dmSxM7da8hlvGWFHFeF/LPUtEMMdkOWEmtYAd3DrH2TwNIhltq1p3LW2Ma
mBRDWVvKODEXFTdr7ItsFiyIRRd+MNuazA+SQRkFFaAQYwQJkNl+Z0QHpwEgEKyiSFabxJONPA2q
Vtw1/hVJEPVamWd7Ww38+s0LNc1kK4zhnJFCtgsheegSKsnXcKaGo6Ble9ey223Ch0yWiCYFHnlX
a4YRye+ml0uxWNj1AjDVrUfpk8dQfNZMGqD4E0lKocV/gkkiAU/RhXC3TfERmV4MJez+oaOh13TO
odWKHk9iq7hXyQ3baC8/lTrDJRFK2GLN3R7yBz9115FKJ30xTESxRMZIFHuZm+YhtkHVutQCozhz
5p3S+wl2+3PFOXkaj/4XaGFveDKiPR2qxzyXLw2lBaNbrTQaNeRGt8G4WHymd5a/3m2Vqu1S2W1T
Zww/twsQt3EKZ8Z33zO0W4ySGYrn41Qa0HDJlOtYd3AMQXxB165oND4c2MjcxnQlqkH5zz46f31u
fJMHDv/b5OgcjCWQDiLV1fBHFtJEmqxnE3BY0BbCIBQGoYUHar88oPhataiSGRER8ypBvdF5y4fP
BtxgjiFUeli3ef6KwV3zgiVWJoZvYCY5zPwsKqNaSOqK6S7GWmH6tbMtYB5/hw9DzqfBYtVdwCKN
Y0aQqFhQF5ePbnsERv5epbSvCJHpAQMEUV2ftzPLNPlKDAKMjJqWawsDsRYYLUZ+kpha1HS4UGdz
5c6SUSJgjgiz6pZlvPju1pXRx7Cwo4ggyTTWLxxSJ7XcWvlH+CVLOuinNNBLalB5Hle03nigOgqq
8/gIrjtbGFEvN1rkjgPC/m2EcgqvLGWYtVXxLaeUam5erPY9Xpo1lnJI1Vcw6TDWMqqiz/pwxVz8
zOK2ZPz4O5x+H/ygK9DDLIfBQRdFPQlcK9JucVt1Q4/rlojgBFTxxQMqXIxKIzlpy4dVlhBpPrG2
GfV2pCV5/SdYgzS5JVKCon1h6VkaXIE7CIf+eorSMBq0BoY/QEzsj6kJdxeZ489wa1elEyq7jJEC
wtYRDUIHnUU2cc0BIZENHDZ8Ospeqr7n2qEvYJzBeynl8ae/H5i394E1K8Ourlj0z33iF5Vs6Fyb
+eLFp6Mux5gympb1uqXIqaZLjKV68cPskMXaWMIbNpuE54COlEcKTDIBJ3v24cJU+jrhMAeuqqfX
giCML9XOlGST4lf3jN6WZUNjr2vgA1BY0eY2WDV4JCbjxvilzlkXj+nqP8UzIqCAeU1pSdMkgB/U
7qT/LWjI3m2OJKSX4oe7oHc0ld91T2+jmMBfhgeCgbBQCYyz6vjecSWcwjJ4jJmbUi0yyJK6gbtS
sr9LfVguCalozuCWG5mhItpT9uJv26yL1fXGkWF4VwdjE0l2TuDg+umMLXnxbz8/F8XeyOdhSKiP
+cPXIanRWhQ/FTlf3r3k3ZiZ+zsMXdjENXHqqWaA76LYia+zQ/bA2IxyimLGrOIxr78cD2hdPlWz
lxZ/qOXHWsyIYicJKKlKTKOo7UMSnlkT+QASpTgnq84HmBs2jDI07DQBUr0Y5owbiplD92G52lZb
1fNu/irbVyyI1ENQETrBn9azQETwDiTj4Flu1bNKzfwwIsp5MMwjMKyjZ6CDAzVciaMVkHuZ5BHT
WDkkvQmMQdjC8arkENr/ZiOxH43gay9cdCpUKVboVYjnFR2vQjICXidpQNMaZYL3xCjeTSox0yaQ
Aqb+1yn5WmyQu6U/+qf4MH4DT0pmPde+FtH5+eglTSby6urpGlmnrn+9em4Wq6FvjWkPYlOiiD6/
C+WRmiUDWoteM1dbMYzkt/LUGvA/G5mgzgAbJYHhhDWQ0zX6sBIbtGwoyeEr39ByqLqQU2QBMbMq
3B93GgwbLLP4BAEtm7cL+xju9EPYUsvvoc9H80voTAPCC2fSw6KeNeOEIKCUwujs3orAtX6HJUc0
d5kKXOli4Ui1MU7eCKxjRaSYvZvipQ8FL5rL8BB4BqkMfTWU9dXs0NgdlIbnrG9QhgYIw/KjnXc1
rDLVLrn22awr0CGH5TuY+9lafx7RXhw8y0cbjsk8FyuO9lORRjcaJ5uJojzKE/kUNclje+ciO/96
+4ao8eHAKyk8MHAzh8RZ9nUnwSKkO29zqtCUhmqtqgsWskLngKH7aM0mdM4CnohfD4A20zQ8W3fR
IeUZARsymn5aIKwT9gW/Td5WaisvuRZR1msvZMFJuwWoUrA70gzgCwPFVmZprEH5/+2OZv8Qp/cA
OZbvfH359NDVSumHIMijSPsdcwvdFmSnBQSkrBizLaVGyN1pMqJFY980LRvUu4SPNPxWUHi6Sxlx
+EvXTTM17HSGlD9qXa1bzG01FIvrFJxb0hD1TPyUzL6tV+1nfWG+NPoFIkvvvX/PXU4C6UY2Ob5l
hv3+nhqm1EVk2q1Xzyv/+GVTk7WWdDKYfzvhE7o7v5L18hbCYg1AgvesiSbAZt9NMShShjcGq33J
QBELiBJlxjj6CttcXhRvJ/VHO0m+xjZihnYuSt0pPbuTYAdVfz8nIpoLyoY8qYdvcjRBT2t56gM4
IWQsQbIbjDF8pA5f/6P8DnxLTcnJTam2wsqBW4p7wjGtIedUqUlJmN2qsFGGrBwFBYfoDRDSCMAv
W9eQAqQYvACXjJSM3iYOE3GKJR+fTAuMGvlttwg0ixVuZVOO7Zr/XiX0mgKEtDDGqdsDK0xiK1Xt
6y6Od9Zxx9VVWXH2RWasT8iFIwKQP9l/KelMFvbl0zmTMHGjnfOW1p7xdsoVgeO6Cd0tJqOjMstO
Q34/pSUtnqoYZIdOpb48homWYuYoi3XbPO0Gwxwx8MT6rn9oa5wMPtBc4RIii3f2GwaYsaPytmL8
TibJQe+B+uynSWvWekqswGGc9gOAwR9Pas3+o4afTpTLBJXt09B6TLsZDLZoDahE+nBp20YerE/e
JP43/FgKvz+bcUOk7oB8b2XdP1oJIZWoiUe85uQhr8tzMAs1HkCBwtllREdFTnVLhaqTlcx/azFd
ZZ/XdvB5q0OPq/3O6nj7vCuf/P9cYz49n/LjKWpE0809VrXu6T2qZXJicErxevR0Uge+gWc3LAjO
t0lB3GzfLwcGD2FryWhRdf9rfzW56NbJyfQxIskdR/okNn6qHwMC3bf6tKbqq+qqVMddzUf5TbEf
BPpm39SmztOaAUDNZfWv7NRNUL/2MLnyR7b57M0KtN4tFbzhAfs6k0d9tGM/7FjtEygs/DeuZ4nv
s+WCpJXjprj2OGNjfUbNP8Pj9Vmojl97gb4FcZachk4dSvZw/x6pmNTf9qSePhAShJnkwb3DxqFX
vCFuot944I/wP3Hph2Q/ie5n9cZb6i3mnuCufJDNex6x6LfF2HD9vPTx11RPY9DKHPW+JnjKaf01
l8hgcYA7MPCwmY++EX1FsEe7NoSOG+U7bMo+XCTN4c7H0HueAzjjufKODcNOYp5NviIKVL5ALM8w
+zC1cnEfroUWVbr8ljFlrIzHD/t5PJn6IK30K9ymPCevbwe+DYct+m1RZCrJezIyaS74n7ldDU9o
mtj2kfWOgDz9hGp8l8iCcQm9gZu3glb5Z/NJpcI5HzSKXpOfIAh44f8dIN4AO3dkhzQcD1K92g+N
7I8eULvD3knyjHYvQr/wL4VqvhP6Q4ds5BgwAofToLZ+daL2vhu9stVTUZ0TzY+VdfQ29leVz61v
MMvS3TxvQTTpL7vpnCK7cd40dnHCUavAzk+OUXpFxTdeIBP3ZgE8m4UMBVgic79Ve45Rdu098DII
oRz4GU+Mgpl9EDaqvS0LvBe8q5Ki9ZB3ub63yqycM7jLmb+K8LuiMS1TLqqoetqfW+db9OHPTKs7
U8/vIZ6BeWDi6c1CAkvpxvxfKXwwBN+Dgth7lsOwZU3x93A1bl4SkIBs3+kazIF/BWMdV84Hm4EB
YHeDMlxq0HEWyXDwATastZ6iZnM7pOvcuyztdsi7iCa1RnwuNJ+3UdbsfP2Zx6PSdkHC/cVz960A
N3hT5cW4Jx7bBgdID+FWyXPnwpdLrRU2uFHxLWxwB7X7qZST3QRbk1roYecIrXi7ZRpwDpV0rJ21
RSEIGLoAv7StR5PymLl79XFrbJX5p3DgTejowdERklStTs4QZcnvOYdsT8rMi5C0td+o1qMNi02g
OvapAnHdzybRdzHh5lQy880o2O0J1SjHSNDQIuwJOICbqEDY2RGoV9pqLHvkWgxXQ/Pf3/BWrOY/
x0k2BwBuyXlDyiPLxi6zNku6zUyItxp68VzuIn0sD+yEQD6WaVFLCdBadws0aXfF1++ZcXTj4Joi
1ywlhwZi+bwCTVsz+vSlYSdOWMnnemC0JAt4USX5RojFT3KDL/hpzvdSXqOVSfgv18+FfhW/EbXP
2oQbUpsvt25So/BYN5vw+CwpkYehk1PKEKANZZQZtIf+wGrquu0Ko4/iomjK3Bn0fyHo5z2yh6g2
6HkeOpOQXLTZguUm3BP+KHth37EoIduhbrOP7vGrJk3pcTZYv3ZxqTQrJWCiSEpzVv5cQgNYNssq
7PgEzc0CiLH+fSeswzUhxCUK+bL7dDWGZniiaUZP0ZtORHTUpJwAe+rtUDF02+Eq7nO8+ymjXUbS
NLrT6lcrumSD4qcafv1GdYWOv6WQNvqgfXdM8aHDuktdXmbJUsGIOZHfB08fZKkXQmN1fhKNTADp
NFkljJAfWLNd/YowhAH811MXRKa1QhLScm5X2VK6aoMiTXLF5O3nZlGYkMEuRc9TrFJGgHiN1O7j
6g8lUFiH0lYMYTQPI/1KzddpandxeEex5meUihhODohtEicZq9rZxSPfyaejq7Nw230ZZfpYMD0Q
u7NQ7blj18I86nrmH18evZ69alWaLMTbhKop2qe93MLBUrH/QqS5kRJcnUkDEhT7pkN+WRRm3Xxr
2TS3l8Bvp77R86uP8V4MOvKohjzD46ok+clqkD0aesmr7TII6DGnwoQihZqllSO5rUIF572qK281
Hzxti5NZogU+REbF8zWW6bTwmY2wTkmEoUt4YUnv5xN/7grvlmsoOSU4FNNebvTLDUgBU9PDX108
uq+aieAmY+BNmvsZa8DjnAML8fcIEno8WFfoEq0SISRxw+TXfcnkgNAm3MMWL+Fk7p8nqE+2ubsh
f3xOVUrZGnD/uMT0D2JCzDE96VaZfmWuvFPld52AZUDjRitgio3fLUeiBNsn1aK+o35c6QM9tuKV
j9lFmqPzq+CVR2Jfo4JnqFdNbyYuohs3sEx3moRhE8VMJtsuKETd/XWXYwZvXpGkiJr/du0ErUSF
E68T+tGgQGDA0cUO1ImE39+EMpPMcV+Wd1zBXdxsx4HrzV881yHTkZ6JOL3M8trU3ji5wP3SMQd6
k53UUu8pQPtcONLhc4/7rPQFy9o5fsxsBbkSCbRu18Hq1Sdqt26DlKM7H+oCOcx2Ezi3PwYoKz2x
JS5DOaCXIcEQpNlDda1A7i3GT+wGGyiQjiCKgq7/xsE9WwBVJrx74Sh3bQ3KYCRxmAWu7iqM9UV0
OVYzqs3IO0+2v+c1byrcyvZAILCWQFoTRN7L8WVRhRY/V32rKv5YJBiWmEfUIA/QdwR3siI6Nc1b
iitS57Kz7z52IHJz/pScbP/16WSa2HUMzS9B/a5rkFPXnNwPWSC1L2exTBMLjsruLe70UZr1XoV/
01PBljoj8yaMwrYOJ7v81H2R+eP8KKP1i1ZUweqUPiJEa1M0aTEQJgcVlIrutVszm4Mwcmaxhyly
Y6Z4hjyRUtKpvqw+OoBPnekZwiTdVTY2AgSVrlX5YAQ9dayXollWW35+Bu/ugOkBPiTg6nSh/Bij
2oMQC7//oiaNi9l5M7Vf2QGpLyVeC6shHjmCzt3OF7/pqjc0g/kL1znaG9wQFVtziIHGWtqCKhy1
JZTBPSYNxteUsyYY6xZcB2ajcJe+RG4oWiRtDDIuIxeiUZHip7kSUWc4OVVLQJ/GVxrIkWVmqNzz
kKd+1QGcZcxpVDqy7qJ6VMq2sg09C0c0b0JrA8oPRbLrFlVKd5lciHPf2ZGvOQ6d67/E9w+U0vVq
iq2kzIFOQiS0Gw5WvdrvuK6Dor0xXK6+Rmyl0tWtg98pZTAnnzrQWvY9q54SQhHK35dIVOjpqO4j
20ycG/iCdfrlIvetjvcKLe23dziZQ8S8M/ZBM+MT5Oucz21Gemnp8pg4VdlT7p1M8yVKzAyjK6Gq
DIUMRoev4XG+xopNfU0h1I4/70nVhsaQ/PFyzQJS6HkptC3CgwfJpAbibeBExlkrQw0iA88xqqht
2Gzl1sfaS0L1/fMCxu0eK2QozHQ2Y/aWE8FT98m+MJnJrCuzlqg5iF0xYmeB/N5yyCJz0Syi3cLV
6qdx5xpyP5KXf+r1OGXK36+cRge0+fRY9pyIQz6rDJokqHIqYYTLmHP8w8HDqDOU08EpffOFu1CD
j5sAsTPf7xgOnb4W5uNE754hvv1R23qATXgkzJ+vCwqXV9YMXfLkoZgq5YNGrh7M3Mg3gy839mdX
SYNbMAdm8ZK6gw5HuQ97m2IzDimHs2cPPHAg9KVYF7GnALcV2yUMUlhunFvsnsev6pMhY4uj1vJR
tg9/PG9kHnwVwQIvDlR2TRdiQe/RXHzWBkgfnuwrK/jpao3/phOjPfc68smf6T/CXD3w9it9plx3
xtjdzfBn4C3hWFvNF1h/Nn8RLS7kh7sC2K20eT+MxuuUg5Kh8UR9yHJm05Om7d8OkD+CvY7MwiCn
6+qp4sEpG44boc4PknFTnItUKwRBORO3UlgZyrZe8twIc31mrXpRTW1J5mLMc3x9qmgJJHVcAUYQ
FopXmsnn/GWm7Hxv+q6oj2h2ysiMvqOzhXnLk02suKV9hAqjzwGm+WJnoLPTkwtVfuF6mj6wWnye
IHdrfxWWoAjBDrv+6TcDD677Z8fgvwXyTMHd+STV0Vsk2FZo34/f+VUUDmJ+X8wiDNsbfwhYD1rU
OU6E+t0OryRcbduPWHveBtzSFfahWURDOanwqxaUhIVUJ5fvmEb99g5s7QmHOue/nOFhXaanRqYB
6+5NoVZ4VMXQQZSGkCwVB4I1rzQGB8GicTs4jSFMmU3FR9yXtsd4AXxjhN771wHR0oZOqbAjYfS1
o0Z4lE+oltuDKO8/BP/32xs6s6WQcOANLOv375Pm4EyAPVf5CEnRev1JgomPUiR846BAx6T9tBwE
YzGIUvbWpDscWzSe8WS0RG4ZAWc2C7oo7LODoiikNnrToDGfkpfH79dCunsdCwPjAL19eVVDUVxl
Blrq1dc8rz2I1Tt/Hb2/x2NjO//RMCwDpDuCOoO9yGR2XSFQgJR0UGqiTAzJ08berdUgEiiSEghq
QMiGuMj/vD3c6JGGGi2sqYiPaOGod84gBM27jueIS1PkwQXxwXiluVV78wz0ZUJ27Y6hMQwmtC6/
PfiDJRiLz0RqGgkhBpTAPxVNFwtKH8W16VrnSNq7y8g2FZXI0Mct2gfW1zQm8plHAlfgnFEtSPpP
vlf0lGUBM722qXZx4I6XTR8w+qjRp5jbIywACA7dvpPQ4zCA8aPCn3fuP2/s6NZxBxhPA8NfHznn
8V9/rz7k00/66EJep+/deBzrKagNX+ekuFw8b9f8XKbNz7rPY1gmbOsRHgNhyQBlNfhr2uX2iBmJ
wkUL5fpnZd3nyyMEx+PT5eZTGgblet55FwCZ9Rou4aPb2jOkOd8vHGIl1lG6SUW+/xj9S7u0QV/5
7VgVz/8PbcI9jCA3MLMnPo5Y+ynh994dTQhPo+o6zkOEOplXKJl5iZekUKx2q+Q5gI0BEZSzZcmX
49+Q/D6yVWdNeG2bnjMPdcmG8p5CwRs1QK32QjpIYjWkTGQ+TCCe2ETy22ZIOExToibRE8A3VNRw
YhjMpVxdYl+EJicAXN/ZFmvb1LVRSK2jqAFRNTtg5pX9qBu2rBYqo6xup6MFARkWV9vD82ooynhM
Tc0fGaQCN2g1o24Z/yduizwmeAJQVtYJrmYgr0qxDL541XtlPAs0hVtbbSpGFmnRuSiPvz6WaS0u
y4LJS6mPAIt41q1QFveC2xk55cj3Xoc6CozrFSeIg0wlBBTu2mujK2b9IDWgb8fgFJnMcZApOQ0m
3qvp4+GTNYsOQTLo2vhCmOP8yl9kwZT1JJvO1xerzi3H69i9CsajFl7ah6d3fRL6x2eJ6wNS6oBu
tSvCJdG7z/xugkcwUCBWOZ8XnHdRCsVkTRD9jENHpPzmY8UgontW3sG0nLQh6hViroyV7zTfqcUN
147BNeeHyYPqQxPfmKmz43OOBI+Dmm5bzwY0ydWszYPIt4ANibYNhgCLQ40uM7wBtAyfs6Jr5CKs
9pQyns557zPFS4l5NOJyqz2WyHLXwobpQwVSDTOclGLO754ChH3ssdC4IriOTZpBP7iLnXBrevuB
7EoG2UbrDuEzrrRDeNuCi46VnaN1i9jjXBmQfrDWiIONmp+wy8LoMJMImBVLJSqzYAKkkCHvRRP1
s7gyK62833gvIER8n0fRawmZHOLXBue5+VHzxNVl3Yf9nYBxjiHmOYzhLsUt1x73OAEXrrplWl08
FVh+8IMh/69bnpl7JgU+9j6K1iRM1QrSV6UFqyJW0/Ob7sXh246lzGrU5BRa7GsRsOqTfg2eFi4U
drua+ELsc5APu05i9wQ5+Mo04JRjsMV/tlUoYeBkI1E7hwb9/rXrD2gZCL3Kq8GVjd5At/Jc22MU
viUROJMg3U+3iOUsx7DJDKLcBxHpb+OtuE7LHL7i0vKKxIRquwTp2suaTTSL9hYqPChZL0ncJEJK
S586RTxhvH9eex8+frgUSXLIzt+e6kyNQp5Yop0pZd3R6v3kr0ChvQR1tvMGLUYoNUvA045DmuMu
DNGeE8+mGJmyBag8SB7UAHxtJ97R4Um0ZqIcjR9hcttRdSjAu+FtQYJvIK/2OlnfhYZntOVrHD74
qx7DyDbKTBhx/0GkhMl84MNGgltTLd8/bY49+6hKg52eCCiFokXdjsRfL8+IkNxneNL1bslv0j3P
9nS+jzUn8FgQpkmZI2lwQLM/f0Siik7IUDBHNAzk+f3rhocLHFM8crDasQmQ70RHH2DMAQJnxv1O
jWK1nhRHiQP8O19SP3/j+F5CUHzuwEuAXq0UQXQnSIKvfu75i5G6I+5S9qQ6uZyBd8Ad9LVzvqi6
dwWw0cZhpBkym8n9oYNpxCkfP/0plgKFD/wMvWxoKYbfoeFh69VvC13bgJOWEVAC1y3SUWiPmjQ1
kn1HzKpIUEe4EXT9dHOz+QaIRNEHG3PA02uFxhoKfNJhHGKqj5W1xNRnZ4vfucCThcz79OCbgHOw
dz+Zu+Ds42OIVskA0Ww+hYY81BGIe0Tp2qSuC9w5Lc7dIeSg4367oNph0hkW5KXvk42dcpihIYhs
C0iFxDmsxUsURmKF0LkIMTal8nLyAf4EvT6+BWcUouQBrNZG1rpi4GChBG2TIwBN9pirJR3XTlIg
7FrWNvatdtIvuQLyNoqwkJhJLLka8lHnjgzeEr5O64yOyg4E+InqAv0r7UNhhuyyk2tW5DidCllh
DJWpQAECtri48Fxr/9rMbJ71NyApkkCdGhE2HK4xJiDyQCuCSZ5wGj2lWf29jNMWkVquk0RaXh65
iHJAK+VjD8erUTInU0OFCCzLC5iLf2odMLqp1abqwmjFobns5SLSFz7FnMvcR6/itoXvjb/Q1VuR
b6WmKTLyV2hIXm9qbkKTDcgifP5EKfCNlsN+go5LgYaWTzIQYe8W+bl3sK00+5GoVu8wpWDx/pZP
Wsw4J1YnUMOwaHsM3NXxVDA9KTY2Ac9Q1l8Bt7FzQaxuYVIxbz7KBR51WvYah9sv+d6SLpZXsO4t
EVPIXxpoKi/DiQOnQdWODnvMFKBA81NnMMbNtaXg6qEpkl1bIrbvp2/ZahVHFUQUx5ogeOxHTbWx
JAcqQgzNHfM9OPLjQZJOl6bYIg3/K7R7XoSQUOZw4HVhz+1FDN3f7KXyRVAnafebwN0n62ZBqyrc
FSCv/1HLF2qFExrCC2BYu0jRc0jgV3EevinDDwDF11NZANyYXv/8LXfR9qvUzvvsuHQVngufYK8y
z413fezL5+my0EHdWCjORXKyQuAkqAzCCzDbKrV1pbjoPg5QwpznLn4gUlTXXBLM+M4bq+y2pR8M
OFtWNsdYJrnc2iPrIMOKOlA5W0NoXfjBO2Yzda0h8e/VFWoJ26SZxnaTSyjHl4JEBJeLQGDV8K0W
JqndpRe0YxkzKBpWCKFMM1mAT8LCMd/MOL3Q1KZeKQHjyGuha5VzyndjLZfqxQUPsLauXR/LZE/k
vjpPmY5I1MmomS2gAT8YGCjK7IBVQD2MH1PHANyO4RlkxIP3FqDeQ2uEud/mCUpuxXCYIwdU0yal
ThZ9h61Q16dxxFsk8al33BH1CP4+gDVlhT2CqUgjg13cKaIO5l0goBBXNM+hbJuZUoUETZzl5nP0
2rAii8eNEZIht8m984FUj7aELIZJcsjgPeVS/SGjh4hZLumvxazdRQrW1YghDlFcTA8j/2FtMLN9
D2kYXN+XrMBf0QUKlnbTQEsRo3BBFGLAnCe1wyfjtmKaKmXLQI8fWBu5AgMAugsJ3xxzTCnSIr/E
2qcQSfaz612x1HfvmAzifymXdbxGVn22HSZGP9Cv26yfUZAV29qcvrNeQUfK04w6rCvYWnKMUOaY
EzymlMqHd63YIks/qUvSdud9UYyRK1neIzVEXsnzc2tpY5hzbGWSmd7PJ5d2Z/LnLNIxVmGbogNo
Bht+Wr97qkYPcFnllieovwTDxFjz7igmjGYKKcitl7Iw22C2u6bcbMcsGBzmep9/PZqJxuKUwJRD
3WeCYCmZ6+u65hMz9Ifg/g+EKFbdqbyk0XS/4i+m9hg7XQYB2hc703uES988p41tVZm6qwqy76kg
YANwiwhHu0m04+suOsDCP8lM1gqnTrigJpDsjS65pu6ED8OcIiMrPiqTd9Z1n2fVOIMtknZXdMIh
iz2a6xaFi887pcAO1TUihp7Q4TEd70jD0m2OlcwIdc+4gWWl2AFfKF6LytiEqmwFxJDeMdJmm7kC
c6U9VyckKOtoUngNuLxypfNs2/GH7zXsEsJA5Ni+qBGVQRyJxs1M4ZWh7UX5rMlEL8Fr3qlDH8HQ
bnA77IOz89J5LEMHF8wjGq8Bdj/AjdQeGI8x9K+dq7c19PhNnoH1Vfpwk8wxF06QNtQ70YTrzNOg
PyVejBLT/L0L3vbVCtGr6iwsP5v08azkJQMCrWfzf55BobW2gZa3PYiMS9nyV0X0Dbz/6hFhtpKQ
ccqxkK0WfkSXQZO6VfrmoFcM6ifV0g4HEX9nwK4lVHtHjc6EZ3YaiL0TBMbfMMGDhGwHXbBlOiK3
PWDiZAL+z5wQWw58ZxaqodmhcqO5rtMHFitCkwbib2RJxowxTpP7OP8+ulNNYu86X+CFerQSO9BP
jOMgRawyV4SIUEWabiLh7PSG9BmNosQpm//NHoNx4jipDmHkazw4y0i2nS8WI7jNqDtrv0fYRSyT
MyeDYM2mwcRFFSINndMnj4/J3L6/sTiAVzZ9jQA3nxJfFSGzv/BJMDQEePwDP9rhEiPCcVpDzMVm
G8fsT1/5ZpvAvfZVdzfeqjvfSelSPtDPKwadiRAxpcIGa50z9r4rrqPgdJpGir5Pv+p5mrVDRCSf
W1Bj+uqm2ez4xUuzN2t86IXdDw4ZM1WCuhuq0YTc1Cgp2gawoWzm58tW+a7AB6xsXPgGUHHaT7+H
pAV7PXsh4pOs+nWLI2J/hFfQYvYXEf5BPwMUjdxvBfXzTQwcngniq80VaEdd5iw8GvQZVDaFy+/K
z2RRKzVqrTns/gvdz/BIPyZpjpAIf3JSXrVvXJibqh54w5NbUlevV3CogOBfyRKyb/LRa0D+Ts+/
uFHiyCnT3fk8Te6qqbEllraid/+PbDo4GBUb0xX6DtxK96ThDiNY9SCdypygUb1WH/ZieC1pIUah
+kq7uWTySPvKmIjY4bdpr0Lwo/VeIgaqmWq5PF4gWxrKEL/PKk20sraHaUlDyre0rBRKqdmHzPV3
YRsVkU8ZwMi7ya3XGhw3kn/CTGikvPpsZrb7twbludTUuLl2sfs1FoXfW0kcnZJdinlHF3JymVja
cGfi6i2xnBFJRNBTfv2J35NCZbdJKnCeFMZjpeOTofSJikynPxS4HT5natiKKTTabe+jEjLmZrle
L9cI2IItHHFsa8RRByRp/3h3k6b78C9U/KFkC6pSJGxsTuCX2ZwVe+bisBHW2Up79xOnS5YZFuq3
XVN6rJvzULRmcBkJrWa5Q9nqMSu43r9fdfFepqG/SvoJi6RZONTiNmCpX9c9DiU2BtVCbLVpBqQe
i7GcU5HVmMFlJsc7VurB7NqL6LvZgnTRjfQqew6oUnx+Lk1tCNmsNe6AvKUljOWpThWCU9pTXuux
DsKbPCFFMDCcG+8DNpm5+bbh45l6ej/ULoziP/2LQK4GZjtB+ZD41q4nmZ8dfIQvZpyA3P+Fd6/8
qDfnzEUsRQQ+W4AqLGvgEMIfs/Y4tHxs5/oXLSIVjB32YXNz/5HtZDUPaqZJdbYBJfuHDMhqkcYg
Aslou+FyOazEKic22wZklWKMuHP9XedfJv2hwsJqwu3IpIUeiNgoE8XBiXorMzBjMkRp2N4ySLu2
wdar+GH/4C4hNp8+PcYKYmd06WCqdTzfvtOnFjxMWyTllWSPk7jJq9uMh4sVpEgWWRNpAzuBNubQ
+CEC+UID4WTOmVa3fp8VVmgjM8HO/u2pkx2sf/OOa8DZuPJtxokSlt1PHg7beLl/2zJbrZYBf0bw
R17OyH6Hp3Rk/NGh/l1SX5y7Dy+PTioUsr0QWcAR/TmGEYRE/ul3XDRzcm4XL+E2xT92Nlk/9TkO
pmy/zGHdVCzxmrbMgvAbVRur5Loz6hlpcIl3QFx8Dj8bmyM3N9GjVtwDFMGSUXkAhmYF1c/skdCI
sM5B6nPC2+AGM2k3ptB9aATg4ejV2XQ/jkaSNrOkPSunQxfa20X8H/HuZHM3mUPU1x2wwz6JT2Cm
GnL0wlYbOyaVg+tg16jxqROvSJjD4bNpmjQK2x7DADuX4K6XweoNz1fClErciJYEd5dWCItjGY9E
/zq47CIZFtZ0KmyJtDyS5ojxIIupCI8RH1Vf85kb1ciDjjovEbO8ydMYs6+wpChfHWZd4zgx3g1t
mYXXUl+6qlmZDiCKvNk7UEI3h9Hsy2Mi7KvH5rGNikdDPVOBr27/PPxbxN4WSZZJomSG9phSXK/z
d3EhxiJRH2V6GMPsjJFsQQE7cYbzofRUdxr5AmXACqrsYjIMbjUP7WPHD15cvbQLokWGQx8dSkLI
usK+JZCtkCBo0vXRBoTvg+CmJVwDI1qrhmI/aoqgsgc1W3tDckU9EyZ6T1j2210hMDNJMt/3znoC
fFotTf0A9KnlZRQBax6wZe40+Xf3/lVTrb23JztB9OinZINg6ThnEY4QJxsUn3kqrXank5py+o5I
7OaCfwpixHDKt1B2pgs4Ll65srGKccTkB11ZdjVj4QcEFY/YlebJWhPyakaoQReNSEbFWbLsOkHe
awJYDtJXkbQ8ehOzFCcv/r6yVpaxr/WwX+6ZhlUuP6H1x+d4AxqQmIW+c0Dhw+/wu5iSFQGf1gs/
jpRZ9p7TgOFzvAQF0ZqP2tZNGKyE7JhkEMAMd9FYYn9+dSC2NtFHAY78iY/SAl5EhVyl+0OGcSpy
sEqm2MsbQB0NfCLI+3bzVzPyixedVrsVIvYD0Ggio05mj4DYizIECKSP42MujWXPKKLCJ1ZvnBn6
Pe/tCQb4djTcZ7ba2VKmwbYnmHwhgpRspTgoqFj0M4SKJQG0U7gGQGMMoVRc1t2N3bbEU7pyvBAB
WXWiMlBJq85fa2+cKJVnJejUGAHOmETvyqhXm/dk4TX5Yg7c0FDh2r55eQ4ggfEt2cCfKFgKh9I3
qZyBNz/8PT9fFWJgVCHW0nAtSjhvpkGpdIQFiWxnND/l2370rCKPKbo651Ih17wcqCOGCP1lyiid
+O0o2c+3lFrKCOgaF83WT9cncpbi3Gn+BjLSaQLxnEsD2ZIbnu00fO2mekqMKqudggtO6A3vwjSs
Xrlx9asRHsS7yzgkcpJ1HAfAl5K3/gaSEfk/siXNcMXu6IsF3kNGBKFboG8zSOpO6gSeXk7VvFkf
rfMzwx6OQUtgY/gJSIKFgpINT1E/QNfd4JNLuudtRWGwXzXI2K18XQV0iifxXZxYSbJURDvKIR+5
BPQYiVqkfX44NaBkYC9xDy9zv4zJIcm8XYS4I7wC+nxOtRz8QjEktrhLTAD6JTSQVCZj/9VxbOB5
t0yHzttfpcdUkPxmV4d+JJUr7aAi+VCjt459YOQOpUqckJHmKImxwb5arN1wqZ60+C6lZIFE9/s3
X81O6Ns9zctg30Ci23p5lsc9fTT4TU1j3SscBrKPp5ptMNnLfVJSFQSTGuO9hqUXvS9AK/82gBqd
IzSnlobF8yyByc/LGB0Mpi2K87S86amtjVJDx1O/1F8b5slaVaY1nZg++iWhPhP58+T4rNLr6y2t
6Sgl5sRZVRt46CdwhZleyGaAWFB2A/OnrgwEes0SN3yMqzU4ql7I1UXWNIhud/71k3L5SeZd3QRq
6rKySrghWO8VEkwb+s8b6L+A425+MsFvc2Ly3GpKuo+TLRk4zinXhqjJpluxbpa8vPYoHXQb3mJH
Pg/CV0sXV+r1mzvYK3Pa5RrnBRxs38t7HkvPh8jidXNGrUAgqyihkn4QdN7VHpUr2Mb543rWvBk3
vx0Nt4rT7+ri0gndh0TzhqM6sAhpshsQ0RaQSosYOlAFWgcXgxxGuLF3riheUwcUqkvMJvEXMXse
t7NUFGWxDR+F0B1ghnW3U0mHufXRJxye0MIEsCl02w8kaqrmB+piDC6L6cd6XnRg+lXOAkty45rP
jDB+3iqpSnHbmaDQhs556/dGN0DfejhOXKraLiujMDCnsiqsUhcHRTVV4bkN3o94db8n+C63DsDz
wUfBDsmepAIdIpZJmvkKnuuWXUSvV05s6A1yLy7S8yptr3z8ZW2j2Zo6daS2VuSxsS6Z726ppL+S
I6d2G1FGcmwoI1VLbRiVTpmwKcaZ4bv93Ak03+zq6WuRvwmo1ug/0+i+U8gsUub7Kgda4v/JAbOC
XRoxRqcTdrhlz+mFmiR3rJkw5N2G7NveXQNRe/sAGKNcGEMR1NkbE9S9ibgQOOq4xt0mij3zWRuu
qA/pJvWmS9cjzI7AC9+gmpYK1xP+lcEQcLPGtt21eN3oBSFj1dIrzxjgDMrA5jJHm5i8SJfFPDgP
wTimZG0mMCNvoLtqBMfzfcesodZS5uCxA6lkxZdhwWb4IqtRHiRXX1w2/g4UQbneLneHognKQOGf
1QwzmAUHZoxBFLuBgVpgYIhfUW9aN7Z0kEcbxLI/97+wFmTgj6BiGpSI2e0zxSNuWaRa7vcr0aJA
Gkd13bTJy0XuHu2+BPK8Z83dHlfqaYhQ/gXG7j8QbxlaYaEmbPdU+aMtLkYpFTW6hABFDVAXPiV7
c90159RuEjuWRycKg0Wbi0LrrrGgMO0Rzs1rfBZndbXk8HGhul+NibpcYy7gLW/zx6C5bck1NOSz
29P/eG6yeEFIB3xDQHZ9xdSp9yyw79DBEK6QQL4sTvf88hC2dKr+X1mRlo3GbUusKwuzDmSgOkHC
UHl2dlCLQEL0Qsydyes1YHGpZIYCbknhD/i1/Gab6Mx821Hj6bf6+oaICE5bNwn1Rn44w6MkiuZf
KKlDQjcKas8On8AOHSaeeC3iYDE5fDbyQ45rR9JdPQee2UguySCPo7QRzjSI+5zOLikHyxJ/lM/H
WTIU3UuwX9tttmDUbpYlQfjlUOI4hPSUOiZluok+ZM4rJ/UDNAmrzBBMSsigWx39EtbQcKcFRvyu
mWARgX6ezmwi1T5VdtzFJ4KFTmMFnnOZFzbMhgwsLLmm0GkiUXJpl4DGo5WfA03s7BJ6GH2RfjBG
KIBXSbRfxGi2Y006bykXp6KD3de1+HHhYSuFh+N0T8qEhRUoj7+BSamsC63BYm8KqWzRZ81BT+oO
I8uz+ezzv7uuiAM+1ckwN8+cbQIEv9hjwgYBZz6uhxu4AovbL5XnX3CFXDadv3FjkShG2Y4VFU0M
L0avjo8IZOTT6TBO1F83Aw/llZP57w3/JCCLHXQsZig/YRJO0fCD8zYEk+60atRPlKMVtQNWTLXQ
cWf5kspbaVaQckL0iXnW1DS6tRDolAa2+lIG2sPi6netwyuBvtr0NTJeZUum1kbFnC+nwhkW//qA
SxewNeI7F8rL2v60KNBoHYiNAe5VV8l4MTp6CyKbyMCpX8ZcJh9CrYFuHycLPyXnEekobetmrxGh
qfKiYPLqdhYbzkDqcgxVyYFoGyINFRqux19L92eur5oRYQdBbKfTWo4l/kz2372edqq12ouizYe2
RQ2gOwRitOVnc5hlk3gC7ZeVjIl4J2mAEGGvPYWCfo0xxM/1ESMnT9WTrhAsH2omTk2tBJQe5ICU
Eg3UwZgWRWjjcWjfTXw4CJH0G6IAasPxj6Q2DrUiM5RX1L96WWRVKi4nQTVYJX5eHHtv5hx1NxSw
boS6+YZcX5arX/Ab2b+XOqxoxFWGMurlBE7FyCfDzc4RhGh1wbqjGt2mnNqMryVIKduk0ckO5Zwc
4r+Sfr+5KvjlJjF2BKkrNriqxeVvIv7PXvRj0mYCDp7V+n0Hx8IFEqQ3GyJwkQZB5WvDvKm2ZbzW
+1IxE4cqaualJDWSaRr94MqQSw+lytgv+GczvM6hQc1KJoCRx+7QLmHdj7NTsmLE+Kz/tY7g/2JL
EjBixBMoysJmIbLds6UmFcDr93WDDFDKKoRy3f2cfo9Q4uIQ/KAHVBMr5c2JGX9NgtjkfW86Lr7b
aXtPLhkbwjaKpvfH3EH6RYWvLtDIZKkNyjAz+mt8doTHFYpuUFnxCCvzMZ4w4+TlzJOWAXW9rGYM
unhJe43MnKmMU/P1H6DFgyl6xzpjWAJMC/EQTyUtrm57dL5CcrHklqk6+eUUvvSDgCIYscJ9gC1z
jrl+PnKT6dOrH3tyfs9YajmmrFIzdCW1nGPLsv1eKkCVOxnyrbLYLczdB10DBkGcvNA8aiUtRvMy
6Pc61zihZVPGPdolNtFThPSV34+46XobWZBv3LeuOITu0MrU8mj1WpHpknHjtqKBhRZlgduKZVNv
W8tah19SrYdr6nKzHSBpPlZeuHv4TzrPrS5m1BlvVIB8BmAbEhoj0LtMz90QDavq2FkYeO3Cwwj8
4lzOqiyF1ulltmvqlndzbQFgvbVe1bSP7GNt8YCwvQ+EsUgQcqJADgEc4/FCKMqwU1cEcXBXFbWF
NATuf8MYDtDg7jxcppLxzFkgsu0JOdg8Z1lI5+8o/9n7FuWrqupcHBQPdXlu6MonBLZyq/ecCa0B
E5rCTdmfGxVEGdVG342rWzV4u3misG63rnVOg7BF0EBgp4Lz4mtmUBEn7iyOdKCohHI7wKZuFouh
MEFU7Qr4c+zfkZmLHNw6KgMgI7NGlIPcyosRTUtIZPlnq7HWCDAHsI3fUNtMLte3HeNAtGACoh0w
hFm1xYy9LL8J5VesT112C3a/jCCBwCFm+EA+efzMETBIrCRvM+HEBHxovlWbSYriIsBtWBX9FcM6
aepqFGAKMWfYzP7zaC25ojML1k4ox559PKtX6OGoPye7wyiM/cfCXW510hGJ5xUlANsdPi590541
b7+8fY+PsP84FJ6YNIt4i8cIzx8hma12vprJNqQgHKLER1sUmOqQmatRiiX/A8vVRhUM6eaqgeY9
m7FaXwZedHRNw6n4+jErqiS+LF8xand/SloRQlcDnQN8mKCjzG9npRet7lNYzZZWMn8lx1XkdOrF
Oo/M9jxroeXP2vhL+vtqZQZB9CgNx8UXxK7bu4Ysj7Q0RrIWJHvO2WoPmUIiJ4nyRavFUUwNIWyr
HGpsWCnozrMIDp3z5HQ4uxBwP6DKFINz+pOYHfjg1GtcAzPSBngWAduTKasVxtN80irlJ4DfPbw8
9JAK/xfRiuawRc90aplvhmzPNCeK2AisVvUwPASA4swpF8bURSWh8ZLTv9YrvvicsR6A5ct/y0Ll
4Y3QL57j9HxJztf1tQXMBal7MCk9vl4W1nRbAEmMyHVpd07jeY9N9WmhhLNzXE8jQUWY1Djzt/uk
Ljd9oKd6oyy92Vbb3mViji6upHTvL0opqgiIOFKpFMN3ATJlDnH7xsptrgLLZ7mRrgagiATXdZx0
dIvq6BOVk3EhLMeYPMheXTrK0YRpofIKOecapLIVOsl5aeGuokNfPEhIe4P4V/WuPfD3SnJcBb2f
iTndclnvP0n8Hn94I0qaXzwBITXyiUUygU4/PUiMWPu3ZnA2pCbc0jVuqVFCZFdNiRaHCKBd+sZy
AMYa3D0MGiOET16LDkowA2F1IgVsMWUUbAd6+nFkmXTysTGWg6yc7+8ExjpQXie6MvO8z92tR96B
LotQFulwJVeflenP2jeo9c7BtkGXUl+Zk01rWNNokQVzdFiv+iHqCopbXe7+2EK9dfwZuS8kHEL6
OiqtpaK+v7XQKyUPT0cOiYc7VVHwizvV8WECg593T3g3XRPnQNvjJhM8IfRvU2ShkRGY6FZIEUdN
tMf0SEPrrQ7+TJOfFXlF0ne2Qai10Y55Llktsmm2hQhR2XCvQZVKu2c9vkErrX00tAprqpxMJUAc
DZRKlEMYWd2h+kIdiIRkzG9hxZpRJXxMLMCFbN2339LLkReMsfWUZDZ+Nl0wXJ0HQHU3hfUcl5A7
1qPaPZS914b/LmTqt+bHtkWC3WJyzftHZXsVhjJ/SP1JOozHsfzk0xFija6j4tJzYZTPoxKp/nuM
0D76PipTGJ8BuX1NnQRqwHHT2CC5NBQxkOBnUxJu8EV2LUIO7KbPknW2FNUqIU05BvxPb6J3THKj
NprA0JUuH0judT7vbG13wHKbmexsdf8TeqON1p/NAvh1Ph+MEQNMoc414RC83E/szuOmOVrPMWqG
w/WFBTJAcstNwK1+VNd9cfoHW8F+bb5vpIl5rp2/1L8u7yYd+me1b39ejwM/YnyhQfff+TxzAWBp
jV8DekeF0OnX61POsYhjA8XAZzIifUXXnLxmoGd3BNyl5+k6xkR2I3x02JqTslAFmK7dNlR+d8Tx
O/S7VQdM16jiIimp7UgY4Fu+vyUXLiuHge5Hb11YhIXRoPA9cOHOH4SH6YBhY5YgMvLz+m/DKXQ6
NguSvSe9xpufScSayUtJ5jhLVZnlBYoKKOwqy4I7Myj1GtEREbt/tVP92LxDgYtcebBteOiBqIBO
+XTgxaa1D10TXeM9LYDffBEuApVQqAm4C7mrxSAchK+O/+uxU2Qjf9bp/ZsApQNXtMO9j+DBM3Od
TPNxS6etVHTGR+cTNDwOE5uc5a8LE6irgw5L5org8R4j1P42K7nxvHbEqnK8JTR5SrGCuPQTtUd+
hIE2mGBvqb4SOsJzemQ+lo85rl366X7fDH5QbAAVwb+BfnjngaT4QlpjoyyZeIS9GV2C9VReE2+J
9e74GTa6wMvSuRR6b6HB/F/qBbKnNPQiHKgyef4qMBpmKCSIavehpnOJ98XXTbulyE++nNchrM+X
+/9PqKxnmRVQNu99FLovJ8/y4ugJMxcMXy6XgtbHg7bTL4pLh9Ukc4i6bMyV5Omfdj6EN12/ALvv
EjK+opOclGAIuvGypmmVy+ZGpzKbe0PVvTNinvgSSeFlhQEZla7r4ikpN2jdIvY41HJRq75zjrAt
pd/Dm0mgnscXQmk1DVSUN2zSe2ityTIyUP30xow1+2QUmGSvPyNkfD3kK2WpR1rNUqreNh848Szu
N1hRqPAVcWksTklCGJXaz0zzN9rAuAy/Emx1JPBgntkdSCjZFoUHlOxJ3uOqj29JSFi0Z4LBZEjX
La3Rm0DAynNz5V3qgxEM37jao8OFhYrjWpModR2Acu7bryPWEVd+3iAq49DCM0sKHxJv3pbYkUMo
uSM9FZH4DDqf6uDmWDFdHGobdW5DIJ+DQw7f3uxPeLnd1Z29XJUQvar7gcJROl4yrFD8I0Vrpcqb
Ts3G0bRJycW/9TC6e4ry4Dme9RZ9ODqxMr+dVCAGVY/nNaIoYBgWpTHPNANTYFDgS62v6z5M85m+
UiJPEQyEhCS7xk5Z4iBFhHizbTtjo4E19QUzQxz0hCh5yyhkvKqJb0dhytSzi28sFUrIgpIelQan
ozswVUpUChFVuiuuh1ViVahbwAl80k1O0PzyAGAsBMVVZ/hiOZRcXZxbYRVSGd1AM5yL+7fSVykE
Ygw6RYqUdQaNV3FKqQRLtZrQcidcEeKIuh++1ODizsulERzh0m+dnQnvGi/F4tpoqkegRjR5BxHv
YcNIlVJ1jLZPP2eCIBSkOc5f45XT07Yu698qpy/p6MpS1gvacG9IXb3qP7+pr5jmscuSufG4EzJW
aOyoJpDO9PzPvwpheuClLWja6QKwt5T79DarTEolUBK7GzLuW8hP3Z1+2K0VqXLNeAVIwGU1MhP8
vh+hUEcbEusQcq32EQSLOOIhq/sCPit8aJ/LTkyU1NGllvjpFjp6b1ruA8JEOQtIIt/v0tdT/QzG
ImqkswicUy0gMIXkIcC2IJ84FKSGbGXdVQTEABkjvFqYPcYA1JlBw357ho1xvutOM+77NVVyhCCs
u/LhERhhfAj7t8H6nSNtb3SrNY8FlEeEwF+xF2KJniPMPFohy1nfPZPdm/qOGoWVJsN8bRx351af
CZaeCXwxuoJZDOqOv1EXliWDYSzl1FUldu4MA+NMwxKsWJ7XlZQxv7Veo2qd3+/KztRg0r30Rn+P
6JGRStHxLhVkUU1EZG2QFQq7C3zN7F8ODpL4mDgF/VyiJTH6gMc+UvqGQ07HhcHBlzIfFQ/3u+FD
RXlPKVVSQuzOL+kKLmwuEI3p5LDonzm55qx23MRW5UE5b3HhiwFjnEnInnuJ0MRhxGIoZXtQSMFq
nn2kxgCWe5T9l7tevlEKjplTlgrz9ZQr3rGUR9a9tlyNCIwUUdxWSFZkeRQ7aPAmgBWMRaThv0ac
ldRBOBHSqjvi2jSOgLLixHaFQ7x0Xyk4HhjajuL2hygsvcHkP24CEPHYHiDB02TR3ztFzfr5G+hO
KPEUHYjootwcm6sWzBd+XQYeq8NOZmTZ8j2fitZhy48Ipw8hZtPAWuOaImI9QnZ7vl/hSonLUtly
/QOE+xwDUSWu3tRg0qGhyYDfgVvPohVH8Cgr72tXFrFMFcY0QiFpTgHbfdc7mxxtdVkSxdoN2OgC
m5o6XJxF8dBsRfjYB6n3nszydh+wslPoulyxm0+1RxaowrvUD73Ev4SWUy/ioTgrOg84AlxWQwny
zieFpe+aaSB/lYEaW04/+RTWnUZEVTgK8J0H90UgJeGEEdts3/RqRr2jdcMCWrs7R9AJuNhvPQFO
N2sXIGSGdKXwz7ISmCWnirM5y9pgC/mZdC7fo9ryr94FtN0k9dhVHqtVzBr3XhrwWWa9UjXMSJf4
bO+HXTPGSbGQV2yAIKF6X+3t+qjt7oS/+/y+rxOEnLHQ8lMuxl0En6lG3WMleZ1Io/1WPGnTdgMj
uTglLue/jSHq81tXYO9n0YHO1zgdOXjrH4nmsS+nYvr+amz+FiKEWD7vX1bPZbWrqHWJkOvtONWY
DJFPXszseLUenmtf7ODMha4ksYzRBBavp+0dfu0Vcn5zdUIpZzn33M4n7XzZn40Mgod//sv4fCNU
HJsiQGGITZDT0szdoFoA+1lEXKSA26AZilnR443cukDxrh+vm77mL//gitwTJKlgPi/tLAOy6xa8
8ViJiSiOipXswP8wKmQMsDYdQ8vUIPaDB1j2G+B6lSzVCU17PEfwzo24yi4HoenbB6IEWqkSsz16
6V7ZlKfvMGYJgcZdCGWkrjfP0lxOjhm1hCDVJv08GuUf5Px/lQPaQp5MqHEG6uigJCK5tDo5NCIw
Zk1jQe3E0pYNnc3iFc5Be82LWefoojltORfMthw1TOTS3GNqYmnekanEVgAU/BZ7d8XJw42b3Z9T
8nNt/0jwuUJWdxiCFMl1jwWrsVaZFV4Ab8fPcURA536vAMKyfJlMXPzFzO8nkBEnsBGpfkckQjaj
kDR8/ENvuAKK8drVLP7I1z16ADYrfkXj1NBtmVPFEX6jgV5lP5TI3Xg3AFX2M5n50WcCO6QMXFHJ
lvquQWVNJgTiLwsqlEVqZ9PTDLCluqa6+sOG196uMlkMOChDL7x7DYVLVjVwymmoV9VrGKFQbNAV
lm6vXdtzWWp1n0Wb/+HAV/dza8NG5ErXkEKHtNDr66tTIC29amO7tPk3MNIe9mqIiggSPukNAeYU
S/0PHIylfj/0kAFhZThwxM6EWvHcaulcH+kR6VbLrMrYjon/iqDTud116y10JORfCfQfFItyB221
T3pRxx4nO2oe7KXl5w/B2cRDB+aj2pCws5C5aUS2ma/hv89KWrBAN4snX+eqi7ezc9xEHWk3xOiG
LbJuUK6Jv2vBmoW5x1jKof9CqoQLw6I4riTVSZ+vk/zlbFpK1WsMqnFbGDlflT08QyeYQDIYCDFH
nQP/GY/Lo0vHN9w0/XmFh2mMvdEyt8zRuK5zux89TeykQYUaI/pJBpxX/FHDNP4dhwiH/meRtfqb
NzsYH9GDwU2R/2jHwTxw8lzDS77QJScZ9EULuoHAISMX5sKmMMr7tjkchMg4FHh0xt5MjYoCaBkJ
Ignn+26ufcZ2fSwh7+AREXEU7/fYkSmeDTlMdwyYcw4HU8CEYmGlzopp3t/hzOE6v/P0XLLJawzI
C3Ub/+UUcElXTX7LP1V9WxruRJBaMiQFLrB/YoiO9DRWVyC6l9TPS+WhttC+ehJQHCIoD+z/+A6b
28tEENfk0MrOeX9LTF2OlH0QwCmXWqSUWwjygx67rSdu72fSaL5hzJRCyzXE/UVMxRRg3f+sdvL5
Vq1i9jkmJQdrwEGTFOqBKDWjeaYqntk2qUjowX8PHGwvS87bO9cbYF3ZxVLNrynu27umNNBRWkgn
AATU8j5sEytfIc95+T/+naimdk4HKWv66nuTVDfdLD4cLdIb8DuqmN4ZfGDyQX7twzLZQlcP8Uko
7KCCbKZyhNI70ixh1u2sZnmSFbj8LVyKQ2wkGdcF4FB+tYUhDYMIN1TmhUzDazhmleYhlumlNj1z
MpFcBRPFOwwXD4zi33289uzidLF6K/KGA9Q+fPJZmW9BLbKrOrt9CyyImVd/KYnlyWQ5ddfPFfBp
jr1WG7yKU+125uEDyiz2/Pkc6KJ/b12tmyOXMnar430kShVw6GHLr237WqITxRrzsIVrW5CgWYtg
V83C0E5pUjjwh4kxhhFmmswN0B2ZEfHv2my/cZAXbWA377yS15oZcJZrLFeT9MJhzcja8X89Gguk
aMJvYHem9CG0WN1GW6WwjtnJFI/DUl7gEG5wf7Ay3eRL5REC+uWdkWYI45aZS6FnLQJVcsMZYyZI
CBUiLz/QrKDJBVxXa7Znh6abxecpK3gPEGvG2qCWyoLG6opoK9kAU8f8m+YnQcdvcfR8n97GxyoG
UmHQ8XmK0/0VbiJU0hUGYmmLLRtZUZrlgSKHynWtgZUAKsoUKOHEh003XIHVimltpPzg0xjpTHpQ
nT6hiqexsAwQM0RAsc8s515DFkHHrPeR1pZ+ip9KB2eBOkA23W1r7YryoKT8sIyEt7ecq/taIUbS
1v/tJ7P1ouSH0CUOA+1iqst67tD5nd90hBYBkSIfPRA2LZ2MCBLaaueBpn+qmDiHBjBXPPjSOas+
XIf8XmlqydQi0OPazF1I7TLHaNzdVrPD811mTALZmsj0stSLArNd2QRR5dCM3bfmKgaFnaB/guGQ
3Ro6LGKVIkPl6++vL2NnP4MA4ouVbuat6h61NwjKy7xswz8ixqGYvI95Jxvrpo5zvU7rM5QGsVsr
VuM2LNqzRyS2Ip3VOneA0KqxYfCMUHs7HEN3HjpdAwnf/aFmZ2t7Rbs4LWzO5jMg7UAJcpWtTSdN
iJmlWrwCPsiDS7EffLTiikJTTEIFLDXK4POta5mWpZCbsTjU1/WJT+rWmnMqdAHGDsktqGsNhf8A
wU1z9+F67b3Kd7HOv/dR+E46JIWy+WdqgeU5EeUEmiya5agyvrPeS6ZgbGGBmB42MEHVlP379fr0
KKr31cKpmm+NnEx3lFNHjOf+LpOfoqEGiPsDFkAbsaXAdMV8xdIXYR7YJhXsqZB2L3behHdb1RVD
tBr9Bte+1jMZ9j4D7+XgvDYDmMZzlJ7eeB4VMbNX1ZANQ5ygrTWhcyWQQ/8uFbJoJpw2O4MLxIoS
88duI6t6FZ1gcBTmMJ4Wt3m6cIdhlgs/gZIQ4WaIXx1pk055l9b5lQe4TR1Tkb9qu/3ywjA6B6fa
5PW4UnvD9mEmp61nrF15eia8ayjyndn1+9ub9JYbmWuMuMvEdSkKhUMDMSNoR0d+uopt3eGmCDWr
jUNE5Rw2il4i6DSt9ktoWx7n/LaHtveKtygCJi1IcfQLs4UoAl0pPEsRvGYPpCxL3AzI4Zrp7Wz0
8TnJTMPd5RxgIa2V8vPfk8LS2St8M+klYw3QenuNFtQz1xXHAsWhyevE4tNVJK7zb+53Bk2lc/Jq
tAbyo5LuPcbsi8lZPhz4DFMRJr/UwbCR7yq684L9HSfrWc2Ia85Spo54tT7H4CFEsug73zVp1sWp
YG00sd56whm1xg86kLTrmFXQquO8aZBCmWNFCldx6xcTZ/USQqhxhYSqERR1L1xz1vHndKUrWIDc
WzYmrkShteKwrdUl1yARsHws2A3Mxp/sy5J6jslBg4rW4BcOWu5Za/GtjLopdyII0NvRvnG94EvT
vfFRECDQtKrTkche+VWjPgys2+i7KcNF46XJ32CMgfaiL26EzgIWUyMlytpVEE1HGop+PjFXdEd1
iH3X77oHS8JaKq4yw6qVvUUN0M0Y6gCYLwCYdm2n+FBPSWwySdBSkXFJPG9cCm1DXksDl8BQMc14
Eyo2wb8GIcXSw45ebVQuiSURZ/YND8/DmvNuq0TJSvGqKzqX7FeApi9fOHF6p1cFnNMZpJKzPong
6UaL+MmIA+8SXTG3fh4FtgI3eFUX3kzNhi7G+ziKMBLBSi4zFMZVXc60W3ys0nCBsC4ZD8BohEZ+
PS17Z8DxxsYPnEST3Dad6P8wzX3rymPssoXQL8dCUc0QLua/SKtuTG9PfIeG1br4/oBPzcHKwgb9
Bn0M6pI1z3Geiqcno1qsRyF9nElxTb45PHH6Cbazyz0HUZlKbkH3EW64lGgindAOTNnKhqYfcFec
Nh/OAiKBmOkUlPUIlG3IWkhoiiXtrIcbLb23DPfgZhx0m/qB7wwmy8PN3bw7GuGbVZ0D0hNfahG/
XjTYL/AJm8x4SxHsGMXh4Ud+zHfR6y+b9AT2qoFwVF20OSzysPt0B8qZNk8/V4G3lig5lfVKrc73
XHVNFisJ4Ac9wwVfvF43W7Z4JMCeyJ9MbTXXJD84ZpQseFkW4au9g1bBBNuljX+Cvx/Ev2sONGrh
rNaOOpwmzwgoTZfk83zYPm/5rj5tgXd/0C99qk8etU/07VACC76A7wL94PNhLysHyKw7DJZcn5/4
B7Ez2GCHwzGfi+sn35kuglUU2B76Tc5IGKVhrr21RO80AV1tZW+BLnuiorjA72WM8E5bQl3yTP7A
rcbT+6uPYlI3gunMa3S9APSp+AtNZfHnk9l+5dOHDZ0XIYXvtJPpcm50NlbZKBA+lPBd/tEy3mkn
F4YM6lzhjBe63gne0U/6+pDTMSNvXNJg86SJizMHrSXHjJgQ7YvjRkvyJwbNQ3kHVPKnXcCmLEJS
HEOEPVQR0UlaenGC8GmBazedZHo/6jtskTshyRfo9x94Bq66do7TeT9+VYU63gUHEEWnsiyLCso9
2PvHb48feQdslqFZjvF/96gYH7Z+GY945C7x+iW4j6QJ0R1D/wOVdnLtj0v5fopTZbGhTiUqETio
eir588KYbAzAOz54QaqfR94+KKVNirRy09bedQJd4J0WUPlAV2owxbqM3QvUPemZimxp+tKucflo
0YUAwO3P6+yF6HytyJcsrekzQJu8YqvGRa7YkyoN55sIC4JpPDIFXuqNu3PzV6jP3HlpZfaTptJK
weTxcdsR62vQlt541MBynPCfVpknn5LSwniIlAUXdHi1MTnyFePE+G0WHHx51N688rILCHDDjmA5
U4d0tSsh5brvOebQR2+h0CSxeh1+QizOolhC3EgH8J0nikVJoKnetTV41ZGrk1zp6es0b55nqoSw
0OaH1UmfcFrz04TWolpx5DIHK2AlfigrBpPDKzdjEhXfWOa4pvsRNQ8EIAp/cVMzm93MbKdtk1YI
x0KoPtumkSa+40ImKdqcUy/mFOywrJv5FUenxBA1AStlipr/6wofVReoKmUBkhZt24Mt7k6jor+w
/hmnJaM6vQKWxJNGH/Xsf14QCBfQj68Yrlk2/UVm/HAR1TdasGgP6AgSac05rQml56Q1qmeSiT+/
9SBTpuDTgndKGfnGbz3nGwep4IC6ZbSiCtxjEI1eNmTmK/IdWTwWZppnGQBUzoabbDRcOeYiGEmy
wZ1jHq4SNGYYZWe//7UsCxkHZVruDRVBVpTlSEqydEA7iXJ5x5ema5zULFvuoZAQMGlzNqx8NslF
2MlFgGPmcIvJsK/BX5WDTSebCF29KrEPB5pksE1Hh9ouwEALltPUqrg+uyd/du6ter3XXrAsovg0
cDB+Ls7wmEQbjqwcNxi2MgCULZDckrZ1lIQnD1Hkd+oXsU7AphLChGnPmVN96/dp+0b5PuXZiaKo
xUocJstQXQsfGjSfK4AfEBk7Gch1A3fk8dwe+KC7Wv/DjRZgFbEy02yd12IUl+d1NOxxjyvxV0ot
d85+4s01h63x0mMx01xG9vrvWsHtq9pa9CZTP7u3tKA22VdB+7D5vRZ5y3aU4LUWW+NhlrrFEKUN
6G8lklhaYSbYXF6IswNLt19cdHniZ3+3iEK4ZpgAAWLzCGxLjf4qNcUBMDDTiXUNVJFPt7rW10l1
QlLYs8I2weW9kP0LlSmPuhlaoK/SvN57T0muIfmR4PT/etl7A/ALzYFrDxC2XnTM+RRjfbPEul2j
SVeHGgW60idAAGgKgh3uoQRt2LM9se49Ol6uQGY8hZSUhYwZ6dzkLenms4w2C4zjrSm6b/z/KxQS
b+QVzRQhdxua/fHHlcTXuKEJ28brb5ltPWqfKiy8r36uYeK0S79XVFLpi4qpttUu6gkdzNbJveqx
b4lUB9TxofDFQffokUKtS7jV9MbJ/DjsXNkWSLErxGVSBA/HyAfZCe3H8Ew/ikK7SU5MUjO4oK1h
maIkrXumNxDg00jZA8Tc4xlHnyXRGgLZkmggmlI5i44PW2iXyQZa8ici/k4XwihCtvbTDPFjy2Ke
2sS26gmv5Yspkvb5op8hQ1pgNHXEZfw9MSieQD+O5Wzlzp0VjbJysrDy+0j/R5ChzDyVd7+T6w72
KUpROI2rreApQ8Ic80EZPH4CETi63/cmPR3G9VwNiXW7PRsKTBGrnB0hnWCWX/NW6QiutyfGgT3a
HLCyozIxSPyt/Osv+2IPIPVpOfX7wREB0MMGkLwPwh0SM7QYQd0dJeia5nLS+o0POZQsdVuyOH6T
8mv+a9NZLOkDqNNhe0mJ+NjorPWcDysLLWjmbCT2vjmqveA4Z1XmBd3OxZ+hCHsgbiqfSvR8xo/1
2Fgvf2eepk7UGZIkWXM+LSPBimNvXnRw8LuBHVV0JCm4uSpMNDnz21lyLR3JSLb8OFMsSDKYUWNy
5W2iw8BKh8b9BS/vOfETtw4OWWi9w6VQuO7UP9bo+xi44KriddNbyf04iEO6jAT42zb818Kq4Wbz
3fSpGLxJv+pxpFeUzuqzoWH11VyQaY+HV4aQ+Xpd4mNZm69UvZq4YBDmg3kj52KxuqKp6ivElww5
zYlJF6sSGyZf1SfsiNIN/5aZEGq29aE311POz5RmtXS/sTdy9Q3Paap9LBRu68mGeiMFz3zR7I7y
hCeOlTgFJrweacsTJuiginTughltH4eZ35F+Yz44Mrv4AW9vkje8GUivj91Q3HM8nEZfQUrwcD3Q
FSEj7w7A5rgqeLZAFaUzM+X3gBUc9qOimI2Waka/hZQKr3H7n20rMNJ45oWmBDL0uy96g80iyEJB
m6e1KF/N1eCJanhiI5o+8SZpTIaK6jibp/q/NaKiydnwa9eUDTgck6FCNRe0nvgQUQ0duO89iwJf
+7p+DST2m5o456sfyqrlvYcXLBRtI0dYwTOSN65i/oX5dl9gDr8sbcr+gQkrUZnaLN59XWVhDx8l
R1XARqUJLANy8w4NAbfQvByZsFjMT+bdFj+QoeuQPr8Sh6+6uMAWYN6I7F32sFpIDTwMtSTbBWiw
iazUbxXYsVD4n6QnOrwx6PqDCz562j+ALwxOS7hlYX1UbRjq4oHUEObKzZUkdENc30fsszy5CsrK
/2Hf37MI+bedH3YaVtQ8PnnUum6oQaBW2m0JHZndUoU0X17lEttxN91RiQjKaabt/rIraEx/vokx
Vaz+f921H/Ukd+mS8RtQWD3m+/COQDtxgEFRYJ/jv4Cj3Q3HG1VWHkuQlcmIJ9zJK/VQqPKh468W
Y+b9drCOtFJX9DkzHPMlBD8g5Ep8V4asOU1xUNRAk2WSNFLWBQNenSfaTWSqodPjOf/zbmGXNrRm
yl6A8PJunv1r2jslWuCDXLJ9Zs1p6dQWrB/szfixVnSkzY0LlwcEr5MKU1yz5R8A3PSf57bvKRRI
R+8dJq1HK01Y1c2BKYAWd97cKqkleqXA4scLuJuCZkbi0gKLNZqdJobMCHSF//EFhWYN5rGVzGOr
x8xohqTqxO2UMLeeq5DEesdSZqW1BwtJ3YpvuRdaerSj0u9+5FyXXqLe+QFdXgFQr6InNXM9C8zg
mt3KHib5QJoLjtSNUpEqruuvgnQumQRwqX6Ukv0Wf27FIx5CKQ1mXKmnoM0+CHrpT/czO89pfTAE
f3d7OMokHy+b0EA8qm8/lU6ET+tc87PuVxaJ4eRniAJLkHqT9EsSwqPq5dxc6wAMSEpEyusVmdtm
ItWVoPYVrtD9NF1rvYf7sioh9OsHQGZw9boWxzpyVwiZ8d7sOrmwWc1VnDPvMJRzR6Z7O2muMj8z
O7wxlMwJzbJG1nH0MuF6KUL7RalE8XDk78799cq+xqgHT982P0wQdnZZQtvM1UJ7x75Blt929tlG
/HgBja7z4OyNMMW/dJt9JxNHkVvQVRofr3BVCOhD7LEyO6g3qc3eBfNyEZkO1jeKQLIwrwraLVDg
2cciivQxqLHZZ9eQo6kXnwH4DWDTfCDRfmHdJLADE0FSOpK4zon+xkBYSo+i5387/TyuTOIMOsFS
DVweLedwCYFJpwdwDb+JQzsEd1HknAHoHMxBihUz3wjxXe8CwnH32VXn+CaHrqvKyV9L5R7t23dX
qkUtc57sWap+Xee9mIM4mIMVoZEr5pkA43olmAUnzZkQ9MbDVeOYp+xSTlUD1J4U1zZYyGG8OPFz
QD5gs/axTBOwt2scDNdO5aR5c/rg2SiAH2/dTkZO363gvGg13VBHAZSRYmlm8VmWiNCYDQ87pOTP
f4H8dTLNR6566vPQjvIDpwb8H/Q0xExK9KSIt5KK+6hbBj1nfB514AtAtNYdwIvxbErsW2KXBxxk
421JGNaZDSksvb/aswcGUT8dRXz3YvcsEuxWDb7bvG/QUDD+3qbeXPO0J8LboMwAk3PffW1SiZ64
Lgp7Dba576X7oHDeDX7B7AGwdlNPe8f+ZrJ0H2GW+GGhjux9eiOVcak0wReF70aB9gWanBVCXRrb
+XT6tCgIx5OTssh+i4ApKJ2LPTXrEcwSav7ZA8fZFrBXw3aNDH9eOax9I2HGyBZyy8mzWZokyncJ
X+m/7Xi52IwAi7V5TZgaUtcEbaBIwBusCDWHIXumvZYVvuCPAu+9DX31zyF3uGhfbNa1q9dWBwKR
V+GEeypqL37c5h4/78GTax73fvELfjgveeV9E2T0jOBRmVpqxcM32EQcMsk3SolqdutU/imITGye
6U+oUsdHPJv/4fRnoRrRJ6mOdzzYAn3QU/Scx/kmfmu34EOzdzGOPpIHbQPTA77mnSn/ir8540s1
JhPHzCsZ7LBAlcJOUKmqKqGJh6PZffSLXwUNbn7ed5o/R9BJJjmEGzxIF5doILCZXk1cfqBEEbHu
Dp6IqpamePM4xyJoUHn38u4B7td6iqo03nVeh1OX80HxVkHODpxeGVFgvZE6UMv+NXccDF0zBaCT
/TnJln7s+hdl94GgXxB1W/rQBBAjooGbTzKDIY39so2MkEHaexxDtwf0+z2d8VJ/D2F9zBl7eh4m
72Lc7UdF8bFgv8/Np3nwUFVd0/67HqcY8rVJklAyPPWPOcyQykjQ/PvIHUil+bZ/0uSGK66y3JoU
7RLK+yBOaz9ABxlIb5mVVdwcGM4uH26WW5jJSMNcpWNAFg4Ck2pfSaBHd5p6E82cRbR16d6wN+Eg
AZO7dzCPRcoK9XTY9oKgsr+yV3H2f7LMPfZWCSDSwlKp2OvWUyxHABfdfNZ+z2Ez5a72UPe4AbOw
BUKIGL8jPTacmdcmbeeXZY+gMkniVr7tU+3iKa+La/RV4x07g+5bKfHTJ/N2ith9EAKc6xfR2+e6
Cc1/DTVrpwG563MGELYi2cFFmgoS9FvM6aNc4mCfqAOkdjZJgpCt6Lmx7Fv68Gm4P3embHJrdM6a
SO/rxX5jQ41NrJi+bPYbQ+wc6bnPAYUFn5FgHUI40IFjbtrQ2UILtPXQTESm1AfDVA1bQg/RlTNR
o3+VwEggsBQ6dgefBIyWecT0JrJ1DbAx0JnDAb66nXh3iafLMVylxt7fnxoS+rkpuIdvhc2GpLtN
Bm/jrWuTIHSgUbfpPAweLNcnIf1Bz1YMLtQVFk8JWinx/9tDYFU3IWREEec2lhKlOu6PFILnPtiF
euEo7H+Tpovd91S5ov+a5qFeGnIHfYRuBYNrCzK76nwU41y0CUY/eyIJcVjRlN5HwMwdYHhiMGXt
4PwxrpM16ajeAtBl6iRshtbAM3ENTlLGKgH4jLhPEHW5CX1u9VRNm89E9uZNvTWLA7pvdETZqEO8
RQpmatP8uhGo6K15g9vJ6IV9+n5Fy1wC6aPQfN3CzmwtrFyp6iFZFMg/kBfYaoFuktspflgo4O5j
oSkTd07RjYh8SCOyByBG7WrRCC1IkV+DYnf+AuJuwF9DjNwUDj/9RSBcjYYAQePDVgDH24UGbczG
nIxvkZoQ3Csw9LevwlkzkYKsfq82U9VHVFzVfBJ23vBioaQ1q01crUfGErZtojU0YEiQSFiNfbMw
ATkUsobqKHImNQzUjSAzywMQQ0Zb8QBqvzxlQ6qzZXIHi1NNOVd7eNOPn2w2JqTIlqA9CvNCcb89
vmwO/L9ELsHc8ma6BAMSsPJzPK3iqRcyy1l/vFb9xrj6GLA3l3c5+lptuEdzef5czoGgZNnNS/42
kPL6fnv/gCnFTT4/ADL+8tkgs1b47XNzxo9XpUb6aoOLR36k97sBzCGiiKrmig9q3FgYBdKLgbnC
zEaY1bQ8fvsO4VQJi/bT8WmuQsLUeqEmi3n6y5gFTu4wptMC1TyruVEFaCAxZc3T1ZphJux/Ivxv
lnSSTa36UtD8EoPzI+YfnhXtyXmlJv5i7fYtJpKtcBYM6XM1ZKNd3BMFAMqsQwnaI4/mvc0rq4iU
SxMR4XVTkHNt6DTIXfMUh4RbcIZT82uP2NqawubtHiIS8yeTJjUGOVX4JRhPejH9c0QYSPcE0LDr
hSW7BhgeIsm6KyDTgXGhKgPUPy5i8/aOkosiyRbFWneay6TXdMn+yqQgfOiXSzW5MKIOu12mT2ML
Mfn82ZAj/Z3952xXTbxf95aC7sna/tE2H6GrDD+l2WmlsJFtP2Z3GAZc9LRGtaH+Ae8geJtrhVEO
TPXpUdS/NBQEN+Zb4rmhlaxOq9AnkiQOXIHW4fhKhD+0oiBw7TtmZGC3SQK7mAz+3youDc7qLYJq
sX27MOk/TZLc7070WY0QZIEiuP+tRBGUPc7NnUx0hc4quwdF+5WdE/Z/XZM7GmjKRQRmP41AbMaS
xLerEDD4BMDoEwpVo8P015kPphsB4PqopSXOrolRan1VuRz588NnMqS3KnO5bA4pyUI5Yn9/jiEG
jFSZdE3qinjAF9ndrQGngO1MHZ13OLgkiGczJfjAuNYuJkUiIXDzN9Kub+p1K+ADZHVaTmuut2O9
nL02gtsgnaH6Ukr4TwIp158pM6KY1xgpbuRxEa/kFdy1KFgMb6eYErU9LwAF+bdSBtwepKckfEKj
O0f8JguQCFmA5608PrqU3RivuLuB2CzBOsqhpYHA2UjG/jeI01gk2/a0anHfQ0PyyYlv9M+7p9HH
akAdahH63s4Ux4T+FwC9uRBeD8Rb+O2XcJvi6aMRLdabJIiZ3JxxeM8BJ/8WUTXLG+eem5uv1Xkg
DYjuqbJW0utF1ObCP9dTBEvxzUDcuRjFuhWaxuQ61j9OaE93kydZ2d4eUUwtgcgJCOdGf+WnyFIe
BNZuIc6FyzXTQbugWUKRMdKjqKtBqGi8Wna5glbOauSR4obtPcCxV6wh+Hp9TCsnvuvvZ2YnP69p
K/x7CEHAS8u4Cdx1xxflHX3sFWdsin0x3QpuAW0aON8RGBKk1qSSYCinXPtSb6W2LXNJHREW45AA
s870qZyHKe6P64/7X18D8rl7dMF7aGJNLc9C8mhXRYGZAnmel5sXTW+NfAsvd5inr6A2jZkE9Y00
CmjiWhS8P7GSecRZl+dfSs9hIDddWD2bo8DeijnK/ZB+W0rHZz8DBOw+keiZlmbBfKwaToIxRt7Y
AsO29olB0j0+GrZyFfQtNrh6N0CRcSTco4x3/QTy3ngeUzsluYXHs66EWJXXqw3nsGYgUExg/BAA
AauASapt3xaapLh1V3eTB2qts12rFc/hBuobYzfoimKrd3i6uhiyjSD57+/iDGj8/NPZSySRdasZ
TpuQykg48IVWTm6iAkmRhNpCJgeafiQb0WDoAu7EOWd0UTLShqfWyZ55Fm8Ksx/VCixnHawm8+K4
uwr0V9Kayw0hiZr9aCaNyxuWzKf+2pBRXM1RPw09A2zW7OsecL2IeZQ77XQWUGgFmNZOJt2oCwVE
n83m3X+aiG3M0+e7iTXwfAQVZCtrmTU29N75nwLfBbj5Dfs3mMH2nna2htzlgLqGOWDk58rd0S2N
GntSFLWKirIr6x7GZxTQhHNcAoD5uZO+/CzHqOQ0QELOUa6cZltbRtIsQ06NJlHIwm5El/smb2v8
g5gpE9kpJ7vTI22dnsEJbJ9GmfNK+1Jl8w4Wt60oAKk9jYip0CIFrdWwUynud+PpYNnOxCc2Yu6p
hVG/5Jys4a8Y/mKAgHefB2u41tiHwzPPHrWhMea7oF41qrZ+g1vaLjxb/ihE2n9H6Fo4TCh91rOv
MJ1sgqCneHSdHpOHKU38axCYG6kC/cL1X/bLGScQZVbYSJcm36+dnMzv3ITKI3HGsUQKLetCZLUp
Uuo/5yeCl81yaNOrp7jQBfOYGQW43Kku3e/xDy5LY/1mjg9A1cw2ClGLAxJtzg+aQl9qULxt0LxI
vGOunr3q92IW085EZwYaOhOogVOnC4kTyoJE8CwdpKPVROSHxht9QDP1YU4kbDZGWiBXbqWa9o81
5i8PlPtotzDtQtoQIBodoBrFX6Qw+VJGnW/dwMNwL4Jv9Z7P4DhptySRfAIYjdRiLW/5TrZPg6T6
fDKrvpfRSlB2hxcq4/TMP0Pt2mRkEhW9SWUArxg7tHrzYupS/IaTaWSHdOPwIOptTUnySx0oIE8+
ODOMJ+YU7+/9NZP4GXGMJFfZBIiMQq+Zx98UEeXtKyHftqUPPjczuXXGlFaeSL0T2GQi0HoWUwpI
aAK3CkbmJrdXmkLHHRw8ZW3/PsuBwIrJqIy4ZMw5IMZneSmldL3oziVXzP1FsLNde8vvqvnzblsB
Hqj0Bo5GdJv2/S+Pf4C2TlFl+by96xwWBSYQ8/vbi84SQoGoxU0EOaiIRKSw9beFptmdoQMgZqiS
ddCyb9M7rIMt8G55JjuqxmbeH4haUppri51O1Zel41aZGsZRMtcBEWkhRo2nNLYxkMjEIecKPBU/
cQolmwRiewie79mJc0C3qz9fFSDuqdsDIEZx5xqU/aDbdSrTg7eftNXpQ2+h5Smh0MTpn3jNK0hC
q6BYgLY74rHoiJA2Mxw6d6Bjcnc0c0nKMy4lcfKUwviGHWoXL8wQYRE8TCicRJ5SvYXwqz6yzbsV
sWpLMCQVKfXJEyS6EwftY+s3LSAFhVCV7dt4BuPeeUPQqFhrCHgeXHEaewHSxaHJRRzc4zD42/iL
JrKsEZqtpEi1/rsA8P+zUlXHlwMKDkjdIybgmJwRxLN9ox6pqsf1fIJmTP2oMmdFj/dHpe/iBPf1
mGykdihF+NnOU89hZWOohaPqGjShcKG4vfM5BWwOcXY0m26s0aYRVzzpcPtmi09eDPxxjoJ9VrFn
KFAKfUvxZQZJ1+aUCWs7sqRLbyZ88A11Zr30XTB+CuDkNUfRlazk6+5+I6KKfOrnVKRimqCT8cGW
16SVgJH9VtODd5DjSh7MFYdbAzTwJDrn2eSY3XJXc8uquoaEQw25jY9Zt/Wxb0zTFYo1APZZGXkH
YNNrAniJc2tgnsqJHRxCMSJOYRemVXS6w445+RBKqGR3yvO1osYzJ/l5nn9kkx8ozbVveWFJY3Su
YVMwozaZLkqG4e8r+Ph5dZtUcTiSwOq+coSaeHURjGx2MgA2DabscMdo3fNvb/7rGwIe+cMyp0DL
AT9EmsJHwz8/a9aIbmLdieSfGyVHbZQIp2UxBtKGRkgvxXA3m+VGnVwaI0tDt+rJf1aXpirX87In
hdPH23aaAa0xpxUmEW5t1MWi3czOWcRkAFLSVLlCKrs08HF1VrETS7Bpke+aFvkMW0cHtoYFkc2R
MugSPqdWcITzIFbP0pE3BD8eO0aF2+YXmu+ErvUN+0iNVq30Zu/ZYq+fXeyqszPCCwoQBEi3MQ/W
C54XIUqgrnK1JcRpeVU3K3xcpBWBee/h47SYc+NyM16PwUtJYsA/ogKo+DpeeAWbg+J2uWR514u5
jEVv8ZH/or1heBpeeAZ8bcUQeIDs6tcSCVHNjP54k7w8v0ipbnm7YBhrbKdz60VsUCUlbqUuuRKk
pJBVp3LlLYJut+8JPAI0MHa069zJOpgkJ7QZHPosPJDTWcYuCwJ2WRWl5QShqdEdFoq2kz3Dxi/c
Ullm3TauN7DmpJMOXM8mG4fFoAB4XVPyG7Fu6IzAsJ7dRz2o774zQK8KB+SvQeR5VYUv6t/hXxa1
Zyrb6bY5aMljLNFwDur7l4HP0lZWKCAcTAJvbLd1U9jth4FDfRUR9Hf/G/ZdNkWB1xFVeAT0YON7
ZdmcF53GKSxeacGD2chQ99sQVQ+6ryPrsuDtPa14O/pwT0l7PEbuRCVz/+GJWzPNpTqvI+YuaoXU
ne5XgYGGzzWnFoK4qVUhWmp0qb1im/34kGPWsNyzH8yk0/xO0gF6FB6XFk9jCI621wsCpOkVVEoU
/yPhMhMUQG1Bfu1y/XqFteEF94a60HGxFocktC8irQ/so2cwKXCW3RjuvBgElDkfK/3II1VxAH6/
RVEMTCP5oQiyhBPWeg3K6yCyvHLvd+yTKupBCSUauGnrnp4G4Z3XbtcwMRv5eNR4aB0IamqcEAo7
dlPv8qvQBHWr3ojl0ty47gbTq3VR2s9MqBFsuwXGZ1iEk9mi3/xBGmI4AKSF8Lemgyuy/cMYMNAS
ocreSEKgt8wC/a31le8QfgzMXSxu10KTH0QDgX72Xq7Uf7456pBMXSI2N9yfdOetGdpDq/Jcu3aW
L4pxy5hcD7ZBVeLnQmT2Lg+T6u+AWX+6WVD9cJJpJ6xFVD+P1Mmd6DsMxSNmO3vSflhfmgcdZzlj
w891FSWKV4iqo2uDSJ1nyEIgeMzHfVmGzzfP+wvVTBqFS9Ux69zzwk4Cr7CiqeFEYBoF5PuxiBlL
SQs56DHPFPD27jDJV4igM/Z1ZtwFL36FiZIlkYRNFbLwVhjtwgyUR5sNpnTlFdByg/4gpmB5dGtg
gFdEjPuwbWFGD08OiVAqTXIHuI6UnWp6BGX8OktPGR6HLQ2/7hqMrXVONsPqF3LuKmK/ZuaHZFIy
vA80ZESWBOI211Is2aPUTGZ67LZWHu3xnJ1pEpVH7C9O+3SZF96l/mqY7BB4jzZbh7eiIsLVsIql
cLdXkwDZJBTMXcwNHrYLZ72D4WzMu0aVSemk7VhuCmrzK9BdryJ8IhU/XzbDUOwgiYY+vyOx1ArJ
UlRqisw1M3RayFoXwEpX7dbbZgHOeEnRnleG3kwWEMVi0K/J73E4NFymVVW8PdS8WqslQJb+JIgL
k/fmq70tPGYLUsUFsdMZV8T9baJBuCYCqz5qyhKCqjOaZYbXjKp9TyaQDbhQLT2g2nrY1gZcJmWH
gYukwve3WX47/0ooOPJUfkviBLPWDR5ycm98cZ1Bx9d4x2Ji5xQ5pfMrDoNe67QLM1pDVG0a0mgQ
6ipXCi2KMeeVyn/Z9lGQMhuzMAPfYpXIzs0QqIZQBwD74vFAfZ9g/bhtCAaLHYLDJESiuAO7MqP8
/WI9N+/NQOgY+j0hFaXIEVh9MGdWVJtphSAzRy5asOuW2xjBapRl8Oh7P1Wr1Ton08ShgZufN220
vaqc6BwzQYNMEWWCQRDXMpwqoc4D+LNVPOd4O0Y9Y0vlFstaXyuduLwB54LnH1L+yIqyLbdyTGK5
ZQ9N+doMjgKMHQtKDw1Uuneb8cU+VMdolk7HIEXcPXGNmI/k8oaA+1kdSUUDZ53tjK9sNTPU7mAP
EZU/og+XanpSgVVNx75BI0blJn+03r6LerkviH6ny9BsxR1jYsqhaiRkntjbneUD097Ggr0ylM09
/Vcd1JZXhERAHLl3D3srucDP+yO/la8dIUmoUaOo+QA8At4lTFf8KBq8PXyARhvC3Qzg/IOgh4bR
OKzxF1H0QvvkLbBDHZ4l6eH8cFPGZWLQVu/PFYKOiE96MvLZ7QioLqHamTsLMG5eu5gyTarqimtT
DBwJr1HonJp84CEpkbkxD1jNDA+jjBwY4RLN2OkFsGp5tauIJOke1aCOcZD1/EfT8A4oTQsoKSfV
3nb38PsEFTpeJVMEWZTbdFjaIAUIE0WlQ2MGOiPWVQv8mXduvVSNpmjxFOKvPr6nuYDjEvu1UrDb
2Sw7Y1uLhmARCDscRNAjrKBNB0xAMZTjzL7kzW5sjFBlq/0GHWxhn0f2bJk3xaOzzNJAJeyUKV6u
5qaRf+LxURBZPTkGtOAU0tJjD82xm5ZeEiUmqLvaeoFE/wOnc1mDuPytJ5YHh/ri2K6EmRPq1P5b
t5LqnF9hjhY4ZN4W0G3jQixnjt8BOye2LKxndDZOgccl9NshXENacoFGUTlfPpKRXoccY3BSdm8E
X6fvRtYhMo/xHJ2MNK9Y2SzA+ySjxSkl4MF14EkoCb9StDniZ9UOO+oAM5FUf5TzdlViFFKk8RPw
fNMrLLycZQxs2Mdej97XSl2IG2CXrDNa5Z+7HzkBpVuVBJ8SmtyTixby1NIGFQCNrzgbpHSj0cxt
aOZ253eDVN+bPfAtIS668nXh1uiiTh/IJCFh/a2yZkhOwshLHs48BH1eV5jZjEKfiHfB6v1trkiP
jelIeBbnVnNhzQ/SBELKX+o33BJeNsamA1rFJpAwZ2BzCex+zEzAQNPf+OzDHVmu05mBEB0+IKlj
/kKNsj7CkD2EhcW+i1bvp1OYoR1t+pUQcanjSXpVburu/7svz+sqi6UdocEXZmzXNkwJErYPergj
hxKGoOIAikwRlFIJO2Z5BNNqpVzwFO4I4vbzKYDLkE8HTc3hhvh22aOSUhv0C4ko5E3UXNbnpl/J
LPl3hnw3OjKvbs6S0wByr/OlPhqpr/DpMz5iutvlySD3dgan5RlfOaHx7UxPtwcFG2nOHR/Q6xP0
1S+RpT3JhQ0Rpop/KFj8UyYd/3rjJO7t2CmhaijYfwpH0Q6kVNhk/9rG5zY23iINuGBZtLAzoN+z
AbVJB+pVe26+b3fyt8ndDAo2vTLAL1ecLxB1FEDSsVDqyKYhoxHiZp9MPsDKkkLHvd+vjXTLPegr
uOrowWNLK+0Yie3ya/3HIiu5WoyGTIWrRPz1GSt4oqQAmUQaeLOkrs/da+1Q6ddbKoN6Y8i/4wqO
8+3+fhNZA1WcubdoAJZinFXRzwtfNfjYUWaLDo4/vApmLR2ITmd4XOQk3Hu/nX0cx4aReU2HPhk3
rWQF7VwBXrl2jDwF32hMp7mxVu1Le8j3Ebw+mrc0O0U8tNomXTJaV7U41QYyOWVq9em92SX8zl7T
LD5nPofJdijNrJTgh3I4w3SC/lXTOUGDL9ubj6arSvsTM1kPYLnjXi0gvhu6A/BXZFmI88uOO6+K
zvgSPGWv5IfHEnRCN57km3MacQPIq2KlBbU0VO5h3rIIGCu62pk29aTjQvDh4vLVkIW7vIgr1j1R
RxLWv9sDkIKZdMQTzHXzHGzPmNEZK8CjptmydWjSBX5oo825mlE3j//znohQQFfiHzTyCdtwT1TP
pfrXDxPmWHAcTCQyKr2VEZGqZbHIIeR9Fsi/m1Mx2iQYMZUBJJMBLOLCoH31N8QN/xgBWu8WoNpT
xUqCMqE4ym7+8JR2YQoNkVaTITDVGE0/pHMfWZY80FwCojak0DlyHkSxe8/BMle1W7Zsc39iSpaG
cs8ZadhssmAAN4cKTcTODtmHC3s3R9+i7C+3WZvQAVZM+JOW+kGW7+8jcFWZ/5GIScItKRt5xJqw
czfJStrHkvP/Z+HMeRN1W5YRR5el6/prI/D2xAuBHbafufbygWwcN8sRc3S1z7oUFad9+GizujbB
PzhvinVclyg1MmCxLwyomsvceDevrccdoyMojq1E72G+kEtqQiqGImnlgw0puPbRNLN8qLdrR+Lw
72R7CJ7nTnzM0d0GzwD2ImAAzzYaw7gp50p3QCd/+ujHgSr3ghaV+nBXQACGy2SXpyz5tSzYPZYN
A9lRgTxxnEbsY6bZMELZn8VJQ6eNlJLBos8D9WNZOOXT5NgKMYdyZiBj4y0K9R2mJGoqUfwxOpKk
eTvP4PJ9VKPAGiNZkBN3yfT0xezdcbFUodbGxb1ftWFpe3h2AS8L10eP5crPkame3dvld2ni24WF
nkrIXRci66IAPsmoyJ9GQs5LBziNS7JBFmKOmVxCMQ6o2hcSAjdr89ZjEZG57kDyp7CnaZWqTyiN
PuDDmVeMT0u/s3hXm91JTpqdD3OwbaYG2LSTOpKQOpSHYGS8xAs47NIBnI5NB5strYqzniVlUE/H
O2CeuviSYOZyaQLsuEryvUjOQAFmLliayTTimVlo6lK5xgaUck064HgcHW1YxVJzu4BFv5NBVdbZ
1ogVfwDCaM9zdeydug65zy0yWfqYTD7swg8vKC0ub82itnwPrl4J5RB6n2G/zyc8Okh5nmeTEMVf
RKsLTjK1fymvl2YphpYNO08NiXPgSapMeb14X29EcL0vEjUhVpfBpq5s16P5cEPlWkt8U/nF6rn7
JugHGY+93SFUl3IsYi+ublgFg9mEdSyKha+7tkQiI97itEEG8STJzCy/tuD9Ktk52MYEzST6qH91
ux0/LlvgTPfIeWctALzncB5ODvzUlW0uWTQXyHRroTyfM0tCNli9Z0LLoKpNIVXUefoP6zFGnLNf
ZwWNWwsEa3KTp9Rpn30M6RHZEn9YcvxmcecgstycEKBMRqaqdY78fe4zz3/o/8GdFS5g+VX0KhyF
zRE0kvX3naf3x7eeqswqb3Ra1zxhrvtddxts+ZYVJu70gFeGGVyUcU79R9svSx6n0udHsuJ0Mk30
jWoTdW8tRSct7E6KuLbTFwz6uG627O9ozCajNyNmL8CTgwhwrVojB/WIA47rxmAO8B6O269DZJiN
L5hkHIrB8QacakAjk3nAMKbVCmdTmD70h62xbKs+Ck0Bpx8cWuL8HgPO1T3fv52t4nGxK4x9V+NU
WOjhyJsUs2ANuUOiSaunMdSbKSryrliLlNS6qD0dU03vAjFEoD/JtgCoY7hwyKt3O1zd9lYzSu0g
UskdTlUxENUxQpoo8E+u+1C6fMV35LD2VN9bnMsyYsEokAHz011szm3HzFbUH30Ay5GHMUdLuQyq
w9h+NoNccJ1zZCmhyT/8BFB2FZjJPEK5Mh/NJcRsAQfZn+eRXmcdNlTWQE5nGZzcw7KDSD6nSJzq
U8CjHkZA/DshxBWIIsfkEMiQ1jqoBVAzRut4x8yySh4YDC5PWc22ovdU/rNZu8iqGwsZYqL/IHlb
PfPkj/i6KV4Uux5GWiWqqxzyCOoOJWlRFQgup2iH03K6Uieh2ZnE9GdkPhTWDnHjqe2x5q9DmRX/
6tx9/WGLLm90//dUBcZEge7OkwycQi5g1fNUyBCkJIchytM/Oxcbk0neYMKbfRhdftkyZfeN2q8I
kX4JlaH5tZd22wSIIDHUQeGU34l6HW8Thb6in3hP7XKLKTx1MloKPNka5D98Ak0tA5In+Aqg0XNj
S0CFiO1RczoJ+grs4v/e0sIRTJUpbd1A3qfchpp8Q4e8pZGAb6/fAEd5KVagk1OOLlXBK4Ne7bpZ
5VgSsceo5sPH9isPaj8wBo/gKf3Kw38vgwuby5IiH+3l/YHxLp9KkadBPd2W3r4Kfh+L6FjEvXN0
GtGXQ/wqnpouryEp653UxNOjA6/Sl2D8/GHykpBKX7r65p8H6Yqrqf1FDeT6qOXvStJjjkyqLHtF
mXYoYDrLobKDqaXDmiTMU990bpsF+OTUce4ivq13Lq4u9NpPTtSy6THvNcRP3AD3jLCHuA0LfoW/
IVXTsYZfX8jUKcwNzzJdxCfORkgcd6t4dc6h3EKQDSVTAPCDu0UvzZMvlLiahg8pSgy4vExcvHKB
bu0BB729pQKlFq7Qwr3WtNwvsiwQy5ktU51Zgfhu+GC9nqClvQlwQP/h9cEZvdSYbwmt3CvJJ2tN
dzXIvDd7xs1d8PXHKqQdxnyawixrCyXrg80IABCEcB/M4QIVPG22BKoqNkxZDTkt9fe5i9O1HJGk
2TPBYO2TNUYiT6wsuCEk58SbWh31CJTrZ01QRKj7h4h63NeN9IkBslev7D7dNlX4dNZScyw3PTHl
1uWAO9tnH0Vy7dqCGQP4Cejm+YMbb7eiFiq3MNuBmIh9mO9RDE7IIlT7USoFukarUhRAlbTLS50D
BbR8Qxzbi8YFmUtXJXzg6Raw7tq2HR3hrVaVHSrc6QLVSbP4d2SEmPZae9Wf4pcV7e2yk6C520t0
QJOf/OOQ/00jDtZE8wTeETloRDd+vWDvbjXtAKFmT3ffejycFri9zbSytnsbaYD9tNzLxeKFjRXZ
v6RHbPaFoRbAD/0XH4MlD8mKaHiEa0BdIVbrXJ7YnjWQ2ULWkz8ctcCIXYqFVDl1Dzgbu6qd/n6t
dNb6EY8Ipdq5y4vup2RJw9kuGbvL7/Q17hG/4xPnu3NvE22fjjc6QjpSI1eFmZgXeGBEZuz09ixC
N0c1k9uwBMZirsLDnxCMbVAQmtmAVHq9XXcas+hhnDH2mJLNaS/EhVxcTrPIMf5GfFI69BlRsG0n
Z2mofzBtHsOTmFMdc6aQJC/H6lCG2YbTnT1iweKp1OKOc40eLNglXV+xXb35tzncLLbqe1Y81Lnv
XyFLoFmSWawnD8pQivms9asLFkMeoCF2ch31fOiwxi3ryN/H/uSQRDQ6cj1kZv4/F0XmrQAi1y3J
3TjmhIfayTiNrlPv/h96Z7fBd7oMYN3uWxLK6tYq+opwv4VxKedt7PYEPqByjDInfHk9bIoHeGHD
ZDPSs5DsRSf2jCSMIq23okOGxVZ+g60QyuQziGT7fSmSI+aJHQF81l4fqQD0IELBO37Ii5EsrONj
TNJt2+XZj39MM6cMGDr/MkqA/JlPaZC7f25aNJFTm5Fo+9hxiLg9OHUnuhn9dRbzb8nQK+vCzNdj
NzOn+38SDwJ/9/JBCxmZ/G69ijqUn3gKwAEtsjcZIb6esygmHgRF5pV3o9aH1+U9UF9BruO1l3ES
qR8aBYVkzKHI/XwtPPbz6y+hvrCr9G5KY+lRtBhn91hdBhRLB5SR3LHnOIR7+rz3FAouRJl83uoo
zMjF3J7AdUqUBd5MpLPbzjdljlgNo0d8VoAsgV9Fx7d+N4wid3D9cE5eW8SwicPptGfQEn/gPiLl
R50BGalpaJem8MQ5MBBdmheGbjlWoHg5GkcUZxK4uglhcu0lVWVfkTEnGdJXN0keD2wYGXQGGXyC
LsU+/nJnM0NxZK2yAJ8MQ8wfY24agMl2OgERWVbD8RcnEIzFoPu09vQIFUGAKnp/hzAoxOWuc/ga
g5K7OWTxD/XXwgBtYDNpWEVavGpknyTN2SXviWtAF19PTH68CAioTsMxkbTYC5+0Jt6iqlBIiGEc
29u+kKL5h4G92okY55z6ADPMOC56bmOAob+gkbGcRydAOH9j8n2eCQuc55465EYjnEyFTL2H2lyQ
LbXeqnXhsaC4SYfsLbfg5f4m4CSC+J7ooV2lxgW4m+TwUe21B8kVUyu156w2inw43EMT8uD2a31X
DxhxRJgY+ClpmIntUy2mT2q/X/8rg2nzClgGxwhJ/7YP9TWipWsJ0/vL88Crmke79lZHAZivHrKp
6WNnQE8oEhGPg3dqdrNS4qBQekzr7C90ZBqDcraH9dPRP7v4bS+Q40VUHspV7D/JDFQqu6u8qaRp
jUZ83Hi+0jY6xzp8sRWDCT4hxIXyUvCtm9Q6SlKmQn8uEpH7WtEJ+RGhfblbAMJr3BEznREvr+Sy
NNPflYzZ50qmNbTipDVmUq+KB3TA+/y/W2K6C4YC8ye4SPJjIPT+4tyjHdm3jFb35ulA2MvzqRLB
bq3K96n50m1/xHeliUhEduwLR2U105nMX8Fh4xKZWAnqQ1TfbMA5s5eT8NaTXxa2i5D4kBm6tRm5
I9hC53Eyf38pbBlXL2wXBquCEGUS+6midpLpBIdH/we4QxofW6cezfsyWLuBiEsHy6bd441buB1u
LHzbbLoUJcnoohbUusuYTQuAzIKH8K4qxtBLRjGYi3vZG4eQYwvPsdrbKdpmC75rluN8sMCK9irX
4mUyDLXuLkwmG+KSkt2ah5L5jx5SfHAkNFMK2bVOCmGyjPz9s4sFu679Q1JSGwHOHm/76P99O01a
sVD1kXZuFKeXYozXFADEbDiwthNJ5pHL+HpBM32sHkDhv9bWM3OdG+QxXSUdlt4hxVhPBA8j+IU/
zOJnrg/4hoaa0IT6bZ5WeHiAbL4xuT1v1EIDAkgzSGShasz2q2GrB+T+2E+SbkqoJrRVD0EYtV2X
AFRXFc5J/4vjWegcjjtGauP7f0urA8XbSp6oYF1/2ivBe0ygactr/+Xwrjo2giTT5m0v958weoZ6
Eq9kiz5czTEJvdZnMan+kNOW1HZBQFBRwbQoLDjx7oTnTBo5m6lOK48MmR4l33NhXSTr448uSMZj
wx5NQNh9hVr2Z1sVMr7nlwcZtAmCFj+4LwIicLQo2H4I9woCnzQiqaP9bkRxnYbRQ1Lqb+uf5L7i
WPCUpFWPDpGnkF09b/YiY9zSznj9BPbSbGdaHiIdN5KggUSOI5O/WJyylL3QiLxukn/IUvAhwcyy
M3Iv771gleBq+TJ4DxS1R2aBhtz8V0zckUyHJLNwXAU0nN5BJtFy53hxuleN3FFdmCtwJ2XmThu2
FRekt6dLSZazpoaVNFy3TytJeoNv0cdbbuYdGC6H3t0cocIMmsED/yjIJJvA9ode9cmHjKiFtPKL
DThLa/BgdH0NOnFFLSGcDyfROwCYhAuh0iw4lIq5Gq0X2PzZCmOjif11ep31fBPdNzK1I7aPoEli
8Qey4Ag06mm0WqMkPcS4HRKyeEdSRaNfO9lOv10JcrzAy2cbtUExhhspYfAM1nvsMuATiRTnfa5f
1HFejP0laOsjXdhs2YYIyewyd6dV4rbx5mvbsa+jfSYeKrTfbHOybXcUhEkJ1s1R0OicaBxzo3WE
SBUhYWNsQUo0uRJDeVU7vqhYC9V6GdGhjS8o2rfOEpadmLp2PVcnGl+sJb7LcrAou3xZ9zZI7M3J
x4J5PZTAiOJlVG+/x6D5lhFaAG3FiHah5OD0sWBlGYz1Dnq6VuXJQt6IrgrxaucyoA512nCYDmI8
n6jPVAYehU4bmp5JnUKmutGIKwHVxCeJQYCwkYbGoy5XQZEEeGo+7dzs/zCOENeFuaD0ABrgJ/wE
Tv0fj+j1/6kgBhQXtOnbUqeQCHJZjAtaoExCadqs+sY+N25bOLv0C3kFzQAWPU0IoIXbExl7hwBz
me1PhdCodk3SrYWlgn58Qzf5ICepGNsOdY/T78rpuo+0H3sizsHfOC2COJCVfjxjIEjir6g/sGKI
t0y/Mzfm5oPFEi+WUZY37xABaVWtXceIYu1DSpgJtxIFku9/OECrt/uXJkEqeQldjpHXyW+rKbhv
QNcjbexp451xO/E0VG0UI2BnnpyEW42qvTzRJ4b44NcBr/Ny2WUTL2wWglGMrkvevR4gdrwNPy/M
8HxHYjTzdb3kKqlDNfynguUBT67GgTDfM0yJYJ5SGi9pxVlgh3JY1qJieecxsYCm7yIxZO41Hi8E
2KBk2zPDlJJaF7i/JkCDfpnFKrdrHcjXmdIe1qhtJFfwCEahNffaog/yjpyX7UU9UMLnya/ToUbr
cyZZ/1mrsEKcKSVLYQ2M3hl8FdCLX0INFyh+MvpdZVm0T9HYehf1DvyshtubU1IELKa5YQkPMzzD
gebMvCAlf98Pyq4kco9XuOlz5TflSAnyfNsTmPkWyPGheZmZQVwJB8mCNUn97Wwt7kIQzYWH4xDO
O2yEO1cM55XCT6p0Lx+Y0Xt8pOSjl/C9p+K8sORIDFJpZIA+RhOcEyO+TSa8MKMCoyabJ5mnHnaS
Vk71r42LvRkyto5nLDsa/Gl5FrA+trWGCQbBPSezNuH3rTSfYp9QEP/FT/IMh5V/IwfIIixxgm0K
aHBRLXhh+OCy1XGegCudyzB1FGEJ/abWkuNyToOsVhEPBtcd/V6TtnN4hTzt8j7Rc5Cc/Hu3pq5C
7LIMSpIBV58XdKrpg6rePgReFAHFOyHh8ALME88dBRSyCOvqyJLajiF4JgG52t6mkJzE7Q9/FuVS
z2YYuQ6kx+L9LpuJoCvRIo29sPFT0+J43ycpUqX+80HMOaX7ebhysb3pDRPTEPj0bY9060KG8Khn
odoGE8+s5SPJ6L/ibbwKrSalfRNrdeDIxdvh6Ig57yibnlaE0OKWHUtITCaD/APgD//8TmvuapYC
wV6+B4AiKWAkI60vkpvbaAfjPwp81dgN0xHotxAA36wZrPBKbg9l5RpPSFFjkj0dIdDVvo+sWdE1
h3wNB0CH6Thy3bMM59XDdaWjBeBZwhKkNJFbvgVgrhtBd5+pWqq51mYJsDeevRv+NXUzFRpJIClt
R7mEkneo2QDlUu5pQrTjbUGIeXtmHu82qWWms5YlIy4LKj3xGi5fdGBpf5PLCz9mx6fs6ZWWMFQ1
gRTYV6lnlPpk17pAae3aobp/lqLS7uoixG1PJNquOulHe0g54A6tn1ufrN9D0N6jmlehk1w3n2QH
/dtQl3671SdZApJwMiqjGYoovhuECQcPW0aonk8cPtkZ+wzbQvjI61uKuklehdXmVq4e+zqduhFr
uV4Seo9uUQfdsLbnNa2flm/yF2a3qMDi7qlSNVEsUxJkTLdGnKthYYux24q/sKVQyzc6qGpvZeuV
l6K2+4f2tTudQztabuZ5ApTIUuluPyMrmem/Syz64gTbgwT1zmwFkyzkJIhFHfIrM/5G2qTm0Vgd
Pl8lpyPX1Z7N9E8i/VWqs+iEFcAinrrkpv45DGo+vnKoTkUXit4xsIdjoFWYIhRqC0qqeCQLFuKM
C01QYbBfgFe5kfrfJ2uoWBqLmpsfzZHTzB443owK8k3ytYdYMfLfwDaY3XRvi83vaShstwAO//nF
sXYlok7St8drDnJrmbiDEo2QZfChj3YjnvlEfJxlsXFKFOvwcHcmxHRb8xo2xxiO0csO56skKyyP
HvKFB6IupNATt1ho6g8Yhaj5/0BUNmlKVpzU5luojxqL/dM2HKrWmnq/veh7ZbkGCob70PdzZfp7
PzV3bhH7D/xwVI9yzR17wnKPKOsdP0Au8APlWnSxLOVYrp5LnirzeZ+ltkloEoKdJTEf0slCsdf6
m3xTyIg/rfp1g43QEem6Jba0GX0ST43QgLuNtPEjLqv3aAmRVf1+kUDyCQO5qd8WQVuiQvOOJZll
4ahN+Nv8F4jyJijF+AkOc4cRZCUVDmObiiCGnt5ANi83vx6+WbZlXR6Qzd/kM1ybW2OvjiJRaiZd
dvyMRphbiOnSOsXLr8bvoXVLwLKN4flZ1rsMHx4Vm3LZeBb8qFnLCUrZuTR4LMOFp3+A5i0BVrX+
ovA5FqRwv9yLROpY5CuhconNkJEhn1RJFi2P3Wjpw8kInRpAUkMXvf1Dw0MrvXdNVNcO4DDed3ov
MdCOmA6xj0FuEjH4DL6YnamBQ7ZNJZAMSJEtlOx9JRA6qNnag5/u1L9loF7U5MlIjaHhNB1XxQ7B
jXbvzDg7DadXaStlLzwQMOwoIi33fYhJIq+tnCiYoiKASOHMdr3mnBocVEWdG6u99Mi98PYE/AFK
MvuLVAUBtZuKLKdsiCijXqq2Mcp9B7safOCq+ZimhzKm9jR9Gpw9jzujW46fz6e2xWCRYQC/Th+o
n+NX9XYnzQbt8cj7YQQefV3avxtUq7hldjAQBeYNN2bst+lNQwTu8nP5Yj+HxvQMQX2dG/fVVBpM
32fkkha1UoTvrBMXHinK3+WdrEKPORzNx7fKFTAZ0OSXGZ1STT830r3LCq9//D+IFrxD+DCm9If8
yleLny8WQmLhWyFV63H87fjIauDiHv9RGqmMXZPEDWKvHjlN87rktLCAmqHhd3/zFmKstg2OlqKi
sH5QeYWcEdpp4h9KcC/aL+csKsSMEGprAItXZA0G5TKu0/PEhLsY8EEWhv8fTpihgW+m/YPa+/pa
EbSqM6rtrd+v7akQ3XZ99qCfzJ8V5Lj4uEAZ3t0l2SVACKiYUEZZ5XbVzE99uhyjYTcIHBHJE8x8
5TdK5CZwmIhsyZlNU+PObWNok9Y39VzZvBYfDGihOROoS1zWqECZ3hRT9TLXsDXc7L2b+Y0bSELT
VvpfKroEKtmLKBWpnJMO0JuHUKUBNhV8BngZcq0i9ZtAzGWdJpx509lPWUMFD+E8m/6AsXHP5qIX
3bXkXt9yUCS4nhe33VtXtur4xf1SgiywRSYdAEaxU8nunw0IGJ1xVUuF6TB0jPQpcNL8pc1voh8A
gsvwQd9xlXt9Qb+6u6buX0cklU6Cy9AMukf03EWneLfl42m62DKmUhcHQIQNj3duU39pa495g8/b
HogkOFZz9COANHNBqgX/IkA+++qEurwwOoTK6Dwt5rKwptkpNnBUe1mLYlg7Eu76Bb4hxXyBIcij
FJmwXzeiNmC7iJhATTl4ECnQG/eMHidcZtMPIeJ9DfY53IMPBMnX2VAtsAMsRa+AYUYupMKVVQFJ
P5sSKgcoLx3OnTTJF8Hdr2Izo4w31oPLIWrctIGHWtJMRQyKULlM+/2KJ6V7c50HoX59GuDE4IB8
SYELJJm0+uDnpypajYtNEFtT5lDhK+jMBu7u0gdx12xvtahdbZSBfFcdOvpJJDz+KGa6AeRoHkqH
/acQJPptYOuyxo5D2MHtYOXD7x0hkcjAcG6yUBfwVgWsU3yWTtPSuMr+5n2B6iDUWC9TWp4huZHm
6K5KWy3Q7qzwA8x5GT1NpSjxL0DkN29KZyrHI6RLumXV85yWaqsv7MG5w/hLp8crwSRI+E7ICXP2
1fEn/MkblADO3to+4d9HmKi+fnixv4vgha5IOvFbeYvdkovH6tjvQYedonvNk0tk0vSVz1KhJmqs
6yDec3YWNi9DmABKH4UU2UJ9p3bgIRMbp+0oj9iJeAIKzUMtoBgKmGNX+1KsIX2qmXubuZzPxyCn
fOqaBZVfyASdo1ldnas8vNdm1ePJgt8MphyuaBcgRzHXDGADj7lGeDgW+5w5pC+FcS0P0d0J+8BC
hAMXZ22iON88AZRmbcx4pKHWqEcuSt7xekzhe54dwFi83fRRoRO0k99FizzUjv8Yd5KgbqqUkzyO
ks5a5hF33C+zk+7ESNVF5H7mLZPrQ5J7y8rh8/zoMpGmhdoJ7GGlYCG/kKpFOJ+ihJXoFkUfPZmN
CV9pcpMr7nvMv8c2SUC08TfvGHnErCYXucI3rXP3Wst41kx4P77oECKuni0hRlbiAqVejqKDUCoY
1ItfLKTqNOJx9o/ZqJq6uh842emVj98QDUQoM9aQX4V3hjvjJnMeFMsVHKqFtRX7hHqRrLujhMGU
f15K9z3APdRrbOlevCwhm7Lr39BNHsqCIZLesRjH2zmqSmh9ZeZzsWNP4NWvOdDM5+NMw+oH5aKE
V4rCP7wiPdPTn5tDbwyEBa4VjbHqfpf8aaA4mUhCNQw9p7nl/10Kh3v74xfWDR70ftV9GGtcEtw4
BQ4+ZqyTXjU5heCXJrGiXt9IHeNi7DJXrnsb76SUf0NVAYVgZQibXvxBne4tGt5q/850Gmq5ycNI
nxD43sJZP0wnI+BnFBfkPzhg9CTPAdzV82PARUxIaKa2aq6PfS4RkCT+BANkMGPu/qbbCzDdh81d
ghfIMt9jZ8M1GnyC0JmraEQxKuJ2Bcva6QLC4DVpwfebIU9RxmDkPA3OjeiTt+LnAkgm9ZHcv4ue
PFZa+Vyyt+fr+udQiEsKx4lte7zriqyt2NLYBvNEPi233l7r2zmuCNsajOLKOjvEb4CqyiO7ATIG
GYuRV/2ayanu0N8CrSzFiUKs2Isdmzl4tg1GtHxmrmVVhUrHioszK44O+sgmok+zRoPD5tEnyMXs
FmQn/7HPGMJXQCXhSwHVBYxk374LwEuuGuN62rUu9zo19Wccs2C3e+cmzIt+Iqe1HoWFrif3wmh+
ImEid4KFxDhsjpfK5qQyc3WkUzy8chnU52x/Cg40MBA0lv6X0NNMNoixMnIjqHBF4bgQVv7R919Q
Cf0nmH77Sval5G89Qtf2IsQkWf4F/AT1XjeKxLFrNNhsonJqNp+5mDbTJP+Hl/HQeUWQEwhEfztL
mzzWqCEW2KRO5k+bu22AmDwvk4qMQonk4gDoPi8vTRHvXGE5NhWyCfyCioSAkkq1dvdGWN0z4XaR
QjjifdnqnFvOWA3HDmkV/SGnZyeBzCUz3K6cKOvRkharlM3rUG/wP+uWwErtz0NyMKD2BBNd21N4
iejcfGVANJsmrFKvQFm4mscaoetqq2iNiLZBh0F+UGdu7OlN6/erp5W8bpKXcp5gZGY2nx3fl9Bm
mLQ5ni4fIC+3Not9ETJkPw3cYrgf0iYiqpHltHe7pM8rp2C6i/1YTNKICMKz0vbivINOYhVhDehb
pv9JmdsINaoJpGXSitBrv0uBJyRYjzGW4rITmpfKLIaKViUCO+LOD4QOzSF4IhASwyJU04Wj1FDR
iiy/lt4JFIq14sm5xkhhccp/ha54KzLLUGE+Ad59ON/89pmBKpBqgpKJvJk9p5TWOXrmYDbKZxUt
QQqBDaRVc7Bb4cl7cLGcSZtjjlZpBh/KNn55mx51ejaf6Ks0joGtpkBhg40CUGZgJfJ9hp4ookYS
7lqqxPKXJhJlKVLVPjXGUmsceZlSuIeY4ymnknnqQCJSl+og5FhSZ9vGxPgwANIri4rNXKmzL1Pu
QqBxbnaNaYp0xklxuxKCL9/WT27Fi/po5JRa/6xMqLhICLGX+PgxCnZYN3xmv9HnZPPRv1JNVPge
wCLNTVemFxt133IpB3SYm9aTFtJHxpGxDdllJ7+O6vXyZx6VJESGIl2a/xxvvXOidKs4fx/OcjFn
uye77rrP8dA9G7WbbtGaUhpgm+jOgRo7qUpvtFT+6xPLK9pGIPlOWbIlUAcqRDuYd6VpExt75HX5
T40KJoAKE70P9LbBQZ2qecB0rcMW/0IXolDnW2xRs1w6ojkbsatbR38yYAX6RP6Mkvqe4VR0bqs+
bIf40IuRg2K2Zy8sFvGp/WKUKQnPsZ7rCzBKNPWmwxbo4LD9GPNi9lW1vrkwNf70p2xhXy7jslod
Psk286gHbOk7iWz8fRWi9jGld2AHC4HfzurmO2r0CzgnF5DTMuy0ZcxuUjH4NeohaXwYhDm9m8lY
Y5FQuoBqNYKFgMOmnUe06NdLng95MaEyLE9pYD9VlgBI8CskZmYoUDCnPTJgDtpJJj/6rLJLc7p9
QR8CGdMFi/ulwvLOqQdtQ1jEJz0KvKHB0V04quF1t7vVDH+muW/Nvd1+KZJqWxT8GlIIGMeDZuo+
G0yG21/qQnlZUvwp4AyFOBW2T73Xtig42THcAHctEmbXq/J6xusxIAlAKdfuAIOtQynhC5D1uZ7G
0dLT5yGWlWxh9njzAZqVn9AWFFS5pGrMbMxxyEwIT5Gts9s9UxSrbcz+Pbq+ws4F2JXbgNX8EauZ
f8ErfDZledQmyJN4MAy+UJU50tzXSFuXRTjUQG1VqB79+k+jhOHIP6YVPCq2uQhiTHMY+UTJBUGA
Px4VLXr8g20I+jF0+tooL0E08iHFkaRd9qaj1XMkpCWDOG1IX1Ux0YW7ysB3kxU8hO/EfQYA3qk3
isM20tmGZjTSyY6ZMTlsr12W3Xop57CMYh+3+pjPFhcDohVXg+NQGdKWHwwTnqw2xvDvi1VDUBNI
JJvHEId0jmSyPHCkvO/r84mwoD0YtPh3gcJ8lMLYjk0EWu/qh5DbOvLtM0Ehdp+dGQFFUdDgrtMp
vz+FncUvCozKWc2OS45+kMkDTmUwRGkiARPYBQ4bSE1AwnOeM1CDtTLSHDbaAje5a3RlJJOtbB5N
5O6iI161MXh8QWs6oZVwvkJCwUGwEpSWkWXTy1vJCVCGkh9Zgv2ubkajf6YZgMNffDMr5QtUvULw
NU/onsdefsHgRGIh9S6xeHrpTEWTf2YL+HpORfbTQEENKdhPc5i2MB3bZVikVDkSZFUAikU7LItJ
/BelSdu1njcsPYUnumMonfwyLHnlN+pE+PBNNN3iEERFqMRmRCz8UrRrlgUm8/rpHC+w6c6skgz8
d2/Y6xJCEqDplTvKs5lUiPsc3WJNzC9/Uf/cvr9ctKJ4IDyjYTJwIQ1a+vsavD3sWQWAq/M50+0G
Pyt5aSOlLupAeWjOhzZMQwm6yimvWkXbhKzignbJu9WilX9RzF2yjPjVVX2JiBp87wHxIF3UxcA+
e0ESA53uSh5KZ1UHpVQMDqIB1aIjaczMMBNg25gb0HlfBrfrNjy9PDc8QPOrb9g3JeVHL9rTJQ3o
rEf0XSZ0ok3qFb/xbUlhjhfz7nH/W2Kgdv5ORw+S8zpLQcWN5KxDXJZh1gzEIhyFsO9Q9McYTaUU
uU9s37IOpa5ZZz0BBxLR+gLZyBbxqOwtM5/0so5DsukJuzEL5pzDF3ilrXcij0TDm816TQF22rzx
6uMcsF1tHBDXBfHK+jimOB059MpJQkYYHw1fLzm3qVLUaj7SH4dac9L6SJ4ba06zJ8ZduA39ko7P
iWPiKNCGqprWiDRd+t3f+cd7PpSlPbeTCeQEXl7bnkHN3ivNrzAwkDLoiM7Ji8aKWVHJXtST+LvF
699gWymVjwc3CRqgHtqjtN+zqRPVmZXnHCiAZZKhk626gmkh7OBC+eVd/VduSPVplZzSsnp8pR6R
0JzL2Xsrxg0kGZ70DtF4Xg31GZ75tn2pYwWRifGGgF3M8Zxgbz8/Er/GNISrWC54S0XnOrVXyuRd
QJhkUxbvS6bQLAmCjrfebwVol53x2FMFU290EUd4jgKOTxX9ujKyYqVP8RLW+9ZMj6XFO+oYpItq
pWnga+rWsZQX0H8ReM5PCI5AUjCGYEe2jiNqtaBeSxk2aiJ6TNIfj/wYCQHHIyDxwn+MRygQeSdk
owyKm9ObuooGDRrtsIkU4syCiZL9O3xXAhdU3NC9Pg0TC20aoHihnXJmRdS2ujGJvOMkgpsb/bUS
IiYvAM64eLvQd6MnaVQ6ex2n9AkMQhqd+RsDhFA/LeioSd+y4HtltieE1bW6NZWYQJqUMzsLQ7UL
msSC96UXqNED/VTUuZE0XFbK/E61hzpT7oJLqE6qAyAZqn6OiFZFOy63YzQ7qcV6KHp2etW7W0jV
/sMZ+9KXDNiCTMzImNwKiyaQMeELaoSf5/XdXq5/B/fLRxgHIhxTomZrNimPkTG7bfmSSi4B8sNd
5O+w8QTufsO6820x0IhnJ1EM4DDsWQLpJuS5/ZBsOqMEdaaOs/m+6eahlEoINeHywcmpEDb7LCQX
+nbZMEW+KQbSz9B40v1OXhvyyv27on5gvdzHn/bavEpwVPgDDp9NEFSUDIpY2wJcqInRb7pxL+ev
Zu016aDQXuiXCQ/IzkJSs6R6Jd8yAgaJnPogbsQKYLpWSxdR373PfDYbaKYxdNj5nNf3xNLfZt34
qTuOntc+/yf1QS8osIjcPzfd65hUZOsQJzJBHGV4lhQhAQ42gCfZCb5i+A2KS72re0DykDadtm/e
hF3W6+WzXS+FoJ51Ssv3FnvGhWVx1Z9Pqg7B5RG7p2VAREzpJK72Eisnh12xupyxlQt72ftHnRlY
OkEOz7U0xWGSEjw2EzD/pbcaDnnesBo0AkNqgI+i58zNLxZwWm7dNrPRbLwVnM/mUKHn+eZ0W1K3
U9Hofv8ZGws1elgIBfbL8lTzVurWs8SvSotZI9piodkfF37DOYMoC9yKOuVmkPReWofdUSTK2/e1
xo4qHBS+VlQ5jxQ8ZqW3sxv35MHwMFNRqLtNGyxU3egNNC9Yz31fOMz1EvsLEQaw4ta9jVFoXfSg
qFeMLYcxG6fx3YgkSEtIPxtFzQzHKO4rK4LHW7yGMFWWkZHMg2F0edQvDOfWkXVMmJ5U5spFmwLg
E6+8lxi4n5w2LBf49gzOXs16A7MUaT2O+VXHCUOCI7ik8tr1atpWnA6wJhk5qEw27fNcoe7uSbS7
X7DZLh6R24TKjkPCQLgJmVrs1fUvQY/6QxjAzDnN28MRydeIJhC1Lo++PPRhBLZ+A7ua6beK8Obk
+y+2OTcUiq6Pe80s4JrBVwNP5KlHf8ZMEXUl5U25vAfpf5fAQGk0HXzftgQy5a+7BwNGRbYlx56i
kn/SnT+PRaLVa3Xg0TDN/fTOLWthYo809vy4PcMpTmsWpcfnO6qeiVBlqnRlR9LT3z2G7ucnH/b7
sJTDHruW6gTe2vW7YUqq42IB6ZT647OwYfhAaWmTsCIHNdFoCyGCkq1VNd651uaJHmFXQd/YONWk
D8s7TabCsnXNGT/aaf+djV99eQBCw7p/X34PXvBOnjYbbdivySmKahLGZ8NS3fLp+yeGHo48e0m+
Y5Ms5L6CS33fBv/Aofs2nW/ygzO3/t4UxRj8WdJB8VphbAmfmxxjLAaP/S+x2mktB34ImI5Zffcn
dpKmD/2Boy0E2uGeTBkCwOdjYcTKf+KO+ubHY85jgU3QHPWEnJoJalO3iBVeAGm36bQaJf5FwaMw
Nb2XRmszQY4AEAbSZCK1V7Vbu1++aunMbqxhFfV9BE9PYh8iY29oXYMEn8K/08h/kY7hXiVcUkG2
RdktOj908RxxtnzXSi7gtfkFz2UM7x0zDHh0k7seVm+oIxeLs0gZKiPgoMWDxpiL4LZ0QwE5UDYh
G46E1zPh388ts3N60+z8b5YinukLz4PlvVDQt/7P1k8ivBbvcaI3enKvx+gcC/+o3ivdxHyBHe2o
Gya9DgmbefX71VaE8Gjxz+NPtisFThC5NIvbC+uokHzHyCh+b2OwXmJvDtro1QOP31yQUoet8zAt
NJUt+8YJayyDqtRehFLibRRpuQMgDyn3sfJXCE0Jc9b2IgT4ZsAFtMpZO8zCKiv9gbBPJIrAnwci
kBrLxlwGO/X2qCmmCLqmk4cBF7EJ5rjalPsKcjRuherUEkGnttVTDsz7u1MbWDWJvwNg+GIh9QLQ
w1sy2PBFiFXFODrQn0EzroE4+tbh82uuyXOqpFrdX6/4Tqb3jve4UrPMd2XQnJU3VYElzsrsOCDT
fTazreN8YowPGGeG0BzCBDDiuHMRNRAThzh8TaWCVdScB1xRXYMG2HMzCMsDCGxmoG/PAFh65Mtb
PBnQLGgon97Yeb9aFIw6IoQkEJ14vduCGaJq75PFIV5ZdgJ1Dx3wJ8/XTPCgyMWWhSYvarNBUcCO
uU2G0GgxP6n105T4T2S4J3mNbb27qh2qN6c98BKraNuroDnQDKe0YwuXiPsthofXS7JO3fvd1+nn
LF1ui2xjQvAZQVSG9H3yHt2qpJhWwmVH2/k97YFf4oZ1d7Y0wieEhDWxwxQ59RI604lOi4PMmUgd
YTG8iTnxGgwfHKiF1wuNeSArqH9tEsSgJFnlwis4H/Xn9rN+IQGtHBc5t1bQFSK3LC1NjSBH10le
OzyjfkyyKAt5qpzQL1wzmVr9XXxWozE6zA0hGvWpkW9s5m9oP++AF61vTKTI7+z6wWTD45OwTE3h
k5FxZpsBoHN+7F6V8XHkyG2/jdxafSJwI6IqSW1e/4JTHG6F3K0MTXwln54eoM6lVyyXvipACXgm
zwsSACuEGjonxXBJbTyPl7yF61RwDvX1mvwhetR71SDB87iNtOaqDtHe3CKSQ0BRu4D+AC8T9LyG
iuGKoB3harkf0B0lILIMb4WetpbJiUGQMS3RNQdtV9cy9Dy4B8Tdicsdj3wbqEgygmmFfYdXtyB9
ZhobNhJ40PcY+AYPc1MjOSlyvTw9gppDeHc5++hiokIP+fDTzkl20f60IWsoJ5ZaGttghd+svqW/
gQ14EWHq2ktxCR/SkGG7FiCjMnIMuyf3OpdfefRjsPg//md1QJ/9g9JCb6H0bfCg9PNOYDBTvtWm
6cVj0qYW9DtsWWkz+4wLXYJYUsshkJwXZXsJmt6GAHUyz1LsfontTHuGmhF/Yrs4hLyO8eHw4L8n
Fle9qhL4HTkCLxAPfMotkFhRulMx4P4wNTynyWYIylN3Ea2Q6c0/sHH7judlKa/wZa0V1n8NaHaD
dwOeZ1yjyy2GUZme4nAF7/ttMEE3sHeUEqdxI7Z+qlgmaY4Y8lQFgiP4GgJoO4H4tPaC9JOZi2HJ
2S0xEmC7+YkhuHQJ5IQKfBSSDsIRX608p6ondRG8tSW1uKf7LmRZJ19vKIedkQ93UOB21+9A65nO
tlzOgSn55lNJKaecRRHCd6CQjLJ3H6RyvWXfLagLKhlQGKmaP6hhV+T1Jggo1iXmAH6RGcS5yE2P
yTtteqBNDjyv1ylYHWXan66RuZ4R8Csu6thfySTZZZCS+i/dHXytdZCzgOhbUXWLN99M7mh+Y00J
hUWXIgZLydTkamKGnSR+mmEwGSrhPCVZ3SthLIYS7NvjIrWLyZ1G1WWzypo/TTZBc4/qqu8NknPa
PowDzG3wSwCuC0Ej/nhUTJwrTH5r4kIaS1iuAWRIwvcmUgp7y9Fd07ta6ytF6GjmUKdz01jcPlB0
ohYUjPl1wmUxsQ0vrlSysHBq/G75NNm6p6ru5tNu6OOscoNTwGX+EW20z5OwIQz9DjjUIxEFh9JX
ay8ZSP2+fP0b7/oKifHrkqm6uANFHmolr2qZf9mzuh8xRGoGuLzEEtkz7ueFvE7XwecDmICik0IS
MkKsvE9mSbuXiJhnIn4dLVA/L2FWEAZLh7Xg0qo647dlnE2BSfunF3gA+wRD241DRz7RXTaCsblX
r81af11g6VOYvI3YQROH/E8sGHUVm/qjtgMbG7o763vIqcTJKRcYB+1PyDqPi2zmfcmgJRy8egfk
rj6HfsCxODuYFf293piz3WGJ43SC9yOeOa1/2JqDSXF8jQTye7mAAlDqRTkoDLtesbBIeQmLaxVP
WS3+/zcC/W6GcLyuecjI4XNZUycjlZqivDo2OwEm6Z+eAU9aJMSsRraHt75rBvdnC7HDgMpeW4Gg
IrIyTnnGbrnyCnzBCSn/W+9uorANxc7jaS/NHLZIvNR5KGYN3W7kESU+NlEqUC4gOLEN7a3iangC
5mnv7FhGNMOsZ3iDs/4xjbeyIDUZaX1/AEfZemw/qt9MFQ4he1tn19w4SSjyT+uC/cc3FX3iVSDW
emAHqtIrkkxBWqL34RbxegOooA6PJmU4G/502tuOrPpEzzoX/iLgC+PB5hC9hD0HqkmvkwCUrTnc
X5+nQMfdQYgUYPkeHJm5cZ7x46/o+aq8IeATFR51f7Na50YHvd1wJv9getBfbXFyHRBxwIt1B2z7
bc/ZBpHCO8jg22kedhgTK6npJZX3j8Ustnsg1iHBkRMcjGE3wVAcBxI5O7dAlNNkSd/C1fOe6XuF
kXNhDpQufCoA/BYzh8nwOF+9f6j7ZYW5ojhl0j9+A1M2vaQZrmFRnN6+LsYrbOWVA019I/CWk7qp
LAOu6SdGj4WB1M93mU+Fg97J7eH28E0RuoGryIZOk+d6p2oNTgCz7OfIRn4inw9f8269JoJDDElS
ggz80y9SUTkHq4evha6WNPzjVeKJpCSYUmbgpI9dy9wK8Wobvghnl8TR1TwbY/zTloZFLf9TRMxZ
B+iB0B1Hr5luVrt/J5z72SPcWDMsrtjTKi4PdNvJx0CVmZqPOcOa1vO2XWcBOpmenBQbsA6OS+pS
octCpb9aPvawHTEo94qxmdNObYsDbl8TzqfU07LxEN7RncAk10i2nIHf370iU56xxY3fsFPkNXQp
EqT2vNppuB/YYuX21GI7Ht0nh5DyeBQcjmnvdE30ksh0VW/L5d1nrARO2ApYjCm9FYGt6zKKChWw
TuD/QeaqdgF18uZ+QCDyzNRnTSc9k4RR9mCqQ2yUMz+DVObaTtqTnFez3Kv+3zkbZjru469DSPP9
qN4FMckd+zBR7QZRV93zQL4WuIvUorSC385BLZL8alEtiYKeOpxDZx8e0YWm/ylVaOSg4z27MZdL
Nk3tdldCPmZ7rP1mtHAg/oHMfCwtBtw9oW1wB43mHTQLkYTj4Kx8Q7KAn6Lawi+g1jr1Ancf4YVe
tCmVlr9A4wcLSfy4FX3rp+ah+7ybOUOKfu1+1KefqWZsdL1eJX9RzxOYbP1IzIUs9hKevPcAOkyq
QD2xVuzHG3e30MbF+33U4x9NvlSLPFikKtXRHHs6lotzNcg726QUmtSWAlhaePTI39iAz15yNOiY
SyAy5LfaIm7hH8fiA09A+RnvdIauiX49NfAe4o3fJCPTYC1KAvmwCHhIZg/P96osR5o9B2f/nhiz
Sr22/y24sPCMPcKdcnuoylHsk1VWlkD/DSIzGwmUdjULPBc0dBnNE2OpZqlylSnPWpPH7iw84t4Q
oeH1cLF5ftwLN4G1WXX67rxH8LaKeBxyFDZLqxCirBwMOPpRAVLh5wrYPnag/2f1G0U1BKRnzxlq
Ezdsm7ULWX4L/ve3z/T81TOvZ1EJVhYHY7YT/OUMrCoUNyz3hvCFCyhGFvIIekx2VephYBk6myXE
m2Ldr5W7eI0yT88y/R51iPDTpGT3s4RJp5FXEQpFusJFe+Us0YTUj1aTfehTLZRq1htfr449ihU2
G8RCtZfIIP6cg66jOvDSwUVlYn4DtcWW5j9bF9vo3/KGyE0JfcKKA+u4kX15+Y9Ag5ztCrISFMK+
aqs3zHPLdXijVBst7qq2gFoQaaEc2d9HoyhqXFGF9tizlGLStscoFEEBRN5sAuHWMWJ2jGF2VXhU
PbPLlvtmJeHpMReyEw2IhnJITk6oviHM3orKOlwrFPfG867hLgoknqPYtPixtO9q+rFVkU5MhN3Q
945IoeHV4BU+Y2/WgczX3PeS8jE9JtJEZrgXQ4mrcYOjG0+aq7e5VPpeeCtFWswG8NNSvl3zpYR/
iygkU96sWOItVkAlkdE1rw5qa0jiTz3lySQQZG7tBBLGi45x1JBwFvEpGM6mbi6szki8DUfC+YA6
7wqyTC85JI0LLWU0A0d9/eb4y//JaJkn9qEaamZPN2gWE13N7HRSgQZtc5B8TYMEbcuoYEve3pOt
mWs+4+Fwsq7YZjZp4bKFok+LelpArIZI8yQz+w9X66m6sArbbAzf7mJSJgTB9NOgwuwHW2NU6Rrw
dAxk2U8xX62TrBRcGPzys/xA7JMxhPKjvkLzWnMszrzbVDJ+MEzfY43IePyWPSuSBrKQ6nYF9XL0
gZ29lTaZsvLqaZEJOXeRaOcpcpnC4nU/O2NEkX8Dg+U2nRCRwzZn/RgO2UBxIUjT1E/AjokN7YvI
csRg+kuTJwNV9h7gjRDgH4Nl0Mfwq0jg0HbDPO10WT09QJJQ9qvDlZJZ
`pragma protect end_protected

// 
