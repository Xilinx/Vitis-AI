/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHIWq7G7ldgNzxGYNsmaBfcIDRMzyCGWhxIB4pjie7S4WTA74C/XTGVupG
aGKaHtQTrnMivNKlR5Ud+FHKnTrNwdtd0gdNaoItOyYuTJPKS7W/8nEOCOhG6RmMySfe+H5mgkJF
oR28hZ3ZMxw2ba5KVtstpErLzy1lRh0PSKCIaHheu6FcOPQEzCiWylju/+4+gGhcuokcVsWf96Uz
y1t+rVIEP/5vafp0JrAJmEv/8rmH+CEC1PQaIS8BnIeXjYS4ja+7wSbVC0xMqUQoXWZtrQPFx5ai
6ZqagQkT+RbqrSZbQaAYOrWDYbdg1yxkaN0psQw4VuV36IBLFXCz17QOg+la0USO5gdY34J0AOFG
bssv6JafZJb+xsp842nbRiF1rEganA67m7V/n4cJFihZNxiODDflg6cCNr62pVqCd8K6MTaJVCk8
xPpL9EdN7B6YKGAoILbOmbVoToCp7vfIZx30AXrLnCKyzOwToYKL7x332wnDjQbr3eC56Ts94fB0
+0UUa8tCcVqps99iEGNKcfhjZ3KF7dJvxKHQaMBME8aSrJZD4qONDwdd0W22s68V7AqtT3GkPFrl
Yc1jo8tExXtVNpAcMCoyaa6AvKyD+06O1kvwikKXtRyC/vGs7ig3xzsSv8RDMQ8jz3dJHLgGygoc
A0lbVdbzUY9shBl749TVJAzKztvROFUril0EL3QmVmNoGxKxV76TPvIIrB3QHikNS6Y5i1QlIcUX
CyPoNqIQcMLyE0PmAb7TMvOqmKGAffkPDI8LWT8IUxM5mxG345P2bNhSwZfJlT44fIZPLvpW6Klb
Z/AAQ6kDh75o38VVdmTvVVkrldn9+ThPD19Yz97rax8ofDSe3plIgJXb9z5yl6H2Zwk3AFVwoLRQ
u3YcJg7qDGcSmejuyBQADAIvrkQGpBLkZpROhJIIOFBqn0RNMWbA0fQY99Ke6+fS5z+5yAdhvF+Z
ARc7DxCWFFsc++bZzDR3Zv4sq6UuBsdGDimQOPke3B3OwvRVODIevPcHnDXNoAChGrpfqyKtUl/E
pfjJNGkf/NuiZTJ3MEPo3VI/mN2AgjoBm1PgGN6OkbWY5VERj45IMYbPw16g+Q4ythRAATAbOxBp
5qc6r5+jHLcnYlNxlPE4+RWB0LEaoeObo/sivdfeBR6XACUU4AqcbTbX06sDxMO7PYkZgtH6HsT1
3G1p2yDg9uQdXL7V/43Shxk1ghU4QekJnIWdn4sINyWN/iYcr+Hdjlj/HMCat7MMYivCgd/pp5j9
RDHFjoiGTJxbiPvkOn16HAtKm921qYdWaZE8KpEQh08MnqaRek8mdoabo2HX0YWTGKLBHJ3JqHjL
0TFffGCNflK6fQrmL11Nen59xmAggXpt/Q8sP4ppunkoGpONSYZYzelfjpFHs7nI48QOXgghVE4m
fDUeEIk=
`pragma protect end_protected

// 
