/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5856)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzHvoIuThoxt7ci09zimA/Smdcz08RrMZ7DQjgCnTxMY83ubh/H+HZnGB
ANSMoQdg9NOTYOh7KcVTcEtSTS4mg6Rd8GuVPy/bDrqZdRbRnlwCQD3RHE6g2cT5HZgWIe+cl07E
pMVwESm6QkNIJzGuPYsMYNSZhpoa0o+47S1JIGYnEiZwwfGGC3LUIVgHEm1yHt7Z7bUMK9Jtm7qp
i2GzM1KRr+vBPYAQK9MnSC5D5z26fgjl98Y50BGUn/BWV1LPHRUpt79I5H0l2/oXxBWKqdH9Pc9Y
xWSG/xpwNAWaIb2UCHSfgvGQ5nM5cSi9S9lR3GREWwsyqzsvgc7KD9sm7SgloBMIXLKZycfm+s+f
z7bLP4lYGezli94d37ulWXYniuR/ubfPYgEF+cXJtQBsLjCvJ6vAHDkvUtDUsv4BntWLIvHxzSI4
k1eqXC7VMdNW6HD4Do7mxDSCvHOtqGmS6SEiemePGzohOcA2i2Ow1Ujo20WAgmbW+Ai8/NVu1UII
pFjLJzWSulO4/ARg2VPe/xW/sQLCzq4faomnyi3mw2FPrF6UczSFqCRNm2BYAyALFW/StxfRTL4X
e6L8MkTNB+/1cDoI+q671LivrWlvO5Rz7Sj/oZ2w2qP+QBd1sh/y4q9UqsQkl0Q38/BkSZOkVN9I
vV1zPMpH45QqC6SgCSNQZuP2J8KZunv93Ja5evop4bMvvmTQvINy0pYlHTE1wElqrPkqoqQuziAU
WOZo+qDXLT+3Hm6NBYtODiTjfZhhr4zc466xHR/4mwDR3kXx14mIB1hueZS6wQinV7Km3nj1MhVz
CcsZ5CAdnsYgxGfSjKLTUkChLSMakqeyapdm+oBTj7jo5OkHDi1njxDltAHfoUUwYPnR5Dg260T0
bNjYztuzFiDxaeYBnhs0Xp+y9+zkQRM3xcaF4jeXCrSjE945r0+jzh4AM6jblpyXyKct2wRW36Kf
sb3fkXo9y6stuplGqRe5Xm2ExKAdHwQjc9qbXDPkNzCogjkbtv2P7yfj/7iZ7A3bMUcSskK/ZGLD
3ty2TW1QOdUmHj/NmsmlbQ2C58FlgRtSwz0px88MiDEmAj9GeHxhh3YQoxOr2P2DfRnlKAwn0YNI
1OU8uxmo3iGsdSjzRgRfjPrr098eNRa2C3nb91wVJMHYK8N4jVDOnPOaBBccSorEB3zO22qw3Ap4
AnHz8B3UchSCMROJjxuCdD875uEwFrrlwdS6OiIcYsnhNotYtVvhH+ZX590NiRpnRZ1TAyvLjXte
iRS8aUqBDqN/Tae/jnfSgRvhTWyXWfG6/41/0Zs9anOTTrVzFnQ+Xyzk0lkBpWX8LYF21MRql/6y
ajxIdw77K89/Rzq+SDnNe2SFkEr59SLoszuaoClmyefKdjp2C3cCtJw4b4zNHjWmZjerg3fYv/YM
IGxGJVPWNTtwqbzL6biBak639DW6XsGwAtkjr0B4p65rMQmzItIQsPcpOTRiqE/fdT/F3wMMJu2t
8rzai+WiXsWOfW7LZa6PB9y9Y5R61EuBMIEJFczQq/OaHF4brU1Raz8oihLgOAbPL3Ctwthg/3Nj
l1xcw5e0XxyI+N8UA15KYNydxVy1lLBsUjKxhdoq7mCsmDMHGikbXoa14H/3iWzgK6UvN9mwzHEa
OklxyuS+OlGWxGPbLYmBCW2Lxsgt0oUd0QFJXsyqZe5PddA0r5lxQ/y3Ske/+82G08izDiQKuoca
ZthRDiEgcHwOHsh3baikBXffOTBQoX1lNzA1dp3w/+60vid8iE8h1YOzUUr8kNUs3x2NKmE+dIL0
5MPdGgzJonItT+Yb6SeNUZLN3a5k/dLarc6DcMHjCZbdCkIA7l+5XJDmrTkd1WKbYE6atZmiO+My
KNvDKdGwYsL+Lc8uv1C0YcMydnXDhPhQ3X1mXeWbxFTf0xhuNjukowkaIQ6VTib0iHrhjwDZ9+lB
qSyMSUoVG81dijxm80VH24ZNH0ucTGnUJ+6LfpZc+zLVt6FurwmZoq4u7f+HKBbZebgYtxfa2osm
USxZUpgdQuEYBRPQ12X5QPKVlz2SvWvcINupOYtAT+o2x7AMUwtbVODP1hccSe+nuvSOe5+Eqgz2
IBOK1UoNcEesiZzZg8AEzrbEJCL1KQSmfi47xU61FDgJNaThWs+FlzX35YIX0Rv0RknN4O0FfSf+
JVxDJqn2qF5H7VDf4YXH3WPQAA0547dvZT7HVb1OydmCiobiejgriNgo+jEPhfUxmeYCkHRc7nSJ
eMQ1rsgcfcmoC9UxqimaahGmUEozMUFBH/uA5rhVFBvEHu1iPEe/cxWQ2sgfEZ04QoBJKw/QVKJL
x/HeznnsNluIvxkwYIlkLHHjCoGLbR0Y1wd4zS4yIyaTt+XU1OW3yjsTTYEJhC7teGUOpk6LeqsD
Ix+RMjdG7QQjuLDUYCqZbQvuxa2WKdXg1fjIiVABk6pZ3ogD8UoucmoRtz32PIOWxqAOxds8QVLA
AaXeC/usC9TES/WEq2yX+82usw9Nj/4uJ1TLYM+xx6dKmMb571XJ66KXEPwbkhUDcqNg37GSuqUS
Yp6QdCRSss3FZ7c3y0vkICc6g5mDvNLBfsqapVhOt3ix5ejp5E8WaPlVnfeGfv5uoe+IVDkNKDQ8
I3t87qjmFeA1P4a2B6L8veOQJPSXZ2EwX/5Chqsskm/oPc5/AYgTKe8/f6S9d3H7ERXGXCgzB/gB
BTCVc5nQACKflu3KL9Uaib+c+GlCm1TTtwNx45QmmVM9buj3tnO/5LKa3CfMmVwjfCofD/38URps
FUAIvNDZCzBE3rYg66YemGGzGAlljBBwnVLuoz6LoyswEdsRh8EIIafRLLUbxdX/Ix9hKm3v+RXe
f699z1xNtZ6KlBVO/u+kLZrOOhJRpgZaT23mmsSXwWvGxK+wU0EcGzwK7Plfpzk27SY1cwfdpAVJ
+Gf5b6ru6KQArmyW92b/TmKS21LHD8/zP/6dv8jzWg9oDJx95povQpOL17Pw69sO5Kh2lQ9mCofS
Sy9e5VM3qZVcKT3ghtNkG7/XVvBHCnvviG45FRThVZzQ1jSbuSuSYSstqfer9nzVHyBMx7Tbz4Id
WiYgj+yX6VZbwN6DwI8Xm57KkqtXV03c/eepy7OsXfwSI28mzP/VGQkDTDJ4WJhdcBsSm+Y1YdRw
O1asN9pUqXLEi4abX27lNdGBfM+D7dznczC6wYrOJCRGw0ieaM4jIRdV6KLbs8/jyjgMqG4GD4PI
WYG7QoqvY3Ut68fpzxD1QXOTjrvk9876uhrkfm3EI1UeZ1DA78ADesB4cVYiZezR2vNUdwWGVepv
YHMY5/QTTuqJEDsg6qwxXVC+om3GCvQ31TbawAiAtFO3byj23vmh52GUt9xAFYv4mJFmoGI6XQ4S
Zz/EpXlGynox8oCHfAZgAX9yEy3FzErDMhg0iAyW8HtQYbMaTaJ2Ln9wAS4c1/iMOKCMPj1oR/5D
amVxllF+aoZRJQE4gvWqsC3Tf0SF/MPsNIbwEg8bHMaGfKV6HJYwFqE/pKBDq8CFZ7HfzqtpISBh
twzCOo1aaOvfSwYUCwwjy3QrC1jnmaqHyxN+CyFrKa2/uI8Hy7kdwVA9RQ/vMmimUXXY1PKs/xEQ
Xi/OIWhSReEQ9jeMrPr+8uKDn04ANmUuS3moc/n/6HE73dH7qO368f3u7A5pfuV0dn0JvDBl2O79
7jyzHkP6K4jGWh9nGHXEdUh231BP0RZzGjEw3Dr+cKurdQss7F0x3RoMva2pPmGQ9wyy4Njq7Jzc
fi/PNBNejUbsuWaAOAXkjWdLqgX6o5Jz0eLCvFKjP3EXvgp9XEYbQMTx85osPwOR91hETATS5gzp
UsN639G7IIqVjZpcCv5DrIS5gkU7yT5Gv3PK3VuxSgiQiUlcSsOiBGR1QfexFfRHJxiTQPxtBlsJ
WurhGet1+bLbfNSGJ2MpyUlQ56IxwvyTRZ9y7jK8k8iP0A6FMOrCE/hvJqLJd31SnRWLn/8rCShG
CfeqM4BKKKC2oS7H+C5Yddsfwb/IxkgOKWZFCWmzCmYT3LEhnG7n2HXVYt7lXNiqtSdxLJX6TAun
+Fw2IITdHEJVlunncHjiHfRe8K5NPNnJdSr/lLM7/IBijDUKY2gBDeANGRVU2QGJk/iDee1RRfKT
kanXI1hNTNss3r9+eMTVQoEXmdNbw7fAU4qy60jt/uksyNUq06pZPwkY+vgsMNauqp81dRV7b8Cf
IPQ3fITVtepEQ+TNqwuBYRJUvxkKjSbhYMZovjLFpZLpLFHb2HF89gXsWtTGfQuRIXBw/12MRtAB
8hwhZTPMjFnP+Mcgjo/hfrRZKoJiLpTFWStpHT0lhFDbALUrHspEtjMet9/fNyvAX6Jrakeryl9Y
RY7OT8uzXj9SOql91F3MZ0J3cPBOEM77pAuP1GX+B2vYGaYlbKA7Z4RwwBA09O4AjpCMj/Np6p9q
ntFVa97lUCyJ0ds7bcqYYAoH6ZI7/rD68sWglPQwShABESRhrIHK97+Ec1YBXB5yDczFASBtWBTH
JSW5tLPnLadeVj3hyEkS8Cmp/7+b5iHBKCPcwP7lmktM6GIAZ3pMPSpvrYdZEP9/94srlVsrr+LV
3FSJNWpjT8xADo2a1QfZUgDkp9brcYv4ihhd3YYyN9wLjtm/6KNzvqdOdecZUeD/IOjzOMoeDRBD
dFQ58/w5PVUpIAlCBdExyGf4ekkfL5VXanLGgGLzewqYyLjmSq2n50wauMGno2PD+7d0LDm5Aby6
z98Eh3FOzmu8MBsKhxzTAZfUcIUW0OgDBGB3F9DtxiQL74xbqJia8jjhdZGUX3AX3DGjFk8iM9Nv
oOIiYnsMLkBR3OIxs3GeHPGprUX4LPJl41k29vlXWQ11WaTwvAxlrC+rtpSqqSgOz1cICt0l+A0a
OpDVvdWTsQpFb6ahNHL045eUj8NGuEzSFqHggEZqSHSHSBzi1I9dekNgIdrPvhWWSPioVjweOIug
rDerYlYf92+jgQWkoLAxoRA2HpGDMVNE0FkrlOnt8mKgQKLNilvCffnaxc2NhHuR2AKD9XXCMvn+
gEGafrMMGYrs8qW8c6nZXI+pJxEjhP9ywcx6n4YOPIlvWy3A/bP6oRqdEohWEVgyJ6V9IECuJ/5J
eL0Gs5jjLY/FROX665+lMRNEOoVxR8SvCTaOJexqYjqWozZq1peNdd+ESgoEsKWY7EsogBrLpgnp
pvUQrb+GqORSZzYXpsiPhMTwmyFCoyg1JMHLdMMg73uOVK1/m72EALFtyYG7Loz2gEGQTL9BxosD
zPSph8sDDMz1/bvDsOtxvjtzyV72trEkueTGIM4QeKO+Tuklu+zvcg2BbN8poB+vXwYKXEvLiJ5B
aza2TWQQ33g3ZhmyMCuYpskoy5348ma9/HvR6AnFjYS8Vzi6l3zMJ71iuozFLQywOIKshheMbsjB
0x/xd8dy0jLarXByTa0+f3Bkoo7yedJ73vxjyZ9oUXxB/SVRb/OvG+CB7hfsy6BoGVL/togl9ulW
LADBoh4BbDAGX2vVP7aLY+ejtd9tuxpOLfHeqalo0+ksWeZkk0u+i1jQarygEi0xfNxCcdJujsHu
uy2BpGgg41UYTjkbQ/8eBNaSYusKIJPWFoWUVLDYw/jljse7YAy91NYcSzqEHkCrgdBX7vnWVEDS
+pu+3XXgJYVJiF85WbvKdxhgVEYOO9MyLzijsZZ+Z4EJsgbMAxhLHbgp9ZGj9p5VV3ifrt2m0omw
qHx01W9rqlAEHhLJcpbU3+U5O+tuUMAyccG7p41OROEh1V1laka01VrF7DlHvqH3meCr+I82b6ez
mFjI3pRo+5NUE6dHlRzEikMeg/ZM4qgq0lAitT5WC3Q9lQET8zS9VhbhsQBLwIrsp0YXU95fTu8l
Tawd1u+B0yCAeusKC5Jq88tCt8JhcP8+hCXDvDKoXpnfsJTBH2O9I3Kc8BwxUyjs4w/aoTemWFAj
odNg9h4V4b7Q1pJQAxm6Glu0Y5lYMtENQl/heEY7zvgblB4Wv+SlAg7TcU70vwxuq0h6U+JaGSuw
nqlsf2kYYqJXwKRc3HTcVE81fgZ57++yeOxVWm75FNLs42/1KOhSO4PnYlWdWW6YKYOsAYEhftty
NUJGm+3kROlxPPcifqwiort5A52qFxoCSQvmIU/JI8XxQZF/0VrubAlJKohbawxi2B1lCvHlvVPg
k1/QhM5UYVguflDg4kLTPMYK5GXZuGAhqoyTH5jpoJrZfauJcJfr29ii2zQA2K/vZvTuIAgMXw0I
b3kp9HGJXwCphsUnvtgT/VAPeTMoMhS6oDCpv21xw71P2xLD+f0AZbcqzmaCdQoB32aNh2+ODQc1
WPIaS0wLsHI9rH7uaOfp+cxa+wh53KzeR/8ETtAUBQHUvHx6+9sHv6KfBW3vol5slnfAn1F4Ca+t
+EBFFTONf0vTYjYrTYl5UJvfBM/dRLEJ8YGYnmjHIcSfVY7+IYO1StsuXWQtOyGggzpGjP6M0YYf
jFUGClEeIofypFxs0AA4aigCqZvImfDE4Zy59Ljhv6ym63VGdXrLFPtreWjEKtMz+GGKpdBYi6EN
G3z0xIqMOjS2k/xQ4PD9Rk8a02b6cPMKqFYbLs6vr1AqhBzCX9gOtrDosjdK+ba+hg9N3nXgMAdr
s8TA+gofaUmBQXvq3DTqTGbj3G8tEI4AST7ea3C1hhWJFOBqRK0z9NBlZZzZyPeEnD1/XgH5WLiW
Lug8+1q2vyOQQjUY8w5EufFn+6JUg/ABiqPgbvilkjUk58f1oV0wUT4zsg3ZFctRtMk2E/cfdV9C
RZsMI16Lji1B9txxIrbtX8j44ZoEfRgX2IkNVLW4i7aoIsNbB3UcJx6bL1vwkj7W/s2re3s0G++8
6LhKRDj1BTpsYPhCiUbMLRpAqNvgIP2h9kxDf34n39omy9qRGx57zOFwgHTdzJUwImobDy3qM7TR
SiiE4TY1nOiFP0OkXNxycpVFKgSwoTZPkwKrmHjUdvJ1eVbZoPBvmxDeypc4pa7o1CaiyyK7fKnv
gCohVylyQjlqvi6mL8rKT2a08FZXsYZME0FvUxskuRP3uSlc92jgu/WwA3hKj0tQM4ApKMedCMS/
8iTRXd7oRD/Q0bBayRI+Wuz2/sfcJ+RRoI9UguzyEoJQOEXV1BdjfbLIiPuYll+ToU32UsA2MJnp
FgefzmvJ3yTUj4qwdyOAlJ0zAYjMY1YsfiryRPYev1Q8wRfHzQ8rD8BFiQIGIBUU5Dyb/4jgS3d2
yhHktryJCM5Wet7X8ONTLdtUi5qEtqWy+cfMXaz7Q/GijIpsMgN2d+rN4CCyIVeJOjsgMP+F4wJA
IUyBNwQBzTSK4xXaqn+BhL5+rRogSKarLO5+Nz9mZlyOJxNSEWGKgoI09RUrm4V9t9Q6fyyD86fj
JAJW6CdQ3LdvuGz0Bilhis4t0uQgVBrA/wHo7RwYRZzfvgUhFprtoo7wKrbHDbjezszkCfN3KM08
Pk90sWsGOP4CqQMbTo/8O1RIpQbZI1Z77AdX2CvBzYpdwnJVWIkpqtEucmqR3ZGmOKGbsT6qqjAj
2MYRc4+gpHlRYMjDIh47gb6rdvPzPjAeAI1hrZA/RhGeBLx68Y5/U6PZpVf9b7aYzoTGJeQ4LMLp
2/WT9q5zlJF8NYvI6XUzUyR2WAHNtVe+mBVc77O4Y3PNtjUNFVXvKm0A/MYWYB8npE3TcM6M+cEe
eQtU1swN5tzKa90+dA8oQa0pj2LhHY+o1xFmE3p5kg2Aq6CwJ0iXN6Uo
`pragma protect end_protected

// 
