`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF7fMQcBGmeujuf1kcotL62DWZ7SsX/+8UkBoWYbos2hFB/4X0vetVDRX
19SdCyw/eqZ2yaiO+szdb0hRz+stj/FMI+QtcSho6WKnetFwhyvL5yPAY9AU2csZuigrxnPq9qQ6
oT8k9H2i4kynNH3YQvzGcaOKO4LsJGn1uCM4cBI3hpOYRlcrhFiDxLy76NfdyzxSTs/Q9X4LKCIm
5PHpjda74xyDLmfaGqnekgfNCqlmiSRAPEfJojMBmpLU+37yC7RvQ7qFq8U9lm0Z0Jb2UU7ZriDb
JRWUusBC2Et2sQGq4Ekdb+uxcP1NdkkOtC9xBGItfNy2wg+NqhE5fLNNkFqrLND3w1ZSpXoGFhBX
9njVORCtyU2i68Ogrq0xmS1uufBquoa7Gi68O1wc8A3bdEZ9zRL6sU9IhS6pFoJ8z4PwO4ATdezr
r3Xrp9zokHf9CFc4xG+fRX14x/fVMbfJE1UAsKiurytfyEqj6jdexGZpwzqlNRUD5SgMcgDD8bZb
aWKYEOnCFnEpregufg9cO1Iyz9iJKRu8JUO0mx5J7DrBd12oKBgDz06nsPfy/YimuPLNNhqHxTEr
GxHaxF+XGuu84Y6FOXoHc1jp1TmnvhdDhH1aqpZXg9ahtJfq64Z9Q1AIbbBxX5i8yiJwOaHt0r6a
N6fpzxsVRovFfWaWKJ63jjtXYbgZU6Erm0ouTcS9rRHWO1tIOJYyYDhJC+8fl3go/A/SZ0LQs9Vs
9DjPN89dHoYLlW9cZ6GGKHWFz5wmenXNY+VuzdYIzG1jziiXhU9Ikyl+pLUYTDoqx4ee4xb3SPDi
5NniHiFOSY7enhMRKoTSqs8RV8RiwIIqFwDOsBDldCXilBPt6nc3Oz74GlYXp5LrHi32+tCI/bTi
nFYBozM2r1nUQpeae07pGVEbN09FkKB2awSGpISLPRwIkI5AurNmhK84ngvH9zHu2uDjG/lKpCkY
4RAs/HNonkcMmlulfbnzlP5FCNk8i6Jfj3S02QnkCwo9Gdi4yL5/lGUgLHRxeNoSni4d/cIY0VED
xyxyakiBIvUkDvVblfA/WficAcFFyaYHlmUIbuS693rnPjHhLdidb6DYoHWzvcV2b60qohMcnBtZ
5DDAfl9V4hM5lj3ZSdhLIsB2/GvJsXN3yt4JQphX3VnyZh6UsMl1Fbj3FvpJIwqmsqinE6KDidtR
vnR1pdows+nM6lc4xLgMBdsP/Q2KaK/RGJZgaRcrdSgfQjudBmR1JsDfdGghI1LGpqI1FDEX6Ddz
7Q0eVTv6ubx2Ho5a82K81q7eRESUsPupBvpL1+thmGk4rYEtqqQ9Fiw1UO2CVsuhZ2bWG7nbC9Dd
Sqd9p+VbdnADCvWIJjQN9q8MJhZ9Mh70i0z2YezFkBNuL6nDQhPpDZM0by17nz5q+DqXmLsNtrxa
y2ki1rleh2vjUOvdkD3dSctcmO5wCay2UfzdLDxhFRzaplCSAbFz/eZIGhDmuBXJlpPDzo4nJIH4
RffnrDbN3q5uMTwXm9cpeE4nrQqLMWZxT+UNJvWQNalaR/ZY9bxAlKoduUGJK2+9zSeU9Om6HSDO
2i/XNxG4KPDxeBTS+wjWg5t+oOmilj90+aoIiSUpTvkQkKl3Zp6+U2ox52R6ktkTcN3dzsbCjQLo
yfXAUL/sdfmtRD9QyFPtSsDkob4YPpHvZeNLDSU6K6d8uA6TsSiIvurBPl7+YuOoyNkfLdIZeM+w
MvjRhVrqPScF/jOC6MC7blEIRQT6Op8tv0ibSgvzjwTua11B7oxuEm304AWKMp+z27riAn0wbPYU
d0KPaiMHdz3OBS2NuLxuuAC8o/NGWEOMuPSAPeSj1mzSIwlJH3x9htZw7Gl3r0fPByD3t4y4yd2i
iq29nI3vz/KchHJVog6aDlBdjDXQ0AiG7hEAiwOCtVioOs2iIjmBjYR2+rUEXkzG3DR6JhJ2Rpae
Xs3eN0P61s17kPSCFvevNZEyP4yoLKFQz3BCMlttyUztcgSzcWTv6Hg5p0/3YeWmuqQRSwuh/nY/
C370GYDaxIQG/WfvZdXCQh5+ih2IrbZKqLNvZIhLGoxDlkKYUWvs8c0ebHW7bqy/2AA126Orvd1T
aHWq+vcSAGKhVfLWartJe9geLSOmD8ff6BQPnP6vgbKMCM/nbtw1etBY/ftq2aqmAnrreLvGqobe
F3WnWqdEyW2e2u7R+y2CGKa2HVHix1jsjMHaDVWgyOq3Glnz+7wKMVyEbLReQQ+KAXeAMVEEaR1Z
EA9ly085920uyYANKi/XUV+8fzRT6AUNYrFh2lKXqzkU/xAeKVkUf93J8j3oETH1OKLKXUugHtZ1
OHWe6j9ZqF9wRGnLNSYp3Tn1OiL2Q8P1GJnUR9BTJy8Shh9DZHdoiDrMUAFgqvkkIB5zZkgnZKlG
bm/SXNS/lMpUNCJlpp7TtAbMMEp+3ggeeSE00LrGex6N7768og9nL6L79pGJtMtKCVo+O0pYz2l5
B/UOm//oQwVYOKgB2w1WMCFZ1T1ysO9MxYDr+gNIxPooyjNeE7qUg3/fD82FXsU+LFVTd5JaQY7o
L5mRnEVgBH2NB3vuAsa/rhUK6OorZ/HU4VKkqWQyV23EQNqzzi8ccI4Wzrhbp9NllZyd3tyVlgJT
BLnu7Aj6/jHTiQPNMKn7QSLZ0yCpAi+WFgeckFPj/kHWRY2n02Rd4MWfsVcaid0esBHRAUXSA/+R
Dot4F4wlTE4pi/5EadlCOFoavTyyIMTZxTJ1orE9F+b1TTL3vLW10UPtn5vt98Sp0bNcmhtSLUl6
+L8Bit5ewb//0oG/Bpg0gdGShLJWq+LGjFzplQwf7YOyge0D1cF4WxeV27DzRNNaVSPMuTITIxFY
WzSC+IAVE3X8vWXNZRiBYJmoScky7bEmHXBSwisFr0GrljEK/Uy3fGqlM8T+xl2hgU3dkkJ/omAR
iTcdQBeBmRJq7qnOuZSCl1SNCvgB5rO/ciWIcTIljZUxJGYwg4lA/RQVFlNxVgARlKqxcJJByNJv
t5+GpaOalDatAH053GRilYYziphKaWbEuTNuezxczDX8qJlc6PDD848MAE0dFeKysDAMXvuCsLxN
Mu3nBgG7XYR36ynOGgyLugDhUo+Z0/pDqrum+SPuJL4Vcq3XyfWKVX0cSoR/t9e7fLTUOfVc447e
2vUPFGdrjRyQsSwKFVU+Q+DwX1D/HLRpmCwy/vZdPGuAqyOIolDsBTqbZpS+sTMJQVT/A2DFGjwD
VRa+pZpE7NltXbPKKUNC95mwW8fkWCmcResNpBATYCANKHR7jFpyHCrxnBvGOniVSbOJkregAW0+
m0nFfZK/heoo3ja2oB2ExqxA4N8VxU0D7BwT4j7xd2swTuj/tqnTVBDgKs2UbTCL3+Cjs+pC2FHy
RiP2YUZgIoTv4B6li+RCzAC8m1fAirmWXr7w/MNf/pKQAeBwKPB+dkLWfRBfRpi7SEbKJQZC0jIj
H3TZQZRi3p97HT32UtnMIWQHR8I3kv7oD8VNT7HaVqOPG3dxrPX1oY8nNkreMR0fTcplTK9O4FjL
2jQwQ4yOdkA3KVQQCJLLpWBKSgSdai7W3KvUuMDtpJa/kEo+jgRxZIJdetRLIYs9MV0PZOmpiYHJ
7EtmHuQwAU58Grcighzf9J0WoiGyCO7uHhDIxhAMrdIs6YFv5kcN8DWTk7Gmds5m6Bua9UX7oOGt
Ku+yM3BGE2ElgLm7sZPutKt3bk8y7SrfQ79T3WH77Jz8re02beiyKPKC7ieUSjl3GOs0lWqeZbIx
Ugu8VodsRfJoNqWcPvCAIvxSfsrcNyRzb8JkvSR+C9kzYCF/y+1Qte3YxgkWMM7lijC7B0G867ns
8wRlWo7HTxzWWFlmGVNPNKvRph+FlKSLmfb9mpEIo4X1OBH+PxkfQF9NFrpjN/FLgx2TH8mad1uT
hGFNoK2L2JTz4olBSZcAo5K94BQpzWpu94SWkwOr2A8KahSmuTJ97i1husQXKIPnBJmxNiS4xHQO
aSr0rK/j89x9q7b+Ea2kT5sGw0VykEGTF3MzKvHXimjkyn8+lxBPKV5ZXF0aVlXZAGKWmShSWwF2
wur6tOTYxkNS1WHspJxNY3vLcN1vYeZl/AugtVqtLIt3fUIGIpFhYdKrTfVH4NsxywTf9ztxUvfq
uao8ixsSEyZaiyfhsvFuEJwuzjoWTbQakU1ES1lr6D0VFu+X1FNVEndtKlAO1ZyKhN1H2BGs5pEF
HNLvt1EuzLZmypsque6CfH2NTHtCxyAra34mlH2xj0LhiJ8YMJgikzLjZq6gsH2EJnRdmid3weLh
VSDKq637c2feoQKpvrSjBi8e4+BgkpDebzPvFOvLj2xit4TM4h4c1D4ZVSPgloH/G110IOmTh4w4
Il+Uu8JgJubXuGDRkvLUXUvoW3COO5GLm4g5ZzawNbv8XLmuvcBR7pUsc8b+MKhG5yIemANks4K2
e5wZSrw3u4tL69KdbYj3chJY5pY6dlVTfxVGAwS/AYJXttsq1Kn3ZMrR8SD+YaRLVNf3JB1qvNAV
tygug+AcO0CDQr1i0b03FRG04aYILX8BppRjsoyC1Nkal9JONpg3bEuyGeqHhArLOIB5CJBYO/+y
wpaZC9hdFN9xT0pQhmKAutIc9Vht6daxltv6SD6h3s1j/h9L/HZJGMipbnQ9X0cib1Cv9YL6GJSx
1k38KIqxlrNgDCPr+IAtoTx7KJADgPIpWxNqQQC3477i1WG9TSN5ClY4zzBRWa7S0xdhi9iQ+QyI
f6/S+w+1Le09JmpcCRfG7fI4Gn9TA3NsT20XWFX5IT6EkGvzVqt7mwg4Azrt6ixpCiLOz61/lYSW
DobR5uVJ9UkV5zLxMSNldVBRqupfguWHL3m7uQb6F4Z77Cxf0NOcffBv+fCN+yJy1eHgwV+hdIqP
CXiJPL2gAKxMJgiCn/KQRco2w2iRkoQWmWalmvPBV4kUcQQDPI8GOQ7GCPrEiqMgZhqJhG3TVmAR
BsAp9DVLg9/AfrX/3w96bj16zvSgidLWYfoEqSog143B8VQEgCUZp+ji3AcXee39MkH41b+Fhz9V
ZiDEhOg=
`pragma protect end_protected
