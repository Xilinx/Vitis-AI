`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0lo0VOrZ7GskXR0XP0vxuG1qSsEV+gLM6DXZ4Yhu0f5PujHxoScHXAGO
SOAmWF430QVnF+y3O5M+swMRLq3wJpBqLc3/XRbY/FUQgjExH7n9FaEOLIW4obH/07d0MIL1EY2d
NnqJnisIk3Os3o/bGq6l5RhjZfRs47itM6Kl+1rQ3sA1VK1vW2s03vu+wf8sk+yfevydkQCerVkx
OxvN/XhUBtqBvYnQo+rsu60VeTuhHKo3MAs1vH/prXXDGxC1yxlGVenO5R92GoG9WQNmCCek4L8E
JI3mCqPVo44tePrwLRvycmzolCqc7ylAeoBq/mabjdwuY+qdS5KRDAeBVHoW5INFu8mvCqQYKlIW
KvuChHiX0qRTuoc0LNCVG/AuewNiRVD83tRENCYKvCqmH3HVJ0xTIheNQ/Txhog8gHZv8nl6NdHw
yuZBfEYL+sZiO8z9bFG0L/2PKI96BAWc81ZrQ7iVHZXgkxpfiQd4cYWxmB9Y6JTcQhwsw27lHDbL
xnGed9JXD+lfyjM7mJospwJ9D4cDWAIa/e9hl1H7f4KyWmNxwM6L4tq6SHIrnGEqJzh7wyKQDvWH
D/jDY5hrxFSFzM3YMqgX0cRfFkvekTCx5nVK3k4Vx5aBABp5Z/pwjwvWBFOzP+pjxHybpfAjnWSa
+IbQlMpG+iZBxRNyiqqcuO5dHCvIFr+dP8ywXw5Lozro9jxbwRsZYbh0WR1OvNTaGk0DlrwgSUuC
jgaO+xI5ec67jBkS2Xv/s0wWoVRRrsHYDNexyXVBPc07Gvu6yGoPHsem+xqTRFzSlHMnWEb3Pttu
Y77AQTSlg7xPurfxIhL0yPuAKpun06BWCmy6FH7UxUZnUO3YHj0jcowf257YIQvLBFw89L7/rgpN
T7QnetldJy7RLY/iOVdz9/1stCfQsvH6f8IEHBfk0F1jEn7dzdjZtwSiaxse7wqJUu4MRtyMQXoD
K3fbjG723/J0J51wrbhLhSUVv9x6mNTd070nOz95cnsYlYPGiH9AJC3qqcSqLXey4mgHcj5qX/TF
D3cva8xj+dmA0O+ib/ytdD6RZv+TvE1byncn5q8urr26BDjihOT/yyHexvzX5UzYnIc3w4Zdaff6
ZE3QeUlrpT7WMND3M8sNozqc1YrrY7V7r8m/WvdMtcfXcW2GjOxikIX3gJJAFWG5nWaiyMVQ0uYX
noNzoTWkvC6NwuSSK7CxLgVUYEX+AYRw/4a6Sgxfx8PtV/gA6csnLecmzmoxs3vw/O8zyd9ywtMg
VtsCBjPmTy/9N5RMJX/nVoabL0ciXv7WBhR7NAJubvCB9CbmddyNL7idBHKLQSF1zmYhQNW93CFE
cqBazkUgTDw4X8hVPRasrga2Gmo6nOgSoiqTyjA23JfozQGbixdz2MfMvOhfF755detbB5tBRjXZ
fr/OnH7XhohKjLMG5eHXI3/wxPmmyI0tTgr1ujm7R7At74V7YNFtCEK4tdUDa16EgS0jgBY0KCe/
ZlM6dPYBuUgEfdxUN5GrHDFF1bKB9/ktlhjYKVOEcElUVuzOXHuM1PC8iOLZ7LrDqrVeSDtKRayN
e8RtEpWV189Kr+afgYwfomeQhJ/bNA0U5rOaeaTUhHxoZGc/2dQE4HBe5/UdokEnoNeqR9rBFUA1
n/ta0H0rwi0UJ04AhNhiegaYVVHWtkX1sCgWzXC209EpYuJ+CqpTj26SGxbO8ymaKEeuv4QdSdUv
yaAZK+Euvmn+Njn/GgSF1N+vclrcrqvIFUFPRbY70bLwvt91fkc2UMgoQ8zvPZBK44ds99c1f4Ma
ElRyPaZOWz88jGBR45RIWcwXFZlSdBRS35h41nN+zlWTiYtB6p2YHHjlEWOB9eWqtTpGc6JC6fEp
9xDRMkzAvvF76TryD5ZMDk+p7Va0qOTboDHqnVup61p3JhaX2JSaKS5beu5heLAFGzt7yhHhEwHp
XeJeT4ClCXfiuwbHj6RdhqmoSP8P/xeVXfDkxskIrcmlL7s24uf+BkDS8kXlQW5F/OXNsxljSwYF
seITALWFRDjM0sHH1MwrepT7fwkJ5r+YigcBXN8Byed7393Zi7pULtROElb61MGrSQX7PrQIjk7c
zgATwccHF8zbrQnmxBo78GhlCpVQHCVnjkLa6gDNz+At4gZmbTea9O3GiwC6J6AFjm2WskcfH8+F
3TDZThJ9+9BGieWKBcBsUX6Fl2RTwVeSluNA8bx4aJbCSTeiue7ZlDBGfdDrM2Bxa34vVoDsyqah
OmfEjCOBcAFZfqSbno/xPZWwma87n6lMmhlHuCCz5g612Bkz1Pjk5aXyOREFO8ufDK+neIRybtDw
4qC111bCG7O9iZS5qreP4IGu+9PTtvyJqleMBTV7ZiznkJeoTA8V13z6eKLkniij0RltVYHX4QJw
J73U1hNppKwC+ScLPUHw3zMGeYlDsK8F+IJxJ5cxIenjJhrNBP6tkROu790FwYnYQjFj4Tgv+JpV
tVO6h4gGdkp55g3sAi6zNTvmXazMmovzcxUGvBTb9nZJIMV44ZMybMhCXaTP7zPY87GEDY80kCYq
TnT0lVe/w8/3czzFjSfuuFg6YZXlik3sPZY9AAH4QptBpxcbSbz/1k6mnWgstrWsZ01XDjGEqaVi
S7sxop3bwO0oHogkl1pMCBLgBV4z5Etk//ZiXjbA3yf9E0rAyxfpcNR3rOA8u1l2nOSE3F1qlRMj
5sHyd7HEfYDv2LK2nOL3M5JexEVg+sKx8haKq+DfsktfCxM/v/y81Pu7IBzPqckEUbckhQfjlgaC
ScOb2VoLECByzyS0uHl1ALJGQdoUgiA9PoKceXVLJorZdK8OpthhFZhGkh0nDnyQ8JJtsjIurbWF
wtFeWunmx+7kfHgiF9O2D+MsHLAtp3poMj7i+qwEY26Gq6dlhQdvO42K9EejN6BX/ZwPggQIkpQY
OB5n1ObHQuBmUNlbbXBRqNyp1wsZzJ9mnnIXFwKcp7xg34wefpL7/MIatndvKHE2P6vXdw63oHoo
/sgTjgzkJlyzMrvnnpJ+0mSPR2hvE80E0qenBI1DsiAGqLAqtoSemg4RjGfDMzCLNnPJ4RKnkxRv
kCoWhWHg8TwS3bG2g/GIALfS0/vgiDBDdU+GrrAGJsI1lIIEU9J5tjp+NbE1JVCq/wjUI24LlRCT
Nog7IQuY7+lSxTds9sniiGeOB+hWabCinNaoyqeKaEmAU6RHMaJ3bP0PEI9NhBdwDU7jDTVJPd/V
QOaB1enZm6Q36bW/DwDtGVyeSZ+MmaUMEu3N7tkL29mbVtKroSLoPtR/lb4C8O1os8PSYPg4HOtN
lncFjbVmATvXrQMl2BgDPPsbYUT7K58lgImBuxJntBMPCdMKZvErQEEkKTsbEzlJXCfsQ+lDuXad
OqCQB9gWbjflHM/Qwfyc3xaAUsB7ITNiC1Rt3dpZ7/iuziNSYaCulUUtBGsu/6Q7KyCquSoZbl1l
4GBWycivQf/dqhgTPoi8x+6167bnuzvFMt4DAzqOlh6UKxtvr8gg43doas4huwcJEAskGpxavRWt
FM9G9G1GLJL94b6BQCXZIOWUetpUQaph3In/sUpaPqw0sO5LCE6AdsR8xJeHsBimNOlXvyIrESos
ar/VyMdIzYO4v+/iHj41XxR8H7JY3MBTIN/ynPTm0oEWiaJu3n59X5mQeREef2RzUG7oNUFgkfLX
kZbLEjpK8QC+ySlWCcJCHIC/WSI4xwEnRWtTqppBljE1tCywlqxgep87ZsCAhB+Og/0rMUh2oGka
PMjAbi7uEDcygEj8Dp47lrPkVYZqMZ6Ku6s660PT+z9U2YvaCSbK1dMXRLXAbwkFaBWElYpiW1zp
SBYqCFzHOXB/shsr8+w+hZEXTaEP7kxrCY013Nd1bjGbg/qqMKcjCIDnHWcNXvgCHc3uFVfhe0IA
A/aB4LonyVVLYm+48IvP5LOSxBCfl7OP5Klv+gMaE1B0vP43f1rbqrzPhXt66+IM2a72PbrEisKC
FTGE8nftYz6Hi0DE1N6/FgROvJiJTP8SlMHRGfcisYOHaXWCQG0fCy5niUt1zZBZs+bYV0f1cSNE
01xkstzxus3wqzgMec0M8TqKBFrd6AyPNvvOaPaBmhmrjdN/59x13YD/uKt3M3pYBHo6Y+kKmZ4C
4ugdg7WnHjoC0Q8C/epw9pamE4MRhYmxErGcm/ZgpGe487OXw5qpDKxvNrYUn2pPAfs4So44w0mX
Zhji/dz17bMYE+6wyQ03o/1dZz1bmlCG9xIkUot268npq8UHL3CvTJaP9XW20gEsP0Sfbp/jU4Pv
qTp7GiL/tNk/I4PV1UVYoEhqoq3txNWXVokKwrsa0deFpYGKAgra7Rb9F0LnWkRt+FRlbFfssv6v
z8uf5o85X60+Ii0qFYZVOYnAXbTr1ZEXMy+rwaPgoBWjxDaTjSYVIHVQ0zSAqDZN3O4w91bGOT1E
JZnSgnhUSrGVa0vVb+TW0qnAE3wrUXMnNu4DCPhYFep4sLD0AaMo1HDMNGX9X/xPkVK/S64nxPxt
Vi3pXS/2AWaHLseqVu7IGyUJeF0UmM9WzSnnN0KGEJNZDC8BtfKH9lUacx7Lfr7voY4dyhEcyc51
4miSBwinB5AbA3pBEy4xqdAeyQ0GlQ/JIdbvCzpV8DKq7/q4Kv9AS3W1x0DKSvveWyfyjeUt8nKm
af7BYIzVa3U4JsBU82eb+RqMA3JkdlqP5jeYMxo9UudfWSuBL2qjYEOCCUxHECcTpXtGrHw+Dk7l
+oWF5sJaivPhEs7l0wpEQwq3OAsUsnllcBhPdMbh06nJTuxFrYbUj6q+ENSK1vsZ/IlzMHCSZj5A
Mv+fraXjuDRm92iQVY3P7SHrGF9+OeSdxyKWTN3tMfVm7TeEGKup0PHl8sC7BcvXv6AJJFcYNaQh
Cj0RGoa7DDHifRIaLG9ucGFX3FlfYycZUrz462+4EZccEihgwEjBg6WKY/SYw/q2SWyaaFD1ZXue
4FjFKNnk46QKStUvidmQmlPtxrjTzeO9vKyH0FrCI53+SYFQNFg1IYlc9TE/sfve3KTml/UNduv3
CJNs17N6rfodOnrHvtvKNU0wmvlPP0OF+PePWagsTAf46u9TMxwqP1A8FtBl/a05ycKMhnvlHVh0
8Td25Csha1UkvoVMC5v6aBmip9H+wumNyG9ztV+dhq6jDAX16R4lmb5y8u9Qvu9deY29SPSd6oQU
VN2y7+ERNBLBA6wzezNe7E3SK7ejnCdoFs0e7y4fDYbsTYIvOFYWFEpuFGxhZ036SaPcFdIZKHHB
SSECPuWB6JMKuVpDFKl4uYDWePoTs0IkTET8BfNdoOcb3zrtkzmsAegDY5GloJ13BWrWex9kzdYh
qWw38BO4iic2buhrPKrl+x7HvQa1wvnHIxKMpZZRvlY4I8kyAO4p4coTbhL4YsDpxj8GV8BIICzM
u46G4oySwgwapSmMmrBaPB6mjvre9MzTZDA65DrodUlDI+xxhIbT2JV6YaQOXF3VPFgKtft5Wbze
5PxyqZzGwL+05Yy9Tmi72EnAwc8q4TNRr+rvkGipd63zEgR1bwHAZ14dOr7e4NhnMVcKKf58whei
1W5HurMqYAF2JN+j4EozvA177qsSYhqILAHPmzrWUsKPA033OWc=
`pragma protect end_protected
