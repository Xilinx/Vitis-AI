/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPSzFjNfvAZem/ebSF657q23aiHdwClHoGTEXbZvHS5Ovens/lzi32PkN3
Bt9P3sjBzCaCyeZEh7+K28i3ko9Z8HM5LF9Agv0NaLeR9LS/E58PP6bmuqtJKQ/Sxexs1D4BOp2q
tBJXrH2V7T53HcsvY0c74JpKgnQyG6gYkg8SHmWm9sDq4Ir9iH96BHh3vtez8ZP9Ev8Z1JRRMpmL
XYCMGijemxJdHY59xU/EKiLt5NrxjguListGPa1DFadv3Z0mjn3zawL9xk0YKyF+WbBlowmR+9YW
Z6rMj4eNAlg9EHwVGBtqt955Dk7/tZVGifFKwr6rAoeQNdIoOjp4EzA9NmQ5qbiLRVWnHhPd8Rsj
PD/EZJjVoXFU1AsLrsaACJO1X74cZ+bX6ZdhlDChLXzDVbYj6gN137Hh+aZsSb3vUDT2CMf8ZVxC
EIhQqyw9mc6RDbYdsVmbrxI5aqN+UYbk4EfEkDnYm5IlaXrw/nbESGsDz3PRvmgDHE5DsyJv4WoW
YzeWd5/sSMp65/E4OM8z6sTNlWSHLtdnwXIRV+YvoYU4vzkg1iZIgjPqUKYMg3Ze1GZoQ1cMLuPz
pnp4g4c8DEME1dL8E6cjwKLpjEeIVQuh/AhC8+m0hdSkXz0NMFrqFV7GRrgrbbFONnYxoDjaAkdg
drjaYTZFQkCZSrVaFSPxpqRl9fXsSEjxoC63TTJkrjJojwfo5ObjaXAlTNxpOL24qjj7TQGnhYf4
+eCH6/PlegETFeZhOxL45KWe4OZ8ynP0u0Lckv9leHoHEAIkgyr6s8kzxJF2YccFudH+F4LUYj3J
DMAROGVG1WzCAVdtiKD/GQQ88LmMQ2KCEsBqhYzb2RpBsOobvyH70e3HWWkQ0txt1rWHrlb/c3Zz
8Vgm3QGzXCcktroNNaXWPnFehdmRAdmyxamaQEAFysYWNWurRdEL49ZPS4DjI2M/Pd4p0W9MnFnN
iaGYKVvHvcgPkQjVOY3U2Pkbuiw4ljOKx0XELbYrY/jY8q9ktu1T2wLGOEDEmJSy7yJ65hPZpBt0
CiQa0qEx1XtPO3dF2qQ1yvW4yV1mxsBjr5QXjXqSdWANyOtNUctYLei9UMn7vss3cXuBvdAXxype
NHspM8y1HMPp8HTyQUmwVI3cb/H07RoCnlWPjEuoKdDdW72dt7+oqYW2dI3fRsCU6pjnb5jAd2TU
E5ZoEyC3vWfH2klH2DCKThTpJ//pDF+91rvK5PHyQJCYQ6sQ9rFBYLknMWy+scUZb4icvFpqvRjj
7XFPL0KvOn7EPoOFx8PEuDP29eonkUbSn9K5ljaUQpAvtExw+kihXV4CdxgpLtNPSLuo3Xry26Bf
Z9GDH5I/GxJeFntPu53iWxLEDJxtTQ59k5ELfr441jS/6xRLWnNOCxxeqW0Pj1c2M3KlwvzBcHs8
hp42Va1xif3I+NeU+EdrB+EoWgTO5C0wY557LtnXr/nSlrqRkKOMhEoKyh8Tph6lyufkyY+v3BYf
/voRcq34H8LgevDDYH52XHIHPf81MfyVc4KI0R6R98jReKJOjwK6VhBwMIfLzZ48LkSSAWPbbcGm
sgzquiybOHjW4v3tCM8hl3GuvAjLI7SypiNQgPUmu9E+dPGJX4YM5O+Lya844pboR5W3Gc+1wwPW
Q74JL8eI6MHfe6K8hgUucMdc2O1Y9Stu5cbNKfTMBPa9FEomByj1CFUMOr1a0WXLHiWj/y3IONKU
Tax7jKOJZzat6w+E75bcK6c5SpuwRVxxPxIGOFYFfQT5ujFXiEeg4/IgylEvXq7RAVKerIfGQD7c
In08q3hr9QYTCvhDK8LeIGNhusi7DVQHP8kexRhSbm7SOkUktYW+gS6vDkrYI5Dfqs2YaDn87VfJ
9bd87a8q+fCBcIETcUn4VFziYT3R6qqPYJQ5XzPSaUi3+cjkFyQksfdYoWJEwxuEJXiBzqHomQf1
29q32wgItS1koE0REn/MYgmLzE+ZR/tVxniARbchQkTBGm8kKRxq7bmEE0FZ4renwUiNr4MYMH4o
hoZrPqRpUe5n1VN5WxaSK0tfXMHTw7hRIVYlIw98FqoX8M0BvmyeKdvy0AOubh5vBa6Ob0U/lxJ/
wYzm1JWpNNumNY/5dcPn6t9G8dxDDj4qctU/U8RZsw6m6aHyiT7xk9cueqilreN0GyeivDMD7ynk
u10UDWID/pDDYY62WNIXULJCDm9/nuzPnUGZgoZkCfjScXI4Ej4X/Z/HvwxMoFWJETnR3y1KwT68
VY2eN5VECjgxvStr0jExVD9m0XDjGVR37JThtmZOpkK8VP2Hhz01VSJrXs4FYjbnE6r1Y0yGYZ7s
rg4D1+UUeV6rlDk5KuZg/XK6Z+9USYqQnnUKS9W5neB2xkxTIvlPsc+MdplsmR7v+yIdBGavAAL/
NRUkIj/DxC3SWFTvaGZfA/HxD+lsFG80rZSq4ytNv8lz7oJB5ZHQUeTOnmuWhKihKMpOyJ+tXUFh
ARJc2KnkMpdR93vi9VWA/uVhfY5D3KzM0t4pfxQ3rk1yB4T4O1CYmYMf7wJsk4s6MQ59x+MffDCB
1q2tNfkkV5343hQevb44rQeycljh78AuFWOHFQIqNYZG2+NEnugqR2VKCqPYRrZapNI8FRHHnvJC
kSqnzr0GU2vBnnCTeO4OKir+87ugOWQHNUYsR9ToIEbbVNU0phsspaowhjMkabGXtqecsrUurauf
1gMEJ8EwcAmEDgTPnx5Kg12cCAvJUXRgvzMvwbRRX5ZA83t27nhe5hKFDxWAGtqwFo8o8qzOIgh3
T4PNIO+wV3bo69bPoBtcT1tghjhqC6tHnLJ6oMhEw+heY4kHq7plIDwqGCUjIEen+92W6cmvLlmE
wwL+Fyp3Es5UCDnzlZpFtCD3XcCSiJd1gw5xurkiAaeh82GnKjSbOp2yPDa8mZ9afzBfJ8es8ALK
QIJphLkafz07TYfb8M5aw1lTnGGxUkF40AsZwlN3ojTo4lBJ61Ti2maG/7au++ApzSAthxdOuuKB
TQGcIVzGLW7j5fPPbhUK0/RLCi2ue38joy3OSvGFpoN8+huZXVlJNGVqe4pJV3HODUeGcO3bn9Zd
2Sz5zsdgf9PBnKfXH2+ljYS/jHr0VvEgH+mb4MbQj5vcUrs+YvXZXG/3vkoBi/TshuX+fCwuZHt+
fvar5ZX6GGXCVAbhPVt89Pe5NrRNhMLufIuit3DQedgRxR1AWd5bvKFf/PYAS5ksw2UJsKuxGtSL
xMIV1OXOrKZqdaBFjliv1Hq4QcI7zDeJHwuzYP36iUI/41Z7/jyf9ZGMW5wqDZ1i5wOa4jmaPhFd
ZdUzHZRPkLlFxBNbo1CK5p+fa7pYkJfbGIFk7uFmP7aoJTAeeOZQ7dEoohXslOVSS84nttrCKZgM
4cl8LH+kd3fW5LyORZtJx2hZFNr4kdpF7Lt7X2Yg9VjSPB8dQLa3jd8Dy5oiruOxsRR6C9GDzJTu
1co5f1qgcn4AqWwzL7nXgHF4UG6nH1exqKk9nu1RM1NA4nfHMLX3aphrBaqSnTGWO7ldR9lKvnFg
uyYWKmnuMnjMtLdepJukb7dClwRpPLuO/+kqhFf5X5QopMYmo0LRKV1vJxoKVrtypTc4GR7SAesA
yqAi5kIuCtmV3weDKiKoSACzdqqoc4usz4Jmk0RE/wVcE50/kjsLlyLEgoGZejZsU4OosBHUSYp1
lRUvwpaGU6i6acgGvvI0O1zdxjcHfL40HYfzjMq+Pm7m6RjY8/zWvhkrQLwkvKSQS6GYPofGmS8/
Cj6bErndmAUb1n9KG7EzrGg2gCtPBa2ihBiAm3jvU2oDTk+hUByaHVNHK/5S9iP0ZHYxVHUJvwhY
vA5dt47teksjzktWN+1UFSvJgBgC/7VyJDdjjcJvg92XDGyveN81JKaylTVEqW5hmYwkOCCEQirO
bC3lBOHGoaXmnM4OzSvYcKcDmN1lAXrd5E1orXqwQ09uh506iPr080Oo9+AQWEBn1gCkkMDBZ8lj
6Ze8TaIiaChEyBUH4UxPV4NMnDyS8DabXRtQYR68UePVDqW5xzMvV+8+n12eZ845qkEcuplbjU5d
C1D4p5sooh0vyXHRTUT5UKLPo/CyN3M4Wy8RntN4bPHpV1pRRmCwhgi+BIxVHTA6WTJGgcuH1eVG
PfsLeXjxBqttH7ZONnawTflDPg77gKCrBK1BiDvNSymX6WCFPrFNA5t0Hrcj+3vAYSTgchePlIRs
85VrWQdVLQ7beMnoWERO+pQerYY+HjyRt2O5jthIxJelq130hMABNUiMM4uS8fhhDgIBOgbOZgGi
XTmDY9iP7nsEZ3chF6Dg2crvR8URuCW3v0635HglMBU19NJ+vrjoT31NbOo+4a1Z3TITKkbEvpo7
2lulvricAPDdz+ESMCI6x3jLyUWrpf0CpL+iDYim1O09qGuqR57AnJJzfIYvq6JhvXyT+SVNCcKN
QZWQweAe+dXFJGZPLwvDFj2Gtvv4S3WKSL62Omf2DhaHL4aaqKmOYiMi1EVwLE6/m2DT2l9yjuLa
bHm111fORS10IKHNKk2FiYlotYchKLnTWBAMXlHDK7BA4Z4ucFxL4d8S1CbfEDN7pU65Wivz9+32
8Z9doVocul4eRd89VJCvsHLp4ki3dTMkgqU+pGogR24wdgXae5FwGOkXfQp9p07Viir4T1I0afx3
A2HANUL9wflruR+HnRbxhhKEU0jU1zu7pW4POCIr77Ui/cJQJMTohAKEJ18E7jySbWMcp3cwoY/n
xP4b3vU3Z4DXUAztT6Ro4R/WrWOb6CF4FG14p7+nOfnxk6CnRw21o7drPbaFWP/33upww5XorQnS
Ghti5E/uQarYDNjepgCwBMc8QrI9n0NjrdkG3nWOGxoWRMRchJuW9oyV6+HHsji/u0NbV6gD9v2c
Mk3r9e8x5U94sjW4kVw3ShvK1bVpOjWtflPF17wWephw3Kj3jyrJ+HYuiE9N/iD2nQ9venjmhTJw
yhHq1nXmeMIUHgxsVuCchhZR9H/o/qS9I5YLzB3mWwQuKSKUQzLYEcsNRRZhlIkvEiKWkzzcSBKI
gP03Mx4RRAiNydv/gqjobpno/QgOjE2UctTQu/3xUWUp9SFzuzNE7OX33Apkz8wb0X9LEta/n6LZ
B89POuPic9zGyti8Ywq9crmIT7w1Y1SvKxKLKkvcAp3x21CsSm++so+WiEiyOUnYccuHAwIzMXJa
uaoVcSQ1QZxmdX5GITWhNA6FniRCscJPNq5vJxE6QetpgYsYDp+Ucfgx7/r0vyGiQoopmD8AaycQ
B9K8XqFKAzxeR2SsoCWi8xSJWagTzYE1qp8OBTqJJqaZGzF1ekanzcMn+O/XuwMFs9uVCZ/cyZyq
hLHRWNa1reg9pv1yFvCajGXwnFkHQg8QIJCx20VBpdn2nts4GZN7eBcW8Xt007kMGOF5SZyrmM31
z6xZ2CJ8heDJZzs/VvH4mK31Kcd99hUIUNtRaV1IZsUzEsaBekAf05rkqQILpPfbB/WaFIcfnLS6
MrFL+EwppmX5dovi2vvwcQVXng4GaKx98sM6H8g6+Pr+W58m6OncDIpdd21no/asHPpkHw3zourJ
g5Vn5orkY8LVBKFAfo1m27/D5bh078VtZmIfR4IODWQEDLpj1Hqx7ND9r9yMW44XvQ1Hth0eTRnC
/YkpFKs9PfSD61qDiPTiFfGkueH/ASWaOE9BVSAyR7tiagxVaOwS19HLW+RDy5Kp/T37PmREixwx
mYE1bA0umhuDVsbUenZ4ePf2U0B7Zy9edf2ipgEeTaaEMr9D8qVfWmEmK3Sp5TDWars7XW47WicI
IKhulLK49RoZkhd3BFesTpeUYYbDK9a5+p7gRQC8T9E5B5bOEeBY0t0Faz+NF67syWuUBJzuZs2L
1i5D9l8O5VnZJeuI7aWapAWJSadIydCv/a0biCW6KnOGCF1vkzCjRybhzarofm/P2QRMIhC1SZLM
8crV36BMsDOkSd56kh8LFIZj6/313vUnzy8MCGfWjr/J0cPa82yt1xbOE8/v+qcl/6RTXyW98ihw
XceoRSp5Lx+FviQnYbQLUWyFM2+VmyYdllK0QIBvmX/BUDP/lUK8n00/nDZ4P71ec3eQhkvYRhs6
pMbLyrukxEOB//GC5fEL3opzBFhPRjW6DwSr8QijT4XIdxTOCctuMJnxggePDcKOnRc+TVN17IQf
OjQ2YOVOzfX/zBHIoqVrPCneEEWmlSSZChgu7YMhemOMgPbHL7HElw/9aLpR8p2XSuJY2XmS7reJ
fsXwAxu65XZkQRgYLi0Gi/G1asyCdQiecZVOGmsFlZ6Z4dvivSSkv2slYtXXuXOkYCRDGLBjHmcH
vg0Imy7jy25rQVSzplQbybPu/O7NBAPYoqsJg6/bc+eqzJNy5QI5bw5q5s90B7Cgd1c7fF9fRg4z
kVcuxDklyZweHMc3usBLuUOO4CUzNbKLzVnSFWjDcA+RFQDqacGsGCGElQushOGY2aqAWGbE+tWO
hIkJW8BelfE84Dl6K+1wN8PB0Lx9QCEarxKhzgF5/iF5zdWnH43cqh4/U0c6+p3KdGmtyz6tTRFO
unVuhR9ybcZliIMBIIkgNpCgzhsr16JkArHuqgOq4iA5ZnJs2uk4JTCQajkp6EI/ubuOepNOYTGj
VDA13WYtFcV5+GI+lykr2LxXDx6ZROVVU0L0D5IZNgFs+sQYFPTfyPqT9hVXfVI2gHZz/L63pW9i
aIrJfbl4lRgXj5c/9T/Wu0QeJNaeD6/I7T5yX+3gxhM71W2G/5JEMzQpd//ZysUQ5oQ9q1mHZEgy
jta9JPzjSfJM1yKTWEQpmHL3/9BfebXKFjk6jFEjPRkm5xj8LKRVWtkpXRhreftOK5A49pgjsf8Z
b1WKV6Q1W6YrjMzTS8CjmUT8S3KKK5Uy1jqQuJ/moLZ3BYfP2L2hiHTIZ7MGZX5I/5OoxR+WHE7m
PvfcYp/VcdNDiMPtDZIA/H3BZu0kIkH2PpSrEG+TN3h/O3ikRy+VvHzBItUCX2TE2Yh2k7aKFCR7
+JMUs4Pd7VQSh5bbc4LxnvmOw1J0rhGPZGJgr2Be0AnTvTmI+2tCGJd4c7n0kKfjV6anM2ehJht7
Du4Z1nxqvGy3h6ibdrKrgbjqsIbuFgxw9E0jf3QD3WzvhzSyhITVapIUvjFCqemMfT8QX2jU8pOd
6CjVIVMgu2Ypb+UO4ErmMkGekIvqHE+5xXtSnBvo/sK+LxjK/O9R3Jxw7rKRPo14kdrm1tFjd1WK
F+ltBQvAYnQCpwaM4+mJFw0Y2tkQ+4tgADcbcoSP3ns45d9kpLbNEsjaTbpqtxjAGUcPhExR27Bk
GkO3RgBdwe6iM1NzwaO8U4aq6KgFPrScynkn5eR+aYm9ggwKpFa1IEnhM6XqVwGIDTl0VGuaQGrl
01ivFQgR2E/7Bj5nkLutVZ7Y8dclI+ST06Zr9lZ+z3ZGD4xMpmEBl/l11NdT626dCgJR0BtCMAfK
TXKRfJoAoCL7Q4aTNzeLoTS3xAPwcDPbuZNEdElpGvIHbRi6rGkxqcxxRc78FS+EH282k9s40jTi
Fi1LoSAbLXFcSmtLKIZISxFKUrMNZRXxCzJwQukfCYllk5OG2lb1GqRE6LULWtMyEZb0TK8rz20p
TtV8DK2J70a1UQ6elvBN2JORWkOjuOY0xPWJv19dfCi4yykiFxOiqhms8lMLXU9b2qaUVUQuHrsP
eauY8Asl4bxiIFubqkqbs0YA+z8LqNz5J2YgN83pEWGNs6wk2C7bcpYQEBQMRZpynGCpZ8zc8u+H
qn7jIbKZLqGXXNYuGm68sSMxN9oQnczdAF8j6AJqQAFznMV8MJLekFvR39CgY2rnCpuVN+vGRtuO
OZHVlIaJpmzZhwQTFPr8H5UancGqiLG3+BnvZaFMCGSXWFKA8tclz6Hfqwfx4p+9Gy+y7ewqX6xu
cB1jUWePh8+Q5bq7j9cGPcBlAFGUZE6HMgBLvt7rIrHVPp9VaTPLqCCw0GHGIwlGD4ccln0jgbVB
kF9Rk7x1fbxpJBLCi7VwNJDc0GUk+gJAhQbNMlf7I2yBFSd/otyVyzVy7pJoTBMeVoHqkOXzQVrz
sue98vH5HMHqMUhpJLytHsW3DJc2PPakHg+UZaaAlDsLE3Cm52KJGtD7NRYeS1egg3s/++kgjP0T
xG1SRd4QTQH4z9X07vo9HnmOG7lGGfT2c65BtfQ/EvPEJozROPKfymxDqAIehaKWlXQXW3Yfb6Fh
45AgYGfDdlR5BYxzRErV2qBhonDooydREih0CKvDBDaco4VF+a+EhocJUzVfMyTnuxI7bULkV3nH
sC5IR6p1WHpEAdw9vvBsgxFjgSfn5S2NlKC+So/KcJyb5P+lp6/9nwmXWW8xio0dqKioH1rr7A9o
0gr69OVIzexdE5rV72whEk/8JQTUB4HIq/70onzTkS2wJKfJsSQnDitv3f7d6EFNy8448xvt1CFV
oQELCUVJbo3vexizNu6/EnFsEqEq1sx/RTz+QJl12WLE6eE+gnl8sNfjT+LLWlLsr4QkSuJ8WbT2
CWIKWbFKTI/BKUwJ3U2RFkRZT5C2ECVdFp2ngMRhVLc1584X3p1Mt5UBW1xnORLmpewlR1xK4F1A
oPt8YxZ3KCS4CthPt2TbgfW4y90YwoJCyouHjLKIU1O3SFKPukVEo+g9PZlaOwV6TpqJIJY9mQgT
PjG+N8oitIrOTMtOPFL2S7Zu3DqWwaVhdaRGLisd4YYMUhZKgLGeOlCDr/W8+rhQVbT1r669wo3A
ym3GFtig59kNtwEYuQQaVrxveX6pM2CWcvo2u1OqhbKH/UL3rxKPdkxDkb/HNkv09z5GrHa8OT2c
+wVOPSBlzSkAnth1Zdpf1VG8YvS5sD49sdw+oijppYrNwse7YHM9dyjTRDhZW8QvKV8WO9viquKP
0lZkzlK12znlR07KP4RG7QeqF213DS9fWpUC9I1EOgFbHXcWE3oJDn14nYSgpspsJ2P87N9dE7Ku
HfFl4TAQiux+4iG/ncPv54wcBck29CbHTdlMiBmWxl5wn5C7OdS1lIej/X+48t9pcyP34WIx1ouz
UiaXOhBkEk88FBZXhi32rWLEmqh3wjuL+iMdj7hAdKcFKtdfsdyuyd1ofnzqpN4YmwrlxlN+9tve
BWkNZZbABzC8uV0hsgEAj1/5V+Y/tyEgY0hv9uaPj4oNh0LuVyYK1jD5xgIyogV5Ii2UkRcIwhuf
6AH/vEnCCTJKWPPDc3yMW2Tho9ly8YQBKRxMRBpML/so0UENZ8itJGKBcIIGDCoixL8rR1x+tgI8
w8hriuTb3I1chu1ak603mkrpC0E+nKW+rOxX3U4NhE6DAVqW70E7jGMGfzNUS3OdWeARIDngJ/AW
+JdxjBuejib0bMF1Fd4PlZS/9Imrtut2w5xsb8K0X+SpTIXcx3bLyEx/xgCx9b6SOazLo4EfuU9/
3BpJgK1FhR/SCjDPtTVGIbpfj3v7kF4LFP7wDyCCfRM/7Qyv8N8LQzWRh9XJDKihZCkLensFZ+Y2
0+D65jzH0tdHqZM+qv7zoP4JT/SPwe2yXRNp3Pc06pc81G7galyx/GUl/wBpSID3JmVvK1yO5C6j
UhvBHvS0mRASOR84f6PxTORQDdJFQt8GwjZd+qLEGr7urSobE1UWbvyJAErpBg0SoW25CiWH2G1W
i7NScPrqmCuKEec4gQ7dGcwAJauyzs+hY+pe52O9WkBMUUAafJ2qjWIEd4xWMOdFBHplyJ6SwFzK
RCLlof2ANw71GZ54l89Q2oZg2qpxcV3Lm0nbb6LvPBtxm6i1XpbR60V+bq+Fn5I5rNYaYPpGz5DP
Inhj804LlMXpeYgWyXh5G1+9BIi5vcVZQltkw1hlRITOPG4qZ9zSDFTMhyBymce1QhGV5FhWB0i0
mflGYBY4I7I4afcqAFCzx43jaBEnAFXS3AJHCM3HXzOCCdbpEftuqjuxk4Kp6tBUV9sfwcAftag8
n+3gwdXEkv50Puauxn8VVpcG/2XF1yE6LZlm84Ga4WiGyGlXSvUkJOe4+zcR60NiK7/8n8st9Snu
dzME+CyN8R/+C8dOn6p7r8INmI6o6asvXqD/oTDSZruNd9bt10L3lbPemtbwUvC0ocqZoJ35aF1V
ylKRP/yQ1GHILZ2zdQCaLolF4mx9H4IRaNGA5mLYHMQfzhe22KXcHgwNh893Sa1jmZFWhBeBErmX
SRZPHdOQ8qObE+/4ZF+S4ixyef6k2+AuIxPonnlHYUTf6WLnPMLSfo6LkKqCavN/+npKI8jNSlYS
ASkaPtJy2Io6vi59/XP4QWdItOJTjDHhaEXwCB+folC02f9AxBC+gWZv00XEM2lc1h8DklApeK8Q
KdqqkZTPUF7Jj/RPBeRqgr2+lYmbarjeqzATSLpxc+FX6assTWQitBM4rocjgZxm6LwpIh3vAB7D
BaHJnqTDxCVE31/3LOHmpVntMgd7dykeP1hvUFU3BG7wQnq56vDTQGcaaB8PsgxF/1ZWiL4fATce
gY/BDdcdYTyPPmsMfbW+xtVxNjQSxd3pQhHE4XKw0YKAwVbcweZimn3KOH5OZZmzhO+wGLZLBGHe
jD7YEPYU2UbLOTVB0w+jVpQ4tx4HecsL4jIqz/oUF+B1nHDqm0Mac/5vEMWCAMRKWG5oadfsLhIt
9MvlEAKtstPfVRvK0Xl9tE4yqSbOFYClVc70gclFt0yqhSovVdAD8e5fBTUIaUB0mtL5XIavF2K7
rr0toTRpyFRy2lgylKzClkZ+bEK+bFkBeFF2A0pYxpdepR3ASZ+zUK3ms6CeMT8w1ionWxI7/dJe
MX+wY54NJki71pE1Si681rWjS8uDJTJqaH/8kIYVqEWexCuatm9puLHc4TxxKM8FXs2A8+oYR9YH
U+VmMRComi/V5Q+Btq+Tw5kO8pxqLmQZDLcSyi6J2DhjO4NQNpDHEt/hxy1PIjlyFJ5BD8MtuB/L
2qYhyqWpRyEOX/pp4BiRhI7zcAeU+C4JR2dNIPjPd7QFZLiVJKDNvxo3YQwnIYMB8pqsxhffmmzC
DRXlUWBjf/YeXzGCXuX9Xh3U6TNG+La6ffcOBWYe1cdRrXq8JGScJJEEDhCWe/pR2iyGCoG/4fyE
Uge6ddWpJbRVSXFwTCVqE+Kwd23BmyXqx/do21FT6KzULn5hZbT3v+HQPdf9+y1Xnt2tfOzcd+/v
vyRWX/NyDUbBCiuJL3Rz7d5OhEQoDckeo/hOdyiuDEYe7XzE63BISWBs3hwNovgcEgsQP+NK3VE2
woXR9wgUyJoYj+22wpvOdx4gPEK6lEusWK4oUtJRbOTEMgotZ1d3FAANCyIBvsDuBHCVOammWog9
C5ffTZ0kMT/iqZgcxQI73zjStIffkdAtMJtItOdYVxA1YUR3mjUYSy2WQrlM9bq5TfkDqMCaGYXT
NsDSaWTVxH6HjukRUERtUwZ1djjLuPUWWAmTZhyQDEcGhNguqs2JvApJvUi3rAQSCWuavQKwvSPE
+7Xwa2sdgALO8WM+xe1wBlLVhLCdV7bECSBEBEaub68GfrdD4KX6rYml1OeBMEzTSwxtCEErKvx0
EADbyrljcXFskSIUIARE9T0aVZYTUPNekLZXAZQoPRp0GmG5r06W+jFlSBlkyPVAuU23+mfNh2Od
Ft8MMCzIWmQr+o32k5KUw5A3I8D3qxWEgoEzwnHSzqSSUKuQRU4/XU2sEry7tKnyIN3Dew45Dexr
mat1a5oV0DWG9ewRhuMi9IGrCs9POiso0oyiV7gTrjX9vyc9KsPHR7W4bQH2yRSmEpn1JHqnhmFZ
xAcfgoib32yLVfgXcZfOiN/y/1xCLDDgOyuVsaT94RtLs6B2umFiNK0os8l+oDfVfnWtKnrzGdUy
otBuvrmZCqXDxoMEjYYYiJQWK/nsEc6OoPCz1ul888IvJjGjwibID8/EkICmexDie5pJqf1RhKFV
zGsRY9B/COGux0zF+fJyeVjRBa2C+kAT7J9Ixg4NH7cVPuX+7xRrLVnVx7oCumDWpCDC+EY16BMZ
TP2UBg9WRGcDpjyb8QUWCEE9PZ4owjf/T07F27FzISpiVndxselmtrIdHciHSw4jZcE/LAmsuHh+
x4kkyThqrYgm869drHe7Vt4WAIFWkrIhloDIhlMc4VSYIuheUcCXCr3lJ+wS3oOAh7z9G1g8Qpfn
djP/+stoVBVw47x7IVETdRMMdyTv479qx04MuMBViy+1xivwEax9f5qqkkgq0kcLXtRt8NRotL39
deP4vtbXAAYlBpVp42/OWuf5RqSEHZuLK/8ITJaIguYlWiU9gZjO3DhTC4pr0R9OoA2oGVC+Hnc0
D5OqYwbdo7kzjC+Lp5/DmFQYVuNNEgoHXIGpk6VHbzhOn3E40jp7Lu9qF2DRPsOu1KH9nepVWwb0
A2oxzQ//HuI04E2Pt7R8+JKjwftVN0hfr+VctN371o7Wb0jN/JHisyY1sssWcl8stSOlYkiRBd9o
574OWMwFbnWHe7hZezc0QYwuTx/3pIVvVyETHsvO9Cka/BtqPkPh9Lzt9TuK8ccPg2Qoq/KJ42fk
qhEiHfvEqNnOrrBW1+agvZ7mtasbog8u8bIljhgwVzfQHhG78ttJ96JIyBDOfsWB/uolXYFrfNFC
WkvoceQdzlaWMXh4YQ3b7LWA0uLvuspMBm68AmyspXPKizelKEIq+FxLT0O3+P1uo0iSjyuJkkQ8
pcpbKVRjN5F8/TATROUKoDDOyITi9bda24jZzaCRgWHP8qwZu/+VdRzDT5XvQ4WhHq8ZvAy55vQd
2ai9wg/UXXpnJ15IrfL7omkCzsjnzMDd5WpqvSWDGrSnWluC9YY0dCVp3mmSj8CKd3xEht7zfNq7
ooFgBHrv21X3fu4izWak+kM/MyUjCKG8aBwwy3htINKVZR42G15cfCZPyX289bTJk5eJUd1dol3+
Tx6Vd+qib/X2liGUFut5GHX1pCWJvsRgK7nngT7JwUjakf6VZUfpW7y5mfmlBL6a2W5TJYlVT43o
Ih8VHbXf70JP0TrSK71quxkVDNtLiSdbx88CXfV0kGAR5uO1vl79AEnUZuF9Vm+uF/HF3YUj2PvO
39/5oNL4ypUu5b/lP7o2xkT1IVw8Iv7nnmUMBxPCFz6WgWxTilM5kf2HIUNrevd6WRSBmsN1265w
kla3l+ejuHoq3EKurkjhatGqOodGMKAVVIULFcJ4Vv3m7EI4rjTuPS4rA6kaCO2yKCFv+ye6vZsf
BflDnPJsIQmAAFsEtIQB1JGJWAzGBaZRm1gQBHisauGSm9vNJULNY6iD4IdSb93sJq1muwtgru2A
aEdJ2cCcx2ylIHiuD9Y05DBqEJJh0PMz5qL4bTiYilmVixsCdLFpMmNAPKjaDQWcuYcDhkpcobLs
hiBI6H6vjdgRKh6RTyoAn9OyurKoGPd7kOiytFNuxDklvn9kULxH6xaWW6UZRAyKh6Y0DxkWSf3t
KozVrQ6lgBW2vi23A3hREuuxkivR/3xim1qkjVJQIMhcbOhT+kh6ydKxfk1DF8rHrt5tpqb6K9A7
VQBJA0y0bJGKP+BKGEkkniH/AR4F6eDGAs8Ss8myhEn01I7x7OJo24GqtlyLkHM4v/5j751u8gc/
HDlVGbckzUbP2CyywSLG30CrGMhTHvNDOXSw8iqwGjMB9MZuaY6Ax9qzy9UlnZAwOW4xoqpqZD6L
WwQBOM/KHXG0Lr8UvKgu5N3ZVV2s8tF0Z+r+SYcV1giC0QDFWSQcdVQvY7FrCjLhoLxpQyNBXv/G
zmhrGyrIAsuDwDGfJQzTEK+2UfQOaBClEnJ5ibt0zRBYbPYt54O+48Ct0VM7eV9lDqZlQ/5GP8fM
8b8S6frYI6nD5ApQ68hxIxmgGbypjOMoljmQiJUn7dUDMpvs+NzkwwdB7ahcUSC5HwUusjplhwHs
7MFwJ1P43IAEFoT3tkGsKG9FqPoBqkx7JkKIr6XVm8EKKQ4pv2FEr4f7+pqp95GHOewnr6gOuZDr
qVcVTGqPYOD1VIbHo0Q1iqQQA+hnuFBQ7yAEnS7LcLyCJUfN+P+HROnAt/k2VDW6WvV0ofjAjBUw
yJmfektjx8KRC6YEpUoxPD/v8AgefhjUU0ZliKQD88pxqLzsMA8odmBAzB7T+/EDNZTqIM053mD/
5hcasuEF2TSZ9HNBZmhJTbhcgDXX/CbWhCoRKHvRg5b5VchqM+hbKGy6A3Jaw2fAqRD1rCAi987t
Uxv1vtNVPKVGB3D8Sm5q6PlzbcvuMS5JQ0zqPk1ZzghoRGbts3s3MxkgRdJmMnEqhRBaeiHGy4O5
uxCN1fymhXy4ruTGjpLV0JRSSJNnX82WHlerrQKeL2Z5YTwLyrng/Ej5Ou1LdWR7mAucA1Dmt2N5
1IYxND5N9eQIOjDTvwrE2CIv+WjVqaVDf0Y3B0EuXFd1/UZLRawnPSqz6OuINxVOBdSzxjkK5OhW
tD7xGOVl2mfErRmJb5Dm6XVX2yPI/++sNrJcJNRXUUdTgMtyNEGDJhbZIw/L1iGZOvbWdYkQ5rlj
6OAHFViRl5KgxhsjxVb+2MuvEGmR4zvXT2V2cJg0eZ/cM1xepaBihtCAvHIqUGNpD4DYoXdrvt4f
O9KnvfqdS7IPXT+H7MJ2+qNIKzM4VxoitvwZm16ZYWkUK+vvvdIUm/c4bWjnUNEeMuniSHnXhYRA
WO5Qo8RlbopTnFKk95Yj4sVY0CaRlRyy3/LSH0NAdWe3YnhDVBiKnYRcG7MaiCU8lsHcDyDsYe6a
Ips7D5Ca7sjIONKm5JMED7JS+TEVbSy7ltGpPdRlSCP3oHAcai9dMHb+LdeP/j6G7GvA+wQ3FdnT
ybVRmI63C39w3w2rs29PduBqYk4YOcpGNuUKLdPNQasOX5XorTe0sG8MFOo59IHne7Wio0WTiupS
jfy2I8JsIM/nqmAn4+hHo7rN6WAAgIR7rY7UoZUVl0ZqxUXQrGMmQyy5Axo0Zm0rRcNiGlZ0F86/
9ih5BSKxsQqM3AK9DGGTKALuWsGV/dM8U3NsZmxhrOm3ZPT4O8pZfr6AysjG9crmFUwGWrEFY3KH
hCE94fjNUqdHEBjUIr1cytzKMPavwsQCv4pIZ2deQ6QoX/8icvi3X7bv66r7UH5PqC4mYZpumv7a
BfoqwpQkFmx7Vljcije7+RIAwgspNTL9q1OxpiNgOUg0AWnGuE+J06FuPmdxb5pkUbxA1cP7qR+f
JCrtExaRZY13byp+cFpu/Hm3YuihLWp0Dht3YppGZnA9dBnqDbwOkrEk0KS8GrzjgijnA1ReQCSw
D/ePxEhHZVKAAPV/LNY1tHvGjlSv0ASwf2vd7aB28BUHaYRpyRfzNrRO43DbpgtCvzkEhvGdYXfM
HQ1yQz2Eljc9z20nsMVwTlOqYIHZQQlpwWZpTqr0/sz7ODdeO6p+hUtKJntOLCK3ykZrUNUCegju
/xoc+2Sh1aBN0AAS0tLmOs4Jb6E0IMUZVIFan5VWeV5vT4JGl9aqifTT9urIssaRQq2EUfO5NXuy
4v+v7oZC8Jnwlv0Yd44l5QPzoViPQ5WEI1k5lmrzXKD8GUU5efBoe+x0C6EmuGpSP5tVYkv0WcIn
lZpU3KiyY+qPimrqdanLbTQltk5UGgbcf8ZdfE1EMK1xCbGpNM25j/Lo9Q0/jgdXJ0nlF4NjYYTc
9Wt3upeELbA86JLD8YWQJwgnr+SgAYbPRrmMTTiLyp3SfgP/LK53khzn5AAmQIoUA4lOZ175jKSD
Y/0wsAPUR9WdBGZkuxHEJd10VHSxhILCZJOZ+LteWaFK5eG6hrBUcn+TN5Qz9JrBxFkke9euVYlO
iikdSSR2IPTx0E4pVqa+tRAlfL6bGiwuJTW6RCVKHnoQXMpiyZ/NDDBpSU/EaJWmha9PabLDpv3e
mUWdj9kdi2K0P4W/s5SzswwQHAlBSzwMY2mNvLUxs6q8HejqH1db246B4vWm4HhHUg4EktqaVdED
LmJV6nC0cVfXjl70Z3elB/8fqPSnYPMcbSNTygNV5lJ+P8Y6JYFBuHWRJpgsFULAn2E/3OgnPzCw
0wkWB6KxsDNPkxQCgT1WuxZU3tp/CksO46uSrcIKrasQnXco1rd9Q3J+FT5FIvm2t+R3Z3AmLwMT
bWCYXtBJZ+NC88gnS7np66n4jcVKw2oV/wmoQRKoFIH4qtnQpjB4S8RKicBI532Tu4Jdj0dSkQBF
6CqZgPYp1r9ukdSOFzj9D7Pymg3iIWBx4x+MAJc5C4XmyZWzF6ZypEKsNANtH5BPLIyB9oi44EpB
cmizg2KsJYaTWVb+LoGxuwxVLrupc8E8y3cbHrQc9UkjPZYlfCfjYP2r6d3rhu93yvGzNEggqspx
XbpEnts6EQRY/TQxZz5eWk6e5oM7vzBSXwcwg7eEtNDeO10kzr5bMi8Py7SPEgmL/TQaBUDXizFd
aSkRLBZE/ZRpSAa7wpId0y79HbvoDoljO8QymnNVzG6kgsJ5rgZ2CaKGSx3O7XoYRE21ydYSSZ0K
NnOR0Jq0BEz+C4ildNkinhdvPDTsSe7csIWCLJetFTJ3LEisMYP6eHRKRh6yGdNuVe1SVMygWRqM
Al4a0e8xIxsmHYMlwlt87eDRAJ/hlJoiMTPz0sXeKHjj4FH6aZzycGIx5Qi6mr652Al+lAuHHmDj
xl6Al8tXSwhzZfbDbrNgeBCfTF9ZpUZ49q2paFu3ZJ4ATDGmgeIV+L3WH3lh/8rpTUhw2f65vIUB
vcnMk12gBKGGdQBGz4e+8xkxMZGQJakD6G6L1KZrnsFdcbgqrT6L+ztZ/1Mtm0WgqdBARERvOeqj
JlALdCHijlUgRFyvzjP6SRzRjAY7004RNDReFFu50KJAGWaQgO3Vuz1SPbKCDIWqd2i7FTr5gvBN
r6agk0WlPes/wRHZlMjzeVxDBbN8CFKltoP5iRPh0B+pE9GrALcs0a8nu+Mc9lX3KfWfxtBnSd1s
7xK4mRx66UbrsmE4BsgZo4QeMQPlow89u7sFyXCmrUcUyfGHNXlfu4lzx7lChxjuUx0ArMT8zq+D
j6SHeoNs844nqyQ2DChKDQ2BtdhiP6reEPjgyNZlUomc0+aOnyc2qq5TnlMC7wXUJ3c+iXK9hhfi
xzKZRo97WRrTGne4l3QwKxjvZTGAyRNwZubb+xIEOstdeHDyp0F2Q3/YUhwUu/l17rmnuVomorEm
wn/TwvXdGVsNYtbU+G0WyEO9FTBDkuYUOi+cOq6spKgNGBKs5qLeR7+UB7o2yg5OLBrL/Wl6kVhD
LgrmEd2OgUuvEhLTPBRE6FxQt2vdVroTaGZHuDnOZaVydRkbdLs9SGzP7MlBajqbIDTJpiisk2iJ
jDV6sTB8AyjYVhaHsxbZUEzZd12bINjXPuw0jcNiNQUTkTDaDCtbaP8DRO/tr9waTDcWX92o0tC0
4J1+gz/DGTXu3st4CCEdxzyDFd7r7Y0hCCuyyHbxUGV1/m2ebfA3kHAuZ1+c9cFQ8dMYMlOCkIXg
+8y2JjXsy1Xpt3AtKNUwmulaBPsi7xnsxYKs+0xsdsAKXsTzh9c4YQAWEN7ldeCfFW6YAPDXKMl3
Hgi1xvtXEOq2rSKzq/Fnk2SLT3AlKm5LT8VHkz0Emud8H6FueqNHSZNR0iTe/PNGzsoTlcWx1UDY
vPm6hPw+UPAsjEfa0ufNDtIi8iSSuv7odwe5b85mkq5rfW88eW920eMDDW8JOuDYkmfy4CTufkP2
tI8DuvP4QBB+PqaQeUxmC4za0ivJK0DZKyAz/I23LZdZSTDOHlDb+N1DjIBEtWdaVk0LS7I5M0gm
TNAz+INo9XjW5WtZPCzQ8gomHpNuTYSqVo8rSFVH1TX1EoAUH35VMPZ7fc0T4sFkequgThDYmSCO
repC9Ma9St5DIwjbo2b6RiEvzqf67Aw8M0coYbbTX6ADIXdUpgqFLr9cb6nMCA1iXZgDDenMUAFe
ktHrSpXf6Ei7KiIrBYA1ypCi5d7VctLnj1klQ71VMjPxEmkSmkXKVHEn5OihGgYMm7N2IISpBTkf
RYPltHqEcvQ71HvI5obIlbuP0NXA3qVTtR3kttsv9uBtpaLwMmcorgp0LoB/tvAVrUl78xF2tssr
qbAoXjqSD8IALiKjkold0zLkRkjgXhFUeHlYKl1HzT4diP8Y7+8YrMzrEwjue2ROV+NtVy2GCcxz
jndd3v7bX+w6hjCJC6lybbgYFUzr1QK6mrZ0mopOPlBWGjpBjP4b64BfuVwlFJcfPTh+fc1g3qWL
DJT8THWgYBOoqTljaCncEvnFJWcenCvwZK/38zfYohG/DNGw4xXX0u0jzf6kxDMiduIiCD9fON5+
CG17ZNcWxwTNExCNXDrApX0qrlSDiHTTLotC/qLj2M5SzhAnw6JHeRSx9iHdWO2j+/gmsFmkLe4U
mUJaFuFlkavrX9lZu2kFbXfEMHhoKAzchQ3OdYOzTQTVaeeNjPbtvcBp7mSb0i0fvuk1mvngp6jp
CO/CF60ehmjXfWVpuPM4K7egqdJzwHy0IXcwVJ+K6udiqPHOndCcgJTDhAe4LBkNTwPIBJ5IYEIf
8Hq7XucZxb33/2EoAOmIoqLZjSaCL1RFNFobM2BMLiuSv9VbrPQyrMbUVjo/0uEFIaegKMwA4Ksw
8DOuQRDf6tJUgBmN32kGhFnQkpUOD+wdLuArz0pQzEd6bJ1mFsWipALOaTDpMBNcnMOsqKKQvqjj
2SxFYN/pVf2iS3LIkyGkRyf1swUQKXclE+nUOcpjz9b/PFhKXogYzH7kCCrsLAkPPFYXQ3dUr32a
nbgc6GBd0C+UFX9t+zO+HX2/bS0yqx4TnQK/aJw8U1F2A9CC3bjpr6B2opcez+aQHj4ri22BOAOQ
vqdOKnvtwHegsoNrjuhT9PuGovokSh507wm0LiNts87gWvkA4XAIZnFzNuk08ztAG3NKePzwOB0O
H3hx5oz6Hg09HiVyllOfnASebqjZ770CU9RzJe0PfISkUnBKNvPTIiV29DBNcmEr57gLm8v202FY
ym0m6PhB0Ad3zqR0DyyMx9eus5BikFDub396jB6bmsWHtnr6sDtEAX/HrxUPgLdimg1W9si3QyIp
qv//7pvGN45JFErgJEraNPgGDH7dASMHaTGInqXQx3nyjDOLwHe2aoiq3vAOJ/kCHoYhWMvSF17X
0iqRNaoW8Femr2PJVPD8c7Zi3QvXhkVyBUJmy6hMjYGYKVRriTBJUnKrb6HPrQfincblALvxEXpU
gKEaDSB0EIQDmttByQzhSt8fBjZYHcmtI9anrNSwO0tZnmlwuDi+cWwNXZNOtnGadtk1B2OUfEJd
HLK8Y/QjwALLilu7S2FiEExQL1LH43YdsHRIqq8BqaTUoBjN6AkWkgBNhwosUxLOn2qmbyj+0Myn
MTZCkDTQj2TSQQ5hyXho2rP2wNsfjGZiuwBmDS4nR2iPQPdIQ7JwyltEoYLpZajml03FZ7GHWbef
mVuBonMuwOg61cFFkpIycycx+CJ55IuoOzO/Q/oNXhGcC41MjuMrzswZSu8Ltip7trJ4CYrKdOyj
HSjLhbPz+LY9pcXQ6g19qsRjrLXldpEZoqn56ubbwvrh0m4xCW5KJRVSZAWIH2x7JpFLPh3vQwQE
EGZfyG+4I68UYI3estCHTk3s9IKI1NH1nyPonSOVRGbzYDdwb0kI1by61ZlyiXhVqCokasbK3APl
0bLKRR+/fId+MQ61QKnCC8dPrWgsFtKNa0Uu4Uznx0HSgK7EYcXXIJKgoviKzKD5yXH0oxs/YMey
ULMXAUWyyTOexQyCtk3pSI1lOEBQKf9EceRoGHtYRrduoTYGxLVVWGZn/xBCufA7jAhb6XZkNdtA
ptKNMvsmUUSB2EgzTT/6C+jTvpQrvjR2K9iIqu/U/v/OonNR4pSr8p1OvPFS7jtgkoJNMEpe3c8Z
hWnTcR+UL3zZvvxN6lho09+OU6YUkGBaie3dnT9/zPY6ZNPLtq/bg0oc62pRmG4DVWips9pW+L6g
4VKYytgtqudEA47MZG4KqiVfplG9Avds/Nw6TUcPFjdoYkoujQs88A/rQwEsAMQIq+MH163+u2RZ
H6rxsMx7DbKB+wvFvLTad0GJCcsv5+NOxrCFOPV8Sa03F5SlQT/5Zqc2BcAGJOa5QVphUxaFXQOP
PP0hZ9REeK/zJWYf68JTmNrGA3QrQ3OkuSARNYghkIHdBXnZ71eWV7IwIC0G4d7ZlThcJixnNb6X
TzO7Cf5Ck4NGZqR2AHEFWbTxZu1orpNqzKnUOttR5ff7TrwnzMKbKsfANQRlMbANLOaecx/twETq
uHIlq8FEeu8ckiR9S4aKPazj7d/Z4K0vHncwusa4XYBDVCjFRja+5cFVNLMI8aJl1jtn2omCQIz8
MnmY/6rvHN7HK6Buz2EWPaFLMOUa6U5bulBuk0nQdJWshOWnldlv5r6VjcjGUXNntzYro7wna7/3
KcjDE8mlhlRCwrdVwzwCM4KLeReuGRn0qj8TquHRbjl53PU0D7QvGYwut/BN9dI4NFEP172uwDuH
iucuo4r/U+K8ZfnsEOdx/QDXAiEL2ncWCxX85HiVMNTfCNgVRZfz0fLw+NZjmOcMUa3CJmYVrrpc
ufq4+vXabWCAsU3U41AHGgngyyAPoZxC/wrgjJTovfDVaZ7FjgEwC5VLDM/bDNBM/BDWNdteGQFO
Szw1IqhpaiCfFjo9EWBImBrkWhCab15LmzN1QmoLCCkQmgrPhN0uZl5++uUU5Pi9t8uCnR3/RHAC
YyEXZ6Q5uTuieXxZCOoR+I0Pxg2udEMh9JtcP+TYRaY8tKoqlNkRYuovNxsf3r5rs+JgN2DnzcOi
sSGULD9qNRxCbRV+sjaLFWj+3+cmkKejCiFcte6nqYcXi3WOe4FPMK81Ax+I2pSqutsgJujkL/le
0tHbGxQQ2BL+hpccjzIGUqVuieotIaSjxB9fjDncPL/ro/bSUaiX1K2tx+amizkNKNjY792Tgg+6
e7mv7Oq1wHjz3zD7qRM5o2kBEFYklAR968lpxwe9oVm3kDo5KXgey8wXJk7N3SmoAjU0MCE3/J1g
voSi1w9FDYEw6iY98D1+oVUEFMipw2WLxV+o3HEAI5rhhTcx4/ExogXDDRzldpsPrLTufxYXj8j/
ys6dbsc4w5Egd/n4OVnIcjHrXSQ/qHPGM4gVdEaX/JY//8jxDiFQQYV68eX6a130BQr63B8FuxYf
/0yM4oEVuuWoANGTcO70Z7HopmY7QX8lsgRhIRrd9BRa/IWfShkW1H4DMYBgjQy2vIh7JmEZSY1v
p+tHIPz8Y5gHFjRun6363rv4qJXqB59U6ZmTzDgEm5cbELRwOSdcR82O2fIBH0b9SxEgc+YCftcf
oz8/9v1UsSez7wIi4fmks8XiNqgPJXvgaNcaSdq2M7Lp4vWMEsDy6FAFr1Dzz5wF0cDtPhOXNwIy
COJ1w7xU1yHIl8IWO8MKcmWDUesRzPAsII1SxrulNitxUpKuyPmEGkw5Yj+M+Ezmqx8cCzykAICz
Dn+iHLpU5n8+rDTnhS4CcQSaQHTl2glcubddDqPpePOeTFBflaWvv+pmopK5Wc+IMx21Fb9n8XD6
r5G2Xxgi1O80AaJGdmM3EcML08zmJvG9aw2CC4xTa69F4klOhHXKE5I25iDABAoOH29XebvVAGxY
w9Dw4lyc6U+MvDTBXCIckIpgw2PyjRCb2Zn+S/DwVt5JGQ5XJ/XnYdaXnemWILld1JAl026wP8nt
j4a3zWaPvE+HTb+FFsCBFvLQz73aF6gxp0eX+nRVH9hQXSdoVbj/jEmcO4MaafQ9iS6qIAQ5SV5e
IfW3b/Uk95cGcWjPqGhsCnKbhV3FSx67sic2FsZN27uIaBxES2mXqdc5gtrfJM/IDcKKtmJ8GKuY
UxiQdRc9XwpGQmpSsP7thSruRoUDjS1YJrNk9qAq9mthas7fcx/TAQZPdNN7PPR5caSd6pkTFpEw
efl5QbpfRgi/OFz7A9Tor19Y1WD/PU3LHNq/WjAvWxg5ERA7y5Yb1ZYWYQ2tS/x9FVQCPqdJhElK
+YON/554W77mTmv/GFFuaS9q+JAnO4kwfxpbar8p7uiVV9FSK5iDXP23eei+UZ3ZIvq+df1fQoCa
x+aPl06x2Z0mAfxqqMCIeb2k/r9qDMHC/pehKDlecgCzcudR3S2k/2XfqxKYYCUsrR7CD7GldenK
F9ZgOy2sea1R8Ui8lgjgizkBjINF0XWB5FdKIY7clJlffRGjhP+iDLsFMIwHRcnjBWg8GRNC2ERB
l4OIAuuO4Xnhljk+xNhTwDYJ862j+/QBQm/2Xc5u0rFSpNDrqntW2ItYot6IcrQafd4eDrQpVTz/
eDyn4Wj9ASxcdm08BZwa0WzuutM/OLDGv2TrgnU+m6idj+njQptEiUsSucvjxp9kWVVZ9ktq5/gb
KQAPaWJ1yM01Y2JUncJzc9s9j3EXXffKpOo0/T3nYIqpEXhPynrrGo9TFc3jtIb8XwMU5qfjzS+0
EWOcDAx/9yxcf2f2aHXmvCtF8AX7WdLDycHnHIGZ9darXcFc/VvFnAfP3rxuAk4EOeJVOWwQ3U6f
TnfzdkAbkHoEpQ0Gs4uieOAwRqW34zE7b5FgZmzNUd5exv1xrXrn9EBD0yLlmv0gme3tKcjSDrFM
1LEqglr92zmM0Vlbl8DQcaRHFAysBI9lvkw7s4XcKyAuHC8VSr+rCJuaGpxj1NkLSqF9kLaR8jBU
5OEJ3OtAIpfCxnmrIFMlrbD3L90JwRA/J2YoL+YLpzLFnLKIeanR4mIrQcsMUiHYM3U0uwFuhFBF
NA/5AM7P88yyqjrt5tnsT5VageAYIQ256/tQMppF6cYFMxlDhoUzV2LRGfKqECAbV0kf6SsQK4L6
ml8290cybc2NUn6xqIuGLuPySgj/XUpRO4rwr7jjKXmj84p4xyT3OTRSO3CcP/ADvHN7nu26xYAZ
yVIYPOPJKxsd4l5Cs3qk6R1ANrmzHO9qP9prf4YOHL4XKYC4Y8GnXrf5Nw8hk4/goGCygHpQqGHV
O3qPLuD9+soP6JEpv8kXXGkJnNZSewY2TuFrLSAP/fp9czGy8sq7sJ4ms9+h59X3vQqHIhmDzZXa
GqMcoP9NHLbouhwqxbnXTiLIqQXglc5n9i+iPVWCaKbsP+9VokEyRBOT5JP2isL8PWe4Tz6hBcW7
XRHKJvekSOgOb6tN4Q651FcU9aJ/xRfKsPhGoGgMxRkEeCAEYoJ1kMlEx3GKcACTtXtPaPenlNki
5hqI2fnSM1GCiZSa5RJ8u2Hdb8phwaJ2Th7RFH4Skxffud0MRLlyHVd93YRW0GeESd+4GbxaGUyQ
JxGirLEuLnYmSYyFxhOZx6u2Hp+Un8x2JyuI8MGa0B9tvtAlH0PmzmdT4B5sBfQkHEpXgglfU2qP
+nqqnLqO9yTzzs6EVc+SX160ewIyaq0PmS27focQtfDB8PPvXvBC54fDp8D8vozTi0c2fGHEw3Dt
QMmzWCbK96P8ik04xExX3fQvwm3HrNAp5KD8+KSL+ZOLqZljpHwvmBa7WKat98dTZUe09LdadjoE
u7Sa3uCFCyC1AfDvL5GMJ6jqaQAHeteorlO/ZEFWQvDJAeqoCGeTHKa3wRTMMP3Fw/aU44pD/5y8
Udof2AjdOQK8WTRcfa04AmjVdTNzEny4LgCZx9in8xFh8UOZAUIDw93Y+iKf9Bcod9HX0AFT0Zy2
AGoYkROyw9mz9uK68aa36Fm8vVJFRvcTBaVKABgzqBKOzUouQHp4EziLxQz3BoJEe7uj3LQljx8H
1SxSsEUUlG58eO6yp+R+gSftYxrCXcMWGganxViJHpjBFoF0EjHGvKBvw+qP3bUHlLcmHCyuWHoI
ceFnCBmGdUYrEum0vvIi0eq1r5cBlQy2rwLF1KMeR/RZ/mQiRi3iMYwsMCb30Days7KwztwgayYS
lFri6YrJevgzsmd8LHo0LZSPFTYt4pUmUUnkGIjHET+XyTGmRIa945LyuBBM5ag0SGARW+5ciL3S
2c+nVXi8QhkRtogfm9pvkMmvWQ2LlmbBJ5gGw4jX2o7+5wrYLT9nTq02Aph18aEohB8Vgm954oQ/
AnR2puyaOGzbFjYAhwu7lb79B1+gGTHcZ9gEbRtgbQQT4Uh1QYSe+GBrQOHknqleFMYcnKz24v0q
dx1cSxJFNl2yMJlnQQ2iQ2nmLhQoj03BRZ0EqcK474ZkVuXcNJRYGxsE8FK64OULed+WtbEMQ4SV
D/jQMtljB+GeCC/EBIBCQUbuLhzYyiV6+EIfF/GAHisCG4xM0rmWL8aiyWqshD3V3ozHGZhwmlRN
+6lzHS/2A1WoAgUmCVdGvWm9QgzBf9UjTU1x/Zawkabdy5P2GizvsJbEJw3F7mpeCD63XXWJ7yjH
VFjBIROLv005yhoXLyllocvhr1zRdSyYJg3fzyfP93QlFsFNzWqbLBIhYQxsPJHDOnFpOClkN+DB
VwDWLmHVdvnlhXewym114beR09V6d6ZHcBYPmVscowe1oDsRr6aDqdh5dUAkgP+jWQQAS2ha396s
2UosK07Wx6ZO/dkSqvPPxMSWAnJMZoi2DHrGllH9ANk3jaUFtMlgOQdIuENVQf/3HDRjXvw2+MK2
MSmlTObdh3eroAqZ7eVgKrhg8tcNxQtKtQnhlLKIoSnH2AqJZ5aGLKBFGdyjnBOwMNK1lVnKObF6
qj8noFjpvo+kvorm/C1O6EvOP8IsrmkOeB5UNqsebJUbjaLNdLX3sMlEkQuvY6Edx0uKsU+C5/+Z
o5GfzgnEDzmQmtmEG10npHsftad9rqcK9jHbZm6B8I9IDRPcd3a2GZtXEvhQU9m/XKqsvtCv66BH
dafiZTvhgqruCCjDAqFtzQVLFAFHum79w0NZdzcsGDZ/869JyTaWOfIGAHRGCFT7YMP/6+MwmTto
f70960pwii2N83jkWwIAYogxf7Nj0nth+YvhKpXS0f+dcNV9shx36TEqZqju0oLz5ug4iLW5s25+
VG4YfrWSmnnxejH2N+mldoiNtVusf3nYL6q3WEFN74S9XpkQV+CVHn/dY4LQlKO5BLu5VExXHgab
2DHBqSOARrF9iqBJrTyMDKeo1+9PC4HwWBdk1vfFfOO5uofhm2kN4We6DFIq7jVYoVxa4KutkOhF
kBWsiRabIjhrIiR3ybVT0YsZCqqGXCmLccql8QLSjEBw9fRU+918Ap2q3ZU4+LSFRKV+9I8pCaiO
IejsXmkOtL9auaiTHpMLkwUvfQ00vQjS5ZL/bAcfbvJZac5JkWCe31u2dK+gvZzhAXliOJN8LFwl
TKmwlSXS6H/H4XT2Kz64GTVcCk6q9vorlF84QS13eIYmdnuW9By1uoZDrK7pzQ7NLYY12P4GI2NU
9D3A7w3+ajVcfD5CFtyE7rZK6Od+Qpf3qaMOJJSJzDiQMlfo5q02cVTFperpuI4P0KXESqepDsOC
HeKGokNzGwgXovty9jOXkXnagN0gTc8nMwsRfGFYJU7mGQ2gFnktuAhG58uZW9hpdQGrLMG7xUuf
NGXuTvJq/nM1BPImuW2gSAgwOHU8kv4NCOxGY0LS+MlFLK2QnZeAyb6A7ktgHjQ/hAIUk3712wDq
RYMz7YxKHsTDAE/LMrZb5su5cvYAq/5MWQMoM1X0lIqvhiz+tTUE5oc0Sce8oJMP9A339Jk7x2b2
G/ndCY/kn8paMr7lxmV0c66OkTbdsq6XyGu3AyN4qYsVfn4hBTTSg5nQ0GjLFtUvOHdt7KIJx1tz
A9wIHP/79ydw/ZA8wamK2dnuG5RWK9RHd4JEcXM5QDqmwF0NgcLm7uTbWHeNIhvFI8S4b/PJdPoR
bsyuJGn6MRp2FIac8alIWRTcf1iJI9LjYSJhQPAFFbv3pp0zqfzJo9ikrvShxF0Y2xSFSB9DFpYx
AAuYrbicWnYhaQqXa4Roz8alMofZouLUnMoDT0BdGNPaXDsiVczQwKz3Gke4Skn7qv6qdaH0Idk5
0JABZkNm41EWKKuWYk4hAOBaNDzVqeP8EjiGoXFU2Kv5cKGFoZRdxK+oKZMtcqIDP+G7uve6/Cmd
9dPIhtnjhZiUkwgwBou7SpXFfQaBl0Zbc/9MzjdnNDIzlclAJJRojeV+zd+ng768QaFdzQXHI3s8
BK6OhC6kb3CREQgzOy1OTyJewkSG8a4UzhesxAUQCFdKBGLHLfnkqhGnBzwqIqFfdbBBT+VFPyDc
O+MdSehPvh0R9CyDSpBtMQEtVnWj6rmctERV49HRNfn9+Z1VYlRFHI7rxFg6gj8Y8eH1KRbx+D7k
7PTtAfxcvBJWr8PiWvvOBg0YEVOberwMKcA/uPMsHvIVpXWU/1ml10Nq6F1mncnE60OsF3Q9jh8L
ycKUOz4p7sEc3NqcZmQ5fOFGiVMkEQXk5q+JRLdaRP7jS3ZUZSQboiw8qWfQAzyGco3fZIdVxblV
e4NHSntwmrcEWmxN4saQdrEdPkNZwIXHpO1VQt9kN1Ldg2GZaqYcV5xXusPoUHntcQjaHuOh3k0g
vzVCIiQPfkqTTFIQyRFmed00tVDwJK1Yw6IolbgVAT5KQglTY7CYVP/fhG40MCE9Zqh+iZ6/pzC6
OzWdVIappzqY5d294nqWZILZ5X55RXH2bKFSq4CRkhPwnrbXzUHKJlEnmTXshOx5INW/4YdkpnY6
RwM44MVoZQLUNfKT6sLQZySUJ4tcYxiP9a3xL+6HWq+olvHeZQXauZTIkk29lwIhAboAeDhwc8Ao
+lzlSTS44CbUfG0xQ9qBCpKQ4XFrU2hDc84f6us9JnUtqSXO8ZKhZBaWb73GBMmKRuMs1m2CRX/q
Oh2xJSDX1WQr9H4Ty7gPaLyQXaiTpD9MLppvVtGEYQI5kFK9B6gusAQ1sGmTuxBLtfa4r4MgATOJ
tWz0c48Dym6O9FLJjV9bU8LHy8tLsE5fKTw67ZVgxZMs9ciZJMWYaOYDlxORq7aHLPYZWL9iPxOM
fpN575siRpu68ZcRyAJi5gKuhr8IwkT1c7+2s2+UwNXdGX7MVLbGIdInInlinGgk0sEfbqozRC1r
Q9yF0ROgtqBlBeSXOtRelAnpaVZ2BVtzwosTyEIgBiTVmBgByp0lk7lj2EdvsywDE8xWPkHlKmln
u176qTcyvcdtYbYQrd3swtnBX5XImz5hyaNH5pRDFd3XSMZcTWaS8KtvdKYzMmKNUWrhBbBo96PL
8rtwUdXAheeZ2PTEzr1admgPg4Bn+1JI858Fzir+NE4RKjkVesKBbvbGAQkQZklr07cy+bLqKTVb
D1M75lWbICml2bimPaT6GaM94h0XyEAqwlXdKblUoSOL+4YjldKcov5Oxk+z5gh8gsDQsH60NoMt
PJN2U+K7rlGT/CZ0kvTJfyehZKNK4iidLX65SdunQSqks0dz2yxk88+kSB9P3/BcwE2lCGVd9Q5x
j1AHaN0BNo7itm4i6dWrBhIgv2RI1ZLPiMpmzAkMvGr2zpycVi7oIFavk/HHQr9LGW+1rmcANBND
qlp5bFyB2ama9l51zWot1O2fZqpycg5gQD6BddQhzPDCkX7U4o51NX88puwImBJClMvpnDbj3usX
Arvrt8WBkufBAWreHFx+rO6I9CRexy0kYvmOxP93AgUJH+aBGEB/haxgdINhyxoCyXE0/isqTqbr
A5XLaA0iPdtIBidyZM/LPRI8Ijyfi6Y7KtdvqYDNLbc45OOAKnHCfYYDaxIeiTriEIfvpFtaBje5
+ENSGYkgfSiyHX71+mrrUH3tt5WMCQGPFNOEEfldv9Wkss0PUoJ3XCZavMZfiqQUZh5AGExDlF9k
6ydV3wHLUQTSwPNBrfRT9+Wc2jP22h/tm7jfszqa2okNqvoBETpOELIb0lPp8ODWI71fPdk7sLxg
1IdqETdyEIwVuFImnKi5x4FpiO7mk+fhk2PTE2ZvsefYJBw84zeEk+rN07TUOK7rpvf2OSb/w3uF
ZpmYc8yBQD3aaGeTfhcm7WO+cwEZlFAt33gQJyHoT+MoibOjfxr54QmZbHXVYWpu7ZwrxyK8IG/I
1AA0qbE2i1SAH0BdDoGjR2Rk+u6VGS7jmfU0/hNm+PlK2+c0u7ywLQh1vw7+hrgFoLx2GCQDYqic
4qQ5/T+nOxIGiSpT1uEKeW6MF7P1FsKD99dMtnUVP96K0Ahl4cYotneoN9ZHOplYOwJ0PnAghuRB
oQ0dS0+vXFxJVWDzdvs3N3yei9aGawtXQqQlEOChAJy7PeGxNiMW8fF1ABji5f9FKhFJCvPEi6mv
TONUqkgdrh7SYhF6HmVfNlmySUX8CLkDdxKyuyVVB/ljtySWxeFlzW+GDLopuJXycPDZ16DoB/Hk
gJKO151wpzkk8ExMm2XuxjDoS8ckTG/MfX4kFpZs8H4UiIPm1s/LS2NNWe0iabUzfN0DtyTbxA05
2NVAniO5sgTgPZXGzfBZ4EJohRImE3ghUDMl9Q2K82HQrb/o4HZe8Xuw1v9OxIJ4XdyNfymlTRBP
p0d71/kP/RztlOhKKYNDAUw9XHVhGju45kMqVNzAorSwtg9DPy6Oc2JZQZqLUfSAEm9/qrcV/gUR
VcLXyBiNufgZVzmYleIL3GWNNFYRqrOfsX9KmyaKEMogV294+rXKwVlOMcDdJhBn8y3hW2bH/9mt
zLXFboDVxaDpACShV8q/gEpu7tn2Ugj7Fyb2DTL146Qx0/ygcEEWL1zRqL1U3V6HX+kP4a6W+3g7
Yzjsq+lUNQhsoNl0fqPUuxFzaflmMgpRJZPacuxqI4DdhOayKcfXDyUN6s2QBLSGATiUwxWcQE0R
p1is0MBKNSYqP5SbRgi6R/6DnS4PYhIo/9XMVs2cNwZDuXo9/Yl03TIdccrnt/SMydHx01KJFtL8
omu27bwAwFA+JSTWszXs0pWhmJCWPiCoZFXoBuD6zBVRZzcchsDe5f1ZOZYQZoZl56Ldazyp8llH
Th0ok6XD8vXTGu4jR1KWdNlOgt1V4HzSygufTm4gR5BfH35u0QSK/1CvLCx/HRf0tIWARn25pL4z
YzLdO7rsDZ448qEcbN6O9cdQgDBlm1EZjp0+8q//BowDvy2Gbnhu6UtoECS/Lnmwq3mO++i2qXBD
x2Tu6EjH7JNxpE8Q/lCrko9G8tiMOyuTXMokXn3PhKxgKep2bbVEsnJ8kzr+TBI5ITfazD1QgnxG
mGcGGm3OAG26K/htGJ2QGOJIRhN3OC4fZWF2rmAvKOd822jTHuNMt4Ygx2+WddRE67UmWm+w6Zq8
hgZ4MJhLazLDtimug3SRyn/lV5lOhWfgw+AK8DG4T5tOtJ946yOCFnsbhajXRdpbSImZ+q7Z3MPP
pZP2s2/waAKgV2CrUOZD2/e77OF647+4E/s1l/CN0Q5HGg36uZM63BVYTmOXSmjPvkXqbZ+XxuhL
i3gRCkVA4f5z3BwPUq3bJtp41eerW2mCKRnDDftBROcfueO4Rx2Ya7O4YWUOy1T5eIWDzDX4sZc6
MUy2YuJ1HSAHK5cNLQNoTKQVNdZZqOlA0zdv7W/UqGGOgL23h8+obKr5tWBQqQfcGnLt+GT0C0LT
9brC+45bSHmTYSYeEml8wRZvUglWisl4zuN3xnMjtun2+bKri3im6TYjUB0VxiT1spLzAc8DEFJA
bRDfLqFc6G454gFw4n/uH/tCjHESpUwFUC1LhlgmHTmI03cyCbgYtVt1e3mVQX0W/UGqO0Y/mMnd
vWKidzn7euOq188pfV9KQ4xAkq/8z4PM5ECDCXsYMnIAyBvwk/WF1qOfT3fJ2vEK+66DX5yti0S+
3QRlDPVF8j/WDjuYIK/ixo0amFwCkquurEmpG5r2ysmTOu8z/NOZEWWQceScphT2Iqyu/OlWP8L8
BVUp6dlUSBGDqcjnZ0No3L/yC4tcNaxtdnn/9lutYrwwIfUjK5kDAMtGQWs/M2rGdS8e+n3HdFXQ
cIZp/T1zhiGjySm5qLsGTmB5rVWhOAr/xX4nEZv4hlL3nO2zwDj0QArs48yeI1G9lbhAizguG2QW
jeVaZrclXvnxvVRPYy/X9mC9YK5/DET6CP1j1zsmmqMO86SGGkkbjJ4qHXcvrhohMCsQs5pgoZRI
cPkNtVMRpG2xTV3irnTf+pRDFa9zCWxEtdn5fMsOSo8rg0yUXpafJvXhNP27048YDXYHjagYggZu
xpxTxE12aCkzCbeGf07mVZUR4U+Zcn0uq7lbVhcQnNxnlZcvJEAtun6SI7IUQx3DBGdEGbHPKl99
Yqd6BbEaJSqS+LvoUxhsM0CxXp/hB1l3zcGP4AlCQq5+oEy9x1YYkbXx5y4KCNhWJy4KvYXS1JF4
KG1SuL2Dv3ou6X4Wo/nSgFkh1w548TT5+CBE5q1TqGUZ6RnkuMDpF+YUa11dV25UGeyOdnmSJCJO
RWc1WFEBdQmXgxZtEMOhFqU/aZWAPNkZKPgW2MkNrTHz+XnqViCwKAJ5cOaWrHZdP4dnvh9SV0JI
sFt+4h2QQJVF94aEh+1u+Vi9fq00pKiQDeb1P9sf3QkF5hjYIQ0jcRavTyi/WVfcp9qo1z5kmiJ/
xjfj2YIdRlbbUV7lPu30MqLgXEYZnCmzMrfDWFWsXF/198DdRc41FnuRu/dbWAiN/1YL0SNadz55
AinV00g2gh3lojsrHW2RzzyjlysYf3s5uHEolLTQbW6HRcmhINbIRiEWOWjxdF5FpG4kK3xPuu7l
zQhEH+AkwMWWcqgpeiNzShdSYJfv5wuOtvgIAlUCaQX34bchskY9QB+1dtblnoVrg8FJ3Nv0wbQS
OFeMtgnhJpxgFx1gS33/DZywxhMMkV7Owry3NjckpPXnzBF0t1t/MVKLHThX67DEVTO0r2cL74bp
Ssy1DV1dkVT35K+un1pt1y4d7lFC61u6k9eF9/Blzg6uYKH6J33BjULgQbq36yX8n+iEOBuqAR/2
1TfnHxHJvhwhivl1yZWhNKCkI6RAW2wrPHnMzHMue+mFVGIM1zl6WizsK9fY9U2Z1fGYURospyqG
67+JY21hfVIQrcrnfsj2dwenp/wlFiytgNbtUSTZoVBgIxYAzgs7N3tHpGN5/A9TuNxVXzjliLfD
tFMh9csFFEbcxFklw1KMBS090yaqWn4wnH4GaQjyrTxguRKJ6ATpQpY4m5fv7kLRP4Ejsm+Ev5fz
TF77y1YFrEzMzQLPJv9OhnrwsjNEUoYyoaz+GNshPeuHuMlgtyiasOV/13HdzHHRVXxaCeTm+sBr
qeBQ/pk2LJoo0Hq/7CYywaWMBXDFGFCqeb+aLFZmcC6qk8hJqb5IF4sh7IyXvqKrMZ2l+/MLF/8y
2+PMQBah4Hf2j2hifYwrV9e0LIl0Aa5BxSb79XHgyImZm4TvbTx7zZ+zLSCtKTvD4Wchuc2NUTuQ
ferwfK1lSxjeoWVsuGvQk1W5hicN26CtkcT8XTmVMNiH83ZyUnPErdeAtWA1Fgr44TljzNURr6fP
gUsmgy1oa5lNmU886vIIQdloXfVmAsGrPiDfJ/hbQ2bb6cCbxOpeSm1CEPlbmHFHauZsZsvwd/Ip
FTwlX8ZrFDxWO1pItgd1TXb/cmE3YfMnznqfBJrqv+wxJhGK9Uukz9ZFWMN3yD5cHlx6B0Rf0+vE
KRdGLQTAbr2A+DsTZQsq6tQacx+QU2HwVDIjjlWZwOr46hsNLLDNgyqPEm2YwOPcKTOsVCbolL/3
gSj7kTFxEMECDmMl4bx28T7d5ncB81w0crrDOL8eNc0BvGiftSpBzFm11B6uILrNVMw/TYhpNKwP
pnOxT/pwxPLVjmGeIYy4DjAQ0del+dZC9sNA1H1BHnsg1NY9IWK+5D5hqZ86LPnolYZ9Q1Fz09wt
I2eSyQDIzRnI7Kl7IPYjbLx5gQPCdbelNZjBj2sWthV/nwQq1gMWZUCoREthXocdf0suFx4sST+r
6TB2oL1O2x34TDn7Usk0OgvZiqkeVqe1UtNVVnFmHKQWXPO/31NRBVOXjXiTSjvDHeAf4c1UzXrG
HWvTJsbZdHBR3eRbhoQij/JdjrVMlvK0QUCfMQ9HrPy8t8IUAcYYsUi+BwaQfKpYgpt4QJW5a6Q3
JiPIZpZlsw92U2k2XzQqqRdhM7dzYpAIVsANIsmh3fDzDpsCBddMEl45iSK7767++DRQNHyN8YMw
qLaFl9/gIM4HHFyLcY65xFi5dYjgt1OmuHQ7Q6nxfP0YFXnz6w/rpFMpCM/VCJ8JIbAM/q+O3q0v
f1ICwGLoaOzPqRED5Sjl+rp9rQYhI6+lZbWhqDJrWlY/jqL+vNvOK3Kzb3F8zEjJJr05x4xNVQZJ
rbSqgifRthv23Bzggw3665j6bFRYOjaHNNGWdpQTw+Mh8lUiJRd0jPqt1XBj5Pq99wWIKYltZbaE
+S4LoaSmxpxhm9WHq36Le9beUVRyrPtYB0rP3mv0XmJGUqYSyqCFW1cyY0jZz4wYFomrUFvLxlpK
+/aATOLaCvnYFP+NgADkSZvcQIPqeXexLSxpwLeUv0o4sxw7oPMoYNe+UQsTxRiMGxSKc+SxhrIT
0KRaRwHmH7QzXG8m6pK1weBLphryg9hpaF5Q8vUaisRkI0SJqGnbq8NWntvT+7CpyfX5nI+EpJ9T
i77YZIlgEYAvI3oJbCjJqiF+dYVVfnCcHRyXwhvF4I07pblcup7YqAdnYLxmKSqPwYlOG7UVCQbn
lOlSKT4dYSP+2rh9ZMMoCj1zzOl23LzUvhhlpKalBAR/MYjKxqEgy6g9KRRrmze7kf9AB2J8z9xF
gmyeXoFOqMtVPzNDyHLr7uhTUa3JKLvh8AWxTO9VT/gCaoYDUD6oDt5TnN4JvIKjIGiN6GaVeQBO
qgsTyZAbEIOh9ZDkb8DoZFWiBdcck1g4qQ2ElSCjJJkJScLY2hTr1caZTVYGcAH1vKDSFCnP0HvM
hGTj8mfu+O8Vd1kl3TfH2IkrjtHlXRti3fmvcvPlpUZjGOBJyMhu2C6lV/4rVboQNy2Jaqj2Fc5i
nJXpVAiY/02hBDirSIsmJYlDOWg/3cU5B+sUEx7FRx0cKQ7HnWLMPqUumek+7sEbQeTSwF46gRUE
Zkeggrz2gZBqCv+g9J4n0aKUnPrDPMC2gpNRCfCkrRjIdFncEyH5SJMOxRnK2bvfN7lhKMZRCcn+
vx75cQ0L11iM+hvbLuz+PM7e5dAdREKjRR98iIk5rC0zEOQyJ3GHlTKS6G2KvWn/4ogFyTiyYp+F
d6pCsFgkqq1abaFMDftmyGTXe93arWOuXyFUh/U2Z7k+3ZKlmE7sWycgXsX1+C9qJ5MPFWJ6kZPS
1jUR8YcC9R2yuYeVftGg8Sp4EBfnAE4ho8blQqzsEAyaYXAMW4AZwg1SQk2jXfWdVPNH1V+RhOF0
jjukqZ0pfalaJqNmRhj24DQekeXVQ4pD/N/xye/okLfByvxrsT1vidtEUGxqKmlqTWtehKsumt6L
9LVsLnILt9pvFVEYq8ugaX15MIDykHVyC/MjnzfoY9aPyoeYqqo1ACKPAQy4oSmKkBC/jBczNk5v
dU6oLk1NYucUZIA4IPfyIIIdxQPBG2GM+OkdDfnSg6EOSz9AkZorUE3JI3U+cccBbUjNeH4SmR/d
lOPN9ZYHpV/AkrThQ7yeXZTEYl7Y1i7+695+HNSlhAjfMvOCipP8mdjWnoiS47+VtZPiSen9N68J
wQm1zPSGoY/fQRguBvppN5+XDtgzVZAeo+TEuARihPdjj6CqAN4GuycnO4MzjaJTULVQRR9O+GGv
veDyh6bSlTsSHeu9sf7Uqy9yw6kvxsaMp7wRYFKxLPjDWG+BdAcPD6Wr3amrEBJ0xM5uW8CYZT5r
25zGqJpOv1pCvPCpu5yU/mSnwGDrbhgHjrOIJaqalC7XpnPWtQDtiAdvj0JwDOHOC6kM6JBSuHCY
Kjf9GSLhc/8JVVIoBBLfTbFc9pL2KoUVi4LjyPoLI99DTmyKNfF1vM/h5b0OQRV9kC12fatpWoE0
NhMFIEPdAJIQzIKHKwl5FzrUE5HVdG2aVKiq6YmneMgoJ6MyL83fIez3IDU3kZLvFzU5KjoDx8kf
NakPB2CmnCj8oll3SBJE+mZYmzGZbEBt2+e+TojOGVUdE0lyRWr4Z1vqqJ8jiWV3OBBxgDARB1ZW
9U2SELJue3uK6StCSs0NqnT6QYgNIKKt5l59W5ZomRLaNIFq+rRz8V/Z65lR8WAqdG/tRPhOvgFJ
1BnzJHbawfcTxyju3FFwngDSJvasnE0yDv6fhUDTEpv/8OfYpzUcfBNE6BJoUrh1QJwAHQjdoCgB
Smdj5k6BAqQvsWtPRq6fwJ7lUubFoNsrRr14qyUNPhDjo00ZbzwiKyDepvQlOiQFfMfxjJzkHCjD
q6l7Q951IboX0lvbw2j7ENMze0OPte6neZUZcXmOu8d6IAaSZ4ecLJ0p9/GdPU0NiuqGKHkz7+lK
JGpGnuFR5KRY1KEJJPgz4hnwCwmuBhnEwNE2906P02kN3zRfcScPewlegK6yDFUOxQ5Z8noEYD2v
msFRU8uEF4zNKbuZ65JBFIbLJxU4O8W+p5PqIFu1U5bxEAl8CUVTSz9NRifoTRhKoqZwYoQzJo7f
WQEn8ORjHiza/+w9Tmrx/DT+5VgopMQ/BkVoV9Ln/exwM3YWhrykofEq9g2ayh1iPxYQ6JGDDwyj
cyYCHb/CsjwBL2N2gx/N5Wj9MZBg/ZShw/vgXotN7TZUgL1fgDKGUreZe1vaz8fZnLKO9vNAhm6i
Yb75ATgFe71L8f+GwF3/KdRMUbwe3ZLONOCbo+nuFqDS4Klo4jDK/HFOCKjmJ1GFr/js3Lv0ldiT
e0Cpo+PFZGzJgyPtWljE7XMT2i7jrc44h7BwVEu4oc0xDQ7hZX8RqFWFag/I9NTkPz0m+XcO2syx
zXcfdQ2UB9Kd7LLzCyTHWZZeVnk2RvCe9KeRILSGTuxvZB48LtlS5iA98XuSAaEa05MoqC4rTje/
wGklaV82+yVyPbB0R7j4VkUCwOIznuRQsSrVSI1ALGHf1GU0OGC4NMGLIj0cHq00fW402PycD5Gr
36mfFa8mE9zYanexrOvxAzwtO5NP2JGzzDpkY+nKXV81+CZbn3kHZEYQBFILUPltsyW0v2EuZmMT
gbxq2stHmEOdB0206wfHy3PJqPwZXeIbq3bC1qDOSbyExwywsAjiIYj52EzBSOmDavY70syGqQXO
E2k9zkgwOgjpB6C9aMfvoUKOSdDa+TZzaDNoNffzDa7gkNSUT5RJazfPjgfRvIJarO1qGAyjIxHV
T+p7wPRIfkT9CxVB9qICMSvSV+EsES3ZCiTyEX0JHUHgZGo4jDOiVuxD3OB/eOOMUigc/WZIQ2uY
EqkHV6Le7LtXhvSVFExciWiCbu8LCqK3bYrGRUMp6tVxHXRua4WBTJRshPNgFo88ooLexJKuEBVR
XYSuE2BmGovcpLyc8ygh7+cu0Er2ghzji8hS4nTlny5nbYzN9Mp1jp3xzn4hpUZIiLizeCC+C09o
6zxH/wnZPuFv6FTbm96eW5J6swfCL9TGzpej9KbCUgeHoHVGl2TfgXN6Pve88Iln7+CwPi+ZPQ51
F0T5YGZRld36RSsC2d9gGLZj+OZRS4lhllPyFeOWrDB5JSwklhJIc3I+Y2Lc1inVuAT7Wy/AkHOf
KbIeJBp9Zt/uzAxDUQxTZar4AXUat493//4K1vLSM6QS0FTqKy5pJqgiw83E8xTGo/PhgF5Nos3K
xH3TMfgG1eoIwHuhcA+VBPgLnnzGAszIEf6anPdtf1GGAy/sQmyzY6UQk0m5w8C8fFd/3ulW6TcY
xlckN1xQ77SBzR+hjVnDYfCtOZsaFwcEbOLrr3viIa7DTJxR2zfqsXjTj0w1zkljKWO7bO+6RKk4
QHtZnDJcC4TOY939EemavnlNsdG1wEl7qEuY8x29Rf88EivJRiE6lDENvGVYthWEUrHSmL6Z+D4h
+b+vMW2BycViZ0HHWlqTsacGdPnqpoWR7Ij0GZXCmPL3qZx7F75GQI3xEYBFRDfzZVpAIgDNtB45
h28joE/UuyxMFjlYt8WaSdZEYVWfKbQmY90U2DGVqorl6DWxJiFobatwokVy7vJkoq3poRn/B7qA
9XYET4R0vMlQg6uwOHr+EuFF8BRcp7uasgwcIKMftG8biEdnbE+xBzFogSxBY8ltnnGpvTdO3XdE
iUo2twIjNXs21YUvkDmNGPkuq7Ngip4VrGxyKNGnU/wc9yLoU5/D5Ea8WoQxm6gfI1BKIX6lxBGp
3dC45MvvhANSLSoPpoCzHnq1x6VsrvYOdvt8//3BEmS8jLgXQG6ordLCmbz138ArPkxMoGDtL6IR
3KuHuD+MfvfpzBfFlEWxMfiyP8eIFA5hl5ladAEEw8fT5FJdt3LtyW+kfEUyMLc3AA3KHft0dwjX
Qo0zXpIPFsl+IbmRmhPlPefimZbdtgxqqgAQW2zYXKxJngmkH5ZSNPuzVPbVJjzihGSDzlTxaup4
8lBD7E1MJcHleXWYmdBhHhQLn07t8/brySYqUdpSk2JOf1pp99ifQKVJF9GOYrz7VPTrYkw/w7Jn
4Ttarql1LDAk1TXUgq7A+6exfF5hvIXZkAoowd00G1iDhclJ+N6QU/L/TRBnJd29Brj4w/fwttnP
EmtzqY+Pg5LMOLrrsIifu6hxPwNbBzlSBgPcY6mgZ7lEBswD0MZwt4wm8HmucB5ilMV13ZfADpzi
vLh6PRgiFqp4A4PKA5T72+Oc1LfYoj1FxL034Lc5CuJQ4c/DlGBYiaTUH5SyL8t7hd2uKHs+nw1y
n2ra/yLLI6nSp90KQP7G5GIT66k3SjbZiBbve/6FoliIWun4XISZCidQ4G2/QOIxGuxAlsuiQYdU
v+GMsly8UGicTHJhZDXe3JUz1Bt36uADZ9iBNjeK5vXcw7hr7+dY+Mxz+TZP2GophI7xrYS8gTy6
wqQVYCY+CmTlnGgkgTDX7evm3y0zEaJ+jFyn8m6e6SCSB1qGFOw2aOCvoAYF5ptNaPZjL1hbZ5yF
z041v19Av6eJnrVkBw3LAidygOhmmYUqkm1UWwomkfc2QgE5NdotB0r7ktphCyaQ9IC6vWy4KDoN
IBbxUmMG5KsbbBtP5PYTOtKa22KIjBj0v4UaK1VgwrjhE7RJGg8sTF86+t62NY1+a5Use1t30Bhw
G8ECKED7zycN5/3rt2PZJwjnyT/gnzcwwXxhQ6f61YHOOYkd/NOLo0w5X9ftCTPn2RjgLvzzvRDF
773HFXvwXYmw+Pfg79EgllszOU92iYuS7v0WieqyX9rvlHyDTiANNSZGldR4HFUxPLsznX3djsHt
ACf9+KBriyhI9qly0zPv2VNk9u4QpE0gjlfsQd+Bnda6qmHmhannQpty/cb7yJXpAyG8F2icF7Lq
22YTc2QeI3q0xCvbVrO8Tsgw9ArBhDVSGPriXSyhLQlYznzRjQa9M48gjtRpeF8myfYmEAN5ivwP
6q5po2ozJP4reDPPy/dpfZ4x/S1ylXFs93wvj/nNpFsc1iqbA8DUAWS8j8o3SZV4EsAKnjF+hrzy
A0GhGrvUePmNRm2EYTy1E96gcbm3MyXM3oDrjUl3FBPBLyPDGqpz4tOIN0YhznUQUCvGk88LVyVN
pHQIHjIuIoTI3XwIWpTsGo80I0WeZaaJ09oY1tXyj2XB/0TSXX7j/Rw/R1xHvn/P42B3UYIOpMbk
W3JfBULaY3vRyolCYhjbxtUYaJYXYoYu2ACRmFvLuh0zrCrjzWkRXS1CzBDJ43D8D56eQo76o+G0
v7dRVeQM0fOr7r/AG4mk6NB0dddUxBjlXnJ8dGbnH33A8S53uo6Hya0Bo28wS5hojG4evaHPoMx1
5IyW2Qe+D6nCPkBLlzYX6vEUhlhnbiQJecqgimbeG0Yv3e5oqOk+unROgSbCkFnXyAl0Xh314voE
dahgav/MDtz2nUUaOB410SwAZGd/ijDTuaBj1XgTPoOr9LIT6p4WcwP//pdnNjIlBV8U6ZCgEOvS
kpcF9ki5aPD+BgxojW6PpVS1+ilWiNkgoi4n6WrJJuMQU8NDhemp5WTxEiZ0CkwiOLov1MQAQM6/
o5Ni4tPYLPo95Y/s/0W8P5rO0jmRf10cS/TWf0qoKHuggYXGcuL/krSdYM9z/Yb21meyo6xx62+O
QqAOFtDDl+Qybb8BWd9D3mmPFJ+aDVLrClSUTRpjgjSYm3JfuM1SE9BM4lS/EiaCKMVdtp6evrUi
Dbr6OsN+TvGDTb+mnaao07J3b2WuOVRZPg/6BWzMreLzxuhtXwRsIv/RWpJ6OfLVtNz8ijAjPuaN
FmUpQzez99iwGga4YfwK6xeuyBO1SWvrknBkDQL0JSzX3gCZXxb7WNSQyEJHJxikDpZtBDKrENfw
T5n+PTP6jpsL3mxxn2Wb4K4aGYgrLoF26ewv+f1uwfuhQQI2yAzvQCWZGBhTkeI+zRskX3p7W52k
b5XDiZWmpkFbtW8IgvQymtU7lyU280fWYg244m9nOTvk5LR3WsQkO0PyCNgbtH2W4iGAhc5TmsIE
9jeZDi5pC1Z/wkg7LmUQ0gyHc/pSiRvVm99I6a+AzKzP07Bmjabd1bn2NR9pb3HvPqWkrD91lAvY
GVC2BbXgJEYOCRiRVsP2hFZ0RxQQQj7p1v7lSxZqiKoPLxBGJBlj+KM0PO5IwppSACX/3ApR1fo7
JcJKRnpsqF3CJTl99cakOaCC3rqofnxSWmQ+ZQLdn7+cJ5YBe1+fXJATNQ5hlZ5IvUQ13syHGagc
+OllIpaPbTHw/b19kxOJl5yX9PX6PXXUL6PPKFrGOXR2F6KptRUkg62yKAR9mK/E7jm6Md3nLnRK
i/1ZKzbgRscvacy7OOFt5WEhZgNwPkKkXW/7jFpJXOxw2rhx94LFGnc6GaLNqwBlIqpm2wdiZQmd
VO0ySdln3dm5IsZ+fbecBdSEUPBGNzr672HpcpNAIJm8nyzHzcpqqVgn78FmgxpEO/8HmQ1VIWeL
M+vnQe6q/aKONsEuMKX3S8nDMHWm7yvhM5XG3ih9FlIbNiRxQZE1O6Y0q1AatJvFQZeWhWw5yxWT
YsaALE9WJWwPnMrWaovr5vclvL0rtNR71lwmWFwsfX/4W1Dt/LOxM1NYtzHAFkg+cE5wvUQtzMIE
YKJI+fB51afNphpMdjVnuUsSVe0bSK6ZkVVEnYF7IgpVM0jCEX2nOHNDVQXUrDJ+2CMnEJb/CHWx
rOzD1H1XPaI2s2EvTG0xeZMnj3cSL1ObMAfKJQjMTO8vls3M+eZvpilM6404tKPueIuSbVCmuQXY
zubZywREmkLwjSFCOfq5QW/Tm+yAc4oraGTn9R4xEUfWoBY48XrsU/E8jfkek349VzErBXvpJ7Za
PEn1GZWuK/HSek9MC9qVv0evuX0GhG6to6trAi6h35NNxAgvn2JbVqtQBE9HRmFP/OEPe9L8Xlnk
JpouRqjeAm0VgxPx/T5bMhzKMYboVob5s3euguHiywgggU1NI++vlYvNEhFZFTTD31I1DEC4/g6R
LqpWkKhBCDHA5y5iVkMG9OAgo2kewPbU2g/XEz5Tirfs2mpDX2PhM1YVb60dqcEHT9yHmuTG3gjN
LmlaHcWaBAzPe4Z+RJRty6LgkiovxvU78LmNpL45EM9DFmg9FOOL9BI8pTtJqhjuz5UcOYM4kZHt
Q1/6P995OI/g+0zHbh7WVqNZwL2Um6kO6bOruxKXttSM4B7lHVlkCUvlTm++MCPyB4R8DoNZubUg
AwSWXgdG5u8/hoQU63cgbUR7FSMSeSJWGDfe1HzxMP6Mht1X0JpJpMMl6m2CLRgeBujBnc+Zlaa/
hU25Vw41+/xIekBnkypIOoJHyU3dFJhPolleKb+OWgWsge6H/bhkhsWJre608MH5pyccFnZ1nxfY
PKy6LFIkOxPp8Cac0FpSEptH/xYX3j23sXCKAPXowb4n0Rij6n0y8sRM+A+AbIAHmGSWgnZ5LR1L
ghw1MjyRTjyaxlU6dQebR5nmGAUmN3IpGSlmqK4E4Sk4c2AP8EnUlcDssbCAGmN161UFZr7KmCWs
to1308G2elHyql5fDOSmWJ2PxX7FvUOZd8H9VlcDTH4jaHvHaBBCLsi3iWkwvLsQ48KOJ+ZIHVBo
0rEYRVIVZ7okE6t07a6A/Tc3sYamWud7BrBB6kJ5HWHwym+nHWKO57xO7ouj9NscraqRMrY49SWT
6fAE4dsf36q2voWQpNqzsgHIJenrskCTVa2QX6CEhx4KzZLtpiM/9g3PHtUcsZNFe8FCucgB699J
/vfMjGhOJEPtOKlDILD4xpLZ6RLm9n7kjF0aWequJ2SbDi7wXv+l0MrAnHNWCDC15QPB8eZB4vg+
bEiiTTA/AdoVtAcrL2u8TGp/Njai3ebVELncJ3/3ta9Z7deWMW2CnrcorWlIBG7uGE2kFbl7N5HA
5tUFM1U0pispcWo4Mhak45zr0zvBznGyAiJ01UGKSgJvjy2izMUAwgPixTZthaY5iDLZ0vFatiRW
k7zKWnaFzkRke6o/ky/90ocegGxkEOUEhtZhu92g8jdoqcnyO3HxorRCeOvHAmcxj8DlXH3EqRsf
Ia5grMJgJIsDpVXrHy/ZOtIzXQc3AWTrgDZuunUksZCrCuJK/Aw0E4uTPHg1TSQWzxJ0UmPN4LrV
5Wk1Ccnc57cJim367jQgg5i2Tu8bZhfkwMac4hQfN9MjqYvhUxq52poAujtSy2ohNDb29A9BBzGd
8SqAB4hMQM+69FnwDPf14zKdBTse9jScdeB8uYwjtL8nPNdrYfiLmgXp+K++/SY1x8vxFyZi6Do/
/YKqcu9BSMa/fOODqpe6tpTnkpWwZvVj6g+DSyIFJbXoYbiSGyNObYdaUg7bz+/xU5FD9sPznpsv
+7GEaL0DdEKr5DubJ/SHsfwgfnLzh1+Y/K3ya8EMQTaP5CNjBuvHaaqlMlPQEP1w5RAmoLikTooY
/D96cmfwGOGIS4U4q746aYL9HyHtDcrOK0aVcB7Cbk/VLl0ikJWOiSZhJr2YDEUOxt2byTupugIp
/FD1c6YgeU6mS2hnbKSmDbWHJ7/m5TsHEREyuXQ+DJtvM8soXTtysZSdyTKyivvbcAjVXwD9SAMx
sgSYJODchYrvk6SeLzCVVyhI/6nTvXMcEDtxHIXT6i4lWRU7RkPFZJaH72YfV7lJ5klXk4PT0kqL
5NM01qOhb8TUei7P/+NemYUFE13WiPna3uIovSuwk0fKk+UvoBx6FkrPwVdXkQRkVpCCHbR/KOxW
oTMCuW2kzqw8mpVVwGmZ7MPKFBnX+MkKQjNNY4/0DpSrzD+vEb4dDKKyIuhuqf1NTzWfPzAhR4pk
t7JgbpDuDoahy2kugNl62eJzdJYSP7wOgk5Bx9Nwc40Cozm78kD2PwikQcZ2LwzdPvaoY5QOF82N
r61yqjMnrJA+v9NGEeNvGNfnQMv2zOfz6R3X1//j706A8bWh9xkDHjpd644IF5mcPqyRZAze3Fi6
UHSwqCUL3XdM/Zw0ojn7WIRaFe9SnZbiTAYxQA2Pv6/+DrwHfl+c2GvR7Hd89vSZX4bd8/5ZlUvI
9O67TwsmI3yoh5s2fbFHnPwX5k8hHC/jRDhGSlo40kg3paRsj7tmsryryzUxE77TK0KrE0g4SKrz
J4QHnx5OEWPzzMwNj76f/EbeRDFw1B7rk6B6vzUBGcBRlJTP0TvVxk68BgfhUZAyMnmVe7zxunIi
9DRRlzP3ge/NI9mz3qYb8RDqd3hdSBRyGx0+UEsbx6m/Ovdp8zeWt7a8IYkiYDTiy+b+wqwLbS72
UM/bTefHfcYO2aGZYTfxNzo3DHOcT+samvI0XnxQRU8UvGUpq9A+j0/FrKPygOA5kDx6PmN+6rs/
ykjBB2K8yJeTLezCcxSEqMKkMBNHXVpeyfUreUqYcTnbWs0YnWAE1AZuy+O8zn7ahekKou6TV0c1
hfYmO9isEigLa4+eC1dovzZfB5nwiKfMbf7vOtGaAVBVRNjTlWdUeAWWmde2dccNkdwM1HroS+9v
SxgfdcxHtEsK+FqLym8ku++boS1D0WJna0jx2JlEXareXuj++R1YZNAx/vclS/y1B6JB/EFPpgdA
ETIMXXLCMXhY9/ktVrOzPt0492nQGqXY28H6TZr6326N3MrMyQp0zXH/ke6Q2S2PscgPZrOHJV0q
8geBXcmiLKG+tDJ6d4ns+r7GniVGOEfAer3sGI/pthBcvyedzEcaulCq+HDwXHooSBGlseUq/B/a
keQheKWgCcaqN5jydkjiUjH7U/xGTbdkFo7gdBhLJYjWELSlaJyh3jyGvUh0yHGuRPd5WSV/0GeV
9uXdY8U5VPFak0cv6GDXVF+jxlpfmO8zVIyjl3ERhd0MYoNh6FIKWHJV4Kr/K1SdBn9EZkw8gOz9
oB8I9I8Q0PbW7ssWgqpUYz9SRokHMkckOEF4+iLT+k4NWLvpxlLeOqkdeTth+whHa0BxLGo4uAcL
EWbJNmg/rGqswZq9mY+jUJrBn+zZlhDZJGcmUx4kMZ6Bpr28BwuxzSdHfj2KGpvTy2YHA2z6wuEN
0xtMKPxmOdRdes7Gobh3SAno+vpPIVWKrAFoedy1lVS6F138U3O4BiNjU5BRLciCKnEMN8469GR/
MUk1purY30u2JQOv4gE+Y7A9LKCSY7TuB4LexDJ2RNqGOyPvTUGR3G64HhLBvFK75wxEE0NMI6iJ
KfX8697nv2Gxh5Ffkuk/sy4t6/6mLPrtvQ0wT6mKMdDsVQcHLXKJp9oWe+lwmBxMBjDakIsZb8+C
NSlFuEOTLf7PElQFuTglkdmyw/u6YZnTGR0cadTCLLQhR1XClhBU/dCRI0lDQ072kqwahsi8T475
XABggPJ1P9maTwklcY389NqtM7xctfIqzfm+4Qnb+uZ4lBDPfXSQvfpsZot8k0Id6cZQ+PtYoTiI
FGYLHWh0ShWELqk36yEjdgTPi76ZLZeIE6mg9dhlTXfKAfhl7FYrOjxOg5kXEqVA/0D+KX4Imj6I
S4DRIdeaFDQPxGnEqNX5drggqWufG93DT8uUIdTdFFUe4dnZUd5lk5bbQGJ+pr/n+QRVvLizWUTL
nTNjQw13qvkFBgDGjRklzvsmnLI2eWLe1A1b+CQIv8h6smEYXbC/vFo7a485XFzL2iBinghDcEuU
c77CG8Y+ttelYmPriIBktZv6QqQGafaon3tXfbDFRMpMIP7yba91P1WN6pQsgavmBdl1sLl+IUcL
q0BH31cHgZxENPa5sDqShv3QYo3duJW+NpUEz1VbsguxUY2Ag6IAe7uaP5nir1c3DAU3U7DR20NN
3EjvEugOjqZYjKLQul6MjCuNd6F+rYbPiS44pRMMY/s0s1DIXgVtth9y2sBDCHllOJtCo4j9XPar
T41Yai0JkBS1C7FL0M04yDt4JApb0ybVodFd03sdMpqVs3iZZgMgMoR2EjZG+jyk2fV1bmXLv7hz
ImCfFvtwK3OviqbXox36Ttkh3ktYFgKjBlJjd9h0d9gcaGNoBNaVspP7kb8ADY0e2Hs5C2CBP9Gn
b1YTUcv/IzhxN0+9+UaMTNuOUMJz0/yHB1XMzPpVQrlOuUw0CBMwd7KQKHSO1rIfC3w8CZDT3SgI
E2a5nPN1oBa6Dkkm67ij2pJdAqqZKUXXJEF2sRlxu5DfNvkHbYFO2ktQ4Iwg06o3p57BrBGgjoif
YOezHbKILi2cOUen8FwP1PEPXZroGQscDBShJO38M/gYcRYBDOJntSt5UQhY9DyyOnLy2WbPy2eU
jGG+yLKaB6L/VDmLKYCpGHF1GyXDvfIIKJ32J1cIqi4O+Mc/R58M2aVWae6gYY5z90HzMp3hbSxF
nH2obWsBsbSXj4MCba3NUo2N4D5isb8xwSvbz4a/vHuPheMH3i/T+AFI9TJnLEpz6RwGKb7TnSYp
yi8OLED5l2esVAElNZnsr2Qrio4JIZ+jjmKMn/f67NdCgZngyOmakIei/rjArRkYneqyRIfOqVH6
wktYRZcDijkPMGvNpkDBe7ml0UWOX3PWY5FPj0Ecv5yflZPeljRP+BxmPDyI2Q4Ot0CRf6N9UICh
EazmgrpKtGE9UQxp4Rd/qCbPK3R9usIOZnj5bO9aWyRcjeQncn7IKQ9uGOjVr5XndlgQhXtOiva5
ZgIxj1LPt57zf1Zv9NQI5WMqdCPlhOkg0IzetSYmsfchmXqa6r9Xc9YZeAa/VBhzODONOOd6jxUj
p8mYT4XN7QwtLTs4UaSF2csX/wsGfLE4erFuHnYWY7WaC+coBMURu74vn12FiIKVTy1r0XlMjzVE
ZaRj4cHhLL8t9gl7yS9PTb04Dkg3xW+C7IeA+Ac2XkZnSFywW8CUUODofMYb2/K5ToPqKehCf0Pg
eHW3zooaX/sVmMTSgRLLJHxkym+eGihvq1GBjh412PDzV7+vOMrwm7AG7G2Pmzuszga8dEsfe9gv
BDOVFumf6iPi5H2rwgHU/luXiU8Ib4zWvlcTM1g9DE/yjTMKNE5hNzUj+AgWJWu55wIeUL10OZ5R
mEvgBqgxMEq7Xd1oO11Rr0UbImestui7lLR45sz0e9lZ3x6xpnRDSBrSe1lS8E+XB26q7zK4kqPi
25mp/aoVAC+fgOqQesW3mRVjUVjMsUh8Dx53gSGTGsSnlFpytcf1UizFyqFX139JB40twutNgeAy
WyByxFvZe107TPzKkwNWsDQkzjwO6iJfuyGi1gIz2Ny+kzBD9Mmey3+qSpJM61PqzpItT1t01pwc
M2rbU5stYv4ejnLIGO2mb5Ml2J2HSODnZCBjwwa3zvxs/A9ucCow06BMCmS6j89Z+3gVIEkMj4Fc
0KioQA6CLxtMxn8tFMYS1cDYHiQmD6Aune/Jx/db9THOdXJxxn1/VN52sA2SzrSm33ws5KsleqMp
Pc5YfQjkmYezhxVwt4h2Kl49U8VTjFH1thOl9/7hVDVW07NtcI1GtxHWx8FX2iFaQ2kWu+Jv4K8U
SyS/b3igHxJ35/GdMbUbbdlrZsndMySCx6z7+d7udLeb7DER3ZOTuckLAtXE/M2b4AVQ7Im/xIQl
Gs9GS4JNoCWQPugo+wfB82a4t88dWG00vlG5S0187T+dB1+/pgDEizQUotGZqeNVa8Xnzh8NI41b
XmTiOwNrpfOYCLGw1jGPB4uu1IC+O2MERvq6aOWH7+P5pX4RopQXDCq0lfKLXsJORHXOXXC5iwRI
iTJA9cnxrwT6v9YdS7HLsayV2FLWuz8ciSdA7pa3UrTW8iZwAtEgjj/5Iiovca7zK6LKVgDgpieZ
MwaOEtSSQgqTZaQUCVt9sABNhgUGjprd/VD7G09vaTbSE+g7QvVhkM6IFyH/uxv8ll6apqlqgrRU
v3G8wfGQVVNsNdC9hdYhmyDudHCFReVe99YzL1f7NyRYSc4EWHa9yR40DXFoA296ekDqoB2c7fMt
sxbAQ8al5nUKkeTI106xsJjf4IbzRYsTBTB6l3pOH/MlIqA2iGhaVQU7+/04zxLkQoz4ap4bKcK9
oIISXPZPAi8jq3DZK8fqiT3in3OtfIlxfOZnz7Bit+huDQmP/6VOZ2PfwqghXA1IL4P5Wo6R6FC9
LvEPMvTGq1iLDZIQ3D4fhyK0zvgdWvAbK0DOgN8U2fw4/TZeoXfw7b82lWsHfBev3MFx0JtmBxW4
s8+dgPXIwL3kCm/7Rx56DlSFVViu1w5O0XyvIkSHRO0duXo3QhvhRkaffjSy8LMpzUoyywUC1JBp
TKT+cROMLXg75MWBx34NItyga+bJ/R0m9DKTIanLT6M6mWJpHQxkqJrPKBK3voeZJxKjrMlk+nMH
g/wD8pGyvMXbg2vFseE9zBFoxwzc6Az5PBGniHApWKRUBGMByiXNJpcrUuVl6GjQ6ESCdFNjw3ss
7LCmreRwO2c+w/7IiaPdtpEYU/Jc3WrVOMi0Pa5u7DdiijPZEdPpKw5brkwD0hbgTixKUezW5KBA
39/5tJGvvfWlpT5NfDddldsI4OhS6DwwVtZRYen7RPJ52zDteATSjM/8pyeSw/n4NzhGUSzN0Lsk
BGamd5kY5Sf8hSYLJxo1xjwX5tU0CGMdlC+6C8+xebs53WFjhUCdPQYnXLW0fCDKcs+ALCn4hw57
dbeT95qpgasJs7NpjiF8oVEo9pNZJr41QCvq2KeEpZt11TzrFeXcx/ngFyz4N7jI77BCKubq3GhB
QL+KKtrvd7IxcM5S0nrHJ2gdHJvMww5pr8L1P9EoRb28laMGF2/DeCnyENhczzNFArI2ojUvi/Wa
qF8drYhbq0C8QwjMZN0NhygVzvzlEk4XDE2cqvmw8DPqei2LTiun7CO3fvr9qdmmqHeYi0vcme4B
IWzrKjP2I6bGhtb6XG1mnng1AA2/7gBfOa0qmu72iJRmiJubmqpTurt4a0eO3MqkS7SlLb3OUrtk
MbbWji6jbAzZSCGYYZn3A56EcthiTrUQqvzKj5FCojDc9See2FjSyVmrcFCErfzWccyfH610Achj
6fGPsuLx0VouX4y5AIalnaAcq856Y5yt2P6QVVwW0JDo6X7o6rD1DiThIg1L2rMlpoSgfPW9BCf3
4OQb0BSye07fOPWMU7whkikX17T3RM8ritZ4dPvkTP5EWQX5CxD4QAiAJ0z8cslq9+a1XWS6zDXM
ypBx3gNJg/cApotpuddZFSafd7kOgcm4i2//yHTNAIPIVqS55Th+YDKxwv5XWY4v1Or4cvUQU5Kk
pgbq4UldNEpEUG75+vIh+9L4frvs5fZd7hEkPIQXKo19jd99Z7Unxycm2elXdd2VHIBFZLscnfih
8wKT3llET6xG8CSMmPnEYyZyO499fpvQVdgtC8j2KknehMz7YmuyowoSzBmmLibyMK7CJb5wCVP+
duynju8Y+VGkxW1OpS4Wol59DojtVSAAR7rlmVfJc9zrHUQOpMMaelNFkZ76jpZLByo1aWVPhnBX
DJqLyWeuejrwp7sHWgpXeaTPI3xqvMrNUn6w4o/y0E7mwTMDUkd8LHN5osUSVw71QvAlNnxyPbeh
XFWv63B3DhLMeWUX4sA9hwCLwaHS8Pqcy0LO+nOhsH3HHTYNVl5Q1yos7GTz7rzR6JVJMEolKA8Z
pFtXU5KNk4elwqmaDHQg/UkF44Frev+BOCAsQBBbnjDOy9ZP4LLC8zoE6YboJf472Erejs0Bb5wo
cQBm35MlN2t3x+uJH3Q6QsbGJ2IZ3v1ewKwsjdVKhHvEkofyS8+Bx6FgnvS5tft4qD4JgKbxXaIv
sH71uhIwNlwfjhvsmfO+q8W2PFI3dfcv5ljTtBE/QcDfnWJFSmz5uc0Ae/s9yRKakaRdejx7VLMG
vEbks34QY6P+rFBft7pSwyp+LQ4qzgnuC/m2+zXV9iyQxz1b/r4V+7jxLOe+IGGQfRupWtffAqHw
lkd2QentEEgCbzlhr4OJSkhMSH8X6Who+H1Etif2gDkHRdTlxUzhToRCN1CDpqNlD0U7vbPWlTms
z+q1SycVb5lhAhYOKsPjKXcrYtbfA3IOFs0P2gtxl7JakJztg408INaomB9JN2rvPFZwr6gpSal1
KOyDVZHRTMdtMftQn2rJLMMGTumdgV0IjFWT5lOOkHTGee+q5UFlbkSNvxHmRt419v6rjwnjH3Ck
GHYFhVZcv6Ci4RP9Gr+FMnhuXsT7wVZjSt7wCYooW/ROK4N00aqECGkdcn7+2tBCZQxBFSfx2DAm
tu4dVDKMjJq0eXhGFLK40BVbhdd2ZUAkQ9XNyxBikHQsKpcjY4P2NOxGNLzrHEyM3GRM416qvGwX
7hRquvQqMmNrODA1hHrjCe9wRhRsu9S6RjVVVYCNXIG+HfIQOfVmDyxa2gjn6CaX6WUbF/hAyt0Z
C/2nn2dNwoTnyZDgOVKaVx+FAhxLjQPztMCzOilqD0PBxjoqhSc1DMxXCJJjhmflbK1ByoZJb1fB
MTQQPfss+qN0lasNzmircCXOcXduJo2qQrWS/ZgBXccVJpYWx3qAfNa17Sgwpv2WtoV9q3DE/65p
OBme8xzka7U3cHPu/lNChcdA1geiv8QwlL9SgdnWotdT4L+siQfwISy1sKPkYZCj6+7dlibwffmA
OljSxB7bXgKQCJYPraOB+Y/yriwEcvQ30zlSjxbNtBS3MX3Yr3iFBA+27WdAqISkSXM/JH8nZ8kj
RZ836Fcar/zEzTSQivNRTtx57ZHZoSNZrsvv00xJ/2s02OwvKiS33+izwC7B5POeIomLJ3M2z4MS
3qtTBbd3ozsymfUyRC+tXtswgwW1a5QLxoa7tCNJ33TPLevFOXrbkbNjZoNNeAhuzlcZ6Me0VoYC
LHuj0K3aFEQNnlW17UQDTTOJ/OnUBtXzOtOANbZqe3MaxOsImp/iDkhoGJy7ffsOQvhpxjUapM7+
VZItzWcuOi/NVR8fc4GPvM2ziGeLbj7kTEA3gLrXib8qlPOX0JiRqfWCii0U89vxMMoMaBlO8s0j
k8qA+4zlL/AWoMTPhhdtnN3lIhSXLPa2GFdtIYq75oWTPllWa+mYhyEVZcHqA0O7JvUxVTB4/Q+l
9UJhmufByxN0teUGUSNNfxuix+84XxJ9NqJCnkGOkHkReLbuvW2v9nsH61zPg5uLmHDiXVfUMmRX
cVpiPgMGMn1Aeczg9liGMmXng9oH/LIFed6QB3kxGV7qV0HdSxPU2PJi1VG8Egh6/Qq96WDuiQCz
nl0Okp0FSKCc9/pfdFUp+NdSet972SJ3yBbZ02STXivFBeEKGPpDC5000bZYvT0cDaAUEMKCdXI/
kgPygUBgDiHjQFfWx+JrtGUw2yTplmX5dkVUgAUnQQjEOkjnREoeZt1mZ7WBbyqMYlOn6k8NKz1M
t8xVLzZjgy+Y5NsPFx+4/jTRLGHM2yp0K7bvT647nR7qqs9TYTEhrUKlTyVnNraIhNzGvoZ66zi5
SeEBi/GesMt1qwBFE835DBH3bGtCgwgrweDm6+2xXQXqpVnRjNMa7nx/MioCp6B8+V7G0a4JdEYK
QOtVTKygwJitqbm38ai+xNpKXJ/NpyglSbCBQb33c72cYmqF6iwDfn0ka0WLBNUzq0AjeLN0SeUw
srMeXC2RSV0zX9udKLWMVI+Shx0audXyr/4QvMYkiDja6eCS24m0/HzTePWujcdaMogWI45K2YYD
xeQIgmHAgvcZt70+DpczVM2rnfPhWfEnbk9vPAUnzTLqOJVp/EwbNCw2AZkH2n7yxA+fVgpBaIeM
z+ZOJcHzL24eYcaqot9GxK7OizVeYN8bSLgWSipRPyKqbck/Qn9wt9SpRVv8mPaZ9IsLlltjwZaS
Bp8d7q4CjTK/w3KB9nS8vkpJ0TvYSPIfi6aNELHTCDTVCZR6qXgS08wDwPQjTL7/kwk3cFgS5UMQ
MPwGUi5wG9JlTBvNTrmdIeMghCBv+CZd/i8OT8MYH5oRu1gdxZtuib7YkP81DW4hwsxdODJV585F
o1IQOYmLTfkIovsCn5JgNCqAaiTDmvx5mmUKfegOrmZ201bfGh/KGEEyMqZ0hXTu4dpJE0oAibff
5/OB6/VEe8h41qaYxHV9nOoV69eVEkR3nO457+5W6yA6VHt90B7BjmqSf69r54l8f1eBOk7VPO5x
sfnIx+PvFLRJr+bmo32hrpLlpzNjZNHsUg/67tYnFgc8gcld+y2vDyLT3hMC2XBKHbAr+nOjhOSb
KBWlvHfGfpo/pEG1C9gGpoyvxob8v4u3ux+UtX4D/QIojGPtNX1e9kCIVDNM5MbtFC+YMAuyU8XS
T96Oj79WbTmo8iXpMBxHrAwULFWF4yMfgOt00tvJO8TJf/HmGM4gl/HXCqeF9m14FugESEMtW4pY
vdINCzOGBNEOW9cs5ddm9QmjZ6aK1B1NxXliBDsVP6EQyw2s8pn0DtZVYKiwySdbcOxAL8/PkiLb
VLDBWUBiZOR4hzBG+TFZMkIyl3AAZIXb5Kc78UxJ92BkmfPtRGBwuawhxlp0BTOLljImryM6b45S
HpFw2jweMjOQn9YHv1V9WQtMgJ8vfzQbOd1ziLmtTK9jec3ei6nolmdnO+0nXF7u8Mrw8dXbMrAV
kfiJrxwuLmcJsy6jnN1TkZ1SUVglpcBoOmet87+Xa8cxK6To+w01Tx3XG05CCcskPibzeqB6A5xC
Zc5QQBnQxqX1zt3tDRrRpCtl8uHGUD1aZl/ck89ABQUCMwyHLufH9MB43U8Jm8GQoNgAo6i9zq8f
SqDMR8rC2cnhspGjWK/AXuYkFGS0U9GF6UPuibdhpf8ENkcZ/oZVUuPHceEgREugpgHFraDTO2yf
riki8G6MWniXlnKpHkNzH0bvum34krzJBxbBbvi6LVbO2mWoL4Cjd3RwS7v547T4x1CvBsn+NAiA
H2nmZmeeM9lvfThXqk+rz+VSSbe05L2MU3pD5Lui5ymUKNe5UM+vl+OFdVsCymaSwYbloaASkWvb
BW4gIH66agc7g1kOVkjrSXDLyA4voAo8pO0AfT2GuYE/82wLYVrmy3nJ1ZNkNcT/n7EA5MlMexre
mEk1JsC9kWL/guZNymEl/rjoDNgYtpUke0nliGTOQcLrNl06gb+pVZhbe8Bc3xr01skJt0IWMO7D
1I5Fu+3sDi20+oztm+XqDJ2peepOSgFwrt8rQcWBytAFAA8rVmRKXF0SXDKG0pi3CoqTIrRjuhrt
bZrgk2rbNdFIwNr2mKWEi1XcN1dv2wQ27vsQeo8Oe+YqR6+Pk/Y8PUp0RzOc93wbqo3dQr4HNLQb
NtrMq5SWgP8hcUlZ1+e6Ivugb2G9YAlEmfVgy/IqxDNuKJOuwJVlVZ79/tWV8lYE5Rw6XamFF7j0
csMbHByJbrRFMPhCBfp3Rbxnsms8E61pDFouAkoQjXN4im1lwsZOIitreNqmy5FQrYGIQ7g3BFcw
wmUrcpXo35sUA/N1zZFWhIen7PLMmULHfhur8vwT2wr3/U3yg6L37YJx9s3qn0dzDIP9jCfXJpoo
qKl14jmPwaevUkj/FEwOq52avv4MvTa98gn65qKh9McAK+4k4e1yItkyKvbcTVeSdi2JgI0fh/CZ
dolr1KQHd4iotTBxEQ+mH/s6CAY9nyegVKYRHt0/lOP1fsNmWFVIurd4Aluwrmvahe78FuiPnywb
oHGsL+1jKs90S5j+HeJpmpU0Gx4DyzJIC6LViuUgIbdPde9Hr2sFyyBfInRnQ36Z/kG4xYnn5yXl
Q+AkOa/Uo20mFN2cRvt68lVqQSzibml8SkEG9oZSzo1khMaB3yERrkR0wRn9BCs8eVVHD9EszfjB
v6Z7UrXdZ4hkaoA/Eod2khC4l6SWLQLqORI4G9oSlLi/JsBmf/sh2R6k6zf7xjNSBmpejOSB6MJ2
XUKRZpL9Gpt2T6PsBrK7lOUPuYIpDUzyGdDxG5uh3g+sXcCZ2Sh5yG3Bffw4HZVYF8n/YCffcIkA
4njR4XzwPgZCkG8O0F7wHtv24fpK6QWVpgwci2EK9U/OF/1VVSoKOQ0da2gnfwbGHqZAlRoXmKIi
EgVn4le+Zv4jhm9+eYsGr412J3X0ipQe+/He3/+QK+bLuD0aOdDaQrr1rtTHfO/a9BXVt4VZSvBz
0ljYSqqICiZPBUV6FX9QREGRYz+prO0I/dQ91xUSLhTSkIgj5AKfvc5T8Oc+LrfbXXM/or3Aqjra
0xPKXnRyBszcBYqYxUHbgwDDOBYDspIb9W/Qd69a0oizoIIrbnO9PxBOw78RXyj07kh2EZPeLK2p
r0Kto5Pcw+E3MWodnx23henkDimKf34BjOFPUxkav8ArGSdc/U1OESTzY0VXLOfeXvKiVIEj1Z9s
rSEtfMwRE6TDwKgZX9A02c4W/XG32DsmaMc7VJKNh0Z6N/d1st2WgN88IQdU54bQCMmESYYNPGP6
6/QGRdZSiVJCkCwgYPQi6MjcJVB0gWCmU5xy6Yj7xEyTdgoOoDIHswlxVDcSyPl5viXKHXARYzGq
f604A5/e8BCYIOYCuyP2HxxiQ65/7BhViz4exLgSk7DhIO71OQqno2249NOT4tbWscDHcWxdMbVI
yI7YYDPaaTpUhWvayMBpan0HsoaVZdd6XWVN4yRnD8tpP10oTtj/bHJftfwMEw85l5mkcqdybeGa
oVK1cV+fHoheQlsB0X84UgfHRPc+rygC2wRD2ZgOJ4/bGAhDcYq0X6lpZtKWPfP5b1NiV9rwKOpU
VJfD7jynj4KV7EX51hxpolrCw0zFbgLPjQ471dMRKUQcehoIMz0n9l+DRwLx1aJUvfEAA4d9hpcO
uBngdTebsH17aM3jzPh/fIAvpCbFswqVPmN8Ybwo5NCzS0hvlZuddlcuE/UOmu0y+Tj4vj/wYBSb
QO8uETw65Nfi6gxTG9mfIcJCaxD9iCrSA7modozdDWxcDxgS94CMxAuauEkEORUcekwAualZrPwD
YnAHhF8VvZJj6lwnctoi7M7BlmbaQN8fQhskkpgZKJlqKKpoVB7AIs/6TnutbIVdCQvSkbuQ9tRU
ErE+RwMeCj51GjtIFLZhfwy+VA1ixyRS63lM6OvFf4/W3jbuBY78C9GFExKrpa9xAR1DdmAGd/Yw
ktVZY03FP6IT8C06HqefBJ9lgOirT3zeszdPZpF4jlNceqfRa3pOSn4joeEg4MHi00Ejd4NENwkD
3Nwp7C8K6nA2Po1gwopD8RI6q7Yg/Qeag23nO9evKstr1WicJ0E2XJmIInr6ru3qigTBrED5+dRE
iPYxHM1byNMK/XH1GTIThNU6m5VGYWwRKv4TqGcvI8NsVWz2dmNW4CTUiuqEL3+/cuC4BDmti6Ho
f+d1vjieXr4uTJd8R1yMWoV0/MGlJ3FOvqfIbUk1jtGK/0v9ftHHkb/xi+VKsM2APBH8IGjnU3IM
iLE8h3tdMJQIiroLAhl2j/paljooJAeAyOp4UwktPyptW/m0mSUI18PzC89D3BCJq/NgkkQziobs
vY7px0RGpTYOy/suwj4RqdvaphLCpFpEebqrimLNLmJrHC99aSjsnUKPJykrSmdvnZmBG1QfQY2O
6m1eEbitzdjZvmgzXYApup94yU5AEXG16jqqgdHkJ1R/CfvO+QAfD1BlNq2Odytp1LT8gouhtO/Z
tBgv2i0c9laga6AWdQD0pwcdgbGjFYBbYDHsXyXZ+lA8Z7Yw4IYiDukLkKLKWrS/JK41tfeK2PJ0
wjJPnBxxTY9FF0INJdsv8+mVV2O0lO+xcuxfixJFIPoOEyJVJ9fRhrBWuN9Sgqv92DseeCfufHgy
TC+M/J4H1vIPwsLNaO5rjqHJc4IfmRvURKtAHJ0hsBuW9AOPc5F798jMdcxL9/QXkGqro+EzBPtt
/aG2zTdzMDQtMVyLhfNq9z+rAHEKU37XCrHgEtD26vV1KgsHsbFd4Jxyt1oCN2iKWGK8sCfdbDtg
KklOgnF+P3ll7jlmISNh1QWHm2XlU7XHS6+f+hTIdzOM6WF9McdjJu/EQg5OKaVYLrrsUxauY+o+
JadMmO2gZeDqXg9CH5KwjA2y1FQfoQnQzuToKjCINRT4yxG+Pj3eNwrKxxTJWwBFbvosAbmqnFC1
knYhkbK6L4Han9AWWcBr6aoW0L63DELm2qfK0spgmuuTBxuMv0RXtp27RRfgxqH4gmMsn6GEC/qx
lEfwJrkOdk/PETdkiwwad7+ByS/gVP5u0I0kn+SvrSdJvsQDvbnWAMCfbcYoTW0aNQLxMzSnjljp
mDK/CbVwTSaKLUfqvYdNLi3kCvZfDjM2REifAUB0CHzfXEPrzP5nZc92AWmrPB09uSlP0UwFFFsG
Jf9G5qfnB2qtengpXVDN17+fmswdDVQA2dUgvz/b8xd7aSSzm3ga6D4ZgYyWwKfb8D3Lk8JskwTa
5ptloJvdTRx/Yk+v+UrrtW64ECBLVT2qVlDDp4ARdr/Wejh+JympPRJIEIDdcpk/6ACdE68fPekq
KOJncLclkFXMh5OIst+0unyyWqaLUkleZFSN+gxupIr/mNvJupYhum1laRIFX/6GUQqfNcO+iOq2
4V0WJoGdMfMmsQ+hjBEpvdmsUuehH5JKMRwH7+ASyPr2TmqJTRFlDrm5kbnjtMohf3LMvwKCY5IT
4DkuR6VY2lQj41V51hpWmcOH1HXqFmAfT2GxYN/2jLDOSPYsv28i/IBQPdjgJYapnTdReCxTUSmo
3zMMLvd5Uqp0NWc7loHQIMSa/2obEJ4TLqKqt+OPuRsigkWyKj5SNv++Wo8WtIMlN4WYJgA9wbDe
GST3SSWQtcSyh2WHN+JRJF6rProNJNn75NhlFBnJQmU22uveYQQ7sO4gCf39aqby0ijKGqUTn4Kz
eAqBasiolPLBrNBKsJrFmuEDbyhcR1kjH4w7lGeVHSEhEvVQaO49nAKVvsMzuBzezLfyqxqbbDDY
l4uvmiuh0/PaV/KJ25KNnLSSeCY0WzLsETpvI6/J1OHhmazS8ua7biyorEeMxNO9ZFOj4axwlHu/
F63RCMVLhUzetBtdV8xycRZdaVcf6fL9BDrgaSi6CokeSpHBjXfWtBcWR1iyGtvfh493/od4sFJ1
8I9iyljGbiIh0/8o5LDUCiYTnenHo2dCvVR4PNn1MTCYtjolooMiovAWgdQr/nNG+uT98kaI6OCl
LmXvkm/PrPRRz9Juuw2VhMsL2lXHzjZa9TE0J3Fu36QPdzfCg0QF01zarqane10QuOgmt4Oz3nEt
IzJD3BxwDjteCYn0Msm9KeXKItrXdkTn1Cp6TyCa/iPssKY+BEcz+8mz3pNXpqd9tNKLlRrdytDN
vVVhNAPTEEzLByhVHCekLBG7nUqIuvXhRQtl6pvQKuhACk92dRa304AHNPzyj+tOPjjqdnecmbxs
xwnlZvPwM7AxaEFw8nDgw5WVCxgILRmw4eS/K/cXTuE/Z13NxJ8fV8rfVLsrtileDfLOOlcjvMiG
p5Q+JVjr0hnjpaloLv78jekuhYAvz2Cnxt+aOftrOh5otTJPt27j8c1A2IPZfoMZwbg4P6xTzLbg
42P1aCjxujG4k1F/t/+BuuzDDPhYZwc5j/l6RGRCk9fKtLxsGGHWP+HIWC3dhHGhI9OONNJRlGav
ef5XztBzsckPFtA9jdg0EoIap1+OujcStCsPRqsL5jDPGWzXxeEjtsEu/XF1NVq6/kIsyERk8Ulw
9thfs1TAy2QTAwpFTeYrCq4CSub4KXcmEBWIEvLXKqirFbc/mxGv/HpQWNdjV6n3W/8//QBs22UQ
8Vg0A2SGZVnV2nlC2EDeukQx/lL9autoODJDA7ewe1U0le3hgV2OGSPEeCIM6VxQVsUZzXS3bjAS
GkyXoBvYj/T5zvRTQ41lhmBx5P+jD4P9qWUKcDKPiViZxrixICamBEGAgzQzzC0qSGIGtgfBuzDb
xE1SQKnFpd2jeg7BXbDlU5LuSwWV4dTudAzm2cskmj/t/RDo+8v+3Tt1Jl+MNL0+KujDCEe+bcwA
upjlbCN2Tjb46e3jTfqaAMLyHUfKCCjJMyWlJbK2xiEKa5NECOc8ODRJfQ3OztUJadAH3u3Rd3cv
yASw0YuK6iMugnddU8isXEZgvGDeIuHK81EAdJ8vULH6Fgr28vdLfEoAqx0zPzBfnP9KQteUQWfJ
Cbl80kUu7LIFWGTSN/fxRUuXf4c6jef1Todlbcm3/1EQZvutyEIb+Ub/mCvmPYtBhsCtNmcGhgrV
KmJdeTOCugSfrfYyXFsnMf5yuj+VxBHWxJL2cO7t6AS/gCSIbD2ruwYVc3UPJY+kUHXA6BXIgREo
AlL26lCm4Rm49cmiVE42C+wRvM/IgLri8sq7ECjhKhUtN2qOIl+qizlss8GqtERBwu0S0gxUmKNQ
PL539H0OdzzMOrggtgmv9DTSz7SrzPqrUOsfYRprrWVsbdt9gCpRagNHBXBOBMjaAimLPAIlrc7w
fsmX1jBrc0SCcPZv9H1+2gRm5/CN7+PvxY4+JDaaOhXoMuMHkskIc4QWiZADRJ+tl42rAm5uWWRt
R+7ubLVNvcNiILTcRaIvtgYyjIrObqbLwzAhzVEM3clm99Cl8RWWL1Wxr9mWYNj2v1pOVQS1RDly
4UFLWYcRMcKn0I5GKQ7P4zRh74jdf3bWaiIkq+puLADmbHfv76FCYSb8rYWgM8+ZF1V4AcnYvinX
EYC+O270TRJWB3oTQYfx2ubIAVWQ6oX0DhvBjj6MOdrYcmqh4Fd1fYe3uPvAv30DqOqzVHyNKtOz
iAHOkC8Kt65rYKOnf89iCwrtdMdzVC7b+OkQSs8DVsRVEboTJc3jJiTYMRxLuMUvgjyKmqDjNLLS
JLDIT6TJZiOfFKw+EoOuuqb0ue3tGmY3Xb7jDgL4bB8Cfv1sRr3fD/PPLHucz36gRk28CtHpXE8R
r+fNK3+gZybcnpqZtNrSaTfCk3fp8PNLBZNn5t4wxDQkcSy5/2E6GJMgW3K7oOTcHYJ03qtyEcdg
CUICI4FXPirlIoZzYBbgHy54eXU+bg1jWYG8bMNmhvclIgzsFno9xEf0uEihACRoe0RnUlKtrunC
d8Ka0bATMDvp37vfzzvjzTymvwrs8hHN7PZL6Lrgyy/IKYt7/nXxlHzSWPkXjyUa007zygJWLhH5
03C+VwFRuwcs80Ibd7cbaAeaaxnH2sneV5FrbQQTi0cW7kng9oO58IvOSPeJzGICH4Ze428NWc4Y
CMKKOUZGF8mhduRN/YvJQt+WJD+qpbVXUcd7K1q022R75QojDfBavAcxEoBM0amY+04KzwF2gFsO
G7zoxp9LnodIy/troAPgvilljTiUWr1V59EbZ8hFo8D0lf22IBsnMmGMEca1wBWr5MhoPN64br1y
zyhei5JfGqrBOwn3hG5BLXW2372loOuD1pa6EXlBaakPr5iQdYME7116x19O3mQ0RJ4Yf34QxhTJ
AO7NaJKqPDCM5VolM0+i0zRwRrxTEqXgTKz8rBEFt19JnUXIxBCCNVYdLVF1nIlJJKz8l2l1Cp0v
IKpFhEsdPCOsGNzjCQlfJnRDxHzkzOd1VXFYxqzcguhf/yCJFL/l2eiahUM0fvcN5XQYa9t659nn
TZ9CWroY4Z0hTDTTjkbwDcg67vqXIF0CYarxWlHJpaBnJymoDQKJKx/9C5XqehJH66XfcJ4QX7zQ
Tvj6zM5zqd2ICK5r4m9VkFuBbvpHvFQdXp5OuMBgMi9DhH9dJkT3CnlW4wwk/kfJlL5ENArbVaqP
YV2EUJXcCXvmoHl0Pdab9cPDry6R/6nzghMbErocQ5oOb9s607xuKwjSJNSCa7UWfqETluvfRKFj
Ur2OFsGZ5xujchcCepqxx4Lf7ngCeOCZIfS5X6IyNOD6Zwec82iNizYChLm5squOm1aBjXQk+jXo
KyTgHmXTbAMjYjqDEUBk71n7ssmTD3QQO7y+GyR8nhd1B8l/RAqP/nGnQZjCDeLWbEtkuxIQBnLn
sZlYpysqEtidc6dc/VboC+Np10EmCDORlTH4ocbz8wXXpeVxoYqnd+hNc1up9r3HP+g7/Gq34KJT
UQ1QlcLFaobBy14KQckcrL+DRp8WIK5WMHY+rOi2fsvEVgXapFib8/pF3uk5EmsgP4cyhOdrhK5L
WjMA/UzYgJ3RBZOuEQJx69fQVfYNPjkcHCzzIUhqnYC4uV5+WPQwdN8qPWTLXpx3xfU8OiJafDmK
nfPrc0JRlfkQj608c7JvR5Iu+4W1A0HXUicJWaT0sUjthiPTf9t4wqUsNwyeM/dAaHAmOHCBguIi
krsW8S1HxD+TepUt4lyUwADBwghZlTR7DulC1SOemRLW8FMDYL5odKju/isBzCZOmbTHd1Ul0Cni
Gewya9r1dXFoGjpztEPTfuWKsl0PIgY+iEUAsNNLV0nbC41UT43DOWpFdpTZssywQ7TZi2TEnt3T
pD6Km6x02dgWfmvmeDQEtc1sgu2u1eX9p1RTqeTk5XP/iAgMFvHDZTZdqd96ATVJKVdjvubHwTfq
qn8ndkVJ2g6dEr8aFKpmgSXH4QhffbSkuqDZoBcBh22K7JMqq9MZPvAXX84/em4SvbmCk0cITC2v
UIM6lmLHKRkdmEbKTL7s5MVhBpuo3ft7I6yl6ol3CFbL5uGT8lZczDpX7DI7y45Eeaw7XJ1njjbl
Q8zq7gfUl183cn/8BmGDMn248lG3/NDDnoA206JDCsdGjXbhcgR+xbZMt5bHKiAJr48lH5/dDkjV
0yzs9NgtYVAzYpz5D4uewBp/LHzR2Fm8oXxXUCVat1Np50iWVMtGd2jwj/q0QU0PsJhDsjJ8/M/r
RT3JG/uao5lZZ82q0ovUcSKvdt3BxY5mIiyfFBnGpXx6sLEzB/bjdt1vyultkDvHrgBgX73EgXRk
cMZVLycE9CtsMJt5RsMOQmCpi+koc7nA3UIHdWq+zVV2eic6pE5cmCt5YWwTQ6ZggFa5cuOYf6b2
VXcnd932eVt9gPZ1YAoesgTdWyOoNbeh6i0Ta23VSJNvvwbpSzIC+BUvLW6FXhnZU0eY3ZePk1IU
n8zgOqX3UbhZA4oHDdwU3ZaQKchoFPNZPFzxYK8KzgZIQeoSafDZxDrHJN81QHD5jpzr/PKeg7wa
NCuYE5QQrQWQMFbQzwwwWTcY3UGMz2D+vmFak4Xc/82hPkjZn3QcYMmbeAR3kmGC2rT3hGFgRMnJ
LBJhYLyXtJVS78IuhC9O7aNYdaOHAxJMn2iuyIuKGMSYL9agVmQvRs7eDaucF+OW+u7/UTCwHH8c
zTGABjAB4swnrY17KygGb94HqvLmrYeC128zL+vYRpG6rO+yfB8wvf+IJN84LUGUrcRPZTEeLwoX
JFmYCrr8OIRq5AlaT+yShc0Ij4d4cu8nZH17uDbmkiJTg1fSrXn8UC3Ec385fTacMYa+9ZgaUJdU
lirLQLCP8qLaadEw68LYbQhjR91DLkxQ4GKY4Me19D3zoddSTCBkachbBvBnBLl1P5fR1l8ABrrg
tRUHik2t8eZsSwKcTZkN1yggFKXPsCpyCHCgQ+Vs4f5+d8KjrsrgFTPd6pLWpWTLGzdixk+NiE/O
Mu/5t30prCKN0MNJVTrCVPidYStLyYOYaNB53kbFAqohLMowd+5xOTqDv6bWpQmaUmxQbDZaMUv/
lf7yBUFDPo2hmWs7AgvQXmX/y3yJgZr+dIWFVxJDrFoQg6VSZRVgMWt2Lq7Keqs7kwHLeAxnYOyb
p0Ly8l8d5IhREky3jJe5dAN66806/gH60TC5S82eV12weaRuQMu0emw4oihmRD5TlkcXfu1I1CGt
j6u5+Rt0r0MJy38NM2gAOlQBYdVBZ+b39gZLDjaE+Vz6FbYiYPGd7fjnvyQ/qW5aa5XdgIrwJeMO
gPyiGHDX3dmd4yQdO2U05DNFIAc/vrEqyq3N8nefKYjoCOj2DmbcQz0+fJs0sSreIMXTg/8K4Syo
sFRgRGZ3MX+YWk85rOJ0teHcB+SHlQtUYP1VMvETkfZ8xeiFdAQXdJFUO+nAftp4E3xmPzZEayi4
VHSrpV3DS2f7XrGaxDNBEJWf9dTMbvIItksk2bK0Nj0v/ocbdEk/FANJe4rIsWSMrgL9QGPplkQv
zd9dgwaxC8AHLAnsCBtqhdSXYfX9Wc6yVekEjYbzvMiR1B2jr77JyjUyQxoEpHzIT6ht2cZEAgKy
PGZKwznE8VcYVZyI1AjMnHLEYZis3JJO8wDrZdjEkxasA4ZBxFWanjJzyztmb8vYEA+wonvJH54t
wYJ6MZPDP9eeF8SzggjcVmY6SnHX1RXLYglZwtlzeJiqTLP/ajRnYD8hEa1EAvWnmr3+5wQP/0ul
Nijfgl6h/tUUSAv6te9bOW5IwfWt83Drf04YLOmprjqKiVr62h2llnq8o/k0E5NWtxkbXZ21Ti4X
vv+9thIKBfkMiFC8eHTWFdR4MtcGW9/tZ4vdoxFX583gJI54cAeEDBPk/5qMC8BDgiB/LIIdExs+
ZMtpuomXv12fl3tpi8HxB8xBN2XIc5NqMYgB7Lq8ni62nwn0TBSgGfKDMk8x7mbOG0sPMsqu+TqV
n2v+1f2r87fB6/lC8Tz2Pa68BJWro9mTksKCBrmHzgi6NTMKXhnmCQICVYCZzT/eDiUb6OTA7CMJ
MEJJfOZMWQpKxlvnJDl03p0VfTbDcid1oIpDBK0FqHLbbZzd0ZohEStiihRNZ6LN3lmcJZsMRSbp
+kRBRueO0LbMay8nSfgnArPQxRBrEXOyhmNzRS/ebQFZ2B6aBt4a0PcVTK8dmg+888NOh/rq2IKJ
VuME+65qMoiGDn5vNEkC6aJxYV7WH2g6/DYEo7zGRJFxVnL3hmCj4uWSPM2drf9QmXsspyPR6pdS
c8C9Ixn36/DDzqHQaNyEBxkjARieouaYR4LojJRvi74qZGPm3Ixuw8WAG0tksV99zYZCRfk2fY2x
Hby5BhL1qdV/r0F7uN2s2cpZ1XQQFz1NQxZ/9jTOmomIpJKm235S8+GzXeRfLfqLmR3NA/SGybnj
P7Y8m2u2EirJYSkBfV0iYFQuhg1SKVh6JQNrjxDXWmV6XGWfF2T72LabD1M7Rz0z1MFw9DIsD01s
RVaTyP1GVLi1CwJmX1YN6FK3XAaoK6cJFVY2leVBIPyPhw5erR0uSDbhaMWHQi2bo9zKk012Icbr
NpgunC6SM95GbzGGiA5Vuucs0SFE94aWbVKStD2yO+u+z6ZfhYt4brEMG7Xugidcn3InqdjPhAdh
YQX7cjz+2OJi5d//E6UQgloc8q7VBHXVXJeJfGst2xHlKpKfZiwwr1f+eGZXoJaw7jmo3qeR7hSx
4eyLUe5NlWTCEGQ800LVHm8lp40yrrqf8yafyInqKlcYXfMnQWJTREPkQyJPpTNAufIC+Z79glyD
oexgA6kdx21PzY4OZy3Kn2xMImnvu14oNzvXPz0gULN1lL/ca82mGWlBCjviX+vDuw9wljqEjAOR
eJZhFZfaUpA8reFfcSNcoVIK4BWqPtaWOogGEM+WxgXAgSLX13P+DTg+VVYWedG0lBAMJwqr+WaO
mBVrxtobs6aXqf2qHRuQF2bXqXp4WwirRvYr4/l3EV+Me+8RE5xDPwg7eh08GF/ikWwMePzrOSNs
kt+Vd9yV569E/RUHMOjqVr99pdVfREEK8WDexei04jLFi02FhqRMXDbPMHcwDrFSIV+gCfJEhpPN
7pRRr3QMCEKNtF2CbfY/bnmvYz5yLjYhbgBv9UYJfl3TkC/JYc87LDByXnnw13bxMkAyYatTyQDx
LODmOB8hQxuRYt3kes1tFJqrKyNlz6jWX9eNTYxJE1HE+hssicjNQpR6K81OjEnTLpr8Ovtu3bP6
uglS0iJqii6x4tc83pP7gfCnGUmhdQfKuzTAVLo+a93gHBdaLOoIa+jKaXUVGNtR1dhoPTGxsmwY
IntK9zgO8QIwBw4tzk6m+vU6HVPiU/DcBpo3FSDSOT1g8QNbtVooSpZY/UPuPg1E447eeOSbhL10
DkCDKvHCptY4OXxueCZOcfObPiRYjv0sreoNqkTtmcUjj9uw3ccWXeRyODwBmw+mS4AA5tKe+PHe
paMuyE6Fj9N3PPGqeI/vqIN4/yXxTVxjdBaeWOQOUoH8uyK2N2s9wD7yryzBs4R7QYRI52ZZx03d
5Sarzab0E6gCM81xEA5UvR2RJ+4vBIMvCtqVCF3pvxcA5+J6xShyFBO23DHJW78iANbaOMOnT3ft
/Tb6PZL+raFXYm/ZfgBgYCIZL25mm3RzgArdSEVn9CLyADf11XT9eR5r4wWyCVDB17OGQmHhwBxn
ParJsFoM/+cKnEIrfLLwKMgANRP59EAnC6Npt03ULEGwihQarXSpCOpqkd7B9sbWyOwDcqOD5CXB
rxDvdf5ZWCevyGjzt5a+AWNCGpmTmMpysIUDIUAP3/br+SRnhFcnDPn1SpXsoZzVrTo7JZtZ4Z0e
Jo1xyAjSGEAvEJ7gNHKHT/OTlcHEw8TLpPyyrrvAz95Q8fWbVX2Kg+EEcdvcbAcVfa0/DPf6Maes
W89mSGbEfUyXJp38BC+WA8P7EGLLo+zl2/JI8Z3E1ydZmBViHhdYGbYbuf8xu2W5o6k0b41C2RpP
df+mXjmHVrDpIOkbDGxKVy05oCnK6htw+iB3s9ewf6NsaDEAIdVPP9l1gDL1Qxq1bJsqKypgXkuG
BGIw6lr92gFWn3nB3qh9JC4SWrDSv+rsSqsOddxKqIQZX7E5L17DELI+q1zVZ3mVGoZA4VcS57b+
P26z0ymjVsQtyp8EqyX/F2NXBcFIqAnWlHaiEwqwbLQ/srlfLOjZ7TwNV+aXyOjsZSqLYDz2U8NK
rCWATbLAbd7/8cOR/sBuDrsZlNPyfJIE5G83NVhCb4wXDIGn+YGjRMc0UNVO/tfIJKju5hXR9t04
mDQbzdhiORkQeTTVzrWxS+Idv8ZFJmw3GPqleVDwwTqYP7GEbElQGE/swuDH0fqvopmBU3fFpnX9
3afmIZ4p18MD2F7Iu5232s1JEj50OpUuoFL3DbC1nkItACcyG9jFr+du2xBg1l+Ev2IHufwXpC99
CId1+2dNMuootPZ6WZ4hA7kxFyjgnxeTemb26Miwz2v0O86P6TAb/nEzph5oMERz1qizkPKnHNoA
7VrF45MfCNTe0hYLteDWjHktgUx6SsBVDieNEx4x6tNI82vmxiAisvwDtZ8c6HouHYoKeG8LWcSZ
rk5/In7EWEUamINaXOPw4SdnjKc5eXEBKUS114X5qQLZZ3m8wd8O7PHEt0WHlYYO57eR8MQhvtNE
WwwGuauMIBwsrE5kkYfNKbbr7uhSIAAE4uPaZ/dAnTITnGKHE2fgdHsRAXlRnbSU/8B7ilUT685p
vozh1jXzlYjaEcYralPF1+2xcwdliZjbIjBKcJMObd5HZarhiA4Dax+A2+njRqXr7vCUFPifyKSM
Np2U2/2dL9syUmQYjNVvXWnjRLl2Cet1oRtAy5VJNwZW0q8a1Ztcdyv+F9JDPryopwZYXXMBIQ9t
2qDHmW01CiKDHJyw/Pe0FCN6oVr0j9C4fhti6IGSEOl94d5gxOXuGwA3H+oiJzXQOGy3VSgStqoo
7xn0GAAg9X3Y/AbX2R01+/cZhIXXph9+ugqqb1z2EHD+2hc0rKWByiO0RvJwWBBjt/di4A2zuXDj
Apesrp+8MbGfk7Qe4rhjkNK68UbFoP/TukUWqxgyf6X66tfju+uJKyzAWFmQEwO9KktKxJRLhLes
VY/7fyvnVV0hZ2OZrAPIJQL7bpH1NIu6OlxjR4mOXu3/69V0IEy0d5TXivURr7pXHrP/QOwbU6Wj
zY652KoZEguFrz8hBicKRbpj1lkI93ZqGTfmv/WMYlxbBs18/boqQoKEau8O2AxyrudD69/HyhBM
PMYlo0GPjv/JUrICSFy1K2QLPGwnjthInTvxQsZamED0YYzoCagtohnJLRyWeI9yP4qd4Qs5YWME
Z4E5r4nynhimPU6FO1AteszQpcyOdGoqM64GGt4Na0aDN7nQHD2UtV3+5lxLfSk277zmkQ1VB4ao
SRJFHrawHQ3/ZqBZmLli41cLljex78dYUuSOCmY7L5rjnm/BU/Xdmkg3PI0exb2mH8j10ZMs05o+
sYM+vX9c6HP1t2o4BypVev+hIzha06BmV1cb9H+to4VrKU9tf2VBTBrhH0wg+KoTypEhORKVpkay
5HBULr1CDmgdpMNAbv1M2vqvbAl2912KE2fEPRKkMFU3aaTDVbWJg+YrbB2+J3YsHPCuOmJ1tto1
aBcxOMwnBI3FDU7dU0AU44XLVV2oGHbXpcVjxksoGpqSF5sSdLVRenKcyv7EscL3Q9qWAdz2osbr
NC7a6DlTm7HpPUIYF4LSVLu4OcQOTrs2zOOLg6e/0bdgalYJV8UCA6LDikL17QH3D8ueWhIFxEXs
8XVjYq5V2+xcFThRx1E/7+UgWxINHp+wpEwTOFtaPmJEEP+wJhfANG8KX8T6tu0siIn2swk8QRSs
DSOlf8oDUVXCr+uKLgR23I1CmxRBLEcRSj9m479VPSJsHjNOhVTuNZ63WKnUDRZwzr0dEkQs0gKa
TNpyd6zbK6np0g0ftdGs6Dx1dl3gihO2zZ60BHOfwhZfr7acxXKw0SnNIlDLZj9Xsrbl8WAElRk0
/xGOkP1WTfXPar/mhPsuWcrQlZe9rGDoGCvTiHLd3Hbj+yDJWxu4G/wRaIw6Zbq6CHBfRdyP2bQr
O3SHhuLGyt7thtg2q6JAjsDD1XMUhB1z5QedsWUi2qOMjcehYGEsOW3dSdjfIfp+pZTLv+h/c4eq
SOqibI7YI2U6g5cqHcCMktjA0WYk1eMVJXYd7TpmYlEMgqmGOQZE6pMo06E3tGLeKscwF/b7tHHr
nIsuNoBlRCAims3xbv/snKv68wNujMfxQkbFy1pGcLtptI0GLcwi5sMiHpyRGz8P4Gf/jDbqtSv2
KMBC/jFbGI73hGnJDQDTbdLumpqwArjJUyXyw1zOXlFjBjIkKOU6LjinyqANGoUQFRoDs2k2GhaB
fLrokPaWLk2lWV23bpVCDGMqsMBWKzeKhCkf+tfsTH0RfRuNYZInJJ09gJ9DUIkSZAkoJ9glWJkZ
gvq4tpJotwrrqeZIa+nZFrMGudwuZDMlsQFXCnZjJHJ+kUvJrIKZH/zuBXKisD/bI8kOOQOF1fCn
jbql+9io9529QzjTv0o/FIBqqSESaKoDIxGhYTQ4eia7PVfBicyI7FSrDZg3DOEpKOmKgheonbhO
K8YbsBuHKkVTTcvSqZtbaY7ljfVz2BklkTXB/WOWzlM2uB2RNyykATg/d5FbOQ9qNaaCbZxGftWW
0J9A3REMKG1wPBdSMks4NYFHptz8WOwRkS3d1KwRNJS84+2t5V9+9XyMvvtbOuqBQc3E4DD6anyz
UpXdZA6fbgzmXly0zcVCCT9p32/mWZ0rS/mTP93xo96yaRv24uDMIubOiMrvv1KRkDMV3/81RdU4
hG3xzNGB1MX8i22yiTaYttgWg3Z/XZpgOfEZoEmAWI7Zb5k3JII/svR6nF5YN6EWvzyV/LtvwpdU
25beK20zarlg7yqVm9CF0XA7VwV/GLNnmXKWaQ6MKYTyTS92F5mGsvMXgUW9ba+VG4XdHb2elYrR
fcjEI/vZbOApSXUR+gV69FqnmGTVkeeBkbNRrynpkc3w9qBrqE/Q6tQCc2F6MT0DprF2CPlUDEb7
4y2PPJYiCSHd3tRS1SQQo+QV6zUxyX4MZr/uk8mZq0xhNeozlI3hzpw4FG6fWdGCrcFaFMChKpjZ
YKf8brefW9Py+KyrUp0BlBFxoG/HnrRPxGz5yNrjF71Zuxrcukt4ilUepB0nqiX4KbCUxtdJT1XL
t1mrbFTBG8oDdbMKQruzQ1LgEjTovmznnfxT+sgF3NxTMo5piFSecq6mMp1gH4XWT9kOJm/Oodx+
gnjiZSYjffW30t/k+Q6xkdjerMnEg9PnRg7/UXqANk5KGBD2q2J0poerfRF7Rcw/podb4DXcxcnx
jJAzmd2ms+5P0LOR7m7OVRdvW3bhm8zl1jsJRUyzKeacAHNzRtwxKgfGo1145V8xoRKz/SPpK6Fb
nzdctMXL2tr/g45VkHhmgl3Y2jKUfZLx9X/1cPSLAkmft261MUCU9E9fzbK9EjZ+Iv97+B78RcHT
wa2N+iU8keKLXJoKBGrafhIAwhzomwfyOaU0elGJw2oxxoj72dgRoguj6fY2uabPD2mSQqccTPEI
TJg7jlUIRQ27K4GHOtsRnftRw2PjcP28FQp20yOtLB19dO8B5DmziQz2Q3CBX7VSlrYpDAL5XZBe
O039dyXranzEm6spne7ebhsdfyIS8Nt7HX69RHHE0l//EQM+UK6/7BEdfDqs3u1XffKYnc+3b1PU
cwoEYEgMFIzWr0N8DrAUMwaq1EpuDIWU4+teQW4r5uJ93SSWn+shIyN6fZYU9nsrCAJsIg5N/1GE
6ls9adpy1OVm3CG4ovoVWq2onWn0p00kTF3vsH1CFf9f59g0aJMW/DyyaZHjGf3e24VzR4Fwou4l
nV5Jv5dwAk5oA2dOhiyZXaX9V+AqlvIX4FnGef/39SxFSC7PqM/b1PHV5p0nD9EfN0fxN+szvbx3
GvtqHVTAEK1xxf3ArhaNDeC/2r4g8NNzQ+QdVznUILQOySrM9mgvlGjKWDL5Vd7/lvt5eo0wDe+m
ZFnu+gaekR18ttwWAS+86eeHCPkIxt8hA4jamvEwMa5nFuXaswmChWYvZK2BH5WAYtQPNGkYIuPo
9J8hzVtcDyGRQgJckO+ko+mhzA738fxZfZ2xcWS35LJl4ZXSGrjyvWkhTv/11ht20X2YBF0eadEj
iE9PypWj3OfymaHEEy3sMKXXnx+9/PZHqMFPXvsLyNJgPXdOtyXqqUiSbDlvNsLnPVk143XBPCg5
5nf8eMIOM3VBoDOfFqaoW7uSu6W6SOhceR37POJIF7xhC/9ODFVw7oUjwyGwy5aTBVETv94WJcdi
7Fi/8rTnCuD6yWyoCcCaiwzlI94PlyiavNCdBm6o9FGg4ezZsB7Z+XdqfpbhDhvNsXgzC9Fu+iJA
aXw+vgklL/gxZeFL4XOemDgmGd/Ah39jzVC/8wShksTrlp6RLhmyh+6L5XSLogGLStFiF0IeyVgy
YJA9XZS+lnWOk8ZHNbcD52NYZ3jfuL4TcOZ+lvJj9qXNlCWAopbrDMsgDL+xni3qoToAkJCB9r2J
PRwxwLuxsAHApFW8uiaitaJHlACvduUDLhYAyl4eN3UZkSDVTKX7re1tgxpcqbKtuzrm559+3qRo
nEhWss8Zbc/9AvX4dhNMGR+9lv2gGkjNsT5K3nYDEYEzjxue6gSnkFkWE1YPbRly3HNvNgQBqSwW
QPGOJUNORLuxK3D17K9I/+qCRMjsQbPDWYK/QGUFRsgYQ7/DEEm3O/Qhiter+3pNN+2TKVMOI3xz
X1uxRmj02yK/uLljJyPcU+EorkDG+YEB7Y7xXkoKSR6Kt77A4wJrBoSy+M7afkOi6pXg3R53V8n0
R1PAJQIlU8m+YWWZBJ6x/H+HiQzSlneKpWjTvEAEFF9LwkNZhZQRKowcI+mZa3hidrWDdmbOkqwd
29lquh0m+15WW2H/tB4tQEjP2FtaPYsRRC/g125Pevwg7+UBkeHASDPn6iTvxKQLPl7zHUAeOKfU
aDDwlhct87EJzKRY+S6oBPCsdwHpJ/ceM3uDBaUJAZ9vLmnDvhTMWE6n6tfsY5+rXjaOj6v+WWTI
wLR1BUoj1KDdcS300Jwwwmx0/JaNg3gbRK0nwmbCoPSv82j6DzKFOy2T1YV2g3Y3Yw/R9YoeZX5v
G8OSlZBrfe+AokFnTXlNbewiK/CjnFOKG55zVKIoUXLyzUF3sBNf4Ad4AfQD4qkF4BcolomtyGaK
xnLuBxVshF+kVmS8i3SqluJYR1Ay6FTBawNn9ThYWoy9549Sy9FXPz1MZcDRVuDnpvqTp5xJBySr
ouaVcTVKdvE2GtmxdDvNVcSwECk5e8jRuXnPxYIgiXrVMTa3VJGTOapcACrx3aTJnDlAAjCaIndq
kk/QT9KCmJInHtgRI54EYLpeJGPsm9hFz09snuNOoiHRPMiSJtFa9g4yYkeCAKVVfKlOO8Pb24MY
o9RukLCWRL0KDFe7a5VP+G4mI0flK8j1+ZPJ5pY+0vqD8CRMw90dMPuTc8+51cyx1gW66cD7856l
RokmAuEMNcawRSzEKK7fko3mFD4kxgc6T2ERzwakQw+/VVoD0lukKUSx3qnb4lRbNyAV7zARzScJ
6Zi/Ws8tcGSDwOpB9y0BiFN/z3nLAWpjIHHS25Iag80LAZejX9wMZ3F9yeocJRXn1nE0uit7ACBB
yFCglEZ5F0YZ7suC/saUOL1gedNdNesB2EvNfdUHbQoA1xXvQWRs9HNToloVvYjUw61dtf6KFFaJ
ctS4i8NMcs02+N53PLp1yh4fPhzph5NX/lAw0t+pKsYvHF9xCKmkvcq/yhFg8PyxlDI3Zy4F2KLj
fvOta9SGfawCh//ApU53Z+1a2/Gz8yJmAihdY2IayN6ypxliAt1m2PAw7STEhOZb0YsYO0Xyim7k
ajoDokYtaVwHyEhEuBq2soLo5wikisSngV21euDoG6e5+Y4F0bIoBU2kSwnDmQ1VUEJPHhA6n+nz
5fVxHva/SzJB5xeFukxUtKRVsavp8Cc1JiftmUAz+fNlPUOMpxKnnFMz6kh6QgvGNwAtPMNAh1Yv
zW1LP7toiqzxJx53ew59IZs1Emp3kgA+5XCI3jYQw47osoHPDkBSPlPsKQzGTuPdudd3Iaz74pV/
yBWvTWxHErl4ysK9fKgEmXLkeuLPqgzyAVllQeeATboiEyoVxSZzXLs+u2qvRhSjnPybD8uB9R+0
Y8JvAJC8naOb0gRLySKWiKn88iRXNwM5aVcjAmgnofaqjE1iiqfUppObw05Y09ts0ETIjThcqUIA
5xcdvMRWSYXSz9bIaPbgw85ts8TGkz+uK8aUOAAJ5mmCzD1rvk8kG7fODnaY0o/d69a13RiTXmdd
cX1PPfoOw/IcTH9ZtmYlkEjOua0EUuf1HtOUUMgV0KEuxLX32UiF5x1E7Cz9ScGEuKaxFSS4lAip
jQMmSfGq2B4p587oBBeA3bPM/5LOtrVTT+eZy3OZ11pByEknTJxLygmTCbKefCtsM72dFiMy6bjK
7795R2EJ72crNUw6Teu34lacA+Y3ej3zSjPeSGOAmTLZj0odNPI39Fs+a45z2rznvSNneZf0gFko
jqikl533jS/6LXRAuyPmMrAEMmsbZ7xkcWLvC3Yy1sTETQBMgLLK/2wBw059Vo83K2gLtqrWRhPu
l2E/V8gIyDAaYtprpoI9Es8xb9AKlkZNCxI1AxKSe3+fOhGUNTCQTwptEBi90d6D0u6Ee+zs4Zzb
9xfBG48annpg5AuCeBH2hjDkG1+XjVxmqP5A9ZYvhmWc5ZtyH1w5dwb3AFwsL1R4Pco9BppgICbo
sR54hA/gxX6bl9OESZb/AK8HNAzWAAMPGJtixjf33jFksa5cwIX/oZgif1uA+heiCJOjXJU6jg3Y
c7QVhkqTgdburb1K+eH6KLNOLPdpQDa/rAaTKHPtI/mmppoz0jWKAwPLLY+RKA0Xn9CszJn9ojCg
Gv7iiElR+z4vbnWji845NhUfjJKapAmf13bflc0A0AiyAsIT7ZwZDwKFovJ/xDJJE0+Wbp4R3U7D
unMG/q0O0ZZEhq/srN+hR+pFWgUMXXzjr/JWvmdpx0FJd6nZmN2NE9gldwG8oNxk0K9UJSLdSBBC
8+3Q9JRtzMpyclxDPdOjo3n8Nuukf+4GGMMqHvPvMaFTFUk+WKYovjUkqzX49irNCogbrBtzZiZ0
xFjyWebxuNMELcjGLWfAN9ZOg13gJOJyK3BRpnKa4ihdJmDonvQojWfbC/BpPsFxIh6Mmesg1Lhc
SUMK+ZcdILhtGYn/uZu9PsSy88HoqYtKI+Ns+emwWUuhacxkb2I+FBurb58fGLwOGMG4D5K4P0Kp
g81Zu5gPg7VFN2NUI/iv5YtmzbMlzmFt9QEOeIs5bA/CpNrqEQXaA4pJR6wH8byNt4gIztk0qkPN
0/hqHQ8WMHO65kNUaBZXOZYJvNhrHokD9uJgUXJZDPtRghKq9vC8Xkr1AFOozuBkcfouCb76CfYp
O4bQhYmxmIxgdm2N7XFvvpz97jPEZmrIN4664H/poossiEVuJ9ZO2UspgvAhHLC8pBjtpWL2Xnze
PNue2pRCFJJKxQt50tvmTMYbrS8zUKuV5eJ/nPNVbQBHyadPYnm0kwHR/hebz6UF6G02iiFZHzYK
gbNf9G1gm/f0UP0F0dZWUpJrP1XBEi7nw7Mq9J9Gv6eY0GkLFvCi6EHtWGzXQyw7tlPKoWoYQu4m
mdoDtMVf4QKKiQt7clBgjOpauDO1Zu85/8WVTbjdmTimRomQNMAYchjiMSGGhKnepelbxAAT6hxo
+5e6u+9MrJFVTo33X7doBUCAd5U6XAACvDgxgracrecv/8RvW+O3BAEqC9hD6FvgkFbetOtN4sdm
Jo1O7ZIK54lbEx788YWplMiQ2FOcEkbChXNItcX4Kjbw2uN/GE03z+nJvvJ1wwzrLxmOCTIJAmOT
9Xh+FGFRIghv+PcAb3TOYUKt6u7r9MXfbJraG85mjdw+ceyV04lP1pa4yp4pQBoctgTPb8z7KcJF
xuLhDyNd8e7RM9aTliVEsbdYfEqt+0JqNthDusPBcxuRM3p/jx+m9imU2nWC5dMrhsbG/CzQinQE
0Pxf1MO+MX5VhN1+6c43cKGB0mvRfM6tFJEAnE1oQmSlZbfkVltpysa+o3bPpKhQTl9YfxWMkEjc
MxkeaWpAVT8ony7rU2XyZ5PbIRVdNx8ISOCdpOuY3Bvqos5W6k/r262R43O0oGWJH6DpQr4HxdVC
SlAgACgcN7t9EkXtJolklYOPWecMs5d5SastnDD5SIJlGGeMr1MddYhamEyEn4erbREr30e0jGOO
C8vB8Ykje3VzBsdKAULoo7Gqlt3NVv0jfCyaOokftVv+3KA2E1TEqEI+DUJZXXLh2qbxicSQy3FP
D6JWDAkuYo3W11rWbIRCf3d4BQF9fqvm3wfbSje+qmW6CbeoKcUtR9LEMxx7dnT+OTIkL5r9F/Xb
QAj7A3Yz5sdErbgL3HrC9IuNMHKqkD55w3MBzqqC1M9aB/Qn6RhK4uz8PRo1V7vh7Oxd5V4q6gNz
LEmSHo1o5tCWU/fdUdoq7gdpuLk9r7fZf9YeLxOQ3OmXT1q4bu3A0L8OSGAvW5e/ZoMc1xQ1K6iZ
wILaEY8BPWvzQhcU3Kez/ESZ71cTPyD2NdZjTlw/11AEjaGfqweWEr31vzh9bUokqMiYiP+5Cr1Y
2E6KpIIAIYCrMn/IQIUXJ/hi9pNR6YrbP1Uv5qC21A/b3SpsC1UwXzG0zlMNYOsGkivUOkxa72FK
glA8n/lWVz4AioMRiIetIC5nvwok3Ch2zmVPUu/PAH8tyDV03j/pW3QwTeBv05MR5xzEWyMx7qoV
f5zccFXYMLc4wVIL5hrZxUuqeiAMSZLNq1XUd99MB/6aQcEliv9Y/FAl6Q1GfhxQ0XlKe3uqZCxi
WGxPiinefL7xlrEKGH/wYnkpeCdfHYc40+xjo4ONHkDbfsfltvZ7yxgal/mUaRdqxw6cK+ttaYtQ
ITVMs/TsUoxz2GAIcsnxszjtTTWq00H0BPS0wr5TAf8n4aqUC6zeA6B/bpEhskr0uYuXmf6pShwM
Lp6OSHtJ/TYPQNjtmP06eaPtLWV3g+MOCrFalN5ixO8Cjq3+GYrpWwgofu5vpcRVLdP/HsxdOMLt
wh983GvErlyCTbqv4ulg1GbKcAd7efOVnx5nstalxQ6sd3T3fd5zRRztaYSEP52Vkj48ay7venXL
hmQEXg0y/N3NlhLHy59dwCb3r5i/uWGxmFAwK1hzgkX5Zen5pa+0hTu43EWMdbSP2vzir2M3tqKi
W6889HS/dEqJUItdDe6EGpvGUA3K8zBu375Tv3YM36LSEk0ZekbDLPwEY7zDS1m2ycCcs5+9Ds+f
F8Zu4s5aYaj+P7fjTKioq59aEc+L2/TGrekInfpRp3UrRLE4ZXS/exQsMyhx1mCfAFW3gbNXwM9j
9N/H36ir8ljnq0IGgKxvmMcW/naoax9XPMjKPTsi74maDO+FzWRbUeiYfR2AhNGM698Io5XcbwWy
zIVX72h700NqRIO1N5TL4KyisGx76f3bDIW6pG8WB781uOu5eg3PP2M425YapdDsJg+dICb4kIjr
d7WNojE9Ylal7CoSQp8/+9VLTud6Oe52R/BXZsTaugu/693YVi3biTwrELLhxHO2PCjY/ujZteVr
65ifBT2++bzbDppqKwUeQUbwmqqHlwmkeenmZvgltjph/JTHD0OYeh3Njfia5ajCHju0YC8VrGJy
JMQDawsLa3nPoAB7iDwY+/ZZ2otI6EaM43HleL+Lrg+X+u46MA4OQNM3Vy/8D22MX8wAyTqWSfaW
0QBUyWfONrgyL+4BxyJjfHyCnsrPW6wOZ3mCcLZ1ghyGRRNvd45W8fSVXkwBz0Tmt7sdBuVVg9td
3LS00GG4RcAimuGa4CHxovkckZTv2wMdMTzd+Y558MaWgrln5/LGivbG4VqPXIMm4t+40ARJtY1G
Q0M2/oztP7dIS7fT/qTCRwV+oC0QQJFUaYTxatS7DIajPobDr89WACwZAWYqSxHWT229O3++FQlv
FSy7DUfhSs/pwOpIGv1x3U6fPbbyUsbanYffDZpvaR7VxHolmB0Tmt2plD1R9lcM7m6uUu9lKDwz
EmD+8/jf19Tt7QFpVN67Q8i2naPu2GapRTjoX/A/au0gfKuexnCRCWwPerVYerGoXeJHxJOtltX8
sBfjA6oEyqxnLPpK7pGoP90YcAUQ0eNQ507IxoRU5AOcgBxVlJFvuqhbTyqrpH8RfTwSZWGZMlB9
MY0hZcRRq7YF9bPx8PtDDfPJ2kNDIsjetOIGCeFmaWtCuPb0M3g9QwuayQnceQRLzTNXm7F2Ha2R
2pWTgghSDaqJIUfL4vecyeG65ko4dUJ9ME550TsvqI3pEQmk8/fhi+97wfsiCymHAGVKPKO5/LCp
ly9psbMeeYr3WeiKUnRnFS51R7gCtdYtVPSsvslNbCXfT7i5KIi6uC5jpLjt4AYSId7eS8HwQndU
cbKuKAUaEXfMQLWrecWgd1ffuuRilcZrBR86DUO9gtl2Y2IlbIqWSgs8+RHdGrnzN1Nl+L4NvH73
0Yo9BQj2QzY0+UQ1l98xajZbU2+Gs3+7xFAvBpBf72WbXdgfKMa26WmzgCEmWQKCHdM6Cj9f3fw9
qlh/awDT4h0gfM1ZSaKZ+sMIhns6MGaU0YeNcIRpcyWC1cMlqTEnNMWUV9wxYJKa4o7BcAFpRxMv
VzHkZUqcAuc4jaDYp7K695wLYyVG8QA44KWVt6NMycoJv2XATv5VtMKPpqKvV3uXWfz6XOlTj6GP
PXgM/JOYSbN1gktDKvvZNogSbnIkGKe8wvwXb3pqSpS9x3T0KPgeM5ZDJPTyGV6C2Le7XYtyQE4K
8Qw+NYV3mUjKU+26lUrYHQmQSGWf4lUvtcpp0iyuQzm1QQum5ssInjM3qOPBL906/19zlI6vaMKz
4/1/7LDJ3uIeYsRwDiLvDE4vWlFK/Rp2dLXaHoY59y5D2VgUvK9Xj3R58psyTCEmCLNkszzUjfzw
O//ynPrt1u4oS4lMD3hnfgKNM5g8gVHXqIwNAz65ysoiPLNrAfnbg4hBpNEzkqhtBQoAB6rEgRuu
cga1OyTBGsmtweqMdcse1a6eeDTOwhJvKsUFTiCQU1qo9R1i99rEmfKqfU2Z8ETnfDmM5pzHqfvy
Es2L+mOtnfcRfbpsLtXIYTekuAhoFJJXAfmDJCT1COxJXKvlREBKGVoxU7bV5XeVAt1uaGU+gNyG
R4vI2Pfz5gPAZbVaJRN6W+etFjoQjoFdUZ65hB1HnA5ll1H9fRPkdXnDDwMMYEfGzljcJRyxL6Yo
BrvxzwR3ld55vDC56ljj8Jpos9ABBRHtU36MIh4LTkUTuNTQbTzV1FcWavdm/SI6CHe2dhtSXck4
YBysqmWEM6v6i4/+roD6g8EtEbMou3MDv7VXwrsARZsLsfhf23ycBK1nLFPamzCQ5eFU8RKWiEiR
OpXO0WVttDqRKorQtk7l6CpHE1/jiCyQv7Ls1KjPotVk0+aAGoGW0wBsCvoHlrWzAaCV2W9F9AD/
7HMk/nwvK8JaWnic5RaWVKn5igWllMAifonKwvJ77BKt5fFE56+cx2WwbSRQIPjnL7jl5xSCXq1n
283+frQYw7ndDPru0+6PA6tev5GPzYf92AMN28oe9MEh6D8utce7b9I1gZ+1C0uRsk5j2te1BTjr
ag1SzbHuThneUlM5numgE37M6jPR1bioeCsINmetqg1oMuXR0g922HDhz3Riypn3lsYt8Y1W0bO/
uJQt7FT+fM/dTD4oQFrzevvGKTPQgEQTeHwzLLOMDOb+Ti6g4ruZCOAO3OQ4za4OYx4RAkWNvM5P
QV7QF1cy4aVDjteLZ16PFmathmBYLu2yS5vJJKO5sLC3mQ3acbvMy1g0J9Q6A8KspnhXONfVWAc/
VOgoq6fot8+sIUQX/TtLlgsX6MJXutpo/2iPyQGLvnqJ3Tg0K6Z4j9YkC4/7TJbIc8VmnXwP+kct
rmZBRRd7/roQKT4LA4IVtlAhRQcq97zu4sH4B7L0KZVC3hG/EK68nTtWql48HW0354fqPt4paInZ
D6dqaGpykqjRjn01jfHUVDjpFRtrFOu6ellRzVXcn2QviZwe6f5kYc6vBw/dVFbB/YV1AYKtRsy0
jSS8y9eTHgKCj2Xed66t7VnUFDn8ef/+5lQTZ44+94/0FMXQqWhAg4XjiRI3NpSpbgJPY00PnK+l
B9CjvX4v/UHjbngZIq+KUT8s7tKJZOiJ4+vhlzQobqHuYPEMrPcwaRe0r98qMUzEIrAccjlGdYRj
qlPKyHwnG6azOSIwY+86cA9+Vxui8vSkh8R5Tyej5u68rmaP4f/465RMreJtnYxD6tqCQGnv02dF
es0Glf01gk3sQJAFwb0HGFnP05VCPFCBsUcC888uJXnLESpoGd5krwPO7sF4kof1IBXLmeirJqqH
PefZsp3tZ8zpNV6E4kqrHjFYaAj0gn//70rvjnFp9c89J9q3o7dguRQMV9qZDZMsJaq9QXFdyF0z
mSCUJywZMfMnwxc9RNnBulrZe7njgQxO4l2MfR7HQ5BQoXxBRqbPgXqbJtH59N7EB5AQ8P/XNUV3
J3TORHVubQWL0ZBvh9lAiuPRI2Xj5TgLIycJW3DbfH46EqoJQfQfeojM99BaYe676MDqctYINai3
qF3KrizAGPWXZaeTWvgqTOBmWJx32i0kauAelBEx/4KC9iyzN8MX+lhT7spvmdvYNNDMN0lVnnao
Sp3MWHtq3a9cTObm3FOrC84d8qi5mecFktCLsLtK/vsAfecW3tKaNSmEW+MMyndjbv0PqhSyGPa2
yeyBvcXQcu4w+4HIzYVFoAKXCzVC+ya/dnCKUIvM6084CMKnZP63A72Xq4IIysFDl3UZ/zAa9DX1
6tpD47NScCETH1cqEst7x+TXroEkcfdba8PTb/NlZAecaxjfssqkIeu5P5eXDnk0PFaKoPt1sDDw
kc6Hqa1KYbgSoZoQ6bGnOU772XhgOD3QDQ3GwkLYFiEZhj7A1GcXkBvdBFfo15Sk8zDoRGjpmPhQ
oyGZb0vmHLYLUkAP3GQe1Y5Qmdyi1CLJwipujmONGm21J6fW8caDdJY6HAUlJtqLXay6TQlYFlLw
53saW99zo9HXw/wgIj6vHxriLYTzNgWyIc5ZH3UtSqDNggYq+bsRx8GHuKxgdsb24dei5cpS7xdI
8UaT0wQLu7jAZXYWB607xAyk2jW6osg/u+zYkKemrTwA2zbD3pkXqwsJ/uA0IarR3X3XC//iPJVy
1JJ3QJ5gRXfcKEaIbrV8uLAtQeqtKLE16iH3XohSoBl/5BksepAxnuTxgIgiyktC3tOR2HgKErC3
T8QrHQpcVXZvpDffH7IrAYXmEMI0rYMzxy0x3B9RCpeOuFCewUsqN2esiAzOXP7j5jgENEkZwMu1
KiKpM4l1j20JhOuFgy4AAoCOquW2sCNlKzhb4ONgQFT069hMchz/posezg1x0kO5bo+mSgjZYbsZ
XRNrtJUyX0evJesJgJlH+7aJCr8qLlzb91Gq4R9gbfGzb48Gobu93l8Cwz0VQrQtu6v6bpIGz3f5
4oX0a0l2EMetN67GNRqmk+s=
`pragma protect end_protected

// 
