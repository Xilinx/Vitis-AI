`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0INbis6m4LNo5fuoc/7VtaFb6U
0+5fXdMnwe75smPOBFJPEC7G1jJjzTejAYkTl7IUTkgZKL+qPo9QsJV8bWnGHQsxi3gvlQOIaFQc
GeHAIu5kCH4qdG/Rd7Opht+51SV6MCUG+Jzw6T7NCWSvcK1kUSxl+7AIlS+WIYISlJ+EKHtGVS9i
EwJnDml+BfWpTB9xPafHkbwEu3i47lW0rm65e8CJMpk2rTZCK9mOmdVwMqdaefo3r/+hw7Ca5b4h
GO5rPEDSABUFjxRHNxU0rEQwMvR2EEady4ZL55ij8w11zh7UKS7xTmM3H2SPBYxF+mGRUYQxl4BI
ie8cyxEzE/n9sY0Sw7XMuDkTZpxOXDjMDwa8Oqk96t3ukZMHsRaYWE8DMlGM+K0ocqBqxcdSU3Iv
1LkcTlWlMQgFM9iQ21MizoJYz2R2qXlwEwvZJaOkufRx4qxc9lssFq1Wg64avfwj/LMQfpWCeKfv
tQ3M3gv0lQN0YI+PwW3glvLH9RmzZ96dgeFeJcCUkjjsfv0w6eHesHPwT0GnWEwvw7+ZOF2DUG4k
CWECWb7nUkQrNZGVLALJjk57EMzNdtiB18NZ5ecbeb4K5pr3ZkNPVsVdfkQls3VMuOfM9v55h+tB
ngXSIUR/QXqznxg2OByRsQUK5kLWds+mTP3p+ILI6DgnGBMBota49LmiQjxyunLDdVoYRHoVDUvI
IB58TTjXKYI4S39JoCLJ+kiMU1pmpQsILMwzPd0Z+0qr9Ktc0qIZpx7ZCzTal7sti4YsroL2M2Q7
7W+GB0AT+BjMplGvyf2rYD4o5kZE2ZzZllhXrUPSVqXtkZ0qEeMViqlnsvIvm1bsQ001yVaAOIh+
Hk+eBfqa+75KCWfeOJqa3+d3aMJ5eNh8y5bKv00/XPetJeY0TJhs9S44wgNCP/ZGYxGtXfckX8x0
/siSgYxoVSNt3swTnVIDCU5tKuB3a3A3t1ZfYtIRxeai/PZhvpXjchqQNRCMVSEH9K1KEBNwJXE+
ZjxfWeez2DckUJ5E/B2eU3seAulkIdSyES1IydwZYaCw8RZocBjGjw0C4yLRUFr/JcAMyPwUHxss
4uZnKsTBTXT4KqDJlyixNZWnL3WrtKLCccx68yq4MUx4flWzmHcsZFtGIYC6Ek1CMvZRjpiwJlFo
MOwNxZ2FwHhqfxfF3TOsoVKeOKYEho1a8wrD9pD5eMvulPy0SerjEgdc/ThZM+WFjooEuVPp3lic
HRp9+nSOXqCQvVoL1mYwYGU1pQlRdf8S4Y4/zSpSPrR6i7aVJ7+Xsy+abKEEm9iPl54fBrcjHf0C
Mxel6DxNX4k5EjRux8fNGgvi9GYyxa7TFYzwRZC/lR0ZVmDsQw5XXFINme05gpcHWZAsR1EUZG9R
uJk8WRnEH80utiV/51WOqlxy9RD8TziieMcVrMuN9bcoaL0O5wi4JkiK4JZPdKNlqRERe9jnKzSd
b+pPLp3O1umTaLQNIBsslGNvpYTHDP/5/z6RXGVuty4VNnkryGRHASNqtr2U7AxGOVK1nAiZD9sf
pZn50CYKf58M6phOUCLP9eqk2T3l1836nC4v/Qp+ZZN4VCzP+8Fl3PYjLC2rU8rUDhXf5xyR1IWy
NcqARNtTuGQVnq98J/1wnzfYrTMjtQC6U+k+pincMa/mMbWU1dgIn3Fp6HxDLHGo2WxY9rGVU0/D
EFKhfU4RST3QsTzwAJcWo6cqbB55PUhXFCDfIkQNKWSs080lDnP2JAg3Fo79H1HGaT5AzwvYdvLx
+d9/bKN9kHHNxfsBLvbkgRZm+24Is45gtiBRcYLlWL1x5l7vDwbeg6B1+sJrcFuAs4gSb0ujYd+2
pRvfEewJ+YrlGsid63ALOg/j9L2zLtwiJBofh/ff1H/P14IulEmIzqYvU9VnQkBhgP64pU9CQ9F1
LR6Lt2ymgxUzjc4O4e+lRVSiUcyrHBOHOA7xKP+nIfme+ofUDNIkkKXH9vMODxZT2rh1NWywq8r5
rddTM1cHmHbW5RqtydaWQCkbHoo0fyVUQmuE1suGtq5TkDB2dfD/YQJ/dFdO4M8o5KtFfBv8dyVI
4JAcFRcazLGN36SK1Piai2iCZGBb0OzmBJHRdC0jQquY6joMH7iXm0Ua//EmC3hvT/0bs1G1Y21z
rhxOAHhDxzY23CJQ4j99y8Hk8c5VgaX1wZjf01SlUL/Lqi/Nr7YUjagS2qaQe027ndKU6LTHQwFs
L2xgE0KHZHD5t3giOwaKET0Z7D7YGGRUYy3m8TXbH+0UJobpjwEKoUTCKVXqaKRG0h9emr6lDiKo
5TRpW25ZXZDX/Op2cHh7ZfotWBSFaMWKjmqDxj7EKjgsZlkTiuTS57yZQLDBqdt7MHi9h4ZRVUJs
okN8DYoCvKJSokQ2fIet59BPQ98AE1eQewSA5WgN5Inhu+nPKRWEUO01ZxC6x1C/Xl/iM3RvceEh
p9MI4Bly9kbe1t2EEsBkRXG7vzIkiI9TRwWtXcvURAo6y0QJ7x8L3BvQdMe/Hv6tELe4uyyM6QpU
nbuMarfiEMFAt/gwuhLm4tHaN9lXfJOx6rYQh1qqmDoc0qHx3qsshYMMRmHrN7bGI+5/YxQK1uN4
kR+6avVXeNxLSHjTPr7HjW9Ljo7QfCoQfBmuV7E+1SxNK2B/PpQjoCM2fsc3jclUxwxhGN36eWgL
hm+cWHmvrD+9udwZyRerW+iI0nvedSB3iN7JNdJo3pJ/gQRn7gSVWXKc4Xx3EFjOc1iD3IR5yHeM
u2OfXj36zd4tabjFcrYamfHMOgwtZGV8cmssYzosE+q37p1Pl14+BIzXUrvoBQV63Ql0ZoVrQOLR
FrebuIjj8G63xZBcY22GlB5utR9DYIRaoRR6AeRFgBn8i14nyt6WE/jWwlEm+fpvPwGQ6StZ0tvU
fn4iQ4btvRMs/nL528vs5PLPHlbX6PLNcKeNAMmOnG/RkR5UTPJ+H5T6QrN591PRPOf6eim6fYt1
8nx/orjcQzlt6a8EZKr0lZrB2b0Kacqna04ch+DZfFt998WfOON9TspTpUoQSAUn3p+bVCsSK+Bf
SYzlGVGNGmJtQ6NMRNifcRLMrYsaRXPjPvXMJVhRlEYy21zl+SlC4072ZpGriIDspxvBgUrprWNJ
Z0NTCEAVmYY/4musG7Maer+3EBVZMP/ntYqy0HAuocvzmhthJjfaUiqODkegdySHadzgMLWGI/ZZ
4n6coR7xaWnC4toRPyZeHMDmGqAZdrJRO7QZk0zMYq/0fOt367+4Hsxl7R1GZMdPOzWXrL35lU2+
346StXPSZ/QVzyJ/uJrQhJrz1zotU7pKOGlWCroCyOhvASFK5uKCtDLnYcETEZcw54sHhU3WVsM0
rW2+XpiXwAuN0QBD9C1Q5ommnbXMmfsEAck0amMouk+UVEZSZMRHSgHRFLKKWCaGwk4z+ceQ9Q4/
/xeO/osY2JS8fb9rq9Ew1nwHQkWupZ+i3laADfwiz4ZXJ0UwArXBGfjV4wWNJbQSl/Hg6wnXSl/g
aT2IDHOzkR/LtzXq4czYLFqFlkG7UsNKoEaGoud5r+QXDE8cNhRn6zr20481CovMuVuqhkR0q+ZC
FCeTBa0tNPbT7B7rlcQptZrzaE37sBA1P/89ZQKhZ5yVmn+6VO5xoRQs1UbbJQPL2gH+HJvDrQ3M
FVRwbEUsvLwvDSvDN5bOVYQRDmGN0GX2aNmesI6wQkQCxzDu9evKnGWxpIckR6cVoYZT9wshFf8m
fSFO+3iMRI5G6BhbP/LEB5rZW3MeRTQc7qLxmjxLCYj3wETy0l7FbvLSO/veySem/oW2SSywlIRv
FSrD6FGVAWaPpfc3bMTOcG2DXL7L+zt112aI5/Rr3F7gW+peTq79Q1haHgIJAdyIvl7B7kowEMzd
LHXpDQCtlo10yRjRvZ4Cw6N3yThAJsk3WAImcGVGkuJh8DBelvhT/vhV1t/fFIpo91LcXo6RjIn4
M2/w6ClAV0zmnfGA2GcqpAogElieDotppzhtfkJzmr2kNXQBCWORvbPXeaLX6zMrofzfPaXF0eSH
fRRmfA/nS2kqrrQoiq2iHhJ6zXY4RQYALrnEXzY8zbO0uxtvs5sH/XzADHgFz1UYP7w0e6pgXbfz
kDi8Jr3KAxQNtRwpOgxpCdOzpqbmYKwumag5XxQ5AlKzr1TY1/lmEzi3VvK49W+2SF0Bl4a2tYus
OsdSG9NiOujV9R1g4qEIgwIP2WZGog2nVqbY1VFje8yGSJ7sjxM/JwmeynliZRsXtqW5NFCtyWGS
H6dfsLh+tEQUJ/vPef8su6PgdDHSWv8LQACrFcFza+EIVUmRbl12gzkTO+B5VbyK+ycL4HaiSq2z
qcxsBmbBRy1n1m/7Qf2cwaGwhYnUvOGrOEEtgB/BoWGskQ4aszhAbaqy+zqrcSy1ZqvKlx19q3On
AHkpVUMeEeFhOQK8NlBO18FNoRQ3XqaAsSifTvDajo/w3x5Eq15VLVV5H3rDc9PnW4g92dRbJdkL
lzXtXEDP8hMcEHGgaSKL5Ok2ufQAKDdeh1gEv/cYYPXXbkwHk/w8JDuo9tLI2GJKhegkHbKPMfJx
bXXtY35HRbrGxBJIIUqzFAQSMQgFlmR5rq6Z+6oaB7W39g/+Bz6V7kolsbnReffi5EAzCmPRGdGa
LdP/lAWFaHu96xJvw7C7VuKOClMkMSALWaYUFzUIaczo5R5/ZKwnkq12JsmlPyo0lamKGvagY+EP
q3Qa6vGNvR1130ehHoPLxs3meu7KarUsqR6gEpGzZpUcpz3ZIAEQa3aMfsAAmf3xPj5oY/8r8W5D
ohoZ3dK8wTBM/UFji9MuC/J0TxbLVRLpyourwXvtAZ6TL4aCPXGvGp0KyAwtg7agiY/zx6NwY4aT
W53VPxp0mVuIHbOBpTZ0jgZl9jHqck1IBkQabwwZx7zl+HeuV6E1eEXHH/jS6OCmDh5ECMfH3R5c
o/OTPSW51T6YMx/jFnptE2fzAZXh61TTT44T9kGUTr+5ZZRXVmWk71X3cSJDbIRJWE6BORqso8JB
HHAWQqdz6lnhqFciBnQ6NTrvC4qbEwNIO6sykgOkXgSIVTYOFUi1hyMTZA7zW7S0Ga2rSrZavFoL
lO61Fi6qHIb4ufrq62fYA9+daeNax9xl7O4Ut5XfU8qdr+wIkaaK7sjSnbt+FNhvkevknkdXNvGh
l6GQ7jFLcg3cWj72HpxCwgsJWx9tBlQq0Uy4rB3J4luP995RaIIxwzP/aj/VBMLtI+Zr0FeawPrt
woOvyyoMsLTGhSOlm5oMaXWtEL/VBhATe5A8p2E4H/fiXxIm9ewoVlWptpV/aC4m0+SianNR83wa
Lakj4mm7vY3TMQBHJ+x0PRloDlde0b6u9GfNl4jlJ72V0JCOhBNIZGv7Jo8UAnoubd3+KXtFyIP5
DQk/HTM1LeVi/wGVOmjsvaaayotIivwLsclDwD2yoZie98ddVDb4eN70s3Nx9Tu08SOClBNscCWo
q43OPa3run1PX5KHDtSkoP7FXkMDRzA5/zwn0i5FMK2370ZOm3dSlqiiAWaqr7kC70M2q9IfILrl
Ws0i3RPlYqjL68tMBzkhJekZggaxTrVxsshbMKOb3iSSU8bWTDtzD1KyfJqr/PmKnqfegaSniYVM
lQ8MKtkscZvXD6en+whRWsvCVFMS1Ry+ItRL9CfVAahqx6k8nFafdgLariCcSK8OipaOFXP3W6Ce
rbshZTvPMGiFSjCKYQzeO2Z61W90B48vJa8Cb1vfsVzlQRlFn1P9DR0LMpCVaRVCZhAGZWLlVGMt
tiCBcUXSnMssNcGmrevQlNFLPslOSTMkVbRfUryZy8WMjEG2m2Du6MtD3v+xYS9QNfcPHadRw5/x
RwCJRvKPadgq4yn2eDe/8SWKCrR4zP4/S3q4cJNvgEVFtTva8Y5ZYNMeJjaFsOjgF2nYGv/qweRo
ZkoRSYsWsf+2dKikQbkusEhfIlhXpn64WJUpX1OFwQ48gwcNcgU2dl3i5pi0ulPy0vEptCMcfB7Z
k2nxSCcBp3l/9fjSQtKoCD6KN/xvctRQqbmCRHPgWkRmh3dyRM6TWUx/wOOzeXo7kewquY125xxy
Q0iZNO+Jkp5ZPk5vvs1UIzVzcWlWdx6JF8uNYJVdkdDXGws8HJru2JhQ/ZJLWjUwvlCRDBJkepjQ
3L+ZqZzYu4muQIzcoVDBr8LD1MsTVbSlu4VAxxYnMysMCBls9qHIE+SgFHlwgdU5AMcgdoEQcbpp
kL+pkPxFxuajJqtHHx+HEuK0k2LmR7QPADefgsFCWuXBrIseUPeXtkywqsQ67WtoSPfD3dnmRJ1y
gMFlBaeHsV+9LomCGo38eICTagebh7VmhuWG499BtnqpTw/Os/u0B6OD+LW3UvMbmp/gG1BJkAZP
bMeQbQhLl+9+6SaMzFZPTmiAunHbXVRvOizmpqGchYRlpg7z9Zkyk27jgj92WE84v74Tyu3YY+hc
1wqBNeiiPEaKLbFpKWitbQ2b5oqd3gjtCsvMveALCXxA0wElevYvO0PZZ3Qp7aOe9a2NzxSounX/
EFhY+Qoh4VmoY8MvZiyW+tsgY7ccJ8OyV//uM8vd/4LvvxMIxkzNBUVY6uDkX8dc1izDYTmiSK6t
plWVVn/AaifGBc5yS1xMZRYLmoIuJpS0UWmHerI5s4gxVF/Megj89sffTsttfUbQCodj8AMDRBe7
EKfwGqd6kEBaL9vcTXE205jDWWNGQsnpaheorl4COfKjln1wW8dFRMUySxQKqfkuQFeMZc/qGQhA
qahgTapc5MjV5boWC9zcd4K86U0QlSepmvjIn6NE5hJE0gKuj25W4HA6dfdLpI5vrwX58mQypmr0
TRv9Fabn24dAE0b5KXz/MqAVDE20tNxOmSQeTxn5eYJpF7RS1CBoBRElkgaxof8VpBPkTJh4i+Zs
JVeDYuTi3LF8Uug+fOE+ijbFMovCrdoz/u1w9iH4PKUicoFUVrx2f3RNYJWttSA/Lc6EqQahGPo4
M20mc5pi9lHKD5cRJNr5ScFjoiQLU1oPOXMTMuYzdMEfoSPOi9uNpBfc82oQntz59bgR5KsvOCyz
FzL0ZN/+awl+mlEc/Wfa2WhgiFuIa0UBpOZ7u34I8jI2KBVpL5YU1/fdGPQ5NcD2vNiroMDKxxVg
KwlO/JUfYoJRfIXLatddBBb1Y0EHWzuHNrnGFE8jJ8Kd3FqgZLaJy6beUELVu6NoSBugWRY9mRMV
nuUPzA6cXzKp1ZsTgaahFCpzSF4wo6W4ewftIqwbBjr8ZXtCDWk2u41O+4aqIGucPMD9MCVAq0N4
scneEX0TtDjj5afi6zvy38jFGCCBNNMzKUCeKxTxXlSh/MpcfGQkpf8XxN8gJurbOWyUbrtK2a+l
RqTwSx4tRWQYmXFLi67ReX3DBBPf2UBe65q4TZNFhLPrn7/h6n18QHsrXfSXxbkbgwKCa6c86Tch
8QPlAA8nfZmJs3vOiRBLgbn/mjUBcfTWPnTGDS+LhSR0n23QrxC+cBp3mLYPNDqL8GafVqAjcO8l
jDlPpKRNad8I0ZjSE/KLyf8pXk7oA1AHjrfM5PipIH2DSl0bihMCxE5iNgHpx+8f8H3KToXCVNxW
SWU+esUoYHkPfCEQo2cgzXJMqZy3fPimYfPzEk3cQpG5QVFI1XuCQOXWxLeLhqBfwW+bUe+MRyre
zRwc8oglbeGL8x62MMRAxnQ+RyYOZFntejOuCDvo+C6q56oNORCCLplxFKrkMc4DvgJke3JGjJPN
JWoVP1qs0lSgWJ2qq1uJX2FSCD/WReov8eUyT8rawesgt6+dX2rwpaOqSeGcLWIKdiY9juT3efdv
zldC5CgeoAMSBxwl4gETdfOvJwwtMnyGbsKH/NBzm3B+qYG7HMOTCWKhCIiY3qFdp1tqCsZnmQR7
X2OIiPltqhI4DF4OB3uFtbiaPhRqvX3iLPNyMsdxmlyXIj/DoJqPVlLppAzfo2UQkwYiZ6gLhqms
P4VFDx2nnjF7c8asgtJc+NSZV7MgcUClfgsMLRY2TYyDpot9ag291mAtzhrmAyx8vkTy9pvCiI42
nFX9W6jDN8RjGSDnKdWz5KXEWBzg5Qz28v8JJ43WM3iTFikTT7BYZLuiH059fznQQcjvYSg2ew2i
J6kkJ9YydxCfD7oDTHaioMzhxKw+4ys2tzTIvWIkS8MtPEdDFOs5kFWu9Bt17tBl6rMWJgLqwsSh
Ec3y7sO7l5dDgWIF7GMDvnx9oNnvMUrQTONa5ZyedUGF02mQD+VK2/Qgc76FE1vROU3LcX6TIrUo
guQaPJBv3g1ZDtUIUFN7ix+nBES1nOjXVq8kildBevYHIJCaUCbDU7KTvweEFbW+HJ8Ft+c6NnkF
cbFNDol3xCkRTDHWluML1TpTr0GX9lCEqFZ6tiKga256BE5xsvsfQXU9W3+YJHHqReR01qZ1ppqB
R+1g76eIaT9O67iUFFqql8VMfUFAkzUYkXXY+0XI9WBVYcrEIZx+rh5XekbM/06O9zxWOWRcobCN
uQmAb2D9RnJ2SK26jbYb/qsKF4Hh7ewkzIZE24ujTfDYblaE8u79fvlLspCz+xzciStEmF3t8Wr2
+X++sUhSlDsegXVpDobiCvP8aH0GYvOf/ToTtLiIv3A8qpGTgSs9/4/QzY/fW0WxMT0Oxf9ls0Jt
JbBbLp+zBer9+Y9rrkduCHnclxrEUTMLJoscjspgspVrtHDQ572MvFpK3V6PwbePHJB7jA6Gffmq
kALgmsEMZO5lwYpz6kqH2drWTsrLwF2Rw5EWtde4QigYs//hl/tQrG9frSf7CmIe26ZdJmRwSSLK
QC3epet0f3yE8F46m1+C75Io58nMnAMs0TjwlwCU+ANOETOjnQQUhTx3ZrTqMzeQX9+ZoG+GcNWi
rcCE0coKG9qVD3m/wUs8PmTE+SERZqsHHKBqQVQj+ekq5SSlm3tnXROWa/zsI3Um+i9O/o0GShqz
8AhvpsBWlfYFfVZzKTTpPwh/5JJljWabt88AV71zM+QydOqMgaCNCrNqaj4C6yLfUnvQpWFy63u6
Yl+dwDXSjg0EgRlz4dN5TqwHB4QDRwXa+NB16GR/qqzyIsq1FJP5f17Wgh3s6fXHKiCjYmRd4chG
4xKHUPo1QxnHRO2jvG5t9sTPtZ4kcnUHeCOzSsoMlzz3SpQwDeNEf8vsZlCuRlEm1DmaeFzDlQ6T
39xuOVOsNm32J0lhjrHsisWWqpQFW10geeoC/+t/fWCdVuefVvc+DvrQLVbWQTQKMkZQyOhAmqF8
85BY45tIT+LPv71TKBCd8J4s8L426ib9btBGoXEUbTJQ8farNTZ3ZyfIt7/2zbnYXBjsMunkCsa8
NWeOSUUaUTXU3fKDgSx7vPL871jdVDJlGuaWZ+R4i5JcK7SQaM380Rf8Va8bMzFfkJ1mTEp/TcG0
tIIJetqd4KqZ1avlrl1WLAu4ckGB1uhHdQAe8RFhftgORxUZZS0CuMmF/DZbO2a6F5QRUbOHAnrD
ejyb3Ig2VcTEMVbFzchsnpblMGO5cTcyOnn87N1tR9KHzTc0bnoz9OQ2z/WPntqqoPkdufQ7hdNZ
E7Pf/9tRQM856zkXRn9GS7bmJ7/lsMeULns319/VkaTaP3ppe8bwnqh6QIvgS/IhtxeBXxHxXvnk
E55JLkpKBmsVJbUkBIwIqh4HVe4YA8/a9piwBIm/rUNSO+pgbFoX4tsM5JmE1u5cFtIajtUgyQku
euNHN4nGycRjJLxAJ6l28XtTsG6fjxaCewnNj9Rzv3qFcBUbTidGcxoMnn6EfG1afI1y6bcJYOTM
dXQMUMJOZ7sv+1E62gXLz0zJFFhpPP/ASPJN3+i0naHE+Px7qPHPVOqEqid52rrlELNuCP8xnnyu
YkB9/Y2KE3DoDUxQGHFmL+Lt1nAWG9wV9Epdd5ffORbLkKmcNszerU+MHdxvaG9u7kNsX10CSYXd
Ly0QTie0QoAYGRybA0FcBYS8qLyrcg+lX7UkU+zNq6IC2D7aEHcsQrPL0cgsJt/eyU/k3eXNBez+
QJUPFvJw3nagkm83pfNfxQvh9Z38Hf1JJHmp96pQtGjNemXYdXqkmlp5ArJ7SuY/aQr02rl3deeW
Cze4LvBQMCweuNa9dxJweJPQSvV+blgRsan0+9YXCQr376wAn7FSXHOVMX7M6W41+rR/ri6XHs9a
2wWcal1j4qrZIu4LsNG8tC4Z12k/1zq7sl2I8jUVpZFF/e/X3yENebQ4XL1f7rw9KSBY7CH2AMP2
LdxBaTJ1YmOQ1SfSSVnLPBo0VnfSkuOHzL8ZOhCXyX37boygZ0hRS9kmgunQSg7uuQXI7I0IYw3N
Dr4OfxGl81vH/Bkq1coG3JvXMGPVskm3Lz6FLMgpkGes2jRJUQNSMsHemc1YOksQbLo7ThwCU9de
NL9Tt2Q7NgnDQfXbwaDZscNhXQqTfGlSLesqxJuLlQ3+RKCSFqk5TIJMuBY6JzBfR40eei2NtZYK
iCWflluS8lnV0xsUdUGtOnlPbdcJXQ8NSEAlFMYkYTCXn/WhlT+AhFuazbvbfqfcM/lQr7NzSsYV
5ocvqMOgHXP5utqRjHS9rIRLDegZaDVDl9wrj3ooPkzRkieZ7fkDE2H5erkX9v/QppHXHCi91JLF
tMNaUQ51h3SRhtKcRMbzqstC/UdHkMmH/6ziLLUG7+RKqMZDLMTHYGG78iuOWiymDLepz4g7NoEb
9Un440AbZq/Y+xOM084zBLQrtSQimRHUepqJySDjY9mL+KoJGSNxGipJLk6VsZIv42f9nEsVVldp
6d4ULlfVto1uBpTOHIZ6vUGhp04zPEJsOje2ln58T5TZyQYb+WFo9Wj7SvDNNfLMY5budZkl6max
h+18Ux5wS1U+09JhkWTGOXct57h1N2SnmJQyOOLCgGv0qn54zdKKGakMz2iLr8lUjb/xrLHtDyMw
HrLA3oz6Ypdmu28MIphoBkHH3gD6po+676U7lh31GLwi3K0/2NzUdCA3mcOrDBzzow9b8yRhi6R8
QlA8sfQXMvqt3SM/ulKF6doUA4dls/BmOcLPymBLh+tUIke8IUii3r/vka7KAnEnm4BDpMhJQPxl
I4ErvYG0k5s2Bl1v912RBDm1wsv9IPlRapYns6+KTAxKcVtSA3zN6G+KG6p+jmrJokXGwAXRah/c
3WHvvhCYMr8M9/DS3ZN84BZuRrdB2icu8IlzTmb4nc6mXcZhbb/C0RcyML2/LvGMBdqiQ0jAAKPN
ZwrZ4rP/yBbhPsYa9eRnNdGl7IDtDaSwNPvaE8qJGY4a6malVF53TFTmjh02g8idVMHbLxrd/l56
jvcAsr7CxD9uLEhAJd6zsQXtF5OCplVt+H8fTbXXlfA5ad+4TuD1y9gY1zkYN04NzVGISyWodg0/
G5eRVEHx2g/DDZ7jI/DLX8I28SsYkqQdJyfUnxAaIdVfxodEb0vAM5ZOxA8gr4578psM6y5JzDSJ
k9MXzltXb6/ut2RQ6spIbK1glIeo7AK/LViOymS2DVFZwavBz8f9lq5vhDJIwJTqtmjE27wjwhv6
HCXSHCb1pE0r5NOTWiiz+cdiZheFgjN/wsbWyv3T5IAA+9rZd/z/og8wj4cSdARnqmnx9f+xzIm6
CRqoZI1nN8MTD6dPM5JNUVPFyE4VZDwBxcM7styFnHzSUy9bJZ7mRnJG8ht1BlgMw2Kxm7ytLySR
UiYIL08lAbm9Wb2JBBSJK2aoOV8JGE7aDTeGVRt1QOnr8tQrjrfqF55F6LIxKkSLxNtnb5abL/w1
IQ6X9yhy3q8oTyo5J/IkjzJXsHKXtPmZ5ahS4uXX+UypXnZmKf7ulF371+EbU8eIh3o3eaSFm+3q
546CONrIUSlfe0nMxyrMLr+50GpNF16LPST4trCojymtMcekWua8f+4BAaxqRojGAkSPdrGSAG+t
fqRPJFKVxdJmDqYlwDyYl0RXs5i2/LXruREPVKx3ZnjZDMM2duQ9GwMw1XrV+PAeKWuDEDhb2cza
pO9DNTUuLEl8EnFxIfYa5lyABfM72xYDU9y6/Zw7yBhzEOdsMSjoQYg7gjeTIlXWAMMLje1pC1RG
4+TXvbxltJAerU28pVeswt7U1nDWSbZyPGUQgojIPNXkD4my6Y1q+SVsZlaxiIETo5IB6fBJFF6K
BpcghSoq0h/7bmtm9dkdI2ccwr/oERHr18kpsTytLwD1ZDqhDQKIbKPlwNhhvQw66DtbMyIVcet/
6wZlvNT7O1DN7PAxFP+NnY7khTBsFstwIiWd5BnKo4Cx7w+KG0gD8iKI9SYEBniQoGQ5YrcSt/na
rtiAFTbjXq4kcc22z2DH46IB95pGXtTIfj4rQDPH9k+1ELJt+40SFRlCWzmFoHBjCLRKiyHmlLFh
jM9NFxKO5zRwZMv5aqRFnvwAfAxnO9QNZwLG0oK4007uNkUJ5oBMgQX92ROgJz4TGTaApZY5mYnt
ebCGaqVIdpKdNQAyb9pRLIpurs/olP6+NmYSsJT+3/8toO9Oc/DOSIa/tYZVN3KcWRxOPeWGZIoH
nK4+Dpiy7ExyUFQ5ESTu7WlD8X6Gjz5UQDNH5YEKZ94HJEWdpVNwmnXOpwHPSarxomzZImN3AuuM
meI8ZmYECZl4KK+EMqnYLvjFbit3Ae/v6peNUeGlpWE8oVhh1gWxPzjqi+uPXRdjK8WzFI25KAh0
0G31/JQr7NIK/v/cCF7YqyWPrgWHlU6rq6Tzx5Zj2ho2gh/Ta/ACUTLPLRNRNGk+/FsBZ+FJCUvm
kjCLKbwnnRdNcUZuCXGO5JBUU5dp4Qye/sOoY/88hqRQwtivVmQFpINwJ4XYko2atGHTFkmRZEBt
uCbOQ85WDJMIEoxwb39jWGH8Py1/un1igVSUY7FIHkUS3wdqeyhfWSYE5eWsmvaYYAbKTxdYSlZ5
Lux2/IQ2aSVBRrsm1zMHgAk3Af8j6ozrlGOzE8A3ujjeArcxozVtbUTlPYhDe6XPvijerT+JTY+1
u0l3pDuRsZF9jqUk/vzC0Q7LgVFTpdoFcFQAfOO5PwKHFlgzOX1Y2BcAnhbUzN9hTe1ldSP4H351
tlIw/vS02zuVKAeXOhACBEJGSshGCLXXXIdzghaeJMtI9QP+V/1ZrHZwuXid/AkrS48LeWRxsby8
yyDm+CxQRFlePDZq8GI862L4PtT8YW+/o8xvAvShv1ZfFBqBTvPrA/f1LPh4S9mkZ3FwDm93RfqM
VAnfbhb3/mUJOq2/hQHN/49PiVbwfY8EFd1u7XsZlItwwV0BFANBbV79TAzUDXiMMIN3FZsYAVop
3CCM7WJCAz8a1olV26INCAXi87wtexgHuFcwEaFPLDvlf6/p9FJ4htknCOPYywsli/H3DpIgPYNy
aDAuJkexpf3HI2BsCCsj7/R6zkagPTWmUm2M9BEW+BfK0DWIk1wPtdflcIiwK7KNlA6kfqxOoAA8
0nua2fJIY5bethvHY5bSQ+lxWtTPWPEYSGGqSMr9DhZrfUvq+KsXG3/zklMO4CTbA7BXkpJE6R+8
nCzzWK9MKI36TxAudJh0sdjfIZGXdy4WLtNMpy+Gyesgmh3ijRjt1aNHb9GYpEWrWXzxOhCvx9yS
5JasHysTdl5AIkK/jhobWrjdfU9z13118miPlZX+Y9ljU+VZQ05qh9FOpXqQvZMADGs76UHo/1ZJ
k39hu86ESkvCPi8Zxnmt/QnlCCpmiHfpcwc2J6zs2nZqBRXLl8DXP1W0d0aC8/u3dT4SWEsT2HRA
leA0iaf1zZPIcU0K+9FQxsWtx1L6C47d3OWaPlk6mzHj7bfN1lfvJkaKjVhE6LyEDvpuWYxLYk8M
EoSurD+UYJ4K6mn835PzV9euuK5FThOB994OJjetKo7n6n2Iz6kE/lsgKrsias8wjOJLza0vYyzo
Z3TojeUKFRlIKV3EdNGaocP8s7uRYJe221zXcldxmoOqEbnbsvqnmerhmAUhO31AUO6ggzyR415N
2burpLgYHesenMxyqM2o2LoysVaAPBd+ADvRC56wxBPymLCx/SkQOQ+no7UA9tV4xR4objdTuocM
mnFbeUjTKV/aiZCinDSyTU/Kfc2UxiQ5+FlA6vHtMxU5Vz6Dw51QDBccme01OLuSH4Vp/BRIhqKt
C9GF7AoGJTxtfrIF/nwdPFDHjtnspCUlTpwQYBa3Qf3rR0FwoXMlfWOYQ+zcojAny+eVchkiB6YB
o0i7U+aXWm0Ag70yi2qP5+AXxq5eSIKpM0zocatLsoWKzJowOlp2Ij/2gWHaP8pp5ua6N2ePZEx8
oyPBHRkYDVvjqd4ZJGsLWplZlDgByGeynbGpjxBwOtAWcsMA3u1xyPEy4gUpxPgYvSiUEP1W89U5
+V85ntLd7w9CB3lRiBemR40EWH+W8a3KEkIvYiOVl7SwR6Jf/Yb6Zv2YqxvZ7jLiHruYqozXida4
lojylQ7jd9onhRq+p4mPtcs9lYWZ6/a/6kP3EaIjjPJWaTzAgC7/emCk9CtOStCZx74lI5UO1hrb
QN2Ny1PoI5OLByy2c/8x8QnS2t13Y2Hx4EG8VfLmko7tO4yiajuXk2cjBgC2MQiwNi7hB7UgeEHt
MM0dxr9ckebGEHdnH8sLvCL8eTI6X2nlLlUS641SZhOu3PF18wZklgWgEOWDGACfW0kUxtkH+4JI
1eEnj6qkPNaIuyDSMK8JRm8JdHRMc45mNchIuU5R1Z6avOzCNWRxIIpNx2T9yhY8WlQHhcWrkZ9G
+Ci8wVcBQnlppp0DjR4B6q0P0mfxQ8wumpk8/Wzsk33bPtm1G+xf88WpqLm8k3BliSYxqIKl9NkJ
rQQGK8dyX7xqP2y3adMy1GT+LoOhzkoiCWzKvaAfbsg82hnS6Cd+cMv/RdG8b0vpMmYiu836t8RI
zEFSocbqaHhdb3SHeCtkwQ4rD7VVQNGiL9KiAr7a+JSG8uUsncHT2YmbVL4c2WyckoscfGsSqfLy
9ECQadnys6Sr/R5/xWPZSQlf9+1xwvIezQr0LpQk2V5rpu1cB97kxot9Ykab97yV3WhA8qOCt8km
LhAwrOaQdA2Qkow5bf1pTDuM9jbh+xSvD22FsiYW6PXLHAzZpyn7Id68G1dv4xfLkPsgcfJpNK3Y
+G8YgK0kRxKWlmevo6lfFq7Ze1aKAgJKPN196QP8hDqEtIB+C7FINhA/W0HXWeqRxP2owLe1ETrI
9gTaB/Yb9ir5Hpzdsffqw5A6DJ40H9N8jTmbgY/HxW++nUKEoFrZdKBdX5BaaD+iRyNEZlNDVkW6
6Fag1MNtmhgvItmtyU9JqixDogNnevYaZjA835jxWM2cpBG25esaXiO35BrrUNmmc8U94ckJm+k7
1XwMiYEUhAa3XFcfhk5z+wqhwhqNl1SUvwxhtZ+9rVFRRuFWC0fiDHPIW/rT8g0NJXqjms93E4SO
/EeD0WMTfp3k/Ifosc/0jdMkhVxJ1NWW7pm6ig+YnzSaOjbK27c+F4N36Gn6mug+9buWyAjVQBd/
/RFTPFO1G1j5meML9ho9OmV9v59QgcfmXLaBij72lnTKS/hZWldjCgCtsPCAvNESlhnr26kxYgnz
m/9ZJ+IVLONeF8g9p/ThQTFySF2SKcwYsIMIR7x8pZI15uLOnEccdo28v7Ozya4SdWL9QUrEcmef
VDz/XjCL5tzY3wfYfKromQWTc6CLD9hCd+XlKhkiRzOm9RzeAdJg0IDT6iHxXJr/O1FPS/HH4lKw
qsFr5/ahk0twBA5n0fsPx0bVuT66tlkHRzG394QeQSJWzXmZZU3yeYalvSZX1yLZDO2n0IXwFRSJ
TphvY1o2rbgeg0bRaa9ASqLCojhUrvyIk/6a5HYpmEEeq6QhdWX0fiBysO01IMZRB6uUcv7/K4Ki
HMhq6sYIvvKvtfB/kmgATAGHGFN0I4+YdXt6bWNXU+76flYzjoLXW4SomcAQD2HZ4sEAAwpkcWNR
q8oPayWr1YMD1dIRt0V5OON8zbaVaGz5GDx/E6vLrhwKE7t4AxMdb3SZymCa4WEGX/jzJBPAywuB
vktv++55XsgsPgjvG9157GuLbg6szTpm/QWgd6xPvjReZobZQIIjulNS/nC/+d1TV8hFgRIidz4P
Vs0JK34fuAPbKQz+K8S+p/Hhva7OcK9v05LhPnLMAp+SL0kTJBz+X9pmOacOmkw3IaiVtsJm5qfr
2TcH3bBUjWZKbEgqpBY1Gbx5pIH4oO3OTUPn/nZgDnr1avJVF45y+WM/OaY9ZypKDfsexK6PIfuR
TFEA07b6XQiuxKFzg1qX0Qn65W13J/jRZD2lPxIBV14ZfhVJvPvfdO1lDNh1yL5KXAomjmDIChqA
pGfdwKZ+dFAlGFiqveh21kdM1bDTgJtO/Y2ftM3AJ4NYNhbGcSRK4GgUrJ3qFNMUhTSqJV8VosVl
CcQ2hT6QVnyNmjBzm80TxOfNQjTXaJRTSeiuCrgSEqoEgWJmKRUYGQ1JE79INjMrJAG8se9yJSmQ
NoH61XSU0CauCx5rvhC+Agyi96K4NAQXegWwM9U6uJbxNOPKo4OFCxS6dQrCmqZEqVEpnw26tVDb
f4Gsbk4UzYrXMKmgde0EF0k8sJTuCUKpaKTQ4dqcQLoxwPraVoT0EOdlhetZDI0YxM7RmYcS4YU1
AvkVCo8surCxRKpg7pRJp7RlLpFXTPzbVvD51D6f6avbDYKvI1byIcszJIQkPjVDtiDMQRCKVh3f
MgC4a2qW7V/bomK6aTuN1MLQELFikTcJnLUT8mYRVGbWXXLsuL1pOWMiGq97oOAVU9dpIlEiphy9
OEQG8bdqiusRPHtM3CWz90fEBMImsCRv7mm3u3noeZiMPLCYlS3Fzn9MDmJf0dDGn6dIWKPbF2hc
fGKw2bhquBebOh0s3mb0TujUEcGExZu8PokcVr1bKwleWHRvdTmXVS6RWuciC0UjUxeN4/slQcv7
gEpamhzbuBFu6zFGeckWWTBCeHQWcrmvkA4kYnX/PWRUbxgINoOYBwtXRnWCOkLECpadkqxcsWJs
CgriTpoKLwSDzoSWaPAunpeZFSVX241zA1CV71+6bcnfB4xWO6Frx4vjoJ+G3bvHAOrCc7ZWCNR4
8PY/ixsCtSPxwJmhwzz8vsumaXqF5J6EATk7gC30/TBLE5lnJXJaFBJWgvEUx0DSLD1AQo7lUrkv
Q6vGwNsGnD8YcchGsgyzP5HnIz+BJP0AccatKv6mGWQlcsoO/7FFyYMi+a3uqqKZ4TAYTHqbV3vD
uvjxmrBCMp4azz5qZI471p68B59VwPSBxscvh5DIc5vhvyDt2ZFmDJ1PFY0aMrPEK8NPv5byKBcs
bY25/qP0SxcZXfx+i0ofmXKsbP1MjAmBrkWXWqwZeJ7gNn1MH/wgIxxvOLI2cAmJ2Gl9iIIFwKnv
Rv8rq2vMoAi6QldJCdK0om+XkI+gKYu2lDRtAy0x39UVPN2oTftlFISc8nMJYw26v7Bt2Q1yvbvA
GaSzGvhwhSQjIbEjLyRckSBMrFnY9Kovlp65P96E3aCzdrSPaMzaOmsBH2utnmmnP3bEaMszjCrn
26MyXImgvolOP5bB9i1lI3FDBSVHos6USPX66/1/KI8LjNUq+xcGqg0ZrFLj8RFRwFaMcs5P8LQS
aGS0iMR155oTgI6pFWZb3NsJ7NaDMX7lsqufI/0/HkAB4tfSOflD8b1oMejcOJPHPx1Q1kVpLERZ
YKX/tGjvjGkp6kBlhXtMFGCKM4vpfKjxIu24FKtnN0fVyIsNeeoFEtG55pjmkFKq2Yp9m6NsTcKm
P9titqhJCB4CNZi0QgOOAUgYceLIX8TOb3juvt+PZOcpyMXQ6bpIYHfedF1+DgZ/29DPrgvyfTsZ
+3PwYMDH+L7CHxH2wTIuIQCcStekrD2+ABmGHWhXu2ZWqIEsOagxuNye/92Hw86EXwNz5jbhzKn0
a8Go5h1jchGHrCT8PDJVP5EesOGsTd0LKoWKXmRLKXMrvDSdfPKTFThBGj9qZBTxoQR2pRBNf5Xw
juafw9o41C9DceI/vJ+nPUyYvTtNUj+XsHWjqjzKXBuSN6KcPclLhvUHo323NLLUEESQO5+nBF3n
NJxqU8wJ+MRBwp9TxELwneUJAu41TxXCnr+aidIkCPWzEBsGcw8U3lUZ0xirko3teRcuOXR1iyEz
gtNKDZ2sr0GeKCtljIPEQ7iY7SSrumf5g1qtgUdq5QUQ9Vh4xmw2Jia0bod+JjY4n5ffmSD3j9w5
1daZZfDTK1j0axVtPycgHzEYS3ab6tHbXBnCODiNrUZW58iXocxrMjZGer1YXv6nrt20ccCIUPSm
onBp9puIbr/cX/CmAl6IW+X41atqSb0EuLjeghbmI+TLR1bUybYxdTKiaAEF9Qj339fBAvWGEvb6
v4ldqnLJDBOWjQgDPfS6IWi7DolkUQAKWCCIMOMaIwnz2OcJAZC09MGbDbIm+us/OqHTYhshIugo
vIcSwJ0Njgvn84rd9WRtNH2xbOYN2lizkN8w1jmAVxrauKXs8deQEsNCeKjQ2NgvibtDfaTsgjCf
Z+qlRv1XF9PO9m5ZO9bASrUyyW101Db5Gum45BAuvIMfOoNVZKKM1U50k0Pi2m6+/Quv0KhmTwHe
AsmsQenJA4/9btt1PdW6Z1j35OdUFmvH0YnuGLqelDOhVSxPyz5xbrvHafABX9CEGAXhhBos+tgr
1RL/6KnM/SOSe15G/vWwg8cVuFEpdWeQ1IiDt83HQfg93dhwDbGBx6y79dtummhnzgduVrM9eLSz
U/ifBPvnShlg5O/juOTtFy+7tuiXpIDwzU/8UAFxZ2weoCua+xPXgF9K97PEXgBmxmvPrInSDUHa
jKN2Bg0ElaspMJIw036uNqm3+2lgOUwPmRuaRaTUrDf/N2QAWM+Zx/nu2Va8lMlHQCesiagXy/Uj
VyyUg0/Ng4BlvyWC9Wpjtl/bYVnwb9trNiSf9mcD24NG0XBWHULmtzpaNg6WjpYZikUNcizDqRDM
hxj3Njd4mutb60P3qrUe5vbsU6m8ZbPwW3SFf6RTef/MLPnoflvxcotjSsTAClTPKS7awovpSovp
7ukDV2ApN/KSCezEOXV4SV9Cw/PO1R3fllObUwG5m/S5D25TJfsv7ua4/yTO6r3eCdtjGgrdafZs
MtWx7c/GV7LvXxRy2ygCpf7vYz0MtkrkNirtZNAM4QRAA298EdTtsLFoGhmoDR3u9DfXR6yhWGIe
AQ6BLdHxEdrCke3YbKPZjmTyNEk9RgARWzHEasvIGgmWRPOlUP3w9WTvvIRVKVvY384WCqzw45Uk
1nHiv4kUtoFE8MsfTKlWI+bKatsDhYdHb7hiHxCKfgnGZzRf8pZiaW2NxcTDk39D8a1VUVoWYJxG
pxtffjWzCmMPPFlRffe0WTrsO3r4nzN3+CviXe+t3QOWgETmiKeN9hfpfK7fRh0m3yh5KkGV+Cdc
uCJZYlxynE7wInOSbI9Z8P5IFU6wDHJlANOinwAe04eOEVpfdPsVd9QMp2u8uJ1qwyaP4zBMXGHq
1fMILye/J83moRKIDwj5eCEmzYBi90dr67dpW7cz2v2MzfWFhnFQrJIfcnyaqnZnc2fZB5fbusoe
Xdt4ri//eh/eUKqOq1lo3fqMhzBtdqsijUdqPBG2u/wBlVikvyLnmybqCp+wRH+FbTAblAu6HUyH
7PAkh7bhqU3s0+0tCLHFP+uSYZotraLwgLZ925kGk/Qcer/uTqPW7WRN3TuHmiVAViDNYVPXuVeX
cxR9dFjNNPMqPyqfbWeQ3g9wflr6TqYebkR4HGhNWd29XQXsqStj7WGdJDXvVB2JQDvFv0qGexQ0
zJrg1E/vifgXGsuU482rA+LSXWa0AcyC1cqif6so2j+XvG7sHhGYLlMgcbtgwqmQEmMzq2f+hHIN
aF2FQt9NC59qPNbNun6TOBSlOXHGC8KIfiCONIDy/tly+jz4zUiuyyNDS77xYljn3BhPxOQMlNeX
kdk4Cxo/3dwEufkgfeVVfMp32q15r/bFP1T4/D/frV+R5ypNsPnPowuWW0u6KCsJRDPUOwJRejRK
7jdYHiBvP95L5i+iZQzxCdgToGEmA5Lrx3E7o+vhzHSQ+Z3zaC/vY1QC5aCb2Jc6XHYpydCFkVDN
swM//QcbBhL2JNf/0FS6YVZCvdJ2uWgFKMVR9hGqOXAdBvNXVOWUGCmsMrXc/XwwZ+4ATveO5hHd
Bkdd2Ph7ztKDQZMXG7mMSCFSFGyqtjXaJ4JAWMAAqjfyVIqefuoI0tYTIle+Qhxur8CX4sXBQTM4
iUbVzJIijyRnXkm0LYKo4bhDRZW8tx1x0Gutk8JKzWRzZP47GNfJG2EZ/j79fSLE2UnGfcxv+e7m
1ZE808YtF984q9PWZoycGYJyMem1fAdDi8poKbmzz1tFull7iIkKx5rT+X8PMjp9BtlY6jYVGiT4
csGEJoP/whgy69nkKS3PFa+V5i1d2/VfgoVKjiUqKS9T0bTTs0AdcL8n1hdsrj1qV+YKtU8PhuOE
7ikV882soxdSeZulL3gZ
`pragma protect end_protected
