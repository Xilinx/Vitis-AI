/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1136)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzFBPvsMxaTJSGUQ33xzYW30z2Cw1E34VRZOLiWoctr9zuxhQa5bdkOEl
pW4TZ4L87AFb50WjyVc7MlUVCv83sw7HamofSe0vrVQ9bQhVLvlgvc2HQ3mblam53stjy/yF59bI
zvULEIECwCEMd7GTqHUXQ4WCOM4ha/0RdP3THXpGc99193ErMwjvnS+z9VrvkQ3wc372v/MAQnPx
qAlpPPbo/B5Zu1WznGAEAVts4x4BrZvHg6FnTnM7N98ednB6hHN+k/UBV33GvEbPQ8FJUtxOmpJs
YldwQRvmpH/aiWtGDpu2lNN0vys1GRYq3lPy3gX19NQKBdfrZnZlwG74wl8v/94ZKKTnQCrdps7p
2DrfkBr6FltkmEFWXiNLjmHF+WXolKGtZgykm+3yDJW4+fExNetshvWnxckFH6JKZeYUn6//7rEo
8jESaDVBdQxsyJ6BWNwSFw+oMA3AWePW43BJv8KzkDc+bMLvJyNnTrE2CtnPTamuBAJ4NNxdzlNf
8FT7z0wZy5fmcJU6DUASnjEv7nie+NsUSZLFQnNlNjZm5kmlIUpqS79dxkiKv2sle9s9ik/Cn1ht
9mUJ8kvYcORfOJOxzzm8ewJANOZ6vPQnH6Nn3ebmQzgb0vXBa5ZvmNsLIPL7rtZ3IZo2Fd9N1gGP
wZIRfqEbgq45e2dlADfa19ANACcNYis9FShih6HysfufkuvSH0Jckqra9XwVR0yZNc1brVZV1BXl
dSv2KQtTEvmuqCyCno0RDxtw+g3SwC44qgtPV3kDrQXtU+Alci/D5sTwfwz7YbOQBRmD/JYSnoFF
dejK3wDxyKVmukfTSJEkDTgH9JEsAZ/RZ3/0s0rIEhKuBZ2mNS0zHJYBMrJjGMZ5vzOsI2e4yYC+
bqDTw906hye5v3Z691m+lLIdYsQQCZvMrXdiBELVt/ELdswPZ4+SwUwfu1cgsC1T0fAlpKuLhzeR
vgEpL2tf3HMnwFCluUqh1fqxIthwYhEspAhzK3zAnEi29tQPSC0gIhHIfvxAoN7x9uBFcdzOhmba
sCxMQ1jKnSuRRWVB04VinqdnCOokj6ZV1veTzJvqPFE5lcOR40QhQgHEpHKndrEQRV60IY++/Ot9
+A6J1mfUVFp5S3+OHjsrZd9SykcANWGbhKvhkwn4mAxJv6WIS4S7kaw4i4sR4jDJpW2yPq40nSMJ
+JZ9bOaWB4IsjuvQxNaBhRY8vYRlEFOaYM1YN3JyPVCqcSAv7+KNrbwj77OyXqQr6nigN9chzCBg
FfOn7fPPSItDafqTYGbz/NbbdP87wOMADbOofFyCNfW81xU5rZGVGMLrfGSjm412FHuEidlJ9XV+
Hlye6XXdsB0uXvF0/hNXo8shXf1z6EaKbGr+K7VsmoVrPIEs412YGxsiB6eHaFyMSyMK+8F4oEuq
sTyNpw/H4V0Rd9rfOoLlVMDRhFB3Nn0lZf9qYFuU+dXAZprh9Fa0OD5UEHH40SEJgk3aO9g=
`pragma protect end_protected

// 
