`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35184)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vHvH
4U8dDqu02lHqx1v3Agq3S014dUO5JB3io4b7u+E1DXTwTlL/CmbkpmLpeDiwXjh0p3X6014+ofMD
ngcgQ2+PSWczLg3iyLRQYDUWjTnU/Ih4xhgZyUXTWwb0CKjBMAr6RqxgQpYibIOVE2soG878xind
ZmXWh+C2TbQ+DLYv+ztvZaVXQzMUY4pt49TQ6JKA4nOil2A9U0pzSX7koZjr3CfT7osWFJXBCG0e
NPEyMKvjlyTwCYrEhTARi9g9cULbg/T71llY3YVlabb/XsVnupQRNlzHi2gsJvw8Sz7fUZ0HLo5c
TvVU/VWQon2hcGE0ZtmtNo9FU16FIZLIkmhrgqlhZo55y9MKY4WkR1yOz/AEo9bJVZLFg5iTLiGv
4twYQTYpdv9QL4VzTFOM4C6IhfSf/u0IE/6eDsyn3S+ma72035UNX6s8AJ9mmMe5BLO9i7MKt4OJ
mqpln0a+XvdfYq3PgxTBmt/6YEZghqe0AJch06UI7H5MGF/xcq6Jhu+FiWZVp8N1D3clmoQO7low
Ak/oOEVx4tppzbQEjvL9uHuNqlXpmY3Cj2WX6IL3T/gRnGFmWfcq6r6WJDelYCVILiSJPS/J5cxt
zrsszSX0y/06QTMtWm4sbkH7QpBKGiHUHA7/k3o5ftQ+PJClML6azGY9z+8l5OnPIc16qRBgXX3q
qjupV9+DpdnU57PoXForLSJzJ2vDRrlIwTG/8N1P7mmyQ8XIuzJa+0/ZoF2Ib38vfY87cUYMrufs
we30phIc465GxZYjiUdWohg1FB0EAulN0n/MwiscZzpofXgAGXNvF1t7B7Yk63ftFTq4I3Kjq8cn
MV9jG1w+4+q+oMEsIJxmN+QuCxUEGAoPdZnKAD1GguPyP9Bglk1kWqfexAQR0oA4PiX9I+6qbHnA
Q8SYp+HwPo2fzdL0ypQQXy7CWsT/qr/y7OWgAbzfKjZcnrECxnRzQOf6h2Cedt444d1UB0RF9CoI
+f4qPbNkDCX3z2dDysHKl82kORk256+2MhDlP8MSkuzjP8FobzrNuaztALOZtlFLT4unoJQ0aoc2
IODI91dFCTbkffUX1ZIjixHWhfuQFOz+TBwc8KVgwrPbVQV75tCRKpwgzoBBJsTkHYsuaWKWxZ8s
Q29ohVhoDQZIShmw1JUojUB4WvCk6Yh05KV48IixW1gmNcIcevrK0BWU+lQHJ1EyUh5GzDkj6z+H
8NqX9cEoZGvvIWlETL/J3k9mYjjpqXxjh+3Qoaud07evUNfciqd5yARiLQZoo/yPRRk9OkAwPX/N
JwZvGoz7rC19KBzl7ArFX/rPYhfVojg25w7hZnFgBqZFAFV4V8C5Yver1af2hAPgl7eSRpUpCmBk
21qkAhDFhzztn+eXzfuUPxbkPKFqJ6Nhcw9PYp36Tn1764l2JG7H9noxOEOers2mXb2LQdIlKTUA
JswswOBpmXVLQ4ngeG3ZsEr2Dy+KRxBFBhi1o/vy4GO9pIdMCItJ/C23O3xiHGU2WkU01RzVd69B
mXDD3Xw7FD2NO9Dwr8KjAaHMBdkadmdm+kKhn7ziycQj2uMpSkAhuvRN409/f9pEPS6goXtiwVTq
jGX2PfL7ODf1ES69WgP6uG29mFXulAwoItIdmIQu3ici7eL7ThzT8jub3DskL6RaZtw09Haqh0uh
yKvFcEkKOqkBDdy/mkhlHVBtSnlyqgbLhFywdJDQPcBL/2ztyr3VnNL4arpM/XhaWBYDHQSQi7pf
+1mC0XETY+koyy5QXPtAR8YmCIjfP66nHCmZhBoAhwODV/j8Tv1u6qKmlRN84bH79uLRwngbEZHF
NFzHD8WmFf/D4A7hw719mvgbE+hJRQBRkSv1vmJ/p3MhouZk8jwZD+XA+GcD8MEpCZInjkg3ZTSH
YZV0uG8I+lshnQq1oOFm767HB+q60npa/hlE7sHFlNQHZ2SYfZiS0NO7yhe9QVOZ3GopvM4Xaoe8
F9/txYueUmBgXKcwgYI7T073lRkl30/8QYSTvh678qAZMr9KjU+FVu3+1b51rwRIk2GJAO2G6Dd/
O624xHCUwJHIHNClzZCl0Y9Z842w450VASpSGCHv1NV4Uo2EqKEDPH/YuXFh6lj2UFQoguChL09/
ut0G1tp3rYmiM7FNQn7vPPqDArWyIHO3t06Fv/ET2XlKuaQrdvrA/0Z6PwFTmigmkBmJLCz1GgPV
epH6Ee4bVppB+PyN9/TTdeVZoKi7ynNsldTUZVv2H3sAUpv5kgyTMzyXlRpWmtDcMpDEtnm/ysLs
de8ZH07eRi3291OsbXu7F5qp8PBl+OrYaNqvWKF9gOKCAN+hmYtB9xzOHL66UJvYWoGwd5ueNTYG
8Mrrfvg6tJer93BMm8gV2l/OwHUc7GORv1Y1W//RzGGTx7Q1Wkza2aJhKOia0EFOx353SgFS04Cb
5gL4oeSZejirbLKhE7LwHeV/y+S/2GpXqk99iaxJJ+ftTs9+wYQ2OUzLSQMJUw+hTT0wFwuYcpwO
WoGggHHIZUhgAlkvN2oa7VPoSglTgcTxgpF70TGqvv995JltZoBCNdUxV4aX17M3H3gw4EUoBOMp
tPHUQP+xCBE/NtYXmY0YO2uw9PYKhTGHW+d9h4t74tk57NojUKImnqGw5DEf1QASY6N+mpvXWQ9T
TWclbBiYMeDMNJuoosU2UDdzFoZA4XppCzcjoa8BbkqDUYC93OMcRVyu5oYMrXorrAOQcpw0L3Vn
GI+zL2uDTJ6V74u/ne2e13i/iVEq1z58/EIDN67cW6fKXoUsI9sL9b8+STHHKciVGGnvspqQFoYp
fhQY9nDsYywQIjO/KzCorgmHSjH6u2PATjHqkzPApo8kBuOfLQH2eP5XrocxIDUCT+qa42BEJfTG
IFO7njBJswWtOJFCKOn43ELDNbOYBaLYBeTvctcCwetRqO9/AefQ9qMIKCUUwH7qJdUxn5orMUqM
fL4pH6YaU+PIGi+ms0okzAN9HDCjzqrzXv92aZE87bkH0EPeeEkeLwbLUNM/c0n5J3eaRnC7FtBU
VmV5bMv7NqcQgFfAA7H6rmMbetPANkC3rJHUZz1RHaXthqJtXfIjVs/G5qkfESBPCH3tQy5V2NC8
lZ2BOtoelnBYEm+czhcWtX5ReQnTw6SR4n0M1BA3E8C1fjcan6dKadX+rIeCA/2ce9KrZEZsvvZr
f3/KJ09o6DvZn4slbm1+yptclDYCGaVr86Znh4fTd1yyEk5LeJ2gLsbsP4Zr+voEgJU+Q5XnjdJn
nJpsd4NedXRnFV0+drhqnWo/MD9gAAJwK7kSiFUTTE1qfrUxoBWvVOMjm+wyGAhr/2Dcx49oG33G
cNHVuUyeH0HSAnAyiEpoT4lxk4GcXkU503xnXgwz/Me3+yfudX85Ad7v3H3A3d1XM0YxYvUwvo3C
r5FX91w9AtnaauU2BbEUOEbtQ1TzOPG7tjQC93ofFrwpLgtYaGw68fOjBqpZVK8gNkr3/dNoUOAp
RrDTXCFnHzo50txaZnii9vzCZJK0LpeG2KuwUdQsCydCXi5qZZ1r1zwXq/CkVYVw1/+Fgg7x5zL7
e7YLsg9Nxp638uPQUqDFG8RgAmt2OCVEP0Ja+ptPfcRpQuvp0djEQY+pwcne6XqcwsuzmdW+i/L5
o6urt3u4x6peLgU9wlratjaunQLkqvC86exUYLybw5XqSa6VViCfhP5i45bPrxI5ivM4srRqHIou
3v+687cgctFFQWUyvI/0XDCz7DHX8Xvva3NlYemEEvIQCfmxm1+yGpov02NRGZev+sDJBOVtb228
qXqI+vVa+i7EYIWR9z28U47zr05iavLjPAbGsLeW0YiwvQNQW0tUSxSjIAWkaHk/xU36FZbCqc4K
700YazIOPuA87k6CnMyAnDS5vaiibhPOLIwbPHBUU/1Dh6fM7Tsjf2kS0HISO1OUiisOItD+0jOn
6RDtEqXtdcrP7QMKfHGYhPG03Q51J0spAkPXeuNOZVollcu4agjMlGY2vSR6WRaEHrRvNNN8ot/Y
7fTZVWAqt/S/zR32aUdlKoD+42V8fwB9rc27+Mq5K4uZROrsTGSmIwdjJBHYzz1fGjMi4xzFGiWO
w+vDKp6slSuhsvftoMaVnxHtrh4qiwrxfgEdEivExU0HYB1f1lkNQpdg1DYmLReXSU+J30Iwz6l7
LuI+rkDOGMPtPWaCDOQcWDfI9cH5USb29AQSIcqy3PwZ5KDl3hXpcm+EqefFOQFPAlR5XPSjC+OB
YFsEsOzeQgQLdAPghJyAuQJGksrmTMtvvFqSSLo8NPIzGOAJhZ15JnhS3cwas7BuVs2gblutdu0U
fC5y5KPixNlJX1M6ZT2MB5mUn/QSaTL1T79n6edUFp3GeRFc6x5EkYdkfVl5Z0gK0RZw4ViSgypM
qiMOIkw9+L1i66ELX2Ye8LWXEkldenmaGr06rK0f4uAWD2WsQQx+mrMfrfeN5ubkg96fZL4iJ36W
zVfuFIRKJEnf7KNn4g/8cmwQMdPJJtFG9/gkxbP0B0PWoVPTCetvZnafyU9gnx9IOpjlx8Cfle6z
A+xzTm1Gh/7Dyx9MMFmGmWB1hlF1A0coHZsBPO0oTVvPCz7JQnCg4m7crdHicbMGlhk/jlvOrjM1
q140bBOc+or9/HefZNa+m74QsikVE4enuiMm/Dzlv0iLR3mvsRXuJpYbP9c0ruBWLlfJOK6kNsEd
OP0bwpaHa+T7JeKBiz52jk0Gnrem2rsXvW24NLDSyNZeiQqNoBmH4+9nrbTMKzMzmS59kT/bYnWt
kEBQ6Bxg5x/IOf920/LylJGpBiJDifoPXISMIeVqem9eY94syZYt20mLsBhaTn/Cfq+y9dq2y7j8
wvg5WutAn15voEx5ancb4Q+lEgaMY2VWeXzYtRUZY+mHG1Dv45Iro4Vu69QzLcK+pNGPp9d7urDk
+F9CYyd48C6LDLDHMfPvmx4ONLOrEQcaoRcm3HRyk5MycWfwucg2T6Dd2XoMIQSRl4Nx+ShyRCFS
xspDCiGaTdeTsdA0c8bvRiC7JfHCRXGmkmuNd7bS/b4+dWEGlnXTlcgRuFmv/8LIaUcLgR1VtZ4E
ieZsuUUjnOnwSFmc71alHPFgU6AQLkrTKgiedgYYwZ4FEufuxV3LZtCyVDAe8zxegBY+pHSJBxLu
N8S+B52U5Z5pt7yqUDzeKNYypov0GkFn0vsoSsKZKDikR3Z339WdU8jlJxYM8HsMocUUh+5TPDZ7
J7jIkNPcG/CLCsFr7KffmhdW9BgoLfxURFGJ/VygxK6kKFhk2Xh10vuPHfCnMSNN93Z4+FD/pevp
SfMpmVoMpGgA8zfx6Qd0NllDYGYqcl8XB+E5MU19LMrF3UPHXVKYGKL8jf7BgQ65hWk1VR4VYMWX
+5PKkvufSODhbpPonsWSODBeyU6gZqbwAQsr1a98tV51GYyNH6GM4piUOtTXnTT28cLONyqcs5jF
W4iVjqVxF7jdsBqYNF1D/z4uCOcrTZKdApV8jxoN+n8nmPvrnHTUbzagYsqa9r9+gd22IYxxEJGa
P2H1ev/zYJDCDJFGY5b5UzRDSr2VI3pYI4Mbosw+pyd8eFzoXpQaHvSt7EW7Z36FM43WCgffP2BT
xMRpnZIoRZzt+fF+ntUoMeqeO+/ZME0cbCPemHrIuBk9Cy/Ee5t9KvOsdYxZ0TBLuWji3s5G7aiX
qhpoTrtPhQNWS7yb8pVLNUV781qI8/+fRpID/NamH+QYWtbtmM4sLHoReomY/79lvbjf4fw+tgbY
F6StpaH/AH9/fW0YHAiyWVudnoQgkl++l7k35kgIYnOcOyEvSQO3TPKxeoCSo1xBeECKpd2zklAy
6etG8W/xlUbZX4M3xIVtLxYosIexloCWb+5J5KjTA26WztynSdIUXFZ5L1MTJ+hEgWlG1esWrnpF
yl4UaT8vNT3IDuwcWEy+EJxDJCEcvVS3BOv4kP8eZQ+rvoshBSKkS0cIp3nBbIbjmTjK9J2iOeAc
pg1eWcn81cV6C0WQyRw8KDYGASLab6JVlo0tAWi8l2orR0E54FwIi5HCO4E9rGKqTov2znvowE54
cmVcggcTNzROKlbRZrQW9bme23RZT17/sb4Ns6Vn1eBMSdoaB412GcJoDSiVS7ELg53+koVg1tRT
ydieEzd3voO5FyXMg/PCJr8mZd7ZGyfpGqcDTuoLmtKXxURvORrKTIaac7ir0yue8C16wMKFAhzP
Ip9z+ISA/nft+b1iGxpMN+R4DTzbGZA6Fl1fNLpxJFxsNUrem7uZCrA9D5IWLX0sQfvzYPHOPU4P
JSvA5oatXwvet5ua+N1JT2TP7T7LZWwlboMU8/MkH7bdxpWfAZi/EoP3By6qDOHVUqYEpz6ayO7/
u+NmoGxzvqoL9r4KTXAWWqDFM79H4tlGAdPK+F5kzXBpN2NDxxYr8X7wEPDZ9VJUhLTHnVSP1Tzb
OSISagmAX6bgQqmlgKR+L5xM2816aqYR5q22ctmBQmeUHBtPNCh8zt2wpPc2unrxUbmhbCssl1gx
9l98YZseAYumLtqi+iYpO4MMCDComjCCcrq0Tg10Le7c2TuBlCBDzHX80nqgncKPGOHc47K68+7j
5jbYhrS/akWrDlJ3auldwYGFsczo4384i7anA7SwMYVlpn/RYuRhz4QKUF2Ge2kSolfjlBS3rqU4
INOpurAzO/dZloJr0YMwxOFcfZso5zxDVYsDgfxNyUGiTxJEW/8iWa5b6sF57csiGHdPSLbEti3q
MT6QZlpSXsc2ecQNguaIHZPDRTmaPwW7awIV8W3cEnjYvfuBT3M8dj9g8lfemFT8CS3WMf0192Fq
EaalXxw7WGqgu0YY1W4Sz4pi1c2q2h7QrqY7YhvndMvSnpeB+58d/xWeqf+BxnG16e1ECYZ+oZBZ
fLoC64Dz/87EPpzCFF5nwPBKJNl8AYJzvYXnP2RKGfpUUM5duKxCg76Swg5BGrDY4uPpaN/6o5vw
DLheZu8WE9jRQZlOx1ZfehKqHXSn8bag7Uur3tO/2XxDWP4fb5YFpaM8VWSaTy/f+950w73LBuF1
VvU64ZfPt/V+5m66oHtGEribPWe9r5tahMdAWAe/7oG/PP8YdX6MVQWNxQZ5yikAJ0KpWdChXSKp
KEa4IAsHkMsneYfEzOZC+JFMLzWnvQ0AiAN9l2aKaYSz9ZEDhCICgw7yFhcs4OHpjHHxRvGV/Q8r
1eiiZqMlnrLkC8CMcj7/Sqsf19BG8baQwuzBu5DTbW1h8GvDPcUKuOa3vLJ8YPO1WL+1Fs/WQNXZ
MwTy4tZeLN+1oe6AEfnUijpdUG5dggakL1NcsJZPhFJJGs7AZO/tXfbSDoMNmRYclLu9ABUn5OaC
tubjFBCbk+/F73+Uk2wOZnJtI8kdw5dCKSUgfp1qT77pVy/ZoYR065v47gkafd+GiIyArO9bPiw3
/9O44vHzC9vQZLLnqUo9d1fgF8xbvJV/hhUGGF1sapi2D8rOsLBydjMr1/wXQx1UOs6kaSRjrLoW
p3mfxvUtw+bITQ4JYG8e+eYgEyxnE6Oiqdn6L+0OlKmlA/QzcFxFTpH1SEJxPkThGM+WPT9Rn2Pu
5/hbb4yAhSrTDdfKeRkyRPoTrEchDkiDMMEAgheQrzvpHGzRYh9XiCJTNq19ZZRzWGBuD0fJta4w
MLz//ZLMl/pMEhdklu0sQD8tqU2dWAM4nGlPypKqxXVSJdIdz3lxZuw65t1Bar60dwpEhGovOWl9
1hlxSHhslpmRGaAi5kcdxPjq94pXJuaJ/yMPXbjYY/UuIwckFh/XaVlLHyiW75b//gkNOgI4ii6F
gH4OkmnaRyf8OGS0cuIEWn5/MIaOIm6IvzTFLSXub4gY98g0h3zN6IY8wAPjeHURwq04b4B1NBmb
NNlsA1juu5NLfuzyg01HGpQnPhUxzt/u6mFVyCLo26kgEH9n+wC5K39BfkCZHSVNmroAmg1TeTVV
P20Fi7B2fNq7nWkJ2Ca3GYF9fj6h2EdMcWEHh1J39Yi7c7mokMwqzXp+BFhTqf3rqHjb80V/3WIM
HdBvlhW6UJv88qSNVsDNY7Bu+vjTIJecs3w8TMZmFQHno7+Jo5AgSOUlzNkzbj1LPMr8JPMPaKeR
OSEiBkhO8S38zoDDLTh6e61Rt4XJAXI75wEKL0vMXiL+jePhBtmLV7XVEQO/UQ5zu+JVFXIC+9wQ
yoZay8z0/6w5ZGstf9jUAbRHhLHGr6xcbbr4vEHIZX5BkBb8IH2LOmCoxmHWySdz7w0R69jDtMop
GJmQ2gJRTGYUj4Z6Q0C0ckiatP0rOcYxGUCEJ/pbgYC3G7umYqUFZOk0ymQ2ckh0S9lEROzsaHiP
Nx+FwrlHpsKKu/L8WRWAsI9Hz8mLER1iy3rKW0NcQT1ihMzvLNiGtr35o5IwnDDpTQsBp3DbKzze
E5BBZSUoNv/xTZ8swBDLwpZXaoZLLxdoVA9Q4vFtO9pWcSWgTjMQL2yJo01mbRYCFuhM8FmzJydt
lS+XOvNu5KU1A2DwUihie8Shx0A74YGKGtznCmC/mbtcwhglLotXFODdOYlKMG048XUMuLeAxqnm
F0T2O1hEas3HRi35TlphYFAXE70jghHVnWB69Hen3VnXVk1Lbi3xjAzrnyWD9ypHGQAvdCMynL9H
F/Ds20nVf2rWC+loTyLgoWdoZLb1nmG6FXaKUbCiG8zujxA9wHtF2gi3dZz0PWBc9erZab4ITWFr
iIwA7+C6Sw8I9l8GQfcL1gBeibNzapl2Ij2DW9GQZ6im/B2HCqb+HikzqSIb13xyaqPL/ecZX+Wn
bSmKBCGKXgaKizPzIUQFGYP/zemobi30HgdbBCdAYk3ZcmEdifbX2VV3FFU/aqBH/kTn0FKYqeU2
2YxPIweAQCsknKry94QeKjBQTth6updqqZimwAagFwVqvvK4omF9OBtsNc3ZWyCZI/eqAC0k0G/M
+YtoUMxRK1V3/QRyo1S3IMbqJR05UIIcW/mLPZ97XV778+rsMtPspfCpNrWT+ZjhSMQGQcOhxivh
qd7lP/PQjkg5pbyd1Sf9+mu8xDy2EdDyBcIh0NIr5PWyUwg1M5dUQZHGjWhwJfwQFKQVpuX7YZCT
/6KjP0Mn1W6FbG97eUNDvcm0XNBUEyq8y0SJBdsXkjzZOjRDajmpGcsQqSj3P4w/1ZaRvi+NqUfu
9hRh/PEJTRWqk72wf6uZV/zHX+85ZETdINyrcZFlDmjfTcTG8WeIWWMgPW3Rn63IY7A5esWeBsvj
wtSMmA+NWj3q+QwFrvtBO2+sQfrUJHRsDRrFNipU4bS+Z87pvbO4/2hmCbjYnlWccOoRUmo6IcRb
qIWi5AFGMPDu8kgFyC0gtFw20rEXdPRbQarpC79QBAcRAaib3ngMPRII41gtOhgBReTUVzrxEddA
xO8dT+B5SoU7ugQBW1NWJY4LrXhtU+PmjbYEJi5+c7v5/Quw9ZMvFrv6GxNWO2qZrwfNBcxeCUAx
9nDEGHAxgf33e+zjkn5mxkYJ5UQb75hXfnbxig98MXcheFYwviaMWpvXn7WGwmJ4HLXKtK6OcK8t
f2/il71AcNuPZNUCuHN+kXHiyx0nYrMioCavm8MX4aQsDfTdBCOLqx/WKgphtZTnsM7etQS40dkg
utNrmhOWyWLI8xecwgjFXf5KUNpoSt9nLifECmaGSj0cGn9HRH1nhncE+gpU7LVuRDF/0fzHstN3
yOE2keyfINYspaJyKoAGWRfeCKPVjrM5OnhEFptZQ4HYoKDknaIr8SzUPM5i4HUTEGXl7HDUrbgn
pfQRlF+p71YlCcr+owV/imTQsE3IcBSnUbcAdYpjnO9TjI8hZcUso+E8gqAuZka2N9ilu8jKiGu6
wr9n8M7yiQCuBcSijmXp0Tq6nXXQgbwYbP5bqu1r9yVOneQlYRbcwClr97/bmrnBIt2K3yTFn/fZ
yxzASOD+zsJzMhMCd76RozmwwVGj7IsZ40icN7oGJdpKtUpvfTRH0fZXkb8WPDR8vDOo4JHhNx0i
yc4fBnkWqnH6sCDAisR878SzdjBiuV+HH2fxxFdf4cAeovO7VKJ7ZIJIKxqHW4VTvPvr8+QuGciV
29RXHDa+rIQ59UJr1N5xy5DrXm7nCaB33D1BrgrWvlRhOCn45nirC3r0lWbpCb6kd79/I5hoyS33
BTS5l2aa57ElR8Lh6IrADhiBLp7XcJk0Nr4ZZhyrhi27zQHCSNKtulKoZKbkgo/t1ZH5KWNqJ2I6
4btZgH53a/oRk4Wiy2tXeH8Zbq7SzzHJ8gWsan77oGEcdhK92lHr0VvJ3Qe/lg75EXQu5M4+6V8B
EaJMCh/CAa+bRyFezoMk6IkeIRATwgvIbaSRD6oliXxyybFEsOwRbR9ni9qvyib8yO3xvbETJkt/
dPSUq1mBKNPfwwHvET5yKnLp3azE8Oj9AP0FLI6ofHjrED85ZczBHFftJYn0if3PhiY4qtcudN/4
SjP7zRLnE4qw8fvpa/Ayb8lCBYq1F09SnfU/clspuI0O+keJdXu0etRwzuXvhS8+Xs4xCMMsHn4B
bnqSlmTcd75Z3M3agzac218LlmoM+mq/3TonOCcvWx3ehg2Krb171eTpvqyj358HZTMwFFf7KuKx
3WO/fd3v/pfgx58eljptqyLV6d1ObJs4xnDCMZgXCIHSReDqyaEbN+8UEsocozjtbFcPJknO0WD6
GQ6skP7RP/azxnLpX7M9d9nX/eFTLw5zTnw1MyeaCaNU365A7WcBd2InWv9O2amVx9JP96Jg83ZP
XwK4GRdAn/dCKv/FE9VvKfm98CBuAtYKfkjBxbN4+MjcVNZiCgK1sxLwrAz/KHoCbY+edujx8MZO
N6Td2UKD6sBbL3olhWsLLu+dNTPYcuGDmXvAxFKupBHBKQFW4PqnuNnQvlKuKIqmWfIbfy3cGX66
63knHqrv0UgOlh4IgjETwWIOcL4xIXZaTyyVq6iRhYoTTs1DHtP5VKqtYpF92GD5g/o1imDEDWWR
dv69wTlIjbzrAa/1f6AaSX0WLrTvtMQe+OT6nukS/ebAndsUIWVAHBrCaVqyCnpgEJojNfuNX8Vv
XoIZkzWOvosQAdts+VFEVCd/NHCJIUakOBSVm9txxvM3U75S5uPNtvtUx3JANxv4M4x48iyteRM7
PLvFkHtGB6ftsQK8ShqzA1E/0TQNGWRpkIJoRFcXnXxKrTsFdDUc3Nfid+s0ssyiybQJvEqZbHAq
VjhJHvBwkIsRDwyI/+1s8je/m0Fcn2ThvohquSO2dsyxD7laH8+U/8Eq06Oq0Iu5X6704pMH5uSx
quzFhbxTuSaLO1sXUPAv/anMiypi4U8VW8Wnb4n02Rfy04nEAZ30KvpUeS9RV4ojXAoYrBPVW1Cc
c2H4zRCErhE7dPK1MB7Xjk/+tew647nDtm2b8wv7xfNvcv6p0x5PoU0S2W8xyydSPUnOl9OA+56S
fldaDPKkGxy8WEfbw4VLbS+f2oQ6CUJSC33ag/Asg3FPXCb6BWBs8G1+9y7UHwDha58Bn80Vmk9U
XTEXlnEZZoxqSnoKL1rQMd3Wnetmi2s4si1Iml+dcGW7fbn1BgMradMzoqf00smQmt4U6HRQCAt2
E5+mj7KRo4j1PRO4C/4mbIvECDMddWLUOnthQ9NesblKQvqQ0HQQdJY5IWALuxNBZaIkNMcMX7pe
S74WxBLLuMMSggMgM0J9HNUZPzkL3UGPBOhoNBF/hzGw/yZp7OLNglLsuUR63yUO6DxZboLkCcFf
mmxYHPnkJh8jmtUdTTK5pne4c/NXoGxqsD4MaiAoTYegYS85gfHfB+thbpWoqd7OonC3GprtwFeE
6Seaz4Ln72BQ+NvpE1Po+lkPuJLVc3peF+DDFAsg3Ff8OmonUVzqEnRgQFr1xxUSr0U3zWh1tZKn
zfA3Yt9rOvud4fg3hDeHD1TjOTZ3b5dftDEKD3q7kRSiScXmywCeyIwTvKWf6i5N3C+3iQyFBWqm
GurwXujYLfwmOOXw/3D8keHPODzvEriclhyk19EI2DxJRAqA9TWNZn8UgXOS0AQmQZsSXYRu5Tmq
OxBzbaFeAUGxOdODyZ29ucU/fcYxqZGFvNQMhAlpBL0hkr3qN43Marsw/aU2nLdW4eY4BQP09UpK
rmdwForFujIwf5WSdwG8tfk0higAk5NJ4TY6F/MmW9ipvGr/Vny0/iS4D6o9IpDwCUFg8mYeXQNk
6vzyxqaJ4l4tlPSTWisSBaWWeM45ul/bU5dgNgzeMI7M6gcgi7tfAouBE8Nei+sQmna1Cp+1AlV8
sgYcTt4Pcah3JnuN3Pr0a1x/R3gzbCPgCkIHU2TpydAl5oGChX2xZgE2lkaW9KJfRNxvooudKB8Y
u9+TBMYURyJ28Qn3kft5o2pHbA4KQE6cXQutv3IVeMFA6XFN6hlt725whE1spAOEi8dSNrCZ2qt8
h11hOIefue4wGrv/+Qm2O4qRu+xlHhs+0zAu9mJKmT6TgHsjidu/LD3iI3qTNOOMivdsHbiguG6B
12rJa09cCcOkhSKz1yhYZbI+k0hjaFYoFwQn/qHADQAS4gSnXdZDfjNPlWb02gCmtWPFZVeT3Dww
AWPkaD9jfXVY3JxBOQPJki7gaKit4vReskWK9M9m+0gwotJb/fJvyhUuW0R7Hp1kQ7jYf/AhJCgi
ByEUJNGWsAWi7r6QylYgbKzK5TEuFS0ZKwRXrzcbMNu55pe32+FXDil6FjsAUd2tHmppOl8MmGoZ
g9NuMEXwxdsYc7aOIQ6/mWpSLHASruwtJD8c3fqGI12oK3cnpw/OSvRP/Jh6/FwIQ7lRCEdb/v3s
6SbSbHZyFgY3Fxk01jpz0DepoYLyLshcpQPEmQeVGT/V43XxCh/5N2J3+3PPxOP/fh0zWKCB+m+0
hMkXjJWcEvAoA4VaGnibUqnWig+6/IxQHmXWKNsf9sWOMjEE5YY/k3XCG6fP918D60ez5r5ffYl2
0D3b+yv5znycYxegM8dbklTZLbH6z9MYQNK85fqjWKsGkQnM/o5LMj92NbWZvsU+2vDYuBkZ/dp0
0gYbLc63w01A9gBZhxBv5Yws79FzQZeL/+jr3qUfL9TN1JsTgI9x89zp6MoXX8tbbtfBf00VGpRg
mYpUhn3TjLt2unK2wyNsNk9aEUW6NOdpbBbwRvaZhg60s/GxBOnOcldFtuxpc8fPvBaNtzKy4Dx/
rALns00xmUny4SobQFjl+WgKbu46M6JkTu97hjx0MY6ILnZ3uTaObrUpI1Fr/RUTHfOhGVTsTALO
ML/ZkdQpLFjxxynWtYxaldV/k2tUfqCfj9vlnCuWVfaeSaXb2Ch5s1ssmEeNgKEnpE8AocNji2iV
hUVuIOf0+A+mLnxci+RjRgxTL9DIBLf9oWzLlc85dhrF8ND2d231KS5OI7JMpAdU58G6CoCZ0T8H
gbH4mdiIHUULZfTZ1lzxllsx79scngS0Ku+QkEfBlrDWLwlXS+pxUqU5SuPZW+By/9X+SBCZsvgM
+xhdyMQZN032RAJGqNn6zrtyz9p3kwB5+XTPx7u4y6mIGt+AMMlXsGS7pnuFvNbNo/KVkziE1Do2
pM4B3KPUK+ljuIOW/i+ivQpQrlcSPelxkZ5gjvTIio2qEV7Pgpp/npDcCbMuF9ZR91I1nBggF3FQ
pFooCydS5U9eVDtrqDf5f/ywa+6I4Uk8pC4D/sHub3yR0yRIzioZZgGU7EFCyZhLJzt3OFaCv3go
YhnsIDeX+/89EqQ7Ji6OMrJFgtXFzcxv3StFfqjloVJ3oqKR+LZJMu2YCsqD12kkZxs1HVftFBqd
Wd7yEgyn1asT1qZxL8fxZFgI8nIA32MAhjmwInPKKwbP15CeLh/hEo5ljNn7E0ub5x0yBEgpN/Yc
PBnxpyqXi9KL9LAp8Mpo2RjGROAIrRnxBAbBNtX0bWCzymoyAEWS0MSfG7s75747aiVTM3QgwIx1
/5xq+nWnk3nbLvLQHfusOzq+2KD/lvyYyCNbr9QFyXZ/rkEMgo5Iit8neh7tJPeKBu5mCxwQNQxw
6aPX6Jwr4dmxq/ZwJ1ckLg4H6E4ORDuF7PINZxornV7RBIqdaoVFQrUHCW0yWqUicRRGHQlh2N+t
pGAJ7IGKGOGjlvNXhW9xeoh+SeBlIRKmGsaU2YyrRzpJEi4E9wfIJZJWSYgg/FlgEo5zziGZF/2y
UzM1m+2lId5b5uc3lufUdDJ7JT2RwX2shGAiKHp2SNC1k6bGfU+ycIF7GQSuB7C1+OPTonn1i89q
vyk2MA/XWbm9K3l4rNH2+7ND9Y5J4hySbRdjct8kdB6p51W5bQKm9+MzrB957G6dsD8rMRoaBmq2
9dI3tALDV98kTr3Z5Pw9Cg7HLjEbeQ3/f9rkVj804hhHikB0OsbcmaAppzGdegb++g+i+5Ea8rdR
dKpoPvdgzjGxKy6vlqFa9ap0vBMywmrYtisG8xmk5hbFUFoLblInl9/hKWBDwPqicVE9pkOMgO0a
dkoHm9dDX+MS+rk2yKKZMc8eliQ6y/+TnoXWfjrwaCbSGl/aDRHMvaNPNbZSmg5BlAr1k8wvgis3
ojDd0VUhSGoptIAmTwq8OiEJ5TC6pEEMfk9iYumbe8ftJz5LGwP4ARwKumWGq8ec1ssYzddbJ9ze
W2mLWvHzrmD7B4uTezo+tkVo5mFQhm8NCLcwK40SSPMnprhZB+Aw2M/k7KPwPJUPh596GoREdgUq
QvvVxDzdpz8oZBOYJ2nXN8Htig9AsBolQ4Sp0lyhhdq/1smAiwScWOzRDMy/0/ifdv6Oytf/mV/e
xCP0eSwKBWgnCQ0TolKGYnN/hWSBRFw+AbIZrHA6CyEbnKLrHZLMVZGksNomt8ixcbTrskYu4Xk2
JVUkxIAlklBRUAc4MfqxO/FvFnrfQF7oeGHqN8G1MSVwPR5y4OD0BT7Smosv1nPbO88REGacfxF0
AXJxxX43R4wwHGUOZleWBz/RAabtnZ1BFXUTX4wLObOVMRP08+GfPN6EVMGRcJnQDuWTQqQktC72
gkB6TURkS3gcrihmxIJkNIT8ym80BSKu2epqmLlTOD9itY+1SeoV8PyWnHhe0KTwPg328Ry0u5sS
ruKwu0/sZ45GGu9QT1yu1nH6K6mAbS4vYMWFudAsVsDJz/FROZzDpKBC66aTw+iD6TGRw3jZBPBJ
RW0k4NX95JMoV6BvINLQ1j62cX7P3LUFcMRsQRCu9PN/U6C/NcOW8AoXM4ik1jeLvXUe9IEbmKTw
W2b1D2C5qv4QZq/cUIzFAP32kEWDa0oEuVWYpkVVsNmQHfmIpekmnuhSUrFgRXSWnkGG2XxB3gcc
3Etyw0/wmGPDoSkrtvW2m2NOYCLZ73PviP+OQXYvCWhzd3Lj+WYr/jv2n2VPLJGhhrVADgZow8/r
NR2ROEBbdvc84T+b5Jg1sKt390QKQLsbzLdFV43amFalUWl4u5/4CkXu5PiaoYrAIJ1tFOsC68LC
jZdODPl9iOtdIjmqfSmPpHgPty5tbZ6l+ckjJXOaXAYFkrtBr067xyFp7cFUj4GFeOqv18ct0980
EDWWLAV6uieynWZd/kzKA6MzJClvyl+e0yIh6v4qagQAe6wokckH3euK1ISvLJbuM43mHdeMEzWT
b4acXy3so78DV87qD4EONTzUYYRT3aYa++hXM/T5TQBL7f9y9o9g2f+Y+qfdRtyWp/KkiWdbmUmP
ZI/OfsKftzhgDdk2uwt0ezpzn/Hpq2EXkVsHg5jU3nptOxT7H747krNjxcS1rgCVWjairHIyzTTc
8Za8np1rZQMynJjLlex32IV3pHnWaBY8XNNpqhFqta97bx55ClX95bWgbtkLmNMP2KZjy8TzNU4W
xpQNcrtsjl1P5am/fX4BmxuRP7vA/2Dz01XIIa2Hvx6CHMLe8GiNbKMOgJVsi6/2vbVgg8s1NQfl
0A8V0F2qs/nX45S9wQZr2rvsqIC1xlKh3NjgdQEt0gi5/bwvcCINE5Zx5UZZb988XgqY3zuaIYah
gWu7H0zFvaLZ/zA/nDYeLf7gOhceWfQKN/RsMV4PJyft7x7Sc0YAC5EM+m++Qh9+9Xqq+9HcHTXa
X93/UyEXtge89zuE40Xi/D7Hr9McAdMY1cd7VbhObrudk5VqSnoDBvEyh/LCnpWbhq9Ou183HMbJ
OkqfidvDgGsXOV2nmRyXQmM0JDFEij1GbaiSG6P4ri25Bgzzr7Cq+RRrDzj2yaQwc3w1NQJg5S79
pVAxbKAT90orLp6B+hWzy8DddTu33hVG89MplAGM4gHJYt7wZiRfNWfnhZRNEhjXvCoB9S6q+QRo
rsRYB01EWDc8QrprddznEptXEgfZssQh2ouydAx+9ZrYK6XW6RtrV5wJU8xcEp7/03S9KFkXxuof
cUCsAzimRaic6En4YWKKHJyQGFX4JwqAFpYnJ/eNR1oHPreC6ncpY6sXvPxWQNEtbsIuwPpFl29p
eSDIMFVUQsKIBlB3QUPXS0zRAxsDemWkPdSemgGs58/39t2Hsbx0RQGI3641hJdxEVjP3snbzI+f
pJIVt7jFoHGAQ7tWQYge3heBskghEqlmYk245wrIy5f7C/2vePOMicygq8KK1hnHmcrGR0CIL7gy
L2nqcVrZMY2Xu0w2jj5CMa6djhyHmY+XH1jVl8ZRvKENUvzUzRXDs7nm2H855dL15NVRPQSJxFa8
thImc8XhQ6LNahKB3CADj0nVPXMeDITBFHI8qTd+hndorugCXrAsdOJZuuVEr4Gc14bvB7S3CcX1
q+L4//ZD5IRIdJuAB3uq/Aj/RfPvWbWcVqcY719xNbjxlr6ccLIH1Tl/a6gK/5S+i/GJRUC2SOmF
I9zp+3RiO9+gfmSSLc5HOQvTe98SNTMBKHkT//glkDHef9jAHB+Q1wAJZE6RChaGEuYwzTChjAhF
NqMbkJZQwVqbYS5OvDjutAc8ay4zIHYLsQSFN4WyDrFfspEwV0GWpS96qlTgER0458vnshus7+98
FMyqovJWWt0eDxMvP0tJGaBQR71i8uU0YFatClzsf6vr2/kFK/c3LeDvikeddWq56LuXvZYrWctN
v8h+9c7d7Ka/tTdvz4InLsDUv3mXONiPOcgynIXNQ6aXYHlsW1iNqlMmUP6QYw9biCtagccklCfY
PUCihaI471Jibe5b2vuK2yPViiNCaDiXMGz1CLvDxSdSZx9eBnwNY7OskmIpEDfaDyKV6iAF9fUx
3aYH15NOYLe2C2YUbBxyyE7tmdNoPq8bsNSdKYsZrYN/Exfb6KCz6cmzvytZC2CzjUKxZqTSCSVS
43QoXy/O/6rX09LrnKFLZxmKcaK/q88Zjr6LRXFQi4rdusjjC/2OfzJwk/CXy/McBOmiA91w91Ci
C6PQf15BOm6Dr6qaR/Kbo+Hh7uTNPWRaJdyjio7tU66gCiUOqBbSeEmf8rGYdUV/HI+BvOp7xs9e
VnzhI0sNwkJHCZR5FB5sMANxAaVlZX7PAi4s2/46psztLVey9VSWtK+jcQlXqiIe+4PG1sdqWv45
h4FQGBD9/vnAujaCusrw/IOaubOUdMI7W90rnFc2V1yDGAGXxoUu8Msz5uohZy3WrvYOWN2O2yb1
MUm9knxLmxngQxtGUd+6p8Wibo1QMDzM6noO3ENaDGrmoa4q5QNUtVA4/TKp2dxSEbCA1/gPBIgt
T4ijFmIcboOou2iGgpPPrvkDpW4o+1EqOOEawo5JQd1dySTIhVeDLwHkKYDC2O7U1S0/u3LtgCr1
gcuz/PfPQ8Inh6mVSEd2xg30q7AMoiNPw6ZLC4a24F/7l40vtIsabqbU0Bq5xqcgAScNLM8p301j
Gj2lKCMHdQxxnib+7Bx7oDyNIz9S/6hGcBIFCcO/p2RRFZ9i1vqy0YT/N5HWu0ZzK+9IgL7vol2P
8jhnwSEoNNX7cVQ2JgpCLoBs8wCoY0800iRZcgf0QibYa8PG5UXirX1WG1LrFGFNnKQevhl26BQR
oP1qq5Ut7H/XeTTbM5RE7nhFhDg+Uj9Z3lpz3uT4WJ0DSijnB1deOiBEfHrPf7AQjyDuIe3T/hRL
bbtJXCGu2tibAd/j/Lfd2SRAmQy0t3qaJsbhuTxGCjbCxvakv+e5FcmB0c2Pwv6Cebpm2qxUaibw
azYQnwF0dWk8wEFhN/x70VLUVtyRUQGOnzV9Kv7gXvF4EA+O5+LYjRVEI2cQMYO+5XmXCyqw4ZIf
2pJGSn8kEf8uIYoHchXlMTXLosPz7KxfShu8AM4sZ3ekRQshoPC+r2eRcUwj9cEhU2q/f5MFyp9G
0qLEod3Vl8GusRS689F8L/ttKXpvU34mwObsUKDhyyuZFYeFnlQC9xBe+KXu818OIWi/Op6GuMNJ
EaTtI3QncN2YoPcv7OtwRc/nQkeQF1FfY9c/XbH4kqHhoThbjV4aBSwGB6C46KhIjTZtYDiQz47N
PuKjzJT1TJzHrqHw8/DWOvllmD99b3E/rp6WyFiamhip7cJINy1V+4dwgObMUP4sZVAJmJD0+upA
35UAL8WOnpAANS0icQox4VV5HpJ4sd4oxfu+YhcscU5CQHDM5Gfo9/6eeflHXBETZqkdpSQLReLh
N1z4hlGJ9B8e1jV1oiv6EvW9itaOqjyLiMfwqnu6n8Z0cC11CUOERyRD4eyZewa+fFPQLQfgnazq
yIWsYk1ih1n3qlUdnEHEy/9bVv61gsOcwzGRb4P7A1BToiJspQBTo4B0csdJkh5ES8QyYR8a7zr9
E16eEbfOqWfJ7Org8Nc6qsZXeUPBdxEFJ6iko3MPYrgl9DhFg9MSzNWQE4SmLtdDEt97qIrC2l2W
kvpmGoRSne5wUioItC1w7z9jTqM+yyE+G5gNuZFiP2mMW3pfUZsUsVZYZ7vTjNLQeQlKxRfsOMp1
UXVwmOcPadgCtXxXjaZM9EJEWJSCYJnf57sjvw2WjggOrmPAgdt+7ICka2Nr+SuQS0JDz47HYl5l
4MVTZoNh/D78aJ0ftjPCE0IwDbUr6rc5VT2XDrdpoernbMfQ3yAuuRyX3yRfC5vzNPkSlF4oTSyh
1jJRgSnDoJYf/oHPsULows9qq74eLwLRlfjk7LV7mfsMdypv1t/i2i43iGqqK/8/U8scwtK3BXB9
VRPPe+FDaJaV4X3IfLPeHeiddu6Mtk7CODHTdNhuVX3lcE/LoyIT8XRKC0+5jgZogcW/sZ70uzVf
rkOVPcpsC8w/9FhyWyPeerbbqvN/vvCAnISOcMm3QOxiQRsLkxUeqPxH/uFwcm8WMFhgZDO+MUI+
3yRp2mb5i6+bBQfBsFc67AbZgrYLg+N/KGOoq98opb7qBP+N7aMxwRpq9NClPdYDMy2PuGL1d0ty
b1mZIGhiUV7xmVu0R7wTNZ4bGcKJwNAmOoJmuUBy8+4LtU7g0sMFOHhsFwsTDAlJEMZIwtOt2Ql5
eI258aaY+tUyVFzc6ZdIaaNMGQ1LC02Jmro5JpK5tyGcOMagkKSYxbyszIVK+hDKEs7kbuxGu5sF
HcqTGEvmGy669ZotPhvEeBKPdvTIZs2i+d2QPbX+EdMaZMBojoW9gmdUbZAz5OfjvZCLByIRFPQW
zgCOqm/P+Y5xa85pFMfNHImjMp840vksTI0CC9bDSB4s2P/5wwIZEPA2ahiQObS5fdEOSWzQTxbl
ggqNS4vgXmQheuN3dpN5eaGtqst+hs+bb20llKRdYUmp0Y9/ekh3DH8PbHQydrjnZ7L/z9GAI73g
ikARYj8X6UgLksNu5f2WmkqbaGsA3yW5py07t34NvgIbY8p+ZVryS0B7R3OWMpNqDmufEptNqgow
T4DC5dgtrXmJfkGZDe3sAkRuqZo3D85cbsXF8ODAE6RJNZuCpV/9lBypDOOOvGat0SfWsHDF4Oq2
XSJfnjZnkDvIP+MRQ03nso/InCcSC2J/noOck4MB9viUR6tfiByR1rAmmAgnovHJ614qa53Xc4kD
W7c7VHz+9QnvYyvEyRpjiMiz5N59BNsDLijSvYmcV9pO8qLY3AOOZweGOCx1XkExgLRj/SjLC+y6
coBwyMqAoSh32OgqRhWPBmJ6XK3HiPlbPo0eekrlN910ga4r4eJ+bO0xam5k9d9+2vXEcwxGg/Ed
dFvHHREoVjDYGZHpzIikq02azHkcmSiEJj8CZIc3L7rvfdBnE2pDTUopTMytt1b1gCJ2i9ei9/xq
u80t56akK2ziTaUFhbwWrF/6ltz58l/DaXcbeiXm1waqG4cQQAROASUHoZQqh2m0qnhcxbhDY8tF
sNCU9OiWVX/t1EynvwGC/f9z2pmsBFsLIDwvT3lbcQFHAv5uGT8QKJuvj/BuO55zeDCiU9qphSW4
v8HqehBh6WVSEK10+3O41mlLUyM289ilqryeVlQpW4k5tATQtWXzoZatToFydiOjaYJx3lDJw3F7
T9A0OELspUT4b86z2nTh+3KrdhJNJM/NFz1M3pecoFOrzHaoJ23IoMOSNfUjaqiYzt7wP8gD+rWP
4rhqSujn01ODlkFbogMS5zv7MUTV1JqWw9jMQT4DNulWVJTLn21lOojZ+ag3koNPncmsme52Rakx
7lOefd5kL04w1RCpvSK32fwGCYVKFMI3xUNEuMSPi4KS8ZMZt/tj9Bo8B4I8v11VNuj/VXzL8k2u
jNPlWZtjkHilbuJjYwZQP2JDM8IeftSkh+sLOLlw0EmyoFFG9Y9tEchKxJoAmzAHUYZ/VqTnEKHw
1lHgRC2at43LWlmMCfKZXp8WOw7Oabaf8haKYOc6w2YyhKqkeTxrpf7btgUuqWepaFeXk9lq+oKM
kmJ7IrJ742KoAEFvQYEEd6h5hlGkIN9/bnXgjjpCIB8n9woZJEVfYec8IH9psJuNa9QUyn5T/2ml
8pAyfyP/2q2/+KlxcUykUcMIaxexx3Uxzr3yMLMfuOeN1xTL4gEBAoKq/3Sgybdr/VKqXG+78Wpt
K8utAbkjTeDAgYNRiCsYKs0qx8qYBcjaub2EZzZMcYctiSQ8zO4n4nL2DNHQ2dYFuwoybKa+rm2I
vj5eIT/n7G/Szgrya3eH1ka0TdSgy2Y8TimJ7FqsRJMPQ01knGrVDgVit89ckxCIlL+/bmr062zW
OIpjdUkXHM+q5m8t9S5Y2WuBce5ObYCPJXRumpmFx5Kw4gaUFcYoTwBJ7hPGf5sF1Vu6W0LCPiFe
l0Bqc+jPEnU8VbQeVMhszlIt8e8MVeTjAmoKmr/YsR6m4SZkzSvywYkHGVpwLvDuTN8CewWHRoOU
cq88p2qI5IXXD0X40dkZFWr8trgoS4s/36oxzTBwUsuejgsCYOtPYhJzZO88iOiKHI4I71QD4fCh
d+f4oaGxBhkNkAoT43oz5Zd+hfm2eUI1ZxuZ567sGHHVllElvU121MichDKuoUOCTIsM4ow3Kqc+
futgEaAg/GXpNuJHdiiPv5PczfjRnnwwg57KthsOQmXnZkbIHT+OjU+Gt6+2eOKewcJ6OE+6TL8X
6I5gL5EKmTlE9ydCOq932ynYukORM2Ev5IbzhjHOuX5HuNhoDPV5guzVTqim4l9w1ruHO5Poqq6r
sGokDxLWwNVsK2KEpOvEt4XmCQN712/MXcHnOjcBmBUUbv8FWS3lGVG7sjyn5JukGG1Vq8RZ+Xhp
SvD+V4S0SN+/YnGRE3NlwHjWFaNg81WziM01gA5ddCTnxso2n/1d/5oAYwGZNO2/ALhFGmjaouT1
I0lNOLKeTlLFXdOG+dctYUpwM9za6cXn25U/1nW2BpTef1uqAHE6hSO/nRTCrkl39MYZM7MCCcO2
+9begZ1MLVVVObtW3FSRRcWVUUr9Alt4CwxWSibXJKbxJvqII+tl6oIXPqbRsFrFu7HNI8eEtVMW
1gb9UNYPeUea7Rn6rHsZZmPpKV8vCrFnssRjBnD6+UCkYBVKjg42qMN1e9YsA9kgBjd9p/WQMl4F
4Ho7Qwj6y/3eilZxOVZTiYtSEbpHV2f/W0B1SPzCFVafshMeSEvABb3qEFZaZfPE7ueVpZHyiVcJ
zuJA6bDh0A9CBYqSUk9ExnZ+/faQI/0t6dvNd1bBjzYMJbEe2O8WzTtp8N5JHcKRo//AevxhITVM
2JCsOHbyU/eO10aliNFp3bAHxJOmNznyeL/8SOcMFuCbnbu3CLBW/4iGTkoqHeWURQ0jTjWHHsRH
/zY7WBq6d356jRHG1iL7Zt624nGNDIdDylyogJMGWDPFWZLDamDnUlD6NwVh16eJGGQnYq+NyPFt
1oXleEzmXIZTgXD0B2er7YdJO3yHrUllD/nWfuQ3JLl+a91WNeEhHIUUeh1LSBrmRtbacaQsn8YL
FSHJZ8uKpoPyyIemTKVkxWQCO/bxKljGz0qYGqbfIkqmMEYfuBElL8YPQzXYwxv2ToH/0uIjPJre
/2mOJQ3LhjmFE32iIRJ1FEyU3lIGanjkIHO/eobklYcQQdt8jZVL/AA26ByghlYtbaIL9AT5wzBD
d1G29Ze40HjNwK+epurk/VPUeOfJaSUDFmioIhsP3nS35PIp12HgBSGzvtvYCrUPTc4upl3UcMeH
I0E3VhEX0DNMjJU0nU3fb+xEc1fHPEBRTlOGCkMK7bY3IctpWKzfeT0pG6EzU/zSUx3ajYVwUp5W
ENGld3EVUB92zBQa6cL1hV2CSHAWJKiW12dWJjol2X4ugVfnPIgP9A/9BD38ENr4k8JEn9X3dh4c
ISEcn+uC68J6PrFPv7NSnhs3wDcSCZzyZjlHDR+QfwwJ08LfkrdtbSFh2r81rmUOBC14b5jc+UkI
gs6eeHSNp14VQlsyHWTBQ0PjaZquwGKSyPkA7uMVK5Yrw+U6jBXOdqp5aI3ZavdAonpCZXhVPnvr
kvr1eQaMhI4O74KoaYIBRXRd9TsxuUhry054U+JoyRv8pJQb950ZsJRFkux8QVLs3Ch/OYgGigbX
mj8gPBQp1BF8LwmMRjor5/c+IgHijKgzUsbnsjKXcgSfdxfc27Yfkq755T5do0ln2JzB82sprJwV
ddzjHw6MewAo/KBhYmHRilxt/M7xXEtmhOZfZ2sh18IKrEq7jZ5jQLtLFBT9od6bsfh/jXuBIEI1
2jlWkpd5xIjRPhu+mvM8x9pS/SFsK2h2lJLTugSiau27QmbFfm2+/CrqMHH/EWGhrUdm4W8Emg+2
BN47oLRgRRG/i7TCLjYsWQeuiP7eMkGjj8CJgokHOHBD/R4S17g6tBdMMhawRGp9974Xcxw0zfZL
b9JPM8wV0vAH9ZMm5yuuSzUKLBM4LxBEvzaFQZPglnXw/fziXTH8EgrcvrikMH8HYsqjEceGRPIN
MUBTUrhFJAUjo8OrGFDKCRLGdBX50VE4nOPtKXonfpQ7HYF7gevRDogCJxuNAuzLIZc/TbqK7ztV
kpsXl99qnj9gLFTcdh8bZwlHDRZ3zdKtpYBsF8H3Iw7xwgqFwGlcoAG4ffcHp0nvJ5kZID4iUAsf
tnDubMEYXuGy1uyhwcJbJCDSWqCv7NP0PkO/bG4i9rrreicnUzcwRdvT4LFVhCEILBckNdYn+b9l
TeoHTDIC8wv9ayAWG5VYNr3zSYAC38IU59YzhPJ4zuqjIPwR5drfo+HJWw1SdOa0qz8CBO3zTUtc
QldQCn33hhD7iDGUSBbblcBkt1sJqBW9wIWL7ftS3zuOCQwswbchORgyO02bUqpqUBjXlmI9PzSh
/O2NBLEuyPtUCOy6b9Hr+nKyxQGVrw7/D02hrwiXEbOxrGTL0ZDZWc3OOSEkNUZ99jouUdJJ26P7
4y9LezhxCB03WMgWAmdMjjjaDWKwzN8qqjY/B+ztEarvOjYg2x1QsDHTDWXMVO5U+NCqd4C/ChFx
wIbRLNe1UaqQS1/1z5BQFsL6/1w60COxe9bFxv0VqspsVon1oGsOjSE6Tv02P4Qx0AuhexEGVTM7
O1C5Twh5U2SlsfHtt5lPs4QK36ugLvVbK4YEuyUVvM77fIOscqIMyzh6a73FKG1aZkOjt9Tl71dz
RqiV885M+J0udHEm2VrMAewWXbdvmsqG0hqMUBcpwT3kC92frFoYd37aUSEBWzGEj4qMhZNr/ETH
8BYsTCkX1oWKtoXaUq2LAgqpoZkSBRqB3hfxtroSYyrJxStq0rkPlr+aDZzwLAUqHWC/3Vs2ZbuS
FwaH6D8otBE1G49o5WPQ8HhRWlJN4AYsJTloFWuCfI6DKRnP8uVau47nrS5SnGv12pVHcnD7JFxT
6iWS1Tj7BGgOE2QdN102+aLBXidsdx895ca37PstKfzTI9IO7aR3jsm9OOAFeS9EfJrtJZnMkmKx
uQBJbVqPlaLwno9U6V0yEehnXFpZJSj4+CaLaGFh+2Xc2BSws1q8lIAx0Tw0Fh7jgYxgDok8bd6c
aO1b99gwWVEAgF3TrR6nSpuXAX0rzeKIVBRse3vGJTPmaDNrppbMAW4WkmDfBR6L636sDmvMTknL
GR8HO0QhQqsahdP2cQvz1KFCfU0tv9GzQFJtiu5iQZoa4hol2wqCM5GiwSMw9aUlIvDdFGd+kCQO
mECD0FSE9h5Fl86J4qdIJB4z4ERof/rbC81iACtdlmxd5yjv6DfFqg8wAfiXumpEeM+C1ifjv81U
uHDQa2ZqrjmpuJxmjVQmRkj2/fKuV0KqP3Yo9TFwVEWIvsaqhrB3A+6awmurns1TwYrgTq6CCef9
BtrHP3m4m2RnQOe9qQrEHGIp22pkCnJwDSsXbVU5ZcxWf524JbxPiZaI/+ZE4k7SWQtkr0zjp23y
4EVfm47DrMMmwpqLEAiFzDt2UhEfhcGOgK2EuIxiV7Nlr/V/Lfe3JDXrIOcaHZ5b/aNyfkuNORdG
UQucLmqjnhC8YXZi5NUVuKbUda4WzUfWoO0+NZxYbwOQ7T/rH4t23Zl3ozGeP7Jvo+yb9rw+/e6m
jVsxPluEWkxCYZrn7g896s5qYDtcBc7w7PtLv2cyVJiSglIOIDNZGg45L9fIYPI+Tly3vVliW23L
w5Nscjb9VZ8z0D22x/f6dopPXqmF7wvKvX7mauenfBceMLkmB2bpqAY4ZgTQJ0Bx3OtGJIzBKtoI
6kZhOw8LcxGBDRqb8rsF1hZ12I1LiovUvuLYIxnahYsPliTizOD4Ttim89DAA3bHjXnz5KiLSzel
/+aljEiGoCMYYbPXPZFgZIPEJWTGLFaTdz/m33M9TURatgC8lZPi4yyPCJrwdwT0AuvF26RJgiUm
qSS5OwHHx/RHUratbu/GdfaLONrbwSeEZPPbjkF66dI5RkyjNPwlVEDg2ueb3aGPuw1ZIF9YcvZO
QfH4jByVKj+fRWwhzv9VKM84ruKEn3+HCktKinAMCeQIogMKUc+hRdyIAcoi6u4OTG16TGI/xZUk
zhedGcuLX4yzFObpZZLckdVBvHZUOnHJLtl0CorXf7oClKeZgOxxwz5w3zx0Nu/4/5o3Fuis2pX8
NZs7ZY+ocqRRPq8OGGBNcAv/XeXWCsQ6s062QLmG6R9Cebu8/E8gRjuBZvq0e0sHhVeOYAr4fqhy
gm9dNbh+ZC1nTU9b39mDBObZz5JzBb38GTm+Im/BRCztCHEyJwP/9S6vUJM92G3A/3jfuvFqHiH6
dywqiUszfyzgD5W6uQNR+iFlcZ7pNtqZ6gRPnRwb8EWZDn7/t5F44ZEL/Tw67Pf1JLJbPUggh6dA
ALu2eZehs5AOA/2Cj8r3CCDi95I9MqXgDg0oxTsAQQcY0k466AdadWOGK6iX4TenfRtN3rALO2a4
ni5xIH0eP40cF9kQmNsumEEDYaJYCcrrYgLUwMH6JyRkKrlVvBr+hWPrsShaeVOl3/Fiv4qOsQKD
6SuAauaHGEHDxSyG9OrjZFfwyDePrdd8guVEKM7CNeO3MM6+qu+sHAQ/4fKYw4jBa3x5PDXGX05d
X5JMQReNcTngj6B/6XHY1tQk8AUQimVXDHjvdiLzV4gYgtHzb2huXxFXzfqd9KzReTPB38RM4N7k
onj86V/xMY4NTPWb8MiSnRKpiLoL/KcWccEivg2W4sThzG122o9oyoDpH6uDbsDTjfBVb0qQszgu
USmWmTlYEM5rRnxyOQIGo/lf4VLZgJnLA5dlmi9raE6uwXxGAcfPSPEFVa7fIfMRoP8RqVvKXKqI
zKfidH6kwtzPYJ2qitvqRUx5fIdnNmZKdEv+9KqwhEJ1V5r4kXe54W6SbLW/OwEA5fe3MPB8+far
f8o81PWnVZEucURaMMleHIMomGSe83V5OzPpDDS6/8cLmRcc49TlSpNfqxAr4I3WqmDBVKEsJglg
gGOQbf5lSZJoZ+ShviLxEa4ZDnfbdq6tMTkT2b4lwztko88bfSKFURBpUd3Wmy854W/t+Ir5w7O8
Z95p4Reeb7rzKk4eVBC2kfKGPyVYSysDztLg1wROxBtngkiQ7HE9BLMS/B9F7a7LXe/CEJuLlE88
BKhQdGsO7MXhL7I80v/M0NFRFjaZghGovMOrwKDaArfWMXb0r9UEK3J9ETDmfW4U4LIAYyOZhl0H
x9iYxLA9uqSDfzo/a0oJVNFvshM6Fs6WIQRV9uDW0velGECrNQ7GjtN1E2qO4QLm6BT4gkkXaGpw
8YqsheMU/EySCifHk6CQN90e0+aDqWv3RojomBdnk2+3+9R87iNby6RAsZ/4lQcS3YpxsRDSSXtH
AzJzoOkOq5Bhctiu041IVh3wCbR3ovsgTr/HE0Q/KeVK3+L04ywpITe0xFT8DKCVHKiZlhnqTvRx
q+sGm6zU4roZjd9Ao3GNFR5YSC7N7fFw3TozR4SlUETe391Na5j2+xcklFUK9b9ATacuges/BJlv
vn72aCjFUrjDDXpFftMrbrplFK2pFrmE6g1/xv0Q1kSqeO5gI6tufiONnGHOiSPUmjyGx8yl3HNi
/TJuM6Kp4Vq6vWjMEcn91i/IMcUEpccr/OJjzyv+QYSSjEwGPFoKgxlF3emH/CsLFwZ1yn0/meRK
Ly/O+8faFb+2TrQZg6EBb7YiVH85L01LoOp91l80hY2ieW5yvDaEsOMy8B0itXanTowEusagWpkK
3D4Gd2OTCBsASktaop3jc4HPrs7GYGf7pN1cuAyUd5PPuE0vTStIKNrRf4mQwUq7Jv7iFsASPLFQ
os4gpVBkCH01vH4yizlnY1K2La5eSnZzrtPMxZVugoref/9iChnfemP+jYs0cQyB8yLRPRwZo233
CmzW8XSwSITA7PFylpnzJzaveGMVSIv11lTbmdGLR0paW9t76ysGb8gSQIg2hoazBnpgIoAyNBHP
E43IWdL3sdDmXt8YJqmT/dyTW2ecah3QWthRsqvJJLNqvmhCRvzCU4R42ISSYZqThGQTuybUNe8N
YUkNHsojvrI4hhTXWTyTvyJkSsMbevDHP4Gfi7eoIDkUiJB6McwxiOKq7s1BTk6xhOsZDhKChGrK
G3qlke1ej+ojy8ciN+bH0DYKEFMJFw2K9bwAgPrzAuGfDye45FCRhMDBdUrJn7BfEZv0wcEruZ8X
WmEfjmiv+TJBCX8Ul3ofIbdvxSVEi0X761ss8nAhUmYeRa+jSSzUNL+RqgJ05zs5MKuuLHEayr/9
1PACX0RMOvAmleEa6sxscCZtHJ6EoA5jjG3jN13THrSvyWvJvx0Pp6oaX2e8MVRb6g44yfmtIUJ9
H4XnXMnx1rSr8/iQYbFxsvC/WB7yaBhBYps9wnMlhy76j2mMKSxbojVwyocGNPYYRP4FbeYQhUNk
8b3Iw/MP5FKO+2hGw1MjowYgZrExlj+Gt5e1yipR9ONkLs34eNS4e/Ntk1BnJ42DovnHc6QDwTOZ
BHWWWqtuvXJyChZnoPX/03ov+a6T81hvgUsjFreu+ZD9bveWl18VCPb8K7OzJb4tbu06sP8lzJcI
bG45Q+5vkMFwt/BMLiHtZc8dM94Lr+2mQHp7TBkcBd22/LlZf39om82bJnNKq9Da/hsh2TaJQHqO
NpaR/UOSamDROIRL2lbyfiGmmG4tjNhYUmxxTpQLwnxe4DANU7O9wG9eSdopUIJe9aieWvP8b7Vk
DqoR+yBhohrEtQrKX2o7eWW5xRvcZ/ro70NVq8rzRmedAVqDoycJO330qSBlvzQYp6SXCGNuvGrw
lZa9Tlhahb+oouK5HjR9RIaU+UC0SM/uCIfcAmz+6ErzoBYPLNMX4ffdyneX93jUNjceyg/BpQYc
DUfS6gghWoRcmr4XJQ+MCOIoqNjZP+ldVvHSlocuAydNfOmvx1A1wi2Wg7mCKpp6aTLAYGnwcv/x
v9LSKhltawRqFMgKEDep0MiAQKUTdWghha6ip9ooR7diyk3cc0LocO7mcEwzHv3qVHZtQSIFVRjK
SNQDM/qtJQ2rcJl5iIMSnZbpwvgAt7DxKRgsDG6oeN4TV3CFEu6vLLobmIQWOQj5w4nU5/Eu9G76
9GGTGrY30ELW47EUEwOmwAH+uPt86aOf9tUft4bAww7G/Av/qcxAoghkozc13n4QOK/9qk/WGbG6
u2c4lEypLKP9Of9uKvLx8I7rsBq8IMpJASXqfGYuV3A9QQkuJspnARfqblcrgmq2ZnQeoraKa4xa
m4TYFMKo8lS+EJ6qh97d3QUPfIV6v5H+MCREXbvDaDZGIPmPeGIJuSaXKwMfFeDRnFwM+jqZQGvm
VsJ/VeScQL6lurddLRymNKkevBfCYrCr6MG3n+0loMvGM1CrxaC/1FDpoOIhNrKPUpMaMalc+ldX
R29eKaivyqWsf2gxxKiPn6txWYJkum0ybFHSJEICjZbylGMbCcuStcXqQbWadXninL1g1xWlS4PZ
MdtWxMyDDoOKDS5mEHophH3xA+6g88Y/7J7KGDyZ1dZLeSwnmSYcwcQtrpAh73k8fey46uZnNGh9
LutIUcNmF2BwUNZkomfyRVcDPB8WHgp1vWrTKQg5T3N7lfvZUrjLDM6ylAclbFUzzq8XzCFV39aA
Oex7ftWfLImOLBQ3kqH+VAAzni3QXDNW0XfROG2/53UExJCMi+810a8/wwcxZ9a3IIbNvAGulNnW
vtzQXppuucx52xbLhC33IYSgim3u5FpQz/P3G7ueT9CcS1PxiArRP7/2lNXQtuFhvf61M7ZaynCV
pleamrsgOI85ETH/4dDh5ramQ56Fq5VRA0kxsavQw+BChnurI8i1lbk4V3cHgXo13UAw3vPOQDfs
fCG1Qe/tMqr3NWP/pORXwXkm8vwf7WycpuzQMrb3Cdaxzij24QlnMPaTEOmbeBvz2sMI19CUw+LH
YToW6Xcyy+CHgkbB7P2iF0VNzzn0andYaxvNlMhkJOxWZ0LrpJozQ8SnowEboh9Qxl02ZjaYtQDS
OVIPj/kbF6T3ccDKRY/nQGom/bmub9sEb+Sz5eCTV1j4iL6P8CrYMxQxon4XvXLl+J1PeF1xJTiV
ep//0a4EDD5UrQgnR1JHrImvk2EFniWPPVZJU69xNDVgt/8S5D9Hbk6gVS1fKCOa0eTIvGHawHjU
QPpJzniHuVa3wUBdPam50PlyaZjyKXrr2gFqnkVd/LvONpyqJwl3I2cWSDCi2Ld0yoZgzPhLNm75
U8LgZjAIlyRBpf1nJ80bVVkBUotubKCmbEN9lPZ8rmEjSAQM8yrdzvwXcs7usO7ffmKZShS7ZRVa
zn7e+is7RkzjIeeIpAMVM5LBrsr/6617c0Er8PAfx0X777NJkgGiHQTlijYJhhYUBR+2gYqMH8X/
Jha9nLZYDlXQQOMrA338fiGd9CcYcrjNBkAV70gJO/DWpH7KlUuzJrbTiGZs2sKmsQgk/8yqmsEo
v1ls3wNjmhc8zl0J52mBtgDkFXd3+mEyRuYCmdmGxYmrnZ297n9sdoeDs3RlP6k81L1tetiJG0Al
rfJCBaRewYku/6ZCBhzFCxrsIALXkUxw4jrd4Ye+YTBtapLhIFvSuB53tWmjkbGjpokYZ2etqmFI
/w57DOzZ2mOoTuWNy2Rsy0ItERqFPN2COnYmZzbHHm7+5cCNJMIVEAnPOSahZf+KMPIy56fMTjZn
hQsRYUIVMidVGRzSyCum91Kk2NNp+EglMqEUACvTVSXtBjNX3+Xf/v5MOs69j2ILh/tvA5AADx6k
P2IDH5IZP22JviN10mJbldXgwR29eZH2q9PhEGmrrWCtHnpcIAmwjPtMpqFpUrFZ9KOopSxP88nK
xi9Qa5pZutWsjC9EmUTH20sugXmA/kdUxZUI8SrhAvEPg9mnqkiYi1RhGjJNT0A3hEB5EO4zhL3C
Sc5Rgy1Ui+du1ifQZxrtVwhWYz83tsYk4531MeMiqrQZ08vIq5fTQ2y8dzmwTFNBU+tyDuYqbEGp
hUyP4VPz+0DXuxbpIclI5IkXivUMefkoVQh2DuG3+I1hAQCD26dI5F8UTMsxH3eOPnIA/4VW999+
ZBieSzkgwlGz6io1tG9DC3Og15/5opr3Y/6aNenadw0kYBxkmwvoKwQlTiSxNLUwkFLEFwxFzqHK
w4noknB6boSfAew/4ofnlctChBGud6Tn84FKshIXiiwlYhmpunLaRRNl7UPRKJDaf/UVCSU5W5cg
bPnPqgOa2peVN9FJydYUmA40lzM6f4aE4xd5Pp9pGJKJLLb8tPXcolcikDjYgpic2+Izh5/0kQ64
56lsuz1Jfa4zsNknxotxkDXOoHvCfjL/5lQvWzabFoRL34SfHZ1mCkcK4fRwjcRNuvYolEZPUx3+
YQTn/xo+zv4LqCgxY2ewEdn1EHsVYWpN6LSStodk6L+n+V32Iz1+YCizlc2IzuTZSGtVVsnhuX3T
F8HmyD7R1Hku7lR0S78YcKU9il9cJjrjvPJlUM2otEF9sZlYanp7woHTI/jYzTWuVTuOYUe0on0K
OmeheWtogvA8m2yROkQCHkDqEmD6UOOVjgqOGzMcQCEYbuwp54NGq/zfRDW5FlhxPpo54ASUDIFL
NIS3OSS/zyQBN4WCuIDn1f/OxkP5XOVQaPo+YQwzCmc+fBTpePOiDMWwctT6S88lhhIEMjy+pc22
bo97/4FzZHfUEblL+1QQyBZmV8cZVrh3tyBRuFAkZYekMhs6HRMGD8LcUxYwEPgHZLXr1LMIKLG5
5rrfSiYRME27182mfuLpujmnXrqUwJIudhtVMf94DzSVsfyLsKyvKHzsn3Qvmx8phsn1EOAT7mxQ
P68ofPdI2HOdlI54E9jUhzs7nckCK5GNvWylbAuMz2CnZbexfDZGOJmwSpM513PG+mcnbVXHZyu0
Wk7pzNlCn6AAtmSTIaQRpIn8+OozU10nVEZTJbV0/Awal6F84Q90oCadUGdxUzidQuIUF5XWk60U
TR/omf6gsa2NyoiuT+z0zcRrKWl6NUc/Tc8MnkzV2VirXK9Q53Rx/f0HUYyic46JCT6VqJyWhbeE
hGP1MHtmE0VryLE7Mpuh1d89ro3IDpLt/HY2x7qlTjL58yA4ntTt4hzgZOU2Wy0SbyG5WsQn2KAf
06APdDxApHxVaMqQZCtot+DHc2wQVaE+hTgWIh4Rpbl+XOUNU/QD2m/kWZIw2u9kiDEUlD7yL5af
mV0aUL3qYjCeuGR9wSUCZmuCDh3lloXAj0vj7lZr1e95a2Y3q+Ox55MBzz2eZn14kOP55EnqWt5i
pZfjTHERqHeOi9NEIjlsOcHWNT811NHLVqkCQJttt9ctkZnhoXbJKCMxzEapmRIHe3v7LpZ0f1nU
65dfpdBTlpROsC+B/Z3M0IfElYNHzl1ZLWvkKVjoUH/QQRTfQnVgcCDCVvdcY7UX+romfbiskE36
5N+7vR83uUcTclIRSs7kP1O1EtWsVq6Qd97TDtyJQOi7KR0IkZmyfwRiNP7KpHMT6DPYe9kbQV+j
CcxOzxXqRTzwe3DPYDA3xz3rl8fbMItGvYGrMp5qkUZFq4WwfnkhBh/vwjZjsnyxohovDaRUoz86
uIWLzdhIcB/3cHt8256DyVHXd2ANJwb8VgU2iAiEN9cYLH/YUSaW94wEsDVJMzsXgJvWWVxkdND8
KG6qnTIPydc7Iprz0gBewf4XydA57AKDi3/JRzoBpppRPFA4p1clhw5e7o7JOPgCE2rGx7r4+fCb
OX1e/+i5BuErXpKoTNT3Y5+6CLTvxuiSrRSmr6pLWv1BI0CGdipX2sGim1h/iCeoyIC1n2EMI+FV
wJRHpy1+J2Ja8nh+CiMKOL3iWVPHvqaoALob3JvVHOLDQPQrDPgFTkyyDuJaGsqj8itwO4Ua9WUQ
RwjecfKsUQRzA4TwybkJsg1OMCGMxnwVtT3nQqPKOLOa0QJJHaK7Zy4U0ZNb/vw1P/YMVRhw5zNe
5Pzbx7e1gHLZ4O8nmy/13Aibr5kC9u3SuzwhZ5KXWDaPZ0MjLj+yVgxw1JB2P0aKhItwQwUfv9XH
8mA2K/SILZytoyvrMk2V/9Sadj1UcbvXSHmEbK83xcpRjJgkY7DT6SZntgJzdzG+eDLg1djOFahH
12drCCjGjuMt2RKhwL0pDCOs8AeBQ/dYP/tiRNw1mr13sDKcEHw+L8+FtqVOzGSUMuhqc0Ynfh7X
NOMKXBYs/Oh0r1fRplaislXW9U93BQMvuVAjFUR42ITqiSWT2P/ws37QkpBsiVF8s7w5SNrAr8xs
ux98hBtsmS4DiBVY6aU1ixcmXJh8j2JBpbyrYI5xYa/lzeAUCBWfHQW6c6yFtRdG1SgpB2or3JpA
2cY+yOXBVRLzvO3oTbMsbxmgQ4spZa1IFU7gJ+CToz9D0rDIkQCDvP8/9r/m8SeLlexNbtB6Nupw
OoUNkEZUhN5YrFVu9SZWHdHHhojswLs2b3KN56sso2+pFjf66R+W2P5Jy7HEjmUEmPqq9lqFhBUC
Btv8ASRGyFjx12MP6bD+dBEa2BVkiNzK7rBmOhg3ImvKQOBfTs6OnByJSVs/dV2dDAtJBrefz0+d
VXqOzni178nXtHP6pWpA5ijmNrKXC1ZRM1kwUj1/vS0FcSLtd+fSYUTBinLnWHMG/U17oGGi/L9X
E4dNyDqzTWgFjlld0XwrVqizr4yah7WgXlBFsFdLVpTbHgUoPxtBUDSbwWp6Wn/vy8QJBji2CVCO
uZY6WugSqKuZRGSX0BNJfQ3G75lQ9L4GfjYmIeyyVgK7TsKd9chZd3F1SS8KnPQedlLTqoOSHMuA
hVGFxApVJSYz7OL8bqO4Xx3lJug8vUAlCfEOzaY7hoyxJZqLTgw5dUZopkxQBBUGSLW7YvplOaSB
R/eQrpNiVS1FqlEba3Qb0VgeQJ7qtkYWLCfWQJJfl04mnLvmQUQuZTo5FemYgIw/PjkKWliniygP
+KKTyL0EQImylMtTqcEOo0gY/GEEBf4w+PzkExhXVnvzf7LoW7gsaJdo6GLuJGilioVtCjiVgGNA
ZUXkSSzr2cnnLjcHSKcouwM4G/Y3qdYK2L2ZmwXwiYVOEoLSZdPm+/f8LBOxrP72MC60ndHp7yNu
b7Ontkr+vT+HqA2aiauBZuWHYsDPKIQ3zhIzmDYKeGmnE0+SqB873ggqNWC+up/nvLqjFd+9FuuH
RVFZKgI3lHxxVXiGtw7jyyXm7lvZjuSFRQSxhtEoDcoEHnVSPDuNyPIay1lR7rohJ+MljeRvX/qU
fehLS7I3+sxBZUCj9uLC0MkGX8qcCFdNnu5d/x/pxwWPFz+y7Or+oo8Ox4nC69u/luZ5Pqmj06nV
vKqXyn2qbdSeUbqW4GRnVakOYTIDi4pn7wPR0zLfYUlHW//UsbUxZ7Qa0T3IAfkrdlH9HBB68XSy
dCc7W0y21ECuvemBMDziGC8PkHWqEBfm64oqY6BToWyorN+4EU0csaEnJ+tPEIXC7Omm83j9SLnN
FCxfAJ59EGis8Yr/yDLGv9eAcmPYPplHe9Hklw7ykMYR5oSsAVZkgMV1gO/V96SyKmXPspUOQyrY
zHVZONJc0st/B9hn742463fna5QM6pzpWcmtnWUbFEhF+u5BK+8JRzxhRu46MvRB97AOzhDcqM7c
9HsxRVtBG649otft/ewGVAT8iuOUpC53r+yYpXMi+k5CrmzaZoCVrbh+ibaseIUkx0lfHGtO4Ei8
DixI/rA6NFMHc7aLdqnZIhgtn+crGs9BVxO1N5G3rXfcw0c8TSLsiwge8+KIhe1Y9A2PvrKUVAMj
o7MW4wk8TIidrK2XjE0bb5OlhMSyhaUPjwBw+YdJlBN1oUhVEWnIN66/0usc8oruZ8gg3caFi97H
2zoS6qs4QRsrCjEiTo21oxNF3y4Jut0cSowWwu5T+qi0T5RI4oDoI3NQjkuMUwsUhHBWwWc6c1mb
nIEOD4iG7v2LKb6TZpYORNFna2+NMM5XuJXFpZDtFXwpT1rxoTp9AJm7PL+ImUFw1Ret7TNBfIj7
WVU7QoJVnYszrgbYoAy3judPvjWpQxyWcWm8OfOSPnShlsI6O0J2P3oNZEy/CblfcMyKJjjClSs+
waxwL743f59sWiajqeYHf8ca6kn+0SOFkdtJP/MuM4ZSdON1VhvJcUSd0k4cqI3Sc/Hnhk+JQfPf
ZC6g0Umtb/7gkWcG0mCnk4OF62e/NXkq7mvwFJ8tL97A2bJs8oljQfzvOfjusU82mqemgOIexz41
t2SbK7jbfrwqWB/Hz4+cuDS6ffL6OKVEEp1bUX5PKrmvHrJBJP2IDPDlN8f9Bq75leU4Okliz2Rm
HTTnp0yFosLvW4lsIe0QpoRqYHhDM+7tVbztCjY9VRK/RtzkcYknCnuMNZnOPCyeci/K/8MlBEwR
3moxZgnBP3koSpYZRigeJn6bPJkqZ2SrbVaGrfZs4aLcUTxR71MXHkM74x/rcKxJDM2rHMc+kM/z
NmT4hzx+HQDYsyPd21eh5vGWdaK394g43/uf5iKIrnuvl+h3ym0AfOct3e0jZTGI/cnohGE9+dsc
3pKNYP9BGxUOEqKwUTL8padftejh0MH6nF2iYpH6NavQGY5zTpCIAYdgl/HlUqiN3RjvGNTiw2aF
n97v/MXQcqM0qA42Ajs7UKpesOwwm/5/DoC+wt8HOFvmeNkY20u2XTnQXiqKZjEYWNEzH+9QbzwD
ODez2JcH8ALbVix+lgrnee5003ZkN+LnpBl2S/jmTh/EqychAB4xj6fNEF8f1yo9TtQqyUDgBLTV
vGc5ocf1fMON4IBsK14ygaO+T53woyP5Z2InwSx+uSwM0Lhixu8KOR/ARP0VgBH6zoJ1Og9/m0Ph
WEUck9UDfMIthwTGeIcqzEsSt8ZITmCojyhTgtoR+nj1Mmbv5r12ikT771BTt6FhiWjG5zWTbaPy
4XGeNnK0pTxwgbEDxaZxEJqTh1FhmWACHsbiVN5n4x8B6qhNWpDxejIQlHksgBQ7LdU6VmvgOs1v
jXiCs0SLz5IfqgLeBVqMKE8AsM/kkddN+mHZMD1uU02wbC+Zc95JOG2KP3qCxExVkg2vZEraTbDH
SVmgtluO0rdVxU79ZJ4jj6st22tc8QnDnicvNTUUdU+YZjpSvdtiFx032hgPurRGRuKUxl1XPoAb
/Jm8YG8r2p9KEl/o2rOI+fipLbV58u5zc2k4cMOv9JmfbLI5EwK6Ww6uAneY+1u4buMx3O3Y7MZe
sjz4yKXZuPLb+aBOYtjjcv+j3aVfwSjyK3DNe3hWCluAMH69TD0/1AZzGwEZwtzwBx1giKH/DCJs
+nf5pvHHuPGp1r4kiARPT3xXnvylSCgGSwS7O7Gnk+DIrrnogQmfmreli4z1IsT7xKfGtJ7u+7hh
P1HqnK/ZQc59LMDc1fkbVnUfL4/mEDy62hIcsAcramkxFAzpPFZIhyAobW6AQtUO8UDSXOxP1NgY
6ppLlT2er2LUOHY8ORjdhRv4u6bfhUhIHK8YvoutX+9q4bON20x4JNV5JO85EBqA7euBvfMv3bAB
yQGUBFZ1JVj3VdKrj+gvjPwqvLZJ1pianikXWYQJxK2r3ThyC0RaLl6w4cPX4UVCtc3s0/dngsO5
JjgrauYbljsSVbngCTAlfH0gT96MWaSfgCX3KvQ+ix3KzMRl8Rc5zhqHy4h3DxC1xInCEKwwJYAK
P438oQWfgTDlLDHm4PR9qR0gQooRUKv+VPcXu7n+CYFRXVsWQ1mcr2rJ51jusskzL3cOalPTiVR5
cwDAViksKFrsNcWorzE0/Kkb+Zmpl8HNwQ13U1Gj0EiKJUhh6lQF2uNDxepEdh7/72QJ8PzCExCA
ouqm3Atdqwt9yfPYQex6CqSKg6O7Aac/4aiqGzugtxBO2BLmHP6es44ieUqzZ3/L2L9sUGeOSsWz
f855CxT04OIsIUGIHQDjQpOocaPAC1dbF4qDWJJfqlft40tV5rU3qoX2u52MPe6v0Tdj/Q+qqtdg
7Hk2W1p5LAEB5I5UzAMqknUnemTeLKVeOgzU+f5vy0xOqfi2/EzBlpgJ1qLZD5nKgWIihC6ndjzK
o3rtupmt15qcIwRX0x6ltl4BMq+DEiA0pHqGuv1RWSxCMUKDXTyif/xDIi+qN5C68Hk12BdAzy3z
LmNxUjoA0XYPgvE80yhhEXC+oId+UG1p9Acahv0p0wYn/AlaFVq7Yclbc52Qyx/SpuHxSsSp9Qps
E9DAAonEvdl+8Bn/xWIiEyzi94kQxbJhU+AF1qBC7mv+euOJ2olF3Uz2rCsTQAmpveAnZZGkTKkq
UcfKeiZ3mt6zN0SHzz620ZEGDEaLZGF34w+39qdi5EarI1OP52542TPFZpE0S/WEOEuUXYzqX9Sj
O1PtkejyAJQH2FAs3t/5rqktUWJkmLL6taLcKbrOhwysepXci7nVs862dPB0S+QZMVD5+zUmHijL
KyE1g3Uneo7oQTdswRFjMxt7GwjOH9hEolhUHTp8wjsoD90xr5S/cyiBt0HITCQxRhNO+dVftrnY
r759qsM/7IB5gd7rMR6+sU3m5xjoz6oby/0EQaM/odcDjxCf+P+299XqpxjhQoxfXF7EC1/J+Z+n
RXY04CSEvsJ0iJqOigQxwSwwXYhKBA8pMoQEdGE+ASq8aq4MG7KXcHLYyF16JdZFnbwHCcYcCWyR
YPA34NNb2LJS2T1nG78VQZ8rBfKd1HJKsKxGnNp9VXzq4AiuDTa4yKtBRBDQzp3DMp6S327/eJ5G
VjVgJCNxaJevLoP1qoLFSR4x0opHmTJk13bkOZjU17f0qTan1Y2GmgXBI1i+HTA/UYUVZLH9CAYq
00A+Xn/AUISwlrqD3KNisAUHGznXzl1lHBMGsaXHtf0KJ74xwr2nKmmbUsOdsu/iTIkuxHFbn+MW
06S2lFrSIzRVNGtddET1BheoDEF4qZ6uztg+FsTQHJpeVdzgLw5b464/bF5dpdxgzLS2iObYJ85g
/WYd2YtYJPbPP7HZ9nI2eS/fI7wRU4dfJtFASXBckbI8m08PZWJY/fi49s0RyEqxOmYAKDKvz6+3
rsBrai72QmykUeU9wV0vgm4ZurzHpU6sG+rgSgVQwYCA7Z+bis9iqr2vxHCHB3oPzh6XJRYGBXFk
NfH9NrUhopkgfv294PKxCE5GNrlqQiO2kbYz9qw8kbpt2z2BE+AdtUOKGbGK3q3feieVq7Ok7Mv1
kcRdDBpS+EdoxcmArJ6ssUuVKlSexLZc8M5WlWrOco1h7Q/5ZxPfETm2hmF82EBflU6AbiinyrV4
ISWZ+5eA41ns9yILpoDUk+I6TuD6VbzK8pjsslJ0gzZdBttNsgipkkcic9pkbJobRI+cub2oBAE3
jlW4KeqYszJPZZLpLCybNAs9H4PVHy7Sjp7CNoI+WGXC8mL9jFq9WYNx0cbJRQDSRPGdnwxz21Gb
a3nGflEbXNswckUqHYUZ0IrZNkQEznSWx8N5V+wwCnk1Bsz9NZSBpYOmWB/vFs63/M5bS5Wjs+vR
EDKjXXE9b3pPjceWFMnfvh4dSfqvosi0Dg9roro31CPlsy/RWUPj7dLXyolimRKD+aZ4eM512SsR
EoOyW0TrKUGYKe+jK9ESes9Hz4KHhG+yEiRCHUPqevPhtNT9Oud0ZXEJhV5D5GEFspdNroImbUSo
9/p6ueXGRQG7toOoabNmXK0fYVRhE234mzMmJoHaagsRrpDv69JDZf7sYdW83/qXWEN08silxQtM
kPTSnXpJ2qHAYGGBdFFkmpKW6J931kH4qFI+EbdvE00i94/LNpMgZpenycufYTq8R6gcGAiv+RTr
CIzRW4n6Adfr35D8HeotHVKrTI9MwCDh5d7HiiQ4rT/xcGgpTaXObzTfg/eBODFXWuJTE83V5Zji
HFK24xbMga+7wXhtj7tzcTOjSUHL1IXjgawSsXrvUV6lSkReIrOTpmE9i9FeMwg50NPpcTRRIk4p
n63QI2hzjQUeD/hZ6Gy0sMLH4UsEotZNh562qf5ZNLUBpeUajw9m4Z5MfSDDuvKxIx4VE1Jmgjum
3hOz5VWH+PBdSb0EIWwIl6viB2+W9HyC0rJ1mAdMLzyMloZ0tvAQWDJ7oRTHVlhAr3AmHU9p2vuA
6/MjfUnQXEQ4JGBpoArg86xLOYIn/pzU0LAwcTSaQPJV6MWQ6jhnTqr2GXfz1NLC/uLFgUefKe2y
6gieZHNxSAt+1xP0tVTvCylQWNFSk6mEysBUVD69MtiDjSF+bPyBujDRGMPKe3tOcYCi0zEtjyi6
Hv0IKtQGnVBtmQK7Dn418NzVgZMcVAzy/7CCa7Q9ykR0s/nCqdK6N9Gcn5IOXPRasGLxmzIwDVLt
0+Ql5ReldAP70LibOJv5qGdK5/7QjveujNuJZoolopSsxCcFjmLg6ZW6sL64wge+/DB01tR/yMMr
UEwEgd0oJsW+rLMVLtgitiBDPdjYoAsjsKeW8XBfvWDh6fRRv8yoBSmVo8pLNa9k6du9jbJG7a3+
XVf/cQDUownykCAC7t7kjVeiWqM2oHKzyS8mf5T4/IHUKjsLXwUDYV0tGOk2r4FYDrnA9nMCVjQC
JMeWo5brIdF2P00Ms1ZL88RPM0ohtJ1A47AYlaLYCGHdCuqm+Q5qSzHZbTgflbYJrsYecF3bXCu4
8ZLh09NiL0Fj1zgjDElAz0mqW6ugUlib/6thlbIiYkXVs807TJpRgebIamf6uT8iNnA3uBzeza8+
iJ+3vjW/NHmMhaaM1dIGsxaaY5RnA/KPoTZKkEerKL6eRYXpO3dd6x/+e42G/K6dPACIsmNfeERY
/EZRsxwGH0VfKvudWS27q+Qexc4bMsljZcqByx5UoyAGcOktpsxHon2HXnfYALGu9Mok7N5T/F8x
ZcQqsd9MVgw2GElO0zOYjB7Ck26IE9FTcZ3/jziXJDGgcLxiAGnZtYA1r7QI/Nbpn8FdKUx6O6Vo
C8Lggd3+SqQ4qtjmLh0YQaol+X3f8et3u5cpXPFz0sQE7GpfMpq6krfFS5z0Jnl3iI44/1IlLOKt
jHDyMntyh6YyUbykufP++84EdoBxTujQpWKdMihkggzPFL+eFkbzGSzeyHbDwownCv4GOkM4HfUk
GUc23bUbg6Ne6wqS+F3Yde8Pul9U9Ri/cvUqFu1lRX9VSebJZQMcIyLJ75XQnmcY1cWK+AaFniSd
wgkT2zaB1f48lQdI+UY5rfgmZ4zFBaS6a2CmHweHJBVr4tMDhmxSCIK7AGEDjPV0XnK60T+40TSJ
7e+R/rCtbvi3EB4Vu8+Zi25qB6C1FRtWoHTfEAmdhUnx/AQ9EYHgi872KchJX0YC19mid91b1NoX
DuAP6ZFQV1lSf4a+SpV9lIa4qZDUAoxDfjoOawChWGo5APRfwz4PKsTvECbbsHwR0ElXg23Ezahr
qU9EcymP6+FPJpfJN/WXFv5uTAM6TDwgVjN0PATaJ0p4IXqcCTwJBvaQgWq+Jd7SYreXYJM5S1rM
lAOy7zFHt/KUOTbJiWn7lRrJAMvXHsuSN+BvB1W2i0KlnOXbO8vbWnb3wUP2AEcUnEbqxukAwU33
K98sFPUmCF9AzNgd9VZd8J+MG2I/Fbcwf6AiWnB1nx3+qRrM7M+xvU+VqzjzNr1MuykfEbYu5TbF
byQrsu4YIKCGtogIo05QU0iCOlBklsH/u7dXhEvI72RmRJOZ53KK6cHP/fV8UNQS0jnNkUI7ryny
ifBtz09foOF6T7VboXcl0iJ6qWItbr/b+uretlHzYQL4sxKYq0FCeh4s5yMV6jpwA3WXAaEIWg5Y
ktX1yuspP6iCfbMVvDG3+FZ1v4SY5qm6Kh2TDF8b1wG+h9zUK5BworiewphANe1SI/EJ3YOIWFYt
570jFT0miXOLVAfcUqmjRo5zbUS52FYQS8EabPWKYsYlJDoWqnusYs0FzbELYkcTgi2cWoqKlGGk
I708bgc899hUctnJioYtFjWbh3hOdODMb9Hkca6rmFNPdUD82poFZVY8eowXzhDCOZmm1J+CQrP7
AFXSf5jOCLKS43MRxtK/uV5/2gIVZdB/uxtbTvMALBeOcAajfPMkTBiRBj6sCYAoc7TT4iZR3DOH
8vqFvYTokUDOvklkOW+yXsPM46WkMTLNLvLeECb5MnTk6n++uuEXgt1Je28x74n6alSLY9gA3WnK
WTXF7FaobjPS5y8z6nXld/aPf3pV3NJj2zsQcY/5Gstp0DfTOHZSADWnCfSbHXxk4apwEfyv3e2V
Js5DJJbsGkPxbxqrLZ01nWn3VJBEJXpKKO47M6ysNI0Ynv5+wxrj8wWcl5bv9/0Uj3yQ47YMLtkg
BFmcXUcBYnjSigqCOnXHBn6ByPXRf0szMK2gclMLWCoXxWdlq0Brvmj0hpG8lHiEwDWBfOixE2MF
Ghv7r7/dRB8xDIekG0xvm0ONqfRG8cfEXAEjFeD6I6uB17vxd4idMNrf1TxNf7PQnlUElqyOPK7N
MXrWjzLti0Oeyir4fwTYWejb3QpfDXAq0KZ2IATlq5cCcHH1v104lnzrvh2RbVEj3Pob903eQyNu
kdEtLrrHXVlVkGoDomkbmnrN2G10CbwB8xaHYTSQjfvlRM7HF7U0V0G/PYVKgv9Ltzp2SUbUEvH9
suPn7dnpYdQTYVIPvvUepS5dSR29w9nnOGvZw7T3xuaGVcEwgW5GwmxNVwEcHC2DhE2KjKrUuMMj
HRw18RoRrgUSf50mhFf5bMJ7FBTC/grSlogcdCQjwov2izQVS39IC/yQoHJmDUgHWfunHsGdoQji
CRndfEJeSyyl/DRoa0PBhwMOEaTOcUlxVbtIl4NJpFwqcaXN3JKFw5kmoTAAhhXuCatkYp0RWmts
Bzj0QSSvjf5S3F5TTp0Xq8hNmNpXHVU9pvq5s7QnEldAqp9NFIxBxZZBgX/gF8GLAiv+TxNmz2zG
xuGVbndxMcPOMnFT2rJ7Me0DDJl99PWs8SgS9zwoz7QJVNTpdrsFJFiM/yaXaojK5ZnQoOShxuvu
o8FPmlYxwXr0ktAhgAJG6/mSnl+twkwJH1AcWgkrkJ/E/EMTEE69aQvhTMZK6Y0bF4fC8hz91gJz
mWrxLSkNQLNOLKRFT8tEobcttlnbgY/z/0Y7GyET2exMLxQkCYd4uU9g0CX6cyBusovkLmUPvhGQ
vAI6XyR0st59znH+uRIvuPNsGPcl5ZXf5PGBbVHD6wlBwL8aOnb7neN0XYydNQ/b9mIstXnCCkwp
repXxR+IX4GJk4MF+eTw5OWpUGmiSVyy73ZUQuHfzmfdWY60Qe0gOAhqv4x2AtzHqHG5u8o2ViSi
9DvRawhUZxW71hKmffAK9sViudW1anKeSYKZ9aisbwJF3WQn/M32VHZtx4HBFca7hScH490jWopI
vkrvJUoJL/f+In6CZ1LkmCU29/C3mLHvFIgVIfKZgBfXeK2uK+YGg++OGro0RnBJBYMl2gepIib7
p4Hd4eoALlDdTTGkGRBDzXGdgr3ozaQVgHe5YYLFIDsvGWcqi8pTxi/JZ9C2/oo0uspV3KmMtCwH
cptxbnl3wFb475BEUfD3umMIhJubSTcskjxXJnarMKIGElY3PrV3VYkfD2fmiWh0V85Uj6TzV3T6
o5vlNxKbdbMYx+AyWDOiXUPsHxezKirH7P4dOLVGjQnEJWVyX4OjFmxsm2LVI0LmstTj3GNdFDBR
On/UBEu7G5JF6Bd56+KJPJZTQTcFiSa31clN373jhr3GBbWFCzBky3pCg0KaDcAtFoGBdlyLA08r
pR1dzqmqlMZ/CLLoVwxb497lcixs5ea3HBimfU5j9dD5UzPX1n6cbAjuEUtYNGT0wYX65OhVAfxF
12Np0N6CI16ORgrEUkKuGa6fRs+XZzziHkX2om/ad4fGONuYSIb969YAOeUhfpEkiSqJWZIrRGCa
kHbDrR3OsqVf6hYrBY8FUJYVF4Xotat3nRR+EtAGNpmQtsalhF9yjemGDh+O9pWp+vwmZJ2B3WBw
GZlqKpxwO9r/DfFfvwR/NtSy+OGZzJ31F3TFCDxXcVx4Z+pFdqylQ4JY3mAznT+RD5abwuU9NG4Q
ScoPUSf/mzM5K3qFqvyUmhafW8OVTnIST4R1EWOeeVwmxl67PgdATXi336ISW2EvcnFQMIvcpLuX
GLtb7URUpXu8RQ09DpFW7YTCAInjr1ECCAF9zr6JRb5DCwt/t3NQS7YOHsxnh5QQWmmxJR78yGlj
bDqjEMZYrKALWrHE8RhF9cY2eaZ5OSB5h85RmppYl9DGnPj2KIAwRWXufLTlVnH8CxSCsqUddqaN
uJ4GLU5Arwuu3MrDL48Jv/hYH8hnn4Pz8GMppP9GvOVL1xW5XNKRBRK5A5KuGA27Wbh4lo/lXStN
8fktZwA4udjM3+OFT+Hyz0O+dDQp0CzNBpWVHSYKGKiz5WEu5lkENR611BpPuWg7Z9YYQ/elFKR5
9HfXeoBXKgJX9dTyXuD1HUbVanlMqKCWzLhKSZvjfAHLOZQYnK3qC4zaezZQeD4s4YkX4jOx2JiN
2GFlZoMb/vPRq7cJ1ETgUwbzrH1dn35l8NuGOOJBMjeDhz3R+1zUZRjRE9oibxED7ZqY2BBSUoV4
Ai9KM900sQKebREKin9KPZTcakMkJJIxbJpcn0BKahp5k0023mqBsy8mXLkAbWkEPK6fGpf3m0hH
SOFTDHI9osOUX16+AALwd13teGSHCZQ1AygwTDb1cypEtYgV0B32ANFDD/Ab5kOcUsQKWV8p30LB
m+hkrZ2FXtCvCV6k54Ljczl5GaJVsYMaTxk5oRGKaVk1cDkg7bBMvkp3pX8PRY8n06wxRKb6uPCR
VtN/tA2SI0funnu17rz1Kvk0K0ilvKmCAGv6MDUbSUqo+D4ifIFBWGvU3j5jrnz6OFl+t0dki/Er
pTpVtv94ukknwzLFd3RByLXxMBGOh35jL574Cam4BizcmHmqB4J/zWEcp7gdGg517cuwbxN5FczP
ZohArlyy0VK0cpc7slgUscFAmUTkKJfbqPiQCgLgHjkZxZQuICso522oXGUEMZyhWWLDC4Eo7SOQ
LEJ95b63azRSYmDUkQypM78dqjXXauseufWFlR3/fYu5G84sME4YOF97cEXzXacDwh2Z34eF2EN2
teVPOv7m5vqR9GoFciBlOtlHaRy0FbC20Li/7+sqWf0gsqX/k+r4FLwOsE+aEneIeAOaotc3ltpD
Ay56oLZs31DaSRjkYHO2a7ido3V+miNxs111BribddNR9TjutfebJgaC52ShDqzg706F8ufgNtm5
nM61AAKJrWdZ2X2Mz/xHtmbSAQ3KBHJMxgPMMkEny83ztn+5pYr0VpQYVoRDHVCWI2+fiQKiDmvq
v6h7Xk5HDffgeG08MqXTnZxsN7MMvJ4egMchNU/Z0zoau9jFZ2emZsIbgaKt3PKoYEnYrVumjCBJ
AlKx4bDyuBuVNoLxczAebBelXE+6bPfOSxH2F/QN33cRqRujY9Oamnc9A617/edgGiCSL+LYJq7B
hCX4dRDv3pfMMafnJPmepPFORLoglZtHSN/I79ZRWLLWKpSRn+2bsfd/essw0UjAAyeti5sqelY8
h2lTGh/qNJMc7WByNNj7wTAE0Lm2lQY9YayrzXgbMSvAeUE5Pc+Ex3i0pxrRUieKImriQeyReIos
9HXq+Dn+jUQb/sXH1c6+/+KknOCDj3BFamcje3l9B7aW0NnyClaL9/1lRXozsDHb/5KSP2FEanvs
EWPOqZLbkC3H2jvmftPP7YOAFhg7Acwx/Da10lJhHdpriiI/NkuE9C3aBoO/dZqZyYfqSeJEmJdM
733PKRy7XUUfG5pbeO0Vyn04V+w72HuqUD24zkW9Hv89XknYJzpgawyae8eTYjGPzcSoxKipyzyf
UkhGyMcBkCALyc6IQzvPdT6Ygm0zAfsHUyYEYsL237AfTcQlWDXT095OKyEgTbDg0+cYBD0trMZM
zQ8veo6yxqCMITyQUO1/2UUNmWqlpKDrnVj6OGH3P0Z23sVzd+hWHQV5pdr4qWgv5iGNBbmDjUUS
BzzOecVfduKNM1+Lqq4GUT2WmcTNrM9Exj3kHap+hWbr7VxiSnTYT5H5FsAY6nm5+y1a3V1wX1Wn
3eBbXiaQKtgdsNl9F1iV3/KYVj7ZDpa+WaPI2NR6/XRB1wXcN1zG/gWbF6hHVK4DjUQY6R6/94zR
ZfisxMjRTCdSt9X/QvOFCezm67h9FzPpNB82v5aG6dtF1Bjtl8zNYZj5R/v3pyvdt/4D9YnOuw+h
w01mMyE9C5vC78lWA1nVnp7B13qUxT4gKHQm5Rx/kTwLKrcEpLB08PNkHyE3RtReKkMTjkBPtfi4
3cSNIaxiEtimhKx401QdBu+ZaluDZ7CVZ1C3RbSv3ObECKYOe1Ras2BGwgd2vfVLWZSa7SAF0c4K
bX/p92cTlssnpEHSgJtWkCYBD9MmWelf5rVrGRmj7OBfAY2tmd5cVltuE6+BPLnUbATRuTi0hX8o
tijOTBxYy6arP1BrxMZxEAOFw6B53FG8SFtkQemCgKlTvj0QlVA8CE+RNcKyHIsFiuQDD4zXuxc2
nw+X2xK0125qTw9ShhfaVRoHWg/J0ZNjfl6bzSL2iSZALrcCdWQ82zSIA8MHRjSoxfF8Rij2DM+w
fc5IpjsHcuiHqaxmkJmzjlERBhJC0GGoN+aRs2tdweKK1DUyQ7dpOuxQ+C+VRA9ndXjd7xUL5xXl
010SZqTZkI5m7VP/sPmwPO25+Vqqv9rhx5rHiU3fB9WG9a80UmenJR2ejuUBoXXjkmZdgc2AwGIt
dcsyEBSRWeyOURfipjqCJq69jUuBBiG8wR0rwWTuazcmf3VXueUHvlPbFDwQHMip0ChvV/X/mx0e
ZZrKgkLxb4zDksH1gR99fKtfjChse6wgb6BL3g6r3gxk/DQPtdns3GVKn+jUETjsajPd4qzWaLqi
W69aH0naFOetILoWKQp0CNg0VJ1yVRloIYgQHzeVNRopjOG/ABFS7oadXrWylHeH+ZxFC3nf32Vi
4TAX+BHAa5Ero9qkgIcVlaax3EnWd1sEdag+bJzvKEiw0n/X5Q/MSUha3mj1B4qkAoCrZzUmyQVc
8OlZmzTtXDTcorImViIldlHKthcBcd15PyXG/lwU7HOQ0Mf8ymh1lxqXMj53otRJCB3D9vBLZpEf
hlD+zLGDbOZ/VqE7oEivYjNhLaaHDv2Cc9+FbDh4cUxy8MXsf1M2kOnf1v4ryWKE6OyToVgb9gcP
t5qJyVDtTagt3ZLLkK8NEufHlYYHmH1TQ3bxR1ZZgFTYfaecqMldQnaMCED7mPbZrGw3aczpG4bE
RH1S38I580jh96rg3dI+RHd1v07ADh4y1cxlw5YDwaPHQ4/7/SBGjVe99ieAtw1eQzQDH2pc0DyK
+9Nrh4gdnSSQhDbp1/kKx662VOKJ8VeaEYTAsJ3nyYI9VBMQcrYDikL1paAoLS7yx5RSumevFeyj
HxWrXtBwu6u2yyT5IDONIMvamDVt6gSeoAu1Xc2BKrMnuMg1qSS/W/1dbD9WSQZdbGu/yind1NdX
CcQyvp7Dz2W2CbKDfi8YL9IIRD7VBcIl1QPXSh+DMc7IoAsresMU7pE+pjzlu4X1Jle4J+Udkb34
LOatBILfyciVP72nqdk7t3ia+mNB1uMwXXI2ti7gK+WKgLDVDh08SA1culroiedFqfySOBItQKO7
/OCrFXK8KfJAPKZbw8dPPN9Fdkem/ZGcvb3sTNtzOKnYSv9yaX5PyDPU5dJgo/Cc91cq8EUS/thb
IHEs5H+ytono21v3eG5YviddVnoPnJBUhyx7+58Sm3oTW6jc6Cd/LeuQ0Ew+NMuT8ZMkibsqFrm1
XhLTxxPckqo18xho/gSitSSncazPuv6qwJitdj2wUuEhQqG0Nue1E2f5a8YlVE0AzIMQOewbV6S3
iZwfzMNcchszLBuwGEt4VZti5/XYl0xDP5zPBg7clHlv4Q8fmak4psLnsQU5+IzIsldWTt8c0zCa
gndLtX/Q+aF8LOMGK2PnXXzQJgvXLiLEnbbXbOhEKZ02oOXAgBtfiCwTZetJw4WZ9mcw2bN/R8tF
825ZwHB7y3S4OjkPttzHLNBNdGESd0DuCa2piKy5bXQ+VNLZfEApcdL4Ea3CAFvwHOyF247SwrKa
c8H8SgUBYDoRFysAjZqyqgODstS1KxTW17Wm94olYzzJgle7yz9y2Fk0eOxXr8kVnqevADwekN/T
NAwq8aGTdMXrWizkwhgUJOEXSR6TyMOuQtBn7A3TdVcMEMkhSuq8N2Zg8KC/rwJl2zUcLZIqFy+L
fX6zKlj6aMP3d2U4b36rf0qBwG8X943PpzOgWIIt/0RL5dhJeHzMIUw0kCfub8Bsl1Bnk3bF5XSP
d1CPDF/iBT84lRr0Thtz
`pragma protect end_protected
