/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1103168)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvl1sgUFyaZsaNGfiPnsQuCLZr9DYFeDh+CfjWmTy29cSOv1k3Ce6aPCuV
G1kpBlhQlG4KUfZp/QCwwC7JOtXSD9O9GKmGJtinECH2gY0gqx8M/mKN1FtPy9zuu2GqzRB+ufqp
qeJmiSBhFo8u1WIrhKEzp1f24fy+ezi2EAfOCwGM1E3YrfAhKVtPzT+DVqb79PkENIvnKWD6T18T
q2P2CjTYM55NurO6m8Xt9tMO8AFUHZTcLwVCH2iQgUQQKu15QqQ1m54+55G3QN069n2GMXIVdHGn
RjQLKh0e82k9VGa8KO1dtU5kqJsoPcNgXjpCNyd/fzs3DuSGltqltG7n6HnzMDC8ZsVhm8Pt3Dgz
ifWYCny30x71E4emt54IJnUY9F65EUjYwzsBzZmztDTbo8e+sz4qZuwMiMclwuXugjLixaeuO/mT
Lo+TIfLt/55VtCFXcp91zKB6KNti611MylRS7g/X5rkFOgLUk5+h0TmjsB1EatedUEI6Vk7/2ID3
wiIUG1nE3gDRtXyUehvEJBFPXVqeRk3ILHS4ZXMSdcIT4+ybOHn1b5D7x+xqFhOFSt02cso9sngB
8w5JMJWJaOsiaaQBwaLWAujZnAFmagOWPCewQyXayJEvMK5zzKCWTB0joghroB5R6l9FJCmUQ7zj
+OMD59/0IQJItNPjgswnn8MK5V32b/bRYfdkNnms5riNDHjRJ9vQC3I0qiilZ8diYRfU+TRrUUa7
FXexB9ZfY+6Zxuji6HNxa0YFQB0pNA2Nhwyvx8MncGtQ+SKPQOzciBC+kd9LuSpxTZqkRmRAdALF
0FmaQAd6kmnoo+6gOHHxySfQkIbGAtQyMOfEl1PExMFCqZo2J1qXByj9UgtkpMRyZlERR15/5pUT
c4pSaQyAXdl86izc9uTzzBs6crNtBVOKKDnJFi0x00iLpa9zkAfMwEcJwpjj7Wpbez4eVOJqavGO
aKsWDnxdjGrCPhCEHzIseBVR6r/STCO07DhKoPa7lWw1yoz+xBFa0dHA89+01m9mJQcTeFiq3D8A
m0GaXv7x374hVGs5Jj8IajB7ceqjrX2Tl24AVduuNQut2EyBv72/RFn0xXiE8y4Csa+vJMPgT0Ao
eIf/1JOuLVVdAnsJlO4d7t5gLe59cDh2jwdKTDlS+UAuvB00jIyVTT7VXQP5uQB/mUizyENYrliQ
xaPPYkbuc3RisKt0Rm5k5hPZHelNeFTXZKjlAKmlAWlJBdyzrX79vnwMh9fMooJ2INixdSud9ovB
rXA2yI5ZFMwZDk+ApmftdkvSfInin4XNGVkDNBp/oArcLmbs/mQwUZo7N0eB0U7RpieyzI1W1L2x
HcGDSQim9kvMhnEpTj8r2/2ejE2X4v0T1OLBz1w0UQgGh9dqxEP7fn4ltqvcqEyMPY1Nprlrk7YK
xqvvdBhvycvoE/9PxmA42M9dJWzEGmj1cN/87M0nJDD99IzNqt/S9n2yy6/KZ65QMUeACLyzxLyI
2tlz4tKkAmbFE1NAO1vF5+sOPHjDPIe7kZDXNo57+E2ZZkR0oHrZzzM0TVlljLg/p4Qa3SuoSgdj
uKfsiKI4pWr5M947qnz3AfsBORsvS+TQKI1N4IvYMHDIWwVtwpsJSTLBSu3bG+LG04rsZ543g9Xc
o4MUGqRATl3ifa/kh609LNNAhcFTjePlBa9UcGqChdJQDdnDHCWlBb5VVdABIi+Aq8zpFW4L1nAK
IKBrwq9xPhHI6tplPUk+g1AyOCfH8ORd4RPENg+k0n0Oa4wCqUmBq5ZXmu/XoNnTLmRmuA+uTQ8F
8SFR8jn0e6mnQJn6MchU2RGj/B6mqwq5KIFi5NUvWDjFj/7S9W60FXlmN139y6XuEQoI7KSixYdq
/Z4xYK1BfKQTIEXiRzs3bCqZHeTOyHPkfn0Am4p73YYNnIKX69nOBQddZ/cHAqb3lM82EfH2n7pH
vTkyR05VuvtPvMKaw65dTigWet7e2FiY4BqxVWqIN9CgURVn/PmFGDE/kDJ8TnV4j6j82okKPY6x
R2wqxZ7D6gPlGJaEL7JNH0fsA/nihpfxgIGt03HWg741+3+4ltlsUWIrPhbrVBypgKNT3CaX8fuB
tSjWNc0hoUWhZytzE0dvSIGMHIxdUUaYayTwoYsV2QW/FH4kNPSvbM4VpeYcFgYrovx0047koSDc
EYm/Hz/mFgcC0vvwXxdyRvKG1H5hT7u/3xCsY9hpUHVKzaYGC1q9BW0nYR8Ip+7BTHyieCCloRTg
6rJzPUHJq0KVXH4YT6GXjWy4D8lbMqRvaN64gKPCkTMJL/FnEfYG9Yo4aABIzdsKX9xmn3j3OE1U
OZV70UU3e8BP0IiXBs7vS8ibaUupBh18xTDhz6F+LriRXgDDVN2HNvOtdY8MgUvSuDODgWkPclTG
OC6f3/tVxnWSgJs1Dyryf9WtlpcMiHDwk4vRVlWOaMLxEKgu0QUIpM4DViijXAtGo085EaZ2HMOC
uj3jRpDi03shYomzVQ1WYPmIJYHVpHOIRJPKzrD2/nYCr6/HKYlWEkGdzrpnHVyEupMJkOxmsBRw
u8QW7nLuGR43eQ4vwp51cq10lwWnj+GI2YzAgZD7WzX99t2Ma0NK+CLX+X1zF7xRER5iLILux43q
KfyIrwL97ZuP9fchQnw/pecb+IMzIirw8CLhM7Dq9pd1OTZTkxpoN6DLd+JWqgIof+a1RsrX6R6u
tY1V4isAkh0AisUGFTldvcnGMt66VCcLbHbf2vIDGfVZbOCXW2CQxPDRIttgFXkk8zk2uYbhMLjN
7dEm3UPyLF5DnViqipa+8x+HyQpGvKKxzLgwFcsFp0BEL/uujKAJPEjfsmdXuSLyKByzMrSzNDCw
o+cF/aIjhbOHUciu+UFol+uQicnNwwyrGbiUyaoytydkFb2xAJ2hHmtpQPkfhY1wLZiQzcviQJO2
WgPSMf/sf8e7KoWzgTtwxnjg3Jnj0uaRXzDw9Pkj3SeXAztZecz+n4vkbRbDx2wjtccMEHDHfKDO
2ugx0SysnMKBZrSG/uunxTupLUaO3TODuvvRG+psWE/wZogd1UD5PHnjEajYMtyTtaGVUWOc1IbX
o813GQMrtCLWz6s5qQnqfuQsFpCt4dtSS+EMLnz8gqEaBziWvfz5+H0cf3eieCnAZs5GK1jCSkmt
fP8io7g0AtdfPLDS+MWt4k4t4Qq4EWRReMy9Ozaotp/Yy/3CDGiP3aG2xnfFP5E9Cf9HkSTUdugT
no9fKck/nySGsSJ4pUeAgpS6Pb4fgAvdojoFDQai+7MjGrVgJk9r3rMZJ3AxyCVyESnE/F8WgTDf
oX2q4iB0xW5gbqs2205Oig/OA7oCk/m9sFCQFxZR6dXIQq7ZbBTbPGxHqk+HL9ebPz8p/8Y/q8JQ
L6stoZ9pTZ072IKm8QZHIs2/Q8DqE2YqPJ01iWXNggIHNn3ptgYS0vWNN4j3RCKBsxMh271bZAzf
i9feJe9WZ45ty2UINOx3XEbFKQ8CG+jpIy3WpIai4Fo9sn1b40O3blcKaNyyaqr1DmgZ5OjKd8p1
DlPJdzHMPFiq9fY1iOyHp33psQdw/AafwGYy/X1uWUKkud9ZVg0purIMMziqblmT1/rZnvLv3xKb
5DFHjMPyF+hIeo5B8LZducs2leflAn1Xb25/Djx4TyZYwC5n2b8yAwhCO2Q7+inBUs/jC0vz0/TH
6rYit5EZ61eRi0hE+lNf0fH/XB8Tuk2FtUHP9Bgbj4conDDQ3SxSqEGY0u3U1l66UV6AqsmMXu4q
h1lZQl3TB0U5CesRfCWfi3rOpLU/+iw64nJ0l7IiMQJ3OLfwQ2CaxgrQnnz5uVcRF3cWJm8iUrOA
nk/efL9uot0oZcd05tXUCkGj6Qm4QTswiWHt4sxjE+xvzlU8wGToDVV9LQa5i4girzRompXJK2f+
2gYAVLtloo57UTqCLPgRCkXeIY3A7OD6NoUfhXDxaZ5/IUk/cAAETF9YyEh1YntJcI9IY/svV8yM
Yx1S06+CcxCiYophpq+kYBD3s+6NJMOE+P0WzVmRJkVRwPz7OwkoOXK/6mvrm3R5g9+snQ0ITRiS
HA/v2lKHPXUsXp2tjOM2eIXkKeDVP97A/nJFmCMYlaFY1IicHKm2FnVk+O4QfecZAeo7PBAAVSLQ
WhVL6DbAO7Y5w+97uPoDyzR+/UWqmBlOpT49DTA83CVfTL1UEHpfcqN1faD7psifaij55MGwjzoA
yPxBetu5PxMBrQh9roIYQm4GjUfJuw4Toj72b+aglOi91FtDkIN8n7ZC/yCx4htTYQ37v/nYDO0P
b/8gTF6b0He9kcI+0oHdDbcy/oY9doaPT9Xlk8UIwWDsWHtuPvnWbduir42xCOPcthCxzvpzeksx
7moWeNdpnVDrmWP9InB0wSLbTz4Tlv2s8hxVUZ/lVnSVqg+JnWuFlnYwU5ZCfhOPGqJ4NrLTgZSw
81k4HIXtK/Pt1rged9/+6ju5nz1UYV1l/5OjLKXOaTF4802jLzZ6P2L1UaZtjXeuwaECRmvIdVdK
j+35xd+7S5dHKP+UZPAb9r4GM4n9ew81peLkYxAo0Bkev96bgig5jcP7mZjuz4egvVnKGXvBPsxU
Ny6+rDbTX8ltBc1th6a7aqAAft+FLxzk7z8w+REDUh0wCz1c1agZq/I338wQKWNtywI6PdgZSjY0
YBbPtjREIv0olsR2d8YSMnisjbJBs198J6KigbBtMWPiOaEJuGtaFkhgdBQuCQzHNylEFHDxiPPt
kzVStJG1r/HVR9hU0PuCwi3MM6hMb2HTZb7I769LChKV772kRyVo15QYm6HhUtbb0jM84AtBldvW
lMIGsczuhwVQOB9KCeHOi9sRXvlNsNAC6HZcABTtRyt4VaYWGnJC8dSokx+kwZEMhU3fJqfvFE76
zmjyAD3tmFKAj/jKVlLr7CBCNQdHEEfv/+NKfW1DuKmvYEvl9gQOYiqdWijXCh8+GlpczjVrOtUT
C/D0E/PPBCNV/8Wh9Y3VZcUZpjnCs03eBjgm3zORjpwuCucxE+vQJLpJqWF781pWqFRkQN3jTh35
RDtaTOaPhTUhvyiLYeBUsP9K343NZFiT9XtCfAHrE8Dpztf0XKOViraWMeTzg1QC7nwe9rlzH/ro
M4+qaWiw0WY4ohvh6w8kB8xOQiIqQZ5f3rYfbJ5vnPiDHTva9DVpUj+8PBhnG5Lbd4ynYyWCtYAD
HzxUdCaAGnMLkCndFuY7Abmb8QKtGcVk5/xUADuo84C5b5Ex5aJm1Fyl+4ysd7NyClkFacMy99L7
ONapzZ6LFZbPlOnYZHdizEPIHtfBTi3DU4xSAe99UMjXugCX/fjZQRdYKOHkB/seOpziRqSvh2pp
r30XXBZV96PI99LLfb7onl/zW6MPGC1gtkizTOHKMV2Gwdc/9TbnxBnCkILDyQnVn8c7PBS3eXhx
AuacXytcMiJaLgOwEQDTAactsSdymX4FOVn0mxYik403Zf9oMDMInNYX73O9OwAsaaP/swnBJOGH
Nx3F9aBrNCPtnfxgi6+dje0oE/sURLcog2xG+x74msHaJiJ1X2/+RuzeK1+UKoO737ojW3BgtD/2
Udpyg5G5D88nDhF6SeKLpKv8ZPMsfnt7nr5t7P0iojm1f3CuV8prqrj8ijrMfCGCBdJmlRxf8Zv8
Pf2oTg+lECLtvXm+vZRGYy8HoM737aI0+sq2AnqrqsEuIXj8xFTsWbSeLLO+ij/HNUmbW/dRmxZ5
j9LKTs8k8roKf1KUz6j9bXWk384YaIgqk31roVR9XtviG6APuXN7hSBMXtd3zvk1sOf4R8mnWQUH
Tr8UBWJzKrA4q2WBMusW1QQ4wMMp1c+G5oKonfXvnhb2qPCW6aPTl322qgRbfLOlg7uK6pPLhwBa
rMqiao+Z1GtrloRl6uNUKgAY7KYlmZ4xm9uHDqPHmYe5bTj8DmNNaNKSO/+zpcRvA4GIWwG0Od2Q
2OUGqZLOW9p2d5UZkRh2VjwOsDwzguDaj1/hnSYf3ctRYSyAezVUhBxxnzwTOLBJlZsh9EDKuqEL
M7EuxkkJXWW9YVw1aFc0YPjimWDgOtjpQhIj/EJ5I0ELwjgDZraUn8fqy1Pff2dos50RLNtbjHOr
vrlSNVxCHRs0FP5oHnhBNIx+c+qysBcnnBUourt/5JrVAzNhocb7Ec2WtKf0/vdaYfOii/sKMZyw
TwfPn0o5erEIiXf89fBVypbflQYnJN409eJIyuNSe8Tuz3oGD+kRt51jfsP6jvAjovHIbLMoLtto
irLtCMgYCsWgycshhfcpFhO7RymAhFBejVWyHuSIcwjvkx1LzURsETIEVhJtMKMBTtcJ4MRN8F2Q
2GFS5l/9KwsOHFZrPd+iakZPV3N5I4EyQbu0NN+BuWkopIytTcGzV6yAX3dzMX2X6h+HktJe3bCg
sp2rRIMIUDkOhPe9Ov0/xMc8vvUqbAlIlfaVpPsYl8G6IqnmajdyBTjcN5Wj6Agm9njLkDhQrad+
2rgKu0wv9ng2LQfBSZ4VRzzNNKTuRYMuh1IVtnVgoPC4ayUKp2n5cCFtwGbANfUUHbdyqy9ITE52
be1BvpqTOgg5M6Xbp5RaFvQggS4rl+xRVg4UrDkkBINQiwM5i/UioRs24dHJ+7NcgShhwS7AiPRF
xDmgJxaRXtIhD8XaeNhXy5i1RCCpfgajDm0YMNfSqM1/5issovdIZ/kMSW9iIcJRl9WhEpZVlUvk
5zjWn9hq8EcfIzikpMDHKb4VQ89tNKoG/uaMnP9x3P3TKrOYuTwlu4plTqPGst7xRdJJEMGECH9j
/LWG8oK6BZYfplZZIZzPPWsTKtYNW4AoFS3lhJ+Vb0mkMdDsvK9ZZ5GAV7trq5JNmnd+h2XnOnr6
8ox9g6IjbHHO4sHm80x2UHXtKrpozCOcJ4ldOiLdxqai5Y4vXCUQYwib496oZQp9rsBues7jqPYD
ZW8pItLFGxJXK67T9JEBkXsuYCQtTTo0kc+mpmeaXOirTKdygIEGBvoaaizwBiNZ2HvXHrAJPQ8T
cTaR7yXLoKKIeBGRAbi2UeiWsc6ERx7YwogQut7Dfd5BIiHtvuPEKcbLAPcwdDswX9GQwZya751q
YELXtW33LiH7E3HWwcj8lRs6jNHXwj5cTy+djyYfdCWLVzqmsGmkigaITcoguS9+LjnvSIUsymTc
wbHpj0yM8YfFEIHFUwSrXdEhPWkg3W9ve7qxmI22OC8zZdi8Ek74+Vhqc17LliTvpRoZIqIN3V3I
ZeSBwX+O23VQErFcusYxYx+ewpYLuEC9K+IqC6S3ZJxYwkZsabO7bmLHp2U6lLDzNQ7hYff2hm6K
WOGZ1M/Jj31dHiiC7HXvEHzj4cxGvqS0GvZUFh751d0YoRNQqN/V74ysVvWOJUvgUFbttXa3z4Xh
imrV7CAz64kwDFxjhnJTlpE09iqkRcR7BnWaKSH1bSOJP0G/g7AFaBRJZ2NAdCVYhFezTFtAHdLy
ru9/6MOKvfxrX3LCn6NHQZjH3kGmZg3eryIQNckmdmDCiHPTMrOy0N7aiufzsCuT7ZXeFK5YCqFv
VbKawwo0s1mrl3uc8Zu54HU0gi1UxegsmYn1IiY/GUdRAcnUZeXgLcPb2zNhnmeWsSHh8fw/eamX
oUfgHBMvN0Pj6YDlbqY8M/rlZ4lAaQF1dOQ+r3wbdIK+GF2FjFR/Inw3aX9T+I4FgTV8/yggLdFF
gp38eW2LLd4GKA0sF5NI7+EFfxVdjZAyb/nAhamYxgel1hpVYgZ46juYIfEE7HSVQWAmf4AkBuBU
qbtF8zRhgmKXB86Xsw/1b2+efiTfTx0iW5drf3uRyqpfACTHPCg38l7YApFa92sE5WZDxUeMnw5T
n1/hu/0R9UQKTfRTXgwPWnegpLLVoxTcB/PX3Qp9OydqFkrH3D8pDX99/KqjsiMulPEdW8H72PS7
dGST/X5A+Ym/CZrb4HRsR1ueds6W/dLCASzKwfbXX+ntiYZGoV1GTk1DdUkJnJc0X3OuX5CYBWDX
2BvtTaMjcygYiBMfeJTEdllhX3/69CnFpjjs25XafPsrMWeP7mzUkITRusnlEkVkRxvTp75+ypKf
HBDqlrYBSeAJXFshdnt1upCZSvj/2shPVLaSAQnchp0gAfbKeX8LNMdtx9MyzOo1G8OhO4QvtfYt
+W9Uji4oA6j3U3s2CGbX3WqiUe6y6zyLKzcv7roAhpf6Tu+6ujXwW5yw80HB2iCjL/g/xYnBzgwg
u2BBF0Rodpspj6Ey1fAgvAWuoh50R1wmDzH50mRGV2zrUm7dCoD2TF65DL7tTtyzCBK4+v0GC5Sd
QYA+Wdm7PMae12gmb65Q0FBXjPzfQTnpfAonunVMaPYMgFghwJdQRmYl2DxbvED1dTyqb4Ps2d+e
VawhvCHaejR/P8SVrd9lFgCuGqURdUtms1dtSyG5Yo0evYI5Chh9C8MQSKyF3YtmenCbDZ0WBZzk
YC8HPyty++7Q69Tuv5Lkkp6w7gSodW3CRDctr9x0eRqI/EbmblVGTibVFWMZaost37OzDSS/kNlw
87hviKIlPCt1JONandj3G0L6092+JsqKrgM1Fh4MK1DJ+LrYxvGXDg7X/a0V5ZPnu38SjA2JDIAz
ZpB3bXlMyjlGKKdLndioYlfqSxaqg09lpYanTGPKUFchkGkTSjxLQcgGUXQeXdVy5vOexWBQGtjg
T1uStJCy7AUYY6wpiSjL9PaeDtTo4y0GgY0eKX1dTWWM7F3DxfWBOLap2tMRlhMSJEOYHtzmTZ0P
CbnMocIFB6QJNOhORaRR+LV8MK6ZH31DmNl8Fp1U5eJSIKksQnR43JUMq7j8/aEGs+2sPvX1yrxO
Ywf1O2FxIjy/vtnYD+nBiJ/O6RZew+OSClmIN4YWYnphcU5F48RptT6HNTs2PlPtBd9HqpF2iYhV
vJRtMtrILXJ0l+W17y4JCatFR9KgSKGqa4sMSndO0WJztXvxuKTx/P5JoFcKAw21kdSr2+CcoVb/
T5pbaxwgvDs2FzzdSf1ZoKrhJOpL0YdPgcUlZKIYKbT3G1oP//prg0lfd8t3RzzIil2DJbLAknFP
jpqMnWbyZmAupqKPbedfvbtuAudGo2euElNt5X4ZkhrWVl4pJ+hotreHqeLfjPJu7dWptyrvGwcO
97xCWYH9L0askQc1QfyeTFwc734xCfvMWJ3j8aQg4CvQ3HQVaUmhoV2pj+8/toFmKIHTfq4qb8tU
78ifkhv1oOrRNWC4965uBBMDREOTxO0q3zErhsrX9XgVOc2WTjT3RN/974rx8TzxVHY88kJ1soow
8GXdQfK+l4VAYVGQNwSY5TLONdLY232aFEeNDwwgOY25QABUHmMjigOctV0B63iw8dhAzmI5ioaw
74hMHmcLrKm574yT/gloeF1jJrnZTKHErGukznvjfyiSp7bdqVm8/kxFWswef0nqjrHHOtIVj7fJ
PANzKV6x6ySNIuqYVBJpYCdX2v7wiAkqXH4BbFbn7+B57N9vWXiqZEMr93s7t/EGujuroT5D0ART
kfKKoDnsNTni/vIajfu2jAnB0OIjnclxQQCutn6+X+raLU8YOONkQLyCnopCgSsh6yW+VYCXwAo+
JksIzgaq+ff4cTjtwj2LWy2NtBNXgoQxPnPqje/5sleaCUtz+vrnKIKJbTj893BYEmjDqAnfyt9V
aKYzaz0FjAnjkpIWgcbT2gGBM+lGzzdkyDearLEmwkf3zi2NVKPXxaVaHZGmhyJDb5P3iemAKaW5
qRcnSUzKvGLGeDAOByIViKcZgGSI7WGdfHWMqELhhRHRj4DlIm7ujzPLEfKsMgIJqJC8qx7rG3wG
kaJwILpkccl1Fv+J4edDvGdXEx+So8GnBQzw67K7JJLLr9gmpnVSnDv5J1Ws9+d4lob8Rpe+uISI
XXDe1+RiVeltGNxjYJCUSm8Cu2eOdoaUF9kTNY4yK863kOmHWB2v5WZNhHeDXT3ddhkJDgziGmLs
9m+n7B2t0P2Ad/Qr1ulQK+/p+RpElFJJiZgtFLDoGEGvJJKUynDliB8/r5CkmFtRG65ILpwBo9hO
fMWoa+SN+Q622lDQTuOlsYTBcFA5Gt5/ssGpXFonVLCW5zK6N6ZwLNIfSok2nEZzzIgYKKZZlsH/
CQQ/oC6iu/Tzehnu2xfEXqUoEAZ6M97vWcngEPkFwj8Sw9NKmo0Nqy7OtnzrVqG/bE5jWqtSJVVk
VJgr517tJEce7DM6sme5SOk/4A4qQJJAhIlP+flmQ3L7ULOEwArtDAjmq3G9pn/wZWiuSzw2qP3G
jSsPc3X/218dpGQEX0AQxUrQ8r//5HU4ioANew8bWzwUy9tcX6WcKccfoosy9XeUp92oq1pDEb6u
DX0JcRjzz0jXBhI5b/hRkz+EwIWbg25EkfO4yYyAZxe3NwU7wgeit9uW8pC1ITBtPKoaW7WUYm71
3xFtsjHWeW8EiUYr+KTSMO8esNX2Tkgr3mBpd8x1qJ5bL7/uW0aENDjw4nMU4xfjThTHXbedYk1i
/59IEn6vLGXVTVutULi0yDfpVhM8CvBgqhcsYlw0vK6QD35WWPspc29GVwrsxy67D+lbI8eRzf2b
Ui1hZFMz4aZMx2oTydS1WU37mfu3MKbMNPcl0IlLJczPAhuMzcQ5Qukk4ATN1qCj1zzEFIv6QI3D
XxBQAA5jGojPf0EsLbg37o1ta9WS8jUzm/o4AuwcDb78FU2OHp9/BVE6RbGfpAK7kalWX3qB7Ury
vsFqHE/WU9/LKjuOGYuU5mykrfk5OPzbV4EMoeZMTmaGzpLsGk7a8uSUyyKCG0gBIOqAdyBRm983
tyvK43cr698bo1TbNWsOep98y9+VnArzsWeZHi9EsfjQeoNwJj/AfGiLH+NoB4A1XWN7FnXjED1/
01ngILf38EQ2UZuG6mr7z3gz3gWKa/OaExS9f/wc2/jGb2OtoYo4ZHMZyeGCGOAR6yMKfUAKYB8Y
kthmhRgEfrPOZ+lT/JrOXlgBAGBpsfGNlFopp4+UeuZYrX7PWGHUTZr4zMfjVwWj3fnIIU+mnaoO
vxaYHjbFjGnlhveGohBMfgjNcg9205TyGAgK2Xl4N9N0oGYzH7ygJfAzGNYfyUBpsW8Pf9yNwBJ5
FiU0uXgotzblsu2ll1VuKR/g+zs9/l3qkQoRuAhKIQla4StzzB+uhwtBhPZktSCoTgAatN57rnVb
Ftv4Mmg6AZGGAgwQ1MtckjvEZCKUGqIBS3RLSYnZPlic3clU2plN8n59JrcAdsqRty63yCjj8XcH
WplifPyR5DGcWBunO+xhPpHbVPQanLA6n12Bmh2Qe/r48SZ8NvdOen7MdSb4D+ByJ9zSS5XHlFsF
HmmeaQa0XI7NVbvxZjS8pCq+rDHR3zhhfvA4bsGXKoU1zOgcNTJopiHw5zVj8X/Z7dvqGWUCVyLS
ZzbofiJ3KA0VTKaCGHYJNiI/m/91HWo/t8sZ6LXiSlvW07z4XrMtjRq4CA23YE9Np6hriXIEsT6E
hZzBKt9I/VPpTFC/2CoBBEMhihsEzIJmEBRmOLETN2HTk4vr+LS7evUXLez7yg5n8hvGBMOhVsfD
oCL/5cMnVmpL+7Wouk/3Y3mTwIkUALL3yQrrIJOk7ZQlqrjhWRlDiVo2BFA7FcNOEU/yrvUu9s4W
VWyvXESN86cf/fUcRzIoAmTq7SwUugLbdpYwIfKpjfFYb/2Uuzs6mKzs4Lb6+gmIxeGKYyn19/mr
PnbUUaXsYFyrJQz7NTlTpbjjYQzLTxlT9/tSHLnEiEIn/ygu8zBP0xsMMQPK9zj5zdeuy2gAVxfX
wIfihsYjsbZ24SDntZUIbJWWiowyrKwPGAyvOms/XP0Pcxkz6ze79LdtEtAkdJ/gxPIf467/Tha8
FCUFf76Ii3QVpto3iyKhFdG+SOM7wmMAb6D55gfblVLiDnDAZ0W1CLK9gNJM/d+fRCUgMaj7xX4e
pl8xyWNPLPXHUdizxUxexNDhJORn7f69JMnh2KuRzJK9UGclXLUYSYqrbJ3nVM6OtPflh1n6wcaB
78zzGsS0Z6YYgAI4V1Rzna8Hsqd+3itWNGx85pG0iCTbDDGOc5YRTyRtoEqP9zWghtby8PHu1wqW
xbbgjOH+cA8gUwTxbEeuIF7kmIMvPyVgUhsdijPrhy8kPZZNF4fVm8ZOJiNm7CCoWWoCYB2sbja/
Cx3kWuWRT2sWIb5B6EodkLoQGYrTRYAP7tA90ZgFTZj//qA58BWNKmoKm5iGHlFd4qTLg/4P+bZv
tkAvmRDWbei5VofNX8+/YTo8/CViiSAtSNlkgDyYW9T1lrPCwTDQi7C/oX9992DL3PKvKEy8CVz2
eegXPf1imlFCksViz4DyWyp2flBtF7P1F/10TNEQfgNRyh/c7C6LRpFaFZ5efOd/NrCRZCfnIuTi
oNGsWbJykbSmbcylZs4VXw3SxZlwbNeu+VSa0bxNj67UIVcXzz0txoq3538wf8M9JBhsiWOW3sZ8
/gKUzhI2DOsDeUxy2GGHA+gKzcytGOBwpCz/2III7jdIhoaa+aHYkQH2j8E7C6ErAF/iLfU+TTnS
ORWy10JOISP/ZfaFY+7QjH8ufhJRG/IjEj9RsxPC9y8Yo7mccbLs/yBNmBnHnGkMD5HWzxnOd1lZ
TOWfELsetX4nLKA8e1EB6k9l2ySuEJWtBknJjyVFkqeK70wLkCxhA5nwlsuq0WsdiHKkTQMzMXtB
QzZUKzGyOmWX6QcDe5rqX6GtJsNEB81nViMMrC9PC4JUYUgC4XE6RukGyZY8QDPlX0vBS3+NfjCp
XFIqRlZlFulIET/E6oT2jt57IJAv7y3pYfKWTbhQyjuD44FYmSqDCfGYX4EPcOkNoBnExQgnkvHr
8o04TMOGreFW0bE3Shv6gIih15OkEndh4yYYVIFachSQpUOpKu7IDQxhv9ZaofvodduaqBht4VMr
tBvRFytgiTSMH65fCq9h99JVLgseTSbD6o4e9I1VcI/ljTj0vYaB+A94neNDjvSrsJP9XBHJqayq
5/5XPIXIJS9Tv9Jqyp9atsyiH5O7CdLKH0cwkFEe5EhG6kna3VgjJu/F6Pz3+bTls4LRIlCRhenz
LauDqNTnDtuQSBsZ2qCIu9qXooYzINtQQpX98yGDMYDnZFSvjqYznQFaCho4cno8i2K9nIgrnKvk
cyEQa2y2v57UShwY2hT2bpw50d+/CDITdB1PniRmR1zYyzwhgWg68Nwl/8U2c9CWm2eqnOrFvBKr
TjkUb+YqYGR9wocSG8cTxMsYudk47IQ96kQEXbo2vwerwKTedFiFD7VFOV9oZ4yyL7kbKmhyDKFD
hiXw8KPXFKTE9c7+J0TOMc4ZraGAsPYitNmDMf/G+nQ9/p8rchhPCSKDJy16mEsXtaDcp1RO1LvC
Ha5jaa6JsEeKNMCo7K6ysSxDX/Nxm2VmBS0gn74CvbxIaQYGhJ4rvuC1ak8qJJgpWs8i2srFko6J
Wsbe7ldI7uOxQUO2ZnRe0HyT5n8/LTf9eRtwz+0rK5IRimvpYAHb7fstBP4iGoO7VU7+whd9bis0
/g8qq8/W80a5OqkfrGdXPVXu05Mjf4/UdZDHtHq9sMOtYtElOtAE1vOog+HV4P3ymNHPF6jPo8qk
M16chnzlzgu18Ygo/MeDUwOCDRnwW8JmUU8sM9xDc+tkTvmI97w3E7JnvMKs7Bd87wpXCy9Kzbwn
gGldVb+fCtjWYRNFNXal8tUF2m984IhokKs+nQzuK4I6RlMT6+1EWe7bGQY9kV5wRYA1d8V1SwVa
9JFWJBGmETmpsc/DFXs3AVJ3xbw0MbgLd7afXiMrdWN+JJt78EJB1Ybumj94gzZhiiTTOG6tbj2z
QvFw+gKdnHvOYYJpO20I4lislX3BOF68r+lSaRkOsASlZvTTHoqgJlW16QO/g3KrmawOqMqD1urq
G/yBaiUlgceaewEGQnL2MLS4GOUSxFs6MsmgUunBX/TyaXLUG5Xq0XnYNRRF7z01X3VX5Uxuyvyg
i7kAl95Cxq50KaVHmyu7+W5QpkH8BB6RHLqAVfrbFJiNDG+l3zMyzzNx1tI/TW923jHDZjd25LJ7
P3c1vL96VraqKeSgpT6C5Ywk8DrIHshBOTf1WL50Gqq46ujeMM8kauJb9IWnyBpnIUaF+d7KOjC0
2/dldE3JH7ZVBdT9bB2uuthyPtjSBV+MIllfFW73GhyTcD/Zl8ucGaXyzfB05bbqL76PBeEmT0VT
UPrFbQpGpYiWGwA1mScj/6XLbrAbmT/40vCZm11zB4U26TPOwX0cUbX5gaGqRtGdSGpjVjxa8VT9
uPu3imRWQIQCBSFoPmpA/SIt/9pyG1lrSxh5qCC0Om2xnJSXUo7gcjF4BpfPmDBzuGhWLzwoDajL
mZYG+PAOtXYk85WjWfFEHuX2rGV0dy9EPuuBqXGqV+CFvft1sTQcKhL3iO43MIpn8ltDb8EOcgqt
UMK1TmdJWLFhQ2ZMTPxidOLMRsUiFHbhqYwRCjgE3Kj4WELhK5jgQOsCB9uGlZMd3QiR7VUnJdHe
yeVdeXGU0WjqrtifUHqKpsS4NK5kMxdbFUQgc29kGiSLg/tN7M6R0hMVe7NYXyD75FLm2KgCtn48
4zRUOtWwYdUdRP2/4kSeHXTUDD8HpmZgEBDl17EO75IMT79gTptxRSzcwju8qpCrC3mpokeQEDYz
0cL7+pAWnnR7NHexdPoWBTjD6cPi5haQsTNVfSNH3p9JhNcMyp/O8obxvlCwZ9w94i5iNonB+qtQ
z6P0WN28Orrs8yVDSBHwOly9+lyY/97AY8Vq/g4g2hUT//DAjureoU/IIb/gIlfxcd9xV3H4Dl/E
HaNnepJK2nKYlE1kcQvzSwE+eJty6KPxCvQbJOeoI36QCZF+4a22uJR6WaTAsoMyRJsUFovmcoRP
9qMGltBCkXd73Tf+AvnbV6HNg2lHWusOIC0L1oIfIFh2wMf6tR04oJIKWsMgKBvtbF2PdFLxmhVz
bY5Ydi9d7TO5Yr9ChZpif/RZrVz5NQW2IdmMiuA09C+36pMb6Ax7tB9pkQVkxWUB2BXI/nLeU1hw
RsFa4Hh0ZZ2c+O/mx/n54/LCpmVReVcROj6qt0rCnKllQFmC14GeMYvCmVmxXgLTfb6Cg0JV+LC6
eZbi3YOkFtvW0OB0lZI0l0IZ1N804q1pJg5UN+nKp9ZO/Geltzi0/0Y093Ijhl09i9IWrWY+z/tR
UbEqPaeLhN8rU9xJVLM/dsrwMZdTTHP/dA1e225hPPCapLbrtnGnhNAQYI0Vk6b0QC04rGecgfag
hUXEPPKmzIlC5ewuiCIN1ROkZTVe0Lvj/RSV9BxJmBzcPJ6i+wJZGftKugvRFm7MXybaamSrYiml
2rVF0xxf86U3qnipStijrSYQyrMGTrkVJ/sSluRotkaH9jUxZ50nrSE16dFif+0kcJNMqhSmjy/6
B+dTfFB6fU38eAVKH2y3IKGC+KNJgOh0bWX4KhZuLBOJZIEgG23cj+LWVm6UMirVJRnLZ42LF1iH
YyEJeemNl5y3mZhOQ9kiPUbhKeIAQ91WnesJozysGHl4NjIjTNyqZ1Pi3RbpKRqRX8HKU7Lkw9Jg
dCEN3uKBUkOwqpLnyCQzMaXCQUfv3Rw/oZ3nuksThsFnTr7ghny0HDn2M7yTyjl7MZbIybUOcyrY
30nSnHoWySk8JNnxcuWUS3p1mtntSoRHhyqtHRoanrNDE54jEe7mSd6u/jt7p9GiS+6W70QGEfS6
7idBSyOyobaA3XpFASL8+AGv3OlIX8aawy6G5eJRtYj+jXpltu/x0CSvHRvCrkhn/jL8c6lvB764
SAbCYHERKDxNqgQfNMdgqgqRvVacdcG88KmANQshRz9JCtVcBAxwvr/H8fm6kMrYIgGyGFBUZRoi
lTn1qXhiD++3xHTmBS5Mtkb1nGrXOpp8LSAEt2TC1XGzTuvbpfrwEcgUGLF3RgsiDoOGK3AskGg7
vTGWTJT/BBOqR5835642LuhjM9rRDwhqzlal8M5/nqPpgEQ8RcoQ+FDzZvH9gGXmDEICUMxUH5O9
deK4x6K3oUDyTZ3XCFKHXVJlAvBVh5b8cLA/f/wKkqEXubv/8NZwjZG0MkMtUJx8VcLwazEOIXkJ
gsGRQbZ6hMUHzQ+2P8FelrOKEZRuMMr+i2lkLRMww5hp2bzM68CfrQEimcLIgRfJ5A8wlSWIie5M
gunUMfKtQzu+UfeXFZs+6mg+ZRpkR8veF1oAhrsCRraAJ8kC7VTBbOeBHk2CC6mGkfYqjQosyyrl
nfXGBaUAYzC44AQak+ikBWTE+H9ePSdP9hx+T0dm/gsWgWJj5n6NksxjA8Au36BfGyNP7TKSR1YR
ghBaWJjawhT10F2cIBb5Ft6s2vWYRN3hE0mG+YHZiA2bxb95M1Bxyx2dw9gYwr6uLG60UmeMQSrF
n8Vjq6yXkwSI/XasuwIjvXtoSaWDniFSw+o30JBmPCGouOWODGTD8Qa+2ZjnYdkrHbsWDrXF/kzH
KPAQsEi65tnmyWoXpX6gXQcAJmQGckBonK4kVXU6lqkPrkaYV8mOB4tOc7iqOWrsjT/WACYzZ4gq
EVSZijc74Dsddy9S/kd+xr9E2x66INvxudfUON0lWGY53YUiQ7yoUxyAKdFajdDYwOcJqQuGVYFm
pRV0oaSk/kv+hrCmlyZxjj58AGTZ8/ADwOSsPpIBzR/Oncwx7dFljbtCWvjNZnrYL7NS3+n02xyF
Euw95NDpEsbSFmip5WPUv5wbIc4hn/jLqoRNR3vPzjgxJxvez+zgpY52k8hbSyeyrDOEfiIbsobn
EabSrRYBw94N4KaBEq+s1Xo5WBzaQANAtx3jKQV0P6t/sDuvPMptajxaKAbv9anUtPSHHR1q0S6E
9JEG9+3T899a8EokzuLnKhDew+YppFcIg/RTJXhcO8Y3pdG5VDp0YA+qnJ6mJznN+6HnpIA1bTEB
9CwdXnaAUxOl4i+587ESFluqj1lJSdwXXwbJgwZ7EnF7BlPs+vUkTpm4Eluw1a6xEzI2t56+QnTi
wkLIj/YJ0pUyyvGdbzxVdfpr1Rl9aZP7so0a3C/ynujm0JI3S+hlNw4EzNLkI5FZLenUmV/d2Uj6
HDKzy1joOiv1lNkFBARAmw4m118FyyZeA+Y3cwKuA0FS76X30n0uZpFGxuxeZSgrMZJzNuMuAT2p
IuN6l4V+dqEs732i4fPQ7xHa5mIuqnfJlvJKEdTlXZ5EQOjbHHWa7jTm+8V21CWix/aO6BwoMXu/
bMQxCPA3jPRoaHEOEwg3dbDdS9P+jJMWqTRCEYgS9x9hzAN3nOqfLjI/Y/aoPqY40NsiszEOIpnK
9GlbtZUdZ+/0QXfoO33+v0ejCdEFACmR6DCKum6+Zu6CMWKLNDYFSe7XrRSt3X7MXOUOa/Kfwa47
a50EzdLqP8/+x7jt/b6ymIdpJ41ImN3CM+0ETU3EiqfmoFCsQ633Ggr9kfTFfj8s5EjPXk0C9yIk
BH6JsCMVmQhn/RIxfP5bVNS9fTr8xIVDp19JBuPIA3CeLQDN7wWRyplLkXuE9a90x2xaw6tWT3Yy
a2jujWvcHYBDF7PsaF6GKqI84FZbS5hzMVPM9kRyRwv063nqRRur+UTSJPne9MoZ/YLTGS1z9zEv
egFC9v81GUtQ9CAEkRRJdhap/cr0I3d8KyIXyb5z4SvPg4SD/0mvzLRfFkQaQ25+9DfBIKCpa4kZ
WU0qlQalQlMUxDIjm9FaBH1LDbY53NlBN4u5PpDgbt96ZUUceioBYluFf4d0aITRXLF46aP0K2m7
DMWNtEIeREEqVcQSkJSPnyzOvMgBCvUKVchB+EK4a2JPgERq1hUMyIA35IH922p64B6aUVztHs9j
E0fdewjA3s0QhEaQt9dNb5xIu/8R4ATdJDyhyo0RIT4erNaZ5Ldclh4QVN2IhQZgi5FSSkpMh11+
LkFD2U0PtAO5UzqraZeGakjzfuNxqEX5FEO8E6DHUt+ScbSs6xJ5CdsXbOrdMCJKIvVTI40oapZs
+gzqD27HtlqZsyCKYaqiQ2hNaSHjfjFUdPQDbxRiabpNqz3/PnzFsFYTLPzI3CoTTDqKaaz1zL+q
rq060zw2LKLOJRdwWsr2CqsJRW9AfvjTYT1o3EpqauJL/R5G6dpx+Aq35RSusH+iUJPBPVK0e/uE
X5DmprciKEyjlSI/qNgxEP7qO+2KJLoZeumOzMEJUhIwCD608Lmvpc5hX03VGx9Oisq1AF40LLWy
E8FvR2dQsqxVqqeSre2gChLMC1FpQb//Di+/s2nOpo2ZVtVomVYT1cnfs9QTAFSFPWnt2H1nylAR
78UyScAwFsrj6I7XGDw9YQ3sm+E3Uu2kLmgm0o2f1x8ik1b5u5pV6cdlzBCBEy7xsz/edsCN3TFA
auPQJdxHMVukqGmZdTO07NcJrSH/waBGK3TDE7I9rglTKNB2SGsxwyLR9W1HiiAVp0XxhVB5cK5Q
bPn/v6yzQybAYL2UrI1yWszEj+hLq8pE0dM5GEF9nzgM2++OKSE+dA6FnVGJSgY+e+9cZIK5YSjX
Qe4zrsryH4AKsLS2+GtOd9gKTEj5qv9zO89UHuYypnJFJ1HvS63TqLbhvxWZziBSmw8jy+4KnZYL
Gw9oauMQc5p6t8hHUTOb81J+/8Zu6FckZ9nrvFbD+IUurGPn39vl9bjo7Y3WX61KEfKVEaxdBYmo
QGaQgtFhAdI9pGEw8apPkM+Obci60aRzYagqOY/XvPuTjvwHPd9FvEO7frxq+BvXP62M+An9IaSB
wtWJ99Ta6N54yDvt6I1ongbESZf4WiBGdJU4YjWKouuqSds8EAv6audMNp3BgzFyN6W9A/U4c49r
u6Jv9N6Bqi47u+xQfkXJXMYB9ZWsxFYw4lYHrzjkBKZ6X0WQZ9YRoa13mLAdObgvNcpEljnIIYN4
oj//E6NaLNL+hQ06db7MvL7xnyWoYtyEItGdvMoLbtZ1fcLuOL0QMdivdkLLoG0wJnIziNoY8OzF
hgIi49RIfdXoz6wx7GWhReqlOMllsx1jr+KMLNQGnCAcsLDE7eBLhaJZiBZkJFtY7nGzucZniIVN
CaVTYMC0BI2/R5OndndxFOil/fKmer5RCAlzQhOgtPHggY8AxrjdLVjfhJP93gVNGAOtrHgol+ix
BjekMPuyePf24IS0vSiwhKQUYT+7PtSWaDFa+ShR05g4ML7vli/GcetT4vWXgxteVwk+8Lvdql7g
k/jyoZMx/Hyr7S6hD2c+PCkS4VMD3nW95qrH9MmT4mXfIlKoejKILgZGNVQITZLE+dhjOOXUy1XT
L9yXyFIxOlOnR77Bx7m4qzDFySJnghKDsu69ifZmAoHvNVyspGR91EfGGa9RcGOV1vuymrzpc59i
xEVnI4s6HkdFuDDssg7S0YV1fRDfbmIJWcr/3Gl0i60XbIYRKZLJu2lASqh1WzlwMq1E+oQfhgCR
wyB/saFzjih2m7T1KBH/UzUg/6svLCDDm/qp1Q+pzRmbCobyoXZiR0kaNLGisLNu8q2fxr52QKWI
AFxvNFNPfWd/xkppjQ2WdUpR0t2VtgPl1p/PgjqtQsjr+bVNEpz7YMwXrs26OCiiD27GkRMzNZu6
Zp3oQXmto4cL+3OMQ/6qV/WPfeQHCI6oyPrhigO17aXZ3Ob7rBQDBy63hNtglJrJ7e5zhVfRD9ck
SQ5cxeJCjvEudAY/gFQJ2zWtG7URChdDyjCdngecSEEAdEuGRwod7nPUNpls3czkmcey2Uzb9qwN
L7d0Ra41kevvoev15LfaphYlaVMu6sSLlvlmZxIAaAbYIkvRgyPalj2Mxe81wbOczIXcS0r1Eur/
HmJWpuTQGEpe2Knt2XE5OuoBdMbYbsJaLEZxdew8u6PAy6es5wefk2S0UXZqZksJPPGXrlPS2hGp
zoLCkeQhRHsMEATzPmziqHIxleem4ov4bcgHKeRUDO/goyg2XPVW62V/wzCqp8by8WFkrLT38Gvh
s+Z1+VqDyesiV799zEq+x8rnsf1pdMfszM3QL4AiWZtZU1fjjyXb33FeyyGTAKRh4M5Aa3Rnmwxp
rzLzrzTS2D0Vy4mOTkJKUXnLbhe7chvffx1pJIQEgFPz+47u+i6MeptG4w2yOaiGJf0LgfpIeEXN
kavGF+K1xvV1URve2k2di9rujBM14TQ4Nlbgy+EKuwXX3mPzqDxTPvGjec0/vs9WpEcvymxsYmv6
OZOA6g+tLhhEIoQJspqW6MINr5L2x/eZFoX5JhWPO8bJdLvFsl/E4rUU/zaMRmaaO0hf0ujledW8
/S67mik83X80NqnAX9mQadDvRhVI/FH7TwVJpjAYr+6gmX9N6NnRm0sCNyGtTU3B5cLeG1T9Dwkc
LxwuN/EM8F8Lvh3Pi8u4EP3JLNUOoNC680bzixDdQ6HvFSzunrV6Gntzvc0Ui+EwnFChJYV/Z5/7
vIrV/XvO3OLTaGQBnE8QPnkILqBwnLPK7ZTsjWeYi/ArAfxK5Vx7jZvId6lyhFbmk+O17u1eNMOG
d6RmcxYjhYBdC+0C/rdKe4PBNqN8klOxrqRqmJZPQe8ldvagUDzdWXICSl6HClDXeMPAYjhqGbhj
OnmZKwg5L0BLa/nBsW7wCrXSnOji1lB02c8ezeOH0xiGucmzIYoeiq3sGRoHigRsfZNyL/8uRMrI
2pXht0oZN8NbLc7QlLNqKF7v7dmsM5qPioXYK+veHhVhNJE19rPrPT0CymiFyZN7R9wjvwvjB+61
Jf961isVGptfVV98GI0UCpKzD2pE33L1A1hTy6c8jMlekE+gcR/AelG86JASLfC7cELgPGKauFcG
3h8JjU+1V5gC5ayTMJ2ywRyDiXqZWpkPrf878P6qJWkQ9UFIwi5O6tuqh66OymuZdfCzNN1rf0KD
r+ICtCYb+BVQ09UkviAlNljDS9iinklwuHgGhlWN+fIHEL4b8719yGMbYen0nvrdRVzEZJeALDkA
ADn++82vPyL+45TtTQa5Il5vlTw4gL1QOyOsWW6opm08CwBgHuAe/RX8hK1+jzsl6zGC3IqR64vb
xROPGmXMVojLCbgK1iOWWoKr7EgYdnS4ALUsC5esp4LABl/qA/m2U11eRjKAHkkTx9Z1Vug8vwWS
ACZXdTR2tv9D4zpLfHeGkp3wV6ywFLtPAyq3JtMxFGVkTfIDFtjbswzfgFhFrhBg0xUtQmjm8PI0
8NX3coRhO8LXx9wkFOL6TvukRFXnqjT4ZJCPj3aF0ZhJKn7fvCsPYLQK/wfwGorVDdjjO2D9p9Wp
BTmN2H3XNnKlSJvDHos211EalfcFzT/WQBes7/eNFDThRK1MOkRdrMMxnSWMNwcnDGfLB2uq8m2E
tSp7ORG8Xp8pYDvBnjK5t8E09m4A5RtrzH1kO7cmiKTAK6YlLRtOvVwh2eAfacrkj31jbMfrVG47
hzrDqF5gXGzDCXwF9t99uPKXz8OfPH4A+cVjGFKjBkfgUTRg4QtTVR3pGMDdls5Vvx33X9TMPFTX
nXmi5iX9ZLGtCu406+S6DwmeCQqm5ZEb2G4yLstrgtwJYP+1pX0e80fMfOgU4D/8nYPoeCQsdDXV
MrXf+Cqay4Acv8gg6+Lht3KLvFyMt0TKVQGV1YsQUcHxykPqnrdcTx9MXEZVGB+vcFpWuQKme0ay
X5/Bh3HskV73Pt/yeo6PVhUv5DJgpkDTwoEfwlUBLpL7bXgs64D3y5sALeQITZEyz0TOtdvRvF9C
eMyJRV9tACudCBkTehsQU1h4FeBA4D1wqOE71n/lcw39vHeTzvOiYygJTOOmi/GArZbeULCt6t0Q
aDyx8n/8XztdnMO9aVVDJKVdn6NE+sxAuSuacqfKfPEQPQoPT8A67JtJv3II3ujJC/rFbZgiGP8B
tYVA7CJ8eOVMrsVNZcyvouQ62qXBU5unwBxEOtEgKVZRroi3H5kn7Gq7GdqBwxY6X9Cyu1QoXYP8
FC/AsQRudyVr1LkjaLiASyiWJsNqvwGUIblSpRQNQBvgrYMDZZiVkq86Un41MhlBwLN55jdia6KS
iX6UGFZqkvj5z3CNH4GgNmaxPo60Ugd3aw82LqGFvIrGMbdBVUsYt75ZXCX3uqxYIkO65Tqa8yEy
AQ5QQpPBoaP8jHHYmLl+qI43pVk4Qf490OR0DenTB3lQR/zElmuwmq1LfTyXBq/coDqH4DI+VPv7
xQM4ZQA/xNvT9kf06q4t/eM1IYdZFLszuaZeSJdCpeqVsQtOWo5T1S85T7a6aVVgSXT/nYB8qihE
KDrBUzEWoN7G9nPNxqsMyLB3vJMhHA7n/xShveHH3Nnomx8Yee8rBivnZPyiZKUdUf5szRKdEvO9
+roXJV1OCeJK24SKeK2X41rwzMsXEm7XDPdFwQkCrW2bCo4YLXoZgleblpSrh0KFQ1YFhpN+qqY3
LCifFsOWkHofd4Z4GNmGj5ljL64gZ4ix4ivqUhQRx7Irac3SY8S7KmvRM00FBY6CrJx9m5qyW0jB
vEZkAgmYXnQ1JRaiNwXlwVXGcTHvOYKaPPO/YDGWZzmv1teyCv4/fLjfDq34rCRJmpdYDqtK3GOS
hjylh5rYuEFmUJJJa7OybEAaDsImuXc3obAE7WN5p8Dk2ZrU1iI0auU6LYURbrjY+JjjoCPHSfT/
K2Jl6aUw4UP5/PDNc6Zosby5sgxNMg5D6SkKCgeC+kc/1oWhQdiJor75XlIUIoocDjfGNIV7buMb
TJU/fcJ++vpAE0Qe+3kBtXtfYo6MVamDy4NmH9eQlFmLJ2+fuSgY8UY0E6syvPLoGJMIM7EAB4/D
FTUro22wn2geuXKGepF9qQXGhBET1mhTK7K31Eg5vhwEYa0yTFRd72wrjUCByWaKOFmtMwEhcFfA
b89POqOaMV/MONhkdeAb3etkFlbG0KCcUsL13H51s/cDsi7nGleeScMlw0TSDuI5YDyKvIEOI39x
LijOshUIhypP1fS2w+DsV5Wm5i5kez2D+PEYcq3/QZukDj4Iewlr1vDa3W4Jrzn/lPRymzvmh9qw
vAd3Z1RfePezTV+PEmGoMyKQfY0fSJkhqrTPIbwOTWDK3xC0UpWT5Ym9Cpz9p/rLp9hJGbH5dBzb
v7AEkKjABf3AK+vOxNoBfy/OY6prEI954jwZH2bzdYoT03XQRGO0yiKQ4HlbVLhLe3/FpmFmukBv
wz+UenFi4v3PcURL5QpwDg6NfM8PGQsbk6h+x0kLgexeOdqZAmdy2kc3OQl8BsOwokjJ6Tafq/zq
vrRVGjHsti8qf4RrnpIPMYfBA5RO2gunebnYxCVBnUwgfRLQjvsmoF2jKcBwcn6UAydQn1ALqSBA
FlcB5V5c5uqJ9Rke0gm+YKzwEaogk3prFZGD9INC4trArB6FXD7f/FaJASZPvLAjvBBEqicY6mrW
NOFuvhEvk9/OJO0CJc42AITh47Dl/jEUPFNZqkl6SOTwPmDCPWMj3wvuMBysOTFB0Kkwz9TIuvMZ
CD5p6bTRktyjantNEm/Z5Osan+BwejkF8X6uZC3AX67zcHjsc6PviGf0nw1XEWzd3jeUBSbDX5U0
JWJJGEUhguUuIeTZYyH/lGxrjCPyFqK9BgkM3tvn/iWg73+Ta798XfU1RLOp02rFLzQPc7EXxQ0L
KhRaDLkNu/Lyxq/4hxWk+yAlErwgvSTYHglKzGb+PlT7DTc8xViaJ8y9k/EmZWDXFCCphof6FNNk
VHD423HcLv1/KZx+pqqBQehs8FO+4cENbHvNmMts4Z0gyFHymuSl3Vtd8zhnc7eyClKm+ji8N+q9
WDMsqbnj7sWLGbBQU9wohxBFlj4dChDvPflVJi/U0OU7AM7LAWX7cFvStVwGmyVRZgZ0FX+y1Rnc
weX4ZjTZ7rojw4VXB/RiJfIlqw85h5thGvlA2YWC9Ze6mnpiXbk5hH25NfxZGexMXbImnzzr4FZm
JULWO+hMYJnXZctbQppICa4TKeOW4qvjTv5tzwvw8qwG1hFBq+2X+JaVxeksqiQAPYOCYaeUwCdr
0r4/uJQn4yqjuPFus2UwKmQbWH4cFI/5Qpf0aDxEH1uu+qtO+cfaJTyE6sW2htSvr4W9eTdved6f
2LfiAm4whsi7lSyzn0ips5V8xBnRLne0m8NfnBFSYn36IY7Cjl7WL2V88qu/cI9B560uK4vugAur
cEHtw/crM5m7040BxMwjFEBqix//o8a2Yb5EBjf4xhBahv3mvGf6CjKSpwrAIxqxgokNXvA4VxlH
HWrLlFDmGO0biDxMkxdvLXS1btG1ar6cfP0Ub1b7IgqrYWZ6Jk5vXunZ3E+Q2roVS7chjscIKfQK
l7iEL/N30D//A/80mXcJoFgl0iU+n/JJ9/gGdfHvnuu+IaXjqpKx6t6WBkw4YRvaqrIrbLSH9dHU
LfQA7R1snCGMpn5f5Rx+y+xEJPSzxxlO/Bgf0GuXnD4wZ6VE7M6jlmTg27AC7npwcBX2SymicDRh
s+nK7ml6egVuzjcAUCRntoPZB5eVr+xCuJGOkGJdoGfiTUQzgDp9QBRLle63sxJQUQuKYwWXbUeH
DuJ5fEac8btK5QzPrLu2dRuH6y0RmLVD749whyxU+EZDMTJHcvQ+Ticd+Dg7L5UDhyZylEz3TF71
r8wNQhaWQHiu36CMXk/OuqBBjBo8aNGDx4B+d/qz1ZCRSN3vEsf7hLUje7PsQEWU2yv2cNDGcyiS
n9kRcjqU1y8N5FI2UhwTExdcmSRXyrFBFooi75xfTtk3i+iWYAntCphSNq6xiIKkhhktS72nxFnw
ISlmUq5Go82n8y3+zp+0jf9ejQSmhv1WG4Wum86uToJQTSs8Ktj51FxBw62gdnVwtuRhs2rUp98a
o2qlPXIbPPVEIflx1EsCcg/yRgrHeNAS6X36le7oLkVMU9reYdd10LulN6QDwqQ4m1UR2lrHe5FE
wSSPd4pWxPkrt4iT2J/fkH02aKt3/CWIDuL4ESwO/ZC91I/Op+74LnkI6VZua2yEXkvzYrh1FuSa
gIZ/tGv6YaL33MW5Zkh/LV/HIWJyOdwDmocBTMAVbMy7bK6sqR9Sv0jX/Ir+LvBOkDNtNT/o606C
3MUQj7vmIEr4FWJ+/yulgXZKqpjY0M2JczD6zmI4Xq4K1SOWV9QHiYYeh6B+FNYcheex0xwZMclO
m1V+uFEAAOP4FUGSngjQdB88mOo8XTxWB1KVh3fVf+yfxHXwGwiGv2Sg5tYF8FqbVZQoz47Kpp9s
AJuCndXZEB6Jo7Jc+1cYXpGsQ3YhUPZwgYPvCaoYsC+Ts7ISOiXI3WdnMU46r2sg+n7CRbrKFs+z
0xWq7sF5ZrLsCL+5dfdYMbvKcJG3UQEQdc5OsIlfymGO4+gC/saOgrTgtUIJPODcxJUhhXXaFk0S
+o84/PgX5jh4Lwx1yNLnD1x/82pVpeuVUWBpPEpmtBBcOR4ZVrQJtZ+vCD3sbFK5FYddKj4m1gwI
Dxbq+mnbsDkkOyvtxa73bp3dzndBy5FOtor2tXY5uZc1XydvC7dh/HCkKTnKB5S+0rxC48NwJ8/D
DeFLc+c6uZQEbOW2G/g9jayZvNIPW2HJdWjDCEpwiO+QtbqEALC1ImDF8PHwBmGR6OQSSEioHIKW
enIfa90tYdfwFnxY/58sqD+ervC9wwV4A2RQZpFFYjAaR7M9TYMxN03cksGqb9zrcaPa0bpU8qf7
xYhef/7XqVzcyY9Hnf+d0YqMC/MR9VI8my8oWgS0zzz+RiNI2oaXVifOqBH7w7PHCpIWhmaBI8z5
ouq75O6+VIGOucDkkJaYhipnCKPLqJu7jhHD4iVqSFAcgDUzSZ4MexmWlRWtgLVahVtjO5apyB0D
xPaODdzliCqaEWTYLwiLgV3CeEAjgZdrJuz4oVpYDRBUuYxRnu+dOhPCcqY0+E9AtNq9yD50DieU
LX0qRaqCDjUdcrCH6qO99gmGo9UjTkYhSNwUEAXMki6XBIOHDqR02prscTOTqA++UFrSjg3LSfy1
OPbD01WPgnU1v/3Jdo6CBUnyf4hTXCiJCwmR4NHrHOoja4SsH1dgufy0AdZsjDkEa1Pzig7dLP7d
1W8h+/KuoQHE4Rv7ucqG5Dacbc0T6LS04KmMuhP26Grg5USNuul9PuCfh0R5fabgPBX3Cnhq9TC3
W/9Y8RW/1izhbdIsOLx7/W/u0zoMQAXXzdNB8hBpB6JgFbhFx1z0lw1CNHlARl8FWDZreBGOyJse
dbegXolkSlGt7N1yhhU9p/NSa0VBy5AbnIbES1LLeGhMkMDRnJC1e1qbXRrgMDeW90oagc6XeuCA
7MLZd8uSXEUPWE3fRLDjG6v2GNSfrVmIT3nr2I9PuPRJWjDSBJ33UAz2/BAdlTCO9U1Cdm3TAD1t
FuOMxZ9+gMFs9NBgG41ukZbDTzwO4SJ4t9rNG9mkyl0FXaQf+e+dnzrNbRLZXnK76QVvRPL3oGDD
q3KLWseRVF/+hDHOhECYG60wJ3CIpTVOB2xNPtJR04mcla6Y4xNKzItxa1AuYv9ecgvta+ZDmsm+
X/u4UUTorMn8nJxjABii+hWBP3xD7d3PpavT94MnYIwl9++P9CCJVRIVJiYt3gDL90uNUE1dTZIM
qdIvig5l3+gVrSZ5o+kLaY8EmEPCfqK3c2PBDbCABpuO/0ZDSQ3MO+LV7f4jdhU6N2PdmbCsQuSE
gvOR+UuSnzqHG2LNJbMgmKCRintxUBqv2udELTTgX1hx0bg0ZAnynPuXhHE8q7+xf/dDmOyvohN6
Sjo3oqu/bjnQJsOnq6fdTSmxn8D+GXhpl76PCXDS6xdLRyaf7JfUPT2tWdPDKcDF/ko1GTUyHXnE
Let4xzibvtCslTtuGrkl7HS02n6iWU+iOOdO9qhmupJ8rP0gCLagD0oQepGavaKMbuEAGGOrJFnw
/sCThGBJWaU5hx7EGY4MxjF2tPn0HLXSyBXEv+tuajtDOhYcx8ukNKKE4kqUK82hF2yf9nsq44pV
nixADNygEghyAIgAa9b8k3Ab+oajjdcTzqNM6NTlHhlKB4FnQffjs5ElW+fimwh9Dtgpux5dVtwT
86D4093QZNW8j1h8l/9ufY5/ISMNWIY32EmvcjX4lk/6SbuTSVq6oSS0X6m2oBmVZ6FNWDgGjfC8
NgnxPqPcrYoFr99XXdnaP49LPYvUvhROBLlygvDIeDZ7BGQzGmarAJFgz3wv8+02E5sHEj37Mi1B
P30CP5H0lxTUko2Fewc7+h3s4KJaVNYATt71vM72wQBRiBcuni9EDksZfcR4kmYX6pMc7glJHkpf
ErAUp42yQX2An5EM2gi79LupM087nKTosmbMnVgBVifsnKFgzuwjbtCALJI++LZ7twBZ018KLMyE
+M0uMA4hh88fsOoNsST5/7MgBA6rvBmPg2+Q1F+Z0svUPkWwXGnAwskE/kuE89MrIUZoXSUOBUtj
VVy3sy+M2Pyx7ipTkIRi5VbzLA/p16oxnZGjpYU2xCebYxhC8zGYO9t/UlqKfQj0RZ2Y+o+p4iTR
Q5yhCg0+1cYKWykhlGy4Avqw9DP7gPI+TkHTA5zffgWmeJOVP34opnCbUB/n1kfX1S4QKs+tPmPb
WXX+VKbPxXF6KeJXcuK3YjjMwanP2ballLSBgdMwlwoBLJoRo9A/6dRY7ufx7TBlLoid5bmyuO8W
IG+pGpdkFwlHN9+1T3QmR6+shcT3hoY9tjjrbQBk/vF4FYRNP4DtjfIiwuoGWOQJyMhSwVNpZC9G
RuHzaFVC5GQgPWPushCu7lJ4kK2dCXs7BZK7PbYvoym0UrHPpxKCCdiO04y4VqbJt/uTs604odt6
MdlBO0sd/LK8CEYOM2Xt+RwxAqqd8t2LsDYcB3pNE4LOpL9iDlRuDWkvz32eRyM45sEkJxhSYG7W
JlYf8wuMpsPLq1hUZJ5vPXdfHn6ZWO9hNBcVyZNAJnGl7nOtU2TxXOmcGiVFoO2htSeszdFCYVUv
Y4Cn4/fM/Hf6RliBy62jlCm4+eWrEZwSNAzVA7rEtG1XYSaVE5wXUmui0MplZDOIlznPQQf7ADf+
/1b1HD2wZ8PzlyE8hh+DvPAReae5j4kW6AVFXo0Krl8NKVezlLxobeQuBtQk4L96BN+XCeDJScTf
fcwZvf8wCk60ogHWTv4p1cT2/TvrwlcgueHLD63ZsfhRABiNgRq5GajCcg4nhafB6fnVnVYKPuuj
Ob5UjhFvZIEBPMlmxuH1L84YlwmNGU9LuLQoRnY0ybaNgy/f7GrmDLwJZxtSs9xSYm8wXD1eM/G2
nqoIVI72U/+ditNb4aUw2RLX+ez7D7hQv6qU9mQs9KP1UGkA3TM+Up8cgilImJPzyBFBB84s2tgU
YC+fGkEbASZCoyV2tuO4zlAEWnojHCG7xzU29EgpkGAoIvtWwcwyWo6uNph3Qw8ow/gOu74eSaOa
CbLa3ISC8SlxHmiPLULGElsPT0Gmu5k58OrTBy4TKR5yeDz8g9/f69ASnCDxNvhuw55i7xC9PwwN
/iXLJU89wg6xs30zS7aW5Crti7nfSCyBIzGlvSlBVeYqeT776zFllPfa5YNhw5pI9s6JR7v3n2Bn
enxuQSo89GW95quYiVNmmb+YUBIVToFoNgdihAAEwM5mi2rfEWz35n5fLqawLGVK+ma8z7HgeQdB
rE1tgbyrtb7FxpuO7jFTN/calw0k/EZkY++hdQRZ92S1aisALbLL5RGff2lfR2sFgVPxVaTPtVjQ
bcjjqG+eh8iBrnCet1mUJ6fJkSS7rtagA4aBLY6gIteQynHuztW3mMBWJYhjS8S738hFgOQ2k908
sk4S9sGwLF6+lyWku9qltNu0O1JKoap8zOHtZw1/mQUmn2cWNLeSVbSjneo4LEHE0pEhuvTQPPSp
WosH8xhJKM+Ql5j5AI3TtxK/PPEvYrqTtTzh9NhV6CG986YVTHfeURKNIdlaGW7N1KyKUczepJls
oT9hpXLW/8hdNKGADqhV+yF+jejEcFdfmhLp2UZAt14cYarw32o7dA9Mdv9wlDX0BNRF+fX1+J5v
l82rXkb2cgHGk9jjjBU21B/2j/REFw0au46HmBYhVzR6WZIAIF0ESUvDihL6+TfPbxXEzC1bTKgA
UI7hZtO+hT5sxN8uqqNlJl9tuI1h+N615tOcK+kjC205CbfpfXm1DPwT+Ni2JzWuuT6O0CS7d3fN
5DgQevmHNxtapCzbNk6q2QG2CXkQ8DMHXEau0/mm4Yf2VTDgYRyDhnMuJ/8+F3G/YXfIqIJQ2Np9
CZNlzM07jB6Mc76mkJTQdedZslTwP0Rbhk4bZwPbsD47VjLSvvQFhxgSB86EEpxvLOV1FV1w4GtA
+TIU0xw9Y4z4YSEUHqYpCHqQIfovrO6AGztbPvyEpilcA5i2UjyOIei1g5i2AGyWU1+JuLLoyUUx
eac+EyPBMm9GPzZXjJXbAX+G0wNH2w+LC4zCGZtIBUXZ8m+W4ee8zZ8DjS1ow0aQRnXkgZYJ65ho
XrVl2Hpu01QnXt0tkaCUQNGrnJhpTzRIpQiggVYS7taeJpUHLB+p8Q3jM/BebEdgEG5iugO5ZEVj
UZDHJfHdJHY19IPmV9sPEyOIoZAa33AHvbxy276yR58Ea73Wsq+c0Slk8qa/4YoYuR1Rez+5MxAF
EiDSaQkSRvNKgjtmnhCBAwNec3aQwd/co4PfBGgFRpag0s4XmmB6OWMRhVR9R57AxTKMlUJk7/lm
pdFymNdbah5Uf01yOXqUNSqSEYFXewYWGopYh90fxhz5qFD+IX3D4e9hrmFDLGQhS+q4577MIkov
9qBWbomQF15fX43yVc/qj0ZECqxeyGLBNFaeMsTjsYTPE+6LPFQqlB/AKRDeqJlR1bsJi1KXMizC
LlCdB2s4YGUYGgriRhlhaj4Mzo5GqK1r8R8tEDBrUqQevL/bqwe07Z/8ZiJQNU8tVAbyHyqBmJva
d/2EywwTNgqseUvJbVX09zDZfSl6QKMwJecLQGkGClS7tWFHiB80hzYEKaC7tAIP/fqia+b1lnPW
tibtft5mQo+4j4hHRbAVwhZ1UaoYWJ9q2XlhMVZIXOit+JBg4mN63mFHOPmKahF+dVQkgwFIjJ/M
B6FSs9dTD9fH4kBgnkOnu6+0p/bIg31/oSEfRZatZRCfn8bkJbn+QQgYo2CwRKAEjJo0bsuwDGxa
swQcWGNxpPWjlZl4FYLtGz2qGWaLde8cZF3RblTDVO17lDL18oD81ai06g4KFXlMlIKdHJnTQiiB
Lxrz8T8i3//KyTUEp/JqKvcl6kwVUzRcQhd6mTYbPdVSJatyPGfuHkwDEau3KR2ClGGukxKRfDeF
l1mLyk/VBt7ZVZTs73WzUx8BWyl9AUGjToNNTLGrNu0JcH8QFuC/u9qGLYBF6n0oBzIBZxnj/75/
mVg2VkpQBl5ArKwXRON8LrLYfRrJGXNxABmBYnuCdXy76HuE+nMG7Lf/lzok7TyWWlB6Fkxcl+SH
ZsGT/nv1JVpCJOTViqGDa2cQAs4FB4+Um5ckcGG3hbnz0tQhd5+1UcK5umyhHFBn2LUNX4b1Mh7W
I7ZIIfvv7RLnBw2w6nWXfILFqYTwNo7tDnnjg9jcQCdMHyzBNLcsXN++/0+pUVFp8KeO5vfoaLmD
oOhS2gp9SzdUd54vOiDAY7b0oEv6hA9wkYizcL2eZ4zbYnQMhAvzN/vDuFrA0PfQpGxMx7WNIL29
U5GQiAI573AJd198DlffSUmUYG36GUyNDIEJ5n2s/lc+suNzaJqjZPY9MR0LOZ8hQhO2zIGbkcQY
z6WyQ4a2YnvxSokUzyMRHsQJsMiI73SehVKK27UskczYSuduF+wdm82mfGjvvdRs5Oz5aJSHkDP5
mKgwsN5MaFtoa0p26Oo+9iiw0FJvuDHelDZe1evJaDT/mm6Ip7VOJRQcImRYX30FvTJ1pdFEv2bO
J5f+C6POoNmAhalTuIRH47zVjNEOI43gkgYvLEPBLFj2KNWzZS0Yvnnkm6fo7/eLiFqH03ZrMPdp
6OJuulfxoJBXhkqeyW8sT2b19kxiKan1faZIY5R8vXZxCOE8IjPFPs88UBDSO55lTJ5+4D93g3px
PP45luzwCCwYqA927jKSoaRWWA1OQEdSYWYMbEHhVgGzU1wJebKXHDgMJeT3gY+7ufR8B7H0ZR4P
dttEg03HaewSEhkwcYE6PDmT5typSW9lLr6VjW2Ibfcpr6VoWg24zHE+EBcB+yaTDvFGsYn/JkEf
SBb+17U0ErwT8Pj+yRzGiuVlEFw+ZhnFnMixFS9tUWpupCJTtmOQuUzzTFGjubi8ycIOjUinz9dZ
MFuE/pi+Op3AuTYc3F8Z21rY8gD/fjut8dlBCnIQs3wUiICoVDLn7F97NM9TSCe9pV251QpZ5oNG
BIOjUgdcmFHzIMEN4iRyLlI6mvojEKqR2l7Ls0bZHf0Kunmss6ZV1zZ5izEE7f7zsop8Uqy08q0R
h2pO/vwPfgleyWASx74mYce8SYdjXu1xGGYOonkvSaE75xiBtfr9hc1p7aCxeuwdhla52uxfnrF6
h7hwwbY3/JmMdKOBaeBZmR3D2VTGv4m/cY4V1Ljyxm8kIyWkKgzpzqnGh9k7j6SzXtHBQoDThUO4
TmjLborFo1BV2WlGtJAxwDX2TTESA/qB+xEkCvjbJrmxPzryCTwFoJdu8kKQhaE85OTaknpIdNSm
JgVsdOFsoyNYzdkmd+Lojra7kwP/OacVKtXkgsVMAfDSYhXi2NvzWf8Yc/f+piBGDt3njsf3Ylgh
zqQCBHGNBgARhpBobUkxfNhfkog0bHqeTBFxb0xe3RMFIvxdDkCpic5EuHn1Vzpz1etp+mhU44rV
E89qJsf5Kh/fSJGHq8U+3Jv75POyav9OuepVwk8UiDb6RHPrF1iH4pprDWY0MmwCycHohXFJsVG9
AFTvZHvl7lHT8ESfUru3fRW2oKOp/0ws7P+hmd/tOJ3F47Rh251E7gOYSg0CVQNSZNR3D6Oj0orh
FaGmjHPu9nfgENmUbZ8WMKCfz7NDZz++gTTkWq6R4b3OSSlRUYIUjCvQ/F66m9C2Ljkd+D+cd8v1
Zh4zCHFSrZKdWacvr/Lt0rYjbkSRjc7/E5QiMazR/Bb7MDCbYRluI9ljLlAXq02t71Tpw/yEuzYj
RdKlciAE1PZ4zsCNjwdW2QWVLGd2MjEZWkuaJFFatzU1PJrHgwUsrJ2gIXS7afHKf1fQ/qznNfBl
uHQcU8IObeqdFGLjUqnRlE9wcqWS/po4gjyl8gpGcET+yfnKIE41HM2rqhRhMTAmJ6QsdFvJ+/IM
IDKSvk3OfozlQ4UX0nOETkVX4eOEauzDCfWBiwBE9J6ktieMMsRNzQEOX/d7zoqUHkze4P5A74ms
Z/KsRsM8xAvavFHV1XXgeSaQUfO7nDu2Qp3sY9beYc3pArHyPHrRLj5JXDmjRfEAqxvgC3GVxONy
mfNuGSq+KCZ4JcbiYD1glJIEBLoMadNjUWa6O/hWtYXmfSAitKXUVUG24+/in3GdSnV9xpzeonGG
tcvKKT58Sfq8rZ8huZ5IeNJtz1X2K6jAF+B65GQI0hYCREyMKoYBu9UPrAY75sRaxTFULP1tlw6E
TvTlYYy2zhvqvG/+EAHb1YYWH78mfEmnHdYNmL9wdME25DA+fVWRuUpSF3gGeOhH5hQpO/TT3yFQ
N6zYeMU0pw95wjODxOOsN62o/ful17txVtcfaVSfSEaHu5nIhGSzuEVpJedETcKc4y7OWz90BLFx
ElEjKFo3crFJGVuMjXWXU5XJFLzKRvC3DeIQr7vjaCgqzI+A6KhgW04D5Ytr51iVgF0jl5DX31Mq
nDqLPCIZRlqZCTXxuQCGGYKaUB2lY9TipfiiPETTmdOUMFejLwUvENNjCnBS5UQfa9SenQrIOuHd
Jr5Ed/Oat0c/eKtj2LShQEzvykMUcmagVvPyuRxxsNHn+wX7iGchYPjdTNhX06BY1McBe5ZQsLwh
1TM5DH+mxgrljwD4L7JXTixiWCUEAN09ACl7phwoPsmjinTZiWOHVZeNebox9HN7G0Novx5VBz7z
ElsmqLM8YZ41g2UQs4DEmLXcwV0+5bGGxCMzrVwf+ntk9oAArDACGk6GqvxumY6nk2dpfRsT4+7n
iLypm18HbIY8Oifr8x7MfkrbvudDRQzj5MfndyT+qwmF8DT4gyfbkOtZj3iIyr2ZMSFakC9wBcgL
SvzNwqJrkou7cBrzqcrZVFMV4VvKNIRDxoUKhZ2LmX0N+7Nwi7/Qc3Mum1ZIgI1BCuJxKjYA8z1O
XDMpDzU0uP5y4Qw+2Ku/+NY6/CsnFxzNc8iRNapqR3z0e/ufqgf10cqqApcWEK9UmwYgXk2nGodG
EFtCasRGNBE3mdBESAomcOnEj/C1dn+26iJ9+eaWPZRiWWepgFrvSrNYG8KQFBsCXNacXse//GCP
jZpKZ1Ylj20kP4WW7fKkTzf9Z/3O4hq1idCu1Uli5Hlq2ceYfTw77cE5ep6q1S+g4bN/FEcJI9v/
t/sqNoYljAFm/TBtNJaBJLAqe89yd2qJiF7sEyCz/43oKwVUb8gZaF0m3+2drgz2XSby/JglZ10Y
mrqbjqrMFv9XzXiWzTpJGqClflsU/eRJmnaBDxwPMkhx6+yM4BUQSVqIsLUuPXkjBtAxXKsV3STo
IbgFIe6Gm2iwNyExfz5TVl+/Pti4kHAU4ISvGSWvysy51KplEBcpSHwmSHjxSkfYz6VwbSFIBJmu
EE/LoZJAUiVqAPa4zDg7frZ0iv24WhU1w6cAUjaTWILZVBC6H4UJEq3fz6+ifUUF+5gf2mel6vy7
20MMFMLFBhli7317jFbAu24m01Z2IGP3yjR65btJ9Ro5rIV1dz2Kc/npjyLN77lXKlvgwX1LLiCI
5BARnDPOXo/yT+4+wOXEf1FVRBOG86rkQZW+UEk30fUOqeRzppqi8hIJ+nTNefRZmO96VcGl7DFx
R6tV5qRrWs7AJVhrh9A0VIDu08RCNRh89CBRVkONrUg+vGDqcsJWdTf92Wvg0eluUU/8CJGFVj8h
ZgeR0mHOZO4Hl6fZGMJIvbuFRJCBmokziJNGzbS3TmNQn9KWI6s8tyw5hxedZiN+t2DbTQsHu8Ln
+wQb3a5sxaiti+mL79JOteVCvvfcJXpmSV6L/dp8iEoWMxapDIbCHfjm+zyasigtK/2HNf/vCqaB
OHzrl9JhO9ygwhTrNAW5CRRi+6ljHIiorzZ//iw5sEJJ4dbi7ZD7ZO57mRSq3o6r5JawgKfaTiWA
r6p7cLwBINLDZjicInij8pDqoa4FPbzp+blBW9BcKQzdMLFlwyHU641/vfVhEfXhtFRKJol0yFb7
5bzTcwrBUoPz+v5cxFxW1HWio65TRCjSzKRUQBWM0p1B7hcNPxHKwqFunwsUM51xBvXBITcvM/+h
5aH43Jtb5CtjO7Q8BPhqg/FsApLkujVF3JteZyl44XY69Ycs6OaI1gfG09dDS5yyi+CgA5eTVYuO
+37/mevtsGPILxDPRE/91Vu4R0mL7oBzA3rqCoggCabuOsiaFyO3YRA+VRDx2yKTXT8zwoVFXZl1
RgiNekOvrUDrNFbv0TeNstGk5oJRE3AbUzpRwzrc9MCgFjPOqkykqwXTyBRfnzcLIy/Q1OnRORN/
VCMMTTUQb7V/MHjYJcOug9ez6ZiVWLkbXrhpyvVdHJM4q+NbaavHsI1uHC+FfqM2Qn8gz9HqT0jL
I1GhOo4EvD2SocCM1T1fSr62f5ls4xZoFhrq7bscz6O7NkDmhw+bxjD62eGOPyV9gE3VT9z1fKNC
ZtwvG63gblqDwoS2Z+IG4Xpf1C3Zt3ObEacymyk2xUyxPfFuCa2cAD+FCd0vLsH4SuUaB/d1XieO
XNRvLTuemHSutSaeIEEGh0CuFKkhAfZChhfvJzpVfJ0en+Vojh/7oZEOUFNpuLHAf6DyzXF23sQd
I+4wGhvtqEqDrvBA3tjGHi5QodSm5i1hUxWSnIo6ylGak7oeJzvBaBG2y2EyK1vJe8hQ9dzM3X/9
3e5LmTbcnZofwEqWhS+1H1ztkrAJoARDcNp09eRRtL507bTvxRCta+9T2H5WTP9RTcePqnuJX3vV
bc4OgSLr59s2Rf8G70chf/LeHTneJHaALfN5qIr1YQOQu88xIT5rOPEjP6a23VyOc9eWWNqqNcrX
vgivAHayCgof1IxR/pTvfu61CM5J6X5jscp/yzk+ZH3xK4wXbcAFWS/d4WjInnMjIHI+B1DpHSA/
MpiyHR6wDFP1xx8n9xE4mQkCzzfBH/J9OqMQ5DpXIt0h/ywDjZZw3sss09QMH8QVuK4abnMQYzfs
t3P4GGZeSZ9SKSINtWfHViWk6nBwHSlUjk6jueQDHQcAWOpu83BpVR9M1IyeBjXeyQobBx+8aR1S
fgEdZV7Nk0WD2eatBWTUYnU3jO6uApW1IgzJ2IYPMTNdWfsAfy61NLTeqAwIWX4oMl1O0qZFORj6
Nyao+e7czseczZQcenN3UrjkuryNzU3jSgHwVtH98SFskwSDSjtmIhTEtFA/VFmxx1F0sclum67J
9M37NDV/FGVnn53oaQLZHpjd7651oXJxn6ZZHOAMYG8MTFaSusJ3RIOL5ZStMMTDO/UWx8vxwbVd
zpyXhWiU/ImGe4RqeD0mi+CbsMMBg4WVj+zF4iWH2Sb2ndpAnyTke5bsoIIqCoAZ5elAHMzmY5Xy
a0DzKD+03GpojEZWSBs0P6JZIzvRYof4lFI9ihQZaMR6jyV6odi4HdQ0VXKbF6NxHnV++q4nfkgf
GUk/Ixvx9Ebic+zp0beqsT1DD+v5EW1dqpkusUP2ZcpJwUy5811MEQnJ7V6qjx2cWDLdlm52kVYf
PW0dev0IMXnDf1qHz77OObIL0BW56UhIcMVHLrUg4xIXlfRBElXH94gYFlYuAiiWqHLTy8JUWorI
b6jLFUOTwoDW+JEw8oQGFM+pCDwfbQH4lxlUxB5hcCksJUbg8lJR8HhOOijJtqFcgb381CJPi+gv
SwgwhtCs7ixfcgnr17c1YzH8f9eY27om4P//b2oAv/n+NYWQC6ng4dzfIBzg/6/3lc5Y+gA3hS6j
87J13U/FO2yej9nvlIwc5o+XFgFVktiQR/xXYqyceiknmLWwJszCXVOQIYFXljaNbMs3QUr1QLKc
CwD3NR7UkOxEmV5s3jNT1qVXm+oEPDYPbJMuWXO55P9ZAzlxkMi/nTlCKWjGTfdjYL4AC++HZa6i
bRevkAmAhfYZUWuwue7k+IivEmCQ6madkDCFkJFwyMiSp1Qv7DArJ6UbMFEEmWcl8l+mY6eKPlyA
DZ/+LPO/8D8+sVw0m/Zq/E2grOL2MGPiR4Ni3S5vJeN6i+//p6sF+xl1zSR+kvb5D1MXQAAZ09gA
UNjxKfAPyI7IvsqIeSXl196YJQKKQX2Sv6qAi0nTP8x7YasqSZb/ogq6hpONwchhzjErkSaLphrn
Iop0uk8VldKFZXgq+42kDzItCrGCfvpDsqLebS7yGd/4qCArSW5UVSgHI4fifzB1e5Xi3Xuzunhf
DLHBuWv5Yyn/SMUiNeAonnQE9fGO0/znh4srvg/G7QSk/qBxe2HYGetUOtKw9LuT4lMnicVpS0bk
Rf4kSqJ3laECNIizipgCNinuejJEELGxWMPBDXg9BpOg+0YNOsUc8LzN1NvaOsnz0Vk76NBDqqFa
NAmEKzGMnjcAwSL/Bxm3ADbikN+xa5Xo/I4JSbO4LltIL5f8BCIwebwF5uLEAqudTpjuKZ+h26y0
oiOvRPmEGT9cI7epj3ZXq+9+lfcIgHbYQxuFpEXPSlQr22a1EO8kpEfGaYR2NKVrPpaBep9MDCkt
9tUlC9QWe9m0pXv3vIEJXh/o+wCDSc0H4R4JZ4IdowkFlfgFpr5lSm3vu5kMywiGPT0o6fHjhSBy
SqnqmIGZ98I+FpDPUn7QKaOYVmV0vYKi9CGg6i+PzzTn5FXjIO5rAX49jhMpwn0OT7FN8/Io+Jh9
VHI/seCwUOrP3TOq4BwcQaZkNZcjsIM1y4TgpgWfqG+7E7GR21AVWbm+XY15NHsdpwKeWnPwXMOE
MEoPepLNYWvMhSiflLoDMRTEXz8BfTikgP7zB4BZtjApI8yCEuoO6HkuzWlN0I79CjK7Y31tYUOE
OJwRm5iewjXEa2+SVRM10l3rmWmoopi5LymhEKznZC4EPHHvR2qrTFqwF82LK7fVgAXB59SihUoQ
J2XiNBg6Qz3TDzW+A4mruT4Xf2tfIpKwvyUHsiLFHulj37OL9Y9BSCtYvqGuQzAlOjG28JqlRElQ
1BZSh/gc8DfgnFUkHobIrvmu5hpA9wH4uHpXxqc8jLYYsx8vtdsRluvnJQ+uu02ey6YEP/hoW3tb
p19w9gWQpyuzRoQR2V0gQ9s6bERMKs2u4+1jy7OQsnOGw+I1YI7giEM+XGAblXTqhtou2oOVL1b2
HcAJ3xMb+bqidRw8UOXb2j4uF6nLB5MlABaw8sGmKsDQfTQiggiJUes+1FMlTZ8UtXDV4mey6j8o
0KtoRNVPvuGns8Jrs78f00JcNKJ4Uabu3RHcxq+597Ygo5vwAo+gHZMAgTdeyCXQaL1Bae7yOdJh
jmYB6Jvbb16OUrlTZkPJ95FgbYvK6ZPhMKXPyPJnhRVDfZBbvDyc4f8J11Ead+Bl/+RH8IJWMMYf
7fxz5V0w4NngpOtC6JrFd3D+PLWMSjw4nJRx+O5EjCplm+5pD5pYy/4yQXqxPSv0xuYbtzE+GKt4
cCthJXmYQWcIjEM0GquclRLdvMp51b9wRX3ngw60pjfiwmcY9FBzkM/qaMrkW0yy2JnP8LsbSpL+
v5J+UPtfDpbcehPLpt2MjZYU5NmJVey6qmO03S9AA3x0F8vKIdXI/MMig8lt79Ill26Kz67TrjTH
P3STDsuKzHt9e8Hwt/bZSAYQPpdI3fsKMXwN/V5JTxSjCwSar0i6N4NbzOU2birVn9iJXddDJXDw
hC7CmPqw96DZdOjBVGHhZAd+jhYIHdPdhdcQbJXPrBJ0i+jfUZ4h64E1BrlB5jX1SY1ImCEeW/Mv
zjPtpLfg+BZPKO51I7k/alzIXUVXk0Y8kx7B600ocZmKtsl6M40hqV/1cKETIv2vGuNDLr0Hkxp3
qBIyks7MtUOXrbTGSqxICKzn9pHjmtPMvI5IoVT0S7l0tSRafWFCJqoPhrTOFoxdlqvQvncHDbXn
HsYwKvs2oFADndfzLCJOad+iJFfO/NF0umw5N7I0qRLbLJ3ve+wsZjZk91yXewX08pYgE0H+ZBYd
GhGLSbhoXE476QhF3ej/h0+P4o1oZy9YRDY77TjmEifthgpHaBZzLZbw3E6FSRpzlgza3ahrFwMs
RBSjvj4fNX8h7h62a0i0NzSSV1A2X45Fay+yQUiL/a9mW48DpUbRFQIDNZTWI9V2ZUcREEwP2mbF
wt27ZDxnsS1uhcg7oK9bsInCky2w7rsu+DGUgZpJI6fAfu4gSBtDzQzULaSbTDHWzb3n0IcTVcwO
9W6z2+3JXSGF+LZ8YcwI96/jOzmGGLAtgXKfYR6RJ+jrR9aZQxcrbW0yu0oABeiZ+rXV2v9DdDVp
urxLOYi9NaCm0eQHGcPZNDbWmILdhC7IkPDabEdEK7v9spjvLGTmyAno3Ic5r3LHgpDRU9v5VI1L
saFqB8Exs7K8fUzPkIHUf5fefZE0lxGXKL2wTrRBeSSk2g08or0eX4faWJAftqPA9boA/WKUAdkV
5UNCvyeGbr1pbKzuamtCz21B9XSk8abHiUnqPGHv3tJtSLFYo10WqGGg3SJqSEK78o9sNbWjy7Qo
U27Th4ex+qy1NBBSN/7feAw4od+MyeniVr16G+kZLeA/i+XtrA1WxZqqjYvyCpJqgMyJsMyanL0M
pMUKu0rBeEAHc2miUAwkZpgjm43ms2EqECKZF/H4cUmpKOB34oZcWI3MxhHhrui7XVSC+ENgbB+h
hncCr3dnZEEwE1lXR39sNj34vPW1DrX/G1WmEBc3afFAJTA2WyzTqEzm/hDuwcvh7pVL2EHtsllJ
GmzA2r154Z8/rNoY8XUgMCtI60fIcm4rlDHyL+/wyw/eXtxX1o6a5xWtioskQeGE9acpbW/ZCKrw
L29XkGWJvj53i/5aQdYU1dvg1ILPp9KCt4zlDQJaEnhRRQLJ4XBzvUTH0O76QSs188U9skmVqH49
5l5bu3gISqG3xAYA2GBy2xuHgh2vOHOhil9IIqc7vuTCbx4m6ludeMq0d50mNoo2zrl/sGV2CZT7
nLfEFuTRtPF/XkG/W0NsI9AWLwZ05Ahl8719Wn4XzT5/6AEjp+8ioXLYcyjX9aeZGaU7GvdXcHuj
ZZvSzR6mxNZECEEjM1/TFxGoXhRQM1IoE3yQA2NSNJ7devva7UBSunJeNEkqCQI674L6xa8UB0sN
gd4A0iQUboby58MsRPqvrjOdNoO6vgEr+k/LhYkn/U8vy/x+VJeVqm4AmquBno0iOMz2Orne2x1g
Y8sFsIkhQrDJuQiH43jqqgwpeoEJLD4RzFjc41IGxikha/uqtZEiwtCUsf6DBFTi/mVXWrZpReAg
9GYr7CQDXhuJVnZ65zRl6grCFRDGuWw859gl2Zfe4xjzvY+bjVsUN5NCR8y8x4I13W/8XvDsWFiU
x46ZTXW5aI0JKx5MYjdUnihEdf2hL3jA667gAJXlFkbWXTZgNhy6VO3MCcKExrLJ02tgkU3B4Aan
8IkFphxkIzibqpBzCpd2PE2Xjfur5fXWs5caySaCHgmS+O0Iq5mFttM/1il+MnWXYz/cbMOg6W3+
s8qa3cnERldR75go4XTu4Mt3pY3DEocrqW5Pa0Gkz0D7LZENZWqaEUZ5Zblr7S7WkD0VM1KYwv+8
VPrRpCwuo7O/nVA3nNrvtuMyxQwZF9fXVekvlDewW2hM6i38597JN3aPNJphq4Aq4++WbkICWd23
5Rw17ymE/TdDF+4xZNhxKdlHo+Brwlj6NHW9Zjnc7tXM9HkF0unuOKMHpXNhy46PLmwloD/CPM6q
7TCVB8ffHU57VUBVvpCx6dvEH9FeaoR54ezthFm16FOUQ1sQwfQzwe//HQEYfyjRrV1gRxIQv20a
oCxiAtbBGNjhMvz/TYIiTtHcIN/2RKK391gShScn4m3h4dsXnsEOVwBj2tBmyRGVdJOLTf1xAM86
U1o5DnZo9H827iqqvjlnaHZMJW6Ihhv8UceQ80mmWU9fsypLyMC+24aZX0wepmQZhoRPPK/nXYuG
ZM5dQSYkyzlo1uy8TNxo+QZtpyF5SdMzEHdXIqTNgG3Vgm+qEHnjX1ydSvDHEYDZas+MpWCr+rw0
mFC6zoL6V06KAlopeaspNoWnHnQdYhLlFj/uYb9pDNMiW2u/Ue/PDrKcka9Vqoca/04NBP7M38Bn
M1SqLjlYb/jjH32UZ04k7FMIxRxKL8k3ID5b7ZE2R/yQEmVysfs4/HlBo+LNxRPSnQMIpF64livX
QZhJxz+wV7jv0oCM1ZPGgpL6P09VFVzTuoRUfwpHVKYzFFkX6hGYJdPxA+iJWBh70aJw1jKC76Py
B2yf/+QumtbjKqSFECY3q8zvqriWihIYhg0QpTGNX1AweCHSO2Bi3IMuKJFdeRk/onbmquFCSuBF
sU022lhMxCVc9sNfNeVv9nbf9CkAgrN0manZF7Ruir6sdt8cAqvK2j3RIHndWSatm3lD9eYwUEVV
5b9fn99T9hMjgE4wEAeXyrPOmiBW4Se1vlIupyznuEswa8BWO1vq7RCYdVInleCzk1KBLgJXOTap
PrlR5s3PvV2qUM8ZPWj9uOPNESVFPMzq9ViWBfxFPmc4e494q48vnxhxX1z3Jvxysh4x+0LhSgt2
TcttpZcs0uG9pUn2glYJ785TRPsM3Ckdok7Dg0R53lyXxePaIdbtQGwDHYS76+cQtBANgxR1T/wC
cLWQmf4afnHMC3ZoFcTl0uL4ovFShFBUm7mkFfts57aeFhtRhmP8qIlwf+Ft6mKpG0HMjlXR+O0g
4kKpFj+sqJLInrxWDUjMnYIdFlZozpsxjFk4uDZuKDqsfc8ZTKUwLc7beIq56SaHEJo5LToZ/JXf
PPttqf7w/hIEGJP9mpI5Ui8uyHvxgurHQwcj/RkVLxcXRusU/hD8DPtxkgvb0Gwfemfwr+9JMbiu
sCQHZJMV3n/HZWhii5bOti+fmRtB2Q2Uq9DnRVX1fdxw4+NppsQFNyebWFkDKM73ZfuXWEywjk6+
yAqz2eCpifW1lWELXQUJLXBLNVIKQDCNxwps/EP4jaG+pgmzaii2ZC9be7bN54F9VNwwQoBs7SAl
ycAxlThEBnHe3MBj1mfySg+pr+yHj4B6b5oFHtZHz+aLuMWRIPleqR4tzLyI6lNz7LkjPGlkthUr
gzntki2eAqflEPUsgdJQd3g4hokUxRytTBV0dtDSTmPJ7E54wojkmJY9dKXkOxqMZI82Me1WJxoB
cSKrfXQnP4oYWMBDFb/xy+UWiz020m04/u7w8Tjsf8KumGMEYFtWTtSdWT4zfn/zpNtZPeKbe9z1
a6QPkgeFc/QMn7JdxCIc6VHajQ6VDg1YKlIQUN7qtV0xeaR3at+pLdGvADrRsGij/5FAEfr1yC+T
hnC9ZGUWfOY8Q703jdcKRIjMcCdI1AODtOMMGzCxvlJtUENOXN3xMRwyV6WNfOwT3SV2VS2znvJl
KQ36bw4B1KTdl6iARLLeYNIJYTyliWzodz+MGX2eiLd3dHReDL+Ci+gxKKhCAFWjXh3eENzodt1m
EGkYNUI///7pX3Ck84wPn4ktoxWElG48UfxuVT6vawps+bnmfZKQL7youM7bpnf27D737DgJS+vJ
U362TbzoIv+FpMa0IihUpbmWzvvjTiLrP0ioPnsI3ZmUOWlER9AmhxaWX29cb6r2QkWXoZOAUOh2
5yFj6P0lE7C6WqDmcUZV3inbwYQtOY90t5SfRr8lFJanQZa/qDAb+ANEvlVf8KtvmypluJ1DvzPG
gYbb6XXRPMfEk3hyQQNFuXhIgDT12cT6xQdfjM5bBtXFUCpz2883W2LTBAEmajbFXnDJMzE9ITex
KPsO7wwg5s7AjDSk8Lv7afMEKRsvotdF+cxcIM9lXIX23yTbNspOjn0A7szBwgZpx76HFll4dlCA
K18TdfbYKC33OcqRLpuyFFhxA7S3ss/i679i/43hFkp/8Xos0rkpg6AEl1WeB4oNilSyydSnt55t
mjMO1qaOt+8j3+nwbK46ESVL7zO0Ix7N/dbAR2w5ADLA3rkmI85RvXAInwPMUDIxThPo9/EN/cf0
1VjDHxXaIVYiAoEKAbEZ1fDok+7z0NYJ0B/HpFU9XZlSPc0mE9q5D9Hrj1bIgBdIJu7+YGgQDRXU
dz/zBaBQCLrJpnqroOy5VIPQtW3/LuTVSwzguOrV5rEIZic6619dOU+kxFQD2PoBdb72HGFrJg+t
bL9VGtgwqSL5fxMsl4Ay6NjFG6fw4Tx+9fWyrpcZZ4du298Mj4Uulmez3fOFFA+UjUL3V0UbHyth
S4ehlINM0k/p04rSmsrif75Zcq5lEARj9neyltnGPGP2G9GYwzGtcYjZuuoZJJvjmndr+R3DfMmq
sppeJ0KKH31JIOvS1oZW+V5wZvBdS7h8eGqrjz/lJrGqVhPA+Ai8P5fR97Yxtlm4MRsAFQVSIu+K
aBSNQxnwLrFtTrWRXWpelgayFc2pZlS2Ro7NIgSdqwqChoOqvyRK08qOMLvaLmAF2h/9HAs1iXz8
i/jy6Y7AWqn5RGlDp7FFTbU5Y9JoBQm3cSPanfNkMq/DBqiDQLQkdxEd9IiOfDln8bg3wFsdFHxV
D43mvauAJduMI47bDlV34US+HoCqYjQwnpfElDMe0EHuRfDmpUM5wOnxJ5xlluI8Sa/kli3loxtR
6lbO660MxJIzpxwOQumThXeXN3S+bVzSJeVCaxn8S8GLnkRaLh8BvYH8hX096odadZpBTxmOXD1h
WlPqbtZfVmeN/qJqSJh1keG3p8DAWfFpHx2U3CgOntCULTkeVnJVgkWMmHJSgDYpfRzl8CN5nx1h
hLVvf4jME3/raswz8gLrortq0baXQJ8t2hoh2fSB3XEPlb6VVl8uLwCSbc1ugB5K9ydP4mXdGKLT
Cj65/TyHanwA4qZVMmejzgturfR0J/lw9TSTNLKiSwAlZpIrBOIGo8gJesyWx0PRVB8l1Dqlizqr
UZzeDjofN3ojPuVbDo5OwQ7tdFJSnW5Z1tswKfmn23nJa2EGUq/SVTHENEZnN+9k7Sy5S2QgWVcU
6GZjPEhv/QGDMzmzUwV7/n38eZ8id5beabN6wOCTn1S+AWGPQFSGfgqTodBTg0WcJvKPD8TqXYMS
ACCf8hdwwncasZoILDLjzm+ML5VlK0g/4hrXGzbKtlCdz7FCI6lMa6vZI7DyW9IoANJO6G+kzUzX
DSjHUiwnag29np5mQ6FkRW63P9ZLA2bJ+fQiYIMzX5yzpYZeae15YfAbban6FdLwcQ/2m+k0xiXN
QwAUPK4Xo41SJ56HwFj22KNwimylVYBztk+IQJ3HUcvjKsML7T8N6aPDRkodbaMh497Rl/iADcqy
uhT6D/UrLxbC+VVA4SxuajAnom0i3QIH/jc5IwRNX9oAYeb8rJc2FA5SSHq8+Wgw9do077oYev2U
YXLNlcyEWTJOzxTEo1pj6BK/zwsmFNPQpyb3Ruh/pyNIye/DmaLewpFxoeYWPt9Zl5h4UbrE/M0d
oWqFc2B8CAo8CQyufqKxfD5jApjoqFYpoBbZm3VoTtauwnsy1qeMD5eXAcJ9Nei6GwEhCOzV/o3a
pz3R5Sj12qCurJZqiGRlxmNrLx2955kv4EK32RsUpBgS+dN0skPFop2coG9vvGKs0f3IEfTj2Tja
Wc+WRPzX+OAFQeEc8mwJL41egfSWJPsohD0ktAim8LK/a8JXPJbADP+orWd/BG3riJV6Wwf0y1lJ
X1e8IkBp++tyd3ylKwlTaj+881bhCLQb0416WzkfSABjrwXJ+UUN2/IeyY35fNyomVm/O8T8q8AK
U8b6E0IH+OQISzZBjL/z0MZmCt28WKpGBtnrf3OE2NgvDBBya2s7XEkgkQXuQ3AIwOpcvkoLeTuE
fgnCOPrOCBY3mROvNV5aJQF5u9A6xrCHy97Nsy2AHzd6tyj+yCuciq9TS2unAhhMloaO+4vXGWl4
/VnpTVcm28v/OVRssI/PsBTi0U6EEIPn2kjE6ifPrnrw/4HQ+C1FzMLfjETBEoNQ8YFPzkmQmgEI
+U754WKmlgotMBIJ021jfbdrGK1dRVmhyK2lzfOw8Y/+Y0t0Is2YX0qIFGGm15XmXNa4V5mjRqaT
xJxstIPjaNcVL6sYR7fIvBevf+1eQEjaY+2A+kuUa2zKyvn6WoI75mFojcXwK60tJPTwoyIL7BLo
R9ia2T0bUMrxbTEPPXmTbiOPFqscDqXSGs6uMlVwdIEVIjlwmjsqZrHrk1l3ukzhwk7OnhjHWanq
6V+apo0NHZELoXLuR31OCw+PB8AYr9QjoLP2PCObQ0HH3Rx0FZdU31IG7De6XH+kg5z2uUG2/3bu
VsMTXeDFADYXXLDkBbb44mfeeC/ux4MdVrHSGTEHYqtKG3cGnKwOxfYKQxnvYnj1b2GPO1REsf0n
mTej0T4qtx42w6QlWRifiqeVQQAvulQO+gVshusecjHMAdqZEEtKGRh2jkm3lG7pN+iV5T8+GUP5
EAldFsxG40F/IlVsgMO+MgImEdxHa1lIzRVvK1nMRxNKWvZdbCyfncHcbjMlqjMuATXKkw7kFDXL
E+Jb8Wqa0i0OaAB6LsXe+sXr3GDRnomj0UK1Tpm3N6phIISRw+FDXdTOR5Ly7lFdkk9NEbdd/W9Z
ItqE695SMjEwHjAoeaCvt3kCQW+wxViHBugrPFYic6FFqLI17X3CrfN+mroIiH4x2Jtwl/lRp84/
BvQRjCCHyAxBHkARKI6VADD+eMzD1Qyk1LFgeuZlJWtY4SRucb2Tl0dVqHV0eV90Emateba7W5IC
zatHl1ogEfuNyXCR/u5XM2OSUz93jO4nkhnU11piba4V0uj3CvcQTy51bV7znFrOpb/HpmpJ7HyK
V0f425Jdejci1ygnJ2jrnf5GfErumlWrbM3gTIH0vzQfSoC1coFIb5TNPMfgfwjkpT1Px2OipgxT
61rDS96MDeEbh0emq8KLx2AxFjZZsJ45N8/1dGWb2YCEIsWTzqXhVszc0K5+j4LLjykbe6/s70rN
6Wk0pGbM1SWQIgopu5lWtjhoq/U8M0stBXwmPCO+8vv/jajovx5j+2bHHb411XBGamRV2SZhHhLm
s18MHHlJsFGFnmiwZK17YVqOVBhb5X+6fj5+3/M7PAph6wIeiCrvsYbrC+jUD/fgibQvbfB0U3p9
7d/oJ11eYh3MxZ0g0e4ypMyVe/UDrgrRq0Pt0cV+y/1IGOvKovC61g2RlPyFQN2lUCvJSsqopQVl
B3wlnBU0ZgBkZsOeZ8qlBe3iZpO6h1hPTyEgyf70FJQs9kNmQm7CQoxFysHwOk+U8RrK4Jo8+JD6
b5wjpvqtUE0Ab/JpvLuN6sfPWDEUnVmOYNVaffKz+H/VBgbjPwZsdJ7Rx/0Ord8zrCsH0eCo1jQ7
BQrtJVFTjLJltXYkkKGdv6eLo3XLYV54fF4h5rEB5SZZXhd802hSV0gnOupMBLnBeU5hYKfgORWH
7u4kLfnSTH8ESBBXJajhsGiQyc6Kci3vndzQTMWZ5/Xj+r9rhZ4qSDlmbxU3YNDB4xShGkTkdKS+
Jxo93UuLr4q9PT6QhHSJO5FVB2X0QUZHewtBdMkBAiUEhQxzAOxCDWQw6ZWsigCbsW03nZx1KiGq
K/C5Br+NnYsb9FwjI226XsEhQgvLaPY7Vu33XafHCLJsf0sppGxFYGl/bI3xY4HYjgLbewmz1pbi
roAsayB9S4lGbLX1Os+QHq1FGWTg6tYv1ATrBBepKv0QMEKnMc1y+YKortKzvcH0i0xqJ/MmgcSM
wOpzX8DVwZCg2ZG6dWBXvgybMgXe+nK5a3WJ6ANtmPUxHz4r7n79XI9JbMHK+yMngeVDQ9sPHNl0
fITy0eHZ+XpnjAF+wBcP8vi0ZDoRzT+PkEGh94N048RiLSLtIislg4NiZ1NJ003y8qY8UnVjB1Lg
oOndgUBeT852vvgEnm0oWQP/ZPQESXizbONfuOV0VlncGGGdwXdM/HHH5RArD5SpHZnUD34t4ioB
8kA/Jj4xouluSqz0h/ghebEAZNHiKqMJ/YDG3pWzh0xfXLoobN1n+PzidIhmQ4MqVkvRQd8bTqnD
3VEjC+4aWlcpPIt5nZuX3F/XhVdXMYrr8gzgWrkiDWmiezMM9sjmFiVv4tmvwGNQx8PRRpG8Z+Rx
1wm5U/qLlME8FMQ9JGgU9YCE26l4AIFs617YsH4Gw1JC0zkHm/vj0Dusnth6B9OtnDjx+N5j+k34
zK1C6Z85OKvtZnBxvnF2uhsTcVQF5o4pU4ADcGWwLebjELB/mG7HONa/KyeXejh4JAK4dxLK93h4
+QkF3aND/huVkv2QJ5mZxICUAwGjeBlEQpDjpPRhAjdho6EkPE4lEZr8g+mklcZZMRDs3ZR3uysT
qXG3K76j1INT7nLGeN9+lggUfvWlsIqlUZ82qbznd5odqJyAlRQUIyfEfGGjc2V9+C5KK92rYRFm
daa2QpXQTkhDO6O7l38+cbL3b/6TLP1uxCsW5Ti56pwQCWKqadLzXSPwVo/MaBDOzg45pBNyh/PT
yR4edMc96D8U8hX/R0XQ6o8Frrwhp+UixgHwIvCoau7iQsGoDeYflSIni9C7oIDaNeP1fT7dhpBu
4v7/DCh01pX8W+f2sFNO/PSqY5jgrLpOdZmNacldHHLqNHZ8n6yuHJyWc363awZ3KftBMNUzIWMO
qvpAgx3SuqvHK0qxPjXKWgstfYT9GNxjrPsUUQcBS9IWy+orcjr1DxNBCYZL8cehlXHENuavBjKH
Tn8NOgswCSd3oD00fvSM77VEcJO3cECg+qAu8UiTSLUtI4kibYeTzqKDi5Ixf9iklC3BBFD4fUdU
Ht+gM2zYY1IEnHIAKkAtFCnjxvd73UisR9yXvkW76zlrJWB3JkjEZv4EJCUUzQeDQMR3RyhHIFWW
QW1cgaH1MVoLnHkhX7Et8DA4c0WUcjpru0IFbkD78++5cMRQoGmJqzc1Fm9U/BCmyvY9Ct/hFsUX
eb70O1Kibvmny3ma0WOR1SBNe1Z+S16Xwr/q4XjHbY9uLFqBP+UG6qjdQrSIZwlU2UM8m5Gmu9p0
dv0XlRG46NUnkcpBgxYhetpCekHkHDdlH92RnTCnMVdHDm/VfBVGkzyTHt2j/b+81Y2prufvSxP/
oUNNjzMZOyORzQBAKY7/SSiYuHzWjdYPjv6iY02T1S30TxefUtrDGhpCV5FHnmlLrT4XAPQo4uwS
pa+IlFm+1JBVSCT4Dc2rzVv1NQ/2DbbU7Ky2ZL1+MGCygvuLlS8kt22uDOjMRClzHM+myjTFlMYv
pNl5VZ8QRPkiAhGet0Z614CA7QZ0f6FU0XWpDeiNHKHDeCIupf+4SfiG50O4k4bHPgm7QgLQlA/R
sc1HwWpDaUNLFmYMFOAJtYsewU8zGK3RGltUOI62Vt4KcdBVkGw+d8ze3+XkhElavG9dG3iPbHkm
IZBq+X2ADwQN5j9WFPW6lGarElfRdppZ8iym3Lg4wldqLv68ymQzZyjQhsWm3PWmJ7pNooco3YtC
dim0USigUJZYSdtSKkh7BNmg/vLOTYffk4oIb8og+fbeYjBO++j4eKNc2jq89j4003cwEydWVsJr
Iww7ULRSGBFzogICG/NyyG+22tFosMjKT9TdH8tm7orOxExxL5xI8/vNGu2nzNM/YYcc6l9/yoqo
vP50J2Mvguh0VXhmlttSnQd/l2UL47LQdhufNmnJwp04x+pb0FQ5hS5P6yu5uvzNMKwyoC/TRrC6
Vsr+l8XWCPJi4X8jOdvHJkbHyfVYG7PTVMdAE9G+GMCt7YB/b0hoAZqyX7q1SYr1lg8yO3zbEcJK
Qu0I+boAMG3c8bx7bRAtfjCTv/jrnLxLajdsmIMd0c+eQfA9dPaDXM8S5DsVJpJuVAh82oCkBBar
jp0BcYuuBNXuEE1bJQFOwdPM9dR02vGE0ss+rkjhGKlJXusm5PCMGo9JTORSw45+niXzFP313myz
1X5xyGqEWSpEfEFKxQnYvXpXTXSPyStQlXUntF1Hg1eAx7tnxxuRWdSMOvsf2d3NwRETqWAVnFy2
2i6rnAbUgzHX0z6qy6aI8HUO9Qu3ZDAS3ARYNz8PH2BWnlvlPiRZuQsjnlapZSt2SK+mZVo/18xY
k8aMPOQK2g1Q6TBvz7klijEgsLlq+NqIOT1RJ4pjdmI8C0eIG3XWKyABkiOr6ZiQhNsTYqJ5un+p
SYOsvrWuxwYylpecKaB4K4hC9q8KQblXImQorV9znQi9hJ0o5k0xq3QQi+nI8svZjRuLnOWwad30
NrjKM9cuvKCwKqHZKBSf8hEI42SmNve9jkatUzj/DeZ2GBpzMYBWDwlm/HSXv5Nvbfr2fwNiAvMt
lB1dCSyI5RcyZtR5qNJ8MSUEWROaPpsZhTrJrnsRGSptxjRbogdEuMuxdZbq26x+kMnIW7WI5MIX
ilEQ0j3DSaC2+ayzMKYx5QhE3pckqcqzkqK6wFC13qhKDIZeJolFQRsHtQ/ZR2gXQyLxQE54QSVw
8FOUZ2QYMvgWpTQ2B572BQS4tSFgPPgY39ctgd2ui1wK8IzmOfJKq9z9XtaFr5lcPiQ47dZi3L/H
Dg4wNTDVeOc0b0d/Jp3HxrWS/oSKQ9M1TZqRqi2CnOYFhvBbNoiVubW9Sw3Wk5bPykfM5rleDe7Q
9LjB4U1cD1HRwVJ5iHFblhlKGfyc6B172pxjqFV6GAyYHfFlW3NP6VbF2fWmP/J4QnwdPmXqwOO6
kzOxIpWmf5xRjDDuevQ5ePfBLTgOZnie5w62IIlTmvb1edVw32efZrM6FgMHg5QmkaxMv6E1dj9L
T7DhLxj7pcvobrDp/PC+A+13pKet8iljlUMeUwfWFIX0eAM2Poc7cEaCZ+7I6JV2Y5PRrhF+eLJr
8kSzY1x8ZYL91XgBYFwLCKU4HpZNPzgi6AxzvHeMBWzPubHqo/dJTn6ni7siDe/whPi8d7OTVIUW
gQCVhtzx02CgdAIsPwOP7HzHXxjL3CBDqBwmqwMHCyKZVS2mCG3Og5xk0uaijlcqw3f71adorkJM
c9gkMGmN/D0J+jZAA5+8fNCy+pxmh6xPtESxSCAb3089VzzG6cdjl2FXJ4lusQADPBartPvxdg0b
ngO/3GxyBAqfAT3oW3VWfTmGbIcMsbGS4NOSeXpjTasUCCYM1t1v7mhBjHMUo7QAo74M1UJ9axIl
x70+5/iKPt+7OF788Hp25YzQFHTA4L/xdXCQXUqiBt3YnStdtC9B/U8wRMyGU2Af4PG7awBJDDJs
WEPIYKAF54kEaOIs2NoDeTIhMIbTBAN5nbrf0DHVJ6eANJVvNjqyuCTswl2pUb9Xp0OJfyFPPPK7
bfQrbikNQsrHKrpvfnHcxb2YMunpvD+wHac4yhojdOLgOk6gED/Qr0w8rlqM20mX5tJVO6LrYOkv
ZYS/iJZC3/J+jxae0cQTEqayMqDDBKb9ztcC5PC/5XJQRmKpUo5nLC14VLyCcTG3y4PJsD7zmU59
RktSTkCTgo6md0TJl0nvidxKilOSp9EHcudrGg/Aj7q40qTRp5qEeuNfC3EiPr7xXq2QIAJ0Rdt7
vS/aBsWANnKsq6JnXgrMfvnf9715EsyC1b3vKXwce7xM7rVPFxiMuwaN9IfsjknOrPELB099tVAh
E1QdreacfrA8rMHfb8RvVRvidRzuJe8P/GxH1PdwJaolIgDSVdur82RU5IeE28DU9Yr18N4p7Wk3
bK0qugPMDOvG/cnrINcudSo9nQeue/Gm9nXN3mkKZVGsaE3J25hObfPyw4xeS/3DB3pfJUqmQhJ5
+iiVh3/CCfL+xXYi/E0AOgt3Qy1eY11y8yOJyz0uactGHdEVz08Dx7l8dMRETSwTHAgIcR/Oscoj
2S2VygA8Zv5WUM5qL8QiFxBVaUhI15EGBd6UogWZo0qf6uBXpesjBZlp7KY3Stnzba6ozr3aVq93
CRDHTXPhXzJgkMWcoAfFhFa7ZXlViE1UtnMq0N3SFph93UkqOK14aaRWXnFmHkb4s1WBrKc2iwVj
1PQUJWIvFFVxYHC1XA7Pf3ifHbe6UJTdGdhKLKsHpYP4qxJI8yNHIL8Be6TA0sD9fUaWozTwUtaX
bGFSzFCDLfw3vO/AIUTEHhSJ5MuSwYhp0XuuvQ2eC9xaP/C5bzhcP459pJQaJciUfmYts+0QZn3L
AdXB26EVT7oXWnNA0moqZBvn4D3vEt4btUhtNNB9Nr6mWxrMvsbDyTaZNgn1AmH50LfKbouMdpRe
+if10u6nMNa3rqNtT6s+kMdEjOOA4fwvEn1mPL6QgxejJpXQhe+PVoC+AqMkyeugVtJx7scwfkJD
peXea0KAevOu6AykaaEUT6SLDbfK15CioEet/+BivcfpPazpY1ZuIaWF+e9V4kDKkcQOUIdvbKvx
ABWo3gOZyErKuIKBDZQSCq15fqrt9aYqEI85iQsvhMMynpB+FNuZ4bdlZqx2xG0lkCCpWsYW9Spt
NXlv0Hw3BRxIpJNEClTY31Sw/gJ7hE+WODr8/ZvJkE3/t3MDBlFxfe4OXZgLtcE1y1JNnR5Ot/Lh
AWuPyvEoSUSzkmQxYVPOIDAcOqJThEudpJJqy++D1NY6eGnf/BzghvA7MbmgM3Whqff5bwlNFL8K
InyArlxc3OxA6zUgwu5CAhnc+waCRt3Qvg81pn1PeNLeQuKxx0NLtW1S9QworDmuOpZB5Ii3E9Zc
55RRXdTjF6ww6lRbnpGmcNTUtqVPn2St8AKI8J8VANkeHlb3t13XpgYBu73ja0HM8F5iEsTq2FrP
Qe4AXvTtJTKbxP/KjA2ZbukAEn6HLZshJOCEFWLctW7S+A1ANbF4aATaGRTP4cl0XZsmI2/Lh30M
cXghNGqtd0y6PSHNJwFNZAS7oS/y8X6mfECX8thjsCuV2hrN7vz8mLAPCEBDRAELEFl0h74L983p
kNOxy8KJGSjg6mLYPiNzgHlEHvvPA3gbabYjwbsaWBaOPFRBgLSx+3ZOQhmC+TDAGdK408x/dp1I
k6aE7RJArSVL0+NiU/m1iYsKaLDvzW9bwRkvIFwPUltZa09v9NIpAJAI8e/CKUwzZ5vqVKyl752I
2NRH+qvZiDlhHmhgOua3EqhkomTKmcRkzvX3Cr0TNLxAZtn9AQwgh0EuExFG2pD7ovG10bvh+cDi
jp628RRg1CWpfSputokvXIvs5sE1cVCB7BL8xoXhvPxizOqKk43ZDR5kdTv+jxIGZ6S1LVCV+4+Y
/qRMavRfooHOUh9bmcnGRz0Zrfq6q+LkkOt/IUfkX4vwXyhXaE6YBB18dUoadPVbHJEDtYk8Erm7
+C0xjAgQE6cH3uIvF6vij7Pz33MGcsTxTsfYuX+g7eL/dqtmuWihLouGhJQpVubyG7xA6L8Uw3g+
3AyNKSoy5nmBnK62oaQSBTXFM8UsewY5BoEjYQe8khKB5buyIkZ4w9ZDu1QkVz0mhsxbeM8Kqy33
JO3v/klCK3TXM56dGD79g/wU5lTY5iWh3cREIFAcwogbK5iy8NgCKcLRE3LVipLHvrWMkgYF2nZo
BEvRP77pJTqV13jxo3upCGio+/4iCkuAQBcBob8pKvgvINORhkC/mKnhEqE5MYjTMD4GcSFHu6Ed
DLY//HAUO8wfiBIAaHUu2UfpvqaEiHivXU2QTPLqV53RIaNP/4JbCI+scN2OobeG2dWVdJnYE/9R
sbZzAsKOXSA23CmMLBwLtvrvvEPrZXXGOntW2R+OafYmcoQwjAM2BFZakzWLKZJbDRODIibutfu8
dQ84+v2aaZ7BKmSrtjyMiUk0MICKD/XVeHMBCc7KxgrweP46RZzO+HygjhYPWcmrWUmHSHSaBY+f
k9QRHGmNupj5MDNHHzWawXAFNywdixNtHAiO2kZ/KIaKFCYFl9AE+pkFNdpOEvHRS+A4shA6kOow
12QdWjUzTuZT5CpyxVsaAqHt6LkDBZ7eTTY8PL/k2SOEbPF+ibEgsnQHRqlVB12eTZL3CDauXSv0
3jQOWXrXi4kSICqxq4Nmh6Isew7cZDO9E06SmOjmUgOh5nAzMJuEZYHEORZHjn95U8vps+X2+r4y
CYNvdsC7KDQJE+SoXdOSpMx8d8CYDc8gxfgmgZtSbG/bLhCvRvliv337BqYKOVrMHOwTNd6VG9Y8
8dJhgNHB2VsNPXlexqCVkuHnK/8uWm9EMGW0Yw8HHtxl3L6XBAdhLQCbVD5iRl82KanfV09wmMdw
t2VXjBMQ0Q22j1X8OnZWHzpVUHi/5gZ2ooh9LF3qmfyQsqzl0SUbxHTDihOh9t9+fgGtLja8Z7H3
7lcdMMkI8kI9W20X34jcpejc6bJLKAmW1SZn/riRRwIuKYhmNdXes/s9ebFgA3NT29hyHUF6XRJ2
24SEuZNEi7L/YVWnuDTKc1T/ss+CY4Dn1sDQAdy9lay86hTsN7C2LVPqXh9Py+0fymHyQfYUq1XC
wpRn/KApXsrpiyBh+G/7C8WyUJs3hBBbYSX6ybUx4MyNJ4gCefq4YyWRwSeZEQyiPQukoZFqX8uf
IBtJJF0kWvWa6zPcbjFWoOSnyWJXNJC3PFeXsRWMcpMmZi79tcd+sIswwOOcNmjJk6PAEfo5aewT
eTYykdILTo2W12PWKBwlRWcHeWtjWglfKLXvenou2N2PwG5Bs9JduYdFcCVL40UD8i+JnVRtqWts
aY4gIJqmehy+4BNrNQwJf6+9Lnf+W7F0sQ8nPyQIOsfkbbV1hHtRoYrDGpbwfRpVI2rKez1Ic181
l+C1iujw7Iedw/VAshgNjNhe3dAP1H1Fwf2dnostsegmTYus6bfOpnGAKEHdqCo2hy/M73kIFa+5
dbUThPLb8Werg+jd4afgtVZmtF1fWJ5ykfC8+4d2Dw+FV7YVmzyeTwmdCLdozpYd9sMWs7BPmAL8
M1XWqe9rGh1wNfG4/VVBWS4/cm2/fFr1vJ1UhHqQZsez3uCh8+FO8Veed+GNgKZ4Q+22TQfvlBl9
q5V+QnTP2q834VaBXlH3pLL4qPhkq0a9dGB4+E9b3VZ2DAzkNu1HYJnU772jhIrtjNMytvAeoJOy
CiHK0jhUNUPoLh3/xyXOiuhPGBc3OAGPb5fOiEvZFw3MTlv6VLdUjovenLfwg/AvR/2WeLgvYe5r
KvPPD+YZoKOUToDOPwM/tdmAkHEZCHUJNbNxrTiQEWifrmHt0syk1qTEG+drmNqnXYD7JVkppFPh
nsEkQbtkbcEDKC93NKfq6UT+DYKuV0L7nEL1mBwpnAAk8Y4Mwy2UY8FHxTdZFmCvhaXs/adVnTWd
xqzgY+fCZ04cer5iJ281qEbVEppf+SU2f22od1FC3F6eSOAOevlzw2ouMhifC/uI6y/9dXcVtYiP
MdsH4Js3amHqLI4hyN5G7tcXOBrHwyE4j67mV7EJpHpgwUo12HeTLrMUq8LSnGf4qsHTExAg8ww+
+tnBx4BIiq0G6WAS8BG4PXyCWOtPQp/vxg3JrJBDweZOW6BH7V8OEkYR5T5cPAzZpCz53dUVUCvT
In1IYIrE6dfU4DnvGX9U6tWW6eppK4MK6S2fgBDgnuFdQr+HtPgs1sRO7fuQjMH0/xbG0Ir4jFng
Ic0oLGGRXes5M0qHz4IE7Pz9jKeXBZPFTdYzqBOxyhSUoRm1q9VE4hsy5i51LMUUcow0ucOrJTAk
GnOHc002riXbGRDUjxIT5T6dcga/PVO5HwwidQrrqqo1ruGadWVcVb8lONG71e8mRGGnL+hczMKx
9gMYvPjc5KVP5IErm+RqZdZuB6VuGcCNruIyEqNpswgDZCZQLGpr/szUANUYHSslE0aDDmHfBi1s
BPNG6c0EuWGF7YpZ+iB2rsxitXTw0UBj3fcoVGOCp6GiwV80fIjzq+h4nzV2mZWq81OXIfCBgoZs
f1iYzDy5mVH/u61HRiQ7uOsaEMmusS/Y1e+ccbhQKbLLK/7Ps0Cfp8XQJz/JLg3fx7d3dw7N3q/x
J3pIUdhOqqlqgeEHZaXXA+VQTW2GpFq4QW+Tuc5HY9gst7OtBN5T5PuZMiqh+oysRQbHjEFyfi4f
5ePJyDmy2MpRJwNVIQDp5IASTlAhpirYY1Iv1bt/t2ZLUvUtPeJ0G9asnla+rB4utipj7Rc4xjIj
zLUtW7j96O23ZdF8B64EXZrlB1+V+rJW2uY+ei6929INQdl6QFezpI+7NKVAZlCuspnnGic4QbTG
hRN3qKshJvlN6wK798rjboq42w+bQf4abTw85C8sa13Xa4lB2aKJtvVtUbvvN/bouqZbWxzrpHqu
fqwMawUgQAlDw5XVRqvB0K7ObijAWzSiCkh9shY5lWdTH8PK0sotlEJSQBax8Hq8+5xBXStdxMr5
oJRudPs32AZ3JZ/+QQ0AxLT9Xk/YsNzp5lCakkb//XrmL7RIPCUX4kPvowGUjA65psdyZFxlR3a4
iwxpatSpJtRNa9269RH4eTv6blLE+2yehjSsaDq4qnyjhm2DrcfDRGj/KxF9CCLe5feMSHStQlHo
cQkqG0dJ3CVHJYyoIee1yMV7Ag4grvuiJ21bv/MCCBUHSfqensOY/ZR1Ut5hX2xTNwGvX2VOzQtt
gEgXXnedJEjg/fGmEAmIu0SiaE3lGVvqEWMol2OezES3k7IDeBuC0hd6gL82t1BeGsH1PnDJn6q8
/2zVhAKRsk766TPyAzfwNsn3BHXHGPD9++pyoljJeMkrwN7YBkOYHO0AJUA8BcoU0aEnuNC9aTHm
QGa1ZI7pDWxmDiGNdb9Ss1OUjj04VlWaaiGzHkvDRi177+hFl7jTKE4ZFm6qMfoSRMdq7zgPM0I6
MMHmHUn7EGtEnA7BEDYYz3WiGLFC28mXLZB0k0sRxZfXiWTWHaX8LChy75KghHX4uCJto9Xs6mgS
Gwq9tXbvLSkVXbUN6d1kr5sUroK6CfJjjtCBiTIobSYcTHKxb5GnPD9JD8Y0aHbSB5ryjfQTaf5J
2jL+h96USb7DS9PmUsN4CyCtnRpEmCDDSGfUEgE8TULqiLFLdV2olCd7SeZc94VlQ8oWJGbJjD7K
IDOlreVgTn/YKU3Y9Oe6a18cy5SphJc4Iij5h4c+dj/+Pcc+n2i08SiE5IFMobrjjvgYz92besDJ
4Febu1J9mdo0z0JRCf5N0othNOeUO3g23xC9UscnxO86jjifp8MXDqAVOmTlojSZFUamIi82YOUv
VD1kujc/+pikRtZ3d6lgWVuwWoO4GRGXmo4UmQzK5IrylIxAfojV+O/+D+keBrq+hw+f92KIAe1O
Zj/e2DMJvAPEQ6D/AbC4EIHBL2GIBZXChHsNLss9E2TmoB2CN52+huVX+cLQ3+KWv/xZUbOx06tL
AnmNDOzXIMgxouLkyJpxY69Ckroca9LN3IasFbHrUegnerL+EdpPERPw8WhndaQtDUq3YEBfS9H4
ssrzCkz8AiKgQmIOvWCf19TCe8cfh1246fH+g/0sjF5C5wrFdeJc+VXKL8yZh6Cg4i60XcilcO1J
4ZldLNjaoJz5d2I0j5r/5RbPb3edAPujHEAEhgCw051+MwU8n9bOF6mK5sFB2zfsFfcghVYPpz9E
DVBgJZ7iwoUTJo0vrvLEbczrng7RE5uoFuJqFIhDRy1KE0gt655xSgy3oaVtF3hFWvbfxwm6L6ul
N1NQKLVqQmaq3RBEqCtiEIJYLEX8c+Cm8afeZlLfKJR1PoIOR355jhGzRqdsVBb3jvziTVNjQlXY
cKAIERyFyc46EJzhZScTLshIdVFeFKFmP6JkL4++95BPF4+xP0Kx/tUgQAlc43q9kTxJ0KAX2qqZ
TaLXltnU85hgznkNwDE6xygGZLQJjI1m9IzoRJI1CbqFqhqKUWU4XyZ7L1bN7re3fpGCbZ3P3+tD
pN1CUsAgQg0uEqYCDYymRjEWF1y+Y9DQsR8gyeitoGnH0D2417Cp3OvzC/HHCH7+wjUFU/E0ctiG
IdoFztSv5txuH/CWM1pCS1xAsOQxngjJ+9Dg/lZdGLe/2IUVnjqRc/quov4MvDaS1MMCkvQjcU+3
bwqjE1eQC6Y1Hp+ZtBYvbwPF724I5yhNxME49t/BU3qfegSkSVaVW2dQwa3TeSPWarYXW25h/JuH
uytFJFg4LCp3edlX3yHFyG9Tyq9OqnhtqZqhCIlQgKcFA/IxEtb95mhZSN+cQsYAM1h4QPqKod5M
uMtG+szGqjc11zuq1b87TFwKezOCBE/7P7jwoyD56hbeMEp/3iOfEBC796IC0s3ey06TFLMrBFxa
XR/D1wEF8cyrZ31Jr4XtXQI9gAR6YImh2CJeuGxJyvSwRAYP7gykpfUSxpgkrw5ga9yGqHYf1QMw
aEcDHrhPpKOQmw/lckT+3LPl+5BMi/Zs13AiR9AVO3qfmZTfxlUPH88NVre+aFFVYMJ029bq+2PP
03B7mUmeOWTrdBbRgwtFbUoS2fFTPAWyOVyyUEmxGmOQu4gRwUSW3oeM3i2bsXNJmKMYG7HFLevH
Onpo8/K0udf9vPwZdYVWL1l86O1l/bOUwb4WKJSQMberFAQzij0rEsSe/6T0AZpcTkiC7Lp+mx3t
eGQqY5C5U4It1sf35tuHiCs+gbpfbv6AToHINhx0w7s6u5L17ydagAcgAKNsDM3ab/UFvOLkinzU
MKNMkSF19Xqb113k/AgWMreV9UeqVBTrZdyfOftJn0ynH1Jmr+3UVYc2Kg93cZ44SanHkAgwadBO
O0H21Bb2FPbc6H2U4QR9qw5mP3xdKKqqi94S2Qsyow8o2MDL2ilYu1eC8V/u/amIiuw/QhLm21kG
N8t6B6QA+qDs6ZEO7Tn8D54XDlt5pSYAL15EvkLf11yBGISggdVYHzkP67LGzT/JS6ryWRLwcUv6
lknUhEwfr/fSHtg0kpfYAZGSqvd5Pv+WrbtStZVKzp7p5Kdak767YG+0h562hkG0WSyw9nGP9xw2
UwrAfrJBhHGQnMNLoPXbvoIqS407k79IPj3PyuuBxb2QgIOK7yItSaGDdIHR9ogSQexkuKn8qwjY
mrWDyYJ1gz5W5ZrMxkeg3LiUIhmbTsE1ZEmS9xFTCsinpxa3S/hz1Gb1iJGQaSPqAIV8nqBOoZUE
y7ez4RDnYS7xpkSAni9e73acVAfmTFYQmc8eWXbp9e0412P8RCTdOevc3E1vWIH9MRLnWkh6HtSb
latBs/XDIv4RN0WoQaf98I5JGsqoBlvEv0OuuGD0rnuwQ7rGWtV4nklgxv5kGNhVLlBe3hzez1jy
9IGnqQY5mS38ciCpKtZwQjELiBcOMABmf2Kk34ZvkH19+DOW2Vv7ucY45APtEdJEkcF046K1L5+G
QiLC72zQlqbC8nliqwyMp9SS7MC7/M+pCYA1Q4kay/daBx5p2hKFYLR8yQ6qupP4vPw3HLePUROj
ExRqfnexuY5Ex7y2O/3pPw0HUf8Jv2r/xACWzvoU4bOBWYJQRnnWKSL1r8kIc4UKmQ5Hi3tXOKkH
A1Eo8P8CQRQx+D2Qbf57+Hu+2b3F638zNiX4dzqHaXeR2nnOzO779RYlKye5AVnt9JdoQRVesiOy
/x9BUFisFFRcC+O6+oo1wLIHx8PmSpwVZvbCyBzZ4AW4DY1NKMRoUcZA1xQ5TcBMXOdvsFES73Rb
070z70wJS9tMPR1bQ0VXO+kROohCAw/vPObZOOX5tqEMves/Z2G2GmrMDQFlv3K77XIMy6W5renD
mXZie+4znhlRSvyOxUihWKacodgRD83MtndPEqRURa/SK8Gy7327vlaMTixcnFhIiSSGZj0VuvZa
w1tWN5/u/kNPvMbiV+DtloDEWB10FsnH/JbrCy5ZghauL/0cZQnZwxyqHBD6TJ5VlkcCfMtfZ0Pw
LvXsgAA8PE84QdfqhNpn8Ks5yYmuGkMXwnzDTDi/5gNJzQftDPVzcchOrfLMYIgXBbNkOvgobQbw
CJFXTksIApgavcQnW+lzWfVRnEho1HuujoNkU7nBljv8ZdcIbfWRDZTbRoCbMsy0oTca9k9o38dX
O4MHKWn9IMQSrdM+FQeXNddkvE8SwGH+UwCFMZVUVoYd4ZG5N7/JzH63doC9qJC9RzvbNclGeiS7
bRHzpXkqAxexGOTO2eqR6tj2wpkP+zqP3mBeDv6v8Lpiem0MSA8Ri5kEjLOSVlAsdxMtZupHSxXy
TbxiXConZg2KuKBHBF0bIEY0rupnnMc7OkI2/pqEkOwg+U42YCEu84y8mCNjarWe2Tvyzh0YAPsZ
SZcdKkoqjCQvzktXfWRHrqaicQqTQYrzvITuxchAhGjhymo9iKcqgMPKblUPanGxpBI53JGVevC6
sK4MWPE51pN7+Milloh8FkeOqmG4U3XJFf1atprjEaAAML0QDXCA9+7ZfJjkRMHKrhg4NfqNUSkO
70Wv5JJellp9wMlItvqw3+nIhtwxn563PDszk1cI0PWxO6kLKP/CSXsUNAFXrs70BwsADXqW/xG5
/RF3dUPfw+IhuVgtUnabqfqE2M/emeo6b7DKFM0Tq1hzfO5rN2zgMRVpo5NQ5TtM70BjaHQz1Qk9
kX9T3+E9AHrHe2ZoWXIcZUAX9syL6TnkheAiE0kJUMzyXGePFrzP/PGOCeQ7zc2QVhW8AonY/6sj
eSQNq5y5PpWQbh+685BlbX0mwm7FzZxAWEFHD7GiXtYL60OgGiuAjYfVkvImKSMsNcG1fNTNGKUA
G5XIxUrLQeJNyMBor1Wrx4KZR0Sv3eDSGqETqjvMg/Easqofo+c75G0/uiEKdjDFIiu/4LVUcEre
7mJNr2F7Q8kB+SilENrBsofev/G1M/pJYmZqUCY2DCPUW2t1e21K22Z7t66kKeFwTvdXnuGmyXc8
+Qtbnsy4GkNNOuDCWj4BRQw+fPAERoHT/lZ9NnjKe/TtkT2Q1bviKhz6dbZQY1ZOttA9Tr7Byoox
ZR1+QqP4vet7buht7u+uEhV/rboN/gGgILZWx6eMg46cxfK3gv4P0/M0jaqtID9uO1f0i6qYPUb4
rRqRuVRNnVq2ZD+oVp0cwbGX1iBdu3ORFJdpEc/ccVD+s5ZfHwEiBNnyLj+IiyizCOp3tpAC1dxx
gPgzsfIUJGZLk2hQCn1dY4gjh1zLmFfXdFlXdxjBJVY1bc2o7Tu8yCAA9H5qEzxJHuszMC/Qd4JH
7JiSaQASH9hkMurmycX6VTzRdkV+/QgVWFxX5T1D9TsGlCWahpEq7N5/Vr5jQLQuwKBlbde5ULfB
Janqs2Lul/1Rwqvtfaqs9yu+x2zdL6KlQ8/FL3mKeViUOSvhY07071zoHDYgH6UTXdMYikwGXtea
HmkQcQVGKPFMy1RvmgiFTVqnQUYiL3HDhu7pbPhLTrlGtimBYBDH+B+zMx4chMT30W8soOL7DqPV
GIYjU9saAi6CbcYppjB8rnij/oXWD2oSiiGPYlM98h5fMVT1DEoB2UTWHOeLIS0/wT+zf0lRJpAB
jmHsow0u/OQpG5Oa0e5CLfM61hqypUYUqGHhDqyn3tbq2Xq00PHW8h7ZjpZO0iNx1BOELfSCJCTK
cu86odmrogKXIoLcz33RzvidZ0qZ1iGK/41ZuoKIXim8YddvDKRDk2SmxX5FEtjqpfaFhovk8KOy
WOaiowNtfZ66UmeQPq9JY7RqrYX/eVP/aMYme7y26s+eec0Foy6XE5tKpWaS1X2kFFvKOQFv0xqk
+Nk35H4K9q3uIxwsAoYtaXlPlEiDOJWRn2b5EqxkqQcgP7xmNk9Z6ujytCQmYQnn6yEusK0XK07b
Jc+d+OamPdf9bXNzIT0zxCrWEq0/aQb1zs6Xg/Ai7isUcyinpZ57pZwrWVKXA1N+GPi2sSpKdfeu
3vJpsaqW+KIfLg4t0StCrqO6Ck+oq38Nw69SARJc56bbIItWF38mvp+0yXB8bX7RnEhjm0FZJLeE
+3w+fykQa0nIB3nF7FWSOqve+FG8idgkK+YOBL1CkA8JG2BJYjRVpfiHvZB8j8SJ8vLQwbZfbyyS
EQXwtE0QBNSbmACzOP/QDcUn+O3pDrl6oK46jYkwS9vh6AmcZ0WXSEKnBYncZeaCF1Ljhmi++3sY
nRexjyQOJ/MfvZw/tHRrbZXcYqkecUUUTMmGkGdslQIiITbW7ve/4WJCXRiW8O4JVBjq88kKapIz
VSyCxznwK2NgFXTN3qWy8lJjO7+Lc+FUOlRHf6/kveSAdgbXy7J/iLx0WAHTg5ZQ/3OV5isl74sA
21QpvKaqWR6TXaR+mctLYv1eT/AWNhuRe4qEni+LO0qV8zIS5PZXbTia9/Bvs6eeB1ZfzNUFDD66
F1PhgpEmYrB+gUU4aamkqHpxXHuwwLPKdhZzl1PI/SVR6Yv1zkamjhDqst7B8pT7sYuRLcXUB/SO
+T5TKb7GL9y3u8BEl2sm/oT0qYCa1Rj5fI0GGGV6LbxcCEudrekDRBrCDNcgsIKuvw+5plQBWi2y
zhg4eK2CAClGce21PJrvqsdWpn9UA/YywYr1iR9GUid/u79aAI5TEHeSwUFssQsINndcces0GjpW
WXqVFRg7QqRB8biVa7cySq+n7p74UskiHCiCr0464HOcXF6oNisHucEEWNKYBN74fQP55m23QAI9
/qD1ChMvpOlnDoRwxmoELM64iYXhn0yde2/8/C6Ag/3yaE+++xeJRGKqKCFBNHKL5myuPM7RkyFi
xmvS7PY7kq8XNvA6zj2dUf0g7VO85SqMFbr+7dj2SC6KP1CspcGgL/ClwdS+J7A2qdRruMFQVnDI
i/Md/hWOv66ZQurbG0JL52+834W01nxWVyVYORPk93eZdyk78g38A4vdRawRC9JzHFqcaldKpkuK
OOM0z0UuJZaxyt9gmz3tMZxM8yUao5lav8VNhr7NOqly2TUkOEjVNU8T5CcWbX/ETdWqRo7dHu5/
4dxnXwJ0WNDYNzaODUFIrUwzRFe5niNCrZxLDOOEqnF9mL3m76mPGBjCOjlxIG7J9wqCKbIo8sfC
psUhgOfhlTXm/F4/uj3lk9WiPtmJxXKqC6nGaUwwjPXPQ/pXTQbkMh6P7JRxeXP+OFqYNN41bRJm
95Bwe3VyQXpBY/ZCstBxx2SyU5D3LsXsaiIl4dX70FCbrO1u/lXZCAbNmb2MANpDWe6MwC+kNq61
FNtCPJ8/rXNzNNkaJ0GRjG+9wSD6YTKmw14/jYYDxuMLjpovQdw/ysBsxTrXSEMCNE8E3SVNv+ro
pF2/FRNwUxjoiHFeQI7BpEQp3nfkv6/5sfjCkPzy1q14uFZX1PDtllSB9F4rqS1QREi0WhJiYqXj
5H+fuKdgbeY7J57bEVavz9FH8DMz+1kw2f1tJUBXd/o0cSSbqJ/eRIFkIsHI8fCFdqp4Xx/AXrIu
1QuSk1EmAiJ6FlwThjM7o7X5Sn8RdGwbH+GwyTyiQ/rt+TfLNdu1YwtIswsnRNhMovZKpjsPhzNV
avFFMOvjttNBIlJ5mmtidEoI30BhtEORuIkr4bX7tMUbB4QKQxB0zGLzRr2i9Du5wIswVovTiM38
kyumCLLyNv7biTenNWHRo5ZQG6V6Bo3fl4lmXkkNPZymm5MVg2GloKqmiu5B6JGYWeVn+zDkEE7d
cMqB9lcYcWZ95X1Ihrsbw0fQkqvnhR8USaHJtN2tEmEYfLh8CT2NZdhyfc6mrQ0sgq1khT4aQg7b
OPKBQ2LcpMBypSlQhMF2aKmJTc56lYSLZConl4YR2e3XBDjWWH0MHv4qWUX0dzNYN7jQBVrYDAPa
5M6+9UX6C4KRfNHwSXcsDlqjg6lGutWzjaSirbHQkngCMpURY3xf4cXNbwFnl4M2Tqt0WKt4x/yK
F2/mfXYdnbWDACWxUpsUPFVSQT27AKnTyMZpLbd938k6wF/QNMhjnPIlkKeNYLyPYMdLUyW0G0k0
APTx0fvJs/i2SgdTcmick3WWfhdwfkV62ZvkLLE6kU8/8dnOSU1teU0c/AZrAl3GpqWi/8P1tP3F
SueRZgPFtm81J0PtpPJbMaw+oOMh2/tH/CdU7SOxu9M1wDy843Lj/jpXv2p8Vzl5JfinaeZWoWav
iuLZj99NM+IOvvBQvw/TO0S35cmJeCTw+v0zK3ZcqcHpfoegbutx1Ty+vkt0Dsd3+wtDB61nI26q
2qDGFVLl+MbbLQEMQkw0QmzKMS0j57zKBPUFN95/Zk44CmhmFYWEfRAjrVygNjTHzimzgcPGGgiL
5k6m8r3ZXJxyWhQAMAvRxlswXNeS7uuTCmqZ3b5NlavvxhLtE9VgBwpuibtqcQezR/Uj5GwahE3F
O6VtEZ8HCiqmDfFF5omq1Cgo7zaAUqnUzF8ir3bZISCnwqAeM02pIzyYYBcmwEcljsIBNrEjGKY7
mtBd+PiRrs6Z6DiJaLABweoKsPaftljfQe3DOspf37WQfdGPXnsOmW51vfxGbod8P5R7/PSSdyig
IUzridB1+XEJy7aGPu4c5v4QOdN8KIjAEQ4GHyiV7kn5aRh61rhuGWJfZhFdBTuWgtDEMrhcyZHf
Q5YVPuPppCr5Ci+fddwCu5ATtkrsVMToUewxteXAVuVt1h8buh5+QBHCV+U0l3byHgYIPaxQAIZm
XDJywfPnsrqz0lIVXyIcylYXNW2S+Zj4sGyq0aD6uUvqtEp4Ddm8Ksy0Yqqx+3kS3nHUF7nzcPAR
VkTtUr0stLP7UtKHPmOYM93Z1+SBusSYMmzHeiqQJ+KNqUk30uK5qIlWiDIQOLCDrLOZ9w2Soh33
LRapEpfCFY3ACbLzoNPywxdBlOOi14Pnh9TeLHrnFM5D93hhVzYXou+qz5Tp+nBhcOkU+rAw21ej
lE4jSrn1EGErEcYOV8azmGrI2k8dl1r5FMoEpfRkObTXNhCuemM1TaOs0rS6TrLJqBWIpZ93DfsM
yv1jidoRdVU6PzGcf9tSxxC2GFn9DKSzRY6KzxYXqYZd2FVNmZ4oKXiNfjSCdznq9Hcg6c22LImd
7JDRZHyLyWBb3Wq7Rrn5Lre63RGg3NqMfctlxr6E4BxJQoGksNKWu3UyXzzE5z/8Z25ADFK9l37N
L3iPZQWhO/7DsFEXlJBsj6vJ/5HStD2d5Zfnpy1oZI5imh6CeEnm374879QDepIUjOyn0Fx8qE31
sigRz3Yx31qDNdFVaScC9znRcmiRLRn2j7PRIoNUxq/csXPTSuRHkNf16DCKlFD93FOe/SohFBsS
s9aSXD1kgnRkF3WGpkpSIEg2Oj5RU0enctRiaglIDb9G/e07PQ3wyaNVbwTpMOG7XURyayD0el4P
x4kTLsoExzTiArFLWBeJb1iwLyeqiwXdEU/c05+cduciPKPp1Du/ILbrkWyie+cHlK7ll18yrFZb
SK+CHX0MXwYV83y+chqhrPeoEIwkDNL2A/cR2BrIKyWIG6cmEZ0Wbtcb+LMHCyEbK2UTV9yTtg9C
s8+iUb+TzsuVFXDkG6H6DITu7cp4CRRwTztXvhk8VxCOsqsHgh+zXEnMBo7htnnYGWFZvU7mz+IL
6l7b4EnpXtE3dXWVG1b3jqSmzog+IiEz0ezkQXxBJzl1aJnoJ02y/qczUsoitvfp35elPgzbD+Bw
ST595cFGHMR1HciAlKMDtZWO2YqBJBiF4XK77OkdmEVkl+wcvnsUvdx2rDPq7M9DrzQYjXayFiqB
jN08NUTqJuVwx1jhV/HYEkG8kaFJoQIRy+2+FjUDZkQSXU+TBIWFhccJZsRmG+66ZSZxxsQwigLo
ymiN6InShcmy70xYke6Kr9qIHbGlozrLxDMhYh83U9eMjY4Ik9Qadj/3thS/8zNdRvjxlz5BWc4S
3G8qSNzYgDQDaINgLdMqVxOTVLYcDhMUa70afwARf9WIeQf6/lnoYQSwgZgPNkA/LkPyFOJwPiQi
rhA7tST9YUiJytLiySQ7+JGPTT7736X53W/usx3vOiK0GtccLgR6NbkQm+jGk/+wfqwCgQ/SASP5
vyHnJqd0nadPi/4vN8YLjrf7oexdjhtM9uTKMrSiMRx9MUpM7yxv+cgfp1mnz6KHqQkuPimm/fcV
W7G1WyxdUWP+6AG4OTHjHytonKa7icE+p3Tg3LpWgN2dVTkm4hFxA8fVtab6TK8NXX8Hnb5pdBh5
XKBeY0tIuIyOoVKOWbdmqwoRykM0cI6kvrME9ZmSu64K6xiFFUw97/Yhhmt0QywHwZqX4VWUzhS8
+cL0NXPU5fbD+EVTEXBJBwH/j0fqBXBEXmHwvCLM4noQIGP60+/iDg2JVPkVR3aT1lGs4flV4ZoF
RBgR0l9kyiKLI2sAVSPYCkrJEHeoPbJrZiJeTeOwkYO1UAaE6hVh/0JCELTqv3YbzCK4EbDU1F/U
h9RLjdVvJYKfRz36rn8LYQ3jlKVuC9U4fNNMFBr7JQp5lbQeuzFMixWfs9nAJSYwHoI7xhh/BRzN
wLd90V+RsZ5qX2991DoD+F1H3XPgF9TsUzDHHGDN4yI+vwjx+sxwwbwVdvQxqpfiBwRQSFkCmmFD
1fSOOFGqIBcdf3K98Vh+an9ttQJnfInaJy2IrjpOa9fpeCGCtufIfriM4FNUvGFdhd3cKla1VpAI
Fd10ExaOj4XRnvBmRS5sRxdXWJOPbaVOkGHk7wC7sYv/PInbE1cyfgvDS4Wr15UVXXBv92B6swTo
ZXRwQxqwbbg+UbzXBPeANv0lQ3vjL//P/0F4cKLtyWQrQ+8w+HQaJv6ppuirGq/ZLUCT5+kQvl8k
lfZLfT6tgluXHxGLja0VuIEcApSXZdYdKRBZmzmaGztOmrmmPmjdO3hfYNS/t4LuIJN2IS0YynX9
T3x8XMbQQs1EHq7o3JjdfFWotKFZ45te4Zp4jclnM0RB7Om16kroqatsSOziIOA4Un9ePSoBy/ot
afYvGm0Hn3LeBxtAvv8n6wIujaImj2+R2DUod/0hKHgNqZ34vkVZAeRwPiNnudBq0xpYIkZ3WX2s
RD/x/gCr+v6ZL/Hgkk5yiW4WDsMhd6gMG2Hzu02eILlvoPWavjYarci3nj5KRklT4Czxv+lrYR5u
WEK17/vAbQUe/WeAoG89iZ39m5VrozxUVJx9QxDN62zJlu2Ia+yjOo9evZZyRhqlt+xrtle9RfhD
Vbklt/H4qZuTXhPW65M1v7RqMWLtP8HulURjnFOEnHEGyQV4n40yymXQJ0y1t0Y8zxFVK62cBS7A
rwkGei3QHaZJnheo0qrIF9gIhoFPfuqNbRnUjLMvgGnMQ/zHOpoyLjiEc03Z1I/3AvVXpq+yqpZ/
CffhCE8eymLf4HItEddC7a8DhfbROj812Kq+tpNW6TfwelVPNs4mcq2mVblIyZ6MKJkxKtN0oV10
7KKKrnwfhi2BhkYbQiELo+Dx8XUhJ0/DIrpswh1YDgP1cHpB/ih/UxhEsLwI7hA1ln1uKUcTrs+3
zK5MozFWHExVPd4xs5vZON/J9D+UIE7msChhAyDm0J0x0rdneZHEw6SJ1xVp1ruIrE/3zlUdHC6s
0czRI0MHnyOj0yNWm0hZG22ZoLbHTH0a6h4eQvZTm5G8YR1Ey9GXAFZVJXW6ev4tBi1oSrHU/nuG
HK33bGeIsDV3aCabcg7QDkuX1uOXgjYfxAoVpSU1AbMU70ymWCdmJeOZf9muGNzEabyfSMuiSY2V
Gbe101ts4HiM+o1pwf7hrHXTLTEuIrwSO8OUJuR6nmI5ju+PYsLKM7zVP5NAdBmV79cps+XM7D6r
BPbOd+/3HHk9JSkaQEjff5DBQG5+XfyNV/WLIgHo9hfth1VeXULSjzi81Z5yrc3K4QGoFh9DfUux
pEumcQgPpexTT5KhUkYvgt+gcnfZnrNKN9HrHt5tw0g7V2lQUCDZzvw7nIxK4wHqspyCciK7Z9g8
YhkGNUHbt+Z49CCeWM0naSPewHKoitBey9qp39DixltnnwnfQNRqWGdcQZK7jaL5ZETI62U2Kpzh
qYWVIPKOQAcVg855vsSRt05LsWzJ9QGp+2LFFqSi8DwSeRQM9oLYugc4GQfVVsRc9AiSJkNG04cE
M5WsAU16LdfKoy5BWS9h2klC2iWxVrgbCb9QJEslVQtpOrMO7+4e2xtNsK7AaGQPZHFnZyEeTUxl
3f9DUAE2+Fo9wI/ihmiomHmvcn6fle4Reo9cfirR5cwhQJCDc33hRwzrzAEYsHhDNPf3WraCm7Ow
pf8hwRnZ1hnVYlsEbScNhakZuqsTfDMHvDDafPwImd/8um2h7g7s6Ofr1Zu7848Uz9B87GUjcw3i
6Ui8Jgc3YIKj9ljlP6WVWPzXi8eBb+UYAGLPEM6w6PuQ+el9TLWhrZ/Fh9AHw1AxiOGJAtVFuN0d
wVc3SoNtqesq1ZqN/WNy2BLoNzeXM1GwWPDry1iwny9BLQS85UuA1934+FnoVkOEqBv4eLDigeJe
HerXTpXZX+xWVFRoy0SGlxK2zaJSmMqG9+BGOtJbSuLWS5w2jYvP9UWIAOdpEmoyyNt/hwfHWyqb
jBC49mmLFbvCuBa0vul2BVmv5t8yvVgs7I+ZWI+YXLsX8iABwEokybA2jd/SjB5eR3AhPWS7vyBt
cRhUkSyZTUK+FNJUBCUWWFT+90oiJPjc9ns3gIpoV68dP/x8eNmaB1H5zoFdQTptEjMVEAJglVZj
wtLtoYWRMm4sdmWj72xO725wu7ycU+Og8V2BrUY+jXLddTexGl+mjb8J0JuHu0onbplTogbkeez3
nSfuG71jrljpx959SGOfyfaV6+4GLRGTSMMpvMjHGvXqvZPDs+057sGATwf3pQKjlpZHb0Rk3cTf
zPQfh7l2LRe1/FYV8YknWrITk5pW4oKiRNy6HTyY0umqR3bVjxPGSx9AeNCHUDVbZRkNIvI/yJVt
PlSVYMk5gB08c5o5H5J63sQQtYqxl9lE2anYVO3GELzdansHEu+znKr+Mrk9h3ZcGAEg5CawvLtI
Nm24L11pB+QIsEtJ4Kv7rUOxfWfPu484OjWo7ZEXGh8q2tfXMXsMylokrwFDO7UCOMSMn5d6v2/Y
zsAD0wfkrZchfOC40XAlO//cZoQ81+xTN8cDqgEvbHbKbHq/x33ewZFZMtZ393HhXdNG+m4NQbUv
GqwZYgyIltUS82tdsKwQmZHHn7LsUrwhUrZ2a4uEe6go2lDwstOQHYhbgNNnxKs4ZjaYOvDn0gkA
+17CFRaRJLs9EEe4gcocKq4cEDzisyn7htirvDJbs6DDQq0z1vxt9ulLfpIgghNbngglIHRCIpWY
8NVJPaK+6CKR5rNohI6L/N4Qr54Ozizkr3MmYpOjfPeY6j0JZFAUGYsFIfFROvaWfTCufRLIy6Uu
o+D96AWqJyOClBLwUeBt5bU1DkYQkG5hXjFBL3Q+KLRGtPI51jwNZSTZh3L6Gfp/ISYgRYE9GGHT
ZZztoScxCQMHHfIRSAMofckKhZRMBI2cB5fqTGQl8Tp8NgxPD0+INsbB8nw2YNGLMhya8+cWjSwv
dhqQqFv7VlqWXtuCk2DcmM15O/quqhXi9MBVtoZ1AhY0WPzAoWFDwFDhCYn2fDvQy5huJ6j3cukJ
W6f5NBYNeLVP65i1DnvcpH7yh6IWSK+LxprIf2d19JeVB5AyRUHPnbypwM2Srq0gFJN69RxsyrCK
+igKos4E9QtlEEX7psfhiiR0QC4hYeydRhifyXWAYuWMvmQddpFvBRDOSAkBAsjVAS/fjfnQlhis
FSJu+3mFUwnOQZ69YZc77Z60zRKwbPh+BYe7Mx1RrvQtxHKkDaEF6d0BnuiBu47Vv123BoEAr/5K
MTWtJQ81zhZgD0u07B49QgYMwpbi+VV5x/Hu/W7OSPgN000pO7Shv4QAdQoO16cLSdSvdGa007wO
PmJU/qpQGceGsCTBViIaohZDcJvuSudUMkcv512YziaRMBHAt3tPWc39Ox/F6NeNBL0teCfla0Jz
IK/gSs37aVy9SROlAPxNypPk8MvubuzoRDWhbZdjAhC14RbiCijJ4rOZehSTOr6k0y2+mU198Kt+
NV5sDT6jYqHdCunQrVB3UUtYXwLr7AaAs1P3TjC6hOk9oP+8wxTj1fIFMpUf4uUMQz5nxhV/87Mk
YeXQCMTfJK2j6Fb+fxP6hkfpspEtw7gQmZR4TjoyPG5Vxq0s8WpyA+lzVUQQvuTvRiS4MDWzuR+L
VUOeJmyUA6AC540XOrwCOS0+i6WYnowsPi4VtYJnaW8l8nlDksyv2Ndb8gNO1HaItfO5hzSAv78C
UPvUK/BZ+v43a48XYCAVs94gwFxtkGspFdmpj3h36z3DpoaYYrc4P4QZiUtjjyYYuTtlkEgkK3+m
eSXUgm6l+t5pwV+JV3eV7fZcbZM+dQDPQOi9MuUmidKXb4F3eikT8ifCpN+whgZ0WlGtBm/Rw4Wf
z2ntLX4kzFjMVe6XWI2aBo4ylSAnbT220BIVIc7NOyF+dzsAVF+9X/Bo1V8Dkor+u6qUbjlO4tKI
ql97rpXRkpJth18lgA38qkrSQgtkmfMgVWH4sfCFcCUyGR44o0ELweCI+8nA1Gg+//jdgsGBKVSo
2ld/mHNiBLpWnIYu+FCMuZYhomkJQTQI0IjwMtl7ojBnFZTjRfeMjl5PERpr82oA6A5EpS8Nx/8D
57c2eBEDeI0+wcMccyglELSJpKhZlKi5zxkQ9lXnVV0UJ/gfl/mAozq+3uGvrFurMT1wI5HrjqRL
eP+QVpjKdorTscTZ3Wm91Z4X1metDGBDXnbng7j0i6tGyrsJaZSyLdtNaxQ7xxmnU5Kc/xgJT8KO
skRb9Z1Gu+Q4c2nfLGUeqkwWLfIJjDUvkuAaWxcD3MQk8w6I7D3UbccQl1uJMiEE2xtmmxLPlLCs
bazixel/oaKRfQTue+1BQ3XPEa1GqfBWwVoe9d36sgBRy5Y9sm0z+DONWWkjv32jNhq7NRMR40Ng
yzcEdvYfbPIqIVKTjzPiautBpVdOKJxVDLS98+v3GTfuHcU4eUo8yv5wHDSN8MEQ9Cf3SxCK+Oam
lQ3tldTPFnLetM5Od3do3Q4YEH5BSkfZ45lfZCFvroUuY1c+6QpGTrpLj5iK2AMDq2vE3Xu0Pkl3
4uymhcixVpXcP3CNtAMbzV+d/1sSmUT5047hy5DPTl50rTvIfx9beZc2qJtMJsk/HjtPW+LY1Tvh
7Cat+o1MWwHwtRuBQnK9m4Lmrrn5eg5hrjRuOOKp/8G0Ovbkt/gzp83OpEg91z+wkr8zZOvD9slp
Y8BhgeVaIN4jrrrrubAklZkG03l410+nCzD3omBk39Q36gsQ89688LW2diROA0lBtL4SFn/T4uKl
h1qdyiLbJrnNt/5VmGClCCqj/HMEaNzyySR35mfqWoK0PSLfsMRuAkEkdl9bTukbAMqLiYqH6fLQ
0iD9FYmDjbXTNpVBWaJ0muXQVoUT1jSghQN6yAm1lj+RSfFvvVids7w9iwl98WhBFSfMZP0s3GDW
JVAO0eyB6ZS9qzAmlc+TFeRTZHnCIFBXe0hbG1FM19nRPxqLHi8cT+pvE/f5YJ/4Gzcm2HOmqqgY
Ll+nzgOi+dNx5h7cMkpXie3kZwNBrWz9lWcTv2xsQAo/pcNU92WKju11qLabfOakbn5xB24csV0l
goLwuI4+OX/9S7LdV+IDpWZT60dZRwzLS9XTeyvjiTt9+Buw1fRx1bLm3sdOqI3U5DHvWa9FIDfH
E9cflDfRdWVnzBWIxlHLQbI/OhmUK5iNwFUu/3NgBNaOnbMMZaJeJaM/8t8eaCxcqrQhI11wZvYD
3HFf2pUrwSbOG38mkmPFAKSfh//mx6hpjGJslJTb7uEjbZw2FaG7f/6I+tIkRo8YItKzw+90IDWj
6YNvwkZFzNxHpVsPQpzjotJr8XSBgAsU+cdrmDKqmNL3FhypvxreMOx2t0osFqzsRPBSV+EnSZjh
n305nfYNAObl8mS9vR0LgASdacQevO6WSlcstAXgTMhXgQjCO981RogPT2WsNfx0KXBEZB+aHwm5
cW839lJvvjCiQDUeC3nRzgFR8IF4YF8ZIruWEfKOViQXcsedTWpKm6jFK5cR+OOu9GpnWgpiiRT5
fy9JmoMnmM5D4tn6PtkBxPptQsAoFuXflUMUaFR2kD7xuZWtD6lESudUtI2ph7ZdRUWfgcGf4eG5
KolUJyD4wuKY9Le5PuXo6oZYmZzlXVQzjeeWA4ujDclv1AOTXj9rzQqoTIUxdz778NdsA4U5UeO+
ePiM+HvhaONTeT8x/kFvuMv25KRR9AuEg/b5Mx4BcToZdWxAckbTOPsWT/0bfdGbTGxjxynQD2F0
fWqq+yrTPiyDTYzaEkrRdmQ0RcMQ8Ea0tLUQkr9i5qVYEniFmLhFBJKkzw0wCi+YdEZouq0haXDH
DXTTQzpc/ZnLi9huzqxMf4PPJ4fR8mhRjDa8wsh7z9T5zaKpPjGMCig3BTvN5WD0d45bLcv8IYJ9
aX09bzNS+589C235NsJOvImsBvOLQK8OS4PAvwUfSZ+pm1JW6efgPvZt5gsFUsUonO3ouOH4WsJl
bUWW4qGmmnM5x/YnxnaFlWCHeZThFjz5G5NXLxGbpVHfg0YYmerEeWbIyx7ka782UZkWD4Ov8gAc
IBK8QyS1lDBATK6u54lxT/pKjCbEfivcBLMYENpxjvnzjF6yptrLIM+l04S3y7r2CP3IAeYDNLmS
RzSIJrnYvEjQ/wEhA3/wFbeo+aFv1PhePtymVzXo0Az6qgYBQ3PnYNoqQY3II6FfGOvPU2zpsT8a
pEeOtrtW484TabFsEERrMWX8ycP3bXDwm0RJIy3gQFlyAxNXSePURN6ucWUH9M2DiGBFDfpEa5y/
VDO6jGduCQ6bmAdfs8v1Mfb5U1MSjOYp26pi5UHKpwmIkHuEkvnvo6I2qM73+w5Bo9b7C5kedlKK
+GGNoL9aIhbcjHqPRLDMbrZPi9DYAtFIW9Axzv0X3M2TBamnPajfWGR63i25NbE+cqfzSYUJsYwO
KJsM5GmFSpNvuGqZRipxdBJv0IHClURkNz1dvrll6hcJZ9AvvyegV/plqp+ALvGAxPUNIaaIA/FJ
JJTOwIH3MZWlTnEXvRCI9Y4nPrJ0wcGrXbasaGoB/2ljcsxMkG5t6ZGCoJ6xGFgiOY550xm1lOa6
BhNicykZ6Br3F7o5jvlY0qTeLdDckMUc8Kf8sqGvrVs8rycn0mkHOvsNsfHfGr2i9nVspSXDgv3z
pv/J6npbY3oL7/GQvPZ2AVqLRPJaBpO9bl8GWk71qshNoY3Z95W4t+jzNHB4K6Raf29rxfBp6A5b
lY5Px/+Pv8UQ/JY/Vn4IT8/9YHN/2FDV2LKyRF+oiM4XSZXPe2IpsJry8KJj/i6Df/H/wElm/+79
UI59Nqq7zccs1VZClyFI1iiwIGpsUgLs9h5QH61ZH8qUVOPW8vA09+GxX7sr7/Evd6xrOmSfb+fi
G3edEMlGhMpEnuwQJ664QZzPWuTjGUKC4z4YPndSDwtCp8HAJBpDJlF3sdbadg+zLr8xArTxSjE3
U9494kx1TNzd0S0aBKYOeA2CPs16TCbD+HxAHt7dsApgzDR4u03RLSaDZnnxbXGIbCDhYDQJRZhn
4i8gNSdcd6WLxqt3mMQV2h4+hMksq6jobnjzseh6F8q4N6lk1xuCnVoDwRVcIgyqSQoRzVBoW6i1
czGoafWfjUroTKd7R+HCRX8LIRxiTXJcyAeGM0uYjqHoNnAxLGnx13DWTNN3QAbzl+5o9I+u+ot/
uTO4PsPviiySD5v/1xkuvcxbAGYjn6cgDA49BEQluf4jLVyFtlZg58Yrrx+n5wFhH0XmEFOYUjr6
BUNCXcDwxRTci/M5e1T2m/RWGIwQ7ZkvWFTRKZD2P1hIwe2qr52PMwPYGN7bHTksBMgTHRVJKz7n
wuw9b3TCH3WceyzIUjkmwDGRy3zYUui8aKymgeJO0sCWKzAbV3hl6/dcKYFKdqbKgA6+AlqDa1a4
xNgAq8kJDuWAfkHh0HvuL2xuNFZbveYWL3lh6bZC1V7j4nvx/WYjLTw1EfJhLzAEonIPhiCwcbyq
CK6xOsR77SC+Vk2AvCbk4GEZoscK9SkGRWAwVfE8SSnQt/yoCRjPq1a4Z9VCyL6QXI8LIaqNhUEy
EHIrby96J7w6MKjBjkdyszlPBuV0S4BRxcgg7hA5XMjPMArevpkvr1Evt26OW4sfsherUu+gTNvp
67J5Hd5kSGldPCEAx5nvpGqABgL4S/BKahWneyJvpYiTV2lumLD4N5LEsc8pEMiEuXjMeliaPSEh
99j04hpIvYYBCkc21vYqG/bB5zIEgxYqTFCB5foLIpO+133+p5bN0fgsdj9pkc4tVJAJkLZ3w+YX
DjuEGMv7qw2nvtUgMIE0gA3y4Bl7f20+1aTiXA1VC0xxMOjSSV/ftXJX+ivzkWztSa8pNv0Byb9A
CdeqUqHnfFGvylimZFxAXnWP+e0lDClhiOLUQc30K6Zpzq7dCGulDumEtyG7gBcNl7QG6vg0MI7Y
PYqPsxUycsPm4PiGL7RajT7VU4/LXfO8UqUfHtatzNwsnnHt8TPwFR67vJFDjVd1Z4s88eMPq9g6
7/BfVRBueb+jCS4lLE3N3vQja2nlsWFB8UdXf9RArLX0R+hmsGOtz0lEVTJkO48kBPwLflJ2znZC
392gc0lP2MNJq7ynPsLUEOPRqEW5dVDTCNXQLl5HMq6inCv8M4duJcqy2RZpFt4rE+Gc5QhNT3AT
mVhUy6MXS1sI8biGgz88K0LB/uoHmBJHrtCts4xQuqfCFASLZK0WvFntb2naEGmEefjM1SfwPq1E
5E+WLsKCErFmG7sJW6B9YjzT6dlPncvvjaQxx1cuU9oUdDRBSlVrQ+qSNNoku9oniaY2pObRYdpr
qxm+g0d2+iM1NgHGCYnms1v81dauUVN8x48ifnZyBI+TF+os9i/oAPqKbzlz04ynZied4+pUIrKc
//C0ZeeziFFdpASa4lu9CXnjQwgDu4aK38Co5eYrp9DhMPRQyGA856h64peaXelw86M3Zi7dlf82
jrcWZlfSzPGz+tdjrsIfYnD3gTbSEkOt4WdVikXt7yMZsGrwzR1X4eY/t1Lfzh7KZvtjOmqiQRVe
ljFuvwEdPE1SAetz2onH8fWj6EHV5jycfdlfIeME1/6srs1ktbrhZ6dPMpu3hS99LROGQ1k7L6b9
pWpr7PTeMcbPMTyy+vslq3zFd10RBe0ptHSaVFCM0sCxh2dAJArQ0hgHZ0Tyvt6/tN/pld7tftyb
m3+7RXATJt+hzXZHc86aVvXVURhFG9+rV6QuhZkHLRvzbDLqRBJ/WXvQDDlN0ksI/TFJu25rMvMP
4yBwhCP8bqlRvC9eS0rUQICYbtEKw3ozpTtN+R9D2gFrqMUE/6uNkphjXLK6w+gID0d5wJxHQsi8
GphopG8Sfo9sCIowfTXgKhAAyXq/jAzCX4Ij19WwU+fojKsrVvKtAHNprxtSvyvTMmZjP1XSgvmj
xGcyT3uSUzPxUKCpVauipiin9+DU2M36p6XgPQEkzTKjbBXMVskvwfQb5rD79loXogoFgWkjOrsi
2Tdj4187GCBvudRYkGcZxZV0AYn+agEJr90yKVt+Dx1DofV9vvhu6owlRWQJUd5ztMNUPiBHQB8j
VIsYEoAbpw956RoHPRX4bCF2shTO2KunGsq8A//dJTh8lEfLI11P+OvMEnaZbs1Cq0I5/lOgIqDN
dXc+Cs1WeouJ92NhudELFsixw4hCVrsmQEJDB3OHshUW2hNBzZGmi7CrwzPkaOgR5a8Q+FQrt4mS
P7U6dmAs75N4/56lqpxVsuBwn+ehgJViUfm1HIEjXvMEkZQoMgPtm0UTj8vZXgrtodMnqiCHYAhI
LPKph+9ePOZTzzKT5+OM9eMknu9kg8mfvmGKqwYDdoJWyASEV2pyt47kx7mB/laO2G+p19m1nSHD
SPh0kmH7DFuytGMDB59zhujtsCttfCm2kxu73Ph6O045Cnc5OfGLexnDyEtag+djFWM05Qfk1YWq
DKbBAhwxO4pFEcT6TLRxWdKlp4ynh6ONoIn9JWMyn5qE+I/eYs+ftZuRhPQr67m2eXJOWHRyRrnX
nDxeI3OOBdN8d8XnrToHMsNx5jNls3/0tXr/TghAP/cOve6W6l8ueXiKfFPqZrYzW6z4F1DC18n+
0SSvdEySWyNAH26B23DPWbAc7G/JP9dfJ3uwyTkWkLY770RjS9JJ4X7smSeBvPPyOokTHTz8Hhio
Nhg9KHcVFx14ap/IiyNvIa1GTZV5zKKGj8enOUrpuePhU59b4MMNS035UodIJc0269VpssawnwaQ
daWO8oErdrtwnu077SPR0OCQw76n4L793LKUn3olPgDwZBei4WV8VKIRLgEEoKOBI4s6R3/LHlqF
Qj3Za17kk07ECCjrm8lALev4uyyhmPgfOlBO6eHEuk/vEshPcRrH0S9YXlpy6iTuXZLoxYbMDAFW
gaFCB5bsuiYpYwM7SkqQ6gQs9uE9cDHTa1JJqMyj7N/RQJA7/EUuHoMR/Ws4qN+qikhc0XT3lPv1
tFf5ez7UQI4/TM8B+dDd1Pp3i7zQm2TtlWvxIwK8aQ/ug+cKFAzRTFYkoMSI3RGCiOxSVItzp1B2
f6jJh6ET6+eRmyKB/V9ixcLCSjRpuxXUGM0axx5oSXvsl9EVcffFURpecwBHBgeFz4AwxsLu4Adg
3vIoIFrwyjbkdUqBhxeOVNlFxJ0lwPdz/qdqPBJqSMN5MDoUNr5WsmHzfX/RnkZixpAPReuRWxCo
Prhc7Oj9Lyckc7B76gdIBUq+F9NcpYDTj60Qz06QlMRYjsp+1a3T4ATgt6X6feV2y6zF5W+vNDMX
7qQu0TltScbh7pjxHAa8ORJ3J5micH2GX5Wdc5kF/3bflgpRnZNbDpIHijucpcbhmqdLoipdLVHV
/f+5z/5lWdCiI0GMhwLxhm3WHj8OUX1UUYYMS+/AioSDHB8sde6RAZuCoGAaDQCy/ytUZVIRqVth
VGw629JJGlbb32W7rOFKozM1d3K41XCjxE1evixUoRkGrsBYvpzrHf+g0ecEqv5PApo/mIWXcjVe
ONfnvkKWfzpUBiGFYgXf98oiK2Fmj59OTyBYlJRhF+p/Oav3PNmp2o55kWGijCAOUbS8oRBMSx+d
VXvXRz9Bk+RqXOJArQ3fTOFbWeEI/Qd5d9cKvcJCsXUHiuMbQeH7piGYV8T6SlonM/p1qv/rXrPE
VDRnjwXsHdjOI51lhRUFflyJA8ovIPWif15R5gPRWX4Y6AF1Sc5r+F7M0bQy1oBwKQ96lbMvGepQ
c9B7PiKoDt7hPt5Q8R/Jr73CcHFfnvnbOc/KwlKPb3D75Uq+mKdHRnqR32QRRe2bMAkgmsN7agJ5
Rhrcq+W9ZNdpNUEfrPHlx4k9XwL5P6KFheftIAKeVYR+ZpHFCbe/K7rGuD6YwGHhp3MC7qTGhn0E
64hpX4MGX5Vx4eXyoNvmV0ZrKNcaGfUHQY1EjYYz/zeYd2YG8XeshuBuGbKQi3s1OPXQW0bcXiJo
GhSfCg/ofynbUDRFxZtG8crgrl8qvW4ES+BGnbq0MORZNUdCsj951KdrFjGa+1FtQvRyfPqojf59
zSJTXiVSDzN66cKR7kglnLmPDGoxMMI5Fwf6VpVk5qklH0g/11eGdWplosX0DZarv81HuBgIQedB
DJfUhkdFPW3BPjIML9MdTOsCMiCIj3X6f12WAqp1zvW046Rt0Of8RpwjIPKxkxtz7Jr2D+AlfegP
EpPZMenng94kEAyiXuoccQnGXFZA2NztypZAvXlQebrE839GQo6wMoSik1qvO4xSxgSdEMDpuYNv
K07wwpSbZvm6/RwfJzkqy+0UUCzyXtTA6ZJs4YleLTxYyq3DlextrEZ9YJKo7ze6j6YCI/hE7Lqu
evPDg7ezxC/tjCXc4oHZe1/ubiay4RBuCom0O91lXzZGNTCHJWGAPHhNsQRiaf5JUPhrEThEK9Mb
EjYq6Pz1M83/+LhCesJy9KKdkLhIwi0VmlTEAMgcvCV6eDA06TSysfjv3dkf6aYA3TofLGZcpYzf
axYdO2DixLyyvGlFH9PDtaEaX+Ftt4NQnrnBqWBBoCXR2tBsGyRmOhQpjr8R3TTtkVFAEu/CK3AV
hOIpA2Y73QbMrgD1sUgPFe3Mnx2V//OuA7iO6Z+DI991Be5Yaa6hqP29U5ZgL6QYr+mF+1REJqLb
nx4uIixEbfDSbkJlrDacw6Tdhqi1iBwqCazexC2G4N+od5TUX1apSPVWz0dzJsUP+BiuwyyCbpX2
wh3Y13TFnSNPdC6iTlrgO8QOkAStIjxBahJvyP5MiARCyn8DMbnXz1Tvln8kC/MC3UyrvwfxpAg/
tyvBA0pgk9l4M0d1feSHi9by4gJc6U0kUN7ehkFBXwgCetzUwbf42xVMdHHKiycHVCtAHB6s61t8
oUk0sdi3SihWMT98xZ60fG/HhZuz39+kmUBNiOR3d+TLaaC9MSS0yPVuWHmgXI3XYRFPj7p+LOw7
sadyu4RLYbd/wVrA7lWjPJte7Pg6sMgoQhRbzeW9UVl/wOYG2JAus5UxAXKgetwso4dblQy88kP6
NpcIG6eYJDkJasmEyC0kwsF643tRt2T86hjPcqyeouZRyt3OJt9E1A3Rd7Hu3Ez6UxwfTDJpexvg
VjxhEEgMoNg8vWr+mj7FirBq320ZV/kO3IeYAXXNUj6Ba2rcV6IQUS7DMdSIeUW/o48UqAhzsX8d
Wxi62Dzp/1ZEiVPbpQ/AGa94RTz6RuF3sb7qwH5W0eii4zFig3rEXXWXOXdd4qRMWUXxc/V8UsSc
xdKSUOMQ4l5/2WN3Si0OwnDDlRGyT73naPlJy3vuDF2K/YIe0UxKX3MvPOn8skddXH9NYp87KvS0
PC3//IKAhq3POJR166BA725sfg+WSMTxce9/az2lW0XkutHmR916tny8AE79mnZ/tksaaZDCc0YV
YE1NGoS2qJg/IS5/fp0hh4QXro+PPZIejWHAW8PWRzYcq7TTodOs5GeEGzR6J7JomH5GnTHK/qAl
uCukfdULRor93t7hc6+6eugsImx2nvO7zHjJXGjn2s31oaGVtJRPlZ+00LD8RoqeLLXCq8KyZhua
Di547sx3rOtvRHgt/yeg1RTare3Zlc8vVoJ7PYD6DoZ8VMmWZ1kHu2wIomPJY5ZNgXxTPhsvsZMv
fYuD32jYB2ZAb/L33S+TJsaW6D3JxfunPuCpx93/nHkMBfJxpe49Vuk/iWKWqILvGo9B6fjIATpy
EtnarnlVRhFmkl/7iYod8FPoxDzm+flD2dqokHnK9TFN1UO4Iu9i3DiuziSgApVWvsR4R8wNzD45
EijOJGQvwTHrCrdH6OLlLU3am28wVPhwVAouO1L0Wyry6Tez1+EtylaZYAk5M2WDDVnTgpL0j4RG
W/5vwXEc6ZS0oNU5bk2O6XAnxXRvktQz3HL/z8DekbPiAXSzrAa3Vw/NkBh7WwGBlaIuXR+DyBj6
0JvWoAxbCKByAppJeJ23kApy1YlMoNAq2ZPzqFuxQZBgd//+B4b6ObJzTtg5YWiWCOm73/c84lmy
fWHhHURqe0maRXUXGOQUz4yyueaMKE4YTP9PaUTHRSMauEYiYR4pLnj1D5X4waVDqh1acw9xHVGZ
Jtz3dZ6XrVOAv0oTgrXS2i0E9XRUVBkbyqazi8NArEWa4I+V5I605XtNDqDeTqCIz77fkrIAJqTY
XOsjaVV9kWAiec6A5JpUaFZCAFjtwdAqIWyDQMeZ8obRJDz86l5tS/ox9xzg7sFyKKr1ZXSdJ93O
+l2V8GJEEIEtplZ9M+MH8sb5NwJ/dKUqvbMAP4uc5vLRfnkXGclkHa/oy981naek2tFP4x2iJyHv
z2ztk9PCplNbZ4CCUVUwHIJOPsMZRMw0PxzJb5aEUBsqDueC6d8nHmjVteyQ+nj6XrshMNe5RCJd
W1q0abx5ZO8boRQ4Yzq0ODWSd9ChuDrw3KIdS7oZmmkBN3Uy5Dfxq8sB3MEuk8eV1rtRmhbPKJ8E
EC8TCz5dUy7yiShGPGPEIom7v8oHh5wL+ZBul1GEHvzzcqV/oOGctNBEiREvKK3FN8tQ2O2L3byT
ZLEoNOZaoJ6STva57qN51owHDx+IdA6tJ2D8hvriPBMmZe4PAwbE0uSS2W6F2IvGvs2DyMVRiYfh
G+7uT3mGCpIaiqVuCReJjadKv1QEw3Wk4z49higcHEpJEUvScSOkk73cNRj9ruibFjkDBn4kGBfq
Dc7cWysR1GRY6tiFjpIGMKkXA3xJGVuI7Tv1f4n3i7mtIjF+qWdHbAIk27LiSvT3DrjfprAaZoxz
FObpEvvJM8anvsiiXHMzx/aOoIabq7n1ujpMSz1ayZa2XzOUp7QM2mqu5WOnXYlUKiR2cMigxzat
m/Xt5eH7BIP/XFT2vugVt8Eu0wx3hLWgCZyu5Qrz6bV0lRtIdoBV4s1Tqz0Ct4ti6m4sTYAY+7WP
sIlYqbKvlxnkLjmIicicsbYGU/waQoINhL7RJUuzwOWXI8c8r8gISous8lTlJ0H67nRymLtKk4CV
eedBY10nU59hVwiw/HUVpMPzYYcrsxMt5IratlsW3LWcHky1KCFbAuBxrZ/tULQj+qAViDJoqR24
KveY/ULUvo/ZdVClL6LEqc66ym/NjsFvx/QCd7zJ5UlfHZUpqBTEUbVaVxnkpGQm+xccka5g68yp
SjmJtsQ3wKb4D7YyWq9BxTgn8Yv66K+qfsNFlAjQrHGR3VNGWcn4KHAC96FRz51oiaExc7QBPk6L
QQLcYtKsOB0D7pkuqxXHOU7KqRzffqAtVv8Ho3Jg7c945OHA0aBGm0d3fV4yvbV0Y8wxybWlq4Lu
z+6uGlVl1eBabqIDz9hATSPugkDF1CRciYK7JUqOiS9IJmpvwx5fOriRT6bXP4TBtByBpXpSep5+
d4cyvVm1e7TtK6Ncx8+pnDr3YL+gA7SFZ7i1qzCdxcoQxnme2QxuyAqJPoxDVuWYNxpFM9P1oOIX
/rX7h5p+H+lQ2srmNkYAnluuZv5s0xC461Eou/NMrxG/JyL8vzxwmfBgzxAPVzl98QJVKCC8KH5v
t93Fp1edJoIfGr1NJ2lx0COd0xXeGJxxK7HPy2TlYNi1LOIPjpn41RsZjiRJnf8aLxg2Io2fpknJ
QPGtIAIQxt5hdrAw4q2V61eTMMym8OnK8xs4mIEa6aUrQgZLNuFXXOMSs7A4dWL1y44T2wG+dbOz
PmaTlIOKNuj5cfBTJlFMKLk6nyXxyZVr6xYpe8xOfpllipFb0DBNNAxhWI6AUQKl/Hr208/emTBi
5N8/lB7GcMjpl5ql1hNPYYDXjQL2ONcyHfuUHBxwBDZs/QJVJHb8gUmMGygjmF6TCHZONVvff/oT
pWeIW4ClkOJPMb0BzhM+vh6fdadGfaVsxGgeO0p62GoYRAv7J2+N1C40Jp2STbBavqmq+v8cGvMt
4qYqy1++8RIqiQUmnBCjw8aIHWzn1Ot8x6zuMDDsnR9km6qAYmaRs8OTa+9xECkwJdxozV2iSaUy
ExU6zYpbm5Eo0gcPnY9QdYJ+8e15mTiWzJSgxa1qt+VA+/O+hZgQnPKc+NZycQ/vN8pMLtwxzQnJ
gUv34QQTVC8/boIxS6lsCo7NIWf2RomV5oEoy2bLxL4FbOqeWBWXPTmfCMXMtUil59PcJYzqEAmY
2VO50ginz1yo2PJHaYnrwWqEJT1Nw9idk1H6YIgvo15kVw0CQzgRQoKnL30m2OvX7mnPUYxDXYqn
QfL67Cozf9U3hXO1tkLFQIZo6wlQC7gm434vi/rRapID/1eon7WAJQr2D2l4JTmqIZj8NR7+12He
b7e0/M2+OViRfXsLPrzwL7EyO8IN4+DMVhtfFJO7vssrFBGZWvpomjHrn1K7joLkXc1LQqW3z1L5
84cW5KXhIFmhtHu54YHfHKS+C91lqqM9FUphiB//XYZv5A4YCUlC6FQLEvjtYCXgbVs1jorgSFnc
soJ8SJyflDKJox9cjLk2Yv2bdpQtragcbMpUYBYBH3OtrT0BfVZyKKhp+29MemXYeCRRLOirWqtS
V52gSVYWwnRmzUBozLIrQUPStNWuJkzUm+4/NEGAtKYPhe4oyM1t/pUmdAVq+FAdg60v8cUX0hA5
y+3wx5hpR1pRlQUUejNE+mHRNkRGKlzJElFAOZhiHMH/9aX+zzfVcx36/ldyKIA/rD16LLftvQBA
BALfw3uhImyPGg/4kThdzM0Fz8fKcKq10pBg36QsrwkuFOndp5BbC4I6NEliZAhsuxBuM/GAR9S+
w4yGNeq4Nj7UIPGo/L8/r24JU8GilLj/csIx4cZDEg5MdGPWJDosBqAYI6vTkORhsSnEo2GrahG/
CJHUy+wCvQyDZDXul230PMfvHZjqMOQ6ymUzrkc3QwQ9FZ4LToPkPucMFLyvJoQ1YgSkgOgiGvDe
k/LaIkPmOnT8ebIR5bChJyt7nW7nXWEI9saAKtmB5ot0BgOmPql51iqwci49m4IwJnBRSnyGSDr0
9BpeXVBH5QpCk9f19WjzMU7XV4qooD1LTODrTwAyY0POQZsrrOV0Y0kwdqrPvXOkFrYYvytB9ENc
/80rI71Qutsurv+rPjgFKj0Mkd8b3HqvMZVks/w7e2iv4axP2llaFs87clbWfYj20ijt9gTgW5uv
RB0nAz+oPRmH1y4blPF0vc04kcMqYBRjWgBJLlMYEJFNBMv1/pzxfiBPVee67CbRgGzU3+d5W9Yt
kUl0WrouSl9TMaw0BSqlm6uQ76aVP2Bk1C8h1PThhL1p9uNTq6rDSeQajMHsK6DkxpWToFvG9W3T
epOHT4iDlLk6Ibbjape5ru9WWKpsbYmdjYHB2D3kEUsnxizsJFFgWMXgeVt+FfyVkEmCuip1Rz6s
FDJqe0hguxqoo66pAnx9rzYgVjBYMcxJ+olF4GiEzFC8J9AoOEUU3hZo2OYtIoy4qag2B/8Mfn2F
BobsfmWd+lhEeJgnoD/LROV4gEpBgMQzVIkh7jtiqGpL9pczIXxSaE9N6yKHgdYO3f08MyytSDXM
Jrw9JUbkLROxujcMUS6g7KiLeW9QO0W3NtRty820WfG1PkJMVAelWAj25fyKR8FWYYRbvY91dG5J
14wg1RJLybJEaVq6GHR20YySwN6oHmnoIcOgdI2sofMebMkDdEDthE+nKBUBrqNycmZgxHP4ENuI
dLaX/aoy7Zsincnu53zNQZLyZDuOZOCkZhNI0hM5FBEFtKc0a83rdEk9qrQbNuFoGtEWmP2MdmOZ
yHgX8A0dM4tih4Xv794tjdDRpciNIkjyf8RO8Z7YP+XT/VU3T6/gB/JNG/s1OzAaFyfuGp/ElPjl
ngUmPKyVRPgnEttQtVkJiSprChWpM4qnqEsCPfQXFbHMAL0hdzL/6z9Nr5iv9nxP7YjmiL0greqC
xsJLKBdA7DTusFkdrhzH7c01Xpm9pD6zExql+N6zUgOFOl15U7jcOMlkgtc9REqukWytyttOIfEf
q6QzRVsf8gb4Cindfdi5q9CfyFOZ7odopfYM4l1WFE2ZvgtwRAiCU00JiL/vk9y5tAKUjAx1lTDI
bkYX3QZRaOh6TtbugQs7xY1eirRwipCTFq8qA0oykEPYBJ4mXlzzZVx9TyZEdJVouEQ7lgSLF8kB
VVGyaY6iZcAs8/wqcaU1RYpUVM9rxISSi6WSGUPQDtCgduU37oZ2tEZ4t2SGX0flVs2MLnOFSHoC
d9PL6B8z+ynsxOkK9fuXbdqzl5pZOnmuXS6j0QZ85N9EhKWF/k7vjlwPW3M1J/SAKMvWOQClUCEp
Z2GBkOEjm7citdDrR88rsNlV6ZGQB8sxkXAcm9XL6yD/kyFwoEEPP2hXIZEf9tiZY0Okss2ERvM/
WGfgRboZnYbqsuUwJeTfYL4oFpSlQBUjYrXx1U5SQwqJ1kkNn6pad1mY0dzTjWWidH3A9hvuZBEC
iybXT4wWr820/dey8O9OOiupbZteTbaMq8a75FSmgcSLMu3IZGr9Qe6IXf0KE84jdeT+oHqWarY+
fPtVoAwU5/BZmxEL75dZWIkbh7oPWPKVkOqtvUsLQjX7dfsdmScgQPP+DONpteOSzQz0vzE3nSzz
mOyvx/Ee9zXesGvrOiquiMymi9P5hfGI1zlj/TbxD2bkxNMmWhYINMNzvEYnKjqXMlKCYEkgzfWM
m7QSbcSmhSQ4LQ1bcfCky0OQ6foTfewQGRT2AJDUWfKIUfgfzNPl2AinayrDEN4d4wBnpBJNRMqb
kdJnWVsUOGM91ajpD8Mi0if9WYBjqs4SdmZSALcLsDhJrgK1fYYmU09SHQWrV6C70mwtaXCFUwB1
Sk08YZj8QFV8vFUZeIz9c4MQ5eWZXGXcTpo6pVQsN9//6ePmVw96H+uDXwrMVJWwggEoQEWbXXNx
ZhAkrHPbFV2gRZ6EPC+8C0Qojjc5/KsP2z7bRZtYADmUUx84sOHBNzb3xO0ii2IPpkHr3R4nMqXU
1HXiRBuxUYkq3F1wuwKV4QniTi4Nat6dVCAXMweKhjcV5zrhvhQ+SMXV3CEi/Q6RaSIuyyn/tDRT
+luOUrU8hQwEq7651MwqQMSstLhaNemZj0/r3xAiU5I0MmOp3/zvkxJ5lOpAjGv4yigQmHW7jhaI
WpHiYR96intNKJpMzPTJB1/Fxuj1nf8m0IA+/lTR3XRVG6Vm+fjVrRmge+dpMa9/wnIZdmkzv6u7
1oHzcFISTlx91Xf+5eT0g5l0U988103NRcujuZJ3VPSV0CqSVaYycErwH+C7na9KS+fEFGPuLGX2
RuGHqxWjto0mDGafP+xIIBWwk2jpbBOzXXBQxyVA+FHbLGltm/6PQMuPVRN3NVY47JzjPjfwXgIx
V9AXm+2eSLU7THHNg9gFq5m2Jz3snjtWE159Zyc6SCbfHQ2e4DJy8AuL3cPE026aod5XFsPXv1nT
fTmdRa+r2ODNYoGZ3gUGiExs5r9LPgFs4nXEju3EmhJxTtD21XMpZdxt2UFx8yL04rm+nD0pR356
6b/LUaclHa0v6fABhP3OMim73p2uofEC9pkIrj84uxzvMf3RQQMWQx6Nmj79C/gKZRzE+WWBYQl2
yMGRu0bF+P8DZCUDgSbnZj8i/G13/cJhgGd6oWB8eaOl5Yj27OjVSczqdu7eGLidS0Qb92BBpDsT
/QseHtzTd7Zk+e5J81cr7eKGYgR++gn7FEhCsqh4nIkpmpqPVGMSpXdWr4LV76U3QdhIdkT94Hxe
vM7SzoXL28Pk9H4vbby5qHuGxucPaB6PGFWVxTjFFTVNwNCO+4pNKM9mUaGXQAoEETBfcLNIg/q7
AGHZMrF9lMZ+fVPEiDMl7WunfwKikXYZB9gGCyVFPukaLn0lU//wU8rQUrADdRRjS+UY5m5C4/TG
wvw9Xa5ycehAsqRikGtNok7zHPlpoEcvm7DcierqlJnMxzv7633pifwujdlYXchbK6Dh8KW0/4JW
Z+0rwmRgVflOZXbAeK7ODDZmV3PHOu9m/ux3xVM46v8073rj6GMUfss8L/mMwnI1UvjLMRJaassc
YDbWc3BpaYxITSWK0MILSAVBTTsAZWbdc0LJGq46RgDtrG2pvR77PUmDdkEGPZ/HYciczWmnlN01
zumHt6VeVEskjuE6ruMMpCQQ+v7zZlbuV4Ku0zQcbzxLupGp0Z+aghbBpPWqq5qQhSvZqZh4EWiE
uI76TdhVhNp6QF4WVbpUfSEB8Xko+WNaAUxrIHIYoZvo5+2gNy3EpK8RtVWhk7P7QQHBj3LIouiH
fAF5ImdrjvY6T48kM0YXi9K09gk4wZv9gQVUCBWFFAhiHaVel+CXAquy5DAI3BF+UOqbSx0fVuaC
yMhSRQRuvdTd00ws8Sa25PQkQv4wA+ezQMEGpInp+oyot+m4cDmJzPRdrrW34pzk3YyZ7pddtR5o
vDiDrWzYWsUj3OfKWYkR48cfNgwryy81cTG7+AWy9zNiwXdAU3/CfxFPHSRMwdggd7z08/jGVGe+
ho+3AdB+ITulz0T4846+UdnSwF3CBPAWGgwqvGsqBD3xKJKr4f1jAPu25UUH0Tlwb4pfB00JMxR8
6u++GTkogG4X7nLbdG3jv0PkxXa9ugqeJTB4P8QrA+KEQT5JiIWecWTSC85jXsbU8s7vw9+GRana
ymYxYXZshcLkChhk1OflfbbrjUX9pM2HMMXQE971rmo4PwsUdv0sUtCb6QdR7IO51uv3kVQm+Y8n
ruV6zEhyje5sKjjXtl+w2zaJPaSG91wiLVAXVCWIKB/aVjVc6Vx4H8ZdAcKA8nOPIUQDq3JFrdH/
dQSUS4gTCEXPi8tK0nnluO5rgVDEqLP877gOzGOnq/ytl+BwSgExOuh8ewhPhhv5srKCgF2NNSdo
Veyq1ujEryHqon+aRYronTWXTcpvKnuWz4YChQEyaOV/SPRe0/y9hDImlmHqKaVTvE4hFLn6xVmK
dAKdTEt1EIYkfU1LmDV5oh3wmCiHARHLpwCMxlpcVvKeGCSF/Kd7DE8pkdQdDe5KtYXjItGZmU/v
BzoR6YvSSL6d7SFEGYjBJAbPN8Qr9PITrjsb8Yx3CkMHtYxtF43P+OKeXN4+PhH66yhRYFRNyMvb
WiWTVkjKGKnqa/pwGbLpTM5Pgz2W1aoC4BkuOtPwkSzKpNauXeMra36i01hmyxib5SDQebFKm3oE
040fa6pM09qr7Aa705EAOo4/ZgM6Jl+pvC01biyfJDcCOBB+btqMfKHI0YSgC6IVSAbxArE0LIc+
Opa2b+fJgk8K8PQUvML7lRpfjLtQ1KXiSsaKYYcaYyKbWqQV/XcNPdFJWuflOpM4hD/OvedG4TzC
25zIvQwLbaeJPDVUJ+S1QJHEQVllLpUIwvq3RpeJZpyVZbSr0wK0KU68lFSjkeYxhOZr8hugPiQ1
MhUxo3xQ+euTO1mPXcw9axOrHSy65dSpOzzptWa6uvXn3niLFTRdHseiSY0cWfFhzEr21/6qGTc4
vXIkoejaz9NIZfLDKRYcKOGMLmCQQz69ru8OEdqQt97LiNlbOcukwTatmLlTcUlpKkNtWW0RjFL9
6FRsiIKi+A6b4BFFys+Ac2YSS5vE5UA7RLwaOu+P9aGp/AFFHMKuaqd3UtbbZ/67cYzwReAY3FlA
2EessUtK1E8HUYOrQH5sj/plpietscDf8VSy5qUKdujqtZZWydEnNGgqRI0GGhaECRp6ONWky1CA
asrycdAsuAFrvfmcrK6G8qIRHN0Z6qoR147Hcu5GvLAAMmGmjOBO23v+vxC7HYMMa43KhE6Xk2HG
YEAnjpdgUlN3DGbOcbBWLfqtgaKMovgabKdnGu0evdHPiofXCs7rsJh+HPGOry5Bm+9/vOPYNUyT
XpfM/pSHVVGg0qMk3r46HvAYMtMPb6OKvX+2z8+9eTKYbu+MQ6QcZdLpUiIwlhJm/58k0dGnRRY9
VGr6HDkIOKxKBih+JziMhcvCN9HTxU3ckqzO2uyVp3vO4SZHB81OKIB2X6HtwmJtYlpOFWUfRvlu
a8a+XRUqnq9SB2iAv2kfTgBnQlf3ENN9F7XTGUnE+h+PEdguPrVJ7z+nxzHulXBGPor3RvTEv0yz
5UW3gc3XVk9HGIONdXseefVUJLhVwCwvEcgmO879oULgbz/wJiTLenST3sjBgllRKf4RV77WQGvW
J+amUoKjO86XiLcAmXGo0vURANbDrQS4U3Ywz5dQ4VtKxBGyqOMm5ElDmg7YwEAWID3LrEy0+Vnk
ehFm8P+uH9ogQBuMPzhw3XB2MM6oUX8lyoPE/lQ3qGqw0SmmmXGb7/NkbOwqQE4tcN9aqhlQRXL0
8xtBAkZr8TttJy5oCRy1lwRjCGVn0R8Bz8LHWUjQq6WgMOnBmxKVOb1xkfzulAJO4N8Mn/CjkIrB
QQSpj6r0+Zr4PwA4fyAuku188sb1ZN3qcRlkos91pxnkeebVmOm2RsSv5JGPp8+DItr6byDn8vuJ
qRh5jvLyfRXxdueGX+wP1V6bmoxk0E2p1MRMn0ESa2/wgb5TKHLDoin0JC9OR6NGcgmwSuz57ilw
xfPYrqJjlBZIZtDRZ26dsbJRyjzVPFoNPMNsgqaHJnEMzVbGnlQtRLih/HxhdaIctjl2ovTy+vuz
DiPJMuHDceMEE1IsqiTE1EOrzmA4VlIN5NGQPUa5Mw1uWIWyWjEJFETr/5w7S8Pv2f39ExVWC2i9
iiJeLg0BBKaTisHUqZn2jENaQR/qfV9rAgxe+tOGh/2AR6vCZfmneiml7vDqgu+ITZzGFsHJOefF
78b+bk7akzFhiYhN/GrW1Ed5Hyb4LgWZwnH0oiRZHnh9V6YXQBJM6aJiEwf9BfqvgmehwIC0IC2c
XW0lPbfAfartPlgyRo+mFpnnCbSvdOXW/JEWs4hH2e22qd+PUIi8nIHp5+tpnk3XBH7qEatno0V1
MWHLwDZ4NbMR9I7ImPQ1q8pR8AnsgwusJYJIwHzMcMypHAYw1GNZNtYfeiUiFaqBOvN3ZdK12niU
6wOlJjMXrtW0mrezG0KgxnYVuOW1EKWdWkmAfQb/dxOOewhqsb2A8zjzJ3u/8s7PBsaY6NnPR/H1
6GsnpMvqh/Y+J0fFXXIuPbaRH8Oe1nDK1Mca6eHX48YYapLjbDoKBXG1NXsqjX+nJbXpYI299n9F
thxq70woFv6/kdwyUXRfiqb6eImLrbXPK7dWr2wO2W/OLWvczWCw8t9IUIZ/eVZ2RjCTazFMt6mt
jAa6FL4e08Zyle95Zwdip63ThMjdl8CmR53l87DQ8sadtvb4MZIXWK3wCqq0TiTe4TsEfKcGBl6B
nNnklIYf34P2JLeVNicHgezk87vre0rvgdl/ifNuyUx3Sp+N/hcwwwlK3nYgbCq75YJFzbezMPFv
mnSPZRRm8eA5niCTMs7Jobwu+CKUQFSMgmHMCFd9C/+pPQYNx1X1NP+wKpQ4utqxjq7kB8pZiYRJ
HEXOBzT6BeZzm/mIMswvhF6JzM9oSDvBlKpDo7g5xyCVPdS68GsVeVjeNt8hV+G6A09QJXe3G9o7
XfV5jnEgff6i+EDPTTlUwwzMR9Cx0+Mwf6zQw1oPGJD7RSKGsbim/exvH7vV5KcA3Ea7sykcqClj
RxA8OzJuWqx9uB7zmzHNs3ukWcRruSr52x3LCV6YW95N4UfWovQVFA6HZfgQmIyhNlhOTpNL/UCH
o5dMl+uy6b+NXpTeuTJX16iBgDHdl8dIk7JuBkgBEWzVW15TFmYZNnXo7/BcDgZPATmLQVMUxkgY
JM808dmZ0L034T+GMPPcW4xKFZON92l9/L/hyn7jdndiyVMyE5OZXsqqbVLrymcXPIAJj7iepnPh
v2RQE8JJ0T1XLzBNkxluhylOa3bLqONzV/ZFYJ83bvQi8Z2nM+H1QzqCD7PtobohkHVvws913RM4
EgJlO2eln8CM9W6vfv6xuFjtF0YqP+1GOy62dgJxMD1dpjGw3AZ2Znu4epM9LipI1i9UZW2uNzXK
T5Lmw7t+BuCxFZ914IeoRy+Gm18tkA/TV1UvW054POJuTjoUXDRxZINQdMugM+Nk8rZ+GO1mRepJ
+rItsJSKO++OAo06FfdEYG0evWF92HbaXBAFA8l8vQLBJIspW6GvA7Vr7ESNdHuBCeyp9t9EHvKY
oN1Ykfff/sux/ZvcNilcjapkDNwJvGupfxOGAPCEgBl0eQ/U2VtD3QctoSvo8vRCbyoinvql/5Zl
82WRDs5rhxkthC9bySLK0noZlnatskcqvrBbIk7hehBekNKOYIKulYaHvNFlY7CqIsobJ+hPnukI
OEmKJQcG3QI8Qo2EYubqn568441aKIf3GNs9N/cDJavVqX1H+fRXWXfMeOmiZLMZOEZ3h1sOXHcs
w7U6e0QNI/OqJGt/Oe4q5qPrDcWcdKu+7lOKdj9Ts1o5sjueB9KJIVEA9WlaByY8I3h0sVBU1pU5
r7d6ffufeledX2KviJfpyyjTwMfLwZ9aUp4/pjwb1h6VIoQ6DQkRrNFCJMX4qMvwELai5YvtboFm
EFK5fzdu8DEj0FOkI2UwsJNRbpbEE4rXU0PFeE6mEwDyrzFKzAuHvdel4iLpJXES1Z3CjpQSCjIo
AP9z1sdnW0opgWNO+1PVQOBxB9H8j0kkDM9d9YawoW0Qa4T2jXMPY9f6B0sf1dt+XwnVuwGGJGQm
8eiUyTZWKSBYyjAQrGKeQ35hV/0i2Kfda1URZUvcnO7CiCRRfi10iGGrxP1e2QZXvSAeeKf3ewH/
XHs5/JYyazmp09ekgpLfNBCODJtZ3iuG6qqifsPsqG/FuSxK8h+HtoOkgBSL4HCxyMq1eTQ2PiSS
GmMM4bcpumwhLPqPyyKZ//pmEV32Pi65P/xb9fHVPBqZNQdXcP8QBHMzTAVROWNMBsUJf86YFI9X
FD6PVKJ9KJi3mL5da/JsXD+xgPeolb9BVFPhFi7j/1XqMBYrj1ZymCsP/ZOYlPiv8V3NQYiqrZEu
i+dDNQYLaPVN50CF02dpfW+dDHYH2QamIMJMJhGJrvEAqW+nKMxXdLzoUKMrtRTLkydV47LrbISP
LBPY1nDFGLzAso8Rum7vqPuHM2Slb20gMY1onRPUcrO5WMM5CGuhlyl+TMWja1H55kE66vAqDqGz
wr0zs47cz3aFAICwgKlxWj7uesA+EmFBRn4Js/D7uhMbtj1hsuf+zZ87c1B0nxqan7kce4smOYjm
+0quoPVHhZnsRHGdaJs69yblstKyFdBT/hM2yCsBuoR2T9ya6xh18Ah9P0AeIIA2xUHMWQip7XuL
QQXpzBTugUgpu8OGQ9+dwBJSiPG7MkBur3RkgJCNHbweis8SjBB3pxWUTLQWb2DM89aXzSjPSkpI
ifypGtnLZ105MUmfXysCp3uKHPiQL6rRTYwx+sp/yabE7JabJMslK17mca6w7XzUSLOMupm8raGZ
9N7nicXMsybVjtY5lBv8WPZ9/MSR7oWmZ1kBKsVp65Voebx7TNCVCbQljvEkaIHr5jupj9ovDAnm
Dou31BQQQViwXwkPpQaszEkwKA+OedqAAa3Bv2ad/Q6vNS2TcymAde16xz66bBl8IFjnNZnRMR/K
qbwmxmlV1sHKz4vLh1MvUGmvlaqgeWmru8ehePBhQ5I21bn1+Z9zAhRdMV9gN2Z3+tIs1Jsgz5Ju
M5umXjHGRHnlRA40+iEgaso0CW15fF9rUCzIvea8W1zx6kcSasFqhPtUuXA5tjpZv7VTznswHCqB
bADy7WLXkNWmG9HLAbVFmA4DdFqy1bPgffyFFhcjUyXlz/koeVQRRLOo6xHSGH+qb+R002wNcQwC
PfZ445E9WKVU9GJhsEXydiJ+dPlRpFYN0I7WALsDeI4afQ4zcNsrjcJElHJ9jqG1wIrRxHw8d+Xu
q5+Bwv5C2qAkpDURU8IMKqHrr5i1g8vYLluH3guUZ3WSjkSsEMRG8tRZy6vKSJxPGFIVnjoJotJR
BIsyDL+IHInothZpCbunztPfwXu+wq/orZH4Y5Cjy0l8pePLowOL5tN/iHIM9O8C8tWW8fKSDBr1
RpTGx/jHt6E5pL7a9WqIYkwvgo2tjjWIPbTTODiTy6nQnS68gflLh+c65tHEqTt8sy2XMIssmIBp
s4+uY0qWY792UrOHRlw5hKjrlHN1ZWBsGq/ffNhdAee+v9A1e9XGRjy+tk5qj4XHz6c74ADzrH1o
VZp0qdaRk3k3gmUOMIpn9+u+7lljYJXJ64CIiuNsE/qxTz2NJyXHkNQI9gOX8swSc91aQEM8Uz4J
DBlCzxao6GqjO1AbWbvux/Lm6vm5bYM6F5ucW0+cXBLsPk1G7ZWnDS/t2HSKEe+Zz/OMmG1B2Y3l
WEMx00fRMAOIeChi+INbMhtYlEnU7mv1PcMG5WHNRpPEdIExLJEN4GbcIjNix8U9H+75fTdi8MT5
QpXzKLfx1fxvEH9n9DUcj2wANgMyS2dPV2pNUA4z7DB3A5H5j0HJww7pPIGcSjIZo7kdTSDaSILy
JvQ8EcGHNA4S+8j/C7cj+hQe4CuyDWFWqrwi/kzkQUSvbDu+XWZM18Y5ACn4SuGdziyxIJVhuirF
nHtk+NMU19Bhfu1RkyFEiyTc/DvCTw1B5w59BKendJVY+2g2mtBnW4NiOR5GpTIusMIaUMHDwoXQ
9vNewb4gwu6KS/loCDJI/dRHbBfOAbMaDJTzR54cbQBzj4DayDtQcR4KRgKzyQjrq5kad585R0Ls
dbZbTCJr1lGMqB2X7pAMq8/k0Lq7MffrZAVjXmOo2YyU0caiJ+nlSvAd6rsh+DGHTT0TbQ5yzBXU
aqXnSgwB30HRgrL33hDr70FGyuIDc9rdc/anJNYsP66MBapGgX++6sm0NExnbfOgwgOglAouPudG
sr4YjfwLfouHDEztzUc60x1Cyw5kllv8/t28RxKVWclUBnsoMLfyWPCJjUzK/kIj5ZYWWnjVhWvr
Nvih7fRQGrWVOb6DlNP0Cq6yaz/BndusK+LF6uGOWT48Lc2tl0Zwb+Q8pZF3/55iXRsTQfX7Gf2s
fbo7WL9e8IXZMJg7UFXUPshPnJ/z7w86DjuTzGTESVcPnTVtY3dHoZbWC5enH73G4ANfCxOuVmZO
sRYXP9L+Clsh7tZa8USmjmfYk0H/r6PaacLg+eKznUTnG1foLyLFuBg3XWEPMcsTtbK3RQcPzkme
cNvs1Zq85emcgC9+cqKv8dRnMUZfeeAyX9i8lft3MCnnhJKG3tJxe8zw3F7KOD+EDFRizwN7RELF
W8TwnQ2z6g3Bia57lR/XKyR+URVuLELX8Mpwn4YwV3MRGur0lQJH9jhp5DKj2SDWxAC49Vx4Ut8c
+UWnPrhlMTUmokRBcUpKjJtpoPztAvmZbZnM9kKUciAg9eGhWDL5CCPA6CRyLp7jPLFApk5GWyZK
aaTPys/vtbW63XKdUEmWPcxW1ofab4d3yF01B7nRoN8I1hDwHph+4mCrkLpH0XSAijPGXZ1g3QLj
kwSwiZdLhP6ot3BOR/fPUzTBoZXQqq3M5kpb23m0zMZvVEpiLOZJkHTbgcYwLvvpm0+7Lt3uMgxJ
95rtFZ1i5nmEEJbzYQg3BiYZ6h80nsAFtaYCKW9w/Trcvpun0wqqtYNrM6zcB8byMEqge4VvoKAh
GsARl3zmNP45Y18LKHRIAYafPSC8E5jw4SCGrTBDZ1FdJwloneh2td2sAIJ4dGdRY1Igw+DL4a+L
LizlRcOiffrtjX+U6TC4TujN0WXzNsOj4U7xfSlHIZyI8SOxBUlGqjvImMJi6YJNmHmSVYL+U6PM
DdEdfIfYH115qmMvARXk/0lybJQbHUvdU+eg08F5xX+kwPpvd7x0R8Yl8d2v4jGLpU9Y3EuH1rfh
CGcFFonCjxlkq4NABZ4YhUQMqrxTtPxqdb9zqdpcMAjuTdFWDHoQe6vRc3tytGGU0wWEumJZMX8g
phxF7JDjACZ8OeZm1C7v42PzOjOXRDqJPiEfqxIhj0FVJWirxmxgVHO9i7kDNj2oS/VGVfwnRY5z
nqW/z0POX4g03j1qpJd41E3+5CPh4iYGWpXUGCEPLdujggD+Nl7sME04Kf7SjyE8RgIIyEWM3LDM
+0i3AvSQ6x6mDUPcpZw3rniWaLcD582cixnn3/NwdC7NSNih7FsJWnYM7p9vdB/Egmrjx9Tpqz3M
6zKFqpwhKw/9oeGJmgdNhTVDKVhwS0bUpXHKfGIbSTJ/NK9aQ9VC2lsvec6qqd5ci0Ol9Nu3z9c0
bAsETlURobdXFa+be3VPxenMS4UZULyGV73fSEJNmmKpBmpil4XMF86UEwAHbQr5gxasfjtZvOZ7
SIQPPt8w81wUmFoGItwY9LCBA0WLxW24ES2NMBAEYHemKezt8wGVpOsS9S1FTmwVI0c0Q/oOgarQ
cXwuLn/Z0L8Ci1C+2JjDe9O8Zt+/6BlCD8CFMJt6tg8iVyAPhZG57ICJwrzf85Ciyn636PXzB5UQ
R7GzMr2FFrtE7PwqoIHvKM9vr9Sg4JtrUcC26Bg1XuiDhB9GOVaIxjMDtVih/Uffvoid2Gur2lOb
meCTmDlyf2xrHeNl6h9Y7OkMtt8ZRdk1QdXVYOiWCkI5qvAub983ZTUNSwE5XapJiQy8BvbjrYK6
znXD204XVJHuZGvOQV1b2Pcc78Li+V/x19t76FAnp7QTjImCn9wEspNfp3Ztz272/EgV6iM1bhx/
ivAkitYH9U+8HeZEzQoXAbIY+b6mK90AWIbZyd3ILj5hFfRifEUb4EsRYY7ueWVnTkJCjs0V1mWq
l+vxcsfyGxqZIIxxF7qGFudDz3Ws35+lYhG389Zbmzc+tOjwZpVQ3rRJA1nFzG5x0kPcqXcFyl5w
rDnf3Izrw9kZ8D3XCqVYwuQEU0oKO4Rn/vfwtmaOqK/m2CgHQ1bYLszRRprPn+RIM5Q2lWxJkI4o
7Q5d7gGn/XvZbq2PG+5Jqv+Xi7SAMZW3R5xovQ8G68pvbi2MqsIyQ8XpFHdr/0yw+Hah3DfAOCmd
gGw7KqF3FNTt8KdSeOp2lRdAb0AKHmX7tAlMF8LT5l44kUxdDZksnEknuaM5mlVoegbErOMKLPlJ
yjAknWwlB0jJZonFM4yApf1FVrZi+Ce/dCQS3rwOlORyXCvn9v+cO4LGzKVxWDVSIVtU5QgZ1M5b
iKbKIYg4dPHiwFhK2Ji79xYxdH1+5F6PrIjvXONru1QqOoihfdAViV1DhNqKPhPs03aQGY0Icofk
SjACsjZP/BHyuuvINjkirdXyXERB/oRUmaZQgESiYolVqiU3dlxwjcUa3IFIDtnH/kP6ul40VqyA
05JAY+pLt64+Z4cRfPUSULOkXhBsy+x+RhRLNZpd6ysBYJX3qU4XfRHe0LDPtUlAXagbkAhcDOIH
BFEKEEyXuo/mSqvbiyxtsTgDr4ggWknaJ4U8jAXAstQ7hKn1imHxCrxMZ0xsU+mEQpgOqU1cW4nQ
4PcUAH1gAEdATn6D6LiGdEJGwDbWuO1Tc83FJ9HtK8ZE5hAwIhQduQgpdIHtaKZpHP4v1OceFF1z
VTe2yjNJxjiYAQVloWITV2HOn2Rwl4qDiComSuLL1K2CgIWDuzYRsP9+NZq97iovlcWL6ZTFDIPw
8c5wptL4JtmptO0Z96BsMqXZAnMcjq2UxTn2f4OPErykmWdgRbkse8zk5gd6f2HDfB1WpxqqgkUF
ZxVsiUxXyQ3oHKzX3HfWyVHmYIp/bLsEU261ESn9MMjSZUd2KqLDpxBC/V0MujRKXrcuUO8g2OQP
U8Tz5FN3RTVgcPbkk1TaPmzfk9egDX/Vw2D1KdTxlV2vKhURUjkUD9kULxow8wW+6yBfGhe2w0/g
SXzvJ7nK3bWNc5HAzjyKMnWDHb9PlBY6rT3wIn5EFCDpVn2omQFZa+wo9PL9iwPL/WkKIvA7qGvY
BKuqoKbmpzvFtt5yjJG2fuOqYYsAdj86Kr/FW5MP20wgcEnIRbYSXzHJrkxXmOZmxacqWJFjRBgX
YWL+SSV0t8MvCXyIqYy6Vz+8XyjfUNHTWv0xZXpkrUJSF/yfma9ij/ev0DagYHKzBV9WECMXbxna
xaNEEmbcGkpzbh/K9+KmXaBfiRFGec6wjMlEJWOCG5C2DlTul/MmntxeuqiMUIdRMm9BkVedaxSs
Z+Kd3vVpTMhf6PoJWAiXlbaMWtJsFbOWdL1oMKbQCWWsCWPRuRnElXiNOY593GtEokzfXrw5qg0u
tepTuQc0Oj/ciPdByZhtWCtkrZFYhfsGRUIAVSCYHqn9yDEpO4uN3B8KcahaSQqtM9xIfahYdr7Z
4CwHY6Z488mmJ5R+K9jMxtZDwmMLoLERV4shg5bvGBjm0sZsXTn7Gph7Vf4yLv5aML0wlTP0p7J1
e2NgQjREIMg7hXiUJzW6bVm+k1E4hvc5JbOmcexub6Y06W7Wolqznb7n/e2jME1YTjmmK8AJmjeb
krwc6Q0sRXi0NqlMkpFecRSEYJ34TDdjs4Q9wI59ObtSiK19e6zax3rclNaKu/KvfpOfN+7P6Ug/
MzSUvCUn5q1tplL77Ut4lwQkBXaYhOTmDTJQn41d5knXWyEzs4l943rlXmwtmbvyHiLGmbO+OVCe
T4aahfNGgmeqH7knjApI2Qb00KNLT6cz/S12Tuw4y4+5nv1cGOJuR8pD9mQCsmcihrf9V1r2mcp6
OzGSN0P9RxuDTCplVptJ00lRRSCwnSU9FENoGQWQkxKTmKCV6c/+jCJ+TCiB+dopR3ZUbP1E2Hvq
6oIzhwzA8eRLYf7iC7ufP4do1xLvUDckU+kKTRWOtZ+mmmZjTaWXiExJwzx7yJkbYRU/6dofsosX
QliDIWKr1wLmAt56Ea0FZBa6UlaYrrAABod5z/iiFyWS0iLYsYscgidobuaY2fiw08VzotPkaOhh
4Pn4bz1dwNRKR9ZGJSEhPiisdRpsPuzvkhHum8YnQbC4IHuP7p8EkzS0tX/oXJ/yeLdF6rhTKyeu
JdmmXMjHP6E5dyJcvgu6qgnFXXRC3dOv0moikac0DGukD1RRiDf6q+UKGeBdpZQc1de7iFGDzrCg
5/yLtaJJlyQZA0rj6mymEZy7+/HmkuTCchoQckYJheMjKpd3EvP7xGWMcsBbtYzwXKeoU6KgsiLw
IkzqLgwqJbgqxV83dek4/bY9sgKS2S+9c9hjGNQW8gN5mX42PPu8D2fXxSMU+X10TqdMV3jxikJa
96TuZWW0d2kHPxS4FidBUlTL52XrVqQhnNFpvltmxPM2546E67soyGH+n3EoHzG7ouWll8phT8k/
4F+Mg85JCDuri+hC6pZ6SkHh9meVOiUJ2XCZ5WPC1k3t76TAndb2PBgpDQpmzh2enw+9FBg4vsvM
iCg0CBixV3lIad6ru1JZa7KNJfeNDuxSZ3eDUtMY8VcaU48kBmAEobZn1BneXnS6HKUIHWqshHHt
/udvPAvJwiVQKQakPDhSP9yS4z6OlYpFp5km8guMQltW7cDfnlqCZCTn31kPFYa0nzCpLXxylkvl
NyZBxp1ZEYNMHl0y4+PodTpBGOoOwvMOvyUErYdaqZ4r9IlOuXW70mk3HZ3Q5uI+nnM0fvq9ToiN
1lP0uwpqgUjCs3wsG93UkcsbdbmDA/l90Luiq0Bh7VFE8jkVVxcK8rfzrrNrMFyOFka5A4OfjpnP
AqtIJPfCuJZYWhCMIx69RSUrb6QnjBS+jXzUSRDhdHW8RnppF7Ma8h3XWBTtK4pS9S+d3DK/qHx2
6jQ/HrecRgIv0MJW5fD8bZRPap0r1R7za5po+3BB9gw4ajm0UjDyFDq3c14gIMj4Sh/Mbmtwau30
RYqaYjyhwtWg/xgbD6GnQy0WoeSRiUN48ltVzs/QFwhTnlH+HCh6nDi/wwbNLr/UVzr8Z840nArY
BhApfaRwzMVtv0g3QE/e7YhHyhtEW/O4pAYGNXs0eKsa0t1tmWqTQ8qujH8FLXEtaYcgqmmuKOoW
MV1RSJVaV8XHvNKxhJyTL2hxiquwruNMA70tLygQOk+DzZjK1+RtmBM3KW/GIgO+rNJzAqEIQ0Q7
5urg5RSJ3/tyNyFWSmyUCeA+dfIMHG6j1KH70RnZqkSqv8rEmmILolYnu4Jr+0dt0HD3oF4ynC4e
YqW5OCgvaoyilCRTNUuS98LsshyhmuCD32V8DeVCeNtJxvwcerBwQ40SjfX1qMLsYOBa6IxvDQmf
SdUiMmto4uX4LWAlHE/z6Sped/685t9MMUl6ZiNb2pHCykFaS2o+cMTrWwDB2rXqn+momxKKWD2G
GVD8Qt68z1Oce7ZvYTHFCBj7/bBuXVcMGtONwTDzNGNSGnW9u1aYDv01LdndFBNG8EKUoKLe1qx/
fWMbjR1/HZJ8iwP47shEWoXk5mhyEQQ5b8w2NN/dDSAtav9+UUMFqcJl9PJnVXDI6GqsFKm/4DgP
KzzVFTqGFgm28XuN0fQHbQ6s+/ni0Mt9zZYWbigLepRJrxE/AwE5fKb4W/yG2hkrN0oFhEwbE1Qs
b5CyN6qqixxA0+V5Vg0U9QuugQv3ppL21hnzxxo5wkyyC2AsUXdZ+6IYsdcuU3s+KxxplFP3dvAA
sLNwd0c/uI/MY06gnwRyvK3f5WB4eRopFaPz0Ec0W3aK425Xziayzf4IQTgAEd5dk50PWhC7gDMC
7z2TxzltW13oKLZ+6zhZr3SwhpIKzdFl4HEOXiq3t3TsCpILExPkUxdSEv9IASj7D1SyHqFDBH0J
SpkWp4qN7LZV56L7sQDj72v+phzY6SeCYPjIObHHtQTd4VlPaGXzJu9euQ3PNz4W0DR53/x2JLiM
wN2kK/UfAxmuhUrOOiFIkR8XYNqQbknvcfsRJ3qKY2I2QiKoRuqMddWTOviVxhlWkmbf8jRHsSj7
yp1kpkPksk+sF0EavihCjdy2uSz869k8wtY2CrSo4Mo2/KztanJ+oyHcqcJtz16JqzcWmg261nzi
dt8y+ZspdRRvD5dj3ioWbi6bREtHoheyifDimMvEg1sMnxFUJP57V1unELhVlTEYkaoEH8/gnIvT
3B9qGRA6VoWTaRgJcUj/Ocq/evAGQTWouhBtGhmVa9SCj4HstprN1ta6c/pM2kAjhwV7xQ8zlcAO
JHDaWHiurw/BtqbatGwh/Ln5QrzNOcM+8i80CtyCqivQjeJshSRJbenVyTfFEoTq/FWSGMPNASeE
jZSwLf74JUyfQLxGdvXyE8vefFYv/WcCMcKwwzfhb3JHL8y1mbD+piUFJahWJpnHFWisrDtbsbss
rrPXGQ/TbdaLg/PxaPoZlDGPaoG/kdUokblsZAStjXmZkHoTKoyDYPp4ErjEGMqvHElW6lhrId0O
wzCo7Ov2fDQQsh8DAX8RlbKrpYDiXt90C5jTYDCamom/f6cX252pL7sAw+YLlI9TPEiSN/UEaVIS
8n0KYRu9jLokeQfcZb7+2kf6va6FGlRZ+dR0uAf3wzB5c3aZM+1UoiqABGncZQbjSPMvEXz18P3S
aIcEP8IhFHVo3AbuShb3ehV4nfCxx/Ae7yyoll6YnSAsJ9JqCM4Ni43DIteXPzplyRdNFYaDK2rV
UkH2nfkPPdfD+wwNT/svR2Pj7j2B9BpgusYYI8S9PQsg/iVCBixArtLz52my9leJziKz1ddfqT3V
rWdsVTIdGgoTBwURdaDwdeToLaaOWjFwKR+xlUl1jfvLC5QkggjFf2cNYGvpGvpNI3BIPalki4i9
NUAcH9hDLa6TPLvwLbM745ooPFfedRUPQ4kRxvbuIFySyk5dMq0L4ASGxHpHNKSimnoAaTRLu0qr
wefEb/WtAgCZnKjCpQL1EOsr5XZUTddK5bJ+WTc3tRYH7z14tQYASFrVQL64Sc4xF7fIAvhxvc2n
gUiDfiTs0V/GzxEzpmwJPmE2Nrnjkur4jouUdb9zeYJPmkNyzT5T5CULEqcjvy7KNlJzj/WH4e3Y
G8CPsoKDapAU7uNk7kWS3LooKsIsSG6IhUK8412nOWthclqGKOvCGPjLp69n/bGlmn6eiqBmzkEv
O1fZaihnFcX0l3SSmpYsdaraPGiDzwdkOKxKzeakjPh34rcZSvphOwfh79ZCrZRZ9mq0rygBi0px
xvebgwPLJPc/BejbhP7NRB52B/pCJv5FbAQa5Uwzsc+PqSmzFkEjsFU0nFWJNvwYff3sJfUpH8Vc
NtefwbA8xJBttQICZAOQt1yf7R3YRPYn9vCV6u1x9Ym9KD/CCMU4LgTkoNuKEzL8TxWAwr5Uck7S
py34dGAfUKyWHVTso9252Mpm6VXTpfEKeXkzGKPuXRjhSbx8w3uIAjj5qe8SafgCqZxR9xSqEGuY
rcu4Atw8byFdUbzPeZoes3u6C8Fhpr1wbnbWfsoQamshULXM4G0ZGvBXBjqJoAX+2ww9wQtUHJRB
MVoP0Hwn3xIedCx3mJH1en7V6hFoi+S2d6IETpP6+4LzA8tTk4FHHh/LHrqJi9KPq9iDZWilp0R3
J6gFWvYDXi4amEmOBEgd63QseMQgqoZPo7/P1GdvFLGCGlHjHwI3fCFZv0wtovcsiW4qaDvMQYGH
oI3WqsZYZUx2WAWeyD3ipPqGjF+Tu/wVcknKk75WIdrOTuiBiem4T6/qqVv0vaxmBIE/ZDxC/rwL
Xxqee415enG0uKR06lJ+GWYTXfRki+f84wvqmq8qrKrjlzj3Wqbb44d/CgPJxG0J3yy95afeqa0m
Lh2gLgu7oFfzUCqZrda7ceVQUi0l8ZxKXoBw5uIpVIg5KfOqZyTi62NWao9SUXBr7iZy03CvV2Eq
rzhITueJ/5fs03m5QXxF2epFefWlLmtkRBx0lJ9RlFHZceP9wkZHenzaCAfFDQd6k7XiKJ1N3uaU
aV+eP3TSlPLnuR6vtLmOa/9VPBNfGRevOTQ8rgj5xUFztsErnpd4MRawX3c7EoGdD65EZXKjKQ2b
a/5O9sy4RkCyr2XYu01LIasNMHP2YrTQoUyQhlL02GhNOs/KIr4RQ28pLa2g/zdtRGpt6MsfNR8d
Jsspof9rNExGKS3aAdIiXY0oQHGoI7jzRy449TI6+Qbg3qINBnK60+pYPGctKYSYsgsapXbmg7Fw
M0MS9sijHs2HYsh6Nv63cOwWvHUSiwGuqA/s4UsO7na3XFDLALiZ78ZskJhGVRVysFJsmpofGsuU
oQ66aEvtWXxKxEyfoUNPBr2hadaoXnJokdlLlvqitTG56QYnv/khhKOx+NXbo5+aDyzimkbqDfLM
mqqsXoDO1liNwXkRPQZ4bW0NxaTDvMn90wpsnUbnDAb69IBa4BvG6siY0oRZdWsHaPZCIUSYQG7C
myk839bMTCJUb1K6gIcLvas3TKHhotS7eRHQgnwWh98ExOsyXFLxV6Uqr67LctoXONSOgHIt6ksD
m8n06da4vU1qNMalMsXLM5ngGmYlMi9eLLIvwj32XOOpmhBh45knk1HMv0tdx17tMrV7N3ZyTfea
S1Y9n7Dir06rDpGJl8YPeRpSelv94AUhbcbNjPpFp0soLC+AJ1xfK3bB5zxPhIQG2t3zcFyfo1dX
UfV1t/2r/r6DoiVjhCArECUOsvpdvoaogb/zOb9xAVWVcavelh0dUrEjtERuruHekSI7tHjOTD8h
8c0v6WSuEwsjBAOSNu38LpC2NyJ95Qa6jdxI+EjeVezfxfSprmslfhFgitEw1aEKZ+GnujJgTkYH
3UXVskVVcBWMO6CImB+YcdrSK+C1sm1R+nvznhKOIzxTsEtpAaQtPjL6KSfVksaJU9fRPPtfVC4T
d1AzXnnlp7sJ2Mv7+aN61E62SB3w2xG48fZb36UDkeNEDImDvMEp7HSN7IILdY8vOnpMcSnlSXSw
iTUaIqQMdfWLa+TYiTh9/lr0W+I09mSDW+5IEsDW27U5EY9udZI27xasHqbi+PRljvyBm7jX7z74
1GFdIoHqiekOTu0QNyXMjpwX8E8or3WVTylZGz3uamLyujBlaKe8drStPajFDeb+QYJE8w/ZQ6mg
4QcoRtzU3TUkWy6kpE+ualqYXkOx7oDM1Y6UYhqBN+Wotukedhqks+ELaX1dKpBxqL9tUwcd9ovk
yd2gcqq2z0AHGsZa0IarctFr1OGQR8PGc1shwauax6PmJNE6ELav0dwrjR8V7iwCcsu3bq88w+kz
CJojoZjzJTcpgH4FoGvDPlGtBXtrQghVad1Q01CGUJAutTiKM4L5RjIsFeTR8/6IhlNGHy034r2w
2xhtKp7yfoljiUThP+c/EF5EqrXlHihti5/k8/sXOSNh9xwHmnE/GT1MrPaGpe2WqW+H5xXjXlak
pZT0u/8thbiAFaxMOfayqXTXOqu0dKzjPKQFVPzgXHy1FnqArqAKVWhp1uT4/9HLiqeItQ7EN0q7
Gw1cPcG25BHEUNWoqJ9Ya3S3I3nJyeZdWtvYHXFijcVbjlkTSDkfXGxMqOKB3qVm4mKpy7ECGmyS
j9jDfqwzuwcH1SdS7MdqR3s8BAysDUir/UgVVyqB416a9fm6mD93rrpSUmnYfkzJhSzg35ynvkPY
01zXxGufH2clJjVxoVxbO82Vz32CEdGA8Lfp8Ml8CrQLH+I5tLCd5Vl7xTlp0vkNUkXBNA4J7t+t
DbciYXJqoE5FY89HEkxgWqi4Wt9QjGDDktBMVAQ1gTg4EScFCTUG7uqMdDkCqZSmRQKthJHlTJ3M
UItSYjZ1dd0ZJox+8O+1VoplityruguMUPyyYfcECFfn/NYZFAsYly+wXT4TixM6yqlNTNDaLPjm
As4zhqcSiG1zAzdoYp2/rLk7DL7+eLQRRecqWuNVstS8C3FgEEBAw9i+xJ4xbPSWHjtW23oz+FH/
vewsI5WiZ7J6VMwlsDfXOs4prMB8uRei0f5Dx1PZmOXPcRJvwOpWZSzhjU3hwzfG99xQyfctyTkO
LvVrcS1jrTni4L3RBf+5Nb/E2uY4k1JTRYRoBLopezTseVFseHo9mG3rrOOOQCHXMmcTm6mjz+9e
PUU755mjq5QW6KYWBA94N92kp8PBhmrriP5Au0Vp41BfExdUL+cyNNUHkD7DC3uTzSzj3vo7jj4i
6QcRaHz0IQjVQPmvaPDKYDpV5x+kV5eMlL9bkr7t39+Y0kcx0ALRy6IyJSsyrszZfFGICpb2+Y2r
+cl0BH8H+bZxMo0UCIigiXzOUrzmeVAxIoalfSETw1P2Oj7tK+fx5/pFZiLpy4m2AibDtc8K8Cu3
kQnO5GAVklcvcbvGthfUlqTJCK4doTyYaMR6zOiIBuk2zJQZM7EiLq7gOQi1AN3oebJl14jx5hf7
nbb6g/4MV87tbbOiTkzJ3emnw00txSBoRxmZZ/j2jr3xNXDuwEyeG71blm9cOhydyEufQF/ekAoj
4aeLMAghB0s7O65tEFfLz0QXqonTwiORZFF6rSckpJUIZKWqDDeqsOD8MgaeMZIdeFbKpfMrEKwa
tUmEhNbYVzzrflDHiRtodm1bP1F9RTH9kZv2fiPB99Y0QzdywuCfCqMEOh8jySUr0oGG5Owg6INz
1LLINV5z8o9hE1Y5XSfvQAgsm0/gez2o+BPDnSs6Q3GtpvjFEB3likgtGk6gPH1dXjVNhE9+XZ65
622/D3xhAV8MGOUYmtHEXf03bkfGEQnw4KXb0b1ff29s6hBqz9Xp7fC/CW+SRWQ0VRxq6jxgMN+v
kCMbqIFRyU09T3avD/5cTnLoOmouRVAhiiPU2IAt0bN5DlY3QFDZcLZWl75MuyEBUqkCERdeqj5E
scsb4fqb4d3+Oc0O2qoFFmmZO6+Q0PlSxEEpoCkGMEj4Xt0pn7v0EJVDsQi5OTD01cGNkS7Lm6Mr
W86cfNfBJtZ+xPftNnhbTLYf72lDWii+bmB3P1eVb91lFftgGjKAqaurtcgZUcvqUkytK7id0Tcm
jPmXbh+I+qo0aW1Ij0bQCc4WDftz3tDd1x8OcAc+TvK0TM/35dtcT8Ju+aqBtkexRozoMIsbuiA3
oi4HTfoW4Sece1vYnxRVQTibQ5P8rWommTGeI5gnrfKn3s02hYHaimBg0BUhY2QtVOkLwsERZNp8
kOpqISro6bBia36+91hjvIw6/nO9eQDoDBoO5rNdKIi+orBDnrbFLNjqzS6hOw81cWCJ8SxlquP3
nfXkcFYCKGLPHB/VV122EMmIaYZcoBx1tHKjYVOF0rpF5wO3vwfaSlChWZq5bQ6ZdelwSD30Sjlf
37Ib8r/fa10d3rJWlj2cZlcCSdUGpLVjjZ2OjGm23shGaeTHAY2LtH/z7eoMZmk+6rv8ifjg6mLX
sej0OdEvf1vN1ILOr2MRdcXYFoNruMLZhScvGrGPEtuu9/vsJs3M2nW6LCTSGY/Uqfd2pL8PH81c
Vu3yuxRjh7zSCdNGz2lvCMIzAIP9SmPbzd8NiidxM3AO3eG0rjloOQOnwm1i6E6eAzkFSpNmHpwV
xxq6CNxdi5ERy2TxKi3UtV28VTJi6+cQrnElXCtXU1znMQqkKRHD9c5M/nezFY9XUfU0VVgKfTX2
BIMzOW3VfNSx3Te0XUxPh3NSO1rjCaT6kqr3+M19lSy2irhrhQVXKcvqZ4W2v0l5RCQHWPs42VEx
pc3qwft7nt6AWF5vDSb8Cu5mLvhUG0C3CKzZOZp6PiAlGyUXrmc5smPGBPDWcwPNYgqEKVZ9Pe0Z
c9hYpG0QOVZkvBmrIaM1kiExK4oO0gZmcauYmzfM7cy0z9YGZIgczRZlAf5r6sxjoRxSQyV4ONW2
VjrZaHPi83EVE9QSpPtHDOUDW5/HokVXIqX2YiWovRBoPuXcI5ZjF9r+6ZnXEyxROPUf3ntdb20R
E90D2CCCetCJqPsZ17b4Hl9XLCSRQlI6cJLM5NK5DpQ7bF2gFmaNgQpW9bNtTpHRm2MiulhK8//f
cv98xg7+R4YK4Gi7aZUWEAjyScrL4Lvobx5fIrkTF0wX+CK5C1qTXppngiYjLEC8Y2AUfvOFKcgE
MPHgD1kFgguc1lvcuZs5djO9wWnkilo7ucxr+0jhG+0io93MA5rlcOl3djUkengrIsh9QdwfPEh1
wv0Air9SrMFN6ArKxr9jKGOQyGA02bm0cdE1s5NAqfHelyeVbj3jmZoYJGRISjRk0ObkLUJRoyFy
sL+SsuVIfhGXse0iaZRdr2OMUmoroQlCSxumxoD7FnkYHE2QledBLD5GkDAv1Hcyd1Enu58XUcCF
/rCLHLcBMBF0J0dR3/cGoHa8q6CZHE2fTTd3W8iZy2jxnJq1xYr7IaJ0/XmAIIoUfKaPQ9i6Z+PS
qWKcJviLITZPMt9kFXJusgKQPA21jfsBECOgGESx10jz6lZ8lRTime5l49be78OcSI7sy10U+DV6
koBfeEExZOwpaerQwYyppaxEy4K7JrKdQDo/u7HudXTrgIOUeeUUXi5zASRQnmlI4GM9cyOdWWXd
68XURRJyke4XRR0y/tUcwram0ziPoh1xT0t1xiifmzAvZBVfed6jzIO0GhzIDN7C2GD65TKFuVAp
Z6G1wjbTrb8dwzUamNKmczIGl8C0wDIXw4tgcjEWoTeJcWwszPJiMNrscx1Yy9+/LgP6oK7t6lxG
XKsiMxVFxTCZBHUkSqeXbla41hd+mylWlXyVgTlpIqjkWCqMGdarkqrh4laJkDjvWB6zjiPwyKYJ
FVBpsvQtAmWuCN7rt7Byur30QItA8bAoJkF1MekNBmHdfaigcjFaFQEJ01SMACOOJD4U2N46Mj9I
wXg/LLOpB+x3iQG2LwfmodSabpjtxt0HQBgORBtQ9yVh+Ev4ptonnJfKaV5CqYtDTAcbcwJ7Pw2Z
S9soquKj776igRnU70KZA0YDX32rCg7ZB5So/WrN/68NEf5XglX6nZkE5H87PtXGgktc0kQkf92A
Od1WCE9cPoahVQ7+WvPCyXhHhHSxiV/h2XJAVy05xyP0tOy4Pt2RcYa7vpXEMTNCoAV+LBrEStiN
UcK/4U+XMzKIb+QCOUazHBPj2Nr/LX6NzbpFya2YnmaQKmmgTRKxA+5W6Tt37FByHuq2WBCXsYBs
wgH2+d133higg4bywFnYk0E9t65EIPJ88byWd0+DPWZOxreppmh25MTuWwvepQsYB8D6/ZGjKkcp
93Cvrb8+G1g+srhnxf3VXMsiK3FHjU0bwHcMMPIPFJ2cb3/KQPgOPO/Tv7BaMQIMAP5uNsuvxKUm
qinLbcZKP7mde2Gta0GtG3SQ19tC+sPstWKeEsS4iMa3PsDlBheN44BeliMx0v/n+jmDFtADBl1G
UuChUJOxrFpAbi2MSr7AG/SlQq3+ImcYEyN8bxBlzlWrSNO7HdK63NVgOM0lEi+ZjDZfHQdP3Kqr
pFZgq2bVB0jBTVVvTyMFdBoH5ppLvPKd3Yo3PWaG41H9IIgujK8IrjJQowuTGSEDY41tClgoshxQ
wCKc3BY71EcsGpiJFg0PFmxs2E0QfQBxpjamWxhZ7XIOIEfLmCbDA+XkbJ+eGo01cOxVl3oO2QPl
CLDAAAxvL22/TeVbB7AspEZkIod1Sf2kNEy94oJQHVfVxK7ypsXjxY7pc7gq27d7jY8Vr34YSZVG
ERwO8Do/uO0IZkeCqP7j50N+yE+5QXE7DwREpvaZ2XATkq66tIPuHUytwfUyKab/WIWBn/VmrpBM
ebC5EdSsF+ZMkVvKtgRh3WerCtdyWc8HMakeqVP09mC/CObEKg4E6BKHiuE0N81OlQP+ko9y7zKB
T98kiPojbSHfNkHblRm5Zh7yskRi5QXMMXR7hQK3C5tqNBJyYGwungynIQkaWdAcOYFEpREpw0M6
raVCh6SAo/v1zaV8BUfF9HhSXApHfUWwFwdXun9aRSsaF3DkTTKllt9Yj+URU13DKK+fPTV8qXq2
+W2dL0K1EPAh4V7Y3QiGpvVO4CNpqNJPHJP8fP1VvL2A6Fc7ybJZn1hMEQeTiQ8Ck9omahpx89lj
w4tsmaw44Zp0cRSc0rESP8gu5sMFWrMGjTDkcvWwYMVSgEmxa1NQlzuWmtvlHFmW+hDU1kvk+See
9rccpCaMzOR66qHlSRoISmKrs7Y9MqzZ6wKV8pMlt4KRJl2wvR4g+idpgWYQaZeXLPEqJ/CjkBJU
KnfCJprZ/EWwq2hoh8auP0Ju7SEIoEB40/+1lB2mfb2MKbjdYvwx/+WbradJpkmmMPBS5GubsrGh
LXpDo6zv2qAb3Dw138DwstfgkfpVGJwhhfKLMrsSWQJNIjFsdvcFNI3FIKWZFypbF1mpGrGqXzB7
gEohLrqhYZ/xgasHRBJW+3mDUm71vYdLgd5Ki//kNrJNQOrrNR6uZgap8moYkL0K2pS7+fYigoaY
giKqtirtBCSXL63YTDla26PcuMXDF/hIbpk0Dd6h8NoqQLI5/EWiEV1FYwM9eAinLBTBKnJuc+jj
ysQvmLwPcVgBuoEE6tyyv5+y2B76Z002usEtoqkgmJ8vP/zzatNgtkROF9EbdleeXXEgiIQOOVD9
ju/iNoR/892AUo8cV0dnMUzcx6+LgevJX6iMsp8gi2T4cE8HYyUxjkwFiLZrrphjFgRKj64PJXL7
eV40VhG0Qs+1/CXToAdsq4EIE/xLVnzYAJn6rqqCkZwKr6iaU1rYD3XpwiudDCW7N2UBOfWS/rx+
PriKLd6eJPidGMy5PB43UgOgf8lqmlbF4havqfzHqPiT8+VA76nwlNmXLyVkoUVxpn4QEZbWuPva
k00/ys3lfFs49sNwbvT86p70hewrv1Ny8UwaXjaOWiJjbwPKreDov2k85kTjWOx8+/np6jGfJmH3
g+JWWzdjHKBqaja3QxStjllBMYNkITR24xGlrgOOlujL0C0JVUoaoZA6CwEUbNjY+0gxoRLBYxYr
58mhou07L7s1y9OqWab0hjpZx9c2MbDH4n4Io+kBHeshjZi0+WoZHcEa2Dc+wKjSOwo2noVaHuTq
Xwbm1HK3XhNjn7uWB0j27VjfCgnawfLWRtpTQ5FNMUN5AQwvwhtxdzKBrBYHeCEhx2oZiFj/opjx
98Fy6yKEJWEHi1IV3Mosy91dIH9nybBqB3qf67H6S672bWFahKbmEBCTIOtquxBV2d6p1PTAFJw9
UVueWBUEOMQ865JcuP5yT+fAfqbLSSY5pGaDPM/9wrh9RIuuWEhE4P5+mjKR/iy6+20g9REISegT
00vlCMblmkJa7AHEHsTSQc7O+MIYf6QaIL6n6hkjLiqhe02NYmXnYxTfmrVIjN+JVNoUbcDPjdzp
8IEvcsRP2KmfdylccCgzeUJkMq/tgmNoUzddfMwKfdVLsYVu2RVFP9xOUtgDPQ/4dFd9dlmptaXk
SiGGjc4P9jods4B0RCljVOKZYVNybGLNRnjWdE/RFYZxCJ8BFwpnzojRjclfxT5D95j8lXaOtX3Y
6C398jz7C7sAKPVGlUywVVwQ2eCO+nwToApNNsCceGYf7mBN+5tJqQC9QNV7deIHRmcSwZXIawsO
cz0bhIfA+HDUqEzUXxZxlW0zhlxxP0ZugNJ+TC+OshWRKUVEwSOEqeUL6uhrUz8Iv2gmSffqwNKb
554jm7gorsGzVTW4xyrJn8auE27qtYfEXCjVDl2ykKfMfejnEhjflJEei4UEfCoRqZqw66dqhPU9
2uU1k4zxVOcYsVTxKTZ0Zexgj+CmLSwvKkOhACsuNN7qhWow/6imqgD088AF7nU1FLTWgBOFT5g/
GG2C4h3JSqDVkymtfESdrmt9LXgKc1/HogsYtGQnB9rLG4ybc5fPkL6eAM5uK98RyP3sf77GvUX+
z2U4dOD1Q/hnkybcGVqHOpeWE6ysGTh6OQi7+iyXGx+ICwPDAxYU0PWf+vTJQwTe3AsxDom47wjG
rgOoBFYrFePHysknPokWQ16J4PMuL4GTx8FotsdsXcUyQL+uOBpPW7bq30gavpXjuXNN2ZIpI8Au
wiFuApXgDrRoAR20zq3qFJz8WiKuijcsF87FMNCRvATZACfKqsmw2axT27yv2PZt/NbUEOx63r8H
aLvSMoWaIuxt8tfu8yC2Z5sXMm3TUMVb9miOEfYhvdamSt33hLh35g1tLjsFHxGUlt6PWsGlZzrp
LmA3tD7gL/tt5GEOGTwwV4A7GR1O3ElCpspKM83oHRMXGxkxx4Z0PRnG+U6hpOOdYcJOQgzwL6FW
iMScXSDiM9c9kQbObErYa4Fsdhv6277oZeCPTrhgJ7RpzxVn1NaJSyZRXkKMCiLbDU5fvcweMKQ4
kpeM6oidlD4v2uf45yxVYUoF8/stuz7DrWeXnRDpNv2Zz+vnYR7hjH/YoQaXpdiMUbZ/z7reKkHV
TrR3dFLLjI13Guqat9mvfkFi/yRdbQtpDU0VwoA7dCD+i6ounvPT+2UwFsopVqzaWhad1ZiI9HHH
5EFUW4m1Px07uu4l7Xq7DAamiEpiIt/5/Fl3JaEvoHWZrww81lK4NTsxwfa4KOYAvPwNjUKQC+Wx
vf59RigNHQcGBQRGZsD7WNblgk4bZKwjBNWN0RpSFBAgu6Bm++0JTlK6hLEAES6orOrUPSggbqsr
ByJi2bG/Z9QAR0XLoAr9P6CJr89883OzILKKZK0PFob7JrntUExdLmA11t6Al0Q4FXZky+G2gsZ2
zlgUFUSZS6NtHfUgRfrzHSXgjFKOOd7o2ykR+6osfEqgI38qiHYi2vxQJt7xceupqJ6QRmnd82Uw
Lw3/yVSiPznm2HDVjW7BnV9CXaqCq4O66x6irj/MqHanlSeMsTx+eE+yDgb42O6pN20f9JvELsVn
870qum2U3+U7EA+HtjZbWI6avkQvnY+Ynf7ZG011HkhkMGNNqypeMLm21KOwPHkt+FNNweP5Zllb
GvBWTnyqRq1xzNIEkfJgomegdR2KXnwJY2JiP7lof0lZzqrexEkCmQNzQXpKCAsTZkbU9rYbwsBH
l21H/eEFQKYrnl4Nrj3bViDyH5pPciWPOra4/Ds0dF70NT817aiCkANcEpkJ9bJmjKKKPTZ1vT0m
RUo6Dgk7R15W0uAa+uuGLh5ar51EZ2ueqdsMT0djqJr6g/Jh4bviRWu8qzzFyw85J2r5EsAyeVsW
5M3aP1WJq7aZaJl6ZoAfmw/GP2GTvYIm6qZQ+tGdli7EK3LKwENRR9S2h+UJNG51NAeW6W3oIkwh
eCBvdX8Yh5DZe0cna24jEOv0Lq7cTOO++micC0i1nJZEMFGzHObTHTswt1RHb4OPGGV8cMWjmxAv
uzVQb5o9EKCx2o/MJvk/qEsOdh9GCxV3/AGtFoSU1hb2HxwVNGowUczzu2tiYskBmPSiLQrUQeoe
cHw7UyGFakIkV4Y66QOHMXz7EvKWjfoQBGr7hLWEb1aV8DAnsflRtOvRxzjis94R3r+SLSERkH76
d+OBvH22O8Q57FxFBcebGQ6vsWJ6INrO1C8Tc/jtI2uCsZjJnF0WaAQo8abTDtFqgxuYAOsic5lG
BCpK8V8c+g22vf4ZLgy24AM71QYa3FHMYL5A/W/SiXlmzD4VvLNrNTEhO2AdX/84+oKDWXgOVxd0
gizyuvfNn6f3RVpoigMgnGYJWj00E5cAOHWDteeASR6pz3voGOJVY7fjd4Vp8Md0jZ4n8LR0/Wrv
Ocnor6rSqAf3XoDN6mGra94r/e/qWfM2XSmjUT0SCkAkUYuEtz+9mOPE1g/DjcEYBnHFvzzSgmT/
ccGRqKH6gSyy3vB5SPb1cUarnOK2H+VT3kXDJBax2LIXiUMWPtYojCiKzwRHQX3gJv9S8JXBIdE2
ULZZDoTgtszVhC/Crv6ZSG8Y+5oX3Cazvtnt0QmMbrl10rRXU4FmzlikkQsKKbDvds3il1ownjtb
ILNNBwgccqFL17/Qyz07JJBMbIyeK1iVyPj52aG7PRjFSp+xe7OqaEoItdoim2BmqX3iz75Pb5pY
xhQPC4J0FIpixI2zvO6CW4AJZYeO9/8bX/R0tedoTcqL6ajY/hQx25/KL7qsmQ8VjTdbs0aTuDjw
g62CPWEKSv2gKzeQ8dbtmzZ8r35iixY2J7BHpQh2k040XHoDyzCv8bVEcgJ1oOxK+qDXXgZN/UGk
fYILYPOrgQa2NTUMFjiUtDw8XhlU15XjPm/y3nFEUPonYA40Xm+ipMZ+SYYODaQx+4vtlNLmTSaR
lH/SoIetTIrZFb+p+JImcRdYzaoR0wfIzPXhKwvBItRpgx6vIISvPgHAs5TqMpj25jU2VFOgppS0
4n5D0AdCcsXlP7t0xme+MqjOdHWaQq30vtKzdmPuWofiZaibY+nJFglTu3pwhn3kO9OWaf3bogyc
IMDuYc1ZadOZ5SW0V+XvADBHN67r0wQ+oySKLITY8vDtk6orXNash8k2KuzU+P0/GygmHR87ehOA
b8ROgcPIQmKJTzVaWGt/CpxaWS17wAqdwN51UD5HhgQT50LQZp4WkiZpTF4Qn4VyFQ0+DxFLs8jV
K8jJ7IYiCbuXPT05wAk12ojTRLN2JJPS1332nM27Bf97d08bFff6SWEDSrcXJcWR6BureHmMOoCW
/ZdEhnZsn4Fs/R2E7jdsJSaa1fnS5RvOAVybfh6wizzvcSsYhVwH4nIku/IlkB1abkb0bDzxj6px
1EtjJHyXHa3q1scKlsY72wnCH3CK5G58LuBDZH+MPyO/AoUf8d9KVzDuutiwJewZu3OEoo1BpWOp
Th4yx6KMTFodfRV3xIFk6liXR/CnjOYHt/S2nvDon8tZopvc0q6NJrShap3fTlZ0cvyd0gsXQVqe
WAE7RRExZj0hmDnoIwfmWX9y1ngG6SlEWfJetI/oi3KCAIlxDAAnNw+dw2wwl+hCPLIv3GvtA8kU
1mv+4LRgbJPsg80y8BAlF7E5SJmZmBeFPQKHAVqQcGFxkqOxD4oZNjV5GnLMVOBL1BQ2bTXizcvG
Uiq+F/VukQw+lnR2NmEzXY4DKdoO/mdIyAUukJT51vbZ3nnRVY7VSQlP6jez1oqWi/C9P34SBZEg
UR6n1GiFj00AnO8gLJIEZ9+RFXwrTxgos4FpcrztMPgWX+S80AGHUkdEoGDBT/zveg4b7a9XHNr4
9vaODpskanByzwBXy3HykR46WSzfaAVZ7E6Pz5vs5idVqKXBIYE4Ijapgwu4vaLYHW6mSqu3sO7I
cvOySEWcsdhXRSecm7CRRGRa+frs1NKhhv6x3/57hiZM4LvL1iHP80yY1K77yq84xQpFzd7qppBl
6TbBAvIHSSkQMjRXo5x6fwWf/2iRqAJunciTJhCfQHw1tajjgY85uCFcYmHDdAH8Jb2d5Y2otHZm
iEGDOgkAUnXS0+tWMwrx7NR76tWn2IFn5hYQg0apJ7MrcJ7MOGcqQgnCBwKu+wAxoGba2wNZPwZu
5JN13gBKk5tQBVYH/cMEkgo2ZJWockDtoifMUU6gCnkwaVB7/0fldsMraT9Ij8qlbCAF530hcWhG
zTha1AACi55ZHEjz3dC9UpTqtkQ86T3NOYHE3ikEBRRM8Qu8JcnL9vKk1fHt8hzi9e8n0zOv7NGk
v6uj4YoiaE/uclmVeDh4UZpiK+z9ohu/AyJ8sYstd79lfCCi3plpt6i9Zqd85epz5mohYXLY8rYk
Ar2/rvSOZcGESSwoAUsFQ07G9FiK5bdGg1gGEyG3U8ZPwF+0vFNIMbUie8PRc5npmCsUWUrOAGCH
IvZ57GFPqV2SZfo704f65YwPD4nOXp4c2wb23GfoPM/WRuPRKmsmIa57Ezauz/4j0C+RfM2QtpmC
bhSvy8r60Wbng0YTty0u2T1SB4nfjApkE/24USGZ7TBK22D+/bukpgRBGmygv7ii2Pgxz5QstF94
i+8kYZIf5dCEkoRR+QUDQWAqjxQuXfevt6R8NWjrUmxwYG5dJxGv0sdpDmlY8pMMhOWUf/8WSRu+
EhWAEneTD9bcrTNu+0YIMfGu+EBPPTQCl9vvtzujxoGrEwfIcL5+Bn+3HyF4rH8WP9pyU4I7AHTu
uXnSiOSF7A9vVLxnxB6frYyWZ9WBvbE/AdBl6U71JHU6I+KDbVcksTI6wQ1LWSTx+Ws1AjB+WQS6
MtbEQ/iRg16XLIaQOmdzCPGcG3ioQRrYCzojF8ixQ21IeiAfO90kg4kVaZ2rtQh7eQVBZycNQ9A7
1qaWUa48kOWQgdyca/mVIzYwPICwvzL+0Ls5hVM8jk5TRS2Ws34oZScbedPUTYefPKqL4pTYNakL
qXurBumvl/F6VKB1W+laX4H+seS2OdfdnLSvSndMSxeEjuoe4yEMiMdpFVvCCG1no79ahklU+sDH
v34donPiQ7vwjjwQQJ3+Zd01cB0CmuPBjMl2ansvylV0P0/6wVymdVy/Ijq0WaRFhvxArPjxX3UZ
7aD2jk5f24g78u6RB7hZrRKou2+HEj4ChiqkCbIVBQ/nJ98fXwbN8SpufArhbXRBxoXRD8nx2fZy
T1hmcA9xA7vg4zHFtVsUZ8Qj4sXobLzIeraUgDv35ah8wHsHB85QmolkJxgQTudT52mO4zBDn+3D
hOaCgewq/8Zr6D4vf+ePIK+E2Lh6g3GzKyiY21IOA0l0JwVOfID5xpGcB/VYsMOL9a5XhAr0wLa0
hj2PXPFZc6fdot53r0gR1X5W0s9x2KUnKFjmFwGmgYhEq+aGcZxYQa+Ju2gSZ6Q8diA2mR/aJ1oE
YlT5AasqF2VrjXqD3Da4en1JOi73yLf5F/dp+2tZcoSzPx8EXAbZXYpP9xY1o1Pkzg7WDBeyNIPm
FXkoDVDh3e5ZOfxf24gsEcO4piDn5eufnWQhQp1HirSSlwbt7J3tfSawcnOcyD3yOw1RMijRc/jV
AD/a0n32xmdCK3urg6AHsy3qClRKEBI49Yh6zomO3UzIoKHtWR5yWBTUnuHuF72owJ+DMhHwfSHT
WaYwYRYQVYXnAkevb5+VieFiGG5/fp84NVYe9bYE+y0KI5P5dNZvq0Z2i9op14Ni3g991Qub5p2Q
96aWOXkISzKACs223rQzFjGSvcKrGwwqQXhAiHNGG3nwn07U/WbhVhB56pRIFWN4d7OxXpAu1OJm
+2EpdTIs3QiRqNok91JzDOFfaDZD8ZcZ5Lf0H+JSqpjmOY9o2JfzUAJCwfBYaZulQfDJOKM+jn3H
4oCdhkLpUkfezeusjKMxJoQqaiXx0VqRI5s5zxSNx9HI+n4/gY8lUsgEuaieSL9ZpuNaLQIZexFU
nROtYB4xfLFz3eX4MgkdRMYEDy2lgXSeLETUsQu0Kk8juZE8amHFhfpcPH20X/F+6OGDrJMZ3+aa
g/bxUxHWgd67xxz2cA9/fgCf1+DgewfRC6ULEBE7QJOIPH42rwGqJJ3ayrDThsKJbAjrgJpY4VX8
MfzTeu7GpEkwBAZLEqtjPEXMWi0gEwRdol3S4bfJfH3zfhL5eNEgRtUqWC24cxxemENdfDPkCcIi
HqrnKNwlGdWzo+ITInWRemPHWjDJx9X8kpSXQd9r5S7FJmgyN207GTzpxDNADcDudGcpHrsPiqIh
Znyv+UkSwc78tVHuDJj8dl0qD+HSyKgvQWEx1JXR9c279f+5kqIakNqkk9kPCKDWmS+bbtkHQFHZ
jMfHa+AzhUJkIpaCb3gbaoclnyz3Fnd9RkxxgLRpp/lF+rBt+RRU7qfrW9GfJ01oKnk8WZs3y1xJ
NIi4gn85JX400MXo11naNOF3fB8KAxjyevuym3+1QFjLTXoLpvE5ktuxtc1fh7/shNmhFuL7y7hv
bqqNmlHZDWKxfv7szzpt9wDBIBfaBMku2ozOPiZBNsWIEgiOotUlxhoO1oihcxpRREZr5gImWpbd
Z02eAhY6WyuvzgPGIfHR4z1AxXSEud/gUinIHjTrGdDeTmC2x12dnes60Cc043rQRxvvg3PwiAN6
m9oOCS31eWS41nF1FdYQfI23jCZpXWSLsBXuOG3EHMysm/5pIZil5ajNfkaOLjYMxP6tVSj4h5Lc
fncvRjytatNepP0foEpkb7gmeSML86OAF5GOSBZ5T3LHsxnbm+n7miSVjNfSfkOW6E+DNSTm5RLF
9q39GU3uSDeFXkfuVljxahsj0QrqnVspEfD88rqwp7Y7HC0UKIQ1eaJ8IxQ/ktDeH1z60l69PDOg
IX2PImdRRAYOfErwQWgjy2ShOT01UOaFW8emzM7OXJJgjHvmKXxmDd7YB640P9vznTULeRsMw54L
khUJAdwmYNIQOpwJrXubzzfmWHgduxlSCmnEXIz2/Har1bQ4z0KbRQr9bOQTzexHgv6jgaTK2Xqh
dGoMRB673jWN/5L5ZI58aob4rAG2P4RNxIWqIPqRFzfXf8eHiRpE3ykRMSZ87Oa8onlod/aGTxTn
T3/80aNx2jL/Vkto+SS+2M05vXRvBlpz0g2DLXLaj2kqZbKrRfbngktshArj2sO7JAiFZgDXMl+T
MVbeIfhWv9pcfeS6OVLMrpxCjUKoustr3U/w5kKPu5ZT7FWdPguWpwveMFTvpCSaXzQ52qP9N4nA
VMZzi8c29gnrTDbdrWznuin3WJpzNH05xLJSS1B/5FmGYXeVgz+ye5vVs67b6Y0USgNMAv0vMpk1
QeDqZ/fQeV2F/gRQfM9ARRmU5FZSFMvjxH31ov05E75xwd8VHMUXEMxBbzLgvysSeP4YV15ngBnK
awyHyoED5AUz9A6gOEuNanHdEINr5v9S8FSiUYpUYcIsm+bLyO3ZtSoZ2UUm0d3g7qxJ+Mb19jwe
zY4GM8zpzeweI0YFBIFsq+HeK/VqQhrRMv1tcl3bW4/E68Qrf87pGXrldLE4jmFBnJv9eVgpAxSN
IcZy31GYVBDjkIOFeVFJIeOlmCkJclplYgnjB1ldgdRc8exb8zZ3p/CjercPDzKXADEGOov8nmIJ
zb3IOlFpU+jk4sTg4sVsVpn+iy6+soiTovBXla3Bgies7ZIYNQlEUOBAq6dWBEuecpNfYj3nJ6dG
s0GSptPQLrz6pWIQ0TDvLGtenh/nBbkNpDH2Jp+mc5DwD+/XoHpqLUHv43vFTNEdH6c3gi7EOHst
43Ivp/35HgqiduJdonSCOx+WWJ+ACOXZpRuUIpq7ubcQY2ZAvVL0xwlMguhAKw7Tuj3u0YYjGSSa
3bBJ34xRJHDGIRbFANBsa+et5ZOy2OTStTfuMyXE49ZWbmDGmw4RuMk3HzLZ483hHyw+QvjXlXw4
CyHngBUXYiPrX7NKtwWOxQYrHcx+5OtySXCxhEuee+uDMY3et3uXWniYL0XrtRwFd/79jIZyYrtT
NKctc/q1bRF6LHOUIVdIYP9rvH9/WJhlN338DEKrmHg7R950oaT4RQK1IGOs/fRs94wfRQSCg2QS
e08rBTReCG02BjA/v495XX21OS1rFK/7bQOasHjAYod6uHwWIZM7EAj8xkm2UHRyXkDSb7qkVqkh
4Ihr8h2uT5fmsrQ4x8oRelreESinOO5Nb4zZ/6cJHumY6PJXxAnYrtsTgDzn12AaxFtqYmpocIBy
NtjtHQHt97M+C9pOe1YEnhz0fqdHqalFUR3LpjogO9Ve9LUj1QpizSQiDbay5kvXGLmAtFUW3jj7
HVaqcYqCmwR2iFREEDai0fc3JxJaXUjom2VpgEjr2hjCfePhmRAp+J+e0IrUYx6gQHsjst9tL1Tw
4dG/g/vQgGXTKoLBKH6F2EVxeSzL5PNnVRSvPGD3R6r4YUOUtFuSz3UGEWKFjP0wMjD1nhtL4O2v
jdI6yAiZKd6ZJcyFxSjPKnTAdDEGh7FSy16xYsWNO9/gQ2DKYY0WzNbVae8zjrAex37L7MzXBBWa
e9vbdMABYX/yNJ4lz5fkYqdPrZIv1UHumiV1pm4tJ6prnhYzUsLugYSmE9+q34O01rGkylZRiazs
D4ozXHpbuHSSddPuAaWENZEyIlJSURRTMGoTS8aMcTb++7BsmN5ZDZ/9OTl7BjOhM0UA3Ft/AtR1
oO4o7dKppQRflET2QmxIgsF+WPkBJRSowyv9zadOESJyr3Ez8rr/v/hvaXPzI3V/EIp7yaeeDVbt
u2Ic65HqWrZQfDl2idEpiLZO05SGw9dab/Z5+KiPLqmqcqcBGoqtB5Bd23864Tk6SGIeITvcX8DN
3yXsMpvY71TUHs5/9Nz/Wt94+oIWDK7I8FEa6EklRGdeyYgEbxHFEluBeY1+ncZrMySYa3U48qD6
Deebeuf5Y2MugXP7frVm9bL8YauIXaKIRKm1Ut2PHbbee9C5hI13DFsoCUUOr+9nSERPbJGMhKpu
7F9UYAtn3tC7DIrQCmwVbj1fjN4xA1n46UCFQA2vAqz41IiNCRq7xhnKp4ypjgLFYbun15KDsDO/
K3c4tnkcpAZ5lfiwG+iP4H4TTlKSftfY2I9jFysHR3guBLDxJ7eAiPLVIKIz1rtuL6T1NQzmnvvx
c7qsultA310b8kq9dk+Dx4k7jkXLMJx3DMfOvNO70kGV3M+Y7pRWR5Gh7oMdl9ZAL38wATucARA0
tniDM7vDDvXFv+n7pkFgQjyTF9A59NMtD+eeQKgnLCZ3X4yBwUdxKK9QC1umaAODrEoku2Gc5vYc
ZZ/HUO+K+ozluSiGalj/r9z/Dm/SFe7xyG/gf5wKjeXURUXfLt4t5Dru8ctU0rXDp1rMLLhq4TJl
AAap26ANvJnZZjnhmMMkWA+zUlk9Cm4MJiuXcbQHd1X1keO8JrihSaCvZ8hGgiuZ3LavU/BYfYE0
svAAr2T1BGLMnuRfDAFm/II+2e9sVLHmdWgX7iXa0Sv0voqdgSCkEz+l8J3JFl2KdNqS9Y1Qn/y+
cYJAY/bjSXoSAHz8xvrApa0+586Zpl3GiM61HlHsL2KgiedOUw3PEaRqvlZUDrjCSNxE3H8AkKH0
VNDu/ww2bqFP9gztvqUUAt0tNUDXTQmjhHQiOlpbURdXELwigLn5LwRPzE0d1X8fQ2g1iJfsTxMc
psqitp7Q/dlMCiTRFk9nOv51eFF5IIO61YgdSBY5zj6MN9a/JX07k7T1yUCKW9ZiDQxp1kN5tFb/
WdudAHuOl66TN3OZ/Z0aubmmXJegNCDXPDNE+P9X6Xg7iDMNGylasK54876Kw9KJ7bmsJDeRE1bs
bg7W1j+gTZ9GijNZvA6dV13azQlZWYvkapoLegXLINy6g36Na97fVsQuBtZ4CscV46eDWIYu5dol
1YbTGHgRLZS4qKmnNaD1iXSgf9+rVPLHa1Jf4lGwq9yJSyc9PZEc7QwJUNM9YjkHh2EEZK4sp12W
qCXbUppZW7GY7MoIifFHtIfsZojky39VLFxro0qlG6fhAhTp3bcHhiPSvawvUmCicyD5EdbvGkiv
M115d+zZnTn9uW7eKjQ8+NXg3cLImNPPSlIekZd6IzVQ2Ejj7pan6yCgPyyPXe7C3c9zhBpo/Qs8
ov2ccRcFM3QH8iCp3gtIIiG8UDyTOlLuVyPWokPhihwRQvsrijMiW/C2Hgt/Io4jWbT42H/f5VP1
5YPzwyoZZwKNJy7lhxA+zXNJMdD790hX79dcPril0W07kq56X5JROZQ2kS249ALzYG1fAUGnL3AS
NuD0BLS4tNlSJzwlW2rPmyZ3Wzj3zajR6PKJ4gdaHbd6c0qI4EtFFo0A1L3qM5DdoVM+ij5aOCZG
kXyiRI2kXvbLR6iD0tqhqxa1qgsLwwb6pOwhSAhy7uQBXN2zUZTz6ZAKxRZDd6ZqoFU8u686csYL
ANzXwxwBE8vDa7YFnSrlAh18cVZw2TpO58HmECoyYyvDVOw5T5SM4xB9I4w8kNynDTXBFeXsLV6/
npYiWFPFdOpv4wNDpeuotNMiC/1yZwffuro650SRdFFvOKsfz3Bf3HPDPybGv90HnHHJA54VzIkp
yJLQVprenLsitAbz9kdDnpsV0qNgJxNslE7CQu7mWlweVtHTyQV36dWoww1EdATvkC4HpdL8ZeM9
9RwZbWvFCFIlpDBFF8DwT++cpkObQVS+fpnbbeWPBMoYO2ZkwiZ+5UAlEg/hAfriHCPhisVa+UWB
uttp2Fi8LoRJh8MzAwqceD7ixou0ikbaqCwQXVIhV8KJIB6ZIpVQYbKHX3y9g9hgOoUOLhGP7Dpg
ZndK6i8OYShh65wE6mz4UiY8WzCiUSIdiJDYAoPnBxlzfGsqzTGu3p9AafJnJgASfv09FS8zVdYb
YhEzN7J+XGlxzScO4machhl/+RnIwlgMKTSILlt/WdB4xAUEgmuu8jDgh7en3SnRvRMoyYbSLOHV
lavezrSaHt1PTTpRK5zco+HIqy6fo8KO27ftIHY9RUAgMcMybLKFlcZ9EEXqY67Qbf/T1umfWaIX
mgBKF3XoXXtbFObIthC6Z844RMfI4ADF7by9aB+CfEfmtnaP5f4zESEnpvmp50Tg/EpssxLxb3yH
GkLdJC4MpxTYj1VG+1VfVZ8m8wmdujME6/NDY+unQWBuDscuQLoWLw9+EvGSi6UaNiryYftFrzjE
nKoY1r3xRSaFdDaVtwXgAkgfUFO+4KYG1phxZwg7loU5/RClg703oUlAOV6fJeoYWqqkz7XMGyqP
asDolgpI6hBtTstmfHnSae4lbK2C0IzD+/m/Iyp4r325+V+G5PYh5MEykSwAOXhhypGYyKyL75b2
4o+Ma/AI3Vevy4mi1/fRehaKPrpmfsrYvcqVxHH/jrSMkvWbO4JUOhlxz0j//gk6qaaoti0fPvpR
kP8LGtz049O2oAq61vFrJI7EEdR3jwnt5yH3jHpQWqYwF9iEG7EY6gw9hr2+ra236CfDU6PKvBZf
fIUNw1m/qUAe1b9X2tAx7C7BG6A+Bva8JjoafacNrA2yyG+Sl6wqV7EnCZYQPnEi58fgkO4OpeGz
aS0e55CkMAXXH1BLO7DxBDrrvep1xFTzpeqUUFIfArm/V6xcHcaLlAXAR7ndCrV3zNsNsT8xnOdD
WuFCSa9Ra/7+D11GVcupXkgSsGEZsVM3b3EQltVR8qPi2X0KhyD1PsFIhP5xUKFugwLANTRIovhd
KUibJS8wkglqVPXzvaUVlWRN9i4SsB9Wy7LKHu4gN/kJpbIAi7oQgOtl7ekl2Fod7096Da6gM+UZ
AqMZ84fuaY0tM9dNfZpILhJwRJc3rMrkXpkYO7eIwWe2gbM9Vpx8Ct5fXrdHRvMJdL8Bt8KFO8+R
rdhuGx3cmd7/Xy5t1VxtZOZIjTirRqrCklaHvNxatbsXyvelaDJ5SsS3OiG9XotSIR2nddQfLTUR
Po15CQFbAFBEi24sT5v1qf2hxPBRj89F8BNX4W7OMd0BwkD9fZ2L/hHXMXsbRXlGkMs2ZTaMYmCN
Fc+foETRhkz4NBlcsk7TocSz80iPdzPbErA5km/B+TdEFFuvyFppXgtG7/v5/GlOi2L7ZlKUQhgJ
DhpqEUO0GUxtXoUzH2JF2qwhigTxyEkxoEh79e7XNEWjD+ZXfuuimE7iHmRH6BJamz3ORWv7BaVk
rVIwmI0NplX6bXl8DRpBwa0v0HKgx/TFZEIr+SXHAfiIRKVdnah9cHjgocxfWFX7fgRrhTirM5tm
Xom1fRwXV75wJ5jZGqUQS7WSQQOPnw/9/5yNm+A/MxbHE+/lL64ifNc52NRKunehDO8/kB8NIWMM
9YA88uRzdwWsQ0pK6tMQCZ6y5M86G62ARGkEoraM4Tn4akMYFSF8Pev8Qf/lT1Ql/ANgfXgnow/1
zFgCTm6EF2Sy8ZHTLB2L6+J5sylQJ46hy203x80HbzumcEHYq2JsYivcaZct6R9GHXAsSr9/1/zl
YEOCDykH+Ci5ERUEBQOk+GBvmZVA3Bw00ehQqYkMU90mhbNye2Emuli/zyJC3FzgZfrk5odgQB5H
vHVmjj2DhlorIq0/iXZkN/GHv+6W2JQy1F1iHF5A2AxdCo8u5dwTZT4kHhjc+onxjx5pWL86zZFo
bWVRKjcDzrSigQkpVM1MEaUioEZeIJbASxr2H7jYNoC2CvS00fKEeg3/JT9oNHtR0tFnxRhz0NMS
oXSte2JBoyZ1K8Cbt1FCiJokkfGlLL4/qp0v5iXvHPtfYted6vAeZfUWh8MgAsoLvBfNy5Npy1mO
34+oNecv/hVYGsAHceUslYuNiGRbojkPxgbHzdpJHOnjXDXobF89tdaPXYuUd8ANydWi5vHG2Sv+
6rrGryCZxU3Ji+uAesFDKWhtfqF5PX02GFzjArxa75uOH3AyOgCAabrzqcVl+8p517cePYiUSvXH
hpUo2rRcLlmvAGAUEs/7vHTFCq66yIFlARV3k1ivIKtWViS4GxmoddL8UaQPCxfvrooJGamhrgtC
PfAHEn1GSVQh7421L1zosxG/R7Zl34IYFz/avF0bP9myeAHcdrg3I/Ny3tCF4JrfR54NginAhwUN
SFlpX+e2kiN5xVtCPkM+nL19+Ttl4NgdT/JiQdny3k0it4SNF7MuvDIT53LAbh+OBRIHovtnzCAM
IgHHBoNcrlKNaS9jA4AxA8W4ZhqGPHHuCN/OMrMie6P30pW4NakyMD1gdXG4w2Tolg/IFCc6QYYV
lAds8ZJ3BORilNP4LdWRJp4QMY6tuOo80CLyOZ3oIPFLgjZj9BRxRzcsEh3tdDNe2xDXBjeTBFGn
PRFFbmurj4t7v/bORsh54pdTJnZBiCpJ0w4AUZb2XS3NB+b7g+9SFT9zrjItyHQOIPKlv4DRij6c
73WHp2L3qsODkbACAIMTLTl4+XelMLA4mIkYiT2pScOM5HEqt7jaW8+0lb8/G8iNKspsvroK1ZdY
ITeTo+kQHkMNcH1BffzoinqEzf0co4O9KTBp6nIsFfPCiPDQhZhmHkexFGaPBZH0SFUMfcflf/8Y
RhRbNdjwWebBd147zi8bmtp9odDIIyI+AKrATuio2ns7lbrAaNUQbvnqKtjkHQVxJCtx1sPZ2beb
OaWocFX4VOoQRHV5chL862X+d0X8384zaRz7fMbO5wqqwwrFFcYxBczMYa8x9e5yXDmjKy3J3iCh
6OZc5UcFBv7Kh7IuwuwlFJihwVMS3VkC3+fxg6JzpZi7tu0oG5D0133GDxA4taTa57JqvGtKj42d
9Rusxtm4axr4hgFX5L2T4tZN/qFM61gXQAjyFBlJt+DB0r+xj+KUvMzbel9DJPFrzICqFfIGEZyG
ZeIGZL90bbRA9F82nXpl+JWHW6QF7GDRKLS3X8mw7UgG4mK0V2GU81MQO8rTY7lCcaAWgib7uqlg
tFEpNWgLZSOCGXtNpvwiDatq9T/f5Jd8IuJl9ZDjf6j0QhxuolgLP/59G8/4ERJydVCjy4wcAB7D
9wZ5han0ElgzX4gAWcY2EYrc+ULS6l3IwSofVfNKltj1xFfeD0RWsylOTmUzjwCJIy1+lB+737aN
AWHT9arA+Z7MgC9jUTyVNRITiQf6eLC8iatx/Hf1ptXT4MxrdBJi6zq15SbgGZ2Q1UUOzS2ZxGxN
Jrp7vwTNsUdSJ1TrHBTKhPyIf8gBurQCTqGrJRRNrBAXBgsaeS73qEwE5C0tGZaLJiTfb738HMnJ
YUBk0/MbjJo4m5AWAfRFHeblhRf7zLpRQ4uBWmgeoBTkAQq/+++3G1eCjRVAaIwTkLvJ4s81raUb
KO3lE+lIB09JxmMpx/ftQXp5JqYmCQB+vVaLzONVfY1s9+FV9YEaqAsLg8m9DXUnRiYqXzJqD5v8
a3v7UWiCM4K6LCa10/hE8GBWBLXsmrHaHKXmbPV5/p7K7814JKLtBYxK1nTa5M5zRr7sqxKNb174
yZCXuWMjNdXR/mo8frrYXFvrYvZawiHvw3i/Io2kcaJ5k6lcl7Wgli8MKEvM5hvX0S5guSpHeful
mbgECmuBjOrb4FFe0aqf1hwsELRZwb2U+ypTGktRXaujmL1DNzZ9mrJjzLxxR2ieCX4XM8myeVvd
BLe9pGCCDiuoYOf4J0cjEyDQsHj0ZjIWuviEj3ZLER/x+iLn7TbWiMmXJ0qth/NVWRjXp4a0V5ce
6GUK8C8R2jG5kW4j25iH+8AzoKZUwMD4xjq9VTxhXHxKAMOBlYLipfCuYsVyUFpsxPKC60NfgR1x
ExVrZhTauFVuEYNJ85CcRHWEDc1W3nc53KgIKO7cQc1aOs/nUSOYQ36MrrLzeaogojYPtr7XK6Cn
G8hn4JspVddHUbFbyYVJIGGW7pqK2mvbQODP4+PLJD8JEK9ZTmg6N2Du3e9A6Je3YpUGAPLwrpty
h4lpAQTqba3dSlDqoxNbhLgBydJUGkLbhvdvtlm/OcjsD2rO4pi0zmBXmGaoa+xBdDMmgxLsSfP8
b6soobYDnnRb1WghoECTgSXSlMprjcp7+1vAOEsRfsPVaM10Z4whNxhWPVGT8RDV9YdusUsBIgDi
RwkR6Vtf8csNxqrie8XAdZmUxR0e3C3yKOUlRLmhuZG7mcWpG2JEeWYXFzbvcylHwC3HDVYGNFGh
RGoe1rg2/qqdOs8K8lFrHz/kcLLEdMIrYbN4J5I9VbAuJQ1xAlh+H8aje+5MtfWXDbRXDHPxBa4t
lfaFzqgbwpWM/Zr5aV6nIBfbL/Yre39+kg5FRdEC9ErRTzX3iTOms2j1Tp9tAWm5/CrzOmSqgyGK
AGjUI7vlBJrYgTHzKqF7OadYC01xHALf292s3GyhKpkE8oHq29OZF3QlW3Vgz9bWMz764/gpm9E8
DNTmj5NcXmVIpTecE2vH8jLuvTPI2hFhvv1xmjQopYRoSTqbAfq+GjZUCxVnsWv0dGpRqw71IdZ2
Lw7/VOg3anXlwrvwAh6gwdZC2SSWClGUMTmc2NzN4ujZJD6WeADGNa0aUOf2cR5tIySdl54fdfIj
+ehHX6gw5qI10mo10b8+t3ukXdjVr/kQ3fB6mTSBrBHeOP6aFhbXfx6gsbwa9dgEET3ANB0dyiRc
7X/mxNisTXz4TcNsKyYMo4IcNiz6gAODetBL6yPBWrRAFgG9ZDKUnmL3Lz6kGZwDVkGGHCMv3QK6
D3JP+pXLmUzYNeZVKrsHBM6Al46CxiuV7nWPy7w+dI7kG5hAbfeEFQ/C2h0FQL6Klu9h+6djJxL4
rVDsjehHKTaHsy05WXWLhtRrzgN7S5pKCeE/vLWGM7zpZfqlHbm2+nFGAf7xSPaJEdjdaF5Wyctr
zZo/URgIJBH5IQai59Ln2zVWzUFM1RDwIQDnu/7LW4jZ2kcpjQUvvDsHAZEF0/60jK7DMS0juW6B
VmfTxwSYto83xKKMixTKkjVrN3HV8KRPO403p0SGxjhmA2RJLYDGmbWzaOiKuDZwpk3uRsPwTTPQ
mhZtLyvm57zCIZk0KjtnOS6OgcUGS4a00zaJNXliS2IaDi7v/xT8C/IWOuxfad1FrsYYWZ/9rwur
I8jvi7yKR08c25CO2oTfrO1970ElKSMWM7bYl5PhZoET/sdr1pEdRKb5MDaDHEjcBd8v7xfGNi4X
dNd+7ouUuW5r8pw8GWtCYKR5yl73gRC2GEEE+yIp/uO/G+EcrkmfwHtKaokB7SL0xEzljhk9fPbl
ixbPXCU5+ARHHU7MZ1rLXeZ8alXkeAKmbOhTpHZ5QcR9z2Z2lfQSQ8bcPmr4vcWepgEEtAuCiA8i
Wavr+4OXTH2S5fOBGdTAmmjTEIU4HlVDjZBH36CRK6NQ8EZyLRkiSfNBbNbnin7zev2YqY3F7tA1
/hQRsAK8vWSg42SztbS9D/FOJQUuWNFGMZYbiVm7pTNwKVH34552CX4+OvIV3nVpITQb/pkTDbXH
8sjxB11LXny3q99fIWeSl1ofK/AUkjmCeeuPvRE9pe62yEMtufFa2bcm89o1b5UeCld5exs8HN4p
4oS9reDg3x+/thMBDnkXnm24Sh0GGbHEHkqYtwxli5GbhxGZIASbPsirkygeWVrgupzwI5JjDJfb
FTkPIF03Z1StN+Q/I4g1iZE1UlYFCJ1Zrdfl6mCnCLE6yRtD2oXaDh+Sk/4T2qHSYjj0rXfpmfpC
Lq7aSYcdGKowTtcpCdtDLF3+erF8w3ny89HuhTRUosiqra1Plfoyl89Z/YOv2eB7Kqb+GM6xJnZW
If/we8jM3oc0nwf3bPSQsf5jjm7fLTyVMzCe/W4DfOWPaLdx5dksg4T7hf14skru61WCBBtN55ML
ClQK5+srilkrIJaSpGgpnwujAz/kcMoD33FmRN2YcrcbXpkdca2w/0vrcSFokj7yNBPH2gbUV/NR
IRNzGfqHt88CWofYeXlaTZMY6KvMpszZvGWZUslJukA8PcaEakeGPmGXtKhelNhL8t2BHnTFNs98
9tvxvnr9W8UApQM1qAkTGUifm+UP1xv09W5PfDXs3n9thelApzNVF048xKECIYOPptdbfiAbQM0s
4qm76wzBE8Wv7amQbLhpqyX+KJrHEHwE/gqeMemdqnZroa+/ZW5kFtyGXPQnd0Y6ejXYvVSq91MF
GiaZ0CQW7MIe8xShgybnFUUFJtW7MytK4G0UcXkQN0rdnTEEMYeGyZE5xyTSBA/ZMGYBapnzfCez
2vlR24zbItZ4Qu7NBZXUgkthsGsSQssEsABsNhjrEtk/s+s4o6xIoDNNY8cKGGPUZp586MsDXwWa
+AfOTDXVwVywitj1ZnuxwB3tryp0YCV4Nk94qPGKpIPf2CDUmsYDyYrm4xDYakp9w/0NTWlKdTVp
P/TUwC3g7YpMcQWGoOOacTcVGuVhBQcqcZyjhEV2IEfcpKuX6PMnOo1FgFeFvTwQAfDZLmFpHwUb
S3S+M2LEqTj1QZWlv7CoYrxWu1Aw3H+zQKn5Fdjh6b278HNkiOQ6sRLOBTa6eTsYQJv9uFm4oUhx
1OY9qzpUGDNRgWLLeoMJoXKKBY1UD+pG/4ICuV1gzHxsiCPiRoJ5kI3DOlGrknCAfieSwtxKHy+D
E8VU+hfAXOieCv97OmT8l4tjq9JP5AWc6UuUYRdgJW2O7uZFfOAOHnZ+Rb9C0+B62hqjsrJlUhZh
8Oz+MUAxeMnDVYwnpe9/Um5XHUVUEKEj33mffUMHzhvCcVCCsy/AcnxeDaG0dTZPV08G2d4BuNgW
Rbqv2K8mB4AD/NW/LZz4rt+gM/vQxYGjkbB8YKBBiCQ4Q/0wqrtM9amNbkun8SlTMSZqjJjmS4GZ
iow3HeuirxyQkHsi/SP36z96KTC/R2NqkfSWc5Vcn8jdZ4F2WqZIuq5Rft2kjkMSW8BvaB7xRsD1
1xQKT9ZDmlO4ScL0axqS/eNee/8RD33w8k8EA59nENk3Za/HGBc9ulhrsRRKrTHv19dk3WXFgpeb
LQUhfWRy2CKqwlI1i4J4EC8ZPM5mgxBW2BXSVy/2vQpwtDveff7FOov4klwVa9cb/FavdHnNpt+R
RzxBGlKqmWSG/lB3JR43MyJ3/9923ZKV4ZkP+JifbDDevj0t9r3bfD6TbnoY4c7L9ged9eCva1PG
vbgJvpjxMUqk/3DGxitINOeK37CSsyqtFhVwuwRftN8ayNAPqlGicNCbT1VHaCoC15QkDmOibMHc
VwENh7MIDkK0tIc/ZP2I8kUupQl2WR1qSzrD8/o/Rb+Z10iNUytthaaKu2tVidW0PCv19+bBrKe+
RRUJsC0GJdUwgDIKyi9d0AjFpVG1vjQ9fve4Jv+EWazMHyMlxTxINBICJJr7viWPsct6lqHLsEMu
/Oj8W54CoIr2oBPj4SfjEBIX/e8rCsIMfXPUGdROlIBmDUUNdiiwE6FRX2OxQLEUQlrqWjMtilSB
coDWKKoVHG8uSLTvQXC59Hp1AoDOYYetqI84nfxtIgiDqAUwFS6yefoxkWyLmy7j9z2LR9JT9npO
OftHNfroK2s5fJGsuEqxAM1WIhYCKK9UUAIh5aWoFvfMjKf2BesAKuNlO4+IIBEZfl5Bd584T0Wr
GVWToJhiFnNSan1C+ZTNNROAjBcIQKgDS5vDCLo/qX4fHvj6ANJQ7YNWFKOkNpRM4AUnDKxXxa1v
NBPXVTi20RnHE/dUJaMi3QXUDu8M1ZV1XBurjp6x1NK9mucf2aADjI4AwmiC9jZcTFD5nOq2g6zM
KJPdtpUT9D4kdtLnIqNnUBwvDktZmTTWPF3L0n6SW2+/qaIhn1ogiQvq7tGjthhES80Bdk7SO1aq
23joCkuVbrfKseRjDkL3yAkqJ8qDAG0cMnSw52en/qlAW7SgArS0WiKQYS2Pz7kSAWuQEdgVYtF/
4wva1lodPjVoN9P9NAh4BFD2trrkcbclkMz56GecuGyveml4mXj9ZyuZawGCiSeNBOordRmjDH3g
SUsyAcoJOFA7o8kCeCq9Q5+5rJNAvgD4tWxxNbGl8h9gwusXZRyd/2LJ0oGsjLpVViuGavIj57Wp
eFlvzh58JbPPsdYGS3Nl45QTeFhCHg0n6qJTFWrhh2pzpk1M8SR3hpefFp+0+Sn/0hLtFnxmJWsw
bwKhi6Zff6fQelbMLGz5IRrKeH1li9y4Wt8lOGxkW0QCPoS67ujeLZip75cs+CWCsJ+pQmE2hgSc
OgVcPBnkDgS+jiP4AUx3Rtc1IxRs9zq9k6GZj3W4wEkqU0RbRfGqC91U3xpHRcP6wCgRDElfkIMA
gMMAf/Gkbb5LShIcF6ySCbaBwWIOryiDAhOKSY1JbIGE0DXKI+Mcc/mQnQYLWzYPqZVhzTciHzos
RCpQ2XPriLMLLtgnbxEubbgCEILsmH59FMcJgcpm8Cq1bl1vVBoeYjr9L8wSogxzZGoog/P/I2fp
E+MxPu/Tg49LMCeIREnDjudDoAb4DD2VciPQN5NLOlYkNER2JuNnEjYT+k+Ykaw/LqgJhnLkLjN/
RVikvrk/A73nmVdDoN6ANOcnVmR2xV36ANGcvLs9KXbIehV2NuSrhHCfuTh6WMU0J/ERsgKZy7qI
qEtTre8R/C9EEyl7a4u/1vp0Vxb7u6L9+BJW3xsXKzXx3KK0FrYwQASWV1H5/c49M38e4+UDUkhE
EguUc4+6R4KQVZ+T1pL3LeVPYTLdO+uFWWf8XQvWvSmTqoxLaR5AouNNE0DjlHo060ApigB2+VXA
oi2fN7wiiMwVzISAVYu9yHQEbiEXFXhAG2HxSi3sM2DlkTB6icL4CijeFxzYJT3Fy7Umsx+hZwlW
xogVRuC8t15iK7VbDOewd3J7688CgsdCp7NsZXagyKt+8TGUApmCeYvPzwlRDXVRdUAaucsB59Wy
9sDruR06B8lnPKDssrUOD440OhRQyM4piHH6TxPzQa+pBIAtrNUTFFpie1P4XWg/Zc5Uu1/uBfVI
H0wTR0V+autUxYH2WvrUPNJ5r/17n1NIkKC8zT+w1BIPSjPEipCjHnurQH0i0Gnbti0QJ3fFd3CM
kRvb167wApfwx28+myw6XPtJ38NaFGmYzsfJES9RkKRauUJW9uS+kLKcI93k61oSMiR2K6sPXYpX
dU5FYjutOcpIJUtScmd89fOSBVNnz78vZcU8Pc07pWgtzjsxGuEZgdinYqkzLV1w/oRIUMRyAm9k
xQ0EA89tFDAEJ4+DlJLPKmsw4Y+JlIqepPbLlRj1Z8Hk0LYZuk9F9HD/rLaUrdKiqkEKT3MMAw/d
VTEjlpcaBdF+Kp3wnOoeDnWdVc+7EORV16Z8tUCim7JZkZ9mXURaEWf8evaz4/25D8dNLlm90alz
fR7v/+ZdQM8uDy9zDUnZc310lhpfRYhtXXx11l6oN7hjgCDIMefSU18XY7gLS1F+nsHylLo5+rAZ
8fEnO5fxBzEY+R3VG2g/kPJwFZoH1mRL18mhsfEYZWu51VmeuhOEphP7trjHfCnAiEAGaZUCq1N1
LTfmWQbZt6SO+GIQohgKjmc5MdqkGV2wW1RZOOeArFKhLTOJ2iAYXZ3BOsxFBOL8kXtOoXMLw1Yn
lCp1Gfa+lM2fsRTkAJfAspqW4coQyOZgnrtsLV9eodOCh7mivdtrCOMhWV7ORLwMqx4KyrERXlq5
/9YBZaygiwGK4iPjOAbokf3ISffx15X+/NtpcXso6rbd3mMeb66ItWaqoEfBFBQDSFntDI2ZJZdQ
4XtPqd7zHMVVb5xp7+ByyCKh4Fik+CQLKthsokmhMb/jPKkj4tcAQdUwEVjggaBDWVtX8/kBGS8B
3ZSwT8ERDlcykB0E7kvWqEWozlk8YkcdWzbpS5Q43qDfI+RnPhXEtjcUOjv0RBYPI1sX5x1SNkmG
43RuhrqvjZpQnkdP6tXX6S6IDcUxMnPQjjkysv4wBjgXjj/j8xwg6H73vASzcxpWKioZTev7SdLf
oCx3bHsD0JY1KB8SxZ8Py1SZLoAuF1TfT01JO0HgSLCTkQzI5YH3YoJuI9ptbvlfCMfG78vaICND
KW+JcB1+yPoDvRtnp6qs7QL5I666M/h6dfY7j8tkMlE4IZ5DmbVQdeoHwgi4QlettXx673LFOUA7
/W+0paebnEe8lmQ+PSTlaF5hloeK7bUMjleEEDJMsUAaktsMM761LlZ77A9kwXmfjgD/K3Z7wIVN
3aZhqaGTAJugPWZdct3uhPo0OJwgNNjeOq5A9IYoUbnqyW/K3Oec7MLW8+hiSkuiLv5VxSt6SQan
Dds8JjivXp1EhCiEV5Tjt3Bb1Yb1ZF3pnonzaxdewPcMwVInM2+P68T8blg9XKybzMP8R2Oz8Q9m
SDUf0H63vmS//EwNhPaNEwpHcUZNpWjkAMrC79xqUauotq3CyhSdVGXhQEE8P5poihn60X58iOpD
XbZoqZ8RPsFESnHY4jhjDRHQNmwqg7uWfReysRKSEtr3Z+4wuoRGLZlDwcTJY2hKJwuWgMJIBzyN
db2iTkvMK23+6r0fV7ytoTyLsMS86suPzvIGwaL7GnUytNp98h2KRkbdiP6YYFaBY4OM0qk/cxkw
qkm7DPg5ZACGSYIONQ3qAVhbHiFaX16/d7+dSrd2U9nOIn1W8FX8wD1pPim2LpokhM1hjNEfb5Oo
ZpHeblYJIviHdXXVsxpV81dhoJnoi8Og9BVEJQpz7FtlcdBWaRl7kZsGpjjVFu0vI204wd9w1Bha
kr9RedAbJyOIYBNhLcZK11+GXAyoytz1iDMideD/9X2pugrGWtNGhQEe4O7385QmmKyAnYLN+gfK
D/Lek6k+exlsmAiM+jsHhhbw4xcVSY/RstT/2+1aKtReUBn1Iz37HjLX6GzoVstEQel+RG1IU4k6
keIjFQ/RNli+OBapI1kkOW18MjSGTLNE72yTF1tThQOtXCynzUmO2AAuzzL4C/IN3KQvtg21LMNu
mW8EovQOZsAHlIgW3qQZLWfhI+zwLH4ms3Nnz0JNQvOq2eekHg/5dorpFaWI4cfvWPwZWUeQEPhi
OKsUXPSN0qaJ41fFHBJ9aKlY+4vi5s6sJvgluas3mKKAs2iO/O4KiP2W9aVCZtwo4Z9BI/9SQSHT
5Ft80ypTt3kEkXKPnLUCV3Hjs9mibr/rM2JxZcUzMC6HOg6DJATBtlQKLQiSGEAe+TnorD+Qisry
wH6CzZZH/1LDbZ/Rvlav5th+gSlZYOXjapyH17qOw5mp1ooV6eXKIwDSB51wLMJNhKwzftByEidZ
f4vvYDcyWBeFKbOT9XH6CM8sJIFngd0VHU+aErRKPqD+UrBN/e9bTQomG5o4PKixZjKDwRVO7NZB
KCoHJhFKd8j9l8OnFXHrHu6sNn5CYAhpQLbTgGRYQNAZY/UpAfWtAnJ8pwD+tV6FTU28jQBFISKu
1pFf88ikgLjhhHz7gJQa/y3sxY9QAf15+tQNWS/MShwiJhSGbhskQqNjm9XiaIECHxCzIEeh3xkr
hV0ABA5EmqVDrasNqzZy1ncLaSHLFtYMfhnF7v2EeutGonvE+zj/4UEe+UhY0mkcr/WnEcen8dph
XBxdIhCJLjxTP+bf721p09g14joUx51jndy15Df1dK4XWI4WYp4xe4c3HQrVkcXNJE7jvpBAikuQ
m+KaAKkpaFJFOGsKH/9SD+72ofKBg53khBJ3RQcCc26Gc0+tIvIgnwPKsJyOVeINGOhlWDAD3hQl
s0qAt4Y7UMWyE1pIP0KJ6fdf+oUwrfOfDutRLsiYvy5tFQ1FSOLtHRbXaYlwdisUtwv5n5q3DOou
+qmzsx1PHM398KH8FAOc9ZU03A9EKiUJf/DNAwstavDmSkUSsXsLAB6SqcbfMdcTXXXzo67O6Y9Q
ICFIOqigoxQZCqnlfLdNDjKNAmtVnonwTF5swh9etSKWoWDzumR59C619AxraDGyWZlf4I7tBcAT
vE01QZhvBz9rxxuNQS9Lx8R2jO0yGrh/v8Rj0RPTo3jDyttomg+wREV9tzoQ45o19UeS8DHWKVBu
GIKGaU44lYgYKASWNETv6BzLygM8CnKJ/ADQ5xonB2Oib+YDt7unbMy2g2JA6CcxmrkxcGp+RcYc
GRZqBliQu8wuCjm0bSEb6pWXhjyCXDD4fa9hX+TzwFA5GEpV2pGTOsoHNr49mEDVspUhef515Iqr
Kad+OnEKOUGXoKCjj3fyPQiy8YDMxFUMaSIvVGeAuZXNM3cjL2It8kLN1xsYpdHsmOh7LenGNQwe
wG3P049rai9hAkKKMz3EtyIo2qI/Hz0XCSs0r/aOIZEh1AVfjNSlaSUfvWVvFNwz7Q/veUOX22zK
NiSMwkGlm8WKd87oxQw2617HfyLdoN6tHUhQi1KFnO1SzVN7cPR21Or/pQi+Gtby7sbAa+LTxQmd
HT5R3UmG/Fhm6knVDfnAB4TS0hgiYQ75jLTCkkhWLl6caxaEex43RUJluW2P8nCHNKSgv9K8lhDO
7hG+b2OHiRuU6qsH2guw4vxpP4pPuY1tSt2bbDI7dGD4ZavJmCFZMWo8STozk/IWmAGCE/CiNDIi
jm8UGCEWRjbJv3Ibp3LVhM5oxD1t9MVFk48D5ssSz0ghXwC9jroHhnMJzdPUH6Lc7xVM898RuKPM
GookxYhQTN2O+MZeDwiFYRHcSKqHuBvWkRrSRqwGBJjQmJav646b6H1kgvkmqcnzypmxG0aC9nKX
XKVbD9jET6WKBJjpE4MxaZBvTaBUw8jL1qkLn2Sr804SJGKKlSMxOi6n63aoxEOFpwGBGZdwRfc7
z7NHpVAhnBLhCa81ScxCofDRGWTP8d9a/LJl9JgqPAl2yr/uZrtOG4SpLeMBqR18OzAoof0TH4sw
NY/cfzAKJjxMepKfYkIOQAxtiJ1T49gjvJo1hKWcANxbhUuretOmY4kGZMC+kdeXrI+hJAKsTfaD
rv9248rwtw3YB+uPzZY+/rQ4bPNRLcm/ngTP6xXKAKbRqLTTgk3YABEniywZjFCaFA2gTwfYcmEa
JzRUYUfq9ddXp++wrr/uGq+bjEPmsRr9eB/BVdxN7//whQBW3KCfzMljqnJTUjuciHUZoivHDzZk
j14Tf/frpwdQ5INt2J87YbFTgbLxnnWbgixbV66YAkB8GJmo1PLSkHDMNrb8FLevRG7YXqNu8mQQ
vfFkNtfKecsQjtPenYtyHBba/kcljotAv0M/VbErnQUTtoNLqhCXcRATSrtdIOcsVwyVKqwTgOWm
yNbzFg0zopwIxLyc8uF3kKbWNZ0EMGIqHZ33Qi0WZ8YRQ5MJsfmanIHAAAmP4BE57/3V1QJGvbqy
TPoaQ2jbAsRUhPCNHGCtPBPiR381F1JolSoNN8OtrbAiLykgui/g7yocsMs/D5UL4ZkB7LkQ8nWZ
s0DlncHGVEYHQH8hYsswTG/z14i+acDsrokpIZd0S70CQMDN2GaaiDkV25ew9tm8ROFMHqvmnDCS
5dceBOQqgfk4ArNsy0Ank8qCyY6JpBySShr9cgoAGt35B/6DH2mG7WnLu5KX7jCq2Gxy2jDqz6fP
+334IjhfTbw/lhYt5UrblR9E9A13sI3kZpqQ3JSDn1XSjkxa/L1D8dcue4kmEsBhKMLiV7cYHAXu
9ht06qTs6Oo+XbuApBa2PTgf0BUFmrgxrLvGYE+iT1V7pn5y4nISWqkUay2Vb63zXBUdPsRy0Uvs
X6rXhxHe/rxD92fUw7c280oBXfargsxJVqSWAf1KRaave+VTetOsDlbf1LzKqWiX7tSEMPJJiE0U
FK6t3C8iXBn3RkgNJlGvzpIfLbsyhOOmxodGOFxtJt1QMJ4lchn0/IGPaKX9S8LXEG4cvsKbaBbT
f6Yd2bkrF/gHbW+NhEvCw06ZGvbWIABK8adbHkQPlTk/xaeYGOcvDm8n16QdbdCNTx4pj3K+GdmM
EilNfrJFYOP0Dm5srkDPzhPgZZk41B3i647iE2/PBeuxcMstEQ0DubPiP/uSngNc8BNUlgehSXWs
5U3CPeHueEKlmG8KzKBBRMB2lWbRAD/Q0VXocLt0Yi+IDpqrV+O2svhnhGp3Tno/xzkg+H6SFDV8
qzmoY814RIQvEwHOFvKO6reD7eZZhXk+1wZ+qee96rjaSJKTwiu1hKnPTyCAqvYqhfVuu3eLRa6M
dIMe4Nlg26qEtf8GVxAdZvEjKSNXEpGQwTCKsA/LKvZOBg/Xmys2e98hj8q1wJCqpBKAxGs1Tt28
YfsGDhNfPoEublqYpoDUpW2HZ2TIzw5zq1M97Hil7UM17dgvHp4DW36RVtR9NCQvxLn6Wd1xsCfa
BxtJ1i1iJTUeLp98f/yF+N912/Mlwqi+TyDMpdYqkEANhJNngxoLUMd6GJsW7hfQkovKlkBZW3VP
or+YGdovjbIEoJHo0rRqSo59EynbUq949GOnIZg4yS4weEoCBlno7o7bkg2rwOSk9RYgUIEJA2aB
kDlZjyUfOAqkdJnUqzadWmiqySneRvCVOQtJnxCRFWUa+5S1rCH8KQu5/l9PQFpmtKnlnxU9NAkd
RKC7PhycDb2X79TyUNZxYodHbAzUyVE4NLaXeqT4WuBHkNuTo9dTW/LElOhAsfTqurIVvMJFPb7/
uepULXEq9Clsq+Ysas5A/tiHdLubJGErkMKMbNwf19a2UL4/EZWJGhcSLYCAQxfa2ijI5u3UQcOl
ypls57hEFSc8XlUAeQ6h8j0AjKhzbs0ub7uilUvwKu4cEDp270cwjd8Z7p70wwBlI8AjgRpYSsEP
WrA4wHdaABvcQxd6rWqqmriPQePnrYSDNEP2vCGyMvXELK9nVOE0aa2DmZP54VtHA8jpyxtSsMLj
fQWXtWcAUt6v+DbgAGRZX9YIkSzoY2rmx4XP3jmvwQblXYWgIAMgGSHclA8gI2YtH2KPUd8d6h+O
w7/Sg6qpVVt6/Cylp5JpbJBTQLWnfrlV4rk5wzAiVHUM/nG6RwttUhvA78KDoFsdIJVLedo7WncU
2alo1KusbkyFOYCztpjX36CoeKqeSK3Bbrc/dTDva4RkByaS7HBPq2P/EOfHt3SFn7LIP7E7rV4X
yKZ9uncBQ1FHgbQ9zRbvqABgrC+vRnS3LAhZznkEmOXvY76IaY+bB5+L4pb5xi0rIju7KbCiuM6C
GzZznvvv+A1moccK3VvUCVOHV6uL34WKtMFfoMaBsFLW+To8GSf0oFft7U9dd1WFcThukLWu5QxI
eql/vUdSy2P3F67zVZDXtMeDStIyGiRBHPSJTOQ0ZbIiDRxxNPXsqcPLeq3FNGDND2tyh1QyirfE
NUMbkWOKs6mqdYjeSXFnM6va0HJ4jnZ4lFeI25X2Vyy9AUIytAfVNyTeIoKdeR8yEwKr95epRWoV
4sVxECBFVm92SfCnR/1qaGW6+uZyCqfmI1PnyyC+5X05OH7o/zgRRjkyaxxu/o748/R8dB1hvjfp
kCrRFd3g9/kQmNpx/MxZ36iq+h8pwUGAOz2dwAWfBZlU64nkSGQBXFvGIYB11v5qx/HRPPKygt8V
DmHpmFOVmapbv5TEP6bzp7v5/68RSZddOOnMwcc3AfKUtarFr7FtmsEWg2fkWNsYmk8uuBFqqVRA
IRPXtr0Uda3tSA8pZmam8xEUW5ovX0SvArrj9cHX6kP5T8QRnFHuusLjKfYohxNg0XbwhDj5f5r6
7Nb/BCgqIwEnsO5i4Dzu25sxjbGppnXTHDeisaIWrQjcVZWZ5mWLaCWz7R+McnSbmKlDcELyr9c2
IZaSa1m3G6mVnLf4W85R2zVMenUI4JwUwTcE9NXr3Di+O97shIJXO5i/LjykCshtGbwST2yFle3T
O2OwcASkd+7XXvJVqxVQAgt7CFfqJPdkRISKebrDjQpPernMVuDho6qaD3yi7YDNgTPYpuaZWQ+V
u/JxUp5/nygC0RWjuGOCq51hSv9e6ang2MzBMM1cm8XqW4ZHWqcNrLjfkHhMDtTZqWXqD8IQ7rHp
4ZH+Yn3UnvWNOO/lEuqNCXGQOlRDqACDIKD3ryga4fyRjQ3ZkXIXAPJcL8lCC7Eb/h++smXxWTDB
JSKHFH7aiULYVppFChK8mRmr3jQhnzB/Os9UP59g9w/wUbJliv+e68QSgagXOFw0nQ727Fe9v0EF
bb+TV3voWKG+GQ4ShYtBRUPSwl+SYitw4lZfzvQzEIWYVhsJqNJLmSh0FuG+V/ct/KNke84mIttv
E8uaqa5Tjb8SULcTcRjig74VgJjD/pndvJNlAPuYKGjRj120xv/VnsM3s6LrIqgE5HESU44WmiL/
Nr0DrweYro9pzIIYHiAvqAQ6N/DQxWNqXFaDkp3QwRRzBDQx3L9SAYAtdKga8se50TCBalSNy8eJ
acGZ6D+trISrjQjuYfuo4U4EGOS5LpdjKshMPXDZrdI50eLKWkdch8FGP65gEyvDgpJsYGwDu94N
IqmJPeNoNLyu9WRSE2HboiTpt+TyMJgiuexHPoBBXs5WR6s3q5ub5mDOaZtsYkM9xiGFE6/Dquna
/wuMbIQoCvJX6916HkCTd2jJxmxSYwAyCx4FnWyOvtdj2HTqP296EkwRJwRCFFkItxycyWI+YlfT
bo8sWq0BdQp9NDya1xSz5XMtmezS/SgTHioEGDNyunhw/NLUPoyHlb/O1wNrYKrooQoE7FCT5El3
8C6ufLhSk9eWLh/atSFaDEzFbGMRZFbgDxMHFKSfEGqlm9t2VK0HTy23LNT5UnzZ/rPVDGMfNewk
mf79l63+wbn3NAsd8vMfvtZVQjPBsr9VOqEohnSLTzZc5pL29TYoXFHrU1FLaRRHk0FEMVVc2DmO
BKZe5rH7JvtTA4GK3lkPXkK9d5f7VHZRr9e+WtC7j3Fqi/EUzp8ENd7eUrQmf8nMlgkzkDzenage
da2jXVLhqvCX17L417cZKyonzT/c9Nv/9Kjpqarw/09ej9nI9cioE38VILBAYS70dvio9R8tFJm+
wsxY5TTU+NnhrlPkiCMGE7ZfHTvFkFtNRzy5Ek0b1HsIm5PWqHZtF13xg0RoePOoc3IRIAlWmkun
dYPG1XUOrEWuIrIcQXh5Q2NB8C8+Gwqf3ZY4/hw7jQEkZvB3kcOZkhFKkEwtR1TNs6F0agQiGJpP
Xy6xkmWTLvgU82uv8d697UD4clOY8O3jdds+bmP1nQS8CG+COETOg/tTF1B8jCGGa9O6Wu49mNv2
ot5HFRuRZIlCjhv+oVaniOvje1IbQj2LF5YXWl0prf7dACRMMGMJDnR1OR0U+v5gZwl3RSPn+sEy
PvQw/rk5updrtT+KymMyf+/jG5shuuXM6oSMwKIysbDzxLZ+qRLhuO9IPE5O43ZA7X9U39BlZn2G
kPv17YRTrN9tcHuHr7mLQF8v/dGWSWhWn+BpU5YrJ7EnfHrQa4cStt3MDttj/PE9spTXiBmrLYpn
YCeUDbv2e7ROz49t7ZoAYts2swxqRrD/B58WzerssC9AHYHY54sy6KHnktYWPfQ6WN6lQGbEReYn
tqoP9n+CVN3Q6nP+imQBgdxu8Zm9ujjn99dFrSm3r1+agkdDeZfY8nOKvtfpyRR0fdm0hMlLK9s/
Q8pcwyvFAA88nHVl9eO2inD5cvLeRv8nxVJnDOkp9VytpeEab5uvYu365k/v5ZgFH7bbA8R/fnoA
kEpNpgJprjO25kd69DYccijdtlUH6zZhy67Zl27kqBbWri8jcPeWFRTVOq/NDjrgTx5OqScyV7lO
69mzcLNTb0c5Ysq/5wYZP/qAKoiHo9Ch1SYmgWbfXQi7KfaJCArk3TZzMKnuoCgmIkRLkC5l/vqy
DwAV8wq0NTjVUxb7x5J+gnHUuaQdWf3opCS9D1imbRqjP2/evfR2Ix/+chZ/H6EdrATaSTIjclry
XXvcn5uR/vmbgy4FXDeqsb5UJrrqggRnmAR3KbgeC/cXl/Ck0ezFNtsAqt8YLzd5WAq+zI/PRpDW
UfriuCQTcRTxr3zVlkuJqf2O3Pgo/GXsecu7jj6C+hqLRRX/lhEs9OyyqPdOEYf+VTRS9FOdNiF9
v/GqOadtJiTNHEiGTmHbOIRHOFJxKQKzImmm1OXjH9wDxrHqD3rrAmPe0CuBFYauuLtZ3fVXy6FQ
aElJd4a3K9u5bCO2DKfp3bOxbt2IfI3+0sIHKB9CCgxReolCPUgdfhX/kwiLkYbJPjdw1a0Hq6Cf
r0BrxXKZhKeyg7ZKfvOfeT3Zo09wdnvqOskyq3Rn+K0oGoxHK++g9YvPHZbT0AgU5fLZ7rsAAZEx
JqOWmOG3EM38pBOLXjOO4dg9DhPI8QhOhBbCT1qMe04YTeKQfUx/60eXxw7O4FaUqES1eyVEDzPi
ISHLDGT8jkgvd9B6vWmWum4d4LkAVrAQaC2DsNNGb3PhiwzSfPBsDQP1wy9LboTzp4YIESx3kvBa
hQhKD4VcA85231Go12SvWIGKGcxFJ183yARCYz03bqCorIaqDQgX8FAjdE9lS9iRj/HB3x3paM/q
CxJbfSPyusGQPGrCzD0R1ZZnFaf2GgJ2L8WL+6H0Pr38jm6SdM9CxmJ60vR5lZQs/cd+uGzRLkkX
W11LgFOPH1KOa4eTu7ZNUJLjEFks+G/lGAxVAlKsvUg4vEMVZuqoX0Ynifs22B45T1cOuVVKj++c
mxFT2dmfjXnO5AoR4Aoip9KeFYknWSE3QZEskPP/pqG1z2HCLyIFU/tvDAZPQcVcPM8WwzNfZ9S4
LWKRSjRs/rU2aa1gxPTnH0VckfV2ZlhNEXaUdtH5YwqkREDEJaBT7tUjTy5rZGMgCXNQOivzByJ1
mLH+RPVdD2wxHAgKTD6hd8cuA0yXZ0OXT20AQihoWPy2+vrqz4PWdT798MI6mn2AoZkhhYHS9SDB
7teqAv1uVrqIp+nq/brJn54Or5hG7QQ7J847JEu+LuNJqD3pYf3IzUofk7uMeiHlLVbvuBQaAuyB
5h0NoRgP5eVnqS+or0zVEjYSUIzvUUVJqIr9EMwL8vGGmruJ+5b1+gqzR3G8Bh/+02ucUP61OdET
kftvmf2ngEs8kAdvw71H1sW3yHZmUJG3GdtN+qJ9eZr6KyfZrQim3pBOHJcIphCi9qAA95yekKwu
FyC9urQiBLVetDLpxmSwT5nhZOH7+i/soxw5bI4RVEtR2+bNAO5rVlM8h40V9QthKw57GgyoGI98
YVDGlxE1Ww6DjzcQfMZSPdBnoks/2/jheXdBdJ+kCjzfm3WFM8OWP3UEIgkzVlbxG7pfOBfwm+Gz
ubxpwZpZs6/L3r/j+CoANC+PazcjYNK8G17X/O2LWipDLYyP42Csmq7aVZMwv1emv8PQlm+OVY9E
yB+To6WkEUc8YGgoFPRojoiqU5jzjRUQbTjaqi2hS1s4pL7aIcHsw9X/r4v/pqf1inhiVHFvcwIV
HYX/XIDvZMiafzJHxzb4zDzjVPiYoVm48JhWNApo21qM2aUpfCkSHXnPXx5SMY5KKZq/tKbEkpG6
yHsXQKJiu5YJfTVBfT3N6CyRolsqHff8pF0RtLcU6ikhzSlXDZic17JZit1Co4NpJUMBRPQXiy0o
fOmw7dg1JcTNB8U42JtvFXLmNDLOGSvkC1joouTKnRUenjwy4yMyDRbidCwoufrVXvNmrQlU/Xw2
OOiNxt8qiQqN2HOXfhTiAv2MIR8mcwyiEa+v1DTQvuAYgR0DMd3vV5gJ1pilR+fnwhN1jisNGb9n
1Rc0+e61EZ86ZTsxQCbTULdnL0QyU2m3sC23RfyY/4Y/qzLUhc99ehKeF3rLj95FZshj1Ax8ZZEx
XxmLm3sj4XQ303qBfMAFCtteA0hLSJOdqFIvGK7HQPwrZu02oLiRUH/JKQsWEK/igfTi5S1o6Nqz
1IA6kxO3/A5ZFTiz5qrJ9Q4SdhhxQ/EaYazsqbO9OIYoza0pwBdXNehrFExe/u9WdeOfiNFZFN8P
ZVf0mS3b2DynnM+ZzK2wObUuzBaeH7kgcH3o/yuuvm+E+85nHpk+fpoNSyzJ4EV/J49O6UXteuW3
+IKy96di6OkVQ5KWE5YrhiZuv/cKG6C4r5kPhsbVIA1k/BE1wF3QTkKGvU4zKyqsEfZYkn6EYDiN
O3VbnvUP5lcmiF94+/nhhQUSMVXVDDMTZoPuV/BqywX3ss0xIngKQUuzgMFQ21AfUcEp4qaZFP8K
Td9BM9V3tk4ZcNozH8b8G1veEaPx/Hu6/mDy1zAMQGqzFBWwYowdhQ57F9uakbhLF0AP4Ee7enHf
bQPJzbN6EmpuvjDdqieDnlqYi4bLyggEqznwIAnMdV2qrQhyed7nprAthDj2sFWejIEVEafTgsCR
TQFVwn87ykxsKujOndJ0HcCzHfBy6zotYzYL90gN1XwXu2INY5tOcsMfhoLhx0/OAJnkFNmQwoRJ
v4pdFHVNq8Rs+Y8m1ROkA+zC4AvMCkLVZKeTdWpbbaRGQBBSdZWUj38PO20JqD/O9APNo3k6GbLV
5Iok4NRcCASiAfSaNsC3oV3tLsAH4fyE+mJ7l/UJpnk9Pw2ZVlV19BkbSKT8kfzcMDtwFhm8G9GA
fC/AzpOulgY4F4JabuWi3H58IY1s3OegX7d4PkXmKwul/BfJ54tCitBa0L5okrONp3fMsW6qTbSm
l/a1uwcen9NSVmdXxLTqyB1wKHwm5UQZmUmJy2mObvY/O46HdaCs5RX12JEhXhz3hg1QVw3pWCAA
OG4dRWg8bJop86OJN3LtdsBiua8Yzu2RZEFHWf3tcrs2sFDkrjKYc42u1CYmKOk0JhwzTAsYL12/
Mk0mQ0opTRepsMWCYWkQL0R5Q1wszS7tvtrWKhUNQ2+Ztu7QSoggFLxFNbwySI/chYl5HLuXpreE
qqjlsPNES/84o7iLTMYu/IDkSkiO8pCkEchPa21fio0fpTpjWvzKIsNtTfYg3qVlqK0U4dI3M/Dr
SAroaIJmjyIexA9TfxzyF2xURNdgBD+WVE3WQXW3Be5G4IBb1Ihc9ig3V3er7+lQNSpqxpCveuk/
xyVN/mNkHPFbOnKw+YP1V0vimkrYE25B0YDqPZ6Ve2tDVKrCNa1NS5MVLoxBSyXk88/xAxuroNQ4
A94uX06OPQgMDbYDd/W2p9ATdjwl14nO+TcywVsMMcpI/JtRbKxBuMvYltpCTX6VxOGwWeJwxD7h
YpoA99Bzs/GAFqZV2na15agsG3dMN80zM8KDU4uyFRevvkVEp1aZ/v6ZScrZFnfW5ceBMnWrLrXt
q+PNinApwvRJsCMAXJl4LJc1bA0i1OAISAx7HRdT/U6IUnwE+HCJKYT+jna1HtejpJEmEQjvEgt6
nxgIHL00xP+HA8HlWT8lzf9guh0ZRi1JfeMBmtxLTBci7hMg3VqVufIDKqG4mEGmyvt4AdSww2K3
oHIV6jAup2b4yLDwmzIDGv87fcphiBkQqtthz5saG7UeKNEwQpP+niujmlG3KuibJpbL3ofJPE5H
ipu9Tkq2XhDzzF+2WjlNeTBw/Rb+JxQHpWxirWvBBSVktSyL14b5GaAVAmIRd1Akve21UJMx6SRo
Uezj9vpPtwmEqxYznzzdtmmargQ55Ud/OOiQ6lxSM3nGG4S1ikbazkHI4IkccUQgRf0wJQHJVpKU
dEHz2MeHivxWpkWLsplc0sVdZdWqtwAbQrbFsrHM3ep35v13k0sl22VqC6ZCJ0JffAfoE88Su7ve
JrFlgDLkvtMrIBoEvOWe/Po3aOsWFqG8TDCmMkQRu5gbtkngp9UAZsKScOQ/9tKYEzB6POb1ESz8
inKyVt3Y/tuoL4SmYZ+1c7/R2iP5LrQOoro1Kru/fYMv8YNQ6MAPGptC8rNxlDM7hnZAVYzODFpD
YEL3+LsDGMzCNGJe+8rQhpxD2hgcieObUHbZ4GuW+Lf51jVRzxDavIDTW55szKiYTI+SpLJTyJnK
XEl3A+Vy/pleGZsvg20x6mUg5bCYYqtkM6QfFhr3gTJqdKPEI8mYYsBXfO12WB0Dakv0j6g39vSH
9JQx5e5cfrkA6bjZEya1udFbNU5/nc2/FuZI37oYe2ekFq++wzUwky1PX4RdwrElu2J0Eot3EYYb
JzrFT0XM8WA7Cv+/v9/5VX2hX4gqa3YsRotYdcdrr4uQe8q/aKpKLGGUEg2nAwgQCzQobkjm98xO
0MRQElFJWEQC5g3KWZnRiPZ5WtW2a1rlJOGdRLNITc2LdRHZs+7J+LsLnFqedBUiRLJ1ot7xig7U
h9qDpoUfzPa6v9QjbyYcDCLZsNk7dYpFaQaDWoz2Rp9BYF0ZlMZT6QpgbP2GPzGzXFhj5lmq/ODE
olI+dhhVurVmOCG8a+1on2NpOi2DEpVl5nRtTvIyC+25dHHtpFPr7QWp3Mpbtz9b+p3thK+Z099w
wNQWEaFukp7+38E70PyEfztFZ27BG653k90a+wanFFBepSywrKnW7Z4woo/BMbAl6PaNxE+jvgC8
RXg5HHLaaWG3LYKRkxbETe4D4RqX3eqK1UM6YDVxVX8ijkNsQQm3Tfa8kC5v5aOYXZtl3Hs+PMsG
PeFXi8wCysv98jvDrIqdD+47MH3xRwMznH95oxcnb90lfPv3wam5yDUEdbXoEekoJ9T6VmVhNkPJ
3tRttg/sqgpILFa/5U7vqpwf1OnUgnWxCHga5R/eQ311qo/w7haK3rfZOJhpAY5/ii1U98Lq0vT8
9FrcHdni3NaccpPw0B2RxWlQBSXDOUifD7x/QKsaw0x26fwoRoEA6cWQoSBrpnFujVQBwxmGyJgd
Gde9KisuObgfawp18rx+yfedu6w6tCW7fA9FRKGlILdEL1cSZRd01/M35zOgwo0A5I1PHcWS4+aT
fWN6mlHx5WltvYXbOtyLIw+9EOx1YSA4rxYXl/ac3pdPiMI2FFD3hLb8MY34KDR1K44lFIEa3AMz
84m8ZhIkhRVcw6RTM0fn3W6hLjh/Z9rPkXaYODPXm4jtlBBiVNTe9ulCLoWGZzqQY9+IwlR4cjsF
Fp/awL5Rz6v0e96MY5bLQXQD+1jL0zHgkHq9GTFbpQXkXRV/yrZUlgInKxTOaoquuO3vv1QJtY4L
hvpkaoRZPUEDZ540jF28b8GWtAuEn+r0xy2hp7WACPZW0S4qnQGbRFSQQpN6oK5bzX8jI7rWt5nV
28iWFKB/pCKWZC+wUuf+M3AjRlF20ceWPiBPB0UMcrJTGmAnSSJO7kujzxyNaB00wK0+AN7DlVn2
8upGANf2HC0oQd7R8PL3Epmfx9HwnXtDMWm+2FukwNj+giZqImLnrXrqChcDSKeSTV2RAFvDoICF
KCAXvdexNGeKbDKNTPkKZ1dcz3n4QS6De0a5DplbKknjzxX2QubTDRAaAUrkHwwEnHEmI46iOXUQ
HqTI/nJZEobMYtZ0x+iT02m/H68FAEp31AwB7+ty+do8fxunE33x+ksAb/aCJiotMY+sXh9B7gX4
XeTwBi0Kjajl0bGqRMl8Ff7ysn3Ujp38Ayqzs4dFMGhdKCGz6jbOpdJ0zApk+uCMUZPvwVFnWDPo
uH0RYI7Udp2WN3SeOs2BMKJUxcJLIpnHJutL8R4AFVtRn2iWIbQgaCNZKnS48UaAerRWksn4IyZc
pK6NhiZNcjhcFAco8nzfXBEyEO5g/OXf4b1Qh/JXxt6erwK8CKMJyJmrHpW2oXzDMj0p5lyDEmuQ
++AUaPfiXvAVbklX1DVKgadrPwm8NLNyZVrx9FasmXrDtN3rALqweaZqUwoWjMxqh4xRgGSYUe8C
ScVeYYs+8J5uFgpEmMjdLkIcTmqitfuxTMG8o1cqOWjMDg/Qxz8123rfE1oDvEwVIxVFRgHyI/nG
xaH5k/16k8rDG6iPn3j3q0rn2no/Q63cmK3IflKp999V9uTrCAze1ftHvYaWt4+pgrVFJ+um5xqw
Foy+n0bwauqkNLeXteekTrzo84ZqyLb0uyHpaTjiRCgEdSfupC1ybn8RBHtARYp+1dIt9CQElPIV
nilvPAwa6UW4tS9ggYZr6+7PsItyUG+qCGeyO49fmbucm53W/XArafA5Z+A86SGDuINv6HLM8iKY
XqMp686p7ZeZI4TvozOn5Fv8WBP+IOgBrJFBwtGYiMMr1xv0HAYeHHXbAdWQSt2n90UYlb2pPy1k
Mc1GoG2+QE6DH8pCdWEEXHvSNevdPhDhxs4K7tjAPM1in0eeaKiQeXhkJx2tGArWj+rgY7YBO3pN
4BLyQrMxDNZI5E/esn1O1DZhaYyyDavtr2Y9w5D8pcJyMfUc9yK/rfSNSqRHSqKkqk/zW6KjjeCE
MzyWdIWO1yPIwX24eaho64UpkLTMIRTpkscsOlk531hGaPFD0ZHaLIbU3sJlylC2pK4+Gmy975EX
MNBpMUE9WYzlHstpyQybCYq9WPuZHluQIRc5mrOaP5AFmDWKJ7qPBJvy0yVqtrjID9Ba9gsrJpdP
GsLBit34+TJIqfRqw+Iqk+nwlu/xLeWktDzVaV9siyTeXLtVWOaP7Xf1HbfMkOttlA/sfYSMNaE+
cUBusvz7we9VYQGmKx7L9CKY2Iv3yq0lxASAeQy60o88IiAzMB4fXjn4pi0ptzTqrLk21DLx/6xE
5Z/lqW7azPHbco3bEVozTyBgAGzGsaXA+VcpI5lHJNYeFb9t6e82eurYOogvRWlt/dfVexPO6Vbo
gJoI06VhD5muos53sNeUdIBWQMBNmEX3vHrj+OZm0gmvPpy8xoH6RghO7Pqu0SilXk+1JFnZ1D9T
Ph1nEsrmlqUhyPa+hBVQUXCiFGJ05GtAoNspex3cqhSBtPtiA5qYpJ5HGuXrjcO8hINb+NsG/c9E
TsNA1EnAPFyO6ySLiJbHwVn2LCslLUUxcZ+ydEO1xK5jHdLfeGA7LK8f8ViXnitmWTQyUqDZmcuu
iSdI1gOVzBORdqCVf6hb9XDAy5SM6TK8dYcauRFxtMnFFIc0iwOmEgW690AqaSpnZmNMvsF6VRfU
wir2YH/61hU5wAYkSmPcc03fOmafJmHByXB9W+5my2GStAwkbSNy/1QJfExVc5J3KJRGbtvsOkIj
v/8QLJmO3R5MTgqAR2vM2TKDsVtON5lToOEljmDnt8c17vxJMOwWZT2Ded1e8/vhdTd6tf/hmXeF
/r8Eq+1xUSKQYgUG1mDz7+gEPspG+BUSjpEYEGDH1vqE5aCjdQb2NkiBF1HRhZzA8UIM+L/1/lWL
ZUU2NGu0VSjgC+ek2or7DdQtxY9WnZxtEZ7c4tpMqlcm3yrXM9gY4+407X5o+PW4dyVzlpHB6X6V
j23KaMnW2wI+HfQg7MevaqSxahIjN5Ks3u27a0LT6FRB/WEG2Azm45LP8qbT+N/R1FPkkLM03hbd
Hbc36biZxJEGXI0F1jkWqkmlH3hwDDDIo6WszIexCYuEd+FnLTR28qp6aSPXmNNu4jbsxUcgyAwK
q5/TyDD6wv8FHwddw/BSyvyt/dffBoCWRgapti8yZOe+I141UgkpkeCs8Qymp+/+3kGydM59Ro3E
95fkTA9kpLh0VqxwAZ1d8sV4HlMhv46esU7L/t7RIkGzbtIfhY0THO5NQ38PEaEmQyBkFXzvniAV
XyahLT+pGjKlSFIFDhhey0rOGjYGPPGXxJQhOLXYBpD/da1WdNxAoSl6xyoD7yTGmASIBfIdp+/4
367CHmoRKqIV3LIw6MSUhSubwxZjvp3Eid03mIuMLMVEe+slN7IrHcYExckHyUe+27sP4XTEWKcw
UKaaim2QCf0sNCOFH26GNKUKTSZmdS8eee3VK40W8pWlGK3WV5qA9dL7uznVBdG8RWs12SBQas0D
jJYct7DW0Y0Gqg/B4FhQhnMyJNXWuYG3izpbZ43EhBLd5m25gvp4ARLawuMfmTM4jZkwRXbweBDI
DMqwUJ2iij50HMkFeY76fiuaayboMicbickQdA5SFaKaaHLjmuF6emkhIZkL/99djX8jJa5en2xg
CoVmsaz7GTYk9g4ZTzRO/RuHtBEOaQsJpw03DPTfnrUA8PzxE5VEzRnS01aKNqDYDvHqQY2+QQ4V
v3woVPkOpTFYt09wM8WMvvC2beZlum3C+1Z2A5tkH7S/CvTHuBmgL3DGUvxtsiAzKFzeZN5k9M/G
bXLrX+J5wyIrMNT0BmWbMdbr76I0DVoiM/9apa0xicBkmReHZK3NCXSRUi3n9M3voXFzPo2uG21z
YdnQIT8TyDfXSZ5vmvSUqE2pklB6UBqfoAAAqAwbz/Ny2FUm3iw+tRY+1mtm4cz6fuqJaAfXkmD2
8/XjDD8PUY9oXALbMSbGdcsewdiaEJ2F9zm5QAlkH/5vHRywg5hMFEvZV2gMMobhjWN5z0Lbz+Jk
p1aKpzWPQacHo6ihj17L8g1zIBp3ZeCDXxLi9/ay/Wd0OvmJnUQp98xlwjnXGcX+T9jSsUXgmr3P
1A0Ge1WqKiO2d7WqP4G1Bc0jkeAPV46Osjjly57Gj8Td9YXCkpKcuICakcWj6a4SZLLyme4fO0+z
qykYL5aLgTwS57us7UbrJ8Slquw5ysrIReiIrOz1ozlXXfhwYgSZOS0hqVBU264sJkAEN3Qn7ZPd
xX89TH2OSV+uABPui3dc8Y7jiNRilQNRivk3quqHvOEJs322HiHW44wHrqGg4ZvomLPuouOKWdiG
HJHQf98eIPrD+ksHoWyZO9RM98EaAahg+a/9icbeHwefkBB2fGZrCl1f1WvHgCsJIdnvGP26D3Ng
1DGQAUPyZZfvAi7NlO1ba0jHWImAQtZPFEh+3cOL6XaWPS4nRFNtocwiLhPPMySbYApyMBBCN0+O
RaDZGVqY4+4YocdSigva6NY0QaXNMYNGlwRfzUAYSjvbF0Iq/ia9iPNUaIcqXdP8KccdRM2zPLRk
2bR0hQc7NStQTosEu+k0Drmm0TpKYYjOvwQ81ev0JrAlK65zuMjfT61iD6eyIOLC4fQr5CqpxFga
xD0qSIuHQWusHX3xFUKld4e8WYLqbXxAuhZe3nRQTbaICyjXlSXz4+AwCKzZc1QXH0WDRn8/iGu0
enLuzYrhFvLp+gf3Mi9jaVLoFYq8aA+P+jFQUicatdvrRxZcVhfPpiFve8WNldiXuqtBSp5ttT7b
fw+sewCbP6NigNfkTjKr6Yn7KSzuw3q2gTsBHVb6pzC6AjpQM9wCZEsUvEpKCxALV99iGvNykufS
AvMhFIqUVl3LQv2oeZtRcDxKiKPTFwPfSUBCd6qVM5R0287NAk1gbS2rlS4GdkFex/WDm1kbR9ju
69UeVT59QIl9PzYpfPD/vURBAxikr3F9V6PSLnsxuXt9Th2wjWUZ2MfBqkIs2AEsX0TycHqJcAG6
cPjjfrKzccX9T/+qkWTQ6+1tAHJWM5fq+3d04rKq02SkboXN7cGLRmL6pqjcn0qR3DhU7K+100ss
NSE831VHl8vRXn322FomN+67gizUEYSL3M60eYBdWa7tc503+CDwyxZfc7XNc5tV5ui09YMtaWQE
pqjcx8AL25sSBrcWw7N3RamkKDfDtqEs09tqOYgaa3xeF99PeyAmT9A8SFrqkmFtPdIKLc/RAOpr
VKMkXPeDft6EdBaRcEXgoIxvvZcNyR0eY/WSiActBCAsTC60KM+8172IkkYkLnHFlVLZkIeG5tG+
Up8cwGsQ2GlHAUjEJig6XYqbq9AcHCXvI5Sc0om2mRQgvpnRDe8sWUBls0BnaeoWoJDVF5/kqbe7
GLQ0Nban6+eDYoEq6b/r3UuDvoow7uWdDqPwbWhFPeS6CsYYSU4/9wE7ikj0zXvbs2GSr/AMeCqM
hhScEls50/nyrQIyac1aQNw8Wy2IMez7sCMplhjY7CBcSsRSu3mAhgbXUTXxoxxZCipK9Gcpc1bi
1ABChR8HfDcphklF7muxmLSJYshu062tm6EJSCX7c49U4JAixMHJ5i3PInmMC85zWvDg/10Im/g2
a2UWzPUuw1dYuTnk6GasFuRX8FEzMm69UQA8TPLEcABxdi2ce7UxOz/S6z1ITFgOqMU40J3Zoxv4
qG64/abVM/304TM6cmddPrbI0tTz6ODVDRWjk+iDWbCpQjUwf8S7b+nSf06QhtZGhuHAno3rxOWw
PGzAT/+IDu7SAix1B1H4cQ7VbAbx+TysRmNvnBA0ymZ54QJInWak32gXHX1PTAIoSrkvSxpD/HdJ
6pZ9buRWVxmEqC5QfGTMOV6HRvyzh7dQy2ONg+gL1RqCGZHq/DzrAuUPoK2yhSlNfLViFRy+WfdR
Ipy4xWw8BUFJKB60z/K1FYPv1IPGxb80XPjQ2k8tgA+V9l7GzaiUWVO/W7ruZizgyJaPirf1MZZm
Cv25dvMw/EL+yCH5TcG4p0aOReRIHQk9K8q5+aYyNwZuGaETx/WQ67kPegLe4gC59G5mYctHFD8p
hbrQ2Men14/47UZKasWUEJ7iVpMkf/bBKeRQqU/e3JLA1GNRWjMFViua039SzMgRS5Nh6sfrMEOd
ypfEEt+X1zM5mwvM0zZ+zvvFCUcp253bfLwxJkoGAAHYUL08qg6PZB1+yYiHI2F87zQQ63+IgWgj
Zb5q2BMPdBitVDUc5c7FtwkwdLTXMDmFSwCgvaAJo1HBoOwek/vaz1fS/Zak+OzZiuBdqwR02yxM
fE0vjYHBrbkc3a8chg3ge6J6HGluMAXge8h44zi7w47NIJmaZTY2qjAJFjtZPYAsnpBujAabZkVV
HEw8M36pZueI2mdkoCqzD2CQ4XzvWU7JgRm4x79kfkn2SC3uxZQ5NT1lKdNxPCJqIIxirS8FIqQ7
vROMYyq30Dus+Cn51lC0/h4TiNMDDBPQI1DalXPwsJJdpg5UfDLiXZKg7fN5s1oWbyUSlvvkoYGM
BOhHoDDLgwTnC+BWcRjnEkijiPkys6pGzdZxL6ddIZ+4xjV2exiogdX+uBDMtTU/YnUdrrN9rsbc
HFXMfeewQq9Ne9ufSax1HwoMB5J6SlBQkiH4QI5WCJcbcAOQIGm3yh7I6AHvX/Dtmtj8m3ijux3T
uDL18qadtQ87SsCs40DgxPH8tbAAKOiafv4PGTGu1zQPY3wrw0rrOL5GtGI107e+VAeyjdnp/ITE
gGqpG1RsANMaClxIGaGQNycE+PDzIyVXTU841rlTYocYtmku6cbhqX7ctU9COqXjBaOoiJ1hHj8D
V0mNp3yEh5H4pqkY4BssCaTesmSm61TACDcRuYZGJBGzNAelX1V35KSBJ8aO7Z+MUrEigf/1t7Y0
VluAf9Dk9dEs6InX7XZp2DUl8JsqundAmC4FsRyQU3O5TpDse3DMds1sXBsCcwHFEw1g5vorIWc4
6DP/oh8YtgdCk5VKXK591aKxviA+THonydtOUkutgOwq2v+yf8Gk1xB8ptXUHJC/hTJF7vucux8c
QbVEpJBPEREvW9ZxzYW53V9FrmQffMHZCwgROFS1HDlEXod8fjzFt8BmPF8qyFrE/UkyFifTaFj4
ALvCwBYTecZ+9ILHytlHkYwrMASY6gAfHDi2pbTrQ792NWsuXaDJpAS+ufvGMLx6S0bwYkJAyAeL
PfiIopKNdFVRR/j1x892HrihScX0bA35NrS7msELFY/bmwKGIU5EwzmThlxU9uc8ztsYp5Lca1Zl
Tp/yvIdPFEo5H4ww5rYyP9PK5XrX3Ut6XmK3kP/ZTwDZFwjjwl1wRFFDKqn0Ad0b9tNuUR5hwbJF
IJs38yywRyfMskkhwRWDnPwyM2eHAzWSvhj7yu6Bfs1YjXGwgQ1QSurpr3DB8dV2kO1aN/TRGN+F
Rvwcy3f3BHVNPDb2Znus8nxry72rm54Ld0DDaReruXXVoT1mj6jGGv3snv1qXtQfgNkpdiRRQfXj
wA92fYfv6vLEz0YxNZkEt4BIvk5eJTouPwvK3GpwGZVSiZmFI+/Q4uKHYiUkOjk8Cn2v8G3AHkkh
TktfxWvGL8W/H6EPhkHOumazra7NXxhWSKmbaULQd8qvPJwe1wa5l6Yu5+Fco9Of2HVIesSACRIA
p1i+tBxQSzBXXoEQ3q1uQQzRWott0U9hsGJ5L1qpbbQJ6Qr9X1+B0XYDMzsyE8fxSrQbUd4EgFSO
iqCcmHMPz+hkil3BFRkvnHNkWDtcCTcnBWgFgUqCjziquZ5Jg8mIdLSziJEjDydcuvFEY3Sx2Q0Q
ch8xCmTSSRCMj1dR9t+d9QVCzjvdSeP2VpvCv0dLVRe/3NrwbdfTVllNRjFaExRrBqlz/sLCs9Qd
ZPCsfxoR/U7hsSyqVKF1tGzkA0d2Uo7FSn4K5GZVIa/f5GrCzwFhIzOQd42pXCKaf+oOsH5KssJ3
b5TUA89+tMzjWsh9KtKBUVeYij9hvrgRFW/s/oShKoUVnTYCRV7E8BOpWA1NZEIsgbcX+tKzCUNc
tUFNsOHqn4x3RTW+aKu79+WurJlzsyEY571sAwdXcuhFH4j9H2xnCNOpnoPLtWKM10cjHxuYb+Sq
0etGxzBRpy5mv/FqLOMJ6hGYjVMoc6xTjpxBIkSdwdeSdwxluThZAV4gKVMOzVLktM1BRnPusWnz
OH8rZ46qvrFWCxV3w/lKc5XsyeeHPBwxtWjOQj8Q9VViVz/PuWraAbJ9pJWVOKp4XrMQkCUAOyj8
dfTrM+4G2bJcArgZJAU0j0AYRDIgIZ577V8E6XJpBNghNyj6NDX7CP1YLjURz6FVLKusS2ngAzji
IOc4Uv4+AfawFlUUcFf6jkyNSeGmypn+d2M66o26iQBtNqBWf07FByFF2E0bVbSV3u0o9HA8xWcj
0nFirXB8B6K02kQZijdit57fDBX0X3Y7LkvRhRKwfYB0xHPf9MvGczHqN/DE8dWBFEsFEVetXn7l
PrXB44un9PMSxcJMMZZX/Yz1CzWGl78oZEkiIYMMeWBLqEBAVlikaFJVuz7CPjToojW7QHege4OO
SwGICZgJxpQ7RScZlaiveDmNRrXCvXxTJMhjf3lquTFwGo/nrPxmGpzq6FyrdG2T+ADwu8gKf0+e
z6tlt/5kx8cYNcVVkyRJjOM2Pzb1rtmdaMWtaplMnmVOhvpZJivZiGzuFKCnvKIlBEpFTxm+/EE9
lKcIEUPIuK5YB2ynkX1dEhSdWRoZuBwzuvsVa3PFYFnBKBi894QAsDpNV2oFWFhqbc2umb93k62l
I2nVEzEcWOxAF+sXbEASYOcKPQnpAaMspkTfcnBE0xWS8kF+0N/0iw/4B6P2Z12uYVfxTvRHVAFN
ujyOrDbV6ZS57aoliBPf/tx9VuoYkPgB6XmSbZ/QHWXIzxkLQaKg0uHWmN8gCa2Aj7qEYVyBscT0
ORHRFXQrL44x7BYq2Bbv7zvPj/dz45XDxne+P4iISbickgSSCvObsNdAx9xP5Mnfgw/Oh1Q+gEbX
rKnkfbO9YzpEDhOzNKTGDYNroPhcRCeZnsAEVODD8ELvUbF97Wz+17ODBGT6bDiVSwhlT0WcMK7L
gH4k8I2WtZ+vF4XARCcfbyAX6vPR00u6ivypM4SxBAhslhigRO8RNpBMYOPoPTKq61N3NNa/gmEZ
/e5eqXqwiD42DzBJkLyKkcpcr6oMOqUWSS5L+UZJv/kazH8fuZSQ+MUTDy13xNktshGmC6mFCcSJ
J2SwvbigHmj7mRRO8KvTA2Zn355H1sqWqU2zmEuVKmfU0I3UVpswJJG+T//oJ1xtzYLObSPVXKUi
/FHpLvDix6W2MFqgDLi9RCud7TRG931yH+1NTjGKamGdXdgPIMiCMADLgyR5YqQ/8meU19ryB+td
b91mrkDSqus9Qu9P1nWHifyci+bw1oFlNcnW2uDSYyxC58dAhO6JaPsqeVUUm/ISu/lVzYItel/2
mR5qpQb1COzewHhMrHD2QpFBDFdo5xMZM3DxwRCVSlE7/wg+z1KijpRZR5U06FvOWJ1Fl+qFd75q
p1XNExLAXY1MojL0KKCYgrCLAXqBFCXm29koYCsbayrIZulBzRRQeKb+6O88LgRrXc5r5yvr/fya
Qa03uKaFZPXnSeR9Zk8gzZ0YnlXpFSVDcmhjhFmzPHJPxuum753tiKTIuMW8R/3WCGGltrPD1pWt
PsXEUZ7NABxyZv82nQM+hIMjO5tKTwJeBWVeYYTa9iNpkl59rpcgw1X2VlOf+VbxUXOZW2Xn6Lhf
SxGeLoWUaAjdD3eazKnTmEnIH6Wzgj3+Gvi0TFX0i0+T7fcGHFQ7YzaHzuB0oeny84LbTUW2Y8NW
PlB7x/rAXzaDbuYHgbSWe8XBKnGdTs4RBvYodz9CxRomzqYIMJbUV3zVmvboF5uGhB0ibrqkPU8m
snHHOzQjpQWnXhU3b6mBLc1XgfRP+RGHTwSzyHGraNvgN6koTUuTQl/xR5AMS+eMxkt+qwKyQIcp
t0l62PXVoWajJg8rT9ObANExFOE1yBC43Faej8d8lJR37z//XfmxHhGtGJgVKT4VG4Xrr5JV3Aeq
UnfqHcHWi+g4OLf/1uZXg8bhmVDOMo6jGCL+mqnemqmWSpRH3QN4DeMnUgScBfmkiLozyO96NwMQ
LRrv8u/H7MhnMb4stFCReDa+WC6g9pprpThn+hG66SQRs3mp1Qkw9piLYsvt0tP6eKaCMWHz44Zc
zFZmkaZ/Qlx5q3FkZSVjfic2a9R7ICcgTr/S1PulhkwogG5qVJccZIMlj9ZCXSEZ56/TjfoeerBg
ozpsy6mT2l1ivseAIUibAvyqRGR5Ne1MGKoTEmPkgJaqU4i40KSYiemol4gL9LeifNv6i+SLas3e
dWXYrGZ+egpRn1BGMl1uX9cEdCG3dXk2fsC74Q7qbpZaEkARtK85R3CQnnzAdXp3XHkItbWRfO24
KtgZFj9ytTJrgHvKiekzvaRQ2S8W+XF+ButWCi/616E3O7AuAtzwqKYLOJAG/SfvmvURf6U85wYO
p+Z2cdRnSrHcKXaXKAdvsVsuBQiFALS2fAGTaBWNTp9dUS/P4v1Dq4Uyc4HHRe9d13ncLZZ07bwV
97zreoz4Hbr1/ongyp+KVBQajOADUf9WdmHZnbkHsIPk6BqwJo1urxGac7Mb3I4i3rd2frq0yFKo
hl5VMvognsVAnwezlTz67Dw0ucLYkFeypwHM8+WH/YFRWndm/ZBMsbfHUXmUWNy30WeE11aXvcRb
KDu02ey+bU63DJM4mAxZsS6WiIODfYGMbsQ4iY5AgpMqYEUuhRiN7IvkccAo5J8hdwZd7Io0AZJG
tul+QWg8LP8al6Wc4S09zc2VN9YBnaaWYjhjSBESZ+DTq9sH+fd0A5dvb9RbpZHkGZ6iFCrgU2vb
lW1g3jzdMx0ethn+wqe2KOockDGWdCPaUPRf1IgPu7bmHLbxHqBJ3PeLFjXKNNu4VzWidhJqKuUB
U8tEes9W1vY1lcmAl7Et3ZHExDmCQTPgunPAIfx7gKQPcaf1t7tOzeefZLJsSlqQhTA5y6QkvRHd
pGvngmXTZtQM/62t4qvqjqogrK/0dfHeqlsYvVE/p7KVIPI9iTBucekuZY8E1RASPk0Vzz//ep5A
/X7LfTZmUxqToeUxqTyXuSDTPJoeaHrnlZ7iMDuqBp7XJLPYS5izIPybu5h4gxSFRsc+L1mDf9/x
wj1xEhq7zQOHQAgNjUZwot1Ur6aLrR1Mp8T6S9BYyVH7JiLL1NZcbaMYgD6wcFKq2FmsjCyOniDG
78LTs70j1GJtPxJeXpVkMCuSw2j8aUFCeGib5bf8zdf2YtmoDB9/zkSFtVo/tvP3EIOSm8IKZ02T
hx9i4wDWg9SDb1HFn0dnEqBb2B+jtODr1omDULiDz/up4HexTEi1D9EySfxGEaoUv8RAWzkw0rxO
ZgcUVrfPZgQtG7WXslMmPiqlh+Yeqb7nDQLzYKb/DgP1aOSKpf5WJxLJhiEF4Sr8XvHrtimQScEx
szl4WvSgjc9RCv+QLqY6DeSLxvd9e75SAuiXyB1RV0qV/YbaXkjHpO4+OkksCYumqhjxJez2lDN5
4c4D6oTzaHKrQHYKPIwisa3GgbboTLj1tRXIn08/1atsVjZ95KYam2vpTS+WkhhCE6MG0Od8v851
1x+jlEmBECz777t2ZqqXT1MtsHLVtdO1vGTY0wlY5aa15oR7rdjzxDImo1WRhmmBZ5k+6dVcLieX
gFQL4CbuRTGvVA6ccyD/LYZ28u92Q1c0mGR3G2C0zDHForNJJD2zKc06EmZ9vvCz/f4YUtgaax77
Pfs3Ah1l8VdtGsr0zxkuwyUg7E+QFaULbuPOSrFclMSOQDt0hJQFBH6hZQIQMgHGR94465M3Z1Px
eloLWqHoHf2TIXYDSljWe4LpQVSD5tZ63Md4DnnGkU4AzjY8siJO2TFdTtNUCAQ+QKW8W7Dm/iyu
EUGx+XaaNGLpcrVoKdh4K40kLtj+xbFIi9tm80Z8Ll7Ggu/9YQYNbACY89EsmARx7/uGzphsc1So
LViNug0e3yKxq9dYHgSFCdTiNqeR6wvMrO8bZmcSBx6zVtnVrdEskDHzXu1ERhmz10+aZgVkcgWJ
5OIOaWV69oELjRynyH3yCeMldz7xIbuNFpwqtn1cN1Vf6MazkspM6IEnRVLIBX5V2JNgBYTPFCgy
9GTUOrhb8bVCx6ctH1dCUM+Mnt2Sup4rrJ0t4vakSN/KpQwLFRO0lh4Qi3Cu3VY+vpxBIssRzLJV
UgI0a8I2NZTvZIaQqrHq0+h0g5RwmmTBDcUfKVCxDzg405bCVcMJ/8I+MGMqYNa6Hyn+5j4iKitf
d7N8/4TdY5quqkpHeQ0s6bAupWG3GyIXQQ56R8/RxAdXdrFVEjb6sjvAVeMgqelUN2Do+eQd9exF
ogHDTE/dChXJDihZjQfalcSIqb9vlbsySLvOrKfO8XoPF4cjPfZl1KFSaZ2R0UJhkA21IXqx5RqX
jTsDyfwdICR2NKMCE0A9hLJHHZL59dWYP6CQKQQH3wWv0x/IVEgVBUoFNTYctTa8G2p3ln31iB1y
nBnvBTiQsVRPHjQhWcjqZKNpOSEaVWoru09bqRjWiTjpkLLpyAVAQGiVDV1dS7TS32o4u9Vd04Bn
GbBacEQqQcbUGYN7N9HlBIHCy0BeWa4vBrOopLyd2zOmSQA8W+cOz7ZqNkmCEWXKiyoZZTPrQWKF
u3yhTQKRYwW59hBDjh/n7f6jUnyB8usvcq7oN7+Z9v6IevrH8xaibTYHyWVs8iglvdLNYpwNltol
Zq8yEoIE+triTaG6nqIcGnBWbSxwYaTexxNpohepfoc69kXkwaWR9Sxy2N2mmxh0p/1EG+873cLs
Eh3WXWWb6P6hDSlKY60i+TPdMyDcJjvJ7EyZPBYs0E+h9bZczrAkH6Oigd4TRkHsBUBVNsIoncTt
yZf+38ltZf0N8SfLCXCRrEhAZtJ2manL+3Zu2Zb3aL97pnO5sjW+q+ZuyQk5Ihcj8JbZ+E/SVeuT
gTewlqJjx6u19vTcIbSifJmgGs54vB37QaMHlVWpuIMH/t7k19htnwyBb056tKrHYJ5Rr35iC+f3
SkC8fz5AYr4c4ybj6TTIk15g6mz0cL5HQ8qZu8IjGb1UKotydT9tfB7JOGzcGMCs89+evscHrXeS
Ode1NMJxQk7a+NAU89CBoIWUpFfu3al7QHhf7HYf7ao6VcPVj65bOFjpaLYnlGQEOB9seQNdhDX/
3OjFOZE4j5sGX4cAVLGf3qPMCs23QIVM2UqJnxGZZLMFFQLxiI1zfozUVLtjplT2sdKK/RAhNahC
B+bocG4RZ2l4WS66SXn/hWXHGOnBQfyEgWNbAT4APJlPXJUD3qbBM8dPS+JXmGBNJr4JAIwC4Ygd
25n+QIb+TnkpNVzRBQaRoXJpw8B8SMOP+S814ue9bG1QyInulM5jQisUBtDxOCwyt+FkarRVbOLS
9AuGnMYTQTLCcPfdynlqbK/JUpcaYq/LUBwm27Ry3hDrVwSRixoKEmWJxu4qHsvHAcjz2qP6an7v
Y+jaR6FyYKSBaCjT/Ir4Pt4ZqlUlYw9DyXhHBzWGvydT1kcymYYf6LrEbztIKqoYPprJ0AN/C6ap
du9u/tPy/G903ThZCXV+yZd71SKYUE6KfVfod31Rikyxu3e1ayrbsaXAxMPPqBAUBfMx1pcOMQph
Gd2aPBo1PqbSLRBjEWqkVAzbC+8AYzz8G86qgCqNqOOEBKm8k0vwZvO+cZRl4uo89cSMb+DqjQHc
zPX+BwbZw0bgFBfJwMBsCNCebbpboFMlitqtVP0Splm6+LuuJlzgKFor27ZOEatXP/J18wPUp0Op
GM4axuMtphDnLleOZzLusOrZRZpnU0/MvpDSYZIdXL0YWeg2Dy0RDnEuZ0yKEnVTDGEEL8PriIlc
lURNYFDfMH9RDh0jPFkr+MCc36TUeWEEttcBL74UW7Kw1LJ5crfTLxa4iQoYt9/1MtfIABEPmp47
5sOQx9w5SimNvu0y0/VJNSaqaqSwUa3YV9Yr2Ko6vxQXoO9q9qLqBtxLRzFzSCc4C8VOJFeU6yvF
iGrb94oBXuuDxNsu3u4hfZF1rg2Or1qqdCSbfidXKaR+JlVjdFBaBFBXUCecXaS27QNWO/yDJxbD
2dHK79QHI+5/a8SX6sm9oNK2FBB7XGjQnrYwznXGxff0KRsAC9YmtgyKFd1v/nUdaxH9wU8cBXYX
QAPrgwXG8pO0J7BCZEgMjfUcrJEdu+Ft4LE5Xby4/iRrBTXRl8F1tzY5wBOkKfMiZKQhrHxh9c0E
p+Tlhz/+5ccpczRwMVg/lqGOSNTITXLWIVO+mefm/Nmog6BQ2wdRsuSr7wWpWVGEYaFIjB0A2ueR
WJH6HFhl3sZaVx3AG4I+Ni71FXuoprDsHk1BOtdC7Oel4o3fr/aFFwAyLdDJwevXHp1V/biU+aLQ
VgafgXgL3OJzER3fnzZvM0nrHVT5sAiwzuhL4/AGpz+tctMENEDiO9IOVsbAHzRVZ1o/CwHeTBat
GfTbHbgY0qOrrXBeEH2Ogb/iwFv9bWVPjEqXdHGsUVMnHJNQL/eNYfVzvKWID4p5SEo9mwodlyZg
2qKYSgSpFWnAqva3gECLw6BAccIxhy6pl+Z40SZCx3xoAy5Xl2CTgqplSXcVFSTi4G44U+6eUHTC
2j5x+FavrWXrSMkg3c7bNF3trqn3g57UEt5XKjBXMPecE58clFiWQ7VwKx+DUZ1hj+4KAIZF6RD+
yOrWV1kTb7mgf0kS/gYyOQUtXCy/DELLMBxVchKkTz1Tq2gfNkNsk6ucSS0ieDZyIRznXNUC7mlV
EhEgzOGpKdArkltKvBDA0wtLeVwUfj3WQLc4bvEusbcpnOXGBseNlS4wDuDteJwZ/53fNgRbB7yB
hIQdcGLlcGm7Q6oJy+ogWmotHYuU1+l104znXDfqSRkKFID5Yvp3J+DTxAZVpQ/v4Stcy9b6Xn1B
L6ruK3hz2vfA/qD3T0t6UIYJrFuwY6DOi7EdYjGy+9LT2enoaOXiRoISSgQyt7PsEl00Ccsa9WyL
ExU0JFBxVKDFGZJSrYc2l1Byn1qDBUBAzIqXEwt+u9C6s8vspJl01GRdGlVvYSgu5TbDwNWDfQN0
DjjRdwF6IW8krnQG1R6sfZt0gxKVIasZZGzbnEgxd+YL0THOtbkv9Tc4e+F0DWSSWUF270UZgLuh
0yNVb9mSGexKC7QRVYwWfbHmmZFFD3zem5l98jrhH8wXe5wbmNmlNm29tc8Ak7KkRnmUhXs86Q23
RhhzzInA87bA2i3DAc6XFCJjxCKWVZCjKEuaX/omMk2AD0KPvoYKg/BIBsduialV1FP2BeYMuFkO
0F82Sj6e4dAYVe6DdM353jxN8VHL4tlb7PZEXQQ/xClQ1hU6ZR2dCchewFcaaajGW8kyqvDuTeNA
sW8aA3syyxTi88sqteOKGR9lZzjN9TB/iwdbma9jsBauSCJP6qSvxSmOwHBW7TjqqdBjKCXvXv+h
6Zzp6DofiGTfBSFeXx1YKI2xGFnx1IMgv4fu/Ff9+BYvgueekHkXLkgLVOYsVm3SPQQ7/ZRVChuG
ZLSJMO6gVQjkQfQ3s9RMD6SxkcQLb1gvtn4cuBw2jN0mnw5mO7ABbxqScaHjA0JSClw/TsU5WOpE
rCmJ5SfCyE+JAKICUP1y/rL9uwIBLdm52vsZFGdkz129xHryt4x0oFos4/UQ/Il9SZU0nPNz2M2E
Nb+hNa7xINF61in4VOjfFYKz3niFSYHLA/dZ2uGY6XcElBa7Ub9Ghq6ijnEzW5eZV8a23UixDC5c
NJMQMvMQsc5L1GzCqyvj4UHggnePiTPyYQ7Qb/3VMs6E5qLJoXjIHScztAPHyJTdZV49aDYGkCm2
21j0mRyViWikt8sRKGoGqRPaaQ1tRutyvOa7sEIk1TUvx4EkP+A4Y8NFAjB0FqCSP5zfHQRSR3yG
QRe3sJd7YBO/1i7Bwweo74NoUNrlW/rk0Spwg8BDUO8Rcu+zfXgMxJBrNdT37j8n1gpVo8N2KkRa
sE+I5cxV/z10bnYkw40wUUosuOXt+kzJQVumkv27SLTnmozK0xQjwkxzvrkWRemp3EaJO0qpp4CZ
+G1hdpuTQsfgLQcTjI+CUJ7FF5pS854dxJ4vsg6JDDUeOJI2PfqMcptsTwITUMI0hd0oYdiPo1lo
TBV+c9qQdFcM9e9hfi3K2aWXnzu+pWdzcv8NqXx6fA6sv0fKfB2reXaxjR99ixswQwomiCdcgMp9
orEgN6vQgUw+KIrRiwY6axlOWvhw811pfjMeqhSCB8dhGapEEy/2MLJ3Epw3Ptwhy6mCR3G8hKoS
1PRHZAGLINUPQx2HWPk0m34HRA5w3mf+Wl4R3LCjTx4yN0/G2Sxnhgz6AV+Aj7h5skADrvaF/ojl
LZdV3Glc0Oydz4Gx8fjeRAeoL4CWB9VK8BEtGLPevQ1CWCcyjYZNw25HBUlrMF34ncJ0MxqBIoX2
pAsMBTeIyzABNCl+2KiGoArN4YgcFZgUdZsv6GiZyjBKg/sejmOfWyprSFvDKPDhV8Fw1ERBxCds
fUne5LHJJc+3TIO/hoXEEWEIQFp37H5Kn+uR8l6wtCk6NN1BtzakRx6qM3/Y5dDWmjpzqf3Dd/bE
2oy7+5mDPwVp0fdgBI3vCvlvVTQvOSmmPMGwP2tjZrmPfFTFJTRVdU9kEx2eXl5J8YIe6intgNcm
Q2IBYzrM26M7Q2pWaV5yctJDjPPVqqQ6EkMg/2nhqrdKnjs4eQzdGWYTQMH4rlu/xaZ00lyOfdnn
yAFMKy45ukUNZhkvuG2CcmO9ZQY+XXcXiKStgkv/M5FJi3qy6cCUfZwfXy9AOX1wvlKT8ZsO9+k7
tjfIoH6+4e9R2PzyHpONr0J18KdiOJ6NfM0EeTbtgS5UskhdZ0ka/qc4VXIdYPvcJyN8wNcKRdKC
fbh2G5WejFEgz2SNoqjYvxHK4a2SDvMISs+X4p1uwpZqtLXNSJ4VXHp7c+gNtnPhzuL74G5N2uco
Kzce2tMsY7zQ+gV9UaIZMAEUTW1B9ofLTnYmlT4SoiqwO4lXPDCVkp09AXEdV70Qi1XgcaN2UZon
0FMpeGOuHBH61g5x8OANOEYwgq7JRBauTpo774EzwncqwODNdiWK2T9sMVHbk5XNGStV1Ii/2cai
gYRj98NRyBn7Z/pn+MmZMCMYXPYVX+qp1RyqiqOSn166YMeSs5+h5RJyuMk/qeE718zgLHc8szCm
EelquvoxUTw2oEhfzlC70tst2iZJ9xUjnLCuai5UqPBnEdr3MRGRX33rNkhtgs/1FHgwHRASKOSP
FZiUtpHVeyaaUpCfxwTuIuFYRXI55nSZPqAQyY/dmOsiZ9lidrEUX7LXV7emlrdlMiyg63HzzLLR
Oq2nFIDYAzbuDP/grqHYw7xJQFgayNBV7696qy8YQunJJxRQs63w7Ibdh0gwuhzE6BmlRHMLIfqB
7+kn2vVHCNWRh8th9bVNeviDLBcnh3BmM9PtCRlPstUj6SaKNhLFs2eM/rLKsDIo9UJ5B3Y0pBqD
osLf056VK+o9/mz7Y9NrxnMT7m9Yqt8Uec4ePTUyv87pED4sBuNr5alM7pQCtsN6bqdeRujvKeFv
O6TvUcWJVq/EZpxeRJinND7vFezUaG/oe+tyqRFifxNBYTQDfTKi9JfN5l2jEJkT7jfQXg1AnDPq
qCu0fawcpALJTV/fjwFWoXwZPWE1v1tXH1QSQI6t6hSU1W68LyG908JkPCV8yYqXoC33GGau6qKx
YnI4JC6xGmH30Yu83yqR//DsGRZmJPMM2iEfyA7do0Bn37vaG6rNXtCLPrLG4LcA4rBgBeiBJhwm
CdIp9mcrXms4E5Nl8j6NmIxezb23s55M5BVZyQOheZBahcyvqJW6WlAEb3O8+r+my1GxZQHbe3Xe
Jyqg1HGPTnWRGrBBsuyBInIsPdQoTat8dERz95xZ/DM0Edv22wbG5dbGGQ9EKGit7BtxjiWudGIZ
7fDu/KJIr5Lt0xQpPExJR1Rq0yYu9VbaD7QOD2mwD/89emjlQUaRM+zmt3f2RdUYzoo5Y/EcSkvD
QrQKL4OVkdWYK4rw4mET+2ayn7kOSy+uWkzvUiU+VXehGA2jRFkwWSkDmxcbZQLkbINnkyD53lXo
x93dvkHsZiss528cGmsUywDfsWKEJn6Wx+D4sWWHTODAP6FSVhKPmrFYd00qIlkux42LzdrlyveT
zqzUyE6GxQZNSPDxm32BvHpUiq7sQkgocAGGf3U15Nl41Zd1OG/YZscJMCHU1rTY19l5GnWcZ/BQ
h6B0wsqhYFvsnJAeTn7d4DzantMZbV3JOqwmAwftkWZllq8hpcFSCNAn4TlKbqJ4ZyQVmb9SavWL
vaDL3rjyXQu3R2Wt7+jQrL4Limi+A0FetvLpw/gMAKHXnV+8wp9QGy9tk6soL8kx+WgPeTDlVVir
rc0CKBrMawyaZFgkF3wtKhAwGV9LY91bHGSid3HVinhDxp+Gq5xPAIEGoeJWTYoBW7aIqq6kDSE3
1Sajb8G256o8HcSDd/wA+KyH9jQjfstFKWc0YJFtmhmHgic4GfiL50z7ZAe9Cg5/lysbV8dfUDAj
4adP0YubfFgSbcgmaJEELhVUYFpDNQEdeqHt0CTAvGGtGTNc5CJ3geMSdcWzF2RqceC3SIBYoMQ2
5mRvEh5eC6FThwR0fBoyf3JQ5+szQD3jlAWhX6LwY9/Eds7kICrHCSq7VSqn9PPMddQfom1fkKU+
xXOHDJ+wPLFtDOOW6zpvDeVqyQ1THGbWe+b0LPnP8d2y8dQcVCB5leVYbxe94ZBZ5LAVi1ZcmdKc
BODPDYxpkGWozHonyj8o9qyddZI6bhldqTNotvfw8FTJJCMNLM+kJXeEUczgQeLgHRHb/Y3PpTxh
T/hm7uzZ81kE77RsVr3xB2y49pVDRoQr+VwcsA1OXlNpYyiY6q4Ylx3jBhrw08G2FHje6EnPjThA
96A/nNLvMtuuSnmRJgTnQxHWM2cbIhObfJqlp1a4CbVnnYm3xtrkJlezLQrx2hbEnN7M/NR5BspI
KTmxZ55EXTXbT4K23oImotxuuOGWHbpDGqx2eKo7ABK/LyoSV7kJJwnOtFhDZ1J+DA/Xm2q2Pn0j
RrIKu174sIY4dDA6vozvE344YBolp/osphVeO+5PAu4cEAesbGzTX/OT/UXeKGQMvgMc5glB47ci
3v7NDAl70lRLgThyJOyMHhkkpWsTsB/bxYQWUaTW6BLefzkRB1YeOgfJNyjr1d03LBEG7v60qNhh
dT+xrKmc8X/fcT6x2oYInGWO6iJ7rDVBF+rK8Im5gwrgggLI44EcwpBpAoUmQriLzEm7jX9hUDNG
PAoTekeyHTql9jjXy+RpWoIfnUl7t7R5DQUVcPcg081Jhp8vA9CZh4xkkaZ+BkzbGd11s10MAJVn
rBuRR1mnkh+7HU6pElM1F1m3yDk6mTcHX9q5l5dZjb4Zm+zPO1Z/P1+fDgfPelp6ZZqKm7CbdfQI
uIdIW3d2lkcN8I+SiUcxkChO92gy6xITzS76rujdFvdLDA7nNL2d0isOWZACtqgK9G3BRIDe5LrX
dYHuFbqFXLdYLvOkIzMPaLT/BUg5i5Rnz9t0UeCTqaVh3OqYI8ye0zWqMVDUie3EpaUH19lvgjMw
41C7NORpQyvZOYuLCFIDDHbcWecUw5p1OZYj/ifLQmfWm1ZWq8tvljfAK4SN17V0hP3GwI6VQWmR
PLSFpcKxGBoRv+vGRU8FUIqGEoVrtPcl0jhNFqCP1gsnjfplPD+rBG3QfGp8DKJBxQ0ldhuqQTcv
zauELkFx8LTPucqfrGUpVHUlKywbyd1Bkfa0WBDujFY8ynmSoB7NI0rpJw4fDRY1sz3gWuyzUiMJ
v5Fv/vY3Ayri2QqKPNAEhHLKJASDS6s1FTSBmBphuECjjIiB5+U9dp2NJi4KvFLS5QfhN14bj9/b
UnkR+a//x28Ft57pe9qL2sk4iiIgDEbyGEshhgqvcoCFrJO+noPyB/LRiKSX1oPKiaFWecJAhv42
AmIelzb2ClKeWFEbTZBy1UfdI/fgXnSz0IYr3mjICwO6wAPzGfO2oOk1lmdWWy3KXaOxSzEL0ULb
cSNy91mM0SE/Jxn799OznEUC+MUtfCEhb6iPYC9D2PsloVri+89/Ckm8VJcQfgZXuhfC7WUcDOs+
HmvHkHSGbpKtxWcYZsx8Xz6IvGN50g6hH+rGo4v13U9MYIZQAKrc484vDz/fAF2YHShbWGOpqnkZ
jjZxbkRwO36n3oQ25gm9dJDs1GdizVLIbL8MpIRc3TyxnXd5zQQsmqVVIJDiqXSrK+dgNBiFVO1E
EiwU2ohzbXeZpOgeRqZQxuvl5VmfV95ocQM0VSFU0dBIB0XpiwUVzs/YNxmIWMoQ9xZxJ+Hl6AIr
OOAKfTDgi3cQO+4bY/JC3g+vaplTgO1IlCGV8d8PR7qO+FzD1zzl3TqjS/6AUTjib7CZwPXlne15
OV1omY0lVO9oVbir6JW47DF24Kqw1EeOLlGeHQOOzsc+jfKcGJPJI1BrJ6tSLrfQjTRONyMkuIZE
cFuJxjPfQDZutpE1/NzoZY3HTz1uZM8q85p9XWDbSoj7y607pQtCgvRzFYchHdt81a8HgrqxmaVy
IVHIkCPnIcWjiNZydeDRNycBG1HJbt+SaTaZT5elDWjZPd4ZNMFqehr/nOtg1zSigjbhlho7bpS4
usqvYXyXMh1pvFalJXtaO91s2H9g6b64nzL0E2G3e+BXqbFMGhex3JGaBO0N0s5tLs/V/SAeyDMz
4rne7XuslFyQsBiMJAyyZHnNIYgLKcjDxflUkRhaTulmaHYjzfsdMw+TSH/KWnaUlWEvRqjZm/gI
cSOI2NztIsxtE3pFrGBlaNNaLQCi1ifq9SPB5JBJiX254b32DMbvZ7SOY3T82ys3zV+/S7nuMwhP
VTTe8IoNJEPr9AhrT/FsFPDaMhcPpk941GXOUDuDJE2sT+CH70z3thxOwglviIq5dt6G5Kxw0A2p
w1X10EgSrg7TEPqiFp+1lGmY1d69h1n3k5PHI09lhrp+ooRPhKNd+OcC2NZ+AerGf7Mzn52m9ZrJ
PviX1jZDP7OA4sVsJTiWKhtb+ZDKnPEx7vwlNOpI9CLtg+FKclgP779R39xK4APcX5PZ4pRb1APF
aB4/xgJvTGUB+iWJji5VsVCDY/UpkJQpdyZLw6COfX0vee5YVgJfdxglJAremGVPFDWJTToTrWKv
cMXBb8bNeQ/F7EzzG+y1xOOeqPcBTnUcIq8lLRC1Q5qxQ0YX9sDTUupmDZAVwdLaPKAAfmEMAN7H
tlxYCs1eieVfLlr7rrMaqfbcT0hyBgRHqapRmZ7DLXg1RR80wxeQlKuMEFvsheunbNoCd2XiKe9L
/MLz9uPYY8zC0wC9AxlN6/fLLbdu29BfgZYBglbfBP7pQ2x9EaGoe0xoGO/ovffp9/mLIER/LZDQ
ICzHfKb4Vka92ov9fKiaPnwHK9liyPMFVbOBF4EU2iF5IGJKixGl3HXJOT/0eImUB2pps9bqgMKX
ajShOVWCUPhPYfu/CQUASUwOkwgrbxxiRlxtGfE+2LbljnbqCVqxiTFeorM9jtHU8aq82IqkCqYI
r+xNo6p/XiGH0exX/f7/JQ+jMAPO5s+v/ZSErb4IUMkSGr7snTosU3Q6O4v8WUap1xZG5EfXfJad
BjnjttQKzaMMzYSjLywSCwMBxWjbW/lbRSlaAoqVtZ6g0O8FmBYioLPAnzEHza0LmegFMdtkcMGz
hmne6J3XZCUjKD4rRLSem3HeYwwKkUz2R9Z+upwZAYKJOpmRiIltpBHdvgfMHuZXRlyoYFkGvoPO
uYefILij5NtoX/THg+HHT9bbGG4zcR7l1ztTxud0xOsmLbMH4VrhQp3Fi/66zvTwQB+63E519C9V
XHxxXwFWuVI2Vl3QRRxuo2Jhv3hr3sTPdNJboJg60iS7geChq4VUKjJTJyXHFky5eHzist3SBRVD
KSEpzBx+Xl+KU2woGjFZ4QBhUZsX+CQsAdfS586TcnFSaNh2YsUhG3+kdFl7m4YgR4WCEgzhpYRU
DEwHRW8z3ChVUR8PP0/4Eam2KXXZYnjqLtNPMPMlmUYpr3xAhl0s0AQSDvG0fNThUu2BQEt6DVLc
+o83QwDea8gyP2/HlynH1b8tpG5/ORNYDHAX9l4a0NkBRyIZJm0+FB6/ZAP4b8HxbZpW1NDMzNy6
1Y71K3PPgicgwhPHTBoIUV2eJlwtqyko1XT4LKdsgHD3Z4s/OpKaTdjLjGbtt1esXTorvbv06sqQ
HPdDg6IHOIityZSb3bxUoP7jyv5pX+Uh+agm+1lcVaAYm181Ya4+7CTEIk8oObYRjTDf5SWrwZPh
lxe62LCr4/w9g2jPaAngiBEmk4X7HUgGRFLfcqz3NoGluDfqhTyOFlEOY/ZHsbv0pZJZ7FopchlC
0XM9hAMuAcFIvPJoJ0uGXvgpjYe6ycu6R88LUH+zReqq1VzFwOd1FXcufSE7TBQm5f0UEI5ZWnQL
o9zsjlo2ixtwu4tO0F4neOYnpFFR7nimD7K+0fzatSjgR5pzmID2L38lhJxkbCR+d3l90cQ9iBqP
v93mm6e8jEm6JfrYOMEfWJ43HxCNmXv+/g9x5AM3PJx0yDfpkDfk1Rj2lPZx4piOo/nMBxHFysEt
2D5jCXPMs9BaRrF7DKn2cH9GnX5UFhmZV0TQK1pv4QmCzTmei3WrDRLoZkNqDldXR2On5hCn5JEc
tR+FC2oPSVAzepQt2Po4f3ZTsEp8POV0EMEBzqw/Ft62YxmblIdIpHCKCujIgzykrnzxnHTpM39Q
Fz+JaA++dbvcdRDcuC1nh1JlZd/G5IqY9hrj6Y37M4f5Me7BE4E46W+yI9AsL4N6OK8AxLmNrTV9
MkLRp5XSnMLIXWv7iRV0hle/k5ScDdmoxfGN8EoeJ2jGB4AAQNjHdRGRSg6OJDaQGuU/0wPXBdLc
AicoZtKb2YEhKOcr2EQHWu5GR0jM1La0HJLbBH8INBEEisU/GuroOzidQhoxS9aDlx7l4sQFOGHT
6J27PniM4b3cdbAnkkXDqCC1Y2476DDmmrgUyx7p6fQGdD3pTpqplKMZ46G6DtThxO8pw3CizJ0f
s0UVYHwdUPGZhwZhx1pw34/9N0dqV2CFkyOsEEyXIoPtJ/4fImhY56kxpyVDw7AEIl7nDYc1tZCh
JyHlBvn+G4T5d+L6B4xoMrdgrrWbITjB+k8Ge7F6WJ0BD2cYfJQhz8Q+xJQmfISUi+4MrzF8G/3y
yRM0BE12TWHadFKn9SbZeEMx2/f5NqN5Wemy9mPItr4I8trNzncPUDgo505oeIVtFZKrl1MvCZIl
EjsMbxSU2jA4TwtUNtHbeHcMIEqJ//UVMfPTYECKQbuku1hr2gIyzYM8cI/OB1IXSAqpTuPDaNAQ
ECEvYNdxzaTqZXiMrsYMHkYN6F6dEAu4XdB8Ns11vH/nzYQ+uq5BvYvgZeQtUrFrCVbmOVkcuPm1
J/kgwF9T8l+TRj6uc3SkWd2XGaFy/wKLnODFLzVxptKPvEO7T5lvSQhTYLI6I65Q3Ba2VJJUNXd2
iY9vmfk5k1fkpBQQgRvUsmwxYe/9HyiMLo5/1g/tQC+qCsWTRiQ9dn4hnQPJa58gwaPFDGTO2YGz
kZJCzOtfVfYJivkS8crWhi+895QgMNwoBrOHDk8SY5e/KbdU+g20f6AZI5028lEVndT5qT999XsH
vLpMsF+cv7Jm9GLW+59C9soEENGxLvAwVKoaNTOd9hdwsVkHsjVVDdt6yt8uAym8xZcb/2qSNNM8
SfWWLuxNL7G+KjBOXf8Pl1IGdb6paMRpJHjvdNSsjPnzo3n6A2koryc+YCydAxGpOIvQrOT2QEzV
1zLZDWheU6r+2D50ku9+rEa6U88IXKRlgmMJNtYsKyc2KTL5u5v30dhmqvSN9z0O63C5eYbp38M8
NSVgOubggQAYX4ObpG/uAgDwxggJqE/EXeDbYkyXQIs1jLE8jeCHuCZ7em/KSPJ0en65MrgI6vnN
Y7S//7Fq6zp5KFO+c8OTXSyeDQwp1kjDwYq7t/nGhaGInz9AV/xeNuZ+JVUtMNDf5sxcEThaZ58M
AN0wYcYpP65bdG5ibwQpGSOZK7Af3+jbs3/vj3ePCBzFz+xiJEshThOeicOhSLHtE31jFP7s4DWu
QQ3zzDeL/gf8jSTmTFHeNV0/PYeziYqIqT5QUzHwuvhFlfYmoMrkAwrByEvoOquCamZCD4rXZ+ql
Jag5JtoIDnlSai2yM7DTVbmwZAtzF7PSGdhFap2IGjlCTC8P0zNqoFgA7UZvZexziPDNrI12qkso
V1K6GprrAjQB899DzdVNgj4CfB8KZ1p7EVw3Ka6/8Lo0OElI83ebk7Llj29YMX7DbYiX7iXL0dme
KLmHurDCHbs+xIPPOxgvjE2nM6H6bn+oAXCP1kx6f7iSKRGe7GMIl3C9/eQJRA7CWA+eoQo7Q4zW
1V/qNlVdLFvsHb1Bb/dHPvsWbfzGb3n0i1/Z4rtH55dEv9CUfC1w6TjbGUzlI/VquemJEU71asTS
+hnsC8f+7dlAx+6GZlYat7ymY6moPx7TJCfgy743gX3XRathCpSKVWfjQqPp5HMuoX7sVdF7fgse
5dwevihLbroStKMohJgMUBwz2qhE5PooR89jT8meczwduNSR8fjcc0SwOlk1Op1piedJAnQkJrtb
s8l6QdL6kQnhsNZGHz7j3hGt8LxOg34gDFxhujYTF7xJE7FSdPO0rI+Myh9y5yF5AQujMHbXi0br
3XGeV+lsopaIe/JPbZm8h5Cw5AESeCAjHbtqf10TGiIAszwO2IE+s57tdiKsZz5To/CiLRrzr32J
z8ORlWecATE+yLZ2hRe75o9Zh+mT7V1aLQevmMeYq8VHfcXI14XZbXN0FEJu5asFV8NlyhKzaFwR
GdRwxIgYaK4sftt+7dAgj7jWZKQsw+2w7TZ1wLTVf0e1RtPxVHpBVlos4+J/baEz04nbEURwCbf9
Xu+GX5e2p2QcL+cWVFrTBkKtoBPA7mCrjX+5dEvpU81qXhen8NfVgdiuUek5gssQIIsICeJoOWma
KzEh98iNK37guxntl73M2kmggXXNFZcTojtfsiIdnMhv30G3YcyUpY9y1+Uzpc9meZODxdkPp8QP
4TaefeCgLoyExVUvokWFwpw4zCuhsFZmkvMfYPjRAgTc27KY2X25Pt9eKRmPfCAMnLhof1VxC98S
tgMS8vkUW7Y27qHhP0xTufINRlxVSFmz/bSWO2toRPjgnK6ZQ50qxvRGOOhgssQycoh4lhRbbAR7
uPrfMrt0NDaat9HWCqR+tw87vl6a2O3IQupgABNCkIAjvRMEpfZSK4EHbxZ62wXFElK65MtIPi+s
Htq7ibEHQdAylSxfRDoPoCeDfX0PjTm+TmussnClgKCY0wiz46W8NlQc9qn7WnJeP9SMKTCPgDbt
Yn87rNV4fWHCBmPeqUlATzrFowgk/rzvA0Er1RQKr7PxGpaxUsRiKT9mFdAl55rwZUNaQtXT2gzL
uWLJmH1KW6rW1diVf2S3AajjUe5dgP02co+oFZcl+Xrm9Fub78Ex0z8YxPYmfTuK+DUJOiD1Ez0I
Uke3RTZbxubRIprGWxIuc7HlcmctHDLkazQ/URnYs0D1aLB3jUmCqbq6eDVOMhXdFuWjovo0jQdw
DIqMxW20xUTMhlG6EdVGEm6nv5IS40SnsdRWRZ7f1pVFr3aHp1OL+FDtlZEhyXQhPBL/+OHVbRC3
3wozjJGTWOeNU+PSAc5BJ41rpkPAH2FZPKSkM6Oj53idEdmX5UsoL724TKwVH5VTXzd56aDprKRe
+BJbFIHV8MavCVWfgsQF+mjcd3xNDg+lI7UkX6l0b6FQaGHEsAYbCRFkoEijvjCNP1g4IHLYRC22
SKKPXshuQkPeRkc+b9Uyu3mLw6JbYrsEhEQ/1jGUJQL9ayTLqVwXqkw3kBFp3H6kfi3YUDT/TCne
p6xlpI+Yb8Hz1tJotaGqYtYAeZ7mQHZLrGKgpRhAssx6wQTeQJQRfzHX9RLcX8kL9w1EAex3ja96
C8aW/Z2GCCGi7tW/T8xqG8pc2s58xAfNz9AgG+QbDSIeRdbhe3lOWA45zdb/SxZcrNLbNXciMFAA
7b1LaIlzGf873WHI2O9jioGddaya6WllItGxvKYKfdZYiklfsyI/Zil/1Rey+Px3cdB/n3bXjEhk
5d120ml48nOdFaWq7v/COtaIY34fHHkPrdTQNVWnoyMxCioKMFvwjKWyoGKgS/VC+5mj+f7yNpRV
if1VADaqExR8jk8cSRvVWVR8dEf18uLemkLBK3KbeXNCynci55yDjZPAqEWKKTMstIa9em4WhULU
RbnHbVFIQ/28exBWzEdWlYWzKGuBO86ksg8IpdflqAwEDPgXlOkSG3PZ+nIqM8pF7m1lsc5hX+P4
roovnJ0vx5Ym8cnPhgmlIFcpHTNbG+huB/GoV8S3WN4TiU+n/UL/hauVR2H5OTl0YBH9+AitnPTr
OG2ccH4EuZ5lUlU9YsrC38OpL3MtBCzCCNYNX2ccg8JhUlSUdZh1+eIYmcKuVt9V8svdLzG+nMIb
Mzre7ifEslZO5RH4uJb/MaoCuF9b7WZpqO4rEG8X5C+1/lvk8ulmPSajUuzVLzvSq5dpXTT37UaE
dKOU77N0dT8wl3vDQYLCc+JzULo7HSOQQdUx+bYfFVMQb3iQYviKnb9ooBO5UaXsh05TyvN30mSO
dDyR6dLa0smWgZPD+n1jWwMqTUJ9c2nFxfALlbJs2ChkfTctxJ0fmESiuJhPasclg314uqlwugt9
NJB62YVAOWIWRp/gTvs5UnL6Eqt/10lvaeKAv2kqJ6uPBofQuXTm7C/MX/+fO110YTAzn5ajTUIr
fTljfTdQYu/QA5eBS2I80D+pxqFibfvVZmrBbxTqt06gth9aQmxcVPDh69OtZVCXXzVutwIWp+2E
pIS68T43ft26gF8NVWzbkU8mflDHTnwJMXaWSQRHmTZMOoYt/Xd36qHTrTcyGwENDmYPouHpG9cw
aAHCyWHtYKCpQ5Qkyyr0MVQHtjDpD25MliyFx30jcg1XzNaGYMhkT7eCEmhQh9Y1hkrSgYY+RIYi
1mv45/XF4GCG1sAMyh/+FJIv2hs3ygAvaJBULwgE++5eSCGnj63FE2tRP6DkPJE4D/9F2FpDHqdE
HuVBwdwlZowOOoAdfFNdLLSocG3lW1bt6adxTLdEo9nOJsUs84YnbaEF06vp7krroGjtiMnpX1Xl
SCkTuuUHHXnO+JJrv2alZbtfLeCxjVHEnr0mfdE726rs0VprIwXLvuXEwR5EikZv/gsraEeTPq/w
k6aUSRAgIb6rDA9WfLMHNvDsB4U5t8HC+8cQ/pMg/3znKSjufoC9CYGrwK3TnoWHkQIjGeX5N1dV
m52WbMioG60RI6c7ETx3XPj3NGwQdXKz3HqOW3SWg28xTBAMLX2gHXAJfDEHzdDYN8gHN68VrtO7
pfWzW9rE9Ybqk6cKgm9wQhYbm3FQ1x1PtOAcasFUGTLRNKG8MrTBrAXWqdUtyRV9b9dsElhze5D0
RWa5GXWa09psRqS80rNURZyIN8EKIFg1BV/6h9U/8Agq2WHOBrFbQwEGRrytfkO1RG3yVl1YJ7Yg
ET0hBjer72muvaxSS4d9iqE2FiyRjeiPVGstQJwnNPH5+tKjTJ4NC+R7DKThLq0/24CarCeQCn0s
9cCmUB8PDp7fNaMWoEP0w8Qcdxlbylv2Xj40q+9Fd27Z5ttnlbIW4Tu1Xi6ASu1JIzVyfZlMMDYV
SC1UhLQf9XDPP117YNgJmYR22VJfU4SkGkuBYE/IEHy2Jg2e3zrOMPBp66OJFF/iu+pd+GKUDLu4
D1A7b6+8q8sA6/6fKNyJUUQT8MLn4TUoxr3iUjqpm0w4zxd1a4iBTTnYY6rDYQZ10S+S0WZb4yVi
V7IvX8GWOQQHE/ZEdY2fnpfg8/WjWkq1g90kFUfZxWUKiFOfu0Y+V+fHuznVrIf8R8dv2n6ulZwd
xsqfVnsIN6bdnZ44HSnN7pSlrKjEtpLofslrjI3CHACd2rc4nYPubEIKVrnYIzL/GPYtsxDxQ0wo
62rqLfXQNomElyIwFkiVZEeT1TN4JeGUD6a8syNbH0V1R7Pi+3NXJTwzkbCGGcPSDgFWmsN7myUx
4P8GRLE5qONN4YdtcqBfajmj/AldlzRI5aGL2lIr7Mc6fLKceoa7g92+AD5sSoji7kJo8mRaUwNQ
2LMVwwjfo5rSIMmRVbJpcSGORv3JN2fajEt2oR8vGN6tj8IIbkRZGC5qcmX9IkdIKH2fgoZbovyW
18MO8gIPdQSVUzIsFHF/CPTllPFzRU/3ASNpwtijMsZb2ayxWCW/iN69VEryHBG6+r6gkph0mVjI
4Iy4zJYPMFmbngqFOINv3VSFxTfR1ArwSMI4uWTQXCpPn9qUlKjB5Q6YOJPPSkUB7uHSzxXD9xtZ
TUC/XfJKp1IQVe5cHaFKI1T77AxL02VH45wlVYze/iGNwLmkN1rOenXGy2bKk+DwrAYowZQ8/AwD
4WghEfGCNcg7sye1UI0dsv0sMG7mCMdgZwXG+jlpFqaNWEPtYJevivd1f6v/ew8Ga0HhAywVtV3G
K2vawviEZ8N3VdXzbo3dhgdZSda0dMS+NqmBxgcvycFSMuwh5ldRIBXdZmOCifSrkI3S4S8dv636
cEf5JwaSPuQeyKdDCG9Ez4o50xAasnoI6xop/vBuq7G2fWEQspuWiI20AIbR9jVfIhG46j+JgL9r
IzWXUk46E5sqWo21pmFvpvCndXihAtpUN0RoCUOy8Se0ocndKF9kvcN7o4tdtfFoMHYsXAjRlVIw
kkl4AxijKdktvRDUZFjJVbFvRw/dUQw702cCtZ9L7a5EolzBkClkMsvHRAXVuh+I7n5kRXqCgKb9
gAZUtU0G4wMsd+c9K672txUt9qhWMAuzqfEvfL8cDmxKa+JoUhPApyd43/SZ/Lii0CGQ9Ke0wY9h
W0Mx0vcBHRt8G9QzgDH2+x3erdvsCevqKKAKn3j5KY21TK9LrCNE+cWtaN0b/bvqcCIbN9Hkn/fH
/0ouvH+cZHmoivZkXfCzeSRYo8wE+ue7WY3eRbf9Vhx0JXSKWv/uWQlwMKcXibDstEmD54GFuIxO
r62T8uioJ1bokSJV5tXpfdL/PGNxbI2hIS1i1qP49f9HpkN0KvDblLVfnGiNwYo3jPyiRlD1e4lU
3idETxhggVzOxPmE6Z3XOtvxcyWi+P0kJB4PtVPHTw783Z+VTfySp8f5p0IQ28RYLGP1ndXtaVgz
eHtMUXv0hAUpJuDHrdf5LFTPRKA9s7ZVL1WnSgNt28u77cnaGYCCJZFfddf7D82xs/Z2aaYy2C7R
ozSxWfOlFHBuAwnIlb9kBptUJf+YJElQhDIDJLhTUeMzZAggrPLU1cFytOH6HJ6/yJBAUR+y0ONl
WLUWlr/deCfFiPH/HeYrIpL2ZYe8gioEzzeHIx4RB6gKrYdNn2PTPu2xXAXTAldzCJeX03FBNqbX
/I1l1y7VClxc/vm9CDGCgRCsYDhCy85bTK41m/T1ERNJKD1ARHJQO5ocTuy3P0ywhbRKtGebgdot
QujQFV+KrR5PIMPpYw5ZUF6XtkXvRr6SvgIMgxbIMM+3hGMiwsx3bSNhKJONkTjAXfFTmya7jlyV
j4mucGn0Xd0tEwEh5TygoEvRgZLjIGfq+i0wPZJacqqcLsbGim0DSvZT0mY9qhuUBCgpqbc8N9HD
/2laN8EsEKKiogkwcST0mP13r1LF29vone5nUBwFAI4TBz8CY86241/OCfDdD3yjIcdvN23hMqvw
tar4Ee1+8OU2yJUdeFxpmOmAXsuAjZm9q2eegHDpWBh5Ms26DGbUshLX2GqnTJUVN7o4KWcBbE9E
VInxQXB37Um7mKv+X1iUjM/inqjN/DuiGpBkBqk2QsqOuf+EkCPnc18OEDVq7mzEy80x8Aebg2Dq
eX/UfhuioDct4osPrOGlLTcWt/GSa505pGLh7gjoSqyfvq3xne3ycPQdinZwFla8rWBKzrIbS3tu
aLHU+FCWHcToyN2kkqOy2h62wNZ0ZlnBTGucgxPR+9oBVzucclm+KhrGYI5FnrtQHKRsg2uC0H7u
rVD/xJkPZGVbf8Ql8oyHbMcPiuZeItDLIuRczg3yPBco9q5R+AsmVDxwNtqUwr8P82g07gkwysoe
TllqNX/QbNrJ+0lt7H+AwBZGJopoFujXhMpDiIG+VA3cKDioro2WMMqHnAGuYq0DP3JoTZa4CqxF
2B2Dfb5DdVU7umXoUAGC3qU2wkuJdLRqjVp2hdf0feUwt+7RkKEJ49+SOlBrW+x+TqhT4PCUVQu/
+bKd6rs2++yWMkR+r9hEeBkDxrN7i+nMOVXOf/fN0+xxJKFw81rB09eVIe6/GG5kTyLf/rkBjn88
yeZRrygXJV8arfeSYwcsofvzVdTosK1F4U5cDQR8F0biT9ey5kkiP9ma4ZxxICpLoJAVf6OzZUTT
DD+0KUFonRLROe5cnqz8U+tE+3XYdxTVLrHbWnKURoBWbGfg73MPVm/H/uTvtjkOIKAN26Q06SDy
hPiKalBdOxkKh9SYvtWX4lGB8mqKzL5SwY7JisqcueyJCQefKO02FsFy8YFWJUAzo4iXWT0Xcocg
XtZtHKQPldPUw8y9p0x+fYd+QPp89smAN35VTG5b93L94Tvl15gL8JICDS6gs2ruLQR0wdXL4iBa
bl9hS+GCF/32XxSCe3jv9wB68H9n31m6e/53Hcr1dx7MeBkyvDOuVCPdzJp4e+fv46wbRLJyT8/G
w6dGs/86Eal8jrGJJp2gEvxbpJPk+Z0PxVUUmZfRvKCENMyr6JrkRICWJlCPUtzZi0kIWcKTTe8s
oTg4VUw9sLutE68a69KPBiNg/Bp+yg3JDTlyKo0LeGFXygTpPsy01+T1o8NF84U407TgDZ33rWSJ
jN4a33c5b8jvIxnbBnOwG018EYXZFNP9pXGJUFEStqjqK12f1S4n7sybQ4aeUwkwHUhlHxGtZKqC
nDUmkBvM+VoNk9/i8D+smPvbvVQtGFA/RlcJv8sxFCxvvLpIssAZMTZvzHq42FF5OgF27oj/LYLc
5ohY4n3M3HjKrlwUn5bH4Jz8qA9RcwuTOy0YRrWXmaZr7k2QhMGDFqW6dt0vxiGY5G89kjnQMNKA
O/QDt2eN5VxNzHmLJ0ixm0LKfFjXL4ASPga3fDqAU+3QB54EhVUWWHxu03p5TGJN3yzg+E8lXiaE
8KV7nE980AMApZsfcqvtPQj42UPm6STThsExZomF+74C+9CXTWTIshrAyrwazv33ph67fSdaTXZ8
I6fP81VybSaiGWUQsIo+EbHS41MJUJAL1/ChXv1xDDpERlMbFlyIUsIbpfvziuIA/shzUJiyQTuH
+AsgGIO3XnMbnLaBAHBgEANnLLMxR2VlPPFW7pUBoG5oZFnguHLeFVJrHgV5Ogtt0rQfzBTxhJrb
uOdYVm8DHPSVQ5ittPABCKlFJhXGtJyXzs5LCwPz0V3O7teJBWMrMQ6ZK+s/c3/2A8En2fOBHa8C
OlBdkeJnlkF7RCrsp99aT+8iL5M5ICUZyC+US0rOk444YpfMI4dBhvfTLKi/nMZzJa0+AQj2GnVd
yDH7jlofxpQ4id9hH9abrc1TugNf24pyyiTkzlYKBsGy7H9YpR7r7cNt3gwwIxI9USjHXHI+QGH0
6ZguwIrYRtpKhBw3J4VHUzpDH5B23tp8lp185LvqlzB7CQ6DAUyf3kALi4MJwVWkqhkOJCFcXYGz
yNPErt17zi/lkMuaqy16YJXvZnBL1N7RuosY3rlgI2yeoWUYDEYBIuUzmVuP8kl9RvFslAeL4qiE
ODM8IYDyi1oGiWvzMCaRaJjfqhYva6qX7rlnfSgemnsWYgydIQ9opzO2Lod0oX22vm5apvx+y/NE
Cm88qNbYmBUBsj28Ha9FDpRpM1VWY4tG7e75Q71WxR3SjK+Y+h9fiIEMEItWBekXHZvyNDe1Gaod
sXC1o1IoVdpOa66gXhskN91xmQ714rc0RvRr6ONQ4bglrFtmCqytjF/FhUFK0vz44BBDWaas2kXd
J3p63tUd9KDNfNBKG5abQbxplFppKztVMNh/2uxp9QbZNeFFegrL7tQYRZH2k2/3U86xDZlmZegl
TsUeRIHgDIUIJLVBbT+O5/XXs1vOhrgVpZcjTbRsYoL0b/ChBnJVy/7xYwdX/FuHt+o/MJfK6xkc
auabt+3/0KfGiXRL0Zv8bvhC1Y6LeJXqLacSjTIHfqZX9lXqoxJqePCJsEAEQMJ8dXPYJ1Jboy1L
RyU+uw7+DjGKYltjFo3TWhCuejICRU8iGjEKopps4KLPwwklX4a+q/q7LDImcCavOsk/CKzaokDl
gBYiePDN/rGaeTX8EsQuAqW7ZKxWKFiaZBghDhAG18gjiX0rLgzzLkLpnVrwe0jFYz8AQYVta+2B
IqUd3UK+rW8/fkcdMQEgdzJt5qTyU39lfEwV1QfhmDhxYqAFxJmdGRmR/Xzzlf1SSiTdWB7fBpuD
t3Ip14PaxRRJ1nmN9dc2gBf6TSiI4nXRmDoqA9JNphWAZifT8mZMbTyQs8wpymHQzc60f1R2bzqR
4SWLwVlPlLRmsioMuMNJDztg9KZbfVX3axvhY4h5Aoxs5lr9TvZIpkUHZO09urUUUcz9iw7zU8ra
6Eetxu2OTxfFQ0/Mhp/X7betNvC2rebLVuXKxzRaQn8sHfwag/m1IXvGMCauT0H3GATJWD4bIqF3
mEH3eVtozhp1BRLvWQo4zi9vWPmnnjNHrzjSkmOPxoG7Mz/YMyLbGt8Au/FFigna2oBbDIOrHYsT
lI7aYBG2O2E5/JlhybuDVxrnp933t99zyB0b8E6vWSA0J+djEKDaD7hS0ayRGWqRz+/eZw7fAHfM
MVOVkgzMHO0vYpSgnzAQskeourzBtSytHyLEIvBPxGnZtiUURoAo0cvXk9lh4gRJ36haSyCjEf64
jCuYJUAqKK9zlns1MwhmUkclxkICLAxjpxrokje7v5Q+VoPln7tAtu02ywDpAZl7fQaxD5jaJRRR
+52a3ibINYSycuVWzAyCbQ1ZD8aaASvEevq37RlJCfyz4BPiZ2PdBEJKPo9QCPYzkYdFqof6QCeJ
i1MZtnPmVX4a7WFoY5mRY/ujZg0r749XqwBrUp8ob/MbCTco+lNq9Hh0Dd2k9zla7h+O6SkqEgzE
e5eecio+TUiZQUwsQoMAMVQPLgFbPXT+4MvTsbFBTSZX4/DcFb4mTaN6m9FR3jD+WiQ1nnQvJXvD
DGPD5UgGgswOU9UHfcCfEMJFDoOpK2VmxJkX/Jiu3W+l9qgb4Xkzddv1OpioVN2xY67ltQEamSLo
Hya+QY/ByviJwOc2KoCvaGgPdzR1twpqbPcxX3F1dFAOHgBazalfxzYGjfwPUU0dGaKGZL7G3Nte
IUfmkjJe9F7pyU8JNA/7eP/5u1AYReSA1PoySe4VssaMzNEckzUCUTeylOwd8ZC/LngPZy9wHJYw
eCM+tQULJGL00Th8PSnPFA7WjLD2/7IRU4QBM0UcILmeEGqh+VeiWP10LErnBaHdgWOmbGRZsS8Z
kEkMd+lW0r3p7PDZRHJPHhwNkJSkLAs9k2RphhFaHolKTs59B+3E3NAwKkAiir/8FSzoZbe2z6vN
jbXF2RHZk10aqSbxtbsVITINbRFsKPadPaTftXExZ8vMAdIOE7PjtVXm3z/etpXdshW9R2/WpC6c
kT21z4vaV0hKEUNbuYlEXoNtgQHm+R4vjGQVvU3Vn7yKbUWw+1Q4SO82iIczdt6I6DcqV26GTdoG
lWl3ir6EK/O3gq004Oxekfz9RpXjkblILuFxszhvAnE25zyEoh8ySVWF1VL26REygm8BmD1sNOqs
zKJkdf6oXjdg6rCtuRkcHGIbj1zMiH9rl1tQSxjreC/3mCV1nre3UYrv7QfqANuPpjj5PytNIkiA
K0dYk2TxsK1T1iD40AM9k/3JlbobzuOSTLjxeqwR8kY40XhJY358NGvbzNMXvFc0hsU4a/vR5Tiw
SgKmapQEv5Cqhg8QmPCekwoW9Apm3O9o7//UGFX9Ri87FIjsLqAT30cISeKd2NEKD8ztmlBImnz5
uWatYtR5E+CehWH/iXuPMKrwIM9eiIPl4G+QSCtu/17TbuKdHS8DVljYHAnFo+PvOoBR/QtwRnuW
YtFOb94IuqpVgD/wYm8EizSkjTEKsR2AHIoVv2Bb07QKkIqc9hiI4yyPV9ooz4DeQMWRic0NSYbr
2yNG6sWQapgbs5mWg+PdARCfzdVJZjACbOz2IQABVdQTWVrAv7HGLmdUSGpJqC2MZOqCz/9K8YTX
vzud5QbBi11IfcOgRo1zUw3rkIbgdUDhR4Uiew5uL7jgN/bGU96Od3aMw7+kLnz6iAhAl1R3Ybbo
xEgzcyUnIeTZ5o3fnS9YSfBJlijTpr508WDzTaa5Uk8zP5d3qg15JaPU4pA8MGbRCMY/p+Gy4KkV
/9rpDKxC6W6/9Ee25zK4ti727r56hkPBFbOJWT9Gx3Ny5L3QBse7YZe3u1aK/QEK3HP/EgxJVrcY
2OG0RFr81wFTlJQwNBH052pEk5++LEZ3ihgMdoayECS5IU7rwBXKMl5B2jR8egnBR7mQGRAtwPaL
eJ1R3CrdE/YpUBEcujNWo1dQXOBTLMDOZpBv8Br9ikRM+VbuxZUVInxkLsdyMMDyM6Xl0WiWVvge
px7ucmR3EwE4POorjCikrL39595Tep6YIeqXPJWHkkwUaJPdIq3IR8doUatZzJsa6ZeVCErwQjji
3caglgRvvXMqwOgaiiEmLQnKJu8TLyuEc6MFD4g4iG1AiZNNtLnYOzrrLCUF51ZM/ZDc86bvOFzz
E17JpyUgG0JxJ1v9vn0gxSnyOxGD8qSitvQinY3W8m4rnhqM0YfLBlCsntElvjAJsmmqAkWxPftC
4rmhOtE506Bcgt5Thy5/fiqGpIeTUTCNAZK5h+xExaLUgHdqIUXcOCEKhlTUyC5PuCxoir0TwKZc
+Eh9bcV7s5ta8JVHL21uXqkRFlirg1T0Dk/A6s6qEpemvu42AJ2NmGpcZxE4SvZr0TbuhPotLYoQ
EEmPN13KX7I9VyJIyxn+xEK8+EWlC4FRcs5EkVE6q8kYbqZMed3jkk0PwHksofTYo289OM8wqEZW
xqxSvImzYMEbXLFj66yNzub+MrU6Ko3YYx7i9AWOghn/DzT4V/t+0gFHegwp3nRkDwohNtDHwmUP
Mx5pp/6r0r+mLyiwJG8oJTIlYQOOkqRZESDAeOrxNA6lXsPSGN6DRCX4Zjfuxr1kHTnHsUdoYatp
zY9FIrT4JEVmhQQuGekosmfYjVA+H6QRQG53mOJr0DB+XV2/U8pTWDyJ8Lgv/ZWtZX9z5utIqAmh
Gkl1lBLmUVOvuf8QcCh5ItbhpIxAiNGgvZFrMz3K8uw/0DfC64V3jsRDyz+sTDHuVXrZwXNcYu+F
JW7iQv+H0GK+jxH/O4KHZ5M4PkhSbJOo1iKWla8bnyJ6zoswnYqcB1rfi7+7SFNfDoWopnfCzPeW
XxFh4m9uk4X8ecsu/RrziT61eBmRMReMa/o+xuxP7gAI/r1I0T3sihvEV2KMxYP3xbFhBam76LMC
QE59OAj15q000/zwMl/JlnT26th1fiDRFLVb33hwmahyMFArlhU7tfvStIJKqfBGkBEmQTYMSlzn
l0fpDnprMOkTjhyxBbqL2FVrUak7dNghZKfCZRK+bLIMi/IpDyoLTXAAoTwPsDVCsWrA1ydCT21o
OwmrUVsr7GuJi1dvdBwzo1UHb6MHA1kf5rnmz5Bioe9IcO/En+e3xECFRU0AKUe61BT61fef327G
vjMUgJ5HjaZp7X4GPXSEbquj961yJ1CC/3uotsJDH8I4LW3zkF4REP3R0Aj05DStEvwpgLT2I/7+
675ZEbmyjdHVD0hsKXyDrlxZC9BLjnuOlqVxMPZVMZ+5rHNCMObQZe4UdsV8GBYrQWDKQ/9u4RBx
8I3XgSQETiEoXWEEcJLumiSvnEa9xYIRkvrbq7TWtjfOjJqcBZ0wLozMyJgkvuAK9BuQ/w3SLETl
4kiOAL9dVeNjgKpOTHDhUFY5puoKVoi1mSJRjYXRJ4cN4j9/3aL8Z5bhoOyle16R3STjnQDd3Jfs
c41mZfgSJcQWENdhEgzUJ7HP60e2rMSKOEXVN56+jmuYc5qItgIw7LvoKEA+S9tW+03T1o5pbIE6
Zs3dVWYF/VL57PXCG+oGC6tcYGRC2N3qZEBhNcig4VDFD7U0nLtf7AAa+oBLEUerG9hoa7ZGQ/Gw
xmPTExrxqlIbVTPztpV0WG/RiTreQrmV/nX52J1IjAOH3JZb7uNExwlR32xxKCLjn82IA4/SfozH
M9zSdJJTl0XrPXUxoPSreM8y2zJ7bZnWlwWoafuBLqmsyk7qLxe6mTVRXI8O5j2GZwS9QUwNnLbO
WDh/loNZ9BmmZqyuAzfwCpWmIMPHH1L+uNZS/aET46891LQYStspMe6gbZCmhbK1CunjzUfkzu87
slkTe1yigOcA+tKXlRK5sK4pgADQ3Dd4LPTivU0I1W6640YaRTx/qwMHPZPvlU2uP6KpHfOsygFS
higMWOhBAI+F27/qHHgFL2WMK07D3rMn1nlyx2SYBvN+p8Lj2G2AX5xwsMTflP68MZ9MRaHPqE5J
TYaJ7CJ5afzl0U0p9r1yfyzKdSeDXwUeHaJyOwxffxvP6ZIWLsbxYNkBLNKfyJa6G4zqjxTse6an
Y6FebRMRDCF5YDOFvI98J6UDSEKbGAogiOqvN/UUahHQZdg484h8pkiFMCM5pkRGiL57DX3kLLav
Ib6bRgdUsjernqNpZx34ctjx0WxjYjwyRCoimj7A5UvKdNy+wjY8TLGN6ZS3Qow0Rx9/hhM/mXHt
c1uWPLHZhQAkWlELVA6cFhPXS0MidC7b+1bVKmPEiIXh3jnODyyEHVGtbTqGu5pXj35vUH5HiUD+
HHoSJF+/D9Y3iWdg6PE4eMe8ZCiLnFXCzQKCGPBKp7heYoibFZI5ux6JXzmaAht+lThzNtQrmKa6
H6yE9kpK0Q+5Uit0hmWmxToS3K1Oeb4Ip3yEo89lLbHQ5x5zsImVlrpFuDzoiY2XKVKSkvXuYUv4
/jBGiQ3Y5HVrc29Vtl7y0rxvDAnRG/ekoDua9LUE6r4YvRdqgjqvEJq6f15t8fpFCdhDh3LvY50l
xomEg7sjDSH0cFP4uHc6nV5uXQjnm2d7VimgnmG7ErZh9H8HyoqxHcViv3pKNAI3kYuNUDDKKtch
GhYdBU7vqBtDUQdo1b2j2W1cf4mBwvgrmhXD9Ynw06sT3BlcBquAIJRTuv72duE7dtBMqzvd5f9j
kvStIi+ZOGbUKQswzlCEKoh6Lp86VkxkIp4Wfm9/BAmwJX/7GjC45iphyOVU03mdlpmIvl12ZFPh
6ZnxUczFBVn7N4103f/hVWyU0h7HIoF9SCoJHE0Aem97MMs6h5fKGcC/7iqr2ZPE2ImmkQo/wXhs
hGFGoos3qeGCHePnz8+iG+C9d8B2x0D1Wf22i/GHthaN/h20D39XFxlHA7RT1SESJYqFCXRSBP3Y
VpvzgxX8d+3yvu6vyIMkXqEZ8jUpgvZgIeeuIKiF62E3OTHSxEbjT+CVYQmd1/65md4iluncL3NL
jZj7MKaxVV/w2arp1rbNINb0Ss9XNOMvmq6e63tfz/BzIJuFsZOqNYRavFX026sBWva+iZVR79Re
LNMj3ocrvmY3wY/F84TWqml6tLqfg3cUwuchvuyFkMWvnQB9IFk4ufaC/7RVWuvW4E55RInIbDSC
Lv4FHhDmuQ3fZd8Gfn+6nVhrKRLvEtfrOs1p+N30b3m1EFRF9vpyetiA3oCTU2q0kOSPMiu/FSTK
iCND5RamHb0zPsWeiYVo5ijr2FSU1vWduDNM2IUYC7ny6S6WCbXRCH/92L6zxdOmyqHPp1Sh3SAY
UulIIgK7h0/0KycSVeZXQB0QaGkB/FJLL6N/LrACYeHSR1V7ojWAR6ggeyg1rkCoSId8y3Ggm2P1
rDbUQm+BJ5fVvULVn4bK9XvE7BJkwCXXKLTh7iJC6lQooEnU1J109VfgV+EcPUGmWbbQmpXWyEhT
2tXALn+E/yrCW/er99OXeOt5MAOlkZwFclxaZ0EmZUDuHmq9yqVTi419mb8Vy4fl9v8EYkquYdtA
+ZltWGXvLhQlTCPXsdkQniyYMlvM78XDsmBFndNnRlSPBviITpfgw3+PVO2P5UyzAfLj8lex7aGC
TD8wqknECAmgm+4/0+fuHcRAHUyHs5qOF5fQc/usMVbiNqQLvtLAw01mvbSSkeMhW6TmFjDJPvl+
r0pZ41TIfiIXbqICSYvGqJE7yBPzxTk8s0L5X8+Fv09jDJtt6JnWbuYu6Hssl4twZ1uDva3Jtsdm
jW5+QnTERS3xKfu4EPSNjEseV3KcU7wi2dMLuQ617Q6CiH1IBdbmbhL82cqSxK4o8W2rFREEEEX3
Hk4KHOOrzPFOmxQNhEWS0C+8gP9Eb79GbAoXjh21qblfyFoeB83I7YVLfjUm7Qa8yV4yrcNQ+cFD
1kIBHcKgVrtIbV7OuPEhvsRQ9J0wvyvMwxqztj2zGb/cd9nit8V3vqngEHXBL8I2ngZ4i7vLOF9p
LlVvlR86I+cmx8F37ZgIBSESnwCD0BzNgiwWVPFeDMRybruTNEITL9Uo7er33gIU3BGxqlJXfkZz
vPgL1DOgZydS3vE377UviQTF9sVyWDA7eYLi24t0lRPWVeeabC5l4CbIFgIS/2vXE7Um7GykCko0
R7jvn/ZG9Oy4Wxgj6zpVZfLqcKuSEqtGJRHc/OYn04xoIqILc9X26mUXxJZ1Idaoe91dGDdjETHs
CIjrJslWVzAG/1H6UmOEJNVlb1vR9tRG9gnDONAro+tcjerhKHD0Z7cpPEOCZqvdourz0bIa3NFd
zvFW07QBu4zUyAI7o6je7xtQkc+jXBE6EUNS8dauzPZVqreujtYanYMlKcyh10r3lbQ3pN714N0y
kPIruHDyDnVnvxC5Hj7+j0f5BTr26Naid/TKsBOykAsEyfHi76HI65hC3MZ6kV12VO/tfSAKp51q
/krpZKnjVcNM1OxOb0oCHKGUmZdJtxy2bbQfwDP63DzqUbXuEiW/L3JoJhUe4pvcHNHgjrYwnDmM
/Xn/NjsaJl28g3u737st+1r8JJ6DL2IAsxqwNaeFUHGPDd7wkKIYHSKnc8T2ic0aFqizzHui+E4w
gmETHKUTrzFn5wjwYoIkC83BKv2wiucV6WBsgsVMQruFDGi0pAodZiLRz9lDOHakZf31I4xEboWQ
0YoaBvELy6b67M8vqDn502XHrjcZvFAwgsTr+vb42TR3AINkoCmo2xzv7fuBqdw2Vjsci+1dGIwP
sZu/6vLFeUlMbKGkjpsfwILNldQiYG6R74tBSPg/iD8yKyHPe7D1MlInIWApHjcysfuZjvGACMdQ
6O7tMMU0qxCve3Rk7LSUHcfRlbY4qxe2h88/X5As4Jl/3SObCqbBnC2wlZtglCb+2F1JBVKmAQSV
9z/Pd2A3AaleH+4QBsFyh142s8nOszE9Fz4hc4oC0Yijy6riusBpwEx2XSFot77rLdESTCjkoC+s
N2bXUY0KV8srbnbt4ZIXUd9Me4QstbVDH9CLuAPHPEnCKBSnO+zL/vzGmZQwTo5LiCe1G3vyeTAw
5JC8kVBOLwWT2BhW5Xb5rxhM/bW4u2fEsG0X8FloNRT6IWD8W/3DBYQzGLyRCooLvHKKjOWeWbFN
Su5S1gpXOOEHPjhza3xY8xh1ycliTG15pbKQ/ohbn/7kMqWvRDiy36iGJWo3UUjdfHKsaG3PUJzK
YXHltRUBXoQYOjGzNmiu2V/FcHY4c4Qr+U+g7nJpBNRNajrYSJHeItJ/wsEBgGheqFBXh+9FhI3o
gEE76OWYT8vzO9X0Ag3yIOhnsN3ZInKWUf9loA8MCcq3wpeiHXD0+Uh3MqQ+iduv/65UlGi1oUYW
JinCzRiaFcS9ZUqTN40SEjPDoSCUMLN1o8PlFstN/mMmqtXv4Vs83IaRelkkX3g1XAJfvhRNbCl+
npNdUPVSq4bXFlbtKEarqI1R5Lo5JcCRB2xp7EFTt6pejgLfQaBd03uffZ1/wkpJfvik36EW6/o3
44t6tBpdnN91S/JyBRU+VfyuKNwCCk0t5tG2N+p9wqhX5yATXEwDmV7y2FDkjxNGcTTR9sHUDcW0
2FxcWOrSA3F+udh5NEO5bJr6YA++hwlVBEavhlwfP8VkZ2Ea5TtB3JVBmkvzUXim3bdhwhDwUpSe
L/XPl24iQRBWLhjcDI8V4d89dDHL9nPTQaMBcjb+5d3JSf+X1bQTu7LFnU00i9sCYUeWcqE9hnCM
i2RsrOlnzwIlrPAjA1fEXkDwJ6otCq7aCYEy0d0O0rppZ1JdiacImZ2nXBWnBecg1ieEdhX3MvSL
Bdb/vr7PWkUC3uyCInXy0Aj5slpbD6uOyn7MCeLaIrmcdfIgtnGgtl9hbdLpZLSB25W2pZfkFFWY
u3MgdTAdniJAffajb5iSB2IxlVDDQq90Kp9wfgSNGB6aK2d/FTnUqzPkFFhWoGXTh0amKVsOgln7
HQ2a10p8z19HPkoVkmehsQGIF5VYP02B3Ggq2fumh9uxuVOvI+yiGqBkqH5tyU7HtMRNZNd9eT9S
c3TocU+cl/ldlaxhRRWjD3E58l5NRK7O15VTZD3DX5A99SOSHGEC+YpAuP7Ir5zBiC95OHEgiqwV
5ptvLTTQxSbufjxQvSij5E1htwMuRQpQ16vxbF3qUZYhFxJKTQ1Hl8qt+wThKjCPyQoCemLS7Xqq
sd0+AV6EmuKGyNZewxOekvEQsqwjwCZjDW3dOsFDHMOBc03hAtSODGKJZgtpSc5MPfyXfUjNT1Rs
yGewpdmkhiGqm96s9bcVARm4wxeexFbeOxDVT7MvvXLKuqdF+C9Slv+cE5hE1t8WaQW0qHgj8Hb7
+mFIPFGpD2wAtcTihGtegbBQDj2GDH0bA4mYhbPVqXiO0UYuRCteoY91rTmPkiIvcqXeQtWdGFSz
HtZhO+mtUyF69100qcHTH04+d8DCfCR1h/Cwj3sfK+pbJQdf7t8rI2it9tU34vtTRftsvnH10PfG
W4zk4E8gkESz4RYrygMeZcuAiS1AHy9fBph2QeuDyRby2GgJRhZLUYH0pnL/i7M2s/jF9NETCM4c
5e+lV9XwC9sNOvHiIRWwkKStbuzSMYid905l8xhsom1cpBoCsoVqEbHavYcdOy8JPUGg8CpzTWxl
94xg1RFCo4aD/ZAfnVLskJlHnwcpFpb/3saVkeHJ8kRzYw85Yml6ttEs50SqnufWa4X1XI9vWSlM
vLtIoz9SK00YlSQZ1aQR9/J2CQK824VxLRW0D+tBPcXokQJTCFylBzMWMuFDoX7XVbNEsib2uooL
Q7cgk30QapzZ1AtheM3G5541pYw1qNGE8xmhhD8iU3DqGqZ5pNjagmSVDoO1mnHlULxVfMIFVqkT
zE1tXwpPgv1mKOxWSRGnMem23naDni2CG9RlfS5BugmqxM6QMJAEtyhqYftwM8IoOVIMTW/2sLUY
tbHbgbG3BV8+a/ISHwwPluspyGqd8JR82upfk+Ccs/hOLvwdfbqyV2Z7zeQfN61D9B2pB5Qcqlq6
bjSctzf+jMtdtsdnkQzyj86RiLpbPmEkWZ52HvPrNenK7TvQvY/3USxmQCK4yUQuUDCnOTQ6urRV
fEW9BaEg1nsAWEy00+rn06pMYFtxwH7fhVQaCvsji8mhMR42EqRhWwkA98VxMxq2mLlR9KWjtmXM
y9JfezN/kk6DGDbALD/VnSLA8t7G3ats97Bl2Jbptu231qMVYkVXCKkp66Z9FCNVU9veG+iLkuml
jIH/cOx6P0qgtqmsGeoj2YuXze4nWikRPhgBEgD5RpmM8GIbXCyVzfn6NqcBaWDCD+OnHlwKKnrB
86/4YHoVl2DskrF8lGLcfiZmmA0nYSnaWQCmQ3BVGDU8GCvWtTM5tzdgATp+YfYRQWEDzOjnd4Ri
gZOOuGqk1jKY1FwZQSrSD7A3ORCmfGeIZG1hWKX5H4KebzxXT81mE9q41A02HhOoh8mgRWIVTpZE
/chTaR5MjgO67ZyAPJ3lSwLChiMvFSGI9Lal0ORwTcNFjqtjtCzEByicM24djbexhCJkJIGsO8pc
E3QE/lErFEroiLdlM0e54yXs7+lyAy1WdiElNgniHEzls5fU+/fziv5/d0WC7Q/ZP/5gz7Wt17EE
nuLGdACYtXJW5kLFC1nrjWGA3JFmeaLEyjAl4EOM080TySLHZ3n3JJ5Sqh4pcR1jJeTUhpi1R6je
rxKZVAS5jsmTw8gEBh3DLDbUH3UOPYOaE3pTIU6w7qKIFwc++Nk6Qn3mYfbi8AGUCr95H9koX78Q
5fS63/bG+Z9r26/dlDehMHwko6i7FIids/XEWtslJVIixPpA0sF6hFqwf5096i67VjMiv+kzKdB8
1eIg4LwYdG2v8PPqJzscgdnd3m0vArJPfplNvvv8fNX03nPBo+KGTeqmRccpZa8pC7WRlfAJsHEf
NDVzHpAnVDVqpZJZ4fjYRzEC78eAcIy44qE1BuSdQwMk7GW4SZX9HDW+vdL2IpQT2e0zbTcLNDLj
EO9QsWzgVXnDhq//Jee2T9U3ENriwkT1Rb7wSgDoUQmucxKYH66KvQrdSV5Rkte5kaLOgScNv2Im
jAmGCJEuRLAcGRSgp6Vxdmmw89RXwUois1sGwjx5uQKXZtoD5KwAgVlA/zBt+Hu8qmTQMcNkkHFi
eoM4ZmbcVCcfU+kFU2VoK5ifz82Yq+r8cyazW+VE3p+sGOqdPPfN3C2bAZjBy/ymQepr+umtIXas
H4k3QweNnCU+5BKOxxzGSyqoqkyw8kJchlcHBM9IROk3+y24zOJ/vqnA9cvFI1g+Sfdg6IEtsq0K
r+JKM5egP6LNhu4I4J1P7HfEIBuPXdFaMqjQkJiaIxqbOhnq7v87sM00ILk52ZRKBwbW5p9+HG9l
HzBf7mCtL/yt82QwpWjNuysdQFcyvAIup5rIAXqJXC90fQZF1RJPMZMrStK7iVY2h/O1EangiHtP
i6IGo6ncd681iUDzSWD06kXPOEL68bKcvb/kcLU6oMNeIj+bLWJ4UdJG4EYQpYLrD/jYJRtvU4y8
lInxoqx+tO4Z0KtbkHTVGWKoakCSVUFp4pd8vvn69J8mE7jyfHRsEWFNIg/Yo/kdCraljf+ERz1M
oedEwh57E1tAHml7NUz5Ul/OK7zh6cA/c4EfE5tTHMozZvQXA7e4gHeCUplFeDkNL1K4/7GloFVj
SNJb7mtejkZyordOKOxtnEv0cSxuP2kUGlfkGF14pke2aWtzjj13kbQxZeTEgcerz5r944zoMp1p
byMY1XaP0pxD9kbIqXavxJyM1OK1ENAX/a44hvvkNG0FxR5KDacbncKbkdxsTLsJiXh04HYO5eC5
QoDgctpMWHYV+I4TSPdbTMifVSZ9oGRGlb2FfEbmbCNFdbLHWZPolV91pEfLT6f1FZBiRkDlTIMz
vntQJHz58gilsCzYqWdSVeN7aLTu8eRVUx6b6zdkTDFrk7D8EBWffTcVkiE/FkwobEnLIvwvE8Ab
nljwXmIeVU8/EqZc+f31pR1vIA0Pl8rqJPyq3f45qm3V52QBfN7EXA+fX1HApVt0iwypgSPDCWUF
BH292ta48u7D/SYxYzxpIkwgt7UEeytj2zWXme5zvyXxT4zwRRVN860QDBRH9N79hHff/5YSH9l9
x7ebW2Ekc5cGFUiY0HbOxmls9TopxaXIBpc5Ygr7lBCGxaOeN5I8quUy1oyo13wkKgF61O3cPd27
mxJcXdU41E8TgOpU31N2nUAQNEbPKSe8yf7TojoMOTXXwXPKISwFN52E8F2qYYlDI+TjEKtz3c+G
ilcWhxDG+rpaBRe1tUW1SevhmoeCEOKI/WqfNx2vuk6gWq0QnnnCbW8cfdONYbPsQE8YmgAz+tPc
oGlbn7YHu5HDWUZgA+Sf7st7eMSiVqcfr9WjRCWix4+yUdTN0w16k7iwF1DvS6/UgeHlm7tjLLUe
mymjBfMnqA5rLemxiHPn9UbTHx93V0IrdLlsuEV0B1EWGQnKuj5aNRYg56Z7QrRQmCWnh6ZnIxSR
fF62fJkxo/gJZOb6uwVJlbeWUzDiRfmOC3GIkUeIELfgbkAyuX7/j8NTk5uc8Pno9xosL5U0zp35
ZKdTiscy76vSI6mMKh4HJtQbou5GeNtLcArBuKaTlMUZl6lvG1y9ttRuwqbT7EqemOrmMDXE3ZSa
4bk7yJtPs9FP01RRiwuUFm8VEpRbG8fMLvI2wd0iobh7n0ywtj3+drm0qZOYu7QcRIIlhW3f6hQ4
JsRDmfehTX6Iov4R3DQuIah6GV7jvCbelY91HBmaJJKuoKfsZh/ymkxc2Ivv8d68hGHQtFSdHSkn
LEAF5qPQbSRysB6V5VeABygLvLoGHilCYMc4Br028JbusKDFS4LHUko2JbjfZilioeHsjP3F3uSC
HLC1P+51/LBJbIerjxyqEHs6BaxtI0MZlffPuFQWcibogc6z9aQVUBCDTbsfscI1w4egq0TeGPzA
F9fnjH1yVJMxxrJ7Q/BE427ejIw4E8iLQTrzkhIIPtW93GN0pqQZRqDik1qpJWinfnk8wKNO+Ewd
vvbCapF6GF6mGxPc53kz3Ze+ffBmmwM9a/FscWkVoNZOyhKmEmzX+acWKHD+j8/SdpKy6AvzcDv5
xaGM/Rwam0BV2Qz7Mm9smmQPeL1aPFKwnrXUAOUrugUV5Hgm7Al43G1dbYJROFYYeRWL2mbhpLI1
JUsgMeyE7yoe3afUNPbq03z+w2Vj+FHZ7/LHoL4V2Gdo+pDLGGKtd4dqN8yyuun2uPoCltr+/LVM
hAYIskTCvgCwU+hn+qOvyOYj7Ai8sVx2PRcjoe2F7ZwrR/RM5qQM1bLCBqqWLAzy9jxJly1108sO
GZbegguB+zWZwTBhearnN7uRRY7xDOo1VB3MH6OxFC6gjSKqF9m2tesOHKCRU+36iYLxG4DKDPXa
zBJMTVfN8MegY4j78YMEDd7fFgNKWYHULGrYBA569ANrlaUN1nCw9hPDPxygBTWGl803rA14hzdJ
MvEvw+iCB6dE67CR8wOLYfbrHaS0QoTjk7X8yWu4g7tMEFePZ+WvmDyR/n+j+2MjPxLla/d1V1Vk
8+uPhoxoPNI24COs3Bp7ORRfTPG3qOY3qwuqYBpKkONWUVHYNGx/ZeJdP0Ziuz+OQufRhwnuBrzz
7XKDkFN3Thp3Y0j1fyEcB/i9YAzOOzx0z/WLpuqRGmxru8BzCmG4L20oq4q+BMZJTgRI+CQfdAro
yitgg/H3NWO9JSHJK+GFSfo68qAPRZnQlBJn1sQg95bSIK9c01ADFLyEnr59QCXMovXOy/9/DOUk
Zk/5JwnAwpc0iz7oM5Jj5Lgo9PtUd5vUYtZk/Antb8v8JSVKPZ+y19YP/udWjpATIAXKbRMTuFwi
GOR8kPwM91O1QVn8tvLV6yJgDEgwUT2v+k35IPqutFXMsKlcPN8NR76nrF6nDhFDWgrNyjqZRafR
l+UIzs/8IS0gyazxZHDL3yVZ6YiCiJP/21pENAwbN86ocWf0Peaomk8uaTfQwM22fHpt0mG1gZXM
ChW6RDAtW7xglWCYtZlOr87ZGJ1fkFMFQ88w6m7IMRAndxTERP9VIgEA7YlsNnTQwjb1GeWCxmXz
1EhwxH0MaIuPcSqCosNsMsJCb+L8PtDtEfphY7K5C8hrxbbqV0LLEukD7R6QrqYAUOCQsfTJQ2SA
NtPGQYzXkeKAlj6KJfsAShbYn01TPEpMtaRO0ESr4Rnh4lZHEifnxfV+90j4vuBVdOkxuI45T7K4
O+uePnYR+TOVvAACW9XXYv9cyIl/psQdEqxztHUDNGwzHOg4qDX6n33xxqnVvSV/2KWAO2s/nOIw
MAKFXY44M7OLQ34dobk5K06nVlQoIQ3Lc6DadVcXs2z3FRporUbOeWSoYiQpFqUs0C7mK04gnQ7O
9JHNjZDljJgjEr7+m6/AAfmIb9r1qRFVF4YaZMJRlWyCOyjYgGhRAOPqr0RFH+hcfcmhLmFfKjkN
hv4vYQ0aK5PgF7kzzNGzxz6/UMTmy0uCy7uLltzMW9in996lQyLxe/BI/rdfTMGYu3UyACp3SQwZ
e+aqxYT9luT7YGmZWXnpHKFyyAxjgphUPYF17T8D0Z6+XTV6A8tFRQZ8TXLEoTEYEmNEVtWI2ksC
uWu7AzrHNIhCpy6IQ6uyMKYpeddItRlcHs8wyQ0NflcUbBWbpZM45vwE0HI/WRUFBwJVtgynIJXG
EKZa4c3SaMvmpfm8FScOEErFH1KPddWWiSP3S8nFvNTbik1z5Xtt/KkIvKZKlY6c/KHF8YAjnTFa
HaUzE92q0G8Y+whpK87ol2ApIFGLAd9vQIUwrJ4GThStY/S+m/3NKjWTKZ76QFRB0V54q8TOkfh2
PWvnPmmark+MOGGkymxTFnEUQnwurqFMhDAKsEBze7zTxIuweEh9W7N593m+TwR2ZODqjy5WPIqW
aYkMfMzy7vyl20nJ8BaRuVYejf96OzIZ+NKvHwmlgadjHfbMN1hL43jwd2rnZHpZpDZcccab2y4l
lJNLqKjM8l7vZkggMvJbVzbmElEdblgtTJ04Mpo5EUNJbMfgE/kx2E/Cky3/VNjoH1A+wunC+N+N
kog7cFmJf4hxSoEYfptwermB/EcHJbWFVWsq+Zbupghryt+hzSxtn1fHSfrCWPr2jnhBMVhUovSv
5BKBCp4joxstY1igvBIhfWp9d44XG+G8P4dEG8XJhEv0Kw9eTGHvVK7wK9WNqv9NQEuJnN6KU5Em
n6LkA82+zcA4fn6lgIV5YdM90ek1xphqwBtY+HuYemY+jOA+6XYjijY6uRpywhd8OmYJEYMiow9F
G73f5LDzZebhEqRxc79040nK/JcPmsWhk0SyOK68DkpntxIWRvNGAqjBX7UJw1E5T1uJvHp+zokY
TN4gN1WmKy3oIFugoz9mIWBYy4EFC4z2gAgvTCP5eYUV77Ef07Uki3N17AfufXg4dHebWDBTNf3k
kgHbYhILTDiEn7JAvIRhreCcPwHsYyJ+XrCS5f45WkUuju2fozzu+hrhTmqk16wmWXMLarY3Ojyk
/Cc+g8in9+m2hZshBtoeXsA/XV8+qjMsu5jrNFMfOvEX6wGWwCudOTUjgvOLezLzFZFJsXQkPevf
jBGIKhvLWEs2W1NlNChu3NXFn0fKv4/7uUd7M1+0l82wlBF/8Y6x0LxVBeQRYynbcdCkqPyWM4k/
ECZv4HsQYxg0DMXfViQlU7JLnkwcK2a6lLjWananBtmmC3NJpZgPvb4tRXsTImJY4Bnih5qSSkC8
xO8ByaQmxmuYxhTlZtPd1PexbUKlDSF+Ww80/MgiZRIZpGxwG2jrMvwO2atuLF88f2feMIoYWvqX
YqYxvKbYGK0lCEYRaUb9pKLfTziHe+eRRykRLVhda8v2BP+CX4LfeLRUtIsUhoEBhQ9srjz7Fbbq
2XJTppzLe4XgBz7j5xPF82Tma4nuVkVfeshORhcZXQlL+ctN+qt0G87BpmpJJROycD4p2dulsRjr
QTA9ICkrC7VWodcbbVagiBtFy8n4Ao7vSHyMGT46WKW8iWydJECTC27tHBCiA1yCVbUDlnvTH9UP
bszlikW8oMtf5zz5HjujaV8yZvgDClfZVJrI+UihLdYEqyzDbqm/EnftkzXiMvhhhabmgpKSLHuv
dpBqW/FlNL1oThyABbVR9mmXtsvxinYvat5oDBarDg5LzD8AIR6fReTSGK8JYCxnChaQolnbdr9s
8wKFM2puJjhGUmG7uwT37fP+pv4Ro6jMNDfZw98mpD53JVFaSfnp83kK8Pu2taDhrwgnmsZ/7tTV
dTQtDCmJsargkeviS2fBl/5v3zPJc0m5EtBzTb7T9P6pVGaEZZPzf9CFBBXz8rHFRyuPy7mQ4m63
LKxzX5topQRWDe7r+bCmg/tQzyUMaHwKFmBDoEu5J2E2Kldx5LDbfWpXp+L6u+q0b7qTCFLVYrK5
vKGRGG05JhPWl3ok9Kf0SZHvoFm/UlEkBI765qSiyD+Q5nqigdsWvRuadcPbQ7FG2VA+yIU+iqHA
1d8HOC9MBuzBaau4GwMblFc6mLoQ7kp6qDtwWKqq0PLEs5BMEEyeRy8h4dnvjAXkoRZwMJkT0UAr
cxwzv//gvXYiCLDexam/BHHNZjAXMNnzjcO2V9nc9TUwF4Ft2etIexNdysQUGT06XqTmCB51fYOK
370Th9DNarSaTxi8h0kL0oyt3KHbcJ0okkNdkz3g0d6+xxUUMnrzYBUP9ggX4Rwn+bbOQMnmP2qX
d1jdJ6TMVFI+bgxjuP5P8USt7LBp+x+0bWj4aNjQVewVi/Ptphe9OMQORXnYLJ5c+I17OPe4I2Vd
1BIItkbOsCz0rLFIOfET7wq2JI8P6XDp2hbtqu1cLxDAucAgm271HJI8UVEUOTt9jIRCelakR0Hq
sDmOkRajpYlp2LQi5S/9BzVMKI6YMT3tsAgvWAENXsYNvsxCRS8wYKH3Tjpt86SFXFhJ60sTSzLD
flDzhVk1xem0UOcjHzqt0BvmvIZ5UPHA2OU1uD/f4HC1bU6i6viIfws4AmJ+Bd63NdJ3jNC9KNJl
fde3Ntyw7XC+pr/h0nrNkO7cvCiAK/EArV1GsrHxLbzdiZg9LRjye6pe6pDTF6N2qDtsiQGbjMlH
7faMHY8KAILIcJx6do8NEg30VXPw0OWVS0cQMw95vKbjZXL1dinv55aoWtN5+cVIcxqCPf5+dTCE
XQN0V3NQypjc/4jNg/JeONjMr8wcK+HMj/GvpCoIhEymcOovmw/IHynVx4J7tHah/TR/tR7KHsQu
jO7yW+gel1Dvo3p5PkU5fymNKuz2ZNPkT1/A8SbLJco8L97PvDAVWTsfYyvjC/S3mzbspenabY2T
MtJCCJhrGR/YccyIMbsFn1gU6xDLi3do77gvbrXkaI9aoDo8X/uD1+4uRZqKJ6GJ924JQR0FfwEh
AgxhkM+quOadpFOZXhI69yfGXRQLTj8RZP3rCjwgr87cCVFGnUyJd3cgAfdsUN7npk67SzNAf/Cr
osABPnl1eKz8/sGEUZxvbZ4n8fjX1pVkeOHyqNtkqOuCCFITsIOSc4Bo1/+w0OMqUWmXcs0r0l3b
gdXPPwlfzpYbx9O4zkaBac2PH5EK1NeH6SjXsyH1081rVownlOmeLBUecuKIFCRLANRwKPwC58ea
/KiBOu398sSLU7Z01eKSxjUR1OSyKMfvD/dupFvPFNoUHHmKfJWTi7f2UIAjCJp9rI3hXUBPl7sL
fEVi88jJbje5qkQ6AvdFo0N5214rLid6P6bfbXNAHeqbRLnnELX7z4dY/6gVS+1Y1m/OHtECrn4y
4BWUQDERxvCtk4giyhjmHxnbhSmAkvo153iQD8VeUHeO5EK4Ch7KoBqZ9A/DTssLbohdY1eTcFQI
3VsyxOBQzfvRs2MHavcD6cGixqTCKWGGf8o4gNlxrmSYRt/CYjd/zoT0e/7T63VT9U8Jk5sqb9AE
Jy0qeuLzxY7velcKWPakolZUOWW9jkMkYQ2HuiaZQVre+VfCI5ZHKO69YJs/4Kv9VTcoRxC9Xxg+
qraeyM/4fdc9OIQ59irZvyJ4jvL+kS78g4dS2DX7jGfZjMOfJT3ft7/we+Edr+FRNs5iXiszeJC0
YEA2Vko5ewOg6jMXYS0f1HaMIo2RYngpKdj7TN1I9Wh0utkS/VI6U48QQBKcDzUjbme8JVCqyVBp
Dm2VURtdleHwhUKW8ezVHdZyeKw8GntG6wCyQL3ka5ZZqWwSKxOT4soamm/b7wMAZ5kyybajCsnK
Kp+JRsYA07LhfG3zSJZT+WWHS2hFI1aGEn+H88gwI+XowQ98bMW8gBgxWmMTeFq45ILAh7/V9WIH
fsXmq+1p3r9sSg1EYnb9kDrTLxn98rVo420vZgXgodDz+peUH3+mcjjPHG3+WkCwIy71AG8QTT9U
k8vFaIb0giLYu5SAdoQZYVx38w0GQNJOBHCyMOicBeb7xliVmThPvgOm0zMkhmfPKeF3EvANPakf
MwhTN9H0A1KE1Wg5O4Vt/AeL/avsh3ToNeUo8ijBs2AYAPSSomVEGafmq/GRigCMIR+6eYWA7mSW
2x8cndZGwTCyFeJxkCqWtTyS03vm7Z8NjH6cWMakNjHwTupfVG5rgAhxSLkjMdQ++0G4fmelrYEK
/7KsLBtosFvxVGSl7R/2IeB2goN1bZN3be7Kh24vqB6Zi3mdxkmw5jkAUedL2F6WIDhOfZW3B44O
FKhXzFEFhLSnVhZGexLFtq+JAGFUi/apuicINRnHh8DCe9JFqzhtExNjRu0jiHKBfd4WX73Tph3D
zATqlqXyR77pPpXzQYYFtZTKS3OlVtiS3uhDFSKT0gIoU1VMiPb28+djWnmgvLcGpJ2wo/ML2M5P
dwFJUERZo9hBaH0LravREgPiscnhkWheTvYi/mXgE3Dp8jJjN9211Qq+zQDiAkAEga7VFH+CdjsG
Vc2RTPSNI1kGUW7COSUtRrksjOeICJqA4p1rdA5cddFvIxgPxDDxD9vs+cq+2kGvHr7QIErMMRjR
mmr4fu/WXG0HDauNGYOum5H6pak4u/8lURXvTuJ3y75MsL8ZMb4ffW4ZrlnCIoBsIXW8+7rgfW5i
GNyDnU9qtDXAq0lmeAVhWYKT7CdYv81nX/Ci3iSMySGLgnoTtOUN3gogFxHVBrPXaKhEgb164tYm
5L6otnR9t3rOJCK2gBiBfSCdooyPnvMXqhBQ4PSt3ePTytWRpJMGI7r1ZSA6U4bOV09HaGZhlqtd
iG0cyfStKWZ0S8TxThN1O4ZjzmBNDRrGWm0qN62FVvyLZVZ4j7iZw6N0H6+S3e8Qv1LkYlKfMwfd
dYL6AlGquMo/T/1j/G1R+Nk4USKJJa+5u29EpS7sWUNz6HwZH2f5zFJWJ1wc+OFa2aHsd8ZVWy2w
YPRbcUNrQf4RpWRT+jE6CpO4B6QFAhhsktgJLwChJuKqE8PoJoBHgabkQx4d14dsiJTtI/y4wAxc
Z3yc/jGJEfNLKcc7wrP5rQ4ECjvpvcXHw1KBk6iFPPX5MrdSBufQktvbhQDRMdI315TJH33E2Hw4
Nfn1auFCB8dFxbV1riYkTfyi/hTewH7sOXAJ59z5UoQHuJnCn2MbU17B4+gjdQXK1dhrWyHoUAYy
dj85l3MZUi72RMv2UOurZYtFPQbsn6ik27/9Agu+Vh0NxJfkA+VNuzbw642WE80ZciLt2RHEKEmb
PdGZMe0CpIyflA38OKZO5uC6BSysp5ejPu9xNtHEOitcNr4QFyxOMffZWatnGhqt/l6SDO/wwjg5
pkMyIQyAoyC/FST5abWyOnJjUbqBuPbJCo7zxOC5rG0Lhb5HcEZpvZmcPVCSZ/vYdXLF7iafo+xy
iJ792iqjMZa5iNOTEtm83pcWItvm+HNXBBSHXyzQK9z5ALO6TU5weJNeySseo87/Tj3u7PCmq6Pl
pm11RteCQO+6PpoAX/K/sMUZRsv+xhtU40GTIXHzaDq87yDmJ9Qch/8PohmAjZ1/ZodhuW4odu9X
PFjZi702FC65699JdiCXwpCIIUqdxvX6l9PnHNb5LtaaI3TbRxOy5Gn4vmodSG1qj1ZMnhYwEsUM
jmx/n2VZm9BeK3Ukay+/I9+WaOW3G0+fb2qmXw67K5xfv1SYTAJpNFZtdrAI3bZciIYWdnttg3S8
FP2pppDBLxLJ8OqWdDRNiBsBqyrvT09phHu0dbDWqUvDChBnC2cGsTp6gPjiPGmg2wNDBH4bb/th
CbQ6m6w+czPHYhoeoEMCUji2XMU9lAn4cD/Fvzh15jjnASCwODYASiiUznVJ2qqna6x5xWsubbLl
ciORL1qKF+/5bReze7hQcQqC+SYb7OcmsosvKrNx/nKr8b7jFN85RCFKMrWgemye7iv933xH5QPy
a1cEmhRErzgzVoZkFSaVZitLXFg0d0ehN+re0icM29F3uzge5izNbRmMWW7BUq41v35twRI9Iijt
wDMeA2jQTsa19lGuIiCMxtu6MOFa86JiN6r3ttPfkS4Iaox7RUk5VA+D2cPut/ExkFfETM0rgFrZ
b4XmgqaMS0+ifse+mkBC4C9Jtwifm1zlhGlHyEqxWijcH60iGDaBN6LrDSl0k028o4/TQCv2jJHT
B+SuQ23DuhBhBJkY5ElbBAAqHFIlOVosjOtGHwp4ki18qd/A5ZzQNG6TnG7z/LrW6suo16HKLhAV
T5SoDTUruxbhbaXzz+pgU9WsHYLCW8CnVBlFCJ5fpWJuSs93v10hkVW+zP07XoZqYVsXldrky3IX
v7crHDPuL/oWA1GAp9YNneBQUfepWNYC/vUnMF4t8wwMd/khmpxs/vbjb2eKvXLR5PgeyRtaWyCo
OWnEXVHFpPMXnlAABCD49oz3WGm/QSJbYeA2Yt84ECoBBYiiiEH27UEqEg0nvRrYfF7uBQKRfFr7
6EUi59QFZknY3k2g2k32wfRELh8gqMEAei0jx2qN50s1CiL54iAtG/ptBOEJqXBFVs7p5s36MGnq
X8zKFEV5bO8rNPfyduC3m5ogF7+48gZ6ivmX/wJAE/nXhVe4+Shnw6jIKMLzGIl3QGXcn2t0wg5t
hxizpFjZomq0dm79m1fNi/MqMtWlasr3/mh/JveBICGc+wumzjdoKqAVGk7klXUW8vPxAgUR6oLu
+XB6oteB16uGCCvZosfcwLgEolGEG7IQ1bNFe9V8yEWp9Mxo6+7EPJarhX89MK/sXQLQ2MSXSAsg
1gC8dZLhSKBu0W2jLiXQw4tWK2J5wTKOKQkPUrqZ2hJumQaA4VfZwk9uHT+WvhC9EH8DqOFxIO93
u10YqWeB8xv6dAVrLv9cYx7b9enknZr/vOC68NGiEgJieyhEkNlUsRGzLP1GyXQ6xJDQ3cExIcBX
Yk+z3KZWmbq1aas/x9z2OWJ5b6WYCOLt96SdgVn6EO7aSB0PWL65OPGpxJ6QRHubX+QRXdnSnXgh
oRDWSbrkYPPKSXclBDAeAWRO5b7xOZ8cjfE+GahfMGpB810sVOeNnoN0IspaRDHzJQjvPiXwDVZn
5uu5vCbrOOho8TaP0ivUWqGJ+3UPKqsL9IMLaWgR/3HmaNOMuafYNInityIyzQitZcrClF0Qcg6x
hc2CXMC9u2fzSkQOs7JiUDU3pilgImiFU7hE40yc31O5HYoODnDf8kwaQT05ZrZPbCkv61lLihci
OXOKTArV2TJD0uBj0rRqnYCeFTrNRa6pABKI3P8shcJkhFqQHSycNEUOkNaDeYc2Sd6I7Zqoro4E
QwazKxGIFi+xj3XtTGZucTf/YV5oDw7wOrVsa6M3eNY6uBSsiMsMOD67DTdJDjdgF/PSxBQUaCvr
DSk3v8XYbj4HsPE1vgGdYXcATPVYhcMxeIm9L6eqCfWfITvR0WRZl1IjgyimIRh2xtuJp1ab8XId
aifVKxubXOGSivFRT5PD9yzeXbSDZm1qdKEI+Q2AucedxxAu78gGeswAnaW18OqjIgSzw0x4hben
k/rLQJrW3mLxTRhdHvTzDy5xCGMpkRyHbw4PgbvYK+vlSfaqbEhIjxclCXQ2a0bb9XArgAmJ8IZz
rtrmD8nAlFT/IscUU+mG8aE1BhUCt4LSABoKW/WfxEZ/F2c+ytOzVln2ZhbZufn8yuP1cY61v1tq
CeH+iUEt68VC4inxAfpomqS3olPI8nzdB0uhuGJjrx3udvTaZbgPRIUikzKBsP1GXd7inKlBUP6X
Ui/g2AHNNO19NP3iPsh3mi0aNKDN75309t976+tq0cFH7Gi/+4j41EEQMOqvKBE7Aq4GxvSjeh2f
vCext+SnF2ZiXkmEnqHQaLcRhVyaoPfXUla+iPkIzaf5EMCACU3uRT3KbFkUqoB8u9Ie4WHyckIw
KuBUwjA9m9bgdRvLsmqpgdCkBZLqWwhYDaUSp2WaGx8zWQLReO/9cnn3WUCHTtCh7OlviR+w/2jV
LL8EzNgYqVtKb81eubS+psMrPsnP7Mku0cB+pDPMu+838c5jIEWNSTSjW0AQggL8CPMlyFsfq/3U
FI1/IJFDmDTExa1Twk+yl2u/IisFurY8x9QBXPW2KmlbtivCTZ41bWEGBEN9tAUQVfoNYEV81eiM
cciLB/kYcfaUB/afVndpXLzXohD4JjTj+EC9E9V+XNTg0ENHLlSJvb8ltzAV+Q/oyBgEgox4ws+q
ovoA+SC5PsI1QAeoHi4q1/sOltSCyrCXMwNm5mMd19zkHtW4PxM1qST+53mIFaQajx3fUbX+goy/
7+ew7i/x2rNi7MPTUmL3TPJAK/OsFZt9CWKBOndBT2zCKTIbsOTX0sJSTFYw7vJkozVhX+vFOzLM
VpRBkolt2WKbSK4ndSZcLlNH2UWxH8DQHifr92ZA29oy2SD9HLHpgVcyQdZtPYrmqMVOqC6rkUU9
AsKtIDxewcDWYWSr7ZYsR12nP1i9OUhtRqO6oDpMNRFKDKTiheFwzOdopScjeCJbu8OuKnpOEZDa
8iELPUA86u6t2guAMd/kIuUfZc+SsT4EfKYtcDzYOdiOhkkGuE2PUnwuRlPd3xplwLxNmRENxhvA
UgeJeQCNafk/yuPLC4AaVuCtIq9E5Kw615YXmQCzzPakey9Eica3JhD0blBONnyoAEZSzU9iJ5eN
Ufhlpn/JaIP+lwnb7Xj4HaMYnSm0unj8bRTWikIRM3IduZALufqJiUquUKuykVjUVEwvhX1EK3cw
Yqo/wQK28Dt+69JsMF8TOFVsi1rIUc4Q8NOO9S74ta6CYJ7Cnfn+Psd/bYd9EZnd9MI6+kkfZw8y
saARRCooGCpo/3czhDKTRatJ2xXqQ2yr1dB3dXeOz2K6P8pG/g+ssAEOW0wWPpgUtlZnOvUuiAN0
LtfHpnLVr5G6Iq1gFRRx0MRq+wh/XU0UAtfn46SkZ9m4Kh5wVm6OuF09GKgyUWxuK5I707Te4hdb
hr8lFwBp8Lzz4F+TT/zWgwvff8Wv8aSfVJgYYBpfNvxuwYOymac/zOSiqaeFrK7JWr0lnpM+OpiK
KIqmiiyZcKJiKMzGUOeDr9h7RcnsTEsmtpuYhw01Fxa82O4YAZBJ/369r/o1D00S1SXPBNG/avTX
qdofIvOMUjmeL+kkeucMuGC9zheYxXpE+DII/2W8PoM4yLvR8c7+6QTGKTstoCDhJTlhqUKGLi0i
A1vjPUGdvxzSgMBZIY3dvBWqWmFQEI8bgYQOXge5Z8avlxG3MBFgLNqliTa/ZBnd+8GLRW5zPNNQ
HOBuAa4bNrjTsLoh+DQQN0e6r+3hYDXt0feEKx0kGABc6fJ9Q725F0BUKapU9idxt5vQp5XHvEV3
GL3HoJG1pyjvnL22DQMx9gjEkrAlEMQbK58KoKHd/Ozxg2C1f4I4vCnOsR5t6Trpe/oZIcg6unzj
6T7E6i8/fLwooh/9XW5hHDCAYMe+UZc+mFfgfRibFKTGR6VWboGkHiABCmlvOXhrX8Ka0qgn0sP4
SxXR2vk3CArry06qNOGDCC5Fm/GngK51h29E+ECHVGgWlyKT0JpR6mLIkCOoTGrxZ1sC3Mlm0RNI
J9zVee33bO6vUfdB5PFwlxNwZfX/Z3J4Fy89dmN82RHnMCIOq/qXt0S+IcCQElbdAA6P8SpxXvUM
ttXI71mDhSM+aWIwvQWjemP+BR/OkwzYLF8lQaJSFZeskJ97g8infOuvihuDckN2+YIH9HBBwsVS
/w8amtuAvruOD1WMR416AIQ6Q+Ei9COxdGsTupW+HPOo86OGs2e6/67Zu+Fyag3PrrMnGE5lXAYG
WdLN6mUdsC+2C+vGmwIkgLqccq8TpT/2B/b6xlNDgCb5gubIBWXJL05NQyWo4SMi+3Mz0FxFRZgb
rmPcsQu3eW7PruOV9gOMGj71zoZjh7AExs6a1veRNrm13ylOECdVgl0XGKvvdpbjV6rQ0737RHnA
22xtQkIyb1vF4eVfIvD0qboESsK+r1tEjsdmLTd8yjEZ8Op11ImewgkpBwklt2RXzw64W+GZjGox
sqCJqLxw+TW5Pl9Lk3tdXrXW3j+jDMw+pQCO1IbkZEKgGFMQXNQ3dFTX/MtLE4XSF7+i+jZOQKC4
ah0w3QPmylBbGg4cWX10qygrd5bY7NVqjhxXV6/3IdNdscqY4BAZg6Fx9TNO7Jmhz9LlwBGdrL8I
DQO/7+ZwDsonMYFsxPAeKOX+Ag92Y8hOwdKAyt/MhnsAZIeEumA6nZT9YlEk+5snCNSaFaMgJzsC
wUyhz0vpCM7KmH++GFks/dw4Qx78vHI3iOgn0X9FWnUB399uAYo1gDb2ihDYzDSYYBB59ytQwofw
CO2NHc8tGa4IhbjSEXrb0QoSvKgpBhkAW4NMbDhu4Kn9KX+3Ky4Nvzw3gkTevOlq/9PPzuU1nd4R
SUM6GPOjsvF9L2GaGI84/F3v5JHiDgXKozixkMnhAILARWem/iywqldhkyMi3BFqGpRsrmG3ln9v
M8PXb7UYk5Kltaz/rgjQ35BrDaeWq1l4zk8vdJKQF3O5JUdEFAN5sKiFCz3xbIitqG5qSp5B9ZrB
hzVZiK5JoOnPF9sTIldw6tZK/vKIVBrtZFn3oQrzh/0tDnTgTmGF9vutGvr4nRNn1ahGw2qYsVRy
onvR34743In4XcAycKqPSQqbKR0NDEjFQT1CUabQ8GqGiIzmkiJrCTyPPKztr0sZn+HwGyqykNIR
64bBkDD06W4A3kR1f8OdCB7ifz8w2xJ0qwZMNzAEZePBK8JAkdZJSLMvYOqgniQ/Fs5/Zy5VmFr2
+jdzcd83aNzYR9vYTVh8C6IQWD4QOosXNjqCZHN0rO4VA2/7k9YMmSD4fIB8jaYv+wud/OoWyJNX
Avd4Pkvr5Ix7Dkn4zm6ZcPRCEJkLhja7/YkdyV2NSeTa9GSlP31QOoopCuSzIa3amQGYSJu6wYaQ
3DYp4x0ysXJHZ5D3qgeMJscrdIGZ0caSv25wAnEwh46WjzFOK0MyvEqutElj+7ei5Sx8SJLduI1u
tU4IA2lKXSiB/lK4SS8DBHHCDbF0gSS7C+lezt5/o1o3AWXRYS07ytAXK1yIQ/MwdfztxVmP9Gg0
fhrcE/1yCK8AsQm7d53w2ARrIe5XQMWR5TX/x8w4Popd08+ENWHxnVgaT0D+feduyD6ivquVw3H5
ofpvJIxu5SCQj9bZ62vll5IKz8II1dLZlDA1j0xpJ9ZyF67SAXJDfXMz3WhjVb5FEgZIc3oz+PMd
3K5Aw5iu87azbW/Mf9q6ZyF+07alTEHF+A5Z7pw/5TD/sBF/GmueHZbs9+KAuKDGfbqE2mA3wvew
jzhhCtbRl8453bUTBhXD80KAz1vDR32H5MRl/EO+xwJ/+3JZzJ4G3Rsd9xmr2UYEWzCMaOGuzuum
+hAU1HnKxGGlzuq6n11kYf1dRTWvBAUaZ5BsuykhBBJ94Erbqph3NRP9NhCbFFeBCBw0pqNHx+im
OT+V+s0WhRss9LgnnuMHqORZjhM2GM0j/m6fWNTA2CwzMjscbD/13QScCTZyYyvT/uDBrNA6q767
w8pvVrduDp1m5SFvmnYvREiMAXCj0gz7kxeZ8q4jRHfposv0MClH2GGHmoQulurbY2S+RpTSaDXR
S35Cp4GZbs20KiCSv9igpkQaCKeOJWiBWz6FOJJnWwPvnse+jfJrNMiUatJxVGiqqGIPDQUBf729
KzWmslYDanhG9R//gkIaX6EMEPWDIyokuit9zmDrgw1obfBjbuvkS+czZLakJGmPp21nhywNTRc0
C8m+FFdMOSJXt89UYJOsfIjT5b4HBy2D3bc4bQycXRqB5tlidAwUSL1RgeYgVPwQqmCITA7/gtkN
Muef2qo1qzyyaKRl9F8Dnq5WM1BrErNviMmK2dS400zti5qvxvPcN123zc8mJ5g5uItrLKJaxz1r
8bGvI1DAy1J1pZkKDRS9ER9/e0OFv6sYL+Qwcj/6u2lych8XB5MJCh0GUwk6mUd4xID/ewOeZF2/
S3DYYQCeN+3q2OYFVWw+Cw42eZwZiZO3yivC5CQuZ8SXyuzajaeLE3zmvDBrp84qrITWOahoRdIQ
xf9lDjcqj2swEzUtjElF3LfLPn+sfQvGQ5v6zO7xNirBZtCM8T8/E2FzaVntU7nHDqkteE2o5v61
UHAMdvgv3gVQwNOcL+eEWSSm1IEckN6jZtdfxpi+eBruMNY3+IBlqx7VshmiS8PAmjwC0cZhhd5n
4pn35Qv7O75XPmqfJDIoN7chIoReIA6gSFZfqpRxBPUXzNstQqyval9GO4LaejS9LlQXOw1e2Qty
MAvc/GyIYKPwxHj37ct666N0dJmphb7dZ646lQcqCnVFtJpc2vzTniskuBlgK6v3X4KUZSEu8YoB
M0yUUdDm8v/v1o2LS+uJdbBLp/nz7ZXMeZoHcjtxqilaYx9fj53Io3jGMSWcjZi89BOv/JM0q4Lj
eN0EBlZ+Rrx/hd68vvrl3I69xamTNUt17Ga/MR5/dbK58T9rRMKToZ1rFKLU8pui90hQp9ntXoSU
T+S1AE2S6ghAyD74q+vnQ6TZCHPRZGeXTlnQw0CnrzltoAjKKhoc2mudAE4AfTlb/odjZUDWSDEf
6O4y5Dh093CY8dfHM85pGGJ0XVsDztdZwdJ2ERa6vpRwpbE0tXCPEo8xtwBZJpuq8Lofi+K1K+Sf
cvKvQ2q2UjSGHQmOlhOMpOaI8569puad7EG/MesKqiHBT0ZqWtu1ODFQgyBqKZMb2WEzI+GcfzeC
daWQCyQJFNn/LhO9lxOEmt9vgOmdJgE2srwDGntsjJxZaLmJzSWLVvrAA8xt/CxYnMDKJu44Ityt
Wl7k0TB4r/zYLmh424zJB2XI7e/ek4wTOqeqof0jwtyXRxQ5TnQUzEffcm6MElqU4K5NhkcyT+U/
zqCSxfBSZae6/3yaa7/+wkQeoYjPm37Pj2fcnk+vlzl63htOMQ+qh4lUYn4Q4TD9jwkMfOW1u5Ln
bvXVd4OF96W3aTgnV59slcmUVF6wk6YUQy3MvnC3EKYMYgBrQfB1qgbopUKqN5UQV4JmbS47O7ns
nzXAsGsv8c73ge3xjC24gsyoBnLocvPHmI9KiUksPAJVcIMAUNCTUTbVpnGVyzSqQ6tR6ZahAUPL
uKsBYlU1E1MawVO8MwhKd0nurqIZ0NxRYcWI2hQy8tzato/PKM4KqR1cftuMWmYPttzQFGS45sl2
hLMPDRsTyCm/wz66pqa53x7flX8V4Yn/TTfaB6uOmUl6wMZFhycja2YgBh/vQxepm0jUePa5Bipo
cQTzaANPsP3HmTjYzvBkwCLJFL+NKh4igHNx0m+g45Mui1Cdx3Tgg8XstPg7GraD5PhTBD8UKDYc
xHGQvhoZSq7JGd2mgU4+uZE5hGM6x8G6vKaLg88flZ48NDtbSy+eKRQnI9txcxM9MiuFcXKi16SU
5L+8f/nFsU4Cp2FN9nc9MT00jSQiFCtMJ20/ogJJLkjDk/RLlSc8GcJOs7YzNo//aS+02AlHpZZO
keAOIvhlunfWI1/QiVJYLIHVSrT1bg/+OhUuyNbfoX6x549/Ape4OjC99bTlHXbc4iYOODKHzL8Z
dcYY268PL3K55ZZX9HP1wUCNX6C0oRCjgcJ3+QAIuHk+TgJOE+IoFDx6chV1xsZjgzWC1GlPj8Tp
Q6WfGbn9FOOA3ROfzj8+KwATJm1l+KoB4b1ZCA/fgJIxomBkPKjFC9Mtd3K+aR0a8KncBMz71BuK
QN5RZyiIHtv2dcZ+jJWhib+DmGjR974klvA5qYJad4wPDdl9orioRSYwq7/i/qQiEPGC/1DjWqZe
t9WzsLWkk5rshyIFXIaSBNYZKQn9dJB2S/dPADK5J1XmH5H/uFFHUGmJVozuoI1sakEFfmDN35na
/HaV/f9AY2HMYtqul2Xv9wgmx0/vPDOWslduGPNtgMRC5teA0F7YaFsdDb2HLb+9M5zCBz3DMvXo
Ej3XkUUTkJHuoNiw0HXXalto4BL/TrUXqbxIfglc8/ErOiimmqvWfIRMu01SNszYIY8VCV23dHhM
P8Hbt3Pw9aoG8hudadCVb6qMF/DmxOHy+GszMwesF4g4LMIAdUsaKKX53+TWN9ZbSxBkj8sx9Y9W
QNlRPUiEGLNRZKYo4W+X3zMSeBRyS55qlAausdB8J/X3YI/tZFD+cdh/gRW3ebq7soOS90p9xX4U
gU3NNAaqWgBlA6hitHMSwcfRnizHUKg+v7SiRXrbwJ1oVsPQlvsghYqwBodvw9EksLOna/n194BZ
uVLU95wvx7zIToFG7dtGC3XI5vgJX6VWyUwVLOWFP+NRyIM87RjiCuha6L5gYP0+jlcVBQFlpuZ2
f/j8TJE1j1UmhGqL9Xyj/386AZxtA75ASSNT35PuGS1BPM8eakYvuEbhjIkknWAMwN5LQhUQjCmJ
FpOgvHJbm90ojaNLo2UVGt7qLjQ2ugL34QmRA/u31cFtuHC6LUWQQ3gSTJT+7rAMg+wreTUFQ6RY
RyZEwYNbnUaZhH2//nQj2oHdjLKxfH33TmnzGK1lwW+6vF8QKd24q1XiGq5zsXNK6Kq2H2CLheoc
LNLgu1I9isQpB3o8tx3V9OwOMRI+TQadI9BU4/9PUUl5v0FdvkfIPxVZ8YEa4zOJUz3Vi1ZQlI9a
Z1/QCWgwV4tCbjmn6MMyi0yNY+19UIsO7FCWJCrMS2qOFfAEIbnF0Vt84wzcuIgrewDkqSVrzDQS
DVvA8uM/4pxQddlw85nn8E0AlCE+zcJuTXgcXqomYUQdTy+HuWQhjHoOWD2h/nFUug75hyinY6EG
+b2hdrKqSZcZe5lj12YYUg6ly8H+qPuEwXvWuOwYcJzc/l+EkPlRcafqGxjDEt6+uEeYzg59RYBe
qoBPDdPYoZ9azrX7XEo60iJNnkF2UF5DTXBPEovMxC68taA/HXdozk2dbGhxA0zHBzl34RI7UFY/
KKLcY6Pr1SYz3jBNG3dYgwuSIHx/EB97ja/eg60ieh3YKLZ1i8/TQYEE2/8bh4CCrwz3vewdLBeQ
YixlH1JDEp8xylDi3n7yf+Gr7gFmep1I6dHlmMavmS9K5lDv1IrY9W12iW0WobAZyHk10PuV+9YR
8XvZDPpqdyJfzxdoDGfm4saaU4G2oCJ/UPZq0d4kATDJ6wk9Iw/9t/sH7UF/YaFM9J4RvuwlhoQ9
i3Jx4KDbBFKPkzNOjdjD38L6CqIZU8Bg51yU/CmAZgRVBfZhoeI/aLACKU0t91zlXxsdKnW4JqB6
3T4/Rc54vLRHq/ggqp4yy5G5aA7JYVIPlVLyZOEBYy2NTUAtiP8Z+4ukSn7dSj/1ttb7oUVEmDoA
MdW2Z+4gg9ofyOevJPlWYpl1xx2+F5TS7Hjl7NWfU2pbotOxrO6yxhpctZsc6X0VndgPRmAK25d2
k8O85zX5DbfZcKwFPm02iVWJoERsTLPDJ2on71x01062kQeUU4bW061ICRkn5zEe/iE7QHJPpUrX
QpFvGmmJ+c1+6ObFbITlvuPfetjR8c8kWJTfDYBuQ1YWrkeZ2RYVp/9owYdiY+5S1UgM/5iTzJEi
mtZ15OhdOChbl4QgHKKRL47iqZY0qp3CplvC4s1PCh8zYQAusF8oTHd0+BfGCnLmb3xg9KMj2NrO
Hr+GruS+9ANdqS8/kCBX9CFS8uJrY00w+gTg6L7qJ0nkdgtJYqLMwxPMHHxmbgP9Gj1n1DmBFlir
9GZh+Z0Wwsd5Ir9ABlgxVhHQcYyz8p4KwfooNGf4T1+/7kZ3ertWxyuM0oVjhVWkfY/x+t4bYFlo
egbTEEzlpfo1XpzH34gV28LnCBcliuwWT+S5Mi6dZ8pWIL8Dg7gTlMSstRPmiaSRqq+7kxgsTVeh
Xkr2BFKLbIBKlbeLAE1JLq+5pSWiW0EyWr57V5b2yLgUdReXRKDTwmerdg6wIZz0Rpk4myyCCYID
liXhqgu2J+jgXSiTAEfBakiUPEP5gqMKPpFPAurbA7Y3vZzuSzbTqik9FqZXpbzRe1sVN5KQoJ8/
PC+HnnaCCt0VD5aHw5PHKXakK4yVubWNkNzzf/lxmVRRvGOdOBkH4NedBcluyF2dsJAEarvtbedy
FeQgQy7fHzLPxjXSSUcn3VJhfnKdhKM7y9La8A1LjWIikEU+xSViLv9CC9WCLpOcd94G9wj+UM/p
qIZp1NKVPCgf8VjLSsGI5zhC7rKm7judRtGyH9NoGxkDeBAhXH7FwQwQG1EMspE2nrLMep6+8ol2
L+yfFhpJFIRu+NF/VBbBvbr8ZRIIqbMf9P97VroxalLKQqcukJQtw52daoBVBPI37fdvHqmlR7AC
2BAkOUuatRNmqz7asvr6PrphvdLz6UU/Qn+X6oPoKbC6V0Wp2kkLsdmtAKIJ5VzZshj8nV+eUUd7
BXwEBkaFX7BB9PuiO0ZjnAjLEGCQDzNI/9C1t28s+SFR+r8kmVKjILUfoo4oHEh+cB7vUXyu9l2K
UbJQr1pvyUOwEvA7VDiX0Eb63YY9PJZy6L+WmL6dFMyF8ipg0NMAqIKEr0fRxT+M6acaoxsnNxvR
s1zyBSLq+kK2Bws8Incl5y9HCPysA/fBb4XUa6zRFjKXMUcEBh5EsLgLECzwpXgFwF+zHBflfdMo
rltpycoXGJC37PRo2UbuZNVwLT16h5FmNLJhxu50d/1rvCJ6RX27V5tRWmzeYx70EMXRjZPsN1LN
KaCHnI2/YdIQqzKQsxAG/qeWVGl1vLi3mVII/TYGXiqDNvO7CCSGAdNOjZmUYXTnK5s8W1Pdh/XU
aB/fVLySBreF5VyOirQ/yyNtx3NAyqvUnqyDEjWOQXufwoJXq4483qdVXScocRVGE5RolQ+UdoMm
0VykkUClxtcJz4ODbdQ4orQNj/39xf8Zyw65cuMBU2Ba6C0Eq+bG/gkZDAVoaNgazD88cnLg851M
G2sBwqA3DQGNee/yqZhwoYdB0H4C9nLZRbwIIr3HVhE33meLG4XPGFWZOg13oa7JnMrqMEocYC1g
iLWbd1IrMqTqzE0euyEdVGiLTJAHx9Bx7q+0OECh7oyvuOxGhBJgUhh5zrcCKaEOcnHRhcE7QH0y
sgMSk7cYHqyMVahzvR9s2fM3qlW8/fEgM+ZmLZnPH1ryLRpwjHNBqyQ7mR6IESB3MmT1hViDiyZ3
8AQ7+jWU0RZoOzb5JlBm0eEM3BrIrxBVxDJ4dBFcJVfikG8EkT5xi9P0hhoMLtY/X1maFooiYqNz
4XmM/NIQQfv0Kwx6uDjw7HtTVriuQ8wUBBZPznXxEJZNkqyoFomJEHWg33bWIkcuH3gAeUYxlGMz
ma0T1lcZENSQ+WVZWvw7mBOOixY3Wks9OoC75l/4HmBhoiA8dsb7qbHnhHX0722UOSxdhcVcoVi0
H2x9JTjK9SmIhk6mCfWaGtna20fVM/IeBB1q3FtHFQUQ34OWLaNgLyVPm4iq4lHVHfuhXKEtwR1W
WdgqDWovtpJ7GhloaKpJ9xMmV6IfdlRAWp239pa7TYm97ewOEqex99nbrkOKBa5CJSGWNXBlN7z6
c5sm9ldPm2lUZEyXsYiFMGwfBm7pvsdHlkbuQ6SJURh21R385lah12A3AXhWQo5GtgMgbZACLb9M
kNJtHR5xj1qetLfTMzY6xqMfuoA7nu6aERnuUon9P3Q/OC/G4zk0nEnEc+PJYc0EstODdo5hNNsF
7/at705tEFAxBXLLI+lzT9JWPcOmv5Lo0rUBo+hV+gzl5XVuq0f4XvdtdgRCh9+tJ1Y++e4x3rJu
K6+rFxs+xS1GVuZy1pQW6KpqNJmFHw8ciIjYyBXeI3ntsZzR9vXdSVUXOaN/Z5Tr/+QRN5Y4FxE/
5x/W8Alyt0rQz/l3nG/DoWelp61dcy9a0zah8yOi2iz7loAZb2jVonmMnq+MVAMhklJ49wvHMuqS
C/qVL4ORtrkgU1WkdxN9KPD+aYHDiAiJN1oLqTamdWh4v0O8pu/Zd81Byq3FDhMih9hCOefifdpm
SlLKd3iTq75WfLXXFKwhASVX7NGQK/h5UKwirrXBX/Alg8f8iBCgLmWN8Bh9dQ8lVA+MoG2nXBSK
mBREOPSob9x+nXATAs+cfErtXpHNy/JERJ3PTWfUkgxalBVSG/AYloLwW5EJE82atPwcOrH+FvyQ
OS2vwZWyu/Ri7qFnIQ9v5+Hv2uU1e0iAlaM+SKDhjay4xFMee6xQD+C/IKPEWhRhMqg5x4lElXRZ
Tu3kGPqeINxWC4BPyc5Uxkb6ugi02IQtqScKzzrRjU6fh1sXRgPIRGm9bw4DQQKc3Wae7PRrWvRL
6fjAzQ6QgqgULeZZo0M+Ye+qntQgwDlcCGlBnfiOS6BJX5XjDY46HbOjzSDjMsr2OMIqvaMGnP6I
ny85C+j2wUVr2rytTpk4CItKJus4VHlgcRWYElaUjdnLtzsRG1y+OXh5wYuOznCEJM4J4oYrk1rk
qMajd0GtTFRskoaoF2oj9JJhuIBg1nVZASd4RqfKqdKaXmK/Yw06QxppYOHv2qLruEYA2AqYnjuj
VSo2+zRmncpRHGaRsjYWFK0UVe4edk6IJyPLC/HrrwU1R6E+ndVWC+H3+inbIUQaBDnFq3YInUun
DLMDsoL8UzAApSqA2VlSTVFQb+psQsxBNWYYItmwk6eTTeYHD6EDu2tk8PScE7tE+jIHfOBsd+gr
2lIO2qq9lCdc29yRZBh6vdGZtflUB25FrKD1WibL7j+DP+9wGng405ZbFj5HGN+Rr8z0iG/TghM6
9RDvjej8SawXWF41Tv8SNd7mw+5wL3ND69M8Jbm7mAZKAq/I7NWzg8BYXq0zw5EEwG6M/RNrXbTh
65bcTCLIrzcX841KQsCml1f26OKZsyRtiPNY1ELsagR2as8iWe/0jCgDedd5qapjX6YmRyDQYXDL
uWDOEhp981020bZZHEee4WCWAzpuF016dudIf3oPYSNcQjWsy2NXU0evqEchJrPUREXSNYH1grC8
kvqDRS8QODtoHjrpoNoX42YwS60jYOEtTjb4RLnH8q2mM47Mm5V1iUozOb6EUYQN6pA/WxV7pGay
ADNfd2pU8F5WCgn+UuLuUKXiIhzOm7aIWjmjmn6MMitiBNtZRy5QpYAzhoDErGVeRUvwixATebmP
cfvhOmnIPUsNskV0q8+YHDvqogDS5DEX5QlhJx+3fQNrDcfIrJuZ/X+dwHFac9SXIgB12PvZt+KO
ZOHk5LtMX/RdfrmW2EMoLt1MG+J/bSTdBcRK43jMB/kTZyCZZSVgGqEOIfjopEzTG/ep18HHc/eC
725uGypDztzwGMVJTv8kzDB44P3UA8VEJcUHzrgv+Rt6BiQDcZKOrsIw+uLMkVxP71VXwTBm95S1
lIJJ0dXKXVYYVpMQB3FGk8gx0OHS1vc31JQCQy9uS/d+a+VPt2DvHDnMYDftB4Ryjd2ysRGTEktP
z8BUoKy3lY9Na7rltK5J7m+Zt+HXJFZKtMDEAviAvvfSkumOJkalMEQfwMvUp7N+Huw+zh0/lPqe
dW4iHI580dnvos2n1V2dX8C+AGzg9XyJ4AGvx0h/CLZEDyBX02tbDqBkoFDPu2JxI3qrIrTswAfU
ETgk1NTcLFh1eyLnVaD/DfZ2Ou+nhTjDlI8VmG6CR0N0qayPEdcQoemar0b/KpTRuE1PHVbe2RLi
1Tq1uQ/4t8o/s2xg49dXF9HVntutpLd+Qjx7K5EKIS6uR/qU4EP5E8kukWqsICE0YrgvZxV4SYzV
TCHfk7HbqZICSaQG6QAT9CQFO+bpLU4dfRnYhrox5hlLo9YRA2Y3H6eMab22cLOJSZX21hkbuw/k
XrGQcOX64v8b2d05rnrP6Spp6/6SPjIwMFHiXPNQ1Zpo//72RZxfssAhaqmAFs17DyGQwjIL7kl+
yfo828p7+LWyt/JinpcuCX7/J/ek3ti+QU5BiOr9TFUQw3v+WOoiuUTv3Q2VDvSK4kd6B/TCUW3C
KX56GCzC5x4SjUyS09H9GgcTFbJM/brQejf3uAeOyPhL4XXV0R2G8YYgSzZ2c5I4J/kOKBzSf/wz
GBT/I5yKYTbLlSaC6WZoOj5l21dWX/sEHTAMv9uErnVZxD/ctTYK+0LQzNPx7NaEaTuujiGNjjwM
1MfdSTm5R98W8M5KW5D38FJ3TrfkhnVo2zmep3RQY/xSqw2dHhMGjZu6ZcFoIGsPYqrQ12sP+TJX
SQjGw61UZM0Tm2yURRpJh2ZtYaJUbCuiFJQ2X6+2IqT3sfxXoIrDMaYRfhOTA9sg0vWCT/si+DPH
gB27EyrFcXdHWywhoIKDFqp0/ENENHVlt0QrfGFR1DePaD9Cvb1eH4dU8V/ApCDhGIT/tl+vvQ9d
sjaP1cPQvfBG6/0UjwGcdZ6OoqssK3yRmZo6bk4wgRZR7kv1k43V1eWIzanbdNianxF8AYaB4N0I
MsusV0vOhJfL3t2F74qqU5K1zPSq/JW2VCLZalRtPDMjDdTyDNuxkjwdpdNNngghrNnlKELROT+V
jPwoczZzS3n4rDMryn3bx5wcCW1Q/ZTZT1/YZRAWdTcUd0/dd3m6P7NwUdKpK8Us1mSOIZDokaJ9
kgGTzO7l523BrIqh7Bqowc7SSoZENtJMXKbJIrMkDbFKM6zq+yNBb9hsylksBxjtj7EZU+brkYyb
NRtMypNEVTC/xBI1GQfwo9d8hnAcZYK9tk+vCoUZhtNALu4zOsuKOzR3UPTLPF8cfi9/1FMbrMMB
dvEJtuxWbtXbE7q1pnGGyJRsuAQXrOXGb8KD94lxypX8mNSvz3CgLF808ISso8qaI2FrgAREBF2I
0PW3FoP7dqAI76uSH/iG6qqsq1iv+YpT9oI3Oo52cE6hEeb42/i8XfwZ40+bfiERWbyi/rNEzad8
Ewg4xLZpAGuMs+oB1ySYPJFQKSFLF+mBl7kAJ/7Gx7chkEME7Lu5lptIZ+/DDEIVFYe24QMibQmn
zZ4rS1RvdrUrkANNXjxU7KkaBQoFvtGKea8HVQMHuPK3ah9W5i54vNKZY2CEde63gTQbAagcmIGj
h97w4K5o76r/NUFN5bjenU9FIucrajHR2qd/+FUKdeRpnsSIvGE1djBbSPNqMVKVBfRMt0ueNmyZ
YuD7+L9wLjEBcDp2Y2fBQvzjRSPBx0Hi3/hG7ov3plRuowMX2ca8hKLK07n+Ctyp0zcBbQyd0l/z
JcIGUozEMpPMxoHMzwYJ1UJrZg98Cd7uDGrvZl1oe9xxEEb5Fw2itCBkUMQmNA473TIPC5sX0f/W
TtZ3Yk3XiAjC4BPCcaA679V3wtp5P2re3pLXvRercQaRATmYelGrg1VLYRnGtWCspVnqpSxkN6mW
B/2CNppzyJAb8d2CTrvqjZCtpTiK84G/64z7vAQsnSnTJuSmK9iUWqbapbdrvQ4cpSmcKKw9JlIE
PHYMVTxIOaV0vsYGPKza8pbSEKudxmArI2OIga4PbH/ZZAfkkPC+YzZ0MT/FJSUk60+zCq72RH0g
8nBnFiOppJZvvSU5tdH6yJFKJSKrxO6md2OGxSEm7+xBabpne2BwVWvjmzfhshvk4SYEm+ma7LJH
ImauJYr+lpHymGLRXEGCoOD/xre+D5rLo6uu4rZ+M/bdaldtEX/wtrIMKAOQ9zahPpB063V8YZUz
qTs5+SEXAcbUo5yizyi+hWB3Syu68Li1likubndG01Q+oKL017H3/R8lpCbHXsO4ELZNrxYWffqX
+D2inR5uB/DPpOuqjFPcDJReUdCWCH3ob+YLphBv03TzLn+iAu+LF5vSt7aWOIxY/YLvlbbaLMhV
oidqUS/GQF2ZawZEpoHtj8PenNr/EJFzPUiDFUvbvVXwAuFa8FvI/EfYxmH3ar3aWheeJ8mwXHs0
qRGzBi4yJ5+vEkLiyO4tgfr3UpNhoGacnB75Fuy1u4KzOeuN2TmaAjCVD7usPt2LAMDtw2AnnNbU
76zVvSEa55E6moAahxwuzkD2E/n97TqWwWT994JvDl6XND+TWmUCss5Ohos1SW7GkJ3OeUCC6haD
LhvQJIoQNRtngoqwlkY1khuglGtveXz0H3zMOagCzcujEnYjWqyEXJ03sbSMXYFu3UqhJWunAazK
PIz5wYlKzzUDMzHrQ2gdV12/8lHOFIzratnLbMzqKSJNIrGlRUun7EGOii9+WloWflgPuWNjZmiO
70LNeCttqs+QSSE/NL8LOHKXOaVVX8rrY0z+dt8WYdt+hkDHD4XOkENUnAiposQjPOjYdjTMfiBg
fJ14mtOsXkmcsK3jA6rKQTP2fWWJdYAWa4P6gI2SfD4AH9sQVJAlNvv7rsY3Xd+sPDi+TQNO8Wr4
ZyzGzVtsf3/Qpj+/J2G3ajCMf6iUFqegdStazq4a24iH8L60leuBYJ6jAiLrRJ5jtDvkibOXU6Ls
IK9do8pGnGlg3jMoQyCjweBLCtxWq+LciFQtt4TqzwlNljo+E1qMyR/caJhO32vvLZfAC0FYOVDZ
kd0RM+8KO87LIP9p85kVVKCV/j2hAfKIdsV4PCgqOlt9fOxPPCy640K80T4BEvC1nv4deV84AQBg
lVnDSY6T2b7sJtxP3AOhVLUvUTpd+kp3jYs3BVkcQ76tnLq5TY6VBNNRtjjJBs0EJll5JeIMIcpE
UsVM9o9HJ20QuukJks9/ftCTaog5zJZFuL4uN202PvfeomZa4QqXmvltQREKnFkbj+ztCJ3oM2p7
aJ3mCfsC6d2NezzePdGeLZI2hOkxBMN3uSC/Ivf3EqOoX3ep7ym7l1AzFpUrRej+ncrCcx436Wnw
5RcPK9V82LyceIOhL7rslh/BW1CcQbgxrDe3mjvxlzCCPWHoFEPK7PHSuQJPP/mG/Y+sEZhBbfsr
a5/+Er6x7cE8prxEHgaubbYdaDRrHHq2MOZExbRKHr7QQv30C93Ncuz4Gfsax2hRxQB7Lj7PvAbI
m9MpqNwCd66ievcech8c7pk/OlPlk6eB5vStLJf68ei6Uth3e6in6+yr3UD9oCid+5vuxlKktALG
SHK93GBOJjdzDP4RL285nvv1JTLLF1mZiZosz92+CETzpjSmR3a9kzJndo1bhF2cEMSpbn/gZmG7
hGPUr/JZ5qffETqA5P/NcQeiWx+xl1udogU6ay8X2RAo8hBOxQuNr3xc6Bx7w1Dvm+YRhT9wYSaL
JeO3j2gQniYW0BqNsnnn9yYhJKI4L2Pxu4oAFKwCPh3a3zMtgTKTvCFdIaQVxnpAwyzQDxJNptTf
5hvAjD0bNC6SpgEMRoJ2ZwYHBr5j6feOuiFTNEc80Z5Kc4xNsm2bUjlpetQvGLo96K7ZfkSnulvc
aUE7rG16/UOTF1qxovG+LhGhVByr75P5Jv7bBC7qXFquYvzwiIH1z8hsD/+IMacA7yiYR3xXfQdP
W2BpG4UxvlQU1qJW21UcIdaYEDIO+WCdcuYwLpH6HMr5c/L7C88n7NHX26qC4d3bxM2OsvK2Ti6Q
hrn9gLEOJJSOOpKu/mMho6nLYRINERflqyOr/4WDMQXHhiRx4ZOa68oVd4zHxcjjGuG/gZWjYkB4
kLwXmq21qTGwR26F8iKH2sgaxRwollFiZr2JqQIY6c4W6u6yhR+Ok3if17rG9GKH7bo37Wo/cjIq
q5/vKBSgHYFbbFIayQ4nlVPoKPnzDf5Rjmo1MyYx6UxRIlh7KJCwzZAB11+prVA31lid74HYpXtr
zmDMxUyjnaRGuIvOhY7a/JjU7TBu6jh6bLJwl/X7xHlyM3D+sYYTtilSHi6OJfDhxYPLZPKmVZ9/
W/gV1W+lnO7b5MHclxpJaE176nrVh7uNpBGhvGIlMwy7gDnKXX+K+pZ4B+2jyYDoQfMro+a9qX0v
zBWbqjx+qPvACngIvIN0H2O9/CcGdlX2cSlMuTkZSHwQVls7u6pNqgZQ+CWAEpL+oqLA1lsMEy0n
C0dXYMUxMMeS0opNOI/4Nql7Kq1PDu3KsZBlbbAuRp5rkBNVAe792eX4GM1FHAkGzZyZGyt3d2iM
SYSXS8yYCOUKF9I0It07jhk8bkfOlrEh4OwEZztHnoWPJT1L9/k8AH8uWOo4fwzf+52WD6rOPNZT
sjcGEHH2tE5CEy3RLKPdIlKFQz1dd9CmSjmz2rUbV7QUSyCNxF+t0Suv5Fn9qqysWG9jmZh0/ZVo
gMzSlxnga+AkIrVSRA15MyTsRT9qtds1yYBXqAPSlFK7CHbMl9g4CLov58y7cM9mefGiTl1RD6K9
bFNNoliBdHnKgjx2pY5zP2L1oQ9F6Y59FMnUfoVrEIDcXIwjOijhlmNXojtgmppUUmoDn4G8vpBd
YGzpFLC/FA10dPSnI+59x+n0Mt5ByBB7eoTdKI/VD7KWRgIrJRONX0yuonV15b+XxAm7slLu5D6y
0jdqe8MriVoh5MO1pNsd8j11a+bwpH/9cPMRoqmb7GSTpcGVQm20LobZxrFW4wSlkwQDBCew8gzo
OrmfgLBlMVdiNvPwqNOFcLLbPk8e4mMfi2CU9K+wb56Pb4SxG0A3kOEEkTJg0kzPuI70Y1bRAPic
jEKmZdGuzlKGtvwvpQ0LJkH1OD0A86F9qXBn+DdNDYuiIulRSn1MGxt8/fPjn3q6Qy9VkjvRUzox
0J8lWrhxWGF6j5OJjsmJFbMCvwGsWaeCR+ZlSyV4mq6lsLV/Nc2vzvdWwW2hv3sB65TjupLJBv9l
3Ea9raWgg6gG5mqzxRdazW5wS1Kx5agnl61xiySQ02soSizRffKfP2fdBz3VmblRbL0tI3GRbVnt
VJI1JV91oISIwMg+lLAek6r3YKXpB5w+3np1PkXc3mT/xCaigAsfQiB1BmDGkTh5FkpOWn2ll6/Q
DsDVnEGhq9rAKtbn14xiX5IQHO4DU3CCUdMBmKkMaQiDWob5gPC96YH3ysSeF4COyV0cnPXJ4MK7
RHfm36CGxwGt4v+fNCyfUOM/Ehxoc/I07+nNRa1fppGlJ0g4DnGBfA50M08z0Cp/zbohxvLs7LhF
XYpnfAgCXw9W05ZRvC5m+zKg7UwvzihquudyUurnY0oL+ztd+ock28TkB2zaOZQxvvTWwfKY4GYf
1Z0xtrdiJwKiioNjUArRjTdQRhtHEHyf0Bv0MIWQZXt7QNOHO2pC7FBLkrv4gM6sHp9HLy/eslBM
SddRapiHrI/DNzVxbjXTAirmn8NdN3WmsAiCFeYT70CP+ghWofPY4f5wJPT/X+UPtPcj0h8UJABZ
Fbik71LlueBvVwQT1keNnuWgCbXhZNIxDy7Bh4PLzxy1RfveN/AX0N3FT7e11Kb+anAoDjA3ztn/
Kml8VAbIuKYHTJsHCbXDOfRNPRcahVSsj9JQcLtcqvveZHJd1qWDsKsS33IDesaQCFAeWge/RzjL
Rbz6Glv46YbRKv0hlrJnYzbu/LmWUEsH2ZAvLMyClwrZRQSgK8mfRcKlY9G2SHoDeGGtfFkwoGz6
HKWyvzHKxGt/b6vMpCMHpSZ6xCPQZhSbVOtkU/bq9GCPWVO5vdcL2ibNEWeXMCuSZ4SI+qyg/4it
0MqmLZ1kZU4ov5FC+nWLZ1aaGZqVDC96HrevRVUOafNYnCHaoGZwH0huT8PkoRblbm6lhg2sCn4o
KVcuBbaC9kWFdZeKO+aWqQU7gydeOIoDrPI9DlfouPZFczuOiIwlyzCRlxT8x5ESGLVigRtA09tD
WreGLHh07FOnFyBRG6uXq2AXxgKidW1Rt3+cFDFwTXCq3V1OGm/wqCNCU2IofoBenjgMdxIXOVAO
RvlQqJCz7Z7noggDnJ7zIxUS85r6+XlPQEMz7yadqMb6e123pyQP7QqjbOiXLGdkUk+nGcz1luOP
WnqOecNaLGroA/v4mvhI/IXkK/i39wyWGlOOFg40RI5pFquonYV6Aej4gECulziBjAaHEnsunr94
yx2L1hccips0qMNvlemSDbyWzbxkspQoo3lCM5Qn0jIqvasdfyjF8dK+DqGLHE0TxWpoLzF9zFYu
Q4+nV7jL4l3uHzXz+tU0y/lfDs0RRpy5afePuqgy7xJZNebe6vfigdEED22MK1UWYGXYnVyzoMyv
PsWm/vGuip+8wLrvUoAjqfvgx5sjiNTlLE9TakPv4OSyBQWz3ViCej/SJd1D2ez7rsq7hav1uO42
2PKCIGFHZcsOs7w0S/UBe9j0nu+PSPu67GvqrOMI/pFpY1SM0HZSVEilAHnim/QsEmCK75KWIsLy
2qOvtoSaCkKwO/sQpsIpmPZazUNykcoYekd76M64KCqfJW6jLAVEgysUZoOBk8hDAhQYs8uvQYS7
FPqAuuxWkCBMqjpsmuczvMURjPIuh98i/ca2bx9yCtepLom25NJmRlP84Ts3yUPVzeplr1nKiw7s
YE66O+Tp0tb27nmqdrJVHQ0TJl+SBfTncJJLZj11Bkvpd3jqBMgvl8SL0SFzlGbVgKsX6z3/6MIA
q7dyXkNDNZRYCx3JzVygD0YCvrH/SxSh9QItW+qjcmpvDZRSK5toHuPzCPjc56yVqQHM4C5Vi1/A
L4Yb6kPthUIv2brdk4Msi7uKBT7fVXIcinL8Cv78PRo4mCd6+Eef7BXzki5hW1GX1cLcY08iURGA
9VOimQ3GRIMIvX34f20tuMNDi3mQYAKPb90tij5WGafT9GAaVQY3zdZsF/fiO6smF68uiqcwu4Ir
nCu4kBWArQAyrxIb4+hsKLAhkGzyP+IKOg0UANzjUnSGuGTTLZ13oBW7YPew3O2B6At4CVpqRDzh
KAN16LFVwRpFrlEtZSlwhVlBFMcvRzxZAR8DZtJtm3aLXKiCa3xd5itjEX+iLlReslA5ObE3bO6e
MHIWzgTJe7oUHDLE4uWgJLyfgJUBhVsriwJHRpTfjqV57tzU1qZezjPsd45DF+KVIKZC+cqI8IcL
wNpjV4Vk34BaP13yIIoHxIQ9eqHVvGRStqH0NApvQk/a1r/4iPTXzZMjM4T3cmtBYeLA7M0bqK/v
w7oIA7CmNRjly6MP2Bv59Buc7FrNKenjh7K6GquUdXa0okL1JGQM497RIK6bm3/UbUZ4FhilXFwR
ntmnYiBVGEI7zpb0lHkscKifgd7r5/yD86pByR7xVKMBeS35iqDKv5bVLl7xKgx3lfCQKv7y7+Mu
s7dxrh1MtRQYUfmYFS6hxiiMy52BmYgdd6RwHDMO2JPPf36BAG2g/xXhnlZcscJ5L2lPJTIPIADX
9M+fuwzE2y4oTSU3ZwKKaC9MC0EQl1W9nB5WdWLGf3xEWf48fh28724XYA1JLFuW/K4kskbEj6yE
aCk6U8V+Qgvnj4zYO0FT89FeyzQLtXYt8exzo8U0UCh16NqnZeeQ2QfzEZGcaQ/2nbO9cn50bFCg
QeY87xoad6/+5KJhpBZzulSefy20dXq1bfIvExN9Agad/B4gC0LfPeRCcR54qWlLFP9Z4KMDd0L2
Sp+lChyGrWT5jKY90CfbaVo1W3vjPNEvVsAzCG9b4fOFuEwDv8J3nPMNttrah2d3lwL2+3KTyCdV
RpY/48lnaxWAH+m4A4REsCJdY2vnDJZDjNZzb8lD7ZqMG4yPIpf7LX9OLQS2u+2wDybK3jvcd1pF
fLBrqUbwh14px8HAYmXBpRMhhICmsYWLS8pioinOG4Nm0ppIV+cR3kFdJM1c1adxdwyYtpLkmB7A
1J0eyvpRmVTBukEYBfo5N9Mc0dP0tt+36GjzL2B/hXU8GskgpLMgFkLPW+Jx15swx0QkElGTwV4s
ojiBem0p8SWPIF1a+f/4JWExYQ5ZWZZeI78llODEZ3MgftbLqeZ//61U2nQeTS+HS5sx3mNOzdRs
jwscOaMMa7syr7DfKhLvksJRSvXs0ozvuFt4Qzwf+27avGNk96gTsIY/9XrSQNDYu0BZgu++iAef
WBIc7rlZbu0vlAoE3AySL2eq8wDBJfL6rD29AoS6EeoQxcD96VJNsx9MK52SWOl65sGc9qAyWivY
v4Rx2uClVNTzwGLcuI0ZeOTdEgHUZBHPxD/1+SnjmqwzbLJIbDIPU5vTnJDuiybLC+/jdj3lqrXN
BkXWzFeB8MtaVcz+jF/ngYSRI6SsgkQyUDTPhbyrTwCb3jpz5Zd7CPRek/Xp9Am7HCaErL6g+Sam
F1x6fDtRCaKg5yEQvU+VgYYZ0erns21vD4EofUM+B8UdbqKMXVDhpUXArRkMHjNAnpQjOncOfKe8
CEjmflX3+ChzgF8eOFGG/7+ZyQRI+q/AnYhMa5RzSU0J2IALAUBk8MEAgTKfboC383u/lN/z9XXz
NqivUAgMg2sA4dokRXvxH+o+txJYqMJhmVcZNDDFRdbhSxeGueqi6inIx1u3EGXQKUvFd0Yh6FAB
QUlj53R6A5bhG8R0ONYs6IZWD25BqmZogzLs8ngJNU8dMox5lNcau8PpIcZObwNKaf2xh5i0G009
RhnKwu/UaL5h86KGrDr0CmxDYYLZnvb/Z/zwnyIQU8DgMv1jVtbt8W6xBUs9yIzJevJ1KSGOV/tC
n/HnH7YBlmLNIYsN8pvNq8AeNngTLA6/RbJl7xlCS7kuYe4xruMJFnK83gUz6G2uGT/u6nJH5xDP
f6yluUlS32/xN1w6Ot5BWK7ilcwPOazp14BFKw58pU14rYyjwvvQwFm2EA/SV3D89jOQryOZ7I7z
nrR7dIcSrat2/8JVIx6qQanJ/+MzpVpvIbiJAxDcy8RJKtkJMB94SILkw2Iakh7DxEGTd8+k6QHy
48JZPbqS1tp7cX9kGRLaAu7xWWGrEUDb8xoDLIl9m5I44RK0MtZ5uJd/xPmLL9Lfy3RDwP1KBy9q
GRjpuhZbA8mORBjjaY2cd+PlmhVpK1v+tGbznA7urYXZbQ84SvT80M/OcztpOOMwWqqte12JcGSp
+9d/9d1JKYjPH06Xek5Jv9fvoGnPM8x4OhQHVR4XSxdCaGYjhadMqhVmQI8HtErqwRPfV49ECV5A
4tjxyTwwWiH5OoqBh2n8WVxNKcADVtVdZ9qaWvQGodii2D/B4CDpVu/1soei2asWmJgPAyd+78cK
5FA8dqlivkNSvTjq4KhmwuzhUmGOTGYmycn2GsmOBAq7lP3cCsxY7x0ydMDpjtBUS8NpHSTGRuDI
Rk2nwwW+zq4usSHQKvcHVk083Bkri6j6xMnmZWiSLudDobiFOE2tPDCsmmEqvULn7PfEQ+LyzISR
yd9aRnqS1pFb5dE0sGld2Jq2ghkhTYgUdx3pAvEs8pJFeX3Af+lrSmRWoC96yKjbp8tEYuHrhdQ1
W/zzvzWiVWX+1r/NiCkO3hkUjr7hKQHLCtvnAw5BNCuIaLQPVgNAVH22LkGbpuGGEwQ3vJMscVLX
BjFMVHl6ekvRwDXwMEaksnKORVfV6fCImcxBYu2Krcq5ZYKd8g4WKXeN2gJKa171fmbh6xNF2F3v
RRb45UlPbwKUYHyYeL/1teA26Y0BrKFmXNjAAWuOwG3fKRK97UWvdNvRjpFgnPdCsXa0q6tLTGue
6Lcd4m7rOTyhyefk3f+BfZE4yITJ60cwOkoLZ4AzGKNOZ9pUstepvBUZPCEytjkrfqhRjoyO64ge
N9PvAoxrRBMgtSyT0vcTNbdxbpnTYg3FFKq6ufh01SZ/6FCOaxnDZgc1FFgzhL0BRiPIaTk/YXuK
2RzB2m89pFPDP3nVdpYxtHhbjXe1xGr4NWqGvw6b5nIj/q+6CxwBnpjcpPd5FJe7Bjj6IpMVbey8
rPFwDmixIYcmYNdSH35sQcpKcP5XWX7x80tEXgWHNWLmgHkVP1oaO6fvFVItHuVacSfztSpO8G8F
CXAa75tFKG8htM6kl5eTXLLNFnlQqMRs/OmhEbDbXoNh+cSLdwlDgyTyBxCwj3rB6RUcFP665xuZ
+B1Xw8Frpt5YWIJx13JiGbYujOEjS9XBk1roBU3x9Ts0gxPOyCN3L17V1u8VLUPQ9qDmzAkqtjmx
GRfvvRK/NThA2UrCXaiUq2M+UFNeP9TsRNp6rikaVAHZVcdNzFCMJLZHpul+D0i0JZ3caxY+OVzL
sJyvTq+BU64p8gaOE9q3u6pPhsPf1WPwbFYPpcRU8CobENm1MmQEZaE7U7DQm+wAzxsgnrJRes8H
B7eSOHo96HhWKTBXI5fX/8In/nc3eVy2gxpqkVxIsPe/+lgd+MRqwqNdNspv/oxk22t36Q6/oBeW
e2NE8NAKG/P/U40JNw0H/2oOsCp/0sAI9OUc47s0qiNjjWTIQyOEDcqUOtPvC+B2fyo2oshKJCKo
lFF06gCCF9Ns+r1UbBSSNcz1TAREOgBoARk+Tja8Z//Ic4DY1cb+tTVmw5VaZyLGIDf6y/AN3sMG
u657/mRmtPYKP70L6buWM4UM09hC7mFK/0s804blB0uljABnb958uNk1v+3AFB8ApIThd4F0eRTT
9OKHwPng0Ge947Pxm+lJzjB1Og2Ux8eGZDEvpk4YpJbD7KTu/SpFliHph7bq2z9NPS2s+arh/Sj1
DLQmIB+IfpWYMRUpvYKdtXY5mL1O1+uNqPUtEBWCqbIEKs8PaBfDOQ5gLsPPWq8Q9Ihk8r/l/sFx
PDPysEEWLbODqXb8AvtnsCsWtqKj04Sl9X1Tg38eoDk2MHUe0Oeg14N4lzV4VCSjcepOX4WlQ6Dw
1IYuo8py/5/BRRlloI7qV2Q2YhC5X11luwQayGgdgyxeTScPHaSe4nj/nMNj/OadUmV0cFxJZ4Jk
td6TTpFloABZaw3yPL0ZLMh5hkSmlPvdxjWl32f7e+t1XhUWv1VdIkHXKIXERSyUAXy2BhPSTW4z
ywuy81Ogy09cEtTzBJ263Xov3LL66sP2Qo691vJu0zE9y/TzqJ3lxkGZmVeOcqBHvbAfoVqwh2L6
TtSKXbniSXKP3w88BKP0z6SnKurcTz+H1f9WxZMgx14HnQEEGOtzljdKFH5k+rTH/J7jPY5bYsVV
E4l4FPUm8UV04Pmwxt7HWVjIIu3pQXXXpO80pFi8rDWbDXQH1NpvEYS+E2Xn2YQnHexEydRDcN/p
2rNGOPJfduLEfhe5VTLqFIZn6NW7ditePGd5DHeWKz1zdQefm2KW5Skk7yaOQ+rsPbMxQU0BvfTE
PiVQCU280OSDXvjKqRyMyRcSnK7A5UQeGDX2fsAsCZp06qiDvkO8ghrnn3cwr8hRQcxQ/SUa3mH1
ZRx4KXsE1hsw0BQ1Kz9r7lDGCuJ5h0aLKMIlDwBfkUMVf7Z+S81vCJ0Ad8bimZ2RCEdOCagKb/SU
GXr53CNRxn8vyq+i0POOTgcUrlQTLfNqoZ6/KXakrJZh+itCGkS1cAR5LlXVBkAoMKWObPeurX1y
jqXVimLhB8Yp0pHj5wa5oswmrhZRv9kx62dgsztdo5BJWaPlYMS1YXqqHa6V45xxLfsdsKcmFAIK
aDcaNa8Cj1RJPvVIyNCgeEBTqY7LvawCGmjk/byIrKuXngXE7T74tqVpVMKvR9eQ3j2GfGPKaNSE
HIl19Qz3sggz2FgNYELYMNbQUjfSnFok4oy/RNGLzRM2K/yU+J6Gw7tIm6HsaxJbIM6qXPkQp4dZ
MTnOuv7GoRbuOBtrE6C7iULlo7yePiPPEmuFt0C2DrLiulwzhPbE5ft2X4wrhMLTVvQCW5hJUJCw
q40GYOvVFuV9xfhv5I9HvP/kBsqaP1Qvvu3NZDAyyh4JNHmvJyh1uM47m0ybnLQVVbQJYC2+lAKS
MzQUwVuy/EPMao15MBNcOCl3tFSBOeUGpIY1m2++rNcDtLuqneHzpoevG+IPHwNs2921/mX0qKay
ziN7y2okeLp1HuM+zLQ5ZNR5iDOp1EuivIJs6FNbMA+nD3YVIJQ5CQAmz54TCziCcjE0+02i5+1W
rdHpXq15R49udfvBo9sPacMJD80LJb9iuFGF16IyxnBpN43vE+xc8Ki9AS8Wf48LH8IkiLanq7Uj
jisS5r4RhQ+DJ5Cw3Jmv4ouNb0ACchwRT9lmSXd6zMjQ2BIvdMnG4DvI8clhLYF4BBeC/v6sCCBa
P4ys4FB5xUIlCPMZc9K9grbT2tBzG+3PEwY+EQHf4MjhWoiI3f6Y+mXMpVSNA6tVqVrhgKWa2hPF
ofiLzOPw13HbVip1nmqefBZ2uFCFutAMM0vFa2EU+KE0Is3s/85iRrNkp0WocVnZ045xOw1vqJJq
g5/rZGXzeuOIxvuripEnOsalfCJtbyJEGsn6T+i6NoeUeiMigKBmtjMiWw1bbPd3+5V8GrWSv2nt
MPSiwTM/hauEWknTYRHx6ZhYCx/Wj73hU4Rjqvq1IzUJm5L/45B9os/zPyS8wE6tum0r+DZV1vEL
E/yKci5Y92coC7ixbO2LtBiSSm7FnoYg8dQXFavCEsFjLbGmscWPAstH0z7+d7ysuJp9XRAEYAjS
iKUCYVON7iiBxjxVgO/wwp7uqEQ0TPpsm+66CGzbIdtEpnEu/+X5qNiWv7/F33eYqUIkzcJZ4aHF
wocYG4QiepDqUz1qWC37NDmYXbMmx9eAwaEC2TGw8lX2wocaNECrgTfh4Rq6BrLe9sDRsYP+AoWj
GuGayjqAZjWBmv62XDEJl+M0dkAeTJtFLDb98pXEecC2E07ka1TcE/D6d4PP6q9p0uBlI2Auf4qj
4ncRxvd8BvYbbiFqIvVw6fgYjUrLQc9RvxOztfEzyUxYN7bKqm27JqxkS3eiMCTozO9MefxP8Ro+
0V7vxWQw9tWzoCALzoBiuuxaAo9wKBd491jspgqSX5cVupdw2CX9YAlPn7aVguTpzAdv1xaFxSKc
ddBiVuMMHEqr2m+ayNX0prK7O601iqCl1FO1H1ry2I2V/XGpLgftOrwsL+VCzI5f+TGBu15eNMRM
5/ygC+tsmaEcmTLV3+l1gzyKNQJq3Fd0i47pHd2WAAxh48Ry2cGh35+farep9lZELyVmv88DB5GQ
SQ08fp1QZqdewvDKTJl1v8QcSkHvsj1SLNMzSOCcJZMetB7+ke5NNPvcx6BGDCEeHEJS/Uo3lfMr
PTirhnyKxQcC679U8a7aZJWxbQQEuskA1I4raKqL0UBGBxwXJhBe/H4edLWnJB9YoNWp3pjoIoso
JKxpNvXC5ay0wdhyGfQODG4PHAGT/5xwnha9nOYDyEkj4CKf5URKFXRM9Iv2I0YrSnmbPzHFU8Hg
9Ky1gqG08Db1ty8tnCOwu7JTDQ95zYb47jCZxOlePb+zLWx6y4RTekiPIeQaXNckroA5EVjmRNjm
2E/Rx1+pfsp92LxC9i9AG4qtEp+/CdGAJR01suannPF4G4Aq1iEIrXYiy3DXMJi+PpxQ3B1wi0JS
AAAWdc55LDZdbbIPvKg+5prbOTHhrrbTh8zr6Ms1hHN3ViPbIWWX/4MogG7zkxuruvR3ajx+/Soe
Xz1jh9hZsNz/v/40h1EibGQy+MWdPmmG3X85En9w3OGiuJeQtAvf6idmBu5z4nl6A7wkxgROukvp
rH09qb21cyp+qUlEc/TRvY17uaSpxMMFHwAtJoSfLCDrzDGAqaJxklA56rZPq3MfzQqTPwg81yTs
EbVxel1skrA3kXfGZZ30tf92nkeORRPb9PZCrQJMemmzCXi3a5Kk2TF6HfUdXWGym2vea3Mqyt0o
ydVFf1pRJXYWDDHkspc8QT19jyTkQ89hQEHUiydX4eE0wSGe5DQWrQyx0gqwmIdDxgqjnbQlHtzp
WZyOg7VoIbLgATH31KA1x3pdE3vDDWaMsD78RxsFooxNHV6y/psCVKt1m7vZuVbLurfjtBFy43Ku
xNgLugy+Aiio0D6xRGJsOyofnHd0MmVgWYD2hvf7FMrw0beI0Ff2o2z8nJEAyS6rfOEJjttK/j2H
Fb3WbzjpyqWyisONRHILlfVvAgDD8sA1BD5UJACadH0yCQhZB81fqH0wX5Hh3Hgk8fdjcDZaXQTj
JbSFndj9dqHSN4I1sWfJaez7pCXTKrFw26AfvUbO3B/+QwwPEuaNRY18BfXu8DNdsMiLsQJJ7BPl
78X2YtP8PwCQNWHHSJ+DZbDL/P5Qglogu1RvATztxe2QJq3rkdIl8HwyG+PbzP7fRowprPV0EMB5
6PGJADx/OyZoNIYnQg5LTIW2eOGRYxgjfkkTf0PsMXz8yDMyfAzysX9GFkrYDtj5gIvOoVT2epdT
Pta3E5I4XyxsbnHi3ttextpUrFNapfQsINH90xCAqLykcmkqp8awkfKDhO/KcVvYdFKLs/jxURz5
mTcuMQoGJmrsOUXUkP4tPI75yznjuBLZNeonQFubXiO18feKXHl1ivPWgBVwuqX320qDM9J4TI99
rGc4jNhjF8iD0L03PYydaKYdxCP4bdQYpZx/q/GdGgSjCT3QsuyDTxXi46B3d7b4Oc7ULhEcZiZ+
6HoGZQ1vago0j82sEfVD20kxILI7d+Dz1iQtGzA3C7+Pl/rMMmFeD0HPiU4KLFbLRb4Qz/7FAfnQ
S3LK+nH9c7k2FTq1kC1QljCpCGx1mY5UGWRVAlJA7fm8ZPIdHoYr/1nxIl0ZmV0wK4UkgMiBvoMn
K3EaGYtPKF4rq9UZN4dxcHIntjKOIB1871ryAdrGFLuMzyge3eeVsyJroz83OpxMzUAqQU21ouVT
KnzDyQeOEhZbeDhqOptDDEhLcJX6k93ZZt5FIjvcNw8bWcNCDlTO5SjTRSKMloCMdvLokcVK1AMN
jf9S4lOAXoHD8ZTvyD0c3MoF6KhtaB0liKUfQ43oZrVpf1KD+znXPdWEpYcjKNitbqJndg91y1h1
0R4EmirmOw3obFrqgG6MSJ6hkeIT/pVFdkdt02YfHVLjtgrb+QbU3J7nnwN0xCYIyq2DFuXHVV5K
I9Ips1lkipGuFHW6ymddcszn8bJCWfgTZScBm6e+/DA09aWBzVw3lngvgOdcCCauGxK7MUEY8Orq
SDwVG3vQgdX9pRE3vnIInYAkaVz4cckUFNXZUtK6Vc6S62VwSeomG/c8yxUDUIdrpKcyZEbse/8o
q1A3TQfDB0GlrI3IH6TeR3Bc0c6q0kfbEFgy/05IRNbf/uCffuS4ShlDDmob8mhLUFdEV3P+1x1l
EMTymAzTtI+4lYNNRMwhOHtMg+dOSdgffNvKjBO8xgDUkZvMMbGM7LhsYShuqfvUiKt7VJ6EgpAY
H917fbvTeWnOfCg6fB1FEY53G4ZkKPb9AMSvI2nnxWxKBUH9HHSR9a+3QQPd/6JTBHLXdPBzSS6v
HY86OlMPv6bleXh5Ht+WqrYGlreUoFqWmeRqn9ahpatqH71ga2jg5u6CuGfdpqeMG46lL2ppUVpM
3x8o02WnCMakfzdjjUqxEgNQ58H3chmgHPsrQ55dPmtQhJ/Djo7r+M0LiiFTP9SzRijup0rlSKuN
7qvng4eaJiifWf4F2ccIi8R92orN7v3ApybNie4xNt+D6GW9z/nlvtkWxzTOxtMROoXcaI57CW0y
nrU/lWq313dGm6x4baClT8r3eM6fo1Db5Yk31JsSh2SZNtKImvLZWwWFN58h2+05KbWyB6ZHz42O
GwahG7n42sdtIP0W33LB35QfVeOQQHzWpD+gu8P4YllLe3s6vAtZNpaumCKm9VB5XO2fGMdc/uD8
WLw3xoYhNiHS8N0ukk9l2lt0cvqN1K1kiw9dDc5eHhBOxt82+my8dekeyQZ0VQQSMrpWDl+AGk1Z
l99urhyoZ3mMRJXIvLtUNQngCvKf6Pd/TXP2RmW/JTZ7jg7FaoKx/8xFN6gRf2cDVQIoGWb69oPa
4C5In/2vACErP4DcPeH02mzdID17bhFFuueyUrDAREey8TAw06W8inaD2Q5gSQbU0BhF5LpEiDJG
Q5028iVQIvsskf4xtcl55Ev3H1FKiOqIjO5ry2S0uig/A7ekvp2gaUZ/yAlen2f1PCvdqMXMuOba
2RLFWKCYTpmjRVQu06mBdnyijzpXU878DkEr9BiS6ME6OzXtH5r5UQFhDMRZiF8l+jhJd7aqfEIb
r0nkQf9rI/4aIjuVieqHTv5+bxEnXpIpVMEsKtXpRR85HP78SGZin6kGuVLSK1akaaAS0jkVX7Sq
PU51uvxGtGjD+6DQTZ9gwGK6EVxRt1SzM5f9Brmz6CMXbmdFA/juCyJbH/xiU1OIMOO+Y2xwcKP5
+LeNfp+HQm0q2XlURu0qn3+Bh2sKiKwx9KjmZTEPfEroGiFnGuXyZPeEsawJvQKdCX4sfRRl/lKG
CcNBzPU7VpVPQmycUWHpnW3M+390LMQAw1Mhd3Q8615ufR3Lo9UB9BsSmO1Erv+KEz5HU3XQ5LK9
TpTFajl6gruSNtHraf/mDk+kR5uFezVo5hQ4VjQAMQWQb6XJlguF54qZx+Wn9fDAG7ujcdJNwCIT
ljP/LxfIegkuluqXtQaXpWtAczOWkb/XP68xxr8pWx2Emdx/kLvLdkqpVjq+1mQviBUYOBKHEfVS
QYvrahRQmZIEF0tY2GLuq4cTkjG55CYiebuw4E2s01pesa8SAkRM48CYFw7HyjLsvVlML21pte6P
AA7eWfaJM+H+cVvvBNTTZKfUEHt5XY2ARx7pLbZp4LIoleeHfc2j2I4oJGksBD/LAo+A+8x9dfr4
g7vooqowyk0fUhDs638biZ5ToEfA98gglyoZ0QVNwNFu/tq/s/0UyVmE5kJ2iZcNmLkoSryGC+rU
yTLGYCioqhz1WE0FUww9tfrsrrNaBIIol4CtzU1jpWqIMwSYr3Ur0J3OTW7wYLy+U8jHBS6lnZoK
MSYJv/uHipYo96VJeXEIIq0B/i9DzFnrAtyicE6CjtzOLbz/TkOOXNEA/9tnY/t13Y/hQJXV9gSe
mVfy7/DOYpANwPQcn0BKOxAY1Srf+UXhtU9mDtknTYTcbjLV2E4uYDpqPlE64FCnpXyGgBRJRrLo
T23KIcq925YbB8AC2ISCwpfVHLQ0FLaWsEMwqcVosk/G7TAW8t4u6XpeY8ZfsXwAXmVLBn7bNEWl
lYtrV0VF0e/RmNDHiPWGapr8MUE68xLKU2bTT213MgHkc7wwMQ6BtnDW1OOZ074SCNTrWIVZIEv7
24Yg8StbpKpXts6xFvl15/TLMcQhIItH/LHyFSawcv36OheJdRRnMvdMvefMFhpiRpq8YvEAWYpw
bMheDlLR++hckc4+mW3gduvhlBB8UR0z+7v5cGvSlntcTfkIhivSJLIgnN8oC6uD7RHi8nKgvywX
NJX9ui4PmUITq1EOhFH6+xzS+RbGajkS0Gw6JbLoy07Y2CU2uqN/e1vLLIFvHjhN3CmE7XPt84Pc
rjMA9eAYP09ynBQHGdVQYj8JpzBdiwaY/pAKN2vzKOW8wCxIlgIo6jdUf0dQ4dxqQyJfzMFfp0H+
C7xCygt7fm3utKXlQWsRSU8mpMb6mrmZd5v8uPObNHKPKXLPtu/47OpWAkweO/mEopBME0/4dYhS
urWw8JFlI41t2wwPEh++mMzA6TrxJ2DG3pu2C5fJlS/afv5ATfJ9WzWZnjLbce0GyfzWtp3TKBQ5
X7mmUHYvlMwXSzc0QuA+vGvHrjhrw0RuPuIPdDm9ZwghFSvSARcZtOm6QBBwWiecvGQMZRf9k7sO
JbMgNd+nFW67DbqPcs/aTPEz5qr+bE5fj4wi2CUdjncLgZoz3XEhEkHR5ogrw+9eXHOGdTEnBYPc
oBGd5eYuNKDQcmRz/g4mDZry4XqHe8xRxBnSNWFU3f1odW76cloStVBkuD+zTMv689/U5c1KCk3x
+lTjLCeKV5EOuOe3GFMnOZERg/BzFSsGCCrrkSgRP//ELmIgbtMrbiHtJ2Ftf2zZdhaKwWK5EWtY
Lb4TV26EgOtNOqAXjg4/JX+4lt+1TjffMVankmfkgtOD1JpkwtZLwJpwqbzuHz9qZXJPStWsHOtl
OSRo7G2fFsxlN1RkuWKzIdDY0XyFetTU4THwJeZLES/DXZWJF4Ep4qmSUEvj8HLI7rPr7wI5eS3G
VK9c+hazUcyUf0fF3spgoK3PwGjVeimI8B5TSe+xE7gEy9/8iWBRW+2T3njis9ECgzry5bMx8Xoq
7Ma/T0wKfAHnw+YC+NUroADVfpEoClVXe61fukxXpik3yF1o+N46SQ6nL83XYOesergwLXaBKbAG
xSiSAjTO3q+1Hds2V0Br3/GKHw50tLHHFZ7mcTsZt9Ju6TkLtCrkG844U2kKCdWGWBRjrdI8znRm
ozZTjP72I0w6fM0AEDOv/ELsEfRIkFCudbeRDxwtzPYxenFIk3rt6+6ZhfT0Zfe4b/d/YDujfB0Z
Pes+4GCAxq+HgygTieiZejUUwt50JIJaF9xjLxFlZExlOyTe8dfcxfGy+gpxqtOtReXO060AX8Dg
H0I/oppsbea2yOupjC6oSKxagCiJqTCACCls3JEBB5mV0/EHj/jRUlXDLM68d2EHiNVl24w8j1qA
12EWyK958D7/Bi3eROtSozxOWGBJOP6ED3Ui9UZOSMovy5L6NdeocDH9qnSlSzfIPoNM2d/chcqv
wDTYTAJYeK2nHnDIl8zGiDh3WXBN8GA2eQP7dJISvNJ6Qr7q75ruibIpVLqHcq7MI6StEyeWQD5n
oTv8H/N9DfyEcybqvG9egR8pSSkq0QcujDCYyNgDYdpAPkHZdurXeOyZeRhfs9kDHVsyCVV9HZnk
Vczd+TVGAFQDNIhuQODWNyuqFB4VfyqAC/5z2ZlVN6w85V1o0ZzExyHaSjxX3DNmFW3slvOq+wqx
Lpllp2bapbpWARhM5jr7hgOjXXy1DNzu/qK+89PKXxBUvvgO4fo+M/sb/gyf/8uoMHu8FXxQ0eg3
J5cqbFKh62hZQp0c47kEN4V70/0biaD9PkUI/yLRlM3LGwB+LvMQdQ5h15u/c9RxV1+IyxRk+g+y
7uuDJfbsT5ss2gAd9SNWn6EiAR7G9aO21O/awFppCBIfhN0m23P/0dYqMH5SbpQpsv71zfGezj6T
QT3rcaTvx6T+dwwoXr2DAXFEKsO1SlPhDgMOHtxkpN8pu2pV2mdZu3TM+vEV4TldkViogGo/t9qL
DLWCfKF8R7pZLhL2xhJrL27AsH1BfwmXdEIrxRBHMWXRVnHVQ5h7gzvhdAuEc/RxoxJB5UZxPPjz
iUIgDzde8YSxRv1RwLB7XqzL00dvw2xzmARLDnE9gpwU9zGcritx3uMsiRNZHan/RG4VU8V5cClm
YIIxYvHof3CdLpd2U2AFKk6M/twCsVa45C6Ra1FdrcKED1LZF2uGfOi2Y/N2opBH1spRm5ny58dF
rFIaC1Sxt/ieQAsxrzI1e9D01YpCBJc9lhdFjyRjmIlXLXz9bmNqsO3/+k2JxwR39kDZvItIjXL6
9VuVST3pz/NXguHLqjfo7KCdzCS/Z3oYefC2NuLPR2xWwoV0RkhcZ34iTXXhhqjWMDNsyIl63XfV
hhExWUlvGmeYyRuoNsRzZyt0R/wyi7Dj6sN972q9yQlvwymDCrHG/JKuz35lWa+P3EnXJo0BSupZ
wXv67wd/oke9PIz+GrPXoT5ogFMGaiqbTtQ8MG5AbSxm7DcOSnN4FfJmFL5LDP66JpqjluiYFS6A
tgOWWaOacp2T1jZyDi/TVSNj49qzJ21WNRwxoodME8RV4BEcme0iqJ4KRJ99Mev1o6/XskQP3v4+
2QAEt0ov7y1iF37Wl2xCBjB4O55MUl2LwcMhIfXOLlDyLlXBkbRMPwjKNCGKUHFN3ryq/Ql7ZzUG
zFxbjd7HWQpPRKM4WnKpHlb0jTv1JtBSWtGGnnHLbvosOdahjM0Xwks84UBDLxJUXyRwxCkxExqV
scucXEpPXUN7+PYkUt2UXfdsdSp19UilUeplzZiWM+v5x8QwGU6zEbKz15MH402e9hM0TSJ7M0pL
MRtNuI3Ph8yDejihulJsLv7AWLbsciobREGg7XGXOv9kpGxQzms28ZzVlsI1xXEhb1658crlXOXS
rWrB762anpZpi4sfvOng5EU4tJtXH1kiTLciq1AeIAZm+oz0perFK4qzRb9/6sWagR8q9aih/jB0
KA92dXEDOKpdNWpNQpKxjkOvcSKpWcCLlKAGcG2upAyWA3RWVeiwj7HXEI6azWvt/xVCreVcklQw
Y/dwQlzNs0onsGZs4DgzwTx/IuWHYB46YXb7Pyli2/c17EdJ6FucW+nAXzdKJHD2ct9nXEpq3Eys
7pvp0PWOof6HnXjiXrTN+RA0AKMLELr4VjqEmSLToU4mlOKNcGKuc1bCJJIjhWt/6uIDXQk623G+
NTNST7DzeWjI77y88e5HjeECrwM0BtrcTTt8Uy9h9BbNsRs3NY87r3+lQ6C9OYqWIWFtieJgE2A5
ZVHpTL3uKXps94SRis/tCs0D5pkhouRxPjza5YMlzUj0rU8yRObTMAZW/JtoG6pjDnb8wcPtumTc
0BvVytmxSdYRFcpzLpUZrYwAZRa6N/2k4g1l6mPmgS85JiS74rqCZtmVXZuyb0Hm3I/Rtu5Bm/ET
eJsHrs0HOBeftN9F7rp1Qla2AuxM95B7SJdoBa8HgsTPjOeVPIM8SJthpxNL68H9TloaR5VkdfnR
4Sy6gPmbQ0LU7SPgHzp3giYDv7IE9uehSkrTxoKP6528RYWT2gNROIa7o2OFyRWv/dY/T53cdiz0
WblpoZ3hCO96jCwXJb1NP2oEB+rB6BJ5bQhRLhZz0oVeksyqceUcKo2TrUoLLyShXh+VQn31iiGa
NpNStpw1maUXuAV87MB+h06xAPrxzP7W7LpO3LHy3veWLS5DZlofvCSKh+L1qrXJOpf6kHrDY4Pb
Kwra0eGtoK6Xa+74sEVICy6xz4F3qsmitmf8cp3ulgexZOP9CYK1ptshVa+lhdnv1wjAxP4x4tzH
0pvQvYPjMP8G7fnJaq6D2eI9HkDqXQiTT1smpSwLl41hpacOdppRAkMFkga3mho2l9+gxXHBtmBN
vzoXg5ImnsVPx3Nw2pMPgwMzUkGJXc2fa0WumqRGhM59lidlDR2Uc+ULzXAD8rsL2hgrzD6B8SsB
1oyJztinLsEY406ztZO1ben8R3DG1vxLA9jlQIGeZ6vDUyFI7auNvxfTEWggFI0xTHRmlckXZ0HY
pENBXO+L0QWFSfgGfmEmUcFFtyefff41dZ67zFgx8W2QeKJgoKd7QUeeywjOjhtEiR4WSobxqhKG
QqJV4ELHTg+ETRK0aX3MAAkGRXvVo69XP8ZAo4+/fE1q69udiaCMhIourRgNgPvLkMvKGNWoJQT5
6j8RWfrdLFdcLuDo6agtVnlWdZVWVA2FoxZ68Vl+L48M2+AbgS7YpFM3iLG5H6lxolh2+AqSbtl4
D1B8mqhLWw7Sr5nWJncdWE0QWoWJlqyQxKjuVEVR779/OizsMxyUVBaYMRwrYIzKd0S/arb2+zn+
wxLI4G5086z4OVxGJhDhs2EXTnrBb76GoqTuZTSPdhlZOCgNvzlONJyxR+3pwaZuQJrHy7ze2cyN
37Sf93ivU1tohNbiHsVeeK7fcEccp8bkQiUvJe8MNu86qAHfJN1Ye+QbHrc+Zc2lbFx6PWMi1tB2
8qbL6xfmhjGnBSq8HwxRYAVOmnPPwMc3PmZZzAitbQyYb3VojrZKZAhUUSdtkjUuv72Cj0crRf1T
3/eiFE1s84ji11Zs1C14nRCNf+SWflIG3vyen6lwGUse2DdU13f3E0CEvqeRyvNDK8ql1VCJNxu0
8WuvY0t98cvFwBSY9Sz/wjTI6G1cmkXohkOGGKf8gxvIKL9/yv9HSnNgXBvyRRVDeI7nCqQsupwP
EyclTJKxmLtsJ0yZiCYsXz/T3+lAektWeBelWig3vCbkYZxS51MKWRptgTCZ8bUzqtrzJ5GlOHQy
Szyr6tIXbD+hLfycO07XfAyaNoEMelSyZSCzBypzkO5kNx05htyHPGDMEotgOLYKWf3oqS3MPTOr
hQ4pw6T8qSpHDlvdCMKafjLR+FJydWLgfELQlyROUa5Z88yt0zHo0oc1rlSbSDMSxl5Ajws4XPNy
qDwHVzEOWGdnT47TJ9CwW+sBpbypDH9nHB64G96WaXsaTxZLBWc7fb3uagBs7u/PKzdycbV695YK
LbSBo80+Z+W7j+84RFeiUYCDc8MUcRUM8sGg5Cu2cSrS7kIOnkuo0rDloU6guo5m/6TM1xP4iTpz
hBUhiXkneZU6W23JcMLQcMFTGStVRHByw9nuGHUvF1hZMS20E7y9yWzyBsrcsX2LkVT79yHC7WJ0
pncfFMaLVp6yPAUDzYzSGNE6iae/Hs9e055q9CivYggOb+QC+8nI71eP52hAMbyGx8PgmU+tvAQy
s8nxz72u/Fd6s2EpSWBAKBBS++RtdGLZceDrXJDDxVdKeFxGgN9AtkLyoiYdRkq7SxkUsc8bGMfn
IlrAhe9S0jpSWqsUhO1C1hNd+uLkATTtc4ib4tvVdQnm0ZWRZ07vyAebljtvrrk81DuGPJWgzdI6
07Mpv3JhKFPccJcl5xm0gA21OeblIdq1d8Ok7s3pE/VZNAxKG3gIkszj2QHhJqcH2prT8wr20sts
EuxpaVEJXmsFT0YvtDlV5Vcu0DioZ4CuZdpapMMyyOJUIIpzOpXvk7RPnSvyCR0WKf1/Ubs8aRqJ
KiCEOocVADlBYmNNjL1MwtHejAc7FdMutoBcM/e+W8q4dxla9cpAdPi0+AwOSAkcWmQuvTn8smr0
42Ml8QYq3+Q7c1h1UchL1lMCLi8YndwY4JhI4GNuxGwbgrCEVVSf4xecxscWYVK3YJszyYb5Cm3O
5ef8hNhZR9U3HGDjgdlczVwlVHZu8LuipnWNFMA4pdOlLicA/kNFpo6U63JzM0Vu7aYML4Vd+xjG
KVTDx0u3ZC5mOh0ft6zhG8p2EJ1j4KClUup0r061+M5m74i4zRTOvoTjlx0b2mwD9bBuaW3LzCMS
ySZHi2u/IElxupcVt0fpCGOI47v/x44dyUhtpEz5s8WRMtvWIfif7KrRuSQzLVssSCVd7yD9IwHA
hWOhzSdYPhPaNRTApaulxELP7AZUNdyKmHDhe0MQtPwckE4rZqWxQUmy7naDkNQzMN02ia4Sy/TD
y8FuHPqzADTU+oZ5/4Tdl4bcel2Py9oYcQam9H2jbUO/KG2xfn5hg4UHWn24ahTJOiqxC1wVlKTA
kGzK1rWnev8yNBB5/oo7jfImDbXrkm+6HGWDG2J/NxAiOLp7jMaPGEJWf3YN/tR+PCDeMiE3G0YZ
lG+2J7r1BPULdd3tzThQMROsG6AyKqygA7Uo3WS9VvrymqDYNCfI9rIvyrKZBwe5I1Eg/HZrQFDN
a3CyNIpnNso4F8CyDD/9WOQWIFMD14kxVaOb+2u0hPCO3Pv2J/4jTjsR/WTF8QgMroLKmdhxTGek
rrzaFA6ovXyk1/mC8B5FOgklwxa6cBhEEjiZSILeLrLvVZ5BcpHHy1JDpHyGahxp/rhSVPgKNOhw
aABRbZxqU2SvVSXYVfVlLBXdOqWp/tSRzJDLmHNJApItfqYHVwGSjzMH0QxVx99/x6bDhavYf3Of
sQ3ldFt3Zk4wdM3zihrdKHaXGh/hYEyX3zGFDR0kPoaZ/8CJdBJnTY3Ad3FKKHMv0I3bNe4WO/O3
oVjm+IBYN3xpyTvlOjUJaV1TFCnXtWEm1Xo2FSOUavz7NRZoq+HO1CbZR//On9bwj4uzCuP4dN3b
NU69zHm1ZuIDCamzqFKldLoW0jHkl5Ud5F/4RyKPKADzCTbd2JyZRTg06vSkImQPLN4x0/SIdo9P
fgy5VWQyADSO5l9U2hRYlYj0y5PoSrtvawwrtQHCd6zUjW45l/fVeVOi7Zoy5FX0G2Z0DsVu8jW5
oRoQaNgKZNdaiPmoi46y/Wlk2HszcRHHH/+f9HrUtgA1M9JTW7Z1ajXTe5m29TZbT8ln8gOo4KCC
BD5XE0tIE8NYS8YAcNJSrvASort/0lfD6fFdSauuoLNRhERl+mF8bwFC3pGs0Pi1vK47bI9pOIeZ
E+9sIRV3SPzVTDBreXhVXJs9vC/OkFOXAEnf4td135Hfojyl+pE4JCpdIr2pLxZXeDbenCuaDZDX
TwiNzLtIIb8lDHZSocDwB8+MxNz6qmwRyUKTZJWFdQ7a/eSibIq9rJug9zChIOhWnIafxfBu8Uvh
LO5PQxSLTKSbANC/fvdpoNTh3+pmZ6jAAXSKAtRDN+cZGKrP+MdQpPU+fIdYNpBfkXsp2ZxawhLY
KjjdJ1MGupxV+sU0z/1STqc9rVKNH3Qo/IizdboxwlrjsuMgx+yj0rpKqwu/BcZ6gJ86oVHB2ZND
97Aa59PhhjVizDu8YLxk6FCkElf7eJpTubNMNHDfB3Gg8gUx1wlbyLcZju20iAjgK8bJXgt95hQp
mZkqRI06d35akEMQpTIv2YIJ26MTkNRpirKws2cHnr10NxvwRDUp1GTFvnv3cmPlgB0vqXKyhK1f
VmAn9ls12tmvXj3rjGzhFurfr5EA08nvTlNZLywn1bx50kACSxWYA+6ZHgu/Gx9poWICkt2PwcD+
AEck+85idR+kB80oUEiSosS2EkfoaLDMUL75Y1vipiZ/ZJi6Oi1xMPAKR4UeVECcqdzQVHQDE5cP
HnWCXDtwudZavH89zrR6iqsl2eqgbFuKodk1Wdso88bLNFF8u9UnZRMBQfuBFpNlHCXq2UZ+UCYG
lK8dJWv6WvMnO9UKqKhzsJhEGfyvEvtH1RkjBAt7ZHvXci/9Z2uwj/hhDAykbBxORphTsqKcySIf
Z9GN+IBE8dujqGPvAcBdH/7G0sjexgV4IPchsCO9LPYYaJr0MrPaRdv+L4eJB8kfJHz/MV/mxQk4
Jjwq/8VBksxQTco39pNPkGJcgI0+erMT6YHwA6LzPKe/N7VCUQ5pHdHHTxFGu5gdWuvzI+osLtOB
P5Pwm2tMVXLYsaP3eXflGL9gRKKLSOSfXVdu5ljdScOGu/ogRcJjRLI2EUkOcOnVZYn0h0zNKiA0
hSWU/vBvVO1M4mmz/Flv66mjNR2nLhx3LypHPoFxonT3ap3ck1/EammG3d4P5st+mX4u6bZY1gIa
SjMexhOvwTXuGSuVCVaLrgqA/HmwE5jLc04Jfq054tlhpocDSCNdYoBvjXo9Oj0VjowVMh5lt4AJ
hP6KyIlR3/Opr34yBNdMrgdBVxETuf+jGbvg3dUoKj33rKCh4kkh+nMyrImp+VJpVccDdGBFs2Ui
/nMG6VBs85WlDQJBZSNFXQy64Ae5wOPR22UyqpO4HR9WLnsX1dd3MRfn/EBBd1Y8IdHB+gny9dyL
40ICIadX3/SHZHfFAxFfKH7BS+hhOFesGP6wsQryjkHn6+nuAVxeYdqz0BNYubZSH/pMH0Rt4Ugz
1yFW2t6//aTwakAE7AXfJJUudk5faIn+ngYpvjwY+32eN8nlcnEz0Wmmd6uF3DniYZJkTk2uMqnW
LOJavAoAce3HIg1sOOuYBsSWKsP1ktOf/YWG0/FhV5eZPmJVSUfCmd1waKJ1iThFiVx+Ui2nOq7b
xFfcpuEXTCs8+ZQfNTbVA7mw7sgg1Ta2gjfPKjE58s8STaUY7Ybtdama34hqvJ3UAd3u94HxKmbZ
+siTZQM72nAOAdc5ntQVHDVu0e9YH7O04Dc1FfM0RflajDx4mw/7i8Y9gOAdsvbdPsBYv0aP/idP
GqOC4/pV2nMTDW4cLLbG/HL1wrUWxes938tthhCXcfoQknlqklaTtRn7J9W3H1JNqWK8bGrec3lI
NKu7enkI3NQi4pXOzujtx/TTQzK5uzw0pnHgPfHa+CHcI+LsDWltbHtBIEsUoOKojDniwuc6rKqf
E2F1J4OjvSL2fjjwI34QUTkUGHfKsaLtAm1Vsr1RcYzDnthvGWi42ctEBgYYir7fHqGRnXC6owCu
BLf82nMw4diDZB1dNNQkhApqeODPRwqrpuM34+sMvQh62ym+s9R2P8mGEl8EqFAsggSwYQz6y9R7
BpX8Rf3CtabinYsAlrCiNxaNlfWoO3Ud5lxeUnbY6adwYzQEeTDNa8CWIbpitLNE/yXcyCKPbf4p
jkoFlC/ZNK33J/nFexQ4nI7NJP/Y21pJIeAy1g/YJmzD4rPGl18c3YdA5CZMiA3ory5FMZtlHVjQ
/vchI5IdGFzBsuq5Ckdt5GGl73F+3ve6/rqzewopbwcPAv91OS7+XsJah2OF7dMCex+4zJ6Qjs8L
a9e0Fgtz7+LjqFg3PCqoMlQhHl6jq6+k363YzqnQ5DhzZJLJZChzLOXtlJprBVEomktmjb2kMyrK
XzjFx7cGG7HN2AMyrfzKAjJgkJ36IfvYC3+7doUUaLwPRNh6SaPgWcgPFv6iF0n4bc8H+eDzbiRv
lHeAYB8C0v1hXc+cODRdKhME5Rn4Zz5erD7t70XVJU68k+yjRjE+2nOx8hDe8ZHSOg1M4mkACFmG
A0uGOIaUXLttqnPaNzJ6On9hA/nAg9Yt4gRlfPHy7OHEYwpp4w3xFTHei+Y0xQ8PKNF6nbtmkgv3
4dbemXGwoE8xhvBOSmC04TqmrOHFSWkKjATkslrQmlVyVjOlV5Mh8TF63qG5Ts5ShT41yf3PsSGw
ytJZcbMjBuShUDLQxo+KqKDkrlO8yz01G8jC/BBp/6gmrLJrslIixAJ0ZE90Y08rrkHsUZ+BoBZF
+6j5yopLC1SpyAzJdxo2npkEYD4iuGXpgYopLlDw6uHOB4XT+wpoA9DRDRIlLfgtaP0IYtFNNxE1
lPfJlQHLPW6TvgdoIj9URM57Gw5xMJNYdU645Y0xCYAgtZnRqKrYjcL/uQHC3fveizujOOXHwHp5
q14s+03A09H3dda/kE47fVcFJg17qTSrH/DL1ymrBZ0l5OPUjFt34kZlr25xnPPHc1PezzQSicYW
poXxGthygvwPGqN/hER9Nly+3ZfcWoiUqwVa1tmI99gtExoF3hOj2wVBcitzhEDne7uSo+TOfcWU
FlBDtfhY2zQ4jRYMu3tiQucipXfCnKKh/lzak4e8EFP6FvEu2wPGfHSKt5zUQCLNxZCuY5GItIE2
z0JXWC330N/UIJuKjiXjKQBbOtMtazykRqcMQqkGphDs7NBCIKx7f30+QP1VqOztRp8zoia5McFC
4CSDVVJTNXtgZ4OMAeQFP6jTemsashz7/02C5R0gDdp+1n97rNFxsQKeUwX7likovqiz1DIP9kkq
nJP1otMIEQDOhKUAkF/EAaj2DAcH6zCGXM3sjXhS4GmVreXCVaOXceZiKqrA58wolb4GmP2mV6oB
ThW5F4AEoPRDw+1ljT9PQMGgCPFvy19AkTL+7VZ6YzMQxYG33svcqe+gQF9CPvxAknDKkE7nv5Cs
SSlezq0hRTiwTxoOQqxRA4pCwa7YjaMgnZyQ37A76zC/OrG2Gu3zRkYwYC8TalHyr9SWsHqtDD76
ZISz9Ksp3cxq3UkPR+ElU/cDx3oYd8pB+r8s7T56GT4daF3aW5FwwuJCteBD8Ri3sSDenR/jF57a
S1OhXYxaTPqG3t65wzBI5ZZocAtsPQF7v3YWQXMwUF1d4GuR4JA8OFJeCItE4SO1NTditQuqXrCA
Tiy3pPLPKgbxR/9fuk2VMEB7oDCWmPzFC4Mda8rVe+yWMr/13QlLAb4p1oHAxdxmaMvIBfqyXis+
J2U1kv2MJjRcPP1lZeTHcuO0YWXp8f5iKZrPq4ngcfi3AgCQ4S+O6WeSgDwaaAoC97iwts+YCKQj
F3ADoN3rLk3BJiDE1VxE3r1HaHr+ZFLhqBno+NJ36E78rV5y2GzXaqHMG1t9tUUzDUm6Mym0yPwj
PyokICw/24ETuL/2EixEFwqlXib/my+UKMMbMPtm2Apx/Z+DFn2iIG1bY5aNnlqpTzffL7qM3583
zXdSxVF7hem0kvCTlORdCgwXbwLjqyOcOmGHOXLCUBYfmd3E9n8TojZIvKorFDVFp83DbgRxBtGd
ybNYqotwDEMX0saI/UYGnrGIdHzQYwnFo9wBCuyB4cc+xNWx8ha5JbMUL+dt1ajOIj3QuSALD3g2
UZB8ciAr8MwDWGU1ZhcDhQuCnHBI2KuX/C+5cu0/UzSWGS1xd4GGGeTkw5eOzFt0yLzoKOxv5eMt
2OSvue3bOZVg6Iok18q0BidmD6s9zoJHL/Yk7D4JbcigTpyGIMyUkXcsINQav1vkUlEmAFm+I2Xf
s0ur1MrH/965ouekAz8G15X2/7aPk6IhkW2rJLODoF0B79oXourKGKeNnitqAFRqARfNT339nP9Q
/nez1nvFWIRC52uVP8mFMKb1zsDfyYGwPvtUG74zznYC6Wcj+9lf35EhcJGSdwEJwfBOIz5dKjlR
hhF8hIqQFVTso3NQRQBXZ3yp6urtWpJ+h8CLRwbZXLBqHxfodtaggILBnjqPsvcZmNhEvY9t6vHB
8GZ7IywiTYQzDLhmXo814a5hc4n+v9/RjDiFpKfKCqTytL9Ld5cTcRctmND5QaT0W7opPXA+8+FO
57n8SHjsfdPoJjz9hKrUJgVdMY86YuDPpNT4MeG7mFzGfXDm6LsP70qTt7Ga4Z32/a7y81HVTwaW
HAkbaruDgmPHjoRw1Nh4u5/4LEbIIunhAJ75KVEsBNhfaTPwfUER6c94McrhblIYhmIpsMg4dhTS
l96tRnL9wISkEmFBIY9xnwS4er50hUzJbPdROFpNgcRlwGpksEDeVsMrLIKWpONFkslfgBuMKtm6
5HG0HMkXKkfLgUtW4Dh3jLxivJUrJzm9esO+quo8mMpY+eKL0Rp4Ltt5wbKq5bYZwsuvvfSGqWu8
AfJm+3uBHWOm3on1rbl5EcHmCPyRa8QlACCkQoXHSKpOcNMIvPRqb0wGlrmVdx+4Z4Iiy4eJvtSm
i0RthHy5DIRS7J7brNG4GxWpVC7yYvTjched7aCv65Zd0RYfwjoL8FW5UW1oLiH/3fg4POSgyYvG
knlxfJ3zTiv0yR0G3BhT4K88zDkkw91zvPXngdhfLtYwbPnGhtxAew/Cq6QBqlV55xxZXf1xEMGT
GVSzViuZLtR33lJMn5bDbNFERA73VHiZQ4QeHxWD6pDs3OjB3G1e8FAiYDdm2iEDh2YgVTnlHdI6
X9nFQF9mDSry4B1P3BH1/uK12MX/oOesMkyo6p9H1jH/rPVUl9M9sGKQeDoVIMrn5w4NfeTwJa2a
+/0hYg2vmbgj9TlHLBGBm5RagY7g7BIzTaGo18vDin4alWNCUAgqZPx5tCWCP4tfX6uO0/k+veDZ
tXdAlRjYHb4HVxV/5NoorDC361k8V+xpu6A9OV1LoAERBG3CgtDCN7/a2frHwmdhnxL+Xx9CSXxX
d/6DUfp9pHqh1PSI+4B93JnDQLjajT8NddUBLRxrt6C7UVzZ+2hV087RskJ9gXnd7LPbi9WWA2PW
ft7cm6oYq7ZRXoEgvKEDcOTSlfUd9Ff2vCLWnlusyIaDlpdlyfgLjfE+bNug6tZI3VKDnXV/ZS10
JX1wpBxQ4aP7xvAhDcfqqNkxmoYYGWvoxYbQw7RM8mw6Q4coPOpvawaml1MtMQqhbGMfCn94ES3Q
zfGC0dJf66LKZ3KLIOIP4pYhVkv25NjjmNlXTxBJZtUzyQJN/Hof32Fgs3DOPfKGvQYduZBEWZLr
5FUFSaopm9XWdoPuiYNjpU3sBujySQ3x6d0h9k9Ij4j1lXrntn4XT5qG8K2Df05liDfSyxV5P9Ph
NCMVOSaGS9Ijs6Pm+zDJiq/R+AXGhfWV+j3v8nistKVKoMVVxI+6jv2DE5SomvOvOSjMSO/4IAuv
G8PAj/D3plpHLkKdeC+WyIm5C5D2AZlSAFjR18VggPTfFCogAMW9tIRH0SDc+AMOc3ZO/3dBHBzA
lf3xXFzMlY+WtVAFH/zBHfzWRkiSCHPqltfCnz7TESF6zA8KwkSY1SfCFPebPfkR790MbEHZCnnB
jY8aOGNoJ0tv8/cv8+6owz22cx7FkKY+qtbjzpR8DSqAu+aNbeoU2tZMnzwe9Fpngq+1UugtxtlQ
izrTZYEjFtLYT1Zs5qx+HbAq+oPSo4nwy44/w7fjao6T7ndETv53//yinz0/34Iq2Sia3RkcW9Xg
zGRpFDEl7lby+6/FxiXzhU8jzSwaFDqTHnV88BaSpriZ4LphgNlI4/9LwcuE6SkbwoqU9VylLWWx
o/pS8MeUrl6DINaK022gDAuM4C6Nf53+92I1NfUJymE/S3fXzOO36Olp5m1wBeYNKZWRhyLjTrFy
wD0n4WkLo3fbxbaKuFerfteEmqgvhLjut2iLs4UpbeA07/BmZoK2XIWF3QAWNLG3evz+4vrPbySW
63PaoQeXysdoRKFEZg+lnzN7bqFPjJVTUyhSu2ZgFMRSOLVTEtnkmL9mKJY7KqgDyaINWNq2bFTE
GUFYwkExvxOiyRlrWXyYOZF/p/wuhZo/6dp3Sh+EA33ihJzDjAroTMEN/nDu5dgmQrHhPM8j63WN
A+vbiCZvW3cMLl2AiiLGmcB2/AtZRoewUezZmNq9bK5hpqC50v5YM+Gt2uyaNhL4937vZmhlUo5g
OXP7LcatpWCMqPRs5YlMaSIE2HXtpjFLPWjMlk8gmuWx/R3SG5llWU3sq359I0PbYOsyAtjFthiP
8eCnYiGSlnUoVCcHPJ1KgzWQObmLbao20ttv9pRH66c7sujQ//Pghw6m60mpQsP4TRXxqCluM9X3
iLTlE+l3bvcMlvLxtnj2o37Izt4ui9ISN8FjV5p+/UJTPB9WNuJb/A19YrO4bMbZWNAKr5/lKgrp
UcoycgmxTJpwypoGH+c147cSPqxbfAO32bYXCL1cHlq/2RjkY0nAVpjUQbFBN6DML2j1mmWcdPPi
yoqs5ygRbbGb/ZWzhfSdxTkwna4ILKmyumL6nVt6kICvDclHYC8OWP1lfJ5SxXxzpBB7SiQ5LadW
V2HbfJHSeXo/RX+KvVzO5uxY7OtXNVY85uXsGQS086rSQbYUPiTzyW6B/H9o38/6L9IYdiVAmLlC
25IlHK/9z8TQlgzD3hgB32I6F8kqjiCcvJWPjvGEIiOZeDz/OnvwrYh5HTEGd0bOek1GMfApXne6
v+Dk8F7rXTjnffrpEfqnKAKLeyQ5HjmxnddLqjlvsnxoyZAVcdlPR+UM6+TxR1Da0NHFubWeO8Xo
PPvHvoEPh8Wisu92waX2jUVEaFXYFdw6S/vuecznLZaD4XHKvr42dakqRg7GsXp3wL7VKOAwHz87
hvCLwNPbh1F5Hpzmu71MLsMNcXickhpnfSY2t5d/0TATOWAKa0JO2to5GqWrnq5hra8y5L+u3Pz2
+oKVvCNxo1TIjYJAHxNVgirqOZ5Gg5p4EgddazWrKaW+Q19LVy3PqWx6QwXUZK7bCYWDndgJtlvj
s3osjsBg6nt6/xs7RE3+uLxbtf13YdmnXx4ox/cBXKPl1dTM5qmVj0ZqBlxmHz0skjz5jOMyenqj
e+6/UPRBz/kZjfSYw3P4P2C6tX6VCH7D7mlgoBcZaJzq14uhPT30Fdjnua2eB9/+cRDWHFlAYu6u
gHlX1l/S65xAxUkmFxZRB4xyO5mPRfdLXsavUSNmTOoHVFZpWa74jgD+aBTU1kMMzFSrA9Tc0lL5
GHjn1KGNsVXUc5JrfnZo5xH2HnkjUMHZILCuSMf2d6TRONnhvuZPvWTKxKs7o6ALqagJ0OHFnCnn
Q4wbdvmeMPQYQHR3ZCVBEt4opPFiuGqO5H5Uq+COgh6dwn2acZVKtM7JNJ4ejdqIeKmpnvCbcQBO
4CJDWvZ89/qnV7IKI8yVmtLw4He0v/QstDQdJ2R2aoh+7DHSfrzE+uzdayWmSMIiJ4LUwAaY03Sm
yOMkqQLeERymnKvCpmQoxuHc2hY/NWPhGRpZmpEy9I4Tw/gRfqAtcMO2fzvthBM6iG031Z8Dpxna
s1RBFyYe5ot9fFftACrYNxkZ0Xm22eGHb9ONaUea2w0iREfITJwcKusUkSJCl9Y1GwRsL+tQzkLs
UFIurVCYp/EsuT8iuwZzvtlRTqBLeXlv9SBT9O77IAlHVUHTLmmvug0sJUk+RgxOtHyjOhuW0/6q
C98zJjojl1p9szl42ZEUlqCysY8t3aDD+OhsQjIHXAmpYuPQGzxKUMgR3ykkCBTuekKElgGAz2dk
YDVmJmgxTQzK+PiU8RUyBjoCfEfe9aqPEKIxRRMLZqm6/tG3rFjYJ327GJSpFCUdYDIJ/BprY4zs
dVrM42jnG2cb+9nM3skdUL9aSsutyiw3MGj8rGaO5YwH1ZcNCVFXu9f7cIRv1DpsiGAbPTYAl49W
CFFLCnko9bQwh1+qPjonCXZbF411H5+35KE7Mh9Cex6QaX5eq6gXSrJi46npEzySxC8ED79TrViQ
PxxwyWh1VH2jZxydxIOADB6tdTAxgguz5tAHvXJpLkE2kx75z/0krXgydwDRHYjxlzpLpqOn0Uiv
tZtF0UjCguBmLyRFPF++OeZiXScKvKapqLkFTp64PXDJgOs8PbTlK0ME+knDijpslhzTuURo/c62
f/LOfunpkPFSwN+/nT2KIcf5L/r5EFWbniTDsl3ieO2aWKkb0X9uBo55vJZCq7B8ONFZ0tn5qCs9
aum7kDIGQLL3MbVT3FwmuFR7By2j8AV9S1/Cp8ZkyGmSzyph6K+rjIRYVRhYK7VQqcTt9Whn/QWV
wOERUX2TvNJJ6Ojdfj2ZO8cxalUTez32/JjYnnYYo0W8sSnUucSSpZln5Qgjwo9kzjf1VhlaUv/c
2Ox+1wzoj1u1IpsfCN80cjQgytToYLcBc11sM4z0GHY5hZMvVxSYpb9wAaB5ZznDNbM1WbkTcYMX
fdNH0vo+Di8CLM3SFPo7shXklzYf7FFS1gSkXyP4i66+3OnqvBlyOKi1XohAXZK3Zfc4HjeAUG9s
LSCZ7MBK88G9SuDJLlht0+m8zKc4wy+sJuc0mnvmpBrwr7Fr3WcjvFxyb8HGK/c82iYSlw7vBGNq
CANf5wcNpRRVj86pWXPgJ2oX7jPVrg9sMtxuwQLxDi85dFLIn5EYTHsncpdPOMEFfqD5Lp5GwJed
/LyKyDZ0LIKnJRUKZeH/2sK4Ipc8zY0HrSwSwfTzEuBnyYWmpRAjlnvGs6qeBjf7rw/Dcf3CWCc6
dqaXFTbOvW6BexLRq9vdFSWVHJTy3DfQZJt5cHyBl7qef3jWqZ0F+fGyyxbmkswxYLs5TC21eLGA
v5r+Pj3gvBrsQ4cXhyGMt2Kr3DJPL+kveczkkvBDXAmJHNKIezURlnzLxjbRbEZDf/8KN8o7auhS
XOA8+JZepow2bUigVxzzzRaWanvm8m/2B76GQFyue4hVrdL6gXdcOKpfXQC8qnbZghfmhLuMfNAJ
a0QqXMbVII826oHIj/ufaSsh3ILeHcdhzUV+GHtx21kOKp7y/vfqdtOUx4rJQFzAuAMnYPKNlymd
DNuf5Mssny+GIZ3v0F7o0MR+m0LGdQ4vIy68rwHQj7kI4sfFn5oUDcVkvpC6ct6ei4NfmMwEX1I5
+yJbwjFD6Qr4QPKCXh+854IatshWli9483Fe6MshjZu4UYOJxkEw2tukkxCqR2vxs/U1929C4W8p
vsURPp/TJhPDzIoFWuzj36AYoIiHp9AdhOyBg1O9E2dGGPpmxG/lHxtODFLnJHk2Lazd3/38HUt1
msew5ozebMPDN7IhPtFU0MDZG9AiZC/kil5cF4rFpyhsYeiK54o4FUqx/pAi2gvn6i/oUjnhu7A4
9/pVI7wjk1fCXbaYTe0PFhTq0OTLxFY1Mjnwo8ed5z5LI8p0mKkcuEDcK1Ftegu53MTireNbxona
3p3CN7Unr67k2rJG+jwk6pVA0SCHF4fEkKf2s7lHaws28j1jRKgd0g2mdtHRanqbqNjxuKEJuvXp
UIZSm8lpLOm9hNzrJTXdvlfqHYaPf5MBhpy+FtnyUgFRq5Si7BtK1A0xSkTmz3SiiZC7m0a2oSt+
aiK5SrNBWVgCdcnHQHsceJ1QGWcFnl7F11fuNHMmdEc49pnu+H4UmSh6sgdxrB07G3/YUB7Y0eOJ
GrKUYNPjMvwm+PGeZjRd54XK08/brKQXFLIsU61dv2FSZ4vv/xLkRHD6RePetiRs6MTkxRKHZyqo
pJP8xkULfQT2hiQYo0VJiS9Sx6KGWBwHQX9quHUOl9wC6NYzyR01SAfispr6TCu4p9RbQRrjg8Ak
ea4IxevXqGjnh8dF+3XohO5W2P6ccWgRdJO7Bngk+zYpVFFcWD6kTe+e8tgcJkOsTCPlEjR586kt
AzRNf+sg4+6CcTKl9GHQB0yeOK3tYUqhApCH9ZEcX7xRWL2B3vjdaOopTH7eFrnR6KEXuBdtfBoj
erJR4DXTa93xmaJwy6V1/hhNNaGfLPGpFC6Wgzu+5h7dr4Sh0ov5bNmfLowq/cOuWrkUN3mSIV8x
v/GbJLcSsNcL4KHlX5NMuLHr3J8rZMB9RSpY9n7SZISzn75dZ9GwVSApMqDxZSoYPtqhMCIY33BJ
xUR0RbOn7DSILqBOYydT6T35PEbiPEd1+C06XIsL4CVCKsvn8mb/KGiz2cxt+kFaeaiMAf1C4eRz
AadZjNR/U2ZsCvzte8sOm/udXYzcMItSobtoW2dvzy+JoamBq0m90d/kwexPy+fJg6COAchah1hj
pNL/yZ7UU0TThaL+PO2w/M0jnarw/J5OtmXLBN+2/InoFRNAE7rWL+fzisGUw8ZcER/l0KHnvW8/
e5xnHo5WMFakj5nXTNbwIogFFHBEW+eO5QJZ2P3BeDvVSuJxjAkn7dIo0YVJXUYW8GoaW59Y18mo
6Ry2UGBgMT1IN+0eZJPnvQvsJygZoOZjEgDrHE7SMTnyocZfGrTcmHqw/Y5zEkeiAjmElad5KJiM
D4f2P7IejjQM+z5TKFKydG48SbTuN/qHqRbpXzBaO2NJxMs0OfcT4FUhqFGiE7LQ2yOsiRgzqnz1
MGPAhxuHEk2IfV/cPqsKdptFUvz5sK3rhqkV/N/J6/I/OiNdM93swGIDcd0+VgazZyjBl16HiAoj
o1NMvILLn1IwLRXgH6iRDG2MBJB9nbFVI5ITUSXSLPT9AJsdIauGvP+2Rn3v5JA2jTa9gPBvDtZl
1C0m1LE54c+XDmaC0ULcrgbUb8Kffx/SluNBANc6JTqYtfCwezm6sdJdamAZk45zLaEE+bdxj4uK
ZYyb9VZOHjQ00jE8qFxj+uuRiBXode9CLNo7g42VJk766mG5akllyfWUj1Z96BsygLtxfMjbd6et
E6ViRLVzROE073N4owjNBt6sozm4p8X+bw0tXI8ENtZVqPKuE2q2yl8kRrPIfu25SX82NgMeBdN5
acQPG8vt/XSEoDOP0o4ElmYWnWkGKrlc41bXUoelNQ+mHC9HXodT9gWsXeci6VwMebbd8XVHzJiT
JvjM4ZohD3eElYYs8lRmYE+t1DsI73XOfLCyLvr8HY5KdYyVEaz3hEn3mYij9kNZZxMXt0gBtMtp
ekbVvxQK/KisB2WMoRo8sq1eJbshwj8A54hFUaarUvvHi+mblrKfO0MqNeRP0bYBPjxJQNgeZKVt
dfZECNxWBJo8e6dXQGJbGWWcSaOFft7FwITxFRUYPBReoyH6KKOw01YMpk1CxKCPmKH7eck8sfpF
5fMuY2kIZEogJfzTzkLhopfW4XuC2CDAslQGoi38V7WER0FhY23//AFLIwLC+U29eQVtj/UP653a
61imrsPNclw5838H4KYCTVARP299rqBOKkjFaxQoA5DL2lQX2EW1HpFF80PrDHX/TmnsjpQbthid
s7+gayDyjn+Tf/674khPTW2T7W3PBgJPqxQeTI8DJ92G+0tAG5O+plkwKgWfo9038zaXnlEtfaav
ZfsFp2FP/jNB/pDinJD+ypO8GRZ/NUt2AyFTcR1lai00EhEE5ADE9bbdkA03LR+A85Riyp1ZL7uP
ZWukMKgcn3s17WRcAORaWbnsCIA+deWeF+K1/U0aRtuingFlWX5Z00esxYrgyL8OaB+aSaWJmvod
DdI3MiOrArLYyaj9wp/5Eff5b+zdDlzHFuFu+plRNo4zJoNXrCzGGyA4VUEXxYRw0oM/F4G0LDIl
A/nBVubCCu+mGuYqE//o86M1pC2FpFyhc0nnXcETmTlcdXzgzsPBSzNY7IzLn9h6QWsVkwLfC/lR
iqsTPAxz5YP16/sSpCO9nuTYkhqIaSTOZa+eF+omJUzCUuL+gIp3WucZusU4Dt5yoWDNa+RTvLLP
sNTMPJkapqVMqAuDscbguzrQnp5tMfQl+pvzejQa67jWCynCQrYESN41iIxYu4R6UqANgpZuiqUB
77dZgjJfGaeq4+JUTo0tjWcXTFlpD6edcNwE9s4Ye5qwgm7a8KWLufPubL9JkY6LFQ2XVkQRy7xd
Sti/lt+VmRZbf6POVhZ8rb+NyN6P9o1Fkk3BvbWm22zh8EAJ84s1413/wrXs3NitVjz372jArzIh
fOw6CObOByELDpxjBPUEO7l7XWytH0iGcMbZD8tCKhZ/oti5PGrC2CV3wrW8zTV8IAHg3RJ8gSGF
I5JxJXIu08A4zzedAiGz15PlMTkw8nD5rzZ/5wpQ35i1a4sHQVMy3YKH/t/f65zdyQED/L0elEYd
dzaUNTmCdcJghvsgy6cUM1HzaBiK7GRSy7I575bAjjvnt8BMrbZQ4gUuTZ/PvESu/0OEpBVhiIh7
BpE7LxDCjhNdRDZa5OQuDECsq0xTgzK7Bgn3F6tgafn2AuYDpuBoVsg3nwgModCq9VzB8KnMrAhs
FLXYnv+/N16y9gSS0dq86w8f7AfzyR51iRe2ZOSerXPr1BWHLwi/Wy3Pp/BtYHiD1Q8NqoIK1rhh
cTmtocdNzMKq+vTNnhZm+j0ju5y84DLxOzPjPN/WQ00FAlpzmzuJgRdzH8OIehynLUdNSa5K2tA4
JoM1xAFFgSMk5xIDdrU9XTIvCZEupqfxdhDFyF+oXweX+fkGUMBkFq3QP2u8qsE1wl189jP8NwDp
hdeP04DaSPZqrmv0MrKubxKv1fNre2MR2PE+VEGbwf2/igCR9u9sRwk8VSqFMlyU5pHzvS1AyJZm
LriyBPngufVqtuTl8Tqve9mg/i6ktJsjzDC9sZ6qMsS+b62/JFDeZYlOt4Zkpn9B+crCpzr1yyjP
mawMYegEaWFxZJSq6i2sXdI2s9g8TocGc7LzZEg7ZpXcpOge5A0kErYeEjS4rZYXLDCgy1kJmk0h
andqtGioGFfjCHOQPvpMZrC7riIvVrx46T4TQUDmZPpYYu4jkm5xIbA12eS2c3VNnBldkFP29HFc
oVyZJGFNvNsDFLZq9Wa5TaGPe3TNwwgVkg4MIHjVURf3nD39LS2Zn0yQVOfQGoWHX9O1r05shg3l
knyy5O5jA45/QZHiOlWBmzUyZlwxFKcqlUOqDpcQ/sYWTVpxEj6nwiArfPB99rogP9G79A2uRUgE
M35iS8qZc+aDQvgPeHp6wVV0y4fcDqX0jXJwZ+q1DR2o0rOcWoRkP6RkSkeY7Emh5sbV4aBFkDfV
4Fqrw734r7G7aaoZC7zg+yPM/vwGWT0x/W3bQeRVVnogqZYEa8NFhfagqY1UBvzfmTBYWx3jS7Tl
E0OvQJrEoeGQtGVIwhS+VszKEQBL3hGl/8niIOTewA+nTnMWfRPHz3tsnJL4UJs3D8L7BtH/sTAF
JCPp2NE1KpBVYL4MEyXcC8/Wn10u0zs8hUME8z9SrbaQgP+h4ezI9xqK1HaO5Cq6DzUjAV10jzfJ
egmNYYDr3Axw6Vhhb33J7MpO1+hxWPPlew6qiv0iI3pXfyQA3atz5+R37HfVKmRuXvQEvQ9rpjK5
Hc9C3GyT08C8y2sK/q9owx0aJX9k2Hl9/0THt65Uo6CdS3otzuNyR4mFALaAs/KUK6qNyEstzZo5
AuOOKE4+Rh+yXCqbgFvknnDofOM3bjEL1PEeJOxSS3hnsIgeDEzAKbl+VzOj55HJtsKiI1aHYHMq
/r06aj0BCtnVCxCGPRQ+4YvT7RuX3n8TCUQZLY/F0GHhW3PrbFgmuYb7kQ/CGcJaCgSm8sDaGirA
8qw2HZfIcTI68s1FdWx24R6Ds9Ukf45rwq+Br+PMZy2tZGMeEc2GWH5liA2hIfrWJmiCuUtj1+II
HvMxPR8BAKpfwqfZdMRZk7hAEdGOyvcpxfB+KxM5ecpwm0QY1pPS2ItPbnC3T0QGHi5z0HTQlmaI
gcb+FBV1evd09FmlCzkQnVuDeL0wh3tWQgWkWkgqnLmGrYi+uVatqSLn0L0u+5qQcok0R8w/Fbvi
DPaM3bVtWfiU7bmeu4PMVVjmUnvI8Af0QrSmKC3veqwHAuPT7PwwizDScKcuR51juItpUTxI3nIV
LrYxjBhDwHw+8hSzcO5q1INSeY4sKaSYIzzLyES77eFDyOeeHT9Cc6H5JOrxlp9MWd8OlDMXqWvW
SPNHC4siNiEEPi+RTT+aRwTHrxv93U2zuW4dTPByUtE29vL1TKKHjzJtkuHgpxd50IYnXUUx3kLI
l+zd0nT0OHnIhT8UWmc/BFuGnhQ88djeYZwULS/aW7qw4EMc4hb3KxBY+CjcELXkHdwRHQuxqaK/
sif1rliTB9pfjbGikBiTzzwgDPuK2Gw8DwVBHpUGtaA0Dtcy9TQZkRGV6O0v5YKkypdksDtp9WX1
R0NKtGVe1FEsMA70QxRg+EOSfqlgf5T6Wo8DEdzqsinU8qUElyOOJomq+2uE13j4q8ljSz4acB7x
L4E34ZFOx2XSZBOfbD9ASs1qCIiFeUa5sEqfPHg2c9Tpt8085vg96mpAjflBHfhEgOr0Ql1QdCr5
K/PbCbR4+tyxZYag9av51yVmEfv6gqDl5aRJslat6gXdxzIMcUYIGYvwCpYZUHiRwr+zfycW4Gii
7iixWtqTIiEJl73KgbktF1Rm0maDxzu2hM+rPJoFByTMNRAZuMgOk2ANHzN8iAppa55cF4qhkeRI
eJjPNa7Gz7wdd8l5uuIzQ59OkHJiwJ3ln0QeVupY2Go4dl7MCYN8z1yi12wJL3LiQ7eCd2VFNAEM
0K2qTui66MK68pg8OL/7hyI8Zi2LLB907HvtOnw6V2EYRcvgg+A6tyrxJSt64hxS2kVj+73N6iFU
mHsxP5G0LNwgGPl/2PabWl14G7AAViovZ2ZWXedaxp6lBOQq21QNp984wPzH17h7VDweEZowBpY8
X2nr9gAUq3o3Nw6YuZeU6hcr87Pj/zuMJm+8xJ7pveVZQhM7BPWRL32Cg5pU8ksOGBRDH32ivq0L
B565IwAhYy5CkTBfmaKWGdIazcf2kAeHKGP1gnutuVLCozKLpQw/cKAHmGJBNKL4XMuYILmV+16o
np+T8umzPMchcYoF23+j2x3cWzQIj4RQdJ75+V5gLOL4hFCp+7hxP0mFIpmH/Mx5HdDTR+txZtiv
F7A4ZcUBQRP3pnY5IuFqObKPhbJ/Y0ybc5ub7IMKVRdlX9dRm5LOJukkzowO3Mfh9RLkQh5s3giO
bDYNT5klCgHL39YZduRIEinBlpkWGiIbFVdjstKeS/tiv3wwfgl5vxr+KyNWmZyIyY1Fuh9YnX8x
zXwDd0VSvL1h3CA+D0txt119ZXXgXlz46UdnPqUA2zW6gr5WNbWF8arUsxxFgZCWLlFgqNlSAkpD
uqJwLF9avBoRnGoOMH9HgFxZhysckztc0tEbvKij9HduzIL06U/0b6PqkyRMfrLuKefM1gs/RNDD
MwqYYLOJkNm8BIGb6yZLh7qO0/vcm+9jsy7qOpFYYKOTpGDtp36iY4rORgygEQplpIdjmmJJQtZc
LD1fNfnsiLZuIgL/jVhnrkPJGvJgr+wolziKItAIrL3H4DHHC0rI3RGXqGyk5UCL+tDjSr3Yuhk/
wu0PLzQ5KeJLYN0HPtoV8ZZXWM+Po0Xg+bW9ajluSXRcJum9VBBr2GdXuW1SdLJGeioJcNJvRGXv
XxmLVupAPRiZw5tLZV2ri/5P9fwfy2KWAM+EU1O3/CEQnw5zcLRhmaGhDjxV4T0Mg3m8CltaUkLI
E/oh1lSgpuCKQulKm0YqZhV6TfW9jrtXOpKkHw8bbabFyRVurOrGLPdioK8/qJA6Q7/QQSLSdKMQ
yojuG6XBhHnLIRWsRYf87QMo7LYxpJzpJRBykk9kO/JIQ/PG9nSTd4lgbvr2V5NIZSdwoZAnDjfk
M6n0CoAxetiIP1GPp/h4Yj95sc2fSaCHmkXcK01riX2x8mpz2PLODqSw0ePg0LCQbf2PyRa3QAqp
7+/vmXnDONk9PrDXGn/ZCDOj7jVoP7UNulhDVqgotUyvPaYp3/fVe36g3hKHHNg32umAU6AbuKaL
S9BMM/fnGL3FkKrS5h5xF8tdycol9oAv8R/a1UTIkpWu/7pRMUpCsX9RyXi2JFBykhi55rVoC1jI
3Z6a/aVcFDmel5eNbI4SsJIvMzaymxeb43xCplE7agW9xPiyfu6xxIt+0eFdsqDNI3slIrEfQsjT
w7/kUR+MvwMFV+P67xXtZlAg5dbax9liChfe/YeMXyVynWTEVhkQndMVtINOrq/BaForYrbCWFca
gK70wCDsZFt1U4VQb3JEKuCJTLRuzdTmmrTO7AeEHmKcAQbGXhIYGXPj5KeS4q0bBBXLedBDDptB
FXBJahDWWseCnudRyPKsnwPXxz7NNLU44uTxCFPRQISfQE5yAYd5k6qETvUcKkrWiOsLaaVcWcPw
u9wUXgxiWbZEnTQPKSAY72CbCpR3HnpUONGj6wTyCKeS7a+636URKT2o+v2yCEGwspetLlpG4Bra
hphNGtCSYgNuWR2EpVBzs5GCNYOkjv2PlpM14yXcDaMpncvDBcXC6WZA/IrlKseXJVBEcWLHj7rg
p5xbjz6aUsvZHtFKBRrnbj1bZd2sZiDzuWm4ADhXdZz6yUMAl8k2DDUz71WuhI0dxFYs3/7n5+9G
coJBGWIDXgmNfrJZmT2vTx+liFnclVoCGKBiUWC67/mco9TyGLn89Jwzoyza1jsbgXeTJpDRczgH
kzbqE7aBTItxFH3kZGpY744WgcJk2MOhGisnO1n+vhes5daTM6HTnaQLUNVe1lvkOKgqzDKySSto
NfTYcAHd6KmmBSygJQSqPOlnQFjqXn9VndZUCO53BoW/BAjGzP6gWqMRKuNgx9YBlikQapQWITx9
l2IDUs3evIJir1mbOqooyx1r9+Kf99LybW5ecS66Bp7sN309iRdoLCTA7GUAC4/+qNM2XE6gDP5m
juXMqOBL9I/QgHwP736Oaw2K9yGfB0zuhzSb2qAuf5rZD82EaHyRZhP+hHFYE3KSKljgXZZJEv49
CfoNNHZ5Eklczmlh/CeO+C0m91OY6jMPf/xh4SribCP5jNMvl3q3FGmXQXdQn1hswR/dCam0gi4i
kfSWY89dbX1T22rgrxf/KNMCoqXwY3L5edHz2HTasHiVH6tOUExWTqdPyk9SMJ3zLVgDum0Iq4dS
dpeV8F9GWPUsG0xsLJcKy8/fXj4xyr5UiAFozk5y7JVl5PtTtfY9d5uE29t1rZzmCOhWB0L3Q7py
9SBD0Pn3Z3jzWMkCWskiows8Mc2m/V7vgng577cLgXUZOMVt5RbgGstGF8jRfvCuCQQI1SUuMIdy
8WF46/aG1MjOlx/RvcGaJMGxi2G1HHWc9xoUafWZ+Eubz8fpnM6RtgQwl7xPZujGtKD+d2ftv9Ze
HpY9JvPlnw9rJz+6NMbosnMU5WWq2uZjRUHBDlepvBPkTn5cwwdBvJxZIRebmzcvau7W08kqdhcd
CDe582RztJ1fXxaZz4hiVNzU4LYn7XlmLqA01RJGbAHscdNuylEM4Vw6Tho1Y6s2MOV0jhzbfgnJ
H1ksrOjhjYKSpC4B0EppuopxPDZt+4l9/fNsfOeoRyW4opDzsPb85DTqCU5+IAQnccJExcneaX0a
lr+akRm/g3cqq74AG4jxUh6rjxwjAHp3RH+NGC423d6ww8IAsHAPMLdFwkTduxvPBaq68iRWI+zz
KPHwEtQqDZowN/8AAE6Y5m7ZEie8EkCQ4Hskcjgd76YbjOSTMDUFRrqJ/twNdcrV0kWxjFI7CoUP
IllBUfWBgRKniVTlf4SgZmzUWcXfWhc10neq7K2qgCcSr++GxO5UFTurTzSN0udIYVdTq246fKKC
EvfgKMXOwvaqDlUPnC2w6BdGlnbFH6O2U+nCbPxbUyQvh1pVZ6SSprXhCPLsMZUQSDShFrWFvqQb
oZuApv+cI/xiH4iAftmAMzRc8qn/ZWTLXF6jNmkwaw6+OTKhLFXa+fmvjIhchuz83o2fZWvANFaj
RfE6hddzZpWV6gAKJY4dHZC9kQM8bTLaLzZRX9dp6b1dPpIsx2i58e2HhTrO9+p0rt0jYJVnvEDa
KpPPsgJUVuGkVMzUQvwQcE7+aPJeHmkVl4GOeuJrB2afoBDH3tTZIv4iBgYqhi+pJ+hhMWvSjBn4
MmKuJ7094IIH+s3QzSIKSsYNxzhhBuUo0bvN5Fgl8K6DE02/P0RHaYIm8EWol4EUOdEF9Kxjn3o/
Il27os2ALkL051jXG+yoM4iAjPUjSp2C9PX+jOGewZomdZbgCQo2rqVUyTub4mEPMzonCwaoHcYi
39Tt3/YSFWsLXxF+gtvi39hMSiLmczdaINZmphyhDuCWnMrA6NpH57Yy7s/67NVnz+TGZLhfpvtP
rt69G+jyktsI0yHnOgQKLi+NmEg8KETLTaJ7J9bKXt5wLvykh7R/Kz7pM4cwxeF8YsWkCtULdim/
gZzbNPA9JbkNO6bfsXXE2pamb9h/kJRzmW2hHcTZXMPXXakwH6TwZici4cyg3EoHC1WbwO4KSi1h
x01aJKM/VL/txePLPrKw+OPjcg8MBw/KyKayLbZ7VmbfAUC8kjkHs0uBTjfcThaMUTucHMr7UBJe
FkTCWVDnGCh1+MYHpbPM9ct5G10SmXj9cDnGRTBbVGRUdtK5Lzsgws7xQYfxSiF6rau727x3l+2P
eH1ZsbAavD7RP43OjL+hk7ePmPHgEiSNznjX3W8V3EY2/Bo3qXqPsFGW7zxY36CzVwglTQjbt8CU
m/RdYn8RpO65TFdyeuBjMJX9ji06O3MBRzjLPojG5QrJuGOuKBJh+4T/aDV5yfqiRxT6A35UJ3N0
8MUFQSL35NvzDdv4xAmUDJAjHKj+MWlXReGEPtnXb/yg5eqAKmxoSlPSMmCwl8gkemRL1h0F+bXg
UKYcPfISgJgtmNkTE1+dnKl/cQEMoi7zkyfTcU43ZLGqW6DNEN5dTRdl2BtNpemd0ScuepSClZQZ
YzSIFW9Ae92XyK9tCmUvGK59BUttj7V9H5tSJxi8NXmYQCSngedKe0Ph07XhtgRTDEZCuJ545keb
zKdQhCUruwitwx2EXwSfA/CxmrYAzfttYsf1TxbV8So1ilsMBSJQ10MYkvpwrOJCeK3Za2xpnArG
jNZH/t+NCIQN7OYC59sAg4YbCYkD0zhwNgUvHJha6cKT3Bmc+J8smcmTxpdZ/tE477um32r9u3tB
rjoU8AIhRcOmmQd+HV3ZwxFD0MS7Cvq6v318ifjz2nmFei2K+3Py+AgLY83+YkUWdy2zcTSCtpRw
Wo+QpyPShLn13XWijFT4DvvK64xywaiknF3TwLnm4svLJYI8pEfLynhmH9St2U11dbZQbFO76oap
zuUzyMKUiGQFjj1VfzT9X0MWkb/aVr8bALtXUjMYiyHgSx3eEblD9sm0v0zIq3R3g0sXTOt0y0Fg
QN9rZWJndodmQ/PzyZx3WjRyVSTMBtLZ7wiXncpI85gc7B3SXKujcHnuGgRPeNHYOGC/8ZAPK3yW
5I1ePIY5ImJvvV6Z97DXiRaeMrlVZEAC9kx2i0hjwqqH0B9H0ix/DJP7etVP7/3QUN+PUN+kfs9N
Jqfsp466KO1L9BRD25BLBHxsAPzVWsbpjTJb7Jdu5V07I/adzD30FNrKw7kOLM7KxPAF9RZZmyks
ap7kG/OnP5/mUN+B2AkogeUlk/JH7JacIPKazjKOhskFH57NKJANf+zXXFM1zVnAByQ8TquxGhKX
neT3MBOGiWoV4sIwcMyCmrKNanzSlqR35bqgYFuM/WWN0CBEfvT2/h6tos7H763VZbgT8riYCncy
dLV38e74feksrUKQfX6Ot3E/ViTVgF82pi9xiB3Jotu+udBJObPzS/6wcybgs4NMTVEQOombTDq0
vOqKNHJF4DXIdXvlQQhO3ePE0PSlpq3zU4RiFVChBd3NrbYJVMsnkmOvYwMFd4++TmP3+jZTdUJa
Clshm/P0S6jftZMP0xO5VASeLVizQtdbddw4g9FLPRAsdB+wealP0Eng7+jfYjmM4fyrFLNa9LoZ
80b838ND1ayfQGMagGDP/apyrfpEfa/6sd4nqkTU0iONIADUINqd/qOVw0SR+mzczLrQ8uLMKj1m
4lxsVGaWRgQzMRcDUk7Y73YL6SxQopYjSYJICLgF8TtT058fkL6mLM3v3AkPbWc6hckKQTOOwpFA
xB0EwHe3iP+7sH8Le03Ek+t5flodNUSJyAxLCrG6BNU9kq7pSDzNeh7uLOJA6PaizcOSYVzrrzG3
gDMQSUafiSvkAuOUIpst4yF020YxQ1R1Kozd8oPmN1nlt2hmHLnJo7lopz9s2WOe7ZspO1E/9+C5
o0QKcWiobok6gQ3EtKGME5PXwA6hVTOzY8v0dNiOQOVyPAr6byO32KTeMcvyzzjzJESTApa+7vRW
PTPBC9ZxrBeyXFH4Y1PxSHcJu0slztxHvEEW3fLvuEFeJmlOzx6cxbeGv4NzbDQhZN1iHlmi1+7R
JByWQf2xoLEpI5AtU8M3l57wiG7Lt1iAhPldU6nHNyrVpYcn7sVHhIFUGAd+tkMT2gyhDcLg8yzN
jNzz+/F+0Jq13kz4r/FPUeFraQCbG1hUvnC+GkjBp97G+ogeboF71ozmwfXbXHB2COJAbV7K8aGQ
kY1kGh4uu2w1W++ReRPhKvynRh9+y3R9Pk7v5+SVGGdlnjFrXhx+9y32X+7cD2H9asKUdI8uQ7a6
0jCiCSgrTREt/5BX0W+acyCc11uCPgJ2uf2b8e01fmTsblb6k+jLSPUzAZOjKNOTfDU7cPgyQ0Va
tpDUiTQf18nGTxxoUUUNKnB81g94j5FSWg5hr1qtSCw01oxhPt3ou+uZHAgJbzjKbAlxrVbU8RP5
JVk73TBxytehkp2+wmTFIFpU3kbxXVm5OEIfhNOPnb568DYZjGFWTIsJEMqd8yxpsmFX6wZU0SI6
fq0aBs6YHYixXihVDLP9v1D7QGbqqOld9ZJGNCpFdxCbxZco46rrW6WOB8t2r4sQycSUePZxD8oD
r3I63WVYvAx4mP8/6rfcwh0k2iJ62jJ+Eb1YrHJLbBSggUhwsP97EWjAWSVbYGcLqMk/0zznB8GE
0fnOByKBguEZ6bh3oVslWzVcUiGlUzcxqItbRBO84lE1W8aQCyZvswn6kakgrhfrkXRcWtcDTBrG
64ovds7jWd0h8ExlrXHv3EFh9CWjWVP5ZdPI25HdHXR2eW4bZ2rjnOiHKbSahvDBJ2+WP/Z+VqAq
TNN1KLFB+5+QGQ7lBbOchzFvj3wGyby50UpixzTV80fx8DdQP63EPGkwdIvmaOanT3vAHQZ8emQ5
vXImTH/emP7u2Eqh4QgHXrf4suPErmym3Gg8OmmircZlXIt1sZ9AxPG2h5S9Q1vCuquoqD3iImhT
CPpABKvcCEz0OG2u2Exu/IxmzQvliVWRJzVFWhmmtdObBeMugdG7iDc4LOq+ubd77o3mSFFhdkvX
Zq7TpVqPDUbgLMZnmocW4BD7mfrPhMHZfkGPQIMXfsUJDGYyEZqyIpihk9cro8WO2pm2DzAfWPM9
8GQTY+36JGeRTHJACRSpdpz5LtKHOKuD9BrHftzSTpKnznl/Xr31q9qxawJmNJ9BTyKSaKeTdHon
FV5x2fFPPchDYotFQ8uUeAOw+eEVAoeYAF1614UV4BQy2v31Q0z0bEWJmzaK139Q3ZljRScKknaG
YBL5dtYWLGCr9gwctFI1U9oMCYuUL0zDxNlw/ggtVzCZPUZEXR1WtCIopAK1kPgiePisUDXP1h2l
ahe3yK0zwZ/g1DyMH438orz9Isu39zJQMKQ/DoV25g/daE2hKxp6VGzifJWfATnZxBdcPNKDvNlo
xlr0803YWx4dnf1kOtD3O98He0Sk6T7fS24XZtJz9Wd6d8YpNibIy/c9GRGSRiAk5AyPssuxA4EW
57jLiUemuLhv8fG28GwsBL7uCBvlAljg7wHOiP5Y4/8gmJIdRMkzXy8aInwRZ8V2LcqbIuX2D+2c
EHnsEEqz3ZhjaCqBu18gdmW1wp8U/vjK0Bfs+KRZ5np3FpwTkQt9/gaGt9nwlF5wqQJw4EddlDoG
FVRsNhQfXdjYbNZv5/7sfjxmzG5cx+0HjGZvbHXe7heIWGBdP0SCiObdYfffkdHNb6uoFIh8sQtr
J7BlSw52+M7QmBK5ij7ExBLvcCihs5+b7Jctd0mKort2nd+Qgb15cgDMYx8SnoHJAPdCPamusM/B
U40UxbpibZWP3oevlNLGiArRXAQLiO6mZwidG/wIV6so7wRtHPncx81DRcxRrbu0j33ICUpstH/O
ut4qkWoHi6Pyo3JmdJVyTnNaeg9trtORuiOsf2eWJK9Ykd4xzoaJi39bLY68z5BgiShE998JiJQA
H+Q7902jKMJwAazF/HKDiG9lNgyTJkvMlfe9mmf6UZf0EKac99Z0I900x7gVVbrQeqz4Z34+WB/v
cskWfHtkt5cdNhz0FvDbJ7i443Lpq1aX820M7AHaYYlzEMhoziYF6nWY2jSmNpy8TyCJet5mt/oV
6Js7JLE/2jWn64Iu3YxDaZFMH9r4Z7Om7/R3sAYV1aavKdoiS0vrMmYHi8Qq5siyiSE9gEa0axdd
omvlTq8KnaBJlcHVOoH8xnKyU+XtcJkqDA8Ex3mTmo2V5p6QGFEqP4RgONSK2lGY3XsTR2j9Vg0O
2TU3qmw7bt3sSmRO/eyXAChNJi72DJIMb4D54/RG284/M7r9Dq26+NQtEmoCvC7MWCR54pUzcMwb
DEJLD79hfn0V5mBHB4i8SKb5gL7eCIgMR+/G6KytlWMzii/7zmXQKcsAUHIEDNskM1AcZgb9frj9
5Dn5N+gmsHg9EZ0H8Lx7c/q92B8QvHiN+1aK1oCcskgAHloww5O3CqsbRmgR670VnCpDki5CyT0E
qFteiwbpCDEi9MBHRrWvPmP1/+xhtMAYl5Tv8F0Hx/i2nZzFhh0ZGg3E2zaf0FI+bg9NC/1OfB/k
8QK62KiAQVhN65IeNeyR6NwNjZCHnprwiqL5NlSlUKB4Lc4rezkO8jQX9eIrtfBOnkJnuypFdgIV
Cg/+O58CGU9sopO2DJAiYMJCnPawUkfmSTOGD3MwftBNtzoH0UAq6j70Y9ONUysdBJmBShlSTCyl
JrxJdJtZVlUvvN2qa8EUISACG/U9QICiOB6IvgQubYqk3EezYBG33bjbwBoznVgORzahhHcL9Auk
koVg+dJLs1SdxjLn7E+Pt59fI1kLfNz6wu8yFpDW74/KzgNAfNbhkAcw1ciq3XugjxKx7I+F4RfF
b+01EvrghdpXLCs2mMe/p1ZvZxfkKrx90jgQagY3bKf2qhetyOEhu0ewVnS84Zi6jFBN9/GdwDKO
VN1umHD1QeeVg3OebzPD6pfTmDfXTT4rovFVF1SeGiDCAZ68jVdYmSDdyBB1ZD144bxQp+kmg5AA
jrTHsgIZ/UDtJjDl8/4Wi7u8taLcfJanKxJDDqr/kMbdgTvc4+aqx8yihqjbNImt6O2HI56BbOTS
PcvkyFKYz2zq3EcXzboIoM6UIx2pj2hAM+XMf3M9NKlSie/yN8JMttsWsm9gpsjmDOd6SJTtoRha
nxHfk+85USqWLVmSTJ7grO5lv/CxSdj8N6NvT5QQXApfLyiQzGWUtSaXmZd/XQ0A0hSzl+087or9
CMIxqz+l+xwdBlZKSnLknJa2W5J3eHhd4LhHQHj/mrL9xu4+EM5EQ+fdHoxsdf7n7k9eXA/dL4D/
dQ05f7uPBI6qzRjFek2/3F7HN9AOkH8PSKdXISl1ZTDHWnsWO6st3hEpE7UcPnA32e/Aq8+8Aly1
FGzUvTzmp4DSt/ejiAwjlS9pp4e8R1kF5tC4JBWWkTt8sraFbIa53ux8g0IV4W3P6qF5UMliVZ4t
8PLJHxp6yI4+IBcqcLcO7kD2HwuBGf/Gbfa3VZqTsBhz3HjtN/12INt7hed62AfZjNQiq/9eR3+C
ebvKGWNCEbrh5ZAOi0GwiiCrXw7wTPZsD8Dz9MdqQrX61KX2VJyCR9fw3tLeVZsdlec6Oe79IhNd
9ruCmfldBvGQ2oDNjUuHndR22amx/kGsJw/0qwfEIC2eQqrAlPHiMMK1AwC/WIK1TazINKHIHj4e
506UfL0SlA82z5EFNqMHflLvmEeuj9/Q9efKkW+T0X0pOukDMVFJpgOMx2lHtW4RAgB0k2znML5w
7D0PDinngXaRGqzTyRGUUZ0foQWjVmixsf1tQ/Xf21C4CzD1BrOGxkqMsqN5TSKLZRScW/5Gf5KQ
G5IIuwrmoQPEzRKrYg2peuLBJdflkHi5ZTdt5ReoBboGDQXvrDWTlmwShjF+ch0gOCqWcGRbmwg8
1GbFyWMElGl/B5cj7XB6OLfY7v3HN6FLHT30I+ye7zezz6uYoCmQOS6p7bySE1HW+jikx58GUfCY
3U5skm1k5FSzXZSaEyc2VcTNKYbzyd6+R0J5DN+zb9rT/NtEkYNHMtRtfemDl3r/ykkSTYB0w8+r
yfXm03R2PK2vo66ObQo9kSJLczhruOmuft+/h4xst8xvmgnfdEa/tTKy0qB9Os97iPBPZuxDfJ7e
53k1/Cp5zcaMydnYWMoHs4mWEryi2HoKCFPMQV9/M7gpaneK0pLq8drbo0CD9WhxzLyGjdbCwoMi
IEWc3vaqNXjZajyaEe4uScgE5CyHM9hQvMixXft8U0y+BaXQ10WR5BP9fAhPdeqxN+Glns+kU/Xk
M5CBDuCsj8OEUr5BDLblcNXqypY4Ln+1vr4PeWExvMiqP6aPCoc4SpprYmkvY/tkX7uGsIudau4V
ZlnaBtVbm1Ac6ajNzrMN8mhXjOrdzEIcZoJa9BTaKJbjntc7NksMgJla4MFCdGiHK8XmMQBwuE02
oH6hkCSMGmVGAZwBJVz86eqxFn3gAEqVvZlqVcUcqlPIlrpwkc2TmA1YKxTLaHbXjNWZ/+5x1X6o
saqVoV6MhofNc+IBS1UvH+sM8fXSJJ/31je2ov0GAyiNT2UuVPnGTLa6daYoU9KIxBvGdrQV7rrq
xgQG+UMH2nPEdkhZ5+/V9QqkxB1iNb2Q3HxGqpRFn+elkcDDWTu9pGoI/cLsJwm6b+0ns8YiKXJg
ToM7qVaIxIE89HU3XeqmRVZc+vp4OOA0rioS/R6dSmOHbPXjruSlJaVicYrpUpi3wgrUIwHDaMjF
58bnGcfGG4ysm8n39D9gtSS0MJ2e4vPPZFAb1an3uGJ77TWooOPuu4TzuLxF64KpDJZJKv0bT2wG
IxR4zaGN6r1ImGs4lJrFjPVKfLUCGhJFOIA+8ZtIPfNmF8WSrlfj5l0AC7MgvlGbL+YDh7yu1gPG
eIni4iUy2i4rc+9vafh4lr+n+UqLKOVqofKybH07vRiNL/aRJBEOT9ZmYXS/iZwWciR0/ULYxyMh
hex0gbM/jLpnFvoYuGlcm2QFFp/1CVFHqHVwSjpzcv4dCOcJ9O0BhJhF4Q7kLPNIHKwJirM3heKY
6hAbk56OjSyX6T/uAdL/Qb1EuXlzdWMcVAARO9qPUf43wbsnQ0HRJTJY9sO5x6FZpucGllWR3Hs4
RDS4IFxO1tqliUrP/8WrMCOcmbieBHHF5SJdm46ATtgA6PqjwHVckpyz7DMP0xQ0rPJVrjOFy4gV
HrsicaCtWlafr43u0LSYsWOtIqwWzhO9/Xc0m3ycZGA0thzvXRrkFKsUoLwH3eJymuYm99FG6FBh
FMevgj1rItvH9ODpckwmloRwhLjoT0k68+iH6rZvkxptKpNL3/Ou6FfMhaoZYreme67THEOmmkOV
VIjsDcPs0JxNaCGFiusmxEucH/7HECGfp/+g+NsrydizVQKBju31IPlu7FmGE5C7WZXp9zAoXodB
ZeaYTY7Dl00om6Fado/r+3ToM1BCwVhfBoKRkd7NhRHkuqGGFEES21hxUPP1V9LYLXDlv5umyG+Q
VibNQZJ+vNMEOTwZLoRg7mGTM81KTXZuE12KxrkNNeklYqh0dfEhldWRZbX3AlJXOJIs8nEZh5kC
Eu/oLZIOemvEIs+6dCHbAJ+6jq09QD1QQBV/b+Ss4zZbBrBo+aEmTv6kcOyKt8HcMWVsMfdDa8Xm
d6Tnd1LCyFPkYRdqxIMDRmhkbaOPcfS3w6AVXrHrVos9g0PEaCUnHX3L832LseHg0rhU/XGAsJzw
Rfoujw7WEqfinDxO27fJ3WNKOBiCdN3pJLpVcqzoHHD+4+CTfJnycQsHdEJd90tOiw0TMxL4JrK3
/pdwUP+53qfbm5SQPiKRNn2d89yh0aFe2WwFZte7hqtjMjipWsGeJ1UiFr4jdY91Z2XrMw5xjlCa
0Cd6QMCLpj8Sfz27cPrpL0fh0Ii3FMYlHhEA6wt7Aw3bidIoAXOR9WpBcnn1KTqGbP3GldyQZCJT
MpOQdNYkfTBYWq5VgioPxp0dnbn72p7QznSZmljARSzjFmThmYF3xcJubYgXuWKOByscODpDc2zE
CCP/GHDHuT1YUwVX7W9NzZmMllRVW0LPtoV47R27bDozEtcpMoGEuYu+ZIOhfW54aCWhEZqrt6y9
mluq1DMs5350g6MLv224zf6+V+nn7eWSkBm/G2XcrHzmU7Og8cKbheHDZKU3Jnrqh1qbT/iioMpi
fSZ8yoFxDDytAzIihM9vHHSm6ey8nlen4y+mv1QtfK+OkoSC4RJkH4rG/MP+ZteCvsXH5qFlpfEA
PSpCchUL/aMbCwA89TC/cbyQOqU4jze0DRBixQFjtQyiKOsNQQv203n42ZgU5xBRARLUMjSrUJHu
qNGwe3PKdygr3OLfLYHOOXYDqOg5u0AX0lTvV3HoUhGduxy8kruwVbEi61gj6Y+WvqCjUBsJfe1D
REJO0MWQjSH37rUMXTu0qAV+RIQqGPjv7TjnffqFS0Vl2Z/Qntq7vxPTHO5BjlauUOYRaLDnlbGG
FJ0pPkM2JClnrEutjtEWYf1bFLLaKsdsHn5mTxkuJuE/MGwPd6LN80RXBBphR0bPlvl9aYk+7483
/ba5sp6zEsKh9QLlm0VXS7mnSIRiD8F28EpxbSRyZUvCP0qJBO/tzUjSHuTSnySUdI3JM+mdzTf8
lXqtv/6Qa5g5cAp5yDKx76ok3aOzITj6GR5y4t2OSw9ACc9Zy+ASQ1/5RZJLPLMphQhtTAaPAgij
Dw5p+y0jXBOCG9aj+1vuJLuqliWNd0DtkxHj/yNaDDrllBJa+VoF3FLJw1oEYjEVm5+mx+a7vZIM
R3E2RLrOlJDndW2ZdjQ0NKSaBNSZsDefdsAZOah5ui8xFKvNQ53puYb8rs7g6If4dFWEAA2VgohU
PD2oP8QheTE9wuKngKN//9Xc0ir2SAOj90jGNOUUUuiay8nPQXf7KleX205XT66bHnAaKsCRX97g
K0A9BU4VGC/Q6Sj+Qruu0775iKMvjJTMupMiExhVTEaOr8EYNqtERnESPn2Pa07aZ/Q7RyFXZJZG
ZH/iD5t6x+RTNBpd6TniVmdjOgjMRuY5n67ISef8DpgrBcnQOM0YBesucTB9Et6kQcqBp1HJphgz
/I7ANRVJ+zLVpxRoRQFDjhWJsn4ghlsejXgsc0gGOr3fK1ocXMcgBSPyndYSRKf7X8JDNyIvOZgm
2zCt1eI71qvVfmelEupI7+TT0aC68kShEaDB4o9EU1Bu0p587ZfXqHZQT7QlFZ7et8+TeDtybUvw
25+TDL6X299URCKJAqCQLITQtj8pmwxHhph/fqrYBZDZnh9YBpTp1M6uZKarbTDbukSz4ANSHOeo
mLLrBUnAGc6dlGZ31T9tN3mpB2dtXKji+vfZwjulIro7W97WCkn7pG9vWcMcuKnH7LZXOa3M/Pwh
YaY2PHLlQYzy+RuuRaIb0egVQm5uD+dnIzBnKmN520GzNOZO/x94/dvTkYxl2HO+FtuzePGOtQg0
kyAOWdpvMFtlQ/WRUOgyqFB4TAwUlVDIiZbK0L9h8dAaGXGINP3II+3Zj/D2rhU1FHaI0OL3ful0
7vkpq7Xl7NPioZV/iWViQ13KCRMGzX5cgQt5hzHP8c2KZROkOIAHgT8I75UxkhiEwnsuBLHtibvp
/qjCaobfH5+GLcrJHDT5R/z5uvK3HisVTZMSo5jzkGVcr9pM5uLgLkuW8CBWEu3aE6H+hQukAP/p
v7Y5KXnrzDKzyzsf1ebMIKUEJdRqCtCUEmKmmrg8d83Pfy5htPwe+jYNnAS0zOB3nHqe7WMejivD
WRY9d38nzujM0DoOd+GvSBzBd2Nm7bWYtXW/b8opPqCN/xVxvibg4iV1aNea5YjDTxyEStc3v0Xr
tAx0ghwxbNdgIaibMifLJO/mPSst5y6DXdNMhNDUsg+3HvbrVG6wECf90JeY10r1EyxgRyYBiGsv
2OCYe3aOJw5WXQ71NWA+pAtzcTDIEBb9vm//ffjFUL4PFoeT9M0PkTs2j9XmuOevLgPMtdblBUmL
ZFPY8i4E0a3gNfGith+rONPUq4wcsNcY83ufWASwijs57PDZgO9P8dcFFJsAMz0gj3Ak136eoz5E
qz2iQCcO9r1kDZ7XeW6pw0060QlXxObQ4T7nbuvpfAdR/yigEReexv1qRN2tv8c7DYSrU0MyPiYD
m6nj4lMZBJ8IFXXKbMAJaiNs18QLqz4N8EKkXELgK3TnMMoUqmTqN3/HgWvp65Mkcu13fEXWv6Ol
NWgk/zfZANCDO3DHraS9oiVN2RiPDxjXaAxdCVtAu18eBSWrBQscozG+sFRb3Oqn1FMbPsmKF9z7
xuhpU5WSMW0n7UFaidGg27QW89QwTYdRr1AWu133Gg7DTt9h58Az+chKRvB3oO/+pUKNZTmtmmjy
Ig5sXsN7LPxh4wkwE8gG+qDNlBEPC2V1zXwPOc/sCN1/sa8MJHsYaBSH3c2KzxAt3KF4HdzHBlQF
zFO5AOT8r7xUGsIjKT4CtFJ2inJaKrm7+4aRrpfHNR1ur5wpOffsOo/WOdpApvoPSFxJ7B8g/ceZ
qrpbbTdsA1HqLG7zaqhI/TQs5XsSyYbU6hVHtLhlmJoJsqAjip+iBNEwFofJ5erMtVJm4xHHgpEC
JCFQvhWSTdy1BGDba1wy+md5g2Mc825Dxin+j4kPZ0Qmnp9VB8yGUgEP5+k9wyH01kb7bI2/PgJN
ExgDglKNn2kOQOns9q5VvgbayRhGCkmXR8otisJtBGx4dQlR9pc/sT8jSciorkkTtO8skvFI5tcE
sJcGvSTREBSnSsFgphpWcCcL1BQccI6XcAkRvKurHL0lKAiFEcZzx4/puo8+m0z/Fpp2qrp16ngU
E1Mj8xdDHiCCQDoIqo3F1BwR0b/z84KrY3WK3JabJZEXC6cmBw4aVd00dh2JxTEtjNJIaaMpHxPX
pQg0ht/H4zVB7VDI3oKu2KFDVCuF4qBWCmPuKhvqVizuq9oRFfuXnfl64s0PflqSqu7UjOxnXdGa
owhcoGva+ENftWw9C7TkGaNTEn4u5P58KpCtyO1IE20K7qsD7ZkB+fNO9e+ja5tIVuL3yKED/4KW
QfkdPawfXDr8+Qrgi8VznTTcnidNDvsnhyclvPs+AciOWPJOyOt9d0/mblGo6l96eA+Cea2zokkU
ZAIEsqffRknJBWEu9laFyjrltfesct7mGQD4FDJK+a2u+km6YpuWTuOhR8D72EFwTO5aQMlfCEXv
ztakvm8MJiQqYmLeFz5lzW1YWlYYiDvSodFVZw4OMgoSCuV6gGdqsTQtDrU6c6iSvLZfVpSriNxE
DhgniQJusSXl1JvGQnPLR5pj3gcvfszU2NzzRuwfrwws7gFNrum0MW0p+ZtwpSzHLxewexc2BMfn
4RhXPZT+KF8f+uhFBMrL0Il9U3WFCZPhtfdSG4QBiDOCOI5fc6Fs16OfGAZsRg4hDq28b24TJb39
WwmtVGh/BmeyZWY5T10h9/o7boNsMTr6vnonTk47yINX8xS1LzGQDa5Srxmnnrqqu+EdYnSGZKwJ
9wvSV8gIaRVaI15XWpiR1Q4bLyE+GEz10rqHvzzR0+jTn5nh1jXiaqQuHt/T2VtPPQahh7mhFVtP
r6+MzbDgNkOnlSBmxGRR4tAa3tlP0q8IGkmipWU7RnIHZOto9u2Z3yZvuNFz8f0a7bFcCs2vUZsU
oVITbXjn440jBcd3AOYtdGv4MfrnyBK4v4hsWZtmU7X1DxcWg7N7wpBoLBz//poTgeSZfhdMG0SH
o2nnIR8bGILbOCVaR9nEuxUIa7ApctHLD3qaU0a1ihgdLqsp9ll4G6SSCdsN9wwY5Wv3kxsgiolT
Mj1UT9nk8USPW2nanhiZPCzf3yT0ITG0Pru1AWl+bEc+8xihog56ZW2/LjCtcTkwAH+xRnHk7qlu
lCchW3tI9qwzQLLAnxPF7zaGem0l+DfByz1k4aP1zD6ZuyGkI12aE8lcOf1flh07ylyu6WReFhPU
Qhw9tsgSaLuGkahbo1VfQs23Wrqp9VmQBZckkYdQ3vbiChnAdaj68n/fGLejMf2XcKeFbz37uZKh
N329oT95S7j+W2Iy9+ATdRye+pv7kEegSEWVlOEyGg3GO5J4Cs1859UVnTXpdWvLIAxypTcCVeZ8
cH40H+K+Do5ex9MTA0Ol9BRyVWPaAa0Ck9u7qSKgLcUn+f0ixnexnFNeGVK2KWrVUA+6r9QQ5PUa
zluLZcPEQDDWKcbESlxAGXbC5oEsEhCm55CWeZTRgManHW3Ua58Jt+6v+Cx3kHfW/k9CRyt2ycGW
12lfLHXngj4sg03gRly3cbJveIJHntPpLgncaYhMOcTopoJhbCQ9qwghbqhzYQGKBBfCQaDCi15G
TEkYwYr4ab4Hw1pC5NBGk1t5r3spRQgmELjlsgrg0e23TTu2SQutSnh/Ko9O40hOVfji4lChjdhs
cdoN/YTne+xqQmh3EjL93mmDJUTiOaUmY9euGZ2rdLDeNyki/ub+SK+stMI3JRPEhakcjt7JuGCX
r8jSquF6WzDeh+5MpbJ+l3YdvLQuVO7xICeFaO2xN9LXd2JV5BgkiTH8Btc0X+HxgA0JwEq/KGe7
CIo9rboipX8QG4B2pgpoeHVrESrUPk5B9dqDOSPCQ95cNoTCpGvfNbFXvwHCjqFTk+GlByE+iHOe
GnQfyjOEiHFHhlsNS1UAjF2QtW3/yY5VKbtzD5Y94p+V0dtPKk2FeQdUabBEi92pdMHU8Q1Z7Eh7
gEtj3Rt3tcFNh2YTaIw6UgShKu9LXoCB4FOv2MpMrAj6J0OhEThko0XZ62N4g8UWXcflRfWPlVv2
rUGeUQqhjYm92aGoVfC8KmPTR9e8EukOKMFukoV0zv3m5uczC9vbW03nqkbiJ7DC2WdXQZpk30YX
0M432scpKKJqm1LYHfO0RbN2NotNh14iKrLUXJAt8Weiv0l3d2/ugsmq/dJp4xZfX6XR7drPXMMW
17Ci7jzdH6O+MVFZwKMptWpbddEigNNk+ddXKCS60oUAwf9Sg5vimwL49sM2UQIbqOU+/xcg5LPu
SKzJNLLrNpMmSzizVWoJlvL2cVo7lYl2w/RhgXrU32FNgLZytOr7mRnm8ZIMy5a4YHddZm0tcBzu
5tC0/J+Hw5uLebfM03Z4WvrUwpN5HvTBuUooF/y+W2KiTJwD0eo3Jmj+WP34gXdg1V0GowyffhD1
YsxnwJQiKVUNpsoDeCqrPwyHJEC94yR0qaeP32PR269ynWMSacSiMTaJmXT/vZOX/fZH/GWIuZ3u
VJuSLAijFJHH640bk+EoZ9a6mlh4QZojX4Z2B4kJHaosYgHaK3mAr9lKEiO3ZHrOciS7y5BvK2Ds
EqOUUmPMB74NTKN05n4G4IfUWKXqSYt3M5mDj9nWzJiy0aSjkuHvIp3Qkv49v6tarTXcROmyuQBM
4AAzGEnUSUtMVQDctBtGCUHJ/NnDkKUnlsHkJzyRtmMtlBwjOI0oVCa+g9vBMJb0jXBPjZoR+81p
U2jj0IlHgkGjjxZ8aZqX088DfgrUl4SGN/afQGtkAzMI/jXpKQnG8kcFGabAz8CWvVdkjH2mid4u
qs2qkXZZasDVE0yEviLsLXXW8gDHeUb1lf2iSu6qyrhMvCv7MPhxKgaZ9VruVan5PEwtscHnMfvb
0VGEKnrIU4Vt/Xlk1NTRhnN0lWphWAbB05S+oGTh6vyBQL4w9wgUa9NbHtXYREXZGJEQNIuvOL6G
CZ1L1OcpVzN7jKm3vuLfDHt8VSttBJBZ4wP4uZrNezYwY8bqucaOulYZx0N6rZmGP7AZv0dZaTiv
XsWq2wQzFVfxFloa0r2wYnHncAmYh6VEKbTApgjVsXhufvERfaPS2lBlGUGg+PuY7XlBWnm603oi
w/FXWyf8MytLgTNIZuA0N2nNvCAWngM4alnN8E7r8DZn0/UFmzUKcOdvH3Ho28SVkwLoZkFyK1jW
O0OdtQls69w6P1nDw/8Iu1sCOC53P1dKH9Gdfd6bFEgGvIkA14pt6o+6ej7NfXXPac2F1OmpvIZN
9cwQmiOGEPHJVuSB0tgcNL0MpNfjSXkC2NNOhrFaFlMmwtHeX9uxl0KNU3hFyNBnqRWYzvMKYWCo
x+7WSqofUx9hnvpZyME1vDXsxMG52sJgpnRgt0t9AhJRA0+guswlaZfBhQV3ISjG7pJVT+lwNPIX
/jU5crYrw/gdXlQAAliU/WO7FujbqQ4VaXwQXGBoAHsfB2TD/ZGjmnNySNwBx0708SNsKd6TBvmT
uBRHq+McGnkp0nTgUAmsjNqC6YxlwyutOrUHMU0w8T2PdX4BmiPZ2BYtN0u29Fc/wZ61ESfETotd
bnBlw4mw6pHYl6hIhCGCWrV1+Ms8m8gMQzJuA0p+3VtvHHZxPAVjPZO3yxbeqGbvDvhjrXwFpagQ
ZlMzS+zDLHfaRmkY7Yjj5BCwGs11uJoJy2LIWEhyKuY3zRvMoq1wKeGoKWysArhQkysEaztJuQq4
shxX3+JvsiNoLf5+gD5reqJslLrJlVs7aDHipcKrCNYvVZkLUq09pb+gQPSxg7fRuTV1eHk01ZpF
zd6F5KaYM8bTDW+qjjtetPBlEYFQPRs44MfsOP2u4XVOu8lWPdxY0tZCgPxvLXXp6eM+N5/Wz5+2
rAQGLq0W+u15caZLqPKM6YnVPdPMdcyUy4V/ARPE3llXuTI6G3qKtARI1Z74p2cXqD4251gjEE3k
CFS166xNI1S752ay9UzzIRuO/317skHla0K0jjZY6QGxeRzCnUzqQMlZ+rseYOO7AhWUXWnYcKtI
WGBx9JzWG+ZJOCiFlQ1Obkl7kQJDIkjJ1JZ0mmpzEiBVUfccEqtP1M/Q8KKbMRPeLqvJZeC9nclK
+/AzRIUI3OtVmFOMboyw2cjVZ0wZIWNKJAP08FeVumai+ne3FwLtmxgNBRF7boB5cu5/rDNn4hVx
t1o/gHfCCpR+d+IC8k9OOyxUqmB1Ef/LjivThdoMsqWLf1k7f14ddeoNL8+4LtFXUJ6sXzgPnNhM
39GcTYCxk5dEY8hSfTKHrCr2EHWdk8eTnl6vjVmGHQks4CSdTncTyTWhTDdS+FY2xqxLPY3ogSC0
gBJdPQkOqEmicDoMB+muDt//pUFRqBw9OTgxyBomBlF12dC9Hig7iJmArqVvB9Y8ToSM+0DSeUJl
GhvqL/Z3fOqtufKLGsTCiLJXZlSyH+NOqZF9II/OfTFr1FIL3A9B67mLgtialx5RXAiNl1QDOgE1
8oPuXt/h0AXCgXYjPwvnOe37cCMGjv3fs6M0puFgl/tIl6bwp/A1VytW1DvM44AEner5KdzZV7Dx
C1T05PBJ7V+i2LMJZC6od5v1eLiAmUuEbvH4w+DQ3ewo33GB7hXEVzYebIC08R0N4urHAa+sTCU/
69wRbNEMT1FC46Uk212xMs6NCDXWjAv6fI/vi7JCzhNQggI0uj3zX0NKcsbOeFPB4wWjaG1hNbSo
n9dXTdXwCUnLc7NHz19PRf6ebcTjRtJxAurHc3iOnFOeCg57hzYQIxiK0XeTr/23Ikq5tw4vt+b0
q5YLaIPrTpQYHx8fE17cd47zbxlWty/gmd8j465Pt+3TRPYyHhDgiq65d5Dwz2zi9ByJFYDcxFoX
k5tSVxohAyrmfQsS3OZhgMNrAXyoAyJX4q4lMG5LTNE+DEhrzFyzKzumCoXb3H9Bqipi/nOoATz3
WGP+G/WKbPhuSckHorlKTtxydKJd3bd/018zSt276BUf97a8viLKwRAJVmrXfEh/lENjn+wBiBa2
AxxdrarB105J9H8q4Kzqj+ihDUeDiCqX+qEJ/c536pIZprefp1Xr7QlUiaD8P3N0i62nzNiWLJAp
Wafui6bA8HyvTrS90kpwHvPC2/tgIDGV595U42tAXHKULLa1Of9Ps16hjLxwAIeIOTQJQEL3pKW4
322KocXTDmzcigAFOOOCn+tt86I1wPuq2/J/S0wOTEjHmkZ3lGpppG/T672uWLQgDuR8lJ9ujQED
7/Ydbni/jZASm/qgnhK9lN7ZrtB3yRK5NQFDBMxscnD+f6lh7vo55vEPTESZTUGTokpaloyCYSy5
8Yk52wmU+Bp3VI+4vOTFo0ML5f4DUfebrpVe9jMgMjZEq32U223rBO7fxwltqlQrAGB7AbZJLJBJ
xP8f09UGEriM6oM4wtSpZT3AvbngTPILnNj4Io8AwG0fie6l3DVetBHj5OW3ndENv20bnI7oRgsC
9XxhFDegD783vl7HiX6IkmmPaR5X1c3htXyl/HEfu7RxiaxzIEPa4PLJrufvR+EoeyZ7oBJnrBA1
OheYQdnlgSSkauKlAddw+dyYfm79+P94wOaw/f7IkKuUdX9yLkKNYHBGW3bjTKCba3YJGGmeYbGI
ZIwpaAbc9Qe8oXAUyzb4kyqGUwwsg/lQEPZw345J22q5vTlBVRW3GTNs40p9NivMp10a3+bFNLLd
kCkNervfuuUA3Ra+hYZW9xWZNIqCFtA01Ey5K5OR+leFUjvwCCUSU56TRPKUDk29NccJHlHxuSRt
7f52JNIc9cqqF/36bZkGCE4IExsndbVkwcxJocsYTwWLHqxb6r3RA+7zQhZx/uU3+lxPoKGFOpys
ejDOn63CDgk8bFWdA03V3h3cOgnZwqrttlB90re2yuBcFiJ62Q1RPNz9E3Ri5hrkZIHGOK0Zbe7w
xm2+Odn/oQ9dPJRADjtYAtnvAqHUpPo3qnuR0Z3LsQcoLWbunBWFaaO3k1otzmkQWeF4mkYDVtb0
vLX23NdFgyB5KNOLcvL/MqGEQNZGMEngtkqOiXWv9X+2OmH52Rk8SYD3oM9HdwJZRjzoeC+0BqmY
LO7y91qz1g7rmA3K74lRkTuQPibuYShcL2z2Qm3VttC8fHcfFjKc3vTPe4fvzHl+NW6yY6EKAXpY
jWGRnmjGlGgjxrA8FrHdpI8ovNuGaqHSLtRGYa4Yg0Lp3HrSvsaY6edsdavtKldr2it4czrK3mb0
UlHdDasc+roTivkCZKq11ioOHXtfcAUaobGNAH1pB5vkhDt5R0vUifeA+5n2OksfkyVXSehLemEa
ROKcaxl409PCNyishreidOsC6Ras5Tp4elLTT2fyOdwsqyZgmy7FihXiEA7QrCSRrELWfnLTILCk
+3agL2Y85Q6rB3gx4LcONLC4FrNf6NpjVM9Qewb1U445cpHZsWErJLJ6urjAfrG/CCqECZoACdxr
pUwEwUUECH3ltMjnL+3hmCqCGgM2Ee4twdpOyUsDkCxTL2IQpiXM96PLfN2qSgx40urzAyNFSy9C
Dppqca8qz22iCPTAULr72c/pdPsM6RCQbp4XwA4bUSHQ7Z14bDh/VWLqZFWBPw9KaYhqZyEABmEa
dEt8q58H4uFIpkNIXcyDLClvNh5waZRhz8EFIkj+bTb9rV0kUM6C9lU8syBSfFCW1wrsPZ0t5srt
Mv4YWBB8LohTf9Axc6EMyOiCfrnavTfkcQUWNr4jtOBI0Rhti4snz23utojmfsPeYaVr/A7n/rjl
6sBykFgK3d4wmq9UfspWUJjdKLqGmo9C3ejM3VgLcTfsOMzfhF2TNPofq6wTB81r4UnWMyMJtI8+
//UHAOvaAneQEotHhliwbxD0wpghH3uZjLq5zLHL7KvsdS1B7aOMbQJzyKsgHEyNzccFpRUms5Q6
15NYWe55h01iug+RcC8d9OgqZ3bIXDNGLsIzvRyW3eUOmgRiAelbA6F2JXf/AI1lKFkqd2CiG6Ov
OQ4hIWji2k/vBK6vwW98uBJDRzizrt+MOooKz09snvh60barpytcPTXey8qy2BcepqcdU50GF3uX
W5t94mb4lCahb1nUcRGvNzAOrq8HA/bHPeRuIvcMQ4sesCLLunYuhsDvRosu2KWNOEbTECE6lDz2
ckv7fY5YT/TOcQw5d4VtBAiDLXNjIpNXSLV6VYK0besRLo5+ohOEu1gn50uFjvDqY7+YFyLa0gby
3GnnSCwhqNvIxmDRKV8qmiBYdF4jbyzU/rYq3cWUx1Yt0Rs3MdUmy7qCJ3V/2EbV9FnqxA8ZoNgK
oOvKF2YQk59A9f5VKr7irLFA4Riz5B1kUl/4AdiYJhuqKA+YjoE0Dq3ak9jTB2/+yD/XUqj5zIgI
z5EQLkiZvQIl/pz4Un84D3Zk7gJuG+Cmppz6ZlAsUIAIAc0RCV7C4M42RZKr5xLq9joWxjGrV85L
Wz/A8QUePnOgYmagDVvpUt3uhJ2/GICi4DykoJSBrQJKH5zB9KBB7fcj/NOh2NOflgG5GUgxgf7B
NvFNd/X8kxff8roAW/iY+xKw52+emQs6pytRTOBWqiDy84z3QgGc+voBBhCMbY5SKprbR6SrP5MY
LcaBzVJlDVLegoZkgmi8C4PU3R08MJXZC/1rkZZeG3/3phpQ3Q9XsKGYepV2sAF7dWUkNT0RGIQd
ZgFeNS1UwbJu2RlAzSab2lr47lydGCepPkrtexpAbUSXI9kPqW0vorbP/3PdIsRj7OnUUawNlSGD
CcsID/3i58B0gHJwmDdeICz8SvvAUEk6S0taW1jSU7hmkW5g32WpVW+wmmNqb10PRkeWXRQfEDeu
LtZvHwDLH5I/1YcpNw/jzgltmlBbcFiea3dsSFJLbHSaauc9VtER1ePP5Ha2yT4B/WSuJ0HC4qJt
xtoqCSfrX0TJJMxe+hr653T8bsHnEEx0b5+3RehHlgD6nOAOMHi0EnlngiUB8HoDy3NdPYOVKsf5
4syBvpiA4DLLUls0hOf4akgnYiq+vX0zh/dKDt4ggcfaGMsmmRMvBzdfVnokVniUlsh/8v+G8tQo
lIZ6wOUansvCCpztIAS2+O4c+vNlKdLtpnKKH8AVEXRxUWeE/huCwkryDs6XUcTd21el6axXmw1j
u+KoVDB9+K9Lb8B+vpVXlfrHOYUE7ZdJ6mkV0+Kb8ZgQqfeoTnwySSBFShWBcaoyBrgXfESjoLNP
Et7szWhMJAzGp28vclea92vzIIX/FJj7OU/3u8YTEsFWqqx5g/QnAcB/TDE0Ye3pb7IWeaCNE8Ef
y2rjuOcvZ2LuYtR9BfUcA3swrbScqqqDf8jrldQqWP1Dp1DxEMrBJgXdLwsYSzVNdR3M7FYfWQDS
FKGwB1L3nJriG0E+AOfb94e7BqttZgo3YRQYT1zAWTwqMpGhwWryo7rcOcHap2Na/P6qUo2aJSSd
FnOC0cPUZ4/fKmCk7u6+Ojwz3TcMuTYZX3C28jf2MksOnwldz3A1sKaJEC1ILJRWMjRKdoPcZXVx
Q4naeSdOHEdB5RCPwhJutnl+liMPsAz9gab/b8GpxmnPeJA2OZBbQAwTyTc96fJ+89DITk9hofGZ
qvAXSDWo1uRCKsa+CSoHK4/kUoC0effdeojxgAmUGlE13dfu1UI3PI978v5JThwx/QGw79obWT9r
GyOytFHVDVKaLz3I8yRj0yjjn/JargeWDPCfuhbNrKKMxc49cQ1ry/FAQjzzPycXwpfDjEqBzqkw
L7U86N+U3azeu3XR6NaauQscElYt5crFitG7wWLQJav8U/O7HarjTICWbvUt5JLrjGtse3yQTAWf
ExlEe+i8ZcFK+3LlJU641gQM9Yj41lrcUlfTnEccTCqZIGxEY/9gWbgIbpVyyaHd9LsJXeDnxjEl
CMiUFaxzRezD31Nxe4EZj46BWNlBqJc1L/vIeHKL2LHNZFTq+U2M8RYUvELH1iFt+Oh3uraBb6Pz
nWCg2yTIVBAKYXLNoTRw9DaVOFqaob40MxwbzwwlQD57+UFauJ4qa7EYdrAEc8Jm9Bw97rnkqXqq
csy1RDf2uXlsuU5PfC6SovTsSNzshOdk89aYh7NNC6JqWkWdQrckhqF00BPxyEW4j7izFkXm8KXE
PZgSD8zlaHxTmja4JbQJ6Iom2jxltqRQ7c3AoHkECsn6o4m1ci5ID4ywVKEblE4NOFLL2zg3+squ
/RTRJjWSFY9qx5C4KLi31pxQNEk0OzaiAF8eTeDethuC3RhGecuohlF4Sfuou/ngxFS1Jy+VDiVv
Uk+ZKeERVkyesMQg6njTqbgNkj9iHknpvRL68TBYCWIXJA5geUinPI6c2tz1dvjMicDTpm77dyfw
UnJsZ6yIDh/kKR0gwF7CEaQwbzTL8GZZg3buInx2EvG2ln0gI8srkEuLuKRwFbUhTo1QupJAZwzE
xt8JFXff/M130+ZAAex2xvQCh7A5HC9m+0NcSdV/uydZUKv24N3JljIdP1L3kyvsAQtIJRwp3e4b
WE8OGFl1om7tIXD3x1MuqnFyBHj3FBIHMTLEPh2e882pC3PRikbDnivIwTan4VTAkRpYOZm/0TuH
JGUR/Lj3AdsyXXEH72f0oWAnv/U2khO2445SrS0JOEeyBFwLYSVl4zS0h/lCT0T+8Xn3DSgjqBcT
tp+38EwwgHFycFMYMN7j/v0flcc2LbHkNdILr3xfS++d1HZoZFQn4CROoc3HyaQM+cRk2IowVqt3
y/KRy8QthgN6T2v6tUP4lxhTLSygQXGojUW6auENPX0bh0VYEdTfYrH3aSuosf+BXP7QZDixGRST
xWG0FerKHJjCOg4HKsBRgO2mUdMX74JMyVRv5DBEmd85cW9iMYvQ31HyMcJrGEXXWHkJT0APGPJ/
t74TJYuloMP1W5aq6maY55Ejx/Ye9GcGT0kF5sjsNgQQQAIfHQOA09/lb3HTybIFQPJMp8iHdvIV
H1WYfhlZi5mDw+ezbEf02SSUeoA5aR1osEvcJox/a67qVlk1Mg9/4JXUG3g6uhAvXh+HrAJHZ3gk
Rqncpe6DIjRyAgrlFaiImKx1iAL8wCPekPW97SiWL3aBLwMPPdBe7WX3h1MTXGG6oJOiM7Fcpoxv
WXKvUIanRNLIIPlp8u2kTzbh9WQwCGUm7QC2Y+xzmNQ0FEVg42wWkcNSLjwYv2bQx++LJTsl8w47
DqverEmd2NlHNxNuWJnPCmjHGP3MBVxLWJCq+l8LcCcgpC3zHnpg+wperyaoODs4meYzme0Gxxib
D+NTU0Ep1CuuIULxjtM0ANiv3dNMNLwcg8l6UhjhuIPT0t7zoUDIPMroVQ8QhW7JAwhC2bG9oXwx
Kf/R3ysha5mTzvjYbynI3pAhqVA07BasPa1M/y8GElcGnYObXQiIND9wD4eDsqp6uKY6QpIjCIoe
u0dwnq/7x/qrjPtUFsKB3qPeSO3iFoi3HiR1M5W6bhSqX5FU5qmff5N60DPtt4HhiQyoz9f04/1A
LxnUjUnfR2DwWu7Kkn+YFI1+i9v4CzbAIjQQTw4omGRvM9jNFYD07/hZ/yax+reqSADFjEWb4RlV
CAP8l1gOKMq76n1A1KtLBZ+oauvv+OCfc8uNjOG1r8Z3Ri9weUpmdmbn3wks81SoiId5qYjvO/g9
iZ2GiQKqxyA8sBf1SwBuUlOS1ouxOP7kYYOy6aLdC9g160/zMG4f3ZYeiw83B3K5rVvJuWBzzL7j
+PKDOW2FQZz0C3Uk2jq/3DJi6awsg+OzTLX/2EsJVe7qxQUZ3OyFvGCud2We2DDAzf/oBzQf3omz
N2Dva+cUbWVXB9XuCuMbesy/51eK09lHcYVe4Nu24BaGZQxKwQUkn4kRh6rU2kNGkVaN6M132nsX
gTX4S/vTEZccqZ0q4cBO9Yt8VAIwmTmovB2FOc7jvTwQDZHiu38j9oSTpMDZ3nN21+6yVut5mtDZ
JgmKtV9jZESh/GwIZC+CbkdvOmrAmcp3A/Jyp7hNh+UvOT8rkG7VzOrU/Hw+Q0XYJSv3vyuvTWqQ
S6XdbhjK+lCSaaj82Pw2HDI2dtEVamvRLebxXF1ir3Z41T9O0chmanK5aum26yRJqdpZIqs785EV
nhpOAslOPZtgyfCYPwDRPvD8flRfMPuxq9+HqKeVYhjan5wIa0rLHLLNNhAE8kfl3MvJOTsEkSqC
V/As0Df1krWFPve8dHLL4+08F4IWtr3HeD7yA6+Oxk2eUSKlF+bxPnWzKlKv8Blv4AXjTu4fi5MX
ocnuQwCoVQb7SxhaCE9FDhiGI5Zg/eyhgjxDc/IjEEXSLI54BZDC5gCt/VKWBCxagiXG9zdWdM8h
TrwYft7q25D0gYF8KGBHpUDzIOpLKGkr1hMO8VdoOHQFe72deIZjMMgbV0/KJ+AheP9py6gN50lL
OjrjQKtZR+bVMmCCdwt6QBN3MMU0BNe7lEkS5GluEF2hSRoyFwQZfBQ+tYUB9kIeVZ7PJqIYgdU9
Z1WKKi7jSAgNNC91F0dn5p4/7ZHQUbo2To8WB8XSxF2GLUJ8KYuYtPEReITJO/oNyX9WaeqZGOXF
+a16dIgHsLPJx8DA3lhvxMaNFcNuua8yFfyXgEN6a+Qf9/QhV8aMyPkdCZqx/HT6ZyAs7bLkRlrL
ghjBSXIpC0Gea1nIq8sYBNCcq+nmIi86Q9fZhnzU/L0Q0EyKBLcWlQ0Zmz7PdynJIlktUn1ihmfv
/1J0g/8ZPj9ISpDJ7bdMrnq9Ocmk7HkrKG/CoujfedwPXl+cQzDIQR787Dt0TnsC+VxpAmW5IuDe
LCLe7Fmu5wSGSMVh9KF2Eqd4ygKGY7+gXTjRntYuiNTT3Tx6t6uAw57Ec/ZJBGT6toxjJXkaJbKO
7WpDWP1gIA5Z6+bggWOxtOEgDHiz5qn/q2DiKB2Ir67E1SfWDQhyieEGsBzhvhfYIuyAvKeBnw/N
+AUkAngzET3CBhVVaaeLPVNO5aM0RRdFnBhyFQb/MWOfeEdLmmwohevRe7dp702cJiA+cT1M7BHd
MGRyQg1kXnx69N7PP/Y2zTUPPJdNz4X8B0lXpMdKQOasJ4voUSQLpSELsOI+2P1y0tbPUPogmzcs
LEHRkB+TyH9QYsNsdhGXUZYaqpYFW0oGGWgoNP4iDCaBVLka+v6my9/JqssNlOxWdb+hekSqXPA8
kkkVkw43Yr25MHHvpG8zjAoS3eKgKBr/hSRbFCpPHQrxAgtJxm5cha8mf2e6LjBCZKkjKzx/rBO4
59yEvZ8NQejH+zQihy7Q42MV3boNAh5r+PHbuL8Yi3uKGoke5Su+xFHvPEJoA0tyo4XT3jCAih6V
+GDPkTBSwmQyVo4XB44DMFaw5gPA08Z5xHJHV3UlBSFa1g7206V3SsKyqtuEsyFVwy7eN2ER9037
gW6pjTic4zo3Jq2CUT9Y2+YCOzhbCBc+rkHH7pjBbmXUXrs15t8f2Fod9rnre6rcKwrw+KLJdqkH
e8QRXA0JXU44OC0bqTMYcOGBP7R/RvZb4I++YeP962Xmcmu0GEk1If8vx1N2Q6XQxHPc4m+6ptK3
uCfdFdid6xKZkSOPXyu9NHlmMRPpwUbpO+lcJDuj9RLQNjITVoFPhgaSDVkf1ev8F63y6rvT3XPZ
zf+0BuAuVmt5vxxkPILq5oRSWia8PvLIo2c0E0ur2NjaI6bSSj2coF8GqF4cvjCTrWJhI5mPjc70
MCBRmJpu28QqpUMbzc6U6Hz7qbmHun+b5v2VzdHjsRB7FFXUmOe40NF6DkIJ1M5KkAwWpuskm2iT
9xf7erjilv0+qDOp8cFSNb3HzS3Z+medSbRo2SR0Oz2QLo4siixAj4oyyMG0NjQGm9FdA2ro+Ht+
XJQPSMwp1YXFP9ijcN4F8/wuZV1eAy+317lWUOHmFfcmWDH+Bvn4hz67QbQu5Bu19/zrNIzheZls
T7E+JQwV2cCnzAz1aaLwmbDSqrP6HiG6Q8cUAMNIc7mEA6picabRK+kM5PGUJ+KjZ64hct7Ed8j3
968Ytc/tgySY75qG4or7M2dwpeA4PwT9GPL72nIldAfRm80MpYhYjciZEkExc4Www2Dvj5jL1DGW
nExrfiKoEx/asmU0GNLm99U5cgTMUzDr+ss9rzIUlBHdrn0NjM/x5c/pKOQnOAXxmnbf/Muvfpok
almIatHBFsmWZq2wA5HvdeljscI6joeR+eYTLavCveiHZbCNoKb5JhCLa9WHqzmAuMcwvYMpnmOD
eo7f2EOfEpEPeNVMDzWuOYFAtVRHP2yer1H+6isac66K7QqzEnruM+J9ZJmVFpx1RKbfHVNivqq2
9OTZErmmP7N8WNc+2f3oPc0R7eui2zG5TVOKdC9k3tHh5g8a4pNe571RwmkuqZv3WceOv0LjtU5e
Kb1ZWpdN+O5C5xcQ5Je5U+zIFZ1m/6T3sOeQu1Qjm9b3f2ih6ge2PC4L5kKgly5RVTVNXye6Jxf+
wMi17U6sW2ncz0wyHNBNj15P6jABRM88Skdoey4TWYDyipgnG5XVxhsuETiMOFOYWzwuJHgU6Mis
JlHEU/tgAeCTK+TXvJMZ2HbRyYiO/u68r41kGQl/IzjMa/dYFQBeMcha0w/xGkkn2vFZMQq40pdb
EneNn/xhPrdgMMlE57x2gsP1W5wRtqcs/5hRqXuw2lwgo3QStimOqycrFGXN3x9rmIBDDWesV6cy
TaFMJvZ/UOMdk/xgC6OlNHCX2EtO1pf/SMwpqC6OONz3mCDZtr9qkmvCC0Vgt6Xs3VgZzALo2G9M
AwMMD1VO+/GEzs+JCGjb/PWWd7m3fFE0d8/goxHPIHnALrITYPesS2mW96eXRKcYUEsBVo1QLr5F
IN1BorDDtMnpUXu7E/c70bM+bA9bakuMddsCDz/GfKcD36PvUalbg4GbfGEDTtKBXmd2J65oTWJ/
8Ku0bR2EC+p7OqMePcDoLjwBmgaDTsQCq/uiaKX23YhbMrQtm7vdsEt9bwd2SJkK7HQmb3LT+MjN
dzRqxOZAfabHb6F7dgsXzE5TNuE50QmAv7Obs6YxOQuIpc6kOWF2YLyyz3pWPg9ZQfG+ggY6mYQ7
DJ6oWxu8xGqvEahiK8BIQoo9kp8vUaki33jYXycjbx2+3AaJT0u8oClxBvE/JqfyvnHplm5lxvKq
XE1Q0+PEceQa/7n7iWbwTGUZaI1l9a8sI1hUEKpxDlR6n/BDe/GNYhFwYS0oWuuBMxleB8ADsFnl
y4YSAimLfK5xYkKwvesAVWnv1JAANn/yzjZUIMfGx/5a32bJyd32JCHgjsUmpoTeoqwHcQym0daT
R5bW3KN0R6iXtPOvrZHNy7vcU0HL5Pk3xf+mzAJD8ZpjPQSkKPJfftXDT4wI/qQzQ5lb9QXiLMAu
n3ZM8RcZAR/EDD1trtCn1OXLLS1pyD6htGI0L7vsIccKQCdkiFsnd5BVnanxnxIrsDdpvAWLm/1P
qqhi6gN2QpxgAogbv3tP8kcT0KFCzR5TAxHFo8lGRd3CKNbjMW7qYxv5jK9Yid8hTJR5O+uMYyXU
h0CJI65cP9G7aQRowvQaiQsf999h1Pbt08MLQPRMONLZq9oQQPiEJmpMQLsFWfYdetLTXQGjivqk
i3X+Yu2GnYfAKKWWlRpPa5CaJrnAJKCjKsFgcfcA4EOQmm53WNZx4HkWq1vRZCmt1ABMuKkJs5Dk
rcCC4VLe1p/WY8E/gfLLjLY4+6VDR8MycuSZAqlul++2NsjgaP10u/sz21nb8YkV13YAigHNKthc
S0XHNiKwYxgxHnHBBCK1TgHGi0BnnCuEFAv+Uij0qoR4sUKLtNknP340HCDiwtcVv0HOejZcbayS
dLzgHRcpu9xbr6iu2K1zYJB0y5Lq0p9wlfwu7XrKpBQjCJS2gJZcPXHsZ3g0RHF3fMs3Yabi3kP8
feOuRTRoHMbAmdGcJjVFXeDWpLvP12qiuQNlnJIBdWeNlAob7zzhOemAbqYNRQt/0LrDvoolILO0
pD0MrPd3yTaCABk/ARkJwB7iBVSPWtmAb4JeQnh2WhTVaxpCpdWkPLKM0hitk6+Fwl3Js5fLN2OA
ctvqxl506420MLcxwUd6Vj+TvP70MmEshbjeZEBumvZrTnHT2zWQOSCQxWyr9KmSdDZppJfhbJyS
S4YotflHQDA3mEX8aLK8jkj1yOgTpVXrL0ohVfMJ6wzmPqu6iXNDVx+Ha9M2KJS2BgZH0iV8g7uV
cBv+9rwEPXJIlHrAh75GNM2jhAECusPSMu6GGvhIGHB7CjLyBy5k+RiBc1ocOXMaJbwgLZxZtetu
UxbORUygnzyTB/pVqMby+e/EpRieRO5zk8GEoUoBUSvRCFF3m/3gbJDMDrK376wAJPIR4GuPFdAQ
dn1rxzQOk4313Wfmmc8sNxVjOFRQyUV7G3S2iF4jjUD77UXKOsvzplpYuWjtP9ArPlQqhq1E7zMP
DHLWTC0l90Jtqrud6WJzxFb/yzR1tKxt+s9HKGt1AdVlv4nM8EP5a9yqJng9z8Wn+NmW+7AZ8VTV
Qdrt1gvlN4qJHPxCk/Axmkvgkis93c4wXKgFfQfQ5qCQmQDz0TCe0cLlsF21y8PFCDSWzhTnqvKG
4iMC+7q8p8Dsti+0dkTB/H/DdyDqH30k/NP/eiJEqhLf4hY9UcygBt3yXNYVhxvIJn9CVLe/9o4Z
6WdHupeClnviDXq5MGUzT2GdGZH2IXF6ye5dGToPSZqMC1GJZamV3gT/AzPqY5njfPRMZYhw7N3D
edatmeWVd7oWnJEyNxhgAkNDfhU0YwhgV3vHUWN8kVok47KqscC5BI75g2Ie6zHanSrq00xJ3RdV
Ne+aaWdTesQG/fN9pJ6jqMK5lcI0IVLRgwSldz1H2TITPh3GeQpGRNqkIQ9luhsBIrEUv7Pxi691
zSQq92DDDNc2VBXOpCFJH6gHQq1uGuoyP9UwrxzxZXawMHuFxlNQIdVTxWd8Vynx+XMMf/SSwITi
+k2/yF1ugsWe+f5g3cAc/IYqtyfZGcoTjznRNUFa1mRzaa7674nb4ERZgQlmQNViX0ziSYzrYpq+
6xBuAbmABt2Obq71gl5186uciv8bxkDNwCWERE/b1kZ5sKkHVQK+H3tQ6hk4hp0bRgURrocHvPtv
ajLTEI/gNeOqlRcmWfWwLGEhrSsud9dzRSIEzTbS89TMgOEdfY01JSD+98k3pUNF7DrsQ/rPfS2W
JILgEMQLUIY5/6hcewZb3BmSlQUnWFQGRqt5N4X/X5ZLEzjL96W3qNs8SGeIwp+1JoGXTownFjGl
oxDsOLMvuntyFB6WEn7s5avCFOJHo0+Iol7ra0X+bvbdiytZt7K1t4niUZU/Cd3EFYPaiNI7cnYC
tmi5Xm2FXwwd8Cevs6nM13UI5uJKWvwHaocb/eo2xszONNIumiaQPkXDFJeO8tFCpyJbW8BfB3e5
jKbfNjJ01vOrOVolFbz2RDipqlFEGXHOsS7NIX2sTm5i75BMDeu/gHGrl/R3tetawAqebiDoAf5g
bClNImJ9AUAvpevoPkIf2iv/waAnJHbnJTJH6TDKGuLyAb0pdSMjHGdDsKy76SpERvTbgouSpahu
FHxWMvWcuUZKs0CvRqyZkZZBMzojD6EvtJVqwxere8LAY3YvbJjxUdTXb+S4XOfYm+gl0LPwyl56
5sGmG5syIsVqy9iUSBAYAjKk2KFeagWKzwfLaUJn9F3Q7+MmkNlWUV7OQlQR28uAiywo/E9h2Dx4
4HiBLKl3dEO6retMR0jN3JlUsCbsc1GY7tYiNuoTuVxyZKiO7tYcxJ3jR0vzMfdCMXfVowJ2MB97
g8rtwTaZOolLplg6VxwOMbxQxjtFlqgqH72C7Ivp1uBylnw8CVBpv3NEA8lsGDTsD70rEUMDeDNT
gtnRydZEpe7o7tsUv/ooS8Z+lHIZL9HPkTpUHjq88mYEZVK/o9jvfQfU9ntt0ouWs+f6/8KQ9BCp
k4IOQjtxkVDvnu198Nb5U3CvwYo4YhwNGR5QKSJ3aQbaZ5sQB5zDy2SaMHmUIy1z7Z2lpjwSvCWf
L5Gz/8weddVQh0Li4WwgY9bbe7LT6CA0k7T01QKn6yu4xteuIVo00p2hUoMQkkK8Ja0TKxXLtahY
uqZw/hY4M6QcjhePyKhE166sMf9cAEyl+SvkwpXi+lt06J8Uj8UzN78VNX9gDtg/ePoEfBZKKLM3
DY9GP6m5QZzMZj1WwhqbamCLehoqdlqPH6WRAw7RN3Y/sY48Z0t6sfs7BnLaoHYndHhh2diTvCF7
KVtujrttHvty3PRMZQI2WR2hLhZ9Fxmw5gWjZzQdKZ1ZzzgnwWzI6gv2WqSmC/Ls27LPxL8pSNqU
tMpKWxOODZOVS57f+kROVF+5XQJwiIFhPr11aK7q5Wuowz/riPCcyrWZpYg8D55mHedp35ucCyma
bRsg+NpNWQoJC7egNAbboAKXqVUXUfiUaJmJxSJcQ/QppRPNDIAwsbW0sc+xQuS5W+52R6dAuIUE
XzbO04mlB/iRhaXfs9m3OvV0ls/URn78VDdI3OUxLzGMlaOViRu1/z7VNqscBEm9Za11zMRneuRa
WXI4OCWz5tMvpwdXyXXC/UJhTPoHEG/OE0oUT7+rTO7vDawwZBFDn44Dleu9vhl2VA2dNqPxwkC3
aDMXheLt02mD5N2mQsDUVXcIysdOLdIg5btlJC71FiR8kTx6CwtjVmxp3RWv/uOQ86rch5F3tom/
EK4cfXt9kHAp2gQ4woKXO+hLIj7MMc1Bb953xuCFVB6392Q1PEBK7vA2TR/Kdxb3yanVVKb8ENGV
1/anq6fyNd8Ww2I8+MmYQTvPyr68GXZBQr9Z5sSM+IAg1qLPjiaKbnnYKUDQRUC0LgESmb7UjHJl
voC37Ur4eF9P8wljbqQEk2tZzYeN5Jz7FFJpPMGSIwKi536qGB1a/y2IzEFPgXF6jLDE2RLkV/xn
Vya1KvNsUZE2VfkJTgWYk60CEvlKgDm3FC3nr/KgXEM7A8+KrZFDY0TaKLyEaOfGT7cCGbMWQFOc
PVBD5/3MySj5sFyzylqM32fGad+oC5kEIPVtZAhD1eJydxhIEEMXebxbZ3lJHVS+eAtthkQ0uRif
MCz1kf2wow3sHmtrsp6sKGyKaxbm5uyiP6/b8SrthT6Tws5soqup9A041qBVJCOWiJbS9SAhiRkB
zDczD/g6UlthOhHPCeUUZ9REEDSAUey0JahpBicLb02r/8OSDtJm/bjm+hBI+iUNqgcZy0ehAdpA
CJUDFiHfV68JhU1Yab5an5XUpJ0j2U1RSwKYtXkpfuNTal2ew5yLJ5hZ55li3t4StFPOy2Nm8r/E
jiQdURLLdBwxIZieopV+TzcgHSuPZm0f0gM6g94da8H/ra6sPS/QsB8RdDgdx8tZ9gDudFdjWJdL
UA7V9n9kmyThHuXj+fx0nIiiI+6D7IgPwE9M0zb40oorQfwbZoDb3YPrcJrRoOMBKb91a/Mus/YW
ayTtC+sjYyp8KBQXSOdnJldmtmZpdeHmsLngJxvukZjxTKdKtgQ/fNSp3sZCibs9/TFCh6d1F0DZ
KgC091pjd89QJNOo+x3zOun9MLBlddB3xWoi51Tim/smyyslM2/kCoPmV7dOdoLyGxxsd70cnh1A
+xzGz8Nmti4Jr8oLlGJ7Cv70w5Qlx6K4vY6m0R4uGEQfy7TKO6rHCwbUOAnsQUesrlSIW+hAB023
6urd6bSPuWq/3R6t5d96Zyn9lx7eRreIWsP67xP6ED2RyInowjfARXUWBzziM9CFsPwoUMgEg5Wy
6FcmJ1+4FGS7F33H2B9eRrkr84LEYGjMDNWnsDKdwhFYMDYlUckvhT+6LgzQqmvkfwnmR7pZnOcn
cyQ+f4jD6kVGoM9FdbPEngcO6Z0ycn7APCLoiFIs1f2YKOyfFoLeVHQNRbYdyeRerR+ioMWqQD3y
gxPnQmCepU4ncpUhnuPOBx2gIzBhj8mBJfIjBu6813IkmoLlnKhE3pJjGuJ8TQIs96BB5JXDuwKC
BhWOqv+/frYJV6c4VnSZEARelB28pc9icVHliEw8/Msvb4f922mwAA2maEg1KYHcwbVtd0g1U2fj
OA3i57VvKzHLZZ50XoaKopuxAZAKTVhinBSoKEZ4J5mjHhbCFizW6KamRttQdho4IqsIVzSel8Dv
1jdLJMBSiMwUbkLRwIYjeLzK71/gQCmSjYY0H72Xq1W2eC70M7LA2VQZebDTIKQgYwnUUO5uHwMv
HCY6UKgTYBrmGnZmGi59vvvHi0vPkMqtCTWnhdJqDvltTlbYBRgRmD3jPYYX/1eW2SeaDOTQ91mn
ztEdFbkc5Ea5sSH0STx8jYFAmBvOzvdS5Q9BCmzAoVRWDr/OX8qVnXDRJbAfXKvPZJFBriayvISZ
uSZ82DZyyC9q1BmP9MNyfpLTU69/IgqzGTMr37A5Mrd0FkoP1Jm47ZfvJIfxvFhs2rFTwcXC9niB
W5b8MmpOiKazM8rR3zjlati28nWqhU0kEgu67V0+g7LzUrT7MVUItU4MqsGQd+E0zp6NxWtrLTq0
IiczQ1d6jesxkg44KMOJZD3aLL6zkbiZMxe5LJjzZKfHi0e8mvGDg1j1taqP4KICOBCp9HX/g6DH
NjFOZjLwH8au9smE275064GsmUuWfyhNUHE4beWlUUMrNUzJokXYdsKvWPheo+dw/wlHvXJaA9cr
jpoWCkZwv8uW2TW0hPFHwcpDH6PPQ42GlJSU5pj0v3PY2D33J+Ozi2QtnKGhTofisw9L7cw6KNyY
FrbOkMmCbSK6VJF7cnzfVlS2XXiutTEu7lnlJkDUf6ZM7A2wrLEQLxocd1Rit1HnNP95bg0afZoV
DuhMRPaHf2ItpdHJYpW9rT7gvxDwi6ftlOpAHO0WJmG5O0F4NBr9E4KCtJKtzXaDUOSoBzjgtWXy
lQV5b0A52mbdjdLjvhLgnd7ML1NvwzHe2EukDjXSiwHROTTJ+OydVkOi8PJEanqBOuizogg4A1ZD
uM2u8A4N+t5KMEWnCY31UwqWivz/6o6VB6sQGgR1ZxGvZ/oqUq6hUBOXfMIVtKoerAlHQvzFl3iU
aKUyg0sYTAR5zqGWBnAK6BE0LeuEhS+XMSydxXsRnk27d4wrX3sUK0txQBFJlcVg+pHWyLOrKDcW
ljfwNl4shnrxHbP+IMQ7moRRJXJefk6p8mq7d6s/3i/X0RBge9+xz12tDT2zNnGeif1OiuoZoSg+
WvAU8YY+br4kkFgCaBasZWCL78wClUcQYu9dvDps7MYdvM6veqkgREd5hWPJdd25LZtDNdIrM4il
0krzXv1bjunV8U+YikjYiMur6X9UyukKlbxp/Rn1IZw+2WLMD9erR3bnlLhUK2/O2nk5AnE9HKxz
JVcwDHbsfB06n4Jod6q5t6xaqtWufb2mATjgbABa0fIV5ovjrPrufHP0pO9+1+DV09KShSTT5ZVU
TMb1bSGSDQZoVr/CKOk2z/Q2WBLlVehQT+qDWSz4ki12pqrkhsOxGubU875UaihNRGPPERX1o+wU
Yj512wo9+srpqk5QOJwjle0CqaAFv+PsqLpHkm1oRx5/6skgsBCxeMTO5zc/VY73yB3/20Pi57/1
k1IvdBMdxgvl8ZEOiNQuSXNQSjKe/WzoD/WVHxsqTy2ce8gTQekgjjK5UMk116DviKmdqSeotOXf
cQmgPpzmOddxEeWCbRr935FywEjkyfgZbRl4s4z/EP+gPqoKWZNmAD+VZk+PlozknEzP4u6XuQ6f
aSk3hacWDGNQx3DUWtQ7AiKWoKqDpJ9cR2vgmYSNuQP7jlnarVlGTa72NYsypta+YIiDRC1H0mOU
RzKzeEyt4PaQ3MarBEVTqbBuxU5Os9iSV2kOm/YtVRMK8i3+zDBClZYA4eFrTgIJ/PJq0Ud7QGgO
JBX/pAwXPuE96rPmlxwyzIlu76VaOd3jEmTGD5+dH1yjRVLpTmD+1foyBnYdoqFvPdE2DTO5Ervm
NoZI5c8D5aaH12bbBnaZT7CchVdxXoAWfCE6iAgJaHRzMIivtopCtYu5IghJ2NcyI5njpQYk2QQ5
0Uo7WumX2n70yqC4A9AnBwBp6ZG8nQ4sejcEQ4+LaOF1vsQ+iu20tcMrsXdMcqwsyKhq5PVhimyT
+B0VLmuTWWciH+W52LD9RO6HBKdQ2HAVEcHTGUHMg2HyipOMNPIOpFnSd487mbwlpMRyBdDi+d0N
qSL9KcHKbGIS8caiGxcvitWy8BnknucKEcByzLuzdqnAVOd2ymi7Jg2fYtx/PNk543edHKCchOqt
KXMzymoWQV+ESeg/yXQulTLWXvMaVxFyiBCLeOJ9K0YD49HyCUvCtjqe1AvhvzZD8TwlxYZySn6y
G3J4I0wYw8lb8l7EDx7ImPH4v/YvLEqL03idysaHrhIT2C6mVm1qvdFYbUNZv38PwQAZarzlomHk
U//1SXcpJoxNVAAGPLfFTgvD/F8AAmyYT5EsB0TtkV3AOI+Kt9Xc1IKF+xBKgMJXLB0fBGdl5iad
rzXW/LlZUJ70HcKqQd3T1a1NEsMhCOtkywaplXQgdNmJhYmSeYOfHSnXEyvH8RQBH09GwPUukUl3
HB/7L+cBqzQEk0eqbWP2MhGTl0bMfIHXGplTc8uwhG5KE3Pb4s+0DQH8YjtiUZQQPgYowBKrKKnZ
hmPMqVRwp1gGtCr9f6kkQw081F8UOQ054f1FpzCDrHmCTyfktQNDTIgvdeu9Gg6FfkGvUChpfOIg
Fc8ixlWEqaiuanbhTTpGfsO4aoUF7bnXv4SZy8b/h1d2aglPtiw0LM5702/1J4PlhiLzwhMqheg0
4IGKy1owN4JxCSucRvbWS5Olun1Ra6QQ4l1C12ZlF7P3+lgzdpKubutrJY5z8F6KhOeW2C1iRSUX
1NQLYGFLcoc/Esi7Rd1/0UmGwkm2TbptByR9Xk+ImwhFluLuX+ViEiXvpwDec0ds4suLY2c5/wC3
feW/FZnvLhRRZIzlHA5NuzLeKr5els9lzgNUV5/YxC66HEjVVzkeQ9Mhh0/Dqul/zJpIIforVzZt
nMbnFxRZDmf2BIV15YkVELW+5izQevL11nullEM+dVk6VDUjRxfF7bkCG7LDRoz+/fM9FwrOOvOM
ReCLsOaWdaNHvlMnDZeszYHLawZByWMD1dqgdYXAVBQbnmi+yCgoLujdDv+GOc+bZL1JSSJmtUib
Cs1sCQk71uCP4+vRaQJWp2rhVEKuZNvOywE/5BWKw1cSkfaJ64HJ2YefqHlsDtSyyRhd58jhZb08
hWw/lu9BTFrZEgfkkQDpyooUpN9rENr1d7UqQ09CxfovFxf2e53694chRR1xmETdMz/b1vrrXF+t
xoGJYkidnJ1fIz8/ilMXJBB9d7lV3BfsasXMzvNxl15IYjDEnvEbU1shAy0A4IxtJbU8e1LmTaYj
88s52dexePbvRmFps5KEFmxLA+OHKrbM4GJX8uB753CodlC30gaUf/yf90rRQXrZXzAty0YfmPtx
Uxqb4KU0M+f6hKUAMQxK0HlG1xIFGmJyr9SSZwb2YCiuV+MjF/Y3cmEPgsPD0fwh6hGxzTnvK0bl
pFAvbapLcI9z+rzmWbr+kQvypf8Zy4MMx2R3VMxvK6vlRE/L4PKNIKrgGyFi09+MjKdCyZdxfIh0
mVelYtonNJEpdsvNiInZZtuet1g9yiMZTPtzX52Sj/Dg1QNuOpYzdeTM5zPrGJ/TOEcUVn7SZe+0
wr/9541Doby60t63O8hT5wYZNWTbCLiGeWVUCrly8ZNrfF0yRSx1vN2ehBXJTnv/ZXoOLNmKX0uP
K77BpIIL2UOBaYIvPkJPQCVn8ZIFQUpVom0ldJmJnbum1wsgDtLbx3On0bor+8ApwSPQ9ekpt0wO
h273ZsQzQ8pRa611Pk/3ue0H1PD/SMfQxUeIcSEDezxQ9IDT9eeTpL8WK3oCxOjPyQWyxk/BweEG
ENRIFvqJY9y5k19woA+F1ltWy3rrdB+ApV4FpyTeQtVrC23RrDGKyP16VX6dGW29+DDjFoAyhf/n
d+VWxJGpjpmxLfCg5fA6h+KuvbtlQ2Wu2RsqY5UjhIw+xg0ckvf9UKQx3q/7ts4BfPlTeZ6baOHl
r9Nm/BPWTHo/N/8dX8SIShP+UsqY01zPHx3cClksZp/bZ7c6qlqXse5J1mu8Zb4veoiso0/To/Yh
nkc4Z2GuN2kd/KB6RCjCKCbUDvMBZ0j+j8dy6rMdfTu/FEeIK7QMFupuqRVklKRKgl0gvgRbnM5v
B3NjYRGuGoKWadUt8pCqG+tiUxT5gePZPp0RFRHAKIvGeL69nwliUG0udr7p2Q/MOoIPdg3UStDs
RKE023da9kzbN7KnSpKj8fTabnDS0Eqcpue7Kl6IDyehije8SCBZs4o5SnHzqEByr5U337NVoLJi
f8xHMrvYUeryJ92FC6Rve2Q+MfNXuqBpFQp/GUPh29uGkCXRWwdw4Y5Mel8V88aeJglktmEBvzM3
Sxr8c26ZLB0d+WGUwNhFkY8T43fOYoeUMKuS6hKs06WsNdbxg3hrk8zzVXVGym1IramCEvvAsZxz
Ci45UXjl/a5JJWzT/byC7MnN0y9xzwY1Sy9leGDZuhsjugFHuRDTYTG69w2bk3WbIG67cBXQWfrW
VtJ2dTXsiy6KpiW8uQ5XXuPcEX0z7XLrQNnsnc2HKH/ufTTrOGLTRgIYsbvQWjFd20AWuq4o3zUY
S617eNbXOEOh37dhC8L75ABsPKAiKwHfEfdkjqVR8dKfSM+HoNOeeAHInqDdnxMyAptbjUcbtssd
6Pk1vUQrLhBTGdHfTybQajji85oJw7Be7iMnQLEmmeol7hQ73GNz2Upf2Qgk48ppEbFd6bEXIK9m
GrBh3BxJHphlOAderIx2tiViWP8c9RJ6K1JCiFe+eaJGBd5VxLiRga4Rj0hGPbuX2/Hf06t1hFPx
yeUrdhvbJ1yKBTKoLkENphF9WhSmVZkAVN4e1OMYLWTHfMPj5VGXpU8YZrm1G8fDWp2kgd2aCzzW
M03qZ7aSAuZhUUs+WbJ7rnKv0CbP2Q1YRTt7wJEK7dYTGhfWFRaIxbX73p69I+xJB4Gnw2evE0a1
RXMx+jOR+RYNAB5RJ7wKVPhafKvdwHl8UMwqD5wupiIu1kYpzWpzn8hGD+3Agr727ntbPIGyWePS
zyfQhJH0ak9I0ywS07ypI/eE0k0MmtD5C47HZKYRg39gFdqAwjJ2q299N+anGk6JlzcUvZSBtbPe
oR4rzjS/UkaS+NfwvJVXl+W6eCF1+e7NMsC4Jtxm7yEHeFenoOsOO2zfowLMss4ZPBRymNUYRsPo
Ux/27Mnue0ZS869GCqJJUI+TbsayX6yapcZskmtoz2N9j1uvWa3lir0QF+Msi6VGhh8cdytbiKyR
fa7WE5aPwl29vgkyTxCxvWHFYwVNASdVw7BCJ44gXWywlk9moJMREVPRObH7FdkpYyZ7DPPR169I
2hBPLof5HQ4Fnj4j4N3AV2IeBpGdWNHbzkNVviqHrXoS0ujn0NN9AZM0gnQIk1vOzLc8HKfCbcpI
pLTNDZYHeW9yoeh+Nd30pJJexFE2ZdQZx3w5I7PuExBKppGIw1GUxh+I+/oN9lotBYepkG0OZHf5
beQbRKKzSf80m6i3lWwX/YKdL6NV0xeN408VuGBRhHZoIhayJLcLEu2IQMeXihgM5Sy411/FC1VH
QKyNBfeW/LOFa6CGZREL74zGyUrfmiV1ADvBbaWSK132HaGFH2Azx6KE2tF9UxauqBVokGDm8ebM
CBzOtLWImEFqUdkgBfSPbNicHpX+gzEwtKPE0u+Ogms/pDB8xMpGS5YXj5kExV2+rHKCasjVRLqu
L4xVH9hRVeGgX7LWCUgab4MzFmKafknR9F1lHpjs6cp/ncnk3oEig4la+YhUXEoQT88ywoIH4Ujw
+ExNQbEccUT8pPsCSTL3Mag1R2kNEU/z614fl/1PrraicXESD0yrR27PAO7bOTqBieyXPQsWQbWX
dosC51qeyhrnxMoX/J3Q0MsfVZ00Zr8CvacbJrpUpi2I5jcHJeV6xfDpPAWgNJV3+LX9WRuhgA66
SlD134P6Mudd+oslSqVqygwM3/zv6BCsK4KQ8Rt/+Uqc7YzeKUFuxHaWuSvSLf5emzWftuANcASs
EES0V75n0G1t5SHfbffBi2dRGUVrwUM6KnCW1Xj1FY6Z32HrpTiJ3tZKdYuDXwt7JKFySSmwMbCG
vv1epYZG1ZT739LC+Ly1uwzZMoJvoXuzc2eLy18PJWGyif3FhmOZHLiIkBqLLA0UdkMyP/HRdOoE
/EOCOpfHXdWI5jgzB+y9xX2ehWiBVGf5gqs8BhOwstNrjAmqEeDPd3UWD9ZC1ZIuqjaE1OpFYNXO
v5X8ObWk3XXExVprF1NQh8pczeU6V0yMl4pcvO9F/Iw0iwRHY3jteQQydec01wQ1naaxl/cFFxCH
rjnf3GEo43wrc18Px95fVr5wL0xhiE5EMX1uFvoLA5Bj/CBrlrELm778UhgBGq1wGFtDoKJMUoF2
k1tOnk4m2Ft1les8WPFRB7ixGB9/IJegAogGSsXcFQHk0fulYf7cDgfeytYlQe6mvrn5C5DRQw8n
gTIrfInc6KKiNcQnlX4J8g6L2OPm30HPgsC2C/DNo2qevZsdOrBeyZLd/6Y2xrSeSTccJEsssj0F
2pem50BHEjbudsIK6J13AWIZ6wPrN9CKDjQ/imsqi13uqrUo16IO+h2MWKtIEyTJYrt8C+PYET1o
a3NGS5rpEKOtklOFsAFBn9hmHPR6OaV6GfyLt35X+jIbgK7D342on9ZEr3js2Q7xkHFwxeKhNNaA
VWN8VxDYThZSpVLDt17gHIVTnGK3YP3ylsiatBhwR/wQ1ee9pwaXek2V2pmZ4/ixCGRGPsWr7sOn
HzKhKPatY1GN9Lmlyrqm3OUy13Aogn6IaY3ayocVZIuhXw0VqnrZJ0JK4P/0vMmoFUteAu/VLVB/
uTNTHWDL+GJhJd6/Stn6bV801zjbIGOlAUJgim8r5jSWgDwAWAIg++/cPxv2fubE5planDY4hjMB
UmypzwWNmUMqSwAln3n8/fCdFzZosiQqqZFsiwXJ2bw6ZkvUvd9souO8l6pwM/7yKueCsDT6dSY9
LF+6H0cQqqsPZx0p26mHcnkggmyOq5cbRhDfJ4r/PVBxJR78mn/4uqG3ScgcGjykzqtJQMELG6Yh
22mAaZL0/BqIP5sbZrvCHCROr++1LaaGe1TRp5gZSAlHS/pj7p9d3u52OOrXvzhgsiUorm6wX7b1
mPnVSjU+v9EwOk5YGUGFPHaWwyCJXu9rc0l1EQ9Kpt7cIYC3Ge+LAzXeJcsMuI+Mk1dVWCFDuk7f
gJCVRC6X50lUU7fUz/Y5hA/fB4CAQJBRloHlYDPyfxQNQJ5G+W6ViW37wOFimgwjHStLbFOrv+KT
NHKSrvQQHnMfhs03rBz0JGpS/bk8wU05ESaEndRtZVJocVc5XFoiqWAHK5X9tpMKfUpWMV+7COvN
1qMOd44tuVF1gWUEvrOxipaWdAFsWl5PC4vdwE1K4f+SMDArpjcyDCCJaw5PMrAE0dBgVVvyas49
gJQtWkQgW1FygHOVA+alzaLfyEPeDzCpxUzS3F85YHhDTHZymaG4Eb9EWnt6Olm/cLQjM4crpyGj
BIQEufbHJryvyxe8IqwRUaHZr1jW/eu3VDeDjGS4taw4RR8B7NupckRYEG1HQ+zwEWS/05v0/iuw
QwtgYX+lByYW+D2WAN9fQPrH1hktVcXQg/dNaDsoZcBOFqzQ0rZC/4AAbhpODoVQ1qGY0ZYJTDy1
Ht6QS3YvS0MJajYsOBn6Ous1uCvVi1+d0y+jpeOBmj+V6rZiMuQmgVyF3vSVvI/4kayXagMbn5TS
dRH1hBcp3/C8J0MqawAqZpk+RSCH83GqTQkxhXthaumg7H4m7lQr7yWL8B5R3GoD1qo4PHjsrMlY
srE4bdL3DldIN1QPV4+pYBCmjUi848O5lR9BKHHngxASKBpd0w+Ckw40qWRg3Y8IrFQxOM0bUk2u
2knVLg2JQbnqJ1pfCsrL8fnKBfCtxF54xSvPv/wmJ45AkGSPrNuAedG+uz3yJVfUPz/P7fCVH498
PRF3LkFb1pBAaQOrTjJWCN+vRNvS0A2fiKhqGiX3i9Lh7U9besGv9XdrHGNk7vKlP74/Dr+L7XKX
jaf/wzoWFLodrbEHTcdwCzhdPtFgAw0CJXvn6vg4rqpNmBPke1WyEksA4QfLsNvMvSzprKnspLBa
Uw6RN33yOejMegrKDK9frRHhtbdtz/PLvsBaCeHLKyV6Xu/3QQxKFnNHd93lOVuw93xZz7XqSOEr
evsu9FrUVhcrqcN47fwAqNntOnaNh1QJk4I0WqwElsswMOEEcaFVKK4qxY/dLMtlG/wNHqUznlAr
ez1pvIDtJ35LHCleAbelXM4wfH5wg39izSuaf+6fqECn0LhcRIKLf6XDvd/B41nGIUZvp36iZFbf
rDMaxIVIDYjOFfc+G/nULI+l8XO9MCfHkP2JDjBc503K22nxk9ue5CCVDjh1pm2K6uv0fvf7x3qC
/FIfWP6+dEUjlxhz+D+m1FHV/MesQn6p0/r/9gzRXpx64aVB+zLhZfb4/XnMdzhRGniVga5E3eef
hBoGexXa2kqZ/DvNfnn6XMQJFW12h1G1DzTZTuuIL7DbzkMNP6nhHqWnbJyHgFCOK61BOvyHbehb
6CxR5pU4qri5+HRoAeWpn6DNgj5NXekwv0fjC0/m8Ad1+m38G5+jIbXU2M9RuE+vshQ/czPaj/e9
5qD3ya5EnMZW1fxM+CfzHATrvRfVt1RilJWxZHnwcQbSS3UsHO3AushBRWzYo2WO/Et1OabMF0fb
0tBtRkdaecpk+5zdxidxcOy3QpMeSM0IfL83JydVFLghOftrrovB2rAQYoZSaoEmvBWWc1mchaBx
FZU//j/IoRTS36Q8hKcGAesrwGnm4e7RhfpSFPhlzmqG4kNpRiBmKIYmSEYDR3Lv2X4QxdSej0g9
0ybjBjqKS90q+xToPH5ALwq3DudVsRqmy2WvmMofm9i+3f22ef6ewsc8xIsDn0zm4+lNcHLvtgs/
AexGA1wirpFdRMcqVJ2/Y5I3rPzwGfIEw2W9Vpvd695yyJsNXTWJvvftekm8P+G06UynPoxygKQh
IGp6CjJ4l3mf9tv5D1Cy+cnyiPQtSeX49Vhu6TE8aJCTGAHrBjILxXMFYzg/4AudizHSylE56UEZ
PocnIH3Qm3lgpkgaFI7yN7nY223rHSMc78dKDk17cm7pSMZLjO8WB9ss4yEP5L+HF7lPpaoNgzaN
uIWdthjxNrmAM4Xlay0KC7XOZUroSsksyFQoLFtzk3ZGUIUiKrSeBorryE+yc+6QrSY9X8YF4kqi
uDuBOTVP5nqODb/AjMXsSkdafA4ltEAyvt4n3mmrQMaV2UY+uIt+F+wd06mQrvkj4enpIM8893G3
MCAH6Q3gTUxGvJEK2oMne/Nw0yk99m5j1FGAP7NHFbNqA/0b9muROXk9fUPVETX4iqx75F18P2BT
Zt/lQuzYL0mGthtTA9x5Oa+Jq+qO9hMs/FhbYFg7O69GzP6wig+SJUk3X1pubkinw3bAQso9i6Y5
5w2mqVqdbFUR+f8j8Jel//ILJBumxrlr83Te1/m0OiYt8QlK+IxNXYG8FZB3H9MyTVM2ikbRpU5S
SR05BEi8euoYYx86Gr3yxUEAlgtTKKRlKzN1y+gK5ggDa5OBj9NJZvZe3V+hjLP9nyK2R1Hg5cUP
7UFZeo4pLWaoNVtuz37b6+rQCJaXWd12bEB6dNzI8rtZL6J1qsyOjGVfrYaOsHKaoZ2MY2EAKMrF
p6wT7Ii5+u+to8u9sC6/JGyiDg4uqA4q92xNHtI0lf5hSPRnoDKXWcasfrKt7ktXMh8u+NM+by2y
IVI/E6DE2ejk+3wT4e7lMTButoL626Fc+KU9g2S6qOO527dx6UwSwuVmrr++NHmvKAfbuMuuHY74
YO/AsOV1kJsn8w8Vnme01HwhKTYxKWpvMLKIaVVUsyYMhMAYY7R93iOe/PeTKgguYrbbUC13xTK6
+GH51Oz6uzGTMpEUFIdZgTRxbwvIl2jKSsyb6Be0BkL5Ajf1wtZ+MMWHMRk3N1WgM35UoWiDCx9s
loX0w3EIkefU9eMsTpmY3pZhHX1OKosoN/5qkmEQz24isys/4Pbc+jOMM8YoWuNKvXVtddp/M8Tq
VeMIejgYz6eu8DIySz2nW1L3v8aeYBOskdRNtrGsHS3+kWMtZXE/MOUMDu1kkd0WAhlsG4EXvrhM
8hK/zEVgaBJQ6rOWhX5P1DzNP77sIvvjDB1lplPKnyrWKsjfhaB+B6c4AZo7hewfLIKkESHppqPj
46LWAWuPYnJ/j8lQVWY9gc46+MWD4t0T6Xsl7TS4UIbMvu+lJSmUFtoVcku7rV3MwLF/MSKQxQfF
f7NjJfOxtR2Y2fO1wryGGNn2KB2gpl+clfkwepxovn/Bj6RMCf9KemyOUhjjpzOEI71+9LCtQv6r
tJysTtRSwcUzBEByu+uSMR6x2cytaNLHmKZe09iHtrIAu81MlrNoBAEjah3ELohPULTn6BaBtbSD
3gBZKG30e+LZHlZb8KkLyBtm8GXkrJ6Zf8XA43nXtC16JudsqaztIDhotsq9vXCmQHFVMFLqvEc5
FlbKlhuFUwrDKolOn5flmZTu6GdM2hQ14/2FM3ZqBHXzQGMEDAvK0wyMOu3BSREX8x3vvbdA5IdW
gpFLoat0ANDFiPMAYleRV3vK/b7/gC0ZU5zUdSU03mv23VQ3oE14WuPuMYt+7lwd7yaBkoJibIsl
sUT5zFEf54nRpwTH5jrkJZfqi9iVbrSSQKJ0HBZmmx/oMIoH4mXZqOHA6O4E6VQL936679j6NtjY
0SJeilVQBqJ9RbNVGMgCuL93H3ovfnWV3cMt45uef1+JcFwNg6u9TYerP2/mJcuy581CUGCuFk2E
/yuOziH4p7esutjDf0vjTsFPWdadzVKFzESFbaDGkQKfBgNAPuuSuonTaMSGUHltb1WpRvHxA4F/
WO3AzRhxWZ+iKpcCMfom2sk9JSlWJZDamSfxN8Gbb6trzcf+/z0ie8/yAPGrWfrIHWDW+Pdtqee7
MCVI750LItEIYoUNRIZgbpB442oRHDFvI6qIz/LkNe38heOo3pwotewT0hdnNhvtLSYbW1bWAqhV
f31i4e9U2FXgGU4r7PcKLhhVDV8iBONvqcYQLLHUTyPT2VTJlZPAy/pHDMkQcWPKavYxUkxqWxAw
oej8KxvvRtNyvR6BTMvrL2RGeC6WcPxtySQCVh7oPs/kcbZmovkClPmXHWM4su+niLeRK9iETvYT
Dm2Ny47vVCd+5EhtBSknul3Vy/2O/2EoukqE9q0aoEZSfsL4uoNKUcyofX3cDRde//wbVI3n3MTQ
OGMlc6SYNnsregugEbCYffhN0XnaGY1XEGoRlYh66ba25DZkM1/1svjXHu2p7Soi5Ss/6PeHj7WY
fePCgJOrVGFuJdY8GU8Uvh+MoCG3EURMoJYJA8tigfBA3rRQww1eR54zDnNmFSn+07CNx6UOqUAr
bgsif13QUZ7Z4QMTcqRbB0wvIlce0Wyc1ZRl9CNUsh7KJ3+VwLBWSnMpV3/xuyODYauLQRBfVtpq
9JvzZRabIhG3N5YBHwzQTbhxt6NF+Ml3cxJTXgXYLU/7W0ovwjSqu9ZpNLdNzcs/e68LVjTzBCVf
8Zk4eF3ww/5cR0VYZoL8SHMjqSjoXlvoR3Xpy4FXKbZrH66ETZyy4uiQDJq3847M79FcC8EKpjeS
Xi1Qkcxnu/veCnq7ADi+Y8sfghtr96FfVMxiKL2r9iz0al1ZFN1hmiTpJ+Y3rvRXBPDQdPKt0iLp
gBgc8VXPdIffjCtC7vgxfhxHgBAFjIn75HzPzrfvt3M9Ydnn58Rw7KWXyZqCF4TDOBUBAzgVej87
UhVOOYJHpqyOhvJUat/6CwByhlvXx7qoWOhh49Gj45DiDxLSCI9GWQIQ5vflIZnK6+CqfgiRJvTT
kxztL6HepA2wgoCyCCgcINbBDrDt2TtEbR60DC3X4uf+XuHujxXafpmaJPI8KJjJP14Hz70ByRqD
hpWpBT2bobZY/tDQV1GwoBF8AzK0G0hCUTG6O9PkQTKHd4qploAPXaJN1CJEN7HKGajyzWPsE7DI
XCEXDNv4UxbGi68wL//KVmrx6XsmxXReJu7Y0pyMDx/KxBBOZo0pRreA15JebWqx4nBF/vmAFegr
deaG56ZWPgdBi44wi3qF1q4m9bEEmyxcCGMkcBfIhlG0+BcXzjy7jnzFMhnt4iye0uAv9+lnmbpP
0CeO2YFUhI7uZQh0ZtvYzTfsstCOsDiYtrE1QYZA3teHVJVaBZEWt40j4cTUuhEv9uQZIaDwlAMj
7Z+hmabpWASP5UvlA4uU2fPS6WMokUKW0DZs+Xd4g1AQamEG8YL7w7SP3VOgcQG9bdLuokKHgf2C
H2XRggdf5yXTUopd3ge+6pWGDhy01oE9EyW2+AZVWM+aqnCexWbhTCwE6lT66n4ajTFoC1+DR/sD
WJTp4VrP+X4/rcOsdzjNPz9h+/gRmBe40XUoHiPgqfPDFL/tESkdrQMX9+O+GIFZ8zjMF0XUqnhu
OraJsRLJJU8gmGkU2dl6DsHpA25kig9D82QQrnSBgCSN/wbx0UHvC3FCUV7xd+M2jL/1iYCLZvva
34qKnZEPWilV0Je7Q2h0h4WdbzFgCo6b7mPWT0q0W+jnff2ZavAQi/ny3uahBjTipqR7tDVBYojN
Q933fdPLK/vVFAbH2jgaE1f5fvArru4BS7L5ZKRNK7waAuzDkvgzITSXm4q774AbcnJrvPVV7x1y
njqHwK9aIMski7SQiipLVIT03i8FJeEl9xAvxPmxP5G6xPUf3E7p3se4k9f05zSRlMysc0i5LCs8
TQUnAJ2QhnlsLIbjdF+S+HXrdm1fjgTwJ4ulX9Deg4AJ9TEAGwYqO3cHYEjsdP8kCAA4pr9d78c2
8SPbY7YBhG+rssYU1jgRNlOnAmJLSmtdBAegYimxe5zckv6zXw9l/kVUidJIJd0t4N4anFPCyPzn
Ui6mbhF1iwqNpGD2rCePA640R7p5mH4O09h3hBAeDXkjMUKrybmwmJKjsBpPDtbFBDXs41cxpA1J
CWjcBUldqE3ePhBLJuJT3CP3NKY3PAJC7t5rOPoNWU7Zu3hE1wE+aP84o02+nYVeI1/Bv0up+bai
euOeueLdm9zmpgJ34PegIoaEDy8mMiAUCNfF5/sImpBhbIWcgTeeObAAQYozHXcs0xUhjG26jKEV
DvDlPDsUuet6fQMnWd04wBRenMfbSIFoUmzoLHsE9HNS6Q0opVUNF43xJ+MWAeoxX8BY8BYZ3cZL
6FIvubHiXdVR/QagYqy04OjsQjqmvnlKe231Bm1U4+xu6x59DRF+IHY4fGp+BrTVMRVe83bH3o+r
BVCeXEZpbecXWEV7rKEO9YOy2RPyg30OLM9Yun7qGxsUpcvrsAQjoS01ePkINeiWNK9/XGKvUr43
vVdu52zpGHSJeSixd1iByRj3rCjCrMawYzFzgAszg9X+TQmW784F1Fjf9PbHiVM0hB8hTPBsrOu7
qVKT0uKI8u3Sie5Sm4U6ve3MAJE6oAXDNNZjn/s7xi+5lGzBFmgicbfHzv4dtrJgxy6EGjZdvYk7
tAqkSggqeQv1gw6c6il8wR4W83myOqr84f1ok4HbscAPxVhHw5b7uDkteDBETmXSHa8IvP30iTbA
kHQ3I3cJrAMQJzWdGKp3PQf5Xao+TrA1eirF4Knwb6hIIVSxnrk+EBtiYJ76MMe1iLfhCTTSxQj7
mZ1ZyvG1IEfowrCR4w0/nUiWYkwJNoba1n24D0R0H8XPacafzHRMBVGXeWmqYC96afCBe7RwzFLh
4JqkKMU0P9N/RVyy1qblNKB1TmhTtN/YFT1W3QDBHtb9E6qBjBPsWUe/nO8xEwqepEC3EJa1w3M7
YNbbcXyyORqpWhm7SMVoBrl4swW36IQGZ7JeZzV9Okh5G+LpwoZfhtoCC9z/2HynjP5uF7DgIXjM
A+ot2nbHjkLXTtWjkJY2n9W2BZbD/9XKhBGaq40VFb3cec6jXCnp0HvsX+UTeS5AmmuFu1NOg4FH
jiLdTEpP3sP0pC5Oq134HK8qMkhMEkasIL8t8FzxvnSquvMf14vGKatXikSPQKg+JxAbWj5YqIYG
EwgoUcVFRQ/1N5IQUDu0oUPVvGgGBgbLTT3bUIRfKSXjN4vRX6wJwCyfD8CS7nZXvAU8jRXDpZ2D
ar5B1QBtX4Nbn3ebF2iuetneF1NzZOpZgd/0ScmFApSyBzJ2r85mPxnhVsiIOyhYiNsnpRZzORzi
5zB1vJqb0vQYy0yxveetYCi6EvkfN0vudDX3B2FX5clW5Czww8a+viePsQFkRZkB69wpNmBaXC2f
kvS6UoWf84N9QOHegeqhj0B/j3JVpDMFN4QdkjnjnmUXkZErt+SSNDdjKDhOEIFtroAUDq4+KnsU
DUz8E8q0JxIdujXqMCKZCRCJd9yRFP0T78Ecp09rTrhDUXYSUULhvX+4XbrFN7KivVtMXQehj/hF
rikpAZ3fqU0vMvZcdL91i8cIGo1lGUP1P+SwnyJib0/OQLGKoP5nAJtSaLrX7cyMSfeEZmf3KCjX
5v96aHYRi68sGVZBVuzwlyKivYQNce08RsO3GEVg1DnXyn218Pi+eyUZ9jSTCu4qrZtuVyeQu/uh
57EdSjqNkZ85IJElAVyDu4qgFa3Gbqs7EhvqCkNvMwzhlrKEbIQBWZZpr+OFXYqaHgDejl07uGN3
EZGPSbnxQN3JnkTiy6U+lDTMM973GMBE7Ly1RaVt4MUNyPfZmquhmZT8Dc5WKGSeJ4I83HHOlsYT
pkKgKGn5aR2CobKNzOAGFNRklMIB6F99Cr7zzhEig2OhHzrVFppuW/7QwhJlOTiNEUuLTv4xbBXn
yB7EafxMHREVpi1S95GJzEAFtoXkXFjKPu3oSx7E5U7BAtOJESUaQBZ7LjBkBzwsgB8vDkdkf6pR
9tPlJMmkSZb4+7IvwNhm+HiuIyTkMacnGwkaXq4zwaMZr5NsEq7Tl1dmO9lLWIVYU0Y3yyX7iTWq
JmApkflAhkvnwwun7wkBTYqn/QJCF+PeLXhxmEk3ousnu55gpUKekt6KOmaYZXJ2juyiL/o5Woyq
6GdSTlO9I5VCkX+3VKUnIAtsGrprXKXTsCQXh28+ZtpcJh02Nkq/Y5e8ybncHQXewQOEbyiDgkIh
YS8B1fvuTx+dQQqmPX2XR2FSD5s4tidmDSyQ6c3w4GrxP4Ok4P1zKNLy46I0JYIlrUrpRPu4nTk1
f1gNbzpTCoeAc4muxmzt7zjuWe0SigkX1dFgG7US5JO7XRHjUedxbiwUuZWVXMLQ07acflXZ/yJW
M9siZAkiIoo+M12u2+c2f04ldMd3Kugn7P+W92Yum82mAZF1XptC3TD0hJemFMRaw+/g3BuZAxoN
CtcNjYrifkrf1MDbmOGPl40etfUWE/dBA7/aBUtg1btmfh4/N0eCfJjx2h7MibSAanafUr8GP6dX
xrW0ZIvvapRfFnKWIL4tKqriYGol8dFbSBAz34NU9oGZTiDOePbXddGl3kRmgZ4ksCBIfXvnpSqP
scJiO0Ieg6KoTms/mgepS7R7ZVvBfCZZjM4a9RYt6X4NR59T3byX37l2xT6X8lx4jEcoS9TEOKEU
eMiD2d9sctZQGAGgNKMZ+Bk6QDbOouFPFVT6EESq0XO/EJ7n1NblS6/uJ3yOtQRWVw9jKegDX9lB
OTVJ3jJwXdcuNWnUKf6QyWuXFpKHOMTw7EmOFnVLx6hDwTLIu1p4nYXkKiXvJJe2a8ad1NsegsHN
iEg7NU2o/5xXyLcNXjxHT/4H9+sHSoQZOD3GHjrDBQX4dpgCewRaVj4euOHZmVWklZmgFa1b1a73
lpWe8VSKgnDdFHJOk0RwbiZ6CKZ2GUPwelNdZPscGVumlwALJJnK8ycQctBKbnZla5JwrC6qDmHt
1WQ51zZMebWBkY4XRDIZ/9yTS6ak2DaiBh1qpvAHvmyY/Oe2ql4cUVFQh5zS3m8AA4eKsEB4TU99
lY9ISLmiTR1Qi/RXPpe1BPSeLc9jfZhn91BNI9dsT9VKsB/I+YSx8BSws83V5oHKC6aG/O0KtJ3s
U5GyUM9OcxXmD090dbOMqrR9CE8F/XYdx51jFjnOCrqxRYs6/iboKWVPQAA0OCuZPAr6iMt6buXb
99OZqThraXGvE4PN8zAEmpOukJq8Hwj2VeLh2yDAmOrHrYCaMTP05VAdlpwGVpznCaNDOihsi4qv
5bkG7/F8OD3NlFtAhc+fZpXIc3L7GFlEHHYg4BEV63iQfc892EgOSCGLfxmDuA+uRxZ5xR9kdcod
bUB5PPmRmtxW2paumLAt59eS7IQ53BCTkvh94ucEM5bGAe+s0O+X1QW9WWkl/KnYqnO5gDR7wkA9
opPMCWgs4Ec+2ZP0hwSSGiaxj7y2+pTWBpnZ2t+LgIJCnqFQgWztYc7kpR6y+S9DAn2iuAgPRApE
6IEu62dzx88kCn1clFhu80X3JXBcfRcQodU4gTI5VjYimpLA4v+6yD0XtWueX4f1pcz1h8vLZ89X
Y1rMhFFreVB///pZMLLjo+pCu+Ln8JLs/N4699sBDaFzW5ao6+CoFnO2/09iO9Tm7TconcK+GUbg
RWm52V3rVrXvMcDZmet6GXYs+yOGAEz4C2pD8CeLAcXk0zsvjaooqLmMX+CGosnJOfet9b2cW7zH
5cU4naXbdnAX5o5TUfPsB2ShO6cS3Ohcr06FGutiDCGNz+eQGoZYgeqtUpmT+EY1niykiGiZahW2
FgKDP3FUztswGnFQ2MxAMgbZOv7Ary9OVdJHu9ADg5zDuvLF7qj3aGPH2qwoBjsl3ibtgbZ2BKZ0
WTuYPZBcAGCxpDhAPyqNgInXJysaehfPs+SxYhD8JyZ5zzPympn3DC6KwBneunwTAkiW6Ovc0uxk
WD6e5NokNhn4MpMtlsQIbRAc45PiJM0OmKLlXjyLsjC7NA0zjDCeEr9e70M95Lp2iht00VULAmK1
qxWw8AvgCf32VE38aB7XvAzM6IIJ+Th+WeAeF/2qgaV72BcKphF8uBaqqE6p4FqCGK5S7vhGlT9A
tTbFfJ/eHPVgNUl3Llv7uOI4LM7xqjgkZOnvZ/zpZe34zAlJYLDCXWZ6yDghnweHp+x7r2lS5+TG
8Y6nHPER2V6D4zjdUq1FFQCv3kHnJMhkHMtb9Qw18vhX8g7C8KKad+sskvJUz4FjxBC1YATy0rGv
/azCPvxaxUiLyMaD4pJ8h73heYf5e0Z+rTACnROwNo9HPMeZxRiPt5ouAX8a8SGe+7Saga/7R3Ms
S3ZnYR2EORb6dDFpLDqPQRzazBDW+MvmTUp7n/49YRZzl59S1UKGE2MmObEP8H+Zhd06JADgCwUn
JAkDgBodED/CS2U0Q8AYkYO6/840XZARm6+5rsMEFQA9G7izKE+zCk1Wl8ByCYP9w0t11aQX/Mbn
Ow2tnJMmGpEyeN0ckPt8L/7lcAtjkpz+a7V4lPT1iBb3QdZKSrL8JeZUpC1UvvJl6vJzxrJ10AcC
pWPHalu+I4Yl2yVm+b2JfE7FhSZQyJSVGeBLkIkc13r6J8r7ZjdLZg7V38Suuhom08aG8R2kgrA0
tv48zoDrZi5TmHEcdSrqb4/mCsrXR8aI3yC+QOQWqTgO4vKpV0vBIdje+WQAYeD52q5c+a4eNjEX
wAL9DL6WPCiMPd0kOM+X55IRWrpuVRXkrLTbzCcDGOtDHjeUzP3yPuG1s6EWBXGEORsaFOnHDWn+
gS6DgBCuILYAB/0lcJvzeF+md7qL3rjeOmYsXK2RAiLP8Tu5VV91zAtQ0kfj6TCNaC2Rx/AiSRTg
ah0B7T3nket5+gz80BTxvXDyznqYoNo2shHIc7sHFKYMILaJpBJ7bNcte9G55v0IgeAhWlHEdaZ0
he42TIszSGxZDdmczLGtAkPAwCWzx3LOlPjsZcdwzPsM7k6D9A3led/TbzpLChz89CWgCts/WYHi
jCs4OqfnlfzYd9t8w7R2tCoYtfOdPhx94jIzdcpbNbC5RQU8tmbBZVKoxAEEpCRcLZVMMUiHLYoI
QSMVj7ODHKT8pyKkwc3S1xWXJ1fkHcLjYXrbjBjW4EkJLb+i4ahvSwdPcpF01yzPbP6arsGZMxQd
GTap0aYNGcPYXPoEkz/mY3myj+Q220f4paAFbp0nrjv9XHmRNLX6EJrmkSAgJX/byHSPEwTDAgFs
l/Exq4wPmITDO58QHn3dbh/Co6Ol9Sd0MrCDgtKrtjyIBPJ0mVcnNz9uPdYWZTOXF0lN7fISJPUt
MtHJ8IotC6D4qAl3yMkDsybJbreR66w8ApI/ahJbIMdnYPeU2FrbbRp3LMgLjaVVden/VSEAIt6J
WX3mhUkEhZlEypLVOF1CV8Tp5pHgAZyZ9pDRUyW2O5QrbpjAG1FnLCTs5PfAtoT0IFjaXisALB9A
HZZNkAZhHMq7P+Alhim1BB14bkQMedPDhWaAF19gqCZJDVYnESg0sPiKlSqqGVCF6Jl1tJkzln6u
lu/HHh4D9Rxl0pYRnMQOAZ9mq4bYPd7zlriZnKPe6vc6zz53wj/E1E/Ro6Xi29zHxOXjO81cC/2K
NroOvPMkgkW3XdSMMgLVKfSXrV+kVGMwkDOzkFPkhS9g4u/lRJ5/8OtBHH7MczGvU1/pbA95JFvP
QEO+99P85mrk1Tic1mbFjatwBiLQaKhVZqepDjlGgCimttL5Jc2d6GXlQoVnNKIJpWUl0rNtlDon
6aoErY7rRc2lGLF/uzB7gC24YLjTJJ3JZeyWfx7hLUCdS5znQlmdTFLvcbofDaB2heQSk1xnYX+R
oFTJF7YkpV792YzwHDZ4QlwNQSJ343pPnWsTNM85Bjm+aypx7eBB6A1D6MhXyP0dgPw8ufrUOqBX
mCasJzpGFfhCTBxvJ5PofO/z5cGG5O9K4jbabGcRPSVaGz0VGuqo81bQeu64rv0SMU+FpJW9q17m
d1FezaLlqsD0TZtAJKCqoppv71xIr2i+vuFC+ib/maaBxlt+SaRAZFknxHZEAoBmK5VVPpW35mkF
l33jZ2qiO0zVmHhGpDuiyWtQJ4rth16yWf4UVOYwj5AzFMg75yBYrSg6XHWUVcdHcuxB0/mLW49t
erYiWAj33Yn2HBeTnhKq7Qw5y903csNPtvNsjAM2IefREPZZss09bILotnXKkh9IbGg5L0ETM2E2
/84xMMLCAS2baq/FM0wKFBxnkHxwtHCStR6j8Wb4f4GWDzv+AfAOInDenf+hkO8EYDEoV7mwAg7P
mMBAeJ3aeh02mpMSxCZLF2zUJjMf8KHmLedm7yribluJmHpa/XZmAxOslJhzD5nI+Wn4FdTYTq8Y
x0PJgTOlEn/Cy/Nd725Lb7lM2dgvHExWPSrwziSdNbW4gkle88JB7loepzt/vP5Npq99MtI/maW1
Yd+34aYwGEKO3poy7csbsi3yUy/NkJ59kc1dHxcbfwl7jTzs8VnDgnv0pJO9XB/HCBJ5xJy4tibX
d9e3hw06m1C4gqGWz2JurpOBj41Zf5S+IjGKeNyqp4AMyUhW7OaWt3PbFa0RtXyt31+tm0IUd3Xz
v70e3Tu2jgz0B6NCymcjpvmt/i0saQbQPc8TjI9QrYnawsUIqhISMazlZoccWzh+VTqr+nHYfyPB
lBlpHB+eIPcmdh2GgS0DO3DgaxiCIqb2Gvq7kKvqE1M563VKGzzoEr6zJc2DLomnR0B1AhRaU/s8
zc7ZiG/vXk0ZIdbgdbXbmvttA18yk1XNC60iTPsCmUMX/PG8WUhzJl84S1SW4hsVj/8PsPCYAeNS
0ameyrCPzOaDhibWFqukxT+J8L9dmpCj5MNcAF3Jm0KzNLPOgylnN8or0bdZwiA3QLSRiGj6L5FX
dFXKbeKSsA9iO4e2cExVM7nYEkpXFeYoGumsn1EN8aN62JiQiG8UlHlSFUajDtH8GgE5nOCQOf1F
11Y4j4rmJk4RiJ4Ix7pe+0sWi8nSJ1ByXqC4ugoThSAZUXPKQV64XjSH8b324abkhbF75qEVS+2p
o28cEJyRI1P3F7+hkxfyHH6WH1CwC/B9E4mLI2x4KarNYdi0KdblmK5t6J/pzJDqA4HeWlDLNV8G
cSsu4Og5p/NMawzH8Ke6o6e2xdq0QpZt9lbh0I5r5ykWITbVBfeFOFiYjWNmZ2Nxsouyr1DmtVv4
wLfEC3o1MIjutUJyAS2T+2EnjcCGfddEKozs2brG02tHlVr860TDWtiubN/XvYrxPStNbUZbTEOs
FLkRenVVfWddMoS4ZXbDKheXIC4XoWQRjzdtQ/XqbF5rfZRpbL3z2fGu2rTpQaKHG2bPRWFlX9tf
nmQFq1XsFmIY/JUJymN2ZpiEMMw0FbRrUwag+eDmXkuWWY/tOphFSDRddfSsjnPgTlWw3P+yHqS9
4eJOSFK8n4pMNg8iB499oF+yFDuAkDW6PyuGN+Gfbm3OdTO4qRsYmv2AHDYT3dAoRJy5q87BkS86
7mxOgblFgB8/8oFlQ8/TUgR5AVAdFhrTiH6moD0rq9LHxznvCb0cH5hDzuDoVGbAGFrOJUtaEgxc
myNJNzgAEZTT3plrN7ilk7RfGo8ggxxU/DFB+Dn7N+Q9WbXMinZhw+DeEChXsveb8WuUCrpAEObL
LLX7YUso6lvwIM7K+Bvv3kkksqAH1VL/5Zj5HuKMFej63fUyLgrZwb+jA9JUZ4CIgQP4NFdRW9kI
sbN9ZsYI6+b/PtWtzqIvPm1LdWLCaYHO/WShQRUJuv9R/KeTZqNORhRFsDU6SmQ0Xp7S4NPDyDdR
tnC9S+dBAtbjCvMVcry2GyPTE6ZYE8OhQMO+ZI9GCZVV522pf31lABPFAodVi9/K/T5S1gosfdY9
5hY9opvaJrlcgZAQw0NjITpttaGugpnl9jp56xz6cts9NmN0e3w+dh080Yu8qrnsmSEKjNU0Vi7d
U0aDlLVpHcwUnqgAtNnnueIUBiywM3+piKJRxGyx7eICIxBnZUDCk6g8rkuOzGcvK8BVxabNZUfv
eNjpcrasphDjvNvixP5FECG6sBSr9m03T7+nmnmSnt2LBgNdNKulnhfmbfUMpIO4R0ch1Pkqpzsi
CdA7C99dNkzJr7s76manuE8LMmuaN+sar5dP2rK18UhS3dTO/3s04sabHnAz9fVxzIhNhT96jCrY
wWGd6T6XXqY69POVkZgqLhdIs3N9NfCr3kJ/hgfVPEpZeH+xFMevoIqpK6OWWMGPcAj6VvWL27vL
k58+Kkfi+RVoYRDcCwbUeaqGpYKRCJ1Og2cKNo8pgz0Nd3Fy6xXNkRqBLGYqTZM//Wjm8tgH6Zi3
fTlkw39FjmlrqPkoeYk+X1i30MWe5oeH7XRhh5dD6Gx9xVysnMeoqYC594BlvQs2fn8ULEfVYGDy
QUx/OCgN7D8/JW/Djp3SpPOff63+Gq05D8HVPimVumkvFNk9mVOXdGJiZfnmC63TgX1gYIf85IJY
zmlOfHzJgdUr8FlMdd8aGfqhUUTafHMu1o4t8Xg906KQecf8dGm4jYPXwnjBgOlZBveg2zVEZUb/
Bc0fJ9qJeE8kvezyhfYcGA7/hSd7E/uehVNs1MO2OvmmbdJMF8/Vb7BsHkMnAoFmyBy/+/9LgrB3
+dXu4DstScog4+jSGmxgl8oJZtKM8s0iR7ODntR9Yb1QHUOe5T5G5EP8UslQn63L2HGxGlv/pjHg
VgByE+9/5veCvdmwVOpJURrQom6EN20AYJXYxTAXOWbqO0NcIOX3ZvYEGf4OLmCuQwOzyiAEp+Q3
ib2voDbi/wgxPowGD0M2LZNFkEaXylpgNfmlWNaYg3mlrYD3s2wzKUaIysaWZsi3r0Ud/z2SxGQ+
Y5e8pgvWaHsdpHmUgvIsSjbuCeSiVOsCSMVZfEuTiakwS9cO+j2WV6kTqe1EN+NphV4Lph0Yc+4e
x2FmFDidgjxkG2p6rr1m5EuFalKix9NVMJnc91bI4rm2ycWc5VE5F5bjCNzIa3VJ7D9UFBSnJ9DZ
ULJVEyHKOCmMg6nyvgVGcWfAk5cOGsV/bWcYKqS1cXWAHwwB3jatoN7BsbVPG1zS78ttjGe17cgu
TxiffL4q2RkIFI9EJH75JikMecnQXgtExu+C2drMa8ljq5fWt4mG1wJq/YmTA/SQUn7NHYBvyUhH
oLJ+d+n5Wptxu798r1XWPfqrhEK0CS+1BPGMkhl1ROB/WK6u8oVo23pY568vsxKtjZcQdv6egooJ
8o++RfdsGSJoCRFl3rqbb9NNz8UjEfzzMFRAPRGNOeQnFronsz4Na+rQWr/AKN2IWqxjwWBOXltO
Q8Gy38rvh+PQiV+xOpNmwTBzV7eTKjfKV8h7LVsI3uD21/hG24+9my8jxEJg4qX7wGV3oZ0V8ACA
aN5UKuove8NBKTugKGVAg/Yyoe8pzZwCuFzvdO1aSgko+iYZUMaifotxqkisoMaslb3MnkSM56GJ
X/qpDVnVIg/i9yhLgHF0250PJu/6s9DOrq9Sq1i+Ogb+8nmd6AOd5LnrOK6ENI7xkpV2dJWjm3U1
eJED1aYjMm1WSHFWi/dnN0pmlhogI11ddCs/GpBi+QSE3gsRXqZxeo9e2/H5xHTxNCuODTqxcvfb
4lXJ/4C3Avcs+RRMYj1ypG1awXcRv+j26tFmjGJyMgRH1JIC7pGg4TVvYCTEE+e2+sKZamNi3tka
1AMa33OGnfFzR+HDT74D4UhdJQVJ2q68/QyW4hL2nW2UfSa38J5QXofy6lkw4KDWcpyOZ5y5tgBW
wU0pXGNJcJwoGxZacTNv5mP26TJPKXDJ0lOOzi/sBSSxN4ePT9jPfEBqZHOXobIYOzGKnycx8SOX
W3uArgbeL6WDfu5/rOgZDZOVlk2RguIDwsCKFqOnul0oIUXyLSBAYLGDJShGszNxt5iSeHVvTyGl
TbAPO4yDxAZgBgsaOLQBuWMU7huuQL/AfHiqfN6cG5aGBXpIUUeCGR+NRTPtHHoxIZtEtx3uwSRd
F23esA0MKdqcZhktSQXzZRsYbgzJdUTFFfNbRryy9S8K7VXpucRHhJA8HXBT35FN+FFv5CHEqDu/
+9ghIvfQnwEDkeLIU7b3M/HfaF2sP9GoEM3d77PmOBgubFGco4F34CsSEAuq1nE3rOeJb4+mlfcW
hoIwF8i5Nk6+T1sZ5ltgpBm4tFB3l0HLtE2d39ecDyPJc1vOH5OxMpByf2stRf2LM14g37qsiJC0
WQWkBTFjb7FMJCVSthXXVFhsAIKh3gtElmnHe9+Fadw8uFvx/Cns7gtTCJcNmdDBedwNPpYn92MU
fLuOfcP5IxBcxVP40mYAcZusMDtSLedtjwNE4lkUlJfabRdKNm7JjmiDk8Q7T9YB1rNEh0dTeqJA
W/9+zK2einX/4LBp9KsfpF6cc1UDPV6VyqUT5TefUXOXrCoNbxSG+Y08lqnm7suMHTWKiGedTkO8
CCymsOsBgyM286ttgiqf3/230ZRrvnkNKhNgVbqzOnafT0SmN3XkLc6H7j6Wvy15nwbbSj35PvPN
qFw8SXI4eQrgWMTMsJpg1ZIizDc0dSIhL7L61fnNGtuvlZag1wg2qbP8f739IFp2c64JzNItUaiT
8tvDCSmN6mO1tkh0Ha6OwJxwVRRyYwFde5/fvcZoHHbopspmmTb5XBhRJEBuB1cFpcXcJuBs2r4W
rd1MNLry/u5S4NdwaC/0sho00cQTikO8x4aKJ47+ad6LeHKJsU+u6AGtXew2OmcHWVmg6yr0V37A
r+c2BvnDnDIdyj+5TukrqlRROXr7K+pTnw6uA3y0MESXKtRok1b8Hv6UDApAfctZ1P571JHsyMp3
DihzgKssoRuDouFz9Y6E8OhOl4ZcL04nK303+VV1s3RURD5M4LbvcwlBzwsUJKVU+nf4o831laB9
LWVHIkItYYJMx6Ro4TiCoap6p4NNr6OY+6uKcwUY3WGWJINNC83flBrR2s17nzeC6v9wUIN2FFRb
QtaZVaGFti5m35dDx11cHRrSucT21PWjJXHuBMkmZFy1vMs7bqgtDW4LuW5XKtf3fQkkV6al9uM5
p2h9ZYLdl2pih7dnEx8ydVUe6juXKzEYslNNrAaUK5173OCj8qhvETsKMTTpNvnhwFjA/yuEZtzY
hNKR2UWpl4cLd5rBnEUBVMwCcgHlHmur/jRUkqCYY5K6aqneHjV4jKzY+ECnva+fGEH6vGUzP0g8
VWFco4xNGp9mQSxBtwmZbL9bft7rBGVmWbZ7WIc6p8ulF/M1ToVv5epejGs8LD7A/ZRZID38DCsX
Ad/VBsuFMPKq8ICjoG13Pl+rYQyyYXmWAAM3eD8WIFQn2V//EIgzSq+hWfheVQCFD079EG1nXSgB
kGOrFEw4t1c+UW6GSCdYzQskBhBjtsktnNRpfDLwpL+uIhJmwcq1QpKmz2hdxaGmybhKRYjw5GN8
XxivnJCwrkzZJ6iITVld4QSnYHejtcqGlNoZK2pNSJ7YAY9bn5px/o/2MR+tQrNs19l18mTCYEze
hToSDXNIcLdiheC/HYjPHv9OuKoVFZs1DrhxPdekh39TxIjeOxN9saLIpmFfsKo+TrBmSvPOw2cq
t4zgBpE2VAHpu1fbDjsfO23sPGSEeE2polqNhP8h2Aj7bAa0Z26j3nVq0w6xpFlIa6AWLiuwQYPz
1WrqGRPfosf+R+kD/eW66xUXcLjSeYUNLQBxdSqIyQR6IozG6na0otq67YgFZm9iKUZLZld5ONkQ
DC6RfLiMoXuh6ySFIis9gE+E5ImPjLXoKmqNhO2bCbYMOxeK8brx/ib5iVHoxpXOEzXiJm24H3Jo
5YcSengENl3QfIP+kLHeES0Suy0W1rI9g+XKfsM/p7l64mq7XiT2jbHnNcZmbVX4JZgFJUJhS5Tg
KxMdciGyeg3lw2ytHC32KhqqInPApf0sWIgS2BUdFlUZnrciNj3FcjiECLNyDQ8nSsDmv6p1JRs5
iPlJ/E0c7tt0xqbucyFxpbqWs6jFOO9octH7ZIK0F2LQoQz9dLwq6rXwDuI54G8YSZ7A/+JdkQmR
HhEyWCNCfHk6sy7m6P1R6Kyst+hGhCb8nxVOZDmKneeV1Ji93ciAdz7WqjY5lZ6Ig5d+OGXqC9JW
SKH4HULNDWlQ1QPktJPnVK0rqar7CEYrYaw8GNJWzKgXRtIVUBhANrus6BavPdg20EJPWTgl87gU
m27ICx4RFoOVeneorLGFyisPVEO/KsgY/fme93nkA6e9Aj57PCEWnBc/zUxbxUq5ywrwRQWMKFpj
XQf4rxHjzo5/+CVNujfJchFjsGwMZO8bbcsi8ycj9Kv4wcQC3ZJUfipYGLt7y02Zau1BAWDlWQwu
CbJC13r+TAfdDVsoqyNgYMmDH+1HTF4XE3GCYmr1BK0XbI95No/Rfozpz91toeeSBeFizVnxjaSM
mQkkQjK24+/ISNoAvJTGQdpYclLZU7BDndHOHwAZqoNTC/ILkpnzBTI0sP7RUn2KxZch2jEyJ0sN
m4MOgC7gnNMza1jIR2NXp4fO3nNwGntwNGUuHauUAU89kjRQnI3J75fE7i2UnSwkDHB8kd5zGhSF
y8fZJPr9inz/I1Gvv7RX3AlsrsDoG+TcCjFiZGdAdguu37NcNC18dRJ2mu0D7R+cpfOYgw72P9lM
T3rRuz83ONus3fOev2/AvDYXFEbE/iRtT+lhq13VRWB5AqEwOeYdpQgmYDTl0xr8IzOwK7n5R0QW
x9Ww78DEih3Rgq647ATAqyGeSCyPb/IAIcwuei8udYKp0Qezbg0xozu/iW8V72Zeiwn/8weceirx
S/H33980oV7sRb7QIrnBvnzTzBbky57cB52Uz/P9Uzf6I9M0yGr96b4PLSjAiIlBXgnX8ItVSBlf
r3E/3TstkAyV5OBwVP8NgjCnT/eCCRz7IjHKFpQWsF64aDoMTeVnC9EwZF9zuo4PK0mM8Y9TmRnE
JR0JAgcwY7Nq6ZsLtKyANsuFFaYFT+f3Sj3OpGVCILf+isYI9fe3Ys8MYV6CNJdDoCJ5IHwc8cJH
3ML8SACTH7DMwJrY931FOUR27nyvPifoY1BGb1wNQzgvC/pHssQ02ZdfpLFTMoPgRF+UbAiZWTRP
pDczc7W+r2+73+w7w+Fyiubqf24eAzSd9C8zs0EkYRwUI/60pxGKzGlfcNSG8PnZnyiq6h4Envof
NRLhvAgulRkAjC7F2O63FDDtux8QxHLMmOfuVymVAzRDw6vZbNQ+BtkcXWZhN0K2PN8/zUFxNCo/
iCYU7jw2j4Wjenw/9h8HA5USNKT4jnsbkEWgUIEGkcMO2c5zfllZrdJvokg1O70rfPZYLV0OZGfo
r++aEBmVwZyKc7AGmQxb94TalPY729eXqikotwAfax+ljVBPApXTwHx6d7/kIVOd/aOInzNds9qd
DAmpXpcJqDnFeMZBPlu7ZJLLfqZaqB9FupDzciUERz7zA0qntHFmwks84iBwWkleInhh/cx3Ocj8
Q8mtdBjqJGyhIUE2x+wvVr2ptvkpJe1yLggLw+MxpzJAk7+a466hJX9LnzD+YaeBvodeAvsrtfWs
6C1+OmS6VqnTcjP/e38KU0F10q55zZ+8J+9SiyqUUDhDojoAwqPSOWxhXm6AI8eUAIUc0cULQIKg
/6LOri2WEnBh9114mjP0nKwCcNmcU3Xe1u5mWKaHkN7EABWiDATUBwHiZiJ2npxj3nj/SqjAHHRa
ompDG67DOsD4jMC1fWcz3j0hTUGWVIzi8HZkTahMcdqZYmPscVmWazrUZyElS4LtdouAD5SDqiom
1MtsbpnKnfq5/2/WUbDygJuWHeHCmJbjsmXAK8zjrHp4VDvzNsgowhwtkkO+rxjmavA7AT6uAL+3
3PWZVZXG2MtcDAQpYapE+8g0Dfe7iiZ0/i9h+26hYbcSIr0zOv+dCNzEFKwgxnbBGgm7EXzD0XIv
j0mrwfsggthsDbGNPH+kljdJqwgh/RpcU39GORXRo6Ubl6un12oujtPFXNprjVge0IKj5hgrL32C
bREbIRnlMoL5rO4NH/kqi7bLLFeySyDnlz2obyvRS0pq4teuaNj7EpmoWTvylRcbHHNyQUfwcogM
Ey3iiVQiSrLZmMKb8DCDE/DORUP9DupCNbxQyGkA9w6mC6bDY/bFC4eiF8kqTYfLI/9wgJ5FZ8ve
BJ2Wt/TZeOJIabaIiR6CWckyLmu8MVRFpLMqdxzVLs8NqSEvihkfp7c6sry1V1AAhBJTC5dyyUq2
k9L9M3TXWX+G4WUeOukGO2x+FVoAdE3UX+iXbncYqYX3zCRlXKlXmIf6KbE7KXu4YNidzI41GABH
bbj90b46ctIkw3mnDq9mxd5jkVnlsyCRyV7ZmzNSE2dUkzZi5IpQmUA7uAcp5Rw0fa3MoEFYsVl0
b585m+uReQwC0U3sb37qxN/Dq8syiYdR+IxNinlfPJh3ic3CLr44SUbNbp8AhT60qNgkYVKOLRtP
VQw4QtfTiFn06RVEhwGuq3tXnh92odyPHgcDqjLAQg16zVrpX24yTYkafgVNRBOy894F65N3yls/
Iu+e3bsCVCo26X5VdAO2imZv0pRtw/y6mUiOoktca2DUxIq0DXyPThsjH3Mg6Huf9lBwaJnrCdD+
e1cQsX/dTChFz0PuLjYP0Q0ckCUMr3sbZi4rM36KWq8225T7wgPK9k2SuicYdHIJW21V36RNOod3
8gax6n6A82/DkHnY+ZD8xZyvFp0Rc5gCDqcXJ3BC/mfbYDOeEXu7+jMEe9FGCA6Gn4tn2mpRodZ0
WJjBLTAlB/SbB+7M0I+PK0FpzbbxSgA+5CNNdp8YwuCLCzd+GDYp7b8mHmO1d/PRY6uNDcumLAVL
m54yYF3t0iSzhR6Syz0pb4uuKcy0TKhDFD7jkLkixybff3ZnUVSJEUZj0UCf05EjD4i4ybev5QUQ
SGDx8xCHWJhYCYMe9kluAbiQftOATdHz2vOgsPRDTPP7AKCeSuOIcBB3MLgfQhzPMLOBwPviM17s
S9pPOL83PPif3330sJzwGmybS2jeFJUdHon24beBwYon3fhB5a0V5/exSuvtO+O5vwuO5bqDOGCl
h5pigfRZ1+m30CwZv88uJDsq04svqLZSOn+AgwXI/BumQFzf5GjP4appy8xJv6O59PuXUhuG1qYY
3FzFv7Yx+Tb9/ei5y+cMjlS1yAQ30rgbwb19M2B5JZsHS+CcL4/bZaotZeICGraOmRzmiL8m/F2M
7I7iMhVyom3t903u934QbNFYxTzvDztGWCjVpe+lTaDVTRBotzwAEqMtV3u5pJFGpT78d56svD2q
Lyi3UJay5rhqh2+76BGGtDPzzRDjf7gdqbkJSSharh9AX7NwSBlqTTgX0toEzrnuYUJAl+htFPG4
3mymfkwUs+5mXAueD+JhH09UFkeb5onloaYNME9/882lzr1Omv93Nvh8OGc7H5ehrR8ytM+ORX8H
iyyb8aeNINj3xmMu5GstRVnlcTo1pmYRnCQFTayYcgOi6Es7l6MlkP/nLFzvvDW35JwrtPzLruJG
xQHmyjg5lK1CCcblujoj/ZhUp+QWAqBO0wYWyloGXwEHLlW/9TPhesyXUv5CIqo/upBvOCeO8fpT
XUdsxjaMWgP1MPhNZNXhtNpole+5JWwCsIeFizeNclZ7qbCpA1URuNacMKAdvVDUdmbvbO1+ARxQ
jR9H9WstOsghCMOuPacqrhASNJ1KGGaVhX0LhfPMGhHnpduJv8SYdBIOGBlCjwnvIiFQcjLM2+ud
41KdfJiLq3l/SMKD4c+l/BdhCLvdcNEpM9ShGyzfnXZseBURo/+qdkEdMAHVWITMSONyRMr1nafG
/8eKANWgZCwbkxWRr5zKqVl0DIRvpg78lRC5FKUxIhHN87NefogA4fxHgEXNjmPorhoRcsE8UM5M
5wn3WfGe0wYT3YC403Ku8KGddVCx/Y6gvJQJUCbc+SzhYCk5DoIQvEBjlhPxwwNs0nnFjU2oN92q
U5nuDGQFHs9M9rzlyRO+P5I1O48S//5GxruT+u1J4eEMj2s8fq+HZRllmPAnKmrFyex401x51ERP
Gc3eweIM196LebdfGV/riRVNlXQ04ZpvDQ9cwGAPYjofsZq99WwJLGpgn8isoNn3cupmGjWXuoCL
YO6rXdNSNutMyCsjtP4nQR+5SlTHSLK0+O6N2uhnpBLU/4RCnul/5Jo8XjBU6FMmUHEHTY316Odj
hZZNUCEAEXZe5Ut2/ZUDQiJt4nIVKkagUVvICEhed95AfEg8rE8cDhQBYHCbAZz4qzCLxYiRapFc
+tbSazT88oS3azccbZLG4Xt2e0y098H82XZvkl72IHDiFiW14tAj4zZ4ORmUAd8kcQeSZeEVb7Sa
EYq2UvVYHDu1BFKccnh+4pe6pghZthaOkSAW2o86cwvu6KQz7IpWSN0mieWAuVMdLPXIuCMSaL3l
aXQi7uCgXVz40j+/737bYPkV7eLpP+rAwSUjmMapSlewfmiskrvsJN3DFUHHr0Mh2ic53QGZzGMU
yUWjgIlK+EHeepXFT3bOPNN9O9XMjDSLQ8b+raU9e2abnIrG7rXDiaQibpN75ozd9EPcwOlXyZMd
/H9YVB7I0PzKk7WqCerHWL/DYfSTfGVhb+z5ckVoO7A7jyiTcCkdHezBnIeAOr/2pkLxZ1Hl2aV3
V5UldX68pyitbEUJH5lILrpVGRGb8UsxbMmunWgF7dul1DqhMv/uTzjeyTx7Vlg2VMZhIZmizgP9
/9Dvg/sZmMRuVsiwfsie/Hrxx+L3M0ttQtK99GTJwHkSWsVYO6FM0jWz4LIdsLnR3IXEZmXjv3rO
7F8E/RHU1lfhlTmehhYBu3EruriYWJIgqREn0dfZg15lQcJb/ZuDfXGaDs0y2NYEI251TXSGpT61
67pYDOxBw90p+BcmyAMizGtd9zqpmSCIkuDc/R1cNtWWFK1+HbYxPqsQI1+CyHI052mU+btZuhi/
QoU1DYKJkMQqReKEMe/Gfa6XX92ifj0KJvXBzJDQMEHBFFnt3o+J0uzYijrp6jf5KnmM7IJgaZk+
/ab9Jdlrz7kV+XGTB4Vv9qB/XHdhlKVqEUKAyD1mIdhU6nZoK0YzSWJ+fl8pNO8+/6buJM52BIG0
DG6gHAGdSRGpuNwJYEPqmEUcEHVR9PsSI2QM7gwc133jD4mN7jjx12RSBA/kZqxRVpdgApmq9bDh
E9jgyF6aqxlEoFIMaLB/7NtRKcacZ9cBI9kgebOV0f1+pEtY1GrNkV75rhMR2sZTUaIGvFzKwojn
kb1Dfh5aF6kzoqy9+Mx6Rh15SObcNRTAWLcXCrCKvkw5bIbqOU5obAwLNyd1T9hDAwIykVyHGd89
7P+jN4Km9i5ANnlV5nTsTZ5DFWgQ63H0pRU8OA7NUgOxinQTOVBRs1uI1hUqGADjUqXKevk7x7Ma
cz2ufGbkt07XD+PUV1QpZE1YWRfW9mYW9CGBw2O27RJaxaGRGji/8EE+pG3XI+t+T0/4wWDMs82K
kRax3y6CVqnc58LQOHu7H+gLM6wTRAVg0TQ0gn/5jiE9zg4RcgeoqoEzyije1HS+4bH8cHF+FcKg
zE0b7PrTEjP+oHWFqN18cpKBGttFvQV7eT11b9pYJxb4ki6SKQJUYjS4RSMKtm42dQvVYknHVTYE
TgSzeNBKCpNB2PFcTwXB1vSmUT6x2+GXqrtIQ+FgSlT8xaqnGUPkz9wUuE6VFcuiLw/4LoVRSNfP
p17vBtVwyMV3yqVinAGcORSkGCkxhS0AxUdjPj/ROiwnat+lw1vHL6kVRt+6ck8uPjYcVZf5ZhdY
jdPDW3tMrTtOwsL/pRe/0c+/wzEFe2FRCaKSSlPsT348Qxr28B+Q2dz6+b81VwADUxfUncJPq5t2
vkOPXkL1cSoevZBZ7S7PDEYa9lO8R175w4HRQHXfq1mfZzTL8K274+MACn21hwOsZuCJyFSobIMh
goWYHRVXzPA2P1jG1w5HaH7RfNhw9HcJpYSguq2YSTM2NvyyqwEoANjuxFFk35xXgKfJHr8FH17p
G1tYRSEeTPt3cFmFGrssALR//mx7TW9yqlK0iTVQbQQ10Qkn86ufVnS645xyVxX0ypxxAuX4DDhw
WDWHE+ZWxFl4bCr26ryQQlmidCTr125Ix3AdajQAyZ77wugUYBL8MLtl7rzrBS5gr7F/zj8lfB7H
Zs49IVIbxOv2QaSRHqNsNqXgz/P67LvQzFRCKPMjp0E5uUkdqx/LFOiVkrJ9D0zb4dEmcS0VFI54
Fu91ofAbhcau4sBJM/+lscVRh64NZ/CvVYtX2Olo6oojlu4StzOX2mwkIJgcdhrP+K1L2+8mZdg1
L/wzN6l4SDhvBURaqLE+6qWAIblmj/2RPzpcVVcmpctIRdVURIITRHAWBwl2ATkKeNAhSgxQGgjd
708m8QCUsVI57itu1LxG+uot+pMBd2JglkBTxAlc3pQ2F/jsFyvwrop1TcOV7sVSFTjYoDVKDgfe
0A2IK2Z780FNdcU4sZzOSym6bz/Htc6wjTIQgsrVAmX9Fx3UIORv3gahOYKf1p3Th5GjN0OzPVIW
CDgMKKJZVNYbshT6rmBo7IispY+Ww0N8MtutKqygIlgdZcUlnxFOFWLWmjdoAOMsaghjDwh8GRG6
jg/oJTN1ju4HQCpS/XVq37MFz2hcmhi6SyhA0uwm8Yfr0CA+xiDepcoBsp0rnbnBYqxzV7TlsJV4
XhToQzPe6liwIs/qIrjS19xGd+tm+1AdJqC0Djkc1uAO5OMoBhVbc3nqx7sJupVDfYhGWTCW/U1t
8kIN3C4ob6KXdj3MN7Qm37qPcyOGo5FeDTR1ZiSAc5U1f21tCkwU38WXHmtj9AmP0Fxn5BhrOZXy
H5gAfNDF+NUV9jn5y8kI09itWIJ2TRelEQzSbmJoEwWrbUI3r8jfrh2iLscS7KkettBuF9Pat+qT
q9hNZDnLzqNpcfcpGd9H6pHtS8tNunj0O2bL0VG7BQOxaN6NkbGnwCKAr80WRLK+2H4G2MMtfm0w
gDX5qr2V90koJDYOT0A096FH8zV5Y29kGF4XjWWkYvu21piZmTWPLEx0v5IJqxdKfQ81k+PgZLPg
vltgK5m7ixexBMn4nVzpNvW1Og8DycYprZ6vIjmy9A/U2BNIQL9DSLIZNQmMVcuX8KpSfvXAdvZP
tTHRq2r7cGPQ8pOeo56Uh/Ca/Wuash5WrAtNqSWE0xi7pJ4BHasP1aoERBr/s9WajZBxz4CxVvVd
r9K0yVkNrxHCq5kWMS8vl1xiFUW4rjtiuRByjXLCfyT4H7RTYceiYDpjbJMTu4re2P+QtUYXtYNh
G8KC/eUhho8msZDialDZJN1PBAnS9lSttAt0e9ZdmwkSdCqkljehyVMwic+lsxPk3Nb+g+Rdgp1R
aK510BNfNq3OABFVn3wYUjrEB14smpESdk1/ng4XjlQsUYeYbvUZKuX2hI6yrqwXBpyXaRclP/BP
qGMI0ahFBqAkXzWv3OJNnGWxPTAn+uQNs2VHqSO3f4dAng+NBhMtH46hdigTiK5gD7nJh9AT6CvH
arxhaRxNXWCQnUWpPe65f5Tm94GDUkk0apQL3c8k0kKmeywjmO5bd1osmeWtcs+TWKM8qIg2dfGn
1uzAzXxhbDqiW9NJUU7Et3lR0VzeW395N/uDRQf2lgTcy9H73LTPLYcV7qrzu2lDAaQvlnIbx2J/
cCdsDhs0pypvhDFJo4S3MtNRp5hWnX/5N/+UZi8csL26PtA5tq8mLQCqDWY9rUoOkpazey+gxu5a
+rlWjZDwmN/pWQ314yQJfUyRJwqC9MWpsgV9cLahovWqgwZO8snLL/D1EpqjRo2h1iRilNaK+Cni
eT+mxpM9N3YzFp+zmhTlL/dbRWS+Jrmhq/SfrbIVSgNOHzi8Il20MBlDa036CfXnSXXYNKq+iv7i
0GcjUo8+kSGI58uJeC8yjSyt+0amREvlpvnvUn9oIDS2SwD9gfMXbBF7BSGuQYxO1TVtXL0GRqV/
uWHPeTLkl9J2w+/mGQXVrwYyv/RqTLfHXe43NZKj55xFamTgmiiyq1yUnCPqdhI9oo29Hd0Vv8zm
Jt5jMksS17j2b2zgSU18H4GjOFSfS0J8NhqCsltbhHC6FCgo14IevlsGuaYnLwk4r2qr5WqKb7pH
JBgLdkibRT+JFOaHAcijmJTTWLAlUm/sj+4fnnLjc/73PWsy+q2Ddu+KruzG91aKqNanf9OjMADT
1EX0g5clEI0NZaTj2KIVsGmQHjIFGIVh1ldOt+1drHggf4KETHZ5xoF/7S9LsH//4gaLsJxcv0zZ
vdNBCOTjKZWKukhYe6A+zV6gwzerVg/4g3P+xFPcw55Doy+4lY1MS7V1IBvhNGJS7UHiLVaoJ+qa
oZisf83Ja8yQS/WVunIn7/7oS4O3VV4fsE9XXclEl6cTlrWK24liJbxWQFokGfx87C/MlOGi+fPN
RI+KZG0O/AgQ+SzFFgQ36f8jxXSGvwgj8qGeWiR+sO6tTKuRK4lL9w0QeeuwOfHIzfPq9buvwM3F
nfAUMEjSUhARuUIrWnw+KDkGjYOd+EMx5rBPWwh9LE2N4vchDfxt3cALqkPoIs3XbOKz879EN+cn
EHQ4rby78fLSCxPLcMdbnNtthDVIYhV6uaRXhmunIY25SdIN6VyROX++W/JRo0lXE3U1h9cgGpOo
oPVedURe/kfJOpjCSHI1aJfTjhrilFtz7rYpJyqyIsn8RWmJFVaBiKRLXDLIiW1TM08ENWP7lmr6
0ryRUzmT/KLajmyVhFYEZxqjfPPwf17UGjwDIrs5Ef6E0W2dvU3pMUtxPUq1HiWZwaLWTHnw3aD6
dkP/soEiOU0ePROgPIZrPvyn44+YfZvb4aJPD1eGIYvhSusWfuBBCx4M2fsUrNFLTi0rg2AfPIdr
+BJbvMn6+C85uT5P/2VYr9TJ/06ylJb/pCwc9YDLft3PiXSiJKhqzlik5hoF87DH9korqDUI4Rep
DmbLOjilzK8k1sdx1w2bSknL2GDhwTW+Ih7jb6udEnF8uGce8kfKgmXhKYFoRq2+VV0GlD+lyGNF
4PF+NRiX0f088IPKoko6XNkAdBk5vp+xBYQJnnaP/WbJnbTI4oo80V7suTC+Mpxuxle2+HOppMKd
YVD33hNha+Wwy9uA6l8GfnPY0KYGeZMpQK3VsTagSrLGnFTO9wLSUia54JOFcHmoYzWJDPPM/V+M
Z0mI3TfKPMMf4nAcZgaj7YhTbcOZPv0f8cL/eLo8tNNgaP1/jlkKUN7PN6+kCJOvHIDbowAF6KrP
1C+THnAAt9V3ObXSHJgs6w14urlG+Jfi7I4EXLLHGU/71XffArwMGa2u+zvqWomY85Dw0iDzXiOG
QBPZrdVLZCueb7JOZRHDamDsQQmYnEsSYi5XGxYIqroz4yD3JSzDPSByoWHRjgf9uJUVUXrXI2IM
BdSX/R33uQMj5CI+fFc4vhlm2R8eMMM1Qtgs5rdeWntI1+PnPI2SjRYFPvlShDewuDRdeVHguzWJ
KtYfvX7r2jpTPDYXhflL5JsUuqMlh8eioj05BIFThMqxAmh5Z0SRjjHZP6KmSkxXFgutYBjMj4cg
6RdTIKaykf364pwY8ztWNlPgOToA50Df4U8vgc0XqJEfVyVxTJvuOf5npM4A0YlkE64LW5VRUY0B
wv6mqyn3XAW//Z1h3EOA6DtYr70br/oentd0ThVqt8fKSWo0y0JksnULR6sM/Dva1AgcAcJRWIAX
BAzVjHkgZ4dIrkySs9S47ijkCIohV4HdUwQFxpYSjDzVA6CJIVUWftMYMjrsjBz6ukmQpOtC6Gjh
58I0x0kg4fWOB5F7l6E3zpb9T7i1ZKZlMvFJ7a6Ofme6OBxMcNsO6muP95Cah3zqkeYw0jTD/RwY
tUf/Pg3gWalI8R9UcV+g2VeG1vkEXJDlK6UdVWSKNGJ/37UP3JulmW5dZSLKta8EggOeaHaQxchT
7uFeW79ODi53+QVgCJ99Pl3OpZI5uPwUM246iVc4HOXyh2DCcSYiLNaE9wKhNrTJ+6wjomqnw14c
HM2A8cULYwFHXZ9LHIsoyIrWtXRNWC1F07xGsLE9CMB9ixaQ3iJvzn8a4ksJxMgd/T+fQckHg3IW
GBBrIGb1ol/lZ5AzgmQ53tiDeiugzyoQPQ1mpWCstGaPC55QShPvMv5VO2P3Tzh+iSO9M0k6bv/e
IpO3Os4RBBZAfsXgOZwwanD6OAKKM/GeZgHFba72g0+DyIzKBilA8NvNJ0a5r2aDoiNoJ6nmLsxo
c8+vtwxz5qz7smEs6k3fheNB0ltQjgAtlAFr0FVIJ8cy9896GUsdAVKG9dWblcLRaDAis1sgW8LL
g4vCrhbT2mtCa4FGtjkJ6nDtREn0hFSaa/tG1m9qEtTk2eCHCf+b7fQX+fLZkWOz9ckP05CROX9c
6t8IksZXnzn6BqVpO+GHyd2FrCcX533lw6+mAMdV2CDOZUIiEM9a2n3AKfNXfePCmOo3+T6p1LhR
b3D6hPDvQd4lsL84BPXnFJHAaHJ1PKKz8vGVLW48jRZTvQZhuzF6yfap/Sk/UFN+sF3jX/1PdKdq
N3IlV4vTSzZC1brnAYCtLTVchmY10QJn1opqOtt7+LcxrySqGme2ONvE2E724S3RcRozdsPZHaWz
MO++t6nKmjBcWR6naKrtiY2bCK4mSozaX6phS2EMBUJzQiIa4LZoxKfjcLVggzHG0XnoRCQO9Ez7
OeWV4GnDzavni2SF1WZHqh2m1kVzX0GDYR/WX/CbYOMuEJ0AHEPR7nEDMNj1fwvPQMArAcPhUhUI
r6kc483mTvc89v1cFWgwZTzEXsOAROMfh3vIdvouyxD9VDpDXNMAUkOmYQGDdKGL+YbiB5XP31AU
O3aaNipUxOz2PHE4UHp4SR2lMYtbjlG3gerklNNjrnSDqAxzFXWEheljV/5OjgPMBhMZ88mpDxHC
4vcou6zdhPel5xDAolLb1Cu52rumsBl+EQK7EroA55q8jiCKItT6DVZQqVWKMhvJ6oaqeQvuvDlP
M1pczYF5r0WjThx5KrA7bU/srn424xT+93RwnHjFNH/LMg31gDzZcrSMwWK+xN5LWnBPOGj1m0nP
VG03IW/gXF3JojXoLgbfWQeplx1OzXk9VsEpxRSqJbdzVPiKcLr2W45hYN70zdXyjsVlxUjnR78O
4U/7vCGV91A/c+2FsW+mYSHSLS8v+6yjfL3cPk7zaPflrjkzuzAEAaCNNqCqswO2rKFLWJiWglPr
jGa9o7ygmglYky+y+q1cD953RjekxFcrPqXsLa2VkZPJ80D7YQm2ooLktdEK2/4Ya/kXwcABov6G
kXabC2U2qMQFGcFA8MiRlRz2Q3yqNJt67Omv4UBwpVCipYrc15Lc3ZoNbYOZrBaDIqaKKGoHpPg1
xVS2V0DOk9gAwHNnZFJQA5wSfSozCH6dqzBE7qmfjP1z0MOz0ZcefKryAXC8HCf79Lhcp53Bx0TI
k+jhhFhA9SCkJnPHY06wiXQu3Zc8wzYm5vjFikqCr9d96+h6WqTWdlzNWouxmD6/LXkovH0nYABX
aqlzN7VbhTNgaPWqjk4nJhajMoqefJHlUqKEMBpfNSXcbPViQk7NineMYMPYr/19ysrIViLnncgg
XSi2LXExiKyhoQ4RPY4XJBz4AUY8KVxgs5DFyK7hVZY2txUw1wWUQGyie66wJENswFLx8SaQibfP
eSFDy7xNnwlMhmqwgdi3Fvk2zS6TasBtutI5xjRfn0SFs915AjIJMwmI9tFw55RN8gFtoAuxI5P3
IrITBXz2SoQj+WRpySRJFln55h1G4eSd31nEDVOBwF2sK4UumjOye3rjurLZOsQrIU37WVB0RwWU
BFPSJm84LAj6xwVDKyvgfsPb4P6P0mEjdham5a4QD/B11RqWy1e7fKWWPGarkmyTc/Bn2iefxtKm
fvhAvrowdsySizL8iQ6QW7ip081etft5Q4un1oKqZsqbw6V5Oi5IPDIyfr3FHHGwrf6Y+cS4eUGM
lUbaJpnP/LiN3j8Swn27acxdVyyvgEvqOk7GKks7LbJqOHaEI8amzfHTt2WuqVC7NjU+c8Hk3FpH
n3Tn+78XEu2wK4dfy0dAy0KB/FfJP27MB++x30ZjBCb7bnMsI1/b2c+G3gNf0qbKOqeEwxbfnAW+
EGxUDxZzAMP4xLf3BYMB/7yZx0FwSy/6ZKkPZRVgtnisTPrGgzcUnEo9QuZaItxFp/4D9fc6XlwZ
o063X6nPnbcPNv0FCJwAW34uKjBQ8TM6XX51waEdXxHp/y2u+kFoxVcNZ+bfdtgTXgXsv6f00k0h
kXvplIUm/iDe5hdoZvyztfqI9SGx1f86yQbTPLrNK+yrUTdToe6ju70S4jLTF2mP6S9hu4wbx1tG
oDlgMF1XXsWQPsVPlncFvwPuKNjRgDwc1b1rAixPM9imw8uiNbbZwSQM1OEUoYr+aPQ8memSWtNU
7iIAJ4cS5023OT1ShuHm2GdDXfef+BqNTw+8aQl5XlIkH0tvWuu8ZnPBGScLix4tbl7MsuDk1/G6
Yn17WasO8ddg3g9gELV0lL3c266UELprUyHp4hrO+2US7pi1RXaR78ZAe1+BbCl9Qc+2qHMUq8Cj
8TiHSVq11JjrqiVzb+oCWzGZvJEhtqvah+hrSv+3L5O+tWyyX+dizITvEUDdnkr8c4MZ8Lg4zrfj
PwYD2R55ujGwh40HK0a4O8Y7hBCIe6XXVQUEXoc79p05KQ80cDTjsxwBdYmgSZ9NcMAtxZgwxKDA
cjJeL1AWUkBhkO/3KW5zjGvSgto44vVfE4oOpcPipFgNynL4dicKvzbDFGUdPL5Pct6ZqzZY/ur6
jbqr+EPvIXjtgPjkF+bHpfXxz7yIYkDzwXXFwBdUbrO3TvPQdz2EmvFSw5N9YbfXeLQUKGmxSizK
F5j3oKWm4hBtUGNgx9QxOQe93Xec23fZPNeUiAdADHdkm+RVbbA9yDGxfx26cH60jVFMbrQUCabq
2t33zEobk/TBNW6PKH3eVkaDeboZXbmLt+KixHMkd7ABR+nYvKnAAJ7tEdhG41SZL+FRtjTKj0Sv
8cO6x5GXyaAzGDlUwmoWXyYmunMe/A7AEIlO0vgXOgNPpeGmy/DIA2kNvuHBRVsEiSlazOELuTri
fiKJ5V0O4N18iwJITEQdMimXoT0CK0G44jQAbCQ2n2nnYtX64bvSkFpuPGNKIEZ/rJE40tIkAKgV
Hzo2ySvBXH8SAOgXSI4BRqVCo/dDkPVk4zXpFL7Vx1fNsJ276ymRDs8dEwY+ZysNsNA5MeDNe4JE
mglqNuDo1TtEdzRZqI3L2doLXa1fVxl5ZvPz2K3miMbSIryrqEj04NdHww2iixpbsr9QvNndIxPS
URb/Sg6kBSPMVrXqZpe4HvOvldSYdbK1lGB9RjJAbNtsJLhH0xEAaBtkF78RNavEdtPJGF50yUgD
i0goKtty1UtZz15yogy5ysjPQQ8Zo0nDg24O8vtRj5FbZqIaSoLESru5loOX0aqtzjx4QuM1Teei
BvPJxXR6eSjJaaAj9z/i36y9UbGui25xJOxYXQ1JON4i+tlvPa2EKDTqHbvLYgu94MZAt2OjB7Aw
PkuAkSI78poUu4/uABA5ep5AX/elfduP0Djgfe/xOyG22hMSsXiMonG7Rt2jmxfIu7Ssj51tX/vQ
AHjLantJQYCAbeaPZp4YjttPEyk12w43MDY9AzA1N6lLg1Zjclide09fB3uoaOJlYKAcPr7rriev
+89a7PnQ0h91calbujezV7Larfa05sYbMHpHXzLOoLPO1NaN4aLO9MMTfulYPjKyEGtRipQignyw
n86+woXfzqr5JaMMne+eydntTObQkFSXxYXZilYEJJMJUkOJggH3OBq9/H6nYK2L2r01Bcejh3gM
kkCj//WEuJfYHrZvR7dUWv7qMtqyoJ8qicfLyC3WAINmfUNksvAZ84+VPyDoxxKvnXnDH9lXVhT1
ULsQ7033F22FpjjsVjtaq4ocih1IoM/qoxeAG3264GBlrDohWkKrh8WYfHImND4f7FmIH0kl9A17
7Vyi7e1cGsyVEq54WyZ3O1LPjP0IyB8m2/AiBVok2VXziYw39Ml2FuaPedwbg1gqYZK+RuT8Xr5w
hKsCmrJuKGq41e6Z4k0ui7TgYZEdgZdJ4I/Cl6kxhZvFLxxlIJdpAnHRomOSDDME4EVosLI1C0im
GBLuviJQOZUa/Ea+GmGxpGSLsvG7Bk45AVj2o5oZ8UoreLSRNyrzPMK81M12tU1jbjQ/eZsdtgi+
GNk7f7eBVIiHGcI/IAOt1+oMCMSIj4HL7SM/4cKhtgs0rKu3cS9MDNKxzoYdKv5aZIXlPue9yPtb
lgza8GPra+WfY6i8n6MVu4JXgsSjWVoHNNUY03020Jdh+3E2Mgn5qQ+Pll2bOVwBalUb4FhZZvdJ
YOY5Nj/nLCGu+LOb9RicDMO5ntSqU661LUohkkykeGpRz/qpJcmKEeDIfLB/Y+gipE73vczUioqd
CNckbO7GA/77ITpy7xXtg5KVn+X8HNzWPIHEaFcllfvUF4Hst/Xva7Bd0mBxlqPzlcBmQ0pnMYCL
4P2yXaLhkEyqb+pxNz4XXSv4Z+vlUQQQ4dQ4efIj7GF7WVL07Dg3qBpHP8Wn/VIJqNa33Ek84X6U
NQFKR0k1NVncmn7n4yTS9RoQS+ztc4xcylQI3TmBuN31U7a9JXCzrjF14UaaEKzJLF6uiwVPLmeM
KVdI4LucpTbEB1mTo2jPDqgtgsOI9Bxa2AOeS5juk30VJptPMLPF1GfawTjPHPAOWHJ8+p77PGIq
8Um2NhVHEUrzGGlPvXBh3aIgW+BxPfjYunI3J3Y/574MoEW3lWeDWaHDHiLDeK4UoDf38k0ZFOTU
pzG+4FSUd2PtLBpwbokOLKyrz+Uw1Xgxu2vLadMYMhYC7rvqkouhmH8aoDTQbOrdSZuXP+UAW6A1
o9r8+t3aX1jY+J6WfrajZzQD2plhtYe6469o2vOWzt2H6C8LEJdYVpuJzojNHlP8ZT7JwHmrPQXZ
uPhlVFZN6ZvO7b/bPNqa1quRh8BHyDc/xLXA8YnQsKqT7zQmnNOKnJZICj05CQxV2iiC3TOfFgxC
thK2rtgZlg0S4a5ceT8jD9AhAICXfRyI3IjdwX7KG8/XC+H7DcIc49PW1NjZ322/RmpTgB4X976r
LORKq5NCom8AarTCbhplgwc/tafME3w8B04eQyXSxMvcnr3FLCXGHMrVb3Hjj0kNGQ4cqMb0RTHJ
TZJoJTgHsprvA++zdmoV/rG3sDkRaQyA8Zs6Q2w7fhVJDeQUcReZ2ao/8KqeSY5VxdpW1kqONKaP
rpVRsTT6RU21/GbXRkrhxPyqggVTBvlhlyTqi9xEUkSQnnwfTOrnzIHc+ijvZqAZPZwfVMQBHnU5
qTDwUFvjfvs1Hj+PJ1//0sZzolWWi66gs16j+plylMZX8NkvAwDvHh/aleTk1j2V3gk3q7y6nnob
dEJ66tux4jcBOEhUwLa9NpifUgxibeGD/x167V0tx1LXeGG0VkAd51EmLmtAP+qxiwmvBUp4pwUn
wYlhCAC5js/YYN9IkvOdTl+MfSebO6pH1xypPdrPj+RJainMW05OsKa7ZuAWINQc8Aux2YZyE4LJ
2Ae99bULM/snPGiGONyhy7RZFv8fEko8yrXxdyweu5LSOrEVSTyEl/uKQNHLeWO3SreB8rYJsXaj
6jENAHXlAHwuCLwLSnuzdz4P7nzYmsosrRJwez2wG1eZBLKiUs1KzOB54Qyn5WkmXTFZkaTAi/T5
Ayv3jXo/X8QGB1auN5tEZFM7bCJEQ/g6mUCw7aROHjqTF/KU4042F7I6KqG0oH682fOnLb15PAZY
+5kgX8dzkEyXSszT490K2vI6P+EhO1R7cYpc8tV1tCcPyUolvxIFnRJb4mk/5nhH2LTnSw+Hiob1
vcKFBnyrUgfZ02smFAPsssXqPZ/heR4duWXi77uz9THGj5GAsz4io1OVqmh5KkIn/vXKsbBrqYlu
5DotCuDDeWPOfFUnzP81mbimwjIGVbkdTfVoVmquQQSHAC366X7/CjRget/rKTbOGSZL2HEFshKj
tpyro4OrR903wm0ap71jj73ErMwGB7pyH2E8C7ktIcXwlqaK0+0n9JnC7SDbqUQmCG9YQ3v2DXhB
IORoPpSADmbkPX1YBHUuCFRu9/IWNNqcwJOD2ruoiUWf3Aj0MFOQ68xR9HxMDoMeC+Lwxc/fk873
0opVkbEXj6ukQgW30JLotjbUhaK/xrNivynNMMkOWZ8ooQ8ZWc4JFXGvNAdAhXCHs4gOATZv56WI
V7LxjVdYBALRKPHa0Xdg8KIfyQjlzfM9iTCEy4dSPZ28XP32cQStL9QiYD5GduP3qOPMva9srpRO
+MdPvVQZe8paUQvqZd1uUqC5Wqxyo08qcTJNvODH2xI2xyai/28zZ+hZ9K5BkF8hWOD0mNi8OwrI
HUcMCYapl1VZa57WeWiic1x32xg6GU+to3sYgTua5uFiEKZOlrVohVGpYQPw8H7842PKhrUNEb9p
0xvIFgUluQM0xMuz4IlUUn9YZETfihpAp7AewpGfwMy9VXfk2eKK02hvjKR7EEn37BnPZz10pnPL
8Y4Ellr+KvdbmZJeOyu2wqBN4/MrHLtgzaiPpXuZ0SLhpjkOm4bTPKwLUAWGyLzp+1hUUBjP4uhE
+mT02bq6Xs4TNiRKff5n4DYCGM5hmeEEIiNBkYIyNs/tjtfKb/cZKr1HXLgoFAeRXxD5CezKwkVA
cP7CWYy1GfIScUkfZpO4pKi+5G1YbKi/+cqaYFH1+hO47voMgY2RatvuWQp+WpfPRpASAWSfxTtL
va4PeM3waaYbu9cdR1kFhzqdBWyymlU95ANFj+59nmiXPUcHFqE7yG4UhLPBUp5tD3QOrR5R/kYN
B7PeVKr0Zj3gFcTVvDvdCT4lFKUFygN9nKf1FQg9cKePI6IkpY7Gmjpkji7SMdZD5bv9HUkVCpe7
Hwtq1qE8QtouiLz0l9baCkeUHn9FLvwGDHLvlKr/UM59jzi3/ivWNhsaGr6mc2GDnJJdTSDMsn+p
7uby4y3agY7i95MoubfmvK9tGPVqG9EfNY+SjhEEcvkrz/CJr7PUBZYAiWjC6PanpOIqVOcVuZ9/
qJqyNXoRP+sYh0oeqSMmsAxRtZPL8OFz/cSiund+Rew2y9Gbffcw4R31T7ltTSIF7L38wByx998R
9uWph2eJ0H1lnRx5EJP7uJnPbgnUI9T/wOGJax90sju/TM+sjb9vYwCtKvrE141x50tgREVqmhZb
0XNQBsZxxEiYRwAC/sUjX3mCOh9x7pWzu5KKPpz6luu9Hc8kv3DEsK8T8TO20mXF3vgbF5F1VI+k
NmpQHgxuiIN3HaMIXdE5l6pwUqKBoyIM3Srw+MNmR8tyT+XjSPhOCfjk5yFfqWQqUXaDCRrB8qxb
AnpAU+eHXzKb88qsZQT9ALxuce7BJpHAAfU0rZzcSEXXfoFrGSmBL2N+AswQiyBtoQK6ukrHbioG
OWtWh9t95Mr6cxcQkrd9+nLT9LG+FbT0t/aJDC6WWoSwG7/+0Cfk1De1hIJeqDe/yMvTYv0Imxum
iJPfuoyNZ6ITBX39hIPm7ixeFWuNaU1LbnZAWWD6abaUlksoO2BRHgX6Q27HKL5Y0jwXMk9aVuGS
OhQV34kPa+e9XV7UCrEWczbv4Nrc+/Ay8ccCskQ2H4Bgi4wVZpal3cNQQzqwTx9JbUIrow7AOpuS
nBsxOGgqWj9PMT6b9eR18o8hr4FuKAkuNRiINqY4prs+Ay+FCubqz35Ptu6dp9KG6YTVbareDKJQ
LUJwQ1wyOF+rPItRdPe3XiNR8QULVovLR/e++zq35aTMw5qsBoaRmoVwiMsYBdUfsUIvEEX2VkDz
8XAcCRg/xKBP5hIG9WDYHeQP2x0roCQ5NvFXUO5rQ0Url01a9y+EUqeDsjcSJXijDS5VW3ZgGccI
fb+NGNH8Qot+M85BlJulnCTgyFpobiushJyG4pWmHdQC+XDF9+TIe0Jy6TWw+kewhgiACgJWO77V
0GwngqT8o6xhbBIwhm0bCfjkyvbKiD/djW/3dBEswN37pWA5Y2Mupi1AsVctUZNHJpQ4moyooehy
XRD2MdZfHqtwSVyRJtE1XH5+WRVxSYc0DhRIUhaKKRAbA7I6mHYbDGBe0j+tcM4Fxo0sBayl2PI+
6cJ8zdE2mgyms6sPGFBVE+xGyGmJ6wgP2KmyBnqGRpemaWi77/m9sL2rRSANDvtZP30fJvPdtdjS
SqcJbDSSEGJXUFa9CZ958iomAAnqnZomsaDRELK67xW9Ee1iYWL9TnSyZhfVYbvSSV1RfF+a0lGe
jDOjMb5n3g/G2D+0bLimvwieF67YPbLM3O3oVm7OQAjmrpS7//FeBUBJY70qkoAPTgnoucAQurts
oo12zaC0Gj1Nlc6q7/yMW5h5jiiSU+EM2ZW/hPK3AZvIt7sL4hOpVrmz5qxWeOp+/FR3st9JptR+
CiaOtgDL6qUZH4+XS19RZteBzPGBCeCQWs5lzg8M2aTULpRzjm56I6IzWshjO4byTLlxpF183HeH
ZGAM0NuH1lK04uUDb8xDGyi5b66aDXrazSpx8O6vIO2mYc6OC0I5OwxXpMssW26UYzyq2Mwxh229
OGP8RU80kIo9AY+/1aU37N++1tjARoxGR8fLQnQnfYjtK7erYUBcyqBBVtSm6vuQoIl/Ve1BKjhh
uiOQ/vLxuGv/1e2J++IOHdMJQd2VrsRkIOjOo94zSy3vaXPOAAQSw+MN/pXBgqC3SZjE3d++Lybm
VDal5WwGbxXj5SFG3WK172hjz3UCaxzDp6O3eyiN4fFNno41H/0oN4MBWaCKnhLTfuIoqjKcrH5A
2gGi07YZveyoat1hDMd6HqHs023rLSC/Vb2Bz1skWJ30V7LKvO19mga/tNd9ki/hxUWvmvkCtDRR
2kadansJewTkzkUvis0HXGN0AAm6/qXZ+FC8nbkzGqM7g75ic2abIdLNajDyervxb4fvx/uAdSrr
kQ4FoVZrbJXamEc70l0AEGVgfHAVkoDcO2ugoGbiqYVHFLM2TETYCDYxCcEWJvmcNykK7FxSlawW
f6AodPDZdjE99mPb6C4GlC2TjZ84RpEDcsQbprhQ7Q+Nv+cApZqlzJxx5g9cSI6MbA0lHdWor2wI
pQ3AI0bigmOZ9lbMMOFL6nriXxWv4BM7DEPiu/fSKv0uss9XKRIh/C3l1fEPs1+Cs27VQ856wJ9M
xJmEJfAQaBNccUpSEB44pxa2WAmToG/6R7OSawDKPilR+uIvDJlVmuCUp1HWkUlGVwkG+tJreI2y
XiOU1baPoFE2xgyyYEJJl4APXIOWYyBQLz8HnnIbj6x6/87TMiBiX2OP0tuvj9lrt5PXQmH1utER
AkNDQb0oBpFWd1Z6YDpvBfMXGGzV5+Z1MWK68l3zhXVrO8WRTw0zoOqcLCKeZ3SQGJlsaxePBk0v
QrMvfFsVunQsnNnFlEBlU5Z5VMWlMtZZryu8Glo11dA+ahhNC9XH2hfpsKmSeIl2okVBrdHUaEmA
sivZP4WKaOGPqPeGThLwkjHjPy72IICHpg9zwdmDrh3G2eIvAAtqtD+abDR3jRvxhttjtNT7RzWI
0dEI09bksDYL2l+PJ+c7llNqN/cKG8piUaSzFSkrraYg4tb/rdw4KB0WwOZQ7iD2OYRqT5LIKIoD
23V6/hEqNSiXkboeYl4QMWQCDx52BVj7s8BuXrmiSXiCfX/4cDpJxP9gH8W5wdgadUSDDe5zZshB
G+vzaQ6ubPKkwtdjeXT3URiChaiYECD0hrrSyBaXlaiNICPvdDyr6G0yYVPGn+uW7dI4qQPn1jEU
wm9W7av2eP4Y6JzjNlaXeUIq1JMO/9Dl9hZjOYjeV/WyPrmIWddA1evlTgbvqIZrZmHOAzfH/NSS
i/I9X6wEEsjdnQMpNVjePYhtdJGoxeLTsWEhXDf+CwQ3VTdpdN5ntxtwqraLypVBJVPSyqsORP6q
aiQFckr6VD20Xptijf263yt7UfsgkfDGm2/ZnX0EBk2Uw6jdHSf7OfmhCffZSSAEbucoONOx+IYa
PHwOk+sQPVg8A5Dn8u5DfBQYpRksS9QmXHZxi4ZQrTIxsg31w7uk7vzGV0qULYAXxGBWODf1BVwb
gTp/N2bsCnjsmwegDVflCTnTXzWM5mAm9dnmdqI5W4ofGEoU1ku7NyJp9p4qrvpsNREx8mvQSb4j
7nOrPrhAp4UNNO4cu61wQE076K7JTgUzyXsq2VWBU9lhsfDFTsIViIQxoBZ1ELUiwNK1xEZr7czv
NzHghFzrOhaVHrGFGx7xetDGtzZDi5OMsijW2gnXdWlfo6nvBiBB0ql7iglU5jJ3ogVf/XTT5AhF
v3wQR8MrinFIh6MMKvZmCN0dJ7+W2T7XMi+26V5rTtnnBl/j7yXLvLHgAw/sfpDQfhkcydWx886Z
b4dSdLe3J4jwYksU2i9zfpE2gBE+JcXHiOfp67VVYfQrMpFatWvRCjwYR3VdyCJrERWXaRYHYm+g
zZgQWFOdbnDJlWbpJjW6aqsMSkZcO5wpwFTtPeFAaEf9IHbs33ufVPfLNNIdrg3WRS/ThLbQ7/MA
IvjXJ61SVFW0BbKa4rHU9lb+n0ozol0m0U3tuge/BsXWvrsTVmYaSWCWnZH+KNESxTRWlWV6Thy7
1kr3VvBK7qDfqTi0yN9TMyVYlj8Ud5hH5KuuCmvO+01RC6QNDH71aRHhB9HuykDAZggIubP4EjY0
qjvIfvVCWeLs6XWUCziHEPq9rSqzxeFfoMOrYzB/xeOoCjC9nW9zOA173Tlz9cIXlMLeMyUwD82e
c3SgxcW9kI7IfaDr8LJ0hk0xrCCdIqyVXVn9Z/RgkZt0eHLB9ao66v2peU4SIh1DQErwyaJXRSDZ
N9SrYPPvee6ZzDbfDekGjxGykuhOyypmifXhLmsJUxZ/JjSPgVe89K6LVkxb17OplYNpVh5hpPdr
YGhtalBwQSKErPV/C/wmIgCD5eBdwoOhC3kFSHiJ5NCloRhnsvHw7QzLPerTCmJQD25LkqrTJEQN
h9Tw2s6mMtwubxd4AYRvfcfZ7plxgt6uUl4p3UBfESYfrkuNBD+Ddfg0B3fViqoIGWgrxoIKG0Bz
p/HNq7TRgKk2IEBGtjWh8k3KcxTqCgOVX8fwwzBGZjCRjwinS46OkAfpv2MFn2CWPhsGwLaG4yVZ
PVRtFgwTy+KofzpPt39YeKFLftovO8zap/yiAgk2I/1whNc/fDLGBy6SpDUg72pHSJrw4/ssoySn
nem1pj48LQQe7WTbASw32XcUN2Ew1BEoDS/yU/ufbBS0quXaqrwGZ/jFlkYnHuK1pc1jys4hDRbx
s3d3/kZEzgL21O7lE9b03qfNbz9H/tvwQGeOyrwgw/yD4QVo0/9IGu1GyRvghO17XLJ7f/nWNpMd
bHnV+IYbVITxon6g6syn4HESYk48oL3+9r1qXUeWLPUuX8yqFhwvDZapKjFVPvyS1H/bWrQEK9+V
BimA2dBLxT8s2SBU62UpUQ0OQnAn9y6wEZOfqCbWqBKQE6cpr4K6skyn8YO570My/PSpkyDfhJqM
ZpRuHGKi2s7+ngnejEOYjMNrZKPJ/jFeP9iPREcRDwTckmnubiB7FBWC8jVm0soZSSd/DzzLGrjf
tmZA1Dzi2qYZHadOiG4O2dfTblkw6wxvomBlAqdrWbggiZCUcH8BLOR1NR4NZmp0rKrxlAwYMShp
7Tu1cFIjVmTzLqhtI2yzACNg+cwDnyl4udAhpLhCfj3zaUkTepNbFQ0RiIIm/+auyNasYgTSGeTF
GUrXQXUCjPM0CYs1iGFd++3UXrMLUhajdBBLGbigdqHaAO+2a8HRFhIsbgJSoPE+o9VpbKwvKPdv
n08XiYPxuSaqbg5i0lgO1zzDZBXnu4b1txOtcF1j4Zg517+mmi6+6M67+q26W3fcZKdMvRfaJI6y
zlWAK1DK58GFxnHSSzD7B9HI8AKfePGqqFE73pv7oxRGCrkldvfM9iB8UT6yD4ZFgiUc33o5oDNB
GzAcqILH8ptmgzNq2AHJUK6HofSJQHLEfeN0Vbgff+VGa1fQ//vpAzG6wbNATyma3KYwsC1a3WYy
g4sXcsftreajTGM8x2kvuPHMt3NRK1wpCc5sa26CA9ncyZTWVVKfyITPziFMH6RttUKsBIrrc/ZW
NeNxKZIwCauk4YRNi8eBw8oubHqCuomXkVrXA9qdhmZyj2FiXpx2vnK2ORk2krXvW8ygPGl7pEWN
8mZ0lNq77sjlfh6gMV9Ty3CvOgMT2fy1ll6YTDKb1aYXALGov1FShcAovpZGrG1516BMLcV6rGHm
MX7EaH9xgJfrRyy2Qs0TjInpbtSGOE2fAfptVzBhS7jtFHJwW1oOy9ySFF0hM2nd88U5z0quO5gi
7i0FA3wMxfr6hzDAL2gzWYA4XJApwAxX5j1+WiIB2tRlf2hKnHuYf9yrRl2erfTbdN6kihVhpYS4
HOrOzIGwqy1MUuDgI01ljsuGOR1K8wSI3Ux2d2N3yKMkZkipEwYBzD9Unx2yxRD/lhyDEDoWQW42
6Qyy7vKtlraQvo6VOiG8eGXlAJBhRmS1Racijf63u8u0GuXVqK7MhlToFdutGRBY5uYAnnnuHiIC
WEephaSW7FRrNLoOGY+ikoMzAVUapH7sO/kFgVbvPgZ8Kb7hivgBAmdgflHBRcOdRXJCt1ck1UkH
662BJrnjnNyW4cVsgqxyt46t6QBVjRrlvFnOkNyNBd3/hL7Ojv2ts+GA0fASRpDhyX28FHPYeQwh
P+K2yM7JoGKNcGu3z8CGjAIixxC1oN+OLNPEatQ0q5+EQ5oFL/GHovZ0Sr5IpLpqAgbS3Sq9SrvM
Xoqy9ZPQI0X7KjkHQCiVHXFCqaInyMyAzLRZJIHX+hc26P7l64bmjhVTmq8VdP60kdO+90s6nRby
6LUOnHt/yhaVYtWUGp0nVN5E9ume9pLCvOhnibKOL+dbeM5yx/PxPqQ024M69NIVc7sxrTsyLJ7m
JZ1TMJzmcopCveDkWZ8oCNdkR08hD4Xp9e2tpZVh/RUOcsqEqG0iJEgIIKA85OJ+pqFey4APjfLs
y6W67WJksKLvCjEQpCY9cCcaP83td7ygM/F1gGRSrz19xSokl8CQHEadTWcaFTrzrB/QRizL5iMm
Mn5j9Yf/tLV39ynAICEa7M3kG83UXMHmMVH5V8+keOgcuIHqY/20rsKnGnhq1V4+arEno4BQ/feE
ZPRGSbjshXuSUycxrsaZkvIVk5MgZnXUpl4S9AFS7Wg3dJY3t3sO73tFiyZo0DSkv5H17/5I6ZUn
FFVTwxFmu5ZWXsAnFXcVoeEYTOa2M+s3Ti9X9V1anErsR1AlYy+EWOj8Lys198WpO0htqx3INEbf
9C10WvCLrLRCz2TxN+8OxvqTietIR/oq6OFrwSIUCo3obbvH5HcsmTZbTSMBkuxMB1S4Kbv6NLGg
WkAFZlL8ny/+8BrDNz/4n+V6e2U8kNZdqeiPELpTTYVFHDnNFElYQwdZ+Dwt/BOz263wS+Y6mTo7
soRm5IzjGoCv4jmMUxIDII2+Z28jUSKOqh/JO5uyVOcPjefdtW/v3YvGJzZ7+3VTD8Yul4JbgSrZ
Y6wU7CwjMCzBY+BdGbRhdbRY/jye/VZLWRxnybOTWYcj8JrSvE6fvhFAOvKJzAg9eoThk5M7gKpi
N1HncRYNLKhz97i1clK5XL2kIx2DYBfTvctUkJZSgyHR4gPQuis7FQ8apESewAoM9fLQK/I5a+fM
uyMhomxn2GomOFKSp1Lnt5rkotBErdP7th3cMg7M7FIwbJWbPK8bZx0YCmaXoKy7FBYsVfkbow3G
lokDOiXL7kAaIO1sD0uvxsr9HJFIf5Z56d7/Dzxm0QD2y2Vijglp0vRJNLsvxi5CYt5DKnIesihK
rjmAwESDNA2I9uqq4y6dc4A0GCS5PfhW1/1Vl2ixkSngs5Nhu9eRDY5bC/OT6VaoTOKoI/pxj2CU
5TIh4k5O16FSJ+AOeCIvYJWNUAVI+ssrh4TWB07acO0FJu+C/aTvlc6zfd8HXz7ycAEbZdVF6tNr
TSaOsctu9dw4rtv8HVJeA0gE7b5nqE/ZysA4/lTHJ+TMsOaL5biF11GgBozweGoFediAo7BlgAPc
zbmfRYDHRbMBEsRMEoUd59vsJ592U518388lsPn3iYpUmJUjLPUS5lZkKaNJKZBqxpdOsSAB0GQf
9cnc0VFSf1yPgM2AWCY/v1TmlvVoC+5GHkS8j3PwZ9hAbA+AyNBh/DpjNZpG2IadHFBZemwhk1H/
Zg+kyrF40lhVv4+eV4awdKAhy6ZPN9T3h35Hrhag0kmOS/jsfPOp/dgqxeJQWMU2FuaOqgheJ6PF
+gnhfdRHoGTC8N4yhvDLAtqXa8GWiTxEFsHA8bfJMmfiEp+bCDWbEOxpXTFabyjDtP0gXidYRR8A
6OU1C5GSJIIaIm7dwoQILjOz8tVvFL5FNLqdivSKnLyVfkRjjuh+5/APnrYgy0y8EYh9T6sc3Q+q
joLoLLBQIVGNKylb/VeVbtoASRK9FDX4L5aNOhEL25NW4AoL3fGFErikTxUm07iZNiV9InOrLsm4
c3zd+tSZdWTyYYSWLVWX/10ZvUVHBXUTWZKA8MN04fATacD2Vf0VbgrUqIfqDMEuRiTfjE5WN1Ux
biLfMbiNLJeTEZZd4XBz9Z9hfQHg0Xb8edlKPfyDd1u6Go784DMhkmHubtt/FQl8CL4d6HY6um87
xYdY3EmQMFlsafuAPPohNtB1CpBXWWrZJ7aYt/RB4kZ17MHQ/HVzmlN/n/Xi3d7VDtKdCVsq2D0f
VuAIMtEFdPIeWb+aEUDvfLgqbQ8ozMKBTtDU2vJVW9mSp6xBgYalxIJCW2QCaZzdkCarzpBbI4QA
qbbXcympCUyU5pSIyjRlUR/bLlDFEE0+IUhtf+vhvxqRoQF3S2MqspOpuCud41Z/+EQYUBs2/RIS
g0hgmyJH/oQhtZ5GSkFbL+48yNUbVWI9is4EZtOebOgRgcM6KV9mesIrpVJUYCQdB7mw4s8YuFjN
WCl2gFOJwWJGcY/WyqnGmZnHLP9Yt8Z3LyJenSHiOowIqYTNkPp4XQGsr5LbTREr4p31YiGyfoi2
qltecn0UJ2bdomyLRtFWcxNseZIkrH9zexjPhcbUJGhcpIEqztrtz+//L0g+Vh8F3kg5yJaQUVRi
4dasd9ix7Jaf8O/r9DJNSDDHKjqTfY9NAxP0zJ2e1QgnzNZOfdmK4z6CofRQm8iChvplcG7Fb117
Zxbc4ED2NKhUPhswP8c6sFQ3TtzxScXjFtOeqlYQd9xEr2B2n/w4OOhfOFIG760ce1AG8Q8JcfNz
zeVUclDfMLBQkmGgqfO97aEVPJRJ2/jwTb77SXs4w+8aDg8uV8M+yLzBkN6O6ENmcnnBQ2Sf9woH
y8kfFhsU7knhIB+oxNvZB8dBkwSr0MKsO5vr84r46lB+VUmXUsAmd/rIISdR+GUmxtZ6vFC9FIZx
5Gb5BBEnxkN/hnoJ6F6w7WBQPRx1A6YqWUQmuConkHYA0lk3tQz6GaKharp/2pivcTE2jkpvhgK1
OPjbBB/FpAKfssUWR5cNA+U4ANN4NhK9ltnl9Dx3CvPFKWWMt7W1iXyMf5DDzpKhY8/0fdpWcL0V
JdckHsQyGUEjp79QiGz/WpY3lQTqGEJAkrZSX1BnyyCPhAccnaEKSn0q+D8U2gstUg3Id/5nc8ZP
hVoo39oCmXk6rov+YEoEiSCt007dJfDQTTB9WjGy6kU/YMTCVw2BSc/QGAh2odtF0gkGuIzY7ICr
Ybxkd3mc9RwHhjqaoolOyeXJ1/DADdj9zFQiv8IzUuk69qSDC7TFyS6K79Pxsgp77anYJq3QxvHd
F6YrayzjL18lYAHUH/fK4ZWa1Rhodq5/1D77niAb1/LMSEeauYYR2r+Klp7+IBdOcSCDWk6UW+Re
OcaKU7nLOqBH0I+XKbr75C9fO3S6O75UdBL77TVTVI21W9WgFXYMAkzl9qsRwJ6fdPBxra4w8q8h
AbP7ugLPWp8Qj3SFXjhkdegSTVFQFBZ9d6GJ5mIhO+B6UW5p9Xz8GeNlEeLqRbVQ4VCQ32FWwQ9J
O/h/re9pGrcSSItNncZHNrCdR39jj48JUspJXL8IAUH6dyW5zJFBOT2XnT9KYhhwMNrwfnlGCsp5
TwxG+7BMHgW5FY9wIe6DC68yjVzKNr//70JqMSS3UCTr/UP5gcN0eiaT74kiDbQ5BJVHf7QLZBm+
jevwJs49FCo8ihONaoQ3a1wN1S+IpMXLT1IQwazF4VQCa5NRlTUg1UNDo+AmGCC8eIOBkXumv8Mp
V6BWwOyf5Y9Wjefe0z9jxCUajob58fUhQ2ZA3q3Jz+pbN87HoSssJnrf3ISG5G/YSfmuEtmhiG89
bPJYcunkE4eknOomuws+WvUR41WUetyoHTHf/6SiaOC8DeCdAJwaN1mX1twvpfK5I1wxALEqOP/u
8K1SBmukU/giLr65xXT9XMbqc8orVBpREWi+Gq/nOsXLCQSZdkPuWrf3l5A/PF2S30IXCzKM4Nrg
KlI2RfXhkfchi4u4dtXqOjW9YUshBGCgTUizvzvj4cfKbI7Ht2ApMZ5UsW9/5aAJ1YNSoiQEvUmc
kst9AiXUJupUsDNAXDEfyxE7jCazjoz8tf0U6SL7H06zTSR6wP/ePJmSVO1dr+M9m6aZ6AQ/MSuS
K8nHkn4JGMqXErGRjU9qlD5uXAO5agFvH2Mo4vy5/9K4Lh1i9+sKwo/MHFvILVikvyW5mKHyzMXw
4m2v9votYyKruqJrj+9RFOTOrGHZ+BaYcclH+ttX6E8rWdvK5gPd4WWiDujDdY0a9IEk1FBoGgv5
k/k1/hiXyz0ykjUUqod3tJ4E16jg05Mqv0E4hGqf5sjNvmi+WTHfqpdEDayiFULqUdw2B3euvXID
jQDpPqwDhfoD680TT4q6naNZRVbkSDO1et6StInYw4vRB5og8blL7edxK+BTB3k51kyCvr/uxU13
ShfAPxhRIWrxzZIbL96XyhuLsPemXHt7O1WtDeCAoDRGmK+JwHi9LcNpnnCKTDrxV/+hynhNaFdC
PfPXhfaoFXbLo3W+oXvfRh6SLow6ntrKIqIhzA5lr4bDfEZmXnNGBYozZmjGc1db2Htx/CiQ22JS
nuPjMIGDcsXZCakb9bsM7Oufi3BOttgUXz+VpQQZ+8EXNIPtDDlEE06nSZ9eT598R8Q1jRp5dyaJ
On0gy/hA0ZyHzQGgNdMU9ltlEZCXQy08U/ixcAtVmc/pLiR42nY20fUzLcgFJrHSlUdA0cEwHf5L
Gu46pJTw5KQSCCp+rLC7GwZnIC79VzJKukpeIjRB9TmVM8FKqkPcJYtqd+CDRW98VHDn66WzZzLw
iG19PpyRX+nulevwjiZ9skCd8Ae1lW2IbvlENSHMI/LtgWaoknPWjBovhQyGVatTGHYkse8a2zwC
s8gxMAzxaNvCMg3dFEHvAuwP+77uYVBr/75qqEmYauhhxaIthRRSe738Uu8+t+DSVDtZXUcbajJ4
wGbYxZ5GBzE65DOO/KlwtFE5xC5gDYrbdH2g3xBQ1klZ4L5cABDRkRKmOGu/tOwbnMO7ImeI5ND/
i+wCgl8PY5lBZ+uDbgJ4IJb/7fcLTJkT1d8/a9QyVah1pnvdmzMfvANu8cF2GhX0FumcmVe6Pp3c
15tzt1EE8CPvprXpEtIHUO6eWFNI3f/6h7eI5oc48hwXtsDEsnl35ojq0tOvozkLALRruwHV68Qh
UNkKoDt2Fd7SYKyG591hEWZandlvC0ZFY4O/YcyeF8JG8RvrDjT4wMED9Ds1TNv67/mjBsfQjBxj
ISsrC08/gMl7eUo2ARL1Dm0pAysr3hSyL8GMYor+7F2khNtTfdVzyR3hLmdC0gSbYd5v+aPdMi/Q
FtQLTk8jne3ivU8aNTnGgNw2v7GcwnTU6c7JJtZ5kx0kfJ7lfPE/DLZezOZhgXP2S1h00coob3HF
8Rfi1/zVfZVmxhNXKoAvwCoyhjEuyVfzEkSW639e7RQNJFxSC1YZhcdfAW3I3kY1oqcorcT33pnE
+GEJM/V6+pQMWQP492e0+VDSlx8eopWldQ5DZF/cx+DM/C0iBn7O6iX3TB34O9BkvaeIR73lqJHF
jeahi/2a0jfmUv8ysjPKwmEYm/mZA/sf+Oc1O/7ubvRlkUvy8CV26MfyfzEtjCI22WpRKqWlIe3Z
FOSaDeaUluEM5Ke3hhr2N+yVLQMY8gREVPSLXIUR8brE6dElC4JFmb+3v2Sdc1vzS7LpgUMOqVO4
6AFFp4Z+dA7oCqKOd/IPINtuAXNbyCU+1HWdFFgvZnv6N/N6SWrEPurvzvN/Lgr6TMCfQlTXhC3X
MHKYuTkCGcibp+L8qunwcz/uVjcfLMPcBBy2CqaUVkHy98DhtcuZKz1K4+GcH+iXFMGL29w+QH1F
WekN8a6ijRScOKuLycgTCv546CYdw23Tr5cUfBXXuR8UE3j7EejJLb81Fk+NXpRqOIaQJirHEb6I
7lRJgSE/jvcHlaQkXNQLQm7VAO8uKgnh2ssJEEkQ4Or+YgylIxBSFgxNMR6Sl0ukIxSTPRN8AFBI
k7HbM/TZDAlWq8dlaAXIq9u2z7HEF1e4qi0IQeVKHZ+fws5BTWbzfCJ6ONJ1nryYYyZbu7umsfXn
95MYlFkRhjAiX6sE0NunhMQuLeLSfGJZnRSWLzoQwW5QvYrYKSYViYyjt/c/NrBed0cPLOptKW/h
m/7MKE8EiwNih3ncG6bWxxwwKT1T2UW1OsQbzttxISqBQwUtjETagEQ/5MK8/+z4Z7kSM9QeBv3u
7UL5uaFtySUMjsH2BZcknOH5lPE7T3Ip1wJId1VD65cC80odPhMjVPNupPQm+ejFIAEYz/zeLxXW
LHhikNC+WI5ig+k7DuyguHGUgO3K5n1C7gB6sg7PsZg29kE6U0zbCL8T0vdPaOQyo6L901yAybQA
68kjsncXbBx35Kmv8gG6aqMUk3csKeAebXIhbP1ZR8IfGBzPLWrQbTRmd42SAf1WnfRFnmhajkT3
K6XOB61zptNwbcyQJDxww3YrasbXvHN+BK4TRFszwWJo1ed/yxZxbkKwv+y0rv9zSozmu5ptefUO
07fJG5TcTWVMtNFs5n9t/PWuzQYRYlykjpih0Rry1qRD44ixrjlWEFaDYu9wetn30RNQDgzXhBua
0ToGpLAc3TxR8gus7wWSqaKT2P8MBS/9+2nWK5Lyv4v6AzU4X+Ffao+lVRQdWFQ0YS5jLG22/8/o
+aWNRvHwK/J3Y7gKaU8qFFUPM7OLFrLwLtCIq8sSW7s4H11UGN0P1D8XzScoYz+cIoLSKYlhj/vg
cgAr66v6cW6Mj2R6Fjp5ISepIPXlhUZekJhQGgIVp5xcf5HaCHDCyuKKeEipGZE2WI7zZOYOXOBH
2fOzWkU/JMBoQIWUKyx3y3BcbqUkdhJ2Gqw9xAInHaX8E0GWFz9vfMq9fD+g3PstpE1LGXT66u7Q
9AMzgEGjRjscpIot5nlhMQBXycAfFmWIuWXqSkqsZjh2KF05TjhExuygUgOFQ+5Vs7YDK4LxSzxq
qyHkXnNZkojOQYFAsxmYR+IaGcSvEazImesuTKx1R/3CJZ8D2t4+mp44k02pMm9o45g9VO3w+gHV
/1FRHlsjJ8lt4qqjoYXd0mcIjDTvoAhe09z7arQrx0V2F2eV+Lu5gVDhQgKxf8FuoB2wHnj7qw0N
ns6dtXlFBb5JBOUFnklec1PDtLLWQT2EM565JTWPzWt3T6bci2oa9QbjfSyb0edE56yAYVYE0ZMd
IlF7B+mHyxt1jU/vZf/RgZBOohJSGcf5We3uMouKj8aXTsJOS6+grSdfEUfjhOjXZDydNkhIiRr9
CigFWm/2/jDWnvI1CBq5CzsKeNRe2usdgdvIdFWITqXpDWKxOvPGgLJIh6ut5ao1bG8a4HbvpxP0
D/UvFSusYu167S0ZO7/0L15sg3zJEgaZAsF8Eb9d29tYIlZ/VW5Bw+Nz5DthUE4IAOUL5XF8ipJv
JWhPGs5jq8igEm7BMrb4TDOeNdkBXFL8adZ9VbrYvPst2mxx1KOM3pX0aw2l48GW9Wjw0XdxWNV9
D8YiOf+cfVqc9AIazfXQEIasgUGU5hHBFqYsS1O+LGliOnoqWz93i70DN54Somcn4IGgXTiO6Z1c
7BLgk1n1lmBSh5A/rwgEgL9BoTBCsuNn8aLJIm4SHtwvTj9OS1NEhy+lfR7e5fofdqV3GtaEy2im
rzOardOsyKDzGjzclPbbdmLuNg7Px6nqn880pac6qGiZ8NaAPpjrRi6SnJyD1V+sWucgIUEIOKM7
bABaStav4CAaryjHqg0gAte++FjEwGZcfADaVnpBUvdK9oer50ZAdIS8z9qZX53hVqpOylTqs1AO
t0gxRHFXEKIx2o8gExZFDBVWjs+/rsXorCnbI3/+8uxPOlPyNUQCSDjXVXFUw2zJV9GjiL2UJn9s
D+gt30o5/DUymolzO6Q+tuvjhjHHg9zgr+GGYNRQAeGBTntP90HNYrki/LI0JZXDYK20Of/D4yhh
XOt747jmvezgPogyoFqWyfintrAKuMg1c8HHIO4ovLmPhfDzLmitHivlfmAFPMpAaG6smnfWKR0W
wMUVAl4BAbFBoIllvEgePHd/PVqtgdMsR4hnXqVVnzJRCqP3spkHNJVneB7vajO+VkByc7wUIblC
YFMFKw9EcalH14xQT+yJmYRB1LKml2o8oTHyvpYQbCZcQ89KNzOBA7uOFkAJjva6wvqRjsufSTZq
Gx8KAjqyAasfc09omu312ytWAxe5lCHelIq8qcle7yP+V5d/l9g+EzNJKxAfbznrLOKzm/Zcr/RX
9c/VaHfWjO33aNjsMk+ug2hxU6o2MFeV3B6R4z8c6U71Q4g6MSXgc4JRVZoJyu/rt1qHvVIFem+9
qcWE4BrfulSThuLvDctsDN/JemvxclbTAFbOVJ0X5eoykldyomTb6WKz+dcX7GNpbZX+wN9OoYFv
A8ASi4EEaCAWn3WhDqdtZckJlOIDRDQpDsVoStPfv7q/oXLcLetk83k2AHbXgHGx1FGaJSvkCGXc
oMBVRqK2Wf8RyQdF1i/Tm2HKrwongUHoRbxeZU6M499rwrggQVwmv3npn940EcJCbIqZb1GtydDr
UEwGplVdgrwqTMi8zDryl+1vxo04thGs/5TOSkeDlOAEYvWUGv7UiJydYBA9W4BlvpBzkPWGV3u4
LMz9p7FbpallmjTUQoOWUH0XSWZMQiUVX+gzYVubWVlSm4gO/4mwB3rliefqJJNZFUOrGX7E/8Sa
TIm71HhfbZzLdm+n/tRBUCE7O/wxDGpsBe+EsX7TseKsG1mDP/Gmx55K1Ash6nBtbiljD0eyHgDP
c17RH8vkTGHdBnyLpxB5FP0+X5m8NxDsQZJ1jcThRXVEyWcuBgbZ7gJFpYCFKIQ63dE9db50jTkf
tlJoKNvU1ecqyhGnSuOdT7TFPj1SKXU3WLi8T1jZgfnmmP4NEILTza3HGDuDdYSy3pd72CcP4BtN
/eUxzmlTgYji2c91+0U0qy2R4ezbaqgiRkPPvdEg4OS8CNK2JPxKQkRRZ1b6O8QeO2mGYFr/12KB
F0ctdvhOJIdJZ0kru5ZYELe+EwdOuP880ee7JtDpQWekDpcZb+h6K8c0PBF5u0kR7GhwGKkbezCG
UzpBiGLWa562JVdqT5o0JnFaJtHLBJmp1mp4icTDMqJJ67cgfg9E0Mb3u9WeuOV3b0bxWL4U5FlV
d239N/4pf04KmX8wyYtXS3V+z8jCg1+t0vpl0oM+4vPTAvDvhwBHBMBYaB9SeFjxdPi1R1oc7LmK
+DOSYsu4peUq5yUzxMKBIv3graxppLEuclC4ihNpqTdoxdqzBfRla0DmA7RxKKz7jEjkoJEHb4CO
dXrci4yPuYg43pLyDcPealIvOioSFfi3CfzBcelsbG19/JkUMIiLyzP85sHL9gKK9RJSM2YqwTMw
V4HE4dSvYByah+YZISRzRFXVTu/NIIzaNNsAnJsC8XLrOA0DYpZ+6p2s+sbdd5bVqkICe2HfLZ0g
8R7kXXQs7cLYnKdibw/Q4kLsYTtZd/YCwgOL/GUD02bu88DiBbAcfDgmmTEw2qsE2wggv9N4yRc8
akL+dUhdz9LDXX40+IaAKj3O7iP9v2UuwNf9+vUk142a1p6uCsbXHoN5yAV/E6acWqqVdqG4Gfw8
J6jTECbc5ZEJVWgXNIVZ/MgZLXoxaY0JbMFpbzeqoE4CEp49NK8EdJ8Bc/UNpoXEYqGprD4suT5A
XjNZAvI7Y1IaXDzoGINpcZc8HgRmgAXn5nq/YvMtEAFJGnxU9vRuSqfCVaXAlA2Jlve82AyWsRm6
7fmUlfrKXhN1qaRngxROvrnPjxcI8NBIK5HfFzztbWI7HxZ/lkL2eSPGw773XnaIz8lNIGs7AGBM
sZgP7shNkPaasDaKA1AX8r0K7+Req4roZzEMnGww7K7mJYSX4cif84zwoPLtHB8rwWP9JFc0oEI+
CeN3xVA+WJcfJQM2RQPz+pzVEEE24/dnQVMRBEj+V4VH3W36AK+L2zy0QMpTFUiXNADPWMBVfokW
sH5C5eZUj96c2CeMbiZDUNKiYmGmd5cyUn+tVNLPeAjMyQFzCuBCCgAZXMEr8X4QZnL03/MKVUuP
lq5GTvQBE6EVowgVbqi5zFRHWk5pds0oVZQ7b7r6ppFwHRBHqsOluRlLEjLTmECmUMP44nK4iqjA
vl+ICtUHk7xGQG0aoF2S0Ts6nx7kZs2OKeI2x6NpMIHYAH57adfjdvqeTDUDInpUuM16vXfkjIj9
VYrz9Hn12E7gFIqprYj91wi8t4BoS7sSLwBuK4HOiFUX1mWbG/fL+0KTMx49F8JHPe7YZor3vpmD
1qLIMh0Kr5JbJq4Wjqg5lV8pG/Z8LkXp8c+aoDznyb8aWnBBB9pdt2wfeo951ZZxjtMggKCXrj7l
2/YxrMMXSTumoREwqHOldz6LRB/HLtwz81AwF5kYClG2SNNahXNR8tvPJ4acQUwYiVog4vnHyo3N
FzMavhFGaqFM7uZok+cflm9kktpUU5wMcWjteqExrTmMhSAja9JGwzvC45XAsASNl3zp4/CtRnb3
6qaj/fvbQQzHYVbbsVkBSeLaTSkjaNIePo0EOk7Zu3wraSQoJT0eYVdqF6oFF/GcWbC7cimEEGd/
6bhT0eOgDS9ZkH7UC05JZTLFy8QeLCiX+Ehv9sfq6PAIWtcaiCTBsih40CcFHvsRG1jv1LkuMLGr
kZ9n0/yNS1LKedY/R90ZzurxzJrAMT4LDcOPe4RDiKWKW6vwW/PUEUV0gnk3TEgmmjOHq/uDzp4B
lAjCyiUvkp2lH9iHY5ihF1gJe3L5eBNMoSK7uznroYWH+CQMGz4oM4tO5tjTnJavj8khfNx74P1g
Chcnhq16S+7uat3j7GYTg+RY0Nq2iMH23mhwGMUjadITXwv/B7IGqCGX4Sk2Jkxnpdpw1B/ajfFC
iA4rru8wMuNbYGlJq8tC5wkaen8lkg4EhwztYGSaC7SGDqV2hw7HWzekN02AOHxOcJm58LS/oG2m
JX+uAIH46l6cnf1Fapfzicycc5mBOqtZM8E9yfdD0rnkfO/BuN84kA4Ux8M+dbs8zoE0sazgljOo
tOHkQxSUf4NKlJgHjVytbgsbkxFrM3RP4kcrRZYgUHgQK4AlEo0s6aom5EpLX9I4vzJsUaVtV6sz
fA9ibYt0rvKT9OtNZqSJ1KhXsGCebGH8a4tGWWQUsCbOCTc69VZ3kiBIGKCF4z3vxT4AtH/gIqnz
JAPort2og04KOIcGzh0T7kaLE5fPHQl6N7Y7uHJyT4vQQLvHRutglGI57KaDtX9jPdQSZW3ugfeL
kMmYkCO0hAwXUVMxm0xSz7Ffo4tqfT8U6gACf7hULhJpNN3vI/XXBnyB8AiWoQdSAqCdTYzZbss6
W6/yGyMkDlKGrHzxQcamlN1qsLT9aKnJWTPwUNAsMS235MxqnLUX54MM2ptlnKPOhJsXzJTzXXey
s7kG/ToE6ljFXqrc8tBJNWAzeb8/vPutFzrYkU8ePSbd4wgb0aFjFbqEDwyhHfI4cbeDVYpU+E46
pZkV6CPTP7q7OkamB6khMniaAciUTUXz6m+PEN7q0pvd/P1UwQqSPJUePARuRztVXSFdGSAgpE2S
1gbPSjiXLFCTwAypj3X3J58bQ8XFI/EAJfoeCbmWqQ+xoePfS1jTrzD7WrFi17doAbRDQ6neQ1fD
lE9O/4FsSP2xyMjKbnkDAMpXudDgRWaaT1KKJRhbmqkv7Fyy524Nnq0BYaHdok2EBGkB1vueZgo/
9CiH1KVYcg6XdUyNq+X7gBiVcVUO/DaxWINrL4HzZbZ5rcMGG7DfPZlWnG2AfJ9Hvj7RRuaLhz/T
r5knIw7nWtPH0QMaPpX3+yVo+9GI9xFuv25w7JlHnIuugqxXDBS2cqH9jPxKT3S5ktOjNA8EklpN
AQcPZkD3xOin/WV0XHDwel0C/Bjr9TZMlsUf/Whxpc1nhmFTVD3uPTyOvsd8Vq0Ee9tmI+cjxQAd
Wi/c2swvtmsD0NItDPMppicWAc2nmbmbt5dRyf6U6JWfyw1NZiureLId5fsUyy8jNDLnAtYVZuHV
4ps/EuZFuc7ufT3J5zqtp3QcmYrj/5DCh6bEaVWNPbwkzK9ffsFSNg7jy+lRK0u4uoAbeedukbeC
mV2lvf2/ZHfb7kMN02IHD3Yi8lJ47YKaWKmhbA7sXyQX/0uC+qVbXtd495tT2d/7tj0lQ5hkDk5H
eeafLMsiOFQ6i11CdZNyxDIWF/B7PovC6tolUCZFuo0JwIImsok1ZQTELojRjXwRXLKEG5cXaqmR
2IwgHLQccX/ZohtxPIrEJSZWWm1gRt1NMt6uYUbVMnCpNv/IIhM44uvx5Qkq/GoW6znE/WptTIkV
aFGxelSE0edYja9blh58XC7sIBSBfxS/kYCq9BPQpYuHR58HhpPzS+bfiwN8FAVR9hMia/1fyVlz
Nf+KhwDjS9lY9CvpfRKl+CC8EQNbQksyM/G9nAImj68cPYdB5s28wnIuwC+GBUBVCx8U/aiGg/k/
aMPzb6ryVhpZKpnv8zK7hOSswqFxJ6a4WMUCdwJ7jjSM+kP2thUHjMx+gCSrk7a9eORvOof8e95D
HWL3Q5eRTqBsSgvDOiGoJ/FdaIB9D0w+FAQiPvwbTJwsPC1E7QoKrNJkzNLl+SaxQ1Z5K7z4I4Ai
qXhhiJKLoVs/j8PjoWABNTntQ3KgtUDWmZeR09X2Eb6B0JHxo/13IekyH+IHng10lD8mkp2uo2DB
fP6QW08wGb8dawi0vFzJOwhE6KSYswFSEDidUwjXyIJDy/r05xmQRlofCx0hXaowExu1xwu2rCqJ
I2HFVToUbM5LNANFIf78kZGOlR5YHEveMlx6A7D2s7TIMBBTwPl93AwaX7TUhJtzT32CCYcwy/v0
D/iHnr+OATHPqIgczsEEd1YyRu4bPalcT3A0bTZAVhzEOeeLm+Nf7tb6aTftcRTondPmwCN9FHNd
qXLVSQ5B5neXUGK45SR9D5X5eJB7ErSD7+tn0YofIrxIk6aGsoomapcRv5nP48fP6s1aDhPeHYFk
c6OAU1sx3p3tyM5iQ047Mp8xYJgIeEBNgKmDrr2l8ChzFlN1FiKYC6K3AF9M3Ln+b8dmxhulBT8D
bm42xOkP/tYweQzzfKLUUYmFxnsTTTVaNA8vYNdIS8rgep1R/9KsnjuUOfAmUIkGYqjRP2iDVFRd
eiIQyrJQwEVbiz0pHJfMJs+BbAAzQ2RtNHKmbK7MtADw0y6AB1yMIuO6cZaC+ep08oNYUQer8Ld7
Qt06H8OPehC29DYJmppbBsNUnX9BTywhfey8onlNgp8tDtGF73ii8iQmxCKbjWUraYqepAeYBwLq
0f7+K417Cd+sSfgISGzPFUZ+n9tW7HKfonu4sDe6Fe9DedX+xgMHXX9TdViVkda6AKd0vZSXT6uH
wZsqiocZ3s6cWxhjatfZ2XavXQBkpf9yq15W58vNSeAywlrnWMoy363jsORsUHuuA2INBeFqhziw
NPdmhJj4ORjI08O4r/dIcXymJBBPg6K6dgcpxYHbFicHpvELB1pJ3CdkVacPOmyUMhn6B2ZUoihj
I1NSQU/UOnKe4CpQP7KN8TT+pKYiWvxmtfz4OJDhXI1g8jdWVyFIGYAjK+RjIxu7hxsShWWle/rt
+SwywMSniWftE/KUSi7jbkLHX0VL6YsqXz4OSH5arwpwa9jfl3VvBDyDh4rSIwhQNOpahhMcJ1zI
F4nSFs7sd33O3wxHTzGGY6mu9tOPzkfjx7ap+jFIiayxkc88foDTQS8FcC9eTsNK7o39C0Eotoax
gdUUH7RATV4fqZucMJF0rTX+gaoTSFXjnBxs4bnw/NaokoR8O6DUA/S4h9iSScjxODypW3IpwAXL
36nvYKSTGr5mO2HuMtpHpvZ+akqTIF0UJjgG6bdLZwJAWjRzc/fZ9mmdVkWpd8E/GI0MHL+p/A4x
mSbtVFg/JQYP55lPvDHkpHMyEZFLGEFJVi8ar88mCFlE9JRm0d6GHvPMI47PMHoFLdZuAhhD7+Vk
QCcQggkLI4ynPZCV4ehXAfC52u+BF0HafS5iyUEpT1TZFlgwuqeAZSiKx8sOYmhsjg2fKfK7ADBu
BMgqvhPuBYqA6HBTyjJomMYd5pzFLeaDfRYt/wNunUGvWK2WW2cXvPEesMJLPj2KEkNY4Q9fr9IG
DqP41jnwW4vtm+SN2FuP/lRaC1IbE32gpeZaDbf0vkzlcwvLf8LR+DYHrMo551QCtbt9Rnr1Evk7
GQ/M0bAqOuOy95GXB2HqGhiPuU4HvABHvr6RwDDrY9fnPo95MCeeDXxu9t8UZFh1gNca/YeurUVJ
k1EefnMyvpD2pXeClFy7Vt8Xj6qcDD1tbrUCkLoCU2ECr9RM0PMgKwwtIk/7zKKN5v5FMKKyMNqL
jI9RedGA7ZGqPSwLyS4S+ryo7Gs/b5TMIM8Gvmv6GlR8eqNUaOfesOjBNzcVcEexE46xeCp1z6Gm
UdZHesExjYbShmiNLcrOAsUVqUPaegGhFzf7cTQjLmmFWNuzszWgP7+OjyGir8EtgzIwn3H7Mu7t
P9+OKEa29+6949BtAjqzBgx0+RYZtVDpBBEdfieuk1eVxrWlRRFVomaIgwyA8HU/Vgwsfs35Oo1+
ERoq4IOM4nwWVVqbMFnWTl+VbTmWDnIGbRkr8u6Jks9h16N4Li9mrf59cdetDIh46iKdK+MDpreC
hVN+ouHdpB/0wZkeGh1wdlFel0wv7TDKNlxSo4e8EIolcvQk4pP6pV92I6mCpgsH0S0GZ+/w/7h5
jgTPdYfHHu+fS8fTB9VtQNEHc0XIt1GadurvTm9lZ4f9aqGubgDWk8nNLL5c602mH+Oh7dbidPQs
VZbebjwi5cYdKZ/MyIPtjhRFC2mae5D1oGMptrwjknCq9gCjt3XT9Jup5NAczeOa+l59Ffj+UkI3
b2ml/iZjfYkv4RxbJBTXJKbwR6X3YfIyKY91eauajFKv0G9PaadTioOrtXjQHIqi8zyKGx7N7ORH
qvsnpNwpdu2Bvzv4WytqDUVS6F5LfuC6qYs1xAsMiEKbMlgVp2qV8yEIUusVxMQP8xUGOw9rHDun
CBed821b4pS5GoGJinG7zyfvSff9YJVp+8AsKGfDPOLdcwszt6e89M122iGGiih3n4iMsXJqJLAZ
nT/B3Ri7YNFSx53E7qebeLbvgQwLi/ZdgtdizrPkli80c8EP9t7GMwqf5nBpsKJ4zFYjS1S+X/cn
DPVBp1JCk/M5wh72D/x12OFSM6ECcRuDHMgiAExGGMQid0iRnAlIWi2uCojBzkawzdmopmqI79XL
Ch5EAo1/6s6HXFNX4xEoC5neDTwHXPqR/XWoWZfkABeRJxBDhWGH4QZ43J5vqGY5MJ3WiITVCliy
puEvX7eJ18bo7rigz5SJlXCRPYAZ9zoNDpUfsBA7mnuaFrqqzo8WAGysR8FsHTAAz4AIj7Ms1dvK
iHxe8iQM+LKCIhm/41ha1Uv0ZXw584A44OE7WmchrOy8+12Lv+K9KDsfx504J6//UFhjhJ3sLu0o
GYM/1iDq4z8o8jlaFJKKfkoI5jImmtpUY3hiKaHCv4U5UuuGzV0UQsxnpt9qApN4yIi+WFNEVYwq
L7W3+mbtR589ahFp15q+6cQjBSxf7JGwLjOwskwameIqRKIBl4Jhn+huFpo5I2DV8DZTxXCCyH26
4Gv/uYkMs8NiHvGRfDmvCRL7D+T1AwMaJdEPvkAM1JAVRrvC+zS1edPKBTndIpbZ3rMdmdiMn+Os
DY/or8J/ziU1thx3CJWiXIKsGDcCAAmt/cerAwH7TDX857C/94lViOozqWryJBVpNCrLqRWr436m
hN3k81hF4gGCLHLzrTcw9V6zNHLD/+gHP1OLe7wQaKGXQ7WUCtjcnV1ormgcSQFgwrxbh3O02DRp
wO7ELvBICZbLQxByr2sgi02rGL2L0YmC9v6R9ul07W5FY1KE6N8kcuZBg5M9tElK2jgMzzJRU+hy
L2e0obRYuybFHlE/U9qbFS6/Ig9leQGuQDWRDqIKP7do8UOrmCoZ4a7iHQ1xduxi8GH4n9rmSi6Z
6W8dP5y5Ysdth+8usNHYuYM59lseug+o441ys0y1SNmyIQGJu4E9eXWGwGICrEwnbJtJHQlT/e81
ldJQttERQ4sjhYTi/L45U8HJT3Qaa8OLDey2Jy6SNbQ70DH2hNs4lFF3/jj1RSgZlMrcBd4OCk61
5JnLqxwOQqzuQzgMFyAR3JlBycy7Gux9JdoA0YzGIAMTDDdr1MjVAFZ+rUlZtT4pHjEpcWt/0uLd
Kr6msfTqKm0Swhzdd7hEyUrjBsc/uoiZTS4yhXntdPUoBLdbYTpASvQAbV+eA4wvJDEoQWhCkq5t
z792d/0Bu1esRUru9OhFq2QJg35WUwtvjklV6Cc+HsWbNgEXZjeJNLdlaXkcBtaREB9xpJaKpUIK
2n38sUOE4XrW7Vdc5Yc17LpWgxMd0m02HYMULTbDIShVgw8zgB7XzIzLv2eNpPaSuFDgH9vvUQ6C
l7wl1TpQI1r4k52tNDVAWom5oKjZZeVQ+ap5KhLf7CkGCvUl9EmWSANmPBEs7lQOstUUSFBNHrCN
yZmd/Dv2eBrQTfw0uDFB1MRCHLQtYeOeNyGI0FjJLJje8YyoUtFsR8LnAW4S+maQ23PD8nCkhAxW
aXv8zOX2X/hYFBAttyqkE5zntjlzRvzN149lWaJpfWLqI4plqRvvYaXXPTUQXGdaX6e+wa2/ooL3
5No4DjW64sJqOE0pVSD10x6E8+QmnHHBl4mcYISkhnBrX6ETX6i0BfXa5+ncSgsSBO4rbFfjmhrr
n28kQ29da8L94scGgvt5Gsbwq5RScW1FvnlYSOQiOQ0dWL0hC7056c5sC99uMfZcR4qRWT+uZJvP
yjgH/bySjEWsGaPEgL1I/vtcyiDfR3lLTogTMFYty+rreHQbBYg+3/Xk/Njo1q9Y0EfK1uy2Mpei
oS2xwi2TEzJ8J3zHyvcx4rOLI12m9+lbrjfmqzFPOFSCUBoR4Z41JnJMKQ3aIoy837PCIcL4L/N7
hntsc/os3fgDurKr5bTKcS1tfMbDu5rI4eu+TXtFXyKAMfJUKeTraGaP8IVtqYjJ52Zz6IgzwAd7
sl0ixt1WTzGhxgkBja/rOzrk/T39nRIRU26zt96tCLmoPvCg//R3OGmae3dj9iYcgu26fx/iZg/e
0a5vi8RcvyXdw/QhMxe6VvegpvmqcL149WxvPUOyZvo7mJFviDurReIAfqL00DWJ3fFNhSY8Sn4S
Yo1slPi/qWcIIL4IiMGmbe3jUI2nEemkrNqsoAP8rovk4VzV3+NjWpDKUlnqYHjCJLOASYuYayYI
DjpB0iQqD8qp7p/+2IN799+GYJ40HRMSAtK+gZG68OoA5arto6Lsyli8e8//LT6LqynkdAlwuqG0
oGRtwdUvo702EdhjFZezp8kVyYhna+pKs+r5x1GTKcn0xxN5XAWqbvZmvbwsc+p2cMUpQDvGG/IR
4eElWNW/4RJIR/AHSU/uTokgrEEgwv2m43IPBC6vcgAwmXmfOO15GMRfAKBG4oI8HAadV7rOGetH
B0P5aWPrh/C3yaF6hkcGdW1a4JiJVY2x5SgJ4gjqCpm1kyDf+zXludwvz8WwN93ll6Q1nb+MvR9k
AcenDgJGKgrrPph/LEXcTZFSFExa5CwoDMFY6S4EEmb8rhYcu5J/t/riPO3MFakhL1qS6k3UFs36
jR0Y/tplJ2HrW1cUM1ZCPuGsAnI2lyFE/WKqNVrZG7LpBhbxOs2rZPj6+vk/NLtdSHzssJcLPOoc
6qcTQilRhDgkyyJ09sZJLIhain+DEv6HzjbWrPKCagDw2eVA1RYLwIChbW5c5CDDYdBVg58XilFq
kn+F5s+y2NkyT5o0/lkil6Lgv6DI1ly/WZx7V040ckxrYC6RMavE2NifbRLLWUOgReUmSlsTUbtP
tsS5JUACUdvtweHsHr7V8oZ4BoxBrGVTbIh4rVb7LOGdjhsD+3BjvBuoRm0yu76OWtYhTdBM1+Mh
74RDh7hckTT1k42a8C8dP+b7GAq/mLHHw8qw4s5hP+3p3WfdtWcvZ4hwomPi2sIki6G4M6aM/q2+
XFi8wR++vDSwZKPsX8CaFebxQ2lBTig616ZcIa5812D3NIHvJ8F544fzSTwmJVOJFepSZ4v64C3D
07ZRWYOZXCycId6CekFnB1mScRgrtzpC38OLM+niYmssYQU3tdAo3W2/h4E6Y2xfasEEMbmLvwSk
wDqt+4mYdfuL/XWF8+4rxo7ieDMxyLPqSjoQIEyeLEZFRkOLPGhaYqIpgoJIIDkd+0d42gf5NYa7
O6CHmAlV0ithiuAUudrL7MoUeagXvit5x0j9GxMwXxi/TKTMfJpLl+sPGHUbL8UwOeoJUA7Zygvu
1YWkBrJqEpH35TgnIOJT/3hbO7yJ0fboQMxS4DzRKk4Q9Mmdvji3Zqpqn94cksgldJLNm3w8oH3f
lVOtQILYCTFSJQMjQ5XIG4/GAZYC+rhdRwa35eUGp+w615/b4qxkj44aThDt0iKwFSPf2ksG0I19
NiBR35Tj2s8U0XT6b+Lm92RBhGUE5hfjzhKZLY5B68z2jP0fBkddI8HzanndtE9/lW/vmI7WAWDo
c9/kGOUdW6q24ICO3laoWzYdobyfVwy8F2dFEK/VObzNGk7RP2JX77hmiwrr/07z2leUC6gSFl9l
5sAvQ8MU6p50U+MCLgnP4aiDEbT8n6YN2C7/stkNl57xX7VrwfeROez301kDFrYgV1/EtRpgRkt3
0c2a6PIDiSaW6BbyWmzIFd2vaw4ZYO4kjlfzb8lufXWGa73FIX7APdyinn2ZLx79Q4TZAzCsbnuN
h07f+uIqBMbgSz7m6RXcVwWXfzLxY1KAPAMxXLYGkv4Bs8ELRS3LD9rMwK/zzfzpm3kvVzqcHBFI
mwUYvaBAw0YDihE4fPQkrlmcoxEcFDmtLiBaffJodQEUnE2tbz6demw/LludK3pP7+0+L5TOxbK9
VvrNDYlzpwPVIzUSSiFcJgJkd+OMnfJiO9kp58Njazwv7eds+exN1IHqnn2cvtfiov9WSUybxEdD
z7nNm8OjkFBco8JSsha/QBg8F86tW6/JbunCS9pwKj9+SuvwEmlv+klNvJQx+F9mHOPI8KP/lZyF
yuHIcNTVrA+8Qq5FF810ctPUi0+cb/fDCG3po7djL0OsGyf+8Er8aTbQEjg71Zl8xF9HqkXEy7aa
xD820ThvT9dF49f/8EwwpBhqjbfKglmQyBN7VYybSjIunmAHvpZveHPJUEtUeI92R+D2sy7oFnrb
R9tW3tevkRsHbLo9r8EDCRuAJ0HB2H3Q5d1L/QmGNFhdbDRbUCre1ruTma9ZotJyog3KwKJvH/Rx
aUZAIJzOHvhfQNBysbCZ7SbomLVUpRsOc1lpZn+aeN91WE/jdqHPAICXo+yqcKrKMa595m+dthMg
B/2lHLSgy8KRhRQb8zAdxt9t12yXk+Pyr7+60LYcLKLNoItxi4DDQN7ZFcz6S3xsImp74cWWhj/s
CLUHmwTzsZ6cDbyDptIeErPwpW2CJkaWzyfuF7QfQoVoGxTSjvac62SyVp5xqJD7nzhDwmgFb7bz
/CSFZzYLQFVe+Dkgfdne8P+rlPdALMj6h44rHo5JSMFMBN8FjwkcKxwKm8SbCdox8c7BfbboSEMe
asMJjHz0oe7vUKd/nVNCUnCrTUMBWERt4VxVLUYLp7EINJ7n1ozE3pvHX2IzG5NNlWxC2XyT+cob
94Sl4gczRII4fTTIOwTz+HPQMObRRdKEti6Vq0WxRKi4/2FFAkvd3uPGhwjEHV+jBpS04iuN1cra
XsAvT+iuZYpjanHyr1/NRIjbW4k64htUTgeVvKQA4v6Y+6WYv2W+Qd5I/YVdUUf9IBVU3g73qZkB
QuwBum5jISqfis5DCcx6JWmkwv5FAWnV/bO+7gbhdHIX56p4YrRCcj9IKjHadXTECUgc7086TiT1
9j+cysFzLnjTwx28/n0NMyCckdJ69a53OuZ2+BacRh7ilom+R5v3w89WxUyOQM2LGag5DNs+8F9B
VYfEVo9KJgPixTE4J1eyVW8aMuCHVERebrKvTclAIuj2OR/AndKhhfjPFlx3YniAq9wdL6E74KUQ
9JaH1I8a7zLlIFM48IzRGQAdhihypGMjT0kAXQSa0j3VBrvVF0jErEYh7ooslmvrAR6e0f0CIPuY
g7qW8ZXVsrnsavtwMLytHnwhxCMJN0JrE94I7QPFrmI3Wxw7ipd1N7/tHFxIlI8K2UayieC6uokz
VtXUbcHxu7bqVJGOIiNifhYiSfOnuC8JUUeHzOh1JEb00rzCZ/nwQ7vZKVSMckAoAa1mpqK0rRTP
3ezABjPdnjQ5R2d3yUAk2OqnT1C5p02i6KJhDDFfrhGfbBKsrwWNjjFIfA0a1P/dhiBgZ1DSZJke
ya+DvYPkTJtR2rYRaUEsey2U1Zgkww4jFTZ/XLh3V/6KrQgWOdvelf2ycm6bSpEiv3JLWdJJyvjv
nQQqgbObOE8j2PEJlDvBy7HwWy1AyNZClkkRCDlDLfZWUBozRULq5NtauWgmVeAWHUUf4101BtXU
By1AOSPMdkWmdqVupMydtaf4/oDI0uQxel3FnIYWvTIW+BKLSL7YJfi3q+6UJj7FRJsYzz/1iT3Q
YTMJotUc5oNpmmX9rUCm/iryvHAA/1ZtnFxU+maShWW0s5XSP3NyG8VQvC0/hQuSHKacG1xIcyfl
c2JPxzOk2WygharZ9oV8Mx6ErUfltsTTSAy8Ips4VFctViNt3I1uz89tKmVQ6Ov3dnFcHXgc11oD
bP0Im50oCKuk8mO+3LcDjcRvzTpRuq1mT8q3mgsiH/7W6Cmgo1HW247+BZfYfwBqwU8AZB7TAGvS
YRpIoBG/53Pv+hg86QAFbO2t3XouP+3yG5Rd+Jg4tX98EF3alHbsbjpENjU0F0d+JcHC7APAcTgu
9SjU+9/kQo4keByNeNeL1Iur0U664X4cUK0sP3cx0/fPC7sqZCksGt+5bIa//Q0pizKxQYZNuzbO
Muq8l/BKsHyHDns3q4IL8GLekb8rLMxEcnC52+h2e3VIItzPxRWo9nzo1FiJ/ixhRc6SNNxbcKyd
n1s0dy44pxKNSA7k2hrRwFBug97SSrRnL5kO1uENY8XkhRd4fzJuUKP4yWjtTqIEj+NeJoaa5edu
0DxHpZwLXT+4I31VBWSLvLnZr9zmDIK1SQ20bhXmtOJ/tcVsjVoMahROycQav8kjfedvt7ckuR3j
jVHOXxi35oY23IryD1+B1nmXyzXDi3O/90+qBOHmfNrKFr9jzXGQZSPDY0JxwA/+m4MRoDqqjPq2
X+Ryc03uJpdzshRtcJZ0VySxlSSnY/myf2xxvbsxYRBUEvK6N8lQUpZ18N+3p+MX+1XpyvMYyK+R
IaTFEv99dzR00pNl5/b92VA3Bhr/y1WtiEp28XRi4T8BeJrG7mflVXoWTGOven4su8DaO3YPvgAM
wK8VULJf2y7BasQHvLq936x9NcIuQM+c9tLu1zZ9mCRVNT0rX1RMuncAQZtmPun+utUCu3zSujYH
kzMexot0X8pjsO0qbhJ4Y0uHU3+d7DAmaXERuyz596wYYQQaRWFk3AWMnWebX7PtktGP2RxniOVD
lfHqIYosHGsNtbUiND6g1iTTdOPMdC30jJip0NFsWUb+iN4RpLKGFoe0aLiPUBKlW8x5d4s04FCO
6Sopj22mh8iDnN3aGICc2PLgIM3+Dw/1Q3OVyAa1L6AYk6r7sV0Cv/MYzyyCIZEgUqVxJHaSeKAG
jOIfYW8qIhkzkFd2wmRaGXpNnNeN4lqQtRFhcA8wlqJm7V7BKCBzKGBU7tdHItBiEwQWr3Q4iMwi
AcPi3ZLPrV/Y/gvfPTxFRyzPEi5efn5vjJWvrNWO+m5yrHFNN3O0fSOgaJvmZu6mYTyFzNe8xPW9
hhSFBGYxvKRl2T/cd+VeEHWJupiLU4fCu0LABHA3RUfD9EiB80CUdU+r51UgYa9Ppscl4D3w1pMP
Ll/sU/6Q3sx/wzVtc/FbC0QPCCTwN1sBQrz/IOIfBo3vka2RKjwxV0h9y2B+v66klY1+xb5QN7JL
YMXXLfNvettXcBvbrrfhQL9qNcTAw0CizQXHdWWwkJVuTY8JyunQQEdEOsbqb/zxvQkOPw1/GDgi
kaCRDI3jdOypt9RvRkHA4IfJvQlHvk0q+MuwIqc3Ms5L0RSTHvy+oau8z1Z1McCP05FfQY4DftQ1
M7PKtujHYEQu11nhF2XZhqNXVDVE3s9Dh6hhnPJ4qeqWV1qcgHqqpcq3bk02Ju7/Zf6vlTaImOm9
tIPRWwGGQPdrIgxgR30C57oOv8snPzXMrbUpsTeFnqMIDNb+Cfz0Q6mRuuyMvIE/4wc45p1XTvH3
QWAmggSwGLet+U+lPxcH21T7XTd/5KMf2yMwN1tvDJspEcYf2oqeYp6PfVjwZaB9rzT+Whze5fqb
bDFAti1+SS/7BYbZlOyq2JsCYsmS/4tMemU6NrhkFjr6fmgmXPqgqYRju0VCUGPJHygBuxDTvvfc
iVmmE6ZwqYF4IgBaUyus5IEtdja+dnIjlDwo2Fn/4e+t9N/amW89hxGtW5kuSo1KLOG+X+eDpbJM
rxedDjs+PH2+Lz8c41T7gFinQyec4rw81gUhVOSOTKCAJ7Dnb2Qfck5Tr3fLDTkUmbDxM+M2HN1z
UyPzjihTFa9Z6/g4yVVRZVdDm5PLE8YRFlRi24al3IF+rwg4+mh3udM4kwICDZUFJAI4/CvhL4lL
CWyr33oJz6KoaHrkOUwTcMVjNMF3eal0Xhh3PTDuDFVYlFBlDj9WHdX+GMon6SeYir3GDuGY1nnU
Ixl0njvYwMs0ZJRwKnonsUnlIU48vT9yKcnbO7v7DDmLwXGtQxjB7yYesJo8DUwDs7HAwnGDi6Ob
pc0/msPp616m6rkDNpDsc1pkoD3DD++ZC80nhLqCRvDI4BU7+xms3cUQTNCi7T+cXyNHn9z+4JpM
UdUg4+1Gk4sYPBE5Nfkgs5/0aEjqjzZ1iwO8+PLVLZk7DwURc4AeqbnQ2kuXMFyYHt8KA8gbxp/m
5x1ZLwk3pMWT9EzP+PCgEBBTFHGA7s763bZOxdS38lDGctgG9Da+5wSzyTlPOLCmBNYRKENUMG8Q
HVH8QGPXaR2TB6SjGvGzyq4luZ/baTOH6+SCC+0XYf5dpBfag74dYeacTHeC8EgeR3m6BIK/VP2K
dV1S3IPCZDcPJwysMQBBls4yghJ422RZR4UrJgftUe6EK/jWlK1oi447OwF21GI/7pFWdDjDEbFe
DxDnxS5mx4ac4iMDmG2JckeaF9VsWzvoQZjBUKjr79KlmuwaFSr0/HkbC+7nFdKCLoNDfmHiXbWX
mnCxA4uo0HzB8fUzJ5G1/vd1WhKYxk6z8QgyVeioFH7eW0YtA9PjYn8e6NvNbFlcdgEQ7MXZgUVS
4FBAI+WWmBmNkFmTenKNrrapMmrqDsJRcENDwc09mp53cZBhX3LkNtgYGOjy00y7U6X1kVf/NGoD
WGzgD4J2Ea7OZ6fIT4QCpDsZO2CVcCUYnxY1KSUIDFUzG9syX/K6xrUzD/MUnMQew2dzkBayJYCO
fWvySVtpZpvPhkhdWnlIoDELumkedMEroMpJaNaKTxAO64z0lscezsKPnovAe/Zkp3VVKCw8Y/U/
i76El3g55xgIqK5GS05vEJhkAHsGJd9UWy/LERqv+W/jwDFODirXru6dvp56GGyKp820UnjM/inp
9oMRZSBxL5Zn/mHS5/acbQOUhew68gcpC/fXVW7OMawgf/kYTE4zymw78sjVUlsxZ2ZYupd6ArPt
4OdNzUoZ466LWXQMUrN1y8JovahA7wPaxYENr52cHtq+jxFtn4tpX6n51Kj7VFkJqLvrJ/8OBx5X
a+XZ/GwZbp9KO854Xk+UaqSnmUE0YTaT1iG51jUl+jE3L3XPQ/rF18YAlsojdPDAiTWB7D4GVIFJ
e7VNDiGNSdSM3UTtoYk1a3Cj6aUpIUuDs4v/9zctj3LDHDh9ZKCqnCWYzHq8XV+3Uq3eU/P7G+kJ
PsX1NIgIava9BtuUSV7T8BKCVJc7FTT3iOG2glpXmhDaocZvnBDKrTe0bIzGCdzY5twpZ4oyrYDF
CRAIGhSa15kkMq3EEiRTdW4FDmp7+whmr+dawSOtUpyHVcLZ9iyTFkhGp1g4vrzGvNt+mVqoZHnS
VZ4c2lsSgPjiyo/+D1EN39jjXX9Z72k7+xjaZHAB+Z6/wXAtpxM6Kt+cOxFJoe43Lr1kZezZ2zXV
CAr8KpWHF15ez5RRGsvffRXFR01KCgozjkJChirkiuhWZhcf/j+PXZw1SqY+RglbxmyxyIN8sJ1x
0ukdWZ9EsncQlNO4X+IV0MSagpnWkzvHy//HKMkmIq6H5b6PeelgKVPafC5Dsd81ZFp0K2J4tYq+
YJJqJNW4yPBz2O6SiQvG/wCibFNu4XE8j6/orDbXad/Lre9fjVCfDE9y2V3jT7vdjBkngiQAaxr4
XZ7iJxNERa3Bp8t5UravuOhcR6qeIcEH9xFdeCWKkA8WcQ9ajO1Wltil7VDfwePs5yqfb7OqISu6
KJwtEs781SJKKcZM1BAd2IRYCnpVP+BYY71+5fU26kbexqy5MSwXYdmU2+YDhe0djx+aF4RNCgzm
eYt74xHKHXgjLIhOxJTBqu6Q5XdwnpU705tysrMcRwkF+K+0lEt9vBFvi3Ik7cegFNnWL1JMXsOg
JIhA+n3MVvsoYm2xbncWABcxPDKUFB9/917F8kxDCJ55wqSNdyn0umALdmi74bFNvJGeoti67FQB
fcEKrtkug13/UcrH3MdklDEvjaEE8K6gxKe7xlFJ7oQY1JmlIVJbOLEHioL1rO2000x2LvB5d55o
LwMZ9TVPsktQu8+rzTR2egAG3GqREIkyfvcO+l9oLspjSPaXZkQDkVby7na3A23rBsFrbYKzbA/3
PjzA0xzjp4JTy3GX6w3cls/p9xfKdrJ9TA+3oiHS+S/KWYPeZLz0EHZJJPZrnnuqmiGUyPVqTY+S
EzKwZEhwHrwGjaaatjFX6bIvQLzTRMsbq5jQJLErOtsPuYukObSv2OCNltCrtQHIZ4an0ywKhG9F
JM7quZpekwd8dT/4UV7u8vk82dE3dOXXJ5wncFlJPChlmtZaPVeIM8BV180hi9Rl/IxrsQxTmTXe
U9Bm4TO3U/43l9ZxYg7hCgzifvOqbruyNkMc8iesWbjEt77qL8xd47cz43Ao2SCs8A1+pyrWBDgQ
9P5davgeJ70s/rQ6/TTY+QGx9h58vJg6unAqx8StIRBbqv5p+R9peKrp22WbBdVlKjoxiaaVcumO
fYke0Zd0rLPGTvKp0TAB+ES54q8ykCSSUsoTnm8cpubDuGDdO7BulEJwiujlIKL1gg7CVhYR15fS
IY1MCFxN2dKttePj+2I7xrY+RIDyWqyMrAMLCWgdJ0olFcmiJlMDNn5Dp7Kq2zMjCQjMNGlSt1Uo
fQJQ0LXPn79bgZ0QkU7vNR8UI0LUymuiwtZgrEvlBm0ENVkQHj9gtWFZnn7qlLSX9NMfJD0KU4DE
Zte7xc05ASb9GsbHofeoc8W9hhK8yVhC733lwpds/OGRlbpA2segwvNk6xvThKZOIULH524MT5/F
RT355S8bS3KjsrJPcbUBeQYDpiB6ilQg6vw+wQIiQzfQlkmUBd4gXYyzUmvo0BTTNB2V5Cl1OJJW
O3eUE48j0Y8XssA6Mz8y39Nvcc0SptdiCmTAdKikBLdR66U/vXnlAsNByK6TaSsYz5xakJhDs9Yc
M+6VdG7naoTzkOMW99KeBW+YZXuQRdgltH583VeQIvLbQ2odMitVYeUA3y7kyO6o3BUMZi4mtHox
a1BrtZu3JVPghAgrVeQN9ktNvcnONYgxqAaX0TZ2XT1zO5kVp0EiqAfIR2yZugzDyrwKlG9JcgZO
7d5snehSUzO/PnE7f97WcTkB61xe5Nf8TosHiNFCm1FxGVGhnX9mIWncmy3tRFy384mxJBh7GFL9
cw/S5b37DFT9rkhAeJwBCNheTEkoIKv9bgmk94H+lqKhkpmM49sGQ0WivfV6RZH/hSLVIq+nIWz5
N+xF3anbf516WfUzxGpibELUZj+txPN+akHrASqTJhCiC7iExBcBzdxVIpvSD3/ijmwOZL92KWSq
u06HYWkEyDWgurv7z3Em30NgotSZNmOrA/saLbwOLnzNNBci4v0Ii5sCrkrQv2cVPUVSQzVoYMNZ
aewY6TA8zupOHEcxm3Ou0jikyuN4zJof8Ayx23B++TAkylLRcNTzWS9YVZyIN1R2xsXSQX7TwH4s
CG90PWbCqJyobRFFl53UDEI5Y6QvagKBP2WUZDYyhHmW0D/wMI9VgDKimF5aF5KlE2KHnq1FNT9I
Al1ei1HVkTgsfPPwLW+Tm6GU6x+spT3RO+SZKxmKejXj/l+ZUluYvDpbPZcvmvJbR9j7X9qWjF6N
JDjfhKZikVgN28L2NJZv7OlyduvA36X+qmTEUrIDexDzKIPljEkKCOg8JtijFIXW7zZcCBxT2+2h
c5/wHZOSDmml54nQXeOzmDIwzvFoLAre+Pu4NKO51QvwzMg+1Fws60yY3D4Tc1nrBQ9BlznXn/xn
kcvmUbLj1/cjP1RP5erFQ1roXpjZRi85M74Id5DTIij+HFkESMKb4Ec+xAe1UM0+seOHY1YPtUwE
++cnPiSXjezONImiuQ37/6+EsBJfTy9H05yjoH0zRc67z1opn5DYVlvv4YXbmxS/35qgk3ZWWHwe
YOftL2qUoeuh43q1Z5zudsI/ISt8E/xQRb58BuWj4PRfhZtL6WCWAzZCGxhX1O07KXl/4kb3ZzxY
Y0k7jAj3tYViyU6nJNSG2JRNOdfQw3v33u7lO0Ray66IPefXwLdXck0aO+IshlD8B6NFYqQOHs6q
DkaEXlZL33WNAgggrxUET3EoaJqOD+FtmhrrkiMKxLwqx+2fW1zCuwNz510flWGj1Ty5ClTllN4N
AKqyClJR08d49x6m9kiqOUExPy/Gajx4rKVC3iepvcT8XXyuqNzzQNgHFOZ7UWampvb8aALpQ4bJ
/IkwHptBgHEa2iUzVk9my9HOo/pkKbT+mAqGgcrk00jv+Lv1XpRJLZdQlU3aBzjbYsES4LC/ijWL
KRyWa4D/UFO0WzenDe2H8y8qWyp6ijAvaDDMEmB6cdxAx8xKdeRK6NEr1vvs25Vg5fD2Zxx7CLkW
1np6PaNRB3/dM5PVtwi4XRwFnktn95WgxmNie4/IFlj8u3jbNTcOS5rpAAw2qvSErKuuCIq9XZP2
SjCV3CG22AksCm2t0S3H0JhOHiDZbsxvWNK1anCX3WTEIZ76GzEQIihL4JSxbn+7gZyPhE+jQFTu
AWrNKtO3UpCs0i5sfzDuYoAxNBMc8QpcpT0wEriCTHjmu+WS1G47Q+lPl524K4f5P1sUDxnR6k3r
czuCuiqrDGnoaIOTCGDM/Fhb27Hy24YMoRzQtkJaL2yerLIbhQSkH9QJDrbeAElAfFs6B4MsBNUz
MrNKQgJP1Q4s4Gkz1HO2+oWRCxtvQp6u6Ix9Uul7zXR8Csrxqc782NTZvCgpqYxUcoIvwQdeaao3
V6cdPlEB48uq1ziJh4nnPEBHJZ+zobzgGNj2zZxxktV514AMkOXbO1vOJi1+V3ClL5EuOy2Ktw6w
qPyqhC5IU2GS6aqXUcMylH12J1GPvy0lVHDGGb5OyE2jDxtxFxANQJPvqIORMdEHvuqOszn0DiCL
vamc1kClTDpRoxQkLySi4+zK9wHg0iTXMbkMazzJ1cDxSRvCk0PWE7cw8c6sq0F81z3qtrUA/mao
ev271M8oy+IJ8WL/r4OXTrGg4lSIIAV2+yQG9RiHDnxrjjlwahe5EQvC7v810Gqxfdt8EtNtPBmx
1TfFibTlVU64tIIhlSB3wrq+HxXQ+R329vY56ofDXsg92+9AzKPo0b/M/NF7Kf5KkSBPcmBMN+SQ
HiPsEsnmbuUS2SQt3iws9Ols6HgCSf/pPowmaiwNqTk3sRpcYyWgJi/MGGF32/7DyCkZA8mbGDki
5Yj45VNkp0Mn8+IMcJIZODR3HbAMITT9hcuRyZzqejrz+GGDR9v7796NPcP100pgDNO5dofAVIZ1
ewXQ2qa7E7n48ZPMzB0jvTQTMa4YiLEP/8wscgjhzaWvJgY/A4ItGErSj5HEKmW3JVigLSoh18Y/
ZGGBd+geRzbxglz8OTdaRWRbOsw4Yh/brsv5Y9L8sMRZpxUbg6RsT3MDAH3HYg3zlVf3xkpfx2jw
CFuAlbu4g6Dq33QlXamsdp51Bw7rWkp+JWgm5uaRRRjoYw9mwfmo1c4F9Jb9hGCossBKUoCbOHzY
tXd/+zrbCCgajPFzUJljmIoB9MFG4wTa9vF1jVsnWnOKJ0ZGEeHfzTWXOSNeyZptabAIiXul9xke
6fDnJeuRvkzNU0N1tYYV5BBPS8JoF5LPk1n9A1KtvGXi3cr9A8uWclEh17stKZi0JsbWprzCE9J3
I6OCUyJhC9dvjjz2vpXSZvqHc4D24gJCcAHEYYHxDpBOFbY/I4XQwNqdhXl9ZR2A/EBT6CdXsWhw
cf7TacIitdQ+Y83eTeQkd589O4CeUCOrpQgAEN0gkRwTq6iCaAWrL/UEi5wheTmSZmsyPbiAwvg0
PAh8mrmGckkVXLW1CPx914yMdrGv1qJkLRV4v1zh9O7wY5csPWpu21zDWQAhZCQUeU3uCiGRbydW
7/QPUyVQPX69mZzszbHwn58+L/mK+P3owQdhD9W4EMvEmFHcycD0SJu6cG8DgB5zTsB4bnZXXpHA
tRQPJ6+H2CZ3pqyHz5u22vp5qO2wJlNjbyvaEJFiL4lpdOAuVTwm9wIVFGflzzX/d5a7/Bf8u7Ph
CWcMsbNpIW69n6twXvrBbyRNPOgw2GPMj2Ud6/lb8iOTsbGq20N+KurISlQUTEfPZJ2KzvIfpTa4
EjdfuiOcRUMlO5fxirI2HqNGMB2TgMiqac4/4pfELC7SwNxxo7GgoYRg6WbjL3pd+D7DOQK94DGr
E5NOl7mW79TnPIqb2vizHze3zbP2uaMeIKfSxCo4oKjtdtjrboEW7EBTCIaPdWRHd5qSvPgouk4P
PTukMN2WyC5qhxu6EPz7oz8cKOTTSewNz6BGsuSftGyjTMDoi+eWEjaw7uO+hQZ7pDuKmPpbF9d2
cwsD6NykVccc+CaYldKQLvUZypHSC+sAyxuKPn/+hEgjwz0DoDxe+pIusXccwr/t1iHOn1t8mTAI
/iRSTR9td+DvBtKosMQxmSa98BZEQtj8Xs0Xzy/HU2gdsboTh1/7TrbRqJ43vrLc4QYPeQK6wGK1
ufmVN9b3LNee7Zx9yGP23jef9Hxvakbz9Qu2v6yAftq8rgzXDCIy6FXPU+ZFMvy44vna4ZL1AlY9
rbzA74HXTcXOtKacC3xtmYM0XaR89mCSz/pEBKRgAJZMwtythLX039X5zUypSMHbPD3cZBiLyn3Q
NynWjDoeJlDyCo/6YH68/IYaQH1zo9RAfLzKcUvyjmBoUbVLP375ntlbvvUmt7jjFwxRadLfKLa3
m7EiHpa6xCAqYQVeTNcDZEMQsVEQG78qsGWWUZ6X1BnP2+ZJLnwepKr+nLK4CL9uhkjW0/tV81h0
NOkEAjyYJXZaRaR2dE3HvlpzK4g7g6McO/iirsJefY/gpk0sRyhswByi+jBstOwXh6K6J3vS/J04
efAjH1amhtPO2tL3gghN0U4d5uPhevqCMdLqJOQIrnIvvdbR78xZgllmcrIeUGV2hac34+Q6JkwW
jaTHBwpgmG8rpNHr5xL/xrbbPZpWCSLI0Y/JujJa8M28RkM0bMByvQlNd7tYC9PuaeMGqWfr/1JV
pkhmGw5nwFdmiA9upXR4FO9HJZogYPYP3LkG+RuY8ci6qocyJeOhx6dwk49zrFULMflBTPVj9446
O16tFrPED24gPcXDhaaAm5LhGtCXF2IMoTxuMd1Cn4XsK69tR3FlXrLUIiSrRch7c7H8LQmUDGR5
yqK/OljkZ0KhINg8hBqPfgbN90CrkcSphVhYG2DCB6je7HucegPPFnpnWmARsvFXyOH6ClEOSp1o
doS12EsEcBy9Q/3IfsKuAaQ3Nu8YN0IULnY94mb4N6ppYvJNeDZo8zIHu+mB0GHls7wNKs18MFYL
1eS3E0Ov2Imxd8hhpB3+NNLezyUBiIlzvH2zuc/1jT31chqFnr9NfBeODzUysyFrPY7JwaWUVFYj
+vcf330qH3Rkmyz6xdM3guV1XPMxqbNVOn8pTbhEhLsaDOgFYZr7TjrlQGshZP/8q4aXNm3q+npZ
zsvd8/gW9eIEknsgyVJgIH8OREYdcdShyiqlv0si0ZBceZk2Y7eabYEaSW1QCFEajkKgWu86aCJU
kz0rMjgZry0/EKRZmDrI03blKkmi7vT8wh2iDUjcd6HhAg9g2KNYc5B2yOtgXD6s5m+16bTUTlgA
xZq8YD1B7fqkOPeXHBsiviHqMI1SiAY5rX3B/hhzyuSBW3RG1J0R6wzV9Li7v29fHYR4HFZR/0h1
TCU9Ew5BSG1TrsQ9YeLMLKKAurr0nIsXeAce6caolBMPB1DvFN4bs8UYsojMsKyltI46w/f6wzOo
xN/mM0kJQlqoHAeM2Y7oMcAHmOmhE6I+PotvFThCVHb9xoPkjiOZtThbKyv3HzqQurYFhNUh+PGv
HviHYEP7Tnfz5amCRyVAXQfMAkRh175hL9YAx4jkufvMr3u8Sf/C4JlAEPbPyi2ZD5JB7GAgZgLn
1Bk5p+IAWmgiC6jZtdMVDk0ebVXLWmCVwnCLxxtP1Z5eIEPghzj2m4RC2C9VBp3WK7MYvRrU33fA
qZX6KNzjixBFWURA1rxjSi+HWNv8k+ige5EvglHq5Xod5ZSTVlB4CUG0ryWF/UdaXlIhURy+fREr
4RLpwqmlOBdxGrNju+c2MShMiZ6psza6ckg54uypVkkG5dMGDir7ROOKt1VisguJHGredBHQOTkd
TEe4uRIVD+uSg9oQGafcyt2QXwedUzYUhRi90aTLM0tzzejSKuqlCtwFKOivxjyIUsiAzL4+JMyR
J8Uy2LFDx3AMp4VKvLRrGrtiISLdr4iJwd06V0ifOhUhsfpjTHhip+jPGQSo4u5GTnpWu9mnvG8D
9KavUVsDQ02jmPhESjHp5UW+wK7fX/X+hva6XkolUkqGW1X/W3xyVm5PHc6YXOd1uuGbfPwHsofX
wEoYw73PqUO8mPzrdB/eib0bAZSuRujtQaBBy3DQ62rApETWgDwWheuFv7JwoPekEhyDuHDBtcAQ
SZy23izs7zX8cWrGq3BRk3RoBko/tbo52UK1ZtDuLgNG1iflMizP+9j1QkiAorkiWq+S6ZgJj4cY
S1mOnYAIpnqRfx4u1EgSpNLh7UUU9rPyBxIl8dkN4rlO73E+OHpxCX6nRWM1bWUifFhwok3YJMPh
6S6lMEAEfTmN8x+reGPz4iCfDo4MOp0WLSqetY3CcGYchGh6uU6A/CVLCXOlmOBD5YWdXZBnQhLA
IkzzuJtI4AwIEuYareqk7RWBJTU9arF6v0WrjOl1+tRLhBXKuFIjs5YKNqr9vopv0FQqeO7097S1
JhF8/Wr07UeejJv9nhLr8Sg2+kM5hNnCOhc5L4VbrZGVXF8HVcDmffpvac8DMRbDxwAqRE0gOf4j
ztqmD4vFwGb0Agn4pEc5ndwoai7D+2Cn9VNk9xplDh8BHvT3/59S5XlaN3QyTnDNxm8vr9PbbJOh
da5D2fPXmqXdR+hRxxy/76UVkexXijyvBKgSDSiLnRh4Lhs8ns0lsBNRiTupmYGmNzmN7A8lhvg3
LUQ/2l0t27ksytuvZDzIJ8aENbYK22Qr/Nus5uiee7uhneTVUcykcfpsrsvajcrxFS6Xt3KRHf9K
T4dxufbJsmPMi8v1vOkiAjotDA/NSojxAddvDt/+J8mhEd1W8C7UKdez36kSZM074jCn1w2oECBi
uONPtqNurWhk87Cd8NEDjj02F363nOqlOBqqvR/sGGAMQk4YVUEF9HU+SBnUUf8jPFKQi8080GcD
Nwz9bGoOaTQoldZ3pXFJ9ldeZB0gdRMHnyJpS1SL1N5LtuOnM0fQTlYFXKY9diIGOlWBTOZeKexT
Z4lZIxPtW7C1p/ADUVsH5uE8+ToP7kU+qHTPFwMuDzeHeGc2Zu7dFWvmfOt9RfLXuuon/KJmTgJZ
prLv3lefUqa/pFutyJT0zTx7ZQa7JJ4VFA9o7ZT3oUrks5hUGM1hdclRY7BztQ/hAUKi1Ii8WzzP
kgFEiSlVF+SCx6bI/KswCAHmAM/9Df7N8Ze9ctWbBY0aC9zQnnPOSmddtMmh8E6VVmQ7FGB6wVYy
ZG0AclVAYIYcAV3SY9dJoGw6l4tCj6hJGrqz247RbDWhCjlL/3s+Kf/ur0Cjn4pf/sW2ax/I0ci+
Gm9wcO9KLtekywPokjqOnFxU0SQrN+5rmF+zY3w1vizAVn0fiYWg6drk3C93zPKY58OuIU0hJePw
3rY+Hglj95IUYzty63WHi6zs7jgSp2KkJfVIgXy02SlpuTT2RJCGCbjGpojpawmpZX0eiD/ff9b7
XyJ9G+BPHcQrA3BqLqBLMquFshmvNAlPWZ0At3RSaJl2n6cJaw/NXSbdFCuQUwwMdshxE5Q2mzzO
rZErXAnkln4+ZOquKRPSDAioZW+vKP8DY0Nh0oHttbnBxUqr87yL/N0Ig4pP5zAbAWjxB5VPhF5X
nt1+ADuoiDUfWkY+Pc3shH3RDuI+Cbm5arxVhOXTZujX9NcWuNqv7KhNZw0TMQHEyxptqTUmaGmh
U3r4Kp+arrkiGaXZ+yoHDsnQx6QIrOHvs69vbc5HgUfEqwqTfeWxcAhs3b4+7qVfuZhAu2mNroq7
SVYfzrA+3dwDzFs3rtQjZrijCJWJ+6VYHI023+ZdVzE0V0PsvEYnbJWdFj9wucNmXdEgIcJDWM/7
qmUNbDumiIYTtcGViWPC5bT55te4l5w62YksHKGtk9hIKkKrpIgYCKXuOyetDOrzolCYaGi/boTL
fspSc959DbzSMKXREPaEfN7Ay9XCRgeiwWaEXhJkOZtojj+c31HqCCXMDgrYPmO5TQX1xlnCVjcs
y06NljeAD5zD7wUw7CTC/g5bwr4RKhp7128JJn7pAA61psWyw4zMuIJdRI6AByvhnwbzfodsZ7ea
+8/tKqadxF2q77fi7F3sUXs42V5Dop3zZQKZafgg4Kokl1IR7Ck9VXymCkBNyHMPX8QZMG5JnilU
bqVVeqwomesnk9KxGxbmAqjjKMebz4unJgsMjSsJ2F0nbu2cY1JkVcOH7LuDGpemLSen9ZZZLPQW
yU0cwu8ARB/Dj5i4TYmTN8+AU9jDftr/XxmQr2lRFjzy8MxKOq9DoaXudbmEptn6/GTWTyb//4zI
dh46Z+BCBeskQbX3Dv8GiTZOA6mKkkYTJVWSu1N0r8XLVIe+z6867TSeUQ8rNvwHg6XeFWqn2Xon
1INm09N6hK5+qVEObNrdt/5EcvcQFszsqwShiS2MIGRNt+SK0lCUDuOzG7icnrK4JfrEvQQkGpvw
/+MJhjEO66rKRnv8tiBa1Nw/mcqmxR967oNvOe2yzm8ZcQlSPCZsSAfbZCHw0JL8c0Pq60SmUmhy
x5N8uLV1jTVPgqAUVUDyVErF635NbFoYNmOeWGnaKV6cnmNbTe8S/yG6sK/p6c+NbBTXQBjktj1J
6VjFirseicVzc/tQWwMAVbpUIs0/1NUsJ9/yRFQ7Fw6KLTPWwS9o/2BkwLacjr/+EbSTAY17BcMZ
YVtaqAND2f+Km/X4yzrrRRgm0YpiolWVFNOKt+8jzaqLZNvi3Lh9RZVuas9QkliliavjXjPcAdJ/
2ysNuzwlZDDwfYl+h9XaQ2LI14CGg166ed87j3rt1owjU04lqiZYLhFfzoduxbNPmmmUKnGZaPDh
GoKi2JsARdJZ3hJY4B01hjC/uM9bI16yceJb+Kq9F1SLSrdDdih+zQ6WVqimsy6aec0G8q5Q7aXu
/DvQzQihlDgdHj5NBzGOytazrB1bFdY2PAJM901QKl92smchCBM2bf/nicV0SLSrFNFITcmqRl+c
lCx094e15XmPYbmN+PVx18MneiCEr2Vun2mqP6/XBdKKVR6Qcqyx30RwcQCRLPTO2fhmiSmrmhuG
jrWnCDpQUelHK3F6apHqvG0Edep8l2rc/qFduOt3uEp/fCykJMar9PEgrXr29sSaZvT4kjPhU5PQ
HhQw21PeogRD6YDjSoEldWl+kNiC/BEkKCO9eNA1Fe0nJTD96X3+kwJhXFfbK7DkHXzZxTEWoXv3
JicXucPkREpBED9yExfUK8o2bbdv3yLtbZ3Zh7Ru9RccERFvW/4OeHIwY2uA1wI3tllR8OUNoQBn
xBwYS+b+OOta6BZEMrECTxhvgPachTi6Da661S9wmO4uIxtDJYBuuvdJE6DI9aFN8kqKzn0/i18n
Tiu1snCYcwgQt3/SsW9rCDcMa2oHfdmHMv3UvgS4zwLM0/XJo76YQR/MfY3Ln5U3xfyYn0UQzmqv
Iqeu+VtggspwOFseZ+gJdpqTidFVSmBYFpOiqw+YlpW11+gN9leM4lBM72aWyvzozr665PJAxPsJ
p4VVaZcRUqDiqBTIK8OO2oegwL7UvLSAXUcA96hkPM2+GPB05y8+lhH1baBLqsLsWJjG/xDx8wM8
UQta141lqmhoS0YbOKlo9dJc/7bJI9W4jzx3OnT3LyotvWy2ZCPCWDc0tG3tYzAvcG3nGi7x+55+
MU9mFixkJI85xv4Xuay4uao6F4/6mKvWjDwsWbgAwxqpEpCrm+PIh9erD5gOKYYMkIA7qTr/dclE
oCYsQmVxZ0hYtACtEXju+rZM/O+8AAusukql15bY28ol7P8xIimcXz4z3DbuMdrjfe4TQKSZ0bq9
VIONzlSEO4D/mw4wXdIPPeW7pGFIIafAku4f/p0WnXw7/r5a4umSRtpdEl1ni/aF9cnBb9oZD8c9
+PRpQBSBTpeup3SRz7PT76WXBT2Sa5xAaek6LrRl458OGAePSg7LvIerjxl4RS5a6ASj2efGSHz6
6ps427RF7NtDjDYr7t7+hWytS63XVuur0afoL7ceVzFSpX6gu+nk11cK0sj6l9syIIC9tV4YvP0b
GaCPd47rUPMhTKFa/pOkGZ0o8J43t/5gZ4qJDS3W8LlN/Et2RiP5T0WsM6cyzidlEtyoVc8ntqQi
/xE36cDdl4eItp/QZM6hy9oiDqzlCI0i+lW7bLviin2BrVNYTmrj5uTAdI8CV9QiqDU9KDWgN5xN
Cw0qwryBQSx10KH1q8E3fdPMga3qpimRF6iAnjnFNnzWATzsKbTNWXZurW/E2/SboZUQsVKswUYS
Jr8sKfav10pSpvw12J6yfWyxZzNMXuwarfRokkRFilNINAWMVLsFNNY0truL67Or25w9Z4e8mAKN
kEd0NsFbIt+0qEClJ1OdaUCS4aQaGf5aAHovIwM0dNAs2P3Wq8ieurheEacLpFf1rCpfhxumC2dH
IpNy+oRxhhY/k9cE30iZS5TiubiEgVdVyvOf6kE+z1qaXLcZWzg/NDy840wsCsV4UmWoVve/Ys9V
key+UXSTf3H+eoqh9oaLvFEmai9ioGcvdcv8iTPc6TmbWWDhrE06sWyTBbL/3vWO1HPNcyGBd9tK
A2qRS3spoUkEdIJZaQdZ8I3mmd8qcwbO5lthxYuemxHtZnzcQHb1VLhOjO3KLameeNjw/MDthwf5
GJxCCpQe3v7qKkvRzJ47ai7dKwEbNVBBABHBTmvXHg2BfOZmaqfFLsBPCe9Q8iWiim4ZgodQsF8Y
4T7heO3rTSCIfsRKtFLhiozzPQ2LTBbhWRJR5N7fIm+Wvk7uhp4yp3muetah3Yh2AwQ3CAan3uDF
oTbiJNT9y+/3KLE4OU+PuCD77w/rmnjedpFn8dvTTNbN6oZnIMHCO1OdTVrBo9EvMBWrjGn35Nmz
H4lvk5M4ed8DEGDN+nduOV2dtGpbw6VD9Rq/sF+4fdljHYeIEy+41vGh5ZKRKTiSzyK6Hfs0JUzX
yMlUgfoXKsNE3NJWWblGzqc8LtJvB4QFzCJ/2OfniZU/HDJ0K6L3BYS47t9jWtsHkW16zeZ/Ifs4
ov23kfYFAm86OsYCpnfFPCfrUaLpPNcwZF7EXKRVzxhfJlWBvbpqZUBDUKsk6ifo2EoPZyIyD+NP
oLpNv6g8asrVUaTX8rieYeRA7lRH9MYvcXCxrqfUx8HADyyvz9n+A+QFjiUXkbkmlqStdTtlL22H
ksjEVrQ9AinInTBHJHCoTvr8+Rb75TExWf9PmbzegBUmARq+UlSOgOSInEdQ0JqaTfmY2yFZn3Rz
5hyBJ+dIJEPanMIVnK9OesosBogdlBM1fs6/YM50MiO0sLDCcpnd7RQ/ZYo6O0AKpcKKAS8Q0Piz
honmtw0JG5/S/US3sP1+jAGu6isiwm+PJNWGMjtHxNYFtmxkp75BdGVb1W2NTaApZYBeJJki/XD5
0U2y7yKDPedtfH2ctihx2+h02ft/UUpCQqKf5x8Wvnhw6RY46AMo8M4j+vZ+KTvOoXoG+m2fbzev
SG0179Stq8c1FtWHt/CbDM7BLpI/aveA58RHyAJskRKbYD3xnOldZikTjV6uBWJh+stPSW5fBSBw
hmOrEVMFIXRPZVh8CpycIlixVSs45XVFhRhXkQmHp5lQUfTsu9aw6bnVZDwzyBbcW8S/rE/D6iQA
Ph5/J9FRMAJLGqQ+g0CGn2t4GjW5BWD1LLWVfXGDsVci6ohYeQZsIxD3AkqK5kdb4xJ4zP3JPxp7
PSazjCBzYEeDbt8JpoAS2aT+cjKjQhmZ5oSkcmLn5/Gjt5RfSC4n4EcEM54/5r/TugvfcHbiaBdP
xM9qroVvxr6KlcDLX21RTuRA4rivPcH3Gt3JTktsrpBCqfnSFZTYdPTPCjh5TYIdHE/ZV+/sA12m
ZRmp12pb8AJnt1yWOoSmMbOfK+w9EDKJQTUIOSZiwLJfNQ2vAkOgHbGUiXbFQcLKND35CZ5or7rw
t8xOZAsUJTGIAQv5wRJo7TGD73O5iDzOCid7QZpPeyS3I95WKomdepXPWdrRdEiLuELcXtJPD9qs
QumelFsBlnxgPi2Z0e455BFlw9m2xbuu3sHflAvg35CMj5L5iq3VesFmGt/6shmLJthD4MWyWBVu
iGVs898J2UeVRu/fT6C5eKv2ItGeYcinajC7DAtIFQUvF+Olsy6j/axNN3x41CHrUSD6Zi2Ai5hD
gkVxjgwqgf0+6HppXtWBRX58IJB9ZehHk5ZvXms4MAD7+GTwzuJpL2gBtwSZh03rLiwYzkq7JTc8
Vt4z0bn/EsZQtLvQEp4/KoaREnHIuecNCRmtuOjqK5EztyKMv8mVaUDL5NCsSlN/afCu7RTH3grn
frlRKedVWe8B925HMQezlNYbKC2ar4y8M/cGyV1c5Bw4DGZ2tMtlYZJcwDt2+CnKL8IRikCl8rK0
eG2on0p1v5qbjOaUnZxQ8ltnz8w1MocUG6osocpwrEfF9l/e7XkIR6L3ni8W19krzQFQh1lbwfpH
CWJ+SyIf5GFIbhY/rIkoqMePq8NFr60TaoJpjXXFg/waaGkuhPIp4GxihvFZHNfMhhBkVo0MDOMq
ujFg/cVrFM6IeYZiSjgfIBIUgvBJU9OubprpiJCSAeAu51Vwyj21LF4f+MmWiqG4a2ox1VVvI2k4
9Wp2I20Cl8Dm0CjaTYyVgAm+f/9bN12MDE0doVQJALA543vNhyUkhopGa2s+e9yEWMzcKnGQI0DJ
uhVhOOMm0RscD7ZkcWWCB3nDLATJXRv3LEYsVSrmkT4V3EOPPg8pvwbWVFFOH9w4r2u0hYIVnIr1
/4WrtOBKkUb+fCUavWrNEl9h+YrmbVIjEreyvMkZKRHNBIyvTMlrDtQXMf3PNUS3aXnxzQvRoAHn
bpFt1vb6v44g9IwYA8kfSzDxalF0Vg5d0Nk72KSGyreI3Tqj9sbUXN/AwZKyUWbz0AVh5ay/Y3xa
0lDGSukCk0wxgyhRLAHQyj5SYy6gCyPNPvuvSZUP7pvfv3GknnZoisEr33mm59/3G5LZjp7ZwF4D
3LcGMmGrXQucyr/g5wnAtAKqyGiBwxEJDaSP7YsSDoxbzEGy6xafku+7J/7P1YbLbS06napiDMUm
cjags90RKZYlHcy6MtibrBe3hMTWeUTUBHBsGYEvGKH8BWTW6shfORhfOF+lhJog8AXFcxdu86t0
AVwnhV7lifPC8a45SuDIi9szoqy8qgOnTgRwHNLP/htvuC6k1wfZwQMNNKyqnzb9nnb49SldiZAi
6BCWhGyzSLpamtVCsZUHx+GQzxvI4grvC36CumyZVQxaRqdoCJlPGIZAvlps2+P6PV6Pubg7azLg
F/Rf12SeGrN2BKquhMAcmaTioU3/ck0YfdJstaKq9ESMUWvvQhhEnHNoe+lbtgWAJVAh1rsKo4hU
eKOxtd+QrvhsjmQmxzlpHSuTge08G622VkeQqFZPnJrqjQxlIdG5wLWa+aNkUfAy6rRrcQVUjUVd
N38mgH6tf8AK55Q+L2Tm5cz+ojZynK2GhhM64FxxFxBFZvwAXwSzAGCo+9glnqqv9T1VrkM6Lr50
cnMrpns5qZnxNgvK+gc95rRkCMSkKaYZuErrwRVnvLjqvBfgVnc421B4J81voyFaYooMQOS7gbdN
dSL2x5BfZhku7jvcBULJeWVnAz3DqnXnyk/wI4HF1H1qIYBD7DhwnF/ERDMPZegJPP1VJk6ESEKU
Zp5N5msBuTiA4tykQnshFWtnCIx02Kcb0XWdjG+ZVqnlxDDpYRPh/cq1tHEfqiC53FUYZVboPAVb
0C11KOj597jubXshtL+qDy7jBxDm9BrU0AMjb+PAJbLlZ8H2Lt0+CUkiBjJI5a0yPVKfEz+sTH0v
TJXUj7rFGKYb5z2BNJsEP3lp/fqOahU/TQKLMcmvgZ2Qe8W9AJ1Vj/UYMaUjTtzlqktqvJEFvjz9
niubzgkFp/tSW2CLweou6PZG4rCci68Eektvu1upx86AJvo3VCmhjbCysmIWw6KHI+iJ/V/tnhgX
uORiA3k8hZJansUEOcLckceDo+DWzRTZaHugLlhsMsHxA5HXSp6AdHDdckNSOZDlwNF0dUBo7Ywt
4Yz0EGj8IDJyel0J7AioaDyP8NLKNmZKWkRvPxH3X+MteFSSull6kabZydzqX01Ybu+F1aOEUeVS
5P++Ht538RKpf5Gl8x12ITXCSnDOP9R61yeHHc9I/GVQmVBfcsH7CcRgwbUwkz/iiijACL5Vrozn
qT+37na1sXLmXNwDOFHS0Tvs542WdZv1+PhHCU4/vxm33gfPk2P544ak87XsYT6KiaczWR7WGZjk
jQ5/3ytSr6yYoIbrMWJ1KuMzw/HRBD27JHXHO7Itdn8/iyrKxA62BbKYUD1dU1haX7ulCWPANQEr
IOHt8584NBBL2HdE7M498Dw8iHsRdHtD2/uHvhdxHM5PLbYFyeXCIXPb0gQf0oYWJD4ZqIY19lco
F9kCbqavd8u9av4dZECsavFIl4nuBNEQFWWOQqra+LsIM++51jp/EBxLlNh0ugKk5+fyyiSSNVF2
aGcAD+Z7DRv1V86fvTjKhksGWjN8V7zbn46MOmcXG0mwT1g1kvuTmPY3WreEQwB7rkTFk6ljEhQS
3DdOWPU+utKeccBAunqRrKLkOoYo+XoPZDTCKwHJ+ojcXu5AiXZMNEtNjF+IUQp7HETs2wFvQw5x
RbwtVKKUEhpmSOKmFTca1HsJsXEg5XXUz3IeZpHgSo4BpEMYdKgdXC/KX4H2uaRBszaGdlAB/7RX
zSyN3g2fax1eztk6gqyyuYjvazN00hCs9TlixZKoG1PqhQ2BFMw3xiEEvfdhGSZGg6ABDeObY57R
1v+RgNxxQbpMHZByuXpdFqBYJ4C7qxJ+qEj8mTXXr4K3am7KAbU5MTrRbMbsdE2v7EgKCU8Sz24d
CA6LPjgHxBgBALB+9fELqsp6yi/iyJkQG+NJbszbLtM9DPKhglmBa9ILc8R6Ar9h1I2qGdw3ZoNz
PDC9P0qz3uXZevLggsXbXHi2XbpCcIV5EB1NpTcgNNcNLcHS+/OK+OtdirTx+QKP5YD93fkrjBvw
Dky/rQlgF/wZPlc0si/DWPZ+XYGiKBn0FfMRvi4BtfC8AUbrFGWJY07lhunijTjgpOpsV0tiGxov
ex469Z8M2M/ejZssZl+xYE55gq/7ZaD97yg6FyM+cOZfCQQbgmLANL6burNnJnbAE+++KISNLRiG
InRcTIWXff5vbfBYmgFhb98oHBCEZvWbOMNgNAi/8M+h3V/EzVpW1gCd1XjcSKe342Wls3yjqiER
o0ZQG1j+Exu1oeR9KIfhly+hToZWLar/oXQrRTbCJiTmMH45nz3AZeLdWKJS4MNrJa/Rjuac6Gem
yVVJU/W8l2MmHXC/1KgxHlnVDf3WRDVMmLGpqu9n9utVQTbOmOQ75/MJjpUbRSxQPsy+TNwD0Lg6
25ajOHwUZJ1M36HsMB8AXRzXkYK54cepJwXQatSMKnIau0CLrc65WgdGJEUcHgi1YCESYOvG6euV
w1TfXTzGl2rF5rC0M3kxZiH5mDQ7hBYKEF4WeQSqC7Ub54HL6QHQmkzY4bNvRHrAwjJSNQRcbU/Q
L6w6+i+y626g8EYYHJlbn7VLgWINIq9BbCAyunMOK1Yt6/MXL43q1BR3aJoB6DqPqbyWpaya0U3n
4Zukhi7sGcuuht9q39yyH/nbXmqYj+pWzXa5wuIGAyQbK1QerRem76KcbvMbL8E7GHf5KNZzbVSw
4avDRP+OnnYahuYyDe4JbwwFXDlJ/L5Ur21A04EudJpNJGrKM7OSpKNyFjY4BCTzPeTrgSexZosy
5vvhil2nchb2BMIR+zbAr/DR9ZHDcarhr2l+6YH9+xBqTj+WTVamawy+Ws+oQRzjUeBAw/n7mG2e
LxpqhLVveHmEOXLGw6EV37q354x+VKwTFvG+s633N8/pvQCe6aUFbY/LzpaSTnL5/ibxfEO9K/pr
sg/OGs6Q7YO072YTVjI0UodMEPvRWdZmNosSbNwDBvCQ9aXcQtcudzN3u0v97XsUWfU0h0pmGHDm
md7PW/uOWaUeIUvJrzeUi8rFtlzhxo498ePrH3kt9Rjri35RLUeRmykYs1sYdSh3yqVJHyD63wHg
An007nvir2yWEfY3X39DJpwuD7AQW2I+uo+zb0i0BtHMYXR6YHf0OGcZQ6hKjWCtLHWGe4Ts58Em
bjTfO1ecZ4P2ZWwwqyq455uZX/MoodZF2okd6psiPIZ7dRgeztNiW0RGRNAzhdyUbh9hrsJH35NP
7U/8+woPOPjX++0UTrSdHDFdZofMIyGQ0FcU5VUODgexj+4zgjLWXTSwRwe/Ey0drwms+oHXF8xh
Kvk9vNQRTmnx0a836wDzneBtnRELvX9T4Jv5N/Ul00mZGJf0TUEWcXZayg305qYjJAjiizjIka+J
l0bdf4CS4UDNW7mU0sEnGlxFHsYdxuGDq6FYGbM+hbgmywGJ1Zq5B2Oe0qFe3qSwjdYAQq+Ro81X
GXsYEdzEq0t+aBz6RS7qqVKx2fHeOGVrlzLQf4gEFZbFUpHMzjqUokGxrESVHaTB0T3/EIDSH7Ss
ASE+NwpimW/34Aculq+Q4pizxwJ38NeTtIZzxsh1gM8BWG+0Kl2Iut7oMrQKKZdibv+EDXCk5kw/
KrdAAPeA/RxbszRrneIym397m44R9/fRv31UBo+9qYrSGQoISzie4UuKNhkfdC2x61hAohwdyp37
8w0plQeyiVa3yyMKcBdynvH5iQKvOoJqx8OmGtEVr/FDwYajWid2HKSp5SsyE96tndMToGNvH/sn
UjcQSz3xXR++qJ6BSdh/X9ke4NWAI/WgU3RRolmFN3zXzaoGDK4mhz5SJfewtaqZ2JJLcmgQPYB3
KNlwzfATiA61rZ0lDoo3ePjmQ1vpqUgE1R4RgQvHrQbPePnLtbDsulYwJh/k/wEn6l33VxPxoQES
w1RAYlYuU/PBylEI7eE/MwjEXLbSvGBGoDxJ/fMwIDj5SdkJAfBXtBTypxQiqksGaf3TXeICE44Q
KvaGQwgvPQfgIf0o0Zk3EjPIPBqwVwnkDR+ykq+KI8OuGqqHfYEOTVfZkxKqJa+QAC2VDCffMHaH
/5hBWEpdMqTIGIbQjXgKw7QiUubyrMJ7zqdsytLCS5D72jlTMAtc4981DmcWtJzkLIJm/nss3Ysm
kSXZ7igAlqSdNEhj+BriXSF7512IjaWqx+qQH1uyGW+ncOR36lAIzBWDp8nyfyS3J1uT75ogFOUM
MmjbdpShhaPaAG/hmiv04NNq7bIoR0JdH9BTExGWRGPQ73zRNLLJfvOMZw6wJyOIeY60ySUFI3R7
9fQybCE36h5eSKMyBVuzNwqpheXASqb/BkcYTxqcUjTA+KoJ8owOPo5Yw0CfxeoswnTsouFekx8J
XWvhw8+giG376nDXxz/MkmpYevdf94Vu/Pc2JZwuf+V3qLBCfKDmCQ8CKwzR7umyJMz3vn1PjbuO
sZZSBpuxguhZMvAX1JtAjGmicWBN6oD39Ht4kGljbJlM4fujsWZRF4gP7bmuiCKwTqxYX1ciSqF9
kPwLR+aWvnHbWi3u06gEpIuw0Igjh8zT5UHVYlD6431Gz17LWrMgytiBPGHA9GsQfN3+5UjVGaAp
QGHaXwEQscDSMavRs7LyW42Fd8zSTGMY9ta47IdJktIfzVuH098OTuFPVD9/zLvCe1f2hc/9pjw8
Mk1wBWKsnrtabNHUbVR5NqGgvjWQSpTccvdkRRDEs67k1k3Kd0lsoArJUFK/NUuAdZdNEaMKsKoS
ASBkNLprGAT13rTeMg/rF3UcaJyyNELekvM8tgPxbci3b5g87b4KFV9uvzWVwrARiDkVBCzC+jOl
/5oeS7QKq8bRyg5dpMXWgCRXLY4KgHHvIcL5Fvb8677tzDZTeVmAGWICPHzsRFEWdmAmXYZs1js8
9ztRmKmAAZf8W1jt86PVD7BIbkKZmSJ1xyi+gO2xweBJrwcDMkwGWO8j1cYib/g16e0WiRnEs8hA
PL84OpQSJ6MKmZb3Ca4fJDXI3LLRc/ASL2EQv/2/RFeDotWRD9kR7slnp8fWnxDH3e/jl60SJMOy
39tkZUuBmsRgLeObCqu0r8WsREg5nJBwxXrPDZWDjHXSOWqP2LwDhZllRmGhZhy+C9zS/YyxUGbD
BCejhQK3FdIfl9DIMXpD46uq1h6+BvQLTfkXqvVf/qU3QlMjVMYGJ/bWUaa4gvov+8MJMwG1YOgX
cRcGqMDTv9JVSKMfEkHrY7vynmBBbl4nWE9atNJ39E8+ghKvchC3RXmV0BLUuzQBnAUP4LAoiOPY
pb7McIlcmgt6U94g3uYsW3oVarzofEwtLKmP9On0ZtcGf9cUBsnwIFp3hYAtZn6lajtC5tGwUcik
OEvrxYCNOUlVp8C7iG5RA/uYHUcHhiFTw/Wd/tOKVTWMCDNjm8vhTt3tGWpuf6PVPriHn3qKiPM8
85MWoooV8krLau6A7uvHQggNCnlzDrG+UomL7KnvU5eAAZ9eF9vI7hKFKGFsXyS7StJuK/bBvVqP
6ipr7orSdXZaqg/NFqU20gOvBkEc91eIm9ZivkIKDJ/FfZGo8Ek31H6q16Ac2F+gfqcJxUMBIVZb
xZLKeQy1KHQr72nXqJL/toMmNg4SsoW9Ce9dKUgAYaFUPqfiVsIaFSwe4MLBKXQ+PYSmQ+RRTTVE
NEa9I2Y+e53B61Mi652pHfjD2vX5QnXRBGnUrgePGdrU1AqJ3rxwCUDK7zadzAffgmkK246+m8Vp
XI7OwIEh4mlP068iRkBflHPO20gP/Gnjg+IZwMylnZgwCx8B2AlzKC2CdnZ3x6hCMlJr19Z3HSoA
Gk0MUR3FYwWQJnuef3OA7hq9xch3+Pv1X2N5w9lwCnXoPbezRFHSzJv+lM2rq+QoF9cmbZJnHc7P
qiBej2cWKH+oZBFZJMWQzo9yNmLyc+TsTk7o2F30MBLVFpPoJaGKFxXVzs+v4OWidijH3/9pG/SS
vMI24BejjtwO4Ci56gQrnTchRLm9lXSyX3j2MdTpJS5suvGPU3R+i3Sm9rbnMQb7Z3G3gNKSwH7c
To91P83KVT1qBcKt+dsB0Qy9yG8/E/G6yzzTyDo6/f8v2ei/47Gak3QxPXGb8iEjVhsoy8WZ0oL4
ahO80JKjPI523Oj2fboyd1mOxiFyqebwBLQu+5+rc/jtcBguJK4W+U/0vBeqk0Orc8yivWIHJ4V1
iJqmAaltLdxOj9Sk1sEA7XLKEsSX2NRd0Sa5oUHbQyKou6VQbN5+wh5tS18GOsiDcJmp8P4QpSP0
C6maZlCrgROj6WbyU6XJzaS+aMvRAfZFPCltUeGGcy2egNZaJawNgG6rtPYiuQc7Avvf9g2qS/MY
XvJY+XAKNaSOD+1Lzb8A0d5dq3Ua1pVW8RhczkEevE6FQ4FmF6IEtKxG9Sc7/gnJAW8CH57tE5GF
EmAbLiRpcySuKZDHgXbjXwBDyQjm8S8g3zSLu3FzJKTPO70hEqGjxc2KXdWGftngxJMuZDFPjJEY
QMXGiBSJSM2wTcfb4piLl6i82n4PFMF89+L8JAXE+tuO32zxvCChPxGsInJoq8yBGSt0Gd81w+ZQ
2jks62oOqwVy/v2npExktKcft7yaP3sF1RMKX8NlF8LNTyb5f8CAIUEV5Vyh/wlKlU2rTaywx7eh
iluA6ghRD+V07JEPA4d205vHa5N1MR9mVYZhfqooAlciLo+vkFMruTJxV2jAqbSJhU/eueUvUFaw
RNcwbS6VZMNAO0F7CI3OmxN52l3kBnBVWDfCTLeYQoLQqQqtN0Kosv6/Y1sd0xijHcmVUDCUNfiE
p4/GMpfmIJ2pyLbY4/j4FnIUyLsyU0S+3zlq0ROpu4s5j7VJIPt9PzN/ftHykm5+0F5xGlF1z4/2
5ZvD2942yzYLIIA09avjRuyGmnLBU7d27bjaSMeiz7hnoIGODJBR4b4smKRMNnQEncjnr/DRuloL
JUr2/Lv9vfb3WEHWqY5/VDPvMocx/5GUVh3iQS1ijAIA+AIME2qP6xkmbTYew5wxy15zmoS35tvL
SjatGcQ2rvI3SuIgs97NSjvCspNLJVwioYcdmTpf3glCStH6OJprRqs+Lwuhok1872MYS8smbRvx
AVZoKkxoYFdGHgeH+FnltB7bE3jWPEiwzbO2B6PDQRw3rtDpYlNcE4sVkB6nmvS/EafmNhPvGz2t
W54nJHsneirNhpoywWjB0f6pSNhVlxuQoxIb4+mo/fuhFxILvznaQbKT1o55cbnFQOv9WxWxcVxI
WfCHYkJEJswgFAukhiLuaW7IRjSaocpbD6z+2gLxZNWfEtspXREnfCM52oFqeuhUitwVxxagD/91
uuPJmcDB0VlrDiUWu2NcIy51X/Tl98u4W+JHlaCLjLrSdWTH4mhCBuJEqG63t0L/sMQjuWugdh7+
RL8/h2oMpJ6Di22cSecPVZ2EGsHN7kqNRd+xnbF1WMNqOJBEZX7o0iA/jVIJS296wO8ZNGdqJgVs
ap9WpA2hjNsDRBL4rYNvTU316fj6QsMXd7pVVqWRcKtLGUbiMKLxKvkECOFxmlxc2qZEFDiw2S6p
Jk3aJZn1nrw37cfbFlWT3SIwoLY+eTTCXdmcfBGH3y0TaFqPVc9ZVyrJStIsgGvaYUHJvLb6MW6v
C7C+R6jBXs/9HZmW8rOHWrHdnzBy2Rchg1vAVoHqMp+vVYHnmXjOQPr7YGtzU4MZ7tgwpFptyF+E
ddkiW241ebsxL4fQiOac2Wyb5rsO2S8oJm+tHbp2j+UBPwxrbulYcLlaS6imoMbUDYYjBAYq70ha
YAzqhYkbB23Ly31iTcqfKQqROVjUlTc0oHC/ZTAO6sWZ9q6QR/h+g3TbygNZSX9ftPqOybVbI6ze
bMXXqAQFWT4kjI0YeUpBdSZnmajtJ5psjAXteDzWpq3nzBfBjg28Wd+cCSouVEqgSD8ZISvx1LtE
W6a/kOTj3Zoq0EaC47m3zlZmmvd46khVcBrNRkxAwHYKIgNytviBqkjGZVxmVc7s5PSLca5sgwY9
FMjlSYa6TGAjgJOaE6fO9N1rqyjbT//DcHkMBK6Px9wSmSk6KDeVVirVjGnIeJzseqd+f5J+ZgXY
scjq7aA9dHerwF7hXiVkWXd6eo6EAX+qgxUH5lfGmUsM4hDwhXd+M/OwK3iB04LebHf1n28J89CJ
V6vXgdB1BJpLk6U5UkGT+o0RxGCnhotp9cfRto7f3FLcAGYiwxVT0VYPyqMhQs5dVN76bSar7NXg
UD+00O96VfLIaAZfMF3YM5XGOgtFSiJCiMdrlRhXcWa3HaUdeLvqGvwiswfQ4D/qHE88liAFem8t
TROf7DPDwu2xBlDtq24n1bY7eakLFjUmHfa5DmbXoKIvzQ5/bjiNHh3gfB670fucDitTobAp4Jqs
6WFVT+1NbvKzOu6B5+l5p/ukor8i9yanRlfVGk7YXDy2RBRe8N5pi7IafYn8UuwyNiwm4BS77ln5
lbsltuihGdU3IkwZYbBG0MsfibKqbtf/lBxbrQRzQ83n7X1yX3bxP6sFB11d0mKp6Z2KFtFkKXwj
vVg4Wm6FVfgY+9Oo3MaKZB6hnSzOFFhhmLpLZaTO6Kk1KR5tU+ojUnydRRLH7SgpvZp/Z4GQ6ZDc
tBoBhVdvFOXVvfZ+tjFcp2UKyYrzXCNeyg66oRkAN5o2OBd5cGr7CchyP65HZPwWOf4SAAmUGZ0h
A091/twsfxqvtEZH6tp9uLWM3Y5FqoCj+YUD3sBR6rB9gqbhUrYbh1K/A/YrJTn8saRL/TaOWbM5
GmgEYLVRHWemHO7BOLIkLXOpRSNZdMXRXB3GiBdWBEN4fZSzrbPQAFcWghsS8/2vsZSljVDkKJBo
12JemSc74GSSBtQHdWOaWLjxvE/aZZ8g8t6J9EA8GZjXZihaQrl7dW4v80QLMgL9PZcrqEwKkKDm
eqid2aV8qcQZaq3me9zOBB08WddrREEcxAIJf1UYqh7Pu4rPghtOelZ/ZdPdlj+1vleTKKNha7SY
g17PKBYJv+p0tcp/UBFOFjXsLP5LLI914pEdy6IvXBIfdTxzbzE5ZiUcNpzg4UnaBmf/Cy+h93++
D1hyvlqpf8q6BxSgc7Jhcv7Nn5DiYStJSeyNkww/tRHcj9S90u+elzHkGlB+NzB5AXA0aaJ9zJI1
8LVeDg3l047lPwfveaEt+JucPpLC4q4x9dHfJ6AR2IanFOR2pZ0uihfVuRbG5kAouuA+H52S3z+z
lgX5REnevLCr6odhMXIOOCuDrRBeKldp436m0S4ms7oSDjA9tUn9totk5G1pEO8ckCl9rFOBqxPx
3XxZvShlE/u1/26UTDe9I5Qt7iT7BJWzC9Yq/LQXh8ArEi93qMZXNMVTfyT+O44Ay+4Yzsx/05h6
H7J7x9AG8wYlsTMtF1E04n/P1pFADIlWS+Zq27JT7DukG3sZaxNxgqJJxtXXr5jgrl8AkwqE8cOo
Ux7/qQf8TBzZAUuEpOScCOVpdBS0rp/5dmDTciMiYyRDeDl+Gz8SauzQvDtLSMuydeYFwxww3tis
ltAPduLgUj7meXIigOwJKaUggo6BiPQTeVq/taKWKT+GZYROv+vENfx/UcsE5PzpYoHgJA/OEYER
vlPVOjony/XanMz8zUufY2aDKGO0I0Axa5lH5f3o4olgQP03/lK7DhMskfaZF8rrvkHbVDmJ1PcU
4UukZ3bJhU+k1YZgpNLZnspV4slG+aVCs9ndWghYF1vqX8GFjSX3vIPT5CXLu+tVWoznUlyX0hAa
/gqiiGuSWcm4ULzjp4z0X9PJRHR5KSZMPZmwkmK1b3uCyFhtwVrMbnC46TzCiHNDJKp5vSQgRNt1
n1QKDYki6tUaWHgW2JobDIJXGcn/RklH7nWsIpPFg//HOz5O7O7wk9+FwHJRCMR21FKkS/0P3G5j
H0sR5dQx90QNapoC115WnWL2Kxg1T0SVKlT4hEECzr0t3JmXpYF4TT/E1BGCPsJg+mJW6/cJ3eq/
bOmT7zk1tGHTEIaKYm+taMqZI5OskTm2hcZIj3aOZTtmjSor1h7D22AdK5C2dtg0CfArp+2kZtFM
nN14siiFTWY1ObjHCaPaLieG0iOVMOddlY836TMYQhUM3mFEI2PRaaCVvwDklwaG+SVSnGj7OWOS
U6nD1yqTp/YF50yRJXLruDbYefyTyDjdzfYaDV19lH3wn08pa5V7GYQqKJOPVIukreKzwCmsLvto
FJU4W0ydJTR1TUyyYpO9QWSlz2svFsShTCBvnmosh7xxYYSXlygdA036QyG5etIJszFvpnhlXL2I
S0fmSn+K9C2D6uY9tHkbKRW3KBcsUUuSgdfK+kd+AyLxOOVzhpRqYgKyTbLpPL8nZ47GwyFaEvyx
6ypcXdNnzO7iMVJ6ryP4VefGfABG+WPkun0msix2adbk1IdjVeu3bLEeQMrqQvNFQae8ZH1TMh1q
CguQLAHlKh8UrOlEWmX6Y4nv/WK+T3ZdFou3FV/2AYUOd/tbsBzlAQ87q+kYB2EsQzhsx+gMs7AI
uajjb9hRA+YYi+I+euigR1xCRfvhj9a+ASm7oLh+q4/NReCBWUGoTXEGl2DBWPlv7Csp6xbblETH
n//ycLNib4JrPGMWvDtHU5V6kzNrxR4+tYd81Dj/htsqqpnTKj24vGAxcNdfm64NjpklrEnbn7+e
U4cOFqy0wKrYgteJ6GSEvvtpc2FHh7cdy8pQweWyBmyHok8ltnt4/XEHS8Flp7olcpge/107ziAW
KyrdSubLII49vfdvWW+yDNHpRMxxBnTlqK/p/yT36K2squzPobjQ/hwaCcsfAgR3QfSspH6aDwfo
2vAe71/PjSszM9zuwI39ZNWB0k8qPy1WPIg3gRfVYAB4r1BRttNgMNDBcqct5sIr/Z41QP4cvAM+
f6eSm2mz7oXRNLqCWf6K/XAS4Biru9eNIsCB285RRF1Vyxr1W39cY+IxNAEJgSXswJ6H9x/KL8Ga
0l+MmSCxWCx9n7d+kym2qB5kzQXJFIObCIYjXUprBmAnWcijZweTToftkc8y1Kyl/9PiK9E9HRIp
pR1JqVOhf93I/nej0n4vVqsyuUQu45kaqewlo25ZQaHUKNW8KZYmtuKqKMcAmGmhPxqYUysLBVb+
5pWBml5SHBTemdli9GomKq78udsEQPeRujRzgI2A71TuTQLEfPmRHm+LOCgwwBUSQHfPny/4EuCn
HhiQgwmfJ0xAm1ff7X9aLtQz848LpzpI90J8nk8hF0GoYQ09k2z77JUj+n7vtvIKqZkc9nPv0mY8
8y5zP2Je+Mukc257qShshQsbJZ5NVPrqyzqTHT6/max5YOX/RbiMk8C42UvyhIzybZc1+wIBoND8
eXAKkKF3bHJJmlxG8T3GTmCwJHZoqqkx6FwrQ7kdJ4U74W2LeAQTT9QGlqTDt4jRoYsaIYRtDNSH
KfQHV6SKcMWgl4g0UPhKuATyyE454TFQR2TLmk1Mc9j1US0qenMC4vdQm+gGobTtzYzkqEjI+ULY
CFqwXiBxHHiQ/YcFItbGnnj6aFV56yv6/JNbuvJiJ9DXYyKPWZEZmgTOlgPZUQPvoK7Tw+2rpQme
+nM0vStnEbGVMviuYDQwqHPUFHxDvQpT7xuZw5GzYFHaH/ytHw6N2oKnPhuo0SLpAiVafpKJuHKy
vWZ0MHwKVudNCX4gXMcVe+7BxEQmhQXLQ//wz0Nc07SpHbIQAL7wweGyXIbP2+1A/GQJhh/sRLtk
jbb5Ti5+vaFen0UIy2J7cBSKSyikJSaQ4T4DBJT5762pKG0iypflDIno6VToRGwDiZ1G93I4dpdo
ys4QX7OSB7QeERCIr6WFlp363ZgI86QOVFr/JrK4MLCWJnv6trdLEIaKJGc1vleRx9VnteGAWu48
x3eSYex9xwZgePAUcDvNaddDmSnp9i0o0BAngiLbGFO3/bM2+Lg1DivxLNBIIL0T4awVu3Ng9lVP
Gl/QwrdkbV0q+CY0mjqPfV+NWfsiXVU/arOqNN7OIJyp39s3MxT8Fy+hoYJ1hBACKG/yg094D3+k
p26mV8nyASceBqHZxh93eww6SyyJHRchPuvUmecPe//gFdJ0m4cB/cDWi+o5Q3c+q0O5BHy/xfjQ
ki6pVn3CeW7RGJE+o4D7HjrY7RCNa2LQKWdVB/MfhUkmzeLUn3tha6RWle+qi+4viQAtDE2vR8jt
q4B3ZEgVYV2x2btb1cMxnL5Jpqd7ixitP5g8KcvmNP8UIdKxsbCqrZ3B59N7RVjM45UOd/KuO0/t
vgtK/HvqOm2m88ljHBq6EcP/iBWy4slnw16YmlSx7uh+RbC6c1GnIXm+B7+y/PMCnmPcwEZ6TOH4
AVkk2powcTWp9c0ZIiwlXD/cdYw99H4S9T/DEYsQM90POp6VuGtx43JFGS1ZHx6392H1Q8Jf4ZI8
phW+SznNrjEY8s7m9C5NxYj4pJJBIkeoLciIxw34MKjkpZWJMljj+YY5uq8pOVXnB4m3RLycGWzL
/Xchj601FsR/ZkLsG0I4w755nCEJq7IJD9cV31GZ3wcbifeZZiakrsmf7T29xcYipycP8Y8BDKIM
tnPSCfy09Lt/wRPmoNrojZ960hEGRkbtXTbVRresZ90BGjgvgTG7FXMX7UDNJEKXTVhfo9hRc82x
GWFGEcp+Y5X5ZY2XSmaXSPw5xup14YtoeX/COE+kZN8aOqbZX7hSNeWSutNNSvUDQ5BB+6OCSu0U
TVMyPMSJuPJTJ1tNcqWdNgbckb34tkYFi+tfhD2yv0UDHanMFe+xEMYP+M07V+1eh22gm1RjZVWz
8D4IWb/PdPcJ6o6qsVj4voUKgGlwWQsx2LI0C99DkMYeqOJ7dUCtzkNQNCuM9sG/uQHI/9swc8UD
cNtZi5+FyuhRB8jLqrvnoG7yKsjrx6UIe4uV/noJnEibNhrUOUUbCw/ZIwD6iyxN37HM7gSc7fz+
7+UWLl9nPdAqJn0QF5/iqcrj+3jDbBAQc2vmFqHyRiA32DKxTH7kKFSHg3Kku7Ays7SvYGk2BE1K
gMHTuOxRuV4RS5uxSRAAsc7M2YA/mcLuu42rRzviNA1hVSA5WsGQLIYyiVjJSqrGqU4uR5J74Aik
BGgXMzlDtoBv7ErdJe9kN7mrPljxfKo6s2zltLoGijL01ttI17eCvBrVI90JQQUDvivXw+zCgRdP
QpUBCiHFPQqp+I6kBZ054unyrT1ggAa603kd5AgMXNz4Y1ZDrJ2e5JqNNZ8qz70qKBm8OxiR7iSU
FLXdY8gcRmK7JKFgvM/IwO02cH0DsO2qCqhuzWXfaDUXC/0U4zVBX16JbaODkLz9TO5VkF4qRx0f
eYg6t3dUbVz54t3/JYC9KWeGUvaXLnZOph6tAOiDTKdRDFO3r02pFGb1tJ3y+IYPwoV3GNFqBUeD
92JwvybAAIYdcrfjOOelohvJ9Sgsmx4L0CyzX65ikBCs7/J7qkI+FeJtWIpND3vHSRBQtVAVLNhs
Wjbbsstr97h9yYdz41wQGIk6lkVRn4t3LTzb4hHI40t8jcsafaLQhHQs0/1DIkj1PcpuxR15KhVg
u1fFXe1XbTzE6uK3vt1+064Zx7YJlyQXF6nFJB1sK4L1y06TT+sgspqLpRt8lXg/8Pg2kV7zAhGP
DOkTCsDhTgawfYlayoi/BQrvZQMiiSp7IxcPjkJmXmbQ724aH8G4lQ3Bp5nmuf5MHEOen5Uc6fh9
ivXY31kVqJbRHyfqFxrEdvUd2I7d114Q60Y99DRUY5o+gRDc9/9dn/pqL9FKG5k8AkTvsC3LJPq5
OifI8qdi+iQKZR1/sagYsV1Tke2eSEztot9mt7Zk7ahA341jvHJOrNoEJ5InEFPlJjNTZdIJqmBt
bPr25FnlViZNHEL5mrG59dmiY8abvtz86dHWsILRKrNtdm4+F4nfz2RhDCaPgfSi/uCwPWEbJG0N
P7o3raHg6fwTu4qOb8ecqFlPDPn/hxOqhAdQo38YJ/Z/MIYAo6bgZdI3AZFMEbBsQq71DyvR7I1T
+qxhDnSuP4/OZn8+SsNAPlVpZFt9Rf1rtTyMe0OiqJX7L0MxNK/1k6r4u5nD2A6u1jWvmtzhSNuQ
bPUDAqorqN+f7XlVcSvinxVilrVxLMSNb5ug/3zvP63D7mwgM0D8gz78ix83S/yw0RGtYMqFIPyu
QfhXNnz72FzHUjI/5C+ceZHvfBqeufcijGI4c1Ga9eqDEKQHMA/CKN6kkI4LpVI6WY0g478gAKhY
4Liknar14QYwOhYqZWiq2yJ8HyelHPzZ97Xjug0AcSNP/siR0uweBThRl5uHsPJE1CaIsxlmiohy
lRtik3DoIie+PmZu+sks7mg9Kyl4IyIYkx3T0YuBOXp3xgIw1GXGuBXZO3O5xpcyg2zXJDsw8Zln
bbOW97yai7W9sldUBHWYzisKqRyZSchz97f3zBlnHsx/4odc+F2LH9PP3gmnAd2ZezavMkPA+z97
yMKi9ujRzHHFixbO/OD0HJunv+g3+KMnGMCBo43SVOveca7WhJzBFUayPph4nU2i4uRgnzLdhkbs
sAB9NcNxxzwAQYN45pOy5qgnX8gYXpPXcHDQeEYnVEOZsm7/ufMuY8X51JJMtObw+91uONXJhZKu
agG4UxnCeLsp7pukut7Q8S8TPehX1qHahbISmQLMDpvHP8Y+amftewjfdNjctOUGIxyVe3R2NjOU
5XSPTiPcQEi9nKvBWl12b2IkNPmROXCIChwZhgOfWJYBfggoKDJudrNdt6APXfOLeNCepFO11BP+
NaW3HGxSkwWRKCcRsPEkWBJurZBFYMOkrlpYdKCaKPWm4UbJcskqALLlaYaPVRPd3tCcQGy4Tx24
scbKY/kDsL5pIvzxiqw4B085YzuIlwPhN8JspZLOc8UQ1zuT0Cq9NWbn1lYViWeAZTfgbGH+kjPq
rzo7syJxL0YBITNB86wXCgsCxsqCe0q+kTBV8XkZCp79dJAi3Qf32JntnGUiuPMd3VFN2zuf7c1G
0Ggcf2SFhfklI7+RqXhI29k5909Yn4I8uqmfL/Xk6HlUw2Qa9ARE2Y6g48w/7F2AJTSKXbf629wz
BWQwQcUTcr6FsQn5WB8Go0TC6KOCqR9mWx7WkAvMg2U3RBceBhk/VHP/I8MZHKWCQ00YO2GXx2YY
mHEju6Ail2dZp8v7frDQ8sRYqjs3/qMObGwIQ5QCSC6Ht3ZYFiuZecHSXKVHNHolv1wo120hf2rL
Wuv60zqEIqcZK+eLPhB6L1GWB8b4Rj/xwxAt8YjrrX25PDJYQi3xdoBK3LDJYnHo52QHfxtm6osf
6T0H3h6MlF4pSqpuc4khPlPJVkbXAMHwzvEZnoQV8f6f0l2/B6BR17c8NwDJYE0V6EpqcG9SXod7
PQkWdkYzeAJqZmfiyhyfyWR/1afujurp9ph+1ghn+mVNGbCMvi8y3kdq0osp/HzDiU3MH5NwVHpq
MlXeizVINXdO6thkRilU7RCIkrHIWYJ/LhP0iJTWfcgDkX83iVGleDoVSBJCg+jOVyrMc5BN6cx0
CxlKPPQlheNlR1s6Qw9K3odm0P4hZa9x3jL/DJ/Ddyp5l8pOJf5J/QWJNt4J+NtstYY+dX+1Nr19
6M9tWKV85l8ktqymMrnKtW9iFcvPj77RVYj0rFdSswZlFiFve0sWhQ+0DQp1M2siLoZGCzt148d1
3RYYr5VRkKnh/upOr3Hno73b62PkvKNN4adOVzLyajRwnsgk5AfbVQdzQQQz9oQOglmW2FiBIrkt
x3xwc1BiGxgRVqlTeGJ1v+YjQbWs4aWAeSJ5cbnkDTjeS/Yv73MBxoAjKxMFzIVjLmNrVjUiPBad
PeFZG+9idRfsUYVWDa8vn4+pWIqTK7Lfop3q4JRDQT+l8JeTnApoynx7wTcarX6u+4Jhrchp0kbT
9FS9gj9epfX2kgXrSH5h6AnrI0LoJgmGv6/EjRDnMIGYNN7kBsbZcSyS+N/dq6pe2a9L2lXlMips
T0L68d0DhoNXxAfdnBJPIAJfz8WOYJRU6/B0D/9SSegsiFlKNKYwhvDJDGaIWOA+wt6z6ejZX/Ju
CFTjpl3pFVpNfIKd/X8vvWyGhhYY7Cq5612/ZH8VBqsggRzV4WYnGxeeq+1HsmscR49Hx+MN58iD
7lFsNOH81MJkALutVEJX+lJAXzxi3Qujc9HCK0muul/Hw71ln8BmNFma63xCBaEL9vVqYDEIoS0E
WokOjItmruA6ICTCbwLyvflvNVWzbeM6oklrYBJ8E1LJFMmKTS5bVG11ZyvoVHjjYPRVzzvt9K+l
+GK6bb6A+N/b/e/nQLLJODh5tjrxlawaYDniyXvHEJ+PiihkYZAjt/4dRHK7xRAh4P4T7YfJGMQa
KX022Mj00POSbrXlARXoj4CvOVhhME6XR08nBErMJ2GXDCoXBWbDhmvoEruL+oumUt8tAXzeDZqN
j/zLUvRy6Inb45k34yb87CZjrTq2zA3Me85bI7QmUIKnRu3jHyS7kXZLzkma3bvGBgkGRyKKsfbB
PMTgXXNMpycnAnbR2X4tkXASEPinb4FcjAT1eSe4IZtW39rciLW6kKhTYVPJvC27UmIlhA31QxON
bdCuWKtfFZXcChoislbpxGog06ETEoQimttcgk3naNDBj+1I7yxwVfgDLarTTxV6k4N95SwdzKQs
zwtvyuEvzghv/2G8wJJ0zm4OCE1edJPw7HCU9L6lNg9Th66ZU72NN5pSTqQMAk0ko73eLw9UD4FE
V2tOp5EH+Rfy/80NS4aYl8Jr9rUn0BI2l2+B5i1TBbvjLE0UIcHXZaA9IgLnEuzPip/azi0PF5mt
5XXE9bup4ur7nQlkUcwJNVhlwFQEu+wylvLxsILgu89BNvEI7DvFM4x4ywl0xPSNtqz7YuPHTsOI
hJLtjBne3aDREpcTKvjdoMAyunsslL1kv3fNMdFQ/PMAFMq7DOARQyxEmI3s+sObB5Ig+nyb8M9V
Oy8CDJd3X/SYj4VuLtRRRTj8ImQ+xMw24xGnnDZRCnICVcfYe/Fgs8rGLGpBkQ08X/dAfubnXwZg
DaBOnitQKVOwM2CdyqYdM/0GqhLR1U9UJH8QuUP+uuyJ1RO6LY+ZKdGBKt6qSilC1aX6aRbTWQm9
74iFhtbYnAFvQ9sEOjEWh3LjNdZEXj00jXUx9vjo69HOvI6HWaxGTHF+FS5TezVftHOCA1iynE/f
4NCbv/CCwPLnvZL1eSZTDLmm6NE+0pB5BzX1ZPtwlkL77uGsIts4xD/FAhrInyLQ5nNZTnXO7Es+
zKdPJlX98cQ7qVPnETxCrdr+F4UITnlc6FDI4nqT8807+98pRBJslEebNTx50NR645xiFtJPGZ0Z
Z9ATk9uRia1Y80AxCLdJpMZKiayQOc39mqJrKXB3HV124pnBOZCaptY1ZFCMnZoKBNIDZLXIwsfq
n1XDzAZRbX/qOPrs98fkQXzKulesFgOxAHIU533biY9drMWAFeYTnLM9uc7pGGhUAjDRI9AXdPX6
jvgPdeXmBdcPeMYvevsOyZm5zRGbGtCem1n+LoMtuur6+FWjxT0Sa28/nUAWT2CskY6X8/cvTtbw
wAxiMMJfE0IhXNnngoIjvnmFmBzmNkRMSrI0zVMBFuSO3JARyybrHAXL9nbi41wxZDk+5Ri/v0jO
nnn+FYwEf1q3PuHRO7n3Ig+1qIZcF0M4rws96GMCU5y3qJeaQB5GNYtvYeN1sIzqdu1LZWutau9z
WaLk/oMBOZHDmCa77G6zN+3kTVuWLII9FKUJF1MWkcqkQB+iurKNZ8f22jc7sYZA8ZgdqFX4IBbo
JRpPER8GPxQxXI2LWuBGU8EU+8IhVtmxOqc7UXdY3kaMfn1+mWdyyrQ2o3wupnc8CM8H0jNepaHp
zNVMvJj6RtmkX2Nzv9V+dAnUkPjuTY5mDqHFconZ9//B//9MgVyJTE3IfGrnHNwUHCbnwaAsIYwK
fUsqgcAt+n4VY0mzyiGnTB7JR+JYeGIAxyb+qtPWdDAVPMVGq/teyUTyxLe1Uy6L8H8uxV88mMLW
95kxQ9x0vz6SDEbiry+ZUxeho5FzO/ySd+IyzggLDAOUeHtULYr1Tcs8Y3ElBlFgsss8K7+oZxFf
P1gvgjLBbch+cx1iJXnAqRbFC81+WjhvZeno0i77oDgL657YoL4aMvjCgY2Ny/NpWRMAilOKAXiB
J6Kt4J2ukDZ5UgRSf/tjwZZPvvEHXRG8FXrSudkqWE7lWbVKl4HR96bqN/87SeVQFFexYSOZzbj5
bcpYrp7cYtr4pK5UMxE425f3+aEYG/c2I8Q8WIgM5f3EQRkxbBMVNuchfw0/HX/p4688cx9yS1sY
9Ifj9hB33RcKLu3dNbKa+M+gkrq+QvNvYzKrf4F/Q2G8DAjPfa+fJCcUWbE0mdM6Uj0WtL0cqVTa
WoI34I4BeNOMam7P9LdlWO8eskJdlnN4csO+580Xayjw1m8qZZjo1szjpDAeell+sriu8Vl8EcVR
Gg7Gv44A9shr6/lKsbFm2CkwegSfS7p/vcMVu+ZEKzWXODadqmHxWqllj+lLH2tPaCI1X064QowX
cGYc7+74h8Kggr3aMzm9W/wBrmBJV2nrmBGEOoHKmr5PToRZHc8tq8oMfVtaQNevbRk6/cBx9Ftj
ZqSVCeN6cvMXguvaO5fZakOc9scslnFt6cakRGo/upguRR/4AOV0n1G9vJzuRmo8TSQyCS2Z2qEJ
4pvhyhtdCWQE38HBspEps5IiBBYZFV+4D3YjnjZ1cChZBGzu8ahcq3UV6IN73TcG44HK2LWs+Ktf
ix8qytb8+QxAKhZdWirotj2GhmgPQ1JZVLPINleZItyjdF/a1F1js30ww7+l+VDYYYNu8aJ/0DeK
/V6yKhGDwdPjz32rnCKbL1TqUe5ObOR9MMn9x3m7WPKFI/gMJJRtYw5QGuM73XI6jWxO50omQKoz
ITc9hQWUSzFw2svuBgesZiZEX5WRn2gumpj7wJGMw+8fkrNgWj0qtWNM5cHDMqhL8dC4EfwuhsY0
jXHjRFkCMBr3ViDHVU4lorI3x/Q/x/80/jCaVk0KXRnOxlIeqvdqZSRhCUFJzW8gZYC4tukN0T2n
7DjClNhxl3lP9eP/4OTo3mED//mcpg8R+uCKySo/vYfzZL9Utl5s31qS7FxUFDY1MzDznkYEZDoQ
HKu/RmGs0xNO+kemCazcxQo0sh8iV8avBugnUH62AbS4ZPnv+BxztwUYz18QXQLTmhOpTDuz84qp
7vZFNqvoe3j0JjSAXeuWDrxu1xJFhvUSmfi4q/GK92rqdutg8SNaygXe3zpOoiXY7W/9Uz3KrHpm
1Xl20a7XlAMdQjijX8j6dmqKf0r44smzL1C531maZ0f4zO+Il2NHvFI/6iJMOHPLcOV4KFDtvBb4
Uu8j34NCn4qVfnFHwNPaIOER0mU4YdUmYVqw37x9GS0woGkWrKLRHzW3Od7zl+k5dyibZG70kdYp
enm4oPZvZwQ2Uamy37leCHb5dMJpznraSngBhLZNDxAqrO+epVdsTzsGm55UV0WtkD1dgwxUSfE9
8InQL8QPhqxfZLS9/xPz4+1ywL98tDYl2hBdNAwfL+oglHi96gy3ByWeXkwyXNXfQl8CVmzELRJq
fpYqn+dZ3uBdODPtxBb8uy6TEHjoCvmtAz8Aqyir+loJYi/IXi5iyfz7BBAAA0SOE2jquAAdCpRv
UslnKd0V6zBiWhpiZTwAbitF3NLHuTOosAAC75dfNmTQpvQN1pgDF+1PRlb9TWBupQ4jHNk3ffrS
DMMMBCWbojhJugm1murkWVO6jcL89tz7BFuiocZI3jbwc/4om7rPa6/t4Eonzc2UJ0L08lWXuimr
/EhQDW4HM6e9n4NmbTxxzyJQz6Di8lmlSc8zE2J88QZyWdxgJoky1rZffN/gGqKxZ0djlVbEmjQS
dmfF43OrppI9+mYAsHK4lnI+Wh9qc5EORjgpp8Wh2c5OxgYfiR4MZBQYUcB8h8kXnoI1L4LxvD6w
+42bUEipja0+KJHrUMJExZNTFZKmBozNUYByeF+6A7Ys1rQ6Sf6v5FPKllwVzi8kbJzA+6wXX3EY
BxFcSE/AfRDE+Nhxy1eMcpZ8wh6rkYnSkRnfBDvhro+TUdUC+HKbBh3C2HUTpr3EbVNoJvpFHBMs
cNCdFrl8FfQezg1lZCBVyQ/6iAmbimzgBaIro+gpO6v2Mi07L28ss+xFDbnPvwX4pZbJtMuIfPVa
joXhaRofrjCfwx20m2wXb2T4wzEoQu1poqQqcvXaI0wWoFcK2PSH6LesugC0zgJZ+EWBCseDiUzK
KizKWL8+xDiFaAtyQnCQuBrdIv2eeTF2KaY6cj63Dt+Ugayef/Nui5QPEgB/lIiXBdfb3XG5HrCv
S5xOzIs4RY0zS9h5LDTNMQv6OFeDHTnvxDUhxVS2w74Gq6d6fqp7xnZoDz17xfRPBd1CbC9TiTHz
IlhqorePUJ3XCBxPDJ0zt0vjHwpjYiy7MOCT/phdYwS2FnNxwG43JTpKdw8kAmt+0WQCXmwN3Iy5
0bdyPFFZYvcBanLBVlFEYbdieLQUJYdzOXsrAtb7xgiZ74yuRWHrskrxqEQ8QEBYXB2N7TO9LG4d
FGteBaWk0wahyIJO+ghXYP32UZLt0I2IcV5yID5pi9o+x8stm5RsfBPysZl/8Qe3uzIyBUgb0vAj
87YTTzOA0DkwLcqI+Dn6xxH9QpP6QJ7j7sa4+yhDMaRLARVYeUptRFWrzmh3BUu395wdBLqiYxx3
AKntTTdSCcEe+JZfAzmB65XAx478WXL8B2K69p6HlF767r2Qn7Kp+qGuo6GvINbEiDRI75IPwK54
YkE4El4telMAFovw97L1sL9w9YtrzwByeccJtqX+2529Jz1EaICo47O/w6tA6ObPgASGxyo7ivte
0LEzGNKiPXv8PYRIAd2t+xAyOjbdI83CgbnLq1cUUYxgFGf/7WkrsqF49mBuFWMSJ1JhRW0NTGHw
P8gLYzv6FLEamQyX0TBd+5dR5Yfn/GBQtYZU+YOdCJ6+F6FMKFfHfm/UOXcNgyGNXpoDkKfb8svL
XrZWDxrXY7UczjvzAQ/fu06SfYonMHeWYm9qkI0kBmkMTJMMCPlJH8HcJL6v+8dg6MFNtS4tfnf/
kzy48PIvppGyZPxtkq2QlTNrOmtCUQwZT2lgQ+lIW7FI1CbNK8DH2VYtNsNrDxDMPp17YnIYc/hB
vPt8GKwWLffa2d1DPxzaYpsNrhCylLXHyyU3JBLok5iMyzY8oVfl4QV1PW6PSMjSu9l8znI+1DS7
7f9SDr4Q7GnWtqwCaaD70PNf0IKzeRh8CEuDkHwdj/MZEMuNFn8go7BLBfKy/6COzhpJNFncHBN5
psRdf33ayRD/Oad6Xuh4ZIQxUYbooyu3Tf7de6BpM9M53pot8WOFo8fir6ccg/VNOZZ5quO5A7qG
vjHJaMkhKc7Q6hRgoRYor+yXhgkNqyosyIer740E5l/xOMz3e1RDQ1rq766Hhu+Hyx5SydzGomq7
59dZ4mQZpiNL8lTLXax1M8esNb9ZQS7peTAvwJe4NbrUsKxR3TJ2MWgPngjARTb8ORK3lYR9pH9c
/RT/Aw8jAjMhFBdd9vF0nXPuBTANkzdnrZC/W9OimjHOaW87hLR/gr22v7lfuINv3J0+8lCMQ7AJ
SzzSAb8kdOfG+J4thqH61SrBPsPrh7CSTOg2sYv4B3STRnSgKwzRXT3tk939ZFP9RexpGQYwenCC
qqtVk1JUUVazavmCYrVnSRN2c5SR2roXrVS+8qAsNAoqZn3O/nDsJZrmOGRhKYrB7+sFLGsat8Za
PcPDlM4l1m96koaKGrNe7d7c6UxxRMx/h35rfP1xPST115Kuuh777CULJn5GNpLqWgLeGleFIX1C
lXJieBDQAV9OJnvvhOLK5GiuNEeEk3Bz0jzHDNfCLaRM0VtgRK4MiD+GHvybeFXkP+uqPOReo3qy
iTLoo5UtBj1qcDUsdBjd0B6uLcN5AA4Zk1kancaYY50QtRCIgKK/xY72rz0zWgai2/H/z83gncMU
/p3RIHgqeOPlOOyLMCn5MlaIGOW4gwc4nR+puxApn90u4RJDvxbLwRbT/XBtr6fKjNoIay8xw3SM
CXbr8d32angcbNCO3A6w+AnRb9Ri1v6176N3DynTLB58cDWwadzFlTaCItiuIBbVHePuDHU7U/25
mUbHpdhGnocKavMZUGkkoVvDvRxufhNy7bJwKNTbpcGfWPcIBVZlbfhnt0kv2dnACsdgJccPDgb8
QDzQzU4UklwrTeo0UZrE03lzR+Gofky4iH1ZFONzMVlpXy7ghU5va8+lgwHBbv9RSyYUe5r70Gqd
e7MA16jbLX0XoF52T2C9iRi8MO0TrCQlwLmzxC4N9ubAMtLDhKG0DT1YEIh76Iq2iKgXhifS2AUt
Kh7ZbYMIUaEznJLs0/x0ycnUWqOfAB/tWwoXZZt3yGQDKziOI8BT3QrU69p73u9Y5zXczTWcUg5n
rrQvhU4OvNxeN6iixsLQBM+FQMmyuI81saQVakE7MVSKuJGFMGAzagBCMGyDdGQRfS1dHZm+HmC7
BJkWlkrCCuNNVRWsqUNTqESogivC4Bug949/w/sWdtQQCtqHZ+rMEiEckW1C6G+2R6K58fH0Difk
u2U1KfvB7PRGcVUjkQVTnEs6T/2aUBgQi0Lo6S3NmdPqf+cPNA0suTAmUYJRe8Bseruuk1uBl9LW
FUMPfy6tNX+Z1fCG+IvI4pR75f6dbQYxIygrHiSyOpLTU4F7lzRdKBbGFy7lMAP+GqS5TPSwd88G
NEj42fZriklImi34HtnfLXwqeoP72bwrDS1/QYd6ONzaPhUil57EODb+m/PQBZfCfCm3tezjv9uL
hkyVnVcrQnSBJtDJSJRmTz7/qFDnMosgk7At2cPVM4aCKbAy0aRfNMNtXgeQcE0nf/RbE4rHWuuL
U22jxMTFdsNn6pismXEzl0bNtP9L8B4BhPCJ57UijD4EDf7DMXou9khp5kJ9ze4mf7nAmDZsqXax
w1LT1tpO9bZ8TAM+pcm1OGkwk0HmoBj+k5/Z6KCX1g6xcEF31vu+gnQXdSH5eev9BvLZJRZWoNVB
pCnitl09QKx6g+i6KOVaDWh1rggP34ROmRh+YoDlpMKY0j770n/1Wry3ucU/tk25C4NSa74eUl/4
lp0ly4mBBw7j6vnzUcfZg1eaTe1MmM61EVox3YtquMoYhNUX2ND4pOGKe3aegwbHOHuWQHE9jDSs
R020wHFa+cTgdC4Tcv11UVWT52jNAzlcD/mS2vT418ZWxwjcO2dx7BiuSzffL3fK0vM3NGaL7Ng0
pyEHmcr2U2csLbATFq/n26xFEbDnHvKj0fDyocjYkLVhuCbNQEtAx7p5jYyXCLAYCEzgNYm+ZAub
57+vVCB53vZEZ/UycgnB5f1Qlfv4qW7AJbCk/Wq5G5mF7BmC+Se5C6QJoucg+YopM+UtAN+exivy
CLedtU3WO+GhN+q98P/0rbnE+tZ9gZF5p3TkYS9wpHC03bJI6C5mpp9MK5m9xroK2k02DZ5o/iZe
7WzqQ6rTeurAr3CfyhHQtuv5evblURFertyqqyEn0HV0cCIlD8E8o3z5mp27gsCO9mPSZTY+T6En
x0yVXwLTRsnxNZt/XGfydE3ud7jQQ3RcgV/Wc2o2E95BIfOO2CkldSEUUN58laFu3X44VqJuHpXx
Z1x5FAMcCNW69x+qEbq834EPkV5DIDufWlquRN7njKt8ob2Hey2g5uduV73VSzsAsv30AJPhsfyJ
Qe0iL3FbZi2BlKzkNFHYi0i48255pTDvUSnROiTUQvH3eLUo1Af92X/ODHbUsajggaymuPXn/jIW
ACW1zxn1LCyf6TAM5xfMkhXt8WDhDdWolWahfrDZiNYL3ms/a4+Dlnf4hoyfuw51qBfjoJjRn/MB
zo+XOP3QtcN/t9cXDoayfStwHBsvWHR0M936jfwTnjmCNfZpvQ+W5pgppeiNhtgG7NeeVoJcf9Ks
/ERsUaET8qR1cOyaOcYp59EcaOZjRKqhUogbgIgeLf5sXvgjQU70+ExVxyJ7Zcs0Okuj2xyKE7Pg
qrUIXPK1PDdGhiP0DoSlnaBKKqKuQjs0LlFA+IaXo/f8fJ+ilrXBOy3zBS+OiL5FP7teAifuPn6T
7V5ZZc4N0f+1pPbHyBKQVWEHj9kLZi/S4WsoaHpUdvFPUQCFBCzZ+H7GlB7EVBiNZBeMC+oFk087
07pimhfDbfHSzYBWV6dqWwYtTIZ8X9WxMjqyoeu0KKm7htHChmer8vl5vWjqxyKuwb6/QRR8Y6Wh
Zedlcwn3xn5lE168VkgacFfWfZJk6hu5HZkn6uNVgcKwLKLQfwCBheDqcLU2KbAj9T1YpG6z7u5P
GFPcBnobxnh+yBl73erg7UevM9qhatTqvmeI14wXurBdbCbLvfmVDZYpDV9Hn4T6kIIWHb9R1Yg0
48wgVLUl/AdaRgpMCjCeuyx295p6lI5RpCN8I3h1IbSZZNSRXxRht8PUsQhiILXil2XtqTHGX9zw
DMt+DyP2n291c5IIQpew4eKpImIQYV/N7wRfZ479eu1ed7TxFHy6plqxB996Pak0j98E/PrNdsMD
mU+UMjxETF+Q55U9jkJ0OLmKlnUarfbgg1Yzf99ZVAZOTcmchAARQu2hxOAk79a/UEAftc4lTKa3
daOOngeiK/H5OFPtDgYmGvKkGLv09KO2NRJkaqrCCapm8WPKdFbI8km1j+uFrymIHVaFnNJWj3Gr
yxPRamprFlDvfVkMuytPcb46xY4G2Jm+Nkq75CPk7RZniQaQLoBBk62U895EiESTM9IW/s1tUqhC
4iGrPu/2jTYOgIHg7hMxBkKXo/86Cw3/5y1uo66HJDTiZDWNiOhFGMOlasHVx74hLqQp4212Csob
rQIEoaaBuQH1GDXlGZ2f1blqQFQAIKU/T5EAeZiHAyRSgkPqpXyiSOJkyAQZxkWPepzCZhKV8/Ha
OJ5h/MiiQcvsRNY9dldmAfuLZfOYQkkUuozbX5Cmbz74lVGPucP66R8C/nz33zkYIBhOOo1cPNIE
u1by7GEuwosbPCmrEGHprbTuz1XSHLfj3pWJT0hhDNtMvYcqGKm2OShXA/b+MaCmoqGdahzbm6/9
A2Z9e73V0mXnBEX503MTr8Swe7c+G9k/RJZjZyjsJR8V2/fYvCcnh2wWyj9wD+XdKpn0IXXFPorG
i5J1mJ0qEokmaELvNh7Ch26OwN4Jl/f+Dev2E95AaqgE/IIM79Obe/oMUawEDC4DEInfYmcRf7Yb
Pyn/mLan5LK5qQZiZ6rC1Ftt2jNGM7Z14Oo/PRYZKLU8w3FCvh6JnyNrc2E+Y4WwqUFlH9uN0MJC
T2uWPXfQienVnHG7nEpFGBYhw00DGGsye+i2YwUKiYZpyTHvdJvUemwH6ZhnTZoXcMSjaOKp3UUh
YqX4DFH/Ncwx2L5N0b6K4r5a17Hv+yOLgDry8Q9iTYBKyyVI9RijeOgFq3uAbDpkavAiHRf2WBvG
YUSjaoVPjnb5SKf8RJVzwAC2zFoUqJDYZ4QFV3ifvQUUHF0CFXtWWpPTz1uGKMp7jifep6h9u9CO
tyFQdDdXwocMlGP4KSMQEGdsqhtlszwrfjXeVxKMwx72ZxYnyE7mK2+MzZCnWY6UKi22irfDwj7R
GjF1M6njS+tD8KtHT0PlAdK9ir3DFd8wK2aKB0UY97N/FAbQKB7Dju7y8nN8lAYG1Ytig82zQiqN
q5AeqNS9lNvqfHXHgvcR8KjTT0sxooHX5KK3MIU19cBt4G2sSCmdYWwe5SOXOdJPMs68xPR0MgZd
Ml+ZdEzsQ5EKJN91q0BnBvcldWiGxIfZFoqj5jUZxPTE1PQA9kG/uVyqr8PCi8FQ9z/v5KEhtS+V
bTmjm8mYSMU1TCS7ImatB2ICyC50Qe+OR1WyDjSnlrPz93zrlWypltpuS100IYEGumdbX/pliabz
XnGhpSWjR0J325JtGkcsnvyE6EhdjiSYFTJpk2ZVnUkqI0EfNWejxEnSex1Aj7ofzPHvNJm/jgYA
mXb3q1F51bOAU9z5Kue3a0kp4SlhbejzlxetiEKWhdR1o9VkRJkHljtP/wkfUlAT0vrr8F4lgKn6
LBbT1AiPVXWRb9N2f9QMw/lpc2xfzql0gUBOH/kZWfGll9mFCs9RIvlhkOvbyGjhdJq9/c3MchaJ
/K8P14ykyrLzgy8bxMfHcRxbjoVA3XCL+X/88oyE4lVTc2yZbggXhNZzSwKpopq2yHybmRNsLTj6
3K4Nm8uNIueuz+vqulWobem8wy/Sm4hm2PLt9n16qxwMbNwy+66sJS71PtqzBpjsQnt9zfi+YW2W
hrxLYZ9t3atJP6f0WgcJuA+jMTaJvabfJ+xZ1UjwMpZ9abHUj5PEB1Gadh4o642jyHhBgvoGd1VW
h0FUlKOO/ieWb0O3+cPKlhY/T9jCAJnpqDdyqoFJN1UeHoBcJO0O5CMyULK60/lK1Iq/fV4AuoeQ
H04VZmdZl+yt9l9hG/+QRp2+WZVeH4i17Q4MqZvmljA4010C537HvZmg0Dp3zNl6RLY/IUtdlvW0
mt3zbO6ftCjQlsSUzIiGLnEGp9sRA/g3ZxooswaLhrL9F1BJnmisMc4aQBxs+n4Y8u30xJ1GPIv2
MFuhSndoo7Pn5SGKo9jkGwUZ2IOuM6rTzpFre5oVtgROVn4yr+A4VfAey/wLp5JvESWCEfxIWpXt
3tAqGVtkjaOJJbhcd7MQcGnxYymcvI8cZuNwzkx/MQTQEf+SGSGD8fqqdq6fQOu4TOmnIqerHv/5
2eC4g2JplQDfPQp/eamibGgXAxFaX1zx+Bl2l3svwiv1OQbScwI+S9/FUjZiY//RU4LUpP3Ztpv3
5/L8WmV6XP0TIx5nkPXEKvpxOnSXMFDmTblbrbYguwIvjBZpnCxFwoyBik5KDsnZdIgqUPbeLdc0
BKPjQz1EipAGPoNuYQNB3AfoGfOFWPVr5BTHgRiEaL7bdWvxMXWltGuHFZadJNOI1m8H+jFh4TPa
8ATD5784cmUuM0lvP7JjswQC7IPQ88U+Nnv+Ga0eme81IA+rl65QxCOFW1C3guWIkGvo0tZLwJ57
PsFJ/KFtETn0UdXSBeVq3jQdVkQI7SUvRyoxRCRktH2RZfGciVk3mSBrCWYHyvkOXV4jXbBMfIPs
vqBjQl2XucJqAy/C2LzC9kBNOCWeUVInl+ahJeiFAX6dVVgi9TK3wfwE2BBX7bNnudS6S4k0Xvq9
DuWXGoMZYYmwEq8/uHWRNaxhFtvDmJ+M0zJmexBHJG2QiyJvcHTvvULHCUIniootxW8uCfcG6HoP
pU8VAtRAzAh15My+F02Qo8TvM+3S1/m2ram8RbooBCsQw9znOkUHYuw49vj9a2GCaBQ3LTLEbnHS
er38pECd+j5BxZgrSxHgjcxxTRwi+YOo08lH9XUgh/KTEVuT+C61eGWpCE1jTduiUreheSJL89bF
TAcE0Wa74ncnxwTAuHKCrn2gEhz6/3sh2OF6aazmcMNLMGQp9APK2zjA9hhaHoZlY4KF8JPCzPw6
Z+ggYyJPWs23gmaZPp9VDg1nx4YYOxmy7losAIVUyXUQiEmG8zlPBbxRVni74Gvu41r3K/H2shYs
t/tbGnFDlcyXwid5RIH3skg6hVlDSeZ7CcVutA1S3D6N01vP5ojjP+1hQMaInn4O6Fm67++HRHuP
pzzUwHVJTVIpU8FhQKeU86xLE/g7rrwJDVYQ74l2yev3v0QvGDJamBnpN5hjIiFzsnFZYLPDbchf
IPCsH3hCbSmkveYIopBcT7l9F3ABuKUNZ2qAaW/r8NkT+gzpdpTN2COTFt8lpKbPR+0Ws1mUHdJ1
Kzp2R4/jFidU/VwZ2TNOdTwLJ+4RlWMsRR32ih5VGnG2uzNfh/4kcGCGFj6jLIu2XXm0oIQwOSRF
NOwlyA/7ttaQUJq1tX7OkdRPlrgpt7pc3OkYSz9Q7VNZGZqep1tJP49T2tPSTKkwZs83UeaB6RQs
UHVSVOxN91Xj9GAegUf08lkBFGbZmGLsCVmA0iKDbnQmPjC3AUPrR+68CankoY48TRdB29flDqNc
Sz3o6ZNkDX0wjHbngzcc5OaLadxOglaOJEw3NK9lV/tnolhPO9yHSLqIUkrGfFWfJU5v1bQt89cF
s+5PjE2f4KnXGjqlefvAAW4Ff78o7kT15YC+tsbkgRnc/Gz+KtlimskvhTTrakRJzTnxs6Bc8tvC
VRr+SA0alusctGkK4sMkch4R2mXiFiO8gO0MhNmzSaJrlY50BBtLd3GuJafh8Y3xAKtPiYDPYT1x
JKx31r4fXDbG+Wi3zvex3cHVTDGOihUDF1MqB1ftMegobXValHOU4MdhYjPpSko9Q8rj+LCNXCay
Ipuhd9pDUF4qm0+mHG0OEaZkXLGAAxXdNATAZjGDjGquoQpKjCFrU5uRxixByNSPOQ+fRrsO0zMX
+cKluDYcla/Jgdo6WG/K1Oj4UIhhTOXR0PV9mhimqdkSGQBR/Q00PvPlplJHknfWyiV5lBw3hGSv
DaZgLVGw61A/B8QiMPik4QukWT6gzakp5vAUaMh/DdWCnLDRO9RZmXZwz1fCNhAyHWnzR9lnwtMM
dQ9ca6y0gCJHNz4cQkJ0QqpFAyL9YbtCAw8Oq+1lBOKPkD1yJ8BwmsPyW8hhmYA2w1Mu+O5hHhdB
Kg9TUTvHCE0mwvKCRVjagunT8ONA0vSt0QBmZ2GG0Y4qbVvSxCU7BWuepWNPeBpAaik4Y20jF8jt
bqk+RvwywgC+AkrF0Y/m4EHkxVjzmyyTz+oH3INHsxCHfBJJxSa26/fQ3sI9Dqq02+2OgNbsHzsE
SvIUtoFCAPjyd3g2uHK/jnakHMBLkJJBLIuhnuLpaAw9I04GyGl9MOIW7iJSU7xryydfrF/EEA3l
zvV27Hy7j5Nzad6LgZtszTD4k1D2LRd0B31X8o7vI4zfY01wy9BuEFqnlVDKn2B9cjUz7rvul2O0
o/4DRHBdc2sgcUSOtt0BZ45To/9Og9zg3omORIqFMiRdNhRSO3e09KyOd2Orq7rdHnStCcwWavtu
L/vh8Fn4mJaB0bnteqTyv5ORD/m1IIOLtxXjz1KDS+Ehui734w3CWRUbgBH7+0FymN6YTm4oj+9S
Q2LD7SSYRMqs825w9BJjIBe6gtcEIhDG5EPGfb/f0sVqJftTIp21PdLioLNueN7AlpW/l2AEpBK0
JgWUhI8kSzj4o174BmwdIHT+cagrz1hbbOKto1r7KUYw1sl6hyX8RP/zKr/09+S9R4aE7cZtdWyp
EZcEFM3gpK18l+GtRbe+xYk5jg4ebWoC1xLAvbdQVUBgSxR/A0J2kcBZYGiVg2y2ypVOt0q5QALF
b2lmHSqHsSWH9nu+w4vBp7C3W/WMF9QCC1DN7PX9o/uJFMLR4494PpHJJOe3aPdkIuO4bAEh5SM2
TxoWLWkBeK8y/PMiuwRtgS83Qtk5MzxGkxRv+5/TnS8fdp0zhP0u6rjDWWSMyRllHUxS2Ut6/UFV
4MHQcaOXYKW94hnYVhfoihMYUnl0sVzSSrMyYEad8jdiUNifEGJCWZmxw2xl2Gf5wfjpzDmcoCyr
wauYwXxi+//bVLgvQLO/WyxkucuuqobQmaCA2ZoNV2dL6mnXACPvtwDkd3CpVJlXb6wAEECL5TVC
5p0TzjN2hlMg/ELDw0VpPoeJ4D1VANmawtcLDe6IrXYskiRpAFxg/lkfxHAtF4TR+INQ+4LZvphO
6E1ixF1Ltfe96wgJsxV+tJshWQuiSv18wvhq5up6eIb9xphjzdHH+/sj1kjJFQf++pgzSNyNOjKT
b4dkyuiA9bt9+DxjUglX1+ZR+ob8ydNViXQvmXkk+taoa4upqUPzHHoIJiruAKla/bd7GLetO9vk
08ChckXK3RZYRZkh13XQ5sidG++60A+qv1s/I4Ky4k9mEmrJPsZXqH/hSRIgp1KIjsIbKuP4FBTG
6yWv1nae8uShnipM6oHd3I9qpGy8W5vPXdp9DzcLbZNfj7qxez5wMCowTzgSjMXCi8qCe7jSt6Fx
8Y/NSR7jyYWusIvGLEyFZ9RYplbQ04ROm57BhZrRa/LSzXI3FVp+twoirlS4o6n/NwWCNog8rP11
O4mS44JePGFxFXwa6TCbdTLVcUj6sLXIPh4kjOQ8gxGI4gT8o/9WCAmUFU9KeqL51cG9C9UE8vSG
cWAUA+zk8AW3ETxBjkPv9yA+P7oV6kNruEcF+K3MD7V73pMsmLIo+fE57Sn8N77hnm1x8zHnMv2m
+Cr/2CrAs2APN2PHYHrPrZ07juysygVCM8209bGnaUBw16TCuARVLGGFiy6waVAp/r+eSOHbljNv
Hv+LUaUsGOC7T5Xinqyb3iPqIqDBb9Txh+ULZO0CDATS2EbmmlNnUZLvnDKlEK2YpuQxC9hXf418
qNAR5dhEbgOKxEkA57gKkwGWsooA0Sl7cmQyKqitu/E7/3kSZq7z/ZsLKy2zRsN0YUuOBwU9voLT
ZllHv7tWA7MTQSGkmrUctVt9DT6q2kjuiiHn6hXHhYZrq52L/q6EY93gUlHfzN8/Dihj9eu9EXZS
Vc6SNtCHa8hjfx3z7p8KYGghdsGhyzJ8YYM05wbs0XUqo5/nHWMRisFE+cryFpGoDY0RI4r2vzsd
/MQLLiunLdfCXbXoQHQyjD1+3dOWatuLwusXK61XOgw2l9TBtv7Iz/fkylF4JkplvXH09LN0R6jt
aZjoUgJev7KSs9CtZHlxaSFIWYmaWjQhtOsGMlF7QM+6TMQMqXX38QcrK0ZxbdCO5U4hAfv9uDRP
HVjTdSoTu7ogdviCljwMh/PVXDzPoRqW6GGjNbXhGEKrSPvCs9C2X5Dc6QoBXsEvkM4zr8jHckQA
mC9oXXoXTk5EslWtzYuKiZfMzHvSlp8yXxHRpLfLV+5EHLQsDAM3ODnaA0rUTUfQs+RMDjas1YFp
gS6EJ+mdr6ebFWiU2lAONkSoF2frJjuOCJ+W+3TAIySk19UDIIdQmsWmUnQvfc/D2vfCXQnUMR5m
vrw7ceiVhylRNd3lL1obGX2Ird/C/Z5hUgP+3qsRkIca5A5PEt5H8INJ66+9aEqi/jE3yQMny2+6
lIxxTP9Uhvs33bprrT1PqnojzkFz3wvU5xlZ1C4jWtwksmmI0lXuys2s2F0gGm4T7YsZkdNQRkCo
VYwII8qnN6u3+H4XnrkEfatD1Jf1RHacQGaB5zkwY/H53SRWyj0zlPhpN2JfhQWt0bVh6ZQtdC4Q
5JcIOun8CN/UkYiFTwfGQDbUxYVCf27ULBwRgL8cahZDaabMgKErYI+twcQnRV91tHoKFklUECzk
djjLc/qU9UsRfoFPcN1N5GxJOLnMrlnr6tNyru6wijG7g6QY5O11P8oLlWayY6j62Lv2Qxq3eNUH
L98OX7PNMmIxAH1kLWu0ejhS1PMDxsQTUZWk9ggZ2Lw/8K8DymLEivrMrGdnmWwRbWpbnIQ89kyI
8oZLCpFNzTCXRchD98Fz1AodWsW6G64Z+xb15/YxxcYzXJQiquonlVBRhHFw5HTMKK33wNyIfhN6
f002zVVk0ppC0j+4g/5Qht4VkyVEnrPhe+3cuYN9cjdrU9N8CcEjwH5ryC2WbqJ6alMaV69V22Hv
qtC5Qx9Y39qAEJJvJ5jLAdVdIHKtaqR/OC39PCvwnBzaSz4T38RAXiS8bPAVt1bmBfMXj7qNj1zQ
xMGLX0xx+YPkEXbuK+t5CfeQ8W6qCMjN7Nzy4DcOJ9rJm6//uM2sgFmt7HEQi5JkxrGEd3Pp2Lrt
n+QNYcc9Zi74wEBUENDSVHfr+SCt9RMPfX+ce8X39evlnt8g+eEt9jlrtka82JFIOH/yLSPGaiBG
qgatQHsk0NW560pSFjEFBoWxc0/04CwKh5U2edFN9aNpGJDF8FZurqChLQtntPQjosISwEH47KOv
bQsXZsSUghS85ha0ZNFgfxNjeR6fWAXT/sp+9dfRwiAux27K2EpvmyisCbInIUE7myz7pk/sNGYO
RL0v7lluz2vOT2tJvVRM0b724O0PJAeI500WBZ7+4jnfo9CHfHQrbO2qhdf55pgMbwnkN6LS2quR
JA8vjTr96kJNUX4v1fDX1ndFAHJKKQIj1kInnLJo25DFV+Zbf5QPWydBSb3kVnh8OrJ9oJmnvQZ6
ci2rcuRfMC5NDrjpk6ZieVMyPFPnpqR7ilEgpGgtsVdZkyuTYS4L2aan5PVrDV9lLi0nmmdjZSYc
l3vqZLRiuquLlvrQ/UiWmQMGJBrYVDKl+io68wnpl0dISNlR0dQrQ41l5w1xFqkAqI2hHfi/5SZR
vuCGqoNE9S+IQIPvLB4rwVcw//OOdk8fh0Xb7yIQoXMmbOngCyPHdJBam2+tEJfCeMrbm3LT8UU0
09aGXv6Nqd982vyeH2vcFTlTbIVN7DMaPCpZ6P75uJGP9rV2iwG6uw/qdjaQZzoydbzanLLRGhN6
pwjQAH+2Uj9+2rBeeBrVXJ7FB56ucHcOHySl8B/4KsGA6dAvStmm9igj6zkl6ulvmA40zBVhrqBK
wS/owxZgwxcSeLEeZgicI9otlMHFHHkBc2emLEWiEnnrOB6LQP9iJm4wgR7Pb/1NizJA4vnMsNK+
Gso1Vlbj6VPU+myc0RnnXjUkYGHYGd5lY2vdg7F9p9sYncAZ1YQk00Gp0FXh7YqzCbdkBDC+9JOV
Y7aMPV0+HUgvKXG2ruYbjs2Num+KAMKDTO6ybTk0CP3uFKPug4ZvJNKTU2VYSMqEXOEeIVpdEUhG
uqQ1lAmthhDSO5KvQXDuKBfjenIezFaTyt7arlEVvs+AuFjVtPv+Gm1aj145tk51wWROIhtQ4L9W
+voscDrBXPZs/bCP12EMSiD6IyyoK5eZpOxtWn/dVfoaQRCeTym2Ad5/4oMR2hFzYLbO0XE+pxlC
t6K413odd4GCgp+Em08THUZMZ5ZGr85JlKr/ELqh1qIJ4TUlIJeNH/prqZ3UvFutxfu/XxWmQKYw
kAGWcWWfkvwyrYN95rgKZsyJPzCj9EeaxLXDsSuiJRWQ6k1Rml/Eg+DQP9tKQRBM+5pMrYW9Wpka
LseKzesgeXQictwGbUG6L4pskWmynX9dBNpdnkcPCQno5OuOL6lm5WHmIUaivlcJoWHSIfSVv39h
UzDKmpmyExPF8elEgoWGnP+k66NvC1Ovbrk7GCWDMPSFEjYaOKymOZuawzZKpGwNc0S1tkTKFAvU
ARbmhfwKtCUXCkUhYFoErNdnTuX+VROwzbATTkaH4936Lgv7STRlnRR6ZcPdRouoSBXfy2PeON1C
AwraSLReXYuhy1FtQgcDUwDxKoLbwfSbNb/FBC+RtHBbEFMoKkET/GDhLfYgWvW5C+SPFBpbg2X9
lael/tBgckTHux1TZQns5Wd89f/avctWfFR7bGTaze28JdGVcXSobW2xVlsvb+ENNgDk9y8RAs0X
CwIXxrIHgDtizwG4hW1kSHslDnfDrj7t5mYEFX0ubhZ2ZAiPD2NmWSUDtSrLSjiqUgEaEbZ5cs+p
znZZAVM4mU/bR3XXB/oxGvU56poI8jpuwTZ7S7/GBTUUYDhCStTiOki8W+FGi2613l10vRvfxaV2
krTQkiKUJY0zsXlqketFnznRzCSuSe9mQeUft6pLe/S6F9j/vBktOigS8TOpWL9/w9YOpcK7XBLG
qCQygmaS6Igth8VZoRSkCbxjKhJwBWQsaTUSaQj5BW3AV+cyBShlo1T5CY3ssnSMUxtl5IDFzVAT
hcWvFvrJbyQ73s+25dL6OKrsQ6vzrvCFCAydsP5X4Yb9I1SCLo/rTMg+kZ7qQDU2IGHYK39S/fxJ
dFQzc2vO2f8rZYwGdJpsP/W5FfXoS9K3nfu7Eu9FqIvAO36PlrC3B9m+kRywwj67EZk+xmZhcp1w
txY09wpke5SfqvoTx3mbHNEPjnOxf7W4RmyebG8EDylOfkDkFI6VSXZit32iftPbVcOtZIwTzAQu
mOiIzfrA4YWkbPH0IftqsK9gbtdymwUxMUUGJktm7FAZQFyUPWqlhDUz/XDsqd93ZdSyoGDrzWG9
L9ZN1yDLZbmkO9RWJ67ZO0QbE2CEMKXoDjowmGuMmytemWWg+bPL40QXWvbXHWHrGiakTTofx735
XUyyXOrUBefSB1dm3B58K0QdfLJz/jBalY6JYl7sr1LuPY0hAEEzscwnJYMFiTMnc6ixN3YMcWzd
SUk2qS+kT6dAY5dzlnqfaX/FTYWGATOLQ6hKdpOmQK/JDf0Wm9J3W+BlqRS4AN9mJIdrmonECZLw
yXP6z4Td1mAPdUUyOySavmBJeqJGSZwmndkVkZwT/gmZFUFWrbc9JzBpq/N8zcV/oINuXLDBaELC
laajQrKc62xtE00fH6S6m/MqGZvAxPH2b/7TuPbsGOYdIRdNr/mGkd6qBOLGdJlP1CCR4g6s7eCj
sZ8PHAk6TsO21t2/VFYZ79qUZ+7hF+J74xbMvyTyZzKF7aDHFBxE5Kv4zSBZvFpVBN2VALXl+zw1
Q7cLV+a/FaCuCE1BZSpuXoCrZNR6+jIAY7fVuqoCkajX7TEU4Hk6m1H6ZrGVV9rGItjVZtxa9XF0
XNJYtfIibJgPRA6ayOyL6nzoHNxEUw5W3b+nFwtjE3vnJCbnxljE+3nJkkRT505yEWEtWA+KTPGA
/dHznJ7O/z3OMwMxtbmyP4d1A9fI5Ir259MlAM3/p7RlWJOPr5mOu6qz9SNd22vle542XbLkn9cO
RZUc59EXV5CVM4RKAi4Rfwbvb9sLdG2uX9CJcLyObqF2avUX7BaYU96yIGOuopZssOTzw0BI3W2G
09MNKq29IajthhJ9qk2iW19f4Rf80T6VJktpcWqwS9JR6K3e8ZmDGv028tbGyTNeGJobT962q8Yt
NtputunTU1P+8KpgBFA1B9B8fVvq3Gc/aI9b1jgYeCf8aHANdGr5BsCGML5PfivSpf1thQVetx2e
mJ4R8hl07qhHQRRh93cY82BS21OuLD0TFpXco3X2dBtxaOdA5W6ZmObxjMRUMms0evvlu0JEMo40
yjgTBqMj7nihd/VRZ5lc9oPD4gkSSpiNO7AGNPhDBlpjcivC6FOJNAhm7rPxHXi9SG2ZgVhdoZBf
USKAUBcKa/BSnjMyhhe+FccCpsNsZUMxbZfKYS30cEiohPBHaHuaEj+iu9tB4KnonyxtSHblrYOc
1SXjJ3agiFWuJXzSmWehhbqY6LzHmqLzPUQh47WsJzKeh4ECdJThStBtBL7y7VLyIiBunD0Bt+Ki
NGwa23vA1fmQ4qm3BWSCLqd9ijGXkqSCq7iIdtj8vTnkklldk92tpK4l2A3SOD4CJMtg2yqHKoAC
ij/jFptPvsCArsMptIfo8DpwpSr+70Dc4GdBo9pf9c5gjNpwi+Kq+nU0ArlvMzyDZR/6/My3OG1N
dgVdg6aul6evzEHlSouAwcPupS/iPCiTo/6/jTFwgCVTRdRo32bRbDG0DutUrkchHpFIvKzx6fZX
4ulBVvgmsbGTzO9l8aXbVIpOKHCviXIvHRBBgqohvyeUl+L4eAuvYqhwdUs8X1NqL7wMVIF+VteR
GDcJuL+y2JrKoO6o271RHj0DpFTfEn6olnykCK3DTVslbcAV5iDb2XhO6dgnnCY2lkn1k116Imfh
dMH4MPSil/HHMjevrqQSpugxxDG0CYL6nNsXF7KTGQzHNevhSHapbUcFNY2nPAElyE9f8GPNlBUn
zVMz8obK2JWNVXDzzxgEwKz/MxznPDnBk5Dfz4+L8eG/SKTSz1sQOB0TcMvPIkdGkKNdQvGWtlpO
iekNPPECDCg2ijhSZyaUl9WmQAhB3/mL20s9aSUjh0A+yvnvfJtrA404K4VmB8sjxELduj/3xxIu
a/XX82oJzWsEc/YDCDOk9XrIZVAmIHKvBBUe+w3q4hzPrY4G1bKNOrDnfo8RJz8JFfABSnMAkBTc
BjManij35UU66TlRfK6rquFN89Xo1NladbZCmD/vLkfKthu+Fl1Sx6CDOxudVohcapmNRAT6SSYQ
vzvoOUAQQznwW1ow8A0+uZ9I813DK7xsy62RTI2RzotA7IT3vUM4HBlLwJnfd7Av0/EPgLpjJBnc
TLI8Qn7qsyNTc5QZHgWo3ZrFRhZrfIplOdsDjDk3/tJGDX28jPkd1vWETlsVyBE0uLMyq+mNxYVH
mRnpn3N4zSpgMb3xm8yyJ4/J7WL4CYeNo6nYl7xO5HY5n+UbrrTF5Fddtp+iir5Vp3l8b5fzbIoC
sTROoVRsDKa8qvgBXFcwOpABDsQjxz2S32fdMhYZAc/wPaRKIRZLoD26B8jgwdEamXXGZd92t//d
IIESmF3LItYklQT6p+/I9NcdLk+IFMDJvV5rq/+8/KoZaLQIUSlPtAbF2ZdvkIdY+wAj0IXUbcsR
n+6q3CLlDuaxptUEBkgqPnRJfroruBJ+TVd2vJrDZHRakYByE7Dd7aCgGNUh79Sigq4S+ebtbEk7
M7nAAsoWp1J2SUfZwBOwQkMSy6iaH20dXu4X9D3d/bM8mnMbzt6awgrj3RA1OnxA744FG1mzCxod
4yXXO8wEVV2tMBRgqbuhb04XrtBqWVb6NBN8oWAa26oF4kW2rnEOHuZMZ/+OPcZa83QUgqs4qkMG
1tyXynHZ2vujQMpAakDrdYu6vOaM17V4OIpS91bBoFAAjRQxZoxUB3x9gQWoDmkUembEAw8wiXAF
OXloRYUWxvKg8nufUrbli6LRU3X4qnAQBhURNZjHT9Rp2z2RCyBf72Ff+eUwQBGah2U+cqMQEXma
UKiGZOLTMHqdEk9tvfgjMvDu89tzRApbg8IM7M7SOirixNS47/UgpkVfhkRx0J5yg9gvJeNgDAf3
YZak6co2vaNPv6YylFa1cZ79FqKer/eD1wJLK9xMfrmCXYjR2oYP74GmQoSeZUIMnjj4l19CO0oM
+DQVjs8p1NpTedtLmCRjrsq1vCvvE65SSMLecP1RxLEcUyE3shbF52S9t0xzO8KVrE4gyGlSWe/c
S3YXyCw53fd3jvf79u6RWykbaF3mmzXLEQrr8aCfqSxEp3/rJvygiAmZsbQSTJrPKHh3fDq5v1gR
LYl4MT/VeXay4peDTfF0yUcOYIqJfzsdREO8uTNRVq2uWH8aa5X4zBgHfui+Ker/blJ/H4q1X5IX
mjReLALuTW+tgratZ3mDucVS4qrKcUXhjdMuXvIjnNTpFZ9pV9eBoGx4gVtX3o7ECQaEqIy/PAm1
YEN2nA1H6ZVox+L5PUPLBAxQDAMjtamDSISgqW8Olx15pyBr+l/SQOwTFKCs4fpAizXve4SQzSbo
2gDrOdoEx03dZ/WQEoXQWnY3xfwwF/4FcgDLUZuBnw4TmxacZr5rQ/jZXJWeHAQAUbDdq//rsgLp
D4NVqyCdJO9StJnXQSK5iEKo7q06BPLaRW3BVI6xKiMGVeVxNMEYBFKqnq1kwHvGp1fj1P3TdW+b
sgZxjL/8HcMR0w2wMskLlFo1hznMROjk83qx69wPJcllTmu6vNcGWBxzuZNCUjPd9h+TF5H05fQ3
7PUAKJyr9exsEYzNyrCZtI8LO6bGiJSd/3a5D3a3OEDYgdGYBcxJXq6cyH42vqSEzpZWZaIrbeku
HyMWEVONLh2xUxsdpLDO9uUWAmLgmz/vcli7m4yIKyibMIqpOOytWWm61S6jwXGWkmsgeAyhn7P4
bzb6NQ0FwMnnL1tqaRHNZqnS1//wrmePUdPnsPdJjgpvbMxzijVN5W/Q6kHv4eNrkqB3DxA/a3+K
ake411v4cEalpHVORhD0Go1c0oUtQs5sDnk2rtOcvN6aHBy2ojmGbg1kSeWvT3EOzV1Mr7IElirG
UjMuZSmXEUuLw9pJ6bmT1J2TAQKiOq65imI1oW7UuOrEfpcQXFPUs3InwPAldsYQxsNOMdYdrutN
lTs0fqCile/m6WA9RPxJPSV2mHUd+X7lImT+p2Tkmm1VK40qRHia+yIxtLEyeuYD3fk4oik5dIVx
i+1HYy52ZHBibYeFXr9TmeNzNBamGpH5wxp940/zBGjk/5kx+gWmWAJn5D+n8wR0H2dj49oKTOMh
hJA+dNi5MvymjhP4uoJSGltrpbMm2sIzdn/ECeU4pdrR2XzQY6Huyd6SVR9FR2VMmOq5XcxT2XHq
tTmuS1QIS+KiQ8myxUPmvIB2caq4xveTEC/dkiJP1cgXbTmrBY/e4//LEdsWq21kVaMIDx0l1ESd
Ss0HIymyw+keYY6Iy5rzk5XQru/jWJjF9+3azNZpibYc/KTr9Q7dVLc1MI183ng+5u1EeD8xJ0GD
3uwcZhj34kHygihJNGYnnwtGjDuVOvT6RcYZeR2M2aR6f/X+PKrmCigRB3Zdj51Uzak1KGQB3jrj
0l/6KoNtXSSb4ecA02kzfXmxmUHFh5FpxWw7DdCQ0kn6B+2cgtS1yWqMlpXCfANxQO88vPeeyqW4
EpEkPLZROzzK+ffELdAxnduSQ59TORM3VxQvPpTDpcTAtA8fCB4EYiZ/9AMewDcGWwQlFTo316ja
wLnsyhH9dI7ujfnlRT/uHblR69nrsVa4L2jzOWn3Vp8JPru+jdcIwP8N8e/7VVQ4SIe7hNi9Y0zg
iDwiigyGG/qX4XdPLUj0/J4EB84vuVG5Mwm+GmBT0H6RKHSJiUPRiEQasYrm6ko+Ot4iWHera5zl
Mz2+g0gfp7VQDOVpdPvuo3WRSeK7dq4xgWwd9gsGQ6VgEaYG0AhcST3QNcAuqydczkdVVsE30ZAi
HdrEEiv95IkfUh4urTJP7EF+2JCacv1xMQIEH1EU9vLmyIp8maoIZ8SpbIivEJZO01zEyhme1WmL
/THf3TOw0l4W8f9DYJ8NlqJQv3TYhg+NDzET44mCMvUkO5QshbYeaV96z+HQCEnLcqRk7jGiCP2s
cwX8rZiOKSjeJ7PF9uHludSHn0v9uZf4qSEJ6KCMlBB7koX2isgGEXYso6HKxdfu2ry3TM90bBal
uGTcsdCWCOHIpEsOS3xEDbwnVJ/WmGmUJhF2IVxQI7FTWF1l6CTnaeUiF+n06Y6WEzIXdQyxR1dP
sZt8bNwLDLQewRw5tmdh+5dkUqrU5sf6DNYzO4HZ3bfi+Hm93JdUDvwxANw4efSwJuX76OReUEQF
c1VGcN4ZKhqYunbeBoHVTQBtOTVbd5fbQNeeOg9wtvelCCLizUNPAkudBAmxrOcip47MXJUYGK9a
gYNxebN42O+AChci1ya5gq+rTrsqDDOUG7+6JN6YSHmH4nD1dVdbcWwtnb8tUSp+0aDMTlERoCcK
MTMcSMQFMPLoZI1hk9sCycV1XgXJcRZzNDtDjQM/v3C17U2PtKVe+3YbvHrzXMZjOnT+r5U+6Qwq
zIwXqUe+xxEDdAISMNvdw469P+eI9NdT1JJPzbaaCfnRVDKPFb1UYoZaLPx3W8LY/xtVXz/QZC3J
Au69hpxsoBBycyFrAhzQEeu+fbguni2WUVzbzPAHuddco5WV0bPbS56kaB1YrqvvxiUSCkSKm7RF
c651pO6UGboo/bmEp0w5L7aOuKkbiXrWldYkY4/+ZESjCTDUW/Fwum/WBPPAacO0JOP5Hrgi7Xqz
8riFB5YgF6PPv7IZATaaaMb0dowrpgqOgxl8pL1MHZH3IpI1x+tR1ddW1KhX+FsjmlmO49jF6QXZ
x/OJX5ER57sFRj5HJBRnjLIm+kVdL2zQgJpDde4GKPXJXzb5OnT5doVb9zsKzz0VELYHpv6Diy7C
JsZJqA0fx24temCvhrOo8PdaYtpwZvS9BOKGQDlphenbhVpS/81hFM+jb68vCvIiiNXoebQiBNeF
1v0LjRVbAZvBD1hP9KICn2xIZ4VXT/vE4Rvq416BMDGDsqnPHVGwCCCTYTLiFBSbOJ7bXcr2H6mU
3pAfYheWm70eJN5o9W+OpNrXS5SyVWfwGw9aW2NwxMS2y7cGTP5TzuAerM4mE0qRHKzs58Ax48YX
VtpTk7q9wPmqwg+vpHEhEEgUTUhaQONeEtUowAvSsfEzigvSs0Uzo33NQCjEMhNE07g9sFIkdcmW
R6L+86H/47N0vVrlqjDqgsHiU1D3TGvDrtjqdBQKREKhOp5NDszHxEL8n5jJTK4X/dj+OUw6XtMU
1LAWDBdG3dwnNL8TBhVL4Dm06qBkQ6XflnaepYJBLAqvw2KHmm1c+P+CSlcgOeAO+A+mHvAN+JkO
+7hG/2m0s+KcGcNHwb1BvoQVbBlTBW6NSpG4HdSpSNg96pJz5AOCfcINTD8/64vx4MWkJG4tFK7U
N+1vfz5L52eXT2k4buibxLKQkcKW8QNBgsIlBgC2l1thQKfosWSQ8xM1kTP2r2RMKY2ldvzwVfZd
e60VG3riqDdV5eTrYKt53bFfe/xxnuU2p73fncULFoYEuMjmtsjcwTeriSoVOVBo/VIZuYHn/dPa
iTDmGz94+B38eUjJZPPOAHHWOrA4OHoS0NsrjaCmxO8U31tW7S0Kf9BKpvuTeDgtaaxeYUcilpjG
cW/LOAjWOhWhU28+zwVd3qT4bZR7LHKuw4dHIG7aUcb+7jyhnEgLGfI9VOwvSdhZXXYF+oZAUhIX
I+2oQlqgMvzHbUFRZx/A9W4Au/LbYjBaYU8P7k8MWbspgeX+c4eCzQd2iWowDcBB1uzvzR/KgaW5
ywAV/sbYDGb4JnRR8ADj/guPV3KART5gSS5EtzWOHZVQKbSSPLRxLfnT91qihW8z/LhtWMfKmo48
jMf53opuODpbBIE8LB+ORWxe7/wVI3ChpYZQZHyQFj6DJ3VK7CBxMmlf1f2BVD6lFEjpQYG921g2
g6qyAXUUUwKiknPrloSxmCWOcr+YWf37ixVjtsTg2itny35gi25ZO90kg1m5HTX2GZksZY0WnW9R
nOY5IykplsLno21wQ8nSRQW2QU/a7baobsAzp6G50OrxcVogmMdNPWws5Z3IoKhTVkCTTmoaXKpn
nZQ82o91iClYs56wpwbKP6cEJh4VPFqUJ3hLc0WNpkDI0JdZVTAvAvGSxqEc1s302evVIJjx7Q2v
VVFiAsyhaZQlTrErTiYfwnxIHHTpM/Ws+XVQBNQINIB7I+qiUG87YxNho0t5wZd/LtozeqljNo85
lQeBc1NcyMrnm7QZ9nD5biZulyaQjZPrq59lJ5tJbKDTTLMKorv9m8LURzqF3dsNOY60WOsspP8y
mxeEAXLXqsVNvjwonOI/fP705s/tmFWxh6nIl5Oog4DgsvXjYXX3O4qkSiYxZtOoxns5UiLZPL49
Dhy3J8pAWUN7SJEdK+alCpPqn7pb8eqfQb1rU4kHhGeRiTiGmyuB/CSGoG9BtJewJ4Eyk2pP2dIT
rdywWtWXbdHqqogYVLNhkERKko6bajuxie3aRMYcUbndUb3LYULl7DdZkfZTCLKr4DpFuKL1F/75
AC0GPsdffHXVu00fJ18uG6WfYGW4Jf4LeKo0s9wFnVHmH+geYoQ+CSOHs4I69qW41sPDB2UvBl3s
vS25UVKX6go9Z2oUUPNi4eoSA37NJaE7ZxmVSJevGE1jBDVAE99rGRS9u4S7OMAnl8bhY2sMxW6k
tPeR5T8SJhnyzd1oPZ2Ap6REUTcNBkAkD1CpURRCgItCBTEAX30jb/FHfF3Pt2vEjFl3feox/Bjq
2ERg8RyEx3HeSyMGAg0qRtU4zMdPy2iZndzsXXWjCt1hP6bXT0b2mV6KILyZEbhL2hlNIYPpDAAL
kekY0PWT2QSUcSAITiyUmCvH+hEf1jLxK+sH2fYDGPRCdya5pceURDR4/jth5zsldHc7NMKlPZPY
nBdwBlpDasEUPvi1gQxNSaUh8DQnYpoN1ppKG+W4t0ow8ggWiJgDBdZAz4Gsg5qiiOZE14Xt1A5Z
15g7OfQFnDeYl6HAkLn9YFm19xkjmzxo6VFRJxYssBmVUN5S6uFaRNs+XNolaL/geA5YvuwLagfY
O6UHPXzXe6MDLjbOQXuuKXwmDVq3E4+8eNd/S7kcYVFCu1nONzbJC24HTVUVE761VzbnWPJx5znv
Cy5QtWKQ3yYSCQl/CPUihN7vYUMt9mA00NUjUlrHempttyKlrOxxj6glWteySmLbH0dSDUmCXVU/
4vodYgVP6x0hhaSSd7Bxkt9F3T9uFlpySZ5f6LT6NPNXxfitrKI156gZ2ViMM9tSOLWzO7EXgoUc
z1bnAWTnkcS5iyf1b2a5IB0eznVni+L2URz2F7ChBuHVSB9/YnMtTLiUhQZfB0KEULij3TN6uI7O
T1scH1zwkOJVin41xYstIpLmR9yxhaSOR6EnNP33KL0hMBKurjNBBcADg1rkSGLnhbPwdnt4HnaG
GMevavvMjM4BXRGL0w5mJW75Jmw1WB4IFeq8JNHdZrIX2u6w0hxEohqB+BDE/zokglgMR9XUZhTJ
y2i4vkfcIutW+dcrF5LAdyUPuAPD1IXbthU1kZY7NCXoNbfRYbzBW2BbHTyCnj4hHxo4UOSZQKs1
rEP6RZaF7+HfZ6DTyopLcJ3kqKE2rb7P39UyWzdzIXNV02Wrwd7TBwyE8cZ31uwmCQtX49VrFccQ
mKVZaa9z8Mk+huxbqVbm5seIwbiEo7E6ktiZ0DA9y3yyVvqDvv5/KmT+d8uqhOAx8mL93TSVqDdd
eLaAc23khHzUULQgcWoRN8I5ktgyujhKd7Dk4M9OT4gf51M++Q89Gi99AAlsWxCplospttYHMMW9
xVjx0TOv/vnXQGpxY7SI5BKVf++KlPh2TwL0CaBmKVBqx1YuYxJ4pc4mK9nlhZ6Riq5iA8IFeouR
3b10Oi0wIHTVF6QZjEpm3dXIg6jOHVf7gykngIOUSyCydy8t6ZfdCasP+ut4j/GMwQPCrsYcibiV
zl8IgdbU8nL8QX+3iMKSMWcQjpM0mwqEG2ZEChIuRe/LtYq/ksXPVAja9bw9qlMexrL6+iZAg+y+
Hm+TBMZxkkQf999bkGrdthM8BMjc7WSi5EzURzEidGPU/VuRkyAOPBctwW4Ze06Xl2zeJ/Nsa8VP
On21R1c8tpEHJp5BJppIqILETlFQoL1HpAdKJvjEajaZ83P+Q1GdCKw9s7HwnKVhWLz/BhjXW8vh
7y8JxWuFnNMLhDiGZGQGO5ses/M0kXUHSJ4mfH78el9X4UtJ04oX3qnEMKC7tjIVVcrs4T8jvSLH
U4oECq89UEZcAeImgQ2yvg7T3VqKDFajLK9Dy8WvsSKn+eszKTB5l3cgo2Pae385uFTMdbOk61r0
tyPz2CnYPRXVWLpdonEgYCImAm3LvLM0CegFN8Eyrt/afZSTqz3c3fMRdcSjSL8kRy8VvsYLH15G
0g7YRpTWHm6wH33uiSDpZ23jIGn8Si4rtn9npkHjwmfthXHzJQnkagpC1ibzbmOA8m1NMKGS++8n
y1VsXqGThKuTDRCVqBSQg+4Bkyh7MkqTn8gesB214gg+dfivpyCcHzdkPumNOmQEBrttsR8m65Ez
0lRmstbQL/q3x3TMg7ggniGFu+nxL9+3S0YoFgZ56110M9ZBQkt3MgcQBi3QuNkvxG7vBLC8EU70
FCfXnpMwpJthv5IRDjBVR6nS8fLlmC9LGc058+/wAlB8Qhe8rG0NyNcm3XB4eJBIjHMu9lXK7byz
38qqWoGXSEvQK4xaTdzMFc4G/4oGkWnRBtkW8Qfi2JWrJLKz7I3eKPxRRM/CF7BWe62Y5hmJEPv1
Lr0np4tfm4fse6ySuYkiRGa/IumuGQ3ssH2SvDh6rtIYlhq5Zt9w9YHJ3wmaAG5D1pYYc3dnT8LU
GoB73LBb5qGfDirAbc9ozRVJ8BwZCOZ67vMM6OLR8tLMra/9Hf32LySHQqDpZAsWGyoFrA1lRy51
OdSwXsTMy1+ym0S0k+d5L65u2275ZUySdlbTv0o+p55cpb3ujbgh5x492jmajT8vVvTsVyRZmftC
glgAiAMFY+VuDkWNA05Chm+7xUebwrihGOVqyQTGB4z17IQFVeM7RPopxY+dXs0D2b+/2afkCRhq
/hNTxpwwPqPW/6DLbvofcJGYZNb1eZzPzk+DOO5sZclyTQldPmYU4hzYwqS+fyheKxU6OzNFouQW
1bQWJSdOHwmDBTOXbTXljq0xyMAgcZKDvHy0RMpWO4FpSl0i2G3Zs2JK38gxwS+zRLKvqjAZIOvu
XdweH/+ibRIckIFfllcLZE7JHWE7jdv+wkU5cSijTRjlzcgKotZS9zaEZGdVK00f4YDbStCNjlIx
jGTUtfwfSNX7c4yWHxY+3fJIJoGopkf5lZQN/pHerkNAd/iGWgWWEtYyzCLqnK++lPD9V5RzcwkC
Q8bg1A0GxtpRVpd8ggP3cSQTlzcmlwjzcKI8N11YrowiFEaJFZ98AoPtpQRfYPwj0rGIc0Le6zM2
KBGQE0a5bm9fGe7k80mPXD8x0mZ+4AtVnsljRimReGj+Bk8a8Dc6TJBC1PbM7n115Nigf1Cp8ho3
eDlJOeMt+OnLhOX3GjM1Wgl+XNR7rP1U45vWZ1cVGq3nw2J4kEeuJ2RZZOR/DoG54k6TZvWTjBC3
iLk9NbSpDPbKKmLst7KKVfPvQsldUUd1IH8NP64RgADs51bvlR7lZWDrtANAWjbkxCFGIk2qH2ED
veQYJ96B6lPFMuchc2c2Uli/KEkMFbWrGq0XAtJZ2xYPsoHjwSUslE3A2r0L/e+D5Oc8LqbcFnAc
Wkm+FCAQzxwbmnxMFeuT0WYGBO2GfmQO4kb/s0cVSuQSMuhn5YjpsqMUsT5U3zCCrdG9yTpsyDQT
MBd2oazH0AfFH4nsjf0m1WILlCHKDR8jzcxJFigrusEkHDAP6Xd6aeZfaRrj1JnD1rC1L53tRSUc
983MrIjOe9Lbqc35XSisEcFWhy/qPX/yeN0nL6bZtYhEVsWYfGqL8y6VSQQTTEiT7/0GauFO/XbJ
l3289TxAWbT/2CYGI7ARxxtyvQrIr6lA/PytgRk+m7HcYE8vclNTHF6KITFaYM+siaEHVuR4rj3S
AE3TVBtK4J4ZO8Z9261+7nHfzaXwbv2zHNL8OUWXbOTu9xKwxmOhW6wjj9ziJBrnAFpOgpHxYHqG
3k3/WKlpJHYyKM2x31qRVdLXHlA23RC8Vq25bni2vMNWNhun0rNrKUB+kuUOSSkZ+QGY+CF/z9lh
TuZ9Hw5TdEURa8ZVlS1Z6eAR7ffvakhCLFKkLJuXVD//39gGPRyTfau9vWFXQDNw57Q1aCLYIktW
CAjJ+xMSm/AUdNcq3yljd/e5EdA8bOt1p5gkGKnTQIU0gL5MAPgOpi7npgEpbYbaEyuoMuY1oPYg
6oXvHKMChJxmj+s1u60usfEQpBEIKLXp+3HRpyXGM3NtttLBNuWxjbya1irnw3N/DbXk9nbmW4KP
q4ZXB/BSJc/C+UsAnsG0nlkW58b9BXx/YZxJ6i5/elDOqlbSO1AABefEX5N+pK4VId241Snm4asY
74M5IsFVEEzlgUW/VNbJjrEaqQU3PzBlpnipsS9JDd5xBcl9vYA5Wg+zCTROGUP7qwTx4cLS7WnG
8gVr2HnqUC/Hr5roUugWNyFbpD8mTt3ZckTN+ly14+ZMOUWtPnHAGI4x9i00bAAASf48EpBB/tuB
OlWDsa57aNUZCIoHDGBapiS5wZ9F0D57TtZtMpjos9vxiYadEsXoja+z5e9d178K7Chw/0jQAxxT
ATVHK4USmJ8vw58ZMsI/ZWOZJOWcR/Io/h77YHC8/8RungnfE/DE9KPRL+vmIk75omHFpEGqdeju
OZjRHRuW8p9nSNa4AzD7QKf04En2SvmSGumpdUBD8dSQiK/Meu8Sz/9KCJlqE3XxhrnXBkNBWgw+
Ithj2xxVv7I5astKSxuNOM7QIEb71NAMY5DuvICtgq5EMAptuE/gSpVLqAcmH0Qx/rOpxOKinCoP
3T70NbkfORoXS+nVTlJSMzuI+e0YauuUPyw6xKRd0+cWk33i8h9AWKtFbCwHti4w9VVaQDZFWUZh
rIdRwxwHnzpaxLXtrLr9aHw9hklS1H/773IFuPo6GPLEs0JMTn35qoFCtGLSm69tqhcWKrIbUoKH
PvUh9cA11+qJpYOdyrhupXuMcGhE8qwzB7OpNsjMDO33ewAVnTbrYC9G4qDdTsz2QD4cbHVo4WKi
lYitObkRfaMrIf1IfXyut8P1pK4jsKvFv73jlWgy+XDLyGRU8sLLrcEOIgQFOPnWX5eYuAi+3+B6
Qy/KSDs75YUaBRfpZ81bw2N9Pp1NurTAhFE3N9xzlPXWr+e6L5vefijx77pqwuJ5KAbBEEDXa90Q
4uMwL1AL6HXGRQ1mDjG7Dg4BJ1DllTdasOQgP09G8rfP6S7ttRd9BkjiJUSlhnz513h6c1kRVrl8
33N4+cLgCIVWKB4NW9W8odQOXF+2+HLWYQ/FG/vJo3RJY8yXw6YOPZeu+H+GS1v6zE0awzCmgqD7
AhDGZUJMGD2jHIGWDzeCtEj/XQ1c68JkTOiBl2K50y3HNDjMWGP7yyCM7ZyzmutaqN3wv4bDbNK5
7FD5XcffPND1KLOHuiDZ5nxQw9RIPltrCVSdTB7K2RYaGtEOYaTHIsmCyo4sW2iN3tPJoJZ14Rxf
2BcUEgqiZCNQbQ5JJuRqmjf2+6JW5ca2/3vB60MnEGjDiKf/VpiAOpAItSZktAU9rglqZDcrZc2/
awJRh93G7fV7WUHqZg2IpuXae5bD8q8uxSgUa7Ba9FqHGdmKwFgxQ5PsLNje1h8pcBgYWn7aQQ41
XKQpGmgEeasd76HfQ+C5pSeEr++BrfScPlu/kFrg4vBbIUpW85WtXIX6KOCGYgRoUGIJrwEUcyzM
mqzOR8+LaR9h3a8oyIwUqLGsVLijb6jQTZHuwfJ7cHh/GTVmhGewWICGkhCXg7nmBc8LQJ46Bg+D
eqgVCsYyHU6cMCYxfCDQoUX6rlIAE/3V0/Yx2ImjzNoW99QAtgwf2UjRgBsT4VBvmLjvwcKE0Sn7
k6xwMe+HjXh2pFxsJKaqawvRb/jtCSLVOZjEmhSSSeXSpGDZip5MfA0Dv8ExOO0GOoA7tH/Qghr5
2bue7llpK8fF0LvmRB2r2Nc494I4GgUGf2Il/yVlViaI/IYJ1J2x3meKuMPMy5FL131r+xkK4eEp
BbTfeBaFLw4v0Cu/6n9p0A/9Ss4Ad0bhdwzyUcyutTKBFDkXqqv4//VxRnpR1AqK9sAdj5Won36I
xn/0xy4DS8Hsw7yc0z3do8/ZYwFH2sKT4lj3VfnfxRRBNsf1XksnBwhy/zksI8IatHfIn4UpxD02
pKqXQ2rxHgF00SpXGe+C1fkd9pffi0ON8q0ea/NtGq6OEfz7ezH4TCLdT+Xg8aFau5ahkYjGor0a
CNP+V7sCvQKHeMrEwdtcAN5kP8hCkFApPQZi1Glab0LkbNcyMZvwvu+MgDA1L96CMCdz8P16SVGT
+UzkuyN/yTttg7yQRjaSzLyU35R1ehAJkv2PVOHugPuk3jW3ed3Gh16jb9U2bkKkJ/R36f2sl5Wu
A45XqnszrMWp101Ls2fwF2iMOszG/6MtRWX8UoJdWCwAg7cTFYNxYR3KsaUQKDl7kyEHfyRtqPH4
zizKOKq5IUGNJTsOjdjKoahSFfz19C+7nuYMRFViKv/6EAZL6YcCM9zWwuOilX3v1psabiyN6Kyb
B85CJgWKXkzPqEeLbbnmaYvg0e/1K8l6gSMMZtd5yzIl2fjbdgJcfJp4LRA6bMzdQKqWxtfWEOgn
Lv+J/TuSWOOMzuGP1SdlGwYgc8MdS8OO/O+AhWb0wu6r4n0BXGjKjuqYX0xNGPcvxhbeF+hylltv
wVHUILYXqkNGUQ8RIbKWutn53CY6gaEvhUr0nUjzPk057zuB0aSmZzr3c5Sef0shsLPZ1/9h48Ux
ay1wipAH47wjUuU5s9kjeDU5DXoU9u4RSfdaUxc/xLA0pspMp8XG5/lq8tpwVUthezY4LP9CCl4Y
zQ2HRJko1GtemdF6q/I88wCHCoz1Iiu7bhC23VU3jUOoPs3N5ZAaTcY4cTBWBoWt4lSwi2IBArl/
aTBCRf06rElwgR2TR8S9XbMgoS6yike9AMZQUmaBcoT7gHw7+K+RtCRsd6NMn5A7OiDv3ufiRP0a
CnX3WNZ4NpBYT5Vr2x1uM2OQzJDlfGQIqdCexnkaYxnOnT4BQfW4CoeVBcSRKWSZ7kBhjv2e9QR8
KsxEGV+IRwcw45n5mxlA0p6vguy4Z2gYLs0/VFHnYwMpxWaIoWB2V1lNcxFqps0awE64tZNOImk0
RwQ9M8Dpp235lbkxdX1aeue8gA1w9dH5+5OQZ631dY5wRgC3ovt1TIRtKnN2aZlrs6ASxK1062eh
8SDfVPI8LB6cTgT1x1ZHjHm/iIyylK2L6RTip6gSXSnK/QJ0SaLFxzf1K5e+foFZSJkpGtkSg/Gi
COwEuq8RYX2r/Gj1rh5la9YwgUUlfn5XgM7kycfuO4EUnIaqYJjTKaJYVEsbAGUBTcM2lMyjMUfg
9ta12/U970mZkHiTM6cqcPko6ZMljumTLgtxaNdmtQVHzmKWYYchdI5mnUMdpZ0tgByOHetxGCSp
piuDvIz0LyFtN40gtBSqCt31sKo76VPa77Tf6RSkL1tANii4cy0dMsVk1E9FL/OwXkigSZazLDWU
PFhCd++18ZPQNeUIbX+uJg33XfP/cWhM2l1WXosZhcKGEnYCDCqo7Zra3gw9jg1BkZA9S+AhhnXR
X0h/tU3c7yuQXckGsEttBKXjJKSH4E/B5RjIG6S4fGjkibC5APGV8jt1JK6V4K5Ehg2pTfnfYMZG
IRktwZdiMJzIhDcadZelHz5jo8jZjsIBdDfcQwUJvjIn010Ii87v5g3AN3WU9xYKIJ03txVK3vhg
tmWPvEUxrR8pptlWaIJ2Xga4pviNlEJtvFELZBRePi08+QumsKzlq40ORg4Nf1GykZbD1AINlhdX
LJMtnZxsIz8DdKtj9f2M02mM3+9S0JaecTLTKNkv2mH/QQXwS8HCJsOtiVKwRBFnIsbJpwn2AKLc
YbvaNqMzwD7SMGAv6gnPFx1fPEN38TnbGa/8oer2uMltBWsWnyteT1DKyVNw0McheBtXEp2jMJIt
tPws0vDeXZzuniayKFKCkE7CERY4nHFl8JfuNSmRHUeAGw4H40IHeDE6QcqR1YQ8gOL2aPcn3CWG
a6kd9N4TYgFsE6t4Q17C6sQ75rwC4WYUzNcMTw31wfVsrxAXMpxUKJ6ehKobnDl0W+m10qBMHJfT
di4m8F8pULOyQlSatRyc3ud+14bWvE94sCrQsShcoKNB0xQNpJSsjekf5J0jbKPRXw+6QuWkti/w
x7aAZuTav2PrwVZAqJwnffYHzdAbtbLLYg26goxQ2ysYgmJph/mfGN1pguV4i2BhFhBAPsiG8t6Z
sNZDQWphKR9FvufIVrHAMl20AJwM/ycD+7D2AHckFNaLrOQyfSsLo3d54UT1Ca4ronres0Yr9/OP
RQ7AOgrVb11voioc5lG2PbQ4Oh3gZaXBMRIFGwuxyqRPMwLhZUAxG1M0k5oIWQtMBL6vJgBMQbsT
v/KXkKe5ErRUYkG43yXPZj2PzSlipbWosQqmaoXySQVTviYcvo8Tn7KN7pVODxprOlO6zGFhFx+3
2rlEiWth59ENkd72tKzdznAYZOptN0SpVJsXPq9WoYBfKTZsAvZEZ2QUgDDRyBhOzNZmShYLH09y
SmYkr565REuCTjj031GY7ru4Do7mV121DD9YThSjMfLylwlC4M8ajrVnD0uF6oFzWJzrfji2pXII
ypNkFG++p3aqrxOzHVK59E9mnUBnRJnG/og6tQjjmKPa7Isa8JAqcEqro0nQUHN+TzvTj40wff49
U8WIgM0I5Ak9gnkDf5AxhgHD9oYmX//ZLfNJc67Oa6WylZLLZmD1q0lFUYMybT8WejhzMRXoPxyW
n4juNzfFpC0QAvM3cDQWBqQksKpYKvIbeAF2H/5zTWkUK5+880n4zcsHbqnHtX1Bj6TYHb5wXHj8
DbFGwT21IRb6ZypE9UE9EYc1gNmg4oI9zByTHN9R0P5yAyYYLKN0i/3Rvq8r1FNd/obJkFerdM5T
O0WoSXlxcYdHsvC85apgjh5m21NqCYqJqRcdLbMYxDS78DF/9SIPeWopFB90oTKP8q7w63kBewPH
6v02F/wbLCW07El4ixo0rIHsc5SDLA9zIoMZHL4eZBosOmOHXW/X9a/tMnfR2/r6UnUJhepGo9ps
i4YlBxVYx55m/ohS2gpUvXwXfAVRrx059/ttUkVGXTmEe6cvFvyLsH2VrVo3D4iXj+wqfzDv6AUD
OVlQz54CFfDXNmxjs2KtbNBTRb60mullXw36N5yQM7ZSOJLGLc+FD1d/5olLzIbsvlLcY5t2VbIG
q8CMDV7zGTCBZA4lTlj4zjbNfHH64Tcb5mhjhExHlMjhqpFUn4ISbsS4wi78joqj0s0uNp7bxL0/
96rZZpFtxGjj3Tk1fTJ5A9sxHS3aa0AjFNWKwh4ors6g0Lqqm+xjq/4na0XKD1OMBjrsvgmGSomw
zbQArAXootspBxF1hGuURJqpErp2WoOkDNHv/jUuiEAkILoR9AlwVrx5AqlJY+/loLxim9qMxG7A
6DI4oQN4SCBeJJ2MDOQwwE0jGE/B8Cmw+gJ6raRKjDM4kHixAUJucr3TroPLcnLiCeynUiB+97Xi
aM2nNPEubxxzHvGXycJBkm8ecwgMUk/D0JGtm70oGKdDJCDFfU0GvHEmAkb8NZwP9KwsUdKy/Cv5
hFeu2ybpcP7SXuK6w8B7Xg5VPhOjuL7y8+1c1WRnLaskQXQJP3akSVjBbmPt8JHenDn0iKzcBzZJ
zQJAi+uTSZSr8oQINU0Fzd4gjqhCM6brQ2FB8YaM9GRnyCJQToKeuH177QYt/4B+9sjhHdxH1p2i
ImA4fkDUBsG7xcs39FnlTJZRo8sEYa9iz9d+WBmheI+NBEUQBKPjD+FhJJSIuUMHOHaZ0fyba5L0
xdE2Qn2KeaDl8r9z9r2cAHaYUyB6mYrSerKRpLbMg3Cgk0Bh9l7ShbA5AHHLJNSmh+7KFzA48h3E
NYwSYWTUZkizFMhIpmgu/8FKMLfqfNAaBaIR5TTB5LSPBaWABR0qAMtnqfumpUrrra/W11UwlkDv
DbaRvx71SsklierZId7WovbxZ51USz0CALWM5jB5AEJDdKC5wLUop97rRkWiM4nNp3j/P0jxBjH9
KXLl4UUkhXSE1VdZLPj1XR6fMP/RNurEKHTJFsb7rtyM9qBvejWgLAoscKj8xOhGi5K4sQ4gumQW
reAyPnPL2xHYvuIakvvKJQ0Uyo/YK2y1Qxjp24OZ4BzZU+isOctxMbCFUzXn5Fdb6pMAN4nRoHyl
4VpP8b1A0rOlseRALNl53OZryEfw7bfGYebOvg5qp1//VGv0ucDzE4X1SHOL5NLshdilEZyEZDJh
7A2UjHHvfgPEgvwkzJCxtKA3R3UNzGOxrusalxXWupxdZbHqKvuoe7AMQaJpNrPOBHDx3i8d1sZi
yDHDDJPcwVe+N9a/8pSvhPycLHpuSio3qcaDdhCVh4GmhLV7W6HA5RmxOMAENpdfIjjQ71P9ffOD
xCoKJ7vffMc4waE0DqlpSmgsqnkDjyDTjZWbbAS8Q/yLzHtAi3dMhuZx+CuHSG+yRA8J/nGAeoqH
Ndyv+iqWT6vIFZX93HT6zNYo3OtLzVIJhLAvQ0tAdxITzerXlegyYhEKmVwy8g5MRsFIV1D9ZpUS
i4UlQehcMEfM4FxjjLXrBDzrNXv1MVzgNPBQewE+kwXZu1mfJQ0E01pvsvCSO+BGQI5xd0XXEtjO
cXmUqBeVhsDHcgGvPQnSA5pDNkIL53UEvfEJ/zsQ55ahCi77G73kUtBiGwEQeYPnzAjiT6AY17Zs
sjZ3L2gTS5Dnu4W3HVj+C2yqr/YLdJUZyS7HMiVNR6R9X3I93amCZqJA9KQbbU65zFWlrktuWmAu
pjLnXMzj0mlez0sycEZYrQQFkBLaNeUr8LwfuAvgyXh/yYIcsujEnepfL63IM1Ei2ssgqJ9p/FMO
lBiQPfvofa8PpvQOgG9eC0b/aP1znAwtwjR/CRwlewqwWzENsvy0MzZTh/OEk7XQDqGK5Mj3eFNF
F3LCUV5ocvaoIdcnlZgYsK7pGymFrmayeBWJReIRyYD5HmMdaNzPhSsGpJwxf3fpNvd5APyKL6rq
2HY2a+wmwH6BnDbL6jIhJij/JIL3Ta1+rTfONeQGVWJ+W9bpXaW2xk5+jnYYC/A25OO/nL49Zgdt
g59Qcs6tJj+4iLCfYEKrKxA1LfSRr73RvEfZs+LaJ1l6F3Jq9jqtThzrCS7X4UHEdHh8SzHPRk2m
1nIuemLjrk6ft4AjLZZEWcGO+aibA4umVFoB/ZlP3qp2k9iP+Dw5GKS/k3sTfMvFxpS4ESKHuJPg
7WY6of2FBR5Fz5p+2im2RseW+mw4aCHM4HH07MJKbqtnM9EXMEZgwA/3obyDfcY9zCfR8u83FlIk
ySfFRUrkm6+77Y3HQefxcg6arePY3cTqMumbz8ucIC9/Hg99XuPZzXz/MeIgmHr31ez+j4pLcBgj
t81xNZ9wLfUEUN1ia/Az1kuLhGTPIrlLY6vFPCIn69Rok7oTBKjjMKNNt0fcVa4+S2MX0XE+0VDu
+zdRX7Cve2UeXm9/5ygzPcgL7gGfiOgGhvIrEQvYOHFuxuFNvrVNEGNDfVjhBXBbAHwitKXFwpIp
WhyBz/H1owGe1ScNbroD4XBt5XHUeWZk0G6bEuacYYM3sADYln9UI6yh3ddulduRft9hdMa/73cA
vGbwYH3Psg7hprb7Ngd4A1hXIcH1QiyA3lbDlnU4z8/OKnahJug/xbkpP2mg5LrR4W/aJBaH0Lx9
aY/OcOsZF3uUUnx3X0IUGmVKPl0pT05AKMZ3jvzDAdWTeBfL10pvYandQz2XvAEu1X3LEU6Zuqa6
GiTD7xszwZFbvwoSbh3Aq+QfHzyjQqxBFJIuk6u5JYUxh9VIn1Z0hWnWqjv1BSSO+eVVILivWXFZ
/ApojcCKMYT140fO750Mgu+YRe5tnGnLFhUagxY8IuWuNSEn1wywjafKwQySxxB1dz0oR/Pokx12
aSJFrQ+HXpcceCzN22SHjB7e5k3vrGBkv974wZ7jUYW+x4E+0axiAvtVvum6vVqcig7L5S8OkM+r
rBCn3hJV+a4PDREGxWg2o2Ay8dqy8OQuT8U68j6MHefRvraF5Ax+Z8k7oIg2PMYPI/xvEKLMYWqY
yBpgK0hgNqErd+ZNjjEUFqBYCDzR0HNwrKZTq26iPitUmcmTOBO0DeQFY/w8DyB4NzM/+AXUjHm9
w51anIGo8bmU21lnsL5ZXwJtAij3K1J/Du4Zn6f1vKySlg1KeCRJgEI/N9NtpZMvnNWqu56gXpIh
wTpo3zjiSDWpYxkNkFcSI2BU1awf+YfnqhFE6NtsOCf9sn8gw+mN4uMxaalHvP30XXOs+X439UwW
n9rNdOwFWC56a3F6oqSV61BADhQYssLmBLyyxA4bwKPl/l3p7nckb7RG6kvSyGjQBsgpM8UZ1nRk
2d8FszXyJsO3jieVqcPPJHMJPMfMi3uc530a7p24KrgHi2vngn19aUuM9wrrV/UHN4t0c/UybImu
1E4hAYznRZJ8iZhMV1ro8qU0h41SrJ19JAzAtUbxcOOyScgYLRLb/BIr9E8r+muGIfI1ppk+9y6x
psRkl9wWhBkPRMcpVXzVOkUKFfvh6I/zJx0EUMD8mItnDYFAIGUKbQSO4+azwtfIHJ5SK0uNE9YI
cTw0drjlPnrdtmAQoITB9tUJfiAWjGnicnklOs5rkqntOxAFskZ6v2nSxNQCa4kD5fPg3sJC71IG
Wea+tB2IYmIMeo4Otm1hDkMGpjhSCyZUekeeWRXCAwHOLD9T6Y64adFdqGBl//1NDnoQPFK1roc7
DMfEaTh66/vJGhEzO2QavCTq8MkwjMAFyox0vq2He/Zr9rj+HhVkYM4mIipjp1g5QHknhqOT6+UL
+t0mLdkEXYMAMPigUGDLaWaKvEybNlRLBR74246acqGjMWY+iDrlr5rWDmhi7/SyUvRZFCtljISl
8RMcHvXEPfCPHX76jqaQ7R6zbVtCZXfYM1D6+5n3OBII4Jw91aQKac1lhlXimjl7KDuBbpOAnXzL
x0zD+GJ349TG4hELa3dyGowXbct5WgBq2uQ2V/u8sECWxYYiiyjd1GDhCgj8JanmAirr3TA6+ceZ
J+m3PaW73OjOOvBw6x3/emt8YMw5pnsCisIYaD/J/wVPqgnWwhIN6QKRCah/q+b9gLZZgmxurRX+
Vy1526GWinM8cFvqaqTs8pJKOB+v04XNR+9817EhFCkL0dUfqeFZs3oubxGM8/tKGkSt4xmMaRuy
h/+cMkLX0tVL8z4M5LyPKraUuRZy/msI9LMgdAFdAahD1sE/0GbsDEUObGbaolRCr3OPHtub7fbk
IZmUPVwlwAJRG0Hv5Y1KOkw4VhEMXYoB7e2R9rtQldcJJYzn4S3NWTJ+3CfXQ1XUvsO7LcmGTc93
7sjpEF04MCxhy4rFS4Z4CGlozzLZlBALZ2jAojd0p4PHZnZio3ONyhPXDJuSPnalWyN4bQf/Mnio
wX9KQzenDgj24xIy85/yCRzDztQ+54rmOk3D8MowVfJ7UDpA0/3uBwR+ySnQ+HAHQVzEbFe1Hhcl
MqC+HkqbgLBH1cDlEWPlFqamULblHdHSFrgLoYijCIpzMgF/8r4xEPYy4Pv4wnuuDe1YIbtXWE6l
gzmCFc8W+JeVgYsbn89hdL6hWdR6HtLsbRiyUIvkYvlJKFkSLMuaSorCTIRMCB7VfKciQudY9OT3
coES100BoM9Dmru4ZJqFslqogIrhChHF5dTrpWaiYy3RvedWsKaH67hEqu02h5DAzsXUux9TM/Lk
ChyM0ZR3y1FGMpf8O8H+FYT5J8ohkZ5X8GOCYm5Qj4TjXZzMpD5wPDjvv6UlJcjxqAhm+iS6Wv3M
18pHWc7H9Z7Z+OUrfQOOsBjDUnyZ0M46GRiacW9PBv+MusAAsQy+2kxY+xVcMbwgPeE92dj3CqnD
sENL2nZh+vXyOQpCIqOU44d4NxnyVfo2ywVrvayELRb99mgMdcutkDlzi7+iZJMfKt3qB5sGlUzH
vXHfTuX29lirgS9cUMGPjpEWGAUgy15CZoAoX7Wc5tI+kwsxRLW1b2zjKrL20EXxSN8yKOVGsEPV
AUhN9EjuE4rhIwyoRjfjTwE1n1HwZuFihmGTmi0Z8OU1FfWay4nL/A9hQ3zn0xxeHP6TSeiycWxC
O5J+X1vzV050wtfW3bsHPcVdnBslVQ3z3Dq9pXFWTxvTs0hS4KEBjnrh8t/fHwkek77AYRan2qQ0
Ktn8SJYGSC8RXKZP7JAlGh1q+dN6brTGSH/PjFS0ItWFbWCr2kGOfuf96y69TvnDsNJsW0Z70Y+P
bgaG7ys1MHK+khyMBDxba7+Vm1b4PIyEBiWeodXmrp40AdOvqJzx/QNVJ4nPbRJ6YsqF3pQO1Yk1
fVIvZF0UcQkcbKTUyESvatrWCJ9aLaW56LRhrBRmqPGl/3hxufZoXp6IRnzK29lEeQ/Zlw0zLnvH
diNz5hFFajrlaIs0YuoW3NokfyleQKIhRriNJREgQK+TyZanfSxFm3w/cquKUJ9T/v4/orunUxwl
hHe9IRHTqU9IicrF0zlYbEYlBolUKCmIVIW7PTRvNhf6Wieut1yy/aJ3qFRVRjs8puPvimGsU1ju
Zqu5K7ahUDl1BEAg244uR4p0GATKqfYC4vm+UVAC9DGuyheFPxMOOpu1oHgRpVivGWZAs/MIJV4A
WngYGqOcoBhm58qQaDb7Ddr3Q/m00HR4M6gdoRd/FlBcHHk3JCukO9jd0I1suadKGhbkdlI7nsA6
TsbrDmWimuXw35kZQ+p4rkn4ORFHQKVTNRLh0U5s9uWCk6z7tFL/aX1aqdbG3KjFq+FDjvCWl/ar
YlrFfElGJd0wis5TsH6iEowxHfLKryfp+IhiYVA9bN929OBt6je7/jSiyLvqJpB8Vg4iZlVK+rAE
nCW5Xi/e4PBOzXFrsH5hV5rlb3LesQUVFA92mN9GJt+mlXLz4PACgnW2bWPXItulpm5wjp7vRhgV
mqaTXWZWHZuaZGhxMsi3nDkDxFOR3yqnuNrjueCgloBhh4O8jFIwF2OXjckXKoVXpxMwni5G3I3k
GsLpp7qa5GhL2xeXyuc1kI1I0HPWRF3fxW2GJGuse8YlvO1D6D2xWs47UF2B7nVOy4twKRO5dFoM
TU2Juvv6RlAy5izA8bi7Ow3Kjy2s0bALS6hZtcmfhRRCOVgFy2Ms8Vtl1Kq67BGJKmgxg2715KN2
ZsnlHSCD9uMsQixQTHOJ3DBaDVtu3vEnNVzAAsByaSIB+8YDAF0UuDT9k0EQEI2mmSTip8SIRFLj
WDOvuqbINh3H6ztPbu5R6ISh6Z/6QO00cxpM7kEdmH1ja9Woe55XS56vdKqvS0rvjykKZXNwrzH7
cN7PTJy3LJy5RvLo0RConEerYKeCsewDs2lQQRH0ZX5p6S8v9zOWL2a4qvFEsARXgGbFhvXamCNF
0SEJeHDIVoOpK0bKbbQlRCH2hrvY63le3EaZAIYswW/sD2MI4HaPgJqPQYGx60ZpzjTWAo1GzGCl
Z+dp4cwrZaKH5diZzatygxkvWZggRpU4W+yVq+rUhS0oOl6ZSNrS60PK3cBTeB++mFTbjiBWAMTl
b3oQ1efdQfUy5SqO6chhDnVJ+VQIWj2OfTRYoCShCTG4nnkbPTbZnPa7/Ayp28gQbTZsWYoIGSgt
ALbKqlgTXJw9ClkDTWbaNwAXMac12shYXwsbOsRoipInGjAsU0O+pvYoaH3VOIQDt52pPEM10YAe
hzbe8sluogr+K4PA/4VVLo8kpZGij6SkSirKOaFxgvNVXZVe/Un78BT1L7gPgO8bllGc5FLcz4E1
jTt98R5Ti4Q+yNHh98aj+w92zXfgxLj41BYh3GhtGLGh8Ii713hDrEAjuve+0lzNj+IxuqaOSkKB
8fZ5XEjG+nqIh0jolOQ4/Nl2qLz9eHf7paBpH7+d2LqpD4kH4wkRVdJsVJ4FxR8ulQXeVfojvr33
a4OcAlJRx2+7kqXDf/OJqBOClCFe8Ll6QjP/wYFiWsrO7I+ykQGfHpdYZmhFQ9x/1G8e4Euy7Ybx
bdM5BOC9OJV5yOJmhWf/K0NJuHPiZDV/MTcSIqSKvNOU0N1T+bvknVB6oas48qahXtH1+LFT+iX5
vKEBd4sWe6bBWN9lTFuQXNY60b99aX6YU4iN58TMVnesBK/WDsiTPSgwPMs9pWq6aw6VdnrEJfzb
D+GNY4YbzngaPQS3eB/2qO4cxzsR615Zcv1Q7bE5EisOZdUlbR0O3+T6iok8z6kp3EEELP9bLphj
a3yfGnADLyDC0MZXJKvGcnXH/dPiZixH+W29DNuNp4KQm0yW9xD0dD4ZYGWOTF8b9t2dWoz9UTJy
x4TX6H++SXtxdLd6KhUqfDH2RvB2HIWMExvYabLW3JOICTsnr+FrwsJfs6VxyChMzua+Hk/k6Sad
LUwVHGkesfS1S9MPUT86tHBjncTn2KZTG2ZkjZULwy0knXD5ndVpAP4sm+1zqIRJ5dwEpLmzE2Y1
4l0qrC8aGTr9qjSMP9Q+uBY8Ow6pDdyUic+Qqixe5zJ5gr9A3oHF8ZUf+Ze7UykigjlwBj9aj+Pw
RlMw0i37UXKPs6CDjZUZayQyOy0j3wP39wT5I87MtEvIGUvhDzpir+VoQJ0wqW2JwSq+maQ1Ns+4
27NyyULMK6Mb3plVMdPQx6iK8+FObqBg/JHePqRtQsDe1+JkdelZ+fwbTeiZcUXdQHzNEDYSnTW8
71X1FfjccDnghPrEkeeS+NzA5dq3jvVLAnGZqauYZuhUNejLxsbEeXTCyFazi76Jh/je0tWlK6z7
FuiPIBIvG1qTT4qbg2bLOqzXgoMg7c5xdpFW4fNiPNtlB1YliPCl9yY19yeEFaQDy7FXXQgpoMTt
MJ/qWLrapJ8R1R/8h+5Yn0Lk/IvV5aQy3vfiWmgYS2K5sSZ1k5QTPZgiICFMa6EeYO00w1gufS3A
L70kpFaLUTDgeXuy0D2Znvdn89S6Wm9QoDxJX04gUz9kSdfiMlihgGhtGPkIU9rKYtSZPANF3/sY
Lr4RWDDXeTyrPklMcNxYdjjNvqFL/1Vu4/GdVTMDK48kD4VG5PD4GOgBgxMNoQBborgPM1DlkA81
YEaDl72i4IUuC6FzsoPO59/wZdq2TJeQ/9Fbuw0iUhLODJcoxwxB5P7QtBziwqFByEFeV3T9uqZR
BeE3a2g7n51FYQeXYC2JG4cX+07kaqXrXOtwwaQldrodLcU2vVu/FJK8Rj2pSk5sXFq3Ye847phv
EAymdvToebYKWAnNzLQBV7n8PG7jIy5SKiqhDu7NqX44YFqqn5Bmzc2fCzciw+7V6bOjcPxNv9DT
F7HyF+/8fPo06zAEAKxT7uzu26e/JpWZn0KN+Nm6Y6K5rcYeCV4oZuBaC1lHy+Cxv26J+dO6jyff
P9HAoM3XHZyMQWDTIijP2e3YN2NJNpInzcRJtXrqintNrpiWYPC0gIBCKNBKmkc8M3MQ2TlwLr6T
9P2Wa3xqdbYSy7KQWcQQsECdPIBX2SdbrDOLs5NxyWLkyfhK2d8V3spgdRpQC1Oefw+GUOknP9nj
n72UCElCeAzB0XcXi4gku7FYIu351Degvt31pavTa7Qe7z5RlsKXT1QO1M7QZ/8RiAF6eupYru81
6FueI61FsZrpmQakZLYHJiAaUAjKbQR8EbUr6440EjK0Zo6Ieh2GytVeRUoBZLNndxdQaKm4Zr1o
sZTs8PSpfrVV/IoMQ6vTb0/4+Hd5oXm0bFxKyEmyJSQdw7Q465b5Rd2FqvKU97W/HSiCCsS0xl4Q
lTXBqAad9KNv155ZQMxVg61XQBs850Qk0EFs/Bt9EjYxIlR6uBjF6hrRD8puzrhCpAOEXGGz3I+U
Tjo3Ybh+x6HfBF29FkkL2oV2yGv80HojLOgHzksVXomNOQRaErhXpkGhcYq2u5wxlaNZs6tStVxP
MA/5nwRJXdfWeXVINqIuz64Ltal9Yd9/sEAijGw8CmgMWJ543qpbX/7nw2VfYTNHAUR/i670quMM
lYeR5yJExM398gyQuoynMdDDvYEo0llzLvY9xKPfKY9wrd7/XTNjuSi6oTEXS3+WXgwAJM1j6QtV
pXJybbQoqiEfdDhWbHXYMjjEBFLl6bn/2Yh0l07cYhb4RhATMJyk6LyLUAfaLjmGykGGXZnCE8Ah
E00CWafNTX+gmvmgQ2QEZ/jLkeuvhtsSpMmmDKUaulChNjSRYmPml3CW+bEiPWIMBJSJz6vGsVHp
9S1iRYQM3JbkX6PVpAxn3EvM8POERvIMYGNcY4Aj/pmK0yvdP4y5w+q29e/CjXEEv8EjLopMH2vg
eAWgyLiQSGL1tyTNmmzaw/wiu9v3EH2rlQJF6kCPaeHC7czEINgAk3EhdoELZ6I4mvyrN7P9vG4v
oUK3BV6LMP6c0Gm+fPLK5iGcE973f8BJupyxFnqGI4+zJy8XveOdjxbE9nRkrLWyoZ2SbYt+ICp1
0GuthVkMV20+nMvTjpzABDQc6SeX2jWcqPPGJxIuU4MVY+fo4dM8VZoYrIx5/R4Uny0Tpb79usMr
TjbF0as6GWvQZO/JPACZXyZGGiMZx1PVYXhCeXOEFTcmNZgWZMzeuXElwKd27Bn2Qh9F9Qt8ek+x
78RoodHExwaqRTFIzNV3dckXH/hWd1YwHxB9wXcq6Gg6vArMaor5+uNuq4ruRzA1vc26dNZIGbXV
x9swrFWOChS8BAsUKLpWNAcjAct2CDNTW46XGwr6USK1SWDMrupfesSnjpCZhv9H3O3oZ21rXP6V
eoGufq0I8mKTQTCAB+kG8DgfQ5K/XR5y93OQTLNXdIbDajCdzSWK6wTfUX5FGacdGGcAB0tMcgTu
9HAH+3cgVf8jTNaAs+/WX5Kp8ijPwdNo8F3B0E1ztYzdiGkxA0Tx+WaLsawVRsYkTsBKCgqZxFIN
hrnkR2NC4m5lUk06hx6ZqUrEd1/2SDY3tzwFvwZZYp6PaNvEfh8vNJxEnszot2buX9fxKZwOVNId
NGP7DOcVSfWnMFSjZr7CSqisYxQjwQIIF8j9s3IEbaurYUT2fRXnDAMjdE8JAzG4kFFSsHX6sizI
sCo/9PmgRG6NetKE9xSYThZpGAc7jYnhliCoRzwHGokig31sFqQP9feJ+jMFwPtXPaXW6T7QTyY4
WnXknhKMsTnwiM05uZHY5empJ9GxtOfmK9Vvy/2l+d9kr41GoK0sf7Xc34udb6MbWUqT3W8Izipv
+rk9bp4TdpaLnQKo6uGwvqyOHHYVDYOjvvFgV9IVJBU0vawuWS9xq1qO0CzdTIzX7ElI6Qh4f9r8
lMwutec5Xt2JsEt1qiAvsYt/sV5zvKucW8TTtc+GcmlTDDqpS4nkv+X5snZCdwu2/ysCnXN7X6tj
z3kbw0baoOUuoFj61nTlkcUitbxX5j3j6cS2XJCeF9ALJrkMSTKStqhIeNW6eQXUF0UiDcEzAvTb
RDDRUjcwGC/XkC+tl/hfMgmft3hEuh3v4chy5AVmHqw7Plqxvrq7n+drHXAaEqi4ELHmjD1Dw9TS
LA+j3cF9zggzVYVYiE+Utocv699f8HGA1kiLAWlFnC6C4kaL5GYrmUEEPWIxPi1b7HheF3rOQ8A5
GL+5e2aENMvtt6gwCIdHg3m1tlMV+2r0R6Q8NJGJsUKuBgWhErtVENy+wmYi7N58ayLyDDFe8WQv
1rLkf09vt57y0jKPo2/bJUXdvx0wrySb5lB60Q2wclfO10uIfZVZmuHa1dXqsUV6m8AmmNjDrgFn
eE1cWQyNrPlFEy0lyazGVcq1dWVdE9KYo1LMbgFpRCmCk54qUkHvuyaFYDcpnjAZnPypOMq4Fz8o
CbuNXmiLnjmT3dwJra0XI/QLy0eFJPK1YYS2U3JubTqQmH+cX/uUKqogGjT+leHFN2+nAco2Y+SX
uwCPrepKwhpb/79EctlhIrM+klfGPKF4Zl6BPpKlO3dekhqr8zfBKWzgkWXoI33nGajjVAJaHbVN
eBa0YZfH0nVgqRE5ID5U6yAPJYsPYlSQY2rIw3Y0KFvtYFJa3XdFkw03pxGkjIhLs79/yvnDfR3F
oDtRukqOZiZqD2p7gSqreMfYtwZUG8Y7695mEUSVY5rXWEV53Np1MZwZU0OkPJyyVHi3ZFxbwnu+
ar+2s3xC9oS3A3TpeUrHG5EyfgIzDUuYeTXYFgPheAha9LBteoOC37uVWBhcWNJhhS/oai6oedXq
2HmZXXzrWGVjSMEQaD+zTOZYhzVjDM0rw2XNgZ/DgvRCv40vVl80YnsJoNLQCOqB2dfjjVcEPosB
/qozdT081sgijaiJ9VVrxUEXNTHwVP36HoVmEg+H+iB1L8OkGoGGuJIqjJ5VylPK3JgyTby9/FYO
xJp9uwFCLDrWwuBTraPAJyU+zL+SPVlOsf7bJPJvFXwHLzw6JZBnH+QOHGEIp5PPDUkrqlLtiog8
ePZwjhHr4mV5KOoRiV9beUFtyNckZ+lrDgjw2Xu0twRxkcdBqFRQet0xQwto7FhkgprDSjthgaPl
rm5ma8ZLhDmO762ZjWYtF5occ8Y5/e15DQ3sOMJU5nHBE1os0qFagVOMecm2OREziMzJTU0WZXe5
kVB1pDujOzr18v97dQ8wNZJ2O10LFoAFOARYgLqcf8eafTfirupUaRzybRs03UiMqoMf+pxpo2L+
SMP5fql5OIWVaLK8WijCqeazHsQnbmcv+Ft4CpoGivN4r02F9YhOrRg5tqb+/dNNxINFaw6GT//t
LDHhdAn+hNoZl78OiBsa/bUvxmqCplwo/huIj97Lmgk0YNsTsWsag5OaGap5mjaMulbge9tRWOmI
2qA84rKBugfEOd0mB84esUzIR0XyxWr8NYCuq7fU6XaDNSGmmkzg0Wq7MfJrn8PnY0odYSIl7O3a
gGpBMBa7DOgTXZ9RyAgI3WYakobXdv/IAHYc9te5zS0lugybJPUAlIt3+HOissRMdDhvtL0/+qQx
EEh0IuTVSzgiWAGWOGetynpVXXhuZyp3Xr345KkLDLyfsjr6wq0vF7DvjoQJ2lNqgMQRs5azxOjL
gvJXGUtpj6JcUk89RISosvHa7zmlKcMIXQHrYjllQBSn2YWvi/ns49yALcmV5pK1BR3BXq6pWhad
B8aOjlt9k67wD8fnpaR0ZptWxkObduND/12MlqF90b8LhoaLUhi/psV+/wBNBOZnKHJKcAvcQQ+r
Z0oCiDA5I2psSy/7/a0Jb4mxl+Eq71KAQ+hSy4NwedF6qeMKzCNwvjLzbzzCXYf8LL6by1MzLCgr
CjcdUlIysWm5tHkKP5smc7jVHe3gkdgc6nNpCTM2CHOSmgUlUpS/ag4FndbdqDlPbCFoTzP0YPVA
v342odnIuve/3PXqQH8+r8e7GimmgJylfKywphcsSepPxqKa3fsxHYBgTDgxjTBtiaTRKKkEBCNL
AHLRKWCnvRSwMvzgT3hBDFMOFoPvAatV4+OxyAne/qbvK7raaz90JVARs1eANgyOJe/1p+WPFNnz
4dPy+6Yrqxnx08WhI5z/fVkixK8tSc6POapmWYpTmLk6BvQ03+OHWLLaU28c1MzQZJJ2519cBfpj
CwA9UXzz3FpZ8nWw5/PQy3AwPkkDjf5Jz7IwdJsdYpG4D10EVV/KlDQZ0qDbwRqNPw3roYVU0amV
Ms7YZ9kr0NguBKzG6TAHg/bVNZVpdbLLs5idSRVcP8xrFwiWEviL24HqmFOYX22iSEZ35QmnXPQz
r8SzN10igdbr7j9SUFij4vTV6itpFM9hDwQpt8NbqCy9/8PG/6ix1EbrpbC0P4JNUP05QlyaJcgB
6JGvRbHW4BiV7WfPrFQBZiuu5ddu1MFs+yVFViN4XQCgx4n4TNp3w83fgUWBqYx3+YcXbOpqDdMx
/BUw2DfSt4fC9sPSmBA5GkIhQKwPYmkZZstMDkgvQ1o03fsyfod+dBBG2BRh8JR4f9GCOos3CN45
GvlzWygvRzHMwYxzQfHJqCF/pHkUdEtkh3ghyHzAO5ZrpmK2KItVXMPO6WK18to3TF7X9vrFjnUC
vi+4tdugkY8V4nN1yp0EZ5J8WVyH3YVIHPe8VSLcc0R1R4eRWWD76qgwrjlLmCvdG8nvhBUX+CLa
4MIa8M+HmpHfqifEZ/OZG14av+gb5rUYKffV0NeBBR5jUKaQby1nJC4uDbj+C7q7Me4gIp9ZX7p/
FJcRn8ljhV1GQLECXcg7q7fw3YcdoOzRgQZQ2N9A889XXG9REkMz8BbS1T278WllvU0o9OTqdyn3
UqVy+k5SV1AyiNgOYV3/T6YNzVqJT2/b5WScC6Sh7Ld+p4bmrZB0hPt1pYbEq5e0YruvZYY8Jwls
QMmoxMg/Oy0w8ObUtXpcS0z787hCAFB0QIIsEkP/GmFBEnVWI7Q6RQSDUkx9RkwJ/TturEmbziC+
thkYeHHMXsZ8MzQA0P3xz33KmvhIzQejWf0yk00Ol6A/TZ2Ju46AR3vrH5w3sAoqc3hTbesTHC2I
ACKcsG1amDUrRS8VdmGJcjbLIk6wywsnIRGmJuPOoxgBy5RuiWOzzR3zgSaWZvf65obVnx0C2doD
4+1BXfvdeJW3FI6R76ypD0ONoGj6sJbr9Sz7wo6Xlzap6YkZVPS+j8LC1NoHZ2LhxROq17wgv3+F
1qnTJVUHdH+j2yvTsPozmvl683FJRs5KnpenVWTcHoHassGB0mv+UnOatXb2aFrw2Sl631pK1RmL
7vQgTUfTnlVBR5Of4hEY/q4hydycTu0bTyNd3nrUvdtKF1t1Pi5wZiqzc2zE78E4f/FQuUsbsWN5
w5TBCtX4kuon9EaG3lVAcbwn8Sb3u5zJxTyuGAvg4GqIJvCm8sfJ3AHYVpyz+RCoHmys70Edw7zy
Pm89NhGVMRS76AF2w3mPtjYvg7mVjM4qRTBbjSJiOzBc0OpPcprfZh1HqdUlCz700O/OVvdoYgTQ
C5onhHb/VoLOm+crJM5ckRWdW+nGjIkVPx4zreAM9lmqn5BuLpA3KEBEsXBdWSVS3VIV5VpHJsWF
CXpXnP8/CWxy3rUlMerIP3CDbfBPcl4NrmG+WkJeQkZOSQVs0/4GoWij3XtRhV19i8ltwLanwmOp
ZDlkliih9Y2lzDIaB0nGE1fd2lVf4Q4ZBALic6Pndg1VnE1+D+JbqZf7K6RMT8sX+W4s2FlKrf1p
pCz2LwsdGaDj+mfu3rwVYtvezfJLFc/m41xKWYnC4Bzf09v+XiM2cgk8eVk/+gkLbP2kUe8Sd4bz
wqapJAz4nJcoEgya2uJK+yfnwKWLEe+a05PJyWCfMElUGRzU26Ew6qiBBZwF5JAzCdcPLhJVeNzF
zI80RVVMX5AhkbWadkJMgPmx5Y85BzTHwjWn2QsSZREV800w2e6+HVtsfVVzb394BHNzCxoVjjMx
+cm6uVY8KXMWjT5ewc53odKklX2a6PKphGmKOTxaJbCcagJoQgNfFdaujrfSS9i8AMNowgHgXCfM
vr/i8NTuZ14H2uswhLIfHMYbjaYHLWUjm2BM9CnfRGUF0QKYMUsWJtAomJV89Yd3YaTI5rqEuBhh
KAPhOPUBtrUOda92Dw3NDj9TXXcsMWlRVsS8lxZu3b5Tt66CJqgrTov71ggzUSZHMlpiefX2IQIb
kic6ByCegCjxH82upHWmhMNJFmSUvSwILAku5jaeNXMg+wsddm9ICCi29gxpRBt1qPnAXwX9VrKF
xcC6KOyCfCyJuZ0jJZwS+K7KL9qFOkjdzKXFlgJK3CP3METVoiJC1m3Pr9Gg0USsc3PbzPdgZgf9
FuvaRxJA3WDvLXCg4sSVe1Z9UNRAFweHCLwE8thCTcWewSHQ4ezzNundHDf8Lqa3bhPYtFcNUdnC
0/bU2+Y45phuFYMucDGaiYZ4YOtiuvOsdlgRNOPU2OYoRy0/NL9JSMc4Erg4JDcXtCtNu8WSFNIn
83apptM++k7rI8mnn8T5JH0+OJmFc55pKZK2zJ2DzSKGtpTLG3uT8HGpJ4GMnxOGAJ/m+M4gCZfA
eItsQLB2Y06rCz8AJ4XkjVl+JZIVoj6eyt/Prvtefn+7hiSY+P71H4LGOXQU61xcFst5ZAEJxtR+
+naT9c/ib+kEUJYZilheHjwzoF5X7STWNqp007kMR8EqebC8z5wK+OP4d2RMaUdDcUHczplTQy8l
R0wlefbpMFthqJ4zq92ibRFr6lGqzjzVb9YwkGGgYcwgiibIomFUTyhtt/ol9LunDvxJ8YNzD1iu
zt9IJMP6xLeZYmhnOVZq0xNXp7e9DF0+2zrM/eVbpC2tfb6NHTJ3bAFU3+8QgEu8BYhc4dniOO53
F21UxjhrzE8CRMsTVij8HfzqrJWZUqlPNrfFOzQFnHztnLebwCWSNBxktPuX1nIRM+VAHI7c/ysj
dd2mp+RvyuYnIieo3hGvJAD3dI/t57XpOIAPd9u3KGdP7fXMTOm8HeAKcUFxCdOY2QzXb04FRAeH
HBD1velUSJfkmMKhDlLkYmul2zgsuF6dyfUnrEPEs4nYuiuJOCFhafv0LAwmG7zE5zvokFRgVZ3z
e5bpiRXiOdNG2/xs5QRUtmHXHd+oL6MG1qa65O9vQL4L903DAAzA3o/RR7b1PePwclYdqEsIzeNz
1c7Sotg9LR/oB3303OS8q+PBp7WPlcTmAZPmPH+7A65U2wfq6m5W0Dje5wen+HPze70YUznh0oJx
Ow2GZJu5Og42s15gmtgnBZsXFEqjX7sf30oU9UwjckjKcR15sJIdip094dZnu/ZeXmRd2yI7tA58
xOPmQ9eiBDigTzATSbCG/65F794HuULNDPmbcNuBjb6AB2DXVswJypYsmdxhuZvGzbnp8L4UdkRG
EfgfdZaaFmqhXrlmAhZ2BeFRvmVmcPN9JfljbM9KrA/AYzctSR7gFpCGqAiHKsu5CRtzNy7wIjO3
+y3+sUi1KwaFqMkWTm/UaVXIYjZzEtmMDSqggmsA+CuRL8US2lX/5DS/BzzRFMAaTPo6BnfF75Wt
ExpRWWPBM/lCle17dVy6AN03Ix4+txQZ3IEx67ffkAxpv5lmWFMnh9rgr8Ilke93wCT+ac6E4gQG
ePVljgFbZjj6a5IaG1sInN93oDoamZA04PZrbyLqEQLrXvY9T6Jw8KrHlXPzauKv2oPEUG8alK8P
R5Ivxk7OxXDhaXUduHXo+CDxwLs8ZSbEqDNQkJCLAPJbdyniJVJjTixFx4fCrWD7OwzbpqHs7iuI
VNptI0ZC98It2oioj1/mEDsmhLP4fGU3ucO8EbYtynnyFAQRHMSEMgVzo1scykRvIuUpeAC2tGu0
kdgy1Uatye1kO82m28pkEiEgdgrg5t493K0xqF7S9k3iXsYd6eqIAQzyqwNjUptSBVxFQrI+XALb
cW35jAYHr7d+RBTihgUTmRhtUlnI8qeswquI3dB8avyiBCXO0aWfuGNBfAFr7gyxyUXcbnQ4H8pk
FQhDnj8jwuSZECiwAZBF5ZilXPN0GMws9mAEA0taYYwSA91rc5p2PE4APN6fy6M1A79mn2QuPx9C
p7GcvJ+kdPFH79EkUPUYtEVwkCkwfNlInkNCZ8vceu7crSiZRp0SOaZCTYuZRic1JHNs1DesgNWt
5MC8x5AByUVrX8rVCoRk08+Sw4Lr8yFTQf8vlEi5YKo95bEiz3/GukAVI2wyWmetPbVG/Ep7G69i
+piP7Pj0AXun8g6crRLUCDEkErBF/Mz3QwGQB7A6qw1nZ9IayGb+kQ2nKISQXS2v2t2m5BV7p2Vn
x3dMopwmAImKYyPS4iyUEUBuKT9Nw4jfRp63WVsiWkp3iLsNsSKE5FTX1jOg4BLU3biiHbJSmt+0
6+GMD5Wl8/B48H5VvZks8XgxPd8/XbkYAE/ZFIZipXOTUo8fTxOhUl7LU12KcZa13mZBdl67HRmu
dUCBlb+mxry/GDjVp04QkjfL8gIPlWeW0SC+ux4U5grY7uRPF88inJ4ZK7Ek+naHb3CnHrsgRzVK
v2U7NRaCWR5ubgaBT13f70LQlMlTbvQAI2weH0nSgWWd2NMKgpe5W4fMQt7CGqM4uujeVjp/E/N8
DoackGEIdtTFTN6AwtivrWVVNUFjDTIC7TAucU614R9kl43oShLhM7n/ZFJIi2GmQNnzqu162TkX
C0pPIGwHpXkTcOJ0dLgfH68MhW3G2sv+Rsyc/m8srxLgsL/V5ZGBOFILgDKJssjL1C1OSNVRxJqF
ajlerzzeHNYCIhXo9hBipe+VnrupvBI6mHIh2LOhho0Y1+DzWjjP8dGGKuOsRJedAN4+ov5CLu2l
GpHZw98GbHLcxjZ/0n/FCFUJ9j2jbnCTWJ4MZvfmWVIy08skNkMMMMpKP+UlO2Z2j6acLVF+edBE
xOrR+xX3JpThfe1o3bZC5aQDryEbikoROJoQ25j1TRpwIWpd1jZtW4jZw12Zbg+51Ywtdz8iVrs/
f00Q+3A0/yYEbdjgswIaxYn2pI753AgjBXKLsPN166zwTQbq77qQNoULig0z2QmujMHz96RewmjC
7d9yPkNvcN1zbvPhVebKGbBpGEgEgza0snMBymgQofyaDkbfrPfW1r3GF82ivIXvOo8hMDSCAbWx
5f0vQUn3zRmbejLneFJwH6pCZntC11Y0xv2TEm7F0AuC1VjfhquAebFqzL30iENTW66WcoVMUcoO
f+YITBaVLjXzp6n+B8dSWKT/16R5f42+RXa2JOD6jRJMIHO9LmsQcFeJgJl0CuIHucItPDSHQXZE
pMXVx8w9BaUGAqQs4hmnL5XNEh4fdgCU4EmjgaVeltNEoaErcEQqkBJkE+eBcvvS4v3np4JjMVVG
CP0FYaMMSabjJWnx7dCWbVgi56lhYt1dqq/NvWLW01Co9ffFir5Yi882b20ipCGjoOAnuh3k00Se
RJeD7KsCd47k5JzoGzYWxW7b+rAoBPNTYQgRJbu4o7FfXCZXyz+U21utNvPmLD9V0hCgZwkukOMo
Ssug6s7MlI2olri3oiUZLqeRKx+wJbKgPDVTrBQeABpIsRw+YiZ1MjIDZ82qUBF2SYgG2Imr8YQG
cb93XrrClTphBjh/OLa6Gko8A1PqEipmpjsItWahrluhE5pNLgOmPKuVtQ6PSb3EN+hccSOp9uEC
PssYmsm8jMj5RCSMAlAqbpMjHcLG56XFvUNAlOCMJo1HTLzS56u2FT4n5MQ0nlYDdmZL4TQ1grYG
NK9/n7qkzcqj0okCTFKmD+q7opKfH6X8NNQ8e3FXNl7Igz6dwevxwIdV0OI8qaUxvnn6wJjPYgjM
FMGpcEn5ellyg2I6z2e11gLhXyFMAxMzC5a8lnHh9I8MtQv4YACvhZMLrfzWQPNViqEGu1v6r+g9
cD743GndLbB8BPMUfiu50NRIhkynMmhnHArTyQgI+kf9Jfdmm/T3hgNy/twppr8NE5EuQV52ZzRa
k92/VxCdKLzLPhwrCknaLvZRyiOSGm82+wm7oKsn4876Rq4pYxwtPPTNe822LFYASVitgIwXqKdR
32q0hEKFrHT8mdhw6lzxG9hJYxj2cs+5r2ce/cmeSXNet4x5P9xRQiVLUVdOIMfKIxkvP/zZ7f9z
GMzVvi/4E0h7061AxSFc1QLicjRh0jaqJVsEv1CHjBaIZpZD+bhuSSmfsL9JAbeMulMFryFFxjrl
0ILgPfzg1kvqLg7l6En9G4HS+kT24tyEAfqQfGoPXqE41gkN4VUMSSjGq0DMsIccfoK5BF7mNXw7
Ya4lTrCVUhswqt8a9IWa2xvHUm9J/iW4TW0TvHFTF3yhY7jgw7h2voPexXt1WRYoUIi+fHkRedZx
vlEg/IOrykHHIFW8HUVydlUU7tKkaUHcchvBn4B8wWaE3jjA3FpSJ2Fxt3D5t84QmnLrmtaWibHV
LKsmAI8PTZWMUOc+jKsXNuyfRLSdWAGRzfKyC9a6rbdjSaF8o7PCex7K3ooYM53lZhy5KLj2Ow+Y
DyMUyTWzox+ULaoGc0x9eSeAxVn2/xE0zNMZPTgbG32GSkAvvCZtu8o/vQvABCMms7ustODbK6wd
N2+KGLGfwuTLpuYjACkTl1JKqAyNGOkmjTqpT2SeAVKHKwGje4FjbjMbbZSNs+oMusRcoWxWWuen
pV6dPMmX6l3kDAo0+dvm73wfRKSh5PnRGJA6hNf/jdIPjmfjg9o7+o3EfR9UPYsmN/zmDcy0pL/+
/vmu5Dpyx+eCcG1aoP28Nw1fudCywV/+l14dWjP7dnIFvIe0SY+kc26axmuxO1oKBdTO4ZvHOOgf
YGNs6ZKVMT5+OaaKHkLQLMP0IIhSJFhtBpnX1QmUEl/zq+5x+IaWEIwUtRLqMbpazqUTYl7WnCrH
Ep0x/PE1tnNI6qv4Jem6nOG0NqeHaUfPEqAwXJu4hGTfD6cFDHkLcl1p+lyT06Fomt6d+VDZ455B
GjVpsEVXPke0WcQma/UcsByU9U0+ERs/+IpNEAQ9hy6y+ZXbrMsBlDo8BeJhqumX8UYFpmGbfbX7
7AlCZqwgWF4qwytCCq+0EF6tit49HjHvd02yQT7T2V4OXRWk2tDuj2vgootQXkKT+6tF/NAARY+E
wEoZKkqjB6S2gVN+JNmc7KdM9naHM7Pw/1PhjRfBB1Z027vDAgQuyhTF2bKpL1jogObielptaSg/
ZCBQq43gFbwSsGioBhmJIp+GcXh13iOJCj/BSu7Gt9Df0/FNAYW9S7kkdikaBs+2oNwCIHk3BZpG
0HMStnQL0U67tliS7uCfcVpXmUo3RSWsn82uGpy5xTwq0+tn1MaNRNwSj2vdFeC61Axhje6ZPAMn
54MWzOkaSraX2pd7aa7oigj1p/mfb5+2WTVeThIzBplUY0YQhRl54ckZOWCMyfsXQ0s2f9DPQx6u
ehvQU4p+CbqaEoOwqx1OuHrPkRNEJhYrMOTqmcngABvmUMGveRz2fKvY3Zv9YAl5FV22OwP7uSXa
6AL2H+DsU0XI8bzetTEkY4KxGqRq/v+FeehKxX8iuXgqp5JazQZdP/anJN7FvXFdNP7CPZBWsXas
Ldj5R3/YY47x3KIh5Fk5MNF+uUftlDPmryD81IMsWsK7NEXAM4TZYyn4VRrgmX+5jUIbSq6wr0Ja
/bWq6GF3Y15ybdpkxTVnhVPtQ8e9ulsa1Nlt0qIjkqB+vebhklm7nx9BFyBQURPz0fqLfpcFCJN9
7EDnJNJ4EkCQPW9UGAyqHfBzMo6OKlAEuz92Ha9q2T3D4DhW3O2UM46XKm3f1nxd1LbVZFgoj4Bz
mk+UyhFIdoOdIsiJWvssndMZCWF4EHkk8V4jEYGhRCJWP9oTnvntMNhd1xGr6pAtyAuYNt/iS5H2
eWnLte9ancUUxXP7brrk6xR3C25tkQAVDVNC1jFYapYBUhkAQOU1u1Ifg49xCxE3JdEG1GvR4eEz
nZUP/1FK2zcnH+FAzitFBsrQsu7pyAUUOpRaRm1sXFuHM9i++WV/q0AO2Z5QyJICyKSMQVb68Njq
2yxxNKl/5HZie88WcHgCCTjk7btaX37Fta9DveahqO6lQSZKwFDqTtZxplz/7DU0m20yG7j0Rmak
/oDLY/eYWGg85+BINPdBCwfu47SLA1nfo+78h6fuMJt6My367ajcIafo2w8XW/iHxw2eWjaTeHev
bc+yqs/fDzMjP7qd0HTNf9bBS8anobK0vXL/fK334LXlXJaiXKeTCDSP/ERdaiRYOgLgA4Kdl+yl
8gPZqc5py09WIm3f3D0zZhO44K4U+NwxRkOlRNEO7A2AAprvRiZ8dTm/wWnWBEmCLFUyu/8cOpMk
U6t+wYWTV8gmMlck6boAjWeWHvGscQSpQgDUmgqOSr7vwUyBi1nlB6UVD1gW/wjdO6uoJBnrrR7J
8QYARTl4ZlDqj7mUJvFZdxxd88urp40d97nRadSorbhbZ6Wvh4m+4RAJ5nx/OMeZgVsPVqph+1kg
Y/oMPld2wyQTw+2YHe6MLQ05ADCWsZT7HL8BKahLBkZMSUrZ7FIn+EmzrYNJnRjqUNEnbpNgIF3a
kPDeo7qKO3IGzNb7UzeZweC9zwCInTzlrYBWt8Y5DNOiBNPCGa32jXAXK9/dIFwSdAyXU9cPLhtr
9nK2FtXr4gJHUFGyJfbhAgRo2gH3c3C2gQcl7sHtyNDHEhy85iX8b4JA/qb567m24Dscfv1Sj5X2
mrx5qMcr55R3mHXC5ZIru355arEurqSxhkzZ2FabnPm8S9XbssT2w0h5qbPu7dbeMRrRPeWrpfZ4
tYyHOYT18jWU4swZ8J5GrSJ0qepplVBF5MMfo8cG+liOhJXS+jUywNhOlK1Q2fOrfMpjcOIPP3DG
88UL5Hwxo7o6ZjKBJcshGm4J5VV4EpzEV/OtWzzOh/XduFS1yre9RxF5gvms76N9+d3uDkluzu6a
t5hvK4oYcNrhHX3I3hrLex+V8daLBQRHYSa0QaK9EX6yGIoyMRxud5cXY64qg2kWRPLCEKYg29Wb
YTLK+z+Yy7g9R2gONanr0/Ux4+lug2TBYckHgysmFv7aodSSYXrQ+MVGdd15BWcDgc0r6OzsAWqc
dN8tvGLzF7X4zpt6b66YLGKyUWpecAKXIRnTkSjFMfHWLehwI4NlZ9mcejONACoNC3vgGn2lAZY8
/H9qQLKKrg3lHUKBHJySPKpU7w89MLwDbYm1zfsB1j3h8uzwVB/+CAOEspUpwcasGOOTWBAEFceu
aDmr+0IWlswYZ0fLwW3Mnf7Sfc72fabQddcJpYn3SHpLtO1iNirCw7KF+vlKC6jYQNCFzgKoxrRn
8gcJAt24omMAyUtbLUYct/ByfugAb+erRm0cNfJi9Xz3RSnW9ZMWPsq/NBc8WRZoOHNoYkspKycP
a2e56X93sn60lwfI60n1hBJ8Y3Gy1yVie/GvF7R3r3qTHO6MxP1wFfXbl8GBncpQbiurSZ9ug0QD
9XQICF+bVitLpQfitdWHqQm6DWglFSAQkRoUbju+FBP8HvEaRZY9zB/d4EfAM2rhGAiu2EdOayIG
ti2h5CKIWBa9fHCSBS7Mf2HS0LD6dUNSdyvl6ueOGTrAqaBJ6Ple41Hil+EHROp8mXcV8Cl4S6R9
Q8h0a80DbFk9O3pHnATol9+j44QrBakHL/ZAXKuvFAXtohoZSttkb8NWD/mcIOnufpJ4H44RJ/TO
zriX8nLHLSAcYpQI6FLR/jV9D5ExIwZWfCTn7J4EY2XDO0O1BuxcK8dnROpYT8rbxv8hjZqq5tSn
L+2aO+RaaCVThM2htXoXUzRJ1W8uUjA1FeWwWWzrm1PS+JluJjrkVUfZch75hlwqbUJtLFZYqQlU
YqNLUToASUHaVOFhy9hVyPKyrx8TsSv18fSnj3TGwS3nEMMR7H4KBNLuS7kLMLAE1BOt0Qbeokz2
AI0C/LYds1+6istPeuDQAwXFDQwtSP9uINnel8XcuX718knAKhomHmuKokIRyd7Y99R1UC7/1Awp
5wjPtFWXe9VwnWLb/l+68B7SUJTjRHYmoyTOKmxT6Lpo6dgs9iuVJCyLcUtDEaD0EFpz1ulE3tKd
WwHw/WnDkch/8uaT4/CLTZ/T+UnxnXEak/mo9JiUzVbKh8GhmgDGOi+7tywh9OraRdV0EyOs32jA
TGmULiSGP0sDAotiSftsKXC0u72+QjhSt9rxq9DwC1rRhb/IAsmBibtk3p06nRPPdXrhlyyM04ct
UC+39waKz07kuvExB1APKORt62ceCSYZ5hUzNYCe5hY6x0MlpXymdtWUP8gQ3Ao0+xD3TVDQVscn
anRbW0xk59JMOdEPe9I8l2yrfVw8JsGyuy1OVyEpIL7EvAJtlCjYnxaMlxs+YUJg+ZOtNRcavMxn
uKcvz/EB7/FFoN1xl8TNhXpyCexkXelvqx8V+PSLRgHfKk+nk7blMQ1Db2AzfUGbRE1cZs3KRbU4
vwKIJwFASeqNprv/bSYHQAGJr7GlHqeuA/hokOI5L3A+Uuw24ZhJAJlNNioLk/LqDKqBxxINKYs5
AGgWOYQ3CwXTxS5pNmWXeb20AThBCIp165hsZSlHahLgMhUd05WtJW5qnlrGd42Q0M+E4CFuBPGR
1Xw1vF2EXXL5TzVu4EDVQRWGTZlapZGa8rxkeovhsNZ1tpfDKxnOo9TbcXuobOdUGG1H9ILS3K/b
+pifOw1Q6F+YUt/GBJkkfV+/j61zNLKNC/kdMBemtvAIju2OgZFvhyQlF9eD10/e1ZLwsHXMYECk
irumUJulsCWukCj6534COYk3EvrQXw/wy4m33Dk+DumQ496NevvzfdvYigVY0mA1s7k/6mogpDm/
is+P9j+mMZcfDKCUZqVI8Cgjky20nfpM23ED0j2si0fMa286Fxb8Vk0UmOPQNZsZp8+X8cO2lwhQ
wQgAGWNsonG9XSqtFwVZUOzUwKWFd2kOxNEFCwRAm+HGCW+hpJpSNJ8QnBgpHoRP+pGDgzWvLS9N
0vne4tKvASSu1lBbzHDgR4g72pFt9oKpEm4KIu9CahMZEGJJnQWSD/Z3iMH0G5cZeKNUYd5xpHRF
J5AsGxvvRWtqDaYsgNupxBdM3/sx83AVRxbUnfpd7Cr+8a3oPYbYBnLR9kT3bnbv+FgzXQA6HSoz
kWxcq4WBLhH37fARamodvuDXeeH4vGMOp3i4CUz78MmGe2Uj2U0MuGjI7sDn3r4Eyq5HP2Q7TldE
AYgDQfYrscDd4YTzheJl+hjrgZWkrW1j9AuSBPG4/ncFUZs1oJSqIe2uT4TaJ0VNk0jzJu1E2nTS
sEe8tCxh8BuZ+P6gqlPG1raOB+9IU2/44q0R0bX+iPP9f7FLd+DSTiGCd0AGHhfhxV+wgclAwJNs
wSzw+zocNQh60yCPTNY7o1YhLmJ4A0rcsc4AwsXXxQz8yZxLIeqrPEb/+XdDCai1W4kSoysQ0+TR
HafsvwBewvVdT3yP3QlKK53zlYVjShrms8Hvcj7II9T8SkmYM4V+UoS0UDu4ir/H33K42PUVF6eE
NahzNY699KRGjzBIqZeQmHcvZ9XFR/kMCIILRm0/WGC7zB0U8AAWx1GAyBd7tT2keEnE4aKKsKn0
K/569xBP0nyDzDp8hq6bkUsSEvLF5g1yUpM6p1msqAP1kGI+pYF85uprR+B9K4U1LD6PI6zFoLc9
3VcvFYMm49Q+qhEb6IMKMRHG1i76qZ7huMFCdz7kgp1dhk2INwfXS5zQBcCSiLrcJtQI5aUugval
vChUJr80e9fInIDTiN3UuCy3FfH4xW+2KpaBFsExwoxkfWR9tfw3RMdKVCLFBi3rfq+qfkbCJre+
31OQvviWfPFWKc8PX/FbiAMxbWjYuTT8Yuc5T8ot376WaV3d3F377fkXis7Mlxn1kBsmIQ/tmTuk
hZDmyaaWaJDm73XIUZDRx+xF+lv08dBRSDCsMRQRgGy1dpWA5DAMO0JORRiYaU58ZKXOm+E7B/iS
dUqqT/fxTHFbqXTlcHtMBChIZEG78/AvXpshHJg3vFi4m6K2hRJ85zQyKN5qBG3ZOuyVfEIkWPL9
AisZToj+5hIqo9PdTVeD0USuo5uGjHmxSl6gSYZACj3aTP/ZK6g7iREXp8hYEblwZSlE8o/eoFKr
QAQgggzVWlsDO0KypIbMpiVE1h0/fOqwZciNejhRjBMQg1Zqa+xDVSKEm8KBuEiw19VqPP10fCyC
FVjtIV/IVC31CteoWfR/KQFlSscWqIjDD90M4jgtHuj/eFUTeOcKQheRSRPP7xrA6EQJEP6t/VTH
qd8Sg253RY7+omK0z6KggxTggrcvzqD7S08mAq1vYoUyucFQWBqH5u4ZnMBs3yG1c4uxnvBzIQy+
sr1a00M4Hj+Bp0vucGU8Vlu5PdiYdx9DfF6/noLJhCXXJxPuTMk19hc2OS4fbJcu3rDEsFTvP8Hc
XMsLLQPu0AzWMoEpEwt+9gNqbmzew1g5U+hOx9/d1z4NE8a1TtwZkarFJhqX7BVQZidRjFjBP9u2
uqX8KdUAKNyBkj4i/c669xlytaKBaulOyVORD8Ym9i2B8MRRD6DSRLrOoJPMVpfhlMSaHNCROJRZ
4ttDp4dxV1Q6O0emmDPwVr4ff1hVkSrGssa6jebIJcZZ1ysyEJQFco+dtUUHVa4RgoGbZRY6mugs
5Mwl9CJVTCcW8rSazr7G8y16UmVXd3U/ihDnin5xwCsYCIDnzP5yKT1vOxBN1iRDf41n2/Bh1zVZ
CANLkK7fJJyeYak+xWHFylwQsCTMu90s6l+SPKvcHKf8f1A82sj7/iIiP5CN7bPjUJJwM0vgynqQ
ZW1OgzZynorR1Hnm+9hL2Fft3OYo0+gOR/TJbrM/hEjr7ZcLyR+GcE2+RXx4WmbEvT8+LE63c/Xf
z9wCJZKWkmfXtu7CbE4mVYt1f/Vrx2odzYJmQHUoLg8+13kL0gsVN+++oUokmtKRuJodLYGks71g
kO9ECp1mzCPhE0W784oBm2yFFPT4s+pIqTS2AAVDt7G3dnUBwUEcpmhhAwOEuzfCRSxBXMw4Nw+N
UAZyaSeXdKbE/hGCVKlga6hH3ZJ7GlCY8C0xqnTeDmHZMGKWobcfBcKedJbbstFI2/t8eXxMmdVK
/mL1Npqog3EJpizYmAJLUf1biIVSET0ofkb9uyCob5Zd2ffbZVF+7r091iA8M/gyNn2DZWi6PXa9
u6hyAOg5go+rfffkP7uOv4zCeR/NfKMcVmpPIF2ovyXa0eMrIedDpYINeaq3Dm4cam3nK/LjdMJD
bmbJW3fmWHa2o7Qf9xhXQv47P+Lop4bMtFgsR/lTe98l/Ca/MfyxLn5Jkl5ZFAgLC0QykFoAaywg
wYTEJrhQk5AWNTK9uUHhzN2D5euO6OTE0venoK1xPYYFPh35DE6tnjFnI8cptOe7FrAPKFYzeZfd
fb9n87OriXP62GUCwFAhwIGK+Pd3QKZ7wbvEkJgeAsIVH5PZvpq35H/tR7ShEQ1E1Xxda9CG7wjq
/nxEdXN1ApOzHJv9VVldQY7Z636jdVSvafZ01a8iWjzgCklR3NK8AeEQ1A67T7UAbkwUeATRD0UP
8G6Tzs17gldnoPVjIHtry5uiE+vSO2Pj+5+v/lVNvyHmMNkvi7L20a4RZPKpMonqKrRDxt3Vt3VF
IZ5LeGeoW+owsQyRrQYQpFmm9g653As9kffP77MxjGO9xJ/Ogi4hduzRAZ4Nma//xFEU5luCUlIL
bGWAUbXaIdJgpamXAWA0IVmK6Jxn3vsCtvPEiuvrwb0n1j2QCEgKAKM2BetVEO2h7PiaxA6nTjyz
E5ndBWYsOUT8bmuRgzcxczlAQPvap7hsnU1RWcMPNjFqnJ4ALTUFnnWOJvs7atpLxB27GCcdG4mk
s8QO6nqC4dcvOh6aYcF25k/7iHRj8qOuA6OxpY352pOxUhcj3mzTq1+CAANUDEz4/b0TuXL6QhHo
q6Mhi220TxXu40yvQy6er1mJt3TFkdfL0iHGHEtJPXnqOI6AKAk0Nz3uLo2UUpIZYcG+CcPOsKrJ
plccFZa5ahHpRnF7i2dX3kHNrLuRuQxFCAcR8LfqHL3fygfkfPBZo2UeQ+YESgg1w7N75YD7qejE
HZxgxXOmIweMon5Nm4w2x3yr/xKYaffkxgU58p4WJlbZzt6OEH3G0L3QAdgBqg9UXLFCOuzUYK9h
AmOOSYI4r5B4S2BMpIo+xPq4ED2yEGfSjKhoqthA0mpKTXVFs2+4nDRm0DG82XQEGqZMfhH8jA4N
djMtPPEReQVTdm0n5faEUHdq4AV9Zns3ypeWnZiAZYoEm2M9FZofXuMDyDJYyvbZk+E/B6mCJD/7
NyeqHBC64G0MtUvlamKCazLZilL9bmhiIpRF1F/VM0W+gtQw9Ev/W+Nb2qdwDQqwcoT4rA5MZujW
2YrqKG80j6rqSB/Uie3KWSxCL975ivilAKeUYg9r5CPmdLjkY48uz2IYS7mWGsEO6xtSdd3fugoJ
robCB6e+6lvf5o3gQaMCkeHJuvMx5FVr/wPJrrCgFROWuf1TN2QRBkdNetX0rJ11lGaceeGvD3EL
H3jNwItl8AkYwSGh8tbIxlPrzFLV74QT+rIRHkfND2b6PY9Q8A0HWqOUsVT9EtxHC1apuKapFr2k
6BcHaixL6y+QgPv/ebUitr+ccUAUmd0iD95wcvo3f5qJoSLuwGvncnt3ppSoc+W5RP9wteWTiFKP
nGpZG6uP8mFJ5Xm1EQA0+0uz5DGLZvrG/I55AsR3Y6fY32jrufKD4bgq/hiQTwQkoCNlM8FWqSij
TshoN1rgb6L+BHEWm0S45jFGMInSfwGXO3mbShIijFsVkn4r3i6ZXz08oQRXNtEezWDThq35bXQl
WFB5exG318rCC033IoBz89p1avqM89Ceb2tNDFvcXCS7sKvK/F1E8scVA+eowKwRuMoQcJECFmXJ
or8NNyAvCodVtJxLpyUefDNYvIUPomYST+DU1Tq+YeHMWJgVUG/o7XsRTgiipVQeTE/t/W5jiagv
g//z9lOHBgkm0JYx9IyAS2nobiL8GAy3l+YnUJBrqG33oJB3cIjuc0gXKRMT6MMdBjs4nfrgBgIE
XPc3E2ip6jmo8AddlIQVCelp9LvZyx9bKM0oDJxe6HXOm4sWU5Dh5rCdPsRlvsqb3djfbqqqg/+S
QULJA9t8kN1/K7Q8sMY7U/9cDLIuqYXeWcubngDntpG0leNs2ejZxj2WpjQhaGjKt143LdEx/mY+
i52LEQJ+f2zyllpKhl21kL7StiCZf01CzNnGvedNo9CCHl80T6Juy7N6eGxcg81uHe9glrVJh9+A
01V7d7x9ppuUo2jznu1pOjhq/5+ASeS7kvihYqHbjG1PdSYZyAecSCecLT/hNTu50mKfgWoi+3yC
GrqqV72cbxFgpXB6C6WFWN3UhFxUpX0HE0g6GAEBhw5QeG0I1L0mB34DwZrUpwfYCNtb0gZt0+yz
c/MCsKH0qDz1lA481FKM2kbtSebPPaOWtL9FnWRsoc90QLZNgJWYLe5RdvHr9nRMOCGCMg+hiVK7
DsRaoOrmsD6DLsHOkbWLfpXPNsB1swQreNu7nYbaYbh+NMD1pfxsAk0h7Plyr3gl6228nrLUVoGy
Q//Wl9hkOaquZY2cPqwX1IyxEBjvgO5QGTKqWAmNgDm6wZZkH7YOwU/P3/4XJpCkxvtyj4yA+EJZ
OICdqMQRXMDyedPda5u5+by1tfLlGuaob9F/rxv74bpFIuOhk8sWa0zZfSCVIKWcNYn0pEXVEPjV
My9cQ1nrdT092rSbTozS8DDV6B/ABdN/vxVZsdoqiEhDl2LfmsmWb22c6aAjbISnWuv5Uo0eFLVm
Fad+8yU5Vq/YYEkEhdFy++5+3NML5vyDn6qXkAizrlhaZW1/oulFdFaJNG4cGa+6XfTobe9cDSlP
DEhosr9kO6prfjpfwGWANsVf1l+PdLGI2lZ+/g0ff4pW5riVOpYkJb4/lihQr9Nh8QTm2MOZvh8B
HivurXzijj1QgareNq9ZCjaShbTrBo1g5OsSZTOUPlrl92uTGUHKvYKYNl2j7tTu8ohDep1uLLTG
dvGqRIXvHq5VAMHeK1/Ooot9qOhlI5H5OK0+qWIxfmUeehiFuMf3S6SCoN2iDaSae1hhFfiwK7rs
emwKnyT6RRLwi7ApAvla2lYl/ivjShsmfbJPr1XDuow7167YOJuegmUg84Ii5fWGA+iY8xrtTuqY
ahM3oyyH7NmlS61lvOqMfABZ1PxBI9dLgHiMuOzDm4Yvfd042KJQvzJP2VXrrC/ROyLx7M3/I/B5
txaAESIbdmGrS75nhWSZzoxDb6kWNUMSMFhOXTz/RY5exBmUF3H9HQCNeHrLXsDU17ZZwTglAUgE
+L3R2tQ96m41kZL/CSdl5vrYggS7RvrXNm/Wj/uMUo54Il0QDoZ4+F60InNh4khdVH7N4CXGdaGO
XCXdOVwT6XT+EwxYlflvTvacdz3sDRSceNM/ZVsRAWkmZKDBtTPoFN591lkAg/GZZxz8B3FkJ+b1
swdkVS3TgpEwxpg78qkgQlxmHSXuvU7vPTDxoYQET+wrz6SCx6cd9SOjtgIUd71shGWOzSimMKHA
iQUVhbJH49ZChDmr8NvihBrAD6fkszKeAAieemaSKqEmga1VQ5G+nj4GotpdWkw4buI4lRLWH8Pl
cqGytxZTDCecqxDicYs9Ca8hZIuRI+hSNrCbnXyu7rB9UC0pE5F2EvK/pkapVjcylDuUiAAZO9qr
Dfev/G5qaQnC8Dt2m2kba1MKD6oFQxpNgnZIrsXG78BOG8CRXHVSzEu8O2j0J7wEQV6b9l+yZe7X
zT6wlYRvHQXGQWYn+3h0G1Aw/SZNWhNxdQJnxExT8uXBQTatTpP+1h0++hn10h9MSecm54Tl/Zi7
m3SGECJUfaUMU8SlZySPx1XYybY/hGW5KK+OeAPg5cxYRj6w/4k4Kzd8/oL67BGNx0v1vV0FslKQ
/UHd73yIjmxWg5yiqe/8lW23ez7xkRW31Lq18rOkqDiSj4O1MfGFHNCPwSZknRKtmXKffQVd8Mzy
EzP59OC4GzN/EEB//DsdnQb6YEJVOqnZUrKkVhICdHMGxthmEaK+zM+3OhzA44v5hG7q1xLnuDFt
+YaaNP4989p6/df2doCAtAqiUiyUfge7jObl3sI+MOXtxTKCgshPr0e9unK3ojmg7qDi6HyE1oOB
9+dabRroMxgmhm7kS4SgBR2VvDmytLGJao951Qj29pXC3elQwzFeBB1JHPAJwQLSxb5rtOAszbfk
Cx/cGALxpCyjICK/SH5AbD+LvY+vI/Oslkf0ujG9hWx0rlnbHgmFPAaZwaYnDSjk3Yc6+3HrPzV5
S3DYi9NxLKJ8SwW+vOdmbYDEGYcEpQ09yup4VBDMnqpDkSKwkgj31sCv7/OZ7JR4Q6cS1JcEVFaO
RrxmXXahs0VegCdyAwA+ViANdM2xJ9V5/NgnHrLjvMH0iO434WcHorReEMJDOrea8U0AxLX6VflM
FBpOKNV9OhYD8A6jt/ZSsLmC7GoSuouzgFaLLDmipo4ubdsi3TiGmyoI0i6zMuBs4hPSUyot6yuF
FsceE9uQBuk5mJpk08UWhx2MLhWnX4N4PXGJhFXcMXatFisy/RUXyqlPcMcTagRnPMIKprFhwD9Y
whnFbl3a9Ecix1De7R1gw+WVU3SEFRX2NfUqLMA9mFm4oVSbzhnYXzm8JgVCjVujjPwlXYm7zM7u
Gaf9bQv88T7Q2tujnlA1L927y9etbkq6z50OWVj1tJFT9rg72ncTpWE7eFPbHOBJh3DMtyvx447k
bTjVwIJgjdDeKyQ7fjSNBO8h3Ylxq9Gk13TfdQrQwV87sYMVaFvgNyPeGbq4cyRleZJhWOhEGGZ3
vwf6c76qZaNlkHAnlFn/42EGvziQLD+cvjYdtGR39VlJ1Cz3GO7hB01Z7khd232uQPrfDEQpX99O
IySwSQjKOXOf5KIaiEHJAVf4AHRJNscFzoF/VBCssx6S83lx3PaMPdUEckwM4mlQRdxsEmHuuMp0
fSQZ2BbYTVomCfymwHmrjOmkUY/C+6JB0tAcB6xN5tB/qs3T7PTaPbNN3i9Dvx+S13pEfSrnEsiJ
FWMbh1W8+pHeT2dPHRYXOcAMxn0VDBpREPEUSSDqo4vwxV+rLPBGFRFJXLd+rlfGW79tDaTtJy0f
7VN1OyJagK2EfCNmX0C9L9E+UUE5d+hz77BtYsgkPL2WQrMIvCJlZaIRbpS/JlKQFW7wi7uVxMkh
ztqcAoby4kJGEYH1BmIJcEtZix6I/wMUXomPAj9e/EdgS0ojaYf27HLEkWgxRpcLlz2mhaxkdN16
XC8biWwp9brGdzN/SFzhaqBj7uJPCgZeejOvePLQkvdpg+4p/vHpX128ZWkJ7Kpc/GkuJsk0MaLa
kyv4XEqYjDjh9PqW3G2Kcmd3s2Cbc7+1leuOWV6dg+SMjqcCnAJ3cBCH8/LChSKiJC11CJNLP4ko
Wwb0dVE5SQU1Av8+j/CGNMAYGeCW6Tltu9/5I0x8/Sg5TJKpgkvldHzeKJKqiaf4tc8c1FRwnfZ0
UChD2TMIdqsFMuru89xD6GlQb1LZbMnMisFxac2i6OfRdrdWZEatQoneDcbfzEsXOa1yA01ulMlE
i8D3osa03KTcoEoWlrWlgf72UTSBxsjaJc8eM/PLe1JF80CNvJMriikefD1JliYvfouOyV9OQrIv
odtD5593GB1JDvVmjAqLgmZltUarI3GlX/nWQQHkHbCI0R72iD8hAK1fSazzaEXPaMewutppJCgk
8KXfa/6xwYtj4NbDeDjlfaD0hwzbvZdI08auEDY2jLH9ZBIQCwwdOqEJHVMnTTHHP/uM9ad+L+og
oEns8Xz89GS1PYXdfL3YWNU2Iv9k79Hhqgb6EXzhJnc7UVh+SD2jya4eZDypTrVPhwfnc7RFMZGz
LiUjZHve3QqFG4R0KEeGTSem854iskQRgxWTlip3sPzUkKJVwk0UChGg3qngtIgYeEcqvJdEdq+i
cRbhPykDWba8+BzyksRCjhTl3WsqitjvVKT+/IxeIXU1R5/wJXpc1BUVXhNZRjrZmLTDLXvQ92Qu
nnx/TOjnvQTS1UXpF1m9YhET8Qay1tHb/6OpqpVFFpKtvcNhsH/bvKqrAGJnStlZG+I1IgU5TmvH
jmc04jkPd/h3qiCL3vtzr26jBPadFECO6l+e08TtTFFb00rsj2vyCAYh4Ny7mzrrtrHVjRRcqBRf
7Kz5vFSAfRW4dULpgX/yM1f13CvdNtZCZVv4OhRnmog0q34N0DbGGU0kyV6RbLhl7KvC92AslVwT
UbpgSwVaV1qKf7jbkSw1dlL09yVAkPP8ObLjFOefJN6aIDw3n3u2ns+owuJzkLkVb7PEW04YzPFr
2oNCuQT2nIDBdtc7pH22i4isS7iwJqhED25xdgfjx9UCY3YEI1W1pNw/E51iNXhLYftrNM3E3H7s
WRIzdOnjIV3Vx5qA4UCu2da9ohW93ws5oHIo9X6nznPKeCG7RB/2tO4vwwV1+N/8mYMDSSgmmvui
E7xhM1ABH8O5nO5kWlUQWD6H9mlefA0XSFM80Q1bk95qQxjWURXwqEeuRl80i9aFyJeH+Q/4DPl8
BS+klQgGVjOkNu8XQGsYwuhgWNDVHdc+4xMirBLn/xdqcWIVYwtjJgtUuAdqIHdC2+wxVXYJVPJ5
sION0MxKKibwL+r8XfFCGFwfNocD9Q2u9Bv46ALYGHa16FgQXSHVRi/B02xhsRFhYrXt+2NKl9Zv
tp8Z1Rgfnksl55ymUEYvuQMUSoEkufQUP9lzC9qFn9YqnSQyQ2OdyXGzKXvTOebGKDMe7t9Sl28I
9eGskGxcHxYaesWzs6jP517/EH0kwJvia/TDxDz5EW/CI0SyyY7CSz1pxDhoP4B8DofdzzGKvt5L
1wQXpvsFyCjj1mHNt8vrDeS8DYogEvC3tibO4H+4/E6ADDT9Sc8s7agx+DE+ltg2NHOT2JpFefgz
ihL+Ahz7xdxnUVc2zYoNLZRCOhMVXHpx/M5vR2O9j7POgZSbXToWuWd/N99tVtcU2oAqdPSczwBr
z+i0m9M7Q45Y48wpH6PqKR77sXVpA6oCjrDBLc4VLEhRmBIA9JVCTurvLnOp4NLOXhVYFR36N50k
SRrAHIQmqtcPTXkGbSiXCozCNBckEwtSVE1SVHtQXLzgcGgjYwDtMhWHy9mZhJt5tndepTsMNYyt
IQvptDn9gDfhcymhKmTqwygeFXgrj29PL62AWIa3n6Q1hJuukP68g/8SfBFuR30XMhWKiW9Cx5OK
zF511oE4hkMJ+IpHxjOqY27GSSRHg/WT4LN5MItHlEG6R8YvHywam4v3InUPEUEg70GBAEJELrMb
1rzsYNiYNBGwGDdasgYnerNpsjmhQZhD2d88YTZb9wF24PnfvvNtpZjKEZf7B5atDkmrxnHK/fK6
EYC1Y0gNGhG2GfMxnVWUI3xW4eZiACXPzzYjCYgdr09yGuFBgr38e8B9muK5VNnQ4UAoLBQkFrgm
zks+rrzjLL4sZu75f33oUMqZSv5TPzkfKyubMVQVTunCeknEcrPO1zasO9dcJJeMH5YMgh8/v437
quCuQWwSthyUqKXY1sawmreqSf0QOjySk3IAYMbSnJmWupf/8k3E3kU06oReawPdfoeRGg8WBR9E
bznjb0kQN6UL6waJsoQzdVEmDTymlNvR+/cyrkptgfMGNQAgrwHpVsSEUdtpkO3KbBUcPKdy9t1p
6WR0P2wp8/py4f8rOwQpj/Y+UiDFVQvEc5wkqkZ2uTWqzPllrQQ/JggiTVIdi0+esKSRsEmEH2cG
JqJp3q72IFmPIFgv5wJwsGSnDVWU8SklPfiFZIMowigCqR5PMhJ4h6wBoA5161cVFi3BmvGYdXBk
0rXhP5SMsD4noD+zLMVLu3ibZx1osi7231rWYCQYA8V7tjWDpzFXIyMjtEsrJkpzvcBaeGwp/lCu
VAbSEpbIDLSRNQiy33Ce8zJWe8732AoaRK7RByRdCHqLcLVNGHy4/JLWDKh1fgnK0kTwb6GN36Mn
FiJZR/oLt+CJ4k1cIHIW11WCBaYrrkAKgDqGTmyNTGg7YYoirXCxvj8qOMvecZ3zRfzVYt0J56c/
d7nCpPic49wbDa5HC6Dgkl8/GLMVshaKLjLmeVimNjs3reFzt8YOZt+DbmEPwfyO5vgtLQ3jbx8J
W+y5dTskmjsjsiybMc14hV8vZf/ih+Y7+ywSlrWpBa8ilhNUvtR7mqYDG789vxV1swiwsLamXQIh
e9Pv6APgUtxKebz2h2cPq1gPRmE61tqPNwmHhn3qAnYUV3Q/TtMG/axLrCssr3h2IW6HK2Fh4pc0
03+MJc7VTFBCr1fWsIYO2X4mNiz438N8SbSM30lgXw9G+PsdL+RvGgazQr79xespewJWsDK3hAGg
SKBG0gvPEZ6G5DRCew0p+TphkSlRPWT7AJkIu82ZSmB1iaviJPEAUgFKI1aPioAtCdwe+8CTJhZC
jt6ud7Zkn+Jqs0W1RoLOMCUgqpcPA/KQXp9L4CVgS5KfCJp4IchpPW05o+AvsdIwpbvzZ+tBKN4o
Knly02hAdlyJ+Yej07RgOKtAjIYDwpG0dqU9VmZlD92JFV5AGmNgdjm9ABaSNU2g9PUqcVyApdCD
u3xCHc141ydnKZn3eZB4vDU+iHB9WWuoqafe3dwhzD+w0F0AjPdnjBHNcG1bOizzp9LBKQuIFwLu
R9XCAOqR1X1H7Ik+SOX2jdpCkmBL7ZjlfwU+x3MLLahzs/uqwIBKDG22aphVOk771GCKFE/FlYPg
JMLOuAxBMUI3QShgbNE4qORU8TCPnaXF2sh9H2YH/O/tKoKp+bSKz/wFNFyK+im7hVKyFx9H1mqw
rpT9+yy5EuoQPNucmyuIuoDQDa6atqPmhuFY3OyA7sxSr7Dw6YRt4/1aUPMllOWkreUBdwpIBxME
8PVwXAAkxu6VCGvwtS/uufZQFvEvimSLqsP0oF/C9TNZhKquRRkJd/b0gdgd45Rm0aNsn55X1VlF
3t+o438UYQnGe6kw9onclsPvcCJiPJ2w0oLp/bLcDh1OZEjd3iAvvKFXxPCtHFTPNFTB+VY8hYfw
TrSBWFQTLAPmKn+cxWz8JckMka7CZAnDLdcJpPuuGz2IzTFQIUF5oyjeiBiXq13fa6VUjFxuz7h3
N2P4XtY6f97108fakFaByFpn7X/c14XO+da/T/c/S/zOkK8w8Rb3fst696UlwjuqDwiOCsMucFeK
JWmYOM0EagTEEScHAhH+YLg6HElr5S6/V182HZYS2YeCvh9P5/4qyBUnYjTG7BeECROCxLdVb8Kk
Gebhj7i+3uzhi5mNMV+oXKhMPuuyvsbiBz5FszO1KxTLQnbwtSLp4Bin1p/qbF47IXY/wVduZrsM
2nKFfMuBdpFpnfhl7vDzho8bAHW1rw2fN+ufmKzyEnO07N4TGmwkP8WAOk3PwxlQXDiprVx0FwjR
TQl0RERuFhQ2ONtxoYrzHOcKhmf9Ps5KUmO31JNHgeqBlZoTQFh0jUJcZL59uNAA+FDww1GgFHTa
QNW8DSKuymIUYISEHAGU8bDspNb2VGYd35r4HQmcVqRL16v5YZUyr2DSNlgij4CbChipNL/I/IGX
GgNJM+FbZlb8gy8gb9hhvx5KMcNZbrouJKSemevVRdfl82z5TdKfyHdN1EpHm8svzQ9EmGU0ypoO
+8MKiQ4sofnbcL3mxTmb5R+C5WEBSIa4ZWIzurzo5pYMvEd9zS9pADAm/IEAXhZpV7w3CCzZEdAi
zDERqU8zvKpTBKx1f3st33lPC6NTn5n4gz4Xo0E3AdVqjRpse1cpkXdsMz6Z/+twYaaq81kuR9vB
PG/EB3Nqz/deng/DNomAwnStgk4BosCDBhd4LjWQyoJzPoqCvBCa5eijYzliDPApojIJfd/k/pWG
E865T/GX0arHZVNv1Lh61Kx92IW4pBtxMXMAJxAvPicbzE2Xux5CiBhnRI94OpBvGYT2k1f8rxNw
7VMhgwTkVmgV+1WebTruVZ2nKozI/kEtx2CuwKSo+bdmQeXlbcgkdSGzlEf+P3ZZ2c5oKb13ALfT
pLltvriclV2a/7AhA+5vDTWv5RV5IzNvLZ7F39AboeRLfQJCzLQqcnm/7tMiNmgHgwxdu1b0fK2K
R0uoz/BwCu0zmlJsxo0fj5qEaU+X2CsYwpfkqGm8YkvGqy42x+n66bmG01HAozrjRkkDv2k3iOwg
eOkOZLgmHmWQ9JAdXQDKpuIljyo45o66cB/pz+Hhjx6tJtZFT+WVXxPiL6myYvMLKsoi+Sj5KiEw
ZN57zaZdgL0VBo5M6x4lLOWO5UrytI4fqCrG0Ei4m06bOlLbr4esvvqbrQjxYbhxQskAqPklZg0A
q8UKszQzAPqnPl6xdipXqjPdjmUC2su1MfoEg3purGjZcY7neyJB4zuYE/4gfudp2DgLUN6oW1W2
LKMWGp06y0n8/ZMC01wYXHBUn/wzEYtKDp/UpzYq+XYDq3+fRGGbiXq5fDEmCK/jcD7FedYBHu74
Bv6uEv74mNJG4kGspjlVt0FN5KbJJgXuxh5EN5knuDR66ju9zXYU7C3XDliLgcY5FwwGWTac3moq
29oO5mThx0eoEQhBcj2uIKcDkUW0T3DTO+VuvJIk3AzT03nM3tUnIuhB5vYH/Xhv1Vr9ufVP4Wxb
83JLaH8L7nbu1dDUmq+TlodsoxAqHj9IzXtGvElpzUK/41znAJ2pfauyrEP1GvHwH4zITOpbUYpe
CjCFuB9S5UB0DyNtLSZi1eJNRtCDLt9/ZmZfJ4JwQVhLSsy+0mNKRls/JmGY9wFZr7K3ZOlrx3wq
yEqsaFEvfPpCv39SonRTgX+sn5aeyn15tXDvUSty0OkwcLAFqlQ2bFugi0yaaXxzPHrFYaDl6LM1
mKqfTZqq3fb9MHxS5ih91OpejpYBGEyxr48Zk8cSt4sEdJl1D+29o/4hUB/O+G4P3LHDVo9L5j8J
hGFLakvvwoX4IL/0YVg72k6etGtpw+/pfnG/2b6gScwJKQDmcQL3+PmuZFQ14na66shIrrN7i7BE
tbfTWZIIlYp6zZff1YbM1/24b213/cR/5fXeuvdWKBraxzSR5+j31Vw8nl1EUxiBg+YIwP2ByeiU
11o0zkK4aIY6bcGCsENotN+5cdxKWfhBZbvPU/xmMuyMwqb1XCxNxkemOLDoWOXxbBFvGQsFtW4/
Luux9hXHp8+0NjLcMveL1bIzqJ1txyYWnzR5UPa2EKw21LA0Niuc5dzbr4HVxzV2/YIZPKTOV1yK
VSd5EwxTnh/IgK6pCHM29SWlKnEGNA4dFM3nt8d+mKmS/o40MCz9pUkLrAJsDWUWml8PBcnVxIqm
5dmRefzy+BS+FeMnfGd3YigYJZqMBEppRr/CnybbO0tq6IDQQGZ5atK0/keAxzoB0R7QIC1SUR2p
neuOSO5C/hHa46NmrPzNyOL9bU/jkNSO3JIoGgP03MtxHIp9DYK9Rjwgj/X13HXPbDiOFDnU+WM0
IvJBh4OBwDCaWffp4tQx5ipeDlxQa6124IMCwDk51q0/23Um5A9GDdfaiCRVODP0PvpRRF4tcLfc
xrR8u6R4obwdJnZd5uQ5E5BQCXwhvFQJAPhCIr0SoTcdxWJvybYb4viMVWooOc3JR7s+sOdrUM2/
ELfKJontT9Ep30kjUqCUWHPH/PjkpMt8/bLvi+fj7b6kXQPBFDiquQGG6S6Il2gNQnalcV0ME3K9
Mmk6RzkKwGjqjsHNmIkp+WDP0/B27BTQM9xtenvbpYNv3HHI33YGRZoCA61chx4IwlH47bk+pBq5
WD/oq/+E/KP0G2D6xN+f74w7va4lpfHqDNOVx5EmXpJGN+BASwI0XNlgdttfIe5Bt+l0AqF33FN1
KPQHee5cAx3Wjs7/fCKx72Gll2U6kBQLcnYQcXFdC8+YEw5XRM+nFxzfCxFm/IxQG5K8KUbVWOop
LwIyz/dGiyp34D8Q2csTf4A4jVf58y5ZRaj2qG3f2qdA7HLNe1fLqhTmNMYQOiwrfcR37vU3jgd8
z2Ez/u52kRFyFiu4elKXgbAqfYuJy78DFnHTAbeo34/s9uDHoKbFJJFBGSIrOThvbdpjM0BGrVk+
FbqgofKS8doCB4Gwzl7kEIOGU/QQG5jor6z5niuQtJRH5Q8w2eSg3LfP1UySOVt2xzthWL6vcshe
7vwmDWTAYNbaJSSFlK+xiDZUWCBDdYShgKuB9pZwJOT6Fgw8dhcFW6nB7JCTPlyZIYtCs4HTms/h
9LddUX0i4b5nZA15gvg+SbcOf3K3txKoykvTytXcgEB8huPlg+saQ5o+HV3P/mJMxKN/vvp5L3zs
R5hPyKQwgqDh0fjOBnfGG/BrF2zlzSqT3zAyH04yaRs0PsoQyBwbGmFY2qv86zzhBEhmr0mMUY3F
E2J0uai7VcgtmJnKAcpXoqfPbQCdQY0KKRZvXf+4E67xwuoyUahcB6XYNNLJhslAsPs21Skcymgk
JzrOJzEekuIzPLv4HpYtPvLHkjthZo2dj84RXOTfa5V6IoFlLk2XWTLNLgZm2Uei4Uw9qafywS5Y
o6EBPez202GnKaySfrDzAK3W3y2tucCfAQsUXDtkE+dbUNobOcIwp414XvQWY3FGHJyX98S1cAiF
Tg03N46HaWjzv1wusiJNc51fv77PPmmRgzNylHaq9/SaqIWYJ7iwiuUnwtgaInW2tkH5efqwxE2y
Sxn3wAmGskE1X+QWHz4POnc6cexhQEere73o5IHxCfl1lHa5MZ0Fmw5GaoAnri+u/j6THOHpWXGX
diBofz0t8eHK/9Mf7AHhXDxX775VJeBDDw43EpITWListsOEPeus8AWm6cvBYtVoCAUwXS7f7/rz
WUwIAqgJYsEaCOrrJwjzuCg+ESik0t8NzSTGwk6vpwC4BaxwvwM1x5xS2qM4Auz2uZ8PZla0wDQ6
gY4KN6sye4AYNSXpYYPZ9mSYYSk7+UTx+OWHKCZsVFt3j1CbUC5HN9nAeDnLavjaISpxdpH3GEAe
hW2ijhaAEsJKGUEPPzAtpVxqXOp9V/iS7/zfm9LAacf9Krnnprkb7GpIhXhsl7NKosekJNaOrUY/
2gbXjckE9kA4tifnNLhPRFstSHtRnLAmg7HMRss1ofE7Ih59+qnHb2bSgUPrVMwz2X1CiHDpdxE8
vajMGUV1AaMZKVPZJVAcqDUroslRvKtsWN0UrexlaXnVFaxToV15fiYPQcyP/loxFw8/abNkoLPq
gnm3XYqZlfZftbx6djL4FaNkEGMXQh90TB9eGf8uvBkK4J7S2pHJmPC2h1Y19UG4nZz68sjb5Cmq
8xTxVYq3wYvTNCwpYpLzuSDZVMJGingY9WMOwmIxXLgXnQVTbbtG/0Gh8M4pv+WksJ8gJYWaKdsw
5ZOw00iw8CbaQ+xL0vWLl/ATG+vj/Nv6Lvu4Wml3N59Q1Zb1Z5iuEp1R4PBI0zXHFIA8Ovxw+Ecz
SRazSPVnCQTTgb3j81NO4XYimkJfnce05c6tWWSEwSwSitKX0jhA+RjvFlEk+3UX42hgv+FdpTsr
Omod/AR/SY+rTqfkMHTi/p8vEevLZ3uaVDhUOkUhIqzFZJILJ5KX2O01UtnvMLH+6ODv5hF0vcyQ
cVYI/zHuzCVHzOztGW6RB/XLO5X9GebhIzKKFEUyZcng9kjMUhCgrMGDDlbEB1qeEMg7+ICMOCSH
MhFEG4bE4kKhl0Vnk8p4jyf+r1zr/TcHEQyFOgx/vq4XrfF8ey5+7qVumryN+DenRT9FdUKsFX6B
VIs6UrO+mJqpeOUzt625oM9zCi7fBWbnSAUolRNzMNkekPBb54eMf+GVGsAU4dT/2tA6grjWoYcl
Ep65NablTa8tH5o8XLB/usM5WiIlHqE3l8tKClZJqIAfN5Ezi8iA1bTIXXHjjXqhOshu1e9L2Wuz
sBXBWQDgy4wLlC1K5BtpEUCQjk+ogizzSdiZH8oV2xWT/UYqGIvTMonTzkOXIm+KHol62fejsVO9
drcJN6qlu47XEtz9QefcuM1pXiKV0W1RiZ6D24RTJXSJ2tHu3RzbopQfBqthoZYjLTHMPfCByxYI
nmgCARo6df9SddNxSkEBCMUY8/jarWIYQSiJWqPq5gIWQkzKY30GZ9F21HIQlkg/tb/vq+/QWlx3
IEv3irEAm139kFsUMHfiy5f1viKf5o1kzHxBLn6Gv2rJjNenLUy1SKErkJskjnTg54XdMU6fwEQR
iXHjQcE7tolF3Tzkyn0xlpFtrKxsgUh5fSzxuv2pDZDbAq4EcT2G+5fL7Nd2ntbOQ0DuOFDhwGkW
F3KiNQlCvmyKCc/i/gaHxV5rOyg7U5qyvcuPezPm2HJqXIeIL2Gz8HVbUiJV2Fy16Td91vOT6aRF
Q/bffoCCZJ+xqwrbPL+UdCQWdlHy31jjZkkqwMejDXp3Ndx4BaS2CtjCLYYuMSnqK2G5Kp8swbHP
fZkhLRJ+WfRl+Cd91Y+ckdKFfdFUfNMfx+WWmfR9MwCIxb29TdSMpj6CTZLFVMJhGi/iQCBSQzGQ
hed5y/UixMQ67qV4f/uzDNbQr3SSvWCItoGkWPzoVx7V6wg1GgB7XAW5WuqdXAM9RLnvDjOVS4za
UQcSiWmmLy58oEJE965uwMAhgWKTuG7lf+FzjA0KVGccbpX4tfY/FZUdE3esX6QI2adZNa9MhXDG
Cb3Hga2x01I3ksiY96JyxRw1ExMiy4y+eTwqqfH7RdXLeiMij7Zk2muLTXtfcUAN9e6X3KMWnTXV
VGVxFWx2Hfg39eIlntysX8vS5OJ/ROBVcClKdfrxRWWh+BgeR9L+z4PfGam66MZY730kqwm1TgyX
rYg7GsrM4hcCPaT/wjWxASjqTN5YKjQFUyk8b/YTmawy9ntEPRXRG8FTlw4UCLfJZkTwUnXtS7I7
FRb/wIUHLepJwVFZ+YI48/KKPmdqglCHpOr/n9zYkuLZQPSiJl9AbLbesFxvjbBIMRj98vzSh2Cw
lWTFMv45CIxqS8vhWYq0mCRDIBs/QsfR9PqHOoWPpFui8yeldMlBZNCa6vhOlyKrMjOGSuB0+w75
7P6XdwV2rqLi5RhDxyhUY1+KhoFw1CO2FKJ7dhBZwro69ddkw7/04VRvsB6QXXgbEfTELcG7Vr3X
22w4It1rN7v2kP1GAXvz8TzGV3nA786tMSC+FgaZM2gKwJXoVw7Je6/VmlNrg1Cf1ORUbK9He2uj
sZTceTnAhZfEd6dxablXCPX5LAdDHtEyuXot7MA9UVAeyhl5XLWsM//QfVeBKJYZ2sYsJVnHKPxv
roIs9LXd3vAmJmYjPnuk2FA6qiPZ2wqg4AxxPPJO69n4ogldhLyDZE7i/wbqFbZT1v5KIHD0EUM0
zPZ4MFToYh3VVj1Z9SSvHJ8dzvvP3pfknD2xNxI2JA/KQHhQA3CL1Luc4zRm9jDrLp6bRoKS+rDm
JrE6jiflZ6vgZE2SLkJ+zp/YV1UM+VMR0L/nop/E5vcNJi/aOiPle85E25vNPm0g4QaPGYGfmsrB
CgB9G7u/jr+z8R2fJDZOVlN3bhKnWZqaz9YM5gOgw01W+WRfQDQLbyr8Uo0YashtYJ8hF7F/zjSh
+mVz0dduvrL0/x6ZvgVz6i0BxdNCU7q9khDrhbO5xufCdLmudD6ajPInzUnQf3gZQmr+MQWuXE+3
ExIowGF3wa618hGsGyE6QDAjq5IAN3inRwas7qOq3ySykG3edGqOaN1bca7gkZGAz++MTQCvlXp5
Wf4LgrFbUxJuDnJSyAjogQl+XZIuQ/mVBhnp4GDjSNOvWGFqL13NhJzMw0DfJdxd5k/3zaWeRilD
HbFsFnvogWE53IPZAZKj6+Q3mXq3y2463K+3i1FXUCJMz50FpZ4TjX7TrzA1sTNdXHWDHI+sxzYA
PjlL/LzTQAsdkl97jdP9MDbDwoxSUoi0gDcCqDQtCVCZnlWIhIMpu9Dq+3q/cRCGAgfSojJh39Ld
JRmZcR54lssZFBcNnLEHXdlba3g72Aisq5XSQMCRl3Ngzf++XNvv8DXysCVANxgXJlXNQyFEsI9o
2LlokdHl8Na9mx+4vCwRKKmu/knqIALLKtTqN8UemxMe7e+g4QDCvj4eVerzy0GpCD5QjSTG49kD
wwd6JggP6nhrahY8J91b3wciYKtyrm0ZU0u7Tc0D0Wadckw0EpDRefO41/RuPcuyhi8Y3YCqLR1x
tVwUTtaYbZish+rV/n4cqrkOf5tcfRrONcxp65flJipzf1katy72liGWbbWe9M+l0IgeN6AqStHy
oZr0i20qs+Un+ohJTUaV4tmK+ZCKQYDW3jVgJGAfpfBVSvYAFD7VZg8zWBBRT0bB9VRXsyYFo7hK
si1bSVApxI8qJcq2Q+rTc5MzJLPGmQXqwbvNsG5ZoyBmjlTBzgHN383aEZEK2TW8wymNWLlsCqkx
/4uAXFchacDSWnEAJXwLVCTdYiF+hnWPepsiqIjw1CdVBW7ce+U4k7rqHO3XcAyTk6rlkGd7E+kb
MTuVoFKOqRKx+OvehEQkLc9A6TNF0H9s0Jyypn84JhlNjl/Kj16O25JRLevFC1kFXtNE2TQkOAur
w2TAtkMu9pN5jpMUZ8u2dwNpTRTT3WVqxSvShKYzgmqlwcY0czsiqfQQbvPmssr+SXc7ok8ZIlKz
VSzTMWf7rQjddcSXSCEldiN3vxxzz3Xhxp+rL20MfLs8JcffeWaDxfEZSaAJdU1pyt7gcMHPsN0R
ChV2BFL99Kn3gu4tQSbhokppxRiAliKA1IUlSLJl3K8Smo4jfFQlTt7gks7UeS7r5+PJySOpYUcD
B4Y52qI7zRDRivLNm6x1Q7lj+yp6qRU/Vn99QqCAKHicZ2mSnTw8neOyoddxsQA6Tv6Ww34nu7Ke
Ay5HlKOBxkaGobUw75BHvorzWjazmlPGjNQNMr4Tm5eEc2/Fp/CbSHqd8JDae+NG0q14JD+onKX2
QPLvwFOyFoDe4duCwoZEDotfKtTS/q2p2qM4xJ2yB/z7NwAKW6lsJZ60tfl5eMdJk7QoLf/7pA7z
iG5XYwA36IWkkTtQ+dfS9RtoAe0Y2s29E9+3S1YOpoEX3AuDoyqOUdiNdWaiSxtS2VKN1E6e1clI
40H+J2hTfmhBhsDNt/mUCqPHBJLW0OmeELmc8Njknyz6l/7OmynmT7LBfxfG4XBx5o3pto3SW0lX
LAzbk5TNLq3IDj7H3bTB4k17rWqquyE+8bC7h5PEET6vOm/WXkH9yimidaBDCftnMTOZRn6LtD/l
MavPqLjfjnkfb4bwakFOqgjoiFiG7HGKffcXkcqyZQAdMY+JYcl8uHLYBdHVoMvNfsQaqnquz/RH
uHZ8aAvUqk5c36PWq+q6lO7mjnvN78r2jkjnhXM/8lEb8BITBMigE4rRXyvUY2EtzGnBAExydLGK
/INvbhKXuTrH6+6ev+6GR8BKzw8buC7yE8VmoA5W7pfO6PNQIh5L6eu2FF8LVdDjkBfQGj/8y+UY
rPxlTwbO9vXqFZ4GIjOLEG+kBFNL+xYv5toh+sETOSESTjH9rTgwoO3HqVVU0Sj6r/vVFVsyWOq/
AmrgeHmRfBLKmHzQW0kJd3xLiaV85oac2wzWnR0XN3wUlHBbKmQuU7A0xs/ZtL9ASjzsygVXBqWy
RgaWbcN4rtN0Mx9WMd7iC9cyYBeiYAvvXfE5TXwEsSSQZzAAjfjmmsXk4KUBKlOFNluS9yJMFUV8
gsfnXla5ngpDXPM9IW6k0T06EmO5fdd0G0DEBRiEF2HCJRy9hhq4QnOpAsv5DWFPQa4bEP/6kz6Z
TzlUCRCAiYTJXRPgxgoEz0YKYuYfrAUr7TOusJMTEOmsbDJsM72ezEaaJmEm0HdXjgHUAHtaBCRL
wx30JjZSGEN3pbY06sUDjvrD57yqmS6Z432gn4Tk8OOmHhLdn2nVQw86rSR13QYrDLqnLitApm6Z
XhNeTSb//Cy1qsmQddp+abm6CfRjGjmf5yVrjaav0TAnyU1W3ZJwIoJrTaN4F+E6/tVfaUY0ttnw
IgIkDDvTca/oArPjbgZCVLrABAvcqBUVaUiMlZXSe6uoKERxRxfpZH13CR+Q5WFH+F4hu8yeMZ5r
RrYnn/TlkV7ncarvAkId6uAA/BMQbY9C0HHbr7xOvZRX5L/S5rmce/FhhxYD5f4IlmS1JuwlyzdB
vNO1CAtsMn70CPUu0nZIxJxdC8gG/jhhPgB3/fGE9yjfiZ0FFUuAe7CZb9TraWMimiqGIwZLmp5O
EGfjRUJw4/wXMJCjZHrij/73ZJtuO+EGwGjqCkrYwkVk5sOxy8hk3GhY23N7xUnHpskZwx35DRNh
mqE3pdm1zpVViU4irUJyLm3YnbLmSDZHKDkj/3USIO5JQuSwg0SzoybISl6RdAG0/mr8hSTuHZc/
eInDeXCe+Twkq3kV8GLGXqTMcYLThgJidi7F3MkQjkQB8Jy+fys2rAO/GoYvfyyz0wWtet5Ygj7o
4xXZ6PrGu8uluwrWVOuLtPFRACMpo6qfBCi/obspB3aRqPxzs7b3KH+nlnrpaqrBgV7hRQZ936ib
ORPY5z8li51vobvArp39YeHnbm1qQTq8UVBiAhk2xBOe35xI9DjIeryMG7rC33DdMsrxG1sMvl4m
8ZPrUCineqfF8MLfPThWyaypaPBGFLlXkt0sDlYQOj+0h+fwyTT9kwsSGd7kIRV6HfI91VM5PMnU
gkJf5iNM/ezKteKmG0SFkFRaiV0cRrRtvTjCjZRXj8qUXzbneHtwoKSqQd8Ll6ZwwuUAmUHPuUjJ
LQLT6AQRj0ZSSuD+8tTiDhRQehD25mNp0qfRTZiX1sRlyBV43S8POP20QYuzFwa7YAFY8CXmXGSr
d3jbbfxBOaNDUBoQHApH+j+hQ/EndlLb+i4A28ABZCQQI++c3+gv7i9GiSTtQoqlyTkDMA5ulIoQ
AOOA25ib6j8yspYGWM58hpZl50A/j4Z9myyp1ymNATqt2v5zxvXr2AcJ3RgRq4/jeKWMRFq8pJE2
afIwGXgDWaUoDRVUa41/KsN9xiTiQc9p5jA3eQG4GHXjtAaUiLJPf93tGbaH6DqdWDytRbCE3DTK
QL7HjLH8SvEyfwWe4txK4YpXZww4tB6vroGKfM03fK/e1n5hpRTi3LOML5hf60Eq/NVv+2l0EqGQ
i+s8GaKXBHci5201GuXpQjd9wJbmMk8rg5QoTgceOiSZsKXNjdid974wkoVTI82jvUOQ6TYiJs6V
VGmy13s0BjQiMU7yy/jfGU6u/PkbMDGFEDAnJVE+Z6mC79t+tTUV2+L56Lzgent8yY/OLKT2wmlH
SfBstiwBo7loqheE7NoLyod7f0FoaZhxzX2rznKQVIwTK4Cw4i/pwS1i6JANIaA0KuQopocX2h0Q
vkIEftPHBBewZogKSaqpHgepMtOcweKn2Ix6oHcOezuC9y05lgz76bVAsjLJqx/PC8J8edGUcve/
aJmp+0VerhrTKspe0LTEL+BU9wN6b4cdoCM0XvoE61k604g9J6J+G23u6iFyl4i512RPnkmKtiX6
yitWQ+lvV9DBOdbYH7/k/idTGcD8ENfGnVvV1k5l0fFp0b1PvqgzLEx20RiHEPHMGVdWFx1Ggur8
mMnSr9ba4Na4Fe2KPzJZUB8MLy2We968EGBpyMuI6WNxDkQdns75BnUCW4bThtwdk+u/QLGzo8RI
+NLBrecneoLVJU6VcFLYL1S6IajJ3PyQIVBN0mCTxZ6DOUo3OzdS46jY4mXg+KDwaInqDGu2nAMm
rj2/8/1CbDsEqYDiv59ODhSo23YwGQfRm2jmVJ30lmgIZmS3OxrQpLzS8cMJtOjBY/EGBD1JnSFY
HMJDA8S3urG0fvDl3Qxkddf/Uq4uN0Z45f5mFTrPe+Ho/n0jCGRKGRf1s/kWRkIwFvn8aR7s2Bp9
Zs6Cx1ckoge5QqDS8uDu+Fvbj4Nl7pHde97jiwbHhhwOePFr0YUetWcqMYYShh3pcY0c6qn2lK3M
oubdT60w3qPG9vXY12qILsOzeW+fBPPGz/P+SJOZUiB9LcV202Fu8qy3CnKveRrCT5YH8cAuFT05
d+gchfyANvdRFIbkLOk5BB9ec4fZlQ+5zaJJlufxpPbkXo/izgylCR5AwrTR2QxeyOUHPHxaaCcY
8fL/0M/GixOObvkkjo6ofXk9lmLwSIKvAuBkSr1+7X5DlGGKLN8twtTQ17QvjTSET+5RfLh38QEr
TcHrqZlgIl/jWaej0x9pApmN7x8lgmb1sUOdT6oCCLCQ2RrYINlNErHvlmUqgnoqXHwjj3BDnLea
5GV0Pa3wK4t13w2vklP+806of3L2Ly0TvgkZHdRI31ZP0TXouTIWz/9Am3ZkJTSXVcKVwytPsMOS
/M9h7vJEkGLZm1RwZ54Ehd7y+7MPEriFNhbDLWKtCzYKNv6w4nnH8c1j7D0h4CkDZF7xE842H2Rg
+XpEXe/VlapIcGzxJLBUhD4QQbQOxkGD82E47H8yHDCJZnRQcspYGqdBFi71hoL6fjpGY9GXRbYg
kPd3jISKZE9mhXlrWgam+bO7zxxS/qS+6iMHNWjZDs6ivqFzMCZoKbaxaPjB/B9yroqGy4klr0Y9
G5Ry9k1Dnse/ThMXuKV7GjqXF4DXLgfLy8hkvMpYZcxdyLdBjpQhq1zsOOV24Frwllpb+HBNn8hU
V+MrOOM2ZVcOEbuIp8a4/9NuV+hbQn+U7uP9880Pt4yQW1n9aXP8Rn8OM0LYvfNq+2DCyaseI2y0
TXdTiVNVKVXwierEpOl3JILlrfsNe+lnm48LjAuiU6aDWZOGCNHk+O+VJ2ekbiZMYFNdQXs55ly4
4CefO0nVJfI10nOKUHyIVcArk3BO7zM74hFlLbjBTm//Btdy4SnWKDza8S0cG3HMjzR0hE21joyv
IF9r6isoDfFUS9VbF2OWrVeTbDQjF6YIOadfYZyrkwC9tKgghqMc2EZModPT0dGMcZgM1ctG/acE
XLFFM8/mS9kea4LuMtJ6EqruMqpZIRW6KyVkspW1ju3ucWh25iG5QrS1ONRgECxHSjXvurJbQZqP
v9MGG4XWrFa5gDjdpB1FPTmEwT7eYfOzAPt0RvtyZVopxWHFcV0eOrgsSUFPyrxEO9eNJ4tUNakP
03zRyQ/yv0QyHJlVQjT+7dhatrNSOhy75Q4jTmteqcP8dx5nFYaelQUU0Omr3JtUVzA66XFIwIP/
EiTy0kGnvrIAyG2Zb0bLEv1RbASsJL2Q/jj3AWZPI6WzCSKqq+j8BhbDbKOfhJJwO8a+l0XLTReL
uXXkxnum9gs1i8yHP0qIhxg7qPjTJzcgKzyXlJ0sqETjn3xJQDx/JqvalhN8M19h7HaaTQmUGY/2
Sg3a9dnoAOly83wk6xv7Kg1aEfEyGaumz4A3XF+5kroFXPfh0yFCqUvh+H+zKLISucXlRVpRJMLz
H00QZd08cAqEe4WlRH7AYgvFRudWGnH2D2eTs/DyGolIOdLUGyfSXZz7YSXsKR7TBekPH0Pse0eM
pCdkpzlqZ7BMQrekqsDdawvBGnFgZxmY9Ac4Yrzah6iM0gw8EU22PCNQtnw1tJ+Mq398tSR5SvpZ
akhkIyvm4/0q9W/lXSj8XWJINV4rrtFEsu3w3I8JO8ct7O8jQZiFonFAwLRqHxmSk+Rm3G3jpcj2
UpJ3Ld3Uyklgav8KvjuoU7GUrZKG3kwAQRPIpviLuixSiFw5EMF77tXMYa4E3Yj+EI1+vmzI4ga6
zh2+OCQ0ppfBFz4DxB/KPndCzd3bxLND3sBpQnIFqltDwPAqHlBKtHq4qhjj4EIpvvdZOo0u/lNX
GuEBjADWRf1ZT6zjMRcLCQdE744IxB4StUGPIl7HX99qO797qdKa6CQhOqyW+QwM2K0lDGoaSnKe
lDyhTzXIvJK6GTrQvTw8FKkxXavEPLN/e8j8uBchMSqLSJiVanJV8O47Kt3Wv41mChlF8kpTimLb
rd0n663LszBNbzhAAaHsCMBMmQnG7LmNfhECCCABvDQwJP5UYgIdcsp4sRTbnep8UVMnvsBFcAQ3
E4ldoqqjxbdzY4B2wNf/vBU0uqQhQkG8TKQfCbE7oNyvV5zlHJZCa1tgtE4KoFhZ4mddkvcha2U9
6djuEGPYKSR4xMVsi9kX1aVJn6P9lapqp159JhHmy9T3OkUw8oFA5JT+W3IxzSW0JP9CISVzvzW9
fmhVQaaN4vUqzFM88mUSiDGsEuv2jpswwSxjkFrxouuSD/o0AynJiOjCZP4riD2jJOS+Vb0JjzXE
CDdcGONgcisOG2p0h2phc4lMwPnhWKwaw+SAGRVBG1OVrhXjve7WUOyVt0pLJqeAi3EcgrFUtH74
YTLipCZaEAx5v16N99razxRg1slj4Frqmj0cXhcjX2iODsP35u5poW/bPbcvOajv3+tRcf9f0k9h
g+nJao1E2ekawfrQcNhBcZK+wbf6qy+0zwsLUWaoq3ccJmw8+u9MCOOuuou7HpV7N3IhWmYDtsiS
mWFQJm4DRho5lgIfAAOoAEWU/7f6gkG3nm7lGt5AKWVXjH1H6u38oAOuDPVluWHAX1aW2aUhKUtz
c7ok7zR9E+OtiuLsBIJvKJ+wLOGP3MLMfz+nWgbQylvOhZ2C9UYxcOb3w1nLVXrroOvXIKQ2AViY
RBcr6fkjMxsXLv4gtcZ5L5dZJnfpk51CpBmlpA+WFrUx87ijK62Loq+K9/NSjL01S1B983GmpO3E
/jfyZEpgKf26SUMhn9ulS9OhmSJBB3EZVcTcmhj7NQ27/CNE9CNm3rxaalZX7Ou74vUuF3xgwBAS
C5kFCa0zCSf6Z5fyBfoT56MgcmMWQHL6XGen2UGx7pN1wW+2MiruXrC0p+lcDQoVlZfVLNfGp73p
TYOA13o4Lz+Jd2nQy9c3wbzAnOZZS4Z9jZCrfOvl3orX6s2LZCt0XYftMSQeZ88Lzjd/wNue+UBr
pv//ZFx5MuJJnxLvHfYPsMp9VqYCt90oqW8k5r100akoEE4zYZyxg4ck8XiQBPQodV7JlFKlA3Nm
aypWaC10RZGz9/mUnJ4AcvF8p4bIXwELzWXj8jg7Ywc9V8ZG+elpy9T+3/qttFwi3UgokYjBXd4C
Ccrv3WavGdaO4I3HCZS5DnofpOBZI/6raaaFR2jfDBqPhJJ75cuA7XOAjux+dJ4mYDVwaEGNXacf
e31IObiyoOHYp7TXkgV1HKGV+09vZYEOG89ESRH9WgFt05l4Lzz7xnjQ5fNYlQqZcd/e9shMUKLd
7XGovjPVtde0AeJLxOZrGTkbQ4Xv+mWk/54vz17+rO1m0QSjXvR2J+q2fXhr2x8T6BfKwXNCwnUa
wCgJxr9Z5Vb6Q1F1JdC2wDShWJGbYqOg5Uu2ki6uCMx/sIhc0w12blz2iiygL7+tj8NfCHmbMa8E
xPPAOczdRp0gONyxB5spN/4Flb+XDXPOAzn3k3aKJ+8+/Dm62UD5nJDpKX2cDTmuWoZoR/y550Uu
R05o1xX1+b/EvabUPh8MQPJ+JGc0IEBIZhtuaZ6AYjQoLNXvJVTeYjkrtRfRfz05TDXKI59VKLuH
uXz6o7ZYFNlGtiARLJ1mGUtsk6GVrO1EACTpcCc7DRI/GKivYMACOuZwTSSusIe9cunMjJqY6BVh
nJ0SdODTQ6KmLhiag5JHTrXBxHXc7K+bDE0IvY0YQSraDZx90NcpHV/3n/kL447fhVObKiIEM/YB
eq2TU9F3Qqc3cu/lhe+43EyjFqUIo5XD41Kb3qaX60CZsbI05+2gcEYh4j4TfNx4aarNeCsVIHvx
Lu7OrL2Esaz0ye0Kw9psxaXDoKouoEOCEHLlJXzFs/scgPYDdodrSrqbqgJJSKOuhCOV8ANsugcG
weLcLy142sSKv0rGwyK/x7LROj4Nrkfol67rennAivXcZ5bR8B+IQ8TffSlV+l50BdmmER4FC7uU
2w9teDlpZizUwMiWDuO42PwmcPNtLf0YZDjzkKb/R1B0TaSjdlWaeAXjuy92mFtKpvt8RC43Aml1
Y+nrQr0WWtc1x99k3Bes7dDBPfuctCzmSvQnGBfnjD3iMLvYvKNGGuMJtqRBwMcJxypOX5XwUKRt
VVVkGLhP9DVTx065Q86u7wmuQkxwFps0pZXMUYSxgnEEXofiEPdegWrrngLd7ck3mopnVU/fPUq+
jhhNNxTY3kJ2XEpzFGtzxCIkFjOenvodxjYtQhZvaWPH5SnbmewdKonZxmRGioEfkbmrT193oT7x
8PSsescdEIVTs7rjx5OJZlNu8u/a937ROTiO75G+6dOzxocxa304KUnqt5zqF9i1+kbstsWYWKfY
NYJ2jDM7+w0a1u5lJab0AJr7fQWCOJjBAizEn3s2S5AS9lxi6S3Yrc/MlN+b6utX4pvN+4Dmp/9a
VC68XJ6BeiJYeC0e50WHR1vk5VbeK/HYrI6stMsX5rCg2nuCZcs7kbWniwGmF5+8sTgSl8uT02n0
/FBlh/BJEIsxe9rGdkTIYtvhVoLIpVDqjqz441uXH0uHzcpOov76M+Tn59CGrHL0p56zT/FlH64d
QsIgGrvSoh3qTKkD+mhRZfpCzsKP+UpZMkLmsi9wRLj3L1Dg6ZSS5wXdxBB/1qqa3nPSvLeghG4J
tA4tX9t6RphiI2mrPSDJaaOQbieL+NxdwhFDVhlzy/7lCxlyf6ljuuXF2gSsGuWE3zGYOyeT0uS/
xGVvhiSAZQoW8Q4tFujPRi6HUvxr8zV4TnxOjGNXewnjY0NdIQ90gRpA51WnFzIm3Y3NqaJVkGeU
wGCkyqtVqE6n3770R/+6kYTArOamSFM3xzGBorkBGUweo2qkz/AF4T06fLIKdgzj8wAw1/wMoQcj
M37DOc/4thuvYsKtChzkpemwRT1/wupbjlAsAqpJ6sZX5poPJQ/uOuh0QZ+07m9gz/ftsOFNoqgR
eXx/NSsxaJfoEEwCRxBjDMCdx1Cmkp/5ZZ4DLJIR3piOq5f1f7E8U8S/FXOcO5ccFL6gZpHaXkR1
vSXSchO8Es3Tkgcl1c6/6QceQ+knWkp6/jeuFjj0RVZ0gX8aShJFoKJmYBxGlXNjD+YnqDR7byT5
4Fa2Ji7geED+MVuYjaboWpBydV+BZuxQ0x+GC8SKbJORwsERI9GyxjMXj48/vsBqPUIJ618nAEgC
NEcu5+JxPRcPXYlRafHv85kJ5XYcmZ1vGyaTUlw6EJHYRFFljBRsLrBRBQ5BNm6b/Fc9u/UVUa8E
+tRDo7kgmkS6XLLUQmzh4BmN2Enz6ISJ6dUoPa1iXz9+uzzn84N4dFHRIzSRB73czMbe//OL7N5z
P7hO/4b6sx2CSXxA0jSmXjWpWCUHtBHBOkln2yVnhUC4VrIGLkbZP/Q5N400XhP618DBmzzW/2Hg
ssO4Plhocvzap76cb2fx6IW3Y9u4QBhBx7FnOaLn8a6bgADfkocHZVPja/XosLMFU/pCXko2CqAN
kCs7jBbcg189bd5PDvoZVQ+XNfdTVW/U+JrwmVT4YB8IkHJOTRX7b2Q6RXh+ihJNIUyl2WNwenO6
z9ytKE5ETG1yrRhmCc/GosPB+N1cMES6JQ6cbVsbNYyDrLTZsgukoGLtXa0UmvTf0EI/aSEzMx1s
h9PKV2GqSa1hgeH6Yhywwu/f2KqXMjFrGf526U9PAKeVM8LhF5CKXHufgFDZcQj4K66b2P+SLcpl
9TdVCkERoovgMzcBaTmho3Kcb9aiyISLuESXMh7KcrIKCeMLIlxwISArb8tzaoTTgIjLrmyz6w4V
ZTMEOqMiP9Ff3b9RnD4c5e61yDVMHL/8qdSDFj/kQje5N4Yy6JwDVoWNhpfgyH13yVR1IXOeOhWx
o9IeW/kpw+qiW8iI7QztZP0etWT0k0p3qqv54JyI8E2mliJcg+2KRsmY4Hp0d62tlDHXTVXmt0Qf
d7Yf8EHoOlkVnr4ZxH3zLMm/FQrj1TYBSZU5vqniNSUrCsE4/L82jOBu9Taw6erLk3I5Mxol8yR7
UHNlrPGbKIeVwbvyypZVCUtpZMTFxp6X87NWKhDrLf5+rlItYbyxWxOm9V6aQHeD20mhjWvm9Hm8
33Qwuw2ZGvvG/xlT1qPbdNrVlPrp1mbwhN27rPTYnwKE4bU4SZu7fnuGEEnTEsIalNQOVIOMm2YU
2oijqf2Jzy4kHBw9+It/LsdI5qb+PgB4llNkBMakSu6YPxkej3whl4b6EKDktpoy37GNjmuUFtzJ
D0FIzHO8n30b2PV1L/wgGsygtutQe/9VIlL2Ocyj2iQ5Z8na69YgNMX0SXNf1zbbwsF5UIKEM+Sn
IDHzgxE42tENORyDsaAuJNDukzg9F7l1t0z9A2hioaTF8B0VjcdBk7FEAx8ZIwktSlzl1NIZQyEL
N7qA6nApv6K2ZDbDxHZ/WA8ZZFDuyQGtwlmPGKPpvnm2GF8HMKwJ8amUsZdtoy3aNSYryDBRinVq
PEodukV6ZA4jH0RB4L9/I+T6TPvhoO3ZTGmbrcLwqGcYkGUE+/juM0E+lA4m+7UAYjeucnVSFBhz
+Z4AK6dILJR3Tl/QBeN5Tg2WtGGLFmMcUsXCdkcDZBquWMdCdAPRfBOwAWzw6M8+hscCh37MNFd3
vth0lJEPqg9I1DUmYzHVpyawKPoacfwbV1GsVueeNfHcbeotHiNZzqD0/9PUVsE2j2VfWe9x7A+k
bV9rwpyJ3bRKqLdiHTGgoVSjcFy4BvPuxRmFjG0vWGmDEY/rzzTirmi+u+44GPf3qJ7p9cFoxVUp
sDY9pxw1X7SpZNyREXjo8Uhsh6bWDyUYxanpQOfgNHCtAGnh/69AS1tV1XXraQbsJhhM7QBx6ZA/
1G7byYhMfBAqKHE6HLilMtysCkvyDP88FVXBTTN4WDjvVgcGm/6JROIgkyjjCWIW/nn0YxVOdaE2
ED/iQ3V8iW5RPFuRDIgpSzWorSXUV7gXDC7jePW29pUO77IdePE8068jQa1Fp4RcNBaD2jFMGfHt
2y6lue1+02e1IyYsBdhnpceBvWU6NfPPJJy44cBPz80fkbb51gWSj+t56kHOW2bVcTwUWUW6AM00
immMAZr8zdalDvhIQp/rr+76uOjvI00oXAFI5Q/7BoWEYJY9drjDTc28mM8P/3+FJP5hMfvW56oo
NTjipXk0yv7uVsA5OXWeNGdiQNUZwkzeaVieRvbQEk5HwTaXQZOKzbcr42mqq9jdRhjwrN4zMVHU
z/H5jycmbFirwreUqMIpBfd3NnhKdbN8Lsv+ZGHGdiIurlYS5KP1lH5Yb59edUILeNh4JNSTl98k
QesB/vK/lxKCcOit6skZACqW32Yhm+zP28e6LopGfHB03czoMvze3xWfFZLDc6DSdjDzgMWrhqqk
xNBr1Awxtz6BPZcGOioXZUputls3tH2SIFh4i7U4P0q3Q1ngJtcOTxMGet56pay/z0+syz/ElhCT
Pr/sKVkupUGlRAi2CnX5NbVNgn/8wVqWK3uBxtxR9FdegiOACNY08PUZ8h/z3aaHD4PcvOetufMC
tXS+vHKRhKkWqV4uadOMeYogJfzGPYHYCgnK9xbsVdvSkIAth87hTKVRT03ikWjuflMuTylslWqf
pH83goYcGirU2tk37k7udvacM7sXmuEfBgr4xcD3T91nYFtk/z0gitTfq6Kva7p9K/wZv9JNffgc
ummzzU5HLIdXRFPgPMp7EtfIzJllxmQaDC89Wg5UCxp+8YijuqDhqqsD1bun7u7lFlAGvUejZNbs
epSIH3Mcb5zAYUkhnl4B/Qbkbyu8DkgixO1XhdcT+wSgJ3qywcm5iW1LJb1kVc8uRewNdEv3wN0j
bcotGmESa5gaGCmKHReoG0ULJiB5OuUcz+NnValx/ZVMsb2kWh8Af1Y6RwBbBPRhTQugVb8eZrbP
2qhnPMRzJRv1lKBROx4GRhfDiCo1p6XJcLuS2zAy/KUxd04sl5ts24HVZQZIA4KkMFtFMyR6sqMW
9Ndz/Gm8WKL7/MJiIoO5awMV9gYMILoTqpVUFUh6bmNSqXULPrScLQZv/yEgoHm+lxexkFiRyKQF
AXgX/tWUN2WEuQHgzHG7lyphIvu29mNvUOZJw+NH7roo+45Y7wK+hXqEAiWCyxpmU8pGAie6fWXO
ASbHnn0KAqlrn0zhgGAz5C8I3BZ9dJzpxaN+0PMW7T29yRJqA5HnXle08cSklUgkEhi79G4vmq6h
V1OBqyVloh+IQ+XNHdiC1MUZdXYcMKomD7RlWiWWSkkBHxBkHyP4esdNXi/4fnsYqNGDa6PBc4xf
aFfAnE7E1AvUqxnACPv6ZSgQ48tWV/ROsf2jnkt4sEh5KfFBCEbp/Gx+E6aq6IMHHtTjAuCwJACO
aMcowQ+ZbtjgVc18BfOvM+0B6UAJltpdiaCNoiSGbhYzHufpGuuoB8EoEg0jY2q/lapaoQbmLGjF
GrfZl53IbQ1x4IVO8RK9BvtJDIkYIH0RulE0qO1hewyx/IDEPtJlZZfWL9yWI/L7Up/u/BJ5nfBW
eomX4OxnwhYrFOWm1RJDl2XIj931H3GH5xFNN0WPs1vtGKHlW0eB9t4kG2sH8a7zOyr9OaC+eu/p
VBQFGkBqrPQFZoU6jzG5BylNWylDOky6Djv2Ro5apMkiCnuGqrM465eSW173EA2z0bhbGdpFsS3t
lIcd4mIyjQa4QRvoHlArAgOFDlOUZsfiwq3Km/7fIwzyFbErcfkm5SgmLwDSLh3J7kHwtT7uQyjY
shglMiAcCv30qjD2NQ/se3uaHetd+LfY+vUTYaCh6OEIFPrSnFqJouz9Re7mFZt2ekepthBNQSgR
6aCmnONWQZ5fyKlOmhLPeKvF1wdXNwrKFPjHYd/JVXRjfTLFBreFNf9lBx1PWx8FP7cQQVE1Hv4e
RAyjoMDLkLl0eZTGAz+RlGWojHIPFJBdhpH+gzr2aeWrZ0vt3ajWv9dBLNNLh1k4LFLNaTlN0S0H
bItiNZJdleZCw4B5Iw17oSsaG4I0Qx9zneunwAaOmGdXXkd6uMlMG+Yv+vdLT5TnD8uU06BvlQJy
dvi513o+5aiY+T3nA8/oGFZxdH56GPiWjsW1pXyQaiWIGhrSj8nDwhwmAzKuk/xGwP3MwmaL2nhC
GSx+sTx6jZ4LHL+FRgMPercOqOu53S1QOPFaxzXWNZOnF4cHMC0o/xdiQRv/x+NNQ3BOBgW9pYsK
Z0iQK/W6S4A89615jAQ6CgqxDV1KMwimbuy3E/JsxiGrc/LDTwlPvyIcnS9VZOb5vg7e2qscNBCy
91ax7ZfRDXcnD6CRw2grdTU/aulVN1NEfu2B147NTqW02hbXkZVrTI6RPKyzR5Myi64pL3wkAbvu
7EPq1glmhPeiMH1jr/uFHh68X11otr3n25ut7KlXBn0fTbTiE/oZ/wLfWTTFYCA5lAH9/lK/0ex9
iR5BQW8KReN9WOt4eKbKWjYO/x7E20A4TZlFVsZVlO/B7Au0nUG/s19f7lC3MWYBoeiQrUdYpwAU
4xkbVZfn1ugaXpeg6N/rn2GidiCEsqy5SkcanNR2jUAM3hObJmuADp0yEhajWfp28+c3hU6ERazw
m1JABobnFF1E2hdBND7IKfooJrznO/ZnJswFOuzh+zheGA0REJQUoe5rpykQs+bZuB2yJhGhwy/0
jxdgS9nf0uEHaocx3Z+Ww2+bPO4bIk7VJn15Vt1/CcAbgnCH6Q2Wi+oJ9d0mlNdeCFfgCeja3gBj
dVEnIfGW2YsD4DyG+6eQmEqmealWBf8OC3ai+fk8+u59tRykKv60yolVGegoeCAsP4KoY+B9Zzio
Bu1eKnZLF7VcR1+DUiR/5lUalxpla7nmy1c533o+2fpKClHVhccwXMBEM8r3j23Tpi5GRvFK58GY
Y3qI1mGSob3eqvDsrL2n81bP7IpUhpJBRA64VXS5bCTg3MoFoO6i86IJ4Tg6yUBIrMkDAr109Cg2
Zo2hqwRletPMlPAZPcYr7V0Rfoch+CDF2FKEG+fQF0s96T1YrJBW/iFWbzu1/4ao23H2u/jgAVB0
kKEPoKNUPiPhh7wJM7s4hemWC4JA4cCORESEwhqdkWp4uJBFXDV8gR31sbN5bodoV8CwwhaCZ9gK
u1c8Y0l8MKOYTu3Q6fmVrd3PmzlwTbpNVFvt2k5lck8ky7LbfXxPtjtGflcqwaYIbb3peY6QHAlR
cjy5fiDJNXUxWEEQpKQJYmATAzEabE9bAGEs6dAEicekdnDrNXVr7yzKwrI5eCfcc/ieDae9kCZV
gLVueSfH8ekrIkc4wp+OHGFUgv3G8JhE3roQfJ8M+5w1ZjvPjVUMKRUM4WkfwxPgVYhSj7HdUePt
rV5oasU7GywblLqcdRBbasGrKR8p2NkNC9Ys9+IkSFKRZWfyfQjO1lcgNk8lbWPwFInPCBoLwCM2
PgNwPg8u7jPhWBtBtYB1kNTu3eYE+MmycpneMD9/w9LuFCyMAUB0Hvc7RHLfTTWi3/KtEXhbI919
RjfOuOocp/NV9UYgSooxFeCg/6EG3ZQs22BMXZgXSoQq4KkxdnaXjZcXfZ5CQQGuDze3rygdeFY6
Mo6fEwf4p0xZhmrHn9ZL2YqV5iZE4qwGSaBaDMzafQNoAq7zceQo5xvVjyZ3Lt4Jq23CufsIYf0Y
CsInbfVynid9+gRM62t8tcxCsNKLX9up+JRI/rVqUB1PZ2pjK6LowY9aFNcHX62Rys7FMmW53pXR
S4TuGvuwaWW+ZjYpR41NIMvVmtU8Et77dhvuyTmRR4fmCZkXLNzI+d753o0I9NvJ5yuMoCY0oW+6
7PfUWBXeBi2mz8RTv4UbzqXEJJVJumsbavVJQk5e4bTLX6s6FHz26wB9AU6wPHNm9h1BSk73Jdz7
rWlRGwm9EJfgwWS0uyfKV97jvmgTpL7a/4q7odOOpraMP6TgixBIQNvyeVY4Xay8VxRdhYnRgkhz
y+EMSC4cMDMZsl7oW50/FgtTDCkQwHF09E72sCULYpgAGFpPEyw9oUmH4Ss41iit9tN4/LJMykD5
vlxDqvPrXr6RpaeR8ZfC7mcP+1SnyrzOQkeceJvsQoQqXfnbD1YMD31h5mbzbM5PgzsHm9A/0Gu4
lodow1IXydJgldoxcL0qmqRF/PoYgYq02khk6ao0jdE8E+m18FH9l8aCE6b7mMZRoUrEmbA/83VN
b4MK/3Vl9WCGG19S8sXhq3IH5W+vxRcV19gcnN8DSmZJ/rgZYHrbt2zuRvHTh7TMXvkBZ1o+FnB6
jE95CT7OQlpUVvmbmLWJXta7Eqi8fnPSnAz77ef863C/Bm2CtAUz0ewCI8opGDXHy7dgTMfXE2TS
pCg+nHuBvWb54KzHUiiGktjC25ygoz6EM1gmIuE44YJgwf2qYuK+KosVqMYwiklBFQ/vhPJQEABN
K5VRzb/xBYBqPmMoRY0XPewRumanJeJqL200ntv6bUrsU6f3poF2gk27daEcbZu/c25skWK+o07V
0IFgjL6eiebCtGGafmqnvEJrDM7sAdkyUQoNKvnOzFlAADe2ea/9Ea2ovn3HR+ndnh2q2nJfVnMu
YtvgIEgDM7qmWChJABZed4cKB2sXFvusYc3BcXjYYnqhbXrpPSRyQm/psLBC9Zd0In7E1kbuf1Lv
oAtpb1qKGsgqa3dgE+ffebEWQWG8ZotWTWwai8+WwtR2e63Ekq8+Tywd8qsNwHEqLoIemTRPtXNb
vbiMD7I6fjVc6wD99adGb/j/sQSCUytbK+9QlTIvZtbgfOdUnwkFTbzd1P4BpVGAkvSBxXEfrL5s
J7tZ7BSoxBmFFkKuwqUYR16sYuTLaS0xNitJCFkS46wb7E00qQou29MVaLW2HmBx+QO67E6P7GiT
p7dPOTVnHrI4pQHGIhC0H+mSQF2/G66IARf4VKhe7IYU64jTk8BUslVzozCWik/gq4L/LUgalIvv
cXSFuwkwdixD7uLTh5U1fR+oyBpAMkmsbs9k61IVUx2u90S+xb0s3vhozn1dcksvc/ca/kjbxYea
4MsNztW9XqA8HNE489089JVNHkBTIFbdQlfbuQJOd7k3THyPLkYalkbNq5oR3aXQyOhswkLD7kTZ
5RAnEVqS/7j//qKT0em4eLfAD96XtRuVgPIj9PcZmVzog8mxNppE2/dy/z6W6HV6RjJ8OucUxIDh
mnEqSPeWkYX5oD8WVsVG0ednBLEYkEAZuXdaQ5FKwummjMAl90/yqvBe/hkAe97pXoEw2qZrxbjx
Xrcs5PH7fRP9VPiVmTxrBWIgIO2a0CIYYbKqP6UISgMESdJSsBF1RkjpM7qM7Z32deiXOJi1JffZ
vsVivYoOGgAGZ5GpYU3rhCCYwyh6Ih6yjqPlfWXDWsUq0In6leM4EZuIPPlad68YSQWY9Q0WAcJ2
/x2jRVpoEetiOflcAvfv4xDBPJ0oTjJTz7zcrGJHp/gnK58J+kzjokdw+XoistNW7KvW03scDGzn
/06Oz7/wgnkoc3I7+gmxDiygpIJ50AvuosTdnQot+M3Umt6AVHpD07+EdZyb/Qqf8RKnrb6QGgqs
sJ044J5aFp0kvrcIKF6B+urRi/jJ8OO+yEYb0HbJiXXACCtkTvYLeoRpsg/4q5Td4R+QZ3eHCBGi
JOw5XG8d9AecFl1uUbdwfr3HV5D49XKJ7owV1hOkv1XV3q51tnkWKxuqrdqkF/hU4A5LgBwHuz4b
OaOAOrXy7/RWYBt6rL4gfG3PS80iIrJpK8EOa1/soDpkIH8bPXPGK0hy2/I0IEEIWcwIbko/upZP
mGIbkm+m+dsmqdrqO+FVpXTaMJggHH0tEb3LypcUSrdM+zApvUlxA9ScqD+FFnUrZxYdI2xjEFko
6RG2xwjSvsL/JjWmwPY4LUhmM/qJY7Cm6aySPFhaB439b2tBVKlBfYacOg0ZMvKQr8J0dlUeTYCp
HMiU0Lb31J/ogWk+6hgP5GdhZcez0Ao39N/dkKBc6a1hJyUb+hNc8Wf/nc6ZFwAPlRB2nY8y2m6E
/GN68VkOoNGyuytdLP6g9ZB0mYeDwpl4gInSVnBy9Cps/07+GDm0ZnDv7TX1tSxqqnCYeHJfBLud
ar080tcSpk6mV4jSyTuHsLJVpmOCPtSK+HGN1cKiZ5nTAM4kk5THvwHnNP7tP/R6rwO2UEFcFGgG
EQWjgHVx++S5HyCcc2G7zRJgdXoDq+Ohdzn3BgENlwIcrUQAVi9KNdZ+UrQ04Xg1KSvCOXYCJFVa
fRZUY1Ci2Ea7ctuxOmILxOt5q2oOnOjgWmFCJlwAPG9LhrxhW4lLLqcFIudFrozFpVBdC+fhI5ng
QbgQaNmCgUlvazqOMiXu9j299aqp+hVsTZhw9/E+PjfHTfvlsBePLzWfumD7haVBIUwkLq2G4S0g
4hLX/LevQtBIDi12JgdyReviKBJ8i38UMFqQu1E+J9iExXD9p1QjlgSK4O1W0lCigAmDweeHVFM6
qUbOBY2ALsxQRAyhkB6br5FYOhiMkWc5ddwMS08mwnnJIEb2cmDqtpxip9WwE33ZklN2fFwvWbe0
B55ZtPy6cYqKdzpqjwYhI7CCeFcdQ5m4XrPioYGQTf+ODL4GqzykoFANnLRFu/zOgKA8noqMCYKD
pTLSlJBbkIUym7n62CM6z5HpWEFib9ZoKdXy7ERdmYNHuqY9AdCE2dUjAQUYEGFsQ5qliOacVJiw
HYsvW7ZOmSPobpUrVbIf0s1BY7i4XQaBi7BkJSoiy0K2Aahe647wf/Wjbbph+gvUKCyvZe+fzagR
6OI4BtqH3zLRmPR5YjO29HoP+CB7X46WPGkcpkN8uJz4tK3CdZhciF6Xm20xL4QXakSIIHqX4y9X
oRA1pBkWND5YCS4CPi5Q1z/jM4dCJN5mQ1wltqMuoTxs39K4srpXXu4gy3wqAu0hGWRNyUCVD1UQ
XmMmGuT0w42BaD0CIMdBLD3JPcrxZfwkF4po4+22FVgmF4sTT7g0/wlUYjIW+F2RleCH+5IFoma3
yoXU29OicGXXvJQ05oaBlgMKPD1tUWC4JMpLFsWOFW1D51iH37ieBdWem0rfuWqHdYlVIcGKn76Y
Tsss+WpKhBRHYanehE3FH4HhRAOjiCbys6/e7rxP0fBzMd1eAqau8ThgMMaXb+9tgiGAgjHt15V5
gOKzzVRYbp80jbzYkz+zKawdE7sem2RfOBi8EYjpABIBxc3mr9HTxO0zHtYA8DJveoerGiOV+6nw
rjzxJCQ1aDV9/ZOavGZeWpbris65SuivIBPgxd1V8VL479m39iuVLFMB5lV8yHUjqNLKMtDCrYZ2
TWN6uf9zffJu3CovcytY/LSDDBJNXBiYxUmeXP3YRGcGfR1HBx7c0xjCjeM9bLlNKJ0llC4enkQ0
/z7F/SX/GyHZ8Dy+4txyEMATbWbIpG4taIw1v12Le0FCeCyPRqVSbGtoQTXDzrdX289tYfxQZNvl
n9bfxnP/OsyV6sYCOjUe6/iH5EnpkMHFA8IRBTAnn0R5np9thZVFC18OtEd6Km3aNoImcNUPlI57
JqvbafG5efJ0yJi2CDNcyzS/+UdwsF+KiAqmJWzysenYp5Ozy2paAf/woXR3b0mbULHlTQIBClII
a/GTqavgodeG8q0LqBy79fJFPLygeO0UfxzsmGccD0F6KU6TDNDQrZx9gfwx5bdqLLGn6rs9JlcD
OiPKILa8OQ270QxiGZ+Tq+BMRbMI+nRvXhy4QagWybcxpO4frxi04OXEhAdvMog6hmDMnBVa4uk2
os63Bq+hvbtPkH9gWkPOB4aAh6uZPfV/QIvmkYC7H8WGk99XsFF6jaxUtuwZKU3eKwbnX4g/xZ5A
5ApDeyCFQTf08YfZ4vzM+E9atWA3psbSxl8OwYF7UyyysthpET563z4uhXHENh0M6/Gd2blLtetV
gJKyq3350WxE83zN51ZiEFbwlJZhkLHabmIH2tzfp3IPMOKTRqtp9CWpn5Pb37xqyoYQu4nIYvOy
pvhFS4Z5BDFEhWSMQiLrHmgleXcU/wka7AfT5iPNuHshjuG7dZo4Upo6DXjIIvt28EmD0FV+AEQR
L01O7KGc7SnK28izEMxJUBrQRLV+aslmkzSmS5dMeKhiG9shTnwo+PET31hCfl1pVB+2Cb3/ISpG
mDsrvRPaZR0ha9BXPcDvuqoDtrhNEwyGGRc57Wy0g8Ynql1in6l5ZF8b2W5LuSsipta4892HC+ya
fda7qzM+EZ9zybxeskgfOjtwSnqOW0ECYuqyi4kntyJVbumG72ASY4YoCGMrZ2hbBR2NqgNLolyU
10rH4UaZogH77xJ/e6ZmHvBonf2w01gUjRDNxOmXi37k73i8GMxcNrXPYprm+jOZSHudP78Ejn+7
TTuSSxWSsMRFpKZWOPX/n02hTaJ/mpbpbuETTngc6lvAax8I4UbiulYaojsIZeTdDoDlfBzc6kTa
yYZJJ5lpmQ5nVBOc+tPQgOdzG02xecVU59HWAWaXBSP+MBMXyr+j3vukiG9VTzDk7WmjwVsfeDR4
YIkMGQrE1fgzQbZe3R7Fp+AEmK/WFB9odk2ATmyPDmK7jrrFp9neppgoOctcomoqKxCEywapexyk
BBq9I3UZ8u3cFgA0rSrHmw2rD57/q2BVovfW9DvqKPranswq+8lnkjGu6smHqBQnilvbQYN0bx60
cuJWnSdaqnT6uvNfjnoDPgPqVV0NAVMT27t6v7w4C2n5//sb/q2hFroDElxiJUbv3Eo4Vdjfk6fb
l9FmaPGZ1Q+XInCPzoGN4BS0deMVC2MNwLoNiwUz/Yrdpv0h/eRLkqZMqLMYp+kxMDFkJ7exjJck
0QPTIpeBHy8L5pWroyPf6vGXVLbxchi39G7CPMYme2BujK9m5XSXfgb3cln2OeJV9trh7OMKJX1T
Mhsw3mwrdW+kQO3OIaEpJAcODpm4xHXiSdb1pj2clA3JPytcq0rJadhMhjrLJfUULq/ne4e8uRj+
kmcOxdu+kYdc1P7S0blqiZO+yJTnS4A3oEdDI4TrJmfOWsuDoh+KN02KrmSPP/T7bffVxI0wmQMj
PLMYuZE0vTekp+Y8pXq6rydiOHmaAiUvOeaJn4JI9lbJx52cB3r6I8GsEpAs8ANA9HzpBoPzEgeq
SsjT3ZY31vjNZk2xf81awwVEO8CmQ6PRDC2YjZZZc/WbkHLo8wxykRNDc6cWYPLTIcopX9OVeCW0
iHqqimZLC2z5GgqDS+k5UbKIqw1twsLAmWM8H4muV0i1Ji7zZ+MZVXC+/dt4tUf/bwpQpHeFk0Gm
dIVxfr0yHqPkcfU5Bo/d0Ms1Pnv7YQvy36UqcM0mgahzCAGymuw3NsSHaKI+vyDZ75+t89WS/Uka
A8VZOo8YyooKaBztUcDNfPIadOKeyPh2kIrchN0ldHDldcETh953965VpOzQyh4mdDM6TBnxFYyw
D4R8iu7XHbt0YEVRuBxAyp1cGVzY+8MhQTzc0nRMmmH3qL6Q4aQXeub/8+C1Abwwz7QDCaGDEy86
va0Kf0qrJ2qnguQdWIig0x4yDjrbujKLQ6sBBFr0RXJf+UE3CP/QvbMYe+CGctE+ISYpguh8Z7W4
N3vhUliXmyrh+6+6SOemIcP+2/KARk+AoCnyDJ+5FcR47PWB2NgbdWWESn1q1VEumVJ+thNDSmU1
4KA5vDZzrmzN3C4lXzEpYymuVEo9PQ3ynlxhzV8rlRKav84iSCwGRqOVbgV943+JpsXcIN3u5+4I
g7e4gIEupzRO1FSTBgI1Cu1P825rLdmB2OzNQQF/LhSq3vxnp043h8zKzvUsmkT/lfdsaVECWDb8
oNu/jsd8uJ7SE3h9o4ILCk3n3156tFC3txS/6RZx9znZ+VyOzDApIr0w+FDvaNsPLfaWpz1xS/kw
02Dd4GUG8tWKCiVBOm+VrjWiratWPYjr8zo8oGHXBZNlX/fgz3LFQvbjO+/Z0lZ3idukWXCXuR11
tsmokP9Smxx0snCocEKRaZ/iM7g30MLdhLI2BIhThgcQrun3zSy6mjAQErjhMdWr7PntHDamdwDS
JOAWoPHx3PtICSe4CUP6lV6nSkeuEKUOyZHkct+u5XlLIC7WSQuy5SHZAnddaF0rsggq0aWiPUPa
IQFXubiiHS5xpTqz64tO8MwK1wScoLl33tcI8RG+JRDXx7c1HfD+gk8vFUKBoYLa4S7EqboxU7UU
L4oCwaaTEN6aHaz0u2cNfXLoBd8t1rMLirl+5S0+d694mC6PpmWumG2x86jnF/raJOEYbuyX4ws3
awjCLXy4qZAIPNGU4/sG5tQVdXZO8yaCI1nlwUZtPXfPXU7hyBr4DdND/pXsPzlq8MZczdvlpxrU
zjwTBfaygUwB99jSplLL0rrq4Eld8Ux71/0eA8YyVDRP9A4/o9PywTI1jrxe8jlZMiG1KxcrAQk+
dugCyJ3B3bplLLzJ/uQBN3czY3r4DQLmsVg3ST8E+wlGKtml40C66Q5QskRetaAvNSw84ly54+iW
rsRXwiAb1sNiAkVhyNqm9TE0mwBxce1V5hrBkaaUcnxncFMVs1UPsCikHH9/N8VMp7wvC5wOo3Kv
Xq3o2LJl92geA9biQ1nM0jnjtTC3A1IUjGOgtW4tNvyNt7a4JnVHSI05BXlzGjjEoSHOekD8iAUV
fT5KxuGJIPBbCaOCnAiM0SJzEiuVgIH4KMVnDuQHmYZ5tnNmNngejaFoMgT1GcydhNHD90PekqzD
Oy97RHFrKThDWHhQgjm+9/ezYk3fFKFrpXReMVomJTreplgT4g7kc35AC7hmMnTCrm8IVjuEOCCv
NITp/Q9mFw0v3+foZTEQG25UgMbLijS9iUrDwYPGyPx1YemYSVE/TIQLCcWznq2BPkKZXhZshr3/
OwrWv2XuVxvsy8QVFTF1sS1Uj3LYVnBXjeAH9Tl43N3DfG54Xz1VyofliEUG+xeZU9IQik3qiRHE
6OoKWVvTrTNOvdCik43AGT69CPU0DoCadFM7FupLmf26bM5BXCALQZOO8jnJGH3WSO6N/92z0mSR
aIWEUoaCtJRiIyxMASjNSfYo9+7KnQfRwTCGYc4IhQnWN954G4pEW72qStTXkLusCGOHJ+cS5fQY
R78otcVs6Cv6SeTurw2zb7NYplZU49LxvYJa9VLX7nYJO8Vx5bPWUpngdXnIM97lcVRVnZ0luSb1
4S+hkjYj1d7eDGgRpFyjLPBmfuRsXglX8ao1T3Djw2sWAZt1RAiNaaPjD9b2FQg/ao2XVzKGjPBP
hYgbJ7e/7rsI2u0ojHiFjAgZibOZm7ehFNrAaXXlpkBcaoa6hboWXe8V5+p5LsHDL4vHhmtz5XIc
TMLKSD/bn8QKVutX1aBswEY3LiJ74YEEVmUMDywLfKJHQaBK9a6qc2S9nxYc2PDZt77Xe/j7TmGy
tRTDTQ7ItJlfAU2Y5xgzO8R8o8VlEv5KI9mHwk3Naf08aRNYAVAL82cqEqtLf4BrWUThGwJWcekT
DOG0RgvJHhBH4+8l3nqX3Mdat36iUmpupK2WxL8fXgtQiLBGkvlUPG14Bea1c+TvC97mEb91hPq8
ThAMMRzx/UTj88jXmr7AiN8yx9qe4FFFji1R5IXIaVA3h6s8W0rd1EFUINnJNRvAucnY/KYr4aFV
yEdR/dYuiGetjFGA0eKdQkjHTG//YiJx33jpazfw4tF+hKsjJcH1x9JynGpq19N4+hn+cvq+pkba
46iS/tjkA/8HD99g9oMZAU7TFjGSr66mG3rTWDFj9zZczcGFDXYQDG/iuRCg3kUF/5fdzi809ayL
+YGwmVecGhV+ziY8cC77gAHlLtP1/YCsfzWXPp7Nhiy6+7wa13CQyD2VPnVwut23LG5ugTWa+ruf
fux9bgEIUNNUJqvG2xeKk8lfIIsZTahGi6RUi2Zu1e5FOIKQR9WQ3dBZ4uqPLgJ3k6TMZqKY25sh
ACP++qizZAA9SFrM4k2t6HYtul5DR1gwzn7FFyAXwvYbZOrufR4BoYqjU/cc8iWroq1kPDj7Nwue
dm8DkiUnHKT/mRpkQg2x1FvNDo1j81j8X9UCBl9UtY/mr/TK+a5atkAN++K8hS72ujuowlD5erb+
ziFQhYgW5L/ahwtb6RGx/mWEoMBGto6PYS335tdOv+6EaCRiJRzbLKu8cgJuQlC2rvQXU84nKQm5
1XKLfjBWYHhd7vj9WzGhu09OZNG3e+7C/KAVpoO/9Jhx4m5WOU3k58cs2LwSYnVFdg1jUFId8zIX
z5NxHz++Ci6QtRA9+QYL43XFNv/MfJZgpYj3nzqxirm8Hbd9iqLzWTAqyYFKIBuWOSgvpDBefD+c
fN2lwIS2SMZYHLQAJp6Xpmk2CJ2knPRpSgSu+yZJIqU+brsL4F9B+CLHsUt3N/E8BoFYl70s0xyk
bn4cmcWE2tIJ+VCRqC/220qOE/aikgTMLehqftBeKndwrwwaDlJMLTBniBLwLS/x2bIAmAzNNiQF
VbMBiLrhHaAhWAPGbtrE46fHkLifghp/02UdXpB+C4WWcL+iJooM6ZqvNtwTwF4O5aMeRCp7tmoA
izft17ewHxD7pKVi3zFir0gnQsm4p5T9SK656MY5/4NVyBaxTKTOBVBcpFf54dBKWUq3+Xw7dhvv
xAW1uxdOiMLxK3z5U/W2TAzXFl38GY8GkZ+OSb0iNxVARU9+G9VuMAzEwK+ArfsYNB2bQ8OETt1G
8/WfP9IF1vSpajT+pmMEKor3TUliKaLWnuorO0/Oo7RZ4pgRBUxkljF4w5fPv0yHdvUGIH5Ouhot
DWYrIS1+TuPk/FvJ2Lr7C6FC3T1DwelGnWdOXSX+TCY0qm9nf6oRqIWc4DC/I10yWQfmIXv0/ZKS
KWpU0Av22tSasxoc6NKq9ko+mLncSJW23plARHB0hGQzmeDPdDnsW6F8txuasQG+lfaqFt3z0iue
x2DGOalqdPW6GXkKJAhyHC8fHs6Rdun0RLonyt5n5OA9bo2hfV3IhGCRnFHTon8tGUlqkFEiYEPJ
M+WvmSrG9wdmh0mYtl3TeU6ZiZ8jeQa82zNqrHy7rEZZec47izfS29tUDVQHXDcN4Z2zyHRSiLOo
hmUxU1oZvIANxKGhIou+y12AMmhwzDUhBQUJfNDTThbvprVUIjCM8kvT64ozMkuJmrbaZZDKQSCl
zTciF4PNxCiDFwagy9+nmYeAArot4AwKC9/Y4jqDHrgMdf9yDcQf7+DHkBn++86zNgoHa38FBEzx
IeIOI/k0Mz7RJsZ7X8KzVfbiJyfB+Jb0wq9HBYhTE5UZNaDMD7Ed4sQQQRsxMb/YJbLLMRl13ZQa
GYc384JCnkCCqP+FYAj1VE3BdPpqm5QpRVYOQ+WnTg/h8P1rEYPkf7I2HXZknqqFS6iVwdsRDACo
Wx5lvLxPAyXU6DF9M8N0WUikAyDXcWQJe2rGK4sKaDIaNF2EqwxnUGQhMbhrpOc6cH/AuUOpwbgL
3ACCkaiqDF9Es3F49k2v65Sw2VAO+kQo0kNtUI43+R6dqIxBeSLfE5sZRHTbCxIezgnbsOTPma0J
jETFSAUFfY8ZYPw2AIkOukJqvN1lUYd8qWVFbUQ7KSFZcfcWNVSPxl4GfUqGQlYeRWqAgN0wUALY
WoSeut6rO0pmrmgHJLWrpXPrCdOVfXY7dkZ4UcbsoNaq4jEBKhyWDZkB8TBdr5JZqG6G4FSHiAeG
yTNd/eITnVXkA1tpGjyMu9dkEcfo28iKM15JA1kq67Ejh1CdJx9MEhhvgVBBuiE6tLaosmSxP3Jx
CqznnF/h6VwAkkvU8BL/gBFpwJoR9eRHjwQHKmrMxU5GRWgKwMDrUCpnSv4AEpureqsTuivR47s/
xpNbTFec4oT36V8XwVhmAGLjpVxJogl44D6sHkIxVHHzpg8oJqLBPVuYJi2AtYnLvnNP0/ZCUZ5B
ViN+ilwHFw+67gKJf8lp7KUva9K3w2FXrR1YdJ3KN5snlvHKuNMueorjkA+sc8FHdMh837VCc4tv
gMFGZ2zh6amgcqFhHSynt8Gf5DRpNAmdbnnyq+Zw2t/bZpmTKzayobMOSkEMIWF18mGAbzi8zdhH
i+xy2msaVr4kBlIRakyZNcKjFqbhDPsUpCHl96zEHzxbik7/hYDrj8j2hIzURFKWqQaCfwn9Mgjp
6ctvcoDxkNyUsFA2Pz+Md+SHhZkqEBLYBbt4dt5QfiA49hf6Aq1K+6wp3eTjuM3IOVr+J2OtxQDk
SSP5EQLbmf67+L3ansjpduj26iDJr7r0ENQCZr70X3fRDu308jEt3uK7reUqh7smk+4BQoYZ+Fjh
q/+dAmkZx3pYsIU2xH+EyPkr9Fq/vjAm4mpBK5bf65kNWo1YPqaKlXaqjj8dohA624h3Faigmkiq
a+cBGH7CBczjhavOue+Ax9LEP4pEXBy4Prs4IqrbP+pB1JzvlalroHzkjn7MpWLC2megPV2I2qZ0
TNxlVZ6Q4w5gMHCarMk8pffwa9wJFmrzYQRsUSu+xsk6Qk77lSfiwicj+EscRPNLj+uSialzIb1q
t1cOjTa/cIieD9qgTGa5HuX+L8TpoCcA2gH4iNk9f+cxJB456wsj0gw4PfDCYxgXc6VTYgbK5t9h
HuB5q12vdJ4HUlQIonWKnivBJDxYq8O5c4k06Mf/eXAhZ6wJG8yO9QWFQAdDkePrO9X+BabMJwMp
qtUxit3siN9VZV38XeukVxYY0CjnNPwaQlXeFDsxpnc+ifhxcmR4Os1e1xMmq2HYffJZof3/b6UW
9dSnDFlkfaHvxxoJbQr866i+r/uQWZKNScLQ0OAJw+uDFbMNG1Zvg56F3pj1cSikuzaFjqdXPIV9
X7ilAZUoX846AU4g1UCQfUjb6H2LL1QQtv/Oeexmp4/0N/ZxQaXFcn40JW/snoKH8vRTbkr7RCyZ
4Nz3YHuokWsdcVwqwLX+u5yot/e7XwHxOmmOgmRizhLs7mxz2nYpxOsbD2WNFFGrdlV1uza4cBEl
cDblrR0haspkVvAtDI6UCRmQ3KPHfigmrylqYHsmhkTuBxGAX06fpvRkHhs6c9Q8Doae4t976CIP
pKUSJRnU4UTsBHKCaLdaG+5ge/D9GWJMCAlE8o85UIJ9emK6jzlHnUymNhrkGCBi46IX92KHG134
p/ebs6ZdO4iY0EfbHuAK/YoLUfsKmqbK5i90wX5irODfhOYKMHnGiTvSNKzbNhyFIajyakOk/Zwm
b+RnVtAgjf/HfAGleGa7RbP9vdIiVpKYHEyak8XTtJpi7AJKxvIglfuo/9gpc9kY362PQ87sd5co
ruD9M9l3Qjom6t1FcMAqgqFmtoK/oy2Frig0+zXT+yNEdJ4Umhp8bt1nF3TVCHRCcXFP0zUJKSGk
U0c7rk8ltDlmO4hfs59KITrHbQViLNY1wVNnhGBgqQQoKcFxPuVFdH8jCeEw2QQ3bl8vGdY4f8Xk
qOxPxw8wNuB+aBmXfuyUqPBdUxVurhLyUdLOyCoC+AE1KabMb4zx1oZIVsbiq0NiU0u6C9X75Y6A
pGitYfYzV5yf4L1Y7jRfEbVHHfktE6JxefMuud6hb8JUwCvkgToz0wsn1jjOeCEEDZpGBnnewfXx
POFdNNsBmWj0sWm5osNB1vBhegTzDcKkKdvaA02yw9Wb29JGRhwDvWWPoD9Qf86SbIcpsrPIwOpP
kl76yzfnW1Liebn00e8IPVw63giwERZgVXCwMPaIJCYHrle3L4QJ6+wLGua2rMnGBA52o28kcPLH
pgYUbAdl+D32TgFNue93e8i9kp6nzQ5aWa9yCmsdKCFqCnp3cfnY3yspOIc11xsWdNofp/EnS9nv
oRLCrJQYePWbsTIflKoGQYN+VI+5QHMAjwr1z5nzkSHqi86U9gw1LxIaGI/tj7OocuzYd+w4jeRJ
nUFCgHm1j6cfV+rBv8OPzhHObBXQ5Xw9JHAMGPvWSgot7dK5+02tkeWp0kxnUrX6TPpkPs8BkVv4
dhh3JwluoO+p3fV1PZWYY07QEEjF7oxQMX4qsEH3a4HWDIXkxe4vVVe1gn0WyyIWqdI4ZNdfb12I
JTIqTFDkOaKSr4lJ5iL91R7oC3PswqddCcJoBzCcf4nPsIoldrJIox86PDhPp/Y6IXnWvddqEpwI
YZMnI5I86fzYIleM88V3+UQUgQxGKVsCcMY9oBPYqC450z77oqgAzbcxg3LzfvZ1C5hBSEsJkOSh
LrL3maY/hURJ5J91/2xlXA7TsJKap073jzaWLansktc7o8LxfCkoEJ59CsbIsbUB8LVIKHr4eZGo
0d8Og4a4XgVjY8LbZ2AfHl7QSgUFFW1lqHMRwXVjugpcL7kqYCga6cUo71oWRqBGtL3EMxFKoPPY
5n6yKeo8Ubj5b7H4z2WvUyNlETM0YuheiVhwWAwE1NeynvP864r0SAzv8R+fxUdBCNm+5uoqhQkK
j2JW8g/ymbcy5ceiICmd8kblOtT6L0XwoipNmJ4rqcVpGsNwNb6lNyPr4d+xUFOgBEurXsjz20Gq
MYDEVKgh3n7WIMLMGf4IRtL1v/ZBkbZXNvkcpR7CrSaKjxWbhNfFpCz6LbZhp9IhqvSi6OryRbHJ
M0Wud+jWmkWfSGG2z6ufKKQGjiy7eC0bC90Bxl2zJOfnMxWof8TwC7Pvhmh9lPRwHQdMsDq5lSgF
eMGh2n+GHMF3CiU87MSiGt/qu3WuFHTR+bhp4M9hdZEGh7bEfxP0CpRFmng0d7tGGVCgCdW08aGK
nQUmCaf1pBy5865RjzfZdy8XJF9tsjm1zvfuEltl4SovfhGYkxgOmBGxWwClgdHuDLRfjVi9lwRS
3vb+M15amb0RAoj2AYEbzRO02dculqMv0ftSf3LCJ7k5oiRJl2HIMedo/oUPveZjHxTdI15mQxaT
Zgm9PK0sNnP9ovi3qqeqB5/Pi7rYHFbsvlgtJ1Fnds7ygP/ZYLLBjkwIrB/D9o5XwJdAkkOX8wMG
GwG1slEbsfA5tCEFKY5UQjG6MWUBc3MyfqrJGpNhVO2DRRxPCyu5HHZqo7iK0sqm2+ZTNTHKKiKc
re0G6uTuQs8g3pzJvyMCnCr61IbEp39BbYVubWr7H1imjM1nFIuf24/LRdVlBElnh9/s5TeMQOyp
1+ttdYqLeKIBRujr2v6ffEBEZrD1xYEAvUEtOkv0j1Kom9NdlaB4A1sVGTaLGFoY+PAE6JVVoKqF
7u2/y0goe+55tTCJKnzWdgsIXZb9MvNCqg43oqOL79atkRRwSA/3SkA9IJKxLcIdOG67lffpDAt4
YEzMr7GcFC618TRFXrqzQC/r7P9qwDfVlSg0TOyeFgCJy1q7tuXsPM7VdLPOU1idpbW10OmCRJGR
ESjpFEi6zqAeBLqsaxReF37b2gYxb59lgVm2yFioYzB8aOTWdpo6IxO3nvzKVeswTLIHaLpmuUpY
NpNNK5sdZhQYbJDa3JnCRPSWTQi0hC123tK7LcWhJuxYc5d+jmDUD8ptHjS8V2CC4B6oWAdt4MUl
D6fX1+xBb3LdmAtF9tNgKR22itdzmtYpmly24qW4IAEtnrC7Y9AHMJtFxn35PTnCaF8paVbqI7BF
I6ihOrF/rmZftVBd/L6hboE9bn/v3yFGgoRtr2kSMU2qPUJ7V7E027b6KVHr+UCu/5gFfIRZV8r8
x7pxlOi+r1G6+b/utQEULdOIrK0OHQNktNrmN9wQo57VFcgok1TnuVVbJLXh1xdhd+hybtScp627
h5UQzwulqweJmJcsHtFevB5BGVMMdSbOraGXlYYmiQ2lZh+sN9hp95PocGvM/akZRLylikYDVuLM
3bn44FznyhMTl/VQiTAYmYV30JUCVPy2ZmQ0qYvKeXrDVowx9mRViLkIdmCslXXVs46GgqyajR1R
IudFukRRGwyJpHXokgv0BJJea5vissihYGd2fa1oL1+kyj3rtUz8ls0v7Y403lzeQ572v/YLkKzf
nk+3CWOCFWvuFcFLoATFnokwSRBCAhqy47cbFH4CIWlL6jVJxdosOXpwbxeG3ihf2YBDjzhFJaEI
I+9hitIx7E3YQH6qIco7Vg6svxzxV8hnAVXcYzw8o3tGPZpMHohU6CGSUj2KuBeEswkHXkREfZvD
HPnEsUq85cGbldjCUdDr7XsvX5ihHrkTcpn9ecOcn4TBQMozSy4ga7AWqrus5lV4J6Q5a8UULFvs
vEhXOSXUaKSslfSfeEZTR0bLGr0veP4zvzzjK9PKqM8GDHM7E9bam3QaOBhzVqo9j9/VBye7L9It
X98V3/uWRhItZXJ2i7NdveogOBDQmSv8C7pjQT27oSqWSBYe71w52XHB+ogIt5EuwcSmRh6lF5o4
C2KxarAokqehk83fSUsHsr68wWb9oSeEGTDkX8ZZaUfE2C77IqGK8UF4aR/P/UJynzYishKbEpxc
0yer0d5iBwynrvCAFFe/fh0ATpOtcb5sW8CP7RDFjTgYdAoKfC96ber6KOig+htNtefHZ7lAsCF3
F4EDovUZweBDnhHRJmsmMLmAl/AVKCiIwPAeS/OlX3bggOXkginQJCAR2RnTx2E+lmTpoqwroXzx
+w/6SOHLxTdoFKZ7VqI7F2eiyIxZLVmrPrEKGrgyOYuPDK1PvHZGtVWuW3GWZyypE4H6soIQe0r4
EOhZoV8510JglN97Rd5qhVPwIfrEkBo6YCIYQBLMGfQUpFlrqep5tm/OXH7AyEL3+Ez5Dy2+ThZG
R9aeg95fOsUMSxAMnzkzw2NXguZrs+CYRolcaHlphhqIFaaae4Lre72MF/prYRLHLbOQlyuWllPI
9++1joZ10tKwj76O6qUZmBWrf5s0W/G7MVbwHeLig6LoUtDRQXhl4tnHqJQshfaTye4YnGKNJZz6
lkj3d+gjQEnCELhhc6ByTJUpZYXIGFyJO2TC2XLlx3cuUKWfTpGikeKIYmyEwIssalzwB43yNVko
KxEWbPBKtCpr4GG8FZzOhuYyx09dgpDyv5yuuzeQJMynMmayiOx/PrEdUaEHNE9M1zHKZtynIrM5
eGeH6QmGTsvhrOJqni56v2fNhnUIizkOuHZwziuTQQjQt+pfsmW+o+ofRXZNsmf/j7YJcfMYQdJf
dzTHDn1rbGjtvz4EN8jblimYyodSOkR/IbvIC0s/wsOadcq/R3L+M7ynJ5FrevQ/MuLY/Gz2ic6P
ck+2Jc0GsydFX+kTbghiOqhLerSaAhRPrfjzc00i0Y9Hm0GRoCn4pFb8kur/+ZS2krAx1x1m9k08
MMFd8oQLf31o/qIv5bBFtyzA9rpuep25zLWLKJGbqrFug7KWy4w8wleimGBNGhCRZU22X0EXaXRv
bgtgXCi43nhewXcv8rNVLswkx46LO2c0CUQ0EmgbBryC4/bFxCgC1VHRquhgILE+SrY4X8M92i2E
kmMUVN662EJbaV74bf5/XvuroBNnoqQGe5nc4ZA6OVaR2XshzfuA3WQn51Fea8Wm6OGxLIP7Qnbi
oz5lr5e/6UF3UMQTKx1noAYkUlnmLEoCOR59vfw5qGWNmrsY1y/S1jkIHnG+5yFY/P4/0fGa7JFq
IeyIG1Grqombv7UednZ7z6HaV+0PP8jraiM5emQmMIUcev/HSZi1ow58O5F1l6KMVCWyh239E2zK
duzVcqZJVhP2H4LaNQ4pq2uObzRDFXhZ5wZgGS3k9VZl3YS6d4BEoCmEY6PSimfMs6CLCCr1SMcm
g/YsVnOp56ORTxIKhHVyILkKWrCCVq18lQfFv3PbtAdbgunnVb2CNe0Y7fQYjPqnzD0AgRUge7c5
jjAWwATGxn0Z+CTo+lb4X+DnplxxR8JK8oePCiVxHPkn1Ekla7rXImEzn/kHjqPK69N4TlJi+E+l
VLBPwn3sFz9tkjfM2lZaWUVtaaH+bj3Ak8eX5OnyC+wgIJsnLYc4Npwik/yevcGB6eednkbKxgY4
IXzxbN5Tr0Xot2f1CBhBNxfsKUAWwvsx+0llbSEbAoi+VgZjk17vDelQ7luK8Jv2PpR2A/gz0Twr
LbJ2yGPtG8oQj4/IXOwMBU2xfWw3MrC/3Vu/1xqQhNvZd8NLzm1ruOcJF7vQBmckkBKgqleFnWy2
alLyhOSeg7Yd73KgVNF4Xu3+IxEGT9sfMtqt5fSXCwgrZ0j54WQk522H5UAyQ2GvlEri2wuC2f2k
WA55QRFGx5Y23jAEAJ33GZc2l27WjvGnvS7nRJO2oSQivq9n+djC7CFF8B+mDmFJJJCy8MYJJvba
wbo0uiu4dQOwdrZusjKkRvuRcMJoa/Y0Fmr0JTinFnm5TWwRpRxdohRmzNr2yCZLh9MU3uosyF5n
Gz4m5Ycftmgy4ga+TZHdXhx0WCFQeuYpnloAPnhLpC9aykUMsRZZne3zlyR61UPbQoNFixBRN727
eWT4YHALLiHmnuy4T1XDhluT4KjJAvcNVDUjOJ43q4/aklRp/cqGSrGUTvwbNdgOq0V/LL757DBG
4/nw2CPRZytpP7LCXzoFTLAO4QeJSXuadk1zseY9O7rMoQcAd+LxJVMCbX1JSfHvEb46Ls6ypegM
juXKshoWTYgACl2k4yzwbkZuSyjhiDY6mT11JBMsmJ1NCWGq3wPfITY2v8cLggeKjE4M3esQ+GmB
uFdrR6vNNKK+wNxQmWUA6ieDao6J9fnHdVFn/wuKPyXg/x8apRx0Y37PXggCFZEppQ+JlXYDW0si
BuYPYbdBdMTkS1dSUUzljO/kG2yK9OZATSUYJuuUq0LibJOIkKX0P6drTnoG7DpWyXORTdy9THA1
enFix5xl/QJwT2DEt68EdRRkVlIipsrNj5db1R/PjBciCFw/2tqroMyQKLzACDHYhjnwgwzQQtxL
VAalkhBDIWTRoWuxAyIRNa+KleypO6bkK4a75Q+SrQyX/I24EOpQuIS1Tszd5N29fCqN0A6iqJ6x
/J7uOgFzZgi2Z5m1GFQrksIQdA9AAsYP12idyFtjAf1asQwhFi5P6sGs8g67yy2jnm0WhVeAHeoD
I9reFuH7VDO2pE7PG4pctRi5bRwBtIMLE3yOJKhGwBfu+qyVqeZk2pTK6sebxZiNA6LxoRc3arDo
vaJGOTqI65yAi43Z9gTje2WNOiVfVVGh9NpTRjNKHTV8h/8h/G3NbkBaoClqKw+tYqT7BJlSM9h7
n//ISogZfBQU+R5fGn/oFWOYDbfkKKOt280uWao1IAwvN6mExCRA3OZUetlcI1iHIhLgqKASAkZu
r3z35eJ/B8D5HpsXWLM2OgXBtCj7sTfVA6mLE0QCs20PsF9dCrJQllhXKJGtzKgYAgbAF6B0da/L
yRLyuL3N3xJKYd7WsPNpKvITK55rMM+LkcoR8quNHtGzgre1flOS5j3qMfaQDyZ+gHO/Q0vj8VgY
0UPDBWIIsBacRONe7trvY3lSSaqEnhAsZhKrYC78EEhgXh5GkHTxJr8kqXC1YdhDuBjjHT7DWvm4
D1FO1ny/OYclwQIClWwC64CfxJPYN2xC12usV5ShDMVu8tkbVUBjwl9konE1ZsbpHsoQbnf0Aq2z
eLH2jKvxFa/h7I/FpswPFXp+kk4f/uK2l0JTjeghOD7qZruUtVNJJjdTXjE1JnIUFm036dWJ02My
gcsfcEivJh0AdwNq76ETaOdTc585a/knRZg87pUgJNNAHo72YBWWmfv33JsO41n9ZwXXd6AqFvFU
JTAgNORR9rItQptii6FMLTLbyZMU3MWWGuAi2/f+5N2PgxI/fhV0Al9LlO5SpANeQc9FRUNBeR/9
LEukUeRsuKRpd9L9wNUBO/60B7jp24T6Q/pUcNzX2NX+LsWeTz8YJpcnLWS6Kt3uMHhfdJWxLS1+
sp7gY8Z84qO597fJCJxlBNdADsFZbjiE67Q4eO4j6+fu6s5qlYqGH+OjAoyDkrjjumQeOlozdJZN
OqNiGYSOB6TsRFwCgNxuxtaazQ1jZj2QGSE+T5sPhbLQqSYss9S1pVkms8g4U9qk0JnqCgNWLgA/
Q3k8tO6kJdsdfM6UBBukkbuMt/uhm4eSVjHBAKhhnWUj/sydjdLCHBBCU1QrYFwbHD6QtdIS3aOo
1ah4NWDeaHAgwFZBBfLAIzQ7VDMFYUvPnxb+YPq6V6KcM9Zr+I3e53t5Sa6PjiOjsbPQNgAC72p4
2la3oq9/Yix3hD6Sk7lXPqLwsck337+/xLzzfn7bjy0kmeyZG9Gr1ajpVrXtmGIX0+8w8zLgNjGt
4OaUrWGhZHZxTJB3nUwCjLY/WTQJKuzyrSWfSgTCQBhAIM6St75vBvGGHW/+g+NiYIMJBn0kNgSk
e8nYuYs/STGRvHueokcTEd8HMfH0irOmchVuuqeowLKCNnBBHCjzGIOn3fH8w//3P+etJvw+RLSZ
IfrIHaClFpjRkrquUn2Uwd61rZDv41Y9HUl2kY36+7MjwXwYXbhtdwmPrUjjAg98sG9yTlNVebxl
Cd7U3hQGukJO9zxsw2uA377YkRyqR4UKGa+eziVnhWFDQfXpTk5VvRD2BreLlllraZ+XBsmPXhIl
J6W2NuI+f3WoUjflvvC1TrNpWk2OQE1zuyQqp5cfeA0HvtR+NvmV6FchfDHvSppUTFFJMRSyUtR1
nW0gkOTKH7l6c2+IkzLuXijCxlz+IFqR4Awh/qZAgC8VsIKh9UIDXUDDnrEBMDPcM9Zijj/MYTxR
EesKmmORfmVGfTxHw1p+T/MMUPrWNHZ25ZD4U0a6lSZZgi6tDWjh9RpLr5TqYJb3Fqd4Xdnmgiqz
L9PvWGPcxnU8ccayPagnMZK4DO6cUKIbrJp69IOsWKGJyTeO/8cSr3qJaKVDohOqWDfvSeqMujy2
/Whbvneg4MVCcp5wT0JEjef2NEXRGPD4hL2FeUJRl2DAHsjGVBn6EtkCiKUTQzeNS/9aks+m7N3n
Y8oFTS+tJcn2fVb1o/mTCmaQouMMAJYTlmaY6YZYRij95ung9aPx+aVmvvJiXWwWgxXSnyx6dEeM
iNi7PnKVUuslOZOeMwYB63URuHeJiT2bgfSk4zQCSf7jqj3G5fLFPXSMYGxJdIkXqfGzabgS12oB
ovUFYxyHB12nLoqJ9pkzGpzlO3CqEVt85kpZmo2jPwZnqGeFEk6ltoqnUE+nCW/dRs1mVAxenlhP
o2kSEmVxfCWHeqrmaoy2oVHZdQyTo/9KxQ0sM6b0RPF9M81aNupOmpOl4/ObccZQigiDvrPDYze3
BQBfMnaUCMRKAr5Nr6gOjyoDuofBM50F2a+Dp4Ijb9q9uPiryTGcId6VSnkCJW+XqkxGHxzqL5l+
vcJO28cJ7l1nZDGfRBs8/ehSxbPcf3zraiYkPqtchLX7YvdXk7h+I82BZEhf16J61AqgiKSnmHKQ
f89jdivhGHM/y8uA6YssCHTdezD9ai4GC/l9URhmioS1r2EBbAwAYvzjRjHyYQkyLRPAeEIUmoAF
38iLIzJGW82qoUp0ocNT+OH7ox7+W9pRRm9zuIvQ1EioLRwXV5ZHEoOZZkNJykZV10M/N8jU5LCs
pYn3LxoMBzb5JWJ+nJpSjN8888/T310kkp/AxHv5G9r7uiI4WIQ8PeauKwCDm+ip60Ph5MXkloHH
pIe8DYUnoBq6RR4QZGyUSq0IeHWgm+SRgetFi00GrmkpllLvdjVh+vrEFN7sGBnqAbEWw663hcTT
vMr3XSsvwUNreZWJxIGNVyPqfU9lXyvW5k6qQwR3mzg1cY0cRPF8SEJ902aUGUv0a40d3ENHqHQ6
qVYCzg2HQDmrqh9CMKo/ql2z4y50j13Ul3zHyheLb7Ew+aP9yD23l+uIE6WTyScyft0+sQITOjoB
yWyR2wy0CHqYFUKKSrsjJZyJruKdZ6DUHK2KnsBz9Y5N2ND7RALd+shrTofynPRgQOYhGu+dE8kk
PGhUvNrxNjtYrM3QAx6eRsC4/jMit49Fv/SfaoGSJGICVFXyRuxuCIUjZOPyJEE8r9jdRblG0LCc
U668w781XEZfIN1VC8kAIZ225e6EZ0Xyikz2qZPi2oklhbirGMRAL3z9vVHMFZ1LHtQEpNVLa91s
m5ZXa8b4/zJHMCFtEjCkKw5lpKtb5bnws3/ipaUWGzPeCNyzKSCyieUZUr1K65Dv+34rQpANnKn6
u1xP2Y3VjY1kycIprBxZA1Dcxz+3E+Q6TBsFqunLSX4cls9Ov8afObnd/esTuKIJ7swUiXF7qc7K
1nNAu6BABmiBlpc+/2iNB47EGyTYmv+Do8A1SlsoWOK64T025+AOqnma1bVmAja/JfQNeqiNT2Tl
1XoVhmLdw9gVo3WDn8DD3BAalheIlO3agtWh/lvYBW9Sz8Q89U+L32uFTa5h9PIliKQe/EjilC4z
wKThKx0Q/OMsucgTLFcvitpCPqcplxEOy3BHhpid1CuaTM0H2dmcbHeILXHT8pzOgP9r9lXN/pm4
+T8IlKc9SqCPxSYLz8HwAfwGAC4EzNne7hNrwVV1gQJEULqn9aGy4/8xMWv5ojyEAmjnaiRmFzDA
XNL0Q+BS0D/wqZ2RJYtUbhQp8d1L9f4kPQBV/WuWzB22GUTrYfjDQzG3dc/vK3SqBDceKkr9Ty7W
jZKK247N8p470dRN5wot6iFpVIr/dMoQS6eBz5vI3nbzLkaovKZJKcJ4kJNW8NCTqafLs7ZfekVf
r2oS84lMbeQi1zBAkbgSkqgscd/Q/BHClQ0n69GCsxu7TNkLHUmwyKKMNxRnsdh8GTgibZk0B3FK
kUV7BSzRmWewILVCIg7QbI6Bba+I3oj9DQ2ltyYjS8xyKX3tLXDH1NXknZiHvzc1RKb9urv9POVe
VOftIlzMftmZ8uPKlgJQ3yHNMsPKpDinmo3PKZGpSN1Ca0Qlm+C4MvL8czJIdyQaVazUqji2eSU6
gJz5H9f/82/y5DKZMl7kUy9AFwxzvDf+Au2Sv8hVCA7SxBVcwYaa6Q+3J00q0CdobrxeyPxVNIKC
y3707OmqpbS4WLZ4j5tGV54RYSdlTXrH/MRRI7j9cf4Uej0WOFMMeQUOwkGmYUzPz++82IxtduyG
eq8+l50cpEL/tZaxfVFBs10bxTeHl8Ixt0/PVuvJ+UQbFt/uCvSClxqUKveg2sSZz783faZMbtcC
dAg6zL+4jKTBs3rYL08+n80WhEC3kpt93Co+AGnorS37DAX7lwoykETws3iAnpYr6OTDpXNZyOgN
PybYkt01lBgHQgvJ3QIUY2FVRf0DENJotCqq1WUnzaNgGvF+BdLLyNotynFMx4uYf+p3nnz6/IYv
zO/CK5GpIwP6H6DdvX99Ui/NSNYysN9h0spx0jiOCFx/ZX216tqdA5TzaPCCP+h2wRfMIAOAdFvg
pK4gqjJv9fge2LsuynzrhtYRnZILTZ9oRJD4W17C4ufgVO0A5L7ql0c7UKIoMA46ZDVe3e1qx5rT
FFaYHnTwAGABgKmE3X43s9hox12ilCCeXiK8CihD2f2B7OglKt6BYgVWudLidTcAxfCQM3foDQdW
O6+peeP/7OuXdvfpKSUYZRTnPqpqXpvCiWf4uWkYYrQVD7TRTleY7zWH+9DLgWNhAqBtsv6O0tNL
UC5+cSOmKmQ6ZrYivmoTaLNvvTTh0dPBLX6Nv80SrSmOB/ZwHnp5raKCJsn7v1z1ul8sNJDIsKip
UiPO8vwUA13MXFoMcs4KMTVwP02PQxOjv3KSgcdkIybLiBZ7goTOav88Z7er6Wi5pWRmwx0EZABb
yjTmSioVDlUrRLkJQrmObKjGzzpoWI1Ot509KgK6x8zN0NDmvyx0bboEEZqolujjGWBXQMsgcA9B
9FkuBDSucimPHfGbbxhVI/+rF+9C+5l6ILTdXoMNCSLuwUzejs7soXVsf36IP2oXkaUS1XFWRxwN
cbdfMoQrucAt/PYe2CeVjjQYDaf7gz2EeYWktPEeSrQNr7/H9jLW/cUV/NHuQD2Qhy5QTf59IE19
gWdIErBj/VLBB4zMKbb/Tog67ZUh2de3sG0iGHVI7Kwx1Qk0DTOQFkO5bU896Z3SOjUxouV4JCfZ
42spdNJCSE3RHaZpqzUUxDUHMNvZq+SWDkp2awLfN5/wFcr+uEypPN946MxJI4w8KxQhnygxHKCO
Xvv/eqC+pffeKYnYfFD37yLWJ0mJxrsAYNjlR4R0mt/jQA2p/xnYCDYAysH4tHrypMm5O/1bxyLF
5HUfW4qkF7tC7bdORqgn4TEiJBplnidRGorhVDmuog01ja0QKpX2UopZZGg3GmkpsfV6brLiw6ll
5wCfnve8PxDkjS9eKQbbQ1jwlOshqFNo1u1nJ6/HU9SGXXZS/62mk0H8KZHzPootnwZecy1+IaqQ
dHP6tzYinMFBq4dqQ3xizeSxoP9X0RU/wvDsyWRqEkjKRybdtdeuIdde1FJZ7nqpRUsG2r+3jaap
5xHA1BcavvVDygjVI9xSbpKalHS5lZzTpoB9ESz0qF+ZoVSK2ER259IEaz/FDBWlH7zwFj/8/1qj
vAslPRXNaFSuxdHbJq5eXjjMubN5IzAq5UefiEmFSc/WI3zB24JUAm1lk5r612FoTamsvRDbbqVi
MQMQvuK1xixLkkjyXGW7d5qEWkj4LFEJujjF7np+J4+YDrRl6UCBfNBYSoZ0QAFormxbfr34XwAz
ZYsgz+0Lgwxg+6hh5Dujn0aNMfKupPdbRA5xTlSqiYMVuRMBtRTptcSD3OzOYQoneFU6J3NnF9NZ
d944GpDA4BUj1tour+/cUOPwhas4vWsPKTixBY6MpXtnyW+WVzmQsqXyhjfKKzI5iDNBfdyWnJmX
AHUSXrYoxyg8hDmsgxWVPOCB4h5IN2KR+KYTBWAiDUOIVBU2DG8p5KCdqCLivFYhN5hYlWWlMLaF
3FyltSl3UdkTaPN/c0sRYZE/rcZ4sncwiMw3JOyRIBRFW04SMkt8rVj+uSstOVjnSJhNjzORpJlM
0ze6K6kAzyDFhMBUgWtCRTGBWrXAz3O6C48nfQAOEiNVMkL+WlMtE7A2EZN9YwBdNE0gHrjPMFZ1
Ok9z6GsYQdSIe1q6Yu2PXrUpd2lsSe4tYAp84vfuuJj00ZvdG1Nkjue0BRzvo9qm2RDcOUt1feei
nSZPa4Xzr8/n+ShVGwiznLdD7EvkEiqkIYnzHk3FMA7VA9ckRKFs4xTejeIhMx6bwqTlCE14whnk
/m9/cgspWIZxA4CVoMd7N1mdslttdl5/0ZfPz7D5Zm7YtKc7zkbQvdHXMdJi8LHBdcJtcgMlvjyN
Y6/eJtlU9ExfcL+UnRCn28QtXt3tEAURmUstpJN9BHjAtokwmIg72HZQpAJYYvG3jIE+3G+aKm0I
WFg8UCxiDfm98XcLik8l+4zkECQbt1vp5d7BEjwnASKqJF7KXkiSPM8nMO6EMkeoWYX7u6VEtZQP
4dpohgnBhrurw2kzaDEp2Q+gWj0x3+ElwaBC0R38crKltKzGt8CaZjdK56TUGkfLbLCfEvbViRpo
611UPOpJiTh5MPaYrPBY0/lOMFiOloKGWyZDAeArQMfZ6poEZvurCxe3tnfJOLblMeGhWEtabUeT
bVVh9tWSzGdigAske8AoDbFQ46CllqThf3ai8lK+JgC0FKhPWuZr52W3uT9+uB6xXpg2n5LugYnD
1GC+CtyS7QpXCeof7eWHzNhan8X7ZVwmFbP2ikOYwrMpxyCow8DMD5XKcMmBNuBy1lNSotKTS003
1b1ZNLGFzhta6WTmpnea11oRhNtqo/R3x6ygq6oqhTfeFdTcSfLGW6nSXmzS/0Wx4i1dGnS17l02
RMXbZ9j/sxeoa3t5eASV1iFC629dDk2dC8OQQ++d0WxF0uhTSv1dJG8k+9q/Utnpx6UFajF4OHwX
Tu4MIukAubPwFZalUBBo5syvaDsgKaHbqb2y7iGtLxGT3uy5KARsR/2izt+g852d0D9bRekqmU7X
PjuDwZeoiXINVSxe2aHz4tLoHJL7x3ako633VGk4tm5s+i7Ed8cu1HI21IJIYpPttYwrgyAOXeOk
Y215Ia16Iuq2o153An61XBKWRcbvy+ASWRlEX9iX92D7Q48oQFJXPw6aScZLGD9o/KRXnk5rGg1E
Q1X3cLbJEppwUOBItO/nGdGaOfoQU51bIlUX3Hm/vw5/UiRVCyUA34iulZ6iZjk88OXsvRjXSeuI
yuOc+OvobUf6F6Pljz9pFW+lmMFnc3L1tyYl3zCDeZc2iwA0k0zA4kYoTA+mEppAf1RdV9hSLvxi
0EFIMC6PcUYZWMrrwoTqIw/hp5Jm31BAgSpVkm3qOBA8hYYo/tvFJXanpzFy59TM0DFB/JxVeNOs
0fMNA26+xGF49yRbKWghUIOTCHKVhzfZBPT4U9oc/fFv7TlSmVzYlL8rlAKBLxjHr0yel1xQarTc
DGc+33AZ3XSF3PimcB6ec+6fxgJPUg7A9lF1U2AlNwkEUEp38E0+Jzs+GdwPon3cehKx5xi2jg7I
AuCrbLG8ubKi8xCQYdE4PPhltmVQZSFo3YBoqztrnbE5sMN2yQuxBMx6ORncbyZaRDMrFj9KKYCJ
sBGe3dXd06r9WthP6LMy4jtPDCK8VoGvXBytzFAhZ5ztLj7Q3HHIXz9++gUNlV/XbfHroebhED21
P48/QIaN7ridBBJkW1i84hLFl68DZcxz2egMBBaLPgPal9vHLjdwzXkAKzywUlF2iVikDahMIBq+
IIBJ5W3ts2HvPvrAWVXXfZb+YBBImTZaXFsEcsW9gew/BXQNKTTPipWQhhgBBLAPj01/pNAEO9BB
+4F4La0Rz7S11plVQoOjWlb44DrX/4Tcup8EltRX70/vHJEJtAXCpOVNxXZhxxKMaqR7MPvZB7uI
UwNv3Onz6M4IG+OREI3wTp/tjtURGyLddamRfQhmNb02gDgMclISJT/CUQz/CsEQMjTSN6zmwd+w
1xXCSJdlOpyAyQNxXWx0qkfzkKH5nYMDcU5SsmtJng7naDxOSjDTud5UCfPnJZMGUlqCd738P4lP
prTTgtO6r6OfvGcGe/GLn8tzzwAkQHfBDv/hQJJCSLMxEsrklPr5PlbnuI1vicPKGidRhWhShIso
3mClf1I3F/95XeumwJdcaF8k9pNEf1ViUQz19hihFIbhu0HVOKwc/vCcgzO3Hpk5q9VZSlScpKHm
gRXNeVWVOgq707vLAoJxx14mMbfX6bf4V91amClh61ihq5+aWF9K1WvRtJJzGtuWJf8WovbzlZQd
Ql+XQLAGgIgJTJ2IMdX0v+Sw/Nns5TvAV6QJEv4ufWcGpmqQAZlAurSh0fJQuldMBpNSo+Cip26n
4JswUdC6NO6SaF0a6DSfa/vDLL0lnp5VYHrQA4jvjEGvjcsOdRuHU5Nzo3ckkArikeR7RWITQbbA
3EdpSNjO93h1Uh8oDfphr6iDMidajOIm0lYXsN0bdzWEQEMmbjXQotgiaz1H0eEeAgu729D01vgA
UZ7n7HSa1iXBQ9WQGagx2BhILNrftB5EqVCGb5tY/9AprJaJY2thTGJXzp++/9ywdm//gVMfd14X
JnZ7HxoQQmQYz1xX1cS1DJsYqFmxP4Oxgirp6iLVJosXIxIozy4FTiFIO/Uww8oVGf3zdEVl2ZVt
vWDLcuoKZrYNSkTgjeVUFs9rg9+yMVNva4H0CrcvFH5vrqZow8a0AEHd1f99CRr3fPntJRMMG5H4
X4kwtyZz95fHmfOgBHujEpSAaOUzX3fvy7i50rwLuUTDZ2LEC2bshOCA06Rjsm3JGoJrv1oAEKDX
rbDbbEHuTnm3tvws5HSDLk+rQMbSgvT+37qEoi5IwCR/BSORuKguzWxLaKjLtaUdb+J2tszjHwM4
JR5fBTi9FAa2vGJr0EQNx5K+YKGpydw1l/GiFxgQUMPOaKhMMxeXVqHRQ3e22cG9ByWHVKtxvt27
/D1rFm1yzmds8KGYT0UxA4CY3pURocsTOPFAMP8QP/6d6TMrchDt+9DUXhdmWZjLAXHvoSkje4l0
KlgyKcXQElegxWj9PjYFbjctYPvuPzr6R7Hl2nm2tz+n4BI6lcE3fubCewM16gQx8zmM4Eh/igyO
nZdhCjFBKjS4thj4CxeLZ1yPIytJpJ5cM5PE0g9QURnyNpPwlA8DukdZGrp0PnzXaTYn5Kgb/+0v
ne0ajlFNr/n/kdDQsD2r+zdumLRHxkMD9x6qbMgNkp3ef5DDQKiTHx+2ABK00YJ92G9Vfe1TiJrm
mHHlG3N9qBXBa6IAldxxEnPGLdI2+VYEqRQ4JBHNBL41ICvYgzzW99K9vC832TaKPWJ1nZoq+WjB
5v+xqDDUWpTQ4ZeHwu34D6s0rZv+3Xd1PLTEueuJB38y0KCmRuTYoCLvEef/3MdWz4dZMhM3c6l6
mUROsmN8q0+V1WQvIJkVvPxa8LNhsnW9lA+dYlBi1rjsMcCRvINpsbgZiQKDp2QXHWTUskLMubAe
mcrS1bo7ED5AD/gqau6F7Ov8QReFHJiFgrdAZ8CrR4Wk6PYLtaw36dc6xF8eLsUDsCoU6ZyOEigy
TjRmNBBCOE5GO2J54u87NNLHVDXkevPQ13VjYbQ3iQo+wW19Y2n4HQsNXoMbZk5uYL1BcSEJUPBg
/0g2ms9EalspAx+jL/GIpdI43xkBC6kcM3MhdlJPUIRMyT6bnMw2JOdQaP5f2YELLbsOaICoDqCj
NwMeHbLwXu1BmAcs0GTgRAOPahCftTwUgfJIXFQITZncoub9He0XSUDnEVDduu8Z2yUnxlQ9LdE3
JRyHrnR31KaD4jhPbIW3iQyeL8i4YTb+CevjrIDuzyPT0gEb4teZih1mZVIT3+/67WUgtN0Uw2bi
/vkbnm+Utr/9Uk53BejKYgeYocLf1g7azh2KJcrLkJ5NMN2yn5kN4CIGQ4BHdpUsIHHc9StG/Bm+
RmqkOJfOQLQfkPLe/pSIUZtlol7pBFp/cdDuWU+W9zIIrBbh0bcb/BGr7lPysGYARkM0kd2Bsjan
7KYCJabm7LRDUO4aqbk32WUsPbMaN7qtmHmp0I5CgEbLYQ9AQirfUnnDbNQ5NtyHJMt3+HUVPCmo
/OLCX5+AmsTA46k7QDmcpb34nk1tix89HsVuMwc+5hPqI71/CVavRzvyXIwdRDmEPCaka0oRBfL9
17KRVnIjCK+XTOcUcjEgzkdN5BUBL6oZc1bcwkhDxaWv9YoX8RMyebeuOFn1Q/wmLP8GIqKYztkG
RYE0BnAjKWevPWhdZh9CYfJYYlQuh6IYwy7zCAq3PXIOsIZH+b2W4gHepw5vlAuMkP/CJyiwZRHP
HSBX9TzOp2lVqyUP9pdOSMx5f4R+WWDqkurc2ELR5gYywDVSleaVrfQBeAbDR1U/2vEu4+gI0YZY
O62hqO3f0c8b2s/GY7EDbmllo9PBDwog4QHXhY92Txw/5cFsyKj/TSoJ36/Gnvu+x4Cww90nYQpy
UrHMTCUH3M21qa1+xOUubBnX9E1v1ryHad+AH15Hx+LoSv5QovFq2EcpFmujBKeZ79+NDG7FQQrp
+rkFd2v+yoWQgtxHJjpYlJdctrFgLtVMa+h043EA+FMkZXg3lXYV63AGheiKQPcBURmQwKh7IP4z
uf9yLbZcTqoCONx2Q3QCPG9DQ803EiAODHg3lymJLQNOBGrmL1P2Ct/kitqKc8spSYZL1Ex+IN2J
v4LKDsx+zm/HW14VcoBWLvkmQpgOK/VsY2jHEE+6ZQ2Zje4O6pLaUUhznJX7Myy6PV/jogxpueYU
/EXMxp1bKrX1fh90O3QzJWW6KlF/8IrdHGBR3fxEtrfNgBeQK40rE/47JUl4td4+A21E9vml0pKw
TdsbRf/QUmCZAN/TgwnrdS79nDsaVPmy/8qYOvlXAfp9BdEDaBurOmmIclQvCULXN5x6Tzu+hO0P
AxaEFVmdISbvQe6i0Ea365urXhmzlrqpSqc3C15yx7ina2HC/zFjxtTCzhb5qh1iukZnesUdiDcn
6lSdng6SMWHx8cKjWXIVtiqS5tC6aa7/he/8m8lEcP8gy9ghzxa5XBycbxOPEEYdWRCfJu2osDAT
o9+Pk6etPLcUJOTc3MjovPMgV47O2ANHHpyXXfQDZUUrn5qejz1CxTcDUx2Am0s0z50tSGtndgRq
ZeiZ1NgL5dcIvpvTok0KhOGesgamB6wX21KxAyL/rsdradZ4HQ8ECIddzlg5j7ZPhTmPgHkOdvFE
igEMrJCs+aIebYuFG2dtqjEWgeqD0NYQSxN8iN3yPWuNDucG+WBnBQsdnFQD18XO57xScjVlLYgz
/QYUDxheeVhOzxeQYOLEP01+3khlkECTfgA0+J7QZYP6r90q6mjqGvpAXIeAsaOzTPTyuaRCHMsd
1xUB3vFKp+Apllolz9Qwf9XhGJ64oa6tAi+UoymVfYrTBzovl8LdRgoNk6EEd+KYZJphpMf79WZi
kf8AeuxxYrv1JcyLELXbziB9oPOajo6gcM6oG+QbHQhaTrgOiunM7zDkLM8f0+TNLTL77lwerg9c
qSOgSvvT0PlwmNM3GRJAd6v6vUiw8V7ImrMcAQWKNN0y0/dz8EkBHNMtj/1kfHGMaPLL1jo+U3Ca
pxVBBOw4m7Oi9yWWZvA/MBWAQHqxNroYpFGP4ezBhASHcsb9PaK83xjS74Dtr0cbz9kY3mIOFbJn
S+1t9NuOPt8vAFB2nu9V/blYtSST+M72Yg35zNEvOGHqVfElbdOgknxxzJgg2+lm31kqMwVBUfri
JdgMrYFsXnlX/pg1rJsueWgnRt8g2ONO2hj7wjue02jq2PMfb2THqGxQfcHfBjJnj/2l5rFBwQXY
mbWqeulkl/F9vjOpKl/1XBTtr5ewqsfG9r/uA12cGdcLXEj4N2qJrC5v8oREdvPIl6WXcjiw/QBD
ojzFPFAnHQ1rk9MZRGBoud/ND+9hBaxO498k45DmzYbwJfhYertd/mTrU+qnIuezD2deUOWaa7oy
Yx+YXAeaic1Our1IhlhRfzdt6kxvTmevHqQd+Jzros1yY2yrDSrpZfT2Pw1nI48H4hhWnbEU8pgP
8RrBZB2cIUo/UrAtthYKD/ecm1iZNibg8XBnnb0BUoaJyiH40LU3n7tZpw+OZHxRReSdyRni2iN7
Nu1ejZaD22y5HwOduM0DPnK2JUYtzqmPjO7ZCqtq2uF4Hfz1HNtxtETXmcJZ8hFlA11fj0vLEIa8
qXhWu+diM4rGxUgYooGedIeHgxfqFNPRiqEZmQ85SDxVw4nVN5KUmz7lHBxegf8iQj/KeCkNMrVk
z+SLZD3mAKjv68ZFWJSWycrqAlIviyyNt2c4wj+6+B15932GTVlU8qALDUV4QTrelyN3IyYcaTev
j/C7MmN/br5DlD7Wv6gcdubVmlweayDpyR0fvnVZjXCRxDGEvOENNaGuzohoHrYhT2yNAVBA3Pme
j2zOS2Bm6Dh7BNxC3VEIZD1JMJpoW46R0UJanWe8lcuI0UNmheIxfhrS6v4IpLXJ50JBlPxQv+va
hVcXq4rCYZ1zkpQuqmvXKxURxmVEA+505BbhZDdCJlMYPw5K7IsqyIllqjmgN8a/7XwOy2sKLmYa
CEazCWz4+mydu1qtgWqNoH7cJ9Vq0PaZXRIL8HHXnzVXQxRKd3Cc0tmlWL6WSeCeTVFokxkxaWV0
AQhO89JIibr4ic6nfu5ZYIekpvjeNVedC9+44MX1ltlNtU5yg6MV1LBdAsUOs1ZZ07LMEBPAqom5
qicrIIs1IS0Af+8BJogG3U5czahuLHQ+09OXWAjflp8+OcGDyXyoUVfEFMx0o/6UlVbzph01WsgW
IRFlFnAwBT7fZQqfpvLK453vL36mp+A1mf4wcBSPftBAgESoIj7qIICpnAX+N1OkzwpNOVmO73Va
z4WkxshOkpRTA5fAYPDpWvKcp/cHzcGi+pgyPpKHUor8QbPqFBmlRdHuv8T2kmQG/qTjCmcgWlgv
0dIwZDqc+GvpUR3Tw6/5AGJFOhxzxYBSktK7n6Al9kDLCr4gPkl8/UhG+rOI5MRhQtO/ZJn0hAQm
sQQc2DdGe/rTEM9/20+ZrjYV1izrNLt2HxxQM/nHsdEusZUPTqmmM+W1nKo8RoY+jjJWR72kFhrT
s0eyYzcnVPXFl2383+8C2XxKfgJaNd/Ppbnpq8atvXwP6yeQpbk9pfEMP+WEZGoqAviaqFwN3ZkW
BAOyGDTkbZskNVhBmR2ExBSGQvwFdFYifjX2lUPGP1fpNWgaVRcaavAEfEhPzyo/eb0vn5uV/Rkx
g5pD5eos8jejGZMSEUbEv74KaKfWY/n1nkXG71jKlDfiID7Tb0M4jJ3gi+CI+htO2QnC1eMAhMcE
0v8Z3O7yBbX/ApD3GUZxjjyma3bG6FdsSVEy3s80abGPe3ejhenwfGtB3HXRpR/hV4Ysrvpc+LNF
GE1kzs0fgiKFZv9Bz99b7QEegD1YTIwyE8vCas4iqVOIM6G3xzeogeNT2b4OnyUMwjCfYTNSWyy4
2vSNanv6Q9T7FzwhdhztZaO9nE7LoB3w5rcbq8lK3f3W7l97q2YV95fqEmGLqJPPPLr+skJN1Zzs
sG7r5779K/KO4R18AzMJmWW6wjqi7rhj+CmDFP/p8EeTFUuemM8+JUTTGdm9XGqH4ARLJ1Y0VGo4
bU8G16BvAMzfu48k7nyQ5QN51D9gkhOMhaPh1S89XVey5X4vUDq+zsAUhuCEi0VNbpj9UxnLDAy0
f5XuzvJZclmhQT1Ue+AXhGj+XzoASCDl1ukI7jsRNDX+bhpJ6IqfdA/Rkscc83gfYFfU2kGM5+52
70xxTb0UAkdfxyKxuBso0Zjenefhh9sqXJLvANNddu8O7amLGHmiDXRSYXwlZb6/zh2dZKTSWusY
OTL+QA7ibYhgWMrv0/S6JYSOh7FZgfycThwxUazKCcjHhEAzwKQedRfEmpqet4SoH/3VzXbzgjiB
Oa/q2LpNmFk4ytrTWg67phYmHWaOHvS/l93W/zs7ujUC1b4WwtWmuBilndQ5a0f+1cC1srCz1r1U
qAsZWxtkoe3UEhJo8MPLVZUSPhH4ktQ7FXOtJnDalybEs6N7BziKi0DqzdBSNg6+FjaSp6WTSc2L
0dhI2R+EqMT5DoKtjkR+krhSJML3r6TwbTvV8HxUSiaoAvGLQlVuhDOGw35Rm3Ab6zVX8Gepoeek
j731UtmAjCswlDHguRFEDW4eiK6H7kBDXb1hTDP/QldY2AXPhK+g1qVI71MFHHBYsc1ws6/zGHJV
Bbw+GIVbq8KLQ7iJ2ERmXZj7UYfQ0Bmmo6Fos8U2tHv/XTPOQO932Ez6NLFn9Xq6uwimaFnqWDnF
3h3k4aTgZ62NVQ82Y149pDm9KNhYhx10CQ5Tu6zu8s/2gh5+GF9pkGo1D3drTR5yC0lGo2jeZ85V
LJeeR2oZaj5F0kpBPfjb0eFdzcENM3gizWwu7hF9+ZaftaY5WeQQpxNY49ssc5VLZYWXsYQ2PRbC
W05JpbFCbgbB8PmTxNy4vhCiNwmIVU2/g+MLwkOUM3VioBjeZBaEuM4dcmdNNq9kwWZNA33r/xIA
8MnbJySRqkZL9RuGg3MHjj9q7IcCrPs85d5s3fuu+VaAVpdHBxNA7iM2g+zNbskwON3XrFhy6boe
oyAhSPO6an+E7OY5CzzjjBlb6w+HanBmTTUuVYQs/4KCPoa3vpzITGLs7yRMtP1EUAMuxmnJ1eah
h3HbuneEl83ipM7sfzIrKhgIgCB8SZrcpc7TS8Q99yIaH/ZhSFhTi1OAVdkff444HqjzaUHL8KKe
12+Vb5Kh12VVXxSe9ZwnnPLKbFAa1hfKlBjW/i0LhdabtRZYVnR1yEoiK5fQ6WtiNCI3el8ldLgU
eO6gwb9vIB3qla+KHz+ynYxXD+UScCiObHEYdQhG7JTIe/ePLubmWkGp3Wfkp+HaN2uQLVb72n6+
c0LVCegSKkbcsTqeDmX3NFP01lMt53mCyACPgiSAaphWZLUxDX/juNrWID/ycpbzPo3MWxV1Ty7d
bivqG3ztd/2u8KlHx75NSL47F0IQXvspuum1H1ZuaKxOX1bFIc1ILLan0NsX2p8U8ZUC7eeL48W9
2NGRVHRUSG2+0XOO6bpxG+TfF2d0QaexyGIXsverdy8X5fJNwS5e6pK0q3OU4sV8E5DDXXK6qE5/
cgZfbm8Ue+M40zOCTnntDU8FwBul7Fj7jREAyuVCwccG9HIddY/WdAuXi1V6CH/7sdHHdErZu10O
4tgh52d+7clrQjudQjUeKZLsnrExMY1zG5B+JsUN0sWyCchjf9pnepmwMbdGmNnOWXFtjlC0b5TC
X9D5E7Ue2TGRTqzqf5yQEK7KiFOC7RQFSFn2lV4RAsVQaXJHcGqnBIrGKQFJHvQGoRH8ZM0KDvOK
jNssG0KkHSo38xnbC/4gDq3K4o86TIUWpPSjGzwKnGQjlzFqc+gSuvrTwIyYkajpSnkh7S0jaji9
WrlAT+b33WuPaaQdD+zcgJg+dIQ4RM+djEmUw/Cx/qWsZE2uFCxHNIgi5bUr/++puDVDYZfhGyrQ
bArvuQQbf9o9NzGT1I4JiMYlw+zNKXZXETrZBt2TwOFU9XiQNq0MpgRW4zD1MGlDd3syKqEMonog
vAb30tfhmmXpsZzh/TwBuS8EOVog1FPWaYfZGFamhBVQeQ+QgtSV+TpMODfPrAQgMuWyijnOdyTS
FzRvQBDNKrIzhtYVFRN20d9aHdTDC6j9Jp6j0vYfNcmUjUBo3lPFykcRGsfs5TOb71wxawP5Kshw
pTQqoYJ+E48BbC0cSx9eSgrEfQg3Nztm6SK/gbM6dNUfitSWrFG4EHTCIRMf4YlVyqRrwAfzhrL7
pSMn82dH0el7IHWktKLFE/SU8K3Odl9BepYe5KCGGnLNNRowf2/p4r7C5FHVavBPl+MZRL2CYyOM
YFnqteWxq0PGq8umkkA4dXmPJCsX/+Z5lD0YRXqqrHq5LiY/uCx/6ckQUOLh6gp/p4lWCe0Uc0Nl
LMVX/OOzRtVb+3cD5SKlKsBGajV5qDfLvpRurAVVXTWQLS3hAOwOtte7yOP1EwgDeTTjDbjzyQpE
7HSzLZWbvfbIPRj9cJxOAdzg2JYbpdtH0Bdp7vn3Dx1YNf4FGNcuQLFvgBNnWQnnTU9voTr+vNkd
SygzhG5Z55DSwT6zUljYbhbU419rMMt5Iun6YXR1GVXh0JO4pG7gXxFh64r0aNcBnNwRI14cs+KX
zUJU50mr6E3v3yi1hqeG3TS1uCsCKB3r2NzEAD45vXUvzRPo+nip4VXwvMWBf52c4ZIArB00uFSS
6j9C07XUWSthSDiIe10MrupvAEaxmLqi8ddYPFnQ/coXqTBd4CTJkF7H7h8o4YwfS6vieju8cCWB
Bz+yBj07FZYsyISOQuCgxeWwu1iAeSgXkawjPh7tIJnWvaz/tIF+NwbpBf7CnvGnAdxnNsIkHhGn
kBgS2ewiULOxyLMRxICOIaKXdxVp0K6qjZZAnIw9s5DLZ+wU2qqqYP6giIPdYquPFGkyPITgfmM0
p5wwktvg65/PTRszPg78GVTdj2bnerSHV2IXCwf/qgUl4W38O41a4BBSH025SNuc4/iJfkA7LicE
rEWOVwmgQYV5R5QUNo9C0zAAvCZeOFK7KAITU4MOlBze7xm7I9hqfKuyJr18MleUq0AM4mhf1+an
BGNu/ZCiDrayLHQf0oI0ljlsPeXCmqaBAoKF8H2kQpLuTds4kCMEu+Aok/z/5nk+82UVxyYBl2Z0
F+4K3oZMHyErTEJtoTWWwK1TbrJO//PZTQ6pzASEjB9POKts1WFIDwuffaaz4ntCIctCu0bUz1Ik
zTTCW/R7dsdtplnd4ha91zivQTJhoYU+qTe9QZ3UvMXI7eHkEy4MO1+75Irp1lXwKxjfSZkCLiSn
MrtPZd9YkhNMNGg0NkMw3c5yH5lmebtbgnPXw721O5c5dNNYywYumKCHw9kJycUQ7Gv4bBySU8ia
irNr8Uh6KD6aAKy8uRL0mudgJTeMDOxAd+YMlWC0NJA4mIsha9jGh5c7r9NDk83DlLCEXiHbMbXU
3AFYZjkpITYKr3Zsh3QG3aECNUOKr3sTpN6yY2z/rCt7Dw1Qet3rM19ldz/kjT08ejLJUDhTBhwJ
SJgfq2uqFt902CFgSrzvDmGuqOML0pXHwAmcgjyaHZacKial9nKpPRpLXnWod5osvX1w43Lq4y2g
KIHzn6KKPy6VJJzjGHsAODghvTF3ONAfuGy47vFNY9FZhgjBuM19Mw1QFOYd8EqzEOtIvKqj/i1N
1JVSja1IsQAisE2FTKrWt+uLCzT/Fcutj9c7KLj2nYIck5NonP8GdYQbx0dwO2foshZWUR1hja8q
A0FFPvFTYsn7LM/10JeLIWsPjcLVdLu8KztteBAi7aqETmmZoyd1MImK5NW211Ps9rPAuO8sYsst
/r5Z1bvn1CTOaQPyq71axmdNolN5nQhQdaZiAW566rzR252FjrcH9NOao5qY0r9c/pXIn+ceG/ty
e+uOVqD7o2M8mMFAq7FYPhgM2B6FPhI3kg7hxeSkI3pwdJaAPxSeVvaTAF1vkDSqafb+IWWBGCuC
oODf1n/gl4iSIO098DNOjPORDDiTTOEwoRInm3fPCOn6ibv0UWy5FabaLtAPPXzDOg9ru7pZn+9G
DToS0EetQzYKy/7+jWCZTCA09YjbTIQhNwEFqFqZC38z/GvpgSQkZlY5xtJSRkE+LmjFq8VK5b1/
qNCYVCF8GpHDPf2IrdQtTQqrD0Vi/ZPRVJaBDSNvJ5gvot87qgSEaiLGkq+JZ906uvSUYO6IzGTI
3DE269nDJhrmMr6pZ7rCHTmBQ47SVXJgF7wGijw22L4EcUb4C6R/5NGxWDae3i+8g/NEHK0qQrrd
HP6BubAwh/kgIhX4/3rfptM6t4vKasSnJWPrhIF/vhE6+aaVYQFXcm/RvzTl20MqNA90o/hAPwH8
Dcq98nF71SXuSBq52iY5zwTCNf3y9xsMpWzFHZprupHRoa09SZDfFn6LxgF2i/qE85jkZ4I/XG5H
7kiX7YGkgAlDVPGDhF4jiibVBIGYIxxTTYW0e6jE+mX5dZJbdwXSe4KtsjZKjUM/dFMveacaJVAn
97cbuVpl8IiiGf3hdYPUSWd8j3I1RcnWNk37+nxEWw4BMYEtojigFtF13NS8J9JA1bV4gLcKQkfM
tnMU0kVNrP6AoFDXTWbsW1Z5Ln5+K65OYMt1EL8oyqOVGUIDnhOrqa5wMmEMrF5u41EKoQeQDTGs
N8eu7bK5W4uyOfWD7FlauS4Lz0OfyP+0JZ5gF+Z5gjIGVZ1elbbNf56w9uziMPqx6VEI5bIBI7bL
27OIuncfCPrDLP9t24Miv8mR2qg3tgYu0e2QnfHNgrS0dvjefQ1dus6l9R64b3oCyyjOZ4eQaFk+
HW4fWsIlr6FIH84MgkPRaruKcRhhAA+UXYRh/YLpH3vtJlOqFRCMCaDa5XZQZ4p9NKDSKlyxFMs1
EarOxhwZS5HIFbceliWmmmloMcd0mTF4HcKEfCQhqjfts4GMVdSm0aElOUIfdY5enDqMUwMC9iE0
s+bvW8WjT7adDp5wW3JL0CNxsGmX4MHPrljRqF3ymCpVfVfjaAPiHdWsmfoKbqeRyDyQb+56AYJV
Pdg2D6KiGF0viw7uv5c3q+pzT6/c54nfB4sIjwhzantOFPtvlnuHpryV3X7P9aSyoiBKv87MhXrn
MjYm3S77tCksnrbbPiKnyhwF+ZBuZdJV90LH6WLjkCcLDBzSy6puRxLreO+y8GlNLrW071VVb1Hx
A1FuJLYF+E5VQYFlpkzO0KOVhJv9WMcLOR2n62UelWMXWrIHKRxYc4WQVNudv3YCiCTGUbnHXE9w
WGUBQR+9KHS2pbt36/LmmRJKNHW4NtGl5kJJWGSK4p7N6OQbkG4hCmV0zdcMbj8ADioff7Qxjzta
XitWrYZwDCskFbVOQAFWw+EU/n98bOGQE6QfBnaYg2F4Lx92HSd8DddzPb3YIslMybLRRTi64R+Z
CFjFk2TJuvY1QyGgohjXgYycIsAbIBxV46BCrzcXs7SfG0N1SClncDQZJZhEUNnM3rzXD6mdZa6+
C7PgTd4MWO83AzbnBe4OoP5A7LdXnLsLvspoN5CU8Op7lOci8Ok30ximkbfssw0BsdmYHOEeRgqy
lzXQw/L0OOqEF9TnpixY1Th+NGPtB4mW/ZTfjpxM6XFUWU2V3EYvKRD9PfbcaJ0g12c7GRaMlaRU
OD6fv7sQVjirrtarAHKLCm95+MuhNf2NkVem44hTBZl9jtQsSZEeDPmKdAcSLrD6UjONLNovOQNC
Dh3LaALCppFF0zL87/blOTF3yZUSxrAZnXlHXy3VuSMynyzWZcfBzYgKqeLc01WNIzKJ6x2MP7OJ
AtUP05lOmCdfY80uywdxiNEik4p9hsWGuSuEaUBJh8QPs28xiTl3Leg7jHjDHWuUkZOzWv/3LFeP
rdQwBgm/UJtfG8uCvuA19LO3rr9ApB0GHBZqeqpJ3ZMHLvtqw6CA5tWzufg5vVDQi2ldg41JAO0a
bHAlf5U7zLSpdyMP4QGeIsRedt6dqLATWN2XeZuMxUsi0oStcR7brBinPjO9eRNMOb4zFLlBcAmn
jxIF6m3nvGrClAWTKRElCksBVE+cjwL5nScOX0iAYdLImpF9pHLEmCKG6Fx4JXGWXjl/0mRWEqUd
j59mcauopDEN6bBsZAAvlAdmUx9w+hGIBOtpi26+XoXjEHz0oxxWfygVh9oUH9KvtkoIJY1n6jPN
pXzGAD0BAUJP1sROHTy/vSJ1+hDZsjD4m4mzVksyHD0idoOMTwHfqvSZ5xIN912iJswdYSMHalMW
bOY5e32kEmISUiQFpjVpf/yRdBgjS3i4kTnigPBBITEJtb77VcasIFS3jdgTR4IH5eylEHFiGu+s
j0Lz2Zp+7kbmD3xtNteeikkNLKVLgUZWE1GBlQcDpKW8OoX+WxpMMCthuDUDbq87GvSfwAJzOn8M
Rs6o6xvh4pZnVDQdAWBf4aV9KMdJtqeoa+umYwxcdMqe0DIZBZaymrrfih6wWMoHE4ook3wIu0Wl
bCxyGidMckB/fv6IAFuGOR2eQVP2VYQcC2lZ5SN+D7NAv/cQsDS2W/ekH0E25fZjA2YFLEjlvnG3
P2EAnkag0b+Stw34bpW5Zz0xLJyTjeDuA+ql0+/Yl7Ct2NJat3eGcboEcTOKl5016f9EI8uurAI1
ePnAQ5So7l9xUNjXVkPqsFVF0P+RciEQYOWVBxZrmKGbiggiIlRdWaeYbXi/G6m4JRuxCvd9xcFt
uSD1OR153Bcq23gqAVqWTfRd2ExskJyVfT03kQBaUIFxjyMDNoobUUhcokaxIbM3RiVcj/9Yl1W2
gxXHEsC7JFV7ZbdB8Qe7AF2MttADac003c1gyWDeWcOy6gKJdt9CCU+9LEaLb6u8NOKTerQG8Kjo
POMYDvOz3abSZXCBAfC8K4hL8j5Qru2Ir0wGj0aLySKk/uPkiZXiijpGtC66pEf7vnjJDHrFhcvk
lydeIZH9ynhjf9Ylq/LEEQoGeuhCwXEOlNsjasF68SphW7ir9GqC8Ta4kqSjJFW+jNQXB0+O0DN9
y8uBEALAXLY/8BeIRY8vqfyGKRuurULtnhWe+pOYc5PWaaXfMiuc8kSYG18lNsw3xqStSLyt3HR5
ZYF/tSHOv8iL/34AZVzGAlRVsY/kVF3rt4bI72f3J8eZMMNN7UEPXU2ONqKA7bwLnxFl3hhv2HPu
qqIMjZZ2uS2PlGRehBIms9d13mu2BlFr1EdoSian/6l+T18TG9S7FtiCk/ygC4641dRpeWx+6aaB
p+zGZpx4kFcODKJclWMkyeO5DCrDVCwMNrqSYoWdsV5XwmnLR4CmbUyu1kBqETrNrBGf2Ss8N0zp
Ok8v9eiheH5o3Jp8hFdXS8CCC7Oo7fTzVxa9JUGW/TOBJl3JtgwlFKW8koBYCl1jZkn52OjTxeZN
JQGlUYZxtC40SAOYXmjRjJYbSFFxU9KpBhE0u1t5aeh3nHOrw0TiZmfCbb4cTxFQNUoXYbpB+deD
rm3IEpvJGbC9Uw7F+F3MEHEaYTfaXuifWaN9XUrMl7kkeFuDH/B6NSRN16MvlwsVCKRwVlvqu52L
7H60cAWaMt/5MnKuOOv/6+EnnxYP6TKjJr44nLW2U8zs2BOyYr1Mu5Cq+UjGGr6p1/cTeeSshype
yXVFXO1JZnPYik9/k74L4FDOuYHDllmDywMXHw8SRpk+1ZhUgFMGZHPF7WPvNKJsCs8KLjHIwfp0
cmAZIPv6iygpzKMqOqz8jObwJgOCd49GjueQeQc4eXR9BraSrSC0dFaABo0m5DyeNLX+U7qfCHQ1
GXG09wSBcDDcyowpY9BqgKvlTXI8Ss9OSBTeumMwpiLjnHTXT+mnz6VHEtcTTS5ddRkq0uB+Lh/Q
yzNDpXFLNQxU3RBVOfrSqqr+h4SQ4vpfWh5dGQnruyVAHYY8o1Ddd6hA0CO4pyNWpEaKH9BXSdCf
QDDXB9Zd5bzH0cmKI9RHLFcmWagXRuB3O7dtPCRtrHYA9awiKlDVpNS/HGVsa2p/7uXdp2MAizMo
Ljnfho7GaQ1pUW31cKYthBBfaRQLuz2RFa6zHTpAggjQGQgasbpjN+j7phlqDzDR0mWDvdCc6Wg6
N+DkI52+08cY8S1TtgqkYOC1WbE09Uj6+wFi6UWRVG6xwE7Q5bXhAemkbk9Gde9l7YvZCx8LaJMT
/1aILqHMwpJlWTBjNeezFtc429uJbjt407TNnkz6NotstKcKdmXQc32cin/6/3tdz+qZGe3gysXf
l+DW4lrX08mxlG1J0QAo5FGAWHNAGjmwFEp+2ViNtj7WO+PPlovz85WERp1w4b4EV/d9vZ13YbWH
4kpVZf0TfUjfLAtYYfaExe351qZKfBnyVZ1E2LleUsAsVNqi3CBYXCT9ks2VECZe2ad1I8D4PKmn
0rM4iSDjjcrc7XPOHW1xB+r44BYgBr/h6QCF1nbfz9NwnyQ2rqflvdPtAg8Mo7lAuSfRTCQNyjqz
GFzCnHNq/CovaqRDHnorY+Q5W43ZRPv7Tu2lS+lGwnxt3mMvtJIEqvHeSSWTVUaAIWlMSA9YMCPW
E1Z6XXdXEjnjqVECORM7t9hGMm1OiL2uXN2aZDQTbwhqo/hwsSFmeRuUAl+pn7o6bAKsedR8huj7
8dwWPcdHoQ40RH2N+5bwbhP2CQUaQxeagRAxrswN8pu2ComOC2GTrxRgYMcW05XyBcnEiqhMuRGA
9r5ixwYHg8/s4jQj6SJpPjiwizbslcgbqRJJeBHdKsEsqEk1rOtzdV8rbcl98KZL7ku+MjB/LHLU
wdiPIf1NkG8kLtJ15CXPek8KrQuoAnFG9DU8tSecX4TO7ndtf8HC5y/t+1tV5iKH9e45O1oxQjdv
GjQu2iTk+0sUQKocjGdvtIRlMOLREvBLJtcXtILYuvtMRKAKDmsm0vmck+ubmXtTwfCF9ClA1XxN
tdBWNUwVqn0+HNgE12+UOzZL1mvA9TOIzX64rckFNCne/aDBAY/9yF4f/ORGMdsISbFV2T6Tz9VE
wH+OD4fOO5jcuvMjodEUgo6SizlvsUOg4mU7hx2WgEq8I9UKYnLJ18CYKFEMvlngnZ3b+L2hOcHV
kPJKEJTE5r7iNO7rlse+B+8rHPmAG4O7s52YwJfNtMf1BDVEWm0GSUR4gHuSiawVgPkxLQlROl+v
yu77Ml7q3qfQdTX+pAiOHo4Age+cV3rJlmOPxyQEdnE/rZvetwnebTxNlUnH+Zadc8Tc5XiReT2a
q5f+3di8KDdGXjz9sWzua9Wx1P4yR6GFhfpcFSUYXxf3+/6lwzn6B+OFZVZiHqg7L/GL3VSkSMN4
eVO9y4oY/eEwOkRfktdwCHqR+MqNMovTnmxelsPgan3POsazN4aGw4QN69LsXuSYxjFVF39IPku5
9RofWxYDnqxrNuY3abkUOm6/Z1aw3DW6DKp18MfjPI4EJ+ndIJ3MNpXcDIID7tuXD4cT0ESx+DPb
+PzYA6TIYk3b5KTthyztgLDdWSzuPyB3a0XY01xX7vVVVvv51Uyd0D+tsJ9FvgAyC48fs8s4cMTL
vOL3nsmCixge6QSHQamyS9a841QsocBwtWahuVvct9Ti8jf9riYg/ataKcs3dbjPmBtfBtRvv2yQ
TttNJaDTbEqk+hoTUybxPeIB1xFbjnrkzVXu0SPmcBIMmuSBTO1Dm52mLZD94BL5gjVhhvFq1hKI
Hqw2cdfwFwYV8iz6DJx++3HmnhfafgCDnedbVlpqvgQHazD76aB4gmH3lnl1xNnBXz5r2PZIcQR6
5B4gfHLYVHtrG/f9Kmj4hSqEFcGijRug9bgMeLSaVDV0O8P5FsqcwQ0wTSFGUc05/2zMdtDbiE60
GB82ytlu9GVT2riZwZulDXtpuzKzoawgvh5zLw+RX3iZy14H9ckb0poa3P16RqLyoSu9ElNZQExc
yJU8Ed0suDL7YJZXMeRFdB4rbm1qsylp0GYVS45Ba99lMHH3o/mU+33+LR97wvYLd1amOQehb2WZ
mqZjCRj6ZqpUHcDl3GliaXtKY8juXXtBWh20ITv35Ed6xVZbCMUbZLxzb2PCIrWC83AtqgdaB6yU
3Ie1fatvPirCtHXXt0A2pnDH2OTX2nzbSngOpl4h+EYV2F3d7/0BZh3FrW+eBduDpd0k3Ia1MfTq
mKmWGXgXdpCKgcF7YFNhg0mbz0O0g3az10DSKCsrrEZMs1UURhWp1SijjGqIy6SmfLLI5Gy+VQ5e
NTiEcxy6R7bGE2Yp7OHziLMvoIZIKoNufPxuxhVMW5GUaOhb7lWsVu0ZVC77W0RlMJOAoZXJOJtZ
aGpkomxWVqLXqfZg9lG8kqBx4RpBF8TkW1P6hhWAvT3vsyNdwq09FIN+ewl5d9194L8S3fEg1Db9
XjWYmYgHWDMK2A9SMaDkR+bORqxA3mrysvt0rLV3E+/z5lNd/t1wwvchIH4llWbbxYC9SOPd4QTm
Tb4uRqj008Mu3rdhWRguPu36bFcPH4aTGCYWUI7ifkIjWH6S5xcQERR/inYtz6YhLNedMwZlLrbQ
p4kBWtsdf4nfiZndBGq9YaQ1e7eEe1eJjIshk9L7SdX9mpuPQYf0zKoL5Cg3YMftU0V+PuIS55nN
GUJBXHZyCReocOI9X1Pkccy3Yr5m5ZnHCRBFyHZ18JlNF7FQ1Og5LtoYK15lzhlwicfuUBxz+OPN
VoHrXuiyuYbjsH5Ctn+7AyhshpE+ibxPzp4tkOu2Onz2NwFjJzCePuLkoO79W/ivGB09knuNZhlw
N5khup8NNVVuF2TycFO4HeMQ39Muux0efiRMmHf3tt0sgCYZWnOm0YV6sbLc/a6jdw4/uCQHZmKU
Dx4PL70hK8ARd3y5oAnIxubkHqsJSr3JTQe8zJUt5wbusTZjKqFEynXWtpCauyv7c6yZyT5kjqaD
gIgrcyXSRQVu+fPl2Arj0L6S4JwnX/wdQjTEs3JROY8AEAifxluw2pbqff0W1kIRbC9GvUGPJHK8
LPmr/er7zO/de7PngqBYLvJzqFR6/sevzNGqOIf4RmmuDH8ZJeW5yDzfDhpJwj00qfskiBK/5zzF
w/jLxiO8EejHXGtCBleF5kltfTNggAtdvz8NJVSzPhtGgh8HA1dmb63Iw/tf3jGHLYwm8HHG9miO
YhaFfSoueMHcLg2Ca70xd+4xEqS5mQy69z1lINeoR+so4E/Ex1BHkm9Z9029Zw2RyO+WPckcDtyf
OVwZrkVPcLdNIFQkylnOQ4B6+ZlcWZ7IzpsDdwpu/0bYzRF2jFiu0TKfuDhPJCJVn+CrgGMu2D86
580DbH+AB5pl91+UJ100ysBhadchEXBR1gNeCuhvVIrkJpENwOtJ1U6mMeFLJJ/c5qIQy0qwA3zW
ZAOn6ii1zLg14F+J0duqh3FQGMJnG1eF91/e+h6Syj08DhTeenm9HkPj+BEtdmCT/bn+BbPQJXhO
GLY7yOHUfzCJAvD5vnvw7xROYMA3B5dtsGtD8GLKH8pIoSqH+j86PCYd+4EhheJ1XlqDaE+lLBaX
iIKqraRy+hvjr5EOxCcF9ObLaJX2QDYBeEs8wTS0gMdEjdl4E8SLz03k68WgtChZdodCSvBjbVhC
W7o/cSL4Rty23lWGwgY0m0ckKvDtp9Y7A5M8Xc09GI8poRgseeMkPPJ5ToYqREaY6tABNQBiw4IN
sIIWc8azz4nWdulHhmNVV9wQUkMEHiyCkNrQyXbJDE7UgXmQbR05m6t1ShfTt+JffrJ+8v3gii1z
lI/9rNKtiF6FMqkisNpAYOwhK5zNtwUFCHxV4IQUKpv+x0b8WmowU8QuYhhao7o16eHA2D+hvbZk
GixaRU3kh5rWV/5H7OVlE0Luqc6RYjE3YkP//H7wxc0mTkA3UOffsDrWULgp8hLz1YdTBYhZVvlG
nYq4/E8dgflg8qe3dG02SXspsw4tURFrhwnV/NXBPY+r3rNh35k5Gr5Y4ZtFVL30SkId4OheSnqh
0OMRTIDdF/D4BRpbye+44IFucu23wVEhBKD3R2Yaecc3xW7eJ4900BvRHOum/WyINhok8FF3p8Gb
BkeVXASS4Oxv207LQbqUTLpNRvn9hbTQekqvGMG92gLRw7Z0sKBY913yRCmRu3YLonJetCKvLxDr
ka0l2qZisud1VbqucyOt7xXVvQ0Ykd8ZVqbUb+9uIUg4Z/NOWQA1Nd1e6x8Y7zh0KX8u4dR5dcR6
JL62kECrkIR6s1p0Ns/VNF3otVrOqKitrwzz8czF2Yl50SFF4oXAcBkssHHsV2IEp1lew30+6t5u
bzyxVMJo6WXQDYKf2CqKoXdA2plpwF5OUNnp/PooUQDOELQXc+1bpR3kqz1HcQka6+khVu62i+ny
kpa2fMp7DsJx5sbsRqd6uo2PpVSihBZJO+bQ6IMQukkecSV0yNHJpEq4NW2WnfSMqWlHRC/9/xDg
k9jIUkEovRS+WBEN+EKBPIsi/ec0lMgP4nSnML/OMPkumOgNpbQXZKUE/VTGPhVPTl3UPOcd41Ap
++/i1fceC7sgLvYToB555zO5X1tGcs42KO5Q4pzQQHCOiJ6cORYNNcCb78ziGp+aB8IxDnmEZwlz
tGwWtOCsyK2RKsgU7Jp14N7RmqUYCr2echlkBwhkXY5M8j9d+SGzNEMfdrdgKnLtsehcu6uGIEl1
haOjecFJg4YcCi2qtVmLrvxkVDOpD+fCvzlHfbiH0/akeSGzE4FigS71lC+Mq4/YQgZlTocLCEjj
+cW8ZcUUqRea8pkWAiuTbhu2RBPZFiX31tGkQiO3ly3pZ7iWu634TaP4gZfUyF2OFyQASN++aAJ2
m/fx3IjiCwdvJi/v2CKE6zR6tIpz7vPeDCx+j6V7JiqgubsYYq0eFtw3+/6dvvAQoJjUREYbsCG8
0TSAHeclx4HFnslod5ezFjRA782tR82bnQwNH1qKd3NT5cW+6hfgExR8Z7PY1nnUA6/xpamc63UJ
uxr9DmaHU4tugF0bzl4ugKeUBAV+isD4FaNWeEaZjo3eRz6TdXOsCovKEdayC74686V1xfLIFbnY
n7yDTBCIJ0K2e2b2rr75cqvEsqRJ+udFRlXRsTYn3MQuC55uBKn9UVdYTCfXKv7vdvV3waAVE6ck
TQCEsafd7yjDnfTpKyW294BpUhyt6Xn+yq6ebRm8eGqI6wVmCOr9EEuI/i8w6xuzMIl0zmPnIQzf
Ddf9K9M1zUpf9KlluOarT5NoKV8mq+VKrPUf1My6Vo5zOsgkkexGw2ZoLxo5k1Rk/Vd1COa0J8gP
iBJXYLv5tDAjuBXAvS60el9dUbpieoQyetzu9Yl6yrLYt+YOLYE9iFT2iahk/VAFEGrUBzcUb+Y6
fLrhS5jXtRXOjOl7c4WuPYwyPGgGzYi8YXEuwX8wLY+Ppm8TuI+LULUXYSE8ODHPbHcVo9mafywX
Y1qCNFsOfyGQsNHCUfl/bTcazcZVLUhgNFfj5XaL2tGdKXjg8qG/tAzVWqUoS30HY+ECK1/RcLHR
5539xxzkXx7BOFQn2hw3/MHslD2RKSyaJtCRM6NgRoqkCFw/prSa0X6PXcQCsX/l8gPCIj2IQ1YN
oN8K9mhh5uPntnzNq57aXXrbtpXwVWjd2Rxh4wKy+NUqx6OSL2FeFA3Nt8G6Ly/BK4U0ejcIwD4H
LejGbeDKnefnpDgi6LBH6O5aGNa5wUF4tM8l28fOMrCwMNc700ItHUKZ6dypTDiUBxNR1OFOYl/b
T+9Th2P8e6yhwNXm5BIElvs+oW38p4m1AyvA4rJUbi+gZv4BnxRw6vGPKRoP/FHhkQIPJ78DFXt1
G2ZgSeXrQIt55Gf6TNfknhP+8oMieGSbL1J1NAfy4NZJQ9ojGvYufQJVp1n0TOIpQdfITBEgf5DB
QWmwTQWMLcOIrHeUEIMcv3u0gJoaYrjWeUQ8C0SO04pot0PaWastQxd41Lmo7VSgvKeWwqdrNmSg
/f3Mzyxip+aXAkh3CKWr0gGWfoGu1eWxj3aVV/9xtB39VJJ6q9pwUSpQEtu6hhNq0lqcMUvmzJLr
W/6Yqmf4mlo1gZANcGDrV0FiGJsj+7UdC+LB921GI1n2R4QRzcmZjT5AVKSSQYYkjWs1/AzREByD
V9fq+CZM0Y91wAOMScFuL5dsyOPzf//xzZRk3pEkQEoIzzxZgxQesQ2MofWrWVAf9pBiDux7X1wJ
VudLdK5kuBdwL0sY92eJ90STnSzGGTRqaPz/OQoQzj4hhKFrsiNQE7j0WsIG0yo5ZF5ur+DWjJ4x
cnD51bk2yJ5y2c9wHCRWrWuZ/ADaozga1skKOvPEdW9PkQLs/eOoUjd/en2RgxI79yHhsMOrGKer
h4w3N+36YDOUcz/6mMp2jxgf0jmI6S7NDbnAP/9gx4UDVkG9uEF90raQctSGTlInirnDlCsHdb6n
pF4WJjkvi0G/tsObE/XR34+vLJNtuerW2AjPmNJ/Jz6hpP9WsO1ljcHzUFQbljc78imlYFfDQsTO
eFEwSr6BrspvWL8bp9deHKjJDajlYndk82B7meV6gFOU7XaPIlLhw/ahqPQy/7SWEEyWA8eBBS/P
4k+6V0ezvTaLFBG3IUZvUoVYmCTT+N6Llh5aivLxBJjc13ZK8FKcbTYvMtAQrhau+7dXc/KfuhGY
rp4/Z/lCqMjvCuUHD45wYI30wgeIMRWN0sGvrdc78PWJd2yhyl1xGNzHTjH7wFYa59RAhWBj/W+H
G4Rj9eeIN3y4/ILigTnf3uCP/Ufcycyz6pJpcjHVBokROisYyGVrM1Ob/N9segr6Qwhnpc+/wn3t
PBH0wUh6Z25Gycq6e/B3b/08Pmav7bKoVgg2eHX8bJMiVpotfxB4VgnjDaPZg4Rzgahg07yhlBTp
HJmHb7lnMYkkxr4tw5mSO43igTXHxBHcvLgKrRD4ha854x08heWXoKVhDrfVUqF3XNvlBAzZstWG
nPRT2RTI3ui6tYU+dmUCQ9pMPv5XHwIj6ge/aQmCegkXlUYl1+PjKlGoI7DeAo9DtvWjrl5suxBc
yIKdxFg4wyy8tD6/xRrgrbwgScyJiLIW7uRCXyCYmcZl2YD1iKbIz1GIiVWHSY9ZO0YTkRzwZBhE
Re9MBXQV8sXd0ZPbxR7gGMP/oIM0WetHHQyNk5vBdTONsbbbl1S6FI9fd6u1qqFJjY5BSA3OFH0t
liumYGUuDsqcxly/JDHH9/ZVYeWQ+A3urHGHEDQ8Rflpwsgvbzhwn7Ys1oENJMtY8SheCcqp+XrO
6tiIRfHUmHcBfvonKSqJ9oA5R9mzaLckF3DLYeuj6iloI576GKog4mwUHkH+js5oOXgQvWy632Xz
uluHfgePN186YFtL+ESTQ+KnsJAFuw5XpIuEWXC27Nx5Y+U9c502+JnuYUJ9DrpE57Yzf3oTwyPL
4h8jf52NKFXjkGfw96m9qz7R1ioyRm1s6Wslpsto4BEymfGJmMVsCZ4PkHliZqw1xupBm1CRdZpl
9kSDGtgDcrwQPo0Qc4QdCEAIMvj74Bd0OvyD2uSMAry0tBWwTCFG/mtFu7GKb87SLNtGNfXWpS8U
KRFWdQScabX1I8qF1ayO1GKVaNd549xN+6j9CVE6JpJ4ucLJtayx0QTXSvPo0vWAKHjQLDWZiX9g
7K+BEN5RJW1sJMEXtlq2ARa04V1YFBrvpreu9ub7ypFexYzduEFgXFnzO+vhM3X03OH5SE7K+cKX
mGM8V9Kqq0d0h00xely42ulMYmXrT0M1ME/tfBTCa0uQvxoBmrFCtXGFlWBfNTfhi1tJ1VzMSy6e
zYHg0sncb/YA5tK5/AgOYLiq3+g+4tuVddcv0VaMRx2Uj1d0qsqyzjfcppCE/Dok7QZBR+RfgXKh
+u5RAXaRAcv8DkU68rWYeaBzJnvsOce3rWpkK0bdneqhFsWu4S7HWoYHaRQnrK7ClFkHxJ/HZlcT
rrdzvRij4nCNXGhL+uGTpQ/uww49SpY15LwCqZG40YVfuUTEbtuPtF7oCLnIRVNil7atu6lkLDBc
x3kh7JZ27cOYORFT2lGiNEoCWlGvIc1vf5ZWKbSoAFSOsvtRJjb7fTsBEhCMSmfkxz4o20V1wk7a
90dV0YokCleUxmnRhKAalHSeXUPEcxdCRCA3toVecTHIqlQF2maRBKoEYPY+4t47QYEO50rAl7sK
0vJcrTo7ZtLUqs4NcLfsB+f+IHpKKFtk6QBse0D32OzGH5RF2N6WOdHQ9w+WGt9n5FeBVLQPLWTC
0P/NLtGbuautt1IAAi4loWM9fQtC8EPinv3SuWPCGTuZ31ybeh2BC88HPeUjnGMB85YhwTRIheur
0mb7vkQDrnQPOTF/FXKIbAzL41R2pghB8V+BwLS3Ttpzfl/WPqdUI2NXBdYRb2mhPmpNPkWvtJS+
OvBxDCitkGXjhNx6BRQZgbpr2wVYvwKyaifXmpbeXeTQrTPbDo/ElqJzer57CmZ1kwKKDGWmV352
NxYwlbbSil/BPdjuAqxxVJsAqYYHj/lt7iF9y84J5lZ8jq7xNyCP3lcn2sYGwHfnOxpbNHHGm/M0
ho0Pf56zjhadlhRxvpRdkxLpEOkTsg0yr4I+iFo/kq55gxWZ+dyJshc3rRrjG4ZKz4HkMj5S+rYg
muuc7prghM11EiGX4KiQI2BU4m4rJ+UNQusT74toQCwExS1nVMs82XF0/SWXqjV9l0vzClEDb8LX
dWfQMTuJ8vmQMkzbgzCU8M8sAJDNtDjuriuowR8h0K+Gj1PL0LEfEBi0XQd537gBfjebYPYhVp8z
wQYDCMpNqXep/BdovoIu36U48rtAiUAUMg9DpSj5XZ8Kp7AUXdLUsopg5rm7nUFneGnD1DVLVVx6
Wy2qOMfZ7vi59WZH72pJHq8vbJpvsPW/Cz3OORPemVrxq8Jy+MjY/uT75JESOLhJsACcY7b+4nkE
rPyUQ8AXwakrY2QoXWbyrQ8UOmF24StldBVlZsiblf6pB1LzP7Ed0rvFgGU/ipPKZ6zBDAofLmPQ
b+F6PctmZf0GdBF0zADSbcxUGi8RtdD0BWndMu/1DJHK3Wamg/FzioQZQkc4MHgF+97hjurZ0iSq
xC5Es0NK36qzZ01fa1AFugAJIXjx69qLoMj5j7hxPyt8QpEODMWA27X1Ms1xQacPXDUXygNrnftV
reohAqAz8HmNh4H8lBWcjRCOBNyNaM6i+iVVqlduvOiU3ydMG6xz0A28zjXpuaTC3GTrqA6bpA6R
QraS2GOpN6f5O2L8ZOjabwT91W8E7BG6yswk7dODBg0kuUnJKlMnsRQnzda4TL2HspjdCYgp+oUQ
8oi+ti2jjezy5hjWMcfnMPM5ARO1iS6TqHbwvNbrWcSoIKKTXo2njPac+im1NgHrO/pbRF/XYSOb
nr7Miud1WgaRGUn5AIbAxGx3idZ1Dk2wz2r75k6DHkIHI/czLZaogm7a9tg/b/+c4gE4M86IV4er
Neram73q2uyMaWUeOEdVqdNV3tRPsb+LlLyRL5pzfdEVF/44X06txbCBvfa/bG6vakDBfTNl6xpw
A55R11YLuwq/hzeS26vHEgXFv8WbiOQY8KKUTUoZ6uSvI91FNtB9ir0t6pXSdH7AGjqtCozEXS+Z
gl5SRBuLW2gK04teH8llZHFkkytoQQcv1CEeHEytJuTX8+UdaWKY7iQDTtnXxMBSS4qxSgJsrJXA
ck6yBTJC9antweb5VioQktCkF7VAnQdPU/A8oU/UzXa1UeQ4yaNn4Svkz8ot/CD0UHTIpLPyOotv
4kRNC3dDNZ3wEdKsKsD2oxdwOv7DLfKbtVVez4oVmFcLUy8BbDA10Hy6kTHO9Soc0cuBuX5/VPj6
cpvNebawS5briY43eQYeX+9wGQR73YUouFeQG54Y6BVs9TPAEpLsdxDScW42yv7nqTQtxZSAmQ/m
u03Nky2egCED5oZDYpq7vjj7N2gQ/yp53chrEGD4XYr/8GbxERRHkPSXY9pTBpm/iRcaOVd6j7Zq
eqFT9pqMBuN8/ybHoKe6YauDwWoJ7xbO592WmDucRuGNa/ljmIPIbOlWqvxqibGECWfN64dJd2mV
/NTQsVA0gUhEx5Dp8j+6bt7shDx+vRXI5V3q+LQ8jzFrCeOiiM6ApxaasZwtVSwa75D0gXTteZ4M
ZXdNRYV+W1m+wRVA/RW9rA4/xVv7nQuDx7YamI5nurx1HoesxDx+KPugQf5lbbllANeFzdanSVwO
f1QQg4IzcmwMCWoPX4Pu9D7nZuSfquy+A59XxLu83FI36/qFIU1rdLFuAJh+iz2mSr2KI8HavgYR
pugimKuTShEEjg6SYLIyCwV+2/tCLKBIzUWB9xKqEObuNsxNGgk/eCoxQnD5W+O39IHtX8a8ZDpn
4mtRg6KhJtedgEwiwUq3tL3jkQUEzPMu9BKpKQCV4Urut8ECzKX+6KsUHadqH4PAVrTtaUTUSF1C
C7GtnPND8UdN0DLlawzElwctcGkgwnNsM1yBYk4MYtk8q09YOWBbs18FVDdSfg6+zaPbEDqS5Yh5
vFi91jReVRe22pXdjNZ5iKBARaoAPOa/tvCkgWQpWTUpYxHCiEnetEQao0M+vWTjglPpqc3OYg5o
E8ECH3pH4Dg2+z8nUUs3ouAgQoXhHQ9w7RQBpbGj40SFP5Vg0zI48hS6T5ihShdsMq4uF1XVVHH/
f5kER0kOPTcM4TIAmdXYge/eoF/A854M3jVlk7xDzwau0l1LcxClmTfQP96IkhYM6oVcbI+QG4pT
dQyGAMSzdqLwCVGBWxn6rF8t5vAgMQ1CLQaAM4K+nuVs3fMWgkxG1fTsCj6jLri/zJN1+RKvW7tP
0jSTR+quxnslxUADGljsR7gRKEyFPWJQoZ3LWMnXvdEoE8Dxwxg2eSv/aBFGGOM+EGCzv7caHiSF
RwUIwiUQrG7wIEB7a/23pNgYVVvZu/uNA9II8wHQOafG9RKewwl9f8Z+CmDd68lv3WKH5Y/qZ/XW
fy+4TOA/Vo+8SPfWtOYEmNDRpvL14LpkJPT3eSGtSO0/eH+TUj272TCbU33torlGzdYnd9GttQ51
O1KUSPtxY6p1iQFnEB7aU6HFZdI2OyDX0V8hMwyMAGWfRM9dae3wZ5HOrMJchRP0SIdTkIF4WjhG
+kJsUHhpfi29yjHCq4ISfdjAu3TEbMDziK+qB9K3lUxUTH0SVhPEH4zsde2Zhc6s2oeUor3dNqsw
spQKDkXsLe6KEEIluM41pJkPE4TDuT/6mpybImIjoYWrZXpLafTi4FqEfp/pLVhcVcyxuQcRN1Co
wudq5wg+KORMar6OJ43MfB1pvVG1L5UEpA3EJA8VxItMEHTfEUD80IWoqDITcygcw2C5k/uqe8ou
rVnhp0FwwLYeVuxLqNuTwCAhKnVfxHTSXDH6H66bEPTzh8vgGrUmHMWciJ7mvdM/GkUGpNbkgg4x
jYiIaM8x7VzGLlAWg6ix11lHFhoOKjPJHF8zy2U4POqW60W8xFt8y7Z82fwZOnvkVAoXQDJgGmVM
S9/zAoWQgNmEOmIdsO/VExASTdtc4c9tRSagUm0xo4owshHyblXbtd5vlFqrTc66SvdqEHg4b+pg
MjhA2fCIT5dwbCQlNg4G27pmLsmLAoOF9OSihKh6T4Spn+O76Wyq0dCcHJYET9mnQ0XuRNuVDgDy
utelY96m86g4UvWgPAQwOu1YAmEKUC9f5RE9R70c28NAeYCMFKg/mSDFkZ3Ho48kV4VwRlx8wlBy
soiGOzdW6SABjGLCPrMKZWlIp2C/Nm07PBIMNMxYn8eHl4EyC9m7HzeAqUO8tfzsSS7WFczqLMz0
ntYNSyGvgBwtexXKBDzWM/z3aiW/dSVrNk1UT09zkRhm5i58h4xnAs0zaPrkVemXqog4ykZPaL6i
5EgBfKEbHid6O/0z6Xmylilq3CoAuVtS/bUhYEBnA1AG4IrTxumb8Re47gjQqpQ6zmWniIvu0uiW
WCliAPfufUUModlyw+RCmzEhi/EfH6bTQZlKqqjn6XXZNOImVVdYQgtmoCAUqwY1ytxZRG+X5vlV
7raFJvauAA7AizSEa/31h9l7HAR/+BMq1hFPRJ5DfKr4hIJz2Jv8CA4dTCk9FBVBAR4/U+Db6eVf
j9agSKcj1bYIOWIj331Zs2AnS6bYp1KhDtjeXt+CT/iRhb2HMeWGbGQjiIJv+fAqrYnwLLSUi7wr
4jKUy1kWPh/BL1IL7mLd8ng+bQEhrxdEhyOTX1OfqPQ0CBLUJBHNkhN45Pn+LU5IufyL5oFmA9ED
5yyoOV4RwaCVJke7fGhH9BbcfgUy2IAi6f4k8rhamuQ5nGo0PrrCuYVXoZFLHoHT7vxBlSQ8JjNH
859KWAnCA6Fm/T6edsy+IF/VA5Kuxkk5YCOF8jmsAZl8SKRwhZuydw+LiNnizOmhNgdzcja+Fr1k
xRZucYMy4U+kB0edfk+RHYkFmsMup83kf624JCqAyVjHtU4LobriduiEgAJQQkFN223K1NgZerRT
6ynn8Jj3T00UCk6r4X9ZkbGBGBY4qlt0nj/K0p8TtznlDGAvx6SoJBWNqyU821+jzCHhtI2AUJ76
Uvh83Wc9Tonfr89Z2+Y1SEVjbnGvhNXWvGIFE+THIDtohjUH2LHbftqAGf9iDVJT77BGRiSPrNh2
g1dplNrFSzHREVjf/hU+jzRqKNaMsKDWmuwXv2+W+z5tqQXzn4mXaN1d/E+E2aGm4qezEs/2ga5J
wU6ff3s1L8eKcFJCrC4cCIztuMrRcutJTrF0Ga5UKYyMe04j1cQsboRAKw3nHec1g3hAlAypKid2
gP8cgfK2FO6H1e4LhlquHV+3Qcwf7biHeGotwNseG/79T8BOueQPbv5yamfIg8pVJc0AYHybhoFW
yWBALfGcZ1M6QwM4sAtw2APlb8Jwa4ay1+9tuxWCvaVWJMrB0lv02ThnPNb0O0l+jOcbV0OD4hK2
oQypdtL3n5FRBF+FK8Z6vUcSXAIbWl5FK1DSiR060vCGa8hL49E+8Igf6M5GHQaj/IwrHQGSpivw
lOvXpWp4Njbq/kvJKUAD9Px8NELyV35BquY4yI0U/SQVFnKtbNIwgOQdISSsjhKye1lyoferEha2
chHFCMUbWe0vIXy7hE/0Xa4M0nJdimLF5tgO4wOxFT3fUfBNw7l3WP9tJ38t+Ic5wNeFfA06yck8
miua1MZHBQwGpgiu0Fco6WXaTvgNShbZ2d8Xm5+0ob4k4hAOxDl00Z+hUFA1gaesg2MYMG7d13KL
LV1f9Q3HeatvE4CqDWdjNb9eA1AeoSkix0kaYew0Gc2vhPZsWjbzB06S4JwiVAzGtiBIKw1uwfkn
tin43dCrSCvo9mbRuE2kvL/cDKC95tB2hie1wGRHrOipSvcRHj0X0LEty4oWYrf/qlixKJQi8HVI
dHf68AKVM3rjSf/jCMtVKKHawNzaRLMg335utIKev9Cjzabeco9j69rIBPciUiNGdhjwbJDrLbWq
5JnXULGg2yiOSRv1PekNuNKl3OSmxq0FRyfy1EnYrQ8+B/2n96WjK6VTHli6DpMcvkhvbR9NGYNB
mCh49ITnzGZf2J4DDwaKQJujzPMsvQTYioseh4vQADD5IJns8HX6b0fBdAzmkSCfL2CEwMJMBNJG
deXAz6SbcqZXZ/uSQ2a2C6r9nkHG/CdTgbJh62b7W1QxPxgctk9CgTgD0Jmbd8VbOU5sP4j2JcJ1
M5w69tkvOxyidQ9k3sNDHv9J9IK7KvyQtRrStk+t7j14BAIC+cqwgoaaMtvvHGj13sxiZnEazYn1
sebBch0WUNqziteoTJQbwuP3sEEJQVVXRk9zULBAa3G3+fnham8CQIagefFNJcmI7cFiMfJNtsJi
tWGh4FDbQoyZYjZ/9Tbvx0zMb4GNFHcqvJHsfP7hiGJEFwZikZbQB05R3OPuRzk/nKzSf2LYcjlv
UFypxowiXynkI0/sVCOwqHViMYsxhtX2Y53ZZ0UmV2qpI+VQseTRlMwf+FNhpGdtC67R2GL8CNho
7vSYYOMzAvjV7zaQkHDFZGnhPBEk228x7HyW7a0OFQGgjn80e8NQF/LJSMUfq2fVoOFd8LlnrM7U
181OeTQRFZV3SQVyzPZSA9zw2MJOi0scBOgI3NPp7OEFsVpiIQ3HLa3SCck8Jk1XnSfMp13pQh9k
5MOe1g59FfOdQCbrEH1lCdehzNL0hr6kxZ7hFi/2/XvNEK6Zj0okeH2+4PCmqImmBeCdXAmnwyjl
TWL4j5knKANCk2efrf14HR0D1ZiiLPj7tsHozT+PuU+Rv6MQxGoZFnTtg4Yuv7MZweLWUjBPjuPe
8QSthTGN6MIj3d9VMUobnI8c2sNfBXzOPDBNxUqhAPtAUqzlZN2IvbAEuIpVxd0k+iSpq/os8LiU
Qfg2qgDNk8vxn7jIXiQc2jlERL9ojUhYPkcfWIcI0lKkmkq7GdhsXuwojaKDhJbuczWe+ynOI1d8
GPsAzvEjI/oazyX36SUniG9HyjjaoyZsMeCGZyjPhFjEdT1JwQSh/Yd1rxGwvSE+UrBGcDhC251n
dlGpAPZlEvNKXpy8axJaalfdSpNdq3BZgbjY270H4YcUSu7RR9ZFUlDl030A1iDmoDxz6pscMLFs
k6S8V6lXp0ktaa3wl6nZ90WV1++L2uW7B2R9IaYH7KvKjmxjwsswBxPSQ4TFF+zoLPXl6eRGVapF
CKKUYKCw0WUZXUnwXgbeMOh9Phtokw6sFP86UUbU6YwtVXoORhIxFmMbr8rdVjJzBipuHCwO4S2+
wCmf1RzDjKKQCU9HScTuJSDjOFZhVDZkKvaWq6SiFlzjx62MRbkSuIRRLthBIzgvSI4MiK1svV07
FiRzSOYDBCX+xmexis7Rq04zPaNGK4Grp+x0QOGjTgBYtWQBETfJ5zvXKUjkKQcs1KrhEULt8Qfu
5TqnpMq+8lF9yW+uXsH/AdYUb3Nu+f5+FOBS7OdXNIkw8nFGaALMjDHD8yOwCP01chjaYYG+3Pyj
LjWdqc2S/FhuQfbBh1aXNeXFKXOxr4iuBJ5Ivm+ZM7t+0kivVmOtbPOJV0yrvnx2jtjzVJ6L32ih
D4eY52QbVOviADD49Oe/d924SdLYX+fKpLEgWZcajtSstr3GeJ4FPKDECXiZ2+L+JtCkO44rszfN
X0x3Zfl4bzXY/f+vIuh4gg1ZEE1uSPmIGouT9YKCSuDk6wzdQU8cLdWCWwWDderb3GjWeRV6hpQm
VmP/GA7qZ92JeL9lmISJy0WnccPbDiJjrzIw70SYdpkldGU5LNoYacENFQEpfWYDHAXkn5dlqQ9j
71lBH3tNkuReAqg8A4MaCrSEEMFRoKCAyCCQhQhbFlu/xxlH9AkemX/dsqr4mUGQUyMJGtiiNfsB
1YruC8f93U3g6MWI6sSN0whhTNafSajMPc6WO/XqGn0fZ2tsNheIaiy5QC6XkjKOhJvSUSRApgo6
TxmIMkJAzIq9I7XmTjz84fDS/8WCGOlQdqN7Ca1fhif87TCZhI8ay2o4fvHL6+AhysofzqOKnW8p
yZKFfT2l0JCs1EoL3ho7jcAfQAI81N+KMTEhMoC5Aj2zNphfebJLMj4A7Jp+DrW6KOVmTiZ3o7fk
6IOeBOQAsnbsE/btDarH8ReRv1Du540foJW/AxA4pXJ4fI1VilNF7AUZjH0qiRVxdA2BumWen6lH
Svi7wl9HynOrNZ5fqfRTgGE5OjpKuj2vbWZsB6PMbQWdTyEnJi9iWev5sf3UhOb1JPSVwvFqyYcm
LhnYrFC8yvkClWErXjgLS9JvuLatOGWkVvBvMWpK12skGMWtpYZeKQXBNrXet0eofpWhdHcZeJHh
y4XXMXsvE7SGCdgG1UBNtBh8LjIrGHOYLrWNTFaiCniEBmrjod5qitB+X9lnPCVT73p6xcHE3xCo
zU72erl93Uw8qTSi9QlGjj022SUIE421OJXEZ/FY2LeX1+NBF+0Bdz1nXYmppPg7a5XSCkQ7e7Jw
rokDJwF5uiOFzo5TUWGPlrNpumQwK9KRT3MAXnk8vlhcoqduoiCZJuWMflk2hRwXKVror9tbQH+V
8Dpca1rAS7TViRWlNSIRhQWxrx4btHEUKddyfJ156RASKEX9dSjbbRCKx+pGQ2bQv/dgVnR2dqio
P62eG/nDmsRzwCZBwjrRP53Yd9NIZzM6SzSij33euqnmDFbXepNu6U7fVksOyMhudfDsLbDU+0Gp
FYuJ562CWf8tRj6X+ijD3umE2xoKvTQE/j32MFiXUCMs0rkl/IhPLv16DuSOup/PlPL0KKuwGn6N
/Q/A5RT5UoygjuFiQfqY1PKSs2i+tKYfEz7CoxeAMb0BNBilO0JUT708Fkul0bOdlCCfgpoDGF4G
aIMkXyaW2QgegrCnP1EOtgq01KCCJQxdkWxgij1RcaM+Q9F3fTaNvT4rguEY3Bq5iZapdST6hs2T
5BXV9f9VbBn334/2mHXM1BIx9hnEYXBWIjQkuG73lHX5bhQtfyBQTy3LFsFItLeRADMZ+nYNWcL5
4JOKMkoCfKoAzCZqevygg4bcckwLQJwnVO08MMtY3GM3WfRxUXxPW3RRm7sHA2nhmwYiljTlQZ7U
hG1ji/uFJDNazCoujKq+Gte/quRpPPN4Iq9uBEDGNwSBDLki+hjy3XujDZAcCL0CsbCCMe1fx9T0
XeqbcjdAN8xi/3N8r4w49LO6IJiOKMWNT10bgVgz6EHOncVr7g7Pb6w9aQSnvcVe/9fmofyKAoLz
2Xe6jEjljGRUq8oYCczhF5zhBM1FSsnvGtv7QB6RdYbTx5JBWeOD2zjMuiPUaFglxpJhYvua9gu9
UJVhRklrSFGCjUUckdPDBbH6MP4MbOlxW/EUnC4WgEb8mGcWqkz4DokH5I0lCdOxJUFdMMQc1bbJ
ggOIFP8ih0B65S/Zas+eXyFRWyayRRgIfPxeDm2NybPTeFTGkXFlRP/7N8uh5MTA9n41625Q5qOY
V1BbL404yq1u21g38lSDuvK9d1pNmpQI/RaCdwh1Uq1RvCXpBmAt/pcQOJYSfGPveRmevzcZiBD8
EhIch6NzAGuB3Sl3+70sTQcC8TNG70FnDxObMV2/tFTq9RGj5ItllPotjpX3q0iKSmFVIO964emd
JU+NluK+pYZH0z2odQ7islKHN/XJnyxdA30UILR1eXZBxQ54h9pAVCHJB78OwUsOmz6D6ovf+Xfk
REKOM1E0ksFkdfH4eCtFlu+/d2w574gU7/c7oVEWGuZ3zyZJTyg6LdxQTjUg1Qn4QYuRV8DC9Kkj
KKmzroOwe48DRA+qSZl4yurRgvAZJSHs6ICgJgwN1MusSCctZ4Ax9rJhpjdqyTftIqcyMz9xPhB8
oQC1Xsq5H8ywWuKQrEAFPaaoAJJLD0IQZzd9L9A4DXOR1GLMuuCRmDb5vk7fmigSCY5JEY32v0fZ
Egm0OnWJG6haStJiFVv04j8TkbxAj4fpSxLeGxiNIEHcQvjfiUl4/r+uQYZLVFugWBJn52l/rurs
fdmxjv+wV3D9wZ7coI3DB3jC7g0X8tH7yZTqVGKkJron8CppiwClhvnk6qge1HEYuUfRut+sFXlR
9wlzmBRHVYxwuQ5GtOu+N5EeLQOiHBimCY4tcPO3y1WZuhD30Hbf0+QuQ9TaVo4Jjx0aFc8YRWRX
rHp0FiWGNaVL1Br89oSodH5yrcTBfRKlDyyp3GIWPiq44/jXTSuzmG2X5uCPCh4d6mlXUYxO+Uc6
fkVFPiMi6Xr5r++UwE7sFB7+8cyyKhpkvPWNkS6Ok3bQZTiYPSOr8EpnABipYuIGlq8HH6+pQkcA
HJIwiHag8D1sUpu/QRJZnMviPNpKjTH3BP0eQOLI2oyPH4z4xFCxd2NRTcyQx03oEaOUK4+PSPoS
yNf1m5IEYB6Csz6P4w4s7Ov80BAktvNsNM8KqHqbr68CBudvLBhsCIgvpVAgipm6FqAlR0PfTeun
tVatDE6v1eUzoYWV/cWpDGsmlaUADTsf5wcfEn3I4gmLTBPnnJuCJBhqasqYTuwkEXhE5POwYdvs
7WqbN4JXBgtIOdO4EdjgVV/0ZT18Jz+lu9v4R5uETc447HKFmFufCBvCarReulQsq/CwRS1lScw0
KZAy/ZrDpb0oSg9rzsTpye3ssUDHLnyMBfTvI+XGiO/JyG3/oXqq3L9WVgsKpcqT+pGHwynymUtD
3K5kS/VdtzXLv7RmkHss8m29riThwa57sbPSYSaV69cqDMnZglbc0Sv9zO8kD1WB/zY427eJJ3SQ
5Q3Yws2GRFk1IyBtTi8E42grfvhfwymyQh15H7pF+WHd8qQ6bSSdTZcweGjo0dGIlKD37MKzWBTB
hi8HUwCW9sYuDD+FHGfKYcrAj82sYSMSoc3Xq3iv+c/Oh6TiJ+hmrMAx4PVlgKFXDkGfWufN1kzy
Sp0aos5lOwilaPHQmieZ6fUxJjV/x6So8zdjXIHyJIdHe8Ou8BPEb0eESJXddBriL13X9hntsxFt
2MT0si9eB80SN5HEwBjbI4HMOTLHOUAQiUHe2rIQ3jPXo1gOIJjr2mpxBEEiEvb0zFuCV+ojBIF2
w90j1UkY9x4Bms9ZgsoFVscT63C1xjS9JZ+5CZckLfIeOeeYa1jR8vLlcYQeQ8RUfF2eVowAYI5f
DfixNYiNTNrTBPrARS3lyEkFEe/EnEaag0qUXKKJTulVMJDCUERsAsYnpO8Vp4tJb6dgUSteawv1
bzDgkk7WR1HQN9XY6jFVqiVqe4F1PGey+lCWPi2Npp3WZJLrjF9lddBIBHwNGCcNPG0/GoiZkonn
nN7cuKEcAAFSRki7Isdj66vnxcMC2UV5/gBpvwbOD84STrA4oAdICj2AyJJPocmTgs3yJ1/Ua1vH
oRTgBLRXBzU14sUUgYduzYDlULI+UfbDscC3sv9tQb4XTTwtzvYRaPxKGowyosWxQWQ9eXHd8a/d
g0gJ6znV0z9XD1DighAB2Gtn67Apttj8dUg/GabbcRegiTrct6ttS8zPvPljKS/3Yr80up2g6M73
3w+x9bZWSmkSiqx7qnp+tS7KToIY7dlCc/BG3XuB4YKKHb13gfSyZdehn+YcCSVKuPJHpvrV28J8
QLPIQ5niOaWbiYqs9cobv5yIQsePjfa+JPl/4k9rD4mBlkMzFv6Bmyw5xeMBVMeUYieS0JHC98Vj
hrh+XFaQkWmSwyTdxhvYAmMphLNyUB2xQr3+dcFBDg5Dl5p4BfGp2SLH3fCLus3SCujGPjaaxGUM
DNi1SY0Alu7QthuE8F7thE9+kg7n49NflwYlp/zA7QvZJo9qv9lUAwrZpoHc5c2kJIOLDC5PqJrv
g6tAFEowHaHCa4gPUppTpNYYHwycTwzpzKlqXGetr1TMJC4IosSUpC3WYNFau4tODvMjGyiGkWa1
9cn2BjmVbzdou9JI97R7W1n1WTwfnaKbUxecXe/w4PT3Nxc3QXj43Q1j9FUPnvIpMNyIC/MHxLVp
1XFJy/K38zX95Zz1Z9JBdYLkZKC8KSr2XMJDL6tRQk3bgOOZVBFPbqDipjV5y+aQMYIIC9QVfCdP
P4J0xiLibm+UvgFRMoGl1APjDqoOywLIkfHefC7wPtD5rrLM0egv2ksikeQlW7bDIG6RqIG+f5ps
EuFTstIxHx6hgVeuaLb/4nSJ2Uhvl5UsRVQ/jdTfQocpo2paLVferj6hOtZhhVgOjCqm8vV2Fvqv
JhTL0HLUgtCp1paBTJMvKA8kziDlPvgJgljTlz8JnmfBkWPRsYlMpyM/rlCrZp1jpgTjXNbkfPH2
NkvHEyoSn9bCDOa+ASNBf5a4V135PrtprW3ovU9J0i+GWCK2CqcqT+mEz6pQpen29hKGbc89YZmt
AVLsq2y0IDRMs4jP9VCZ/a8mGuYfk106HZEfq/zTRkN60FJ68BPaIwRFuQzS1pfj4PqVLSYtQP7L
6m14DU4izPkdXTy/pHvT2cR3hcIMobTtmP7Oss0zLxc9nyAGQ2QHj2Crnc9/T0VCOnJg6NXy1ift
/lVW0RHqz9reIImjO47cQO8dDq7HEFWRk5LlhyJAP2+x/SSMcwajPPi+WoyKWpYJqpmWYvVOJaM7
O0AGZ8a9Qc7sFHOpZ+z40Mnlk/jlI8cW7CwNXbEMQoAUgetIaTymn+AXtNyr/iCcduTLto1NMUDd
rTOhYKK3Msd/Imgflxe5rjbbXFlICUVgEGULY2f5/dEGFeXZ0znzni23n4Rpj7FVeX6Pe97RwDyb
QtMJHmgjWJRfqVQWVKrW1GNAu3LfMflMPALPym8nvODCalreXP2TspOheJJwxPpbEKM+DWWNVK9w
zwVvYoEP3had4eI4iP2d/OCHOogM64AFfLaiBQ+fPO86rikBGbtEnlWANZKaSg+0NW+kLyqpouAl
XQuAtZcP7SkvrejxH42Qg1G7QJi4Iwmm4Pp150+TYLI5xzd8rwJB/dKjvKGL0CcJ8sYiTeFJ7EHW
FLT1EffNlPiwS3rHfnuWDerK1hncU/EmD3Ln2HmGFE67L9zuYt83i+VXSFDpsEP+PvxZ1HBgQ+fl
EzaJtakbLJnku2UuD5Ihh7NcSbZ+DqaMZU37ZV0BrKrjZ9HYz+O78jfR8bqUrOPUmVPkn8xe4eDR
6Pd9AOx0KJdNYYUqjHj3Yd4gBMZZAuzrJOEWo2jhgXnz/tKYyrp49o8GRXafSkNqazxSVvdqcdev
HSfg8ivkd0z75MjsNQ/GrwXR/BPmYxl9/DeHk/TFT6FQHMF4cRtlUJe3T29q0pqNSPP1l+h270Ch
TLJgXViWpKmTF6Qcf3cqFAh3I/rtA6aP14y0rEy8Wl1OyTF0dTEDZCmda4cZcouOlBwwAj1+GE6u
f1vDfJl9fgvipsGYviM5VI7BUXQxN8bYEMJVPq/T3mD9+D+msPhSTKCcUeVs2n6jBCI9HHd4SrZa
x8jZqL48WZHhRWelnO0edDZl8Ff3hYZ9WXwtrOTV0s5wjJvlzFW9qRcONvBArPdwj7sudZWhzPt9
EoSDK2v/Lgkf7+iG3QyKvnTfv9RP85KVyCGMhFd5QLxr6ur4ocxaFB3l77Nhcdzn7bVllbaDcVRm
OGz5zZA/J83s+zVzaQSlerylugHi88LrJYdLDTIGzeLY/2XiA4fIoGTMjHFhcL9oOErakVcwemqP
GDytl4L0VDInPdC8g/zbyntIMkHx/kPDI9DAOWJU8QCEbVtl8vRD4i3tHJJsRgP/TBATpgC2J9Sa
y2pH9J8JmnsNRY+mrskoFZoqQkcIQ6Mvbnl7NDEfX4S+dWUZcvcQ+I7WSUrtoDb3R0XbYNoEI54V
8FZCHQSbZ6s+xsO0siZLpAgfsiYNDPvjUQkxbG6wmd07as2Nqd+94uVZCLy9kXzZXLnneN8fU+Sx
ZsvCz/pOn4nF/wWx/flMauSaWh1d6KImg7Q6U7De8KfT/p6Z3M/b9ZQSPuUsFtkDwWYCrCX6QA8+
adpY7Vp2iS3AztJE2ONSPxX2R7uEyiW3oQWqx4ZcVU4GILtPkAAZKtEbEU9NhBpOHJunYDSVKF6n
oPxpYfIOyW2Hlc4RF8Oz3kL8k5uvH3sUtoJKcbxvXPpCOWVgDntAV7hRjEDdgPHpDrTFYTk9Jg5t
POtVlLVhl2X/S608HCzaP+ECRG4dIH30dWVGQdTEfIsbiWzn8vlXyVUuZTkT7G8JE+d6iuDpS0m6
lKiSXRbwymyH+LJx2lZIdPpO+nrIRcLe2SqYlVfAVfxE9gVPNOaWs3HlFtPf9GUm6HKCtaoumr80
xVOK1pgdyO+nS6enegomAV6A6amu1Io9xtYaSdrTkChjOB4trGFMMwpHyDKXCKXbCaAo/gw/2Y+A
0b6jdd02JQJncHD9f/x6b2elBAOIp+ifkEeT35gsFDoTc88DToCnWJ1X8sLKb7BsJTBnsildLQ0W
tcT5009wu3DxV05L3eX/MLujlBzDrTTYHy/rZF48kC1M9uRRkc/TAoGltCpe/67VdmpXWgKJOlDF
WEgYMeHAzdXLSgA3F/RiHC6liHaPSGZz7j3RW7+7sCKwQoZgu6Lr+0EB63/lqBX5Dr757sySmFXt
a+WmekTQn/XiRAi+FKCAdSY4HESrdd2O7b74B79Gar82tW1NctzE5P7grZjjOBRZ5hjEmK/pAsqM
rcE0qyhLwfE6eZJJSbV0iEQ/hpc7vuUk+YMJArTzHdCrZnPVMRR4D8liJIWzNEx+TO9RlzVe2WEB
onKy1sxU0bzDKRILkPCBaF14DcTsUNK8aLBeXG/RGwTnenBy5uu6+Fu4+Enq0l8MBphKnM989EZw
S5LbV82RkkREOXkpbgMPra++uDYWXZLqGJeca4V6Ota8WQvBPL+Ci4dYwo+uDzcSjHmJpnPgFoN2
70rNOBxc2Fq5pRWcu6kldyhC3SF0un+pIwIB/Ow89eWZitNpTcjAOHqsWoAt8gZ0Ug8eBN67agpH
9y/dsa0qs1IftGzmby46I2GBGuuGpRDdfIpPmTAj5xVEx5ADqMHsYUOUlmvpmDKbTywMwfvc9SNm
5QjqsFwFwH3B2AbKB4iUnaoZujxUz+8gWvlzdtPvixBHRFRwe94XKP3jzz52yvn6dumr3ED2hRj/
XfhtvYcALpP7lHUtPFrLxn/K5Ja+4JgOYHFR+J0Alh7jNTsAEMnW6wcJtuU68qjHQqGNnqMCKeDq
u5eLOcxrld/p/36Ut8i//5wtniCPJXvMJVCsot8gBiu5VjdNSystV9zHssacmUTc8SeX5F3HwSjY
VvUxTXhgpMvXJCe8IIxIk0a2rhRqXZgJLCnv32nvRRTsxYzXzsCiBTNaBqWaIYqul8tW2VXN0q/c
vlQPyH+7z8j6YI9iEZ/87nmuCdqdV9lmfRvQpzX6PLN/RlSgCItCDgcUMAJN0hP6YTU81yPW/RM0
thQ5Gtk4nW2f/JLui23W4124RY+8jjUzkyllb3oc8abfN+R/99YIJl3wYekb1Av+BxtRRqUJWnQn
iV+r+gAyzdASxsp7ipVoilcUDkRrEFubDkIN4CGFxzwr+WbXogQxzHD23/KCylJQPe2h9FVhg/9O
TxZ+clFWAPi9xxgFQYfhIsCDvhqT09BXbZBna1PCBTWF0R1RBEmb6p3BhlMqhnCzPyecCMWLwKAa
Rs2tov6+cGGuwKw10XQkh/jEzA8l0Rq1SkcTHD7HChuMffueM4mHb+JYpo42pXAG2x1GuucJrSLW
+ariwt0hwAxkepTD8PmlqXszEqd6cVtzaLXV0QiIsUlTyu7y3dXIY8I4YVIfj7NkQM6md6J2EDhg
NaZ7V4QpNW4ycDYk18KfIfZgWxRxsOpF0toGgWISTrUUMbmOHnR9oRglebsdrUcyeEsaiNSFafS8
Lvz+EHOZ+9rvvWY0SQ/johW3RVMTCa5ZbHLFFYF5tw/xSeJ8VGY6kQlOHUfMrUwAOPN7fvYt306w
wAI/esXVQ6cuswb4aq3fKixVacO7Kkqb97qEF9GZkdSqzLE8+z9CRi4a9iHWcL7hPpeYMFdYnnGh
z/ncGaaKrXWNfbV7AA1ww7zPH0w/xvd0jX7j7I582WI6Ul/ED0Z5mSsXk9sdrSStEH5DxayV4RQy
gT8epoMGguaEIzPN9mp5pJAVCYxRXLozsGRN43yRwy1EgCjQk3IzQp/oBF61y7uDs78EuHi1uuqk
jgBjfaB8skdbhRfBi4/GxgY6mZMOYNH9RdVlcXJ9teyObdGVUWE9ZruK3yRregOzM/ORyliPgM6P
gQ/xUGBGBJlqhwAgYRrKJ7OFKm+q2oJmrK9Dj3O2cTC2qwtF6vyvJNumU9HX5RpoQQbH6HvU0t3+
xi/vku7VvmKxpaTs+FAXAjracUST5Uids7RL2H9A3FdGIlIc7G9moI+0mARiZ+T5qPlowj62JAfi
E9ATGPqqd05OyugKfumav6UQ7OrNSeNR+jpfFzfc0mSINiHwAuHjN6FSh6823THR/gz1krdNKyY2
ID7oMt12dUjdGUTlZruA7iKJHbJjQMgLb6ABtoKiWEzOs4EDirqG+i4DJYZkkGrLXlNS/JBoGJE/
EoNoECefZXFOZKV9IpdHSv1ueA31r0EcijP/Mm2xtTHHGLJLLVzGuWjxIL+OQs5lzLghg716k62h
UOs5bj+ridr/zbgtgeO5ZOlJpPXQSqgR8I89rnrkAhMLHfXSVe4NrkhKxiEfvWTWXyBbRX10Tve+
snEsMTwPJNDIllKZYYPCmFqax1qyz+Fx3Q1cseQ12xP+HmtXtpf5Q9Il4L3tmCdhUDd+Ccj29LgJ
4ou3hTfXGHadaFmf4c+4iRXeqKTQu8Vb0zhidAhxCzTjnLPOgOfe9IDK+4bBWb5v5ugFxlF6rKyi
LGJgrBHbiAB19ZGlilCEKUjbrUNn6n6E7LEwgKGOO2x62KZZiUx79ixrzIl4I8OV2uxK8Pf77ppb
6S7Eg/o5uhIGBqO1LA+RTbvrysVuRX8wz9L04SzXXSxPKT9aScWJx0XwxCYXGOnQZYeXqcnht/ow
NqZ9B0lgVedDIFJ3YBZirjjKd7mI56yLuetW9veLk2k0InNH3SmmAneUzq8QJBU0z9xfifvRVQN8
cdI2YWfUfZsExlFY8NecDRclOxvr4IdVUFU7NaFrRyhnJl7T3THSrILzo1/zaV3dWmJm6RoKRl0a
TgwRzpPbf7I9nUULm1VOzFxOzSQJpDvYgCn29LuHiD7iBEJ2LQ03eK71TS0bVUCX7uWfx86I8i9p
DfsQKYfFUTTTeNhaNUZCuW8SU+5LwiSPqtGdvQWkDe/pYA9Ar5sfCd7Ac+fPryv29s30MhbxqyED
hHdwcBcxVSPM0CrEI//Dww6ZiqHqKuys8d0TOet8vaOWoV9Kq0XZErlGAAC+TmMO/ZlSiI11uWWa
d8xou+s3/RqY9TMeJHRHfoiZIoetcVWkXbvH31utRJ+Rl8CYgnSVK2SgttdXu8KtJl3p9V//p6gu
E9tr+r0+P2lXdt9W5ZCxyAyV9M7KLewEWXPwtcTcYEeg6KQYYLIxH/Rflf00v4pYBdhG0mvsfja7
aM9XjKRgqsxeenSVayMuAshYSjEtyKdWit5JzVOd7do8dMSiYcuHg0Cv+Cz+vWsiKSC0kZpY4DvQ
eLx+A1vCNyfDn2mXpCmv+lhjYABX9WWG/CQIn6JzTGgQQvmWgf9XMMuiYTQk1rsldEp575zleR3H
tljR/axUsfdzc118O3/h5JX06aO6cfCy1JXVXFKoZi0cG0OCqtIMWI7KawkIXBQIklW/cT8BGupK
k9uhqsQeC7z6TRn1geYMHUjJaCXNEItQIZiXzWSzevNbTdCM1PDkDTEYeELoktZYXraQjZgj9lUj
hWrBt2Wcm3RUOA8Su3uJnHPDTopQgX4k9q448Yfgtd27gjYG+6UEXhEBg4odPyRG8CoaxY4PjzAp
x5Gqd2hsGWrG2XLlWRESflvsH8JGD5iBLuu5qkjjaVKJRdQXS/KuNL+eDuahWRkGsZHCerpWMWDJ
WCjljDZGsQ24EUwGa6oJ5kafzg280WqzfyrIaBxfLHBy4LhDE9a+VnBPKDXvD4PVVx6NR4oa+pl6
wSbhm+ZaDGFbbz/ar3heZBADI8/BUTYPnNi+MuCE6sui1zpPV/LWVd+Gtml6Bpmz9j6QQuDOAt1i
f0zQ281Em1OrKTJxypC/Pc7/IkF1sqryTEcfnh3AlTg/72E+zu6ydz5RfzpnfUG5M/aqazW3qrf8
Zz1LDlltOr1U8BgfWOuRGFbSURmbcew8YnayZ1JButs4QXp1v4g6l+EY3wV9X8u5DCTuPqmZwnDv
GyhnEOW4gGCVbxOSRK5SVGEtNoyUuBpZWxo3rx+bGPUlJjYtVANjixwZLzQvza9qVwcPdszOhMAz
vezJJo1cKWEKbdtAbjX2fGi7AJkKYZB2Z5uMrET0uIz3YUYl1bQQUWyrnCKT1LW9v+PROUTnCT0I
1sLHyizfCQSc+sUC4hBww5lj7E01hpvlvaQb9tXeoAPNHQizK04MZOatfNIk+/Pg+/wG1MKi8T34
XZaxRQOsn4W3eqGpc9Ku4vZza9JtdpEifPsv8h3ThuTTO1YgrwPi2JLfMCfcFhFnmToRQhopRcLa
c40oyAes/4CzdbGXM9k4PEceNp4DfkiZ7HBn8zNJEaVqbtywqE/nqUhnm6gj2S60Iag0kxrVgkmP
xwOHz+Dg3ThAiMnbNbnPYscb8iktaoQEOp+0TP72fV0MOxeDxBB3IONxFLJPN7pxNc5gWesDAJw8
jN5XVWp+/jQvtoEclepV1W3sL1HXC60SkBIjByffUpa5Y44W7JzyUSTv+qU4qbrD32yYijwEBuIl
+ytemBj+Aml9OQLOsGOf0qpQtVMZsrZ5d1OOx9N862t/mVKkdlcwl0+27cdwpfUaBxQvGIfvUbJ+
Gh3z+Fjo4BIirthnSuR+VlxdEaEYj5YscgvjnjBU0vLo5B3yAIiA8X2m/rlc6kfOpee5ZQ6ScrOe
ymXcaYb0Dg2gJ42TmGNUb5NoyG1ieO5gc7muDXoNuzT8WId4gOVJHL0gMMibqJW6jKCmYg+kpAAG
ulCWrnYw94zT1LfIRuSoEbK4NLB7pmhJbdzjSI8f0x40q9ncJRNJVx2anconIxf3+9NkzhwO1+ST
mYFsURVRgdpvE3n/sAuxB6h9sftPvSs2qlwhJ1E7tbCJNc2YwRYLXT/crfwvBUw7Qd8WWv5QA0X9
hVVl+W4aRP/8kG4IdX6QZb+aGFaVJVys8OZKvbXGj7GqyKQPXKoeb7CSnmzPNIFAug7kVpylGMod
3S0F1rXqt/1A479MrOY8RiiuA6HCn/zsm1vHSNY9BwKCB9kWo9M2cF1YIpwco5OCWZcFKskIFqwh
gISuDCMEVQgHkoe3BGJeBCTKQarjxMfkpokjrxyCyw5sfjqrKLZCwgx0ki9hDR7zgsdI2liUoCgy
IHwAGXm3UxoU5BgRLGG7k1BhSq2gyhxJtHc+jg+AfAyyGBmqEUzR7ip5ze/AphEAOas+6dLZdXPw
KdH+bTnR06CVa9CRrTMfGGaDXx1eMCWp17kkMrWUU6XOSJB+ruAN+h/QdVYuPOKQWApo1e8auvz2
sGSMluxpnBcfLK+EPDvHgFO8e83XBbnP+CNjRcnqg2SzwG5iD1W/gQK+CVxLex2jmolb+H8EDSUu
uRMyinvu4x++SUJ5XPUWrFjudPjqDPmDDil+uFeHFnVJPQoQguI8twNYP6it7CiX/In6ZZTmQll+
NbTt1Ehun7ziNgKV7Qyi30Gp13eW+dMb/m1CoqwZ2MBNMLtILGnEZfkU5gseYGZmF+s9IP53rttC
/5FnW9YZaKFeuMmmsLUpgBZWvq5p5Cl/KUGo3ItSVR2rngurcWmFCnaVXtyWgbL5j2ICKN0Mtpk/
4KMZor81Ylki4jmfq3DnanOFlDob7LHsGphgCqwLv629/rtEBYbmbg+DI4a9fFEeSGmpFz/9LSkQ
Fz+HVPrCvNbvAl7+m9W1/js54X6Qho4v5g9onwpg1uBdb+sXnk/VdJlPkM6WKt6BKDqfurScU6lM
lnyZoy4KFqbbBd7f5o672Sy2Lk3wWJ3dYSs7DfMzT/k2bUVeK0th8yqjdjWDCvP49A+IRF1aeFuw
DcBR9xKj3mivR6buiNLhwIv9RQxgy2o2HSTtfkuuQAOnfxvEDvoO+xHiNUc+UVaWRy8zMNHY4zTb
F8cNY5XcSusUT+9A/UTbxc4d4FpC4AYUz23lAer7bI1CayvH7aLLEguhThSuCmbOGCpU2CxLciIp
7lCWF3de3TpGE8ISjCVN8/sGdPFS/0HlyyaMN8CrlF4/8UrUJTN+owklio0g5VhDsk5eKK3FjFfS
oryAWHteeF8sngPEP56RkBlhaUnaVG/0+2cXlUl8ipdoOlXufpBWYi3/j696ZmgtP8hwAMo0wwX8
vSqv6HZGFKa0gzGYUctXc38TjG0mFbnG9BigiDNlC8Xex+P6eWg3iEqJqXt+7He8K4dWVvPYbt3I
y8+8Gst85ZfFqmSx25Grrhr8dbJDEXGbZIQq0LB4WHfA0mvuAFUa1CCRBOqjg3KGYi/vGyUYxySI
lfsfmIe3H/3ZH3JrVSF9f57BOLKXieInUDu/1Nq41ZLGvwZjpxoIoOsc/CkmX+Nn7CFRGV9zL67L
KpAB5gSq/yVIxMr0A6OCQsiHCYv/8sxoRbXO4D2+OtWBPdBp61gCO2XOuo/e/RWTQ8BVVY22JSUa
QkE+UyLiEVuTz+jFaV3/XqViCt3cRTfOpmB2B7aIOnhEQKvnTGw8PHDLetZ8BOI9igkzB8qC3QAb
UUWOA1x7GOq1iXRzR7lvqkt5RyfhnExm1GdHckDerPFU/tG6+pM95TOhNfXxpSwn40oh/qHsqrXY
2O5P/NUtVGBYhnRNm+2G7DV825CLbnsuSbKSSqxW9i4xHx7lqH9oo54xl/Wy5KxKCpo3FR8Ujxg3
Qr1h1is9g9UsAt8l5iGHR6yApai2O7/0jsCdftAp50efaL3ic0ydjrXbofCiPu2K50UcGI3/orIF
STDSwZiYlx8iy/94HVed9EDwvgbg8kyo58jTJrg8Ey0AVBryA6l+85pKrPBHAFKPxs184geb8wpE
vLzmeuh3Iwrfyyw12THG4BLLYkdny9iArGol+QM5fp0LXJXLa07UADUaW9QUPh8IjjtyCUeWtEoD
L6MA94I5sy2GW+wN/xFlUJeWTKUaMZ1bYomHOACz2i2QLJrGPFEUt6sb21e3pKoHL6CRqnHFSVLc
XuzcFsgtNLEWUudTfThMG2Z5esf8/N9gHZeb+kNMiiyIooK9R6WMKzskLfgwL45EGlehfhqwmJ6I
sCipWsknKf8cuC8KdKNfhTBNgcqEbYxqJZ+R5PIlNoKULFlUhqGMZp/ZbPOqI2rLV6fcCq4GUdfl
21noUWL+ZSYtZ+5m942qG5FnpUxtBkktlsSjeQBMol4fB5/gws2r7tdaLtoK0NjfXC0RVeouttLu
z4XxYS+rUd2vb0bbVccZcv1GRv/9Yh7PLmBNQT+h9ltfykiM7Q5fLOXEB1yQLNcb46L71eKLlGXD
n79egsodGRwwtlCXg+lw/CvHKdysi03UwgpLAhPq38XNp784onw4qk50oQuirvSfBYcdZDzcnLc0
z05RhULZqbRwZIddnvHGbJSXHZhbwQ7LHsPYXo+aB7STWv0OvWkxol5Sd6m/hSNC1ilTJ23tb9FJ
EOnkmTh0rQngxkD3dLv3jGyUBCtYfNZE3/iKG/766ggZt4wOTlKKpcOhn+s35bsrQkEoFPw+Kjko
fVchtUqOqaTAQToQWySXqLjnykF9rivCH2SQA9VsGZ49kdKRmo/pnbaIf2sfbLA6qbY0l07kF2ih
O6M9o1ec6Z40Yw0tTm+Aw6Wqq8c2n703qJqyt7bXqaMPyR2Ig8GHtxZ+f9VIjMP5V6SdABflzQZK
Lfw6x+1fF/8Qd4ewkGzL0TVsteI20lYJvNlLEXbvJkfU/2t7xT2V7et/tVeqh6b7HnwZXtwjruuu
DvG8kdNIwcg0tE12fFPPFHPrdpbrJAiwLzvqU3OgR5l7C9JjUR6iXKwBBKJTD4Po4BUC/B/deaLn
PIama9wHDadBJBeMdyHNlQkh3SZXX3okqnFKcHHiYbLxPu0HIeiTadKj8fRxxUxJMY9nrVs2E5wO
mfUJKRj13bGYB+JQvzgrootLAgpgD/i8q5QkmohtFIWykL9osbG/ysuHrqHRZe0Y+m5/2IwlZduJ
HSB/M66cugF+oIoQ+tDIzpovTUi2+rORn+upyVffSlolwOqgpKtWMTrieJt39jp2/fOYrE5kAmeu
kpL7OAeZuWwU4gkMWUZQkzqy3mihVH6TZakP2vFr3Ey7UyrHgctCySMUToNBp4N4fUwAIFy1cJYS
+twfcsQ5uj5seEPPFJ5m6HC5qkWpGZjOLxIWUX3KJLr4Hk2HuDc61G8Ru4sC0z55kSnR7tOxsQm8
d8H/hEntHl0HKn/44tT2pz5msAWWxAepYF/5QEPg33cMN+I2jxTuCEm5Z1b7TlZzW97TyXIlDXS3
a4ZckLW6grjx7fiiI1eKP8c1PeiFDpKyqaTAz8PnKcuz46rDElxTfEBfBXOnMqCVqNNs9Oqk/lGu
j1d0hF0JtvaK4cnLk0ef6Y96LFtZiQ4NhkYlnpc8PXrHWTXP/vgR46RdQfq0k5ZMS5eCJPty4Ews
gKVzj5meJbARExpps/8AXXUhhwTueFxLumgWlG+AjZx4ssLxA8K2w8C8Fvo982HLolJReu+FThjK
S7tWWmRr+2vRRoOxeVdf3TEPgqFDQDdq6sYOe5agDoOpHTcRCRIECKSIdzuTo/pcjZwyqhCIn8Cu
+xP1cJ85bRq/tLjZQqxnmGGFXsK5a3HqIIPqxc+dIfA7XNq98XPTVn6Vy10p6QkirDyYFiyfnF6b
YFmnaHMobeyMXpePEtnQI57rKntN6ptXTOQk8oQxxHWfTrj1Iwc7Si4bw/1xxqSSK9RFYqXW4Lua
DHUS3D448mso6hbx5CRD3IN6CJmFmHeCNhO6S6Z9q4gwOAUIhPxAvASFOhQA5/o6BhknJmPSFHBu
Cm6fYvCf2g59ruHI8gejbWQ7QO/KMlSHGIs52ZwXv+JNssAwXksXkAxnVtBWMr8LaeB8I1StY23W
s6qB0pcmDIr5Kh1R9AFmkZoRovKvM8DfDEFRI9e6u3TKnk6T3X5SqVHYCHaw/aK5HTiKuFPndCij
Wc0qIzPEEMw8j53eQo+eAp95a8HIeE62etIRjne2tvNbjSqm/sMkkohe2DDrrUldDTVaYkNaZyEJ
SReoR28PfgVocViogaUvJEdYq0rg7sE4db8FGGnDYsoW/dfIlu5G1vXojiZ35MopMdArSiNqKDDz
njhVnF9pJgTbgAmFYoDojy+L4YLlS1FP80y8Zoc7KHPIfCg2a0Ex0uXX8duz4TLk/kcTt7KRm1UE
nBUYs3bSm+nbjmpZSVXaJ5DGFzBwE98js9bmXyuZrqT7z475gjh6m/h39O/2oDPDhfpaBzvKYjVy
7WMNRgnIoYLOYYkpfAZFjYAUr5xnghBP4qddWO2zt/4DMbsGctNcjsXBaTsI3J7geujEqFp/EWd4
Q4t4E+tXzynV03nJmf5+7+b4CGzD6whTb32jFB5Wy/nkXXvabiJGp33m1fnn1vxR3FV7RxsyrQhJ
E7BERb2fhUX5yni7m5+AWTWzl+Ex6O4yhyFz9LoYiM6NWE4Kc9qHWHBwrV3Zt9/TPvm0h1r7/4SQ
sNm0y/p+Z02nG6BbRJNIw+iYEAOtTnEbCdEEBwxb1y7aQRAJR61WSvTmYjXICGJM459fszoxR0FS
2yXZ7PzXCNxDlOwvh8WzPPTvdmm+TvU9vn6uvP/lcz6HC4qWDFGk6pc12jzB0PTSe0KKb9BzM0WC
k/xZvCQlWsDz5deE1F9e0WVVlUt8sRCdI12+rEITVYzEb2HFHaRlY1tKP2UwzJSD2kYQcnUpV47W
pZ8lsJdMNzC8iFF081SVs4Tnaw3tgCfTsxu0NyU25gxRFHUoltKYITNJUKc/Hu5/P0yq46WFh4e1
NImcIHRNQl33yCVg1DX25prAFEcE1qg9UG99iZsqTSwJDBxKSOqkh5IS/p+zQQ83aebWOQcrp5Fp
X1qjPMv9ZLUWKRMEfhM5NcREbGVPSjkCih7+oS3xe3NVQHcb9IO6dp1IdY3JZ4QIZHl/p79aZNVh
WG6XqUas3uQRy6ffnzgkEDLE0vWelKEHhXs778onUj/MH6KwOJsE3KB5im+MPfDFc4weDY5rCp4D
Af4WuzSWQGUoFY9ZfVdZ8f7RkJ7uY1zUi894AQQ4sllRPwGYrTQr0tyJyDpOazy+WWASBsU0bFqk
LolCfsyYr3dySEb1nlIEoq7xmnXtV6UyfUH2IYkMqMw2a2my23DRTnwQy8Zsv632KrOLBg1FLz/s
bLILQyXBSy9Due7LyafG1sehvsJKcExhddiw1wIwuwJfhyHYwLhOwZ/gElbLE/qWlfQx868+u8lh
vbJUWODXDa2YsUu+dlM4yR8X5CzmX2SuOKcpqjPC1UQz/YDIRQoll2N0d5//OWxa2yt88ELaGKAy
36dbHBdJeDj0LLXfcj3gLiygWCgRJ5NnMCaM3Pu+qZ4/BOILpSkW+2tmoS+077ooFWwd9ADDC4GW
iciqbm2PZq44RYUPEhwO2QXC8cM7QWKevM9Q81+wvNv44x041Xc/UwHH5s4sfcekc3BTUrj3rzlf
X25xOvN6x29juxVgSl+/nY0E93pqDiJZ2JhCa3YJ7bvLK5jftlD4TPJqlyXpSzIGs+fdZoBPl2TY
HESV6SLZZottsMFhmjFuIHNsaCQPnLSe8znld3KWCngYAn/DwuZvgg29QSaAvzoe7dk8Ivuajw0p
TCoq/fajA+4fSpBNEvDldjWqGDuSIpP8u09qn+uahl5NdQgrMU8fomGKMuNAhCqYLsLMAAdap7jj
j2jtKj1fK2WXm4gpU8cSeVHXEUCUhoRfdW7l3trfarQj5K6fx5sLEQe/qxyqD9DFbrF4CIP3gBzU
W1dV4WfPhcnb3H5gjO2+Y8jmT3WqEAmYVOx0K54Etam6obToNVISapPz6J8fi35j1QOF0H/bIQCx
asd4tVZJN6W5pjJvdhkvlKgYfeV7gATaQakva/kIM4ZU7LMndQqxsYVHR9oUag6IODvolshXnwnF
1twUBkX3KwOfNq6CxU2uHi7zdrNMDREprSLL2UfsyK85sDZOamyW4JeruNtoPKVseEHpVCWEh3JC
pDD4JRBq/NBtn8aFxgvSm3zA+PKBYh01rakhDpluvVXE9gKTsLy9WIoVP+jDOMrp9FSqmRqGlRBB
AVSxOjcnl6lD42hFdcS0Vy7GNfmjARSz0KK98jerQ/Qd3xC4cLiGYH8Ec2jujliGdSWHU3t8FUuY
syzZUuHe8OSIie2FbxzDk8MCpaRQ7xCMh4UmeyGGTt+w6q426d3599OPBfL2QJRzo43JandNZ9Rq
VuBdSZyBkqroa+TE/U6zy0dREbKF5nnm2iHDBWCYfgo8rBZ9t5rS0ONrtDoJUa3E7GbOUXIQp0Ny
Y/J8KS5rfy4K9ISs622Jn6gLAUPnm62gE9qQR94JNsVLNTHA7O8xzpVZf6mRs8uadgBYqmMKMQQ9
JjJUW4cBLWGGE/iqYEPJDvU3aVXUWGJVMngXw+l8ce5Qqmwm+jQXc61qoWD/uxgfCHvd3/vnbbHX
hEwmnItAaT/VctN7shaLoYDgkk2cJovkOt35y4UrtqrvAMyHoYOy/VmcwgzBGX5++a30jzFCUoeR
qFGBFYmfCfF5lxoqL03Qtaace+wZzIoM9ob4swTfagXcw5k30PquV1hvcbENu7bTjDfjz4fijnSW
jLaDgVWA6BkvBuXhyZBDFeW6ka5/EY2K+RXf1rjMbcEy0W6usHuyiUWtI1NNlHUoInNoaMVouzOK
jPwgFnFLxdmG0ubG/sZ6L+FR3MnUzzGXkZtT5Y1TnvoeDCklEU/xKWoiUTjP85o8Q6pLNQ/D5miN
9TwT0Xf2HD8pBhC+EHsSgpmAIVamltG9oYxftlzwd/LsP6hQZR2joQ3vrfNKn1l6/O+/6doNDlzu
oj2X7adX4oV5BkHVvv3PICFQGHpwKZiK7cfo7Lccr3V488ksF8NWdVk0X1+FiJjTfjtVSkIh0Iid
wELrL7f/glHqQBSgLLSt4SXX0uNoCu7Ryx5EIAaIxobJvxABIEckVOvFM8LR+bVzR7tkqCdXhgEZ
aXhZaxQeV0yluR4mm5n4K9Lsw/MzCd6ZDvGV0HJzVsaIpmcjUHqLmnzXwHXXFtTdK9OXqmmVzej+
sMyDdJ2ajjzT58ricLSCGl61zVYv6eaBcHRvMfF9074r7B5fWtmqOW+/U0ou0kDDheSiGddMmTTp
2UcVmES+u4GAvS3bTbLpSYR+glclB/qYZ7tlP7K4y2JRFHAXb/m6uRJyGMkC+l0oC7XaWRowNjWL
gxld4nplyRmqpLWxYEuKBhHx8a4ujOqCs6sq+kl4R/FW8SLLv7nvZybbY2QF+LE+vNjsV1nBx+NU
sfcuxttN7BFAsWa2YR2tF3UsOUHyG5EmfS0htXpmwZ/3M0vkIMSHsIQZPBS7Vn/QMRcWWa0/abDt
UYFfANd9U36S1s4GG3yX9K8TFW3dc7TeRCWjXuZx6m3+84reFTNj0ToMIGhqjPyT8yzVtkmv04VV
khS0EAAdbmr0vgXvghixtou0xEybqaO9y4VMmtkbVJSEXSyzjJ9b5WRlwyNBZba0tJiRRhrtXv3u
SoMybuLW91/jQcT8Y2H8dTMLe/MC6CPJiCR8z9TGg69vXLrBB0KqE9+krpanLvSCWJ+eigJdml9Z
mMhZMLbeAvfmvLP9rkzBW/m/ARhvqeY/TdGd8HExC4VKoUZL1ZP4RYuQlmu2JbiyGnuakuRoVkWP
WQxQxk2RawgwDZKzCLk5GHQbfCA5EwwtKzF9yf4WvzxFDZBucESVYkeEwbS+Wzr+30umfZJDfRO1
WbRjau7BYiPuOYjgROLP61EQbdQz120X3qoOCK0rkIqR+IUKYc59yZjIL8fzF70mKhfdTNrlymgR
QG2YKlwS5LHBjUcn7/8Q3rP8PPveVfaBdh7gQNwi5cmUUI9xDaTsRXiS+W1VoTml7X3oz4EuWzyj
mwGM7vOEuNJtbaNext/7oMmUtKxZkykErPHXNdOLZ1JR9e4WuveRlKXmgi/ikwo6yQafYlTF7b+f
4qCuXCQffNuX6Z8pkdE5mo96cwAAHuWHI7dqiqY9bBpos2wHWM/28sw0qvqRZ3GnUz5lYqd4+FFN
aGAGsM6c5lJde4VbPa6c+Z1IJ1Fx8THP3p2fj9G8wKMvbnmI4xKNUk7XXRIxxbpYLpSe0gYymlL5
Tu3SCfuWHHtN8C4lTPe6fCrflpMPN6u89V8MC+LTqrvnlzI398KhhcBISaCVmIgRlzKg/OUfGxGv
rUfI+oGg6HdXZeh3bL0HqJvldCYMfJe5b8dDtKzbjwxVOeevGMt+r1WtliL2TGK068vpdpJ88bW1
+wfiHebZfEj44xIewegE/2Krg2YbnXiwAT0Tp2lEaRxz1zZyBMFeUGlHEUzkjtfTkzlNHH3nPU5k
SrgrPxtAV6+YcxNZrJXIxq7Gt/j46HdSTPSDBnbpW2a4uz68Zb+IyEnabFypr8pR/Rgo1dqtR5nH
QawS8ydi55mUV8AU4ouHpi+R1NXOGAbYvR4DvNj8mSsvYaX/qmUMbfmAO7h7ixd7YIcoA5zknzOG
bOrtKPBmUZNMVdIVpM4xube+pbiUKS2YaLox525bESVsVk//Tcymb8iL2em8GJ79iXPLBktlpvRc
ggKiN4OZrbMQf+1eBTHOWy9U2ldAbiZpKKBXNp6FZDxfjQKfR1lxmjRr7lb9ml/t8hhr5ih5flRX
ZQ1vIXCfDX4TujJocWt5+g56PztjdrlLqp9Bm1UCUCAWxOCFpDDJ+hAE6U5u1c0yASe/NXx38f9S
by5ZxbCDSfJhvLlfjycoTropJbARt8MovRTMYqyYRd6ZwXTsG4qNYrAjdaOEPBKcTqmWoi6pDr15
hbVh10MgXM+QsPK4E8acIE6xH98Gby5buAzIeTjOwkRs+7sD5UnF4tkX5LoPLcgz8h15uf8Mszas
T5n5X4chT00OGZOALa3+Yc7LrKibOVZ6KAjmOIX12jGa1ykZqrVjF231viOknOCFwSPdkzfWzaWX
SF0qLabLSFqoKqVnetoeCDR+ZJv9efVMByBdZsNR4f3nC1jP9y0CxlnsgRWgNe56qtp4ER/6ZStu
VzkiHcxuzaxNhRR8InFeyPSGJnfBqEEqUJUrLyh1COgkkXA4LesN2o0VNS5hYCQaWIC6vywXz/CJ
tJzWUcnavQo5WA1IaWcCLbCV2GnexM4pb8ZHTrv6s2KfmUEmakWEt2eq8UV1PWtiT2UEZZZ+Em4f
sg0r//gGIOHlnxdUxlhttlRmt0nFQkJmB5k2rXBL2/7XZvNbMT74CbVx3o7YLmVAElFM7sX4FuCq
x5w180xb7RSSexAJ4pm23A+C6Xy/0oTdRz/CKr+otZVSIthVYKbDJjKaNXO345eiOup+WbbL5mws
jf/MXvfPnMmfghkPDXr7IBAy6yqP4BG7i0WBrVMEzNaRlZ+oaTnVMBNjyZLo5MujyfxVnOUpFekL
qvCTeVjRT7m7GAwMxn4wzmCRwAWOa/o/KKQFUNQsOxcyYFRPNcR7SNRIWGm7vE6wFf88zfKCIstH
r7hRJ0ryk7GbN2bhwVV97lFylpbnBMRD+O5HMUiQ3UdrLYND+AMFCYwrXkCekd0ILbuRS31NxNTa
lxvcXXlY+Kt7OKnO/2K4k/Z40pUstZpXtLTT82Xoe8s9OW9X2ZAAUdrDsx5Qg5zEoyvMhgwdOvWJ
4EKjTZaN2JuBylqC588/wADb8v+LJ8IZj0qz6SBFCzm6spGaW0tQ6rw3TKzaeMc2dtW+Vxf1Ei56
5ZTWptnEWIAKnx5RhUpmO2++WilYfaq6wg2khehDid3lsX3m2jWfAyrz1CEjtgF3QeOY9K4QlPST
XGZDBSxJixppSwMgRSQfbZyU8KRBu7+TSq6Yl5VEC8B6uAnZxWS+sDYyE/U098etwOpp43KXFij6
TWK1DkcD8tnws3wCavc7eoJEsP5jNDs6KF63mi4gb1YTgODKNLUFaDxasGnyzEqgF+rFQvF9Fnvq
Ih+eXu0jIG5xSOrwnw3AXMfederIoSeADV5r4dLwjhVQmObVVIqRx9vXPP7uoU+xVE8cyZCh1hXd
NkiJi82s4chmOZcbH2/3+g6sD2s6rl8XZs8DNSNxk6+WNXgDKzVyVi457XRnyo6dUaLd8LZVdT7g
1axg6u4vzyUguXa4ngowIP4BR1UmYcX5VzDrx+HeYgkPFTzsqunpK3EK0rMHmppp76WdKODZExnn
2ktrbNRfEr19/ZeSpY7d4vbKJklGbGxlb5DnI8W7lUGfr7xILCJyrj1B1FwrRVsPOVXUJCmf3NDN
GuLqqI/9Ie8lpWZtnfrIjiE8c0fgwBQ5YDfQ2sNZqJRl8nKWT/ouqDQsTTkQ2SZwVFpaQRq+5AKn
W2zC4Obm/Zf8QgKB8W/rKCIxj8SX+fuD0Nf3Y2H+9t5kNtgFX1vTuHCWkGq2zplO8VXwP3Z+SXrK
2wuD5OEvU88JayXHSILlXJ9XpIOR/C4Ha3XMMM8dDDkpIaSWOunBJ54fsy4WpkhyqIJAEliA6f64
oEIj/HGwKuK0eYmRrK6HqYENSPs8w4M+hudZadALNm6UKZJ1iTPp7FxWDgtu72GUg2NRmexVGwsV
GE0LQYel1MvSq68XLn+VWBS091uojbWhy655wDemtUHqfj1dwwpDl1gL7gbEBFsUXoj5NShKr4l2
+NKNGrs+ONFnMylvozePOOB6T9kMkIVQs+O6xutBB9AS3NwPv7aGWssOorWQ3LShsGvxPS7Mmq7O
aXDlySwhIkEEsWpmo3rQYg+w2P+UG0VsdILZaps7emrAJuYJlA83XJBsEalRKonXof92Lt/DHDBT
NeOcIQOnTNBQgg8TYGDSuVBjSOLKQoqECyd0cIL2qNjvGo+LQujKM2amWQNlquPVGlOyV+lCAngd
I5MEGWFoSmjQA4Ldb/fHISi301Mo4h7Mz4/CCR9XYAUApOdr9Cs47AG2AYWuDODcIRJcvHl6FlYt
74EDawv5ciB0cuJWTcCo2IAqCrDryobye0OJY9tj2zRUVRcK3uAS0z+rWB26lEwJuovTm8Uh6MYf
H5SoclC/qver1IcVgBelbxFvCRLmT90z084WkABNULOP/AUWc2H0IWuCihAAh0TsF/RGsrAlDped
VY2raJ3rp+9AROZ60+2nfHM3kqJzKSn+OkB8SdQ5d0+pj1L79SVGcffYTnRk/Q3tGwee6dQOmq5n
1HmbHXGofSLDif4LqPS0h6BmgIVs3e7sD/lyOJBKni5hXtAHLS67KFfwN+PzJrBzhxrqctj2FQfb
LE71CTRethLVeKZLgWE1PA764822in0+iHe8Y7M6soeL17J9tCvqfIesnG8nE1kdz7hMpQ7gszRE
z4lsu7PunXascsC0oTkZPin6GPRdiI+t/j9YXYd5GMgRDV1L60H9eZz7UIRdFO7QBf7GhX5SmYv5
dyXepoBmAcdYJMO4CAJs00lIf3pm6R63rBjQ/9xeJhW30Ve+2vvIzqSCIQTw9cCmhmjV3dzmpW3B
MavkQC76mdBX1Ipd38diEVTp3lvkJ/UQGHejnldIjNWd9bmyBEDP/onGZrBDxS97n6BzqYWOjXb1
MzElnXeHuLGDtCiDeBr51fU8ah7pD5QONKJX7+LN3dACPoI24Kq5Cxn1g/aU7e6CkcQZ9+7MQ/uz
2JoRPfE6Vs1p0eWG//4xHnSw1c9GqdO+ubBv45b0o4Mfgqug3LW6knrIN88Qt05k0pTi0xIGGGwo
Sd8P2Hui7qb5tbjpMoRFLuCKbX5mUXNlwe4Wlr6x4wkxg/NYE5bQCz6CIF1j6k6J6W+OXCaV92Nf
ySRQRunbYuu/0v7r68FG4Pn1WDtj1btThp8XguXeyzTmYnTjbYEkFfExDFOMRinXs7IHS7NmjYci
R8MABmRg3c9N5tmpALDgQ2aDEfy0OXXxVlrw0O9l8hhoKD+uJsDzcST8RmMOpKjmDSmi+EoK0q22
4EdpTpdRocn6tNocK5OaAQDfb/RQOSCu0BWjm9UM55MoU0SrbhoNNtoo7rwom57oTn+yt3uRlEFS
UCSPoi3Oz6HQFsxM6ds/pNPqx5k28EMhLVmYSJryRtl7VTe9KPbmdVpYfJmy19i3ScOsttqkxwNj
8F9jtiqVv+HiuPRBO+ObCAaHboj0kHS/y2qy68qg1gSpuV9hGhcATwPbnHBvmHvuouepGFvfMXug
cpGA0cwxjO5DJw3Q0jKalh1TE+L85ZWDqFonG5MVDK/Lt5NYrqhBuXF1M98op/cOxUlfRBjFLDDt
L3/1CDaL2IcqSa/Pka+ycovpHl1NWZFWWcoCj6opH2f/D1Q5j1nT67YmSzewK2NUW+rlX8XSiq6p
yDxFmDMhZGAmg7jHkZgyBY35c9AE3Pqc7BViHHNhGcWEWO0OrxL5pVvw2zUINsRGewW8zf6Vi5ei
UuodxNkumStoILL5P5vwX99bkVTiZ/CiHfNOwrh3Hgp4GgOKC5aWwUq6P91pTqgIeaVcS3n3xYRm
vEB8i8dtbsKp2T33Alb3WyT/lQF4K/nsKNvsFTI49s57g3p4yonn9k6hrdRATB9iU50sq8h3F8+I
mV/oSI8gykVCgQ5C8tNjTTFKUe2nMY7jQiJFOUI2fhlgp+cE4IlhfzI9tbgPxDaL/MEKnQzEJkn0
N2s0WW+ygOaXFdc9Ftutf9XruRB4Y2rKUwW/9Pm+bfXbhD8qWbPOGuGFDe1twlsRfSCvS9uoftJS
LXqaPb4HxenyzL9dZJrqmLPGoG7GgRnwfJ2FYXWKcwXLjxPVBwjwt/UR/7XpUn69xGk9MGj/Xc0h
7fY+f8NIOdF3oSpndE+OFSsMfi6ni827pvycu0zte7mwTEvT+iPc1qLv8YXwfIYoYPK0HN9zuwdQ
Xx35YBqiE44YHaK6UaraCu2Ga1pAcrJtaYpFNcYHSd+K971tfb1LTQ86UgBEmUTrl6pri/GpneLA
QhjBCBvlDCPYbRz6/hEsl3Xv6ZcKlYRpX2hNRG3BB6yPGnScqyt+DXI62KAJ8IYISX6Jpafi9TXm
vRFBZcKGAwfiP/7H7O4v1f89EC8xU6ALVgXGNV6hjEaZK6r/azfR6D89STNMNPGPW3WvOYx37RBr
4txP5YDMYpwgzF7BGFAQF1/4NggF0yM+UQmrCkVdJ6y3C9O028OBELHh66SBOa3k2lhff4ifyE5S
+kF6zwvPZLA3/QkfaHRNWXBE1z6zzBOuhb9RU9W3u08lkdKMpMKdDA3qPdExyjW6uxsaRjDmBrFL
PT6TbE+i5mNEyXVM6wWQYOZwIiw3gi4ZacRVCrMQnAc/XJ4sWnvNSAIUJb+/be7LJQmes3WVD7YV
nSkMcZbWA3/r0wmJdoho0kh821mOhh5VmWvX48tG90xHXG5eyh4Xe4NhbqZMZsC8/hu96u+VKtoS
m3mavXTQ0BnYWmmb3y3TRbHUMo09c6H5NiDUrZfyonjAp1ef/n6FVx++PfHoV31fi/OTR/7tCjdK
j8RD90rSysaCPA35pxPTTex1JjFNaPJ8QIKM0KrzK4uPNYv3VBr4pvZCu9eC/T3BmjxkP4mMmijV
z8jl7oFP/f8j/boxdwlOnERSeheTnDRl1uFZ0sJQrUrB6zHSXjngxNE25Afk53Mtmi/u4f+PuGBe
uVt1yOwpjLkgUGbP9lpD01AE0NDC4ork9+SSG0f72YFzcq7WgmaS250eTVLeyHpfaKQSUW4RKFVu
cjzi1jXDqumRtdCE2BbMwZhjYnClk7rUULAryYYPdfqS3L1fPNFETD3zAjl144PlQ/2RkQZmm/JJ
otXm4NEe3tJEi1JvPoYUfE9EVlxGrTM0GK9YlQcJVI0X5HToXuVyXP8T/TRHBQtiYOrSLR5lNAiq
Kxca+aI6dONg+6l2tIW06P27e6EQWD/hUV5sycDsLrW9k1gS4mlFUu3iYxbbI+BC3C5b3vl0WS4z
nlONN93gEvj8FkKhn7eUMZBhzMeRm9uat4dylcTkyRRhkuN4dDPbv0gLH+XdVv+uJdWqUtBHN0/f
+EtQg/XprVN7k/GD1KFHVyjUjv3R+K/2H6wfD3YpzQQdcUtI6ADDqftGd+iVvKnUBsEV0YECOlon
gO71EXMV99B3Y7Al9odwQqRsPVDUJMA1yP8pURrvMN0aF/KAKz+KdUa8l/ey3hIEok4Dtg+b65Hc
ULXPimN5crZPgezxp9qCiOwwNnOpDX1SENG59+UzqH9AXAoMvEMbteIu7fJUYT4aYCiBRj8zLsry
IEaFzDjCzSHpCJEROlcNWKKTODaetb07r70okGyB34ympN8z6Zc6lt1wNX83LVhL3djk12bbgvdp
lS6/wJK0WUC43nrOIVLAfIYOKyP4dMSEJrHpxJ/wVtHip6tgJdU2xqiaC6DHspHylvlCl29/Xmsw
oECr2Z04f77OlGGlOFC+S5cQnEUqw8tqK0QI9D/iN2yO4dTIsXKUJs98eBCBdqXqDvYsw2G7xtbC
gYtTPXSceM6bCKmpSubENnW9Xl1JKCWL/dqOJjIqpy9sFIWzh1F1qSpY9x5nENFFRyrOqN/xY3DG
NJeqXBR8f+xI4Z7kmcfbIZAKXMqNu93yUALgxUgRLyDQmkPc0YQ8Oa8BLVPn+cZ0EG5cwY4pbZgA
FP5t0/as9t0fi3lerJGTKUPpC6Su4VJtU5/tbUu27weq4nNai0tqOECoRRZ0Yd1PV39bfRfpNNLX
67Uh6Ne4d33eHAc3rdw2Q0b7KhgBdxkWaeWPI6eIaeFI9GiVDQWJYAqsAowy8LInHyfP9xM6k1Zf
851sl2yJzqRSALZtfPRTa9LlFGnzHnyJoBuHOl5sc939F2PCNxZv6rlxCKvq0JCQ772dURFvpcap
FKBfb8VGnYPH7+d/Erx2rAXoxCUosnMJrZxOlFP0XIyxSAcBh0oPBMxd/2CKEJlHmXCHmcw3RdG/
5c5b9dzaH8lWk2IG3+4eDyw4Jg8EfzOP352D1ilgLKjfv+NqphrPlftvngsIiVIqy08WclFSupht
ZtqhtWR+U955ONAqFJHKy054Neo4eb8oqs0wyQe9SqUk/Q3KQvVlUeGNId///B6iSSQnB8ym0Q43
1eJDvmeB+TqJo+nOb96omSvfAko+3coumN6JugRmKO89MYdZymm8PYgUHGQcvm9q/tURe7OfgkhF
wsE2rmPAT7XOsUJPGfJe5Y8C9zJgVE05kQ2zyVdLKGMchCOhlLRH+b8K4BtRRS2pVrNo3I8QeuUm
e7vNBZr8N3HXUqYjue+ZRnp3ukDAO5fhs/+kz5H9mqft5ycLtZHAWIhExR2A5nZFqcHfZqHMO2dO
YYEPwPZOtjhHMpzQO8WSBBieEWqi3y+oQWWg32HwR3oMbFkWk89LWZv8lkJQsLayYGsUO8sY03UC
5F8w6BaJFptay+SjV+avVhZAJhHrCXeWVqjNsKMROixy6eNn9OqQ7gbC0RqgzWmK5wFkNyppJv8D
RYVPfIMXAn1wsb3VB1nGjaxtxPwUWT4htf9Ex1eQ39qVLueml6q3mph3eIGhvwoRyaQ47wE+pf9U
MACDawqMZFWKNxDdbfgWr+qerDSH5o3LqgHsRlqz3huZNFTmlNfMujYpmzv4Ae3kV5LS8rCW6Xy4
XrB0zBvdi6sG+CRXXZbRUfMCceLWyXf7MEltxXHAQvBH5bpPe165360HNp8bj6YplwyKhe9/DYvh
R5NEi8tsrYvi4K+zMsvm9Mwxuthox3vtVskgQBGI9/lwEvMcaccqRyYiw1cJtaapEIoIbC+w/xLL
fB4oj+OHIVHbakXI59GP7HnANh1mm4A2HF+ocI5q4qRk+E5oSktBZ4b4wPm9CVRpAIGqZm9BOC3j
WkvMiCdWKoDNp6jG8H/omvMtxv0hEQtmoeBfC3epJAhMAtqx2PqNVoqFwV/IAc82oJAruzwslpSd
lEazASDt2mBBtIYvhXR0gmudEU9n1z9AUz6EJ2N1KDfg0e9mWtorm9f50GF6k3nPnqL+QHjM+M/5
aio4HHiDInn/KEspmHwloDiSzGh/MoCKsmE91NsZrvv33q5d6YIEJ3OAbfYjBZzBbAZDf/2Fgjon
lJFc+u2AlnQ3XoK/QdOGQjh1RaJQXqPGjxMrOJO29YUBFe23HlzbE31z4PR0uaT1MdW/4JvS9KBh
z6/zKIC0vwD9iZTCjAuEGZ3O0rk5OXrzn6gGVGMAtO4yZBhqeWqL/nrkwr8sQUtNHqhUd+XWX6Uk
4F06HLhH5ReVmQfhwzhgdjlLpB0ZNUGWQ1ge8TcPL3KIV6batNtIv6TVb0uQfiBILVTrSzOVR440
PpTu+/7/BCuG9vdXqiTyViUF2ceO7GHAwZFbAdzuqVgP7dBT+yOsnkNyn/43F35z8U7peC9X7N2G
NaTNBZTkWChIgEV3e30F9m/8Z//tu7VgxOOCJWKouEY1Hd2Z6nO+xu5TKxMNz5ahxOtNNrlZoWCg
h+dVAyQXbyiGNo/BVoaVUfQ7mJkf5e7E10IjYQOf0IbLEVlKQeFS+hI9tzdCjODS9G8Le9eNvEFY
VxGWEGk5hgIqAi6qRSY736pg4RPvAZ4LwhDaFuWcZXzXfgH/PT4XfbJfs4UnCAT0es+qnJgOX/8k
BOYnm5ypX6YXWvvtpFCPvh+IEI/C1s+lNHTq09w+gen6rCuDo+Yt4nAxk+I1wa3vGaXGO9QZ4s3q
30eRa6JUd7bnhA7a1maxiK3l4SVZmtjXnNRnNXnYHsK2V3qbhMAVvgg426RhjySZvHPHq/sYODWT
TGVseBqjg66jWC9uIQ0AZ5uHIukBN9stiHu+bX1w48RqBHjiRPiYmZjDZuU0RyhjKEg6iiPXgES+
1XFfSK6xpZOgaQz/37GJksTcRoXGamk1k3L02bhNY33jzW0iXLHS6EAtSMzIaTlfRkObymxhZPzn
/sz2fnHYJ9DakLP62vDsziLRhIpeepW+lHFT4GBHzHjcizHpiU4glHo5n+RAFPa4PQxINFEQGT+a
+Eela8+HyIY4qocyUvZ4lPgwbI6RfzFgPHMyVOkWJElBdIJ25c2R8+KwhnZkPjhFitOWlQk916mu
b7guiuYA02eRirVgbh9nEfKhuBPQsHuSW3vmKHpyspR5Y0MTSlV00VifdCYnYUtlAUdy2sdz9bpD
YAmxMW2yH5QLDiPS0/0M+P/l0MD9KqkuSjMayFp7a+qjVEv+YW5/PiNFlWHlVrmeL561+7ehBtMX
l5M9ZSoR7HiCJ+fazB24YoEZL52s2xb3ZWMcLsox4oSBfGkoWCCRF+PEBt0IH602TXY62vhmSy2p
DcrJNhz8jB8k9yLcqkAhPPwHzzyrcENYFzERqEcp8wPQLD+RpPellty/bu/04kIAtLBZIUix+Ydx
czWn7lTN7JNIh2UjHfrvMk3q7qN8eZwlTPvlZn8Inn+L9yHyMYzQGNVc3pO4MydasDrnahGoamCZ
4wAQFe3NjRvaesyYSFbFf2V5pXUDbn0LqTe5ira2sbzXpoADGpcls0RtO/HUb60sITM7RHs0sXMv
Gu11ENAgHqKpaMiH9qDqKhRhlnTnugOXi6hA1TdY8kxujhqh57SATSV1jYl7qPT+f18YExjNkvgh
1osst5LUAkMppe99MwcBgu3TEIVQa3fHkv/7RJ0kyqEpa4J6lFYnEgsCE0PnNnQtiAq9vjc46Tn+
CYvYHsdq//UZa9s3NXL+luuoDO+hQ6mm+u6cONMzsgG11KN/PGSX5yf17L1AbmzOGe7Xz0Znc5Er
4Oj9dHCLJoksKoOtOUT4N9YC8DLIdtPEPxljndqGKp1TtLSI1gbsqOPw+R2PNehtE4O0ciKdFyYq
FXwumNEVn1JxFNeur7rcltvt3hkkC2ENWyAv/I7o1RQcM1qJX9I3kl8qF7RjiO7IE+eaO42K9ol4
RVn/7yTiurxfzOwmKUDN1RMQNouoGt9BYeAhDKXcbcd7TLtyEmLiK1nM/QD+7CItob2OwacNQnkY
Ozdba7k/ExkhuqqHQvWE8ONXXQ+7oKyNhfAJPtirmZqn5lM27ibwhvW0gC4LccBzmM6DRLJ0FKQ2
7nL6kw4zHAzWx3cEj0JniIT8sjxk6ugOWDttO8wLLx4sYPqOayCLNu5heSXJODc2VQ2hUirwI5km
3dEOTeJuNrduEK7eo1RZCjy02YfoktDayHPB8/gKM1Gn3CrHDwI7OlzXHE/7isgOt1/1ObKHDppG
doTj3cpz2bp49qqfI43i95oFLuxiWVzBIFGcKs+fIoesIQI7Mr8dgBO5TGu/O1R9wRS5yhfIlPMC
N4MgnxshIy2MXgwpCp8yrkanK9CsKQNuJzTmvK7+s8wZZKt+GhtljqPqvxyicJKEWmaWKR4RzL6a
O4cZpUrCtqLuHvHFW13oIpeHFqEpmAkbAsbCXaDdkmnlolus70rwVmhAwTMc1k/VxVver/eLFtG2
ANBEhuvzFx3KupMV2ZGzv2msFRXZ2tfM0XE3GIk8VDt63ka5OHFbY260Wkv5siQLP8U1rzhx2tZM
z4IH2lJX9J1CQMcFYWFyLTMwDrApAEpBYYSgIxKTxHPg2lkUyHMIdACOgQ1BR6XxHjcaV0gQgSfW
XGEhV15US+d6P5YqvTntQJRhlvoQaHGYKQyYLHHRHC+W1xD7vPklvKCJdYRufxCiwDemj5TxKGZ8
kNmpTJB1BVbHURzA0y7wJOsY6povoKCnWkd5qvx8lkZU4rRAgeFu/E1tY6TL5zt9/XhVODvh/Trx
iQ/wA2GZ4sC+evpo6Od7JYzR5k1M8QhsucaE0mHUnFIR2p4RDcclnY1l0g5ch+upOXo052tux7/a
DM4OIR/lFISFTPGhnOt18R6nOxUmVRMOJVL2OWwctcSg213HSb3dbKZd1hKFnIqtSu9mz8gCRXTL
BfuQli8mPl+f3b+tAOG47I+KITkVOcq/WZd/eeD8DoaHjytYuJ1VkduoN+k9NEKrIMTC1V4agC/c
OycsJ4k5LK4r5OmD0/c9doPN4mUl+Rxc0ioixBZwbQJs/TflZYzBpApyX8y8St7LigQ11ZUoQeBQ
HDf4v7tO0UKKkIq/LgtHUIbh3gymNfw8KlzIAsQOLr75qNe1Bb9x0X8SXv2L6bQBrkW7v9o2m61u
DwgzmSoF2WK8LumufyczSEl0OAS9uHSf5M+IisxENul1f8FyfJFTngQ6JJUh84e04VGjhWMmm4UB
SCvClibMlaDH9imcnFctZjQLWpmEIjlsew0Kz1TqLP4IXR9lDq6UouvcwXJioPsqY8g6IDKNyJqO
TyhHYaIm5PVZ7m9mZBdhrQ/a/ZpJrjmsB9S4kftgKjg4WstDgJqigbIcm0VptjdGFcWOSEhmSt0e
TAkh0iPor/h1daGGdNB6PKU4BlbpodwIbDY3+5FMBdOYbfIGkpfC6xpLlNEx2sMGAniwGl/IfFiV
JkkKVLEfaYDblw9yaFkCr+1ZWXKyXiGqHwRFBqvS9lJWY8u0yGiZYhFUrmFb2WcMYGyUWYCMeovn
SYtm9Kzr6JLEma/Wh9lD63zm9yflw0xcUOgtLleWHSb+PWgJCgu3NwDkqkI7PJ3KN4nZhHeeZ5QH
KCdnDWcFStmpG+KOxLS5i7yk+TurhdA1kf2653B6c0e/j6aLMBPZ3j6L0S3y6SEJBO2YiQgb/lUR
Rnjl+xBvUt3CsVoJRV7FxTM3TPx81hNJquNnBd9tcGliD1FqUB1T6mzmtSa/QayO9WSQx00ishZC
HfWbW/9QAWGN8rBtHt0wjqLpzbCvEH9DMa74LzOXMxHFjtBQ8WFOaac55UuL0GHHZCARqT2F533E
EtIaPqfUWPQEkIj4wlRsA0UJtLGfukBVIcvPxSO4nLE9Ef7bEzJGuBequh2YnKLutBg1FFj3JijV
ba85HugXqCckRBO1mz9HZ4cuPZnYHBbJrYGaYPFwLWlMOjfSAjFdCvzPd4Sp2/y4cLAiSMjIEnXV
5p6sr41TcCuUE3zuT3j4LxJfG1+Kgegh9JW2wc+fT/6hIknJRG2dwCqfEOi6IXSLEQJ4hPjynKO2
EIWQMHoTZ27/pI88Ag0LeSqndK0/+QuH9m6WVkrZaT4gqYaZ6gcQi/yjr7BiUDnIcWjrwVEQAg1/
+C5FUmVjaIoLr5rajjOnLcEEXAQoV+8vTb5qCe3HJjkeaF5DFVQrL1KNZKX4HZxzt37/ALgaxmtc
OvyJmAmGE3VBNAxSUO9LjBZfC61pWb20nzTkkN8Od0vM4GVJWPqCxgpk149wLdDQO9IcFRCWCCvq
3NhCYsfQnW3TcPg7dksOGlqOXEIC9rCDjxnpYNvncAJIVy5XayyKh73eL2vlfLr7QiytemSpLobE
MQoWezo8L1b73DUU/nXFsh+dqAY+0LEeSgEfndNMLB/8ubJ3fOdgv7nEqXzfn1GgUzlVIIksaRN4
FbmNDatv4IS2EWMRK9loaGzMSAV18a8F6bSPgt7RhAhi9aT2BT33qrbsN58zwqStOIFKZA7qwtFa
GiAAXbMAq1KdDXMhPPfPKOuFIIRV3W0MlB305vxLBeNiSoPQ/14iSVHDI1fsdanEh5ljRYPsucOe
8a5Crt93AUTYDgBX5/EcGUco0r8Wh5GvWmHjHqTkx+2oIk84tTiAlVoOjfXeeCKfPyGZBK0Mmcc/
Q3vChvj0Kj0TkMFdkJFUGtq1/qbUzNOPacoorqu2MJH/BfeMYF1T6aDe0mseYanzr7j2hGPh69KM
geWqpG/SI5r/IGQcb9pkReMH1trN0oj9a31I128dOTSdVCpZt4D/tBj+fsvD9bVy4v7SAPGaFhxp
55k+OL6rtrYFEmgHbg72h20SkYv9vre7zpRLx/JOPfPx8KIVXsry2akRzE7KFVzH+9c2iTPSY21t
LkL85aKr7IGEV56Alkcf+EpP2mfE6hOVhVJT/WwLuC8KoAMpRWKCGbHahPIoIEDXGqvEoK77uBR5
VndCOJa+h786Qq8yPWRpyhETjU8KFebG58rnlQJHCNB8GJ1v+GtXRHZmkJV51inc0VU860qD4UF7
DbzB2U0lDU8yeJ8UvPcjv93SW7TzHEyRgwd+2dgarF+rdlK6qfURyEbdaihnlEH75/ZCJ9J9QtLK
YPb1Wjv6Fpy2u8pUTxeDCApamWSWjS8EdVZ0Be3B0s7wPrnn6x+fG188DoVDjk+rU4rjEIBIB4Yd
yd19y3+BPLzEDJHj1cTEU2c6LsmxORMp4nMhjRhq5g5LGYrxgT2nY/BcDIJTnjPg7oszT7CLc8ef
P2BRL9i8n7ejBC4XrUhxD06nu8tK8RwDOZaqVDt8IPZ7sPEjOgdh87KPg8fnkMwIFUzJiu3cNVK7
QgMErff9EowPzcB07QbvklX8FUCiRKSkDSKHCi3jRxgj0nFPyGcWf7yM8Ph1Ab+RbeO7qx2nrE5R
S81/wNGRmE/7anadIP0aJrA9EDx3fn6pHNG+wyi2MoBDPrB0lM48IrMhCIcrVfbEPXV8imCLWyUY
sLO6evhLAt4uLG7Q14UAVLrdgOAMULx6WFpMslxiXMbwf6bKscbRpDV6hwZv4v6dfg26MwL91sLf
RZtaAd2oojN8tF947JJXyCFvYpUE73nrKDSmiekD2Z1ijexpGNpCXzAWFyqtMq70vxo+zDcgMcq9
IvKKbjOl4lp2iLmY8D85iBYfRQLX2gi01p/+/gyLM+eQg/IHDBgBWhS7KZYyQ6k+h2CB0ZGcnC/q
zuxES6PRo1YTKGzYhdaM9DQN/h4RWEPNT0++FqyQoVbUaC3NHF16CPPg44yMmjcKtzEle69dd/B4
4ITxr9jKJp0OQJnfDWNpOYeevGODiReGdlOQMrIOH8hZ5hzPMqz5QH39HpDcdwbVLdBwO28wILm6
p5Dk3pDGNCktuRJeoT3eRicWiQlrSnuKb2SIVrVk+EMYH8h2p7mH/TPxJLr/dMlP0tMcHAH/RQGx
e9hzUBcz4W8JP3dMsK6OaGkG9WQKmWLnzpLmW/+LTGVWeDFmX3HGILj0Wap7mBjfBn1503feoi/U
XyCt824S0zLOOQN61F7qarmCNi8hwSqp1C7TDa99jh7AR71dRa1gPgNOYG2iUX6HamwzCfDGL24H
ONZ45saN9vVUJLs6sm6s7tfv87CY0kHJYFAMBYrKeeW6P/37W2MSHx0iGrv/H9BqhNAb5Wri6z8Z
iaIXLx2kJGJwGeQajp9UuFNeQ0CR89AlBniN74OzaHvfRBpuhp5bHRVqxpwur4PxcnmR9Fw5Oyvj
IjTqPPzHWMwX9EkU2tl9VnImGtvK8CH5r1GhCYFbQj5dI0pTzh3wVcdx2g32Urj+f3urz6IOQ52s
OFOspOodCg6hCSerVDPprnE2VU683aIo7FSVGs5ewHemz5Mz1odUtS0KngWMDpNWjwB3ayDzdtIb
kaVoWUmyZWVCGMjlnQuB7gYN9FKxD+uiyJ75889si/HrMVQtNB8uiSNSadHQJ57kuWZ4ZufIV20D
lrScakJgRdY72RSNzHeEPo1lOJgfBFTQyBIfXLFoFCZodlDfzwT2YXTxxeHJBgoRkqpzY3vjdHXe
Jx6QI7AOzR5chPLny7uJuJqQr5ugWR3FUZxaiVcf2st69Xwoa3R3hgrInczCB3BTBrNNVESzhdE4
idQ+fLAmNk6LH55m422MkYZUUyVvH+64XNg4AhSDuOVPxjzT+qt6bQ5lgz1vfu3DRK2ptxXbRpa6
E02U1rk/8CSdREtLrWkD1N3teF3u1iReA9y2XanGFReakWJsk8C+0UJxM07nMyfAxj/yqApuLvYd
WJn5eWGb/udJMONkjjLYDxDujVGLLHoCszVpyQzPoZ50JeZh45gKCsYkAQ2bd1PP80UJonOKcKYq
GeiQqMguJyqL9JqVGDTCE1mF2yiUxAc/RHoejtO8wZwHKlpuZV08PfEUQiNnCusGGKHIvK7B0Ild
CcaFctWSRzFCysWGCtkyN1X7yzjLb4j5JWX+PbYTm2Z0u8RDIjU9HTIa8N9Ni9MvkSXRb3BVuqYz
iKh+Z0FA453idE6z0t1iVl9arNUYqPbUxp7bbeh37wKZxU1IVyqjlabCMazi8OrVTJB1TXoKZVrD
AVulWb8qHeBBo5l3iZbQgn1MJrLmMhdvhKYrAjXyXa04ER7UnWEHvHBC+SaJUChC6NZiZVkHOyBf
8O1a03PUDs3+cdlcOLq7rAOPeaHY1ukCFkLXxOK4Ca9v0J7PyvV8nbqA1sqSr/W+J6tNGEz+dhBR
mHeubmc3YFMGu3wKe0kLISUxOWlYtTLUFVaTKZWNH216zEFsoLSld6vr26r1ecBll7o3BW7WPPWT
y+vZwoXnk/kzytrNQez7OVlAl97lVUfpI7r7uflM6IX/stw2f3nCW4pSxNAElwoEvO9HgR+Jzl9T
pyu157dUogbLSbgvymeZ7omo/JleDcmdPZQjBwlY7Y0nq7x/cq0vsVka7kwhtfB8/6YjRjnu1Z8+
r8LA8t8bdbx5Vghm/APF4Gy2ivuWoMWntv1qt0N8v4i9WTEKk3KozeCbsRDii83FFAXCvLnqcC48
RzHxTogmmkHjoB1Ii6khK5HSAcPBj8bp3UTPE96/Uq97enHHKWBsWNShjBka2+Ftmx1HuyoXiE0a
GlR6mBql5v6pt382dmahDk1hTEvyFfpMeCmDo8U0FPHC6qJyH/cbBZHwSuvdc8q+ewKYcy8XusMo
tL7gitEpW+PBgSKP3D1LmXi/X96uFkpLCgOkheDJb/hqDPt9/k5aOaFL8gADjyi838AZ8Ejjj+Sb
gj/rhiDi3qy5MPy8biolO0Zficb9WGK/XwZG5Gfq6ULvXrgiIuWzgdUK3LN/nwTnzR2LLb2lgxO8
+ocwEs7H4EsrMHPYaSQXX4OCv/WfiWr7hjZj1jf/JrgqNUpJj66Ht5cFJxf6sm9DV7Qq8mKm3GxV
uYUJBWsNZyfv0saVgyuurXqbokoll5xdjxhHYRoq7x+n3uphAruQFnaX0+4+TryfJGscxh0yeoV0
eF7s0WigCFgGcfmxatN0WiQnzRf1kK94zZbOhcEjMb3AxYTh9leq9NscXN21FuTZIJHGPgRFHAxp
sTW+iKHZrVxgNxYAqFKQE56aiyzmxghS0766Ph/TCEkTp71PFlfEtpy0mLZegNk89C/vNP80Hm13
nv+68wJfuK29fuhy4sFb+AxBLLVZ843wX2NJLF26oO4X8qVgZQejJXl6pnt/Jv0acaniEVCharQ2
y2QoEkXy1wX72R9JoCfbWNcEKowgLrGm6kx4K+0zYV4JG2/3/g2I+EcQxBdiHFrO0AdE/Lj2bfeL
vRT1e8GvSjcL1cvMaprMiVkXOUBCMj3WIK2PZjTi0C8WqsCpgT4bPFATxyrij4Dm0Pv2Br8VoPJr
TsLHcbABRig0GGLZfelYjh45hXEoe8QaPilRJ3p35SIGuNH4QYH5lCuRzbYnR8ZSK3oWKa0MUrph
TmPyxLn4oPS8sZZp9kIyh+330b6bhTEUMwOC1WC17cjzv2h97wa22euh50Ms5lqdYU58QIbn6L/W
wo/pFh5OjC4UJHFGamrovKhv+dX55SBHi+Bd3lOFlKGYu35/zGTCbk54cXzzb4eh3DR+cNGaCHJQ
NInNJbhprhgJAfrzKkGeL7cWhOeu62wcMKlkBIH9Tl2N6GK52L1GByEbiviRIZtCO1qKXRBcl12Q
ScCrQkbc/0I28lNbQ/EAVAU76yGT4++NZehDRnv8FqkeUSkp82Veo3hcn4dFbDHL+2nGoNfz4fPk
EYrC+BJlH4V2F2Blo8KNoH0tvPkU66yTH6He0CjmjG/laKTeKbHy1966uN+piFaSB1YcL4QLswfu
BaQXRlsQ6UchcgUoOYsWQFAMTazC7o6zh+MKZ668T+dRdOcCpKXbyLaVhsVgzf4m+qkwQjH+YpFT
01rtXYHTMWvLQx5U9Iq3yUghEu6Iz142fm8JX4Q7NLaRvwquwknDX55uY+xTUp4R0ODrFUWY4k0D
1ffT2TsetTerY3LqEuYupHLl55oWtHd6VzfG47JooKNXG7P9/pDpawFO8Noq2RQMB5MeGLMV56T6
yyM37CmcEUfdPxeHSIZKVEPKhVmxDmbkykfF74OW68WFbQSJ58jCFameKVeTPa4qA2kEdjd/sM7a
ye2YiaVRVkS1A/mm5wl2S+/xsWstVWa/+/uXsZ6Gf6r3ben2ojvTCHdsdJnFk97nqK6QAdYOqB9f
M2zhgqp3sBt7JDhaz6T95bhjP5KYcRhjXEGO6qzFvX4YxUtQntD9kjxejuNdBTekeeEG0Iut0mwl
Kk8KubLJlYetnrNBYY1D0GaEoAxg0m7OWbzvJBj7lSjILxLzuFsLnlnIChjHAx2kdnMLnIkCSh6M
Qyb4xIpRFLsVlYnqYAr8+hvmnVZ0g/Bv+m/iRAlBA+wRpTUQOaub91qiH42Di5+WCWWtiilXIPb2
meA1DUNxWQaIxodqcgWEOBbh+aTcNKSxu6fDPUJWS/BiSxhN/lgQIIdA1ynMprsiZGn4vlxgPmW/
yAqV6sQ7qhq3afy4yTMx1Vq67hDywAwPlhz7JwFZwknTBGAMEXBjhd29NeqiMIJdC9Zi2ead1olh
wwUQZMU36yPb/M6FW/9OFEFNV+plEWa8uDZZfiff2wA+hs7gLYDSftMEu1yCpXtHcZSr+f2897sj
XSq0qZIAiwDZRuNl4o7nBvMYZRbAchKJRISucYVhxZJcuF3xYFlos1E1cEajkV46SuZMp6CP12qB
jazP/4SqVfVYxIcbrMSPcPOh1+9R6PVU2JGEl0cJg/pr+AIvxyi2Esk+GA8YK5tgL1NODNzikrR3
3JokHVFt7khZ44qAfjdXjxpyKJ4R+v33d4N7erKTzz06PsaxLLjShZxhWAJBlVV9VNhPUL1okZwt
oEj1jIW/V8tZourNUTofp8WNicEVNwziqVTkC0ckD9/h8EAZx2gkL8TGqnZi4AyJy6CkjvsgKvfb
CHkE5H7fMI37CirG+BHILHNlKwv9VHoLUH18ENtuUm//hC1+yDQxrtdM/fSoWgFq36+pA1uXjxVz
E5jL/C5g6Wk/lMfH+8HFdNYPHuE49iVowumFKRfadtN/PHV52Qwu9zUgtCK2c8BORYQ1PnUjYEUK
HvEmCYuYmtVIjdnP/Q0xDcIm+Y1j1HvoLzp/TfklShiqeYe9FCB6lfurDQXhKFiNeUr7iyVEQqE5
Za1Tawc2Js1qItF1PR0APgfW5HNDyFMw/aBR1MFYrJlCFaRo0aibIEoYPtv0LZ8vY4ZgMixJJhvs
rtalji4JqQz/GuU4MU1eRE/MtR3tZR1mSKCunbmJ+n059+fZoLUyt5bX6zrUcTuaMmm6dR6ghrQw
1mL2AgDv3EvDft+jlNOXa4Gf8Suxp6V2AcNOOyl2nwXbYnWzhbeq6Ee4qneT9EchehD1JQojMPeY
vQQb7CaJMwOOp3sqEkgERP1Y8GBF85B07FnnsatmemJlzw361KngR6xAn+hk7ohyzPRG0uRG3J9V
oWdUbOpLFmu6MXMy//HVQem1CrapJyGL1n0hVN7bVvfrFQuQQDcnWGOcBhyAg5vHT8YAGc5/qd32
yWUoEeRMoJCGHtxdKUpMUmdsZADb8jZx6wD/iQV+hlI90mRh5ulxfi65QGu3dyRjP8d1uwd9mJxa
ZKKcYc7M4/CTY1C6dYco2AzWKJWg0p7qymyr/SSpsQNKTzX9TNBHslvEKzQugPBP6kaL3jZRolFN
V27KFUHwnooXfWwg40i0bPaRTv/DPtIqBF6yziy7V7ob4iV4ga5D7ApPVC/COBaKVWm9RdTZ8ScS
CTdHWfHOmUYqlSHJzWnGmgN0OMmiTHq17AoTzNf1m3hKSRW7AeFzuPF2jdeEbL6U1XeZoMtmvae0
l/fJZdSpUX25RZb2BJUD4zZWcTcK9VkixV0Ex9pyO6tbagPZQZKmZbvTLPL09WeYLmF7k2V8B+OR
VaXvsHLixgc126n0f04ai9bkO7eRT0ymUOTjzxbCM/U0vmuBiS8w4OAw3xDT4WSMuaGbVwjRJk00
7SDScwEd/BVV4LA+OIj1GOyffpHBWNNLlnrn4iX7pHEJJJYNUS06oHDLdCgCFCh7HY26V4DxUrl1
o8rBJIMgnSrzJZsEm3yRwppj8FRnoVHTWhEEKpo6xXt3OsUks3CD+xStmSbDiJn0wqrY2SqMxi2u
GiRZPXi/tVX3d0bkV/GMMcJEOyIa6s3wn3ngSrfagGBwaCdwI/geh35t8YjHWEL9pb2AVoclVW6f
NXT7UCK9QQwa2/8JIdLUDMcoNfd87mbO5LwdYnNoNVmOHpAMvRQh1a+pls7lYqSkGI55NQz/t+th
lApBqEIoVC1FL+bGJrhgZP5kckR1YmW/34aFpbsQjTArvsixiJgIW9EetR7JgeXLNQbcpwsE1/n6
orc+AqUHaprL4MrHuEBGAy36KAKEXoTxe70yQkXWsJmLYjZ4SQgaYKcp9XNAUQ6WEjD2iVDBZqJM
k12FKmlZuxB9JbMhUeG4wS58RYw/78iQTjJCvU/IePLxL4FsiOHQNHtFixhYJR50tX0jcvPmLLue
/fKMYnaj2PKZKYuODt0WzQo5efQHjgsf2ac93Jd4g3hehrVX/4CcpI1xj+25mAMoV9T/P7RkZMfU
UMJ2A9BUC0su1B0rB7hnb7nGppYp0QgdC8Oix5ju03RiO/DuoW90sIACDZM6k1jIOC2DGSCGE+dR
fYtIxwcZ/YOhoOQth+FsyfQbOh03R3pD0QLpnWD3U5WntM/yUOImeN6fqlhCVXveABtXYDMOjL+i
IP9NOudw3bQDjFojXdwpj18pbLHOWlKox9A9NsaifiK1uLwvD9hDdeuzi9onv5Y4hoC16aAr3iiS
nvmcmU4lnp2yfdyhKcg96+TMw/aoYi8Hky/zjmC2MQhdabUNudZo1aWMxB+83dOMwlpCR/tEyZ5b
EYhF7l5K0S6t0uxjBFgNRYngiUkw3CrKpG/xAI4UdgBqjYzi2NOl4r4mBf0BiRzboTUbUMLoovxl
emZO++XCIOHU51c5qBL/XKydzBOoSd3NWlkwRvtZGuWuRHREhXZfK+aKDli5oBgLhMTpoxiRehwi
yCtIRY6SeNekbK+2AZrsPmzfOr3r5ikzMK64NjAjrXGZuCuyXjxdrsqsNsQJzyZ/gSXWCW8mcap1
J261EWoZuAXtNH3xwtrSCiZx3FpnWssMFmyYbsjsZTxq6Ep2LPehVK2Qtojlq+f6HYZkeb+YZWa4
ZQZXYzDTuvEb/gFi6l0cGTgTf+0n1T3h1JETeHU3U6LQiBisAD5MHGtSWfw/0i3JSbQPMtbfsuOU
2Sz1PW1uVydWp4kp91FSOPuDDIrWDr/oLjx/MkndbMXKFumdf2lUIdQQirbnXs0NchSEG3LiTKD9
oYKr+IfJ7EDdNjkhkspJUTfRxnjwzSqZf/9koHdKHSb/zZ+9jhX6nJ11HkKXi5Ki6Lf5ZAWHlJRM
3sSE4LxY2DgNNYfl5U+X7yALTHJr7K+JuE/g+/Mdz0oIfpDM4ISImQXahnfOeZvhhhJtRMlsv09P
8NhaRRbjU4O+/L3A33JVZnpoU2sTo4ZrJpbarkPVMZcR2EjjlF82DxBm6GzlkbpU2S3TuER43Gyi
T3ELEVus8rSv0VYnNZEoe+baqYDxOO01mmiZDZhZciaPBXLSXpALrLp+dVBsACrAIxDoXzi4OEwW
rdFvx4rZWRnINQg25IdEwesmKNN92jNjEcZu6kZpGqbNlb+bqZfBVctZA8LI4evt0W+PT7Bc+Zpc
9lr5tYycSMGlsgmJ6x6+M0lkA18pTnymMKa/9OznaybH1n31jTjBnqnUD3KfTcFKxZjD15Vl+55R
GBNOO9kvlSc2I9qgiphVEupJaf4Ezd8r7naEAW6RJKC1wKdb3YbyYELdw1JTGGlPEDw2iwntzpKb
OLtVHPe0rzcJo3IrEmBXN2/bKlBXpf5/yy3/8TtAN0wjulYeHAfu4xrAIo16buZJNjvLTdZ1h+bf
RcGr9jIqnsySqiFOGJcvUa+DXuwUKqKlskn7fQo5hSUQHQ43EbfFd3a07q6S5kVdcIfOU8PpAyxJ
LxVVIOI9p7Bms16Ew28n2Dm0Zha4Ofs+iHhY74/9AjXFEAAVY4rD7H+uRlPBYftX4cGH3WvQG7dr
/vhU+uvwJiNOQmBsrUmjkQpVgEPewdS8rrCwYEIPGjD7A43wJtzMS1q/q5mUHH6Cu2S8fK2NFPcM
YceGdM3P2Oj9KgwGT07Wc+SsGG4zwY/l0qq9QTbhG7larnFYWCiilNmgegla7a5h+ElwcRwYCGFC
uE3WHr0QQUXuYpf8Z5mVtpZJGeaZZoFgZonPMAezNyw+GqEBWl3SgQ271qTQvELRzm+SeCj0gP0a
bON5ereOo+WTqymnZEs0KzyNl55cxmXK7nulPubLKkeVXcSG1/c6ciQsBhfJzISmLvbLxMMOPvvc
gxmx2DHYtMONwacFbcFVXk0I5cBLMepKPeae7mARsJ4DwAc/95byTjVqg0YBRKEetYXlD6kozPm9
hpsgxrV9eE2QeQZdpXBJXbwhZdH8eGgiKrAVv3g5GJAHAgcOzHC3vEwDh4XD8tqobVZZPH1dU5oC
JMmYyL2C6GN6wzGu59r3YIWSaHrohEnm4gZZDGvJdoWwO/sHWWUuKODaYU7C9BYy24gWVznIMJmZ
gU5ZgYtKwMvTZc/XKPvwFkL4VpdDRFNBmhyd6KArmlBW8NuMcdzKLmpY6HStAWkyrWbTrM5kZTJG
Cqk7OcSR+HquI8Su6fIzshpDmOCybG+R7xNKvosNv8hhkrvup8T19VJu+0h3Gk+o9Lty8MSgBG8Y
ck5R653MS46sBYCBMTNCrDcEFwR5SLzPJx/XRkrNnosxslmfHX/gjR89XD+08/xSCRDhNzF0XVXQ
tWL/61797wLUHu8QnCQH0zC1DYgHGE80njwEjvPdB5WbCPxJHYnGZTbPUmzlT1tdf6fHzR6bxfcO
2tP2HdKq+wh7QcW6eXzkPMtZUNyyUYA9jy55CecbHHsxeOA+AsV6ViAHc0p/5d+ptMTZyRVMeXQ3
bBKFQazaW12hp9UttIjIlJAWPmYUuXn1xCJpy7azuuCjSHjaHvHWxE5qkAkZFYLOXgB5ZpEQXJvc
m6pcUwlopzTFmUKvD93UNICA+ZSPPOQ5lijdhMg4+JKnSQDSnL/ktTiCuprtKcaadYj+C5lYZzTD
/WK/bjJLoG6kLZbndIpVUzxNDI2K1p9lj1LlW8Hp6lRr8OHI+B4tdzIkcMu1rD8qKOf7CctRcKQx
y7v+V+rkOAN2XMjf8j0IqQh1d3wWvv8ORqRq3YN3gVWDscXlbry5XnDgzGAoeVY/ePUnGZhj2HD4
xBvinwOciwIY1hFjETHomoxlWFQzVuIfjkPZo8FOtlwq8VXmtNsMQFGnN6c4nS/TZgTv/VBC98q6
9nHwfZ6/U6+7vsLfT/IbB294wZXbZD9Ndwc31aXpLcK9UpWORd9idQ+7B+mXFD5eogYRKkkJZWwg
dFcc5dX9+ySVJi/aaBj/chQ29oM92jJPPXFGDD3p+R9obA0r4bGbarSQQit1PheA8xwDa6SOMKWD
tkvfa6HXSx3IvoZ12JyDvyw/bxnzlKBVraFkMyjgbNKd9xOY5/PgpLx5pFzQrW2M4113wZWImNjQ
/9pajLn0M4WQK4tQDmeWT0bZVM0/c1AQNdbHLMPDZ2qUlssMu3C9+JFJoiA6yAVZvRapqv9VkOk9
9gy1GpNqlXlbTC/HieBbzo8TR2FBrXenLJYyp/gdYqUAo9u8fTrhtDZzLSk+F2DltE6r6hUOR+Tq
qOcPqo1EGrJWMjC++Xi6POnr+sqN2AAjPr6dDDTVS6PQVzoe+c7TQyb/7+PiniAsARBZdlQZWWGZ
aPwTgebBNLEis6DU4oGAgFbCyFP7mC5XEPLNOadzg8UE+DTkzRCv8BtSF6P7d0uorM+vQookOf4I
Gh74IWPUJllXbZ7naFUiqurIVKX1ON1+lR7ft64UU2DyrOf9/yKs4O52LHRHbHZqvxHiIBmJT0Vy
X6fu/Or8Ao8MIanJl/DfsnK8+NLiK4RKBmjkhe+UwaT5TchN17srw2KulirC9sYOUPjSd6FZ0j9p
vxv9j0BXifZQLbC241I6b5hv/MVzFSfj2+oq6aJEbqAfZPIQ9i+ds/2djFRhdCoj79B2E88dRvhQ
jy++PUCkYkQjCUPZEuCCP+kvZo7Qr1SRTVzqi3swiMwP3KTTjLH12/mmjBSouun8ONKHirMXfEoO
luMFQJB9bva+7v9nhhkKZ0stJnQlQeIR7ANAo5YV6KGp4MsnhKvmyXGDBUWEM8F4q3gQY4N9KXnL
Euyji3a5pfMuF6YFOf/IIg+wH006n0I3l/0HUnbeoAML3jIAV2LEscaTTGjG5VGJzEjnKHs4ZDjt
BpKagVuE8HlB8fNbfaoFq3qbY+ymAgX9H2aYstCr/r70Q3IlEqo/ZvIF9+mjhpJx7duKFtE7+lBI
8b3gRrwUISNgwyyoPJ+Xr1RHe7YWbUgfYxT7bKTsWK3McQf420on2f8G+ZsF5pFbi8p7psd5IvFt
cmAyXtZEU87D51aDp+IILNs86cg1VOLg4mFYQ05rtdFLRunEt5Grtr0JR3tjIaF2uWj1sR0SiJV9
OjqWq6kqAX8KZ2lI/ZHoMpGKTVDo0/qp70Gkf0mFsljia1fY795p08fhCiX6RjiwF4dkJeNMRlmO
izcRZKbZLJhtr0Rh+aOOXZCv3N1iKODC5rJWoVw1swoAIsa1kttZYlQlT2Wkb8tffjry338nyO6A
P9bX8xjKY5ppMIkcvad7hSYhWDF8yCjfc8kPODSTnNnc7v1nXiMDINLxkDjN3AeMCTrMoNp3st2d
DgBx1RQd95x64yv+KgCN8cm5WR/DjlHWAL+docgWUVE/RS10a9T81mU6+E0t37zAGosTJzShiw8Z
cvQl4byAYXkOM/J+JnnRiNelHcBgYHB/7PRTlzVmPrYZrMZ3yDL6KAmVmoliRPMTSsfErhNY9Ygl
yxF6V2RkvHvzXYeIk5tUqen7KaeryGsn2iLqXY1lLhAnBNKC5ZHQxi3cgmkAkssBDRAmB7tBrxDf
bLE+3Wsmd0Cr/UJ8G/gCSdd+EuSE8dO0eWkYmHdrA0z78xfzDFHQi4wVB5soFI2Y+RLk9mWuH3E+
NCM8VZ6CtZRCMI2nSK0eJ9SBAviDKMwKEiQBU7xH0PL1VSoaTtBAUBY6WeZypdWVd0EElfSLvG0c
cGvajMD4JuEbz+W7fNDu1/O8nvs2CgyQ7tkdQDTQFCnPcHlU1KRf6Q2xgmkPtmv9+OFSDpJ/SZoM
ILKIDGb1woL7oVLVK7S6Mz7sRK2Z7Untkvpxs/zR9kdziEnZ57bOEXMlI6Jtkr48wp8UVUYaR/cC
IkXPa3N8OhVHVGYEuKQe4aAMwjAs3NQHyFajjv3e1frrNxqven/o5dFMi0VP2dr9arUW2ejDcnDQ
B+mjvUSeJ2h1n4EfX6U1x5f6/YsiZsWDouaAt8UkwXHFLa4u+at3HEsUDZ0NUPWHgQhWNqg+SsgC
W7aFtZp0U1B2jScwJFVV2EaOUG1bpbPumBgyUJorVP0ujePywt5S3FjmhM2XPNk5PtEnq+5G0eOO
uuKkWZoWIPNS9D5efvf4ZzsYcJ3eIwiznyxesBXNslRLw9CXE9kCFBH2FPdEiMNCRiBBAknECBik
ZXHll3ePEVhs/yxx9uK0jxeJi1qSp21ms2sZftEl/ThWc8TCMqw7swaBPzrPXykLB1qDsr71hVPY
xDJIbG4KqVfgQNmjChbCyGqjHxHfIdFirMC65GHDBuL/wWKP7Znj4G3r1BLki5Ypvd/Mi2rqn+ou
Xsc2pc0OzyJJZR8Tqm2KFPnf5QBuwQ9KY247eB5dk/9xAgoVEuz4FWIDw8qL6ivkCtgMyIEscu06
Nw7nTv6SfW4wbektcejuX20QZRjC8aITNlc5tiirbq0ZI7Ze+HjrdrmxAKFNHyB494c2QxcR4Inl
39jKBEmW3k78csVpz7SmJYWzyVU2I13ePMDlvfFMP6YMHAvAIvTKA+mgvyoZGi9bee9T294T8Pye
QHm8u7Q9/tBKGppJgUfFGXkQkj+UwbaWhVTk3+jNAN1VQFAidwH6SuY1I1aF3XTCdS/lz3SZks0m
yJuFUxXQgxVmdkMetu2PSmob8l5GcR6Y9ZPSteYLgfxlKZL/81mx+SJM0AwOzlYtpby/2jvDqq3T
uVOOPyVzkbtXZLjJFbEZpW9VDDw3WAYNeGKYElmlOa/M0LPiF1yNoFDQToee1nTBgveCOoD/qqxj
c7Nu3kCUW0n7i705OhM998larYFr3yoJCVagemdvQ03cxHv7gHp1fgfqo9DhS5vtXvxDyD0oUeZd
DU5Uh1UWYy/u4MrzqbrUXHsjfR7OYnNlmo+8p0/pZT7Les1pAgUMZ6xj5UZOv38qqqeuHFAl2WzZ
h6NdFe0IWeRQsREsqkfxAkSlTwibRF/+jh1Hr3gQ1cPdxnnkEkdtvJcvzKv5bqEiH2FtqdKp+rZG
yAc3g2KHmhQGC1KzEXTbZB8mS1SB/GA7pGmaSNAc9uCR1m+N+hnU2weN+7p2+aYT6BmsjHmzIEMA
dbPuymR5CsQk2vAd1AHP4rujqWghv5hqknI7lpuu5PGBbt3Gam+OJBFlSxRz5PKZTH2Djz8umtdA
6jJmsjmGocaSRpO5LnaGER4V5LFKArYJuO1Yo6/RDdQEgf6RKWBZ/tdD584hJ9DiiYXxhYi1zWu0
hTBQBtxE+6U/qD8GcTkJ0K6kozo9rvfETSkk0BUJRP1QY2nZcyRaXAzq0heM5ymnGqiBeG6Uwf18
/Ae771E2QhP3czouC/H2DujgIUvXLDvOSTtISweaU1VLPf2Lj7ES7H1kHvhur5w6R9Q6pDOR/nDH
U5d+S65QZWn4k9lEzkFC/cys1vH+1+CN82UrqFYQRwd1AzVujZnkUATVBZmNDtXSmxvsFGWK7Ch9
N3wm6LWDPqKAKMKQ8fNzJwcqvVCxwVGyOgss4KMBiS3M51kcBy0xPuDKXJ8e6moEgjMUXk4biPxe
ECoYOo614eIYmr3zmz+stBLgXt6cLD9Tok0YZt5KrsRZph+9MpDRtU4pvclhCItogeyN+n2aMCv3
FEZO1558rGOHn19YJm2bKTuRK3sPBedkYZQX8fQ7PT5Y0L+MfY4v3d3nup3h+q9XxIS1ApWtOpHS
uvF/+nPpmH7Ft3bJSbzA7aPAHa9tIipGuajqCG/HGqyh8wp8TaYy/HeCc9XVxD4WZbJz73iJHWmx
Fok+VaIFJL2i/QQyNhiDN4lGGgtE9gZbDVanY/7bIhi31aTz81hK7nsQMxx+DOfJpY7AN7BAgXbZ
ejIWP3rHSAGj6iWFTAlxLBOV96W6YipPVSocW8xsVryS4nMEzlnk4kSep7SZsST40WLAwe3K8xu0
rj0gxFCvFNTCJzXAiPbNOVLAGC2CBbbDg1gtsHSHRXg2RsJsHvS5jTMjYNfckBGtpTlcZLRjcTSd
QzqO0APDZcukklDYD22rTz+LC54MEs2DfQVnKVxXLT7U/8rKISsLaO7NUo6t1zmgwXb1EAAxXagm
1QSE+dst4gsr+3aLvlnT7mg7fC2LcMLrAcJDmnNamtbOe6RjcdjMh/a7jsXSY64I6D+fHWD4TIph
hr333bZkA3Dlm+H60DhZuT4fSdq6HqKsnDItH6gITK/QFCZyDpwZSRIaRc2NChLmbstTHgV7tR/+
KwtCmEZquf9JyFdCJINXV2i96hINdeI2IEz4Jgnv36YhFyfZxDXgcwAGw04BRG1kovK2tc3VOhTD
PvWbIoIVpXj77tTheZyiOCPIMZzbZenel2qhTGI8Sm5aM0WHTXQVP2BpUSh7VoIK50bYXDKIwjqL
pm/8z26at+KqhqupJVSqMjVbxid8L7Sj3ORRI48ZAmEkliHU9gv0coeb41YHEreksLVHq5rapZck
PKGqJsz9D/kQZzFmO22YcbJeEa95RYGBVw+JOolF19v8QnU49qz0IkgWX0ObGF4srZpbrzRKhkPo
jIrlxxCOE/e0G4Eu42GEKjWQbGkPUhV8YTrOo/NgvBYZJkhn+mbMmh9Aoa1CEVs55UTWNyH0tSIS
3P0kjPWqq8stk8ifzgnWCODrVSboxm/TEXzCiMFPeYagBGz+jGeJheO6JS3iZQjAEflllwg2YZU4
8qClgc84kfsQ16/G6l17x6uhFCGJvR3HU3ZskD4zn248fQ8/U9MDgKw4zRhZwsVNUaVXPCnQ2JKv
lLbaolIfNzdCu7ZdW7Aivz2UnfXtG9s1nCEfp6MEBipW+UlbYqsGJ45Kca8dT8mEhYUcamZDV9tQ
llkM09F3I7kEMErJo6r4HCZfoY7sVtWnpWCLbvLfKooXrzR6ChVkd9hlx6EWlaX5aYYdA8cEGNrS
zyHzYwHJMlRV9BxMeNvCJOafUY5OXt4inEblmor3rGxWhYc5c6ox09EclaUI3X/OYzCJ/HV0a4u7
ZD5/9Q0iApNPzZru88BY+rYAKuTLSm86IKG5TF/nqwhWU1vCe9qLSX5WfHohMXC9NNCD3y2Bwe+i
avV9AtZfTJW4D48yjEyaRiSUzMjZdjkoR+vAFClo+q+0AZEMo7+6F99vIFwFhSWuBkgy0zaKS36j
nqAvLkSMX/XtD7m771NpHN8tiBEKEInTFn+rz31nrNgE5A8GDcDM8XXL9kpZiRMvTTHn6IO6uQ/8
dnZSlYnDySVIfHz0UEW8coPWoy8OZMGEhDWAGzWsnYe+Q/zyFZJWucNaV5BxNNJDh2v4tGSM7wYN
8/mne6qiJnqlYvLW5h4S9f/3AUdk+U6ggaX8CDiR9ABJ4zoqpgiGMWqachl3PsVWzeAOUc+epILN
HxAsa03oGFVKa8zPj/x/jHOGJNfwiXfKXjyFwYkR8jAnuOSpJd2c3NmeC8hSKE1d+X5zgGN4AxF3
gzJTsXvR9oxaqJYOxgsx3HcuAdyEREdX9JGrbhuSU/1J9IEoWydO6KZpQ3x8TDgualny6xG9ykmI
ou6FIV2t4icG1Uo977juacVLxwjYotXhxqaarFTQ6Cy9MbDmupe8K2kQnWLaDgS6nz5Z2JibYAYj
CA0GItiJQsaw3FAn4hZgFLNpK2VQpXbeUByRjhGNyntlCq2nfkZ0JOm1wm8tKhvcN1MPBgNPkvSi
TxZhWKTXRocR1jSTWgTPfyiopnNPrwiXD+r+RYvTlevNRYfnrpY/pD840GGV3Oc0bc17+CXECEwW
XoUkHG95uVYYAcLx63LT2lf38LBQk37ztB/Zs1LKZ9Y0ccPaeQsKi+lT2VWEsUo0LBx9l4mqZRHA
ruNDeZjHPY5FbO5GIT6MDO9w39vkYm8CF5HAtgLuLsMDah8uUF6vqCuexgQTO5i9tEW0O3kha6dS
sPKYbvEppCwCl9FNVVpwtjRziy9Nwpx+c9srVX42GfTW2gEIelvEHvVVnaHrYxKlUOZXOf/6Ie5g
byqLhG1N9vdzYIi76ayMA68PJztQQTyzgUS3vxU+2pw4UjD0k5I4Lx1jL235GW1cuwsLkaClcBe5
X1PpF8Wpct2hocdPA0AVa9ahzvoTALV6FN71N9/nJ7HVmDwMXiKbiDOwd47d46yuaUd1IgFWIsez
eQoGAHEztUu8AWKEF6XSgbP8Jy/+mjGFWJJ/WVzVI4SaZOqI4V6KWy5z5GBDI36KLlU9lY68JanS
72ZDxSgj3R6EhSrY4t7m0gHDz/kX6R01ukEAZzWEhxfbs4iRrT3zWO/CjKi0ANRRiwtIgxYLMg6L
iamPcFqzRjeZtBc+7l3UoMyARM12NVfxXZxIooifBVHaXixbiSTVgBWkuRDlGoxNlDRcoCn2D95m
qGi4hV3OxFJ19qZSrLZS0mdFqAjHpgueuS+DXgYGOHganvk4RJJDeEgkzoyOw5cy6bwmO3LRa54O
THn+radalJO4KGrol1xuCpmbbTXWI1R0z+RKaAuTW8Tyo48bFhaFFG0XqDOUUkXPEGc3yv77I6jL
3W2Yj38u0nqMzrz+FZfGQUDN43wMEaBb/ApVkV3yobThcdIIbgqMD6BqjlBVlOVG+CWRTa+BJ/Vs
79/FHfCA4lkkzKeENcQChpLwLx4pzqIhfrUaRytBmaeJfxczqS6KN3FZg8ObZ3q1mbe2dxzr0JCA
0wJO0sZb3Ehqi/Xwx8AgCAs3aLcNEFgqOGYvUBumqvnIi6D8AaUW57xPCOA5A/sBwnIToxQ5Atc/
81mbmTvULUfGi7bA+iv9qyU4U/Chx5XlX/foXTBbZwBVFICtoIBWJe5BmBaWnoF61YS9ClT6B5RP
MmbcvdexRVMhdSZ3JmNGUcC+XELqhHMfV20qqSHnt0xZ2g2nM+w9gpFD72L9vRZnmYG8IsxuE2ll
qcYYV+mYUovF2MG7eV+U+T28iwL2D9GY+naux2v3tj19Tv3AyZHycPNa4LE0lN6sia+rXHDwACU4
x2AZfrVXKBg5MBDRE8cyZsaSQ7YgF8aOCTQfkbmZLiwcpc5+c/2Dq6dcVWT9JR8NIa6w2Z6sLlMa
r29qaXxdGVx2t1T0MwvNplgK+pQlmsfO7eUBCA01SWHSyBmfgNbmUx8FECWwqQyLcPttcNgcpPze
ArowzVcb5AdP0im1pZOZF73I7LEhke73KkRjti8cSEmZf+8evCpbncmqP6ghEHnhKJq82Zo9lEdW
cQ7B2y5X3JWvipj7x2wcA/dLtjkWI/PEJjYN2kMazCoJLXti8Te99+pDk0CAWw4BkzZL872p5dDM
LZV2mIeGF0Hmfvl936i8v8pmFfxRLzOt270TmkZeLp+0fvfV64mkAt6Km6mnhhyWzESDGXyCGVhb
hOm3tdhEIXL1VuR9awsR89Za2NMuiKQBqUr4ShI8amjfTdHqPiMxSnwBqGvSexE/TwO8UnWIINXJ
owngODE5LuIovzU/pgzr0YPVnMeJwyl4D+7oeSQhBX6j5x9MDCX+8SqZJ8Ep2PtQvYnZNny2ildi
yiXRWc3yfixy1tXIgdvGsQ4K5S0pjPIMZmvHfQba5Ql/9Xt0FaL92RtVff8k+y1jU16b5PAVlqKd
5LUUXpu6Ag5YQHJvKQrgDqMmfxtYyT5MrKIe6yMD9m2aSrdu6kbLzZmXQDkZRFT1Ftg6AJGd1eLk
IVVexh6ecdZFZUmpmv1yLgBNondmVWZXeqkk1YlnOhx50NGyTeGKm4YRTVyutMW8hKz9Oz69EnwY
bnYchyxgfD1rW0UWwIcEjHPYXqmWUK+sH2T0FrBfTNmtLK/36cAPZYHurUQ7xaeDIfhzQ6iXX+H9
0soqSzNtBX5q6EqzsfM145Vaok3ie/kUAN1r5M7QQY9xUw6PxCfIjjs7LQyOOMeYln9Fney/pOkb
VvXrFqLvBgPLPOgK5wAe+dRC/3+SUiuOPScPU9cBKJ5paubrkVFQBsmoticNhyQEBhZ26jmo6GBF
t4mPZFHuMYoNdpQl48M9roznJJmuY5yYyKxRYaHbMnUbkjvQabm3rf9+jkjJcg+2beHangCJ4t4B
42pZJhGiyfOLwlGuNgHyILgyOJcH8Ka46ElkXiRFZKweCzYUpbKa3hitxRVzf8k9sgKQYFyN2VGg
GY7alC8d+XjS5uO46kkvQJ9+dubtNEinaBLoZk25LQUYRObqeB8EYZQoNLvQhY0CFpGLkVDTQzp9
RPtnGytbbT6GaqNWKZdnQnlqmkHq2Zcpk8KQLFMI1uRCbBewk5iNs4XF/fuKLuTq8Bqc0B06rw+d
+GUkwT/XD6vHGaoLR/psrOs6R69MO2zw1HvLMwJHDtWTKJNS7UGeFtZlkdswWRQW1ySlzq86id+e
2kxzjsXxH1yWs87vGlmY6p60ZA4mJqisb+YkrSscFrYWfSFkuGMJdZi9gwfOc2EytB7wvX8LOPhz
NPyo6TZzM6PMZ0wQ5PTMXVR3CB2QGEf/r1CHZtO3nR4cpFrPdBE7UxZqMi8af7Va1SDlMuy3niX1
vAkRWHWfqlJ/+zHnq2embDej0HiyEI+kLk0Yz3ejM5lMqlp+7IN+LoliofNvUSObjjlDPa/uj9+y
tvjpAYjIFW02+yHinfC3PEr1Nx4CrNpdMuQFFNWABGdbeZ9tVb+8gjTbtD/6BbP6d4nsN325LVa4
+kUsqYNIUKVcPEqDEhNKXF1yGvNEuaZhO8WY4LL882m1YGCFjUjFqtI5lsO/9CyR1vtACTIK/3qz
F9GQ0a/E7UDjuEsLeRVx6sruLZevvbNbiW3HeQslDzPhI0iu/IymNI9ksgkf3D8q/pdDbpF90z4f
I5nDQ+vbh2bkG1SiJ0fJ+rTRnwirlnSR0Pdbu8uwI3PhcqEJ158uuKyPgqWKPQvJS0eogUbHgTMK
Ns6SsQUAb5tEdiSQ9uUzY8gC4BrsIbWtU3kKUru2O2GXGRhRuTOXLCbOscW40nbrVznyV5ZF9mjd
7Rv2rgiB26hPIysV2whB/c4mEqQBez4pMj7VKFfLpcPkgUPWsLv1epO6RwmOexTrYUeAvz0d0bC/
+oywkRVGJq2ZzLrOihjFuVhqAHW86TW8V7+5pSxcSXEAJRQsXhpev4XohEtjmSYuvkxdHsfG7xpG
XaqiFyesk+X224nYwG3r/9Z2TElMt+Dm9AevjHxpDFALNYmlF+cjbklUjWIChmJUWYM6gVd/lYhM
uilqjkHl3wJnStBoQR5YrDYQGH/k8qXxdcrGSmn3KQBB8RfujoMf8o4efWnjHdk/Bo8927/w60ub
0mkR3xRu7j3nwugS37j/oIGnxx+iaTHj/MMRUc5T+z/okAkemelRyRSLDQKD1YZOxgN5VMAygnYk
UAQsBXrAPw0h17ESY25mOYYbDTChZZEcupdrMdyZG3bOP0hMdbYmYTQUG4jbK4NemaxUw5Lj+N7K
EX/UAZfn9n/r8ukT/tT93x2LmNlHP3ZemVRDY2NGfcY/rLpsG+WoV3ER8HH3Pz8iHvSzAohxy+yn
8OXzBumxMHhEaaTILvrOBUSmtRbBQN0Pvn0+F5VXKg+XyRvHGtbwo58SEFuN5Yu+etAr3kSxz+l2
f6kR0KkRs1K0+Rj3EmwlDBJ5FTnwUCfMSq1c20uWRYD0bgG6+2h2WA/tC8/xFZCe4/5PeGDUDVU6
meQ4EuHGqEB1N3JfTFZ3As7cNGLnLqYMw1yEHabwEp+N0J5Yodh837kApLBhg8tyoihw2UCdGYKV
/sOPbcBBJPFdV82ckC/vqCj8BsGMwVio5zg/YFaDudqYo6S0qo/CELVtynSvFS8j2M7GbQ+ngUtw
HXLXCog2+uuHNy+ADMeyW63a/VmHzYsiVf65+9O32Ot0nZJsJACEialfU3b/DTCR03lOj3Hur0/O
Dnnc5aDNrP0ygssO5gz9DYbAKNy0gDrAQD2Vg/C5VQ8Dqhp2D1CGQDyoL1QH/xa3JWf4yR2O+MJN
Tuxltsiuex0J3AMzBVbbiN8RQBjL3oFkombLGYJDmGVen+O3/A0scftsD+2txGpDPjJysI91cGfx
j0PbfyNrraT5sB8IjbDTWFcajVk0tdg2LLX4qZ6kidoftLHrUcwdA2ZOYphrQLJEQvpaWYz6Pr3h
mEIYlOtlq/QqoLziY6sEpkbOQWLPI78gaHKAJTfoTeemJA2rYHhMARbLmgfDimgSdBqlVzEId3AJ
2DnzU5/vIXhoAvwqt1W5MeSPgpVVXL+mZq9s/8UX3lhOjlxq+f6nxyiwk8U7rzVNS6OQmwj4lk5O
zWA7idsLpwF3oleyA7AJaVedkkVaMxrFgQuJOvD37xCHWciOcqFJh56TZjzOJ1i+HbJ45S53DNWt
HRVjLCvGun42tV2EJ/wUAr/bsnVeQ0jeQaGzUHG5VB9hjAFu0/sCWTh5lBDWjpYYq2et7ZVm4mHm
focYq9EMpgMplkuAHOBd67vMRebics9hK+HuBRgw0ctvu0biDt7TIe5z4JWnkejBGC0wAStWXJQ3
MZcMKZ+fi8ZNp5/JD28djE6k+N2rgjTFOMM3sqKvonlYk+wyYRcT+Or2Nurfec3Q0kHfyvY4LIdq
4cZphAzINqYjRpdA5ORfDl0l2g+GKMQRDVWMH9S7mwvH7yunrcSdYmB+MhlHEGT0hJjfeDif8QJJ
ttxhI334jC7WAL0fOvWvpm7R04/sUWfCAJqBuNZxpQLw0w9ZAXuk673MdRwBiP3899PvnWME8Yi7
j8eAaxp2LvDyBsEdjhnhidZO+Mnj2Xng7tWANqmgD7ZCjAH1isvKU5j7O2ji0jiu4FowN6bAsGZw
RDbZCKSlyC/YPg7S54it2UQoKJBE0rHPR9L42Ix99mIRxZ45+o0x3verFX1ml0nsFkQe+97hMWb4
Huo+7AGlClFHve8vsI/oaHt9nq6fEXjgqmCKRc+eWL5wEV5zM7kK4ZkiwC6AZYncrXXKT5y0Tm3Q
CFEVa+rMulOsj2oIfzwaxJ11XX6/2+Q5RcC6f4MTdYqYcCXkN1Nh6hglJNPPy2VFbbMPbVcjaa0/
RplsCN0qXmmB7cdh67Dhk4mYCdGXoziaKen1ZmCYWPf7Vy++q6JFIjZCZaODW+ohVIcPASkLbwoN
vQ5CxXrpnD5azim6KrZqc8G+oiIxGidH7r16//vmYpydZIoX1ls+auBp1oYuX5KPRKE84ri6oycS
OujAtaNPc0/RyZ5N2jGi7xMZWVMsFM2YKNMAC/LB5JpkLCz7Q+zKStm5f6yXhT+PGY2Jcm4ku++9
yEPG7jdQiP9fKKZco4q5vVDVv4UajIWe79y2sIjpcFMray7HHWy20mxr+6meTFnsuEWVYro138xx
tKVxy4hf1LHQ7DbLRRcFp17zS3279EPWQpz/lNvdj6xqhRj4tvyk6Z+SpGHsIQRNv2PyR4jI19iC
TkgTV9uihv7jxJqAxZM+fLtmMlZUnEHVO9pwW5Fsrjnl06nnItKBLp2tO605EBEBV9KwbPiObWt5
3x+ntFgyJBuKQ39CRNXBKZd/iPiuAO2Lh5Dk+qGfjIxcURsCCEMTq8utntFbKvwLjntmFYrQlfS4
TTGchK8Tdy5zQvlr1gckrO9v/v49SWZz+S3OPhrfrIzbnWPoeGc1OA+z/6/vq+hJopiiEzWns1b1
VN+C5o8u9CQs+VCI8T0v7HMNNRhznhJ6j+/Wz1Yy7/P8qCyEKn9dFfinlr03leidzgaxJT++6i6l
bI5Jb/AtsoD3cFcQ2Q4ywwa/VEDfNX5MXjcaIWRDwkAeMyv6WMGqHM32aeBwW3VKnT7n++GNzMKN
6pOIfBuwDUx/6Ih1GBkFQ9N0iJjCGgXdDhL1Kbvg91SPpKECA5WSKBMOsemu9FFziZgLl15gpYBi
ARUnzOU0uwWdYTe3dYNn7dBApEvDUxmzjktHwUoVy8Y4Tr63F+Ke83GTc1l1/24oDkKoJVScqgEA
IvJxZ30t2KzAa3IP2wGphRxMSblJZnyDVlO0Al+YeZj/9qA3APelfdXyjbZT9bkcWwc/RP9xxNom
93mJcYAVUb8xXgsCqmduM0GV+WaPQf41OCBVHzFAa7m4OeKgFF2DIVH8OTyeFsnjWMLghnBKVI1c
rI3U/Zdfrzut9/kW2cvzVipi6DCQBxTKTfJpubHXYcE+Hmj/nMym42LWT8safSJUcWKI2Z8mbHe9
YX7tIB5ox/J68NCk0GSFGv1vALlXKYAn90C3Kms8aPgk4+2PQP7987HgwYyYAzz7TU9/orbEAkSv
TSetOGbqiFzC9eBXVdzUQGzq02wLmbyZF0BNMVopBVE83FhaJNp/835kLSe5tnC42+PapjgpTHV0
CuD5V5XUekWCHV5DCR0RlU9AMlyLPUG6r1VHPkdhIPvNTYEGfhBzxBqJNePrc5Kn8DuDDHxSuuV5
UHo39g3TVVhyUddXA1lvX21oUIOoNOBkYn8PvYgSjioFXvJEztpza/nJP9Viqv5+BLI+QBxMys0r
8npb8eURN8FV2NZfrSCoR6cig3OCc5DIt13BaX7y6MhWJl3YTBidcmc5YJ09/qTISjmCQMwsDIc8
UUdNzpDru0rsWECE4TZ/SWFR35eMhx/rEh/9BKXkrj5dRXDN7DlKSLM0Yd8J80Np96+7evfX6bdA
Ma52zUUdZllp8TkDGkQVVljDd53/3HY/ZKcwjC81EnjRMrxgxC+gVcdN19oXL1vBFj1aIK3QV637
O0j2woe9RaqBCwq0dVHs8biUw5weBJjbbTCgKmecqxxO4kajiHKqbZUfvZ7WqPlqpqs2zVDMaeG4
bgWaK1DaFP3qTBJbVjRDtknM/3ouAVEfIn/gi4a1qZ7pRpTLT6AvDEYXiBrzArJpuxxoimXOBQkw
009ksguVaE76xFSxDzmeb9tIpw3AEL8kcKLbViZ3tmjKJeMoa9uUT7CJrpB+g4JEzdtNwLrOC+7h
P89B9xR6TQMFdlFLgmIqT8a6z9Zv34xczi3BNPn+7tdr/s7xJYHg+m8BVOBPphasAPB64spthzXs
jaIwKOLsUAa2O8bteUKt4WFWdLL7tEkvwLBk/rOGWkqZlPqrIIveQeykVtyJYOd72MACdesf6T4X
+yY5OeRug9n4PQViZtXiV5AmO175PVot2QSMVJv37slulN9HciJeibfrNnG4c7ReeXVXU6PzoerL
CtoQJdooG5Fz0GKwQUqduc2PqHpdggBtn0fe0sk7z4GvHV83By7zngjeANZLOmwPP4bPQaOW+KzM
f0Q96MWpTpD8nhObP9BfdJKA6UB5Wo2Rxlx0NIV/ZLKfvwq3vefvEoxelUnqbCTfuK4aCJHWHEEX
ugSQHxuQQ7nogFtHrc/Pvq4ofFD57U9QOjsqbSiaUF7S2IqbB4y/ifIrPHFllgWpV5qKIzhca4k+
8kOXnBu/8FWqmrYqJ40SPaz1u4s3aEPxovCyjSLhF9MGxOOGM3ZuJ/Qxkz5QAsJ9jf5MQUAwlUVD
WWUA/sxyMVYU1jMZkTIWJcOJ1Jh+uvA+jZRWKNhIdZYsqWxIGgCIqbG8Ww4JYZ6a0+zgEOOpWDwj
wx+TUr8on9uwrrb68XWaWzamkA4LG6jCWKpjzFKN1dVIpaG1+ebOQItp9Z9kW2tfpOo9wu6w44+A
stM8CoyCiskuESxV38zDDtxc3kx4bAGHSmgU2VTXOu5Q+O+bS36icJfvOd9BJ8E8OkCEBFEd1BgB
nAuYUWBBckmr4g/EcM3txpp4+wnD26hEMoSTO5J0g0KzU0vEmPVdlamudaYCSVVv+74QfQqnDjtk
QM4hnYsrl/F7XPHceb2hcvcIiqoqIvf0/7bQRIc8ntRzHkUmNMhC51rqnO9a7bNKQd+7IaMiwsap
shP0gmZGKo5u5wQMDPW0qNmaZe0WRzWOn+BMJM+dswG9YSUg9hLw4ha5wuWPGwQXsJqoy35InEp9
E1JUORy+Mw5C3Dcr5hWpNryUCwrihTCKteUWT/3gAh1ua4agDYlqU1Y2zOLUXd727KVZxYTvNQcx
oQBeAuu7rI6OhvR9jkZCaPKhKF2qXWzP1tEaNvWPelgW3hHgdMhOdSJ8Vc8fZ6FoPOgZrPCedztR
7LMcBgMgs9YdmM5MNMBnyL6rKxy2jegpA759aqQ8BgTAoIMNEkICce8AWLMQHFdGF5vmt48yLEsP
PsNcd5H/Yii6PElnOycm3ZxaXR5UU5JyBmYUgMxMof0Im9Qfd3SNOcnXeANfgxjsErF7LbtASzHI
rrV4Evfc/9pcNjuzVvfe9NxnHqHsUpdmjs3uixMBclxgdZReRpqnDln91eIWMStDOkl37oryCqbK
Nk3DTV7MVV7zGgwt1Vb2iYpWypB727pseATpoYqmSydfgwUo/C1hcrgD3p1niaZjvJrxIqXpRi1q
lgJXAc1N4FCcKNyX0PASs0wlSqg4cVcyU9bkXR9+K0UvL/JilyNuzSww6NiVohTFM1oSeysmicQF
QgCy7f/QKmatUsZwYzCtftqmM83fuE2tExzbc+YzgIboK1JrCLkTtCb5yDM7bZFuFnrQG7VcsgpW
oM3Uqkaz+f7hF4EzOg45Kp5EETPGSLNQ57XoVY/G60v+JNiCfFP3Go+VEOtNk43kuo/KY2eHp7w/
yIj7B/imOv8buceyZJMSlnwJKkFUP1KFYaAev+kBdG4I+Bit5aDzIVgJQzEQi0XQ4k52gsQPmrzv
TR5o5ulHhAwJYLCovjIwBSRRV7Ye8XougEasyWNktQu+qosKt9Fy2Q7RjskXBlkReCodVDNAqxjp
LpsezpNzRdwv7R8l5FUE7o1OdcYG0FlnULypgbz9xBXp7WdpoNtSVxLAAiup+IBWdt5GoFr0wJl/
VZwP5B43f+KLMeeIsz9X6An3vo4W+bO4Tasxt+o9KInXNxqsHK7Xj9mPxrFnk4oqtNIqSSON9mac
t4QOyRdRhyH+PeOAr5eE5x7b10l2sOY57/FoFRC8tB4u5yqF88w3ZayKqg0QFd84jyQvf6lAW/oH
T94R8MWKCoN3osagmf9137I5zL5xdHIV/Hpe81Du9J9Ue3unXLv8Cu+lTJZ7TCXTHZXd1PRbvmv7
ybFJKYW+Zp5eb+9X+ROkULKsAtZfRmg5zKKBSbK9FNVFP7uernYnMJlbe5/V3n7VWQ8jWkZdgfcx
u24A654mF7cmye8mfO0PZi33UqLcVLGXgJGAYH8osv0VbqaEAWIQbVSbd1bIHqxAGdG0jcOwMqzQ
keAJMB3IjozCyExLa1pA2ossRuARQlrnVYLTYzhboX9GL29AVjvB6Fs33dISHV/eAbE2yBrQW3X3
cHzHZHrZjIbt3hlXOpk+TiuINXE6XKMGhJw+IV/gSErEfQqjQ9hbtUCeNbyDQ+fMJ3+A+wnHtwbd
VqsELTJLnx6zEn4MspwLnOuOV3yCgq75pZkZSlFqOf6xGIHbWZ7+gdCiWRtYcZXAg+Ppsztvuj0/
dOyDJL3uF7EHubPa/c+r+nzz/jfLYGjFX8iTXbD9Dh6yVH1z2tvGjwYM+8D3nzzZOyMJGfPapEdh
CCbphppIIlReUIjwsWJfh+CEII23/0xHtLD8ubbR5MGbb2S+3RJmWmyaExlCC4L41tlwq/rCMD3c
G+1oOyYhkiHPd/tN05/EHRUtAScmG1RYivQppT2lHcRTMww+HkjUbXVr3Zdovf9cJ8UIwGy6LS70
e6CQgBbu+nPFncKNmSf7cDU3XbRE2SGIrxBUFkBwQ3bphDgzPQgpJXnzl3BD0B5IZh+UiwAL+6SQ
0HoeBLGNqpN88bF+mhs7DNz3vGOKDOPvyNM1D8sko6JAwBaY8Qvb2VOFKB7qTalFVCOmaLiJsBTW
mgvs3VGSkLND2Ptp47fw22vvqrIithFu/riYXLl0oeSmAFU8BC991dHrqwZ3rF3moPZAw3CZJgOZ
nUgmMGfPK+mB1P1Jv5ctY2ebxApKVoflinMZYiNljPp7kcsjo5UCBYQxKSH7LPmPRffowK/JJeVR
9xbqPBDt7QP0CW03i1r3cu1qdygpAcroxQJBgu1TI5rN2KkMAY/Mi2NO3foyj46pGiZttEqcdg3e
44+9jJr3B+hcriJ4IyFhfm2d5A2+zZR1Yha0WnlRIHNSFK5Ppv1AKIC29dcZynpObTFo4gSDiwA9
tzNJNEKL0UdwOwgSXApsKyvg5uFHzeR2RnFvmbXt7cnCLgd1JBqF9IPncBG79IWEvo0DiesYsnIC
ENQEdsSWnsbhNfZflRiE9AjOXTObZaA0ETCj58yaANK6Ea6/hvQr1GJybrI/3QR/GmleTImSuWd+
p5oGe52smUgyHYHS//Fj4pNj76LqvafqAkfoGOHmr2atlNdfIl9VpktWRlgVpxQXG0Oz3xRrVhBP
DLCNZHLXS7SawPEkmwjzduAobn/DEeU+LpgloooZB6CF8HUxiAcSJJHQGo05nxa9DCzqOm6ZpjVl
iuEYo14L7cj55/9GhTNg37Ql8kCY0GF3cW1Och0lgKk4GfQApLikgnueOWoXXU3gOVnUWBipiOva
yKc4j/Y2Fdqp3WyRRf14+ISgwuIZCyTRhg0ximGffnTA3QxHv6wCDpubYpQtZ84v886t7wJzgfNH
JdDojefHVoq+gDNsKfrZmhK2thT46uYCY3D/NKAr2VvwRT55vkxEkW7YDmVHrhoEp+uCfdzhXd9s
6JqkurYzk3YgEBysIMne+O2T28oM3Dqe6SosmHTuWzW+8auL22xkXQmawTVb1gy9Ahowu07W1Dqi
VE8oHzMqXXvceBFRy8BsUCdoEEiOeSoIaICwqNopQGkpRESbpyjSotAeKU/JO5H5GS+44oS1A5S3
NytLJm6qCD/nGvv8UgYX1zCg+0NRd+aKPtnPML2ryhXYnwctD0LUBP0xzuwe9PfT7FsMDz04ajKf
WqyPTJXHSbnbvAeHob3IRHBzdcswWh/S/3T4kr2NO2qTnfZBkAs/ot2BNLU8jzeAA6K4xp1pVKRv
YMdLiR81cTjmUPyDbrKs40Uqblj8lh7uo0Z9A6l3xfFxutqWrip6YWZLpSCMsRQPXrVwaEWPP0oY
tswZ1Tynr8UwWAZ/RCsR1ViRFPxZ4i+VdODV531+9yArouPmRiz8fwKorKwtgTTqOfuPeCia2S4B
eh9V+ITZ8PgzwDw+9PdYb8H8E1mVfCXtMY+qWOUIrJQpNHDjIaSwdaq6ps9YxFcLV0Us4jYKPwNz
UTcXrwJ4E34sPb3PhYV6nYZ0dNesCQqCfVmQKkND1JDXzSlY/GSF6fWCiUa8Cl2++QI02VxVsrn5
aNHYCzkNieg5qykithbxOFU5tdSr5i4ynCCEkLynDFz0jEnlsXUEdGKZLjBy3HuVst3hP4xVOHRC
o2rHn5nylFexOYqmX5I/XMNeNllH7LGCp23xCrW69Px5bnT6LPBLFeydTsKLvrDwzgoBdva0XKs6
dpIDtgw/Diokt4WbI9gnu30kXnvw22p+m1WcsljZ/GZhl2xSCtptgGrlrnO8DVmHLl6L9ECJcX4v
DJQgGV0oWPjOcjYLK1O+gX1jOrQ0WHD59Sc+t6DqpynveKjha7B7zCAuUC+b9BSbIsWncamfCvv7
0lF4I1Khkw10DsPcLOwal9mrIqnFXaXQjryxI3IeAYnN4nJonbz1SUZnc5e+F2TDEMi6ycpuiCSd
RgUooNMtOxrSDAdITv0P25HYN+OnYEjJb9Sp/9zNrShdTk8bPun7XSty3VpfYpqx+hmMZyMm0DnU
c3GWx0CTeyVNHf5Wm2/U+ufzPpOVgLtwEb5TTAZirQVq2G52MeMzeTQD445nXDAnDYkHPNx7Fv5m
1pK94aKxEs7NbwUbJN/IXc2dEm/hnjjn5YeqGCvTQeluVxQZY00fUnYDWJpp54EP/8fwtYq+hnQW
yXIJJJU/6IH8PgOSLi+nXVu5qetlbpNRUMeUof/berVz3zO2JR/CSMIHorAI4aGckKm3Bzd5HhSV
EV9b/9jYNW4S5A3O8FgnmoAO/9VznfYHFLO0GEzMCqnJ+FFqPgWCAZhjkCQcsIS8N5or4THcU5CW
I7/LLJcud9HaU29RCJSkBc56XowD+vz6MVKLgyGnwHDwtQBCUhQj2nfIEdz2sYWSFEC85K7SQZ/G
WbIS3WEIyBm0f2w2Mbecq9Z/oXWbBxTGgDegKdHTFl48/gU2hmkHMH/zErrZO/7GJpnEW3u2gEPl
OpNYqEPOO+hYpznlCqYODir5bgzxbR+iPxkt2J/cJY41+y/9/2mSOK0oQHy+B0qOLAHbf8YGa1RS
GzaU/uoseT9sUW00MMf7A0yi3mcg7Kq63Hyioz4RyIPlybeldVUwygDe5aq7SMiAE5DJjE5id17+
GgnhsDL8KttgWrxIETVeNXZb5Q+dKnjySseaqYaZ9XKTR6zjtXSX+QpgzAqvUYdCDpuCG7mpvRIX
KniRglMtc72HT8MaUxT2VsSoV6eY7AjsaCciaTtB9hD3i2YVbQJYF/5zBOhqxEjOppAvSGewwHL+
BiyLImDyCkIJIDjXyXOiaCn3CNA4kYXxv+cqVdiyHbkt7A6p+KbAybzRX/qTG8BtZvieMOBrfw6S
na9xMgM8VOy2x8Ybr+H+06vDCIq7VZqKXxUMbe1YmBqpVHToe3cTOaP4jjBTcfwhXag8c58RlI27
C1CgGwYtFECp6jyJxjtyUyoYlXLjxlQO8J/rx8MEoDe6Xjyx31LExMIcLFjgJOOzuGiTX97aYQv1
5RGuSz13E8P8j64Mkb3jvoFjCEBdN0ksJRQZX7YRxcTDAc0CgLLk40u2TnQuAYwpXnyZiWJX3qtD
lbS7KdSJsu+L6UWeZjtNnXkCUe9MnzRc1CGAhLgY886mr0dxKcYH0DpirsD6ex0f+pfHCJBvkTCS
DT+X4vxmmClto6TJNknRdKLFZ7/hqToHgLiQZXD3XYez24BuRBCRdqE4Ab72UotDjKQ0tRvjfM+b
cLRdFKWFGwuA+RLSmMhEG2xVJTFoEW+vxOR6I9S4cTpxxbi66paZT2L8p/aAOR+IJtk9W70ACAh0
Vf67if5rPFxop+rYhybtOdoIEJ73TV1iwnCuk8SQWkVPlr9zsjeqfiYe6ari1MQVu+fcVflAoniI
FjkRgzV1Rq4GpZA42xt492+6fJoSzYX3P4fyFaVwfysjfTYC6YBw2zqAh+Wl3eZee9++m5WOCy73
Ij/U5lDCKQp227sI0QLrLTOnv+dcW2F5zp9bUF2PHMNl+6OdstJ57hz/s5V3iDPSd+ivSkQIaYRi
8/S3+b6cGE+ns5tKXsfu5xg01GDIHzlCnqmM/GQyIhT7tVyeaoA67Ox108k2SjFGsnqFo53F+YSp
kObu/qOUCuONA5KK0I7ICJlOPktFRRFAp+maSmRiXgOpVBtLtohfMliAAEGkyDLZQ1DIOJJBpwAJ
0Gdlw5uYsCEPFhYwlBAZOpfxAAv+4n3mIh7bBHiwSQRV+mtdTKif+L+PqhRVXoHGUwKyl9OhU+O7
1ZuxAlNNe4o30/ymmy5ZvLqLmNdcjPPSTO/AO37KIZShe4teVzsSU6KkrHDMNoQ51tPkU1YlZxtp
jXxvsHPfZ45o3vmdnNwlGpWHIombY60pjdw7CP22y8aWEuURxKRIJ3HUAOYr1rsT8rQU5mgkH7uv
x9+LnecnlmasrF/In25Lm+nnD++I7n/tOSygSojDrhH6j4/d8gvHhkrOEkwLQMqmgBCNQLn6Wn+F
3OGbtGl+uhG++WPkZuf6Q4QMN2JBN8ZPrfhqnrjZFQl18/Alr32yjkDpZFDlHiyNhO5aB+Mxxq4g
La9bKggmG0ENpzqX8yzA4DdmrJVILNRrNWeoSvO3HZ7fW2DyFCUHBu3dkozFUu8E34s5NEvr34r2
tuGbUEqp/82wOHT8giwY+Gy4fiv5IR/zax6A0ik9krLhMVB1/gA+T6yBnjmw6pY6lw2AT3SUEcGO
q6QnAJ1jERCzrOzyj6Zu0roFT3PWAqb3AIj4VrgQ3eMBHCVGzosZQKnkfYbJT8bOut6HNA8hy7G6
Hzbs8VV/mQpieLWZyfG3mOs/MSuSEA6FG5rltVwR27DW3a77Gvgf5j9Pjlrp6uziJZf6J9Y7Xqkl
R/mC/ay2p3FK1/rkXnEOpIcPBOTf71h61KKMTWV4D9WaSE4z3NPH5SUIHIvAAyZ5JiVbDo1bvLjX
rPH/yW6Zr+wUX6AIrTL1rnIS8g2OvsljW9zmhISnBf89Kh/8RaDakr523BCrVnSx7KX2duVpQnwM
ME7dhYUngalNp4q+KOL/Jy63Ju2gF6rLyanyPirV9i6KHBkqskzsdzNW6YBqtRQrOJXaWUuEr8D9
qVZQq4hJv29gG09+UFOZeoRdDlJQlQ6lAbE9GceMnaVuZJbloZ5QkpwzFoRiBwWx/k+lOdab689c
qnr/jMmT82VnFGxeS8ARgs3ieAEstdRLfBDV1BT9chmok0CgOPeKC5euw8od1i6D6sn4D6pMNgb2
oGylOxuEmQucd+nUblpggiBt0UJDMlzGUcVlL0FPPPsLu1ryAclUAhyarGiixTuXzqmtOg7J7Ozw
doAIso+TaON2t2j5rOw9IjIERe+3/edNC2mSXxiI021s+9K5z1Bvqd1Md5h4krPfT625acxiwrAf
aOAZjhfgXpgCUwYs0Vhblhi5TVOjQxpT7pQiGwfrrJ7KZ8e97urMzOossV6TG5hRLf8EpHXpslVP
fuBgXzToRfV/D4YPuwWdMKm0bUWuDsmAN+CVmtLgUQ6rO/pzh/P3gQNBNf9EtLmuJkHVRKDKxNBV
oEvMXZ0PG7/dHTnHd8j1jHDykhCa+TZ6IU4fgo/dOiIe4mEFySHedWmatmSabWqIptfbGfTxUwHm
B4WSxbYDcd11cQmqLAHpJ2eODkmCbqXmBuw5ws0DpXx//lKJbxnWwKxsVNw2FMGbr3P++vrG4dfU
rDMTnD80uh/XvuVONh+51GnZ9hLAY4/PZtSwPB1vdRYqqItBOWlM0KEfBClY2DIk4/YwYusqY8Ur
CV5vYG0RluOGR5c0kmr0GEcVX7xDV/mfI4tsssaePm8vd0EbKlRMUOB4A2eqVLCsVaDCHCL/lmTt
fG8HNlkrhWSGV8cKXeGgw4xTCio30idL9mG5dcbGaL+GjDH0C4arVlKzqvpYVIpOoNYCXjn4UXsg
Sow5gH9PZEz/JG1Wgvsi5S7dY+sfLV4Dhji+x8zs0Jj0uu6+/8bOwIAz079j1RLA9IyxDf6rcU44
P+XhXY71Lzz50+o0oKeXX+LoD+u6gVo3wnKHRfEW8o2QS05T6PQbjHphG6nt1zwVgN0qbsIuQPM6
+UMD3E6XD8WLk2wlJMceoJ7K3iQoGnLyiZCKAEECjkBOZN4SdidCSd4kPcshN4GrauchtFc8gUB5
r8yvwAS3Sc9+8gmuSgg2iAEF1eXiOcp9Duja7rnTBYFGhswq+6uJAsdYO27OG+yVysA9aio7BkdS
ZGgyRHLhiOEp7XGgwaBqc6CjD6gwpyDOJPTdPs6oFX/CODTm/VTeCh6M6e2Lly8PkdelXVUSR4DW
pfVVSCbX+7CTZ1mdAaQdU4cEKMwyiNHTFKMrsb1OnOeyeKH8yGPnmX861dcE2Fu1wVi3HsQOV0la
dRWJb3tj1gYhTQVpVl+wOZrBbRYdRGFupxk7elOee2L//DtXilx9C5uN5269FU5C+VwNFC6u/ojv
xEcsIBlszxbF1ZtIf+yfH0VXptRo7klOEm49Zm1ZlgviBDS/nBa+2Sn2YF40OyWGm+XOWLn15WTd
IpLNjzM1cBSz+9igCtnhpF9Jo8AM2tixKMKvtc+nDtQvp4L2S34xTlSeLfiy4/DxHWpoFIn5Frvs
5+E9FYcTGRQMAzOq8xnGJMMBKFBh1unu2q3AV0KtvCBem3BYj1fIXzpxxpOD8iJZqqR2lXTyLrKh
dO84OxOYEQLYlAqOYK8bcAUqEYo9jONDN7mpHoGnybkre7uh3A3kTujV22nCiE6Hju7aei5LC0jJ
gEW4I7ricEZwsvz/Z2S7MKrEq9vSV7gdn1vc7Ht+oI4THD/LhSn2icoyYRXpHcUyQ1FZToRwIR//
ckoi1PHS543/cDSAkDd5dvmyplWCLHqD29nkBhO8k28FNRtPt/w59maal8Cecz1uKWRUU+DRKGyM
RyuyrctRr6Mj/3217pQHjVnivvx6amzbvVmrRWkzhk3lbVSmEfr31m4XvtBjb79x20Tw9ZY9MjF6
JKtcLbhRoNAck/NH6VTJrkm7Lni6xfyDcx++G0KJxP9twT/NaQz3vYMHNM0zE+6ERJDrvLune9bv
7XohwYRNVyXUflcdp0jsNSoDTUSMGFHkfZtnR254BzONvMXU8ZJKZ7HcgDFvRRxuFYKo3Gxpf9Mu
yBEWjH4OPQUqhwnKg797h9W0anlU5VZwyhcArWp47qabrcFFe1idoULcG0Zadq81FIBNfyCfin4C
cnI6X9nXIZ1i4hYJIRUaV1OOrbbm9Z+nL29r5onBU62vIFhO6vaDYltxQBOjR/JR2yviraFjdLZG
9gRykXwhW/+H2MvAV9OsRLRCq4X3b2yOL2BPdTR+hG6PUJtFCjTWX2CjhBTxkL2Gkp9SUZQXGly5
pfvEIaLZ31xL/yqyajxHVwpPRvnJtMebRpc+V3/WodtbzYGplMPZOuZQV5nAaCcKYfQoFK2lZRBS
R3Hh0FMVhX22k4uaz0zAnlK0A3zqe1NGivg9UpShZP3D4zB2h1wt+y7zvD2TObizzdVRaMUtDur2
JkuhXPlerxaRPmvWWt2YoyX9IheLP8wP6I/5FYWKu9DmR0JFvCTiDXvVvu5SCMs5An9k4852AxbZ
x42k66OwKBz6p57m12b0rLB5ZZSjpBBDIJ7pmnDjzwLhH6cZgpXxAK1QqX86SF44hZVGwo1aQC4s
pBAm3gR3nIRbHdHA3H54lzJ6L/5u9Oc6ytYxYCdZYxr3HF/xPHh6DCFlydiI59NNpb0eBkjqctvm
Qg1vA2AlD3a+Q2LJ3R/4M+jmdLkQhpSap3A0L2F+PbZv31C0jH85XGqPSgJcMr3Ei9ZQd9zymG7b
uuEwbm1VpSV23OsGVr/JBQc477iEJZywuqTnY4WADCkRb2QM73/5BDX4GtxrebCk1znnCzzWrOr7
Iyv7j5kfeggXNwaSbRKOuNn2xwt7WmipM5gBzYhhKP0lA+xM1++UEFI3guzEviYtw6X6rBtHBlEP
EbO5LPONwSU1mVAkOXR2hAjfGX10noK526WmwfgqzGmMLMiih9E748/8LTXuciV61146mgC7hktU
GCdV3MRdeQZ00YfaRJ1/Jnt4xQrWbVYVnrZ3l7DIWzcNZcsl0lNYvCZZ/7N8Q/0lhQ7DHqhn43yu
EBnW7XCVPrD5GOa4LAN1M2GrfGS0zn6MhDqEghmO7uVFErIdC088kiHO7I5dcDz2pdFgieccCyjK
z8GZ9BDa1h/3hZT9WvVRl/Z6stmJEnqPJzPzcRwsC6saEswaGGVC/RyS0HShjpWAFtNsbhO3ciis
Z8H1iMWpM5BjXxeVzLw+Lkw3NlIf7P+L2rnjifhfsKPK1meTE2zNS9Zj9eZTY8XsuLXhFybmh8yu
/ikyfL1MKDZP+GMDB/cDWNOzT+zfqBq2RnQeSotGUjZg7HdAebTCLKft2ItEOpXoACEOYw8XvWff
DCoeeNocMqa7e9gPU5+4gfco8QeMDBe1ZILj1gWvnBWuMBYAgu/gjM4/atCMTIBHRtQFtOY16+N4
op9O+vAcfTpG3y/LIm/I5nFHGP7KjPWrwQLh6AAk4EM4a7PueFJ8sdum8Iob9QRLmflZ/OB5fbkJ
rv3CSlHU2+RBEM/XcxetWj53thiEVN+hHmpc2iUxJQCwYSOpoSsxdqgrdOzNMyIEoHg0QoHV/zwa
dcVwlTTpXoO0/ZkYoKsQn5LyZiZUPwQNAHjvmBrPyN0dkRyzhh7Z2OJ2PpgVYuGO2mFoNlvb1KyP
UNgO152c4HT3rHgUtRnJIlNDfP+BaMiasW3l9y9/r6VyZC/lAyoM5UYVI2k4YJnsE2uGBqxA5qJd
+B08Vs/84fRcpzA5N73AmVrKK0Cu0WWdQYa7LaRYjXtxrlM/wu4ItdbRXRJJA3twHDrRSDPXub44
I3GaMldKOyFTmjj9GoqqASCDFS7Jz6c9IPtFdh38VOn9azyWZZMFJzgLWaFoBke8kAPaTV1zzXee
LBex/ahSzLWUFWO7YcjGc2AedqIu1wR6JZrWyH+Eg6xL2231Vc3kCHEdBNMbykouwgB0t4x0LqtB
K6tcsL/CYCoQYEOFdw1l8QttfW2XeFWCd1eWUil7L7VmAQgYIgm3/vCvYSSIoeF4qzaEwG7ki0MN
ZprbURy4vESp8fs16YV8yZIlmoHzF3mZVqbGfy/Ai63ov9ztsvhOxy1ZAvdRF5WGb1G4WfCTOtOE
d9B4dNG/t3BOD8L39N65aYDItxdrOJgHhOcGlPh88jnm1qk+oCk3XyLnIvo0yjUqtVmEp/gh4nQP
q7lC/GA5xvFSddg6ENK7e1CxQ6ySFFmVTiAW/EFBWTjoZCCvVnDDE4kTs9W9Cn8FrfoYWGpjTYjC
CXgLSalAXtzhdiqMbzJU3aFG2z7uMmiBKJda1+m5Hsvq9UROKpQ9ZNmJPUx+qIY2B4hxZlnzjbSl
JDv+eE3hFegXZkHir5BiWMduN+ckjhL3OPWn0qqEazbNfWBHzQtoYLn+pW0C/j6Ny/Ji9bwZmFqN
Dzv7Y1QihWItocDNVB4uOdsq5Vb6m7PbLaU0aRCz/3O1zv4q11i1KjFM79JutQURypgT9NY206KC
yThXXE1XH92Wpn3gCw7qhxW4yleiHAYmAhMal9oLSVU76r5Bl0bzAvPhhuHXxW3vH6/2xIJ7x+CP
CT3r9wA1T4xT+gm30j5QniPIE9Zmfqn5Rujp+iDD8yrUTUBDq1AZ8d89dS66uSz+/NB5djDsbiIE
T99qYLuzMPAWZBlDcALt0WzJRB1xrdj3q0oXG7OoauSWiGdoAlBiSvqAPMJJ6pIxvo4mKoo5bzOL
THX1VfjoHI+lVjf29NEIFDI3EgprqyW95agQSuMmOtynKJw3h9iid02VFHjiognuSw2QPz+v/N1p
fKTl8hiXXkMLmrHJ+GWZMMFHJu9aRVTMRhI3L8EM2CsvF2GHhJZ3k2KYlCR3j1xPJsOLqNaiI0XV
spiTjhbcswdQXizQ5xEyWghlg+iwuT92TLhrPS79sVocd38T/TrpbuCF1gyYVmla9R8GfNQDUhUn
yYIX+RnTANCNvGHq0rsEZy4nPvG2RWGRQDlm94u2TB3oKLdXVtvPADhcp9NYAUnZAjOeGmnAUPEo
HtRwA5z9ezJhBzfbiNgwEVagXULwBORpKu51q4lYBHW623Y3rsh/Pl0PYeV54fuwZ/HN0J41ltGD
kQNHB1S634i50OMwoGCbwxG8m/hlE8dxdN+2oEeSW9w+LZvL2l+kTvsVwOo6BfemRIXZ9FRKdJww
gxYbTSa+K7prRbIt+/uZi5cN0hXqFRp51ik0vaADCzTOslet6gTug/pUO8xNK9BMq5KDwarHWFLB
oKfobRorBnPfdoSTOq9/8SXhjJXfgZVQZSme0I6rUsI3DeUtuQnL9l9jMfmiePsCWmTJqM+fO76B
j6cn5KYKfS3PI4WwObGOZi3qETvC8GSRn3YZdahD4YgqKmEPANLXorBrcEWBeEPT2wTjDXRneQKf
PR4XKrb5DjVxsmYdo/nud3+y6rj3OvLRRyoHflj5CMYHfqSTzr/AcqWNmXVLEILa9cfwKlTYT5Ls
jqD6imW7ARgsggyQamM9kd/zoKNkP+aHyBhLokJngzsYLP3UJjI792MZ9+IRo0Sc+LqPrue9FcCF
Us+04e1DsE1sxVc4Xl1n+NMU0Xw+SRfVyUU0/n9+B5J+dg4mrK/0eCFSZNZkQ9dbtca1OkvXvMnK
eoCTBdQX+A4mFWlW3JntQ0hftqz0jTFTJ0jOYG27Wjjc+8v/i82EBid6Azmm81aOXCp92txGBYZy
m0HGKSUdLpNlm2QNUjAkiBnozu+wrzV3dTy949df+VssnUcMTypNWVMgP3y9bAcyJcmuor+FueJ0
xzzA4mbekhNVTCr5FT/MJ56qgzy/sJFSuL+YSlu6S9QYLlLqHpkM0VUM3mExczXQ7X9OYauS1XGg
kYRXgfDWLbJIqvTpQkHko5utpc0LQpGECkKnzTXtfqf2UeeRwsUHwAHJWNBk9LUESi1hi3PRfSnL
4HCcH/Zdj4H+uNnnNhU4EWmU0Fa+x3N5uLoXptd9lrPmaAvb+safc39C87jya11LveLHVBGvQyN/
yHG70dohRyzziVWgHhjhvbQlR4FfclVz9tvhX3gICAKMCXgdJmEfPcJNXw1xrmjZETiWI5tW7YD5
nz1KdLb5mY/GsU7WhqbEqN3TsuOIZpn0boan/phvAGZ2aWABQ64PbB/13yymOgMxiAK8TPnoZ9J2
Jxt8ObfX9sfJtT+ZB3HpMeq/u1AfNDJTE5S10C1OBSzugwqgdEdOz4Pm5D36UOXtqhI+xkUKkszU
g15CKHIQ+aakOGuqQnmrVmDpgFxY6UXErcq4iw/JGBnvjrjrQd48kD69VOlWMYEZ6e+qdyVpcDSg
/NJFwJ0zK7gA/my6pFJDWOcqxiymDqVxQqS5YVN5DT0xjdW7aigb2S2L+Q2ArkxFHL5v0e7xPOKd
gODldCTKyCCmr9SnJNd+GEQFB3zD8RAvHNoklzFVNunof5pQ2hHbchQ4yXaAGYSb3m41h/3a2fJn
qMyP9Okcm9qmZ/6wFlht+NmmID1Hje031/Ba6RZZ+yTc36DOWH+DhgDAxwAmAqs0c/IJDabllAN+
BvwctnET/DP1LJ7ZEtSnMtX9Uz3sx8pQJSLKACGWWpQHhlAbV98h+x3ozQGQ5CIRZleaV6DrcdGm
Rect1zEk/VCNn62VI3Ryah6LbMNb6JBNbWjy8l6o0Ad4QpsyUL+25qlvWSnLIlUxf424rr0B7zXb
2NFvIGEa7uLzEU7Q94Btb57V8wB2cItlGxPPxMwYi6gyGfepdyzxcSR9z2YzZf/D6+8oiNPfM0Ku
jolXwNux8aQ7pFT4homSjS3o1Lw2Z6mlgKpN9s39Ku+HKedNWJKNOoZNbQa4so1X83CktYhAGlOl
Ggcva9m33Au3E/sLOVhvgvPqeUqhJ3jDz7kWSH3ZunVeQMolQeOTarinXOcuRWqTlKzzckGVxd1k
+zlhUxhmZxvQeI8YoZLguoHDm0qtBFWu/AL13DbYBoYbUI/abfTO626gGUs/ltnDKSOmUIkOWCBy
kvBMoJ6Pen5JRqvWCusUsfsnRQOVGQkEf19/JWwms1MG9MgMxVh3Z669Mf5UZKIjKHvnpm2ySj0O
+5IxivAzyEZ1VTFs+ztRo+fbM4A49qTgWlBqCEWS8xzOL/icI6ci0aBThow6EI03hzn3fLjr6eRl
L1rRYxzRJPO99UKQ3XiPRXD6GucOn2tnOBLTAvxApg2qgOLQYc6yiJwAX574hOe0lbjQoNoFJbGo
EMg2Xgax3rJ4pAXXMWsd3O+p9sgwlER5l0om4U2SvvUkuwONjhAN6w/fM5aa3DvAb5Lhs8vzyx3m
GKfZRq3UeXHuIqtxrBjAIHxg2FJUkPgZcKXwPPLSuQQhTcDlGl+wlvEh0vHWvZ8viJggY8ZhxmX8
s7zNTq+eto0QnhyzW/XU/XwplEQGl++GXj8dMtdEWAsHBXi9sekMmIijMwYdGCHRRDBhYFr/L7M/
iChAZVPB9UQXSR7jJxTqztJWO7Wq4ORqtAQKA+Z1si8D1C8l6nG8+TqWG4VBMI0ap/Wy+j5ucW+x
gMt2JC3oGO3wJ8y8HqTB7Vg4V2DjQgw8OcWxCreXcAxTkPcxWZlttWnloj3Hdkn7V1utV86rKTlM
v5UHsLiVkRpbJclLpjfDhfIkCiFMW5rUlrliT8zrYuTAywY2Wy65M3xh9EXwkCwtUmqbgdcNw2gW
FIa62GYSeDI9F6gaRd958vERdHqHEApHqRdQoKS1Z4Gog4ksNJsBE8+U0WmEfnqXCkFtp+kV7rhu
1PmDVlq+9oibgzdj6s3GZQ8IFjNF0ApfcK9XyFo552CQYXSEH/7dluNrb8zXAJNf+LJAF/W3Iwar
+NJnBPCOwz0mskryr7nDXHRAkDxwmRnO8XsuQbJudbxDoas7u0B5Rx/RIVCRDixPfqvZjf3LdDkt
/eP3+Q2kixnk8Lo/cRs1tjewFa+tN2tFK47kv4hICLo0shEtV++RKWD1wQECbGpnTv+fWJxOHJx1
avjaS8vH05tEHw5R4zY8snKs7FMugUIOhDV3ibzuDt7o6XAtQNZdfnp6c+QLD9J+qAKdcbrbM3ZM
qXnPYdYka9l8mgWXKTdBJCQuGvFm6HLRu69Gqxs41k/Oa5Z6DbbWoz9z0LfymGCEM54BYGFtPKhr
3JhOj31ZBcl9UUo/ik5tmoWSR7NbJ3OYgVPFMIopNkaoHJoR3g2GWlShU7ZHRRXhHchSUtRpaBto
oBAgTszyuJ3ORDkZLEFLdbNS7AnW2LPgKNF0uwrdKFA988hFIGsW8DiRDOLGgDKOk5l+cH+ePqSb
/Rta4b/IdnHAJiV3EY68R23+tZPRn9ug2woOeVQKp/zL1/6T8SiM5GdBp8SdXFwk7YYc/jr7jFG+
4G9rHCxUc1drD4n8bqxJqO0W1ZxGSbkChKNKPCeVq1rTKVCVAgPlFG+WL2jn/DPs9m4pAVQ0HLzn
xUAaHza7Lighj8HkQU2UPtH2UQ0mQDHbr75kdBUYYYmtY75HHwGOOgsR+1SIGx7DgCUiANuTqB9C
wtX6cC8srDHRG9zkYA4G2udP+JIzqox4b2Nkjnpn3zbrX81ciLw6TCUQoY2azJfWCCjFFDMlvndA
JGqDnRSHMPI9KRhbBFV6+nOef2nPxrkXRHjx/aApMDX5UCYCLWiFiR7xu0EiuyKiJcuPy3oXVHwb
w205WnlvG7NKLOP3s2VX9DXryzExNJmGZTOr4Hi/jn/fuslYfiah9hwzMX8kjdTSlB9kW/irOl+l
t0uOrMysb2eI4++YwS1dNv7Vd2lYjX+LhlNtSDSvXwE6IO5AhRNu3fIGjPzUqbcT2S1UIudZxmu+
xHW1PxFZTdfJvNPX80t1Cuxq49tCollsvsugPov2MSazj723OPh6cGH2zJmtpZMtrfd43ndukibs
B6h5Z9Rjr0YqSUzf96J6o3o5+Iyb5AcmCnv68ymnkv9wybTQCSYrkN82dFC6RzQSAxZ5dQ3YvUIW
7kpUun7NdkybTNPVOJNcrxjR4YboO8vm3PDIvvrbqJwfeZjEkMJPC5si9SUrv2IlJbs5Yy1uyQqt
Jn5vOIjYxHgHs+P2fBJD2TNDnGsgX0dBX//aat/hfUER16+P9pcCiga45ZdNTzcsFxQ4lDB5KCtc
fNg2qVQnLnop8WYVNQ4oTYbx8XenoHgBV+cEZZqP7TnBanDskvc+ruyToONvsUUnta5MgZ5mdDPB
mIQtczf2Y61S3Ti2BVLocYf6Pkix3XIAnaawRlSqxP66C8zZVfrwkBWMw89oo9B67wxFnEBy5Vwg
wLp6lc11Yd0Vnk+xGc8hAgn3I/xcNly3NJMTKyYBfFEvmdg7o5a54sy323tm7J5aakGYYOrnN3hA
OlTS13OwhCdKVtoC401na7tVhEeilYT06VnI6RxXvreZiz0a68GpUa7lpt1gu6S0S8xLCIYahoma
W3bPgQJIOyt/NSRxULbXsn5pGPHOlQi75JWW39gD1dqXfO3Zl0VcDEtwOsRV5RZTcBAxTfT9oTTt
xD+zvoeoPyPufm3kT14qJNu/KUzbcva4fa35MT2HPx50+BbvCPbR82gSGOSPLEIF+gAJUBJB29k0
EwWAxBP9EPDSaJkXwIzEVxhjjU3ov6OJOnsEY0G7HB8Ku0il4m2JypZPYTRzGkuUgKaSQ5icrjVN
tbVbS5ZTqH30otV1nJoIiu/MKZpBLdk4e6Hn0Q/VwJZD6xnEqH/TYntXtVvgO6HxFB6bmuPVgbd7
WoCMm0gGnGOjjtPF+DTpvfql4xOLEn+ZlkFaPLlKXGHdVp245avyrWnVznx528fB4FiMHLBNd7hZ
Z+xih/3rkNION6Uoak4BoOLbhF0uVKfpz1sxHz9mMiGgVPkTg4H0gnSnZLTNSoRrKqt/qZmUqu5s
pFwAyykQPJT9fNVpm8akw9dXoIwTI5q9FtLOAc7kHSLH1nuytbW6ncy20ZGMPjgbe50jQe9eOBHZ
iEYD5I9QxoM5nBYd/N+/NV1BE/5odddF0QtO1691m9RE6L+2RkoCcocRzI/9Agd3srkxzTssNhC1
ibhn1K1W/0LWRJxJXl0VxJ3ZYVsCMuDiB4tOAJhT3yDX4pFJM+Jy24vex+pqbWMmaosp/6+tcAdB
o1Nz+gPJR1iZPt+bi2HM9N8RSxrpGsLX8M4kgDzk3WTp/riSx896S29yvvvsffcYU2mFy7S2QLiG
ccrLqV/TrI135KDroaeNDWH+Ql3IC8pafEFXH7XmUzQVxTO5cGbJJPKQR42kHaghnwOg4yuDk5Ai
Gf5HstNLNmtOSluuQj1BG9xgR7X+Wz2uIvTfVFAlmezvxDzJw/H8RH+Y9CghlO5fZ7OyOQzSYCGj
fmUY79riuA06kHVg0JfP4mh9ejwW8/6OJBl09c0yrBerRycJ86JwobWDlbKQvaMGxPnYYSekr2aU
Em67WkZzRGLU3vHiPWFgm+Jn3t1mseZiEIcdCxU6L3CqrcUEXLLK8ILKirpua+PcRM9WO/oUlIxn
xIT4zd8bsvwwF7ufsWo8XOc1u71zbHnpeAFPsyypJGQhLK6ZNBm9UoYbVmztalw3qUt1JRvIt4vA
Mmc7m/gzo2XP9J2ttX0HOHsDyxr9fFBVnalvdLC4pv80v+LAHXN4d1v22GjmNL1C0WVA6PN1qKbj
zjDQFPUlcoa4OeIHArhuWHFwec0W+BD8HszMjjhvU6vOEfMkDAejOVgbstGv+7xJyCfW5c755aQL
JPyKCOworlh94k8K6ltL7Sus9mcdEPHfk7jO+pyAMTiphLuRJrw4Jsd9bLA5TrIe05a4A7s3ELhq
/8aMfmUq5WKwJBOMwR7eZp10RCiqHDdQvu38fVveafEd0wQpRkq5mUT3cl5yoppOvS0H2+PNshdh
LsBxvCFQpRylxo0fW4SaMsA/F705UR3Z3RMcfl2NG52vIp0ecKl6B/aVh2S/vtmMZWyDVjFBrGX1
VBwY00x2FoSOzwqZDZcQcTDIwD2Kn7RdqQfGIoJA977qeMxzyP3kVCyOU2oz2GcH59M7UR6jHVaf
3d7Ogidlvkh5p/BdkNQ81XTB9/IsSxPrb73SA46xFJ4rYqUoDQsZ7U3fNcgMq9PO8Za26N1h282Z
jctBhm+TpqtkVWndL8zh8jCJ4N7S7fn5YI1dSvvM+sY6hcEGzZwLX3H8bYxAZH5FBmB0uF7VQM01
5B8l34tOYS31PYQf8otfK5swGGSBN3cT+WP56SbaD3V6j/nIj9L0/j5SA1uCpha+hinVl4Ercskf
JARdcHU4aORVyWQZ6UX3/gpT7Amd81ooZvUhX0a626eKK47+pndp4ruL2rehSskUzXrPbx6egyNV
G0bkrfFw1uP8sSHzNVLfuGidG3vlk6+HF1r9s7L7BLXs94Lamvqwrini1KgLcauk0RpuVUiJ2qCY
aqxTrLseVGtlvK+WU3qZdpvQxYBDINRYz3sq5iqFnO0ImaFCFdamBFqIEnFmHKg2avrvcbyOwgGU
WAD8Xwlv54H8wLt13c+N+4f5fli0BLkC1/0FtDk+yd+W7ZFE/ZaqAbbl7mRoA0t2a0CkENgK+gCD
0UrFIeRLKmysrU1HA2Hr/skIwtg+lf4RHIQS4IgMdEnRpz4KHGA7akWvJ47h0jBfH6aBJafmKBDo
sIZQ5HYHo1dB94RccSkJpS2A/veBHBQxEMjMebOlKgoyhpfmXHpFwljP1WjKLioXY6pLb6Rt4LmR
fnHK1yNIRseH/vK5dDKQ6oT8/lCXAgWWyyUgasJ63KYgQ/6AshPLB0Tj+/Nsys0bxpAgfCd3cFGc
zImAVvJRhBSiv60sFHJ53PltwW2kmL9hxsrPEAfPnWIsXLS7KccRhgvyTtPCBaRrYb4S6EF+T9cL
uULVKsfymMuV/iA1MyJ/i7KR8YLH9c4OqToFJuwgglHohPqVmydQiv76n7wcGJJJTxsjOLkccJhm
oNuAyR18qm01K9jy+HK38SeQT0tjcM61s5EjTnt3WxqqwYB4O9f13NKl/YkYCU3+YeJEwuyGRRGv
v0iuKAxZtU04IXLeneC3zjDeXuFX5/Q4Mit+EdKprs7vFHJn3ejXYhDkkxiJiEtEWAjaEX4dqdmh
JSSWKkziPNZwpsIEAzmD2DRPNGNucX3bwQpeaVvXvdqN2MGYWgtB3Oebhj3uFHa63KJb6Q/ODNJ3
Kl6gAzh56KQ0b0P9Go/LDYBQ3vGCyGI4DTE2JNm+6f3y+atVpLbWwrOQyIfZ8fzPGawIW8Z5T2Gg
+lKlmHpRA1+isaIi3noiSh/zTKHEumvABiCXAcCm6f3tVWdEXtAoz2hu+/sNuZUgZ15Hw2MgIwsN
VmzONyHqpWz9zRrlloDDEdZrwodfa2IcSthTigGeTkAwgr5YydMTscGeyyo82iJJz88OF+mYf1v/
gfjPYrG21xRbMui7kbZ9Oc2Ghk+WzyiCqmhjTa/akmEjatxi5jmjRyA7yAfr79/EGHcqT6vYCp5Y
RDVTCaNkklpRyXA/FmDkGZvBcF3oMdKsppQi0Z86sJwcQZC1jXb8hMIyn9sLVa0lTl7CBWTekGCy
fElo4E2wEddkeakup+iDzYOHdIgANAZ/w5e7qNl1/dueWEXcSpMRePbFXT47FTRPxft9wb0FwTBF
8xwVpJMrxD0LZ5iuQ0G71vleJcOslAc7jt2T+izJLMAECNBq/rp98192SfTQYrJZTFtdD/RuYJOf
rXIWYTc4qKUXpALs9EslqnFFBm786HAftGMd3kzUKgfg2QKvX+F2c/kwgWB+ySKU1U4PSFaBY5Qk
4BQDwzbWbc7gVaYqy0q1psIhhy0wqRSjdhSaoGgS7IVyTsI3kuj62iDuSs2/m6lghCc6V8qx/zU5
MWYfi4H9CwVUjgr+6TSs/2OXlNz83R2GJPevEdkmJ6u1LN6sZoXWFINo37P2TtklIitf1xr+VAHy
cb29Jk3hH4BaodlmnR0AoNryzyX//atso1BVmPgRJWA9ju4Q7zF08YtOFWLDsllw4yqMMY6uK3Pf
G3tJvHltyOGbmDifghuBwLrJh6Cwr4rxT80sEVaF6RAuBXfYsVI1U6KviL5C2IOcmmGaC2vdbA/r
EIDoIWIPjho/WLN3E2kAJCBj6aVcO2P/H5EwqSwd9bKO0lEEgbnmRVZvZTi+3crKdksFdJ9IilIt
uVs0EHcj4NVqSOGEN1daW6RBYhgacI4rHp+epWieEGMbkbtKsViZfgIgd22j+8wxL+ktABWCPERV
9eUiigojaOX+FVQ+hRubEtOIjXwKxxKz5E01Ak0UqNEgBG2avVEcI0zlvuAM/x2y+V5fq25n76rU
JwwgfQKDTWrRsatK3o5FKGe+L36VU4MAfEbALhbHCJyuadY4PH5+3ghqTO6VB1KIHG3gBgdfgDU3
90cG65hIYgUxEBr8WalerIE6VcVDFkpH6QH24GzRohYqoLtjKzavwWVTxkZoy0S+rMad92FF6QF0
2RxNNC9MqxlJEuDQOxvTt1oyUu0JPY/xOdRQb4ZQg2ZrmOiqk4eA6r1Dn+2cmndTZ4ARiRvEm48F
VZNZtCrL2GlOEZGH1FUHlNVgUCT7uip5Dpfvs30iyhkbHcnMxhrMO6PCTx91Lj6M6Ku1UYqNaMpJ
d8unNXhcCtB6FMGFz71E5PyphII2QtesTjNflHjg9tSPj3lUIbonTbhWAdKxpdAoshy3RfltN640
uhZkBcAJoXVzD6isqF5LB9gQ+ShMUfJ0QuIs+K9eiaZN6DUOorLOK++2nsqNL63o7Al0GJ/JdoyJ
FlDA4P6aA23nOs3g9lAignsOSOg7fLKOQhu2Xq1SGQWLNqBu0tvvTVyuVOdpyybzL0ra4UV/6SH+
EUZ+Mhi2eDjtNq1jYmP2TTU9qg5UPjeKg2mjRYJO4wwEpcTdJN1fSfleSz+Na1UwjLunHQqR63XK
sd7hp+IOIH0V4WVoCqavFOy9gF5NvPGIlzI0MXusGgGRK7/V8GPTyV7CZ16B6w1rn856NqLcElJR
TlExfhdMbZbxwX1PkQq0uulLw+sMlUjyN1HLWnRp/MXIHCFMIjC6JyZ96RgX4kEBh0WlZg7d6Dkf
Yiir0DCXWWnTGvKuC9VSP9JHUMyb3dZ6w8fkhw50e7emnwa8ExmrVL8FRJ7UrD8zHEYBEhcYYlD6
qcLw9p1cINoattTcaicXnD8oyh8Bh67ou2hGinEEdWNKxDFS6+LKUvGJWEGE2A/dUBrkRxFJBfuN
1LVFn/EUq5nRLi3g5uClkXmh8k/EmAtv/1cdPbu1XTcmjxRcwqWwzjmYibL9qc3ygMxjBtYLwNzw
MN4JIAVFq8OQaffPCJBXW62En0kxYNZyZAHQSALBmZUlf4cKZJaJpytPSR0BvOX70CuKkiB1VrFt
9zwVU4Hi4wJe4r8H3F1PFRWiM4xs6sunzfeqHXT+Q9ZXgZCGNWTkjTn+q/mL1Bfmo8U7CALp9MlP
BSOJIuLg480SP3HW+iaQR72KJcC8bT+mgdVIMAZ268y57oev4NXpRJ0vFv8goCj5jPQshhtYGmZf
LoYJufODh/V81ZWjE2YL5cwNl+ljtNDKGO9bROF/mi2Rf7gMsypwvNPa/tlV/87f2FvGt8tuRQ+T
/SUY0o2M6hyCPOQ/oKE9oNBKov+PTRsdHPE9LREVdCF/A1qffWBOAy2gpplVceSN2H92Rki6Fb9C
gUMI7ScH392SRc0+NKvGOmMIWzlFEfdM0KONL7cCUVUCqjk0s0+KWFMcD6ySdy12dCq63nQfeom6
ip93Lba2jWUI4jT+0/dPesTAb7ozlJexhy1HC1xgnSV94hF4taEVi0dcrKQh2YrSYc5oyf7mYj1k
i/pmdrxBX+MTFpznQUw+wYaOXP4P1k30f3keoBTIwlkQDD8zyomA4aswcc6yqms8AII1qGQD5sc5
B9ziIRHv6S8mXi+BXuBIsGmpCZD3ebZgiod6mc12klr+2reyQqRi5OicjBwrPKNbeIphyje1mjyp
3dkxhPlBbq3yCbfiQ9DzP+QRhfcX53V4nPrpFa7tYk0DZOBXRevpIL0Dh2UdqlgyDTsy9ULYwrRt
sYbnMLrTMbeUxgbCg+CJIjcnjoDl42LfG6GMncYdm6cgqRGdnfDZp32nayag/QVV0A3xjM/Z5308
iAbuf1lGZMzFFCpyBLm5zhPpXFAs9LVAujpYRsouIT2cnlz22yTRE9Q9MCNHuhM45GO4LX/ac9p/
7DMeQvlU7xkyq9qjjqH0LSYW3oXWaAxKk91aJk+lNsg0mB7ADbQRTRmA7JdZr6jD3nN/KaGMu7KU
3sxXHIL/dSmTTrAYoB+Xa2vbxZTvm3Ancn1NxAXCFlZFtjvJSokSdBa6yzn5lO7uuqx8rLaeuQL6
Fo5/2FxnwLtsaIZVCAZV/zvJxQt5tXBegnoNiL0X0M1BDlZhN0O7clI+mxBmvBAhC0hJzZZeTNfo
hXnitllA/VOUAVNDaJn7TcWDVX34dWd4oR/KTt15Dx72q+HMbq6b5VIiXT5mPiKAw+bQjYNHFtJU
jiZ9gH32ECb4SDYCnN42EQs3Jhs1fzQuz50qI/ByLRmI77LrYQF+YpQGjrWEJRbhu6YjsY76XvUI
5BMjf8rI5CY/DIj1Lo8D63hr1Rg5pKqK/L87jktKkItIGYqR6iccit6HEMXeza5WFtvhTic0uC45
m6MNF4E+pJdoPIkD/vE7odAIa0NSTz4VAxpPqXBNM/febmUOfyGjYfVZ2ElHE2GUfGhjuftEeJwS
x6E6nTSW6cGC2jwZ3QTTa4NQVLwUnLPN1XO/+r9pqg8Mf4OPe1kij8v7sEhrVpdIcRdsAbjjNypx
syg4s/cUp+22WC0Lqt0GL36RWbwFyGRbTnoPt6gbToCGo2chnCSojYzKTR9Mv2ILx9Cmjejs77vH
widR1tYNdJp2OTExW+bfTgGw+eQ2i2/daq+GOuASDqlsxsfAXY/C/n4k2QltWx0XJRxsWnqFug0u
YCaebF3ajuKwjZMtTri2PspFDs6bUrd30K3nZivAqe5p5g58s/zaPQAs9o3aLRnEjrG0sAqGeUTC
nbFnWNbOUULpX+KcFxUnlnv1Is7Okz6WqK/bb2fR6DwkIDqy3QqhR85e3mkbKf4tcQijsmJ/wShJ
cv7aGtYvH4BBhkujLSgBe/UC5xyO0JpighfAI/H932zP1bBHFtYQrsdlqvMDsE/Bq33BxyKD826u
ReLpMkvhtDpxgw7jk5CAtnyhOmpaQ10acwVtpG+ovDkF1eDF7QLjVmvMgczZCEs2+r8OVl4DLvjw
5LHMldPiChT5ICaV3MRLqvfb5L3g9wX5h7Uhbwtmq7fW3nn0nay0iUk25Y/Mf9cqEJzBmLDi4p1b
SqQMuu8pq7an+Sb+kyAl3EQvxfAM8yUhLw2q5/A1PhsHgzD9odi1fcPtjBjMJ34X7tJvRf7EWl4k
AgaGLlCGgXbonFDIWVWPS/pwthqfSQ3ZYHhVSblYLm5bweQGRTNWAejzMja2LF4N++mihRYK2kmh
drLnInmar1zwck8o4wTnQdgZhx15/o9mWRGJkBRQ+bWfw4Fi7knb6Yg93IeQpXHYAmr5Nc5HqWL3
IV4paFNxw4ls4luVruXRxRlYRoQs2/aC4xIl4s/ZrWibcqwJ4/GJPsnsBQTRj6WFDm+oDrfO87aU
+9U6VczHLQ1KGizsbrD9mquBTz6OY3BdKEHjOGQqBrjm3XEEq+jQ5SNguWTemWBv1lpBUAf+qHJu
pQCI/iHY5jZo+XfB+cET00EQwvdmGQn6TQkSk2ixjhKCv+zn+yyDM1flJv2vRVrX6axTQ41xU8+w
GVaRXlfhzAER7jTnsdDLGM96jY0phdnIYATWglWn1yrGUmDUIYNd+UNGqiRPBxJh8q+T3TV/2S5D
urG0EJ71McFjGWGHohSuZ7rZhWbOY4m8jOhrMu9x4x9GPwPKLto5C6T2eYqndWo3Q7YUdJwFX4WO
TtFj3fP4TYDr9qeOnEYjmfKqy0whaHBHLYQgoipho+0y7XEUxXGo1ys6A7CUKHDbaphcePK7Iz7R
nv2fv94t8E5wPxlEhub+q38MGSq1zahBoEX+UGDsV6RsSO/JZi6BkQHOkcxmXE97zdfvXfe6qKrS
zLTnN4cnlDOou8BwAir5VLfXp4/VHdSh5+fIfMSoBT+SD/QRXAZdG7E7NjEzfeukxh1XROqXcQaL
yqeBn7Qvs88C+OFGy8Bw3WVpNhJwdO1LxzzrSWPJOBBfF0XuRc5Z3bjr8qH5EYWp2UCDN/YFPLcs
DGn5L83m03FyVFGYmk+y1i5wVH8ut3I/Xq7VqhmaGybHw6ZqDu5GEw7CTjtmlQ7Hz4b95o9QUjkX
rnesn5yqJakgyVAxnipiI5MM8gmVUMzul4gS5XzdZyssrNPCKnT5x86ghXA78gZeBHYQqQDs7bKN
u27htIpuhBGVUpTv3S9TMxxjw+beycKhYKerKwHwiNtQe+F9/TSJ43rLGSQrT/lTMuLohOl6mM8v
Ddis6X51Q7RpTa6j9YCHJY8cgn3Da2IivVwVPwib0u6zBOYivoXUdXf2SJaCJ7vWH+a62jfS0ZrP
t1dStXGnRtY7Ppb0xr5JOtyXDeo/Rwl/CALR/yYyHfgDR8MEfxMK0WhH4vyp6exTEVU+MQHi5FjZ
3UKvzKfub2mtJpn4a+VGa4nqhjPGvDH3QqMxpSbbUdqsMRyRZZOFdYQw8CvZLfQCd/r79tLG0cFZ
0tg8jEANLgK+eBYRaPH4vmUgZDGW/jAb2OrCGC/52dMBDobHtxYwKpAh1az68oC0t8kUwaPgxOSY
tXAd1bq6FYSDPGOzIAzEiHw5yqsgncfTnsPrsskUnFeeCI0TotFIWFd+g7Y1290vQcKeFJx3svGu
nIYRF2gN7At5JgCjo53wqiZfZq94F1JGkg/Bui+ZAdad8/aYVblxa8wSsBIhNZRpbBUr8Rq+rFa4
5vnop4+lPQvWEL1wX11y28eJJy51MAZsS3vnWkJidQ3zwV0Nx7D07HkzZQcD0LkYqYKgQd3FiwiO
/I2et3OKwU6sVIKsgETw/wLR0hw6JxXQ5pbeVd3kEEJQrHBFW3vFgHTUYrRMpmC2OpWPWmZlk10a
O94/BkMUW0HfnJ+CFs/yvrj6rqbYN9u+HXKqGPXRc7Ai/G9gsoxqHI3Ie5QIQOlhYsA0Vfi7ki+o
BRvX5Wgv8WpvxQeFHK/khwpyfgdWOnm1vqzdyrmNd6XTMEuKGkh//0x1BoyYXmsz6w3TcUiZkEfs
S4ywY4zRyDGSkd4KKVqrwaGNpczt66ciYmSR4mYusXEJte+WgEoVQQW20UpNSjHYEWo78GsZW0Eo
Ms0y9ZcQRKX1MIQBne4V7A1qepEX4b/3zeV3OfgOaLikWStabAAMV1tCUY5rKU8f7S4qm45JTzgd
C+mEp7dil/m8kP+DcpR+IhYf/p4gGHDEnVIhHcMarxgguc5bujT+7k5wE28yxOrBI9ujs9sFNzG3
46uYqW1N0X5ng7gtEkbjn6HMpHMbgkqy4g0iBZogc+DR/fvlxUWDYDSt6V4A12LSNZfPzNmuc/gs
HJTJyRkHOCljJQJ2rfP8nRLiHDgr+EZrJvOYo4lx6mocA5TU132eqguHfpAbKIlt6w7QBxMtMEIr
Jc+uS56TYZj/vR2TdLWsncAFEy8aIm9d+66z0zJjfZMbB/kFdGGb4wajf3gLRKK8UMQE/ZOs2L3X
/V3tBR3orVn3zAIknjjKwvnhLMy1SbMlSSzXjRQHSnBR6MEc1tp8UJnvj4zoJS4OKmed434J45b0
ppt5gNMWht0TcmL2LrGo8lJS9yrs7HrXyAbAc82Eb8go5OvLwmPwsOcHrPEUE0okD54uWPeEQyZn
gYHphW7j1fdZ1BPbUA1bYlyS5kD5EmGpQ4UuoEGif/XUs4t36O9Il7zjcLplPMxRy85M+kDsMK+B
NkYSUrNAbxD8pr+d1z/5MAmD4E9O7Q8nSZCq1y5SZ+N2Jp+gj0y1hxuQ+fIhIKujYjf7/GAfxv6r
CHQU4okg9VwhbhZDC6U561jrbr84deqVYDPcV/xjg5wqlGBOpWeUh0ngGyoL0LluGi6eQ5fTCKVA
KgkDch6LPKWRBj9XG5HkuUZKl5RQHr4SNQqLoupE1YGH7QcOL5gZlSmyvcSTsTSICPAtRsh6Cgsq
XoPymoNSUzsAhfzbt6BrmhrrJUDna6Yxt5VaaOK3cSRignDWV+kp1dZjm5a3dqm4cB9mwxEi9wNh
a0c/fUnODiYf0ydLBtMgYFopnVq0Z5g3TqvzA9w0v6Am255PkuAymXNsY5FLndAL/+YHfKoO99+1
O7WTmWoBys4hodx2E6RYiHRSocldtkI0Y0PVeuNpQ9CHnxrgQLfeMMALG+F4vYcJ9ZHylpcAOA/1
qYNMVdHlJUn3QGTSE5gK7U80tMgj036+mP8qVETQrcYfIsfYgqQoieLWGPWxFojlJah8apjqJ2oF
Uoq9Yqxdv3ctZCSIZ6ZHf85/0AVs7M+7eWP/5y4qunDZCcGHKCwG2KyEcgaFN0ZlZClhZfQrfElG
ZqqrwPP3qu+174NYSdLXDk5oXeiXeh8S3l6Ui+9XSc716RIO7t9yHjDYKPTH9r0gRlIl80d1TWPd
W2LH3IbNXhBXdtkpiCxwFnpEB0B/fiF5tmtjIMYDlEtYH67cQptZUpp5UhFu+HpgKJSliZaWtzr1
mPDXg2Qf5QiSKk8vnC0aUHcpthwrivSyos5Ch3HK70p4hlxFktWJzo6Cm+vDZFJPOCZrIWlzR3xt
hMgWXO82TyrEAkpf4yF7WY1bkiwdlVhMFx6RQqnDD/OKGjZLHcKBhrkBQp0tXDHJWSF7Ctc7J3Ye
6pXI5oZeLCFCwXHjQixRLyh0VA1JylEOVlgm8mpzbK5Zr8q7MfsT1lMyvNJfVfqbiHmtoE/NPRX4
EQGYk4Et8ZcwZD/GVzADGmsoyMj43JJ+DpDk9EQK2yTkxssJ04rZCHrJjo8k0lowCRUP7WkIhAd7
1VFbXnP7t1NZRjLm62SxbEi470cDi3LZNmhtHyL8OXqbiLRCe9359NMI8bvQPdbzklfH6jKl6q8B
wE/gl/rdgx7f2Sx1l6j01e7ZXmfVHZk7QlgVHUBAmYVeQvkoHLvvm2QZLQaw4Y/r+MN+xF4Ykl2S
a5zEyAoxeOb1aEtOC35yzAZkHFu99teYS/sPM5kJXbQtyiIKz6yKNXbijSGD8dJFoN0Issp+5+Lg
LdlMWl8OZLQFRHem9o1RbphMeuBYn/Unc5aTV4GArLwgDNalajfIhI27QhEVn+3uKo+0TYBdHibw
nqAkfQZpEgQGugjZ5a7vocF4o1eD7F9SGGdbwRfpYEJ5mtLg95QKcwrQ1pXPJ5MrSfnmxB+1bNX9
MUtDv0Vl4j9k+8bFTNtUKT0GpYJDyKK9DfMS7fOHBEN85aq6bav5jov8fepmriFwnO/6tY2yLF0S
xZYiRwF4T7AytKegX5yvISEKvI56/YkpvHwT/sjottl/4f6sPJA9u5wQb34hENRm6zvuIfwh1DrX
JWI7BKDWDs7RboAVBZDDZ4KY57QWQB6H442BzRGqTdR0FSXLvRxOCLN2CBakvNgEnUDSk69nELYR
cM5ASWAABzsM95eYvzXsITS1uzT7hqTAWt4MexESLCSzWqsL/1d5q6dTZ3CoNMRG0aQxbYdAQTvC
tpjZQn2kBuO3ph5nwPyHYk8EgvrQWsE0cW5oe+oQ9TyIbdamayuQ2M7voeS6f2qQwYvRA18q8lYm
PYYUnxYGhb0J4z4zdPI1Zsa0Cfb7HtA7EtDfQRp7KcF2WkH0kqUtq5ubmroRzw5xdyyMsJOrj0TM
4sOPtLMr22+sJVSI7XbuRUEGh6/OFWUWFfpBF2C9+b6gisDgQMob4xopryq3kUOCeZgaNrWVkkRr
2eBdmC9HyS4Kvo0X1FlZ4YHlHSVzUW6ZAZ378eLFvYdGdK+jTkaIUC80c01m1gy9vW9sMfK+mH+8
990G30bP6YmmzXlfjqd97Cg+G1mrfOJNONM8L7zMenEYiHm7GqKc8UsRoBkmEsRaha5RCAQtcP+F
C4Cg4l4LC5Ec3Owm7XQBtN288/FZSesVJsY+/W9xk3g/mWVNCYLnYXHqde7sWb/5wGsPRBIGyadp
z8IcQbduxuAz/UentakzmiCfex8AtM39s6lMyHiuW/st+QGMlirrWpGzagn1ctMg3ZFn525KYmJy
tHmZLXqsUg1SdlXGSJVtfQoDjZhiPhhegtTIc9n2lWZK6svWKv82o8BhC14aQNbljaiIAQtljG8Y
KhMvvqYADGrDbVhCq5d4rThfQ8IL1Bom/vIRwYaocGG4TNV+MrVQA2NjYvUzF3H0payB/OHUtyda
kQIHrO8O+ZsTHuJXZDXKrxhoI1+Lee+HeaoLcQJcMUEytxMiNFgZmubyprxzM/IrwWbzVOTbhry/
EQe9nXAhrqrKrcISAEUl4wWXYd5ROUsFTaEyOl01RwyzagMT4rzP1KMXYVYsTRlXRRCJxu3x3Fir
z9FU6YJid0rpv4/ul+fBQpXXsCWpzXH5pVuvXCJI1lvWZX5QxpgmIeyGX5IRbw3MmTgsZkUz1oAQ
DwB29h1DtXjSkq2rC3NM2JY8wJ1OKyLTXtizx4EOUgh13g5YEcN87M3pWJ7ZDLOILDqI7vtd+iaQ
bSahDfWIoEQqH4boCX6kiuWu777cWl7eZKUZqVl7vnzQOdZY5dG9TsH1/q89ZzhNXECSYQUyxUYn
jhzo8AhzaPuBVrEdO/P68G5HINIg1xWgqDbNFJbMAjVmqptQn24ddYaK5QVVi9oLXZ4lgxSO4B2+
+GC107LVF2PBvjrIH81wc0TTIDjsPMQEySlwR9Cmt5pf7iCuLxjolSOxKnYjjz3PgRd+SYyuzDr7
Jd8viCm0fyLcbvqJ9jO9rSJ5rmbFYqVBeKDjYLlFHeiKps7dGb0mV3HOpeE4RJnZdlEODFPBELuq
29jj5fXLsEkZA7vxehFcyxDViX5D1FIqfSEiYOVCbYnrkWc4l5DZa4WDdlNqHM9uTpsWiSbMRKPO
28/Pt2+lkI2ltyKAa/EOSk+WHb7QLNcoB9Uxj4Pp71MRZ5OzPm9IRA1ZaSM7UpoWaTJuH9xAUi1Q
HIl255+IAVkBSu93jWdTOOKVeug8HLaMp706wQ/y4LrM2NLj1jAMAbhamhHPm6/yw109bhMcDoYj
+f1lqS96oATPk8R617yRLPSfkMcT31sZkWg2bXn+Ib+GQz8SoTdR5DRHMHerfV3pm6osq02jGB55
nmfSiDfsvYlMT6LvhAAkQD8CMs83kH84SiA9kEtnUkEm7+8gX82ik8pr+IVMrvmTXA5BYoWTktaK
VTz6VXLwSWVlq2pHZQtAHPMgoAV9f97RjIQKkUQQtTSgaesiJodO2F4zE07bzzpTZDjXN8/iMWIG
lNix6x1+elEEyAIc6Nq3ijQ67EnCiTUb9iEZica8Mx0rKXhWF6elWw2z5rO8IpInSGmTIQRIKT3g
jdMnKOVLVF/hUiQF6evB7U//Si74dLQr/Bb4Scg8xtwbGcMTUgCTMZ7TCLR6s9mlezdkFIsAoJ+k
sjNf8vN3dzsx6MkQL9NPgokdLuFTmqiC5V7r7IpSCyy8uwEBjeN7Go0PwwJ2Ua2bWesrT5SiS/1+
C4W0k/5OEokfvOmqQFWlfeWwcLYmRGkosYu4jPH3n0Jl0EDLMQCOuYmbK6NOHCLqmnGNavmnPkEz
B8pAr1MPuOWBznKsecOwfrlirpZ0KPENHZxbrKzdHfn6EpMghllqmq/5TKqASKMOZZzsrxljOa7/
E7hnXmC4JXI6xSl4oTvWXSbIF5nbIdNENke5nhh52RIj3+uEx9/XBgblboi54pelwlI+aLxLX8R9
cMmKEAnMUnvWe8P5svMPe1bL9lrXEvO5IchGpDVZqzMm11z/3ch+3SVb7dBtfyBwxn9gQe5xV0vp
C/vsD4zSogScAYDsouiCDox007dBUCIuTLodK/LLUaVxL8n+BwY0ZDVhHp01GLgo1/46mRgHRGwV
Jbd7aGuUDZMyEqdKSuQcUhiWQgZdvrTKk9+mfUz/pmcAiXUWIIW5UxnU8T0sCwWRpTaMbDq/Koei
6PrVdoaUIrGwFBg+sLlUla2yx8ezptZngOexgPlDfKmYZpY/hPc3kVooC2H34pPDmIxaCh6LZ+RA
tmo/gi8INRrFe0qh5+MQOq2/LznJEvaG1mJYP/sUjRCZcQVZ1GzrlUcL8Ol1EGWZifR67QSBXLZu
uwmaRu73Q73TuvDS6NZZiCvPd2MG503ifRuRak+2a46nscGRfUqPl+VkvLbUvxyzAHdw4BKhdnjz
RQLxrqGyRgxFEwkecOBdqTBrz4chRrIT8y2lUHwGoKJIh4/BQ08Z9FJjdKXkwIfiihLQL+1TFMBN
K3TUtK0Q0fqsftNer0xKK+GhnrCSEDRXMVQjMEOm6VUOl7P7+YOzK+f6uvliQCp93CW/VSqGl7JR
wfuQtqy7Ho0qM0m7IwFxqrva40e7z/Iddq5+KjHTJgMaqDeslepuQ22h8Yy4sGO4/wOFKlsE+FFg
qDXrXyBqE+YRIE4SMgd4FaJdDVESZzcw02qXZFzno7DJndaa+iIo/R+kakZi1UCJAqrirVCGUJVz
nVni40+MpXOIMsZiSrKDkIqgPv80IHJmW3eRFUbZAfAma1hcPZ4XT6OyISsclYpQZdFDTcXttKn2
seZO/ICudvxs7mlpi3VX/73FfWY2SYjvzWr5hrafj9/r8WgScVwaZnuzy/YV1zS+rTjh+ZKv4qo2
jFigeDFTOuS4ncC/kuZjEVeokaX5iO+VnGCTpsi4HQge6i+AGMztWi/IDixR9V+8dcM5ODSaAAj8
klO2i3+XRjfMjVqK0bivR83QKOXXOX6/hz6F8Rk7c5nBHI1jLqGNYD3k3pUt90D0Eq6wAW4r/for
A/nd1cZPrGljZTf68syscVE2/4HvOWdAQuyRAyqj3pBw4KPHcdZ5CGXPKmM2ePRmIUEtlUpZffem
lYkcQNh6IxTUMppFaNrjwe2WtF/lDOpU1jLygjxFyS9nJQD2hhpjhNZAe+82LFlSAOunvzPhyymw
axr8mvuymAAcDi71AaVgyjkjJEGa2OLr2l8NYWvYVaa2bvWk+3qnX9I9aAr7buFGrzv+BIXOVXYU
y81HS746sBQyq8FZLBEVNc1Ghuc7QRmfVn0HPIbCyrnwnIdkuXzikn8j+aqR1gUFTrG4AzsmMqxN
wtC73FOQuMJl1YyyJ02RsfX1oSEMMUNXIISnhO1QeybwUSFzAXXIRU1nljfNjaXkYLnnPdngdAHx
bZ0bvOJuiOLcTC14EqadPJ2qwMYChZ4CG2GxStmbZ6fdv+536YORh12g1PC8lvCGmn6qlr6pF3/4
vyY6HgIZkpk7F+sSu5tXGHub1BVBKvQEozDmXDYcS2Hyw3FwQlEO9FHtx8oyvb8jwshoOiFkbuey
Gj4CDHzbmfksZzM0u6K+ZhBpHhQK8YgHPlmcmyJyFV9Uf2wX+wTr7IFGkXcaDimQC3F+pB8Zw9D9
3YJMzstW7iRsUa8c4wUoa7xDGOoUHF6We6SZrROCrAoo37oMh01cjB8BIfjCPTO1UB227gzWI5ep
1AuolIC6Asu/7Nb2YfiUoTdJz5gOpyxf4/1cHA7W2w+G70gbhJ5UKYeNO4vZczBlE/QMXYgVpVD/
KfJtLEp+truLwyJk7TRRtxWTEbIJXeR83zEJjrxMsBdyHE2yIRZXZ9z2R4G3+zuEVl6NKR21kq4O
VGSgdFpQ4uDXW0bCY/aX+YR23UBZKX57YK/dIPJMK55mtwjueLoTKNTwAl8ogZC+nbqPnBQCz4bv
YGMjCEyCB2Iv9XFMyp0UNagggS/3qr+i3vM1F6844Ec5tuOsuhvXaLpO84Opzi0qQyCXfQGcRy1B
co5ZmMWCcS/uxIyd/aRcnTcvpY9vD0CKPI0fy2OOtCWIVFiIoj/poNkrL7z1UMgbu4GksohQ7RLl
GSpuC+8yJ8fbqnZKiDfsnohOx+5sundWZ7YF/FlqlbKVwTdGAgcByyojWupcbxX0muVny8eoR726
6CZJei7bAYcEp11J1DRKnd0XCh30gYZsHT3ZiGRRMM/2l0E2DGcQZVhO/ptgHnigLatnW21L0PXG
WrBVB6GyzkoDHc4Mf/ex7PgwDeccRpaBZ0fh6Cmep5WpefuYblxPAHUj5zEsCw8qDXqSsK0KSOuq
UDTOfaT90VnoFe+MnIU5Vj26eDs4N5yyW6U1tGB8HhxXpJ4KpTmfohfXtEi6rMDsFDqD34PzhZ7o
9emzZayDkyfiqs6UpcRfnYL7mVBJ61s57TYFgSRp80soaZkIZRWXQQxqlAQIbThokNucOdjo5g7W
6PT3lKyzCpNTaLDdDG0UhJTJLqummdsrQG/K1deP2+yniPxibKwBmqMcgECWUUKdoRwTy5ClMNgO
PjyI9uWB+qeffjMQznmMICUFWfdnNgGSDQdEz0cVsmnyY5PpsB69pZWZQAzjm5p8JmkPKxF++aKg
L+EnegQ2pyuZ0J8BeaLgiXcUXkrM/NEF5vE6tkU5vkcJ99AQv7ZwmEXn+zAhegyK4wnlv3EkRxnk
eto4eCgmw/7vT/KFofvXtijyXAYM6avEImdWVGVahO6wcY3vUH62sUHbGXEnVgKPPzQxr2NuV5zz
hn3Ig011Bxz5hZGXwmI8ukVVfTywxnNY7ia9LKBzQo18fxPD6/lvKbCJQ4U2I9khsoM1phwitqTU
AwbLEH1EIr3RUKfy8/2nr4hSOUfGWaCohS9TQrqNupsrAphgMFlIpNi3p2nydWECd7Woi8tWZg32
9WcKxMnygxTq3yviFzgq/mrNAZQ+7Sqjmmpwv/W6a+Xb34UpHKiSdnW9+ptSfYC/FWLnJxyfFJWa
PQnXwP6iTxiqBPcwz6fHPnCv164iBoxQ7DVBIiY06H+GnWEveJ4oJMSSPLi6c7+ozRhE2mQR3BNd
t8yauWFETr2xKtcfpXJziv4v3yX3bBv8Cypw/8a1aUQ0tVpcDf5z82a9yYGWQDbL+Jh7J0hoaq/3
FVgD+a3oWy649thm8fBH2i+XCsIHiUpvfo7US7S8xBMYoRzMYF4L9C1nBGwj+U5UpLI9Qe+Y72Zj
NZnoVTEvFTMZCBMBne2AqzCfceqTnYnK1BlcYSIzixi4pYy0sES9JwmOZKciGeFi4oIbroyOwoMW
f5gFxzRHtQUfX8F4OHAPpJwUIxDrOWaG82zv5NJX2XDe5lSu06sV3ENi1F2wOmZC6+KMQ4cAlr+m
G9lrUtrLlc/aUJWy0vDqSL1RIpTlrwMGHjyVX3/o6ChbCn3isdtvMK76xMmUgvGk6dfS1ZjhB6N6
rJfVSJ9wjuh38xv5QOKLAtmuE73BxdOBJr8gQ548H2+8FP6Xu88Lq2jd70tdrRA+MNPhc2vBRsHs
X/L7DDGg/mBTbQ6K5MPghiAR1Mo2gD6areS7UM2C4I41J9js2zTvk57i6NzM9eOn3IjQFWO/VODK
UDrKJdo5P2yh6FOnhnj2bSJ3tlsuGunEv5VM4vHHpAUB80rRozdLgu6I7HjtmOX0o6JL2v0DrhQH
KdGt7DNUyMg+MVUz+BEJQzK6YxMADoU5J2AdC+ZZT/7mM4DUpKykeZN87cPIaG5bqz+wV7oIWZOS
vvxU6bb1Yhni5iHpyKp9PSl7X/wJ7V4RCmRtyJf687KK5dc9ChxO/HVMsnnLCFquaYIGwM67UtCX
OZOb3y/uHFd3rYW2bRnm5iiHa7G0rv+E8eHzDw8GlGdmgpnYqqNsICVtTCqcM139vK1R5IMnvY7X
S470OjUVmpwTc5vM7JXJSPZhryeyOXwhS99JveFELjL8kPjgNVpglPvMr+7WvDooLDY0i7eZibUU
PENbPhzeXKIDPE8d9jD9H5A7GrI/f7H07Sn1ZBhXpI52Xj22SrI9G4GLGB+vR0Bapd5i2PVNeKca
YPNCCOqntIJR9yrochpfU+msPQJqvRTC5L6lrJNbjd5AkEZCLK2WTvpnX9zdz1zvgCIBT1gm7Ow2
px0RCeF760Qg0po0ydxWIWda4xw5h1eQZ0+0wcvAJzHmmCCn3EbuKu4VPGnczfjID5ZSG7/b7VQS
I/cGDf6P7e0wFoeJi1+heNOxSf3xvoDCABtgnmWvLzCFiWqF+e/q5l5oW6tfvCowqzboCfhd69nL
c7ArpWiS9BwvNeFK0jzUnMPTkUtOsG7mCn/1NQYsec8ntSsgA7TkMGGRDc3Mou8+j6j31cZfAa3Z
xl2Q2iA0lEMsIEgWjYRsx5WimzJ5bwv+O/Wm1dxcIJfJ3SMTK4MvOGr8euALDT1kV2W6thfaNCRP
kaHIOPpe1my8m/5oKnXOKl411zeyRO6d/wayCXuYNUbKlIFr22tSd/zuoxyryFKCuSpb9/C1cRtg
SRwxGdJK8XuXzNdpe9BnoEPAj///HyccXumf5zmOsp9kKPpkV1lSw9JPLUJSCQUkZN++TkFF6rHe
rVS7DdcyPk6Bn93lw2Ed6yZRnsC5b/nykvtI8CBofcoPWUnMXJo1PSlCjImshOTqyc8HoIcrfiMT
T7W1tSbaHq6GpH0T05o4Lb3jB66WOLaoOj21JLnu5KQzo0/bBWlATUnqPtarx1BxEcJJO/RlomUV
4txIkYRByjHTsmCbZGBBX+SX0DQDCL72xFpe6TSkgmaHzYTE4NhxRj2+Q0s5MM1W4/zovkZhG67q
+8+7jbe1/VyakRte104CHL3LPmvGUGq/R/M368LV2USCwIhSr0llrpsn4lafqZdvg7kcSY7av9qd
0yYHaE9O2n3LWA8u0O7S/c+kJBTcKSBVYHVUL1+KBnt5TwXDpwz2FGxo8EFbrvP9XpzhsA2297MN
zqaLeZxtP+ShPlk17nPtFPRCIl/yqjPymERExS/uTX2BhQCPW1liLRrP7OvMeZrZAcClRNIlJ2DA
B3umZHr4ijRP4w3u1z+g+um2/CDdh5P8AR4Iq9cG5EJ13kbmsMaytuYk8lH1SGgoMKuRDNWh7A4F
12Tlk42ezPF8tgcApp9M3cdCgHdW8N+fROVPslVPfyvF39GJZlKkbp4Ii0FfR/euioVeVMTBYTY2
JUuK/GDnkL+dU/TYK+hrr+DmwdiaNzmElcIw1UbamjluBolk1dBdF97Xw45RSCR7df6UIYY5CZS3
dPXZcEvwJcbafUnSv0civcOFGKxWsVzquORUkgbiei+8dnjAUYN8F/R7Eam4r+V7w5icfAPHuXi7
z+ySO/L+CvA4Vl1Ei4MKXe8qgPwYTfcsOldXuVXhq+JO5BixyBUn7bw2ygMBP2r8YbnGMIAsPnJw
UDrYUEAULKMwnmVFYRWW4pA3R8BJT3VNNI/6ui0k8y68L+ICEX9sNr1yUbsDkGQBxUe2dUWURr09
8zEQ+XkmWF79FFtWL3OF3HBL3eyLDZ6Qb4MYiRsyvS/OupjraPe792GWarEjj2kWTRM5twvA/FDy
rifmyMgFFQ24h/V5MF6aYOHRfKq/kc7CajSHrg5i4aoF1GbISWLmowzJAtzyqkzglE7QxV/w6F2K
zYZve6tcj73jCJGIbFx7g2XoWXH1nthlUFlJD9clQRbliHaSEsbBH7HANWr2ldJhUC/ZBCUMVoN8
gc7FfvZ2ZvVAbPNIHAFQJ5CP9ADnPf5F8kzGOoixDZKoaSgPwCK2zHWMLc0p8pYJ1Y83LPsEZOeG
sPRKUMonGXFXVb01BlvPSQ16DhDwRyRG+oBEnfOu6P/BfoXb4XmdSnmv7qa4BzHIws1tvACeZmkg
kBbeoq1cpEk+QIKYxbIL4ZIbdD3T1U9NxbOdz04FrUXFai5FZ1ZHJ7Ao+2y9uM+gsX6X4Dq17393
mhdW+e5srWyeC3sKTA0E+Smj8nE0vb/rq9F9KKiJYWAPrZvvXzSYvj/+lR/h4keqSK2JNzt6LgMg
HdLboK0r7VHs0Q15MjqLqtPFtm1iopBu8tZzMswvwFSYjo/5CmwDg2kpvacj7A8xmqwD/n+g7jrL
ZVdymufSg9Yw0xHDyigU9VjYGnvtMFIpJnndAP1R97VYa/DjcijGpbNCs9a/gJChC4ru5xeoi0ys
kRyE764vZ0geof+PKUsmdEAnxF3TO2j9zoRtWWhdsn0NdqFqzv8p4kQ8Ueq/9C3ItiD+C/ug3l76
YMWlUus7nMVr6NBnnVyZ7SHeGUGuJgeFW4iHo1XIR1oA6FYW1s8Cfv4yAw9r924x0U/eJm3c2MLd
Hh7z5GYyxYj1JTfZ9FGk1QYvE+EE9XwHYtpHRm+N1RyKKmXyLgWjfQJ33hhBeywjL+aX83j0rWH2
D+25D1WN8hUzlVxPGWlv6mhbie1WxyZuEY9LNQcjU7vHm5ooIcJbix+gixwNpkhc3bcVpIp+OGro
Lo2uU1T1o+A3WlirsLHHcA2AdA8bnqyTuwO10yadcLDxZY9PanRHsGkJ8BuFe82Ui/aFA+3pbMEO
EsQ1piHdQuF4db92L5YGNdDZvkjeDFcAAKprqklAKJk7TzswpMSUS5pR5HwstN5gHfIvjuHlNkP0
NjbbaNRNpkkq3Udy1aIN6zs/GNH+HbDM6Jq2FXNUqjJy3fIF7meRJkKWXJOza2XdH8iWuLWRpkfo
R1SXQ6Q0fM6WoUOrsQrv4UKNP1JvE5ki+HJiyOBEarzKeLQysuayPLZ/QzQg8ltQcejD+UghOKCg
kVyjhQDVBh9Y7PzvEo2BQB7FgEYWTF6WjFHtjBv2oujAYI1CN28MM5vHGDoZWRJAmm54jLfoTy2O
ntWiHhqgNcHjYAcs36kV+HihkinWRdqBYBsaKY0qICIYSMhNW2CzWR82L8UF1UTb/S0i0FTkCGcA
SMlV12DosNUwv8V2TQI3A2uHyhT/GjM7SEZNTbsyg2nPZrHZ2+vSrkWHxtfBdmBxxvprYq5E6rXU
/ja6QNTRQf+Z/V54mjIPZXjFEcCzY6rKU8z1dv2GSVY8ioRJznUBdkLZN+gxsiPDaGzkvvZh7XfJ
YCtaCm1fVhUfd+wOOcl1R4G0IFgEqUq4Q2lIu5s2vC1MGM005l1B4JPrgD82fhhiJPun1Aq35iQ1
1c46v1ftwu+oWEt4ADV9KIQOPRxsqjE4MaWJsFxVFRMA0iYJ/vmyuMDhYhT5RSWJwhUHvwbC/jiU
WBiF90GMZe7QSgA/ijbaVVXHH3h6IUt0ugnZkvkIKjGFpBYGh2tGo1va/W5BlPHf7SmN3tzAWdKq
CfbTFIhT8iPmDu3zGXFDG47YS/zkW757deORKr4AhkA6FFBWjGYrgCiUuE2Tl8EFFiBbUxPex2/T
GG/0VZc3ImUh1MWMmiQjQBnet3Y3TkQcDt+frCvgXHd17MRjMB/55AfuU/sBkeUpFJnyu8IrbLO1
ilG5jsDx3l+HgBU8+dXOQcC+krdtp0qnWGyCbPl+LWQkal6vuqe5MZp0zuTfXWcw0zdgiWoOqdfe
5lf1ps0UwTPvhJU6XZYA6BpQPA4nQlIjw4QlLdlOx6tMwIkDz58CqrgVsJEWEQFw/glctqkgXfU+
Zo3QpVSae+lOvZ1yfTOjfo9y+pcoTRw9LKHKZuIcK/svJfjLQdXsy/2NM4lSwe2wmrYnn+rUBZUg
PI/jghvuwKoESl1WlbDTRZebKMOvroTFo75mZAVVw6GPeiFBl38dv9Xq8JbxSxkT3UEzO55FhUUj
oOyeqzb6gNnte9Y9SJatxCelhZPxdW9VqIVMbsQsHO8zatZ6sp3T1G1ztY7Q/qIlYxW52Z5Vyml7
+dqQc5dJ+K8H82KIPcUTgTQYFvJph0CcvaOLa7P19+5QjOvcYRdfyiAMNvypx/96NhtpKXHy875n
e1ok/xgMbCUtoQ0ni9DczjJpbnYFVjPOHNrLojTsaTjWV5ntDAyptgIlprLiKPrjKcUefSiQo0oj
OqvC4hDQNbm4w0v55V2ZoSugfYA3PfgJtH1niO8uUoqT/npMtzHUvgM0M0VTscGm3q2dyVdxrmmf
5YSsPMMAJWyll0eAOPJ9QZX4eZpl91VCZAea4o5pQZIJTzDj+DXnK/QZDr16nAqGy/V7vfKGphj6
8CvBAisr/TbMDWQVEi308XELxiMtkwqBSgE1grDI2MUuH9gJtgnuA8bYVvUpt79fVzspM2eAQnzY
7t6ZdwWgl1Nbz+fGzFDTuh51ji38gQT7mld12QnHTEKGAmBV0o3VjcqWQBr4jGwsseaSpbqfD5pM
hGz55uAROtOepF1B+dkMhofFA2dsqWNbmNHb75tHsbGT48j8IYaHWTkGPzQMZQCExN91SPEzAKJh
c2+9ELO2EwosUoRbrXC7Oj5UUARcgRaAR+tX2df0QtGVCXhiKDAVGEYfpEWdnWjoZttvDony3AGj
ycj9ahKE+1wW7qrJE+C9OYCX/GI5ulCf/eWaQcFP7LBEgEkEfWatm7lvu9OC3SqT4ySSeWZ7bW5H
c5hbDxi74YlXsfqLQV4LdLBFEo52ZwfP8EVOSSjdyiPyqhXQvHoj7T+pksbeeb3y2vrG8c1HM6/t
LKpNcSwbTA1DFCAker8lR3YyZwe2mKsWMSnvdMTKe2G+Nuzk3Wh6Ghs/FMJeJEUHHpZHrxInYqPK
FoHpRxV3JRR8QTigo1vbnN/zvDfzBDrW3iAuo31nYnqAXdxcdfwj3hENUSzPDjSKfw/Hr6wMQTI0
B9e6Hjfv5cgMFo6L6w0dIHeiClQrTTqkrvZI5dggXfBqAP47HhZPQMBH+OhvCl/4jMaLibQTVu5N
mlINnYbuhmtMtWiJEfjQI7GnNSt1VpHkKUW3zojTMray07i5b8/D7RHzQCvKlgbnjD0nGznZOLeQ
K6pa6ONV2R5LmCCkny5sPyO5xPt7F605JJRJZnaHWHQmKHz7sOr1WD/QwQzlVnaOf85kl4/Zue5T
QAXg4wJOe0tb4cfajDSiFcwhQQ0uEYSC738Fn4ZvM8ILh+9kOSLfBZwbi9xnPhluBSGZ2Pdr9joK
j6zbvnAlRZ7eMrl2nTWIMPiwjndC6vD2fcpju5qBS3niLr3taI+vVlJmCeGgo1NQH+/CRexWqL1u
bm0vUyd3H3W/qpvT1wqczZhW1elafT5lGCVWHH4guPPVJkWsRlmW0S8Hr4M2SPt80X7Awiuyp3px
IHzxCZaNLo8OkocxZ4HRhWrIoIXkdmOrraAyvc7dFP0jxoCSI0+reT6DMg4pmo2tXRgH7eI81vz7
5esmihhSnIJyKl7BwCDaIoSro5qxHoWDr2aHOBjzPFei+Bpf7eHNazp5rZ5Nlaz6aZI3R7WrRQ8G
6VaClfJrBlm9MpJ3hfyl4f6XNWcxZonUzRfiS4+3kcJ5Avmg7MSUd3/4jsK3PKOcrn1EcOQqQnFn
MRgPWoSSff7CYXN6h8J3L3eFzYB/DpVfLNa45mGJDdgOD6xdFCnqzSXj/727ebyQ7UxP9A79AAkh
uxelgeS6gWgKHPFNgKLJBXolwXpzdmkZBeoFfOpe2+SS/0j0o68c3JGy6BcWk2eTbj6KAohhAVwb
qnArcXr5n0bWHIMXKinTGzAz5TLpLiGHgy+D7XP19j6A10Nkomtyr0ET/UAKbxdWzU4iuw9cntIp
pJtN5/g/JwW3BVyMO4s1VZsq+Xxvne7c25NeFxyTkGJrsfClto/vymCXSwSkfXzHhMgoaQ7y7Tcy
A+5w7YYorONyIVFuUP9SN4i9Enl2caFdN1L0cpVJLWPkCzgN49rxJdokOhPsIWt5tWPy8AQZUP8n
j8z+ZyUkhxZ+tL9UE9bbr9G8HsFih306hdWHFL+FFFGIwbhvJi4slopNhZtFgtah4aqzE5V+IuWW
XbJ3v/EqNhqaR71MLBsP9p411GQktw+Aus+yMaAcXMKs8eHAn4swnzU2aZmkUegY1U4V11jT7jG7
KvgJqwkCek6N3uRdhiqyt+1Yy7S/iCX12uTU4v/HV9AIAncXWFk4SKQIA87x4Ba+TVh/EEbL5xJV
dvT9X/559m8XZEvI5DQ8toXnuOmr2fY2+KUGMfAisXDnIn5U6dV0m/QzjDuM2Z3DK4qQI5uCakuf
o5Ydd+47kjr70EOm7ufs/DP2LiqAndD4vCcaM9k6AqCPlyTxY+NrpMOQRceY2xCAC+tsa/RVXgBX
0quEq3YWMQ3K8Vitgmq4XnzZ/WHSxwTS7Ykf8Gx1Y+9tMK/yOH1ze9XxM+aG62Bz8hUSc0LNJwUc
IMgtUDCUkQpKRsgI3BtXL+qHOak+rYWroyHC3fF/55wGZ8VvzaOhCDl9A5QrLOw90nZBDIEb6ZoN
AF+fnLtVRH3gGh9mD5hgtAdAby4+Lsy7jbsBYRfGnkI38rqtQJLYaY6B9pb0DkmaVe3jvluaCCQa
aajWBKIaAxUJtBEbO+w5vVyQrhalswdq2gegz66PSbPuh4XsjF1MbfByme32aAEqUMZHFK+9szsy
SmB/16KCLs80Bih8YMPnnVk+R+OPA69D916a53fGxvruavFhckwlKD9nztHAW2R/+xOFs9RiybUD
Z+J0QiyS1aoMYboG4UC6dWsKH3g1DP60vXGiXKtZjaGWysgxIime0C1SBxqvaNsH3Bnog7goX6s0
y+/Leel52h52IsfgzCDEMM3yFvRZBAkJGZhrrf77CUPVykeJ9em+NaQTbJTgGRAeB5tBkLHK9xAG
7+i8V3Q+9ERE1rFCoqrYJOEfmJBcDUH3U6jL4rRx6zkRaJR+SPNRcahyBh4gpsciEFtbmSpwLgyB
Eh33b+mpCeoONuPQlEsy8S9ODov5zlq+c20MPq/PBJh7wKBGjBxrESx9ALT0sVtSAaH+K/Z4Np6A
Yzb2FCDzwkoTBNo9kw3q8uJnY0k65f0jGXHapDZLa7d2le6HJoRda3DQRVmTQFQ9GSRqpWJtoEvo
bjcRZlZ/7rh5WwGUrOwvoJtTQsdSQ0PAklho3SpVWkr4GgvuJ2zFRq4vYZBSFCo4TXuB9N84fV3p
zr3rIfsLYy07+S9eifipIrrKopfGWu3JXJ4LWTT19UaGUKHzdvi7/ovAfzt5LRQixxte1peS/4j6
JMYiTEpyr9pAnWQjUQcULvInxGs4q2M2BO2oCkZi/OZsOfSOz0fWuGpWvumcDWSJl+7z/UGvaxue
whGIH2Ey6wSJZ965Xx46JYrDlR1uDzvhsk3x4XzmlzeE9bHVfVWkWs6o2XK5/HzOqthBg615Otlh
1cSUTZHMMIdCw1aUbfUlRZ7tD2qdJcKexc2hwv6Q2SJ6kwASIdMLEsk9hzRLlM3S5Sgtx+RZfDzZ
Srv64r/zeBmI5UrdxA5OvZ+pQ4/yB5jqeOQatcrA2mJjn/BRjr3smAtfYluE13elEwXFe3ERlguA
FbdpFwbILcy75hTVGBeVSpFRUFJDo7zbzGwZyNI0eWu7KY+D7QY5Wp+/IyQiXigjpel8sj+ws/YW
ho6h3WNgNanbxKWO8V43/AXsrkKMFBzooir1jm1ORDTqF6PrZfxs928kW6x3ExiaTJ/b8ZgDZhfi
BtKQTep3zs7tj9CTBFV1xUs2O7TOKEq43EnvcTQ8d2sPBKRU4UiKaEUhAcipeXW50IEdMUG10xxa
HYC8cEwc4Vyh49F+INFkfqF3kZT0dAPX6pqJhgM5LY661ullpW3u/WG1gMZQ66y70zRA5gMj50BV
fm8LP9GZI5zZSo3vk5UthsBeL3pU8SrVlb0Ei+AaMH9ZRMC1jHxZ+MTNwPctsPLcAtn1rP6fybdZ
RR4NqX+bXTaop6+3zbMP5rqWyIlo+w7zp36OKAHNzgouECRSVgDjD+HI6c6sTCNfIbGch7KfkZ4+
B/cXlegCprMJwpc7AJJmnCdlfq0o1Lstf0l1laWHphkuFwla8e8FGSWEzKCqyFBW+kDVvAvrKqMi
eEIDEwIVND5/Fawk4mdjiyqwoGGLCKJog3SUWHlC2MLpLyDQtcI+hdmjDVCjNt6J6DHxXp2H8S/B
mTEZ6wWBbec5uhu02/U4utFWx9vABtnXvQottdxKkVKCKMcj5ZhDmVJzaWjX8KPOhGkLS4yAlmHz
A0KbCnfEXkFj1crlB81Gr+Tj15L2tjr5+Mgpd/p+0ASqUwbm+60j/t/taTJfkd43bm1qvIc2p+i5
HGk2EzRdr0V7VTXLw2lN7xGi25kJp6Ezu8lD+K0m8YXcrJcl6gg8ng85aQFUiddqq5v0FCiuYots
EQ88+/WEdxDkH05xCqvQNpYZA6+kgQBSxvGKGAUlhYfXZ4we+txRxAnEcgpNdrhHbuDEInhZDTwc
cLNVneQU37ogXjVkOOrtJN6+JTC86FNUM6oOYD4cOEFVJ9M4HaHW9nBj7eQBMFG9fc+2l5Y5xr7V
Abn35aKmvWocqjJyEHM22C3/Sw1xXcERecpl7BL6zjanX6iENMTj25gBnfPdNnGDaW2toDhimBqp
XUtMaqQkM6ZdOCdVZ1JnYxldD+DdIntt8HswvDoo3yFhX2nX9hys5CiWUIcnLeAl45f5DHdhPQdK
xKLac9M3D1Uix63kmmqQS9/nuGSsk73gnyommNLM0xJYWSxZmOOME88X8qzBHMSmq/TIhq+xpge4
Aa9x8vYr1wK1F9qvKK9tv3RJs/pTm1hmt/OTJmyiC2jxVZ9qGJrBCydoE6u1/o4K1MacbgkSyLWB
vOkYFoxFIhAZz9j4pvIxv43fogJrs8WD358d2qIP0wM0nqUaAhUXFHSR53AhrDLK6PEF12ZJFZ66
+PU+X3VTf1Qn3NuYp4lNAwPK0/01E7KwDxq7yQHRq/HiYZ7Gu+eHvLMzp7VPg5WYcR8YKldAfXwk
eoFjRuYgIt/V9Iib3y64a5sqRlEV35/UAKHdRX/6BSbeonOauuoJ/hTVshd5i3e2EshYE0h+WE3R
e8Aw0pEB1Bs1f6wLJjoD6o5TlLg+rvsBS6i/QInRvOJcyJRtTaBs9w4jE1CU5FxVMM5sTy+/uoDN
nwHmbtxYQX7WXsnEX8+1hEWlQOw4iUPWErZzaHxlOchE4kS1jwEavYNqFGAXjonmI2mYi158rHn+
ds++ZejeuschkTnYGbSk11nW7htU+pjUrOezblu43p4lt393XYtWVvN4jmjfGGuZozZF4VSFg+2o
5Y0sJlyTaZqntvKb6Z6GAL/DGr3gU3fGTlSSLiqQji9rkiK9LGReqhghkbYMRSd1e43zGm2/BWSd
h67Mv3zeH+6GgksP1ul0bbjwSDQxUGXk1IchBH4v3QOmrqOsnJrQQMn1EIip7NrRyOyrx/0k4fUc
I1q7ECKU6PDg2Va7MzmEWjHGqf/c976XG+QIWX3sK6gDBx62BsDuX1IEltZvcWzcpO7sPOojTlZA
LbZkssGGRsV4sVCBtYiYJMJ6EcYdQqe/SZipgZuEBs9Hi2XctaQYp4vJ0zWebBazNMeYExyn8WFC
rhqRNq4oZeltoWZiYRfLkSHpBclJ+sJpysPFgr9wB4uRIY6l+VLKTm+LGVkSuSd5LhDet9Nb6kU3
IPCpMsMAsFC3J9bRuZhPDKE9HX0h8K/Sj9oWSLWtruznWQlYjvMu9Dy9pqVxvZ/sCdJDP7tsIX8X
cIU1zBweDWe+2DTp3N1xhfQ/Sug67EaQeltoHJQ8KcorBRiUP+3capFBi8oSEsky/be2zA7aphN4
VozIyBimjElY4bSTO/2qFxuCcv3hemT4MBybcSiIAU5US8ufDbhu6xCQyzIVzzQcUrV4TyS35TBu
a6w5UqJmWG6Qw3TTvvdBkawvVSimGQZzX9lU7OYepcnYRsSCGdUsiP6oN8mG5tYoJgKnKpoZ7C7+
jXgt/l/MA5Jgvp3HR0GUvPM+ymv7E2vAxo9Qef4spxv0W9BgNv4ouFMGqT+YcVrTQEh/zm4oLIOw
N+nl/IRCECh2W4yfO/h6ktTntHyOHxkxNdcwg5sVGGQv9h8E34WMD+nH8V9dlegCh/2ER0rnW/Nv
litb9ixWpqV7yV7Bsy75PokoXp8qq8WQ+Q7GVmbJQp2zQXc1qctM2+iaVqXmvzPMy3JCG10GX3q3
4/DMfCDkq+WmaDxw8nKUVWs5/QLQvqF3kQK8BzpNFVLxtHf59VAPpXQWYmY0/d7L/crZQUyoTBVI
kOl4ZRPGIheG5FUQdItVAQ882DbB/BFXy920R5J/ZBiM/n7S8s5PuJojFLJk0s8JnlOrxbvh/3Ph
Gjqc03tFGUkw3vBPMSoVUF1xXfgipnpFv7LpHEZpBPL3wN63ssBbUEEvUnXeAWYPkAaQY7kYUitU
35IyCZajD8Tgn/E4eG3x8k2nFRNTasYyiRH74qXByu3zgZNmCvylssx1pLFMSTLOOV3phc7MTOIo
OgGp9eub0uU+vdezZVDKzd8O5ED2NhuuSmELLiRh8E7cnQseWSVVfIRvk/+OsCZv/JqMzloVX0Ip
i9OrW+fuFuMtBc91JlHmo1W3GN6vCbS5niGK3+RRVe2GkithMywT6KD+M9ibSwuyKaMwHN5JpdjX
BxBX47Ti0/oyJ9juK03ags9M74XKI7NmzY9b0lOb7lp4q91r4BLdOO+vyWpfCy9/uG9ABkslYAgP
+MwBZvqZq8UfnfD2qCWIfbZMcFeQpdthsW/lw9VA/aNJti4aVfKiQqdBQpOUwoAmJcvoZmRC9GDO
lgC1N5tm/CI0db9bUuKz/AJHLzcAYA63xIq2rSluMomFCvWXLbW9g5lRuEkKqeekmmtda5qZqmRH
4aM81fL+kD1kkCZuFd4IRLAlgWr9kySBrQUChRZNmPp4oSs1/C+GmPOnMihJG9Z5y5s2L/hNJPrA
JHCaOccp92KOBMeakRvDRObwi2i7tdhFPrGokdKUTyTOLkxr00fH7ctkAYv4xG+AJbgmYVerpbRo
KcM34sU3ubVafXDRYrhzkmvri9npxVDo5iIywXd8a/utA/jE+MGResSiFjiTx7pbl8rv4PKpmNe0
5fkDPE8m4tcgSP8NwZXrTsCff0T3HI/B7/hpYtIo+zVP2csuXxlYXGWBx/J7aiuJkhSvOArAnmDU
GBlQLcefvML0Yvq7kRJcSdyYMYyUP+okMjvbcb04CtG5h/XNG0tYNR7roekaWqHYaBqExhgx6+BC
NGhVIahSNbJqgjN4H0S9yxz10X7iHfMuLiG7O63dBmQbNhHleoo7BJY1w6Rve/7SxmDE1X+PgI94
7EEZVpfJA4/3Rsq95MCepHB1MrV9ZBE9LzNKOBEJu7ltF/1SYT3RambGRSSnLvpo/h56V/qSDkvL
VUSG2BfKB10SPf2/HceW5Qr/Lzn6XDlI4xXp308mANAh3/29ij/+xGyRjea5Lg3Yshuq8N47HBj7
4unotzE0jyQBLaNTOQ9kGo9U7xHxmjyz6c7ygQYgVkrIR4GhN5uLobpyjDsNH6Eqc0LsYJuk+nj0
4W8HriL1aslLv5Xd8QtP1CS3ry3J/GR44f28zarjS6HNBrbSXGO8B+vx8YE6+CuoxRs4EMGs0vdR
O57tY3odGxIu/lYAdyogLwf5vAh/nErYmICd8PTIUveu7nlSxNWRVU0TOUvB8I9ZWbkg9NtBgGs9
iiOZUnD8bbQSy5LSzTJ3XUQp2UQEvGT3mnE5ZZ7AFkJ2GGfQqJ1qJcd7pKmJZbaZPXqYlXIwMBwe
G9x6gT2a7ZiLCloizYI7V8C3hG/xeShUN1Gu7ZlYPCmUymVcuLzr7TSjb6IpP0YnGZlEsw3j5kCu
OzyXKiPzAwkXRbN9EUnSFPjlea9LzUtT3bZdw44nRPYrPGzvC1z98Ksn7aemEVjEFTXHq1jF48rz
eO/DmVCIuuLf2AgDRSvOT1WEhk3xSQADCCBYV/+yJL4ReUZzkCmurFkXkSHWSIMLBm8tIZxxXLf6
wzceYRb2c5xd9k9wQdybyWh1Q44/TuvcDFcWR803Smnv7ti9HO+oP5X97+i4zuyKTf+YKhU76JkX
y4M73bKmpmGhnKKy6AZRVIJRwKf6cGq79A1gIZlKZMjtc+GYyowszXyCN+Fj4HjlzcuuvfgnrLT1
1mbVS84qfd1wZ95xdVENBBSteBdl+K7Q+XAPkXxrgpsAo+kWo6vleIKFNZXitz/VLXyF57S+9AGz
ErCEQPMHqwuWTeip/3oEiWG2KLJ8La0ynukrsewxxHu7sPD/0TFiQTGWaHuBWvFcz7nMrufW8UUo
vG3w+Y6AqPrwAWqSYDCO8FxKSCb3s6GZ2CEli/gA/sMP8mmH8K87Qv1oCPzfRGEKYyQRV23sTglE
zrD3OPDrlBalCLPZ4LGToLByFZ60jbbnayxJGf5tAtnVx3T0xz7gwaY0PwA9E6SZ9JUlY7siO8hR
E6s8fHJUg++y0EBZJ0hcS7X+HlYD57VjRTpgf4pJOiQ4tS3WoadkpotR30eXdDTkRbVKH+7m4CXO
SDDZbm9mDrPXRLVt7eS1RLFr3Z43jK8Jh5skxlvZ58SlRVAvAFjScRd3TaCu+aSEH7GK6KWcu/lu
J4w7GZ/B5J2WNzcxMhFu4yEqaJWLqmFXSytsRRkoFWlUDY/02ZZthMn7LhMHQwcmdlcCeIXxMyfY
/L//WvBNyPkb6EGU4JAoxlWKGqrmGjfUs6ohln/u2VktvVJzfnrcVzUUTBwaeSdlZTlEm8Zp22vA
xfBbNL5YNM/XWdHYZfodC+Mg1jPuNK5TjefTnEAtmLxpr5MzKT/UokY8WT7rtEwsjV8gvw7zlags
lopy01/un5Z10fqAnyaJG4aQ3JiWXWS5ZrTkSJbiy9x9KWLvGxuj8UEDNBuWURg0n7jEFxeRIVUe
8V/3nFZHS+ubnjwxwDhnBsxhm2PveR0n+aSgHbwqKnfVey/Mis44wnYipSey2eawBZALdliQu4Ve
l6NqEL4EJ47kR34tdheofRm0YEtuVDzunzIzbo9EgxK1q2s9W9v2uub5ncOtW1zc3UfFQJaOizbl
00gSxqcqyL9YF2Yb6F9CVJ5OTNar6Frq9lTe3S/QPOiZ9X0oD0iaN9hfLWhuRL76oXM9CfV43CE/
m5vY015D3ljZxePxpHe1wlXWoY+XqcpUCpEuf0TS4wx612BkxJmeMAmmMSTlyZpR64BZ0L2Rtrmt
GfEW3yymPrYoVwf4R5VXzSZOtOVAShruXtmzZvZnrjiueUcNQ8pACURAD+tiV1CWa/y4Sc8m+ZVJ
OMCaoM33gYFFm0EW6cSdTdpu/DZud26WjPBuYDMUJEigvXDH5Q6e6AwNKKT2LxvDHOOCJCBWlyq1
pDCiORS+M3i85ltfW5AJoWY1BCXBwE4ZBMMfGLpE/9JPFdqB07UDP44TrGIal7mk+vLEokvFFA7G
TOzJeWS2h8s9JIs+7OWuZpp3vFj28rkXSzIRUM+e3Kq6Y4H7T152HquDN81nRzQg9rIXQI0WRIWg
B4acM7RG/xzUxed6aCxzdeLbXNEyalZWXCg3tl1UJWsS2u2v1sw5tE0pRmUYj9xxaKS/0Q1hLMlF
woPaUrKpS1Fmb0bQCJNOpo3Hvju3+lp0++uPibgrGIiAFbhFhK4NYiffwGa0sI2Imx3zuQwnI8Kg
xL40mIhVvcvhbUFRc53WI5q8+IXgeCbNwwVlllq8sQddOuKASRg06xMricpBrS/Oyv4q/KfFLkxM
ur67Dd+K4gjL9958K/zAOYgf7R5ZVcTOZB07sQhbt7c15jEMxoQDY4rNo4sQ73jm4LBudTbO7mPM
5YL/ZSXrFwhX5/aQHmBNAPckn2gREfF+ChXXFDptVW5noHhXTMue5rUIsuc+L1aS107nIfLRYLd+
FYf0zTZ5k82ksAJUulaCl6PflNUHJtRbOMEF/6BEzZK4RTA9LN4WnBDzyxbZ8tDP9itBqJyhUcE1
/C71Wscz+jk8sTh1t6bYJId3Kfi8paOEjnOJnnX7mtoRj9s8yTvjgKbXbWtpueeo5/iq4d9zOO2Y
E+e34oRmtc9p760isGKMzRrCYdS/Ctn/v/cfn0LuupIYy5fM2mm+9Y6ZF0ttpu2t7oCu24Wbf+20
o5zuSNSHBhLx+yS3mIhK2rRP0AL8W/TUEaAiMUGs6MVhFq2J730wfgcZ3UZMv+4nxLAYvDvKfP0E
pdWsLQcjcneFG24qJNUbwubutVFpLDXCymqdlB+u4cE49/1KoMoA3NSKvL1f3K9FfGpZtJ6Ctv9N
Idnq5yVVoA5NEedeI4avhIt4ryUE6UIUqSihaLLWQXRu0mHvtj1ptOyWmVY8rMx4U7M//dy3YpjC
E2auY8OEgjweW1C2ninko9U4EyGr+xlxLxUv3eoXBhnC14AsokNxYwuZTDXX63YwYArAnuaKCvTK
Gx6/YGwpDAdZclQdXdp8iHbf4qSB+9TX6jWyYKXcxZWz3C/dZmKpy2Ax5fbPdSZlnvKAI7m6fECd
z7CPCuQuPhMvsP7WBtBHe3crSoToMRtjocZIl2CjX6m4U0doBYqxLVgpFzeNwHS14gPpRu49TgIc
5RSo0jSS+os7zA8IebTLiSNq5eC3ac2nQKseLInkFXuto0T7sNz1YVZpCSdlwWBKaLdUteFQrbb+
jcy7v8EqF70YEEtkPPJCVVdknQ9rFkyNrT42xlkNGELLdLL1ynflO16vKm05oyw9GDh1aj7Tgv1/
F/eloruOyju1EfpAxKZKfMHJ4rizynXGqdAHLy8NVxrcjaitCOG8s8O7KhEm+bA5nw1jXApPgRIg
SLk+zI78VWVybFo9jut/K9XcRl+KVwJ8L7oQ2i4ohCXxPqTDYXRWI13DbVwYHBPkwMgk9os7cxf2
8pvn3jqHknrVXS/4WwNKCJLv+QJo5U0qI8pDnDCdqSifAmPTGCSaOxkSCqz0IItvRGwRTUUpcs9e
FSeKNy/0I6KptCp2T2vOf+CI3HDu/08sJynpqh9Ttj79z+xlJDvPpvPsFnWRm7T8JQKl5VYFS2kL
GW8FJsB3AfcR+15PmdPJqO5q/+mTgkge5CKL8pejST0mBRYkniIJrrMaQcL+Nlz5Jsx/cmLDEERo
JXkD+mgzZNwjd7nLUk0pyXLVh9Vjb21jLO1mwTFt9uCBcpvL18Rd8j3BGU6hxRrx73eM3p999UdE
8Vr6ZuLHUPMidohg63iDR+a17/k7dP/xnFOG/6CRbqgWUj5VK5NuSWXdicWenJcvufAunyT8r0ov
D6x9SM8MggbEHNOaU5O/wEL2sSjE+Hd9TV73N6Gt8LKhsOvfiCMbtT7PFI6ceUTRFnYpyJak54ZP
2MwIfzR7g5kAnW2JvVvhgn25FFcmiIrmRL2kH6QTZT9Yz+EM9yErcAeuZYsGhPrz3l5WfY1T03aK
+7AFR+hjobUIlhHk2Y7cEE7bmX2k+welvxdnnxxjrg8vz3nbN1Xo9L2F9fSKDnyrEo5D4frG1crz
eYREdN2X70kASKYw6f0HRVjQAtojyA6X2eB/wd8wjPfmIIVFsUTs9eoAMstZztu8XMO4EEgktOz5
rVIp2CyNEHeY+8zYTpgUm7DH4eFKyIAx4INhOY3L8Ox2bWmfNUfCfdumvdbgi5TpZs4H3RmONwQC
OCTE+fO5leHk3IwCiYyvqjyuSx0mExOA5lOs5+j3FOmpGiY8DCWNNfH/N8Qmu+9M+wFxczOnlGHj
JyYytdxk+er44y0AgtS84l7/YXNd3Nkwgrt1wM6zbj3ugqLYlD530ISJd/QnP33ydIUSHK+i1iaW
dBN8N3nbYlkWhHd+ilk3xNlNXKdvHHhfQuWJpmCP9GiII6t6hdEzOhNbb4PIp6+nk1No5e34Inp8
GYBwdZJGdZqrxFGyDsol+6ZVDBuncPCQBsPvl7nTUHvbEY4csLntceq7IODz2gFDn+SH7F5gKIZB
qG+WFYdlOXHNctM7ZjdiAutfLqWbeuY4oqUx+eCgERrAGtKXNgdd+qazoEAk9s1UpzrrxZKfJSTk
U/gfiOxe7X75gYd99oO6Z7yseUrTjUXhLPF6OEh8kz5+4fA+pox9xWXDARXFvvq/8ZY0eH36ov53
Q3tcFfoVaXicaclrhdKJBMH4TJgUHONXNBFvdZTRkaTn++Led2qil3g8h2LH6nB/kxWRw9eqtWQ4
96lMkjbtdc7GKBhBnZuXPrNT8CLLoJygXZMb7y05CBpFupX0965nEXTMiAGMy6ZyAp6CJVDpj/3M
xNyOk9/vKJdP+QYWJ/ZwbtMvOqlo4qUoLHINswv/cmkZlaWEI4CFLFkaaqA6jW/jqqs74YbaBlLj
SoVV8QCoffCyfvMZuUKu4g0xOVEkz71wa083irnvjR+kNSDrBHKZfwftbUckKkZzEunsyMOCfAop
jOBSo6GJfptM5Y8LMqyqpdHJyZnVIhhFLcxfixKe+zwzM2/caf+voohnKxqqmuows+56UwQK5KVW
EDcDwHOqj4sbP4zrFfh5iMbZON2WseA4xZ24BOkjkwqSC0WiEswWwGPc/PYRLlpFBU0g3gqfPPds
W95SME+Gsh/cfO4KGytrDwh8illvB+CTW9xysnCd1DpGQA7mzVP8DBAr6JXuD+AIIzQ+QOs/lURM
XELpw/0lGdPmdKCbeYZLMiJlEy8dd+AMOcHHf14BjarClYq5L8JYeNl+OVwBrye+wsSMTNB0l19r
UQzPzJhq4upKCqBplp0RC/cYBGd44HtIoRU6p+P5PKJR+YpyuzGULASyfWASyQTVg7ynxkYGUOCI
ZUuEiF2MilqHoqH2Xlem0WyVUVc0U1hZkA8KNkAJ3ZIC+ErIVPfsVw7hnCM1yJXOunewdfjLnhjJ
/a296L8tYQtoHOrylMj0c+L7ZnT5CymuSwgmnPqjYvCjJKdHJ6THrPSDTeeUgFpiX0OZOOHxGy3W
+mdx5T5iHMehmc6DfFQ7xjtuzn6N3EUJu+8teNIFfwS7B4M4IFycFbh6hAX9XD7Z+jPk2z63D3f4
xZ40bdWqnI70f27mEf3e9vcdMzIeZ/BMSLXSCgDB//ZHt0Yzw0XF0DjPT4ze91v1/aXXFe36wHjz
8p1XH7SmcSOmq+jNhJlSkHnA8zVuAHPPY7OM2Yil89g1NaoLTKYUb/if8eABQyvXgOTbfjkQGbOm
T+5uMgiDbFsIek3o0KTYqwfI9rrdGND7c9YJ1MM2cScUU3zID/bQCekfyv4C4+snTPEhrRLXg1CV
DXfpKLznnv294S7/i8hTeTUoQJmBwOMlKxeyEQ78wDEQGfsO38mFgCBdP+xNFmsDU2PEFSbV91fb
mrXUmHk5pcVzE59Ddc6a36BGytWXO9q7ycpQjeJUgAk8Ac3/Smbz6oGHsE1APuPqp+nfoShLVInm
JOBb9iquvEfE4f5TYhpNfzXmjhOk0Z+P4G2ugOEWJRk/i5ceZiT7kTeoOqg1T/dSO0/5HSQhWiZa
QGjzo7J39VoSSPRfLYj4wSWpWnInFuVHLxHTXqeK/SeeUw9Md6hXmskOMxTQUAECcs2tXGEVCBew
0u1himS+dn1eF6MuUaKLpl4iryxI8G7wDvxikVwnkXU1hyJl/nvi3JyS1FQOlasFXM+6wRjFO/5t
/DN53x4ZrQjWQnp+ezgUxkEjbbkgZiqbudTyNW5O+NXuK1/bJQTVv9/0ctwWYGSFZVg6MHrbdmwK
WAk6Rl0uI5XnJ3rkGzWeYXMqVkeA9sLv9CmQ1t+1aUG5ip38yw5wG4duvtPJdlltgL3BRvkEaXTP
hTXHnrN+YmlPA1FWB7YNbT9yZeMnyEnVFQDOUz8sXBzsu/K5jHj/h/JAbvTU1E44+a0oPm0cTMI2
g85p3hDf2wNIxiQLeytBGhy4qyTPXFtO2eF7ocpas90UpzVeVD7JSNtudeFDsLw/nPQCbyt5rKJE
YRumSTDPXqbO9RDDFJt/vGbnvwmOQzOfs55Qr84SQyObF07Z227GRz/eO0k7iAG2UOZKCGlZXSbt
XBQ/258TzMEl3pyb6o2U4kak8XKiMolwClXTLsw+Alw5gHmH+vt62DAoyC0jeU3deXXiYLowb/xr
rBaOl19GMU9T7QiTR6ptUz9qGN/RMVeje+29VMOlGA4cQNiHmglcohk+P+/wbb/azQ9OJDUnkbJ/
rSh2NNFWExKLNQS1nrmXO7MFVZytmaKWc11CDWI1t1gbPluVQiV6GHmxtWAguNIwrn9YU4AbE/K8
xcX6LKYWxfuLzssPGqy2JZUrjSD3CQ2tNPpaLpFzgnkF5dkRUMSI88JNJwPX/Kd+XFpOUteNslll
8AuFZ933SyBdZa1++w4i1g2uUUTDTuOS4aCTVOUpfuMCP6uBP2mlB3hNaC1Yo2fi2K/KmSDbZaoU
BVjKLBT6/FTms0AHqqYwTBC1ngLvfEmX0QcE96CwRQdZ3YNuhf/QMzo3kx2LnIOANLiD0ddalVBB
WySQLuDH8tfB+MylcnW6rAqlJpo53bvEpDAimm1BG9kL2JeAIMkk+qMmTvb5/wgAMplODUdMck9D
xjYGyWUrlhpYsKylodrEwkqrFEV97TSbd2jaDkt4TWS2PL7+5NLZFUT5oDsetFqwfhuJmAtnHqJ3
YngJMnccJapmX4N2TtE9WrDHJsVUNgTsBwQFwDMrt2IVU0d4DdF79Ak1bLsHTvCdWec2UCvcyIBk
nk1b0H6eRsicxyVZWRYqCTNiXzYDluLaOBiA0pJZgdMUpHAAJped52auZAqrwLkxeYegsCyOGABU
5k/pUZ/pXHU1G8luCxoqkG41xbX1kYoHOvYMg5uV6/j8Vow90wgHXVjo9A+VpAOSTbGeS42kwx71
qM0xQsn2SzWrzySmZZb1d02Y3YC2VkuElWnZcjoTagfo7dMdVJiA/Z9Fs3bznMvH5jupsSwK2Iq2
7qntjlKcV8XTSv72LM1hQVoFgvd/BTUOVZcOEpaoBhLhCIKJrZeibJrBuL5KB1xfDQpPPQ0ggk8e
dcuNJoQpXvI2UXszyz0ABB7yPgZWX6KuxpIj0zmBkxITIAO+0zbnqk8zzlp/ZUBTbewmwb5mpAvr
jGNG/msGZ6+TIpoeViZjdF9yve3w63VMKyzYdzEfjwfcBuKuQ3JkyrC6VehlnDabBXK+WRJX5UOc
yydiZxGB1qC0BMQkjwnanP15SjrZRV49Aiu50pti3mAt78/AY54DkATljT2Cath0D9qGr4XY/SCj
ZpVNcBhTAVkIht82pbTvxEtm9l5tMYdnsL/k2gb/TrprQRH+0mrFWtdgtg8geS1dMB0ykesQJy55
5U3TqcYcQHucjUbUPahlsk0gN4IFpRbVVJlrDKokXbDP+kpoN/60Uk2FxZJJen2UWqTpGyxDvkMa
pt6bT/HLonFGugzzFSughQclYiQOZYg5otNA65+h5jVsnaX+NU5R5M2n/rmrs5HZQtMrJk/SChlb
fvFH3BTeo2g33bpNMfhr2TSQWkC1u4a6R5z1TWj/wqfg8lDz80BiNyIGkniW4FgiyJ9dEF8l3mIC
JoJhnwK7sjOV+CLNvk8NlaEtq7t4xomlnAvdmNkQpC4Z+3l7skQvl7uotPvkLVADaLqrhpwlAGPw
Us3fPSL3pFu92XKjddns1n8TakTYOJi8rbKO+PIcIYtDB37igJrnEcExgK+/WFfopemLt/XDe97g
Vyzjvbj8SZmfeW69iR757O4OxWKENgFI3nHSLWqI7E0BFybj9n9u51mI0TBXS4nM0Egk+X3jtT+a
Ro7g4vhEcyDRbQ0A6MymtzeZWMGHusjatYFOBnTbLOobcUJsW0QpsLEUtd246Phow+VYm2GxnSJ6
aWqDlGfkhecfHdYZMJKtICDNsEJaZO4/JBFZmekuhwSQ7s7M0BzvqG/BYrVp2uFSz4OUwAC9/BU0
8y7sJrTStei2TMVDIm8SwYuSH8o7q76uf7x3Uw6a9aPTwpG9xoSkSAPMvKyHSdKwTTXGC5H8BTiJ
q0FUSXDTqLvgQv6Q5agcVIWSgjKrAE5uznZLBxDfX6YKtmhFWYujmbcBU0IloHVxewrVXfiRj39+
+7k8tOV7ZBJPM51QzvF0WRZnmOsroMA2yvrMcypmABfS4w2Nt4lNs6jUIbzlhfwKWyi5w5NKupeX
M8ZgNBNO/RlNvof3QOskJ6/bPpYHzO0hM8AWNQog9G3vsZxXkEvJGzQNlVBm3u3FDVPXbTt+R4eq
CYUMx1iFLN2+oDUDi+5+Sr+RBk48Evxof1Thzt1KLSmJjzmwHgCwT4nnACvORG+XZFzJHjQCnuaV
ByBH4hT2aRgMiidk9spC2o8B5wF1nJLh/u6FDpG44OR9VSmIBjLuWooLJu4S+bcePaNpMTknZHen
zeNLfUpsfdlCbqldPURYm+/zqM0v76hH75+cnRYwWfVZ/LyJ7BX1RKs/aIw57RfMMFompP9tU4uI
pG1QrrmIKluMoLc/Py4xjzkdxhr+LJ5zrXleDOKIX0U2J9FDMgsZr5Xx8zwYV/JV8tXWobgnRxQE
ptNrDhtzKda5hAbwqrjp8Pn3ZDHU6p/KbqLKpVUamLdqgPF5RIoarqyCra0xh+Ru6Cjr5LJhacvz
UTi4mOykOuMUvcZZsEqaR1g4CGx4dRBdQYXEJHBMCON1rHhId/IxgJJy7tXYPVJcnpGCzywMy02E
iYwnz296mpSCMdNeUPxsPa+a4bMw5OU0+olTQuOQotXVtRIkRgGKwJMqYWYx7bSzbYW6H4yBij0G
wypmQtsei2KOolUBPzsrEtTwEBH0SNLDsqSFHh1B2vxT0BAOCijeiQjo28AbOjlrsP5OP0Wzly5D
9OwjJo5w6Ab3uABJWlo7lvfjIAoOvasmTPujZmNFQTpLHtGeMESZXPCSjntbiv7fPweCieGmrHWR
H/r5zp82cTRlbioR3bEiwSOzS9wJSoy9e2a+cUpkQnJGcv3/0+Hfdwel5TAWY1ceSwu0fZDK7HnI
nqYs2hjzzzZXc5vJlG7Gg5NR3HT2Ci1B6l35iG3wTsQWXrOw7QEcG8GeL+HtAf8+YW/eZPqbcxg1
ipYgnwG9YVa0USd2C/WFN49lkyitBbLR25HldpgnEKwbSjRYgglFzZVPWrW6ijgqyY73Cl1ENbsY
ZPCTVJowtXZZZEDY8Q7qkyB6aEUBKCuEqtFvXdzRYshMAiL7luDeXUXR7u4ca4rAbHnoAwTl84PJ
eqaxJOyRogR0V0XNbRG240iu3JSlgq8deYkonYY+s37V/q8Jiea3nZLSOMDMotYkqCXSn/OK//PB
54OOToFI4G3uOc9WMoH6Go/Mz/cw22bS9fADzuAyqO4yTpLkw1I33x6k/fATE5Mn14WpPLObpo4h
ANkQrnSXeHFLlBTuxoXsXicJGo7MjJ85VxeAITXjMA+/Jd3+1T6jplnaTjcodOaI61qZ2DYr9WRZ
VfnDIjfIP9xf5fq7Q4Am6+fPTxZyM6bWrNKePDw3q6934ECx9DoMrczmyklexClv0UBk9sF2wANB
c4Oa0/afukif8YIrSn3Vhhu8kFo4CqFaFU5wQHMNtFAsqyfeTUT+dLVAzNtOAhbvcqv3aOWhzcdh
fMvyilqpiwHPiKhkg8RknGDjMsH/MsDcFaqyW9Vt2L0mL0lsCNHooEvXK3KQomSQ0n7bzBmJ4ihB
+DhT4alfFPfAtM+1bqKdzUeUo160PHDaxCNFMgygNPGw2I37g/yflUTclrgnJu6o76ae65pECfNW
awefv0f5aShW4bKBtbVfKzLkCOE6SFVVy8L0+5nf0wpuYSJ5sAMuLupZvQ12NdsS7es/dRg6Lr4E
3wLGrB66Z261CUiJVJ3lJ4jijLz9XrqYPO6NKKmjBmM9OzXYE52xWZB9IEpLa2FjrGgwNS9K/1k8
egprn9U5NrAle4ANMhMAp1i9/SiFCCEuk2rh0bLt2j1pno3qF3Ss8/ATbTKazQe1eFxCXUJPtvck
FZeYNgy8koKh40fo07P80CPu2jKnwVXRBtV1ygXt80yOWso3wXFlftP871ysWlvkkHbCBLwFPVIq
OZ5Ntxn6SeRpa7xQ2KyOHlXoKWkYAGxcwSCtYNxEe/5E+ffWvxDTUS0Z0RZAdIZUZiRUukoNhH0X
j8dpN+w/Zs2u70QkjZBPmu13J/jYfFI55BL/RDeiQNH2v10HKhvy5Sp0ygggZS7Vusn5EJ4iRAS3
4joPGT64f7+vE37C9zkbVFxdqyu9ltvgTI1PFFZ1c2CEaPxTPhJENpZ/18sQFtMD4ydKmDR6WOQ9
hGGsgf1vqwJO4cFb5aO/m/uSdFR+3YKMxWdrGOxpEfLui0bU0/YPqBwhr82TCUh7SilHsqY4amTX
CLyYSLLXxP6l84fWC6UXATp+jr4HOJ4s86jCxgyLgR/eSc/C84ckZUkhhMt4jdfvYllHqWFOD4XP
7siupHN4YlSm6dHuaMGfBWE/uvRevHnS9tgbg9cmPyvtqtPmxmf8V1CzBv/76iFVjlfo6tqNZxC/
nLHEPyjuakxG5WICUxA/e/3R4Fjn7bk7aJmidaH0gJpU0GTeGwQwo7vmOJ8TM0pBqnDaDSR4j6K+
3Ar7eBH2lIQ+FQs1sVsC4N9agkpBKXFNxOzloWMyRi3Qjp1LEBLaIfZ6nF+KE1D3sAmtzjyi6S4E
UyN8rdPfPVZkTbR1RyRvwJNAPznmXFHDlHNGh2sp6xuhbkjMkwtd4lr23TQuJ8087nwe2pyYx5b5
Yy1er4OPmCy94zTnX1Ph0LJLS+C2MhHbpPELjTo9ZiFnNrYLaRlNWeLPLRV9Cg5XpJclgWbl/D0I
b+s+5kTbyRggpxzgIkLJKmKIMAys6Q7pKANp8nP36HQqLMJfJkMllH9KWbXWvRVmNTF03Jh/8OCi
XXyG/EflHF3JLSVEBnsPhk9uUywUfPvPjzB8msWZa2iSG3/p2u//FYzh5Z2zVCR3ixJoE1W3do8H
fGkVZOO7AwQN9yCmG9tZLYJgML4nZgv5DEEVR9n4qe1EAiJUr7bF1XgeP0KJptlPZQdpIstnZv5m
E7D/SqxV3NCT7Zbq5aSATZlRChu7kTptSJZ03geh0CnG4pYQgjIxkJckJU+rguKtQ9j4QiiL7oRN
8uBhqhHvp2KneRjgQERDMes5jp96nbu5QeEU/VkzBSVuF7dpO6scV4u3FDJJqchyUzkTJZeW1sY8
2FUpj9INAoA6AFww5W6+ylrpP5uuXV66eEa6qhXVgfNm8N2klnLVj4xThFPWHVaE26+rnTDrc2ho
WT+2DrU0+jyjm7z9KJvTcMVqXuMxMNowDiWDl++4EygDSyWv/yeNmvhfSSZZAKtLCEFb7grSNN6U
lT01R4KYAojOnH6OQMxb5hX0sKpy6wWgkrE22Z5FKgEtY/ookk1HLc50faUop42S+zSLMHg+BypN
Zz7SuIwKRb8riAmFnFamduuZJV5yFSy6GpXFW4H1ROOClfjDSevMh9H+TuHn3RclRzowfBn8P09n
wjHHnlXbu9kq71JAIoehu9uI0YqkKO2NodfNGUbgJyyz/CoRO/cbKQZNwdtmdknKWNZzPFavRr0y
fZ2KCBb3Mm6PSg+fsi12SH30vtahZ6b5BUdNvJe5GWeKZctyLMBAb2ADNH3OMyPi1h/MF/mmnMCz
7KqopZ8K+9+VyKtVq6ANGTuMyVhXW66wlkwM1QbivXEexP4fjruNxn93Ev0KkafCh9CbYiZYCixo
qp3/vSvxeNBLCOjQ7vrIDEQSitguOUVUuZQuQmmJeNK+KS+MnZ/nO5UPS+Hss2st0F/IYR+BIpDJ
+a7of6vSweRphjV9edSS+0HbLxj50xoovMh/SdS3K7WEOfz7GIMWVFC91gDzXMwrr63QfNA7Raee
JN8FiOI+WCRVtF4Hc35tTGb/OZsapXHUB9WABERVDxA2+wfAqxZhckoUtbcfbpVtrgAAjrTH2VDG
wmJ577tTtniiBGc0u75f0KlebR65zXza7YW7HJZwH5WQE/jSVZkxtLsHHASL0C9RJOqljtfDyg8g
5LkVNeFE+LZFVAIXPH4hgXL+Bz3QCxrNmQVOKy4fzlM0SoPao5JsMv/i2FSfxr8zvyskEoUknjK7
jXEPzBu3J6GxH6BkZCcxjAXhp79AaGozOROQupfkmwV4suGG+yo8Vium2p5hLsHIbDghB8eC2GY5
aceKOWczyPgtrXwS61j43LbzuZsJ17/poQLHFBC+YAuUJ5usxCAfQ64IE9NBcej5lUvCt5zNblsG
CesQT2Kj8Umkdmrl6vxeS9Z2WuJYdrt+JHMb2lWWp6xuOIp9WCNIvDPz8qPcWd6aV73iB3GY7r+I
YphQD6K6glHSz5NqgvBPT4MKnChCfX0bzNSSkUR0Of8ZU9+6CyInQXtTVrqoH5INQzHJ7Oo5cDtO
lGnJKUoa09e97VytFSxut+LHTTLeiaZzFE5t7pt2khxmdatlbByMRK14HdX2J1pE0f8Qa/xVR/sB
fyFjqHdsHasChRjruP3GDQ7GrZ98GBnwoQNgwW2V5afFT5cnuj8wj1TYGaqPt07tdzpCYDwUnf+k
qCpKyLG0B2b9lQagPJjcAULjphGskkPipgkqbqbQlT4AvCPIg/J1GpJOoLUcxgTZO8mp6kixqCFg
aNRJNjl0U2fwUAIhLrDBdGPhR6XaX7lAVPUaze0xe6foFhnC7+lxPa+00jYL2so3oY70gXRbLZn6
qk71nRF1MkrpDtVe88IxKuzOGsWA3EnTqlLqUaFCvVSbPoEA77oMyOs1i3yNbx+jDwEqZL51lx+A
8+8onLBBUnb73T7GJ/06SogUERGSIuRRKH9Cn7kghEec7emOiMHC4PsIukkQ3CylT0LSe7Cv8O2o
OsJq46NP7A/yP+rI4E1wTfth08WtWBoY0GE3ItQZzzSqTPUS7xOewe6bdoFSmb6YCnpUe3OtVguu
C86LdjJtnlkkbR7Oz72fQrO666MAHKFv33NWTyU6GifKVTtCclxWfcY80bAdcRD5cigIl9l5kYck
k6PmqsFI6GzDVY0FBdCRyh6SUgjWOOShRJs2dtRnjSZFebA1JnFdKNCOjBsjZKwCF16xPGgtXuRq
aqdwo4JjtXJDHdvLlztUjs+vUTg1HX34kx8B/yQOnRCGqyoajpuYE1X8baTY6A2VDRCKJ/DEqssu
El9qjJAi2UITn7jaOaJXc2m1KyKQ4icWdsKKtE7iCI1Qy1VD/0aiPC+mWDuyizChd6hZaDOk6Aod
KzcFbHvpulWSZAxDCDC39d4TK13mYsSGaAQSfiz7MWsLQKrBAJnmyvwm59E8X9ggpbKAPNdVnNI4
APm+KTqDEkkZOb8fSXfNv8Rvxl2cP4NWFiKv/wc3L+T3/0+LJySJaCsTNEy59udNwUSfRAkO9IXo
vMZIrloXwzobIBBHlW1VIXL9lXTyNynlY3ULF9PejGRi4PmyvTG6+pQ3rW6OxhCLcWYJvQh4G/JB
Ni3hq2BODgl4sY8C6Y4U1lK/BVZxQ8iz7hvaiIIhvPD8Vd+D1O0v8CCP7ULVufSoEhQCmbCUz9m2
wG2W2jz/foCev6EIeovvUtyclSkEZG6XiCaSX9iprqy/9K3B6S8f+lICn9JXcXLPUk+1B6xo81Th
Nnd2/RbhWVu87nHu5s85eir2Yv3MnKEry79v+/vvMvC63Cw0Pxm0BsytiSIcPPUizcc5q051/mxV
fQewnIAYoBOtoRwpqBIbMDEpO288kxwJsU85gXEnjoXLbJnqd2ukkeOWWno9aHPytPCEbNBNtfeb
CwWvzoNyDtGTbprfvcm+H1OeopwBeNmxNGOdc9XVIKAj7Ywiarfjg1mfGOWuIsJzKHjfh3peVcSD
hWfd9GOA1KL3s5UxjQ7hF8FROKiLPZ5AB42dNcx2NVGaYt10YTnedX8NYlwXHHN+JLMATVfeD1jP
KWCPF3VO3Vuq4lZtf1BLw/1olW5DSWFGcTlIo8ha7ZL0ginvII3GGHifsPCyR4kCxeIqLivoxtC/
NYM0tLiiB8krcJPBJuxoxkVKTE6+XTH5wux7SNTe2vZS3rGS2/YDUZH/Bm2eySMGwaTesUmuZgR7
op0R0qJPsLL3hHQ0ovEdkMo6KnVOdPDgp6sYZfkVKFx7qZA7DpjX6bvSr1fpVHBFpPOzt1e72laa
Wf+q8HrqZitl3gpaXqwaBjZEYGy2689xqebxFUdCute2JFYS5KInLS+MAMoozHisZ5soNlSesV5w
Ls6ck6aLOtLRmHnbBHjugSwt+jxG1vEjnYDI8jfJcTRKgUP9lE1KWaZeERe2spUd8TafOT0z9/E9
Kg147lAD+tg82AjQjehOSaA6FvtG6QKCIVz9UJWTCIZwsiGX4/x4xSIBONnQFwjZUVzba2O79oDD
WSS6jskTq0Fl3MWZaJ4UNLPZJMREMttS/r+zb0OWvyMPVqAXAe2PiJK5YU7s0yWdcLJED/u8gsUH
0Zd3vo3YHcnF9GEhRouVnh12ZFcrHe5C2+dWH3CJytNpCcdjmO9rndxAZ/7/8ubsrjdZAvwZoSYK
XZPFaZ4WetnJ6zq78BH48EhzKmkI0wTLVazd9yNtxx0gQhRgo/W+Ddk3F8NG2gktpGy6yN2/Z7jv
3N5YO1bvgrbTGQtKMsKxGf2U137XNZL6+GHNX/2qHpQ6pjOw6jZxH20S1Lwg8cfy6tzpImAaWmfS
B3Ox9+P5jZ1PZxrRBXhnZ5UFwOpwbRQ/DfLtCcRpxf+fuQByfyMZWaDsRibxJB3ER7JGquyuo4+X
cvPjxMbEgBvntq3I5BVwHdkdKdsZQB+wQY//GJ5WIjapMD/AY4F+3umytJagJtEkVMhISihHlXqs
QyxK7hWuji9lp3+U6uT6yJTVyJr0Vh2cX2ySZFaDh8whJW+qdTe7BauCqrF5SwSarJwFs2Puyb+e
Od1MDqkb1cuX9HyUDd/DYtsozWiGu1GHmJFRZjJSS2MIv4Ql8qrvqdgSkyMwVZKYm7I2+0N8bHpg
n5rHPrYByBZVGlRO4aBzy1HjJz5CX59BL5ONeBAY6NQUVKrZVXas1p1ayfn9X2aefA/SiEQxFgXs
buVrbkQbOZZZGj8ZoQZbpDvr0WcyqTnrvFUkHT+gQYOvHIor6ROyYjNZjWOSZ6azl6EBMAKdDUxU
k6r48T3Wrn5B7vilz7QLS9IEXMwGyOAMQCsxHCbfAhKlyQGzIyzJiWoqYlI9zBs0Ug5RRp7iV5DX
tfIUqzmwzYRVqG2GULta+0VpKBx+TJ2mRe3XzkukhVXEv7DRLnoErj+tMhhDeOIeXjjfXYpZD9tE
wjuW+l+AShVUAd2A5msJa/PPDRs5aidmjH7U1oTrnCW1M3JlgQt1HRUCNzgNE3nHhjvYhW2EkpZ5
jHs4wv5/HZTxVLNO4KikdFSpPZvMcBjP+TuirwFkkUxgQLfVso41Mw8xbShVq2vg6HHj49nTnNg1
rVfAlIfNcS4Jb6vxp+jdqh1oqlhxht/u1nEtdtOuflACcOZV+LkVJ/p0Qga/GURdtXJGRkIdVavn
DCDbyS8qVt/fMUlX4f3/O3pHOBP5Y2C0HNaUw6f7jTzKGJYlu+dLFGNsCiStsSMD7UY4VffVoaob
SXv3fsXsZdYymJfRInXLrwfsntd7l/EdR0b9aOi/lnbijgU0DI3mc/sxHe3VaROYUbPMxtEqrYe6
DkpmXJ8kBZm//hQSZZm23hJ/WcSUP4sIbnDG/jeKy9zRML1mjZHYPm9v7sLKplSB8bALPtyYPqIO
8x/KLV0mstpj3CkNHhKk+IogXpnF0Q9h/UqReAQOaiMBz0/i4znggTF4s6eK1WJZszhcaLA8VVJA
wCtM3gKULy86+2u1BjE1WLhDR3jcu1yURomxFR3Y0LzrMdbhFlCsW7HuSLUwW/pIyIT2ETMsJtOP
LcurxD/cf+uQgZgklZt9x6VWpzDY4Pv4AWwIJzh1eKuBAe+L+aA6Zy336U/1Xqjkhr5B5CE5b1CO
7gzTY6nypBpOeYfvTFBooQzizqVatSWIBsuiOaj6nMziS65RidAiAIPk14Fv9FpfjCC9kkbk4tKI
NqriaIjr8y0/nN7DsC8hX688hgdj7mvrZjjWAY2IrH4FUBpbwaeaFVjSMqW23ox8fB7LkgRipBeH
C8/xbQmaRu5M2B6a2Y2ZHRbWDzWGeem/eDES9v0gFKJnTxoF9rr1SO06uPlqkYEaE5UXwjRquQgX
p/ciE58f7jfsHuajtGK7SA8LRHTZl7DLouzPU1UDw62wZ+/BHc0e+sDpgu7JdCW7vT+66GuZvlHP
K0GaqtOo3iOWOmqNHaEbToSeT3on0QCEjjImaC5625Sl8QJ+X/QT/lZKz3F9tq5QN2GvMAAw+69i
JHe3I+qlWNotmvk/8Ar61TqH+P9H8PrOuMZc3W1PxkXLm9IqoFfZh/AMd1lbCTw/0G/zeetKgiHi
nkLrhoJhFlQPm8bk4lP4OTBxl5n3BDgG0TrT26rBEHrmSnlbKCycJKPjkAcyHp5/N5ShQa8cOZld
H1bMWclHXkQX1s5Jlqv+wqgJeZxG49EgLKLth56f5YK0QTYEaH77iaAndGtDuRrMPgXCnj/GN+/Q
kADf5QqbV8wDJ7dWck/Gn4ZSEgaPHeMNNHEHY39h6S5oT1P9WqyoPKZ1sI5VbJzW/hIwZR+SYQ0S
e9DFSOjJH04X4Om+LzZWlsfBKcET6fVmVpTv3MJ1CkaJm8j8uFb83lFveogKdZ0zIBcsBzBhqDVC
i3rIFvKD/IonjVmyvL5/Skd/56hf14zDkNuf97+k5wT6OE11yhSJWGJMgpuFOnr+8rE54ICpRF2P
wQ8Ax9Lgnu0t2sgoftnDjs4ycc7s8j4/+u1Ac8LuQo67BLg/LjT7seBpRgbtMBCBQ215wo7jEb3T
NSNDCrfYOq+LyRmHyLK9B13ZQu0oSnp0vfzmG+Gx81dOTljBmmlGV0XVThTtD5xTr6rxnO8KjBRr
Vh55ia5Y9ArTI/Uw7M2XnJPWzqR2bpbgVkx6sL/fTQgA5jBbpQlJ9om/X9+tpptSZEQVMcJ7FO7A
2xDQwkel+7Q/Owgs/D+FJjdXg3ejGYX9C7rm8+scq5Q8sPE3U4I3E3os6QP0C76KTyHtCBYx7Hf/
NsAPyriaz61iszAxIl1unOB37DCtqI36PQL3Z5vqvoFxgdR9kkehQagxGEM3dxTxD0UnYk2p/q/B
ujKvGOrDOX//K4cBjwxcbYAOtET2ZiDxXlfr6OHSC832DhUOCn0ZsecP/zarN98UVL7+qpnq5mJU
gs6D4Irr19gHMi+OTljOu/DW+vdMWdGOU937quuVBFcQZVFnH7f3vAITwz45tqz0FrH38IRw0Nan
rjDOhfrhnfDWumYJaH6/mrEQLCnblwd68OAO2TuwArzLU7/FsNmFjlUgzci4tDrvnXP88zn3KILg
Mqvzdqy+EmNIweiYTdjyighkFhWiyc3bE0o4bs5FyNE8F1RUW3+dfCWUoUjv3QsCY41IdSr/WO6A
sbAEChtZ9yxW4JxDWd9YDJtx4PUQJZX7Y/H48oZop+Pfsz8m6x7CJHZgyW8zK7N+X0Ipos12zwnt
5R8RkOB3S34pE/t0h5428tYQbyOsiEMHGZAehRFLt992NpKJLeuzQvfHWjtZQZpB/CK9hxIKtbcQ
ppfEniEbHPn/WwKB650je/f9GNEdHVfwZRwJGaL+OMx2ew91IoecCt5gKSsfEq+P6P405h8bjRZ/
+uLvWja9+3yJ9LBLdp8/3nIzoEfArKsmhfqwOXYIL5yCA26SOGM24KufSktu6DAouA2hBLqEoWaG
A3IO0FiPpPRJl4AGaFxLtaoUrMmG/O/oH4XiI7Pyi2FJcsN0OdkcoCTml5X+iukm/YcKVTnmhcAk
eutzm/pCNPfnUtRAPGvsHRbHIJpDVNhLzHr23URZGvu930K3ft1x+FUbiLmfcZIxxozBdpuOZ3Zf
KGfcEYt26FtHbSvkDrZrhZdfh1u5Vlki+N7YiooZpNW2zWen8feGNLjdd1VOZlwLnnBZPCKXTkOw
8Uxn9WYJ51jICrflFjksFdhRLA/qZnEUir1wn2Xc7jYmVQ9h6kwHlLf9EGbE69vhUwDhk367vUm7
0r2iF4X8+qHQhcX6+/TxyfG8WLx6QAOdXfeLlrlMXN+GyVtZL1QEctQk96IbdZaWhm7XZGUK5CK9
/4DDXipytesJYUYorg34M/RALZATlH8sulIS/LO+A6DprbSdVqC68VmrD0DYhh6kHgaHtWugfjrd
wYjxz7oIPqQlQT7ww61LR03DIpz8stj16a1yKV2zCB70YJ+5WE7rx67THCytLUq+2Bya0Z5VRXYF
C7Xd07gc5yrmjZtkvtJgEBnfAx40s27xXwvpqdeuXhD2zx1m9wCtQ9SUeequr1zhSQ77wSLaeYLI
PiITM0qy/z7Of7AxIGEc3edOb53IqWvkUrHPinqan6ClPcrkoP0nj+4Kl4D3gTH4FylehP9l3j9z
5C3KMPQ+4ZtcbSTm3z+Bk2ItSQk/qKkx/4SqAjw9UmoMwPMbTSv8qSklHRvBSIigmaWwgfOAtisa
kQJRG/fm29qn5q39tT1tW9QnCYlcsMEdzHf8qhslzk1RtL5AJqAAYldu5YzLKdeSttNPVvEFWD4M
mafP948TW1CQuWA9nNDymZjeYnbLIlsLNUrUYDy7ztArNsYZf4dTA8l7uPBBe68XGJ3AB31seDcg
I0Hjo92gNXKzmuekcqFVSOudnlLk6OSEZ4p0iv6AzqCry02WwhQ5NLYVOvGB0QvjiKJYYTA0UGRd
RcYYjON3QYNZbh8Rvsy9JceCxsHKKqKpWUu0Zg0youNhS5orTPMMu5oZQBA8/JDqdIXfAmIoooz+
98lJmv//9PEmuM8r1vnUUJfWsef93TachpPFyjJxc+QJ0XyI8xsYOdVPbe4g/43kDfJn3tUX25hi
Zv0PMbM1db9NenlPjJ8CbmVKV9GkDJIhPJE1upsnl0IUEPlf/u/Ak9075zpttDUQBzXFQgBwK9aI
GHdX7lwOwL7Bt76muebUaL1Gqdg1mOk9U07me7yT5Wwvysq2WtWjb3vyEWDoWvuUB3xbqKWRQLow
OPWrngt0aKGMdMi7oYkpZ3n9I+saHdLn0XbIkv8s8DdobFtbCjaI+dM5XC5NQR5W5AqVdQOznn2t
jKA9FEGdTotuxW1UgmvG1ugNXUwIIFRr6hteDJPA1ne5wcY//+B5Cd5YE1N/OhZ1VvbXwlxxrIcT
AlXAe5lUj5zEQF10drIH3S+OqOB28tZOFq4x24S+xD4cx9NQAPYdQ7mkjt13q/84S+9/XACopAjh
zMf8KewwtYv7GHoYx1a2An7p0t6NRl/EXvuyrotn86v6ykG6gI+wHkExVFVtyKonq2lQmQ4M4470
QsUgz/c4nJQO1wvquKYqnd0X6Mu9+c29W24DnE3yBua1V/3CATDa761TXKyKa1FZZWD5wDBbnEPi
sdRMa5+VTqPtridhcvM+jmGHZllsVpCtmamPjl4GmR07zeGQkzwO+PUImdMF1igPrCx3LsoSCSg9
FwZYHs8bLT/girUfOg/dfDWEvG/W3/FZ5e5uR0mvGWUp1M2T5dbsK+VBVlq0z2sgzIktMV5F4tPJ
XNfJBFzGGKXQ7XOC/0DCDMyR286tpxHL93PGw15NDRRFzHZ88lkCbRewJ46WQOLQjXqpGBmjA5yg
z0NSdjkYBI4PdgAHGkTkR7tBzVvbOGeF9Zs55jg9D9jSIg7hLDWSHKese1Urq/upE3quxZMNxZQZ
cpwWFEduk/tIy+4OcamPBKym33Gddc6T1LjPS3DAM2s6lriQ937tmv/rUl1UDlF5ZLRcGf0ITELd
qTbasuCZM8Elr0iVIMmcNUlNENT95tXZKPpwTLDYTR5LbbiiNF+UNKcS/SFWQrpn3Lndkzy1pU+r
auz1gRg//7riMjVWojgWFv98KSwk7QbZV+QPucDeNw7Of7Lf5z8CAjSiOLt8LbgipUAGzC2x/wcz
0ZLHCSzi+84TA8lFj3l1tRPjcxSso5xyVHg2QIvR+gR527jiVFI8uTLpsBiLijGhsP9FT43TeM25
G6FWAyfssb1hXOCjEty1C1osptttQWYL+Vks27NkiRk/Gn5sR0XK7i5+qkc2NRGhDWCluZj+hjBJ
UwEF8JHg1rWQeCxV/ubAf31Xb30SPW7IriUlwE3MVLjdJaqnTgOSrm16es6++/HHh5s2tOJhIAc8
oaSKDAfU3SV1OTYsqPIW+OAUixlrHv9Z1KBbT2XE1/QCKWhDxRFmabwBQXLxfleX5/aaAc0SavRv
SE0iDUdIW3jffGxQX6FE/te0n+9uStA7YJa9ZN+18l6Uz1rz5xZEMFeZnqBXcvINPf71ngJJGRSD
KvLcps/QGfWYMF+1BN8kyGtWM/a5am2D7wfDhCV6ddTeAnNLgCYCZhly5DCnTE98M1olgNTUQVCJ
INbyaUe5SQxfv10kcWKfRSQb/BW8cjv+W/3itO5ayQM7j+uGxyGiT+tDVjqI0C3lwGgma3avZlv5
+WUDG42pELsrHeVf6sD+BoXDqNp3P1Ke8mtz6BQlmEo4MtjZ1w1ECbfSCKMzxJBVs7H3l9bg6Kny
BpEFZOZQk7PcWkCqLKNrLwZ2dtC3ZGy/6ZCfcDWvv4JuAskiyD1xd8nSYz1746U/Z92jaIhuyJoD
Hx6nI9C0HFYG/Wmh4uI0kJwKLV/N6g5f9k68fje3n0+0lGz9rI98lre1eHhOczcJ4kLnXgT7OQ5j
++vLpKMi64iuKS3xEv0Akg4xdVJkbh0fqBEcJ+gQUwZ1pCvn9DFAi+fJQ/Ec5MsBc/zgKVGeEVr7
0LCuc6ycIwiTj77KgFors+qhCgmgZUE8RFKqXfJ0NBaNPlwts3V9eJBW6kRb4wL2T0CiPE5e0Gce
KokbPXqCHNFelnUJ5aqvmSxiqRjgjZcgp9Lw23NclTc6ReqRMsAv37L1iMo+7f52hyRpv9fMNgXz
9FvyrL9bSTPKZ2j5XmhPyFqo3F9eps48wNJt4q6erMZ40S92poK1s28qPclFX64NwipiqalOE7r/
Z1KDEDNyqV6zJEkn82Y2v6a7Rha0STZxllPHw0YYOvALsXQBgKJvDgufqMdyKwx0QBA1OamcYbOG
KdX4BmkuDCJlWDbPKB0MJmId4GlE1Q93OE7S7YkyJEAwGkjgg5kcWjZl4dXkdQKz28sUr8EpfnNS
LyvI2tFKPwNVpQMOozdpqhqB+R7aof2tn2Ifw/lSXvYDhdGiiZdHKwwz6BL+eVnY0T2iFMldc68t
epydcfcS/XjZZD8rOt4JPKw/XWpIKOaN5cV6VDfmGDEROd3E/bb06DW+V2ycJ0waQxPGyN4u+XHr
2E0eUNAUAb1QxfXbUkTMwvNI24XXjn1JSwMqgFxLsCWqwpfIDaUOGb5QQ2grVKQOgfkoWIDk2kdF
ktt4u8Jaei3mHN7DZ2To2RweBUAQa6r4fhQzN1o1IJk2Wb1e2TbmVzy2/zuw289stOkS8FY6s0Gk
HnDGSJa5FIc8skQ//+8qnnALtrQp42kb4iB83Qw479GPtGiQJ2iAVQyXy2nuqitzdIVONo9U4h1W
AuS2BHaQLOfotIX+hSPqf2i4CVqevfJy+Fdzx0PkNU20i4BF/S/4iXQZAa3WICvMtJg+IAPnoU9o
MFVs+V+/g+9Rg7HpsozNOI1zBkGgCoqswSRG/uAeS53BqO7sYLrVXioKQQIoeFq+Q9FyvyaBTIzP
QyvivxdQDF0PBPnGWQTQLl4XvE59F69oK4aA+gnj56aN8iQFvvmaUpDWWgq+Hfmt31dd5ONKxBRg
Xj6vj3nOpudDgAHO1utHOCCWhaB9YA8XsaBa/BUABLhfUfntrA+tRUplknuFii0RTPpQmuOnD2cH
tRjuLMbJroGpIvXksumRsl9Hw7A3ANpmvJHJmEC77NgAyjUvldh3WqE1ZPs3mdYjbjABYOzR53EC
Z0KdFoxlFGdVNpnzcxikrVVGbAPp1G54GnSr9yIm7ImXq/Sn+Ik0/hnzWhKFXieVfCL8s3vRth+a
L/fvmnkH/cJp5K6FOn6VWiDgYbLYRy3cfRoA4TYnCzURFEZo4NYWdxAaqFyBYqOId9g4S1IBB7Ku
0EXZLoV46mSi9hI4X4gKYl7O6GIa7KyvmGyccRjaNcNxjLKMGDzlYZpEBq8h64FN1OOCfe9dPvcF
NP8GLHA48rZ3ibtIgObgsUV2oxw/B746ppBVM2DRk9x1f4xrJwSnLe3uT3+AZkeVHzof1Be/aics
tPLAMm2XNcbosRDMMAroeIQsNVDuK1Vqt8m/N8iEMz0WGE2MlyAjoSVTLNKbaAkfs6xchEjMn2/i
PUe5GupgnMzKMWu6LBzNh674FOYN9PEJFQ7F9b98t+2NoNzL/g5G0L8rQkpQK1O/UovKKwUtK5zM
ij+mdYaNOsYAxyigYdlxAAqgYSbeqIsz4L/7cMbycEnmbXzmnsMLrU5TBJvK/mAzBcyv3O4MOKOa
FnMG3oEqcv29bVis1IGpAcBaizoBY792NM/Gs1ba7FBIYKu5k1Xh84sHaEKTLESZe3LE4RfeoZDm
l4cKq1eqax6Y7D217FWUiI7x/+u0szf9wt2IleKfXUcBxMkn/YVmJFUSJHxQNUIhROoyo+bT60tG
1WvUFzO8Xuv3UNIxUzMwMXGj9h41bcs+lTG7O2AcpkMnyC4Q5HTuj52TPajkcLbL8x6EGnG8xs6M
tmhRgjMp7SDpvsTm+fnfdvUrp2EPPwfNWzYduKJ+P2k/ao1gHgVzlrKaYxfwdFe4+J+wacVtQ8EB
HTwUqNyM/6EVC0zT6FZaDj98ON7iuzBK3Wv2dFRGsQTHuRkoC8yaMiXAozUAbqJyTuqgzNOPXnet
QVaA+ER5GzK0ni0J9/d0UXdsfx2qyNhZKb8fNafCmW+ZqNryILQoIM3MLJ1+V7GR3LKI06aWUY3h
Q9ha8SOGBxUq31tNbkPWIhybvE/LDXq7YvHX+NB2yHEg/I8DNdFnpC7bbFJRGSr6D43ksloV2XD+
iM+lfsYtaz7XZ5RoYKuGTVrnVURS4U3xV1E+2jKbQYYJ7H7k377NlRu3BXE/uqVXgb4AyZxBzuuY
cDoQujTOZpUA9n7Jnlu1q+CJJpeSlWUwWrgWauwzvhgMhisrmE0jTNbxBNcRnyL8CqQRJiPQ002a
gX2hmthI5Fps2CwFGPyQXozSd5ErxJ7jyoYALqBXnoCTngpeWRRC32Ljw9v6pG/uUjV8sLH2xpNC
WRiMhcjd8/FK9IpeIiIlIPqYsnwX9jnPOue988hmR8aBLfDs7rYqBXFkU1Fn9y3VUi8HSpTLVsB6
tIdwMEVFots2JWvReDhKh8i4dLkkOjhf2qo30YcpNk7q3CUhzBSYLYDDq9v9XcqB6WUI0BVkQeyC
I2Fa8siRATKifs4qs0P6nUAlKzn9S+9wOO2ELwtzKp5Qenx/f7K1Cu/vwXZp0e0qKWoH3GXBMzeW
g7IsoAGZ2fyaxIWaw5ki1mWzAlc+W1takTbPcAnOFY9glejMwys7FriJS/7+TeFbz3OzLt+fCNK5
H/pqoK1b/MbhgCqBcDOBdoAO+9uOGdHIenuE1pzNLZM/5x1gzt4p/D84f5AY9wPXeNMbvrZ+d+Wm
AhLVAkMFRXrm1jBhk6wRheYoHnN9gMOg/ajUzGjNwbk9n0srYY4ZvrTOYfiex3kjQy6b4xdB2uyI
B2/0DQ4zY1fbiMlAjJMxK1f/HGpJbZRQjRwnONY70HbtpO2874NXfvEfpXyoMmeSZXQ/A+PfSQXx
omz5SmSh65dLQbD5yDGoP1sYf4B5C5HGaL2UEPUhkzIrXeUviYulE0Ec79bmJaTIcnnR1DuBuhWn
z8WgvzzqbL/qEY/qm5JDwSAuvGdX7fqfPvW5hvynA8XqZJvz89aVCNF0bixwstMkCIDQvq0D83pN
a/xFVoNX6+f3KgwSoDUAFLn8KNBDcnHmeQj0zjpfB86hkdF2tuvjtYnAf4mzpYUPJqKajBZJQaBi
yqrwFZWiYKY82fEHKPUphIqBmf82QLqhGf4XJPewvHgLwqLZK13GQyyr08gBzfuTH5Fl9WI6cKz2
dYTmnvfOpFdK6rK19qBo8tyJvtx0Ue1iS/ulZKifN4mlJIcqATSAP+XAC6+mDj9uibsW6OItl20X
xxz9nesOlw3MERchST5SemZ0Oo0oThC+zteIob3Fh9a0vl9qWRuFlPuHGDSeajE14oYDfJQgBSdZ
+V7Bfw1VoeOvDacL7YnI26bRWSsj7zAVQMyONiAFNva2CgtndIjb2mieA42H+BrYP+UkbnWYm4Vs
uckpb64QWudeCn7ot4Uauj5JiBFYV12ABONc76leQZZz69W9LYgCPi1ZMaI15wxUtLwrk1M0rjiT
hDiJAepB+BC00WVi+O4Mgbx9nBRfetpq+2/dThFfuU4l8O6Z0BeAWbDMTcBYKMC+bhd3K0hE1qaG
KuMwoGoGpFHpQX6m4LlCPoEEzbL/bpcuh4z8ej9M5U/5iI3W3cMEdmaaDqAk58pdgsEvh2X/Vqwy
O58EjbY0qzOMQbMCIqPIy7T8XpaYsuO45rAKwyL8ZXIitZ2W0fZMb5gHnjjiiF/Bz93EAtfm+cWF
6k/5Iv3zE8pEM521D6npv9PEwcdmjoklwYr6fA+/XaN0v3fXjS9SZW6O0pEus+KyWyOqo76BzR3T
1g3nmHwk9Got/651X2P04L0A8oUCkXvq5KeY8i2Q0glDSj+VQkrJjmEXkHDh67kdYhVfCwrAzT2+
BwjRGrNgkQiaPBko3YIegExcTnJiR+bFVntp31iBOCneXsOYw82kqn8q4dATWee/TvJXDtqcIXIS
oulTePG64ko7rIphpyOGKskpRFH+7gMNweqS4Krf1Ax0t1D6pFEzWGBa4QrFyTpj9/Xy2KKMH1Xu
Z9TfQ08yARF2Jagi5jwWomflU3xMrT/XiI+tfV1X6E8ru9r10xmyp5piy80g/YKYWmZ+t+bd+v3Y
djLJGI2RyWWPuivbLoYgEz4NRTnm6ozCLZXFXEYP7XoFEEcSBUHtRuiJh67agp6fcEzx0+sHNQg8
ZKMBihIIipNPZpS7hN9+Rj8RF4DvdyWiA1t9oEo7JMU03sQ5MJUOpdANr0dLeKoa28hl737BDvNI
YCBTYlqf0a2h73wIlIYW2ykHDZ5z7N6sR486IScI6L5jCmA5KGwhJ55oFZD7kPtBPXNlGPStPjlg
mok/DSQFbSrS47OebB13ulkG7eL+6CqePZdf0vcPtDMMJOrbP73Vy3r18aANSU6isgQkbtyHajn1
Q28oI6jmEqZB9qZ5Vj9cb+mgbBi7YxQaqpfqejxzOzuQIdG625O9BRI0uSEhsZ8+YnA0KyeXZkSM
DSqy/JE0UYjZGk5d7hspmqfW6LyPFzRbdahS5DXePajL5+9qyWDQseDbR2cNiaIpq+LB6BdeCjkU
Drh3XXqgqC/x6dbjQK2mnLTPgEPmb4vDpGbjLOBCTN/DA4mzv7bpYblITBtXzuxLAyh+K90xoxVW
V/VMVoQWh78dZFQauF9E1Gkr+nkP4os33S/b9EDl7eloDUXaOMk8gC0d4Kvf44yXqgKbkyaoAUxl
DyW3yXg/HoNTXXD00u/2f2RCJCOSjG/nPw6wIDVDvu4rDVCrb0+IRPMhVYa6IKhPMOl1B7xs9S9Z
ETK+cZRUknvIjE7cvoIUbuBoaxYGr80rYa6opEcM7t9JPYs1kC1QiT0tLocEHQhCYdtMIycSm5Y7
jMvDh+NkA4dn4SSMN9YAyn9JQkf5eNPz8AYTepq+rHploHo96NBGrFkcHRlVvfE/HmLO6D5ibqNl
Xdf1ZqwqugZ3zaGxtg92elNlGkYI72UohhG/aPl+eAqdHjwWzaJYc+WpRedb+j4g56D66NzxoNwg
m7EqhZCNNn/QYyt446QTCQ1mX7qIRoIziXuhj5H4U+Leq6crllCh8XWJ70x/axUBgmP5QOHnDPba
zcOktRiwJom6PkuhhHT80NIH+gh/ySea66WtYATG/46X930lNMzDej09VoaB8DqGkcD8qM+hWQ73
YdbZW+FczxU0pvuYMY8VhqelFnRDL8Caxt46KtbjPfHiTe1r5YCTCqcZL1tXNXOMPHz974tF8ZB4
K2KGkrsgZjuWUl/IJt+bWomCUX88trnjjWtwIoIfTplu4HVXW9gTZUzvTvg5BOThF/IfK/tipgRZ
/fDi5sQBP5lGWwdjCkKK4rmRqAjKAXYQlJCsh2RjToEx3yQJjh0xtUqgmtzwk3anYiw/1ohyyP4T
GVE9RBpC7K9uvbVVMZtgHn2aYn6qcpX4JysTGSFkF7FBAwPWmpmaOGdxC92GkcpjjEwjyw4R1OS8
JSkWyPUiEgihQWKpb7D81YjR+bj3q0Ncnlqp5pga0f72/hKeSVeBbk4gLgDAgB0nsFQF8qxl21y6
kAYQ7ZcKetQ9Cg03vFYPthAvC1ZjhWAI6i8acFaxnaIPDfC+7g4zXTkBLY/7rA1nWxJKaMh9TVlR
TxqT5ByE/i8nztrdtVOENY/8s89FeHItesadmgqpllMaDNvN5XVw+/9RXRRessP6E2cR63I7n97H
y9FsxUnjXJrUUd3fuXY7euziMMaose3RBQLEcpIm5rlenkorg5w7Ko2bPZ4dXUsXd1devAD0nSOU
Kvgi/qi/2oP4qXpsLVNsdYrJCoqEvwLRBszHq+YSB5QSJ/yE4f9NbbH/NtYoKbsPTd3s9K2yPDo5
djgnpFM88dUSrOB0C8rlgpJV+1KAnddKXWiOGYqSQOc84A7biowebwCXpaCVN5ZH/5jqZ62umywn
9kiQy7lBRwz9EVtZ7LvlB2jMCKrQVPPBzJ/+wlozneEEa6bR/o7KL3sCxOeeyHDvFHVCvnKqbp75
QS/oHJze+qsdjseYXm/10ODDTbw40vcRZcDtaNw0e+QILARdCEJzIgZ8lP+bjieDuC/DJ5FqUdoC
39PVZdIg6M3ySk6l3oUllhYsZAagEkh//RoOpS5Kci63IgeYb06byGO+OyHj94S00mpR/i4GZuco
4QwuFQYV1ENPQ4xD6dMb/besXPjORiANgIA5rz+r1oXq9ZWAB5oy43tOxMZAZBTgtlrw67Jq7dkF
GEWw1IxT9x1EA/ssGqQ1XSgshjTx+9QkuimKobjjeV+4DqZqnnrU0ENV1ti5QWbN7TSpsNQBh8ky
CPyj5N6ejP88QlY+KZAMEdKfMIqLutZDwhT2oJlMRiqM2Q/hUANoLm0Doa6XaceXD5ojbT0ikEY4
4tgKKcwa5+UQEnztBrQat8b9eMBg9+Bk2HWtBoBWH9OYQ+/rI2G1KNqrQ3QQI1jPTyQiu0Jo7a8z
TzpudD04u9oilgK4CmZMIg8YTFOsc+CCloNnR+qOETRxw1qsOTvfbx4sPWve5rk2MMHnB9MHtZVc
I6QpaarC/ZEvury6aItA27LxxENJ5NDpvwmb4GZi/huyEHlscBpfilmd+tUn2BJE3AgqEaGtUy+K
qZsHrhTlctvWLxnbNX0wP2nrl4OabQJShr51JKk+onqLtoD8Ku8jOmyxv7oGXOm+9O2C9JboBEH5
+oXT6OdECjUKyem6xpSKqTN4itteM3Z5U3Y+Fjb54P0cq8cxqX4+eOvrPtFOWSdpWYJEIEKs0mfV
tbbw/aj5fLoyS/qCZwHhoRQgfNoEN8D4uOdIWnC1M5bfWs3wB/+oDbkbmTIOz0YSJMUMos41o2lG
yL8BS+PpxXnTOvHpFtKs0hWL+dya4xwb/k9176jAHFnNLr2n8wHNq2iXWofA0eUC9dWSXjdw/fnF
vq8tWXKhrhizwhMtHzsVnUF3u9QISC1QM9LLjnFcvIi4DUsWLeYJrp9tnBzaR5TjF+AtrNRuZnKz
no6ZZlN/z6oEvj7y9P4YvUGntFcMdVk4Fbtzvz4oCgtDO8JXNl6dHzdgoF2fKDtwBeH/lxQB8c24
Ax3U+VuRRpEbOkQqYxG6MPRum/+qdgHyx88tPpvd0WsgHrZ9EqdUU+5zpp87zyIxEd2hgs30gN/2
h7t03KdZH/NSalqPku0SDWkpp9hJQf0/ZqICHNiOJDcE0JxoYu5n697heamqq3TmR2CIr1kKoyAV
deJMymt8NE0j8o2OvAAVf1EY41U041NkE1F2cUX0A3BnL0i9fB7caD1wV9+hLNrJ0NCh7MrfmhAZ
NVV4GaHoO9XivmHpnBriDdLb3fCjT53TMdYWxJlUGfh6YchDxw55RE5xfBDxafOIiEiwNY8lZqaT
q+5QhAqQPTDv3r3jLmnDuuu8BfUZt/ASV4LBHA5RXer8CBKdShKQPL3RrBSan0mj/hoVRtHrasVU
eL9iLu3VK6Js6LU/LEgu2R7dHcEEvUKELpAsk+9iXGkhHvjhE2MiW6Ni+pIZt/fLh961GpNdNlw/
8d0ymo/lMC4JwhoJFcDvSkIYMm4FT8B73KLzY4Hn/bgM01cgHUkCACy41TTGqMDmXMGx4xOX4n0Z
21d6785qnzubwSYSH4EMKAlHtrGfDqrgXkJ5WcnN3yIG85jWnEDD26WyVnSFWT7VUyLf7lVlb6u6
sBYVPxdi44R97JO0lXm9ptPu7uLZyZyWWV3taKNyNVzOF+0XUyz5zFhv0Qrm3CNYIp0n4XJ24m/I
RddMGywLArE8hOLXvO6E9d/LBJLnhtvOs8CQjYUgiFfLrGce09YQL1TXRr9rl49Cb0xnM1yqZIAu
RUjZJxvPSFUe/6v9cenKCc1NN1WZ7OvW4NXBoCyNVQ1w1hrWuTcAqkn/19Y3eQ8AkBi/WWrGhsUU
wscXlhkAWHvGOroGpYhj0A1fjiEUF7Upd4+rg/6z2isvaER3OS7c9xXpYu/WFKrnPfMWU6cguxtp
4j1hHCWyXWwHd87Goo+Z59a4fHnO3boBtVSqhWYDprwU5gO+U0aP+TD4jle/Wt1pIs7mQXSOMCc8
/uDtau9ijscD0nBD3kAtM6hEqHcx4ZF1lKPYyDufWvncL/dTOYOdzNTa9VMKC7wPWNodlfQI+iui
G8eI2Xlz4N9W7eqyvPgZRbAktCr8qGDYZFokuxZbB0O9zUTHMaGpLQOzwNJ3ijDuHyyrcSFMTKmM
7FNVQJxs+cnJo3r+15QxFXJlWmrbdF0FhtNqDtXdb2xI6NcUGLusFN5BRrDC1NcYfhyw1NbF8Pv1
U26gJ6zR7Cp2Vz6WPvpsnqIXKPGB/GaJnytZpe0b//6Aa6iIdVa4xXCXO7273bAQnmcxA9hG4y8l
S5dYXHG+KChr9uEkQqXjqdnAIyoQxrtRdqrAjh5XEDa0I3Rh+tOLLQhTYpt1hpZ4Tb3U0dVk6PFD
WKDmYR/LSWvw+vSaos0EkBfXXtxdf6K3sD2/O6+/IyBgxQJM9zVewmixgPZg+Nsk97vIfdzmWYt8
r0N8HfQtuSOsA3JCHoX55G3GSG/RFsYv3X01TSORLQPlllhn8VuDRIu56vQTGAujd6WADEbXe95y
JIkpCEl7Z0dpXHPshIwEs50p9980BOm1DRLdsV8IQGk4voNIouf18aCdRQ/PsEvqbobLyFgtAQO/
Sg6GjpVFxP9WCxrKhhi6YVTmAPd2mIik1pn0F/l1dbXSGpS89jW4tpa0qTqFjYWHq4J6vks5VfT5
y1svS2W+a4kXri8m71qH0gKLwqW5KNx9WqnQLQZDeqNRtpfxiS2z+oi7yt/9rBfJY9mCxVemgsZL
3IoDSc7SGcvzUiaAS2kXeEewsUDpoM4StbMJH22rzj4YJoupaGPSWKO5ik3yk8A9LOQUVp+0PH/A
ltL69AeMumWisToN+NuaLT3WoJQEPCmCVifz+X129cWArnSF/kixt9xe2WUiCnHOBAlXGtdYbUUM
RLd/XLX3yWsAhlrWizf2HiGUoz5MObUpop1yTbpPVaZQJHP8JeGc7kdyyCisP1xQiNp8Wsmh3MzO
185BR2JanQOXni1LiHtamtMK5Kmmg8KlgSncwoK0/3vmodxQcHqQfrVazsiOwWv3ce0YccUQi/XU
6QZsHWZWs45pcQsbbc1zUcasUMltGfmVtKCegQx8Ibu+t1oCogErtcyj7kVu+/i8gY1/73LxVfTu
LVVEP1OUKbJDJ17WkHIzPbrpPjCcBMzdx6WOCltAkdcVlauktxa9asa6cMgNfgd0UxdeEUgs167r
d/zaHbKX5KEl035L8mOjGNM3hDv6lxwJLWntH8Qwj1tIl8xht185m+JbCK4bj7zoOqn3f51wjH0A
w/wb986yH9c7ebooMP7Rc3XQm6eWWzSB8SeMaK8dvgS/3cv79tstkGN0Vf2m92CpK6sW0T90Y0lo
2UZMP+IckuffWTv64k2QfzVcO8vvCHvGsbo6Z9I1JkjwoARiKD6D3z4RicIuZP1hapodoTGUf8Fb
KCNccwdr+Br5TiWTUCq3QTFkF2RJD4MfjBa5baOOwNp7n5w8IzyUVt7JKVG8/NFo0iflzcb4oqrM
38S77zUJQIw/EPN0mmyUX9SaQyZjsINPMFUnm0NG3ZtcT9Ez5VSe2OfJgo5zOT2PUVtWkYKlP2jM
BVHORNb70ZdL4b+ONk8xsn5Z8RIQXmze8K9yHLSeVuMijojZKRk++oUSHft2uwAArX1XbB3YJln9
OFnauWBH4z0Jv6CAC3rOeJfBuCN6KTp/0Ryr9ABe5T6CiqdiO56WOaAoDlxodPN0KpT7O3wCrKGQ
7/cl5spp8R2uJdHl5oEzv2jfAfeSU/cV1PvbcIhHXboxlMTScnD7siWUCkDcvxFsXNlcdWnm0DEh
7a+rJsA9BaLHxx7oMG1kV8A6bltEBEhDV/rpm9Ch8sujtwZdosnNnPk1rI5RbSVLYTKrFzykwXq7
K9USJ6mgtIrw1SJSKuFHknMZaYF1f/mSDiLrJr/OQ6h4JgFqiaoCkYIy9lAjIrA8KfeirTNRSHe1
PWedlbCGwJCpwKO8dMQ44Wtr/Vyx8qM4cXL2qMSBmI/UbxbnB8SgFLbqjVhU8mfA10ImiU19ilOq
xITH/O6SCJB6EmDSYNDUtHMd/vTPIrNjgv1nXRMVJAxjndGu1Z1gTCGq76yFmjHvp3ulnJn7jZXM
At6pKKA35TLhrFPIWACi2USj7x9s/24c9WXRROqH+pJCUmeknLeviGu0vDBC3R8HP9g4pBRurr5J
tZzwHVJlT9eIHL9AKa6R9HyX9Yt7skvCyEvTxkhY995Zb4A7kOmDvVrrWIbZT6ecbVegVbTYj8hY
mAMqpOQqjmdB08rBKITqB+ywVPHqz8GKvrXqFU+GKkWHWcMSdI2lyORw2KM3QcofugtSuEP+Ntfc
pthvWMBrdKnZ7seSANJlf+obIGU49vxGhAJ2gFlzbBfvIUq67GjxBCk1XOxVAXxeBYw/PO50BaKq
GgotvTbPd7fKheoVmnYs5l3KiqeD677qpRyP7/B3T7jyFFsjge2DhqQSzcDTUXbYp8spQZbEwj45
DRv5FUj92eJRR/CXa/zUCVsS3XP9CV8LP3zjvejJyUfyMgGYdXCCt3BRmxFDM11zFHdBLgheNuDz
5mH5G8S0JEfyA9pzazBN2GsBnga9c2CpQMy11wZDwnE6tzQs1pTEWURQVBHktJ1b1U15dMvtmHvU
9SVwWmpT6t5hwZordE0L9DZ2GVTKS+fJRMBAXnyZfM5CyRPAnDXoJPcq7yXWeDRaMT+RdbqPsl7h
fJUZ334ngSf3hJMzoGvbu6ATpzYN4D3oAHUCcDohRdAUc5T9zRXYeEnDuCrJaNnc5mGC6cc+m9+o
Zp4QQs804U/LyVdsiPTeg0+zumGMD3FbGI25tyxvfWK9yQbjuiLKdi/iCdT86CXrBqWSF0xrJyu+
6ffeHPKd3HJOAPPtTsCcFbYYHhPL/mfAbxkpAt9HTXxemG/9ELISexg6eYUpJxfO2qhG3BcVsQWa
YgIfvexuW5T9fsRJ0yh9Ozj6TUg9dhGgoYHv2ZXpycK/x25OL/ZA4s8/tzzzwmbjsiNjEXhfhtTe
q0Vr/Xl7w0psyOSr7TPc5XAvF97Jcl08fpcjOoORDuZ32xRt1sB1CYdaHPKeG7fzkdU0J8G1qSaO
S8eDXHEaHuSRgmBsk7rnWwlRADHgzOSqL0a7JqJnPR/Kmnc82RymOSi+IPDBWTMKeFZYcb+HaUuI
NGvKxPn3a9XdwplIhlsORU1gLSSJ4wekFoXlNqvGaBXiNt7bLdnNqzGAqO6yM8oUBs4Rdp/hzyUN
xQLW0fkWuXjNo7bpzax3F4R7aweOtVTsgzAOu18d2Lk6fEUJbw8jUUM31y+vnCd7S7KEjW+WzV8V
yZH7GFcMGIxTxaMoQ3YEr5n93AL3qNNbUX4AqtJFnRztXJK6liG4YZEN9+FGiCI8hKrVPgmG78xg
LvG84eW9bl+jaOmEfxXqt4kbgS3v+Sr45wyeiayhZjH7nf1RhDjlMXh7C6czCr3rRAiWhEBWQ+0N
FEioffo8B9lwqIAsyQtbYGey7Ku1yWpOWfxMrqJtllrzmhKAdEsL0jw4ee2JijbPdCba4ZdHDv+R
oPZiG0mHfgqRWHfS68PR9ffJf4qvShgHHfJJbzJqz61N47MHj5R1O6H93Ini448k1lMBUM0KIULq
5jVvyHJKjckAlI38Oc7sJHjNktU3jOHrBKsrEVIxJf6q5EV8zezF2R//jMWDCzW6vTaCpitnfhQw
dHoB/mDI2D4jwVU+/LbxeipCO7xVi+jwhHbqnAt1BnY0L9CrhtFZO5gVxJFJ29Nqkt4Dqhde6qeO
CiQ4jJIHowV5Lo54wViJNMzVZ7EUl4iIwSBZoKVJQZXKAyDuglOpi/Ld6cnhQSitrZFhVYmnqyuW
cPdzzFqZlCKMuHtQL27nJWrvFa4Pv7T3lg0/eCAdsUCP03jzEzyMJnwnYLe5ClgCj65QcJXK+TlM
tnXFBRjY2KZi++bzE6SHfwBz8RSC4pwNo+0quPgNkChGUZDZ5oOloQDZ3FEtrVIH8L6DG+K7ozQ7
3RZ2GpuNkG5jB7nD1AJ8Tq2T04RsBkZYGOTpXD4ToLwLKMjeKFeX5dlLPm/XXF7EjFrEdI24j5jv
zAnS427vS4g5mcbTQl6Nym8ZAK/0FwFw3To0QTQg6FFvX73gSzTz9anJUXUCfaTSMkj+lu4doSRE
7/zQ6qeKZ+pVfnHN2pq9cshPepHFSIrE6igzpJ5kjwPpxTiV2ESaIu2/n+3gHTV906aehjh9tTHC
5SqdWf/jfVmxBkfmR5SbU5Ze40UTFO2thxlTlaU2yVe5/Pf1+mGHgJrVWA0rUOEDBUB0HLZS8JpX
QfphcGTJ9kPI+RRLJso4r6V03RnkNnbYKeotIHG1pCX+ewRhxWD2SURCrQ9Qpmp/yRLtKMZu7NEO
LdJgc54USNwltKLsEobpdscmtlpmPlsf6jnds8hUZpVQO2O2mr5zoTs+2HmXuLGkzqErFBlfTAV2
2Dm9uuga4v/40f3tk+cVA1WVbYgVcwjRwnp+lvBFhMGnLEGdNC3J9Kx/YWJyM/pk6PAwdbCJ6W3P
Zwi0B3cHTvv2p6gB8HdPf3QzV/G0Uca823YooLOaIz1Ac+aWu9X2dv68tY1fvWvxLxmUFdt5ccbp
W6xqcT1d7VcliXdRvKAOOh8RU5Y3GaItDWkZG4D/lLBr+GCdBiolRJtNbBWWkvFm9JsyCvBuvci7
ykvNctgs/heM0EyN+MbxMJaZuGcrpjmbv5KXuCN7QXsPUWlh0AvwXTNBvH2aU21/117U6H5gwQZx
gmKlY40RylhYOoyiaNIk0bVqr1+Y9Mh/WQVa6DTKRNC/10f0eQuGPAyvjodQefHNuKSCEXSqH2az
ftfhtxDSoQPcfmmJatUHaD+9UuTdifK94zkGTqCQTtMt+76a07YF8bGOoDIZfYxt6JNXpbZVNDVz
akCyrxazX/G1KDVyIYQhqk0WzeCwmzhHo2DgYgOdMNz4dzOoqACcDBUGueDjIGgot16VTjkRoljJ
lGi2AyOon/WGOXqpDI84bd/zhUJcXFTkB8xGAMy2k0XAKAxhdqmBFDCPmf8XrjaSawavp/6t74l6
ptK3Qep+JCYaeytR8BJD1twhsuIdhpFCRKJv5L1mO4tqrxKSby8TRRRzZu+rzaJmSYkiewm/3o31
41sZ8Gf+w49+ZoffXzq6LZrBHK3Ha05L1FIaOt9NGTlf75eaFuoyQBnQP4UjtZHbN9rTxazzzV8P
fKBDkBE50enrZHLCjY/Og+pfmBSUp38jFrxLSdY2/HW41MxGs/v3/6yXYLUvwARsWCR+PTdO6JIT
BPZv3up7sZl1O+BcQGIDsn1/fZ8aGfFGRkp9nudeNy8n2N6C7e3C1qwn5/gR10ukrLQfNSHUcy7P
FzQ8+j8+umYKlz0CXMVneUkbhOCNjjCbyEtyMlU70La/WxOwf6GM+rBKHejwUQvCMAII+zNwcwL8
z1gpeD79pGg8fFaNvf86shMO7Ub9TIylIoImkqIFhuBaEmTanAGb4UOsYLSx5D0pa6E9HcdU6kXj
9awy61mdHS0qVx71UY4FUAm/S9AJqLcxMNrQdRK42pSNtQx+WTmBudNGZrxhVuziACfLDI/h8+Gs
9ju1ZnSW3E6+7UYhxOWH4dfHHa41t/r7eGEflAhz3B+IHjb0bxw+1sZunJYL0ftOHVzoCNKgBvjB
3CIO4OhsDKUBq0fPAw9xYdrFtjGqxWCmNUweNlB0hFOzL2d5NF4t2tGnJRrEGtfpoc+hfN3HefsG
HPtIHiapB0nWZ+sOCdmzjLz1Y9WJhxRpnuHPV0gPN+JYApuyQumnbtZa8LgoY2U/mt8xTo23ery8
XRp70kAsDPyr46PnD/psml54fM2XaNiLREjRcu+EbxnbsVRAaRmcE5f2FMi5cijVtUrKV+Slwvdb
fLdXEK9gNS2BbL71KW5WGoAueVs3d55AywQSvLzJ9W9LJeWjnSMDyXfZIVPBJqC6YhYP7/O38SPW
Jo7YENYHvZrg+WhGl2qNLt/Z/0pkL31hNqV1ER5qM8vRFsEp/oPgJbaONRqmaYBRjqAEudAzTyHe
ZLL/bENVj6Fp5awYRvUitniXUesyD92HCmKSxCkQJ8lkGgFA4BUe90GHx3LoNqDTui0FRT7+SMMB
A6GNBW6rkVQu9Dt2+QbKKq8QpRmv/Qz4+9djocZJeaMtY4e8BknwvFn3WbHRt+AhieAtHB7VicwR
yNs8jwFWQcslNByQwFIZ1Nc9GFMkFG0MTw4/vGEs/NALdZaGXw5u1KGNb5WNuHmtrR5wVZIzxqVN
g6aV72IE8gqIlEV0fXuYH9AtLcV6ZSszd/fsIWyjcE0rYCOrjtozOEXWBBdnCjSt7erkyJZ+yuHa
rtJ0fibdI5STJ+SXyvllUr1C5ckIwSs9/dBg+JkVt85S9ceHZvwyM7YakRaDaC0riadmhsCunSTv
+ha4w6UMaZdvO8mFT/nERBdzEu/XQ83oVoBTLVxEyhH6Ubknn9ruEF0YG+0kGsV9lIJrROIuHDz7
271Kn5XxBRProxBWGKqN39F9mE4LIUgxQPdhm4MYzNDd4ygv4kGi9e1f2q4kYZhVF62YnwNj1ug7
qRQ/FAtmvM9WUfT7j1k7xLelfJbC0De079QvFLQORwzUbs11nNBIgO9U1NhsGf7ks8TbA5rpmVEw
gEGq24L8XhM3obwhJBnAGGjVuJH3TH8udYGEwSw2CQW9ntQT396DWJSAPwUwlcy6alM4lwki+CiU
VmzW5oahQhL/pYDg70tknLpw5uJPlcJLstRmDYvBKiDNgCTatNzOFbF7gMUHaC7jVYZJdLncWglE
xSfGcJkdiG+D+KqSq1XaIbqiCTd2mfh32wx9JC76w2MsjsoaX2caf/jF9MhExSZsxWZ630YkHr8o
++qZ99O6wF9fZSWAh+ODXvbK3lfUDe0w6uULN6g2JQUGPTph6Xdkpqdnja/4d8HaYU5qEQPavVlq
7x0WilZ4RoBwjsuvGfIoHQyT2zvW4LzEd96eTwyxeWjefHgangGc0rb8GnFNxFaYRxnqsI+8M4UL
QImqT//chM/NHKK5VH6+ugZp64MKBv853wlJN3HHlFGWPDzBLgB8GkZe+qAXDclqkKQhQRXYzZG5
sTtHHVbCyr4H4vuevuXpmr8Wwt80xsZoiOvw3vl+fwsnU+lCSl+Sv7vaTD2a965KEiKb9ypEynO+
M0N4q4G3c/wIF/3ghbsGhtNerfpnM39PNZLS9Pwiux4WMBimiygkS7oAu31cCzXr/FP4SeMKBAEw
rO2fiCxXDJwePIQ/ujxXoicFHV2JRt2EUWPLCES9F/nIBgWiobARRIFZQ9XwlOUvb2dfE91IwiIL
T1mMbikWFHEcp0QizFIiZELIbt5dN1cqgzYcsEua9thY7bWDOtyIW6GXrBoAHaq/mrbXyAppjdmS
K3+SbXbAitqDUmM2jNasFvs+0lvBeC0DQ4IY90mKaRfCqu/ciudyjRyncZ6qWzF8ITtjveq5zrBR
rBLFJLv0mm4f11PxoNfYQsyAeKhvtM52fcNoCJKcrHN7IpM41M0RA5Mi11E199C0DFKw88Y5j6wP
VAtR0mzknUsxuDq4DSzs+Ael0I/LmHefMfNro0kVw9H2MVaqmuK6qwTUzxcGp4cFkkSeSz/JEgyE
hooAMMmtxZEtcn4a5f6UWXpPSiM4qb1UsFNrFTdQFPAmM6G+t+D009wpMrT/0mTGMLcWz2BTU7ZU
et9ohWe9aouTZnnDACB8AX1KiD9PmBuJmEF0dle4xKFO7DYQYlrwkY6BFOoyddzVdEPlXqGCrDzd
JIhFKHUxPmHDLGDM0y5FnOGkWorv55ZwXg5aprkpVUnLJxLl2HXGJNmTb/oI/hVDIU5W0q05fR/f
rLb7xW7dTPlq2OBjO9zHfrwYK7KNHM7m2/31nT08TslAMukj48MKx+tN8H5cfYMpswVRp47N2rBa
04K0O5wqQqipOr3PaaoI7WuDZfSs2bUslIddYqAe/7/YVhA+CXrDZdov/GdliGKB9KAqBkF6JXMx
h4ZOBJnggCOQsW+kRqzbR/tlSGYyNfqRseQryvNxVW2y+fAfyblUF0eOXN3cIhLhPX4lO6YjrDxB
o4Tf0Q7OfCjKQmxiRalnacauMtPWcmm195lrsRcRUuU2uSF2tp0gtiaWFh3eodjpALWf7vxx5ZJ4
s2IJlDeiFLqtQITD5xls0z6bpw4eOEMg+vtiMWj+dwpNx1l4IWOpFDgdvvnTmbjQbK2mQ1nIg52G
dEbHnfIrq6p+ZomDcC/uTULSA4VCuQ7XrbdRhnSFeCZlEmCHy56KrUICr4BBL0vRD0qnehUPrM9C
u9KDHCBLz4ses6WXIrsfz32ab2R/fgx03AbqK2PoHMMp2wtQ3tRh68I2rFADbFXXKCeeI1ZMihbM
Ie2Z+02SLKOcr/yTDaA5jazSJYcLkpvCVPa3ps9fCaYsq6YN8TNLywDghnPz2jvXXnSwei/o2DEs
dUzkVnEhNcUO5ZqUg3MlmBcH0WVQNnO378SrZV+gpCIqUd/6ghQxEgbk2UkSE9IgjmkDPvlMTkC8
bMaWQekGGi5+vOmvwOTTU07yH1tmT50f9ikkP6bqKdMTNa2YZA3jXY9CcNqzZueNyl3rBBlKoI9u
Vv2wNVV5Nn18hbhWdGXQ//f4eW9+/CncuqFpvIuaFSg6gCcxXeETSk4YZp1uaNleZ9+Jhb/gfEob
MAkxNUSqyhnu8MOio/WZbeGCNDFPCu5VU85NnueB5K1O0dccMIfASmwQmLykkd1M10K+t5dc4Cde
aDsxNEy+7nbj2+GPGeLExKEMFwM8nHhb8c2RDuQLBRh3TF8p55YtyvCBYXRsafDB9fjFQEW9dub3
KtjxWDeNub2LHqKX9Re7oGc88/o4Ty3IADm45KILnAruVtWqh7Bfb9c8tyxr1V9ulU97iiiU0vRK
Sy8ErS9qN5gFSEGCcLUx//XglCm7t79kWWVA1Xyi9aAPIP/CVDXmNPBqt+KDEmbwcojSNwmbKpcM
sDfJSwbJS8Yf7RtKGDcA/rzQYENN7mz2gtonmih+bTlD4xNti1Bb9Eptr3tMj48JwWg88EPIxC5E
jLfwnve4M0c3Rix7wxOJtGFDZ7jGnp4cLXyL/bmSMyNd81IANNFCgNn/NkGJ6tSQJpuuW9I/tj6J
ax+NsaY4sEadWDICFlXLfy36l1sNMN/AEXG2cvL6r6U4mSz5XRiNg0RVyqFHKjf+f+DwXQ6cRUVJ
NH1nYZXOvN43KfPqWZDJDR5xUFYro8kn4XihcBgOCLFZ1BGWoT6YqDyTLV78aedO9cQUDQE9kjB6
Y8Ntn0XfcJt7fSSniAHsL9lRYBhjjGvnr1XbjN1oHn1ZfGdL3djpATo29NsLeEifkla7LB94Pirc
ILUdjbtB9AJeFqWObpkNY5q4wywqQakOjgtshH2cjMFDtoSU1ExRsBHTgGmEy6vaeBmQlzGFgZjE
nBwMtTUrVh3NxJtXA8E+VB9aQiJHXx3hC3fkERbubWNsBHNdgplYS5+UdTuNycUn3Kfqf3noOqB5
efn8K4xX2bhHPV7Wm/OWHFZRxV1cfgJoe50mCf3iGy7KIvfVoQXWT4dOdBLczsrVGfDcTGl0T6xO
HjKHCo5FjWtywbXEFxxzUROxOiJUo6jo0IrTDRLkKQ9s+bSpASobG29sWQVos4+lvilHEcLHD3wc
5T0LoiQN/PRZoHApnbvoXep+BSma0RMBOfmmDLNK5PZvWS0l/Q7briPokuY88OrqcevQqcmYVBzB
uNPRYP92nH2wTDdrFqq5IOA0emfIPdik+d/e/mTCFJl0XTfInXNYXnSJCH3Geh9kIcEUJ0iawN6R
mD3BLXVxUDH0OGTU4SW0lNdIUYpYO3rkNnsFZc7IYYJEOxj6w58Y3bLFmJ1/mu4+R7HWDydNuZ0X
j/P9J0GcZrHRKp6NHAeidKxrmfL3EY/iD3RQyXx0XhkaNhqfaLkhhR5i8D1jj+QJfLH2XUfNJDC+
JZdWP2mTl3RYh20DtgYq3cz4sQnn/ATchPWVOPqT/6tF7VZzgvV6DYxmaguJ/bitJFC/HP4gRyrs
BrKWWFAwvGQnczHpAEsJNbZir2t3fDl10K8cvceVrlFaOOhJ2ltk+EJmEyP3cfMB4G08PIZUl5sm
w30PNihSNct4YW/uhW+pKT39oFYMcUW6XtiHuNhHijX/DL1EJWWl9+Y72clL8dEO2bUSIm0wAuF5
3Q8wb25vGKg+Tz/aXDgJuE/6jHc/denaV8PF1GC+LXQ430zvQJgdlriav0k9QWO5SozsMeeE1Boe
nUrM2baHJ7bJT4BiwpAKVKVYghOSnit9L/gIfOzHELY+1ycPR44xZOVbCCLrrGvHlRJmLzIL/FfX
tAcbxDK59fHc7XNP1l3zKXewUpgK4L0FluETIKDagQNvImcaXUeoc7EHIoZh4M9IA94HcjXtTwEH
IW8cG1kOSBU68L97w9m8NdiJE3rJPLT2x3cmZO/GAo/SFDUN6D+7btQW75659AYT2gpPxd7b4BVw
IBXijXExyovpfHcFsSs/mRM0Z0S1/o8uMMAD6Yt8jlawa49w5HGa5tqqIZZ6xBbmHPW7Mt6Wugw8
N8vrDHcrNpy5eoPRoXVr1HrhO9oLs1UJZPJS95PrMUjKf7qzTKuPksXycFEZ9KrtFazzavbKqWWl
H0Y71Cz78h1PbQZ/VcTo7hGQ4WbbPArDGHpDuvJ0dfH2Zlv2mbJfZBQGMLJcJ4TG6fdvYYL9YHjP
sMJWHV3gri5dogfNAzyZUmtoTpAmx8seBiNZ7MToNCkrkuCu4aqMhLzqC2xn0ORfc1p+kH64aKER
SR+vSVBsM4vqo35aic7Z9q9ejRybYfUvCJRghSr52A6ZTkuv8buKtDITuXCHp/zoPSK6ScEcM5h6
BJp5fVxGs5Xa7xlhEdBQfn5PENXnEBEW9f/Zi1APGyndEPt56GhpsJs18nDCPRpHWmtZHYC7BuIr
yRkBalMYs+0iRT2AvWsm5Z0WmzqqXtT349OYkF3q07RvlSBSIrMLnd8uBZVoeTZmBJWAM7hn7yxc
OVbfr2KdGtdBEXf5nrlQvKbEbvQlGwatDN6d8mvgwpsFQoRQWR9fsjy5VyP7LuQrYhvn/Or0P2W4
nlF1nGlGGSGDjuYJdjJA3lTav/2eCKVYZwGlz3aIE/7ljAI7f56ynI/Duw7mbyt4IhxtceoVAMal
0TQ8vKLpLuuKaC4498GSiPS+bZBuc2QoheQdbKch1pWOXIBTwi4bfKMr1gw1Bjr0Ell6LHBrzLta
GMJ5LxQSldKEUM8hXJnL1SCIPH3tdaPfebrqqvfALPKI0f/EP6iibE33XLgFT9KT8MZxRiC4+oMr
vnpKJ+BH1GCwi9map1MjWbfHq4tdn99Kv5oMa8wOFqZf8G1rx+/JeNyhtq8/CTe8enNTFOZvuY4n
PEjMVNeRbi6fnKqVairMbo/0oKaByBO4w3JI6jD7ELbMb5btInewHn/oAS1YC2Xpa97400mNDd5K
D+94Ux95gg/wOW8aMLbZdloKHJ9Za7M4t8Jsa+JeluhtCMWzuNEpw2q+QYmK4+In5GtU9ZoFi2TD
+ihhusHVZzd7BcyqO5QcTCUw3oJtcamZuHolbY8+ucYzPhSHDj670vAkjsvaanq7v5/Onbg/kvki
iLyOvWkYHysDdKfvUhbFGN/VcPPfp2aVpWM4Cfb1PDq4tVt6WjZPdFmDpHcTv5MLNQl9ttrwikK1
Szfvbbz5cJbIGOAm7mpS57P2oC2OcsHa5Ycv+JjoUtaedk8yUvkAtVNVcZx+pu/2+Mzf6RwH1vPM
p7ubRvYDccmfaImfD7yXKKBDX+kEEbSh7qt+lem+WAL838YyTWD95UMAn++z3Y6lSwIjyEj4HYSf
um8iXcegOixLbYdxqcQc9BWyM6EvI3tMn3/iqSewWAm2PJQikmXgY8scFVjsY1Qrw5l1ItdJnaVv
DtmGszTUJomOBccntCnSHm2pu3xWy/SYNmyXKuv+wClx4eIoHHdtcBYzch7W7i338QnEGZr9v23q
NMZhEVUe3ewBTuODmUDRNVjYFpI6ODBblgBxIT/XmLjt5YH/pqpfh8Y/YU7jFv8WnE/2mNlC4VGJ
GbQObEwcBwUN9HRSV2uMQ+OkcdchKT+GLGy72wduqm3aRAUGqSa+NHzCgCzsDX5ljcAittp3wvvv
S4X11Djzt65NWIMvQ6RUGELAh9w/IVBrhjts12rsIipmI+xlI8zenljh8il9AW77vhPA/+lGScGw
C17+JZ2K5aWB3BjKU17dLrsaq/flHG3+KCUEnisKm37ShwGQ16i7XXZGIFso/JFKiHuExRO2dm54
WyzsM5RkrrAjZcCYs4fZAkGx24KuLoKJq+C7UWFEbiyTgeaVFgImOlOcmClLETX/L3FAtQ+r2S+N
AkR0sIIamD4CUBJK1IqGft1zEEw2wfEL6KcAmhWuTEHmsIbcXOu56cqwRw1gnzxJ8/NbNTvqId7C
fSknbFkP6oCk31eFve4HDpMFoX28HEptlc5w+WH1NEQBbouCYeM+PuQfkPOgggOwmTrHlSWEqAWZ
SubQF/l32RbQTfiC9mzkJ6bMYDXjxXy7p+30VWrD7Zx6kkx3cG49uQh32ycp+tHJuQPV0C1/AYIJ
Cb+LfC2H80v3HiEi+L6XreFCas9Ud4bh8JoWry7nuRfmV2g/iCHFcUbY4ixO3oYBWZHRn8C8N3R4
5ReOOgsZqQSLYbScmhrmk/ZhtYurUV8siofjYKu2w4fIefM1c0uj2LneCyEUUVAnhxMaAZpy701A
2yL+4B8qFRF5xZVPJ8bRNBXOoLuGSW8f018X6bxu0+SZ2rm91lniA6FHvRTESeF4sCuNaTBWcaaO
lsFkAjPYj21IpsGGkA2JzqvO/gJiqs6FoX8BFbnACNkZTQ11rfM9JPey2tHN8UvTiadQSGXd8iCG
134FGX2cOBVXhk5sVUWiZX9K6nDSxroGO1x8kngyfJSJYTVBeFzAk/yyazfGiR/ko9syU5GuySjy
A5kFK6V1F3qpPf2O7ahPr77E68AsK/EbgHlVS2YvjxhkOtRcjaniLxhg+I840YyQarl+ibik1Tq/
rDYZKqSx963OZx5YAVHqQxkavqt5Uagqm9T+X9jGaKDCfrtIl5rxEwXEvwYD8wOUv41HDOaPb+Ca
eKA8e5whlyK1GaUx4moWoYWHkYMvhzhMm56jOdA0BtAvQ1UT61+wnntO9ivIuV8i4NTzNYMZc9dD
oMOAd8HA+wjgCMSMHwI0m8lrUlSQ+oxoSNsEIFTrIpDcKGLUAOfFyZJlAUtUVSar600wWLnBEEm6
uFcdQ5dzCwI7MzMTj+ibTrNXAdiGb9oJDbD/wL8qK5DB67HV570h4RiLgDy/HWQkD1/6SaRG7EC6
loA7YWZDskfCzEwlrZlSxFCWtCs04eeyIxkBIeRf6T1+b9VQBXCwHnn8FhenoSXIOWjvoS+crjXQ
RNUQYYYpQXEfF/DHbDp2HWEiVaZHXywD83UZUPsfMxQsYlHa/iMsgWrmxtSfEM4Z2UZpkXdWRMKo
ACNnZo7YXbvKtOMXv6lZMKoeexl6O50AxwicbKC+qGVp+Dp8sUuraKzXdozphK7alCz4CYfMxx7F
SRNIjv2nZWJtc3tAc1qCAke/aSFP+sgXY2gTeYH/g4FnIM7mxwcShKQxJX2gyF0337wsRs4A1Bkt
b0CnYxeCic9+tCX2QSSftNexeIgBXHwR2hvI4RlvSip27uT/8Zc0u2nnaS3FWJeLKJfGDI2vXW2x
/QY5TIUWuKSHSMViXiPMUColn9yUNfQwBNSEMR6Fbk31jqziIOMogWzqA/rkkEGGo0bJml7wu81Y
2am4yHPakITABUlQdpmCDrkzTU/WOe+RWN9xtk6ZnQruRa/PCD+GPMruLkotLzrfmeFH75BMJbn+
nuR/JF8YujqsAqbjs0qca6SkElyLViE/jYwqNMyz/g3cjrNyrxJ0f2uIG6+kzePTjK1uvz5s6sK9
9hXQnbCJrAsql7ZF7MhxyWgNdNtQ/swYDI6mBT6BhbNd97pAOGlxJlOvBFbBvdgpkjYY5MWxDN2t
4DgwZVUei5nl6UW6PSi38Zoslcd/ClZV8+OGCfdunjIrWDeOpa3uGS1hNDNzurw+7TYi3st2JRsc
DTctVx8aP8XNygiQjFVFagptEK11a1c4IxIzNJH1YmSUN9+cvhcZYuEWPIPFufXpKE6SFgs+Ldr4
n9JQ7pxpAYXvJHk/aE9v0dmlVRbT+jD8VV50VjglwboXV02bdt1xsXCknzlPjvbXHNtgtY2+Byiy
dWFe1NaHEPLqOTeDbXh74gX0hp7p3oLIJ6B2sIp20F3+9bZJSlX6sJxnLDVFIumlVaGFJIS42yoT
/HgZDLmvUL2XaEZacmc5lE/EBBpQ7eET8FhXm81H8bieDq2e1u/sOq05QOuh/4h6e/MNUeAfTRsx
86Wu6FwHlC3ykoEXbtx2BRQFq9tUaQZFmKjo5steeVKqYBuPXkQYCo2GLnKPlFgVWSqeO5q2p/t8
MgxuCDFtzEWX7rcGqvfddDttZOn7eHBWMSjv/kbPwFHzh0eF3OPa6lO077ZluJr5LCFy5HDc40pn
75fdIUiH8umufSMTcDWpm7jIZvj6Gjw30ADz1gPDyKFXjgRdlhGLZZp61rkSTk7bn2A9y8s3ycqu
NhwevLt+G5KDv/eN59NrNKxs5a6DAVsqBD/hbKkzl180BPSpK5O8QHo3QbIW9dMzu24J5Cm8ypRh
5UgQflDeQo8J91PghxKHhyu4eoXiYHfISCKmWSZ4jnpYIJWmHbNUBKoObh4m9wPKM7QYgvYgoX+k
0Zv+gztAlX2uZIP0TXNz3W0lmqZ2GUY9V165QKDQqs+EAP8QHOc5gXXOKPiWmVGMEda4VBXSTQd0
59LLOhchsE7fxZViAYJmC+8snkG0M4QeQKlMRqJF0gdGf5Iy75JdfMSS6Yk5I2Bfu5Lk7mZngBQa
syvWidPK7xQMduU1FiYWLjaGJGRvCrma3FSuhN9lWg5OLBjGLMbaf/fwhoAXO3Z8iEpjSH3A9fT2
nesfOgKz5GuaVQoKPAXzOarDvD+qX/TOYF+Nz9GfI1NvtjkQYbwT7Ir7ftAy8fhGhgzqD+OhPFei
5ymVKWRUuL2HaqFRIVgX4IGNGDXopcHwLmVLexPxlPCS32UZ4PN9g8AIElprulnfxDhdEnWyzpsw
KcPpRkCajUVcD9tLYH46kQnbd12yazS0A+F+5ZAOCRoaJ+exPrxktDKD0DVtP4VzC9tSFJW3GAmh
mufsTC70E+eTCpxsObq+dtCtjGBcQdh2f19dBCr5jc31tIzD8EiMVsqmbI6l8pq7mzMyMVlH+v+C
ulLAHpF5VUIdFFLUu0Y+ZlWKP1n6CZGwKc8LXOIsYgFaiWlJt5bTCvGPdwpqUc9sYGZgnBeMy1DY
At1AZa7Zc5UFIk2lXje34T7HV2q0R/oCZIF72Zek4YVPqKWQX6+eqZj3KuBz0mHRlbMEOk7UXjbm
fRPZzKG5dWOv307+84TbKBcUXK5Ix4LUfNmc+pjyGlKRRkh+T6uJf5eaBIzyUQ37Dx0L75El75VR
aR3QK4StseGA7va9Xr8igYnLOvexpQlb5cAI+H7DVKnCMu9B8itgEP9C+FbIChpE/sz01624EYRe
76NRwy9M80e+3a42PAkzyXvRdc0Ykr7AtzPo5ih1Sgf7ubrWuPhfSdg/SQ5BntL8cc6rEHq0Uwur
jJ4fHkgWGIFIvIIHWyCE6s3STvV+dCFNbbr/sD7LqW0EKRjjH8d3LKMovyFB+FoGJltNkCGudvnd
XMYzKLqAYCDBC/LkXV+06opOGJ0MG9LVSTaE2bRHKqUeavUeCZhCYhSNypS+IxNvi7AfjDpnmbDh
B/h4kHvNc2vxFIp/r957vbBFwsTxIMMP5pMty/eCwkHpiaYO3pGKRfoL5GEindfaczw4z9uPpFsf
rQPOTJcb8O9pZxlxbDaKyTjwD/jAcmD3DjpFtc89o7FqIJ0rduFc57809KcDRIQmIA+yPmx/iEeR
G5ZAlnSWNp/HRljJBW75rhU7OLjRzVxAszzI4DadgsgTjrG9anYTMoEBLSJYMsC7Pcy6WJscALZE
A6peEgceWFsrHdS5pBsNxujvva/hruNeA8y8ij/iU8fPDkMrlSLyNgH6YbkIMys5SwGws/tujJNU
My6mbJIPE51YZorMd0x2VLv2jKR13umtUkWiuTQowQiZX3vl6uEQL1zAoLETGwL4n6ZWrHBUKqF6
y3v2+W4d2styvenIUwcdricLVixxXWTpAiQbTmcAcIQi89CK9bfsBForwuJZIegjPSkIMlYsIc1R
5rXqtrt98ePSZreveJSGiHEC8jScPzBJ2XX/1l0rDJkYDpyJmXJFd+HMmF2z6zRym1RYGlHVtiNj
VYjGN1hs11b7D+a3v4+pQyubAJXDQslW+XXSTF0e1JMf65osz9+sVrlCU/RkQlkkYQqzvCOW50cp
D5LIRhmxAP8laXTU7CxpcU00k1qjr0yW9QhaibE9cC5vQejtuTQLcwBapS7Le/NWC4UijublrxDs
OaEtpzBx08Ws5lWd3sxUPxHkEwJT+G2Z3c6zfSUcmzg3mi6rNRKCdY2CAkwwzWPaACFXdrzK9U+p
xloEZ+raWA5tk6ZTaIJbS8Url2q6hfrwlKprPfid6OvCHsbS0dxyWtYi1IQHuW5c1cPQgYyh9XmV
/94H2p1vOUcCaRkMa1SNGQgEV+RUGCJprlPBy5+txEn5yWnwgUH7oi2bkyM7LB72wCLdjezV+Jb0
Ks2qz5890Ph9iWOHupnJdg7b5Zw61r9AZ7Cfusgvd9Lw/SxqnoZRdEVL4zsle0kQ8xiCkoiJPuyF
wLQWC5dweiwsdKa2m51ZdLlKmYKjZnS4BvQ+gGr98iWr2bQxIm1J1hPgteDSDp7WxoBiQ3F438qw
heCuCMhqND85DhIrQudMnn7RUP/9+K5MVHQFGYOrRmlWi1w6m/FqRmT01B/icjddaTxpsy9nsTLb
TB2CWlgDRn0pVuKuoXNU8OCyPz01sAGKIpySrLDGsMqaQ/OSaxlBMPE/45c/ng5ebjtV+PdNe6WM
EYSfj9lq3fxiBwPQHAPxdoWTiCmTTHyWuXwdxUM+k2+qzTjXBujreFv0hXdTNdEiQ+zZ4bYdcVMq
HISoEGZyewHEn9fKfB8DOzsWj5X5D5oV3VFhTlcFZPaRUB7tUIxoXVuLl7Zjq1lTPuukmRs714wB
EHVzRCIZ8Uz294EpuYx+4GSw/VjMrNtE3+P9xlh7croXKVlHjimrllIMb8A8hu4K4cfaFWUVBcPx
StoOpFEY7Vbv80/7xMV6gD6/0EXS+SQxO6PrZqZZOqjTLacY3krdtgYP1zeBMJ4X2HXG5/58ZicN
kJUJD94caydeXC1nO0IMfSklOjc18SjZObR1jTLJKDZ+1UeEHDXn5nmMTq15N0V2P5Rx+38TF9I5
A7kdzz3eOdUpX4ulKhAKPERBrycr5ix6/jdHIvyRN6fZ3bMKcpJPPnxtYJ0RgfqLD5rFZxfWo7Uw
wymKEDyqotaAgfY0XeQyVU0MA8D+R5a9I/yAu0jjqXY9VEtEae7RNmDBJT2W8Iuh6g5bxIL4x89C
KQcNeUqVzJ1Y6xffXPlk+lrvYEU1x+Bpg45mrOYUCJccONcWfCNjE3/NiFDXDsHHOu/8DIDgizUd
jUIAAVO7Jr/4rsOIZHTGbxAvWvpg6BFthCYTnxZrvrtjK8xJ9OdBfVQD9NwAI3hr06uqgZD8bScJ
CCdCNODmjspgXwrmbWd7pLgns8y4YMAgMc96xnRu/V98fIaoXJDtwD47mNXnIlwqUQKg8wure1Zs
BunKGz/FU38rNpgxPn6nBj0H2y+JnlUVhFu3JWQ/Xm7WurxEcKSe9j+gWEL4aiWTmQp/L9LyN0Vd
71LA6zgxdBVtElRChyNLwYad5clEsBRAN5ADVskwuZEI6Gk2bCsU2uvRQFvRjYpwEjZyldZMH4MW
oih7lmdvC9pds7PVqYKKMEFGP3d9V7PMiGzMrUmFz2ZcnwzISFhnLI6+U6tBz+lMqkwJv6VaIvz+
qDJJnx9mybKUCJhJ9QJsc+QDyGXcm8j5vY6fC1ka4CDsbg4LaZFsEv+Nh3rDmroOb/SMi9bpJdFQ
Awpytwgpn+4YbufNC3CAJo1RL/tmJVz/wkaYxFffvWIF0IxJsas/VHsg3VZ52eRPbkKXoKBAemRR
evyCsiMyEwvBNcSS5Sh6Q2ER0WnXJLhWSWyxXlD/agSb3wvQ+D60uzPZ3e8UkInoyAUhQ7m78uy6
uZ0xvaQ0PAecTyPP5aFWJP48ZZsxtEsapQwH3jFelew7XAQ6qfyro0+FM+ijxJn/KJI2aFwpxS93
2lILAMEIOXqNg6hMRmeMKAiJ6CjzMyViCs3F4Uf79n3RtKrE85JBqTyTVWkifuP7FltPbJ7SdQfm
EDa3LjPje/2tAs5dWSOOVW4weFJ+Nb7siaE4CVGsXSow/35g7KN/wRySKaYRkb35KPv4OsV+QDAp
aRR+X/60iBol21WBNILM5eezRsC8S89fZi+ZLaJsxGhtVeXNurl++Ecn2yae5aoKQtLwnFj89Ba/
kXOEcotDp3eMGgQ1ROeGWjE/9HVuTNnNYS+gJq0cUp3LAtgqGv1NMMU3GSqbIgmjT9QAEYlgSvUc
xDp+zg8m8Wz/ayjcMj2JSZeZI6djTFxVSuDgYjAfYdDg8QyoEp4JSeZOKlj7YZU7WlaFvpHjvEWO
4AcWMv5xVX7cFpls/Su7ZXQrdLqjZE7+UwdRHvNPAfWaBzo2XxxiACL89qKHS64qtFqnqWQ/h1EA
z2YFPAvBv7tbVDyI1wp7rUw3TNoZeyhfet4LAX64gC2ZZnSFOx2q37Cx4uGieFluekvb2Q5Haksv
09Vr5o/Jzi7RmmMu6tPxCtfOrIQxKGoal5ITGv5X4uTVEYbgOg6A1Xawu6erUP70UzrEfSzoiLnN
0u85TkeNP5d+acigqnyOQA37BBfsFrONQJdG2/bm6lPwLdMRReNLylliimd3xbbHtlsjNNBOGHBa
glSeGV+h2ZVjDBnoowTgKpginMAVjNioHEW39HBgCGqQIL7ijokl+qPXgNjMYVCjImY+Qi5ZK3tn
LRCX56VrTFZ23LRj8UWRrxwXe+plD9UxStqq/tbm87J2z8J2C50IEmJRmHX01pkzntKcttIzy6Dh
65iM8MwV5l8EQ/FH/zLFOOI2n/IPwU6MA5EQmH3J44QTT/dgj3S1LUiKzE0sRkHQVL748ObUykjx
ZBH0M7VCxZSTlhK4SzaaPkP804FXCNqPgLEYOjshhTLhKkeFsQOx5ccMDOlXaJKzH7LAWHXxG+lv
hwGBodg080UkrmeK5MEy9ckHbhhw6YTw1+9IpXSoiqWd5fXVlpOnVgb8H7VMd33eqbn86Zubrjsz
8H/fgZOjQWLAK2VdrpTI3LaWf+Dret3IpIQao2cN7Gl40SqQDEQGDiAnZoxeQ/bqNTGivmZ+ARzC
shOdkabLW/0mkmJYkKVu34UyIsW7+u66LzAj52XcC07KDRCuM3fx4l3mg2GLtKzwLOupgrXWH+Rq
aeqtpB9t0vNwroJJjpxA5pwDlkNTqeJzvD/YRvHHFFb3R14nm+xw2qcIH2vJZOc/VYBkXR7IghMG
4XOLXi5E8eGAuAWA0xPT7zOsVWWXqddq9xeRBk5mLwoYoPgrJd3qsIAE9XLk4N08O4XmSpLY51d6
sjQCoSE6w92RmeXp/ljqIjEMC05kVDVhCvKf8LQgEE6w4ZgF7EqLOE5UQYFa1FR6AL/ZR+3p1Sl9
UUPiDU4wEtSGnE5Qsv4oSXBaG0rCYpckmeczVCRTemU+QMcY5ppL7so1Yt5KjrhNt+fgfTNi62t4
8gH4g5h5i/hbXiH5faFARy70WrpY4w2wRDOdoVok2jGQ27/yKdg4DM0b4eQlVWhisNajHwiRu9to
THktjD1iJGGjtMVP6DQH5mVTxGgvBEY/QvFlHesdgBZByObqjsNYuTBjsfOVVxNejN2sKoOQcq0m
dMSfxyHPGIq83D8N00FqcpzNj2Vc/LqfsYLIRdEUp07If7rozV/4/LCsCqLmreDlbxvaypB5FC0m
9g/XQktt7Nve1Cpn7RQgwRkS1IdMvVuLfFIH9OzimSGNEgu1o+xMgRXFuyUPqAihwkDigDO/BhMv
RHCZMjEFenVd83voJUrvFPWxUIOTXD7qliVmgODzGfAgej9q5rkBmq2ztEKBgme5oaip0v7DVn8R
SHsnK4hN03xSO+nnEf42ZBsovIEKUh9PyxCs2oXKXv4b3lwsWIbMeba02tRX8fBcxjSKjL4b/cI2
rZFbygyq255uKrtiMD4U/xzMl6GZasWEZhNFg2E7FAHvjqoaHyQTfCeXh/2mtS7T9ARDGhxMI4ZH
/6BOR1/v/qBHhMfF1iljfuJFflIAfVn0ohlZY38Vt7KRvptzdQyVa6a+R8zLUmol2ijvOsR0mNug
cx9G622YQHPlWSz0+g7/jFY2fTRlTvadOilCrKHVWTPmJ31QTMb7WC0wXdKKGQI8SjBraSlNWpF4
/v2vFYoDn7TO0RF4vnofTGbals6dD3dp+/l/puLGaEDGVGD2LiJ67VgSy/eEQ4aIFSlr4D+X/0hx
kEKhV+KO5F419eTPkL7tFuACjoNX+AkAudoG4JmSC0+dgLsT0NcuZs485rdcd0XUJ1vhSGxqfYxf
fJRq868Pz2gfk6qlnCc7rzlFWk+Cblfa70k/9nPh3Q9OFTtucoRzlYvh+Seq0C+OaSNGYlt7NY42
ke2B73/qrfXkEXPxjaUeQ2rUsokSQAPNhEaT0C/C547avrb8jT5mvM9Iqi70KK2HFpSm4vjISPfZ
oB5atiRe9smkImWjj76OJqY2dXWBirqyhDRtYzy+u2u68VdwYbkpCuWl3uOrKVmsDAqcS2BqpDu7
UX5ica4wwFHX3t1d7ciRtoacBsk3ANNV2eQ1ihihIxB4h08A7SvXC7gwIqZwRgndRvrlB16zAy0/
2jhjiOD3NnMDma1tqPqBwjxPmeMsaH+dcHeTQJuyE0SXxed9QQZivtpgUbPd+Q+I1IZ8z0nXDTfh
4KwSYbvGusCbMqCeCC/NYyUAmSxUoUD0AiAfSJqWj8U1lVxmSnThO+LUcbR7xIGGZ0rHl1XsP8m2
gMKz4r3rS1IVgdwckLIlgyn/136dTQqP3kYDGjP+2yRGI1RserDyi46SthSd5n88wqUwxum08fim
pTh7+B0z6/I9B3GdirYgkAO7g19Jb+VI7R5fDqM9t34nZBtQjlgqzaeJEGMJCoKRZjBrKGJxcSBO
C6p+FhL0Ohzx4+iyx8nm+p2E3iji+LWoiWX+gkPRY6jY2MvfpIuBfpxUCjkNc+mbCUhph4J/O5Fd
qVSaZWT+sRRQJ+6qhrIcWUqH3s7hiPYqwdww5EtzBerYaTRLjQdLRWeSkhTbzidjYtTTBpyEcyt6
WOrycHVERvc+ZAnHDs+8PmSDLctyQ2hkLdO+dRbnIGfFoZXVcXAjXSN1S8jDWPKQJ/mXiG5qDGgF
TUt8Dw8qDbD8o35Q+ocdKJYsdfh+UBqyA8A1jU74FGFBpxB3Qr/K32DxRDZODwCoLORdy8Ok3qzj
j8qXsV0aRibympjV2Clyt0kBEbgn7ys/HQUhEGyILDTh+dicHM69hxsZnQrPEPicYVTtt0dkQnqf
J03eWFNSR+FlaBsti9fb8HFO7mYg0o5wM4PI7w+Jy7PhQ1XWrLd9cM+iZn8IP2fymzJyOGq7Hx+V
yaZwt2Q9hcbsfvwfvbSfBd0ZV0G5X35sFLSREO173sOeBVHgs03ba/oe175RsUABwRea/iPrI0WQ
oO8mP0feXgPB8pGM22PaO2IrQL7faM5zmI8+H1PYpEsx4zaXrNdKbhGspMfMLhAp+R8bjvn5y3h6
9KXAVndhSGACyi9Qmq1PkRG275NQ3acS6QCrEGZzwsbqGpl7Xn8meLY7rEa0w/nzyijB3ZS95zYI
oRSvNQzO4SNvZeC1z0EAwCaX39AHkVEpJk00AFeYW2PGYU0/vBKHcx3eSroCliVVvwgCYFZ5WLBG
PPH9we9ows1CAe1rr+PhHGcNq2gy2+lIpWC3sdmcaQmkfx4CB0cBTRSvjAEwnMwIHsqQ4jBOC7vA
L/x8JdASDfU4CiX1r0NOnpiwfVWuIOy0L+eAH9TTFmI2Obff/9VP2s4CMVQW3DO6nMIX00KT8RcJ
HOfE71pQvdaUgffBLJsfIvXO4nfkikvrUPi5ld+/YVAKKvm7dRjjt3Bq//6bQwVXpCQbdBhRc+pk
qSePMCLwnRuHvqacmbvh/ndPwd9XYCwiCU3oWehzUCoiR50kO5CUAUfRsXN6ky8SmnT564rx85r7
ZQHb63v8BnEIHremDP00jEXxowrT9UCXH5Yq4cCt2RJiYHg6K9xxqLmduH4cS14XVqn6U6sg6sf7
tgc2oNCKrkqmXNbf/pdFDT0qh13xKxJMffoI6wn13ehthHld+LvFly1EntqxLrJYOOAgTBRcbQOA
XkV4ynHe3XYBLdIGRUjLVkwwpUFssG3Q+2HSR/xHXcdcuhvzF+x7jwgB9QMarS0FhmbSAyi7JnkP
NsLdSDm67Ng0LYgpUfAT2iEumDezbhLl6JrqefPk3BcxOLxIyKJG/biND+qSjquGbGm42eA8ze/x
R7u+zX4y9FWtgc72whfFjct9xNo/2TfrZd+mwqFjcswsKgl8BiEkTABGpGcZYjC8UhZgVRa4Z7Nl
kdqcf4t5uAcJHRTsYsaIkea1ZUaq1K+49m06FghID8x9UO3pW/X2NakUpEMhv6vRfNCUhNL8AnU1
DwlinevDRoEVgGOkmGYCUt8eOvf2gSzyyAUtcxtadQ3iwvAK5rxesHUlyFyToNqsJq3AMpeUfSMB
CFR8QlwVufpBTosvspQxISSdYur1gQpsUE4iKRaHXRv9f/2dCDeBOfak6m+Ow/NJzK8KdeiOunb+
ttR+GgQsu6RLTvVKpKV4iB4vnd00ac1srZVtOvyChWJnAefLSI1SZm40fgPlYBLD9OyqO9IIUKs1
Z0gnamKEqtsL/gPPQBaRZmQqQZe9y08k/Spb3H39j5GE2SBzE8ak3Xvr83k1ScKdyLTdx+C1Vg94
TGtilHgo2wFZl72GdYP5pK8z/H5mvs4Lo2mA31l9r2uvAr1gpF9JeB9VHTq8NYlWWpQfeY4NwUgf
25GgRhBoxNN1fJ6pPJTURKxhKqfcMdxif5X0JgNMQ0Vt6pkLMYe7hLxkAkXfXlLJ75iRlD4uMm/H
QYt1O+SA3/R11djqR+lIwA4QWRURJqEiZPmGL3nWbz0LS9qEwyHP7j4ifkw8iE8lTEmKYISPJSrV
9NfY1FKFrQr3Ohl+wOrxlpUuH0nUVg9kZbkzfQlN6V0gOLlXZ6iF8ZEvlT+9CUatl8E1KQtERUQA
kpn2Z8N6qwHxrM130M7KqxbSi5w+9vLD3XccRNpNqi/pyLGp0hfTNyvoG/+VMCBB8QsSzxdl09xQ
oschy+1FhO6y8AAjHUz5p5LgrXSr8aT15kwlH/j2I9zW4QMimVDsVyXFxMyesv64oObJD8Yv9jMs
GHfF9RgUL1aMjtuqAl1u9IT77gj0iI7YvMPeCU22M7W+kP1mRDJ/OqIeHBhgfiiotxkJuN9+SwwR
hnKm3WiabKub9KHH/R+Lzra/+M6gxECxLqZ7MgaLSaFZjUUrSL5VFPA10qBXHo2Ql0Sg42tVph88
I7E6WeecWWm2iYuvBHyen7q4abhVFqdbct4gY8VwEv/dcu5AHbM8x3BXplTc4n+J+SqoGd+pcVp4
odCnqIMJXxMyKiIRABwgBlhitWL5WZc9a/cyHozC6B+P9vvIG6UKzof6MPdbZmTgLi0bamMYm1Li
7uZRxMN/OTI2QqdgNIsr71AjxTaL0SgzTrjTadY9ydzpuXkX8HS8+NdItzgIEpfqOQHA+0jqak4p
hAcdCjUnL8x+XiUrur6TNFBM/qxmu7YCJD2mruNTqzLRkK4BI4fW9xtpggPw2KXBXUt2/COJTk1i
I7zuDbvw0x8ox6aovFVqEYN2CwCgp2KgV3RSQbfT9dOj4+40TSTRPvTwwLBrgsq6IX2JQ0SzW1g/
tkVpvDdh6LW+7IfVLe/MZM6pTJUyF1Q5zmOF93xPqL37PRXIcuWnNFJQWm86Ti6DSxMv3xZbakmo
gvK2NkRiuoL6imfg1kxXwciHKtw79k1oGVgIE4AXgUXkKBFzpIlu+K3thMG3PwyIlIvSYbVL0w2w
CNFBvER8Dp3/zLX+mQQM9ASVuyJMvwzWZ57XT/zRdHM5UTRVygACS3P2KYaYoE8G3js15Z4zdO4R
cV9Uv6engo5D2gN1Xk8LcRjvQsd+Xju2aL3tyoIaVBO/i4NmDg3DXCfcvW5GJv0zyHLVYtYRUybh
Vh7i+etwZ0lZmr4kmGJ01gSEP779yx56pXcksihGfDuHl/Ez799YjunVo6BDQ8bhJSeP81/XgL1/
0YYOAk8DyVcGW5bdQrdFT8TRg7rCcO6phdEG9svMQE/rc5U2CedUfpkSC5YWLLbu9iu1USRjTT6L
7bh5Rl5iWoQfV98YJHcJ2A4sz+An7vi82RGrlK0L17B+/jhIMMlnKfTgzMzpsEdHa7EJK0ADZHZm
CjKAraxJc06iER25seZihThrbF67gMmoH1inAJgwbbg52TwkqpttBiktihm/1j/ry3PJnfdqiQUO
VctNEsN1FEp8It4T7wNoLuwgrywxSumHQtelZDKoWCttntIk3WIzs4exNUR+XBO8VtjbV/ymuAHr
TZm4uK+wzI0vCN7uj5C/uk/6qZQ36bzU3pattg8k83/aGjI4PvGWlUwr9nJcz9j3HhPUbc1fP8GW
pmw++n8oWn8nhGck9XgmKowZZy3xKDgNq9N6sUOAQcXEHUx3fWJs/Bo4HbJanp2F6tLaMHyBLFxe
2jW9UolXqmQ1pms/3oWh9ZgZQnprGLK1lJM/3C1poWTNDdwoJ1FCfTfrUMDBXd/ABzo5cBA6Iqst
pW/B6XV0DuVRVG1DqtUoAwX/BSh8BSUkIZoZiXJ5i6UX1G8aucj5rlaNwqCEGlc2S8rhuCNMggIH
D3+Vc5dN69H/Rwphe+trg1Y0euEPXCwQA9qCiI6npEEOv3vCzBsPWxE/jfXrR9pR4TvWuLfCNCbg
rIk3y1Ryk9D6iQmDoPLphIhX/rltK4M80Jq0KHP815sEiDx2fCjGq+6R1yJoxWiHPvwrnkTVZTt8
ac4sY6fdUGZsD4E9bJuCJC1H8yLqDD3G4/09218GhIhqRk6XDbj25i2EPBitvpMk94WE5kC5tRqi
6D270PCtW93ZO5yrEqYagaaNm9RkGmsO8I76P4a6Cx20VEXJJsEXOSdGV8fJlsprdOHEy2+AaVDD
iq0sJCmEGBn09tLyT+e0/r3eD8pxgQDGkaF5p+mLOrYV+jsjKBidDrTUsk7KH55FjXJnWAi2Zl4Z
E0p8whacTsuh/jdDvWOzSWs5gs+RbBrQPFXOwQjJ8ECSI47tQO8CCVJQNpMSdmwUX3Hl2I3sUuIJ
2RHUlGdo0Ufg3npVbJYDY7QL6/02JC/5A+WrAiyEyXF14DkqnxzMxTKwyvc8KndrjYQHYsO0c/qA
Va8/RHmC/sGHWJax0tGxq/fIzOimB69Avd0uDl05P/h6my36w+OQWIJkUBprCDY5eslNwXTJaaF5
LJgucIzT2Uk42O5VJkT/5NLJww8JGiWRZRXmRhdKh9TMNFnEdoPJTKBscS/jU5AKO97s+hg13zyy
utjpkkay9XSDyfXBaVqeBtG9HPxteympbVZsWkpKzr1lMxYWlnPk/HIv0OXpVmdyVdfwZAV29rj7
OBdU9G61TWSKYi8p4z9eQfuVkdeRRRPcS8WQoifnjVi7D6Jh1/lNC0tGC38xRSakkcKTOXIn7Qsb
XmRFInGuMtUPFe0pxzE+zgymkZDEuWT+rL26yev7oJ1xj5vnSXsOxgeTTWyBeK95+1kdYs7Qr/T3
AUy3UvgMg9yP1z7vo9rpktVd17WuZngu4ZwYy2A17wRd1rIhLhS0+hFjqgjpmpHaLAyH7XxGWhst
daqWUARj2djwh9Q/aFYdaQAtDUvDRasa7Yz0I4BFdanJVCp8Ybl9kQq1XiRJSlWp4X9OlxuQa7hc
WRGiNjOqzyTk6ZsF+zAA26ePcDR+G8G77NTknbfT18ESLXsVWg5Wy8GSS6bY6hXGo8ZgkWORBqDu
jvnPQRLehBukWodeKL988COcSBUlCb0lERDy3XCOwMnD+vsMRoLiNaQWMIUcm0XK6gpsoY/S1zhH
xJrgz4rY9sI51eZ2FWG3g/sR2mcfSDA+l91pR8ctdC9VceBj4W4X/esFVAhtq9S+Lc7A7qhrwFKV
wLUa8DpIOQXSuho+kiIQnPX8UoDH2sOyzH2U0REhgt/p6amAimyaNpBwth8raU4E2CZlOH9gS+Eh
yhCZsWUdJbMPR0aY4ZxPL+ACEiZqKHvWjsBOxv9q8/Obo4cReP72WJrSSBBbYGTRQz/BG/wyRVeb
xIQBQ7K4QVikboWq8+mubkRWCFN0m3OBqLBRxLmcxB9yIws8ANQgt5KvLXgLQXMZuSj2uuDv7vhI
O4tQNDV8en86ZZAVhtos3AUhWp3QEIAoq/wZln+SzOYvDXsST2YmeqN706r8oEPuAuZZTQiwaGik
QADp5IeBFHw87mYyS8FVCW/zJQF2OmLsNLaOyrT8NVSj014XhZ2aFFHMy7Cr9BLXYH0zXyae99Ar
afThY3ZJnkZTkRtXvPbOrr04KaX8Pi0v5+1D5IiAtDTHeY0thpFWdkwqTYZkfLcQmwNkgulu01ao
AWlJSiFK1638XmgRJNm6EIyCA+8GKyLGzkpLdagG7eWMZIvQ9RVgy6F0oiugB0FbF+PKtDds9Sks
yUyPRTJSJOSxC5LxUy+Q9rjHaHNHJDElyDdPgssr15qyNo0As8lKjNGLktxSdRFLS6axwxQH2nrN
oI/GYLlbTKJzuk5q7a0UPnVNHV09fqz0nCJ1C3YsPX5+KJO0XtTQiapG77jit7jcSuaoGamHnL14
qpDmliLMGfExBNBH0cyx/Boo/8jrHWJ+cwWUsMPMDSF397dwVvhyrUNGYDLp0L9hAIRJ/kox3WmW
O8SdXepY7vf39kkwDyZpTtvxKYQ1dKm+3TopP8jTp93aXzg3PpsgDn29YTY9P7pPSRYx1T1UZ9zf
eCZPXhllzz+AcJCu/JAdqRL9qxlkbfjIHK5cK9sY2jtiTrP3esnN6CBVBV87gBhfbqYIoPoDWQEf
jIpBjV9tf1WhlfTDpBDSP0ABUVXMQZthAOr/FM2/RZEDlEV4r5mDdEiUkERJ+yBZAi1u9pQ9DGF2
RVdM3QGjbMO+2J5R4FjhHXdoJebXZAvXDqnAmWYl0oB1jLEW4un+liPIfpxv9D6hPpq/0xPmSQFV
luBmD/OI31vjY8tgxLbVT/UUD6vkCM1FZR2mvwZtd2cmuYxxB/DxVlvfPV9rvwBon1oLl3jD/Ncx
4/y7RjQ1+jDR9M3G4Q4DqpccjgKM1e9vtrI+N1iAKDkWvXwVmjwCe2sf81ux9WmxpN444nLRCwbj
M/U8ZrLuo6aZvcFeTjPiUwNJRd13A18X1JJQYv2mqFKgFAtJEIvgvynlPvKs7FmramlMQduoJPsF
v/sKCEl0TkTz+XXMfl1QIGzKHZguFilMNFvTuCdpOusN1HV/HSznMpJsuEkaho2qdYSPxXAtQNpQ
uS2EpDsOxC8OLk76P2HXxXCo2IPusRPQTprgK3Bxzp2X2n5SFojJdMbpiSZH32IMjobFP4W08XQU
6PYuajHyrukPvHO2CI7+alkJYfHb13a7LIXw5GXImnKu2NCKH+VTb12HItSazVBNNHs+wucQNYUT
9zj+gqdYT79VL8K5yl+NRRSoVMgPXssDqu9kXQHDCXT3NrSGKkyuiyloBTN8vnGJgoudvG2yz8lb
zrmZHu4lRvtUVLjH3DAZbBLVLlTz5y+1s21VXUe/QCvv7REN9d7cJz1u2GlAaiylp34IBfe5OpLi
4Vj52CUEdEn//DbUO06sP5cHrGPMP7N2DrqULJ84OlhaKq8EdiRZJOXm/TajCOK+YWAukPS9HPuh
+Gro9zRBYrDXKALzG3LRH4qxclluSLcB5UjjowQ4HHAq6zPtDAx/E9IoIouvmAFHfYc20Qel6FY4
8pooqRxylYv/yXCIC+giqTPk6DSjT/b4RtOLygRd2/FQryQ3lDEHYURT7FButsj5eFvz3dVViarq
UWJgOzOZSZltNi8jo4DHqizYYC5FKwVhJP96apdB5LPLeOjO6iZL4KKB+whlM0wIDWzGGCpldvJd
tY4wQKhF7mKQkscKV8HjkJuS4qFTNarQZ+54G/5s11fDIN/KNQkSBRLu7Ol9SlbpIodpPKxjrY2W
gx+qEaAbsKVna6P6tyw7qDRyiMwX/iPoEFE8wMgkTMG02oqDxnUsjponuyuPAfCBJ/XmYYBQ714r
Oc+cxQh0d4kwS1xMXgGVTvqrnknOuy1JGKCRVrBhvhwi6mgq7xl7qd25r5qIlRE8POBfWbDt7dva
JKORprKScbWeGJbwNlCwYPgaJSfqldHzOeeTox91YJ+xCOHbZtHuxU/8wIfuFnZWjCdbQlJAqnJR
9LCgpn9hhAJnkqNAuZt3RW+xdt2WF3q9NQ+MbxAvc8+o0seOlgkPWA7/xqmbJWDNr1J400UX83cV
w3L3pX9aYrr/g8xWf2V2dueTeDUN465fN9vLIkfDsTbzs+OY4naQftlhcdysiy0xkSQqXr2mXwql
OWMxQW4XhdoXBLvzozelhJKCf2iQnjhpJTCUlkeMn7YAFQ7VFy5eCmW8avKjklzoRDpD7VkG1iX3
NBGznbvPym/OWGnR28sTFzOZMA1J7cDV9Xse+EPMKLrWPCdzbiySp+u0IKdzjdtA8W84+l8kZo3v
Jbx0z1RagnP0F5gm+f/+GlAHcq6RopUngcuvv0bdDoj3/WlviTFSV3ZIlGAfndbJrsdhRy27u2sW
yHYtOOA8poHeTFIEde12dNizw32b6okJ00r5jibIRfX+0+rT3HWvxefr5Cflc4KtjxVISmWHuFH+
IZaTxzubu6xZ7c+2SRzWmt+d4fSjasKLenMKrIfVuYPx2mwf7sw5ViIv21+MUdgVBYsVqTPHZUx8
H5qPAQaLTb8kJExisGxh+7e1o6jRUz7pkemcOOE+sxTjDwBYQ9KEg/nhDN/8DaZlgo4tWJOHjeMp
7hTH/Q5+WZJWRn+CxKqjX/LETPtvHVB6uJ+fKl8KBsGIZduCS0SnXGx9Y78+znFlXjp68qJsmdi+
CgNDaQbF9KWvyuc8xBWxtp2WVE4u5Ki5/15FyPS7VbhLhOzvJlOdNBKBZPlkmFtHrGoQIFBsaj6f
8Us2y2iMC6wheIv57T0BAa+212SAuuLW8966VMcRUUP6Mq0j2V1FqBR7MKcqN/v5EfgX0WZzzYo3
U58sALpU73jYPGwKhmFmFss1EJqwKDKoY0oXniALqr9p24bv1Klzan+lkJL8iLU1DLeyeJe+r1+N
L/6FwrZETHGLEzNHDP+Tnf2ExSNr4WtliSzR5cA1cDITedHP0T3N3zNQ0ePz5zoHxbfVbIXeqeRh
GZ5noZYYlzdgo7ZC3iZw8Dy3kMMXRpVYrqJ0T+O4oHWveAz1YhPRf0+iSlQr87E64LIjDCGYUnw9
grm8JbAbYgSwaVU/G7hX05UH4Zu4BPOLsMqjoC5M4Y8gUKHNYKmdCuDcX6s6u14y4ZC8fC4TUaUC
AJaxCSbp2ZRshnBCbTEu20+mLjwrCrvI+5KEQfB4ZAWni1qJZwb+Yq08ZABRJ6QFcu4+TJ3urkt6
f1L+Mq/J+mOF76ruVxTuOaFaWryxhhUXCXDMp2oOtpBgKlI0FZIldIHA3Rxskn3cpW9iF5aR+rUU
xYgRIxYKcDMFkvr6AcYJRffQSxAmzRyOuQ9JtaJuSA3B+cLNOeF0rMrVU3CJW0U9h8FwK2aJKYMQ
Nbn00mKpwc7lF0maRSyrQmYAWgrjIjvx8wabP1RDRn9h5VkJ5xAcQHzsxnpKgfHQwHuy9sakEwXQ
1iw8SFk1zGU4Zjei5+FvaVFJpRDdTPKVWnrvZZzkSt3n3rUhEhMEcXKz4F6TtYxU0MBcWPS8nKaz
eCq1ceipMNqxAgj3lv7gJ5+2qXAHPljCp3cA0BU/gtv8890JiWA9JcSL9Hr6HSYGv8HathoQR96X
r69pvpAY/y9VfaqvMAv7VhDZ4fbWx+a65hQPPEYLyTwPhmyMthKy/BMkg56VykFes0JrCnRoTmL2
fgJjE8GkUN/yaIOeXEAXHWuqMdE5Tu8Pf9AaOzEoDXavZZHE6+AUmlIUwDYo++94dH1xOo/W2I52
IVnnee3cLpCT9ieNhvcL+OW5V+gUXQmxbpe2OEbioXFXhh15xfYh60sxbpHdCg++4akpFSDA2Aaf
IGUHY9ZOp8JrXO31aWY9JFyi9wM6tnrqMuVR2vC67zp2F5hJ3zt9TT7O8lPTcjQTLLlzYviEYIBQ
ryKJQyrKjR++pOcCqsA1I643jnqSypisfx3QLelxUBKpPSJTu7DYehW8Oeo0SS2pDVpyZQW3zn4o
/4RV6bAH77PfKuruPpwKG06JdhTwD5fDmO4xOGxJb3FVDBV+45EfNqorixaoHOqMwApiwiYgKCWy
0Wd0pH6Fdbc9Oa/oOFP56DL2nAax4WniWOeC6HQYk1GGKjHAgYCJaMYKiPGh5hwaC7UbhQirzKnU
l9CexHaEYMGPIQsxV0TspeuoDbj43saR8wK+PsDrQez1a5ErLqdEic0tKKDbl/HPmUvP6OcSyozn
WFH7aOb3va1KqLlIDnY+v/RRe3PIgqBJqDwZwZsMS86Kh018a3eo6ywyXqJfSo8wEpwrEeXEre2+
dtBLiHZSmpDZngRillW/urVTy5V8mHhTHmrZmdiSJ8K3FYVD1IOkrKEcOXpB+BLehw5Q2CrNBfla
zNZ9GzGZyk1caO2DDKHftyucTp61I/XtBDrNkUHxF72TIi/6ytRwkrwrqNHLCes/t7Le6al6BIiL
CfpbyWSQOXcQ/xJAqB1pBW5O/rpxSPu6CenYghNTa6vQzPY+cZWpkvJKVSIIW04hImi7/5mR8p+F
47XYCtbbO9JkDNUS00+XfOFfHSwCPm5s/as74IBEHIsR4/8EwcEVb9M7TP+vi/j60n6nTX9SWWTQ
ONDbS/PgxK3sP6OJJyo75hWSTnLUmMDBpD0lQPaC4t46xCcgEK9hs/OmOxUXpJXGXWRP6n3OchMV
G3Mn6NAh1U6foi5iZp+Ny4t28SRmVxCJWQG1m7AzIrqPPNo0BZfWqJIli784E+Rw0/HilR4YCyDG
pu10Qr4jf/zx9Sw7GPqdY3oVEtc6zE7tnSJgvIwpoVx0SSN4/QPWhQGdw302AI25GA2eAQxG7OIb
k+AyLmNluTwB0AbyRVOqtwdeDIRu+z+uSSx3OS+/6NsS5DzksTn1Yp3UwK4n1O9heIShFxLqcag5
IByE3LsKOHWZ3PEHIw+FGTiH5rnepfAKQFo2JEv2gGVUHRA4b8Jn63bDf2upEYpsBJpgRyT55mEb
t3EQ0QsKleXjpuOtRRb0M+CsFrzHxAtlopu1pGd4mIOYFhUrYxvLha8ThfcTdxKIPORc6IZ3V4SA
c5euivD0ojPqNPAqClFaqzS9CWY3oFahw8OB64uT/kTNk5YqsEhhpeFlsQV4m4t1e7odjx5nryuW
vgiPhclllEExmlc0To4hVvjiunK5t6pJ+PQyLoBbCc5NwRMjniA+4cBIq6SoRP4KhZIA2jihLh6Z
2G6APp9qqTxs24MOcvY/3d705N98FOyGoUOngsKuI4DCyBjj8eVFqZbblRcfcAlXS5nRbrGoSge8
1JqO7W8pSCs8yX7AJZC2RwfI8NCEFYP3ObIpxatvbbB5SdedIglMSyBwhs6/vdgcnAm6mCkoCnS7
JZ2sgxlcSFCWo1l7JKPshWSjBMNKmrjk0yuSfYfYmDH40E2d7WqJQXCvu0sejSA2EwNskxTgynoq
sTsAwy0sbTLmWD91A2F4LBBxWpYxqUYwh+nAn7VqYrM4ZEv+x4Y97RFUWP6H58YfE2F725S6X54J
G6KIc6+528x3HlzOreGAgf7Fdr9ZSEyl88v78wXyDwSlQ2919a8lWvgTQmJi94qMlgCTXH3D/WIw
iuwpUzWBk0nsIMXyVI2WmY+4rdKwPEFbiJUbl1bRWk01+d6C1wfg8Vg+Kf1SOuw7JrDoed47Wxu6
TSxFm2iU32dDt+FQy955H/Dd59ACTsEZbJNuSZvinoDKsVo3vMZPyCpekIkyrT11WnngsyjjCakj
XjMzBEVvBziRrC9CjWyOsjqM4Vd/k1xAmGsmTJ9NPO0DZuq0vPZwtqO0dOfteE+ou124iY2SfeTs
3DdyqK6wwFEHACw5N5lx/j1ng9mKkDcOPLHOJ5y0u3E+YYcuDX0i3+853nWURHplWEuj8Zhp/52u
M2p5fCgh9i13fklJ7FsprpWszBpUTJyiY+CIvr9T9OSCORvRhHX+cZ2M2TgXiGD94j6hFZE6DAg3
S33yWI+S9HWsgt0tkyDTy22+Pj9Dcq+sR6iVOSPShRU5pmlGXYcvowE23Guln4QjwXuaSXxkda4E
WnwHZEhfObTt4HC5KwsblJ8KlCeWQbatjRZft9BCNLZffH06eVqxCpNRGmin+e4bLYwc8kkB1dzn
4Wlo8EwfEVTjxWltW3dmWARo1rIMyb8sUh1zEKPhkk8fL2fT33NLrgCmPthCEUoErYBKaktZgOv3
hAzOoDmO/FCKGb/dMq1QknkHRQuE+lt0MQBrE0ubCfTKWxRLyT44kOMPx1ic+Y0dDt/MSGDr0u0N
57g+RlC0dMulFfIhYSw+V1ppazT+rsiywFM+XILhomZ873T235wXSOHCpzWmLkpjEZL3LAdfEiSs
8ovVovYbufj4l+DHiqhHF3aZGceBZv9PxJdgg4+RSG1bta2Y7V441WtZN50uZ/0I3Eb1vhVcUbq2
TMTtORD773f+rA+RueGzP/8vX+7+KmmkNA8ZPBEtJ45JjNlyThjK95vY6cmkVC+ljQSF/VclKi6b
0biWHXBSlt8jwYOmpUTytTbD8sqgUIwsQtWgXolQEwzMf+4W7eCt4vtqS96TcHgj7lq/lXMzNpPj
KjwHWmYKGQ27WUXiHcU5S22gFFbAFfmARZvujBycEZhzyndRQR0bIR05g2+eOf4fD8za+suEJlmt
np0DwgvS251XGWFADNZBUx73mdvofOHwnVKYNKzCt3tC7H+rLyAECSW5NQLc5PiJCNU+nZHMZNcN
fJy07rcMNha+qnTJVQhlAHYe68CSz2Wv2EarL2CnWPklJ3y3dNQYeeBPVnXE+mu/dPeQFPRpD/ZW
aBcTZL/DEV4n4lSUltQaR3DpUGB5+MqKGJSKKkmaAfZwJn45ixHTbBuecCFCXoqabyXKfyIyJkY4
dCpQBgx2RP/hS+wfQDmw8d8DWf2jj0S49esBzsN3AE4pGMMpVMd6krxDxE1saXNh4YOp3c+a+/y/
mzVaodi9dpFzMwDVpQGpduL2hRRziE9MvyfKNLeSvmnD/UQqBvhZI99iA9L0qs0lcnA6YDdpWrBZ
P+DMAobIN4Ro9vEC4a2xw00EGGq5C2wFpYQ9B/nWmEmYEbJOUooR8shJWVLaMD3PCXJxo280HhqF
8h+qEACYOtya/i5MZ0QUhkZuenIlxu8M9bcS7rkwRV/Dj5rgVGfrFJlYvbwEr2zBo/zifJlqGcBi
yQ2ri/xRJvUDBcKrNl5EmlJVB9LKAsStbdlPe19qBwjsAsFhoUMDLFcAlHO3PVmFT00IGOXDn+K2
1GBTQGXpEBKMHd5zbormLmwPsG5C5Bj2ha8OH3e4DlKdPGmZhOI5+air/huOWwoLMjuZryHKU7JL
VbiHVUzH2blHk7i4mUUzs2wiux3cxDKDSp92brJqqY7cA+Z6Ef1AIzZcIdqog2IpuKK2QFdFDKFL
gtuSZ0yPw1cNe5IayMP+U5m3eVq0xkWAdBS4j82CjifNf+YLUgtsRv7s80sxgBakOoXj1gy4zP9e
NY7FHORsz7SaqQcdcWJ6c1aEJkAd95dmatmRZ9x2LWvDvx/gwneTgVYyDdZEJwD+qhYUPs4tXbff
a2bqnZ1osSX3W7x0XcMFfAkUQN7mk07Fwhc1791DL34NeynTUQf0HGfddQIUNzcmXm7F+uSzgrgc
niTF1aJxawrpoUZFQhNvK2o46pj30t9oTwoluTudUY0YwAlFgcNdNJcpV4klK1xJ90HtpgSYdOWC
aBvX+gR3PzG3+CGWJa2CvG54b7B1qPeQ4j/pU32JaTOvfkK9mIo6KM6dACrHgwb58FZ6E3f/kMcX
+Rx/OkBtc/NutPuTWp0dvr+nu/WnCHtUJ78AUO3GTRYB3DyvOkdxcAQnkbb4IXMqviJ1Pb3nVHO5
saOf/Rw49dgJiZboZlCptPWxpoB+QpLIwLm2kO6E+FQ95ZsXx9wclYd9JoBKMmS0h2GiBm3o7E4o
KqXvHXdBax4Ecx7L4Zcq3iOqZ4veRq1eMpQ0XuyJVPvNTvfndMtHpZWuaf3Ho/ox1wQvPZrTesnK
hIZA1zS9ht/aikWV9M/MzWmhMMF+x6RKgJDllKiHHND3JN4lgcP+7vBz/xyOZcUgpRBjrZ24g8M6
KdQfo1lW+LAIOfu7TMMGhQgY44kCyYjhIIosWjfo8X/7Y1B7HsS0ymxTePIx/vcdK15Wz7wDooI7
c++L7XrtaIO9Ogcx0kWgkXYN4eAv0HV1Q8ba+DWhXbHo5fnc3xxUx7vTNTKZMf4DlLRCEunfOCCe
tpQ7CZlTvUzrkRSC2PZ3XIhb4OYS1VsColge3d/TNG+MqpPFd3fHyNITQ1bXfN7OiyEahOj5DWGT
YiA9CRY4xBMOirF3vc2Tqipxooi7Vcd9MqQTiGH6ei0sMsBA+0/WaJMro99Xsxv5azr6T5BhwL7K
FxtCOSsh3HA3sFxL39ZHtOUk5lykI8QPfsLpqJ2W0xKWcOG3UhOHLOBNYcknb0rQVVBJtBYDJpvz
jFF03EtFtmOzuebYMKYF7S6EeSz+hrHGnKn2wAoD4QbzAu/yBm97FU+YX+2k2sT/ts7xVhixBc/M
aEOm6kVB7iZCHbOvXEdvbw8StUyqUYHkEOSKay5YrIT2z42K5JB9Cic2e+yI6AxtVmwxsS6fsTZx
zKdYP8RTLohO3LMVWowzjeVAAm5x3n/OnY728qjhRD5qzvSievdWHMvPGatRKTaNNoS99f+MO0Hj
JapmSIN6nwUs6oTaxrDUPkklXLSlrOkev1TI/8/bPfftq/p6rQICedE9QVfoRJ6yOgbU0v8bhTxf
vxY4qEcHPysQ4GByavTDUP9KO92Xkp1trGnEuLK53pygJuFTlWdiM2aqrC36foPjrUm5H6ph6l5X
SeCBXWxhY8WJEpzM6W6kd44HW24Htdu1Qx6LU0p/t5BITaWd/EPB6OWkaN5acgLb7aUZ8zz64SQu
nnomteKJAjJ342a/WMpoZXtWln9BiqVk121Htlsx8Y7UnERTn+PwtMnylmGlFMFvc8gCP/B9vFaX
p70oVxMMoFQ9HOeIGc0crbIhtcgcwJ2klS5zj3/oS4TWa2kTx+mdRx7pV48b+NrIqV34Md31s5v6
M7qVxnzFGEMLOUw57C23hIsGXm6J7koVL8cr9aCIa6+irU5EFDUPd1toA9kWHbVSOsO8JkK8kG9m
oaie7xI+mjgUW+e05bOFoc23tA/H1EpGLx/b3R6Qjxc92th0miwwdUBWl/ml68izNxWWcAgpM9rc
JCRMRYiYttQ2Pw84NonuVE4EeRY4WmXpjWc9QGKMNsNhL+aj9ZieSDUN2+wOMeC/eRqzA2NweuLP
xq0BRqlQrH33bpdzaV+yIS1QRfWg+DytehltfZeypYgPw0nWilza98DMXh3q8ywvizW7vVmYkWDh
49fT+ZgrUZPU/2r4LonuvJJtTNjUCEzyzADb4DWp2K0HpSzaEklbBshK3ph6Gu3aAf3JeG5MkqcQ
QOPz+CCsC1OtrPKlu/UyXzZyHP1oJNjZdoiLAaLuv3LqBSXyHAnoRGICZOcyPJKlvz7qu2qLKLZR
2/lDCNr9+7v5m7VzVHKBBbaTODnIcMm8bKcX1U7hSXvzwITGtv9hXM2rlKHIjAVqg2P+pYKuuVET
1fziRWjx8CCmHlaNSLfmLmvtyaFFwbT68GYvRwaDkdmqCSFlwOE3aoveX/yK7u7YYO8nXzO+eFPP
2+b9aFf9Jk+DE58+jMUAMfAcseCyHPodWLhGevhQJp/2Mx487ORqJ7aJC5y85V1Ryy3gJWIVJwrx
5vf8mOy2EYz1qpWXzAQCeBS96RTppIOqk/VZa+xeYlfuXXv2RyOZSH/g9bmYgf0niBL6AWXBhT32
H9aHPUFFK6bxiVGIs6TVTc/iGKODeqhgbgJv53VMAkUjNGPpvA8EymB1lJPbdz8Oh8bZ00dG7GhW
o/zLU7buHn0pOvpvQM11Ilaz/mbf+0uzZx3qxuMVK4E5pEmQaUZSTlouchouIS8qOwvp1Nw3hXkR
8WAfbe8b54ivth8aC3bxyE06hqV3HjQ1vjzDXAr4ayN+YZvlxgHh6OH94r+EstjjDdIH3GfS+Zw3
ryNHvKFfMmsu6Li467fNWhiUrCnSceL9dkCcCM+r4kUWVVpmy48HBR+hViiQwK0KyWxkEbrWlwlJ
2rbzoXz7BNasi10nrV2ZIQ6RzbDqRQ01k4Xx0gOZ0DU4rIE+FphnDELu0rESKvyPSInMXJdnI8At
OQgAWq+IBbMMga7TLErlto4n4RlZNQ/t7piSNNx9avHUYiVVx3HQjSnE33kUJM7qrjB07Obkfc3c
5yFzT0FWKdWLOrcv8r1Qs9hifD508f2WLaeXE7IaZSS65huzvfegE5NYzus+rDWLILWhbsSQr+KB
fHoKxDFkNepQYO3ZC3rBAU8EEvCF12S30KN5jpvC2Q2Vm0g3exE+fkrDCAxXZC2J1mv7PrUQJQad
C/8mmXjn6EUFIqEoR2Hn1UIDvGW3+meMSELCGyg+l9TPraDGT58tYPvSQBsJFECEug9ICDEeCJr9
JT2ARGWn/MQYjaR/coaD4R6bPZ56UyqEKkYsIZiwzp8+O+kzOqvXwZ4wpQkWPuNbfMgz5f+ri66A
nJEOW+EC/DfkmJ4tEMpvRKfxHhMggaZ2kDK1VVHkBv7b1F8d3xXN0sbjgzkU0vr/sRiQZsNi+5wX
76z8Gn7+dBXEoJuhY2Ayh6GhY0dnTydGoIAZOqr+otlpuKqw3B25lurEWno3iAlwQb8lQyQfTg41
vU/37BgOkc2hdpgOOA66i4y2I1f+h+SiGdxq+io6YdNnSDX85ZgMTB0IBkDhrR9qID9k5pzIeYT1
2qpArjq4Dz34jLg2ABre5EyT/fZVr1biy8ybkXjo2GvxqVST9N1k4xWvo+AJ106zgOUZeWYZGUqQ
cKudNAaXanRIY1JyzTjbWkPId/FBA3tUWfHnzebXetoIPFdFUuXhrRF5a+v7ChA9d6KS+3zthlIf
IZJ/7LgkNQcOG5FgJW4XjLGHPF/asDZS0Ml9de6iMAthFmpVgAhcdjEFqO+Bbsd25HHurzLNSxK4
ka6FSM16ZnQcnlREE3Kehpm/57k++Qvs/UIV9e9GPdKAshzqlQrEC2zCXuM4lXL7XQzQjS05jsOO
jNaXJNEuwb5z1hPRO5Yb8jHz5uMjdbk7jWxwZ1ZWmdXD5R0RiO0Kx1q4C1nKTfvOwm91SYYnI+cl
PRVdyL36IyKhGVneTBsiTj34UaWMfetUGYWBtCcfaSE/hF0jM8z+MaW2skLPSK5Z/8NaKkZk4t67
XxOZYt/cV1vj+qs3lVDDCGT3TOksws/myMpOxsrMh7dsgrCkcqrWoUIQHrekWRc/ZvN4pXBOAuw3
GKJO23vYL16OGPyXxkw3aI2MabHF9KPcWckwhvUVEixfKwdohXH1O4URLVlvsQFb59jSZO0S1nqg
XfXeClwoUy2s1TYwxru8tkUkgv4+b+dME/9X4XSktVAGUiGQsuO/LIO7lfOCJPXoV/saUcn23JmQ
dQe+K9GlrpGpUuGHq2UaJL2DhZa0fAUp8zlu9sS6NQey3eA/ovt+Oz78GAWYhkz9esvCTyZdrHNT
IEaz0oH5tbH/KXB/SSJT2jKexkuX4ZOKzn17gHV38kKoagWL8LtXcXe8FdwKf+owD/im5dm6JxN3
794bdQKk/DSkJKLn7+a0TlTZurSiVEjvAu5lErK2y7QN+RQNp0K7KdIZ+2gvbYYzmZ5RdsVTOeDj
fEOJlGZ1X3SBVzqee/hmvYgct4TVD9tVyaUAtlas7GC2kg6f9AMNEq1UaNltEq5WyDy47e7NY4lA
+0N6ri1QqcNIX4BbQ4q/wXAbSsL7VPSt5tspO8qPM3X0G06gE2Nxa3dARCHKjmosm5xGBjJVV4Dq
SelVI55l9zFKyYuupP32cSUaNQ0cUiL2V4Qp10xAZBQJwg0DndmVg0f5q8SSqgmBcsToOFTnpBlm
cNVpJ9x029sGoJwaiVYxDWA0pNlpxRV2TAPclfFFVF7+L0+dIHq7r05Af4l7XHzJa7hrsDRwSZ56
IsotEWB35UDW9p8b/FP2YZVsSfCUFK8H9zbTn3TxMRjE7jq53elqMoAu/ILD9p1/uL6CRAF0wf13
FzbdYikBRBRUnrJ/RU08K+HmtcGb0GUuoajEjeLME2t9a+2QUsZyJWpT+3ji0RRWLxS2ves6XrgP
cQF1aJg+/q3NlmpNf3VPg+2f4aqFgPO9Xv4Jle2BQMsHQDFSgHi/LVPH1j0LZ8eiKR1zTFf+vJxr
ImNtM4g/7EnBai25fqA9Oub21iu3QpNAd6xGJyG+iJhIh9O8dzlC34trWazxj6pOkQZlIi53PTE8
M6Cso8a40Bjrd+pB4jl5ChDDEki2mE5A487b1ctK5h0EJ8MC5xDI0Tjkej0Qf1ifE+qThP/m5Pek
oYj4NgJUsnJpWbMbX691zzNhBR63sFtda6A2c5IMZUAlo5VBqmqdJ0CfyohpHPCYY0HgZhF8GO7u
faAcjW0li29xbG9pt/6o0NmWluf6D2raJp+FOWyMLPxQ+9jY72I9EMzCJRbffwI7Zm612afQ206r
2n9GYYRUi4ynUfe8KWjxGtp+Jwl6uo9fH8m/dUGcUYy90BRrrs/au/jtVgIqiisQ/xvSeAk2rSSJ
vXuZ07BQEOHODZGTxIY7qLp4/6qp6qUaT1gqmNIOiDG0TqhjV0rKfr1UXyCGG0hg7gAHgtg9nTga
vFNyeOxdZJJ61XjwmvJTTKSMhytsqYwCg7a02ZilC2il8gbm9gcu+qQh9WFwMpmyVD9egTrwteaJ
DZF50gvQlY/ZgEPrk6gTqccmEKk8n9pMhf2NorYJf70JhDyzvx8JlkK+9hlRpzZelrIJWv3jahd1
KH1zqKwj0z4kjwcg50qiMgw2Q6G2s6OK9YbePWWZwU3HqtiqCHER3F2hG68o8QMs4r5oMWTLKpVn
O9Ai28dC1xVR+gJWerrwxpas3BEY3dU8nLsvnCjecAGH464O1k6gowY1TYinzTpnafahbS8DVzek
VBRgv2Xssl25i4sricRkrz6FnAEQ7k8Aqhaw3j/w9w5OJMnMPUhOS6gATjYlHwH1HWBlEGO6TeoB
6ZjzxU8rbYrzu3JgjO33NpIeFF+kZkYK+aaGWSu/yQmjL1RQLRx2a0fxB0TN3ys6dfLiGyKgSpSP
12vviPe+gF7Jd984VNJQ4Dh95nkV/Wz72eWDNwqd0rMKfQkQpn6d44xMKmxD2b+lLYlfmAtJ0JuF
H63CsRiIZbmPOZqVYAT/3nQgANfPfQqCnSEKre+DqDL9usmExzNMSlHQ4zJkjsbs17C/bkdHZEA9
eFLq05eGgOUPCzRPQXtB7xkAwFnP5aduRi86aFOzN7uS+T2NtkdIcAbWx4xWRspBwQ5l9qrq97mE
a9ktCmWEBHu7w3YZ4V2c5y7QZzXqvVNx++GiSyMwITcmN62Af8gf4+oBVXF6Tr8+e1FsKfpvmDV4
WaqS35bvhzMhFb0idkuVzueVkhcGeWChH0CTebQ9Gbaysdpr8REyamTHODu0oC6k8GDUvmBAUTRM
mfULl7fVxbe6zVqARRrsb9gglwAnTrl/WvzkkZ9RPtaT2ARYmMCs+q1IXps4kEt+70mkhSagWf1u
57fqD4NHtCRChPt18078rSBIkPknxryuGmJ8QZi096I2pmaAHDMjtfdYCaPGt6fdj+ofywlaN5kj
zlBtCpJaBRcxfzJi3oM0wWbV6qC2+yiZXrx/NpA1m6iJVjVQBi/4X+hpuPXvoRlKhl9Ucye600ME
nYvuYb7um/n7QwFV+T+kNKzqaHwt33eXNFgSJDj0joVq63hUuY7PiGO+u34EXk/R+L5gXCVkWRod
uiaFxio8XfTebDx8i4EFnqdCLkU4WXVmJa+wogK+xGzVgrEc2RgrUCg6O09PQw/fpfiqC3euur+O
8ZM6Nt4I5D4YnbItsTrTsYWSIFGwR5WkvFS2oTS4HTibjja8hqNiJDOYSkKAj7t67jwRQMcxylMb
zbm+GXQHUq+dMIV5A0afOuLvTnnJjaYB6/FAjPAplhBmtikwNS+rpj6d4MKkQT2tuKMR5+Z1HYWo
Ur5CDdFYpHDHccnACBCF3P6Wq+iS2a+q56Z1uoONbZkixXcXUJTG5jFLdEkhB4x7/PxiceupMLPd
Oy/qwVUMOeeaK7l/CeHKkl9vxpbirt01EcSA11LQ6ACPWDJ9r0EWSK6FgfI+13Pz60r+8iwvJ9r0
3ZpJPjeZUOjv2SOLrLDRoiwCrJ4aWqoIEShGC3lg5rnN6QfNKsAuntiunX84c0XMjfCHSG5gbuqx
HefzmXp3QFiS9dFq0xMlsuoevligKnIn9lA6QTaaRjHSGJat7q5Rf6Nu2y/z7+HyoVZzKaBflPj/
obTtze0qauwM5nmJ5P2o60esTKPv9eUqAvijOKyvLDQESAi4Frkk4Rp4K3wf1oYOZg71C1DuPR/F
+Ko9+VTYE5ppNDR2uZvRpdp+kV98jb7/SEFOgmZlFGLOMbll3duMAoKMDILqVMUk8y4qLz+vN/Kg
kTkN+6jOkxQcATRBdH2otBjVK83ZBH/Ni59mV02MdisMzUAnEe6HW1sQPchFHldhyl8giKjNcmBZ
wCrcuynotghr1AqViMcc9pfssQUv4W3lCinrapqXar42AQk2DXjms6hdWL17oQrNJso4NO92ZNUL
eWsJXH9HQz80MCCopjsH0T7z/vcXDyVyERiHuvoQgSndwpIXCYWNMIkQKhsCPFxPDJoCgXg1LWPb
38p47CClxSBqBcGX8yKQ5uIGIv6xW9p9sgW+gBSUSDnMBY3PqhITZyQ4pcf+wa23/OdBIJl96KVI
V67cTPlJ2pCq0E+cscuZu7KehHadWgeBKdnag1CX7B/aYBXKjRs+ltCCy1vTZRRIzl6ohq94hRp+
d/aZXivcJybrxHDJcnG2AqZPSiOb/f/ZUD5q/xrkDvPBXDE+FwoLnIB/Ohs8lCjDRCrYOeo5r1D2
A7Q5BGDfq1xLstfpoqEoYpC7oEHBSB+/eVvABStwv13tKtO3ax28ciXsw+jDqufmJm68JnLLLCiT
8S2ZZz0gCTcss5FH0QWVpt/F3Acjh/1fpqOtWoLZpCBtvqDEZuQeTyb2VXwP1WBcLptBgrun+hPL
5NRp2zRdpkSurdcF1sV6VDTgO1SEqcT+d6fBqKGqqOu0DpkdD+QUoHWp5/IEJJk/PJqSCxc2Tpql
ZHEnEnogs7jw7U6SsdcRK7nEdC1OffaQ/WcGAiGoTEUJGfFVFdawBDDoe0sHIsWiMq/Ce+AGg67I
oCpvsP0Q4Q1UvSyzb72HdWiXUqDgjVdeFMiQZ+kY6aqIKLr+UMaugjIq2B8dtN12K5pS7vuTHJk+
m3EplU/EGPJ22UNNKq7yBuNKubIVljfzxkhQtzXGSCa4l6xq4vNo83eZ3Q6wifmXaFGZoYsqufyR
fTQGkFYHk5IGtGpd6vbSz/lgPeZUFCzpfktT9h0Q5x/FuGx/6i2ums493wH8AEiHcVe0HCx8Zc/x
iDFyllaX6gK4zit6s4njtuHjH096dmMVwZR8rtxiNz89RG7JpbPoP9ZbBAcU5lIXY4398cHfp3oz
VnvVeWugCrHWQabZIwDSpWAXjUx7DNiiz8LL7HdAwMgPP22xG7GhF8k3W+4nDkhueTHX05e2JjW3
ouxyI35piSQqkoM+D9miYT0j6EaFOtJVT8qBcXBR2xxzMlON/uLuyn8sEs1WvOGJlTs/x7DlBBgf
ViAtP0HW7BZl3Icie/gG3Iia9zcFdsq7EDWnDF87829A24epPTlBBetczUnMkSgaixcoJmOqX2aW
PCk/v19CKTGrVwMkaxPYg6DElg2ekMNoyqm5laxm6GG7dhxl5xO3EgN50PIavq/AdZ8OKxjv2zFM
WSb+qwYayfbvi1QUHW/3K4gkyZflE+BxHXtjRfNBiQLr9Limf+W93EO2OQIs8yTCb9f4QYiBAiH5
VCXzoWZRrCeOczWRVEVMjqRpXO/RUUjrWLN7v3NAtO2tM/wkiTVeSLlVbGiCUvfAoskF0VN2ZkHm
VGzbvRQTVzfrCutTKICb6eyHq55os05+ZLvuzidOeNl4kXYpcb6vqFg7f85KTfPV4ciPBwX+ZwbI
SwpMerL/aEt0uExxyV7Meek2Ood/9qcR7fwlWhc3R20EEI/K1DhaN7hvb8EakyG3j0tsQrs37gAV
QYC8YtZgWRC9tABSwwLQ6ZgH1S0talpEYYqfxQjH5dTmr+LMZH0f1cZo/R48a+NhYshYLI1HvM3d
NGijdjBB7JvAGhckQmImQJQdSbswbBQvceR9ipjOIKvm/Jgn97L3x0uiSwehorPPvZ5D0W7luygG
Ao2RT7RQdSscaxgm+by6Ku5rFNe6gbW4t42VE5uCe4GKwUfIR3CULKIEkRMA1z7VFQOlU5D/mMMd
x7/MKpxHs3IlBJvNbvEjDplBl5ps0rJE9TA3twW1C+ZunjrngjZ9xUj2472AI1nSaPx3Qwo0sUFg
235F7vc3NSa6458sbU6n9OPME7sLDDE9KIPrXmXM2l8u6dsvHEGePpsS/5G51VhglBjgg+/IlsBO
VTjwrPaAi7vSW4Z65PnDKnQ4o8yB8oW5U9zWI8yiNMQmWpWvzhmras/FyYnIBiQaLQPaspvRkkM9
23fNNGF3/szNn2W5EwqjCMa1558pMIwLx3mL15uvvnYj3ana7cPqLCApxuLe1bQFGBaGMGG8wVVR
1r5VcUNHvL48mVOC3Air+gsv8X+yZsqZM1rIsIOaFfGnMrfPUr/pBdyjQlrukGtiEQusOMucW1zi
UGnnZ/hJxWyaXCuwEw1ha/UBacusrxKS+eDvO2+Iu2uvrkOvsJikcLrPnZLMBGIgCvUKem+nmTbd
odzRIBaKkmcYNuj4GmM/RjWOjfotD7qmGq1EkiOv4tLHHoT/j+LoZVXdNBUjvdV8x2WuJYwXwfnF
QsoRz/V1F/2Ju8gibcSDF+vTVcpchw/dE13RXTVS+uOY30II5082hI1R9gRts9Mv/H8/o7+mU9Y6
u2U8JT5xLQKJY3RqYMtyMN7R8UXunHP3MXDMdAhzP82LDJfb8YpgbKZ9w3K1R9GulCnSAl5YhApH
nCcb83ZAN6U8Q5++yoyHiIOt9grmGaZ361FtnN1916KnT+rPSJ2avyn4WkHZfxHuhjHWc0Sn5jcQ
XjuQdKvxma5tSJQ+FBfdvVFLmcUY0BLUrYGBYxBOdK6TCUGQqk0wIWQkmWG67YhevFtF5v6vmJnC
JRzju4CsWkXaBKP+s7ubIX02MwcvqRBZsinbZW0mWU1rvKISd1wBWI0SKxY00SELy7DB5kiiwF6a
Wv476e0eStXZBfA/ybrWYMGkVreq+kY+fBsHRHtQXUmJufi6AbmQaWKmni+2M6Mt30DeZeG+B5tu
kzdOjLigxlwZZ1cNmnVlY2C4XmRcuA5AT0DPtYUzfACJyhrKPYsmzkVnaLqdzeUfnkMLU5AuAotS
zcglZ2WTzJS+DzvKXaawoGaggy8psIoPDvpRLWe26+LtxSWU4o/+ipe9U7GTOQf8o68VeflVj47+
jD0XIefT5rtKLIZgfnq4M6J8lJ41ZmuLE7BlFnJwyVyt7gx8mWcTiHLDfeMfwUs4ajZsAvKuQRxz
DUuVUWIWLIycCGjyqJeiZU4kZarqECOh0F10trUk9HQrDu442RI9+jGp1OEmvlV2Rjc3HAw6xl1k
HOByNdOgP+PjtrwZQralzPWMwesq9rCdJxMsSjTwdamms9NnQsAdJk+/aCYWVs0vjYg7RZd+EinP
RG8Q/3hxtTWfqnR2txsT6J1CCVx63XRb6qyleFtVT2m7Vxsj1ediCAbap/YPOpv+0BKK/+SoOtI1
Y9rNerYKkc/pRNxoxCo1NhrrP0p2hsi4Hh9wpogkhvVULGMTaHekcczI8p4KgMgP39oOTLyqyPlU
mC8rn9tw2SRfiKeDNGVuUt7+NcwrJtcQGnmOrZbIeeh4Zp5xyohhos1mcpI/cLuRLt/UtU1+8RzY
N7Ek+EYhOo7SdISryQX5nkoNsGZ9RKOoGPUPlGn3oDm/3MtFWrrP1XTYnx1d54Z8Xq+lj6nPkll+
Bb7vy1fRhd1OoF4D8oLMMr07rLdhaIiBc/kCNjbh/yjU9ScmKc3cG05SWfTNkFPjDz+vcsj+Jra8
O4ysFUQ1J6vG14zsTfsLqZ9xH8TsLdNgxgRjde6m4MhRVxVgbug95DwkOE1NpUciI8e+PhCBAyUx
6W/arGyJBJjc7zs4yLWUZ2F5GdK5bYD131Mb5lnBM7hQDbgCTZZnDcWLHEP1B2VtxOHX/+pa28P4
yw9yPNgOjKyH5VKt05yAl+l4gnqzBCjwwS2H4bK0FT5qalsISC8UelqQ7pzvWtAAsrlJqZeL87ow
xFlIBkuGA7k0tkMwuYcqIrEQkLxR4sBwNKcMztq+RCqJAC7mCiNaik/mPGe+PsfcWJWMy14VzRiI
jM6WhhHF0rMMtUUc78wydTKeS8YPgPj8Juioi5+88iJd6s7s+XdTPJ5s+Rx3EumZJacxr6RvRuxX
9YTqF6j3iUg3bhrPkoEjdIpmVAmRr2IR7/LRR/sxpa4D6uFzVuOg8VJPZ5yhTaNiW/Pg9cqzvI85
x//YYq1Q4D8AdhCjML98K+B8l2NRpzanBA+CbOpW8TmbzWpm3F16703OYPD3D/fJQFjF9BbRUxB3
TIHThiIc0R/TnMdiunomkwPDM7+mddTo+Oi5OespITCZ+dFTnxjMzoh9h+UBEkgsHTHoXxJEaRwx
PdzyjCoUhSqQ8D61p5vpWQV2hF+cZT+wKLO+uk/aih2PiC+7I8jgTCxM4JwLOsZZRfPayNopV0I3
CNOugVU4ynLhOhyaW52cODFxBIgkJTDYVcoU0GjY08adpKrDJZJ7pwzdqPMtFo/fDTt6Tco+yYaI
rYLao1RxyTpbRNn4RdsR3ppWXsy7zqanCprGjySc1hJ/8vc+MaAbDy6n6d44Nna7722RSU6APSpw
LprS6DUydTjH95vVFUaYfYa5Pk7bJ3fpmYeYkq4bq0zkic5aW9LW64N40pAC9BhgA8fT9W+M+uY/
lmmw9PIN4ej126OurqXJ5ZaNF1S/ML1uG8iSy2sney7X5BG24oC+FSEVUwN4RLZuDsidIEqjRpPN
GM6TYjczpSOqlSjA2P6Orhe3qtm6ZyFl8WwF76XQGWzEnvxWVOqgVf53+gbFWuBbQwXJQAYi0OhZ
9A+SPk+VIzAh7PObjfz0R3ejije/LS9ztqGZuYxUyZ7icz5hEtKYCE/18mI+r9xgi0yQDkSKw3NZ
hXLpJA/uZB7sdncoTOfUg8TWNOpUKTFy7zJkT/4qMin9UNWRfnoFmhFrkrggsY8YGcoj/Iv4m74N
W9s1TLxtarJq9J5eQN2Q2FiLEGurA/G7mW9RznBzybCLHZhrK3TNvvD+D6FPtrjXZ4CR6sEddTkO
A4Z70V0RpxPzb9g9+ROxNHPZ+50svU8ImL5zc1JST6sT7M9JMr6j01dj5qU+CQ7eR/6Uv0HZyBwI
FHqfmhP8+ruLWzhEU6/1Z6rT/0auXP762m3krfJ5ZOAqZnfnEIf+IWXo1n2nVLKys3eDy9StTuBZ
+AtlI/ECBdvUhDiKQALy440289kOg306QV7aRcQneFqN7Afs7NbDzIGggjCk4aYUrBJM+ykGcjaZ
qj629PsZyaZNakzWXU5GXBpqociNcldHaaxzE5xDu7Acwy+zsGesdEQXSSd118BBIJFTgeOzREEn
6G9y2+M0ASkEffks10VJrlCfHiQCFgz0Yp3GiT2Oxi+TslhV4tRELqSfOChjhDfOdztMyjsvQhK1
27QaeZK2jqeXtHwaKPqrQpGr+VIr4VivCTOYcznKv8nzmb7xdER6sIhLsbBoAOhrpYJMfg/bySkJ
lGXSxvMA5AFyffTOOue6pTbinSq5wdGLxtSV0LwdZARwV9viML2PMIayvICWgz3apFu47Ap8smnr
kT1QenLbAr92nlei1rCFamp2n/cWWv7VWr9Bm3uhv2M7JfrucLoRRJdNf4wHyoyiPnl3AfPQTPb0
w7bhxP9Vq14whMtgYJCedQJQCxllVp0RhnDh+uC84OGZqculqGJlW58txnRmEjfn02iRrTUweXkP
ruBhoLWpBmDtdWQiy313RIzXLiPL/1ZKzpGTnxXnrxkNr/jSgKgZRSJoFcEeqWbNFpeB8+fIF1gm
vqyaqht7W8z+XVutVektL5qOESaHbf6/tT+wApHh1HHqZpJpOww18bstau3TOfwAjfiZt4vcxjQy
u0S2V51nCI5Mr2tN3rEvkzlQqB7vP+PmWJZhcKUWo9MISHc17IZ5A/URJSmQGbQu3U2zxZS120pw
Q+2QSUwH8vnSl+B76ScYGEa9msws01JhQH0XLPoCvIHU3Rle6AkEp1lCfRmbTgqZqp+nlobGBRJl
58c5h6artdnHBfH5jjggKaLb2+Eh2uVm+3a7g1lxL8HJcqZt7JZ1RYyxU9zqO4ktNLjM8q6kxBW0
0yAq91y8GHEWp36drb0Se82uT6jDW6lYqjiyuqBBWwYuD2XRDMmNwf15ofc3IpaxKM3yzdIoyQ9D
Q0FwgRly6Pa9bEnN+QeJ2m4Gk3HTsZHnYDLgzKQQ5wD33L2PdS8viBb9mBwJOcj15dqsHB5VFxU5
OYaph1gMgrEynNlag9ExZpBgbJ40ur0XckB/KF+Sn2OJm5WjzFC/anEI5PX77WoZFTWY0GWiadWr
XKzK+zScnqDBeiB/m70EwjmhZ1+GjNM3zM1YV09WY2YCA0ED8dPQFSePgDihMZJD41W5+nuljgjJ
C1Vnoxxl2iw7AAt4/3l+hC1FmOSfrCoaxhrmnLoOCAkLuCwvaST/J9/Z2NAu0TcejmeI8QXmuLQK
cuL5s9EPnetI1YqjRhUZW1NC74h02NUR4azIy/+TcJiZByaTAKP7xUcNCVbD3duZ+6QdKUShRogD
RiQOQ3ux23rsz5LIwRKTf6c/WkWgdoffnVL6HRQUaSUgTfOTOCaXZzuOfXawRvSwdkGD0MCgZ1pF
/ss4WESSIQhBql0uV9YY9/x2oKlrjyIe0YFc9FMl0LgOwhqFCdv3ho1puP1zw/I9qZMneYyYEwkp
6eWRDFaAAhGE1GObqzC4IwHcbtPPaD/BZTwXeKjQGUNJWHubgmQXb2WBUxjVyXYTmuX8H12OW55Y
45hfEQ8TnX4bC3zzd5LjEDt9/EDnKf9IyY6cDvMGY+GqcDIRNYo8eOGfcIdfM95RSJUqu0b4AI3j
DouxK7vjgFBkufu+XKpjPh8COPga23KVCMcg9gxvQ+X2CLdGJrOmBvDngE0yvSJSCItL6rttkdxa
fl8pFqaurCkQ5SyJoFz9OymvvkUxbtotNNOxiBPviWepqTevQHWNAOeEtN9aNTstEm20odlKpcFt
2BnT/jOkeNH7S4G/WGFSWw70aDHJlIGdfeNJabINZOFwGfheAHJqAcxIfp4tTLYvq0FW9dJIWW0Q
5liNazjmcS4gpuumwaonkcWBNAbV4wzR9eRVxqnIfhzFmnc7kmJ5qLEPifz3rKHVSZoclXB7ckqs
k/m1L7rHLASqJ5V/gfxe21fwf/qja07qFtK9azWRBN4Ve8OLiuVNjR00brVk6G9HZxEu3XVdxexe
dCDKkKJ5JvLGgpPBprxXqBBkrLwOkT6oyBZ0zbdXJdLhJAdcBl5NAYDG4HF4Dk3Ct0YsWr2EtLpY
6//BPi2LmEdTlS6l0oUK6jxmmK9alKed5cSw5tJOTz1q1LNN4tDUCcNXt7cOVrnb3YPtyc+Sw8HY
uijlN5n/1KCJaVj6mkP/XSheexz5FJNDjmRGnyhjNoFRlWvbYcZJwTvy0hQXlw4QhIYCWZ8IRZGS
7IdZ0a9FqsCdOjfiFIqWRQH6FEpT2rfzVtIuzwW813X/bOck60ohsrAeAJsHPhsDzfMjJKsU4CFM
qemwUJ4s02crI4zNIjMx/GBu7Q+DgVVhE3PDTxelyxH/X0TCX7YBQhKvpYEi7rwncr0+tkSF2VPU
DVAUCpZO0YMKOY5ByMfuxqvqwpHKbBkGmp/FWNm7wXkz0N6PGBydeftTttfbW4IZUKLMug9HqF8A
rwSoyF2cJ4o6xzbJ4px/9piZFhg8pHACq9cqtXDYH3aXfQ0t7lmppGs6oEQL6iC9ys2YQEdTKTgx
SNIsErzZirez7xxMCdjyIGzVXjDePT5e2cb3cAFXNe6+IZYe46LXlHUOijjUWDWboz16GpTBNE7P
daimYHeP21OYULPnxDwaoXcM15FHMpE/ltHp/MqykVBrQYxH62QqljvsNcm7lhMT6y6nJcxLINK5
4gpM0Me04cSmMgxEZqlTiKlGE/u4Fl+Mh/nOKf65Qkt1xuOr7y6jegTEiciKFTMrz3BZx0eHpnZo
6RMBOL3bO5dboj57iz7rvPDgt0l/S1Cm/yg1NuNVf/mCK8Ut1JIVni3tTNgqGX9htxAYt+HK6lG7
8v41pZoMA0SDmn5UU2FBCtv+47g/8tt4bbCJMXdDUra54XraDWxjm8CMGl6NN22pJldHvpGlZlMQ
5n4LBGCvBjrBLIvcTUve6OvuVCBs0t93onm7B5c8P49ynnhcp4Vkb2L9s/4UWOMYX+PI6FzXw43X
FxpqUVmA8qPg4fIaTeWODt1/f7HqsJqwAfA8mxAmfxsT9Fy7m5l32obSw+ve+PPIyf0yhWAPoWXU
ks4OVtakBiFSNgb93ZLLZ8NOCI75hIL/c4WS/UXToKcvThK+YYHoec6iyt1Kp925IjSUR/hwdXan
opBdOE7lkngMRLj88dkz3AWTnIiBXwi+eidzE49+tGxj4TvYF0IdFfubUmwZ6OorGOxpybhTmaWC
OP1MNjP7hkFdppPmXp1HFpcjhAGEQxNvoO8SeU9WZ0shEaxTrDe4H0omlfIWHB3IP348Dh5t+pab
YOn9SUEHRV9CRa2+n9osoguCZXlJ1w6zQIvgjzgWgub/6amGf8BUBvzbG5So6Dy3ZKqzXJmLaHPV
BlCSbHqYphUe7Tqe+NCjgVAlAqtU1Sc1ekNWRau4vRLvsTpgqDjygjsMLijTdfPt0gYoYyiokxKi
vqCxT9pdikDhlp1sRwVHTm5P7tfXtKCIWxkshzNeCe+oiI6gpUMipnMtSmpBhzlPuB//qZPubZfm
1IAqO5nsso7uCI2CSnZeR2Z9KPJY0MF5DWSmwlNzWk5zEJsqlpimN+AZY393ZuphgQ0rdp+hddyg
tIbzMY7nWbJGIHGQ3fFOTQBG4ni/d7biEFT+wMX34j+HFkdNCSfP+yJXbBpKNQwgwZbbb//Qs83a
xnNrZAuRLYBfZbd6QiQXSVzAhPKVf6YCA/Hsz+gKknSXdyMSgIzC6vfzYlU/hV+WBchm3fpAUrZ+
dDJgnU65LsjqMYX57M/V2eJ0IWoudXVv4gEKGqwBrctzggZ/DVlfYgHoy0dQCNKvXKe1F/5Qvo9u
3YzFIN00oGKmRsD/6vFT2TUzrNrLxI9B7xMTNgdKm7xf/m1tjHh8ZGGTcEAF1lzA5lsEj6LlA2WW
JY+f3CM1lS2WVsqAG8YAM7nzH/n1dvd1Y/ZVYykoDKknzMoNlcHqnmB+i1sYf2fn1NqwChqtlU17
t9G61uVgYAsxq7Fcr96xSE+FmEAv4G4RBJfJHBdhfB1GL/b7q9q65eWE3cke0dfsK6bIYa5QhVUW
ghiCz11rXgLP5OYrVcre83xGkyDM5vvcBoArsWtrvqokG2X4AFCTmm4Ej/D5lmos71SCsseEj+kt
Kp3a79ZLLvgQgV1d1p7LaZGoxP2dofg6zW0pTVo7mm/pjD6aOVvK5C+cN2hw+40kCwnQGUtEcg5w
kdaSyA2tkoQ902irhcgHqDsgwLuN4q4G+aSe96LzhErw0lqktfD0CFkRQ6fZGxBH5pdLx7izeE95
fgUGf3hGJtY1JLYzcWOMuaE6aFxsGv30yoqkbRyO8k70GwZwvcrPOel88CKPPK49MD05q/z2W1G/
01ZMIlIgfCRKy+e+eeCtTTOT54dUMF98v+vDq8s+bSLGsbyTGxsNf5gFgeiGatujObAUJhXjoBzj
Pxthfv+SxwyV7FaBP7nPpQ2Qr7+fi/E6Lps2hKJxIje7mgGK8oT8NdYNeh/35rh+lqJAkcRR0pGd
W9TX9O+/FFNkprajAcTiNnnbj5Rdh+0dWlPjjfhmG8PC1nFFXOHoeHXF+m6hlhGHJtNGHFyfihmC
fDnNMEYZGtLeY7YR+Tr+5A51YHCmi9h9t2qaiCZR1ZwXk7vCklV+AtAp9FxwZY7jrjRtykwASbXa
jpYqTtrDgyoEJefqyqL63H4tAfev+oPQYpAtTSrCUNlFfHLq1/s4G/spwYJI18GFDy6lfzfd0bR/
y/xeLXRPNAX24X26d1Z3c9fDyig24Q4QbiqOgxMuC0yeaabfLPuRvw3uTT3MCfWfUNHphP6TUnnz
jaftSpSSZNlAYqnjKmXWhDKJVxmxEcSvuy3snJotB15p1bwYmfc7HIB/YQhiqAlLt9vgAViK7ibO
LGxrQAakXnsoeuTH+m7HRuqZNSrlLcIrBy1bFWzeSeTuMafDINBRypCGj2fCPXpxqD3S3XGNFw5x
Yke9btveuCC/0Fn/3kV4y5dpzSs2IzgBkwyjmby+C6YEhx2tAyhbfhKZjNGo0yO6WQb/2KpWEM90
iwqf2vvzgD/3l5Br1PsgpVV8w+pxrs1PIq7WofyPsb5EYWESro78SKsp1Fz2yROmVIke463MGkjs
qzYaVfB+KHInODqxCfoIKJSN1Cqd5Ib7fJXJ2s7Ymwc9sn+MZPRbGaA87Ruz6CREfdQOqBRE2mTt
InuyD2EbJFCcLJsLN2qegBcQ6/XzsyntHY/ihybgcmtrNDVcW53J4hal1RAqNMC1FuPVhPspXn9x
TbjbNIN2yE8FzhDga8Y4biWHght24tfxIWjbI7UQHaB/QrNYXDlLrd0tLrOsXBd8ewtzOzTI9zuF
AkNRIbUbvhqMuvzCTrdKzuq36nWBrlqtvBTdGkehU5/jRTo9GM3yL3b7PUA2FBx+HY0hMWyE+xqO
hqw0/F+KID0pS4TwNEXHi6j5iHJXetHGKNzgyEYTF/XuwehIp6fQD6CwQchr9IHzu8gj8VuwRvWo
9rzmXPxji/CduWyWDtMGUPSJKITuqOviHfL9TG7OQ3XzEvqDww+6t+3M3JjrJMErtX1lzQZ97K8s
eBQkvWgnkjyMkf4NMu3yo9yzWrmO4X/z6l5KN36zSgmU/8VeVFiDtFQgcrEjhbJ3zrhV361yBq0V
7LNzQiyAlpSl3HZbJ4ZXdrYNkA8/hLOjj87uuHDjzRPZN0oX1YSjpAZL/E3qhjL9Fsbtga3H2OqE
mqKyYbRVJqGaQmXg4V2jiD+DG59eb4dzcnfv71OvL44bjRr0REs12HwyVQayEjgSKkpFH4941E/J
np7J2TlcYNBRJCVHkAOaEgxc4y8sGiaSP54Z7THfn5y2kfK9bVr1dmNKY8cBc7KRk6xj3zXVwRj/
g1M0ROSu6vMr31lKBpS5iMUEbSdTpGeeoL4zfpUKm9IVksFvT36JV+/0bAHba4ljeYxv0xnZ9CPE
oHzGPJ15QeanIRdXSBJ54GfGJDecUZUP1n51HSSB8rhEEntc11BhdAdEhiIUztyVFRMjRHFwsZt4
sILzQRUgIdzXNukrlm/jMCOJ7b8z1b+nGmWkvXWO08kstxwPbws7bnZtBi+UcBz3+S/selG/v6xY
cWhjP+20Tfx5+QyBIAjFB/a5BlA6KOEB6a564TKiaNTCSsSMrJPl2qQn7DCvea9TXWUB3Q1c6DG7
XAcjtttepbUJ6/GwvAshVJMHYVv2ra0S19pte8YZfRX3gN6shWZS7SOFHCqFh3gsDaAE/++Ie+Ne
BlGVSHCTY6FTtA2R2FgwolFUB6o3uOT9rH66AsUkZSeCq91LdjGHro0UjvcfvLQ7MhyIxUMr+ECe
jmOkJdvlnDZ3DDWArFktXwt5l2zzqAqJOV7reyRnyXhn3JKr9HaeguggD0bC4IpVgHsWRRhXJfmF
gZvLZJGCV/2eD5q5PmnDyg7vhl2COOOf2n3szoPeRNXWjiB82mv5RpRLgPAws0P/2Nbxpsryn6BQ
V8Gbg0+PB2ieM9idDxgUTME4YlaXAi9DdP8lIYkbd/DvS2XmJ8rfbY73xLCDDv4hTmIcdLLkqLEw
1v10WmdU0ywAtZvu0B6yVvs0XxY/FlaWTQriWMfq5AXhEj1TsQ8Z2ku6inCEWTzEOrTn5RbCrvFM
1ZR3IrEzDhSv8SgxkdXwmpCLMl1N0/IJC9VThc0H9gqlRtdXBzCagUTJiNnLu+3kYq0ugoENB9gO
sbdLqXZTlDq3nlpYafYNalV9giwvJdtmLTt++KhXMgETMLNdZ9x7kwZ0Jyxa2PjBZSNR9XK6uZZv
zdl1oz/3/sMNiHwVrbmoPJd3N3yMnWVzO6fQh3CkTJTvSgbcDUGoo1HHu4lM7i05hbLqZTCPlxr7
eGBWVexTg5gvnY2QTbM/GzeXE8K2b3eHp+6kayqGnwRq47n54lgIdd/dnrM3gwcLLeuyWFwOghWW
iyFIqH76jPj1PbDQrO1N74546QYWDG+bhZbodRmC7piyzpcBl7lPL8PzuENsjAd3Mj41LQf7oJFm
RhgZHx+cmhYU0lkPn4R1IfB9VvWn/EUBlO5Gn8Ty2bUIDTb4KN8FWcd3XzbM0XKBFax3Tl7V0WNs
kMCS8BhVxREuqDvTV68ZYtOOF1v5W651mRkORJ6Lg/9Kepi0hx5yIXdqmlETCJEVEaYefimge/zI
Aoy5yXxf+fJZJu6dlLndLiojUwkf0vol1Tswzqco9PqRrAxaQRExGJXK4Ny81JyKgWRl/S2a8TTx
BfzPAAyIlw6rPYSuPS/wK8teNI8dkvs0QHBXIq0M6Svahyom+Ilt9o5WebUxKKJOnaHg0XfWWBPy
QUqOAhaA/Dpiq92yqpxePve1NgI70yVHreynIGa4qdotrdKaCbgVW+bjlNnRVDjCWS3+pGHFL0Oy
72rz+kcV4JY3g5nlwQbvAKIG+9s9oY/9j0XCDUtHYEH+ZC3NaauZo8rgpFa7UodahWGlKNZrRfS4
GltUnJxeYrzmUEAMC8lLbCNUHJDIj7Mx679SbXUvoYDAvn6X68Lmj+4tp5fWblU4yQHCM3PL4fV4
qh/rWxQAL+J7+b1i65pG7h9805prGFeW0OeDLRBC5XRbCce8NI2qVAlIGjK98bxhmRf+Oc65QG2b
mUEbUG9/7fcjzfNRz84tJIShjG7YzTaiwmRBBoY+f5IVzkLUYLhjsIP8Q3xZQenJwrAFadqIIYt+
5FPbxRGt+kHe5oqfsM8upMmNA7OpAqsjfwp+G1jRMjq42FnNQ9bBZLKqsPRUbCqS/fiewVlgwTMv
Jhyus5VNHfaI29LdFkd6M2Oega3Kw18mmE6p0j+X6vMKvGXbWGJ6IoWcmGUCkUdWF/PwIf3ABUBo
65LTqIM/c2uoVLjrzjtfbU0zPmUwEZR3LBhv02lyLn5PZawEO8Et7geBaNQQsxsE34L4USHqRqXA
mut4TFRM6XGCvNmjNu+2J2zXWiR3bL3oMY8IKyg1cUhGwOrX0dx4E3u0UwZUSzwd1ddEj1ormc3m
ZGu/3qJydXWO8X0MTgNxAH3z3KeChcP47XwN2mlYMdeE+VHxN9IjxsdlHBAHqhdVCn6CAWKqAJvB
tH3WMxZsMQJWjhdK/HeZTefU4AVDWMc1kjcTzT3BvlsH2jOunKrBy/mtazBYGZyabUUe7hFMXPXJ
GDIBzkZL++lDqavwnHDSCyd32Tfz/trUZAdMsq0xfIxaClFDM+WefDsKNP5Z+DQ8D5/w2q85CIIW
+jIUMJyo/1gzldDFkqFO8VcR7YTqXPZrh4iAKKeBJmmhoJsfg3kFa4cdbcsYM6iU2chrIGkJGJoV
vEnPszmw260UdM8a1y4vQgp/S91nIlHfXDdQtQH4gH/nscs0kYWG7XkrzlaJ0GFPBzt/nwAVnqXw
py+R8iMk+yNpoiMoNpCdN0eOdbzThBrGpHqRsqcaiDgsEnRCZDpgUp1/5xsSPsbDLuDjYwGEy74C
dzGvEC0+Lc3rm36ASgzcDnqaxIA/zblC5dwf+xf4rSc+lPxqK+phw493k0t6ih5SyvXETWV6G+Cw
J62wfarJ89XbhLr0YlwavhjLSuWIjY0z8jnMPWjfoGjWVJ27ZOwv6UpE4ADQOE3OrARI8U7l3qQ0
sqdZ7mhgJdnQnKRTcWdxEYYnj4fMfmIwzmmUKiG4vjPqwCQfs6BGdhkj23IYPwm0Flaxq7N9UiDO
5DbScQKZF/VkLvkUdVcjWhPphNRmxXqZtZLHi5FE4QSVb/erp+BW4dwEc5Rro3we/2uvXpahJBZS
fuAiViO8qLTl/5bcvDMg4zNQ11I9Wjm8j/WY1V4zTsVivlzpbraRSFen5g+aaVHXc9Ai/WhTXNdE
uNIjFGh6nzSIQLQxA9uKDYIyonLzDrgiFbQylQW4RoKbM8moafpigITX0CKxJJl6W097zZnC9bUe
/BRMu61/RNb5a6eWMf7IAaBSSDBsmwfHnHccPzTSts2Kmn7TfxkASfZCcCF58s2djh0XLaCTW8dN
gDmHE8DqRIoP2r+QQc+OOQ8oihZ45Ac0v/siKaswLWOUE4YM1HcyfPIFMLiK04RQbsy2TFo4uvOv
sr+mHdQyUxkzkfxN+hYUtTJEjrSYOSKgeSMlisMWJCG8mxfurXXmuKshrnOPn8BZBNjlT99YPUNV
SfMpsZImri35Zh1m+HOgcHQA1I4CKWnNzkBGPCBWjbVyRAWDFqfwwm4A4NWNAevjAVQR16n8FQaM
y2woFWmrEZc1ttjwzwmXFxgVkUnsy7K2JdZukdfPyKWoA7zR70Sdh6GkvpEEqqT2hNM5jUHVPXGU
8ESL2/IRgZqVinp99+wCkXge7q1pzCabiW7z2/GH+1ZnQe9UVxV/6epvoq3bMicdTWof/jtf9iwd
uPPCfFj2SPcWl0uA6eG7+PylUgSI5iOZo56J8e+409dIM05lpmqQFG1ifWWgmSXdvX824x8mgRQ+
OwXNh0HMhPiNU9DiQhv9p8OtZ+V32HpzSmYMVUhsx7+oxn4qKjhNJ/sw93L+5wtUa4d++D4M9WFh
xC3J8Hcj8drv/lsfViH8FqU6pwEW+1czO9UfhgWG+D6N6jAYVWIOWdefIQvGO75Bjof/WtJDxye/
15+Qcyb7c64GRa0CCLciee6uvGMtHrxDQ+mDMPAXmU3jrDJamHHLk5FMfHjAnzjOiaF978efpYDG
vsXngqWF2WT51csvUoXxv1ekPsGRGPo2T2KkzIiz+I9L36Lp/QvDL1D5PWilaCxQnEegDk3JLaJ8
926DEjLl8h7UyqJBODpIEmyTVru1SotnqWOEuJBleLKpWrp0+QTopyjLXwdrPCd/+EY5ecmsNij5
9JsOFt/8rI+ZzHY4b624ZbSYlPLfAlXo0w5CIFFzLOxg6m/c8ap32zVbtJx4N9VYszfliTkUFYBI
r9W6sG26xFiyzOL3sdW6jWCInkWADXoJ89AIXzM9iNv8OaurZNiy9tSk/ApiSs1rdR1MK2dYfQ5A
qdbmTo+7ntZCqSrUfWoXs9KsqThkDpNwLc8RTrivvFePU6dXPPdZ0HtasZfTe2LuNe2zOm/i0pZ0
GvDlWfvwLoQ79u7bOIK3cw540hHMTf4Sl5R7KLx1XRZShBX8vrI4lzomnHx+ZZjl7+24nDYy/vxx
O02KMnuYA97RjNszTGeDh+AFdIWz/ZsRDTdgSG1KiavFX2V5lQDu7WSAERDu5BQl66bwPzH29OVV
q1r6vgEfpB4HUmRBZ1q3XSH7lGj5CMK35OmK66NIrhO0GoVxC4/LAUfZRSV639YyeQuAknMUhjVB
CXfn9Q9EsK9wFa1b64XpMJpdvbi1cDJDISaoJcrfq2Cm6oZ6fAdD672ldK6QL53jofVSAM7hlGm5
rJRBHL2eWIZtS4OEQ6LwCK6OjaauIgFbJpk5fhzAu04A6VXs0yNmpJ/wSQVdCu9gL+Tapm05MVSZ
XHTVwpXsjZCHdUw2FOw2rKIsoL6NduGCWw5Jsa0VWzWFHguTmhbYK5gz5FcyvTGau6/4mtDP9ccV
1rg5Iz1TnDzTrcm9JhoNjkcVuGw59RCG5/iNEeKpDdJJweocdYfhJ/vgqwshKBxAKqcI+GCdxUPi
VBXU2wj9aPxCr4rMb+SbfG1kgbHQmO+8pws2W00beEqGSRXT86aZirKBfY/LVUpm3D//D9lsxoYT
9w+3C2c/6AFQWAoC4lz9e88s7f96gvHZhlnPW2wwMPPHKFv4gwa/OlgpzLjbAshUI0PWEhqTmTND
M7XGGFC+tCdym0ueea+D/r/svKqb/P1a4hPAt6B5houuH0bDYUDWuIb2JZRjON3d6TUi9Ky1t58S
IBmbyS0f8pvjYykgG1i6OR+B3QO9Kiptma9z+d7qHwkqhwWDIwxoYVXgl/T8B+dpJcU3wg0ClMbg
oCUwQX9IkT998hXzb/3IeiNCwS70dMROsubPwfYmjME9Ac1Olg7lAXk75WrJ/q/yEVVcYMtRmAVx
byiAYKAgMuSFmi3GqHDgwj4148uJJA+GXJXfkDCPH1LyFplSqedg76lFw4yeaq3FL6+FCid1JlEb
h+gRRARtQIWvP0AUhHatxsYBacXY5HvHQCtIwfLf5h4vaA7uVjh8SAIWBwkuG5iaaU6FFed9E29/
Almj/J9bZ9Gm7P7FFq8SHMwsQ9Chs2QONWJ0JLXOGoqh9dxwnTDtBwSRSxPa2aORbVQwUeA0i3T6
tBqvfVsrcJZI3QDtQk1kjzen22mhFkuKhqarE5mf5+EXZdFp0UVmcLZeaK2hamaR4YbRa/OHKVMs
5wut3f3amseZxY/0hmz+qZHgX96IUTxrSe0Nv/GnYOFIEa/uqN/FXZMPComupcXU4J7ro3vNVlJZ
WejHHxW7qzjcAN9yS2t8IilHpLMnfZ0B071jOToRMYsyqTFQua6NZF0MrnFLngE/kji116x/zqgR
JnmlYoTNQnKyrdIG3e6PVSpoyVM5vSUaKvZOGHtYeEcLtg84Q9K7bE3vDERj/D+lrbI4yxSyOd6h
oaPkUWkbDdFkjJBL49N9r2pqeiwGI+1CVwATWMhOLZByYjz+mRBXUWKwNZdFFM9BG/Nz5UmhfEqw
2b1lX0bQz7DhYRObOvDStBuFe2pen+xkPrZb8rM+rMM7+h8aETABF/oYeoIRkt6dinoSOlNE7Z7k
Yj57i6E70Q4u48dCvyeBvDl2/3tXur8m/ZO9IoR07pI8TxO0dJHlN2hXM8HLTaa6A8iBPh7z8Jil
DMyTjACqAS2G6NAcmVs5TDOHaJLOa5p5hTA11S/uukOg0GezycezNhx8q42cSiMNkxDoPwDz81hg
vz45EFFw4uP2Se8PbIFNqhUY6e1JM04oNn7AavKwZy5Vyhxfg7IPykS8c4dG6jVp2TAGLTrn5PXV
jPQvk9KrNofoJ4OTXXi8lkmQlNdbXVKU++cgf3kIZdLfaR2qw3QnSmtlps94ENAAvMorAwr9E13w
a6DQTLEWhge4b/GHY7DXac1JI85is8VMKORebrLByhFiAC5SmMasM6Byt60YFuKSbE5QJitHDeg8
OIhLx/cXdnkcLvtA8JuKfPioI0QdGS8AxAXh+fQfXoeQqj0tyH7ted47Bkpj5b8nM5uHpUsY5cmr
1QgFQKWMo8ydw9bwpRVSEv8Z79a33gVC+I4XqDhoIw9romZC/8XILL/e1RG3OYNlR3DnRTiawSh0
UxJC7EXV5fbuWKROan97CDEgGG0ObZ6vSwJpMPB8KcRmqSnthDeEqcZLo1vg1XvmDjKkU94DcUBg
6dQRu88OY9n5rmS9qc26Uoq6vuivJBsDcuXgns4+IWTztCSyWaFtLk6ayPTb50+2X+jx2bP5/CiW
9+p4Gz+FTLrhArdmXnnXesAe7GjujrzLEOR6agK3Ml3UVtPdaJ16ty4uA49xEy8VJvBzTBwKn+bh
URKgPDmfspNUVGfbAfE38MDvbro9TKrtLj5frkNh3c4ZdU3mVTCG6yf6a5KwYxetz8lhIBnkj5l7
8Edw5dV+vXZ2UM2PZziz3KHBjJjTELyrUEPLLL3xCCq87Wpma2qnqBhJZSWb2T4Lykc8NbutCVka
qIDc9U3stGM21fqX2B8MttReSVmMBBrAGqbpz5IJpDbIWaubrjdvbcqE89Vht2wWSINEXhy/QxIV
v9nZDDJJuicp4F/YLUAlvfz1QnPT9Bec2fUpkMCGE5xFzI3uRcMxQYrQV4NYUNYPi0RpMl5wWTFh
tA8Hi0XlwTdaafvQc9rIwRRevUCQRO4cCHp9In9c6JiPXJXJZhsDxF8Av2zYlwq08RG/vfxhjIUU
wqPjhjn+gzS5KQNXOJtYkAJJqKbCYsjua6VwHJTxTg4PCzFfNTWnlNZ2k5Mf6vBCuiKSoNFtGAZE
2XYkiQqXgYAV5TGDYvZPbNaJJ6qBB5To+hESTAKs15Tu1IKBUAPQUOyCh12Cj3o3n2zSuccdQ7Ry
aAr6ldpn0HGon85b3bkbvP2vXME+Gjnbd5dJikZQfLQ1kaPqhOFXSeOHqficnN7NC4oLd8nRq50k
pPX3TwrAXpImZucbjhDuwpe+scsNFXMjieLvBVRUKZyik1FVc927+eQO/BcG0+WxHzZM+2VEZDZ0
9IrmJ4x87Xpf0vbHWfJz5AN3qZ8CbKULgPS4SERTLJpu7oRu6Rt2nFw35AJcADu9dx+5qt5nyTyI
Gza/wu5eoLv/l86UWmdykh1WoICM1b+8RnpIJy3mnbw3ASYANEKw4H91zET6IIJHJi+A2JzpQHvA
DuH8aPcBkO1ikMtkwlmvqb0EG0iVOKWIGfKk24WjKi+T0cPQkBSvTT16O+5iKrehWov9sg5uxIjr
ImF5aK93zs+gHjVmTVGnBi4vngZ+/oayPGWLtQgomUzGfcxykBuj00+FRvhlesxeFg6LofZkLNkE
67D95ZnSj313Sd5pFzUvCIa2KhpxPh4uLt8D0wwzHOTgdaWdlRYi5TEphWFtKIgGTkX8ll4cTrnc
pswuZNweaCzsYnqUfVRuDyqX5w1OZfJzmSUktPqdxmRXcs2kLcuMsAo9tu4eQbf9C4x/QosSeBnf
CbbQGNMAyo+5o3j3qbw6EQJY9WqvkGrplQZ8U4v5Cw982kYZwAuXoCrxbcBnbU4KWSSSkxLjCEia
iDVDWHSkOhOciuH7D9q1V70SLtC4XmGP7bB7WgAr6hguSvCiuqyjeqLHe6RP5dgcT5zVPAaHwlZW
xcCEgSbEwpJYZum2cduvt81KO7pa03358kBHVfVDlYCHjR6YVZ5PQGao2sNCR188iz02iehRdAxr
A4PRCMGTbaEu91Y5JcxdSLz0byKrQBCl25Lo7LQfng5j+42RaCoRlp8iv+pUQGBTBOJFZXmvhwuT
LJfOlUCESvUwdFdvcT9oNeSgMNeYWlk5aQwltkLVnPsP6K/eWOkLK1t5NuRmk84NhGVyvdNvSxQZ
8lCSKVgdT6Yq6znOMO4xqPOPuD07DIXlyjfYNp5Dfi8a622Gnr4o83nPWfEKVnYgzqXstUjC+0/9
hQluV0oqe6/9qd9Eb5jTmrwMfz3AlzOCSaYyXnWTDu3+7KoYvtSIdgFNvpDGMUeGSJEB/5fXlCKj
1nK48Mf9kVXhisaEfmlFHCKNLPErDuLoKFYEsPClOggMoOrKgfsvnu3xwOG9/g2AoHHooRT9wvRJ
eVRQ0rDyDXCYQjivMqZ4e1om2XDRjNL5LER9I7fQ5051hoUtSCzSFbohTuSNR6AxSAqUgYPkm754
iub7PJzMF/uOgNKsktf4J+c5IrT72yidoUEWwvS8H/7dZ6Yh5OoLLQsHvhROSkbjb0nUO+33cvd9
Bu2eNnEEeO1G5x/vvLRpXigwaQ/00nZAg0MM4bYOXNgmoKozruy+ywDbOXxXnuU4s8Kn7BbjhYNb
NthlmOn1tAh8iBxGz7K8nk3xCFkfOWHk8WA7/vyVJfbywm8g1ojNzdmPm3Q4WDWYApb/pikG9vAK
5dA+7Puz25xqtyM0ud8e3WN805nJ/LnvGnXmeHwHqyXoPGRC+HqOhtFUMgg1zXMTEZqSCQjjVh+X
beaddzZ0lPUwj2UUTI9gELZKpX2W8uXO13C8KEdqI1HrUE08MhKsUU+WKuu9adlJkv4EE8KNhcx0
htkzKxQ1dXK0HvRuMzYtvY8xZw2CE9AZDo4N2ywLyHYD6duCmocxIPE5nuLc46+kOYDYKz2aoSsZ
Bf7e6Nyp0z7uBSM4MuRItcf+d+0pdrJuVPVuBxdNVkLLuiFMtXpjBLAe/9hG1MBs1SP/2xHEDU8j
OE5db3gIIy/X5fn/HUreeDQhZRV+FmDwCBnLm5ip3rpzVvxkUceSkBev9E3iBt/nyoXThPXsSqAp
aiM/zpJgAaBL5bpt3EvGB/80OHx6tDGgP8GC2aH3Hxy/qzxRtiIztAfX2O0ZFzeAW0ClakPcjYaV
HfmUkyJNYO00mpcc+P7crP6Q74zR+HZdNXppxIa5IX7eDPFETsHJWK8OL2CIXwYRfTH5vuND6S0O
3csbX8EItG9gAHsi9FOMmLSQrsppNOmQGMmyzojN/afeahMP4nbxYWICiIhzLiX5lx5Cs0UPGRIq
47Z0f6UIIoTDWyJZe03Enxi2a+i0kBJQEZF8y/tLjYlfYp+BJASF/JHcyjF+IGjHv7WDOsE9klyH
7EQlTdzH3pcvzcDe47kEh59yBAKhO0SQ4seITBsyMrd67b38XxNulBuqlHmjitdlQO1RuCb1UNqB
ZI2PyTfN1R4q78RGJPyVoXmHcoIsMINqBQGD2/hYnLWbIHDQPrx4fOVo1aAHJEN7uNPo5eukcUJ3
9XRbrA7RC7K8dfSopq37rbmR085/hrJVN0ZHdyGNfjsK33yJ7K71a0sla6E9SN+XyVZ5BxAi/sIG
hC8X1S71b/DJmxfloEzAQoDHi132ZkjozjBSb9EcFpnLcwhY1zhYM5ruw8EmXb5vzkICg0Mr21L3
A5qos5HVinEVzOgvoVT+CTOOtiHcKyo5eJM42HcGF9myPTbanFC8Qw1/IG5G56DSS40dysRVoMTz
WkDbagWoh5Cri3gX0yjNwja3O8RbAt6qmgQAYxuKQjSEkBkT2Nzffadne/7R3SAz64JFradtTi2a
FrQhQmQQnU+9HKAbO4pMIkyq6UA0R+lkq2pOjTrQSHitGBwIe/EPYAshF6Vbqvj4NBbq4TXbcsfk
E8ICkkCIc8TbSZH9rAUYwoggLRbic63SdwiY1pa+zEV9EyvED9tAQiFxPlcJMGMcc2hCDooFEvTN
blr4NC9GWb5lurtr4yNrp7FvdleAcNlv3xoBXDVBx08posTBB6iOESsPvs4x5DRck1tm+TN6RpBd
qa32Qa3QwXfzywg0yZ6GQzSvef9FhYgOMIRnrvFhipkUeF4nAVK5XI3r+YCwwL3v38/ulVsgKcTN
fmBAeU3e0QsKIudPbj1wIryNkHyTzME3ViPaR5HpepShG4qqVt2GtUm1o1uc2U9Vc4gCMzQw4T1b
22xLlkihUbifYTz/oFnjvjGlUhZzMl2GyJ0a4nsveN822zeq4TcGDDW3/hUqjzAplx04O8lWpCMG
Blp0+HRsWn4ZINyHK38EsbofLZ2rHXkrOsAin9LSrDGVuhCEkPGuN3VcEfZ8VnaOvReDkayzW6Gl
K+Dhv5JT4ipGBLt9ncOcIjCR4WXYVkIxOSqRwhJHTGdAF5tETYnN4twibjHCdR+ZxEfkuEnxXUu2
fruTnRC5q0+5mR6TkVArHaawx9yW3eEbC++5eQhHRhQ+xqrB4r2iHG8ya67rtL5q+hhbvpLA+UP9
NaUJRFHQ7MUZ0O186iJEIL+htWR9HozsygADx7xJSB7QZtnoAjLd0okRN/p1QkWbKWw4obmD3Vo5
ZZIkZCM84Vkt9JIO4Pjjq0KrNj6drrLcay+3dDPttcxSAh65gdDMMFST7UMPXID85r7JY2GIR/eV
NY7GEpR3QKKFi6Y0PxirOsXoITU1H/EiKQVUxt5RI/g0nljmzbNBoeiYCv/TiJkgmdVNEhyK2FT1
xNUrgn3fjBTTN3npTnutXVT818/ZJPXtd0BG4QAErzWtC9RA/e/8dWyzEwpZ42gphPOLBmnN1IoR
+BvjzfaWy5y8KN8VWjD9C7nGu8G9GRnbbqOs/uqC9b0xyRfOzjrvGhfctvVn1OYlN45ShcbXo1yq
6D/0CcMXi86HlVym+HypqBvhhTJEBPc7aMybW+hWaIRnEPi1ShJ30Tb98Vn9t9Yp1367PrhTZqid
uXQjmslTNKnr+dI9J0IkQGb68FEi6R/9gBr+n84ymTzLODLlkRmn5NyyNCK+sdfDVFuZnIPJsfaU
R91mEjJXA/PqmImUpB8uHwaqBvYLYsePFFdLfTUJP0Kj5V9K0yA3rku5GjbyfSJ8upDYIvVTyLJp
VDObJhp0Df2UbmrVk+G20dPmfxHGDFIbpMgZFiPB1J9tbyYPjREaCJnQ0Sdk4ljMPCXrveDKnqpM
ovBDgEhcAg1zhybTpB/rASoElKkPr40XZhaKRMpNtRWBoIfYVKinnrgkvhW4E7Tm4y3x8e5xlr3/
NRYBnupdjUIRium97hi0Rkp6NP8KWBb+SBAws/6th3gQcf6P2T9H2N7paeSUoGZjhvvm3jiM1VHR
rpxdvRW90Fs3Z5uFE417/YeXFf3aAknw5hppm7Tq+LSwIm4FQPWx0vb/ujHROalSIWaqfJ4JVqoX
m4DgMk5OlwHQbURIDhDvV1KfWVagPO2juJDpla2jmvGZ3BhTZmtc0b5RqZrCAMWT/nZ2mxr4GbtK
/lk2s2B6iz8RH/Z6Y6hpwwtHQItI5JUG+aGmt6GR7B1KbUvcEBluovgeaCetkH6cNMoCqtycHiw7
fpjKlNGLHRxv69e+2x9acrEsalhk7egUWLIAalPmyEg9eRpKiwXOo7JvJwZyV6xEcY9KLJsO2tMD
Xh49DwIPar42y5L5Mfjz8CQUSJS5IaDHWMv4q/sNDHGR3n+H0y1QhSCq6qd5MtXdlOFTV7P/DaN7
Dnh+/uqOO90DRq/ohgWA3b3NC8Grupg0WRh22DcNN+eITCYm8/oJsKzPs/o1Stin1rH+s1NugYaX
6d5ivZALRrIHHBMZyFORuEB/g+xfrugRPBS46pr4aQsU2rfSLV/zzpdFQtt8jAhBMjez5f+7dZFE
R+G3x6ppFRpI4JOU+ugBYEIlm2RkcCLvG0r/Fs0rPCnu1CBfbovtAXRNhVSbuRNL+kLAASTWAHi9
kKLbTuVpO/PPBpaV++bGpgY8VDel3PbfF0hJLPL4OqJlE+8cYjSZBUFl3ZFNPtmsZBCSzAhd1wvW
PkAfcRh1oZ31UVUH1juahdUIkt7P5fgfru9wriGv+2aa9lYDT5BHg59ahzNiC2WrChXUmAt83hRb
0fWcn6GAJBLnn4I8hbl/wjI8OqsRx4xt832K5El+fdk3CL7sE7UweaEZm+g/8mZVhAdr6A2yaZjV
2ru9F2LDPEnZXAFrCiON6m10aT4icW7yWB2CbkSUcAbSzZzbjC5U/VZGWLcpKYDzakLeZ+cwmMgz
cMjLYk0leu6/um08Eet2snBp8FKF9KfQEqKC76QAQRJxNC4q9oSLwqYNt56o+80j6Bljp96gigHQ
fwaWVVCCxjmZizzcXf0F+qfCquYn78crY3pCcIahwulsCytBHSWLJLi8gxeVH54RVTsWEVEAL05U
kEYHwlsiW+LuH6C9LndaOwwDDnmGDktH2JYHM840CNefGNepPs9ZQ54hNnhgLAGqT2blTGx3rgOv
FD1gA47SeHXHm1fgIrygFxyM7EIXsSWDOxVMllAUGgU3bbePYOvTDyCSh+hSqTDWElSZ0Gnd8bNM
k+lM1hq1wWUyfC0+ONehIrxmt/SYQFBLtjtCbjT2kFGwwEcDTjYhQ+Z0yDyOe8HfucCVxN0VsmTv
2cG0gDhUDExqV5Rd/SHWslajRVLnY3cTxXnJkWeHqhBpsnJyUN+AX9+xnd1Bhz1vkF3PkeoNgJLz
vzelJA9Jlbei/cJXCwstDhzfSVGL3vBJB8/ke7OangCA3XnKRlPRfmcyUdpTei39GC1Ha2ROhNgM
YewaBLuXXR5MejAKNf961/umGJfU7g2UADYL5EqGp2C/W6PGNGh/P/Eaq3Eot9vNVpkxI5KHvRIn
6n5bvlhZNqbw4YFDP+PZnuBwqXM4y3utFgoeL3GjVZ3Xq1R+vO5/8y63qA0SCoJpaCxJoYy0tsiJ
7staPkIN31UZScs6ILlGq4tSkuAsrvvHp79EnOOFrrgSAtJ5h5ZI6C2NTIg9HBcZ0Luu9u9v1tcB
AjlJq2vvZb1DTx+TgwoAYUZ4d2Xhy1ytC2QXBL+RcbQN4otpI5gxcgFVrQxXtyArpt4zzpq7YIYD
ZIe+QRULJoZYz919DVu4ID/MWK/ZW21RjZGUhoqHL0hCX4zNjOhWOql6gEX07GZJqMMlN454RmW1
aHmTO3U+go82/S9RhZJSvUonjISyBWjAdJ78H79DoQA/W5DhogKmJAUwpVtfcudqGq+FxxH7PF5j
eHEl+c5QSBKbRaeuveVjQ3Q9HYVawlElz9TlnkLvV1H1fItoEUcSpnQzYsxQB9Z7hwDbwTrDt/AW
vPn7eBn/a1NOEQsHp7hBffRoDJhLxTiPPDHiW0HCzoM16h+2yhoKPsfz3mvRh8MHg5VVM1oVgX2E
los4r9gcQwPIgeQOBmw+tY6XQpBvhi1NmkyeHLumTMC+pqKuH4nFxh8J8m+xZmQOqxPIDZLRnUOy
Tl8nFJiXhutaf67HiUyo0Jf4eUNlcHkH+P9FfwV5ZjheRXo6orEfIudn1EIJhxjLm4NwV2Jd/4Pv
qKESQTd2O3IOLLimbTktfamKNxBbv6w5TPxazgoBOaCY4aasrGQP43Z5l4iNG9o6HT5Ks5FSu9y9
YUfClMjJ2YV3H1mmHDIV+S1OB8ZFbDTuC/20M1JXNr5tmzlwbp803wGeGzIPpvQ9wokj6jmIioZa
KxP+bhAkNC9cawa7VweBtc5LoBZKixK9/9uiI2n87Mtp57OxIU/nkLsVxUMox+YB4fXIjcfa21Ut
j2qS7YeJhjBxtlZX7m+XduoeokcGTV6SI479JH4sOEZ93lLeDBPIiaEpabJ648A3tGMQvRYo3Xx6
vPrbmjVQFntlbiKt4Ooi3pCUnaJVCcNf09w01aBlFYvdgbcqCY0/o0U5Bmv+q+XGUZ416baFJqUO
3kYu94JEaqazgBlawDBZYLkbKcY0yqbBElwPCdcTc5l2F1K8FT4amSK5ztRz4yFFtu1ihsVWSh6+
dh2zM+hnYUXps7Ffnr+gL2NkPPm+wIuX6Tb0EPnmH/5lKvYwNIofAYlZR1yl7hVWW+cbnM8PoXjU
zcWwcyUg7jHI26HROjKQA2lJ3zF2meqZK5UGDz5fFXBaFMcuEbasd2+r1NW8iKAnlGMOgq0zjJ3s
940RDJ6SY/2fB+KwzaMZIVnWso31RA3WVQYPZAiuv3ayWHjQVi42MkPtvwmZLuwYRNVWhJE76IBy
evQBNKfThypFnTRVWPf29lQbQdVkmWLrfpM8Pg8tkQ6LJZODCUcx+rWkMo5r3wUPaS3XNSneZC15
zjNid1/TWwpONstU8PoUcApvaeGDnenf5MPSYAOTDGvWD7bb4YJ8uKoRYByYqY7IgjA5hTSczmQL
PoB8ngf5Q7k4t4d+FP1BZJ9ZF3ZQ1Ektm2oFM0nD9cMlZCisy0NgVBJUEXogW+4nSwibADYH1HlO
0aGk47YWkecdJBbr/oQC3Byw/+V2H2ZNiiYtIvRAqO76yF6JwvV104tf8+1PAsgUEbVBP7mfbboC
bNn7YloH2agud+JA9usy33wWtZKB8qqGoSIfV9fwPiSLjv7wbyCSl+YgU3n76saKbcGgbp5BrB7w
cfLDV239irLadVd58OAyjBLtbRilPiZYeou1Cycnye+N8jjXWfyuQRUojtQDkNQr05Rur6GSyHJX
ln3i12J+dZen9lb7Q8e41aRymFkHgrF/E5LM8FCdVCgA5SKV8836lG0LnGiPowzJRaK70cpLWkvM
p6fk6BTBvZgdVdhND4wcoKPL1VfKiHuSaSFJ07FCwmsf5XGPBGf0XkSVkKKv1SHflpVoTbsCsfa7
T0w+EefwEVAOSKx95kB2gpANsafFE09Fe/akmr3oQvdfuR5RidFYXttXhRlsv2TKhkW3FX88vFZc
3qLwfazwx4xZT9Nlwce5V0mB4/UW7eykjdHilLUjkT3+HBZDW+tGUBYGg/YqRYYEShJS30JVy3w0
DWNejEPo7CvEzLjuqUVZfPZ+5JFA67jonA72M8UiJ6L//ccD7n8PAqW/RblVVCmm2zV6IYhvjJCD
TI7eX/2mqCl9YOwh2qGsL+Va7gW5CSa58uu9U5NlLmmbZ6zwW8SdklNRbRbXnUCgWCd3WD78g2+n
cUKsQseXWZZEu3xtksmSPAuNZke0dZN1EXLZjcH3QUx42nrEVKPZu+hI/SEzh16YVt1slRJfggVw
MuJhjsVfbHVFdA2gQhhRvMaNFXBw+B1Ut6TQebnf1CDe0mqo8pcQdNRjNn9PRU15P0CzzDTqEtnE
VxUMiUEnf9HBkfOJU1S22bq4XjZmZ4UfvadqnhYBQ5XluXRsdAb7BV4v87grRNbhnEoLLK4m05Bk
HWHfllVbUUZhA52ErkMVQNaEWmvqegFmkFu9HfuXeSd/QzcUE1WYKZatL7TsXVqLiPEUVlCGPSVu
yJaIc/Hy74EvVs92BIHPZkiyhTWlBv54yhKIDeSwBhKTod7ejLDezOeJ29IhYyJriOnjou6R6qE/
j6ouFgHImfeubx9KlgZsh/ZOka3Ra4wiq65+uIc16zxnhcql3RtBDtlfckxuicWlUwi6Vmn6sG9D
ZLKBclv1zIoyWR9Ve++84ecMShH0ZFqM+PfmcxnwZ9VBSzGQMUao4QOb3kPx4uxlo98fLfkmbCG1
Aztkf1qN99XtS0zAWt8hYJbqnBFEMTTxjzeOVy7ujSuiT4174j3/b4I/JPmO49GVJtt7OCjo7qRn
n3aV+EstVO/nRRlnPhiVKWXeWEv8Nph6YvnFcCf7qvc415QwkfkEofMRFuja3qJxpnKBbd3Zq/1Y
OEm1xwgfk7ZlMMvghtfyRaNq47y6vFuxOx2TuEsxpkHEviTrpLE2dz3KCdlv15qxItaS/4/JnqKi
CsMa1MiHPT0qvcU4SSh5zVMTw0B1Vx34sU7U00n1Z2LNSTVsDQ0Qv/w9fCgzju69fhfpBzkrX6dl
h8GbIEyW73ruBm4Kta+UwkXdvwklpKJQ0+j5R9uh3nEErDFCE8Fv8Xmh6Z81Cyes6aI69614Imin
/vs3rTwqZizlny5kytaco9b5KEojxpf/4iJYZck+rhFZhylhwCbogVXLDJXGm6oP6zDOSIdbFGHA
d8P52ZhSXqQo7vb+z0ZiBYnTdI7bE24Y6qOp1iV6Ro/LTbAoGEZ+4zoT/eeJyDTj0Fo+sQjFGBdK
rFiTTSto4p0JVnT92iGhWUObun9s5X28n5O/A4hLz1ZOHAclPWHuHFz9jckr+O+j3NltSIQWLXgN
pxR6bI13h0UVuLNaK8iIClk10KZoN1xX9rIoesjHVtf47xQlhvafLiqmXOgfzpsSBWHlt3R6wcc3
fYyC2hT1rFqwBqfSdoqmewNBsSXd5H0Xkq2+Yjg9F/9vOOF6/DdkJJTdOOoDck/pLCvZ39xQfF/u
tQ9uLMPeD7H2DseVbyRssSoqnhROq8Uj5mVs62SJgnYelgxFV9wscPIBisy/Y/E053bIoJtSy/+y
yqZgAhdluFiIyu5NJGAxN/VewmIcMJsQrVJQwfhwOKKxw8SD2aAcWOkpbtnCbYUv9kviz063HyTM
gkfBmAHlvPiDvXnF1wXsSqkMIkIbQgWR8kHPxgxqScyrwvt6LWUObEPxgrBfj8/hQWtmSkByrOid
1hJqGrrRzWm9p7SvH/pQGCMZhfq28Ttw3Rvpr88gsx2ankTBbt0bx6phfZQO/yr7fYmJ4nO5NJNK
bVSl43vT53xdRCKEAGuDA63At7WVD/SejE/AcuA2M/E9IV+6ACkLU32jBT9eO7nwUVtgkIThDxE/
ccPPz7vTwb4PNggBjZQHj5KOf8dGOhGfwE+tFG8RSDcIYisv4IvdsF49RkAFF6PK/AjBOg+zqeZN
hXHOEnq3X5YlGTSPpFevHJzOPJK9vtGKwtqzlq1bCBebVFx0h5oIzLL1CZxneVx1q/6MWnSNw2By
JAWU0W4r2Xmx0CgfWy8My9Axvgjkg+lXQxG+u1o9BzqQzEu30qP+wLIkcD2E2lFIVwACFqN4nzLV
UdbHFE0+Dv6Cw5LtAihpW1e78++XgyNP4CoCVy909bdrR6k7VdZP6e/WOVd6y2tn8+59be4wd2WF
uKzxRLUBeVtXTt0uXa/WqoAvGzq06YDMsmX3+u0Tis8GzeziURm9CiB+7DIn1G8vrOtea6SwDr6n
UOpxOLVOsAzyyxfwexheBZEgtG88fcDvpzVPWCPNPMrE7CJdR5lMoP0T/SUXJ6rBNUv4IQbcCS8b
8YoNpcV88DD6HlXoewGo6eBk4G0lsSCgw3h0DIelHey3COvlPf4TPO1MINC95Y6k+Igz7yn6OhmA
mDcG2NyEupXRIeBXElCvx1Ey88WTlrknJkcJ5K1nJ4czQ/O2iNChkjwEHpmoI41sX+obhF0Utu/j
VYn3ph00KfcHedBlnshGLxkWWrTcw5n6+n3t4tZATrwgYDQ/vJ7NwdCTYOBTbd3w7i2aKmZPeCHB
3yy3fVSXHydQN4rXnXb70yr/0UXz4uaJ5YGV1KPjkzgdAOt046DTOLUyQXdaJ3MKhu1tmtnd/J99
0ikYZLrbZsCeqDGoRMgYODHURLo4gA8YDm/wv/xjKhsEo2Qd4zV9t0QBCsR20yDdAoMtLlLwYvVN
4zNRMOjXi0O4ok8sECaSYBwwsn8T9aRiMQ9docW9CwDQ8CUG2KIgGzdckUMZ8pNwalZBAINLvYP1
c7VG1+2trQw5y+rpGMQ6+5Da967ibu9KClF5Gkr/VJ8Dz0hgbJur9i+QYHHX+0nd2XkMcWHDVdGw
TJA8v5YKr4dTeTaPgnSreWJ2IjeXlY5FsV4HGukDqhkv1V9N+HYWc7tkl2fCfooUEZBaFhs3/CXc
IwyFJLnxHcWHSFUq4hounpBetal8ScKn1Su9Txl1W4KXTAeH+Yjg/PfU+PmfwKRBZtFB+Se4i8Pf
nPR0YLU0Pu9ns6NcNymYOMJP9TMcZcibyoOELZbtarYlX9lJaFsMasZyfjpDg8/XT/5YUg0wKr0/
XQqzjxr51jdOPJxvoIY9ZI7dKR3dk+RhynRJfnvPxgX00kyaHzR9upaDvyEh0EkVaIVS4a+5ik3o
sdqmQLofXmgapctUNUbYBGJPgviaOtWAjWhLHDehrJ4iw0j9FfECNUFbJZiHB9YuvHfn12AvCaGd
kK7Uq03jK4X0B4/she88OtTYEaYIjxeZrJlyyG+KJePmz5EevG6ITxejRi830rYckKWULmsKhay0
zQzbL3hC/zOYkbertcDiaoDhs6/VKi1jJ/RTRT4K4dz1Utl7ppOC9IFmL9+VFFU2PdjPpuNk1U3K
VUAxjf+cm06YUzLjPGGmAVRS84c16H66Bk3ZPxsQcprZzBTxyI6imCTg5JhPYVWgsx2KpNoehdEQ
sZPLu4a/q+ac2XCLmeo7ZH920PB0LCujlDVLjF2IIK/XH6oRg6KoKj3km6bHe364/pijmpPmvkp6
3D/jAcJOrenMpc7ewiDJqZ3F6zxzfhyv01ihLI5r6G5JX85BKTEtENwZ7UiMx2oSmiSBcl4O77qc
L7/Ubsl1vWSJVF3jqztXcuFLdo85mvgfjiI6B2cl8BmxSSRKzT+I2MH7Qa9SFp7pjutvmLIepH+E
Gsc91QL5+OdGFw39LKoFd8ks50faNiNTK+vBwHTPxBZRz/F4LRF1bsJVOpC/V3Rz6gebmFFA6bFI
w3JmsvDYzvhl7KLwK3irkmgfe2eaie2cB/MYrDMzm/0meZZl1ESGscw+3VGF2id13DszVOM5kcM4
JQY8OCZbfSzq9rXGXzLVZS5lxpKmT5rVwMc+LTTi5lj36rw8m4moc+KV/xFQcjJ0Locptd1vfE//
fB/KWJolrHRy8S1e1hBbQzI+abZYgIdGewoB5htfRVub+ud7F096x9iQDqDCFSLV7LmZi66D1Iz+
cqelSpuBqadjl+Qkspu+rsMRvZWvKgQfeABlPga2G9la3KIpO33WY5nueqUQEIhtNYLXm4fCSFyV
X/pL06Dt10fGeX4W3hF1y//EdLLyA2nOzsaKyKUYzrsurGpWsMtm4EIMQekj/IPp8lA9ejkiQxpG
ePSQ117pWbdmM1cs0o/DpaKxI0twtxZ3O259NFvt5NVA7vNQ0fQt/SZSno6HhYERzvCwVkeeGXb6
jhXOGZNBPZsOtSCUDw2YA+blxuijk8k6oDQiOmWPvZZLJHezXt8Hjrq8ZfecSHJTlXSIfTwHkTAq
v9cvgksBu90SjD+1MLmU2Hbt3VVB4C9/twxkWjjQYYWAT5J2PQ6k6prz6btG07irvUpXafb3UScz
Qjvs/aKmrk8im3C68MGapuW9DRoN+P5oBIE8VMVTkrcB8Hp2+SAaXdqiBYnvEHgAMtWLmHtAxZjC
TqR6lXd0FlFe/fFuDL1hMWgvKEXvTzzxARt6ethubxPSRdMpKgzFbqdenA1ItwASeEHUE1FVfhTX
1Cey6CDlNz2AgnDC9wAzdcaqSg6Tp9RMQppZ/kqfiATML4EE5OiVqs/p+PjPMSJdGGghr6Zof/Dr
2Osep7v1NtZqtIqT/Dt083o/7rVOUu6oWRgdMVdb6OMHXbqGWTEtXJ6YovIenaVcmw9oiylH1cwO
Zdd+JEUjH5I1Lsw7u0w3MvZlAD4xKMOU7d2l6Sa5VeJBqBVNuZE0tWrOLTlExal/6nBs4j61nI8s
cbAcW0ej0uLTmnuSA6FQvuJnF+sRaVFYh+ZzNAt8tDKE3DeGqJAU5Hyf6BkDXSrWR+cskBM7i3bb
vFByH3dlfavii6WO1GLakkUQ3vENUdWEbpdWvHN8ZQ60y61IdW74pSBbVat0RH4CzJ3o5egTRVn7
XRHskvznEvsArz4OAc2V3SfaCXrRts6D4576/TeNaL4oVwAvygZ0kguVBHL1E1ehB3ZYcNz1bfDQ
SHOmNRsUasZl2VIoTm4mWgX0N2qJG8EK3uJIvDQzNiYa+0riXS9eH1iCoCFVEXutB3M32axRA3pr
XLiP5cK8/w2tm4xEIx0zu9YvV+HgExxIin2jYX+3w6MqOvXNf0kOrn116HjzeC3OgcmtdPT086LB
TMHo/RKMXGex0oQD+foGiLeIVpitjVY8e97UBfcas3hDOFMjbzkFb7LKq6qu8lISmy6/8SPxtsCy
EEKn5nOK9egQADN2SLfYRobwLzpRzc1L4ZSsBLhxTS0qzhfcumDd+i0pxe8efwQ5/jKvg0+8k171
+5eRNLPzViMQay5cF7eOxbH+hkyMd1N1Yshd7jqo+mBuMysq5G4sIQFMqTI/DujkV4WdQjK1jekc
ptD3wd3YwAYeQTT+4ONmAKccX6KkwMTV8YKh7D2d3ddTNXCIHT8uEu4aOO4t6Qys41pOLkeAKpL3
IpSsPVb6l3UHQUhzni8STP2Lt5iaiZuNUhLvP1zhB8ymJPNKlMa6/djRP8AvG4KMLygMg1IKKcz5
KVIfWS0jlZRVliqmI/5ZMc2qmevZfXsMWk192mvKcWYweurUMVk/KhsdJRz+1CyKtegYDVABNRxZ
/p4raYydf0rHCdIByj7EyKIwl5JwRcDIj48l8C/6ihcjfA+DRhhQkPKDIF2AMGV/e9c5jNdzA5kY
HmJBIZLGRp0U05cWWvEqwb76/yUt4S2sFRoDTZ78LTb6oJQn3VlEYAjzjqBBbvkXK+bxKOG87652
8seVly5Cck1vB0o/3hxJTBjtP9pVB04be/9KnsPfngbAbJ0K0fNNeqOhNWxIXQ9H5TP9WPxs/dMP
UYB/cIC56ktG2V23FKO9QlbIQTJXl5fXrGFu+6kyyYd8CmbxntfYnFRPO+e56YgpO9TZlAgNtETQ
ghCRrRQbdCJoxWzuqIwJ1+Ehig8gtUL8Y2iBqEmiQJiM2DKjG2HsMp+jhHgFezKq7V+SknD2KYU9
tXVIeaLFtHztcUEcGZ3UAMbCOB4yvS7ZP1+9KUhw+Sk+vWzptqGQ9a5gcMzoL2MIf06Vo1fRqdmW
8mDxfNKcLLAFhSO+UoHvn8V3+abvKHGjJ2Zfu3CV2554IBjoJV0VX7suFUWnr+Izp5YLc64gM4kc
0gXm7NfZXVQQNEGe8U5nVMK+sqIlQzz5dLv+P/km7bEMVHmis/eFd8RMXWTA3arUEJbmmLnVhJPb
uYF/LJNMafr9bTaD8T/YivvUK/9GnrZs4rx9KvMfJPycN7lwYPvtEl65PpJ/lF13oOMRvol4IpiV
fb6NUcxkWF3ECSV0afNZSUJX3tS/aWRfRCzxUPKevdFnYnqociim6kJ/xbvM3aS+x0WVk1M3PtH6
d2KR+MlWRRERFVPhXbdf4X4cK9QqyUNwzB8/oxV355boagaeQX3GM2g2IGBuxTWWdrrnqdTRZt4r
JUWtXcO53Yar4loO521F9/WMmLFxDUmpy7rrNscUBAjV4S08QEp0gxE1iB1fFhXu6OprMtJE+OEi
iDKDovAulu6EGYSHVGU6QD/oPDYHafy0Ogi6gPR7Y08iZaHpn8o3l83gDAto8OrAZKy88YZKTJYV
e/K6qjxT8GtuR/sdzC1cAauK7Qo6UEEietpEeotIvq9sy9MfkHM/kIlueWiyVjrdYN1bReOCsfPw
fh4obOsX0AqPSGDNoQK2pmPydUKTYKxCzB8G4VXlIWAWYJb8kW3u38a8pfubXBmxkWeR4iqr3TPs
yaJs17vJnmr0JfIAzejA7jNLwifTBFLAsbtwePy+8BuHrJ81G2YKjqLW387ejt31UZscewAj0qMn
PRaXIEWoZcv3Vx+O+n7GR+M86D+uqyELNZg4Wo3SJ3beFDXVoI7+tdkigY+uhvhCkSwKpgThI+ls
FGXrKQhs+8SmNsTIClSmnp1+2T1eBRWfj8tbn7wSQC6776gINj6pH+jSJVYj8WO++uisr86SQer1
E+3xgl9BTffHgF23nss25TojJlKicpGy+02pNp3BZrpW4W/wqnJkvyqibOdf7Mhf9/8hrckMGjbt
HNc1DYn5veR/B+r3ZpQK7QLkae/yCNKraEd4mKZ9pGPmQCItAxgfxJtVdif4mVHl7zPMFmhxfhHh
WKs9Y+qPL0+45r0f0JMpOVZnDTiDucUrRC/NEAf+PmgovPLDSSizBUrn4TgcIqBx5+Y2RmYONqeF
hfUkSn6MlUzs6i47aQzMo7ELffaIwUSJjqSPu3X2awxdi/1PGHWnvojIuupgfRm0so/qamw1Joxf
1ZzGSgRLm/j+d/EkDckeLl+Fduc+Ih+wKmZDpklmtzvr3A17yhqkhFgEX+XP8FaRIzCamNKrnDYO
uZcasc4h13y92QaOxFPXu1HICluDJSrawpPFtwNElinCPdkDsRsLPGPS1xc7vyyY+BlVSNuI/oKy
3lWJIOJmwt3A+IEEJ0qbuH4D+DMevalgzUZFxDkZljfbeOqgnwlRdfeHKtBIAAI3YihLtDkPlTiJ
Z14fXeiDHKfwJtTJIXI0GhFbVQgsBwoRxliG4pL8mWnS5/F6Tx45xQXPNVelASyQz7AtPYkcoTLp
R+7eh5tA1q2nEEtsq7B85PX3JASdz0DRtXwidc1E1pelRrpcTkllAMEcfxL9+GAmKlC10vqkLvB1
UDAZ+oPpRrEViuodRB40YBZCV0CXVtTT6SBGvVfJZ6YQ2UJJ7tPA5+H1BgxZ5bvVNsTJTYGQFJIP
5PP3qOcZZChc4lRzjIOMEXdtvef3wFSKzYxC2Lx+F2IGxIi5BUWU6yLBlwzByN1ECdNOQYfpwRgz
n4lTHMwntxXUIaEzMZVYip2kMK/Ld7Z5Ui+IIpIO20LJ96M7s9jU/hX23R38HKyCa9faHKLGnjD0
jF7thrFvPYWNP4rd+tSCCvFwlumLkWOBuot8ZvFa2HEQO7VNV6TMt9wKvZfvRWI8s2I4gbio/Wk1
97wqorGu/yU1zT4DGdPA9Thf62fyjtBK0GR7MVmg5j7OOzEb8Rvzkfin0J/ZBZjXF6xt0Sz2yEIF
a8qqH9ELktncJgdt1dMmk6HVXrqL53dd4nz8RC0X2cyip5QWv6q42cTFhLg6uLy8xHtHZzktztTp
WY85poWGiJEuaPoyWrhyU6K99KaV35wTXUxpeCTnXAyFEpW9/B1t2pIuUoTic9JIj56QHQkxs0z8
XMGFEmxl3eCseIXDGFdLKh8U4knxuX1dOwGNB2Zv+ZQDooufOHN6LjUI/lBGKx9N6jGWKckE+xnY
GWBmEf7j6fc59merOOHo3/KnwTsS90H+hTCKcCc1ZtVBacscyjn/bHanLlIkA9s3v+FEet6MZa3M
5bPVsHkVqr8YMwSx4n0KqceiQbAlSri34bIKhPwCppgQAwa8RBXsH+YpvWkBjF/bESwvFvwtPWv4
Uyx40sLW6dj8Kkw06aoWKrJQt3yucFc9ph8fj0xu0UHyk8hbbAPm0XiV0vGMHUWxKbNau2LIh+FM
DY87Zr1Z5ZrIdN03tN2zZ7HMdcjPl6UfRrdU+XXQiVNBjM+U+AQ3wFVYinGcrBzLXvjeX+jin0zW
rCNPohOdgaYtDCjUjjy0uiXZRdeRzN7BjyAx5CdpqocJp3CShT3a1CA9evWRQQYCM/Xc1vPE7vjF
5Uxq8W+UhuOSWL3+Sm2a6YW9g+nqLjTLpo1Vm6j/J3pyanRyWb6cF1eQWjVije7dXvzjCvEyjXB5
1w91DPbFJ6Uuw7qs9xB+IjvaCJu9ji5cULVRbSbrWuD2RffJuuLIXXJFcJ7hy4jrqfDlYB1b6NId
zposj3Ca23pHKOEBHyq8WwhFWn8hiQ6CWIOWnzMqVG0r/dIA63NhkVncyEk7PgC5Kr698HQYA5PF
QQ6Xh5FdUwJMHd+suSN1aVK0NPjeuszZiX+I3lk4BzOYtuqXshTzRR6H5hdhCrMQJQWufQA4eDIp
dB6ypEiVeXV96fqrn2zRdcuJ3U4+EE9vVAtORW6GH08QHcJq1+HuooQ92UM33QeMZtV+Gauk93f2
c8AdNVBMW//ZktYr1asKWo8ZvsvjnD3ccsjywToffdXf8oaVN2VK/WdO7J2+YLByOPjhKdcvFznr
KREFi0JU8I3SJw8e1tovJsEpJU+hUIQmgtceHyoMEtaU4kf/4r+HrZtfS9P55iJ3gMnQdAZMHJVc
npj4aGRRDZIBT3kNW0550KfmtTyiKkMjJKhGw9siTLWNz53TctJf1hB0QOsOuK8tlcAXuRvc3K57
sARhifzrRajt2aghQKUjQaPdxErvzQSR+UP8EgL6Fb1RfxHoxdEbZcMJeT/p62EhA5huk/NZUdTL
XuT54A4UCSV8Phy1hFAnYrfHukZcx+POo4NVlcd+VDgWWBb8LwnrK3LMAtCGel70fCczGOzgCaoX
i4E74dyPXBfm4xjacB0FOzbsVKPhnpgiBMbefSzQOUbpXOzMtEd3kqUJntRGtkz37jpBHl2dQkLs
L3258en2rXMogj+7wywlp0iyQJvVjJT6N4/8NYkl5Sl8UwzM+imXLaSdPZp7k8uMb/vehdZk4mYq
EbR/aAM32ZR5wyuGDo96wSLWpN9Vq5Xc5g9eAJeLQu2MDIh8W4cHzsx1ZsH0bunLB1Rxsfpr0EjN
Y9BmjtUq9jmJLFRvy7vhFaSeCFA9T1fjnb6PpOdaowcC1kCHVFP7llfOhovevj2KXtHBrRBQ2h+j
PxbUyObxrSUmckIwNi3+qGTkeWQfUXod90/jbmUxDvTlEK/ayMuHjtvpDhHdtWtqvmGDJFk4R2IN
BPdTtp6NKByyzBjMvDcVS+qxnJGP7enkDnAThMERwOrvWRF/Mp5zNMCv7ZMy6/+Qg+H3pYlUL5t1
p1zeJYqYzw17adFUSFDIBFybbZjNkm31WZDKXe4nz1bvIdORWx6WRH2muB/ryz0winoCNmT7yBrj
iWp8S2qxegRnrVM82zHX23FQd9Po9xOtPN6+O13sdrZZXlEALqXMoSmQu71tTD7QlfYVRxLse8D/
gVDdFbPuN5GfNNFXM5ldtcrnul0/jXoG5eWBga3Cz3aqaMPJygv1Yo9dn3SjAKrHbfoj8wyZt/NV
9+nlmi0ZW2saPdhi9EYIL2BuoRdEX3QxJDx6LS0asL5mH/5le1z2VqZs1LF1L04KITWuJISJjOlX
hInIhg3UnxLTVGhqmv3M4WW3VJIhdLTqRyCZiUDqqy3tUtsfTzi0BgCa7By7SlxWUCEyxy7bI0wk
aU/zxmf4mDVrLcGB9BB+Hf9ZX4Luf9/qwtgfHoqdXZdGboA/zvTlU5EVLFJ7cghwNiRr04D81Jq/
VQt7C5QM5KkIguQjq7Kwe8BGk4nAaHECVIBdaoOwFpp8frga3nFDG4tCEpxzoPUfR5C6hB6jWLp3
f9SX+qS38lyvQShYz9OCG0/AArYF9bUS6KYO+enB+/vSxzi4Eui/OYF+oUqA8/9HdUkZax6HWHCU
zywHVPDQ2d7VAzVmeo1tQixvwmI7SrE5hABmB7NUJIEQL0kURycumY1bnThBsXL6KcS9xa2Fqlvw
t7uq8yoSNqWrmD4Nxl3XHct1sXYdU69R9bjxGMKYClbkLAB+2sVEU7gTNYa6hMNr3qdh1p4FgYGU
OtQ1VJ9RR2sJ7i95/WwGAIL+j/ivFI+I8O2wLqWwaszUrONireqPYyPGUYTBO6h2MSJoXGefBdc+
2YgxoEhjGGI5eN48T8LxnnZ8SVTUmB98I6TvqGNuxYZlgAqQNK9yz8MQf1P8VOOpj0kQ1POcCt/G
HtZXfFHp8nJ16k5xcEhRGQO2jaupzEgKqa3FsL+/u+jRH1p0QVIArN9dudLrOr3AnsOi59bZpCWA
X1gKXLhyoZ4cSHwyoShoeA+C1xs+IUPJk32QIaRfxST9K5eEfg3p9yM7ZaK34znYb0Thtd/GHRjN
Ippp/saLbm7fqm/YAGoHqOtvxi9sCwBesezZQiHL7/v2AdMtA0sqpHnH4IRtNiSQJwrVO/TT/hDg
oh6C4C/kWgtu1LZJorQAXXcHJNN8o5a1LYeTxgx56EmJGcFQF0yBoKabhYnexyYDfKA1YoOCMiCK
wXcyhb88eWBDKM6HQcAWwELM6yd7e4tQTgQiRvHRkibOEjgrJRaKqgbbJHqg6dNmGVIrGS/WA1B2
DivX5eELNOndVgC1ssca2CUmcxeLItVJj0tZk7yy+3tQcvMGVnm+B+PB2hQaanNK+3F5mcqyZYfg
MRR6pfRu6WrYiiIYpYbSAnO0qztaTSlplac1miFH3FjAnw4LtlZdD1lSY4NbFUcsbJjYkyLoeJEm
SoLHnaUOc7Gs4zGlF5Jq2DpaxQianf2zIOrhFN03q07xCYdDIa/4+YpAnvy9fzy3wBSnS5Tc/8i5
7ypN5zy2XYAObxJgGWhqOwH7SVLlWhoyKXZoYO9mEqlMW5GfwM2FG206FZqdfoINB2pMTnlS4Rzv
PjQXx47UYvKe2r2QFgL/ay5Q1pW2NP1rTM4qGOtUoXxxKyURo7QHq1OaLr0NGfikJaDNNdvOk4Dr
cn6/ksvik46Z2ewMugtj+KxWXeVLTWoRePpJ8osRYPlLFACjZdAPm4psGO7BYDyERXv9k6m4woO9
QB12d13kAnz2g0sO2CT8f6Fg+xWyQA3e+O98Jkw+vOLhr1FLq3XuC1x6diAgcEUsbgePxr5Iogn4
FIqNj9J82lCK6OpkW395IOcO22St/RPxaJCtg17I0V3mH7E+ddlggeEkVviYs2264d5xFxqTpdqV
NRzge25667s2Z1F20DqupY/tWey6Fj+B+wWFEGMZy32LJTfxuNaf5Vrn0/m7auNbt++XDxYwwAPT
qAlK8K3BpKR2rDz3qsGzhoQtAb0cOfojb0Snd2uMQQL7Too/TaMhghfrLi90YJZSe9TcC6xWFppJ
Liw23odPK8VMO4tEXCmQyxEr+6+JoSYXzN/WIJNkHARCzZj3yNQI+pGP+eAER7CtwsUi/d06UbDk
eHJWzst5V45t3TMvoanNYu3qggryhZRgOoKurSTrvbTzffQDkAg0/iCAOIaAaMRdB3fITIJiRYhU
s2znK4RTizyR/+iLpUjP00vFJrusHbhBuaTwCGsY+7xnbckceW8jVEB46uJeU5OBOTF6KzryI6nb
0Uq1Lsxp4A/ItSjiMWHaSzPeL5DwtuxgBvFAYgMFikLte+h2iqVnF263RU9QXYQUQszvfXVqopZ/
MdAbdtGAsIDE93nlsCkdF28kZuvRBDy/gDTrkd74QjKvwo+cIX+VoiOWmxuu9SwLacuOCfccZ8B+
TcFmef5n0JhakRtXObG3TtxTzYKJMc/Sm484Kwny+6lx34B13T6A+XVof3lDRT4zORanV1nf3ck7
8WHnO+d4j5E5XnWKewY3PVxcRx75hy/yUM1XTLWndBheDa8Ped8EGRpJKZuPxgi17GghcKFHkO/6
UO8cdY8YJaAFJFeXF1Shmc2qp7z+TZUDgwsD5JgzT6IJqGpOf5yVM2in20R/klFeN8Gl1pjKBVHL
jHWJHvBLS+Rae6ZRto+gR/RdsL350OzvfHuhyjjMWx9vENNfeC55nWVPDo9/kLXr54wFHuLj/CiF
UNVhhRA58Xd3cA8dgtW+Tyzb9egC4WjDtQYQYjztvISQPiLQz3jtooI4fwkts9m0o+8ALUMNdnDV
HBzK+sblboiqOn3Nft+ACdkraB1IFqtRk5bVHRc3pQyPVOJSyG7fdUyuRNld+ux5UB8IJL7swhdv
0RF6xcxCYGcd2wu63lNvrEHpfr1fuBW0NbnOAmM+pOdG6tn7f1TCDkCK//pZ1ClTiTHOtd3a+W90
EBO6B/okPa0LmPxErOJv3WzmOWuv/n6r6z2yg98TKr/lHjMqtMgitwgf+4XobBqrQ7GtE1vBG3OZ
BFrH2ZXFiLy3YolwN9emy8aAynenp2UKy8kyDZTlX80RlTVbnARIZYpxFd27qIUjRsh1lNJWer96
/P+q3LBrAIWVHkZRuT2NDc2Xq+N+9kdzQ8CmXrHPfZHzj6Uo3DfqseHhhu86AUw4GaG7fQhRsLiX
9L3N1Y3sAmC/lSZ+GJ9oBsZS7XWO8BDD1wjWpydKD8he0LTI0Q5K66s2mBMkCK+HY7WNVeph6WHa
3QPIeb0wdLo/8Jmuo63s3KZHKSoYkhJfe6yArPKmqOjz7oIOyneuZXJVVBvOpvyooe3SVzcTzB78
lTKC2VQZJSn/U5m0AB74lg+8opfkpu8SldlBabpfoFdx5GqwyAvj5WFQwWCMNw/PFmiqU6btgakp
HOYevHGgyStJq+WkfEHd3MJD/GVgamrrwIqP4ya9TuOimNARefqlnLAKsGf57hW6t1L0tLpIW/Lc
d6w8xi5ZznV+cmcrIrCOAue5+6eCOXziep2LGCpsatH3wVVPwfhmNDnhDLlA2rrPncL87NYRmHfF
BT2HRCEPfmNihxCRnYHKTo526inVXSRWztZKdP9Hp4BlaKaj9kxK3iHuOdbQWiKY3ZxGCcm+eD35
3SABX7oeUzxab1eZdK5bUKSCP85TAvpWYm6pbeI3LbhWea6VSEFwwvmT5z1kx3LTZA+muiiv/wtM
U4QJaYoCN2AX1686vb5j7/H6wNrvmo5DaxEi5REYFm+hPUeMvO6+/4zz/RYjbqgYf7h5aiZ+oBvg
OkMgVcDgRBfzNuPD1SOR5jLuUp8cOCQudP9w7LoWvg00LKDnFBs2sPdoDXZ99FRxAsKSN3ihxVG5
00t8sNAaPtbAg6yDBr1biKx9drHbNH5Y+9mFjHUFFqepdc/VMeUhGtzZO7K5yu8CzASfp5g1dNCx
9MlqhnlM8otsWPak17r+DE7YFXFfIoe8CPpINoJibO7sckKxdx1h1aKkmz/e5Uhi0QczbTZ8zXw4
K3OJ4hdanhv31HeDDLMSaCQtikAzPhWB/jJRF1hXFUFJeHe9kiBJFNAIYzwDDxYdcAyDAPc4/AoA
AxvfSoAZkwjC9z3QlzInmIoX6LEJdjqWdXfAeYazFf7hREg7+NmeRJX7sTuZfhgnTkYcpr19/2lT
2Lmt2MKdn4QE99C6xyrc997T/ZLFS6kZ49wbJG4FmrgbgN8SHEM+3WyxpvEF3dtw8be8Xl8v5IUM
sqSMGFIi93dSXYAJi1msEj/yhNWCFE7K4fGP4uk1RRt+3iwWbCFt3uoxEq2Npi/zv869x4xjjYMg
VCv4uQPXv6gShd1s0hrNb1NfO/lUrkHIYwXDHiwrn6TYGgZrwEXoba6f0gHsQB+TFdq/W/atSrci
c8fAqEhFwl0KZ59Ibiwo508S2izknQ1VC8J8sXpfq96lpDT5pLAIWqi4f+2Zmi6rE4maclkdtBpS
VNRSxk8igCJ0IQqXlLeWG3GXyBnBIk6UoUw4NLZtsVl9Xd2W6kDmYLRnzWEkQpPuC79yeJgrXCAs
wA1TYIbKtSlJ26yjeJdFdLU+kuKgNtohOWVQ38x/2zzo6Aq6vXivJXwh3VZVLv7dv+PWxo7zioR6
1lZgPLsFgVz1l4/24Oib/lH56jWrDEmGpvEogmymOa7Uc72QCILlQNZQT9TnM5zcL8EwBmuy/3Uh
OvuPVouxRX0F5MxT+pTdajokVBO4W5TVlzqJXxyTU1q/hoPEPVTMKJccIOJRWqiggUZeLXecTk6B
YDzfMBVEowBk4cv9dliGSedaEjgdfam61wS/qPUpwNijdJSWylg4QAlFoOu9nEMFGw7NP2O9dWvl
WsY6PK9SiVfF6y7Si3+SaLJ1x5NTQWBxhpkVswM69m97LM98HOXYLsqmwfHEL712TZxdn+LM7ERH
FpFcOvi1gAtV61G1FbI/cYgiqNSIA9ootSlQAsaLgilpCgI+EG55gha/6H5ErXAdDr0mcQaMr7Rq
5z/aeWGbM226rdr5aFAaCufHgMB9kSMxjv89EKxa/n0GCZE7ySz4B6ZikBJ9bLvCI0bTOjh8TrcO
YT6yq1K5vBjQMbwozQQDhCX25L7nXqo9o7SShF71uHw6sIzUUsnP7Vqw+GIHbsi3ZGsaXORr/l32
mkORI2NdmVzN7Ns4AlVoIRrKaDL0HYwnenf/3YMt13ixsaV94DsnWMAFjB6L2BdYlHXKR0uYSbkB
z+vmQZyFyC6hbR0C1EnhKJc/4Sa3xQFU/+7nQVTnWnkMA9dXB+kIl28pZdACgImu/mYfC/R/oUcy
REhgYGReHtfo8TA7LXQFD1+FNfGknACKL8KNphuFBIFWkcWH3hAZ8qPEJw8XFhQQc5l2GDyeaZY9
BUiXhpgzfrAmTZCxYJ8n2SEWccA6ne3gYQKKQSIQoim4IFCpm0iIMgrAUsP3XVGacPS/FmpX3K0S
o9n5crgnShEwuQ4aSE3M0Q0Q/nGC215KkwDqU+TpfLiTY7RgCjObYsT+akbZhDjA4ktTpfcmKFM/
QwHwJKN1T2WBQkvpjo/9TWO47AcPFKgH4n5mjJZeSZDDDNzPor5y6WtkO+HSonULlK948G6s1/oa
2XF6Bv3qMaJq6QX08FmpG6iGSPg+TxsJewMaqKpTo38fVctYkjVrycWvQ+ZWn2VF0grwF0DPpGP6
3qZIHFOn0hp5sh4h0U60/VScKfjZCaFfLz7SntgW9tMtS4HbiQIkFDmuf/yG2YDpCMSCbTqGe/9M
BSw/WsijbcpjK2zKPPbx7ox26HjINDH7q3UM9jzoJLz2ymOFRJZAlL/ks6ObSNRXp5GxJGPm107Q
0w+ASQ2ThChwVaFYWFR4wcKWv/j0NF10uHsgHgi+Kk0WuW/8ch3GaydLifXn2wtA9675+elx9nxg
HSpm9sy9B5Ufk74IBCv74wCWTjrcJ53EZRiZ/VU6jXwCX1nGWtXKCTReGLubiINTkNHzMwx+AG/R
63r3ovd+teGwIuNPSjI7B95ccvzmwduVIhOSQ9D2yaacWF9cGZI9e/QLqheKMS777fADrMcNDaMe
w1Ez+Nk3yUC0UGpN+19ejg4T/dlG7eMIkyvgvAKWJA5n0l0aM8GqiK0I+BVkQzH5Erytil8vujHo
zcCn+mQqFpXT/UiMzQeB9JyczKyOeu30HYuw7yGun8VV3b/MUDN3s9VZzqyBnbw/9TYeWv4PbQ5k
b/7JTzWHrD2jYozY3CW3tVSKis2FJ79Ltj4QJlF0ls1wMMsBwluXNYW+tL+pjrr3965wNjtNKxNG
hcVb4K/9o0mUmMxks7g6p/w1IkFD58TGLVgaCKqc1ZsUQ85BDVxe53dVmxO2upOMyl0M7zUo6kvt
MxgEkqfB1GKiVA/OxB5pQrJUAythti7nH7UB7SVxR1lyVAxOTFFPS5CKiIp9V1gbtkSaJZsgZAkz
sijDiiXS/g/gdPExH9S0C91b0GNKK8dS8+nlX1RDWaEReSeWvxgHsDAQvd99GWhCanEBxO61PTjT
Qx+CLIXovN8mq4dpOAftyx3HuTncUGMyXgnOoZTVi99Vdp62Fm+xa444Ne9K6WOTPWDWP9OSsmH8
22GzAkh9UYi34HjQCw7cdszAE7ZsWY70LxHdlOb9vNyhK515ovFJksMv7Uxsya14lXs0dv1U3+qA
tR706vDYGWH/17NSIbBUb5UrMcbyErsJoHEK1Wfn1Nmcu/VZ5HP1osk2c6Ly6yMeBmlHPIZvz6c5
PLMcciLGu/hgNQRMi3KHV8xkV79gG1AQBEqOeEiYbJa1ZnfocHrPPy+PEbt127V0E6a5n7pN8cri
LXr8RSxgwfqjudUp/Zc7iUPyWm+UHuYlQ+HqYAeULzCuffD2IOWBmHmflFWg8XfxyI12c5aNpZ+1
4NinFati2W07py5OTh5rVHOG5KvLjBcd/P3G4ENkE0Owi2YRiwqtyN8FbE3DLKPPZCpjMGfpFVja
oi0BXWsXqJR7h8VAzu3yC8PjZOr9rpV8JWaEX1cPs/VbSTcdkomuUBCRPDG2Kt3wtnK+qQYQpqsw
P5qt5h70vuyEF9ZVK2X+50sa/cy0+LCY+KAdytU4cVSF5M8UW3Qgfq/KuUi/DHEZU1mJqwVIEkIM
ChPltyk0AzkPyToEzKdg3j4hRd28acOuxpdw3KkNy/ILm52z9NoehUd+XZKpe8XUcwL6rWis8XuZ
q+AF5AMMRNIEHlzzVj3DFg0bZv9N+aW/1f0peeAfST1pkdhAHhqzXMSJmWohUkmFGz0Q8SZtpnlh
Ds6k6ZwAiqMoWR0UCVrEDSx0Y//SGk9Sw1foA/8yietkI3Cj3yiQJyNsBoWT1+XXXbLYrNfiH2rl
53o8P1pFe3px+EN8JiDpvqZCQeiJvuhjm26LZQbwPYL85sHaIPRvv5lNeS0qz6md+1d0dg3ZjO3g
XMf3Dt9w+mBHRy1u7tOTYiSasevon31PzgCGm0XqP6suYaxLpN+0Ry4jHC/B9boalwuFt+hMLcHn
KWRF/Iuzuy/zy0+eoqj10MFT1RBY5Ud5fQPNQmXbMvSPXyYHa7dihPbprLFG/X8J0QTONGHXcDXj
0wG5N5uKjI009itZFrEP6f2KfO/v+e3fDDnOPpszn9y3boP6ny9YUqaMaZzHgiqAaaZtRjyIAbwz
3Tp1YdYVisP5GI57kznqP3O/E+BuMpdp0kzCVCWHqu2pUo1iqYzEa2BAnpfXeivAwm5jWIacqfyE
RF2cApmLehlGImVigPYpFbIRlYOwsm3y7PkCHJjscTRg+UsawMdF/7bamnTg1YO5IzyNSAlrlQxc
FNmCgvucl55zYMDegYOnL08aaUUy2eh4GI86sdp8mMypVZlhuWaD0g7J0MpWLjpePMKwssQxbs5H
wXTQsuYY5dumCQX5GX8c+cOxo/D1hqGWf25m2wafnP7FDDbKLZywfy+eHMCF2qiHvCY+0L91TSxS
fMRgqIsohdsoJ7ocFu0h9miAPrwzVoHcOdV+rHm17V0UMDwxxk/jJ8IOfc30ggT+uRq/onlWZWwu
B9qU4d27XGkSMtt20FZUh9YQpRZ79WSfca81UIJ8/ylIl6m//a8h2sDKo2R8tkj+m5Kbc0CyjijU
HqDO7MBWD9ha8Ww8d/ocNOnn9j3Ts8DSdPoTwiQc2zaZgFwhkiW2WUUIamgUTm8Z6KLODAWrgMzZ
cK2tRjmPehJVJ+lXPb2Enm4/iYGW3vxUsD7JG3C0syFwCWzN0dguFXhH5wE2Kwn+55xUZsrdFp/P
tYeRIleSxfQYsJAk6FwnbohrwdpkeMGXvPAMLSbIH4H9yRbSQ7U8PB0Svqycc4cEA6oJIkAVO7Nj
gJOjmEMpw6dSyCCspdWcfAibjkIyL3iAWJoYjGI4sJqycr6Tz0crlbicmMO/XveGb1qtdD5sfAMS
TC1satSy3tn+DgnWz5A3e4gmfymFaGPMEcr99FMx2xoHlhC4nhMpX5tWfJd7QPragA6NxPBRdjq3
o/AT7fRyCJV5eMLNjw0UTcN6lmfzJhPMWsJwi2rTzZPlQEIodauKoQrYr3lW8f1nJkXxgU9mNqEB
thKDFEX4P09ONe3s/K37hjNAYbKyltTuvuUVXwl8UlEUJratqoV4vn2xwV3KqLhN4JoYhOx/+kD+
ofNEc6NOra61QFsAyYTf/+c1TP6dz8GZX6Y0svojFqnm2WF+VWH8Qj//WVBD/mEIJhMMjlorpvcr
NdgxV05JgEXOWBp4cevA/gbiEDg+op4br3bqTAy+tE6KGFKVjZAp+P35OHBT1bU+TmpOcyHUlTA/
JQJnSaPBFoSv2YCGFvHMDb4W4cpfBc+oLkBEjosDDmti2XE2Sh0DPfUvp6bmNfZpkfK0BKoZtYKA
YY5FjDyjT6JPrKeUKB9h3thZtgWTbItJOSyeuUHg40utf2LBNp5itdqSEJtckcC50OV2nr9ONH/Q
JJEmjb/6MDK8U06l5yXaGA5al4XW4npwa0EHlgHVu15W7Acyv50k31RWDKISCK4ALkAKRGYyHmTG
DVsAxNZE5Yh96sc50Vmei4J0KWlk11Ygd3TT31jc6HWGlo1GeLSbD0g4Uxfw8EzogdRJMO1BGm69
nXieKPj7Fn2GSDLBkvgFAvdM1u5/09CtP6JsADHYCFBr18LTlvQKJYLvCmZ5JR+/vejIeot+6IwS
7zbNPEe++EEAIIdmCiggRgZ53/rsuT1e3yxVuXPCbb6zA1qTAg2NE54EofMKLcf6Xpzv6kxqkVGj
xuaQcFMyZQVuxmTn5AdTh5VnDX+VOn+Y49VlEBJT+D5rB3ZfdhsB+zMOzim8eKQHAGy7Bsj3bNtw
ULp8RHO4J5gJ9k70EOluliXpTBGuDVhFsJbaVU+AP6N06j8WYVFhVJLmfzf/D/07JH/42xdnTmZd
V91RFB3d+ZgyL76NEoqiEPJ6mrsscfmnFOaWPul3JK3y8LqP30ZII1KNhPlirO6402K7Jgq9ifmV
239yuPBgm+HpSKy/3HsseT7Kho0eeoM9p1KvWhzt7+eSQTBBd55vLi8JwCavRFaVJe08rFRae7Y3
BLj8tgRdhE9XJbSKYV+1LwiQLSzrD19dreDEem2Ecfi+ey0XN+EyooOm3NVG3Dwg+1GEsfCuh+1D
GvO6w+Yh9qahGiGXa8mMbUxkT09D67MzQVSbNf3EdvEGLjUHY6wu8hQKeqOIITIR0Z54knACvYCv
8ZNeyw2xymybrs185F8kKAv7pUYglA8O2IBVWCyHa5gsyB3iYyalEyRKIHnEkzknRLLKpMzt0yI4
MApL0JRyBw2WuiIhhCajs945qkfIjSUxKm6AefT/jGNa/lXPfZWDadt9R6OLSxE9phyBx06KbgbA
sVcS+Nykt2YmbemTuw/INqW4Q/BuIuTE0Z0ADsOQmHjxFAPwmV9u49z8Ect3ZqQ/I1b62FgQu0yo
17/nTz2Ca8D9YEIwmz9RWwVIAObZ0vgxLsZsA9dN84GXzY7GGESf/cqf0oIvcijJzPWDivseX3zU
lhDC5P5A5+ueOs03qAeqKszZ+Ddx3Ptgz8JxntVnCtnYRKskll0zY3LoPVFq3PF2kUmb1zOzBDFY
wlOtWv6WpgPkEmFBVGQ/xfy0Oyv5z+/58iaC1N0VrjCR4FzudYkv91GsOYFTGSM9JTcW0gy5djED
1E5bOOr7PSv79YUWjcXsds2xqQus9ZzZWRtbPAsTIvwVQ8+I6eGoR8IghcmKhgeqp/m2eT/6W7rO
3hXHJOW7B7QnW5utK5n+9jOtVlpb5xipVQuWiFO+tOHdxc10M9h9kG0ThbiZnHCQFqg/eiPHIrie
WuR1hHYmtK/eQSUTmFju+rVc94l921/C4BTAKDyZR8mndlv6HI3yDTFKfL/VdS6HbIM76nsp7Jwh
vOxWb4opXrBs8t4FIydsBFYxCKunmnEqbfWRFonmb/8zOeaimvOnchfqLnOfMD9EyGR1OVVU/zpz
OEvJHqWW3lJH9dtfD1tsZszvWdNvkHOQ0N4xlfEloxY6rPXpIemRDYPEGm49mm5YVhwe/U3k6l1x
Se8mea3Nzm6mwVfHQNgBhxiFs6g2A7XvS7wIRhkv4ko4OoiKS5KL0A5QSPdjj13o/T6tAbFjcTAI
q1xY1FCv7KPEz11jYQGQR99JSGkQLJiZr50xtBjDkOtqj4JsqzHUngTYCyYivZV9OKvVL5N4Idyq
FpU/xcm3alImHBpUO50cH7KenHrXZ+g5SCXM+3GDx/KUfGrJc67033h/mlXaLpAVAUqt5Y+pyCxQ
zJPKLxHjMP1Ka3h4Mowel94YyUh0SYtxToLSxRP/l5PH6LyEHXQewT7TmzW2XGN+JW0kJqJceTE9
SWYu+o7qjtyK8cW9PgXZVIW+9Vj6HFHBkl/sJ/C5CW2oG9Wa7RFVj+Et8RHFKSqXenBjNeJuuvqm
7cD6MZN94ViuyJMKdlWmWHjLOPBVvvZBv//9NnCcJrahJshYHuDyWtukYqEFe9X1KXuXvVg+gpXQ
Qe+G6Zwaod+evH8z/xhJ3ClaAhinMYBYfnOl3h8xbEMrFp27w7p7GjyMXBTAVGuiB7KSGgH2z37k
8vdjex81IgFO9iesMADTx/Pz3VBLqu3NoVGbdRXzMDU3pHh0R8LjwudY53lr8r2QlQKBaBw7UaIO
z9yu+LJZsP1kV0xzKrfgJeCKn+nKyNdbr1ieUiNHJXN4dTQWTLTa365zjhxWa0VAwqHohl6lsOqi
z2SNAIERNNusy681Bzx5VXEr7aq1R/g14jVilNutTZImYMlHxNEt/TMyXUtCBntwffbuaL7iZxdI
eOaunW1CC/MEuHl5Z9ZiHcTaT3UC1h0aN6zovG1Dka0Ivo+pXnDU42nxS9Wq3NKpG3AMHpu+liHR
KvXZgLzVM759hlYc+DARtYJZaC96NEiad2C6v67rxU+XuIl2xY6xhYuYLe8AEKLT/LLZUfgr/dax
VAxf9LIkq+eZGLDKxLC2fR9rn2HR6Y0Wa54nKX3qem5dWhyYU2UC1+PxI4+MIMSrlG8FbENO++r/
8LcOcbIH6pUzze2RXPfvC+X8StS8oxfvAUFgkPol3dGm4BGxJ/GEpnkNczNitEpbXr1MKigAoC9L
L3eLbi9Kgnki7iKsKbSsxuz6ZzVnYiwsSw6I1t9rtX06ukfmV871Y32hcmiN5KNBNt6Eb7D3B+fi
k7J7GWLpX2zoglPvfqUsyti9aUWlvoEJjrZTj3rJTyLj4fj7C5XLCRwGkyjKfWoeAq3tw4I9/g3+
mK/fJyOll0kk4pUi0oNPZmopnkGqGWUgOgXhpFPMaKVEWXdvSfG+cWKXgErs1Mt4sOx2f39RPsOi
N5q/Z8HRbkjIg6p2F8b0gHUttlV3nB5dWMTR/ugZN59zEWIaiZxEbLp3xZoOs6lSI/vuLgkzkjUR
I4o1mfiHq0E5ssxas5iWe+O8WirJIQ7iYgUhi/zDVscPdZ8q+a5KxEbhAmcR240daYP3FuNFBCbH
rZyINUZWNB8COKUg8sQStAg8zqG9H15kX1ZARAvPFZx2pFiR68QPGQ9N9j/NIwpiXfcSSL3Kphli
JIi9njEQSL4iJXJ7yupx0JSZcZuMcDlOnaGwGAEhmSOkLXaPrbhW3DiJdSVdwtzdmGXeHi5cQ6Kw
ylwqO423L/rmFfGphE0NZYubgof7NG6NIJN8N6Uvv/xWoHks7loyFReBLMOYgkjGpH5Rnqdbe+zt
ognJncv081WtGQjXEGmKd3OomT82u96XNyEpn0eXXmqvgobS8OYnU3RtXkaRSqJgKEPsqSwMIXIY
WVvztrdXDv24HMCFSDOiqee85T2vkHQpjs+Fvg7Qw5mJ2iCKSApQuU6mru+ZxV6MPK5IEW5FBAL4
nVWMsTA5PUD5GdWyvVmtrWkp8ZaDT7MFtypCz3vWwTbrCcB/PlEgMWdyZJF5/JC+b1V1SlNAzvLt
FTG32IaA02KV5s82joi91TDSaDqWjS04ubr0vYKbGJJAco8QjyDOv4AqvGlZCOUwTEE8EOFNOduZ
YUPYodbDAdLKnmP7zsoXReBPSq08JJujdboGHQbb/lEiW2L6oIu0W+OdVfhLa944/Aiw5AMypn2R
fy3uFgDcXnQx+202tQS7erbjHZgP4l/Zk2fajyWNT03EgC3b4e0+C9RgBx4BAnBjtiTyPXsqidN4
/Fz0+69cm2quShnuEnOTb2rgf2p4Oar94wj3wYAnWMFxfqXdh7qvKIn4LtdI2sGLhXzwl4UvG+eu
Pu1IwKsMVw+jN5ihCyIIRDAlIAqY4jn/Pt/800lo1sJVU8m7nddC6EEr/JvZDzV1GdwiUxwdBs53
wCSzlOpbWLGUNBR3xNOFecfLC5qxcDYfPTsfUggDUZK87L6k2bxPiv8d43J7Yl+U9jiwCxX1lj0P
1vmkfUiZVJsDOkvkNAilv1ztijFpTWG1WpfEjUNBDtr8/pE7lonp4hXom83jZDGloYVidIce2OeJ
Q8zgvow3HZIHyXp3nIyLSZuI+w/y4VvFSpIupxcW7c8UlrPPxURKMGooHptRinaGXsZ/HTX+TkEo
bbSwcNoaixJIwY6FYum/XxIz3VxuuaGMreyBytYIIhlE23t0qohKgBYRf5xkKggCuQcgRSSvMxia
XkeOUv+oyA91BQ6HNHy1jOkGPEX4sbgQ8j1YVjCYwiY0zwuJIUeS+ykMi4GvwZs4OmQk5cCKEMOr
CU86A22sJ6WGVbETQb9epjbGpjjHMgygbaUB0FlYVP259Dey7dbIAFWJ/sSeYkqpLWJuvm+y0lYL
KAydmbVnEahawye08OPZNgKmT9EgJ9L54x7Kyo7dJPI57BSb41SUfsMjbmDoedWJ5VDFjsI+AFup
mnm6meqFvw9jGkaCvmpMqwkZOJwMxnROc1OT/OOZB5nEFsmJ3Eknb/c6lBfumfcKpqHJmU0FlO6N
YqOzvEUw1ocCmRTlwak9pphab6uuOFB7ZCNBr08D+R5HLiDoI1m6MWu7jwl92RzwAKszxuzVfCQe
Uzl8kjAM/R7Xi3Mnz9hPXs03NVLOq54pwLY+POD9H3agGgqNgoEmPA4F13YadKiwt+I7/FFDtEt4
oDfj1ztcdynfzS/omZ0gGeRTi/BBYOWoTlZDb7kljR765f3WYAKFdq5ziP/a8wUomSrfjXgjdpwG
LH2K3n06eZe/aDi99i7/xD+cDG7Rb875QMAxNAiJhH3OWqcddobke77TmNKN2Fv7Z7x5P0s8nPf9
vXMnjyHGRmyqFoCgXtNwH3BRwDi1fL8F8VqTWoL2GdQSBRl1cx4AGriYRSZNjlc5FyZUEv9ovvHt
sO1ic7HVKsLtGaLyzEVIDU8Snrrg+nkk2rrTORysSLLwA2l55HBtZBhs7E8CoD2rVdwHT0qLWkP5
D1fIivHnUsMzqVQqVsHKYD2O7dMvdjnrsnLe8DM6XPPlCAXUzMsCe9YWdoZdLMYFpDI6+l0wtF5r
5uZ2fQa/27e5ySXoXuiXO4v2dydhrQmMURr+3P8UWsOdozTa3v8SVUVXs3hIiizawAEQCecEUF+R
yc3weHwPQdYFJaVYmhK0jy/zcCIJvM+lQ823JtPH+mlz1MolKFY3utg9Zo3nf4FlUQG6HM5CUmH9
dT4QOP8srsANCD6rr5AF35P96k+HRIA8e53SsDZG+T1LnEEfxNvuMgWWxm1G8W94uPgLbTOpKOEb
qoVC0E9gjh6jHNwfHVBH9v9aLcj/5YLXcGc0gomK5XOgfJHI/UH6ijcQ1U4jj5vPCqaHhYpRJbsS
8O/tbpLpN6iJWGfMlwSVG6stTU/6aEpOAZAYmvFHpHlv3RONyBc6/4ptsSJ2Up8nA9mFvEqxw4Ds
P0Iy2VsxAxca/Qe53/XzpfnMY0U6Y9a0TCIP5zylVIegG1T1iPyIMxwY154EXw//MQbdDtLPKZu3
uA3xjDyi0uwRyydKwrRDCR4kXQkC/S5p8CQZ8BQo4fRnl7/WMNmosb5zGtOf4ExyNcZmb/KioD9b
WDmlRxSsVOhGK4ntR59UBCgTPPJe5e7BrnALktInJg0nBT8Abdcpyh4/5/NqXogdn2zZHQtGuzgr
f431mh5fuS7u2VcICanR1oRFFjIsHtEkRXa5fhUyAkfiFwat3EyiP4El4OpJ9SH3XhC46LvmB9a4
0R/8zN4VLPQp53Md9WC6jW9aezZ+6Ivh3Qm8Ck2eR9q8enbNvmAvrvdIP4/vZt+gkL0552AY2W95
25G2SxNKcaK7fixWduWoNMcUGc4Cc5aI/msmBzzQXznzdIG5Tw81aWCU11J852M8MV8OmvNj3rAt
Wi1hhghRVy9KE+Z/sH7KOpYf8OXtI6vESI5yA+9/yfsVyciGU/IlVzrvnvV+hwiikN564mbD2Oyr
mj2vww/aWlP7+33Nxlvw9RZtP8X+UwhViYMG8k/8q5rU6Jw7z2mJyfrHnQEv5eWPQowD3vldZSWw
1oM04C6s8TDrbyZ4M/540hbyL3fSex1KA7HtwGiTjvxIy+sTG/xECopHSqCzhIM+cas+f2B+y+Fx
vScpZy0JGaZEQRQQ85jQs5vx1LSHF47SUrCnO6OWGLXrLaQTWkQFmV9KAcZ5WXG8+q/M9cdpwXWb
iaXGri+K+IE+W1lqCdKZAakn6lcCrWzKFdCzqqNQ1WFjjkAGkHvNOyKgt0GfyB1nZIBXaeYKk0vM
Jq/h1T83kKhhA8nLZrNGOFkhwZgJuFilw4WgoEjA9llwkFdAzEfZy2nHNSjLuePQwyfgJNKukuzY
8P094NattT32dF6Ia+bG2rWg9v9Y3IUekBv+ue7jr7JoI0mCRQOAhjZz+4m4lpSCwIny3FA1UKub
f8zXw+6s1Dh4kFrZ4xzJsC6IzHndpqYZM6i4bXs/yQwvcjro/B74kWYiJTBZI9J3+87VQZSjHDaZ
VfyzqiaYpQSxwBA4SslRfQExiioPrcimOK3eQcdOg2kh5XVZEFrBCNbHgr6jUATFmbxWhQPrFH0x
cqeDWPdi38VkFUcdkkZyodZAkppcQLAtqhqCqzHWr3VDkQErP7VDIo26wGUfYCi3/owx5lBrQ/iW
GlIqnccjacxSCXssnejqy68u9e4zmKAcSIXfbDc6ADEjgGDx08xVzYp567rFT6XOQ3TwMQ/OrBIm
ZJVcAgfgkX7+RS/4THWV57OcG77NpSLqLbhW8jPOxaz6Gp7nzisnD9XpXGr3qSZyMMAHQltlMB+l
vzYGvC7WDrHEDNrIJQgvR60TStcVEkMjhpM1S3PVEChEU51A4cat0W3ok7Ipb5KSYVerkw1B+Jnn
Y36+qKFLLrGjSHq4cXSSGY6Ne+gF6GTS4bYmcLh64lQkG86DzIssJcIwVEzfFWvrxp+hcOk/nGFU
auwnR5S25Ko36WJXAXS5t9QBJSPXzeHvrVhHEE3rqWB9z18EMTnoN4eDIPo1/tQBQ+GL1N/xmgbA
MrMWOJtRsbPAwzN75XcTDdC7zwVeG41yZvLibCnf5w8R07SIe9aEWeM4PwFvHQb8FKjzeE2kqaD2
iXkv56MbpUsIciNUlXv3Iku0psj9jP6mBgiXiAIILmoWGX0eSxWCYMvVoaoCMYOFpofjffZTMVDB
z/GQMM1SK/c18m0AejfF9DFYTNnPGx7GIAxmWn2xBwqSsIUJ4kLAALXRhw75HszoQMtxLazbUC6m
IFb4VF/DEwsP/eMKrTEidLIjTY9a2WkNk0v3KuGS0xiA9WP+FUJdtGbSFNHKDV5BoZPgqxR2HAlP
yk/LaBp7Qb5GJ2A/gJPyMisyV8fIfN2pY2KSQpa8Y36iWMS+9fnxnOhAeN5ufE6KUmeoxm0yXH3k
mwkDKZKEehLhwJp/CnWlVZTkC2dNJkKATGbfLDbCxZHz85ORV0PeqEI+/XZuGuMjMtiDJvcb0Ak3
oG7awqWk2rErADC0809edvk/q1CEu+hj00bM/PCUk56q+1ontGVObCbDcHAgZMqk3SF0x2IgQWgn
6yTHa0BMxC432vrdCfsBwPgLOO+gIgzgjXIhtDu+Pz1HCSrxuTVShopahF3kGlziDzvj+gYZOq0A
ckKoKjNr3WT69orMvHJ9Q5nWWEfooXK9POI478rpDNsB7m+eHgWCo68nTwzyRoVDtJbO8L71Pftd
AZltv0UtJ6B55y2vDBjCy5Z7CnH3Sr5AtnjiaEbguNzo2zBTnXrlf82uTL4BzzkHNGyCWT1HKR2I
9O8BIB9UxW5lnhzhkjLRvBLpcsKVT3v68Q2EjDehtKVo3/XwEOmolhwukpmSHrQmEb23pwYkFNv5
IjD69cPQ8QLM7njsgpDgw/pds6IHplmkhm5GIwm8lW6x+tg+pbRy05kOQ17x2U/cfmcGK/QTRYAt
LpphUeObTAyWMWZdMLvv+6AJ7IR1F+UETqQpSeiFL4g/tlf4ONyOU+8tVEB3gTzX2VecRAF4XCXl
2y69fwxgHLdDBAY97u6BqTDK7+4jBIgN+83jt1a1RuuW7Ws3w8B+eVYBGkZtFL29QeWH2x0h9QkA
nwwXh2Zp3D/1Hvu0rYWfTj6EBLE1UEis0lIEj82s8vgH5SYLE2zLmFrvTgEOCgghPtd6gDvooJtz
/90xeeEgpRB2v0UVZlyvPrVFOjwUAG9OVUEkVY+K4GrYrP74y0UYXBddVJUtD5bGz/qkkxsZ5ZIX
gWY+SEXnMOS7uLWlZP1h8kj5aa06sQfel3Nab4uMW33JNRW54a4FHS7csxUsd2rhov8AJoJJYf10
S7sZMuJFUEYxtQ5L3Itpxt9QpUjg+Zc6M91BDDkl2rLd7k/uIcf7iYpaqsQ94Z1wjnoxYqtfLdoL
5cfrxXR5y5h7jJDkVv1WWugcgfZHOdhyQ/dxlFLalT0WX3tnaamzdoB19kF6Qc3gczKEnEtF6ePe
o8Fz4T/7xMFq6cTOFqv4CzHfnMUIijEW2OwBNOlqhFp412iOyIMlbKCwDpbnglyj14yCOYNvUBUj
aMJWcA4qs5J9QVFLaMvm4u3IQTX7XnozwfmhudQWPSBZImMdhajqkWouID+/pRIwpiJDBE1a0h1v
Qw8v6kuqDFc890Rru08tHRIA1bof7M3XssXLYR1VMl7ropWTWJ+6Uqct19JH5mcVWLnq/u/Y9FDw
KS6mVOlKcGjIi54ASYSSPEPHJyhefL2ijFsdlrHKmFvyL53W/gxqQgofPcP3eMru+Vpu5fqf66iz
3ZbBQjyEbwpBjqMI+8gdAkrWdTxNnOZ0Iyqi7edfNoLEqbTfgL2isIdZeLL9QfFGll/Sd/+9iUoP
tday6JZ7/JVu1bHATLlXvbJSv8CmmKPe82cghyBVq2VqFqehX3RIesdyNZastp70OZYszSa4fb/c
zcvPI5JT0x4VSAx5PmYPV+OH2NjR7LDiYg5VrUqq2Y1uL1BsA/5mkFbewq/ymqHLxGAYAJ21OICx
go55gihmCbGt61ll64wU9uJgPmY8Ou0xGGMk1Ihtgiqvp0Bq63kN6FABtcdmuvU/gOyGQA0z1Hko
5GUqOSNiIftRmGxY+w1dTvEejM1UgdGu2fQnjn1gFaclMrzHETyGvpAS3B3eIaNylO3IJY4wM+oK
7Wv0pYZWbFXR4LXGpgXm/266tUaVNWOdEO+s1+D1SNzciqSfMFvjk9GfYy4qiEuIoHWCe+gvhD6S
whhJhFPo2prz8KI9NOXynkwQKb/qTa5gfcvKrp14lljbBkDAqznX/dQRfn8mX/z7oRNl1NBYf10n
oO/zGAyT77g0P3WX8uCU7GKqToh0P5fC6uzVEiw6a/Ri1D1lUmilLwM+k+CFSJWAssokFWksdbMu
HmGRoCldYIK+QUQhui4gzPeUWanHb4E1lbSyaaYXdHYIdbhcsdV5Zs1VTT5WLo9LEW+s7NODPw6/
RJAWeCPwuN8G+gxd+sm22q7V3o2s0A5xkLJtxsu3DB8FDAI7o6ioWtN5+yNkLtU0oDk7deajFakr
gUdOJy9T4pSOsJ3ZWn0acRDLvzx3A/njahoWFzwbPDiXxVIGIszf+lCG4eguu6c9D7LiZJWk1Wkq
1mNLRjrqMmbifWd1TasSaUgEn8QdFz2DXx2/BMKvZc/dyAprQSchFu28wDGQoda8MIZEmsxuo6Qb
S/OI7zBiWnck6J2KcftE7CUfqxXDPfHYpQiDm6iennf69qCN5CZLK4u1zZgD6bQBPCV207gwZSPM
Hqgd+2H8BovEHnkGm2GqaCT9o7z9IUIz0grU7xdQQij3lbVdeiD0ewBPxiCOhOTMT5h2zxT7Vv/K
Ere+ES8JOyMglWYmQmjcd+XUWsbs+cyCHvFfm83lW+W8S0jo6HsBJyyghiQRt3CMwTUVU51/6Qqq
a3dj6eRjlGHMVGOWUSIkEYI8OOV+ekfpVPoAMaUjLsb8xkUAMDN3OG+IeY7BOek/FiiqkIaB2F0I
3Kr2AzK0jHSHea1da6ptNfcKQojHcSW/dsrMy3gUM4FjFxlQLRZEoBrTNW17xQ7xhjJU5syXZdW4
Bcebd++3QVMasJeq74KudVepzH9Nu6cKEaenSJJNtUV3Tm0tj1FY0z005v2LeJgRk8lsipre9rof
N/4aocYXERnLOwsC1UUfuL1zektPXR1Lste1hzu8uc/ZLvdqwKT81GJxqhYAe9mMOijuGUUAym7v
D9pzGnk4dS6EFFDInR9QmMAtgqLX/X/q/CGn8E20WmcXZHtjEQUXfA5KcwdAkme3T46MeRMXT1kH
t3JlmCDLCtBH8w22iI9a53oa8wj5jmXabDenrU2sbsvdj1pGBx45lmpjrWcC6vu+OErXpGg8HG6K
yc1hhViOVNzS3X4exYR9sU/rdyEPoy71nQPmYvJLMjv26S/gXzbvyLnNLR9aL9/NKfQHcG6qy6bF
Kbg0SFddWNk4/vTuS1qEvpuHBg/xNNdbXIj6I4vRLjtyzBa1WvBf4PHW/g2zkhU0l89qksNdrB6a
Ze+fCfkVwZpVVlL6NyHpZ2E9A2FgKiuoe5FoDV0W/BMkIUBJgF7ElVBcY7/qLK3UFFpc1fpy3id6
Gfa5aBGXI58A+YUHUJTsX0fH0q9vGH//4Db0y0S/t76mBoL/amfUG6ot+3eKryCg5V/cyoxC7NT0
5ElPjv7UbPZmVQ5J7hXFXJw7Kmu8iuUx4f/m0YG6uV86nFvA2BaDrWzdWm2PG8Rh1jF7Ebx5SQBV
SK/3X744zfDHwgPxJHX36Js/4+bROonhhnGmJX2K0PRg1iN80+Le0s0OmATL486Wn6ig0EsvWN99
tMR+H7Wa0yhWWJoKLfxCBZa0ecaFhywKvhO6y1zc7KV3JhgwQ/pn39nyKN5s4Ea1+QPO6OyHoSDm
hcHYmS7p2cGiTzHHJvws7Mq7D1Bos3Zp3My5Ul49qzepQ5nj+KlpZouauuf8m/38tq+sCRMpWdn1
LXP0L/KaF+HnwpBhnRCDRjVZtneO2BpYVMr4l9ml9bzlM4FeF6M0QZ4sZWk1z19zHi2hsoAY9ILI
PHqZSoSVFZpkvMiHuIRUfht03DaAW6Ru7wXlIe6x+Mjdue4U65lmY4eKkOxTUYIJndA0Fn9i12H/
x830HbiAcyfB/kT1+90ptwFEw4fw3Sdhod8KYa6HTv1mxZvZDdgg2dMxisr4Jor2U82mi7Rlrl0u
b2zlSoa+f+o2L91W5WD3gpdS3tomnyw+SfAtYzdG4acvSJw4FddO5aL/kR4Vjabf8TSvfp+NdyNm
4b1StsDO3U3izPRaJSD2eRqaoL0vmiYIhXYNvM22HIDxOSZxsr3ifC2NKbxBtzpGi9rrhiLrSVl8
oAb9MPc7lm7B/O8vBWnbNtjh918+O2yD6TbDQPglW55nbp2bbm6jFMFjRuprhoVIw+JKITSF3fXY
tMNmBFerJgt90atFT9Lt/4ZX3awCQf9HtlBD429OIvXRKizdVME/b/S/MggZknqVs1stnscPYz11
7FvCjRpXE23v7McBglkFc6Nwj/Zi67WCIKbBcb+fJSZyJPEmeWY9iynvSwE4m80MsrR50vUWpGOh
jiKstfFs3yo8eNl4jVXWhaqijvrYQ9Ic88sAE6vS54uVoFDIJGhRyeZeCSqj02Js4LR+m7M57ZCX
4npo+zgpCz/gASPW4k5sEquBQV9RkOjdnrCypCc9ZtjF6Za2EgaPUmuyJU9rMBEE6p854JaDo38V
Mh5zgjgP5MtITaHREbfCXNChuTCZ0DoJksLGDMOeBW5tXesUpsOUjZKDQSdvwFH/lAyxONIOXFHL
8s+DUFwyBF4V8a07zXfRo2ZZJBmTC+3aKHMB05MelPWkF+U498Jm//YuiKVBFXa4ZO2Sf9OuvZbX
189b8Hu5737oXwSzqwuqUwSZdHp1fhix9uTg8eIskedcEwi3oDbJ+YLsI43O1UBeH172zlTI1ysa
tDABPksIoVeAN4SuNT21PYYo1bMhKKswTYR0KcNJ6Hgkmr+Q5vH5DWnZoLRtqL/Tvnx9BQZgq0BW
35nMfTa3edrWxYu/VwG32WXwG6nooSSye3/IQ0Oytt6fIGsZpcLYOeOk7YOsZOkl6fybDd/bRfM9
qg0R+6D2wjpnliItLmZ6Uzv4Y2VBd0U5a8QcPe+dWgtvl/FbVbrdBo2YlLqwkkLpwFpryjIcEn+w
tDQtORE+GWApBDxjgWwtDnfIqJLhJdFxfnmkHVwCLNt0JLnKvMXVDHM8zYZMu2uX3/0Nfu3BprsL
4eux8WbT6vXHhL1ChVqodLSwTpvhdrm5pjp3K4HF+4wz0tgGA+p1nz8GmKz/sN2UgNXP5nNKdJz8
z1P6ZDZLDVIWgIyu/XCsMHkgCMJ6kWfuy3M+CKo99+al37pmlmFxtF2HVIEzHl0DtuXY6QOe4iZI
BXJo8lHAV9n0M2/ETwS4lHIOV1sI1XxyOtGwPdNMUVkflGzncKQ78aeskpmtrJNtN9PouJ3L0/4Z
ObIKsr01YARGX4tRpWdh92mUI9Ka03bj1JRqEBlkZaFWxFYW3IDUNCTGZb+qGHuv2OG/g+X0Li+f
qfYU+HEK8eX4LAyv7eqnMy/FO14eq+GfzUR0A3J6AiSINMbBEUqPDlxxpzDEvGhD7fiVZowQurQG
Q0Q0KUYs21xWprQnH0GX57bG07KXZjMDipp5IYZo+xsAcLUZnsAdh+jpzLK7oZS1XfR7nyNHtXi9
7ONHzn/x4HY6zBWUZ4U/heaVlX+Om7ekEu/wg2lr8p/A9lycYR5Ymo5mprlRCkZ8RDa6fZ7oJyBI
ucAHzNN6+lkp2925IYBitmP2AhZxYncIbLGlsQbmUp+JHPH9Iu2QYkig7W2WhIwHYeGINIzB8R4i
bASSP88BWsS5ykslpPhuyBWjfZwCL5l4JOwOzdBXH7KjLLo3FJ15k7tmBETmYpnnlQ1jmkfK90pm
bJ9tuNmXcyTZQ5ILGaV3FPx2BzusTRUhEEA56mMHBm0VHaKQxhCsf2GP++5NT66G8sx02FUCFyc4
ICbMIe9p4X7NcqfAg4pdBu5eiA9mgV4BUvLRHRNntfh1ZasKEfYhgwlSbvwut+kBX7JYKNammdiq
GXM3PwsX3IDInNt+XTjKPBIwrZqW/ymQYq5vM83l+MqlvKAcIIiQ9IXkfcpfD/zgY8Fo2w9p8e7X
wbivRccesYXwWzDU9TnzFQL7B+d5NUWM8hx+xqQBB1M7S/IfqesSx9bFlW+iFlOA6uvuY/YLKdYo
km2u6KsMYUB34yPWbydNRKHlJMc/CbW07wR3Qnkk7r8w0ApGkNZFdKPU+4WGpv8fXPphjiN+Y+Sp
DDFaPhmMf7Y2gjWyCx2mZTQvoa6bmmfyz7lG/xX17YOnnKNnzuLMKyOn9VohKd+fUTlrZY4VFhuu
9rxxrYHqbsFdRVNP+hTppxbCYeQrDwbpjIIgsid2rcrqrpRRuX308Pgr2VRu+J4anOtP43nahvJG
0PNgJl7v94XFBjKioPDMQYAm2LCKA9xXFKkc0AI+2elemFyeyLAOo572vzKh8egWQkvvxF6NT7pm
FWbpwNAuBRN7TkUrv59kW7ChZ9HS5L5RdC+/7/6CZjubDCzM4k2iGDNd+qYKpghhBR8DWzcg0Akm
n6QK8LuRw8SBbcDo9cKobFRnGzGwpNgHr9s3zi06Bhck9YK3DqKqDYLSgRV9Ier0b5PD/rsfqMXS
zI3U8Pe+qgQQzkVwnrZlQJcYvp5kt0HSkcVNY6DJwJW1pa1DHXNTojLNl9GK+W52l4nn9fv6ae5t
of9fwviMO0Vf0CK0xbWsqb+A4BFhDVBEHD4f33j4T0qqbjoS0a2wXykbJEQ+356OEj0VVvBYhcw2
mlWkMNQx+QGN56Mx7R3fLn9tDzmLM+fERn8gNQ3BABaSNFHK+R5hmV9o1m5ubhYM6fKDN5664gpa
2ybEnJVqui1vrpmODlpdo3HQ4SCogQbkmAz1+s1qOOEtt5jFTtD0cCL66jj3NFSptzC3xEAuImyy
G2oJ7jgauyhaESJCIVk+Xol0L7EJoePe1zHmDHKUlZD8n7W2F2/ARUQKVfyehFf9ej97JJKbXoGd
qtKkwuTYytX3k63BiNFwctqgZJCXjccLnGI/kPqNyg/Yn8QMlF4pKLPtsLk3tcuc9lxJJHepGFO6
0jFv5ZVQxybW3DY2XcO66TKO4otilT6mBKhgXiisd8s8dRbH6lRMSfykKO5ydVoA0g+wpLdBvNPm
g2MQkSyO/eqMjInippyuvZIGla8gZD1kBdPddN5gasyQTH/JAbRwWCI+GXEtfOGAW8hMjPG9kbut
/onF+FR0UV4mM3cK8Cjed5QznBcIN01bEZEpF7z1u4KJ9xdieUYT6Itum+7leJnJWfEAqNjlHTLo
IxdI8jnb+pQ2KJD/VV6RvXD+SMqlIcl0+phSGMwt/z/f4LS6BjjYKKbOxlbW7M8PBxS68mgPG7Y+
hsEO+kKUixKeGF42MwQers0wMUUn3Vm5zVMbYA2I0uYkw8+1UxsDG9G+pB8joHmpLLt9wWMgqtvo
nxQdIze+fcAqmUqBY+D/ptCZrgjrmm/h1QhRlpdrxa8EUcdYd0pFIoVPqY5+6Ed54Q4iWGrerYzY
Wlih9lLzfhe5+ftzY1L2NoSTbqQmE9gHPTGCSXAp4AHvNFtW0lZip2F3XyPmWYbrwS79U+cJtbqe
o2StFbN6A14E+bU4ea0CReMV90zCMtmcNOpMBZOJdbvcFjC/Y8G6AwLynWMLv1HeIYkAA2mNfu2x
eIOL7IGW/fdqRtqtEYA3RvJX0uGJXzJP28BGmIeDthWIl6aQ08s9zBJD/iyrJurA2iXCEjzQrGEt
R716eF81IP8IE24FaUipkqDGogAlfy5BVrOt2rBoULLVdytX7ycKKLOTwoq8MpDMtUeQX84+W7Bw
My9KXlj20hSXQxIdWTyAXf91ya1Cr8+pULu89AHPQl1o6RC9PR55++4V2cOmNMCbW51SABrfAEjI
nYOAENopv+eaoSG8rIMBnsBDouc34L4kA4Djud+lmWURDhWxf0uhB84Rk9nO4ylUWx9C140kyZA+
xMoqn2sLWWmu29u96FFysZjSfzLO93pkzGclY9TRK45Sub5xffcQF6h3uX5yzhvOUgeZPePjY/GI
4hdC8x84ANN8npG4i5nlVSnx4f2dgGVaAUkKYcIvyDrwSf2F7HeujralOQhpk4EN1WBY8e04VMOh
TJ7bmVXxHo5wlqD5ukhPS5ryl3U8Gk89EaAmKHxx3jrYV91auqyTGC08dapHxqRRXCI1YfqUtrr4
RumiAoB9IQ2J41jFWd0uIQF2mWeta1tu+9AEQaB9y4d0GSM/+CTVZJgrLmaNbVzQgXSatj9pvvUk
hVstAnUCqn66zKxkwFQvBgkKJSalSxkIidFY2g7yByhLw+2VrbY8xgrhZ2NzzWB+LsDuyz25QY6b
I4YaHxe5JTK9EhBJ2mN12B/uaeJblWOoYlTtLcwLb5qXl+mFOJUnbz1NPfxjVLEOwwfiPG+opKk+
0gU4eMOzCeeeASBOjuNCppxYTCcqxhTFv6IW10SQHt3ziXNj5qdNz1ozwTye/fVy0E5CX/nPaZb3
GV+c0PpS0pPyEn5S4+5WsneIcrbbpp15frhRSwOkGEgM68GK04VhnzetvLzI+8PBgk2RDTnDOnuW
7wfSytXeGdbqItWT9MxwYsUVBMG29NLJrSG7o//CEPjU9rpQNbFmVkhUqOH+J9JSWmK4aHuYTC6G
7GwwoTuINiOy2dlGxobSKSngyteXDozUVbYniG0jSeqZr0jKyl6vylAksJP6Da2Br8ELtP8rsYKQ
EjXh1TssYgd7odl1Pirht0ePo2Kj6cezBLvHrCKs7L+9u2Iihu/wtvjWC8F7OXzxwdawPT1Bk1Zp
ogqcHWr46Z1vMknIVudUXOU0EWAaNby3b0UZ03Gu7CBf+eOTrYKrnjGMyhNLLKwxYGNh8srMfzRG
zHM57neKs75uT3zQ3LGfVfBoJ3giCQ/VngJDvBGfONTv8H9FvmyWm7QWe3TT8tZa7DLwaBLnd4bT
wG3sihIE+KCQHV65ab8hSp+xklOFxZa6NnSo9F4HtxhOO/jYbCk5M6x9Mu68MPjxPLAEW6IlyhO8
sWT/bcVpXA8yjFvRqe+Iy1zuVzmZDV38aeniVZ2eUB/m/l91NdRtQLIZ66F+HLgWM9K5Ec1hlnFt
koJZJdnXPy4IUxGd5nbGGhXCAu60ToPIwgWhlg0wZYqCMsvK5mHEC783aQuEpZ/BGKGsajAUTzA3
vyrR7fWoOAsFSNpDhB81yD0JA8dvqZH2IBPH2epwJ0DEYqLo1MsObNriOtxeBeIKX0K8di9N4oAi
rbdoEcYGVgsIG3HzWsxHikIkDG8y1cldSqio/4uBCOblutFehg669LdkBbJTk96HiEC/qIfM1Xsr
FwaJhyVUNoVLQYujz2xsVrj2iqI5iYNiDaooLbZOQDYfqYuvmOdhtILPUzVHVXWaZ0bNW5LD11dL
Lj5g3t9tIPz7f3jvrlcHFy621qLdqwYh6WGTAPe+juA3QnQsYt2TZC55Iqy8ICpWri4GHpx0RDWF
40E4PKg7td/IcIZKux+zhO8c4yEruTMilhjdVhiwE5sKGtFN8JRfKx/l7eFapAtqVdAGYahpHXfg
PH2opL5CBBerPVcAfUnWEAqXw1gQwmMRURltQGqSaEd+qKe8FJY7ISVpx72DEz5QZ1LfPHVP2qZ4
WaBT9pKYbJYzTY9d713fKY27y35VCxreGeXmECspZtTjlO7Dh+4YePsu+cv6pkMnJFnnccrEeF8Z
YyswnBW7ed6n5Y545hVP27MrJVG1k8bQdJMuXe/DRcDJT+Z9K/e63/H/NQNDPnusjIoLCBBfMP0R
8U3+SyEFlAeYIY6xmsiCQi7d8pSeVq5yiMCokvybNFdSUsBQVg87tkh3xWKfxrkJhhxgRDcobBM+
I2wCG2wISFDpkyYJC/ppj3cJ0ie81xeKazbkl4CaUGFEFv5OKC+I0fHwVXLQe6rSAUpHf/i/fTAr
WO1+fYOxnRihm9+3SRFedrWySIJViLFglnoP6y7QzrquMrOowtUaMqNp69tpuptkVePa5pbdbQzM
76EcknKxiRzjyrC03qU5q+feQIENxeLGpCWIT9XeovVQcS7Yvx797JX87vcwKxKeuHC3IDYNonlY
4JwV1arfEKNVlrqd81MhdGdAqnP2ZlBqhIh/qQnf/R9aCGMnUiWTO46lPxdPrbt53Q/OxxGEpaNj
5MJQgkvU/BB4brnrUFzobu9c7LOZ+sQQTW16jpjwgNfO1UJO9pF0zvB9uxdzQrjQhRv8+UXmkwZq
maCEMVrIOSvg5tl2hP/UB/cckbQf2GXG5Zyx4/X7olwFxPftc/Et+JOzoZCHKPlfgCJIz9VQ2kGd
PWtJ93ynQqTCqGCmHvWIN2+TCtLGAO7JI/UDKpylXLHZtvktUfqGnh6xPiVWN1MkZMRI6ZRY2xap
ygbRk8vLkXtJxfRukCC7T5E10oOwhX1DhIQ60/L53OemVhcoA5I/T/qP7VhUKpVQusUo5Wl/6UJM
MOpuIqO+eREA1sfkdIxWYx4E9e2KhTLsO5xfrrrV1eqaK/97ywJka7VI3CQXBIGQRafx2bD/vkKS
bovw1AhKhh1jVAVoIed3G0d7q2peltNJmqGZGNxNXOrT9xCFOCGCMYu575k8oqi25acZmKvdZNaP
+5U7xxczXIty8I0Awn9MiCLl2hi4rir10VZG9JvfssIe+TmCgU/jGVDLftxmY8wlfz9zF++BKZWF
8ql88lj8yHuInByopWfY4CWAhX/26CLWemoiSTdz3PuosMUsxX9qfYWbOow97X+XhQqdf0Q3aEDr
8nRYd+0CglqA0/ALxM+UW8kPLBdgFjP7ZTYTax1Y0/J5x/7X1Dc8bynuxzHflsPYolImLYomlSaD
+QaAt2Hct6aD7vgKwExbv9j4s1Oh+IpJ8wEQqquhK+1qlV7kM4dN4CfulwN+cCxJlBvp+V6w7wlh
Y9k+P3g5XoWUtqk58RaYK73jOUXrTZDBAsA+pxBvrqonMn5Qh6CHlicSOTgWBgD4CRmoiiFcyOW9
Q6iSbKXW+w9JRnCjbZx7eV9IRUiXztEmU5Pakj/2kzZeA6yzDViJtVk5lfQKGKf6fjT8elZbzPks
ZCGC/C8k8MNV8TJdDrlA2vfXb5EZzw4YwnA8MreN5l4XBiecy0tK3EglOXVFlhRhtIe7NyaY6Lis
SVRbzhQ/0NO6domvmQBpJ9rYNAptF6lc4kNL5SKY6sINGBkcFrPVuhHYk/UYbKaY0XQHRpu94J2f
a2vxRisYXsr+hK0vtL9stTM4QWLCXeTudREQte+9kJo2JQ8JS/0PVI4ReaD+XmFFvyHklRFP6/ws
WzW5rBrinRlq4tgRhTM9avsPHYnCYFIoXa/UGqUogoOU5HY3mVSvRjAttki9NuvupzWPRDJdSK8M
oMkUVVA+7wiZypNzSWh4IA1lYXlQ+zXD6FGu2V28Zz84exnNNL5xCDs13le4JEEC04Qb0+/wQoQM
EqxT7os7rTPG+ztq4+pVJIb1l1vYsMfJ1zJTVrAcTd0I/g7o8g8UvXVsndqEN49Fa/UoUw2Gq91P
drDV1bdyknHDViLx0HoxRi3NWjgXgRFPCoAv2B0A7jbdQOqjmW3krq0QRHZfW31tx+aRYkMDk4RD
bLF8d/Rt5SDrbZ5J2k8s0J3gYNzapQwDVA0QkOoYKoDzg2ai25LwyiO0Z6oQpOaR4ILzsyCPq8D/
InnqDe3SR1DcdvvCL9xaPBI72BgV2+oSnIVTlImhQCckrukyukr1l5mFcXM5zlQOVFKNKbv7Il85
gyLE6AQLfhtdNJp6FSKZV2x6lU/Qiq+k2K2HYr18txF5HGrLtlzwan76IYtQ/fevSLSxPB+ZDxcN
GztBlV+AGcmJAmK7J0qJ7H7qKOurKAAt71rrDhQUz++Tm26OALJOsMv4L7kbHINQPbB48OsPADcb
qIBog7UH+x/tzow1FoByZpTOMjEOL3QdG9UoAvZJtfOy5gvWWhK4XvG+cE3CKBtde2m1KYEVv1+1
pI7uf2O9B6QHyWrrlyCyBmWUTsPu27afuJ0g8ZbnayPFmg0qleKkT/JVjzT0dPBC+fO1V2ao0HLd
cCFoe8ZHDVUo36WnUHKLZfXiVSv5HPwsoA7CUrdOFfeLy3ss8Bgh8sPuIkCe5PCcojqK6X6A2n0j
xvWvpkdXD1D8hd7oie1lLile6EkhkmQTalojFO/1I7WHF1/pPJTZAH9H4qjEHbyo+UPr/wQNFtza
ssZ+lwh3a1cdKfW45FC5v+Vu3BBsdT5mSvZ4Kybo/q7Th5SHXldIUYeyJ3siopyVPyE0rofOvPgl
/BnnFYRqyw7gHy5LvLkK47qW/DhMz5SfyLUlfaqt8QL9Ncak2KwfZABeunPK8xICd75voUoRAE9T
9KF67BCxQKRIVx5wu+jBWd7QQj6iP4B9Zhoe76HaUbiJsXGXCR39jGV45ugTFx7Ef5/gNUbfQ0A1
jlFujUM7IO4xLm96zb/L2UENceVkTlveMepFeCIBYaJNLemDkT/v8FzhRXF86jvCHYdrCcnGwJmo
l2e53639R3NQHIvdZpEbcu6JZMkL2KiaCQJ01D1v/2yH0wvER4dk7tWpS+aGP3rjrgC2GxMruBA+
ajjErrfjHcm1AIFZtlfYc9dEasQLOYK3WrF/vjHIccos/0DOn7KeQFzI/IOrjHUi6NFrxHA+SsyZ
jUEXniy/pHuxNjM9Hsv2lsbzyRoFkWVuqWXJ+7wU5TIF1NOltTgIKT7pK5E4zKJHyECwFVxj3JVE
Je5JASRndUOHDkbPMffzffM67aSwxP7unDeitFqAah9oQliLv7bP54J9cCO7mKqJWpLUid1C2TsZ
xWEgPvQ+BMx3vwwn8KmPetLt2bsEIHNsCT/O9vmyEBER45neVuljEbe4X8kcQRYIZy+RIRk7p5SU
5ejTOUYZh+p5+IDV1qEo5eZDyLucAGYVaF/C9ZfBRzrQwfifsbd6JfXW9fYSZe2NWsdNbBVT0mmS
R87i4pIaPYpzQF2BLaF1juChS2J+HiF0MfSUxEJ0aSk3/Ni/n7xhO6776igsPH8pJ7wTIoj0nysd
OCHDb9kE1+GfO46tY+A19q6SUh3I55G7b+24/Q6FwugIDKJry9Gw3M5+Vn+hzfC1FtkJ6nVKGrXJ
cdScA2xrCxZVXyS97La75l5qKgNeg3tojqfLgrT160dwoMZqVZ3/MdJZMtPJRq0sors2uktrUMIH
vCBMm7pQxtCp6w7zZjZM+5Pcz7/MSp5HtP1d7v4u2HJRtlS+iv6bLBbH8u7sMJd15S3ba7iuUP6V
ip0elnDpT1lTXCAU6ZOOqT8IfpDKyUNAo9b2v+lCjqOApBDELIzwvnQFfTOq5eevR9G/h3CBm7TR
yEaoTvaeEv+X80DU/79+2zu4z2OrNZ/uDMg3hjGNg3uxoxBaNYB7w0kQ2PIWHMJzQwhJGwCFcIDx
NquzfAYWqj/pxslz7mlDkbZOhJxar3T0WutSfnO7o83fcmVe5bKtVaecIcPbywA8wX0KkGFmFNn+
VSa3JK+ivwo2+ruMepofesxIVknNreweLQUBv1ag5G3bXsWIWqYcfLMewY1ZAeSlEFbsJhuiPVTx
5ue90636YoX64KBm8REGJQf9AXsiURCywJRtaxVHS2YCSOv4UUOipkIcv50agT87shqZ6hJpF64Q
ilkDzaLYwJLiOwKxYT47XTIXGWz3MnZbDtFoLI8uKKg4pVPueQ1xNa7SeU8FGjlEqlDIlD5e5ejd
V9LETMfZ6C/vbptAI0kp/9ui/T7uehUipbgjBFAYde70M1YuTV7oi3riN4pq68qBSCfvw7br/Dw1
kqSl12tJ0hh4bqXynBeMZgJeUyaA/Z0Pik0mEYyCd6IZ/ButPek4wua9dvxfDy6gp4KSQkxnh148
LpISpVF+YRtj7iDWHmB33yyGWA2XRW7zMxDOTO8why7fjmjmiYjImV6v6+d9lpb0G+WK8C6uxNL1
XCMxEz4s0N9A2rVj1CIX0s5jrAbePRdQEgfcpm1PISh5MWG35lArlLPXap5abm4YDSLChHFeQa8l
Gl1WowyqBEv2UEcP7Rla3jzB/jqdpBO21vGpsRiHJlbBssRM7WuhAQj7ImlTKc18IMtNcsR62ELH
LLOvRD+NQ8uJuK5ufKO5Srq7cUCjCpoQjepqty+xNWKJ6GgUsv2mbwKXFuWObumjefgj4jjOLz3d
hvH0oTMRRLHIqH361pS9gsvW2UKQChC4rlWXxTHsz7fLn38fqE4SxeV72OHuTwBumtDijqjPdM2H
XzKVU+q40VzHAwFG6ZOIh45KzU9qRBTp/z7rr/U5OyxsmmOG5eBbeLGtk4eSSGWB0FD7Ms9Kzujn
QHYqlH2RtVtPvIy/i1Nol1DzAhFIidMyaCWFjEzxJnpl/EcGDKPgq8u/KSXII2mEZeKyTQFGZ5Tj
O+DbHZ8ucZjLkKn4vHCcBEkQQBt3e4gPJkyoPbf0tXKICzZPsEf/fGmBrf15qJ1b7mH7KjhsDkj2
cZ+Bcxquxqutwf6XrMJxK8CLvUZmU51N7afs3LsACD+MyhDPrN778IcSKEfxruHJNjjUJrSf8mzV
t1AwQjGAW4kbiidJ+Epodds8DfdeSMwI2f1b8xjsL4YIZPuZ911aKsW7VoK7CimjXXygsGEfDHdi
EcYJIOT6Fkao3i3zvGddU1ubv/KyT5Rvd1NVXh/UT+9YNJOlv6IIzWO2X0/g7dJf3B4HAg2T7/Ov
BnxfDPIl019TeJxoifbxWUpLfIi1hOwlujYjZ+c7f9JCFEkE5FMJxUVFkhnDOOIIU3U7YA5o7ulI
Chi/7Bv3j7+FmRWpVngzlas3XZo16jxSbaRWH88yZV2wkr/Ju86U46c9Ai/fZxjj1VrO2o5yxntP
YztEg98PneBsFOsYtpuYOFePJyCoIVDEJzhoy031EMDVEmHlOtqfSiUb21XaIDyJm+E/7/7d8rlU
wKb4pbSeH4nYk+ads5d3pYK7w1wnIpZWhvctccCH3zkjenkcBGkbUlUdxiGJHVOuf4mDR8yB6Fk6
sabOPmKvFEYw52EVUeKX2wPdWoxOLYbN7/Ph6osyqIwbNxPnc51q7BFS4rMk17AAIVx9eYZ2c24a
iHrdcF+vsW2AHhvJp/6AQFZqO/axZ2hNqlV2en+67V+cjV7jVom77Dymv8s768qg4H894kdM84u7
d3Ot/ACDR8uZlHykmbxvHM6zfdyiFJiO9GR+8X4yq3YGrbHVsG3XzFAVFl9+lyJ4D0B7oXEeP975
vFHB/cMJaCbQvgL0kBbMWsTS9DC7kUxuGooiVhNzVHsP4pbNixQVfEthSM2c7lpSIlupy4lQBN92
XmV5aAqEQJSKoHBwQbXrIUunXYMJxdrCBU7hSxU46tsv0bIkW8Mnphu8JSIP/zf2QYLNNeKq5Bes
hhoKFAQjNFHU5clRn278WmoT9FSaZ2u0ZAxdFozIw4gdeB5V7/HHjg6p6oQLFvg/9sS3M4QHGCMf
nrSLgji3W6zGosIIUj4W1yCODkxeRXF6AQH4STd7NhAnUNonLWI5Y3mBoCyG029euvAWr0CNzFCX
/5n01VUTK9/mYTe5btxAQoQvRWrxMas7HkBQ3Lt8e9jClCyZ+HzWixMi16fttmV4Clkh+RDjLuGy
hEZknK24Sp5rOkftKVlYPVnAuRW7irCP3Zmj0fYT++rymg+dda+wEXkBIduQHz7VgPkAwy+5d37+
swcfiQborFh+D0/NCuM8DCpxqtcTCWjTA9N3SvNWor/XHuRiXmvdqWmeW2sYbF4jwCXkc4C1YDyr
bMJzVfJfNsRNsc373jefCn7zf71/ZSxTfM0ljQA/tKcJG0cOGBBSas8JVX4Ehkh3yRKAXzCsL48h
GM2nthwwwPoQpb7DW9v77LK8QBi/pJDkhibtvr6DtkYMDlJGuzH51ef7EFBCSnTgWVHe0zKVwL2B
dmkaSCiUadvFl6/E0dvdBOSfTCDuZS/Am6X87+zGpz1R8EdpzHM4auu4Euid+LJTHVQDFikQLdlS
mbV4aL129Vq0N8Uhghb5NFIpWgO8bzfGB+nN1Zh5Fwjq4pKlqXH55K2E/QNyP2dEgUxvayrrnwGt
MzEH2fADCPlR5KbWN6eH3bo8CzeiOr5URf4tOsWAy/jwUKMz33pTzNLgSxj7k1cDx5eC5oYTUGhm
eM75A+hYXxWO8RNxHzEsoh1I1Q2kKraxvsSPMkMM2SVd+6ORgAYSeUcOBXp/+VfMkHGMnnZIt9+i
rZG/DqfHUy18xp5HSU8Ehq23hW2wP95ggjtZkdT2FM2Eyp5ROSLapJap2Pq8oU2kSaqf1oQDwwJp
z/jocNEG/d+HpMlpUZIDvU3FXNPra2G63Z8yszZDtWibfu0SJGHohi1oZ88RG7LuunmKYZUNncQL
s74iJohkxUVNSoYBCKzK2XctFPIoqjiIxhAmOYBQFD06CizF9xBMYgrEfJJZF7RDHaeaC2qHBnG0
GjSBiYwyTJJZcv2rWvBkDXUMip76OAyD5OvMGy+7NAlJdxIE5OpRKhVr7j4Wh8o+gfN+r+U4NFpT
7TybwlkJt1vyG+ys00tRp8Pu+MfUVaN9as1CR5j9BigrGk+88MrfbvQ1FS7Kt7kfcbqrLUEDdKTI
G0TgA6OZMdn5oC6i6zV11k1CxASb/vqIV8RGo6BzT86pPDtSO9kpNzCdrGu9EdDFsnt9o/E1wMC/
ZzsreyqT9yUl5e73ONYkn9dWi3YxWCE9dQgpNJWU0XUHzCDcxG7rkogZbARw0EcZe8h7KysAwvXF
olR7+q8lQQLPZKffatOMKZ6hynOrL6s92klK1PvxB1RYqNpAi4Jr/UbS9H2L2WVvaMRhmHLjhShL
klz7ejHiPqo3K/Cp1dwB0zQn+TMTZxrA5QHzcBrPUH8V5SN5EbcDrP3Lq7bg18I0fdnP/p2anA0S
1lYTR32jqJ5xZWC2JoWLkR6JVQYqx+6/NwY/HzB3pQTsRU/S2soQJNPneCReEKdjggV8GOA4T01h
fOLjUcc8qkfJhNX+rvv1q6RiAxpDQWEpIL1DBztmizuhjWa/58imQK42woxzmeX7aNBZxmlZhK1G
ZPKAHS1bN90OEXNG5Pw7Bd3YH+l08tS26t7NpbLvMuQSbQPp/yR6M/nmw5xb9/H71pGGWtJuzNMO
dROOwvanSlGvY8uWOYrp2lemlDwd1vAqTTxIKrT6h68UAlxfdIRBAKtsu0r9B3VwVw1kEtKPvlek
KomwreKu4+sSUa30F1OrJR4HWjx3dnyxQR8bKqBAhF5WP1Y/q0day/Vs9VdaNWq7lqjk0d3dOlHQ
QHYl+d/t3QStbAtCh92rv/smjoVOTeF2Gb59aLv2Hbk+SjiSrLBBfbmPMhy9mP9gyvvxFuKrvdTH
oHUeZxc4t60Vh+UUn9bmMTmaReAvRnI2Pi81BSRcxYwm7A/Ez7b9//lxLQy5Abx4EpeTzvBdRU/R
wV4WkzqBxyiSuJ0Xbfp2jhgGnarZ9tUrrfruEBK9+uzksoBYfZNn6iwB3enQhnCyRlfw+UGR7GVZ
YxcrJ3qpMePC60gfHqlbxfm8+ec6Ilwmmd2KLOFcZNSpsF/5NxvC6N50viYw/PJyQHBOC9Hw5qOa
RfY13JP9jdYAwUDmsb3NfZnjoDCdkOv4bgLgWqyKKgnM4DrIxg5/MAgQ1fTWOHVBoDSP/TVosiPT
d5zduvjlGhO6OgwTK8rR2ZPtsL5Du3gKY2hYlEVbu7rVZz8W+fpuOb0bTn6F1BTDMTbY8sbkZKr4
Y52oWgvZKAOJG75ghRUvSQ404k5/NDKwybanu26XPyMWNi9/8oWQWlFQof8JDPpJT8hJTCCH0+qS
ve5KPC8Odb+PqInv5A6fak7LQJmQp/N/QvMVsNWxxQmOkra/qUNza0xzYcmvWmoMOYhbkXZlZDt9
oWgYWQ6MFlirmOoJQ/DHYoSzGDAaatKe0IlXDWjlItp7X8DszqLtGASDW2ExArGY5hqW53f+Gi/A
Q6fjNRYHZ0em/UB2ae2J1Hf0CF2/1ljPMaXp6hXXf2rKcximOAM98NqtIg2B38hRs1QXljYTwDhi
01RQCEjWXaQ5a7slEh0+D+JCiWuF7a6Cy9cffqbQQTymL9vIyTxjgZRr7zAN9coWNP0lKqn8y4y3
W6V26zhV/a8DBJXg82J+55uCBKvRtLyFwmE5fQehstaPlWUFWKfSA+8Mfw+yTXnr1MsRJEDOTbBs
k7EEFmu8NxgD4Jkx0lmRdl835lbUoxTOA17vLkNraLBrcYVIVW2pZMTmaXNBD27153xnvZsKx8lC
Y7q+IRPVCYvZaPCs2lIPunKVYwDaEV+NFTpJgZTL615Bwc+VP0eafwWyogRG+OXKC5xhawcXKInq
sTyEbiP1UYcdCL/fBHz+wc677vC8DKckcwsHXuLDwxSBqdRN8dCrb1ea7HhJw89ZBqHY2EpGJ7vV
fmqLAYOvy/RkqjK5sCy2g/n90nYvXyOd41y4A6gP53cCNrrH2x7CILeXB/p6X33DtwPGWIpacnFq
bmI96WrutBQWioIUM2ZX/qAPIJeQpInDQlMiWE38wa0Si4KpDPGPYi2Z7zM3GoXKFErDJ5tjjTpJ
CYosSQMjf5AmgtgGjDhHsxlVvoYZqUvRtbedc2fty/wOa4bXqqyeagvJt2UcZuMelKEYBNyXsIn2
xYsaIn4uIt0Fk32/hd97C/QlegO18O0eDHN02cVTleCFNNpGc3KwxBMXAPlh4okRSVIKC7GFnjVR
7Vlok95ZyCzOfraLP+kAEPVYbI/zD0W0UPLo6un/cuepMxlirRdgS/HJzkn3stUbI6FMZbp70WkQ
B0Pzs1dYZjrXyo/22delQR91H5mQrTnRrKE8sfrFUcXhuIWBPGYaSPGSV9zneaE7CJioBotMzan3
w66mwxtlPKSW8Xj5aEh77+kYgg9eoF3XwB69aHzkBhDE0H+Z7Ps2i6DKDkB+gM2XWlm3XIbCxMVP
pk/hLGrnTBPT12LUf1vvlVBCV8XTMY3qntl0dmv6UTbsiZEYjcdrth13Bj2qcX8mst5LRmBZSams
FQ7hwbPNiKi6lb+wOcU11TQjs5+nNPl6W9hPqLaPvAgI8XUBOrFaMN9zxrGJAB2P29X8Azb/oNIT
xk9fU0riZpE84EUflIcZJD+a5ZMCiihP4SJTpSau4+UgKG/NA2aJl2t3dT7St6aWIi6maMmDvUbJ
B3jlwQVtrtb2ui7ww1OasakqmTneHpCm3G7MOD4UVLNe62dCyrUtdkcCRMJsNYxEDyY5rliPsnwz
+9z2/z5DKxNbrzeEJTq9BqhECp9vmrou/uxt0BqfSVuvKQyJ6V+0Qa50A1P9Cc40sj7rBbsZtuSx
Cl/cJup0qIe2WSeCwV7Uc2gGBojT07vBwHiKabFLqNd+WdHTQNfwK5JGadK7nXDXFfbd5hDcmj/h
8OwIa0j39ofAulQeOF2Yql1lLk3KXmm3SKmI//f6gk0gvMP7rhUwpAlyPHQZLULJgWSNCdyZmmR+
YBUkKIFAyFAHYTWfkkrRdttJFF5WekPgByHde6kkSA21Y6R07rp7LSC82j6uyAoiIV5GF4F5pAlc
9oWcvs06llCwESAC+/2nSL0WxBG7i2MoPSJZik4DqTklVbudPzgHa9Af6rhF0jF6oATu7uaPQohm
AWjifPie5LoNxH16t6UvbJ/upjFe62uOKu1hJxqCOfiKaluVt2qrHR+uLvF6c7xZyT1oe6NKIFEw
VhPRnK6CQmFahPSM0FqNVe2kVgPN46pz4msrIjJxZldEvVy1ghjlaDlFw7w/BINPJ1vu84C7hWz0
Mr5GQvCE3ZPWrgkZTD9qrbrySiC7EJn6AhbrTYdD6NJyWBIJ9ULsXaHOGW5aLEe+WSJ62xyFi4rX
HzWlP62FI874d5rerDtT757iMUi7Ci0AnMvHZhrpWRwOOweJnNQoJi8auxlH+Hj1CmQfRhQN4lIq
W2bkYOuhk4xbliefVYN1j2FsSXoKIGvR5CXZ4E4TDqMOOCPaVeYr3PTpcFg4JfWn9edGSqE4WNCf
xIN3l4sON5rMBJOV6evEKQraYIlHKZce6tdX4DH/HLpTzZowAWwMYTgPHBh+IcxiDc1MyrMgfNNw
v5rmPhOPEA8/sv493JIBODMH8qpeakP6o/dmcaqjaCJhVnkFhQfg5ZHfY0UiWVbpu8PsPinGvmJA
F+et5p6yk9yUPiRfUWgELgefJ/jTF4bfiths/SddPu7e17EgKZcpBNBHGz0uuL4TiRy/sUsImmy+
c5Yk8aIDnqJ3sbLXTACCZ76cjhkEjk2gg9zC3MXw/Dl0jehcTEy1+8E4QsEk8DkHdrfEhZU+k9iL
RVhWfmFVaFC/3TLEnoiZ632uThZR1bsWtle/OvCbB2MJVEdidv/B/ApTdy7VYHPf14JGjMJ111g4
xY4iweoOl274MHglq/tcwGzwhTj8Uqu4SVgVnB4yj5dZvEMjOkpOAdssyxETTu71qjTtZDCO5OSl
WU7qh0257GpHaJR6A9MJs9Wbbm3A3ob0Pz0dE2yxkoxZge3dKGKGBLSh6CdA5LM6vcrbxW1SpD5o
6p6wiDH6Wx2P2Yy6ReBBB+4xP7/2Iqkc3iNH3bNuTuGc2JdwP8t1ggHPjZTpu3uFiXMTpSIP2bu2
SN5J8qTPrsjmzOfJ6r9CzEHPA1h8E3s9V+7i5q/FYHFBfFbU7FQ4wtu0BoN5r+DxXhpQ1VoOu2bG
DKbNfMgTqiw5qrKna7dBeAsBJ6P1uzeek3Lw1hbFBm8CrotCKko56EuDpx85tkAvXujkJahBcXMG
dArx/+pYAfv3U/aW15Y/zvzS51wt5EaJc18iJavxlkeT8h4hD4SolGFAbK2hNHfWZEk0qv7pi3hU
H8eH85n6E4UYIkhAhbbuMQ6930kWiK8DglUcbipLav9hIBxoyG94b/7gOhHtULgaPa7J34Uh7U6C
mBgxZ+HyN7WwZwRt1g0goevcW7HyILft9MNYwEUTb63T8hwZbewAr8auqpxqwme8J7Eo3FKWEHcy
ObaY29ywW886N8JnSB3a+x0kucUwQKOc238PPAiXFwZReXi1y5EMoKKXs0a3jOnlMKACO+mCa5No
bM6s4KfHcB4LYcvYosAhw+gOr7s5Es++QDJn/dlU8OmNURUPypzdSJOz0R3vFzIqHZtSEeiqhDA8
vWkHxn+Vu7dh5qEUfmf43gLyQVJb47F1N2iQgmrUIC/p8rjO3xgcNSgT2y6DfvXA5nEanOGM5dBP
GxCnZ3kOJJ4lFmeSgZ6DFI6cRajAPwpWWfHG9MnNKXffYvWEOk1cKbOF5ELc4In0fS0Z4vISX0PP
lYHtQ+jZuWMpQT76l6oolu7Z1nTShfiaQKNoyqrt6cqv9pTZH9SS0hQCFheYshXjqWdt59WbKI1B
eUU7Gkst0BFDu1Be/kfKbUS23+7kGBTbA27w46Q/cBLveohEpSnJKw8ScIaIhJWZ1tLGyiktiQ+i
AxA8Ty/XclbWycpXIEcuxiSGYrw/cRSrggoSEy7Pl0TlsBxf76AOjaPH8l1OOvf3WOxerQKl5lsj
A9aWeOVJYKl/Sg10FFZBEqJPEx8Qf5tvXFQsUKXXOEy70Y5crVYhWJACHmxmbQ0yZUIzPO31jtIZ
8Vbw7nMvgbpKVCA5wOotUm4psfQu67+Jxij+H/ZXQHb2qM75pY38f7eky00JaONRv1TRuh30hrgQ
OSaPjgh9CRqrZ25fAXE6HAYki3NrTiP9benN1/tvWxWEBkdcgcZuQ6FEU+Js+Dc9iNGgviGhzqwy
RSAky871PWNAWCBfOQQD1v5jdAcsXclJR0fXBBjjv2sK/osf77QKxbtsFIEfTdfa92NOlWf+yW19
SCUNo8ph9Ed7AD0FtIhHcMbi8YwPUeKEv/xF6EFW7H8wT+mN4l8jJSCZjfgxYjk99qGd6dEPhV5v
RuNNcMDYLfcJpQoPsAhiE76KK1I9Fj4nWyIBwmY9IoqxxtzHPmK6Wgb/yvmxddkfDMvnJRx7e0xI
8x8Mc/ykxtYGDBNAwaE6n4z/wk284q+qklDmn3vlXZUKcsNUo0ZvD+sgcUclUBwf5Mtmfuy8IRoG
9Sy2/6435CGgf9hvIoe5vJZkPu10PL1H2GoRpVHbsdO46FeAUsHFmILulTiYWMU6Dwc8wHq1zlmC
V3FEbM6GxQOKWDmM/i8C9Wp5yMhdJH9NYv8TT+4pngjJxjTIVVHZ8G549IWG0agUld3fsiXSLIxJ
Atnf5+bfYTRMhMfWWFFk495TeO/+UXQXSYfOx5t1+QrWS9ataoJN/aAzCTJV8QCYFcfQTYr2U/rY
Dy/IcjVYAAWVdhSOGDGFCcyx3Id1WXCAjWlsEmHcL+IVcsmHkXw9AwgNawC3EsGf+s9CLqoEtxmc
ZFgXIDp+YZ02ZLWRVEDMb5vkDn0l31X6UsaZFgVLuutWZAdK/88DbLPbRVEFf1njbZIA7GzzKhZg
fZr3paIIHZFxcRzr4icgG7q2lBdlSMmmFt8qPrejBTK9LPcP0HbYvYAaw8VDBSGdmIODo7XlQxV1
hsUy8Y+MaUj4tBYqEZIzsApGHGpiuMJFDA7c68imFQ6ZpuaatJdiSQgEYUWIE7pbf2sbQDGNFYOL
UyARqQkAOux3ToqD07B+MBOEH48bgW+2yf9WUxbz0bRGMe+0bCqya30tXiy8+aGfENvR5KUciWDp
KpwUTml6oa3b8Y5F84v4nOIGkBkwH1oVhl67tTMNo3vipbkS/ykPRqZlAwJvwBNYnNC5UyNWZuv1
TeZKL2xs8o31BrHtAbuuc3f9PvtduYx/zah3OHJGFQSws2P6Q0Gu40shTYIC/90X84EHXhBjK4iH
quV9ZN4A4SY94/5DYhObD/SCcwx8V590fYgkVAey765qJYAelwYPAdR9Ox7b98P8nXC15vwv/fZB
jBji1JY+K3AgM/cWoPEydevdNiJVPE9uHkUXhSMIA7nG/PrVmAX7YBoroF15TCL9RGAR+g0X488K
k80j+l82Kc3pO4n5KQ+vuqwI20aP/lFIQZb9jqOxP/siOJC4pcy6yrdwahYv4Q0eyRhwx5AHBrDo
5T2Xvc4HBPmAnSXTHGqVgtU+mEyzWjAmhzY4D9ZjwMsO2d+vEO0Ip8VecPK8MBGtILGB4dHAx+Fd
e4VkCIDOo7YtkS6bCGsnewuCEJ42Fl+jDf7o6GrnRR1oqWY+MPIfTFeXcecqnfslV9queqDkVd2A
l0iggQ/RxNfEhb6xnBSxDNv6ZstghGd/4IQGKtuughJrls3TZdEmC1fQRQOrFneHfNgX9FB36nq5
YQgbJywmDxsJE8VhNR4avepObON5NPUV6y43Ue0NBQIu3YlZFQti1IPARyuu4erXbdGlYQ5suRaX
h3Eou9oNsrbrOHPazOu8KxpyUKsoefKokkuguH12VI224fyIKm4thwgy0itsjb8/Txgfv+RpA4ke
ZMEOZTe13tm57OZ9cWboWn9QXMlQdcQBhhNjSG7LH4S4Yrq729zOFQHacxI4XmHhWPMb7m+JjC2y
kvuMsxs4w7eLXgVKsdzD4lZHAtAdjVTOE3qL2u5+AqxJ9Z0e8Zpv++U7+WV4OcdmPxerslNSDvYD
ZspWcBwZbTAE/XZmnG0LfwS6n1vwBqWaMTroz64JFzmAzIyLBU0Fxius5NbrhSfpW3m5p8M0UtA0
E9lcUhAc8BFiYg8NnWUXsdR1HE7itqrxb9ObVstG/QBFNvUKZPoXY6oOqk1N/fMKZCocczyRNie1
iE2qIiqHw6mVbBdIjC8TJJ+DGqy6GphtveIbbJK/sooEPBxh6sc3K4hnDpdwJ0LU8yrNa273rxWP
UMYnrvRD5KN523VfjGVLb6DkHA32Sej1aJiqwVZKabsHEar5/Du4JYcWI5aVnktuqB9d/BjmEZa/
iyM0KcdQK/UW9bi0vZPoKspl7MmMXNG4fUiLpVlt67wPMiL1e6igyX+0QAqQ37BH9yBJ7EcbiBL3
Jy3Gujv9L/FPeBxxiogVCO3pimJ4cwBUso5zyvu8gjJQe3CkKDtaDr7s02CQn3liDqNItAA+wNDr
jmInClv10ft7Xyay94xwHsHwsY8hsDezDqfahiXv8HU/l6ierATa2cTonjxEjGURGqsj5Z+9u/8n
xv57iGLCnIJZPlgDxHc1GiA6RsrPrEw6karT8C3u9PsV9XtHrnjRC65WEUh4KLYrRPWNCnw/vtmv
FJRWx79kFauAJHPLBj2oHpfMDyfUMvI4I+jiukB9gKfIdFi+cozQM/BVJ7fqDQ3DTdenG5e9qEVB
LlhO4XsrTQOraol9Z8GyncQ6mSUcd0DUefu4IADdHhW4WYnjp245+KqqrrojciHWNGQ4l0MU6gB3
2iEZICETqKptqXAMihPZnAW7ALYM+Hn0RilV3TucIeur2M3JNhPKNtZ2GMg23rjHls0NcHRxxoQl
CDmUfW1qYXpr1bk3MMF2yBl0rQIoF0sX5NwFLVmc0vffggDHcO+DW3k8IFBR49IaLjKC96Ui5lUQ
FKchbxkN9/66A8dwZQGuNRogRbozz2+QPoPIA3gcjeCm4KiDJPX5f8wq1GFwupLNhyzqy7dk8sWM
5w20rrlznY5T/5dupY76VN7oQhlICuXb2VqcMWJ7Sg0XbOqTTvhmydYNA65S82jvn6V4e3rN2AyP
938y/wASVB0KYjyRJd/V8U52BxOT6LuxE0kgKpaY7f7s/I72vkCWZCq+xFzdJiPLZmgHwd/He2y/
hTh6ACuVH0fcmd9Bh5xFCvSFO1iyqdvAy24H8irnc+C9WoEg2epp0hc3lsULUeuJtxzHfxC93vpZ
oapNiLh7NB1PFrtZd9LrUd+ITA4zNAi55GwcowmikCDBnmiS012nDr4UeEAhgpn+huWSlcTNe/68
LKxyQrjH4Xwguol13oBdIv2iSOHG1y6hZJ7/FIv2yHKlplnkTY1WSqw3fNhgAHWfOjONFInY+vS5
+mY++MCuf1hQ5R8yI1zBw/zv2Iq+Mh6dmVsDYCrf+juDYdNyfzHQaBk7DqoLRy8hsSvV3YdUe6NP
V23ZP+EvKk64cu/j1XhDV1cmdjxrJQbaMiZmVvVLSrZhvFljdBIkRrHuGC6do797wNTgZdKXeTAF
1Gr5w3ONvm3bU2LXTD8MDPULtCLavaofpI4REeaf3rvxKnNNQRN58/rirkTLIj8z/gQeDdXu7+xv
msrY+EESmS2yzd5BVtN9yruh8G5xXEu6JM0YpCDUY0sf9fqundEaOlNmVU5MsuXzUnu+SzUa19Td
S4jx0wFZIxq6lJr5svok+RpdzvdeayW4AQgE93Xx4+gc0IDIkhfzc6PDas65eCM+1kh0cbY18TTo
8MYnzJ3XsUsl+4J6CyfyeH3Vyc4J7Ucw6G5tbgm/++TI/rgBOHqdUDxJNpbT2IpVjXP1OpADhqXJ
X3sgiE/fzb2SKyzmI/F3UXPEN+vulmSPGSO8w9IbbhRCwXEmO2xrwZ9BwwPL9xXIBMuH6LPlc52E
EW3j55yhRceRB4TvBidhb5WUoxMZyX4OtDKBPeeiHS4L47QuMr3S0BDSAThknTkA8P8/HweqNRHR
o3EQk52OE2inGno0wJyadREN3s3jL49yQkd8ptGgsF83pmnks1lvToG4rklLP69W1EnMYuAPmYhb
R9DEJiicF+F9pgOQcC8j7faC3eLvIBPRtcbevMtuqvPaapTRWsOVGkXB8fdTAcsHWDOMALLY5IPA
p/dh+7WCFsAJePUUuwuke9HFjcMnrCNkxaN4qXmhBPxbbvTZS1VtsFDRgCK1QSMfD9tGAeWxzim8
kysA/f48lreDniRF11+5pXF44bTac63D53V6sjJMkTxYTOL/K/eoZtaFtd70iwUvZJh+d0KcBDTc
MAroO1XBLqzGwnUrHks8UJipWBw8GOkPE1Xus2gmTklKoAQ0mb5eVHdD8RSNhhuZty83WsAN1KwZ
hgBjcKmUre18dMW5sgL3MUuSIc3m5kupvLKDcJYNkKmMhUjb7EfsHeZMB0qJCR+TkBO5dulYfow1
GKvAF44J9lHKwaxEp4q0nZXCdiXgunNttr+vLPxv8M95SH9pGwwqKutjkvWv19EEPnl+OyMUKVS/
uSs4FHPoec4pm8MkScV+mDwLu1FLW3ADQYnDxRBvgacysj6QeiUcYmpPNKIEqOwjJRleNAl/YhY/
u0eOHzk22Oqs/XRKqdRbYUTvTs1NwzqRSI0UydIUHsiH1Rt06VwI5OMPx2elo2lGVRDsnZfdVEE0
1clxnAOFpiLgBPP71huS295uMBtj8TAtFzzOIIhfWzMttRc9GpjvJjVEkpXOzPYkhu/M6lFeoZUk
ElwjKqHm7opz0FXLkUARMiJNHfaAlqx5ZaXAWHb40efmxAg7rP8meIXpT0676Q2RKtkQtzB0PI1j
kgDjtWaHWl5qPvL1NYTT4+IBdi0J1ia6Ov/oMVlfaDFjCxThhRRJup5vF9YetbB5YCj+FPnRcels
6i3gNS2vuguI4RxP22jv6tmFcOjZz5shMakKMw/81NANO6Lj0PfDBR8xXYa9/U4gf87JJfIdzZDu
y1zjtQPaEHIQIlN/17pvK/gEm7RS408kUeEnsAEVN4ySiybJ4ENH67ihH3BUW6XtVZOQm+w2Gdiw
2oSUgQoYYULXEc3OG0nrdXHFxbDNjZRo1AneH0Jqoeb0/tZbuKqvQmmfKK1f68TbE06Oi235n24P
C7uNh0VMO9JdPiwCOELFrIs5ShMGyrLZCQt4Zz7OrH3zRbSCXzWpGWdnwxKKrqy/xG+JnKiSoV5e
ZXh7Z9lB+aKCn8dYCc5ec/7cdGT/c+fyWmPFv2E/IP7L9V0wjlwJcIHqbNtLQBviSffA+IxLtpmw
THqOK5FRRADXySU9A1Wx6xOwONS3oNZOIk/Kwp/docJouW7b7O9rOcUC7Vrb+eX6bRnckSkg9npA
32D91dNHG0RQ1PBfAXqlF+m9lLc+c75NmLx1JWsLN2ksjmx86Nf9HxZC0bw9Zq+nuKpjKjhFSWuK
nkGgqsA62nb49wH7X6AeyEwNYpmn2E8WmH/EtXaoAamAo4ZssMjEvsZ1Tyqc0iJ0jxUfuy54KzPE
4T/p5L0be1mVHZYPMUyAt6TR03qKGuja+SBVt23dAAPNQdFljS6CDNhfLHqF8d/BtE7QeBRfc4NC
dlhJLQpzk4hx3ygHcXL7e/AR2XmsTsFnYgK2tccrhENGw6cQfmjDUHsH2FKX/RX7jO7GUd424LKr
UpMihiigPF2dzJ6pGRU2EZWJheF76hbuAmTIQDwdM587amotGayHuX0GjgEbc/rY4Wy42PZnkRCq
mw1trhf+I1X4ICyNwyO3I7lW9a1t7uzHDjgjN4N/5JDoUJu818wZKevpWmeKxUdS07S/mDQdH93d
SOlFZY5H3PqrG9CvRkbX6bhna16VqiO9zLS6gjmiBLqtO9Uz4BlcHHWAPFko4ytuwYFYGFT3mXFs
Jsm1ydyDNAanvTwWqDDjyFZ2/95IoCf7JoRSTFNdkLCOJrAm//QTNF5L5nJffPF026+XlOMTHmzT
Uoc3m7I46swxHFgLNzOXcQQ49kQm9uJ0zpwx3mW/LTxuIYkuOuFAjRuAKcVTKpN4dNvaX3ay1alT
LwruQyJe4zifp/AZElJGBbjfliCoZBVJ1XroqVvdV0iew2TN54OU7D7JOyKyTROroDXYfmVbwtsF
H49g7aingG3pHjruxsUADITOW759O1/IrdblVOjNo3o1CCjldbhGEeGzVume6Cvvc+LYALWlK9SK
KjX2iSdnB5YeS5zfPVySwL+ub9x0IXai0PY1F/12sFfqD9qIigU0t/gbt1IwZqkxr8DS+630NWWR
QOTGhryqNBzC9Qi6z4X5B6KAJMHlffmNvNQdW4jiziLY0s2LH1KV5wSb2vte2xugxmNwU7NNLcmg
GN7pk4VvFztd0t/vO7c81geSRv3R4oM91GzscM7RrvGyAbhkqdYj/+evATlX6pu9+64Xz9HlyDPw
eeFoRGAt/KTBV+HpE6pSpqEA2Rb73g1O+CV4Ql6OQ0wum2IygLYRAkpzWVtGQzrMvXDABw/Wgug8
ve+seRlSmWSG2hfHYiyWly9rY6c3F6bsG/2Q/2FbZwsv5V7LPSAzw32L3cKdJhceRcGTC15EsZ+t
HYLVoYXlywIHt565oFE/21YnUnwdWmiHXF1yUUI71KIL87W34XEi0bFXH9K6QEQg0bo0d5NP3TXD
Y3p8sRxl7NMOPWUBU0vEPQ4i6bRu/zF96PeaqViPgdsREpU2N6OiLqZ+7nTYNaRx860grdslRSHz
8S2zd8epvgUFGXNWF7ppB52/afyNAVqpV3K/2/EkeTJiafhu9cT4O6A2fgkXtb1FQC3p52jbC93G
Qxd5Gzl3g/4/KXIEubWyvvoBvYGz4tBSiKUUX1hWdHkW3ccLPAXBgtFVj0TVwa6xGxt4tFT0DEFz
s5fe3ZS3uAG6kBhX1bpdnJ0JEyohmC5+qD2fgWtiyQFuVqxxY3wkX825OFrmCKPruYbmCZDGFXZp
SKLb99y37Fc5QK0tVy/pJAsaj5qHvFsNJYMsIr2WG3lW4DyQnLLCgesxE2iPVs0qUYZIJ7XuXRl9
Ots/irWw7g/ryoLr7cn9el/pD3PeUQEd5bVOuUgr9hvLxLqtxiTHvidicj2dm0rieIJhW0DHErsm
YpQybRLM2l98yPAProLniLhzLGNKHi6Rddk3oXPTm5MN+gHmnUpcy1aW626fub1yiyVxcF65bsq+
9coQbT/AA8n907oUkj1r+7DGDDpGxP/XEbT1fAKXV9tInfG4qk+cgh4ShjirO0zlmYd8lblSRMGF
yKI01JwXKnvauYo8aAmKns0X9h+CUBBzjTBXhvCfonyB7JVihi4jzdqz1f9mU31X1vWDP0yXKHH0
dEputerlQqrBOWE8vPKjJVPi2p3om3QN9M4tLKNqrhRF5C7vP2JRJWrXOop9+L4DpqCuvaYopO/f
TI6QFLP8O7iGARGgfPpaQ2OzR76TfzJIf/U4FELfLGbRdjYi/BK9/XnU8JjUr78Gg+xtF80OMwBE
xaXrCgJcLHlNXbJaa8lC+nekWfblbRTUcbobsiJ+l67jHLNRZTRQB9bpqr6bE+8QlLmeBoghEWag
m4Whl0lq37HPLLy/Jgz0ArhKPqmSfHtyVNtQuVXLw3bQqCofLSwMH4Esgoixlpeba06DE8yaAmKu
vfSg/XoeLGUO0+wOpjetnwtwpUCLPZVB1qw7mcSAr0dwl4yYWKxFpwS7Kbm1fNsDuyG5MojCoMow
d1AEnAWmHIiTMC4ugnjdeMKF/oWo0EECbog11g28W07ALX8xM3DPexZmzwnIDWzYKk+kqoSV897n
NS/RBynuQqQ5YR9JF4J31cbcd6EKWphE+8KeHqBDLld6WfcqwJe7+3YMqtjamQXfd/sM9lmfgo/j
jfvezN7pgICZ0RMb2ge/t8NAiir/vkCq0JtCnT9bMQSudBrMNaInkv8HQEhxDRI3Ur/58vw9uoBc
pJoUpqhZN1gp1XnuuvjIAxrsuNR84h3hVQVyHattyme5r2711mfIKdOjP2oYlFPTcasGNatBsuYI
Q1OG4IeokhsuJnu7Btoz9jWvC1NCfw9oFaA2N71q74bAj8EmtrLNZ7iGTvLWXHX3ZtX4R763fXMW
kbER6IKNvS9zHaeAuPvCLEGv9d3T3IRyP+77VIAqjmIw+CUXz1Bg2oDD/3sh8dpTZnxHN6uDbEe9
a/ax3dOmVcJMaLFq+k5+qMABwQjF9QVqpcn4mZGKtKHOyeoSjB7MWpTykG8kxOzn+taE/Z6d16VY
wci51nIfVkFwj9o5fIWHaCw8eRM6ouj+UX3zbNX5w5HIztbuNzuho64+vCZLPzEXRyCCc2ep1bsw
8FC2YF2B2Rp44Ba/PGrmOqCKRC2ZzzULNiXkDoFJziyLHDerAN4Guu6qKQkjbW9Bd5Tg/5a4LSUm
ERAj2sRWCCdV61CV2dKk0VAWm1iM0x57FYCzIDTd/GCTivMYoSKLaGnOTuwlq4AwlBjCD6cop+ci
d8LvYznoTZ2HtId6uym7ilMOzKfJE57ReFTx/8L3ALG6ShZayFn8LIgePlZKNQynxI/clyHiyrdb
hGjoSkVL1vFUHvFb4Cyc0eaKg9aHXuyYhR9bPkEDrrlGTF9haYn6tFDbl1SXMulg78J/vroh/41H
HrYAAjQDTCOjiJhxRRj+OusqYrik+KN/Yvcbq0bpv3oEpkisZ9ePV2HEGKrUwKrPDuU0KYFhqOZa
dMqZWK1pRmq1FmelZQC64V/CD7MtlkT7ZzWP1ewKBnUpimuTmUwz4gU801iarxjZyoBbdYaYETSw
4ugbpO+xUIyQOhdigzhSVr2lziXnXdfqIn6kG6jBTJITx4T9LD73XVItYESY2WXOW1fkXO47Hfp7
FK28rQeUtJ0PDKOXnOCRWgpfKUdnFVTPH2oMR9rNzNQxwRd/QqdqJAMY3Z3PJbmiTP7wrFwrgutz
a9AKLxT/nXNlsrnQ3AafANa/91bwOazdJ2Li2yM2RpDbbtT9/5ecJey5u9lJ1xKw5TH0rhQyEeSd
D2FawOhIJ+Gm41fmiAsM+40gAZnOSw9SXmKfDL2UjIAd+6M+s91CQx/EFfvMfLdmQZTrm8O5na05
SAQUDAPUELMNr8/xGJFHlddJZP62esXfHFk+eDkOKfIO+NUqhXPhTsgKU/humuhRw6WRMue3qEIP
QOJQRabEIFvBfMxUX1FESsPNTSjvMpIX6irurEWP/AXFfHbE9K0pm3SW9vUSAdtrx7AMKD+rmQof
9tmhcxVEPPn0LZCXM8/pwQz9wk1ERuSh2INxwoW5A+17ucharukdPwbTRBBqhNSoaHrzYIGWbkQl
SfVq9stSGBNJlk6s7F7Lgrvvqv3huZLvedpCb5tF8ChPaIUQP0bM2/WLOWTB/v2SXpNZCe/x4AEq
zFlKtXQYQ8G8wiSn52joOcEsd5t+/QIttMLzGvIRR4sA+C2AbxTJRazckWQVqcM4vARNar6WNQHi
Nl47rUTSglLAK13BZn9/4NxY4TqKpvGb31bSOrnpjtKzRGVFkJvAa2S32zuOWOG1Bo0dBX7ER32p
ybMZQ18qNrS6lcEq7tKySHrLaVkzPMBGqjlQVAC3UpF/z9YUQMvPuxWjcDyxXKO8zsSp5oQpLgg8
vOvLwz8U5o/Y7bZI5BwVqd9LfEqrmBjFAj0Tf2uKrBsFbhd89/pO0LFwJjvi7jmrHd6jM+wFYl8v
8wkbAA5oQrrUMPnxoKPTFH292HLX3WA0Uzdun6cjuB0LYPDypEXfiyXQLFuOobw3i5oM/afaQL7t
fJN9rIZbLWyzAXmorXcvlgQNtF7lOkf8Du2mGUGs6/sw0Jf00UZEDv7HSquknSzvQadgTyvXDCrt
tnQLU8QpCZP1D0cRiMU/k9ufCi7Dg2VnbjiDLN/82Vjml8qXVrPcdjotg1PnvkP0tJThrK9TWWHa
7LimdzOSFfXCLrC4TtERQCdZkKEFZCQbQuHqunyTwrZHEA1RJq7tkrWww1LkwkaI1B1U99FhiH5J
nL89kRa26ZcXWHmUWl4rhW9pPGTSKKSntowgGa1t680MYT8RKJeF9xJfWcFHgx5NFjVA8LK7Xalq
zOWGK8r8zuf581ptBLBgLKCo+/xwAprXJ7bNRDuf+U+bszpkdROhUsKbaZgVKXsBSCjfkVdT5LF6
B298ZfduBfZ9IKKozCgcIXAuPIBWIRaHmkYjqBmcp/UYEx+Z1bke+PTb93VJdhCk7Da5YFbDFL64
3haUotLyMKjsFI1TCIMjjD1tihpeAXGoFz3hL+j5GdMOjNDgcS7Dsf2BtHj3v43KgkyMuGe+DYLf
TNoK3Z5bqOIvp4aWmOnmTnw/cnKfefz8e4H5zVy6S/er5YRw7zIIYaDWNb2lboJ+rnzQAhOi6NUA
jyUDT5sNtlKoLiJMAH4z0nsv13wPJTlJ5khHs74h2HPXHZrHJ0ZuNyQfSRKSheotpvgRAPHLkecC
VIFX93+MlH64dLWwTmbxp8gc+Gm2E95Gvw4soMjWAbmsCDL2UdiH5nvlSZLKV+ofXkeSgSdlDMh1
GbXHykRxTelbcgL+S8Idpx2M6RcNiA6db2/jp3/b51BGsxx6bBG2scIBS16ej6IyFBDhQNSzc/2i
BZEZRErqISJAulo+ONL9eEqQdncENoFVi/C8gXtQxqB2ASBCiBAbCsdiZjCvYFfnmsKHrYxWQcfg
vQwfKVuRLkBvaV/d+6OZ66hO3ap5Ibrq2Q7rnMHVLXoLh90hA2BSiQWYD7ni/ulWhQUntMXA1/mW
/TrscP38v9lnq1etWAq7XM0bTsyvSrRH7eLMX7IOqeQjPhCTgcp24d7pbeY2Z+8RyGCsLcmkkFBN
3Gi53dt5vLi/Jt2lOx3SMWZ/FwAlBUJikPsyomEmMXl5rTlW4KBLZIeewiWGRVec6OD97mLzspVh
KWERcs4WZDGD5CjbdY6U5r0dspgKWvPvNSlML9tuhYwFd63ZWbqguseOCkWAMzC7JwAaSzCNRG1V
b/0kxNb2b7Ymg59KX26F26EoCChhJ8fr1g3HJcLQuqvUCjW3fsZY7txShKMWL2KZztj3qlSdyUXc
lq8mZhnSWkpEdh1Nkg+HkpHxP1AKcOVIITYt6t+EWprN6KplaJhJNru18us0lf74JahNSJfmTySA
pb2LLWViz1IkQbIg5JKMlNNYvttXgY/3pvsSqWtZSJ+VelrSWKaiWhOCM/m8y3Scu48769QDhOZZ
ytheseNY9BTF/mZTFYVHFInEuj9fdJ3l5keiSyQvE2x1CeZ7CvonK73hslzUrvAG2vzkZUxLVOBD
ocI5vnJY7t59qsYXz8VB+dwgY6d1sAUmVVQrKYU2VVKGors051dUR33EA6PAaYtuKbPXOm3tfXMm
HHmsj8mVa8DOKyuFnZh1Pe1MyberRd8KVEvyMv67Mpi4wopRO4RiuhfXbIt9PgO/MN/ZybY9KVhw
+KXYtQF06A7cl2omIkXR/gam01bD1ecPq/eyWcJ0G1yG1+z0P/PK4TX8rtAplWrtxKsgVJwRBsLa
NE1O0KM/9TbcaJ8WHjbS14BKmlMp8g38RYXsCth/sZ1OOXN02r7zkSSjk55o34U2e1+K2OtxUzcr
i/elkREZT3Vo4rxSvnJGUWCBZ7KWb8n7drUxyfRIsjeEZMnOD2uECuat+DUBbfx2zzhglWfnLi9I
//Xvrv1/Qk3+0NTv4+y08aUxLNcKSGid7dDIsohPRUvXaV8v6apCgqto8TeKud9ZxBnLXeLhuSfc
TsUj7mfsnGc02ggjx5G5Shi50lb48XsCTuzB8WD/dSMX5HLx2g+Gdy2B6tFQ06iccuvIRQzog7mW
DFpsUD5vOAbbjI7xsreC8JdpPor1D75aTkyarjxhi/at5zCUiN49IPe/eD1peOn+x9jOgBDLF0pq
UAVTpc3to1ilf1DSAvOiqjRqTvFb/fY+m9Z6dh+XKg4XD0/AAviWozcXyex0FDp8oyogX25BbZR7
HDBXJIpuArhOYrTvlICzTgn551oOL3fckRy1twDOvN2sgUV06UTBev66HOUnIdaqX5bXSYX2qrfC
9sRqS3+tTVjkXTIhJL5ezxGIUTUdkcVwNYctouhoTI7bo290b6JaEn4+6FlZoS4Rj92J1ogpT7mE
LP6ICSuOYm94BpHr3UUfRiO5It0iyQ+7xy0O+Zth1jPKxykHvhlghPPjNe0CDeauV1Z4bd+tkzOK
72a0hLnh82rv/BY/DoLr+dWvocqHZ/Yxi5BPqb31NshTFXaz5575Q6zH6Rro3g98ujgQ6NZxELjn
5ejSehddzbO9ot3OL41Gkr+r6GLFVVBUBFWth640jyWBhZmRzKoybUy9WAY5ADsvt51BAJctA1gt
XMurKwyb8Q/iLIcxAisBjpR2J+yGVniUkUfSzm7KXZFskvsF5MokaHPNaos1wk1Im3sfDJaPXLZe
VLEPXfjHZyUBBiq6Dq2PtCSaHCSkUsKXd3actONVajUvK6623hwRgrEu5lYjwS9I9I33IzpXa6VL
m7L4YyDOYAKbTK54fMUXZQGmLQG9gUlUhNQVtz0AODkrJwM729ttsWNI4xgmlLVhBSAKgavayFli
xR3KD9nDtjZpsKnYvsu/BrkhVnBYQBX+TBux34U2X4GLUikNnngMzFskw3RZjJ/SeYGUJvz1fDrq
Q+0bBbUAGYwuAB8KzGsmNa8Xrv5tc/jyAbO7T5P1OF8zOCUlCy5GOUF8YyvOYfdaYWgRMTPbA4Nt
XJOaQxjd/oK1OIXfUXkIrmIXDtiLwd2rzG9omVdFevu8hGriivZd6XttukLxv3HcyvorcFzkdhpJ
6qublggWMBpN7xixdij4oRhHzmTYDfrnU+k97EuTG7NZA27fQMt+8b9tzZ72eAr71gBxpGUSM7Mc
VndVcyM18t3unSKJYbjBOLCAdV32/5rL9j8bDXTrQR/f3fuER8ViO8+mLJo7TSGz260TQ95gbWGj
b1fn2xZ/QmBJ25ER+YQ4lchBpnknW6J1HT5NhRNVmjerH26r6sldIVrqQaB5xeJ4oTDMDuZ53b+z
FbTrnK+wXVq/ekpNZGIGMbcqDiW2WjLG27WBFLK2xz/0Gnzwupiy7RuDNGXZxK0IqqjDwjmvIGTG
kZ9I/oLQvdXDjthZVuWH72C9rFoHIAHWADMJEQpfwoIQV2uakV1b/YINysCAoHPT4aYG3MBoWwHP
49TCT8gQjgQt5+524sfZQ5bfA7p6eyGc2VtAItDsQuEnkqWHg6oW6HjVqauD7AXyEzvg7j5BC2uF
27mo/ZYm2SjtIQbVJOuWe2A6zX2qnhZZTHVUlq5vxYse5MRObbWpbtWPg7yQNjOK3Ffr6i/qEgqd
1q0gL2se1TfDE0m2Gi7eh+iPS0XqRg5/oUQVl+gVOyJ02Hku6qRoRA/rUOuELMBPJag147bNT5Dw
Z6j6niOPAPKrJvyRopOBqLSyWAdNU1zMx6ifxOkxxxLTipV1fkFezPnMfkKmfj2CFLlVmjE2u9cS
7uyhnSGVtQDZ234vg1VgQ33+IKwNBYIQ93V8eokJt6uwZ+1j5I8F1ROkEcRtfb+Zuvy3Bfe0wnbM
Op1UAnXVpozu6GvOClF5tT+qOwSa3GvbAcJICYJ9CfKtqyZQFdtUqxvNJAyrGA2Km4jGgLbJjhRj
wbY+PnIRgzo5bS1mpVwoNu2L+MtVoxSmrCw3NVvORZHRx/fGWI/vywPCYiT4BFCJMBdklqRx+O5K
6irkLfcCnkwYVAO/ofKxXaJfkN2Tbdcv0vhLP/zYHanxfxQImh4eWA1TQsdt8qBe/38AOb7TnCDy
B6WOM37y4aJEuHdIVUP9jVxgagQGg5XMaqxmkl4qLTDyDTvNKtZ6yrsO4u4KkGFKsSIJMEEHhpnG
PKrdjPrSNPUKx6W2LlPXcIWHyv6MDln6Z/Oq/+WMLVDHusTyWhw+LFoN7y+3xZRXasd/5DZgWt46
hNvBuZ7lae+sWULVrKmpSNsz0SwVQbHYEDun+b4rdqpiZlEXeQJ2aiA11uatZRRS3e42iIxpIs8W
DjfF4CjN3wzI8bTPp1vByrbmWTEnEDV0vyAn0ynzra/KSdpRl6/2RO1OkVwm+28q67Qhx58V6v1n
XfCjK2Bou4s5dQmFysrRiQ5+Ym8zuu9H3r+1y6aoKWCR2m9IgpeonVE+LarBQ57TOT1do4bP0Rfm
FlmBy3h0c11t625+AwoAO2l2i8kby/ezHoVAK3aLfP45n3+ifC8Fx4O+LzRDn9rxB+Pu/CBlFLdY
I2/nbk60qwwAXFUveErJ+JhmssWd4bABS9qKG1KlXfcvjZfYdugwiLTdl7GyDEFjhIrafsCQcIBH
O7PdXIahmCGdne87gdT6Lz/9upyDonLPDF4hwj72G9oLH5YXJE9BOi4z/4tQBwBJ80HH373AQ6MZ
p9Kug55VDd1VmjwsKWq7a9rUpHSWsw9+NpmtqWYpnJOQW7z7394pOyggT+NL4psCzBP50tpc47L1
swABPHk598qdcgYLNIVzFT911U0MrjGnP9awtzfu3iw7KgX1cOEl4cvTGhAjgqxpAjJgOM064tVX
PezVD46+ThhB1VfLrLFgqC0Ntg7HPmkFsfQ17emuF7adASwUq1Iqx08B4FuyXzbEQoJkKwX1c7wC
u+/irwSHokcBkRDYrVDQn5HSgMYO7cE8yqTJtaeaU5cNUePoZaeM35NOIMUBDYV3vOktyWD5ZIus
m6DEj2GXema3gKFgwpd9KqDCI1uqJWQAMgAWi8jylZcHZ5OF5SowSR0eX7Pwam/tBsUvkdzbvWHV
wIsnPTsJZ1J0A/lcKTU0hcMUroAV6wJhk0/pHmiHCg0lWQxqORlwPA+guQonnlaIiEVDVcMPl4mb
MkMbbqg2kRTqFUB5P9Ziq8gKEoD9tvCYWxhOvclT1KQvUHnJyoMTOCrt0hQdOAyNU7Mn2lFjnEOX
pkSk23ls9PtLV3ENDn02HrAQNO7FodmtLxspPg4i/VYVH0Om6XIVKhbqWzUrC3ixQkr7+pqV4Df+
s7TDSOdYg24yOGLjydiKZ7/MgLV1vR3DKXOBQVzBLbIh8C22IDQI7C+pkbyWbZRoG5HAB0vXq3ZY
zpo/4p82Z9CofZitAdRpbBGeHRfcKyFlNwfatuK5Lbmo0Sgt5i3gW1tFUseQLB3yrjhrKamMoHLX
Cf5ogh1XDQHl2w6t7wUFiPQ+bnyT/ZAFIRR8FYAnljDapR6hna7BFzlYHDQbYGCni5UTeTGCQywa
37F8pcEpm6nS+6hB4iiP+7wr5BNo3abtIbdKXA43Z5PRIRKpZOjnS1yvrp+/3brzoV+56IsglmRj
0xOu+HC9Qluak9m3dpPEA0ptHpIyg9kLRlhDqjLXiVAr3Eax3Dh82aC33rJ0TdWTKw0xknvwYE8R
t21lxkMX8w1M19UdTdT0d6gNsUzC/zbRNR5UoM0s6acY3rhJuRp4huKF4h/pFx3kegHEOmAG2TvL
07Y3GBfa1q3dCjbcUrh3k7rSxze8/r6sdKXC4xxuC0DK+laC5MrHwhnMQ97sZZwUDm7NggUeYU0q
mxFhrE5VYIA2ixj4GXkE+LqC7p7/7mGNTSa5OVfXA3VtIHLNPOmEnDiYjn7aSAmJuuLa7F4gtJ7J
xFcS+l6QbglOZBr7CohuEhuYMLa0iKCiUQs0YcrJdsxAlXFUVeHNYVLmSR+EkobGHKZ8tDhGNfgH
BA72t6hPi6iIEqtQC2JH34TVn+9P3M6uMml8rA2qjp4h0d6rVbPtMmBlwvWEmOAHm8hfluqQD+KI
rjJQk5bjskYB0fnh+XuiLqGCjEm9DnWTZbWecFRHNL3JK1nZcHEEQqeUzi2Qycvpr73FRurXt8AH
f2f+/DvhBroeleFpAH69OTkPd07JUfz7pRpcBfeUhobr24+my71Tf8+0r+eeeJ6EoPr3kMBUBWE2
s5uDUFiGwXISJ43+p4NIHoQpiyGlm+0sugeFzTjTIkhLguNp3d0xqIPHdVUJhOO4w8gFZH+iXfAw
vaewv+zXaoUffc+gUfauWzVHgkpS28uxB8W2KN0iL4Xn4KUc9uSirgfhKiqgWXNDj6ZIfcvEnCDg
tHG/BxZkZInZ0aLD1LC4fRX19ggU1BLPj9fuW0+NF98bhe1E75Nj5C4oZcB5eD7rE3BdIpGlpKea
QzcBYYmJKEq7qojeuQSuFiMpKNSmkTCTRzGbI/2avEoq7zXa9JWMqRRoBHBXEvPSklqvvf9124AQ
i/7NOdo9knCI+WU77RftTaz8ZvZ4q/JkU6BPoEgd/iJYNGHm+dM/BVok264VsQRRspi+8RfwVps5
k4nEQXnf8w1JHVX7eVVNowLtb5YE3QFrMqmQeJRUYOfQFeAyp60jX2BZjesb4hofCQ2PhPRY6X7o
nJJcrEcsVe0cyJvRG9ERDpF4Icp4LvBGsTqaNfQe/ZLPB1e1JYbDemm0rYUb9mfrFv7nspBzk54X
e7mGMrkCUVGmgfRlWG8wBULwM67NbOL6MTVouHOAhz98+m3cON3G+97iiE2Xkx6MC8bnVtI/kiuz
cePN3ngRFXj51e+poImfF8Gr0KxgUgYpYV6LW6jtvCCEyDOVpP0fcPtj89Q3YTbPoc+Hpw/2rf+c
RG82NFT0sCYV01o61tXANzqk3L2PDu9ZbTB+FlXDeoTxETqwD7fNW267swV8eqky26C6t5Mmltmx
bK5vOsbrJLkHS5jNjl+HE4+p5pPGBPmgSDQAZsqwIOMvFs/uC8nq7zdbgfWGrXNlKX+pnPRfmjOO
+NgKsj6URjkB3W9GuoXphPgh2XRdFCIi6nYpHL4R+uzPQJFvaWJBJB+sWu7uiyTJERD8/t+OaZJo
Ie++XodyGkzHFqaSyP9mj0RDUXpCks1DB0Y3kYAOz0Oasp3z4ypWtYhAWr6tOiHj6fV+7f5IQG0J
6h/sagup9qvMKGplVPQljU4uMk9BVapew7Xq9NxS8fQLF1UpuH7/OF2ydUF9N05NCcYvgcx7OGia
DjzgIu22m7dvlgbVaDGgqKwOfEeqf/qy+6jwMCTaFDCwE/L2cgsjES/qWoQ5HDrd9Q6hto43HT16
Qix1xb1fMSred9BBwGJ3hIryKHP5YRhn4Y5r7kBGI0UR9ZKDobq+JVASa4ubYDKq/zF3uV10ZPCz
60R+tNWAiouDLPFq/j7/tswjO6aesK4BVziDx4jOgo/FqQ1dDIWUVxLszGxzJbZE70CKPInx24K1
2oW6IdH82KB1JWLe4xXYaMP/xdHugud9buG/k4H0mavfv7jJiF0ZjD7bP+7NUVDbxfLA+hVpq3hE
wEE43UECNZ9Y+xpLVgNDSOBnLhw5k74/GZHizOZ7JTFBRCBxFY4edYMYgbAikkt+KwX/jo0b+4ww
LFvoquQRacq3/QwNzFokeVv0mQnyWIOyNfbHPx7WNNMSxnggt4NdIt9tzD54Sn9XCci26pmiM5S2
BPBatdbGpCAweQ+uLdz1kei7+VQUwozp5MCk7wdJPIqa9/bBQr1qHsAMJpNfhu98gPrqfO7QfyCU
0UzOtDYhpLUC4nOKxf2eeMoN4EmbHxUK+RIDTc/6399LmHw0zeT1nLz4r34mBS6aACDAG/eDDJmd
BSJc35D95XuP/kacvTJWTsD//e52mmjDThOFajbnhwzSCBF/Yk1Sgq+n2ls4zXMIzl0zaDzJ2sM8
9ixe/3gQaCoGYJnbRXvIRBHz+VyKa2hWBhJkQSndz7K3sgQwD1W+oNMEFOulAN26SPl4F9x6mpGd
vfe+LH4BRmkdGgp2fQF4cbNM3QtzlX8ZXgHcbYJv4PmODVFa5jYgrCsNGfIciXTLDzrXK8bsyzEj
Vm3BgZh1isMlQ9O8vyKYMJWRmfWlA2th6FwQ8ZUgd3MobYBXhJIpzhTAGtoLF8JFV0+heudSyzey
mZ106rcJC4uCfwyb9/mJ5IVyxx81AmMx38LJ8dzx6bl7CIZsodI4NwxSGPCetii7JR1MFn4uAxcN
88tGQ/4V+ZrZD00i/6kdqx9q7PRwmOyx7BFOq4MGKZY2M1PdAgHsjgjNMsBePUSxID6yHgQxbt6q
lBDXSYQjgIJpUG/xR13KMgNpQ3dorVvhC26Ztf1gVzDxrOPJYweVOuOR8UsRBGOCKJVb7wJKQce1
N0TqteJkSfA4Kfd/4HSexJT3k6KT8H/xjRI+/oWFYeR6UghocHzhP3lststwrTzjuxv8jhXpp3GL
iEhTvvjLDB+13a60ZDQwur4T1Pxy1flgA1HaRYhOrQLoJn5WBZSEJNw48KxorJlERViXsWJxmzmH
kS/9sVwAXGfZXuBsUHNRqbf9nWNtEqbKms9eICENtXEo5Z3VljipkKi/yazYd4nlKfuGAT+Ppa9E
17U6yz03qDFDQIDexO9hA3y2sY7i3cq4t9344aSqZJ0D0ozYT+mZJ95w3t5gtmzNCIj2V8kl+YmW
K1Zz3wXyKnt0YZeX3XI9ta8Qg/ZrJvhuhVmb2vfUnUGRmXQObuEVZhdqFxu9H4KYK+NEGPv9EvMy
8kSfBeP5OUGXd6L/73Yd5ppwYqcqiD50hJ+fbFb+K30NbuLH+qBq6diCPXyO1XeZmo9XViuR9nRh
l14yPE61S9o5lIe497qwV+Gm76NKDRqOW+tJoC1GmHTfb11iTtsNidMvNW9TwXxOl3GszYBK1XHk
fIJek8KZFu8vLOOCqi5lmZICXLgYjI3MiW/UCCmP/EZIqtG/LhAM391nK0RsFKnh3heuzR4bw5+L
HZXgFNQu+CFqPG8JDX1QeMIuUFlPh42hH2NlW1W+Ok0YqA82wv85tqmAi38esUpMBfu0slRFn+Mu
FRik53J6ujF2sjKMeKa4cFGDVARvNCVj0y24jEy0t3B49lcFmNS1hdAd7Mvsjcox7y3oF9q/O5ed
xijjXjK7yP6+DS3pg3GgKFPSBSuEXIm/JITVG6Ykj62C4Vzb9AvPFEsAv7CzsygTU6tW7L3bZZV6
75mVhn9t0Ks808wXsUqs0WGf4FnljyZmodmcA9oQ+thcwRq87K7kGkqS+aEsUQ3kZXOud8WZ/8G0
MHDHkgw95GcW8HgA8/R4U077lSaU5rKmbsKpWcgVxxJbBFs5y6RMzOlXZHwe82lbPYCkIxaT5Esq
YC1FioHtVFP4V3d9NyFoFUxOuOpDuxi8sM73u1zof05PK3/alEWm80zHAVKABP0lH2NqDjsOl2qT
AoOdGXTTrJN8jRw8EEl1AgCuuD0Si3BWuP7LWL55345Se6kYjGqOA1PQUNRqaSj7k7cq6UUrlFej
/o48oj/81irpBvAFQ05iIaHKrNPc+/weM3114XnsD7h8CAssFjJuJomoy+GlGC+eezsjlnd/jYiQ
y69WgmVFmp2alumoepwhPmmn/EUQmPl97jw+4XXGbOSPIXwNN7orEk4Bh6OKKiAOZch2kCKZH8Qw
50bZfjvug/qCvhlMnWsM1Z7yt2UU/1ai7LnclgHSOjXOk70E0vkMD0uo8Hp2PDJCIdDtIlHvbMx8
FSftpgigST+C6NODxVi4MKHhpVQi6Udz4Zj/3TUwGlQcU+3OCZZZcrNjDZAY5gX3B/CD0310osKj
tMUDic9yogoOxgdmQNYA6fyopmkSS2sz6MDMS0RWU5iRyg/QgtAs+RiUbsZF1KjVlIzBZ28TxAJy
KUTFAboujXIYTT71oy2NM6j7U8ssMEatBt4a2aljgWerHKCbXt0gmAS/aVJ2FrVJh2f9MoBK82Kp
fCKBXpuXI/YdR4maU11PaMYrSKUuqdb4GOhGX5FUpsCeHgL9JnA3xsNe3rTuGplANm9Jpz+NOpTi
jcCdV2J/Q+Gl/vkSIaDajazrVBKQkd2Y9/7MIkYhPWdeCtBVehimGyO/DkhjIZ7SwYmruB1rIz6q
3jEOaIj9/vT3NTXquFJDc8SbHYedYAwtiOjP9o4EzhUYyyKSJYnYpCZDzl2cysDTbYKk0Xpe3/c1
pEqE+40SVaGccmIYE/dszOWI3hOEwWMnEvWAd2MGSMecwpeoQgnopzFS3KYMtcXUXkItTVM35uBC
b4ACAZ3VHyy02AqpUR57Nk0k0h3kO6kiLa1jWv53vEMyDqeNMQyDLK1vvT+NOdJJJQaPfRknbkfH
O/Jf0pDolwCkHqOobcP/ifTp92aSGlML/UHnFgG5mid0ppXvYpcBl4c8uXJOw2/8xIC8A+1BljoW
SfJLrxVuPzuu4mkWab1gPpXR7XyV9bowXAfJa30Ro8dOGXdp67dMfQe74HUTqq5ZTelPGFpxN4WQ
zr9WZK5zJfNoX+cR5sWaHT7eQNA0nDqj4I2Lg/AYPb7cgOqq7sS9kFyX+3sBn5oOEpyug+q59o9o
WV8k3A3doU0bKkZLT1dCO3JtmxHZil2fQiBar50gBNQQuPWY8KCGznL4MnJ8sH7utJn59MKr2Ay9
VL5ot1wzJj3+51KuDTReZ+e0Gtn8QBEEzwc44BdhHDWDnCphdrPd2ur9SvEPp0RS6SvZSbAEhSmE
8gVzn4AFDjGLK1lqBlvGCGhO5S2vQkUHfbcJnLdXXEd7c2Yi2uQ9HmiTRcPKu/aAtYzRnBDk3FOl
Ayavl02ntR8ZsIFVpHUvzK+CU+/8v/ebVGpfijR3w0QfNbIqdWi8zaJS7+Lc8Jn60T25dh/NHHJA
CU3ra9Eys8iWiU5BGJp2wKfiIEGnkGgk5YjFfdfqfNzvb/1wge1K9Z3+A0xjFtSAf8qJt56c1AsC
qUzbYS/mD81rzQwzOtJ7znUDfYSypKuy71WhkrBv6Etqrp7hrUs6OyfaKnIkBZQ6xzsRYJUx/ngG
AvFpRZb4StT9f6Knu1og8QZZh35+RpXiXHZl5V7pxZv+H2BrvA9aedUuSjDcSpR3GZGcGw1MOQ17
tSaz+2J7hBGdDXxIyqSJUOGTaY1zZRDcFjxvt7ajQurq2kdtPycoashhhzwpkRsMAHHQBZ0/Y5oy
YAL513l/2KeYQRrTN7PQe58S9NFTQzYddhBxIBQMPTQmYNHA0RZ8iKH57F3uxGcqjhONtjqt7Hdi
AgmoXKEEIQpSFOat330K5CkI/O8ZbNABrqn3mV0aZ+a5bamsJW9ocGeQ9Dpt9XcjmNGnN3TY8CSP
6OZdoi2KO5L1HE1KYM1kOvDf6cHW86gMg6L5p5GBtb17tnnlN38Lc5MOv3zlxMDmxVSvysMV3T/1
kTJkLMP8nRG94QUHFe+pGqUlCq+bO+pIvKcwP+2gr/w5Hzk6FDZ1FHiZoEEv9uVMR8Dm/eAuecJS
vsFmW8qh2yW/2VXOQ2ped6w2GIKjCM4iHTCuwIzqMWSy6w6Q3Wjw/uT30/2MkxGOAPYxawtys2t7
u1nXbS5ydoAimQyaF19oFY9ankdSM4XvNWMxA7GENm1zf+IYhlx8Xz13ozYd9lh5ciTEQiYbIh6L
OtTewj9AausNXqNPEOk5hlSTcttdwFV2J6WTtmg4Vr591d81J6xKuQ3IsbuKOR8pZfr6KcXMhppa
39KGwjoNb/k36B1Gv6A9P/abu0uJBPrRC/qoLgXfxrER/Qi40mwsHpEU4kGrzrsOhVcAq0yiiuo1
EIxzn+qgEQ/DtZvJsP7+Pxp7V8dRnhvliPPSOHXuuTX/LjFcmRuPEFcgXIobPUAXxlM/ig2dHq79
CJoR/flXa/+qAz/B8dZgYXr9fqijEWlI7N53JTW6xY1mIyhuEDx1/G7S74oiR81eVtfl82S3OIgl
4p+nqLKHc28OlCyNYm0vExPJZ7QNrEL1C6WXLCpYcZV8yNNu+HQld9Ti2wbONouI7GPtxNPne53E
4jAsPJePYSCJ+RV26v1A6KFQGWlff1jDFz6kWwZCsOBEOfzVouNsFkiqViVsrs83ueR88Ilp0LJD
2/n2rOdTI8bM2TT/SnqbYaB5tvzzM9p92AOOYAUszbUBTp/Tjq3WP4n9uOjbS7+iWIDvAJtLBG9u
FGci8JwOJGkDh3++9hUc7aeZrpEmPp8OlNrFsp7dNpqBiS1RGWN/7H/MK8VZT2eBi1PZiG/haocu
aSC9jTRn2ZJHmf/R8mI2n2Gr0qEhvkNKO2tYsqReDSsDWpXTj53OCbzpNiK9czlG92lmpN3DakhU
OOl55J7YhVc0ZA0z1kJu2FTAvZPeopuxCdlWEyg5BulTcgzcO8TdGonZL8/sdRqV6K4NpsOUzlkY
FSQUDNW4mIVjhVtlUPvFLnRVT6z0j+lUBIJQskuTwhj33Ps28vDNyYrEdWHCgmI3KpncHiZeGrgY
CSZinkfPO8SMETcoiRm+xd1EVsJonLoXjrR2sMEnZFtjYDGaTssO4U8ijTx6rlmYt9K3K1uxa70L
a1d5ehnzfqSYAQEihv6UpFO1zm7yEV97OLNZqF65N9fbfvwNuJOn8JaEe5FtPbDSAL2CMorVvUHC
+CtxEBoWN2i2qy/RceMrp6lbzhAOgudv/LaeMhPvObdsT5XTjFvGR5HSzggEJ1BFTK8rROdWVqyK
HL8LIxeKFBKPIEggumVnECr2yZWBIs9P5TSCmiF0itjJzn/brRxLc/76kfVR5nxdNfUZ5I4bHac1
KbpKCdWhzKTkOMX2/sz2YDMhVY0bMenQPuAQKCV4/nQEVPziZ0fmHJH4KfCx/NpHj3EOBQfIpiux
yny1P/NJYVER5jjNkUBDBSp3mRHhtP+60RJ2C36mh4sfzPva511aogoAwsz1E959eRuvmmIuw7pF
5VGYVSTaSqevKHLHK9gjMVHZ+eJAKYCu+P2Aha9V9KpW6cX9YIqCSnDR1XzuhzHb/4yQK5LhiHOJ
A+1Kf4V4+cV95InBf5Xi6pjUly4JCGtF+JxN6zYYdgkhqOor2XRQ7+Vsgrl9rD4eSw3+B8zBUWqz
NRwr1+TAs4T2bdMrEeY8pCEzUrDBm9SOgZdNmAH93UV0ENi1ilZ9K6bW5JnJqoEFZzpMp6kzJwjp
E/CGuajkFW594W8nVJo7w0FYigsAvTODDeqcnBWBW+VCyzp0TmL0xDAroqgMQxKT8PbNIjPIpYt/
VRYawQlBHzL9lp1X7jKh4cftkbUYPN1Kjh986EsfKN4jFEkC1fo02PJDKX3jK4Dv308kAds8skqf
ximIpVSX8MiNMb3LAuao/GLnbMKLAl2Mzc1oeL52aWR8aarzl14pQfz6A1eDPwHC3yKufiopEjwp
dXFCiJlzLRDdgyb6LNyvOSB1CcCFq8zJBxbNQv0B4MtY2iubeCZtjfhXdY5ljMSo07kgs9ldqX03
s1X7ahvvC5RJKrA9XKF9ll1XdAaZ7PPHdBQgB4JusnLS91rQoPXgmx4HvO8YVwJJbV56QyUj9oyu
HkPwyR1D9WwgB1PwXrz0DY6V8AWYtggwLkMnLa83qXxBuuVotmqpqoQr8u5GD0EHh1Ovs/4kYBN/
K51QOlY+KekmajGvGuDOw+TBTv49FQ0gPOJvOF+zVqqk+syx8nHxVp3SeOuft+pQlCWa9JLJS2Sv
pCbMUSZXCtMgWvrkqvSyOA+d4/rP/Ee/paMFaFxLYGIPf4tZhnUv5pnDdydIoVld2tUbq5QZHqi7
ZMvuunIx39GeyCSHrGI+f9krdJJmuXoGEIwKIZdtvF5z/7tL6cPCzjnv7iZBtR6M89+0idaVdGXd
Nw8qXd7BYD4M/a9ORdUqTFkhVixe23nZEy8Lj877IJoZjJUQOSUjodIoKuHwuShZ7vCT/RkUSYSW
3syxkuSGzBMUo+fz7+A9qEd1OhXZ7F/3gLxYLEwFe7iFwzfIJWsJkvz96XZmSUBVDVHYjeWyJk/P
K+kec+HWrjmXv7iAH6hpkWiKYxFL+8ak1yOp0XDWZa7D64uVHpEyVKIEOom1y2jMktyFVU2cnwlN
X23OhpWnZHSekLS970Bz/E78De6HVtZ/enWCN4z+ak1k4LLRmVVJRmNMSfq39smv3huLxnNoR+sr
FObDJa7bH32jVIt2yMVGUT8KutY8v3yE0xDCjAFbW6m/kHeyECuKb8kuP8ZC+vY2SAPZp7/bpj/A
wvsii32foaWv0fLqUdkSNdF3TO60Gtpi/wlPFqRGqimHBuQbhS8bGmPxk0/p7GgxQ/w271qcl2vs
N5OUW/1d/PLo8RYPLjw2LaCgU6r9oWGvRr6DO+YKqmSyRN56qaS0yAuLJyE36njeEsgvn1zrhecv
dOEVciSy122J0Blcq9ZgSvBhjwahtZpCXcrhYYJt9T0t315Ev3Nki4vdii9HCZABaSK+wUBPCF9a
/waNb5ms6zRwYBV+lXbYQCSa7kn/upxUth9EXx1HeAMj8JQ2fXMJtDF2F6OQkJjsN9rr9jksjCE8
Q3U0dFcgzpZbpsYSHtKh8grHgKcO/VF7ZuAvv5gVEf3jTbWwEaiXX2MmMrKv+eVIrskL7OTU0cLm
I0pyZDDYH/HcTHkAal7qY86CAyJTl03QHuk/Qqkt9suxuZR8psPWEL4fqKGE49t4rxiM/hKPNwXf
xh35GzYr8tJt9+JThkBrbeHVa7PQ0OgM14fBW19gQ1bz3rn10+5RHg8fDqGGTSjVsAjmV/aG4K1K
QNRmMKTr5OUPUFlWSUuONR403cLdCrgxmlwUiV8lmwlxmhclLjQlJCRUVPa9s2uQ6UXHhCNFqIas
t9cUoIhZHs6TuYuwVovQ9JsZOS0Oy2uAG1xYWciariDXFUDDuvDIbHEtCeNJYr39sWcK+iHbTEhg
PA26N4Rkn2OVzUCiMwBADC5n76bPrZytEdDqdnLva5V716fIuwxxFdK9ZFcP3Vp0wny9Xg30polP
tnN2ByeCh9kDT6dlyqlHFsELFNYorJmcG/UTKU3QXT2Y6DvfRkZWTTQuBqKFF0ZKSedn8Dahgbpz
aNMKqlH/sCpSMS/fCR76VY3H0hakE7ArrlUd6N0AlB02TJMsuTO+ojt/RXkTeuj0TIznRGyPVFnG
OkEUL8pDqFHsNJOE+LAafFJBYIo53G8kPAs3PCklT5PDOtCvNdHK6/lf0joAsEHZO54adoZHt5lf
CHL4hf44O4aqNyjYUh0d+LQnJjnAMtMX2Eg7ccZr9Gko3zU3vSmDTgU6cfSXGxkoYuUS94+xK++N
Jye8p4YYnOMG8YPzJoZ9PlaDqMaiGdOqGfUkK+wh1V9z4dKzzd1CFqSFMnANvfot3jvw8dPll0r9
W3xfFaraxDWGbYkOTxTy0/pNzvYQE4xi2D035tzD1q+ZQJSkf0i0MNzCvk7tQzYL0weYpMaSVZem
y4waVComJS3rAqQ50vlkRnXLKSBStqjtyCxqqK33quI4a8/NnRtg6/UDwM7h2dmXgNDZ4v/cLfX5
oj8MWnqy0s050E+BG5sX1w7NNFLgxx0MW8TnxwsEmIVFF9kIqernmUL0Xw95n1tXjKc9EXSz7MZT
0rnfeg2+r+wiYBuS9hPIxh8w19c4n3XHmLyJ1pT5KWVZTWSLRbC2RmA9lApWpDXKTXkd7/KFRb3h
uuhvV/m5He+TEulHDWwJi6xBOyN7Rv7d7pME2gk6Y+aU7owGGaFgRVo3apXR2zMs+lB982u+tgwt
0Oh6u3R6g4UOV1Co6Y219FRNoH9QHlH7+7R/Ef+JrOgI8q9p92E7kpUTE/OOqIztbq2e+98+aLev
7T7dk2rtejk7SkoYKXRQEoAsEyG8yxMdGKFtZ6ed2DfRGO/7IvgEH/TU+PSt85oAWyxYQSFimeKB
tAWVHD/33Pxo7k6tuwfDYYBkiPuJsm+PqwRFVQBHk+rk3gMmSEFCJ7kRgE6qBpxDEmQPQN57rvNN
JUXmEtnicF46slP4WVvOFUA21y3eOkwOIUGNevXF6a+/mK1xDO4/czfdm9S64D5q4rB8jhamWFyp
Q19kjSs4js6YdQQDV1YbDeo6eJw0b07UbMhwRcl5ua2UNedX9S4LLj4ujRLC4Ccd0II0bTHOEMmm
xZORhrRUeoyCuEzP2Nbd5vDAZbt3psktZkKAPpAC5DpkKWQgtsDMA4P/Us/MZy4b903S4TWPU9KS
gmp3yS0Rr3LEplMQ/09CRNN934L+qe3vFpu67cGC+mH94DDE2bYfCTwbkLhgapQErR0yFMg3QISL
ntJgIWwrnBdnCk/F2Hhd6gsFcorJolMy29cAYT/QueBbqW7NLAQF8LrfaSIY0vMRPcopBmID5Ddk
BLVdf7W2cKkPGdnmM94PHdOBf3hjrL9yC+qrIMma23LstQGL0+G0JsLGKmTiTT0P5ASKcS42OnvM
DWGrKvMwOMWzjmelgcatHurbR7VjKLe95pr1ld8lrNLSAXBTtPDz8gmAXqzGGHJew6wd7MixT/LK
PfuR9DnYn0YIOmZSyH1uNPlre0SSF59PSSayZFS940TS2AgqRvPk9iGL7x5heUhbpb9yato2Ofy5
OV0o+90edaP0sPSrVDgrg/99w07uIuILrqx1nCXPkZn4Tm9qRyQMNU86FWznmAWkszqNbs83GVha
A+aGPLlXkl2rFCxUgwR2ETafnjy8HoKw2BfB7VLkekOUuVWzjnAgVcMvOXMgYjVruQZEr7/iPDd/
yHA3oFYzqCq1m3x4P1X19Vj7VroE2/L6XISkQF54/pQJVY2HYbRF3eq1hq0On1hdkBo3VDnRE+AY
WFCXspobmaGpRgS7weBqSgsDS4sY1ypUYkxCyk5DpUOfAXpF3kBTy4iNNfaYip+CV8UzuZgjuppn
FyKqfmioT5nDBQ233g9mwuNaWktOSSS6lx4/LJdnX3JRGZarEM4Q96wfTUzp5FmdAYzuodmtBaZV
spTI+Fs7ftqDhPtA4QjNgzYqxpKKEUHw4Z/MITsyx8s+I6Ga/mRmDWea96NnHFZ8pN7Zlv2k13Dd
SmDOqlbtjNG3sT+p3RPW6MBn8m6X2fZtB3Xp4JdsqJ7qlj4TgqCpOEmm1FqW96I/qFuRTIczd6ky
kMGgQyV544JuxoHgzQ3azeOpIDzre69YqLea4aAtOnMbqVT5zbG6LOFOBBUGYS2YmkUWqfRWOv2P
00aNvxIWzSx8fKCzZDRCOG9kkoRoY3riAZir1ovIyf93+RdJc0cvOAzR02Dbs/mffj0JPlYSFTSU
2ChUi3jho9fjdy6u1tn3Rl/ARf1B6xUeKbbWQ3KzMRtzcB7PxxNWY9UWNeXZTeNemySJoU5TCf7r
72Cp1Vg5FEkSa3JTGPzeXK2eX5vqTMpzrHFD/UJYAG0zUDdujZMG40XXcb3ZaQC62RfdKFN5F3H9
zF1Co1HMd54KFS9NIAuDLtosEHbQ+zQUL6BKm6dts0e2z7Cs+5co8QdM+zjKFd4bruVYUos9sYCx
arq/CzatlhmnbW3pF30cWuESfdeoe9g0xpXHtW4F52cyuWQewQiDX+FUWb7ntwGAtleSYtEw3cEd
NpHxAbSejLne+yBNFk91dM3O8ySk0q0uDs+oNyyaR9HI9j52V16LezkD6Yl0LaAM7GXCfdYgaq/K
hddz6MyJwphPsXLgBBPc5wYamvias4fzdGNugFiu76XH4dFPfPUYq0Oz8LpGCziY0uBgLJA3paLP
fhUphLWynMJJ6r0tFx3zjjaGXpRSrf0RtXco0exweFw/LcMVnrDNfXzMtLg2B81iFni9yhLVIFSc
Z6VvAm2CyAG0cFh7jV3s0sJ3LvHdmtaFveZi0lPtiwA4m3jeygn1yduTILdAh8UJwtJtwtHg2OzE
Bt8WJMgIynj4cVS49sIBmLkReVSJM/uEv1aF8LWwtE6XPabq58MR2QPQx0Z6176T+ux2bzYhtpcY
Byd8imKHtickBBwTsIZXm+iUlI5KrUf/u6MU8L2XXoo2JmXdbdhqn3gpzUc0puknIVSSH3NfbDwV
nx9w8JnxDfuNzVDtBPa3w0ozbaSridDgCEaitUbGIp3RTobmj7Lv0fuLICzAZtE7UlAy2uYohyd7
rkwqu4+nUmSpp17WVxDOrQGI1QmDWA226RK77dy0um5wEozodUUFGYbyqLr7gQi8aNb6JR4f80Ec
GzqQ9oR51UjmYanUe6vpjrRgSYDhfSAHC6D6qFPzvuDHhpyq0kIB1mQJnbxBm7qM5gELwX9C4XwE
sffzvPCVL5GkUVi8uqD6RUvdWyIZx/uqOanrrfvzwxQJVOvsnO6Yh9olaLLD9VQBdyt0PtJki0vo
obuKDtiLtiUwJZJbciUqCSCM89DtktD0eF8o/XDjcWIzsdFFVq6IJ2YugaXW5rJ7ByquMCy0g758
wrD9JJwgEiy8A689BIDS9Cvcqiwww10VjGHWuJYl/5CLgusxrZYGJdj81ywx0VLo8kz9HIK17Sno
+o6rXZmA9bXi8iEP4sE78d4kqNqqpJOgWWv5iA0bTDZxqWywB4zHHinD2+YQF9p9SjanXi/m/ZR2
nPU/FWn3wIr2bNFBQt7W168EnWsYbiMyQdGxBiQ5ZdTs3LH94VqGp8IcMtH2CGV+/5BZD+1EwVq+
o71q1zw6Dt+a6iMyMk4LixV4mO3DiiyBTMtiv/OahAjqP+oXZFNJ0Sf0cKNylfGsYtEwt0xOD+B5
E9TGmAeBy8jHMh9ucPG58X44UEpQ4BYw322oomyOSUxMioKQpcwPFgn1bSBbdqn61O53902VmA0k
TKR0ZObMCeO+eC3eueZNSxO2lKQRxJ+Hqdj2wCfceFRsePnH27OJSA8Js64o6xKhwrEMHDGiQC36
6ilDgzEvW8YUbD/r66WV8Uj6FnhXHlOT2yFevCauPE8uYicmZcfUoAZ3uftqRW+7jADXNVcIVto2
zEqROcAURSFs/eAR6vFsD/kZbnqmDd8jQacTgyzImlst95r6ZV0ds+KDQTTspUpE8aYsE+pvb6Bd
JpLdgSj2fI0NBM67ab6XNV2UB3QfhkNobjG8jLa09K/rzAyy33bzSRpH9PuPjfzq7A3sZXS8H1PV
98O+dSyQ60tcJgmyeDKZ6e7SdTzZq20+6KgSO+GBH+YBqEzWEhGZdY+shA5FROiPopeyPREXRqZO
OPbKBM9yva0s0mcCtvUAcjaT8UQkrCuGHHe8psoWF9gd7u8zCuVJUQmRi29dNWU8p9purhgqmv8/
CBm+jLyBW8wQLtMszhfww0jvGmaxrP6hS8TEXT4OWCjexJoG/VNGCnS4TQDSY19gDYb269bkSwv/
AyBG0qQQOvFSofNI6y07y2KLhwI18pQCmDNZGsDu/frEqCbW/RB7cWCgqx7HJ0kD3tIbIdf/AbG3
Z6tAOXtR05LZ3fNzct68xBAQDWLmMtO5yTJpe0HIWEI75Fg1RwAq5xPFfUbGn+yntp+XhIV32jmw
qseVOyGtIzQYGsyqfSysyyBw5h4YeMd6tA+1JJ0VNU231F2PPDWmznersxINaBjpwXiK9fUvZT7S
NuYwl6cMX/Wyi2IaZwkZGVMeHGrkzulMUL/gLo9KqLyfP7/AXt1hfPY4R3wFRfJQ38f2GOK6jdT+
uqzoo7YHZ1VNzmJHDt2artkZjvCYghO/9ZChIEDH8EjGd+yZupz4hEdHn+msCPY5wRgL6WGJ3O2b
T0QoOJ5spTvYITzjZLN5pEv0o5QDWw9rg0z4KBktvlP+caUaDbPw3bd5c0HMLk9elKgFVUM76EIN
x/zqnc//frtYkIQegrx4a2obe0RVMQ5yfMQJMUhWFyM9gurT3Z6Dd1y9miZ7NBi47fqcf44y4pON
1EZQ7RPRPnfJo5im+CnrILSTuTf1QxzkZmx8ut1AHZnj++ucV38YTaUjN0Ln6DLbsyXXLab636dj
bLGVrcRajE1668ptArzPuPQjZD3DsuE6DOV5ZPoNbmzYWJEnUebKUOjjRxvY6+X2HUM24mR6quDT
q09O57O8JY2CPG3z6Kt/MQkn1EL7mLlZ6KCNPUay7ilEe8o5fkLMtn778hu04XgXeP8NV7jXIWIO
G0LCbNcRO8U40Fz2u6dj5z5klnAAXsS18lp03tYzEB7l+UV6KTpHWn4C5Gi7OOiX2it05mS10m0c
eR9sauSPfvHKjoF3fJRZd27iliM54FhCHy8mo+Sx7lhNxNpb/1cWirOXnQo4ITBPcUzswjKJirvX
JYFSd2O1JSmaty3nFgcbgToex0Bss1B7OSZ63j1b0UbfKhtvhy4ELdqXo1e+K6b5fTyz/qCj2oEF
XAXkW/KIKXsp5TnLDGvmaL11oYjqFMJCA7WyjVWL+TTrhCVZ3ujtczlws2q55LwxbrJ0xZxoJdDS
NuWB3UdDKqErzEdmSQxmKwYgA1YP1DB3D2gw2Z4XMCmvdixnqMvVtnuVntGIF5Pksm9oXQTuMZ3G
xm10EGeaYiiqtPi6bfN5dUVLp6mJ4R/kr/G3Xjtxvg1MQCX87qsnQB1mhETGAoIY1TAW/IvuO/Bc
+xNEeQs6wpEReDrmLQqo6QwF7aPLnlREey1WF2kqUk/ETkD46gKHIvTeigfBm5quXiz7y4RJvdDS
BhZnVPVqx2W4Oe75lUgGAzZ3SfT7y5M7KopYiTIGeee5ETBxf9c0a9eXTfb1yKDLl4o4D+5LkXy8
Y/DayNddfv3lf30Cu/kh/RhQ6elbcky+l9EfbcWvafC7JX8kjGq7N/oP/1zbW9a9rKtIHBY3G8jJ
h+jv2H5n+A74VfINw8/zDfT8TtlH6CW6SUKm/XKy8/uf1qQO9I2vigKVnP0NNzCvo75RIDipGFUs
SrZTHuk9rntpX8l32ORl+ZuQHhasKkPCFMeSv92J9E7/ul+qqy3wJp7fSJUY65+1juT9GO7yJ9/Q
n2yrc5VlfIlGPOhOTp5Eso9ShV4sdbT5kKjXeedRv++Cb2PB7z/teGbNrdRd4g6p0T+QGzqnO6al
sHThWNdZ8T+6+vPLaRcqoIIgYY1Wv2W6iXlNCx/Xykn57AtqcblLmuN4xLbSO3tC5t5stBAw01vG
h7uh2oz/1w7zC4LJ86I4PrEUTwFYURjCYmlSZX46f/XfqyeibrfVlUKlb9UmZvKt+xxadohPZiUa
h1BEFx+iX04jyNW5Z+0r3Cz/rKHKWPhYFbef71mbvUK3a5ai5LLnkaqbTW9bWVyHbbyU/nJsHt3g
fApSi4ytSHOi5UvfmnXpQ+YhZyWVmjEVIcVFtTeymRAuCY9CyQ7an5H8zyiH6TIyvO5ZiAFamkhf
pe+QEjrgQDjIozz+IZIRiB4XQBfm/SjsDdPvLPUFDRoN9UiVWj4TftARoGj+mSkMffPqhFHpmoYo
yFUAmbTqI3WqQsB8Jf5TNX/Upzqe60bmsBpw2Ic/mRLrhHvxgrQRTt2F2qKpKcfOFToVeG95RPun
6DEQYXC6971U6JCuU2iDM3qZGo/hKA0dc5I3hDNdB7oWJwNMaPgJA14Fj1WNuQye9nkEUiojiVmO
fmlWs6JEgUHMmj/ToAVtZKjn1TtzlT6mxcjC2nlXch504NbgVPpAGjFkMEv8r9VW9eiQnIg0ZZYP
Qxe2Vy/hNaT27z1IzE6cEKrOvfTbpb7uGlC1xBO4WBzbHRqVfct2CgDgeTF6n0nZcHqMDtkpXKhe
R6YcJ2O4dGAG79rIXmkOxQmuRFspy70Vgg09qUQlNaABiNHhGJqjdUPhfoNdOnqTlHKhpaOSFO4M
FKWIdw76r7MlCrEQGEPMnTXjDiQSHyl7nOYkIoV91IBwTHHFwurkPvBRwsonr90KYHrmCtAvGRFp
iSu4R4el5uFVZfv7lMmfe81ohpY79pIrtnRG+SMggXJWsMqPINPc8KAe7aBURpNJgOTMHBcIkrqj
eVpC7b1ef/qw3oaiMRwCxSe5jW5g74ac84xPR7kaAZU7sS9pIDoIMEnBnVUJzm1lXsftXaSEspdw
gHxXpNjCULX+frUGFx8Bk3dMLrc2ywRFgv1LN8DoONlXyhbs3pLOKfeu5SQLxq6aSKajUG2YHukx
iYvaUntaaz+oGxPn1jkWWePBZq8Vd0k4q6Rgp6pb6J/kafb+9HCDgm38N+/z+BQVmjxDt4+B0I+F
w2WnWfwMvjOOG/V1zq7WdcYemKEfd4NiBwds9dzxMTA3/TUCYLWBsUJnghJvlQ/DFrqYVjsGjd7L
qrsvL5wpTtbYZmaJw7dyAhutbvPfDVaTrPMDJYsd0QNZYKxvm7M14hmmYj3VSlo5DvqBWfKvTx7i
Nm3Q0s9SzIrGihsiJbn3DiTdlgPU4EWiIHHVLQNieUj8sms/2zzCpXWNC/7uJvuve1HAe0iv9Swg
EP80Nhc+2ZAJZVsh8FqBI/DKrl7q7PV47gVa4xFcsPhAlwt/TpJBmUMtQp/P1IZDUausaxTlyuMF
Jcl1ejhuP83kS0zTTsNBPLALfuutDagBmO+GIhSUbvGRzIfnVFLA8wt+n8TvEluRwizVdD4oV6Ec
1EDEGDGNipcL1XfSbClC7f5tuwmG50EVZLi86nCVRw/eXSjMnjdmW77fs0Sg63yY1A2G9oiZxJnx
pyk7erQNVCfAlez2/HpTP+XjiIjBFF5pcETM/8XHApqnZQD9rnwv606TAwfdL6KthHATzDvPyEOM
0xWWFtqVQS5Ifqf6HA6bzw6SWAE8DP3xB8v1qBNtmx0XZuxKXqQ/5eaw7xwV/l/SIiT3ZmmxmvyZ
pxqp+s2sza0RT9szwXBGCV1+Fg7vtKtKhUMYM52irMLiK1Xg/KCqaFE1YSxVDi3zhz3Rypo1Q98N
7Z5kLOFHO4Dxde7PW1kfJk4wdph48EZ01cX/JtZlj1XbeBZGbG/wF3ZlT1HEIGY8NTqYFfer6yfx
KbfWl7xMIYudAk/VvhbcS4m9k3xhixEcD+3unQ94wO8D7WUHfl1UmvlkcMslcAYbCRZN2Bd/scTC
WtR2CrdmD4V94RzOx3VubUp/tBhLTOsFxJECKTCSXeDdsfWSYgIoTRSj/oCddJttryMWeJ0xMiOI
XcaQ0CN+A7c7l5MPh7ZWOo82hi2phV3NvS8saW2Iq8QnNdLt+jnQYB4VnLDBok8wluEfk3E+QHBh
5K8sgVwTkaC34WQlEQnIyLZ5LnfrTN+ul4vozKWMMxcdRu9YBroilRFUv7sN8+vj3vKSwZ88xscb
wU3kBb4z03KpZnl00/atvVHBqiVhZDou35wh6vRZsExICTjHxAC23Bcr5PXEcAP0Vs6nd2HFi7EI
ZZrhddfjsx1wOcLGqYKw4RUsgUueq8ih1X0XS1VikdU9pq2Wjm9TgPU0HGnJWqBD7I8MXxwX9Ywq
XKi0bUll+RDyct6CjSGXza6+ijHbfA8q8WPEe13GeXSsJvnoDcxIuTBvs+pJslOOLwnlQJw5+9wt
U1yZhlOelWxO7cAfCjCaEdXYfCT4rN9fCobVrCWgXKF8QpYytOPFzMkXXro7vIQigI2If0USIrMq
jldbCPdH4JbFq58NAkbaJ4Hp2CVBNxWsDFws4if52p7Py27k3XhgLRAFOr1uujjqXOhLsJI5vynA
m9jOoN61rWitPBv/oRvK3aUfS5jiKLzUsGrpTSnbFwFby4+jQ3OD7JUlS82p19NqApiWMogu8548
ODZRzJsAnP3uNRcVnYFHNseu3SRFNtfHPtyk+mxuuf5PMSlFWpJTbRlrvuqI+3ic+4LprBeY8rDj
JI34xT/OvRmw3IMQFNb4hknrOlR876OKr1ZKKzE17pezKStpUu5s+fHquMRO6m0xlGbSX7zLP2HT
81FZT8XlcR3VtyMATlTM/YbeA9EBsU/Xd9yPE6LFeIXRogrJOlp15Mp2WzhVT58idX6USxmojGi2
YuPMHyczCrvK7+KRRVFsvL6zzDiPCrXhHJeRsAx2DGdK43mQXTmQPiG3+sEi80NhZvqf4ay+jup/
OZhfCpd8Qy9puYIX1TC4nNxxh7UZbYHE9bySpJR0Be291BnRt+hDrUN2Bty0eF8NDQAz3xguC5Nt
/wWIha8WVUjNcW+QtKdti8iNlUmN4rnnOWPLDorI5vrYHoXoCIygdzG/syg/Zfd8WvsT528i3ySU
mqKIz9o+Mfzs6UBGG6ydd34KGILNYxDiwLzESTb6UgoS+A3+qTLlkvyR7R/KWele7z0l+neCEAW3
ckTX/zLK8aC5OczR8GWFa+xZ+SC0B6oiaK6AB+0/Uz4CU/kMIPfcEF65zGyG21CpqEcwNyaQob/u
31Cz7ibi3C0/cI8sNkh1B05e/h0fxTV/ISH7cweizXw/a15dJqwlvuCzkNJnlQNYv3Z61fVzx7Vb
nTrkNbeUQZEfzhqZaqTDLhJudzUxDGGBG3wDfmVCxe3XJdqdpRW3BfxVlrWMPt/TROuV5WcqqTHC
FOkLLtWi1BwaBBO0FRvwZa+WppIIc1tSAprtxaFqOxWIyGg8GIbAXl0phmRuhlm7cuS6RmEiLhU1
H14I6lEJTKejICCRMtcN+ja/mO04AfWqetdILuayTnUvzmEl/+Wk0yqdWzSepHWZvrfA6ZfGa2E2
JkGN1ZhpS5puAvZYScz8CzaO1sJXAghgwFmDXxy6j+8X1eCkVesh6bKz0IuL6Mpmc7dQHvBdMg3a
JiLw9wTRnLRieI97wpVZwd3Ir2UIqZrhjWG6F2XGcQosPOTe28pLrzXgy483EswKkdxZcSX6o+mW
I4K2et2rHNAXiS+hYujIL4eMmy29TYgj2Q0E/IYG+9K49Yo0KvdaS/JPm5P+HKOfchzEKRr7mbk1
uJZcqJP4kZRdZZiUyxLh2pdFMsbwav6ksEp5dLWPyLIHTmy9iBasYAPUOGqVUyo9bB9Hm174v+qp
4/SUn5BhUK+96Dg5a6fEBnzIgksUcgAgOrJq+F4BjnD22oL3+erzBIeL5wPl5zpd+U+Asqrb2BeR
2nqhUueQxZdPetj3woADYNm8A0fgiRyIaXavwdqck2iXLhGyhANINqz9f8tcsJbZNcEo33akKy0Q
3RZJD/WOcnrjW1faZT+3D9FKPRGDtczyqpjvSz8kx0TW39BByrKDolcSomuVtsJLHVoLeFrVanu8
PWj2AfxWdjqBAs3zC9aCl0KCGCBeTpQ9kMaMuh947pI19b44Xd0FUEqOCvIQW6vL+t1WiTjm8gkU
TZU1A76fW0qAJ4sdAuEjbt4/bTP05GDvnCKg1JYddYMoYGk6/gKOEcBfKukxWzzusQ0HE3UNDA7P
4HfbdZMG2PyvW6bD/cgIwxk/pmqgp0bF6bzrJi7MPGpxFXtashd4M9UWJ1i2eLy2fNmwDcGg7jMp
cfXusrKxbFU+YrMxkyUqr3tonRfqY/z6nqvpW3weGovlCSCAT3iDWXHRoHXekt4RtkYcqv/oLvsq
PiJKDqjWMf0riWIXNakf8U4CP3ulZNhLdSh51nZ0vJWwBO/yWQlhpskiEcCKIuR4uR0WXFzKx5dU
HU7taQdYPMfimWDGZ0h5qZFWryrxtjgUz8PZPLgDO2+XB7DWhj96TGRIk71947jGVBet0WRPWG6L
P1ah5IS38WKFnmX/H+zbuYeEKfCfoTIap3UyQ0MQmyJd0keuk+cij1rJbzBY6tDg59KDIxj/VIDd
Cp0NGgbBV1/8G45uF+RAP6ZForA/SSTqozfaHkk/DUDuirmEBs/AMvjC5+DTYKbtSM4+3b79ieqd
+UZV4ev9/Sx1vAj4cyD6denWIH6kNSCB5mmL+h9sTX3XEezNGH1W5A/EMJHX626h3qzE6Gs+ncI6
OIdxJpqh4oiC5trvEtFsaD9CGVfBOJonLG5MTpsjBI0xXfjOFaI+ipuC/3ye4hewGQ2XX+teBsCH
Q5vl8M6LnjaU193Zk5ZARqZZ+K6DGdADBjskfogi2slupPMa9T6C8RONjpDAn6ikuTBZRD5KPIKy
mSmGJ1U90b6DvttRkbPdUcI/k9Gmiuzp2TOlh9FvT4lIpfroowr8P9D8s22ntO7JRRRW3B64Ym/P
BO/JdKYvHc0bdKGavliwLtHhqHUco+zDS83LRsdTmvSamxMd3TPWd1AIJ9XPS2cZwuftegMVTdm0
yahR2cWe+UgbY3SEQmB5PMSR3b014JgacisQ655OIm0XpSq/Pph5c46BhZtOcAn1RQKi1i73jofY
/N6MbxMU3EvdEvjx7UWZZWPaebcHvmWlz0P4Hxrz6LMHeRQaR8gsMltvQkTf4ASzZaWh8bZEvBKo
6agu9GVxWIVdppegmxFX03mU2dohqBcTA9NERbMGXwFY9NrDiJ8aiIIBWCDac4ySUkRljRQlpA6V
WFqAcyFAsYyhCW3uI/zekMpOW54uGVTwK7MA1ZrVgHNcLhR+Ec1GoEs7RRp+H2JhN7X/JVnJzXaR
57M/oEQXsu42MJ27jS1ms6GN0U1ICCGj2Whf6OK1gIa+/gcJoXV18kXUmWV4exO3qOhYUaejGBMr
LpCCU2EpgLjVSWKRw9WGY5hlZuJagYA5CWauystqAkD2Gx3gwcjhVwsVcNAar5tBIe/Qbn9xZKiZ
uo28zLAFcAhl8sRVeM+tNQECnqkQkm/wFGtiLKFfRPq5x+mUl6rcjQ5rntJ0BDvcUNZemPVj7GsQ
fwpixPJje5xSM0CkwF57XwBQedrSJZTyVTmZBCkM8TmxHp2FVRl1fLT9CgsgAyKXGm2/guZjQV9O
fQtekrDdw26oci5H3kbJZrEKaYAhWHLgXs7olrpKJ/8qTgufdrmQ/GDopxCHiz9UWnTz5X4k/BEt
FR8f8Mq0DquoRMG+rIRmLy3qhEIFJzEDy43qHDKwlgri/a2E6ovt5htqLJA9EGbJpu7BpfdnEEds
Qi2YAq/HH14DQYLurW3kBZMWS4nmK12JIDOacUQaXIErKC51SS+NlZvqsmpIuXoV4UiImg2XN51P
F37im23JkegcIZlSjz+wHwRGonoHEghuYgyAmStDym5w/KAcb4SA3PncnnA8ikD7pJbvncMPA5yJ
A10JXn5O93MHM2WyyR/YtD2bSwLsYajib91lt6zPceZ/9CS8wusXKc+X/vuWLh8wQDKmge4GMCrJ
i9xkMA/zPs+dPvnidpFJ5AqH48DXH7/GRCpv4MBe2qyw9PSOQWIziwCeHySK0Fjvb+WxlQGivc2r
a58NhmZGj2zlD5PZgq67VljDl+VUdTO8CNMvgSfRbBy6FebYAZAMHTWe0iOmib43BAXS5rEN1txk
YXM52go+kBzvRIKlsx/6+HERqom9FBfZCkJc53pGArfdAl6Hn2RZNrlNeNXx2HN5GjgO3ZniYRt+
bDin1ap4J8QJTuC8Kmc4MFPFRzOPF4Cdb0/daOw/OMXYY6mvmQngIfdljd7KV/yMDzOoxBcb2L9q
jvfu51knLoLfN5n9VtO6uPtmKs7b8uXDIO2rev8EnOOtI8e+Id+JQ67uOKWbQ0O+jy1RGxk8DOPx
vDewsdSIeUN/lsIzTO2bsyexrFjBjY8+FKV7k9FGVOYPifH14wP6AyyCFtq/R1aub0AhnXfrR+xA
jCiv4QQg7zZZifLdmBtZOjK/Wn8GW8tPFcyyPBOutdeijs6A0MjtPWbwIL13J8qiZw2i5kN5gBIU
NS+dFv6MfmxzEHs0PaM8DwY3dKJG+ADdEgP1PjcaldteNIOJvyn/SFZKiV4oBDWHP2klnMu61JQo
yjpuhIuCBbPCkkNMD4yZO3gvKJLNM8LQi/LxDqWG+2Q5dXmtQEwl7aFtXT5ISxLkn5uEmZLQAcPZ
NOIoKULWfXOyCtVaJBTAm6I4sKoE2cQoGPBN8sh5Z5VIHdHOOAUMUtXzpKl71UsM39eO3VerMmOe
HiDrV/Xi2Ncwo5dG60WPMD2py4Jeh8+ELUCgkhl9vthiZLnuH2ZIMzrFTRDo7V8+AtnyiCC8sWNw
hIeA97iE+Peq0/utZVCU3Ucl6/7kwesnjv1r+NFuBtzRSAn9+94Mkjw0GeP/zib9nfptuV9UZ9Bx
cmMqkrXE3P18YNZpVBPj6h6nNAqAV2kSrr+zuwKYDduf7T3G35u8TR/7D+deHbw2pXIq2dWJOEJX
JFicUoAeAHa0TdXm4iwHRUeLVK/Q2In73aw6HtKT41/ISwNwvA0kNRvwW0p9BLXWfJKVHfiSHYl8
eONFnbg1LlN7FHKJ6Jw5bRqop/WrYfPSKg1GOwNC+YjVKT0v2cW9qM8hM0BlwvClvFNLlM6vvW8q
krsO8qb1TKv89Lt91t5Poil+JQQrsKwo3rB85JSrV44ERMihXbSqurN+n0Z//+nEcDntuqyEwfC1
9Ez4tEDlQDoBwCosNN5EfQ9iOqiMujJ+nYwcOUelVEji0T7DP1wdUZ6E9NrUcKGdsZfbFjtGK6cd
nOhtzAXp5UM6Mc8zYM7PKPeC//BK13ssWhKa49I8S/NJNt9zqL/qpdiZzctCtxRReUCWmnauQZ9S
D0vxjRrTYUrt1dIOAjbn7Ie5rRwdBxoes7qhZvhQo9MXbKX/vrBE5UFrRHk5wORPxL2qasy6NF1l
RiLZMf6dzuOyJv9AsFhbJqrKedDabG5+5XZMiKCitVtRf9EqnnRIjvCKSkfBzu88nlFubWwEtWu0
kKOX9RHiByIpxb3JlMYxBCrJAGG46DCDPnpsGsCPCoj0XH/kSEMDlBQMmBKZGHAnxSEDqF/l8r60
GE3M0MYspvWt7ctdWx+jFFgr4RWgO4/1QIOeK4zjEHRtKutPghHQD8qUqgSzNBT/xNztCd1ZRavp
gFVZWf7XeEkVq+1c7WeZwFTCDlX6Rr3+RPyNSgnevoMQsQGMm/bD1fqWM626P/MiWxQYomm3MQXE
OXhTCVddY/hWqc6lZli+uieVCkgoaxNmW2BrN8eap//QKAMMBH+ofnGOHyjZIGZ904YkznFXTuKT
oGF1WyDrFk91tKxp8tIAyeTUkEnooe0/I+psbjtYrMMWZJn9BX22/yA0xoTM3tlSWnHoCE5u+rxu
f3UgE5rZOTFP5F+INH+3HIaBVMKWfr4ejrFABg8+Akxy/fwS+H0EYfPw/nydUsqdQAT/HppYbFrY
lfAosNSJK7GulvzvfjNFaNWJYZS/+EUeatumpL1Bi5narWCyc4EZS5il2kUrXI/BXEBQKjvMRCyP
Vh9cYowt+wbbJQukXPDzf69zxKBZLbI0je8NuhbqrfKjGZ/Bd443S8dUfBrA33LyWi0CDKulnEPx
tF7CovYq3R8NnJ0zZsVjciK13JsbVImO5qVv814Dkzdnb356sPaE0VX+NXktKrnCZUCZvsA+hUi4
Jab7U5HFd2LDC/+AvySww/iQKUSvnAlVebZ5g33RNhe31YWwtk4v9zCyl+QOFX12T7xHyTT+Sn/q
vB+hS0RSfFHnaRSX8Z5SBs5O5+8Pp5H2azc9D++Gkklk//6p1O5mxNe3h1mvFQaFpaF73IHSbRyd
P2Xu7JBnzI5TshV7QZ97llQCr4IiikoxJyGUoHK9pXPkjx1KsEuwcIHt84nIr18TzMO3cB1DmQOQ
1jSa924k8JKNkRSMyBbvzFaUuHlPUr/pvYuyFaXyAl+LbEjt6z1GXSaZn0vajQKprbk9/6z0PWLr
E0ARVwLHRG7POkeRYUbPWP7IMhwHDU++s9xiqfY53/nCcFXEK5FBuFhL0nBxqKgWr2kbStnUYhYx
jFhC5VgJ043V909U27WqfwO+xN/dhJII1S6MlRZ0h2bUc3ZhO/4GDc7Os4tpAyWmfTmI2dx97GEP
KUbxm7Ppq5XMbBqO5EVkndXZjnCnO0nkZjLqwlkHwtLgceLWijU+aVAImYHaIntdsFcKoKxtveAG
F8/VPp7f8BZvLu5yPXyL+BPJ30muUzAWdJhij7d0DZIHyWs/sFx1yMiFSIdMvT51aowvmZiwuVHa
5UW7E4a3Y9ygizobjzc1BVCNQ80XbZWSBL/CxK/6B1D/kDcCDcxv5E/YfQpQC7j0tkFIWnTrYI8j
2Fte7UIrzd32+B8VMLVfZCrlN77agcSob5/usqAAZZfs7wNWKzZRlzTwpQR1rnQ//2XKogMSFFSm
3CYBXFDEGUBp8hLT1v5Hpd10Y1oyi8b88E50SMgg0QnwtAtNi0bEMGMsVC6gfufvG/zJq0L11ip8
L9GABCxI67Sq99e4U0Gcyi6hqSZJwFb74dTS1jU8t+0A+DYwNtla4U1f1q9cJYVZaIjjjU3xeIXR
2ZVeX+a8XBVl8J8ww+brYWiydbuRK42vf+ENcSOwqcR4wGe43I0GnoDacFAS+c02UX8ogZVu7AIQ
hskH1xE1hBOMhYcjuVU22xPZ9S0Yh56j5SN5kO9yemKdFv86FNOBvb0jF0XOD7o4uysjhnbXa2cV
xG1WUIEfTG+0arRGWgD0nSlIKvjMg0MEUK3FJBpINdX98LXaLUl0bTZMXTaQ09ZzqDY6gZCxhTGn
ABlYKtupVfQSSv6Xn+QynrQvF/5fYHo3U/cH1RqVPy7uFZGJys7Aoc+gbgQGNn9iquc6+1k/hswz
G2IvJVmg87/pfEIJEsOjy/8IXsoef63NomZH7THqs/bcx3CWb6YcFY6HIRzFEmPwrtUo+BaeHmpT
+Q7XlfNeVJ0GcLspUzuzyb/c1HkFunI+xqYyRR8VtNRpW5L1H0jHbvZY1T0u3ZiE9A8vQZ0y1BvD
QG0XKOAvFyaPG/3Js37MIN8+h24+ukAMAc/U5yBRcCVCIZ+AvZETc4yQ6OU27bkiOAMoFSeVjmvO
3WJj2cwzTYUa5MKKX2KH4YkFyZmv/MpD4xX8EUUeTfx6sQOk4N5zA/uYz+ARQL+rUdL189QWesQp
1iLqERTlIlJUIu44Ao6OAOHqav7+qJfaRbUFeEKwP+mTfbowr2ZP5JyKi6/Fn3lQL7R2RbozCeKb
mnjHGoMWcPeuVMJkg0BGiNgRZ6WjgQzw5pZsxDUCO9Uk/PPSpL6yFu4zdeJindlcp+1k2YNckE7M
mUmRJZBAzgeW7ZGclUQv0cYLOd7dc1RjNM6W9qdTmgVzcSEo99yEMfq2hFWGmCIzTmIkypUv1K17
Y+hPSHJ7Q3HXg3v5Zr9FPGs7eqlx2Rm8/4UktkRnzvjyUMksGrM5Uhn92P2UPrDpR/GOBenoS8hn
PexAspciP76Qb+nMhl4HYUWoeHAKLUh9YM8bhk/ft2bt3IfbkgeXokVvd4MeJQWTkO3jqTtKReRm
LwhE/3lYlKGKzLpUNwK8zjY1HsRiG1TxE/5UNDi9McDQ0CCGjcaibiVgWhch4H9RPFr1i0hAi5/q
PVIwyueRfEYK5+AYm/y8+G2Q20wqgR5j9kc5PNWg87oAv7Ddu/z+qet7eU9CvAvXBj8u8/+7fwlB
Z5avp1rYw/4s7Gc18wwgoXzQTb3HOmfnzdTcx/nY2xOyEiJHMZF+QTdhFOJsI0Ec/JGDfEAcMJGX
JtbHa8hMcZI4LaNmlkmfl3rv4jxkSYeIs6VQ8+TDwRMxsEoQ3QRB9ZHeSbEDPSba7m6Rfpvg0AE2
4AxWhDGk3iCigbpsKEr1moyYsgV0/RZf4SkjcHHppWWR4bo895ZRbVpGU3QsRW5aMo23auBAk+f3
rpF+akzS5OOpAtTq2UPdwfUA/hF8ojhcaEZDpICcI7ThRBnrJzen2a+IFdY3BFtnF3cT/ZT4oBz/
RsNORZwVoSU6zXVJx8sVX5Ur66gFKQ1L1+Tws+i5u1poACNPpZLnLjOwSkQKkF+43e4YNAOuf+tP
7yYeR0mgkBRVHe38+6FvxRsv9lIBj+HKzBlRUYSr5DGVY2/bv0yDhJQ9haVbaOz4umL6KVigznNp
9DNxbjLB1WW6r8GtGHw/14mbUz5USYfJNKYOnsMjZuXHCfXgBfvpJJKqZ5Q8ftoSrMCKrDpF0t+V
1z8eKdkok6wsiycY2A3ZzH0meRU32fvcSZkB2vWcLDpWWGBPBsnObfWi3APupmSo0k0npCg554U2
qL5kvi5UOpLrVq4RebarvyeMN+RN3Jtj34ja59nPNM0sOjN7etJkvvYG3v7nsfK/KkdAorDLu9CW
HE7j/R9L4NOG9TOBxQQI4AoGiCXT7W9//j3S8B0fUel/2/RTSE25sDjV2yK2Kv8EwUfj0YuGdyIi
Yv/VZq3cJA5e+IsL5LBkD4BJttY9BR0JLJf+msJTFfCVYCR4hSu6iXeI9OlBXC2TGTqWm08Qgkuv
PFH379SH+6xDX7Jw5VGLN1txI6VnSNWNyQELe1AYK8PoeRmeYlFvsptsAYmBVoRh70GEQ+1lH0w+
PP6StMFH7cdeL3prNSsBl/s8QOUdcYl0s6G+ljMQoAV+A+2krgacBJdNxKjOCtohHuUOso9FisSd
+nwVQKb2SFnsk5LQJAnDR44U34OkvhAr3xKtgKyrJMSuFeczJwpFo7iHnmXU+rzM/q6stRI1Xj/Y
/rN7aMdEAh/4+ZVm8urUuguZWKpip9LFatJ4ptzyA7YxLSckpPDh9+gtATPyTNsqkTtFdjgbdeEe
s6uoLEMAq9mJNfp8ZTjLmtaHMDvoCXUZzXO2idAQJk9kCxQYFbz83GAh9kk/NrT+XrbMHRIMQD3C
GcpQJuj4jFZMQEft657nAbHCBz+cHUrszobiCs4ftY/x9Vw9rG6Lo+t/AMxLbarqE0qlkmLIZazi
VWcrSHpMS39SCwF/fXFmas06T1qX94F8LB29+horc5wfy70HQoDGpEyoyUvikSWZNzEDMWz/8YrY
eBp/nuHf+iSpKZqw39sb+1LHLIkjRLmI8yOpWBqCfE7020EPB75DiJtHAvO5BFVGvWwH1TMM8oFl
TFIg1r7sytu23FZnjcGxRbgOBVaIjIbhTU1qanmaL/q9snqDrLX8ShYNhSWCSIKL7GfGPwrJeQhh
yQZ1T1wLcXHANfPf7wXIxAv65TmfVtuMfs2/juSsJ+1Ikuwy2JlxHPYg/fpKkRMen3hIto0v0Swl
VkRln7OzGMZX1bBA+zFb1Nap+2rzje2YKZ5CKuYFnd9HmY+IG1PztkIJthAQfVNsbdPlvGt+19p7
CCJY3N0Bhrxc05crF3zMPg1OAxzqLYC69GmWOiRXq9MwTcsbd3CkGtP0xPxpIZOfwV+J7HPa4bW5
rYhus61tAWwGcDS71Fnf8whzpOajkT7HHIMDLsw4LS0wiZawzI0CuE3p/oYlVh1BZMpo6a+o+IGQ
0z9RJjWXoQk96GDNw/yW/tv3d6xn3NUsY8SY0pn3tlnAne0TYwa1JAtMIMKTHCwf80cmwcYIAv8e
fCE0DvhBUsoAGPeTB2QLvUuyixGS679B+YcjmsTFL+UZtPAiXRX7QABJhBeO5Ha51SbqQ2YVaz+v
OXHCcODHdXhpzAeTtRIiS08JwOSPZvmdv3xWGI7pHneWfrlcl69vQVsLY2/b3BTQHDrdsJ6OtEB6
Vz8Q8YpSMQZBqKgIyDUGDCZDa4Z2qcAFciOjZ0sfLF8X3IzH8NPYPW6P/6xJbBr/szPgYlEUsgsn
UxyTYn89bcQyM40SvMaN9hYOsZ7hpgPomBgD6YGp+ZfBLoJXU81sX2Uddu4TTHrAIyHT9FceVT3J
7pn4i+FuJ9ewkYiL89Cf6sYgksFkEBK8xj5t3jyXkKlOa+QCKx7F//vo3rlx0UXg+NbSAxiZPm32
XIJKvChmVVVI7FzLMzQVyKXltOtNtdwFjK23y2gFtJOf42afq948Q25uG+KaAhP4dgX+kcJi+g5h
30BZd+HxlHBHtLt/pakzB22XWw6KIlv2XlpGaoDUiwXpZjMbjQDP3PqI7GnGot93LwpZ+cyIxJ8z
ojRmS2JFFMNbIH92v4j1NpLOuiVJmzhRlmv+KpLwa2/lNpnc3RfiNRLL0hQzDGfWYMgCRAsRJ1Q4
+V9mP0scD8KSkIRz1Ci+Iasu77apc7zrXq0jeu5anHxhMUVAUFoY45sXVb+yEy++3j6ybNJhF/WW
E1WkIfnBJ22XKQ2Sdu9roKIBLoPQDpPqDTw70PXUG023upWbDRQWIvtsc4RKACLpM4SbkaVMOndA
5knB0jUyboWAhEraYsaqhAak4n5t8fYWlwNdResIzzZml7t1vu7vrydmfbUV/l+neQKAtgAQQXzP
079Pfn/yOjmRz8GcAkEQaWtdkdkClZEkQ7U0WyvtXp0DOOqL3CpL5nwWAzMdIvnf18f1iZ6yXLyj
VAvw1rz/CeESEfoFxZ4OS8LIhbCWXmp6RxVLTY7nSXLZ6PqkHYGyrf7t9i+3KZlMxBvKmJrRO1uv
6t/43HG8njS9oY3InVYeyU7OISwl4GVTYoOHxC4dWgo5SOzlcFTC81aXxZq2xu2fPEqQRtymfw7K
3LIvWqBkZMSwXqMeyccdVKl3cJ/fDAe6xMZfgpez4mSgt3VVVvDB+EufX9Rcm2pZevLSaewtxxVY
KN3DoqzIq9ke2MN5j/ZiUJakfGcuLUU8z3DdkLLunHK2X3bmQOliGJrCkmgf/uTOpthFGs9MUrEV
rVsk0H5iB3uzg7LLs9aPegBJ9n2f685BvuNJP3DoUrdAe6/WK89McbuwionCMrrw8V0+UkU0S0AL
+f2Kyts3qD3Od8hsa+TRfCe7k+CCVZCKTIRvsLiDVY024N8x22gE/VklUwWjLO63TgdjxgmbEJJa
X7493csyIIW2Mb9Noviwcubaku+Grwru3jnR1uHViM/8qJu6kpi7wEN/n8GEHzT4XZ32/IWqtEZL
YyUhEesN2lIcrSA1MBislDbhVmkmoZS3TY3dsbx+e2D2RPJ1YB0jc2S5Zdh6LYS0zfJRZHocX9Wg
zA5jroui5ETR2Mv/QnP1PDVE80W3I0w69NIIyCmBFA/riECJmzYNXK2KDltiANcqSU0CnbvQ+d8s
ww+3xBOWE/ywCQ458qNkKxD8nKSyusSLWP55iAaN1u/+DcTNdd6NYa459QvBH33sGrEzMRzLFnj3
ErNuN/5QcnhShnWP7YZ2VnxmKVb/U9/nqisYrSQuB+zhp25GKwzKPwWAqqGjN+V+9pfwQJqAFD3q
hHmffdc8S9+b7q0UEeuAnQtfbaI1cAQlVl/k77dQd29FgM8ZQKcw/fqtmIsUAJf5i6PQb11z2gah
zqQS2xDgZcdrJdNN8tRlWc3Vj0qQpj9CkJxW+yIebopl5WZeS1tw4By2P08Ol4LcBqxjLAa7mkWM
Os2MgHDjpcGX8lNE5+W+GdBZqPNsL72kJdqANz6GTJDB7C0WQTQ1HxtPdLDvK94dPsHuKtqQwByD
3oDjX8dG+cfyTiBUhq8Aaa+wpE/lDgk5ESSaNN94Bil4rBlOR1RSMuYsek9VATd7GHfYLWfT763S
hL4S3sxsn74riI8FuUyOkYkV+ao0Vxnrj5+vyN+w0zksHwfEciPvnND5n0H5xNRDbXiRTDs08NDx
Bs4/7pwOoRTDG/XtfO00WHXGA8lNMc7DaHjmV3z22hg9DMB1UgrePBTX7uEyDqeflXQqysURjQlF
YvTY6zHAH/WLFDcm4TBady4YP8zpoQ9EkVbCItGKr8HOPeesIQ5z74eUbjQdN1qYU40h/6b8n9ma
KwBeECQcl6KoSGfcZEaQPGZR3rXiWlwfjdqPYG/mFl/k5UnaM6EK8LB2ZFZ78yLEtqcXSwvdTOQD
MNGv6Ing7VkDlYEVGgH7pN58m7NHrZPaZCOxAO527P5e26CZOLCtZBwP0LXXMRCiA6203BoJDyle
Z3gVzVxZmCrVdLDVxPiLsCJEFEklHes+Mgcg7rygaRumJpaDXZ90aJ8mOTqPfWVoaD5uj75EoU2u
WvUwFxEQAopO10UjOmEjUV8ROcQzHRWzfyZ0irewqlBodaRpw7BPwygTiYCaotUeQ5qFELhoiCe+
UCxuGpg3eDm3L2cjlu5qmIpPVrJjwuR8jNE/R6dPBvUwcu9S+drF7A29nuqUTK3SFnpV+2NaKY1o
zQu7sjWKGhjLSTX/gRIRcLpRYBHdDMB9heSTlGRxT7N9cfttMTITMqHwDSvpzAg6ZdQUjnBdsIaQ
BodBWsmQJ1YAQcr/FblvcQb7t6zN5rnUjo9N8pMqV+KclFIhHaTyBw//18i2ys5mmKY7y9xQvYte
a/Tc+Qkibx/a0oenv6SJZuVPy7bPAO8OR2CtZaDfR5OsQG9P3jUYXnEp/3yfEee1b3eVXuwb5ynL
sfi/izTqYVi7f1icTzcnCkFoMU3ARd+vh0dYn+Rt4GxJ38Wm6VhpPk14rczo1ak6h9M/tEtPfkUr
/dENxINVdHDIVESHrzqe40eY1lqiGhHlNyIiI9+1P5/HaEBhzHs+lHOQ8iNCzV3RmSxhtnY4XOcN
ETym33//DFNMHhxKUJKKS18it5NJK2+8ACGHVh0OPmO3KJf/74SnsB9kByxS0bPUP4d3+Qh7n/jK
3w2s2TR6h0vfdFOvqFdI9MP/MRebI9S2LzqUAT6fAGlK1spdLTJo1Z4PgWcteKKUSA4SPxzHlmdY
eYA9xHU9ijQny4/k55QjW5ZRMj/YclKLRAzXXtVzkBgU0Pr/sinlAOPES4quAixES6qHkOL71mEg
5RZPhNOQ4bwgAEm88cjvBO6C4qYhQoe7YfobRdOikrK32Ukn19GpNgpcPYX3r+r0mmTLqJzFpQY+
20g1hoH4LV1ZaZwMGhxmEvgOnJr3JkwTGiU/GzmmVN80giiqlkXca3UAZI2Zlz1GI8UX8WygKNha
dqwT+gMtTJvc3ndCN/xJpZf63U9kBcwSzti3Gqa7b5BQmdt8/JbwXp9C3MEAaJ4w01RCfmf+t3E4
ifRS7MpuXGvLyn6vDR2yeoJYWWA/vgiMZENQZBTut5c9PLs4fLH+DQTyvZmpVkeLTz5jLEi/lGRN
WweS2PrXnboVK2fieY3ssCMBsmCiWMgzR+lZLBrHZ3YtlGQQyll1szSB9K1bXNbq3XweFqDI3fG4
vfb9q+a84jOMMuWV+z9O1zi+YHDOVeALayzT07hXBLodwlQeSXHmEczU9g7OLjKBH65DpExmXvSA
mw/e9qH04POMWd68qQBKOVw7chbPCnS/XDz7QIElwjdQwYRDh2i6mDhTtdRy+zejepHYt9SUm1A+
YuNc4XgCHpevQWgrDfnjUQvvbpbMVJNollGyXUz56oxJv8bRTDacVDRlopqCdSTTkl11hvifwRtX
8qw3+SFdk9NUtZiDSxot52M0l1e/qXrGTV1q72wpnI+BZFi0FW1oYiDaDFrn5CF0IrpTq7R4MCNT
n5u2Ty4GRGrdeGh6m+eCvaYgQtqe3CIDR5rljnYbnEmkCse5lqKVU7LDY9PGAtKJhOTQXw/YfK6N
VZYV9ZcIuJ8OvIYOR2mlYz033lfceJk5CgFgCasZFxeQwrfuJiA72j+Zu0JT39C+2boqrLAtdIFe
kOUp20bMl1kiV1D66dfw9XriOBz5+cX4IiErFFSz/U5ke6vorB2ui7/8oc8PnD3iEuLbI9QeAfxF
mFjBqk94C1xFqy9ZEUd7AgTVroZA6YltMfEmzXeiJ6H7mMMb6qU3m3Lf3I3wCQUdWDT6A9DBV/qJ
uWlOcOqsmdH+d02ikMp08YNbiZU26+9CKJRnDDcm/G4iv3caK2cFgyQnVtezvDQ+4XuOEgw20BbQ
uYzQoa8lMBGMSuknyadD12CIl/yUigqNH7u1HSQnd3++bbrdATMA2gLni2Z6jcSJEPhcxp6ki1u5
I1sHy07CuEsNIwYIwFY9uVUl46TXctU+hrYIJ/JIoLqhXhXshxQUuL/qspky/cAXfSlNtR7IJeTz
awi6o32k58DPLiw3Ht3VWeGOP12XwQY/y48xTjQo7tpKz42xhmIGA50BmjtetuUugLMv2y9A2PRc
idVhXJQ2+qDj34OKVqK3JEv0hmsJjPqkAFX6ZfFo6+HLUNWEsTIHjN2/P2UjCzYEinl4eFd1dtgm
YIqEcr6OVQXAkkRCXgQTf8+ol5+gKsCOOOSaaK4VqBle1X7AwwC83fcRb3QvSjMSqC64MmlFrA3r
ne6GWMAMx9tOzEteRf8LrIPsZcaH9B4GcvUdK4X3OoqGGuCKV+B+m5m0yDbYbnMJIQxNnc514BU+
URu7Sccz+hhXixlHF68P/8kESJVP637UXW/Voqzzfjk3oEWTGqcwMcB0BLcvMkq4XNkjPHlT8sQN
nBtRwGqRYfdc9YegInS6f7CvZ3cX2i50ula4QSEciGczN4R4YYzxgxsiQDSUI+Iyf8r3hRynrbov
BPsBhPvSUaOqoVb15l07SzpoX4Gn9rz2HGB1lestjLljTgx7JaUOteI+s0YCQez8YyFDtMOXj8w4
OEMKIA8brCstJSCQbtecRpk712pwoXvUX1v6IUZMeAWsuOYNhwYO/6T+EobwhKr3ion40+qNY7uh
beu3hRbcaNl1WMJsUeT9OTMAT4tD1esFWdCJ1fSDmaUpVy+Hur9B2ORxHj5HVYryeSF8EKg6NKjK
5zkiXvbAr+6v0oKFdJENhr2rMqBtG6KLVsBoIOpw4EZJt/xIKV1nrn/Fv8rf2NerjwCccLbOgQYt
e1jT/ynmlKtdXupcAtlDHpOS3zGNhbBYjm4l+6jlX+/m96YhK9IlIc+PUkn/POU+Z8Op3ezLymWB
GkEANs6hnMMmMfF6B8l435CeMg1PlDnaWd7rNvJWuE03v6BHsts5OqukrCLyzjOlwOivGm4PDEhE
dK+0O+CgCmynMoUtI1/aZMsm5fBFay0F8LUHpn+xM9mQpmWaFlOuETJ1QLwG26J4jnFNJSjXFY7l
BJ72Ee3bmXg1wboHEMalQ7Bs4n+c/zbMMnuTNl5IbctDS0zcSgYQjvm543gGMJBqeJo3Hn13zFPC
NZm+y5fSQNqoHI4BWRHRrnHLEOU59Upwu/z1cijNGjmqlVNn1HlvB748HLEB/VYI0W7zgBqBgKbD
l8NcAZUALYHmgc0xNNxF0SOkGUS2b4E34o6NJI1CgI68H6LnWgAEn5BFERxu16fiFuDPkm77MoEt
+An44SyOSyevhWtvip7+1MsjYhIR0+Pd2+kBWZ+NJ/xnYOYwDDkskh/6aOeeBbUkLFEggVwaz04V
ANQSiiZ80cB2DNePBRlyFFgXT6f8q7z2FjB78Bp0ecwafoOF/kaI0jXLp7Awp4qSE5zI4cev3mkp
S23ry03IAi4/Xy78MTB1/sqYXiO4OFJ7O7GKXwZ1Dmc1M8yRBXGWxmcQLmboIgga7KxfY+KZRs7E
k3hfE81MPbsuwn3jhaI4oNVzkTH9btpwx5ddb3Zy8ZpfxC0x7keOJSFlUh/OVyRUx9B8sTKWuPJO
a8L4zrhE2tKx7FG/a5X3aqhnzaI4SfamzxSuf/6kvlvt1kjTn8fVI63QXkc+CSsFAAGC547gbn+g
NeVbo94CGIboudqwW5itW+biQxjV8sGICrjVKpPZXxv2rykamURLso/k0w4ZimYwmCdF14jHnZQz
vCj/tYSR2xuK7cE0ljl8g6fQQSHFeR1BuAD05iVyz1Epgliafv3aUgIHk+1N3EddFQBBqaOsEFaQ
hb8GvwnOe/S1T6rqlo/ZWMs5kHNaML89lhlUEyblabIxGgfNwLEaEi8wczOH4awWiZdaPqciWTFi
StIM5oPQ2ek/FLgIS8svMlrJQXcNmcu9tfsHHffopdmTX1Me/NwLPbCJbbgboBhzMb2tYuj6Jr32
ucELv0v39u7FKsUOqfFtvvikdILA30YcHlAgKGGCF2KIDwLqNoomd028OcUA+jlSQA0Njin6/YZq
aCS6g9IQRnB5pxWw8xrrIlySEFS5Ka66RmZj+cMCOyR2G4Ao7U1jAk42b4hyfRcQT057wJmg8E0w
OLqVufPGwF0FpgEwUoPhBgRyvUV37/fvJIo/f7NOGeGLY7xLiuLSX/7uXTdUm1rd20DwKYKtCYq3
XLvw4Ntq36AcX5rliMUmBTC9ss+aQcHM2qYFdxLN8RAaDaEGyume1UjR+7mUJe0L9QH7TYzTdCtX
KXGzptiWmfKzhKM8HFdnPSVS49L2acSYmve4jbN+n2F5LsSd/hF91Cv4wNSkFUbkj6niMStij/5A
WqXJ8Ue0DNI3txq5mzjFv9Go1vX8piZUMMIXsTqjzgyFlU3i5jYXEOAZJsaRDHhuSZ0JBc6Gw/Gv
2fTC9aXi+zOEaLBvdr9VOoxHsxLiaOBIcV2pr5AfvncRww5gHVaWt8kQn0JR9DEHf0LNqJIMb/AT
215hgnoDQyJvMD/ftgyywvFIH31PQij1Fh82GmczEekmRtX7647QwsFAYTdnIlt/RLBorExkfhgF
kXPzi50c6Npbxx/bk0067dV+zz4aNI66LlTeN99hT644O8tRuVRfW/iQqMcWvPOzKuYcn2t1O5wF
PGS/MRasILoW8f5ysxyEHZs6n2c8QpwKW9BIr5L7PQh0DU09rLF9y+zX/6CSQNAq11BEMnxaG/Q9
/1BKUweLBEAJuSaAiY64BK1rIwmcLkk59ClVvxxxopLEE6RqqadP5RfYd5mNhg923oSCgtStlAky
ozS8V+l9aVBX9C4UUR4hSDLSCYsZaGYK2JlZL5tqkC/BE1t1WLQMDkJYw1sYSsiQebl8Poiz18t0
D0fIuKpeppg4ZTEoSmgAsYIH03k3SGw1OIqmIabucZAp/mTY1ipDoX+e6VmYVdhRyraWPcTSqbLk
+9Mm21c4tyy3N9Z0PGrqEj9dJi/fX/OozI5BQ4vtMc1Ercrps5bZtM6qfM7pnfjoCS65xdjRU7Xu
ec3GD81V6QI70LnNRXoj5pt5p1z6/HBzUq6E1TxFzfMtQuBd4dn78KS8BU8ZEfbIfpXx6t0/WoTI
wxdOqBU4EaiuVkiZ07LD54CLdmMsxMqqasXqAoGpbJy6ZbxchmKZnIs4CMb2ZZVWCieScOnt6Zmm
i6iCmoUdFZdYX/3cyjFWGArA8mUZWSbuM9ZxZ6gBDtQ+mMI85PXGpcBKMfXfZW6f2Pc9uo0eqrMt
b94pw0t2v9ZPdQ0O0RBPSFDYOFcLlx/gfqelzIu4r42JoPzppQ8b0S30EYvoSsw/tdP0RoHgZKUw
C4tLwA3qa5jrKxjpoXE1vwid+a26DE9n6Se71rTgIe3LDkFcUx6RzIajo/66vJJyxmw11H5ole6D
g0jfy6skkJBRuWFbGHTgvmVgTtWPPQon1vfJakGHW+6kBO49vl5z6xIAtEkos3JHbMkESWdQlpeV
geM2+nI1v6i+wSl504OTVWs3NIVy9IXUzJ0Wia8Mau+G42abgeEhViWqTAz4gedmdQ96KeG+QvVh
a3qI0dCW6hdFzpjs4I0vz0dGWutfxfSP1lbu+7tNW8HYkRt4nGLszgO1HX7iTdLXVp+sQ7H8WNmx
NxQ7JqA0K6YwVUUNj49FNeLa0lgNEQTAiCwXxD1NRsTMm10haLnXfO+qwf6ehuaAlHnDxNmZM7Hv
wX4gPRhF786MD/1M40SMWyhPoomDAKPhG8sI1/vNwhXfVs68q1YA0nKRXI24wvZMHU9AIxoVyvpm
ZI8lpQbgG/p5dlSy/fOcgXujTN2g0ih0fhQuuE+L7xBL2h7cFEZdeFG0uUnQDcUZlTEOssF+h5lZ
GGceFkqG55IGuRL4DYZpjTBb1fRhdgCX4c9I8UC9YP1InmD7tVGjwv1M+NeDJFuFYWdSSWE9Ccss
d8eGOZCtLgLrZInGMFBWPrbKBLaFwGrImXeL7WOPofOhgDN5UCo1lGhgE05Y/caomrY9OQzBjPiG
UOW8CxUwGfEfJGuUQ0xPJWRpdGPw2CgLdL1Q/RXuyj2VOjLP0W9UMgEygOu32A+MxcVIuCr2lpJm
T4NPKEOMb4Ab0yrAUXRMvJYjwinMcqA/MiWykdZlZTGE/4aru9A6G7HByh09HrX1/xXLjAlA6BEl
mQimocARw0ylM0PZodGO+OfT+/se8aXho55C7GHe1XqwO8jFzhm03zqXyh8eOeE3/IYQ+Fv4l2xT
47LbS4hwD8LjyzuIFKdR+tnyJqsY5edUGAuABRrN04OBp6SrlIuOKE8d+4fwe7OIgjFS1Nx9QRUZ
Tm+iZh6lNV1mk1Dr51lo9OPV9IihaBWBdjq9/t3haP3eVdDz0FbzEQHr+YF5fWmce8K0Nd+Heee7
Fv5q9nN5jKWSiqQI0PHlL2lrr/W/eEzyi0F2Z4JWEaEyO/Nx/X9pQJMs8akPDpJQ68nVkS6ZbfSA
TtValRVoAaXjwOcyxD3ytjMTtqQCIJ4iV/9Z+2rIswTboiPB4o0hNr7nffCMGDADM6CkoHx1CLmW
O5C2/OyTqFM8fuo05WpoM8Ms7nQQDZOaqfo5ux+2e8e4xIvBroi3ngC8Sit7G84o56R8kWWyDDA6
Ln/lveTrjnTekVz1PIMeI6ZLhyxIQhGywrSBj5oC+IXcPXyuyrHa0CfJe2hw1RKbRS4NoYcgaUMk
UILQGRQCgPW7T4vL6gwqu8xgneTUX8kIVio9WvjbnlaLhcC6+AhGPFEk555dgalrQeNp6hsB6xco
DrZY9NkIAlsOLcp14ZgKtJc9j89AN6PbzPknvzRCLeMqYt5w4O/2Z1dKgpBSrwGv++p8eyycvbyR
DpVWoXzoFHlUZS6LWitKY1BzyPPTTRo2+4sXGalg05u9KfZciA+pfpTlFQF20NWLa1hAzt/CwuBW
FxW1QUhH4YPuwLhHqIos3sQYEgrNEYz6cxPxJPNl3WkNZpDLc+v+YijInrQaVBTNp0OBF4gdPFlx
bnDLXwCXFJaeFshn2kIVTtyjl00/ktFbKxnJV1aNMhV0+AjeNrUgz9q1gd8XUfLPJpC2lZrApwHx
zzh1csIpIVWyKt8knDML00x2EJqzPiexn5ROasaCm/3ttJsRwk6CNe1Mi35PbtVyYKCmT+Wo+x3d
/+XAqDEGUme9R21W1++ON/h526PLjjlTUqJVKh+VQyHv0ya4sB32+c8/5XIuZpB7h27eTyITUZPo
dq0YrE3bsKaHUX/dXH9P1QS5Hx6P054XV63uWJHtHeh02bY7Y/IuePtQwNKpaO/11+8jiihCFhPn
jASt+BjfJSGjz1HmDXOzkLbjIbajySa/9ulBO34bUQFc3yRYXVhlypU2XQI0zOep617Fj3f2F81t
+AX8wzLJkt1+LTmoQSJ8JRlmKCAwv4Eg6BY73H4wTDtw+ctU9FpzzU1kLlPC3pk5uKeAupQb8BjH
r/l0Tt1zw6Wi8vTq4U1F2Iqu+K8FGlgLHEaq9scStHIOOkO+SeD/C5aauEebzvymeAuDYXgVfX2T
JU16iPjftL9Jr5vKVQ3XKC5AxAysfhWbCYMmWBXy92BFhvh833NKr3JHNz5jZ+wurhyvfw7a+Z3W
hJ12XE+fTuPfGIAqbLt0f5E9vpiEKQKaXkjiFJhipKcXoV+1opxEF9QZsfcTt8MCapjjB58Ic+QJ
C5iS/peqU8+hHA5Pik+VXU8HABLc4A7B0QbC/M5LEMFfrnHX6b+BSVoznuvcIbeQXE6WwoFNBI2U
F8nVasn0Ko72B/gDGo4HJxu0zA2x+qV+vqTq4H4ZhsJxpjbg9hk2vk8rrprDObUViG2kS+0KOcZ2
BlxVQ+PGhHmLy7GJuStDdX3rlNcgAITdma0VX3b1R9dhYhZQ3KARXmASL4BpY59Sr0saUqM1sb18
ixZkYZRXVB97aV9XNfCybDlFSw6opoHJVAV7t/rJ6zbn4UDNmqTwlChCGBIsx7aUOPa2Ed1Px1f9
5oY14JQNKkbzNOoWwGsb9m+ONhYaiiMwgolxxXwtjX1zvaL5ueBWJsDDtv+VuisxhWJPhyOuRBLJ
YhTp2r0dnrdPcOO77ii8vFmwDqbs+Lw1nPTEMRWCmth8MqQSLqbAXwTvedeStiydJVH8mzoEDYMr
d0Ytj2KWKXdV3XLdKMrYK9/MT9xB9XO6GXouPvO/V126h3QNB+79WFFBVIQQpxEmICNE/+kCSYO+
3fbUAJ6Ai5Sgz/by3n6jXllRhIscfVUo34OyMrtByhhB0LKP50Ai2yDB6eWgeKQsgUfUNOvDxPoJ
P0Y8a2SmIoawE1XgDuDoarD0ERc6Psrbus9WmVvGPKeYeyUljcXkNJMPpNda5JD8/jbRzJIN2QH4
xLOWtpcvEgm93VBeAFSyWefQ4nN6pYc5t+Mwk2l+0RNyqiUJloiCTwUlkxQBWAQxdgK5dPfuCjoi
+lOSKFWf2tDCejAJ2xrGoX8KaPRE2ZikvXulTyfSv0F8G/L8Bkc0dNOoV1KV73O1pDwRJXmPE4k3
+PO/77mA5pIsVD1eyzJRTth67hdyniKSO+zI62wrXl0ifhwAzO/lMR3unUpM9g5Utpr+woYKx6Wz
u3mUHuPmJUfNLMP0n5xtNQ6nsNxMv+UMAmON7tJ+CbXBqP7B4k0z1aIspw6SXmsN82WAOrNJyiXM
f5aHYvehgJSLujvYrWQ6tkCCiz4Oaz+TgfckFx0+Vz10fZyLQ1xw4DgMD6tg/hbzQ84ym6KdZ22O
E8Let6smkvVHC2f+jFDQUALmC+MTfbw3NVvKJeYsUHRhfA3pd3fiQvvRkfGvM3NBDqePB0f1ut5G
kGfQ78y0X7JdLOZfzTDPRLRMmgD+IB9Cs1MTOguWWPO2/clOzNgVGsTl2Lhdn/bvguhNWPYKA/Cd
vEk9sbB11UXKKYzjglnxwS2TeMDSts8Kz1Pn8rIAUvywOAtmFir6yNSjgpgVir6oBD/rOzYzwiV5
2oVBxjNoogYCSydEqDgB+KtjOqLgx8ibkac4Y3dddkb3Jy3QQPf7RJAJw2UEI+pL1+stq1X365Gd
iZqc5oX7HnCaanB7D38X8BFnUHyiBtCMeGfkWze9MryxiPw7BYmkyE5Appaiz7WYUX92ykVqmUz7
go4qGKUqUAFzzu58Odo1wK6gnuAGXyjwtnuwEuz0vftOCOp87QNdAzoFmIWET3lTWThof5OyYz9p
nG9Dfa2xrY/QZLr0VQ31x2CjqQ3tdRypAxvWeB+q9gU2W7emwlq1fnXYf3pEizPVV75dLoJSapvJ
1HbRMQCPqw4bn1dd7Oy0FfPmlYt9ShR7QJY6jJBS7nd9CSvb1ftL7xaZc4+Ag3bMsnwvT8fMRnDH
7sqdf5CaTJDYhM4Dc+G/5mXyScQzJbOC9oSBGMSOKZ8gg1ovWyVZO2j4sOupOgbVF3/N7a3s4z9C
MsGiRMbHjtCscLWmzpM4A6s2A3k7JgHTj2gt3n79UVfT3FpnxDCn93F/k+B3l6C+OEBRQFawu0jf
9m3goAbfbl7xHWkwUqvIAdAhYvO+ygcvmQam8zjAQL7HQtiYIalk+glZIUIKc0hnj/qo3LbZ3Tjw
4M5XEm/UiTyAoMBkAY9Scfbl7zb3DlN7L3apG8S4BoOMdVwDWZlToYQpLsj/79HlrCdrHs7oh0TN
pSyL/xDPFBZVdO6yiqFpEZaAZMJ932BBEH4g4TWguhHIA3Z+se1Hdf+eR3PiFsIWxKoOCzkzPk59
7h9ntf/ublMQBaCo4BdYd5954EwJcjaARvNHsvcMx4EXQRCeMdY4Jv84f/S7pfmdmjdQDxWDRhSZ
yDo5VdQHV7LZ6Y92N98Ifvf3enLC/Z9TVdMOOAoe3sa2EiR73u2C9DOWRbyF1LKl1R1D2iRJNfdB
op6QHFr8gL8WYEM0nTPxcHzTXWFEnBlAXumqtODSN8jYi/HngnLOve6yakKM+ThmpzyWxgzoVW/X
lWfvWIR2ucSEYGfoyRb6cX9V6iRZeKZ1WmjneN9dgICfMr9EzrlBTBq6gyKHLFm8Wq42q3fRrva0
XJBsTxge8sK5BJUVXgQMGIg2VRF5k48vyoZfKgP49DZn9sdQJRS6nQIzlOx2U4i/L0MqTcuVpzx8
V3puXXDiQAe6Mlvadz4X6/yWzk32CcY5T6pBg8JWo+m5Pv2jDgaguuWNOg6EnqPDJrt0uUWuekCu
cNCiGIB4xc/afwRZjmbdB3X4BbM9m3aEvNwkkkYt3bV8TYTQuSUbMVsfiOf6bUMHwbSO5nAo9iTj
Fw0cQwhdsxR3KZ8IaMJ9gH5WgUQV+yksHnKrG/jd+fmw2tkw5Tes0g3HdkBrU+ONHChdW+2Iq2CK
9dAVEbuP0oCc5s5AwG++1YYxoIuCNe3C6sRA69yGK2wjsMJvoXgv+dyTksEYHW3riLBJzaPnFNwV
OP+y67yf48VcP0UsdUHm5EaKWumdK2UevmVLrNsFdezuSChKgbabeQRhHHc3+iD2ru5uPkSe4doU
6Q//7STAtZLML+NrRRGoj1MLRS9f50Ck6RB1H+l4jOo46E8tfJcQiCHfmAzR0wGBa66wX/5Frs9v
RVdVhYK7e5iqvlzzHTnIPWaYQXx55Jeed1Y86ZX8mqufD2D2P9jVz2XpBA8aSueJhbiwuThv+x0W
z9Rw03Enda9gJyZ/Lmq53mMMZ6XJ6bFlNHEwX4BaGH4U2v0omJ6xJs64LcMHZZiSAYUs5hoG1trk
H9gyfw7+xBNe4Hijk8l1NUko1PMmU54lMGf/lBmThrtLHrluFKQFk46Pvo6r6Xzl5awFg7rQF2Et
mNEYNvWrZobi+kYfSoouGCP45Zw7lQW1sKlruq9k+pzPqaGr84hS+5jsmT54cVL4jL9KVGPemLyx
n8v53S2eoXv1cD2oosHV5wioCrWiZz4vXceRL3wzwr5K3ZQkIsjbYbYQgZa3lS7fV6urxMQPhXok
v6MPOW+7/9mFPRdYxaUx3cEHekEKN7oDQQvOfCGvIOM8JjUq4WAHgKUErDBayoxw/v6Ia+Nwoc6S
f3lpBG2aUlDegXMoqCEBBPM7eWSmLffWl94A8R5WjYxcSr7sw5XYR8/K2pqONEoKbTyQ7yspA1UB
eICvHVRAyBtqjDG0SxPQi3x51JQ1P94YM/USPMYhX5Hxkls0AbKRguiXK0WnBkgUhB9DHbv8aF5i
lE3wt/aKr6QhCMK0qaeeHvDPrvLCQXyyw415RTSb8AIu/3fgKnoyksqiJGGRjNRGY2+qPeRIpy9b
i904Hlul5LGGl8sXmQe9xapfXqKqCGFU21l7v3Bti1k3SM2WCPE5YFBUemWn5nr+xv5G2iKON3sm
anxtLAHWWXPcXvlWrw9F9M6bl+4J8K72vMHBrFDRhYjjZzkpOaE2BcsRHzrQwVaMF0yT+X+JB547
DzP95bBvOxyFy0B7wnjvUVJkawWTTVU1QrFo/gMfVgZxueLluxn0ynLfza86q5sZx811oAOR6YdL
WLJHdM+9cNHWyyhjNaFxgNkikLLquGABpe/yqetAEedaNZAIHUdl+o+F06+9fQvB3ufuRoRRSD9f
SKYQCw3io2bH6VYmspa8bdRwUTi/M5Md/+9roQPnPVEc6oLxAf84Dj7eoxFbgyWoOCBd3L4/D5ds
IOBzKNP/IN3TZLd5fFn06FJcjmJ1KHCH1Eb5Kx0yBdy111zin4ZX7MzVRxei6etkI3mAuKJdq0Q+
sUgh7R2d7ijWdYF5h7ec82qr5/R3MhdkDiCka4jG7yeapa9ifBf2xcrtcEPzV1M4Zt+CsDH+jJyQ
pZVdwkoy0jkR66znuNnosw+k3EN7WwDkRQU4ULckAxxY+8ATdoBh2pt5MH/IhECYAAefm2k83WIR
wD7fg9SsUA4BgRlfie05Mch2wqScA2JUaJwFaNxd9wtkRP+zD7fBcMRbF+xAyA+E3L6P322Ii7pU
9YaQZlNUs6V7fBVglf9qLdIL8qXociDuEAZdSZ+T+9Sd7PSz8odRyldAjprmd6Eff9SITdmEig76
zL9wquhgJ+G9xDdxhWSUorWNWL0GBZHkqVakAOkbUO4KJTCzCVa0LF5XX1Nlx5SYh0kstKIvFySe
cavpHSYhksC7Nz3nouF5oiJmV6IyPXZGOGQ+yMl2YpY6VPUqpuDsY90ldTb2eLDeAkSvOmR7XF/l
ZhodysMnY3uTBzlgZL+ghv+cF7IneFNsqYQ696qOECVvEfq03MXAZoEbQJ/2ZHYP9qUAG4xRvavD
0ryuaLIloX+bZ3G+KvGSCQOLsATA0zvjRqiugu/DbLpLmA9CLcYp3GM2saT7toxQIFMXr3yZNRgp
W8f95RdS/CR+6ApRA2jEqDfJDW3bQxgTD0ZcveGtERWVCCUIbrXz5ZL+LIVjBjL6rDdWbWIrX25B
+L9T2WFb+reLZt8Pr3c/Hx7kAEPfaAA2xIr+/A0s+pNWveZibN35pREggl936en6ngoAuSKWfSBk
MUEcrtazXkzv588JAQ9ahaL0FewR5D0bJPQjcJ7x9LB9iRGeEzIt6xlqkPnj5w3Nx8nafOyxSBAU
oE3cWLoSsh++88YURXeTTrdPMAaVE4vyWvNGAgd48fpvMCmThLhnnQwJTOX/WUVgD438kpUr33ib
IFSAGMwyTG+svBBMORCb2AfqtHgIQliDsFv7BXHauAFK/JdFKBvXteQ1HmiouHfCWeNRZ1mUKGzo
RpRVBODDO6kVQtVskWyjFzLm5tZr+oFYkjokBX5p00FdvbcdvmZhGScwMTzWZ+hCdaLkmVqQIYbg
xe3ApT9RjB0aS7JCHAEdxZs/56qdesWaKBvFwVp9f1IvTlQQ45xS3oRTbrxjEPY078gLdfJE2Bgg
dC6mxzp+1TDBYW6jr9/7z+Gfede5itVaB8N1YSambLS+Cq+idXajSOefxZaYUwvE941Fl5X3oM8V
udBg03ke6od7gt14Hlwwppl6YS4jQkZXpwvsdxwRFJdaybBkIIMNOqgRqSYb34/T/YREusJ5sCBE
lyI2fLJ2aMzGIQYGvACaK1/XHoSgJYPDcFi4Lq2K7abN+0ga3HrWFLNCDArUxfvuuGos0DImL1HO
oO5WnoctnhzxoFwbMfP6GvthyYAQbH+yniHzk8g3xpL7NEyf3mlz06KlLxPg/R/LFn/XbgbTbvaK
7gJWXl6ViX3CPUpImfLYwff7fwznmKzC0sLQqWrTeBPnzfXL6dlDEhnuG9msnfGAB6AoZxQE/bPq
4MwT/b4oqWHxvqt/0Z9M7AuGP2OCBkKoqyY79GSNQzFJyOiwYKr7x4AFa5OmB5frF/q/8y/c4cFR
mX0eOV6/Z+bTh69BY3Uv2VRDkPDUlXybYvfZmJFJn9otdlI6guioFuHSxtA5Fq3y5s9hMFirLytP
IOaIIQ8yRy9FhPj875bhpZCYfhh95kwAFpHNH5joU3szObFsZw0ZDDWOBqhWjuMP3l5Sw7qlCIyt
XIivsJ4CXn/f94LmbN8sHTTdlBlW/GAl7BI+vpI41jnuQ52aP5s81eOdc8VjouNMND+2wUA3OGow
SaLzqpFuyoVvmy3OEIVRN1qri6TO8UoauBgpy3EIcYt0m6SzXX8XkAgOKnAnWX/hh3vUWrnPghaC
VCBGPrXaJ2+IVwRJYlVboAnLVwdUbMYEalBArIeay/jnleDxjdkEDUNaXc267mFY7Uos3YqqvNul
/HqSD//Vk/pHQ8853Xj2VXqLZODfYytyObPRX9RcLyO5voI0jvg+qmSwShfr8RF8yNDx3m09Jk1G
NWk1qxUNTRX4fvMEuLsNq0Rtebf3aFUk0sd9LACCKnSBOHGNi7b6oUVMy3klKbaCEFHWrUPC8XYo
JSCAqkxCEHS3h5hjdZ7AwGHUnW758Si9166Ydo3EO0pFoTgSN5if9AEwzsUWJ1qbxuZVXzQoSDKQ
wSk6Dsa3p2ZCpwVdxNSO5lSdxWy/wZmblLJpzZIewCfMNGjzzkXjMo0YNXXZbw7NHVg+DAFny+mh
uj6VIx4z1vOr3yOM0qIVT/u0Kf+X3CId4HSE4ZRqjoz+5+dRiWZXy9VjjGdLznQ7zynAg7SXP64l
UzaJ8Nlqiq32zP94McF+HhDobeQ6KDGYJ52lw0P6g1KZIl9s+ZysPBaUYAJI+WMIH00c0yfB+/lU
PiUV1Ra6yGE7CPOS1dF7K1JfYpzGRNmwzEUDwYxqNw1CR7qgVZTSAreMy4q+VpaOJwJh7Pkueu3z
kOpyk4pG3//2UqN7zt6Tza87udrUaW1iQSCjTLokoOAwcsKLhtLyXhU2RZoOvpH1ZvvsjqkRnuA/
hPN82ZpA1rIv49hl4hodj/WUCfw520BLvvnSmhk5lnGmwL/HLu0j2qub/VEzpiWY7II5FPJDidla
2XOTuhZ5KQmMGsPEQ6g4QJ7tGX8Mtcq9u03lLFuU12Kkp6ZVLHRxqXHBfZ1AWNtnaN2wexdnjluA
X0w5IfmFBJNA0PcCT0TSdVDFodVcJ+Ety13W2WZn5SlACtKNZZJLGq67walJH7Ay1u5cOEhXk818
9Uo99AD9ph2K9xKnTm446lmdZc9XZIH1dW3udN5cRUbx3M8LZW8g38BKOeYGJP6Uyd6CVVJAlrr3
WVgqiqjporb3cAldE86D0xDjepzFqzD1gjAFwXvoFmKPsg0uqB/s2OJNo7PsMTkuP6Q5G2vEcRGd
CFv8DVo+XQZ5tNFpQ+AyDYPWDFIQ5JiYzsLYGsX6FWPTMxKW1aXzhN45fSfaaEDOXhGMrWcYonUV
G1UDH+9kA7eb7HwlpXwBLaas/GF9XiVw2nES9vwmDXpkLGi8lwYTty51MybLX+Gpg+gGwPhIC5d7
FSYqqJkpRVgKMmEWUwbsXjtQK2TX0J5Ex0jxuETY1V4d4+DJncq7hT0r56aeWAj0oklgvTHVXY/y
j7aqc0f2wou247uUdpShbDvQRFHFH+sGRwwh10/R8qWst/b6aqyNS4CmYogZRMHeA7nu8PcTm9Xd
lNOafr0XF0MTEJy2enQkrXzOBG7yJSAgRsR9q6ySLh5rs+7SRJeYXHiUKMsniish2ci+z0xP5OJe
kcVtyo9tKh02gOi+nu3j/yFs6b6nGd1Cm/Mm6+ZRKISatCJPuHnLRGs4+4OXWmQBGn4xRuNlc7fp
lgeYFEq6ouh+QY8HA+bHndaRp0uRX2lEC7velEekkBrCvrYRPyTIaGodhZLLvQsbM8mETr3VZJ4r
pzjjzzSwek7IiNT0I4yiBf6MaQKltG5FYh7vFo7GjxOupeEXmvbkn1RPzcz1eGMS+PnpzL5yJO+S
qMDW7/HLGhsC/tXcP+vkCr2Hj7xLCv7RQufUEPpL5Nr9xAIGEV0McdLwsMrhCmMsOa2QzBf+5tmV
oKN+iUwH+12FFEJzUY7Zw5l74I2uVvC0BKWss5RFkFOwpZ6gUiBe1pYZO+fc1mx+eZ4+6oNK0lqW
ggC7hcNF7Z1/DXTjfBgcOyFqTkpqCnBjOXB79spxPheMWe3sjsGF5RH2RVlUHG0QlXHKiqxCK3bX
OdB5DNMKJBYa6uitvDnc0w++4VHg9MOwindAiVrDg8BNcRtwe8SsT3wH7symkuE4dKw5p5T6k1Hy
D8gqx2wvnPcBwNaT1G+HMriM2N0LbxVPOeHDOv71JKzEKYV24eg4YQKn5GRhPLMNB22DbvpLhNnt
GLDEB/10xPvHpmta6vLOlBcpvtlMLTGXkjP4IYaPWuBEk/f2QKWm74SFBnDF1hxXivfMGP7Mvq1L
+DCue0qnK0OCYze9H36SXY80HPBeSkLDoyOo0qTPVZ0FMxCyWJyyF9dGFXfg14Ayhq39TAICMogh
m/qxCkt3S5T0zr881xXoacNRaTGbHsLdwF7y5zlzsMt+VipTrNbTwy1YKoKOUMSIthe+nF1Xapr2
4dReNYST9dsumMNk1jbOyBLefMxqxCNVlX6Un55/fYeeBvfkNsHzU4wJ+BgtlG/jyrjuI+rMFcjV
nkqGxPdx4JfLT9qmCIiescYhZi3JHqyhZnCQUPCMhTO+n//+YweUP30d7uWWaB+nzgIuxXh7qwQH
A+A5pY0GCpPOOMJstOH6mnW8MIgqisQquKUbUK/jkV9sttx4omll+rNCKqlphC439SRFtUtyNDdq
audOAoOq6f7EDbf/3qDTszk2jnddpuv7gBL+w3CavqjFdAz1+W9WqoXkom3YJuUKNXBTKmRP8EQw
IQLnBXMcDbM4k2hVUKC3MDyUD4lwTkCF8SaQI7H3M9S8Grl4Hqxcjl4/S4fatM3pS8qlS/0IKr6I
0O2OckBWr2j+EvfgIXj3s9sNnWavQULPjz4btIuOu3+X/iTPjvr8LVHBDvNrzQJsjQZ+g08AE804
FjGTERN6v8haRrV3P3fk6oJo20lBrstQBRTBSBTmTTypygiisZtblk0WEu3lqOgJ0t0dlYA2vw9+
uSc8EYwPO7wL9Lmt4xrtwFwezByceHbEg/E87pTve9GgVEIWkXos3Uob7KYIWOKNHFQI3sjOmMU3
lPcfg3Te00eNRl8kFwD3SNy7iDJY496Gnz3lwPUApoHuXLuYpgZh4bbuz+xve6RwGKouqPAWUzRy
gwInqBBqpxZyMBIXD49bi2DgaagSwvXMiJ/TSemR/5iwkzMC7tG7s1dbp5BUJjBL8eerZ/+nkOFI
KazTq4R7EYkwOPTqPupuWwovu/k3QLz+0YSlyrvVodBmpgB15okPR0lL1TzTnvob6lkUdCswyO7e
27/jdQlfyZ9Aqs7oWyFh1sTYgrgDyMIAIu5F4BQlqLTRcW6IFWryWFIh7YJRfjumMf+eelFZsn6H
QiH/f4Sinv1MUvOt4aEdYYdK6YNc0aT2KXT2zOdupAZoNRsWtkf+dFKbHJwgtK3JQpiYRnrFgmEx
OlAX+X/u+1oASHudXRSjpXK7ODUgQh8zNLE3FYT3Y0gLZh5YvGg3eHjXLUiU4rEpKLecyMx/YbCa
7P5zvK0CFhUloExnPzgs8ZZ6G9YNOtwQwTcC7aGsbbjUJTAJZLyEc3D5LaTEAt0d9Oxj8P9EYgfa
hYFMMPM6pAdUjrHkdZEAuqxbBRaidf++E5VHEOBBmeHG9eIJ32RPhOox80pIs8wmdXFW7faZnk/d
LpeBanQDkFuXG2HZhsne7d2zVBikXQMfkcDHO/5W7LtcWEgeB5bh9qilwmwBH73GOEVbLEVBm9Sc
JjCd9aBuXnt28l+ShDMtu5SgDgcj5T6NV4LK7YZobPOE7e3SK3nW1Y6JLs1y0ZrAT9YmYOjoL75d
PDQIFuC3t0vbf/WUwi1f8WqRfXSdUQRBv7eto3OEsfxgd8zbC3iiTvzkZZXLJp3xrambOY5pJO9G
j5Swadh9+4ufYc0UPM313u6CWCRuez2e0NB+ATlusBkOz2T13PObU2B58wNf5ZD3gAty64rmjE8P
LgKIIHlxQnevZ2DxyhXcPE3jeXT6P5PY/eICVxxYHAUSD1dm/fqnWL3ZkX17LMrmr+uaLMpYyFSO
pS+yiS88dd1Fx+/JdlAK6ST+IVMWwUny70zLAz0wn96GzUWMpVqs3H2PR3DeGXacfW0xTvudGUCO
nl+1A9H/804aTeSxcZIYULCBLEm9GBGyF/QSJcMZ2RVXDwrLR/zWiFAVjkwzC/1fI2xAGQDdNmZa
HFdOdkHSmmURTbAjqM7okLjuCO6ufpMDvdiLumhvW7cQJi3bcFfkhkthchtPpv4nLTgdaqslIxXu
yYdODgBe7K5l2rxCcaBwN0pHCD30DGZcrc0O9OzqLSDtSb0pDERuCMF4lQJteRtY3z9E9mnc3Oap
OLy4VEB7bizmxFN38J+DX/wPkLynckqk89dzZdJqzu2fqc7ENmJ36u0LMwwK86AMrYTRJf4puI6c
IyZPNl4plv5OhAGPhZoxKXJFHrl6tyuNmQPglcodnGh8PjDakl3Rhowig/AJTDCxvymCI2MygPli
+IXlbBgAwC+SZshiIguBoCZU5gSfqLKnfBFVIDmPCS7R2NBSIIGAeBfQbPAW2AJSlAx+fyCOHCa3
1RoQVfxj8kgiaQJzxcPgntNMV6qyEK3DGVGrhuVwZuaYF46NDODMgnSfKeuN3J9tVPG2fFYGsFMO
mtdUyaGwOcaEolXcxLyftSqiJSXpuR+4nDUoHuFUnf1quvcevlTscPlSCE+3uzybncha8gbprX3t
3IfCUxzPo6kFOkiJrlOi1RRYebj0CgWSsR7zo+cSC/fUgBWxhk3BQrN0MYiJhfJ75zRSz3eSozGF
6iNJmkl/dMC+IpU25I8q3CvNRjE1zCR7c22oUMMrzB/iI4bGqFXuD9GwgIUYwhZ+/4w6AT5JalNo
Jnxq7joOLg9QCmn0Tzvo0ACUtq7JGopNZrM4fFQ0F+XWmj20K/vF1gO8oJ4CE3si94/SJVuTny1H
5TMhFjOs7NYP3XsM4uU5/W1Z8tc2BNBxEE3SnZ8ZCKEzFCF6yMzJAFSe/8oqad16m9P/Sp0D1VMV
CAACLlWb0IXV5702831uyTD8eCt8/kC47bCQ/lWNOWtdQ/oU4aESTIO0oIHtYboSJSX+IEuECmKa
IMdzfpmNYT8caFEFdR04OhGxWVwa6zu4z0Pvz8lwRsTxfcJJ5XJju+qVSQs8UwYHU48n7T5MQysL
dL3KVgExsRc1Zg9ZD+Q7bB5ium1NgnOmE+qzS++n5HZVj4lsWUuzD3rG90ZOxw/w+cxaFjS/E/L2
sH5SRSvCa3j/Gnk+cbdPkKOYRC82K1+onTyx2tGQFdkXKjEBMxowi6YEVaDgDgZE0WGMcCtLhJao
bDNudLRSRnUQ7f8e2Vn4DE9iLT4JrqWx+ffvjmExwbkNREOSMpGfEpTEsvxoP4gVdkGSnsZt6hqk
KF322S/YojIFWCPliPEnHYEJhl2yO/8Q6fu9TSHi+1pLoln/67lz7fixI+GlXY85XaI6ihYjQxi2
GnXpzlRVDUJ7l2nfCPQ4ETJQtzAZhbQU0ajlafwNnALJPBSHOEGvDKXWkpF/NGGBG7GE6VpShSPs
EhFlfZ/kMb2rhr5tJ7gimmg3CgsKYxj86X/sR91+Mdq6HB5ySDjbBgQxNqLsmW6vwIUksTgmyB9l
xd1PGS97YuYpkKupM2eW5d/RjpxhLIOz4GlO6iMBTGv9AtkaOTzGuncgScAht9sRw9ojTqTxzpey
wnxv8S0YM2zQXLGXaDRQE4Q/VGN3DOMOYiDTf9YQ6tixHRxICKogxs4d9QQ4DemfCJtWdgH+sDHD
wBVTV09aadYShhaTi01AUniS1VFRvc0bU6BtbjfnddGZOj0hT0Y26cjyss45aC/weyvcUA2YIMkN
50qMLFdDRqlokcMqjbcGx0A4+DXyfYtAeO+NpBIklg4pEoz7ernAemilzOHUieuIxl/dQl7aEhtI
pg0tD0yU9DdZJ1eQhsNxjguD/zENUWCkGZRgrsnJ1LynA+s94xXdHs5Zdu6Tsj9fWlpRUbqukRbl
rGs1c+YkxucLt8JQEUZggAXE7mSTm1ZH6bl+E/h+jLiEOxOP8z5XlbfmnC7b6un7v4/FGrGW/Z26
vEsE7E+kcEMer1f9AwmlZEzIcHogN8Gl+5YUzI8u1MZOOb/X3Z7vesE6iF/kkdD4omPkrS3xHNtP
nud2xYlwTwcVF6Fh+LXmeJ5shnl06wALQZ5tyRTvOOd1nYSKXjJUGPgtLoRybQUWslt+2HG3552X
yeg4uTTZMa2UBqX6YPqSCnIlGnn2XLy5iHOYvQAKVVosZAUqE7TF5cQQNYCBoUQ7Tjb8EbA5QnLb
doPk+hiHRZKSYYi7+I+G8IDtZIRBhesadbuuItpdKfF62G7TDONek7BtNtRlAdEbFJ4E3tMRAEpJ
YhR+wZ88MO+MuRK21Ly2VyBa9ZpcyfTabFK/TW63ANMt8NHnSzGJupc34MXBDdn2VBGGmZgiV385
fvOzm/beIoaZNpNtsZDv9GCXlE8jwkz6yBNHF6YzwMEihM4PrOBtI3UCw3+jMag66iDFp+acEGMB
DYfSysWFP4yEKusYIV85oAHvWuVrwvqwNkdnzg+Xub6QwRKZq8hReSGa0MSOYX5TuP0d4c/l/kuW
6d5LFITc71kIIP9/ay2SSKH31tLDx81nGubg/H/2Qm41puAqqlV0GRuqbFx9D+pNnqXxTlC9Kl6e
c7jdFrNkFNq9MtD2WE2JWmEuz3m5t4RpRdUM+gmTzxpneWEjdJ635Is7JIm6Pzlki10NCYnShqJN
gNKbkXx2Tn+v9VQE2va8VbtD9nYVe+gPFXV+RD2/ycWdZgxLUA5SE2XLUDX/wSbDjOBNbOJyTVjz
alonYqVO7Ui5UaY+oCGFWwxThQGFsusKfmq3Ht/c93W/t9G0KBDoFJnQFkWBuM/Ny+1RYoBoOO1P
4TX3Un820d//3H4zXhahYfh6XaGpPUxJC2LMb5bcszvRa6B+2Ad6neUwHrpMmU6qv3kGCv9WDvLN
VdK4hJPWK2WXdrgBUppk9zvE6pWNlVbZDI8s5790NnbscbYG/Af+3+YH9X4zwuptmyd+oUkhhmHE
MtUaRHAnjLARDJOTKIFxOaESmIWrUtp1z1xbQcjJq5DldGlP+4qbcT2AedsQf7rB0SFAFjXk0L3T
ONdFIwrG5VV/l/YH5M79tG7Yt6gnyz9t2SrborvlBYI9UZaxp2+VUScuVRxmY+fsXdk7jK3mF2Tk
bsYWCzF6QdPQ7nl7/Eph6U9/Ikv29ossg7EzH1Vq2cOHBEDXY1jtdCFWygr8RPLGQohjmv0hr4Qe
OQWJPtJh702GdHfgRuAO6fdWOAqQgtDXWRZIaBIV4JaaTLk3Abbget2GfuQFpwvix4mzoIXdObzr
fiUk9O8JiAW1h7eKJWh5jlErJsLURW1B2t5UiUg6hi0/Z5nwhDNNozzyGrWnKor4o8sQNQ7EMQ+7
LN2CSVSxX/VST50a9Pm+FD6eX4PdamJMEges/U3jy5Q/4XetPqIo6VmTsS2rTSLS0M1hBTzfhadm
nhegu+VIzR/g1xpl38s+hlD0N8PCOcC10I3msq0JSKAXLzKeGx5T0JMxbdeSsBnASB6IfLaprbSn
i4wwI3OmApfp9W106btL6Oa23CfrJqPOTPgwcEobKjFeuNn4YgUXXuYFQiAJIfAHlDwpAKk1tE+i
6zkOHQEYXMgyhXkUop8QjezyTInxnbW4gevpRKnEMyqva6U/YWwseapmVENPoIpuHbJgLowAp0az
00b4KWdXAfPMFi92jD1YCVVgZmwiZkYggPj7yfC7PT6PFxIK0E4ixzCOY8s6/sAi8EwbZ4JD8yCI
zwb1c/wQuMVP15pUddKdpR4RkPnM+pdIt+1BPx8ZKJ9hYNndVavavi5r/GrzM3GmaNlWjfYo9wxo
hpdWQDyypseQtRC3FNBL5Z4EmOoCvZMX1ZLdRPs5885vdHjfo3e7YDBH2LwegEdlEUPeB//+3k9U
iOMhnUiJnzmpUIGxgxIiNUb4dA3l2QN3Q82id6+bxI2DiBExos5ZkFegj5RyhHvzfPvUlQjBeM42
gmm4fvq2V+DKwn1xESRUKwiAamSnGFgS0GUeSPh8k5CuRHgRVJvy32HkULLeuiU5ARZO8bdRIox1
dMAdhAMDMn32kG8muS3JAj8tGon0Ea+IGeIy9+FIFxVgL74pCUxsDZYPFHjeJIg0W8/esNGa9y/I
I387mlvyfhnrsOuigU3/jEYADV+1n2JaoldulWt5+sRLDKXnkkvtEe36zTyLnKFO2mbZD8dqvy4c
noMUGjGxJdFvhM0DrwBW2UM3BUvnbkI9d2qTnWaYfhCQvYFMzGrTA6K1FOIVtxutTV62oloUaZRj
P3hrYK6I9s1DQcU7pLcOY5m9BTOCXcKchmd9OvCJMFjnFO4IGx/u7gcg6wEmXfwaoni+z0stphds
eP++oBslT5tDVMXbLt4MiRO9vC8OCWybU9Y79HqX8M+nCe1kvvHy6Idr2cDs9tKf/M0gFhR4Q/s0
inLUiQ4hhCV8PheRgnI51OJiFIpueyMn9mW3hOUGmJJBP7Fu9OXXwQM4OZQ2jNvRjfcAouQKBMg2
2F0Um+kRPw44HrNbsFxnPcelPdB5hg0C/UrfoFQkDRFBFtEmp6/jzDxn+IiFf+D/K781BexAgFSp
/WHJD7/R3XCpWLg5aghjYinwxED7l0hcIYvq3KKK6qp6DJEeQWBbi3MBRaI3FZc3wssfyY6h3c/d
YRxLjukCZpKs3x/kSI1pQHrUFoBQ6Ho66QkfJYY23btG16kcUPgNJ2FRuolFumCKUYrl09kJZY4n
R2jj5H+yRH/rZMX0H4EbjHcO/ToE/eAOgvpYunvnRn7owcXPJvoOJmz2y5HlTLCCG9YdkDaA2/SU
X23P7NPogrGHf40RXbykNnUMwfYZvNVdHku1Azp0FlA7v5ysXQum01jDJ6dXQuDcdwdH95E+jv5u
lPLrUST+J2XWiPCq0bXTgHaSHeT8wqmOR0UW0oznpl55NVDdBxfI+ewVtI4hrqwBFLTkiwfz1KCm
YBYKH+TGHDLF+OMpZokGkOpU3ycEl38i47abvpeXh1C/+ZhU7C3bn7CsmjiYJWpNLYK0PktPHuzN
wimFLaSzjCVThrv2/ZvavfJfmcpPiC2NstBcXvu+ccQZhCSY07b2mm12egy9f2O3XgJRr89IT/Jd
Sb8qRlRKTmjAQk13Lo/M4ndr02iqr3Tu/YDotYPE/oMf3IV9wwmSouC2Wd22y0Gq5KRnIBCP3SPl
trpmuqcBupPwkBWWe59ZTkuoBtRFlRVi+Ps2W/5EyYXKU7rIHFbu3UgdvMlcr23BDOr10NgUnQsR
1T0SsfIW0kNnMyt493KU4soWwFc6kwQ8WYgaG9EWO1DjcwiOWEKGrCrPUVcjHT5AEMy0xIYGQ5yD
bjXdURQ/UzBLFXbCB/uWtpLfMCbCh2qX7LhOk8XBfPw5IhT547TnSAihFMMWSvNx4iiy/KY3+sK5
pL6lXJZ6l+LAXL7YjlMal4xKQZT43KTSItdkdMqd0fR+1c6ENG+BV3/8vmEzNzlVP3jDEMioscqk
f9B5Xm2VPnBozCzjTErgNZJdpXZ98QF199yEpXUV/jBgQu0V/m8HtYyQbDf8Km3MKGH6FGstZAFy
5by9Y7T/klQgGjVuJtuV6QFIxfDcjoEN1Ye1w/hndsXEjAg6gEXe1ZeTFviYYJG7BhdZCWHK3cDQ
+qUeSrOSQbShCsMF24bQ73BfEe5cn0QTDJZ1nJBsBZtYbK/tIVKgaKkmk5lmKHsVVkq1ZcTZ0h5r
OlymDCjS7szNXBLSy9eejwXxKGmuWFKuVjtPZRlWp7LqWt3fd0hRMW2BtPZwtHr6KDSRoOXVvba0
6ll12JCGUQ92eB4b6cKHdY2neNDiTAYhCJLG6mr5yGeVvd8ycxXRiSHoSaK5cdTZBWR7rpSVvOKt
smWFs7ZoxtVSrOI+kXGLOcnj9VXVwiojUWpPzMoMdcU+d3YHqIjjaNwnbumg2bJWzFZY4NN7BkiN
VxykU31XrSebpOXyc2fVxTe8m8xwC6PU8sx2FyzpRW7bj0Quupiy7xXv7WrYkvu9XibzBUxntLr2
+7iPnsDykV8fTHvYszGjWYJayTHR/7HD4o6e3Nlco4/WPgE21W5wSguf/JVuvqbPgPgZVjvk7Eur
r2cX7re83dM4cP0eGE/SC+SfKXB1WbWTQTVw+kKHL0ma0z8IZbY+r3deptEFctLdUX4621QjnnGF
qV+14A7OBEWqyTHzKMv9QqnSzXDJgGCfA7FaIGTbvBmBsHdTCPjxhWN6z3UVg1c6swV/2txS8O3A
tWIIv0Ux2PnmRkvkV2KQpfIg3m0++Os6XqpFQ84F+hBj7gk8kXS2vZAieBHM+mzdA20J2nU2i12P
9myHrGJpawfrH6QIz5Wy6lKYEK29rAfBrmkNwcz8Njn53fTafcvRwDMc5jnn+PbPSrmbR9rvljki
xSj272HyV9sN4ZVNQKpAng+RxzsvOWvIwxSgy+x/ifu/aUizZlMh9BfeqyQFrh6t+UVpWBm4Ud4A
EYwRCeuWibi2yB/I1Qne5U0OkZo1uj5Q05an3CftSRSvVLDVn8vc3omlmUf0m6P8UfMeYTbg3Cke
nqHwA9ri/E+RX3VNjcnyNNBvWLwjcoUDLmFu8BGM2xHN3BxslMguEf1q6+HKoXTjP7Nke5888ITw
AXLJJ7vrRXFGO7iOg34aPKb5/7HCaQMpGTVqYGY7P4rjj+N4XcJpwOhLkF+QZxuAI13UDWkIq9t5
tzqnXgstqxd/qC9dUPruKa+iY5K9Ct6K9aaGdqNH7ir+NJA4sBwdhH3HUgH3+Ecwsqo9c9MmyO5Z
F1FNzcbwRH+D1vTBQreKeENUmL6AbimItokQk5d8smujRlVQF8FKoKbF0S5wGkE6KIKsMqxRHU4E
8X5h07h3kWlfmbKBJRrukLfKz3Wrnk2N6J5tWZIL1wNgaiBJgTHVljD0x6do8rRf8PyUbuYHf3S2
TZevbYNEOfnl0XBW5je+S4MyznKLGkaB/0Fso7L8yl7qSzK87JcGhYW/r+DKRQc27A52flPp9sef
XZEOeH2vCud164W0grF4dSWHOXW/6Hn37SX8kRQtHvJ8gaAJ+CV1cDZzm/B4OXSytFrbGj6eDFRv
PtEs3jUGA9yXntXbCGNtCzE7wvUV00nL/mkf2VWveBif3Hk0a5t0MOhZ1WNHjRL0D9S5nF6QS9b0
QiV0t5QyrxelNiyu4d+n8dcjshwgbUEe4iwVfDT1+MMU+IidKXCvz+4BcZl2Yvy/KL/B5R32zhzX
ntlUk39S7VZ/e+IHlm3DGk0R+EaMW7sQO7rvRb5Rcvk1qynLwVKS4GazkuMpanPxm3KQdnUqQmfU
OPjwEXdPYh6bWKr6b3bvP3CpiQstc/3aVahXodYI6R/MSHbC5LeHRCzTDI7t29XytebaVWz5E1Jn
e1yE7nZRu9lM+W7zG9i8kepu3hyd1de89gB9xe2H6tKvtnDeiPiLe8JQijfR86nun/1DCJO1ea0k
IuyfCRzvQA81gqarjYHOOn458MyYxI2BiUuKQcegtufdMzzulpiolAWwKNnXd+NSJIqbC43bhDWy
83PjQnmBwOZl5amO4ZyiQ0/AAL/ssKFh5otv12Nlp95okS702BFrI7LP3kIw5TecGTjXQeMtCCxC
cDe5K1EPDsl9oemQ0HApCjX6Mna80ubg7dv2SX4o4Axz6ZH/ZYwEQ9VFxWDPLW+XjlaUjTkLMnBf
ncRLg7O7fLMJYAFB0My9UzCJrF2lzpawY834fwA/iiWgSnvshML09TXugNXVVJkJQiw0Rmf+yRzw
WwCIslbDDo51oLZ2cMXcojctizymKbb+HYJLz78QPLfrvNvtl+iF/p3q1b8Ol8j9b8COdCPLyg3p
aopKD+IQpueQqAY1o8OU48//sw6xexeqieJLAkVOuqo1Gz+mCOrCZiY58uN4awE65ww6P0gqQFqo
m8bM7fU8rvTrWNbbeEGSPA+A2QrNgKHV/p0AlDEnXOdVGWi7R/t8yVC/vq1Xz/lekiyKawb9duI8
Pbkuf0/tx3lLcv8Q1vApdEiLJgXf3StPyurQZng77jJqlePLuzzjjN9BMrniUGU0iYuWiuyLhKmE
1B3X+w4VTSVaQnBckwxaR//z00MyHBnUn8nHXl6ydB97kOxZn8i7nLrmimJUbGIWiqLZE98C9NmR
PhYBErr5ks2XmAXz+U2pJAWvm5d311rJ9HbwaRjA/EVAFxvKs02d1NnP5qrKqZ6ZSSL4YibhMRw3
94Vfjuc6DKRy2JJDrrmmPbZSL8NzuVyHux5Y6/wd7kapesyoHgOPAPdMPMvvVVfEwTDsJp8HKtmK
q367LoINOTprz804EMVetMBe9RDbElEBWOCEz1/9flp/QQG2aAz0IonU9WpyX2jFr9JpyKdmPcXE
r4YAxeF6pLTTELwz0vqg076v56zQsxxtonRTTZYC/D/6MLcFcz8T4idp+q6fndEVPyXbeC9fIa6X
b42wtmZPFSBy/dafIif2RfEKD44IsUJ1/5Zra9MuW0AisRCS/f18OeFpXLGX/Lrjzbc+f2t99JNT
wKeNuuw02Rz70Cmjdo7Stb5dDVQdx41VOFxKeJxh53SARUOZUrff1LSXmdHGuaxIK890M8tnu3SD
jjWcE6XUMja6EiSnglflknPbbsFLauiMUELr+ezbFd4KnmDdwFZ2ueVkQQN9QtZ9iVNEdowU8csF
DI0e5zBDvHBb7ae7/6g6QaEIZW1Ni0pt2rdWbqZTHoPisWGCRaIe7OYZqgeihg4r0gbzaSyR3TtT
CR1nRNQRqmI15C43iuhH8EmxjTG9sLwktbsX0A/sceDajzYcJmMjM21IiSSwWk7RkgvovIgg1AF6
BiXsTeUUc+K8Z5BsdYdzKmtKVloLVVq/MVYRCowAikTp2yvGicaGfT3ch0BxCLTw79B4f52Gcz/Q
gsiwsZcJoPbiQ93rVpnIrSsL0tDZpLfXcRlp4cDce/dBt29YDOPCXM+FgitVUw4unGbS3g/ds8vj
F8g+BybX0cbVol8qcTy5nYnxWU8keEIUzxYEM8O2y317kGpeCNBIw4BE+zoF7nD4/8FOtnF+D/uC
haYrW+2BRQUyKu4bV2Nlivkh1v+82LoGI7zXcgLfT01SGRApMkgZySRZOdNn0I7m/TBdFKlGXqyH
qHVTUG5xb83p/V5emUfNLUyG0p+KYCSbbcWPFI3VCJVfT06DP1RltVt8EId17+sbgEfIYQrqcox2
Uw0mpNkSUDGPPDyUoYBsSdMd9hzfrt6ytl+Y1SOpq6J6JTv/yvx/FZclvUm8Ng93X/2kHV1dEzWL
WmLdGmEg1lvsdb1V/epVKLott248wL0qGitdYT/bPPkXkVyIgukbAg2+0gCn6J95ZkkL8NrpEj7V
eLXtyrDtoZ7Av27zgB7gdwT/ctxcVuii4e9/JKWTx0orIN5mmUYnsIfnyA2a1j1ofoGkgJ6RRshT
tSRd2vEG2HmDq6eBRm9PtOXYEW53cZM4jCeOYZ7nXgKF5Qy2g2QjSQcii5KUClKOg+D2jLd5S3oq
zBmaB+QFjCGmB4WBz89ylPjvtke5MKVhGrlmEn/4CgAzhkvapxLV7z74VroyhDgua1fRmTzluXyH
ofjpybU2yKdTlCg3Asf+vdic5BbrbQFTjepfX/GESGywxK8PCaDs8pFOEIS1Qx0lPHgjNswYQMfz
vlKu6p+12KfaigDWLJmHHoLOrSzdVYGcqdeWzTtfueC08CfeWQZhWbA0xiyKhNA/DjdBi6ocMfBG
lbHubh7tXL5dNwT+uDnLmyOWpnw1gM1DWtjjgB6FHCfu89XP33+imozcwUkc/VZ6rETXHut42gas
PUt4ouRTq+R0ru9FlrIpvXWIW5nndxL+RJvwJZnJWcIIJTQCbp6A/2V9TBV3nPZj+xOfelJBtY5g
w7l+2sn/WhEGa9Ywbc5Avd1pjbJYfJOWDB5oQfk314YfGNLhm5MUcQ6GurCKl24iWtlwGTbma67b
HrDuc+ajKgf7HOAMNvQsi1iZcJ+amKTaDSZ5ICSpc0YFmdD8CSS2kRqB2mX/PtxIzz6MevcnIVqh
ntzQzw/VCj2hLYKcvdoUKm1KR6r2BnKvsQu3kcfOT0Vh5KROiJwHNuEUvzffDkez2axQXcYv0Dpl
kOEdy/0PJfQRXfFRgiQUH/WrbXMSWkgzT3wBPIUiT/0Odxv6bEWJOv2DWG/LjdUrgRQKySmq3tDu
LY7M7fgx3iIRN8pfOgtWnR7VJFF76BCclkPG6D/A66Zz7seR3+fydut0yNyO+r2bxwiNvzI9jJJD
6KXkRh+SM8ELGgSmmiDtpmJMEqPDe5ZHHvqoOXXM2dsHHueGTjSujMJdDudV8k7P4NHgCuPdHWW7
ljCjQbaMd5p2jHFbeiGC4T4sB6y7nS4ya9KgrRZlyBVLPkhfccff9XAz7ie8R1ATFvSamkio6XBo
z+7GwOASGKRiYW0bZouNhtnEVi0T7MV5jWEIvUbP0tgO7cuQJiBPiB4Zqdzsov+MWqb1NwpK0iJW
RU6zSjRj/8YPyIg0ue8sFhX2FF7ieTfjEIeu12DEFpPyr3vMuq76H/C83rng9tKnTM7wgo+JXvzY
JVEND/u57wTvOA3mnt52OmxX2KEXC7p6nuRZBnJFvhB/hiTkVBSRHUnewb6GnQIdenQ5HfWYuKNp
4ntr3MQCw9BQKFsQUpaXUL8ontXVCTgdgFhOeTD95LaukI4HFwkEDwYWrcoewfgS/2JQx0bGWqPa
WoMcZep9SX6d+QHvxXAzqUtEJpGzLhWYW0jw8tKL7hXd49RUSM+RtzEByGJCItx9I3TDRA9LhLO/
nIHR01JU01Re0FsQnBBoN4dggOebZFp6q9nXtwB7g2bApfGzCJSATrOpG8tkvIdPl84s+Tfu3hLH
HF1VGme/Vv9Uy5ZMFXcJmHgeaAv3ZP4WpOstaiB4BVu6+ceign1dpfntFn0mVn516dMWDBrcDphb
GPUd0hc0XDuOcEijnBDcghh33D67IQ9dqt6UmGzT0YPNkK4MYid3FG6tvqwM+0Pxim2VzOz5x8mI
bkuTLmYuId5JkkuxnPR6cPikZZ8Bf6lRzoY2Prgic2dRP2TytB334gN2VBuMrCWhSCwLEDZtdE8A
ZOnE7TNKhwGhTKc+lFVcsx4tD6cJCTzuOEYSF8Kd5XEejy/K4FZ31hky2UfFxvCmpQZS6KrKW11d
nCXleVTyDZxq8+d7pOCW6vVPml3wTJU+DatN6UPk2t1F80oUFzJRXezVeyVqadXvCxuM9KxKa4HQ
tjU1OyvjYfT2vSnOIO0DWfk59BakbBVLz5ikPghsIml+ZGqFW0ynH9Rf4+izRbMTwgI9+W2bFKLm
jdV9+cXJl427GPhnBgReVOop4lBREQRLDM7UIlylJ6I2VgweR+7u2K5r3irmnprXlXHHTi46G0kQ
1CxkjdFxVdLGhGYPZZFbgxvm2qt+bgoSlx10g0tZfhuhqT52rWCGmI6h68hWHWToFsx6noS5yg9q
R3Fr+gw5tLkxVJojmuhwS19+4ZA87nO7rWWwaGx08q5W3NMd3IVLr7KcV4uZV3+qmBN0zXiDiupN
sMMSjrj2GW1eIpzGFqMYO3V1tojAKQNmGP+T/kVjgiwpiHK7k0zkP73i7ShytFR8gWLMC39bCmkC
INbrQBttJnE3LGUAsMxsVtft7msxLEpNomUo5bCL7Qw/4uHILsF2amKMNHNniS6Kzk1bSg0knSfo
0tGJAWDQbmnYlmoB1niCcZO1h4iHda/hAIaL4pkwIS3FMxbZzQjKCod9KUXTjAke81O0R+Sw1sSb
F2SRvit7VNJ+4lC4ozivWpS5PHSRWeSaDO+GZV7+iQw0mSzplZFfgcLjPj30wY3wD7nkpNfOmf/Y
57cBhcT2Yj87DLwd4eWpZv6Ssl/OR92/+ltJgceejC/4i9hKB1962Nw6VgAo2Vh0Os2k5QKhcdEw
Jng6iYjrdT+nuxCrEGr8kjD6Urh3ECvHPTvtTGXKSDm+AxtIF0u2PH/4MYdaDhy08T0IASl0HY6G
YviR0pgHhPFFaAGs7It26FvRE8RgJVXse4UUJHHGlpGz96pX04U/qvBIIPFzxbpuREK66v3D8agR
62x7IXw4h8Wyc84AjXuJu/2rvBNDVBe1jIVStnqGp+ma4Nk6yD3x/2O2xGo9ERsXYPcCSD20Ig53
MVEda0FwJ4VCTd9RLTmNJ4KXJ++c5njTSQREtbQYxmcm8a5qwZKlb9ng/we1UAJem/45FUd722jJ
UegpqOWzl8Q2hwqKByFk4GRf8MMm539lunPHCT9Nav36U0bEUckjtZ9VifN3JV45kALee5hJQKE6
NGRoqcEXW/HVvD+oH6B8MoypPr1OY+UACLE5qGbn+rprtcLVCbkokO9A+wxCjx7fsmGXdbTdz6ve
k0EAddodFytmFKrF4/XakDHaKN4ms927V9bxHOZ+oPiu8WpgOUDWWbKS8rvcP9H+7FDpzanO/oJV
jDPY8kukSZOJ1rzAM4Ma5O6L7BLB6PgpU354BtviClI6mFgiy51S0T4Rj5OwAgtm8VD5AhK/xgra
OmG9XEVAuPItPU40wUb37xfRR78Pdo1DzaiJF6869qsIiuXZWHv9YUfzYdXUn37zxU5Ia8BMfP9U
2U+vYujXcCqvXCGhELatr4tXtF6LNdGQtDldyOUL9se+wTTaBZ3DfGRHO744Jk9SmucyocvduDiE
THZgXIvfQSnE07by7IHF0BEh2/XSpQZfwZDbB7iQxdunZLEgylyIBzE/1vfGTFgeVbP0AElzYCfQ
lnutxcMjuGyX28Z8uaKd+2c+p/i4B9mIdyUBhWpYVI7UNH0lAcdhovgq8tvMRnx8zlcJpQ1ci6+q
rg6HM2N6f9X7r7w/ieNi8yXyoobWuT/r66RJNBR/ELkipADL5ienotu4rMcMWvd16nr6ul4ZYe/A
DNki+iV4Hgd8yxRElIRx+XmQ0s062OCxlVQ2F5YOObPDESRk/wVIGAQYOeRGRDZ0hXviMEhiIVbe
xexXflHJlnojtDDEqIPGfvLiBlFuGsvG2/Ibyi4FuFZxTajLheev8LUd8zwbgVJCnByi8oZlAnMP
PsuLfi7m2yaHxc7QwrZzIrLfbQLbC2tO7yrKq93MzGOk98ZHvlxwYKvC6q/6LrywcgWJ0+kUKSwB
UgO7qJOFCfGESxAfTJCO8EbxDVKqL9fnToWfm0SXaC/CiSIoTCUR2St/z/lCZLnQB9cthjq5Hcv1
sA6cQCv/WK3se3Ejbxj1jyfiSjYEWF4cty+CKqtRSGVXN8QH1wWkg4u/jNKX3a7L05pGS1RHpwI7
c/7cCcKKL51oSWGfEjgmx4ZxvuUP1j2CweQwHdaUOQStOvXiKsRWppWB7O0nt4sk17rSaJ5TWSmo
ZhZkW2cWp+WXXfmnm68R/s9BAchye9JHA9PbtSTrsOt9yBtTq2P94phqwbmGdl/dV/OoQlbvukVW
ZmO37uFslo48o3ahFGtWFOJxZtJs8RHTSvzApzpLIQOjNSl7Kvqmy9qL9KS96RqK8j2xxKWHO7kD
EGzUpAraPBO+CEK7C0sa1VjDS28zqJByqp8DPouGCCoXvwgVNqQjpERUQPn48mT+8/tasu4DzDFy
Wz5Yz66xyK6Gs0gu4xkoy0H4zEVXXzH6lRpzXRrSFE8FC16SDmsgnw1AKWobc1/v/eldQlZfTgOr
mAwJ6Z3wUZyPyzv1hGqfeRae23xNA3qpzQhMQJ0NKeUJbw6YM959nQQoGmJHfCSW4x0Xw4NXIyIF
h1fsCDmU/dsAgbHIoWFPjJdjfRDGXbsp9xbAVvT36l0IaHFRXzh4Z2ren0PDHKQqpLBR6VRgPRS+
EA/7j4P+mPBxfhSDF2fgjvcO5csneXMOI5vlY3I4tXMBz2HvF9btcAWlKAHESo/oFLTXvl3IyRnN
Wi0/6q8+BgHyJrszbPa3sIQA+sSgpDL2ZeY0u/LjhWfmrU5Xw6ywcu1hHygsfZH2/aSekYt2NPRX
EjGTPaFj+5HSJR7ixqkvdhJzujoo8w50mDf9WaUHuKDUpUvkKZf5kVys2vbDzul8nBSyGWGo5VtM
w7MIHuddxv99g9NNpvh8N7pQNfRufGMMg68cvhwFGlnYBi1u5GN9sR76ll8fo6GsEiqNdcgLsGNI
zhQzi+i552Z6lAtk5WfhmgUs8ZoFNX+5fS71qBoIGLFusf7yLpwx+vzGOSutJ5T6NoqE71EDDxiE
x4g9gl+rJjHdkLpZXzJwBXsixniDlv8nrU1feg5aRC1PZt4qP8QEU/+SGZHHG1UIvkUq62bbw2LZ
R1pbe6Of06GSMTAesl1L3bzvUnOAdlQRwee8jiSMFUNxf3ZMScxotxX3bS59C/FLTyxYo8xUDpqx
T/V/WWZv9kxmfwHYradXP1ybeAOkt2NIUEDrJB5lcjSFeHqAdjrPGYoQ5q6NI3iaq2/lba2cm9/V
J9NlMwEwxCHNrV8d7oGDs8tt3suZ4hlKDxWtNuTIXqrWbTbjaF2i4QiTflklI/Ey1ZpyW5R6tMzR
ypXLP2qVxXnX8+oipR1GnHY83lumtU0Lg9373gGmKyFqW+PhXCXG5yyWXuuoWKjiODdYIMIeWY5f
ACEbVjuFLdxz/SIXqzSe+U7qLDrX9z05JkO5xd23276w9nB02JRHAqUOhkUnibp0q34oUa4gp8cU
2O0/r633T/IaOzgaHX1M468TgcXsbrqughNNrggUmxZ5dmsL5Y2p8nt24mmhPEYsVXWvazCY8NdB
iThkJHceRdE1UcZHgI0ZE6aXmoeI8Wu2PRWYXetHc7KaAKr9FNP9YWeGj4uizM0ip/QBAhE9ZJmX
lvvvM64u7E8PxdXUj28pT6Iw1jrzLLEAg3AbNOcoPw7x38COxeE/QzS3+BzTAVLJ9Szb81u6LQ61
mPuYXPnq+urPFK4vrZ+hboOqEGqIImivF1SXR4H7aaKdkQE7iHzYqXpG5DMBpZH4Ahecy4DDf/ig
kwfILNpEFsp80eUqXABB2y0tx3T6QUhX1oGaw+ZMHNKHOFOH80l1soulBAdW0F+W72SSAi5hiZiS
rJrrrXTGgwPGV2xM5Z0SOXCIeCWj40xE/y70m2ncP/4U4bgVr4oCa9j3BQl7oYWNCwhCGEJYv+9m
qeNG6bqp3mYTEWWNuTIbRgf+p7kcdU6QIAvNH+wRt4mM2z73A5qdRh7NRBduZlXhuAk1qnzHx+jH
74ZVR3ji4GrFW5Ty8hPGIJAV2w6ExTBCcrlttWhq03LamHW+T0m8tSIYaUqt0kCSq7ZW8xl1M3+d
3NGxT1qA9TiM2pg37vEOQFO1GHg7MtNRwnGob6aS183rlWUac1KK5Pmb+Leicqx3l3w2bt/CGV5T
mUwbjm+/VmWejnx/4Tcvox1Rfm+R/A7pVo7fNaHTQ7fx1P38Dc8TEqq0Tqflng3euoFaopgsTvrY
jPyoD+dwSKtsh4B/v6iYOSmTdYnqh+nPO+5IBICHpCnwAvY7mQyDGJotBDKSSg9oB4z4BUNhZA5z
/VaFW1z8Hf5kArYLHRqbGADmDJZmyDUcwmgOSVyTKRxRVDDRLUXEkO40RGOgRPCI9pIlkGbJBrJi
/D9//1pSS94uzDaox1JIZ7YloUTTN1ZIUQFFs8b9v+5MzUTDZKMFbythRe2oJ2aBTSVof1f6GHew
8vp6xEiuoPfYaiiqsPcDY4imFi/h82YtfqXIpVwv6VDxP9psYl6gncgNlV5QQfD7WdLrRpl+mx0l
5VzcqwPGYRarnDJKVGBTg6pBPwV+5iQ1/jnR7t6hxpSMyC1DG8htABtj06Hk2LwQGc4RNkV+wxIq
ad0zE3D48F4XtNlPcMKxLzJ3xSzOteMPxq5ixvkDfWX2qI7GWk5GveRBhwF74NIAuJyP4yj7uZgE
VzOXbTUC6xrXpsXvs/XnF8MXsWCI+0WkZmpFJVWQJtvf0DSEmFisqeez0/1wd+6Oh/Tg5e1VdTBO
IFtm8uXt6gQHroT+FE85vgowMRO6ujR4ddOq7+8xgGtHKNIrON6gcLQuEdW1J2wQmqJce/vcP9aV
t+Jy/YATs3ZB2YLPx6vRMgojhe8ztqLGjBU+w8Bx+ygnjjAfz236ryWWPPPD00ylNml37xiY8hmS
y56ynEqEThcRb6RCGvybKJPEmzSWdrr1PVz0JBAlXnblGeGtrAh1m2CWwt2rt/NQpfhAjI/u/V/N
KKW3KuQaa2b+bkp2/rCNAGYnhDA9GtqoYZ49C+nHN0qXMpxmbeFP26XOaOnRB1l4yMZpCWNVRaBW
19w/dD1NVsM0ay3KdV5iyq92Z0001extknnQic5T8poF9CP/H/+hysroWk1cb16aRzjSB9chAqRl
/j14+hjhOeJOTD7thMQYyWUlMlpofKYIU3De5rW2kbpDxEZNUoATUUSsfpZGldf1DhmHPMp/XiF+
0ZS5lVbeNMmCoNFFvHylcIZT7uzGnCyEK7KsKAIC/qCNgB+5+reshbJY3OB+pjspjCS4DW+8dCZi
rnJvrrMbL11w3AWLJVpHgpdrzjfoYQ3RyuCSKocYHq84/X3DVIT/BOeuyw1oo9PC7Kvie/Iiqg7M
9tbJZOT50Yn5rYHuRIJG1w1UQi3F4qrdRlDWpyS4MD+gXuKaOiE7xaIE+ww15dOIUZcEb9juHnPE
mO3mDS41TTpeJaO20upmNbykOHRRLgOdLiEiwOdOZ0THSzidF8b/6Qlbf2rXK9dFrbGLqmDcuDJK
IjNOg5MagjK4giOIymAS7Qx9r+Wv4zFpLiisvYMEK0MAuopnleIJUigLiWS2c3UQQmH72u4AFsjC
XnRyokS4c7aqNfkUQsv4J+EfRhYViEB7MlNnBJTumzGotbpQgTFIqKklN7OtWI4ga6rfl3frZ15T
XUpRdFUC4PQcg3eMCcEA50HWsOuOyYywD26qGHUbBSwsL/rCJ/EGFNZ4eBL1v1Pc2OntivvC9xUi
nZXyiS85JVxHmY7NGUQ0lHAp61SzxRDq3MPWEoElVJrXD4x7G0+G+KweqEcUH9vrDr4zWwAdmx0/
YLZjB1a45arhiLYfiWNCw6bzWsLxiCD5uShunJVvain5KT4aKvVPTUlGTAd6/UtcW7AjaKhIGj0E
3lqe1z9s9Rn+mJ86A0Z5fkcM3MEabDItY6Lwgf/dZG5F2jvHJeQhwxBdbi7045uq9ehr1qYLMp6p
Dh4p36SQIv3Y5gzSiDZkg2NAUdJsz1Xd4vUPdxrcWlYHwi3PfEsIs8LdOBq9tvQqUTjdDREX6+RM
2qruix3upAb98sQj1iQ+uscY6Ma0p2nP2C6jk8e9xFIsGuYVV0PixtTAAPFMiirNsywgGp7hUXed
FHSMgH8tVIXh8M2bTyA4JXgY8WVJAlPJCGKglQCJxkJMHxBJKZCVd4Id4H9BMIHJjjIKB/hh/xJL
508WOFJX3mBlZOO08RZuVS/Cuief+bu3kEYSEdWNKO6DazZKHdvnh6rLwWDGB9CN3b4bTjy/INpD
kn9Sj+1rW+POHjG+RZBmyQO0CJ/VKqNhh3/2KS0+yDQ7hdxVpu3lewHuYCZsGbzmbE7EEInWKOnO
E2Q92gYvoJm95NiC6dnWbJsRda2gIsUFBdlYzGTcXvvKBrfzfzNDKfFLCt/JtaUVWn3Du0nhrcC+
W1M3JtqrlqAoqn++4in9pBklOJZafOHA6P2dh03K4YrB21H2jRQUDJkRwx4qOUYpNZLosRUB5jco
naEoV3tKepKOunyQsuYoZokr5TvFNBptSiQo4dJ+iREq9CV6KV/Miyi/QuZblDRJ2DDaX/AXYhAv
YMAnGtY0KTy9kJRFWtSkJFFzB9Gob+xQahKq9gOQlQDQBdnfnedQqiYwHuH2oLRNasKyRhUGH66V
vzUKsBJyDJ0vKGs479jrURi37ypHFPM7LuJ55mUFmurP0ZoQl3+SfHcL3tN8Xcv1t3iXVfDfbw/w
iCmz1XgCowSTRkACdlXct/JaIPMUuo0f8IUkOxvG+5J7E//qko5oJigS2YQB2jnh9eEwVdrADTel
mPoFJp1/It0AdmWBlbTU4pKwChFnk/s9ChZTwrGBc7WhCw35+i5AQcA90IWBfd8Ke/DmX0IQJcd7
6P1yh3g7UCWtsmPyykZtbtby9wWT2kVwTBqYyHbsbh0ZAYxx2RprSLwIXp8q/b9m+1jQKuEd1lyC
16uO50I6AuS6mos3PlS9L40ODyKdfLTfRsro/qjkHb66+fA3i2gvSyVyCfyDkXWN/BPE+uLKgQqo
zVEVQBZTlKQKl4QmBhjCenwxzKjtyisgTKY2gOwoTnuoL6If22yXE6E8ZA2iw8nmVc0YqT9lGmq+
Zs3I7FkRazpjjJsf0it84sAKQhw4laNl7LzCxOkXScms+i/sztKo/kA7YyrvQz5hJuSOQDLdk0zA
HIT4mwZJzu0Qxi3v3AVOFrwWrFa30ELXLCgRCu1QVpCWGWfw7HPKjzkkl9mf7ckjtg/1Nwsep1Lr
cnuCycjZePpcEdrqdQ0Gr/bW9CPKzIFAvBQyCKqG2rXSGdgjM78ZKMizeHhv2zNkGoO6IfYiQQXV
xuTUsv0qRZZ66m4Y2wfEHRaJmt6wszDJ1pLS+PMgjzG7/fgebpvJU6/v15R4zSc52+MONiw7xf17
dy10BQimdAs0EA75E1kHU3uM9NjJJiXPWwhBbxEhzU384zUvPY0zRjMXV8cIBtjXm7Y31XHX9KnX
Esnk45LTKHFchdm7YZsBh2+Kfc8UjXXjX6Us8mL3Z8d0MJC6JF8Z1LMKRRRclP1RNdHhMQW3A6q+
VUkJNBKtpBHx8AVlhC0HuDfl2vaLfFrWqhgll0hZicP58sJLzozhPEuQ0aBrtfv6IblF2er1uurR
hSnH5VQfkMQ7yht5JyXXGvc/0vJ1ZqvS3VmDFdfm8L0beKPOm/XxWnjsu4oKNkMA1m5ycnw9E8c5
A0wME+y1eIZV9RNJUdC/ozp29xFneI4izrfxTIIoXa4v7vM2n0XMaZAU0xWhpwEU4K0gzNg6Gd79
zz3s4eUL1zd8+x9Kk5F0kiKQMXhf+PUmBKEe6dUPkdgHo7YEIdVZbmevOpcyN776AClA8rWwx/MB
nbw3jDDDTRU1py1vL1dOZrlIHF9G+rfCh8/K9dTGvP+fsFeBCTH6F+wmn4jyiuvCm3GV+NRJm7rt
aCASbwmScEvQNxqld5P+Ls8v6b0sgxfwsMXS3H21Lz6IJvD+bVlUqIjrEtrhPlKNXlJWFocD5SFe
5Tjn/j+VKSmb1y3R0N3vkdRRH/rfJzV9xVGCh9aSpuCPL9dgh0O/JBPyLln9/PpNzSaqh/Dwf/Sv
YcmRMDEVqSfQ1GZLkqJX5ywG/VXUM2t0rrFHv9HE4WCjR3o6rvb48mOgiRysL1lESGVOV0LeoL+Z
m2wfHLqzC7XnqDgKjz/+M1nKUj0IrA7q3EMirnDc7rFU/QZ/rvXb7o11gqlPpuytIbYEd3CgnL0U
h3KMkJQeaN8JMVeZ9QN2QfTnR/33lnmZIAZBx2t98kHCdw42b+3TTQ7YOD08cct990xRMpLNpRRX
9xdVNySToDKCLP0ImdeOrUYI5UIVc+fC6CutyDnw3Gj2lGP6seFhzmZYnxVFzJctH65tgjrSJA24
mpO97ZSj+3JbnMHygeKHuzsC9WgY/30jgWG38eb2Rpcmg4YeJAPFXsK+kldxZkO24TNyAPKb93jX
11jSL1aokvBqCyz0FLW2Ad3fB1pnbLFI/sYskfbBEhAJqdGu1d1aZCEDXNDbI1AhBzS/mkTzKdT1
nCTJPdPw1KbMoh4iURSF/1al3wucu25HwjNHN4KRA6MbLqhJ94Me8hR5VD4Kvi2Dy3XHbdeSLGD8
cQ1OlSMv3ucIUB4qm3g7mE1hQC5ysAfjBUqkPSv+4aSPtvhyJzY8mtSa9kmPrVy6KclDW0UeCWHF
6XphZglMxIIWcHWwUTDnuUsL6Tx56NK3qB0/Et59Ocr59PY/6XCMWD/zUB/jO4n2udWDrvTtHb/i
qhd6NarHP0D8J2qVxS9MbX3wnScoUvUA7EQ6VtyEAdugcAaM50Kx2CKbifKvlSAyg4bbXi/fiC6p
J5n1HxeJJ08OiKhYG/oHraXfM+uWi4hhq/rf5MKmKn1sOsRtRe+TEWAwy1TxuyxdoOr3T6LqT4oQ
MIArMwLGp5fQBVwYBneSLTSH1cN/LStwkcIFsJYQ0d5RV7kjePgRQhfK0h9fL47ad953/SX+X/p4
q7dl3UwGF9Z/VMfhXdAUYf2jWPB7P39E9sHhgLAcTvfEjf6HPqyrSTv92diTD59JsSkwMVanF/76
zZ4PgDT+S3dTNwGns6iUeN9hn14hjOYxTtV7YumtUun6/e+xttxno4HwBVqwlCsQbFg7I1Q5A0Rg
owlAWckrJpVBVtm/WEF/6U8ORczvWmTj+Oyzp0UavvXQwSXA1GPzloRdaVM0RNd+1ATBZ73xFSXL
Z1ZPWfdYh2ZFvQDG8aJw2sXrKcNMzQHGfs3z/w5V6X07oNdRpoIOa531fUQtE84QclAOpUonSAVu
NCQu7XgfeF56JAIKeA87m8AwC+1I2GRhkyLICAlB7uzTP+DOfGqODnvDmnXgKJml1fTnw9oM9d/0
td6GdqtvQtEEIiEnuHjB2WAdZpvBYxxRV80DJHz2QYriPrsGq88SgGROAwfDWsZeyEZ/qZ7Cr5xv
HWUaa4YGmAtJt+4XzhojhU35F6nm7QhegXU13wqJ4wWUjEUaVLEl6NvQjK1Gw/LKHjhpT+DEyEtB
reuTFDXGjPrbFc9mfEF2dQhcs0K9ZfwGl1dR6HORPcsmorhNZEink3sSU15QN15dJbCZboeijPgt
Q82sdrZBZy0mSVyXdRnEhjFf6ktYYxYyMOYOOphfIuJxD757KNmF8AauIWq3hj+qx/QWrUGTDNl8
32jrYt1RIO+C9kqs9gOFUh3SfJNcOIkfX49EX/i9WVF6R1gfMp81SdNpjm/fklgAGPO6fSlDnX22
Mip71tZx0C3cmlG6RgcDn0ryGFrg7z22hHFF6ddSXLs5qd2dC9qMpQzGDdjyD4tLUhAYXh3P8Snc
bzB7ACcz8xFioWBSD2tC6n6qcoXUTMMmTE1ji1+lJQRnMMutGISPGVjYGS6d9EYoLujd/xHT5dj3
KM5dr4TILWJd7G99O3Qv/T7qZE3WgSwqps27A/YrzL1PsEWpdslA/eVsEYaq/19dDkS9k9i3o/Am
peDNqWmU7aRyGw2Wfk0yH38pj8zYuOtqAFWHJXa2apAoaIgxZQG+Gs0dCc37Q/OBXY4jMMw/1Zlk
muvnT6Ny24LCOzUtIlSLBEaVBr24fPR/KF0bab0Y4s77FVbuEM4706VnWXPJnGWPweLtnm1g0jee
Yi2sr55sM7FyKa42PsBISRLjZoBfAE0YJ373jrRfhT/v4CduvBd7fxCJpL1t2MOkB7JntnP8ubjL
6r9s3Zv9az83ulWxb8Q7hrU80IMQSLarskRg6qahKTimq2oFeBUA+RJ2FvytZPwOplAr5QUidN8K
BBcvuGyzfQC1oGiHlxIs3CyRU9I9uFE9rH4SWEaiRYvScc0BPVb08l5P0vSTDL5hCtrEXG3sSTPK
mZeK4sg0la161XOWMdyGkaRHo2nnmQ/rMZMyvZ8jEPeyfSRcNWQ2Dw3+TA7mzxWOYMyW9qGkn3hW
rJHjfB1qDqUJ5gP5V8YXocPGEcgS0EFSRpaY5lWZLvi4XU9IkrrUryRzy5PeZwPixGm782Q3WUrY
5BlhLXFqkscz4NTkSJzKPywLHX/wOng5osGib/nJHFqMnho3SwO02xGFd0xnVatBMsHc4HnnMkev
k+VBY9yLvYDu+xUn+zUQQEsp0eHMOKb1/Bl5lkD0xI0frAi6N79lEPVHZgVSVgJWfy566/fEMKd0
PNaH23fJWqmOUxMXbfFcUnPTysBBTWIxAv6uLNzWQ2xtUhdUsx4Mj+A1VMwIe0xG9R5Fb45WhC0Y
CmyONBXdwJ1tV7Jqj8m6LAnTUokGVSWx8zFmlYeIm6aljVFd3TyzTpPal9Y7CPwUzDbFZO+mxdQ/
RTsQfHqqRwvMYH/fML14KYf+WWcWX6911gAbzUT2Us1mPVeYaEuXlBwyHlZaHl6PCn7tXhgreNAM
GvSONQ6C/sh8N/mkOuuiYvkgegXn8YwCj731rsabY7efxYiVjOtwRf/8bJltzs45sLuTJ6txR+9C
bqQnulWCLQrAQ4jH6rgbJ9yondSfscGGTBjfRK/rGkY8HT+2G/4UQ3+oLP7If9jTWSi/jFmMV65U
ZGmY5jsC1qKESIFfFBdJEOCO3ImWwnoDWfCuHELyS5fyCMc+q4bhyC7FpTGy54GiREKiZVZ8hp1K
WwBIZQBpS7mqXXRCiGdOdyBvoZV4T6RcNGli0G9mP4hgrrjsBOXsKDm9zW1Bef498xxG9PnmaRyn
dpkgowG3lNCCuF6xtV2PkP0RUaPnGeR0VFxz5lQNTPmVEdJDF6z9PdXpxkZwU0gpfEXUBjMVGdPM
7VJpmu5cqqFff7dxY3ims0o+c4Deo0rgckcaem6ZsNxOaKzj7DQS2yeCl1T3Ng4Ngj0yhc6G8ZEG
qSEjaJdY+M/YlRkj22RNw5ozKgx4zUNdUhWSNCMTdag763aIgyynNkOreXuKyceKgk/zaprmFZls
WaFlfmf8/KbiDMQTA0kW0bvPEPqQ90qAlprFnNzSQOBJXchY6V9BIC5rWTrDHu7OJIptsPGOv3Ay
DqjT1GU6lKYo+OcxEtedESCUr9/mb8U8FstFs4Nvy4yc9IZcpSB0CfioNPpKdeZVhU4UoGU9niDs
OgVsQ9o/w8sEEVqM3J37JNxpShXPI3hICACMkFy4ZUzUw73HpiRs596bnMIFQ+UgLjMCN4n2MLR/
Im+2D7FF+oG9Z6H0rFj1Tuql7mElz4DFwwkN4ijXzfOWWj09UPr8G80klCmYp2GjeGku4sRNSTBq
BKk3q9t9Di7H17wHbu1ZwE7n4hu5FAWfTEqj1jbKwecOkZxfUKa18bRw4KHapNOpAZ10BxkKREQO
EupGf4o9kY3lsu1WMw6OicO44vRDEoXrG3fN+1+6kgdEdGLMEmlbYL1DbZgm1c30PzI9MRYFfIbE
GP57D15G/HS31pb5ebfXJ7EmxLF1V40ftyK0HKClCiivAQM4Fqs5SQCSh8w4VWOSFDuBqafQ7Thp
jDQn/bzfOg5QOjWFYxl1MpfPbeK5CVNtqtt8WASR9yT6k5MAQYIo8GSPoXiBHSY6wyBQWFkImSNJ
ojT3VUhv6dD7TZCicCwYUXpMwIErYkREnIr7tcP9GeMWcyD1t4Eb3zj8R/VDfDIgqNNyyYzM8/+s
rCDY22PH+r8KZi9lxrzdKJSYK6TY2ZXcx9osOOipcpOOx0NYebArFRbvmaHKEC61TTWPW4GCt4g+
tnLQr9lAXN2zfpEDj5twKCZ/vFZh4WlP+V7w/QF/eKKyCFrUIYpK3PuUvAmynTCuY6j0ciB9UaWf
5UPv2PpyVI6/9MdJnRX8eSJGQBs2gV1T87H/OyVYPKjv5GJfVU6E76Lk6wYM2naFGf6exA8xmfeu
hPyyNeUznmWg8IY3u3LRqgp9Sj49Hl2RO0LYEd8y4CxNbIiRg1GQ8EZ1xaaVGeIKx03HxtwkwOWT
kZ5G47zKSmTvGEGQ1anFnU0mWc4ES5qkZVRRsVmKWCp2ZX+hUKkMGBN/jOmXOgtlWthUZLY/CaHP
LV6rGtPYWHFLYTU0kcHf9lKt584zuoMxtJEVXql+9AVFuw3q07+gf3CvPTJPdEuTEZBymIjy/Uz3
lr24VmJ42b5uNdr5GWb52Lpdq4VP8MAHPSA+UdtcKc4EwFtmyrytimhC/MecOii4hQQkiLspcw+o
+o1FHZ1Ev5Crf1B69Qunb+0+42zSvfyAB+8jxS06LQ+F8Qkwgvz68bBEvQKrXVIZu69L7gqJkoe2
rDygAalG932rbCTrOoF8kSt8vryMwVWbmlvhtbam/7/HmiQAZgavx3//Qwn5hPiMkz4gHt5l0SpS
Hchi6ot4v94xJg8XQkeMlG1cV2N4S6hoewgJYrmB+n0YnFmvcla3rwJB9rQfKklCJlazQKG47ayi
q6WC+tCSv/Zc4i1zkZy7oQRS2auYUMlJUH3SO+IffmBxyA+ViGKvP4WP1//LzuaNK6VqizM3nYvs
aSYsuBSe23FZUeh7iNTfGFVB9bYXrrfgNuCwUX9j2Rtpzn7EDfDKrpkjwZbI54S/6XyEWUAnnmaW
mkKWYGRicO/EdUmZdbgLYUYp/6F3rnjTb08PLFvtG2lAzHz1bJHgEGZAOuJilewUL4uXr9i7DaGJ
vsJPTCmknxHO/sf56SpuLVKngzd6cJWURmaUtA+tx1/U6skYEUjCLcDbP5YUsJqaW0YbOKn7hK7F
bV1O4reqYjnj4wHmwmhF/H5ktTN9ffghd9bIg1HEqfsimzilEDc2Wub7/UnolE8wCbgAYhhSkOPZ
UaftMzjJ6vGVUm1dgj8oYnwq6t2W0DLCIfL/ujMo8/DszbXeXgJfg8OqkqA+f1ar6w4C50xJLwnd
NlhzUuR5MpHaDFEjYfEBf6qPaJ3cnw3lreAxPeVSHjNLI/lsjO01JBfYZls/OLPHcch4Wb4Y0Qo5
LccCdkr/L1Wgy71hi6ACEvgSu+6oDQrdGpQGrFqaQFTVTh8Z1yw0tdm6oevWobghqhwJaGa7Qi2o
y6sTPS04lDmxG8DSUOVk+kZCQpjC3cWTMnuhpey2yOLfw8SKjb4R0b4CIezSfN3Wk+NPltvik0LI
G2j1eqk2+zHv+n8o+CYuvGDB356p2l/nKwn+krQAUQDzFbTm4gn/vK83+x3o2b2BHp/Qq7mRZgwE
7iM2aaIFIhSCzHn0oFIqSpvUjGEmZvkRpkzA0FhUqVihbZxwsVonywA6/scx7d861OAGbecQWnSf
bybEUQrbZsXmyS4PKKe9gR5GgpivvGPHtet7XT5BaG9iNjhaxtWXBMunz1lMqcIoXkAJTllKqCD1
qu3Kdu7CiOFaoe2klCF2hHno4xyK6dAuSW4HKTEQpvL/C36LUgE5ETfsb6/0uOI9LMXtnYsB3jlh
ceoLnceetjy3uqmozS1Hdhl1XcKr27yQg+Z0dBH2HU9rueIQh0cinkhOxqk8xFYn4p/6OTAiS/gN
2/IikquJtNZsXdlW0Kc5SYMEeSBBvtp5/TANRVWVa6WlyXHzqHJd1YG0add3tfGUHKomPs4SKh7U
aU8AIV679Zy1E9/xRRzs9ZJ2ea2bLpO3G6f2dMY0CgSCf4brPplpuo56P8aKrB8bQQnjlw88W4x7
a3gvP/FZSBC3m2vo2LNrBeUU5P5F4cY3szgK3gR5CczII8TJFN0mIkaJX1fH/kc8Xz7BnudwlQ+r
EilWUVDVCHDUp63BLan2QqBXLJUUaimrq2e0XG1Vo4AOM9fBsgtQh6+ofCQbv8UwhQeORrT5nlDq
WBC2yeaDSRtxNteDiW3djco0DzcQX0V2W/HtzDGtKhAp06NqBAfm6NM093QM8Tl350xQcor0qEL1
GNfg0JiBmqCLzmtm/SsT01DBkTRf4+oPzE0V243yoynn0E4Z5LW8cpmEDg5fpNQYpsMStTb99Fkb
U8o00GkI4ofMkVvAkbJoHlpuDlRAHhp1GTHnTtJzVnJfm1R6179m5DeWzq5OHOMxBvNTK3sRVXm7
+0rILV2a/fjCsI7wK3vz4fNJg91/2Wwea2sVW/gB4WVi9NprYn8G88huVtYHoK7YStCDSIP7Ebl7
YlM+l7VBnQjAeeppkHigVfI9Z81kBLRxr0DcN1oTwFVU01Xy9IKcltTV4lcJP9OYYmCD1zlSExdq
NyFM4L0+B5x5+5D5NMwWP73bUkfDALw9utsqDkGFqAOw2IIhTialQzEcg4f8n1FsB3uZ6Y8fxhPc
ZXnM+BBji3qKsnphoAko3F+LyO/7LTUe8UYcoVVX2lrQLXlx/3JvZgsvYvo2wzjbeyIpxErgkUyh
xuVcZ4kNKRgd906E04rT1Eco54V3JshkI0RmN8buVCTxdBHylSb4cQdLOi5yhnpUWqJkpu9e+GBm
y+GEm54yb2pIYoxRhOcgzIbV0TopNnPz2jumDPL+WqJQCZQCalRPf61WA4XaT78QYxR93gVkQYR/
IGTDZdL7RUT8FIUzbDMswow3dTSIq5BWk17N0JUb1aVc5dsEqQ5HYuOrJlIV9yDXEvrJWNDfRmRy
ZdZGiKLyqyL51Pww8QMuJmZSKNBqmuraSGM0d5wrNs1dl5l9wrntHE/+REJxTTMKx0zhPaXxfcQt
W+2FF2oZRps67RSaYx+lks99yZxxaCAOp1YI2gL/63kiWbegLdJUOGqpfnLFG30LLnX9rnR0itoS
7O4HlI8QU8Meml1TzvoJK1xehPivxrozRQXF/GKDdSJiSTBD+UkpVcZDBZl3HXUlQliKQBCZVhzl
J5knDv36/RkMPkdLwMThz9R8wgjdwDDpu8yWGjYdb+/VIvnbTVMHAWFgu9uK6bz3/maZq1V3Vl1H
F10ZXzHiea43XuKlJssPxR0SeahkUQ6PnsqMIFGvtfUu/xo7jzc/MzyCDR9rZkHp4VjSaDRZqWkH
uRQ8Gcil+pELX1Zt/3yzq0fg4GqBRynbWC0fyH2HnUoA5B5p+qbCku0uulNGpKO0Bh7hYF1W9x0j
D1hAc8wf1jgsAZwPqHyq5iIj1cQMK7nSki+lKdJttjwGPFpnPUNUunZ1XQ+hYlS0LzOE6DOXV20T
PuKLQUUvEW2kb4RsKMJ0EgoJyHiC94p/wWp08kkp7Y2eFe8Fejji1/JZRBcfwLn2mI7y17yzoWrb
knbgbOZXIoy/qJ15/Lk2BnfrWZCWNOr0gQQYQYwSJeBdqiO2+xUXSZtIwddI5COqpZOrJmnAQJze
cuZ2SQoK5rkroeXW0fFj1bWFEVVINQW0DbT3pnW4LSMGQr/EJ+fSvMQ8XV/eWFvxt3tcd5sCPS25
o0hN/cZEVNQrbfq1CptQI3GQsTAMN64bLdWVCJXqPCKKghi+qQKEmvzLwvPyc14ab3qoUsUglIQm
b8+3pPbYcHU7ZpkEFNWANvDZueLKnk72R+8OLNbk6AxINqQ44JzJMUieYvh9qGLmLhlPoaPg4z1Y
LulXsGfWvA2npv5OIxrHCH3EHndnXzyC0dQCznbPuG9oPidq8nvNudLMZ2tUiNdHaeCFkBiGlOnv
zyxs+WFE0VYefuoqBXC7L8RnK0B/2w8E1YKYGsmhvn6OMkqMoNtBnJHisaWQP6Y3EbkID+TsOlUf
3zZP/395zti601/9d0cAT+POvQEhyDAX4bX0a1Gm1Y4qjPYhszGt02367kqeqdr4jR3rVysz4sts
IYRSRRdpSkQRpnD40B2+eCwIbEXeiEWj6Da+JgYtX5XSWlgtpZDIZyNiSKUN12x73VIFHKrfVOCS
jf5TARpH04k6MyU6x1/lcbgonbXEEWy/TVVbAgccStfMSBBSMQdcOijZGjkl5rO4LRnCXIPnPzWD
isknxz1Fwl/2xt6JZG3jk1IM8j+Gp6LjERIdp2tJ1w61F90UVTr08mfvT2tgoFm6OtlRwrcu5Y9l
C4cXLZZTrD9JgSdkOXTTAgvTLsBmNVDIjsFv7hWPIIXH2iVnS/1+nnSXa6Z0Bau306ozqeK05KaI
Ktd466Qm6kC+k+g2192Esr6LGCMKsfhDvG1/Lwxi0spOLHvQ7j9CjvEmOCyL35NqFiV+H13GUZBd
pCs+B+WbaXVVmSH77eaBYbrb9N2oVb/BxxTbliZicXFDvwphbnbAlU7700QkQDYnYl5KDD8DgbtG
ZZPlxaj0ZCBIFiexXitQdB7RpXIJQi6UMy7fYAIB34/zU8doH7yYujfk78pWrjjIGYxcmrRBBfjX
Ef2U933IKDYzqoKp/izTJQS+kb3ffYAiHk54+NxQIyGysA9pPylb0v5eRiBoTJWMvAQZvh3LPVFP
Ebqln3/9YacUdu1dZtc7gvJyGYRRTGsJWduHRAZYDZgAN8kKroEtuBOPX/8Yp/gTKcsavlk8q6TD
rMaOE+yclgdUZb1Ae7FSiTHye4OexKQTEQn9YDhYM1COFUZTsb7KDyrYxCioSprPZTzfjkRCVgGx
1m49uNWgKoq6hysRMo+wMDpxrLRmPOrJeZOno9Auesr/MNGMp4kXyvN6BFGJclQcVO4DGyeqb8N0
knZ/LC2Zd523VUTzmLQX8UCI0RmzX1pgv8o2Ir43ZSLDNL8Rdu0OsT6RufUe7qvB0G4fnaz1rbM9
eJ1jK5CA7eGa5lOOsMlC4gz98jGOj3rjyaLB7fxtqOQEJnYaY6IglLEyK24QRUKNoFRqS6TRXrdB
DPG5UVjZ6VSlEgWWdSW0Edq6/x8pQB0BxPdLuA4rKjIPCzoLw6froni8K72/ZJKlgSFoxsdfx+z6
EoW/Q3y3j00ri/bZ4gosr8/jKHIXoFtO+oKUFMMMXUDa0+cx/3y0A3nKZeN1t/8MXDftmRYTTmtB
wtbzaxrBvi2zLVOdthchnJGXOOdISH+ioh5/70B5Wj/G+b5jn7Btvc5WcLGcJsjqSHzpIXHpEP5f
/ojPqjvMDjr86OB9ko9cMn34qTN0RRtQbwBStCg5mamObj53l3I/5Kx5ZBINYut+5NMrh1MXhdSb
buvG/fz2pZB1q/qtfYzzu3MmAceJZ1fsIkIv4znX9QEiooWkmUi0Iicj1b1IVbF2hryJv4OoPhHZ
5damAUBLdKJNM6x+CiRypONwmJzz3P2pLbsrpqrMoULbbft0dLKZ79SVEVLmSyew3DF0aEmtE+U2
rxlQPNnVFr8FizMLaIQlSocwOEK5LrAUtqDB+IuZMLHVq+95SzrZRoFc+J7mOcG2jeb4Oy9GVz4b
Sotabi4A7N3hMC5QCeij+4W8kvdOUJsFFlQ7RBfgKLFP9TR4CKYsziu74JOqMpYdINtWyr2tT5vp
ax30qLMwDt6AQqMRNOXT+4cROJMM6EHfUI1mkTYnPH1unHsQvPC7FiOoZsd7Nge6Km1mXK+iHI5w
qkWZLE2lVg1cvXBX33FSDmdN5s/aa3gelOLn+/2ohGgLtnD2fRwqmXKck/i+NePvuGyioeN0RORN
QDX9fe0m8zGwlBkL5EziBV9iya68jZUP315nyWWzCzdZyjYZkcg610fi0pBSEjkTM3v0+wQ01+IH
pXn18EvkS5AP3ruy1GdCSa7zWnJ0sW9X7UWdgKNc3YAKEAHBtIH6B4BiCHR9BsutkuP/EW8rugbR
v9i3cUqpkbq0nxiwY3qVRYdHKQ5WtiKHiKi29UTJMInYp6VdwNWdCeNDmEzse0nBSf/TO2uosHt+
z5JieUNSfiCdA4FALSI3+Ym/GTuDI+nyc6GPilVYU4CECIBSidhGrhGDAMtAWA1mvcKK8tx/LEBj
QLpkM+Me936yJ5Ps9VXZjyQHHFiPP14IzySVprpwRRzqT17VhBcOqMAh8jciINFTRPLq+/rLYURi
ufrkZIj2442/aduzTnYQp5YaIK2Abg1V05ZsI/DvOwJqbgCAmwQhuoshFnv0nfa1yoqv8DEbc0y3
bVIRt9HUYyc+h9QNQm4h+vjJWKJDnFtbHM61r468OmfogYRbKLiKw14aN326snMjo51QpL1CBlw1
ksb7horb2ERF+aAlzQT1PBQcZSckQM2Q8EouDvdEowze0Rr+Rm4Qjwe8b4iDmI6c0W4+/nn4rBgd
GJXL3nNHU02NnAIlYoVFyOzYBul3SWdPJfS7hRqeAn7SFs9V2eutVooDN8TnAOKGlahAGbz6Dg6y
WDyQTfVDlE+rIMoLxAVYdC5kU5CvM2gKbDo/ppJpKW8vFoPiWQuynk81WfHkdEsNIcsYVXQ9/bLs
rWiTWO/+v9z4dI8+A22+mMYYzioKY9X4oPYhajIyuKxQtWP2sYp4jZpU0RNNHeHYwVTuYfnWVjsN
MI3eH0W19qzsphd1f4kTf/cM3Bey+uFk9vUEFXLMInf4PqSbP6TRddkMEltRL0dCFZPpVSEt/AAB
HlR8GhpvwRojEcvdkZekIaFN7oylDa/bLznwUbzS9CnD2WMpYGFOH68hHRB3RsDE+yWGUmBxcrXE
FGhxmzALDA898VqWtdArS4bKT7V/af/k2105C0mPmBF2Gr6f3zz26Ric8+YGE1atX5JmN1ssfU5O
XseR2qSwRAhgMPSrhYNvi1EmrjSFkYmJwmrrydqseSPok0jMTxlUkzBj2hLf6uAvLCgHagcQSQQs
s+7Yf4zm8ldVihQWF11Ahdcz1m+dBbZf3ipbOEoQiMK1IAStosM2DU8+Imh4Ads4+teiJqXSHyZi
QbetzoHbVvWEYljgFNTeI2REBUqa1yHjABoZ/uthgXO6Dqhduwc15fiSBHlooUQMpkM7nfOxfC86
/Gf//eKop0TwJGqScgraR8cydBbWHvzIn/3it+4MZxLZRlLk+0iI2JKMQ0amduVOXOlTp636KXSn
JhslVe1Hvlmzf1+gunsJSLIRFQyL9KZU+GAvW/+MmE3tJrVfY3fUrMgQEqh13+mpvlK1YkCcbrLv
95FqPUPDL4Mh+13KyNaIoRKEuhCTOPDS5IlGfaw0Vmj5ffZ+tzBBBv5J/vDaNMtrWTMznHVbN8km
FVSkExM/0nkO+ScBT6VDumVqxD3awKXDZSEHMax4TGk84vRPFEHcdU48TsrpHNmoBfN0sDnSU+Bl
kf+PK5rEgYGtpvqH5C5B8pF4hq6YaxkhQU+kcL4bMo5uBcJXcdyfGVYpS0qLwsSK3AycyKiV2Vbw
2YhvArjF6QaylBwOjzkVUsCi5Zy5DsNy1x6XdKwN/zRzsPkp889QTU9mjMbmRgfNYewafc7zoHds
k7FUsXsY/KHqcaPwtiC+JArdp1TQGHfSWIzWxCTUSWWDADDuh883k+v3F51BfgsLk8AfgO30oOEb
A9+56gIVcesBfN8eiRqoXLbY4Y4nXW4iEGFfIrUZzSIdrxk7C0dM0XS6cjU7oWFsQU86YetU1YEB
aCeDl+/lJeUYFtdWubDinLblgGqFHuuSUcqCu9N2NxI1lrYyRtliY5x3dRi7H5Eoi9szzx9h+5sp
yFx4+PdV/TveTzhyXILP1XZ18E13mvjyv5cFK940JF8a+PBE/Qz1sw/8vPmWgwiUctSzeTLRWU4B
K138DQDWU/oQQ46m2WPCqekpC9eWp+uVYb3M7jQLXKoSO8JKUN1EYFbQ4sIFkGbBkprAGHxfJBw+
owSdiQfguWb85xt4L+rgF9+FWBZJLtTLoi0BE7MsNYMlpjrPbGw4fMD62SDRXUJ3+/6D3xc0dGbk
oNwFSwAg+IqOKlLk/eOUSXUrGOhEIsvjg1YJ5UmbeXVho2BfY8ULfekL2VzpBpbvnj7Zi66E8dA2
Bss25ZkPGA4OBlCeSL9VLvbK6yxOr3NL9X1L4KZ5tQm+4RHwJJgPk2XrjGAAjBPBRzlEIZZSsPIX
VXN0WyP2sotrYRUoXUjbTYNj23dzjX41Dv3O7o+vb9cqTZW2MNakxoRlTUTAR9sgQ0jgggr6fmwc
tmV17GdyNqQGYvd/REFV/UF5Ww8wY7FYqp7YHa10gUETC6SXc2Nwsw1cdi+8iTT5W5yDuSJXOBqs
KRYvgRajNX+uWoFTU0G+p/McGgmxIdBSMeETW+HRu514aFDXIY8WOKYP5UjXbkrO43EKX/Tm/1f+
u781iKQSBLOOD3XLFe0JZLSDQYFw/XvdGkgZNhBwjW239FlkTsyN6UiUOEinly5qpbOlYOlAeeB1
J3jlseZzDn9oxTiS2XqiBmBBWUzWlydzqTnxvDmZyubC5BnQTibewpcg+Ik7a0xKan1N46Fkhq1n
NjyvXh6nOWHQPbon5RjiKOu+HRh5FG5Xrt3NA8PYXmrTdVJxoVxtYDvMLhEu18pIefZ5Djxk7Q0d
+AtA0ENfAXjsYMHTW7EFkA+2vwP6/zKAhcCOSZtB7JBpdtjbYGt6IDv9dgq846KLwzBWoAfRCfd9
dtgGyuavTyVg62GGEwDJmsFup+HVC6P8Z8nQXF2T3jaO6jJF02GyrMRoYcGEe2driMrL7K90+2w+
sy/Rr8twQ3VIWECjVFtk4O3NBehrxMx7Umt8HpNQa2ex3+ksSF106NugPBmm8eT7TllGuWbaJdUt
vMfPAvKv6dC7ns+YunMsZjuHyPHKVp1tWZztseEidNEdz6XL0BkQBLEO8EpVVt5WOXv1GNKToh3U
nKeT90jPm7GLIXd214QbkdIREGsgyYdlZRCiMnFjN/t6VFgxN58hYN659nIYtwdhJ+5aoVaOYmpd
aSpr9Dogb8WveTQTtlxiKQi24pOmw4jLF0OLvPW0Y++K20toBs4051hgf7+Tbp/yskbqX6WFY+W2
yCI1bVafdwu1nhMWIbXMMdMs7bWRzNnoTk86xr4X4ODXMtm0ewENaOoJK4qa/OiNleV8c3mCyDg8
eA3du+xtjUeXBS1cw34Tvwob6aQ7luJLATD9c+fYtUqJePO8RKwd+DTnolv7ljJbkIivzhJuHSJG
dYMhDDpxycLgQ6TV88K5pe5xvX5e9xHiNIPBPJl18Qzsr1YVQCKjfoCwS0/eQ4FMLF7uwpfUAFWL
jWYixixTNpsrfTFRrdimkdJUO75sMhPcpt/2AQhtNAdp1WS5v64YdJb9KuOEfTRW/QPo1P/YdlvF
Z22qYKPCW+xIvdaq1++0Pv3bkleOwrbjX58kJ+YaBcg2IPHczM6P2TPfB7+nnQZwo1XNNPElvqcK
+oQQt22o10g4WVMrRmnLnlNnJsiN908RDArpqnF1iYzTGF79cF6zkI77gUjNMhUICJBJyO1JXnfV
FCNI6OnQBBGTJhO3wQs6PufuEZBYojfj6eUXZdsD8aFmRme/pJZaHFGb9rthW7i8xWLc4yx2SKqe
otQAr0Hk5tIJMvr0JxRxmvpj/xj72ZjGc6+VPwwf1r5rGP/s7WhRN64uH8i6hoPkiKQnyUswC9Nu
JRqZGDCfDhykLTEdLKZYAfFkwSgvBji6YLDm/bze+eJKQnAi0mxutHKbZ/3h5QV21UagPmbUmsTB
9jWKLtwcOALXI9qyxTrGnmlg+kNcMqIqZ2kF6r3+lecf34yMlPxC9IKyEje1F/z4TqK+RpYnPUEm
SzMecxbyHM89Wp3txuDDbRUaawF5aE1J+erugDheGQoqlCbP+QXEiS0XlpCFQUbyQhIcm7AneasV
okVASQ1Ew9UX0vNDlE1Z/iW1+GuuAJR3CFBrAm9KxAOrc9IwTBGkMkQBgSTEPITj+dNlajLQWbQY
9bcolMbHgTS3YahoVcn7gsl39IDjHXwF7U3NohGqjQRtFrnI/9rLElEfnhS7ws+NLNUtsQZgDyZn
eFttiuYTlR5t7Ru+o5Q7HyQ24rXAUXWGZ6MJUKhu+pg7J8G7O6jyFI/+M/2e5eB3l+ZX+e6U/u95
phw0+wDE00GQM+UYPGa4ntE58LPpNxyGVaGkJ+4iCc0aPucQqBsalA1rTIHz9+lh+38t5hVIyZeD
YVndo+LpsFTV5magLaQOalMlaPY6MENUA1gGngkM3bJRhjHOY2VPb2P63/WwHXuLTMNjP4OruvIA
ga4xoYCwJzyNbHr+aDmVMNE9629BQMUnuhW0u59QaBFpvqIkhXwOhZcRQkIJkn7tx3Z68mu87sO4
kOGmOizP5ta2kEW4fL0tPutHbhjg3MiAlAgNvR+plxMvFIwUyFSObTrZhz5sHNw7dZDpRrlZOkAt
TF+7Ixw3nK+bXVfhbxPg7jBGr4Wc6YBVR3tAx+t1kwRZe25ti7PoZc1LX7qgtii9VrG8apmvhwep
rVoje+hMFzdRX4R74OeRpX5QP9QEr79/jMRhpQfeCF6eSpmxe4J8D58sk3uBY2vmlCYP4bnKrAw3
vxDurFTgHFk8VDhQHlZZkiga7lkZEitThPGjNCcCRCJcMAeXimWMlEBT/t8/82rLih95IsnfH65X
n7rk7a5xKa6aOFKS9n1K96sIiwGGm1Akm61GAAm9p5/abpYNQATeBmNBQtCWFYGPsJ7uFMP3hnc8
+OwCq+pH7nM3rjhxJd68hCSFvuH6B373DlL/T0IiABjxIk8wtRmD58ywANKNgM+vvuxW1l4wH6OE
D4Ta1gNjILU8hX5F2zLbRi2ke41qCLXUVleOXyYDDF0yfNltilOkkU29Skha2k2xTu5PBsaaepHY
9xdA9J1SmriKOtYj1xigWeCA2JbbrYYB7CW6UxXgO96NMY4MtxLqAlN1FdFa9o7aKxVcy19zEEJZ
XXvHZY7epHD9yIW0VHkfzkdI+TRJp3EMT4KPURgQzwwZrIpiNtAgX2IGpjBP6EmE6lBw7Y4R1600
ctujDlSKZxM+WfTdBPM4zSXOHAbKkMbK5LMV6GKMIi7K0AjWzIs1EXXkMzgxbzcoqb9hKUnqXWdT
TW8CGq4jfwgXu1URX7Zmz2o/+kh3UBBAIZH1tywDx/sSqn+SVomXQrS+nc2i5HXMY/7Fu393vV1O
JZ4nXp6dIHjsSBoEnPkTh1IRQEsO9Wa+9hdRbtUjNlPMeAV6KAzzkctspJH2esbZR5IizJaCRgqE
YGrFvt3c/oWeWDMz1QRoqr+4JkEBhiHjPWIUughb/bwhXbqKGyg8NzTWT1M492awiD1t4zTRd9PD
kvGKun7MngDkmbbZqM4n7TpQqAJJpjVAbUxqGK+ACC8qND1BwJcDtfeFghwVMKKtythd9ltXHJ6U
8aLD4W8bTF3/+yMzao4df3IFaUR2qSl0x8sJMWQAejdUFawKnZRoO9gNJHWBV+5p1/+ObC6oOwAW
/4kYrNecekyCHZakovG0c2qFX0MP8nRD8JmP292q/CdT0vHEbQlJ3K5R4IC/yY+7r9rsnCOcxYLf
IdLppgaW39hXqtVyldAeZGzlt2gONdFtp0bCkwSeamQXL7DYslLlgClOFJeRTI2berVBMrbLDJ6+
ygkI/b6pOktqQsPfZ//aJ1B8QGnXIsiF2MINlkppTvlN6cZf6kziqHF6K1wlztGVBIenog68Pm98
fyQcsjwVrO2Dh/Eo1KDEdIGrF29AdpOh1mahIowVSfzmuDiS+ZG/QHhR6kAE7XA/zHADZAsEnET5
NFbRb9WnFxZMoYigaWppsUkUSuYx0uBCa8hVZkopwU2XFv+tNDWzKA4yM6nsFpaVKvHCuD2zW1ES
HsFbEk+wzVkEtjcN17KyBcjG8GlTDMqZ+dBfawdX07N7HwoefjRO/tpMzjPOBUVnRxvE02GOdqg7
yOJo2QJMBLdYKwVCbIFL7evqqv+9uWwvXzhwcM4XFhDqDqrw4oxbK30W2hWzibWhb4cTUJlZ47al
eALgPI7/duBKGxHp79phWqirN+yaBiTVMXeBfXuiogupMxKuO/Syrp3HAC4OdI0+zNHlmIkG/bvz
sbb9ZuugOYrdtbhKeFnOkBozeaK57pNjKJ/tpVjfzZpQSjaPOZMHFMn7s7tN/cZE5Tbo+2Tdf8RW
NiIjQZpgO26Z+RWvqAxnbXsqkNkPIU7my5UVaFhpVEJ92FtRDkQQNK670FVDsgdalJHGRsl9AVLU
qPdg/+N47mQsQG2lxyAMl2PBihhwpPF5tio9MNiNR3xnwEn4ea3vjMHYgV7LsZzQuu8CkNRrTA1X
kkMfmx/gHoxoDY8WS1U5mquD+CrC2SVpxMZyB7A8U99pXYjTEO4Mhcwua/2Dwr/YIJ2L1y4TI/A0
sTakMFmcuS+hvpVZ2/g+GeOuCAOoq5pvGusU9UCIwwiWaRATZlpEH0zqwG0aQHT1WBRafxdHQvBr
j3SDw3eXyp/UjGanNgztBiGyer6Z+YNEWVDJu94wnHmaxTEzdBFrN3o5mkmJAsCvQFBXfKUWCZsn
mekBNFgkTj940lH1aDNJEu5FDUH6cpxbB3871LJe41G54Vl0tcJGmNq1hVRb4lsFo4gkhya1bg1z
crp3hVkyNEldew9L4QcNyQti8bDNpJoFZEILm6CfKPa5uu0Cc3i+csUCNyHBB+aKrQm0Fq47bmLe
ABsOR3FPWBIHMMdgFiWiCVz+JKfX+0Llpeam/Jy6qzFk7XbCOrT6nhyCbjp9MrkHlJWIm0Vw34AZ
3FrcMNNYT+wvKOfPdEwUNwOh84hCdlsmD1m2RkbYiE6ZocmT/5qRrAhU/6t0CRDF5ElaElLkjYig
5nCXs/gZE2QIMFpF6bIAsDIYuOOD4WL16QNOqbDp5j3LNf20SJBiTOeINEqBvPNMqjGsBX/tmN7z
8ihK+nuhOxihj5jpiS3FvRLleV/bfnOrvGxdC1rc+iGrPYrG7+z15w9twWsBO2SXWVzGAPe4crQv
r7x4aIgljnmF7I7pMADQiSrm1C/y6ookzuKSE+xFqPAFwk6uy6RuU1AgVFCYg4zgwrl3bhdJd0jp
pMn/i0OZ6vtGBbbYUilpFVeaIimZ/C/G8Ue1M5FW5SERf1qUw4qjQ6KDNFtFCbD4ocuWen7VmWx4
0zDhH1IQUgnZF3lcyCAZEKARUP/5bBXWLynthcrY5R58SsrvK31q90KKDc6NzRWp+tutZ5Lo90Br
FiK8GFlJilmC37NZ8SzkKGMQDyTZ+c5rdgLQxaYquWnRZ/bq7PRqm0R2BZ//g7A7bi9kLSC3RCy1
BsbAgQJFLO/oRlrSJ8ZFg62ETAvh81E9N4RkLD9ZPG0Wd/20gz6VFGlmilKaSA/4NwoJkH3MiaO3
j2cCh2MOgZjlmnNau3UmUvOrtS1Pg90n1Q6v8mC+3jcd+eSjXQSeG8DT+435y7GMTc3NU3giDm9C
BaUkM+k0BivXXuq/SUSvJjbO6Q3mlg/BZ1L6T4+uIzKzxIHpEy300QI92ihmfX2n6iVsWcS/1oMQ
xzFt4kV2eRYeWeuau5ILWXOv+/dEsjii2jJfnhiTjJu7fuAt+4sQHpza3ZiJcMONfHrS4gjMXKob
V8XuR/xkbESa2VG91m2FbeLJvHpkH2zwZHlM/6hZlqi5cYRz6jFchVsMLyJfFNQxiMXO0aiuhTRR
k2hDc/PmO3jMAcm4ga+/+b0kAh+FG1qUQVDEHCR+gvCWrYEWrkmhFbtoeNkfU0juIY9ncRrdnyxs
6Wa7oXlnkKV9bd5nCSjfwP+PVeqgK98h6INxsvg7SsxeOoBmSiDjOY+lQ5XDxdV6pPPsNBHROK9U
304BUhqbrqKt396cSfjaZTLWxBgiQ1eIk9Jr8Eb+rfCLf6sMsNlWlMRTnS7EhjJCGekhoANWmDnL
HbhQehu1Sn+HQSHreJF1u3glP1t1d9oUGBGUA2pM1ZKnovZZ91I8XqNnQFzyaYczE8FBUs/NpXrY
KDefIoPbAuGapAzlWsPlmaUno1I59OYM552nwQtchdo2PLoc0phsqXEX+fDYdzgrkOIcTZAxlUcy
MUF8woLuXEscCsx7hJM5uHTmCM/shwdwGI/0H5s833jkdHvou0zFGvxbPk5RTCcBHl6bmzwJCVzt
zp5dQf6z+Mr47T4HEhz3P8zj916YZyAfo1PffV5gK28bu9SQHVgyUDcjIHn2zyqnYx2NoD1UvuDA
U+Y8qpjPWRuQfaXYn2s7NIjmRX9kvt1S9tIL23Oa8+8GZJ058SvXVIMT3TC04OoMQmzlB/Fgaiz0
pfwamWmDtRaJLBmOPNJCofX41adfQMxg55i9/hhk+FZYCbt8UppzFEFpfHt0m+eRDh+t/lMbBR7h
uKORKFsA0FWVJ7NO06qNB46UEtebPM5GbF5/Q2bK3m6F22FySFnAcTupBe5F5mKnXs5jkWM294lb
qSrr9hzxdD6GxGibIXNBHjtnNG3MPwTehGuim1tpD4qF34OoYXQoTBYC++Sspzkqj536Z53VexkL
N3Qrxla6LIiDYtxnDkHrLn+MoJhr+X3LgoqZLyUlVlRzrq56oaSL0HEV+KIqomII9mBOmlGZhCNi
4zzsELVpdEWNCmYEKvkr97QIYZLGg+46Dtz57dGjysYSmvQlfyCsjrDKl32XuW+9cQo6tUC2wc8e
mhALW7sRW+3SZtktInGxblfFhqdqid8cm6vHSjcEfpKH6cLkWc3FXLTUrC6s2waesrkgQKH4AT7O
AyPnbM1Hw4lh71ECWT18Af+W6KMRKAKFISOmZVqU1IFQmNbYAVBrMpBwH2gZFaqij63VPV1lSooW
ssBikpcp51f2xxX6F5ZOOupnsMF4/N0R5Grzy3xnc/JMmH8dvtvYcJSbNaOA45q5QD28ImS9yX0Y
OD9ynM9wQ31PtZ2EhWBpRakNu1XgOPVib8daz0xZal2yaYOMKJjYVH0evhgZOv1KtsiwsGRuMYSu
0BZA9D2QN8RSL3leqJ9lg/0qc01O1ulYde+VxZ7jICiMkjH9kmFo6aSLACQGj5mZxWac5rkp1Wkw
HbWJM2/aVJZ1VRtxRjcxQWa9Zohjffc3kouRyy2Ac17MEP4gWsOV8UVUmSZwmbe8QnHhe59kmKFL
TC8CL9BO65y4pkgiMWoFMKshTN6p15GEEWwM4EajTUiDTmsrBXjmZoQYUc7T0H6XsuU3/MyeCo3E
bnhtMTScfpiM3KOCgrr47VCzXUIpRR0KGj6xAoudx9h/Z1Ulvocgj/zyFUTsp6CfTNy7Uzdv+AtA
1uShlebwR3QQZXwXeOhj92KjHudFeQBfT3KdExLYYy4BeObX6jmIcIALBqYXRHwIQUXTJwT4Flbn
BZpzNR0R/xMCAi7hPPjzEMUY5SEfB9UpZbp/58JKFYhtu00Ji9/55fWCsBnLoFiYmLb/0odmMjdD
HTTAjHzEPOXwW1VyJa/CAUKXGn5fKMLnsRg7E2qhclO5VsUPJ9KktbWBxR/SDTGsr/BmLiqw757T
jJb6xQWD9UGh41m/j8SWZOxb7ESQTTaYFUpB3Rq4MNIsEDcxxswqpVNZbapAmKQVFjxyBgYePJ9U
vN5ppgYDwKy6kTEspYJXEfcrnXHQtpBQckfIqISLefF/FrzQIEhtAOy1FC+7lCJTDYU8+yth+NGA
bJwoe0zaLZaYEGhhyQyNwLIeldLIuju74utxGu2Gm5W838Lu1PivzprBfoRyDQBU/v6FS6TJyPyK
syLQJhLS0GKFK5P2D93i3tZzP7/LsCfjhWFMooMgZwqmdho9nqPrIGKbWb2dGjENef/9RGQVF5FS
D0r4CGtoZ2sohs+hoC4qZcBGp+Le6rFQoLaO5rwDMllIc7sO/Tn1d1jUQjBfEeDMs8qnXYoJHmv3
ganGVq4+kqYodSq2zsRfUQ0Df0YgIlsaRhmOS7N5rxZqwPEPf7gK7z1AwkFtI8h+B2atjS/Z3uFU
sw+/0Norsfa63SxIwSYJix19JdCulb+lF+OaKJWP03ICrnRzLUdP67WDwmdPmNa9XXAMmQhGfTSE
qE9jG7l0iQfBdsme75YZ3QreLeos2OZbXwlqxPvBNspt0IzzO6vs7OhgZiz9937KydlW2Yff8UBD
W2Q3Joa8E1+KynMvC3WLqyIYJjXIKrUjC9zIck+B2697Q4/F5jeyO+4nRdQzmIaxM/6+wXHbEzDO
c4tV1bmWMMQbPsrRqW8Dz6BvarJ9FaUyV5cYBER7vpGMHQa2DdFEjHhRZZzA/1sQvPdNUKko9ran
1PBSF7X5ck0xYkYPpS1CMrrwJYVvDlUN46BhTVrC22bagYP4Iv96Xj0ZzQ1hm2vwR+OVOhEn1/SX
MfhkmhxtXOqKxk7ujh6GUnepbtEyzhJYQZGqy5uCDpTJyzRLxuMJJ0QME43kRacTRWJIaMvJAPHk
DlTD+rz+9PvY2jm4eKEy07HXmQr8f+tqOouHhYRgLEswAUaUnHQmYa+JgnmBZ7ZpKMTzLn0o7x22
0FvHUbQ75TkSf6RvCTTNY6vnjDsRPfar4NhdgK4J2egcjDUZ4a00xsdTNl6RSNybhrHkztJicNCu
Yv/U6YQBZnQ9dMg+BQ/Sgxf6gN7FuphSI2qCyo//comn830K9sUH6vJIuLGyyUjS4PYfOQRcw1LU
pzyLlMEJ26lECITwBu5nW3NCeJj3tOTmopmH6kbBz2bKCEuOO66LP+nLdtOPfT2Ke1Jy9sa6pst/
p0ZMEoQSsrKRITYD88eKzfHdnhDuLQmy0mM4p+e9iuOeno2MJYak684Pa36QCHp1xn6NXA/V9pTm
rIQhuBYSK6Dnv5tOjZF665JhSKaUrn1A6qwr4GddVJLaGFas9phHiaho2idYw4ZIFme15b3tTH+d
3IuGOGEdUZXVMNyF6bh/+gPAVrsb3jkkYWln+qq7fT2Vb2k2M4QkPve29GJDJBezGMJBEXBCP1L7
qCQdCKxh/Tmh04LoB9DgqBaDGpBLAMnqmkUyVAotGsnBY6cS1w73s1M5JhBHNOKQOhRi+M4oi85C
85J1IieTn67lrgPTqqsYGXRWFND6bNJnKR5c5VXbymxCa/rmnew21D58l72Tj5wh2Xs3DbjUWX2A
LvRJzeFUl6B+MPg+dkXCqaUXyLch6mkBv7Mm3WaNcvvAdCZBIZIPkB+2/L5JYfF+jJrhGA2svIkg
UdXNSurk5+Jj1tnmt9dnMyZYLgsUMmVrkQZP8QfUrq6iEN9t9mVUfHFVAMrQ5wvJE3HZRGfexUh+
rao3xvPHSaBG4pmflpYYlemOiaFdq1Ca96AHGICcTm720xG0SrgHSu6BVGb487OvjmFWy7OEQXar
uukH7wuPfSoAVzoLHZruXmjPFTiDDeWHGSuIMwBV+9JUaYrXDOBXwyZkppllk0JB09Jb657DAWZy
hKFTD7IsiHUvmmqaqb1c90bCbve+2LDQVALoEuRm/R5dcpZIVM5OlO0Kl9pYDa28/VZgOZUkzf9t
APqDOYT7pklHrTa29VBMGLUqZLQFCphOrR/6xIoZe0a58k09uIA9T6nx3GNrz0JTdm4lI/tO2Ydm
Nw6Fh+7jWpFWoFigePicBNAuw8dIgboDuy4SCXa4g97Ov0DUFsnMbx5zb4GlJAWt3CyUld447edy
/JqJZOWv+1mnIHtXT5UzEn39vagMWQmRt/ql/4ZF5ibJzQP0qacHwPoikV5uDE0sFwP+rwAFzsMx
e6nzpW3+ok0R0HwZ8wKTu6i2fQ1X79c3VAO6ox9fea45sqiY6G3mJndBqnkEkG811e4PJNKSJB9I
4B3HfysBc0cx1lHI0HjTYAqQxFIjJSjHqw8DV7umxRUwXJQj12R98/dbYtOXoDatYy3m+TmT81aY
AiwZbfguoE8VhqkFI447eJmImgScPZpiI4PP4EmZG1YCPx3ShSUppCwQX6xQjsQ3dMSKB43+jlhH
kJ065unKlCj4/cJhU1krGsgdLcMKf4g7v1Fvrv2F+5N8VYc9tAqP0roGQb8Fm2tkslBioHVbJ1U4
7Qq5/BXyk1M2VwexH7Zses0ZJoxo+PRzHGBvfCR6YtZpgmxgNv6ljM4L47Po0kitxA6S1jNC6BW7
gZfimDm3hG7VImWxoB+zFYYozseqZLOdEi08OGtkpZag0g8gJjXa8C/8/joGM1WuywXtq22JgArY
zVyWlHkoAXGagGfxh5ChBtOjGVlPjRbAtjNdFLotJJEW6MmoRdzKAaYjAvzznG72xSZ1axpR7UVr
KpyQJP9p/LqLK8A79N9VKeMEgbEKGzOPak/IJc1kb1+z3Y+XM9LJ/EczI3KYt/4CezJ+WU8Hv/0N
tM4634PfoDxgNw/kX9fw0sh4EiqdiBTQE1dSmS15eE0EzQMrBbGXG+Y2T0Rp8ngqe388KAD0buW7
VN//WAQYZQY8q92BuoK6Xh01XjjfinRVyrT5pb9ygqRwhuillqzykU28ZOt505MonnFLkIjYvX0B
21CHBbaJzKLwueqO6Vcl/Gsie5cfS8NY05LAA6tPNTbl8WKoYJ0ES0mearl3gxOjhj1NSFhcSD8C
XZptGHgud6faZvcj8scLBBk231yPNAkNCRG0AW09EW1NY0eqLLs3jxNq8Wly9y+ugqsA+qFJRpC3
WG/bAOQVG3y8xBaojvgowxcPNq05EVBmUtb2VvvNKWbyHEumXXX2lenDHuPM87jghHqHvscCHQ3B
9IwQftgyNnu9Yt8KAOoJInDu9J0oFqs8dZK8ASMN7L0Mr70CcVBHaT6nDrcL6Mtmexve2vhN2BQC
ID6Z+sMec//UHGRs20n5aAN0VPBQbtOh3IfdKNyIIj+Y0hEP79QLlW7x5EqxLRG7IxYR3Dy7okQP
rlvFRR3KnPBqvUGREXJX5gC7/qzDoLbv8NNE3UOadT3tJMV5Upc6gGY+IuaHWGWl3ejSftS80rfV
0j6jLMylUIFPFInEI6OJ6u3tFLyN808N9V/OvzeDpgytI/alQ0d5/XNU9pMZC5C5UILqUEk0jtkB
uJmhArQsoxJn2+hEuPigekfbExtNxfhw3HN01jHGsgT30/aqFGZbxzGb97fMMFykB9690qzw+jxM
5dZBrUMGuqWGOmSQ/Scm1gjuaWtGFmDsmdkNrOpztijGetrxQsAgu6UsjHwJyEGAOogGf0GClm31
4ATaxr8gHzBSJrnTcIPOi7IXty37ozLrVi0J1sR5gij//PxUrcoTUg+I5DUHUZ5cYbxbFy91i/l/
DK+dhrUaAO42QR8t0OhJnOODPbgge85Dgz2IMGTbIX0n+TciGXwHYHURnOlFwgUV0PrgsoQwcbP1
241oQGy4hhpw47DOnLmbW+DWFfnpwcjT7JemRvHzd25nMY7biQ88jZ4fg0xdIEfCZtRlQIzbOEo2
T2JleksGc5KAji9UxaaZZpZlVbwHI4cOVv+poUnlgYJhBIA6M3FkwKVj25YCDIa2Kua9q2VA1qFa
crU/5MuKE/v+Fby1CZDzo1uvvo7m3vUn1tvEhZaXc5a4EM9WHVit/3tNMbVTL40K5zaQ17r2hZmZ
7BxuMEgj9+dNPI1ElYwEH14tJ+OQy2Bz5Msomym874fnYLWhcjG+JcU3QA/tA6PBtVDrJBY7Eg5E
iEsm46jMocWubWJCEFU7zkAVmqU7IMg4vWnavkWkyjlhIIjg/yMvjwplv7T+HLoXCzEslvbxtfBh
rp/oII9XfYhws5ZKSNPlqaN7I+0qG1K6I/tSnDnOcARCSaTkN6KIG905nvZmYzmfizhOo/7Ivc8G
REVKeW5tzyoXJVG+gLjiGb7mF0kHGVeUbSoFrVbyyIt1dCZyGjbHYAgo8CjrbHWEHdiVVoM23hXw
kWKCngSeLvWS/lACQsKLxY2utm8QugUHl43g/drNvuItVxd41/65hMDATqTzTZ3r+XrG/i699KCG
lVu0OTDDGzxijtvLMVqslyc3hzq81yj0rIoPTyTguxtzqzTa/HnJyltkrGD2p7c2F1X6H2mhQRa7
WFqOa8+8vu9cMB9foSTO6aiW9j8OjBH/WOS/P5Q+vBHkD9jG+lLoJ+ktQbjCX/EoMR/rqKTfzKED
0lTo1i4uxgCapvBuearRTuoRrV0ho117vtzUj6jXEmoHd+a9sw+1xKPULwWi955/W1GfxSIq6Gvj
S8RGe8TJc65WD7bRjHjzuDVWol81tyD10N7d8MrQTNjegDxunnaG+oAx0Zd8Xu/fpvFl04k5PgXJ
3pDRJPYxAQoaZbVWLEe/E6/hPgCyZL95W/CNR+ZDucHpZDPUvY2DdUYoL/oXFxPqMjiwpxrxgRIg
Ddahek3tHf6GeXd3zm3Wp0FWOVs9oIf6AR80tJUNQNg7gpSUJWjCYS558Jcro7DoJX516IWBx7rh
xQF0myUXGIfK8rzWB2OinJnrpNkZzCMYvJ1v6b1R3W7esivo/x5ss2IYrRI9Ne8fu7uhhdlAdKA7
hOytHFLunJD4iaarXwBrX4BsNFxHl1bj3pX/YP/LAPymCkP/FE9Kd3UFFxua3kQHwdIFqe2twPIU
zKEyofY9AxRuhqeMfSCUFoEKFwzRZOnaNG0lgrH5yqxGQlLal7wCQcDX0hkyN5LnY1BFEQVinomB
iofw8EOwsIvbP62rflWmCPIH36Lo3l8EUT3Fw1qtITiXQfK0dmZxmfFvGrdUyWkW5bpqFV/vtsgJ
neOrw+Ns7TedNwwqc4p7H7VXAekGzsSDaliZbMAdpf6CXaAbtVOSgFMhBsZBgin3K9aD/jCSE9EE
MQMwMBNuH1rsZZ3GPIGre2XafGNYmZsk2uYBuTGCBB8FFzz2fjWlIH4I8nre2mB45PHE4Awnyq3c
tnr7+2Sga8FsQNMCkUx+KRpb/hvWapFjDOlPrYerbUPJ48hd+7psgZZBu0xAubOIhcMpFNSner/l
0ncJnYxCnW8OOJrz/NLgq1duuSYuTMH70tbJj6zbfgSmLeyYk548+WUNA4Lklw9+E/uEoue7UtTo
wCXYO6vRObXjFnciDKlH7RHnObxmH1EX7PF1j5/4TBQo0y66Slooc6K5vqOSWXLN/99A3NOjfGUx
+6Ya8QBj4G634WYQxywQTtD6pylNWcFRQdYV+XIYvs+nOOaOXjqW0w20HU0Zmcfe3m+5c/hIbEZ6
atSJvy5smNieZzz8xR/b4SC1BiRMT6P4lGydR/xCdeXOpyFCx76WC0KyCrnOsqUBzEM3xrxPmi4L
nuBJ0p/XIlvM05UhUXzVt3mjwJxuye5laDxTisqnP1OT33bN82N70tEqdAbAGuWFa890DLEbrfMb
WeaG7/RbEBNdzn5Rg8hy/tp1nAvLt/qbzJkgCibLvU/uCGubGgapxkZUJI45SKo71+9duLRoF/RM
z3vZNTTORUbgDHoZ2g9M7bOfY0kNwdvwCSV1bndbj4OoXsb9hRwL+NH2dRZTkkIzfHnK0O/szQI/
60OymUl7oYKmrDHr9UpD6RqRuXhmmf9ABbeEe0cqcRea5FuEvojdZowXWwYImZIjiNdu9DHOR7fz
3wvri3QPy4jbKG8z/k94H7vwJhXDaaSjKVy1YURtMyfwo+jpUtvJEVqDIDOh1hLXAZzLVAF3uTX7
jnufY2kVDxssomtL38j7F4ApPGPIE07wFH/qLgUVZFn2TuWLdPK67sZfUDgsMW8Td1fel1dzOe26
nq9/HW6xV8hoN995sPNElWuI1Nsud/MMdDYvxwYbUMqFs7wdgjrsnqTuOwyT0cNVpohGqnFlOYn3
VdFviNOmbKwalkQzAUQN6p9DeYh9ws/+FuRosnyq0Bnr4b0qYfbdDRjx3PAZBwkXC/v6IxThN1ND
LtcCJgvZMajKcN/yoE5agOaYHOSPLLATwtR5LLMuxvADBWS1/4qgU2Y6OqIgIuN4m7W05cP3R/4Q
uFWIp5ZaasnnrV/Oth4bxYwwow7qoyKbJGJbiNYkdscddIF4srVYpLfzH6+Dgb/V5m5MiE8PIupA
anuPdCulFUOxWOt7j+7cPmvLGK9jrm6zvLmGe3vRSPa3Q0v3HxpCszeaNkDUzr0xJR5jtEv9HD7m
Y72jJteCjqBcRWBA3y0WR7BQtcLNJ+Pbsm9zYdKHuOHzS+5rz09wz71rf+Xxll2wvzchVJbgexh4
T1UfDKfeEiNPNkTUQWjePvq3ktKnULWtRcaSXsfx10za6tNKbsUQeBPh8da2jS9yQu8hbE97bjcE
bjLQNgPbQ+4RHn9aghX26QITyY50FAu2FPJCzJTIs9te/FVuCjfXzYfuHuhPA9DdB84g5rU/fZdc
rc4Q66uyU9P6Ax8bNc3LJCTETZ3Nj3qWRDAghM5lS/+A/JZb3lAodNHeO8zpVsbQbeLMKMcZ6QgE
jtSBGpR5eJgK+zOV2SqN7anU5vRrurAvrt8tX2UO6+m+WAtVFj5latvf6IZMgl3pIYb7+sLNfZFC
ZQM4lfoWrS0gRpGQg8t2no2enRhXRwISZ5jBUqpkwH+tGeldrFMTwIaCVJidkJ+m8/Ic/M6Hduxo
lMkwDwuEvlS3yadZCG0Lyg1H1eEdo29cCz0lAZx8JclNcVzSLHW+VsprvMMRYZpyLiBMe5eiSYu6
cYqneFtr7cRJCU23xFo+hAXcVBWALiY/y0+o6vgT4xqDHF952hC06fG5nu+xnh/zP3bQuwnbxczs
S6B+k6RroZKNoIeGpaVJfzHi4kWb3jitywGWO5qrbDjgIQ61HwBnUZXRWSHB8p2E9NxghAw7aZY8
f3BPYAYODoDFOTJ9oSKqO57FPbSV5C6F5XW0QDGDv4XuXZqwBqQaJ76qi5pUB7skS+qQldRLYZsa
nZxQEpkumuWpf2j3sOS9mQVPTZzSygYz+5rnUBexA75Py39Hfb3sneHC0vydtCJjsJclZHOnzgsd
uOEPyIXr4sWIyqeHd+25JDsXSUreS+2OXzg7HAj0Z7VrM2zXlnsQ/oJvgFSRKC+UJWH4bE8VQ00/
E3Zv790XAXZs0zerEpyFCT65PwmIVosv2I6LXadEoaWTtnFmj/eE7TV5fehPujnBwuyRyb1kvWYT
9jlXHLp8oPSLelUr+9yKSCjted3oszFm9TcYFfCVU7Zql40+syoLPYfMIilNQc3mqJU3Ty6M9Tse
iwMT3feGF0QNl6gM+4aVahDjDcUxlX76p0Ajh3xdTnW5BRll4GhzshUF/GhGyQ0ARjfCDBYsJrTv
sTZwkOAWDgS4GfbcfnHkCvH6aUcBiQMDB0EPdKzNmr4reMk63pcK5i0kKiSIGzJ2MYZwrNI5turw
MBCUKLGCUyL3es7ZdmWy/C87RRQ5ik2mJPuYc9T0RJtUYtZCo7OAjE8HBrYitXLvFFZNqutK+K+J
4IogEBSyi81nertgh6W5Oa9IhF91G/KjGjMShk7UgBY2gtUyNJQenEhoWSycQfd9kjuRwlWwQAXJ
bgNsgPYVMwHLkuKcYJW8GrFGs//xsTRl/7CmH23t5/txttpSFI/iHvvCMbxGiNUgZLx/PjBPC4+1
DFCOY6i24FKfbPfKwg9isAkvlu26fl/tozrdnX+DesNf1XReoW6Lo2N8k0upxGLZnMXpl71mQxUh
SoTazIHkbD2mTEoWmSwtmZQaNJkG3O+3jEMwzdYPtdYQ7NrfjK507bmeRUkSfkoYt1qPvfLIByTt
K96YLcCcwc59IjUz0BrjSQL3RIwynox8h1tUWpADiEq4eeRWZGpfHfACYAmlVu0JdtoxIyFI2u5s
1E9s3Npizczl31sMgFrRdTtuddpJVHJcreluf0I6P/lMAB03Aj4+UmWn521Oqu/KGYsF7INdGGNt
H0Ge9OuU/VwsEZJ9D0EYnmsjyVFhlCrgiinIbYXMNhxhBcghRV5r4/oYaroPz7AEL1Ms8F6zIOJq
hmA7z7jOOjFN2KMUEFbACcfTJjZk+41rp3xdCYAGIOdahRINtOh0EsSsDTl66Gv+M6Ofvmt9DTJX
Y5lTsakZ40QVcTxVVT8ZJE+y9DAInky1EC+6HHS1vaSwljVM7YMCHer/5nSlQ2e7OtbA1VIdSbwe
tGlPzdTpeesn+RJcAYnrWq9F4dwLdfAOY5V/dljutgtecW9wcd0A57hot+ZEuCBihxu+Lzb1EXGs
hVlxoYlgDQpuzzpuSGHxRjII6e+ELelDsg3SijjvPXpnORNZe7XqcDIfCJVYPBUILZi3wtzcRBD/
naqcU7QSJZhBcWp+bZUK4v4vg5NA5W4P5u+775bf3MbvU1HXBz8qgtecmLM8ARVRj7QIuDGBhyHA
btqI1AorCLdweCNmmzFCdOR1jaIXPKiLDo11rP48TA7J+Ap3tyNIKcldfExMqK5FEUzCNHoUZeZC
14pbP+tEbcQi5Mr4nSAQsaoUSL/SMtBtwPDuJrTAh8rUBX80QG9c83KqaLKqqY8XBIKIaCieHxU5
eJEDeRqqn7FvPM5PvjB5tYt5zEUB855aLYvVsEW8ovmpcFDUixSYoGkNEvmRTAgr7pcozYxsHK4s
yE7gx0QME5x3iS94rNEflNVF1G8TXIQrQtJatBGJEFe2/XV+Z8zQnrztnHf386yRYEohL4P89S/e
CAtjtP2IfXdOxqJ6rfIMl/GMwhrHpsMbR6+oU77UEP+UOP2kM3SpVC85MhnbI4eSWP5A5RryKQxd
AlVECgyoDowCRZR/b3JZZbvKJ7mlGaXSfT/O1d+Wll61SWfMU5eCwf7K9P8jxbDxLlqAqbHO7trc
5g0+algjpdlkSxJUq80IfmCC2OCchghFqFkG75T1y6A2GqheE0mawJ8CgbQhwwvFtiC56yeaPc6K
hIVClPoMH5Ju8390mRJ/rm23RgD44Ke00DACJxyLiwjSKFd62O3n28Aki45RyJq6lemWMJszF9SU
fHbPeHfgCPVzL1Yf/SqmHSbS6GmpRP0f2+BLDwwBA/L3y4RwkLd16pdD9OKgvQu/4GYxVVU6Mh+7
vq8tE2amj/z1SvgWEaqtFD78EyKGQNSaEFqgLEitwj+s2EuPEL6aNbc1TarS62cSaD8lxrQi9ehZ
tc1hLkCD5v71R8m/hw3jc8CSNtyisgXMo3Ti9HdKU8c65O9h/WBd2ZsJWVfzbMl9chiydQcJKZ/D
TegSY3476pqMILq2J11dWPvdeR8IXaqtHuRVOq1WjQrUZHP+82Pq7pV80UJfZ46HzRyHbhlk6Or3
QPlIqZmjnCwKpJTT9rFQE8DhCeBz60jFSSnBAsNLjiTDZ+gQBeIbMIZ1lA6iHslxAfQbhhcQDxKt
24vxL5vJnjh2Wr4T2veTQaRRr+xAsB1VZX1UEfD7kXtzPlJD05dn0zCFoswu/jVlA7fOmc/vrUJn
xarja4rioAKl5w3av2SgAM61IBZ+uPAX5RXyayL7Zo1kYarIW/Ff3YWFf3a+hahWioz+Or7DlVgU
nerZJggNO3N8BgaRj63mBAiYBgR+evtyG4nv1V9Jrt4Xas0TlAjMl9KcPkuMU6Zn+gJ+9bIHsc51
6qcua4TF2Guhd1HmDreQuwAe7rMZx5WFXSM64d7FzSCXEAQyn5QiEngLTPvB64kXobeP3s+P2UO8
JEMWt9vJL8RZyO1c1T3N5Co3wSsDq31msPmV4BFXgFV0/TDPN0EBExd4OUj81VizhMeS6iauklYv
h51lH75l6BG9rASedgWTSF3xvKwdXHji3T7eabifViAp7aryK03+5S/vl6iavXGZQRV9S1lav5YM
6H/pQ7NALuIuTRNKtB21w7JZKXXtmTdnsobQGj61RSHfmkzpBXrCz6B2AaJ0VfQMOIn4ZwtsSUUF
Ds1lmuVJqJVQAoXBB3YNxe9r7WTme0547JO6egbhuN6N/wPvXDgVBWcnkhsROlv+R4T1JN2IVTQv
Nwjv5qqkfUPRVenFYbal4vgy8PDwna8XGZrDY6jPAWuKxI0zHzgtzJiq/K0N4aPtc+dSihNeLDtp
fCYT/k7kaMJPSZPvIuqtPrXH1duf0Fo9wTfRqV3VW3+/4V5pZ5T65y6drcodhvk8+GigXqkCP3u2
qG5V6QIAkQ5Lx0v/KDFjqbAX0DWAv2JDlC1N9CNeNJI9iJnCzi5hQt6ttlEnwLjhMYIefk5dMErm
+1jFXOHrOcMDbCgwj/yFhPw226Hr6pf3NSZ/z5GB//ILCmjEdvs+9ATxQR3cJYRbkbZ2/DV+Tbq1
hvU/LhAF3zQacyqeDnbyAO4NLcQcIOApYMc1EM0o5RDGkXSN8bHOv5EqJZfMCOoJdIT8ipTbR+mk
vyL3OvBqfvWxi/wJ7jFRfWync+3V1bsWkcBWG3fNdSUnAtVNuQF1TN7ZOwJQr0XqgygFpdiKJuhI
GnvOrpThpn5wH+CFz0MqRYBhfwJuIsjxDECVYEyDQE26tFbs+RNU5tj7YoRUU0PkDExDmLbQj9NU
KgyxXYyoDrcVOtcwjIkRU88xGVmRO7L21HjpYF+p4fcMRUIU0uy48mw3SQHy+dtNvPo6zz5Z54et
rUvTDokQX6hMhZjP3fkSJkuU7jWCwaT1Jg8hV/SCq2w+T8pmfz4/mSEapFpYI4BGEpEkUhS1o3bP
Fu694SA0EORGRvmkmMHfdEjFyXPVBkBGK/Uy2FoHiS8bPQZP/H5vHGZ7hNRC6LFj0g6hdsnynIdj
OSnOEGXYbRcTF7cSDWWHADWpQApzngwIr2Mv3IA2qntrIODTKGG7HlJsWkXi/Uzz5yi7s8HDrD1U
rRB4AU9lh+mmwNQsr+7U7+bzT1ZLi/UycCheLBxIw3xtkNikZ8P07UyANu6msqT9H8sKheIwRalK
HAIsXkJZQTYsMsyQgX9rhtn0gVkC/ifsa1qEOn7xQbG8RYnuXX14g0lU+//uLYugQc43cZDy2LaP
pKf8i5z8U6qn+KvX29tiSazUWrEjVaGIpWW76Qu4Wl799Qd0y/o1J3F2hrF4W6nUqcO09H9DYW6n
0HRUAWs3nrXw6r+U984WYx1rVtQ/CH6WiBkvMATK19TzTmwV6DRCPlhcuDj75gKMKmP+0r/bHtcp
HQzomTZbYsCpcxaYCzSO/fIYzst7Vpw1t8kE4NhMRLcI4+pov+WdH3ZeAsi0fYFgG+o+elTOHhHP
j0qRZ2crX+PJxDI+V9VMjdK+ajw6xYjU07fFlnRHdlnvi/P85WVQXNOMSnUbe/04C8A4zj6tN0qf
uVYJGydL3479ddMuH9R1rh91PORrw8SetdYVwwUaooxx8wPs10QtGjnNT5J5JYq6PpiWwuudnTK9
u7fjjL5/yDvwNfPP++HrIqlUsextLQ+PTurg1hocOj8QhoD+dt++cXJaL5Ku5y43CzBv2Z087RnJ
ZA4Z1A4aBAZsi9AEGOLQ146gnJ3tGIYe4lBEL3tjS95156ySFFXOu0HOR29P1sPvxEMdkvV8tcwi
z02y2o5c0WPgAj8G2K3vwj6x4+X56Ay4mJnved+5JXm9ZvAHQIEbuBWwT49YUw9Lbb78H+jWTY9h
l9yPmCFcwbYDosakTFwUsIPzwhc571ntRxWj8fnT1vcO1qxf6F7t2C2KQvq4mSclFMI+5Msmkl6c
WywhTkfUPflukK56ZN5xq4uMQo28e2UFpYzWcMK0rDeCDXaXLXr1lsPef9iQYvX3V8rX7sQe5RId
TUzmPGfoVkvyMyKmO8K8QffkNbOznypFZIB+acHJZTgw0SyonJrOWqaDBLHC2NNa11dBVXv4B3b4
KYYhVja7wzOpEZvdyG8X4FUXS+AcmxayLweseVxHy3mqn0t94bNPPDk6eIQzosnNdOIUxoLa/5tU
o2GhSV8Qcrvi5/hSKjzAc4pplkEjkpivXGTpyoF0kkL8VD8TPqlUkRNIQh+bU7DQ3fpDmq6ah/Ui
YEdj7A/E2sbOpooEpA/JuYv7aTBYKFoMY4Tm2SNckbs/jcejjAwtRtF9zdSck1uhHbts4jpQeoj1
LgX6AcK/IM42E9YjUPsnkDEAj3rdQe/NiEt24a4+maube03WVEYpqbrLnE/fgBITGj9tWu7yqV6s
zjAIbs8aqCGdMNnZSKInluJ3IkOS0CmMDjXplitE47G5wfbr7VgX5wjQNm1uvnNsT+e1/RtoQGFb
WczkcQlivwu03FOjMnQQUhLuJnEFBya6nfmOkueHp57+9dSqbtnhZmqEPZVOweX7UAxpd+zk98ds
o3UIsaxJe+s8JXLYiePU0GAhOen0e6SOMbCIpo0bYXMtfY4cUnYMA7RcQL5VZhdTL27DnhcYcyJ1
f/yOmQN4JzY4l3TgMxohF7hoQ8BylQc8Vjwu1t5cctzz0+XFXD+HpcRY80lOzKM6wPlL5RoZrAP/
aaH+nSBpFnZ+LdawFdms4tfsGMqE3oxmHvdC8ZVslyDMX6wxIpWrPWq1VouJSQ5YKi7VMj3rPz4h
4JjkWWHCc6eR5S/4gMLTfSprNmnCJ8OJqRXTwDRdQ/vcRy1YDqHrPfhKSv1lJAo9agQI2a5g+9em
sH2rW3NmKsroK1dNa/N9cB7+kSrDNKen4ZqWVDmzUFwBsRbBaRGQRDzbqUIgHOfcEB9xUSivPU0j
r2hdpmCEGqREEXTKY5KozgfnCPx0sL+nitIKWuZNpr4PX1fmHFE/O/dU6BMlUsXvt47ozoQ2wBWC
BgEq5LAFj7ZRDN8UH/qo3tsyGcEhD7N9960B+6vmYl9fKY92PjS+Q7BKaGCh2JAjDcnIEkb/CREl
QHPhuUd7aZwC6hN5ow+gkbnJf1MojQvC972MrNU0DdBlYu4GRGxJmD8344UjUBv2McS8xsBYLhBf
BtHxt+rx9a6izy1J8KW9zyxXIW5sl6zaXIq6Yf6/OpssdaaOvOFtVzEnWF1WmKJlQNs9r4a870q3
WslzbZGL+l+w1eUQ8AlbBJ4dJiy6Z0kuUHxrbk/uXpMhUMNOqebUE2+eE3dGGjyo9BqWLWt4p02t
ImeOwKD9OAib0ZHZEzwV7h5MVA1auMVHpHhO0QiT1okaKOCRNkOy+wLjysIt6bE/3WYoIkQHhVKc
wczXV2z2+GneOu1oZyXEQpyoS4KvdkZrNYI0hGP7hsgZjUSytN1/fAO6gIc9cIjRJ/Q2iTUwxfrm
dvsc2z8+cQve/JMNxMHlBly83ueLVWx4wqLQQoc7xVeKtWjZY0fwzDCqsaF5bT5V1N58waYnEKvH
ORM8Gl2cdTSuflztTFu7W32sMN/sI4JEgx7prfumBdapcB0MMu5L+XIPvnU9Wz3bLxtulaPR8nsf
D0cXcVqDcEZSLFRtmKy0es+552lGLA6t4txMljVdylRXwc4uBDXTvfVvTyhCYfu7UGofAcLkND9f
ukfUGb2jBp85hllXYmqIeXGI1Jp7ErYzjvQVOsfjmjPnIN5IVsr7YdZAMaXvvyOf61VHL98alMPn
s1d57wgROqqPwVPTlWGHuWCwMy/YDnMTSFoJTFdHWF6Me/IjcVwSu6OOGUfw/ji3Ha2nEJSoPb9z
+8zUITkINMrtEPklzIx4OTBms2K0co3S5wc0IQplEkMZ+XKsKROTF0k+aBukNEpfRK0CWg49b3MD
lsqZnDs7M9d+YRb8gj0M6/WmuQIBJzxgmrc8pa+38kDWSyhS4LvhSWAX/gZINJvu626vZk9sNRbX
eqZOVMUV1u54bnfzIoKBKqETAsQ2KXqbGEM4TiCdplbhutDaN8jrPhQ3XI06HKotX9aHj0qBlHGw
9Dx+Z1aieryebx+cg+nzusSYdbJ7eKP0uy7Oc7cdpNeI1Z+Y4IoXyMWIA+5+WJmS1Kp5bC0RfR26
iuN4bhykTS6L9gvi/8r7mU8CLZJ/upTZxuJL7vQruNUc2ZaZcZzW3pNax+EC6motjyh4a7kOj5qg
cStPi7EMbyd53EhGyJz/fd1+L8wCYiSzCGVcD3NCICpkKfgKfnsFEINEaTiICPB0jdKRfO1pEMuV
mj1L8AxxjmOep1Xg0ht4mgZuFQkHIdAfcNihPBs58LdRd5VaMqPKSv8dzRZNP+HxxonMf0+lJGnO
RwpHwdfzFLmbawkv/SoX8P4rG2LqhpGRZz5wPv2N6M9Hx4A2PQ3eBITq+g2KjxEaqNOG0ZYRCkPB
3kf3bMUGOFIvocm9zE6ABL5DMRuCIBAlkdS9xXX6uNOqmST86bimpXCEweSLOB9Rny38zzr2ArIy
MmNUj6tPQeSIokAt7heUovdRQFK6LNl3ObpSBlKKHIBktaRMF47q6SfwDWisqVPt5evX/fHQ721z
wrWtAMQ0NW+UV6ETBO0xw+J06SOzW6IaPCE6/ETW+84mT+qX56Tyu9mCE6zGbj9rkN/7duocENdQ
DzDn488+d9mY4KfPEU8gi/u+SyaiK8lKUQeXLr3wd3wHJVaZNWrAO2dc3V3Kaspveheodn4XoVO8
a1UO69dKx2irLsjxNR6DrmJJozi6KEJgnWh/L4TvxkpfjQ0VfUaAYM4OzLsvht6XFf0xjiP13hEt
UjdhQJMZahBovookYSHtQYXwaCvRW1n8eLndrh3SuPHfUuCXtAITicKSQE+BfLgUgsNIk+iecJrz
/lAVkrrMo00h7xR8WxAaWQM5r+GjaLgEt239R0NfJuAal9BI/Ld2gKm488YzGRIBE4afWg4Z7CKs
mz8asbIPESu6NPoo9aoQJFGrKjNOxutN3yDlnpBzGj/KYj/SijlVrLTwrhv6wSOGhzx1Riyy9XBB
mDWsN5b+hquGI4/smPwMCQqgOIpBN9RdCVhDfiFpQnO+VLgoFeW/iGxlyggJIfBkswEnx09pRVe5
x3B9Csf5UaysIgvvEZXEWV3GjeT460YYcJtzLbw5sgLk/EFFqiVOP3mZs/0yn7jX2Nkq/q4//KGi
WDqr/F2+Oa056uAMHV1QZOkeLZDQwwA4+VYSiBhTaokBaQGAr+itaWBQY3jwwQAf+tmWimQeImn0
sV0ntkYA+DvpU0sw78istr4IP1f0eNYubmVTE/LvTlTWqTlf4+oFmo1MPEg6W4r1Uda5vl4X29jY
KHFr/+nOOnDXyvnWdoTLnB+oF+0eHvGXGZJM2vqSr0ARHX0fSLV8uY/Q/6Q5cD1VZd60RAzX2+8s
H26eMP5Fp5fmCfP2V9QnINas0cpjh7x+RRvIuqd0MPCot+EHGobxQuST5KesOu43cM8oagRj2GcH
Ui84rbUY4sKIAUN4BCuzsc14P2XEKS0tT8gA08fvf/baDdrLGl7uzlreBbVVDnvpSqXXpP8Obq/3
aLblmOrtnE48PyAZ5ndGcpymEb8x+MMlJOT3s/+XvBNKDiysK+E8fi7fQKl8/0iiIaF4XikMMHTF
3kSDABFip/9nk60/dOPA++r3hNNktP16h/F98pqu0j/ZY6rbAfMFpyYvV1yZoA6bG+xYBujN3gq2
QBbbnQWN4dEp+rouIKZRQqSMyGLkHB9VaZ+1FZgKDcfkUqft3SU9vde7Sw/lueWe89mlQcG3H0x4
DtPVJJ3AkyNF7IVBtpEUYYBTfye+km1zdAaiMpLQa1C2qQRI+mqgwcypcTjTQTMtJI2F0WlVPqX0
qm3xL9YTCgLQIvKVgl76vY81noktZmzmqe/rnJ+y+9f2SktsrJ7n/PBr+6rUDb71UX23LgH3/Uef
fuWBa6uQTB8EYTQ2AJkgdVbiG5yLks7Od2CbKNqN4PywkIxCkBSPROyl+xhmE5m9S60R+ASzJz78
9skYavtRRgZZMpKGxhR6aaXKuF9VxtzEY1FW7MOGslf5vgOu/CydJSZgZCYzHvH/IhAhrE5VyLdo
8gT5srbq8YbKKOVGKjJYqUH+1+KmchsALSTzZV5XgipJg6PDWrPCjtfmiofbVtn09qRtVlUYBTRX
TbhJB4FdcAQK4dC9oe4m6T7FMsald+nrNYtkiY0S5w0dWxheHj/BTEsIr654mkw/VxmukN91Akc6
2hL0xrho7Ah2w4c914k/1IFSh0cXQhXoDbByIVjmGkxg7Z8EpUQLBP5xJQ7GDYk4o964mkAFnBSm
HJWsVk7SCp2fHmji6Gr5kg59y1yfq4r4Gc/wvPRLuPDe78i1K3yQnRIYM4VSuY0bx4NRanzGyUOn
dzigwHE6J70HZeUcs5XlQFh7TBYQBaOknCKiOFYg6cxC5hYm5y91P8gjbOJihnnz74jECAMKIpDF
lyjZF9LEopLxrK1kPduFSjqbX3Y6pFsBype/nNC3IyPbwmF8Y7bZfYgS9S9QdwPzCFdPZcTh/h5a
i9kAUiI8FeDWhhXzvQik0IYIcZQUVMDZbqpZj36EfTknU0s9ll+jn0qOJS2v52C951uGIgyjlkQR
NpMOpve60NrOOcLmhMdneoEm150hs1iBtraaUMzVqK82URgYRsaSMQh5paXV3L/74PFS3GAjucxt
5HBq/pm6eLxR4cWQb0Ctw9HDKnPGdjuTbxfVRl5O3KJGjCqcx7xXyBYjjPGEt98KM+NR9Hx83ytc
Qy384LNRbv4G3ckEZlhHAiI3yPI5J7mPTn4YR5uyC9ibepYD5rtDo9cJexDS0UQw/5GUVKEcohtC
Xo3KTUKfyn5xDraOQ8ytuoS9a1dqOTlGjtJ9P1kPx4q/5kU4j9rs9rMnUJ/FlaZE7WgJXGJ9CoDn
xxqoPilMTKH3Y6vthG8P2+7kUq0CcNYM9NHf+LkPGzodCE5/2Smb+SCUDfwuPJf0vap6nRI8zy8z
qy/EEh999iGNaqT9RBbN7m3YzfzBMNhMDEd8On5unexUWbTpliYZzE7jvRMHGHpJMLibXYJ50PvF
PyE1/TeaZIxCsh7hkV585KDdjL1WO8TQ/NDX3qHkoBzU+N3Zo5zOgq9qPlrUONFqdVB1Ak+p3kNG
3/l2V3EHtnR9wjGll3FeuXt1ExdkTOcTCdtTotduFt4edm4ZrwvatyIT91dPWQ4bmokXnGF16xdi
stAK5A6vXZUmNdC4q0JM/qra6KkG7QuvHwNbljoXtyvDheMBck4lFcrAbW9cjjslNHJ/MUvUTvwd
tZZjPLNsN+2dDqSN9Y6/aUGMypWPR0Xrfa99atYeWnmSysaARwJHHDLHIdxDCJS4pdx2B/ShWVfq
hjyo0nPCTOL57KYwuoz4aNdYusVTD926n2WtIvNOqkDjUvSw9FI+PB25yo3Dq8Xlm0XSc0pYaCId
E+OTTSYulbAOsncJ0H03AnfRC4tmCy0V7sCMv6E0R1ZIQDLQQlufHncHaNzwuesEA1tbdUWOFOch
KMlPl7i57siDf3pm2c4A4IsCdITBrZm3sMSlo/PUh8TARoS2dSr7wC0hh65MyYBmtl8SFoqTCgUN
OQoy3ycoX/vmJsGHrMlNGbnqc2hJ6cwRgayaoM89G0yIYIflk3BiwFZu/qSrToKRtBCZYaytdHgZ
o8yaZzphmOYLT1FfcgnLOOAyFVsQW8L+uFIBOz8XwXcdRT5DHyN3cXetN3CmPtPL9JDAgLzbnSN2
QgF5OG2JmCiC0G5tEY3pGTId5iQBoTlCngfX5gMA+kyxhkjZ/Ya3D7ec8Xfg66ghbRzbaZNQlSaC
g9s/9NzU5wxr9hltpywP0IqLFjNN5slq86HQzezuQHJH7jDgcKTApW4CVIqc3KCJdFosmdVWiBeS
Smn/KEYltUJcLs3tlaXEgOOuQ2DrhYRRSPxSFeWwi6qPri87f53bw8jkc0mrdr6rEu/fg8ERwPNc
mmFfZcfeiYSR9V/uRudA0yHXxXAj689o2CzxrKu/RA+Anx9BYug2oDc+FoXdFHTQ9EBvQ/T/HzdL
iWYaakhnzFW/LXrqg10Hp5WSptLO1WdkEGLLfAV4Thn84rs/S9ix+9FY0RkJ7kEQJPFj0EE1NKTk
7Fzcpwk++al0tPdI9Y4pNdG/E6wiYIVrQ9/Wp5u638dpHbWs01sW57RmAGpOmsQlH/SiF58ryyOr
pUI8XIIz6OmvFI6Zb5leyGs2DYwd1fBwMXzJwI66ApG+f1rkpChnA2FQjKrv0hL5JhNMzaAl6Cp3
NL2Izfxpa8ItD4CG8tmKaOBhYk90lG/LIJWhlQxdxYE696PljXWkaZ/d5FbqJeBsdLx4kjt3ciKh
5in0iTYrZAsJ22zPugEYUMtHzfXa2dGV/MHTEMxRAlFx4EFgkYkUlDZxQQZ45JY8L+h5RIdYdY1q
UmFrSDKlXfHjZmUUnePdJkOAtEK/hPg1QFZA0MQ4De/J/C6/a9SL6ckJp/ZVtfzZ3HZT4Ye1rAri
Bq5MOsjbrJsawzZRXSKwmnvSc7HOMZL5zCDEvWXnWB9XCShpXrC289XzATYZIatA355Mv1/RMmtM
4XzfeP3e+/MRMhkpy5Hc9211EtvWVSJIx9pDkh6Xop1wZW9q29tu4ug77vdL7iFQ5lHQNQPmSm/b
inVdb1NRmXcGkDRS2wpMlRF72QHz5FdyFWlmwihnxBJOf58Y5/iUuQPeg0jOyeVib9jH+yiNj7i+
27jGEGWJPiokZstJMK1TfLedktEvpuMT9qzT33zPPKx2j2I29jNEfsSUZ+PHciBimaiRF8Wxfu+a
mnTRqEhLKD1CcJ64dYuM5j/wmt0DwVQcx+/3BLBGarcLukOtJCJ3rS1HeorFtdXhVzKjwMClt9IB
mmXVsFl4CQzCXi0kEsOSr5hY1OI3Zaidb6th0P+a+/KMjAYtx7QEmxwDIrH9HyjdlSXwgtC0YyqZ
5LVFJL+l+WVewhMEAf1VXi/+bOAheODxz9cL0rEOSPlFRDsiPz0i43TPxCh8V9UxNUTgYqoFB4lR
hW+CSW8MaXNKQ9Q/ReaIHzc9UhIdGEHGElbBxLughTo8pfNpSdnfgI5KU4i/yt1CPHyOKsUZi80C
VOYrQTCy8+iG176xHf+ykgi2XFKfx4SEtb1wcgU8FDt1lyDtf/9hFXTBZOU9BZF4htZo+FBA4Dbc
26lKWZ4iI7bMCfJwc6VSQWcmZvctqdUU9t19HSruHdMzmErPVvn7EtY/d1CYLTJN2VYE+8Xo4Tgj
mQ2tQuvrjtL5oSU924K0+qVbzD+dxTGidrraEQB5JsWJaq4eCV2g5kQyh16xk8ybdLn6GwM86AW7
yI6MMijEAIR8V1TEalQ2TtA07U2sJoyl2Uvaie4Ljm4uOUDb0CCpZ+9BFWrNKusvynIL1GMnNaDk
5O0jLCcR/TNN4u+HU/+6C/E5HOmqG+KTwr06vtjATxPVLsTCuYXXvzWe8frGiDXtT6ExJmDfesHN
CwQ7GlsEGDa+pKS2NExEhIducA9tGy653CAk2tWZov1iXWBSILiZupwqU02U4OUTxKT0sxIqVcdX
2EsmCt3paudGLTDAq8R8La/Ia6YFze/1OykpWoBga2fsGnuGMUKwTFh2eBk3K9owEUIBHH8EFlAX
N8zDYa8BZYV0+bVUdDJ4/IIulCxfenvuA7JzUx/WDjU8n/m1pPAqaC8zuAjdR1aPfaaU1YAiSfL6
hi7GKoUbgQfjek0rkVaPQ3aD1RiEcijZ9sIFmySe9XxycW1yDEPyOEe11wkCmdBttXc4FuwBjD5A
p3NRJZXR9mdyBw3+rRw9Jb5xHlOE1nSUXnRxRfASpb8X1AwBBCvMGs6ZKpv5lCgPEIvgjBfy9CkC
mhm/3i7i7deJGRNSfZu97IjpCfqzWdCCoL/0Fa5qhI5OxHrEENNWQI3/MAJG3vBFpWSeEHaYVjZU
xQDUdOBgEzPqsjbLU7SM00jKquw8sPmXX/W9vaSTvfWrTxHvmyrH72G1XXP9+yhKL53dF8tRtRf3
gA38dfJFADJwN8UtwW2zr0NeSC9WeR5oSEQRNGJLUYYIQpDE3M2dTc4ykTjuFr2AeJ/6P61GCCie
VEdsSDOAgd3i6HLNwBgtIAF+TjAE1hrgMUBvw8Ueh/iFlOp0hRx0Lh7nDBUlfcMT1dD4kj5hhXrY
d6ax7VQKqYRm836TEXNqdKtUpYhFXrQ/SIb4EXxU+oddgo/T8+iegMto9o0B6U1E8M1p8qVCqLIk
CKXugrIwjtBAPN1vcCUePmZmcG42qPUgBoFo0NFcJAwK6Kmfr83UnGCpBPIKrJs69C+KIJhlM+OD
lqlar3FWfm4mDt2/NXjAN5IQzV74uoiajLdRLly62F5L7mJjTvIB9XKUAugNzSZTMQ5J0GSgJNBp
iq9dYE27VlDTG/KKeOw+Zk30Nt/7GX8MpMNYERjGWBC7ksuKVYbaw4V1RFJStse1xuvvvSJcABio
BQm5Qle/TX9LyS8snvFOMne2zNO0ezYVLAb0t4kVFctesmT3KvOgdyS7Ivpw1Vu0Z/u5p5AY6hjq
XmYDjm5p/v+BQPYf59WfgdLRfDC4yknLlcLL/VpSgTJuRuWt2yTMFjcwEPN+HMhrYhLZG9yNKVT8
kQ+goOvvL7vemGLsL+4XQ/FYG4OhWvkplHAV0h+n7R6HY4+1L87gEw2jtryiTrr01O8irtQD2OAa
FJe9AT91F30yepUFv9VzT5goOyUnWQ1E53X2EVuZH+aODuAlKfUUAP1eGSlSDa2hssDpVJpQDdgA
idb0VItWrB7ueFugxUoPoeihucSeDyPCoyFZN3T2rLeB3LZiEC+vpM3v1b4SXecCZM16S70XSJkt
ZQlBFT9dwpr+9LmjJv1KU9fwjB5Kg+t/HjNR0Zy8jybewRa8TzDUIBkydQCM+g1m8v73svZFpKnY
Q5vlfsE4Cxefvqga7BCplQ71DY6nh3YVMxPnQZifkwi+ghbShpVY61AuH/jFrFMfaOgudH6D23B2
MignnEQqBZWtj7YDSBhuzGL6JVMww302LZirpojwgS0WTDBwi4fCCufy5V3pMwFSZPX4SCttjPSZ
M35BjSOWDRbIxRITf5PDVDYXephtukasXAeva5E4UGUg05boAsE/tZMXpFjD9IL2XtIejT0yfLeC
sfck58L81eirEkI4KQwdSvR3yFTTaIw3rKbFCPE6JnhURLQCSUUBar//ZQ4EcuBmeAiKB4smsebR
jTbTA6aG4ZyF6Tyy6dzsD/sbUenoizzlWYNOEl8ShGpabxSGtZ07HZp8asoxdZvuAYuv98QEbW8R
sbgxkOxoKTuqTi27hYYFq4NQH7MCAv31yGxtjD1/ghBLQUJcopHAjTuLXQUjvsrqpj30Lh9ktuOQ
kPEB5kTST2lK8adIpiAdJiO5oto5WaRuiji0jPSRO+87XqJ6dtx0Ma+tbSXEJue2lZMtKHHHR1wF
ZpYN8OsCRA6mcvnIiDIysPhCuvOTTQwEBSr7GxJsRItXiraVOSmO96OGxIxqYyO+oeEHqLRvqaQV
cWRegs3HBygWl1ufqD+SmWhXJZD+C0kWh0paNt119Z8UdNwhCjyaTnk4QxnCwRkUmrbwbgg7E89y
pTLDB6joaM6YcMyBDKESK0eElIEb+sP/mG+w2acJ8HJxVAVknU0bqycG/fkaeSRx8OoQJ6egJ3DX
Vhm2uKd0NK/9MAytMgOKNVegAXSuNTVRY7iAhh02ZAP18bQCpi+Nt+Z6jqQNqjnjD+JkmFn6wtbR
f5h9zEfZ4J9pxcS0LDQHwfXpx+Hm90bzoi/NdLy/S8WAFhbgo+FUsIVwa9pE0UvnPqvoarOM1Zg/
BU85NeGT6vCDmH1l1XaP1RlBVRVtUUIbl9VReUqXf0Q3BWSQrJ5zFVfhdEnAAnb0+esCSOp7tbqZ
DIDmteHh89pR4PHyhFS/3iJONqm2NAZ7oYyMZvfghUlcYQ3Bye64ItDZ8P/RTBqJxKZvrB3A2dIr
gHVoGSzFVg1oUoaE6hQDgOPoqVIKPK+5Jj0FlezFaUOfVZeARxba6rDoapvo3bihRKv2UHllA82f
O6MlqsyfpGXgr6FSUUisG0jQ6QOcvAAWv9b4TT+SaO3wwLYnxOuRpez1uTw06gD6cNzQCP90t/jc
ydPIK4UVLhQx0kXVhJKr0tVXu4Te2yHUxghUWL51t1UOyAlwD/oCBPyzq+KNpYBsgh3a/dS3YO9f
3HvB+0PnwFQHmaVUzX5MRqcIJCnhVuWHf1ExV28tP1iUrDvqrNf2Z6SmdkoqssXok8LFz6FoLEdV
SKTn3y/ty2oBpkZyhCTvO+4fsFtWtqMtYoNQ5FT/kFmFDgliWvkvkjz6L813caut7vQ5Tb8Vy1iA
0hJ7AOX/y1l3Ts4II2bTNJG81VyIE6vNzYCibwRbyWGXkwrZ15XavFAdh6bs5znrD2cBqFyeGV9Y
uATIQKBsO0Dygmn1JgRrcsbXS+w6xgrpavaZZZRdeTPz3rukFEsZIq7XWBKEw20c5dOj3hQlCo0A
FQcibeQZf/TuCStJHaKQhrOBVzuzHRIba7QM7q528TTJ/TisK5z4NFEiWylsJDJcTG2q379WBtuL
tU9BpAFVllLj5GFpa3pR9LaM4eevJzXfWrfDkLRx2GVcP+XCatELrxFLEBHhLxEsn+2McVZy1KTh
FdfAjHzVkda45XSczoYMzo6n9NsTXUDPiW3O/ymb6Z9HjeU6rUvsP8rTzSnRct1dY8wQvB+U2QH6
B5JcknEdB21v8TKvscTgip4TUhaBPeGTHpWBMQkFVznph6uE+qcZ75PmLbzyaSmsmztQ6oR4q4AZ
ui+fPvU3jMKtRXZltwuCNVAi4DXWT6RQsMaZmYP0pez+ZSMWTFPFKgcU9VhkFXEH7KrPKQdsSupf
4fCidS6lMVsg/LsQjSfTUnGlAyblUAtUO6cLWlGpL7VNvkpfMk4H4IyRKHEjrBjopgq5Vj56iDnx
abk/NJK96vuyAh1A5NygdQvm1R5ZOsJ8/FgFaw5a+L86yb3vcv1DmUDUjB6tEhzc9nEQOfdGSPbK
SjNcmGjCzld+BTsgCGBu7ZYqMkr3wQHuP/eQ7oF42iMkTX0SL/Qgu0tGf9RS9APRw5mqP2XTpTk0
M2RvUfakZs+S94lt905Pl9ySsK8ghYKSNHQrqkpv5Ut12n3zrQK0g1hSIwsSrTJxaWMcPQkRfEBd
ITrBInBFvM38dddrutMXmKdRlKQJMRbyT3tLUbZVwCIeLbLZPxlFDQHhZ6c2fjbzuOCPwESLphkf
xeCnQierDSDpRAdUBB5RmvhWkuqee/ydk4TUrzNRx6O5pjats/Lkl2ANQoFSI3PabHUwAIJ3Ojk/
hjReIwnt/sHLoAnED9eQNVUwZox2KjZYfk2WSK6MxDvUOsWF7NWssLkSLHcM47tiW8cWRSd9XfTA
+k0e2bBVHkW9ldWFJYp+M4vcYMMvoaawliEMPBnpH2/uqZzZK1RCDl7IMRlrE/Z4cTeHCLzxIaE6
4Vn4GjLWq5/DaCCmowGvQfO+I3WcxfJY1acLrokNqsJd/VSZ5nySXAt5KGX2GJSc97IJEFABIfRb
mlWal+3vqxJwQD7J3xqnrxuSd0qHzWN05WfLlfSCT2hq+2jTmLIjVI/0GpISbF9jvoj9iWmxyMcI
JrLqWUGHezYViFsOA7qErm2wWN8tAephuPtPHq9h6+Y2pIZSFmgmfXvt3uAB3krefqcr/CmHuUXl
pfNdIxsi8xzkJPZR5KzCkTuTB80udT1QIT9qyD/xMYIOFAEyPEnfay96EmzXpIcMTpyYz5MG2Uu9
nx40MriKsN5Cb+u1uU6NH8VmAVRKyrw0IVVZLggFx+qoe84YjBoF35F2MA4tLRD5hzGiZmFrHOzJ
8buId5NWes7Zpe/3AQiAvtibE9PGGpkv0iMnJ/tvcoENxXmUEFmxrtM57fItvv/FHDTRLtw/ezoB
McJDwXzqpv++oXNBSdtaOOdJpU/MfHE4Seu+ypkitHr2Ked9Mx2U4l6JAKofGbbwOKFigcnhqolk
YMe0kjcc7u2qWn//TH1kdkH7TteYBEqabPgmzS20y9ycYWopcUKcAprAPz/sePZKtrFpKWM9Jc/0
VC40lkNaEyyb4eOBScsctIlbO3IxGRKE4S98xYNDdw7T3GMY6mC6Igh1f2p4Z9pp4maYvazDB5Lm
4cFKubG3zHycrXjl5su/Y/d5I9jeXkuEFEBLpZJsHvFUl8Lez73d379fTZbcKbYwLG0RqM4ik4hI
ISzUZqhcPrBL8zqLOvoMtLwdwkHluPO829XTWSWV7A+qv+MCUDZbToti6gtQJGUI80bomWGY/B5n
DWfnNka3tZNk/hHc+BNsDtfpDuVi8IIkfpQYZHcD4GO7H8ZVe7Q63c+vw/3DYiWc+51N/y0gMSIb
2mSUO4LUb3bWQTd9AsXLoyowcxRA+n8K86rQjG0llLkHVymQHpRcHY+M82Kf53Zwrn+1W+3I7RAQ
vrfk47S87s5cW8UMRzIJjjhX3h6GdL5SjVMr1MNrXcLAgatb8nvzIhtxo5KkZhNNvTFI+MUKOley
AD8sxWneEnaCnX5HnmCojJrJnF6zU1HUCFalpj8/Q4QDOsgx85ssK1SdLyOXq+MAsXZU6wZc/1ux
5tfR5t9wjnb0KpIE4/ODQQNQvwq3GeWxOvAmwcbKIbWj5EbVFj4QimbkUjk1wOKbWGWJFFFB7//a
f5ZwqYFummffS60YQZenwlqTE1Wrj9WsWekDqBw+RRBmf18vZolYDBT6kOIl13nutB8ornZCZ+8T
0DZ7nmabQ/seOGgaGEl88pmtcghr4LZzAyM86ObYtlJ8sXnPBVPSktlUVpHOcEuCup6ENclDSMkd
pLugJYkrkM2TRmx18+R0xhP0Z0sEmJo4WsVn1b+CgpPkDF3dho8u5tFDHeLo1d/aUp8niHctisdU
IXZHfGDgiJyY4P/rQjeFDm/L65TJFyKIWayDlhuXbenfHQVhzkQLCddHaT0L/HGH6gJVkYcnwjAl
2thWQ6kDWCCWmK8M44y7Ne2oVswFvzcYFpfnNKlzUf2vU+ZfsUMtOq6j1GleLUjZQKgZBO9Uxv+b
Frl7Vcdc6+SuUNAci3FAqXQdYcEeUsbdmS7fz9WxxrMk6SMaTpyp/xJQ8g6Ym971/UzrOWT/J9De
+l+KaEyFAMGKVhDMI5G8LjEelHl8W/LIB4CS8zImTdF91lDHhldqRPzqtkOiUuqKVvDLClNYP/US
inBh7zfxMixPmRpqKcqfIcCUrcG0YnvnAnVozGs+zNkn66wrO4azT1bE0xiooRBGq4AWg/eJ5yx0
JAXLRvcOZrBDVa5Hdq1OqJwBU4W+E8Pj7uBACDmCY+niCDEG684t1zpfgthU1zthu0fYnqUDn/cf
bpXiXTh3KehKoEHuHicQrwjuUpEookTyYkyyf8hRo7qup78Mj6Tkk4NCC6EVr2bxuCqE2ODveOpb
wiAmYpR+oWvrj2/bFfmRqSJIWfpBRLS4f2ca6HoCKX1LKEPLL92ql1+PQcGQjl+LKsBvCqfQ2Zin
LUT7TW0HECO4gS2Ey2dgsbQpLFDDQvd6v9PEhxdRH0oETiciMqTiAoWWU3D7FM4l5fPO2p2oEqd1
XzbAYrhcFEDdDO3LbogiqaGxgrMfaWt6/RKpX7/pVY09EMrlEWE83l6sc2ydYtm2d1wXup9q3CHj
5ixSkH3Mp1EPSHEhBRHnHoT7V905npq68fL1bd0Xv3jmVfeAKzSZwOHsPLb4mwAdt4rfPTIcNdAg
CDNnBj0Htrv4CwdJYY9F/AOHW6c2gAJt8WsZX9c81AklkrRJcNXiEzKQqwt3fmP7o4bTSKYSAi+r
dYN8/LXw6L50Qes/+Pis8KEVmSf6AKQ3PiDYh4DInkwbOlplJGzKCB9RhWkgRpGydliYwSwl6tS1
1+lM7hd8vcCZYg2QaeHfhSj4jmW2PVlQYqpMajsCByqD5vgMYHzPGX84I8fRO+mn2n4r7Htbb2Fw
b4Sbza74W1do2lSZ4DtKTb5F109oIEGytkbZNGr3vM3zYZjutv2Zrh2AeQMQ5Dv4NN2l0Get+Cej
ZzQ9WNvGOlz6L2a1RxFm8pztsjXSq+ZQcS+Tm6oRKqHdEsOBA+VCWaHoodPK30qGYqlT4PKm2mDJ
ZMwEVw0SBXNDveGgIGxQMKgIigIsWfmCqu4tz2ICa4FqhFbxFYlouFMeywdoHXLfiNOR6tmQzP/6
5Gqmn6J6d0AXq29pugHIj826TH68n9jgqbRjv8Gw0Y+MVtlvO0mxnywt0PygWyX1SxLQCtD1FdI2
CPWbAxR0jMAkkO0rE/NSjykKHR/4iqaj+Zo1aOMWo0bHPZuiTimHw4IeJjNbpCd7aHUv6Qe69Srs
vnCIo0hKWzsqMLfkkpe+Oo25Pq8abi3JMD2v66c2DvFC17cQTe48nHU+7FooMVC63PgFPtY+oSS0
RHo8fn6SuF1AGQS1MDPRLvqAHlWdiA4yJVJtCn5JKVmHt4zxZDBX8Bt0h7tHxM5Fkgyh0uzWlaAP
m4gmyTuV2EtiEir0Mm4JGdlzb+SNJuMY8cLZMSmS1mGs9WtT1isWJiFwzlEzdoqm2sIJTekhqWdV
iWgb+OwrRj2grahPzXyVWVn7A+5LOe1b89Qy0ONztdHlAx+Bpm4lYQXEHf0VF239UycT7NZzNUvv
moW3oGfWXZTPmBOHe21I0hw7KebKQA63rpVxHW/vZF8PXdUbozmq6YkjxJXhJMmeHMQG6uD17gjn
q9newdAOzYx2LAfcdlKL8LJk6bozgViGG1r19nedCqKiNgO7YCWXjI6qrDejdl44is8yujegQLpY
whKOJO3F+fC1zt2Na3PoGp4Xg4cwU9PxfVaDRE//jAWnqtaY0K5yI8DpitoC2eHmWgY37JtRqrZD
XDo/4UlZb0hR/hC26b9302aP/FmbrzxRMxrX1GrUNUGHOK8dG1kmDjvuIwHyd8X6XAcTYXHyAKEP
7MjTmvCWeUOl++si9wRKJAL1BufpomQZcAEmkZI2dWQdlTsBWLlZLB8PfXH6Hh6L2Ijl1IeBc9S6
/qaTkFUBAMSMgfqpn8VyWPCmYGczGlm5sv53YPeMah0vjIXPonHrAzH1hHe1z/l2BiVK5fuK0mNg
VBKn7SG+2Vg2P6wquDPe1gSUaGX1aR5vsZXjO1A29BqlSx2PaLCvmTY1387bsiXk4hJyX+ZJtGRQ
XABnBvOxT7d4aj2qvSJLK6rPPGLtmD4WdFKTjBP1ErIK8XeO89vgRNIENOgN4/ZWVlPVZMO6ajqW
j2Cr8V39VJHqROw9ytgtvcfc863+7m4nQLhpKt+/OHqy5yk+ynYMNVkwXgxLHlbvQX6IeHiCzfc+
5ci8WoOPfUgGVvqNhkDzz+CZNTJul+HrqMd/djFkyLRe6PlBZMgvgqlZTPb97JXJy1T836mCDy3d
+qD14LlgcjqjXzLXBHIlroVlvN9RNYA7l3DfVjcTpl8ZAtwuyUK9juFc9i1NS7ut2vv8ooL8Dbqc
BTbBvE67zzuPMFnhrPLx8uA1IfYJFSGV5DSkTkQyxQ0hSlClVftIpOEYd4UmfU28qT9W8vJ9416q
+t7byAvZTo9OwYd1BA6dd2vz4Zpkb9hbtA6NVY7h21trneJrq/hTM6VXb0tqc7Rx5Y/uAJM4zHCx
SlE5aCIJSb0dVR/u6VENkdsU2Lg2u8rd3LwZuDdh4Vwz8YVDFXXmaLtSTd0ZdYdz9fL3jjQwAiiB
hqYGgwBlq3p3wjv6dcIWMUM+4XObUmYOUrNkp7VOBb/s3VDW5vpzBjRFlRRfnsztGduZr3OZ8nbj
PiUcch4VkxbquPAuNA0gSiTluXidd5sWNlWBU+nqKtcZtma6/Iq9J3m+fmPWAbY/nYyhivOOR41t
FCVpzAICLjmXdkBIyr5UGxCxQaaX5R+T4JAgpkV+JX7VP1iB1iXeVbu0NSx2CA4bgThWhHSAKr2H
2ETvmbaU/19r0ucoc5apUc6w/H6Etg8J3pddxLWpaMpw9BcwuggCgIhBCVS6gvw0Pbhl7kwrN94P
bsXEbTOHQj3FUJpOYGVEtTiQ3ZGeRMUlIEy0RuHtuY2WU9hCY5vIfu8WKL+NXIWaDIaqVh98RTTP
dLI2XV5m2Lzqt9vKiLjvgonnWGpYs2hglnuQF6lLauJ4KHphaoZtpFwiZVxbWMeL66ytJw3xTkmN
mhxV77kbC4jpTB3M5jMqMf5tVreb6t9BSQ2gjQtogc7jnE2ZvnP9Bpe8ZqQ5Is6MeajfJX81I8i2
X3Z5VZZiujuzazE6O56fOfskrRmFdBUnoASjyyOiB2Bof3h9Wkpioy+pYMu7Aodrad/ovE0z5i6A
1NDodWcTfF8WKV+KUYmftD0eEY2qJNyLMgd6OiPGez3rA3kKmx9O/bf8Ouh1WCr8+9woIM/iuvTr
9aJOZuwR1z7k6trRooKnJ7x0S7a/jiCUJlN5Dq9l8H91AgFO4nHGVUCGhGK+PW/46Bhh7vif6a3W
XC/VFC7+eme9/3lhqyENQJfLiNMchfw7ix+h8tmX/GZyWxPWZY45yI4Gwqa3LNxs6NR7m8o5p90K
MmKievtfOaQ+oHXH2eOM89dwL9jvaxMH6FzuVc+6LlUshjD4KU92Cm+4Dr9mj8lBydDdoImsCbgQ
4BjOzhtJtsXrcoU9rsTadCqbYMKc13HPq43Z1Jw0O+/8lbbVwrRlv3uaY3ZfGH+VR8DBC/h7t82G
gaU4FnaGVPDrlt3mP1WPCzY1jEkCrU5yz8r+Wp2WSFNUJpUG+4otRcnapLCFsy+1cjEBAPKFZVXq
nn5+C7VUqukQSxGAc695HamVd+E44ugQ+nWC8gCOEU+0Cq1rVr/bt6Ask88OW6Ghg6B72EJJ7VBx
GPWOcbX3D33B8xhoPqJ0k3TdrOdHlQIsDXUEtYIiuWnBOzD3v8OxMb+2E76bK/vHE9laCJYtDr8Q
2/tgHkUrPATMACcCg4jt/kmYCOwa/qGWVuODQPQfpgTaodTN6ETmP1JQLMwnhzimR+r9EdJujSjj
72ztPAkXxvNLYbDkwe8bprqClMGOrlXtj0G1XMeRnNrFqHhf5s3IODilVZR/842yv+da9YWtn74Z
hK6l0yljNqLleyBF1z2Oa7RnhxNhpcxgog+4NOfDvB31Nfa7G0cSdaYCqx0ytOZW+W4s68Z9JMi6
UuBRJyhG0imOR5HIbvH15a2cb5/+yRvB9bNnQxHvees6so251GJqxN0rxwZmvrn0afkaOADEt6Ko
IoEm/IgtHNWpM0ksvoNBEpPDBKNjNPdmtTRZjWYtFWRuC2fJofYnv151uvvqt5OpCsVxRdhWGmvl
j4MyGrN8O94YYR4I5P/0z1D9mKFghmPiRrCoB2YhLyurEx+xij//xH4IfpWgCVrLA4gstvWPs3dS
uHe0R1e1HWS1IeUWWuHlPLDb+RdddK4BptS8/xHIkbPYsoA/3OuK2FVD4IlBMVik64kzHpk/iNRX
m0up8fJcC8OQYQIG+IfefBJrPrFB56mg66CKO6ES7zxS2LG0C9mGAE38qJ6da1yUkjNN/8xR2kZi
xQzLJUHPlsL25C8Am4qe9VMGV1I7WfARacVVb+hm2gxPZ0DVGdY9sJfB7Sg1oBek4M8jfknF+9UB
UZABZ6vZradTb3Ibv1Mxzd3mjgAAhSAEyAkc5w8KGyMxzGpqqOZzSDKvJW7P4uOZC6fjs94Zdvfk
98w9s3BrBbjEzzRgTTOKaGLOTBunAjRTmk3gvZ52t+puMNEKTL2FVglnCngQrLQZv1hzATejPxvH
xDvbwmuKgxZd1F1eSgeMcjwrDbTUhupL4Zn325RMbH8fL35Z9rUdAvmcuReuWAHEglJf3KP1IC6V
QrtkCaURKj9+k2J4EHLdhpEgiObAke/m3RXK5gfPbQe2EnniAB7QlN/8iQA5mjCu0nwYKE/AVJ73
dT+0h7dNvQKuLA1xj4XGep/bJZgfhDBkrGzcCp2SK+FvMi+w3FTm0163PoZmUGqZ3CMKTO+Mxzu8
ICxiRieX1SZ44RuJnvtptY7fyGVHF7R42ZW9+5o19HXRfuQ7W+/PNh357Yu2TY9tJZ1vRZESi9o7
ya4A9mHs/eE4HLLl/RYSEal889sLOSxNi0xRlyPJyVSl5aQscOsqPopvGQ3Orooi4GenHembHEhI
SgqvXBp6eppZXL9xc7kyTF2Rpv3KVrYoSpI935I/VpL/0Hc2FZ9DHYypmjfprkS+RZu9fOBtNYo4
2Nogwsx0+AwhNkgEbEOHkYFBUwgJf8PWF60i0T1crQJJgIRpPY4QaVLIY5ichzcu4Ufm5OKxvMZo
bCbTFFyg4UT+x/1OOityUIdaZLS4KkPT2BBJxH24s0j2/1gK40/cH7zbSNL1OHfZPS/CljVKCov4
V4/uajNw5GVIZBsSTKTmdHS+htvue9sm5291QYyGD17u8cK2EPe8BB+/lLKrMWKCEwQK8ZF8wlH0
b30tRsRvWRgucWEBkyTi4cj60SaXgbE6zhLHRv/otzQX2aaLXQrVlNuzCv87cZ9fWjm8f/ptqWdd
XuM6WfZpDGgmOFHckQz4KuxHeMykYToaou/hlUExZw0z2pHX91ehbPEAwvezvCXPDNyCunMJ4KbZ
s4rpGgn6i1SdypgoTPq5sc8dK/nIVPhgAWq5JszD/8xXNJ2++tDhio9cwyDRded6UZvxH5NJE38K
r6Jo8aVwrdCYDmDh2OJUmpoTwfI7KvBwxzadHXmfl3jjj/m5yPM8+A9dCVyTACDXsdNnUkveRyuJ
7sCU77Nmn+hxZsGqchVHYk4UMcJKLckqjKQtERY5GLz/giIWo6awAj6IcwB/UlD/lZBklcsNGU4F
ATMs2AnRoDAa6UXwjMbvG/435ag6+eC/Qn8y7FoWQsycNXIoe309g6BPwG0Sz1ojvXhhZMUFyLoS
9iIhfDI7GR/GjY+3Q/h7W5hIosN9UD7/Nnsr0rLcm7QBXJCxnkbRv52HxcoZvR86UN/oUNtFbRY6
q+6OzTdJs1G5D8hOZtIMLjrAf7iqBO1QQFYvAYBFxFWn7D8xJqLI4WOIq/A8byfrLfPBPwv9H19h
OihfT9FteHATIaRIdSIvptCVJP+4ZRgRPNUCmsHRYWQ5fAk1fl4V4b+9fOBk9nSmWWPLIv8sxW29
58knWvS2rxjbyfLeeeCXOcMXq4yhRwzCn+FROhlNIAxa3lhnXkCl9k7oY35AYaBKHllEy0rG287x
YLN8T4z8HBGWSrufpc3DTT7HvUbQn18ks59aFQnaIE7JrGoHUGes8tpbBcVeYMpbcRb8WYFJxBjj
71qlPKISvUm326HXkHrGshUF2s2+isoj4eKYABcGvR46Vd7PTlib6hoWFPqsX1k+MX8iWMHxBQS7
YqR7RGOoksbnCqMLw2OKdEXJ83vqkKEfoGOBbbUbxFIU44nPqviJ+6nIsA5Gl0EGvodLhGiDVDCF
UPadUaIdxFomb/ajJfW2X1P+Hhp+TkuokkQqEygZt6y5E5hEeMEGNAma6IUvxVAfZOmy6hO3fpRV
NfzLn+vZEsScRCA84BIr2PzKOVKMtl3YrUxqFRIzTRClp5sVP5ZxQjkh5SVI7fyXjoEbbhX4KtXG
cvPcG9xVWV+H9v9LxpUyvtPTGGtsMLJr/19k5O8neSRzRpmyj8ZcUF1vherbJhpMb+1lr7rNlld9
q4tOo+AfpLSn422je1IjVpeo14xQPjJHoB5x2w/+min9S13+7s2ycJ0DX6s4fWcjknteOkkHqLf9
AfwCgFq2ttHdDs1OXDfjDxtzyx7l0NU4LuLCtOTgShUDcISCq829ArGL9ynqXO/WuRurBVYvO9CP
zhGDbg2i8uUU77vgC5BiGMqxagk1QZczUaigXgumiI9Ce7g8EsX55RwmY/H8X5vc4bjKVwIgcRhl
weIQFZloAE1s90hfdTx7GxO7lUqwy/NavzVlwFPuyBiE1TONM+xd9OzKKlqQ2oGF4fESsYLXv9a6
Iy2hORCHtPr0xkLIrEfq2ulLB/ZOh1Ght9PpTKeW1nESDZzeK0Q+nWmrg4ML5u/RGlo9L0olgP2F
onarz9mIy6aWypN2MK3UQTsgu/8MxAzQoA9gwxRZxdK2H4O43oJZ8vnU6eCtzSNL9yV9RmCaCbJ/
Bx+dqsj5z1hbHjUmYWJ9ZxA2DMcvyhZ0fGbRRIYEym+OqJxnOJE/XvvN01zyDOxksrelIhzxQlbQ
IxK1EJv2IM1OgnYqZiVolkY+pO8TPI+8fhSourasPMyAtTAuGOvemZQcbCTr6zrIJ4ncNv9iSeWS
xyoRjHqDxViEOw9QCq2Ydto3iwKs0FKQ4KGXDZwPK/2V+XkJdiaDJrOwghHKcQPAd1iNXUcu5uTQ
uiHoESuH7L02nxnFli3SUym23hktbL9n/znMTY+vKuKaqKaGIEmIJ+uY7J82rOg+Olbi0cFm3xh3
3QtKiD/NTZj8zj+aAjaLCt2S2DvKU4ePLX7ovDvwwdL9eArw/cQI/Pm1zp/57xkCkptztBP60MSD
4lEkRZA/B6smEBj0fIdHPjasjnZAWxtIf6H5mVR4AI6/GjNPO+/cQrLdZ62KeFQr/8LDBdWaTCP8
HEgJRkJReSN5AoFVwxOaQATiGJ0SEZ3FIMHtlOnM+hl1hyy8Ad9Gv+eqQGhXzPQKyks6Be5Rgs6E
2Ou0tVVxEegctow4dwYZ/WDFR9OvMuZbQbCSQ6Ddv9/rZ9rJL00vzXc8hW/VfjJzW7OnIi6QR521
M6vCNkDLUprdJ9sf9iEv5bO4l4aqcjYd4my7LgnI87lgCbwbCuxEgoax2v9unvtmMHRK3Gq1Ehxt
vuY/08oFuahkKARktEiIiVe6wcMYmA/mCjCu5IWTutpasV4JiSfTsAK+s4ZIFYvNkNJ2xazxci2T
zbADbqLBnyWJO+OdOllw3hFUfN+agjLJ92itnsfbbC4hqdjbw2Yo8P3R3gE6SI4STTg6hJe/B9Go
4pDD96dMbOxHe/A9otVyJ7uXjUJBTud0zYSqn/EBwT67BP09haJrRkeM45OzEavrYUxds3lARm03
HM6RjsNWdi1Pw8BTASjPEapDcD/ZRFr/0UCJq5UR2jFHhwd3gSq+NcK7VXORTt0O1qS2bbXjc9Kr
FMRrKW1uSfmL+sGxMakzx4eG01GEfEOMdqV8dDD9ThBobyuDKi3ItLzgddCj44hQK99NxJqPU6ZE
Eb31HIjb3kSJW7t9zcWwcNMb59rxxeZYn540mZMxvwxmBsCDdyAmw77hGYOkhKwLQC+GedJMQFkq
hEHlFRqnGGjcGQDSNF3gDHlvBr8MlG8PKipVM+5tcrzdbpLbkU94yTOuoNFWcHYvZKnek94TCFLG
KDp7YPLvknFH0NVoHcd2NhsGc10oDZ9Ci0NkSRpAU7s0Iq0Hji+nptXUfyKIOQ3CZelBU8LGmSsd
O0/dd6p6e/leHLPwaHRLZMX3dO49emwZnOuZ6qTwDnRYMM6BjiWvZtJPpq7cLZjhzd+eMO7in5HW
zSpXVIeoK5MVa+JB2fNzxGT++vnLtwc0mx3yTOTzjzS6w/+o4Tpbzkp6ynmwTYy6q58rIW2LINdV
Jk3uCDa/YIrZlBdW0rclFZbvci4iEzOZzXat3zeOf9D/V+s4dicDGELk4xxAWaYDsi+Qt7g2Z1/m
cIznhyw4GzPNLELZHBnrJ/F6FzAEV7Nip9ECpkQDJW9x7tN4fzwrtzc2EG/58iJuJeAt7RzyCV9l
SI2iYWvooLXfjuDVNCLfts1t727GSwpZDY4Z46GMKrNiiWm1KzS76aFYb4QYFpRxjeOUlTyiEeoZ
bR/ECjhv86oCINVwbTGq8Bon04APQpGrgt1b/19m6Iq/co9qjkLgVkkwmdI1hOFDulFEif6LP4Bl
ursuTRl01qVyu1d8jXytH6aHLCmyug0wt6Po6VlkxlO/2hq34KxSOAl9QDYfowWa2PLBSCpBJfed
Jv1QSsqVzO/cC8LL/HYjnVOOFzq5mNAyxnkT++HtkTqb0gQDhn46T6VlNz0TeZukSJi5yfm6T1HM
+hqpU1kAHC5P7VWSljpZ4/uRVIw48xHzf4eyxheGnA9XpnqddAztX1mwIlp19EHxZP6pab4qS1lG
0lVtd4/yuO/tUb0N71VpDVM9/1MvvBdwcrGkUebZqMAhbtAPg4sMVJZUQQaM6Tel9g0uhYOnZU/9
JC2DYWciojYMeTnVC6mb4Xv6E5LhS4Zowlu+fmFJoxmKV/BYLc7fqATCReKVcV4g0Scda7vM/AWg
OG0i0z+M9SkfLF6idgGOGgg/GSPbkUNYLuDWEkWn6Jk+JMJH/ql+dl/vrPXFRynyViMMsAVBXIFW
HVhpKUTuR9Oyv99gNAnzVkN/yg0yvLHhLvGC3bz3a9WNel4ckEloFKzhIfRmxhfNfGj3CaLgiJ47
gJF4jHvawaEuG11xGgBHLQ6Tz3Met9QhKazOQG+bAv5EG9uqqEPKtLTUqL3HdTzegv76sGaqFm7B
ZbnHljulCsMlZvuPKQ8N+JcVcwFxUKNZsv7CkhadA5jD2NyyGZjKjJEv3TE5fOGHqvbLAWfBjtzv
LDfywj73KqcU9QZRWPzly+XR7v6/AKz7pN25Gx9CGUMmy67lDsDaqYDd5ZBuxpRgd4MGzD/msAbg
DyWy6di4hKlg6mZw977Rl+Sxm193MxR0oOdNFCfJw8aGwgfDTvambagMImfmsWH5lhYfhG7VxVCl
spX7VvcpMMrrwhg8Ukm4stSIfX3gg2JybRmlXnW0oAZrGC6PEufrmN5Gh+gQ07BNwSbue+WJltoC
4y4xEPafivNz+Q1oBengw1Lb+iLe4LzZtDJVzmZy3kp9LD5xKG4XhVj+6ZUbyCaZ0p+XQsw6qfMG
njxT/b4sCPNUDW8QGLKFtG4gf9QtWO11WSG3vPFqUVGVWimIXmO1q9/CJiNg+td8ciNiWk2wI0PI
K5rRBXRcxQieG2KpvypdUDwG/a+KwwXP+6vJF2L2uOoCSBz9I95f0FoUT5qN4CNGkEA9G3DW7fym
UFtJWeAHco0NSUrJcqfU3B2EvMhl7DBY9gNPUWsYgFfBow8s9LcbV1uKvvBuamF4Y6jYundxCKvW
N56FbufOYFUV86II4Sgb4CWh9MTJtem805DIiwEED4mY1qEfEH+V7OSWJSeif9F03p1SdIh9v4Ip
0RJqeA7K+V+1l2UulLVtNhl3EQLSJRhzJ6gYqtqyqNvoLLkaFCmE/wkCwNSYTOGEcHRbpnuVkCYO
sTnrkCZx75OpY/zB3iiZGvCCHbAFfB4KC/g3N8y/QOv9wOWZIhn7z6OlWQd6/5B7zo0+OP4uXer+
zpyvsKAXUN/ZpWxFKuBVUcLP0yW0DnGZKPy+wjqx0tg7Z6lnqraU/Gx7WOhL5h0dMMhcr4FrADWi
jWkOFhSEQMu2coKxmNJpHmd/8b4CYUrLvXDX9TGWBnnjdrYS/lyfoPCZ6/JObFe9rHot43CdEIIy
IUAzG+MACcpkP5DBskyOUIwBbLn+U5vGpvSyvogw2/AOkCvZVZlUgPKreDYFLUySZUD2+I7vFtLi
BCXOPOZvp1stB7QPrXmRMsXlzaUiUn+vcIWyYQefhFnU9s63tZAbr2BGfzi/3NrKyJR+EPxy+yRm
fr+tFr8dxhPtUUTP2vOk7e0gVSdU9xy3kbSn5cphf3hKptulvYEP8chmj+XBVhhFo1BBkdT86H+3
RNDou6z0IOSkDeIRtb7Atfa5m4jU2iWsprgK+Cn+lnEBH9G7uyp7n5mbF8nY7lq+MMhccC3hRFqU
6dviGL6IMqqAKln8WQJMmVR0v1RlnAYNwQotQ1cV6smdVTQMbwYiCla8hYWftGXXFByzeUJBGKrO
AY6UdruLfhtTShHNoyVSF6BnMaQGLB2ajeZuv+TutTuEOCA721tDsn0wDETNYweuD32Uq3dfdrir
cemom6Ij6BGVM369pk7XmLAzb0PIWLwLBGGqXufFR3SBjqAmvo+SlvMCLzZW4yMfhTBcX6XVscAx
kV4BXnQiDQmizOGNGSEGGbemhzhNvsz22P8wySlgVg90tQ2UtMB6Wtjym2EaOoP+GWZcTbXfEXut
m+vxRtzy5xsySe2ljFpdYmxUrymZ9p2mFIAtVPwM3XotE3A/nbPm1mIVJrW2aa5g/H4kH2nYhxvU
/nE2igQiPwotAqQU3uYorD8WtbrKD7NZ7tED37s20XDeM8wKRdOtSvbTyV/PRM0j4U3bNWx/5M2a
sgkE0dXYg5NfWV3SKlKaWQP2q/xt6sGCUNi8PsbEPxc053iZp+vT3if5O1rTdc4yw83u9FRGNjew
zAnrAbKMueSnahOphQ3c9Nq8adf8A/psUBZ4RV5oJYlBGObxWxBdfBJDj7B+v6y7Rc2i24UxNyof
3umvH5zVYmrxbiAMFVQ07wpUDp1yF11xkSsi0KQLSR0fBWwCHt0Ld09hSwgNms3p2pkHLVqQkU9P
XzwLaS/yQ76/bpe9/QXf1/phZVg2sAe6yC0xUQoQDLf63g6zuij9HeMd/h+0K3kiDQ7/Uj3htCz9
zgo/lQMVFR6KSodllVjR3KhrATx1BMYmqVBxqG17Q3aiLtwtx6rbh8+/k9g1qxS/QnXSlRB6Zhio
7ejXSFNRFplfKCDJDaatSPLakMz8yEmNYp7OV4cAbtavGbBEG271Zv3TwX80xLLNCopLr0rP9u4L
DVqqxLkkRXD4z/2DJSjHFY1gN3Pc/r26Uo+sMZqL/E7Oi4UKFgAVXn5XjvApQ25OwxpH2KhSvi/s
y6PupX57d60MaXbB5rpWCXO8k2GfascfcvCFvQrkk1YZrtI8EShcwwRo9GYfiWh6kNUND40yaor9
YmqeFvGGIKE46NkSwo80o2fASZ9uVOv6dc6JPxZSz1cDAIcZEaQKJo4jlPXkegdysZRCLjSpSaRT
iMI7sCHaLLi1AkAcrKh0ws/ATZ/Riqj03fQ05QbFDscmoNJLWfLmiDoXRkQzH66kPfAntKPgKFi3
MVoE+bizggIj6b253rAXxzKkBY+p7kkzQ2yn7Yv75XOjX/SaqldZitAGc7eOAPL7qnqg7KK6n017
vAgNLUhF8a/w/CF6ZbEL0i+Qh2CPwoQbFY1bhDebj/9AKVowHu1H4qmtc4Xu5hzmYC9I3+XycD8q
xAv5Uej0YrZEtyPvDZQCINMU1MNo9jdR5OS6CJvcbNCQUTL/g/d4y4rwf8p/oPat1Wa4KfF6xN7o
LPCTXZiP8ufzZ3J9zyPyeWuMiIoEHUQBU/oiN0I1ifvv0CuuJpUc9tuf0YBcjuArKEL+z9LdggtM
+Bg30C90QCwK6ro4jF78wxz6grhXSJ+/tRkc187rqlcd+b/6pJV3DrzSjG8K1vT4ggj27ViGXfSw
qPU2QAhknvvhltd7Sy3h2nd616MFRegGAjLIEN6cX5n3kVl+R+OLBbAmi+6ZTaeYcYBpg7d12hiP
OQ2CfioyCltD2nHWvpyiVhm6QFB8/0d1MZeQSKiTtx/PTKzNnVuzxgOzxOuxwpW8rRyiJ7V91wGn
LqSiEB9e6rmDAiRZ8ETDAo/8qO3HSCVG4bFtBTBWDYl0jmdqpmah2IYi9cvpGNGptDz2CnmkNbzj
JtLroM8L620+DCKWU+r36PQM9RO6cj1Oducw9tXw8t4Ighe0+Vz+t5HzF7QuNgq1/NTA3oWnQDNe
BwRyIGOlq628JWXGKZ0PV8H8BB7kPb90ibaj16w/uq2LnjG7/0itUbAYzLATyAlR9HT6WPZcDcpL
e7NXzwVnHGKlzDfXUWp1RHsz9zg3MqFHmh3xvtstDrFUMGRuWOpSuxjZhXzRm86oXHHknr0Ao/GR
DHG94fr7+SnDtacWuJlNxaelb1Q0YWurkr2J9RwK0GoQ3DDRWov//+mBJ6WfRr3H3lSWfLqL8Lta
ShEERRyIXPNa8Za2eO2qhTqtChVjY/pbIxj9YGlK88KR1c6xkDFvrGqRcN/Ivwl0EVwues4h7/ej
Lo0w2OsNANzhe6CAgA4Ji40gq/mTUw1HOf8K+JHxWxQ7qqYVImlNRMsJmnF5r5RKXUV4nmle52vN
6PjkHmnRb/8Dlo9eI6bXtbzItfiM8JJULhyFpxJWs7oUeatFnt/+KKHFicl8fJVzVcoHdufdNU4w
PV+ZsET4u+dUJDn06+Sxltaq16GO4du5afeoRxm0MwK415+nYi1hoMJ1AbS9gTOafkbXwXlHYr0+
v4IMPnwYfpnfP/qvLDuB+qA3m3OB14nkNF15MNTwrydfv1QpRZcVbSl/damvljDHW86qwsg6L8mN
lC+xxNuA3qjMAyJWUcLzEe9bOMj/hmfYHJjrFw0FDVQ/aRrGG1aJWkUTr6AmVm/Eoj7YkW4jFDBI
LXJp6nzKUsUMOtYs51UJKw2otvHJ/ZmYtGD1JZtx5jKDO1LU30JCcDRYAnZrt7UDe1k+gOY5LUB0
bn39KyYtOIEN1FhncNroH/ew/aMDCM2vOhWT1nMJWgwOBPhucnOTEsk0dqA/SNQIPiuqiEwqWM2A
iwh0VWso/eSV3wR8ZkVHamAgrZMLPRfcamIfb0xZiQ0rsPA68+AnZVGsHV+ayEAjlhbYgIGs9DQm
6sG4jqXyUkELIVEGiAAi1Pj/X/RZ/Azn0gtRQIXsn9aZkZcFjqLdqBo4w1Q/9BIz64WA+GwP21l7
FAsnpy+gp1xeq4VBCVWlcUV+dQ9ofoj2e3wsu2Pay50nidP51FxOUmOYeF3h1fILZM4FIU3cqrqb
Z3vvQRW7oZ91LABh8YjslAp33HqXnN9q+rXPqPdOHCabHZxMhrC+mj18Kh3Cym+EezqUtxDYDaSa
aOxyDZ5nOTs6MdqJASVRHNXmdH0DUO0N08IIdqnbCAmJCzPlnmePv7eXoRuw2ty+DL4P+nfHoCPk
qpKzM0WeER8uTTbCGpDB5FzrxwwppaqSfRq3/GKfWM63iJG3axgsc5iaVpi1t5zp/2PKPaL2M7s1
GuBK0zHsAk2DPp9IjpJZ+IBV1pd3LD43GgzXK7zh01pEzQWEbfx/L84hvEOoAw3kS30aqnKzj/io
IIjSp7gGiJMCp2eBDHWf+5tTipqPRJoN1+pkdLapH0SmyrqKpqOBW36b1ak3OV2FQ80AU5E/ruHn
SG+u0QpQptUsneO0wwmEO8tITCPt9TE1+66tfDS/7Svyf4qncTu46FzrzPxGJfzR880iHCVZlacO
JCkL2UVBTc4FfZkNc5XdBQGG4hM2EF8LsQxGvc7HfYLOGrGlLsfb4VvIx9S11zg2S9kdIgYQxQ2f
qQXza2Qo1Vke7m/HNEX+o6WYIfc7FTEF0iv2UMtQR6wT5WdjcMoh9ZCHUUzkAg30fRvAKUGR4bVa
TpCTBzsUH81LkTaE6QFlqIBF/31Rs2Sbe1fAEVE4yq8oLJ1JXIEk7NJzX66UJ5gqNcx5zrPA2wLX
TZ+w+4LSYm60VdVRfv8wI0ukmQxR6O0VM33yurMoiimK49KbVR6OUO84CO5+0oA/EefOrEbQElX2
CBqRIyUQ722SDWN+HXjlvWIKfXaDkSFePExktDWEeg3NLw4ZOQ/WMXU7pkknLXKxG4kRI6KkUgXH
RYv/kUKIDv9NS0tTEDjoeXOo0Jkx66U3cjOkwteGXyNIFIoDGDJvjqaqi0MjEQQ/nYlNKmGduFls
+Rk9AJCeyISP6Z09icphyWCj69w1qLCK9CoEDHzd2qWpvbn4iCE2a26jmkyr3W7liOqLCojXZiJg
p0OdPRYmGoW5raL217tRXLRcfHKuMrXsW46Xi/kNsGxvOccH4Xt/kEXgecPXVhC4rTk1UFKRuPDq
pXYuKdNsEo+hdn2ZcpDg8K0Tkcv5WcUkzZcN1yXLCyM6kVED3rX58IT5WHVtrB08+XYJ0lqN/0dv
fjkyNVFGsIFjPrir6sL0p4cKM249NRQwks9C4g4IozsvYAigffv6nLoNWwt86fqR0bQ/1OBCcw79
WN0bA5i2bKQfZR4foFoPUvLRHuhD+ptz9F4BcDYsrAeREJpko6G8c363bk4T6WLnWSm9m81Niuvz
tLBYjj6BP81WtfrAAgFSKQPL5Gq6cXVl+aZq0zHlrPYWpBsEPKGpwV4sWPy6dxKmiEvcuACj9TTk
YFrCG+vD4SIgCBzzoHDadLxeUF2EfpZ9r8oYQg0Hi6W2g+EqHoU2Iy974VWMSAvjhg2dMN5w+RMd
AC2kZ4/Njs8obDvYGJZBe2Eqq2svAJdKW6f53IbtFrKBzmxKiMIlFHyvcX8BhOPkBa7sh5L7ObAy
OO9MKGvUZA/R1tnvP1zWmmxPtrlMxWnZmysTZEG+RJAgX5gmNiRbsBBDNT6E1M7+6oyk4hLMmtyy
HEusGDPoVQN2K703rLMCgsOGEnsygkzyZhvYDTD+RSEjozqn7yT8tBNJnkyJCPP1yD8VNipfAYqY
RcwSDjRSYF+au7zpknISrtWHLEjnkNcDmwWKuLa+m2pjSk6BhGWl2tR9tkpYQag2L5wRe9wKk7hG
SYQYhO3va7ZPiaUY6Uw7Ydl1iYES5G/IUBxWxW60mMtxA+8qaQz7Gpi1uYQ0iLhsk01aaT8LqtpR
j0w1XI+/vQoKDzxmtzl0JyNrBjPBvqKLPwD5uXMkAzPmMn1t4tcxoizAPuPDMWLNEHkHPGBh3Cfc
ZYETHig/JYEdHPh2SItSM6vzLpj3EAsRWxTQS/VwC1ga5hYa65QRY979VGGnC3/RLRqvGX0vyCCB
Xj95l94aFn3xLEbo3qkSn7CDOpnaio56+7hu2mhP7L7mmNjIfzgPmpQNi49Rl+hmoVKTaQbjynuW
Er33bMGFTXISMfM5aIKrQIJbaHE/dXMyghIAJ7XMgStlmmfsqOTS+0IVWTD5WqSXZORNRkwuvs5y
5wq539C3w5mBdvP2GJPJrC0Tm61nQXFRgWpGIOwRsfOVF5Bxu1nzupNnpRl5wOQ6FHlKwSU58ZIo
qNV7EXjKGdC/SjGaxid31AHNFlthGHRSySLgh40eg6jygfM21qaq0W6vfCZmhiKEvVV2G41gu8qy
0zhfsSWJS2MITnOkfJYa9rQZVceNBIE+Q4DlVTBnNNYze6dID1MMIzX8WwMeq+GtTVxo4cElJavV
R58uDLUD8Kptmj7zYlT2AtVkUDZ1u8rtWwwXOnNJJ9niDdzeRd61QIJz+URPAicDFjD8KJBmh9eT
zpc+YtXdf5ju14PHM/9L1DSBIxvVFutbRJg29UaBxbjnwLZOkTrLDB8O8buZ1B2Hlekc4RTtndGn
rZLOrjDqoNI3cuCiGtCvogg6lnjTjjJvE7pQqJeqHJdt7pPQrHVRpzwyEJtqHxFsMzcb9yxI2JiV
ZaELXislvv0ubPltYHj4ve0NruughNkDOY93iy9K3FHvZuENm6J5FWQVEJT/kE+z173MSXRPmIwe
6yn/IN+TF21NhvP7Bi53DtJygRr8ejABaNJued0dGboxJ2D2X3Rlzp9Ay9q+td1SBRkwKoJs3d6J
YxeblonFqyBtAvrPW6n3fH6qFj418kayMsSf3dtHkC2fjv+UuioOpxU8eKl4d+XD0MISKkdfQP+x
srVnp4VYpkUEyoPS+rh8dzXv8jPDI+XDvXiuH+BqZPtSIBoN4SyUmgUwPKUePTJuk3ZQxcqTTGal
uBNDLcwVMe0gd8OwrXKsc4K79BkHDuqXP/WF48bVdt/KjpCgBfvPwHj0yeSJITYx8Zt2Ma6UOisW
uLpfZ3ZU0saMYe2lAq4QN4QNTrhbtyP7ciK6fbBnfTiy9g1YZ9h0mHryToC7tbfZ+v6mpEdWymmr
syyi4DUu79ZUS6GegaO3V0N0aia0TEXurBjJe20P2jRxRnDSoPyugaYm6v9nOj94psFotqWby6Pz
phjUilYYcLFepeKL4mDVZVD1HqRoVWxFZglN3ERsMwddL2hCdM02gRyCruaaGlU8DHaXFVD+/6ls
XYaZAq9FDQiw/sBCQDpcsprPbRIuwBkmShmJD5uNwiMxi5TaiVT9jvd5PZmu0wNAXHnKWld7LhIk
coVHm2PudsiAXYsHBTFO3CHJnuYt4iyWW0ByzMx5H21VFtmIiKwizGerGZ9ECKN6BmvZmQqEtUMj
k2g6CzmPB4ji5S+WgsKFnhynY8SD7vru2ZS8dOU0U254gxMw+wOfW/dMCUAyB/w6M2HMkz5GWc/d
ZcbhNYCad54SijFTnGY/KfJhnJjawilqnmsveSRKUqgdo/4boL5qz1dFLeOX4oGE47/Li+qOQmXM
GgKYpqHvXpkeuh4qReb9x5iWFKtCdNkOhsI/Mg+CuvbL/qqMMp9ViVIrjIGi/vmdVj1gBJ02+Ke4
oyHKYSk7xZaX2ZGkiIjhNBN1oyeutKfJGM+cymcvQLZhdzwjM92d8MHGDg38x2C0jQKt0MFwszLl
eWNdBqoAWxx4tf5bVGTHIXyycRQatO8l2p7/pxPMPl1NL97XNarb+umi1eAIlvkacEII2nFG98Km
3aPozphDh4H9cdwN6fWg5c2A+3KMqNJs6vEzlSylYwT+lTu/aLZnXOKbwQqvpZoAiKxKmborlTe2
XH2K8X0PVi+KMPm6qjXevZNStdUHqz0MJmB6PYFXVJ1h2mHt8n/32o3sFFzM4N8sCwQ7aaMdfBiZ
JD0YpTDJUQxlT+PXKlKsleyFzeLsSZGQn6XMGM4aPHZzzlt7rOTNIk3ZZvpCL3e22ErQ88UN4YFQ
CV4wSnF24CP+cY1iKdyM4sG+CWmUsmN0xhTSGM60mAPyUm03zAYoyxIXIjQj4svFoyXyDi20cCJ/
umIudMk17UbnkE0lJtChnOSGWt/MPyQQWSRi8EcYnuDg70VJeiBzXFJuZwobqdbQ/T8j6YF2EC+a
JYRvry6oTWS7MpVxnXVe/as8aqjJbP4yQnwFDfAwG6DjjXWNf/YXErLI2EOLEEi5Z4tIXIA4FW0t
WAicj4La+PuqXSRSrIsY56VL9woNlRwktL6009oFt2zsnYQmIfB0g43wUL4IpLAkmWEvZYW1EAno
1Nlkt2G9rRpZ86+32sImA9ULkiSFclzlPeVJu3OW44bZi7+VCuLuNKxBteBJ8jBt70EPTtzuBXmp
DixJcRzRlSbVuVfCUctigzOoPKXmdsLS0ZDUeiCo2+mkpiQxwxPxgvukQYyldPH40kCYG/rjWzcT
X53kq7GPEzEtrm8D8h08iJNiLfiT/OfAWjgLb+Smx6C9yIWTJLwMclwBC++x51V3JDWhzMvLDrmP
ihJSm3KGI7XYwapT1ULrrKht4ZqAibZ3zz9kXl2aWY86n5ttedmLAwXG5DIyjj58KNokw3QIAeGo
atkUcdDwU9AOZuwDeGaVJBja/5Gra9Yp0Z2C7cvoPxF2mq7EokJd/oLt1XYcjpfxEcvn+gKu+/Ri
sVxxVsVrg30HU7FKxyYszUr/qIBbkBDbhC9kqivTSEjpoyyh0dcPk+D1VTx1DsOGzIXOzekH4mRC
Shb4MvoNUHXKkl+IMs5xregbeeniyhZbOTEegAk922aut4UkSPlzD/JE1d14KvWrkjePtcnuHBC+
BraRNyZTjfpNv5U0AmoDIwcg4Q9agfOfFQ3SRNq+oqu5KAICAt6awEGtJX97rxESBhUSCAX+Rdvb
RxWmIPJUDSnKR1VWyrGOzzg8rNxuhG0rMLpAZOoo3yRL3+RcjFPzYTEBIoKVeX5i7S7zMLEACZDs
FQpJ3ne2jmbDMwH1/sZy96vC184IYf1tkInghDFgUCsoHQ1PtBFnj+od/2tP7u59yf34sTm0/GbI
qjKBqkLA5wIqlsnlMN0M/wAqfCPCtGX5e27EbUMzSTrx28x081Ez61zX50heG6DIUH736P7s1OL6
oqu+lxG9xVGZWyfgp8Tj6s6TqfZR3UHS6AO9nyZlPqwkeRsq4jEmUQoPl2lxzCAwy8tTj17oPuVK
t1b9o+CRVcm8oQwMe/OK7e1GOWnSUPnv/2mt60e/c1YuTw5QcergVQO6qXFPKOujQO3shppyi736
G86TCWN3udIUi9EMoH4ERoR9RjMbgktkoPw0Bj3f0KTZgEoVC+2AQSeWIWCXHmBj/wGLhuQ53Mv2
hBHrmVIPS3RoM+9flQHWBglLT9H+aTdIYvRAgCont7iMOyjKphXq9EtQWYy6E0qmiFXRoDKTQUxw
9amjLrMzmJD0V33kn/XXDwz9DQ7f384H5WYLoPCPW9NZqsAuIOZSSTZrjNmxjkBW1vISf1LSzHpL
S4UqbGubHs+zqkmtIfZmZdQzTzbNiK3lbyyvCTVTNIz5c1GYPSI1OtgEom8Fhs3iebXyZweAPPTk
uY97gHejazW51fxOoIjYIesAUImHCJfc7pgm8C7+tYhOOnGYQKPL0csaSrFIHCkEP8hrdVxKJBce
Zn5oGGjqWWbcV1T8x2Ys3gTeWBigoJcw0O/YzU6QRKN/0C1NO5jV436IEEEuk61xf+vS+yICw0ce
xcwKxfXwACT5AAKf8LCdCMW92SzKyddbipK9l2/0Uxz9ziNQSJoeiAw3gQLruebmjx+ba8VJt28u
F63+pMMCcc4YhTqoxre7QSyu7oMJ4BBGtJeQSJaUQWA0b0XUXiBzJC+tYOPeRAXadeEKJ1v4xlwV
vR8yRahN2scIlR33SUHV45x3VF6xqhmr6hOysH+7ifLXs8RwuKOVZm2cw+b6CyXeLVGM7iFvdSvr
RyhLzSnJeman9fugy0+LbPBlrQRzVt5RCOvolom1MV7FSakHTh+EMtIs5bk+Vi3mNWJCdS+PxT5H
2ljgcf/m8cXMAPXCIowpMc/pCzpX/21r700hRc4+cF3kJL0PANF/bNy3BcdwdrqdTrVyCGyWaQ4Y
TsqiOTpH4jsn4KgbpxkPgefE0y9H4gncI4n2rvakfkWtUnGFBqJA7VMVf/rzm76cc1rXQrPD53NQ
kVPgg6hI7y/QCtUUtMaysRMK2ok5D1rJp+G9PFcKmqNZ1RQmQxkiblKQJDFTdYdHuAWvIgNTr8Gs
4ZxwuIO+Ww/y2cv17VNlszqdD6jYCloP1qBoOZdxnhBC9SVpfrz7zPg3nUjJkn02/HmoQq/I/Gwr
YrAfZUNCksb/7PGqFV9+Eq53bnxi1OWqvTQja3BCYnuKAURQfEcg9VojqnYSW0si4L2jmz/xZmZi
8O+Q5YfyB/+/v1EoMB+t+7wvH5ztOE4qN+c6mIRErKpnozXyEsG/QAGFuIptzTPpSjZ2f7WdUrnL
LYEQvvtbX7eZff+Dx8LGnbhLkwrmO8Zf07JkCpJARnE4PjtVipSgL+7fnKYJcAaCi9Qf4EOKJVrg
ecJiWRLAHD+qZJaFVqt/PavOWEsYCtgVnhNyalNBNVWxfdj6bMCDDieXNUHDOR28cKvFFRt07QZG
NkCpdLLjwTj0ja3RqbcBEEXjGxmVK4ev/iMCjlyVKLRFPJXhjYlkXK/ZVTRCYJHyuLJvbb3bVNr0
cN7gw3ty1MqAEySbDxe+9lbyMDdEkOTIxr2CDULG0ykn/M5G6D1oJZoASxY2q6nj1FvHXPrXGTyC
LRbBKKLN+8J4X95vwG/EH0TKUe+a0Jn6nS4S0ieV8yvRuZDnVYQ1v2ZWuTRwkrMQkCJ+dsEn3gE4
V+zARF09487vc3Jdy1GrUgNh8YQ+JafdN0XbaYkK1e992BJCagD+B+i1TMRBbGFHWFNFzLUFBWlz
KAxWsCQesjzXngi6F34myTT5sexOFNzKoFqwO6a+80g3JhIgF42CHy5ax4WvP/3YihQ3DUn5YAjM
CSEUNBKU3u0YTM2n9KiK9HFzF3BYa+O6e+6P+PhyaQT23Uh0H6R+OYQ8x2thrzbHkjqs9ibB4+Ho
bSAw2Mq4WkuK7Jr2wKh8hM9XuIhajQUsN11OqDa49Ig7NWzb7hmT3PX1gCfF7D5v4Q5QqA5+XQcd
vH4GdBVE/qecRTqmwLASZKdM0RDLzAdXmZg7PMkon0zB0EmoW6UoBnKar+KVuVHylFckVohIDsq3
jT16K6hh8Hhd1Zo40lYam/MPSV2EA1iQb7ZwvLsKni9dQe6+kpcvQ0VfkXb1eTcopsPyTc+kKgH0
5vt2j+KN5uBec8j4342RLsbseNNwUwwpe8VAHGeTJyS9UdwXBe3L3uvYbjoLBto2mvjCf6nyhz0N
PNtP8dYuhpQ4kbIHGD/xNsafJXwTL5o2SQgmM8bNfx7ANHC5z9MI79p17Be2JSVixPJKvH4MkExN
4tlIX8KzqefhLurzIicnHthIggvH+OzRw/kPJzBiO3gR9ik/MMkaqm6FvpH3BtSe8L5pvw129YBX
jZFsR3pHROMymKuFOl6rCl3Y9ZOYBBhPiVscf5FhIJvxTrSAHjUotbUgu+56BbmWQe4v7x2SWm8b
VLfdwEU4dKZaxd8G9ewSoyENcXD575dkH2zjBHd8+mb0hIAV4K4per1tzKAIuMqcOF0lYcQDEwNa
AlZB5pj86EoSQj3LvMyWkfXAbj0+FZcs2a/Q9QQpD/Uzuaxrn3U0b2gXIwFcpKt2iLFvtQ+zQSXL
gmKxJZq0eN2w/rl8G8sEJNRxfCcj/EHQA8pbodbzfr7S6va9Gupg68LWr3Jpu452PNmDDWZOQZeb
4i0KyoxWsUyWXYYy6cXB63gI3myGCFH3wxVZAYdoabqV7/HvNPcqWBcvBLoVRdQ7DlL1GGv8YEMr
qdEyR+a+6xODnwMRDVX+Sz69MSRZH7SZIGl+aKSDfsdVT4bXGudmwhYhD3eyujlZUIaoXSe7oqGy
ZF0r68NJ/RuUiPfslKCIN2bSrag25W9maKEICe+hRpKjWBavvnbwFI3O77dngmqAQS5Bl4c6EUh7
NYilOHPifgmFZ6ixEUXsIdsd6oXuDMHnsUbL3OJoFVQvuVeSv9IFSSoNEE3AhEsaN5eyJGwr7Wlm
gJ53vdH0+open4fTiAVd6VC9CAPDQjvGtkbIkgO1mAoRBhGDk2NCDV8pof2NlHY+D7WvJ7WQ2lPv
fkBbgnK6ucTNYLi8AicmF3C7+/KokqY85TgEM2890S6Rh90L+ycbTM6q8E1VLqcgo6R44NLOaJfq
isM8ruZ8Jqm9ZcXp1BH9JRXV0Fp7Jrj0qswuKybG3EdPodoXm8MCMKZBxxhzs2yzt5mya8gz6ZeQ
Z99zJn1ig/E6RJTPp5pkTjl9u69NPHlUzXBilrZwG/YeVMJzK9T+L4u0LWV56wwWvwLKOBBrNzzQ
jsq45pKzXWIxKTLFLZ/j/WKX89MZpRCmK8Po2DE/5+tUXPOq7yFKQYxtfGtPtnmewz1cJW3m4YAn
w9QHP8WZvVqDLLLGceMOJcQd8V4clrFLOz4eYuHM9KMfMpPT92N5XrAsuBppWykQQqrVsz3RfXXT
cCCaKXA8XGSlTJWjUTcUOBEpYDPVNiiKZaIRN1klz0CBLFzH/KpTslrCU8PQHvAnr6Zi5/Mq9I6T
Vz5br5UA9wl8dl8LNg2PnuABK83Bmzm5GYclnLtwv4euYtkOes9895rAgs4Yeb/AwNReryrBoe4X
k6jCu9+tCBhLgLViHyrrIT4i3IVA9HKvE1U/qqoy6/QUN+yFC0uWSIpdGoKNh5uY2M7pKdyOjDjf
BGRYoXnl+c0bC2+z7AJ2i0vOppCqkm3EkH1eH98lWuqKFaKK8CDIl0OPF7MB7jPvW963Z8CrXuu5
GvhXeuvmb61HBS0OXhP9enygvK4q+xgN8f5/ABUfuf0BhL7sPj4iEj3Uda6fImLSnkwpL4G9phFJ
1iBeV7fClHLXJdBhC8Y+SpGoTy5pTgTBDuR18OfYRLkYTPg4aDg7/aTb0rYXr/6pHyYlqvPZHcSx
EKi3bIPhYQMJIigmvd1fD8GX3+yZfe4+vi+M9aM45r9T3cS4T16feCj17nYxTSCcnmEE8msIsOgY
YyyqJT91M3BzY0IcC0icZ9p6aYyhS03Avvo6DoZdy6gmzuoJNRkc1gRdHNaMAJN/qsa/6vKj/M8u
Fi0CIdFGMrkxPPBRGi2uECp6u5NAws7JFcklXOflr0/lhoRaI7k0ngJ2dnpZwutSfwQUxmKcxLoq
SNR8Za0fZqWYYdHXN2/8mGicXhKoM8nz08RfioZf4GWrfZV19Bq/3cO/Xly0VvReF5bYPmiw15X9
WPPFh9FRYH/sT8ftjjPMX6xhmcS4s13NmKejZhkZOo30QYx4OE48d8a78TPDGSTcSQTBFyAARek3
94YuX6lkLBZKJw/dU4umoxWk3waAjyLAIXR6ooqBMK/4Yd2jX5TqqksFfCK6hF7Ew8srk2A0vTXr
qyEfVHcYrnw8FC+v468MdMyN6W9E193gb1iRh6bBIbiSGKf76WwD/8OZTJ/1tiB34Smfg8cQL/qS
fZvTt3wqtMmFrnXHNLz+8Ptx5lOac1myKyH5hQwHU4jipIoQUN2NmCHaIo57go/1gkNfnXMeU3yT
p7tEfkJMmENXXfhDUZK7rXn6R80ugOruTXvSLb63s01OxFpLBByY4GqYcwKWqYoAJukWGDLJCT7n
MsaxV1saCwjc509oukiPcB1ozqKK/e2slw0XNQMQ/6zzKCJ10TPY68fq9YUjs5bWPVd66jniLBMi
0Ryp8RmaUzli71LzZiMt4zV2nL1dT9WBqSJU0VwLE+sQn8wH0byMUFGLYz5rBeANP6/5JqkBltx9
yHleU8VBVeL0Uslxxvxu85M8Gzv5moKuEnFj2/0MogDx4hl0jCt0GwM2QRa2NsyIJUNlwmziGFFW
XKwLV5M2HhE15ZBBbdb16y276zkQfNTeNbx9byB+8IjaRiuwCM7hcSv86mPw5HoNmGCfdklISgMj
1Tr95/+KwzY2EmJf8kPnblbBiPIcJAWNugalQlJ6tm0v/IiyVDEEk47mumjPKOrFKtjVgaapdYNT
9h24AnWF4j67URZdlbIkJXXpz2lAbm5XRFxuvt30DJ9SfdUjCU/fJDvGzRe9REsn/EPW1yCU7b4U
b8u7NFDMK471ZLXaERcQhesRwdKBMnKPWiHtUPYUySyMd9ADTUOorBB706O9OIcA0vYzOvGWpor9
rraJlam3E2H34I8wB5H07YtQ0KwSnPYseUYX4qtOJVnA369JOl0O4XRxor5JYe71/0S97AR3A+sX
OV1sBRR+LBCutH93fFZhfaz0nDu0adxq2zBjhZ9K7vh0tcYwTsBRkI15vu/mZGBuMj4r5rkqFvnx
B7JNVRPpHg1Jy82nvGDKglBowoahfPky0xdMo4ZzFgFDLCHzgGi0JCcha19Dv8g2fNIvpniiNOIq
Xmamb6QWdjTrTbl8cvHtbCERcx6H3sWYmmNhDPGW+4QQSn+LrPhIrjXYPaPQyzsS0WSYW9f9xHeK
rqlY+ZJs+u0IScwtjblfhO3cHD6NBVhPRhESerZuoHxjKtB+Rx+KXNJ6zuGTvlTd3/e9620g5Yim
mCv2g+1Blji9+13fABdwZw+htadrt8wy5sXCuHrcMyi+z/kf88SBCow2mwYg1C0QTBCHL+2RBre1
/FUMe1p2RpcSPBE0lh+o/Wml4LvO3VMa3d1WN5momaGKa6VlkPDzaEO9pSIlKTtngEgUqP9vi4Zj
ng7DNnAgAWV5VJzX23ERFCQZSaB+uvSjjE7zB8hpN3/WGyEcZJwFpmKp38XfAQiXQ5tMXOxWZn9a
BNaT3mzqrvdmNeti6IFDl2t3thkfj3JvbZeS8VnA+Yt74nqG2aKEP6U8AgwSkv0U/BRDjgSlhGEp
ryPH8XAHJMrFyX8zWQSsJI9CaS92zqkj0W5iqvT39T9KoxEdl5NDoaHprPcR10uQy72a4XOd43uB
CPJC5EeH4YRe22i2L7WZEiOWvOBmpnACFtlo0Hq8a1/k/Ex2IXlabIkV7K1sfmSkGWNIhh2tfeX6
QexaGWjwkkfqPcRlN/iDVn/O9DOsUQfHh/9kecv24kU3aZFFyeFJhfN+4tX5AKtPCS7pcKh2nxiG
IN+hgaS3Y5IANAmsIaMxl54ZYSGiEPyoFizpCPUscVDQhA9OrLSABRqhRApJ8t/fE0JTJRi78TJD
9EzvnzgFHDol0rgchNjGNVeocPLUs0g2MThLSiqFnHsc1yHs/m/NaxlEiXAxNEEitEfHanrAH7oP
BLJBKyD4jtqb2vSEZ5fOqD2OKfhCEWOVIiWjQ3jRoROAscarO4HDfuIOOVQqV7WsjPUxHFFQW8Hw
m/Q5MLBA/eNylnJ+vNzXT/g8MnhR/ujPRgnlh7iPd5KX98AGr+D6P3CWwnSE2iizRHmZBE4s1h5a
5lWyNkjePyE6IV7RgBRLM88gykcOxuE8iiblELevmsfGtsQysJLEaA7mQRORb/NXoTj3m07LIh38
h5ZwJXPiJTk59BmwPSUAfoV3HwksCWxxP7Oy33WXndKm2x+3Sf5EvBG6d88NlQEmKLKly2Nespfd
7LRzRlCSOpzgbsfVveUGHTYtmKJ+F+1Q4dSuEdx0qHNDc6ZLLkx2Nt6EU5O/YyV63H6Q7U6tPH4F
ZZawln591th3dUoobB7bmGJkOgAzGHMKEdxsK15V+cFdlbQ00sm7R2aSiQnRTRiP18bg7qA4IKqg
z4VhLPGk3gaV6ADxODKh35jkZ6G6LUt+yCl1oY2kfSmkiy48PReczmMVETV78URK+4Moe5LZL5Xb
vB3ob1dlvnYqqU+iHrOu+utm9sIVQdjdShjo8+b4b7WosYLRoIVEaMXbKykBybcvzzgO3pTEnPpE
FtjTrT5zaUvsmK1X2/sctgbUzvT8fwsRBvGIzjjZeLQKCN5cqNAPpKgWLm8wsWubUcII7dBOIRMD
pQQsDwPqfddHqiIJtE4yoCjpH8+JN+QDc9FtxzvbDHSQwUI+H61Ff772737c4YU+Lkfr2Z3LTwnf
1HI2PzZk/KhuhFwrTJaONnEGdajjZqUKFs58kymR9EENfg3krnM0/ZtW+WMe9OSoahWbjSa0Z27d
uB8ElPuT/o/46Adw+kLHlc3KEL2NY5DpmdZ2PMeCe1T9qz9Z9+bh1kPKnUnPcekOHnZjKv1czwnC
FliqoxNp1SUDLuk8+C/y5Z7WZDsBtMe+35yDwIhWENKI410HKDWcrQoZNPmDBreueWbUdg82OEqr
/djtcWWgYwAmQjH8oj/WVLaMW7+vkLpeoGPXD3oSKFhamY+0p7Zg919rHUYKNimeKfClHU+Nn/6n
5NmqwftVhsG5WPc01bSsMRfI1haYhH/y7tEZubWOoQP+GNMO1if7ynCWB5Al+xP3PNP9KwObHH4P
oemgYZr1wk+sXTQ+gBL7HlTQMKQmj6cbVqJW8yAa1pkBRMYkfbEXFVPvp14KKzwPJrAApSn33qUO
jidBoq+EUn+0gxZZ3dFYGbp8LH6UB8RZMDUouNZBTsZXE0zBXIh7sd1yVRhxNhZKJE5Fx4IjqM9q
v11MOpcVhKnpX5TiILde+A8cUCpvwKZovra3mGEol9pyR1mixYSJIgFgNdDTxNm9kLB0UvmNJBKb
jmXo5s94CFxZFK5rwxrbzCIKVXwE7tlw8OmiDH5nfhBcH0DP7O+oFau+rcX2fV6dVvgOXx+gme2P
S/9rz/ia4oi+oUqpNBP4ETcsbgAhG1F8jO3MBV/7eHq+6W6O3myB8KhhChZin/erdqfhyQoX8WAr
3SZbef0HjqAKOWIaHIN4w4+qYuXpWBwen8bU0mVQZBxU39LAdRlxSBCLKZTucEa35nTRaVwEgl5C
Ntoucfg2MDLU57EktP73DvjUegIqePaO/90d/DsqttkuBaUytaOZD2MysKhH3WPBygNq68ZDbllv
0tLvSN04eSEETxIEtG26UpSB9Y0saueqhuryYsnzsjp0IWZSOgseFjuitwFhwIzd60rTq+th5yT8
oFxAUmDqfPnkYVIFa2v18hipzIuMzC9qSmhOcXZ0mzEgznPJ/bHXs7EHWih6qwNZuGbVLDYw0oB0
K2xUgrLwuGP/mHtweVJW4IVqiHi+1Nfl5E4JrpcM0hQkfCnxQuUynEdI+d7y+AuwvLgcwkfOPPWd
2MeKWU/eduyac8dTG+f+zWsXnVjWZ9aIqpEV06adZv0L/+cMdl6T747YL47yiRHRmxlkG2F7z56J
XpklJAaTfXW+k8jExVer24wPZtXNHQ4oijqmRpP2llbuYcWOOAJYt/QeGky0mBF0lFbhJs7/MEqD
I2mSbc7ZuT9qJwgIQEvh8tdwSp0YueRxyfg3tMQInZnXpAPAuC/hxsyIsyLpngKtfQ8Zks2Oh61w
1KfY5FRqVqLgO6bCWCUpxJ4PtQnisyxhSIkeORrBbeTDNMBKbXzm0kcaYE4RgHnfCl2m54ADfV2Y
n8HD5gKl7D1bAqwWaA8AJ9xna2Y+RoX/LSwLPoi0mvOtWryLdgJ0v0QMhPRie3QsUvB2UN7gJpG5
RfYHWsaQ5ycZ4kz8oGAN9N8UQE8dV9ch7KyRvx1AurffqIc0S+lvGLvOTthBUKnDOoG0TRyWZ4LD
0aiLhhnt/SKNuoB/GswEJMwh4fmp+iPs0C2dqlGZ1F0XUqL9RdpNRTddvK/ZTczQ3ggrqzxiW/LI
WaNO4mqZ521UDNFds/iqwYcSEwjBkA4E8uO8qmPN+DdjoRYVRHFegafx/RkKWNnHymwvUpdqC+/i
53HcCi4Dir4E0sI/iR2YJCnrDbDf/eFN0UVz2KEnUBIHXElMTg5qz+3krh+25iiug/hTyFj+1W2g
9SPGrp9f5Bcy78DPrh5+IfFm5uCvkghZHzfGf78VfSj3mbo24NIzXC20rZi9aANurDSa1p5pU2AP
DAINMEppgZMqvtW88xVUD5fTizt+zXKf5pkUWion/e6XxocvuJCTZLdOV/Rx08sPabGiPMYzHI5a
4PX5t/rNnPJxfekPAaJaH+0IyYYAqIazB3bEHVjSw59pzlONYcORn+VZO2RopyhUDCYDr8it8oJ8
FiKsXQQk801MSU0thQUYFQ7G2kXIDHyUdDBjjDR27qKZKCLDovsbIlE87lEXSfxm3iyNfKpC7C+/
kDPkZyYoAH2zXsdET0ZtVFfLOiI2TCj1Lsn2XDkHXZi9BvBGn1m56z3uCz8SNAXIdT4vq+g8thxq
2L7K2b4fZrN+EyWLRuHrjXYO1qNlFQwZ8cM8b09g+njPzcuSBWI2EKuHn04AjrYPM6RUiJVD7CRe
/COBZ6hlhWI0+vgY+14gB1oXX4aXfvtvqi+6GECqRGt/lv0YECmfiAPIHOw+Tz7msWDsLBpKP3AW
pJCXrAAnSr+ItTl04uowECyM6M0/CNeA8FTUhpGMR5HZWnVUUS8SA5QCPqJZkDENHaNTs7Bp/LyZ
DzZch61vuQwf476LyX7ZcSA20TxqZbq7QEhcWX7L9ZjCTCI0N5oHx6mcsP4gZTxXqjkQxMroaOx9
/TzJucIYcDVMGWk2rxK45PuZQOs2lJ9tY0arZ5gBnIwONN5FAo4CKEBzlFrI320vxgPAcrJjZBqg
cHv+ZGo7kyYEz1tWwCCxo47nXh8q9kHgGtcCvRMVrG/Ku9EmKczGiR+DsbYoh2aSs1moGvAumqvj
6WG8/hVh//CWGekdMZd4eN4Q1k6Q8r2V6FcKFyuSBnIQPD6Gex98r80D7CLNjuQ3Z+vrBjHEvmUM
vkfVq+0OFKrVTch8Ckb9hJ0nAOtuAHD05uh8udjUhRRVCTcaGlOtAVf8TBByUW8VVPzYA5jF9uFx
BuHb6IJthBpQt4Td8X68KsYe0cF2pHTn3zmitlJj9GC3c1JwdyhCt4zCrMQOD82YTqvBWLnvUGBm
UNz3zSyyq7SSY0DbbT4G7s6MirJYriAl0SWIFH57ROi58Jcl7MKEGy8f7uEZN4X4YNyMPk21m34A
xwducxbUVDln8p/VcIZ9E2NK/hHoXOE5kihlmS1M1kGoAwT89YudtHRCt4VZ2TOYvL6olD2fmmSY
cWUY5IVIxWiw8bA1IOMRUrvDJikC4VYV2sYeT8qXzdKNVcY2ZuHrkwPEmJ6pLw2LPwal/SDLrGRa
NzBlx4tjjO0nXxdqGJZ6BM0vrFvN2oJhX03MS7lE0QnolQmwWGvKu62namxQrY0+7mZ1a7Uk+X5W
QPdaHYEOgxR/RqHtuUpptiZxCJ8pulXQEFW2OCn1o/4D49nKQGtt1YOdjBU3/rFL/Pm3HX3d0ONq
UboLe/sr3MMsLdO68ryBKeLc3DnGjV3KF5rM75Pe09nJZhNvwAjTMz8BunzhKuN4Y1IdbzPTtqkS
UyOzONDgaFQsT7ii2kEuc1Ef/hdVb4n7A/5zTTtDFo+OXD/VqlYIGJ8ZLAVl9nqFUQruQtoory5Y
FuuZgcayo4aA0uZ0haqNXIbBwnsa56pWjeal9AO4F4RPB7jOnJaYGE7w3RGRtDigF0e2HMb6tiT5
rAi2G2rQaTfhp+5hvFH9A377EYKwWy5qNOAL18u08vuadf1zW2EVaK3l3q6lZ6uiw6oFTMevCru+
Rtl6S7OXq6EgBqQP6T6h1wa8ylbt/H3jv6vBxVST+qzwUusP+22PzkxaC6qF9Q4uucdKplVELt1k
3c9m0hSK/NDwfYoPTBXvWglaoBbOiHcdGAtzaszsHJxgVVqU8vL4cTy+bAr5MgH1FhgPFIF3hT/c
pxyeQJXakPaCe1hsNnxru3DEmzZc2oywDGFIzown8ZhbbujQ9fuM4bUGi/M3qnDDOoBD8xIAJW0U
xvM895iVHGpAqbvgKrJS/fjNydOJJ+f0B8b6t0eV4WhBJQCcPbL1yhaYxp67tVahJqESeo7Qb9Pw
TwiSGpZUaJRDowSrdKvbx0v+/kYzFp+Skce6TAy2Q5LW3l6mjANVa7jIftdxKuTGbJnZrm16hpuS
XNlZA/R8sdDFkI6q5xTEDY4BWgJbtc4bRD8DODtRs7zjwnkJliSKHx7iRGPMwYZjBRK1DhfnB3iu
mrTQn5Mos+1tbR2v1N1g+4Ueu9u5XvcUuqr0piJgpeDShI0qJxkboptENF6GEU3Z/OaD50fAcyo4
tZRlSZcBI2f45UKSjJfA3WnDsVgOOVfI0js067cj2aWfrv0De03qQgTZBX1HI+e6BC7GkUpQJapw
bV9ZTDQyZZKrkGai/B7yXucrNXwJMxQk+bcZUUgNG8RU11ymKfF7ZgHKWCY2swQUl5G61tHcmI1V
lZe5zo//vm8RiZ2BLt95A7IOBXy1KNeYg8Lk45Dq21XdcYftlxqLzpufVnN3IRvY6QTyGxtF6VCu
lWVJPyWo2pz7W+4W/DgWUuaC9eI0aBDvCtXypzbHvnYB42G0RQZP50B1xIW5Dx93I0vwUtwKNHQe
TXp0yLJCi0y6nPv2AOOV/Md2iWr+OzPCTuVIGiqNpF0Rkwt36fjKzQlyH9aBBqtadeg6qD7+QiNk
oey9UtD6aorE0HgL45gHGngGk91CgHddwBpk0yXa2Zne+nWvzQ/Doj7cShDwDThqEWv67catuEG5
cZkuJTXsEClWW48rXbQPV/W0meiHW4/0e3wyhJYRi68nzU9zvXr3F1iAHSmufuU6wrbFsYOYwl3K
Dba1qtIyuMOJd1cS4DMdKjb2IsdoX6YwGwVIET/V6Qam8oDOtwlQEBDUZYNeqVxcVMd2uiLlhuNU
Ieln9bT3UCEJ8BcmVKpgM42PmxLhjlUy5cGWhzP5bS8lNbxGW367bdiCCeZ/oB/nakdzD/2rMBlz
uBv06HqgEpSRKBlfjRq+k8Sa2nbS13WzY/E49EITB7OrsqYo6yq+Yv46Bp0YgxQUY4YrU+OSaoPf
g3Yl9rgkGM3SClZH6owo/9BVPpv0zxa7zdk8lYwpU5yPkbGpFfptdw0k3k5tAk3EDibXRDwrtrRV
W7q4fFfKq4U2JAVeTtKaoVZUqXgADKvv6lXAgE+hzrsqJrEyCVAM6ctQ2IVTngECoZc7bUjfQ7tJ
l5g4dhNnukgCLCrJjnAABRy0ke29wSUpl3j4ivWmeOfyt7TZ/waH+yH0hpuOY9VNz0dpj5EToZgB
4jg+OpuzNXzD78QiFJiwcP/j6m7fUYOIEG5sz/EnCM4NqYAZXxhSRsJ78Rj+JVClbzcdd2EC+dD5
MqSyePlrUaU8RFphIkOSJ6Xxc3lat/pt48lo82Jf7wC51QEHKdiguynAzVAAKVnq1uUL2qG0LVcG
NklpjLB/ipX0n1P3NwWa0WiJwzdrjjJqGTpNFyd7KXOJtM3AXaOPo9SJWJnx0KhXB8qO75M7CB8b
oyDwZzhSFuboH69/F9XErYfMCgxajapqPyC290l+sp8gVUlcNBJ04VPtZCCjfd8ALtytJwjNy2ap
bd5epXssyCKG+ZXGinO7j8k53GELwA65awTQSiDCbLcuyJ6QuSV9KYqyIcS9l68ZkkbfX3nzJ1KA
PghMQtF8qbG30KDOgzn6zA6XsShi58I4fweeUFC8X7AO7+O1/A7G6g27M4DTRp1cXrwSh6RAGy09
NxnX8vKELYArEB9nQ9E/HD5TJCnfpAqJciwjNzCvPM+4uz/Brvb2FfUvudeXdR3wlsGmXP+5do2v
+RUsmgeDxni+HIJy9k7VmgMFFOPR37Yf9l07iDYrimcqhcNMxQsQJcv+YTNogC9RFAV7ubbTE9pq
KJr/WVHSlZ92xlVs15oNcb/Q2C9g/h/uAHwKIglg0ElOuad6xJ/Z2yc7PqImKM+gnGjTQM1fpc7r
K7n2vhdofKno9XVJtZ04zj5hwAVsfeayfs4i7v12heTURGv0xy/2RcblUfMRsILaF4PvQ0uf8ajm
PU0N4pVwmikTrAgh1OdKngrdYbkFaPpdwn0wO6oFglYtyBCY0MwgPAjFUAstYLtcgrSXgOU+jaWH
2nstEmG+z0TSvkim9EJdcxydNB99ie6JvjrzjEk2SMFtAGTBV37vcenWeKv43e9tBUMnMf2AqeRn
JQitx/ZCkKlpZNbD0W4Q8rbzOwFVcXA0H5Slhn9XcytDTyUX12sGGPrixvHrSn6tk5q5yNf33AXs
r42P3AuLW37uPgizG4anvFTH4kjmHFrDi/eXtl2Diojj/TkY3rVFuKt3w9w2g17EFMvpq07Ti05Z
FEx2VP2nx/woubHg3V2H33v4Tz9YVo0KslOuUC4xJu3YALr6IbPhBOx1KlLTN6ZtZ2Q3+TFlREpA
2qhnhAIgrvTgDfBGE/KMggHeWHzJwPXLyi6f9uKwmsMiWpSEeMNLT64+nV5r2xQ7OwGiVn1ZDcsW
W4+Q+LRVAcJMFdOQd89C35oJJofUm5oeTlqwa4hpKdELjgpUn6gSJl9emHPJsmcpMMMB+Fxt1brm
9A+E/mqvuPeBD6iwonCbtNArPMxckVFibl/82/NsNEAb8zIVHpLsf/NbidTPLoiPyWi4MCjRU3ok
PBudiWc+trI4/WaJlXdazSObLY7LxxKkS1Ew7O08h4zIE+2I2h8aJ7C1/+dGmH+SbkBgZU7wdSZu
xAre/hRB/m937L3O71qJesM/mKibTSCjMbaj1lvq6SN4VJnoTJs80xqAHagGOKLS5zHZ/i1T6bPV
i8YF384lWAQiJCIwVZGtI7XPMOWjgHDUXzuYe5DZlTtcTgrQfeXctj3EzwYyqi8ifKl1Ah8dEewd
KBsByLcyqEZmKPEA6A2xDz2vJag45NheHbXIkhQokmgNw1MoLhGSzUcR42CJAmpMERd7aLchyBG+
nksuQQLRlSQkkrk9J5WdXB5Z9wNjLD1IBfwZo202aY2iQAsP2EPiIQyNOHDQeo7SwFSzr18xVFBq
8sjHkOhCM1t3OvXbzt7RxxLVgXuh7Puj3wpc74vV9SdrdIuZHkyrbyYKbm7j67NvhCX0v9U76Usr
4Z1nKOuOWQDNWb6lj2//NfNUMTOK84eOz8JbXHfNMklE5G6gykpS9QJC62Znkvz6jB9SFJj0r6mY
cVqMI3Tej9lS7E5VRiJed8Oahnmwt4Ms5XKVMdcqIIf5I5PksIGUoVJVid3aVz5G7a031gnYNbCD
QIvxmlux7DOufKX4M5uI87A7VxIhLS/qaxYDTpxCpMzhbG7JclO+SDhwv6Cg0181I1KlgRPPK2/e
Hex2wG00DhCGuP8RSdw/gB8XzfCTSJQHhtO2Y8iH3HoEnqJTgOxuSdIws18jZbxPuKo6Eu5xaTQ9
lxMCiKShIuxK3xDV38vjxJiW+PlziIIKLWnAZsMqxd75CD09CVYL8Yys4KT2D8jKOtB3EUXlG7Rs
BdFLKKn9xG0M4zJfT5QbEeZwfQzKnBdyVs5c0UlagUBTOp6CMG6riwczj5TNE/57d0BRh1gX+rJV
pgV85IZjhc7YeSySQfovYLFGbNRd8wCXDOgutSRKpwQegoBE43XZjX4tjVaNYQIY4i7YYk+Byqgy
gI9LMUNkQ2YM9WrMw2daNsh82bHaOX1aCNLPBUzA8r9HYgKEEIJb+RFJ2glwde8ly41ZYQN1MXk3
eaRy84USEmBgnZfw7/dRqOlQe2fgSxbJiYWwlrPfQF3iaCZr+LZTP4a0e4v9pOnWAZjX05tZLvDw
58ogWX6zE1i/eUj0lGm7LvxfJAAOZ0zjL8Rjo3fIkLs/KScVqAktrtMjuJUO8ZDAyunKZFvVmWE+
EP2WkD47WFdTx/0BA1LV467xUQKBOknXQ5L/FmoxyTpYLbXuIUc37tHefEWI4/J3hj1iLpzd/Zfe
ENahm4oW5KhCoEtRLEhZEXF6tD+e3PHtohh1DHpHYn9KWgRYNTEAoOy/7Qx5wkxchvBALKfvJaSY
GW9vD8buyJwRh4YRycJI5Pi56/NBrA396bADbk8vJD5yBuLZ6udp7EORUeaxfsMUjrOhthqMj5i1
ClR05bW8sQcbSkwV/MrHPD0L3wUrWBqb0V/DGEiI8dW+KokKfDMDdDDhpwtwSGsHkQgriywBOby+
9CkwwiaWHQ0GjtgpbHReZ5Y/KGwwZH/1XXFxqio2ys/kn+0UKC8v5xxAlOZq7oueRSpIcyrJXwTM
Xd7GgAzQCu9M4x0r8zc5Of2UmcOBvpi9oOMigixvuSDDcimSmPGjReYWcEIuFmZfJK9oTi/dqzDL
oKgfB3iPnnYx9K53DAaGUQ/kce27Z2aeXf7iA6t5tTThuM3lga8GD2TxtdPKk+1rG/kBS2iiXOXt
PgDNVxwA/bdyuAqWD/naN6U0tTtXcl0qIQm3TwVLBLGq1bdhktQaSQqeBhxl1euE2MfZDvnyiSDY
Nidi60E+h+KPGQkD4/Va2ZPbdeV9DamTAt83lXXBnYEVoQFJEMh+3PIxLbl6fwcQFKsZC3F0pOip
5JISn51p5rMI1DVt0qO5nZDFRuyrhVir1uMpLx9jJcGmdhsrQFOWXmpY8sBNolBz4yY+NooR3Y20
Mp853BBKd1OCx+ofwMEZHQiAnm1Ufaq5migeZkHKQsv8nM8NmdDA/ckSyXqZUaF4uNkd7pS0+dyz
007/2JMCtPQZjSkOric2Y9i9t+8kWpCJ3okp3U1+vwogh4GN1rHJ81QZFdwaoqBSZrQvcYiVFtVe
ZH4tVXN8av2EFj4z3KfNv8hKGT1qm5c0NlrdA/Z6vTMordQ/bIxWOEClYpGmiv1C4bW/TNZfb2pU
xmygdMMoA4eEg5qXMmDqusZY+9hFLYEnriEqv1zTcFpC2d7Kq+LcvspV4kxj7VVAPHDVO2KIy9Q9
3+MqIxTIeoeA0Hbfsihvl4ntn0VAS+s6aST5C5SdZOeUg2/OJgrQm60nKoPO9vwpDDlzdgAUJQbw
d9l0eMqkMKIXV/9ZUaZuqNMr7YXyed6tK2fwihYrTesBiKKzcE6i3DkmiPdUOVafZwenjORqv8nH
K1wfv7aQShdVrpjvNsY0nL2h6JGJHro5ahceBpPL37zOK6tOYfHm6fqa5pkLsh7KMsr8yzuk+uoc
7IIpyTCiEiZfbSGQ42xDeL3vMEDuD0QNV01eBsYSomh0Fx0CA1tuMzWbe1iGaO6BtD1tP62x8m6C
/Rg2LpdSyale5gvVfmmyNeCljRHcTC+Y221OwiOQWTa7ZW7+7rFdSXeODWBst7xcOIGz2imY1eUv
yS7i6zNAdbpnUKdNZH472qLyKAGnK3NOB+CggQ1Eoj6EbDthrpgRVkHqHd6/43rUBRewn1Kw+LCp
1eiMzfOC/OClwIF1IG78AJjBObXjmgjzTFMx3/AkFJVSdb4B7cTfp9tXerRM8JnNxFUuVoqJrou/
FZuiDzdPcfDHhhs+oDJiuO8k57U6rTfruLd8pDvDWzMC0xOKDoQPV7vJmB9GVs0EKslqyty7ay7V
1SEd7k1j7vac1hgaRg/OXzjjk/HlJdEqjae6YT2sqijHxU1MRVODcZEif2D5UG9hGui/yw8X/r4l
j634z/P16OLXBKOkf5SVwt0ccNOAHDjsjJBmEhPHVuc+LFsMeJIJBYvmIARV9Tpr/utdGwiBhxVw
XpyeJ3tekvff56VqMfiqZDCs5H82XXrImaubCDr4a4z0/HsPsn/z3Gca6yeUD61yGoYc+k29bsAI
q5NaeLiVKCYAN+3BgLVLUuO+5B6wMzCtHC/mMRc0hgP8W59MORJ1XMYPyhM128mLR8qhacKaapNB
8+BzEYHs4yUKRHYFU8DoMJrLhmD4eHcg+rrsivT5w0aeGGqRG4VWDz/AB8fFFa2nJ+A5g+DEahau
53PYZUvk97wRlHQTek3ZiAqgw3r7JvT0Ul6s3CBQ4zIqBZfto7/GQQtPhAj11bUI5yzdueG+9aBF
LM0Ma4QnDXlMtfVkTlJrZpf6qPdvJ+8Mu14ruo/+tdGgwdzgSSvlIrXZSqccGraCS7TgG8ckH9lH
WRoTPwVQ+V1TVtHGf45irwPwAFosQOQeKBtW30mCrtgJQXUkTVc9AAIS5+L7+a8IZ8rkusI8Vrdl
EynPC+6FqWkbB/742B5CkzlZNZnCC+rrIdMpIfxv9LAZHuei49HFynGreZ8VIK8AdOA63x7TX5Nl
TAQaJyhIJZK+JkB2OKz8QIZVZfA9/qiqdOgh4c4u4Xyb78mJQ1SoHhHRkN/C5m9UyszFoWzVUNnD
t+2TqtonyKQXmIHLh9sHHNU3eHqF+rxNOHWC94N4o8zEifbXkJiyU8AxWYsHKpHn6y+vx9fn91lq
ynCof/IemYUsDav5RCEaqcRUG4XEV4t5k6/T13TQaST/IZa8M3rmEGn5VCymnIFeqMPMaghGS5MZ
PtBWBkcPv/hpm6qW0qtQLMoYENZiQE3O41Rdcjy/2JbqAnLlUqbfmHhpyw3jzxpbJf8BAqdLIMea
YWsyFINc7SeIqiQJTS9Qiy4aGr6qleCLkIaUIRl6y+f+Crnu/BXkZ+njcvsavwcWCE/tXBFevTL9
cE4D2aMyOJoyfrMqNYix/Eec6AOEwKG9UnJ3i8Mol9/0i+gydAvwubMoQzZW3kmmafr5OZyJvgrD
aEwcFFqwqXbNLJMh3TlbqvPeIEWe1ad6n8YMQyidJTLR7QGPMUBksRMUlPwnxvUtSOI7caXJ9xeJ
vW3DVdYuTgLLPfBV7odL9YO3jjSfw2nAHAlL9MtZU4jmLG+wEkPSxowcqjf2ellI7fJ7gBxjpZZa
AshZBd+5XnnVovA7BcWn2qWhvpqaCaUlkOxQeBXPk0Vv86QzGwizRI3AZ5MLIF+uptS3LcI3BcQF
kyPZQiz/xmMxkJd7eszCI5wcMGFHjAp+mU2/tN8U2VBQavZvkwonaaIGXcarx5sYBzwkURjLmbqs
Snn5MLaUmKZiAah4d+S4NuVtGiy73avyFWRduLOc/RtwX84dcnnZrb+l0lh4VDD+FdlNjXjWh+o8
Qx6qAd3zAbmHdzjS1oGTi/FsGaqTxyu4437/1MdY6epzH4HlOlA10ePwKGeVlptRM3JsY6/hw8ex
NygGaqUSLJQks93ccIkJjcvc9eLCo5x9unKBqBq4vvvlspA18ebToXF8GrpvJGm/ZBfmNTupANtB
M2z9QfWc9DN7CRR7l9MzMDVlpjRBaNIeVj7Z16P5MBFs6bDpUb7I5yWNpjjme+bF1OquE1B2UHc0
TanvlRNBqbZW5Zq2fxTO9Nj0L3n422T6Kq2n1DEY5HEwrub7bPMkt4QcaflJqbNyyom7B3JcXYFw
BodhVFK+YtkNzolCAbvgCJwhKZPSubcLlSojVacQczv5P5JZvw4tO6XhI7dKdzoAPQQL05LdCNed
7qwCnMwkHfzOOIhCqghPXlLH45UtZGv10y90SFb3WRF60I7e55pfXnu4Dj224eCOYFwC3ITId+wU
2Sgzjf5S8wInYEMVbIyBKJCmtlWoyiXBR7Q0xDcSIEAwVVcssT3E+pkko/8hPrw49R7+quM6038Q
zUKJZf8BGpJ82XeVpK28QK1fUyHoNThJCrDSNDscM3a1umaFxReK0uCLffmcce2s0xOxOwzXURxi
yjEvhJcV754SznqzjpO/XtsjD9BrbOvGQ2j8wM2pBPLkXyWbiGCCc+2EC4FbB5Nou8CZmYIuUvvX
uG4JJCRYKax0ja4fqhNAQhTMuvIyM9peH3XsUxlojFbwtc+ECE7mwIggvbW3yxQeaZFdxeXj77XK
J4IVPY3xsQ/wFMId69wgwdpsjfYr3IyZZbCWN/f+neaJ3pREK+O6oA3QA5U12LBN1iTh9UggG8CM
yAPb36m+fAYwYZsYfRkSoQgwMYKXLcZWqYgyWKIRyiLzKMqxE9FObqnV3tCTlkYOEHnfg6Gyrrxm
jjrDLvdmgqKavb9JlX/b9lXEgzbsk25tcrUmVXdIH290Dzbkv/mdVczV0Fltn6fKGfHov0lucdS7
hv6BMn/x4mb8FKMzQtejvHdQbd9WsNn22Jzp87FRy/C7K06yXOK1FeSussA5wpAmh46zOTySncip
DSjxHQSDStS4d9iguyxSlacU6lDBWK1ZyFdrCKmqRM01tSIVCBjqlYnGnfOLK48hBm9iaWfmne/v
LR8PlqzFWvVgOMuO20CJJsiMncp+HrK4RJziWYSHwqAP4+q6sSm1cwoJfeqLhwcy4sJ8REWuVdVL
6aiz+JngylKW1SceD2Aup4CTY0J/9N/7WG58dwfyXjyeNZEEYyU+VOjYnZh0AWEx4itnWh3vYgxu
VGAzl9iOjaLBYdv8LBefJqC186hpsr2G2bQaPVAqsBGo41RyUm7gIcAdcI9e505tivp6/a3Xlq65
AX5jc+wGyHUPlmpPykyUfSTsBu5o2gx5HdeqtvMUbmId414Rg9IdSxGDZ2F7xpdf4GJfCh4CbsAO
0E532/6HTtbhNmv+GabQzxZdSUwAWwhwQiwBj4grewuDwzyPaveLlYsnDbRGUHBTALPiK7UwGEJF
/KNb7iHGR+CS5vxDSlslwkf12uyesTnx2rYDOW1+Iqz01uqXkn+BsPW4va+CVM3orTy0dP5ktDk9
pWTJglslM/MFI3UdUNWrWDi1/3Fh9TbMPgyMyJ9WKXCj9T44GZ2Cxz79ezGSl7vCIPLgdEIwyaxo
7LLznjzsW+3P7004J3qexJpIbxfR1w4cNFKrigjCwnJa+W3zTsKixzKH6fVbOdY2W2Fxls7Kseyw
8nDTT8Z67apwDGZHXjIW9iymMhiv6Fpj14f+z5fmUG5QKDkU4tnFziYpWQUV2BZ7TGx4FT42fi/t
IrJ+0ifzpYeScVEWDrYqyGyLn85tdb6cegaGkqBvuPFeri33tD3cUnRdKx0+bpnGrTKl1kYXJVHC
OcpqzDdEeD7Es3EU9CIYn97FSnvukyt5BwZB2rJlczJeXs48oXWAAqYXDvRnf8uEFpDGSguZqkHV
/8w7uEg/a3JbZSRUO0Q3t4q3PHYInjEYE1pzWUcZPf2j0DdIhfcxtKDr0dnhUNPQDC0i0ORBeSQP
tgUxmnyBBt1tGnM1eYxy0WIe6LyGxhroSxUfnKvIzvXKOWyKsGHWTbr1smvndzKllI4QNIAiu1ML
cMW+4Qr3ck8RRdHj+7LuoXzQxRLRmeT0HywV/kzx/5vlS+n+wusOis9NQrmAWkhvaledHN7KqTDL
YbLMqQKzu7wgNgo1Yy3d1VXHdprS1lfim+u/FlncGfNa68QhJjomrzSLet0AC2F0M3ZVrAzx7G0G
ctY8skx3FZMoF9IPXJc62dmGEIP554/Uu6JGfuFtyCRxtXg/NmTsaBG0TZtCLx5wA42qy4hd680c
Xf3qO/pBc98Ga0Mtkyg8umCcngZfxBXL67AtdD/Y99PT3jm5BG3rKy92OVBLKh3Wij43wifBAdvz
o4CYDsVCSnj0bgbLB6+C6xA18UYj5LH4HBj7piwFPXelKxyl+k4RZBivewrSWixcx2LqVrGqEyO+
T6c82sXpKdtdvkURwkNz/GYLeW6e6y5XD5u6B8CB4iCckOdq7e3aV+uIGZac0nFCmpeJ1H3njcnN
WKjsad5TbdSxVWYhVE3kSLXv3Br6YJC5bHZKqU7gMDJ07krEqPvuk/5XrTC3y78zgpPl6k1BgIoe
jzdwKBLyLqnGmF/b8fbj5D1tuLT70pJyo/r11zE5vfcLRxQfoGBss+BS86Lqmm2GaIYaVA2zHS4x
tiTEBX4Ko4nE8nr3DnfC84DKjwPFu5u6wqw+PCXxD1kfRoSN189ICTG5rhqYwiBpzmLO358c9pDN
CLNAlhVFbdLLLEBoYBWOHr/1hS1qlSWHBaPWG7oOFQ6Xa3tmhiUWd1O6tqQ771Hsaq86tUfcsAco
dfijfbPBao/kzGDlBRHOfk5rk45u9xPaIacgZG0F/l0nM6j2aGVPNAePLQYcnIMu5ezezhYDDOLU
HY+BWm/yTGq+myMw2dqkOiQuUecgDdl96pvbq4eDvIIkqJDhXEKcrLiXvHiolYUC/GuAJb7eU/8b
6vGNnimOcQSEPsX0cKnQEdmWOCljIS0r1UbIvH8F3UOIVX6tgDYg8KGlFZGkJhWC3VCLEQhX/rkr
Z/gDkJBkjQMoohGBQC2rqRerRZzuT7FDjCZ64CJSeiFqbYANHt3lOR10XGLim2o/LFUv04fazmN7
d0SMCX4Ftq1nCoCV7BN/BYM5eUxK06acPPgtHHtK+g/vDjkkPX9VUKdpztTMQl8myoSZcnnYuJl5
TFbMpUkPxmFUvSr/NoAhVNfAPMF0uuCJfgrcjVibkC7vCOA8eYtDyXTpFYkcR0kfL27tBnKKkbpN
lf6250FWYNgWgE/A2aeCfpaAV0g5Zbj2IqalKl102LuygHKLhWNM9YVtkZH8UJ+7xC/0lWPFde/7
ICLAk16QLU3wBV8GVkh8TkriM97+cUwKfBp//bWlvYMW5mEkdeDUU8qo1phVrju3L1H0nNi55P8E
Pu4F4M+4vROHjf317bP/6Hul5rh1fgbtFcrllVzl3gilKZ1fsflhewODOaHcukzes0jnTPrBb9i3
LiQCuyZFFILlpeWiUDKmfeea/qNy4mNlqMqwNBicCsj6cwoa/xTIJlOYSj6DjzFIrtK76HecrRJy
Rg3+C8xRHp0+cYhFElS8qs5XPCXJ3/oYoTZ+teqqNgsVww3e3/PYJPjo4JXnoXovoXDVaCudE8vs
j8vqgmJTpunpDTvyt4AHQRS8VMNPllJufgbV8ReVFQJxZn4c5vcGIbzg/6FNaeSULDHtJPUUT7Ps
nUuOwV3FD7U4mbqs5eBsTBipamc9qYu2o8+X0m6YtSOpsQXjW9+v+nMdOUvaOZCJzbI+FUDzuKv/
FfeGjEt7RNzD1EvvF0e3yHosozQhOlfU0UB23UsbuMx0V5Al1nLdCn2G42SBBM0bXnK68IOVJ3yB
1uvBTCNfANERgeaA1E3CgTIF+RiEhsM9cNbFKlTV+BmaEwpQmMaF0QBYlEQyPXBEdu0rDkZD88UM
TruOmtb1Qdif/wrObaHsM3PPh2En9bEbcRQDbKAc6V9IITVfaI7vegxUKEdgIv92nOcgZHunADb1
tbSzYesmcgBqS+xpd5k0lg1Pjerw88X8MMtPt96BEfYOJz6zyEtL1pK9rAo78kKLcGKMJ5fYbwoZ
bYjypqlDBiio5GbbxmQCAXD1krLK7pLy8SIWMLTJOSGqie1Rb14jNNR4kxj47IyXNPqMyfVuXnQy
CbEfV50/ocWQkJuAJ5v/F2vbfXwF0UjtMjXXvvc1453y3ccJCM6OQhe8+RIqJGPZFxAYVYZVZ5I7
VzDFj1YSjGgwAuuyQO/V7pE20EgpYGGjWuJMSx3Fm3016KQSmaNkAyGhoXGt7F5zSCJwJbQV9XaJ
gQyCrgcUN8iGf3kTQB4ywYJuQqJRxRKHQaY3wqQpb29dZVvhWkr9CbOqbe5bF+Kl+OKFxpJgfIXf
wNGdp9NfYoQUu38Heas2fY3Y4+72jMdI13z4bGImHEhen3ueCjSGXdRnSBgop+LdLrVP2q3cus/o
b/fBQmU6Ef2h9BdAzsUAG3qe/psLgpFSoaeB3kWPg6feumiv3ZNcAAVpmgvCdnvg55ZOxjd7qhkJ
HvtINwms/5veD3cMWkLU80SddnW+irwWXVUkt9UVabPJzjTWdZhk0qcPzmQx48VPBjL8ZhzWAXcI
PchV87xO3CZllhGcYsY363h2AHrkdwsrI2Up4dWUJLgnZpJ1qZkJjy/4ie0i5zXIYweInYUuzDq8
CFI2nMxU+9VRDV4vB5c621rVMIRbBKKUCnxY2Y6Ng6Ioc4w2mbMZsrE89DPtRTywub19Rs4QbsfA
64G9Lwu5fuFf3D0TkVIopUIYHu46p6CKRghW3kVOUqu9rx7xc+VQgXT6un8iruUs1S3wMAqein/d
cc29Swk4BCnYdLK7lp9YA0zIDRjbvkMki1TCKnNhKFBNvQLKRp/2jVuNgH3ViubXrySYlgdXK56r
l5OsPVupoRxbkcL2XvsWP9qRwWKM9/z4+OrpFzvYC5Ra0r/oIDXMQzFu9DQER+at69GAcrB9mhi0
IF1w18r0eVQK6BRvXnSpfh2MJLC/71kC+wFaTMQC3y0ssjU0nbrUhYDRlUbydwF4CcwvWUD7zGtc
MCYkjZQUYlmyv9VXbxKQvdGiar0U666+xxQaGtn6yAZ6FpKUgysm6HAEJqYandgaSm3+vpO2AOj1
Ge565imYfxrnDLu3HoAi+XlF0ak+UjM0c+udbeNuTxsoVo4KnNwCN07LBTqdQPqT0eFDOQVuv8SF
vxq9dJkSqzGkwz6qjWUV9Qpv5UhXTLx60xolqGMx0QtPsobLctKeWEcJ0KoqZKnfP5O9CbCpuLxD
ACOCxcuUgP+Fmm6qpdfWO1mFf0iFHjxdRb2c9i1TfPt3fA1BvgiRB1c6lHpiI8VV2Vknde0pS549
m1HIOajQIz7P3AfMbbJR2F0Bou1asXS8R3keqRY8wWAY3tL+AkRExkb3vKYw47q9K3tNQZ2XH1iw
yNbeY99ErBLuNTnCAkZITwCUT86KmO+JcCzw9Bpc0PZqanVaRbbRexvTbPXwrKHAoYmfj4TsLdrN
5tWTn9sT9wj7c4AdtXrQmvvWZjapHHhe0JpRz+BlGQs6nnDWSpHuP2UfKYBeCebCskxvSCWN3ZL1
5LnihGUZM3S9xihknSKYMgnscpy5zVSodakBDWxO2MYE2WQRklCpGB2RARv2BWjusDNqA1olp7DY
soUTkEBpKWaEe354ympu6yUXK0Z9zDZ/NHQ671QqoHcgnprRSfi5bBZqog6qz4qJIBYVjQNScw2S
r5GgTQe9F/cpw2xO6ST3o7VwYIJArHqnBHxSLHWf/TJlBu+/ItOfGENcUdtxBIKopWxUaCBth5yY
p3zqdm348ojhazrBVoNJ9SS8pZaZ8UT15lKT8UyWl+SjhWDC1v5q0uFFyK0wX3zEtZ3fkROra3FP
rk7MOSNu4kiSyTQkdkO02/VUzaf/S/W0vjWFpjsWGr750QWiscMfg4aaOc5e7Eb0naDK6W1sxLzf
8KzK2m6UZTO0etga/WNSQ2sUI6UIYXlKOsbiMYRsIJo5gFEnXZEhXLEo/P0EkeAuDvN+DEqEyzOc
TcbTSVCxiOY+yp6VCn6D4QtfKQ1bV2CvHSbhItcX3i4FKhexZglO4JjjJZ3oa/Kxu6WerDs69HSx
vjwmYg5l0qWwpJ+g053VHTk4dASCoZSf/OFUPEtXzVSVaLh9qkomeFmSvCaIj1EANQaEhfzQIoDn
FZh9vJAlYQ2JY7/3QRpjYqMw0kAC3Oozcf2FEBQbme7VboMwGSOdEzT4/0V6VqcYe/ywtODm8k5m
3jIWM5h3xUdFtG2fd4EX/hs4vN9VsUXlFxni4nBJWchQFONUxl8H90kstqmwTRTEZkR2BVvjk374
Sj4e/tLHZS6A8gIa8BMHj5QzdAfYvaUcHNWmNRsTWGcsNPwcS17fXsazMeJQ6if/4lz1V76Wpp+L
ZaJ6vY+bHXfMf5YbrAARJ4ZrVuDjqFTZuwG5q0HDA2HYCs4TApvLSJRexxCLE+wVuJ0vXMMvAaGK
re8oeV9B8IVxMKOrB0EcrYcGmZnMzj/aRREOkSc4Zds2H52cYwlnMm5UsU9JVaOGhMZF8s5B2GoU
eBWgZHWZGe8sjpVMbmwoyWfwGfsSFbnUdISyyYXIJZm3sNQ1ytpFvKgAf/z6B+NY3EqiEUYp5+y/
yKjuH/mqg3aWG8YjG13DOSDCZUpZtNh48xo0EvDOab/xFPjn2+WRNnlFkcwEUDQCiXHg4mtY4j3E
Awqyl9Txy8/jKpQNZP3PAKA94ZocUaCQ1tjYhIF4UvwAEk+Rea0Cva9FfigILclnIFrGn603iiMa
VfxtXdPUclDqoDXrn0U0STTtmrFEwW7luBpHkTBooMqiOr5XhrDq3t+2dlUYhMYWeLa9EOLQOIL0
o9zWmC+qFAQmraUnuVlWVSYNuLOsWQLei/I+vJH3HZr1OZs3A314iVFPQoHpTPhEciDtxdo8o3uA
2pIZB6oa0P7bnU7h2Huzk1v+3lr72y1hgNvo6K4o/O1jAuBYPjV+CfbWcpAtoDu0XpwUnENRKS7s
SJEf9IW+DqS2RiDhEs6HbLkPF+/lhScKGHTnOKv6bGIcX0O7mG7GYMcJWnMDKQznkKrZe3b0dgBy
JJa7HEY8oVe13dYqolXYn0jtRwlCkJzC3VUMsUAY2XeDvYFJz/p15jw5vtBEWaPR8cvMyA+0mQ5w
kjkgBl0hH8DWvdn0PgsLd2o1HsxTso8jO6qEV/j9BUN0xie45MH6HwUzl9rfgUhL92KSi+BR5a8N
Jj9CmKAVQ2YxnFbceMBnsvvtPIXjwh9IqmPAmdYQQ9cpG2ASYYB30GAbcA4CzPkS7stHRCPZaU08
5QYoRPtS3jSTbGMa5/twWfrVAVI82Av0j7JveILF9X1q/czqQAerUpKBldsK1CrQD/NnGd6QZWJ1
EPn7wZTWGkL2bdi8xAitGxcXc33RY21TQLIw0OU+YSUeFZwUjvuM1tUlHLPOdp1sV3JbsT1b50Zo
ThH5qFXzZkjsSzKtVWlYPhlYR7uhTVB0K75ikIEw0cVft61IIVD9x/uA7U7/Nw78kvPRwrt2D2Cv
sUkoupvdpW53ZYAgCxpnIEOvJ+X8b9n5idyyDwUz/nRjbCm2y0a510bwj4+ExSnixO9QfUK0PLty
ecfOh7pGePhbmHrXqjhTmXbwOmXvlMyFv8LhLdNAm94HvKVpih6i06jWwPZUQOr7PwUkM1xFfwtY
S0BtepxkfPYKBhzbEAfBOA1dHp7w3ihYId3en39eas+brNlAUS+fO8GpgBwLu1CM9nYepZwsQpy8
ftvZ2Ms6pz/IKjNQmgd3/ZZUt17LNrc7o6AaZmSFKc6pMmhST5dj1HQVGkGuUCh902DjUuKA6i17
/3+u04KuuWBIAJbFwABcWTnThd971Pal8dtwz3dF3wiFS1O1M0omiXgoFwN+RfczZUbmLI4yG9Og
qbLVt4mYnxbM2xE1Y8X+EpuENTX/2TDwKbqQv6Ynv7JN3z243fCap+8oLGwLyQ7NN6ojF67vbkOH
73NrVBYl9jfuwed5agK9ErB0Kit3FSF8wel+YiVKiyN0VbCt+akW4XY5WnV9dwJcOEP1K55+Vh26
7SoRbvzBliDaPlun+6XLjCQHV+NgLdtPfcLkMJkV/bCDXzQ1NtI1MHyJBUmRPxsLmlUewSOwzXyL
EoV/yniv7Q6z/P6XJE5XzwxQqhM/7uBJgkqG3PbTbUMct70ULhC++3pIWlnaXzccHQwiAHtHa6li
z3AKrZp+w8uloH/uGfQXuFk3cshQrA/tOBbqRfzmQbMWq461VYu4o47IjjGFiwQvA49ZN7WvF2I5
1cjQ44i2t7uWLHYhNJ2JsFuYnqRhrBF3qP+oCEsz2swaSP9N4mzuBIM+26xxUyOJQbg3JlQ2vkEU
Aj9SBi1l1h2aEf/E0S8e5BNxO4UrP9nhpdsZzgRkd+ZFFRTJiRt1W/wI0YyCia5wS8RngSW3k4y8
faHGfFkHnqKTTVp3Oy9IJJo/1HZ+UpQKFuSCq15IZOKDvTiYMm8276dAVJmPAl4U12JgGJzpwMwo
olNtrFDq9BPjPICkDAPf+M39Xi3dnCKxiPObfhbO8owM725+dgAtlf95wu4J+EYSa0VlP7+XTdDt
kpjo2smMqp5BqY0SqMm6/bqvke7wnKMiQIbWU6uD3ythF3NK8d36yRPR+ijwc0UROWiBMLx/Uw9m
y3INuM9gbR/hF+Fny7Fu4IG/z3eviG66rabGEtYpBWsdO0u9McRxV3j+kNzyLkUwNnUYQP9opcKq
M9ubfQkYRhWfuuUAf6mFhVBYwDJfO3/avXk1itBMXfccTQkuQW5fM0zLA/ZZ9GGhuhHyz/aYPt8M
sDwbIUEEFIzJV+W4/UCpRSM94rzY0+QjN2U66WzXTehTrLRJ2/MdLOIkWEbFZQhTPfS3J5Udo7GO
QUiAdQ/t8nN+oMuhuwRfjlxf6ebWuIOK5jq3M7PxHPfxFLBgzO3fIIcmvifTgsfB28LpOHnrjO9P
z5IiBZlHMmwYH4bSiFuAEt8Avsahb1EZXzArCEbXU+ILtUeN6sfj6ZgpUgYIM3yeCWUV7RYneGQL
UP+kKF9LHx3m/15Nux/S78gfQkVCLwBdyKCZCuc5Mf48kP/T5jtigEbLJwB7cpUQtD5zWAdG9sEe
wZPRvPAIQpeYHCIUicGRooRK24QFGuJiiG/Uauk3ezpafRg1v1RxoBDotxj/sdBjLZdF6QKkcaXZ
fWojLr0ELyAZwnAi2JhMJ6uYPcjQI2GiuB7vgaDXIxnoFbtFbUnCn0fwCUYORAO1M+GVK02jf5+9
9nvcCeQaAMNVS2LuT/Ytqw3vTLjRKf/XYfe5WspspPlgUDAaSsNfEpSfEgXAEZAIVKH3P5UfE6BG
vR1V4nywyT7+3F5+nkgzkTvHtTnKA2Gdm04JGAYbNK3KnGgUZnrWbbcU7IuPaJZUtNIkUjAccUsH
elFe1zYHps0AJ3y1t/eymYexqgo1u8EVXPglgM1JrbgJ8TllM2Cyjh6dXBl3TYnxsISA5Q2BuDrW
ur1oMY2WSR+cjauwe795O5VtkPbdTrOGv2s8JGT2Pvu5TTPMCG2kNjesi6GM2VPpTf05YoRBfInq
Q93dRZz7grui5Hq7csAl2hyltyWtGqu0u8hYdRQaOBnO+DL8CTwjUvNmHSaBDHsn4SuedQpp+T+r
FobE3W5hO3yNh1p6OVV8daB1Tix8qORNwNY3pyfdA7XHgdjGOzJeb6OMlirC+U3jOgNxZVkDzk0x
o0WeXx8O+c1Jwf6EhH9mlaByY/8RRV+xoZi+kN/Cw5K79JnuiYUvZDtbIvDgVvK96o3jCBEuy1/f
0wal1ohjqGTxmx1M5cbeALZ8x9rQ+ZUpLquweHmHZva1xB6LJMbEYdBTf2ziNuk+EeSuMigIPnBl
63gGTmKLmHi2tT0yXHqujyNs2x0xlNzJ9oW/G4jLe3X+kpzdROfkWhcVvx4tXvRubNMu6qNwTTVo
vlVXgFosUB8Gnrj9ZplQTlpRt5P1Cn9sUbLHw/qPiFrye5ww+2+aRkS9JddTfY4YdL+zV3wAiT2X
CGu4N131ZW2SlFE0GQ8Gc1f0ucnILvxEeOyTMAoxRDMWVL96wb4LfGzw6Svx3sx7GE+KtliJG6O0
CEm4kul3+J6OpISgyleRCU9pL1N4uyXNswX59Y7YsrEnCEyyubj7crFvP+1v78q9PjBFtolflEj7
uc5wa4Sota0GtCRHnWbSttKXYyEwahPrmPw3UZs+ZENE/DLMtDqrXtbwuV2kr9iPnjGdtS0B+xe0
p35R8SIxm37gx03+hIL6HGfTTKMV9cvCM8dedzGmgpXnvJlNmdZp9AK/2IVZdCQ++/yDQ39cCn0p
v4zu8TCMYeqgVKH7iIOi7MKO4CdQ4iw0ZUiQJEB+yc7DzSE4ODlfpfRy0a0ISHo3L7boLLP0revE
EdLjd2C210KAjuNBXsI6kiVpMUEOfd/WirPLJYyDX3p8S9NZpRfY/LInpr6sZsZQClQgfOtp0Fcy
CzCuihZQYZcOrQ6hzferja+3U4m8AmaQ/Caii/k8N1fHWBep0bSvpTzYAIRFH+aJ5tozxJXV6bcw
s0x1RlyAyG/cGzpu8mErfD4XIXaV+iv+oJQqhFWciIVB/B2ILAUEfFUlPu4jLWTmJd0UHlizo69z
dPNuXN/yL8XtMIK/v7JPny0tq5XwAo6c7TqZs64zrHpU1oh4B9WlDVB16+OWhvFmZepImZGUa7np
0I9Emu8Y7MpgthnA0Q505qVjXe4aaLCZ1arN0skUpE/Om4ISePD+IAMLJUR9izMWSh5zAuQCtT0e
HqDyhK3GPnehncv0wv9pNd9lgwN5qp0nw/V7cxeBRDpH77807j9LsRzp0+rBApurKFBVZy9edX+s
mgOSPZCDAnWSNoPlfA+0XSkjgWSuGx4ci78ZelH8ORsSEq2LZDBHSkE72QiCFxaV6GoxJcOzzFL+
81qT2ZZ+sKuLXtHPh20Rh71oJpqRyvG27l0oIQhnXqfn4a6WOJCUFQTDpxDqT/U8upQEQUeXOvmk
Pb+UVNXlAh1uFjwixuFSJV25Os64MrCW2rfn4tefmf76dqwsvnyPrYsUK88+mqkTRaaLxgb7yfja
lkG4VojgdtkqBwuc2WgB+f8JLyG6OFJqAd62ZW++iLNsCLxRYnEVItpgiz1VSAiKSaiXWTJnuQgC
YdtYRUSgEE+/GZ5ICFcoz031AzDXEK86zobAQgdbQmi1elluFsEnLqckGe5smy25cmm8ZQG9ZfzX
d6SABfDTor/lGGoM70o6+tAzfZRE0xCzW5kaL4WhyKXWHJ1XCpeW1IdAsUfhWgGChWvBvbo0FZa3
mQOfidVI3cfCj8x8IIhRXC7FOPsRxq61/dHvOJ0rNpVdkLseCKhuQ/et1d+sizSkQcdckY8hJI5S
49VoTQyL7G+B2VXdSMP/4y2icY4e+WhT7k+mTR0JvZaRxGTP+2J47KWyycDbq/3MDlKsMUmXqh1J
PsMW7o8TlrZjl1bNaJqVSn61up3Ew79FcBIGXH0jW1YkaQjZaeDPTw2L+y9pbVSsxS2LgD94afT4
k/JnpKJKgGCybLAsUaiHrUqJjLKTFhhq+p16N4qpHCvIdIt1AyCyUJiTEURB+L3lUAKAV05Ff76i
dIOlYP7odStS9fWcngAvjDreLGIyfhLG9ERKHs/ktFUX9dkjoklOV2t72eCr2j8FsQvenSy+uHsK
M/rtsA7e2K+XFwR0xa39BKt5hpG1dIZA7yy0T7ELfNSj7vjgFeVMAohXTuyhev6OtQbYJHv/aDNK
yBApdl4GVQ9548tRvos06+TxyxazI0mQkQgfBmTzez8dAkHGMU9BZ5DoljcPZ3i7r3gcLBDZrYHV
QJfcjecYlfJQII2Uthjt7pqumuI/IWJgyLS0n+S7aEDGF18225qzDKtfqfAx2DX1Lf6SFT/R6pNg
nwuyWoh/0G7Fj3ew/I9KZH+bnvqaS7hzwX1U7hDBx2rGGNnNe0D0mStiGUREIUaX5iPEOuKSunOY
n/8GTM742veKusNRh7f0JBNXFLNojmY2M4cMcrDfdsSTkMVMo6Y04OTf72as0lqvU6c2bTgn2hw5
GRF4qlOPPgS1PqppAENu54dBL85AupHJq/eFpKoY5VRmt4iIB5sm5yu5BFcQawOMLxJ2KAbRulen
83uZ3YrWC2t52pzK8NvviBpBPeBkwWHPW3wzvinlC3tiZM0ZDJsHtY07CLVoUqIo83e31RAYU72+
dQf+AmKwNBRT8sjF+Ig0hSdbc0qMFeNyfOac3FC1k8AyTfDjUE9c4UtrS1RPaQ657jERMkQiMVOi
I+mRsidJZ5bpaLIAuTUwq00ESX73OmcVgEZVu+YCdSXnSmOaFErJYu4lcRWtV3SYx37kgvS7dL4a
oQ6e6kq4tGOU5YraWl9oj024E7BSCMClYX+TtJggBqj4QfTYg2w9QrLy4dJ8L8P66hmjONzkeZmT
3gVirbR9nGPV7Y1C4d3WbHB1Lk7/NAHr59a8KeI1oXjKMXDciLgJzNIJWSsee1MmCA5Dgf9Epip/
autd6o2wb/R/G3Iw/q5KLMimnKS01LhLMy6dVTjtnvf48a+cGOnUQoODiod6fs9TYhY8sF7/k2qr
+TIJ6nukv+kmtlMnZAAuEfEA2/xLHQoCB5CHyu/FdXBoXMELtJ4FQoGjema86PM1hCGPsyLB+1hc
MgdselQ6cvKt/0BcQ8uawH4kqEyQ2y5+KYUSCaRCnqxd6M3Z1qRdHZUQsJY7mezpU1lRx/Db/vbm
Fxk1KgpCpg/xQAuEYW6GesLppFL3uSmX9a0f5crAEQWjHpimFtoiO+bd8KgUvV89tV7OK1cCP2N7
ys0SuuRLlY73rbQ1HnPWhiH1Yh4tHqXdumX/xd6eqWv05mi4cFrAInkCuqOuVgqOMi1kcp2SWI4Z
bo1IfQvwAIAGqSxGdT+hhOtJ7UkwAYgKk9H6ReCW73TbnXA21vrSXrGjAMuyp7oMStTU8evt8/yk
SSFgHH9I2fKtT5dtP/HBEDunnB2R0lO0+a8rBsfMsFvZFQbNw2c3QR1D5OxJZygRnvpwHW3r50+r
8TGhRszikq0OdGnKwH1YTfS2WV5oviS9/XL0lyFHCve7gAH8qJAeToyQRmKW2wMu219LaqvGovI/
cwPrmDzx022bWJxUsKY80ekQgX/3Z3lRQ6l4NnNlVc/xlr9eAM5CULQcDFNLkuYxf52B2ExkgP0u
bAdgEfGLFtap4GeMMN59rMB8ljBIhZu/Xh8a2huYAvmuPEjC10x8ssEEBx7VieJ9Kg1IKxfD7pPE
bRFqQclVGmeVOqtduOGMTUfsgyXP70fjucNPty5W/LZRXNjR2vyCDhE10XPLwnULkcUfwrDfV52U
ItEJ//VuI1mm1j0sEGUZ991ubyZ0SwikaSRMj2fffhKgsplvGS4Jslpkqz+7cqAqH6iBVRorQvQ6
/ns207E0bpV5gp0FckVWhhbFhsihreCCdgwZRZilkXSxO81rwVZy87+jmdbehvhtiBun+hqZALf8
ubfT2NoefaEIlq66VCJThm2DvGCp1USR5L+4IZ4i7rBFrMFA82HfBtFw/POYkVdroH50CxScPhd5
Fco0wMv4beJ2xA5U0iiLCvoi36feZOozOUWzKMfxTrP6s+bkR/B4zZJ7sHs+xhNLODO7UZ13Xytu
eiFhOVSwR5Ry7B+LFYrm4yTNVxyKftI7uCPiIzCTLV1WWNPOEpBAaDZWEmPPJJAvD9CL0L1kPhYC
tS0fhUF4r2r1+z6KrRO8U1/tzr4jHVutYs+fRsW9+D66Bo/nP/c8emMO1WfZRd3X6NZ5Ew9QnOP/
UwZ2DJHMpC/u2eRqc9yZqfLaKnnZJ2z8PQFWm2dgI/tMsfe81aEKQUVg1u/NG2ZCxr0MKGz5/l4a
4cWWHTH7j+F2hB3+3pxZ57hLsrfM3eXrp+hIO+BT14apl6/eMmKCvPO27jdtLJOZvT5ObnKsNWGo
irlnOzBL6b4bwOYa4Z2g1JRg3KKqqp5n1bu/NGbdMPXcsHwupwx0xZxjlWCjr/98LkLiYikVq7PO
jIt/lpvpTAOTXEFAJ6ZIOu/YUGou4UcjjOYWpVXnmy54wwTXad21yopwIixuIwVtgz8eXW6VlH6J
T5A7sWxzG6VUUxMZa2YNUS1AjbsMOc6zLPORRBFtuOPp52XVIsO3xo41+u1ZFYZHMUg7ecDWlCCC
he6zXEB+PVgM9lrh/s8TZl9tvvVA6LRt0IkTrxTuNM/HcydWuXWYGRUQ0//KG/d+b1c5aTsXYxIm
HSMtKDHaC5+Wrvy09IYdWs9JiRVQixU9SwggatPFlVQIXwKljHx4dNOhqkxGyPjs3xdMD4l5Ynh5
xnlqoYgOh+vDOE73zz9AT3pvZ/rGRtBtBOrS7bTaCidg7pel6ypGXXgX2Nu07Ft/0+ppaAQ1WTxG
c5EInAsBs7x++3Vx8OHBETvNHvmZ/QIYDgvh7gLYmetA8oLrVQ8zusSWS0HXRGN2xJt7CYJYOuqS
tunjOj9rNgulSUjOQpexp+LzV/O7qeMMVzi2lW1yiOhJ+Jeqzp3vbzlbKEQ2I/9dVPBGic52LkEw
BKLTB1Bu05QGDzO4YQBxn0/Wn1upUD+VqQyXOdZv3Sma5sN597j7CncfVwOjNywfE8LL8LAvJxw3
CY7XkI+lEZocvYu8ksMU1ynhl5uj/Km3BtPOS5QWnHEr79NiWriCJB2UcM8z8Q1dEoCi83+h60Te
zlI31DKPmGH5qOLOJkSY6Ir97hkO4wmlu8KwToWuC6rgThDnxr5e2rn8uOw2LRn7GOHaui/vYs6v
r8+eEBQuEeSDVNPbnneMgYe2LhgpTwiTqAoLGowiaNWqwUQyLVrZyQu6B06WSTp7N7uFdQWCDfZn
Hii5L9BbREpfDZy5GUTrIgC95wJ0m+QDLQYfI1TcaLf5+rupvlNd7H01DVILb0Q1xvzVEo/1WvEz
r7Sxs2lCLhPmj2UEvCVvm8BGi3suU+KZfenwJu9lnIOHpD1f94uiUY+BWtBarAZkMhx4fpKIvjSW
ngxBiGkwvmAwgK/EfR2NOOBQvucqg9JqWLCr7abEZ9YMpgrkKslE8G+3ECb31sbYNhNihWxWJekr
irdWNPNtshANTU167RnuXkuLqh9CueogiVqdY1y6ysTBDSFkUvsekNqNAsf71HY4snYQOJYuUrSN
poWfiY4OlFfhLZ8w39A5XtDwKPf1fo9jKiJc4fXXHZkXqhUb68Iwr6lPXYKzfP4RwBdWe6DNHm8x
LWFpNqX9lz2BJx+7acLWIkykIBG3AnvJUYX+PcQMBLBuZqiq7WIjAJgS4EJ0EEjhvv/lk/hSIQoF
YJnUJp9ttgGRFYV9+7ZkkOFC6yJg8d0KEIAHultY2hbDq4RpR528LC17omYvf8tZ29g3d3fNNDxr
j2mejJE+u+hI1GE1SO7GskziLZqITbTjwQ9ZTW/F5kckhwe2Qrz60a4tt8v5Jc3329kESIHZBliE
BPYKukY0ux06JXrr+r2JQSmXG8tvY4btvr1uMY0wldK5EURLxwEhAzElTo+vLhlV7XhiXECsB53K
t0IM0/VX6QDOEeJwVhhRVz9Co8T9xKrWiXphfY39uVe0kf6CEiTQxpqsX9QQ3sWja9+sEu+Tttj7
iSg8CCGOWo7zzrin43FaavgCQ2ydALA1DmznObYOzzdA6SS48TX0O+Pw3Y3qGyOppa+EJR03KYVq
0qBmRcGh8zS+nd9qYLtHzSgRJFhFHVErHoNQqCzJ5XvRrMUDUxVGh/GYWXKUQIajAhUKjrVvn0ZO
o0gN2QlfAfl9Yd3oq3GpcWxVbWwsTt7hSJk0G8vf8epqYc6QQkCYhbCZGQ/idEXCu4Jniic6KM+P
NNTogA9Bm7cMFVdVSIRXoUf4+85ZGJJqKTh7NRfMVhlYGe1uQ3Et0Z1GPsvXA2ehwUaKk5RQuq6k
nQ07j5FzjjGva7KThDoCvQVvJy9CKeXWxNnL5ZDj9K4X0ZQdQvbw77e+q7RTZrmqB87sXMY5MW2F
ni4GHGMUvVnCwtWFFwA6AHvCjW1LgPVIVBE6eBH2K6u592WTSVbVNJtEQE3gVg0Fhmv3dJfWsk0P
pdSOi3LiHD2M7+wbR2jV9+zlwCz/bJWopa3You8ZhEeCHw+QgBrfGeGSZKKeIqltW82y06+bYAa+
3RslVDjBniBqQTcjjEjZ9Ctap91ROkZnKNH2r6mduYQYA/mxhPlIotsAE88kY9fA2xrxcW2tMu6d
lUPmf/ka7HqY4lliyZG5L1geaSPJ14UaEr8lHCMjCSG+dvO/RoHVzPK7InK5sEwVFiN8lkUqqnmN
vibECS/a6Q/MkRJWu/VEndumCXkOfhd5jGU9EUaQe+QGEHDei1mSm5aqEyjaXofcCgWam6XSPQ1/
3s3FPqEH6rNDBC4Hj0hvb4zXwv5G0DkJHZEiYGXwfcD/Xl7pooF3TkxNEpVq2yrotE/YTWBmdxbC
Cni0FiV+Z9AcoN2lgW85FneuuYHiFwBers4L14bPG881AfHg7Ci1FQReX24/LCk22hVXVGg7Tmvj
ibVSI/na11c3dViu7cDDwQ9gfk+WTw9dBEKa4xH0b9Ga0bgkt+KULyh/SZdncLiMD4N5vVGY0V4J
7yGKy6jzlNpl+oxiGiYlsF45htEOBAyLF0rKClSxP13r2OLwUFETVWl0P5yU+jXqZZ21EOL0wEyA
G5QclYePdBHlBhx9368W8HQ404a6fNHUtSag6FD4PKrMnfLWoEeajusoOvIT2Jv4EUBCMs5ul0tM
PUZ4FKSEQU1evB/tmNo4s72KBzzakBnB6GbtwSF3viIO4Zgj+75ey3mBmnNZaDfn5gimtSkze1nk
a/vVt3yBOx7hyuKf6uWbR3rm36jxsaqH+2EhbBnzroCHw5EW06ysAu012bCk12W+xEW4h8DsE6uc
kvS2zc48TwtmoI6AZq6aw1Sp4Yjqr96nR5eBJxs00OS4C8FjHVb+GrxdVb25UZLuoEGsYHdjQpji
TJW5NdUJeWAe4B8WVaAf3M3ARzHZJWn3tTCZc4WvgjFphsNZBKFcT81MnCYeJZsR9Z2BsbLrzQDt
pRdavB8mOz6tpNIhzIDQt+U2npZMw3cotauI+P7JhuiRiZhq4ERoelKwxbco/TdWTMyGRy2IbtoB
J0e84D73hwEtMISU0pz/f7F/innfpnZQ75sZ5iaTGM5TCfpT/exITTEbg2QCqPf28F8S+LtalrqZ
Ks5UsOWTQYN3wQYxwtRJyYmiJ4GrtAywjH76p6r5LkzZto96Q2Zo0bJWPMCb+c6TZxQwn6W7A3rB
SBlto76h3G27ShrSDG4X51t4MDkCBxuhH3GfVXv12gibGJSx1n+dEq+wn/zM3EJW8g1Cp+XNSs2o
58uTZqjwtJoiYa+C1zkCCpGGT6xg9hNs+KNsF1GvIxj0JUJoeDbWR2viZBB35gGQKa7F5JsuLvTL
Z2ZSgy5qtCe57ybj07C1NRa0nxxPzUv8CMVUe7bGkPfvQoHMECAi2LgPCd39QdWDE7MLvOcYQSr2
PKQ/fq3TlWxa6I/h6zEDJl0NriWU5A2bB/c4b8KIbjwkNeUnDJxQ8cIygVlzu8orBFgTU5orGqQz
vS/nIUjlqIyEE4Sob87bmrccG1LlW9i1OB1mG+pDJetUDaum8cP1PqZZHjwMJkDeBT1pZQRg5QMw
7rdjZDCgfArC9CP2vJ0BdA2eUg9RVcN1ECncby+JPyMmUNeRrELTFRTTgzOr/PhrNdFPFHRDiZde
/lW9kk6oVy+xLcR/xwLpHRoaosThqoXgGvHZ9ybNZvT6WUo3LRkvF6x+tvo6KOgQgTCaQS6s9rTF
KoerpwoFiuP7YgWQrpDmhQFw6sTaAz3vUSLk3d+HylOd9r4GAh2LcNV0UjLUBojuG73Joad1L6jx
GBoK86nQSHN7DgcTeoHlknulrXEIpJiM35v9aImOLhGlVtuKfgd/jZD2n77Rpa9CkVVoB1+c83rj
xaPi6MHz+mzroeDCjrVLisbuHpq5OoqbwZYCJTTvGkaB7847ARaJr6VRb+4ok0X76JQBjrdUje+L
AjMGOGWRaQDz7pPYp1kSw568xb/jxFzEATEYiJSHrJqcyDl2aTa/rApDRvuyqbso2abnf4XzOv72
ix8v1WIRXBwxyli7STioBWil3T9RR73xnbmA8YQl+RcepEWRsuLLtfLWn0u8el1ds8/FiZyLcjFE
wFdQLeVuNND6pdwIVDSELcg++M+oEnbpm0LpOZrR5mhndDdlBVfH1Bo4FwxLdW7fCB83I62lXDQP
w0X5yeOBeTmf9fJcl1qQsQ+NANe63IfbYRHFqXuEjZITYozBFCkd7dsgeGhG7+TVDOMP848K4Cud
6QUWZJ7NY7KQwmpn19XCuzui+9Co/xhC+hspzoiqgNW4d2ilTPwjP3qEcNQLG4NVDqk1/z7s+qZ1
S6VK9sB2tKpohgDR846tksJLDRf1a7Q7iMiJtjdGkDzIIZolrMJ7IM6UZDlgUtFRlSgCPcWsqsqn
l89rT4Y+cm3Q2mDPpMDuw3hb037SCyhgRFcckNUMX4e2R7UUDboogOr662TmknNGOpO1h+lXMLGS
7GHCGnRg2i3OXbO3FValvqdKItRXUhddyAqjyOakV32PJ1e1Pjeny0FbUjcuJDS0+44FIKkIYBv9
BZkIlaSBPFSkkKaDE2IIP51xOITIjzU9sVm29vv5dU2eimUZ3LGo5RWMr4w0pzHLL6C6+4ABS7qF
GobLfN9JY4wytCBSyMHqYKP64jd4ARzKtW/5r6dSraAS1bxWK9dkMLDg8x4EurgujstsayysGJ/8
pECmWIVDL4NJDhuciEKUCTeZAquLX4Qgxs+Dq+OX1n//+SMmkkHluZmQHI5uOa/YCs9a4+Ta6gHv
h4sfQ6srMQw2ae7ARxtCEiBNWcIjf2w7w58vECRPJKl1ZijFZEVJnwHD6R/f57j242F8XaFaT+96
C57dUZ5NvO/WO1EbtWmG5YFpv+mSwX+VT/Di1g/MN172uzazmAPlmx830mQXkfw7kucTTGla6LVG
Rc0FIwktCQCp8jCVit6//H92v2I+mVojLNksaTw8GaoX7QLUMiq6pDDIXL56pjhbpQy04pkmu7mc
PRiDpNiwtqlObNH7fs6q/JV+ruK5fHtHRqPl0AVLmIbwArBJaHugPR4S/H5rLcBwayii0q4mC0WN
3XBFwZ7hqlDkFyHtFulWQyJXXlSBLS5hT+FvROMzV6LCK527CVYYxWK0RyBot/SKWgjf+hIeXamA
AeZMoSTGkgVr1msDpJ3AqAZDTsHvhm86pOR9RMfconmNpXxQp8AHzR5Zy5lXUzW5btNloW6573Ml
Srx1tROnOzTDbHKIaeSziOubCLhIT7fqeOOSrqvZOWfoKxjk13azdOimCgHWKYIwEVNBXjddGgG8
VGXqYLuhHkmgD/eWbs0m2iWmzv3zH8UqDQssTRbXQ3qtk/m1InmarR+3kCdydwUiSzXVPhbphd7v
TjfpVoO4yuTLj302mhNB/yjsqm2Xdp3WectyjKg9pKQcftFLQaK9Jwya3CutxsjpyMYDGGmDUjjO
iHFNXw+ZnrTIf4SBh6EDxF66bDhUlAl5ZpbSx1RgHHQV8UQ36JuB4/A+ihi8WH39F6yLg8TnIY/V
oD1rC2cWRT8VBpRqr648Bl20spSJVnqR3u8k7N2TyghwvdSFJZdGGVjtIVlSsCSKCscJOjGnFJSr
xsPBO5jZd1TgLPl+a+QjbbPt31WTpxCfYHCiQPQ3pFrDSEU+wMP+u40SWfLv7B2kSIAvwQQWyJHV
1qoll44hLcUBSWGU2/BV1y8anjo0IeL1l5dZQYjW0UNCCSJbijjhm23U9hVMLhF6gW4QIsmRLDRd
Yo5et2lvnJDwPgunlbe2ixrumevqwcR8vgWg6a/gBpUGCSTMkCufmwAX70IBejFP92oKofxi1iOw
xvG7QKM7V2algF2NzamSJUcdEECBvyBH5MlhbvJiHCXCAVdm09i2AeCDpIQ5EVgtWBZCO7Gc06tK
NtEewYjY9bdyU0gFmPlYNgnTTl04YLCJxzZs6DOri2zRzbVFKEBoX/fw2qYOb9C1L3Kc55+Vdx9K
+VDjPVJ72i8krqhwmwxkURvvacV5nlBtrIXorfdp4n+DfMZd/lobgCVbNqsD+hkwi3K5tjCD16AF
uqKeWBjXy6PgtI8ljfcVdT/EejlQ/dBiR0+Z+ea3CMMUZkBmmsaNhLtBCsPk8msF3TVF/JrLWsc3
gd3NKx7L5JTheyRLEvWAHvBNbrkuL/5L3FVaT2c7qxXNdUfYx9GpV284VsJy+dy0zX4IHbOrL+fV
7CTT44lTpPfQSQ/ehhEyWU6i9z3bN02+q0MWfIFJNVqMRoaoEK3XOCGpqIlxPHnJBsTo1YS2cBvM
XS4jptiakKLn0ksC9QysTjllk0OtlWVXsGFufGUCLRBn04RxQCoh5nfXx1xNuG7E8M1EoFWmVGG2
A4m44hSFNYd2SPYj339cSeA0UiRqghHajJT0pVYoJK9xrAD1E4GJ34na/WMAhcuUzus8Re6530mG
RLtQevsbMqnvEdM6K5Ws9jnaudqaJuRN9GsXoq24E5Z1bKRWAM2eW41Ku54R138tDvjlo8xdfF+r
CCqeZWbzqL4fNLphEsTfC1BRngmYs9uspa7TaKH6WVhTysnSPedv439KLK1ZU+NXL4OAPCESYV33
e8TQw9+Wuw8KBOcjNjlh7HB7JbWhrSAA69T00eCU1Cfpk/Kq0WnniwxiTNBpIxBytUOp1bUlPDl/
x1UPWDRD2Y48m7mFgSwHw4Dz3lXG0hFPVvjWID1aiCBS2kg0LW2mhpUKlzGQ4YoQhq6/MR0bxj9C
xtLdPevBjlgyMwosYTlYkx71RswHWx6pHkSIEDsEk7f2LNH4dFxZiOCxZBwbsHWL8cJI2mI9qmGh
4ArHA7OPFhU0997oq55dXXJOWx+IkKwc8KnUMbI1GSdyzYgQ/xUPiiKfllFbpAla5/lxFVn1RC12
7v0AVEfoKRETC6vpV/UH1wdP7oT2BlJhTEp4eokCevF0kQvk6mz83TbilFkp3Rl3WjTGgRymWqt7
EMOhM1hjc1HOIC1pjqieRZB1smO32LsorJCMX9ua6GbdTMARB7bSdJb01KMNgoFAVm6Ghl/JHg6I
Xzdxic3mau1HphxNZX4JsxjOmPuQfjo1zyG1pVGMJuqcyn7D5YTK2Wx69YxiOK8cZdcRIQ9pl7Zl
dDihYAkbUq/d3blDRmxk3ZgL+kvtj4e+ceJZUd4mm436IeAOk1kUraDRdsbwEmLdaqZtKSGnBA3i
Dcigil+tYzfUoD5sekL+lFbUt7bLHMENGxUllsawyfyAsxjISyDd97u2EHquyJL9Laijm4oxMD+j
OXCnMvYq9BgxH4h2MlsoZlc5DUB1dVqmLdOQpmWAeSJ3mZZKSSq95DbHPB7w6ISZqv/yP3oKOWlG
gqIIVeJK6JqTs+TwguVNgwwpek/E94JAG/MCujwnNIUK1LxxJuC8ctatyFqo8Zn0jx84NVwaskK+
pivKHKh1juniOGVn4my3/nJLIxBSVkZe31Ok8l4+N5sOCC/6fLj9HlhJu5sBTYkTf7H05aUUaAo6
W2oAVu2QhZCIluMhSp94dqEw+iMTdp39RsAHLBjkAqIgby4qVY+MfP928zPfwn0KoBrhGiDFBt5u
EqOlE+rHfKVEaiAMcEpQBwrF9zf0/UxxkGV64CWCKohkliwWQFFy2EJ2gL5JTfD26Uw0BUMo64Xc
Z9B+GJ7SuSUepAtaVdic+u2qBuoGTTyZ1LCTL7xS0ttFFAvIBTK2//BbohlYkIKNH5CjJxIC5BBs
v9DEvnfXZCVgZPJaTt6lwM4SjNt+y4+KXtvqFie3VBlNboAXSju6iOVRCzRCs0eWuw/XCCgQbNhj
dW0LG8XlPBnjsN39j6LgJ+aicLwRtXADLME0hHOrpW+n5PJ5muXbqtrTzp0DKUOd0dpXkD/qLxY/
V9uq8VwNHZtCM5KFAlhFA7ixWm4+OI4gffw+Ta6qYERMNDPfqAGAL0znQykB8w0VMbRhkBEibqzt
DJHkuebXKkY/WtW8PqGjKriHHZM5bsAsUZy44xPBHyIHzAdt54OKU607dWpKLlG4w8iO029kgVq8
GJE1U5iq2T13LoTi8gfyfnlqcpSP8HhcISSq5oQwVoP2pOUp/HcTh8q46p6XOfBorA7iVnZoNTLt
40xB2xQ/ARgM+1U1fwJvChbXgVMSpSRiGjgVVMb9GbFvtiCdAEpm4umyTPiJFAUG/6BpfQS3/Oq/
j8IV7AvbQTgob6flfPrQw8kzWomva5hNj3oHB/yYGTOLG3mxXPtVItjM3NK7tmYuZuKXBO2n2cSf
KNv8Gid/ixwHiaRfZdbIJ5rKGc9UeaA9/osflxp2lMZR1C8LpaHlBnW8PMi8E+k7YTT5NMBNJofU
0a6ltPIQnNw5Tz9MGDj0e/r84PTExb5AGwZYP5DnwDiSYaa5fqfQXTgnLaye/gzv7geBo5b5f1Lc
CrpG2Y12iBTws4aGmD239D1vGLjc3teXMbeXGJuqWfkw1kJsaKfe/iYheNADV2hyzIK2Dwj3ikj4
5XRg6Xk5tCTzljHCJddnl0Jmuh6wLu1orIidQpKR0/ysc/TGn4j1xzBAJVxOG97pfyIiawC41wnj
2Pdk3gok1m3IEuPAfIeWCe2idVJxAxPws6/KRkNyFQXeVJBczmSPsqBN1lcrOjXMphwDff8pT+qT
8urP/inbYHO2w0NtHTP4uPQcS0r7vW+I62bJrVvV7IgR1TLqAZztWQrJmzR7R0cC4YiJrg7e2MWR
igGxmOAj5DkT1RdMPa2rRv5DOFcCKxcMlh7Htd8HWDFT3qxXS4kXQYJ3zZR0lCVc3JiD5w6mRf/X
QeiGNR+XfhObptaJbLpMHgqRgD6enyIBgC2yLVFmOTWS9GBHkJkpPS53ZRwFmJ/xJXc3CdO31zLx
xdoR9UqkggxRZhGVNNefGki2qbf66VlWI/nFZGxqhqfZCz0SA6bS7GS0N31Zb5m7Bk7GnCLngK9q
YcE29TAlmnmif/kTegKnTSwROpwt8fROliZokojrJdrCO/rC1QdGmyYkJBmMTBX82ATZaNPeo2Pp
FJiGaesKnyU01eFN3S3Xb4380FyOEpgJ3AIlVleA9NLIvf9OUDJCfZi1H/FmJiALRmaWdHmK/Y0/
nHopo9MeFej2u1EI4OnnvuGQNkuZW4JfmarMu7KlJSAUMqGQOAeFpbv+z+p7pclH3nVfuNUWqR7N
ClvhnbEJ4E/owftQdMThV7E88os3ufMkGlwmf2Ygq2DfcZJP3Xgv+ZpVQUoXbd2Ewv95qkszOM4Z
A2zUEQCClms3v6Cq8OeqY+nyeWZyBAtMC8igmV34qHIqUD6LHD/1pEOd2Bsw0GO5uaVClFnNgD8y
6k6ojiyb2wucJpl63JRVCSiOrFsvANNtwCsmBTKkUWkibtkvxkTJy78476nEFTcV/sMudiJnYH/l
MlbQB68wBKQx+p4vlAKIsHtIiMiFDiv1APaG8UX9viLT6iUsow+zbYt5D8EPegAT9F4c8X3+aDbT
GyvPprh/AS3Hw4Phi/0tlPc7etuNHoZdETTj0ZG+N7MLILqQMtHwkQCob9U+RRma7icnU87qpCL/
5Dg4HLf84ZJL/wPDIVU2CtR3SV7soimKZ9LIBZ7aoSlCMLPiIOMki+TTH+cpp8uG7LpI6QdRxg9z
VLQOppswnwB9ynfC2+g/9/b94DwtH2HFsAowFmSggF3RB0iiUOIIUhVdBL7evrqjU1nVK7QARFPG
yIfqFCdAbSGVwVgdbee9eVrpFqN9i4ePeV7lmuvNELY/MfLvcr7MZhE8CkIHXHdywZTRy7Pcq+7m
lyLa54/EqPUnMMgzer8qrwAt7PDDn8Iq6BNVyKIzN4kCHfLCcK7MCh1+9dDLDCEHes+2Q8k7qKmx
MpEV1fH5P0MbqO+h6jFbpWtuAQ8bC8vIyWSxdkuHteeY5f4iQkp0e0+xkGs+luO4X0chnn5dwnh3
iT06kQg+AcTLZt1TO0pE0u6thWQmhG5PGmfiAtR7bj2WKx3oUny/7qhjVZgGqDRkXpjthG1nmCUk
2YMPHhH1u2DGiuMI2S0FGjus+wNtonnz+mUO2SXeb8GQxX3RA1q387iG7h56GHeZPneIUCzVf2Wz
rZeFKkq/6Ga4j75R/eWuPL1ril4xqAhzRV7vRKeiXPKC14AWwZebQjzuAL8dHeFwXSR9l4I5/xIR
0TMT8BMy129Tx8kxpGswwMZIa6R55fXQl1I+QWCouellhvTeVuT8+Rhmzqeq7PqlGmfd0Vk686TB
YnTh/kZEmKhM7wXEbxL2fcJBb4KalaQVicmcRk69pqXL67cObVU0oL2EmclF2sFXT9AIGf8XdeHw
9lcf7A1lt6i+pM1glFZWkUwbUfk1pzzOZWTlYlJXHAhYYylrOkwq+rLIx2XP3jaYdu/HkJRvwF5+
eYV6KTG2g1AwkS/INGWyfRIdTqgw2i9T/JBRLAk4IgLhcH9G17FYQS6k36N6D94DgPRrOhnslKyZ
NPahfacEoj6DvzWpzH/IjD3KeyjelRCzZE+5K0ABMaJEjoEQx663yE9lVWOEtWOKaaAMN78rskVt
ihZV6XaU1geezkDEIuAGb6wDg6f1dO2uJY+CjqLFOW3OBJkT0oDMLzLqxKcDSu+75SBU91NH8Fpj
2HY6iPcawj7Enl657zZs4wNrsOOdke6XGFdoXMi6pZbodCe5nmLArdrF8HXgJQQUp8Y900eWG6C2
k71PXTgp7zGECevo5vq885jDksw52yp5WVMjIqhtsTW16SQ+EQ4grHSWJcDUNOEg9cg7HPpjbeK1
6ookxmuuuXefaURtsfLeyBd4ZJxR8fcCxzHx25YkTJVyeLqzq+qbzZDJhBzdf2jjsFf7zMHRa+eq
FqGsr2/kamG0VoXJktiWpL9Tl97R+/K90a1ivuXaDhdLb4HsJPM8RB5p9HXXEnoGiyli+gpzokUx
oktls5vbKeyvLh/6+1+tVI2s+ylgjiuKZUJFEbspfGjoN5fyS1GOucmmMuIqfRT0TsA6DKI2Nabx
edJZXm6R4BPaFjuq6nJh1W2X8Op+P1a9O9e9UyGLKaizn3nAxKoWXvSjr58Zm309vzsZQepOUymR
Exp50J1iKFviWD9ZHkhrC80QjZtvOthEGvj+hPqmcgmSmC6HryR8BR86uBybvAgntQH3rSEHBvG9
/RNSKq4j2ICw0uK2E17RA1S6uNoE2MPR1ix26kZonj2FRdhvC9yKBjVe+//ZsUKbO46P660HnlpF
ccHcziFXdpgJ0fqKF3reIvE+NGc+4e1cJSSq4N7nzsizCON7ggd8SpqhrEjdzu2AEnkxcf8QJZS4
darMrlSJIN871eVyTOU8bpFRI0tNyuaYPLSKkSBmtyVhbzj86r4nyAF55veSOVcFgT3xToisznKV
pfFfqzESTSmlaUEQ1AtjGXIGS3PXxkB4ew/WCZltI8YaB/DTPNr73/wXHfGHzNpO2c3BnM8GTHVq
H4i0YwXyeQgKDo+YGW+EONGD/3eBcNV0KLkbThbGEJJk3hqDsJN4ydZtNPrXHKkss3fphJCKJwWv
s54O2DHVXLgZHua5viAXzQQHo/Sa+e21xIGgSYRX6zhhzZcP2hKq6i3ElWYjChwTYMKhNAkJGc5K
dVFbxZKk0dp4E6efmdz+nW3VfyGXO3U+TaZV227yJ3GoWLR8NAJkCb0nuo1RPaBN3/cfwO4em8e4
lDc21a9/7yoVcntnEirS0e0fXQe9QGf3Fa954iEJ3+GDh/2a5df/HeUHQ0zT7dF/se8/dU9s/PEn
6WatKLfc2Hl5aL7NqBlXJhf6BS1OTclhBJqpJM9q4Ug47VXMqZ0di49r2VI/K7xpQWBCRjNNiRZf
V9ZW5oUpYRI5CvDP3MLgs9h/M8oyqVuk6kPekDoBcGMDRtcjgbo85ldAxwac8b157ETGZpuYhJtp
wh2AWh+W18lLq68hxZH8BKXLN2WtFJt2wNiBzogQLd7h7xctNDwHcyDvlag/QEkqlC5cSTfMkzi3
6wv31dCRPgQf0HxQ2gbwE2WM8VIEQNcp9LxNFnsKabLf+JHkfJRJ6xHULDDZq5vuiqyq7GPGfU4q
Ltuh1F8SVdQu2tqD6bZrxZRpnzECP6HY+QzZYIFn5oItHaRdyDKao2wyGIElFobLrQDydeBuDLsY
CxduQp1UWDlzkfGxoTWbOz6uXgU2OXQQY7LDGa0C3sCuaxPrkxll3ItN1cW5bMr9JEv6w+qV5YL0
f40aCj1SeMN7ozG66JMvWqpRmCwwHvncCa28gCwz/j2SHBC5u52/wcL74dIMt/BN/3dVSYV/7yFu
8wzBJpeqhNoK8FWATiNgAjhCHytGs9xQwcwbGcKhtH21d2f/tpspBLa8QeTkhdFinU7y8kTmy9QF
xlRbUeky0kOay2GCU2Vj82QoQ83ebmMOq8Iel3F9LceGpq+IGFKzmyBSwk4Uje08pi87ZufAbaln
RRhvoIkI5dR4ZCBxQTOgJ+c6hmS/SigzrBzwSdIpy0MAPmwYQhArT07/yu+lQLOvG8boTv1Yts/h
ZocGJXdF8q4blvNz5lJUl6MbJIWZ1bo/WPu7JRIYa3F36X9S+uyp8/XCIJgRHTDx6RYo/JQMP7sI
PSqBoREssdL6Chrc2baBZ7V3VlEXVVxgEpOPyk1aCrg++pR4ucTz/QYLlwke3Uhpl8Yi7lIwu/Jf
6cjAzLL9sg6IU/Z7FBjn6C5FEW9z9gb+9uUoelnDBA1oVo8dFuKfYP6+GzW5s2UveGfIMfg5W7zO
ruf0vsaAFLleOFtUhMi5fvolTLHvzGCjNeV/45b5Qi6AjTWwFgLjoP55iDsfvz8d+YkgmzzjFZon
7K6j3TvDSPz10wrxKButb6bCTwUpE10vscx3fTH4q5GpXg3hrfkwQsNTzZM4QqnoGkU/Gr06Ma1s
bv6KsLCtoRv0WW4GD88XU5v+hg57IeptRDSMvRUG7SXqu0ba83unGuyDy0dHWjo+x70dU7FDGIXG
EEnr3o4DSeMbiiABCovs/XuHtBGOJc/vJHn/JZW2aN4fEfHoSrHBOveybSbqCD9iKdvZ488xTMaM
XqyHtDrE1hWs6d9h0toYS0mdAYxKnJR6QrgcUL2Eiw3//QkmldQRxrAmcKnt80jkO+HWEmzxl725
GdCzxc7oxWuJmQ91QJV5NINgfDdQH0RSPPRGr8HHaH+JgZi+juA0G+1JwpnME1062q4pt0rHI6ja
f9mQbM6UlDW/9JMPh4TihuT17TgGLQTrP+pVdbvDtOcem9JMsEWMwqd3wQULeORn6OtDeZBAd9bv
EgamvYFwG/WjYi6g6OYEWskN0aN0SAX0D6kOpx1SMYI2/3A128IABpIAyB21lfodfaQndLGjb0eC
NPo9FyOGxfaGICyDeIiVrr4+SsVFQUz0e7nszsFqbVBA6eSFHPvFBdn7XG60EPGj8EXmFGRVRSAx
GZQ5kmWv7NEV1u1er01PBp+5xsPW8wg1lRHCsBEgTH5Ckyai4H/AQC4RfqRQzrJUNhnyh8/IjbDT
7thd+02ZIpqEea1PFcxqjrWG7IFs5ccLnAYIV03YnlTX6JSBR90YlDT9AhxN0Yb2sTsno8bjpI+9
nLwjxIyb7hlh1iurVKWby4f6RFPvwl59l20Q8uZeK10oE3ZLHk6jyXea1vR/YtFSwUgdZbD8X0MJ
AgHHEWLceqfQrV3WsnCfLESEwNCgGACsQDv9HYiGEjfZNIwXBUmPqlAjaPIGlXl0bIaPsThRp0YW
tkhb0hPmT5igJxvrB233irH7cuP96YVSraShdhyWMCCcgdYZRWUoRqgtMbfMu9BQultkFsjXkYDM
waxlE2bm7fGeGP/40lMmgK3tUTuj7IdoDnT0zubUGiX8r4oyMzLE0Pf9AHc9sQrVrd6wZp4kxPrT
oxlVYUlSEkv1fDn5vdqikNnFhyPGGvZUcAVEpvTecH2vYHL6iSWGozZukgzCWuNp2S1j+qDqRWNY
fSBYTIpuAjbdbPrF08hu7LIcfx3hkbX7QX8pja1V7Lmdq0nEWTNEyO5PldQtAuVOkUs7BKk4ZpHa
U29s8H0O/Dlge7I6S5f+DrV99mdLUNUmpJeUdsz9IC+c5Bq3LpZV7/s5+Os/tP0Q+UH/93fZXHua
xWrTjLRMzETTZe37Z3ef4s0DTC/ikZuqtb9tv3P1X+X1LGWaiWrvocb0eXiOEdBE3++Vlrw3YAMu
OoQ5IcrDuApyp9VUGTnxsZaX1ChFZsKipmvEDFWh9IOBCRJDor+zc5x19eJgkKBaAos2PXjPYihl
0f48tTvuXscu7ErRmbLEAScuNOUy3qE50dQRZABdJMi99zhDMSh79YNu3E9C1ZtjHgcLTuFi1r3p
1ePZaKHE0gKWU/ikoD8XJsmYey3l04lN9hvAT5LAOBM7w4IB0NGqkO4KtBRb88BGJrBPs80Ngwdo
tknL6WfxNXDp+HpmRFH6ftvZxImVcZvQkrvdwPdXDAQ2PcustN0g4oTz+f055nhVMtshf4k+ADri
0dgzBZvNdewkrzKvaz29+HkqCOq0CI3fYg7mO18rsp4z3PiSYbw03nF15sg2FWegDvfATwmesCgO
h1FW3gndkQF/sL5fV2jvq75d/uwpVX0UlWdan6v1vTGRPUEedyek2btjbr3JEOn9UYaw7XW6USg4
Hv/2sIt5U2gH2ct3NGw008y0lzz4352ArkE1xMvzYdo8C8mFyEzVXwjxiNM31dCYkkIZMCbnrwfu
wMru4qYR8usp4RmbK7sKO0HuWf/1qZPLqTABfRL4MZmKb9dwp1CaUvCsHTqK4g1MVfGDzq7/SUrH
KEtMTTMfeKR9vkWasyxHN09DC0Uez9elau9Hgpam5qTkZ53J1MjxuktWA/ZGgZVtRanlukHUfYVK
Uw+WEs+vuOZU8WBoVMgqEV8W7edps0B3S0gr4qEkYyhcODzoKOMI8rhDFQ8kMJEut/W7eiC0h1Sm
iQVFOHxQevwoSGJoOhekIIzRl3brTqkfZKpBuRdX9yxO/wWHRBmYOs2p05m/XGwqL/Qh9aKW6ObT
2SKD7mYqahSCM+sNSffP72GOK/haho1RJbTGBjmHaLNLvoCPs0gQoCN3RFm6fV7LFX1/YNzbEUjZ
ThpnxPqvpIB/jlY+v6Oawcq3LnOAYY3j471hSP2RILlCl4nF7qSJ8vE4180N0clwOl4tmkB+BKPk
27j367EAVHTMBBRC6URZo9utbKVI38roy6MUqeeLk6CyVg3QsECS/h/3XyZXsqaNeFBZxAGXIu4r
l0+fNuHp8g92lyBLlubVJX7pdTvACCYPIQnPE+x8FsyApKdUlSJBAHxZb4Kz/dN40AlBNhMBTjMI
YxVsaaCY7Ofv4p6JI/oCWmVdDHQqEvj8HSnrBcu1iWG+eCOOT262/cU/SUAWAZtvEgB6RXTQrBqs
0DNwRICq11EeoLa3kKXRz/siODT1ABmjJ1jxXx5x7ptXeCaX7pDxTv0MaSO6vRZQbzwlImCIaaCE
w+HgeLn3THu31jyYC535P+qo/Gb+0sg9acnB038QENCSm/ihtlWe7+XXNWGGh9EpuIUlSWLvKYRk
UGjzyl56WHiDjkKaays+2I4O5iQJuvQic7uVs0yVS8jpeFRrTLagIiWsMBUZ50pyioTnb9j8a/Zm
8OFufPmlZ/7WkcuDVmTv+uFrdzkprZfQz+zivIDkGv54eWy/cFC5MuDyWcLeBKbex3dhZE9sIzsF
1ehO/p7v2sNaCizSv3obekw57D63N9bNlEy7GR9SE4eWzQ0Z/8S9Ummul9RAoLQy4B5WogmVu4Zp
tBDDDR8rquQp8nEcKIpjT7xJYY2B/v/lwwuc2UVNz+SIESaR+nYHpp4IFNX5z4KQpRtSZ6AHAgP3
mZYScnX1ch6J/04aJ83Q7uFTBywWKWP1iRSSQPWcIkxhymEoqtkYh9cRKmFJde6wC8VHFq/3Fp4b
Ihi7r4pbPW/NRa5FEJcMDiSS8dNCzNP1rAofK497NVFpem9kyeWVWA5uapgu/xukyL+4LBxtjtHp
ZeDt/P+2hPPo7YtjXKaYm8845KwQet4Wv6haR2HbxiMFGqKBvp1WrfKovURKCvCyFslmrHqNA2Iv
AHrByEtpUaaemsI9bxjSUGbOta9c7vL4qK16RxO/kkQqIFGw7hiIDfP2DQxksbV6g/x8VK2lgy2t
rr6jHNmTX8GNHJfgURXo5AzstkV0Q2kBd7Mik+mGMOfW23QAIZL7VnOWsKS+7QGsXIm0nMq7aLq4
Xux1WHIUkyOSy2fg9Cuz2sTbUnnQtOifjisdVydGC9YGqlsvuvpsH3ZKhvRr27mFvYprufPN/W3t
rflLH2fdkWVu7L9FoSMWEOGXbTEM6g1ZTa74yHcafZQai0J1v+Ahf8wiZz0U1bWV3HMlAuVge5pN
uf7Mpy7+qsXEVxz/SlSGdW2tm002ZC6sDmbJPooPOE7z/zygq9/rTCuxz+GNHyfw25cyyNQlWsYD
9C+ri8+8bvJbY4RDZPMSSVjp1Zk0mYx5+diOswOdh1hM8/lsgks/zGYABI2Z+iws26wJ7OftUWwZ
PznJ4RM+WaLDd/8gdaa3GP8WMKrp6RvuNOIH59qwdaA2lB4SwYhvOX/EhbhVwT93ijExGIlaFYZ/
BhmZJcnL2h0WsQIeUD0k+WqbQFRMv+d0g5iM3h0lEKn4R9ZDHYK5s/JUQkI05Mam5EsRvRyQHVcf
BnYYaPbxdjpg+lWKDXFnOgFECe9gqR3mnHl4EJBZmosgxG2g+HBCJhAIZQrRHazsXKNADC5lb6tl
LNYKHv2mT88DNHC1ZZMqgBe2UqQch8/1smrTGWFLRuUxPQKwu2tZHfXADdOSuh/U352hQ9rv5NFf
q/fMhxQCySJgpzBFEsHAYj1GGGl9Q9cPjl7ZiKw5vmJNsKYk35xAiZVygL81FD6489zZ4jPn5DZx
+nkVyvyJJZ2oJAuTa815B41ud781U7aD6/sfDyAMbXKJ/ymAK8kSrylCHDf1vbP2MtPI0QtcG6T3
NV4nojkVN35HHAqq9HVc9o9/97DGC89YLGnHJezC4db9SXioPzPAC1onVHWXOMwqJlFQpWPJ7icE
TDgWvEA7kQ0iXVJFClJ4MCvzcV+plpJAumFOk+WFIAjhZothffI/1rVh3xS8jdB1ETAXFbAN/czr
rIOXAebmwN6JQpRgG16CBUZtN1UL6429uwKo3taQaA6hF4+bLadQf6LkMLYLyf0ox83f1H711LaW
+kuVct7+deqUjy61OgK9gK5qCbKolorzYa79sWE6toU23V4D173BqaFqTGvZZe2ZT5hwgxR4wYEO
c8r7KGTKJ9coqQHHr4Uh8+MHX49bU6k4OHy+idy8BMI2cP5teFzxpoDdkdSJvuvEpmup0waHwqlz
LkmQVUc0c4ZZ+uEUtPN9QV86Wzhpz+qBju7rravv6EOhaVJ/hBiR8LEUpAmQwAqNRVndGzZTFq4j
GvBl8A/MowdRqTXRF0G8Mtwmyvvm0paNd7BxIlrmUbySWB7dOQjvXfaq7xkHiSsAaaxu4rr2UvG7
tRQ/kR/g3yT6DDcCayyjKItS1/RQvXl5yPZU5bpSj7CoJWew5hvA6E4Q7RVBx+c7lCK4XnkQmOfD
xNXCApBvXcCVZ+HMV1/E+RYYqVZie78Q7t8k8a3jpJbg3T8NAmCrJiIUt4AG5Ek/5LJURV30qwYX
AGdv3enOfhvG7qrp8tDz+Th36ixN6gag7NJj7UiLPhHlhkl53ICKXY4cZC7boK3YIWXn9K/XCHMK
lG9PFaiZa7KKrFpchGJf93JxKmAzHQb5/INluyJqzEtFGOLOrsQ/0n1cEq+2C7c3nw7L9B/sRIwH
VK0JZWiRRGVfwy1xlCGTT4z+J+FU/MI0B8TkzAXsxVUjF3H8SbTPhIZyav5p9GnDVWnabMfAyz9P
+WKjOtpZS37vsHzpmqYC11UWKls4BYKIptl7EPMUGFj7xwvRzRZJxRiyrQbUT/2LJ09hLRlxyMhD
1nQpWjIpEW0iy257kVwq9DvvHh7T8XUna8bm2Ubh0rdGzK7n2KaCWAkQ8UAZn2JvawadBTgJVpEB
fwmRYMXY7Aa3i1f3f+nPevmPELndukFPCvTTni5n4vWtkiOvXsiamZKXCfhYltP5+6qhKsqb1u/l
Mhjs6tYj9OwooDs9U7PfZIz+1IVcDZGrl/UuCD02GwT1W/i7Mn54CykFRqQbhqU5+bpeiDWBZDrp
vBLLlU45gMuBNRwnuRRUAboFom0Kzp/yhmPbPUzUJB4NJlKcBKnXzxiijogHQ0DzebOYD9WhSFoj
MO/12pusjD/RKa9m1ve/T5g7ehpSMEbaaiO3dRf0zGZQ5NnDBZQ9wyLpgzdeOpza7pRgULIYr3yS
yGZ89K1QQw1j7IM85Cs38VQQzx+xrLnjlQ3Zyrm/7RUZs2RvXDQ8iAEX+W55+iUwtdsDDrhfdshR
YPdBD1Rq8kNAdPCu71qD9Dj+36gNQFXiMot22SOcjOcZNzqMLzKu9ZSI4KfcfGaC0BpT/EiImbrx
x8PAyB1gzr/+UsVwZpN22QmKhfbYkGhWlBf1YlSqraUJWwHoN9Oyqb9QFBfN25gEr8K/PQN+DByC
HvIhH3PC0+pZiFKaTDq00vLx4CcNogDpLcWmDTsjV4KmSY1f9yQQax4InpGcuHvZ3YX3dT8kNJXP
YIKFjzf6vdDmGacPi9KkVCO0/oxrwXMfabRUf0VQX2RxGPyieLCPQXqS8him4fwg2Qx5MzoF88Ce
Yotn6vCbTi1iPdKPRhiNXpG2ITl2zMMxWYBkjwj5doKP15qT5wOHGklV0ASBG/tpzzUnB0FpTWvw
AVioQZ2adyH32irkxdlbW0JRB0eGIVjgxTIFD2h3SEowrj61hpyFFAi/pLeVnpM1f3LmD2lwdbDa
yLtL+XhcNXMxuBxh6FVyruWPe5fwfVz+Pz2jNecFvqN99qn0nZm0fic0PSuwMnDjNAJc1+eeoZKP
dM0BKc5xGb2k3iM/v0c2OAtOFqDKDnPrZHHhgf7revC9NcJjSLVDBXIob3xjhsV+XM5fAwboRL/7
Q+cu+n1Zw1x/tnQQPEJxkgAJNAq3D45Izn6bK22lNTRxGaNnE5Rj1k5HWnKrsizFq4ph5w+yU6Do
0bBDE4VLyEFGTzZjPB3+HSCPiGCYUlQnYanfTlDYCAAoRH7VwKslCz1bcoDYPpN6sHLgqbYVY0Vm
i6WWCgUiiCCyzIaVy+pqPNEkI+Pc2a0v2DNcz0kHw0k4U6v8RK/ukzyphkIiKYQ2g7qtf6flymDf
FGbDVkbOWJq8oxy8yKnNhsz5s2SUs+1wxUWkzRMUuWvrj8XQaFeC52INGEUEnUUnTfo9dkedXT/5
evgEctQX0aygT+lolHwTqoqXZF+cQb3Xy8OPUkbbWCwrJV/6DOyW3YNirVLkNVvJ/6bNkZvTmZd/
1WyhsEXMXppQDcj8+YnELujTLDoy1bINcUf/i6IunFYbbOSSMp4d1mzTXDk/yTQHaxL1LPGfbVQR
Mt02HX1p7R81cU18Q5bhsJFx3ZcX910au5udRkzggOgFb/VKPMWvN0ufxtjA2Y1c8K8GzY4fGoqk
bJcYhc5gxQ/oumNUDJqe37JUNhGbPGlpQMqymkzD5CaKstIsnEowWe1LofCS3GmfCw9ahWu6HGFM
t4mJRW6lwAqqiMjweAj4RUhyfyQA6OgYATIQOZj9ZwkIJMm0m7Lm0VV9yA5LrZWmqv34bUsEYru8
kLbB31GDjkqZHA+Zw91VnuYqHLLM1TOUDE4st3idxsVcNtY4O+YS2zCBo97zcEup28NoUD33mqYM
gj6mE3YXb5XwKykYveU4kn09HPW0oDEfmN+g0D5O3mqTJyZagay8dte65yxbxCMX4zOXsLxwY5R4
zfBKNFwNYbAxyZet8tTs6giy55pyMW0Txgg4hubGVbxStmciPqsqq7UrMLXBm10tnGXtP4FI9XKa
A7hysg98KV02sfqcCCrq/idHxTRQbn1/sT39hPH4UKFA9AlPgK7sFEWv/xJ68OYimrtSOignjTHx
fGcyvoDCIc4JiO53+luX/9gSAlwchfT5uLwsoCge8NM8vUV8/s0jU7m21SBj4oe1F4JFk4UV/UQc
PAgHeiNEneM4YxyjP3QMBaR4pBPHzcz9YFGlbhxlQyTwBPYvtb98PD2a0u9tymKzzqYlEwOc5gDF
08POUtvOGPdkszhk6UifnCWt/sbbridleglJigolsUwMa0AMsL7+AJLmKG6mUv7ikv12g/EgUzKc
UKdFQgV+ROBZt5Av/Q6B8me3vNYOJd5XL1dJSxug4LzPwUqvLU2ZU/j/08hvxQUWCbW42KgUlG3D
VsJGZdjMIzTilgktC4GByg2jcRRENZI5RmEnhKN+4fV00xLq+t49Y6XviLlZ0j00d3f+/RhxPdMp
hlKEH+T7SC3vTYKda75MQmoe5TWN3GW5N1FpnGSdTSCdWFRRbhonObckKf7IhdiI79UPL+JzhBIJ
4msgh/RuFlGGb9IGbPg3hC56OukKke5iIwXAkCVBYtxgi+xfRv2WdWDV/n/hz5/YEZgKJtUDuA+j
MsZujPaZ//Li6n+hTtQ/ZJVMxuKNmpI+foKKOCu8TxgfENl5xixG6AijNYi9MbxjuSUgreek4d4Q
OsGaIwPjkcaikyBYNcOKFQ+oEWZnrhjfVH03YuE80DRAj9xCCt9rSYxASE2qwKSYsXmWscOSCysy
E8Ykhut9w0tTopCZ1PTfCOAZvYqrY65wWYdcwNAHNFaBMrPFJu49PAF+ep7coUSyCGaryjBSrkW7
0/dV13JHmdbU3avPhzqtPk+iATPfvuAmCqIMm9bqO0FEvfbY+QVzJFU37upNSnXcFyfEJAT6gZK9
c5r7MtB0basjL2+R9eit/visKE/WTO51fJcLg+BNYFmqQmzyD/Z/SxeefxRzflJY2ov/KMo30Vsd
Jla33Oe1EjWwsRxuP8hbn3pAqLkBEi4WLzSLvjG0s7QVKFMutqkibdOCOgbKEoTBGz6jpzrFPCdw
XSkL404KYjGMqSFGDlLLi7UnAS6OCJ1dOl3NUS/5ktJKc38/hVNtAOhks0XMyeYRLcDLzGqi227P
/d20bHnQjwOIUJV0G1bdYCiqxzGjNQ1pjzp+eKhWQwobceKVsaT78m/h8uuV4CsrACulAA/Jchon
OipGjWLx9PR0WV63v4wqcx0OIV4asp30MMIgt1vlZsuD9gdL43X9Y0E3F0rIVs206fR7B/7nQjb9
cmtnHR+FtilNBlJt81HrV2NZktkWNZtoFoylnCB1U1P6O9wWuL4DLnxzuowpvnsckhn4PFlUXLRt
x/Ricbb7PpgmRSBQrgLDaTqztY9O/tzRRI7Tm3kYzRHh1DshmFhaS2psmlgR9fIBgSYzpnYALurj
JX7RiCDrv9lEC9d2ON6iXTTPcWcqfg8iiyMRuexOUPF60rRQzV/F1IUPcsrm6anvs0T5K2T+1xOI
2Zxzb3l1Bko/bq4SY+ISmMJjNYi2P63Zm8E+4ayTxLV3XckelE0lkAN9DFFP/gKLpo/Dz2WE+c4t
6jIsmY/GtaqfL7+HaR0yU45LnojHuNPiIsW7YHEnWKqFocf7Ughk/7ktQlQYzynKssPHIP4AeY/g
6S6H2EcgEWr93GxdjkCdaOijfC5Cz6R2UZbFTDjJd0Stc9GXRDsEHKe9Y/d3jk9258SeFCDhXo/v
mA0wAX7vgV1GMPiqAVV4AzQQQyIEhP3VKj+qCaxEMnR8zzeJFTJvkaqc7PgsacUKdi/EzQcIvBnO
ynYnWE/yx461woQfXrxWjhB/vYisI9ppe/FytpxVKkcS21iPYB6w1zOhPivMJ3iMUlWwHXH9R13R
BEChKxU3xbVsZDXiW3kggVmy38IVIHaVa6fL6B5UYfcDecqiKVDzoJxxD1U4F/Bqn0yf2kKdTkqN
L7U7emO6ylu8E0ShCRefNqp0tF9H8UKWUVnVdPsKE+pwuMQ/pLjdMmzAMneJo5RInlxLhSOK/+8T
+HA32KeYjypWmqKzm9mO30JNxcN4K0FI3TR6V5Csg3Jt75P2666zwxxGDSY2FotYBIzo/5fk/ErZ
3GomiKPtYTe/75RTeKpb/K2lsLoRsUOvlkPXF5gF0CBXz7vpljeRzmvbsjpNLaBqbsQdcoukC/Pw
a6sZHfJGwJDSGf0hVMjvj3Cqb6naosK1jYspvk87cEnMevwdHJoha4bxcp5nHyJrxbtx8K+O4Oja
51IoaZfYo8FNaX234dSO0B/s/zGQ5SWN0/nJxs2G+yvgH9BTytt140s+MUWCDfktYjfk738CLjDc
bkPzO+8OdxyBv9mb0l1/O94SK/qLxzHRDGb+bVPc7ZAurOZUVl/OhTlXJe/Rx2VLNzRwk0Z32puU
OkbkbAaL8/JY5DP6M+ISV4JXEfGNHZudzYPChUV66hUQBReomrmYpOJ6COiSmpj2LDvMZZNQIOx8
j4NgFsXajKHnF4+27bseww8DNzBWIcIoOgU8uyo11jkhMXqnedCZv2mK0ELBd2Yu/DoIkWrbMdBh
h4oqL68zVXEcIwKgmShvA2QankUqev1jxdN4xXGw9IEOIIWmUl8yS9ixc4CZ6tB/O1NscisYUDB/
9EPIjVfZNjoQUQYs7A3Hi/C/kJeqVhBqlI0hMJtI5ve8YNhhu52xNO11txh25yt4aI0BnbDMvgEY
lQOp+htz910Cr5t2gaKEgrFw2MWgzn1p4ui7bxPw3J/QbTo7VELioCNwpQAZw61Lm9PmTFAi+uhB
CsqhcTmboy0aEY6R2XwLfwCGuHOMqMbqZUPnK4xMs1uLaARyLB3mAoXbIoq9agFoJjmxKz7emNaJ
py6KyG25j7wFs+zutQqjtrJtRBR1Z2brhSGLwrreLlWKx82735zvr45NvQZzYUULzEYDvAk3irPp
joUWrHmBGuTDyGoTXp/wipE5sNkjfPDLRmzNL8qvrejacI5or26pEFgVO9SCC07v8Zp14dOfTxu6
byHgGV0b88MhnPTgMZtFpGJ+GziRZEdUFW75HcgUzmPVliLGQ4LplImHwjVN4tCfbQZyfOv8sHeN
+BSWvpfVtbWwBHqzdsDH4i9BRsbiljuEbP4Wn9cWJtgsBdB7dUyIuwWjapGHTnlONVgiak1IMl4H
VQrun0iIvDurQ97HT9wnvm9VvYQTvAKag1kNK9Dgj11C0YkKtb7PEmC6fJALp8A7eMN/R2iHECS7
g4ETV7jEc2fEQAQu8igiTufwe9ModDvAL8Hp0jKmPekDkKRzcGvja7Hyln2obiXfWP3UWZPHcaNZ
+Q/YNQGl6+29pBpu3M2mzE1CT51fPIFZ9JBdm8cJkBgEthkYvE0aihNd7hqjpHh872E1X3zMlGnD
06BQsTSIrS/eWL0upEaceuQkXM2HxhT6sevdeDDfrfogpMBn1k1PY3bsPJcj/gZ9k67Pz64hTt2W
VVRQjHL90kjMautmjiS3XStmXpyBdJIg+5j2M7KZO0MuDeQbhTECbRIQpgC5D1gNG6Jb9BIv2bXt
B6dCigFMu+XsZcdb6QkV11jQIuPTZF5ymZEyoFzc3mReQ8pkXBFm+ThvIExwpkP4f226MXXktmkl
Iv5deM9fJpMGzvBitIjqWbSJHkvuDVlcXW5sAJ1vC0kdedcQUxDikY5aCLOtzhIxofHgS7SvltdE
wI8aKnt/Pkgfg8Rkf60M4Ewe7pIHWghuR9Mm/5C8ve+KAf/os/5R7Sr53AQUd4zHkYDW9cEquzWc
NFr+7u0X3pU9qPfZFypa76Rx6NBCCVKBlZ8zf5atbXGqi4Weu65H6CWA8BOcr/yWneHQD7nm8OeZ
14veLvW1kqHAj6Pl1DceQcFWR44aXinqNy/9B2rKCMiRVOvowoOH4yf1bQF6m4rLefCBJ5NcFK1L
j2sJKC82vS+Mv/F9xfglEZZilpVJZMr7UXylxpQOdMzU8/SF3Vd3v8pXUoRhxTFye7b9c9Z6Ljmi
UFZNpM0Bxlgr6metN5VS7c7d24Fs8zl1mejgN21U0v0lkC1WVFWPIduzG052FCosbU4vyLRnys9r
H9Sb/hidSiN9LzC/cfOGwl0/9K61Y67Q+xwUPsJ6mJrM67cyCgR/FtsFagcrHfKkwQNudeOVuFwr
9IGBFKZXNrNUuWoOEDmHKSRfyZ03tfWF1PKS7XtvUT3uPdHG/eGfAFgknzLTkFXPeNnkaH4/kjm0
7RnrjrL3tcTvUiJYGLUx+DvAsXN8+7N7lb5uQUyG3JsVWSASLRmLk4LN3WUh7XseH3SPX60mWtoK
dUEQEp2zKQRjTNZjqxEksKoml60HBvoRxRE8XOawBrom3otv16/inJ79g5ZvB/p7K+utj/KyZcZ6
3vNUWQQcNGuMZQMqFPtoVnl7rnQ5xX8xeUn8z4SwcXhGCOCQGN4NWyp/pJG9higN0azvIUDDxgp8
xSXqhT6zw8lh9UXWsXcKLNg4feNTTC0izS/yHFGq5HWQfw9HycaB9tfW5qLCllEOPGp8Myi2dnIS
AtwgA/lEch89Bo59FdFncW+9FJOqH1n2AxgQHtOgDip6IZXnGs7AlyH0SboSfm+L501x1A67Ipq9
4hn7rp76aJVfgQ8gxAnf2CDpVTAzz83ZSyKDUdxDgTVNAOfefk3AOc9PTucO9J6CuU8Q9hVXU7PC
0UJO3/BLEH2lsLjkbJcmW1r4us0RwSEFh2yppykXvhWNansylk7iAR11IEcIjrWZ2H2JPpToAwSN
0bn5Af9J7yLFzxcoBVByAcIBYiFQ+6+GqylTATqX72B9OsN2HXj+K4PCUZsdu3Q7EmY6bXoNzAOT
Mhgicmmuwww2fqCI7NIIzBeJ4Ids7zNP6XKFBKA3b35VRxUltHKD3mjIIiR7WAaJBvKcvUwd451e
8qNnPxvKCiAuA+BVdWaFuQcBwdPGPEXY4z7cK4IpeKbTYY/p4/o4eUegeZ5zKXnVunYDAqh6DLLT
2MRw8m1UXOtvchmRvM51FpHR7DzjbCPyQJQoEqZzXRmBjMR4wFSno0synvIKoJzYW6Vh/v9awYNb
bZNQGfnp0hktEWTIzLlVAUPu51HF7CAM6SZZtViVSMU/D8BqbzjUPPJrN6PswPtg74AmV0Quf79w
Ct2CaIyIElMwN4Srmiw9lhVkfq/kskxZ75/P0mRY4YeGkN7XZ4zabN4w8HfU9PD3SHmPXEsOXotM
z581CLnTxAdvBdW17ZlIkB1zrvi+cuaoqDSdamSfbaPjt6TZPuMj5TabC0W1rBbuF5+T1fTDPDBG
ExUyn71xX7HXD8gfTNhA8y/pLuVc74XUuwpFkUsjyL4b47HwvL2G8UTNdGAq/F48LHxcGVjDpgxz
cvAQG0cz0keiYoojg91ompra+joGf0pitUJZl8E70JlQULPNfKqlsczB14Im+lm40cIavAR0q3O6
WVf7kO6OVeiziY+QKK3wS3qlgLirMFZc5Mkrnihge/o+KjqTW/517dswWamO/8l7wH9KqMfUV2a6
1DRt0Q/+U6IXQpZVudn40xYUlwntj7xiznazNtE8uCBrNX2Ko14u4804eeCgHD7C3HJVr0UvrMj2
dLO3pEtMG6fKAm8pVhvlOb2jyea7MUMt3fOrM2YFr+v3vZj60fVXNzxwxc801VqDR+O8dONwoqGu
vNevdI6WhzJyjOOEcoKDqOLYTVHR0//+NBRGBYly6h2Dy+fmNdwtPwo07YkN0G+goCXSE8t0WadI
/hSTfNG5O1wZrxM1K8Is3166fSn5W50ksEjqwfizl52pE8Rj007To4LxfQeKjyBbX1iiY3zILOVh
eWDR9q0lbI/aDrIH8p4rTAnRhWwMfJDjL4VRyGbBxlddvnwtLsHwo8NADYLUWFNxnDVy64iv9mWO
kj8qlUIe89GfSNotZNCGJALiINTA+dumPtgtXmAsc7b5Sm2GvhGCp2r/vvCyttlg8WofE+KNi40z
bhTJzZcfSFpPBv5PNQp89z86RbvF08L0wp+JDwmu6qbecyZCHRc9w9K0KWmzIq18NNIm1RELXjaE
qluJ6Zzfx1qBlib4bN3FZEVyXGvw8EP3RGf6wAJK9Ngq10awIM6rSn2rOtDixtcLoR5nSmlkvrFt
/o3F/p8YoclEqqoM+qTe16vPWpxyKchyRCUvj1+m6oVL/AvZA3vh0hzb+Nuv+e5ISyE5vZxDh59r
zAGGOh4/mWw92RL3g/yBxnxZGdy3R2kZbqedLk2yuT475IgsyfMRKowm1OhME8/L1X+zwsl/FCW8
0xZuSWrbfrtEHnPkHHPbyCaCxdIViljL0jXA/Vi3BTCwx/Ki5NLCLDjSXXPoLoyyJ8ueHcWkpwC3
DUSMn72xC1X4vQkmNf9XONMWevtaCoAGUos+0hhvWZkStxviw+KEjOtzWtn7JMZOCRs6hWhFuhel
3PpMVsK3mjl3ys5MqedKDVG3jzWvbsmYATUQk13L44QihO4USHvJSh8NFD0qgmezNBIL5M3tB7Ti
ZxsF7vL55BnQV4gs/zr2QVJv52m9wZDc7mZFp615fAmgKZ0/bTKFYVtic3nsrqdfTodYQKifm+PT
b385wMZc2WXxoDzqr034pJwq5e4r9JpAA7p0FiYFXR+nBXJG6w5s/UDgPC6hJCheIDyFn4FSjbvD
/GQFcaEb80lTGsx2EdGM2tDE8k6Wqpd1zk7E1piPZJU50nVSSmq6LvF6Cx4UJKmfKSdi/9MeepeK
qGotONAowciqeqGe7ya0aILpbM9DSDZgFY8XiquDtHSxYPnrp7JXkd2XRUlqj4M/L3oCkXd+pSbW
SvxT/2/L21jIV1n/ztlYCxq63OTdQvvWAtrZnEg451JAh0LHlw+MFw8FKwpAqYC91wHhLJ7vzTG5
OLlbS8IcaCGjH5xCiwgpthv2jRrv7UWCV0Quas2rdyba5K/KKD6QeK6VkrRe5gKmygtMxRazt73U
5q11mwwlnPQqVMer6YH6xUUYJ3ItHnGPSGlD/Z2P/l0G4k3LrXkX0LSAAsDG56L/wHNvt0yhVuWQ
WwJeLbb1/LHera3NRlzZBhae0f0amk23aT8R2k6WmK3C5hHn9tv+whfgaah6uyPzc31TTx5f6IQ8
igUfeNwZjdF9dreciIQ7Izgtv/azRh3OrmOqVYOfLh5Thj/jhYej8lN4wX6VSQPv6D1Eqkz5YT1E
Qwi77BUexb0FN789JG87D8vDDQaeOjYt0+UZW3GMcLvedC6gl0X799DbITQwu2FMZSq0DFT9uwwZ
jDgnYYC/yyUTPOPxA7KZQAhK8G68l4/CNrTcMX53+E7Ok4Tbz99L1vXAnLkP8ZmDckP3vJv773ev
Ykgj384bftKT68A9aPm5J/L6EsMEobQxJyaTwkpoNKOWMEc69hsfH73bliEAfC411Tu5evhJwCbq
gTouPa9glXGtTUjnNzUZMP4bvQ31CtZ5MZdo4NWjPHPOQ/2FOIAb0RPEcaa/a5LhzSaZBvr8ONBd
gN3pgmq7/g4cuOj6alvoJcXn8IDv4dd6ugvc8I5rH411+LJqGq5SX8RlT670H2PRIQXpJz3PcTX1
hmFuNbl/GeCL0Q5mV2G8SLg5ibFpreF1sCm68sTD+d61UNpHCaUXT/D7FRNGebAntEL4f1nFGE9p
S+ks0Mdj7mpPYa/817GI+pyqwWUB36GhVO7rBTGvhdPfGdhgWu3NNlqFgNCefd0LXCCEALaHon7i
rVPSCJ9yVy/JXJatFR2+zsUi8fyQTA/Un8Hugrp6Oyejwyu40/ppl/UL+4KJgtcAaLCeKxp4FsPM
8geiU0CqAVMx2BTgnSdCZaGuP7wmBkakSHw8LMuIsd/0N3aJq7/5/MWrKtejWfHh27iMlkMjfmRf
WsKGjP2QxHkcdiBdKxsjPCdcjBrf1ji2awCekC3NCC3cXQx4u/dKmWLbymHilmhCnDBLM5aWQuLm
rH6zH1/s0q/V8HZDp7V8RAYeidXi9K6GQLdn+PeU96J8bbnCw6SdGlKj/uThOhXcrIvFUkQqW9hU
kbpgwM4ZeABktF5F6EO43zPpM7OcLk5JKFBOS57xlaQiBj0KKVOiazFxrKwVqqf4tMMsAkIcBdCt
nVRiWBiqYdQsCYm76KHeorg5mEsV/k3o2/7wrmcbv2sLdluGdG7Nidgjr7AVz4PTWgQWaJngww+q
MHQTDwx0HFJ4CWjVw9s0rzxL3PsEs62oxPseSr7xAYJ9ZlrZGd3pSi+S2U+FEvFvJyFf1T71Bb0r
7RRqf/CUvP6TVEJssrcxhdc7r7EYcdDn4aFQjg4JOcjiYJaaECmv7tq2tbR7pF2NbXIAT4K7oeyw
B1CLTV7sgeqpnqVyHpFUCUQx+75vVwnRQhVjfMcyi5y/hk7lNei0E4TCJwQLYTHJVacjkUOpxhz2
jDWSSxLcRXtNqFopChUZCsOIV6NtheK5pB2B5vNzvJxjLgtj4IvCKhLcxW2fThVrJbYCq0XMxuN2
Rd0zPBJUvMYBQr7xZ2zTjIpzK/bAmKejUpPV1JJNwn0dTIg6TVr6Q+RTiv85TE978donZXm/nRrz
AkMEa5DhlbHaCgKpN4TlKA7um24qQOSeS3Qj1OEBfL0n2PVAJxIV8G42We+PQKaL3JNSrn3imSa5
zgIUv6rFHqWwbxGuhtj1l3Hkze/k6iWBz4XwaaewiYX5YSQT9egN5ChJOi0G+YWHFx/XtQHi/L0/
eUkeeNSDnTkGPxAIAIgbWWAlCzYinvKG6Y/OoM3Vvcy9j1KmsPfsGlGfwLyP/Fuixw/cjyfw8cw4
eV4DEtnfNj+naoX2aKuI0e1+OH7xiDLhkN7Kqtnz5SRrhIBI3jMMxDX/eUd+D4MZaIJ7x/91KJig
9l6DMDF49ePlMk7nOuJkeyjOmW2a3yaDrO9T4uCNM7sxjk8/Je72kdgR6hYZp3BNtTkdn6qhnsIR
j4yhhqBCfCZGaGwDWg2Lsh3cyUSp5HLz26h93pTl2kTsh8WN7HCXk2QHjfADExA/H0WU9fZf9aFa
MohpdTTEriNNyNMhKeq2P/PXW9n+IUKVqIIsOWU+Wz1pw6zFbHKvpis9BmFpMyCdxwncXL2lu4SM
050GRFtTstSb+IoUtxrGCqzzFZ7pe40ezX36DExQqeIZHrhzFUkdQDW2pkqFyjKwkEKIkmkCsABZ
TwFOrJkAaS1A6IeGoi/6ulgoK7Z29hpb/BMxIfiNsWG19ksRDoF/vbG/PtS+mY7dmefWibCxDPas
WMqRC/gXr7Mb0j8VrPeCOLAKdifeIC+hT6URguwowZgXTsGVF2cLRZY72FuuBjaQboOfMRNvwyak
tdqKEgA6vWAUKpOh1gSvocUqMF/E2fUnGcLN76XiOerHsSuRUP9K2b1BtBi2dX2Lb+x19x11evs7
bVtIsDINKYUr6fSinSurUNJPLXQJX1oYfHXpiHbthbylEAau8XR437QBwwKx8HCDVFdj4MdnEtpW
tvzP++zXd2HYlu9hTBQeRqmpsBzElDi/2OQ4Mlu23xkCx93QaJyVh+KPNOcF19KK2DI7lKi/S/nc
g4JFL4k8uAaY0nT/40dJ1G75Y0+fC4UzlN6T5viOGDWSc4zHX629MJt6JpltOW5UCqNoyTJZvJQo
4ng6erJ/6aeZSKe0Mdfi3BexrDgWzx+uEXVHfle/uxGqD/1e5VeVXLLhcpJN2Pk073VLufXsSJBM
ArOI9r3aHFMyA7RXBhGgLP63RhwAcl1ry7fbSyvl6l4hFccRr+PFo6qrbbpdUfbfgQEcnA3Y/Q6n
D5jeUPDcV73AekSwyCcwSgpaAcXQAAlERBUpuuylc7PxMYSd2BZ87N0k+f3V0bNQ16wIXUvvBH52
xTN0HPHtS9U8cxS8MqqDcZb1VMmyT2Kd3Nmidbq/XCIoUskFPaKkiLFkCM+IF26LA7GMgpnp1e8f
rMTFRZOcqcxjDpyiBU6vY0sSsliJar824+FktEa/7CgZ5DiqILOtrnCGvcP3bmaJDyt6KJ7ZDed2
Un4+u39bgLElTnmkT56x2NLrcrn11fZ1xk6CswzSL9/rgSMNaTBmSsz7XOGNJ+b1Yg/h/1fxMJBy
zPBE5+UL07B04orYX/eZyd3bZYR988wYTBMLsjySVW5JC+LEyEr4lGn4FT2BVwBPYeUKdUtXwaPE
WsRyVUx1hUZeML+2EODlYnTXNlKSwANJYQmpA2noqwg3BZCMceMU15VQNQAgh2W/pRYNq0s1oi9A
wenBNZu3xXu8j4Xjrhh2jbCQ6wK6Zpvtc2o66yKt49DtXOdfzNK1lBGM9C3e/64+xc4AabwAfBhV
Zy3Gm1n3ACKu5CttPtT6bqM3xO2wezKnT6R2gYP+jsFc/dqqcocqlmFv/oeN877SsQ897ivWJVmF
rxc4gKYb/JhH4BzmaoI07rAFpDHJ7KRB7m7Qulj/hAUxPWX/yK8pwcITJw5BatzfSHJmaIXr6fnY
HNls2uuiKhxggKJZt94I9D5VY9XN3SuKndwFVwTpT/qJqpddRNYBSlvU5M9l4M8fQpLsRg9fIrHZ
Ch1X0mx91cy+eq9GUxCJeNWCo4Xul71uVOdT1TBMRpUsEY1/0d9RUZF+qDh9CZGqQJg3onSizVrU
wm0IpQiyTW0Jw9CdjlA9dZFdQJqSgXSEOHFdDHWswAc3N7bYQLY8MfNzBZIb1iKmp+NA4kGQj4fj
Ym4yrruy3jTLTJETeo4iK1yAgOXDFHwtbcaq5i+3Ox3buGCLC8lmftvZW4hM6x55Cx/a7wqZRmQZ
ybVuwb+bxaP99mMvhOfeETK6KA5epRubjdM7zUXy/8oi6XXslofGy5Yf0gWy9p/7fBdxeMpGAmsf
6W4ndOeBRNNDBBURhDk2ppL0LaXkrnMT/AaFPrZCqL224TUGqLZ7OrbMFfxz39ySBmDwesvInfyu
UOG+uWRQbTJMsEp1DsTeDFb+ZIb2GaQ5+t1h7XcCE4qK0xA+eGQ/DS9cb+D5KnPqgKtMeViW76Fo
gqewCDuAIfCbTy5oT+j99/ooYO1i51eatggIIbErYXzd81sI5ZgtwrjWwbGfFLUwYhzOj2V8BxOn
i2NfAPXmEr9wKjjXF4D5BrtjyyOd4rAOLYccUHjtatvNDeGPn3JANVulfrx/dXJEP7BC7DujXcBW
lFrlNRJ0jkGxMAOebJBhxHx1Ql4qIr1hZbCQh3UKKHpQRwFoICttPtpo8SEo6W/a/nlMmrJnzHoT
NY+8XBpJuDtsoedBHebkM+8Gg3nNyT0SRLOb8K28eoPDAhQCDr/ON0FmnkBgrfLIS89eOxb8rMHP
H64b1fnZQapTQoofcC7W6oR2iV2glkPw71wofpxRUZwlCNx8MLU18aShtzqXWuZ9XbhKLMyj56W2
8fva0oeGHPfuF7a1bcx+2TRbfBl4rZr61RD609nQ5AZ1jDcuf+nODst81ZibD2gEUFqZfmYQvY8f
XcRfCQ4/sq1oPKPZ4A0W7LBaI/HGzlpTG2c9EERc9/9PpOPhx+mPa9m2GvKyXuAZ2GYrpTgG0HxY
oFuFRsSeWSQ3sxqPHUrVFi+PteQNbqyXhl0SKH6f56X3irfiGVgSG7Ps7NlOOEwZESOV/DNjXu6T
sg7AxVjQASieOH3urg3fs1d23bXzlIm3xzU0H6TvpnRDrmAHmcrZJZCdp7OnnLPHHxFvU49ZOTLe
vtavucRUPZQv5Q2x1sxlnoxlBGwp0oT8Q/cVXGxAps02pTZ1ZFNA+i9IkFDIZJMH1cxeT8WKUUY8
3OQ6LVoE5YcwC4hBbqCiBrp51UWg78Etz6x/o22DGJUGe86BOxGJ1OWpi0I//a3UDbntKjzoeb2G
wmTH15QHbaoiMaN0b/+bgDQaIzyR4RYY3WSXT+WIeeyk0xKGHJMn3lzqCRwOXsd5M/+aYBSyW5sf
Sa/lpD2CF9mWnN4hqefSGxhAVPEJ+k+jOTL7WhPuBvcf1RDwI2fhChwYJMTDbgs8PiXNSX/z5isL
KS2Sfl+QxYMZs6+zJDRMneaVRzkUXVsGXjjM6AUWfPPIxlT4SBUF3V4uGCtej9dfbQugqGvsNC/L
fYAEuiy+k7Uckwz/o+hNnfZXmtLbVVAaPhPIHNypbXvJO88AI5pBVv3hCW7HYoNhuB291OqpjoJD
xjKc7cr3TggINJD/vLWp9KBkpf+cvwg7pTZS2IVe5HgQ2cy6cNVR4Ap88pHxQo2TOvrfadqTeas0
aeVcX0NYofFtzVdqcSMUVPgbMzAF+PpRZuHbBt7C+7uhCNd5M+NIxegVslVKrR/HF/wW20YLCxik
yoOuFSLyK8E03nvA5ywgWsi651v07hXpIVEhitpGJOUVN7f8+HBXSyP8W+ztyrj627OWC968HYO/
JrWoILDc8KrjGFBVChrHHXC/qkNvuK0aftL7kOzcaGUkTfFgu6B2lkQDYaG9FOnscH9f+w77YO4C
9P3EagqxTTHrzgP1F5MZhFll6t4ZZn1NZjn6WBpeK8JZjo8V6NH4DJEAxk+noTACfsd2m58ZpYR2
Ior/njaLDR0k0yU4++Wya7QuQCK4bgkkceCDQuvHknmF7tNY88EJF9+9qfSLLvPc8UDsSkspBsLr
otpjK8e5oHOvjZVa2fzh714ybBsI/xa64XiucUFmBRK+xxIAtOS8JMJcqu/e0noU4tgo7DNwGzXP
Kj3VFWnWLAd33tbotGsq5qXFKrR6fZbqH/0EjfdRoyY3MhKM3ZcjEn5NjAcJTfr6NysnbTUObb0c
8EiFP28kfr1F7FWkx/hsSiy71MFxZesse4TUCoz6lQvVUrDnYMVLNcFBZ3yKCkkHdRwzr2tCQdQo
ynvO4W5yWLBeSOBVNup7UFnKsKmHnLI3jhbtd+/YE+CPtabqI4on5nyUSsbBY4NYLmSFlB8fBcO1
ubAPBXndtk46sYB0UHSNcO/Y5kG1s5JvyWbEYMfZxk/2eNaES4SPuky2P8kvaiO/YoG1QbmNmqmo
tChOue93/bBRXMDyBDS+pg3Yo6Ayvh5TPwfuntBee7+c/gR/eJV0p3EZP/d2dGCAiIzeKE2x2XTk
s8uYiLCMCoJdd7Stb6Y3WCmrqQqJz1/wGa88o3pisaPRPYBrD3Vm3emCgLyoK8/IwOYt+ul68yX6
5TaqVJXvGZLB2c5rLKSzmo1tIoEvILCa+tJ0J6e4vfNHEtkpg8/nB06cw1FZ3hvV6s2aBJiTlqZ6
WimhtYN9ofrIydVSUplNoqyAfVZb303MbhYuFw2EWfyKGZ7M8i07K0n8Na8F+Dg9mSpLeDq+4Rxl
0OU79gQFY3nIC+0CaTBUOSpaQDqeJaKUkcoY6b3P8lMAShmdbWQBjUeKTfM6C7jmKiQLTlATQ78Z
8ukacOh67kVL2QiTdO/knrMNv/LEJLGWVgExgnZk4xDWZ++FjTEbotxP/WTSH3gOyWi83NGxl/ue
WZjeEgg+03EWFPsC9LpJAj6HsET6b9EF9oO/92t0uHyEXJR1QrLJd+TqbjlfRHzfA/W2bNuI+vtE
yKvfC1rMZiyRDzNHgUOYDdm12jqxsnXqzqC5bZest1IsatKY6Fuf/Huh0LeLKJdYdBPyRlrsrQbV
qJ+VFHxQG2Az4JjywuhQnkumwtPUmJEmJSoQfUBjY1oXTe4ZecWzVnEWbgi32aw9WkfN8OsuHTVb
WVdkY+NB0/yGaUjqxAXMpIIHrTIPb0Px2USfDVrqm7L5gYCJvuS+kLjynbBcs+9pzCzk5nfv9snO
XbWaYgZw5K+xeXsFaEPxiJunODxo9HjoVUtWprb5UCqa35m+oyvk9+DiKWo7tRYknPzY2OoihSeC
xmE6vsvS6UFdPchbooa7ZeTnbdIHHHxEZrndaWQhFf9KzN9doCRDbOJdbFvoHiB4utsOdj1hCW0B
7cm92SWuv69K3VkOmE5fm3GeiJY4VikO8g3I8FTVdBg0fgw1wEnXhaKriDxbyxRIC64n30d3S9PH
CDtnpTb4KyF36dbtUdF0pJiPoO/zDKGZZ2LGdkISWer3bv3UubBaOG0RnIf+PFaj0LIROPc/UVkh
d8vKdDYLuxz5Y7l6ZWOEbiZ3GWpnJ7xB1y5waO4tUGthaTmhRPGtpEgzH4Vfyd1TA0C8ujluK6Lm
bpB8XDGekAU/j13mzcVCq1BmX8KbrsABjJ3nWz4XixL9RFUOwLsEohiK1Q17DI7vdzNW2bxKgvMp
u7Pdm5dxLk+aXciFML2770NIIcXieHgJyLn/+F6fByX/h1Ru8QxCN9NkwQrWgMaUrfzC3LSGiPDW
cjowA3IlSh6XMsz92jcNpVyfD3yjAgIBcly0K7Ji2k04eOyY0YSmqrf+AM9G4TS4T7k2/eMl8IrG
TI5kZr72hh6vkx4d3oM26AqjZD2vkvS0PAh4kRsxpJvLupgfCJ+Mw38jMsJJ2IXpKmbBQaEj2O0t
eAvTRrHnH5QkNkTQW35TfbybniF6D3yiV5lGKGi7YgcHJsTwI2QsVHsUD3NlkbUEMeMa99kIDNcm
OAi1ciSz8dz6/r27rPFXOsCUf6a09FbS7CnYGX+gn6G6r2az9jOprk+jmWaVAHbzle+CTm/PFOLd
k0DcyLyy5XXCz7ap1izdU+Mt8mvYGgvmrcxS9yEQCEZN/jdb5igXGHURgusK5frlIydpZn//VWgO
ZWzL0j4vMu+jypklbWE6bRCXgjZComBNv0Y6tMo948LO6Vha/Iyb3grWR0ZYiu1wCx92HY59JfYg
i4CLQAS1OZqdAD20B1ICkwuZhLAxUZMWrznFvmr1YaNfQPmzFk6VY4g0EVfxkreT1NMNvxY46o4H
2t6zTGgUTOhkSuDdwtBUXPnhCRf2vD/LIaiJ7BueelyxUHRuXhJYX6kpUM9x0QyZETjHl4ZUhMKe
BOXPH8Z6wfjqsYxBg5fzauWznosJXSd8R8j2iMC4yXRhumgt2t2gTMAQAUSKU/1EBMxDDzOJdmeV
MD97rxeWIcojgHYoUviVFpxZnVqJ/raYaVCfZGqlD/n9SKnR2FobwjCNbRwYgy3cxVZDTnozyuVg
I6kShYnultbxre7Rh5sEBDaB81I20C3LAONxQ7BaX7cjYOL5vQmKVOyj/kX7c/BNjhioUfH2Z+Jj
hjVQgOggzfOxSFBwPzHD2szR0fG8BlUwCEiR+myfCYU/bndqZ1p+X7LD/21XTG8byNd2cEhG+XH4
CY7sp+4MMFXSfLzyv39NtjxyVOd1ZWoP6ub3Oz549maoEBlM/puVlALSuJoCW6pWLZVwBw66AMKe
DZCNssna6m8gNsZwQaP3LkrRVTdvcZP2W+nS56z62zWScKusOo46NJNrVLO55LEzg+FAk2ddlmhc
nKwlaoX8aITSNRiCpO4C8Lf/QwIisRZj36AGspmocbvuALSslt5vYOZJP0RuzBWUkjxq0+krOZ/G
6yMjnltuLaCMTg4S8nqEMvdvS5pptla6snWmtYsNNVrnoXYugFZe6attZvETSNYdwS7POyNUwFy9
6x0Q7usMrwcSNnTWGJghqfiaZBQP+D/ohySxMo2GAQ+IyhmJZNluzs0oki6BXJqkuBJPKs8WxA92
zW3Otbnp9ua80moxzB/wfuHUlUC1ArGsw83skmyOA7jF5vIiJoDrApn/Cws+6fdjvuyjgz3cx750
ZQyMfLY77+E+J0F+U5//DnuEKova/R0RkoJAfmiLS3sz+kMnCkBPn6SUgnl58TAEa5wPZ/L22aty
DYc0MWmSSYkM75UCRugAvoyDrBDgCLRyi26Uy3mUzWMQBFjCiCORzH30KtYBkDwo8TLzK23QfUsU
WhZJGbMYKpB8gBy2SRHcGHPfPGg/EipAKe0TyPxjWeFOOdq2Ks6W3f45USCenpIt+p3ofr7euC5M
GXdzQK+XKMBP2cTutQLFUrhRToSXSrYGjaAsyiPwN1n46780pCqnXK8Q+cFdlGbN3bVEeCg7yEr3
wk2iNoS9CBSLF3GKhPUwIbgrCxCJokGGPVsXwdvqBM26f/OQBcseOUwsZlathikkdoxQP9oFjdUT
BVrXIIjBxZNZSssxp7lAzDgpo1XFjtyXVLLkMStdSI/vfRgfEfE3ZS4VcrUQkfjd8BcOBHhSBWtK
GGPCG4HTmcVISOdMbK8Hk6zkXuY2q8LxRBrNPCb9vfnxomXFjDpsnnfZOajk84x0i1WKx8NdF1vu
XKDZ+PYXKudcoWxcS/pPxuWSbYlEwOtXNNZQvlCb/O5fdVr4its9xs4wnnsci1qquQZqMHohLnlX
Y/K0S7qOWfXtHPdiQMljsONKr5tdrYkpGFA1afuzFuZA24cA5ISVBduVb5fcX4xkuDkFxp/lVP/0
4Pp8ocE0Xv/Sd0f+OV3C7j7/cYA5OlWeiB9cKsP0oDuUv2XvmJdp1WZvdUIJZFGc5DMqyzd7Z9Vh
FxOzUu8wWs8P/ND+F27ditetOorvb34FXTjXl2ApRZHJ/VybYUrxN4KVMEAtvUkoYJkU9QlEd2lh
zUMV7mSF1c8XWmrDUq3zzub7DROqyF57SDPNNxD12X9wGp3RT+S1i1RAk9Btds6/O/yHVJv9b9Dl
5f7Qg8bqv++CaL6rVaLz6uiYaVjAK8psFPDjRozhiYcnPEZIZUSER85lwPWH4fYrjnKqErN6bb+y
DpU3RLrLcSqUNzrpMbWy53QGiyXw1s5MqGh6iuPJbi5y4sk13WXwQN/dNcesEsLwsRT/mBK0lM25
EAI3PNVDutT9OIVj4BwodiW+Sryf5f9JD0FuKQdkAkvq0L8T+ifSA/RdARyfrsOw997P2uSn/Sx6
bPJ748oQeSKyAiEmfAtabSL751jza5w+YfueJ2eSzT9TeL0hUmqhJvbcBpe+UjWp+C8ajwODykhM
r0Df4jD5wENuaaK2/MnToTZONzO7AdPtAR3FsYSCul3T2rlFBAzxXkZj0v2TmJQb5rzlsr43h/nh
yioow9U4Zv3sWqIzGjDgr0Du1VMyYZB3hjgU1F/ebGMbNrFJk+2VTNgE5qc9GCNkRUW1EyNfBzRs
FS4eRf3L6QXC8GOuDLkL3biZog5WkqwCsbZoKVB0WqSo0Q18f+nmpiN1QbO+syp4hOVQvcv36ZCJ
nQIuQVNQpZflkefsexVk+a1BRXEdyBsQntAEKrYvTYBU6lbbsr1WU8wGIeSRRLXefaZsAjobXcdY
iJ+fT9qQ/H2/Dc/KnQ16nIAjLCi8uQsWomIWDurOZqaNurAy4mDrafjytVy6s+bOmG+ZledCYu4w
RHz/6uZP6WZF75n4+A1FHWV9rxkkrAkBVC4q2TC/cJQTFNTwzZU1pEh6UkKkWo+ZT0draBLgnIpg
ZxQdf1Yg9otphoAYIRAmilTY1NImacA+Hg+VvAlvMJ65Yff2CE2wuTTYoo99hMK5g8KQHzh8vUJo
EqUiFxpEs53lp4O7GyTBO4BDFKFclPFnJ4+PsD152VgYPD7yAkPTEoBGx8TCyNPrcFFoVTqcZkR4
iY2mNAVkuUyaQuszLGL0ewfKGgCAcnZumf+JnwMumVE1VQeCZpiio2sGvS2lR3VfINM9aS8eqj/c
89xXu3bqqEWGlrHi9Lj7rpgWXN61+Tody79fUfo1S3E9uYa/aHnq/gJeb1zg5Xfe8FSGO29rrkFw
1Iyv2Es680J0eRbyqbrs7zwno2ItgrGiBk0axpq+HRGWm+/+FTsmBLUjVzJeqnNPid7l/+C37pFi
W7lSfdWnnlq81GmCaW8bliEqc0YxnKeVxWm5tvYGEIYaizU9uxLXIUwR4FIr9VdiwOj0RSM1cCzS
ZJsLue3JYrWWj6JQYpPG+/7jabDYrESpE7wqmw/cwnNNfWKqZ+s3+x5rDBYq+LnsJW2fBnI2Z5Yv
Wo5775IeJi/VFuA9SxIBECTvDRM6oXxl+bDvoFqLnIWLyocJMNjbS0n63r0Wx1cgcO5vGxcmTGad
O99iwGou1O+20SydllVPIzU2blQAfL/1urVWw9GCmxA4OzTH8J4Pe3rne34ASn4equm2k1SrkvWc
0x5c5+1PAwtTqiC94MtapcDa/bhX1HmYz66gVTOdOhqTpVR7c+bBQEKfMM0McRq1T43dzP7TcWmA
4CPHwPYB7e4+sLsmky6y8w8ZA2sCLeJre3p55v+MAGiitIqbfSjvlS2BoEU+1nJ0RMYFxxk0te8F
mDJGbtRULSLdRewGpK+kMyzf4SDiy0MkOAQQqM+r90UkRiC4ekTsJjVqI+cLLBM3uv55MrfxvHJZ
rZ3nlJR5qbCw8e82w9kd8eQ9HbqJEGvuFbZtPhXKbpWWb7Sgpsbo1pgKi2xgv4+qS3J4nB4azGmp
oDuyo/h+eOS/dRsp6/HBJUT9C18VPTzhkTLWwD9m2GAgxdTTxmd6q8pObv4Df+O65B7KzhX0xIZw
KBo+h2Cf8jaKFMFk3VEuJ+1wmO4D+VQf3zGiMcnGXwSw4FLJFmKvRZpxcEslT98B8q37zwy9V9Zr
ZoO4dP/p5HPQCYds8kuxIPRu522YVIwmNVxkzzAMjcUfgOjx0PH1mR1wYFiWWRa0Qc0vSnwroSxv
sGRCOrX35iPbOQQ5MYtcBDWrrcVc7Yhi4+1A1KfYZKH1qKj/6wYJhLVVn89E84JwPcovBw23Lzml
xnH9WAnFKjIak2gbe9b7As8rJAel3Sdg4jL6YTmKW6YJLD0ui4ERF3MS2GVQNtT2nEFzw/WwfIjZ
iA5u5Sshvr8OHih2a4TqLVev58b3PaY3wSNdsNGqvZgBaW/0NyJNxFhGfg5Xe94F7ZrMvD/WV+FD
ZZ/T/DTxt45CEeSDZfcveitY4pyV78AjnFlDjVcT4ueAXiv32NPcUlIQskSX7tIrKXLNLh5rM7mt
kENR3Hyh4Yvo1nMk3tqY2T+nqT6nN25F+eUNPw4WVjrHjSfEHsXtIOzHX0fwE1QCzlJPNJXYYyeE
xkQEgxe7I51EaMwIQIECqQJ2LCXvkYkqG7AShvSmEwjgtQgB0FyiLEYeq3GJTJLuZNR4NNFtym03
ppjvRrzKzJvTRR2z6h24/m0o3j5dauhPsWbbb+UwSct/SflOco4Vq168VDWSFpaEqlBfL24dMZMM
1y3yHzpGjG18+RT/85qMS/pc11xm15N2LsLmnKiDPqwjZ7i5PvvD/KXqXXoEUW1n1deW7wgjLpG9
I1soIcDacO3rQfFphuigJXCkS1vJB9Q5FThFGamMBBLC3EoZsmHvIYKWzqpbM9siotuzZb0ETPlQ
EffHlHbODHrppuAaWdI9qkASnn34oclk42Cc9hPzLQOkKHRrXtCL8+DSq/6iu8ldj4vwJmPKA5bJ
Ev8IkwHABSQjg02iDCjqxIwwzHnE/m2XwsS+xM+0f2VP/vRuwFOAmM7tLGKiDetcSE1el+1rrCtI
5KxWSUAa/yzZhFL77Pl8rhKHmt1WuF4XmdollV791TvItRQr90adyjQe4fxwU1HOQ21ZOUzTNvXQ
tE6i4Ftqj3BOlfuCnFBrYm0Qrgdfdt30E2xelwKIkLUUhS0MrTInSLt3mIJRx4mhONUULsCL40Wa
uQhuoYLYM5MOcjWc630xq8Tvft8SNeC3otqv15V23V1OkSrS9m6NKQRyKPpHdQtjbqmNgChaPtVJ
lUEPKPN4rWfUdgik5N6SDLJ2JpG3tU685CCZNt7D+iuzOeVdiOEJ6Ndh8aqL6buKp2ysr8FF3osn
WLe/pEXAQ2wrQd7eeKTdywWQ1owwLzGTGfs2saIZZzZXIi5QHXsGEVd40H/62iP9JLCb4Yf3TnJu
hiy2y3wvKQQgPHDEsj8MND9aIta2Oma9zm4ndm3ndHPVbNygcTdMRaPQqIXSYEAKe6xP5nqRl3Wx
Y35OJGtXbat9Ks8wv1zuItyrNBdUaQKuUj/vsHXNtsQvuRHU6Wi9/IWmtsXWrtyA4j3C3cNmGRTM
yc5u50TCN7oPZ7oC3X9AuOuSDJQv+IDn1mVi3o+1dyXlpRR+M1FwqBDEA4+kawdDiA0lch6v0kre
edoQqtFelQLtOv0WJoi7/K4xEak0/OFyDhMO63LwoPpdBjSZ6oNN8wjA3c0JPZBmmluJc7wZyDog
Ffq/WkJjCjCpWYvkkt214xZ7/sUUBNPWPYTDtgXrWqbwFFi2aIeAEl5AiT1CTyr8WfsA1fDarAs4
Gynsr3A4MPPbLBk9hUK0rakeT+XQLXBu7UFBfuzhA8O/HzTqqKmRuQ4rR9i05iX/yokT2uJIpatO
atnfRrImrcgOugE1fw/50L8kIHv5DwZWiJqlBQTD6V93FwjEJNGVS1vcvjL73ZQVZNHpnW4knOrd
+jbp2Ka7GX66Jscyi8NjyS2fB55Jwt9ajOPa1HPbGK0esibXCUR0lRxfXrKsdBIrUnNX89iFlsNU
r+7k8FAQ3oPZj5+ril3ufhJYEGercsWTw2IPCuoWea5e8GrVfwL7v8FDXe6/bxsP9pUMMCrCsaEL
KZahNVf+AnOqaid4QGEaNnpRe8/saUn5tcYal+op9afX8o8HtzHWXM0sCLA6Q2B25DcIFJLQ6+hT
YiQ4IheZ5OthxYJiLP6UMkYLyAXzFIMpwZ39uROoqo7VdnyyZXKPj+XytlZFt9xeTKm9Kw/UTg57
Na7oHBP43UTCwimRsYXUeDPhat2sEtBwvPXSu9G/Dgh/AILGm2h96TbUxu4kUUw2E1pzaxEuasr8
EeX0Q5Q+DzZwW/jxEfLnPTFJm4syyFtbkk074u/JaLRP5VD4kTzCUdUWU1ja9b1xXdeStInAcn0J
eCgUbqW13gjL9bVTGjNOrobO/6plepFVP/WucVhpM2J4q0qBCNfduljK7W4u2GGnBpWhw4Wcxz+u
EY4wbf62oWR4cZgx6QT6BrWdOigdIH77fX8dQbIjfVMTO81O1v6UinRfty0CsSlh0TS4yXhC2Bfb
BoK6hhAxGSY/wTvEv9uqzRsSh0GkSTeSyiOdY3e8UNQzGt7XBkcYUsQGE3xZlkLSBPAaoSrAK/r/
ozu75gasEqDDeQ/wTOPk2vTqn8ntljWWEkDg1bCI/cRr7vcyyqug5z7/i0kR/JiB45aNZ7GrMrIk
KYgePGJFsAU5PLxAkLWMBR5sTyt1b1XUkFpLsQo3uhQaqY06I2Xxyfk6JtQ8mWx59nPU136KjDuE
ZRJ5i+gpEn3t6hBm7SlXcjLr+otvHkXnvKUSONSPYgI3VxhGrOtg/PZL80kP2QqerInXNedw0nNe
UtqxnBOmuG/Milzst55x2HNuuMnurwIT9vyPMRNzEtckHK+MWKyGkOZpGZUfXZiQ6lgzDO+ChaUb
9SluVweMcj4QW+7JIN26D24bNkRiDBeNpo24Zei3stsawwEGrAko31uKF3X9xxyMMDUb/KMhuByK
nk0C4atEeIL8v+29KVZSIYPoiE7lSG6rr9ekyVAqMQCbS55a0lsGp9soTZDWCtVQa6/Abm04URiJ
mSg6UyBhM8NiJKFyeEuh4sbs2wILIUALIJHuyudFdQYW6t0plgc0por19VVJYcIq2rFX4kBP3jIO
lcKrmLfIg5G1ereWYnwvYGkTWu5Rx0a48fwHBETxIG2f3h/q1g2a/GCLTqzeIbZqK4wT62/swAGr
PAfWU0FgBXgU0g0QN2PHrXjV8fofnTH64KWqcPf6XcpYnoX50iSBGr7NWkieUG/krTWQdi23OmBV
2mNg0zGJRBVzqN6t/2aDgZR7kd61bjh+7t2THOeGgxb7xOlZ09aTZXPP47DBtYT8eZ3oGsFXJQAN
u0DGp54rGgu1tMJx81xxGefdd23JpeaHxg9VESitS30dTTkGfptXOuNy3fCI7Mega7SWSUI8Ltxa
RWmK9c77C+n71Awl0X/W7cRGaB8rBm2WXpZfsFDOgMnsgplV1w7yQ6igUypO2Q40Ejv8KA4/VxNt
fxmUjzVr/RVaRq2GR1RPhi0y9cOZr+4Q45goLwOK71ofL2KtCis9iuw1CjdCcGe9kR625ZIGc0pl
tVhMEy6P2qsIo156aY/Liws9h6tj6XupIJmKo14z+5fM5NLOUh8IYnp+dQqXEiiWi5FPdAY4Lx3D
crcuosSGXRfClvdhFoHCmyhk6wvvnqxBzlkJy4+SHdqETbR+bZWjIkCAuZ6XrFpexMWXNxfD6o3x
z6niwZzV5S324JTEYDO+vedPT7oOn5qwe5WmrbNbgzjCrz89/Z9CWCiT3lEJvXvS38CY5Hx2IxPs
2X96tm4uzM1oTppYN9RjxLw6NLeD1tJxZzNG03wmgxjtwl3QQevJ+bXh1Ebx5h/sKL6ewTbBc+ko
esK46twxxPAAzN9ScLrINi6q+WoclNM/EeZKObd+HmnN5yNcEZvgt2qPaeJ2/WJiX6frCZzmE5AU
yG0tGIH+bcBhPSOQsJY3zqd6rVoGClCEdtfzKxq3ExM4dBs9mmdYWRhtj9uDQuunoC3B+5B6ClX7
wo81sNxePj+3HOQZHJqJFdJrN0wP6zv186RhD9svQy7Kd3kX457exkwHu1F+wynWOZThE33hsXW1
TXJ53UQ6L3Yfuvfeea9RyGluFac2+UufyEOmIUaUhTibNyDKPjRZYoXPXAvQzkHvG6k5hMyiUkj7
Drj+7v2S3uWphe8l+/VL+jpahfoLfgfOVHIzUIh9ROuX1wVGTvqbC2A1rlUiwDhhxPqI0nAvpLUF
/0G5M8Y/JvwSyg7rc/5ul+8tJ9SPr6wCw2hZyIPbeZWwQM8qzAv2F3nhUS++5OrVpxTp7X1MvS3K
vmGhglNLelRYvTxLvAYjYHCyPW8BRzrY+pqi69b3/bgpr9PBIAAm0vFAAAW31qnjDYHLUD+ZzhMA
R1Hk15Xsyh79G17+lQtSSWpIw1so2JVaUWil2mxkL5y//t77cUxET2VVf4bxLwwnucz40tkVo/Cd
zYSCmCG6YcYEJSay6wKS1WqxGU2UUeRdsyLWb+tGjm1ufLy2mIsgaGWHTN55oSK2l8O5EA+TBkjs
7qTIDed62ydkI4r7OhPrBYANKDNgKW3TRw8DYkCvpAukDvbKICKduffyklFuAZ3EuS78e+zHwgZ7
llCdfoYg6S1tvYAvedQ0rU8AwfU4XBvxHw7sa+7daQ+IeMnFU8HcKFpb1Pj3MpqfLaaOX+JSrQ3L
Ub0O/UtQhNhiJTA08PM3qBxub9mOZjR9TTyn+crrM2j3OWtmrZ25L1yJXNcHLDXztrbWEHWbuDYr
3pa5tCwNviOyMtEJUlu2NXyWVU6joqtGwbQlncW9YwF/+hl0zE+bhEBRgpHS8pcoGBBBbVtPSFQh
OoqnynIn1YDMUxHxcRvGMwoV+aFRA1+E/Ix5TDkKIb6OGCryRfsaWqRkgu+lQN1tUDwwqbwlgv+7
jYgRfGW/Dh8U0kSgj3Fsim5iI0BUjnb2nXnDPvyG64e3w3trO1IowmSzS+BPrPowxDGQKS9L1+ve
qDmKyhJzGY8N2Ocv+zZpUzlfA+uqs1mhLi4Nd/HzWtZpb2zO7s/wnLP1HZ12D5Zjp8AigNze/YHJ
i4PfBK6wX9aRoJKC3V/hp+Ci2PvD+k3vDp8cxFmgVKOxo5T02VgBLNgKT1isJKWSshsrP7Jw9U3G
ZIUoVE2ucM8HRv2sJd1qlX3H0suaAh8M7XRRzAOSvJiIDPff9lnuMEnargL5bmFh2JAaCJ5LYLST
bQ6byPteGOVRsLECf7m49ONWlECI+uZwk2nuvOqpfV8h5Lxyw7r3EvjjR2aDLa4Btsu++7XyOW54
Vz8qxSTlgm5DyK9ULQYkETiWqiJjOH0S/oKvWZTFQFt7vh3uugzP2AiwzqzOLAwUqYzHVQmbGkRc
aeNANbk/aUt+8wQK2+jCqOYta0QGR51dfSptqLpLW+3SKWE9YVq1Co8Sp5UQqORRdhLKSpIyp+uL
Hzw3i4h8xiYcFMZ6AUsLn+35XHtgPUYwitYTo+dhrgHhmpdsx0Tu5uOZS2dxuMJ8WbOFHfAQl2SW
0NWqDYfBkFcWYJsGVNqW6aPUKBSzv1yad2MSspAP0Fu3NB5CqoWgYSYVrDl1cuNqwl3ws+pFFM55
EVZ9cGoZErThE9ArOVcVSr/fu+w+6rcbDegq7CJEj5ii5BatRFNoJput14RKfg5PsycYWAIth26C
bZi65RqsxeoRhBroL0j+QlfpPTjA6CWZ3rVTlh4VgP/bFRl/5Sfc/9qg0JZ+R2Bw4y7zEA6Zrn6Y
eYz5DjFb2WJNJS+6GyC1nJkHdSZkW2/oY6ic2eaOWzxINFyIugFBG5SUJ9XcVVqHtE6TZMihY94J
u/przBuTlskesTmdtz02ld9THMD/Vj+aVccqtUxdqb8X4/4qCGNqOmVk6uO1GHCQEB/u7D1x2RiS
ZwTBwTqcbGmASjp6sADjQVg7OGooBh3IvnrDNksR/Mp+mMQBJS4b2FvoPt/XMHiYx7mnJj5VQ9ek
Yrerp9tbd7LsZZJdlEYNjkA+qQkBvDEcVLojyd4eYI/CDZ4cnKurUlQh4bxsIsIDFn5CnxzMKKNz
Oe026QOPyhLNv2uKwkG7b3e5wvFuO0GvXe2jlFkCgB58sicV4BNbTyruo5jsWwgH1nX3csNJ9wAs
kS8+aJL1Z2ruww15xap7BuXtwLUFCLhSh5JoAKhnh9qLXa1ShVQTrQys5MPTg2Fgsg9aJUXsjmhT
ryw0qeSbHkxkRw9NgVs10+9tnXQbUqoYODf97ntCHbQ+dp0LJTw1iFIVb9X3rhnmgtMt/BBFNuoi
XejNkto2TvCwwARMcHZj08YS8gZSGT7xRFOEPLeP9vw9A9T1VrOZGbNtTvTR3kvgV8cSj/VYNxo9
W/sWyRcok07IVyfCjyrpz8oGgduxdgrYnC+frp40+h2x3iGCCukkkXJnC0ySTwQPf3JyM679GY8L
6X6+5j02SHevH247oaezMTchUtjsiOEfcvrNTJwY4hG87hjY25Wq+USFE+HhObHJVpGnJUJqKGVu
KI5+hmwWUeW5y4Gqe0MnQND76FJ8vNu2yGzPy0LHU/OI9xTf4PkD0pTh2L8B2bF+7RukyN/iKWfo
CozdNgfQvuwME7aRth5gOVHYLbg2524Tcd2EGkIivdVNW9BLsxCz+ujO+b0Ie5fvuhKeCWNjAWOp
64eInLYsS1LW/zaIWzd1oJFD2KO2YV2u8Qkp7HFWEaJ4eCIaK720VPD7ZFTFxOStyYS0wlEZS2eY
jnVB0kXkzx1Tjr/JSxbFDAmRt+hTciGL+E/3OPBcGRmthxgQEF1r8TM86EOBxi/To4/grDuAm92t
DcbDxy+S8YFypFlZS4GbKQVfod2er5mDjfW00p2F+qd/3WVXo5vGAEZRa/G6wPb1gw6lZ7wU7w5c
b9vCZqad0sQlwVoFKKpNMkxDX5Ir7fbt/3hf/rawpjhfgqwMVqAR8uhTvOBVOr6fJajruA+5hPH0
X4lMJapxeMXSb1vYdf2o3VEtIeLklSMV1YWE4PcoyzmsT2pr0XedGVVyGy/S52Rhn47CWZB1sm0s
MQ7SVe3UC6nzTFVNtOhamY6bM28Qv3F4w544TpUgLSVSQqUo6DFMCh4wvMnjt6aTulqa56AkFjgu
b+PZYD9bhMRFXnRwhrhP4ZaVhmQPcinPigrj987X2LSY+wW2De/pQBD+3hMw4IYEIG5YkwwufAEu
0mvn9HKSF/zlSAQIeR+nWB53YISTzSPa0vw4bS/Bu6R7E/8gdjJkXBQLror8QeUxoGoerZe+MJG+
iMV5zw9BK3UZEshPeoC3StNOmc7e1yLMX4oEJEEhg1IqdEsWc1R1DMjNgPIYrDdVUd92iO6bDIC/
tqwKhJEvGFXF2dLoLEZST5e3/wolxiQjK4+rYpXMtjevDANMwMVRXhSasrTef+ZEXVXuULlWnTPL
Vl8q+Bs+ofWarYjLkAYtxz1XUrQeYjqNcSKFXOx+u5HzTwdRt0al7vtD2opCYInjqWzbThe90Cpy
NTME2kn4R3/Er6wEf4WvQLa8vluPx+sBV4WPVY/2FQaKji45ciaA9pXAzu8Hyqrxf3Imacz0HB9t
X5n+jll1n6MNtU0yPQTejL7MSpquOz1hPG05fsTwa3b43IGHM2fbeRdEI+ABsQOINxNTs5O+gSPq
CZWGAyna2s+fW9rc9Osj0q6zAMOGCGHNC8R5+PTXDCLcpc03S1HO0pxvfn/51syxvfeeL9YRXO0V
c/FoBcWOBuN23LPSLW+Ll76b+ZbXXzBGHezL+L4aMhK+myxtbUFuAJ6reA6NM52Na3mYMC7E1IY7
A+M+/U7FQGK3ZTEiSsDmLBmnoFvx8oRX9ECtFGa/jJTKtfp1+d/sB74MwuCJ8ue0wOyhGYimjIDF
bZFjwenJQ1+Vax7Z6eXhXFKSeZsXBSWZgeh9KejC3YNbrevOswQBLIy8RsZM4pxiQ+mCALeTf6O/
XWP2+tPKpQiHTwR0GFUZCGBrjfuMzMmAKY06EBfWt5pNiiTC6DRuwY7Q/SKlsKG1xNke12tToX6h
cNvPbUdOUSlL4kpV5BY/AkBKowrjyYrDIXNZpHFfAVi/U2gS89SlWbE0xYCcRQHuroQE1LStgYSo
rbMXyrAZJq9a4asFPp0Unu1pNkkO0sJ4RuTVKfZRFCETrcRD9zrpV0Sn9VeWXthEGthCDKnPuZlu
WPnh+5ZAW5jOUyTn857bH4ehEV6XuV6N/Qt/qUd9Pj2syjibqvLqPzJSnMelUWSgQ3wJtGza/oAT
chvoztcOWMWgIMQ+VRUv9v+x8ymKC3oo8UfS42UTeJKfB+uQnQUIixU3xxctEr5qIFCfMYYosLnx
qgELDVBKAaW6JbnKBAUzoxsWhp07NiwFaNqMXf8Ij5ICGbFFaSWmOE2Aym18TQvf1nvrp1OwWIQc
N/8Cr1W86OsnXYn8pqz9wSeCZ2lPpwOJeztVsiPPtPp+9mCbep9JFtHsgn5wel4e8GxzWDOk+eRk
3+FaYVCN5Na/LDX2Ez1fy/0v9i3YGMYOHToRqnvGYDPjo2qDucz0cD4G1pEE4T/S3HphZRFBUQt+
OUMLRJEeAQWvjfPayrYgpVpy1pz8bI8vdKwUuiQvTNpmlmGg3BPS3+7KdOpcGSR3Z11g6UWfy/mk
XAjZJgpRM18NwxRb6GjX93LOsG4tCj0aMHpkx9fBlxU7hmKA2UDQQU7z0jXNMn3ZVpVfStTYK7BD
SHHCsB8ZJr9pL2UcrHq/419Uo6rOukWIK+SVp1yeDijUY40cmHNeWjvHDj4wQYThs8DGeSEdcoqP
c8Pnpt307Qp2aAwnenDUcu+x6zygaDsEKpOut7RsMSxSidUALUSfz5z5Ne2BtYcmwKicYkQc7f01
5jTDQM6w3XRo9HzkIUdOwA3D+r6PVolDOrSaTj0Vv7htyMTSNBr/vn0N93EtGt6Bw07EzIaDiccq
NMqKDB0F75VN/ITbfeZ/NyBfPcGR+5HeT1JNiCVjbCaOqqjzv9AMDhK3kvTcCbOLPZlzVWwkIYKg
BtmP/pqH49XsP8QQf4ILvMWKnwQMh+PNCejW7rqoGQDzEJ5Wqf8lZ5neugFGbi1nJ3tWi9MPuA3H
zmG1WkUvi4qnPbqJaABDV4CbfHGUpXf70aULRoaUzh6I1kKxaHj1jojjN6D+C8SKFDwGVjo/o+UW
M1T8cNDGC7zPTePmnVTW6NwZSC4t9webish5vOT+8cUaOrdxfu2lb4FuXTP43J6nQE7DXh8YAwKb
buGsHtfGi2/RbUBV/LHo6Tw6q2pEbNFmdIU1hjgCi2wwXCCM0YLvqLLMXuIuhRKJqGeAQpYda5eB
gFAxGaIWiDsHR4PNAPb82mCSHWGYcWV+vwEsca946Izh9pialZZc49GSw41RXwrcVxYg7N6jx0zO
LS85bJol11AVv5laO/EPovJLukgXn6CxRrCXWhgJ+B2gm3L4cc3PrSRnHt9z/vDJDwgtpxUYuqix
RCWyq0rNz55oLkMJajIFDjsYd+LvBT/a6qX2IKjOMgmSO+ZUU5iEXPWgd1zouD9P8YTY/CaiOrp7
iG3LuMV8jkmSpHJT1O0GVtl2IGAWQhPN/lMNKkMA956LWo578iIzDpdcfvejJwsURONK+r9Ir9S6
sG9WMfXZxx3nojoPk8c5iwBIUeH+DjFjCdl4suJjshfmRUqv/2ShhEgYsWmpRjUPWpadhJZOcTgq
1Ps0uOp2+/keo4F0F+s32xx85I3LC8mlt57ZLRbRcWAgbV0ml0dfy+wj8Z98c+qegKo9nO6j06j9
Igz6YeIM56mYi3jFoxrVESS8scXjum7tSFz+RPz7+7r+sN+QFNLszOYJ5apJ5JMdM2ei+XDQmktn
Qgt3Txlzxz2zuHlgasdsgz/GV21KIT7wP7RP2RA29zE0H5s5K7drT0GUmSEMRyNYET2a3/MzKjQG
TcraQLJw3YC5sq4M7ImCG8gOk8fgSjA536AETffl7+QxrcXSk3suwBhnHJhqoQQoPaoGjNmkxtrq
gU4J7/vIEP8SlrZmTBuDeMJ6f5IlmwZ4qKbk2ey1bSDwtIozwRdFRQmo7obXmbJ6gXafK1Sc0zsV
ACwnoxwv5xSxBg317rYswyHjXhSnBriEMq+3MBS/yhxPQOJe/Rae83dbmZJplo1JR30W/jrlZJNE
dlnw9vIdQ4AW1h/AulfuAfTVStsJBCqBHclwdw0JzaHrPdhli0vBxIo+DN/SaKW9YUPVoAwU7ou1
8ILAgLElHBFz2zQzQQEWoN4Kmv+nYZEiBLJJh/aGyrjEK7+Rf/IKI/aid1RX4CUubcGD+FOqd+ex
fi+34724qREplU6eFl5+lMWoBnXiQKLnCsG/Y79TKEI6CC5zW3F7FuiqQNsYBau2KMyHT5x+bZwd
G6hrRLCM0oCZ5jv1cv1Fzuq7dZcFeJZ2+E2Bjq1NhJnb8bif5E6mxrQm/73P0+JEd/Du403kFJMy
2FtzN9N5UsZIHYiAA16+QiKIMKcyKZApIBZ5qmREPDZ7PBCeY5Ci1NYVV02gxkgtbFUQ/YwhMQSi
fNANzQLXSBxz2TLr7DpwpoQadImeb78mqAgIj809yZ8siIcbN01ld2PnWst/bTBrEDhRz93/2BV+
xAEBxu35Xm2ohEbk40acTdbYTpT3kNvjqwOFvzicehmqGc8aXhYkoL07McjPc8+gRVVcjzCyvqsI
Ux9a1Qp+WiRK6YK4MR+jEP9uR2Rn0VmLieTEUsdAGVMrpWNqQL3cgZBOZNX7FS0tViyC+tgQwBR2
FOTtS+7IJdZOlaPye+aXA7luCXUZVYMNgEOS/wqJw34O0yAsxBAFyUvN+2Ln+hdxojUeSLMS1j/Q
nAzDPd0vVoo0q3C8zoTLLM9vQQ+Tmum8jbLj8OGzrP5mxlIAMtRwCow5FlT88FY2zWvoB/7McDZa
qBNaXl6Hf2SF1Hp0sTb4zjh0ov04+B1CBMIVQMTYfroMIxD+e5vx2bEJul29IPpBGSaDApGkyzNn
rkA2UqQCCqvydtmvpXyvzx1K4Zv/htDksW24XO5p/LGecbHBpyxxX9UVkAtRuYT4aF0y5ugELLet
Os4v9lxJAyBm2H0MYwACb+xZc9X5Rmsi6+dfwcAgRLr+2Kpv5d986f1Q9DHE15wWD4LBmNfSubHa
cyQL1kizGy/7wWW6c2FkInKeVjyqyU12AWg2eIoIt8IorDKZOVf5NQego8y7wqEn0sMiX+VLkitH
wAkHcmSTnqrh85k1fhKkDZ4riFSWeXma3LmQYEzyU3DHhmfRiEUKK9J4it9/nyvSKaFJMWpdf7CR
7xWQvWyfxSTv+yI4850GMCE2qu4XBzld5MUkbLmaEkaMrTheNSYX53zDQd6MfSUE204va7Asss33
lKtpVV/+XIaas00vBlGyzTmWUfniIi4ZmjPQMDBsB7YGwLx595Y+Am+Z58ebDKiOCZgwnBEvp5S7
tTpOMTX3hU+t1A4r/Vj6Nk5oTU/Vt0lWn1ShGZ/o0hjBCgMhbEoTUbdtXi5mLrapxAHlHi1mobct
zNn1ZA9Y+VyrpUN7d2oKGrZvV+jQ9Efz2vOP6m/2/c0QrNJECCvCZHNZYV7p8hzUJWg2CiHiK59p
WT/NQoguzmf1vVZN39doQjqf2McBDjh9UEMu181seW7ksjvoVqrfnESXXOoOPsxRsOjwhkju7Ax+
8LHWUwQefrxvnLYoJdGfJha5cu4Or5Xb5m4a+xPG/bbboX9pNjFnYtmv4dFWtu7zvtPmKrGPCNRe
PCFyJZpoVW+i39FTPo4UqzIbzYte1LY0sUKRu+uV1PAGU4uQ2SqLzhXGb/us/LGxOCzU4MBOerUh
p9hj7Rno7U5qf4CN+bA7ZpquwAwTbQQRi+uCgbrLzIAdWN6QSYC61lGd7VCXSauI5NDRrL/tejPO
Hv2Vxm6xMI6cb7Plxk/GabSZO7JBcoGbhrMJLSAWVQSbr+JRtv83nCPpXgTMe0aMV+Npi7sYIBLu
Pj45iECft1bVBZfcXIj+bIrg55FupFA2tGmmb4pCmSf8Tjy3dn1T2UBV1C5FOFl0kYm0WuIxQ0uu
CtAHdcYNK4V0H2KYbZ6k/J6unsCEHK//gG1/qiQEe2xrT2loinHRK2bTpRl7uDRqebJd/FW6sacs
ZjMT81lxYZgcAKU316ZUgqupitxHAXoKZijdlNJUZSHOU8eS5UwJJa4XRnewJnF6tbcjsM24fDfI
hildKDrEtOpjpPxQBTIzJ8ADhQXaskcT/rdien+0zAcan/BivkYhyOT5C56BxENWQ1mCxb/AY7w9
JXY5nDsNajk8P4lTL7E9QmxXrmHTGSYnNMtDRtFZ6JJnvIm167W84QAysiQwKBluHCrMoQdeW/wt
xJykN4X9TvZ1XKAnRJvBJduPj87y3OBeJdEAhvYyfw3asI8mvOjr9x4H1acHPXmNk+FagenKk8/2
CDbS1GOYHrvy80co/c6+XpiA2WCVdLVVSMhvfoDFqvxLni3c1APeeP9dNXDfAyk/kMZ3Ul64V6Z3
NIQAE8peydcP6YOaZ0aTziphCN7Z5ZpC9RemUttDJ48RGpKNn+OO+R3n9h1TJf9pVeQwhovjmg+j
qlGyojYGZIZ6bUCPRJI3cjWOr0LqpF8FBPaokeve80ugGvgJrTRZXvhrOzy52g9CawXxfBMP66iz
WvKnSeBPJOnEmPBIuIWDCBFBnWHTzJroEX2TJrIWK0d1OtRdGAnzelw2CjZZpxvetMCS45WcjgSu
knc8G78qbIJcS+tQ3rrTFa85b1BdEXj+nlphyBPlSjSdsPF9uP0ONl1agZn7OaO7GCHazOy3KNI3
uqhHWaipgq/m7qhMNEgt9y6vU4Xj9gX++6Yl8Vy0JE22BF+WBx1X3bkO2p4R5V7C4MvHLBQPNLqL
io4nJPH4BDysz9fJqRbfD/qlfwjP75zA8Ue/xW2/BC1r+pCaJzDb8GxCUHNfdsnR6lsqCC7QfMSB
ybADKLfcESd3BxUk05pbd0Ohw0EyBbRBaFbkPYwHgzxrh3Y8z0sriPlmYdtPLX0N9YjJFDCWayTc
2SWLtMx65yzWDVL7SepNnOSAZt7NwVYkS0DxIBIJwBF789MXQlHXeI/GHbhCi83duLBzc5qtkUnF
iZIodMz/hxXVZJm/I3pj31TgRXNOslXAtBn/s8kBbNHZL9XJ/zmxh+8jq8fFKH/ik5x8jlNh3D5C
t3DfxTwWNAy4Ta01oKl7Qk38G+Zvic011UbAXvrqC9d/k6BtdDflpXHuYKV061T+hmC0It8GNRwE
nFX2pNBvi6dDVXD61wvfMIiNCRmYuQTG2+fccAwX0V/OkC5xMjUj95Udod10e+5RSIC4+M/qXvOr
hXXy0r1pZ5gKqjSAenmqlUVf7wKmHKv+c3wFBCylVBJmO9ThurDXsOx/6TEWwKe8XXqQ7thxl1AX
3P3a0pvV33TR15jYUNmCEkE3fB6ovRLfIZ5Kj61kILIMr/eoQmIcu2tkj3x/hk3vDjghuWVoFuTz
W1IehJOnwraL+tXhxCPxmw/xpV+tOBnql4Gd74UvLy5WwbhOHU6WBEsqqIImgBDKM84EgAVZDEDE
u7fssIsa2l4eU+SRj9L6PFZvoLkHgC+Exojpra0U/+HUWyzn3L8SfZQ0zSd+aCX8r2qMzoQ5/ti1
xbmvwyXAknF8s/TjzOrvvpOl5liMflf10vMxeXLNbqDxRSmgvmn0c9v5+8m4+O0PfSxUd8OXIyON
2PAXgTKLNN2ixmPBQOFaELXQ9YIy/4JLkKXvo3X33u44IW49+/HUQvn7yOVdVOWyPPasv6v540Fs
gE2Nn9pasXAkEYtTGMei0WwrzaX4gz3KMoLHUr8o/V15xFtmPVOryzUoZ8tfJiEfRcdjgPERRDTi
4UQWdsg96mu1VB1r3JqEXJ6WWeimGMKBIejAnzVgpElSeRXjEEB+H5nVFEoL3V5Ht7Jx2ez4jcWM
G+TUJz/bWx6bWrQOfqqtMoldpOC2VGxpJDZ3sCvetEWGbx8JN/FQNccS0otm5D7Y5Dt92wfPTkK+
8AcBMg2oIZnmwfwjnfJHxsXtusA5X1n8UQrv0Bu++ty1SHgYpeOUP/wThxjrn28L2M+JWi6GdFqm
6yE3CurYjLoQCQ16YJdkb9R5eu461UkfqRF1GVEPdRsyveUk8Ybh/veRJJbkkAtOkTZfoRJjMcTZ
eZa1Vs5q+Q5PJHZgpjlwCWP0l8giFbVq2Gkgaj+o/YeRp/vI9ZUSy5shujGg0jHKhj4QzzMKQel4
1DF9WTSLxgY2Pq9toNa/2Xzy+WgX339GK9wlIEXDUNmp1GrcXaVVc9PCPt4Mh2vn1ouqrEAu+U3r
FBcTElxBl33vBHwP54nN8EykCahYJAIk/Ez9ulJplXELSMk7uMHUGWpPq4ex15Dz6tAOvi6WV5zt
uMv4vgn1jGhM0Lu2nV87LI1qNXDrWbYRexzF0gXyhZyhIGQaAVZj17j7bG+GjPyqmG+e7xzZOapp
xht0j7cfs1ZD1bNzreGE9phlSQOZ3FxX7OJUO5SptjEUuObIF4tnh+qVxICmAuRMPIJ1gPNLZNgP
JjM6SeIUpYob0hSpAXWPQVKTi16l5nP0Q3lDcn47qBtsWK0APUfJFs58JWh7WANnXuTqCmmOqTNj
qg/UOrDRMYPy11uHKXrjRYYNyNL5g0piwy9yZBd5POR1hc5zjB0FzTHESTNHOSKsShV/ucTdRiZI
sZlhaWW9iIsj9kd6p+TmcP1g+PLfaK/YsmPzuWAqYKFPle/12er1oYyBvbE1+iNYS5+RD+KFAZ/I
N9RkO+96DcZvUSvCBOJE4vJ5/6t3O0cd5SqsdQlfQOVLZvyLFwBe78s5VLssfW/IjwO1Py1s8DvH
Iq+a3u84JYSZxD8vRDduNvmuTOcC1+MpjJG1EXIReeIRES1O8I7OYD8huOEQveGYdPBYvR21lIWb
0b8tanoZjNpYvXCerSNBA0DXb6vh84BHWrpgLGoK+MkZWQisgTl5WjLLP46wvyfyerEXL3ICd11p
HCBbHMoDQiSYxP7M2brGOxEaubcgmjIqrNxbjrcCn9gdOxb28ZagLmqUJqfi1D88/DokKcEVCWLi
Ex8Qk/dxINuTmDFvH/bm8VrLCHr2DfiLqZlv6tRn4aPT0YdMMlIXoB+mxvwfpWNjdGkwlfgCzAZ6
wfRMoqbCLvXLCowwhbnkK6uLW6DFtJXBMjlxz9DoKJ3lL3QJSrVRgMDRriFdEyfgJGEqWancjaKG
suOAyqZFEmjp14bdrUXabHSe/pBmkcgu7e7Z3YNAG4Oe4YOrFwSZcdV2aIZW10VwZle4d3HzxRSt
1RhtofS6U19ZzDinDwpmsZNsIDQwpI3Q8s32QFVjQyrD2XL6++AuZLYPYcvk8CyJfsJ4kY4OAQVU
jDrTyZlF9byKNLb5XBl2vY//G+d2FM/4eQztDHGD2twsFWTpp9Dpdp71L9Qarl8HRsGaMo7eomYW
igYozjKEFhWm3FggDShzEeBdY2yJgL6l+K8N42/+2A5UdGJvvxBBxdFJhV8+g6DYjO3IxASnbaD9
jGxIS7rUqXC4V5UybrchjUVEwusGwMPF5zirkKJC1ZlMj8rR4bPB5v6HYAdsXp8d9LRMYMYpFBAR
mYnHy0bFclwybhi72uPIWon3kBxzoKjMBEhfl8Y56yxmtIu735VP5sw6zj6Xz5un2xFY2NCTGNz/
lNOJLZ8Wlh26dcbm+61NunfYNBi6UvDyf3T0iCrnj4bqm+ie/52DryWlUCdx9Ne6Xaau+ADbejpZ
PC1cYcOTvGNCkvD0RYnCLf6Ofl/NXpgySYpuilcBguRoT7SsBqk8Ae4EexmQKkQnJE77bT7oIKkf
1XcVJgj0DOnAK54xJ4MpVzEFbswESiNUXQ8LPxOAJNk4aG4sWSvQZDAIHG852MFF5PmP7lvqkSEU
tS9Lt2Mu1ZlbNfMvBPWrEVE7UIMksqbX8ukWxV0pcR2/1ZqjJiMlQK/g+694EHPcSD75unzcegDs
qbASa4N/ORvvd5TmYbW6pFOy4yaNy1MLp1myPj+EByrZveaet3xAkkZ/YWlPvS9sxMsXF0cu6i3O
yeJtfn/WWGsBNIpPvINFcTzthfVnsKDT/oW5rTUklkAdmOz4GslZhTW2vVd4ErpOyiHBopcdAYfD
DkWGKhuEsPaAoDaaoEnNJi/kdciQP2cTKUUvas2mm4tAJk9pWycDkPb6GKYkrDS+EB0AGjhMENn0
tcTjHUNaaZdPYOj5JaYAo6I9EqO+q+FG87GqEVfBfPoXdKd8y65dG9LLGTAI5nXULcV8Ch3Il3N6
6/Zk24/dEWd+NfqcTROcd+LwmhYBmlFG7F4Y6+YsgOErCNzlS+n/lFTJJl9EiDLx5331lWMNOZzZ
yqYpW//pAQO0Zx2BJ5KHQsJ90QhwZO0eLXbWBBdq6IWyNmvORGMQneMs+DHYvfGTA9Q+UfVrTkv2
hIyJxNEKqbakX0dtbuwvL2EokVomm3oyfPXekqBblBQcmT+ST9Qs2vXk//yDitBwH1I+8yejRYHW
eptIGE43owwaiJkwHw+q7aORvC9KwVRdXBwLg1vs56thZq9tpBq+103veOyUtqhFWU5u5dENFwnA
8NSla9ybc3w1ztPiL+ZHzrNLuBIs9FAmLP2CQwg+XU/TsLVAUkxs17z6bnAa9m4M78i5PfonhTFC
Tvxy9rBiouMn13yhfVulhk7ZZQytXmX7lND2lpT4wi6UmhforGxVQAJkkWru+fcUIolDcGcmf1uO
iNlpfLkbBoIY7RtwVC4RK/58Msz/yMNq6VeI6RfzKJPPwofL/Taxe3Daky5omkHzk/XvDiK/cpew
5gbtaEwiEhSF6sT6TB7RjWGvAlRU5Zx4VlTK761KWK8UxRQSkjxvLgIA0KDCYIO2sBFejjbPQBd8
kuo69IWwhdXWC9X6G7rvRK7fJKmNCq2wcWKYhSS/lJYF6vzVAFo7RkI4KAGawFub5ADfRITyYUmM
4Ssss3SbKRxHlTRhnt7+V3Ssrwto6bnXWfOFg6wBzRLUMl90lgF4r78yywsK+PIyIGtIVSWnIvJY
k1q0ERx4e+JMXFSSAiSjVZlBONY0RH7+Acw4jM71Y3dbMpc4EbL2Pkb5mSHDnxnL76I8gS+DOvtp
H0mc8k/PF+Ap6GpM/I6Bs+eEsamyPHLXRFQwWzfHCUpG5T4PSNLs3tkt9uXHzu6I1CLKKoLZiIHt
xTg9tkpLhQfeRgB83yZBCvx0Fmmz80iGtIWYhJXMx26ptCQfIpa08BbWeRpaIDrhvmCeoq3n0ADm
mf6WIEXDxDc7mWKkEOSOTaQdAf/+DKCdMx0sKgNs6kO3pTy83Ew/FVg6RmhaopcFOJ2SOPkAUWm2
FIbO+uzcz2pgPPYlrWSp+a3MvluKqSDweZw1ynRRj8qo/KV2G0xydvlNqMZ7TYhNmMyifUQwFvWg
pD2KwEaCzZhUWRvbIEMxa6vBzvKd1EEDSu2jDUibgsAcQRtTBtOrW0CvCe4+VhRj1SSkc0mmXxYz
LGFAr4QwjAfO1Uax8HwAvuIf8eZsgA9WJ1JosURUssZxpe7en1qwV5027HA9Pog9cUxpcfexDddV
fcmmlk38dHYfiRtC7f03i5B7HkbPpja698yQwfVoV+VpdnQh2IsIhgSSxRayauhkmPWVGXuMRXwc
LzMhrExNHozWOYqItwy3vu8qu5RlxeaU4/cWKRpnxhAMAbIAoDEJfKpRUi0/q/8ZXhlTi5A3rDNc
KWcW+LvchJOSCDYhE7K0PEs207OGeG8yb+w9lMTYboGUveHvFv5F8281b5VcLMEpwWCcEHddX6ey
Sv8eXJqQnAWYdbH+YoxM28VPI4ZJT6CvDDFqyj5AsUkM4U68aJfRj7u4SBvMAWK09f4nrpBqFf21
KaiP0fstVG25xXKZ4hL+SWT+LJRg5iyJ/KVdqERn/NJdgWOL1r7SFR9HA+wuTiInAyBF/40FpgJu
f9REZIhSUPWEftLCnmlE7tPAcFCac/tzF86elpPOwRLqo+aPGBXwWE/S14S2OzFx1Ro0Ud1qgu0m
MRzu8Ll2/dGSvrzh67/Zr++sm3b2Gr8t9fxGhVOEkfdKBH/5YGJsQn0q3KPa/UL+J+4jZwG4MKst
n0fFXnSt/87Jg0knIVfUxdovq/tI7iYpLn6O/nrTiPwhGh3Ig3yfC4g8J97LiLL4GqR9Inm3yzo4
t4psWxJF/2Sg0KAlxdhw8nsNQqotRcKprFbFQnAVXlbeYyutDqDY0P3EO1JCB+i12nk5QuWKxhe+
gdxLo4p77so/3kXFLGq1ao2JqP14bF8zZIKuDVEWdT7GqfeQKCM1zCgGiGvwIY5Vb7aRQEkTClc1
4aKwNkGQ05HOG6NST1sLIfUXop4HgqvERyJdN5qsdVyfyTL3ADPs5Yj3Mp9HMrSyRromjHJvp4ex
v3NusPAdbfNlnyILTmVn0gLnEfAnL/ngLJkLDOgPTnsrD1L4+A7hQ6+9pdZLojtsJ+DgJTO6ykkB
Bwxjyyac+9VRVK983U9zyZ7Foi4c9WlAFkcjJYDhcgnGgt3PPJ8bgwRaVyI2bgTTrc0oyzI9Gzkl
Rf0sZAf5BZ26kPtHv0gFZsq77h2OGYJ7npiPvFdFzf/3heSd7QV+rAjzv0tU/kf/PLe59vlrvUBi
bOuPCrg1UCEnCYgd9tyBv89es8c/1mEddsMxnMtRC3hcOxFS7C4BsmTlomvhfHBOpaKD2nsc8gN0
7PzU7DNzk23jHIEQ7fcQoZviTW1cxqZYR424q+vPm+GI9aounLjm4RfYLJyFSWa5ijTAoaoM1WJT
h6E+Hp/b9icAar7C7/KGA9cy5SD/AYvondIVYLtHE24PnL/rBc2YzVlh6IkQne7hrsu0Lx0p0tL8
uPC1Nf3GxNMPHV3+mUNoDNmXFK9lTjEr5hGGPKoi/Wnw502KnxAHzcFSMXOBlisCzi7/c8qMxTVM
L2IEfB+7GJ7TKx3hojiLovhWZufwo1B0qvHO+BrfF0HRSXclZ+OApetde4MDvovBoGW5dcZ8gofq
mcl0+D+kOl3aDh52KVNJbeYUBY3Bfkmvmxzhc/y3pAiC74fKNjIoT/1LpDmBKaT9JnhfYbuSNZz0
Qu/0v/r/QY5PONjs+SrFwbfz1blb9IqDc/ny/Uyi4Su9CEPgBnnLEy647zLWKjS2JIjX0HpjPAgU
jX+g9jePA+p9pC/FszE43qeDa8LQT1MhjT2OcvYlg52j3OwyJUpbFFLXMxrHKjJEr5fwnI7IRTVb
j0TVI62h44CDYm3a1UvyfvjCB5ZjSLiqwN5k6u2Drwx9yDM6YfYjmiNMmTtse4OzDLZerY8CmlEB
wtoU87gEA1V+UVwsbVeb5UidTsUpOhmb2pKmMWH6AoH064y7FBYTVvMuP8Vex4Iy+YxymbFdDHcN
JQYh8u6p/l++k5UHNHAcC5QNd5rJRz0CM23e4yTxhdx1doTUh4raWAFfjyW5buRRMpL4Ejfb5Dkp
lbMJVcJ9FDXsXsqzkSxLNlSkNlc+//19i4qdzS+OklXK9lMKRB5wTi5uHH8t6RdOol08UIzKgHV3
vCujjl37+S6Adfh4etB+OoE4iZSDwWtQFuOPwyJOE2Z6X/D+6rHRA2s21skUEoEXSr5li7ovWqUi
XICJv6VAtlmwWlBRnKvuPs30zmB8g0sw7S4Ab+Odmh1MjjHLZ9X98oy1HH6D1wPcxOYWYENcRrt3
7z0RHOTSFRO2pHCxOf2y5sU59Ziq8I7gOx+7f2gB/JuYdiCc4JxJJf/LawgveZ5H2yzNCJeNVGuL
GWWU24UWM/be9S2htM4orLka42nfr/dP4CgFbKVuFS3VIePUrw/vnnqGwHgJeXk3giSTrOQf15h7
XtlKEwR6zgxgnYpDd8QZNV0fz+Tn7B1bRJ2dpBUaO8JyNHynnXRwwTqRxRfwaxZ5t39KwS9vBXP2
Mj8+2nISmS71Ak8BwM76R/SN2YSDAu3Ft+K0rwKRvgOrSJ84/sk7WADiWjCGDdYKwJHKGLNtAmRW
2JqR1cXiOZqzrf8gN5frMhudKS9cySkQGZ6jGWBgrkX5m74QLl8q4UMDT/Z5RP8CCFpLCA9TpD9X
bqKqKwhLgGP4D24XNvfIoKzsXP1QuUo53myYY8ejd1XjfPavUfL8T7Q01YOMqx4lWWVtvMWlLN1K
QUbUBkFD/lQl5LnxVerNBg0FNuBCPsS/kZV+ILK5BSZUnd4cftDfnt4UYbiYF6pq0T9qWVo9PevZ
d7FbHFvu0746ofX0NUnqZTmc744U/B0h6y/17O6Fnm0/y0CvzfrY/U5UNMffCMwrE58k+1hUDaoj
IJ/SFyKE7it4C/hqBMAN8JmEFisloBYS+c3lrgWUhdJ4hYjvdzZlTuyQLVRHE79g5bRtcveLTCxq
DAoqeA4/cHusUFCYeTdZCS/otNztmjtvo5OriEzY1Ol5YRiyTfzGLnRal0AhQJplyEbFe16qr8Vm
zlchD6A/qjPp4+O5I6+OlCCaaBK6UYvzoJZThKg0jTaeij7gj1rMVmFO8xoMFG0bQS13Awr6f06t
hD+8JFuInOb3kKLvjxvPQn0oqzF8C8KkOM2LEeNavyj50OYSde7uYKFUroUB9iK8iuGKKFllOoMP
9pcMtOucqtn0Wso92ruuHSPsWpnkMAiFU9qG8aY46pIx7LQtGRSKzdw47f64LTlmYupVL/akrV10
3NpDUfEUn7Q8RGDxekEgiSsai4DrB0XUDs5DFfbQ4f8pWMrO3nd2RuAbLYp3VIM0q/hpQ7B9p718
F0Ae2qm2w+EGm+ASiemwiXoeY/gqhx1p45U7JG04PUYVPAuQB0tXcRItO81y4NGt4wJeKxFpgxcY
li3mQeRHKHp/Wivln2+2a50cCXtubX6VYx0ODApC1t+qxR38PLbghWSX3f/vX2CSVvLzdMFfZRy5
mTLilgZZF59RL0+U+0pWCousmt3O6OhKO/xNkbIUhvAHw7i/M+ts/7sP0/GiRQ/lKp+lt2lbeUoT
XFt2cXx2kIKaCN3xWoJA/bNTzU1VmUXObZPpijoYlaMFl7tUw/KWEqKDXobI3Dxljmd6gzEWsZTk
D40rOH1TvOUTUFGL2mt8q2HJMcooVws+WQiDASxhlIA1vYIxvjnXyclai0kej8VLwETwuf3AiyXr
/1uPSfEP3EAyw3qOTTlxSHqBhcRXAKDvjVI/lvyZWNjmcyoct7zRI37WuCRUNcNDeorgShk1/bT2
F+A5hZ2AO0o8PtPXNXN0grYncT979ygrInhZSSAxY1keK4jz2NYlXTZFedZGvunSIHcyA3hxK4BF
ShKlLHqdri9q2/7BUT9XTjq2tQBze9lc6qbQtOLr+ZXBQKNWNR2MO34fMxfrtnThE6YqrINO5vWW
f4PeR4dk1A3GRnqeyho+IEE/iTjFCsyHih3fFfE9ECuNQ24Dp6ESyf1n37kW3qkQrnvWlH7PN2nz
Tdr4ObEC+m9HlQU/FNSr/Ymq/E3yh/RKzA+wjNTxJ6SCnWcQoNK91f7L7T4vL3SceOQLUt5iSfPx
9EqDwf6wFrLEGMKNjc7y5rxGixEqR9kOqouq2UewGcQi60MpvVkCESp0uuu7lgypfua0OGAfzqS4
Aoaol8B4hhs/KTSiMcxuCkiaB0Pc9pDEJtngJSnRMR2K9c+ANRyOuqVaRumdQyBOqkDiu0uHD2EA
6PX475KfpNwg8TWTMHrY8pUA/w8Q0j8YdtxvGD0XE6m/dtWCSNOMTe03HEnm87KSUJE1AT5OKTjy
bWpZbb70ceGthY4MYyWe38j3CVsKwB6X3ZAwG7wA3FPgIIvrc4Vzr+4GDHBay8e/wXbRB9DTvjlr
vAxq/zap3Iw+o+p+gTqkHNCx+LbhqAIiholx3NNdcwAWfwtPKkvnqlgxaBpwELMMD6Em9zd2MXNv
vDjC2mTwWIb5PTqCKnIibM7uKVUeT7fpAL6SaqAIc+shaoNBAKjcGwggaZG3v1Bhs5olSfUASZVZ
NK1EpymjypUSXAzMjHyzW0mKBIeUt15idcgpp9GzIh5u89OyU/1w9onNFKpEWdLxzrrNTsWZ6doU
eZZWiGxY9g+NmkSAjHFYR6kEnH6221LxlBHVl0PhscpALLevA+ys5txdOvn4zLi4fGYsYP+maMYP
VvJ0yFZFgvmTGmcnuB+bZftLZK9Zx7pSZydwqAWtFJZMrZv8zI7w3h1d8MEZg8Bz2xoELogD05QR
rK5JGT1D+EY/pcs+c0CqJ9midPUK3x+6z8sD86YvKTVYE4yIbjyhtgO5/ks7yFYZs8hmWhbuzJWn
XmtnU7lKMyShuMpr+8/Ia50mL/OL9zbGZqPK+oXREbc90SOHUc/Vezn06Wp+XZa4vQ7Bw9INU6C6
NyFlOpqKkQEVHl3mgKowAL8G8DdmAp56gb2idYKR4TdwWJA8yVS8YGcbHaA65QZJeI7pfYUGzA6i
qf3H8bemQz4xzsfKdksTkDNorvnPbKC+bISzc+WcDNYO8y6l31BhuMVvuv/bXEG/3puORxQVoqu6
h+D+Ua0tnclbHlw3Y+LhcHfH5WRKRPlljmLwjGkKLdIXNZoIH+oZERphTHTblzJJlHMELdA5pKoF
/x4MHStvTthNwEiVC15hrOdrQ48Si05ANyfjA49cag/BwAOraz8NsZ2qU5JuGITlDIbxxLmVTzN5
b/EjsllaDLQnzrsVN4ao32gfMwIEoX2APufbgoxZh10FD7el6dWsh62LvCVb6F5aENbcH3HGSQ31
BXpvMjQvSUfaHhTOLcxxbKjEXuYZanbOYyx0eu9eDuex64ZIfK139926m7nGyGhTbjqo5tT8sorT
gHBUlEhO3hcwWmut9u9AZtyD5527N/cBBsHrlIE2rH/JZ/qTLCoKWrH6DMirdNLwCY8NkNAXHokF
8jbHg6rMw5xiOLGN0YZ19JStYXtdPN+OP4x6cajoTVaj9FW0iKTPAeuIEiKWkmd88LtsRUqJOadZ
MbUMSJvieH2W4howga7O+XFM81fBnG+AYx1yVaue+frRJebyA5QQ2M5AtIynElwCqezscLZ23y28
4egNJzQVNXb7+9o83E6xbrS3Ru70bXr/I2nztLJlF9fu5jPP7FtZs8o0irx7TjnnsqRuy/W4GJAO
NjloN0uE0xEjzl7efIF5aXYfIa6ZjkbftiCsJUQa/XR56/7EB6Ga3r56Thx1799DKwB+Z79rCiZM
02xav+8Ncwvr/TiCnW0d0nOw2xfEGTR63HSuOkx2FtEfMtrBpC9pmzDMfO25l+HwhHWLQvBPWUIR
OvYM46qgYXDHO3/Lgux0hTHOgAgoS/oAHtaEftLxd8L9wemwL0jjxOXzY3Aj8yna7Yn+x2dJXfRk
6iZs8V9w6NqgvGAv0tL7bmQJGn61j3+MJmTZL/fl7dSVliBK2ZaOsU4+sqxkGmrJVleY1SJ8JT5O
lH2WJLCDug5LKSzpnowo/FVH5cJK/EYIpAidZLeZYrQh9COSpu1m3VfTMlwZdm6Bujyg1cC141v7
3z+9XPRvhMZrh4rwlMa6vH6dX7S9D80rDnb68iqzqCAkqUL5lYVTY90g0rMeoccIzMUjyMjr+66p
8RuNFrkxp1srr5emlKkn10ojmGmJq6uq9Sdr8piW+NRUp6Kv+dz9rIGEcqUEttMiHq9N54Qz6Pdk
Yp6i6shsIZmgxo6YeJ7UVM6dOM2BtkgLLXR8+4Y+0TXdxdgFg5BN5czVjVP59NtlntAhxIRFJNFY
9ovVIhr+1jpL6EWIWgqkEbdGrlDWdP3dO5G98kn3imwMDfC82XVqMAi9++1530Ia/0nEZT5JR/WN
TuWzedsk8SBW8mf6uHLomKl/VUmHHAKbbXHm6Cuy6TaLyFPsnFNo/mQUu452z2jWAw18kq6+FaN0
lkcJ5tyqSBvJkYMWu4+AFWiTPpiz044FDrDCCIlzNdigRzuYcCqWAMUOZj+rza0LXt1UaWe/XNgA
uUYgxWJo0hWI4pmLuI5dZIXLAlAsLEvHjYtBiK757rx79apXb7uOTbuz9/BNBFzsebmzuGerM7pj
F0sa6bcslcTz3cBoRohtDXpasrD3avGewjBiLD1pXF1oT/tkkiefE6Se+WFQEOAG3ptBTgFEH5pW
Rkzfu5GuDB66fwPmdHyzBkdikU6gWPlX8HaT6gLd+0XJzm1TtkcoR+2O6y+W69+EZyrfDoYN/jgt
GjzTT8l2uYTE2Xpr+pHoyzeUjHzyOtvcw6XyT1gKxSLfRYzeDpICbkBqAm1Jwx4T2VpPxBJZiSoF
scTYrw/pA7vzr7WIyOKgpbLqXMGaJW6MuEwsmx39klNk7kqgZPJEnIoCq9k+qbOl9hrTNjdT9k53
Vt+iliMYvizMN/v3bW5HSqX6XSADVJqJ1Vp24VnE4FGStRgItG2TrIS4jeq5U4tAYm+GpHrjynjW
GGS56QUpeliseoyLAQrA5F1hd4PhACgcTTKgBuDakDjofaI6G2VJy+jmz1eek2xaCokwCUHkY1Ce
vSL+vSjCiiuPC+kbu0wNyzrdEGJvVl1vNrUv9ejdgXjGbx2ppnPoqo3Dpyh6eYT6BfgMDKf7NrTb
92G/WdNfIRJgv9RyZ5+QDFPPdQ3uBWOG/Bo6uRHHk++KEeTlBFTz5G7kAi5/XdpNJSvILYnN6rdY
looFygR6LPmK+ulj7ZNPW92uLMwJcpzoG5VRVJl3I/tXfxe7QgtmiRLvJ31+dQ9n35OQFtLdL6NJ
ohVaFFxGT/BdqdLldCbHRNExkk8Eu4phb9A5R9we/aIL4V65UvWTOSdo66Z+8OAERyVQmKZxFla6
IX1UV5JB1Nd3serRm18f7iGB56j9nzbVFU6TutrYsB5xKH6O/+M8HKbbTx29UsV8f3fl3exa2QoH
mjDE+sig6SgY7gQ2E+lq15XodRj6dfmrIMS8O5mi6VFkFbdKNtCGGvnCkkJjzQHn/pDgziEoTVaA
+4rF/0bZE0uvv/2qy4pMzXL7WfpNEvhIt8B1RXyc7buDRhZak7haoL604fKWW0pDrgVL3Tpp1nb2
i1uJ9HNhFXp1PkF/1BvjEBbqse594BQdoeVd1PT18aT/kJ/yl7HFLWU4CorwwMKc5+KxmADqJn8o
pJkp1nqDXmEFiFxKppzRl3LeoQTFhBW3J5BaFJC9USnqaRZFpyJMrw/4uRay3V1uyiOmrh1ckawP
khfkZH74FfbUbaqNRQZQWuTb/GKLXlbcaZo6/Mt8ekSKKJo3siXEIpE34K3P7oR/qCZpiMLmaUDK
9VMhMsbvdJNMj9CuWlFgmGwF0G/MmcTvPOi7h4a6YlWYg8q4VGoNHxDo7mrsOWONyALqa3z8dj2b
VJIpLySfIcbp19Ulvx2+Ax8eB1ZFWnvmbPMbpYyezh4hluxnP6uBi5/6gC1P2nY8QVD05gZ4YLua
u1qa2kDqtvfOcp7pyO+6KjZXWJShgYQ4moqh5r/Zqs8HhHdkUpYUW6ZFI9Iv0ZDTdzwiImmf9KHE
mHSgzCYiEawaWJNMYvZpX6KExQ1ceWeekms0GxBBnwkxozXTghlWXBpHuZKOxzx06QVZY0G7O9LJ
sKbYsTAbvENR7a8tobsfJAsrbmVAi/2acAc8C51Us6CHz4NIuJW+wyYy+vca18lXsmINRPJnMlVW
hqGHWt6WttAQEXNOPo09zJxZC7+vOVIG+5qyFol4CgNhWsQhjpnoCKS1ruXQsbTmyZ8QBS7g4Qnx
tGfXDOvpOwaEY7P2zlLrWKCEjGz/mYaK3bWCTtB8mQIawhhxCABm2oerIFAqOOaY6HyuSYeifnjb
Z2lG42vI7A5G4seo9fb6XzCAM6/iWI1Z0vx3ACjKJiXvhvZZ9461c+CcOK89tApWPt3q7+86rF5l
tkieShqmr7is7phlPDhmwEpLSR1Rl4zeZieb+HojHIFqcZdyPApZNVhQvmh7oMyH42fgMAUttwey
RQ2Lo6xVTK231WuWoykpSrF8/cyS91ZeY1lmpWPq6u5L2+VojjKjKTvLuEC/vogijJkDffWXaSNY
yYG9mZ84rDAAM0UV1YYJWW/wUHz9RXs30w+0vS3oh+V/AK3bkPpRdmDc5B/yo5pcDOs8x6AWrhni
I+Jt7MBjuLP1YhK7b5tz5cGOE1+Ir17YlfzpgjSJrrIFFvns/Ra44cOF7BobAi9+mcf0lq7mN3mS
wwnkCpsdKJ28kxROYeilVIYRqYEDgXUvlBTApHm0TVfzoUajXOW77Gwecxnd11eULqawedXiUs7B
3oQ493y7Bk3eyKyg3o7AiHYJCC1RahmUMcfmb9jlwCviTW3/Usf6vFQsokEXjRiF13qXs3BCWmdF
cUtAVkykRz8DDyNXO+5k49Sakg7Ek01JuoD3AOIx9/jE1aBDs7YOr/t7fKlT8P2HIPqtmYCCJbEz
UMRz8qgr89pX2rMfe982L2m4OyO8eF/i6mBXcpZuVHJqK7qUxgpkYTeUzqCUPAD3Al7MOoWI7iTf
7SJSyzQMc+0wkjHXDz55Y3bQd5Ka4V5NQ7nU8JPF7Jf+jUur+PlKfEMxUf4O0dNx5xSHrpx2VYno
LVAxWUApO1Ac1h/HgCHSaTHuS42wJuQmhwTH+IgD4D871OIX4/L+P9DNszPEHEpxSn6FQddx9uvx
hIAW1AjggejIwsYzTcBirNKYnxPpAO+IZXVWtAyxmpheF3D3CZoZIYT0UvlA8j97bxBVghx79gJo
UcXdRR7X6s+dukl5LubvMST0pFJylT/cECgaVuZ2/H/AfidWkNTa3jg318C8TeMbg2hW7vhq9NW4
9iBqppZQvP062QKkf50AAUWRaMfE1R/1Lk9B4HYbpxnxLcvwAX8eA+M0r8HRculwIZd5LpxY7+rl
vq70ur03rLAaXKSKRenPtOQ0ijHj01K7+UyDqdtxfRpaLxKoNWSqiSbE2hS+MrYA5WxBv0/2Lewn
aOUftO+qsGTf00qnQtnFIUXRgTNSqMIbYFydwBcpGhnV88Hlbb1Nzx9ldxM6uIoL1JWkG3SQgvh+
3xnLfTG2JF9az7+hJFlbQnp1j+fmhT7UKXMw8ZEifOBrPPKtJumKjF+mUOJYCqK6NHncqJovbs5v
vvSFGFrZT7kdvbdNxw76f4ozoIAowpXsjNQwozXaL27aUWqRF/wNyYN99yU/lnX1H94jGJ3f4FIN
QABebFSdQKz6lMUzfKM7N+tos9CgBVZRS3Z5NlJSFwfdeE56ONXChFrgIzEa67hpYHGH0AKMLCd6
jv7st/GkbchjSLErPCyYEwkXg2DHvvDcx41/YrfuXahZbfs/8TNDZj+G2d/vfMRahIJngPmmHGig
AR+8Qvw0HKl+fzfkzMAdlMWZKDJyoD+9ouDlEtI9TAwADwzgBo71KgEJD0u6uxwioFy+9gzRs5xN
QsFGhS1JzUv9rR6wCo4hSdBS6pLpRcDOu+HVkXnuS+HNtNBlhD4oSTkEA/aelGSgsQPjP7Lv3392
GKPBWk/M1iuilm0qMk2O1mhBcplXhRW82OA6XaqAU7Qx2Z6rE1rjhhjXCU+JSX2qOyCE+UzJEH9T
DUS3ubTCAxXTRr7Rut1osTjJmqWm0A1nOD7rJnnjUSrCDo97PoEBX1aNY3zhUdrpQXN5s7OT2Y3A
u7zxv9kpkSTAGmrDuxiit7uhRKpBNaByhnl9GOsGHHgcZ0WisB7+Ia3nukIVHSIj6wcLidVn4aEo
BLmZQtLyLTo/5kvB0iggHUHcO8zuNFY6wHPBp7LiJuaMteipyuf1nIb5zqLaQmyQlAE8F+CjIBMD
KcwyC2s899BeQbvEgzfK5R2DazInibWijo2GkS7MVR4eDuEjOhJVpVwZ6vF2ogooj8c47klYkKer
/2Q0ERWz0UC/RkixN1HEkcLut462jKeczEqUJcQLMlHiIw2GMBsCRsOCMhNfeLQCXXSf3JCMhVvq
JbEzht2MIZZ+6nNyhDZ27NX8a72er3ikbMgJYOA1cir3xMSQVefi1FFM2TveoIZq2IeEt4Qna17C
z7GGlcR0H/8cbKtDCyYXZvdFMadgrQ0WUJ5QUXCk6SGWHk8rtXDa6WuTNqC7UjJSVZnvfQKWoBHc
hn6vnZWeIgl0OQDLZ3BJKkyMVPRNWLTieHK+jtFNkqkbcsHzbp76HLY3dFuis1twsxJC5zLGUlVE
XT6fPqVXNgSxl75We2hmsnPD5m9QlV+KORJ9GsTSqBnBEBToQyEJ9Y2qNVYuDZaGa4dtEwKXzwlM
mEwk3HPE9tdriRkVL/B2qD7y/wpQsu01GVe4EqQ8FQ2Mj07zIKHA5yQM/13BEDRtyFUEpQ0ely8/
eUQp0pKZBVStO1Di7sADEW4VfBZIJ7s6BGv9sr4ijRI4bMyR5av0cA5AadE/veIHVU/ipZslS6me
dNPEDnGHIQ016IyHRDCruBZTzeqfJQQcJnFSOtXUSpqeRuD5dT5cGqmyDSi7Z96HGhsjKCZZwoVw
IwXVe1+NtKdiC0UeYQkvjHlwYIt6r4zHhD72zQGMBAQ7ss+bFr1DZYp/WZA1OAZT/RR9xp2/TlxZ
aHBWYYCukuqfhCbpWNhn5/B7D2ZOm50uSsPwsqr++NvQdDAYTA8IGsjpnRlzYpa0F8ekS2Rdc0ly
yxVbK7gzXw327I2nLYaRliaPsgMgkImZUgGrtTwhlGMQAW++Dwk3mcF/F1skbWueXoVvSGdtVumC
6CJY7grGMp0FcdovIj1l33VNswN1JpvAGmvCF726WzuImZ0229rkTE+l50COA4lD01a3B7sbc/uu
LO0s50ATWZjCMqqptP/0ixvcc0pnwrcwAsLsVxp1hE6KvwFQJIyo+wAWb+Ev/HYmr45nkI5xduIT
HlPwDtXe4x4fWxsUCUgsaO/SpXoFsAZeIJaJ9HZOb4zhuf2E4z99RCICqxiLA3h2+7/LyVB/ewke
Y/pVKXThW/ojZroYrZy95D3QFCjuqj9alS/QFZ2V8dAYqs1D0OzThwfynw3k/bQnUg80Hp/q2nPy
ahWjOc6RydCwAXcTtCiKoTsz+O9EPdu0vyTBr49tt/7rL1r26vDAITIv2wUUxWXtdSGZo7rTPtTe
e0L9Gl9l1YsxjI0YHQycTo9R3QZgKPJUdVUU0C9WW8GvcOlo9pFnz+H3Nr2W2dqRwsC+BXTP8nBB
pseDidxZj+NOrFSLULbf/Spo1JGxqpdNVKMdothFPbji1JFfmHKPSq6EGDjb8nm3MHrJzaTcW+5d
tUDqwBoLzPcen6SPIB8ZmqMRoTK9ZTK6KzR7YTmHyjkkd/tRZ72zgVZGoXiXrL9NoNQPs5BH+Jbn
2aukFVwCIabnBd6PWhuzxZwbon02PF6RwTV3SlbL/3YWIIp40gp0DCMki8JXTxWnWLtKXw+Q/7k3
xbQE+Yr2YDTujQITlLcjXBXOO2mXbExYb65XxholYOL6mZaX5qTFxYCrGC/mt4IfCUSCPF8DdoAr
EezRPU8lKfnaB3RTdsuNFaYhDNpfxj4JfJXFkjNcT9Us1OojmLhfgvWWfSkFnUVHGkoekzOX4e6B
bxRuqbce+aqGlcBmPLdsfCc02/rv3u/GEM5bCL2lcNXUv21Qhj+BZFBJp0vb1OH30q+J6n5jwppd
Gy9OLdQwlR0+/UNYqc9eDRdM1yKNLaDxmMd/avRx8AGnkhN75C2EvTcmU4ac0gQ9cY/sXts9m7YK
PA3A4adIxwrm8TPG5Z29uZgQ7xvtN3G4ewCglwf10A63mQH4i2ZnXQ2Q8O1slk0upb43Irp3d6zL
LeyL3PxoAB/1FGjhXjE3iNgnv50RuA+H/EOSIiSCZ5HJDRxlPZ3D3xt2YB6so9cbR9D4gMfDHw33
clF+afcvQx36dMzNi7EmdMOPQdmzqDrtUESxXZUY8SIoDfCL7TyoJ8ijhSSTZnd9bzRxP2dkROJ2
8A5oexhOdu6HaaRbmM9QJtGn7DOe3+tJu+3Q8ydjBoPi1tpOT4GWeSSVrR03AEDbw4mGEribO+Z1
o6jXcmcPL/j4s2gHr99xPZqNCeeotyDxgVLxB9JUP/Mpes5PUfw0wgTnnXuecvLcX3O412CcdoAr
/e6RpcPK6CNl3szsAE46tDnP56qJwXeIdKpUfD2oBjiXmQ2ImDu4A0LuSAeb/HbeaJ453aOI46ms
Jy82K8LFxLSXXb5AayP3UIgPU2amgrZP8YhDofS3nn6LUj97Ji7IUnYCiYdnrL/o1pJTSiIb8lBN
1tEJe8PzanCnF6NqxQe0PZi9jUVfFXaxbVmTsU/SiRYIG74NT7NFgByj06VCgIlFDndAW7ImO++P
6eDIwPYX9Bo+C25+PtW1Varp9TaFr4WNvvFyVjipg9nyKpt36q+p/uKY7Vy+PX3MlBZavXAJxcck
cUoTBMWdAkN5nim4+Y8mjRojWDEpBDifgyZjXZrABxhop2hlPcjrsVSi0t0qI3W1uFUzn3zIaf5b
JYWnKeDvmcsmLxuvvpCKjZlLSMtUkQj7Cim7TwSPNkedGky0KhcjbvzRU5KwrUsuqUGR1aIWgxUm
4p5vobf+9gdiWWMUMsDcKRPiugtbwHWHnhYcYioEcODjiX8dASOBu3bdycMn6Ix3BTmmuTmmajlK
A9xTAjn0MjqiA/Wjn9mQCuNXHceuQEwVsCHZVNpoNmTv3xfZ+H2btLJ8YX/8kv1vaMuiAn6tbRjO
zRBOmBzsRKpEZoLd5jVHgaIebe8qb6b966gl1ws8u4Vx8AuZKjByqCN6qfGuTYehoUU/eIKZjry5
cxofaEXZwyraQ9gQW8P3v1cLey7O2ABaYtu+mCVdA+x04ZtAwcYxpjWG9ei5kc9PhMzUUyXu1Zkv
jIvVpXLR6Zu/dciV0B5kFm1M0DO8RoRk+t6Fb+/ERTwb2h0S8Zurcg1It1imoatElS2uCqxuNTYl
GWFtIRUxLZCsp5XH940SMepfwL5MOC+tmO31IvNS6XoKQCAmysIoBuLr1leMY78aOmlXpWLENi8W
OOss4xYN1j9HqvuQM6mKHS70hGeHmAEnoa1FxF4H+vz3oO9WDJNbfDifoMvK+E/pyn9+Tnpk/35E
mz/3SimexcMpHWAlmSloomSBWa4c2Tr/7qezkDjW/zdk4zsffPwp+6d1vs6UqADQ/vHnDSinE1WF
mQJj6WxiGxW50w44pezJrB7f/FKUryM7ApeEMCNFIimWhRULYy7hwe9GcbF1OnLtFO8K9OBOjpMN
7vC/860X2DTAJv9tXGjMzj6fDixPcgbZClbZoOb143JgSTKwctlFiO3mRpeSRFwS+WzzdcztGhxX
nz/DLczEFvS1yYqM94xyVBGBnGi2wWMhizvCF7Y3KcxDFLVyi6C5Cqmd0O00TnNy4o3yP9kSJV4/
PPNygd6jxwC5SP9pq3xsGxNsPN3/IGKQDKwueA3bjrKaBdYRkJtplfA4G0wW1K5ESuNrHlMxqirk
8991tf/uzg4zPHth7NGxWxyJLqyRMNRNpJS3lfPixweZA+ez1YO1uOQv/sx5YQPFItzxUjGtfQA4
7nJjHwP/W0wXSd6fx3BpdFje2pFwcPxkXHe+y6xnpXvLIi5R9rUzSKjWcT9ywFibzUT7t1ZedQXZ
DKz23oIzGEnSOkgVSUq1ATvfHKu11sgMhtNk+sALXmHQQeZQ4ecvvwrklUgbyM8rwiGc6naZUVzY
p1LSjDVl30SjSMW9kzWMAqKVgaCTmIcRh5P6ezPjhoR55MzsyeYQy4F47p2ugRxb1Hlc4jAXOd4R
It5BQ3HSpz2gwx5+KMZ20fBd2jHxpa5mmr59vZuWsuzbdkd8ruoRo5NkooBNOd70+nhNRo3ijeX6
exVedVDzxcEmHIZj1zm/Opd+P8SOi7cJFk+ntazfHrGzrEENkIVudVNKYhoL63xXo6csmXJ6E3aU
UQgKVdq7FN6+yGQUVu4UgVDNjF0Mc5pJZrIzQLbwIFdz5h5QiHjhhQu0WVHYKhsEZokdlGH5YMVW
y//Tlwu96FKaQn1rQFY6isHNE0aI4O9FhTsC19N29x7PmKXoyBtUFAHugBWBfQSkti0QD0/Vbz1q
picnwkGGQ7uRn5xKrsWw23ygVegOAwjtVm0Ynn+qN7myXbaYXgkU2G5gQRumm7cGQYpGvI/1Sgj5
MPzLhr6I4rjSsoSsZgXISzOfV4y2Id0jPou9bnL8DV1L0esMX246YzBSQWpCP4imgD6Hi10l0+92
F/aVn/VD8UfdEs3NTIB+hFWX2IcKGCL4bgZ9NjVmKhKmSf4Ers+b40bacuS0759zwWw7tMb0tCgJ
FRnNN2EHJyLLilLmerwb1fW0tCaoE9l8r0F+BD/h6FFm4HsxdaV9isCgXFcfnbngx2yE/Vj2cirB
0otETV0FyAHdnZKGkKqpsobJGcrszNaX93F8GIbBak0cQaACUYSZHZPFFCID5kPavu0OZ2fwC3iv
/1lJq89yMJAmJAkraXK8VHcO/izGfMxTky5Bi3BTfSfE3QBJ6HfVEclBSFV1I8OT5NZRR1FY1Cr0
dBS+8vbbQiM7/+JfmwW6pffvT7mycLF/cRgB/W1W1fq/4ASlmcNlGPEWA5vqavbR8ckSahkUIjSx
xtqKWitS3g3CBeH521SuiFSIvbzXep5VQUwRdjApt8QXhN3zNVARW10GIeceaTPasxBXiMAv+hjm
PTBXp4WD1GkoBJ9YtuB9aTuY3wm84g3QARQqV+f6PC/fOdcI+8KxN/zN6hpMdnPeNSUy1mj8YOOG
gcuGfYcgu4cazMK0Ae3MNUYsGITtT0AQ8LO+7zAmjJ88djVvIOSqJnd18gNyvFNHGrIqox0Dvycz
3YllEepyzww0IjQw09XwwmD/0r+ffs/Hok0vxFtVZCqgeT/PJdu1s7IFHxjamD287E5wqL1hysVJ
RBSVf7wdubMSG8nPiRsgjo3ylSvEuedpcxEDzJo5AQmpoRhlBCmD8PcQHqHMBawLfVekCYT6HQGg
2nkpalgr1dNL17MeOK4exh24KPhhZlg2lkrFo3PUJWLK+RdS8RWYySqsivg1myS8NLAB2r1EDPlZ
ZBeP56G6zmrACTy4Iz+GLn8BYZjqugwArpJgZUo0H7PkgdQNy5y0edUuCy4OHMIcIekn4DsGN7hp
ZlbZGQcWrI1LBRb0W+lZhQJ0D6vVRvdQjq/Yc+BhAe08VTuRcy30ToIYwEHK707KLQeZZG9QWtZc
tt4jpHDrAUex/gJqc+Y4GNuyo01K3/8vrr2OVLBzOg79rBZnJRLjvcELPF3Kj5R+sbbVX+qWmxM7
DPcotaVtzsUGv3+UAEJzHKetmwHzIBMR1vz1GnevFi3Z0M+KfItKK0ZBAORLs3tSI+RNUaBpqznh
pVBC6lebJcN5frg1+QPDVfBRiqw0+TKymQkrfMXEVHRdDKpQKi7m/0DPySkli4B/WFAkxzDzP0a9
qF7H45Xil4XEvAa+ULtoi+/N5aZw8revJh4jHph6TYht/NMozQUDVHBSLy7f/ivanxrnFMEeBc2H
ZXohuDTfmIPJTqrzYJfkRPiZLpry7ZG4CNL8nKtHiVkeQ1YzNi/Mrk4ube+EIW//gmzKRwfUDJsb
YvS7qA3t9mVKfat3hw1Cq/lXlNOQcfhjpMzhy3kW22LJBouWZG6BhOAv0Jq49rjXfvbc1FojZxRc
qurzcMLWDvJlMctDCtRoDYjG0WEsXfVBztN0O2caXCbivJarAHxU11mRhJr3cKxr2A9SC+E6l3N9
ZyiO0f9agFwSu4SezlIYdPLKmqKe4jw8dr1lU7M0UmkOJxWmYAO3e/5byDSseEsxjlUuSLRHj7Mp
inZPjbcYtJ06FiiHrySHcSNaPukT7JmblLqo9tEilqiSTxpmDr+TpMq7k4RKpXoVq/hPUbFmAFUT
nSe5BG3m5LjwIsLtkayq0+sPy8YWdFa9vVW0MaF0+QvKDegOVxBhSpOAga31kciZJTlV3tvX0vXF
vgZzCStRhqfYmnNcFxUySlTz9RG5xj8xMW1r8RyIKICTCfrZkXrcpPbJDsjov8qpeb7ufBvGP2uf
s8Dc9LHHr3UhXeFdzeIqfuf3jvEoKuW00Xcu+EqJKXx0jjW/nhQZdROG2CHH4YNJ9gTaSetoQNR5
m2b7QPRGxT4nm8eg0GaB2eOkfD4nP5elq89irMs6OJBtRi84Hrl8n3HfYc3va0Im8mw7seTi/c3j
+7cNZ6ihxMCm9c9wFQS95CFawr1ugVkUaB6Vyy/S1DO24NGFlWRFsAtwLylHLEHsAp2AHAdqMSwX
LolduTTfULPjIjP6p+VDHiERU6crtdMlDYHqVIf+dEYQl66oUWHbRMJDnogHjHyWg5YOHHmkFsVe
SK/XNp+SqDxzPLCwRtCGqI5LG0coOfNBYwn1F3cxCagr7ZNPGDPtPGdhCCmlcs4i/fNhV5qGKX4V
Kl5vVeztiT0zAFU4qt9ZBU5XADYlqHV/xksVdFcDMJuvKrvc0ZbgXl1ZO9jTMRpHf+TrvZBUEH5U
qwbsVNu+QzBrLK6/6ogJFHZESZgmG8dQrOFSy7i7hDO+cZXvzgpQva2wR3EYpXzGpDq2Q47B69vJ
di5O6EayHX2Ya7g0aNZoc3fETgVQOZ99oC1i8tA2SlrQd1sqSAjaXZcMkDfrJBA/XM0GGIVqCGTE
5snrW5EMrHpzuZZ0nSybpZXfQag/mTKylsY2yHJrnHEEOe/396WFMr4hvaPVII6IgrMkrABw1TLl
Sh91rmfGuyx7qEkAhRmjloN8fNadZT6EUIIYG1OGSbwse4YjTEu9oCbb3ElVHl78wKHYljUEVI6L
AeQ22QM5CTcl7vBccfIlVFlKFFWCdbe4GdWqOMFfTs6prvPdnqGGVNl8gxvWVXIEjBAyXmdDmX7E
uFGPrAFN47d28GVq1djH4sXgn/QnLTxvlYLyvPkgT9YscyjVvtq29YRn5FZh0H8g+nJSz4q3dvO3
RA8tFwRkFok9EWfXbjS4gN6aOC4RgNq0i5kNk6QbP0AIkhXzYgvJ3L+b9NPZB+ahxTK3YjWwjpAj
/kCkznxasJTCoB2NhPc3MEzjfijOoLg5g+r92iZDQYZgkYwAcxfdawozUH1mBQNm2RGZX9uOiqcs
zdaElz+t7/pNHRqLhqUUjNc/DE5RewQaBM//bscOMz9zdeD6TrOpNOIpdr9YSJDE6oF4Hpa4fYWv
G74ttxmnOoP0fZp04TaLWCwOBI8237TCqDM8qgLaskVmUJRVatKr9bDIdSMBid27/UWR6HNxVSaD
7+P8glTOYwE8EGBxU8oW1n7LJ/LqmkQl4U3ozOh++zUYqQlGAXAa5DLEPdJqPJpziZrJkWSkWi2s
FV2/Iz7LPalNm1ivLglLgmE0EwpRBe73Qbx5uT+TUWK/UhV80ZLcZj6hU2iYSGCqyVc0oI9AnR5d
CY0astWmdZnqUlRPnueqlTZLlUkGRo4ZE1Q7XKTGtNjzaz6Xh1VBgARQksbg4IFZsNH8B9MzDYJQ
5vA6qHg4fNtcQhlchYMUiZ66gIQePkK5fvQ/V/7fLanbb0taw7x6rBSy7pOqmK3FRkVi1W64tALd
pUdbF+HuVEetyoUOfjfGy/I85L3V5x9+eLLWjJMt3Sx54jiKgKGUkpkwJn/i3faKd7FZqdrnW7lT
YosiGWDrVhsn1BTIDLVtQ/H6TBuVfkiX4FSduA7CKCAr0GEs8CH1aCgQWLBbCh7YBMx4Z1Lli0DC
w8fU+woik6/AvbB26SMW65RquYVmeT+FDM9ZDzJWcbiKHA+HjaXD3y7obog2C5JN7pKvmLFatxze
kbagJRXO8SF/Ejl8jLLwxYh5IowSZScWLydtHOGknOUWIo6bsVbIDEUfdB6Cfud+9dNpGBMeVWZC
AK6/RXhv36rWuTXppFymNVA+iZf+KZJ8ZkpswBgccRaG5OXFJZCqEW1jmsl7LYdIybMwM85bNeyG
Gp/VT5O3hu9ZSlVXDgLKm30nj3IgM/ydKNR5M7euKtAHPpj6+f3eMtcbjnihUrBW/Shp+NjZLcOP
C7Qj6JzuI6zOfJE13dKbYH3blOhoRh2CifKYY56ILDPvdMQnRbdw/xVTymo3smtjTNqt/x4XVP7Z
ccSbhn65x7nevZDuzMN8V6T7vk0k1KxxekhjV2rpslb1c43TmG/5BTx3LqRl/BwmzwJdWrrFF6KA
lDgIp4ErN0eWG31mPRyv5kEk9lcTF+rC4ZtMI44/NqXWqWRFyGx/MTDAlKBRqWjpfB9RUXaIWZvW
inqI/zqccKHzTkhpogX3nFCaUT0qDtK3ysyIPHI5NSCKgi+EkrXqEO9cx8Rtr0joIB/l+Ke5xzeM
GMHRTtVcC1K8MQgSh+JKdAySA3cbHDYQhnS3aM3zrugnO9KQ0TtGDwBTpAlpdkHWQai/v3HgzzGr
p9ZK41Rx1u7S5cin9i2ouHf1QKKBp75Hf2hBNZr00PghmN+/8b5yyEl6dpQU6r1hmdj3DYBdeAvU
03G2RuCxt85XS5HdQl4yyIKzdJ3DhvM6h8UvIhBEtOa7GDY45X/n8xbZozpe2rmO+Yc4XkVgGu6d
kF+AqbWbrFVqM0mxHlLqa1fX5pSu/cu35YWQiK47g8N8SnqP1Fk31E7UIcepg/M1O9BmnkqEklXl
vXVm6BDgSrExxXdVAkNgHKxagaOwyqIJM4VNfovzeiaATpu9waIzf1s080idG7o8YstxWfP+YYoF
zPwtR5dnqsVBSHLg6H6l1Dp34cb/b6WivrCTR5/hiDN0Io3hjAwZqa7bEPONnqwvnp2gCxDkoBCd
Go7QoKxh2Ea6BBMoVcAHvOZnCHzFO726lMISzsSFxToyQPqzhUBJmJvuvUCRRNVzNAFkdAaib0h8
oiPbbWyWUsO/b0vC7MQjA7oMTRwte9MUAO+ft8sZW+vfto85tHQmUg+5kH3uDwTECy/Qc+GUbWc2
ms8VlzTyJeoEPGBqSyeaI0wdSgYvizTPbwt4vzeLld+iNNlbE5F55nFUw/ryjTcU3cjglh8APh7c
AWuzb+rHdCNEfRVp0r4zadXuCQvZxr37l0BhzjASxyrM7DHSDl2rQC53vuaSX/+CTOoWqKfrFtMQ
wMzroKaagNDqcei2joZ7MIvj5hn4O6zMvZhIBGcfd2qkCGY2wZs+89Ne4DG5yzxZNuH2KHhl2hn9
EcFdOG4ShSx2oeRZ1EDvZBo2nWFycmzsN1YoORoaPDOaShHzl77q6UfzRUsBkEUfZoW7mRM+KuDv
jmed7FBoGdVAL51DptEwnTyvRIPMtIvkykD8Wjg+Op1nZxzwBRT+p1xNM20QKf+/vRxFLX7GOgOI
+7/q2FJiIqS1DA0yEp5UNK0fWOsq0Mw3oFvCz/vePkoAlylwp2JbLlt4wMpglcz2k1hQ4/Yp/ABw
OS+4/Kds/ofI/wUq34mp0Ve73hTQDjk1cwi42vHbHlzXbjjwbatEJKIFyhTKcr40WcBzKD+NLU6L
pDkFPPyJbCWMsHRTRgvyWavJdfQXcFL1TVIvUmd9Q18WDRq2tb69G719aOcBGXRoxpfw3miwxQQF
29MHOfGEhbHPqYYZUbn6hITajlH2HbAzv8pGzlYSD9XJJzV0Ny//yWDKPei9YXH/JqtmhTjTCNbt
f3xCXeZ4iy6e2akjoAyaIkCTq1vNqiu7iBWCRSJuH5VBNvv/8xe6D5rq82ciqUgBcuF0L39nk8AY
2LWwSXlhCUptRrj8Wj/qRQ81UszBS3HYaJ2XTkObPJa8pWB5J1ZVCehm3noX9w8eubELvNcYJz7E
Vd73EpfRG52n1sAUgHqqpsQbIOYqrZPe67c8lL+9cG00+jClX2LTVWX/RScleFd0PMP651BteT4k
8BnVyEOLcMO0YZfZkH+KNoeRWwo9Ec2Srqfu7J0SIyePThKqvdWg6p/TDlosjWrFIEC1lgqIJEB9
fV4WWVzrdaR0PJKrqCK/A3jcjcBVbceuMhs7K9sWSPToE2B7Zz73afzPh6f0Pe0kfnfODzr9jvx1
D+CerPca0azRQakNRlqdxobMflrUSfXM16AEIKpq7RE4Fr2Ug39X8weyMdvlxi27cVDaF08m/Qfq
Hga9fbupchTxRw4vQykjqlhWQJiVPTG1aUxBJng03oAFcsCt0ufXfaR4Bv+LUvbleeuNXfvd/Bpq
eKLuWS5V2eouPQ3763orUWPpUCv1828Txw5yYXobAd4PG8RTavWKtuPa+VJcvAvJh5F4Hr6ZW13V
TAU2vW9ea7DTSb2FplxTVCI1LzdOcThMCvC0HBtpdk00neIlprlkdYl2kSyHHIhi2BUfRtTjiOKg
pfIrSVwnRYFkCReawomoKHscmd3kB0Y60Qo2mRu8f1C7mPwyld23XFvpOtchowXP6Wwd+XcL2gUe
NuYya3y8s5BFU4urSFikFlQtT7KA8OS57rDosZPsoLSfTnkBbkuPEzQDPnpz8/ZPTCC1iCI4WgAA
MetOu5zWmLQjWMxWyGLov6hgqV6e8umECurLyTgIEGLutRnnQEo5M744z/5aIykGLrvO8ymQYlKq
N7CZnSSNafmMW/cRZW6vBrFkJ3dzYNsQs/I/KWEne6xlhw4j/DKszRft9aur8xER7LQ+bjQPs+LI
iWkz8U8Qt+oMaqVtyBHRA+sj60IPWwjl/e8V7oowHcom25V7A9xyu4mDh5ayu4fq3XDsCfil3GIu
liDNqTVnoG5x2K2GPzUnIvAcNA/QQW5tj2hLsxCuq2KGbQPrnmepOWBe5vyrUHAdEcOJ9UA8j5aD
9aSsSWAsw2S7y6fnE3HAfglY/6mMEbc3XmDeeMk8Hl7OpkfBtEHpERsUTYgnnXP4hPddPPB7r/jL
26QH1uPIqXW68NtSY55PBty42ry1k4sVujuD9mz2V3DETaJIYue3OCZH2fsGzVz9gubuaIUyHb0q
8Qjr3x1rUYAhonoIsPvWKtYYluDY8zSTEgxX6moQai8riBmUo7x+6tG55nehrPSgGdo6GWa+X0er
nuWrE6bZs1mcHELaV8mc2DYX3N2Uht8v50BzQgitrFPkpNmeF2TxhkvwQupsjZQiIsE7o/H2Ge7/
1U9pSEYGfkSQRHPv6wJWFOE/of3TXE5OjyXyQUo6gY19i4qRl9akSS13fkWTrG8UH25ePE29LDyT
/RYUXK1iaOAuiW4kz0OZIGvXDgmLa5JglyaDSpXY0NhNNLYKbTvr9GUya3a+u4Ilqc/HUyQ7cCs0
w4lAZuo/NEnn7R4ecXjSH14x30g/RgzBtrtgT6YDkCVnJm+MG4jDLo9eDiH2spjOgqf5RtnAP5QE
Puu6zAn1XwITBcNJQo2nMVHGP/WoXxSPyzQuZXh2eDkm76/OAQkP8JdtZJHU9zz0OZEkkoZqd1mf
zUbeWAs5OlDFZ4YaDEYYabe6vT7afFyGS4k416hR2EGu5mSVaRnC37R7NalvbWCl7nKPrB+dcioy
e4+LGqcIfS16Gc4Bvx6OcvnhoAORalzpohaya4JM2WVytN8eSZSrGOgmWUvt3PAf6yKN5shv7/fB
osqtAXTiEiKtCM89UKReGzDnQJefvUk3NSMA4A7NSPCFOUuRwh3kiaBprhjCtCjFY799wjrU0YHj
h3esr8JNZcK2ZuzweKdvJG2PySi47E5puq/v4KzS0Cik7np9KWEwAoPM4mdOPoJmat1A5gDFBFmG
WYGqFnYvwOgHAB6LHmrogf3iFDWee3YJsUpSoS7bQ/xPHXLPFH6x3poqBupsR9kQsixGmOVdHuGz
zIuJ/bVJ+IYt2/8OnhAZvfVmYEISdHhJ6slcAisi1wDhzX82MyD6oRqvPF0VHPXA7KgwEQmhXXwi
5HpyicV3a2jrFaAEId1eoJ3gu5z2Rv+jE5dxvHJLi9v3G53aqU6Dveyk11a+ORdVuOuOlbDzdGdR
F2xybELYK/aVGh38Z2fD3N39hXXCLcTlcnxI9bzlSiHGKJPubzq1ta2VoUXDxaoyVMdG5WIpOKwl
8yPx1E55eQXRmuVveFaabHrd9RKYwagMLDSW3lIGVffOtBX7VOKPt4JOvabxlQneGSvwZ8K5UpXr
HnCJnx6cFKvDnSa2M64nWvBEuvW+WVJeJ4wG2d9W5cs9qQlAcRwaTQVRS0wbktDg/BjNrrGHsDOw
nmB5x03qqlDPdZv3+QhIeyad87I52hAKGyh5/PLUrqmWKoe3ix71WZ4TBS4gvleuxEKrIadax16u
xpbB47MXtGrPQNZVmkALVS9wbqR7KHVYoSW3E3vXM9CgXJ5cJ16PfkMJe+Day4NOGwnv5TelYyVP
h82CbYNMAy8MsOn1DCyBhdBMRCBIHNha70eM783sPZgATbMLcsdCoUlv/8loyUJaMO3BrwruC3/4
yV6YX8V8HS0l37G581w9sF3l8XYAl14dQtuu8GvklRJQe5VhG6axi5vJsTx05Uz92Idoa0Ljmyys
u3oKdTJjd7PEveUuVPxTnTTVzSqYHZzathIoj+gHb3HLuUU0VUCVWEINbNDSvVGpBV47kBN1QQoa
YIYEKojJ6WNUhLtAkVzAanOzlFGy5FfRvOlkTxwMXbanqmTqAiLZ6Mux4JboDOWSPsHIH+AR7oL3
AxJ6Mbkfn21HlMvn+j1EMofRC209OBaJyvpwR4LtMqHLpSAMIwalFagbTqK/RWRE9RkrU59/an1M
qO3zh5sPOI/CCWaIyWTRpgKlaBc9ZTEGlBhEZ8GkPN6xz9aL8WJCzTegzg5atuq1qYoK58OXYxEE
T30SKiZQIVCMY6ZOd8o54MjDRvTnOdWa1YVYeED33wJEn/gPeyWcw6YP8E70rlTvVoFlhkVRm39k
68SFuGXOApZKzZwLdSiHhN3iIbjA6Fvzx3rtGt6Zetiwob951qIgg+HRw6EtMVy2NVlGVh8gDf5G
1QJj3WM2djHBIpes9ekFzIsI7Is+UvRaJQDiAV/oeLDolBrVenPwYXJ8AZMzz9kPDDHa8tUe9XhW
SnP9fyjKG8ejWr0ZRHzjMal3vMzm2brrLybx2CLCT2m8d3GtoYTwDBxlWPGBHvHZdBxOXgV7tvCM
+8y7N4annz0o86TG6Ewjz7SxHWNV9kqJSBPnHtdauLBdkpcw/srHqKFVA5CdBPIz+Uov41x9p3F5
g36dVvCs7tHeT6VkUOF2FoKzTQgmI6SNuxajuSWGKAqXo0TrU1mJa+kDoVeHFDSm/W7VitV1cx5D
RfGKMTXTJrWyotJaA1D2r++Yh1BbfyTlf2EovBblvX1f2zkKDKRHPhX5qZ753JQ4VEYeLU1ec2k/
Tb/ifEHwm1iivHZNLFIIHhnrKWvOxc54PH30S07oTl85k247M7r09BOxFucvVeADxC4/Igjd/Z95
ES8XEekOpVcz3KrItpEwyBS/sb1mrShmTzUrIo4PkYSNpk9B+mYtyDqSANR/bjF9OWFHxJ7MsFjs
MJExBFcItjOBBB2EF2hKWBe+ziISs1j26CbXaymIel1FNgpisyRGsGyGC3E2oHXiwAFHg3FpGCSE
56aHT+dBt4g4eOSo1RsOzW+qB8WwK04rpx0isWqzN1lv06ny0C2B52Oxxd1rn2+hwx2qaTQi2jSv
/4A9pQda15x5k1Ehk5B+aJoQOWclWmsP7Y2lHXsQkgbppAJdXepO/54Oc1bha35Y3lwNkd19T9Uu
Woy8NetKc+8GfbtxjdloZeE8ov8FbuTA1WLmRqI+LYa8o6OhdnWiIEYys8KrPF/1RzovSiOS0V//
7RVFhymupFTMUJZJ0wxFhzXvwD8NuAN+2JPuazqEbiE5coT1azzoLoviQXULvvRYpCGa2dWHqIAu
rxCX7K28Vsscy+A7SXKnhsddp5rOyco+GjDxFEcCFegUvxpH+GoyErSA4iEMwTpWZRQeyFB8PQr8
z6alXlbq9QF51k9EaUHR4WUc31Why9qrecp1VTx31sqG58ofKFxYpxkU1Tq1l2PqbVFsW2ib8nxg
mqQfD6eTgN1OyM+2keAmRDavO1trkpje4qA2ZZ+pGfLuD5jQVdov8H9vYd3wFGIu6PbWRY6mus0M
MhxUr4xN6N1b4iXMuhQ4Ve/e8g3lNGab+wriNnDdcgpiXTDWtSaJLwlwPSh9ZWi+zmIuBQ56SN4G
tVuKcpCu1wn1irFhlj8qUhXC+mBl0qhb6/n5xjlI7ONdom3dATIvY1eMhBVlyrwO8v8j4T638MBa
WK2hhseg77zot/lePcnsMe2ONhw+qH1b5wHhp7rU0DpSWIb5LXp6xbSAGolDSEv8Lgg6m7sapLGO
AzECD+buyDPfDG9WicHWSz5pPKb31pTl9CoN00Lm2Ys+c0QnoUkCsUVie5sMJzdD1XJS1GHLXzga
VgHXqSX+KUnuXP5t3T13alGZNXaZ+r+8DHd360Mzd8muNkarXC3MEqkw09z/muLXOJMawzx0A3jF
TpepdOVqxGqareht++q3IutpOxN/e6wnHXdPpqJfernL+cstXbWwjgKq6lkKIOo1OM3BFnbhN0Yw
iLaHNShoCAqTkRNOGwSWeP8JHVaqh8j68K/Furg0ELy0ZvrrllliV5/jYYn0pbXek8/Tap/k/dCk
X49d+wi+A3I9aT41I/hQe5nS0CUY1CBvMWAIl2SKgmJz7IwiFqHSgbASOREsq1e3i6fFYvbcTNJY
IUC0pos5kZdUlKBIB+URg2hOdKVIsmxklr/8iRhU2lAQDL5qiobyGE1+85MR0l3RATOl3ZOd2DOn
7I1tk48rmSwJ+vdVpP5WenOqW/vvcKBKkfnzzoWiJYapvdy7CNkZ52ffHJr6sK06meH/db4URYA0
JGytcROL5KcMo0KLe3gawU3OPF3YuUV8AFsapBsrxauLI56U3dcIAUz8PRCQGItZ0U3qlyqJTPE7
OjSJWbOcBI1UD30GHravY6RxBAoCs+/vYXo9OYP4B38CC0j8yGLex+jyItmW0su6Ic547oEphFIM
32EtJ6x/gprJ8BBzVMlO3KT4cV7wlHQXlQJnLSwWZUFfLorR3dcsysYNLdig3kB4sy2yD+reYeu9
NyykCi1ef8pPjEG9Anr6F8u+hM1FqeFbr1XycTn50qeAdCD/KWYtgVfk+Na4R4/01eRIQMWe3+J3
PIWFdeqDpafe5DcjR1G0123610GvRfSo2fh1tMEUuF3Fu8w0ZDxd2s8Nxx4zsGLWksitt/nSXyQS
62n7FMzVENRsaqvDsRRBxFF2OL53Q+VljC5c2TEJeHt6pBSY1p5N9s9u6jyro1Bhg8yO7u8GhaFl
0JyDGXgP+uLRgm9gtyvH75/igiL2o+NCE2Q0ilod6MbUSnnWr0X9VwyDmYNwgl6eZ/IieIYKFPf1
qFT5mbWexSCxZrI1KCkZDv+6qQjsFtJJy+8BP8sdQR458PWqGpK7aoDSgd7KWZm2apaRWMIM5tPm
KQz+a4KUkXQKv34DinxgBOeCWbqXUQYbXrA+UBKiE8x6DFNrvRonLahjmsM3+R8ymA0Rtk+4AVMA
M/O4+HVx0iH8n+R5MAiUhttzvyfNG1o2pegifN/veW/A3pULxvSxXTq49KORD1TFbE0eUutWPUIo
qHnhtzWcMiEGaAuQFoROcI6lQm1MuzQUm2NKlbcHj6OEgeNhuC1uVCaj3/YVEpVoKRtTWr684CQR
YK4ioVVRjZkpSZEcyBysC6iBXAuNUO7EZ86SWom7OAf7ghFeyMOk/7lx42yd1gMqRqvg8I769AHx
svZu5jUIVzHn3/GiiL9m821dD4HgPQ2ug4CW751zHRWYWURZO7ZT2CcrTI9RBXU4+ke+OeEe/ULs
Xd4vxw32v0yHzAvvcjKxm5GaopF0zI/0r2h0IcdzDMyrZOPp2bCJMKLuf3pa9t/QTkjz01Zv/sbO
KsKBhwr2Qy1QYDuRMZKy0JEMjG3zt7SwXHXJndCzfj+OdDfoSEdmm/dxiR0hSA7i61upYF2IocCT
4HL3yVoBDKar3M790b+zM8xlhnrAoZvgJa8ptGh3GCyS7zmWBCgycwzZcXn6J9FxY1Stsxk9jnZV
VvoObmk0c0Gf5rCmupYIrtfJDEmApDLgNHOMBAAmJxlxd5imdpcwmY98E+b/FSXMpKYfHiS07wnR
4/KBw4fhyRZTnx0Kh+RapDj8C2K92nm+Y6xKJZQLcf6Qnc53vyzyXI/jCEnFPpC3kzWBdF8OBn5I
vPkyAwXO94yBThO/L+DhqVmAcaPqgymUghu2UWMxOrpoT43Wg6fLsLv5G1nUqFSI+NZ4kY7G0Hjv
qWcO/FsDJWTBo+B6gHr0GAd368vPX0lR885BY+nrylH1twDDyaq7ZAqcTvLKtNLg3/FvwfJe39Gx
9YGyg8LNxgHdoqdLcthOUoGu1b+/4QYS3scW4cOobwRh3t0z3/R3f7hRaVz4t4Je5RdfZa2awLTs
+X+ChIdM8b7sAp3UBzxDhnG8ynwCH0cYfUyvqEenhOKyvbjYw/odpcc9GCTH8UHWAn6VzNh47NRy
ZzlE3T6MaIwx2JpvbHHbbQGnaQ2rpTY6plJv4pa0VXdnEca28zOFspW7SURhxPuRzc4f0XFJl2Du
8qZuG3xYwoQLSMgp+X1oRkjjycfkjWsg5LdWZiGPKExD637AXXlzvIFyZtulmfLiEj4jy34coHr5
DQxAxYiB2ZGSd/X8LqmJqmXT4xC5RGRptynKRp0Rt3o22yXr9KUl4Dbf9P856Tr8a5QtFHGa2f7W
EI7KSpUfJ3hOHojf4/Pd572I/9m7AVF7MoYwM4Pgoq39gSIpbQ/CgO08od74iwKx4ZYYr74Eu/ZI
oRS4EPR1ChN2rWZPM+HW+XLhQmKNLJnN8cJLmWWMVpGIBbw59sPvlnz2sI5vhrDgp5umoYpzgcUa
e0dp5si4l/GuY/75A3uqUIIvW+9Em2X0bqTdLRxT8zzDws+eDZCL4hajJub2DrHpN/bqUbP/ReYc
T8yNwd751cJhkZPRdue70vovfHoT8qdVsiG34vDkP/Prwy039t1/cXu7DUCvVw3xwIy0sWPKFYBv
mtJM6wsK5PkQDiyBG4YS3HyoZcHA9z2bUgf8qSi2yo0/n+L6MlrxF/k7qCXly5AcawffVIuB6ZWw
YEkOVB2CYGXQ/LBvHllQEf+Cf0CbCkWp8REE6vqeKatjz5A/cPV3jwCa6M47+v5+Cbc4QkhiHiT+
YkppE5yoOsj2BvY3ZET45w2uXtkFLX+y7+qIy+1VZPd9q+Q2NgV2v6NMCwsWX8y+lnPVYUytjK2U
Lv/lTQRJ7Ph1TAxOmsU/sA5emzqOLm3CueI4rh1QZAv7sgTDut5MtfHWHILKTKSGSIKmMYrO/spG
5W/xunoGN2vJWSDCyp10W3UNGib9EuJgQD076lVIo8etrhDpQrPMr3hJCUVXdhHELbpRTVQp6Tl/
dorj/XImD8PPxIva6LOX3nfLbnL0DXX3i55pjwoW+ek0leJPt3yxDu4ctGPh/zgaXWePgIsSF2rD
EZ9LEd9aeTzBM6M/NoGBHWCIF93qedC1SIZ7cPfI9tAQ8Er5rjQ0GQJPgQLcr8qebxPSARMzgaaO
ZQZ5O4N7TBicI5qjY1wiGmCVnsNFHANn/yiv/bzKz8Q8m4UvvKdi2KhUGZncXVBxxAP0siZkH80A
UHH32WfDY8Ieyfenp6fBWAQtqsMM+nbl3CMefO6q8cAXHdTn/SYUrIqX3wz0yuZAO9gBbhxNDdlZ
sKOpjpbVkoE2fCa2Gh0uszqng++Mq+0tUAg09dNp90jKu+9EuUfkedk2FyyDSa9to9VxCoAgKais
Fv0gHc60lo6+bcIEY9npE6NR8pF3JX+rzO1SRLyY2/HJH22Gy3BpaNMJTckGHjB8TLaDHIbrbMXm
9+Lvc1VO78/U1Zoz168HE4uB4x95ZDyX9A1cHWBdDS0bl3Pv9BRthMH0dpXZvA6p0Cdk0kPL83mj
o9GdwsxYsE2DuIc+cmyIXxGzaRflyBBrvPmC9/cLzTTiPODGrs6wqgGTsH34FcLo5B0OCC5819r0
9ghg9uRvxq3cxwBnbPPymz9fVTYrjIoh4vOKnTrUyLCxoxy/wuUkJwcZcjcgviTE39XPiTgD5+wp
oYr8OE+KJ1MUe7raZ+STfORNCbUXSr0KSqyK0o9W8nfO+hNq8XSCJtSlpquyXc/JKPtN+mfaydjf
nQT6uXJucufvihSJdltgSiWYJCO1aczElkHTMn32z+D6YrdrrNaVBYQ2tJC6p7lC92j6UEQZgKtK
MNKNL7WK8zUmX1ejSUg8ge0Bg20zL/2aXud8knRZCMQkvzG5ghga22uBtP1y2nbA8BvMRLio/SOo
MKgDFbDW+7+6wW2g/elZ0FVLHR7Zbt9IPHQoy5E13mHc2Fb2OHwP4TJ+yta6ahFXXP0m2RCwFx/S
17XiBQuMOQbE/O5gBILxUuRtUFLWiOk6Jz8UQoKGhiDuehYlGVQ48CgqzH0eKOBMIqX+XfEDf/p/
uUHBRO12cQ+Mb1ia7XID9Cq962kR5UBt6iuqvRo/i7VZq7UQmG5mzmjNb7LGF/XaphevzKfN6woj
tE1vWQlLuIxWigP/NrbDl9g5voxqvilCJFa94uqirTfkNJhnryHwCUADVLLD0IPH0pbF37gimDMq
f3xsRoFfrIrcj122BJ5LvJ4/Dgt8emip3hpF8f5A0IgCC/Sl8iGLCiz7v0W9Y+5kGCwmwHo/GKXm
oGxjUhZX6J9ByGEBA2Y2mxcTOkewMpuFOTfiGt6N5zNOrnwY5gYxoJpM+rmltXn2S2eWnQ1ITfR3
hgO4AfO8SVcchTdGj6tAHNmGBqXoqsj7bL8f3oMAHV9+E3ufTd06t9sJ93l1zTrG4LKYaUptieeQ
hbnYl8Bk5Hnbtl5STfTGx7Arqlk5mA2FHMK90n0r0sQYzWhbKhnd2gEVJJVpaOaD2w488ZXwXO4W
0N43jLATmCC7oSemj/Jbp4W84qRipyLmC35zJIDZ1Vfwj1MxsF1/AalwVB6n6YUwU6iPwb72xjYv
8EDgFFzYKDE08hWfDiX/RStm9oBYzOPWRpb6c5yEqYsGaClHs8nUDGx/L55kKi6yajvLaRLvIHwn
emPLmH3fOPdBtNuVT10ITBSK5Pidkem+IL4u0yb4VCd9eVJU9Ccd1yygCNtAgLlS+akFzIwIOByD
0vdp20Y4/lT6OGDLOv8/zcMdCU/n1awhy42v2Z5M4cGVwH/cO9+f4W+ZE1IDtTZhD/zyHUrVOya2
j99kuIbXe4FxFV0sg1XVDBKCeO9mzK4OYABKKXFIjjbgrtAWTLKkNQCL67iKGOme06zh15R9Mo9F
rVAEx0pdhn8gTgJgJFWD0JA4A8uXDfY6DNwLXb9pxTTi/xpLkOsrnD313lVVzG3bgkr1Yq2smxja
p7ReGTT7m7sv31CNN6NZEvEWxjJObhzhaAzhN/OGh9f5V6wMIFHBmDOLAAJB27iIJ3V7sEdfBEKf
ZfHvXNzYIkIBMlFy+Y/6TvrQJvic2rSbSSl8ELnqGCPJirtNgEEstiGi2nBkQUVvgxvVSop3/afA
jIv8XslFzzKU9q+S5tN9TVPQDTEb9hgusAqKIFzss2H21WPvHSlwxx43Tl6LSRJTdd1k+wdr13UH
/Mp2L4WwuvaHAN9VhroHMNTyAlsClmAkDPu74TTL70zfqhhe2xIoOciBrmw1AozNS2B5Ti01Dkbm
qpbQd8JXnBNjYTugRvO+7TBoc2SiS0JJcWMir5Hk04ALCR69ZFKiIphKn2y3fpW2XQghhOs4jYV4
qEM+2VfBry/YZrvNdYdB3R+CrsjZ8CMq2sjLEYjE+57CLGrweLTdmttYTXNmmCMfv+9weS9OpQVT
u55gOElTK/VoPvMCNV9+cLg05A+tr7WO8rXC1JNEkdD9h9N79sGFIAd8NpX+ijAVPQgBCO6E2LjA
VRP+8FY8TVViR7iGFmFLz3TLUhOlHCAKsATWiuMdj+sPeyorasAkqEZWzCI3DEA8vqQMhebxHR1q
zjqjmsAhZ0lHII+fSjTCRCWdYyVSgpU3HCi9AJLVK0CZrlxWnV5Rbfjoc9NQxV6P+YcCRz4AA0NJ
UWHNfB1c7sZIugfVF+6E//EqaUce2LeKEzaZrJrj2P09gkL2XkqJYCdEjwb7tuV3MbnZEl6zrhxV
CpIuoGZZDAAVeS6+IMigusNVplPfy6SK5Zcj2ALYgOQ928MlhSDLGZ7DYxsZKkgcODlY/Sw6FUv0
xquX3KoN3ajTbCuzTj1CHcGJpwrzjqblfioimvNLWSp6x0sgn6VNGRkg6vntqM5Nc7jFdEWlW82I
FeBusRXtp1S8cniLwLn4bjiEALR3UzKQclVH1qnhFUi45VqAyKaUMGqbTG24KF14TkNH9Jet0JRP
5WJAl+2WI+XflozhNQ+OIsErWshi5tVxWTkVqQBpzBt0/iL2RfiD7xyThyKBi5O/8t74NZ6JGddp
zqAA5zKRabQrTfHzL/a1WWTDCYw8vjopfzC7olxuQPx408cQHqlsjlS81sVGylVwc1X7D4cn+Tpb
Jn7XnIbZnakprNclQdd+r4esNNEfqu8LTQBvUjJM5MEIKunFW6I+R+uQ2SHMH0obxTWJwSfk0rQF
xUUkHG+MZJFTT3XyLoQ4kf8u6uNZcrl4/M0MsNnapRyC6mgBNA9Z69a+7A7JyibTLXozDsxZ5Rts
SneHPiHWQuuRLR2VfQGQZd64EbYQBa+GtXOG1/bFoLYFVjhmzlAOmiNvg0YRKPsxydNyY835KiUq
cPGzi3WnP7s9pMn/bKBU6h2M7f75J0PXt2ftxs6Q9l2aPDjCE6ru+sbc6Wm1R1E/wf5eTLAPbn7u
1ZCy+UE4IsQumAy+hQxZNo8GIa1NXKPJdNdG+g7AQkSSo1G1ErPZdIg2PknjSv7VaC1HQa040y4O
h39ix9rfqr3q0aOlY1DBOyipG5Q01uc8zegjbX9egx54d9VJN58dBMVZJNijAIWa5eEU1IaOkKV1
kExVfkrkwNEVPBjEqyhauV0VO3QdaKwTMIH35SIRKKsWWzxI3XcYB9cFTzv+2DxI4riS9/6x1fd6
uVDGLSGfBiBcj5eIemsyKnAoxnpT9lAhcLmbkf1gHfpGahEtU4qSjdhooAU28qvU6V+Kgbv/F4lG
6Gvs2r83ZK1UZXSCKi5GjP4V7u4jCixzKYLrHDDdIFIV3WVfmnXWd7K2qDAVT7bq4D0JQKyYDPT6
BH7gvl+LX3vfYpdeuDyEpRMSR4rwWC/3xJ15Mi/N49QB9egrxRlRYvc2w5ApxukZ1DzDvsh+5Dda
Jva2/v7eezE+BZlg7kx+7lkTsa2nPUTOybVX9JYzcJFpqpzGyFMwGliJTOQT5wBfb8dJREkF5xfG
FRjYulatg3aQlMxGk+bmKrCwsqqUdsHGPgkLTEtJ5g+MkWEJG4Co0vAbV5ICyHugG0SJ1WW1NE8+
slZSGYQWwV5BDUWXCQOKUyYIteeTfm8E49YLgT2ZJbHge//oVWRGUY7r/uDoN1Saq0wc4RN6RLDM
QuRMOvEdWLN4N92PYoA8coGOt1TsHxt4Dzdf2dOtukNVT7TiYnNLxZxMCdVxis5fSNp5QmwCPluv
FdBTb+dQF0B7N+xAhZ41xcUG6f5eePtfF2EkUVckD4Jc3nzm+n+XQej1Ye8XPM5aQYf1s/L1GtMy
8Ioh8ppMLpBDmA0XvKEJ57/X5bvXo89xe6/SS/wylUudT7KnAWM6wxRdEvUpMdRVxsriYidIC1fV
kS34CiBOZ4XMmkxR/HWcxrRdhzr4iCizRSLxLhhnseGx6u52d6f+k0g+gDT0Gak85fuZHtFAzkev
WLwU896fqozo/BX0l8PspXxcoEHlob/lJqSpfLFyMWTMOY3IT0GgLe4+MoiWgBd1QBxC5JEsEXu1
tOseH7/IdwO4JdA/kLaqWJ+SSF6/rAUC4b++22Xr2rOT2+1hy+rNrHxJ6ga/Jm5SgbQVFdIB+GU5
mJVUFEGn0I2So1rpZq6osjwxsHkh+aoKKvLELxu2qTCaCtfZtXTd0fT2QhJDiNkDh96RvJF6YByn
NexxmtllLbIBItEZU5z3zyAD/5wc8t6h5IQtWgTHr/KKWdwKA9Klz3nyyhu0BZuwUCZr2Ad1hyow
687IiI6XdjgQDMLfM/OfH50fCTmD+ryITXaLVn+27dNHyv8LpKWjmtNqb0qsDB14gQcTnHP30MiJ
OaVfNKP0lBjsbT/2TsmmTak2CAIEDHmF9SRtijr+7SlcBkyIofWb75x7HoD0hQohaTDTZ4XTQOHd
wMvXUX+zzZ0IfQ/ZC5F13mrE6k3afBfPkkfiwiYJZYMid134fZSYV/yATnGWRKHUBZ/sMJKDpmVP
dr7UbwZVDIBczQSr15klFnnaTcMNybvk6dDdk8Ct7ACRrIoehugVuiQ9ru/VlCMwkGJ8H/trmhxx
QASPSFdJ3Y2lmfukuipt/O+exqpdG26bfECo8vzhBsSo8QyIRt/nwC4to4GTg8cMTlZOQDZg9WCf
/RyfGbw1ix/ZjP8/axJQqW3aWQYsT82JASKO7Tyt7tAsRviUe40+RTWtnGfW16XjQwq+LS6UU6m2
sbTmK+mUJ8JvPMt8pl9CXAxXA/s0rIcriBwYAUFRZncgpHbscZTd4gemEhcgSvdAuyyOJwmcSufm
1ldO7s1dzLIfbC0ehaWeMNteo/Rou8/KDvEEvq9nTxY0qL77DcuNvxCFENQyxbC9EinBujs7JYPU
S51++gzbvhJGxCD1cZtSYokingigOzPKaO7Ax14i8bsb//tZbKvzp7xgItMnornWxuVXaO57HgZo
+6hBY+/rZ2Z7opBxVfo8Y2FH7xTAFO5C4ZDAbmBIgXxjCRxmB7APpBnUJu4Oq+0+PJlWW1m2+wA6
o5zU91UcRIrdG+vv9HzZGp7UTgF8LtTheBXBAZjqdJl5uHLUJaKtjF875J9fE6/3lA+1cRdmGXo+
8iPBqWvnjBgrtiOErFnYa+CIUy1diOiZcskVB/9kgpGmwr1n9wCvQpXDG8uqtdCWogEGeuEjbOHn
4PItnQj29ZpqLFL3c0axFNpw2v7Q7wz9xmUaV/l5QED3vxX2+TFEs9V69RrUNRt+naV2KC1bWMDy
o5mRcmCAJQjEANigWuzLqP/j/U8lZrr65BA8YlCzcQ4HMhBkT90r+anyN49RAzJ41gThpKrunMis
w2QDK02nwBXm9y4dG9d4jKFa14QvkBFO4hr/WLwlHq39/z0VwOX3uFeqCUvrn24xzxAH+O7s+ETW
M8U7hcopfEu0IovK1kQVQaRRTdylNu8iR7SMtF8n13xLQ3FBI6xo7qs56ccyV/xx5x1Gf3aQQAHw
erFYmEJIk6dOcc2b8GqSOCOt/13l46mtdERwwF8p1jQJbvdlJtWH3+JzkkU04XFmTrTMxgu8ZEW5
35AL3prJrD0e0Sr2euX+HBsqo3GikgfyS39KmSfCs7VW+QY1VqtsMjjLx+b2Ls6kKNlhST0SEIgd
IPuQPQdt9TpAweTS5hhEi4YWmsmPe0M3ckVCp5e/9MD0QizzNVx3SgFCdLNh5AO6etT8DkcqdJ49
N/olEWa8QUVCJlvwn3SooeUCjpx+lEvgD7Lkzjwq8jLDtGAJgnvvH7A+mUVafB/pjWXft8yaJZCq
E087MWRaHSOwYj23CCLf9rUyvSjd4ecpFOIxzWGGZ8RnzpgwM+feIYZxHJ+fDFQBa+yF71bEwn/R
sP+3UycprVaxHaTxoKfdUtHzO/OCB4zHccSOn3fpD0fAsUutLdNgIUWTAjjJxpVFnzEvIbS1enDg
N1/PrrHZ43xJLSPaUI8+/Qwo+fPu84QppZwODPvFCwrUleD8yypeffZX9KOxsEIOgO8vwoXlnkyg
lev4xbvJo+00c8REHvS047bYVxoLv6DhVBp/+8kwJHcu6HjoYBCRDRbqHUjYbe+OItUNi7I2yn3l
dtVrCXX4Xodt3nuaGTauMnr9VGDFGlvjmZnT3MUpMgH8PrfHqKmi0jZvGfqfjw8jGZwzt759Lmtv
0eBz1kkw4UmedEJkOAvHi160Cv09PIludx5B41o4BLZG9yNje0XGyWgzW6Ejo6njyFB2vGEMlObM
WtDPPUTQu+zvlDJ6ZLH0995pBe0tA1+3tf6DSXHxyOzvZz6N8Kp8GL1VW+4rO63bMr9hOUFHLXBm
2Da6maZ92VAQ9lZnsbNNJgyAy/++eSf8IdinnZii8ffmHo1JSTR52CDgD2Z20+L8Q854V2xau2IJ
InGFbHUGSn6e4+auomrWIlfY/BEAc9g5zPzlYh5x+4g72ADjwDmA5R4btPFNYIT2hggiYOfjQrPB
rAg4MHCXa0N7WN+zWSf+0dGSmVA0JY38S4lid9bx1lzf/NHazvfOKnXwUV3hQh01OV6NaZhnHu6O
OSVKNI8Ic3ZQ8eDo6id34kHjjsjtM82dJrurU7j+GLctbvUVr8iYFZ8UxDLbwd7ml9jaefI98b9r
5xwisRgb7ZbwSFvSbjFLm0Q9UZcIVwib/Jt+KtIx10T5Ngup50SP4z0uqjPkn65ULx8qpU/+GH4+
iwXbdPWi74phbjGQMil58wBPyyhdhXPAmJNzbF3aNaUcdK+9VLoHHCaW5fVtJApeQnh0HOpowGRQ
7fLc4f6ELaeRJnqt4R1n7DPRXXu3IAzJPLv3X71GlJiszuVEETj8vbj9gaQ1CM88SomrfxP9IK//
n89w/0bhlKDq8EN70nCEyAw4U3H1MnLewZ4ZcDZZxZ2O5UvGuPIoUnf6ODB7OLeDgIFtyYiebg5Y
6XkirYJz0/vtBnPgCPokxRzTS5OfOvR2bwrhvdUZh6e53ZJQiYUMqw3xd9kDI3Lsm0jgNJRfuUQT
a5axYip0tarClOZ2jJaY0qDFG9KiGOQuqT27a50Z3ly5A3wiSugypb+v4vrRN5JkoDfTCwZnfdnM
Va55p9AGaqoJZpflY+EwkLToxzvy3bsconTGAgXiLe2COsbNKCWX47TGBHmmhpF4p68GIF47a/eQ
6KVHXtfY83Srj/RfkiGYEsuxfnWCp5JTnCsT98ka2xnL/Nb4OWUi+DKfbGUIRlsNdum/3PvCbUfD
FcydP64DqZW37hQzJ1ZiUhdMMSR61C4UtP7IKIHBy47+Q1o3PhyA+Wkz6ksnAzCPjkkrSTPjVaMj
0aNWnJUie+VSzrYxVW2fznK5mAYMBW7zuZsGI19cpmzzQVVkzSfMbZLQ4F2cD7ovWW0p6vnN54iP
ZK/LGsid/BopeyNSo4D0UGUtWaRwnGd1ZRbOUR30XFgMRMygUG+0Q3ZjVZ2z87kycainV4/eDNa3
Q3cr+bYELVz24gu0SsCSokuqjFnycdp5PeFoESo+hyrdJLwdnF72U0vnSD8Be6BKzpJb04MwuSgZ
zvEIkw0VqKkf2wqUtwv0YLiDHeOJxTuMrYn+nd6iHytwr68/XBm4bX+iDsWy7eUNuztAhOdyt2pt
uls8HyLAOTwT2hqikp8/MUmw+3AFKfFijd09KpBcf6v3B0O0hLLbZ6WHc3AUCKWj4pTHskk6Ghl0
9rzDa3l7RdOi/i0gjwd3UluQmsUvI7akMORwVdhpOmlFC00zX7IamADfJLApwnhN5SyhBjxDLaZb
seTm6NOFKoyQBMJWmyOjR9IpFrwjQvBLodqix6P7nwOHL/HjqFcJKUekvZh1IcucI0qPxXr0e3RO
2t4G7JLT21K5sQLXBkCYyWAb9qR6B4Ps6rFE7njzbMqt/oIX36OKq7P7pmze7KaiKd+PoeXQ9Hfx
Eo7OxE3Frku592WtauYhVBniUtY+Qwsa+xuDHWSUY0H3JHYlxt30Jrpidps8Ht2qaEwSBe/W0sga
8wcXQMY6Ym2PeARFiqXeESaUIYve8On26KM3y/wcttGaSAMYNKDGSQ4wZ+cWjjFqsjQaBKooyzRU
Tlg++9NjZVhsYSpjbY2XxlFWDn6z9RTqQgF3xcTWJicD0zslodby7Uxxm3TgAYm8AEA7q9qAN/55
NTj17rpJTTObOfQ6EfKnA20CLWf36WCg1eIpbkgTd8QMH+vOyhCHNqi9BfOB+z8cbitWPc64k8TW
Y2L9fPam/hbczoJhLIUb3xxVpRNS2BpT9g75shQhYjJ4I0BQaDh7KjyD0TivjaeEm5Y23tAu7pfp
qcSESZ8PkoaDP/U0EJOXqH/2CZg5sSu6bxa2G3xSx36lTgHdAuK9QKf9GPbg4ub8LmY27CzGsnj7
ZW8AfciM3u10zBYEoUtYL4DMJkm5pmRh6F3BZV8Gms46KVove0q2URXG/yAKB2F1/Qve85brnoUu
lsxPxVb007Vi+oMsYyOD3P41D315VKpBOz0nvp0tYVkHKJ0jelpdtMcKdgXT0ytKb0QRalbU96+t
la9msCzJTpxQY5Z67F5KZYRfbNaqlfLyRQ23K0LiXHBdaarADs4Cmk+hrXzHE+oeq0XHOTGTOYbE
uJsIUkgHIDk83QsLGjfYQUpAVN6h5rvAYgsZo6kAZIB23HGFIa6wJFmbzxHuPY3XhOIM6pwbNErd
NB+Sx7gc2Jmv3hz1FjjZ6kFmzCYsS50zeXMPaaCFgsKOxC8tUESUO7luTnxndRvUwVH+T5phKOXW
9g0G0ijj0bgltK2HmWcDDM4AxGIsBU7b4cEAMqyp3lzDlRDRFgtH4/1lCP++DpfAx7+3XP8MlyVG
9v0xtqUDA44skOtXe1mlSdBRsHW6QmObMf/yvNIoAY0eRJ/C9hvzAfsKFGm8OJyM5CW5yM2u41wV
tATk2IevWpKSBqZ6gLGa3LhI3UXKXZxo70lJPk5pYHwLAI2Z5up9mBHvyXMFXXIpqBBqbnToZ7yj
A3sDpfTg8OG3kkympdzSofaQ4L8GdNAi3/NivEbZ4X2o7ZCkSOoPWmG9Lfq0mtRu2yBkbHYHV/dN
veuP9cTAuy9DU+kpZKz+ziYLsGUwlZk6GJTUV+sGxJWOY5iEMVikCHfGhOVrvAggmXrCKLa4ySSs
RdBc2aNt70dyFHFbcxik+KWGZKF/qtAgc5J+E/Bcn1LnB7zIwBIPi/XiB6xUIkzMQzLzxeJEct/3
mUzJE0x5/SPv7/oxmeGQzOdmL6IpBTpBiKrTeNJGkrIO3N60b+YJtXFFwbIfayz9acI2XHdvTc51
SETKkNf8Ij21+Bzhp3togBSj0iMgkfKHnFOJHlxOFi3uf19rYFRt8KzujcXs54v8kTI5Aub5TJw+
GUUjtxyrxE+yeKLG1/FuYwtjb7qPfjEKmLKxUMNIeikFBDxMMTfZxkUHf0davlsNg9EaJpgN3zH9
hXiN55GlF1NZ1veO9JSuscwELPJCkQ9BAdeGQA5tDa5k1RGPO7ribgPyuQsMyIuT6nRg0YhLe6JC
ciHr6kLMbU5MTCOqo+wQjStbmQb6B4AsWokBvAyIfVs2AVDba5amgqhCvnU2/1tg/c5XyWomnB4B
tvrwv0eSN5mZep6ROVLLlvbDnUosklWu+6vBmbEoL2LitMQ3HAyHTXqW05gM+COf0z/4xCbA/0w+
Z5Q4bITShbr6eTYdNIU1pmDXaEHuJaCHBhcaiiopHbLsue7ojQpp/+V19GwOAH0MitQjFvBKuekg
HhuTcHRdhmpeq0egSVT+aJLzuKi1c8esV06QcTium7Hdor3yZp99872fv2uJq9i0+dpIbImV9w1x
l+mhcJZWvgJKOERhlN4QMRlLxJp/bqNwscKz86Hhd9u2N3OmOzX7yTviR2HodwDNKppAXYaChtAQ
ziI+d4dOEj3CsLghEfa/+6otucFf4ITAhU2zayY7khy6k32BVg4tg/vZuKS2f8peo8EfCd9Oa8Zx
MUmHjFvg3RZpZQW4KXg5dGxeKk4+icJcooB9gWwOwUy4IgXUMpCgxfOsNuOquHxxhz7PsdV6WQy8
at2KT+PtJqslO4KwG0AkE8lYVIZekU/JMKbgee9BYeZnqRn7sCtJWnIc4sGJwlgbCwAq+CEiGwpK
9cEaR2fX8FQXaBVQ7Gk/eH4+ggd817o3UeeVPJ3StPid0dv9Qd8yvvnGdH9QV6/mK53GwVUzx0lD
Qwj5VzaYXpOQXU4Qt9f1jNu22kTscDN9Vv0V0fp4Xd9lMWt9Re+Hovmz3ShBF5Y7oKgIKG2ZvZxT
MBFinmg0Kl+k5wE9xig39pJaMtMUA587H5gt7/3/3CMJBVgG4DJaw93hucBl6gFFJeeBQrp6+hGM
aDnnUDcPJZI8+vi+hdmADGfw1J6zZbG9AT2SKCwEOi6UestXOkBd0ur794xpH87PJ2YSnPvJV5se
/cHZEaYbr090FVeU2qLMtJFU++jx9xTCD28zPv6v483H5m33Uhdr3+u9a7dGqdlwVdGyCls7qZYt
X6Dyvwho2qZyVdmyCfNroGYlroyWWni9QQDUdhyiFKnEzJ3GAjiEYZ2xRUVW1lA+UzUTy5xwJAbv
aIzW4jEZx66+5gAiem9CKiPQs+0iunZhTF46qSoi+a9caozcd7lb2LNDaTD+MCObU83OS1yD+wcg
f/MBKxtGHMJmpHPzou3/1Y0WHdygjHllbPWDTiqBVLPFehGOJCwx5PUrRpZvQOv/8Um4m8v9mtiE
8r06tXw7yuR+chOlRyiKAvS/P8iLorfZePtpmOTuXzqnt1GmyM5b2+Byo8Lr1g84geRTnkE3GKCF
ox71u4gfTd6MiksOnkqB26zlC1Ot+jV8TBkzJ8SWIjauq8FmXwo2FD4rZQiSr2T62Rut4vXp4IAw
dxkOJV93YLi95cfBCj0QZ/gJ1Y8K8Vtb+i7Zqh5BMDT27T96xT2F56vMUMYdYE1jOVz45xZhnRVf
o+s7FF5hHnuKqGnLIGJ6gHRJ9zXeqskvsGmkikNrOfML5wAf42voly2lKV/6LaGC0JMeAthI5gpM
Q57HTHzCeFT9tpKpjc8Jj4sK1N9g7cvztWeWWK2mlwq4LmblkC73AHylWmN3W07LXobzv8xTFISC
gbM6ZW57KxoDNVv1xHygO/nYLxZ6QXZ3XGE9qu2Cw+a/hYbp0JH+aEoEd980iDKPZSKtUDwbyjEY
6g1Fc/YmrhzfMZ344f9qFqAOK8UgDMwe/yNP2LflKEz3nhNlh33hrWf9OHeLIWQfUBPGcnsWHuKP
OySaAui6BjtCIYv7n0p479zT9GWhKgPPCU4jINDPv0Bei9z9po2wY2yxCWL+Bf4/r2qVRgjBJcLM
4k4E9Z8xZa3Zyv7MDtB8V5COdHMuTbN67lwA2xzd6UOnW1HUQ5gYyWObZ/4ITVP7W2ParfnhbW2p
ybiyMJ41OVrWLo9vxbR9Q8e7Fdl0SrFQBfxNGs7IXxEzNwmdvB6PO7z03C32rUxCeUdxtUTuuYKe
0cbaVaQL+ufsyN0lo3L7kuqfxIdGtLpbyNmUc6G0451PrIpw7rQ4v8hnlgFO4Ls2DjJEVPP95Cw1
FVWywFPNKH4ZkdVPBtim/hscafP3cy8XM/hOL+y/rHb6E3YvTyaPy/H7D+PtRBOIZWusHud/ezVZ
qsN8TnaBxD87qny3SSKLH0KoqkUILCGC7DXLIkO0VZTrSUJvVlnys3MdTS8u6esSIZme4lKbp2ve
j1lpU5jVEbDFOWG+w9c6WZyMhd2CyR7hR7nls6uMCUt230zDE3hNn0YLuNv1TiT5USJ1PSyZrVQs
AGLzkj7Yixj9LJWn5wV0kZKfF4HhC40RnUpJE7mEqzVujvUpIdGVHHtK3RPxsIC7ASRSgxsEJLFn
XbTXqqqLquvFOcRspuIndb2OLpGbxJ+Xjd24DPHup6Y0P+oGEe8KtXFj+lYAOnnpTnhZ3/zNEGzt
2axQOJPQm3o+LfBVCKQizFXTJg9TmENbp/0HNDVkLWO7tcwmWhDGjdaPnxZOhVgOP69me5g41hJ3
yoV1sLfMbBYcBGEzVZSnR1P/RVKCBHDeBhXPg2TBz54/eMse46Df0Ae7Gnm0u20PC7m6wVXh5egU
ZH87rHuMBcQxdkUyrHk2mZAzlO8wQP+/tO1SSYmAuWMOn3Wh1VicZVsYATtyswFsBkLVxq/3w6FD
FmPlemsN2Vgtt4a3ENmF4Mti2QNYWm5u2xEiCGZ+7tCsyA131LIWD083EvtxVYV8lNMBa8s67WwZ
GJgj0H2kvEKM0pCUTDJZHviQyRFjDi5/+9v5sVSa5UTy+jM/ePKF3bn4FdqnkHRippX2GLffWYHN
FM2M8AHUDVz/5Kj1xer/2B1wPqH3oxXb7YubpmoTsxbWwbj8gq3wPUh/QjQcr/Xute4TZ4AcjOeA
4+DFFixpWJyie6RODPKpvD0BjcuPKCCND69THSUqaryEA1UXWJyxGLhf0XLGl4jwFMClO/gHgICZ
ysCWTyk6A6RoeqriT8X2F2BcUahD9+p+tlM15hmCr5iIbpf2SosbiASF7jtBIAeHFLhkSRS0LDGB
YlJ9u8C3I/zC8uaFV0pJ7zVBFt4RGs8fpxr+MxYF8YG6+evDnt8yRAtHq10NTTqrBR+U73ZnuLW6
q5HvrluHdn9axp5BNLkRptbKM6p3CNhDe6l+peSPYaOilN4Rrt+Oau7fMoCJ0JTQv/hAFHvZ0wxL
o+ji21z37EgQ54scvijPosHLXcxGZhx6/XmZLLKnzfjqHB1ZFuNpO7NXMxjJCafiVg/NjVj/GJgJ
gxFhql5DIZ9kksym1DImlyDmeRrgnxnyf0OD36AJf0vgCDzcgl3vDHAm/R1pfKR0isT/ZBSQURl5
cvCaSe81AxadyrQIIEFbh0OdqwGdABzSkUdQrUL1EtsyqAIu/+9etIXDmBTc/oSeAbllP//xrvxp
9eKSFBz0VYlajpqzxUgCWIIMigzkMmfEcsZEwxF+EVAoOf3RpzJ+PvL+kgf3XhOWgqaCFAo/V8nZ
U7XGOzXNXKX96PB2oWNPrUfjm5zsVjgHxdgZEIWgaSAaCJC1lLcaGDfjWQarOL+kZPVEml+nWz6V
kZgminq9D+hAWeeJLDgu9Q0VXBiXOTqPYz6aDoAYGLitbq4eGzQvb7ilsQx2pl1e5Rj5W6aUlujt
8gDytqtqbvWhrk6MzGUKVvk4POlst0sLgvxFkZ3dit0Lk2NOTk1GQC9Ii6kTVJYSsBIR8USlsasW
/vvuvxuaYExyXztoJrnw6Yk2UeewN8sUuCPqaCzI5/YHE9vsXIqdBp+FeKV1OU8fvfkjz9Bxg/lG
Zq+EyZygTw3peiS7fy6X2JtBzstOU6xSegGM4Q+6cWOLwizyu2tDpWL3JpPmc/TpnCjzSxPU1rrr
Da8RQUi1qYAFzMRO5UQxn2stagfs7Fv7kewjlhYlsuJsNzviAzlWl7wFnxRyK+TRbXAo6vwoe8s9
8yCGchH+VKMRSOdTd3PN2G9XiWApTJH51dYQUS+ONpMAH1iGyV/2ndVgTD1AWOpoEDnjEWnJN5T2
5Jr6xjjPHlMR+vvTVUFvMG9By7aw1JocbViIHhljdSr5Uk8f/85GwKNwYPIT2MrdIkT+APjfymZq
u62qH00qHeZ6N1cRB/w/ATZV/vZ3ohgaxQjVrJeOLQLRGxO3lf6EPPD63/1sBEEWhJp4u2rdW94P
VYSJZe9sYTMIuHBCpwfOdQr6BvuL7vj7AGCuCImRoBHTvGwQ0mfmp8rulUyEsLtmvaN+ImR4IRRT
pRa/uT3UWfAW+yFVZPosO64BUPD0wiMN77pAgiMGM6lVac0vGzemxX2eoDERxgOJgwfYUru1wkXG
ZEwtq4WyTe2JsUOGtFV9CSgOY4haSj50bxPFsfu1gsU7WoIqfn4CCA2G7ZecQygtWjXx28PnHUnQ
S10yzu+0n18lt/QnHM/ZOsow4XikPHMo4imC+AVu7JdkLUAeF+W7ZcMJzo6L+/kW1yhDvVf/KEUd
rDddsfDTTWrNa74e6hbOfg8+w6kJ5FBMTIWZYMVSy6OjHndgFEcycoNM/ZHMQDDIpytQVYDGWQdJ
sAncokVyQKhp8EskgH7Ye0lV5jkdApyTAO62k6+9+m9EZ/6b/pKAWTolPsx1BMzkptsISKlOdCbT
4hrTeiQHEUHw9g4AFCMx5hqxb2gWIcEXQz3+Sq/aeKUttEmMiATXRxllxrR0aE2pF5uHled/hKOv
4UjHluCvCkRxo5WUEDZuOdhEbyaikXHgrWXTmXzJq5J+fg6l0ctFklsvaVy1Okx3SCyY7ZltEFFD
Y+1EolGFqu96kikKVzse6kE1qFPf47lQdEVS5cTl/0bb8YNBFbLosktUknREj/vOzv9H3H/bkUx1
sho9fUwC92hhXKSzHG7D1ZeL/o/K4v/nT46gH27FiNJuyVH6nVcbOWp2Aj19+bCNG0imkbh0abYO
TK09tn0+mwheR/2KBbM4xBc4DHw8g4pqeJMcRZzggxXcVRq2CCf6HtWpK8RD1qF/zE0kamva02a/
dqWg+qcDmA483rU8h0vU4QOrHYuCjmPMOVD/xeRy1TQocDl8jFgNUF92F1Ac8h5lB83Spoe6Fjud
mA9Nx7c9a/V5kDNmS2rvsDHiD/Vlo5dwWilnyYGvloJRYlMcwMSCX7Y2IhWcLyuNSFuYp+FPHkau
wN0kVxdMzTz1zpu9SCX9F9Y5ZdK6o8wyShMT1zwEgILClBe247swbQ4uBjgvH9q+K05dS9Ff2RlU
yvtgVkOKpxMhjAvQlGweQs7bV4JBvPOS1MRl4tGjUgaXZZ3+mN39dXKdLjb6jpaUKmayKpS5DFW7
Hw1mXvNnKzhKeSq2455VCunnZp502sNvY9hHlNuHFKfUk/uwOBC8L8GKaFvnV1+QNk6j5WnLcHSV
mVWcLyT+b+LhPcD4PVjlAzERzuvDaBphklfeQgbQrxHmtydrvXSiRcit8ZqLPvHcErtDiZO/xb9l
FHGoPZl43oM6bdnsQ5+p4n+bzhfYZ96gMAcYXLxbXhvMYBNpVe3bahpXi+Yw4Sa5pH9Y/dNJ4LpD
0Ln7r8nssJSbYY26RZSEPM4cQAYtK0WOxdt84OXYxULVWlkm1gx/+4Gl69Wt+aArWS85motcVbby
vbxwuU1GHgD7Pg31fl+xjhcsa0NfCF9Yf5sh7584btlAxn47IAEOOyL9dcO2609xbM1g9UOlH9v5
eT2C31DoC/B/jM8cPG4x8UHdfZxP1OF0pYeMVOuSvnjRuIM3nWk0kz9hP8bAMN7x+0wz73xgh58M
iZRN2Ix3eecO0UHqM20TreZ5zg0Yt6qUfwARlKUAdo2Vp60W6E29PLS28oTRr557w5/gFuDbt/eh
naKOunHt92glsDl1r8IGD0mlbkslU/bG97Ocy6chnvy2mUCg2WTWOlnnv6xJ+lHTOPXnDLqmEiJp
ln33dkRPDB5Db/FVkT4IkX8n2G2bxOwLsNl9kp8ysY/+8Gzg9L6X9Ip3tHC8YIAy1PM6ZrSb9nip
4tlOeKBqO4ruvUhVXelVwuEM2SnJ1HQleHWPZyBUe+XtPi6JFvrspMPrsIiIvdC6AkmHaxuAPxv4
Fp6c+ELXeo28CT+DJxpkI0mLI+jP9J34pDatFPglVVFU4uVhPZ0K7IhdVdd6rHRAnPnCicKb+h1h
1PLY5THs8L/IhMOfz9p/JhxotJBQMTaAIkKWqHsnxR4NwFhJGqI/WyiE0eKyyJ0aXbxQj0pQFzeU
cE/c/8oSoQ1uUV4eSbx0YcF+YrSQdd+7BgL9zaHe2OldkZEP9MpXsrWSKvZdtGGG1WBpjdU6VnSb
WxjTb9Nk9bqMjkmpd2bXmvwIaS6mo4RSBlFC+VB2vcuMELZF1elwS/cShwY5E0ara1aAmOhEPn2n
uTr6a2o4Tu6vyT/9DPIZQ2UoiMvS/yDYMfadCSqTgfIOuP61kek+9vBp9D9GxZwNpl+G4Z+YhcLc
cSxhhRj7sD5qSu1CDtSHa9d0Y3BKCsdJ5a+s1Ph7W3o4F4g6v7rvc6zItj8xa4AUCmopI34Xz77F
SEagyYNoLA3T2hDWl2ZGfbNXhdMpx7KYr7PJmuU18FctqrtHAhssnLHkScwUf4zUd2OssJ/pJso0
C50e4IIUizpFjXUQAhwquIyVOpf5il4U15de3IMbhitTBxM/uKyeuvjeoUtvS4m0nPOOhXf5AeDd
q2ICprXf44b6SxhTHjNeCpIOiR/pCxZobvK2z7NeAwCj7nX8TDwKWZZ9A09JqLExzL+FTUPX5sN6
9HT/IilRI69lKyY3wCM7IsYFCF9tUg0oEkbGOLQJAdC4DP042sb+88ds8D9NBbuZ76UmyyHqwDVV
vjDuaBVWXfMqimv9dBgE7Kqc3fexdsXU7Eh/PVexxvKfN4dkoIEvHXvoeXYXN7d68a2Rvj7wRgfM
OAcNHLbPKy2tsV0BOdJVR9OeGyyyDj1pFOVY/xbVid+buUTE2Vp+xLl0P6YeuVi8adUHPzE9WX6r
jHtMfwGobCHhh7MYuQQhp0LsicSv3k8/kHjFjlSxP3xbnLWGnQ2UlNd8GSNVcZuV/3iypaYlt+o8
KW3yL9VpyEudFSca9Gxr3zG1LD7dLpm+Q7DlAYBEklZ5jPx1rB/Qk8kOE45CP2NjCWffN6/OjKur
prSlveNYYAciTjRMQQgV/z80KIYVO/EWEGvk32RQesRFiKeAVnY06oM0LJjZSDkUeF7fVTEfKBG8
eP0lMPW9DaCdQLoy1UxE1WUUtEhMItmIWYrP3WCRh5uOumJVKWqXfPKKdqtqtg+ARqIcvp6rv84r
pDBEGKXIE10gHXqqIY0nu4KDR60Ny+NQ7H8Chnfe8dxlyi4JZQxh7EcETuq0B1LC73yube0Pokiq
+39k45cHQPry3k4jeXs2ewI6jd7mRfXcHK1hWnKVXmACZBBOFTCdyc0jSOl6fUYzgVBGl9QeEOEm
nlySAkqKcxvaQuVLpvYxMiY7vznd8Hz1+2Eo0Ylc2oticQsK326amXy5+6sM3fqLQ2kdK8a046e2
f4rOMk2j0o0zO1dy19vAQfntiD6HZwvV8hVMuHiulnYr4pDTGnzy+srZGq6VI/bdxFOg0SkSiHuJ
mRiAJ4IID3NWI105Y8pZb1PM2p328Ej1hcZ1+cQ+8AQpCDRoBuq0MyOZerey1r8EAE75BBVzcc5S
l3lnijCezg3fvt3aHE+fDtyjwu3byzCJ3CtUif6H4CK9VRp/V1gG6K8F+7RWYo48l+NPLxuKj4k4
lqWt1x0jREGtziB4oPs4hSreMe+J5HMKug7L25GqSmvb7euHEU7zJabOlkqjhdCygn80KulYCC4Q
7/lK6P7FN0IPkjCsWuYjlj7PrHTjc8MNqXD7F1GxP1t6v1BANE+GbSLu2wis3b/hGXjGTxZodyTO
/vf+zDCJnmGvJyntDa9ivcbgWgS9hNICrGODDb42GHqNWkL2Q+uusrg3mYz/FwdgVKFvNCPqVIlT
seHWUOhFy8+432eCfFCfNECQoxH3UcPJyUrUuO2f8VukwYCKf0u99v78x/rtyfRVFdWqodTc9oyU
d5ooSuNLuE0WajXyzIFpBjlXuFNTSRCOEMO1PG4+SU72M6Ul4Ur7Cv1f8S8g9AHrPJdepfCs79ev
iGhkVKYQeZlEDjelpcDSMVwAp8c+1tHeZNK5Uv00QTmntBhxzoxTiADBFepY18dt4LWGwzYFnjoQ
g9pJ5V9sXrT4UaiYaNpdllwza3mAwXNBMuWls2rbE3RmTPp1qw+L0f/qeqwqDNY9XzaOUAWkNati
LNsI/LR5KGXEXFIJF2NyfFvlerABaGLyNe4EHjrT4RKCOsH0fGrIZebtvBMgjHV7mlMla4IKVs5I
ontAsiVRUUMyyevyf5yWhYlNOve3nEydpRZ+FevQH6GoHLebPKP2RJTsZj5TjJ3cHcP8Ym1MQZIV
adoqkB7AnLDBlS2KIQnPDZ0HbWrtDG8udRC0geD2NUvapjPjo1gaUg8awzIXbDKokMb6epxtOzpp
d6GA0QYf4Ho+xdLwVVoQjO7oDhYJngQJq5rkLatP4SMZTuP551QBPUAL8eu8ZmRmMniJqXT8cCne
AjAobX1lctbD+ykvsSdQzWUFDa/YAfOKVcCv9laXIdl8yCeilOYbOEF5QSKf7E6q3/q1OkrDPmYe
wfF4t6xIin2BsUza51mDE8WCXLS24RYG+SDWhmmzbRncWZh+XXO80BXv+3sN0dEV6OLggry/IAGG
pQHc9izQKbs6IxczQD85xSa9BBJl3FlvtlMqaIZMTFHdBO43HHc1XJYPyUnsL94nUskck8H5IEFs
s5jHUK93uXiUWGONtqKx9tqpFzAfk9L6LPGzCT+mRF8of+xGnI0wYYoxRnWo5Y2LelFiLf72SmiN
F2/Zy48+H1WeE6z63PCrraIBHDBKYz0+BDx/gbgNOhjjeI+Slb5DPwaQ9bqJ2ihrPOa0GAcjhBey
hg7YlqMayi8SQUda+YFQQfz0nXRcMLP0wD2zKJj8TPKaZgtiVtBj415iKUtSnz+vPasbJ6oYGkGa
Ll5unKBhmTeRV0z9zdrrokyK6hMi746mPJWTIEgNsQDr89HglwTDd25l6lNjlJvxrhq46H9Uh/gb
LB1pXVwxuTBN2OXfxg0SeIRTqysT/fOuZpjQ2rbZIgXa2jXuGxcnvrkdBr/JESwxxQrAEfK3m/Ox
igJDXaHgJGNRzRnTd0GjvKGCE+6n7DVuRjWx4RTsCr50VkXi0lbMamOYHNNabbeuEtluXfV5ONKm
1Sq6VwQpi5Y6FOvR0aOXidjBILSfO8T5eXwdc1bkczM/JFjHyLHZm6lgChenaumROw0DqbfPVPs0
tayNJLlk0qFcfSjUNT7Z+8nAoZnRn3/ALIpRGmXO9uy4JUZLF+8rFS/vsDHU6FrQwCWeQdpgZueD
4B70LeLgWSkj/BhRCXx1S7tQmRUGzE4nvB1mI3VWf0DHP5t8V6lTmm/rqv8gTFmaEVru2YbSMCYV
LMo0xVgZHQdhncwTiYul67hzF76hLEoddDVuam9V/Pl5cGrrMwhU0qQEM7zFUo4rc4fZ8SIfr7Jc
gLOyje/Zd+PK02DzUDFlKpd+5Hns8LIv2pMRG4BW5Rk2anHorIWgtGFlyq1g65l5e2hdLkMTZfVG
d5ppmv6sVTIPeACodbDptxX0Q1xkUBEZA6R7bHZi3nvy1CuzYYrx0WXAJvlVlewqIrzTtsjmNbpK
hSMyeJMAalBJQQJLJgDl6lqmrb243sacpGg7Ijdk/MgEXM8u/ffGARqQNjYbQxY+nKcEhxQn01C0
VASDLN9b2SslLCex6w9euaHT/CWpx7EjlY1NibTYxIhxPEK0Kzy5Rzq2rWG4Gr9re87RmrBje4p7
rPJALTxM2RtBfY1Gyws39cApkD4gfSSSeOnFw+OBCfGCr4i1r6G5J72dZ3/P0/p+e5MvIKcdHK/D
2Htv1XYom6pcGaRJ8i9PoMbW/2PBXeSCWkcWFC9NlwCDDMrqBJlgmQCau4RIblHhtELZpamG1D52
LZ8UxjLGWSe9D8sELH1iqiY+27QftelrE6AtNqcLt6wbyBUFEFadPkoZCMTyniccrpymCnmWHDdO
kv0UyNilueBx1xhEVRdTbqH/U02ZrDCMPLgZ4l54NtC/w8XKV/WHA5erHMSJ29Fyg8kNA+yayi2T
iqOgpvsM1egm3IT+IF1azrIGQVN16VrfNLBnEukivPdd662ZCpICu1pntMtEbGBWzNKBnnPsyutv
2VuA3g1+CktaQVfAGtd3KJwIY7cU+6LekIrQVuMHe4mSI8klCs+RekKbrby3Mjo2RWmfQODXFBBb
TBJIPJvlx7UYgw9xhHfZiCGZ+12loLF1Av0qmdkg8hxiRG+bjW+BXvmncwBgja3FoQGsg0vT/lq/
XDivGMnf0hOI1dZzIbPlhreYVZEJ72WT7zH/CgOd9Ly4Wdh4SULOR0bXyzKBb/A3GcjoF51XLsXD
dbH47NTFbBteD9EIJotT4W4KjcbbBBT5TJEFUrLFZHhB0tm7aDHbdiNEzDVoP/XJjPN3dUZlb2nx
/clMicdzYuPo3olkf9Dc204Mr64EBh8i+veqSWs8IraM6zNJcuEUPeJeR3+Q2FRDg67uC3G2sy2V
RjKVU/wKW9CcKAhMjA+sUMMRWAZBzXPAiHf74raGJORgSDzGLi3GN363n/VMJlFGfAWgWIFrnqM2
WhSoARc5GU2kekyBa4UdJ0AXoBChkGkvNnk4L5URyJr+ExxBp7CRSBC1nswACuxIQgJO5I6ZPNSL
yPXrl5WkobLN244QfiWguWdTz02gE68Gx+ePTkX9DJ3pAGgv7K9ukYxebWhwRinKcEYnjVp00Sak
DrP3XqcIUwXAEElyEIt/WgtF3jQaDvOkkIUysIOSmgDJLocx7ZbFu2fuWh/wSoEq5Hd6K+OqjfVt
kwuBdogKGJQwmWzxx6qAtQT5s+SOW2ge7ybXOnJjbNihH6C3kb3aTmvMUU/K0gR/0e9BNWqs2wXC
DVlcQMnaO1UPUAw1k7z5fQdEUzFOZ3KA1wJA6icntF3x5CfpVEdYQt4YX2bQOTQquKcfKhFWgQKx
UPP6PEvGv7dTu7Ib+9BkWlCqKUrF388ZuF9jMLkjYATEokzob1GnzAf+InK7BoO+b4FsSw/SvQiu
/CG/d3Y08RAFWnc5u2iwzZcQjnRYYo1/oBPeOoprTtAbtakMabiXyhuLRC+GblFoghrQr3fOUcl8
uVPAeG2QL/pgoz0TIWL1Pdm9IeM7Q6Sdkj6OYy+8ct1QQQn0+nNB4otKJCwlCsbinmbt2BH46XOy
c2oYQ6pUQ5vUB2HZfVLW2v7HCZWDwhlYk9u9cjbBAeVqMVia88+AXqJ1EH0SoRJpBU2tW2IYPvSX
sJp9krteQogVqTzrXd8MOYkqxb1CbOtSTzUAS8NUVRWZDB/PCTk06PR1GndP6wEtrqoUxOTYqVlQ
ytEHmB1+i8vU2zLy0cOsS6OTQGq+9Oc/AxNxHjsQDRkMG6iPODU+qmEPw9H5NuCNY8dkpJix4ggv
F/yEoF1r5vgTnZR3qkwm4j6BdZiodOdfNGqzry9pr2SpgtYeGER0C43YTWJrYRNtMFVjQJtF93fF
oT9a7yXfvf8P4QpAG9srhUfPKaeMT1HHk0JRryDYC3OVjunLW7h608E9SVR9UYqRT2S2EQvM8N6A
96Nqf+K5MloYOLoBUaxt8SJDo9S6VKrkFlMDURNTjQZx61gUHhPsWUVKbDtCGHHO+dZ6JKhU4bgv
ytfOKfmNxlF+vVNn8/6kmoEiOoV1wNrrEy6VIi4fhxkHVBiwwGJhWsNrOqrjQE9kh+imU3re4Rfd
ZVGA9l+icLWh7LDfbw29EeYSjCP7xe+lsoXT0PAEHCMakyKvp/D/7Z4u5o8rna4VdWog1HQmFo2N
QtmHFxebWPEsEAXn/GxZSwR9YQJq5ZbIOWa5AxkeeAqiBciO0pPPXhNUC7KwDbd14GHepQNtQiWx
+a48hw6SPy5FeY3j539cazj13OKX6HydZttd3iFyX23EnAubKBX3QHDQh4KQXjwfQJbGiVv4fBW0
7PY03jp8ek19EZbTUflxzenNHciMQuIrQ0sDBjY6TsHtgMM34xPGMHVCGPlKMsWdzI6yODFmwl7y
9UimAY6Krp1KYA4nJfexvvNTltzbmUJE/lpXSOsoKotg/x7CtLngH6MSs/tTkcwGInrrTq8yKcvs
Y6xxtGpTzVL29cjlrZgIge3CNjSJ2whCN9zjEiL7hmnWMSgp1n90LmHmsBgm+YTPcF6hEgqlBNW8
JQUJLhtkiIv3m2csrd4sSWgtDxzpGhBbLQBAWSJ0PlA19JtiC+yEOJ9fiKGRf/S+JxMCAuhhXj3+
Ng2lLmV9N4Ncn7qTTG4Qo86TYKaI4qR/GXL9I1mabRW+otMuNxh7gLHtxFO8VlNrtvh+v5zgA4Qa
mEJXzyl93CW0RHyonYKNX3RDxWK+rPHUABKAY8Od5YJ9Yoj8cTRlejh/NXFpepl1QbuNNT//Jl05
w5qBL855Oq7UDUZ0u7xpdQ8ezmEoG4UV7qSGRa05D2GF6L0K+iV0VUXQaqq5lBosc2Ky/gNekr2u
tXwARMQWrvGWHin0RKJvEUXAnS49ousxNrDGclDMBwJbsy/2id1YquwhzD8UowoIEf6Gm5SB3KOV
3Kivvaw6XqBARxxeHa6u+3P3zgRqMajNFFhaHSTaXvFRhBD5zObLMjowki8c526aLlQgM0Ixyafo
h5u+LQUohhkCre8iHsPyOgX05VK97Vb0bDn0ni3oT4cVKNjLUbfVf0A4nWGjgimfxRdLRO8d2QBl
9lmQAmNAUIc0yfdCh6h2HJixlY2kGKn167zKopyTx9UIryMt8jtZIWmf+r94ZSeuqqv/z5enUQ+5
FYBfAUsc3r2WQeSjrmBpx1p/KTNB2FGqhDW0AM7Nv7Cd04HFfQDXjBBo49spxUZrcZZ4oxZQuy4B
ZYfU17UETpw8CeAP8EBu9MYQQvCVdoLvXoxAq1zpIU0bRuz9cbrZdNcr3a51CgnKgqiHVh41acRP
ynSqH1MiwvaybA/eT5BrBW4hsejfQ6nMk9W8qYl9kDgP5mNqZhiX6zMUnkmjWgyCvpF6rEkcKM6G
AvLQeibINknooKa9inDRsXCNRK20t5CaRG+6Ase1CGf6r7hJ1QTrFW2lHGxfstIOTSecWccYyoPn
3musdvCFFZeR/cKPRz9tsYPh1L/kJ0blKpbvl04rS0M4jq9UWlPP6/juk9l2o82e8AhoGywxpKjw
ZiUaIV6HTlzGqMiEgizw72pS+t0KQwtiAByhrvP4yyCUAkgUJplufU3A5lH6Znzt7fgMfBqJaeh/
HaRUl0XwphYw0wQDvkeJI1F/SXy1+6zvlVJf7SrUid2YNtegLBJDDQV6DvWNxA6kTSdmmxv3/9ct
PzEWJp76hucDs6VMFqUTapUZRDNtESqkH7ASNTe7CCNI7rgHCHpl74tgBBF59Gw5kGL4GtPNgjDl
3fVG+2j1E4thuTUI8arpatw+nplEaq3cJdvIvRKXW8vOeesCXZZc2nYf1JSKtOlNcuQFHXyK/vye
USMUa1djgxJTOaLtEuAKp/kK5g+TA7wATKDEVHcXxkpCmcr06NUw0ZutZ6TNoxbzAOn2903yxAlK
pLO348HeX9PuCpn04KIm2+GSMHeZTiA8qFfBvtE/Ns4967yqhWJje2cVon3iDBRa9DpDP8eeaIun
HYvB8DypUNpRh4hmb51aU3o39zHEoAz378bujZXakVjL9YPK8QsaLJ41Gv9DDnsLQ5M2ZDThaQNZ
gp5f96KY95864fFLbcYhyITcbTD2tHRfub3xu8fBiVXW1g0x4h1F+JyuWTI0tkTCU31LVX5gxpT1
M6ExdmVAzA9ri9FtbrXPgn6r/sJrNrNdjWkzJlioOcFtK92E6QfSJguuJJbY/JVDoVZf1rfzJe0x
tPXRYi6xSRek74ffpvDma1Gqm9F/zj/BUVic5W+bugf5XXbD/q68620dlYeUPFmlvHIZqs2obewG
6Y7opifHEPc+S+gidjUQIxE8xgDCFUH8IhBMWxm8e/jCm+sq78qGyUw1uzCloGhOPz/BC+AHUFEP
szd3mRoroue0fYXDQQxCIUOGonYWeaa93m4Sj2L30tSMHsJoOZ0WJ5J4V3WebNSCmqglftlnnBb2
JImGWKIVoSA4PXamQUKJ2VE4400DpyUM/dBVX31EBjjsbNSX1o7Jr220yhrJmGAsv31g/qRXF4Xh
bZw6LdDZ2a6uRIRszXC0AKyHSIyLLqr24kk0M9RjII7Y5i1zsh/dPBftuTVTgWSNQy7xVXsFK1Xy
ZtKevv9wq/zPS66KxKYaFGrhehPFC0rPv02ci/LmJP9ak1FKReJOScV1dA1oXwI4H5MD2coA3SXU
QHMSFOCD0U7TnvIrPcUaWIuowlYv//EK8cbk9gZ5N2lhw8nyBUIPujfH5ZElnK0O3i2+PhDBJIwN
biHI/LW7xWTz8kcmP1ggRrEihyz3xEw31lQCFuFgJzMlraoEj9rmiHeFmuHix8lggHynfnb2Egrc
Re6ZxuRXj08R1pxQju0XzdKpkuV+kNnVq5X64DB0pwncruz0rcnCkkX0k8yCg+C0+6/xdVsUGyWK
JUyrVIj+nO0gU52+kXJ3m5ZBtsCLZvwi9RLHdjRMqGbMy7tf+Dqj9JOlHJgWsQi79Eo5Yl/dX14F
NCiRKbMjXwexE0fgYVb/SjqRtZfnUxysudzo5kvksZm6kS2tvbAsVHKuKD+nYknQziVeNV0OwpME
fjaD8pX3bpTG2apnA9V7f8+s1IGYZg8HDJgyCFxmp0cjr6EgxwFaqvM+fJBEcO827nbcfVitoSfZ
mr7YpaNZ4bMd332xWueq0YuJwWeTnPBCCu7th7vIGiyLuVKp8i+DI8cm47yIPzL51BYQUmPfiETB
HI7YfBRZXqwcq9HMy3INexXOyRpD6rr9TpqzSuBdkd0zj/83niBLwWwAIKm2e1C1Ok5rZd+W8CMt
Zks/Kr4itrjD2RZD5LfT7hYd6smMYGSIk6K5vOtTi1//L/07QY3eE82r+9SpQBad5ommVp95crAj
qON5af4FY59YP6nwe+b9xpmEBGF1kSLEBdAr0J1CySWWE6hZfuToxBGNmUppq1o7Cp+gEhFzqt9x
vOFl9TgQs/FDem/sZOeC7um+rRlXTCW5S6woJIkOCWXPUQkGwfqZocqCP2y0Cg99xHebUHUIiOpK
fqUUrVKGnsL8hYnw36Nmyt4T8R5I6zu7InoE8D9OZAUeDFZQFa3osIUwPf69rRGkt6DDhMG49jrI
9qMJLp6S501UcPRsatgbwCZF7d/p+fsL1Wx4CgvshFVun1EhM1c9tbyri81lGuxTXZgHYmu5ElD2
c6po+XqBYbLYTNl7MZywozJkhrWMnBGzzpHB147csWt3gKYvUXMQ9WGHIWDCZnWNpqxyNbWOVRNp
17xS5Rqde/fAY/3Schj0tjdYs7HXKRk7ry3eKv9cNPgmRP4CVjYRXE30uiRd5PuMR9OQX1hnaRYj
xtxIex7nZfatoNKp0nLNeroHOCwx6h/FXkapTDIL1IuQWhmzZGXb6ZfQWEkzBXsH2Q/7c8aWVgFk
iWSXsnXy6H7lm2iOFUeq3fvyZGcfZZbdRotaYM7BAoyMSwtZThOxFvNpNioofRp20ok4FWoaZTdh
dT312XfaulxZ+O4Qy6hVAKwb75agmO7aLgbpql5WLrBClrlKL7geBMQeLMKjDE/iQVXPmEXu5Rhv
0dBbNrkptXwHO7g3NYiIpotoin8fWgIsxj/eyyABtN6++w8LZfMo2zCJJMgHBCr5MhnEIxzFYiPj
yc0pQciIKmp4h90ybOzB0c7c8vagLpoVLho2/uEH/Yl5jDY6q8IXifE4RMiU73ESTflZPIDqL/W8
ZMCsB/o/lYQaYILN8aJ1kxJC99DUPvcJjaXQTtVV+DnhethuNSEGjDYW3q97ZWi3r6F0+OV07cyN
oNbUR9uVuZpMAL9vKSAQWOO6VmjwuaLXnf3b9J6JGdC+tudtRlCw9aCrcTOkOOumQ5iB6zrKfN/3
KuTF2KRLS7lVwZ/LXQ4al5C0KLtkaCyFyYSoM9Ti6XJBNF7RCCqeBCpNvI2kY2GV77RlYPqASo48
n7Gc+S9tnwGkl02iz4Mesuu0TmKRUpOqwJXupeTGSCvO6pzEIdMf9pyigMsSqyniBeouoJFkJXZK
5jcis7YPuxXISnxbsOT114wHaKtENUPDCP55p/Zl/jchv0ZJLnOk/B9sXk+kZA10Vqj6oxaztMHn
snCaijmdm+Oa/axhZC9OU6/55Qoea4jJ3Db7/sHXbrFZ8EcAiSDxnBEgDJ1Q22Z3sFUQpw+jt3uM
72tIwh1g9CTmVJ96kKqvghuFOFY0sV5D6GURzaOscIU+RFKEWdweB4RAr0tEbpx6mMlrx1QarcJL
1wL9t5Kho68yZi9Wx4Eg/deqVPVDQBtODzjrUUb+qDXc76tEn6ynsEbYAqGf1nIV4hvUkStHYJ8l
WR0hyqxp/nfz0o6fXxY2Q633uc2QX9Sgp3lTJbNnHKCJGl0qDs92sldcxJLMiEuND0JAxQfbt+RO
5mkcTt+XrzzSzPiKF1TnOaradnu1rYa5rrhufQF3R62wTtEYfs3NMWvo528ObAVb/0xZSRw8ymi3
MK5NOfQRntTLtF6LEyjwQGzfdgQSW9X+Kq/EJCQfB9o5Q2fLQY0FFDi7ipT/qkYpJoAFemnnUkdg
Kx02QRrK3i34nWiCSgRWrSUfWgSEnvgSsupdaegjq9aDEqp9+kZWoUtgrQVCTLpmgQtinnXuCj+O
tcsjHIxNvmJ/eX5dcNsxzDdK/R2xcWSmOKkbaa62PvDjOg3FVQWrObyHvhaZzhAvDJPT8Fwjg/Xh
SSmBZz/KqodvufyGBxRuMXgd+61m3bM6j6wONynTgdEg4oftJYm6dyazN+s+vJ2KRi/XyxINGazm
MK96S8FvOZ6YYJn0mGF94JlhU6lqxAiyKbkLD7+lcKfncVhrN6uDMDRspvn/Sl9RiL8DZL7JUen/
9dX8K/52I+wYXWvSCyJzWWra3AvZfEG1OUsZgltjpphdXmiAKfxW9LYSc2WjPG4p3VxvPjumU8Xt
JgTTs7UuyFguisTwmy3O/XYQcp86Po/vlhLULyq64Bj1s3MlwKkE6Hc9x+eqApbc9f0cdRC/bAG1
0KenQmOTUpMi2xJncm6f3c6t5PhyD9F64oNEv5YZ85YZyg8PK50HxskVGWlK4TDzzeav6BdxXRPY
j7Uq1hwhPynFDzcBPzMs3scVu4rYo2Is2QqwmltDWNXfgH7m82UEsRPzBk4DTKbZxewjBQAEigz1
gRMHKM6qOtQzBhJyrcXWKvosoZ9zSMJ8WojZzWihUqYTUvtkZul4o03PU+oBkXjXTxZ7mN+QTLP2
NpgDtfrFL2X/KDgd29edAOV13jGC7FlgBHWkFE2Rl230+YDg3YfBVgMp6ammKNCRWV/cduHnrD5y
p3J2MO8uu8a52UQHV2yNeoVbsEBDfXbZz1MsXcmlG6eWlOFZi3QH3Naxf3N6ikGsSsBoQV1v7f8h
D9pqb98zHnegiUIYwIULVn0w4diy7qyKELd5n1Ye8nVFhTLsQnKASXPLoStfdVcvYcNs6h7kcKU8
y15aAeF/2jGKwueUPse8FjraREhbgXZzGHdKkHXRT5RykTm/DIP+n0HDJPMC+FdGuKMNIbpVlZ1C
4cAYb5H9/8GSwdSh8fQpRCLUvmj8+KF8dUsjpiO5yMOz4YYt4GhFCBJ1n7FuNGoOHtjU7duVhiSl
J5LwQzoJb7P2Jx9SQGanKAfP071O35sK6C4EDdVSYqFTo+uuIRT33oksc7Hf8Vpm5PQGFejNGdHb
KxGty87BCHQ/GG24lg5MNNY7/Ed9ho5yglKwkGSJ8yilAtEqz9ewezcTCDDo+HhSYBzR/RRHB3xF
5DN13KcSX+OuTqwkVKLdXNBj5YdqNzIaA635g5+8Nn1YZXA+Yv6MfIN31WAPc0vFdtyH52Ryc2uv
fSxST278mb5aVGweZ0vqL4kbOeaeG/Qnr5QeSGaljVxmhAnFOtkqu4+/AQLXkQhe6yUmk1x9Vffc
qCsxL8tjEKO3CoKMrEmV3A9BQ2YzoVyRFWylbBac4ZBcAUrmQPh0PtCkMSNRsffDpFoSwqiwogvW
CITTxTjzrktfFW7bxM8RtFEI+KHw7aWwUTbgxDGgEigTDXENczoWb9IU3mzxRZ7GVCRJaLGGhkzt
HrP/RPgZn+2k6Lz/zCvmg6Borv+X98k2t+frJKGyCbpDwQI0Nwt1cnrbAjm5Z1lqhC06OZmqixEs
2M8jDjo/Yc2CCmvA3Ub6zaZJrYfkNBsba83bhoiWabXuSfvM3WtboG5cJlQOdE5mdEY2OMlwdR6h
K3IQ/Sytxt8pG4Im3IaPqPqDN9k4s+eUYC7rDIy5WtOaNnY2FO7jWuNc13MHmA21oViTUBTdtpb0
C1kF8CcR5epyGzWMgrUtk3Nt7zlOJu5cYXnUTMW0hbiaY94enWc1fYMfqUSXD5eD7U+gkDLgAVNu
bz7SLDnqQw2Ei9IzxH2gTK9pfWNbJ60AZUJo2oZCSLMKXbiwMGZUDeCW11IxQJCV39andJxOkCjp
1oj0HI5JQ3f/zT5hWw+oWkkBv0ZpRRfXaE3i8MSpZnD666gbsxRyqHSBgKV60QKH+KjL327I9cTs
EOGLOYxsp1J9RjXe/u3iii8k5y4GqoWfoHmkk6AZh97qdrBNDpPaGwzh/Y1e8PUy2NWK3S2Yj2JB
QnkWSjTtF5/XewQ4vO81eDMux/obAOnVBBDcIfyM/GuY7itjfDGfcJGoLkIcHZcWrwNWcu8S7uGr
rnTnIPCEcU74EVxz3mCAev8kvwfvSTvIUw+TCpExKoD1MgIgF7e+YrIT5ujfXHVzhvrZU5090bsQ
aL7uqfbSrrjZz0J/IH5XX4jofKnVb3chB8h3rj31q6q+QbU1Ffpfh/jOVqNk0tndwcN6RjVMm1O2
os7Ps2P9k+0T+sDHJUgQ9uA6qz4clF/c6S16YRgioRceDRkh5HzLTJhinr/Cm1f04EwugWxh9sUT
gZWlN1ScZH8CwZhsSX8AEVJ8kYZPBmaXuGOkEr7Jjc7EExxZWYS9D39x5g8+bYsAwKmUnUC+hg0Q
U6kONryBHLGPckvajv2q3C5PyYA2e7MQP7ifATix8qe1T1PIz+Lk0eBjTuXElPsKaURfwdrRPBvD
hq5gVS0BCcrL2Sx2gZE4Rrb1oZKrG8z1aqfuxjmCQ2A4fqo0c4NSg0stpFtS6cUJylsE5kggUcsV
pa2vSgQ2mGiXeLSKeZpfSvVKnfYXz3Y0/EyDwgrHFI6pnrw2RqKddlvzmA1+p81LLbtMFLHcRESB
obmp1SfbTGMbgMAym6M8pY9tGQXA22bKYrl6zpEjebkMcrqybdMJCXpv+EFuR6q149ROFBOCEQj+
fYTNdRfdKDRgWs4IKmDM25+KOvNk/Br/5gtLzI7RcT8VXf2L/4No5pF3bDzEzOPUhzUWCH0u5JHa
oL1MqjEWmMKFDFJiV90eiQKCok+2tsI3hiQZTPrhJYZlWZowJgCMkqVj/YH8bOYIKf++deDONnVL
pEyCNHZzTtZbCaRYmYd6lqqgVYiq0XtoWyettJMQnGgWTJPz2DDhciz9m76bVUTKXzhNo1H3koPS
Ymf7/nbQvVUIwL1+HiJon9BcZ2W2arVwfiY49c0Zhaa766xC8v4G9Uwq+2VaG65iTFnho/mhQSOb
ACVYv/dh/smMsFUILmhPbwSJheJZAHMWtEYklq89UIrFa0mNRRu4NfcalZb+O+SaNUQn7tj55mbC
iksGmbqFbMvTVo2VE7J8FY3uJGw1DMu2NMfxeC+1NXi26lPK0wWKO8QHn+nQs2pI+/vA8D+owzzW
OT0opnUUA6rVlk4rbZQRZTahFpW2QghZkvh2V8FXKHS2IS364SBunw98mjUkz8o9sCyn2Zo0CncT
2MU0zOzaU3Enz6gYubAfoR93AIXwIIndx92HiKmwO6IJ4oHsMh/Ihfah8LAp83MTbbkM2FCjjQx9
AGgZGnl9z5nGknINUc3I7wKMsaWi2o8qWsBDp3vpEDTy1WTkmxOGn4NwR4cdsYKhB5Ak25cAG5Bv
xdrQgUOh6cqHtewl7eB2mtqpuwTJdBAYGiROgemkUE516E3aesT2z9wHZAakaxfZOpS2x2yBz25s
vUA7XnEwMduuAKMAFGnMm5GglywKY+aLsr4lwNDhwka+O7PcaGs4Es8I97Uxf1hzMp5NSuitwViX
XYRW3ctmnMRCucVXWCcTFY/zJ9+dUaofGVYxGgfKf1xB6VNLbTZaOtMmHaHQkC1bLLZHdEjkZ4+x
epTUtoEFuNPM7k66OZmsu9FNfdgb4GV4c7HRouFBDCKMS4lQEKtdtsSHxQfPzgbeuc22Ol2poNFa
WP6GMwpgimvOqZZDTCR9D36yWJ+SEla5pwWPBFsx5F+UROcKLowavyeX1T1UyoDNQAtzLMOLk24F
+BG10nklEuYsjERPBdq9KvWYYdUJjl6Jud3JxnXJHcEN0SoD0wvMk3v//L2qXJ2ICnV6BrSdiHsB
cJWoXpmMMl319MxOC3j95m4xd+HmJGj57LxSkdWPzOIdZBn1O2rSXtJAGjNTu5twlfrFlJ2AbueY
yYAxzpmj6VbMBP3E5DO5e88qQHJeo9T6NfHnDt2vqGH4SbUzgZqvRhgbViK/D/IYIDuibc9VYT0m
eHgfzkJVs3bMqG+OxDSLFPtbOH6W2TGAcIw1yd0gvAeLYv4jckTV4Pl3Jl5BVTtfTSE2PyCYibO0
CmEaLX1NGa21fnly6yjuA+st3Lj6kcwpDu5TOej2aDguQsBsQjj3EYfckrW0eiBCeVAfkSvK3Opm
8GD2u3O/VOLjVEaI9urzhUDTLfYwHGup0FcWdA8S98yr+iD4LapLTeIlTHXigPJWRkNWp+xqy19F
sk3zmfCiis20zMDSlKkvpTI7cjsee0+nNCw3agD746NrXADMGJzZuf4iMVFabx6YAKGAb5iCMnRk
qs3pxmFRYN3dakSvlChaQPBv5xAWxhh+1CMnAfP3gbnOa8OMayH9CKpfVJprMU+s5MfnrnJa9Hrq
ke4TCX+bALYOSXOIMBSRSBPimqIurqD4Xmj9bj21beY0nCeUWGlVibNCIgmgdH+3FuDWfxSnmMY/
gNISugBUOtEJeotXbfbxHxnReJQBQAL2Ov/ojaUUjw/Kgnzxw1XiNnxxbg3qc8m5AXcdxmOXNGM/
NpnUHPeSIYcbd3FmoHw/pM0b8U9ROZze2yceuM+8cC86z1Ozzq8gQ+rG1rjV6YnspRYN6wCNI+iM
4Vv/VqblkukyD4P1M8H57XjyEwHfzZ9B24SB9HRyCl92Z+HKd7BaQut/NZ25+xxIp/OYQJWrLbeP
3FLXHDhsiXA/aQL0OtTZSdu8U5cDza7y8Mu+HrKcEnv14KZRAtbUQpn082wOz9yIh0eP9SY3LFgo
aSK8m7alCqNattNqUc1NyHuT6VaAW5WEOnAo7XhmKnH/ktt42jk0nY7e8uNevN/qOaYUBlCkL5i4
x7j42xDtAlQ9tITHL4nUGUXuVRmDNOwZhFWZ286KbctCanleVyFHptpGTPB4tA3DfuvmS/sHiQKJ
E/rBqAiQAagbkX1NXCV7YDfoMlOy25wnOFvhIdqwts8on4vwFR0E0vKs3pUExTO+En97/ZRazYFY
CXVA0KvRu7LBtsNKhNiSXr2mnFBSnpDQpHl2iHsp1qgKBc312p3qgHkmAsMJvRuPUjWCh29J8w7F
eQ7K4j+WczSqKshvJCKjI87gRsLsRzY4QTUTo6TjlZXieWK7mS3FkvpH/9RouhZZSMfChM7l3kd8
2JhLXObBSX+IIYPoSundKpdEs65u9eQu1dR/oJsH0tKeZuUIYIUL+sJZAYFg6CGrUuQTXw0yZDO+
Bh5ngALer503oVPAAaXjiUnmBN2pQiNHfnS2K9CuHZuGkwUQY+9g/shGCO9x78AOSqpGyS8IQmS4
xYT/DDwHqK7+m3ib2P50mk7dUbXrkMejn+qcIogOr/70KLwpcpAk3yQ8xqYggDjFIkLzXBWw/Ov6
q6QR//0DnL9JBRYW5TuDr7fLiNY3Rm9fMHt5BGXVR5PX8bABpGDNmWuMsusbgnShpFmGvsrUXmnz
9VwXhkrPsstGhmIDiUEtnKr9r4WXJcrwqEJkkWFLKxN6V89tUhQXP0SGKBGAAr98vJS1rMAmKoht
3YxbPSGs0mbO8dq6myBtHrxtDSKq+9HWa5h8jvMOYSMdfrM3ZTOnlda1viq8MXeEbhWgiFmVOPlL
1TdJnHkKzvZJDRYqKY/hezubbpQRaHBMWksR1wz0dEjkiodHMlDXs3K5YgQGSrJiFiN5b77ZTods
M9hYyQ6PQZHKIvZJXS2fG7Q07FcpHjAnFOONcDIb8okTRUCQGHyZ2dbrLJZONiVwWiY6be4ZWUol
YBHbLPlWuEiulg2NXnh/icsv0zxTeg3zvQIA0+N2KLvHZ8aVhpEBxjQ4IkCpM5SGukG37mTqa/Uw
VUHN6FkZfsMhYynptX9nupUpysKUFkAPqLevoQO5LK43YxQO11ElqUJLBWnnUtIrv/smr0x5Y1Ey
J3tM5edtTXVArei5U2aYDIpoGE5Sh1Nlp7fsqIxBY9god2X4jjDHvhWBWdNmJCgQfJj1OfJnwoB3
OODGw+kvVEJKj+MU8mj2qN3Su3nhMgumWomiYqLXcIJCBfNExHFnwOklZ9fVzpR1qW/kvBhp+Dzw
1Q9ZwACRpbWyvewF04Avgl1AARbAGX8MU7g4VJfFa+w11l6MlTMG8YXTw7VRIPfin84m6b+5Or5l
KNSa3GUFE2h72D73TPjcXFg6c6OH+AU6+LeBbI8lAs6iLTrD8qvj5em6zrObBX3HMtNelALNdMSY
h0+xbzYnCoUCujjJxKjZ2rX56owNn0cXzlWuOO3cHZQ7VE6r7u8OfUKcVXtsy0a0lZAzA09Juwzv
H6POWjBUk5LpvxK+G4X/4DsRXcO7abxlhG1nHOlPWlaBM8KhpLNraL9abekpRQRblPJ/8X/iJEYX
2LWI1NfJkC12YAawpyC61AHYClaz1CgEVYLof6R8yhCNCLEK4qrDd8sAtxr4naCKwOOJ8nGTHjDg
BJwbJWEyrqpFq+HdWlm+jcR0UUqevkaZlupGDHhuFVz1qfbsdU94/1g90nnUJsG0ztl2eV82KMRT
aLg9Mt8WNi64FOAfyLYYmPeMsw1/YLLHamC6+AzIPj3WoKFwadsc9xwPiI9mOXRlMUfpWdxesbqp
ngoJgYojBBK5qBD0sF0wsX1AFczyvgYxz7py8BHN7bZd//fQ+323E1uRHzjDUK1Q/IYh0+JTxkmC
piT1gp+jKJpUVJ4Dun4iDt8IpCoqvJF3zmQx7GK2Ju5q8Tvu9kEWCzoMf82MjryvaIwGstTmJUay
tk91FXzgB4ZG0TdcNtFJHyjNjxH9xeyYc7mEnighOxeLCVslkgq3bZcGM9GIF9Co9Ar5QAN+2ZJ5
EQP4/c1WW4+IYHI2uG+E5tiWqWKh2xrMS0Qt6O7+VQ/U8MLxYC7J5jNr8RkqSg5lbB7ht2nVH3K8
EMQEa2mNfx/oKl2P+/DMreskJO+Ze0z9512ts37g6mBfQ3mBV1Fm9pDvOs/dITUh4vh4KPTSHaIj
PswxIp4J8ApRViCc7oHWg0/PrDeUA+kqy185FvcMZA5sHscNFDlsng0qzKGWzuP2D6uKZLcGsiRh
RX1b8Uqcd3o/5sdscUKTO+qvyql+95thqn8TkJjCSC9ohC4cDcf9vqxRduUqZOgiQmKVVVlNUCKB
OiAOBGOl2UPUNKwvCNO2ff3Gm5r6NKMi2nx7SnYcy/I78h7bZ2Qm82OrTIZudDA1vGffU81fi0r0
pfZbk8oQslHV3dqmbHRkog4wnObdeNFxYXIFqHH0UfT1SwDA1NHozv+a1tzIyB6SlId0j9y/bWHf
LwF9xAIjp+MfCKoXW9UtnbJg1jjhjZ14K5sQL3It2XCi80bxjBIp2ZXUyngsgajpoqKQ2Igb/IAm
36b3+gKvrY50rxNU/5ho+Hedj+uSWX6pO+wJcls15KkONFGc9DmmZ1efftyPW9tmlhLi8dsiSdgb
N4+SgdOYhyXMPCcW23ahGrcLDXGxTFAUJIyAzPulKiBNRUu753UYFHDk8oBNmopA6WTaAvd4bIaO
cJ5ZBRcWTKcDovPrHQ00AfIa8R6wDvi+pUNpWiFJ3YE01pqtDSG190hmCURBu2Z0LF5zDRNJO232
jutjP0ncXRFmWDpeMSQjQeK6eZd71Ksbcm1gTN/VmRgmxSO+pkbYGpMJfq2YcYyHbIA1k8Iw0psE
rvSxWgEYSheMOLEVd1WNQC96waGjSomEyp+i2C+i3pyO0ZmMes6jWVPW298U80PoAvoaiV0fV6QP
BTn+Uwb+fhiadHMAAnW7pTmWYE6EE2FwkYTOAsNSPulrWkIYWXs9xyAGOvoyCUoEwfKav3nx+agM
6NkHCLoWG1I/vHNhDtyAKwiqagF4hxr+y5x0fhktGlSgz+tMv6Mx9T+WaCDUyNvjuofZUHOpgTCG
KRM7ii2V7Y3cc4A/DhEdDa+3Vg1gQJMvajBGjf4iZ6wtgjyJZj6Bh/usNaqdqyramWS9UccXWZ1v
C1lX5ajHJ3NwtwvQZZb9qtVnOMWVB/EGR8n0j8hZ5fYwCeHjuiRiHaz7msSkb+bEp1/rQhtCXtGv
AVHSzUIFos5B3yppbw27IHu7h4ZVJa6xPljNQlU+2hPIC0EdBgKEztm2U87efWAC36/b0KQ1t7rg
bT26utUeUiP0Mt6UfMH5ZtfNf9JCNLB5dRzQhQkwMxwEroqJHqepxTDRw+iQOpjUWw8ex+eSZp3K
W2cHzYR0MSpZfT/mqXB0vvuIU8ktHZh7NXJhJ40HbZvgIaafWAwtFHNwC4CuHKe8QFzKFx3x2wHP
HwGdfF+WLc+Ts14m09vUyJq7B7+AAvvOamKPouPZ/INZXAHMF0RN9cDpCT12/aHniaAzqrOV7X3z
Q5CWzvGTIKJyOizc1dEK4wfPWiuIObxrDk130wcUPdBARnEyd702c9pFjKXtNxrGhpkmBMvJY/Aa
kAGdJ9Wrh8iI5BN7YJY8KaxRtnDieyoGNBi8YBSoYD9Zy87PE5O/ast8zi0yXaJmjURNJh9VTQK2
ietb8YJNhsTNOSlJO9M/eU0xP5V2s3y0BUJiTgSjKDy9dzIzdHWX7Q405NPvxX0/X9xSR1+L7dYx
o6P6KMLXzT9BS5s6S6IFoh697WZQ6pcSY3w57/UilwBhWu/gqEnqMeTBmO88WattX30ltVq7gH34
A0lEzTneS05je7lkZnljS+0hsJ+YhE2jRsL3Jbuin10bCtyLH9vqx+vnquaaM3Mm/WDPUT6D/bM6
wNOIc2JNTDsh0GkjTipo3HpDuyWYXBn9izR3YnicXSpl6TpepNOsEA71LLRf1N0fZlaVHN10GTVe
cN+mn45UBhEEXJ/lpTYaWHvnpW2rtyQFAmll1HBMXZYZ/p9R5EvmDXecIb5rCO8Qhwk2BA5zSkYJ
wd1dLOIAwULOdLTOV3AgcGa5D8E4uK3brpYYYdrG0wwKkn5HS4+Uru/mfMY1O/6zMX3nge506O7S
bDKL4QnTUOIn8kB3d+WujVo/rt5TkrMoQmpuGGkPdrHm/eVboWGTP4nAy1HE9nlU6YaAIMIvJWng
cF08Ttok/amY4ZYoQ/QN5sxvBCY2EFZRyNNT9thuDpmcfhZU3Il4LWFCXir8Fb4R+1s3qhFCTFwJ
twzpHWb2KktLJMcoc485ogUMDDukkQCc/pzAL2QohBoYbPjjF+Dbsku3cQYW3FJczBiH4rmOF+Q5
d0kBm+3WgF1SpKe0W81rfq0ueHOyzqOVBF8Kf+X49Zf5VUjT5q7h06cvAfT3uO2u43O7wV93Dhar
mCgi7aR6ydhgIG1C2Xr+qiNwtVIQAG/0bsadURDFHZ/M4FB39CVdXFvcji3RO/rjEoR7RY/BHt29
ZcwRlJcUpJO93ZXPXKBqBSYxAiTDxQWgH3JGpQFEHt+QCkJCeczb8NfOLE4MsZ+d0fPp21gsH+Cc
RYWzmWfGprusS7JQ7YdBVR/6FCeC5zFNZ14UFZ7p/8tZ9pHnziwkXw2t7V3twhE3KxCUNz+CpgTZ
PlzX9bXOMVDJSVpQ/GQtm4dKttRRoR6VOy7tE0TphCcSUY99YjFhbMyp+PaL4vNNhVOtAxVlEpIq
PYQL2HbEVHn/jFWOoKR3dd0eOixPYgBCbQhNT4g6BD7wXnyAm/7hut17zioX38Zn6w8roUWeNuaT
sZ5vk5x8kKWZdDmPFSCw2hWARRsQKmxisROZn1NnnpbaP41atPOGwxH7D/BF60nvtinDuvpMtuOM
DF8CsmTz4COfAHy1Yg/Epl6npEhjapYbHLKmNnwCYN3aAMKTijbiWFIreniymmDMTJUyIMBbUG8c
AzlrPUiJ3TTI7YlflOdP+r+tIO5YyxF5J3IR16BbtRDAAaid0ZOZdvjDf0i82osaYCK3uA3VtZ8I
osSBOkbiZCPkkwv5qGFq8NknKxdku7uCeCBCAgdhP7DFe9vmcLckdG2jaExveEpbpsoWzXZGgs/z
y9LkSXyCRw/JzWha5Tzbmza6K7LdwQggVbbtNFBpaXbHnJaVHQtAGssI6wj445pB/Rjfiw1DJcV5
aVoxImqox8nhAq81C4N2tBpL9oOMT1B4+WWSwKYMldcshyrMUAIoJ66oZ5ZBH1/TWBqtJSWQl/gX
UJxi0bD3XDwcafmieym/rGqiNFnqmlOfWHJfPPi6dweSK81F0LqlEPPiBQhGj3QmtYat0yRRnlLA
eTmHQ2mtFfW+OmUvJjTLJ5ztxKjKx1FuheMlNOLFZryNm8gjdgEfvJ01tHYotlFB8kv9QKCKFs1V
TwG2xnVoCdBH5D6GWEK4QrQMJxJ0x00/YGemnvFL5Ujc4xyHCLfDdQMPgdbV1RW4CsVLF+wwRC2Z
21L8uTv7FSr78v2mYoXHJOwo8lWhR941Dyxtojmm/LeyZzfA1DpWqszcUTnogMYYtEz2l+26b9WR
DFCWblM+0pJeF3CBrsvz7CN/ARvsNaOHcqy3nBkkrdppcXyOd7J/Lewj+go1U+6sswi5stSoPYAM
dRJitj++yHhNWHzEnWrwIGLdR/Yp9T+tB4CjmQDfSvr7nGwiCf0Ro637Y+yyz/FRi2TjXRQHQDzd
COsQJtO5xWp0+z9/csQNXKtuAXtIjr3xqSekOKQ7MUqHp2oyPnxjXDV24v//qVGvjZNv86+PJS0g
HvZ5uFHKqUYLw6FJBc9nykksxqoAmA0oD1L36N4NUJLcpgK/R0sBdTgC2+yNRIJvJiDLhch8NC8H
TTE2MW41XuiN4bgfI/o76T9EkCJX5bkQkXtWLKNKPq7mZqpGrDOHS6K05rOjKC4GPOR4WzkCSSVI
phh8Qk6WhJaszrgqdpfPrm5RcvksUGjygtFFAfyTAqjI4A3XKOZP0xUQlTt1GK8u8SYx0oQeT/ES
4h7GsguXSo1hhWaLulzSBwkEaxjtEwjXJa9WfHsmJBzP38MvSXC3aFXEkAXJNC22qrCz+9gVxpVJ
F/W1qTWP45D0/XBQ48RTNKVVQMTwQHNW7G2YZ8KusK6tRc+B2YeWXA5Tkp29Qty+UZ0jpa1xV7LA
liVriiff0Y7r9zyNEsuim1puAZ0GbIbtabhdit/476Bx5nRpBzvfQDJBg+QA3uX1wmbzEtOr2yid
Pk3e4OwHKA71fdn5tLZ2uyli7vgLdfShflNMGn8r1CUj/cTDzDi3M0mrj09Vj49nPAZrYmHnAf/4
TcFBuYJtaAXXdYb1BB/axnxAcPfiYsJhdj7kgjBVpALiGSgk24IsPRjjGpOmQs0CwtRZMba1Iq3S
/mUnGWFb9bcjNWwMr+wS9+f8Ykv+LZhKF9ZFws5+YPz4OqIf0DNXkLtQs3LdQ9PP3W/M/PEkYybX
xiQaXA0/46eDsqyGHiIF9oCYchiAkuZXUs2UvWjmSgwOZMuMkN7J5PyE27zzI2Mvzgfg+kTbvr3z
uobsFH49ZWOPyQa2aN/JmNcoSXl1EurpNCH814BT734nE+g2G5/TClDxYYiS/dCb2thyZbDgTnQp
5cEjEK37Y5NtHPP0qQ8gLOIQkjxOaUM4ko+NBRxvzIIlRsW/TSvr1aOBF65PSaibZKoO71xsd2CM
LBmIgPnVuSZaDj2QLFj5IZyoRsiBw6Tht2UUjfzk/WWDROgEjZJP3odaaM3Bnuebsfxisea0+Wxl
qbxF/2d908xoeW8z+S8lQhWxPNyvBx7yhPe740qPBbvpVPJz/FD1AsMtDWDVQFnCoIrUddLGn6Gs
SCWq4VSoi//LCKVqkptRDCMW2sEdd3uM1F8rbvXUiahCZLp3I1J9rrgtD8u4XXXWOXZ1hlWS7ebU
WXOMdew8X8jGsRpu55S06GxaQ8xEbmciyE5icRWAoWMUF+R9CJ+OlGytDQ1jvtbWVobenw12unUF
eosxNSvqD66eybCOKSG/qFghObZXPg0kqA9vteT64CRTzHDnCxATLud+87YGVD9G3Exdx82Gi5ku
JVLua2gD7xzJsZB9SBtyfLrNrb2INS5R1Zj5/rxLB6mK2RqFBK8RzFZ2KXEJTscO1z1ITN742VrX
5p8NpCe3syHU/AjDcJoMWzJzkoJqjN+CaWJxr47c++6GMnOmYLfGgYbFA0cm1HCAXfkcnur9bts6
ERWEaftaDh4CiIr5FEnn3PCmwbnL97tYQBO1r7Y2ROzU0wMQcnvIrogeJQKpukmMwmqxocIdYyk+
oBnfqtkhMKTeRnt5jUg1yx1phUIKrB7LJzqWL4XiUwdPFeoqcm7EK0IbcrvPeMPGzKjJG5uOMtxb
OHMgPvSelyUNL5E/3lCHv0fZYWX+uT+l4SA4mRj8qHJbzLptaPscVQLpiblUbfpK3dkL8FiiFbas
XsfdJYFgielnalC4lPK1gRDh9/d9R0LsSqhP4JYe4vxyD+OFQVREekBMYWEjEAMRIknmK1bhLQhn
vmnag9cQ0YdSzlVjIVueEITa1CpM0ESpI1PsCRivDUaNuWsoRNjYYxzgX3Lz23yFXyJ42LI9M5O1
g9CaS/vgB91wuel1+GbG5EMNGI5lZS9ZoNL8cU2ku7pBluqAvk61l80+mLRJ31D8HtAO5uPupcL2
rzDTOrmteUCa8X1tF6sqP9P66YS6WwO4OoX7ZUufE23uW2Xi98qmuNjswnoCYv0VWLgBU+mvz1fy
S8uBsCAj/NuhKr2OWBxNmNDOHxELQabGV1MBeyDodGlBPZONxRA+LYNaaZptRMKrBURHYJ++u7NL
wxr3H02t6D/rOgCB9gK+xkh9lANoA9H8OzoVUAkvcY7Qrenn5g/jzV07NrxljBq0XeCh3ckH1bDF
c6pZxdoQHREHswR65cT/o7DqdDtW1VyHQFND5wYs/gfDWOBkovw0wclXAJ7d3r8qmzjEZzg+c7PR
P4mBQfeI4lH0hU9eKtH0A54w6WWsA46ZSTJ4y2qBdtz1rJ1G/fdsC0ScvTitXjw7Q8PAkGtSqcvv
4BNUeVBQer6C/rrfT2bkny3MuwZdD2YFBNS+Pp5jKCvbqvxPEwKalo6GUY681roujhYrbViZFxbk
9WaDHUT2oBD16A3lpWm0HRQYAJ8rJZ6FSF8C9qeQyKVCOdYR/cvMyqwhvcgMXtbhC0pNVb98jHxX
kVSGR/8Pe4g90do8A1CnRUBOXuFnbXnfJATZd6cAHEd/NDCgnvCvFrvu5qK8awDn+PRPIy2QWV/H
etCgXnWWGxAG0tsmV/jMQeZI/J2G3uAMB0aThy2Ctyxlzvrgfuw8S0fkNDV+tyqelZXpaJQCovJy
iVNEgcaSG0tJOnow3uoJkHGhjeQSlEzDjwu7Q9xh+LVcvu1n/Xye/rEJ0VXqS25LFnCRtcf5xFRN
8TJ6dLSE+gSUtvl0MwmZPJDAltDgBogDQm4Ks1lGFJ5FCa6tzoVNLfHqL6ozRQoNCg5l2wsYJukX
2LtGQ0Uspg5S6420IkfUZfZcduaknDJXsy1k/5tQAXznKttcmAx9r3dwUYfRGbHyA+eKcmQ2sbLE
IYwyK9OdJ5uwc4o6OlrGEUtY8NoYRoyBhQs5H3LAVVW3WU29njcfLby8jvvmIGgaKRpUrqTU3wdJ
beZkLGluaa+GT6RpOhxVXPLv9MCqtfMZCsZu5iZl8KfoBgEfSnlcOD/OALykS87xgvuYTas8F94A
7FFL3t1MIXVkA/L3VYhQNfNSkwtzlp8UhKo0YfD1WomxwDNuYRaY6+A/Wy5e9zO/mXZD8rfeRzwe
5sVtZ+NV9iNYWUcwGbdNdIGIb6nbCvkpUFU6TJAaknoVsvqy/EKDI2D3Lntt8Dvge/U9vEhXP5j7
sECvyZ+jq9Vw+04qvE/WI94UcDQzSq7GmEYj9h6yP4GE29fB6QujFYcOSIRfPeIPtaufz7cTWRgu
ztHwdknvxZiA7RV47OBHcA1SRPrBj6RzOxlmj8xdXBeZQkkaEGHIytbe+y8BmfCXvLSUUeLr0fOQ
bFJphTJdvBPvtoFh19bDvoXTQhLzO4cMIM8Y9XTrdovYCGLRSXJ/O53W8J4/sMWou7zn3KMIy+u/
Ac7BF2u4W9CTSVBHApoYhFxrmpBXhHhxfNwN2OzsJbVuNjnOS/C4/trkZ68xloHBMETDguiQ4ecR
YU6FVGphdvYIoBTGKVYeUCDhMUwnnoGfBj4izq/kX5yG2fWlGi2NZ6yALlYuIYS7AL0rT5h6qDs4
d7efoqVQgQQwKhiojD9OxzbjgnJcGOWq5escIzf2Zjv5xSH+Ogq30s5dmRzhasLbzrW/FMAyk4Eu
k9e4b0lUUuGZ8MsIwyixlIXvuZ7+8vJrKAvA4zFDea2CVPQwEP737Sm/1pCSTczSGa0eJ6HScCm5
SHWLmX684Odk3SB8oIza46nZsARSOWerleOwSAyh9IvojPKLRUDtZbOVe7Vs8zO98r5wb8CQWoNE
iZWSl9BEJTGlEMIkEfIrOlSTPcb2Xwk2ycoS/BqCARUiHvJc+qV/wwFyDyqQXxuC155LXH4G6dwS
CZ613/IsA8hOztuFI42x05vZa9vmhVkvtH3dRhNJpEzU5J9KahHeFt8q7kvObquLuLCG3VP7iYox
10cE1x9XcJpjDnRAqDm1AR2QcnpQsSuEr+xe3JmhGwjNVNdOGgcH0TbIarDNlRUBa9P0nE2aP8Hq
t79/f8oRwSE9uAvT0Lnvh4nhXzioRgoMXp/McAF+7vPcH3qiKvAskutjIFsyQIZ4ygtzL5TglEgr
KA2kUYjpCvq++kaCHbhHhPHbM/5om+IiKT9YytElIBkNA/z5UuS+1eD91P3oYCr1kMoO9+PdssFi
xhTtUwNI+0Q4y07MxpXrCh77p33uVW4QMvBj3lWHbpgqyBwPEH8O8QCgEJNUMYC/abaN2x95qbRB
brRx1Tmp57D+uRxh8EIeWcyxagWRQ5Al5LUw//4OQfRIThdHFR9hD4I66PsJ81KG7Y2LOWxdws1X
qW9HjhPewex6xp+lrW32tS+sc+jr9ir9mZATp/H7wXUdXDghk5IbV0TegAWMRrocxPQtnXO0Qvir
d+Mv7qVJVG7mnPlLU7t34KHzZt/nlw770oxzEdBRtTQxbIn9MQrQxwFonF5NfLxwJqj2VA0KhOx7
3E5/YwPRHt498WBVgoek2Y30rCmdRVHWc+zrEYi1o5ktI5lDkVajd4Zp328gwRk1mM19sZUjkj+t
TRdAELlybhGNGKl50LU6WeGSBMGEgZenPjSPVpX4a+JPClFeF8I9wlo9e2dpy8wkY0nGatwfHARw
fG1FVq3ZObg1fxFNx8ZOe4Orehz2IUIPy4pRiSHB/EJtnGIfcHPU/Lj2pHIIlCgSycYGAJyrQm47
3iKSikS8SQQvTAM/YcSUzZZLvfQV+pN10pYroUYYDeBpSbOPWwc09HgQ+Ue/wcvOqA0fSE0YEGFw
WBINxRNOsOvxH3+kCxZC27rg8bvQk4YL3b+ON1UOx7+Cpq6PYinpzV2zvlD5af7M4S5B83K63Wrv
U+AZbnbuPnroz3n9uxf/U92lEQSZHVJulXolgTRQMdaw3gJFE84SBx3/2mlUIURqP7iD8jxUuMxy
hcQvhkrLymnBUl+fp8RvRiEZK74StnETDzq2o+bW/XpvxkZLkOMCawfoS1TFeNvU7ia42Q6pCtFj
UQ4zfD5teXqtqf5IoQYypGDiZEcx2+/QXQ8/WsyS2xB1Io6S5X8Vqg0n0mlzzoqIHQkT7jK1aUrP
ZJc+2IPKm+R9aEj1aaxz+XZfYKaWdHnEFyJqoP5VXsn8LYxH4f3+OpmqstznplNB3Bm7HWo6tybM
MZYvBOn5sQSF24DcZCYRIdvJ64o0xdHXLLcmMET4/NOYmzSH9oQ9YEL4iMd1abET+GnmY49nrZB+
leDI/Oshh4n8QSXYHfzbnkIwGNazYU21e/e0Oc+IHKG5ITLsNQ/4UiJrXWG094dIrgUy1zHj07vS
QpjtEGe0IuWJWoKPKJwmQqt5baWq7Kmq4xXrV5Rx8xJfYuH9yp8M+0sRg8G1cyP2Ur+ofTPQGZ3b
3oR+OFpwXXPEFrONQKM9Dvr/4dk8hw10FFTAXcl98rfisxfTt7tcIQujLYlALS96KQsSnuDWQ1lr
exNUpyhtPu/8mmMekyEnVTM7eIpx/jeoPecAbbzuuXvoAVC0MWIDe0ww+D2JwQO6aW6pMDFT0PaB
JGxI01Wq/hQcEJ7hWLY6O8PfKoXPCMy+SwqR3srTZyUXaQkvV2fveTUtWvN9poGaunGBGI7QfbA3
OloHH+szhTpcs+WrW3xajxKRZ1I86hzv9NA/kSGh03wRWVgVnvzuXB7N8k6vC+qQJEKYnMpfM7HU
D+oPL+OB7zN4loD+AXB8iXxeU00d8iMX6amG4N8ykYUVo/HswoYcJ2TDzm4V6AIXnC9vZ2ZkoW2J
nS4YzuBYB/9ocLTap5erQ91qeYB8wHHvYmBy0ru24eNH1ekviiTZjw7mSmbV2OGoz9kkziLkKzJM
Yi+DmJDnMsYAIe2VIs++VF28Rt0AR/ynWH4HtMfxSh/kY8CS53dUENDRSS5SQQ7kMOmQClaz+SDk
mo2XI7qHwpkEFYxvgCJ6WVtkRX57MhmF19GhYq6/Pi3i3SQTTCi2HG2jMu3qfKfvuQEDhCeGMkI6
bRO8uOBU3azcarSvo7FNfwfjhU4cc/5MyMb5Tb4QjCKQr19LYIhIU7mMGvxQsFeM8SnXSF1XlRtb
1S2aJchr4UntLBUGYuwMjp3NmD0KLs1eQuErwur3G3hAcCuNT/4hl31ttfkP3xYIT0xC+IesoSGC
ZkQMNYqayaF1LbN79i4goeWVCrW951B1C5GTeEgCIjh1XeSeHtYi7+bukhRqWkrz92KD2bRNb1f+
0lnunDALdl7M5hPR+Mvs434YywLZY8TE/h/d+mQFFVKCQHFv7aN5/m1idAgM8SUkfjmAO9WMcDc5
Oy8jcqt9r9YVXtpFmmvuEJIEZYii//t1H0aJks8c1xANS0vZ1BmE9ycFj/R6i/tF2UZP7EVVnT8m
5HdQGgJ976OXzdxkWyotaCCidcM8pI/rx/0JWktQ8bS+hhUpWbWPfZ+iys8FFMUKMvoXU/gu9+FW
gNeL4JCINVn70s05rADkpj+DWY03N3mpmjY/20SDjeEzwNTRi5uH1SGOllHyKKKhMLsCQD1YkiFc
zA7DKi4lrQIdd2LBi5d4AGQZnInWYJfbs4q33kdGuqZzoyRWO+CcFfHK+ZGpfdqUXEFthC9wZQBI
CizcAU+niJzRj6YzKdOJguYRjpwz2p+tiutIweLJT6bPikg/4w56kkj4mxG6KXzb5B2JhZzAL2HG
3/5JGuaTkqP7YyYaIkS/2VcSjhQcOZj+5uo4h9y3JyfC9YjIIHELVSJvneya+79WMbbZsGlDLHWy
RP6fmSF57WKtZTE0h+rqHTecJ+szYflcJRyBOghCl9kPTeWSSi/Prkx0dw3LQwORInjZLYvCbyKV
srqXr2lkWzwQuW6dNQWXLx0bYQ3HxURq6DwvfXOsAo7UFWFnyDgfQea4ztU2nn8Chp+miWdaWnsT
5f30mdkAKQ0/X4+baX8QxI3JsgY1fZkjX/Gpa0JR529qvwqP7TfvaUqzhiqgFX8f9KKn0ufr+pPM
ALnd/hI7Ytm/mXnTlDI0ksV24vBbO17pRk4E4XRbC1yNEQqtYF1dx4K4SZ1AoykQowINCMQUhQFS
Mo4pcp/T8Bf3uLXlCeBt9d2P4Ot3G4AgUTpexTgsb7R+q3fFEe0i8SUYryZ3TToIGSMlsJWsWPmV
sTK/f6z6q9MwjAEcKZznjbjPWX++tamrk3DK7KmpZXT4RYxihDs280VhV+biDJkHeq5G3pqRpIee
eKoGLAN8zNhl+KqohjaZrYB+FzSGxlCs6h6o3cBVj1jVVKg+0qUx2xuQJ2IgAcxCXMpaAP4ozdLo
/JCrXqo+SxdeiRo9kdipFgQ3pp19J+l/FfygYzp2M44egwhOxd5EcHXImqZP8UaRu+f9zBkSii0K
5svcp2JwL3cqiGEq+CJBshunlAifJkHVpicayyHHm4NfBvkDbK2FxBnuy24rl2k64tHHqSUcB27O
dIXOdo8sEXN5U/wTxr9+DLj6J91ZtDRdhEuxymEikPXkTHxt2gLqYuPW2fcNDQjzi7AHOa89QjpO
9vbbd6tnNHV7nL/qlfRsfiJYdvkUge58yTjE77dZylV2XfrDctQZkMy8AfuubppkZEB76Mm1pnRl
MZ90JjN7XMruUSr9ktVHkdkDQtNXXo2kSeQ7DhUCMtug6i8lLkfv3OWMSSi+iF8fLzQzRWPQ+lCN
mSEDuF3J9wEVSGBLZTcHTCEHkvQF2Cf/WgHj4kI8Gu34RpNcXkCE4JVEuCrEflBXMumpHLmaAsrm
t4NPxUv+QBSMVyCIfLKqwUPgGOxBdzXaPrMbEMzX/S4+Cx6STr33VIszoEmrC6HnScMe/Eqkn0aY
IavE6f67TkKnp6M5GC+6n4pUE7hNyjLP9e4g7niEytZZboI0Xt9nLiKLeIIr8a1ZnrB/a1pOrgwd
5Qjtt6OhubfKqqJEeRn/h6veEYbKbKHfnsUGNBMMOKbwgW2zuGua4TRmAgaGbIZPm8qzrYcORl+0
SPXezTuQSXQFtNTxtq5S7Vt00Sz7Zx8a4KN8nYbmyTAwpp1qvskORu5SAzZ2m+fjtZdRC9EA/ntH
aolClKuCT+oTFGI1y+Wr4PfKZbRjOgJ/Q5Jsenjt8trnxZcXAbjqKLMNpY/sib+jVhJZ1v1Mb9TE
psCvOdSTf3644FxGNtMCqfgw6HHm2cDyyMSrXMUFkodDymlD2GnFJU01eUgEWc4+rlNgKP7U7y8T
Njrpvotai7IMY5uCR3pnYECwn9TlrrZ5O9v61KSLU0SoIkOlUtBVHzPg9o5Waq6Zr+BUAmj2s3CJ
wvJgY0wBzRhm++CdqSvpzypVONODTneV1Ga0DWf35yihYn2vUOOj16jPZSAKURI4CMZdyzDp+nfI
mr4Vwamc/PfCZBz2OWfkATCDlYdGNA99T8z03grw+7i72YMIuZA6mTi18Yk46B3yuqcISzTEYvU3
HHSoNL8vGs5+W9DquPwrL9TlEArBklptN7mEihi/b7K4ZESpjD1xFW0KAMMI6GKqsqlkVkLQdET0
VPVi1vq77qRY8qOwWhH3LiligDDgCNTT+nBR3BBJVerz96/N8XKSPl++jGlr5qjMAC1T1R41iYEC
U0tuGLNPShyj/dTVr5TqaZ+wlOusQhtlAK3HmEZqSXKSTQez9IrDH0ToVzHO3bCtj8SvUa/XmrNM
xM/DmaclGkjr+WR5j/v4OVI/nOUwNi3NDnBSA7oWxUA1dUwsKagPdx247utPNkFEZ3xUKAsFQauQ
QAOGkOk5qQs7veRGyg49/vibCw8/9y1nXvP77NfZubi3W0G4QW+UisJbPQqNqeHAl5vgvx9qmfw6
Wy5wdcIskTUf93m6yhOZ5rBkDfTKKJAnBmWKOTqYHa47zWMtNLmEDY0MxtUuabROyJpEB1G9BL1t
xw0PRIYbArihFh+DSAJlvtl0RZZXml6ks0WmLjwTZS1K11L6/5JqfLZDYtxsbbHtYck/rhaojU0F
m5xbH1noAHQRu7IBT12a6L3Zv7KbzdmD6JgCAUViwQ7ovsgdLcvvaCVc5VE6VrMtFRkRGc0aEpPe
f7LBKG411Q+WWAgkhcGKi6P/cs7yRtfeNUgFcEi9Zibc9vvGQemz12W5g2lhNgEhcER64gwnXwOv
GG7UdGTtBo7Dsq47GPqRPxNGxcVFNLKXWT9+TulcSrJac8A4sK6PBjc7qiP4b206C2k6VPDkfzAu
lu24ekyuFBVn+RPCOEogXRRbeurJgAVHZh7//h9EkYs0OQdnyidBY7Wok4f7NAkRcfxebxSbbaE9
ivJ6oJ/RO074MthPzmW1FIySJ3IHotuL8vvHmzaOiUKeP6nf7NK6HKN3DvI5c1FT5Or3tiR0rw1U
ZrFjROUJ3yWWNTSuPJ8wwBjGlC0IvAaJ64AnuxcdBn3d1R+Xqe3rONUlGpQa2bpwNEw8ZLCwdber
hI9ioE81aVlXbDISHCGVvWhwNIRejnoVl6J5HIG31Xs4KhwJHchkS2mIQEWWQX5HBulZsV9JxfFP
9DfKahnQK0E6XlXiDqM0WF7TCdEkpYxYfTPzy5mgcmYgBfpO7MbKHCHTMEiKcUQxZjKgLs3zohMd
L0btvMChQnViDvHbhQsZm3l8mgZ7v1B/hVf1J+kBxf1v35xCGgvaYHDv8uwDTOYUXFy7riehe1mN
TLzN3PXZonWzDWJqv7lq+lZmfEPKkX6tCM17w5KauyPdnnQmlh7r2ItYy7e9/1QcVxFwu1BQ/WSg
FE9OeSgDWROF74yQ116PfnroGq4esR6zb4LKLkNF1/CBZJs9ORL8F+5SiUSZjlt/+ifB7Q0MXw33
8mx08OI0frujiPs3kqePRvEXkDU28hymzwVt0mt3nTC2ibo0CZHtDlTms14iWx5PS+hhTDmFGzhg
RS+9IviJl/YMQAvqD7Q2Y0g3E2uidc3uKOzT85XapzX/0SZgzPtllw82sqR61YwcxmP3dcOpbTqM
VnthjYJJ7VRTJM0gX0AD58WTxqaaCFIyaxUHQ0EABIM2Yg+8kX1yoB4Jnl5CZAVM02SDPlyTksaD
6F+9QOxibxUq1/ITPEhrX8FyifuUTgJwvwnl2+1xEv124n3FNVqpcCczY72Nx2SVf18R0ZYkwIsi
5DgPBBjTJgBHogKWW5UK8GTBKlJAiSHSxGBLKFJwhD95hpDbqQmfCOYUQPdZYtqPAScGrNVvI8V+
nB6xMZsZM0+IOasRcFfMfTXqFSm85bB9cp21qn9DUV07cpLbOxPqukb3EIOPc54hch4cFwXMJvJo
HjjH5DSU/eG0RvKSY/JwD8W8RnnR7TEdoNS2dYO3bJe1Uiw3+zc96kQyNGSs7njw9ph6z0eJuHb3
HMC2C8LYZIqW7uas9FQgNW2J52xr+UUN3cD21nVrJpbg1SEtIzLR8uqH9lztMu+/az4ePweeaWPO
7bPfjcRv2+5BXr0NtPBjosBuULC7LXoN4Z585u6i+8piDB45Tv0wnzJpcWi+WizpbLGNwO50RpOF
QRDeYpbyOo52v/zO0T9Tl/D/S6M/X/hEu3E4dDgnpDiO1AbcWFrxuf8IaTn6IxpP/HoKHMoTekVP
ef4+t9Fi85x3VaftzlQWpgpYPhtUGFvgwClX+mGNb1Lv0XkqoGiF5xgIV+70ZdP74+zYhfVhk3jK
OOyAzlk4lr7m1yeeeQ8tyL9Pe4meor6ic0IcdaPUTZk/GBx86YlplltK/vWz5y8reWFPN1cPdpi5
aStbBCJyBHhoJs/B+BIwVpgCkahmfN4DoNydNK0dByfokZzb7TH5UKhiaEIt2onEXlg11cfEWFeS
Q0DLhSAqBx8VdR8D6PUfeQcNoH5eOepwiXkLN19l/kHvJq+F/8eHlAHi0r2rwfbCvXyg96joZ+TS
0VzAEPgWG1fhWO67ho8Sqq7NfqwECSiQc+JgAMz6yiWIYAIqJOPKEeTbpMWnJvshJSaTWl1s9/+A
FfKNRKRfjm6IAR0m/ZQjqDVb6GC0YkyjClMS30/Gm7248STfDR3gpkFq/aGx9I/jTcUDTn75/Cjf
dGPGkGqignZRiZyA0tRvi/j2IMkv3nYfz57PnxNHnyKicXoG5Q+J01s9FP1jwHqjs02Mdwh2nvqS
CoHcBeZrVIWbTExBfZ80MDGOSVO60z8Jl9w8KQgFaU8CKV+OA82XhUoiDLTjEoq4SeUxRmbwXt+T
ibX5JaI/FaVS4n1poincVL3Pmw+APFIQAQreSS7D9CVt27B6fZoxG4P97LG0JnsZNvRwOpT1K3DA
cUuoPiDGOxyL5rcl0LMgYvJYHBP0ljoc0tnmd1HwFNg6I0etO5i3dl3lu6ScIBeZVjCSv5HLGvux
pAnFQLjV6TZuO46XCQUnaIi3llA0Qa/gYY13ij2jKtmRnIvcIHN0Rh34cNItN7w81ffq9+cxUUVS
YS3v9aNqXvc223cQp15981YyEk+b1zHeFGowYHyoBKZpOHTFGqPCq9x1kCAek5ENn8b5DF/ZNuUa
GLzLLkY6dIk73Yd26y4ZNPJLjv/z5L/6LiAhxU6tu2E54dN+gekauPVywClZkwhNRiLSpQ5acfa4
Y80ZmGLxrn7shAPnN4+3+JbWmanuZLA6uM2yCP3ZnWkoLTE7m6fZRL7j5c0zR2zRwJQcFZX2Y8G4
ZVwoPcnomi4uaJHButZJUuo6Gxe8nWLbHIuoReya1moFapwHkI9iDbQMNyEpGlc1ZG0kIhE5i96Y
LqreUtFJPZxs+ZRMrXb7pgdRp+qVy/LtdbOGX29MgHHFLCjipBqcmj6FFNt9OVTjLDgV4Sgm4wV2
cWM65yQd0R3VCGV6Y0w0nj6tgaBPbn2S43IqxaSUVyyWOhDMIf1y9W8k+fmXaGiHYC2vcIUaZlr5
EO/Hv9Vk4Mt072MUVgxiq9/FnY00csmvlJTGpVtlPZRFuRxU3BzfS7aqJUgHT141ZTEcGgovwjYS
66a5Kp5dd26QwLVLcRatpHUwTkhMe+vTcIDUeI1mHWFhgsEYoJVQrKI3bH7tR0WwCuMdY5JZ5XUX
V3bmirCtz8vccUIO8sbAssF47oOih6SlvUR9Wdtn58qx8S/1KAOMURT6IcEU2p0qQUSIlLGGxH2t
iiHMmHhePofxcS48/UeaO8YzjVCWWdPPi7SGTAkxcM/4WByyRfrqYmpuZyMksHgwdNqqiroCw8ev
H5SS4nQUBGJdy+9zwbVb6bIpWO1dJkmTUSmUGykoPnLkDIFudMlBURWq+w3TqaS3+uJRsWld6FUt
/OI47pmzssQjEQ2eDFDFi0nY/J4nY+01jv5hx/Q71uQj4rzhaHDFUAaPtW/wpCQmfaOURhLwTNL9
liY+hyWdT76CK8lwaQlrqu6X8pskCl6HkcPK7FXt6TgQzlzqTnp+61l5pM948Yj1lnGJcmqV4qCr
y33V1Z/lT3CTPW4mipKUTPN4t0IUETd3Qe2kHwK03YtqmoAzO0HrHzwq5bDpGBUwJJ5ggprC2N/T
+4UYOwoNB1JOAOnpGGFeuGv3e4HQuA0AoaN01WigKbkPfmKdFVyD6WRL40e56ngEmb+yv+w945up
/DwsHVBFKj6aSoJEnZ+aly/tcQcT9R74KzgC0QgcdHHpahlBa7I+gqC0SgItCzrBhGe0IHPrvDlH
RE0RvCp/ExUcEeJt1nyDW02RGkZw6HFbOZCWQWF3TKf8St4stabBT8p1OA0EXHlhxIMEuXGomEz1
tNIeLoU/8m6mEci8xkmzG1mry7y8DEvUyMDd5YjkXPwqN71oP6r6iLx2ZH/gcusharLCdlR3IqA4
S5wPX8AGqvU3O0SESWEHr7M5aNylswkCtlPrJCCoJ/b3M7trRbbzwkDZo6vXcRGvfVrrFVWBCj+M
BXWarBUYq75AZphJGPFujG+V5aLD5WnOXe8FRAu5jB/wOCkXprQ+fZF4DTQQEXZv84obcq6B2GxJ
3WGYTPBIQLvBBHidFKC9p+L/IWDRlKXZ1uFaGfustbfgxbDKJqU7cSxfiykLCC3PUZavOuV+ygR4
a5kgxthJs7k/VodyfkCDjK9wIAWT3khgXCJu5kE+b4Ykhcjt0EhAYQpY0zmKK3azkorN4yJSHHQx
0U6gDzmtrs9kMHTIPI8ZiA5ufQ5v5RSkkuNhWIKacad8ndlAvezaz5+0+mMHPIkK0zEQhOYMJWp3
VbNyo829Q01RU6ACOfYAsr1Ei8a4Mw2WrALTGonJGPLbCN4NjrnFGbgDzMbT/eceSejw1nSq1sqq
XYGdBwhTOFwPeFIr9WWk0N8I12GGiqBGh9+iRPPQuVamP8WPl8iPhJog2NMpTh5WoRaHoEb6EqK8
bBL3vchRnTKk6gIyKgt2284jKvBARFv5AjnTgsfqRGoXUr4OGlsnnR/3lEoyJxKrkd5uf54KniRM
omEQfV9Lq+LV+mCvagjunIMPaOFj8vaylOwBiTdyQW6TPa7efQteC/twTXSCDnDRaBGkOKT0R3+C
HLb8AB++4b7mXTHTdamfusZYbls0k+bVOOmc9Z6N1oM1qPVVNWgNF2WS7rEpdDihs64c3ADsgaoJ
3tLfvl77cO4s6I7Vm8FXpBep75TkfO0KCuN6wufZSI0foCiHPolRMZia8qA8IaJds4oDsl8c/6sR
OHnu0bn+0pjEdsH867AtYn9UNuLkCwzJ7NUW2HIizNqJ8G2yU0aOvrFX0cyust27eX5C6GHncedK
lU+l7a6xbDQxZ2f2eulweKaFmPzlJFQ0wBEsISMXUYCVx5cJ6LfnjpyFqJN4oDp+niYXCnlbneGZ
Qq/S9sj+9fR+8usFh7hThr84iVWi0x9eMDcs29A8x/7YfCBRqEBUmaZugi7OwTIe5rCUaFsjhEk2
EJdXFe6j48f9DXi1RDzCr35feZGzrM/m7QzhP0bLp/lDP49RQBCNt8xh4wH7S4uvVi7uT7DGFTMF
ZsacXNNgfqtFqGy3jxMaB/dMwuk2l5b/rhHe6vx3s/0De2U/XT9exlXvByE1x59PK//erHt0GIX3
+wHEHLAlYq6hKICEKRLMiP6oP8kXWXtjpFujcWvA2DApOAnr+WxWlbK07gQ+q8g5jxbY5goDiN5p
cLkyVl5eePzsmPsMCZBQjmJDI6s1g/DUkv2GzgvtrqRUXroq8iMQ9tSiDoDxqDJkbdNOX583ia/R
y/iuHRPcayeaguhfJmU/pF9WnzTKxgWI3bOXYibD7Gq0ME1GYFY6WMcsaAogTHGkndEhtUsmnM+7
HcOt0xsAWkE36VgoBK+R3ekEONDu0kWuF0SF8iRReZUHQTRNFWGIs8KgYLg4oOayiEAaruRm8BNj
svk9XiUryQr7pB7tfiXPZlSbiD9CpL54EmgwP+Dml3zbwXnQQJrEcXGfyi1LjDtQiX372JofS40w
Z+AFFEXP3qbj+Nwr3TsHP1/7Oxljhswt/gk6KEyEFO3PQOO8nl0sRf11NvdNHcLzi5MSSNzfeVyo
MjNY1AoCr3mWJCa8CqbtXD/gM/9u4QybU1sI32UQcGlzVbQw45CSRGmkVCtOih+NGySiqiscbDI9
CAm7kAAxcSAKcCijyaEJa1P/9plFz1rZWPcHvRFzQRhxMde7KcOssy6jZ7Skuvi5hZTrsC3+l8Bm
TNaEB4gjvE6ukyvc1nG480KIPC6vAoZ94fYse18ZkegJSpylP1OANDZjJDqOirahJV9ndw/F1lGb
ifonMmbNGhXMtIgsAFbUFaG/jDgv6MovHhb454Dnqg41A26ssOZ8vkmjoqcC3BVu7a/4dvNnf+G1
gTKh138W4/Ie4X/YoEJhx1yBHAsmSD2BzEvZ3yPLVRKoN8b+/2b/SiYDubrr5J9p4aByvxw4RfB6
69WDWrDJj4JtJpQp0nL2OXNveXIlpApmj1Fw4qGr3KoSBXnbF0Cizxk0C4Lwm3VhN/RNndha9bnU
gvvaJseWUA8JQJvrHFX6W+/PcXBJsUQq5eI8eT2R1qHLTLVoseA8nKk2ROxxIRH1ivwAIe7scwsB
ViKC56Lxqdt/nkAG4TbOBLBumo2V60lndwMtrkqdrT8PaJgaMg6q7tbz2a5kBPO4+ymDfy800TVJ
aNX6BsJsXGllKxgyh0VCfoNuS6mVXXIVR2rE9TK/Y7/9vXufMZJwe+iZvV4Uz5vT1AbNgQtsn72j
L89VVKkKXRPig+v6g5SN4wP4FG8wtM+ERMboUbTdTHuI/un4TPAfmAf7CN0a7gnpWevD+DHyOv12
91n5GIvRqZ0wHEz3Cj+HpCsKlI3GgYmHlL3LDxOivZ4qtM9wgkQEVS33IB4u11PXEZkyN2g4T70A
7iq6ZEXhTD3gHeCQjwQ/dFxtMRqw/kpVOGqJTtrtCwgDv0WRB6loSp62VNCG3N/p+xCHjagvfwbP
qz2a7BoC/gvpxzf1Eb5BRnPFzDTt1cYsEh53xt/1GjZp4pXu07bjFkBJI2OazofJZL+UsXKvd+nW
RtUjyH9s51TTpixHVtPmGcmz7ymoy2fCuzcl1FzMjODfUPCD/DJT06Gr9Mpo6KVNQNJVJoAlIOLd
bF/snBZBDtGhnf2sy3QRAY0Im+L3m90beKlTTlk5Zp7I75S/n2RN57R6M2Uq1HGIOAVxIL8ti55t
gsbBwZDOSKQl6LUCxA3cuM8r5occ93IRLtcLs9i7MeDJoouth2MfS346Jp5NRCb3ZXjRVdBQ9iCN
ave75vvdsiXelO2A6fj0mMZK55MKpYM9fqSYXWk7HGy1qjMKj1nkYYrseOw4ixd8e46LtQttrP25
VMJYGYQ3WgKnUJ97wAUWhzryquPqRu/PUcmURtBvOLHepxwB8lFwdCZuyCMLNFi0DFc/Q1rHSa/O
mUvjtJ/EJmBWW6Oxzh77pVEbaJozZvgfYfRRJg1cbk2Lj/7iOi1gaerwcpSesctcEdX+MVHuaY8E
rgFdMRUqEfBpFQGzo2yqA+FJOT+sNTZ27+bcBmP6Gl3ZQm0eviKnouJ7t0zRmMJKIWoWFjg6tn9+
WTB9+mW2Gjx8d6rcW/dNWZpXwUF//IdoD3PX5yqmJqZj77kCyhiATjNre6rfk+eMf1hk87SwJB47
gwWDp4w7jVHV5YJ4RITxHrnuXs86rva5MIQFHrKTzU7TlCdZsAgYnsAsb52JdqcFPELFGaNPnCLn
FDugELcpjk6zdWPoZtgiSCqXrV6mPW/gOOlrwoOOBFE+GltbZn/9v5QCXfxuyJB8hDF0Zv5ifdLS
U5osLHwMF/kHfIvmLliqYXQ7jRz0Yu+Ul+gPkVFfClTvFKdY7Luadt40ziIgAJyPlzH4YrtI6Wlr
HNbJ9v9I4v7hy/v1fR76C51bhYDHUrMjV0FVXVur2PgG7ALSIg0WMNtWWpKib0wTyqyg7tXbj4wq
toPK/NIvQ3E/sv7wekWTXONAlt7d0Qk+ZaiSNp/Uv+GT/V/OZdR+8vCbMbG+Q7r3ud1wh+RPj+j0
dPFn5HVbYIOxXIYF16G0IJwcl4rSHoJtoiMKSzteHf3bigoAdS6J4ncD/FM8cOmiPTdE0Oohxo7c
Ba/iF9orSLCpt2jTAHJOeiiA7Zi7tE2GDswUcopCMcqeWpMByjYs0jb/vdQaaRgVlqI3cqfe0Y5U
E/VrBKSJXYYgB1V6Ulbm3TjRvjzVm/uz3jb1kU0wRSGrGa77DVHqk+NJOw54iSV9vH7JAvBDhjiX
+79bKKq7QyB9SZv09No6mVL1Pt6oqU9jH7j6GxGcx956Z97uNbTtRunV/mxoeD/wkcDBpNeulqx6
ikNyS1vWDeBXx0lB7n/HdLGGIGcugt9ptJicytykoyC0JRIOGsI6It6z+zaZLajRf4l/ISaVFc5o
GYSy9k5g21eDglO6p160JkACYe4MJGfb0BoWelJXei0KM5AS/0mC034bMGcoB09I3M/07IH5/IdL
ksHzXxMv+K1W/c+CtWI1lk29mX/EUGxkuaqBvO9Zklck+4iP76rcf4gFqcKWEtUnPnbW2fIIGzSF
imNkncpHxlOItu/C8VSTCCfppcZnu3DhJv4YPfwoEizeYGxHjkuk70rm8usIpWLRGiRd6xXakO8b
/eTFfvQS/TIyoLuXzS1u6fTSuPt5iGaEpqcsMuGdA0RuZ4VKl20PnnTzGH3eWSa5/ir4sbDPyb0p
7h2q/wNQX9z5//0LSSXJEY7uH7VMan39vr1N0oB9EtWVFBvwBdOFevKJTxyMUik+aQc65o+zsHth
MBfEOxBnYRew8jAV42Xm3Z44rGl2eXnxQkXJsmjLKGk/lSgWuZt7z0f7k1zfbY4JCBMwmRr7kZQ9
F4PdjEgxlAHuMYVEBCt9f+jv79ByvADGFyphdNiz+dLfJTX5By0JYPYTaoDDPc0dn/EmkbuYTN9X
ewaDhjo6FAtjTAr/+YXMjgQWvHnH5wM9Er1RU6WTryyp6XJN049SjvKp7MHIifszPbVuVbpRxDiq
ekuUBCOdC4twAXGTrOdlWy1VFRMjDtNg43qU8xoS3Gau5WvEPQ5qGlMtKCEBN7UFOyJcvvhG1fCC
4GWS3w35u1TQbw1EYpGG0oltIOjTYj1ErOzkj2LYV7UaTkevTxcOE/cveB7DMwodnZb0OkTgUnRI
dlOf6uWRN8mDfKkdn87O+7HGv7Clhfqfp6LDnkBYbrApXT1DMQP6WgqMmCPQW/hTIDdPtOa05fR1
iDNym0gSSC70/Kue34Se3lkfTV8NpJG7VaCr37H5Z88HkhnhvE6vqwKQ1TIvroVoupAtMnPNrkFv
KkiiGPyAnyE0Z6u8txhizwNCXQwEI7yWlyQfIRH1g8HhSeQVoK/4A4Uuz55VsD5zFP6TZPRtjzsK
9PiMCeluWa6rfimgSnOva0yKNWUoVXJPxMwDsYt0hRkNCN3SAC9Uxfwki87JtojCPNRhv2uTGxsM
V9k9ToG6vXVrbwe6+nGlnm++2rZQFmXL1x6ek3s+tG/tRK7R96uUmhXnk7lxO6Q1IPPi9X+EJPX7
j7P0KXGVUVy2RPkbM6o0D+OHE5tMiNih8F4ogE2aD4k0u+m290tZkV0VlVYgxl4uwSo7oBFH1onO
wh0eoeM3eQRBaxfXXa6rB+fbgo673ua3D0kIamjPQPfRyLVf9p82luOFr3ZJhrbU245k0mhoMmKV
LUkTy4IXlLZ3cgZWWTL6OeZo0i0h9AxrCacFi36n8UoU6AitW9Ev6yhpbfFNNyz51H5Iy2AGeknT
tHhgW6LxyyYtVHPTGPIKd+UR2u0EjUx4xW9K5MaQT8F8+RBP23/VLee5aDpMk0ZQ33f7y1KtZ9RJ
BwMMunx6T//TTWUfk4RxL0Wvw+XIeQe1Pd91EEfRLI9/sFhMCA1DfC836gaEUXgWiqyqGMuLqaCl
pTbu8e4LmWR4wUlwJzeWabnT6d7tA1nYvW/4qEDMaF4Bbf2i1gOiyg0OSRHiO8/mmbWNkOQUeqvS
QGZuu/1uDOPmsldSSm03qEA4mJs4rw56+eC6YrvkMLGhVb7p8HsNOIq25kJ2vA5CnLaMKmeeYnlG
I8mRz66x9e41oADJTTl72jqNWgrr+VMar4MQ3c/+9qtFc45A4AiA5wYRj0IBSIwZUQYoikz6dFYf
sq60l8w3AqY7OvQsQjkvT8007DQEoom486HlH9aruwREURLu0YgGlhOB+PzGFsrXhpjr8v33qPaQ
qrUKras2FRyd8ao78TB0Nshm4q6/HbBA8kvjzMz/D1Tq1hAHzIPRj3n6Wrhe8yD9vId1zvPdi3H9
Qo7tZaxf5VCF8IFdfXZ5QuZlk+xFxbjtWbruHVjwUf6hBCL/gXK2a4mpu82lM1n1Wu11wNWOELQH
2o1ltwNLfBtqaGkPNlGtGmKk55EkZiDpKwBCCJaElD9QxA4bI4a5CfVsgUyJ69L0ctNhnhdZUyEh
FSGWHWWlkC694WNd9o96yytReUtjribgIjthtUlrUg1uJaZmQX6kFITPdh44uqLonEEZuktLi/vM
FCmX6S5p5EhpCg/+QtQNr/URuFE/VyyYU6US5cBqXcbrXuPSca6V2D/nm3gopO18gw2WJ33wCxz/
QUEaObtFAM/wgt1ZLYjUcED9rPeAQgyu2VYx8dKMcfnM6siUhRUfqpY8NP6xS7+B6dpwqGKV2JYi
uA6ErLHNVSPKVtPDzctzLT/ydeMKIo4IFkYatkb9dKe2xIXGkTaVxq0EngUecKR3sHl8aE5gc377
H/QMIoiUoPOSWrooptG1iiNYUNcyW5hHpe45oYF8ZpmjQG3bI443exyOlp6W9kNBbfYJqm1YWx/c
Mw5TRg0jjbw5pM+FYIc6/nfXkfclI5wjCcvIL+LReMGUFPDQkhJjrxAGCYNlm7aNjZHDpK1ZgQby
pZF2QU8R4RVZm+UBzBM6BFop7g6PYCevIw5Q05Ka/7QPmpcaHhmCJZ7Sc34iJvzUoP9DYQoU7k1M
8aRqHCAUpCtju7WJ3r+K86KceC3iK6o/vgaTGymOI/SspN2s2XcPCkOFntkBOGQd6oNLBOygYeup
yW0Wj1RPbkR/q2AKVma7OnlMHgN1uNckiXg5QLe4KsdoOV1E41L0muKuX6103VOb93jT1eNEP4Gx
JP0OTBQ685Q8A9hOS9l8sl/4z4p8pfF4eP20P0nqaz4wv0EX1bTjuMNt19mNhZJcgbeON+4S5jOp
Uj9tGqwGiY7e9NTMUWO7TvuUi+FEGn44ffPpl3arKNDBmpqielCRLaV9txQM73IjE9RyMfBIiI4/
zCckA9hTSfusFq4feHPQlmX9h0CmLGDwvvMGCsTINZ20HW8N4rdq/5q7NWY/7wgZrMYP7zVQozxi
NiVvoI1Awc4jJ0hU9AVgIOkOaf4D9lIXGIjETEq754CWwtoY3AX2PzEOVJsLfRoioND7304h2Q55
VUiny8vCqMaoV6N6uaRsGUHuA4ibcyNQfkHr0zvApF13On7m7NjnNf0ML1/Bbf28tJKkQclNFr68
OmIrLCmX/7vssB4Irlg/mHDISWa4rDiwT8ZNLlWjTcjn22qMqXabUrjMC5LZG/5w4WdjrW9W18Oo
tjbV65fjproCKzMDnVUaT0nJDk/MN9fsDvtlV9U+BV6IUMEU4CRSjHNm3E5od/dxeTwX6KncOai2
bUv7JAHGzFuc3oEWWg8j8W3feQiAPTyZfpI5G8s3KVh+y5DZlsZZkfm5mguBK4EBlDnD7wcaSDmt
fRJH1hc8YBwCMs8t+PrX+5b5yMOPHcrx8dp/j4dYmZCfguhPvjPhBlzQIu2o0rXuxBoMym1i9/Gj
LXvbW4sLdC1Tk5slfsCkTyCSxBzhEzF21E1RoMfEAgKVDisNoUZUW1KxR2JGA92yg+4wO/dqdlv5
x4af2L4v8sLR6tMA+qZoJz9x5b4+QXQzOzy3eBj/sI7MwVn/hDPh4LyJp16MgWzm2JqP6+coDi0R
AJYcu9jw1MlP+J9zLB6Dpqrr6Yx8SysTJzLUdTFpMCRoHCUJJ5/ea0AysUB3STuW0BOQsaH21HsX
zAgXHMmYwlMPC4J7/cWkdIiN5vfe6q8JNSocP7yfsEZ/ntQZocCVYIOx81kFZPzM6eZ05j7FCKfM
JxRKgUzao8mYlua91/lMIuRCxBwHIAN29ZHqZlE2Bz+B163kElowxr5jBUP+tx5wY78hJTS1/4ER
+Uj7sSSzMzDDqjMEJlukcJNUZj/4VFIHQOAVbmUA8y9FcQExiY6YpfyU9TScHGPNxIDmS1fNBNgC
+zdrOgYOVAAtJiNzYfeNZh7Uzb6YpDYUZaTWD0OcKgMFStkLrfy263f0NXE1vyNNBsP+8yZM18Bl
I9O2QFBoGircyEobEOcVusknlrnC7TvsuT1ayEm/WunmcgsDmGziu/hPOZv7xVPLS9unOxMaNEsd
XCqzMHMedoacNiec3fkOLYhsqaIxKcDJHXBrPAwjheo0vNlPeE5CU1NuAY5o2XgFNSuK46wbaewX
RmPetHPZUUBoyAA3lYwxU5rxT/5P68BrADqa+H0OKk+cn+jiFfb3FGCHXZSVArz5+mB7Zjh4GHuU
49cgQzJ8F9xRQ3RTJrEjMcPRdo9FzC0h60bPAPT4YCJLv8n0izDNxtXwWkh4wxL24YbFvmv7nEJ0
Q9u1GrXEg3LxH23P20f7sc5b37y3N6p3rP9OWpweqN36cAA6Yy4ycyatBZ8pWj7HY3Zr+c3D5QRu
6c9zBQNi9pXkHJkyadtJ3Pu7XYZpgKjawDuf7AYxMKiteN/eORdm1j88CTByssBbom8S0iniF1fC
Fuo7DaKF2dzf/LWH3OhZy/BRKWpnwCMnjrLuZJ9CMC3bnzYAYJuEcHMBEwDfgHIXu4ClLvuFLRin
U37bz8TgAdw4gM8JvgV20HhE05JArX3KWA5wzA6TZm6ExX5vZ9QWf8ZVXHmRYQhYOWBEkZVjVGMh
zZkMOZOUqukvjqnJd811U3xJjtJ2WPqc1Pm5FJH+ztBjOwHgqcza3O07kBVGhrIiREf1gSJsdVF1
WVmuOvcedhrT1MroKqdPLnS58OihVOT/jxlNPvGxtgTLbyhHEjBSUKZl+GC0AvFj8l3JmvoXQXgD
hkPrJH6hl2fH2AxnCwOlZ2mhfxLX9W+1hJZpQzGZkuhfsATOSLtIa2f6D2NI1rsmrTBZ3Qn6n84u
baAcm+LqMSixNPFsXEqgX98ED6/vAWLEsAIUbu7h4fIdmisq2LX/25gabTEs4jQ5SYzSqZrK+/B9
Vo2JY1ZmrDICrpqQQeWtakyNXIkR+ouNZtzPTNc7aNP+eqKahZsJf1jZXNwkiRPeQ/Yfqy2Rs2Xi
mmnjfb2hnp1oAl/kUjOr/pzj8jn1lzXLbgtoUCeeasH0p+p3UL3lRwJzgXHHZCndjI781w1IWBXJ
ilT74PlNKlgxYWrdjHRnq6Jry2JdP/nLjys5Hs+UXoKgaduZHWwLB4dr+jQ9BumbhZpku+1pXkrT
DkkG03SC8FTGEHrSlbsYmyCHt6N+W6xS58nuNEllWjctIQ+MToox/WvCpB/yIYWei2nLuff87gT5
5PsodY4DoKIjh5ZmRfb4IsDSXYDXN26rToDB3uMLcSf/HbF4nL6Zj9TPS4OOmwbgvP5wDXO6UTZj
5PmDnwOjENwpgiRfVZEkd6e0fmgaLpJEtxszEaoboLxD5nL/xsFyVoz76RhiGXO7Eb53rFNjtC9q
T+rXV86j2b2c2mRy6HvyAnapNc4aDcqb+TOzYItCed0efxbK9dA+bnqINJJCzTh0Lae5VigScGKG
XMaMJAoLB+qwq4e5Q+xfORgt+ELDkTbQBMTpA6/DG7Pp2DxEVWyv/tHcV2HOxarZwcqO2NQNeu5k
iGKuHXIvmZdpja7+YMB/wwYBPzXMCfQrmNJs7wjUectEoETCiay59ozw+v3DNMpy/KWGnZLOqGSp
t717So8O2CcA02qOWxGO3S7HxiR9ihZ60+kM6HfX8WRzlOAos52pMzE6rUfOp+/5ar/oKogSGMz5
IRxufSD96gTKcu7hssusk/26cEfRLchbiKq73eswKj5f/ozwPMRW0p0EeNianhxbxstDQ+zVShWw
W5FQFsZJx+PuROx2+gi3t5eayFy/AGPDPl/8JvW6EKfdKKFsQ+MCOcAza/RZpDYRylM5+Jm31LFf
mYjCAm9yoPxGupH1HmdRRvOzBB0V2JSu3SiYydUGnfYYYV8H+FlBsVjvyWmdd844kSHzELUMXN8a
YiF/NEhZwoA39LOsjY9pcbFlRuyI5q4Z2S2T73DtUv4HkLH+dzHRzt0ZhLkYUVMAZ7aRvHfqvSPj
Xcei2gb2aVhj5ilDzye8QNB8dkk0nz3dHh2rCRn6IvFMgI78wkrDwYMwMc/wOytP2V2/QFzMEe0c
9F3y1jbrK/g8th5GH67JB5Bwcz9aLls9JQ5YKPsznr64uGmiLrgI9KwAw/m6sqsQl5K8yVAWdZHP
8cghPRduU9Xkn1aVHthe15Y7E1hnkieIzcEZnEMpxW7v9f6y9fnbhVTUB47MEOR0koFCntfqu5WJ
j51LNk0F57OnGYXSpo3y/1dlVgzS+CFSXwDxaR8aiNmz0jzjd2pmQ6skqwc0t78jhz1+Rvj+Jhno
jDcCGZqtP+yh5l1Cek1OuHx/08B9/z13L0KOabG14CCATFLPaH261p5gyIhQcTDefiwIRPMbHDr7
3T31FjP1/rp6USTz6LuLViPq6F9RCfMGLqr1ADXdFZyYA7G9Q8BgLoZJx2+tTMZVdP/NZAtNF9Qo
1zgbPlrqkfxb2LXdAhgZVT3ec/JAlghR16/EXzC3ybjmTvN9WQEMY6P+5oaQEznetMXe9QGjdSjQ
yozWFK+v1w5cPeW/T9gb3fU1u1OfusqwDz67Rg6QD/ExA1s7Qs0/+Qb/DzeOWisUSFQNanEARuXu
hiZfFnMzh3vmuKphLnOzPUZpt8PyjwKN9lUa2gDim2Ih+5OuE6dPYc4JtcKRoWkZKWLkjdXat1wP
Fnf/ArxoupNsID0yoEZk994h5JB0egrgevjXIx+bQ8KUkI0tHk8vrex0wxWKyIrnGSDh8IpLRw09
vKiWCm6NXBOgooSK7ObxpjnVG+grmuq5mauXeRitHLob2YvcohO9zOQpxmJG1wlu29gsVlFVOtE3
/JCMZ2rh6jsN+fCdXlK70xkbLNFmhQDv5bz2RCEDe8JsMr/wuCEohQeD5ACy83kj4L3hyrivXjHF
grV20eMTgRmpJVaf9MbDwHEHGITAKIQYJCslLwtrS/SWGx7ZhQw2sgOXo1cRdVbPUxw356GU6qmZ
6k+eXvVtxfPDiAhuXqOWhh+hPbsdY6gBlJn7/0cgBxUioBP3QVF1kCh8ROFTN7y+24Gyxf45CLCZ
sQOcDsURr45tVHXd6cjfND0XiriCUHm6HTILGRvyEgarBz9CU2W1hs4UjEDKeCPsHj98yZQp13I0
nyEF1wYQPUxszM1qAXFFssgRx4vF/254ZGkLGB1ayKzDCPIwfvRcTY9GK9VRcRxJMoXjIlO96CQY
9FwtR3PzT4C+ZS6Uww+KK5Ka7XTAK4f4dXbHrWmTMZM4KPhw5pgvJGlouOe4dzA4uyUrHJzxO68r
W603q2Kfj17VY24l35xqkp3Q0gZw3D2u/8S3VGyqZhVW9MwIm2c2nOshLoPYPJr1ljyM7uwM3IFV
r0MAudTqV5dyb5uLllEQo3qRPVc6Lxb/oSca6Jw30UVl/lQRTvsvf2YrXN8JDImwfvt0DdDhN4nE
KZxL+BsT2nO32VnG4zb9yWwpkYTm+aIGz99OcTrcFlA/mhOtN9QE3Pni97mf5PFJltijXqABrpVA
Ir4OZotto6h63N33OckzV0vl1Ca88op4ebq9LZoO1NMTD9K9x5chifSYdpd0V5UNEEAjE0jBiZM6
P6X1IlA/7lBPi/aggBl1ysfBrfSZuNkS7nYAsG74CIxnxizQE0kBhyJxwVVBCntvJomkI+j6KN0f
FiBeV8/k60MZe8jknC86ZhIvZkeWLe+QdPi9n+JfAIXE+3UjR60S+OrcKBzpHUqEOT2lKuJrdwtV
bz142DKgdLL+Xu4IHxkP2Ehb3OZXDjHGCLyF5dbh09WRsNoG42HDsxVwJtGUN59b+krJ1oVA3LVC
Cj0+Gdm9WwWlSgQ+8XC9yOA/wvfamjQ9dMCMFwQVn0vflPO3iVt8YhC+FsVbSbhl+PzSroBU96wS
xq0BYLQImqt9grL7HYge60fs6l0vNFGU7SpgusSUFYwCkFHsrYTOCKOaCnGk7fq6mZ8fAkACl1VB
Qm059KIpFYvDpzfhbutluFMq6CDYfHKBt4fB5E9vwYmqv0q7oG4/vecX/YnQYBE4MvWSyC/xJDLN
X3YrMVE3LAbSv4+Cs1v8PuZRAhXyNu9rfJWDbYSPZ3jKTq7fvUfqiU+XvEMqrmuDmXB93jFwW2zf
AVrrcVA/NorpMbC8QuyteTgSStAArC7JP8S3ebePHuKH0jKQcaBDVC/x7Jfk+hiNlR32j2w6RlLx
rRaA4oV3qDUGEA53VOCGYZB6zgV5+U618Q9V++AKad4RAaQYMDlw+/W0OIoufFcGwKlknwy5k46J
VRnEWLF3KaDSBR5kExdkZZsZKh7bbLpXAV9HKi20XBJUeNRRT6R+LFBxRfakBuz6O83Paa3LqoRd
/ukvwUvvmSzn86vasSsiG9huuh+0dSJuSFimc+cPff7kTu6XeWETaj8QoQyyWagHezgKfoMSpTQ1
MS6kOyLxDaqH+aCOPtRP9ENAgg1Gc6xKXjw6WmM26eFgeJnBNwOt70qkymJhRWlzoLfzmWyOSiNl
GVzRAG8GeDrFD7KK523u4e6CUm32EHodvqUp62GfqHoSCDMHfPmpFS9Qk2obb1BtYuVPanw8Lp8g
6Sdxl6LG9t9SAxtTYtqEfL4zoRZZOKG0mFwakqsQMdIeUQPfRBSkwM6BtcQkFn8iapdv1HmDqSxo
RCaHqgtC3GvOPPV3XBIyuGQU9ZghRMcz+OYDhZaRDf7GpZi60C3JmAeQ0LK7CoZvWYQF+26XEIA5
3rRNTvMbSEPzSP6pTBqcuPyW3VQ5yxvWsqpEJO8IE/kRMrJ4xgKQY3sFGr7rm+daU9BvPS21IJK2
cPn8BUT0bqjMLv8/3tRl1ncCJ3hvQI8NOM+PUkQ93TkqjGUGYS6IedhNb1xy2CifSEYsMXLKh2dS
/aOUP7/vbmRJfH1FNQl0Kv+ZTjfBXRMHQnAoOESgN31KayEpBG568g9wYLKyrelh0AkWwFnrV9Ls
+hekgewS5IIFBwioPeiJL96jF2JZo0uuPj9GNhfpRQEpsxPv2Ta+IYE90BNJwXQ4D/q8igyyuUiD
+DfNIPPMLkWH+D+AxfXdyysyeZMWNet2fnf0nnR4zRW0Qz25TesqN0XlZlbjHES96mnVDzQyY2Dd
PL+f2xdersG109D6nOs416H/e1BNcr6JWHHYnfS62JRFqEyz9HRKjmIuXae07lJGN9bGq6Q8OqWa
Y+OgGFonUgg/joTsi++fi0mepGaM7pbsVFblAwWd1Kh+TwLduW8Idnhk3ascfmktfYuIrGiSv0OS
QSMAO1eMDSTJAjybc4w48BoFa/5aHjLp/P2zYuRZO12F+WjNkqcTfVSLS+PruDzaIqpXkBl9epEm
ebnckakuNa5CNiEhhfbI8kYqNz1p1Qho2ZeVXaWaJSATqASYDyvAmd8HP/8clFbCJfYnwG4wf5da
4LegALlvQpUjXNbiyTX9V3ChfeoitpdIOcnLCmdWmN6yNHsKSZthsQ83FnbV6/l+JpsQ9NNAEhdG
IE7FBqjVMCord9OMlvYKXnPKmN00H1vpLi2H1dqKezt0O2MLi5cyb49Hn7M5ZWhL8Nu0vUlRPnAq
3Ou/k6EAXOzVWI0ruaJaAkYcsrHecjrtbrAFpHSOMRjstRP016w095MlOWKyg7bzhTqM/3wQKRFd
RypQtptNna94GxG+dNZ4mmDczg+6qgYhQyo+47gxxl2vc7v5sxMoF1fEYogSmQTHqiNHmqNkBjY5
HaDIowIvpSiilvplBFteIGmgaB0q9wshr48l1XV8JfqTh2Jhgr8JVMgEhkeSk23uz13gS1Lojvam
tUj/vCuqyO52D0Qis40b5s49GZnWdVc7p+P7xH7OyhXN8Qa5hvXxSUxAynphO70FH23f4t1qPwBq
fQD9dpT4XG+bXptTYMR7GA/daL/rr5Mr2MT8bntTX/yF0BZ5T+/lXCXXD4B2C1a4XgJ0cFVotiwm
g//ddtFN3LTkhiRl+z/YkFfrJtlMHvd/CamgQhJZT1VNO5C7nWsHa6u6AvR1mG9oCS6+fxqXH28p
/KLZ9m8Bj4re/eN/EztugcOeKWSTocaUCUjhBJ+1jzH0lCq2FZkNDz9omSQb8F2nwxTdl0q/7/Xe
OVWX+a1A3EAsjuBXhWA1i3FaqnvSogtO/LCEipFZqmZKtsmtO/cBV8KSCp0UxUCas+iGemsX7kgy
SVyA7reQX6yuRAAJasJOa2wzAi9Lsvu4xGumeRW+9W2cGo9a331nAGl/OChPP3plUN+wAlONZGE3
QiJCPy1gL8fsTF+q5AkvyeH+RdMqc/hWfImmuX+rJos+oJDTvcEHeK5QK7RUCE5P0LdF8KA5m8JF
u5CXAPLMtXGHKSrRE/BBbR++I6eDhxbs9AfFvpyKaYaUb2oUSjivnyAAxhvpN2CBQln4lCyYT+Ta
gicEB3I42m1UrQuDYjtF/AW9vrxi490ebFRaxNMMOGukJBKiTJB5vZOlZoM2xJ98W8OcOQ5hPT1T
10PB2HYsVSEK3GloNy/zhT3x3HCFH1LJHEHsfuenFefupbWa2fQs5/eLqPvU4WqM0jn99aFeF681
I4+aBmmJjkky+woXaVDXXpj6JJGLiLX/IokWZk1eKeoSDJKm35O7iaoo+W1do0Z53J7nQaf5wqzO
aNWc4ADj5hUG8oxwJhR1EPea3AdVhukzjlLWSHNc3EMbnmrIkxVSLFdEn5sFF3XxJsQPppPT8/HG
UOtqZh/sQijbL1xob18QTwTJb2ASHDJrTTxZOhMsWKcK8t/gPxBpbcm2ZPVLq4nuNjY/5HBfViyV
gJUNKRkuQS+9MQXUqUF6RCe4hvJuEFt7moZJ5teSqKwCbzgjVku3FYbH+Nz2S9W6L5Jykull2q3l
ZZz1XeiGR0po7Yjmmc9/KHNZUF0REdCMEAjfNlnTu8Eae/6JJf1WTedIvJFpvo4ifVJ3T5XvNI7C
Ek3tAVDeeQCYqX9MITFTX9WPVDfIQzqwdl6UX+TlVhe2dUxuYGVPT+sM4e0PrHZvB7H9ZOn4Ka6X
eoVIuUo/hCF9hBQvPm0LVEuQwFn92o9k6zdQuYkpw0MOUxIy91+SzshknANkGFUyOOIG7HLPjd7Q
D8haY52/HBxc58HU8xU9m/WD4+BluAlhmrWTTa7Gi3O12ijsCbBlz5K14avqAdIj/QC97tBFRQqO
ZkmLWeRCCdYmCKnPas8Ewm6Qgv2pgx4dQelHJUSBruoPBCGPVIZDfslHAhF9lS5Tz/tBQfRCbIKP
qaQzN/iu024YOtQCbABtE05divbRJ3rH8DmFHqI19JOikdn1mUe6cR1bPDNrPnNvqvhRu/w4O9ti
hPJFWQyaJ0TLcLyBIZ7hpC7+YIGMgZPFa9jtvWzSFp4WPqRvk76DpQf/krK2NNjbPN6MxkVB1/eh
UzSBtxWB8GKRlVmP89tPdreoF6AMDcgYENvA/fhsgB+873/Mz9jYQ4pIFTLX3k6UTxgPj3UoZJ3W
atE8cQq/nHEehQJjNLhwAhWzebUH4lQ22kNWXiduC8FlEk9iQGNCHcN9ZgmivDWqMMJArvOpxDrk
+oO72iawybWyEYByptmUpDCrsBw41CIplhZ/ZQgQ4OU/2dIM3j4OTlSPJV9DtqmrlFEDGmdVPJxk
GKb22WViO3GnNi0Qfs8X/ByUqYYfDSzK3GlOJXJ2trltSNmy60XKzgQWBtFeFDAGSe9KyOlrNfpU
KhZRc4hikoXjyf0GAwLvGHck+yzDrDUH/Rmxu9COqV4nywLsNKc4rpIt+ZLCnUzW8kob0jZle1jk
iQNriqXk/zDkmVRl338IKJjD4C5U2mnCWHleXAwFTCV6tnZYyt0un1Qcob6iBHCQaHLt7BU37UVa
fkEwGygzQT17QwW26fi+F2SPYNw2A9otT439KgmUF0RiAPx/OLAwKNu6qjBxEmi99R6m1lqGdZpO
msXi6c15MyeSH+aoLuxrOP2SN6eUBmiVVx+wa+ejimCT4RCI0GnWVfptQMAIucVTzilPRcuKlNqI
6+Gxrtvmgw3ySZ2jygNIPFQ5tkpmohFECt+ow/yCmoi24w/0WueVnWIvvl/iZYIWwfepFFIg+BaD
nDs8edadef3VwyuQ+4hIsnyKiOp1KMiU8df/Jr2Oss0StIfc09eNksRpCUMvky0DWNkR9usECV5R
SbrpK0Hjfw5wpy70JnVEEyDwmGLspB37F2vADkimPgP4IECXO5xHOewcj55lih93tjNm6Jbxsp7u
KbhAJZgLDsHVg2u1h6D+hk/PWkXXdnTLltMkIogAgYxzV4rtQuL8RPWE9RgzSUuRGHq8zhtsjK9d
BdocSEsxdwaSSYjcuo6yjooWIhDIRzmTwEH9MR+LisAMXywBNqYuOacGRtPqGt52udpCzA+yhStN
xK21XnS+Crh3LDViAJSDsZVKhe+6l6bftBv3pb+OVIDT5EY4isBGMxrs/GI/A2xulh5UTztUbSae
umONvNHLPCJ934dzlVjLnAKVcVlsh9cxD1qFzNLHu1cSQMlJEjGxB86bf046aiHHl08pdrhdrRcN
s0V1jCGszinXcXKo/FTQxdXZSGKduFFNze49ztK++ZamvZFO31/Zy4ykit7E9+kDnEXfG8KgS6dF
Hhw78nGGIc4qbWCJ+GzHeNLlbMPZ/6Ifqu1JXSaAEObycn3s9Cnbz8QjRt3b8lbVtB1+qi+QXtsY
L/CCW7wxa9jOJdoFp89AaGuogq+Nd/jyNzO+iPEoftwALmmxWIx4JeFHbXcZybQ1/TZGPW4Bu9ZI
6S83p8p6CPreNpfYDxgoxIKpmYf7XfR7bieX9h8xKxh8FtVqjlzsT1tzsFXncc6/GYBGbAgKgCWY
MJRFTdMLji8dNFsamex9CICM2HlAbgEplIRjCyAU+jYL7jGIgcaGaWXiRbUAGzfsBsY05bfL1SET
KkcpIhXwHL8mzkHhLpqJoJZ2Rm6guJnAkAC21cnKk2Ak7zG7onTLEDFh5kgLuCdUIt23gb9CwblO
Yls04W/hNeDiOJSNcf/82O1fWG/rIJQiKgx/fyPHsRppZzqgZDIYmmx74thBg30qFE/bjcbB2DGq
qQfs8y6u7ro7C80FCYCRosmTD//DGsbXJUDfjJ0Ls0VQldzw3Pmoi3TAEN+DjVLZcGTEWX3riDWx
n7swuDhkwvvd3N5csw4CrqzgJWIrlgMcy7K/v4OVf2vRq907QHfnBJGUcg0PdNLEp5y3Z7gLRQKN
9ZSx+8g2GGBEOASjOLwAdtWrSoHKle4YmHe6fEd+qiFmN2Ir+OnusMAQU0sekaeVlvJcXI04bzyq
4hiQsX77guaaMJ3haHQFp0xeCftrM5WzKtY3J4f8PbovsJMj2B7Wr1Pk2SKwNwHTFJaglaELVhgp
r4qhXdFc0Bhvo5ofHgz6SKFTgrNjLSkanWXdEsIdetbuT+be9QEz1E8RVwO2Ia+ryX4oywlDh4Gw
6LazQijKHLJo3vvMQM3pqZouXGeMLd2cGiUJN6Ag4u7gjhrGL4p0GPuM7HpEymbh4h1zOLgsQz7M
t2To2AymjLGxeGMefb6t8y3ixYMTCwP2/Hknftn1G3TkvlgYxJ4sC9vZ7K6ks9SgprCVwOFTICB4
fVgPbWl23oLyrEWcV0Kj/XoJ8OR7OXhvCPMDrbIVPA+oP035nP7vs8oS0MNqLrKyLNglrIl8XqSj
Y6D7MImwJWTOp5PHXRMhMvyIiumLttd/+fGkhNRVI56TXNSaJsp4mCjhmiOLQEeDUWXUHyqG+TRZ
PWITO0QPc3dhM0arHKAc21fT8Wf2FS1z23TyeD/fnMOo3QRmSA6Hv9yraU3kkAfwLQldfsGg2/y2
o86MJHAfpIIrEo2ysUbE5PlsE9wYtHxBi0zOmY8BKRlzkUPYHW83pPMYGMV9rozS8bo6AgSMDnTi
g1+8xMNOjkaDOMrd+8Z330H0EuP4S8j9P0zM9xQ8vAKWpdBFbXRgj4ioTCU/CYlvfmILrv6mQv+R
PAF/TjCg29jioE4pTnRnZrvjoobKBTzl05g6MkZTaZtzh+d7eCz9iOlOaeyFZFF5BcKTHV1KRpwa
ZmUEy5ibw5R+U5XLf7I2FSEhRf3GGDg5RJWJIrpjE1B4OskFo7zQS6Zr/ex1pjPiWjPHC6fid2Dy
e74YdYHpw1/JF5TEH8Fco8blKxqYmVO9LowsSCRyiX3WZ2/LbXBaYGoofnU3W6M+fuO081+Geetg
Nwod5JihG3Lze9tMdsyypIrO8lbxTOPFhWsUPLmRE+BM6gPrGQb1XEVBvY08jOQjYauVxcggJ81K
KEuP4FAL/ihd1i0ptVEchGQMZ2vQxMWq+60aEKPvH825kwaM2zudkvF+8fIVA4Y7hwhLZRCvf58C
Ig7Bdz2I/e74g5Nq0ZcYwNIa7G0nq4cvlEnWYGvmqES4NVwtb+hFJcSbVSXsviy2GqqMpdmF2fOU
pzFjhwJe+4kbEp/FGuNQDTPA++/457be3WLTcjbPySMdXHbK6cRrj0z286hYQqjjZ5J6s5P6MbWc
pIHrvhTLlumBuN3ElqexWOhLuB2lhjxmAy7yMdVdixAuT5qSPqDMTYEmAJ/kqiBHu2xDmMVlL2mM
Mp1ErhZNj/tqmjRC3SFITw+wX59NDFfhfd82FxoytOyGl4Lz1ozWF4hkQulAYy7VGRo5x4BXRooE
LvGTvicf1sVP3FgeBq4CcyxrT3DqTMpKAXpH3YvUFOC9Ly7oRBcTPNe0ltLMfkzifLhZXDq5YtDb
/R/6hCl0EF+85MHX01ENcjovTVT38geZVhjbHPc6L3Y30SzpwfYCjy2y5NvsgXkwgqR8xzRRJWFU
3T5WIaD3jY40pYhtm/Y+uOQoeGi1W547JDBc+/dNt9qtGgzl0Z1kscdEOteHspEyDrWjXqfI8mXV
e0z/vL00qKkpkemCCd+Mv7hwZ54rVH4+oosXAFisFV9w7vYqeiJQ4h1YWtBj0Jj5vGRc5Ner0MET
ijm/M1gQgUARLvrfmKgcLHsadkM+MhhDjw1kR65e0FH+xsTaVaKG34T5ME624Vvw2UkwAAJXIx2n
m+/y3lKkja6bTU2lc1QLob4yQhXuggXcT+4Hm2mTEUhzhUqeQZI9L6MiMap61Rb7kYJeGkIpPzCy
ZnLjyJl6hCY6u5ttTEb10YxHYd7uw4jGfwR8DgCSAZyawwc+diBbZfuFWvs/nvc9/HOiQPjJiN1x
ig3F7lSEqKy2XuXExEB8mFpnheTGdLgN9Dav7+4Jig95MVACFtx4+MyFSaMxfJnRBTx7kJ4wulKu
mtwqLy5M0y83Uj06gSHrl/ErQwh6mGa8l/FwrKJwuyqB588s9quSUQA2wXLaKJznXxkbsU4jncH+
M/RRo9QItOsi+/texczhgUfB39YdARwbgakCzrOs/UYVER7BYNOofKgcCQ+7kMrQkceSfD7aXfF4
HFo74GY2Tv9Q2b8nOMi9yoBQJVUzdlVPsr+vsJ/p4f1meIxRgq2xNKsXYs+sDbXKocDhFgKD5VyU
1gTBxlMR7ao5vHqgJARBTUP5g370p5C8XhZFBp70lgiO4+pGN7B2/GC0phaVFbWViXnJn7v8Fefq
ZfHmUDxwmLV8i0Vbzp6HuCh0XaWjBAh6jxeqaY91li3f3bdCUPyAPekZQ2UnP9RifB/83YOcEciT
jWHH7ZqBSJ7g+BsN5r8qHuVny0yVuYeaQsEmRkEqtnGlnFzi8nLSet5x2e5cecIWRZFKzVilc8Ki
OAxjRxcoahAsCSlkAcvK2Rrfco+acM9mTvAOve+5qv/5oU/FUXYZ3a16sWPQHN/8xyz6dsXcKlmd
Gi0dMjdpZYEgD0L9aYbnNs4D4tqVIXyOlUj8c0hkkU70A6ncrAQRfS5WdpnOPeeUUsAc6IpN7v2i
MPXbN4hVH+vXwyuUc1yK4MCebk4jdSx5SqJhGVWBxTyxRtohlKpchunMOhQxs0q3UiBAxJi7JoFD
4fCLbdsxr6Vuz/k5LWwoJFnZPpYHQuxcP7xBqikm0ca9Y7eponvEVvqiS+0EOB9v91fcK4ebyhZ/
KsQRjicIfgPnRB7QwYHNPlMl7KJk00RUHtvJ9+iBTEO2S80+AT/1PbWglV1SG3ERCvY96ZI/CtZJ
XqrxkST76Xdf3zK3Cp8/UeRPSp6KYGdvftjy3AgEA5GyIUz6+icGZMdt+cLkDH4utA6d2ZzKcOI+
8hlxR3S5ULEYh1anxdgEPB6Uia/RODH9tN3hAM+t/r2haHblxhGqrdlhu4gj3vBzvK7pg666U6zg
G70LYopegX9+J6Di6ypq7tc7YEbEMXASfSJKajD93Werl57LVStKbMNtp4bFwzHUDievCjwdHVhT
VzccuV3KAOLCFIxdWydMCil9OAOECHG3OywfJicILAPn6Bkxlgejyqj0uRNu4cCqEJGMevKJ1X+d
/DsSYAqBZaNvO9MoWAcepfySSKr+HzpA0cRxRG1fdAI6PZcf0B2Q6+QEN8hWNU0MJXGv0A2xzoOM
FEHGvyisZamNGLhmvgL5ZBgAhoISsh2krzeZbj7tDe8aNjds53c6vlu5dwpUlTJAxBafFzI1jNGy
7Upt8BIKAULWC5xMPl3pRrdzoEyG9bjFrG4Y8jqNN21+0V9bsbsUG23QiW+DdXgtPHWrL5tTT5MW
Ty+V/AOK5YI5wOZm08rvk/eo3AmjF7b2qCn9Mg5dMc8zXVXyTY8PqxvOmxc2pPR/3LoBk2+J6Suk
2Ggczd2Av1d/rXrP3emjhs6a6GioEasyCrCfJMqQGF5L5mr+sTgsedq1RCC8jjU01mVvsTqvOYuL
/xjFBfDWR4NJz5CISs6ZZ4CRmHGeOwyhorwaNPqn0ri5O8PJTsX4jwW24xyho7TwsSFjvh8G4oHT
Q89bp3X6PROJ+xgH3X+tAtWJ+OlgojXKkI5scAtaY0POoBMnIXI8zBimbQE/122TmfX+9lGJUlOf
fwf3cOoB1oaY3HJdWJ8YqcE9lt1lU3e4bYwWNayhwhpzBh0/HAcAjJRO+hh+jJgCMdp8U1TQkhRa
YNzVQ6jR0Yi/y+YRQnikWPwxB8Bcy0OHrJHCxt6EpYNqSzXOW974qabWFghv+SEGlczg2+Wk0XjA
8AhGsir6HQVnk9A8BfTX7/xYCZtRsG1XgmgLjIGbjtG2gvTK5nbrsj+Ch9WCFCRewMkbjAraYCQ7
aXD6Jrv1dKEN36htSvMeI38h1Ecb0fkpBbb73jeOzyN770SgWJo+G4oZKs/10QHs1u0ZDEOmB6wY
7q7R5AnPqva3WTunWWYhNOvvh8wn+VFT2+KIyrn/Wr/phw5cyTBLvKwOquPGAwtDUgkzG6QXqfaH
6EPpPoLT6T8r7nxTrvBADA4/ODXAfQVxT9fx5oBgNmtg+BkyMbZ1rLJf5Cv/9MYnO1eESlCRIbUo
iSDn3USZ5YJdUgQpZpLWa6QYi1jGSpv5zA+4sLNa6KnlECL2cxP6yX94FlY5XMEKAiNAJFGKErgt
OYSmUI/mZB0xK5jvqQwdHNt9dY3E35rh39PquTslvqSgt2jJoAINmz5WzYGqu6g5ge+OjUEiqO28
Zp0fdeGErCrJC8PCgYazxAb3rW+6g9zy7uD3iKaUGE+gw5rZXxrzVPklnGgJhcewcGNvYNSD7mF/
sUMFusHGYXqSV1TC6VTDUPNAmnrKbKtVf1H6xjHAkfL6I4FtD3XCCd8NRW+NvM3+iAjIRKLGJUnt
jjy+asctHZ9Sbl4RaNHoogiXZ5TPjluLH3RB0eSGVa7W2jqgvjZyG8CMDd+6FKhXXHR0L3DKS+6D
hh6MklPW5KeyrepIhphX4DNneUJCNYHH0hnqWjD2Y3Z5DHO+2OOAqPECpOq12c/AbXLcwJ+UaYyW
JJ3ebxN4i1BJGQdVMQ8PPsLVy3Eddy1/vJcE3gfCHvAJIWHw6b1z40zkcU9Ymn/QwdYwCzL2X5H7
6lm+B0cF9DDvaM9k9rOG1dCx+TvFzQDcNXLaK2vpY2hv9gTVtm7B2nry+j17kTI6/ff5AmAxpMUy
h9PYJ2UJGPFLId18674QydpMg1raereaDIAnKAWVJtMlFVyrhRFTeauOmsBlwqIB1M20ClzByKdn
6P5JXVvF/KU8gdqU++S8p+wrlYMymMq562jYWa7I7dpjApz4hrdcV18fpbhmUY0pAxVILSSvNNBL
M0VqtF+VkkbhnGpU432c6ZJ1RfVEq6lBFvepGMdDr3erTbGWXMvP6EuHq1Ha/eiQvWfBqvAJhIl7
PFhjw3ZI0frvwazzCBUZkLu3ibHZa/vM7sDtoTRx3FLBWvJnPoOKTXgHC0gucFdYmukZk1AuPqHE
LFaABz931800bYl1VDxggfs1hOlpAMy5ZGGBUFqB2v/4+b0+lW5ECAgBc+vaw8hO7r3dGYy5RWEI
M8aHxurRa9ie7dMGXL0xYIr96puXVWIRf7myrYXl4RouDIfROiefoAhKzXuqTSDpKM8Yh/SStOC+
uzNNEl6I5MH/KR9SaxPjdD0eg6CST8O20GB6lwiYhWjbuk0Qb5BTqEv6oQ7DmqFfmBnCPhi/7Qur
KtMmDSJbeuvZNeC6QpiNPQzLdzTY8z+Dbog0DYwzRnzZ2KxkVARiRTcsbH3ah4iqbbLiNQ9KWiNk
AeBIcvSY/KpK11aer2r/s1ltG2jdxm7AVhHX53nQ7PDtOzDLSMpr4ek3rJY4b7J805H/slgsYi8z
ftogoRJxD8fJUATMgMt8/t5AVTloGfmSwlsVhJBSc66SGiIfEar7fTcQMhKoFM4iWkenwXXoN0N7
bochZmzmHHSTySaRDaeQaYxQXSUIhIqfBtr/jNCJNor/bamOianFThHqEqLx/tTfF4digK0GsAN6
TtuvitUhA18glB45V7lv5yRBf7sBJ516kC0k0tqmcKXFRMU7G9LARUAma9hLeTjo7W8RrtvX/thG
ElDboICBk0PRfvSDXAa0pdXydFTfCX9F3Hh2ctl9SoKbot6AU5XcAC8OfA/XJwsOHY0JKPvlSuh+
myyh93uIN+4l3P/Nu27Mwc9XOvwlSdyhohDtFoheAxXMHU6U4Rgq2PYhzEOmjxd/XDgg5W3pIuby
7USX1lNDVCUB27haLLauw29p0M55ao++slAVlStzOWvzJihyUPKZDQXqOjtQiQmcVzeVQ985vUdp
VUQA9VX7uc+c0rhjEbfjdRdw7gZD6LrREtVEWP5lu8oQ9CasJqLMSzGEmqcVsFXNrj57rfnKlk1W
l4+mmhig6jYXXFj8AOQL2PxbgHG+7MUQLkDkrJOiAPd+26zMTggmuikZozrYcZhneUlyzS+MuLu0
nmJOhH42xA1UYszJagTSNXjBWfhA8RI6mFOSDiQCssNYOhtnSB0dRm0En/hbnaoI54o69CQaNZgv
OguBRS73DRRqtQfBAOv6HHP2KkrPUtSu9ZTf783gFDDpAAQljvDAc42Sh7hBWd59+fc2HJ6T9D9H
e4A5BmxLWxbysPBmtN58DavavksSsbSTDMehPJbm894LHGq3eIJySZKaTUnI6n5Zj7t7MKq89YV8
WMXc9pRIYu095nFsfUF4dob/o4y+qomuzl0B0xfn6I5KK3UHUqFWzC6Wg0VZXstkP9ZNG+A01uFW
sWA2WrMyMepV/HUjJ6AeoUm9Bky+XSgovaBSkfKOqsWkyybFqYi4pYEypN76flZXHqAta0Zfaj/C
NnzwNDTTZublqsE73h0G4M2e73bb7mzMSsQOWzw6J1OCSEfNpFAxknfonmTS0s2xrItfkkHuhTLn
ip0eRQCtPIZW1IKCfV9Xl85Fxmby34NMZAsyyWdfzO8lbt941WmoHeyPUNRn/VojXEOGUWTbg51y
LdU1qRe7lXaAPZNfznjVJAQjkEE8h2LeruTe7dHL8rfNG9CgMpIhkrO8ioL6CJkGLm+6fOG/3eqZ
mtKecsjGubkroIRdmWIZq/YoPPV1x09N6nux2h30nYWQ+sDVMW+grQ6yNlkMxA8kBzA2pB9VQbg8
Wylta0r0pmPAV/a5b5tJlFpykll8NPKVmNvkrTlnImdWpfYM9hMw0Z/Qtu1PRLAsKzjVVe82SRt0
Vuk6a/FV+bCiOeFlrlflbSf8pHOysln0VPxt6EgvoBwdEA2q74eAZSaO6XDQ0DGxdUAoMdm0rkpk
ou8AfOPGBixPvCmbLbpqCYbYtei2WYp9ocbiOczhbLT1+URabhFj5/nJEu+/NxiSTEoClZYIwxyi
MY65bd7fsYwVJt9aJ10DMh+AZprjDtvh5pVpdeTlec+p22/EcWeVEfkEDFhd4HagDKJYau8cgeXe
fvmG1knzy2RhrrFBbBc+rK57DejvVOIVDeRQABB6xfl6ZuINtHT3LO3IJMCCacgy1OEgn0I6nrBB
DouyblZm1v5nnzjgUnzMI7q8p7jhVR4+Kdl0BPtw24Co4edp+MctC6ovoSKW+hQaLk6FvkZ/tEXG
FuG/ySoVbNLgtn5sx0VWydzp2nIVpG4Bcby3HrQU8KIdmvJUxlUStTxC/DQIFqbtbAsHI8YVul2X
ZyLa/A8Kbeq07Gmk5tfJ+LJMLU7tHMUjIG25aTv1ol0UAByCOa+Eo9XkgZiAmrWgmXGjbh3gFj81
twnWDFDYavnnVDGT97dUhYob0YPwP4AN09PjjJpzVbQRlA8OEaciIgFzSwV78UpI+FiUhEqpEd57
zJhNyYY6055VVP+HTggees1KrxS0s3pPTnj8J/M4r+c5nrR/jJKmGZ/WVgtDfy4/pAlYA91dKEBq
MYkvAaGA1qHLS/kCAL2AICCZr7kp1vIHYygTBxoeLDKt3SOycB6/5AW2BNnhT+PYOw/dx5F56lMO
Oq+fh1cAFrPwAlDFkuUBE6Fd6bpDCVhKqi+EnISWf+EBS4JMKvl1vLOD9bbypNY9GcfIA2YmQ179
7WStm42XBKFA1wo/terEdWKInrRYYw8PcCZz6pKGXOXJ3LJRgj3Z2sGi6eyCn5O147pB82uU9WUc
uUa9AnEMhQowDnQKf/0XYPGf2iBHdRec+S40IhpEdgv8dCvTLQjz2XDIwZSxZpS+pPDtybJ4683X
CSO1HB9+i+EOVJuicz6L/8o21ZsCR9SS8GQH3cgHf7jhdgy1Bez3k2KQ95dzWpdy4xonEkK0H58b
y6Th93A8rauVprchTGh/IKw15bYWAOA3rrqORLjrOWweUdnnBKrIyzeFBIUPG+FQJNTFJXzNVqT3
4nDDwauPcTzOrKEQDIpgRLPLpRX+PuLaAT2Ix+RceXY6WqX+TelKPZfRy8bp17UUfCQ5JYKtDQLw
eK55ep7jqoL2kPpv+KG/CYAov1Dc1hwzaI3hTYOnla0HOR76H4KNBYy8T4Px1CXJ/t8GEx4szGLC
7CGhjC+6wkjsSWrS6js6PanJ38Qh/z31t0fm+HQrG9kKh7JyGL01DjG5jjnBzm3U6F8+Ikth8K7o
MY+ApGuKxG/0LAE9QS4jx84STDQa6AXIFLc9Si8iZKGneHLQMZyuCqHRknRuXvbK3Wgn8aatD2MH
STbvdDO5HsANZAltF1/IcykPSS+wIg81KYes4IgFVZjvcUl6t28mH7Evk5NuLKhfX3BUitQOipEg
ztfTDwwBMYQxBBMXDzFNapH6mTRmYlosz2SD0hCUQUF2DA4Z1rlYjaFJsEdwIVYR8ZIZDyJnuAFj
kh/PeZVOI1QYfFj6cKjbHXpi0Ezr9sb9uOIHZ0FxfRo3piOk6zh9kgw+fhSCQkZk1Gv06BPiN/AQ
YXwgd7Zwpsij2otntN6zqskewX59oTNXIHv91J8Qp/xzA//rlnUCoeHj9uXEYv1eLR5skTMJiDWe
4iZeQMB/mTK043G1oaGgfiAElGkoEqzrO6kyXRk1T3hNQ5fc0s1maxsqk9iNhzo9W8TKgVhcZlEQ
qA2T2xJT+TyWxkgQ2lHaZX9w57QoOpCaTxIoijUmsirQdqmUNwVNdru5mBZ6cCLvApqfGKDFSF/m
wSXxfclOpxIjccOSXcdZOIuIR+av2CVNWhiyEvGVos2X7a+9FsHlxNzzjSCINI/LxHN/QWPvegTq
EENcx9UiJIiQvy71NJTUpoAjCxcHalz+81l+MUogKpUDhETZd1C14AEkRY/8nKdbijuqhsCK9MAa
dxxY9jPGcq7c0tC0HA/RuoUqKkJRf+YsuPHaycGqhs1FeTTwlC5VZ5kYBdXyoFyMCYqpt+hVVOfl
+EvcKEru/ImTazz1zNyCQt4zeTCGe6dcgz0QpyRNBrPwGIguhiWuCgbxLztiQVfniDGcQMhGUCwi
EBnHBd3zloOOB/NGjyppE/I/McpF4wNeQSUhzHBJsQH3Dp1iBYpEGzvDIhWwA/q8m92XE4+Q8zMe
fBgztqNOcAOTOTga7Z1N0VgnuPqBVVU64HlXDEhIqaVBe+L+tNu9WPGe8mGd64M+dRsx8+uDBi8C
0gE20LUIExuZBuQVaJKSMLi9El/jWC4+d0va+egi/WSgesga1Mu7VBldQHuaGLPBI3+jODH22X+8
62zJMkMwDI5Kvdk7vetpnnAFqpX8yZgVkfcq3O0Mlhfl1+Q6JYSJj185cXa6lAu9UYUXB1xs9qkV
dYDkbJIVjUGOf4FTWaZi29gACAjy3TYhcXBy3F8J5xNKVo0Riiig1Q+/X+Kx1moJEx8tTkg0FHXB
OHJdt7xFX2ltLG851KY3MP8UgPiEvpseShMvRv+FdpG6MSr16ITsH6YMNsFCTI5Y7TD1WdihwczI
Osy3F8UI1nYiWWYKy0r67DBBTtEvPMBx193cpwf8DMKhkT/9LOhYIxMpO9TBl3mB6rNBAb0DcYCA
XCHw2pFY4k3ASAEJ61rKQ8YS1Rqw3XHUalT/4RKEqyR2bGN5ms8a5J/Mc67Jp43Y5MiKHn1QLfIq
ySGf91MFxQp5J1N+uFPTSvKoX4TZZUF/6IAk81FxSWmuGJkWQzvYOj9ybI7OwoJxHe2vyEadzd8N
bYOVJ8ACp/4yfNSHZbaj/lbh94cGUb2JIKd8Tf8p/txdrKR+vVhc68OTN4FU0Pz3FEMVX74EnJ9M
v7Rsmc+j3KaRFgvhUTvIOxi1NH2wuJ7/Plc8d9ZxkM1HL7PDPaGPAAs2ry6ziuM/r+fL3Ud8fExV
XSeai2HyKrFbcFQw2Q71oLlfvIjxZWO8C6qoZkB9r6+ap4S/6sT/vPiM9jUBloL6xrjc5SfnJw0w
sJnwnVwoxCjlxqzB7DD7nMK9pgTqIr3mDqwJUKZdKSjayEVKnz5vWCaHTfhpc50nYff8cdSFzyQg
g3dvd/c0L28Ydb/QsRF12z5jRhZ0ek4zVA2cDHlwYZ0D8vbi6CFA4NHUr0y1KE92i+dHEIw+KvuC
sq5fYgoIVIC1h1xKQlza5R+S2KRaLTd9WOiP8GkSllmrCOnB5lIWpmrxdGu2sOxk53KXU/TdvPMo
srBUt51OFm+PuSvMI5t+yRyWpb/6M4coVsh/s2KMrr/7IJAE8vm0qDF+MLlLN8BEdUoUgAoPl6lZ
NMIQ44d4oWjyYa99XEknB9hNMVVyudcl9ENjstqtvqUhTlSMjRV3YcDFVmNP/zf65o2OV+v2ZUmo
1BjCKuVzEY4ru3kOvaQtK10CFkexf5+GC9YOJGOH/5q1CJ9h8E/TpMWdUDezkWbwxqgP5dNpFp7N
FBF/W8Hg4Zm6sII/WCTl2I+wPUZih2TrdC7tD+OgQ7J7QChEGGb9PrJawXuygODHZ9PjuC2Maw2D
9YliQuIPr0gXhhsyi8R+I54k64id5MzJXokR5AkWi7aWMoXxXnX+IWYmBDeXi5byZ5McmI04cQfy
ioGcB13kOEXZ0LSxcI/j07b8JABPuOZ2mw5I7+SHKuMAeI5b4ZWIp1T905437rb09yOesYn1PGZ7
2yLyJIgz5XPv1UfF8E4u7ZCBTQzpHBWeQlRxNsdhE9ndQapXIkfKsPHNn9S52zW+aOKlmu8y/uHu
/oQwZ/jteI2w0NwT3be3qZ7KfdQv4G4rK9w3VxUsWp2xp0BUnTrvPr35efJRmccHPpuv7kNrRmAW
PcxJFoewHZk1tb3tHHJ4np9iKewchZy4BfgQgUQEHliKpUfeyLPkd+XMHAxaN2tCA0g953vF4ja5
B22nc8nyc2r9K5Oaq8ElEjLNtSeitVtiPT0RoTAh2sWjBRIr/DBkNGUWhWhpo0z9LDifNY4OxpN1
6gFLijBzOGzYKnpjFMdO9ExJaIWzsZz8L3L0/b8Sp4TSmn5Wa+YJvX1HqYTDwdAV+B03f9QJ56v+
ApzXsLP/lPSnOETck5Mo4M0v3Vxnw1BmMQ5dQ1g7aQ44Y9tv0JEIfy74CXmDbfLShWbyYp9+wFp7
Nyi+cvHtmABjN62hz+qvNL9jVsyEzBQMJsC/JxbcVjNZoKTBpDXyUu5CefkYdV0GiZ2H7kurvcTn
JWgsc+JQBWWGbsKaSHfturyyPNkn200AdNPqOayviQeM5T45eNz+bQV6GsJyfCsTNwkdce1BGNUm
K0ViH0JKI5wwAuLDU2S3Cv7Ya34wqmYCryUXTz3zqMIU0w2Drri22Ml5clYS1KNHbl+LIwiTQboC
/YBemd2lPDHj9vE0DJfN2OjSLNYIY+wlpVQFGl/MasHL7Mzs8jPdUfkCSPZXgvTH26HxHsrpSTqW
r+xLgng+KfOv91tq5XiJArC904MJenaS09JNavXmpgD2A40a9jwK03UaZqFQqtl+3LIQ4WlBdgO+
kNtt/Vlj8JggsI9Z8K4Mv12sqY9hwz2QTfrXaitGoe4p1/LYcfoIq430Txg1d4KbOvOMKg7DAnA/
zFmxC6mXMjSsBcJbnSrjj4JsFmA8wMzLFy1Jeix1UMik5HZKYx03zUbVoqJjvP2wcaAmo0val49U
M3LjHuphzCZp2lm6YjBoJpB7v2nLstzRbC9/ORm7Rsy9PLRB62oInMCUeaaXgzh+VrgZtE3rSQ+C
h4kM41wrfQzlgJ0p2KY2uXH15GId5ah7/QB9odwRoCg5zwdk9bUSmZqljEtl/xtmDFlMiit2cxVq
ciqhYxFdNVnDSx/pIfIv5SQ7lK5Yq6/OGvp8/YnmZ35MeaqnYix+6yA8IbMmW6ervlM/T5QpyTCO
maaz/DhVHa0tK1MWn7Rj5bbLIcnUHDsHLpPEjt88V7geCNYx1gFRgrERcEB+izaimfJsbGCqCYTf
nerT2/kbNKNHcwmWIxz8VfL4dgh212ILwRQ58LqTGgvhm8uSx5HouhIqpGu54wIi8ZkEnjDoRx/l
EO6Xf+lKYM2TrPR++X3T0/h+boU3uCCgzGEMyv1H44aub+h1p6HKFk+e0S6Y4g6dmaEuGfOkk4qY
EKIxiqHIdZ1P/UJWfyToT0kq8a5ZywYdQiTiyU2TvvxWSRtLYDpUP0OrLl6Zquy/zYn+6fmLSdOM
qdL8Hc5jAX693wZlFFqWU8Chx7xY3C+ecEGUZ2c+DTmbxJWhgJDZRwYBrtrjDnd7tWQNgKcblYxq
I/6MksMyGcO0NRVLunJi15Xlc0/5BAsZlB6AhExp+2+WTGvt5TdXR43buJQ/YmOMISPS932e+42X
bBkIcPrgOGyDO12a/u9rIjBTHWiANj54m11PeqRRU6WSRXHMYPzKov8E4IkWoseJSLqOYSiIjpz0
VPF5pCpJWTfi0MdX/hX9jXH2HsHuwLWy4MOm5AyWxDhaxotSO5wgpiohPgKPbVd4V5N16cIur7+x
QJvfO9tPoVrNxcv2bDcyeYdiFR7Lf5ZMckvz7xSGYI7da8bJ2Ohwes7mPy21cZAQwuEZ4VESyapH
FNkBtrrvhCEs6D0dLhP29Qgd63ll7QNBYP8a62uEGDozwwJxxzLMU4qDdzNyqF6SMFqsOhpC8p8g
VADz+m9CDuh7SiNS6nrusAYiPPTotRg1QtzvBK82HAGLVWUSPHFsrgZWlBxKF+ky7fb0VbMrVmGL
XWEWxkOa1Vq6R4pnjTz2KzoI7udrUMznOyhz6TRtSVrNXdl+5Mo/XkigtKamp3GgFZ6M/k6pMTh4
3CCpeTpoe3teSTHjEgYKaPaXGnl9ppjtxOZHzedwT1SQiAcE/0lRmbGfyjxd69zOGmeAjhWIVu0+
0vcJRcz16C2ZTjix4H15ESMuXFlgNr466yNVOFTXru+r+FKgfSF/2ol9ZMYxKh58NTuH7mmfE9sf
FLi59HcymSk9DiMJCAcxDWadz4n/EAsnzHmIy5CqOojWmaDxwChkBEfuf7IydFCoD4LqobnZNQzD
oPhKzQyu23FjoS2nFeLy9+gL5yJeX6L5GJt61upsThZ7VeG3hUl9WZFiWveUmt0Gb5A40oM/gqI+
sspMOnywYSOMjoX3VYlzFUTc8S3vy+DJeFIcR1jVsTvRfHOIW6Tiex58g8Gsol6WKBHykANQ44mg
lumfCb+8tL2g/X2mYn3lB3fixV4GWRu1+kKd7uyVAXKhwQFbHUKDmXw5urxihOXc+q/yYgb0imV+
1kt75UNpjlCGVNaXq8PAmgaQzEqkn0tTymI/XKie+q0gPrFnBiDHuzaqy4QItwHnbwy5vHo5M0s1
QhBWsoG4IDWyoE8PEX9LAzjFGEXmy1TCg9DFoeeJT9cZpMavOnoTE8IrTN7W1UkZawIFOFi3Pvst
mjBu3PyJ8TNxqpWjl+557f91B6mmJc4JtNhLCwK4//nyEbEjbGtiMVkqVkUOo66l57k12at8ACVc
NTCX6HiQb79CD9A6PCMrEoadeKV7Xwsm01PxmTgfLDXpL6wAYEXGyT4Ojl+UoBhOIKysYqy8kDwN
di3JU0ixo+dwfa253wdPYhrkPAeElHUoI03Y1o2swx1YyHWnsGXe44efW20im1NPWpc4GLo8mqBw
tcuLTF0/DwgCtn5PJ5p9Wz3y5s0k0GxgZ/3/KYvtK+ylhA6SO7Cx1pP7Rvedw8Z2ShtBzjIAigwj
oEHtukK2oGUUcmmkwT+y9fx6cckYmrGHdP9RIQ4+lkFysIH6G7nJpH7EOacwGL7AqJQlmoUesrI6
w4B+e2TESTPBIkwhQ0JDfaFMVxCHWwW+XL/aDmbbTI6h9DbZx7xot8o14uMZcyk5uI+uLev3ArEd
Nshkwtdwcf84IrLkx6SpfpUHINV+lf2iQVcQJMMwiBljZprLNXbIwjgQweFS0EiifrWrRUd41D8z
DDfsEgfvH3eoIJU8k5597hXUSXndEcYlg4+YqFVl5IoHIY0rH9+j/HS8NG7gbOXk2pmpafDEJidi
jnaX4reLzu2H8JTaw1pVBch+zxQalVE0cib5wvNq4UZb1hsYUeNeH9KBrMPt6yA9i7Kg+QHIyTBP
7q+OUmxRHyZXHZarMCeYZHKAL6lob50GPN4cQprn2x+jNrI7Q3xGYXYoFbMfsscFK6xiu34NEVhG
VKxVJa1O4YQ/Z7W7Yf590Y4zqtjvlMO3AbEMnqyhnaq2S+FX8vml0Hk2h0XCVyz8Bbaxg6uzPsC8
dxOMzOrxqHECVljC1lWxvg73IjLScCXbbDA75c6F3zh8JCVZxI5Zg/BBIZ9m60vf7dpAYTuK6aVA
9qTwcGEcMsuCho6RznsXL5qujtJ57pTudSK3UFt+4EAHo4j0IoayJ8JiEI2G9x+sRYXsh/gYtsow
JDGP44YOl25cxHNWhkSs2lqEsgiS/HYNBeqKv6uaNRlB9InKYEdJXDltXQSWEhN5YjAOc1JA2wTR
LFFq6nADs1r9GE03rYqD9HdFPOfWyLoXljFhD4unOHmU2VdKw7pv0oXEAcYvLMGLJj1EQBx3Ys+x
pWzP1s5/IAkHxV79oqmMR5kN9H+3WvUb++jvHPhWcGQ5yz8Xdqq9yEr/LB1iImgUBJ4oGkZ1T9hm
dLol/toKgMruX6y/2u2nkPaJPQmWsJSnf6mFn8aCzwKElktcsx9sxecjbfJecm7Shw+CYQm5MKjw
ejdQPkQCdRH3eK4F1gQFx3yBj1eZFIunBYyiEaURDx8bZkmm+XvabyOTWN5XTRfWVMzaVezaCI2Y
pX42aGReO70SM+KpHT+wezMqjkLLvcrsUx+xTSAmAW0Ip+0bd5brKt0iE15UxPA2saMQyUrI/9Yd
hq8Pfuuisj4vnBeL5oYQ9PR/eHbqmwKwxa3uWxsARf6Kq6DlmSw9r+guVO2jSEZSQ17FObt0gaeS
Ki3ncllt937PhH/JgUEJ/fHeXU8k3Bxnk1bXe5jeqUgXFwqJojs9p28MaZi3EVKr5B3Fd+zsjQdc
vh5dClwvWIgINOUHTX4hmOqquwW/oprP07AA9/bwAOc8OEGwU/trV+gq288SBIoKp0xr3IsCCdtC
YkUt1q6NXWtqHNNEkOIkOqMOoiv83Q4Ytud9j9G6Yese8QN/Kk+aM4hRrLFqDhPC/J/qfsil9KaJ
sSnRAp3CJqjR+65zUKcKRQGrnBYxU380Yr/kacqP38kX1pCG+8Kws4DrrxOYCQvf0shMAmHkswKw
8WglcQQ++PZsvk2+cSbyie6Cs1tQLJjxl7RSBcXChGV4uPADLgFW1uojFiNSI04dKZat9+AY6YNN
HbwWZU30UTRaKApDPt+QP050/QeEdLDiWuIjChcI3N4qda/70wtbujAgBctFuQ8DsBfTj+wqd2VM
6HB4o5lORy5kp38a9fEoRLclyQLMiYX0tGxjsUsU7KmvvTdyPUZZJrL4+fGr6bQA10odDwVsRvF8
9jb0VE4gBpg5v/It5AClVR1N8xgqJyMt8sah6BM0wWK4DyfmXS92Euj2FlcbnrGcQ0zN0tn8B9/E
Ek1eGNxQ5lVYQ1fNSjwZnyHOFZMbi2vhXGZLm+F7pnf19c0Y2i+PauiprWoZcz9qpw2LlM2kV1pU
+b9sEB5PMkxpkiMnrlkB5JuuJxaFte8EL7WeHNNOwGus98Ru3PS7IhfEx27UsDDTLJ0rbwAw3F3W
FfT/n8K1eFoE9O0V6xRcF8PMgISlOfY56CiLMiwNDqIcaepHAt7p9jOBCgC0eprUGRQLD03muozM
6T+QqliOQv7QKz/aLC0U2zdzIjzF+Z1C5zYIeZoYvAk/yFrrdQK2LqnektVxW1cXaSH8Y26RAIh9
1e8jDnKYpApBX5RZZt6lfbeJf/0e7HWlE6LWrt2MZWC6DzqpDlNXChJQa49wAvXXFp3Ja/8n73QV
42GteDjmlwpTwh0EPnWQZX9KktjUL0sl1j7bzTJrCr28k0ER6CuFE5p4h3HeSnRmYWrMKY837PW/
2MuupwJMXc0hLIQaCwhnoEqURfx3nmSqsrRHOAVzU3oryLhoY/irle8x1gvx6cAMi8d3qhaQXGIH
JKn/AoveaG/qv4EMCAeDlHctsJv58LwqmwdwYA4GtdCf523rqZCvoYJeutm8c1f3c1sXJ6N0K2lg
EdTboPRAAAbPQr19Cj2zmuuH2LW6NqUPgmB68r8tbLyHpr+h4TT6/PkpKrPEhcasI5fU2qhoBeAt
1UhYK6SxMk/SRdchkNGdCPDjPryLdXiXVT8/2GEr1VbcrVYbfTDvUvluFuJSKK0OApZWf9aEqDiy
ftgt74rhITleu3YACrNPUmFQDtpIHattbJp7exPcJtX7TSco6twgG7vkbbuovSUAOtznzQzrkYmC
2VtcdTqv0gew33ZA+teDdasTjtyfo0g1+FgXO/+ObyMxRQaaa0o0qsTd/CCxIozYrKcp/rX5EthK
p1OLnl5AXXurjn7RH4hvR1z6VC4QqP3GgSSdc4x1rgPF0B+YasVlfe+k+pWb8jjJjF476bGhPTeY
JZ3j64yX6djsVwgdw8IQgwpemPMoXeQNT7rq+q0QeDoTY9rd3Fupu359d9/0uhZ+0ghAEJjtWFQf
PMeplj33ldYhGTCBoCYyRpmajXOVhoVqi/SLW3/FVxZdARiQEB7z2OYlwWltfxvAfJEeGi7lM0yI
AZH7yQ4be/r8c8UbIJu4tnU61V/WVobWe6Rkzow/Oko+3JvVyUhCEi8lJb51CLFutB0kFDL+ac0b
AuwbtFoF6RmS/geAev++7kLp9zGbCGfMsGp2p6Fmj2SFVWSVai6XYZxsyD32iKJhaBHba32b1d/E
STOH9N91EYfhJQjhPPKLFW9vez1fIJov4YEjBq9Q0Ut6Zvrl2EwFxmRZueFkz1CdYb2zV6SJ4n59
GpoBG7qf6UstE7ik6fd5vzExfc18F8q77OOkHgLtLYiPA0GHRYmuNnsHxSUu2a0Uf728aT6fnOva
O3xNE+S1Fsfw4nhAuzitND3cezsQk3ek7SRhVuBXMJH4qhy9nHHn9iARV+Ujlx0XHkvG9x8awNkz
0jFz5Rh5Lc7+NW3yp8nzSVFmvC4cCEXFivb+UJ1HvuIRrTd1ONUhVJj6uFSoRWqapLlFFEJTE8YR
pSPz9guzOksUJC5tHbwcultULRQzAblb51qC7634A9Ipd6lJ3ZMG3/ERixCBNCO0xWOY5CAXPYML
dusGOIBlefzjacmFbtpvbvmIKB2gfYFju/g+ebUBwjoUE7yGdlcbJUJ7LIobxP4mLwgVn5b/jeED
btE01oMvk+GGnF/2TjAPkwkSgcBcx/r2/pco0F6gkxwVkkcCjgNR1oIGOzlCLYkvHoVX/3x9lF+U
csw3/RQ80ZC8f1qA56tK9YZq6tuG2IcpPHFQHaXFq8l4snqCvwyh2X0T5tIqedoDgs49rwC4eU4m
vesnkIKf2zvl0I5ryKOpPhwh0OJwIHprILl2rQd0VauSxOi6OJovt7QgUBher078rjkuu78mRPDQ
ljjotm5cqSc9lUfA18vvY/CXj1P7HAo03Q6fziJZG/dLJyOiRRWA3IFMWI92HO32C1GKvJIEFGQ3
ab7kbUBBkuOBgA10yowqogUu3dPWw5GorAhtLaP9ru2QDEQooqY4fsyxiPVt8F9rhYYBMb/gzDv6
hKrwnyItZY+CRQr7xdZB/+hvdvavvRvjoCYnJ7+7nmcDjmlnfoZwtERs7YKa/8BKzUFbeWbfnlpJ
zCClPAiET9pFMC6b6B25zEX9vxw5P1RCz4lLwJBM2wrSh8huY3sSkC3prEZigXvGKelLK4964AD8
+tPF/jbF4jFcFaV0I/l5p12B2RE6nWwvkmagF8ZNz6wjuY80+uM1iiNnS24VBdFXKR2unOKDRamC
zVirD6kbAuv3k4bt+BWpEkW2GfbsYdrsR3ABrZqFRfKnSBvMRM1W4RP33nZUL3BjoeuTA4jBR+dX
7ilbzdCCfNtsK6zHCNsT+GRKOnD3h8lerHEHoDoVjmLcWKPvvxpbEsUb7mjv2RKjrbyrCG4o9SO0
jfa8LQXDnT0/WmokPzAfXvONhIGoPIzICp2nQZ/VULpksaJ4XgKQz9dI3YsNjqOGZIGpNliCi/R2
0c9mHq+V4fU4mh3jJyuoxNn/3uLoO8hn1RmkJLxbmcLnB5kemzQ6+pEzzI1Pr3zjxvWH1PmfLO2q
HwhYUjJNVLJldQTkppz3/DSuysE5pOBsPP/xOvGmwQldEtOjC80q3FV5WDR+U75vwXTOWvgGsQCH
59EA57zM+/LhWLnWBsm7vqKGS7F/kRJvj/WCWmm5cuV5OnDzwvl6gjWz7ZtNdhbg/kc3eAPgloSu
gBYmcOZFXXD2TWd4fPItfWh9cEGjpTZTM+u5Jgi7wrB6n5JtAFwZ8VVg9ZbuyzN56DxHFByCpXi/
xA6Pg7KZ8HztqlzqJpC9DZ6vkOWCcAx0UpOKwCruJdQHZRpJn6+KQXQttxS91ZF1RtD9DNriQgnz
9qb+hm5tYwDi413uKNQUlLUqlmiDlIVvFu+DxB5QstnvIRwtUfNru4hh+HkH4VOMnjbdKFzgcMjW
4d7yt6N+Zv/k3kZ6IM6I3dwkftZlD3cM5w07BJJ2eqk5qurxADnuoFrrRKK9R3nA0jURe1/3pWQy
KDVO5F2LlnAo0j1cjKxiA6DPOIt3isz8BJWgaZSJau47uOjKOgcinnqWSYdoClI7SiIwQ1EPy+2K
2hbAtUIOrSBRIq9uf++9ihl9Ope9FAYxAVeTFvQ8Noqow9fLN6r5i5SLV2dvFhdBcK3wzo+YX8RB
pyk8/LpDaPmCjMOKHXCecS77rWhm736A1NzHOPzRkrPRTc+0Hp263qvLuOEhd9QSeMSGGqLX/RkI
z5H7GgqA193FBPykzm3z1XGobFzIGsU6wy57XUK3I8GKS3+gcks+ztF2eLX+Lt17XgGYFbghoMUY
7Ff3PNJvf8ibu71ATsBrF0ppKqMdGUd5xCpnBdfLsczJZthn43pLSY5DFdNbhFoTU4HxLfWN6c6e
PZ4curoHF1uurW80ueYeXOZF70oBD59ZWk84Hcduh+MtKmNuv4qyqsiq1yNi0x/rUcosMPk+d5jh
M3Pt8UtqECQ5eSOTB22BKtSmg+29EpJGSbbNSyR+V/ZZVHatxs2qp2PgFGEjhhSE7oaT6xumYhPg
4wwKSa2pe9cpf8Y9PZmDflZ2qG0g9SEi4phd8pV+mz5w7ryBelUKt/fObjhX/to8bduEf3L9kr1Y
7cEJ2HsK+8jMOPRAhFO4sEmbScJHFkG6+Wnc6q4FK5ZFpk8nVAdfiOwgxafvJkLEnTEDe15soG6c
3+Duy/Rme++meVI6V+KWzJFjTfIpbGnRpi6lwngIshYT9dq15BXDWovjIyqP9UcW7ZcpKNwSEkOo
kk4kKk7w8CdtSH63V2i3RzN9hAc4xSMUa83C2sgV3DtZzWQhlttDGRLiHy15y2tG9i+Br5322SB+
C1/8EcdKlu6vYlHHR8n989prCwsyql7upPZrosBYVe7MLnH4Xt8VHmFd9moEJceddErO05xZhCc2
I0vmBIkiWaEIrp6eI2A8JkX4zCOO7I3yb5mtFhGWKB29k0Gg9Q+cePECmvs8REMmcZ6OtHb28n7r
hiHdT0XByzuTdfYFBYdNZsIvFq08/CFCeH9aTxIiap4RO/2tFiSoXoNlYPF39RVzvZl810cKbUKQ
39XZClFMb1yhJgLYcWJKrfo0nGw7EU2bA6O/I+URomk7WeSMEJhDhMjuGw2B3AG8AwOamGtM5ASw
Sf6qsXEiNdPgvnqKljLStSvD6K5q/fJE3QbwcqXjJbuQ7/MC/qBflYK7rc03O6cG7YZpFPb/eRD3
xWNMswA8AH2SP7DAfZUy/VBwfpq1AkayYj6YOKZQtfCUxRO58fqlp66ayvIWOeHtdGtqX+a0FMvI
o7SsA0fGdbCBZPPoDhhcB+arE4seyyFSzEH6DtWwRw53gNv5IVZBExUG9czpIitUoSm/wuVhYiyj
yiV95pjwGdS2ZTBShUaVOeZbMogz5qniRhvb1TsUcgJFjT/IPAgizpUFutPoUyN84ZJb72CLAUG5
VeewI2i3EvTqsgsDweQk9PMV0zCAnIU4xpCyHRx9D4VFKSaZ7DRQ+yRzsw++IT6yzWz5BLWSOT49
279F1SlAxXNUQqcgjvF73Ju0Pg3gLMyh3X916rXoNq5aITSnAH3w04bhgAvEHPK+q2CQPOJ58qeu
LFkIQ1DHVsGrVBsKkJTzIuBO27cmWwtlTzgjduTOwdEgAhXufZmdD2CPnFeAsBtIKKGr6ZoLi0Dp
mv8UwldBW/XWr/s6Y2hbkR4FvUG2BTi+RMQqjLSARRCcmr+HBVe7z6lDTUz0e5vqirRXuiL7a7md
JGODh9EIxuyuCynRK8iSu4OO8KpeoPYMkSFhDQPfIdEx3P2Km/SP1HF9kuR8P3pC4QOBuP+H9c8J
ITAhGItLK0nckRKBacaX2OXE+j528+6NfHX6vdCT47pj6w4X0S3RBtxzHBgnKXdeirvDLfUPR5vL
kUcXYyIwLNjtWJ0slWD9LNyhXGHGhh/a+b8hRyFdQpI1q/jZXb60ADeUxBXbBwi/lInnZCvjlaxk
W76yRqe0askDsC8+AGueNb4RILB/uBx+ifkrhTksDE/G6jpStVavBLnrRctoX4SDEdqpoHq1ful9
Uq6GHN0655dwLfX1AIfJT33u3dOHfJZbRdRtQasX0Iu3vwmJWWmdPBB25P381HSUuQT+ZmLhKX9m
EJx0pHNCNPdhPRsJXDjYh5R9o4n6IdPq8g4uPC+YEWVaK4bKzbAinSgJFgsd8sNNDyQ72efsHd8h
IQbZYHcr/Z+p1ZUIbVDTn5LdRyPlCBebBHtcI2MlX4VtVZpidIqVseUjO15jn10GJuA412Fj6A9V
BKS1Gp7i5BZG/DO+uaaHkB+CGgq3kV2KfI7CLNTlSIu2GOh0vuTaH3PIo5SIpAmK6M5pKcGSds4Z
UZV0BnchMiHQzGbYdBWV4Zus7xQnY+1mTwDjdx5SSgpPVHPIEdCZ4adOFLjn/XUPx+0voIyPIzWG
ipSGi0EPvKIBYE+Jsu9dn0Bst0ASep+JYeEl1rO43jsOzLe/ZBdh/rXQFeS28hn2NBOnxCHi9llb
03weF2kd87JVvc+plJcNCAXdIBi1BfWjz/Gz+VHQTI0LO4GwfN+HcX5CvsiVkO4imhWFqjh0Q3ay
c9+39KzpGWV58YD0LcLKqnP8OYizbNAXdce1odyYO0Wi2sWuR3ZKkCpgYQGGReWvcKj/3u54MuPp
M3HbiPdniH1rJYnthgk+MgK9VcCQHU6UBv6Ie7F/m2Ps43HLyul+LJW96MOxtpR6I9DuGAgf+rEp
WjiMCpDDTeReaAV8YXN3Zm8t8N8Yw5Gc0g5ktAcQ1aKFPyZ+69GT86ZzuZKG9njGlmxOp28Neq2R
BcTsM2puU2NzXR22jDgu31C2J5TOBJ5xO70OJ933MWoqbXOoq9AOuF7PnAmOca60bXmFkDjgpw3g
Fp0ZNs2IedHiyz8xw1gu71zW7TqpW5cE2s6oE+04Da8JEOAkpzDfKKw4ecoHteHl4bK9rB2Gdr+e
1Fmw/NCC/Y2bwrxFNNyMF//YK0U+PYnR6tHXQwoaqy9SmVNGGf+14couT+DRzjEWEjVJXNPzreYk
qkozGQTvHe+l2GR4Km6BV514wQoxrU3uE8apaVxH66dn77kXHw2m+Th4W8jsMqA5jka4AFJwoFFO
r84L6p0iMFuHI6MsJ/PGk3S8chLkGb4IJDKXdrfCwdZcyxS/PVhrDYvwSJzp3PEVFRacRMzRVeP4
32t6WldFNbpFTqz33SXkNAayG6MbkWGC2EtaopVrs+q0v5kxAxy4uPM/wH67fWjiSWLP7r4ZbWrR
Zc/mcVonFTy0/ibXU1PoH5s9C3plYS5kr/oakpEZTMrPKqom72SqWa801tNJdXASGTNneJnEKZUz
SGz79XG7mAcmPAhFCMvHENSgZy4y1+laKeeh7Xo3nfi/thmu/8HvLM1r9ZYp5QmUnY6tuYAmgyQ4
oI3v2vvCp2YZNN0rdn+lsLmz3GN+5f4GFWtSoHmM4YRna4giTMxcg/omBcYmTbxJcqyttEf0ofBR
O21IoWNy91mGlI9YHwGX4Sp+FOnn6kRRAjSRs0K/85xnpPZ2WnjmKRU6XGQnNp+1VBWYNfY1u/Ap
3Wq7o9HE+goiRyFxgqCmdnRLJ13Y11Fd+1M2B4SxPpwNc2i71Cd7Zjl84wuVli398U6gSGcIlYlT
0lSC6g0pnNUVq0JWKFgxpCyAxvqegUfJkfDJ56s2BCqfXFQ0MA9fTSdQ9Koq1TdkQY1yzBk4VH0+
VFp79hrAsN+LQNXyMBRUKs0zk/SG2b6ZhqUZpccDJVV/OyG5zJfJac3H6yzWKypuDt/rEGBtuvqc
FGxoGkMSSMNldm+F9thjVH9Lyskodg/bsMZF5di8Ec5y06xx9Mr1Eccrx8MpnhpB6jDFe3+PUqoB
7pWYYY23o/16bf/oE4YXnu7SpT9UDrRYYoP7uYfc2B0MwhPlRp17b80tx0i3j4jMLZxsQKJ6rZAO
rBvJTvoZuXXDjwO5fkZ/Af5pmhBgZGmrIdH1kR9T5RddWYSdeSfza0tSiOXDaVk1TeS5t9023Wn8
Im5Dq6aw/PhzOD6Ek7O3q42rTYsbI4MY8pOMYiQssMTw7DRTOD2UMmc4FJfFq/bxy7DL8zCHX75k
mZohTkG5rm0NpQyB0Hav5vD/Ake8AMoDxny9KQCeMxRsSdiiuF6aqNvA/PP3hbTia5yKM177q+jh
Hguq7rD1sHBfhrV1LZGU2GFUqBV1P4+C8ZdTn5S6As85y4//3aLqqaRaYmMcOqf5glCf74rTIVZb
l98OPLXHYRm6s8XmlJETF1J1iwHs5jM4+kMH28v1dFXznyFH1OucLtrqEvVZEoGkHRGH0WDFy73o
rPc4c4cvJnxlcoLeXJIDUtgr81te93LYwHCohBuf9nBodSCIJ1VyNb2Gs20jlukZrXBgSzWKnaGj
kBzbH/7q1KBlY2nreDxCnnQK6misjDZH/RSvdKcDAqL87Pt1ZCZC+N4ngLRqyHxUc06LtNlOGriD
w14P5qNwJ1Parfz57W2V8VOkkXBRzxxmM8N/Us3h91WPsHStaCBtwIQGXSyYpcL/aw1hza5P34/s
4uWWkgOoHYc5HHmUPcson9vRGkyM94kGCHWQxJ0XwRl0WrKRemSpomcw8G4VcT0oYvZ+mItorCo/
rvFVmuXIKLBG++Pi1/CO8u1XhHigUbrp8aVFf7wrrxT15cbBsQ4S1oLjsgvwiWoBr30yXMv4m32X
0bTm2maYz9CkeafVSGlNdL8gs1h2qSOILmNvB8sAgQyHLC17Lb8y8eMnQLRbxmhlCSAS1V7dGZGq
u5lsCmTIkOERfHltZthnSNqvqb0Kxmu+Hgsfqhh/H4vwnE0ESLsRbaymUk7mp0u4SlUbvzXJ5svl
y0QK1n7qObtyOnjZKhfEr3kVuyY+R9wClF6wcsCVZOCas7iN3M4ol37EY+njn4zjBWitYnZgwn8s
1vysS1czCVtQ2eqIthi3whBJ1yNEwxupaln2yHRjp29kinn3POcX8/KvhreniU01RQNCivAGEVT2
F+KVXn1QnWGRi3Fdfxq5vP2/w0TJ/Mg7xZf6kxdSJxoooQyMy4GR25VhqlnkGO8b4GVgSf8kuvY6
gQgZiG5iWYFR4d8pfikKQ4eN/y57QfzGl58oLRKZ4kY6ve60BoUDA2P4pBk3MoM0pl7ppwtEGzD7
QGGL4nPZiPlBe0FVL/rxkB2/ww4K87yoZ0jzz9GEg9J6jHcbH3muASz+LRtJMLRKPOaLJh7Z5u5y
cDJORiEhoz8QOjtw4WFgY/cXd6te/H/wsUUpg4xqnSieJexa2gjrrEx2LG9UImrDdqsjrd5t40Bz
i7l3546PM8cA3vsZb5ihHgKyuJxii7AOo7VkQxN3tKhcDihWErNWsz0IK6gd15H6bbGAOYg+12Gm
L39jk4iwbfobLvziXIa2kG9ZNIzO616BGnOFz5EDnp2Q1eG6rmSxIokUsm8mmho5F49DFSi5in+W
gzHN8vP114CxA5FQyXIbd+tccuM5ptuU588bLse3a8yutFrrxLjV3CvXBJo25TegFu5dXo+WHygU
4HvlHuXptZPJ2tmP9awt+rewoVsRqCwCD9Bvn00p7qOTd4avPUAoexVJPNMdKNlsUi7b0K9BdkMK
8cQ8HZOnzuN5WwNS9hOE25Z7t4xA1hw4rY3+QkTsjKH+BaD7xJ3C9yeFDU31MDuQbsnuzI9DQEkY
F1WrUJFYfnjsac2+9L4PggN3zFG4bopUF889T9OGBhDflZwvlbkfV/bUMqtS+bSXjA+q+1nF9r0S
uq5wY1KRS5joDWvEB9pO1UVkthGEcNyxfJW0FRufc2yml84svkrsnC1Mw+iJ3gztcJWh4yxgQDga
oTkVUhhE6Hl3PZPnSItGlQzkxAUX+j2NfRUKMEbDj2CKev59o3ylBU8Z6TRKOjnsAi7FP6vbWm+V
4Z5VHhdQCoh0i+9TE//Vf/NsEkMqtTKETTetKLW16cMKvizx5TfMLXPsWDp/+kASQhAssrqHrWaY
jMRonP9967VTg4Qd2Bme6EfTXASKxgRpfttr28umvxOLgurvktTS/0JxLxMPKn/qc/mYbt8syhch
ei62X8fQNidUZtZnLF4XZh5P+iSkMUqf6+MEXp51bHvqvxK/dF19yYBvYhywbkgfUPPkjiHAxl08
tL6A8JkbpqFlNoNmD1sJmUwKw8urgeclVfCbCsCVJ/oQayBUMosi1OxO7D+qkiR5fKP62J+u+Uir
xkyUDpAzdQEhTHV06M8zUodWPo6E2yQgCDlVE4IB78j5ZxVNzi4Cdjf9MxTSE/xf96c/28pRkhFy
sXjd6CcIPo82FbuV+nFwJ+y/PLYfSBFZDoDunecIiz3vp4FqKwob1ULO9AIJCXx9DTvuxdvPMaNG
jc+T+V+0TOlXON4jkmlbKRLHfm8oktmmflR9Mu0Udb9pDbUTgWqCMj+1xkvLEg9Kqc/xJtSg7SOE
749dhBn6r4WCe9oth0gk/MnsBgK+x81epxAB6USKIaLuBUQ2a0rmKw+yQG69F5FMx5/rLWrG7Su7
e7oIghD1/rO4mWkv1Bnkk+Ojk003ta+om0GPq3Z6jlZm/8YA5O/5H0atFhN57edho+kGPgMN9rn8
IOFBeUj8Kwxzx70ePOqDLUU9eX29a01sCTPmCKqYisBOwdGZoFVToPkXIVqs/vSLuqygqPOJmq7X
thH5JiW3j3GWnZn9Wc+Kli7mjBBIMF8GC2dR85zGw99Sx6mLd41IvXdg5oBJZuQYGtGjP8Ie5Mz1
LJ3FzKR+pZZxakoVlNeh/3bVXEFmAK2mKbmoB1mLC299VsU8CvQDwYvaBZiGfsHAbnMuNPqc7O0Y
N932ZPg/FeHzeHjnnh8czApvNMJr0Rs5VR4ApangkPIXiCyCmpekeAyMzQf5UzY1fn5lcCvmFK++
ttOLT/cxBF79A+YMap6DouhrXVDuneCLye+umr6ZBidxW4mvsH5m5p/4Mrl7VOowaqHV1QQnv/c7
KTn92dK28rEKe+U4Ukw1aoBr0veRcFxUMK36AirPjAA4cGGtVLXQE4I8I9pa5Jit1BUuRl3rWes0
La8BhGYzPO3/FDcHFJhzFBv04i6464dllOPFF5HJdR7+BVVqZCDIK2NfpGn2g75Ps/MNMC+9KmtU
pPlwkZvkz6aell2xIhWBv0dzh/dzYx7x5OgKByc178ZhSmRu96ogbaJLLOydztLpHrGm9qUetqu8
0Ee6IQg+t8g6rOk+7hlDiH3j6Xn0keyBmwPaleYbuUjnqsX4aC3o3EfK1JQnbK1M9BPbNskOntyo
LQyn8asPpqXYlWPI9lWz+cug2TXcoGQ4WuLF3UsKbVlUdw4FH0W0AkTDbnFc7RpKuFMAKiTilXRV
TAkDI7dJgP++5NA3ECT96RBWbbPzqxrW2yb75CsnFrCShc8FCLKtD7MHzGe6wPLWwmzLYLLDe1U2
BDsjIspdp02ZQgM53FV7lecnvM483NXL4amglKTGzkVHEiI3yjZGLZ81iE5rLbc3Yo7DbQL97ui4
8gkqruKTqTRcONzQaaUMXygLnyuwucXrCcSObdvDAqm0a1fVWwkYmfHv52Ro267sJfX2foYS1MD5
y6XUugyCZ14KyIWcro39cQ17KurAGgbX5Tfhj2TUM/ag4Mp4KCxNH8ukNduUmlZtoY7pzx2hkiTR
I9f6g6JVF8YeTul2TdBQqup7OiS71CBg87RCigd4IVDLh5W8cAJr+xJsICoInpEfaazF+WDFxMVv
EXr3IRo8Qctwp9EWOqx5KiR098xSY8Pin9w4gG/OCLlUoNlhoUrxn4BWC9tr/9xzokdzyUObbXe/
+5Ad3LWEiklJNsLJleJp8GO4f3/uuq+aG5S/kJY2FzxRVo6nLGy7NkDmb2lnqvJF4dCB08ageSWz
5PUQmMAxv0vLo5OWOaM9JK8AZWYMN4amDYlfCWLLY43AxLsdjUqZViYhrV68N3eB2g4nnnZ2hlTO
mYZOWzaiFhTof73dghKE5Y34/IOuw5re/FG5VcCrlxNT3Ob+DONQK6/garUWTrLjrvoV4J5Jw5BE
FZhPFgfZbQXLPfc0PIdQRBAM1GMfcCusE4qKbFk/Pg8WLkKdexghNOlf+i/LrzHeIer6VxGEEStJ
ittN0WjA0bwAQGm7ds15u3YNp9KuAzGXqqVpHhXEUyDrdsysuEtwcdqIrHkqVHAF5Ra6Xw0j3s3K
dWlaLAKCKUgvlUZZJSuitPe2sbr4ITa/911R3USJkeLqAmihgl86XVpoYMHQEU5n648sv/Ce+GKG
+cWznYVdPncUyG5P2Ob505fTvIIDZAXv7cVNocOT2I00Ma5GVTdKbasBSs7gmP8AxHTDphDgx10X
w+CnjC/ZzxwD6cXPoaNm9x9s9klyV8JGVkuzujrB326K0nRx0yCl6sZVUlcPcgmxVflXIA3XhcZ7
Kxby+WsUNSF71RQrjUrzEXjYMIxvRHtpsGKnDc/onhA3LX8N56FXkAK8TuBjSPibu9M0Cp2yjGhv
bHXysPbyXWMI2DIUDzTvn57Pnak09m9i15AXWO7h2x+I/h4+67DjHn7vyd5EtrmR1+0eGHUN3rU8
Vfy9EmnU5XB996Ag12smkywdhioKQzrJazgtPr9icChzYt2msjG9CeUi9BmswXrKsDssgmd4DIs/
6gjg+KOtCP00k7fAekdFsWmH1BOkMcvfq+M8xodOWjXptKF7P/93Gzx8plUJ8VqiiX4SjYnCnGjT
7fbB8yhFQ8G6OaYtmvp5F74JCk3Zgy25ePY+vq5aLfvE4Ih/KmPa+bFSKInX5fKgv7gY4lTbHM/o
+6f/jINQmWQKPMvRyNV228rbJmg4KrymKqqWzVNhZd95twzOO5TLlJFMsVpUgbbyB5i+mdh2wcWH
PaicfOtJwzcM5YBW4aeB0oCD+fg51VY7C8kU1GEGABfvqpxihIKaCOFeB1BFbFEexRlxW/H/vU6q
DWWxlNyIWAOWRf67PI6zBaEJDRHIwzzoGSHYMmEhG1dQsl749y1mwQbN7TV1a6ddeakYZAj4JLgp
0IVgiEWynINFFcuB4Ff55g3JQH7//dutwi08rKX2fSM7WqsaeZHNFh+AFKcXmpiF8tgOAUg5U3ZO
xSB3WzOqBQEFFlN9je2WzbAhYou3lYswz91xh1/Mub1rhV5YXBolUGDuzXUWS5uPwq90We62G5ED
r/ciq71MVdn/2pYJ/imWVpZ2QPy+My0cUkOyYO9ILPdV6V+kJIc/iMkYU8cxnAmXwqkrDkDd0+T0
sXI4VjBm4pzZKmBWRA+JscRr4QtrrIFlO1SFR/i9+zaoTjhWSdhFLOjNy1cy5z6j6ODTucrgoOiY
UHuzZ9oRpF5MNWL840x+E/wkH5mmCE4JhM3AkdzHir+tkmkZccfwjbFHWkIejp1PXqk8qPNPVHBr
1Xq6Q3wBkf1sj5JiJd05yP2vAcys3NbvUE2+Eg8fZxQL+kI+QEDutTLQZvMBdudzhgW+Rd8KhZJh
5usMtW9MAZ2MbGS8P2CPplVdMSW+TKDAuqrmA6qIVnr2XHQYvy1y5UuHxn8jLOTDtQX5M5GovM4P
sEKIzPDilaAxe3OUsHG+GCY6pds712152ZY7RjNBq+cMW1zO06bXMYmmW7TSO8UeveFBA97G2gIn
oRTUOE5UaU5K4qHFz05GZvTbHHw40PIaU4YAqhV/c0tHeOXmxLYH6+oJ9tmRVkA8PaXiMwE6VMyl
Ls3j0hTIdK9eekOESDYkzHCPQAYcnXnGxUucdQo9guRVs6YZtfeP4f+0L+zdFlDPzqNAWUhQtvH0
ZNzjBPZVaiLUjgVoJCbVaAXQzq+ycNRaCPVXvs6vcFHOxzuhPtEg2qc2ybWLXLyWMHpv5Hdtfcpn
7eB9wx7w4kxiBWuDbaqdOK3bWPHNSI2Oyc1JH7oP2zLh4jMloWVqBW6EzUYi1Kdrksq6p+FW7LGz
zo8XRlRBq8VpCy9QaGmvyAvwhzirRpDYdpnHxAWYFWitKho4ia/0SGumi034kxmSHgUm+cWLOI7G
WrpUkh+e2ucBHmSV1BAPXfBUTpWeRw5z74777gvUOCelj2DIN0OKxn68pBb7cdqkIix+DPDt/4On
KAsjr1jPv7f3EIXuKsffL/0N2ixTNVQgEYz5VOBGTPx88GIsF/XmBqgPpjycwCuk0/E8JuCS60qS
idUUyNn4WAGx7MjNSBglSRhvPDr5CH7WO6wN1HRiiPXbLsgiR6rnSNMFq2+1Unl0xBpKWPXyDuX6
V70AQ8yoBLC1vOjeqDbglzkPqusxDuwT06EE3iAQqK8yFytFCun7dfIL7e/4xroiPT33z/I8OJmr
KimwF7ODzxA5bSLL6udVo9SinqtTWCaHDOkjqs5vzXg6BtcrHAiQP1W1XkUpuiaFPWygsPaujMO8
iEw/v7dW4GoS7GNO/ZEruC06hgjcq3UOXoh4zKq8mASQbhEkCESlenMW2c+M+zr0J3kcpINeUj3w
4PnRu8y55vR8uorQ1g3MMEBE8eZKoSP/rv6mY4Rqd6zyJ5XAnFBEO/QxMTWBv4lpH029Cx9Hnww7
5+aVFk4RRPaGublmr5vJt61hdC/Ix0CIX/UvPlutV87xOY/4fXFq7KWqtd0q8jKA6tU06QJRtm4n
0Bltidw4p4Ewwel5SCStd+st1QGLWs6x6Tsnjf+w9lMY8WbyybDj/RnNYjHjMWsNef8sdN8jKCqc
k0bPeIuoiqndiRPNKetyYTwyf84UmMFAc0beq73vO3EcKXnhunp2dGzwtMlJqTcsyYRrobT9Ygm3
Z94VUxZ9BiKDyirtPE6+iYErf7uBql/MDOMXNSOXA1KynOCO3a9M2Tn8FTSzJMypwRN37VugPmnm
J1gL/W/3B6h5tf6GB1C3a6f4FjD5Bou6+tf7bR+buseumZNbEM5yqAtip3m091qrxmhm7U9t8gpE
8zqeARAJuKTnFOtBE0VFYXZbyI86/hj0TRt3Y1C5/rhWW0gkXdOqVRYco3sF9YKQPZa+B9tV6W86
Xzf89qjv8Rw605NaaVl9DbXQ1WUoYyn0aoMiTQ82bJtyUD/eFkFxUxYyr/FAW59kbsbPsU2JQyAB
+uzP0g1gCmYGoaBu+q/SluA855JxgupjZUUmIJPNq/IfSYFcceayKAKO4dmOfR6cPisrGqP9FAAE
3XXw4Mvk4B0qXk2LJaKVxn2pR0bS7518wieBX5xUzvEYO6eKWi220N0BRl+DDib6ExRB52SVhx5r
MQNMcvUCyUSJti4Z0KelLjJqnVZmaPfgRgr+ZbAEqT6ewcuE/i763B1tSsQ9/00weFtWA79vTKnd
BXMIQlIEGtq1GQklfQvaGRSNEEwGvg7UXxf6NOHQuPn7RL0c1P0dmjyzN6gOrOlZ+nykOYu0w3v1
VGkmSl3+3bldm7DL2w+Jrevv9Vvgls/qg6km05wiH7VvkyowKbUAj6yzVPHpJwtcDfvJhlgeKYHr
QCUVtsl3TjddJ5IIN+B4NPQ9XbltOuJXjFZkX1T/IY9uvG+Vq9k+cpDf07Zwtpjb87RzStN2x7Jg
dG38aWUlaz9XXtU3ejy3EtkHXDDimLEIsYZyeBP3ZDTB+rr/Zw+04IgC0SlEmTBq4BpcnwVt1YWZ
Cb278hhbLy49dDRw82g+wpqaFZiJ764wdYS1NU3/MHuOnII1zzcA3khbFvTZo3WGpNLMF9u7+b99
2pdSsN8UN1YQfGBXd0nW1L8B2B6pY0LnhYzhT0wHwD8hl1OjtRfNFNi59c9MOe8R5uP3KB7WGN2e
11Yh7M7rN+7Is+c6XFXUrtwM+0SpNFgNQVmcz60ce//DnkuobMS7EURnybhPXyCpsfW64qYzpJhp
TU8RRagwQJBfDuRH+Z6pzABLIgD5u2ck1il0Gs3gaXzv4fKUdB7u5V0WepJMp7uFaDYyHV9euFJs
jqrqeEnv8vev9r9JkeQ2TSYcKAimztfezvI+ithTznedv8v/DaISJoUjaJPDEYOM0TRZ95iORqH6
Xkv5Zd10mktkueXYs+tvgcCWOe7TB2M58WEN+/lf2Kpcd4lHkgjK+bdYGU4/Ncm96cG6pYYCP2pB
Epc/ohsjApSsIo8XnEk0Bj+BvEFi/BJ8ISEHHWNzXL+mK7oxvWPsf8YqMEBKTjN1xCPYA+ghafGL
sGgJ9rW+JjqSgeio5PyJAnd8CiAySuIHTmYf1EOGzo0zjtn1hBE2NHPp+QOdtG+mkJ+3QD14a9sY
Wc1S8uAprrdyRJ+N6JaGy9TBCVvAuEuT0/1xsODghE6bOlDWGt9DU5ifHshHgxwQk29QWlrXj3ej
1ReMPR4rxJqH7YG+SoCkEB9eW4n5IWQcaGOR7EuzxedCxwRtEYY1xvU2x35YT02GO0T1op7bzeOC
uFREuQWxnxzFXvjbzQSHnUF+4ritxbJa61UOXrIarm6koRiLJb83hegcyPgYlC0TvRn65cnb1SRx
4Yq0XO+NFIive1W2XKz4+nX7ekjpQ/Z967uJvotOCkITdLCQ5WflyvUreE9bZv+Agp0TQg+xodDu
yFZKHX6BGHc+CvuoxOGy3985WYxev0NC9zNvpDs0IKhSmvCNv2ig4lQJb4T1nl3xf9JgbxtS+J+U
KBT4O6IEwjEMbq0UxwwfPuLh3iKzDLtriyb1Z7fgM0v79xOkfcjf7FZcK+HPeqGH5JNvyhwQ0OUm
P/niWfAhmBEvBVCBM8lJOM95rX4C7g4yoXThvt26BCYeBO1gsmgmZzTHKKmvbreiyiaa6mGz8Vp9
/vzhUClsC3bjRiqkuVgWjnntpEsu1sVxTMZKxWwVofXdOlfqaYQiS/YJfiTzqYomtaAntlI6pHwd
7MjqqpG5yuQJu+HHHeZoBsbKSstgMO3N2eobTSCWLIlnMg/DoVYB5uqMXA3yaRQJmLnAUCyYesjP
LvWcuBWb2m8Gael+OhNILhWLuM9N/mW99IdtZVBPGLRJgOPvHYtjtfiIuhTOpNfUgauSsdUVsSfB
K0QGUBzwUcIRdLPxcvFbA3Fmjdkvd1mTFTQXoYfXxG+nfmNoWy/S1b3nr8djRmxGbellmPo7JVBw
qxvxZGqn5PH4X/qIvlAq/3EHIYNukl1XkxScVbE2HI6PEqgy4AoUmscrWZTrdn7qzguViGPF9tL0
5emQfjDjLI6WpgmOReW9zcRPOHCoUwBNSgS2+NyAYFBidWrQFraoWOKXc9vFEMNY36dgOyMm5Q0Z
sr14Hp9nYbw/nXYZcCQPcorSdPWl08Zk8HoKaAmDBlMjcI2fc/wr9NhrbF9ccQ0CcnFNa2mAZMwg
/Uvy61MfLSCijCjwecnqOHO2Pk+Trt3LomzcTXkMO4Hq/p2U/DxoOfxtQvlMd3XJClyyUZCqCzjM
3gHHeISvdqOaV6kCxQF7BqbJIpTKbzqoDde5oCGhoxaFdtjx7WmRY3NH3YOa93LoXj2wZ9oouPLC
aycnXp2ZIbQJQbvX7gR3RbWbEzra4RiBtDG4iNnVzFEILpMQmopoP86BXZSob9Un0tg5J2KTvsK/
KvOm2Ag2q9srQN5wM8iyUqOGsCfJR15AMuu+G+U9KCAduuNu5rwG+dgQD7jE+Nc4JmTmDS3DKp5m
ai8FQ1P00fo+grgyuQI0fp85sFoGinyG3N+H0lUXjVeXnkRBKzmdFZQLGIxqxJBZivDkeA9mDNH+
3zDcZ40WbVkqjxcBPuw2NC6NAHoE/yUqlYOcZsDNmh7pzRZzVk6DO+aY5OIN/twE0FdPFYRJxIVb
UMD7Uy9ieayfoQQfcpW4nwR0FVuWJNKAffQs3wJeB0UD9LioTo6LyYigFwbjzKNvvEUxfciMevN7
eI4W8/Ztu5oOFfkHzEySms8rOGuT8lUvF51s2SinL2040KPPcXeI6fatBUf2w7LoPbQ9Ne5pbpkF
3uyfAlbl9wu1kmvzfTlBkt6CMDU9kJL9/z8Ch7JTo7QX98HEPXWLnPI7qT1wLPP4ywieYmuG68sl
MOGADgMSITDgc8VSCs6JSDWODusbeFrLcnlZxR19v1vjtJMqdxrcVhAd9ipp1U8gfOsFDP02/ulD
qSrGXonX5uhT1deyIGpLiwhKgJYnl2Anb363eiLU//edVpJEDZTwxbaE0TMo6vyQtrRVSX5ENa03
N7zLo9eq7A7oYHYqpeVVMdRK6BA6HY0p9hY6Nu4bt2cc8U3/+Gl8z30WgKpdq6JZCNtkHmZ6qjji
zFWsZe1BWnUxTw/p62SpuE3IEFJHv2J7rHqX86upiJx3W88XCSVIXfXH9yYmtPav9qdpBa1VfpgC
zAisqZzXeMcgD+YxinBXLUaI8aRFOVEtt8PeIlDql05T8ZLO/I27XytSohCRIFbnIrpJ/Ialjt/w
EyN0UehPJzxaVaLCxqERK989NlXHgJf1+764Ig85OYgZG8h/R7br+zEXnVSgnWeOcUTetEAcSpID
sikjcz6M4NzIdFIP8YwDAJ21l6/3oBWTx4s6J7oDABIG14Q/FCoQNb0l+OckT0ywsNZCNproZ9mK
R56w0tTZOpGhC8h2nddrL+cAnxVXjUYzTsEFG9v2aK9HDdsuN+A7FXvGi7J3nQ9SFd3PVsC9tHm9
wQP2dhQePGKQ4Cu6PwCMOgwscvKfae4zKInELXz5/mo30rWf0W/twHLVcmUpPG+c+ZgWWZdLEkst
7zUAgVCJcrxCUNhXADnehn84FMFefw9HA4UBxWeGKIRhnkpf4yH/idz7QktftLvQ6ZH31eHL8xfC
H6svI9W3MUQ0Z3hBpWogkL3Rn4s3wkDOyIB49DmTIqRj1vX/BrGarYUgEAi7IaOEu0rREsJQ2vIs
7+qoZHBdmlGHp+TUtNH4eV0TJ4K8HhXSzDOsjACOSwhTHRrSElals0xUbAuNHn1XGhNv/0IBT4/g
DIKFHC5DXsqaRks2kBw80GjvsJxIoKP8/eqwxfKsREBFOywAGfmYTC1g5oYX676dYcK9Z1XM5UyX
cJ6zFEYWIKd/cRT2LihUpu6uwox3b5opJapE7VYeejeSAPgiT0/HlqTFqc/22BpKVsffGxtoipkn
0w61QlJAlaHGt2BmgzRdflz2Tr+2U2Bhp4tjKEKGLif1HQuDUeX+3gV720ZqwiDRxNYXM7suD8+c
CLaLISKmTRk1AtDwfcIhBACKLWB9LhTvJOf8wsHw5PrguF28xPIedNJ6v2NlITddbUOz6meNIeau
3tHOqmz4G0ldQ89b0sHowMWPPnEJJwlMRfBUO6GXv2txlJ/knLCmsJsHfsKSkg/13OMeO84i4icz
/xzHWYFm0HqFwaHshOJmzVcjT4WNUzMtBiR+cROlfFkqfeJYEUb/hArfE/7blSqFuZDBkgmrHHw5
KmGbHkPfu19g+lXmzmqAi+WwDAebgan66qJYjbML9g4JDk5zw5+VSGGLgX2pp0oXY+9ej4GeXG+7
ptg5TGhxttp/gENabAY+/2zctzXVxLgAQD0UEyaTY0BtmFQ434EMij6X8POeX3X7hoHTwOv+21EL
TSKaUJNsmSmCQJc22++M/4TTh2k9cvlAHBfSfHi98jHwmMrxgMsbvBrh+MwwUfQXLqoJGcY5+2Up
kWRl3kMNTRKec48wPWDh14GoBmnudFhdBnV21TnO0KC/8ftDfD0gJ6XDJTrd3S8WrmbTjVOZwnDW
mgUiQFi65AAARim0kqDK9n8o+VW1BKmd801aHJG6oaZp/cbLyVZSKx1I5pc4u3uBvO8N+j8cUdhx
Wkj68Q76p/QI2V6WBCFbb8dqdQnmx4v4JzRmFXDDfnW9YPIv4YrEDCsA/lBtZ0t05C6EbE0h8n84
PZhXl3+DxqtM1MGodqn3LGQ6IS0/NbDo5NVqOAXyeXC6ASGpawsYCa3uaInitheR0Qdh5Trm33RC
yzqUnS0Gpvhs3kZLmoalfKV/K7zXAykAarA6D5V1TcX0/MAniH7BgHW/RPt2o7O7o6ptFarYN+Ez
EoLCRWcRRlRFezEa3CSatxy5PGH3dfQVx3Q6bPbVEg0QZt8irbht0mfjLIyheT0mynLGuTrcpn+J
YcvxLisYcP7mFLpNmlQWj1G75VGw47+CxuQdsVe+K3HabWSKtVgtIWzcIC8eNWhG+lf+Aw7nkx1F
r8as+JAZ382Xw68gEfizjx6HLO4fukiuFkobEzr/Dc08NjgbtR8yo2LYHc/lI/oZ/vt65a5GI2xF
3YmZKKOF31ANHe14MX3+A9n9Vr1lhPPzNYDXXfjyZHHmyGAefPqURe3nUGXj3Bqdg/i8kqLDwI5+
/WsAsedrCdHhO2BSYV2wGg9Y2tmYqf00cDKR1bdQrb7QzXBS2zYRi5j3bYdhwDokiyr//K3KfH2f
paVKO9qOd3P2HBZcNY1WUjiZMTfk2joLOojfNMbXnLxmpc2OedtDbAsFjfNKxZyBJJLDE3QgOE4F
HZ8DOdMygbl3fk46eJxPDqZsqapwAFrWr4jwIwLVYWlEvaNPJrnSAMlkxwLBOTvKGV6P9dQ64WdI
xXAN/IUYqv5TzHiSuh5Apz9A+mKUDtcgjhrAVI6RV0AR5mMI0oAZOC/bazUl81dRmW2P/FPMhU8y
QPbwGVtCTlu23S3Q5i+Hh9k5jJ7SpIZhS5B5zfSGyF3Bpu/UL0+BGmCbIoirWeddAO3oA/GIjaK4
5URc6piRJR2P2KaOaEiWylai9GvbndDmuVvCtU8vOCHDxHf4sPL/bJZorH/NaqkpRUVSqulV6FJt
g/ggOCtDyivACE8Dv+wWuwrNbEkRmDkIm52wtHhqZLP7FGH7dUePla8tJG+/AW/w6qwpgDMBFT3g
uVMbExaBIGbPzKB5VGcIMRUALePYiF9ejbQQuOPn0sBfLbjxze5aECR9QwYlV+Ra2sm04evLo3wO
mgFFRaFlwJRL0elLtjKcZVNo6qujuhPnSQYDu/Ht0yDPg4w1ucoI+v1MEQSHaSHhWiLd9wlrLSFj
0xODJoAHNI0zfhoGhsUbEgQif92SQf+UeWPb+kWnJlUiJeSczcsN4DRCnOT3lQTNPipv4q/eYgon
kRUcF9X/NCk7jXhsZ+lyzR8IoAwpZDHaljdbZ6ngIaY/+tvTl1mtM7C+v7JYXVnsc6BW7GKVmLD1
c1EJhEm/saX0MIB+sViaOp+wNoSH/OVNIReyUepM0BfohtKUmNiqFdYLanwJjHMqvWebJIVh0lSq
68rYGhuXUzu50xJP5fRIm15LmZlFun/DGWMuH4xe/TYyu/I5vfhLU4A3NqLU3djcvwcHR7hRb3vq
wXwkjvQbhPnGgjJ/TJes2RZE0sZhppj3F0DX4aWR70Ff7NjFkpEaUYmL55mNHlj5s5NxXg//Qr1h
IEMj4eybQ6atxviHw7GA7hO4pIwVe6/P55UYB2riOVXWfsUQJGL5DsPPCSKzPBaljvIAfA51KjWi
X8Mawj83TvJqzJ7NPo1nSgOjtZU0HnsYnV60NgF4VZWar4iiUyV5vN0++7+RHi91OknEi2EV4aZQ
2mxKMjOyUt4ZUJeWqQJ9HZiv2vvovoT2aVoKwooqzbYGawOwkbKSrVfMLgKixfXMQBE8+zOQwiwl
QyAu8uoUGk69gGQliZoDqk0wjas9vuez8XWO2KqZ6UNQlGVOqzZGqqvNbXP5JzKMw3v4jdD5QP9+
92Fia/R3O9fmfTNzByEdBnhJ1E03r93jgGm2wPHWY4uy0CrkJFbu6LpYstwXb/WupUoeg3fBij53
op3mROJnNeH6AXTq4J87MDV87wVuWu6pnNRs96Was0FAhq4/KQfGQVyfiagmSvdE/OIXA9bqmBIU
tURCpAOsRYv+FwNeOq5DezpyPVSpsr9pY/0+IbGIlwywmKktuCcAx/E0/kAmNvO8oL/uchFXrjbh
AWT4/O0ZbL+NHop2srrEqzSO4sHGjQCCeT1gvF0ivX0eeCNpebhVj5aPNl3sUft/JHX2YvYHKUmw
6yJB72nb7XSRJ50ujUGu8lw7WclcTpbol3e7q9ckIBd+fnRVV88vWdjMnWey52mpeUyCZ2F9DeLD
r74h2rUPBlfe/PN6ITbKnp8Ygz0glXEke4ftKPA7yn0w1xHJmSwqtdFte2FzJJoczpuzsnZk8zkK
5rBGUg/fxYWYwvo0NHTANes9d/n2LEGI2GDQOsHLJK8VsY/jeKtKeD7WIKh6h6L8P5m57NxIaW6c
k0Bb3QDya7nYl4uCCRJduA+6/1ARgjBdLoO+3L2tBjTqay0cnw7zSfOEuZS/C1FUOR/Wf468z1SP
W6hTBF1Y/76Vo+cR3nYnhLu/ozm6+HhStahJM14Jrf4i8VM6uKJezhw7V7C7fee2vPrJvACNi5px
OQCSm95voer0heuSs8Fu84im9VbrHTm9/thl5A7DXde7AbOyMU7hpmJBC+A5OKCnVW7V1+JnsYNr
eywDcbdPmHjOGls4BUho1ydJDbywU4YYKU4HvhWDqZ2Vtmg48WxN17eI8w/8/xTJCd1UDQmh0AS0
nuRxSac98KmqNraxra44EnEJ3LWHKlo2Yz1uolpb6+11jGWLVGVf5oWl74xa4lzzplrHE0QxERak
mVWm84wHM18tJRQAQpu8c8sHeLwxIVH9g9+5joxplgJSEixoD76LGIsvH0FEEov0/QzmS7BizfFW
m+CANUiDHwr0W/GmBJN8ZaI4yGFlGLBHOimT3NUPwZP1Az/taWGGHCAUun7B1e/J3zbp3lw8jTF3
EA0JDGsLZQdyMeBhq+XcxRId1KJDIkSLSewIp35wRwwnVKMU53vsZf6Z5fMZHGR9sUcWekC8FNQR
4aHtZBAca2zkenK7QSgjIQ2Haol0EYXu3FiOtPcPlgjGfOAEXoC8PLO+zihwRTr+JT0hUWGdLZuX
1U3Lx/L9OUySFOiG5U/B9c8WFipiTH56oA1UPZaXju5kU+OA0ORd0DoLIzSm66etnbd9YStHhC0K
SAYMUbmSg6Isp4xDpKGe7xeZDXke9oLetfESK2ekggLI52EJBe30dDvwKm/MyqBpyKqsNALyJJTT
E1Kd67L0dqwwawh4l7BW98XSNAdMmOYK2RRrotwcAeK58lKEdClA2xYTqwcF0TCJ+WRK7Mg5s/Nq
pLIXG8Y4SedOPes41FB7Nklo5ytY5di/UPWNQc/JNzEF83MQn3N2+ws31dN/T0aAYcKfpAUGhB8j
g6AfPOIcg8dWFXSxCEGZov3Q4tVYcJeF0Vf1vL2BHNgThCKOZFUkwHEPmbl6mmyuM24s2qlvi7gf
7rkaPn8K5kncZt5uXqP7SWieW8/M/b5otAaozeyVXu7WpKx/96eTUEgEkuPDxRTH94wIK/dy0NhV
6Y+PWNzOHeXkaX6wdCjX+Sxn2JYscf2h2TrB2XWHL6u4ZoJO8UGiseW0by+EM3m29Xmsy5fUr+eg
3MW/sPlf2Tex1/Eb+RtM0wY9g7MVhKB9vjzMTACWqe2mSH4xSC6qdgQNVzCo5uuUPFrOGDT9c5ae
td8GfUKIQsHiMFFT04cU8EoL/w0ftDxYXh+EbaLPtth1iGeo95Lryg7O2vO2Vgd33EH6OFPqIThu
poPBr5nG7bL1kPpECdGM9O+3UvHbsS1x1YmqsFb6iD9nlQ12o8f7Hrhj31hvcVULG9o/DTB7Ukk2
uQRzNm0q1IAQQo+2fp+74HMA0sTK6+/IfTEykVea0pyZZHDY62th7Jsfi7xKVBwbFHMPyKuH40rL
LbclopHx1m1Mkgg7Gg0KZrVCT174WEyg9bsg3S4y659hn9hbTRM3RI8bSerAiJtM0chYXPF4d8Oi
JZ+5IvKETj6mGISoilHYUUS171CR7GS2cf//2q1WEB0tlC4E+6q1M7+yJPMfAFLVF9rsMh+Vd3HB
bSom+GEoOm9mAVK7LAUIcZsQp0AgAsdZc+cXOawK0xuTgouqhLAenVMzY1uFZja0t9mawSonIY7B
wdaZwTwrPU7rxmbJiNxyBZcThUObzy5F2xk2yDjJ8wLwHFGRQhYNYXS4FCe6MN62+630OmRrdG5m
vfX0huesvMyvc/DuB6fKU5M9sLa81mai6+JVO/twshGhig1RbEYzCSDRhO6nlAR+g1v0L1tkZoYF
lpXP/43aOX7vWgJLfGDFNbr5x4gCGwTzjeSt2nVzv0+UxQ5hZ3oqWvnHGCavNpkTS4zVx36Uc4/q
mEZ6OFtsL7qTuo9PKhnMqdvwoDiWVwA7LWTaI/c8BEX9LSbfzddDEpZwz5RsHEHPe3qdeq497ogL
Be36NUh8waBk3W2s1P9WGQFNwYWFVQs1y3ek7Qq1B8pENc91cEgRnJMUEBm1qoCkF0dfZBUIKsRK
L06mvIATj879Z0Zs1eiH8Csqzwh0JDkP/3nKKLmHFon1AKtTCzkoSpXqSNrTt6zkOeO+PV/dUnPg
WULWsTd0MTOfFm8z86gZbQVDzkXNF2zB0RPDuLydiQDmICxs58q1FwkMf7GJrglAKoXYhmFXdaED
trkUvWHWO4bGxkee/11Xp10lxLLnb3LNQSHrFI8OKtIgUZ5c9t2OkoDADhoKND1iG8Bra5ffQuBw
o5ym8swHnGsJYB48swKyC7z3esBZDoklCuo0MbGJ1uvC4mVw/VOFpTgeVsSbz6UZMFR9VvxGLyOY
0WH2jHMkxsFbA84BdVf2Pjc0kb2k5pjzJu8guwd9S8hN4BR7FL6JLCehSKOKLmlymQ5a0GXWVjIQ
1dGCVogajhzLzbtq+x5Q6vNHnZZFot6los7t+ArWViO/2bumXU7MgY5sygtj9l9MwZUIlW+3FudD
AY3bWwYgG7ZHZGB/fpfAVPDr4dN+NcGaiYphJqWPrX+qUfN57P43JbIg8R3o/OkULY/XjZ7sDFx0
gsOiFvYA5uXZFf61033ofnSK4Kgxbe52gfzy4QH39DshQ19tBYYRQa6xbM8eCYDdrzdhaFWYjw1z
Tl5ff8j02Ja4DVXbG1jZoTAizUCuLtmUKWx9cl7LWot24WRHecumN+HWPfiujaZDCV1MpZwmH2z5
ZoljU/FRYE1N+RvtJeVjeV+qxJvaqEuOUqiPbdDqWd72mwBWUoihI9gF5E8uxI0KLu90AYhFJEW1
icSFMSu4Or73O1aKHjBY71R4rJu8RuaLMyoW70QGhMX+M3jLS4bKmD25PUibAjhI/agQ9PMxZkfr
VKQUk6W0n72D5MymrCpCEElUYEC7+dy+g92xkmk3tsSg8D9M6scZnQ52JHYUVBOU6q2tkIeZ9ep+
+6iWQR/34W5/H4nY7rWBdbF3uo0hhZCVPWwD/FoUUD+cIPSjjRtSdK24bPCzvPWpfkW1xE8V4IwV
DrG/YQHof6dgTDEjiXJsY4fC6AJugaz2VHj3ajHjZuIGLruxMds8seZvw3FCV70FRw7vQkUeosoM
QilpukzRVmLwwVjIbqK/hWRTZDIumsAcBh0Hp+RA8GgquHZELJ6Xjlrn2UVNl4RCuwjSxo2uFnJn
KZJ4SWEn7p9RBOVG+SpTizc/8yCaQNEKxsfYG/7MdJgm5Ey/szEcgj9CjZwMQjhnB3mGBfxUZosh
gytkUMDRVbdKWWBAqnoEbIZlTlWxGw9sXblW0yIyL7nfHlWz9bytE6C5tQPwg4LXubQNHKAnrap/
juqwYI281F9FOc2IwTIOhlKWRh/Oos0dZaZBHPe20iRr6BiW4uT3zQF0sN7QNxATR303QoUqDfNS
giII1BbMfeV1thF0nokpY7JxAugmghoFn6wepcF9+N1MlKOGov9VLT2pENXq1uUfqBQizD55WSmC
HTRcO5Ct2fjLCowJghUCvQSH91bOArrW8PZidhsgSSe2PisawK75b8pSfSykPxGMbDTGLf7SSpRI
4yg75iGqmQYpV768WYJhTWWLjmhN45GjxeO9q9kK5SMmG1rwe+gSX6jfTUFNU8TwZ+BAq2+xct1V
In9/FCldu2E+FsFJCCMLaSfnB5OnxllzWJPv5xfXrUV9syAtrrKG9EX4MrKwTxgq89pJkRhRXGbR
+v4PO4Kkjp4s9pRxJydfSoPHryPekJd3eRw5NH3rIqA+MmXs8O9VtwCYDZgawjoXnwxVDkW4UVtb
Sd3FMJmJbZAb8/gycauXZg4Ic1xHyPPJNkNqZXlOJUo2/jO+kV/DgMfqI8QPum/31HkWD4NJngTJ
dvppPn8PNdfpnlCj4HH24t8MZIN01Rn+Tt/N4eHiGznnyqZFncRgsBk7uQ6i1EcrDrYGdZGJ7sxB
LB+VaGWkMzeE7p4G7CG7kolVQ1FbyeFPfhyUW98Ve9cEZw4oQgHqTVoa9c1hncFDk03AFXXBFZZ3
c3mT7sM++3zeAEZlqK8E1kdJ+cL+etuePcxlzBBxt1dGowi5ycugbWqBe6AVofq+ggcKv7/sbwEG
DDtFjuQR01HOzp2Z3oTpCdj4bVoMxyjzTTjz0P/QEPR5doEnFKWXMQdf969K3NtlOm7JXulUfCW8
BH6tjCG6axgYH7Nsdq0NVgLnS1piVKqpVpFL2JXOLxD1CVYSeQZC73duj3uOhxV+82THNHA4syBV
8FQWN11mumE6VmElyUxldmvR2HxiUMOcGL1l5t/FYqVrNM5Y73dxA45RphHqmSZvy9q+NsciFJHR
MMr37Xz3VV8HkJRHrdHH/Blz9t87cRddsLQXeNKgFHyvzBnWOZo7mUVOdZY805xjN5vGlc/O9WfB
ImTAqG/JoyYx4Yb/epFiFOgmo3Txp38k9EtGefJhf1wbYB5B2lTOvQGPPhv8ZzjaD31Tbd7/EA3k
loFwe+HnEEa21Qav45x1iGvRZ/A5oQv2ETfn+OCNu+n0mU9RurzHPXHMdb6dOJ5xOCdKfEKqgL2L
RQnWtotBg9niugAsFoIsGAkULLhkJAD6Oc8XFSzQFOcCwAfzSICPyoKSFifz3Z/ZupER72pw9Bo3
bTty8Mx7R+fKtqjBOvn4k44cxTuuKaoYQQHnw+4OhO4lPq6jQnzkwGSVa+P6lu0y8QQQi5dk4Bvx
wd4fYBn02vSAwuTYd+xyijlPL+z4VlILHGLm28lNvx/vcypcD8ildpNnhM6Ch6qba9BL0v4QenNn
PeV1opwcQ+2vQIlik2EfyfKDUMC/ouF1lv2l5TU8e1NIEuJJJmnryW2TBSVI9zFzQTjlDE5a50WT
nt1dsEJgmbwRGczbusTrbB7wy4UkZ0fgxOd8n4fPRHZ6EsZDpxtrPT+u54BFODipJKHkj81oCUvh
64WLPcOCnjLwfpvvvV4503dzZqyz/8ss75wXafUD0vNiFY+AEAQR/piTRcOkkOCKuivfPTa6HAbH
/yGDmC5txG72bV/mvXHPAHL9TZrgAxs9EO23K9YvlcbjJbtrxupH7HdmfFbh9JYMJaBPIj+ktjL5
3sUHeNPszmL/7ZsALDiAqDaB5jZhfSMwAuSOxq5Ef710LzZLb887QTZuce343xw++KyqshYL1yz0
/WeB032ts5ScraHKpfx3mYTSBTBzt22moTqRjPJIin4LGjMQ3FxPvSOHvwLcWGa5ZJdWi4XaYRbz
Ji7pajXEhpKCiuW+1/6fx1o95s4eMElptnQ0MlclcYE+xboXMuZn3TIdFFcmhKTfduX6SFkiUg0q
MN5I1op8zkCznKj0jmY1CsdA1AaruWTiAytV54yHFhvgIEAnocUTmxUcYgGsN/vhf4qw9wrbZlh7
wLlAjT+ZTJwLN/fl0JeVEq4QdwsAfaigdUOwfE+/a7wmoXot6aUxAcR0OWXxCResifscXp/YWkVC
MGOTyT9Ax4wc6WYSO3by4w2UlvYLPg5GHrDXxURp9ld/yXPXBc26AdOlgcvobLSBV1fTf4ggqNG9
UnINCnQnuxtXCKXjHchcpoxLtN+hb0FwA8jvn/OlOtHm3VYc9YCFzl0UC4lApaG7MfbNDdGycqgB
kBbwwDUnmhnYAkiNbo9xnxVqP7/uYBu5XRkwN2XswLV0uil+JUK0tFOESTU2J9psQxz7L1kMrqgW
xU5xo1aQfx3qNjxVu2BbgajH7364BA/dtWP2NeJKArofZtUGO2h7il9fZSc7lebAgGeBV0XLYAnk
mIzhLA156rirfNx25hKANr0TT3kI8FZoepWlaqahGhab1tXrrFKC5hV4ZElXU2tFhr+kunJNLb9p
dfoLTGrfoUnkD4DHfb9HgvkeKb/yKqHt+BBWwKQ2GMsbOVqlGU5LuXpq7F1rGunBZ0dQg0S6LLH8
ebUrTZN7oCduLozKGea/vQQnwraIoyv13ukoAsT2nM67R3p4SCvZcTQLjBITWPB/9WjVEZBkusbz
f8a9bNPn5jgRxm4EcMsPABnFnTb97zNZWASGr3ttX1iNxRS36wovpgLPY0dcVqNc+8sLTt5wFTNR
K7PS21WAAVOPz9Gqg5L0GSRSq1aDweHkOdf0NtzvLxRKyB+kgjRWslvp9ZX9HPnTcOWdjbFZz0jI
g/rOqiY4aQzbzxomqLX9ysiOCeqbVxyENQEL0j3/q/2IeKbjapL6F6BNi91CNs0OA5c5+si9CQkL
NaQMsVh6CPm5g5Je7o5FgYqe1gDnMMQ4Rn7QKiz3hg22NXxCRJVJhEePv7MURlJJvF6oqGQ2iM5d
yZLWmdG8ybomSa6m8DaJ6cMVeFxbg7y4Pti6jTPxxpCEUc8mn5SXMv+epUTNGwHRdoZ95bvDLlB2
fW1P85W5IzeZ/BQdFd1305e/XT/ftyunkAOUIssgkCQFjOiddLefA0OG+VCe5P8t4xGI6SSd+uDN
+MNEI2GYDmnJkkLb6Zo/i+ZWJCZJuIx1BYHQK1VVwNWI57Gxp7cN2e8tCYu8TOo2yBczXDZiEo4L
tqgwxolclqQ6uijgfPZOGaWpvFhVCzc2GoznocYgoJ7J8Ru1OoDVVksndQ7yn79IrqvX3u/q98rD
NnolzO5+nsD8/DaGIOIv1VteBTvG4A5tSDCu+WTZbn5K3LMQ8Lx3qOBg6dnuFJesvBbzmWzVtP70
g7ySEfth6VH/bUp9tu+hTiFhV++grjCW9RYkI0bsuLHf1C9AxjrXEHla0qjYIpNDygg65VD0Av/i
+7cxHfSRp88526SotA94GyuEzEc2P2oVh9EG7VlchdAMptSw29ymNBXrQsBerXkQmXEmkAsZ1tFr
7nLRuM1cUwVjne2mNSm7JiOn4Evf5z+QpoEo2mSFTdPjnLcXHto51Z1DZovSfzjKupYPbAvQ4hW9
VMi2+U0OpCdD4HtpIjyrqyWY3OsPXYSnn8GPZuWEj+eOJbM5tNwEpP+L53gOFORz6g6/BC8oDsPN
jaCr6OMgd4OhC08iKX7cW1SYmyk6XlKE61iNjlNADuE8cOUAmiSR/3dLj6zDWTE9i9H66vEq1sdR
6yHsuMz6jXxxfmONHs7wLXKYzntKWXEkqzk2ufT+ROiBgw9EDtpJIBiEUvnorFHBVCxooFFVfDX+
e5PxExs/VbH/2dCTU0SVbjDMFsQOYPMSlKzTnmtars0ZRSVaJKbSjv8DvVsEcDpeeQENCGcWo6jf
ZFlOqi+AmiYExqP+cbdbAXYOgR+O4Tr3JKJ4liOH4FavEU7UYj48KCQllaHdG8NMCC5TWUzCHqb3
Jo5jRo32sHRebcGZTEMXPii8POMgszhN3dpf3OLaVvu/xdKSLH72IJj10aTH/WhdBreVArhk5Iev
ll6IFBOCwlkfrB9vcC6kTFi4UitvYw5gkkwN9pJCbvmpyZJc98hd2r7+z1TOhVEpd8pECCVCh4IO
EMsWf8ZP2F5DRO8NuvoWKEofiUNENA2qpMW3qRImwjhbE8B3Be/Yz8fMIdLqAMM3XieMXjRT+CsG
E67Axfz2iT87oOV+CAy7eKVqWwBUrUPsrkn+N1CDPpgdGq635MafOQbfAwSJMz3sYesDt7pj5Mht
gkwrM+xWNoJMLniz6PgfLpUmXVL1NL3Kog1gL2aK/oyt+V68qy8cy7blBKHfL3D31REOR3SxEVQm
54IqO4cK/X3D9HDju4pR31Ofv5XHBcnRgyv3DMScxgW8r9y+5Ui6tDVdgW4VhsvQafKTgyCWnmRA
cKTfT5GAMMJt35wOdGLqQ2ZqLS7bTrSNV1qcPv9PHaD1uistuAt0a3VNAItF4sRmMCcu04/RoCab
64aqlL9Jq2JNhFKGX1wFTrhAP2gpsKQewVWJGhhPKtnj9llcKDnFZ+x1FyJ36nhad0sBCqgPM7Uw
3aMc6zi7S6LlyeKRs8clP/5UbPiSZ+EDIYgKC2hqJ6a98gchMoHohfdrhf9acoBGIkHJNsBnNY9Z
dZHw7V0M7mwS0gB/VljJLm8CjcA+Hiw1HjF4z/tqpAW495iqvV5ZcE6umUz+vdEWk6onzzL5O+Vx
UB6N3kDxbVW5RSxhQMU6rGggkG80f4uMzjVTVcEgAjMC6CX724aAAeK3KnFfBUA+Ln5IWj4quM0I
8Niyl05zr2CiHk07p5Lz9vt4jPprIC6RfX3BjAranSzp1ZJon7Kb13OcKk/lXePoGpbwcELDbec/
tH7sNcgb0qksxFziVqyNAlrIUi4ogqWkFc8pVL7oQ2N5EX5i9gI/YP3g6F8cjxNAPuWuaxEjaXO4
GsuSKYLLSL/ZoKOhwLH3aiWq7HLAh8liDvwgs3MjKeOyjHQ3wy82MYJte0Bo0r84sQQ5gtbSzJtx
p751Hj2N9M9UTOiYDebzJd0H9M0YNy7rAyT16EQnmcLZOhc9pvHWB8DbsSRPUdxrYk29eoYDYTxx
5ghcQEbLDRtylOVNmPtPwe/uXI1VpezhTkArnuKbQ/5KpFkr8IgDL9xPuBwy8yfKlQDiVRkrL4HA
QpH6ZERdcFnnOZTyIHzsu+8Hh7edrvJzsbNJnwCVrGxTuXJ9RjZSgeWl72GiL/Oh7ynZo2lUBgpG
SAfWy0f9M4opZ7UoWtEQoGDF95Ae5PqqzCfFr7kg3Dl3XkOLPjVvpdgvAaC9rMKI1KFMuFM0yjeE
uCJyL6jY0OxxXR2+ALvoG2iof1y2sx/06Cq8Si4pmVorm62oCaP8pkOJRaegU86DlyAApv9043R+
7cF6A/efWzc9Ywtyd9LKFeGORCgwijVZbijk6Uot+N5w8hw//uFm29EtkvH8qDgX2zEUdHIuhZ0F
wdKon5N1dA69dfq+JQDtsr3AsegACHBq9jeYRh+phRk+yKeYsJVBXBFkUiv9e4sIkU2zzYrBnJjw
IOj5n5q/uKFOi7Wby1w5hzWAJCz2q0qEVNdOhXWPDLjTymSeAeFRvbluNx3gNYazAuTeuqKKDeRc
ZsR1I6b6EcK4pcYLJfarQbp0RWUpYmh0d7spFVB33eJy+yrcVeDsCkBJMB4q3ZbIaOiawQPotpiF
y4nvWlj18xk44VyDt7Es53cTzMC6z95J+P1bzqrjJSgsHTGbKJg2o0AaXMDtc8AqiP7borrCqXio
vrDdtPovf9K0H4EvpKaRTQOYGdLZI3Gxxgg0VeXSrcBJObf1uoVZY6CcPFctwxsAav1vkR8taAUG
zyrloZGx3VJnkp/pi0skm+tDZ1SulFP6mSqkCzvwGip9hmNzlBCmcuamNrU6v8dgkfo3+EaAveqU
X1DmLozx92mj9f94l7zxWs4tm1hAWos9tnBqllMHEicx1UKAQw3mqBbydbxvWDESEg+M8OpPH/rZ
t0nuG2rZWCZdg7rNd637SL2Swv8tpvZ7xcmUZtv63ThTJCjJjmkLvT3dVOuR33jKwde5DtsmtVuC
mOq1otg4IHH/zP/7K+2kciBO4fakeXBNIuybtRb+jcRuzATjrSmttN7vWVe4h6xODnr0SHnUtaAA
4f0G8LbLnfeqQwbRDdmwAIslo0MtWfM7wh0K1rKXf+V3tqUvE292LGQ0Qt51QCcuBFQexff+IZLK
dmncvCoQu+Z8HIWxpT3ctgwZzDwm5yly5cjIAHjVCx9KqjvKABq3cbVlB3Qoy6dsxyA2VVCWy1MJ
DXZsTWnN0U3W6NFqyU4Oi1Yq8Jd4OPAAe1EXAxupw1k6etNB3nR35FgrqYcbf451xMFGrpfUu379
5UTAEISy2515E3G3lH17orrSHeu58zEpOF6r0gekLEUfqLv9LpkGFR4fLkMbT7UMx4jBellFWCuz
yqiLwTxxfoc8faGoZFBwNXf5mH0Ukedytpv8Nbf4gcoiy5X2aOZGfdcC3s8QSH7iccGKMqg6VvIJ
kHeUguIEAMKcV7wuEPhQa9ttwq6CJ0DuqBGyQmpjdoch2p7poOgTVOrANnA7meszJbOhgiX24num
DGbFb2bAHWlit+MEosYGb+pU8WGtDkqDVteP4DemNy+5EFZqfSIiQ6r+h0rNJ/FXMWmECadaYyTI
N4H/5HqBBwGpgXLNCnuEJi4ZMbmq2P9Tbz7w3B/vXgfIOzmc5OB175hdc8fonW0Ks+SRmMQ0TosZ
GOumAvLbWny9NCbqHlT82vQ02pbWdYP6DlmhvwaRbVUnvG19YralINtllytfkqyai5gOcPH7gftF
0mQF6b1IUbfQLRLGj1Qsh0AuuOG704FLkW3dB6CpPoka8Z4H57MosVN9GxZs7xNG3dkmahJ2WFee
mHfOofmUOY//Yh/WXCnQqEm9EhYZI8JgxpERN7/X6wuegaDsGWw0G1i8ALtMGtYwQqSCPdOQ9oIu
dmJaOkNpRV0D0HpSicLQ6bV+J+BS+om845glr7cCQvPC+jA6qfzeTdzN8NojtibKAo3063l7FpW6
MzFd3GuKYyYEOklGHJCXJBoXlFRWVOCYe+25/FeaSpANmG/Pw5MOuN2GXxMDbyvxCjaKZzEn1HXR
ZeEgRKRGJMaXguk1isiys2lmwqzzmX81rC9tWlMUvBgi0UvevKXQaUWAMxaBK3O+r/Zb43IC7FTO
/suwvQ1q61KWSnqK0yboJllcIG6Xz7WoCvvXWwfFc9gJazBv5CI4FgQ14ybYZp8Tf1lP3er6W8zL
vqhrd3rMFChxj0d8xI7NkpkxkNBlUO0c8LFkhLzKzYklpuXkvjMssdJ7lE808bAqZcrBOP1bHLfK
Dfipno7FnOTG3K1L5P2Bm+KHrFBleixrZoY7JKD1/m2rItm69cr5n8gBl0HV2wMWwkRzXS4ubcgL
3LJh5aYBhAqWdcYIerm78IL7pIFi5H/02w2KxA3DZ/7p2nl/DGtH/6YF1KbFRlTGCNfIWYIHnnrE
3SXRZR9j+R6w/EjMa/c64TPh42F6JrIPPbgrwpF6zJ5IppC+XU/JFip1ANwtQ9DMIvzKbwc++kEd
ZJqI9gv578wXaErc8x2XJYfISWf3K5K4SFX+l0w4WocUkSm7koVQi/ZPjYD26zxtPRN+qUVKl8a0
84Vn1qayodBCJfL7Pl7XtcMOKh9rMjjGVKXHG85oEuYWIDvC/nps28r3lEohclvCnXy2GqkCju4c
0KuM7vhHYp7iwMzjvWLfj5rX48a6V8ejXPfupbKqvuINGoG4HswQMCaHokt6Udi9C496vbqRuzFj
0iBkEHNJ8Ccu0EY6RtW5PJeWqoi7zEJz1AgStyuMHbveXZCvM5e7X5/+l1nSDGQ75/XsqJilc92H
VPoMSbk7BjttqN7cm2F1WRHlW5FRg06He2p8OcNvkYrpQWJjcnCS5rlE9ieXSSdCYuHxjHQ47MF1
Fq84BS+JHSNRQg9rsXyEz7FGHGXwrqUcjDBpgBMKfM+tMlt7R9l3AsrcJsOES6usYDXRE+56stIT
S854Xu+4HiAF6+FSKWJKUhOPOsjo2DrT4uUDGkzf36120OIh35wmHDamb/or/W3GHVjjcXrWdulj
/e8bIaxh/AJ9gnU/zJ0DRS+gS2o6n9E/MM3yRGKQQecNDnTGzJuuaMf2e/z+17mHhJJ9k4nXxf+2
p73X7MIW5m+WVf0CbcshTH/WJlXMDi1cBf0b4kU9tNwxzWyUSCGbIrSkJCSZHMfWJYQ8WoGnUp1F
Xag9FnRKPu6BaPcL+nUITwhhLb2kuZgCpYWu+H9JhHxF7zKJoKRauvhFE4IaD53whj6hAObO7Efk
jFpn/4sWAIhbxEVsCSW4bcG4WBSGy+UsBTSMi3EitWa6TjzvlI3oIdfUYZdJfa7n92FEPjE7nVLI
XY3ptHwAfAMq+/lT9fTFC7VPtzcKufLFB4uOTvqJYCCFqWphVJDpO+dphVbAi79BgGhx48urdY1F
HOXJbEc5DNrmTz46q0gMk4ZJAD75M47Ito/iLmaLct0RyFpRlqeUT6GG0A9HJdHFe7RkcyWgxjZL
fPn07cHeTb7yLBEFDuamObIKoUBFC/v1DGCkk0e8JFcUlEgx4b9zCcLecdanetFMOXspVRJAq7oJ
7Y1e9Z4o0mjliwBw+4pvnXOR3Zz8+8iiIQWECzYT7QFYqusGRbBNMn9pQebAWVzrHTFbc+SYmanQ
4TNp5XbIxy4MSJGILOludCvQSVhRsFfeyTSmp2A/Nwk7/XlG6NpbcDr2yinh5GwoW85icbLDofQg
h535zbMkflEd17oOjGBAJvFooWvG7G7fw2Um9kAkEHIVS3cpWaVHLBpMZOpUnqrLHcCk9GR/RmWh
4ZL7nwZHZO3YYVo9k0o9mfCQ9wdUwqfQF/56SUH7e/9w0Kou4JhNZwJD8We94i9a1ASZw2SHFSyd
U9agNKCsvKZuqzC+J0RSJGIoDbokYFjKOXJpXU1jmXkPqquXGi8U+CqG+xMrxTC3BRwQ3BjCDLBk
UJ2Y15sFEiYnDc0/VfCxBnQNL92yxXc9h82W2LRCK1FKhcHI6y9YOYMKBSPiTVOMzHlhERZOp6k2
fst9aXVUvfSvDa5Cz9jXLXygnaO8NfKG0g8uCwg8PYm7E5Ubovt5u0vWGH1JjG67Cov29s2aqqMt
FfwUf0Z8RCcyiDtxybQKGl9MzdpICynrc96IVNDB3Zf/gB3TS/R84XabKuAZIBagw1KuKd1Cbh32
Is2lFT2xU0FWjgpTt8WaI1sgWiawTAXRIePCsHdhhj+p0XmbpJkvn1Nd4TjfuhUwTOnn3DiWZTYX
YBuyWeT8wchXnMRVeSX4iAmPpt0MkNSqbEobJnup0io3DKhQLV4TV8rS5QeHyRPF/3KirgxtSUB/
D/5GfZNLgHw4oX9jV/E0BMRGJMw2VrxLOtoq4nxfKuNbsiTSM2WMs0P5RAgemEYAUfic6sltvUG6
LoHRF11E+HIzGmHmtW8Ci8sOlJtnQ/2bP9ii8BKrxRE4FKOZWHafyNpGmKdu9gjzjlkvU0ZystMD
Jch84hazzhvKg62x9FPaxt91TrBTtZs/Q+aJsnQJNr5O0qYTxu8tRHCYc+Kb02hkBcAU1vS4WKSU
eCrZ1ZNaqIa2C/azxENEBWda7HaqpTI8OQsFbUCZx3nz1c4hjtqklfJiPi559Cwm2fJhJX55Mpk6
pMWN59nzvb+cNPQb38YXZhOjmfIMts37cgwn94Vh6yjwk+mAAd+M2DuVylqEMgJpbE2CiXLiLC3Z
y0ThGlgnztQk4rNzLPNVU3AT4jkg/PUFiJNZo5LZGtG1/lgtFucpqAXH0DqE3sGSdRkf9vAeCobS
h+hDCK2BnsWhXvbamp//90Xcx+6QCUuG6M3Zu7PY07MaCuPwAfKE1azi+qPtusuj//YvWVtAPpxL
/9UwMsTRyWUDv0LeJMYVUskzpfedAeL7YEbRXo1TCUB1nmh/RU1PAxx6dvG8lYt/boE1ag91Kpl4
uVfzXdgqxYrcvol/H7xVntLJR1rWYr0X85yMhDgw47XISSNpaJkcJ/ycgcltmcL0FYw6KFHGQrvq
xWfB6vLhQqYqVRRoBO7l3zKvZhN46EWeML5Xa5BXKZzOPafoMUVc8xLpXKwhPzr694zu26ZruO1z
n9x58KVW7AedhttzHzK1dO38M9aZk5lv/ctLcOjee41CWzGM7vzfP1PtsxFjJ8NUboGSF5mRLQIb
BZPUGF9jCR1R9a1MQygHsDppZihFQdtQWzooVdeUvaz56UvhU6u/c6cUrH7gHMS+bEFUx0SVSZvk
Bxhywk2/LEsvKMjrw5ZYiXbKN/xW9FJlUDoZuhbvYLw2sRNINM8zFr8sAgb3d2+ybbYtAbRnGjU9
YVyfSRVZcWVNHsP442uFgP44JLAemp4cGLvlh8sQ+0NUFrIQBKpyoM0Xz4yjqPSEjdrAhTvBV1kl
YlDOW9bDch4zeYd/GhbqlexggIKhE6BaeRzAqbIfJ4SbD6Kvv5sGqQ4m8+NzOaQnuzuxKkKk9vXh
ElCjGtCPpCW4agCXULRJnoCmGQYJx+cEjb4zHOPygQ0XPbBG48QS/OJMp1M70tUJ8Md/EzTRloqf
gLnSl9SSCj6BaU5lRcIC5wF76CKnqHA3IgFTfxDWH0KWcB3djGAcfytgaReED1IAf3HO4H+D0131
fCWyW3UCYKSUJvmI0YGU2QJX+3vWDjg8L+n8Qs0DRmPJcRuP1eXf/5aZp8jeJP4KSVziGE8EECku
JGpNJBTFuLrLYetR47CpcvmTWGebGQkHmbijUcY6i3opMi4JYSgzSR1Qe4NBPvEbRdQV65+JUCvz
HMaN0ajxwZsR4eBHd5r1l6ECFAnE0Mk6ebIKCF8eXo27jtRy/f4iEXOqaA1PoBOsxwEkKnLkTPQo
0sSMink5DlSo+vVsrJAxp9cYaFC3T6rbHeveFyOnZAshwPUJPvHKh3QCX9hzYAgMaGy1FwYWCrGC
iswsPnlIHckiSLAas8TrMR6NPcCA3FS4b8JhwjPXyv+1B0djRcZu1Leh4L5si2VfaR2+wzvYLeRe
waUviddryOc/8eFsMdiyJoPE2yaKVtsvT6FAEvd9oyHS6yT3RNyrXxe7MPw4LbQt7oROAV6ZzRgC
vBo2wqop44WlqO+bwQq+najmAdKpt1phPUXhV9s/Z7hCCyrYFWiGHJ6i/79+YM4xVqDLP6+8MM7T
ENJvaZpRsYr+MNxITJCUcWgrb1nqchr13VpP0fVApmQOB4mZvtDLfNVY3WOTYozT/fh4ViDKlbCI
Y4c757bf87lvzCD70vYNIPiT3s6R8VNu/ygJgGaARjfRnkxR+COJIVNZFBGb/XBHIytxTMYzIxYS
MSjRFD7KnT694TfFLnIOWoYT3Feurt82XRH8rTZmp0NU81ZotHDQPYzBxNQWg8jjFjaQg7YOnza3
WdL8lzSLK989hM46pPvwLPJxp0/28cM9Uby19678kYh5L56Udm8NWWP7iPppc0qupZZqB22BG4Vf
2abQRM/ZFcCagB4NsCgcU+7jCF9+uaSV32ANSgXnVPSyKgQANPevsFIrljzEyTX7QtwzblAMZmRF
DnCOiy5T+4LIvR2EAtHqYk9jzvXccnLxlmaL+7KMZYh6A+M3Gd6MkMqEghVF0gS365ES3o2GdNWN
2yLOCe8/k2dB5dPIcicU5z3gOVFZ5JUCkMJ+QdvqVXSDpBwdk5cmO7lfhV1mjmceHMGTdgBXMFiG
I2FjUu4Ckfh+bnZ95CVBrqUf9d1WQ0d6UefN/ePkxTZxg5qhujysIkOXTIR1r81Am/PhAXta1Pyx
M8ck1ZYOnJgg8BW9vn7kO/cmdYe/AEjDlPxn1AzA0jTKBtJXLSzbYMOJ6FlXxnSnQ6H/miRf4FoW
5fRN2QRjD82hBS90tpRlst1kUAT1COFiNAN3+l6fHrmL+9zxFSiUpsukw9rxUVmG2Uy69jp6fCTX
uEMTamW24dAmmrQTKWngyDOGg7rRVT5mFL+ZyR0DG3TrcaUbkkVo6VpvFbnODzW9UbqLI/XUmc3J
71iUVOXSlQJ08cnnygi1EjpgvVtXOBuQ8dYtNesYLoDrjz3nJeH3znVFmAZzh10zch5KJh8YkTrp
Yi3F6nNZBSgk476cYNGyZ9eO07vuZ7I8DRl9SMG4mIdd+Unt7CCdQYBh9yO0cE2dwEtJsY2FCgIh
Vicn8relIVVlK9Quvb6ihAa1tZBxPXcX9E69hmI7OLZi4eX8T5IVxvA+mRYHdtE+sASMu60Vs+IE
u6l5Ffzshr5WfVWh8eFQ3Q6QQ3rqNVKObgZMmC4fAxPuXaKQh42RM3xl6OsvjQirzMYwgYEfVakK
ANsJU3B2iRnaZzT+TE1D+DEz9VLHQPH6QGFSX2OJMO4Qa6bRU9a9QjYIB3a/f74yvvD9OGq6YhvZ
J5AfM/1rXicXbYCn2PCW73FE9HzhFTO5jY78sV8mNkW8B4kLdfPoz83UB4usTvDChvSkjV6Cyany
fQCs65tvv1TB/zSY+7ncaOwDdLQJxZktUeUwO4YRDDBbvuum4V7QeYSxjubsJC8goA/RphLOH4cY
Dx0dxQ6FiWkicx5wXEheiBwb2o9Rw5xboNn+eeOV+PvIDt1VwSwAH0GaEdeoRwely5NOeICfxN29
x3sI+Ml8SB2Kslpqck/7hmGKfuP3mvUUKCLZ3QdS8KN//HbN07Mb/lLJWW3xqtUDAiSrrmdafJjX
FYcYQXc4vEb+3tsXGTyLS6+Sqd1ZQOFqebbxf6HoeCB6gTdTDV26W96fV6mD29RbmahE3B1km4lz
85eSC0LtQzd75CAO4hPpFAAfpZ6/66ZLLwO2yfFlWH5OeCxvHjk/kXCgnLG0Dy/1D11u4Vclenrd
81kJGZp4lMtcSWL+soWjT0RaQHFcIZIfwlf2Cjl1Vob3BC4DaRGUyURVUyWTz9EOjXSwEkGN9AQF
+LUaeXfGpYANDJ6mjX0t6PpEanQ4opncFe3mb1QwTV+dBq9rowSNJmHY9NCuLF5nsbFIVvUsBPDP
n/6Xkxj5nY4K2HdOvfDVjXypWRlWyCa8PG7tySscV/Kvaz7J56BKylNTfITkVszX2YeAOsPTYqt8
WVEb+DqJEsmGZ8Y7rVjd09abD/TcuNmRRaOC5raywbWBbDdVRhBM/irMYOyOzUdOMoGtfOx1zFzJ
O+4mzSKdiYJLIEGzO/oHSihKALf9aqV19ucgeWsyDc/iuPa2u9yVLmyebO1jLbWwLf5EbjKSJ+cj
O5ElB+6VYKpNNTDQyT8tvntaqznYaS6vzA6tBLp61Ie6CHDIRzJlz4EdEkRXh1sQ+FSG8FWi9w0f
tiiegHpk986bUJ9nrYAytO7XfH3+Hsk0gxubATgPTWBXj2/7jQ6RrvTg8zqEwm2352A+AQWzCs3k
deQx78qiGQdouru+6x4bFsx2T9GztHr9lG36QzmWWEinGuf7/hkyBEBNLclZ5fCgy+l9o+T5QQGE
zGF9EJJ0dmPoPiBzalOR6Xa2SF0hr+Sz2wPiptoZ2WtTRgvV+mLbWErritW+yz02H9dt4qdN44Tw
+HZLZndoUv7qJJmoZfG3ympB0VYKOY8vJ9VDJ0//u0loTfJeKID2HPSXqlw4kXbjp3X7PLtkirUA
E9hLpS7ZwGB5kEROrpy8CAqoHZvTAU1qn4TOXeokKvmKF7AF8Em3h8dNykXWliJ1tEobb0me6e2A
VaAO/R1G4qyUg6C6cTDabFB6XPt5XfemqqDaxBV2AyBxLinO5sTNnD3YCxwKygVqW1rbnHVmmVht
V08DIIBGssi71KbY6lUdGcjMwW0K/L4gdHg9oTSLn+MgW5ag1ZsiUSuVoQVMUrzrPSSY5I2JlaRa
mDs1FuH31mGIhmYSW5xElLNRfp7tTSfSeSQFlP52/KCg8aCVQSUqT9NWezg1c6odOWlrvSjg/lfh
hgP1UsbtRAfruFT0t1ruWmY9sN4kmxeLY0Q4bdroRhiF1MtVZD2FTlmoaJz1xVpecliO1CyFIRQ9
ztm7PHOxfd2zRcrwIfBVKpK3lxymlDqcdcgFLwdkAjuKcsTfbwNin+XrRRBqesSbBUN6LM/72vug
UmWLeq4ctNX4I1kSVddoSruoQJ771tpryzgdKXmP8gRbeW9ApK74HETsruXBaIMUAZdgFlzxZAeW
8RgnO5cejnYoWBSmPZF7wPkbxVO3KNNZLPTs70zsgU4Vboy5M9qW9Le0UwXHidsMcX4FJ8/kqAiy
PjK8L9VmWCC93xZ+Is1njEO5gFgWU9xmyu6BgSLwBcpU6tP1j5RJVvr4w25qt2sJf7UNXXlZ8RaU
AEuHV7uzCpIySmoeyj9Drjihou9pjliBSsYhWiftGT8xdqmBSOChZ8Jmph2OQIUiFhgNWM1cX3/A
ymti3jl2IR34m0e39uFThfnoejfEvxRr1U9fVJwxIMBGbXdW41eiG5PgD04nJcIeOJeJ4BzJsdxl
NUsocDpkRN2jT5ty3NEPMp2EHzy9G7iutw/RXOSptJKkOreLuRqCU9N/W42IikxatCKEcqRf/fOx
qJ9Tk0PQb+hHuEssMA/n3csCNxDpgYRSO8SAJZhsyfDJjVUu0eT8B4L2VRJQDDyrFeKq1NIwC4y0
KNuQGp+aOc5xNMyVvuV/RDoqGaHBCSMqnh9pfSOaBgZ/VVY1T/8gEqwjS3SLcyISfT19PJw5rerX
rhtgNN2sv0fdBmX2YsYE8Uzx3qmJv94brsXBD4KlnQs0/afDA/hefL94SfvH5+DDA8eFpYNjSXWX
daHsJklghaUNtc6BfVAF1+j6kY9s6MWx7vGosX2saTQE41SyM93vTftgAa9soIniZ5hdiyoiSOyb
PB76LB5RzvfxzQCDeZvLa5EnXt3hg2lfphVPm9FR73+mQirvbE7mb1FjXQYMkt/rG1GMkUZmYFKE
q3fbImoLphMtiIQZJSSynSjDxc2G1e7+EiRVLh9hON0e59OSpqEfAkFilJ3HT2kT3Y4uiqhu0TeM
72sVrNVxT5oOJr9i7upqg+t/noH+Fdo9ipzuxFn/btKY+NigKersEgTlbuQHjy0Vu6opQ1zZQDwa
2KDD8Z/wMCfyXyCC5Ye07pOJ/zLOf28M/izHKqwaRBVpJmsTu7ADnQLxK2OTuQuwafWv6/dvrxjL
6rpurcd+2YnMhSuRc2ry2qWOma9RudbtBKoNY6BF1iTO4E6EpYFKQigHoRpWDYqro3JxKW/0SU0M
pw05o1hLxgo6i9xe7JG2+SFVs/U2LYo22Ubhn+T3ATsHOEfPORoCNY1Oep65X3eygKW8PQIa3B0s
UaVCulYPjTd0F4SSBgZ92d0MJSBQ6qldHWnSiBPkxC2XSw0rPGF6uo+Ie6HOD3P+i/7gVvMlmluz
0vxQoqBShsupE6t2Iou5M0z6f3frBptxPQ4tbTpq7+fVRchhbTEmTUG/jAVEX1C/PQDZhlz0ZNuF
qQ9K269fLkyD3sDqAmpo+NAzyDfWTqXEo6dJqHrvYY7wxj6ZbnGapTSRoG5m074401rwe7weqhuR
Lyr1TZMj/SQrjNnFZw5EbtdAOfGu2U2yFrlUcR+1mqVenggEcPyNGnWhSYl8h4pvIqm2NN3TzOor
ZHHkQeuayhgcTmCpeCc9q7yBPrsqvMs4SmSQss2K8Rr4nyTRUawNIoEOEA/j1P73PFBQgQSS6LEk
hxaPKSJ1UCgPI9BJa4I9cl8Dw8C8ADYc8pQ4MsuRbkm4O45ZWhJHfUHNnNICaC7yIHcUO+o0oXbc
3n3qOuwDNt5HzIDGNk0NPywmupIIa3/myY72isVHiaDvjlqdltg6pUtO+3YJxcyXGca407UPG3Z0
OAycMtwDTHQKbHeACQdyhKmIvfY5fkM2olQlFbUcHxBmv7Itvt/mvA58V5ljlU7YH8rFLdlxLeWZ
X7IxSmROYiklFpMlk/RnGdxUEEv4gWQDaNfE7bhbscHCDZSbe4qFlviHPzvK7PvkyXeT7Nf3ed8C
e3VkZYy7jBJe8akcaGV4Z+C/dfsMzQy133gyIoQnvvXQFU6ca6MfaZokLMd1xv9gclLmqpFEgTDp
3/ihzbX7zKJc+NMtUHfnChTgBJFHNAog5ezoHUWXtIzq6ohJruAZbFffSUzU8J4iqVBA6/DcGHP/
refOJgQ5Ahj2NrqYA+OrcETt9mB3Qko/OQXmNDA8Z4eqb3ImjnsE95f/GKSQZ55bDuD/QmpQ8c+N
fd7YJWKPR+P1s9IPRNcgIz6Mvxqy8vMEn4Lfef3E10+9EQOEVGEGOKTYFN99vLH1+xpeSwV8z/EV
kyUb8dL9Q+ThFauY7BpX9x5QrLTk2ht71aWUWFHisJks8kuY5EhNHHWr/hFWemw6eQfp8OWplHAb
s9onZOH29dcGH4fcNK47MOm9rVNnIS5FoYofKi9L0rZvuA9q7UAI3Q34TzV9yvMMvtUwUrrGHw8H
pSCcTtdl6AQ+kImF5Q5eTkA3dTu4gJtriU995jZFdO3V1byxc32WqleBp6zr8ohvXmYOgNWIoVTG
nyuw7N+YkllaGdJJcVTmQ41oSDgavGODv/ptT72npYh1xNlxTkNnXHc/33raEhkrj/DVVSly56fH
8zcCfltGxtEYUwUcpm98HNLK1AfZ+L2Lwbi5M8qXIfyJUZjBxEgYeCAOt0V2Kws5cof2Cyyc8qGh
gNRGNNDHQknLr+z0uEeyIMrp1hr/WsqV06B1G0L6tmiYcXO3jLn5pYc5jKta4b2QACd0R4LK65nt
mREj5Vg9TnAGlcr9B07ZAxZC/FpgWQuP3SoPUA5BOT53Bj21C8jt9iU4Yq/f/clKjdhOIhGa/vpf
iFhcZvC4rmLt3wgqu9awJTBidHneCrXpCkZcYmWrrZv9WcL/jJNE5YvtedCdgwMvYyX5kpan2QMJ
kN9Zl0umdBe5g9JPEcl0VdZIM1v2k61KWmBvAJb0DYNJvFPtW0vK90N7XOgsJYVyve2gCMnk+RhP
QpHtdlL1NcFmbt2UobJ1NKqXqJ5OsXVJn02RqdMyiv0bUHTY+3utAhaRgbJuNw9KjZNCHftZV5ji
i6TZs2USZtGhFTEz/7LA7R4/4cDWYwwOd08/e3+8EI7vbAJcDSic54mneJ5agbMxfxbKWEwCOErn
c8rttYJzFupFdMZMipKlroTDwcR0/JhFG4Ecw+SKYbQbgOUKbzz1JK4MUAGwSmDfR2m9UnMXxruZ
6tZ4bZ3Gigs9TvkXT2fiy5X/oGHZqp8nh3VdPdnxCsMjoWltDs+r1MD4+zFoSzLi4+9VloG6P9MT
n2QBiXKvetuXpaZoYoF1EXLKVB6ss1vCdrAzFgyqztTL830RkL8vrhx0JVh1nE9p+hbg9c7P+cIJ
DL0pjiOut1U582QeFLs68esq5poYcecbmXsuUN/kKWdcBuXr0o96eUpOqAfRdManvHzSKDWaaySl
GUiXVeG6do7nimXnUMR9/fUl05P8FTlQlY5CYs174J+GlhGl6EqiwIoumDIB3WqzagWv8GAELDO6
zQdVftBqU+vfV+gop6XdsbG1lMNEONiZhLjxOqF8LvZ3cWp0nZhqoHsUwpxhOWbYp1vtqVLiqEHf
jZnmcWQlB4KPVwZdzYgcmPNwyQs2NPjYyb71JPlXIEXJLEbsWw4uQKOMPLjqrwrp/Rqy7ZiILxqJ
Yp4HVk30nBqZLyOsSOAz/b3jaJXcxmOSv3lyS2/9LNZQIPbs88tpraaYpfZT/B1ZqT4162xg7jWk
F0NdObPJcwmZXzQEtnxK2OteGLg8oFDqM2wJ9tET/z0lkJsUQMaCzG3G+a0RshEthp/re8V09+nQ
J116ZPwkdrYP/evb14f2f5oZp3S7sJ5Q4tl11mwW1r0M/U/QUgV7aze7Y/SCPfzxYAD19QtviWnI
OgyimXrsHx2dli8xngMUHFm+Y+CEaKjnY70R5EQZzz0THhGpFMY/WlkKKiPQDg3QIg65/Xt5TeR7
mRwRQLnoFR/bn9JMw2nFqQZC9YmDlbm4XTU9GNXh9pZqQplMgXbREQUW/oYxbFadHaMksUgop/3f
uhMPFv9ScOXk5MYnO7xRy9qWpEtPPLDmmjNtKFpneSTAr+zufYuAswV5r4mqI7FXO2fxFkkL/ZKX
GzHOZaD+I4z2e+ij9a41EBJOkmFqfUhTrd8wP+85vJQ/JGFSStyByU9pxninkOdttR/mG6sRfiNt
gLM46Vz1mFZTKnhH+12URLHEtqPF+EdZrSKSTIllYGCgX5mjaQ4v0AhwhsWtJL4pdbmZfylX2HkL
kT9AwboKSHUbtJ0phAcpyYM5LXzfQebnINXu7SJDRpHgHu7FJ4uVuMqhAAUEqcMz9UOWwt178Lal
pt+9E8bAaVn5Cs5/sKs3kksSEWm8CqHVyNTzcXRBhmtSjfGWozM/hIHfpl79QqOo6dm8xvp9rdBa
O/gLr9iQp/trYRhxUa65136EEvpKhuKpqyM3BPvl9bN4GtO6MEeVaNvsvycsWu68i8iofDqrLkah
XUlnR9Gt8mmXDBnL3ga1jfoFQjfOcNYg7NZ39k6vEe5CnGS2WTnACPPywlrmoXX9vJIMS3kONfwB
5/ExJkFWhLTUt+Y+KJn75nTs0vkxorbJzb+8TfRg6FhcnzxnZvxjzKHptTipsuj3mtqAgksW373/
2XsS3TLYURiiBXfCiYQqcNwpQpwT23WSzlTqinyhMWbhHOHJwvNYTdTu3eBcc2FvfNoawaOC+tkq
CcfcEg0RdLmJ2E4LkWYfq8QXYhwcDt6D+kJ37583iG148H+w/6EQwAfXUGK1MexzK8vcCAZeMS5W
5ecXGvduJIZQ3gFxNRWyBq7wwsOEtR42qIt/QR2p7f6wnlROiMkhgnr69lGfSlr2IRbpdoOuwZtv
O8O/7PSGu3RwYfQg6ZWvx0spGl867YRzXM6yJmJEDn9lT4wdxkG7Ahqdp9CwcjNu2/p1KWdy4503
K1LqDjpVUkX6t/6BK6taS0HuXKp9N4NUcXaX+C93AC4JoJRyWnWx78QtcK592bbLGDBuPRNdMMxs
v0intT1gP4cM4P4+6eemkgjl6y268wNcUKZw0FI/gMku/XHFd55hVb36iZZsibBaMg8teAz7IyU0
sGg8y+1alJPfq1i2ZIdw/57dT8piFtUrFYcwuhaoGkUO7B5ftaaCIm4U+eD1d1+WMUHs3fIAkshf
J37fbBkoyZoo22vtuSvBylaqdL+ih8PN/8/rmfXi0XWCLQ1IS7dWWZUHPrMPhkK3s/SdlsUXrLtz
2JjUM47oLWQtS712wFPa/t7IQ2bhwjFHrhM5RswmCAj8R7EmLEIIeSoWed0gUi+4OcwJYMa5/MVQ
oDA3kZVZsqhfXSBrjdcbkx7DgA0gNUg9aS6EVzon3IaxoTFOdys+AxJTJrXyEQPwsedkIKl11I4I
SpdKcUeHZn5ZlbOuzzRi2h4+6qcYKWm6UEi39AVFY6Sm+UxbE50XTsCKPri2qdD+GHUcXbhWXV9a
16aR44/D/9RYIOeuU8Q9uRMUgBRcoEC8sN4NO9AobWfxc+iAbSCuKaAk+ZLHWFNcROzUGu4zczWL
FR/kwp4J24DmtOAGDMC4Mm8s+hCaVRjRfVmy+bNVZReN1cfgwPdDSRUVMW6GAgO2IaVQ2i5hxL4q
7UCvN9+j0wVV9lqkBiJ3Dz8ASsp6e5zcvdKct5dgPIXaMgoY9HbTfhnPlvYxgU+YeAsj3MpQHgwU
2H7OyBNnMf4tvs5kDAdE2sAr72v2yNZeI0p0fv1SidZqlcLyYXjuXjykZp+xyWoSqAf/PUaUdy8Z
GfSOd1PWwYkv5KzeMRlJVVHCLAe0vEOttbtvEV2Ed6acHmlkekrBkX/NnE0Rz6ZoTBHI/r1WupYp
lAyP6ymKSiL9vY0kTtB8Tv4gqvTrnFmmtiwx1YEpgplF4H9QBazHfAJH+7rxFThqFdsTssSW2Zr4
aeKa6i/joDMEeiXKS4fMk0wvQjLWMH8evAmEx6bR782ezj9BQr/KhLrxjLr0+Zj0VkdfEPjxLRBC
aM6irHrCokAY/mKzcY7zZZP9o58s4pYJaTCGNTvaAkVfwHTDfVCYOFNBfOvj2RHhG0jG2NLQzt6k
rkH0rsv5QyGtgM+rZggvBC+smCtRq4kGMoXKtM2iSVBggh8anJ5Lmtrl/2GAI5vWKm0PRncFon01
aWY7pBFBA0SKfXsLaQIM7Fw6j2MZIjvxVQXVLpe4mRRczaI3ecbwEZbVhxPaJtIcOxO4YzKqzjO9
4XZvy0MKLWL4jqDM/VxfQEKDG4KuSyTHHPx9vu3THvaDQ5wi7eCDZMpQNRUXca66w/kwvnQJw42Q
/IIL3AlQ8B9vnvcvvJQB/A335Vf2p/h+iJB+OU/LJO+0CremMEwSnQNALYgqUocWGntDRFD4wnRs
NjTnbU+4uayMZVeS3lhEzgZwTyFKvWZ5qLnjkmkAdg3CMiwQTKO6L42xsU+j8plsBX8YUrxYp3De
Oc/FwZWl9MMxb19A2rtSpTk0057rZ/LSFxPH4mnZOjG4SthWdLK7u1QjF6ghCod7PP4OCsCb793l
521CIMk49+460q6f74V4j+PKZjexeDec4J7+mDVHtrDvFeWrkzKBJxB0Vir/z0o6nxy9dKjPk4VA
+l1S32ndeo71d45B/l4EEKf3Bc2CyqSPSub9DE8Tpb2o7PVtjCQv/r26B81svYLLMeFNBWEJimBR
eZP+xLJm+sew9Tyg3y5qAs5uR/uEtoPvHwGQAN9sjaIHWH5/i1X8DLRCeZKCx2uFjWEREyptWMcn
pDB8CBVLF2VqeDliY+xXLHwcCMkcHp/gBUVcKGQZTV7v8UZgyd+oyeY1/i2pUZyWXJUayH2nB2Sk
2ugfOTXLC/d3cgxzcaLnUIs4lRETW7QIOfO4Wq2olCvgyRdpW/VJ9EyG7U1XTRBWAawlitVT+0cj
tUve+JcB0HRea2m9fT9pcun4HdQjoguBc6SVcPBT4I7pb8/bDKyHdmOyQgmjJfeuPUmDezvzBjtL
ilbZ35JrpaOKO8kmDU7gAF243qCoyCEBMfUCijbLOPMDaqN+viGQLmlPMz/5LlxMmhUhYyLMOrMd
k2tHhHPv1av2EB9O+t9Q1ora0++W3+UpaQsV7thV8lnDfSEjzegKTHpKij/izfMNglCK7Db+odBH
64jcIoBXxqbw10pe/9R4CS0EaqQHtx3EMzA9KjooasYCB4ZRcYLnBDEpoUdyj996dVbwubtstpob
mddBNoK6j/y/vhMOj6qvB4rfxJtflNpkR9sw0f7n3rPhvPQjsP9+BM2vhYeqX7fAPPXlTCAVRBcI
BweduLIVin2STHkSuzEmBsEdlYziwEfi+cPUYaXPuggjuB3d3lB197Rrc6ik3YSjkHPubMv9zixT
8BECw94AhdVaiF+mNELE0ArH+uvXeqP+qabIVqMCdcSh7hvi0LmZ7n7j4f9uYpkGo54RDmGbARut
Fj01gmfK3IlC8tnZXNvN83RfWICSRCgDcrtroR+kfXGZByXuXbXPIFrdOi45MA6Tt5pvg6HLkNRJ
Y5vN/xAxpxgeln/Exn+0PIzfYx+HTynGuc6V/8L1D+q8GKtWggonXy2mODMh81k/evCc4pK2HAsi
roXddK8kxtPNsHatwWgkpcJy4myt6FCExaaGTSikFY0TyFZ1wZgMARaXP+FMn7EBvT2TyTGgHrh7
zNLQAqplO/BvEsaSlQWENAG7tK7OFAS5RrI75t5BLMqw9+DhLcp/q/WRC4l2QwiLq8o9i3RwNq9a
J6zPZZYBOPtxHvVn/eoRvQG58uj8DyReO55pkOx+nzTQBv6X6mgPvE3cHp2mYDSM/EHgF/TNR6QN
UQjIDqt95pB983iQGFvzGHmIgah/Jgi5aUTrLlsDjkdWbudmkRcaVxJJr9vQsrZIHpT+WjFONZpX
qz2VvFL6VQG0NVQS+JRYC4wsKNeOreYl34vgOIaKVG9Sg5d2U7CbATATTThbW/L0iIWzpQEFEATe
vlMV++65dSFliBldvAcVXJCf4OnJ+XYWKnxkyowYSxPpOWvZhALAwolrh3y1R9AlNEggqIZqkwRi
grzmMJAJ9HwitKuDXnUCS5+PBw50BYOBySRvmeKfyssOJfEp5zA+VkOpmwEttZWwUvih+YsfH5gl
9dQoGBuzGN9KRZzd1tzxlYmNV1Ut4I0OJfYil4/mDWmjHztfR7lNgEumqZ48KROuStsJ3elmt5pr
3H6K0+VnNB70D9wiVzspyN6iFwI5z99RY7JEW0K/848mwZsErpj4SCm0u8lbwM+cysh1+H1+rCM6
5bFWWzx0lkjFC0WnndSjk7+N55COo4cGAgzlYLqVuuio82HEXou1EDzVKq4hrzVo7kAY8htjWTiK
ydZIbz9h9J6wRifIEIg1rm52MpFou3DNJ0SsYLvf88W05jkhpKwexe5wn+0hkRGGCsTKlhkKfou6
/+X1wjOHWVfAS1rnHO8jUCRhVdUYA06w7h9N3Nrs0LGKZJ3oxhiD+mnT3GxSvt7hPjMjbwFtrF9i
Ig6EV3w5hr0GvVGg6G3orRpOqFKYbbOS3NplwKXRFtJks9howpN40q3WH7Ee9GDV47H09VKltPUr
ohV9zCQyzSsbtUKNxR6nY3tTMf1h0athKtkBQX9mTdL/37cgiI9dH6+5wZHKpNk2OkF+xF07aNky
3LSzRkQ2rfj5+FOz0DgsHCQT9JwwYZrrJh1RCB9rd/zQeXsXfiSggkJkIAtmUeU3Zem9Mbl0hMCd
R32w36KEDyK+iP98teLJyXItcUHXHoyv2gKdcMGaQpejP4fvuDuZAGJ2prtjHhDk9LZMre4kMwrI
Z9K8OUSiyHPI6zVTHMlg1SeGspcyRZ6tIIkErbOwBjMnUpNNzMLuRYeDS/z7ZChLNbS/G2F8Ec4S
5nWTsRj/jC7ERwAqX7FqhK7cYphrQ5ffJQrJ/QDLeFWBe3YtBEttsPkurJkhGUsEU7fuSze9X20R
o0t+Rat2qa8VSJBmjhDHGnRNEDdmuO1YFMNMpCD8JmrJ3MmOoNNa/1Ye15FlpPmr2I4feGibCKBr
B0PyX6yO3u8TV3dYZ5s3/dDNvlBS6UV4NiZerBHVdXYeQPms6JUqiKpf33WSmnGA7GqzkrIg3AIO
Pe0QlaC2eqncLHz82P3HglGBBKaHPxj3lZeHDltWsP2lyVNtEA7igY+OtqRHwoHCE8B7TZwcUfJT
RfeGNF1BFjdanf+dyxN2PztsBJkNrwTEKra1aBkrmu9MH2ECjmc9813CcVVrLW9oigKrVq+29JO5
yWHR3Z94bqdC9OWV8/4VdecA21kSz1nZDrBP3QozdkI4QydzSrnEImb1n639Ux0W9kePKgf54ueo
J72tkyJ7JC9rCAKNnU46j/rYNCZknWXBOKvhboLM5lwjwkWFX77dOu2Q9Li8wEf1oeHO/OThKDGU
i/VyYTK8OAynmjsWX5tUciHhGmgQ8yuwCKTXQ+7sd2z2tV3GIw8g/nCnS5KhcNU/owthd7pwegib
ZK+kMgBhvYGJGLhwe+t7v3o4c3pFu1SqEixHtdfVNhq7h12WZgZ7PVQ09VWkTnkMUGi1QymwOf+W
D9YjEfHd7CiDoF42E8yOo95AOZpTpdZLNORiE+mbhfoYJ9zz0vX27+GGNCafZ9kL8ZmzfMMg2m3t
myrrXXJUtGokPoxO/ONGV1rDzQSvN5E0sOL3dueHsjJ78WCfDHa6FYoyQbJ8MBN5ujox5P97mard
/0pgr4z1NuUOiispHyZcxZrhvxdWok7TiPuOToA4mbsMBNwuyen+CiZ5NKeTA+YFgGZmJGr9Rsao
prdszciHCaHDQC0jz0Blstt9cizTsjp6nQhwC2RYB7yBzJHHhqhMpzUcUFHz8hLXJjQOtTKMRKPG
0003KNuI+m4wp4OgbvXCjSopOII0VmmPiGtqLZ0wUbawN+e767pa91ZmNOkOCR7pEMQvwX4yFd0s
C5xGhb8PtCUVtY0AyAk7rzIZ9DNoufl7YBJywZDAmTqSIXfmsE36qRyb+hLjejAF640psNqNuWLn
5kiPfqjll1XShty/sP+odQqJriCtCMeAmsl5FhXSC9kEV2+87kYWVTjX/ZC0OiKvwMEg+oSvA8St
zKcMyQ1IXR2CQLsRJ7/v8NWg++4Xwa4Ib8xnf2dngLzKkY6gFLP9vkVkrjjJuNH2ypJ+BeD7IWXk
S1K/DbBrtGmmEE45WHPPD5fg/4I3AExdA6ex9jcBjtiVLpdaVMLy6TtfVVHDkJ14dVZGX9S5HcRw
lLKXhNsM5onwpQuy/O1DZdmbsPNV5ubuJDvjdNUnH8/eTeBhmpSKGuSMpRdjNf2o6IbtnPTBp+Il
9VGncewHV7IPm5gaIZFGu933hN8XAASfeoif8Wqc7ltUi+HwNDhvZn2Zxh8rQ0kXqKFxt8V0739Y
U82mQgREIiAOIBsLvUDY87lpL1L++f1I3hSpYfEQOJxac6BxdlguWLkw+8cNYXEUSIw7KpkCOS+n
PzmHu8QUh+YVk7MpD1jc5/KlqeinRq8yNHI96UnUK/4pdAZj2pcDlTf4NvYE2rX39MSyHJwVIVb1
w7fStOmx5LIq924VTU45tpy4arNNk4o/GFDfjZ1lpMUQsygdjaBlfcVB7PX6wKV5FspHRByWqxGg
WV85BvELqG/4KqO/tiey32zvZX51tvNz81KwCuKdz1yNQ/WM4sJhzi2oVVGFGpB2aB+/EWUi6PwK
e4bD8JBxtLWyADWOeS3S9gFQ6cxAe5/gDis/npNx0Oe/JY2kn7jCthrtQU4qrp+H2/8UqDFSfxTn
cUfPk+g3v2EQ1tCtR8D0u3EGoZReMjMKwmHFf7P3T8HA/Rm+2dNF1ip8ziHiP/yD/vlIoP8IuCXl
wSV2Gw3I07JI0FMUJ9lCOZhrbvBlkKQ6dToq/8pkanUj33qzxgKM13dVDYxdOe8ti/WC42Fz8m7T
OglRr2eQrOeCuruVmyyBSnp9fU/EWSAEQca95EEK3EFcnuwdIvBTyfCrvlWQHpsgBAX1MOr1CCLE
9aloxbk2biH2Y5eD7LitieU379j2Y5k00oa50SQdqZ7qwgjfa/Zu5t4a7by0ChvJEKnblzlJ6s7v
2VEBS2EA8gb72oiT6VUrKmyIstKmbRrIc+Bviuv/r3h92dkulpca2asC3zPPgkxBo3WLmNsZkrHI
5twDEDMvthNMbGFMkC26dgheNnsGkreJC8C992Mo4kennkc5ayAvqjAcXRc+Jo+5ofGATQ45Rm0S
35I52h97stY7RljidHHTxf+JykVKbjqW0gYpf1PCGB0iuuBsiXs6HFxkJAPUhAKvturw2pqRo9Eu
kz7/Hpt5Z4eLCyrjhVp/yR/SKOUHkcEnYS4MrZXuxxHr3E0FXJL+Nw3NTKDRIfVvgriE/0NZx/72
MM5Zqft0vb1cqxxCKMPBz1q7jLZh53fGMT1nhdu1pQ3R9UZBmVSc1PLngJJgBlZGlz3bpugpf4xB
ASy9aYsn/PocX75POC03tRmfafFWOjvyYGnwbnD/SBQvwEj7ASE+/uzcgq97DUMHP79DeZDlncSa
m5O8ECNJRyoW2yWYtyLT3UwffVjZf6i4sIeUYjKr3wQGr3cIFxKJTzzjIUNg6pZcpXBmgns1VCnE
JmTA8Oe1GSAms5W/t2gb/UP4+ynRu14en0zscO3+SjLLZSYNTTL+ztwXZ5/bQQZLWG5Z02glQdH4
bPAi/EAk8LDr+aubqdza0NQJkvmgW3wvBzYTX9lCUfjz5ESyJfsKO6MCjUoZW7tfaRSa0BNScA9S
MnAv/OvkzsDkc7K404R9+X6tH17j7Qgi2+YJmR3f+E1fVkHTYeBbwY810fyBXBbyuolJMI8KlBLy
uTCAf//GMpam6PkXzRN+nvmnyPUdSPS6d70iaPaoAIzA4EcDHz2KFVS3tRAe4w5+T2p3+HEvE/z7
LgOJy9eudbRZNVOjVq841s5Eqtd09hsXXdkHo50PFv4HPMVuJ6KqxjQqL8FbttCghTZI/YTMaxkf
wEiFGyUDWLUxeZVneE0NE8Pl2ifFPisBrZypG6yrONTDRBy3sHLNHXaYfq/ca4R3UFSrdDchevaV
bvHBhd7Yts8s0bAApnRmx6he3VkwcpUU/MVbJm9k9NhNgXk4HxEYpdMrXEERCEMB20ygdoqOhi1d
qGmeaM7l9+WT7T76gZi0+jgaO1APQP/143RGRL+92o9y73LD89itUBJT9u9Om6JnZpBWh+HcJDg+
TrMDXZK9Ndzb6JCETMc2pmYBku+irfGaPliXAgo+V1n9sG0LR3CiF8Hlusde3DFQc/tI8yexBYRg
PHHGzC2/HLjoN9+Xp4ruSsPuz16TH0P1kS7dS5wUwsHjoxixBjAGWWzMV/gwyv/Q2oyU2B1K19yY
JW8aSRnTaUjUau3EzqwjtmULSB9HDC8x2BG/bo1g0VmyE60a6eMXvkpjWDGb6GM1lpxsTrYzrN5j
C0QS/ouRnzOS4wu3tvI7YnoBn6aFESZZU2tua+pwzNx4g+VyAEmalR3b/h4etIZtwKuh7vLAO0Zi
gMl0Gap+OtB0JzA6LRiUK9nU7TRWMYBVPWoIO9g2KjzveWXrKaV+IU/KAK4KF/ujhmwZNEIJ89Iq
P4UanqGwX+dbJjaUnS+4s7jjNeJTrSpRiPwHys18cuFyxZ1EVtHcZJmdnbBCmpzuCuPHPrPXkMHh
tp5oVUHu+wFiy5hi2n8+O6O4J7AXpONkwn4thjIYqQanr88gwGGqoIrWO3SBvjAPdsC/8FjA6qI8
QF7USkyfGp7FAjynVPkAhBoXy34qQnpGuOsbUzYgiS9cXg2tESuBORJGZaYorvOUNN15fPPDOVO0
/CXCN5AkBIiQsoXe+sEeV2gQYj2ydFyGUjBsD7w51s+l2+TfFovFNQnoPhfhkhMmSQz0Xl2PFKX0
m30vZMZfRAXlnWUlKGqne2hVX29C0pRYYUViPkhDU+uaxyBKx7++Zsp6/U77oJLKzOAQPCcirsNm
FOo4oQGZa+EQs+x7qZbZPTZu1G8Wyz5vGe8/T7gNWRaSXMd25N8rRio6gyY7WPjOMiyBtuGAcSfx
+YOxIKRdRuEUIrMdATQq3MyvkS+9o7mWga4saDrOmeaphjusv/2VArSvb2YB3ANJtKW+GY/cgJdV
bv/UzuGgj/sZr2zpD31lR3aw4iNIXVViO4Xe9C4ZL7DILID0kqX2lRNUDMiNrDd/679D7RuKDeB6
Jc9oltaIZq+lnp4MPiuk/2jx3hJo1xc3j1sKEnNhKCR+KXVr3TJiQ42TcqXulDgpSXdXd62IKjWj
aYH4VMJjG2Ww3AspUUk0vi6Lrlb4j8bjHoAEhCftOX2l59EfPmwJDYB9sEP26hZhh+xeqDQpB4zH
RyO7JYJMeLiQVEckRvUjkUywg/IfV62TveBscSmnoQYSiuF8So4C1JOvpYZw0YOVxTuImAYepQat
/0G0LfSwEi8pKSBNu1ZLU/rkQXG04gBeNAyaBjn+tg3o/hNiYk6bMyRl+R0APf1iRwvjqruSz3oq
R1ArZ/hoLepvJlnl+wXW8ZLfhZ6pvumXpUrmTdQfnBYbtR07KeioEXuZKQBN3aL4NcrTo9dUYpYh
Z1ti74Q3vNdfynQD7d0z0xOWSM0C50GwgBqV/if7IMUdbZjI1TWnOXbOPMIKaMcSwMeTSGhAmR6X
R2SOCPmlaUS5BpAHDyjqMc4QZMugXynKgXIcOSr4F2pGdE4H/YjOPcThvNG3ePEQds+pygcpuUW4
Ypu7PCW5UBuBBPpk0HARt80CGE7pklOXigzdjCDfYjzVNZzTcG4fCqiup4Tq090BLatXOShPvDls
nBM8vYFuaBLx9ljlhISkTXCKhDLKjCfXUJhxD8nj8ca9MeP5p8CieyEhaYFymTEQrQghT7RE4LZs
VWxzmODJMlZQ2uHF3B1qKUcwYqez1MjgWWeM/sxv6GiqoSQP2u6q6WTWwElapTC825Jh4B653Qql
KVKgzc+iYdr7WWgJh2/h+I6hxvNFsr9xHigzWtKOhn/DJQd7PxMHMMnGae1ApDPEPMUh598If7vA
0ckhB3KhKytN+Eb5usvc8HFTpIcWsLB3LXngddTR2J//QicTUpfhiKZFe2yAPqdDzxFnavgBFTSG
kMz6HCK4q6BARd3QLzHo1SLSHHhNIQM6QduIOkkPntTNeOFDhoyPdsXynaaa87y6QEYRgu4BK1ef
tiZB1DfLK0eC/DF/Ji59sYtiOS5ZfOLnbzeFYEXX081108PZ8hk/egUS3wTD9FiJ7N1LaMVOysrN
8sfT0ypfVjAFZ+c0oEhwoiNi/znvP2xGNXSI7M8paXqHIgxeZ6O+mpdDVZIJAOuC136cbEUwFA02
JLwE1Ceg4OixLhnJ41LaQsOunnbXPyjDOAvsU1anEWWh960zYBPigg+ds9lZDfMD4hwsH5hrOuqs
/5q+YdH3qFQVORkYm0dUzc4hfK7s3aEwQKnRfncLvD4O/lByYlBT7J4fIuVHvHaEO8pHWQmRHZjZ
qHOe4frdYm+onrxY1Yf5TGwbYuorOqxsYh547uWxFD/75rFyeO/84qkx81dJnsGUvJAAe6c7vqAV
2h81rWwuZj/70Ny4aAORXmMj8vh2cXHDBS7HUYkqRcnW+jwCPOmheM5oTK/B1eBzdgYrVQjvzeOd
UXaqqN1mtuP2KnFVuRGPRbGo3OSwYnr1LPIVilzRPfCo1N1andzPvFCivr0juWzBsKCvN2+JbCga
/F54amzTraak3DU4riTEoXH67xk9pUjdg83L8Ir+y3uqNQScDh745PDH8m9JlCFsLHTd8LBg0lwf
sV1BtS6WIGyZt9yh2EQZaYrr96tNmS1L3Fncvesvb4QJP8pG1+NXLlo82qiXxKw8eh6iqhWbc8Nr
5/13NtS0PndVwxR5B78pb9oJIRTi0NPMUZ43f8l1ulahcUfHr2fKik/vcCJBckkGHM0WA3Aw6nOO
uo4V3/ZsTuRDwKCcUjvD6VUNiZswQ5NoRgi3xeVIyGL+6291Iqbfjh91Pp7sxG99bKGLzS4ShPO7
4eE45RTRhqDfq7aaLR48R/foCn6cIT1s7dSHR7ncf1AT8GsYqX/7dbeIk2o9Y3G/k403RvMoFZsR
wxz9yhzHUTZZz3YVZj7Tns1BXN/5ocLe7rXeG7aOu0EfDjJ/YGCJPDKQQw+H3+ddoXqZh9ekqCsl
JD4dyMfwgQW0YvwmqLdSOIU7+xOrZ53E83jWHYhQIZyPpOpjZTcxjhM+V7Joxc870oMiyN88tLrd
gMGLN46gdew6Vcsw+zckfgIJOTTAys0pcbWASZbsreXVhK7KiiRBWmdt1nWHsc1OBACX+daM942t
N5gTFldv906B8MnOYpg+M4vNbcdlSgJ4HJUaySDpPk+LGCWxEP9Uw/H2NLI+4uqxO/Nlsen0RLk4
wJ9XHyfmn4zGQ0PmNYyPPaWNqivMKU8k1q/XKFsRNkXdfH6MYOruc1XK1VcGLveNczz4twbeMWgU
yv1d7pLs4JOPWqPZJiAP468YjeBrRt0BCnt+2jw6fWYlJIQmPJanVRkNXYeztrLKQYFAdxGVQVmN
Gaz4gMtog0BTc6vAnL1y2K4tU5Eh45GO4h73J1DslR+6Q83ckVhCu/bZmwJzH+r6i74MD+WXDmFq
kwbn4Y235r4S5DKSkfNgOQfScrGgDxTyozG5/wN70mRulyIcdsYY+ZP3rswLTJGI4ccQPCGr77Qq
7PZxIMSpUAhzwXUvxR2p/t+2RQCu0EeehNlpaM0t1Em+lIIfSNqPus16GVJ2MLs604ETJlNAAEBa
kIV/tKYEnTdUwuwpqbRY2TwGJJ9FeGExbxrOgj+EGiVaa1MH9CMywN/wKtnzy7BSGzVzpK2pRZMO
Tm45zyXcwxqB5QVPlObX8w8qtdVzsSmZw/h3WwbvrWHXjgUpWQw6eWNeh/ZYjrjb6AnLacrhjCsL
Lt6Hg/H2HRukUyu7syg5iDJVvFoj5tIrvsNXeVgeRZF9UJJA+wgyi/KYuZAfqX4LpqQ1jtfntf3W
E+06DNQL6P/UKvXm+DyOubf9J7pwX69MTU4Jal5Hri46WcVIu1FODasLCs6N7cUkz4Q65CyVx89B
1XxpDA4uoW/9tHg8DSeUUT+MwVTiCc5klfAMFL/PHyfX+vhAQMZidqNAVehs6UZa8r/azTmt8/Hu
0Kq8hkXWzVsKDjXsYNS8AzALs64KaqEDtd2f2wlJWD+MCKZUL0X7gsTsepAQf/qLxSz4CldFynyu
vwtcIakXI6RnhKIx7DztMNrVTynT7L5R1tLOHPzPSWeimUngKa7CO04OJN2OXjIy+U3ZmMTPia9L
rMRd2HMl95Dezelw7gHvlQxb+9hZ62mA6uARyPuYdLj/H9U2ojOBWVIo+aXxFUWsHmptwv6wAulk
l0cNf6kKc7ar62a+fbBWl36QEgtgaiNJXJMn0n/L1OgHCChYvMEORwrJl7zK3NpK3v8QD9uDNCN1
Hr2Nkm9gv8EaSO+sxEYkOo6bGp+dZK5cRo4QM1ycivGNqQltntR2aY2uuC8i1Pq5THbEMmzh18i8
mfh8h3zyHZ7q2qz7ueMgXRaUMRnmkjPFQESJwsatRFrwDrSqLJ5ZCxhxiDtp0c31digJu1ehFH1a
CJbxVhtXO+bYOO0py4Lz8c4ntViqNotNCKh38NoDOC4fRDhiIL04HteRE5cmq8jr9MwaN3acFvAn
iGS/KbXj3IXektmGytV0njN8Y/YP5SAxCo6pIYXfTf8LX7I8zF0NQ58eElYZyRqXG80FDOlg28Ug
2WlQXeHsJyiAiKvgcpjfSFUUUQcM9EIkk8i+bow3u/UGI80vsjeNiUneh27WzpAXI/dOJK6UQLUg
PlwlcOwGo4419iUCiGq5UMBMn2NuKGjk+6rR/3hNHu3LX+MS3jiAKMbeJhhAK9cczKxBPr+j3rOo
3WpYOl8T1B4m9JVBAj0R2QaNgMle97XCZDUcw0ntsV9xXy+/tlGvnEMBznNny8ipcZhGUrcmOPuz
ET3K4oty1jQUG+9/u+0CGKe7tG7cmj9LS19ores8ISHpaLGoJ1DWVlAeuYsyJfeMS7ODTBf84KGE
Jumhl4AGH2G4rhalj5a2J4pDHGJqQyVsKRHNnUpx3yBlsHWeGURm84EAUsba0rfmIV0FXlthYZxh
UGcJesknawTxQ/cZEKaT8LsV7HgmuI49HRUdv+Af4Ym92i08oXmAaFoHzLUeKKIaRffBg2gx7F7H
CGJD/4GZ9fMVTBVILF4IBHXVTGAMMCCieZy8oGO4yKxnfRY6i+X1lw3jNHOfAypWrzCyZTJZQ3Uz
O9FR8wl4extcqEjnQf7kWIeS3KrtM2bCVqCgklEGll83g5WXW4yzUKMYeTr4BEFHeF6UJOpKxtK5
h4fRqpwm6YHjsK2nofoik1f2EhiwncXbVcdjsgcdYr0hCKwVPJHaATqg/yilT/dVaJ4fALldtcQ+
qxZaGDZ8g58XzbmL7+I4KnqsL6/j5E3sixlnr4oiNaiZcvQYkFNKnNYVDjy/sK7X+bKZ0zi3YFCO
3ScjUspgkZlbrhNfq/s2Fu5WDHKOpl3nlRYJfzGU6Nyd84/Q0DntKbADijsW067poae6DnaFzTvt
SBVx7Ai0y2/nbdxbHo06sUKUN4ThDEzGfBSuM6pV8f887o1SflSioVjOiUF3k8HOB3Sl/D9+tnUv
Rel1eAc8hDoqou1AToIjVCStuXdgFpeNtvsNRyj0EPOhUEDC9ZuHIt6eq+3X8zh/dtnUjvsaWR5z
LRf/YVNYTWh7JtkIN4XtaWTBuqULfJIJbp3VymdHuPK++cZxuPHPJppweRgLSceRT0f6Q32sRwAK
x6itmmu8wQPYitHA3bgfEgrDuES5dfUr9UPQUzzTts28xPZTNzKB7WD3gqf28eeb+q8/KMAfbUTa
mD9FuNI02PCfZy8LtcmTwlF198F/obxM/AuIGKmkf6cTl6l95k/Lr9wm7iWngIUlA9j5SNEiAQcR
+4a9lIaIndX/pgqJJPlX1OX3WFX25eSRH3XE7Mks1Qu9ux3qiglskDbN8fIVTZeJDfiOtJWxVJ/Z
98WIn6fBjZ+AgPYhOxm2FxAqmuQ35Z9pXkizumdkFZ3Vzhk6Dq2ju7S96jVUD2zvENmGFxCQgvPP
Q/+mszk7fsYMQtZwSUbZOqg390Q/Tu/k9NzD1klApvGnPNlmshSUMPuzgPKUi93/pdu6SlUpWqxN
9HTbU1j3/qvhb2beTqr4hzVAe6DTQi+H85QUHB7yi6VkWehYQke2b8SBHzxqWaUECb9B21L6xc2M
eQX/wtNmUymOngu38hh6VOZlb+AWYwKC5mUAGgl96J0UuCRPyTcYbJxFqmDzCQArq4cIDr93//UP
/hJlBGkbIoY9HUuZQjwHT/Fuq2w/Q/E9TqgF2Ki/z1ICcNRj23+A+QFOkJeZWS/ShOs/dEs+07fu
YA5/eMTGtmpOCkl7oZEi5pc5kzouiVD5sSb4BhA6ZrpuO4ABRBGGIZ8QAEVFjaaFDdmDLtI3qMjp
JdGJtwifD5lSHjUSO4SNNi99i6Rn2tZg5acubn/uMon6Fe9d7ENp/9r/1s/HyxJBxQ96s1dsrPtS
lEVu6me5hWvJr0ykcgRCaqghM9bpWBT5S085HghJz1EaDWO0pu/1lMhuCldjfDFU881molWet+nA
j8COy1MLzJyZ42T2uoacMcMkgJzYr1Ohpc633msCf41CVhwoQajbF5XIbuIrc6AJJEBCwk++B3Th
555bfnD/OgBBT5MiXYyXPoDPIe89B3Vm5Hb/EMjU9ighEXY9Tz+GJT9glpRPfWO67+U9SjPT6MAS
5XptTB7ISh5cCsNdstkIg4oqJtMC9D33YvsqWNIMHFt6SM0A4XhmCtNvrjPAb32pnOtf7LRslEzV
Lcsa3Z197fr53lYQhuiCWNiqk1f2kKwKUgRflVhY8We9jmeLHn1ymkNojlHq94Xo3qRtzZecUtWa
e5+SbXdAfqBvOpXKcEM0LvgvR60EVwYkkAAa4+hG+4kMBgAKsYIY8I5tj6RxmwuPTNnVqrEeHbG+
xB1oDsYavvKpGLZnKBCz24p+k4UaXjeh7gjRl1ouHMNES3doemsubEUZbPXZD/L1m2PZ7rIv3HhD
jxz0Aq+viuBSHMUAzlK/QfhOWwUerG8RRqBOqsaf7wJqKrZB29oKf5VBx/nL21FeJ+Q45YqLBoSI
9M9c4RLAvZIl8ptV0+ZH81gE3xuVUKAd3xMv753kbdh2ArFmsFlG3jtO3Os6KOhrCM+kLDR8v75k
BxFWTbhZCMWSZlJnLHNd1FMa9bfeagS2PtvNKP1K7DkWTzFmAN4mfctFDopcTXhrCTbElE5B1GnW
2IWcUjV1VPLY+w8TL0XEERrMomU3hSH1xAWA2jIKuqD4MqjogRWdnrtIZG7/f9PDc6zS1hsb3e3z
YAKZA6UTQ//iQpLn4lf1NtmsfRt/h7gdHf1+0ASKiNrMBTRBr6Tn3Vy8kjzmDSjZ2JX9Nzs4bLzs
4Nn87EjKtsjFW/i/QepXn/sXKgV5lhv3ArvafVxuVwo+58msCQ5zG8RRpnOp+2cdK+RCff+dmYBA
4G7o7SwYiA/9N2gZdn/YnWK2r8msZgVRnK5oSqhlWyM6Ppf88fjIfZMQ1Uf0ceEweQGk3Je2TnPZ
IjEHtcQSv60l9uWW8ey/Sdey4SzfBObGYvMIZ4vMM1bQXUuynYTSG3taVB1cCrMiHzNtXXybr1v8
YtE5o9/rQyvd7a9OaZrN87bJz9VAVWSKAMVHEQpt/RACgV3HOjFn40KBrsCH91mPG9DxTXd9XtFx
xSXKCM5y21jQt/lgi4cVk0H3bgAXwXUuYAjVRmJ0L9jG0U2tescNjbycuKaifjuwYfHSL6/xxwYt
4V8m+GI8tHuv8TcXRrwI09lZRLwbpIK+Ynehww+ZyI/RE90TG3oDW6GlcQ5igeT3veVtb4oYp/IT
zY9+czWpNxRRS5L2DXqsELfbuGDc+CdZ8otxvkzGiUt4dWjK6v8nh8VB9eqoXXLYCwoBOHeNGhXM
O0VIrrJbgUkNtKpjjN1j25pbKH12cxZ6LkyLrsBEHuuWuvM5dhTmiRThEBkx3bYmAL40JwktaJaW
E9I3JzgWrunQtbZOeEb6wGhqKfjFYTDjT2SbuJY3g36V1G1Jv/fLirYRbPBTxgR6ar9SW0dVzMcV
uXmtYXBqjeq1ULIux3J7EH5ugI78m3o5vYK7tBG2IrsPqxDrEJQaWh+py7MDGSTd9jMXy94VVaxY
Jrp4uJvgozE51kfcUwz/S4RnzozwpR56Gc+yEKq/qD27Q+3Xkigf0I1mbgUIjArLY6o6tw55dUBW
n4IJikKd/YG5m8wvbVEUVzirgIelyf7jX5q31O1unz6N0zp0+AYCxfL5DPhC7OtVyctmnHLt7bMa
AFjmlqjpB02LBP3xUoTuwId11oQ+WzW6HDEN/k0LqTT9/0r2Z3kiQ6k74ULinyBX7azRG/YjBEU/
brUZ/5u1Vwi+wlakD4OgvwLnWA52sajHguMuI3kibL4TwIrW1vCaK4tmUQyJRvmV7kP09KRuEYIO
qr/rPpCXjGo/k/D1nfn/L13Anzgdj5Fi1jO2H9ASlZUzjq+JwQ7ToYGbLTkHAVpMeIKzphAZcqDU
aoDJJfAj2k3DO5zeFjN1wnRn7DHTPUExMdGm6f44AIF5KkXn5C02Ijme8U1Rw/5mgdhEIbypzsET
akbwt1wJZsupKPDWy5LGYS2ZB5BKL9/hEbsK592dQSpp3n3r1EkEyLRErNu/9t2hMrYjBCkz7U8P
+Xx0ERzyot5rMAE/rsftY1eROG3P1bv2rtOSLFuZQOHToq/EONOHm4uwHVWxNIRj84dIizc0+lwu
EXGIM5zykH9TQsFkOg8Zz77N6PH0T2d+zJNHZauaFBWRAs3ixOIRUUvgW7xzKaBB6jlbKbiAoNgG
ToD9PgCJmXmpsQr/5q9qNz6u6ReHDx8ZpRjIg2ZUvOuBuhWmPwQI/GUsblgGIVmEm1ekU4PNL+Vp
g72iQRIm44hq/xwHahOLcZscbnyKpADe+JhLbs7ghqkWAP69TV+r0H3tkgy0SBzaSnQNKSaRPO9L
rv7JDVbELbzqMEdmDDlIqgidVQXrdtgaAkE5fe5es9VMuQgOE7IE9soF8nCBjHhV/IbSuCnUESJ5
iRphspBKZlSP4sXGB3Z/nglUvSxPFLsE9pKr8BBgsXCPLFvf7NMPxmpIjUccloFRqwZE1HIGQ0Ro
k4AzSC52gZ/M6PjIzxPOjTLWHRT/1OYLvpLNqu5z0m90sSenhwFOMwKZatXDZSJubLqNxTIDJStQ
viQvpN2OsMrbPxJtrDfCjwCPCT7a8q4OGMv8FeQ/USk1CqhjlsDJWZKkS+5RyfWQtottddLM0jTe
fk6CS/6kekEwbIqK55RJSadjs4oc3+qr43m4R8ojWrCeawRVIUCX9WocNG5JEsXbeNTrln+MMxaO
vrYYfAoFcdejH+FLvm9vsqKVsgrhmyzh60CHa9rnYK9SmBbg/pnQZHni1s6T79rZ/KO19N4AdnoU
VllYuFk8uuGDAZdW1tA8FbMjhl7TX2Lj27uqQ7l2iDbecX9ZA0g6e8MYqZbWk8KBZIU8vethwuky
rHTc56dk8h7fldlZOjjBRatRLC6NXkRuyHeb7FSMf+HRAL58ouHH0w2AhTSrenlRlMS5rG7Nu+c6
1JzT3K9aAi31imKwcmuP3Fv6XUVXBqSuIuBK1tnQzkhzc9OaX27NDz5suimOEyTOalmwgMWMitp6
Yyg1KtKF3i7yF7tmy0pYYZMLtzyVeI7T2/nYW0R6FOD9QJ8Juv4l3IntGguBFs/zCpCcI0kxwSNh
Wy6nHUXF85xvRj83TB5gMHQCmdjpad5ve9J7wTukzjtsiTs5h/FaVIcCQ2NHdna6mCWJmwrweDPJ
rsk7/NgvGumV7dwiL492lqIn/unAlTrScwigTnIWErHniAq068vf7qybmDYvBvhTAaBssKmL1gQA
64fpBsh1y5WJ2lTocFRy/DVvohlX9sTGklc3fRadAhQu5Td8R82MgiMYcCvZO6NJqyY7G+xGpbF2
2cQ47gA5Soy2JBQbmM0Z9ZCTGz5j3LFTN4r90qaIAjVCouCWxpilwwRRYnQ1ncG5aQ/SQ8bZvcEK
h1YWp+e03uHtf8UD5i2oCIuQBNnZ7PNK/opw+t3GRp7CSGVP2MY0F9gAB7WktI5Sj/gdgQbXN+Wf
698zqZIsgNj5PRb8J42I+61sWNkGFW2QkyCOf4sQpgxzO4nvE6FUDHIpdTmbXEJaA/4war5eZdGd
j3mUIfjmMzOQrlkTY4ro1svESjG+RmTdPjGXlusH2v2J2W9KU3kvfnCaUT81I93fqRRM4h6zzfp4
cDhSy4XtW99jt2Fw2H98cQ0pfFDo6qN8kPEvyvkQq1E/sscup82wLv25aJHi+KeBwA1Z7ijlZrth
FhUYHB/GMBiNMCLYqYxmlCK2Wcu8m9I1ZP5Gvb0jJJayp87syKUMVqWL+Dcrdxf5zimcwA+cbVy3
dsvT2ddbsBKiVFSLNxEvNM0NdzNr+iujqft6Sw792iruVavZPIWvLtK/Vw840CXuC1UKd/q0vje2
C/sfBGDY8Jir9AJtDGjkFDToqjfaDUSrQGdbDkLephqJfrJuoydh1bkUCRh06I1DgymXNTV3bo5+
owMSSyjzTzDR7u+mM8WIA01Zz0ESPJrzcHu9kTbJv2mLetU+9I8PfSkLpZ5dAuOkorCAcefxFMTo
ZREi/wCM/7E9RRwXqexgYWb1HSIJh005aSVuJdaceJzOKhcREil2gEozzpip1DASNe/MM7MeaLQn
NjxvtOJ3s0uThNIaNyc7cC1OnagoKL7fvU4nUvfF3HlCPru4Ow6t6cLm1wSoHmOAuWIm9T1IwrEq
wzKFkp9oY2sGIh5yWMIX9wEbQDkMQ7igOAVhaGcVrWr0/oyhuCk46g6aCt7gV8MvhhEwkOUxCmDK
BgTIPxNXEu49TNM0S1r0Mox9oTwJk1SVNsIfZnuQVHnkCCSMONxmf7YjJC+cPecg9qoaQGypCiRH
JFcnqsiGLjX6YM+TNBhRWrpprfD14tfdyXPxrLn9INsCH+PDpiTNgIup+Qm/jxGnCvJcZHS1ngM3
K6JOJFhl3UchlNgki8DkYBr8SVkpaSKNcYN61nc5WiFE7HYvcO2a39c8ADpuuLghw91hudyDtDM9
A1+DVQs/uF95cXz2Oe9VJoxQBpA3rG9UWIZpnbFOnr+Xe9Q9I7P3M2SSFsE1epN/SGyRzLNyXGaB
UxkPgsNgaHTCWCC8dVoNmMDOUClPoXn79rEiWvRMTCSfBgyvOH3VcOWCZlk1CJADSudOFp2Gk+JR
XHPc8sIN6s82miQaRz6F+XvXoHB6aO4nEwv77p92/C6/OFIckCipM51YYKiOq7IaH3U798j7kWrm
qt/BGRxYAoCh14qXhu9+GlK7qOvrpA4FUt1ZmXndkzvnAx1Uk0vCD9796ATKOU+BuWd7GWKFRO9p
WDS0xkZf0+Zfm8mvQvRp4cZLJJwidINYzNu7GjlcGKrl83JBcMqPn4d2YnpOrvULSaLqeMXvQiHC
PjzxVsFEBn89ShKscwKZdYnS25au6HImkPbr1uMuhTltGQBeG/Ry9FsLhXRjl6gitHujhS0yng41
Rup/hVsAxlajjgP4YRUoQsFXCxCAhXgytDBuJmvWdrYZFp88tZB86TEhNv9y4ao/S4PkkiFZ1daO
n16U2mYmXSj2PPI0LyPVnt8bDafOa3QioUBI0+IIRlDSh+8qHr7J4g4OMWHW4ptAnAFPf/7VOFbA
m9m/xL6mDuJiaiYmWWxglhvLcXhLHcb1v+6hcFhg7vyQiLAWO6Wo2CWc4fRv7Wuc4DPCnCCheMzn
vAypDkyuv6kH1g4blVyxolQIqp5aq3cVPX4iLoaaJhdzOFnyfTtZ08r0n4/DOt/ZaFoUl2OqcFH2
iDSkG/D9ctK0dCC+LBxrXkGNdVXDiHDlDrN9O1dIjTFEWWMwaDTqnVC8eGjDcCppC1JMG+BFrHd9
haIrFq4QBuH9Hu2qVAGGVIolBrTaLvh7dWikqvHjJ7E8w/jASp6b0a5i9cyVlbrBus04HTGsJoN4
rmVlBAGKXA/OeCElZSy9D6r2AMPcpxTFHbXqKfl8AwxXoWYqAWd18/rAGOyPt7eRAhKoz2gqiN3B
qBQDkQy4lT88y4hGTJqDlldvEGpBzWjJ/mcEQkAdP1L4aWkD+Ith1JHdBLn3YwgWq95E2q1CuoXD
N2Soj4oJXje1dffK3m0hyQKLoOLUhTUK9ZQdUF0DKxHVSx8E350c8f2EwGx5x2xGBDg4eS8GAot3
umRpPjzHxvVkPPJ2Ha5vxZMoUQDWX8ixhZMPsGkk26lLbD6QHnm9DAL0fBuxmzVJB3QFsJx5YgvW
pYvkulXqMoZkm0Hx9OBpYzJelsRE79eQEQYHtgiFvXX788qMNbY0bY+Xz49mcPKz8xpWVg5dEKXl
gqN7xsqukGcVZhpHNr9+JFV17CsRm7g/jJ1W4WTZQ8v4KJuf8GQSnkOt0NPpt1sYX/nDC28M7RWC
o9VqYzYn1Wm8KxeD8il3nDpwO/lc6R8P/RpZUFPa/kkjwBFj93tDkcLRKGQ6KjdzpzhUiI6yJYdo
ekUopj0wWrY/5qL7xBxoKGdvjmBj0EICFD7uIZCg2m/UrqLx0zYzcsuowHAm7b1cdbYbOY7DhSbA
Q2iXIY5CHF/Doepq+75eDVuy0fSFF/MWvXNyAnx+4PCg9fkIlOpYXkS77m6HIsAjYHr+gk9oL3ez
bqdDDDbMOJkzMmLMWyvAswRKLIJs3zchJctxopS6MatOvkV/TvtVOEodxRgER7cqeuqkaufv9wNu
csSnsBtzKLqI25uFe9CM7/mm1jGgL0Fs0QlyTvIKcmFd9eaC3A9qMK+pu9X5/l9n359SAIBQ6T7R
YxX4hS+btMuhCURJQaY7RnRai/Ovle3YGZNHqLKB7hQIq+IzNoW6xai+C1RE1wXa/XBYi+U8VTNn
U8SFqNvH8M+fHx/PeFKdON0kvmkUVb7a0mlnYhfKsygYWQxgkgamU0kGlRmmBsUiACvAXQfsVOcF
Swi1TmMmBLhgRpx3b8U9KUMEP6uLfxJGP7SWWm3Gu28FulsRRIsRP8NhrgcrCcJZK69y4lFNbeCP
ulA0W1KqaLI/PMByqWy9AG4wEDvGPOiCr1pXZIBUZzvWEElqKm1NFnFtfF9fyEmz9rblHsOQz6eO
xm8GVJ295ldLNOJ8KFuxkFWOlAvdTbHDG7mBEX5uaJ0gTJGoHlr0N7mXb1UTwmmx62xbAWNJ2a1P
wWhVovh42afXrrMgbqtrWcowDkTpaTyshN/B5eVfCgSE2jQPhNV+jzMQHZJtAoyXiIJ6vQuIoT6Q
/9+z/xIfvw7AUxfE+aMCB5Gg2C9Tlwfk2SHWZ0W9Eyn9P7WKRKSfbeymyRYDF+fbeAfJrhfK/6pa
bZEygY/oL47jrBz9E19GR5MNbqQOx/a3mELmNO0BrMx4NG598rE9fzYjFT5bkXjiM8E4kEW7LBM7
LfdfnMRP5Ps3gKcP5J8sVJUboQaUPOPXCmXdbAXrRSSDEIbOCZNUH3lkizuXsHa6kWflntjjWs4o
zN9rcoNLN5Qx+3xwqP2cRx9YkG4aYSyad/iFETBFP6nlrwBRIyNnIr+JCiepr3wVWF1kkQH++9Bq
YXva3puv0OuyziqqqiuayJeFS+/twQ8L5ip3epdmsaCLMKPFEaAaUxM6NI94ccpzFx0NflMtzUc6
GTKkm62vVQKlGZ/VNYxThWeLDKrl7NlKGdD9ugKqWsi22JaHFNd+PquY4WC1xjM9uRYlfXI9rzab
WWZyu5N/Mn7pGEv2M0bC7ZGwxwmYbb/SzFo7fTUfg/phicjOHWyZKNg47RyuGJL4KaI8FyPXlqi3
HWKIG2Vx+hruh6n8jRR3xDaB0xEh8xbeIuUZglzb3el7lUPC9POq7JbDsNVL468H1PSyOvHWdTpY
qELUjQHF1jPv2bijaM/WOHl0NNY6gnFpDq3rb6Q/DVCWd6fYBJzRMW1AZWLt1B2jlIljOOjq6gbb
4SYl65RL6hAaql/PpPyhCHth5V93RkJAX4yyS76t6qNkbRP0Ci1NSYmo2oosRcpM6Tr03bEzXoW0
oZNuuZxvWhztChXhpyhSQVAvaHgZ8IKK0N7IoZAQXQ+XTM+9N4gB5rIyLa84N05WKFMCcqsyFZm/
sgEViPYaQ/Uw9gofRV7bgiGuDYZuOGqXI8agBqbeUBxZB9wy8RfUTHJ7127SWiwB9A3kGVGpqimT
tAPhO0uHwXP/+YGqlJLpPxt0L7lobUsyoAyXWEa60ekgVHL04THDJxNAkVI364261+9Djd/bXw0D
HISdZzPsUZXHiuWheW6AIR3BaDSJLLT/C+LGifpvWMrq+XpLmJt7/gjLE8P2HHdwFL3HVvA7HrB6
SgXM4PlRFxrJrBDs5vcP47wAad5J4RnIhyjl+dyyV/DJ3TpWn4zTL27vBps8wuyDpI3UPZWjriQ2
WFLHx38Ggj9LnCxVr5Nxn7GWqxNrmsJIblKKRh/wYCkTfWx0JK/bz7iFx4JaA3kv2NPh3YfmxS/m
Qy/oO2/MwFBj2ZTTZmjoDbmmd4CON6+/usb0CmfkDz0TzNSS4cZzWdfE8LELmeN3NRf7Li8TrEtZ
ekC/dtIDbTKC4j9Mt4AzWuBFkyYAAAJMMtTwvNmRlmw7WtF0iA4nielClpD61XXQa0nKODIwptQ0
0hFW23jclC6aOoOuh5d8NfT78INHmqzYqovjiDFFDBIeZzf42W5dmNxWGmyy452oY+gGRjmaTtj0
3LnNw+23QRCfqMwnK0WWf+u6IGNui0jjjhuVHDGltrbYG/vOUgCDEFcXAFZQXuhk1FFRuh0dNGn9
n95pYi4NgWxlQlw4QLCVYTQFBYq/OKpQeMjplMKtIWqYHUOSgxo7cxSuObRzgrxwoT7147c9rDzY
g8aqpcJWxrgTSzU8wxXLjHLjdh6DrcPQ8hUsaZ1zNvZ7N4Nbmpi/3MUJ6N1Kbqzpx7Yt/8dyM6F1
lp6sF2KAf/oEbR/ewr0yogfQ6suGuqPzDWRfX5Lt1b6WIEzcxtoHL09M7mwCR7lkMuurxzVNwjX5
eDF0uNV5mV5ccM0JRnSZMUAKEwUowjR6EFuQs5iu1FLWwF8XEcPfVz3KygYJCS9bvlvtSnemiHRo
UscRpdXDEL4SpgU43RSNXlKcfM7vd/XtbohBQhAvwgZeZmXPKfwiNU+D4hM/BEIpGeYBaLQsmzRC
MsJkvRJwv6EjIinypUbcye2wBJwjGLhY0NHNHZyUp2gYTgqgAOc6fNJhcs7QDPNVpgJzkxz8ioZZ
fYULOlvEyPrLRuGPi6EMVNFos5yhWaApos7kmNNrmyLSDwnKqMo/toqz7H6S97v5F9td39yC+UyT
Cpu8cs8tCOgVYeLtV157kbK1kKTs+4kmxV7BufVHvUmvoB54BHEnTBF3s6CC6Lrcp/WmpF5O7544
UISVISmvUCHZ46qkQDo4kZB1X0MNTgvxpPG0NRKilY4kmDccslJyPP8xWfX3+G8b8JqrRHoqJ+uH
LEu7O/8EQgXuxRAF4aq/UmS8B1EVKJ4C9ykvJ80MxhvQdosutMVZgp7ztgAW/ov9d2pY4Q/Dbuob
mzb10YlbjvA/+JesUF7zNNiewXZheNksfsaYodRvLpwZkVWccfcf9XhshABXy/zSSi7t9hVWYmIl
zXQg3JsXpN1HHIPoiaI2K1pfB8tUL5Sv6deGK+JOC3HaVJL+nUySdmaQfn65+NNRbLPAjTo87uqd
XQE+Fxoc74WdK2L4DbWHfweoCsqgeEm86bLWCzGCNMKuPKFWMcaNzfPgRCB3wEEJQ6+Apikkiw4t
/RyjjgSaOxtZgiOp3TSAWKi4k1oIoPFo1vzGKGOoQfbE6gosNPqBzy3Y4vvekrzFeuoia1Lxi0jN
GLHcvg9l0N3iRZlCqqmE1em5drVunoqbE44HEXM9RwguZ6JVqSx0Faj0ZEMdkqGOrWCfkZ/REmrM
TEC/qvjcQPgK1K0hHg6wg14ywzqXr0W7MpSsgMJmNdEuil19uy+FHtcu6PajlIvLLZhCnQ3lM3KW
u/mYp3o33yHEzzIPgkkxKZJpg8FHM024m5FTuQasWbv2AWayiZBU4YzHhzs4RtXsHXQ6kosuBaHT
8zOfdfawsrIa7M66r05/TJXdaCnXiQsW06aXug9wVTylPenJEFhQjo2++wNG6UpL/oQrrWkCASQD
m9WFSUVoNIGWc6WZfdjz13aO7xxuDOqaSpIhbdLiA12mYHkVnuAHoMKA9v0tjqO7qt+Kx8raQwKO
WHcT/h78AFAP24i+UxRPEhUNOMT5An9OjGLBa33N6p2DEaNBVB76uNd+V77WWwTn2s5LuxrDsdoe
tUop3Q8SMe8q/HXhoAWO6Ho9o+hpzdV/RDID4APofxVvjjrHs/+vATtTPRUxXa2JyDND1QBnXP6Y
pGYq5XZUBoi/kJ5uDFHcgDrgnHFVwM8sJJ3W5OCru4g4KvtHNUVOfUGYbywLIE/PDEelSuPZCDI3
6+Y3Rjz+Ri6k9KyUaIPzKKwrk7CDYjca4iQlbTFrXrRh1HapCGlz27GiWfCPetAALrbUVzrjROJx
TnaZB9b8ED39WFgahDHmLp1snYLbmrZrUFF4lrJVCpVezoJMdXTT0xNTijNpa1sAltZWuhLPF4JQ
WwggDkOuClrO2zNc5DYI/ChNjRXsLbPcj5ugWNrmIqgJOaGcpsRyLmYaqe2weBivkG5K2K6E+dCw
OaA6/SGeZAc4QloenxPRCfSIxFth/lkfFMkiepMfMqV3c2luz/tS1hgaHz9F32/FPkYbuegGUAgl
QEfpw9qEh2cD2OE5K+ETs3C6PMx7pLNs3NsSjuJiwsZVkPCipEwS+jZf+7t6Q1gcAHjCc7JHoQU5
9MXpYS4d+MEUXEQsJUeabbuUr03tVg5jkrP/XSC9WIzcGWdasA8V2/RkXDu8nS0KgH5fZGWt2tOL
loJ9AGx5wC7/7IG+tH5ECqhDf5X4V0W9XimN1XJxjaRyEEgesbSSKOJePRCCJy8OfLhZC3pe4b+/
BhVAUxirX8bTgqcElG2+vZVWx7elY+T5hUX0BK9oZLAavbBDoYs6YLamymMAt/ZQZw5wFfKRORKe
oSyoOVxanRhnhltkSO1petAenfpusKsNhXZlGo+brL2JVQTkUMGoys9VXXmTNeEk4/B/FLXz3Fwc
vA4htKF2b/LADlTs71qQQdYcbvn5u10wiC9QA40z4HFlHNR6P7QR4jwUpfgJ7qs0viIo8DtCfmBC
QDxb7dbBf0LjRu+9ZEyfWbN3izGw2EV2zJLzsLY5IR6eQmnbi6TQoiFBDQSH9LQBTNVv6JfY1m8+
9XeWpyeZObFd2fJxhvm4XXMXDciHLknMGHHHvpOc/7nRvn7Snb78uFBIar7oFeYUbersLBNRDDt5
dgFAcvBA7rui78EnvLFaFZJPAWZfgL1WutU8xkvwpyy1LZfJiPqLiKIRO7cD+XLQPcdfofjY72of
x2pYi8cKth40ZLzOtEN3MPKaFHpGqecg0pnDkm73Q0sgOVEcQJkRHXhLBfmIg4QEJ3MEY+JJ5ouh
N5oq3e3e7dv+Prdjxp12c25mPMH8QivZp57EOg2F9qgguJxgKT74j5mP18yV8TMCA40Fx6xkHrox
FvQuVnsh1a8+FsxEAtAhwtHle/eG3dlq5Tp1aeL9lkekPtfbDMAeosnYrqWmbzZ/AeVk6xbxRGhz
XvWp2BpI7uWJBgXJLONGsSZVm7B5MKQooBoIPSdtFm/FkOIIyI7C2QqYzl7IFo+wPDbx4eRctUYu
ilq0CR5s8ahyG6C2YXpVU4zwHxu7DKUlTkgq7HwXH3o38dms0f7/BWq0QsCGQ5HSAWhl9NTtt0DK
Qok1Pd8tNDooqOCkTjFNW6KAqi15zbOHnqzjwmCdpwlvOTk2HWAqKfa7Hi0zMEL5g01blDkutzKA
l3o1hhFOVS6TkBrBK9lHPPbKhzMwN6EJ6L0b+Rkw8KE/cEz7s4/TPhWq0yWckcG+NsobDXXBUWbG
ZKoK0v91MlAuS1EZ2QmuFdsKI8qblvoiH5qzjTRlmTtrEVMHWosKHOpdyQIv9sheVj5SPBQ9QLFc
PwZ88ZAW5NTUuvXO9kKuTsxnPGLO8vN0HX6xL9AVJCTbVqAam95clM1tq96l0DaFTrXQMjtzy4nj
CVU1Y08RoS1/Wtv3sVBxIoINDXZhBWFZLqV7M4Fg3cGQbE20dzXjenjZA5XVsW/tY8EkB27kV9en
V/ltuBr8lu2CHJplX42zdz/COw+iUo1nmA8BdBEn/GzBErrFB74EhTlNoxnIQCvkXSWiPzXdyn6r
DWIRHvabMA8JcFvQOckV+HKID0rzIy8E85kjvDa6iKF9tiqKGUJsCQASfECdA7O08AmatgA/Zkix
EWpKe4ecoiC97hjbJydMTvv9aMj5ae+Br1ilba97cJlzdUR8QSsIZN1LRH1yC66nyQANMi9CR2gk
kLO8aF2B5r4hTZuU5C1XsXlSfMxWpCdZpZHxeqYe/pwePtcoob6MT55mbg6awV8z1m6/0/U6kjoP
SiPjDWcLcbrgod9J9qm24P90CO2nPjqPGfA/oi6kpPvfgFr5FjOYs6HsBchWsVnh4rypHrbGfICa
pSou3LQOsPBEY8Z8k1efo/K7qSn3EDMPPLWn5kknYRmaJAkwxr8gH34v31MJfDo5COw1F5UrbixW
xQ2wmhC65UBkB5XBYv5YtOd4Jl++cc45kGushOGRi61pV8JCUVsQYPFfOVhiu6I5+KVbOfDmZ1eX
XTm6ZYFMDCscJNIonm1Mx5Fz3g6f1DEVFmqtMewMQn6wnT8+ltbuTh3VaZEiY+RJL7zySmAmxHOi
UDotzE4iwreq5RQX8k+mp216xdy8m+qcAMwZc2iThQqKoGxtE8t2uzGl+oStzLwieyAwIovqXq60
GBLg1MPrwomVgoefXy0La6aWDc10J2XBeBiGGG3UkdkvcOx4r0fiX+RGxLTr4omyVftsd/H3zbTp
JWzPzMjfepmwPGnqU3pPe6wLLF7/i/7elzxgu1b6GFGVvI17cCZqVOi9kH+/1JS4zRa59NHJuxMw
YiM5RkLfvymTmvFtcN9sj4GZVKoyAlseucPSwSKxFUg8z+9O6VgNslnx5AZh5+1R8zt+pulhqh/X
a4hAq2Pyar7PfwTCfJcYp42df0Iu38NN1mvpWomUr2uxHK0Z784G4ReqrK05sWIPRElJvJtYox1l
0/cOuUXT9Up1AC+Yrz+/IsVIRz0OrjFTiwFpO/qYPk250nZImntfVf8CPzYAa+BbZ1UeKs7ndK4c
KQFGAuzO8I24x/FmjPbl/h91nG1w4MJbaxwt4Hqaj+gGYibnk24BG8xuyyQbMMuR0MMAO2h01n8q
xiB9rzPk/rUxpQNEzYZTAPKcqqsbLMlJJqdQuqBxtoY5nsJD5OAF391PNweYW/0L6WpHJU0hQGqd
OnMAa8IByUtSVTdEl0dUG7kJmIjkk1RGOlPieYKtNZZ5UWWB3dUHRyxainOfsfMcH66zuzFrZVs0
Tkz6uO4b1lBkXblvAfbHYgvP8CTj+6EQdGc3RF/lMCeBxai8Tz2ITp4Y6/HPn7eDKi5AYeflLSlS
pF3SR75TBI7I8NsMf4UPqQDII8cwsRCY+Id1E+rgL8h4nekfnrc8Hjk6RoaNCXEPYIvxTtIz3xZu
oHoaao+nlhb8lwcSFPths4djS1BFqTrmLzXx3KEhavB/ST2mSy94ZgY7zpHO4zk5gbSceqYwDGHB
2cnk0Yc8NJCzxjabS1OIxfb2vk+R5LM0U04JMoy5+3LcsY/l88ceXgVFa7pQJ873GWKsWGO4hfTr
bSMu5CgT9Ly+tDTBSP2vkIw2CZ/EisvBAGvFsJ60oQgbb/dPNAvZYig9jc9rHiJTHo8tbeBrvTwB
ZQ7cyHDpcGv45/3dW1jE+0KcNPOaathxpRSmd1D9SW9eJlYXiZrp/8w+yX5W3if/VOBu+8ECNoL2
nrPWYqaSsWFfx83MnQ3Mrj7WHx5ELgp5aeX/jX8TkAY2sDZozQdUF/yRqhqqg8aPLLivnm/GVlet
lPbcPg76BewMQKY1LTHW3CmvCERRsWJ7LeCzZKe1TNST/XYkNBkxodfuAZE3Ihj8armrvgS2pAH5
3Ojfa82WbTBKfnLzOPxth3HTLRXbXOdDjhsOKdKJaFoBD81QncpJ3ULw7NdIuI4iJBF9n1WX6xe+
nrmzBF9C2ayuTUWqwjzPxxk5wPx1oLDTmNDa6ZstBS8lcXLFO+dlukb9tp9RhKmtsUoulgu3irzo
RWfbvEuLxebfHSozmnmPIh6v/AGuZipCqyFhFL3EXLN0OqoyDSVQO9otTSI5gAhbcKsZuJX6UCxt
B5h2TAhWt7egtJnh6Ns45/KTLeoxMZRCdtihQY9AF893iOc8UskAIBE0YV3ITNfo8cAg4XIc6o0a
YbWOssW64HCbfpjJxV308tOAqZ3lzjORM9yra8jl1PVgFQbeW6q625OpQMzj/cu7HRSurORBVgEa
dck4yeGkQNPYitWhvqged3Mq4DqmBp3SHLnPZ4t3jz3Tmqw4xMyVnx4aSLxoNyFMOHmz2BJTSElY
kUC17sN+T5VtU1FIbZsF3OxPvkl+EwjGYIGSnSbmVr8M1DEHjwgU+ymJYoqpTPGPgrkf3EPU7D7V
YKs0ZPHshp0f21Dwogmtt94ILyzaioE3meUz/kEdjc1Gk33VrLYTr3fvC0fsZehF4KHbMFZqjW0m
CB5Fi5xT89xWcAuH97XLmjUACY2qWer9A38UFmWBLd6s9YOUQoEkPFeiUYCGzOYcdk4VSudNOP0t
EOGIiasXLzgvkFGmnwOcRpCwDE2h/BVstwhTljmx511xcwacTtENVLsWMzjlJaHt5jR1hfI/Ntpu
Hii0t2A5Ff8ujDJgGgiXrxKNybrI3Ycvci6JFTCqxEQikYHW0h5R2OlpAQTKHE0ULE8ZyULKcczd
gMtyJ6aPhVVWaunGeX5/vY24a4SxUtiRtOkuVlBm07ogDF/L2P7rXR20UvVEiqGJSPu5qS5sqLn5
WocdXFT3bSFhVXzL7rFwqt/cRf6jogaSxZS98OySLTJG8Rjjp9g8fU+cMU0XEBaKufvUccOdVwR3
3D5aC3cQ01zzzyOD1rAp946jdWD3BIyGqjmPmRAUs9beNG7egW6c6Zh2AdqhS66n/evBy0vaWu6n
P1SyuznTRuevIlderqv6i3MkGiBVaSaIXETVeG7fBGK56P9AEj847dN+ZfZIiAYnU8ANpmXgErjT
NCilAF89ubcnlJzx3mYZsamTwNhgFBnDd5rqU996oWYDYMUIfyN4ZAiPuV5mf2ikC/owMIjJ9/p/
kEwZ5Oz7nQsW4mOfyzPioy/JmEKCCZH2xiFa3bz/Bilr3TwZdrO6EGRrHXQZdlJpFaQb3WIx8f4i
xcI+2bre/FsWQcU8Z5y9JdwSOECvPKu1jWmVfSzXCEqIVNFxpYFHKSzEw3AyOLn3NNwCdhXUksI4
CzATgowN51Bkvwh1U/n6iyYLDE6HDOy87TcvijgHjY52MMuiNotTKm4gUbfUWKzan/U3FYIPVrXO
mxcxfr3tgoi0HhlWC+YKCB8Kldnx85HQr5OONi9tl+tK2WoTlB6sBasO7LeG+AaZ9tKtmJv/ZCZG
MPbcvfHCUEel6xdRiqn/NKbm8xBSOXOLUJtC41THQNMVIKRPaUxMyL/ZN3CauWIzR7Z0HbMaVG8p
lmmGoA/8ByE2m9eyTL4/8FLgj1beAq91gN3x4M1+HRW8v9A0fbDndJ0y2qmEohEdob/3AJCfoDl+
OsCTxO51oa+OZ3FRCebu7Ie9HhJcWK5jJ68j8PhBJ+1LLnudZ5Se4usnPFKOcceJpG+UaWmAehxf
zopnZVDXcfPSZcQWMhtClvCnXrVLNZx22wS1VPUlv+2Ro4Dg0IPrQCBnVkyLIApoD1tPQlAzxyo8
/evhdcWlJREEeDxxpAhDhbsQcRJzKN9cBpRNfPE2mOIdyHTPD9yPV/vV48+cDPPhdmumtLHfWFgz
cbLQN8/97Gy+yQbzAo0JjsSDWfjQaMPpijDn9F4kVDxs95PnQrRzLdmdYphaKUUCMkMojouDOiTM
YTZauPwrYUrMMveJVnayZZoyrpz8Jmpqzc/oM00jzZCkKrllxPyWzl0tTw+KCu9ErHSRAt9zcRpa
dhQnFqKmZq4X5TpSkF3HuxSJjVN47sZiCKUegLEchadJPY1VyXevpfEtlVymRAhJLI+NyiiNIu/G
LR8yryjLhsVDQ64SUYlIJ83qPeLGYu99UnwNavnvTSx53OSFWQllL2v+hu8I9eybk+G1Y5gsouMT
htgX8ls1jqhVur7AvWZSzPYBZDXdHJVrKEHvULe7hKlRPhYuCxd237XIYS0yL6JMpLZHpWJXPL47
4rFP0/NFBnFt1ZKEFRpHyplj/slyLDbRloGCbrA6iYP6VmsSA2pU5VpT+XEEkvFS1SdNq2JsVIe8
QzbYjJlXWq2+VtLKy6cwVRv7yg4dkh9/Vqthlm7Tt4yB+RyUkrhuzE/1TUAmgeUcTDuCSnmm1D0E
xXUy8eYpxAXIQM9EiQILZ6A8cB/32lIaeXEmainfo8J2ZnMuLnV6x1vsJt6ep/zdEaeaTI5wGN+e
q862lirAjXBEuVXAVKVSzZiXyYP6K0qDcj2KwJiI3XWSd7c3qdjnpzHyHDrDIWGVY6Rqg55kKNbS
iL0RNXMHIvrEKO4dbTGOHZh68GAA4P0hZhIku5k42LQJNK95yYYb6s0AmxgpE5Xxngc7KusrzIoH
lS7Zb8LnUSZsInTV3ofpSTC3gedHWtTkcKRsqKnEU0SPnD5OF2O8Ok45RjyhqiQWqUU35jjWHpgh
KyAD9MKKBT5Q2m01B981t9dZj6Gd+nQ4BtU1p50RQD2ExsPJRiwa7NE1A+t6j+q+mMi56yxv6SNa
loVfD9SvvMCW+khnrhcLe7RjXbU9e0MEYtRrsEUGKeZogx1Z+F/9Lz4ynFSI20eKO45+YJqWj+1M
vABsHv6PAHJfK3u2sXVEY7NE9Ko8RID7Ov4rLUuCe0P06WjHzDhsV0tl3OAfQ4qLgv1/mY5ZNPqx
eAZfj/wk1K4+GaIAApGPcSbl3RZg7M9UHSxWu3qar8JDQ5Ym9uWmM4hKAvSIHV8yyRmRwQiLjx3V
of3VeITA6VM0CshGYpbrx8POHllTlSs+1vHTczOzITOrkZ14gbL6PfRkaqAKeO/1rg+1xQp8WzlG
2TFflde+jobSya7lqrMU1EzXsvsf/d5PofA7vxy2j2Q93PJMOTDSzxUtrSLvzdlSoxs3Zdt9rSI3
myoWBnUVA3dFaj9KVHoPXhwWrJ0aw6dSzoJDqbQuV1qIcQqIV3zmEWz1GqAHmYvv5dxwN0v9Yeby
z8wTHUYDtnvQMPKUvAACUJHtd55CN7QiNmjThh1WUdiL2sJUS/57Lxi3upzGsX9NNHDDvSKPfH0p
TjCgF0sbntWpAtFSAfJK7Lvm5ykjHwuaw+lAuyN1kWUZfU9kvASRKivb9HOWu/OcK+IZFLTaLKky
YwulkC151PsNa327hvr86vpgaUSo3BKTOIU8gFTnjfP4LwVLCX1AtbYOIc8mqZfovyFYCqO5XhLo
1yYiI9BS15YBj8v7GYY5f2AuAoO2jkeYnnAkkDWa53e1TZehnY5bx7Ymzb9wVtbnX52s12C5H1Fx
u1BdL2H14csCDq3Yw0npthpqU7AdlRU2T+OvzIUY4pRKd4i2wxz+jt+z+Zt2HkgZdaUaXMiRmYmu
WuE94JsT44uxTecLUdF2OHb9T0c1pcXm1om0V+mpnZWomwzVazjFOuBXMtqNHwyPP+0zh3FdoWgi
xdZmB2vidIxjw5x4et2eW2u5nCUuRuJz1i7i+994y+7JTAQCDaxyuoFi3wua6Y5xMG0DXCKRtenT
lwz/RuS4I+H3tj8uEVCExKfC3O0v97h0z49r5PxflazI3lIiqqn70xhe1DicqcYJ7c89EvH2/ml+
Tl1F/rS4GcwyiR1QC9KRnO08f4LnOo/dZOY6WtUb9QBnb8xeVvHRam61293qih86c59TVi2D2qEo
sxgznmmPf+p0NtYSAxhqAKGGy0Ho6HoyYzZrSWtDgFJ2jnGaZ92Pd9Tk3qYg0QLvBqe8z92beV1L
PIpE9ZbfzzqRLcDYqjZ1lPyYPxiJfKVt2pITLlUttKVfMewFmvPiZRpgFxm7HcfZA/eRRYgSAfQ/
Garmvft2CIqX0GR4dB8VcCAGn8BUzIxUJyDzyet5YRZVSmjQ1rOKnz2Pw17c2gBE8/7p1xhkrlI5
a5qlAVD5FSk1QVv0NTTObqluyajLy4tJxWMxsoq91JmrYUwBgPNc5JaEAZ6R6X9O2kXOu509GuUS
G2CNkJfSnN3jdKbF4dKY2DyMFVb554Nvj5TCrZqsNkbvQ+cK6oXNrD9NA8U7LaJUx6s0Mg6WGLS6
kj9YeRLY+CQrQC9JMXZd1xlDb8+Ys4tCRI0dtVecZlULcgW0PUiSQXxoVgyZex44G1aoOPrzc4qz
OlPWPeoxw9uiadidiR9L4SMxTNb11ORZRpzGD3+Cx5Jzl4O1hjFpM8SjF0j5nLwZvNMzxEkTVpo5
liDMJ5LocB3hB33ap0ZaprJxFXPQibVrO4W7vleyHsPZyFs2fv8G6Yk37SDL6aSQEesvuVIA6jgY
jr0sOn/ceEUROim0etvOAAafuVDGAn4FPlAljCdRTTgL4dNNb81eY2bMBO8lP95RvPedCB7Il8kz
d+BV2EvC6zY+4a+F5Pjq9BOH/oEybpwoyCz5dUGFfCe7XflaarSFLm8cY+Z5c2SUVDHl7tzKHWnJ
Ay/sLFpwTjgpigZQqtSesUQQVlu3y7wt3+frDv9vmplzrnq1UDo+DYmU34jl53YVbqYzpxbuyz//
LzrD8qPsSZCcX41x6pnsqddOg1gbMivCZI9rnhSRlsTQ0XvIjmMWMR12HRqFKwM7uTZwBPtm1VJA
TbB5oLXlHpM0PCssKwZMo0LdF6m8TDs8okwoOVxoV9/+oUDDG9FkuXgkWwhSDutXx0jEQAjdDAGF
zsmuqVTwoSuLug+vddJr9tpG2GowX87CUfg4ISyzfLYro691Hxu9sC+F/kt5WPTfIa0sP98WMVrD
cME8m4RppD6Zjxt1u0qhW0Un74SIndRVUbQX3H7latn6Lk5VJVdJeG8urZT2nlxa8hKRJ1Da15hJ
7g92WeGYrAAUWkcZnz+NdNerYrIDci5ZqjfT3j9qPWz95vFBym1fYnIgCKG5PAmqKB427C7AsgM3
42oUmvwSfpE6XjP330KnFQi8tuvS2iVYntXOd1HvoYZXUxy6cnu60sZLqI1x4rc/CUBMJrHI4t9j
GWgwk2HgZkiwvPNOSc2od9ifg+/EyxHgSvf27WtwLCyIPLCOrNS6SwvmrLlfJSMOtEcKOdT4T0gB
7AxDWeSXJ/8K+gvLyaWcVKDebUZE6y/L6hO3rtB4dpEly2+QwQ51Zf56e/7iDhcecdKrPztq2Pe+
Z+2MdVDfRdemz292rpPv+ilTIambJmXY3URZ7BM+StNB1e5T4FQrPewZcXJ5ZmHWQ6nkgw33XK9r
x9rtK43sk7FSZRIs2PSFt8O32K8c2DJ16JbONvCfb8dGS/pFSYr61OewUKm66ZbJfQ2757OecEM+
13a376UPxet+k1lrTCFnO8yy0WG5sJxY0iwUu4Q1twLTgDZEswWfy69zSMw95e6s18R3bpPrDWlG
Ptuill4dNmNZ3ltGWiPHD/Ekmh/tDkrA+DFOtinx4wO9irpcDL2lHEbXhBmrcSM1d0IRt3ydZmvJ
YKHPBgiUB40a1yFpxuBIcFckUyumklwkVO4ftYw+mdMB0ky4ITNv0QVAqqeI6Fb6jmZL8YE22NYc
IwdKLN8DJWq/fAbRhyjBUI8xX+rUXF9KfFXkjJANa8ydSjeYExLAakBnza5VLDXYytREs8ztb1tH
J7n55N2ypFaL1WG+mfEfamsDMZoBwnU9pXKm8WRZrpU4/UqDsuFO7stXu542YeXYm773dbeSJjLS
h8pdGaCrorlUsMjeY+91618k21/Unq0RYMcm4rd426N1GRU0TpIrp/RKGoPOaALCkUcTxjyzhKT7
EznMjpSWgTn1YVoJnJVALXXtUrIdssuBuutvYBC7ZoWnrRdeH4lBuJekROqNtyY404OOfwVmqx7c
tfwx4U5QlVewrGFt078SbfBn+YELN/Vt1iENSg4xPFmUOMGI3nL3wvBafqWZ5DABlQnaVJDOfSlq
x63fASmU6YWmJOp2SYzLdAQR77phweMakSS0QIK5xpXLr0PAAn3kEEmOtK/z/r5O14GWzQmT3OEm
VdhsKJjLsv13Ps7mprpwkVrU5RbBS54MNPNZvVNWr2bx0u0VUL4MHI2o5GjebdfG8hFeXiojC3Y8
0FcwLm6VP4cz4NbU4H2H1Gr5zy1qV/XX4JWIHPaiEFq+xOAD4VCtjwVwYo+fNHjzEuundzsKXAic
aWpzGtUdONdRTJCOqy53nw8DTqTZkz72++rs8HNxQG6o9bOs95vgntTzY7AQFgpu7DE9wbybeRhL
IHUY4I8nQCOLLJWmhCXi2TMqUlLgMfpFacguQGImMONs7lqM+zDtC/mEGh76qMFnKxsayzaNXgGp
iW0l0qe6Ae6AXNkLIsT9WsyR5UBJGjUKEBa+/rRrEDeRevgcDbYFQQY6B9pJZttZfzYTx1g17B2Q
/xftCdAfWPKraasj2JABMtL2dHEXL0DjAZf15kY1mFCw5SEiLSjwPx7Ptk9NjsMhrR8si51dEIoy
i/5rvKHHHTl+22heXGF5NdaksAmWXkzr5jyPNjEV8BXouXftg70rRGH827u3c3s9yK7UwbwEAaBH
pU7JYuq2BJGGLrrWW61zdqa8YcEDIfiuhLRGoqLP6YijNBQiSU9mYib+CfvcB2UxCGpg/nrfxSsp
qBSZDi9IdepgXuDU4Bw6k+vrAySWAWKbZqSdDWVsUyFYvOLiKRPVaP96jzMuDfUGHvHHna+Y/8uZ
i1vXRuf0LtyWo81lrcZxufUDzblJovL5lcTAFrP1FJaoOEi/6r3vC84kXHjnw7NN33YDupA7ycKL
zqOk5p6bcAyPAtseT8bqy2yxywqRKiTO6TUqgz8+sYy79Us+18uYm51Xie3VNqJCAeJPwgdfB+kl
EVEvFr75PCIRPsu9UQ7C5UYuw/bprU10TgaLkfHZwa5kNG5BIjjweibK4njGw8hHAUvBS+OI0il5
Rc1ZgW6ZEz4iaac/HDaXA95LhPWdb/JBSwBvRpWmJntpxkWny5cv/TX8Vk1XvavmzZEMnJXYO5wo
kuKd7k8hQvuZiRY2ajbTEoEnvNqv/Ryu81GOSCUM/T9Mscy3Sd152xU9zgziFurR9HT3zzWWWhHm
qs6Xi8UqaZhu2x0O3KEgxHS0OHXJQ0LewNhtnaWLTZV3JHkSJ6HjrwZMKiMXLZaZeklBHR19crHa
mHthhpjWyHzdYwg9IUWMxAGruqHiU7LMiYNi84+1aXV/nvuAy03QlrKRHdi2TUej4b4m/XZJschd
ye4D7b7tRyjAFVVH5/R0J8lt3wQaaI0vhkozSAXR4+0EJ/ND7agsMdjUv+aYCGN+I8M9pogp2EIc
mqDQ0SDIH3/OgxfIIiyXlLKg7OVchagPQTxD8Tct9+v4x77LoYL5V9chZ7vh6xC7i9Gip5swgQtB
CE66ImMnS/BWQBYp/J+yVxLd2qevwzWzMT5vMpkdCf+2WBOowkZy2ZFHtPjYpgL9tTzUVmf16nem
GYN/Uddk5yyGqfPo36m8gqo3kQR+W0O+ilK0falSoPmFXIAPOuQN9xu5q44T/WLKMU0PaZ8tE1Nt
hldW3gJedySWIU585yKK/xfbhb2DfY/xJ0Dt1V2xwo+IqEPQbj9aO/5iL5/XqrDW/xtgNoUBpWkd
Q1wpEKfh5dkomUm0XidW4TmmVRWm6hndIjvC5pszzDT1rBTC12K2Lq4dxRqHHTe8uJnIkh7UZFvK
+NTn5XTCsNQsNUb4crCu5UwyobPZvje2yJCBWRW1mPlHOrJ8/9aesqQkjl8LeQ8TAozVgllEmLGC
3RowT8qYqdTOPjei3gKlCoWpLQB8ml/ylBNYRYAGtngOsnflx6Fuo1ShqE2Q6mf18GnrjlnQjJJb
M/EAvhei6sP+n1KGvQKLO8pyoDoT7MEpcJEHipBQ2tJFHBoiW7lzw0zY7V8ZEz9AfDNYzFP67gGS
L1wiujGc2FYQ6gMeyUpJAInrvo8ZQF7mqspiB5HDxMDhxG7HoPzEAEyvWG4JL8r65owcK9LfEmrA
H0LZjQJTDFBrpvc6Ox5QzYjD8J9Eo0Rh+RYeoJTNEcpn5UmFD1Qxs0g0xhDWYKJUWtwwPzuqetgh
Px+xLzxLMxqgN/fX1To4xs/FHtBbjX7Lb/Hpg1m1nFjTurxHZh9iKAr+/HXelWqOw6hXE0fwgtUt
S7T5Nckr2rAvpvsQ62zV6VQ47ssQaOpFHD4Tev9FDvJXe2UALYoj6sDNmeke3xy90NVps6nAvZVN
Ku0r0z5fUhJjK4pCA9gNrxqBRMQMcKRKnxbvb7tNu/kJh1934JqNyiZExP0Vk3uSjLJcGGNKSyp8
U1MZUINF0TEdE3qLXZZa7h/BoLmM3eVP+PEHNolM5T5CtSCj/Etu/RQnqq23LMUKiLbRIWKz+/NL
uEzt6iatwB/KMR23tJFUYOrOWvrC2hiJ4TjiAS9DiDjQ8PLasNWtbZuUFSVfAMONofOAiDDZm9cB
QTVrPVag2mQvO9KmcgW32UdzOFqWcLnFtcn0eeiL3WEHXXCs8dBFE0+/KgIWFxOQvHfoIDPTw1j8
4itheCxTxHdL2kn6TCgfCfSZrViW9Y0s9BvY0D79j3igC20e4q6xgl1JTvWVW8Sq/y0kPEcLmkOH
mMm0zJ3M+c6+cPbSI6z/NuCaW6BuKR4zVsQOVpnoj3T7Yba/sqnzHuiXgt4KwBwbGSwyh2q8S3XS
VA6cVXRNJ8T9RD9WzvQ2Y61lM8aWVdfwC8RkoysiArjshKudK8dBaV33ozZXNFK+6W1hMbjPq5hI
9yeJx0dOJ8vvzvGyTwH0iov31KDPYiDEySRV4WN43gugvqeiWV7LFugvR7kWIaXVW2KxDBMhgEgn
Xe2zrwZ2uLJ7HGg9QGYEgBt8zWoPXvR5B1ms+lEC/FzP/I9uhubaV+NM6FPuxSVmDLPgnAhd5y4v
WkkAQ10U+YCIndodQyzHJ78NZj1YIJWor+fiydBeBBKX5eF5R6GKU0D+qSTZcaZeKB8SwN35bAIR
JH356iKIj5jGe+s4+3z+V58yO6QY7rVxk2GU9jW+Pklwsb9FNx9qThmb8/869dpkfrYaKzyuAQ6a
kg/8xlav0w9j48z0+Q2bbc546qQJiXKYitor+8eG7dKyRPHXRIrINqdGvhlMBFsx+LQNCEioEO/D
9pf4/b1G8Stfi0voxoRWkPhJJiRODrRQCwSINPnXmnxWCaIEMeEIV70AdZe1zIPrWERd35WIYzkz
GAM1ljkyQ7mGHF6hxeald3/gWFKssMYXYd6EN13oigQYtc4bJrgg0ynmoTbKJ3tBwgmAWNmI4KsD
pnv5x3OYc17aoYsvxENGawK9+Duoc1qPHGFHgCTsqjZHstAI7NS43R1vtPqtd0OMEJBXaY+PlL65
T8BBW1lBCTjhxQh9Fd75zGdLxdj3uHrCY3iDcjViRn8LcD+9cMXsT3NRKYyM2K8ZRGrKeK+dLkcM
12Z38PlVuVGResr4jx5WVS1UNysrviw1+GcnlIc69MnqHCqXg/iOtR1d0QffpZ3O+DWiUBym4AYQ
UVG/2/RNASrHvbFgOvVJYU8EdZ4bibY3eTNmizY/jN8mT9Fr+/8hVc62iYNHgaCDDDhAm5elEXR2
MO/FUz2lbFy8bCaR5Kecgg/mUobwr07vmXbVv2iS3MEL7KZZPw+twJAabI4HgREWM0zxQKDEZoAN
SwtzopyXcyjHxTFsFVOVUvxuQKTES56I4aOuCY9BDn9ZlM7b1IyJ/nkLf3Tf6qSs5Yhdl7ZeGury
EjRY5s2a5akN5IQJfc4j7v4zd1ake0AI6zfGSu8hmTCLHpFzR2zd0v82vL0lZnwEofZTvZY85Imh
iVXD3dNpWWLHZc93HXZI1nfGKmmbwmHSnlFsSYe15Yq/n3zyRHWq+ZzC6317oAeMahoq5z1oj4O7
+yXWZIN5hsmIXFsdZLegBLGSyYhJdtgbiAelm5JsXA4FTUC7XcwEmQwpV8Fdz7aXM/tyrqn2MoSF
ADmjGeDRGp5GE5/Iixp1M2TMSS7GXTpB898QmJpclTjduOEm+Sqjx2JxCuKsvffsnfle1R47fQap
24QNyH65jWQT/HjUgH0yZIv1look20lr8ScSaU+8s1r+5wAzIApq/39OieSvIm2NgNg7AyD1KP4F
WOp2ixpNIurWA/GSeMoSm+ujHML4cSDHvVHt/pUurPyMhdfK363HlXLo4BqbeXpio0C6E6i3FadY
gC1oFEH4/w/SkhHQ0hbExoL8DmlnUQe6P4GkOkXVtQFkzRKK4sVBCVO0ex8vVcAIXM9n69MH+2tN
yp5RF/T7AY8q1dEgjNoAoncpWwM4PJk4AmatWOSD4fvQMKQT1QGpeBBUf+WQxP7+nlOMZaCG9++F
l2TGFgOA8s88nb1TR6N+r4PkUrlWvfmFnZPOOWDrf2/F2sHgoP0lZnpAj+X0HRgkmEyYI/8vTF5T
jUbE8pJGwhh6XuDLa4jcxPwqqQYBocUdMGLXVXZ3deQxTQbfBHKgvkm5oJtA9LzadBeQxyRJuPMF
40nUT+P34EkO6AXpIVLlNOpkxZeUHaPwxWRgwCWtGwiIqBdp32pji7WUg4/xrn2t9SVC3Q38omWd
3tSwDZ8zvB6OhSlnFk9WcJ0W/vuYu4yDDhjH0ALc9hTPz3B/kvez6JUe9D7FYZNi+BTzmwPDURL2
PrgX2On4/FsWAzZFJw7RjN4nDzz05pqqOcOehlP0rNIh0Bw8y3Lth6AcDzLEALvq26raeo/v8kh0
NkLENaqFcWQYvOCcg9qVaqrLNv0LdedsQnMyEiKqeJGAVvy4hoiJpLhN++GpNAdaBb+F4wltH1Fs
+vyWmRbIyV8KTrBxvHX5YZr1AdsGQpBLEHxHr8TPQ/wOJPeMap9koahplofDDQ4e7nkOMWvqNArE
gA0GJJdjSq2Z3KdlVDRpZF4xc17xpGxyy/YmqJ5pweu26WuIGZvigUFOVg9PDpkMARcJCRhGEdmb
Xl8QrCwq9l9C1FFhzrfmLdbAwikJtoO7EB77vWw5ulROohplZEPkTUR79Xq/KyVuX50NBLUp0+fb
59D7VmrNXOYeggNOhJh9Ld4CMjEH+Bj4/AuaO/+nJLIM8eBIOS83KV12yVjd2CQR42AzZ5Rd5i42
lb6rcXux9LDC03QAC+6LFYOLP/NGirqinjJ+8C6zwPhk2WzACK0euXFVQPu7XrgqdR7FBrAvNAX0
gfe8NqmxkTZnZB2yiaJWevy76j9+RTPQF35d722SxBCBK9rXLkPtlXgkg3XqMx4NdLG2KRew/FOf
6yBlAZoa7t/aa3pYAgqC9x/IvCCRDmlLoQPTTOHv1J4H4zlCqQiTxLU62BzmLN+B/2ekrNwu3Jm1
spRVIGj/2sIev0QtB7qk57QpubF64UTnKmyYKQG3Q17TS0xGFZh0MAtt+V+t005KHQ7wyfM+fkK9
r/+LeHPxSe4z+mWa6JW3UoPGpIAakyqDgSKAZ02aaZDhg3ekFf6TznIjvRKoMfzqLrOwInOZCxLP
4nijAa+jx8MhddbMKPQLQaDYOxI3snRkGYdjDaNyphS89VSFXxxno5YlUeI4LSGCM2rEltIMn4GA
0egUCwV3w5gC5DkqW7a5EBQPKm0kzVZu4gpUsl0GHaKuqrgHHH6yUJ/GkzDT9FeTotYwGhf/lfpj
2qTXsERcAnP4EQMyrtXqZAT9Tk5k5zQcbk8XRyH5N7U3HTbstQ3RslZiN0XLX76m9nJ/NG7h3o5m
lT+QSks3yoTTt0l0HH3rCbjJItZ3wYPKAJV5jCqiieJTTgydKvTsVTz8fUC3eMQdZGgPJCS2Y0HY
VhTvv8YV7danS7/Pn1S+BbI6Ap7zRRHen6KRRU0tTb5OIZomujh6Uxm9MGWXncgPdZmM3Mcxgal5
Q8s1m53CXLui6m9n2UTusmmcHKLA9fM0cwcPMN04l9yn6LM7vvMI8t0jhfUbrUVhV3ug+/tW8k4I
P7dMrs8SkV3/CRm/6C1CQzcbCFL5cZ4uGTQQW7vkB51/4JbmlWDy8gwyRAfQhE5RPwp6Aei7jnyc
v2FYbqHidGocIRHP+2ryaFIMv2yAExh3DHvhzDORXF5kEAuX3FOqjWmnsPxBGq4SQIfS0sAgJbm/
eJqrpgOHkJlV3ifMPyLAgNB+3MiuqZe+2BIPN5N1hTeDmbgilwXgMPSv6Qq2rj3iDTT2o3oYxnTD
gH5a0yMKfPEkCAaPubYLaOVwSv+tXpxK4Fc3o+bWD/R8KJ7ofnjF4DeOwArueNcs6iWDr1Dg272k
LIG+QDrtgh/UwsS1APeOVKoZibVqEhJtj8DiCavZFqFdC1RqSnvjjzbxVH6AqFHKpfVQVjgAAfai
bGZfZJawR6lvCl6+LD1oISwEE6YxBbSkYLj+IqJ9iWfiSIU04kH251+hqMjp2iPrVAc1qwnK5Yf9
LFfhrVd6ixC2ks0aUPYnem3tzMThDF3mK6iWJjBnf0LiOp04onkZuaCey5Ry36nVLltiGL4dhZVE
zbuGpSQgkVqngFZ9Ri1+LfD1Xnjq8JvJUVayuagCQqfduY7VKQ5D3sNRG/3bJPhCdC1Jh8a2qPdM
mdtJt09Gas3uuUk3M0llaXB652YV/H7vZXyaWPuFKYiRl8Jyo9UfbEAR/SdQhnevI3HOFnlCx3tH
x6yNHggKzgM+AnvGqna5Cpc4sjY7yA1wwfsSZ1f3//y+nmeHqnqC22fbn19bcwAmL9IW8aIxr9jp
5m55UBbZPd9aLWm3cBMc8pPYKn1RcIjS1tC1xMbMm+/KF9zRZdFZqQeLbmy+dNwHXoo/rYdF+4T6
MPB6dvkgbXLj9wSOnqKrH1h4d+euoFlDooYQidNDkS0pGvDDi4Y+EaGFvXUNtiPSdczAO8OEuPOL
ihQ1ZbwCteqcc37jxBkMvfAM0af7lR4zPEhVXB7PRctKAUZyldwQMVsAnwLeMB0SE8cIEe3YsrsZ
6/1eCKTRwqZLhY9L43Pq/lAQYBA4NTJXyejq+/qzHNP6320MZ0EeXBAW3hDwhc3BsKUTaxdBlUGW
J9OpyS5miUaDTEQY5LVnXeDTmRoO5ahH40LHhZJXbW4BzyTKaKzf2fqFjsWCiFo08LsqggkW7pd4
m3bi7UpUL2yMYE4Qr+5TV+D/0XTnYI6iPIKLD0W6TWhf6av6+JK+HIiUlqBswol4S9y6avvyHxCh
jZLcV38ePWuWw/jdZHMwuZudJV9w/+T60mYl3dFTaHTTeJnpQmwFLctoQWpjbtHFspaZcnZaDRRa
8D3F6/s4ZOYl75QORRfb7Pzz+Pr6gAdU0EVQNGsRVh/Mit96L4o8RGMG61D2+FNukvv+22ti5QOf
SRoVa56LRDi6JItLbs0OiMqlp2lPUa27OSDuFEOwW3fO3Ndgwu5XytWe0jfY5sogSMc0vxrRcH9q
E1A4C3rffYqhuoeklr4kQSUinU8wMKMrhjjeAq7EVH2ORQW14SD7l/o6I/vbXnwwovXb7tgAAWtz
X3V6MIfwgumouj+3FkR2/om94/Vd7dcrTqaeP2N2YELzAV/LJKMz0Ngd98ODhE8N/eKpJIk8W1bs
NuW0+8YH9SFvanIEDRm9RzKkFdfluKPvyaJjStxjbjqQfV0yQyPjs4k2mFgePsSz94+Gnsf0M1G2
gtm6Npy6QamUAaJ9UQSj9KfubjEgwen4x3fcq+9vcpG2COjTPLkl2ZhZP6fV/Lfgwk9Q7KJECG/6
hhfCHJCJhI1nGxugsGweLoz/0vaNsDu+16A1tMgjeV2BZBFmh/LnquMzb+EYMlXQaNGe6LlZG8jY
yOmuEvT2KaRs/RTqp3yLK7wPOC+IpD0IDMwZDbbQIrFcZD6A0kke4Zms7izyK11OAMPXhYHrIYhv
SLgwS5PpB8k0veeElSAEFWx1wqofJ7V2TKQJclDWWUuUJ3fRz72VQlpTrCkc50yIJQ9uc78FWyfr
qq01FFyR+gFUnUpk2OUaAI61qJkkgUrJzMmllxHKutkw8ydzxbXwZeeyeNkG5vz9OaPZJ8Buwq49
rVs/mKDgXUYQbQQLZyV1WTO4Wlty5Yycf3a4Kr/5SXw3HNe29d1g/+jZHLjMZzvWWA3i9002OoVd
PV2ZmarG6ucoux/8rffwUGHOXvqxV9QvK+KhNbpwseRSm/oWceyN6+CMOUSVJeVY1KqcALmgjZSo
7QZtU9/cu7CSDkL8YhDNQO99bw4pakqmKdRAc4rzXxkT6GHnIPL8/+oGgNh8mMQfnoCLjtwMYIQD
Dl+T5ksAHu+JBI/Jn36fYB5dDkpu3LXAf2+v1rzuXSweAEbtfoPj4VVskAv/bvgNF4VLb52c4nmd
Sk3qgP7nv8ag+37FSDIGd2Ibxk9tlj4WMy5GRGaR/8n9r+L6GkqAndg8yA5AYwaZXwYHKHlMcLbp
93JQUEFPKmONGzEA+4oH2pEWwXrprDoSGvr5FZ4V8w/5Hc+L2nyHOoK1j/Qj+UlcDG0kc6LAU6N1
kNojI8df1O+AilZGoQC533ab34qUjoYTEdGMMjOc5yg+fVJlbJYLdzcnm0d4NUUjDjjRZPPuHYsw
MRGg3DmkyQ+K9y6XTuNIxNVFTLcOwB+U3vEYaQ6B+se8//yzCsdqfcxu+MsGxeNQBbXo6vU+09JQ
KueOPI081AHghAcvEVJbS7aUA8twUycTtw01iInazsnab6LJ+KmpdLBvhDSbpp0pMQu8Gi38Lpbi
sAaljypQqth6X7IYH6rXkUKlQ8q+Aw1fsjVofPARVcWb+1N9xEGPgP/5L0FIH3McgZXj7xbT7/42
kigBApUllFg/zxYUBnezpNTiIqsMuZlKxKRwmTJ065oF0hq1eY9RchEAGSUBsxTGxYQe8w0gBuDQ
tOZ4ZtqG/mHj2T6SJGd9t49xA5HPdIzoa+zYZtn4T/OyAclYuow2gAb74ZKQgTCBXM3jRx8ehWaq
SpppkLnSq0BYAP1Y+8YxOZNPZu3qCnSUJde3GIg3250r/41R6eOnvZPmxz1Q9j/9sHvSxRysyPOp
RShN41Ft/SfpJY8cDF18xciokqVaTa7+EQ3/4ahyvM5bfpswmzQ6kB6O64FPTMc7kdKN1VkLKOS3
jtjw/MsK0wjs1aAIUtFxvtTi087RDHEAe7OkSf8nhe9mts1V2gNjig+/DWXljHWsF5c7Av9Y3Yp8
7KtEu7VKYIW2ZLUQiPx0Inyaq6DQoevNy9JnQAPrkAlCeLyi1iGXuRHSZSU57p6pOGLOrQf/zl1S
WFNgOCwRp1kktpavAE8FluJ4sKbxgg81FVKgd4ASU80V+C/MPvm/uNqConUzIG5pUL67EhkhpoOO
WHfTQmDagLic6t8Z9cuydtE0CUel64TpFHI96v2jxppGMHbDtrJK0sx9vc86qwfym53WobW/sqTG
BNroIur7A9JumBZX9edriEaLi4KJfyIzLqNxa6EtJWjzySbn6K+btDP0II9NJktqL0TDfhkKX+fm
8Bb6AtLNs356x8KoELCfgOw3V5o5HtaP4LpBOQDqxmJIraQcAvA80Yw0quEeiWDEhcVadc2d0gTa
JaPZJmVmsNOGynafQfTudJsODibTxJsd6/dTiMt77q0pC/c4bVvIm8rHf9hR2XxG/R1XybbJbNBi
noVQ8QYE+n9vna4Horn1CJNgapiz6IFMJh/1ws+X+hr7z3htyn12PSAZ7YW7iLJpCv8KpbR3xob3
vT/zpGSv0/du2it/Mkk7wdyMdBsOD6hP570qo7PQAF8hKLiatrQHsFLLLiXuUZyEkuMtvfL/nf+P
ubGAVcIDxXlTxD3271l1X2poMMlfvcpyE0VG5e+9Ae7dqyLU/CiKmY5Uz2YUClux6qyoaZ8cgsZH
EMSw8Owy27ddz1rPPG11z9yz9sDh1iML3sAkDQuKCAdx283BjK0lsY8FouDZufaD6FRS415HghRg
vP2H+0PMqeKJPwvk5qNcz6E8DPGXRuuGPoXgGCsyqWzejjvTiqjIHZ+wB6NQYFLMjtE3b/Bbm9G3
uNYaJICM2HDLmRpxWpZazRSDGSX/sRfgZ++CuSj6xg7l+W5XHCyj0dHOQ022K4SqD2TiWIDHTXpH
AHxNb4O5VDhik1+ij8Yh+wBwVPphI0aYZGEnHM5GzJSmsn3zQFY7Xb8EKi1TNLlFuvPafXDaYoHc
Jbc7PcOveCkEdAECmWUNyzrZRGzW/fLMhkPy2wovhDGI+ZVK/c7/7WSMmxlqa8Yc4rt2oCJdkBeY
OMXMvm2oIRaN1aKhh2HUnfoRITrnVEDErmOzUduwBguYKfUWtlSQNfZ4Qvbj3bp2azKP7B6D8Kta
mb7HCrZPoZKBn0E5EAWNf6ArA/4v6IWnrtEDXP55Ic5LfSaJJVLdzwSqwISOR5uY6QXy80V5NE8e
CJg2SowaAIp5YJjnbPaEsC4NZyOgzE2WcFIHTfNRfInFbEwF1Oke93c3gvSLT5YAjlyKm6mdkjX4
/gbeyqR9maZo71XHAY8EjQwTKu/tk0F3kWskpiKgXrp83tse4hvu7jUX2xnMx1ot5TI71ap3Xk5E
Foa3a4xHo8H+CGbf2o2LglPUfzdaI7xfQdEcYcSxZNoTnPw0CUq4ixEG4PHcesjSYNDQsJjhTfwU
ejMkBL5JA3ecBTppnwWW33afh89vjxWQyC1ABRWzoDOnIQTH92UV9nhrQb9Sg0r+6+dd+bsQf9dZ
XMse0dmESc2k8PEz1dBvW6NCG/AznHZ0k4aFgmyWTYesImODVD0DKIOKyVkF82pwdfWStzwQST/C
v/MpRli9TgjShHs5z2nvnnTYvWAhFiVKOQm/nTDd4aIz9pZxqsReJK/9JYXmxTWhkkec2hZBFoIc
3jSKX4VW3A9JppGxbdQ9XS+5c2Zy4Kw2ZjPrVtlm4kisluTp9aUrpgRZaaRXxAOkDehL9daUl0gi
LR/Oi7z8k8Fxd4xQgQ4voEjOqu1ZbyKhfQklvNSywT65Pho89jYOkQRaTpQXC/UoVzCGGElMg8eQ
bjm+gQeG4aZOdGPxOTdrV8wVkzH03WoXksD6MX++Lc2Ff/RASiboyEfd5QWFbAUVc+T+p90xpxPq
XEAfcYicxrPNpytKIIKmFhhECRuaUjyNYr8WzTJa8V1/ZoQuG/KQzjwc19M+0F3CL/gDdAtJgHiS
LbjuL8gsB1q+VIDFa40zUJU4pmTIEHDMDZS5aKC1O/T6bQOAKQEjwEe29hetPlzsbaGtVvWf6zlX
Sm+9q89GM1h5WlCkn5fPfHLvezeSbA9bht2zS6yQJAcTjfTYAHrDzSAXhckktEBd5F6VDk2efFsR
ld3KYvApdiUyP8eIIODsOTP9FdyHJdkWDHhMG+sLXva4Ac3ppsudZuyNp4c6pyi5yeJAJIw4MOOR
Ba7BttogiW68ApuKd2IkKCpeJ9cycIeZYNw1pOftsmG+hufqQQWjJmUrN9R+vL+9ySmYj+eVrKXn
8/H+X26Le0g1KziyXpC6+yihAtyIdYDpsCoD/6TC/VNbtHfahTdMz9TmgBdOG7p/EiycL8JowTKx
rFAabT3LNbk74TPWTFijL6aaUTlgKSq9CxlfMVbNcitcJQA/gWEkEpar9tczt+8skaw3+kygvXal
0/s9ieTwZDAedOAUfdrX8eKI7G5ZtMIF672S9+69pL96EMqeRC1XpqjX2LASZfUlj/SzbDjQUeld
fFP67urBD3XuGjkhYT7p5FX/Fkk+hRNq90diWdpXkTPxv0ilX69Ugoxuag+XNGXvZdbhhGMxy1By
8lWo74AzJ48Zy9gGW6odXdjEhDJcUkF/zxXCHE8YS1rITjeVi7dgx3z8ULN9nbdkAFwiLRyc09yk
0wugDR7tuN3A6sbc4oCXf33LJCdHW1OS11JefiCmP/NKL3aJDanTTgedZQ4xB8uX3uFooppWKw62
OLyftuBNjL90/TWc+riEerYyDBBj4zZ4EldW+Zz2saJZksRib3/+Kmw0y3qGnpaEdIq++bR3+hnQ
CcBslztOK62cJy61kvyhgSUF5d9AyLv7zO5jZiNncrRtV6y3O9zYrgPYUfNkLoaFHgDtVbxUlPEX
+sXC/XhoR8PqN0vN/M2WVjlj+Pfyl2TfZmQajbeYf1a9LXKC4pZhXAtG3iDTaQxcP/k9/eIWTuR2
LyOMP2/9SYYcV+k2O6tbujtOrfsa44BACiAPNdRsEwF1F8CASUNIYISQSCqnbAWsUH06ydmEJ0Kz
SapAMSgETnve29hI9FamwYvXasRBdF+cUlkohIIrON7TooeVVONV49iI44TuCPpfRF0Pz5t6ISNh
+FPj/PvhYTCOJ3XHVlJ2i1IAk03k9wp/f293IlxB4iGbo1WyFjwIFPT+WNDVRFVdW9RVUqZGBQCk
Om2uqg9toDaFYzJoDA5E4oGMKVfxePYw3i5sXCRiIWRAaJCcmNOUCgMA7G7hn2xEXAdipG4fzsKc
LF1BmWTQ0e5wRcyjGZUbc8q3zvDYLb8QqRXjrTE1nqCkvIh1vzwjL8kHnt9oO2DsWmy8obCWSbWz
IZaBUfWw4KJfGRMi1I8ozD4PLxm2+GvdN6+1l/bPlD1egr5TzUwyTcvu5yDIO7sLhPGjebCl6ftj
WeOxfZzThiSU3oT0lIQNen9XkL1uHUBGakkEcUeduDiAQSJ/9HSwiQqUKibQ+ijuoxcklYoc0Jgr
5OhlQt9NJTSzjb8DeSLYbI202GSvgt44OiX7o/9XO4Lj66u9Su+Hf2fUDahq8Tyf5wlJ/xY6ucD2
B+PTw303JaZdjmoA0F88in9aZ/wNkDgroGhQR6EFxdCycte29AthbIIlOI7wPqX2PZJvhprgMbMF
/yvXC8jDwET5vUJkbRfGX8s0oz9Zr0CwalhFWD+ib2cLcz3+rr8/6SLkpo2sIfVyL2/gf17+kdzk
eaJCMNxXXSV0Z7VMKq78NyXnRj1s4MRlDucPkbDOQnIR2CZnYwhig6YFBNvONxHjkWk+zvPj67c+
kK6t2t2QrfjinDs1jhsRwRjC+0mORTe0pc8njrpoxIDlh0Mp3VjSgPwdyYAokOdovkRbIVJciCPe
k2Gyd9Y9LMpqvXl1R/xcnp/gnNYOT3rAKl5SLlbKKsr64i+9qCdyw0VOlVpJoX/e69JyldZHovyS
TbHj43C04p1j1yGZj6gtoteOkXKkTgeBxEt5VZIGwaDwZtCuftuXqHyNX7jy3cC872TsD4tLD1H0
3xwzDN47+3N2c5+xtFKRA5CBBzKOhhSYBZSGq5v/R+GYNptbUEP1BHvXtoTlu81mIfsqHmfSpDaT
hkvydukALYD6fqciiTwn7gkPV5oJ8PJPY+AJiDWDfL+ECA7VX7NFw1KyaQcXjNqiur95COauFI9p
Xx8aP1espiEy+nUsNnHbqJjd72RLDmqK+xdZqCRdYlwxPAGfGzRBI7R+AUB1AASppZ+eq+lmA4tV
8AOF5YX3oE0fGyvE5wCTIHSIYuZHe+TrHfzcZBKpVTJiFhIqBEcInVocBn6I8WBx27/KZR6lFIJf
XB5O4XMY4H+NQVVL+pXEqssDLfvRnomEwvnhq/g5tq4rLSpbTL0Ff/jowuWYGS9nCUpQVPQwzXjO
PwSSYScNyyshTACRYgf9kxa5jsqqFo6XvagcjeWF4b+dKPJjXv0lLeRNCoIUzK+EnOZlWcHfHIjo
lu/l99SUDVq3Mjyp4tAikPZZFaV4HU1YKKDv+w8FQOJSzgazhUnKg5/Ie7Qn+/OtzXBdPU7xXvhG
0n+GQkLE1RD57B17B1Jr0lsyy20iOGQuexR2ydlCkV4SGMM4VeWvKxsr6NF9y6eJH/wg0ybBc8ya
EUNOYYc96O8ULdlX+ZUIjc9A/6ph4ephRzIPgtjC6JU4wKMdqas+IeshhW23FbyqxZR/NCdON+IN
UPTYuaLSJJExkNca7WJQ/no76MWYmC3p3VudlFAFAdbYjlXu274ZuZM6KjrhC6sIc/eRij5hjazs
6xuSfg3CVm1H8rOdZMy/Vq/Brqk7TInDSYhyyMmQtihoYzVE/cZbopSMpY4F5uC/SiNRGVOEX1NC
XZX9gLqvRg7JGk/QfAuqNWtyHjc2EQUiJAj01XzVCrPL5mV1ZD2wzd0v9j1rjo+q4Che7GxFlG7w
EsDDn2JLubhwXgquTI5avac2mto5UUZUrqlum4MrngyFsDtH0okuHbW4ZxqlZfGIMUZFIIaQqIkI
I/Yc1ZDJSUPke9k6iIDbUQlJahV3QMgr30QHn2FH4/xMzvhc1WLCEf6n6XUSBlJZAscG7qIopiyB
jXSZn/muJjkxdHikWYXqNkNe4jcfOAscL531BzHT2hktLZ5fwvz167apmdLH945V7vRFSO5DqiTI
ff9/lj5YkKh3f+Yw5Q/BK/e2CdyjtNkfp+unoScqzfMS+R/o9+Xm6eYB4KKxE4lSPBrQKK03zejz
PSP3jo4e7RMY5hCskqenjl0dl/Y/QQUCNgz/BKuzbgYKERo4GhxiSiiSTv/58AtiCeKqJssYKE6l
FB+QHS8+/uRid9HmIdnew/m0oQUXfcjsblorClDXVeeZjrdJe1D1TCdG/ia4Uh861A5jY1x7CbgD
w1mYhiz2UI48xzjXEak/LM3yRM/ygAlMxuNtMReCE9e9vFehpL6BFvrWvzKS4P2G5Lc6I9I5Bl+F
mYOI/BgG9AOVE5VNFdLFZjxf/6r3gO9xpmzkytznpUfqsPm+clbPD6gVLXliomwVGUl/UHzi4smr
HKmqgkDzEIXCTckB428VueSaal4iiCPnlG+wKVH00QcT6ZxKBT8TTHDP4NtVFcBR8FZve9KgJp9p
YfhBEbGL7ncG/FYat3dqEyRBaZw8canKVQvjrAb7WypI9gYk1fKOUxLcP64IEEaTzislUGI4FB4N
UgOg3tLTeaXZOGoiMOCbVdULvPtrdRrtvNEqheuoy+czMVPLXLAHObfVV2fZgUJPKUTP2m1aGkEw
F1FakrxDh484zgdgszPP7alAtfTLg4BDPQlEVh5RirapPV1jfDrJFZ+634q0E8foopV5WO8zK+/d
Y6in8AQs6P0xglImYJfbmXJk+ssAxf31Ca2YRaQ5OBh/hQF9UTK4O+LVr1YczOHLIuyeKKZyvWKD
WYR/kWIbPsDDroVyN49aQMvEIc8QZcERX4RuWGIr+oZUoU66OKILKhUPizjhgjnFgIuZnlnUOgtS
G1IA7TNLIlOiMNwjbPLg26CQULtPfrdArzMpAQ1lQKGRZgERSIflJGmlCyCOcq5dZRBona6P7Tsy
xRdfLDUSYPV7EWYALvZtXjH79nAWTeStANcjnHYs/aIJRlm+/T4ekKhkDj4pY0q0SrjwiF7FcN9t
fYwgZOEEUyaW8oUFdD1OZclkyo3lvcQ6CTzfJlfiO/JvxgIhZI0oos2i2Y1HuiSX0ByGGLg3huys
XHAseTZeY08YvzRP2DLPElYPs6rJVvOnM+S+T/0on3yXTQOm/Y3iTZATJ07QyfjWdUTFh4EF7gnJ
6xAHVUcPq6bqu39lYQWQu6rdPxbMgNTaFnF+Fyuz16//oHnD4twK2GSPXXGdJOxmfMJMydh1FNNB
4HCha1bNghsMFGvDnxvikLhlGj7zY7acubHPGPyEeBEyx+qIySGjNg5mDblXjOJPhR21cutU3U3r
G1APMY248w8h072kYZrSDBSsOby5EhGNZ8gq+o4h0rDpdrz1lfC5STxcul1SnWPymJzg6YPPx+gM
OATc8b4MabxC2XeViGMX1B3Xpckw0ANElqF3v1mOFWMeUctMoxykBMQ8T76KBmKwsDKSqOjpnfjJ
oy4vUeFdZ0RH0YNE66BUGDUHbbFQNJIl7pDsjF0K2bfn73CHe2xaYXJP2e/Vbj4tsn5m0tbhfS3k
ZJBf8eePOrtnqpz+aBMd8/3IUKv2UjhBoK0lvrTlpA96+URfnWuFHkP/h2UaFiI8AfAljbMKMtLu
Aft3FMR8rRkTajmFKdtS2kRY/NyHdt4mA+YlejIQlXpfEc9XauzA+8Xo2NTgKsBabEYbo0q8u3ek
ZvI8TEb8dRIix6p06ZQ/J41RfpAq8VgcGzbtWyWvIyCDKb5cC2agbLeC0q5lPu+zJT9guQv+KQ3o
PCTAslcq8PwV1mT4aaH+o+jABeXY5kYMbuzcDPR4OrOB6MMoTMSskYFaW/utKC8779vQft67wM7V
2L8Z/SPWl1GcnxnFdcljrOQn0qDZPO3MtEAGgOGl28LLNsyMSnd+ZyA/DxGGlvPv/XCI+/CWDNRl
6SkXluzPdfpfyln1ocMFm2PlqmWUAWz+VgOPd3nfIOpwnpiaTKrPdRRjgHJu80g/9cLAGyCDAuVf
9Th6EyzgTAO+yixKqRPyxDHv3iSQFxmTBVNn0HZeygK6L3BjB7Eo6axYoKL4q/ADCbSEc2nmWzz7
1nOytyor4qX/8VqyyQd85tFzDC0EOWSen+ezovNJmBjDlTqy7A0YpJiYLT69ZoaZrH2bCb3lTHpK
22SgSemWZydSs104zmUlBKxTZ/f62Ixq0q3kNXMfb/+UbxKWK4JfRpekKFdLX7iRy7rzS9r2Kud2
plK5ms2i+idt+IfrMCUK7TY6PWk4vce78n4K8lUmEOzoUtGspW3LXlYhVxFXBgR1jXliKMGu/GeD
kLBlUOrlvxFXhfjJkyvAblUAq93A+zTl66UzvyglG1EFhfr1TI4i7AWDgAs+lQFTfJF/vJslfacI
xs3sg2W+SyX9xVxcK8VLpj9wbj1mMfAdfkmaFRVtM2TdslxdhvRu/wmUs3Wv4TU8sCxknO4aylxL
N9k/cdtSoNAcujpj23bAe5UKksJcOBJA7eOGWSUXfDwrgAX8ceKYnB++Y5S9opm6kvugbuALbwqf
pt24HaiMfZB9wxN7O0n9rNJlZYj1cj4/5CCRRtu5g0DZWIixmxyhR/wBrCmAL5yqiyM6h1DsS0nx
fXAWACXu4TUVgCxJkZuWqyuGSMkCh7svEqsK4Kg9WiwYNAz76o08embE/NVI1JYDs6gD6TEfcHKP
lXkARH4grPj2R9hoEntf7mNIFq34Bk7LkKddwpY08qZHrp9vFH89Akr+XjRbTQPuJzL2p5yLg++X
Z6ms57D5+Lh8UAbnle1CnGLgOnUUe+UXRpbBfIuYFVnlha6Ui+9yv9+Ay/RKrOdIuIQLwfXsdesw
N6iAyeO/DZzAs3dHMf2eApjCIx7KXY++YyjCnc9OSbZj3j3+bcernnMyS77wEDA2r/koHmAhuIqo
40k9s1PZ395YU0vT+xWDNemueikPTvTZCPP16JW7caGU5mwqVsO6p3LQ90kgIcVjJugipitlL1OS
aj/vrSfY3pSXL1I7TwOHy8lVDGHOsQED/qlsrLpIzGX/oaAj5dV2pmQKu5wGoDdIgrkZOB19MxWj
44OSS/N7AY7Wjf8umwB9sBbNWGvpGORF4rQCvenKuIQoDcRNctoXthoZrc5RYyEX6aXujX4ncIxF
zRgJOQ/ZbRoGRZP5Vrq915ognBLc0VrPoP8e/EiGp0ok9ZrS3YAtlvclp6PflfKPR41yGyu6+E02
9DOBIS6PP5xGs42cBmRzwrmMirnSLZSczyn2E76NcB/QjLtmog/1vz+7TLsVdaJJFJxSPLU8320m
wC4dMwgJcpik0ulN0pX/mJd4ERMH48hKPoJRBG4uyb5j6LiaVwh0duvPFo2c1bs66IgoA1FROWmg
0F5Fa9TS2wejntYm1N8PXVuAXEA315UuqJTG/pIOyuY8j6LxhJuTNE06JzOBgbchfatyAKCD4PvF
ShhPm6m9j+iib305QbSmoiU/XzH1V3SaQfWRSJViM4jrx1PCYz4oi+iMCgY37/GE2e+Gb+WXu+3o
OEQ1FgJU4TcUvB2o4aEjYOX1LzrYp370nqypzCSUdNM0AyB9gJO78iUmtcFWCemRjaQyYhZoTc82
k3qmvw+eGdxV9If96l31nHDGT8+oW3M/U7dE28PfEzRoLkpG7J7icbEXJaF+sR7HmdcJZrNIqMgl
G0A88i8T3JKv5+GLzkhY2kk7LxD5nXfX9TJ/cpVCOrmVle9LmfuMx8XPybTjwui6dTmOnQMqch49
6MvYQljupKqN3PKkG9pYduB4+T7n8sqBIR00EdGfHuI3jfr0/doH+s1vqr9yaU7AFBZap5Z8mE4o
hAS4a7nI/IBAiXvLiYmuXluyTaamgylp27JqqGGuO+bGUty3dNQ5Az9VQ4q4Ae9v3T0d1dEs1+N1
fHJOYV6b6V8Bduh2/YxoY2kA6AoVMw7vE6f7qA2pIz7wfdMTyP29qxyMuLxx7QVbSOLfgyrExdE3
zxcfPBx4tJ2qNXWFQGP8SK5upGb+yXoIWoVrTuc6SB/HYY1M/0Mr9/TRoJW2vk83IZrRXGdEGvO6
5JPeC2dLF6AD3COSwJmNmV/VZI+sKAkTXi5MBgUeYRipFOrczPsdzuEO1uGMarXM2ey/cYwZJ7Pg
yitckLdLbxUk4mMuPOZl00WaOpXw6/AzveSv4T67iWRDFiTiPUuApKQpo5Ce82G/DnSHi1tWp12/
Pld+igtlnQXxhpHWsHBI9t8mTeTxFT33jWxgkpBMf1v3Jq+BseciZks7HeWoOrYh/TQK4Oeg19wl
NI99CbqaJryhMzTCjtX3Ehmq1xJHoyi8JMxvs+d+OjGMXSAwu/zxd4CSYWIf+HCXz/V+PMK+Ic/1
j0S4kYPOdzZv6SehaxX0tRHLdaB0d/+ZeW94TXpFplIEEbZzDzU65LRI3zDyEIjey3XxPwTxGstk
A4Fenaz9b8IBRPXGLE9jCpwMmf5LQ3IKKOab/UiMcZZjgo4+XxvP4lPYJFewGAv5uue+kaaq7xpd
bsatZ0qk6sboCijRdnfEYdmaFCQ4oVJyKwRB8QakuINrkjZRsN3z2TR61s+LpcAWPiF5419kc4P5
hhY2p5AaRRpLLWEziW2c4EhIYqxnK4qsFiKILeZz11cHpfTWzBi8D0W4ntLtxrj3aVNAtiLUE2P7
wMPl4slh+UlbqXyVvAAIbG4iiEFlzZn/NnSRkmsRrUJLHxFF5wuX4e19lO8MGEMxP5aIYj7lhX7T
3KcRzMOdNKi930W2bvPOAcTcDEJ5E9iQo1rFODNiTILs4X8yA/dWltRhXDDK74FMoxAPC+HkHKIZ
VI3d5I+RZcZBxNJpKUT+dPPkdOWL4GVv5eI7tukhnOel0LlRxi4gLGH1Jx5XXiSY4pDp1Hvgh3w/
7dPU0dw3vlhbXXGlV47+e7woqTVS33mI5OOKEXQJAXU9AfuUZloZ61JnANrEgGEH3Anc40zYaHPC
7Yj2UarW7tGP1l8v8wvlnXmGnucAgQhHSh1ILoT3IYma6k+zHaqxgpTSfgJrXef0zi8vYuU+fPV3
86hiCanSu2KIZDT8ETtxgzK51s4IrtWTANQBqRxfh/10PwUxDC+9SVGDUr07P8aDxID1kJJxMwOq
pHevyb28A/fYk3OpoZ3aXGj3CDPYCDKvgfMJ0QJCr7ZsmE4n9b6OYTD9ZySmUnnoesE0ReAdDRuc
Dfrk4OC/6CY1zdn70fVZy/SQ08EpIV4Vre2POhHz44UvNnSbm2Xx3FhT6Kt+zs6+/6SLruUO57n7
P1zYZ51+DLbyeU7jY3os+qJox0HLD05m2Y+NFx4Bkf2dmo5T8/zhxkfT/4bBlw1wVHroItnKy2Yy
PIDQ2PuALxAp98ctveUQDSTUVq5d1Cwm/baScnkxWUnvmj6CyOiTUndBPai4t05iyfGXfjQpqWIu
z6gQjDbf+1Af9MjDoESNPvmgjExiPP3NDDo5FtZ56yAr85geez7tAIGD39N+hvZn9S2Z5aLiR5LW
M2LZJX7PYfC7eRoAC9Q8z8ykz/W+I0Lcg4x9Q0sHBuqYKBi74R09sRZDG9s3qCXsUuRt81pOx4Ee
9VRUJBhwZObDYbdr2sr6wUV5FYETnK2CVGYvkGg4Ya2p8GpEoGpyU/dnU6VXhwygg2u3BJrb9nza
8p+TEoldlnFnFduCMgLZhwCc1ptKXKSL4NcINGQpOQqaEHvoPBB5pPMZfrX+B56kMmuvOD1Co5JU
mivGdrKde+3CryJQZOSK/x4rrhYQTPqlQt/DRhx4XboSq36tjRndMXraguQpe7LmXkINsD9izX9K
JOg44JusJUrFF9dM8UJ+Hok7359NLH4YGr/8fo7xzJZulBvjwD092fKrkMqhz3dNpziT+CduvLtn
8j8JvEmDC8Uplvi7ND4dm4V2Cp12eSPh1ULfChzLbSgfZKSJaZq134VXx/W8Fk/wbYkXxHv139nl
QSgBztCn/ksHB3X0VCzhehY7hTSiP1kYpJbIp8oIAsvuynu4wD+0sBtVZyPFkuPP7Y4cPytnDlwp
Frq6Dm35AOPDtKh65pUrDlPGjDz7TdP3YTFyYtmw7YTeVIM6vUZDzxPuVMDpQsBaKwEz7/KKJIWU
AaHt0EqvWjmqZ5vJoB54NvWdopMcJSTfSaCcHrmgePLkdcyGW3qnnaJe3XMz2dOq0PDLakvm8A52
SNGXlPG9fTTSCG8oLheUti2ZWGD5+TyM5GU10zTxQNWxBqR+IPvdqi/j4v9N7iB66KGa980phXBv
5cn5w9HZQhlAVyLnwWyj1iZXvS8QwM/CKZQZqMhj00zGE225QtQU5KJN7EWirkifVtxZJVzGb8MK
tQF2cEBS5ynl+DPQCoKZzgoLO/YIVJRn6hea3KB9qKzKVvllZHptS6/puWL+QYaaRshgdj/pypYk
vWrwcBYXE6JFQFvQsgYqcJXz5q2AHAQBAtWDELEkSf90dPrG7vTmC3Lti4SkYegy3GLZP1v1bFHZ
+1CCLGLpbfqy221PZRMo5NLWB3javQVu3NYjNd1LnBJQZ5ragIfMNMvWnWLMTmZc366yQlEB6YVm
9663QJ2sOGkbrvGyX08+b57TeFVtGZZxm/ByVHIrsYf7sEuuLDlNldHvqJ2324Rb93NvjpRIFvU4
TapaZ5ISeykJ1vXI7fTsPgnaoZItYe2tfCMRVf7yY9DCBaK3uMEkRST3hPMJcHqmvfK3POJt3A7b
z2sA/1f9bUa6dxHdojKB350F5G/DTyryphLDEBlpKbGhhig4piJTZNLg6w9zXeIEryoF1TDL3rtV
lyiEpQR7EnIlnEGT2hYEF9O8QUMXEixVPqQXg5Bh2Xq58DD9jkRsumTNxzGFaz9BC4u4iW9bmd/8
So+MfVMpXyH9Zu8mdd2KzmiCc2tBnCh1PgwxQ4D2pthJeUJZBbM4dF0EDUgwYpSVEQlTEGJfKjmv
SHk8ZsJjOv+/m7jiZMbZ43UYkGko4Leg3gTMm2VQqLokJOu8M8nhMoVRFDmW2TryX+7Dd+YObe5b
p6HC1V7KIW/6+UUBumABbTq2rYeUc0a8qZKPOxG8RXBd5cXBILDzrJdfj6tW41YR9nFUOVVtbFqK
eGvxC9OzrGVaVp3opbNQ03vtmd/NkvoaZ22RolIHgBx+VHLYgJmx+jYoV0VofYriXYi79vVkFAr9
q1LmgogFvlENbSFvEu7GT2CA1gPmc8f/nOj4s/1A7QI4LtIx3lB6fiihL7sR918J7Pwpk/2m0sis
/Zx2E0Ql7kXSrqD/4SeNQolQYj9SiF9SiptubzKSdzpMMbu2yc1Q5xxXvlvESf/eiivt9skS8YOr
40VPcn3rb82IKwFFVVaTHe9FDFUpaPPvoIlT+AmzkVQjVg6bDQbE5bwOZBHQW7S/Ey34Hee+Gz7+
WY4BxNvFJF35vJULl7tnMF5GKdC0ZE6mIEq/O3RultZXTuSgdC4Oy54zG9gtBonpuJEXwOp0sVqq
7NA/MadSuXXrQtk0Wi5RXx05csrVHv6PxPUcGq1CbCL+thCGxpmdTyBJG1rx/LVL/9oj3z46akzn
djzgUSlVWaqp3gY5WWl2gwltM6n7Bb9Vd3JKs4Z14cB8ljJoF0ZXo5VFu/5sDDqpvquShzwn96ok
AE7Rgcm3JvKYksoLUmGKcZIpZGA2zOgwezA/Tos7kZay3I/PvcD7a2Un7X+HeKVhDiCn8xPGndW2
5bbEI2IxjAiMiznAg0M3d5Qe9rSE9R0+0TNMFyOWrjpn2r19oI3qHY2vJ5Vz+FhdGOsaXKTohJyf
GNl1OWjYS28usOfww7qhq61Z1HuqgZ6M8GRjuwXzWpO3TUKgFRRo4KmnlY9c1b1uEirV5Nrg5mZu
oyTkVbpeNR/O+mKM4gen6zSFB7TjNLhO8tHDdsr/zQcs/niEyeRez4+I32GjiXt5r1FMVuZwdT93
7AiQe0NltY4gtGzYwjO3a/+qUFupV8MCl8QvLNMKocAz5eDIs4kTlyqwRa1kkZLsIGYWWUGfqdN6
F07umrlhbdwZgRQXCeCLnf3zSG6NqshpuFym9cdtdMJJ/uTwL9+ya0NO69qduYHd52S3bCVN7y8j
QxsCsranZsP0/5t/BFZjQbMfduEM35OyqQyTBTVsc4VjYVTN1qyCDs0nBWnSYXrKsBGb8dUW0F8s
MRrAH/vPTbD7ZdEBEvotK4WEja1ApxxuxwRSzOQ1bV/oCQEcmTsAZjjrPgrTM2z6Fmj+yfRjSMJg
5aNgMQf0RpnL04m2daFBZs8wW0z/GRTG5jduYrjqW2YGMsWqDN84HtklhR9BRi3rbHo6Ol3WwJKz
iGOwem6koVszp3P3LhAtLO9awDuJhQio7RgiAnvpWSio+8ejQrUtcQObnJlsK/z0t30s+V82b019
GwX3b1kekP4wXIjx/P72hLldKV81w3PRXYYF7yBFnzXHhcAQVSRyoFN8A56x8wZyehx43HzEnfl3
Yoo7qKuSKGrMdqO6lHLMjlS6OyFjhJ7+OQhZY/gJyKd5i6AtbW8hz2pNxBeyQpOcyGoerygbyrmh
F2u0C4PO/blZf/1CURufel2C7AfZtZWIQwX6GzcVe/Xl2yJ7swjn9CE8pplP5FZnUjQfgSdLKC0N
uMeiQEXqs1z0RFNWybaXwlVpS0rpeneEJ0o3PO6cQi0UL70OtdnKO5lz3EjCBMAkmIOAOgebpLmk
XbNgW0d0fcZjlZx/id47D2ylvpC3os2fpiJcql9rf4SgDTJGoiUPthtuazmMM7UDZuZQXRciBkdz
iPRFMy7umGdJDmsLYjl2B4bPzqICn5U0pUEMt8d6Q/6IqUGpdIjolhVOBjlNKMkzR9aZSuTzI9Tw
kX2zOObgEFMtlTvnjvWWIwqoCqtELe0J6yl2WmxQ8kL22aiW3ztMpuuuOA/i71bACmTnhne669KH
oEW1mDXnjs4nlXqxFKLAHHolWJuCoInKO0wqUqbEanNlSYoN75uS/ZDny40qKGQ06g04cbHmXX59
dqOmkMPF64lXqdAkoTU75PXiDuex5M5gsZvxZSBB55Ox1rsNl30GRgtxSIDjKiR4E5DonBFBut1j
63tSvsGFSmbEgdQKqjFZR8zG7YC7LxQKNkf8yKEO5ISW2N+5LciNZPTxHX+xddcD9E2Lzun0PQ/i
fuB+sCqK9+R7OVrqVIE/TfhODTmstkvnfATlJr3wS0MuobWQZXlSr1jAMGJsnhuzuxHQk7VwphN9
6avcxaRTUD1Xa+Nzj+5Op6zcFZ3LunpkoLmit2gOQB+6bt1XslOreyFv5qgLmYq3bsT7ZmJcLaT5
QD0upWfn1bM8iRvbEzoIE9FkFqeFwFKJNr62CsDZHNmQcDeeO0EwxteDr+pd02f2iTGFmCQxneUi
o0BT0Zq+aWvCvnkkg9Y+G01GtBiNIgbiA1yxsnelG1cF2fdDUKxMsvOizbZ0I5VgShAFkK4eyPGe
x3xgunaBeyl4I8jlHMJJrZaOc+MhtXT0pOHp+ywshcN8gmxwuoTzChYZOdwWXkG0HUVaclrdtGr9
xeQxesVcwt9Hfb67xPGykt4Gp6Sst0qJGS465pebY9zrOlPiqAXs+6r3gqQI+emwpo5Cb+u54jsb
fKjBksUUkoFTx7QmOSCAG83Vhigp4N18jPmnk2RKT+9Ash8/gehjGR+546XVYutQrrNwV7w4HMGL
fRYBj840Msxr82AjSJBmxquBQ4LEoOj4ADKmRTDpQ/P3ujT1aJqjJ76Ms3h7PyXDS9m039Tx4IUu
K3TqYRmxUx7gTUzlWC8jOkyzkPHyFKd7OBE341YKh8v6qDSOneI4RUQ6y7d33G6iv6jb5C60ZoxN
4v+ChzbtG1ap3/jZtbqMfP05KW1BjCvRLTuZ6K0C/KZ4v+U9L8Nt1vWWUGClmocLYLBp5CMu7i/m
2dFqbhphcItJjWhURCVIPV02TaG+JW045YjC4SpaMroMRwetYRpeEO0/kfEcORKY0iHy2obHVQup
7CxngBZAiPcti59RjG50Iu3A7Qxw8458C4c16j2HiyTKhSS1PqYHHds+KNBvlwfUO8PzQYvrJE3S
PtmxBHYsKdyzV5ucQl2bwo1RDRD9inLiSoDXIF144/z3O7T9NYi/13Vz2+2boHqI/NjmquTxruSb
jV+UXAQj7Ozj1kY8jPC/gmlwCw1kQ/rVCY7jKAwO+2XobCGnhQhnzDU6d7AVF0dHLy7DKOLya1f+
85CndMgYQKKvYZIygFcmLeRetVTlnX5uzvseq2zVm77qcGEHvO5p6nKNNsz46cDTj54CNDIh9akb
IUfyWVScLPr8LCTdc5x8qxcOBempDY463saniacafNCAVZJ6JB6Rw4kWHX7NC+l1gBdqXoxmsp64
jw+U6t0PabSRoJmqmM3cOTnRa9kJx3b25FvXXVVI2PB/9jZ/vVnffqphEuTsMogiidEZVcLgCfba
XH+NcDsmvLcqkMPUDVbLqNfmrzC2bk9JhmUqloG3vF5jQRoDfeJbVsE4s+QV4P/KufPYw/0DYA5h
VGz321q7BzKBVJX46N+bgHCeSlxS36Awb2AGYDLTsChIF0laYrCPVf5i1T1LV2oK2wbaDiehqPkM
gLYO68d13/t3+uabpcCXOIjL2LhFFK24jjPs58XTTZ/+lEtQiCjN+o1kkWgyt1WKrQy1UPvjVCfR
J8TZwbUNL9jh0G41DdFwteRfT5srqnAANrHQijURZgmOci4zS0kAn6qvViO4oZW8IF5n21ZvNxLG
8wny2WTjJEgJ++4QzAdcuHYgHqj949uh/TG+MGQ+bXjhDwlT5WK8pBO7VBHNZvG6M74WYVXOdq6q
/MyQ/B5gusPEqewwrkHFn4c0X+3KItMp0ixmcKvu+929V3WjngKE2UY7WWak5NlTChMO5A9ZkSrF
cWdo4ypqnAwSLf0yArWGNKcQy1i7GNcy/5Brs6bhuOGhPAUf1Uinm5YzG6J48fznvpmvOmfMOk1d
SR8owZ1dFUCTIScSq7GdSMPSPyiEwiDPUU99AAhlD2Ez9vkOMgWCrjQ8EpWa6p2nRlDimh5LK5ex
wicN/xSja+zgPSQAIUOfZybVamF9mZP4o0Xb/OxGsTe33vHYj4CCW5sANdxdKRqsIEEfFlIA3kYG
E/OSl8U9LZrmimFsDhIatP61t2pZWhXyG0iKnjoG2azjbEreLnR6yyKfmbf1J/0MqhgS+aIVqmnr
N3yoHxvoQZQULEuFlXyQNCG9pFjY7k89sv6/IUEwaihCjY/+IMa/BmJZp96r/o0dD5fLU2uroDSU
qo1k57bjT0ZxzoBXI1REON+p0nQf+EmvUld/kIhgbk2ATUQMr/iAU3El2gJKPKoBf4BQkicFcIf3
ioHRf5D2S7bA/lwNSDht0awQpvJexGtxnW83iN7xvpSGBZXzT74ZpHTvGB2nlurd4iHNWJLI31aA
g03N/BkJGiIp0YI8tJbTY4t0Vw+bBrKhU3tx3ert6V8HaQPE2fk9tdxmBJcDfBG9GqhZBkb25kr4
dHk5vTAv/1tNiTs+w8xIEqdnn10w57Elpi1JsPuIXWWmmEmqTtiuWtVjesfsAxNJZW10yGubFh1Q
p3FW6w1ayX8493sq0h87WG7pGMCJXhab7aGDXiHQNJjiajL/Ow0iedQmRU9vcLNtKRbnrcmL9BS8
WPUtL0q3hfqGBXyf9/9L8IV+FGfJp/Y6B92RW/begP8hqCVIF8XneNv35m1hoD7CrQRQZy4pj607
E+g/FQjlLq7/pXWbnjWhRYbftC7Yr2pD3xSA9YwxiRpKpogVGVZyHufXkQi5SpKocBCH8Ws8jQON
brVg5IOUk8Ot7DOxr01ki94TjqS2zryfKK6pshXMzaFW4CDVMGNyqofwrFO7AGc2WeUZFAAKSOtu
eu18DUjvlZhC06+Urb7S1EjoRD2G4UcVz06BkbF54sPFZwcFmdD8BYQe99MK9xK1Ih6q0N84tqUP
8iskVr1xufUVrFkaCZ1QCBVGAvQOvEmmfXQWalpEij8Ws1EMTXWWZH7yvsyZym8V6BFSY7b8fSfs
WiCJn0R02OyEO55SRd+IqdRU6gLx56UZfHgAWAwvyyAu+NFokP4TPxiHcE9A2RiOAEo/cdqntuIg
LTT78QbAaAO8zr+cUhGA72dBjxqnY7Ffq/cKjP5HXXKzuwuN0EkxvR2YcN9KsKsMsaguMVk33an7
VkNlNlRs8CIdPmlJrTyUP/cJNynxyUoJEGjT2OxI+Hq7LFOdL4wpIo/ddxw2sIzg0fX8RkMwQI/a
Gg96ogBp50oQb0V8325TbaocPSXgZIfk2dii9Hwtwmn3KKswO9c3/2KpLhjgZ/aqaUH28T93RiA8
0lbcZkLaX1rbKlgmw5B4MvxqRGGsQXvSqVEPB99cKPH7cFtMRdvGdekCFyinLC/rujnBSqRd8hZv
B1BDgs3xbxFhhVDrY+EsqPDp62NchW4JnWdQDt7vo47fVyUdZg8nB7DOvTxBEujxGU7Mb0jJ2fKH
/TDaOwGMFFEIzxXCMIBZrK2F+Kt7wUK4rtWJ6wvL44MUXS9O1DaqoDiwLWC+dcA85sh4wpTLGala
ymRpimvfTk3QZBP0gBQBV6QwU6/TTfedN98GQeR/yAPDMAgDHS/FlGZTEDbFQbbCxbra+3f1DYhX
R6sbqZbfk1CMbeOj9KlyAN2i7ssjNZIrXWx98/0MMcllz2/lzXoCu6DvT+q/l+LfwQCpzkV31NLT
Og0mZaXnoSaPuvt3fU9HwRPY61evLFa2UMjJHI7Z7BnLvxI6WctveDcTt3Dg6mC3nFjFatLKv0gJ
yBi2efBzrnlWNYBCSpfqjgFPHkzUP0ZkdNeO4/xUxGukoNYz7hvmkNawSQSnr7S9RKjHK4PSC0dr
uSTmdwmuFMGSX0JWZd/HPwIBVInUe5pHMRHYM9zmUaK2AjpVJoO2jSin3ddZbL7nKZaDSho2mH48
MrHIlh0mvu9n3YGiu/ie9titOhCh1O8BbI3+OlJWQRSHFP0G71jVmUnLLLspML+q0OZaWES1OrA/
gUAIUy9oD9wpM5L6CdIYqxAWE2SpidffqsEeJZ2VIiqRdDqtffYpGD86DyRfkngk+HeojuRa4OHt
uyzRaOkeAmnpesw+sly457131id1C5LpJ8KG47hZ8bNZGWBcsUsDe9COOpbiu3ZdfR34Rh4jB5lq
k60hbTWGMOf9Ykl546ua3kZrEymp6y8qrjZ8kmP/nKp8D8qn2RyYP9tJ0Hu2+VQQZG9+LFO3q5oE
1NNBb8VZqRCxRnjNK5KbzdrI0RA+pCIYjA6oa4nh/+0gusVp4h51O0piMJpRZdt/v29JcU2RJpBV
tPapAYxqDNkahRzWIPX3KciNyQcjCt9BHkaQFsrs3N+dMX6g0iqQgKzUGgZV5CsK3kIUtErkIJko
7GTe6iLZSRhmCG0VIJwMAr773hhj4qGYSjbbDAebYWpPdI4NoNzRayH9jrMD0ix4msYeINkiYAbr
htccQMi7IgEQSxyoS6TZdqXNhfAcjjHVA5pA58LuA+anNAlxE2xIC7OWWNYMUSihzxy+yboDO7l5
1nqo4IS40SS8O2aGRnICJr+y049nnayo/DNYh3LPtR0xHXJR5gP+o8KPGoYtUPOIQvevjYFS1tNs
BiLJkdPiycrFLuL2TxTBMJwwPlxRgy3/BIpcQWt+MyIgChnbudXrnJw0jzGK9Pa6UflSQr7LflAn
YcgsRfJGlV4PWXtgpIXVmCqwSa3rjOguXHM+x/qANZSmJQJTruJ1eQwVX1LYfKaXpcsrNpL/IlOt
zl0w1nBAFYV0hVgUL6n/O7N5vjE6mbRNqEFwduRhHmyBwhV/zUXxgSqXr8LpKujkC1kp0RS2zsdt
fnYjqeNCIpK7+4NCAQA4zNRjHLHTmSY6kPq50ZW3C+MjVxUA5KLPHTe0Y/AH8iZl1uLkHb553Fv6
6hSVTrh640vwQHUSybcHeNP+ezWIuEBj6SMkTnPlMNh5HRzWJqPkTAxcdXhCCDK8eTQGzigQdjW9
X7tNWmxcbzURaG+EDcIwInUauz5ZPJm2aU0UxxSqPxSOtVBwrZlGtU10ysxDl5Ys/oeI5Hw6BPgj
6FMVdtaymtGzKA/SNOMn2CRajUCe8I5wOA3uzq+OnxrPrSomW9iVJakW2ZpvIIKltb9KnhdkFxrC
qemEd1TNkYZaln5ffVcuF/furmHkOvfOZMo5z6yoMF08XFJTk48lV3fL0sbojRl79mUPNzazgQRO
AlaFqTdB99sB8Smw+JcJLsf5BcKTluulv52D83C4AJyuaqinbxAG7oc51ZNtfx/5+9r6Dq7KHQ2m
MrFVJ18M+yO3e32TxokVCe5HVo0FlvwpKrhs5KkV1niqtpfe7sgQy6oeop5E6C6IqhrCateUuCeh
RuMKIGZLpXd3fZFAgGmOkpW5SKIFyTJlm+5I1Lm8jBDI/XMpKmorCIk08n+PRcR/DM4mQj3EJq+W
RJuROoTxYQJ2efyWyplyE1x3zmlPQugZlc8dSN+W3+oeYq6soJwyAhrEBtNESGkN1DnRqkyZZ/cG
pAH6PeMWtgPKZFENeu2cPVYw/sgiXC/Hpe4aZOrzgPbrbxWNkHmJZSp9PE/RKBo9Po88QvGQ5SUP
tK/3eHiBj/AHTLWFOtfbpkX8zaNBJ41YdWZnU7alxPFA9pxvmN0SSygJM3enq3SBuLpIvAvYQvJD
rhB2ZQmNCXU34ktKzgcGdyEJZx3szjJguhU06+nvTBOpCYYmUp+pV9uzgY9ZxJSCbY9B24jqB8WU
h9e8pgtgLF8S+3wCpaEP4KG/Q+tJDtZIG3XUMJlfLBQO37ODJvyHR/rZAOg9nSPn0CCDuUYaLLfN
csmf4/NpRlb8FyCcMuaKDDs4lKUIj5HUJJUD4GnOzyhW9k0fjI95k/GF6KP7kbbAiSU44Vj8yGUx
nREe63kc8o44TJ+q7EwI/gJxbN6Sqwb+LFZ2AACvbGJeN33wbpJ8XeU453z71YF3vP58OuS6VWFg
KQsvHKFeBCiwjXG5aUwnWchIaSB4p4foGvKUOwG1WDmxCRD7QNx269/q/fMqES5+pSpKyXFd9BL8
zchdR7K8XgBZPFj2XHapUY+s4GqQmfToc367YqSg/0ihdm5lRBQ42Ih2j6uQgT7QmuBkKNdEV8yT
F0FZ3pNVMr30X/p9GctsL48KwOuFn5YSoJDS3ysWLdErDOzxBMDjG+yJY/WDUWm1H3iMjQbmo4iy
Scat912zjTl8aCPdk5nDQDpIzaQDJrIBOmItnH7+iCl9D6soPei5CsG3R2vRwIIFm+7XA51w7XLk
1fKKiv5zM3e4EoL3if4OomgurM9KJKs7M9D+edkTAV9CvdT/SE+VbdmzcqZWuMm6E6N5KtA9GJwu
ZgVJgPz9ZhYwEm+oz5CbMi3TY5+wk19Ue6qJ1YI24BDrK1Y35hPHlMW7buWKGH2y9RI6BTWisW1j
B+PyXTY5EEjnys9+krlD28azUTRFUdG48wLyH3sZ0V3UUkcCpXih2ki5XjsB0iNdU7McnWoVeguv
frzVlnI/CRIl01m6yR/nEmCVa7WomvQmRlt6FW/5f7ObU12pbRjG+wL9NxhqZ9STQEm7soRShG/Q
dJe6ppB4zmIV0UMl+t9hReKG6Db0uPS4gtL8DDeLoBc+Z1k32bJvFNLKfoky7hPBUb5pyvATxPD9
GLLaT4HLY1LRWqbG5AhscOLrKrfZNY7zzVvlqyqqc6aSncInlbxS3/gJ1Aiyj3+8gF5XEwaMkIVP
Pc1nug7kMOQqsgKiBxsAb7qqJszvyLfsvam6Uw5j/eJVPHSxdjV5VR+ylUEgX5o19LVbpxQeg8Af
l3W17iOFql99gioGOv2ysfmk3q78G9kw8FcS36Nq9ZUfU8ufiU+ozXvs/WONjPaToXqv5t0RSiKp
6t+UV6IDGU+3dD+ITMCBb9v/786ePwnMNsAyOy1DjA1XC0+JctGm7XM6JpLDVkopExfhjyOIBjPg
Fi442ibp3CStNuX8wMsjdGsIUd5wo/rebdiO0cPfdyWB91ryxLvH2PgPGYJmQM9uEB9G8veYfdgi
Qr3ytBIIDyk0XupYSEjJ3gdTQkTLQ6gYFNvnufoTmWl33NGXdqxcSJiVVLIhmY1wzQkqYqNFQybg
IDGoKNm2srfXVhFoD0/tMr540+SKfh091rpUxPPzx5PCFhQ/2YgpQPffQndUJxYmeCDmMFTiOdS/
4LBrF1DnzcYyZ/t3YxrXqfwicYsLrsGlKdxSw09aejZvC5UlLoPjTTjFSuKOZ9JHwfRKcKSwFhfG
6e2TaixMuU/tHx9o5fu3BVZwM7XF4HF8jYk2uQh4LVxBxidY8SRrDRD8wAS2a7ZqGi58BLYFct3t
7ShhKTg7+LHADLfN5x0oWelhSscZOpC350iLWnXMO8JhwkMirW0DtvWTgKYu7u0JhccrYplrJZJ3
G1Yg6u94/sJUqr2eLV4ShyFH2fGc+3pzSQ3rPvHjdcNmOHSmqWZClh9DGRGVcilXHa/qKwt9WKZo
n7FxnBZeYg4MOjlB3LqciKJqSksnZhQ3hb/kFpZdVe2yCLBrgTrQ1UAklhrpbvPC4MGOt2piKWSo
+gfJ+jkSmyvC1tberXJAtqHIyl9BB2OfPeKlyW1sn8dgIq7dtN7eSSOq7GSBZXkN5vygf+tFjxjg
kBMrncXR67X0GHm0ShtnkiTFlE8vKjqgES42TCQ4wnVUA8MLrRCJtH4lunWoa90aFTFatuclaI5d
5HRUAcNOxh5NaUhn5auceEJ+XMcUk6l65TW/d3sQ7M1zgKXCLYnbQYyYjfBBgRugwqkNeXLLTMCT
Tvkn08aLy9MDvBSTeJ3NU1nmcdm8b1FTPYdTW4fVxHMJdSo+quBB3UNTvCGm8UawvRdHPS9mObbx
PxugP175ycDpBfdTo7msvr+3riewGfUuMqhwbCgUc3pHmYURd2ZzxCQR0ESvtp/ADbl+Ld/o2pF+
V4ukNkoTffGnazDY7NHMh959QxXY9GP8NiDR+AB1NY1G8uAlf19+6BWC1HDlgEfScQXmJBw7B7eR
j28PHp7jhL7q72MqCq0hV0wPa/c8tVNERgvsl3j0qqR5BEV1OxE8mbds7ojy1LfF1wxnjt7iVTPY
CRAjNN0WR93ZIiNGP0TrIKtGp/2jYvUER4IjRFaS38ipA1n0hlLduAcoM1vpASAB1eQQfWQ4gPNq
Jwb69ipktYWvgPhin37vE7ys03hN0j6ZjBq8CpA8v1Le/dPA/Z5ZMyCbkayYN5G1gkoD/c+UGqiK
wIzzWj1cFuMsAWJyt3y7n6tL/+pu/cTC9MC5mIIu9DfmYeDHh52UkosrtsbbbqC7gkpUO+Dc7g4T
VymSm+nKKLhhPiEj6qrzlualy0FDwOYeb9XVuHnnIXx2WnRLgVAhxDkutOwZZ0HvwUNuR6GF1LMX
2SvtSnCoIlA87zxVzCm1NSixSGhmbZ/PyIP+cGIIIjxpoXFcwOnnNqO6euDg/mE44RsiZYxB1BJW
azVLdOvcn6/1WKW+Pj4IQQAMqd3eV8oNB1TPlJySZWjm6t8G5mYWC9Gea43slerlBZIQzwf6iC3v
qKThY8m4qAYW/ae/5onoet5ZdFGiG59GYZ8HunshPrDNqDTNw9xC5iWbedsfOJJW90/flqMMGxNF
c/0iC/VyWu/vzk2U5+IaESB0KkAYH3yXH2igltXYrQ60Wd8f3NRDxJ8/SbU+Z9F6F07khaUcD09e
EevuljN3XyxdNdsf8vzMHF3TZ2PJxEpHtk3m9e1qvMyD9OmTbMAxF0mBUAmqbtgDjvUEtyXp85Vm
nFt0RttmXXRJ2C1w9rvMseEQi/rGgn8dTbk1ryY3nKTHs+lgVPXFnZu7KJg2uezYIdk6nALL3+FV
z2PDE+Fo4LQf+kgNJ8/VbL/q1TtDss2H9D3zn1sfQMU8YtkFJiIBaBzmUM5lD1CJ2pVegLMmsL3n
YV8Tudo/o6Ox7Zzi1KDi39iEBKKnpSL+aWQkBHY7ob+xAEEDJaAWluKhrHONusdJzmk7JUWTtD8e
YQNn5PXzR49RrCvdBqb1uAeTY7EuR1jwRlltiNjEreNtkuPfYPnoIUbgTeaZgxtBJVXhs0OQUm+5
AFiGUnDFo0ofT2Tai2HQgeO22Ne4yERO/7R/eJxeTjV4tBxs4Q0+YhmffEfinHHz0m+g3heHDsF7
Se11v1krhXqbGVxlO4YS6MYkKxZAnyF5RWlufuplB+KjUcWlU3azLExIszukkkP4BRb6P+/5hSZU
tRLVJHEusx9Lo2VYBjqOOe9xVnvtV555F0ScbQ6HO95d7en1kQtszq+tgV9epFUhC1k6nYU2XX1a
9+B3ATeyqyP45OS96kSPxmrGa6+GNUMQRwtzfprH+JPlRWddD8utwcxrhyX7a/LbzFUwbIgYrujm
GppyITSYl0+fFkrxdTEVhhT9GHHQWcMdAZ40b+bEN+o0gTd2KwwlpOYEBKTpf+Efusd3ZCWgnuCj
KFJ7gat/9/+UGg2H1J4FybOUP0j9zG39U/Bx1IjM5oH/S8IOY5ECvzac1T7OoPSAitt58OQQCMep
Zlit8LQwORIgMClEmRST7q2LYsN3r8lvh2RSRFV5uhp3l/L96qgmRsAnYxrJPqhlkRm8N7TtVC2S
YyA6yC3dIuOjNF8PTFBAG0h9bnu6eLZftwAShYYKZoshfukwy6iGCA56ibyzT68RsD+VDREq2ieF
8Lujw3Csgdds/T3qMdL4zlx1GBM2zr5taY641J6hcuaEOncK5lE1TZnAk03uK4cBpcsdgAEAEp6g
05bVBARgciOKpJ+Ekrt0088MXdxK/uG34w+vAcmjYiTrQQOAoaAdh9wEUpvcanQuPJsmoLT7tsHO
uJVTuSEAAlDsqrM8hMp3UGMmnBXOQWETKlNp1Xz4cICMIwzTYe+aP1P9M+rMrVAzKCM1p4PZm/ua
iZQ2uRCzx1thjYj/MInyJ/J5c78v0eqJh5BY4hj9yviAmdz1CsF68UIxxaEMNDXjhZ7ydBOGLpWL
5s76mxLuLtnHSxbeJ1vV2sSx74VTZ8pLxDJE8vAu+5lRHJWeS1LxBgBdf8jNtcCEf5RPwRFlwOHb
POb/GFm3BDRUAyoHauAHDz/bu6oVx3tLhaBf+OvJsfNEXvLGC8wqECH7ZDksmJ5QMmllrYTKGXaZ
nXmi9WiOV0cOs3MpX0c+XJuJe1KeROYfvOqZNbxVcYXHwwGZ2MknV3cywrQUOACa9vexKehVN/if
a9XO6fwT8WbK9ScWcq6mfKDPYXyOYX7oMDO3J3i2wXQB0uTuIrp1tnwwFI74IEzy8VR+vqRwtW+F
5FWKQ2+YiNPxSDynvQYk2AspusKZOqU4GgUvcvlRFFdsx61EWTEob1jyop2fI0ZkIu0YJWxT798M
guPbvDYnWXrlD5DGhv5g6sLU3JUpZaRSqD1/SkwVwX2Kr9fjqRSFS7KsSv39/p0ATfTdEYspvMCz
p+Kv7MtQrWKUjuIvvALhDaiy8gxW5YACjvraRXZ3JUqMGTNvuOyFDCIRbBVZycCBs+N7/ep1rRfN
LIfQVIJkQv3RRR972wn+kAG8460vVxAx+6/HYI8YshpzxfpEaEDTuE4LA8gFG29S8xF9RmovwXGK
RQ7Kq4xJcEC9wYxUqDYGt+18ZzhzfJpjg9pKKLf/Dmdd5YALSF8UVOOofnDDXd05raq5HeH5zLc4
9V+nMWPP/uYFeioxKp5mdbHydU3O/HhB1J3HsNUIhz469esV6e9R2NzDTBkdqNaDTwxPQ1/fZ+9K
YGTHkmMG/pvPhlh7YP5g3gfpnNA53JpHwCYLtxRn+PWcWuRkKTiAyG2IOQvWI6rqi0h/LKC3MKLX
9g/6ILHECvQ4iVXhmfUJF1jJIebE+w9UiQ/pM4cjFgsCdjWZVralAxZa61Cd40ftWpKB2JYNNLtb
fBkRA+eEYNLxMTt7zPeRX+0w6bk1Ezv0nounrmZqK10whrbRI+SIu6a76w/c8eRCAdypOaxptRtg
M5auKUQ/dHCzL2AN5wmC3Op3CJcx8GL3EONzK5RcOF1PFCC3LgkqX+0cIAweGWSvPBUsGcEas6L6
qWL3YzjPsJD7Fe/AX0cIgC1Y/NMiX/D2/ODCYv7DQkUsNaEXtPrmnc+k4nXKV8naSkTXfTGWnm6A
+IbllrtJH/chNrSMAxixAhzXA15RmVUbLiOB52QbaTGbFLiwyEIOiHWz312UTonMp8bzUsIM2OMK
6mANhd8wMtMO1i3XGYqB0dbSux2gt4fjve/v7KY8e101N8sgUddu+zz/a+7f9IUSAuKI7TkUtDRb
je/9VEIm9tVahX7ipLJv/QQGkIuQycIsVfRIGF1AoZsvY8/wbRejHCKAWGUiVQFxi30Z8rXt822L
CzNhwbSlOBBOjLTTwXKJuAKb0h+Fmf/NFIhKUWzn7Ne81rwc8iqIUWWvhx8yb5p/8snjNBik9WOG
ce3K+b8/N1gxe1BUj3mopWYuOSrAj5JWiLUo3U6Pm4A2GLXjWbnxCvzXbSJUu8VIw74qu/jrVrDA
7ECU4maj71wdJ2rwr8To9mX00re+5wKA8XoV4cNBNo3ODssekk/zptvKoCM+o95X2iMzlwrU28AJ
7qE5eCnD7Q5W7CiYWfRvuyXaP2lnOEOht3lTT43iWmzpPpGzMo3oJVDZt3vVgDVR36UnXtfJCDUB
XwOeyqxKoDjDyfKPdUuVxG4KLBnyhU0AOFnxXr+NgIvQOZtBiIcnPmhxVehsB+p/D/SRk7zPTzm3
eWqZ/Psu2H47iiKOxtVE9Z6O3flocbuNTuZb3qSudYySpRmVfSZdOofV9mjXDDAscBAesdMe7A0i
vlC2415JJycfQioeZwxeXJ5xsRw1IVg1KgrKHuJBnUx0J1g4n80U4M3X87oJApCOgQu4kfWqigci
iSd065JxeUhTcWwiIyDjRljvdDOXIXgYbhJofK5WA3rY6yzSVOVHwdC4IhHCkYySC8YxtIEo4e01
I1jr1nnX30J0leUOxApd//2OBy9jCWXLL+w04hAXO3+zX0LM4YrG7ohU3uxclEALNmAipyyuMCcH
CYFvyaAPWE+nLYFxy9REz1dajXtF8afkNeVuoRxEMcHtjKDybCsnerkBzzCNoL63WpOLRXw3c8HW
HkwWTx/ZRgV0PvZ3U3E35bKXob6N0FPUxHAw7HBsCBWnE5bZWZGoCsCE0nRvQygOduepQLK2+QBJ
GBK6VjwADAn4bbSDdmUjZUDNdmIhw3VjBERG1lAJHNtU7cFQeiL7cbS/9kPT0xb4qTX8pwfZKrdH
WUAssYgk+IhGefW2YPcO0ZgkwtrAcfMDCVpqe5EiZdYIiut1V7pvpvOfP3vFjAgkAiywzisr9Xkx
JlK191+xGqfO7NGHYXmoanW4Kt4DEJdScYVKTZVgxApfuwyA83s4mpC2s9QwJyxnJ0fiIk+lXBKM
EikhKhmoccBBNmwQiCoGkZTV8+TxnWqCqcBBmiE9eYqGyxzbA9/yntJ6qsv9s0bRbbWCEWvsPQXh
npds3DPJvhqyAkUDa4he5YwJVSdCXUi0TERjk8KnE0DrakOhGHrkg3P0Of0G/DLGw5odp/6u0xl+
TK6xH52rdXzCfQfIWGziVhNnEMjgEFKH5xKPN+qJk21sXCmGWdXkZxQMvfpoFE739Jja4IiEJ48U
92HtEkBIs6RN/MqYGUlcmzuWnkLbS4+rr+04Zte25YFzKMrHfSAgOKkKduSpFfmStd80At4LDPJV
nGuGmyQI2O481BPCLjKIc54t3rpYUi+WtLaUtoU4LGPieHicSohhdcAoyb/kHcpcn2Xxgv/ofDtt
BE1vAsVvLCecSq8QWGTb3o4FyPjhIrUqjYozY01AbxVOAl+9KGrT9b+zCZgLv5fe7fowmtWvRe3e
0jBJ+FVshb/zxjLdds1IQJhrgt+ejFYzflA7swGvoIcgZLts57lWfaz3LSHyu3OGHnQkcpPDHbpM
JORdWEGwCWl1scdYllZHqu9FHh1mHAHGxrH43XErxYrsziZChxuCsO/bukubt7HrhsTxjMMNodIr
W0+kQLh3zjueOED767goyMiM7zRmuuf2/4GO7QTL3rqdnkAIeHXl8AKt0AqIr8vnAQDa8dqRi2nl
PBHKJOUnNu+zyZpsaHVBeiErJ2SdEyPERaYkQUX3qlBowQLO86hnGzH19esdQzOcKUj7acz/coW6
WFnfQQl7BTJckVKw5H+NIFqCOadVZu2/QA675qh6OCJtnL/T5/YbVT+3foKEClmpP1dHyE8pqCMn
FyRn3R//fv9hy+rTBFqdLMEqw+dgE59G5HTql9Y3C8cXK0t5vEqRqPj1FvE3aCf4xc/R8AIdxJ9v
yP8kfXXFwJykVLgJxQ6h1AulSMQonWd3XnIIYmgmS3IqZVeNSeKn++HEcOHyM4TjPcbRlwwK+bKY
S2LyjXMYKwN4xd7tiqDygDz1jrHwOAubeB78gierhjoawKJfO56Oaqk8XPbLxH2C9aUJVNPytjMm
TVSsyAl/Zt1utuNQva4QVnOONOQxjkKXqDn8lKWWVIt2JR915593FjEpEscxpxfRVPodYSF30xV6
0Kavg85YaMmq+lcpgBDA8JQtJEcVQTGLcWhb+kVaAq76wpcCk0Jrcj8QnzHiTLvJa/9l7NucZOwK
0btOwBxbY/kdLd4MrnzKemGjVA1gvVxU3xeR81xLNsJqIi2Xy9Xd7bwxgd91blCeynPU3QzYYTtC
QcNcIR0Qju+YuJpgHnD5v7TyEtZijRnXew10JYXCnQxSKQ5kQGpofGa0+Et0bK79ObPsjdy5EzAL
V4U8AdsJ5M0dolpQqAnpwIrhfQ8Yep0qq6RWrf4acDnP6lBizhAM5afPVpsYlf20j6FGQWN0H9ky
k4cmMiM6YQ0ynQb+3Jjuen7/taqjXHRjrajthjgFviL4hfR4yQqD/daxlVAwqJn5txj3R7Ymuqmj
BcHnmzuy4c/s+uJauVqnr3jyrI7a4oCkL+14fRjU0dvOkskNwTGUxrHhYMZBTLT8Bu6p3D61YPUv
JSMfnwHtvCKJN3ih7plavYKHTMtyyS3yArXp2oopvQDQMdAm34mV+7OZmDtEhG3q4CmzudLLctW7
g6x3O7L1PUj3EVaSFOGb653FYLLuEjz/3HuzbqIHxf1pLQgDWEMIsv3SoEumRv0rCHeRYWjc+9L9
T9S+ulrOE9jxdcFeky4HRrcS5zbEhH+GiMhnCRdItlzpQF1Tkp0Hnaun9jC2VhwFFQvUS/42UGH0
bBCUhb3baP/Qk5DKz1EkVRWKF26L5rDz/W2jndMZlnZ52kpwMRmBantBprjl1AELPPEtbtqHnnOE
DCq/qB2bB+qbnVYQee/XVrq9rURUUYpJDOlhnMryHq52kxBlC19VCLCvKPxEj8gtP/WSBOi64Ng5
L44OO6LY8Tr8bp5NANJy/JY1cC6ulAlOyt5p90FLxDPEXa2gt1InLGI07pZmVAeS8lG6sN/4fIRD
D405d+/QLliyhIRVNQWDR9Ose603yPeT0UQJ1V1fjIuBqu0xw6tKkHA4KFHVzPHNt0Z5Ro/fnFq9
ln6xn0UhbXqF991A8VKgeMllyXWk48IbOJmzct/JFlojwFV0WM0IlG4WhPEN+PvvyKUKhw1vYi49
gpx4MrebUCEABKTWetHHzGnq67rewDi1KKa9pQaoJE5PysuNUUMvQ1K5kB4iJR0EED0IQ3Bnh2BR
YJrVz5HbnZeZeEoDZpgfZSmLcNpu12zskl3XZgELYcexGLQQCpD1pU0qBsH8KcuV3+Sd8pjBTSCn
tfxOKalnFX9zaN/YNJlL959kCmMc27+4bxEp8is1Q/q9RcmpKqPMZQ9iBlpxJyq9/u0GfbKuxzzD
JX4rVCjyHx//MBzRR35kmoXan9eYAM6p+V28cI2H2ff3TX7/PU7z+MltxbQcm1sXoPG8nq14XDK7
xuO+jSlCKB1n78nr28eZNDjxgYRd9KhfiJmKunHuqFSLqibuuhfFRBRwBuuyGbcnGBWWDJnn5JX/
kIRambSrf/lQdha3HGHZmIUqRytlDf2l+maTm/tD9YCpoFwgbHKlznnekVKX+JF7FQwNA5T2o5T6
Hze1lfO1lrti1HjAQZJivtgMaH7Tfi8iyypavjQ6ZofOnx6pK2wv7qXTVHymbmAKcT8BFsCUqy1M
dmxomc3uf1pbUGIu17gxk2tAgvU5Cl5YNYuIN8Ov6avhF77QZOFmeS9eVQ+8urMWvLNQaqthC1oP
H/NTDKINPZDKjTsnJ2rBHhrUqSgNuQmlDkwnTMbs8EX/bBVzuIhpa5n8rHJSpHLvmpFkP0PJHDLC
d1in9ma8sMHtBOiVXxlTOsywzuNX/N7/77Lo2UK9uo5mG+/MtNUNq5hVYbMpm5ywCY3IQgeHg5In
1sJpFwz5lejihMqpmCTPoq4ojm7e69B9gOxzPuwtau5Y/p+msAItYqBKUj2U9uWPAS1LZtvaadsg
lnPGDQ3dP0vL4oNOIG/mSaMKCMIguLvw0JHLmqWuvVlnlBONxZa0luwJmyFEfQAI3NuL1ASCNRA6
jcSykBsKMOPFGwUX3vLr92EPMNxpJvDsxv9W1b2I2M8l4l9db/XY5v1tHbA+J88a261CX+iTOpIN
wHruOstBmiCrD0uTYh3xECTxd/t4twU/+DNYdm+9pNefEtxfATzp8TCerpR4/vUpj+wD5wxRnHVP
vZglGadm77JexAz9+lAi+e0ZkxreEkafq/ol49cXwN26AoFXjYYtxio2PcyOaTBsinSeyGp1T7FR
F7rve9jWw2Bq/ydcz6Iy4tEJiyGWVowffeajsBVHX+AGNl6qxkUoYgSPeCqkPZOdk4nRXzWfIiHb
SaPqOecz30GcHlCZwVrDkZZAmriezc7vcomRMtJoYynjBVkJqK2pOq6N6ZFrfq1Hr9IV4eGFX+9H
2pbKdrw7rmbR5p8mlU/bs/U0RBdidiLKah/Xk+S4Pm2rbshaCNrL3uM2gYgCN1rVWdPi5f2vT6pO
C1ub8ko8R+bKFOtKGadOaFVKlvmOvGLa4gdqcRdtx+qmfx5LWTlIZM2XZx7DPgJ6j4ax40jjjvUp
2zAKOsP4IsMEkh333OdRuv8hCUZPhmV70HzrELVeCY7Fjgzow8uzi5i9otzV6mKuwFqyPVDsMEEc
aR4BuJaZy5eimfjmyD4T8F6twysLbGVf/T7M7b8kjS3/LNzdjGyqg1YxtIV8hHz3+sB4e2l15mtd
YbH+/53dwgaNdsW06tdEXkap5GUl9tVC6yxC+7TDuEUTUPt0O7IN565e/1JR3ckXMyluNLi9LJug
dyRLa6PKTzktucvh0LY0YpWggEXA982YQaiq/XMNp9Eg4OQYG6q0GUU0amDHC5udUDCig1M7w4yI
gH+jbqFoXyQPkF0gjA6af/J8T4F7n5vak3C2AVFaSOuqCFXC8+VHwQ56sJIUoqqG0VqoCSndnv2K
3PwokCWRHsH6R7Rt436rQlOEdYQTKDlHNx0lFwGYdGsTd/OCPUMC1NcA8q9rHbXfkrM65G2ehTcK
2aCdCsyeg2l8qLjNycvIEshSiAf5in4wLzNKsPmtkD8uA/5LB6AjVCmyYFD0HolkUTQDJZnKEJQi
g4Vsbv6pKIKcjH7axzyBFWbfHnI9Bwia7i7V6snJXf/OsvhDgtTd4t6y8+6yTv3rH8XRvJ5N7+l5
xQlEFOqDmboDUq88aY0EEmHA4fwYWCITdGwN2DiPSIHrDLZio9b2fuk7Ek3AIXwYvqBHoXZqXVJP
2MpPUOY8o9M1ZUZVSdhnbCyCxVeGA9ehfU/wdNJ+fjdMRvjQeFyZLYE3YefLdERW0btW6SbWj85A
1GcIZnvxG4qUW4td2a8kyaaDZe0l2r9CrApFINzSpY/ArMmt4f2QGwjfzeSyeCC5D1d+2pN/qsO2
IP911yxQplh9s91CDbVSYgjswiVm7973PBALypUJHlsTopBGtlcgjlBVTXWMAJsLap4KH76fH9Nl
lPDDD/Kzh6j5MuNe+Gu99YjjcLLVpwa56JotTWRG0/Goqsj6n4XXvleZtMYILq6j3R5FxgVWD58n
wgC7sBukhjOEclVqwWMJLZGOS8SiMcXYrCVVYpJrEOdUrKwjmttcqO1y7YCN/vv84QH069fM+x3Q
c5l/cJz/6Em5Qw/NifEUDXBbPEOzTnTaMNgQqxfnXdHXVkACC71tWa6LCK62eBrq6ogfhZdysf+J
6Q1naKvfVuCnfuwaQ/mpaGfTdHdSqYDLwtssP/fZ5ZRiAyiee7Cs+9RkgSKpZjYJHUxhh60hVP6Z
kpRJvr5/WJflCwAjxyMBlAFzaa7MH4WsZOBlkwzqUDTWnga3z9iWOzhIEWACmm7Jtq8CT2+/bVZ7
fZ/2UFKTTyRni6K+i1s5WjEN7lcEJeuf+U8fzVbBJQAXQSTO5cRZUthI0s4Vch6MDHApgRk0x4Hm
75XTzNkFdElTtP1DQMNpTuyzzy6Qn8Wwjg0Zmd0br67julFIc4l/MHMXu4S81H4ZEjL/QSYTQcag
cYxU4llO/g25/PiubiJE7jex6zY5WLIgTagpbrpw1DXMgr5F8krhdjSjd3l7qiSDyP/umtHwfOTG
fVqYuSWeOrSCVjM9Bhdjl6tKPDiFydKkhlthd70SxWpfzNqb7wjuXNf5O0Uua8MSJqb1zH4bcmIA
2IvoacrEKhXI8I+kuZKreRS99Wt9umwR7cNFjHjXvSbAYENk+NLK6aZYumj0VUHyBjJApITkmpCI
LIj252+yJn1ysdJ/JMSdvBLnnN+Qnxn0KR90SvFJ4sqHVtulrqWlTBS4LT0QlJ9bSBsXnQ/F/O5Z
p3nKu2XD7mgFRkgGqrXEYUeetbvJBUUywRZvMJUQmlRp05hyxIvdHdIr7dR5TakuDGG6iqwlQXC0
qeRKHbK43WENIdHpaZLSIGFfJaZOmQuUb7rRSgoSbc/GLX+z/WpeY9BGn2lLfVflWKwZIigj1Jyr
58psqQFZIqujyyHUSh7HDxh6jUSuVs/4NHY8P5XKIIpsF3eHK15l0yG0irSa+XxhjG6vJGmAJbWR
eog44kRkSsCx3z5cSHKI1K0Xrh2d6mRPME8lQOx1KEE0d3oKOnAXX0B6cSp6hh9cqj7k1O8E5fxO
bvxMTce504+gocfbSwPzZrObGpBLeplYu83vx+zC3mk19HMJi7ejj88x3lhFeOIhe8HdWUtf4Heu
GytM7JZRC7b0IKdZIeOhKjdRxTE5e8R6KlTca2qlt68ikvNhPt4dW6tb4JDz8LbqsAcBB1N5VqG9
niQonPtsK1J0cv+Eds7D+7OfZFoF6UbrRgu1+HBWG6cRb+3MnQALHmDTseW0xLN/keiMpj2/b+Iy
R9FkFQ6VTSlqH47N+l902OfGjFLtC+DKFPxSW6D0gpCj7MlDpGHI5M8aIF+/EczIPeZt/Oiqfhqm
OuluTgeX7VlnSrYsjulLnrG+XqgGu5t5HZyKmW/MsvdgOi5ip5a0kKJnAhcyAPmuN3q31C6/pxql
HwbSSBAw51mCtm3titU3A2owfLFb4ag2/S/e29eZRvDwjINou8GfvXN9Xj7n4teIM7jYvTZIRIpr
ma7hBm2pwUWMzZuFhVFVweHYmwd/a6vxeu9rm1ymL4njfpZYQ7USd0LXiuM5QamzhNNuzXrzJjik
zrbvtaKLa3hPqrbqig6+d+lAqPy59V8imMhXOodvvRquUN7GVeVffJpjC9jA9G7zfWnIwNig0dHX
IxezCh9MEfFmpl0Q9qE5eGqkSvqDU9JNf5V6sNell3Ji/DhYzm8FSihY4XBFrkAUcY4LHSTnMDYa
nZQ+z+T0SgQRx4g064iS55RG/qlXti2To4j0frBwMLW6yWYYy6iWouTdy6lvD2xeqfjUCDYNggny
sTQCyDXnNvCw7Spr9zrH333xgjaRPnmsT2Uexf+QZjrMWsBxjLutoUfPzmf8BLoDR3NiKhvDSwjP
Ph+ebd1fRnU8ocjf3HU4wB3nwBDiPzfjxoW3RF9lQnsN49vwftyM8vBDCKzzEYqcvdMZhtVP9dB6
uWXJqvAO4WQ1KxUInG5hm662lfW58CxXXFantVcO8idCNl9+eTzsC5RXaGQRV+E31wW+wMDUFwsy
Q4lXUAmzDT9ryBO5voH/mVJSGLtod9G2bYpkLZO2Nt3hcSDaeM1JPIQZrs2S407w7wrDZ0sgacHm
43vfWCVYorMdWjPdfpU3j4vr5IrkaW9CJ6q6fJbgbhN8Eo1PUzsvndYj3XShE+WtCUNN27oNmKOY
wVXS/1THlw0HzcwGH3KzrFtbcjV69D5qWOotfhQXObJlY9X8Cxw19fRwky9GmEbb7vHvkrRl5oYJ
3vMGvf+HKRk3KQM36+NFbfiZSEyQRAAmLuIq6PKNGthUCH0aOiFLpwADOAIED/zhbdYUv4oQRlaP
6NCsLeVBa5Gt+XMBwjp2L5BLUyg2eQPbX4yPOZojEugQ8VjZajs1TfYxRNud89m8kRdnW+dtngYj
txjnCbGmmqLcMe1rfmuDNsk8qvh9GRWJnz2kOAptrYR+bLoHKFBNdQXdMsMR/GRd02oxFcmchmUh
Ri+7fW1VcD8s8hxFR41LlobnfATDxunpd62HTVYUsyKCQAmt3pCtau52H4ClUnTYnHg9bN3U29yR
g9fKzP/xaFzUzdIvsbA3m0YRNuzaOm8biQrPoqtme5/U0M5oLbPaiarcqLiIpGCHdvVBPqFrPO0z
T4p01w+VvbaAKpIZYQK31WbZhm6UTgGhYw7sr5ltzH8qczNb5SGp4fOQdG/fgyicL9nUAV1BbVKD
nF9NBRN1LgnyXSYgzQxkaWA4DleQF2+mETwbm/Nuq+USVmAzkyILRZ2lot0Er4xX7d3i7N1X0pZN
ei1sKT1SJSJA0+K96k+yvuK/12ZzPP0MaQII19kKb2P6oWsHysRAdaPCZXMZkti+miFSMDEzxWX8
/V+8XpJUocEsDQEd3wG2zSt1B5vdZab2Zeyh6TgC1darxhkaf0QoEr3jYJyPyAQhqfcQA6Cae+ch
MYSeego8O/M9XqiDuYCrJqw6rCnrRrmj4Q1Y7+63cr8x1e0+Nki5ThUrDlDFfZWtG5Ejk/25gvwG
RElqsetflX2wYSeOxj42yqF083m0JhCl0qnKgRX4fNkzMkT/Je75bhzz0hzdb7Lmzy1FPFgUzAwN
NFwMnXxG9sRVNxtAENh9wer4AE1dFBwCd0cA6CVkA6PyU5cAS2efAUTPB6Z/JOWLAUXPwdJeSIm0
2QtTF4zCtB4lc1mqlAwIgsm/ShkhjkztoNmLNrjpYf/b5tEeIx4blCIswTv5lPj4xk5e17MA9s/Y
ucjdLp1H7T0vb2ezh+v8nB9ziF7FkfvTtvt1x50otb9Jx8LUrpZtQ7P1xgfYlHVAOO2UBhK0saWC
fBUTdHjNUWeiOR3z6kEbr6YQhkhWkMA5JB1YUx4naxaavGUDq78Gr5lcuSEkA1O/OD9mm5eB01N0
DPanb4f/Xw8V/x3pPFIQ0rjh9hBw+BbBaT2zqyDkPew+xze8OdtYQQlilQf9DbbhCL/kbOXxL9n2
xfFVR/cyVVP5be0sZ6SDbb1fbG/6DfcaizmwAMDSJpOS4+pqBi50ipqgEuJdwt9FzSqlakBYvJJa
yvDLbcJ1G55SoM1SHU8WCdCQuTugxU4u7dTNvFQEf6eDP858o+IA0UVvOYrSbX9ss2wBDWpGQqLA
LbG36jJnrXld8Mb4WYKUUA1U7rr4SP+kSlhOfNi82eFVIOibw8z2AHB+jAkHH0dnakV+FNDL01th
IJ6nt6ubwrgTwA7wwRisWNMykPhUDnyeiutzqD5sAoH/82z3FRr3ysCE+idiMGOLoBx4hWKjVI0J
uY6rzw0WKkPGBWT0aubSMH6Ld6hJ3M6OWmO9xXVlxpxGOSCiXYZkHcrYLVNJHySieo2zVZdg7AlA
ecsAaF/Vvh5YVLIdmekD4tHC45SsfOpjfch5yX3gbl1E3XZtlKjc95X5svy/v/UV9OBNYQecjfvM
fU0kZZreVzKTCBcotoNn/vUS9oRGTM3XfXP9T5/3lMSnjvCFJgvb+wpZaMN7Ji+lqI+FA2Kwt5mO
xW9budiPdM2zHAVlgdRZ+KQfAu8rx6u9cTAs34CmH4EoicfGDcxw+MMm+W2AF4kd1LrgUpv4ANSe
fmXhojJyGhKygnr23FmEXp4Lyq9NWfQMJGELsi6JQf5BzCdlUGoZhJ9VbVNOizyOr559k9sDiYQ9
FiE5C9C9NroqpOy9i1Yw77piTBp86+RP6kK7DKnqCLz7ytuxu6RtBi6tmq2d0HgUjqDzNP84C/CD
cgnueF++zlxajRnPNSCO+3U63HP24/6udNikS5fHzyVZOLXkuH0IbmdAGKwjQnLylvi+uuKpNTdt
KwXCGsPFVNxOjHPxhah6aUXBwOUIBMoBzSq9MD8v9pSHl78wBJ/l/3ISXK3DGBbctcTYgesdSRdy
3ydrFNDA0CYlupoQcUI6WVxz/lCL5P5QN7F8ZBVbuSc82LculZJTHv8JILzBxl4fyUFmjwMw5w0l
s/BbwyhDtwCTKq1B1ihj4Lmtv3NF2ZX/WySBjWslY/elrRDwjGCrPNCf5kdIDvyGTLEcWTdjg46I
diRNgvZLdZc77CkOrYYPO1dSjHyuT1M2IMx2m5cts2+Tpv865e+CODIpecqUHE0t2ofO0gQ1HcDK
mo2vO62REgymsEp4fLZOSPDch/OqRGzUzqGrXxMbuG8zqyoQPMeowQHpxJkJZR6Br1JvuBZKUSYA
Vr6AUcznq1+3RTTvYYEWhw8rjjlZCndlEDdboXbM6pa6+4IfG2KszYa0fBN0bEmZEuFYIjV6OTkv
FmU5BUMqWD5mA99tN4g0zeJZepcqjE8fHLGovlV1EvBVxbf4azbh4+c0x4DsO1bFpBmc+Jm+DGNh
wf9yI4LtPV5anFEt2cdRtcXp/rhFqM0mvSTof5Sjd/y/hrpC2QvWBuXTWQ/VqLDDEhENPMSE9YhN
BerSAhiYHBsI2HqZa9LHYz13UIvSUEtwMoGWtf1XEyHj9v7zGvRncjs2GXeo919PKgwkHT+L33wp
Jph0DGGYJHNP0Vn4giVu3fc2mJv1gItBjJheKR167fDCvt9vNn/HlGcNPdwGl6+rvXv+ezw9b6cF
ymi/LZ6sBz8by7B3ivHv8notTsMgGKY3sPLXwbd2af1WEnJJ1VIU48023YaATaAB74cKCgEo0CuF
ka7/y4lCKbZJTbr/c2k+lE0lc6bGx03CXS/wot1GyJwtRwXRuVpf2BblP/GcwowR29MhFhCMLxQq
cqfl4IkHJojreoH7XCgVU0Cf3OOlrwd7Y8JWeddUFRL9miYQvptjEtDN1BZAGaVHvDlxR+QFztC/
7oJRRzb2vwKvsi2hrnF95nwhBAqfNCYFEeQsOVqfH4vCx9vMTEZFP4ZbmIvr4mPEWRFu446/BkRi
jEejgIl5AMvYdKKINzQkS889ALbRhM5y0w9peDGVCr1bL3fIDMeLLzPOgE+rLCw0B7ZcWzfz/aUd
2bTU+gV3AtK9quitZJxHh7duc8zslrQUUNSHwhaD1QlBWX7brNPbJgn6xPJ/ZJjj6gQMgH8wVEx2
Ikuejo9gW8lOuKSrma2XeBKTB8LdJSU/J1kn+4+0WCrf6Q7bcwQ9Qs5dycFgwAtzvMFjhIlNWhSV
0euzrbMVGuHcBzkp5+QDXyIht+1IiOXrnQq4cKnHIjZdlvBA20JHjAAt7UY7mpoZUevMwqRVt6+I
WA8JHMR9bpUWmjxut/en8AfdGgd9BKk8IwTbpdu/+1ENkN8Nb48mfM3O6tZAdA4LnoxeNgg1d1Dd
T+PjiVGUkc4N5yM3Tj/4DNwOEwiy2ccPYmFLuYhpwO3prhNBPEp/dVLUWruUkvyzMmtwIZ9aGrim
51b3maXuwl0e+jL7cm+9FmK7Rw4JJze0Q9WC7hI3jHS6+w7ooJnE+PCDCaYy3RRoq/rHANNu9Lv6
lPzHuIzUtHR4iMqRshe4sewt9EnYMGJAolLKQ0bmFbq4iuaJud3iK7H5A7rcoZLhNUJBUlDKK1i0
gXIQP33K3sHIWzy0eYQXIGurlj+ojamRUGlZ2txyxGfZQmI5VfB/d0C1ZHPI+D3Tcq/3TGslgGtT
9cwbw13niozCblzOBxopsXfByaOZxrcMDVjDHvh8KbdQpZirGFkMoTTCYVJc1MIhJRtcXB1dSpzb
6fbnvup0RlBzeC+oMDdzZUZCtk0LQAY7dYlYXow4M21x3xbCKDG7kFSpakXOHtc9+lKHatJbAuLx
jpJjPT1rk3q0wOnHbBemG3Q5MnOkEEP+VIdz40coaAs+jAUAiDB01VBZcv9tk+Nqcn3VGcocEtys
cgZxSdB27CaxPc26DyL5hoq14ThGdm8hWGMof8zJH/lp0gUUkP9wZ+wxv/sC4rm2B3oy72GxCpag
VkpqzDdKuemVh9TgjJbwWGU73z83BWZvFmNgMEhZn7RAXd4dBWhKZsPj3+FRr1ShwwTCGpW0Jphk
d9u7X4e9lUzqM3or9HfITdwMwG4ndSA/cNxZE5z0rQqrqTOu08k1/3K1NdzCHfcbpDuwMt48nthp
yxG0VxXqKx3ELGci2o5gh8XmQL0tct0oisfAOXlhF1bhJlYwkOjgT+rD0Z3c090UBqeAgkMpJC/i
KAxigGKT6OmMEPBb0hwKwZSjO3XqIB8frZTHrK1sYmjr97p969VUDH9KyP2Co187UWjBSJjGRGJO
f/fJg4Sk38vQfOwmkLBnrpw6AARgDNtFiKSPiXgFYnTSEQkVPWVPwoUJZi07bMsLnhZZyCevjZ2d
Z7jLGV67pBO/4I2nI5c7PmDGV816pu3NgsDl4oUY5+2qKJ7CUn1wrVBOhxaDLyKP5t0B4lNdr4+8
UXm9yQIq0YZxX8eUwPh+9Rw3RKQngC7oZV0Fen2x9CNba+4HFuLvWtR7Dg257RRZBzMc+T9rXajH
M6PCKeB3k7pc4UChJMD/gclAG6BpPl1DCufuIqxBg8E7fsGBy5x9MzfrY1KX+xMZHCZyaxzUbPHc
UHTfLJqAg/CiIzGQ9n+hOwQGBrtj1zi27BjBz6BirQjfyaC6CuoLmCQc1+7oUNGr9PQTd1NbJgK/
XVCGrdCVqAhyg6VEudmYs6wgrPUzejtKv6fXvh7KGbqVT1H1h4z40UhE4pwFo616TUQti7Hwz7tr
xUN5GfoXCvSqoXW4AQoHADCnaNap8t6sGkBvIXoU0n5p9pv5AcmJDgO3O2CXOtgJwrVT9wbCYxVp
JVUN5VdOv1LDaK9r8n1qvzxxok8XyWSAyWVBOz/oPb0Dx8Wi7fy2EE8deFBdrAyuODJ7bt7ie6nP
py12FHbh1s3dT1l7zx0RS+W4+DX64WY9rMeZFMRsQVzjPoyxCVtvFRl0AKZhB1Qe3kub/SKZ87jW
QVtkxojinds9E9reQ7SDLIxZ7MUgmH/8A8O+ydKBkCOa5zev12SZW2I3sdVUmfg9NKAPcQb0VIep
AwI4d4M3NEiElwrFiwG0P8COJYERW8iHXRg79kVhKKDmkgQP6ThufQMfzEqS5dl3KOcIc3Zh0z5u
WjKQRoRl9japcZVRvWvv+ZOJGiCIRp/Jy6/kKRFXosOFVmaCSNVYNdhLfr6eBTHrl4OaWBxUsJlr
qKFnP1ldNf4bYZ9XBgrXuUb7jZ5QQ94bjY7zEzZ2qhYCFXOK+F2ktsINQDAlgX9dpkcmIRF+MEry
STPtOw1vl3V+qb/GufnsV5mgPdz7Mvf7Htv4CZlMTVL+lTm+WuR18mMQBQ/heVUWL22qb4uFbo+p
2igSAsyAHxIaEIr8aSRf+58ZqGNgpt0iuELhUKHtwWVPtylnYcsf8tkUvfMCF9QtL3F7dD/XlToj
NIbmTtvmBbrynqT93/Fp5WITzeGAFAY3+EyoGNa7CQvFnTneOveNUJS40kk05eA2VgTMktHaYEAQ
70Y40PjuB84YyJGQwOILwSQRI6k74T4G3iAg6gIJ3nK6PCuf7HmOwzigSAvhIpHIyTwOQqF/iRow
eg3MpBG1Nm4yOS50ITlbIm1oZrCGZK18Yq6nQR6ykXV5ehP870S02iPRHYHifAtWzk53A4WzvMcg
k6z0Midge9GBczBsEU3WrYJdk1UgrlmOvbvb07A93XNWk6xvNCfRmONvpISZVZVDa10kZzjUue4Q
wIbska9cSDUO51uwqtftBHKH4ygCbKTXz+Jxwei1KBVCnNMr6/jqe7bkl2RHyOdLmrrY3IvPXS8q
dsVB9joiCZefCaTS1zUsWszdigtNAUjvq2jiFxQpumCr7xfDAg9Vf18eDVh4jDoai/pK3nwuQy4/
SYgWYFCQO/1BEVoYyM9/mCsEDynhg7CXcJ4W1i+sIAjvEmQMrmLwjNGJnPgRF0emPKPwL1AKF7ib
T4YdRxEhamJLwl7jGIGF3i5717m5eoWM9ZSZv0LJwY2kYg1FXQ1xEzrzWp5U4hOFfGzlJP4G1SrO
dvx2qwRUEWo4rAR+Oznumg9dcAVqvQdeCDZmAk3vELlRH8U6tOvFq1XBZ9zHH0LW9ugGInPgnYfD
m9YKkAnpYIxv/6iI+SyUyEeZqt2rrudvlW3k3U6mLjf771mCNhcUDPMMeTdNljUq+4YP+DVO4hhf
jFWbOspIkCExEoThp3eVrqW2XZzepbs4on630Wjg5I+sX9u7NL2YOAu1O1kNFWnT2QOx2TZdWc7/
dDgh4oIwcMeRFAZJhmpvnmwf8Ml1i5GRll/peB1lsd0r1rnRU4iIeZP8aApwm3KqnwFi8azNALdD
lLy38+0d1aJeJEZaM5dKoqC6+ohP5JS9Gn2J5sVxG+G6Uwvh3DQWn96zi8zDkAf54Y1cjgDW4vlN
Spfy39Uhq1tqs7NKitAhp1hR00Ym7q0dpgC1uyMCBL/Vx4FXApJqEnQK87X/vN1LDnYLB+ol55AM
p1vJcUN7D3Ni56LedqYLS+WaJTEOa1tNvPuLrjfmN7g1lK5PaOjYbR8yEiDQzwvGRdhoxNRR02Fa
JZENHyUS+uCcIz7VARiqxEBibju2wCwAJ/2S7/f6fZMPpVuXG74S6XuJtE/M0SZQFkfbt+uuNy5m
ZYHGEYsTXrGkI57FWL4cek1CVsa4Hvxtv+t6KxQTDgJ1J1HrFEuOlnXSYASxrtF1lVinfOhq7Y2S
EPOXPtGtNY43RVHk68AMpgypVQ1MRjzmwygPEl33XVH6UgIec5HhPp9crSMrHAWgpDGB5I/cdqbm
O49YMtpvnhqpXHAwsMUeCqGt2fQtAtKnZImqnWpQJVMJ56zQEUvoRBySSgtEUKxtRp+eQ7wa7Y4x
blsD2aNSAeonfQocGMAD51jkQlfweJ4UTAYmCsXBcTIqlskDM+ElFdNKuiB3oAT/8WeKZ+TUytsr
aC4xFsaRUdt5GLBz9220FqrLxSzqsOFIuuvh+qNUBE0EwvOrdVo9JeL7mZ49xS1AQNbVuvHGYwqu
+bnXmjC4A2xC+g+bqYDB8YHo7ZLOaVqUW5qkDVGDGorHthjgqOm1WxDCxs2VsFhY6nlljxUydGWr
wE03s1FK8/xLZmEmqcU0cV+53u0dHinbpd/acYlIVBDorcs4q01db6hmcZz6PaEzMY7LjPKaIvw2
6sezqv/J66cL4WGdNYhW3kAUzCkzxi9J6xSGpLGASvP3o06uMyvXNj1ve81zVA06xmiddgIVTQ32
aGW/WxBeUOPhVafg5KS0FZswupcoTEHX4oxYP98wE9BakYfreuLk+p+6ZFniUBoCb/zwgnVl6P9+
BSxicY+CEyd1ugkk4ZQfOPALTJWqVVJIaakrXrVCSJtiT1sr/QzyZcaPEnGi91IwvQXRF2doRtfT
DDVaGTmVsuyfHnPZv7GpR0SLO30pidHIQrVWGh9YYXOZpqDb00jTaHTO+/hmNzBOCaFF8ZxnXGhm
I9Xy6EKZRSnaM1Qb4EIkHb3eDkhG+Es9uCsKCHI7X1UqRmlk3NYv2/Zo4n8qIG/Y2DOsD8MsvdKV
5N2JH0Bq2TCuORS1mNh9jbxAFYIrchAJbmm5LT0FTN7JlbmZs4JLqHdk7Dz7zhYbfLk+WKTmmwFr
rU9u9uo2iyLS8y2wzfnwZtCboWnenkviK5YZtEFwDcb5QDw7WzWc292leMH3ZZZSuDrdCjWBuXto
mudltroS5fnxhKoHXpTX/RRGNLkVhzasfh32cAVTQZMu5l1EvM4XDNFK06tsptYuThB/9+SkjUmY
n0KpBoHlNMu7/zZmLfT3qwDgVPhVTN+RE0yRQ/cqOhISbC9RVSLRjnd9bmEM1xtf1UuFFtzVFiZy
DzzaP9OzgtUTMxB2lIrHyrpaAQVnIhZQa3dCWpWcwpl8X8yyo0fjpZgCjhiEQfzG6OI7EgA3qU5H
5RAq0m7Td5SX3pjTvhymI+btY7H1hq9ydiEXLWxmrpcGOkTKFJt9mBkhBOgNefPeafQj4Top1rQY
8sEbQRajpz0ArXu7d1WPnOnVbdQl70gdPIh8MaNJUCwKeUju6+xQzUIiS4yzTB2sQ1zty1j4oDf2
brmPxyCDNFUsaLJR3AFhzw5kq3A5rZ13UXfGLAbm4kTsM4/HD0RAC0QksCrKboBc7kTlEbn+1iRx
uElfVjP9rtZ4DWW2aBw4StgRk3vxXcE/qN7ohT3xygQVNKnAt8A31JEkwR7cP+CGXfRdn0cm19Ih
cerBnOzAQUreoq2XAtZC4KzERCAeAa8Q2U0ClT86/YOfeE4X6VhTVQQtVa6xgC4u7GrVWkg11ulI
Hxp3cKH1A4wTU5IKvb/mUe9+Br4bnc7cPyhYUb+hRrJRU06mNczfxljI1EnwqNPbxjiCnQlaJZT8
NP2a417S0l3bXHwQNNXTVSBSrsUg943d7SrbiZLx3Tpw4E/AeFGfE2+CfXW7iBZJ197xUsx9nRCO
trDeMyM4Vcbr9MUueiQDWJVnwrmM5uNxA11ZK35JtHqfV4uWY6mk+us7lzFa5BzSNVthfgCcGHV+
vCFOIXEp4QmgSFefO7G3FN1Ts6idkJQTeQlUteA++11FEQgINao09ruYrnwePi0RHxrd7zy9yxB1
G0UxEsq06SIzh2QgYP7lEPboaMjYFYj3xTVsdVh6hC0AGOOp4MyZ7HmVyqvoTDOrqyKxtXBwG14e
y+Fgn70zcikYaXrfLmm6dBifTh52zdsFU3j7pyQYX55G0U8PUxqIkeWGRXE7KcvivzhAUvNa/TrA
W4rN+hRc1uUAdSbzWnYhUCA1P0Sv4YnCW1Nbe7zlO3/wA6SPdjMw0OLunNfoJEypOABXPkwHsFdn
wk4C0PyrpKak0Hb6+g1ZHqOVL7ytfouYFPjqinu1IyMQdgUQK77P7RY7QgTDLtd+Eps9G2f0Jy+a
OqI56JQ5I1skeKuYOVrfEL+oKq1o0AoUfy1VceOaG40Qo4KIgp5ly3pbtXLQztduxTwrfI/yL7zI
QH4792BHjQ+1zxAsiRLt8VFTyubu/jYWjoFUVsPbRsqx5as26nQmQUxYgJZla7wah3WGewkta8EJ
kRzPND2vCQayK+aMzA2HhLajEpX5wGUTHVB1gUvybEC+ak4JBfkqrm5jkRsYVVcNP+HD1jGu/zLS
lf7RSp8aG+0gESGT/ecYxHtRbYRXfjrzui/5iEsiw2YxapNs+WmAN0nQ+AL2WhB6t0Lduh7sLciO
Qu+SaWoO2NSa5bvZyKI58wOgySH3/csnlIq53R0WoN8IRpeMO3oqDCGG6Uccc/F8ePeK9e3Iln3S
nDkrKjc4UvOYrOHiwIlhF27jLfU5NoV/i5VRAQZ6IxXDJ7GKGcuYz9OMO03qAjJsKlectC4z3m5V
L7QNM6eIdPIK4C4xOiOi2Rz/+2wrxnPtujImKBHNNPz6HqNDsoXUE+8X86cmo6Dx1kJxagHjFOWI
IVPTL3qGw5YGaequ5IdAviozl5KQ7yS0YxcIKhceUMvWiqeAevRE/IIU5KW0NJvtugXTkdQJVhOp
G1cm2Gw2k25gfGZLp/MxUrO6qT2iiaTDiRG/7ymW54FJz6h71X/TSZnofeAu/VfoBb4+K3CSdzOk
TDQBNOto/OWy9u3mWsEHnrMFUc37OLALs+BvBxodfjwo80ZOnLUqYEjH2E5/tlFmu1jmyToGfKSf
Bjp7Rt9IuSB270FG7m5PEDJrIcIuxdHUywE3s6EUJaUQrkhsJTfW7kWgT8mHI/DWpnXmM4nO1Zsd
qxv7q3XekldpfBlJx+rSZnZAdrsyJcHKDKIaOLbwNYAccJqS6QokLB+F3sBvG4HnR3F/8Vu7GWSF
sYambTlJ56gEScWAEYENCQ5qTzGoLFNUDVKMKg5mBswccSIL+AUp1wegKXOjcSBk1c3qep1A/uQ6
9+b/rJLKD1aW53cUgdmlMG7xpAkaKl7no+ZTkjz1JV/Zhy50kgxGHPlmN08ObNaxG9XrWsMIzg9r
hHtnVvHPz+O+FS4CBIgTYRLjQwzCrnZ/NjD/qTHyQDY6QS0hlrt6gTQs31qHt78nwy1y2pV91Kiu
eqiaVicyklWUcWspQLJvAmKykpKRRm1UjVk5tfZt3OStq5CszT8kZwuf1jNGMiOuz3xQWVri0Z1c
aTeTCM/EzKWNPOES5lDGTQhg5nJB7hS543KSaJCQJjlP+O55n68XPSvwYEZrpXT7WN6lqyVQj5K4
rCq7uK3QCNrPuAEkyKyJD5EdDVQpfLRhXFCnHM7Tymnrz1YHmPNGqmxHkf4VA0nnXZ7HdoRBf78k
shv4LKgCHCQm5/DAOEuFjG3kiZc2ydhy9QZIqTjJTqr/rIX8yyjWLDElRQJ7Jpv4YJZ4gHdaU2Am
psWREu8PWzEYPZ3ltDXAIRnwLVu6DtftvvWJble6UTdFVtX2uWTzhKnOHKs9jMsTLA/gnaGCW0h5
k9aVD6N2s3u8kii0cCp142hzlyxfkbUxV4Lqb6nmMVo3eRKm2sW/7YmYgM+QOvD1tnnabqTqoNeT
bPPrSBTk6AJAIt8UAycimKLmCScYulvnmMojB0nvlt6hsB89eJbGBuGpV9Bv0EZmE55/stztabZ9
BrteGfumO4xEstdx2L6v8+wAqqhyxxjDg0XDo0FtQR7+xdq4qznN76KhXtPFaUNZry547zbnoOMv
DyaumKz2LHpGFXuD746SAyjdKRwC5BZ4w+JRsGC2LV8fImHx1TTikIhIU4tE1xhiQTkuD9eeCvbE
JWwqKfNjwBMPhp3YAe+TDVRy+5fLD2+I7x66FTrKkmvQJy4Q2fGS6ZWVBZr9GbTyxeEGQ1rKL6xc
xzJCTzzTH2QEqPKo7T9Br//BbwsYcraL4kpseYmgSNE8Vtgkn6W7k289pGk4CoYI8KgW+A4Y4p33
MzcaGxH5YwSZVJYnEekcXbAe3q0CgY9/MPTN+GJJuMgw1ZDACfCT0kuLYfLAGcOVbvtTqpTsEY4b
SqnPmYgME7OIxS3CqqMksQd26aqwfGHAP/zRW7hmABheuHoz1swT2F0gksmjsOHp2Sd3SjQGo+E9
kJGe87Xfo4cjtNiivF35B8CwkESA9/Lo5eBgFD3FNsSa5hQV9Ug+s03k5NbdaBcbKAy9Y7JikENa
SzNyKD6qxgBZENgm5nCh2qiOqNN7AfdDalkiOE8DEY4TMmCN0RrPmmH613QSDW1gb7DvJOEqsbNO
d4/JvASpzkzN0KGUOT4OJ2N6t0243SGRjK5hscjhtZdd7bM8OIRpmxGv8kXTqvg3FRLtUwweapLn
2fTwhY4XDuoPJrIQhxzBL3erb/vgdVRd8yqGTxAWe2BJo8DNtvxOgiU0OWGpZK6vZrd2THWLr4Hj
FH0/ClyoUN30/JlV4IMAHXwtPCTYC9XBt25rMC9QYUej9rFdLhBjQjdAcKZqA5ImJCqHtyMESdiv
4U0Le7ru4B3yZWTQy5FXgTfj4x/9F7mnWS//6uEc4uxlZGZTGKlKOxKwGoIf9h1I3u8x1x9xgDiW
ablec/3T7/BrFLHJgOmRO2sdlGtSlwo+alUW9evIcR1DOx7Fek4Y3nH6LBkOTsWrTBMqdSyW3KSV
uznFYVRRw0EV0zUIMnPh5GeHjHmnQpbh20j603Gp/fqg1kVjhCP3nEpVQtSvrHatGmDn+yT/W1y2
iC3P2nZuyGj3V0a5jkhC5ccVME+QmYiDrBDhfHnhTBhG0iiY2ezaYEz1Tx3eLR5+dMXATNelv2IK
Je0yB1nSjsZnIhCu88yju4iudU4p/pbjHzO3nh/9rMVFnVPMHey6/9jyCUGjixsYpIWvjumnDnhS
r6KjkypYXUQh4OYZYhlLNUWw3IwkT3bwNPuTiNJImWHzySOVE4OWOHYkizbtxpxPHAtr4hzN738l
5/2+egNZISpig3o2TmPi+ODHZ9QalkggPhIqTDUmJ3KQApBgf2E+rgpXxfhapg3Bbc6W7GHN9hDB
6vLDqarxqFgmFbFkS8vCeKcou3Kr5xnhRUkxRAUEEc4LCnWFIHX/TxmEOHVoMcR1SoWFwzPpauqf
0j/BIkqhvWUd2jKXtG9+CDjAQEmyEwTeEhjRKKe6tpBdqroHpncXAgrngUxt4TLqjfLIG3DFRKko
QDUxep4tQoyR84x5ehiF4Tvdcup7LrjIILvOR97pArodgF6Ch9vbZoJLjny8cX3+SlcCLH33qEH9
EBU/A+EHyqQHgUqbkW86QKivYVetmZ5w/RzKgV+5EkundXTTeIOCOl0qh4MYXDaw242jOR64pmNE
vj/XGeE3oA7fPfYPBV6+N2zI0Wede+M9uceW6FR4dYO1aPJEGRihYugJf8V+DH+jYnOmfCDoJqS3
5xyiV5AE6SB/5uxRJ/QyA7qh/BNeJwaXZpURgCI7pmtwPMe8IogW2XfqepF1Qe1jMYBQfp8uqiCx
M/G1dGEKqN5AjOkcIG7rOzxeUknQMVXBtFXFidYxTIT73IpVdO6pbyIprDfRpdKtKOsulN2r85Ng
ogy0EMraMfZtzwuljDXSnSvyhH9ic4T+blxL27kCuuZLcBiwHAY6QI9DfXkDARuyB/xdUPxYCemo
KUX0z7uV+ZIwu1b6uNAcVJmf13uIfqbQO93yrXgImy9oe9fTYj7Y/b7TGOJf14G76vSoRQWa/Bxp
qghbdtoG9MXbSdqDapx2csiFUyC3ki6pSa62srgyQwwpjgIffyJRTqQxjGru5a1r65oj2+4zEEFc
5aVWqf6tAaPhQzh971bLuV0UTkZNsnkeCIem9O/JKVyDTqnpvwMow0dQTuvgvhfuUq1hZm8bflvo
vylcaZfK+ShLV75bCA7toBNnmvxCQnh0IvMk921zD5xd0AUnsvIjazBRwESwyOMthBaeR50MFa6i
q0htc/jLaDnYdy/e2VUKiK0MexDNUaXcLCyPk0HBlYBW70t1wm1/msnMuU371SvD3vuuRXbO+H9u
DZNSxZmUil5D9rPxcfVwaHlhSWyD6LwDan7KbC31QlQyoRZ0F2phdaHdHBh9qdMUoQEiAJmOUQi9
EpZnPDf+HmZJshrsVQW1j9ggA8IzCHlgDo3ijkrAbK+xwtS8GGpk67n3f/pnKexBYW7sKFw6wXzm
QWMgTxTcZ4vqJZzrghASWUOu7Z32pLgJztzF3tNKN+2lEtv1qv7CZ100vPG+KjmWquB/Ovyj88lL
+/N3TOOZCovtKTaQ0dk8k7+JSo7Su57CKTTkzLAfEM2onuga9CI7lnN9MdPSlGAR1peeeOaASRfB
+jJzLHv0YSjQy5RdqtKI4P5XHMFZURSeHktYcxzjHEUvgpgtHOnrQfG3PQBQxVqhv3bMvzJuFqWk
/JH/UzTDlC+9j82twCwirn78RKEjEC2YZ97KJeZkKrLHCeEd9/zB8qvfoN11tDGxF7SDnQz/XyHc
H2Sia/KojSIccYqmm73gblqOW6CYofJvPFMjsHOn+nkZH0vx/rA09x5XWNkKvCj6E+bsLXLDN5Bk
chfkzK/LJGqYQX6NNTeiv4UyXZ3JqYba981TrvjDS6lwNXWuP/mW33NMbJG6NmCK3D6cDnXkwhme
NkRWGDC9ZaICvrmHnbruazQ2cZlliOv/tSHqDpr+bmsHuWlIPdkJv7+xfZyiSLQ6hjLj8g0JZDzO
7zMVq/mH6LeB0omK9L15igwML8xXDmNnm/mySuGo/rnujEcseOk1XvhBVdcFyDrXGv8dsI7cx2bJ
XuHIgMX58iOGsdNzXCUfh6LMmr61r0SpZquxXwEaUsvvaXykbMxVeku8cKhY1jgFYzK9ueacKWwi
gbG1aJKH9u4QQnMxgalPYkjImd+S4i8MKt6iPMQmgAMMfZOSRsMFsB7mnilb8lR1jw6Ip5h17rWe
BdpQA/XHLl8/Yq+oohAeQzYgoQekmMI6J0J3P1PgXubTasI6u89zBg2LIkzQ31se2IPOc67FWz0D
KXcM5LKqB4lxfFKYiH50IrkWY+/f46pWFB+EHETin/cyV61vI5eJj+lGe7HBggeYdgm3VscK79lJ
NHob1phDSNj/YqoZJ9jwF751zq9+KkNHiS6nYywb45vFLBEnbtxQRabODwqYB/fvSthKpvwG3io0
ulNFkUvH368SPwfQYQOQ/9Rx6o7RtJXIYIjg+BA4sciZpRRgjU6egYYn8NI++Iw3zRRQ6VOiTkPY
mU7kB+WCuKjeWseYyygJ0gki22C924XV/hu9Viq2cElKxXiwEUtjxToJTZATZcQB83Uglz3PahlM
lCr8/JQm1X1xUKljwbhnYyQeWZDSYOpcD6a1dxMeO+u8TuixeSZy+rEGD0mJ/HXZS9OgyNTDdv/r
w98YNqQPJfWcZuqS1kZtSrAy6WUnwhLHhv/HU7u9E+I/djL4aAggkEJJYCizMIh1wGOv7q3KFidx
144yAKZnG3+eXsQ9nO1HHqZmVMsrlOI+gDBVXD1VX09Bg0CF8Fa6vpWGciLBfWV/0REGoRmQXcxV
tuXFwpOT0atrgjLwka3lYDDdMXcyifjz4Z48HuZ5mCt7AYJtMG7lFyC963JuBBewwcnCq8U42zaP
h7+RSD0DhlaqE7Ic7HmDeUnPgFK51ua6K7uZ11w1Txpqea8APG+Acel1xOeQ6gQ7j13AWdKA2BF0
K192B+RAkCgUMoylOXE0JisC+y/ZebGm1R1/BKdjOKiHGjZHL/lxLPY/8RRt+JGrUj5rrwAbvBaU
X/x2H/Lm61tCicDqcTW3qZkRZLP78O85MVHF0kKpzRkLIVEtscs38HfEKyKUNR4Lu2eZiB3b7jlS
GW3WXdVYcEf3oskN8294YnxfAJdsEFMHS5RBR/9QRXiYF21aY1C+uf+e9IsR5mwyiamMJDm16Vqa
AQbMXK2PJ9TaDSAFZqoO9lhc5VUmkituWsBpebJ+qAUVqkpSa5PH2n9mYwGWC4pvNJJ+MB+F0f/3
2FbW/k9CfVURMTWDgN40Sp5Ua9JSb+7xla0t2fSookJR6cfr52CqS7EuTg0eelFksp41aZy/CGlz
5hU2krJ8+gJMdseWW39iUbiZF7Vu9dtiJIEQA2oP4JSRMF9TkEuDwwKP3YW12RNTpEm3BN8jFTsD
94WlYZn6w0KA/YhkRUE701moDEXekMc1kEMUN+1iXK9YMfO6KC6BLL+B1JT7eHeE69DmCiPWmgxG
E6g6BneoSGd06c2OZRYtk10JsRgISpx93G7xhGzSaLqKXEBFp7R5lLTezBgZen/QpeVMu/iSBMMD
KZgyXGccHOknM/VNmF2cUOP9ku5MLwMIfMrR3jMXjGXJ9GANKvWM/yApdmctbANLuUZrwWDFqohO
BfLso2rqxusUh/Fd1kYw87Psh+Wnqr2UoYXsnKmMcuSqJE9mISiCvNsB2hzP9Zzg6lWng/BQnd1V
9UghrUY/OZuxkR+M5/7JXRY2gpvjeHE2BProcfF2NVUUJXeKk3R8SlKItJY9ddHpbwXftR3t8H3p
JvmGt7jyHT1gZseXvh44L6hoQ3QbLs8Foq1ZSX+Gi0oQvL0OiGV2KKYBiIrY+xjXmpk88fRBM/zr
ck5hTNM3/LdiEl+3ej9GpE9zvnyLvU/yv/A/ZApDlCHAWZUAOS1HeP9zRG+6pNX+d3Nd3SAneARf
EsltYRcR2TakVi2t+Zet1L2YAG/2DG2z2oA1p6rfgFIb8M6PsJjae1AgSBiPlv4y/d5l1ZoNGn4f
q4CQn9ufvNXIlKA9VwPkSv8TRHQzrKwaQq7N9KOt9+9BfuKtMOxcoGcfpoNEY2JhsC9hFEAGcfj4
lNYPYXIXeg8BHsGfnYvQ7Mqc1Dm2gRYdTnTnBG9Qw4EuDKzH9TTmzNVERWGlU7QdBh/UVJYBg6Gf
/vFU4oXgGFfOpc4KI7NljtGgTvmlLZMvtWY533cZtpBqJIdcmFAKGQzRZq28u/4hp7SWfek3GQvB
K0jbOzZwXqYKtoTlpldMEAn3mCz8gz/7xvtIggYX4kFqKMOMeRnxZDw9rgO+7144arINmbyyD0sF
M6n/8vMxgMxbVvRryp0/E+nJq049ne3cletQESDcP9iSq8o4IkPJltTaeIRPBmJClaLXnjtHtNEW
K/61jHweK/5N1MJ6048anuTHjgLqjp+dHNOmrspWJz91YlsP8g/HmjJt/EmIwHn9qdo+omyhVp30
Zqae76MZWsdxNE3UHULtc0jRtSci2aN935a20w0hx6Gyka+IZISpTfrjFCC2lK+6V94msrQtzuAl
UiMczh330bEfYe4aYAQWADI8sgL0xlY0Y4hsZbZgjjVR10wN9SKRSp48MVG0Iirnd6PQCQ2Ao8WE
0gevtRI2Qk7uscgzXhUIHz2tc49H6WiNolB+ChhoM+dELmSq+5RCwLl35Pm9kRMXkJWbbDgMywU1
ZpqvoJX2rQNcERc5ecHBZeFTWX6AEW9z0ejl+XpQhxScTIAf6o5+WoR5AWe+itB4KC/cdG7PkKcX
5uJFUeXCJthr8Pgn54knoCceTl3d6rOqfUhs5v4xkUsDsYn91RmhQhy5XCloI3vTV8sZDtfu+XCy
gQavTbYoUAysG0OaixGUHVl+h3O1WTxuyyMF9Y8eoO8SDs8SErWzkcadnfeZyRVfvU1A28Id1pqB
1RkK5gj9l1O/NOzxNvJzB+2J6LXTVQS2RFCld1HctrjM5BZAUsYzO2QKXGxhdZOgiQGw9veCmObp
/gZgqhB6CCvHQfSLnjrZIUXAcMHtC13784aBlHjENnOqIkGk8p5F4nEYsQ4cHb+0+A+36chqcb0A
L63GdLOF369f45FYAwc/SMI4atudgtqRNE0OF8zPvFNTeHXWsj3moAcBODdjMTyMTWBncu8LMBah
wAYSJ8drfT4B9JAWYF8975Jdcgs0pXPOI370bLSt7CKy76qceprZNSCpIjbqUFxrKRvyQS34JPYq
ozlWH02W95ilSiR/zjG0dJlwE2LFpOXgRisUd9xcYoebbIPyWdBSRwIDdL+bmLb4euqt6qUOxIsk
UFP4apEk2Vd4abGezHVOhD1daT0iahSV8+DlWgSRIJ305cFWaniAcCfm2ye5Sm1hBE3WNRTfN8vX
c+TcqCWCiX40U5NPHRq1ebp9dVNneTds4DBhLaUYwLDClat7vuOF6zJ0suYgWwAs1TKU/iM1mxbc
DiDVLrzbYhjzMXX3lP5O1A0Wq2ehynWi8y8A8PtNp0THzsSPirQyiViqwsO1MrECHH9Nff76AW+5
Kk0woxqFeb8u+6flz+gKh1W/l1k82tjE9BL5G1VuJRlUhZM0uPQKazBADKTCLkqcEesnWf+96cct
VP7ItBc5oX9myaRVcB2KWm/nGa2eS3q8TP+3kSZKqJFQTYufxQoUwSNfRPnSfpHk4l0eLlwFsuLL
6yeZkgQyPzSy/2FCZCA/9kyFmANWxF+2lz5wbkfFRdC5rIqaGzSiaVKYHszheb3GJfBVarUl0W9S
ac61Qt5D4zLq48K9YUyzJkfPjjvLGDoiTv8sD7S86cT+bBrOTV2u7gGvvhEnjYMkM7SfhfTWP6r1
GcvXq3kyoHc4YoW2CRHSoyv0yH0XOmf4U0PDPG/3DgqZCFZSpZI9HujHyVbZR8fWIK8Be0Jb1GZn
ogAolap42ahDESpu8vYUeMcbfcNFPzdkHL38gHkOw7jSBIx704nthyhiOKWvBE1NgaLoTJo9ur3c
9TA1sICMTeTaG1sfTfSaJiaD3ZLGV/Ed012aAEd9/VUiqITjLKJUAprqxtxwm+bvopxm6W/tEH2G
F1svzAaBqEvK163AjwUN45GwaJKLfngUu8eaPKY0y3uCrVZ2ERneftULXp99+Jq6t2mkkSLmEqeW
7i0uWQcSBPit967xiGD2Tlw386mEqO7OpkLIj/IyH2Qiu+iMqc57J0lXDXxk/obfza4oJ6y2G/0c
Bsfh84SHvCr9agD+1c0A9v3txrG+7hnE37dX7BTmHAxhajNIB150oScXAt/OoG9l6SafHoNVUK5t
lLaLsyuC16dZigBmYGN6oZ0gAb6Hn29InyT7ACcM2miK9zkjYoPTjqtf0iVTCuty5ucwhnvWkKri
rQt+s/3Xx9oRhOe4STVc4pSCQoBrKvcHN1b8gMSxa/eRjXctq6cnJYtUFuGLluF3AiwE71GlyZB4
A/+3ZVdchInrSo9TR2UFaLU43nG5P3clyx3Jx8ERhIMblRBdW2m1+y5A8/iEYObgYqn2sagBuPH2
5SydTqtR0ydhQ20YvuYCRBpiQoTY9gXq9xavDZUEuAHWqjIIPOAFjMqOiBqrQOgQkifLZ5Asby/J
C9aml5iIhaYo6DvSg5auMCN+aB6DuYGeANVOjWFL5RohTyPwFHPgaxAwHI/m7Nr/++65/1dbBlGk
3YRULQkdQyM2qELZQTds4FjG+q5R3ANr5ETmyDGTZ8+KdxYuWrgRyphcnxL0ZQBLa13+F/AFoJLO
aSUd3N+nKbqoks2+gPylG1bxMaumFyMSo23+aDw8IaX07U+0kyGToP/ZLYA37Hxt09zRSQayynZ8
8mmXTBRwmf7CJJHNSWmGdduZbyNFMFfBUf4BcHIWzOMwz2qLIz5TMsWnygmZuBfaaXX87+29SUD/
DVFM7kD+j7E+64gqoluBWV7A62O+0kCNBrgqotGPGmC+rVf5f+MDA2tWC9Oxp030mD21QwCjsxsc
V0tp6wtaTAilxEWdXYsVNxkd/HEMAu13NXjxYzcQWyOLgL3K4enObUW5bY4C+RLrqqMp7J9nJMy/
vjDHO2kwtFJJ+jbh87TP5xWFHNtVhfZ7XTpdeBOU3xoXkqLf9m4tSiB7H8FjEplRJBLhG96Wu6vP
Y/bAWiNPf8c+gNOAqFG7mG29b0n+E1nrUOT410SJMY2vaCIJQEQpETNwx+FBkBGYa4M/NkQ3g15w
4j8SLSKmiDvIi1JYoJRUvtG8SbPN+yaokEurXTCK0/L0huKr4aD3NBuIluf7yAGEnOiEBpBvbS8P
a0P7y2rWVgqEn2N9FXclPtv8djomqiKhXDWqi+r/2+FVsdv4ze5pHoX0wiQygmP/L84YYulaZAbq
z2N60EUYK8id7zEiPCNnYNSh07kBHM3gGmfJifvPyYt29ZBRKGlN34xERKm3K1hBcVIQeRDJDcY7
BATZy/wHDHba+rcOl7QfTzUcT0VJeRLoqkbfcpEMBjvVDwL58ure3+x/U/8nF6oySas9gsX1nd9g
BZWfiu/xF7dEybZN+HyxLsE/YdrSr+nnWdC/5TzZezaTNLlFxtGEy0idnyMTVPer1UqHYuLPPACW
imEDXd59RrcgxnF0fFHBb4wRlOwv8TZlWnD946SCwQ2LbA5pJhhRMpOdq5rL/RWjxhTDkIYnmPt8
SpNElJQv5mZQG5F7SZhBG4ut4WoCys73GtqtndT5QTXvLsBAXoVR+ROrxRJKG9J11HE7N9MdRo/t
bB5IBIrI8PWnc0nsufkTd073z6h8tGVrQJmz4qKVrwrJ3OUuAWj29hcQF0ghpbFRc2Gp1gnFia6r
naG3ZSXZyvtGVkhmYNZ2hcmMpcQBkN/1eCHqFYsEK6r2hY2aSelDU4hUy2OladtD92AzzNR0sfXE
abQL5vmS6gpcdSwHvCv+N8B8tl4FqP0NelvTLdviuk+imG4AmisWX2SKOylbS5tbM/8DQ6gsChdH
vkhhCC8QZOYmvdylH/lMtbG+rN8bwseC8966WpotEpbHgJLm9PDWIxx3s8EAMtcfGMoNQrDM96ot
OWIM9wXWEAfz14GRkJ0CyOEoYi0qOVSBMQq67i4msD/F9h1/1HF5jG12wgH+YqPDAm8qMAGTFYq9
X6SU9RuDyscgs6UDZyXBs5GSSk8+5OSNhCWODOGOQpHfdUualsOEfWiVxovm2mEBx9EGFe5aZW8h
fohg9yeBDTNOR6zA65A2rJL4Ta6R1DDMT0he59pIiBQzr0Pya/0JWr+zqmhwaBnkeEa90/cM7hTH
5Oy+rdDDk40pu2GK6ZRq2tKZ89S7xszNVmWQZpOSU0eLWVvCjigPqFVTHtPtQoPQG13rZ7E1I8Mt
SpK/8DrIzGIlKKPA9jBhQ0NuZ9oObeKhdCYYT4IdCjdyRrTlcJUiIDp65w6pyEfhuGfcvsnoKQ6R
loDXUTYiyfZRUTLELMu3PD/Sa8zH++A/XyfKTLMjnWU+o61z0g43xyP03CS/nIRx36A6OS2LDnUg
H1ITCTndAjLqOcSmZTG7I47tY1yMLtpis9tOntE5dS8WV8vYuIlC1Oia4JJRglHFx52UCR86wZ+S
1/BGnN3Ua9vAYgby6ZrOOgQASuvxmhdk3Z5RGvkTVVQ4pu4ExRptzti0skxOl6ULCtg/KQ+oMamo
0VmWLoP2WPYUuUgYR5eUyezSbJQeGcmmKauRCS7lIk9mgLQAtE3c+l/n/8D34jds9OmVtgJvPl2W
/r6azgI9xds8w9fKGio/9casCB8MRWvxRoqxGsIcNWwiu7K+9HdRFZuj1MxFObkNy6ci280EII0I
Dsk7XRHVIe/KbnHNQLOxD867PeU0rjJ2Du9HG9FloujuHpUSQx7d78ql2RmTJzNIRz4xnlZ2q3c6
kJZHCCK3wjoWMPBaYJ89MMfcgOlGtTDnW2kwI0f4+BrTZJYpGRCiapg4tguD9gLso/g2JdiG0DtE
uVOTy7kdkYnElNZPiPmxRIT7agv8k6rnZ76q3U+LlPpwtRc1/aE2zPi5X720KvUpIEIqacpLGqaH
HDEE6OwHZyC6P4EMYDJ/1sFUxcFulC4SO2a6T69FN9FmRN2rVeFrb4Iz7EuReWcEL9A4r14HFHzL
FZbkCUteEEuUpCDa350aafode4cb8CCRuRS/65w8DpofMG2D2+yyniKNS4ZJf0Xsp/cKHepJhITH
QyXOaJ2War2nwIAjXrHknK0VBbl9ySL6gR9TWqA29dwbQ8CCRGhVaze55ZE5/u8Fm/d53bxMl4k/
jMuW5CtY05L60gLbruZEjNJJ/cwTeIqeg2wvZ4VSm6cC6b0YTK0UB9MRLnjXi/TokB5VWM9SHP23
v5TRZh9JJ95YxELpe9ryQ9ObxmrzQANfan9xjCm2qPJtn2nje44B+OyMFdvzCwRqf+h85ciE64U3
PNSZT1zG6PmnU75uU2XlrjkKEEJm5EHIF7yn54nSj8ivKcmKNbz4dRHQqdl9SeHhYNNX9xjQzUfc
V0j04wyvH7oeq7WvslvzKnSuFIVbUL0EZWRclq3PL1jAiKVlh5wgf+c0C3MGCj5IFm1RKGhXJRWx
UCLs4u85fdGhRDEHgzkAQX72NxyC06gXEmiTEOqIciJ3yMIwqUxFZ7XkQNwyBOt1CH5L+0xQtO1T
mppy5Zb32PcSDApQXYu8vm5ebJnwpYmlN9yf6+At9qbHH4XPX4p6q8pit0QXQ4dECAEzEWHFebei
nOS5um9lg64lPkAZ3vvq8W6fHfkPDh2jaf7rlT+T7Bj41jGcqhnZGqqOPfKdEyQ5/peEbR9YWfVP
dBrIhPoxhA3Xu2lYEuE0AjtPpdwkR/lkba0ousQb9gbD5Bc7uyDq4TS6VWboNz5uwkpjPxWn79c/
2X1zCWpdIqp5MiB42oS4f7QDFg0O8IcnPytQYsdZucATTNkEIz9D8+x0USiVIzjJO4ibiziC9kCp
GYTEpgrklD/4ILGFceDKiSMJDe61MG3N3aXJJ+avn/fx7mNRsQfNUH6QbuckULEOKoFJgXNptW77
YhpL3zzuxXX5IncwBW0wZxRa9aOkcQBB1SjeutYbWtNn7X5MAHy2af5/T1nIlJQLuxYoPgZEKHco
GvCVP1OTPsMA7DLZRkua2Jg4gtDzng4QuDmqSLLsHN6r4sX0NgUZVYnzuaV1U/6abZ0auQ2AMJ96
NQowKYscIoE/PssnAjJwj8nFdTmU6K874p3md+c6g+1BMiZofimlJSKSzZM47HbOYeNsRvsJxe0W
ym/g437z3bwm9T51t8bxpBvggey1fJeRO7osII6P5LukUtKfWLf8GvAjMIPVARtmm0thTdhNKX07
It91yBZFFaSNKrti7EePTEkKqPHX73CsC9ZZPVPmtkrkwslbuDdCjghpHkFUVF4KWEHHyk1BZq2b
ZuNvbOkJeItpUXkRLsDul6yj38pU02bFihShqfUgnKMhP2NxhoKYihb5EpFlZEZ8HPbCScmZf+on
nCDYD2az22F50+1hEFAt4V8jOHDd2/p/vtgKfTcaFEbtcAheb4HpGSR8gTic+oYubp39Om8CzfH1
bBpV7ND1U0pX+RlyHyBDteZ0tOcA/Y2fxd+zwhNS4wJeyTk2SPtr6r6cR8fYXKTixev0awN7Ihzo
eRqK0QmBl+rubVzsPbbUXr3f/LO1j9zRDol6UGOthLT6CpMCn7PYQidNOw/E3J0Qd6E9+raA769R
EZ0C4S3deEBnBrHVtKwPj4Gaz9DJ9OB0JkDHPKLoPnnsJQSU/BP8FpbdPT50ga7Q5voeQIKqyi9y
GmiAdVGW6wFOL/tF1xDgtuVcHkLAiH7NWrCYRR5cNRVzfJ2Dotilsfs0Zw3vU8YUcnGuTAqlQAW0
H3FRdV6trr09r6h2n4UfdEuME8iGf0OvI6/nOsr/Qx2f+yNNO9f8oLH/a1u3UXkQByo41C+no/fb
PT+Q5AEnSPi67Y0AKThugw8IfPePoa9ZPFVvH0R+LDWNZg6wgTavXjlUE2s9FymvPHejYRk0C/H6
rmXahotJkAI3NBoOE9PTwuCQU7ULq5KwbGZJm9iFKm5pXkVl5oHR3bq++wvylk0PBxfnspjnfl4c
G4sqj54LZxv4QityoJucqy48fbJEjXavfjYVKP/SXNCuhZ1qm6ZEmlZPv9m5eDxF1KSvvZHGoJpu
GOqDAJa68e0INyPtJe/v9aY1/Ep2diwPbHvDQRDAGcp5i7irhOgvAZLKhhCy7xTN4ELYNYqVWqF9
kOGXsX0/MoDBlWPCKx1HR94Elw5b5kjww7E5rsYAU7Mk/xkt+LV/LWGkGU4ehabu6Gx84PGu3yoK
f6AcZyCc70Y8wI8IVUHpn6OrEIYpyTsjEoezpu2hSChaKi5W3bMqi9t5f5wb8Pk56AYK8McSWLdg
1HYwkG6wSSKgN1ahz/o9Apyw0fhLOCzmBPu+OMNmuZew7PBdMTu+UbyMCAlG0iQWCQeKSCROdVeA
F/Bme0Mhe6rzPKrHm5E2ZJdUXXjN7RQG/fVSdUuT7LpJEBfrWJ+W0rlUaL77z1v5GKKGSbUnm8a4
p9GuPROOjffXR7W/LbZ44U4TkKRtfjaLaYI+6tYPp9vvDeHMpQdK/jsnbMwrr3hDuRk/O4et3xiF
cbsM85M5ToOSb5pG+PlLbcqJ6iT7OvEd8itBmR5iyvZ0mURHtwZ1i8pXB/JMLEkMKWgOO8qrnpxX
11kIQ2lo+b4f6qet1rQ9oapTASYDGVifTYzLE19FAymZof1je2UmoIOHkOy4TC+9Rvtl4kij1DSm
TCCm11HtzXSyIAvQfbxTxbsihdQFsLVsJR3A+U2Re5V/H/B17Gy2tKmVrVQ4LgT6d4NFe6pLkO+S
1xpRazSnLBO2dfdiqqAong3s5uXt5KRG1AmbGfAjglqrH3eh2E1HPQeNvkNvkBtMtBNCfxX2hyXn
LhKhG7d1+GkkTnBqQWINu7u+u+9kSAjBD5Ttvj6SV86XVvj6xANH0VJtl6rX+DpezkofwiysA774
ptklAzU2ELRRLFIdLmBegvjDRysdQpndfBm72/IXVRBhb7aZ0P5m2ewg2Y11ldCZw+3gc0vFmilC
TGapxXgpXoQVZQqC6PG1zi4WFYNXIbodlQXKPhB/f2eYNJfgUSNfFNnj1XxBhJZillI11CsWTIiC
dg1GBHIzJdN45zYxe49MktuC8akUzuQWB3xAtDRTw8utmTeI7JQTxkxfxvbDYyGxrJQEwodIta3A
DfiaTrGVsPOryeEy2Tj0kfAtw4PVmVNrMg9dBmHgwQiRt6ao8aACHFB8icJcLfsd5jMyXOlPSSdX
FlJvaA32imFs3vAmhPHTMflLOvnvhVNVQsDpP58f6mS1sRHtlSyIXscM6ts+68HR9LLta/CLMefK
Snv6QahF1DRYwgoXjXmVQ6zkgBoK6+xnvBgZLIk2iZtIzYrpoizHCN2UpzlKm+6hEaETt/1pFQjl
CbocNdpKGtWbp9myXhZPk8k3UCLY3mddwnQUGmEQG5Q7vX3zO/gpc+CWyV+usYIQMQSKDFgmqLE8
SdsxPqJRZ2mN8WTVTBz5nK43qS8Dcf26zpk35SBkr53VlYBtDR6U00lEaqdblmoKwLzPFbcPfuXH
hdxk/rI6z/B2udMAoLXgDjptlXuqjmMHgwMiB6ieziPREv8t+vF/OaYwA5D1vDPcid6RNN6ZqsSz
NPuRayNbXNHvc0MZ3YVhv1kSbuWHlkG2avHPpT4sUcf7uBMi8wQeaTnD46STfN8mhoqMB27evRhH
oMaHJi+A0UbRJjqlFk2+OAiWlDoZPy9vkezvZpgnZ4DzEIkXcwg4QhfMZ3W/8J1F+9aJbRodyP/u
V26fouGpYzkgvQngVPT3eWbW1CrlCd26uYtvt3EG1a/i3yXNO2xEDJyXd6L3ZDOZZy1Olj76GYhY
WM4wqmjLZSGqDE1mgEv0BlRDd6q83fFO7q4wmAIC8OJGymBXtNmtnAOJXPAxvRJgCRBTbzw6m52g
RApGCz1hWFuYuFaTjfdpKYdmsELp2CprZWoK3JYcG9DHnPI/VoQUAP/R5WC3CRWaMqv6vNu2w7pw
r7DCNF7QZpb6R3U5+e+X0lyQNB92WtfSL/E9BJnPyukaLK9k2qdi/ZqbTIdTjRztrZuHmCMjnx31
+Oq0qKemx76Z+bq6Fx1fmIPsLC6+KqJod0kuXEy22sw0CSWN0akaidszM7MrTSUViqE7pf+8f8vY
JqTVg4rE/nq4Fpdri2TOZmj4xGCspxIYyYIBD/Fad0RMXjZ2By9uWU2wn2n0oyZnau+4f1Ch7WH5
0q/+omb6uIkr1q6NRMAB/uPtlsOApPGYs9r7D3siKoj3WZLNuyqYRY09OdHQa5sn79UN4H1piWhN
zzWwFXI8Z8h8lyJqUehx/IPCDyOGpGoAxgvYr2vG4AFBec0UBSdktxlti9OckWTK6IxE/1J3NM2J
3hwx8UKUbVxTSV8R+f2drtGpihVxU7JN5DGmB27qyOh4r0dGgaPWXF+vJdG3G3QmV43pYlvTMuxf
K9fypA3f6l1MRU57o1fyHI8yi1oA4Ac5yGYM4Cyauj4o4PIrbY+NhFX9DWHdH7nP1UbJ84iYGMfC
3rYPdFklXckenBlNDF2eVxqx9yLoJPZlvqE32GclpVrj2yGkSy2dz7QeIWTwxATp+aM0DVmVAVig
BcmKW8dMIlU7dSiAwYiAlJFdmZicd9VpAL2FTV6GRwaFWXm/JfEgk2WkyIxIhqWwadIrWskJ/Dla
ie40ix4FnPU97KETSCLBylb6WRDJVP7V02QDshNtm8UTfTtjDbu5llDU0/KkRPXe7tR79L7a+c+n
lUWtcxgokqnGOaOHTcL9cJGviZu/7EvjQ4uKX6IpA3UxZnT8Uic8pyw27LNaI4ibwELCQ4B/t8q9
RPLm8IZrzbQp+ccF2HJCapFSd6uoouWv0oNpdNuZm4l3ug0Tx5wNIkNIRTUTOkH5grUqJqXk94OE
Rm+vVYnqvpjkp86F/R+jBDHkZ2GdfSP2OuVJaGtKldgOlgMWFZoTB/dsiOoBS/E2B8sATPpzebxB
GbX/GIXvMi0ZnYmqtRZnUjXTj5OdkHmF4/z+73hE/Yy4R3fdzFjl5rQPcWTkhh1xbucD7+fg7G1Y
1DGlPChGTAYKpBJ8ce41zebGqMrikWgDkZiBjXoV4Ywa7jxwKis20clxQXikGcNCDeesGn+jHONj
gc5GLSh99/mBBLijrT0arVaU0LcepzB5aWx0Ij6JcYSJ+ZoNkAvWrsiyF2Q7YfG0/Hg03YhAE4AM
wRi6/Z2gFM9NSQ2VFwtM4HgKaI4rzxzRZbcqtVzlZ5bOcVkPfwfJyCIhSrpqvBvIrjf+fhJqJMbx
rg2jH7ZFr+W4zsx3G0i3NKM4tdWdQ3j0kq1oRDue7MVqqXWqKhvG9OUo5vNMI2/Kq2Ffk6aiyGMy
wLUUcglyjnzHV9yv7fpt/YRmB6q2wQaFYN+mE4BCM1O5ER6skiOS/I9k4t7E9DUlc6yo36h2VelG
243JsgT9GQo/n6RPmi1T1aFxhBnO/8OtEV89uNb3+Q/11XqQO0cpJcMjeVP3mUMoXK4QMW8unsOH
U6gb6BQsOKmvMhaOb/DS+zPhXdqn8yJh/NXNC3gu0WLJJQbfPSxdjKPFybKM55SjydWiSVseOJZA
rmS4onX2oqA+ZgZhnSs2GsklVe69h7khJMpeRWcbk4W4KajmvU912Izbj1bQ+7r57qDU7ex+WQ7F
hwcD89nKGkv8taB6pn9D3Vbo26/n3sdZ26HXiJCbAyXK6BCXr6SmtW6f7JqsFwinWMWHEVUcnDk8
Tx7+w0cLBOZWz8KHY9VBJJ3JYbM1FGOKoTZuHuv5StUlJVL+Q5A6OBz/UWKcaNtqgk/tMvIDH9sr
o1fAvjBtQb9wSp7mBeTQIkGFxaK0X8EKjzaMWQcs4Ln+QVqVUL3bU6jwdXNhmVcyhktc5KpQHWVo
ejJZGppaZHQT6WQoJKKl0VeG4Gxr5Wnp1RPH4KfGKsCjcJTzI5gfu93fxIF0xPChqORPACxqhDOb
OyP7DFZ4SKLMIm4w+j8XtzducJtIh0owz+E8IjPZaaLwd7ATaMY4fzOZZ00EY4s/BtNF7vdYCoiu
71TEaFqUmswUgM7Y8W+KxOugK35pIvTgYcvzePyD6ONgj3+ommFPkXklHXUYyRXV9q6dKSpJmfAn
2hfJ7BxXrGfVPIZ7M/14iQ1noL/XPf0OALR0R50bvP2LtL/SK0K5eX8DeMIokK9n+cygSrWm0sno
AG6xRdqjQPLqOz1NZLlQj+vGslkpkUEGizb8hJ6iFDKMdqVzVQvV7e8mSzoNVmBpoNodn4jiIUzH
xHqjj4YDihsuMDuURqwzzHRnssuwYmxp5/IGHL6kJqQ61YIAh7na6WJR/hh/Eg+L33UgY/r7xCXf
N3qff/szALNThqiKWud4X2FfsesRD8wsigovVdbPaHDmUnRK15nB130IYGHtUaX/gwBoEqBYrU56
KgTp9LHGxhL/Rhv7Tc997fBJta5/6vK3oGBO28/SWu6E8hYbMobHIIPodf9wPjVRB3cQF/gO//hL
yUr9KhLM5wlXALsD04dD3Wb50hgTNpwbf/sMTz+jit9eZxO1nJlKBRPLaY4lm97f3n6puGbU1wNY
otMV3vng1y4WysVBvAu2wMLXO344H/emecgvHZruS5vBdHkj/kmzHdfLwaS4w85ZlalfWvV+/MOu
tw8x8TKUk2ROwNuZknKveQIyVK18M920VbNlf6yKQB5gt4dpy/pAICvRrOZTeDa6ZUdaF0QwUFLy
5u91692voSMlOhH6WrDvhMeMlaErzI9dHc2Gwlnapmy6I7VHORbS1KAmj3JmK0Gy/XF/n8yXETy7
0S0pjahLWLw508LtwbVi1vtNmqyItKAOeADaF4kgbOqNImdtZVwjWHjiQGV8F41F0kePExxR3bmN
Miyd3+9nAhD6kIUGW3NKyXggx6e8CGzRQ6BcB4jJYH0fAUIQfWrQ3GbjS7ZOmkC3xjsfuvTbl3PP
qJxmhZbbWdu5H6RoLF0PAsZYgV+rVljrcHuk58P5xINtYw4A4gaOTpct0f11+uxkQvGqVdE/YbkG
W8uY2MJ2aSfk6l2lW4ghRer8HV6SUOC5tH6Z111YzAcY39/bDCXI2JSqI0M+02RsMUSnVZRD4GxD
MpXv3tWF/10axz0kkh75daZOMSAzsbVfWGTs+aO4q1b11MsypADn16or5R16eR0WfRG80IM9tPfW
vcdDviTkstbLsd2LtaZ8NbQ2Q5sJ3BVOygVKkjWRKaMjblXhTVewChkLKGkY+lJK2tfZ5z7qDxQw
WN4T9CIKI9hHx1sZueo4DaizsqBTNDP8aDUQkbVHZ0VF7F3GfSRKlD6FHPZqO7cZrU5n5LK6rgym
UTrHgJgS9dpqCOAqqJESnedw5Vyhv73Kq86ZvYWoP9ZrCxtqsrx/dcenAAdZ4uzo6IkGPI578ndz
I5AFtUhV1O85yOTJoE9tOW6tKuPxxTBKpbB9eyrZRyGiVq3gKyLUsNODDbdj1bAGljL7XMox/dDl
M8QiFgKA3q9WvMPd4OJzOf9RJu4Z/GRPjiERN2BDb7fRstle9NSvbOSScyA01FV6tdJcBkPbHqMp
TW0z977v2O34PEJsr9uudopfYvBuzu356DX6kr0dalYRXjxsQQKkg87CCJweMYdS1tEkK2XsyYgU
onlaF2jcd++ClWJGW/h83CYuX7MoXFAT10Tu6/o5Y7nG9GGrrhgfA9uXc7EEVooJYK6dS62ZlQAJ
S+duHRy17q5M+vJvq7EwJPL9yYZBIpHWX/6Ve1oY8ElWiQP23kZQkNEEbdNGNC26gNcPCCtWWQqV
n85VgQ8TH5ls6DRoBL699xlH3sAyxHOkbAkBJSHoZ77rOevR1lV+KPjmwih0H2p1LUgs3AIt332C
07lwoKYAKMgLjurlL5tOSaEzA5+KiQyE+uWLa19fLXlPy/y97/vZf31tNVwDt7exBT0FEoordRky
7FrL0NpuffHIa9S7ScD+aUuOH4FNVSPwJiGlwT4qIadtOmN+P2FGGy64TG0+yNgLxBJ+5Fz+6hVD
5KhdsREfrBakaI2Ej4BnhukW2KXNDz4BHXqi4Hj9oHeuxzz8vSAbKu/iY9i/B8F0rQzNXZ2Ls2fR
N4qu7ag2OR2YiBTJUI0Vm0CA7iqkNOor5UVZ/TYRvdiXWdLAfXI4jnZ/VMhhgT5gkj7pLsZeokSa
tj8DJnObeNOOKugq/nDbfT4+ZclOwczQfG0DkwR5P4BFKKQV/mb84OuM1LtjcF7Au9T3Mp6AatdQ
PAps+BO8EuOCN9B8q/JYj2db8+eyTEcUzn3Xjyvx9nwA0v9YjaszOXB5ko8ZuMFXvRda+V9E6pyg
ad58DemJZlelCJQzsYmZEgpMzPKuu2niL6C+JnLcDO3XInMppU7hUngOjmBrN0vFNCvsgQFQRYEM
vENG/RzjHC3fkOdLnfLneI21sASpKpTWM7miORxnEdNsxYULTdj3QdCOfbFNLtGZoG/MJoPpL1Mz
QqDkjCmAPyhlul5V5lTZVM6OT/BYbLLeAyJ7wMvxGHhv4Sr/6QGXFfG3rE/5triAbAyvsvZ3K8LX
DnLAslgFopcdypOZKrR/u/WRiLYurgdrBKBiWNWf/U7eGzfzQ/8/si+9Ky6YHVzRVaowBF7Ne26c
DpFFegCY3m/lZ2cxvIAVYovtGEhm9bWgfP9H+C29FWmhmOuJyqi1213SotoGX5AiOfRkolHwhtIf
ag1yHqo9JIpp6+Ril/T+Rmy0uzhp8I7BX1EUUr6ILkk6sEJFEchyRr0ZE8EmdqH8dtANIPgBQGvr
EkB5UN+j/h6gySAQuLiSkq1owsXd47Ve5u0D1CTmwLJHXXRwnpHjEussQqMl6s1tYy6jllQIwleH
Okl5NM4oIM5BXYm8tNlESgvqYQ2nZzM8BltXAZP88Qhq7lxjVSQofU4Yzl2W3si7jkm6hbXEmubA
NcazTn4P0uyd89u0xrAK6eLrDm2O416DrbBjd/VZDX4RoFhSSDB7uCdjo1PkTUWsP0oIT+jASBKI
S41JKyrOYPAwFP4ifn7jpDCxlTndAgISIGEohKIm6T2T71n6Mqu6v3K6LqMg5WxcmpaTcSv0JUOI
ttX3xONWb+LbDvKb22talXMANjVuwXh7U+cMOFJTydQLERY7OCpkOWrbaQUSiXUtnUerwf2l3zZW
kC8BRZCv/DF2HqX5FsLr8goXAX94EFgBFlOWJ0e71MG3FbUJj/zPf1Dn7hMrYaXqAqSOcudleODv
a/NACZMBjiX36xH3laNx7LBXCFx43mqU8itIEkaphibBJIQCjm7MoFVnftvtpijSnkaQ3uP5bH1a
6YLzitmU0M3hNE5+ENnreStq9IlG9vdiCzFwnjV77qKU006j+T1lNBAy+GYOVuxinfDI2H1iWb/s
qyhn6WgmoLcSOyPeJzYDCg+U2gojJnTsUAvf1Hkm+kqwMMhhWlRzsfgHWTI9fPXSRsNr3q32sR3A
gmQ3i0qUlOr5Cct/cE8l4PCNXmWg2eqcGKzBwWsHlle19Fel4yZJXiiUvfJTzh0zS21zwHpz/sjH
zPFwiIGc/rivH/oELLx81z6Fi0blJDY2VKEeVt9BrJj1pQwWJlNte0V0DpgzeJb6zCXYij6pTFEa
2mcThVitcMitDcvXXqQ6g3Lnv0ifJZk0sErV+3K3rCyQ6VYKWN+wetXfdfTG2mAxtwEQnAVxsTZ8
bQggwkP3KAlrlhyRWqmuHnzwk9v7ub8lkHL/mrDDeLhTJn5mr8csBk7s/QRD79NUTH94eWvgp0z8
OXbBRbpeAfn8vsSo2Qdz0Gt4uG5s1T8nrlu4NrY5In2ji5StnbdkwMmnDF6UMC6d432aTNTJSxGu
dXl/7Y1RJKOk1LAzd2m7F5KEBAUMbIy0GTXKXAp++syfvKn6geEwqkwUyb16QxArxY08QGD/rOdQ
+y+lGgodk78hc6GiperKoLfSox/Ao7YN6U+m2w+Qu92pRLjPcSg96Kk6YpqJRdQ8Jdi5MK+HcRA3
kO63oO9SZmoyADuwVqlkvQ/mZJJZySBPwKnMKSeqMUfgbOn2jp4UTRTrnW9ewQu3Twq3H2qRBP1Y
uKMZQlBW2jF3UwybObZh1DuWFXpQlqKpECGItcnfWDB+522O8GPtKiVg2d0nUz6cq5YpjQCR4W9Y
r0QQrQNEGe/BbGC69MBqDBQojA77PH6m6yAWdDP0hNbPbWyxfNMVHZEj150HMkHhY+1ekJ8/cDFv
7CKe3uuGb3C44i613y91xScMnkwI873U/nOQOiDeqKhvhcudc6qbrx4uY267Oh4MYLo1j9lgwqZL
lR75uui41J6NVOn5kGl6hsiY++6NNiObQ3nMrT/WSTve2EERN64wKIbmnHPcWNqTmAT5iI14Vjyr
jTk78MV4ZEubSdvI48j6rqV7MzxmYoG+eExRrFuWTFhANfi3j8o+Rh3/LVDCP7E7s4xyVo1PajRx
jOv+JtY/BjRQawsvcUL6XXIofEKd3YMJmOLCI8KihsufByqnnOUILn49EWuZld7HTPniClDrMKFK
8nC/j6GGP62ZQMA9rCoCbGrdjh/Fuqicfbli1TlU0UB8J1K4m0DD3yQKWrL1xdVEGWa1Q7nhrweF
WoS6VY2Kw4HYGzcM3mMkNZKUwsxbRKYuIetkh1SY/gVqTTyydyWfXSK2Q/KaOdyITj85d7AEl4gH
uyMxoioqXL4B+j4etua0gy4WK3QHdODuOJjzLcLJ99N9UE8ViXXeOAabdDQUV9pVtBWQiidTYDJF
/vlfhhJpyc/OBbO0igaHMX/oHQ2+KxnAEvLduBIhgqeD180EerbOw53Rl8Yb5TyNylWtrVOacJc2
2C1P6K9xOoPmnyePgJGpL2eSMdfVGIQMOQYMCUR5mjkQB0ymtN6L/y8TVpV7NGbRMgYyKR/GcIZJ
Mfivkkt1uIlrkWI5KOptiUBXAsTTet3AJjGkxJB6Plre/W8HhqpOqRXz3Yx6F8zC4fncjo2I+yMj
shklrrqntCt/xc04LPIMrGAUc04l6/o1Mty45187/rxmgi5y0pW5lv+EMpE1m46JFioW3GRKXfho
MRJbGdRNSlXanY/tKIj1ME7zpAfaiYYsHkpoiu+hHgbvDRLqJJRPMpVW9IVA3BzmFMl9JZLDdEkX
6+fWypNedIK2MpVIFfcvTztBKYNYvk478I7ubrZpFnQQ9OeLwcUe+lyMoFa4go4wJolypNNVgVFo
dgPla5RTulIkNERvGSXaAzM2aZXA61Cw8WwYcUf2mIy/INrYCirQkDfaSJfBxrBCZVPAw1PzBpUg
W1ev4Pz22uOutnEaPWajQV2zV8TFoiwg2Xj8v9vz3FsSC2RtlDeg7EPnCJcCv+bjgEWmjnXGm+02
1rvYF6ErCREcD5GlY6ltsfAn1lIzxlNw+SQNOdNjtiEQxQHqNLIn4H3T5l7ctJD6rfhYx5dRBh3Y
mxSbU77c+KP//kl+n/BPmblgb0woqCbtmGIZ3XShPoH/pwrKhyx2m3dO3U1U+RBgE6hr9sqAhepY
enNNoR9vCr9gBbC3dudBfs8GzVM0MTNuG7ZPvMKKhQOubhDWqZVataX0Dgv+pfJupYi7FaC02ldx
oiO+x/Lacfi4g+YPUP4hHy6DiuELM8O8Dx4VJP0U+LX8E9YYI1gLByXlD86+HdkSw0Jy0rLF9KYT
EUPXXj7asnDTKUmYXE3E8BrWyZwIzXTwdYi37wIGToAPwDPkM/to7R4OxaXXasF6O+qxEv7hpIcf
u23/xhcYU6Ca1yScGU04fBVQKZaZVrvnkboUlaol1GNZrh9kqe+pTYniPr8Gju4fsz0R5X+3+rpa
UstSnwS8GmkQwU0HBGLt7CKBL436ZevNSYIPybzWHij8Dk7N/z4at5ZfgoscrkGTbCwGtvVoHaF3
OL2CBbba6P47dlSRdBfiUwiorHH+nJsz/RKuiUZPZ0EWAlC39lCmkuWjsR6C/r6qMmlMuoOfn/YP
xbPwuDBu5OGZwl+huaVg8L6rCeTo/dnkNw9iJbMrWzD603FuIwLbGBLLDKsDVUjWuiWkbBua/4Lj
TpVDadtxGGze9DKn/mH78hT/nk9caIzNcALAlttNt+8P2LTjsKHqF2+5nqQnn2+CEYj7AK3QPEIJ
mU3zYhWL529A3wfCHE/uhL65E7x3GZczKxS9Ys19WGx7CLNClVjJG9DmxOCCdTkZcooNtYW79JjI
Kp9FC7ZsWtWEx5gSPOm7rn3irnEDSfl06qRqLjdXOmX4VHIhU91HChbUTM2fJvL2n28tXlU/gkWU
5quNyCVBpLWU0Ow0tNWlb2F6FGnRckSoofxryV/j9o3sLnAnc3LjzCyI6+cYAlbJACR236UvLes4
11Cyq503W0IvEg4VXgNjf6xsspCGGOCkBsCv7u803N+Wv68KVD0U832S9ClOcXQUQ6giAeojFug8
JP9i7aLuzWUCnssO7nqsiq9ruJG6a0EE9mgwnDTcsyyeL6kI6bRpufJ1E93ZivMNASDBUoFXI3j6
bZ53YpKwPGxhVanMaCgUsKr9expfONi/IT82rhuIRYzKEytTA1A8tkwkMGP3k4IDsRrsu9ySptvp
70OoKpt1l6wBg5opdQVx7xt9yuO/TPCsxT8dAfdQ+WGSG1uv0YnmnybdL0G/wAfw1IKvQdHoGoc0
7skFi4aSbmbhRzPBKQhI6IPUcs7p/2g+nqFv6MXfUAqXGfcs81ZC1SleFJYMo9ACklqWixRXg3zf
F8Y9AWT2RIVMN9Xx2Sacp9G3grP+ctAYI1GI2c7xFqgx4jOFc6AQqIs2GS5zYibQL768lekUnToX
t1BIY2cN1cuJXBdtcTSgprXCspzqY5WndKEhcdPANBIkQ2vQhnNPsQGbBjr4XptJGmriuBqqFCKT
TJ8is+trppXGLxIEHSKg2KE32hqnWuPR6UR+RfKVirSNc383WI6ZcaXdqg+592H6oYLRjR785OMs
R3mHeycyScbTxfFPizdZFKqNjJGyPh6uDYE21NxAfBkHwSeRS3U0FBfmP9JtWYneq2MuUUG5oZ1A
zwIjOb/nEsPuYJjO+fDjFx7YmaQnUoWAw8AEtxeWVi77sb8bNEORoyMpMLFSY6d39SeMRoBS34oE
f0poxvbWNDAE0lKTqLwYhH2OF9HgdVY6TvIHdaQj7rbEarwvRsUge6mHfVppPhdnm0iGQQR7Q+JX
q39HddGmD4WoAuU+Ei416ARRAk1Pn66eNZ7sRu+aSIRM6WGSokSxyRnYdgkdYORwX884MNTlEeRV
r+DkU+8a9TQ/qvJGl5vo7RYpNsbdzk53n4M/FEXyiARkvALNEmimOagsCcTJDLZaY8XJMPm9ofte
tKEWfDGe9YRjWajMpZ4ZnCbk/S4+tDc9aEccfqlHsshwibzXBoXtWP+g3VQUh2/eZlcZrmGn9lWM
V6mMIfpe3cxuCykaodVDPYl7qR6j4WuK03EkDOs6iOBICOtSwYzor2kGMdsVgPxlaTaEPEOKe6/M
xzriUtTNauhPuYXKZgyMolxuiyCnPoysF0ymKQyD46fGtH2wPnmiON98seLrwnE1C7ty/YSbtOuW
zPTZjaZzfTYhoVCtVmjOq4DfXL08ZF4QfRwcPmnIDWlnf+cW7GVCFhhWK7ekbhRaQT//V+WyxA4T
9Kp1l4iyZzVFVynMTVRTf8wyuB8U/QdpUdSCvOeSOrSaTgGdo5sy0gHTu6QgEIfeLrzmo5Y4IZOj
xvXHzUFUuEfxfIzhez1h1+mbynD1YlpquxfnsfDnMqLjcbMdjaNTAmFqHS/daDd/cVXJkpPPogps
zuhfrn1Ldhufhy0GqZmF2t8zDPH9nVe80E3z6yz7YEBXrjAMDOM2QLXYL+7FmmyQ1IB9fxl2nHv2
JlQSQIMipm8wJqrEbTlbrdEwcuVD1pg8VTGkg1zyDUK66lWxxd8Qw8Xb0/3ceiur/nuoagVANa6C
9kp4g5Gac8aqQ2w1wVRof7CekuMni00VhykQxGJA027YbNG1BaRndb4MP9vVZuRNhGV/ZvUafsTk
C4oc53Sh/g9OvCAmjdFVA3BANhBR/iXj7f62ib7ObTAVehrdVMceTxTy6E3uzzwy3Nt82/PWI8dt
vSjFFxP5lFUiBpUJtAqfRo63d2bIiOvkhA+FNbNV2QQ2GEBI0PYH2/v9d+hwi8ad6kjAfP7QQ7tN
Px+d33M6/nI3ZKBrBo1xSXCm8xY2SKScgBjc3htmAxMu34JjYxVzLt/QtoCBSTUPpBfL+BV64O1p
UJ4My8KB+inGboTcVrucklWNMsYzoMX8hgsvBaKA7EJKihsPGfpG9aWXlJ0IjKr1V2V1NlgIvENi
LK+06iP/0YXGomxy1dEuAXfqQReFxQTJJddRVhLAwPa4+7piFV6HU+hrvatOY5K3V0jXRK3y6834
EZYL1CRIJZO046zZQKOSFQzIXDB/wxRb5eVERD6zSSffgnGuznOTBR28iuGed+ClMf9Kw73RbwoW
pSiZgUTx8XM0yuC6WNGfap4wJWRW6JU+4ozozWiujBRUQpwCmyPNDJQSGKTOwaBrVQCO/QORbBCi
gjBwao/czaoKM8saiEcD1KmmjhwqoRj6VVtv0hsRdhLMIEb1yjSb904Yc0xwF384IPo/OY7z9Uy7
wXwASgsn/mi/iyiiVOE7PQ8r+g3bhKNpsoYBla1BEWqB3K3NzXyCfDtUW3Vm3PouWRgi8x26VpAq
6j5jbMrs6BvahvKvZoY83B/aDhEPXpCaT/V/ivPXbrqpUEUodJZSONlsT+xNGqBqLb7ll48PJYyv
HGhHqHo+mOytiGYqss9QMUFl+2itymkLDbxuydcYfpdPFvDVWoj1VKjCJRgQ99itnsOXKM7/h9WO
qcFn2T2FjWntlSvovhLWB6PtCheILU9rUdj46OIFgvQzLK5KmR16gwuGXC7/mygIqt3XrGFacOsw
QKWtGJwE5wrnkNCjYpAjVV6Lu8qym8RXLc94sEZ8vLNpSoLTAR7RUi05f3RBmyGPykCR1F7tVSaT
qEYg+pkAh9XpOl0wX8+DTN5ab1v28aI0C4LhnWt6w+zCmXBStqLgL6NVkNsAPDa78zXQ0LsTAVPH
4g57u/ZHNbk2DtDWKl0821I7cdqYSSUrI9ep6wvdjAxl2mWc0+tG/wJvzw3WU8NqH9c94fh2vh2q
54ZRXGtvXHe5aYVvZ5Pdg7Vt7deHEI98u8TC2ihTQeYVTE9VbnfyxErnt5aUiKFRg+1LbRccVDXI
4JGPyEQHLR8+yaMdoLZz6dUthnuABVrI4D13jjYk9+zaZ2Lmo/gB2z+8b6kkvTE1xbBrPb8o/7Fx
sEJqF5unHol9q5E2XkC06i65mPLnx5pONia66h73JC5e9psPyMYG6OrU+qvvfq7zo97ov7PcV1s5
rxm7ifSOer6yjZscxE+Br8xCcRD+M4Z0CHlW+7QhwagKxfglCS51AhQklQOLmdTcwfbP1Ws3IF7F
NG/2K5c8HMcs5CkFM4z/RB+tiF8E/b0mGGfz6x+ALu953/o1WH33wPsaKgVzNnasvptUQ5+jY2EG
IODSmK0H87sGdcQpzr/ZofT8XnQ6fZZJwuS19yCPJLNTN28Ky5w/Z0vIkbKjEo4h3FF87PEjg8Pl
k5ShHr8CCgYps4jXqkLxd9nTuzRrABKRVhcWLuOw3Nuf0/ytIP4NKuXi0eUaDCpt0oWWiWSWwXy7
u2Ktk+gYnQXc7OdU3mdNj/Uc+qFts9BWFd6eSbbfxtJXoveI1IECy0a2r4hXMPPHg8nK3v5iFGGW
jzdDnmdDTCSprnUvMbbR5Ws+aMtykdevnlBteGg1u054/QnaXTB4rG/TRoMrQWy33XHrmgWbAZJb
s+m9dB/1eUPplJnaGi/77q774R1RuU0EdEBFRAELb+XO4wOeSZdP/HOttPXiY9f/j3Le9mNamqnu
0ywFSk+MAyT91gJtF5c/xHBOzgcg6xU//EYkiAqzmwLOCNTQl8LVixN9ybM9gZqQhpsap976Nhbg
jSEd1mLyjFdhHFjjW69Vrm7ThfsJi9LSPAo4murV655YavFh7vkFdWSQiwDOUzsrKfGfqUrqPGh+
i04l+yCoawhTV8VxcMJtk9R842zMfZRjNpeJjqIe2ADZjzbjcct4IUJtdemTEn0Z7r9Pp1JkXRBJ
gXgsi+bbC1Leol3OKrZsgfOCHkhqENeeEtFukrqYl3IN4c5If5dEzse/2VQNO/XO7z+AzrFBHAfK
XG3njJr/RHYqllYo95gSykPG/st7+fOcfluiSIFngLlAPYTxk44uPAyTt7Xq+7yiGDu/7YlWkmFx
iPDEBtpbHhDIpgrb58aW0gg7EN7a/tUiz73xJZBMGLYbGiCLMLQkIJvK8xyJjoABKUiawd6umQjg
tcouHPMpx+bMMb07VC6DtGxi04DlQDfHiBY4QQZzO8StCerkr+zA+oKs2IeFZiIYlDk22wJkd2b4
rdccPeUfk7UY6RpamN29dTO4LFkE5qW8qTCMCL2X6phN2YCXbTv4TU1bjG+17xiZ0x0Vch82wXY9
D7fOr2428c96HoPmY6WKNZOw2XN6lmpPqHLwOQPdtDXKNtVstk1VGzTS1uxVHNMD0CTUQ3Q5HOzz
Il6bpESzkxFY7IIX08FTNFzor06/tOuz1F5uoQixHq0+l7+RsJDHFQoqX9NeHI9A7rQtbhYNUe96
GGQXwabtXG9cRogI4EVFhYGpJ1o5N+AH4H2LakhZdZU6RvzWvFFv7SvaPfrSlQFXEKF0xPm2erM/
do47y/Z8r52SlYfCCLHm+JiP+gKSQ+2J4PXP3sWQ7Q6vhJYgMCWLojduYg6/X28BVmF+S0LGKygv
U7scDds5Cq9DkW4BbDIkngb5EoEDbjoRXLWqIII9VGbGP9/+pNmNN6+oXIg3lP85Dca1qB2c5nXh
DfihTouNRRb3HQ0JmR/IVNLc0LMR6gdIH0ENchSRDGRAXgaExYI7K4MaSAsrawNfO8LlkvFPP1MX
BI1peGzyFp2uFgPtNd966UEJagqPNmrAO8ntXcJ1VuRI4YLRrVLGG5zI0dZPM49T1AXqfkesxcia
XaqbIda2RLK5OSXrr4s/DKdaqmJGmg7J/FjoSn9qitTqOgd8Mc48clAVeKjIbVA5kVRQi77oM23Q
/9PePu4N6OyuHd0Do4BHizmxiQ8oXqY6xwqsrxit33wk5ruIofLSFlvxIogLNEQHvrSzas2echCJ
ax6Iw1yM2bCXEYpn3AbNVA2dtXuIDRo0EjrJGS7i67RlAZMKHNROGJyFXS/jcDHTyIXuVWwu0ghz
a4utLFFFmzld/VmB49gR5+dln3wAOvP/dG7lLPjkU4nez7fuUONM79qykRFRUQQrYVV5WWH2P6pP
QU9jpdWbEKPPjL4qzL96NK14Opl17p15iDkIgOeYyAnMu9jU9yxoR2PhDwKAOFJYnBfeeRYJh/+D
akQYslqs0zSAcj1rPCBVuKqhWqVlrMENIn626XM/ek35rQwTZYDBsL7qBLholNz8P6K7sC8NhEHy
wAKEtj8rfyBeOzAIASPbd/fmQaMOWzzL9XTfxoNMe0YMa5/lOyUY8RVKUl9E+RlJZ3tNjJuA7bdg
vUtZ86lgxVDdWN6tqXUWLcTPDlQU5QCyYAdl/KBDNv15gB61I6P8VrXZfBuV48wdvs6TfjTxSwFR
63lzeT/8vkdLh6luQvcth6XNf/VNpOWkOONcxgRdMjxyqukwy8iUgIU31OUetmiiLQtxSxhG1GIu
b5vzUmx7UYo+H2MCnykGfDE0DUYYNDjzQoMQ5ViuFqiQ14XdHe1Nj+awSgdtaMn1BxxR+8OE9WPd
C4cyMq774vO0HXbPzNJPDb3+jPuhsyFhPoTgHpBSOS+aQKTVP/EPjUFMmlPLZ873LsmbtL/9f3Gu
uGs89VbY73zFfRiu8pcvPrOlugpQ+/GDEJexIXb7zgLk679/Kdvc8N2YxQiWNZ1Q2wgyWgCxg+iU
J+vkkYkChr7q+2CvYfqBSetvh3UV4kP4zUg84XKYW3VD3H9Uh/+UmS1RhO5yRzBplrXpEjamXKSe
/ILGxn14b6Bg16/oALfCzVM9gldbR4MELASUhlvbObmtQT+uTth9OLVsh54iw4WwEJwyUsj0AnFC
+/R6jDA2H748IbHaaIKesGNT+fvJVZkb6Oz3/Xa9JG3D7lAwMABHvej30bKPvLck0YXKQ894boYd
9byIN4r/cVBTMxqoHa0Z+7YytycfAKcqpI5C9YC4j4PMhDWzpKT+hmHHzTDmUwsAd/lAJpVN6SEU
S4x25CiX1UcOvbfDoyRXUfmgEbrF81IxOIFTpy42ym1OcIlmqCf5yY6PL9uUqhpUlW8Xxf/vd6pp
jJrPxzZcfugAocx0CYPCbucxQB+hP5ZSlKjyoQ5Dp/txx4G9lF0QyhBKmrI9vIiGKHQmr0fQ2Ytn
FNRTySfknhQHlyQZrtr9i+TGdk8qKAm6w764UE6kcSBWPchy4BFJmGQFm2r0NALJPd55+aCrwUeX
CIKmS/ri9BHBGSBA9Yf2tacujdndPpm5UqIiL0TNhwxWnKhHNT+FaHolwbzXtO0V1zfwyty86wzt
UMX4Cw5dBN43Bucx8q7v+XoTch0e9ZsWFwH20R2TqGbq3kOdmquEFY/mPcJYcXL2cr3oP45W7zFW
ZdD/5HRAGFPs3v5/QSgirIOMNodgDc9cOhIQXWp92w9ApUikI4DrBuZqnAwmJYtJYzk5AX9zU/Yw
jilso/hakrQDJvJqKgnR2o8ANEVailBsMh9BM81hPen1FHUT7We8nbUIetgn2HVIpNgUb+NfGTD1
U2igwM+Bgth4K39zqW1XgTtDyntGF+gAoLNRKwLv2LEjBIcCitM+GTZ5qQrDgpbG9ZgVw4CC6X3A
FdkcPcdbt/cze0PXGHUHhlto9aA6fre88bsfw06ZZPY0V0sfrwueaakMsWVSZSQ6goUP6ga6xlBw
bAnky7sdKFIp+kPJYhlVDyomlOqv2MJDR0Y1+Yu/bzI0AJzQ0MTN0qmCmjDqX4zo6gx+vW6JeT5L
wfW/qbeOZOutK6ygdUiACybvrFHo2jgPYx6VF0AkR2vfDeOFbe5dh7jInUZ9MrkT3YYrMa3G+r7K
UdHeujssFmyTEv7htjq0S8aA2Kv8SjqF2VWEghMe5lcEs2BDQ/uNY3t6E+impOw0S4awzKQZT9Ac
1aszHnaPVYoxRmTkDRksb+mekcpt5KDaECpMllW4rRhZRXYuuvncQm4oLzyoPVZSiH/nvjI5Qrdz
b5gFWd4G4jh2DeXc1f04gR38e3PKqerJCr9NHvIJhETIiB3RZaPGTOwxg7P/YG13VgVkOwHSVCQo
qUfoMhdQEKOiI+wQ5CY4d1wtafZzyVdlIiz+Bgzc3CU3ryycj+MgmQLqWQQaI9x3Vn91Z4zMsPpG
g42L90nllKOZ+SmajIvHamvmBFzOS9OcyVc+0UKLF342oFmnqD2m9gKyNamtj+NZ69fEwu5aTjtQ
Zfy1T/rPyv5mZptNSiRkqtUvN86Bn/LR0pWAaFAcMuY1AKYCtV7H5Qitga9GYGDc1G0J4R4ToEbH
dX5mX22WByC91BGb2p+jyoTgc315IexqZs9SJFTRztRRLeb9yzmuQZGiUdIV7WUSTnhX8ccpT2ZH
5MV1vI+T9qDtF8fzish2a3PYsaFOiDfK+MsIq54TU5Kw1CiOAMCWWuJOuxK9bDPqZ7cryOwGLQLi
R+Jdc6im/aSoqrcdqH39lYMw0TH1rCpZ/R8ZzBtL76lRTsO/J+jLaRtsdr6ImkYBKlvs1lxNPjz4
DBmb++X9xT1bVNZZitxnCGNzwsf7KV37LcYmuQFs27FvxQm9dTPBVgc51rdzc+hPvLeZwakIz1Jx
zpHPUZ3OORACtAcG3LtTDtXMwUFM0r3v6l0+Etqe9+qKwwF5sYAKKVZJrpiXks5wk0/AfkTHatZo
FelOxtZ4Y9X1wAdWtlia+rHJgQv4i4y6CDTzWWapTpr9yRHfKLli453CpxriyvVM/oTRJOfE2ZGf
KADdC+ATl7arYVQhZeoniF8op5plwCKoxMUQd/gZPnJE9ZZBQEX410bsGk8YTmUrfiF3Ew9dkXfo
Gj4hK4MD/NFaXYXV1xVRvDDxfw4uqzBYXB/+kioOnGBziasW5xkFwMekuT6UAIN3zejWJE2Pxu7D
cFC2Ky7Ais/E2EuvCgbbunVr94zXheThdKdeG8cu/wQjx2GtCqwQDg02DhNSjJy7ukrYzulrye+c
OlA9Ay/m3ux35iaKxPqF39RHCp/mjiOr5GvplGmxK4fGmNp9n4NiwqAyl1eqruhUus9RX8CL5RKt
QyS5z0SnZOevS3NV29yaUn/2xRdMV1h/SXTVXYUJVCkf++CvW9vqEWLx3DAoLT6VVkmlbpMqB5UR
6QpLShP7QlWL0y33TZbTaci3noDd0Gil7ifeTn+k7c4/UvnFUSiHFFmvQgEU8NCGWhMEOD04CiWN
eYsJR2ct5bh4U3rwJbWa51ISvPdJA6vykcwv6WUwbO+MflZgeabMhlMFxZxxputuFJPXgHpAvZ/O
qpRQ7GiHsOL3PT6yqAOeBoH+SaH1eYDVgtEbUSLkD5g0qn6N0X4oCUbBTsqmmCIwawjllOn6o0WL
9VqHcG1rJueznxO1xW3SfsfT7fMxUjIWIFqo80rooe4Uy1aw92P7NwHJhwtMhxo/6ut/9BdQHOkS
QEvwC/EOfKpbP73zjRkUcW/9+dTUBdDhq5xi6gTux5qjrplxz630nCMP7Q6B5+dsJOPhWZBux4V1
ZE6WL5uDlheFL1FJu+BqnL+O6JeDxtTZUpP1+8ov+K340otJLsLL0fbBA4VF7FfpvypMKmiGPlb/
jIkuabc5i5xdqyCMKl0RwPGkzxwcs2qcjwqwHkp2riAFGwCmL4faeFcGC0djv3HU8qeNHs9XY4tA
XMg6jUnH2LRdIPfg58MgmLwEZGJQkqm2i2jWjl2xI8c3P80vBF5HJ0SpbTm+FqKpOMGVjpXDNi3n
4QnkFqnRht4Q06Fr2ESUUn4n/g/U8Xp9JzT0pQ0iAmemTSFMGuJ/nDoSoa6gTRzi17uenAra4Ru2
d3D3mR8gN/jXWyjS+q7jJF08fyrJeWjgY3bHGeh9UkrvpKQyA22eyXg5i/a8kbPO4itgI6uplnFA
MgEiIR0EYaHYiQAcQAlvDodME5Ni6JiFvogA4mpk4bOySVEN0TW8yiPmmk0Xhp2m54xdIejs9vBv
r+fh0kQUGMvNVXXDb+Tnaj4DbOKx+i1Ba7jVpQ4itPb5RSr5LGa0Soz4/4NM82bd52Kq6zLamSMH
9TFlg7MXXdI/iHEr9SPaVW9PpKqH8tJxciwPv7aFAEn4sTbprTM1MhhvNSAFUa2ZEQhxwhh/saQC
ebFdhhOjeeR4cq7DXc0H5OjpmjR3gbxt94FLiFis52YcQU3PmLLLrBPyW8l5p304mGI+e11LPXs1
12CIj22zjs4XzdgTo7K+oZOLw5KLvmtAfsltkHsyLXTFbPWdoH6Wel+n3OCGe4GxgWm1UvRxTxxj
UfYr1MnYobfmxNvnVGlMz8kgDjkVvtC4ipjmi45RIwPEMrATTR6SbdJODEbYO2EgIThDq2JTOXc6
V9/IsLgcWn2PHvhYY5oO/DEnFP7y/wLkgey+NXqwZPbFboAB+CC9F4Y5ONSqBb6WNY1u5G2LRUWv
odCMGg1Mzp8fu67zL1sTdYEWB8yjQG2Eoxs4bbnkWecJBmSCxa6KQaADkXfTn7JApYUv0PwvvkQU
FciuX1ons+2vl/J2C9FX5hXOCPIZHRp1TCE1q0y3Co1bExAKM6Tthn2nGt5OKds3/USaSny9pUrH
CwTs/qQPDphgbvhJnhDAdtPxE5G5TYS7XyuAYJAATkzvLZR5ecXCC1ytoHDO+X3ff1F+0kZFvwpa
CHegXVdRPPWoEejliaT/l2Ndk+TJN1uKMHeu2FKAMzxe4mhSKiN46B817BQ0Genyjh3sNOSu99aS
E+DgY7lrNSSlFkiv4t4/pcN8clbANIEoTYZeJ3bO07aSF3n+pIjlOr7V596dCTmUoV8da6FiEeSD
rFABvLN3uGfh47VaaNcG62xQ5hGvtTVK9Bz3HhmpgbIdzxm2ZIHoSgc3fl+JYxIUXrCcDvR7clkB
w7Zz5dFwQO2NIeEV1iWj2rRQDher8Ht71HhK7kj6ECT+J1pjuW27UkGg948Di6g+MP8wb7pToBFv
YMyLz5wN+K+QLEOEzmD+mzmyRf8FczKwYPg/cbhSv4Bsoi8CKdp5zoFMqy1FBd37u4kFHf/UaH1b
tjrduihNP+PEL1rIwI27q+3e2/nS0F+MjYk/pTK0fTFGl5AgD79MYCoR1ATy7SvjO9NSLUSPep4/
j5BN4XrSl+OQuCUHhjGQS3tuAt6HRJzvnc+ISKS+xay7bzhCWgzFWmHYRvBOJ72sqhGGUmYHRyaA
X775UxSkRp2NkowD3UXLtfZ6ShKikXGBG2JZWQVOVidoY2WYsA4uIaynOpy4D1G7FDsgaX8gnDse
01ENCcSwySkZbE/yaPbZ+XqZXzStnu81B7dNsKMnp3Sxt9TSmiI3EYglLGzogqFfuJU49MKQAMn5
65r3/yX/3kbdaztIPAlGKwk/K9zxnB6s86JAJkqvNEcU6VxP+iCgIAMj5X9U6I7GBiAEaNkKEtbt
WkSAmK67zGbtD/v60fyai2iBtX391jTOCq2oEstoIhmzVz02xxwyAWVa6DGupivvzS5w2wRZxSoN
mS0PkDzhlTkLX6ZmErEQVJmFJU20bMiABnBEz5Jx4qrWa67kOtKhxRfTyTwzLG3RV7kZoeFoRkRe
m7AFTvEl+M/02B2bVC4/OcLf0ikNWBKFQOSniDCXlZWQyy2YAgIrZ9+53IpORIaJgR6zVnyNe+Cc
4podXb/caQrGuCfj5i0c1PC3yOyuOTXmOlRM0uif+zNLkBIt3743U5rL+wLIBXCeghtsf84GC2XU
0kV1w2+JIyNiNNwN1lrTYXLMe7egMnKxkUKlPY8n5VM1XCx02aTBt00zRzrqQcjEJa4oWdGOZwal
oy+tq4iXkoa3psBxlmLcZb2j2D5Msl9yGJigl45zfP0QtVF6zuteLoLXTjy3iQyjaPMY9DowUGcM
TkJPzcvUs7N5w2E8PcWLXaPCavnwdF9p/MQh4YSunX0S8BTTipDrBe/ZTODyTWTJN9RYl3jKqjnC
GVRJwzH3/Qw+ujXV0DBelGk5NJiehlxBuuSOiVBvBRGAr5r9O/WFtNp7xa8HeFfs7j+VW49p/oYI
h+Z988H4c8ZN9kW0wna9JjlCIUZTHIF0/pxQwYxuq3oQqOIF4VBCdXHJiioONh98W6u1uvGV6wLL
DRK2a5rYx/JdM0xRL5xyyTN4nSddQCMYMcojheD1ObStZehz92LDs59ZBCShNFVkL2SVIGmFzwei
OWZmf8KLXB2nHnjHvM/iMUTDX+j5XNaAsDQKVyj0uwlqCG9LigPgzA1tetEbyrHdg638rC6Rtqfi
seA5Nb6CsXvAtT4qljmhHhkeCEpjnFnyLcjbGXZHOk91YAKTixZvXts72JDOhVoFW+t38qCiev/7
QEP9fwr5+EKtorQ/pKndTbzNUxPL3YIoPXAr8GY0nPZE1nFL3XQGhdwbc1IlF5gsQkRDtLtxvAf+
kqKgx6WHHTo7nJEPr5ym+9yxn/VGQpjVaaDN1m6QhWCzp8Tn7b/r9NPJV3dyHP2jz1IfgNBcf5av
asMK9nqO5dDBctShQZM5hL6ugm//IN1TTfnuiWkMKFnrmN1CgcvX5PCnY3naXyJDq1QB8tLehtKT
QGRTJBNDasVndIS8ngmnU/t6KWo0sQ9ACfgzpc/H7waMn3Jm4TVmFaI4j63YEHczWb56Ke1UHC8f
eHb4AqyBRpW9HBYvbk4VdtISpPvsK/CSuj7Ie0HbwBy1J0eW1u5p93KIu/fkhVmDQx+gLVCYs/Vo
LCjZQ/tf3/L/O6VmwHuETWTahUqbb5ZQwpA7ZBnKm8wNSKrXYXKT/VpAzJEKxy5f1NLmA4PgY3lV
iQYArWP8gImnTBZIgyHP7qsezGxTdcl+W7v3INzmdCAk46bJMNnaDQbIKEzxP4WIt4BbHhMks8S5
TqYuDcYlmJr9vWF3ZTDJJyMhK+NoLSW2pSFEr26RKRZbOA2Brc2FE//7zQCPl2V155YVedekXfTo
S1YutpDCmgMuWWH9RJRlblx1VPPtln8av7cj6m6c9W0zbjvP1Ob4cYfcG8XPcyxUs+MfGiP8TsQX
Wr1VVDjHove+K/Q6bUipkOuLlUaVlJX3FUtIn2T3xz7XJz2ckv3BdAn5fgApgYuIZFq3PPTIBcAJ
zhF170uE+bBQZ1CX5xYcBPVBAra46R4S7FI1A5tXpfw03wDpCLHmj/lwcWRkgfMld8QWn01nzvHt
gxtRj1W6Y7AHEH/HoGa3DY8hzU7QvbQjQqOImY1StYwG0727vYMHxmG95K8hlli3cGe4/WwNjko9
WpX4liwJTTf0Gu6ebnwhxhhmzfDzJsdyUWIDNTfwL4ca3qLyYTB6uPKEO8VVNuMDMgeFEm/lGe9z
wzn+fG6KNJbXdUNfeshgCcyu36/AvHu2jRT353ywEIM2MROMdIQX3uZ1XRy3D86gaWSgbjbrCbst
VK8JFHJ2x5er8us6Flf/yfXSkEcIYLtyOjQaSNmVR7AOpv7bpAWFkVNT1KuIVH+nwQfRY6emneHE
6zJ/YBBGffV+lBZHla1/ZzInIZSrvwhsO9eGYTwPVqt0QvjAY8U7ymy6V6vuv+8/+dIruUo7R0Sv
KTTFioAtxkjUiasi+EvTvT4MHjFcaTaKXzm4whzZFa9gOFo07eOA7ueuPXwUsWDmqFtyodu6PypK
Z3fhcCciV/QBwprGbtzqcILaRqsFvQ+RBJD7soifvxcW9NEB2m+xQRdfB7BJlJvA8Rw3fu7M4sN7
LAgenl3XY0iB4Qm2It/WMDU3ww7q6TTybMz/I73O5lak1RUUxaF7hTommFg0QmBlpXu1KURhEQRL
Fpnemd3FEoKetzsN7N73aPe1AYlHZATREeZL0lbirYALaVZhGfTUr4WxjEpmXs64EOwYtKhCZoa7
kSmrlNyZj46XuxuE/QnEWFrp0i+TPt6KgdzmuM8t+PgwG1/k34u/RT3SKon+w4+Ct/gmYDTNmulN
jO9RPb0iIpmm5orlEqebyiYjg6SsGGZJSb5gNWNehYNhO1vYYaBVYu1grjL/dOcwsBw7fFa7ECu9
B++/rOjAQL3ia8OWiuOd9ys571QAFLZHqNkrefjt9TzonIJ0Xl94gh0IGwJMh7wbIcaqxvO0qN40
756Qegun3Keo99xh8YznY8DCkKLO2KIHvwZ77H2gUa/PoH/UCgETOEogQkPE3K9n4rQbMg19hpci
YVk1UZgOmtBSIzOb38XgfLtYpugIQ8EHpsbcsEcTx98jWXyMPl4AJd15Bmx5ubquexDqMghukdOC
H85R9lMVzSQNoHpRUqmxhegKSfA2c2XCY0ZXKKsSJBPH7/IFk2oIvMbyM87UnN8bYQOad6nVQHSX
0yjvEKL9hdU9v8ksUqpiMGAB48R9HAybAywKwB+h7LbY8Lgu1rTDSq2/cge/khMPE0OBy3zBE82g
0f7F+qvgBSY2WT1ztH+n02cbJcUISSIIE+mFG3H5i1qjbt8V9N2loYXyLp3edn6kSNoVAGpVOWrn
cd08VwUHKdTGLcd+3JLHatsdt3AhZTgiQfGTxfcZv/xRf0UwxiNa80pdMq8IibFevC3ze2AWUUkM
X5aCkY3T2nNmGaWRBcwu6BHdb365WgRDVDnur5IQwK1qo/qZnibrWjPDQxpdwQ83xnh06Pn3DdC1
bNunYz5WDBKAfWisi5GWOPvPPGM8hS5SgOs0ewdVnEP70xjgjBeWMC1umQZchn8gwhv0l06W6GuW
DILz2I6U4RiticS1IskFK7UauBbP68H6MIKOp6bIESqVSY3uoTVwqStjFC4fxacjz1WVhq+6rzzL
4AXr9KK+0ct6LX9C3yZ7f8Et4FMICnHSOLO8KnL3LpRie//c1vu53PJV+6EzkxXOUVih1kgT44XH
VadMQKH+rBjlLpFeNXAThUNJk9hK+fJsLJrOJzPSwgwoSrYsdG3tB6dLqEi3X7WuVY4Xjr7aikM4
5Ly/wYuoRdtTmEd88MbkCijclax/jF4Jmae1/CU22SnVy6JdtlficOGhZJaMdJ2T2HV7faqFMatb
htpif6g17f5H3QnnmATqDV/6YPoc+/CSfBGBwLYMhXr/sxutF126MqgmSRVKxSmIBmuMVdGjJbwm
LHNE9nky73BYofrSOvmtjztl1TdgrodgaCpGLS6WNNPyUcsbpXKgeAOlpDvekbOT9czYuxZ9OWI6
M/yAo5yCoMOS9b4wABHo/sCr/WV8knc/0dYlhspcA+msa/37aAfefu2Q1sg4+WAzdcxm6uoIip99
74YWOLxsjFw/OO42Qkjk+FAho4ssQu7aHJNP88CkFYs7AE5nlAGbYgcHF9hM22dwUxfyD/zH2F/k
MZ6Ki1/0KRv+HauX+nmbHE7PusEMOcO6U7U2CwTLaDSibQ/3Oc8TMkdW/pMKZO+j3c6WaxNLAoNU
EtDBKWAfL1HyZRRJIwHHhacSrebLbeah5iibcAxn8D2hD1MGKQBHst8QyDH2aM217TBdSXJNx2n7
AoKV/Jjek/Otbzp6iuaguM/tZy8K7RRIvMjctaFxPVHuiHSZNFOChaXm6mCF4vsJAiMhhZDmAJjv
4/N8HV1U+QrI6P2bH+7t2B49qxfoXN2DLpqCNnxOY2FmVWW15g3eBJeUcJYeaCSOHwqXlQzd4G+p
XDhd743uFgIOj1ewWRCeozbhLX/ra1RJSHkqBTBok769dnRcHMCqYsyOpPxqD5Xnxo6RwPNrzp5K
8Vci3qzzLW/BBOVANUmqbqPq0qv75mPa17aaRC+z4jpDmU9zXZWhFh6Zuu3u06NWzFRAL5rBodUt
nzQ2Ksr56g7vFnuMltFeDkvn0HjPOmiaAD+HTrhMvl6JYYcpX/H3HYKyMG0raD2s/pNdy7UiftZ8
lCjhYEMCtYERO0LntCGCTt1GBOeZNoOtubwUqpZM3Wy57Pmp00ZpvA+M0oyGnFipsNvG3up2jjX0
SCgYCtw5LA+tXySFnGdoWVTICQchMdz84Y2pr7BNvxJ5dNdGLUBSQQpdIk/riujdBVAGyrdeHsgG
QW+aQD6+oYdhteYtiWtHgnHNQINMtytBxUCykyIKcSAaqwbcC3XjsTh/gzB8afj1mnUMN6f19nt1
iTRivw5PKXbE5UmSbeQ3fCQY9FunH8TZzCYxC9j2TukJHgjD+H46I0TQH+tgeONH6U/lgYLsIJTc
+zMifcI8ICsLRTcEJnouMM/zpsfO5lxrK/y1uQ6OIvUt9BYkTQsnbc3w0w66H7g8O5gR54pMtc2Q
yMiz3OFmzWXu/CFNzY+OKzF0v2N+BTxPhK/c+HrCby1PcI10RX8iG//W2/XHVSQvH/OI35WToAY3
wGoq0nU7w0+1w5NPD+2ANBpOxJeE+Ht1EyPtLi4BVUbi+A/YAFMwhCf2HKumTDkIHIQm+21QnqMu
6SH2k4K91NmYCxNTDK3eq6SMl0MJBT4ekzXPkSclDUz/hbicQrVFCAWmcoaL4xq6d34rSJtmvXxT
bDBxUckV+dZ3vdc+dT+/dR3FrumtpWWhko0XQReRF2UbzYnXBKUjeH6PDIosQ6tzZyWo500qc2K3
0FAQN94sc8TOA9A4kM08i5BSr9jikMdrEbL9jgdyWPZIOABRTcHyes+RJCm2ygko0SPeF3jKgo1Z
MZmuWu5REltgtVWRO6VCAkstbJwtE+jGNvdFfWqXLK+SGst60VTWPSjz6klekKY3yP+h8ygrFolO
4W9iYqRrO5TSWGNqK3OqyFFORMubNPft85wQ51r1kqeqTGxBn8MXaUAeNa/HBP2jw3OrJqOdCO8E
rM4TAhBbRv2HNU0kMBP/mUuhXEoZ99tqROCp6HazhEgpSksc2pGQPvkKiau2R8Q0bdywVIvjTuI1
Owr0CnT4WvIq9P1rYIaaiN/llnvR7hd9vUM8Pr9toaVCy/vOmbpYZbezxKBoYLwdLfIrGrJE88rO
C7sXszTnyANBQjq2IrQT6Tjt0VqDFt5ZD0w31Q7NQEH/i2LxN0p7lalj9SMKSb28258SCayQ0NWW
I/El2/R1w4OSfens7kRmp0f6EcqaMMPOo3bFGPmpba2GPkQlJ//Zad3Oi4oW9AbCnJaA1rqe1g8o
e2A/xbJvWGa67n9c05dRSHCUbXZuF0QyDc12aIt9lpuWmBc5SFjN/WEkJgqJKxXPQN+wkj8URTmU
lTbM4bLPucX/nhK3nVAOPux7O2RvKUYvZhGDoqtFkzstsRBED+LgUuK04I/cnUJ54TxbIlOwxLAY
hm/thLkubY6FpJIc0rSYMOkw0lV3xc7zQzxEI/dO6gf7kUCdHQkgRXJgFx/pGVyaRQ1RJvqOn4Bn
ZxkF4qsFILvXgMcWTjcb5EzRMbZHkAfYMXjOb1lew0L1VaKZJ4yTO/5nudtGTZHiN8MDWdRa+XFb
DaRing5E2nwJaNv9AwEu7UlAmOPcmK/fAM3/+R2f2TFgjVRohijLVREjtYKA0JNlZ34CTDvwAYeI
PEGR+RaoB4MDqzMRdv1ZGO8GQmOCehPhqPYHhyx3NoQic7KOzfEO3O24Xdb7q+U4rio1JsjUcZiw
EXtTKo8whis49LgzAVz8Lr2O57i1ceZg2oUqkORCDYJhPjMxxSxB4RXHhywfrEvBws0ccMNtdbGc
CzhdaKwawB0kFYkoE3ZH+ay4jb+yZyJOYKPWOgZ5yfPnHdpqWhUSrUhxR1ptvpR7pY7G9JIAa78L
Z2AQAtk149E89O8zS8n/jJyvW4ap2dg2SktUDWXGBfWlqdNJ7IwzLzGjED3B8dbEUAFPqrrQVOAs
lBdFhY1h2DZdXA/INz0q9f5c49cZgfv+hjpYNvgxd4vNbQN/vCw5ANMeXHX6cteObVpdL3X8SAzT
fVJdhe5xnQXL6wwVWXBuTfTRHiCer5bCz0QL15qQjIaCFqMHYfJiFY+NavC//jUAe6airRDyimXK
ROuMo4jdFd4yEO4pm0eYqCnalbk6K2lDf0SCGMm5i0MpWJuI7crafAJJR+lDSA68H3p01yxn8RTq
j8Sq8+SxEgr9ClzZjn4b4+AFgu5I2BOUA+XB1H6sIAofaa4m7phtPAznDxgoibEmU/jWcVzH2NmA
qP3uGJ9XZ4cPljkkYqctfRr/jacHDIcadboqbpYAB3cPsKPtHd+k4xHBkYPou9WaIPeXtT5KdyyV
iDXdfffFebaNyXvlZ7M3fiTdNQKWKAa21AiSEFxDOU69lzhXByUhC6y5RCilyIzb9orPFnfWsiM1
onfcEa6ok10f65MYv6/bH6GrTvtPic0yBN5NuUa1cl2sqgo7jcKxg6jlFKr2r/9TkZzs+jwnAmQV
xWcXNa3/3RjDGYYlmFcC1U6SglQsV9mrl3L/lg4OQRrHy4vPWaL3mOATIi2Js942/E7C925IGm/Q
TKT+Zm2k711itj/vHc2vBABy5KYEox0SZyOt2DLKidxpkp/ZX1h82aOPDwd+BaqgHfdVdnXTDpwI
8RQ+rOw2O30n1MP5hnyPJRcdj4kE3emNz/0jYLg4b/KVkJbnXX/vL9pL6YWBQ88Sq9iTOEkqbkmY
NuJe+yCfjQvwH46vHWat89/PRQAv36k+bYvfMHP/1MtiO++HmyRBcomA3fTw0sijMaAIaPSlutqI
xJsgt9o31DVlIatuEnoZG+wsOF2vstetXmxlA4LmQkgt5MKYyewBaMmrCJB6OK4gRwABna8qnSl/
gPHCYAAX7Xd1ozda56y9nADT6fTW0AcZduvZcj7cJ3DWkW73XFv3o3LD0B4PN+rsaqjT5xWGiDun
Qrh/65a598gELh4AiXGuGVSvqy8nWJ6B7btolVvJ5KmGRNhftE1fPZAZbH4k6+RF4+N0B1qzfQnD
nFI+/SfObkNeoRYcbJUXaEJlTQJKZ8KK2AUSus3AnSRuj0xZUB/lV9EJPS47KI+4YKz8tSlNw38w
J9viDGNqK9rT6cpwFA8GE0DoNKA9xWQcasAqzVkon9wR5WuRBy3lSwCNd/GDoe1EPG9cyJHt9P+y
7jopvWrD9L46ZYLWLXpUx9IYPOgzqCtL+aChOQCedQwkzjAAmM7E1U6zjaj2Sygx+WpgWoQH+XRU
TzDbiychvDNh5HttYRElH+cv8gb2FDArXQQArhqXhLThhth81jbHKumrPrd9qGC2Df64y7pKsbG3
CsRgqPSejFVoXpQWf5uJR0BT3b65du1SG+OVX5lsbW1eFKrwY+7ZdjpQENYEEcY2pFHH7WJUyc45
m4A8fOgT+hqKFaF8c/jMM8iZBLHM+9+DbFw0+JFMEdRlX/ecrF3Mnj31HTWAFUjckr8lRPhE9A5A
dbi7gi2mjGTtBK8hmPRARUqnwGzShqgCUT6jtttF5UJRZV7ahz0MGhNfbZLWNUyR0SM6FfCxkSP9
tOSE8Z06MvzX1LvTleiH3SfUyl5OZPmaENKawFYzLoCeISf0nea/4YrzRBlxeRdZUglkgCMruNnc
FeNDRafkaLidC55ZDqignW+hjD9NFPGTUrZWJk4F3WQkZ0e2D2qIAGSM1H7EFY2BRbmB/jBcdLX6
xB8GjIvk5lumEJI2Iz3d8yattcodDQL7nDVshdvb2RM3wAWYtOADn6bXKTTNvR8mKnykvszRns2q
mbNEXhGeU+3jB6jtXWveMSYv2T9Tc3SkgHzxxkP5ZxqzNL5VrXzlw6SMNl3051v3Y5k0uCNdLNkw
Hy8pckfF6UP+BKWibcpia7ANcn76ORDJdvBrsYf2b5hRr/Y+xmwFIMd+Ik2wKvCNnTL/oDRnAHY1
GZyD3jFMa4t3tK20ef+f0U/iZTYHSI+rBI7vIE2NcyvX5r5o9szVGHk8qtDfYsxQAdfFcFYztW1f
VkXTYQnEdXNbhzSNzAletTPd4qxMwHkaAJj14RE6bNCKYXizHcIPVy/8jmd82t+eXdFMA9bO5Wjw
e3Vml80VdlQyLZmHSfc+eS6NAMeDOFNYzTFW1VkIZWT9ACMTFI7bn7CWsP2eFKbgmaRU+w7nsrmS
0sRmEEC605rgk472fRdOJeg8694dc1g0gwSVQTmUKTVSl2Ypt6BpLRYd13ZwqDvfUnBdWFWTMAAm
Kv7/B/svyuUf3GMkCfPPZ/lXHTqNntbyjB8Qb90fWpbxFtwiWI2W8uIR9yZM22PdCOfihp6gR5iR
mkI+N2f4iD6Z1Cdoh1LASCv0IrlLE/8nhsxcoRhMft2fKgxRJyjwrJkBlmnKyDbdxzRcz5RMXVjG
sdIet6KJBx1+M+bBbCXSIdzF9lhB1BG9obHHT1SH+kgRyPS1nPjHNh/Zpbmidzc0nlT/+FdTZK1v
qpyb4YVIj80bxDDUpAXgjuJt3QlMUyj9nn6lhAlWhHDBB1Aiz8A6XsfggRDMfsu8EgG4OQAMclPj
rFZS45t99r0gMBxx3PN4tOC84nvmwkGjLxk1Lsgl7IviOS2NFTc3a3U9w1TGXMef8yYB0KpgShi3
dl4NnZWSJazKSaCnB3lhFfjQUTfMKo2k5Qu9yxPos0q4jfr2/Wq9En8XlrFDW5pbbqPtYSm0uBuL
cP8C/twfqET+xmFpMFNQMZhK7sbn58QKzwkpEVsOJr3X/Y+4L7S6dAXsKEQe+HmdOL96F2uBha3J
MNTdhM9ZE7zwg7rGseBMvcgR5sfz58yOv/+s9IqtT8ioi+KBN926T5JsRwmtyiY4SUKYAaEOvdDG
GjO2SMBKGKDJUd7/EUlYDrT3XK7+4kwtv5ztElOoLS3IXfBMToT7w1r5DUUJbxHydPlbxEK2fekb
uxXu6wYUzZBtnWz/yKzYKhgRlrImiB4JFGRpoc0rkXbEfNRpR81Dl9xRNLDqCiotrKKE594x8A4s
isRBaf+onlxjZi1eVattS+TrXo0cWpOOBr//Qh4Q6aOhPsjDhDhNLAlyUxx4c3i6sI/LZUgLhHnE
ozzQHlEIxOSHEC+wRCGw8JOnObLOW8/J26GrwS79H11XrX1Imy3pRJ9YJjWIxqQei02lcOOaWZsi
9zBOOB9Y5pl2AAs5sMvmjq4N4E4x+69YkTpQFhz8o/JXJACHCnupwafMu7GHWcDlxGl7jCF7DvBf
ZRUEc6mb8XDvvAlbnMloHH7GNcPZGfIHNZU3246F5OC1gF/2IdMzytfHVTTnDUZfn8ujn/qKW2d3
pDj8djMXtqYDNKzn2x9WFXg8dZLu0wEl7JaKv/45P17DJPzWGFlwivFni1AkxKgJV/l2w1wgy9BP
cdi3M132XpqS3BHrD6CIMSLW+TNRoSE39HmUGj9FxaiRR+GRUo0iEGVdd1OBcgKowsQJZ/ZV7oW3
735/Pfnc9pwxUt7JlZC0gaUgiUecssIivvqutBHESmFv5EPCUrF9jUzHvh/ABj7yv7TTi+zP3fRf
I31Mwf8Mtc6i8788EMGx+GLqqj2kWkwN+DUhU3YTr9dBjD1rcfocLsuRAYQNV0aLZlWVDq3GPZXQ
pU+4ojNhZ+1HN58NzuyBC3W8TrXkju/hGnd5XEYbv4LWCD6zX+B1DEvxIj01yCw2nCgTlNUzlyey
7uAs9Rg59BgK3XiU/2Zhs89SlTxJ4cy9TSrFuD/8IAexFmLHOqVo2/CzK3ONxkem+P3oSu87dVCB
TphO23eZ1rKGxi5FmXItxLnor5AU2Vxx7+f7/yOujPBMHR7lgsWbPgFxPWjTqqCs8foIQ8IKGepA
e/ISX7HNLGI62XiHY/Zs/LjXNcIBCERCPNpcojrMxXHDoBMR2TfPJgg3+uxuMUAoBn+KPqHpjSgv
hCTqNbKjDbcDJtFWwq60TMtAQyVA+TBaJAZSDSdK/5VfVgFMaowqJ8H2MIh8BgPsqWu3x3w3QBys
GxjS/kuE6rdvAcbjXGQ4f6p60+0fxOhjSX0O4IVgFgaQ6i6/IasWfpH3CyQbN2qvhzZEoUWxGKk2
GTDRRo/LdRoKDXTvbubUsgZ0Dq9KLDXZHRRe/ADreo1XFVYnkXKSp51kyP9AE9rFawkl/qywXsQK
dhkuavrWrr8vQr/tSIHBbL6haTNDl3D8tD0+LFfLD70BhBpgVN141jFhehfW0l7UGZSWuKJx0XZ6
JQqWS3lp5YDj9Yuc/bO64WvD5mykaRYKqg6l3zfzNXOnrLkcYt7cNnfVxyZbUGKZutPeAY48iu2u
14Pn5IFGnNrg4hF5aW0csUHNcYpWpRIS+vumBGbgSUsk0xjk9PUGcNQ4rhRdkpiSvF7+tbioLv94
4k0QW9eOjv8FFkKiSkyGepe65KPRBsPERuWjSEFcECpLi0ntg6N41psDLrKkN+mN+PR/yk3VfqYF
MMtTB57V+AfvNT7aHl4Ec1Q5XjcdqDsi3pdsCMOCWgtEeJ0TaSnP0n8Cr1iep+uZsGjxHGrwqpPW
0hw4BaePdYMZIy/pr9u3i757yGlcrKaQfLJbAJMTolKYtjxgIQv1/Q3LLFpWibcpScWCGFsfrXKE
aWDvJmQ6KVHl0V/p7FHCmKExR+JutvdvnrqS2N2ImGcQSJCLzlRZrsDKR2Zp0ILXjRmeJdEPpC1D
xdtijdG8xgLVDxjIcVQAOcQdouN5j8Zx/Oe/X5t6rUilj97hu98iekqweC2Lh1WCOKKMRchrriox
BSbQpfL9O2U4V+ERlUpt8OSVck+oeptNaNluDyyGL4oIENlo0FxlGnAAymvO8iMvC0cwMrCRkJiz
vRiiv50Uj5shniFPKhFetaJpLKqGFDP3EurP34XeAGr3vTUdq9aISZ0hYBnmEdnGdBHleJlCQr/9
XhA95Ql8WwEn5tkTwhU8ieluAgm9fganCxfb+Kly6Nr07EYVI2dHMojV+qd+9Ggbl41UtsT2nJ1Z
BQvPrZAzyEQYBvIICx5wwAqX1NQ/6G0D26Zaux5E0aoaxl8M0qJXsrg6SFF2GBF6wUzNbz4Bmttx
kTLAQ3RbuXT8tEhZh3TEo9unnpLhClS8ptRz49Sh5lP1EO5Ku3/FajujmqZzhAO5VmMRWC7qIlR5
6jiph6ZWFjblwkDvQOr8hTUHjgHWuh4r16oX3UO+5kWdZBdS1MToNk1SRlhh6e7LpcE/Eb24TjY2
ye98OOuQ3fQ7BQpi/Yo3MH21k4uW5t4cwLq+CU7+peldquJrbxAg6oKWAQ/sUctkLImy52iv7tl9
YLsYtXa3o/EWT93bcrOQ0YdW1X07oFPqRCBXbtWIBPSqEiiYwPscG58iQdZRcAGJ4QQislLEH+j5
/PBohWVaQQbgWD6QDChWwhYLJyjZZQEWPlsGO4VpGZOUUaGYr+g4YBnIjAQVKHTE0AKy08xgq7Sh
hEwuulE07hyuDYX0R/JUvf6a78CdPn1ONAl0eiOcT8qgKkKtryrBCua+NH6ohm5CFllGZHBwjruH
oP9mwRaDLgKoLdYvpVPaUovkyH+njHJUGBOLE9BjI7HdyD8t+4LDjUdoQQtN/2Opmn3jNcbt10PL
CyjD5nwmq9MsdQHZnC91cNKDkSMz9SnVWHZbHm24SoMxaD4TZ9V9SNtxsNqaWRRhNewNlHyuZv/Q
LrllU6GZHtCXOWEJs8fF0PxGuJI10Jbh5Ob0Q/65EBMheXgqrgINUsV1j6/Mpm1dJMoipt28uSSA
cBqbWi2Dm/cz+FtPXLc+oHqEv7HoSJRGeh45/7Wzg6TAWAD3Gj5BDvXweBbJ12jrd10Q99+A8RRc
ueBVy8HnwrQWZ7nd/JnWiPkGBnnNhRFfEEXZSMyehI5EbSNsnLe4FGcONbh8JzzjG0+W8xeLENZq
ybH6OMXnO4UynNmuRXNKyzMQlBHebibgjhV8jHwnJOCeV07nzdFHyb0WiuFP3j5N43v6URidG42x
t9SVlXT9Q1AAjByL/SPXuXtZga19U9YZZBTp49GMp8pUDcyg1L3uGpbAxSgfSU6n6mb7rYThxdAp
yXVDm2eSiJIglyyfktG8q3V9q8NjjkRrP+7+qMTGEjY28qBFBQWgwRniL86en5JDBXS+kI/p2fou
wMDbULD3TjrtxNmjUb1U18K7+rx05E3GPP4Fmob7XabpsWTxfqIfsWF+X+ne/ZCtI4kebob5wHYl
F8DknSQ3OrfjlYcvE8CfwAmCFyRfWYaAbhZI4GpfHCSpDL/DmxdbSB2m4eezjSq/Xi7fNmYRTmAm
H02+F3x8lwEcRBSnETbvyj0Xe0KV3Oy/KSzTOUboA3kzpN3A65iXB00EcGlTwPa0Ll/oKdzbUWKa
9lTFR7QFHIyI8g5s249ShLWrDtEWs+3Rp9lrFo/d8lFMCD0SxAmi2UhSqQIm0xiuCWnbvmTBRqot
k3T/tHdtOWAt2aSfPoif3Vc/aVeID0sDLdWUJLFuWpYzpXH/CLR3zmb6Q77ZDuR/+i9j953avp7n
K8fHp9rBzPCZsGbGo38SUqsJnyDjwjaQTF5HRGIGmH8RV4aldyXWxdyd32M5eQR0eqP3SRzmCE1f
DZOF25iCu1dmoIPl85/5PDvUQOBCA/puQ4czglc+75zwz7uKAVW5SyYSl/z8JRYPCXt9jr2KlMsN
d/JWALMZ1pcQKafLi3O10v43KeWNrM7CQrWVzY6bfr3IQKCtVMu3ZyasmczhWtfGJl6w5QXvvs2i
OSBfXzl9UzvaamOvEkHZgRPLKDWPoBvUYbI9PrTdE58mdwyM5eOu+U6cdMsVvfcpTQJUcApt0BwH
8FzDlKZhvnFUg7fGMK4cwNGIUDyaQN7iLUUisONg3mRTOlkJw/eorqDJA2AecAplQ9uXOHM/ZiBR
UXsw2AJKXnheqisBgRg/+sUq5pmRXnABjbm+TSA3uf3owUNrtkm3bbrsgx0Vnpmb+R4/qN0wOeg+
UII1h0YraFw+zZNtb0poyKqI8+LD+F8Bw3qvia0zwiRZAyTF0kr8zjUe/Nmd7YqQ43ejpK9tQVWJ
5xyLhVurItpjUZ+bLGqdawghQb5R5UyShOEU6IdIsvzfjDVAyHftXd6TEdrNt92UexA6MWjs9j6v
2EZFje3X4/TrknYuineTP1QQZpKHXMtFBLHD31x1EKnNtC7Yvso8UugMPGEPbP77YQb1ELyWD549
5E4PUnT7Q4XjZMzrtGYIvDfbP1m07P253et/Vt0jxN77zhZJcmqduTTJtM2yESSHn0Qj8vnonMws
PcrWylgd2gG8brA1G2KSgQHjvnO9dFOhWDXkyi+rTQSPpbJzI0FZJu2RpKnCc/euhfNSgfcatKdy
ljzYXOaAwDXcl6stE/8RwG6tf3B0CakQ8dBwuBD/xqUI5sdQzcv7Uj8EIjqK9skprcINLbb2ykmj
O3ZH02vrgAOwvyyjSdNe+plt+XJ+mM4cA4vx8yxrty8hQf8uKqXO6tX+b+RxxpQprlvW3ywh+l6L
tYJEdWHZqOqCoV3C1TojxDkn5kdQs+oLpkyM/5HXFf6ReaGwVfX/GDgPeIurHLQKBUFTl+3t6ZFC
oOolkMwxuJZeljd7klhEbLHuXvYNEIMD37fNPtMZJ1sGAXs54ilHoGW1H4ELk4FGMZ0haf2f+ZFQ
SQfYWOeNmH+iTqC0H3on3gxF9evQY07h7LXfxWvnrOeT3FFy4vQaf8tpCKmNThSmyaU/z4K/2VAM
mj/5BxxbfO+lh8r474lREvp60ERYSGaIpeSqVk+4RptRb2OrEbDqFvi03UVGPD6UWaUEr461UBYk
qcJhXWoB8rQKX474onNi2fWCVrAqRcEEyVqtmORf2SpaFXH5fklduFX1U2x0L8GAU+m8D8WOgNI2
sl5xUPsdkAja9An+IZ5Wj/tWPSUZGoG9To8htvj9TKLckw9nRo/LQoH54LmBDAWJm9GqIE9hYFcO
7vY6FPsmD8w4/8nWm3xLQDrZxhK963eJqJObJJKYaJ5O/x4n4i0BlVummwpZpBXFMzp+G6HWFgHy
XIckpBTlXYuYPyZAB52b/8T3RiVAD3c6TcogbfMsOQj/MRN8Tij2kdnBF+B9l5NYvGXhze3BnSkV
R3yfeFp6r5JhKifVFH5Jg8w7Sym58XJaoHvTqLPxrrXgMx9j8U7d6mwCclUOWnIFR8Uw9Zwoj5v+
a5KbgaoF8Xz7AIQMi41QEFifyaz6izXO3pCSHXn5iEBL3qYukmGKLxI9TLfPbbszJo9wxWSUdBao
g78pmfnruVlkjMq8yWaLaStadJSTZ3Y3RavjQz7aZtR+zskuj9kiPd9AJ6X1iYgGR/LDkl/l+Kqg
KiM2blqcfoaEz+UIaKSU84arg94GBrT/O+W+H4rW0J+v6mM/v340DoLhEQdf4IAadu/YwXN04Zuu
JzH3h4lWSHp7Qg8o+T6cproxR9DNMRsZRl8IL1qt6XK/khdj7hnYBdK7vg5Xcy038zW9HJUlQA60
YNHuwvuHyUz58r17JikYsPVpAEj1pNhzFUkK+WvboYXk9oAGmyslZu+umrkrRwh11G3CUxEV6HZf
gVEAyQlFOqKHMEZjkqZvNMs9wWt3Evce2hp1v7frYglrzljdSsN7mxm4MOk6/Xsz15YQ0GX7q5w8
FF9ytRDkWyojJP/+6u8aXWAtJS9cGsUJV1qaxBZ9v8LWf48ZcBU54oTiNrxxwLkGxxhS0bJlQ6HO
0fhMocBP/l4PvpT7DY54lJrRnIf0Em6TWTrqaiFvxU7naSpVsHdpl8tG6VbNwh/U5t4LNGtn2+Rn
uDrVpV7LbTe/mwL+rMq/Obn8O9LzQ3PdOIU8Zi1JpbIktAWhJYOnFTBNlrHxGrC9PTTnzFCKDyNp
gKmzFj4nd9LVKbX2QMpVX66SfIq65GWl36IpKkNboV49VDZu9qtR5wZI3ZiSk+7cr4q7pEr+Gkc8
1SHY/4rp65KbrDoyigyOKyNy2rcePfVORjytcQ9rhrgJVwhJhI1TZNACwH26SoqorqMv7M0nUEis
Hr0COTeY41KPqFshJDazm8CUMRgyt+0aEkmqDnWZc9Qm9p0JP/3vLfW6Ch55nFIUvCnNIqZcHZp6
fmrngWddFk179USA2dCLvBpdJBB90bP1IEX7eHR0q34CrSK4/rkMktB3VBXVCXr9UdYKWPq5T2Gb
w1I/JvxQwYCdr33hJON7JHQmFdIKWRX+AXxewxDwujSrp8QSsOsIlQZ0lV6ZF3MUmcvM6nur8aCm
Katnjz6oyd5RptSZz/WKIG79p9TMWnfCj6FidatS6gDvy/+Umyy9mOYatlPLGjcxRNUbwEDpvpVr
14LL5FsNiuyWrOaMkuAoP23CrqaOEtPpav2HU3l1pSBZniAdcJeJGt/2sjYvFmt9wV1Xb9yIwz4n
sEb4N9qW07Qqj5QeeOiygtBYnYASv3tXCdKGJTYEgjZcUQEVqpzdxz/elj4aBcxriwVFUY6XBNRA
2iZdMSjlGAzwbHGom16GwrCgEnwiDRdSvY2w0VfDLGQYE1wd4UBLmNcVx0l01/AX939w4lfRaoeZ
/mXqEV++B5mTzFtwgKbp7k9fApliKAClhwKEtUPHkhLoLXMz0Fto36aJ30/cwe9DndDEhd5COfTk
aVbG1UlQ4cPiob406Wfr+YDDv9US9IPG6/hB37/qH6DSLTsq38/buNPPDC4Uibopmr5YA4SzWzSD
VpFoipPHPySoTiUAIyI665yUoBqXxkOSGZtbZGhUSSVH4+oLpf2V+kkIqxE7cMc0uf0KAqUxdo2n
Egk0YUFS2Uf4JbfeKOYZTBb8QMLWmnM1WSdDzutbQyg7pk+5oUDFLI7uHLtCSL/j1ssNJ3ihZmrC
adHJCfeUh916pwgtzJlrZQYMyulJx3S+vU6QsaFZ/dvVb8BhQV/dSL3AGAM885WgFI3W7EXSK7Bm
scal8KFXNEwVR/526NLMXilFkHt6yeNwYRYDjCFPYL9jyJU/loLqZSgsu6XApMkEbjb0WEoqzABz
jzXSEguVv2Bqad7PO7wP3EfcetgW85cyXrt4jtxFf0V3zTlS41ste+a6Mc/Dw3vSEf7SZoKJ4DIi
I0dSPaOO2hkheYxuKtrPH4v7tVHk55BBeexlj3NdcZgVk1cSTn/sMDge4rgEI/SGTrckk28GDrZr
PAkPLbZRkDWMnB+ohNfWjg84mjII38+4Ma/UiP2IGvDmMFKz9zTUggWy86EpZwQUSzOohH8m1KKP
kWI/Z6rbVyYGRwTFgQju99dEuUeH92tU9ezvYMPXhrcTnetqaHlpa/2gWggk6jC8mCBSdvwdmjix
qLmm+WTwHFE+zjXIzhL2q/Snl1OPZAlWmYFpGmpmxTDum0XoxBXHG8qYUHOOMOukH4Rz0WJngnUF
ch6Wpct+yURb5gBVqZfJWgKcTxIHdpdfeJvb1k7h9Al+EcvbOMEQtKwrKJvlpOAtVXfzFPhD2+eU
pTficOtAw3Fdu9I87Lta0Y4K32S6weZZbeBI3p+G2EdTyj3YDJaUB6HshBB5cHDi5+6pCl9CWJeL
vcjQobiW/bQuld/GMJFBt2w0sdyj7r5xO8u/UyRYrWXd7eecNmR/alX6e+cFREMyxFt7fTYEPG+3
tn04aq49ik6aFfjCHOY0BRfKCY7hq3VUaW82E77qzyBUvVn/cqu25GzL0Au3McCPTiTEgQapjJW9
mTLUZCU4cWmJAg8e1KcaoZ7J4Sl5xL+McA9JWSHQj+N2dP/mgjQzRcPFrmNUJSsv+KZrkl1Fy6fC
ovxztJBVIVT7fGzKNytWlS38cZTDXLB52WTe9C4xYvMMlvyVDqhgJ2QUNkw3ZPyZ7MNufv8rP0X9
7/ZdxM1q3sx1HSdmnmJDNpmlTf3o7KHoz56tkt6bXPjYaLgpsrNNCdkO4ALtQgCE9iUc/62s6v4c
e4mm3xWP5Qgab7hUnkprNeoUkBV6BT6HiPhrlZgKJvxAbEGAZWmiHNAoOlwuaINhl2sWLLGGaPHy
bxJuMrVpP9LLLQTO1frWj7JVzk45pP8hOhvyeQvEAKK+61WWOVj/onQDf8Z+rJyqZL7RK1igNpjg
l5R5yHoaVy5P4qaRdz2wMDBhLTUfwUU4lR49k+n8g8GukqtKkMiczZJ5aZz0B6PQs7OlI7XJCGqp
NynfKOYd6hi0jLJ7/MBfdw617ZoJXUSRCa8c2w1lAsFFUfSGaGrhCBrsBYY3xzp7H77vIL7LkhtZ
cPWWRHjwLgBw5Z1nfSPT/nr5ttbXd2ChhMG85g5YCSXM9FoRVZs5q8+dnVg3OIEqxdXKl/hXWrgc
5K8u40DompbsMaMTLWJWRDLIHzeUToi1fn0HOEZleNR27TtdUdGGTrYriXcbyqG2QPsOLFkgprwG
fmGPhn/i/GIYmeDpKqmA2QCbt9gWI06CzJPhfZRiUTfw0eXq59YRVcq/rKwlQU8H89eJYv/Fvst7
iUphbXaJeKrbYWx/fhRULHNJsWraabluJY6o15TITtOQ1avSZ5OrGo8OO4rUfjnBhJANb6SitjLE
0Jvusm2B0eoQ0CKk7MZdNIDeBSNac4arIqoralJxXs/MSR9T/vReyZu1dfGONtniZhoTFyrg7wp2
8RrJizQnCjhGGNN/Vz85YljsPc0YrQ2TSDtUGI9qxoXhXOGIY5ej8fw4mIMrIZPZS2ul8tEj7TDV
x/KATblwkqXqBIqS74iJgB6EH+D9E15aYM+PvDh3x+F8kotnNIzwNxrqbsCBXtwZadnwc0uC5w2O
1B7lnPA9VeJxpEWYf5e8EmmAYVfUXhWo9WCgl4ORnbhnKws2p5dYGn8iaP3hzGWn3FmU9FeQPAJp
1E1aRmbfjwZPH6AicIkBBPZ7WspGG7X2/iMyJep3tuVoi1HzT+LWnSKLftNkVY/L965lDTSr8xf3
5fOoSsbSm1Akt+MXRExDYvcce+fH133msJEQ0ADiz99YIkYBPHofoqEJtN0nttP1xd3DKXIgA4/x
cuswdQsxvs38B6oXCXRMH/OzIUHscjW5K4Pfb6JWZmtxGwCABw1jq/KrzrKan3MwQuTVelacve8Q
e8ajCOwRT42o4nQcaCQimcMrBHAdhcnyw+WDa2xNn8UHjEO4FX1NLyOcm7Te1Ms4YBHY3WoXXiV/
pX71Ffg3Zp6SB1AMxl63M7ee8yqyAswt4ucwj6G4YnRb0Vs10fjw9JY0gbfol2+XLT2C8ZjET7t2
myMGfcCdzgQkWhShv2lWE7sAMLSbMRIyswnP2uYFatkceue6D/NgPd97CTVWLj38SV/oxuBppwow
xSBNDDdCKI1XXYj3Ud5qsg74PFhiInTAn8diUodQW1WXIC4WfqB73edpkLktjxGCFOeyuhDOq2+C
m9lJPj4mNOQCRCJQcJ8ihtLwFWLyiXfG/QeALLxq4f26TBl81mqGPJDYIXgOGQ5x2AtkD5k27moi
+Tj3D8SFJZKdFaepmxcgo9HIVMLUz5KZ39znDv/myfbLiQhwd4lb41HLKyDbPOZNvco5pDB7fL7D
1vIFAsRrt3jfS9PMFUrx1qfbq2UkXgSfxYDB+PY7p0A5GYXM4caBmuAFNpZfgY78lL5Hf4DxvEK+
p0ExHkB5ecqWd736rbgO0EJyIfAci8kzWMjkvXoOUqlR33BSlDGn0xOmsiAsisefG/6oDMxPB2ha
P8lGLQRIZZhvHHvUJU03sBnaQzA6KSB/R5Ky8tBWpO730Uzh1eTOTie2p4449iVTFEoRZataccL9
p9eEcDd86t6FYDs1DSZn7NKKQPBZCj2HvccLAD10pC04NAjXv5XbxzZ8Z22G1jDXRF+74FjSQORz
gyRIXKfc2fqRtk4fUW/zzilgSqRS2mM5TPEO7MKGmiFFJMdFTrhoEg8Fa9U/Zfo20T95xqmjNYtO
HkHrsgCNS27ZjEVkPIU3OclMvYj2ARHvI1tU7z2NTr6WOTWTEMSs99+CIQy60q7LaVXl6AMdoh1S
uVBxN/xt/IaXzkTiA3sOM63PlCmxSSx25ySQY9flTPcy9d4Xq/+XQxdRxb9d5ZAiU1BYWXUN+I+h
GH1vTasYymwANIU+Cwm4GG9wuqCQwQZPKl+ju9/Zxl3pVQeBErF2Hn+HXfivOHdfjeY7ELnjkhzb
MXLTgHBqUEqKktTXQoGU7ATVRP0xMDoaunDV9YpvxvVhR/ZU+N6QkN6kYmPQmcr8cQbxbufvT3R+
p1XVDDDA8/5Zep+xBhGEHmO5rxvMNbixBOSdupGZmeIsfJkYvEw2TAeCtMRL6B5K0KYYD0rTrs8K
x0ktx6kKaPajwoSxZEM+jucZIrOeSv7ORkVkhMZ8lSi9PhL+tHV0rG/tAzmhHVTVaaDd0PQhiFB8
q22DWCZL+uGoUvqiSVTOaq9IHtzTF/KML59nZMd/sF710NkDi6g/Vuu7AmPLvV+eLywtmD9Skr++
a884YiA22VoPZMgCuIiTL41V0trjhpnIzl9NumfguthH/tJSCQEM3F0jbJSLG9XWHe1yjdR0rj0T
3NEr+NXsY1FikVZokTnAhjg1TxPyiUDLF//UNgWwC0TOKe3fT0V3scjXzJnAP1w8PrjO7ZE5YWem
lPh6mxT3jj9JcemLrkYAhlUXyAnSZ6ADGDwoVKP4tfV7qQ12+FmS1ooRxefjPGZ8W21slhoJDkTY
2OWGMTMoc7cz/90zPeNDOEtHq07rK2yLuiH6uOaDgAOMdTq0pOiRYqn1QNkGiHQpvHBkDWWe3+vG
jDCaSL/yOBq5t4MaCN7YmEnom3Z5mNk/bdHiyfHkXALSLKKzJvjDsCUD/ADvRouy+IlPsYEsdlsy
TfU1sL9alHplPoRc9yqppjQJ3akjGcPB7aXj0NnSTbVmRx+/eXecEX9P2mJvqoDls5Ldrx3dZ9q2
iPKAzZvPPvUMpWrSt1kjXJeZ8rn0nW2HVyFFeiB8K2VP3F0IUTcRE2YpxfYL0CgHzhGIRT0QHWxC
N7SyxsLtI/5NGLE4cKTCwjdnoNLhb74TNhXzjalJ0TYjmFdvs6Ro/wwJSi5m2kQC8iuaYqo8mu7E
PavT4dhEFWG5jQnSvvwfpSWjhbhk53HLxpr8mrWzxZyD05uI8wBOdiHChGTPVtPkMA8aRPrHwK8V
g3ez9Fdt2STh4bA5NaDcEqmOsr6xwPox3L4rDch4HbRW017KHblOjTtX0l0aKGgwyx2fv8IBtXQj
hJdwWhQaB/eJa06OsoDvVPTtFKjoFgE70AqZJeU1aDhcIsFFcmXoUkORG2yJwzm5dyZ6Edr0qLfC
KX36OkBoKWFSxDzO01O7KKmEyvTP6AyGDgN4yC3TvZkTYtyGbvj+HWiHAlcqlfmZi+5DgR1m4UaN
WlAAzVVCKnJs/bqw/8ihzDKDaT5cBBaJDplzjdcb96fnLzAiIlM2Yj39Q/k/F7oCt7sfL94bNYkQ
F5MyOJjxIhXWeIm4Vt1RF4THP1cZa04lZ3x1mWwKyZ7GaFqj60IPCa2ve1FqgT0vl0RKgcfOkzQA
mRTtrrxbLobl+KzG1BU/6vrpKOu3TLe8bgrUXXxv8vauWkRbsiXAPX55gBMg0x3+M1YSl3o4OL15
VUc78eKiaPPgFyRD6bKxjhqIHPkyMmH1vNGb10BMsJEMMLQFr6p+tCm+vNHuYPhuzWe73ol0vePk
e7IE90FzBOLeJ/PH03WWzGTeSqY6ZWjFsdWj2A7324TKq42C+J/fmKfw1ML0YYppbST+xHkFJWg+
nOzaCpRUpdG7iquT9RtCiZIDoYenImKmbTQlO2pSB2+SCKIAKHlUWDjiI7v/11O/BN7SOpYbute+
pT8xD871iKWkfVPkTcqvS+OuNKauu9F5KIKqGjGCGUcvVOSoQldK0GjbF1zjsFJw6Q5YfntGrUNJ
7yxtYNSlp0B4u8O8I1dOZe7eUDopphwUV55FA6u1Yt41nOPN9xosoH+MhG0mJxrcUWtEiw74GO3A
j7RVEqDkTzxIixdkj18wWSYftKhJMEvFncIxPmwkCjWLhZqDmDry4mArSPwY0KgodFpDR1ps+4v9
HfQM3i52Aj5kwuN4FxjUgSwjg8mkA99ypZAB4kba7rVxLvZ3P4XCOkCPdlwhWzzcgdkX/OZvH+QD
AxL7ulAF9oNNC5+BgM3AwuALZB4OiktPpJrg9R97gKJKTW2dwHug4x7O9uBayMR7oztCmiBpKs+M
8t+ek3F+mS+vKjbLxEAIeSFVt/Ti/hPYcBo+Azr0YZ3pdspwi1W0GcE+JPawD0X5seZDw0yHGe3c
F0SSM5lYRaq6/agcHNIdK1tkjkQJ56qn2pKUv3iuSnycxzRcDUr6bRIBZEC4ZtyDpnLYt58n8yf9
oEY8OLIYpop5+c4zh9kOK3gy+ULCf/xIR0Od+e+Rc1cSIIVO6qiJscPNCmTbrqaeK60gESrtU/W6
J9D0yp00gqee2lziOPMN5Rfxt1uWRh/Jro7wcgRvsplaEwAAuP+2X/yuDGm/fCgeE0kITq/O0H4m
lVkRZ3GugqHPdWMWCqTmmLUHAW8jG9BRrNGvpT02BAsNY35V/ieduSKJiFQyu5XSILijpH6e4i7e
PNh++J5o349uBqrVgD8ajW0/Rnq8YWMwWFqdD22f9hXSoM7evJGaMQ3HD1TJaSNUzxmCTQiex7E7
DlpXxzhYdNh5anS3QODGUlci/sW3+P7s/9ninwKpTLn1KuvBCH5zY5krYGEuM//wFbIiEEJXYmzT
3UznCJo104Pa+xum33z6pZ1afglwyU8ebYIsa31ixOcLHRnTXRnrvIdHJVjaiS7w584E97bb+f3s
mRt9Gfgr0KouS9i2WkIBNO4PjZdjqYVbZL+26wcPRBsIH51QVaGWOSMgvQUHI0nwYLHZSxCGjegd
DCnMS3il/26FG+FRChskU7ptbPUq4CSoN3mVwTHXpmtPOatPYhWlc43eNCFJjTR6j4fqhyFLt527
XVXFrDN63/7DYYqljvDagoqUZ1cflcI4R9Nrb08OGnAOX1f/KbmVgpMO3V8GHIzJ+wqHWGf9yMSt
8LwacaPQ0G+5H3RaBre2tVJi9yvkxUoai+SOuX3pMOFphETjc8SdStoPFt//3jIsD7/9KV3204Kv
wDltIZeN4+BBD/WNrYAStFc4GbHPzOzcbevFX3Z2vd9lHAlvYsCaaS/rDSwdLLIiNCqeSzEDacky
RJZYhzmrGadbpmWTqkmTrzZ4Wb+zXwOdGbcygFojW1Mh7TtbRYwEtZIRnZwyEqfmOadwvc6aHJTB
JYJ97jY3U0ULOIOIyUwtCUIL6L8Myx1dAc4seSOx2BclJA8OWZYsNjEwADotePwY1SZC0I9Tsh5u
WwsRXoDyTz/mjnN6EAVMjBGfLlQoVvsVQN1Xt8t/l994khIAdlBV86hSEj/8kKhmSAcr4iLaWwUy
GAfzc+cvEWCUpxA1CjDJT4DJvsOh4xxAG+lSrxERroIi/QacoVwYTxkKBxgSIgAdCrEDn8SbTG57
AJC5aaVSqh/ZLfjpvIw912pJvWBzOrOkOg0halIEMH4L00Xjhk6Or4H481xob6l3bwU0ej6TRGLd
vZHXmsiQCHR+hNPQOnpfrWPmq8jw7lFcKshAtVDHyYBObXl5vc2ECRQL2ImHadsDhJd5Py2FksVu
PinU4DqB6EENzgoMDoh8DWn+RY1NjWPxzRgyp5mEZ+1U8QYCzYtteVLTz8/1erwBsehDgkQrC1qy
WJYW7Z4blHyAJKQNBk8MVSfPwv0a15uuq65ETuQorIOwIsQCrx/hGi+riwXzIHvudaqNbUJlA1Qn
6Whj1v86rRZLfRpRK6i9HenDGOMICOj549S5nY7WM7d05SvCABTuvnWAToO1IM5hbJQVzIEtyBY0
vbg/jyP1UuCjv/51mJT6Ipovqj1ZIKzI9NBf/qR5sAR4j7BZ9pP9V442VIswMXhbzpWRm87DgTjh
omr+1VpFLq9xv7SCoTXVfBjlb49U8Hx8XPoaFVM+1gfwJb/8WMS0fvh5TzyuzAMrzaoMDTsAaIaA
5mu8B6weL0NbfAgXDHchWUMBntZ1MkSk8KVGMke1n7URd2/r4k+YYVT1fW+UWqvDdNVXXFoQjFzU
mH8P32DK0QoJn8vnaqZwLDiEVixDE3kalRhDevV4mnG4xIBW+UWMpgNuDZue+BCDTOmC8bFoJVNq
r1Y5QGCkz8LGYPuve3+88zf54yxzjggkCbyrttKjkFgohX1hIEmbVKOeVOJx33qqgeNTXbrvquHD
et2xDO2+ZXj6Axzl7w32vPX28ZiYX+caPfthxo+gmwkoiLzje0Ngez3wMfELVLb6IxpmkCwwczhu
sDBhVoODJ3g8I4tGzTky0OpBbAfmBMT5zAU3UssWW5LIghLeiwBh3Fn8q78WeJ98D53b+bZLnE2h
s+kiMZQADOaEk46nG3RQH8bePQJEJI02OuqWpxP0Nmce8hAj6iGKhzFvE05EhN00ofT+W8dRMRj0
NC7nzKLLLDBe0V9ByUbRiCEsYP2n6KhkIDefP/Qf23DkK3XK1/3jSDIdbDp7XmBjfDQ0Q/MgliDL
weSgzmsdjd81SpyxtioiA6Fwlyxgsxjr9ye0l9yt3Xdht3W+rbB54LgoPjV4SeAQgWl3vYhbyVlG
S36ycgJA8nvB1iVa3QUrv42p5G8KxggRpMstyL9KtFoQoe4JusUOEvq+9xmsJfr9TujNAV8Ih4qA
dgPLq7smJDKbkvPCXCr5J/wIKpS37PJtlc9vMo0gZQ+Y+uO/pEVUAB4xOYO17ub7/5lNiFTU8+7Q
tI0QHa0JBLuJSFrtO3FqcRqxPBLvhlMD6GYg2SyDLA+51SFJflCi9W4EHTSlsfVtNkYNWDpoCDOU
l+saCdl+zVYu71TFSzLaDgXEwVREjHW8hqKrnqF4LVcYBk79ehEIPLcu54f01IiKddyWGfOiRcFI
2cvk33NKQ1AnQKJI1CRnU5OT3Qx7oAjPh3hiFUjUu1kCn6v0wNKUAcYY7+LMmGkFMxWXmzMPIoSX
MjZL9OsYhAKsOjXnaRFfNA63TLoYgI9PognYSTbaWOq8U0NRlSlM1KYUVFtRIeVxkmMaqUPVWGs/
89w2D+A7RWySzzwYxp44X/CnKqtJCJpFrEHtMtZ0zLJ/e/tjLI0R9rfZXEWFNV2hdhbxzWtqHbQ4
8gIkLVs61BDeG78e2oxMXPErCR3RZH51wUWqvEf7XnwC5LgIWfaGUCJAGKyo1qbG8fuZq6fJ9QUy
EiUJatO+GR4JEa8+UtShL0bdF9RfvhdfIppxEzq1708HwA99k3JBNvSdbxNFpOTaaV1BU6zrm176
c4rObtx574+Bz46eY0Vwrjh7NTmMEtXoqkDSACDDuhP1/93TmuwYv+3+q+7SogPllN4bygDN9NYL
DjnVM7bmO7BOeqNA797F7YkPhXdqH68vCfQ3sDc7c7ZyLttN37spx4EbtQ8JCHUa14lwEbejeQyI
zis1A4D/zLHmTwLVWOJ2k92la4BqmnKjYQEYyj8/oIGye9RWwcGdpW7Q4LxcR09cIz1VKgda2TEQ
9btDWCQkqwh6r2OXhmzSOJo/A/lEQtqN+5t5MD48rEKYjbEWFcIlTZyHeNH1tsvBWVCPANGiRtTp
VQkQbTqPvBnaDZEHLRj9Mt/93hLg7T/by4BHqAL/ie4ZOpWj3DKYFrkKO0nsimpaGjt1LUj6JcvO
QVB2t9mr7C0w2LypvETC68XJ+DHVcUgNOiJQbR3rd3p9wPI81FGfSW5XOUTytro4AkGlFpZMcXTo
zDuSRgKylT8REUJYc6VEHTvEsGNmehRbEOlJFjNYyYlCHemp9boRkgl7OXtADl1uHRe1LDONTpOT
3i1DhN5C/CInAAK1Il9wicFlgyML5b8X7AqsCN8nepD0bW9h6NQdfPcDu0xB5+UDlKs03PD14QhG
K5i5xDnLw+Nsn0wdKIBFDZkxZnfHW46tWo70MVkrdb4CIBrwB96doPvXM8cf1uYvoT1OFzmZfGO0
wX/su5nKU1yBIZ+vnRmbl6hpbK9agNe7qQ5RwSJ1qZ5MH2lrWB65eZq7dyxzO2GRUdkJHT8Jtkqd
XnF9TNBFHoH2Yu0j99fBV1ORGr9YS4VGOOmLfA4eogCCThF52C0Sk9TwDNKlHXOa5x3Y40K4fy7v
BYxJ/fTOKxv25/byddS3zIIO48S8nxZP27hYbXT4tEIYieHNqtYaiuHzMXc5UakzMjrjUNFfoV/R
5o+n6ml7Id0d0hlzN41+ZOYr+BzMWSP8pnd6VeQNZdLcprkusvCCnuMzRyEsIkPV+Vd4+qGa2aB+
L3pVrUZ66IL/fowRc6hzq7ghoWrifbVJaFFrHnAqCsUSU4OmWDJZMuZu8RSPvvt8suBORbrxe6Lr
JgjC0nwQQyOKCl20ooGTDiRGKNIqBevUeR67aAx+wLsmWTah5AbUdMR66rwxLJlzjt/ywkY8z7pj
R8H8mBHzOCmiVqT7Vo5q61oMwtXlB/EJ35ugc2xIH05/DMajYZ31a2O45MYHwaWZKwNWvdI7roIb
LJ6eCUcsGxopu+yKDKHzDEMdJHkaPnFGfP8wr2oKD3rkNbgiVQgF8zeF1zRT0SB4DrP08fUh/1eT
F4PCZt2jEJQLwa6vpt+2O0wjwbTTYA6ee72bZNg4vFTXTUfxZwWzmG+yXIbtcFYYWn8EUqItKFSn
thcMbGjxbwRg8W4IXsupWUEPEov6oG9CIt7/jngssyVijgGAzfkpvyxG7aMB2XzPtbbt/wvd+PpA
fKlXs2xvETZKBfVbR8X0ZROfnlPRamzPGj1Bl3DDaVq/bpGzT6tC8F5WFfMW86dee2zs9zT2uTC1
NWXeCFHZ5zOcXlUtqUz9zIwK9eOiYrPJnIxQK97vVL3KL+x9aVI5BPSbHpwQSVnDK0BSKK/I3A2o
GdAe6j23joN0lPhF+N37K6DGuyrsjWhLSoCIMWmS1Yf2X8KWNsb3W6q+E+k3euyd72ytKIO4RV5u
KqVSuPsTqRgwlCjpY6laFk5W7i8LKHtIiOXEkgSPwnoEPuYQ/QMbCl25lob1qRoCSDs4mVLGObUU
J3XSqPWjyLSULhCfKcSQjGr+eF34+t9FLK2tfg5Lcap2puV9OxTpXCBuHWHppEC/PcjP15SCrKEk
ekZFshFMcFy2Pw1uuTPscakLK2OzHRF6GQYO7nD068JKeuJv0rmhGZSV0KoHxR4jLI4K2g1Hp+c0
6Q3Zp3HnZz56XX4JNLhx6cZH/41TJG04KyvLrZzAES05slMIDlUJjIqTDzYRfPWc7HL0TMK+x0C1
3YoSRxJqsHrUKP6/HDYSpoWa2itzUfPvRr389nKdIkUDhwGcygZ13dH+r0NqMWE2Fv85cxNSLG6T
A6fIHWoUQPPyY4gjs6Z6XiOx6EgjwrTW8GN3IxmNBpc09ckn8GrrFg/UjV4prp7yfWDxLag/lCId
z0GNVgbbl/Y3sddLQTzyisSnlst3DC/4ZPYwGv2vqlURnw8jKgnmAZ2LG6Nodv0ZNzVL7x33Hz6/
QXfzVydFZJZpnka2TVXhyDu7QBXdQoW9Lgh392tNN/g1oPd0IT/UJwGFpiZBOOWXnXTCy7hn+opa
AI585XgPwp2eK+kGhuiYy9QAc6TefUg6tFF8lvHG0KhZWptoUoHuexvr+Gfcm8rA48B6pTebaEjW
b7Nt+wqTLi/1ziIRfj3KzOP3F3RpGLOAy3QepowmoJbTmQw3Z0D9joukiIM1OPVhEAjVpSCb+9Wd
Bapv1HSy69fK09a+yNLwsSnyETnep3I64JE+4HcFn5Z7G+M+7/Sio1MF6EIsN4XnF3gZIIqm8t/d
s9Y1jF3KibcTsldmS89ANc28OLvEdt3SXFqru2PlPvzEE+IphfzOSHp1zODdfXfHpdNamhPj073J
JULIZUT03zTuIdFvfZm4iqid/mqsvAMKFsTDdBeGaFGQETt7PT8QiaXggqWY7IGapU4bD5OR5gfM
2frY42fTaYX+Rho1aF6bRKFMuRV5aAsbyffZMtAD4pgc77jdvxSIBxlY1HdPlferTUGrcq8cooz8
SLpfvZK4HzYVGocuKbNPY6IyLRYoig5LGzxMOOZDESIDEyR5hWniRrKB+D9EeQs18arW/GLjQFIt
V6ysonsKN+mHoQw6ZL/jcZZ6+0ndZbzrUG9EkKhpjUZ7jsQuNEsaY3oKfCQZHJ3VuZf24iZjcfIB
+7FWcVZ5aB3o0mM2jhEDUU26GRqTVz9m8sihC6KvCBiEiWId8aia1gxVByaRv4qxTN3rP4Ren8Oc
9iRy8p1D89YHoRjzrClSLhHI4wbL/2oC2vf18CYMMkdDFovp34KdhAEQzpQKtwQxAoKvQt/EDe+i
iDYJQc3yfs6Wy2M6fcY4p6Raf4NGwaVyhDY/eO1XK6C4udWVFqEbO7U3VuHANl6ln5WNKEGCP/R4
HmVYD2BTas4WP2qziJFEQLGW3qdRFDVyXVhk0xJ24oCqQ5B4mRdcqTgAtA5w0lDWuoyjjty42it9
V/b9q05jwNCTWc4EHYGtlUrkeQZpr/k4nK85iVpRJoWTW07WgT+dFi+5KiC/ZUXVHOP4PXGOXlXN
2krLIn1LpVTzOPr6sRUDSdwql0Cn9Rwu2LgNtOueKWIrAMjsg4XkQpyso6LDek324/gClc4fe8w5
yghGiP8vqwLJv4ZzfnVoKpdF3DkqE9xLMVElFUJc2b4WcaVoOQyJZthunbFaJMbx1Ppy71PG3Eph
xA78v5YNODD6l5HoLoxb2i59clnVs1ANVZf1N46hpsK97oh7KWQeEOeRUbZmMJW0CYVQ9ISnu/8W
wPv3dTPekNsAZ0mDxNoct1dLr7RxZyR56BXM8EGSH9PAalfQmdUUUupcTCha3vDnUwnTJjEGuHr/
KClHIMYP2Bc/+Pj9Q6zctlGgK6T57bUUysvbqSQtR8NEGEKx7OlkJUnBs2ERsOccwTSL4jKvWZmu
qudXGBS+EgPn23MP81l3RrqhmW5dr/bddq8Z/OBB/XBQCrFXFT+MHY5rqM95xowUSuhdpKMQab5e
Hq7PnHvG5tpzx9bj1vbGW2wgBYS7z+dxpDQsEgetCIswXy7lPjYCK7R12DsdIDT4y5HT2ZCN2d2Q
l+0e/1Ce5DXRxgQW4ot5W4Gve/c50Wx92A+mf/DoX/rIvmgESMp2pyNNw6dtFHe7nujkAcYIHvEa
Gm7Z10/hNwxaQcqIQKn6OQkOeJHH8ibPu8EtY8CCbTmxBOrX52YY3xIptsVstBdsJs0LxISShtK/
O+ZulsLnR2NzFtjA/iEXOhANjgY/As62H+n5ETrDGgOLOdEEYzlYif7qmQZC1KIMWGxjhZMHCNYR
OSCKH2/rtinM86bA5uKmBPdt8RgA+c+XpeRU32038LvR9lhFbRJ0I5I5mjTO0xk6sO/psG8dB4Qm
1JjWlc3Yt/knpjv1yKvEAicLmg8JbU+a7qAqaFVgjvhXkYSkqFPTUSXyxWx5Uw3s2YNcdMpAPtiQ
zzbXNsgK+0r8J22SYql65C/XDS3LFSbpjNSrht15e3fNVxwYueu4BgLNxnWKr9txeUSMF69x14JC
aXnm4NIdVhYmzCUdy9cfz4TOibfDd5vhQjeSKHHATQ4dCxJlasLxrGvPEtufkspB8ACkODy3wVKz
x/hfSEqkfeRXYwqpnJBnBJNjBU+cASV5UynV2DIgu/NCUTDeWoH72Ee92Mhzq0Hj5wsMo/v/Z13n
5WlX2SS9/qxF4f2lfnOEk+/YqEn0haNGUFroSKMONd745nUEUIprIT33H6fFYajvuPaTnMlte3MQ
G3R1y3s01PE3MdgB8eDw/5gij3i3g7dovGaLtlz71g/XBHjpQJqXXygVZD8hqawJVYpE0k92+MbD
CzSPUJHUOJyV38bZMFnNLVID4k+Udoh/sRQQpu56bvvOlwZc2FusdQqq2k0oBupVi2jJhcTI3i1i
8++YJszQPppU8o9s90aMDLeD9Cbvkx4S3Y/nu8N5zhEfB81jtgdzRqsqtg2wWWWi6KJiL101CEeH
t7QSfGSH2y9/FIUO7H0P70nGeNJ10N70JzJ8OW8CP+gwU/B4fkqmX6iFQ1NnI5zqSU7HarQyns5A
h8ln+9TKQZeqaLXv7RtThybH2P5vt24U17vfdR4spnFkZVCJtpV5lsLW5LqCwkZScWA2nLEfpdpc
thmtNeqCZOEhEODj9QXxhMoRY+xCeFFDuqksbndLNNSsCynTb2/I7OaXn+f9k0NLuD9Ot47jDGGf
UZWyyI+HX0rysDlu5Hr6JFUTHqiY4J5TPa3nnfxryBMHWM/T8H6+SYwymBcz6wfGYY2aazoXzan/
ei015Jhr0xLxRWc3L7nDmI6FCbXES+Tm6M4pWFatVzmH8WTO+pjdSgdfFIJTZeeNDCtxtfCG7C3y
cDBFkZL7n2ys4SL+S66LZhQVjjqKkCt1KSKWKxbcu9Y2AU45juRo3p5V0rKN+SM2AVgEP9HfzVjz
3JRXWQVMXXvyXVfBKkKa5oByxjd0khIKI65wceRh6pytp0I29o8W3UVX+tjUhma+kITZavq9qBk/
cYz5yHWmGFVJoYGROoLYtsNNm8dNUiDF2pYCc23c6vjrUp63khcuemGJsfCJMTZbaJxWppXrmzfr
dt6ePNRpM8T8DVbtieSYhYf+McJ5di8CGgd596vOSjc0al1jiVgBybP87Q5jpp6iosOSGSri11tS
McL4OhqulCpnUIVEFKR3t6EZi3aNmLzQf4TylMqlfA7v3squiMl8d/Rc0h8k3Sr6jzz4ebAU46WK
SD/YPd679iK6YBF0jFmmqzBQlqj5s/wXNzWT18ahJElnoQR5a4blEtGJH2h8fnDFw6afqicPi3Gw
USfnQKPU2pClNp7ioUzGtbg7rebgQCYzW7Ao8p5LdyNqAyxu+TGn0cBufgAwGZPn54tRU547RIde
NtLTsZC5rEPTEq7F1hiA9oFhpg+1rI6ZMkuAqJIKihzrjCYta/c+5QcpFPOsXHSCQjIPIT702CcS
wI0l2xoW1qtxN8EWZtTrKqxyBgQxLkgKWzNK6r0RRV8ZXVFsAiGys7f8A0oZMRZFWsTHBXzmb5EA
hRzCOr4Hh0dHTkSJzaspLFoCYM5pifH0a1u7znB7MzkMwyBNKkMorzvFFrIYAa4I2nZHWGzwmwDk
yotziXzFqAhMKzgK7f69Nyr8s5buCad4RreY4zBDZbnNOYWuDS1YlnQWiOGO2rhiPAIlDCozr37U
r+29oinhjvvsliCL1zjV9H+EdrOKztkR4Tj1+uNzSuAPqFh36c5ytsDVmB4adRQ+AzTNgQ3LGf1G
etEsZi39/RhC5TyqJtmM0jyZ9ktBoZCid4Sch9i+YAVTwtREY0SgzVBW/OAibNZVqRwCb8Vertap
lsxckwyBxfhGmhwNzIbnfPdZCuuz+oCwYc6zdcqG4zuguTiPJ/RGUietq9Nf3zaVFExdQLfWU79G
u1Y3/3s2CdsYBKPUNI/3QS+06OoSfY7pqneEont/1shUOJ4m5YYH/1nIMG/bnZH1dwkcn4OuRXj8
6P9qzgrDM6b0SMqqisVqLnyNcaGbXD78GPW452sBS5EpDQg1pdRFKHotPZVtVu/7GySPP7rgqDx0
nP5lNmyrXy0k8IGbamxtG0sJ+BK3hWtDlFEbVcykV/iozPReJywZ0zbNd+NCZRW1VN+1LvUMZOui
aDx9NrSmqZZ2qwSXR8B3W2wMTsvAgPzjfnQsWBQiGetyL27dBQBaHubBcScMMQgHQ/+VFJcdJ09O
zoR4LC8ZGlvSAw01vFVfmXWPUyF/Ck0Th7lylk+haUILVpZZKl4U5wdm7dqYl403GgrHO5oYOiZj
MIJfUr33rN3el0T35zDgeTGla5paB0d39g11B95iVh1SLZ1RCa59aZkK85t3K8LOY1OFWIKf2bpW
FUoqFLonTfZrrz7+1LxYQLDITIn9izQpLhn+pj3Q6fOulU5JobXxY7qWU/fPFFkTuTJ+qvOf4ixP
926MSIv0eGwx3uglWS4VH8173aokOgaTCL09w8LCJOOD1Tr+NOrwXKNRhS3zL1CDVZcGYSDDbAjp
2jdGsrf3vWz/yHpjuiKk0EngR7YJ2kFoxP9csFgVOTvObJMNIU05sjqRYbTW0iVfGPALDHjQP/5R
GRiSuVwduMyIpvQ4GmPlh9uS2WmVDJTPrDlgPA/rQpqHj5MHiZQxjrU512nASV9fVaJ3hNrLO04U
c7KSC5E6f6O+zk8iBJEJ4T7y3ADO5K4q/oyBfDU/SvDxzYz0fl6c9gIXCEDlSPBamk3HPZ5fPnrR
DRmZq8TjV0ySRurolge9k6PXfilWN1++Xxw/GecC+kzm3KTXDZaOjSDIia/dgbmk4zI7FVW8NxgE
VXNN5dR3zpHbRLAkVrKuScCmZ0Zev7nRdeZw9FFeoE4pAC2Ggs++T7xrHhoDZQMD1cG1r5eEP8RJ
CgSuVY0Hnf6jMmuHDlzi7TL/2ZSzkX/Aj+KjaQPdHGv9oLgrL5z/giX9EFc3CZSeQN0RO+GGbbYi
Omw8EgwPfnmHroX4MjVdm2gmtlQuQfjp22dZsW05HpMqFlARvkUYe7NYra9wFJq4ZsC2N9j2E+sA
QtmnbA0D06/5VmH0OBnPvcPl0ilvAKUTWrIluSMB4SnA4UZkfuOW/CWKwUqd/T0RrB+xBj8/9eBj
Myc3R2XxB6Z2iQEe5zEBsvAFxECijZuCTeWaWzMlDbLpo+y6wqL67gXuXmWKV4zrRuWdzyY0wJ67
JWVB1NuJ9bMOMGGaAHOnIzWbpzrh+Z9UMPQo28xo9ra+3oj5QsPhFeM6mdDozK5vKZMRfa0TECZu
OajZK3h1oK1o0RwYEW0CJmajxY+Bmu8VkiL/YXllnTJKgCqTDcuRxookjEI/79iZ+MvG+xYmzw8g
J2zGpGrj69Z6FFcIegRl4F0hCsTGRNZOYoYR4+wDCrB3nxf+7uCMH1nu4GmRNDr2rwL3VvzAM0Uk
gvUvM+2Jir36VObujPHVQ8hTBCH38eud8GnP+w7SCqz99wGlJXOgFK8dvfB/o456pq9PV5PL5016
CaANlRryrH8ubdCFlzwL7mf4MR6DVv9WYa6a55WYG+eJjXzMcWNw6f4YV1RZFayZ8aE8U9Bn4wlW
hoExmw8vPgIRZv7Rc2wKvcRU4KlEWfEFG3BWB8KOu5LanICuvujoELl8ibA8kLfSI31vDknVjfi7
mIvXew3ua67bhKbHlP6gH8YAzR6kSZH2CJH8Ztn9n7zYZLdgMVELm970CxsNn4wF2fzDwjlZp62A
z+VqJnTVgQXpIY8GzHmxUbL23VdBDavPHbG/9E6eWiTR36BoB3wR8kN6fxN+uhYOetJuZbmua8gW
AvJcoKmAb5sClZySpyfyvgCUbpYQYYgPVbCba6gUerdBLbDgASgVDNUWg5EDcLcpbH8Flk9RoZrW
960rMIwkkO9EFotZjmpVuR83p5OGXUzR2iUyF18vEI8rJVtuDyqw4hxFUnEjOcJUPF/3GQfE1xeU
TTgacyacXfctAC1T+KubPlzT5+FWwoK1Y305Hxw9jc8jNujh5TWpc6U8yK2TCeYY3IgtboosDno8
UaJgKMoUE3sCGIpwcOHrKsacX+r4oDBeSuIoqa6y1G2ZV47iLxeWYzJBhYs7nQQRt0aNFHH3H+9a
mVCPaIiJKZs9NjMhpROTYxNBq5lIuCVWY/eyzCb9EJGhY+g7aFIlxo5rCiRgkncGeKKmFPvvC7dj
/OPe54JtNCat5gJqh0RTj11ZyPTs8z5bGq4DWKEdEPBnFGI6q03EGbpxCEqXwCo8m3zodutpfeGb
NfWojAtCnjRUMJ56vfDSU+wMe1F6vDMsnrRsYadU8qj4cSZwk2jJbfpzyV12gq3Uq2RqHWzCRN2j
0UXgFn1YPuDO/raXx+E/92DZ258/uOnMzhwYs2tDX4ugmyX2kZKwR8UjopCMyKx48/lWZtqdRRlB
OcShQKm5p7QRsi/tpJhI2yRY11ynpjJsjXgkNKXaESOTx9ANZr14uqC1B13X1DD3zkGxMuto+PvM
ZLk1V+MjIJBcCkjMgX6kDuvhoUW+mFGoyqFtIRaY09KgwMUrPQleYA3bF861nFCCCsb3rIc6peqT
lJZkRYdy/PCaWls/RaWANKgT2Q39lDB5o/iL786OaLkcI51LcPswALDDUDxoO4ayb6UsqJQnA5Ff
HnpqR0xkYkZscsMN1wNFQXsoOrgvb/u/lidabJOyceUNkh7IiRm4ywmbQOed9MLZx+0wDMY8qP3z
4VMJrlGVadBIksAL+URcpnvWvcIEovne/vlPrIJhCRc8B4NRhCjIBRtTiy3mrxVEi5Bwj3/I34PB
pk1Mrco3FBx+KZBaFuGLot75xHlNvL1uFXoeLEgMuMW18CYiqrC6LcwVOPyb4wf4NBq5aYzjZEBx
b2Lq3uzKpLJhVli7sOBMe8Toa9I0yDYl3eQ+Y1FE9EbnlMu6s3Drgr08F+2nCdQFtikKrWTZ+1TN
PT8yE5nEL0qqWHWc+j0tkp6Wa82fbP7uir27uyP++4/Jj0GarcuemQ5skCGuzeoaaL1vEYC/0yvs
R4Vhyld3RDpCD8vZggdpS7/qzVwRRPdvHrRYIi5fkIqQTCgJh7AJf/tZIzjOcpdw5tcNPF+l7smq
yJydi3R96g3DxoQvhZo1+Ie8uelBpU3ScCg6jYo3OwGvub0Q30fbR5JFfm8hAUyDwxkVtFBTdwWc
fmAkzGTeSWYQtL9QHTpraQ6h7ecvQcshLex5q2OhndVD1R/Plc1Ec+MPNg99PdMJnzkD0OEzuZKl
zrK161IczPq/dSZ9hU2fIDeNnzIKDBri25DqM1uJoL4M26e8bjbwRm2/4ZjwB+KvjAXn/dCkbt2c
VCj+XCmplahul/uXZnd9tikwO0eailjkCruBsZY1ox7AHsM5TewQdMzAK9Ho8foXU4NjAISmAtaR
T0P5B1cjkEZ8MMlP54R+yaXJvtDp6a6WueME5Q0g8fQfE4/2rL/Uz288TpOkC5AYF/qXcZhjv633
0bn8kYPTS0o7CK2fIHtTxgSAjahVMPNAjRmfAqK2WXbuun2WcHVsbPnfjdoHMxh0oDGwzjukpJIr
CURQiDCqa9fR0xKFhtj6cFivGjFFTHV1k1FwZMXxvnWTSfZvUr2AECOg37ThuSbx+QIZViiAmvdD
/CWSXD+03q+yGcOlGfqTE/uN5e9PLgxoH/ZZpzTypB9N4ZqnFX10rz0T8HD2q9FV+kflEd9lM/ZB
vhY2gKRd2LVnbKKXvuGPNqrQOIfRdQIJ2WkX5PPHdtrqzSe1bVW+t/UCWBi1QBQJFV09cClpceQz
A/I2YtlrZoPq9VtQ2w2sl3yQ5FoumRNhRAZSq+AUDjDP81ZoiWnscFKogtzLFRxn8k/Aode5YSKu
Hl+UwFasAYiRADQtt9QQqkw6UniFI7x1gmSqzsVuKzTEM1bwtdMTKekwbdmu0uRYAgp7rKt3XQnB
KCDFDmQjXLd48NqC4NnLk3NdTxAGCyG0TMmYIY9CoicaLLi+ZiVcuqtwGBWtxMF8kcpzRSLC8+sD
+k0Rn1O1IxXBmTZ5Uhooql8a+pREKCZ4pMV2cBpJnVKVMYFprBdW7FIVmPxX2IR2qSAzTz1yp/NN
Ph7iOqU0iua3Z2lSL7e2YigOFLxLDXKah0t8lH4WtsP46HvuBAUjKjk6feVslRdeWoAn+in6GcRv
oyqRcFbBdvLs2IlFWjGBTQVPlaBP7qkXxu2i9KobjDFnmvmeKTsjbmk0KZw+phQY+cEKDRE8iXIA
4wq9RzLaZEjBbX8422XoYT+OVRNnCar4euobeEzQMm0H36rFWBnOig7K0WI4+7NfIw3C8KOzWy1l
lsGaOWBB92DDxWHUoiyh5Yj1yRUyOB3wkvqBiPfB4R0E6yXRCHS4wZQezUb+DvDv0VFkDzWieak/
aJCNaa90QYKjnl7SdW1t8A0sT5Bded+eGlyZm9pQGzhUXRlFg83GqzUn1j06WJ3Sz09LixlnrcMd
UHfcZzVvc6A8liuXUJ90+hT9n9rOLdlXAY/D7GOvqUHLVEC7RmU+X6/Prd7QPAd7fRFkSBjdWh8Z
WNgcHLVrOMHtmRaKhOvPTZ94EkphvNxQdoHwyux6twC6v+zI26sF0c3hW+GGhsCTsirFiiiplY05
je6dwFa67wzRCXaI8zzt9rhVt6K7Nhq9a1tVFv0X9pgnpJm+LuRGZR5c4L+FoKpDixy/STgcfvr5
yYXKnL99GhYNppjkyqV8nG/jmhfl8GhhAMxbUYeuwn6wTph3GFhX1W0HP2EMLKi6cVXpHqf6s7ku
2aSjca2AAzSyE79wx9uhhpruCTnyk11OHdgBt6V5nFVwnvN8VEqKlk5oELzG3rTtXkaLdBLswnYz
nX+l4j9y9z0rv+63VTCUa7fJQ72Fet+lxREwQhy2kogEivRzv8lZaAs7XCBG2bhDd6jz4g8i6Ht6
NDGIb8jWrHrsRD6HEWG9hmfHlPudyZqFhkuh7VfTAyE+aD+hFhifyJ/bdgPU+rpsRLtKfj9Z0nWx
RDMY/+npvAGiT3QAd69M1UwtJF1PZSmPuz7YvlZcR76Hc/+vM7xD1VfRVooED1o231jLEFjMVP7S
Snp2v+GgRheZNIatdY3qmwwBjOAzd4LJJIebF7TsExrY6LKEUBXwx3V+BKjQHrDEggymjCggQIiW
2Kx/KxnHWyUiPnAp0K90rVwDkfYkQUSDF3iMRL/Yj7VUInMIySb3wItPlR8KOQxdDFVDSjPvKYLr
bX4ybFf9T9MKrAq7lVAOw9Pm1l9EdjPrDvV5IAnhhertrQsYBKs8VATr796SU41N1nq6M1FPCm5s
Uz2EKxH8sqU31nZcJWTyXgfGn3ewLfjtTSaJpNDX1sqx5u9iH105Jxc0hy1Rvs+ascPXc/SPUM8F
aM2O36FvbyBGXtLhpmnPR4je1clV3cXkACAuDoBmuYF9+60DEYrFyUrCcC2TRKHb4/HVe8Va++D1
6Su2c2EAS934ZxSuCTahdodwcJxcj6zWY9Dkjc22kek9BZAz0enHJJhEIIla4htyT/vjwc8a+BQk
EU+SjfLV4lofj1Qm/u8+Bi15eeGx9x4sXs49mvSR+4kJY52dLEqIK7LY3wltWHSCQX5OcJV9l8XR
B3ivKfr4/gTcvDLGYbKiwN7lGaOeXZYIjl4GxWFk2oJNqjzr6cJ0SC8jbGrmBqNrdRYUSOP9X5cm
JW3PRQjxCu7+VnNz8dedbXtkwwGgoVEhieq3TAnbN5fu/EjuQfAOl7osJt2725DWdSmVoz3PHp+Q
Ofj0VCwrM8yKd4AO4/xqZvpAosDy2xfTPjW4U5ipcWCf5pdsD62vEsHb+r9zwlEDop5mKQolSqvs
iRdlBQt/WNomp7IeY55UYffQy+AGSKMxsbV6LD7wXFuczH5nCpR7DjafJpf7gWLxBHO+6+Ug7974
P/NB5LoJMUF2JEkInBdd1vbn2xI3NXHA4LfRoT7s0Il5i4AgM5+ih3LHEiqmMbz9HXOawNM91onn
0ZFHRSekYOR+t0C7XZDp/1x85U+iEF0OJUub3bhztNAmB7TvMeMNY1yLxOc/TVrbrYvoIF1hyNVT
wFTh+ulnC4xvrXNHy78FnpaaYCwCny8N++p4t9SZgH7bGNPrGJ6ZnlkGh6e/VRl1UfP6aVZPjnzn
fKr2ikpeA26D9hqas83+lZk8QbJrxQGbfsRf8t9v6U+ps5NnVDSqgxuRm0VJYDrlKOm5VObDaoGz
tifZwUPnVmSKeiVPrCW5ef/X4MkjR3msP4GlGXdVDlLf0XxjFN060/4htrp3tRvWJalhKHC68r/f
g8o5512iROxQ1/xvewhggAGu/lI1AF7r9k+Qad5xp+mG4OfotXwXGYstE3rnEAjuaJ0vqsYCdpKC
lqQxBpKsLDSzvy+Y8be3UD5l9gQFP6ftsh+kxtH79PtHeODJZqv1jnDVFc0DOhw8tPugLzv82XXD
HEFsbCmH4kTwPusVDoaLv4E66Dz9DbLW5T9SQEswrKZJYRn+r2DPd0yrV5W1vRqsWzas9IEW082C
GODp//q5pL+KlUzldw4sMStWzcpV9R/HncDUUDBWb+S4SlSopeeMigLdBKyUJ76SAb17ErFau4aW
vVKPSaffZd6MDt1Fr6/Ck+Axa7MqIhXAqMIsyCdAq6PhwJVVTYueyICYV512IsFF0g4bJOmAyFWq
XD8uN2Ya01H/98l9zNoTEggemZK/s0H9ElFM3L+GQg0EC6Y7jfO+1svjYMS1eS+cufjfZzEqoA1T
eoqwNbVRjlpn3Lql5ZR0EQh6DYDSMwRIr7UyZCkAGaHLa6TxnrKuQU1Rj4SCKpzP8LiRA+Av3zNp
fTiC+10fT/zT5plXlwDYNgp3yZudVzgHLrkrv8ymD2hnK4443RFLl94xLdzFRSqvxromdhrmDFxP
v9ytwRoalxzLtfFt7CBFoGo/DUJe2PHcx30YgokTRBUfEjiHgOqTqTjJlUYKMDhXV8KGy5ITeM9P
larj/4X4Rrq/Ul4NiNbM040+ZG3dl8tG+p3wnkiomplKZkfPihYfEpyCvRK1pfTFyA1S562ulD8n
SReZw/03kofyk8v8R5Ik8zfloWuMkDwG1Bx1q1ateSpYfQ1cNevpR+eSb9c/4FoQfJ9uJV5wSE8G
7F+fFWZFy3ZuffenCFy7YwpcJVk9zyJ7+u92+XUjmCW78hlWhIQIqEfAm2sp8AnnpGNbk0yEBAsh
zh5Xd2uaKDbANGQN7NdI4rzesKO+3D6bHyR9d9sCRcwtMftXdtOggBSsrtDrkK+C4mMLSVw7xzlD
WWTsGuJl24srz+ZRAW53fEZ+ZxhTq6EfBdgjr/qhelKWajKkW/SOGRhRQseRCH16KgjXUIsrAk7E
ctAYLXyuzLkwLLQR2H08bEkSeHBFzxFotmWbaWgdxl9L8ViVOXmILm/sjk3Vi8AEtQr9vdvH92l5
qNG5U4QN/uh4UW06Bv4eeQGXOvnhfPnJ+/bBrdCzq8pPUtA1TV3t3/S3Lo5E67AvYtT0Sm0P9T8C
cdwN5drHWhIqNaTnLXiey9MJmor03I+Nw0CLg8n4RmkNJtN29NUJOhOgqhpyzJxhaKSB9k+0KsCP
i05ld4UsjEw1fjxi4MLYMHv+nlL0jtER6bT1EVx9m2FxygKbbV4L2QamncYxUPOsodGFT/CE2tQ9
LGllo7uAQmzIAT+BoWwuFqRWJhVthSdK0kiXJjSk5/mD/48QJjTcicLMDqZj5zIWzOlwsT8XfLMI
jYnaNHjEke3gZ2GQDrwzlq+4FaSCwUo5+f2SzIl6DXB5im0jKLtpCGcUyVsXaAdy/riy2PgDWZGt
QVK+qJWVj0Izkq9o6XKMlslruGLLIJxHvkLgzLS0y3sNRuhOdIDzJG2boIFVLKflfEFv15h0+Spm
pCb5DoSkfW3XWMmX/LED8Obe+ipzcBCRlNmvrK2FZKVKmZwsZfB9Z6Y/zlHv+vTttTpTOXi4E/Si
NBWqB2/yMZRY1P7WvSIeJBnwT9SqtkrEVAe7FRr56EFO9zGt1fwHyAnDieZvlBzN82S0EQMHB5An
cEPyAJ/zfGWmTESB6vML4zyfoH8yXe1eo4O2ZIVQHRqp+/cp3AQ1s4GAgoGiC+dETkkulFSbbS3I
W2N7hvccXJDqDEGekbocx35bSqPHisronJuKBLXo7UUQuKMYhl4hw8Ir3XOy4gxcpDhtE1xoa+U+
Oy1aOWpMZ5tfmZZDNuFonCs4cuXKvMBs3XE42y7V15ymnyxrWSJmOfxXQ9PMvq6Jz9MI7aHqvmVi
HE/PoZ5XFHOMieeObAb+DQSq6kSDlLxcSAFl6nO68+/3UybjvwKRkQt5mmUggiuOBl52Wf4JlMY+
JQph/ZbMMJ7kM990EJnc6n3iCAj2YgLefaSOE8iT2MN9cImwd2q9Ns94rR3U0e7xrkIdm6sKDOBF
K0okzTKDAIygOPLzzyBSeBEF+nc5+lJ0Itk+4f8zNDhil7nObkCEf3ZTddWqgbvXjulXSYsJY8Xe
CPdzaxUG3bkZKlJnAfunW7yH+p8Do8IXakmwX4J4xcDSGVCP95vgN5Ze0eY7haNWoQOjZVGU5NFf
vluYxM4TshwhCPqe2nffy0gsrR20m2lQjE/5YzHcTy493243mPkgQ0cYhooEmIoQr0X8153LtT90
lNuw5nc38BedDXWd5cbvB6DQjUCp8EMjtitIaQFUDDuniYKZxPbL+/+lvxqa123X3nxnPlEqG74o
G5xCDTdLS//BxjOi0LjEnexaklVu4dmbwuBiX9JDg6TS4to16JcI9AQGZI8o3ZZu+Nvt0yWKqQZ/
EXoQbkJKl8k5Z1/nLSU6OgBIStDiX5SEm8dYtCd+lvzAr38DQV1crom4LAi3mGUeshOZoAeR5qQb
kPcKmefqZps7GUO01f3GMT/HpjpIjKA/KGfglUVJYNRg4yChP9813RLcz1C3lRoeuZ8V0WBczoib
ttZoHtu5tn1xmdUFwdvgR5uDls9bn24Pq+mPf/MNPDQVTQ+9/Q43Ymkthk0KekHDOEtHS4ylTkt8
9DTTPvHJuWSc039ewFO5YVLJwE4qLCrDZOhinK2wZPjBlsBATfJPtT2L8ywT+rChsp8aouW4yE+F
oZcTMCVZeOq+wRZ/kqWuO61Y0Z6G7IReTyIHhQAhvPBs5/05x+BUJJObICbZQhNuX7v/5L+LX4e8
+v3FWxZFKFAreX+ow4Hy8EPIZxYo5Ytv1lK7kA0CqeNEnT8TMbJOKAmx6mXn1+IbTzCCqh+irFSL
QkFXsK3kSaq5qpYS2nzXlTu5mUMJtTL3oaOn/cg2xUkwKt5FeUDoVyUIYDW1eItOUA1s27BY5wek
jaJ+fjUMU6KR3ueQB8pWPyrBWZ4MfsLm1ZKCjaZIzt2yqREeCHrVnSEPvolTKo5k3VkxT7XXMvmt
8gzuHBj8HK+V9IqqexpXVHbRgBBYmMFADK4gt9KM5EdfM1FZYtlWwoA0sh/p8/ovcyKPb/wqReMS
AunsCApxzFcPFSElrjbAsR2aS8ful0htMEot7eYBwkkwNWtXd7KKT29XMn96zOHc7StFpu3LU6yU
efBRvI8bO/yyhnMJY/UXCKatGudsQxWp0hXEsWO9QdHpDW6W9ZPcJtze1sMi1wWW+Djak4qOamfC
h/ZoIZyMkGqG3zLT2jkgvAAbcZguIFLqwtFhy5iEKkNj9ki/th1n/HKlsbr6Y4BjstotzXh/F+hI
fioKqk5aEIU/qHCM3an5L5DX2F2L+8EjvM2rkEJm6tDqDvvRlS8VaBv6x99iIOM104YipxE/5Fvr
Dskm1GPVQ7vqOCl/6WjTWrjTbvNqfa5l20V3S+V+cstA30w/JwpXh8JeL36nCOCUsZ1o7hzpmbf5
tG6GK0UOdo3j47PWDg2eWNAtJ+tMA7KB2gyQA6dkJQCdK1FAk6pRXG5izXIdH65bY25DIfJzck5f
Q5wXGWG/g7LOoBtgIv3BVfYQvfmhstGKAYpVokLw/9blkmdIWqLH1gHJ3lqcyCw1HNfj77UvB14j
XQpC2+RxdDW0HnCW+qSyMIzQ/XXuHsHGNhWwhrvswE/a649qdgzV20G2xfTKED66U7/cgvkaFzTl
JJ+TC/NEP4IPaRtHoCJwcDI5ngp8D+B73EThMlNsDOBZNumVNcwsMgcutyrWgEskHqEMhK7ERZc4
7zwekiV2aO4Xg2xnlVSNJOa1KiFvC+y8RZmqtzpiHpLkk+3iDJujrpKAEFy2YyCq2e7YRbP5d6IE
JmZFkbJTXBzt5uO+vsVBOnWAmp35vJe4Sfvp8tmbNV0ylxyEqY8oXPzHj4WGjGp/kL46bl0HcAvd
MEKMnUdPjLvLKULOeug90deKbaZFOjNWCEK2S9aW3T6zE0pcv5P3nm9ggXTbb9jepK8JW92Le2Hk
meg8wSOl8CY1+DTdvoiM3NzXqC/EV+c1zDuFch7TIC/y3NZFi/IjQFsUn6epvCzeyWsw+glddMc+
e+vtxjMRTxmksR8K+4BsggYMVyr7t/y3j6zr/xnYVlQrUxP2FQ2VO5Ukmktj1YxKxS+fN184vcet
RoqRMB8TLckmlbX3kHuHXyy8YX+efTKeWRSu0X8zV94Xtho9Gei/wo5QEjm1t2qaJwa/6NvDRX1f
wsbNM2BjhUQXFpc7mxkz6K30kvos4GujMO7JQOJg2bb5rwH2MT09it3Hdjl5lVjUlMdGSN8p8M4v
5zmBHIGJ1CdQpCtFhNbqJ7qdGLytLoolmBgl8qDM1rB0XWpCf0NpKpc1s6TEEozQ29JOgELJcnLJ
BYHjmGb2bjcBZtV2wEEpfpOtLgMtbmwxqdB/LUW8jA/FuT61dTgbpU9ogRL7WhATmdr14ObfNh5L
japy16hRNxj2iyzy6fz8HNkMQKTyg7WrEbxrS/zVzYFEgY0YfJZCshr0gi++G9x9K72rvcF9WqsL
+nKavERLIiabyp8duXWhP08REWIPcI0K+LJS/+LzYyxHh6bvq9KnP37IeOROItYVdhT9/MLGS8ez
6cu/Osb+cwxSbDmY4dyy1TtU58JEUCbTD+JLx0+4JS2NotKod4QkkMHvWSXY5jRGhMtJSOId0WEl
g2Jg1CORUxQawqg3VPZ0p3WNV9BkIcCv9nCwssDYfwxPXWvhhyu6UL9PJBpnxptfO14S3TNWRyB8
vM4r9Y36GOSYb1j2zfThXB8QvLnjgeS5jayib1/2P2yAGl1WY637IiTgZzTttBeAlZ+dSXJODxqH
xb6NHAeGI3DD70MLt1iuX7cej3PTeNuCvENO0zUrH4HxzkNIyxWKtfViKBzRKq010yjstxqF4QHz
wORuU5BVnAwR6v4sJZBIsxX9K6N4XAa+jrFERXbCF65wPVexwRSCv769uwlP4f0cQPFIuAXxsf3z
ZdedQ9WzjAv9i7ryuVmctX563xDfZHN2xnxKCjwOm6elEp04tZbGvOIMfvcMqdpGp0GAEIHO7wB8
Uy1h3GlK2Scs2iCXZLtw5pJtZVOFqKkEkF2qvrZ0i5oGizQFq6bALTOYkePtoSY2S1GaKKCqJ5Ge
sxDtzsFQMtsyX9cS8L6gJ7mr+1H4Pk07guq4+eJNxFEy2yNivO5uNJGssSMwR0t8+6PmVb4kLcTW
YjVBt7s6batLorGtAej2ecZodMymaxja6fkTpbO0khWm5wL/3cAGcK5eE7VbFCyP913XO4VqRNZF
wAYR2Ka0bouFal+PZDaaELzDgvh/TjEAalq7OegBSN2tBBYnBKoeFgJ1E/7h2qW2F0KpeW6iOE8T
EDrIGFLIWhpFwk7zDCRI2hTuOV+1kr7mYbPW4ljmtC6vqo7qviXuL3Xse7p5RpUyXLaQAFn39s4B
HeUGgVNeNEl/O/qPNlIM13RI3U0p55rOqXUedn/k6mmo6TlGvCAWuS/H7coxdzy0Aj3MiryQkmJv
Oy2Pgia4irerH0E/YEUJ/G5vOmHK8uAJ453mES6xMBzSsMtISxaKTqF9HnBl+DgusSpO36wOj1OQ
tvtNVrXb36I8JhIFKG2NQ9OYSLzMGZkDrLz/10e92q7sV+P+3QK9/AQsp9gHodUREojrNbPQSH0I
RY0AwbUiGGYkSVIO20JGJhs7w+NTbV69+YRQUlfJSALlr89RQ0eMUWjsxbEAyBDau3AWFLmA1ecI
UBTKymO2f6AU5ouUXi+NQoxiyaSRUXQQzTOD12gKXZ91/GkC5t2DjrVZ5rYJglDQOBScSwJwKuom
TUDi5kX5vSnwA5qz1heERnu94RxiXipzr8TyWWWF3TMyXcAbmpQDYA6lpii8l1Dmtdvw7Pcjzk7Q
xBS0L9NGXSqweaIYsaN2JQNTqDy8PDoFBYTQmi/51QmDhlGRr8ApWGM1mkN+W1Mj2SA2fRWqWWc7
S1jDXdX9fasmmkWFCdM6cHRE7SheLtQLyptP1ZBaTWtPi7uHZIFIrgzlzYSwTN62J3+msvNA4SG3
Ic4RBQH6JV+IbUw34LclDugPr+OnjY+B9Ouwrb1xeXR5a+u0bIADb8MmiOf7HZ/xFAFdQodm2eF0
szhaigdIfXOafYe9+EbeU23IYMwUskOnaUF23u9NMBp/0lIBTV4wFcmZ6z0B4fxSli8G2qw6KrMJ
4iCZMBs7zsB51GvcbhKjO96104KW0r3xw3eBpBiKEJ2grW0A4/f3Yq89AaBDd0/3Q/X2ew8q9hH+
OFUXhSTa/Cu7jrGZqUeKE3j3qNND2czbkFZ1FLAE94x1/3nYgdsNkOpeDyMnzQwDYxUXDJJQ1pOc
L9H0rfnZgIQg36MmIvv4KGWHTn05Rxe+NChk1lXNDX4QF0f0lrrAwmQ2EK17+pNspypgKsuDMdty
E7jI7AJ/bKzkwtGP9Qcmz3X+XMy59rgSz4dvMD4XZDk77RRjgqfL09+84KiG4+aR2X+eLICX4K/c
oL9r4aMfiTSYEf4s7PfEKxLhphsBMlHcS8WRuG0d/RL0VExSD4hFOowIIxp/bPkTXfYexCMXbZHO
wZFkkDR4i+4o+Y0RkFNBhww1VQZp3uuM4hzQFIrU/uAaRhJYmxnjQEZeHP02w2/mHQc8XZ0SS53Z
yIn+zuAZFVIP/6fgcAEik+WwwhiWO0oph1p/sPP73caTfNl49nnr4IzaUI9HQFIe6RLuNcnNYb4q
jaaPdxH7pIUAJRRLD9F2Bu+qHFsObIWm98bDLVsh1vUamyfDWoHhFWUZnfen3cZjguCW4muZ+PGR
Q6b0o9WqtbjTpdWlgzQo2yHxeo+g8qv6GeKB70x4Y6ZuCEoqn0LMv2AnTI2aPrsQM6bx4ZM79i+e
IUwlOeN1VW2uJt3yqz8rgAK7+e7BfogNj/5fmliqQK0lbfikSv+lpJJSOubc2n8dE0XRqbn3iKGu
GcxvXPFkG+GvvUTN7FffrEeePEzb9H6ILM4wYxyxwEcte+/gflMPy76k0ahJqE6mmP6WeJjb8b2A
n6de0YA6foRa83XaouoZ3/uXwNzJbcuYQAdvRa+G9CL0FxQ5TuqtxwypoZ4TIGa/JridlkHEXUTq
DP4Lk1cHiswfXyUSM8NEQHOzwlpinMHzkwTX1EoaaF+vNn57QnAy4tO+OSnwAdGUeCJ1I9PE6pII
Y0AAaiPGsW/lBB2P7wFvoMHXI8y3D9kon078lZF/WoSNvBlBd8Q11IXuZTKvgJqfPUY2Hbg04D7O
jaDdZuYeXI7cEa9iBNG2NM84rdJsVQqq82faFE6r4mdSboC36shUkm8N9+yKv+Q+35LdxbMYwmYr
rcZiAzwg75Doi8SEj1lQVBOWnZFc1Ot0hYXSHydzBI3alu/ag2xez7fDuKVKXveNsNxC88uO8EbV
2AOvQATOo3UmQd5TyJoBjd/ZybVNmouVxh+F4rQX8aVpUw97uxyWfwtgItBXQ6WzPmBXq24wJU+r
gRvPUY3CtUTN4K1Ho2TyPcrV0PvXNTdPexlH/af0nBJKC5TkjILX2jGlEjrHGrMXj7x5NxOBhmoC
4x2R1BeKZclw8pRiyZ10emIGnH9bghp5J/jfwSDrxl/s0CmMGWUcKhXnJ8sLuLf5qrfMEjakSBT5
bvlw7KxURNByi8mFU6gxqp1qVApMeGMT7QC8KRxoyJ+raNL35wXgL+K9Eg7Ib/zdN2lJXsSWuAb/
6NzRdjdnXtXz/5kRo9D+TTfgM1xQ+Zm+uu1LVZF3Ht6efiArdT+JWG20yovD2Nh8BG957s8TbbDq
6sdpyAKKHKg1DRblC69WAAX4/59Wdb+dIP4ucbaQ3RVYTBfGXpplNM2LF4yf88O5eNPVJUetVAlp
8x89tWeLeE1jyqDTeki0ImDMgzptUj2LWEE3yp9OYb+llzBNMHD8EVdpJy0cWrx0lNYkWDuqLRhP
HpwJVNooCcj+11B0XAY/9gxNJoXcOR43nL0BibB2y2RLSSh+XhDKfqSTh9VutxRS+GVYRpvVtprr
ncSTGDKAsuKvpzEZyBKALaHnLJ95PuyLmPCKLMWXlS9+gzuYSelmk8qNrQr4eWUtPa4OZOlvGKDA
yKFcMpKf9CUuSz6JPtiz7yWqM70sblIc93Vct9UCDqZkEzogNZ6UDp/GKRi7yAVnQklE6odBRTwb
VNU9mFHlYdS468nNpF6QeYTjdDba2wqD55cquy3MEtzKyBQeBsn9dtXtvKEPO0KuOD8zVMJsCoGv
5+sQQ1aZtUokPGDkXXdjACKNt8QQBeOtjv6DJ2OVJBR7LglJ8V6XAZY+TLZhi1unx6hX/pXPG3XC
8nox/eexPVcsYWDCwiqBHTXDohT19roq7n9JRAX5ouIkVVXlnLdESr1q7pT5YVQ7sAc8EI+G3eoq
3fj80Qp7aEeVbXWtg3/dRLNJfAAeDjALlWEk9r9M5w9u/cXMXkwlvSj2Mecxlz/P1ATT3eb1Lpjo
Q20QlQ4XT+FFNaGaPcdwR8shjo2+oEEw9Fw6QSoAacQxY7+ANjyebEsD1Q6Ah8/aScwB9VPVTw5R
H53AScVobMi5ak+bQ4CtSmnMctgT7A6lMLE8gUKBH/5piVP9UbDPv6TMuroHtDxFGDMHLoYopuhu
fWL6E4hsdUchU2ZdVggFjU2sSpZfLjz66EyUZ6FZKnHc3YzoYi9IvlsVc/Eg3qqw4u6QaBmJQyho
0mp8bkzOrO34RtSXacpUUiVIUo3c98vbxDzyQB948H77mtfKSguDCUl1TpfA5uYashcDzhXY+OoL
J96FN6uTRxVzCvvt55gciuUaJJ74m1qrkTAkRxprYbmPpJo7peJioGF6c/z6d4r96boju7NmDYl9
n4upy0HuLWullbJBHkVZJQhA4RfSZ4wRkaLs8HNO1NVZwKXLfzuwNpGc1L3jznR/EsRc1tsn9XLG
v8agVRj988cFS7SUY1WUz4kO6aIpiBGAA4baUBwmh/nngAcEww9X4nyn5c61jmXJm/6pQbmqILme
gmG9Wy+G5XsXA33aLYR6FBp85yc4xkFCOm8n0sWPz7m3O4/JrydzLVIqeqssHY2OB8J2ffwT48xJ
4bQExT4agwdVFG8UPrKJlXN/5kgBQePy5Ye6CLbLp8TUWlxlsWUlKavQS4bKPhSNhFDStdcs3fB4
dykNB4mB79dlRWdsfEFihX7Jvoq2mwM50M6dYKzbMgD7izR2SRuxdNsFBu1t2Vr+CweBB57Xn4NM
ag3xN4Ndju9un2Xgom7mtRQOsxmXTlsQjbjXmi3k8gqb0LL7cMPPpo//yziARJxC2SX0UmUjnjyK
dscVYdA8U0AnFMNCEXU3mhP0sSBKlJA5Oxx6Ysy/Quy/wkHgaihLr+3/tuwTkZ/8ObIs0oQ0Z3nP
ZrIfhWbseW6PdBpO5EFAO4pCOoVBujlQ23fIvd5ntkl9Hr0Q6sD7bnLmRTcDABJA9eYBYlIrtSzq
GeK9nxXO0LiFxcSdn8eGDlyI5jTSSCsAyTSH9Q+GVeBHUWS6KPWCkpYDopfdGgblVYD3RzkPN2ar
Fi7ueN1hZ/xxP/OdX43Se/TUv1tgCIccm/LQAqb/7KAEM70N+qZNPgpWoGVAQmpPQw2voRGzRVUm
8t2r2Q4hv+J5uP0COTQdXGy1EbG++sVcoBOo6mNR5ARYPk66/vTLodTXxzLKof83BmWXjrOrQVdh
01fCilXxf87XK74TjIYSSCXOpDkIFPoW3/7ByZWzWYirxI4yw3V96w32bVXXeA3tEssqrhabYG/M
0cmi4R4SgbK7RnjuOwib4SnkhWoczfjkF4sn/917X+ekJYUJsU6d8X5R3KIMg05rS0zD93Ur7N9o
mIWaAA/9Vxd4K+RK8/3bcQGxBXpzcaNMIN3kt2QsIpf6rA9/7VZuXLcgVaiejN9cgJPLRMCHM7ZJ
4sYkX/xzZ7/kowXxXzlql3en1ndL65tSRUdQm35Vb8H6q4G4vj6bQdso9W1L/0qJTnsHzPuafnt/
tISPA6KygC3lPszA54on2JCrfKYZlaz9NgNXL96L15d76uH+9rzjhkeDa0OfFYwuYNZK3S++5JSL
97Ot0x8d7I4L83EI8f0L3jkn7J1h5Q8G9WDe+ziFnM7cAIE2dLDZqDk7mVSOivSBwDEk3D5EJcmm
3/1nkWkkriukMNs+cmSoHJnqVUd+no/9u4MrYLUZroU+J4GbBqcpAVfjBb+QM5GAjvYX8iZHxcQD
nJNdWiIw5IYQvmGuVhUoaf/x+aP+Z7R3KWazKPuytIDOgVfrP6MWlWcnYD+rHb/Sn4qMBH3t3sHe
OBZ1Wb3cRmmpfy5lIRIkFFp2xArfYHO3iNRk1U41exuzytC9CqvK8TM/yLNcQGYkzInPTmf70KeY
GV4nJsQcj65lZG8sDn8Xl6DaItQ3FRf79oUVGodAFrm69OYUHHIlL6GsLBLHqnnQqcQOnatov7D1
tt1Lv2keg1YZQitsjSVe/dM0LTuPGN3WGCv814u6HePyGNTNuEL0kp3zDGqmjNw5/9ZNb57xRh6z
+7UW98mSiugDBanJoaNDxGTLPgni6oWCLK1OzAHYsxfP5pj6i2S9Uhq8HF61D5CwfayPCQhCDC5b
nkQkRaX5Bq5oEYcNX75mMpm6h8cS4rTrJPnpnkhrQSVpXq/26dMY7kVC5C2IZg74k1onOcdNzt1o
AwCrN5fOcUQiAVad81vjQXO0da9gkqxLS/HneU5rVT/pbhp2LMYgS/XqBA7nwonzS6RnIJ+sF1qf
XIVoGCGo4FHngdVH9miZumScN7JXP2ZD+AWMFYjvYeJENOh3gOSTIITBWgh32kM1ifLPZyleoSmR
J/CMPPnbKngDRkW0+vqWeJbB/eDbSm3Vqcr1Ff63DLwrCDNKhJZf8hn2Qi5paNsscQ6mck6BB39y
GLZJDc/2dOtg7T3Jwl3b0WhnM3MTo4i1YbHQprvHDZtgQNe8tQiPjabqaPX1x5kvjYmS6YqLIHIS
p3qK/j4R3hZsdfPpxbOH1OmAP08QnQ3xCt6/qtw8wWTbeNH02lLbxff3Am2DbSEekV8Ge0gfCrZH
gi9mXJcg0FPCqvc5XULXHp0r7JWPOOvRTXZbAtBOsSU8IZhhLFer/GGsMQ8EL2sem1Y4uE3XIvCZ
CMtm8uL8in4oi5yfbfiuAcsV8o0vkgNC48gQAOD69zdSmlIDG1dv1H7cRcfTEJJLfonLSw8EkApP
UFgjVMJSRrHzxAdFtUVM/OHyPRHTLvXSVEaUNpiT/pmlsSyTn0SX83tORQltyGAPo6venU/+jTsC
QlK5nM9MjamxlswltsUAtjAwInPy4k0Aj9Tuvmd0VDZx6vt/MqiITmWlZj3oacuSH0zKTdwcefaW
7Xx5JsRzFv71DlkZWElpOYnMk4jNeZCUhKE+86DZrlT8WyKcM5iUVNVoz+5ate1/hbcKaBXFGIZB
GxNuO0zr25pS7U/rfxeTkBoF4COD4q7YzR1ZpQKGuwlZ3v15bgLFqDM4gCXUdMGrM2LCHufF5wC3
vTVHtcx6Lx3HkyDK04skFWafUtOmb+i4+WcubTx5wKmo00jHV5qdwZvAdgYW2ykttNyCu2e1Vr9z
7X1NKKKXSGnnuRBUTSCbHvItcWnZ9FRN0kPYj8DlgNH1BSf6LeQDxOs9py0QC6Q2DwdpZe0XafRj
kUuRjRxcqsu+uQWQHzivLYLIy+N2W3ZjTwhHo2DDqkejaxUtmNCZvRmDGMhX1z2sCpZiMeb5JUqy
rPRgWFKlymiv+5kXCXqincDBzEJJwPhwNmYPZPwM5Cvk/sKpnqYT16mYSzVit4RkX/PztwCiEo0K
hs5bquNFWmwkx4U9jNPSONDpzwcAQ0ODrwNh6xiNFx944Q5IiGKi2W9yXLpYhtqj+PIwZqT3dYeY
i/WndyrTMwAxLjh0GXylzE5N3XnDCuK3ZDFumrhObCUWnTVqqy9qbXX9b99Hi4l9UqUTAoQd3z5g
gI2jDiCzYmRKOyTb5IUtCYzF8MhejIkRv1DcSBviDQ4g0a59RmbE/hjjpMuJ3D2SsqQbYz9uRup0
vn20dOT70FlYYvyqwzgwbo68ES/QMQZQp/ct+bjZZF3SrVKaha2JjFzg6oM1CLpqM7mx4F746xhS
ILCEF5yuqbBjuqPaQpGCW0jsbyihgg5JORIbMMdSRgp8Th6S6OoeC5mgiE9AVe5Ng6Jou69RrhL0
YvJRiqgsh8C9Nb6L8R+y5KvoMpMMz2vKj2nmof/O5Kuv45c+OiB01wngtBmkiB2vFwYp2p7F1u/Z
sCiifqhDj3mtUHJAuROtlrQIkUaDv88JqnjkUg3mkxyf50V6LKXZaYsW4nWWA+lFNuSSFWJWHLIr
Svd3FrexKdxI9oLYsbz2Wvhk9b8VS2i7EquwwNYrkMdVcK8XmtORdxAk32hMBu5l1oFF4B+aROhg
PEHJK3MID/4h8Yw9Z5QOQo1APvqVKIPTvwlmdP5d4qmfovk1lJ+hcoWpGX42TzQeo9KEF1vybPxs
wZm24rt/cK+0JmV7MkzmOkJlL7ty2DtvmkDsu/PHHDWqX5lq23qCh4BVPsBotzSo/nntuGznJy2b
IFbPYahhBveQmP+kYEg5DfizZ/8hnU8zZjt8DQiWKURKKVjjWiy2wiaBifF7K3npgvSfvBwkIY2T
wx5MXURYi0vPUQrpH8B7rSCJxAj0TrMo5mQcnIXwW7WpeByItX1n+/3YtiWzJVX1rTEtAGrxPQ4S
A+wgk1FGJ9f1GiHjDavAY6QhSxPlqtfUbly2zdD8weUCMLNmSMXps5lcE5tVTBd9xZ/lxlw/zL7j
YnCFokbMvnd54oURqvaBJMML9Er3ekghkA392EOa//KmdBBqSvmVaIs0js1JbUhyxHFwVIUz8JT1
7gG5BvXe58Xd7rP+36B01UBjzIeptgSMQqhZLCzflTXIaub03KwnQaPJ+R9m5oOZ7WciUfJ7Vi+Y
UcIH5z1rPthXPH+IJKTK85sqpfPyJrS0MAQEHmBv0jwl2G3VMQ8g0oBSIyEGBQENv2XQoR/aJ29a
OWCC5JCPGmmjdYIelaLKANntQZHdyq3HJ93oCu52gaQ7pfE0FvY3c6WeXx6sGdpNe+xYZ2wSc9qH
m0niXEv6d7F+fbM0uIwoQm6NkcmCVIupJfNLgtSCO+JgxI6TJj9TxLXat40eatKPzrkx+eNR5MVQ
OkP48Zv8bID27G9t5UhFGcXqiiF/nj5yHwZd/AruVkQYCvFKvZXn4zKJRiWmp+S1TuDvagFE76Hc
z7EtRqNvwcUQcreXWyxyn2ur4EoLQ+hJ8lSzrYp3FVdr22Vvkzk9f2cumuX346Kwi8+/3hqHSGEc
HjdDNNj+YKEvxZA0PSBwlqljD1FZwGybi9yrfLysVmzblBXb3SzLzDNMaPeSojJBCGBDTjqLjfSA
l5o5lL0f0qWxYkdTgVwJq8JphS4mIKyBK0ZPpcGE3lwUIbskK5o08d+o6Rpg5mylyJfLE6zWo96j
VJnFjHN7CAseQclmBGmMd6cd/YQQJasa81lF4bd4JyP2W72MFJD+/4inRlL3+wm8rt2YG+QumA2B
fBtwByYNI+rq/86Atzte2uCDs2zgod5ZrsqN+PDl/aHvBw0O/OWwvcMT7nkTOphQmm1sRIregsXR
e/fvFu/uVZ0WT7SzIdHW48YQF9IyiGkQOP/wvw0pA8ofUbd/s0yoUpHIFAqIF4yiDSKgTjOJVGnM
1ZS15a/Qmw/mBE39Jh7eo2DAibaRtscDpRIZfqHOnRquZZ5q8pTLGA1RC6FyNSzdSHoRKYODS0j2
c//QQDmY8kTLCocU5nxjKUf5RhxFMzx42GRzDKji0h2ILD2lmDEnWmaO5IauGdf/74CDjV5aHCiN
xft/oGQhQOvBldH4hFbgXrUjZUP8wRbhG9k0J3chZ74/vnyS9+zDt1Jr4yIWf8eF02E8odZZu3a3
ivUOuZvNVrGyltXcNEGJ9Unxsx4BlQK+dsNXAZnL7gpeqT2YtlEctmaJVbHZhszkgMBX70tkzgce
ccsQUOr5KUs+dX9lg/+n+Gc6ULCdcXuyE0Xitg6EVF5ompeLfmWOveiX+GJQCRK/lRgMn8fqNrYi
BFCTQRlAxOekGns/2z4m8kmc8OuEji4OSRaW1ANXDojSCPAkNalf5xhiw/Je+wAKd3DfHMJYgM2V
1DTfFL633bg2pBjZ/xhZliy6gTEAiNguOaGfPtze18I8yfLMB9G4+fRqaF82oBdEEYy2AUizkP5m
uuof6jJU5P7ZMfnd76oyza8+2G++7luy//JsPOQtTB+60uj1mUCMlSYg6Cc9vooOi1zXPWLi+XFR
FehdrxxrpOSI2+J1zzDrj+B/Ugp2KqTnx2CxFA5acEoTtCdjitRVqG2VJZWJ9Xvsj1WFyVS58Sn9
LBijluV6tSOTreFbAUrU6EXdHyb6ajt3U3UPxdnliJk5QXD1Mdw3uNy7uCQK6X4AjIk+g0N4XN1x
lvRIEMinZa4CCKhCXyE+1+7zuw4xZDeyelsbNRdYpN4INMk40m3uZGAU4FXMw1pxVSHmTcwyE7Me
Oym2CyzWlbgB2SadhIDkOCAD1hZY00/I/qpHu7ptefFTJHpWk1lfgLAEeHFKLAXHXSJ7w989pfWs
b8mubR5yexwo1x9o/oE4gpCzQ4jftdbyFHfCTd1qKJ1t4oLnZZyidLRfgBPPBahlQDM6qkveE2Gg
fPcg4uj3wgKyRdvGxHMAy7x8dc5R0IWh1fOiUACd1Wz0izPilkLj2IX3oQ0Vdt6QC321O1ulQYQT
8sKGyNQ7RxCkfd5GrUX7tiNUpWxdB3Fm/UR2jdInPR8Aazj3zkPFbLh9inGSOHNk+mDRdyU8Hahy
iBm/NeEQdxLcrbLjvF7K49eodySAOl2XA4sP8qA8aKV0dzzGkMus73JQ7SqcmqOkRDD0ECC6ZgCb
iNRmNiZU+Pclc5GIDFxVk50rJR/TxWJTiDMt4k5MDHfJC07egX4r7u5OPjEQNId/5koxyx1aZuhX
QaV3b88XmT/E7HCi6jaBGe6xv46jg/u1uAfq6z89D9DBDhAhXC+TuTGDwikpL4jzbaUXe0rtLS/A
ghpna8wIrHjQUFEW9w3CwqLe9bBOZ8FTGLpnF9UnMBZnmhVAGA5dN56yjziEL3ER7pct4QQNccuk
67XBfFXx89J+NZhm+ZCjYhuH1vEHHIUUsyV6SmG/MFo2JzmXx/z3hTT1QOEyApTsosdjs3go8q+W
v82X75+9AzSC/cpFUZVbEEvFJV0y6070kZ791aQSkKcf/GG70Jvl3unv/I/0RHy7ULffFzlfrB4V
rG7tjZxsmYKK8tOZnkmx6kOAAG/hRgHsF3n7vLmPKgXQDQv/3vK8LuNr4hwX21KlLXLYtouAssev
FJDHWPmHK8DyC/TZSStYTv7R862M9YkZSxD+0azqV9JqpL4OjTpUix4GCsAV0422UYtb+FJuYBW1
OqzuGdJymbZJIfpahyrQDtORbimPSPDZc21gcAHoSizgxzCk9NKfXF/1rajh2FBWYt3s1Glf7FZt
fUAq8ezH4k3X/9UJD551Fb8XvLWj5q0P1EphULfaCNIxTyDa/1vJIfqjgdRnvTBfz1kBuSh4aYGL
0m5Eb/sswW7ulkBJ4HFceNvhjwfxBQFoEUdRPLYSovIfjtH6g/BQM8WVWs/6QMIEqXjIIiaWw1cz
A0tqCU2h848qF5F6gQ3PqX0ycnuKG6N/c5uDByZrrgxfQ5EbDdv/lb1PrDHV1Y+U0zcfdBtJ+iuq
5Ob0z9uIarBYi31RDOaIEI6+txO1wQuEz+G4OXplnta4GiOVwvK7+lGaXitkHo8usn4pIzax5j71
OJc8UfIK0WPdGOCEVXmylH7c+VaeCGMjehEQI+u/52mjuZ/TUlRZvDeKa69bvbEQjyIWhD3q/y8h
4Mh9MfDhsLMqPpmAjKicQCbYVVQKUpFEYyuOyUmi7LvdeJEGnqKRlltlzBfx/uz4Kl4O+ZmBE9mY
2iuMInQSpi3KHRQrfarzDq8K9p0/z8VTbXVjrNdrVBKRkGU/TeuaXRWxpU266nj7BpHtc9uNQgzx
0i+AA4alUp1c1H62ixuyLTVYR6VVD0DFNHFLCbFTtq/3BhvIWF8g0PziFtv7d2XuoLspSojxL7TF
6G93EJVBNdFsIVi/HdMtvxUvEbWhBFMZdro2dheVIAU4NuIWxhgcPLsCzUM8GvvZQVyB6HemfDri
3hMObpJvShGajv6g38Mo2lwDdh4amZwG1+g/3l+XBfDy4Vq/sGtmQ0Pl008/ZNhvws20nA1OqeTU
hLjnPyT7LTM0/hlC2s9QL3/70WrLzQI8z8YCtoN6kxVw9SV7uxRYGSxyfE7LomP/dWR4uB9gHF9L
nbgrWxHHIubD75yr6dXjSc0GZjfkRNVqyigYzqMPe2dWbL+cVwhAqqVyvoufumaHGKFFiLkZm+0C
d7O6c/7qYcjjKRxPclmRlZAaffUHqwXTKu/bMAGOT6yZ5GHdOEUlI0QqM4jmnR6u+Kb92yvP4PgY
spc83PqhKaerHCaikbkhX1UnBKPF7dLQ5RNKLjfUGCd0zG1yJlGBcsRcA3x22/D9KW+ki5LfP1io
hQiadPZmrQIXFJGZtjuzTpCMn8UcWqhfkqLWPa8JkuXMtxCTe3jTQMBLxaX5SATeoE3BhqyHhlVC
QLHE/x/tfz2hw5LxC10Bf1HzsYM5jlYjCQrxVSmRBC7sJHzmD2KD6df20UTXsu17arePbChfcBt1
E6Qu48vCUdYEnCntoWyzXwLeL8A1JYzUI6Z3JaKy5i8o+eT28S/hKHaxb5T6yjFs7KHjjwpIXq1X
64J5YicMi+ntIUDOl4ATcop1qWoev5eNo1djAUeN/yvjC4WmXPvt/v/BWGzxz/BdErjJkZYNhe6H
ZVWUA+NFxkQN92KLmH84mxM800mGplGJzet6wunAMy3n4Sj8Vl7jW8UN/tzT2RAiVeepfwn7zca1
NlNBqgY/NSsdTVZpK7Flmpct6Zdd2dU+rZpShMnjbq2VjKe93gmIqd1GCsL4URH8vHa8FO+xogJD
TrU3S8pCcwvF0EFGHnPRRLEQj9Jf2SxEOfKsv/laCLzVMRZKpxOW9xfx1oh4mFOfxuq/duIAWklN
T46wJPBoaBrsHXY9piI/uvgD/sLA4mDzZgRbdKfcFQdXZWZHRaesgTJNuDAw+R8jMpFpfRlx3Lgf
qbGn8iYACaFDMtqsBQ+XYJjeNu64Bi6l2gMJ9Ma9VljjgAqmYGmCaFcVRwd55cqyYepSANYlQ3pS
6yt+b/9s5HVtGXiJMpOtqakp+TusNLrOMInD4hM82P4uZl+DOhyyeR3kqv0rmDldISmWlCqJ4jQ2
U3wmF5UGiVN6Xp05eiSsEDFgCNT03mj8+SScPuOk84LS0wqUvPq4/LI1YCHYWLl4l4MxrunRcJkC
r9sDTcexm2b9FpdZ0sWzEyGWrn1jY6H1JaB8OMF0V+1aglFPH814hc8o+n+f9MMWFkgSwyZlRw4x
bip4dXT3SfMS2LCIBtIyHxPM3ei9Q8GUru9OKx02eS3SP9q6f2rG6KW+tPRzbb/ZybgrTQAzcM2G
ktDdLUFtOzw10X/VK9EaSls9sJi9m6Alywwcr2EeMFrwsn6ObGO6jxydqqfz1srwyXUsbPU/lWlU
SPxOevcIY0SUX/Jnx48rWFyi+oCBMHY0izJfo+pbbbA9MSsTaQooZZMuTLQWCSogmbiDiEsSdKzX
3CmK8gNvqoQN67d5flYzH+AkqcX1E/QsMIygQoSsDyAEVluqywRFui/4QHrbG9DzO10LqDfgVnfO
NUS65txNvSfp3XIjms//jHGhql7EQBhYSyBppwfmvcf9LoMZNLXL6vH/CVHuAWLeyT9LkrlH6IaB
7fJbqg0QqEKsP7Bc/0+QP6kE3/V48EtPLQWllwf/3PCJ5wTSqPNKKnDtiItrqdmtSYPVzJZ7gQsT
S3BU9V3oESis3duwUFiMNcD6PB1raYPfiwTWroGsQk2o7wPffkmlQu2Y0uhsoO8Rul1T4cUx4DTY
zSvG00KUucitkzvCLegPEL8OBTa8nSvNikVGurfRWQW4BCLhY5uH0kzEVfX2ZmJraenS1POno4o/
95MuT/I56tCXvIJr0rqkvSN9ptnUUsCy2o2IKGzrCoP/fO+aqgV71yDDRjhe/kC62zqbx1BKClPF
7jn576yfFFvLk7xQI6xdC7SZRIJC5vMJkk1+QHO5w1YzH7R2Yi4At8Gj3LZPlsqICqlWfgbo8fSm
H0paRTK7LDjPFQ1bUz//lyJT7J0XGI9MYRSNYrYqveanOzbrOmr45HuusTe+OiEk3IcROsg6sOXm
ziOhiyTyVUIXaRjDzFPwLDAkh+KhfJw2RWB6wNTRp9xTsAKFJ86LPvA01wm+A1O6WQGVKII83+Po
PTuyClkLWY8C6OrAb6Yuuu3z4Ea9mZUvr/K3yuEyPtzu220bxW6O79Z7c1U4poyhPqvfwlGFSjeV
CIv821iV7crBPuwG4NfBUKFAtAcQNjKLvMC0bKDoXrGkpcPMlADpIkxz8IMAqIA9Tbf6R+g9R7dC
UzwqQiwuDTzBWCyL6kKXP5HulfhPP8MEyBL93neA2oby01JXllhxJUwn5EnMdaKcGiDO48coXkYl
MFTd/Dn6y8UWNSACskUpPnlQoa2F5T+ahROyq7oJpp4er+vx4yDxevNKHP2aBdK8iPI2V8IyzHOk
vr7JmDw/FqBKpeNdB8WXG6xO6q+CEarv66cwpbHAdDicSiRqqaVnNq0hSQlgzfWtB3HysZ4PDf04
pzonpyRK/V7qmgQMS5/vyrTp3LMMNGwaw4mMoVekLO91nj0Ou4Rcvo7BTKTvXP8FGyvYXhXxiZ3m
5ALqiXM10XFDdat9a0HDjjfW4iKTKytYEd7tNVIc+igrdFAYet0wIokJKEgF9utqRirakhqywg/Q
wjPRWu0UTN2mdrVzVfjuOWm/PAdiVDUtGBZ+TvZFMUMFXMRYjisdRV8AtwQkKEPfEbDYTXx5qt00
I6OYhPueAiY5GAgQTjWNtGdCRZ/+Msvx6lN2f+qm6mVVHvl0EcBIBP6K4uPvevjvxwaERyKUuDCY
JEuz25t0i6krWP1OrIhI8abYzSAaL83rJPJFCIoDoY04I6esWsIebg74rL4EjiI366KGHHfgh4js
8DY5Bt6WKPUoFrjI2D6y/DPsybcExUO2Mp5avaPWcWw87vtE492wznx3E4mzZcL1XZk4ZvIlpHo0
qQPIRydKWJgIQpEsY+EtnTmrfYrn6WuAi8j8C2G6hU/D2B3wkZqbhla0C59YXEVirC6UKVh1XSV0
CU6TaxCszagWRyw8BnV8sDXKFlyii1KdILvYutu+N8EaTESyILZsFqDJ9EjV8XZdygfvkAj2P+wY
NKh8DrNQDbAwxFJqNPRagl5HCdVYCAwUWOzdgDf6NkrCsimVuICHnkrrywZcQvQ9op+uAEln6/UG
UFSVZBSNQeZtEKVADKnY/yCwIKUgKwNpuJbgeO9RQXI662H1LQ0xEQqUBEk68IUI+8YK8rQAjtxf
Ho//alOOu96cbiFGSFwUK6dLKTQamh5b5WjFq4E7i1+TZ1E3+mJDJXUhkGKeBmdOBd4XpY8497Nn
MM4tphzrw/OOws1Jy6ub/+KZ7HDRVJlGzjX+aRXFtBT+2CCDYWhpMTmIb4WO//mg8BOdSOxbBvMn
7G/Jb8EHRFbRNylfxgrZOwVV1V3men/ofiYoVnuUnhNPPRmXQmGNsh5MGwxXg01gsMqPMtHf5F8/
DIot7Xtag8JgG6ItNHPMNv1/X6baf7eGuJ/5xxoaAnelYd2KVfIu6EOLwJmRY8MK18rxFxtp/IoM
IRVwv9GkBMiDkIFQKh1oKYzQNG8mqYvfdktF74dQKoyzU4OsDrtvmPgrPidsNCOc/zPzI5jZLIHp
PavN18T0a1KQtwZsB8pwxPLwg1FhWjnE+uurzgSCFCEy0x8rwdaqaZDAClvfuB+fXJ+QTOoEOOpD
qjsi/MLn7WaVH1YkBxOCgPaT+ZDiwEPp9gkK9cf9TEmEHaO+kDz8DjO9Wp9XB1e6mZjKvW90h3kL
U11rwEssAjjQEhkvivieoGtk8sr3WtpMQdPEhE5BWs6pmkBBqN7tGsXh9nPNC1/qukIW0sIbZTKq
PTiL+y2XfeIwUgqg7QDH+ti5k6fDPG2w8mSdDBfX8i3TcrxMqE4fJI2/CNkDj+isNbtod5136Ky0
G4BOCy1KSKIOcyRJk2KaGBsxQLrTBHyPLsj5GTfd+J2v6s1e2jgiM7mQn2cGimgJGRAJOozAvK5i
YIDpWIOCF5JIjF+YzyPU/btggzeSaBpI1YGgsWayvHh8/B5kVgQXVXhOr+7EXxVoLU0D0PM1saN7
SxT7f3Vs6t6SAQsZwtEW2lRkIlmBNSMGrxEyWdzH1MzlFUV+y8vg9mDL/bIeTSqpE0PaicqN0O4x
7R9sSRfLBfWZFHHwOofRd8Mah4QHBKEEnEJLe2eGCfWSVWiZbtDrJamq8OSOMnRNAt1DyWAgQza0
VMGAjj5o42Xzt+uI6FchOVZTLHEbvpE81FFadJIsjrtsQbr4TRxeTgL+s5gZKRd6X24lJhrXWbam
acCR2FbMJhpWA2OaXBzSon+TUkL30o0w5wIoLseSPaFapsbWbFTAMV7+8XViJ4Os9FktGIt7Yk5f
bOubDjPsu0iOg1+EAio9ed4XZxupMZzl96S5TsR+xPMJlf5uxbnMGr26mxkpXrGB6F9tOPyYZQfi
TfZ7ZZsrvGh7idneqq6paWnnaLsrz7WceaJKTr+kCdLrpsOwWUgs/tJyu8NMAV7ZZcleKVoMbvQZ
rlTBfxqOkUIhKiXJihIZwCe0s/f6fqZ1Otzp+nKYAZHPw6Wu0QPibanTVPmgC3dhRnM25c+aikFk
JrttKQ08X/VGs6FKbC1yHAXqLWjFM7CKNldQkB9NoBYCN9HsttE3DTyaRENHtKrAjpQGEE9zT0xu
RSKNxd6kA9+k1Cl93aBEFnG9FkAwTVOmsquCaxZrvr4IQyxz2vMPD0ivOuABQGVRNnji/D1mK2YD
OUC+8LZweH/7GSwyHf7xH5KmetHcd6XfAT60bj2pJZC5XLsVMvIA5GS2auxjg3wSOEA/e1iFbRnV
Igj7Wwp5AjHkUTbhP/8Ck+Hs7cBoqsCjElf32rA7bxzhrSyHFUxu6KEoH9scSDMSaXoh/W/yT9dp
h5BEM4dyUnOmJWdsIebCHXf41H5JOP4gc25z03Sxx74w+vN3tbWqAQzhJmU4mP4QD3q/htk3SSPq
4z1VuND/u6Fr582DH62VD261wpmtOqf0CgFGHxZUPEH5ig6EYT5dK7BRrpPPQtr4gEJM/PhOfANB
XwKlW8FK9QtnEj/Z0cqYpDo6MxxtP+6cRRsarjuMrjUIi9wpRuXxdkLhly0ktHgGqqNLw7q2KXL1
gqFMdAthnLpz1HfuR/00KQuw1qDW0rPXnN+F218r1e0QzLXA7FS8WEStWm3sgh3QDaLXyyX4mPXy
ocEmMFQnTaZfbEimLNcsFodoI6zz/xhI5jaO4RkVztLFsFe2reLKjxOzsyKN+k3R3zSPyi7H1KS8
RMLIULa7MMjQLm2wdK93NlGQYrmVyFbN07AbDRzadjqJWJ9gNMJphXK3A14RIUk8GAKtajZOeswS
5GtYd1R80pO6i36sh3mJzg5t6cwalkOyVibwXs6vPDlsrXHKdizzAwUa8n4u689Oc342Z8N3a2of
4xwVR/qMaMHEUzqojMnsR5RoZXZkArDqDI2qMQDAyeof7+iWnwBc+OOxiaBNgkV/HSQcI4mfms66
xbuJtL1yuioUymTpeTzaRtNe18M8JxwKKuAZyPMcCgXiLi5QGQ+C5Z35+J8Btjmm+P5qektfwPb6
2HtjttRFl0SJ9jds1DHEQ1VPozPYYmDkLk6JFRuEjBz3Z1PLN+yNt/MMNfzDfO5anTLobXeC5wUX
OJlRaSU9QiigwwX1yNU4xzmircFWYCl1kFpu3Nh62hCTYc8WgveTzWwxieL67ACclmvusT+HwRtW
nbwuALK+j60dRD/8ZJn2t8YHk2jSfxAOd6ldUzWv3ipKh7xKH4sRLyk90/yhLVIHMCZ67kAd8AND
EIuIQCvstO8w1IEGDTmQ/KIdnASRX+8UnE2xmgzaekxKKZMdfVXkTv9CT7Wk+qdpRkYZ+HI8LAsH
FTpeEgJR6IJfSAy0ZI73PIZNqYWjk2H6iwqwp7y83pwtozZj8PHDebTubWW3wdZAi8Ck8xBy+EZo
58MsMItYxaoUylD9gaXTzUTSkGI8LloRBJIKjAvCPAHdqI0gv9h/g3HYxyWS8FEhQxKDSBSwnx8e
QfNKNq94WOWkXjbxzl7wvPzzdPHC9H+4d3bJU+lpUmf61cfUWhkkxSLIZA7kb5MDaSWyQ7ZLfgvU
kLzx7xyjzX6RabhqkeurSA11XPyiGXs4YQc3BCAwjBBPEpZticXXB7FQPH3SeurPARsn9J26+mao
VG3Z3canWJS/FlXyi7zpXq5ekHMnDZogP58q2O49Pv1u9qgS19KNDOXtaapHm04CSJZyKwS1bdw7
gHy4WY8yFmOAbUk0+li1a/HConz8YAFRS/FV1XO0LXy0Bhio2x3GP7pIA2lku2PvwlcpvfyT7B/f
i8MMY37cd/ymbeymuZud5OW7soI+UctX4TULnR8lpgA5YA0cR4GfSgzFKUirqP69/lyItNVxzOc8
a9bLPKEU9aDVOa8zPj554nhClYylyqtEpMZKnKg2tNRN7mo4+dPXORRpALEWQE6Gvy/fbJoVYLwh
kLbvn69aqxgj5OjzC8NBPxuzB0xhfMl1ZPujiDeF8Is/i2rTB9e5Tr+xAvGHSr9tDraE1H5Gk9fq
iTd9JDmLHqnYArz+Ga6NiRSpeH/lRVDMbG7tTnR8z/6ScyqlZYqmVsX8ctLMvEwpszjqmDmZQTd9
T3kpgRT7ZnE4YsxY5Ur2HGOAye/oY9qGBYSi3yKT8g7lJ6lmUnnb/CbNDRco8Lwn6/nQ0voNBhgF
fllzpFXR2WtEIQQv87YbWiuVZgp/iXBXbB3imXuUbsiSSElzlm9YV7wT2vfHK/qNl+lnBwCcTIpe
TM8dC8lPE19OFxFzWZAF6lXt+DfETeDuC/98HPe03pUC+T73NmTHORVOrlGoYSCZhAx2+OG3FQM8
iBLH7qYh9hnlSHQxGvYcM2/kI/YT1pUZ71Q3LVTTG9/1UOe9eyT31hCMcjDwbpn76f5RtHl0V+/u
dzoG28HVYraKOp0ucJwx1x3zAm5KWXHGRnZvtASx7GdmDwMJ5yE0Rv9yv20Y797VafrdLWd8DELm
wHP1GSnLIbHG//rk0VK7A7PG80oYNc+jfeWe1GIVE/BNfCNrBQCiCzaEEJLUQBYBB2gYUMANqBsa
MglEa3waLgQrvL8z+uGUIltoPl+yGOA3XO0Na4/eiCvDgED0M2sYtPOdpL/LuOctWy+6On48Ks1A
P2NL7Lw3ziqpt1wppJo2mY6FIc9ec3d/1evCi7qkNM9eb7Vz9GUJDOQtT7RS+wBu/0QshvpDi7mX
DYsItT2dhqkeim/qnAdYhxU9OPUX+2Y9QXCOZ45jvZ2Sfa3spyo2ljeAqsfSPHGl5pQqXGz6DSI6
yG8o2arF4h7kMFMUJp9WZ2BKCooua+z4+ZNfiV+cloj6dmeKektmBiGJkwALPJ6m+2ECJXwlT97s
+5tOhkh0dV/Ltzuhbx19nJM86BH7AYSrb5g1jrWVmMWprzAZ3Y9Fa+ZcFJUuzT/5XbL4WwWlOnb2
hpw7bw0kiQNNGZsXx2bhYiUbed7zWxQWveKXvl0O7br1wO2BF6nefq6M5zQkFY4c9sMS8ahDkX9l
1AM4hwVjcdreCow+SpEBOIosZNhs33u8Gdj02qRPElZqyFtR4GpvxyL2rUYcd0RcJbvk8b2uzd2t
TNtmrD8TDbLpasysIumjwQUiHg9z98XpofwHuCXs43JEUQ1+hXbwZFYO22w3Fbuvwp1TkAktZYmi
896AxusQI+0D5J5y+lVEfCcLghrg80cLEw5rlu0Rk5v9DNMGMPZLd6CGcZplPqvXPWBAfaGr+vPS
2MF/1HX6XAbeGX4iN9W/r0q1A1gBTu9Ult7lIldPem1jHxXOQqYgPddo0e1eQBVrAiNBKpxZpZ4D
XJVDbvg8xLYi82gCU9ucEKbzOwR3zSUXX3RTkVTl4Bt6oZMVsDsP81UbCnbdV8FgK3/5RONfViHM
p6mQj7GqVLmCMTHew7C0lEs9fENt5N4hsL9eMet3Ec9w6rhwJtmCuZcll8poMyfc8dJprBNjiV/u
Y+jVMQ4Gsfirgio2wtX8mlkPySQpfsZHeVNr4wFnu1FOTTBaozuRx6ALPEYDcZWLc+NKnG7j3LCJ
lDWKp8QOuxR0KHpfQ37mtlo4YRlNFX5wEUnbwDVS28ayCcZp0A9m/EIJObpNdGZucIz/Z24DLPs/
7+lMzvdkIsTepkbc+PAkqjFhebB2qgQymkc0hKUkRJBf9f8NqpET7SQ8PWoahzbc2TRRAkbDIRfk
GIH883cHb8wm0+g59qZve/SDaFJ78EsBjdJhnD2U7fScoOOf4J+k8ozYabo3RMMvn6cNJMobLRzg
uP3R9hXgqEWuvEJUNqO+oGe97GX3OdPNIhTEvSPdBHrZ/TRZ2tk1mn9qAddUW2BnLBQQGVEbexxV
JwLN1Xgf/eWlC7WcQNO3br5Cf/DHDGUwoMfYt+4iPcxruHQur3Mge2RZ91B3yI2u6rDLK8BbgWuQ
xxsFqlkwR7YkehA9U0dsx6xCYw9K3Sq2eD7mFO87lU+QaqODTYfV/7Wv99XxZz1bW8uv2N2EOOM5
aQfxY2rX7/wdDK8B76zKwWpboKJui3r9632YQ96u6vjKYKGJxenbSrtPHsfuSoxJIPteRC6j0+PQ
H38c+HIbpx6ZfjLV1ZWHDz0ZEUjoXrnSX7fvRBS0cU0Fp969ufDbc7MBDrKAvXckp+Z6Wo4BZ+XP
mN1y6lyt4Dd1NkY1OS/210jz1E5BdEhh/zQkx7LHqYW85M7nxw03uJJRIBi0cVQRbPlg9Wp7DLiU
J8//7i5rcCneECG2Dzl1CKnPFelSvMPuqYkpMyI41Xc4yM7vsOsI0r4KCXCJk4/LKwboZRPL04eg
3dsp5PnHNpaXhYUWQIuudRPA+6HWe5MsKxFeRkpKOL5KS4AukIkwEg131EB6q17nTPuNQSPTqJfC
L2cl4QNTVR6GOt9JbBQDlRCWxsV6S5zIBkN8xuZbpqVu0qZX1D1/8/J+E3kAO9HEPxTWooOLV4u+
5K74uwtk0WA6F6QlBhQw9c90c+rLO4/79kBsW0NyLG/OuDLQyaqKki9GsV5X/dK4GeyWOBbDVRtz
0QQHOcLalY0VHv863Xrfq8yqdrG/+59hqoHdEjufMbryWOBzBlmII2mQTl5vOnbJsrNTYU5qn9/i
DgQbB4Li/amcjQaqaCvvML+VbKCbiYlLVYlJsG5tdm751toRmcctjFrpRdBg+vBDgwxaf/aN96Gq
M7guRs16LHAOION2WWyyo5tFm//gQEXU/cXKOeWyDg06P2ykOzOco4adrrg5cm60J+INrx6BJcm1
AUZAnmXJnfPR1XxdodXzzFxDH/dg8LVBQsa78W9PrPpfUyuGFuvyiHaC7Zg0dq1KXqhORlhWPKov
fXsrxyWTtZGxfv0xJzp2DxeRD7/ZAjQF+Mqrwmt8BH4ZpKMUGtNjFAE70TicoDv9hgsZYNvn2Yo5
LX0mMs4a55ZfRydz27CoC4j/N8GDR6dG/TOnK6mD9+/2BRD/dMTVg2IyV/jeJ2m9LRSpcUUccj0Z
fX+hfCUB6UF78vNGW8yIagLLBS0iOFMfnBlNERYud8XxNAyfhBnkM8bkvs7mgpxOHmCzfSNJtLMa
zyZrKd+iGNCa40FcGIBg9KzkwggOR0ZVBTsG5d1r4UI2ZxaXm1jJhlAfFtNnzXe6QWAzlu79PW43
gxBpIDrahVZ83WVVo3k04GWYYhDihqSj2oVlEJVibAjAWRC6o4YJDZt1lxgNKSZb7Gy4YzOH1GJD
ma04kgcKThvg+oLykbUu45O4bsnyE+mdy9yRsD5bweez981/OlHXMUrjIrOP8NVts2NTsbTux1La
se/Ovfb/R94p0WGRVvWEaQ7KXL2ZX+j7n1YDszcsfJ2Sv0m0OM8WAIXnEX5n12ejhRVE5W2cg5sj
3L6ZCd5Yal3cj89KmR7+Lu5EuBOwOxR2GqNcdyS7O+1LMHbKD8o9nJFexo6wtbsbDQwNS3Bg14pU
/h1Nk4sS0VkH0+uGOeYeZNfEjY90aagpCMHU87N5ycx82t38sIq28NBtg8hA2fGK9KNzKCJkossj
0+Cga4+L6q6hThWF0AIXF5jcBZRwxt8EEtqVomODfJLx5t1DQ4MYxezAj80MF9TzyajGkQWzHoMs
BwcEdONO7wqqHnHLSRoK7gJvYr1Ud+5hyxs9WfamKVoPeGSf35CpI9K8smbqWY3FLiZOLSso2J+O
TbulG/ft8UZ9yoqEddz+AMv51+cwG4+R7epE/m9C4sUnbJjMHxXAyq66BYIjzbrK4sBAULCOl113
SJEPAgF1r4fAwNgGGpkOJY+WIvWF3P0fgKHfAHDUU3aZca87JPktOMUzEuZJ7ZEnXUiF3UE9ZGT3
3sxXChV0bbvftYs8G+J/WDcCnZzVNgvRVymXN8FgkUAeVlF2eihvRYh7ieTPmzerlXObI7YcMTqg
FP4GTehwIX+TMrDJ/NSJ/hFfjdSR+DTmfVPjYVyTN7juGKpJz/5RrjkqFRqwl/SwTBZvOHS7lJdJ
4njVzrZLA9caLPBF9wt8MjRPwg3RW9E4eIKpif19NDl3ubupcmeV2Y+3jMS8APjABpiuqwFG/xWY
e6ncglBkGXGM8MZ4enDy+mqgth4FBY/1m4fmbp93OvAQPTNvXqzP/0Op2Zx/aYZmKe31TH2Uqxdg
GYRweR5wJSnpQUX400EAay0JPTeI9YBEiZUqHhcVmSP1txsg5DA3pDq2Zzvx2OAgKeZMs89ne7fi
HaXDRzWOyFQeo3lS9BzrG94CAzJXCwxXUyZ0mK/oZCJ2wYSATFIPaE5X77Ie+te7zK7IrXtE01M2
nOIL4lz6e4ENnbOGkzvFXBosPh68r5q5BL/bm57sIcP4d4I/eDzqNWYscSvUv9FwYAz+wora9QG6
mtbe4yePpfwqXejO++lPXnYJDvhuZqOkh2Nq21Uf/E/coeHbL9AAy0/Tu1F10fi6XTLYqV1QFfnV
RwWzI3Nd3UNFmvjT3muZV8J5y/jp95gz5PrPmfJpBUYWrAUZE6Hdzqb2hZgQSIc1nTxWNOrGih/6
POOkoSUg+KTBqXd19Z55XBCKqhTTGxsHivW9o367uRo0oq/acSUFmlc/9ilslniluC7/hlbSBlsC
dq3QIomszElyyoe0UXlo3oNKjwVtjsFKVtUq/niU4VOpbYVqKJT8BTjrQ8oQxDYV5K0TAenZuhWa
/cyupdPu3hMnNKe0CJM1RhSLjtAlFy0Wgwq8fUNybz3W/1/tRH6S/uEXv2dvEyE/T6X7qgy5mTiP
dWj9g3Id7sbnMCHe06pSfZI+6tectYnYOKxgvGjieA4TDoUZl7qcUfYx2efIZ1n+Q0mjIvDdlwsr
cOQHkUWw6rtQYXwyG4cfAKttT+GooDJVIfWE75XkqlGRV9F7xqfy/S2LJp0ZHFzLUQQc1c2IB/Yd
Woe1NhgMMJXSGG+fJio41tknAZjPOElLgzBrk3ubzX6/UGNRG0L5pOqN92KnnaksLMwNHYGevL5O
Ha0AlfnpVwyCKAzfDtYLu9HlW4n+8VYS/lOAKBvlBx3llkVBhYQMJEEdYWuZwDVPVhQc8OU030r+
24TKAienj0EZtCH+UjWMF1B7n40dgW7BmFDayha+LCbs5+ggeSU8XvLlKdta2r0rl5q2RoCllb1y
5gXvtKnQJ8Y73ujCbS5gm5m6KeTmI3W79FvjjHsT3tW8fGI1ekxxnBOpAXJJZ8d9XyoMva7Gy8fr
sNRzx4+KPlafZ1lXH8wp5XQDn4B5kWP9iClj404HWF9oFmzHjFth2Mc4o7rwaTm4jz/kK0D9Zc78
cRb8qYIHXAoYVdIKlkNAbssLs4xLySdJ9ezSzBFTZlFmZY4yZ0Yd/L2449yXoshKqexgNxAiE2ex
8N8o+1wBhbfUbNAxrPFBEO4NuzS5V8N774MS+s2VgRHKqGDy6B1mBtVgVT6T7XPsKc9UhiOVdnnI
U/3CsVCRL2s2pY0qvx7Ldj3ADkS+5c4QMEd64a7v8xfchYw48c89gWNM+S0C0cD0aMjdE0KAaT6J
cgUVBWwqt13TMp3keRifW17kLMjbaYA222xUsyxgWnaF201MFUHZP8h1vZ/E5Ch05yW+EpD9N6ik
TSYZvTW5WdZ8fAZDsS9Ul8gkCT3Y5mVZQ4KABCb6deOu8AgjcjQHjAbPfM0C1neq6cwOBm2bgvoP
B+r6eVWeUHniiT/018avzsFl6gRpGL8LOsB2CkTb5NDsXZ+k+DWHOPeFwmxlOxJpVrv5pkX6SMuN
0jOQeTObXwxfDK1MtOk8BW1YkBjneoh5BzN/LWwiGRySeoFEtpp6BjFY7YTwvabS/hobFF1eGzB2
6q9ezirWNBJbqTOMWet/NqQApeWqwZbOdlj4XGFd7+Qyh94GpN1BoHa5Q3bDQJ3BP/61qEUFGvCW
YYmWuA2fxm7Cja7qj/L4mpdNex+WGfo4u9hMKbOJGgoa+LtOC8SIM2+cU6444gd2GumePuQD4BsI
JqsuVKbFPsSPeEIYWInFqY97cQODiAdDnflFAWmert5k9TPR3GPaEa42A5zLHv5K+Nq4/z1MCROc
KKhTqo8x9fAfUk6+YuihjGRIBocNvuBXjM/3XeLhjtDL8YXsQqVTg26eFlo6Y7TEAd4z0/WdI9kl
GPe+6fcXNs5hQtaEHOQSGdPbF3k7uNzYQ7D2i6yaYHgSEISKIrA9v1WRfe/Ofok2+rIdD+xASGIL
ZD2JRWnYZolYmA6wEeAwqFYdbsSULxUXHnBU4L7W8pQUW+QoTYLlov/RXKRiks2iTNd7Ygr0yMlx
zM0tWRHi0vr8MLPcZi1goEQcKNGZpycnc6SpGTgd20+1AZBYSjqs2kTRUvDYHjX5PNdE7IE8FUM0
OuZnMmYvoLZwWb1BXl/C6S9yeJf8Y2ZN2h2qBis62Lg/dvyCs/DqCaQysaEvd4PRRTumjar0uWxZ
MbWRFyUAyq2akqhdsq+ppGETDLN+MSQXtx9HAPwh6ZJlXpj1enD+aEEywxgAams/whr7KDgVZXlU
wZtoyyBIKt3VBVzaVaRAqkOOfhZF1iAUMeGPWxMaOI+MsX0BBLZDIap95F22gnb9Tnm3cllDzTrn
Hi0aq2GEPrghDg+tLrga58gEw5sbxREeBFibcVnpiQ+K0FkKYg8iJ6vy4iSuD79Yk071tO/n4KTp
itBJUZQQoBaP4EIv+UiRlsM/9K9p77YlcGAYWFXHpWHX9sCavIqbC6ZUoBmDU7T3hJEq1MCbMbtx
vpbpMJS4SUcYwLwCkJp7oXNA5brddSN0lF58oEGnG+iO7ij0H0D3tqDJe963P8BUMhf2o0A9L6eU
bp7cC7QKYIMAOIpkvZqAD3fVUXWZRONZP2xWTuRs/Qqw4Zbz1S8CG8sW5bbeYkmnVItUBIvDscf/
FHv4VoJsy3dbq6EvJZPyX5wNAmSTSGU4gTSf1NopOLiua//AT7KT0x2PEfcilouG3uHcqcSv6eG1
vSG/AmLPM3Tz1xbD1vZCUecFYmzSpwlNAXhNe9ynM96PRfe3SQysyWxJilXZTGFjg2CMIpMyuu7y
3CEtrbMY/upRMGJGBCYwQ7r0B+WzS+nbg+5DiUd9FEP32A3XSBfo7ADv8dZcwejHRQBk1EECFVvf
uRTEwkWN0redB5Lz6zXmBQ4FPMw6wDmONorOZwRiubn4IghfjkCdRitt4epFpmPCWWrGY5u+RczI
Nhsmbf+tmTKHpCsQEeGOOfjIwWTrJIzBNLn6bru8A7L3va1z72gqSeiGaW03QE3IWYGaF13RbzZv
X3vRkwRnCeUP4DvIS7oOOHYHsgPwQ5g3sB1Cyw/mBXRekijvhGWlotXjqsfPrCPzWeVs6NOaAD5L
z2dAuo/6HtndTAHnCJUYb+qDsJabeIs3OO3Jrk8CdTvS2RkxrR9uziry0ME9gXr1tC/a2nMfGUKv
0OPgoG4a4ygTPmBVBZs8UQyIKbz1/SXaEKQGtZt4jNAngpIwZvBxIMDagVulieUiTe9+f0UEgs5P
uf97GnJKkJSwR/IRzgv1cEzpBy7t8kU0ML/07LG0v0dFpx568tZVMfRAMhov+O673sGSiZUetulu
25BXlRBquZ8ZEVUObD/lL39EDYlyihwtEkSwaJQK0SzB+yLKtCQOEQW+ilstTOkuez/mXJzszO7b
jbw+zwhWZ8t9AVWj76gfAt1osxVe4nqdgU910fVbq9gJd4bXAMoBjkklgePKhFLNOVP2iuchyzCZ
FwwnBBDVjstlMSrjNcfxWDYKN0Unsaw8pG0YfiIMstlRY7frK9aC0tVA4AtaYsH7dinILbAjnwWe
tfs3TdCZJgh5u+c1zSffbP9bpTpxk2IVqz6qgnjzuazmZ67woyizHkoEoi0it7LpkKkMmBxHFDFN
muvmQcX48RTmxz3uGYBbPpEquxiGnaDzU3kQUTDcyeuHx63NhYwbt1YLeLPIky2JbB+IgblY6sti
7C29S+/aiCHX/xroWoc2RzERxZKheTOYx3PXxD4tqNcj86JMKQKo7Qj7JNvPrTali7HItmc5VKv8
e3ZURJtK33/VL/h8+Pec8nlB/pLwuvupAeWuJCHs11EdtTboh7HDYY0+xjaoOudADsEdo0njDC53
exzewRmSEb+AnNxilMeKGvnfie62vz2o/XgUIhkX/LsLCXJltZbg9tNl808cBAg7TGv7nJRS5TrN
x22++XuW6EMjdTa9hiD8MspfB4XrbmBQ0XQ82LhRNiAFONo4KrLIPwp7a46iQJ1XSIMzE7sXFVDG
fNYikXVhbk5fbi2exWIAKEbmenuUOp4kvQd/NK0baobo4tk/nuAb1pQtymopeRYcRRhKqgAFyEVH
UTtJGkflIiwgNrqs5alnQFcYQwRx/6+hQH6G7Y+CzHD8mcoHsvEZfBnob1P/lrgJje26wCrLRcvQ
ihXszPl/cvCUVOIIIKZZUg0Z9Msfxm1mDdWUUPqh8mvCIWQMFO4S7X7+ETKfmKPoUdvg5y6XZ0ev
rw1iRTuVnhfr+YCDZY8kfDRFJUqXL9gfxyEbjFhdqle5n5xhLbXkdkYY8j+vcRDZtjb/hKSBXJG/
L90pcNobBpGZE1CuTQ3IUXQF7SdsCTNS993SbjBZuOni0a1k8tsN9X6OFPK3RRyMgZg8YZ9FBpKW
Fw1AYivKoV5ZuX8g/yMNwPKomvXNQC5IjeH000oq08C9UwIMTbUnO93kV6G2SBlsZZhnQIDgF6cM
waMprTXbfd67HtrsbEVS2N8MZizEwCOpE2FbNzNntRzzmwQxOb0qAFwecOMXZ/HHHA7PA77yKCuN
A4pBV1fTJqvqMzUbLeU41UrLMXmjoB6supgbF/rK+yhi/hCFY3fF54qvrzJ+F2hedRnIvG6X50D2
G/BGpNdsTr0O3XCdy3asvzKAYR4svy4D1G8t0x39GmA5xbNLHfDWaxYsEWkrc8snV0dWeZN/UnrL
v+rGM/DksPTyl9qsCLrxyQCAnC/wyM+xAo4Qo5t1V015TblCK2GBQz2uRtNoRumYV2nUSL0Je9SM
5p5m3MrxLZ77CU8rDi+/wKa3kznFgVw3RTwVwkoBvoMeZ8qtXCFQ3ZhcF7GcWyRIXNQD6qJWUl/+
YfNIh90Ady+WiyEzMgczRrXBN7TGeqyOddYlCtkms6830Jf2wT2UUONMY2WX58ipMQVMGdqztoJg
EUF3KHntfS1La1dkgP8FlVCXBsAj2Ym/HoCcpfmdq049Lph31V3+IcEC+Have1tv3+IhJzEXqcFK
oW9rW+oQnxVOtYuqDHh8xI2ljbbuoVQNgJcd/M43aEgNNM7jFmsQduzX9D3qt5Bk7pCNyRyEn2l9
mPD+9geYDIBfYn9o5WfMi76/mrrdzSa4QMHYupx+tzoPBYq6j0WrLZHjQ/UQ4gZi14F7+0rDVpLz
UtQTezqp0kyujlDf7CTHTR/lIpVPIlWLJjOLHWJL1OHqf/ESkz31nIefPCDByEqjxLJD7wOtLSU7
FhBED77izkz/ncAgcuqhg3Mc0VXEnGnXvqqB01M2LB9IvO0fHAJZ5VkFstRuqw9RG6RTGZzYmKIN
UsIaJjaGzSNE6TikFsgIue3C2ynazlKzQJjjnBbvJW2jQDPTk4EVBCFHV/OXR4Z19DiR2Hk7X7dn
/yySCfN/3fxwFyPQApliKF1uBV+vIQPggiChwhXkMjg8yS2G0/QzU7Df7t75MLXr7nKTdCfoJfLo
c9ZFIIH6ybUZxbozhowepeEfEJPjuleuzneU4SVLKx9xNZSYU+k5BL/EGNt2ivTH07h7DVObA0VI
XY06KOQyJSB5qQ3edj6bawBy7WkYaaf/d6NjVT/Tu9d/A30mQNfX9ZTIqjdWi1nyrx4fbH7lKRKp
gipvRufGHoy0cvqbV31UDVaE6Y5rvaSc3Ysyq9hMRItt/qXtrEDUMnEraozku5BLAftbfuzfXNfF
/lxIEGo00utcOt1aUIievSx57H4hAJKvtrcdwrluJson8/RtNik60qZKw2A3nsXiGiTSpp7zf++v
HbnWiVSCqm89te35F+CumHJ/uZ75MhftfXqTbgK+L/B/6pEdRtKLzNTCgiX6dq07dTJDpYr58+cR
men+b9Re1kQ5eOXJx2Mfg8Qw3SVQglQXfkWlxntfJhoMruaUlELnkLHKfcPKtRzq8kTNIH1antFh
8hlK/opcG9pWLkH8a6NCASsa0wBr3zXwE7VZz9k2RVaZdNKKoHHk8PY/UcgJX146+2kRP1BAsaPu
5ABNW9Xlc2R/awZg+ufCbuEbJu4mo6uaYo6UORXqhfvlMXYjdGrSih3LAZfrihVk8cQUyOsVdIko
I9ea5TIZRMVNV1BWUD8+fXf0HaEfkgDbllRWt3lQm0edYYVC6dmyUiKTnsyp8vPTp8FDs7rBfCx3
7pTZ6wCx533stCP7TKdbfwwSl60vjI39t8nWxDn7n0A7sawt3RcmuNVMyGR5rtRecnDy1RBtrLP2
jN+xtZq+yUAVRprXCdMrvD+8z9jy4NRk5PewKtBvVWSu8horkrajopeY09dRg1jG+PG2BhY2yoiB
NNkinbkk9C+HPzs+HdUb3737vyzoqsiuYCRJybrDo1OgSmCJgezc+5E5+dPl4/I/8zXmB/tDxWeW
vE5j56Tb2Huqh4cfpJ9YtYpkfKSh/C7v/Ny+/K8wJaBxl3OPWDpSvBMnP/FT+bwwl4rguAkxszyQ
pLL7ultmEp7d6rwsbzZrrfilzGy1Ufq9UxfukmFoNzY9ISS4Dxrxe5uECjuMaTA/Jo0TapDQAeIL
caArrGH9lWNaRcgMRj1sS0LzUZTSsbYlvALjGJb2kSvYBH7oS5HVnHXq/WRisA8pemmq/By6NF3L
a0Dubr8DOwm5VHbnYm6uuT8dmFCqcsbilt/CyzRhQlw3yEp7mECBV0VciBoOYVoYfucspeN9hkdR
jhHIRp/sxHaREOCyNH6j429Up9A1QbBHrRbGwP/wQO3LMqu9LwR8TXwDVh8k6vbiz91IzE0dAmvh
QSKwLc887C3RKbe1GENqcKwshKk/03Q1Y6FmEHyyBv1Dt597S3R8kqKL3kG3YSqjwskDRLKlBR9H
BBeK8Gu0ThJZALabnFQoaeqRXwed3eYMKMAoYzizm3SGwKSsZCsnDS4Nw9PlIxk5lhBVZ+Bvxck2
IKhj4wRM6hCfhec4NDa3ETfFldADd/HUgihwrwrDNn7NMS3fvUssB2ypUMx6mT8HEgMuue7P0iIu
M9G4Gw9cxAcrzsHB712sPQ6Xf0YosN1AwHI8reA8Uev8VWFtoXNXAdMM0URoJVqtcbKglqhZ7ej4
k3o0ZUbNfPEESTU2se8KA3hEWhUXnqc/BHneizGpX5KKmayXaPH0bfuKyX67rpDc15D2qTDAuyDS
jomlf58BlFro6Ox8iMhBDzgYnQN0K/sgGYZa9/AGS0YQGc7c+0gkhNW53YZ6QDt0mYq3g2K6y0oC
M9DHAqvjH08ZEwqv+8mXCKEOv1q/qpUlRFta2cuuGEVsUwvvlM6WYHuXuIdXTGfn4lGgv3XmVOS1
OHYN+cZxkwO8ofEU+7dBuUedQiHCCsH3VZsgSDsFFbf45XAu7SWJs2iCe0K3zZEF9uegnyIsaRcU
ej9ZjuCBQsPACjhnDy0Aje6mGf2mm3Vc0MFAuFvP6i3cze88J1/rPRA0XRk1VPcNW4F+YziLnD2Q
fJzYtzkNV9Jy/hfqUbj/6U8/FIk28iSIJVE5hcxlo7TyyUXUGlwdFMKBXLkPYaIJQ+4E1udlAsdf
DHTEYfsDQPS0IMEh0smweOT8XseriGQsWoMU0TiGga/s4H4VCglY1gsWyjOuA/+qL7+BEe0/dZkO
FfDvgeWwghcdLj1PYbO407Zylm/8ZEsRi9BAB/6yWNdc7/pTSAnVyhodFS3lCTeNzwXcj92HHYUR
FMQGeXhTIcD8HJtvKW7dAmW4SQweqngPxvDTaiARgxjODS9xgVJaD4okDY7mh7LgS7WcinOPAB04
FIbz+DiEE6Qt1wTVFXn25fjLs2bDb4RScTxumkeKgGEuilIl0IQ+R/r1iYfMdyXskpDvAZXhBvUr
feRmIMlex4l55sAccdxeZyxks6cvaBap63/c/gKqVTd+g9zf2Njvk5UWdPxlcmAIh9enFSfcNt4M
FYezsU7wQYlmgR+pAg+b3c4hKNAllr6eCc9Msn81wne4zy74rC2XzuTbPKRksZ2OILI1T0ePR6Yb
wMr8siCBG0YLyO8jMyHAjpgwlvh3tIRNG70gZJvsxsCjVv6iKB4CepOSd2DyXoQpchaTAOG6L+TC
MpZsOHwliLS/7R90F+fjwMf+F4tsE3MTpkML9MQXPWWbFkORyWvsyO+kdDUr7wlxgOAWVkrVXeN3
xPoOMdEySzYk4LVL5vKyUdQlVplO8NV0SoUlFalEqsKX9DFSGhgOPRX2kFCGPz4mtOvbNBMYA2Oy
5n2l+nv+A4UB+ZxYR7dqPymndWbIr55a7a8n1pm++JgIeQJqWmYjnI3xzTjL70YXtbKPe+TdfSpv
SeBZQvVuWjOspY3PIkrDTFT8dAy9fdWjYQqlAvR/bybK8QlnlQgINIZUGIHM7PnfAsghx3EOHy3E
e9V9tRoydQlD3g757Hik79qHkt532e2v0T6+/1XiM35v/89185oz3gaSAf4tUQB2u54sRRuEECK8
gL2Njt5bJXtMBXJheSf1xx5NGCCAedSJZNkjm696TnLmN8IX7mmQhTBWIGzCvE9/fwAUWWdQPq1s
BqNFhCn0oS1m+8oieY9vQVRYZ79uIdwQ9U16BJNt0QdHUqrimBAlqHahPVzoiwcIP4KKQ4mkqvOX
edApYTCXLoCGtJoQE1ZqRzaYVoyzcA3Se9o7juVY2+TId/3HfZLkUj/pqYDEhP66zMugslnSX8fE
QoF5zMX4G0dbJ+Te8R5u1Is34WHtjEOtfUNh8x5RS8sD6FJtgj1QKT1GsbGvHDHRvo6knxQ5yljr
qFykC8tRDGm/UmG6fdT8EnH8TY/o4SJDmY4ugzNXJH33LPURmGPa8VYoNqjvtCJ1CNYOd6YORqrb
SLJA23ZO9yKQWTexA3ve0KdeWRDv0UPiqFrcYD9PRQcI/qvzFN4yV1b4s1+2VN+N/I5lJVECxUYQ
Bnp7KbwUFZCjseIAlj6DnAD9rGzA9p6m2Cv+D52GUYicX7Ov65UO2uxp4BtS++kPfkrhuHo1hu9S
AxGeb/lDl5g7SXAiqeai8O/ylfSlEh4UgTlP8UZwRKV+2ihj3CM+TyhfN9tGaQmJG0+Z0SULN4tE
t0+DHt4Tq916HN/Ts4feR3LarHKmRATOSyI2gZL9KX6hKbEbuyWPE6hri/eCy6RH/NBHIk0SA5B0
OVHAOyqi8sn4/amFhsajUtN4M1oGdLdg8AIoCY2QiYI5Xd2+yYWyMIIMYGwiJwsjLofMVIeF0Wx4
RdU5tKwW9J2u+cV9jZ1pIaTij0u0/QK9eTL6/ZdGL8aQPaNwBtlo7bI9rQAW/fU63TUEWXg6DU3r
R3Y3ns0hhOfwPseQ3vOb830QYZmabHh6wqeV1h5BXKndC5xJvdz0i66cI9OuYVIUD92MJjjhVa8R
Ys0/9fNP1g/HfJUP5/YODiV6KWUxzeujR1LPILJZNoPUTbJYe3cdWiZycihyQVi3HIPdbI70/yvG
jx7p4LEawb2R69B+/wga7WomhFIOMnM17EfuxkYolI7zEb1N2as7Z2ecnHPiSTUuJSUhJYqU4hxU
OWjbpS5onKUB+84iloQEaYSL22Es6TsFUWhUJBp5cQ4BJLayz1/mtfOp9Mk08eWaXyolRklEZra/
PfDRq8gtEXG1Oye+S7iGXZbFM4vDqFs5mejfqyBGZWLBKX7Sr6DbzGSmidcjYRnOA6F8H7y0x/eN
7xvlNbXlSB/AvZQM3UHiobdFCynXcSV+iuYf2b9E255ygbSOe+sQqoBOhgfu5JC3mmcS5DAd1E4q
M80r5C/V7PZFbwV4J53fpD5oWKrXPe4tmAwQJvQ+QyA2JKJvh9Mw3Wy+XddXmx5wgB27wawQ6Xav
2Y2cC3IQ1IbcIdBM9xAN3zQt9IBlu2Fz+WEA+vFo6GtzSv3OntKccA5+0eQ67zMjhgeG3ms1ixwn
QjXfEwagxVNK6Kgxpd5rXxrsJjbH4ZueKAfoYsGd6KCI4SptsQt4EtOM4Imfv9UpcCq/9wGGrTfn
y35iRP1dhl1EQaykmhY1QQv6A1CeQX91PmSSMqW5Fq1i2hUyNBQzEZv5gskFWnJ0hAj/7V44ossJ
wpve6OL1Wd5pG6zQowdQLdWdQI1dJLs5We8CejPRKahaS6tL/gE6u4p3sufaJrNzpV8R67yXR/h+
weEgkVFCcQPLWui+45W0tFOdJ9xkXnRCYnfiEIQC5jT6lnc5Nfigk3y6FIg1NPi8Yrbd6GjpZXHm
iepdKhflg2rV+NJ3KPxZQuKmbxx+yGRjsZkvCrp2qfoDsyENMaPDikzWukCOjoBULNdn+7trpsln
JvsRbokLiiozbTV/5kI9bs6bl9Py3tcNaHpUZ/P+Jw2EO5tNHKR6bowAtTzvL+sDuJpjoaa7tYGX
xoARlzMvZBi+I0Lpag4Mpz79R6BiUJ7f9C7wx4rK4/UDCgsB/dcISwMy1MeuWg2RdajVf5xFfpDO
L5pXU5WW+hJ/JLJAw1n/RdTiezbX0bjwGexSrDwN4qYGQxeaGiiyCXQIk3pgldq8EXqQy4nzFW6W
MPTYWTPjEwaC1Eyhqqwh0sJvcA/Ica7jhf0R5Tqy0VdKHeD/f58hPGyr/NfvRIbF5RNRXdWLhjw8
dGrted6rmd/qeWNh5pr2rBr1UCE8mmdeDVuxG/at9gaKSaAdRkTKJh9SWL6JfU6dXTajn01elYSG
nDA71X/uMObg+S2KIwWaQGcA8f/8sDxPladb4lCpewfRuzaRuV5XYotVI6llgOKRMS5TIrBQv12c
AkbALQRfUCK7DPQZQvcB3Hz1lMz77V/sKIF1kQjSb0ickFdjN6eKUr8L4WijHeSW5wVvJ79fYIla
Yc1wbAtkjwpNEYrMrldRwJed5AXM1e+YOpVlmtWCd/hll64WRMV0ZEH4O//TT7lzVrdGkVhEgasg
LsUPlapWLi1WXec3al6L63BcmqwRlThsPzoj5JB31gK0RFuh1yOnIRXn58KbpatZhTCl/ZlSV+3l
fosytK99bR8bBRv1taNqbuga4wujydYYB8f8yE7u1ZXyYo0BsjQeKSMtTaAzxdJZUY3D1yvEQ201
hdQB10lotcQlpOkGPtrZEfjm6dJgyroJgqVaGUvQXg1CH2d8WTEhg6KloXa/yGBGvRMStoug0J5i
zICJtsPY+6tddREkurBJsgKEYBu3i5JLOv4x+RXjNaoFzNhA5A8udaCipY2VD8d+IPr58ivhHL/i
ERf3wd22Iw2l4QV6CnI9pDdckDOhHg3kjdAm3i8Y8y2C9y6yQ1/+5/mDo96e24ABa80cL0L6HMu5
guQlUq5sDbpQRWBu9sCj3SsY0lubzfh8081uiwpieCT7ifBmDgCr9XiJN8vTDPWOJgvC91HeEz9T
oqcYZE5OPQE4ESQ2yNo13WzxJh7Z13+boRniuwYbplbcw0udKVB/pEbriOuIEusErja7FHu78D9u
CVQkvJDTqP271rn7S6Tapo208VQMQ4JmqsssW5B1tqxdq8wthpRUXCWjQBaN3/ERvip/Wqm3AGFU
dvHUtVhZ3/NwTlaHDgHZFQCFwB6GuhPT5OfjW1VvtF2cvMZMOY/j4NAQQnSx02ZUVXJBk6Wr0zEE
Ri8zM26J69uenlS5upE0ij3xTp9nHH7RmL9nZjf76/bF/KC7Ozmw/ekp5tkI/JqVRq2Ov9fb6U+x
GMAlvGcpq5ohb0eCG9CosGuiOAPIHYJamDHy7LukNjmlbqW5l+qceY1RaSqPX/cG0Ulia62QjqsM
kcYHWcENuPcN+IVshpdqCd0wkN9bGA/FR9sQ52lRNOpWzO2CatZHoz++aVnMi2QM01+Qkz8Py66D
q+LZagtNNYc4w6NEYu6AiR3bLhogWIYzrHuoP2HxyMmWoUL3bFhvo1toBaC6kyMIIM9S9QAtfWP5
5PbgPGFfKXKq6RWEqVyw+y1lXaqWkV1s1m1jAFb9gVrerbpF/CRsSHmsgTQbn45Ley14kty9fwrK
4JNyAy/Mb+VzXiQOXVeXzJ6vux1pJlvayON4dj8D0Bc9paODynOt+APHpbm02MKU3f5AuPGpuALv
SD0wQcYlIqzWEsQr30ay8ntoOhvGJleTdzVSaG6XSJTaZMFmKwPCdg8nNT6zhpt9h+4uGKKw2gcx
QNGRwXF5pV7avYR5lJHZYCQ3gLqPJBISo6VUB0KaLaG1Nfa1cjVixd0STFqs58tTZT7xCp1ra59V
6KYg01LelRhMH/UCWw4ApW3Z3yVlPxaldN8fzgbSJU7nsIB3U2YKx3+Q3/pQ3ZG0GJvEavIrow90
mIJYNM0oTYZIcy5zb46pqPD/ea6d6W0rrPd+YUg3ImL6d6875kn6KH2A3+XV5LdY6+Xb+jIHgpxf
l+8VYL6vWC6MJ2M/ArxMHvXuMjmW5lQCtdN6B+HFjnvLocFGLGFlosaI3R76IGcSUX4gzVgc300D
ultbd3awQgIS3I7/jZ7ZLxOXtUJkxgMw8+BuleWTSvUXkkkNYpXlq2t03cJu/rz7exJDHxyhULV9
gux6aBP/NN4wZtwfgfQMNAf8PwQK0I8+ohbW+HU7MiOvYNwEqINJZGsdK4cuaoA50T5P/cbUQ1Zc
3wtJycCBnysBC61iYQWYf6CsK3tAKJyE6NzwpUfvCW4nktj3lhRiEj+XZDT4vFOYegrSTlt20Oov
XkhfQ8C1NpX6XwQdKe3W2zWt8OvqBIvZmwe2XK97TZXwxOIYnT7w0CzaVcJkavNmJm2ItK3ZAktJ
k3YYbVFDJK34JzODVLRiMXmbj5g9G1JIRdnFxfzoT0A3w2CFKEnh7nSh62WZm8c0wp7dP6Il5u5+
Ntm0ronhvbg8vtbaxETT/Ordfs/8Ru5gGYL28Wu4DQeiDrW31LDfhm4LbYJeuAEvwGs36lTmNvtU
S/PQRblYQ1uLCx6b66CcHN1SIOBkbV2jcOdiM8BROZl9G0HB87nWQWb2PnxF0LuK+XmY6/Fz5v08
cAtd9jYgv2dgyGaYwBTWx16JszWnoGLJSxqxxHSB5oMOPwluXUsc78FTCzCK0loywZGE2onipCg4
8wZLvwUAAui2GiXD2ujCXjfr3Gz8nszHdx7U6Ctx5QLCohfCe9WIvZSxZU/YBNIy+aHsdVJpCp+i
AqP/rWbs2aK1yVy4egk1jMy4hIHHNMn90nynksY8Orp2myPXJLNFm4sUQJU+K45Ygw2sPUVTwnr3
Of6oP7ndoIRjc1kOxR18sAOoha1SW9VXCOCyi3zl90DkvrCJQnsz4AIfK37y+iHirLwfkL8xpz2I
CwOghI7mBL2oWW1qzevwUuEn/zWJ+CDnwIBEMcDwCvIZ2vgKNP0F0FJ06I+lA2nND+3LVCXiXb0S
Dd/e3oGlww4heZAFGf+KR6cEfA6ULENI79t+Kfv/GuCtZ9Eo+djplrzOQvCInlYCNkwRbesKa07Q
kDJtXgcLouLDK+vVTO5m/TKBJ+xKEfIJ6ohBkDIYmr6dqW7Jqcu1+qAmTlTiqf8AfPwepYJeGxlL
9WD8tw/ELYzX4avSEQdutlr+MOB3beg/D2KL6nPFpaTZ4GTtDP4nv5GdlxmHZ+jP2yRRAdu5VuWd
W0u6V6pNSy1TAfV9Q8m5QBrf6Kp8IpaED6/HAywJJnCAPjJi6kpxp5XlxnRGPxH/kT45npjlE/SE
2+/9FtEO/WYUY40+J6L2G3IEGIDmjb93+SzC5Bzu/q7hvrS+UPEekk6uwIodqaCbM2iRJZn5UCvX
nxzZfxqjv9FTOFlCBS8lIuke2IS+ovVuUKFoSP0JGt/cxT0z8TlduYwbMNly4Fz0HLMWa/DgbvR2
5ABP2eg7SgawHy/g4MDw0kE9Zh/CeoIMSv8pOpCJgJ1AwpHqo/OoH1Es3OLElq3eyunoPNamcclp
zo5sgpr/KJXJm3DZkmps2ScBRmQalwBG6WYs4Lcf+13CBfnvLyqQyhA8+wgWFxMGjGHmojTZNTs2
Z/WfFKVvYjEh9eO/j0II0aowdRaNuelrkzt42hiVG7uL7Cjb+en0T7S+rKhscRShyn4eAnWj7I8W
BXI0cLd924fXbj0nG+9Fljmq2fiIok4atjylz1d3VmkONU6lQ7VUKRVBs+GPNFWT+kMdaOcT3oBE
+MSJTaciI9dI00SEJ03R9fMD0VmtCs6eCkPPLZXqmf4h067pQHux/tyt3HBGWMMMdeBYeM9jbyMt
XSBdWi1dCx6F2I29V7bWUAZ5Xh0IutHam/YeAdnv18/rX0fKN/uy3wOuzlFQUJhNwSjPgg9N0D8T
UNvJCkLJqWjsj056A3ZUi+AGzCi8Ih5OZZA2C9FqJH6h6dzSRVpFEbChcRd07RIfo2uuLsGf6B1A
D7YGGP47YIiixu8UM2Xpb4pnLXsclnkRQBy4kktR3X+upLAiLoAEKM23K+BMIM73Q0sBRd5Zi1Ly
IJAJ2IQ8C4PMoG30NdKzhP0O8jxGNIxg++DhNiEV8Fs2ocseksITsOBVuzfdWI32PxTfzCC7GGpF
95KqGM0bZx0aEXSKLzTemOTNjCiUp2IVr1hXcWCDy05elrJVEP+zxb4+G6WqjRjc+3elvpS+QL/O
Z5r8JSJ7jtxn5mNZ+rFHWqSaTqyYc46fUTPJjPNOx+G8RUaxHBgtp9AHaIL16I5epzFIJgD1uPbf
Ho49AnIGPSVZimhoK/e50HQ7tGub/uw+FhDIsZhoIQtZg7DElzA3ML5sNUHRy7rjE7KGZUQEyvT/
pda7FhkExmh06Nvt5VpkXxpDDpf2mm6ICRGdjUGydLUrPcbhYxn/qtA87/Eas3CpDirUEWmvElSE
bFAdGeWfJ9aV1/GY4htCdNUOOP1/6EGk3sEw3ReHZx1ugZuBFcmC+48QSMKZj6A/TRnP+xKMotJP
SM28244lNH1KOY5JSbC1WrEDsVuBFy7zZnjcHhWzUdOMmPK8MJtDmnRP8CFBYNomGn1jdoxIoFmQ
3Flj12WzkKvgzNRFUidtuBwVEBmTZ7/RPQdiR+baB7jl78wMMvUtRpS33aqZDz+Eg8byfemM7gVi
+cy4kCgjkGzEO+DNKEZti9hBs05lChVvWBS5HCByCc6nLDKS9rnU2wxrtwrs5EzAWH7SWUrXIMrn
m9y5xEXLCj5BVSo/BXPWLeh1Vtf1ynSNCuJ5h7jJVsdC08hDTfVRGqeix7zirPAmfizTjfo2fWwA
N6LRzWi4irUvF6O7AUIsxVxmvydaQqM7OyKrvfd+4CSRVaKqZ13d8eHX0wvc/RJofLuu9nHTurzT
ckeEhXAEy+dLiAOKznuQr/R+alxNtukdR6aticz73JJAy6GPvpFzZbPeDaWXHLzxTO7+9mXw2JMl
BKXU1vGaTeO3X+YjtP2ve4xZN67HFniK0xH0tBe0J97LH/fj8f9+G5rP1H5dv78PW0fS32peBIwa
uvGPCWFh7xCL7obB+x2RWcmV+XfaIPYtN0pKOrotbAezWQxLntJJk1KqScoMZCWzS8Hc5mNweUlk
2dHceSYd9/qnM+awYvWg/aq0O+bmiK2+Y+e7sybizBWcdaMFS6kwQQdKL7nn+vr6xuKk4jV8scoY
GgB/OWLLgpyWcAwdunHVxIa945vc50EeMZ5IxBjYXvOhQBHResNd0Rwr1xUDwb8WndpyNTTh1Evt
az+7kGrab1ozWXd20VaIWBDhRU1JXXX0ghD7aGe/RCDjE125GT1qDTvG1gC4m8vwtYcZTb4LREJs
GSLjRJffs1nre6z+bbN4fsLnWNgHho9dG3JuebhLvc0DSlkMbe+JsQlX3Lna93BwGJp2CDu217d6
56s3E+jcc9Juzekl/dynZ0PBB1H6X4C3NhMGTaYg0fEhfbaQUvj5sMBQqXdWOhUffMqx0gBn/5GU
yPEyC3wzE1pupyk9qVxA+mJXSpqNqdcNbUjC65gbvfuubZupUlT1XXvmfN5FaqaqQGZddIrw/XE1
Ss4vtm2AbLNDeMcjQJZO8dAV9l5tAKhud3KGfSXnjwlH8J2kwWdHDlF1GvrcZW5T133Q51VJBAq3
FRVzyEC2ndS7N8/hmjeuyhOhgl9pqS27kGQyI5Q97ghRR2OZLs+Hwzw4sElrQmld5Eqm6xcyyeoT
cVnEtBKLuWdneZHZYk2oSCsDWnTeKC1XIhdEBPEavQ3AMPm9GGivq6+WAFkrJ6YrxF1GTTp3u3HX
JsZ0KTv8xaJ+WQJhlI9dPCytDfQpEOvOnkWJWZGzoGKtslZy77Rj5ZVLR8orrlcipHTopcuUQNVx
8Wrs3bP7JhB6ZECqG4TmKmUTbYpXenyu7fn2VSeX1eGkaAlvNhy6nEHmH53GczDUkylTFoUkudWF
WmzPHbThEmZiVaNUdMjw0yz8LiI4oLF64xFo7tHuHrxlkENrf9YRaTAf1HIICHFDeoOUqaBGYWNQ
dDn3yQ8pcqaSi1HWSvHpR+QbKOKCQYeKmyHVAB2C6ljkXOv2i61v413nSZARuf+y3bpSnqsRpzpF
kFjoHkNMI4CbXXzeuWF+hqTNiUj/9LsLOEY5puYY94KNWioF5ce4YkdbtMWhNcUauVJG1izXGIFo
eYHnFm+5QA4dfXenu5VBxm5e+MM7tMTcsV6dFr6NgqV4vJ3OeYYnITCXJ+c7SIkXEQIJTRCXYrD/
u+lokSQcOIqQwa/D28qiTvj8Nlac+Z2z68jWZF94eY173RyZtlU2yGAYFczxu53luMUCI+MemtX0
ZZE0yEm0m/bFP21g62MNJ6p9ntWO+ojHp+eGrPV0BZZ2ACKlIWKCSxE7pxVgLZisGgsZfPtlpX1/
COa+bHDkephP/HvR6PzsuUSkY5ajmV0AsBNuy2hdNdn/DcV5s/sijDSguWA0y5cv/U57cddha7J1
1eISYfq/EuWrCWp7KGY6JDyhFYRI5Zm6bBK9/OlfKPh/D3MUSxS87Hx+dqZbK71rILqMSYj7zv1u
MhCF2AUlM0a/k/KOWc2NbqybRKQgdRVDyeQp/vdxaLC8061ZCoLSRsuam9pGr76EuzWeQCF+RaxQ
j3s3dCoCxwDoWQJA83VlpVdnSNCJubUuU3ANsqHLL4Tqx+qLNDj7HchFu6H8PG/U6TS/dy++cls7
/WBaJXH+WQ1utbc78YKfKmk3L5A5m152XMC3CC9rAEhOYD1GRMsvqPfR7LIsjwem5kmBPXYPWL3j
STKhpzrhyKlKq/NXoSTRIYWRcBkM1J+SXLIw5D1oYLIVv2fbgqRXN0zGhfK+4N0y63v2v4QiF/nc
XEKd5C62YwyyN1rkpk3VQqIXFaOMjTcK3/ljgTJrQjWv8UKTJ8cuniS3ROmU42ZDbl5AlsjVmW/B
WyBehG9x5uFnRPsBBhu+sCSZKLT4e50IA8q0g2RD6kfOkmnzINRggqZOiJ3Vt71ow+5wR7FZiGO9
wrg3t64J7N2arUSoXXbruqEHtLyjik9NeKz2bqJa3bIK7K3ZZwTbi1a+KudSHwDGTaqs72eIy0jy
Vq0NIzk1yLkBDpeunG2huqglyvwmP7aRzt/aWvbnq0dQVZq1WJZbGNUbzakT7qvc60HSpKkTWdjb
IaugPNI/6ZAvui5owzWnmic27BFXtIP1/BFKaVcbZivkUDwQvDnjMbtacjmzAUFWoynMsgcwWyjB
rQR38yk+qL9ImspaBOAVLiXxEyQkzLPkhQkNaxKsHc48I1zlJVp4HYSlaas3RJkwS5WvdPnrxCxS
2htUvjOXN+CKlVU9UOfc/W4NFII0Ow/uFL5WTihjwsUPfiRBUQyLjpdJfiUu0YKfhx9GKUzIRQMo
1vD6XEYLgOBPVcKO6exktODGpHFpLCgh+GxCfYGcG3Q52dKD+yHMro3dvFxlyPUTGtjQ6ohVC07m
tFTljvwUQCE7pmcIesYWoZsdbYeX2zBvQaoIkAzTq14cD1a8G4eev8Iqsj3+PfQwgFyTpggp6Crt
xg+0IuenfBlfIToV/fXoLbkdLtXgEwzzdnEP4Bc7DnBPToU88XbGCGtHL69FxXfeZw7cvS55zkSM
xHaCmsSfWC0QqACujoKpMNIa9KDnMLHGAi5za6emcOM5kzWqpHOivhF2JLpKAro/BYUkvYgbBYGg
+e7Q7BJQP2e9Qn2+oEd+s8pmVGsMPqGfXFxNkd9io177CC8kBEqWK44uLI132xR3tzEf7gTRa0V6
Sbo2lpmPgcky1TC7A6/X1jtKtYCrKEjULqdvV/rP/dseODFd1e49fVEnYKsNKzGAz5pRlBoVtEc9
TKue/NuTCzXTs8WGJ606pXLlS02XmdLaL2zC2JmTysjVrDEmcr6Gmy+neMr/YsdZhQy3Zqi1pnga
xBu2MB7lXgB9wwHVdly7PhyA8PMZ/yStcw8b3PyIp0cIUKe8mMtwc01qtE6VTx/gTBSh0mU1oLsb
duurbIyoahtjFnWyg7jDL/+lCSRfvLb2qNGx9sv37kCDHBjrp5ldZ8Fwduf0pb1fpUlcw6eK2LzD
ewPEXaIoFl4TFAwH4bdG1ryPdWituA3JXornFf3EHEFwBGdhvjdE3y+mKA/tUHNY5bK2aYm2PITc
rM9d6dFnUBGtijCRmRuHqFBzykgGszv2ZwaHwsMDSAfH4qWidU2o8WOWK/+OEOkKZTtKByFM44tf
4hAMm2FNn1HMxzozeY9ARGBum2ed2J30O98Mu+FPDXPntQ8MfL6oJDwzfZ5PIL82OzRCrgmGYG9m
YPo8g5sWUs9MfOxVOA5SHOAQ5pxVgW0if5kFWXC8fRUc1Hyx8zln6ficMkYyQXHmVpR+bOJoclSC
1Em+sq2hsSmlyVAMB+p//c4qUQ5EEA2J654gF3jvko0vtmBopqlri79mo67IYuwAjzwVkejqLyK6
qspd34BBlrABSnl/YVhWJgfnO0V5EPwONq7ki1FQvKr6s3Kc/6WefgC5HdYn9/JzQqiFc0c9H84m
dOjVrnrsvmUbDmSWgbcvv/fPjYzLsA+ADe/siUuZmtMh5P/XJAaZhBTi4bsviKmKVRdQI/YRG0/z
Rq+bnGhla8yVVL2leHZvTEcVueSo8pA+uJ6kou4FTe9ZF8vskO/5YME/c+d/jCvGhxhOtlFt6oJO
KFKMfFr+/vAE4a02n9gW//5yYkbnYdeWIoB7Fi8PNgiHWmWfMYy11pYyBsyPc/176zSn3HA10x8S
lmcs/IJv9TdwF1fAFf7kd7WHETXl8m7civ8x44f6FtkdQmieOdJB6v+8Ty/t/d2F6PRK97wa59YU
xoaa+d5HaddCs0uEhsVnIl1Ab9L55Fe39vXkZF04nF7sKXU2cafMv/hOq2gmXqImGmCk34yHvDuU
Kt7oXJU1dvB9KSSolg2XwJbD57VPu4yUBlWR9f2dQEmGJjVvIt6HfU/Hrla/gppknVD5pfiTrXBO
goCtnjdFh7CIVWFuB3tdzouazJroMSFTfg3VT4+YPYVsCRspTHiEB2suxaWlRJnowTwePrB/YkZh
7QaOF+n6LtFcspS71BLRjfPlTG7olVCIGLSRn70vIuuLSck91nCYF5WFjZqC/PCAcnlu4A5+DG0q
jtcnsfexMnfDaRSJpcz6RLKlBecODjBqxq0G/6Zwn3kzCpsMuUbwd2rdgMcvniISNgp8sGae1Zdr
jZQMiz8GPzwt70CQz3i32Ne4wZFA/GsNQ+mrMEMiZEPXs0azE8J5OdH2e+2oa5CJ7/Yv0N4AOmux
q2Q6GTD6HqasF304uDAI4WxHftSmt+gnbDC4zTslOEwVMn5lYrHeUfS2f74WePHTlKqzgLFzlFNz
SZNiPB3t8rb6fy3iF/VITq7qUJLf5fU+enejxUx1Q/VE9yoXgnAroJ47BMXDlw+MlMpyFpxQFjTP
gZJ+45rlMfwrQPNT+i7Joqiznbv1ztAvWWqGze6DmPcD3BmkZsBZXvO1I8ACDSdGcTjJUef0kvo8
fZylXywijkGOQJ9p0eXsJNNIrcN5KPmSC+qZNPQdrp9086ymyGko0/EFu1b2C/Z6NY3g57qz+wAG
k2UTr8vMx0gt7k5KGl+pKygxyosVLd2vjL3o4TknnPF4Dgeh/rDUzPWlkvfc/7OrZGOOcx2nW0kH
hikaBmlNssh4sY/25GE3iygYKdXUU+OgDx1znt4XJSraZ6Aw800HbM1JmyqrNzvmEdGjA5gll2TD
6aBBhXavE/UYDDTjspGIa3hbZs1suCicHIh8YSISaghY5JR1HuOMncDdoHoAh6B9gtTSWOfiV6YV
DLdk2O69ZnCoVCkj8+NF712oaw43Ww8yKkyGOfKxbDPjiHn5+7OwMBMacreb9J7nCYzKrcE0pchK
Ak5JYbruLPp9W3aStYBuaK1WVI6Gh7uHGyIy4UGjgIA42075ejozJ9/LQbyfQtZoARN9Qrka6Lfy
qge6mKfN/4ydzV0QKvmThGXCspoYlZPvll4Nxntp8lwJkwwtNAMqmdCrjsBwS9FieC1JndgypEJR
/17mb80FnzbJCYLD8WZ0ZcTwc70NbVAXgU5A40tY3g92o74QKxgMOWzv0aAlKjdyRdX9x3lf9Z8u
F55CbpORP8nSu0VQSP3YWSUwVHnBJMjF897/PagtGeRZRZL/oXWeuCM8BI81c6h8FsUGfS9enDD2
bYOJsFn7ROpjWf284Sr4QyvPud/ASqNAPN+jXSpFAEhGydrq0bO94u+g/AMDNjAHP/3ejTCBYbHL
t8/jvSL6firJKbwSFfRQKrVf7pvlLCwFYyqXTL/QOQyW4koirvriIFJy1U4iYSjUmh9r5Tvf9ny6
T8jqhRTQBFRlzAeHqoU4O2+3e8VAJqnfH7iE8Qcaq1Ts0Uyyag2ApxGpNC13y//G5hVELpJlBsvT
9ozx3XtABa18lduqA/9+V1uco/i9FFQ1bQ7QfLxF405Dz4vKo2k3S4BV8/JJJy8GN9REtojXG6lJ
v8xkk5SYZ3vee1be373aNyzo3lvtlL49uYMpzAw2Sj+6nNsFE7bWY0n/z7iUrd3b+XbTKAcyoUfq
36HknlfQqPi+YqwETpJ/4RNBOEupLZK6aekF0hrIZ2y4+Io5LuFuzHgZ1fPkmwviYo3NdZOaZi33
ROZWq9h9UL/13BZTreOC9WhfT7KgfS7ghdE6y6p2V4HRZYJi2qiAErOTRSM3k7lrbOOurzIIEtg1
0y/6vfzBrieBph8J2nEspU4QZD9hXjd9+EkiWIQZPBZyGCbx5mjM0FLiPo++rUIKrVKjq6YzYFjx
chD/V9icfvRgBFTMSDcVxneSgNieMGMbalYxwdKQgyIFLjPx+lSifsBaoqmFsAquqPdsuu3Ne7vc
kF5hFDnDIjE2sOIlrdJ74q1m2RVT6riKYqh3nJuiAroXLk+s6QITEFSi1l8zRFhnbU/8nGz74G3L
sLETuvRsCNT3G7tK8Fw6Riz4awn7BGzwItNAxQsKOE4PDIuvby8UUIfZa08M/ig2cNauy4x9kzRe
JN76g0E1F7MClMTMU9ntmFUeO3Qsxf0/uKuUMMTdHKK0u6s1lTVosEXNCb0XvFUX6FPkvxc+lV++
BOyp+EsXPyEJGSbmh1fcjk7Xj5sLuyJt8SS1I3lRCqSglg5clsyMB6RXibIYiUPkfipDKz+DDs2A
1EzqELJphGmzyDdP9Ab/lGT0VMADuoUIpFTcZGRgBaCVTCqw7tpjhdIYnbS8NDTh6DlIfm0SLfhA
PZG31g+ZFfU7dXZs8NQs/sZiw3DRfi4ZHy7TvOUlEbVPin98UG54kEiD2EG4JaOXIsmPPsBV55vG
xCYPCJoXYxgtuDJ99UHl5IQJd9kpKuBD5zpfv4nzjkRApgJ9uK0sXGbL84H7/eE7FbbeSFAWfhcY
PEOFrUhQh6C1awaajpt6lYV+6iuEQX+NFLpB7pyuuhCvjTxTniDH9eDkU9pNeyNSDASHUs/AImSO
QZ7p6PeM+0R6b69FYORTnToy9uHE//Mtp7vdGw/rXcdAr3XgWkD3fb4mvtkziDhRnXIiO1V385/Y
pthUKViCpBHza12pB0hU95lvlJ3deTTWnZQoySU1bZppjN5QSUqSq3KaBODsuUzRqZXAbyii2S9U
6P3zJgqYMDdxBJzDPG/+Ww7CJZj+T0Et+PZAE5NyR6a73NWwmFF7XgnDfIAN0pbYI5ZG9bwzZ4w8
9HP7RYYvSqwEVI3+214nweaWG3ejyKUtV0DnuxzynPb52ecyZrAMvC+iEF4T9iKVZzIMhlW9GQLA
yIuPQtcm7+PFGBl5MtXI+gsl2VJ68Q8r7xP7TR2C9OLUdqO1RedC781/kMASpmAbNVb6Ts1m8j4T
6+CibiRJt5TjLJyJvRtz4undKbVgSdWERavkrIJBRVwvY++nOB/0EDr9W+9Qz00aw8iz2hNjaUre
9BdLy984Y+5z2iecXFpshRZyGj6TC3biMu4qliSgN3xbAEzg0uxqOSiYecBBz8MjzFj85mgDKnQg
iTdOrQOKDnDlJw6yrxwJq42yIVY16l3ZStvLA9xcP1p3pUCy01U4TWzcRBD2CCt86LQPFlRfZaYc
ZbhwhYqHAiUrxkSnVVO/aZtajX5eNFpg3/7P0/IbU3JAp6qxUUVk0cGPNgz8iUB2RgzT3M6ytVI5
jJge6RUidfXDAYHVeT7+MyY1QhKt9DuxKfPQkdY+ZNi1+3rCl+aIi/SpfgvzBaQwPdTfj4raoQnh
UCvUVI1iPRP92vqoXFwxXVgBZbSDDYQpCSSUt05c9aNVkiB7h1Nrk9x0MNgSM5txin34hzDQWcFb
y/9/YXTX/8tP6fIhqJRlb/92fJdX/0/Ghqgela9V7JIpjFHwUREBCKeRwHHt8ZMgf0o0qMCdg1F9
FUQJSUQfM7uIeA2bo873c7xDqPJrlYPzN+ZY4Z7DOVPGBprqhw44hSjC9+wpV6SY4AWPeyRzTbpC
F6S1sPfCwbV9zoPceFb6WhcxzjLzOxGPkuf73PQl8NHjBsGV+MQvEkdzhSN/6APUntuhELHYRzme
b9KG8BV+u8zvcRGyaQ9wcXcFDDUILSDaP21zkjCEMmi0MSaM5RCyAMGG7i3e/7lHAoE1rm9WAs3u
hlYnrcs7QVv/2mNOduM+IXZdRiJOME6qzfIUefJmZzeJE8zwEcKjx7RyN4Yc7AOWpihWdIWT78PK
DeHenHKTvogNu+zEeo1tr76aht7Kh4n1CQMXwjq4dCnu95stZ2xA0yQ1XEIUOT60ertGCQpIk8Hw
nauUhsvx73lxNqUbFOtPPZZcMjzwXEcvUz6rROrYash0/orQW2Jzgzs/fxdk1ppwJG+VaVx++uy5
MC8SQb3RAZjdFtquCRsWu/pNJF4RoLqjXp92nZgA1C2dtkPj/WFpKOS98IrGlibo8xexM253KJhj
De4ldkQVNOVpf5TovHx3Z+ApWgduonQZ54sVP2iNy5ZB4IcuYRZlF2oaNHAciNZEFBDfrcyev1A7
rpC2L2GVx6kV6cLTFe5u7BltZdUrgdMqAoCLaS1QwJzNYE8CA0rhP5hjCEVCKEfy2tarDXM+lKOG
aoMTlpMN+egLi2IyMeXTDVCJrYe62o2Gr90S5xyEPT/yzJY0wMUFjoEmr4yuD00UCIugyRMtdDo3
eegJdOCUSd901GMmf7IOpZwYbJaAM6RcpwKkxHlZqV5FGmQGrcS5lJH2LmjjoFsCghVW3Uj1WXNs
+AlNA81UJvtlwUpHo0yNho7Fj3B5rug7jlyFDv7rYSpkWCtIdaP9FyHlMOU+oQLRaOikciklnj2U
/dEdzAymXm9UdyAqUMouFe/gbX8rAIT6s06HDY0jLnlN9jJ2AXHzpd6kax/e8bU9kk/2MIiEoU7m
7M1DoAv8kI9jWvLYrpEso06FOZbt6miZslFCu78i7nZzsBojx3auPxhvrVQhdnoeMgbbclGt5L3F
v/ermPWg8ORzgtqNQm1H6rw+kFdH693ikVzpgkYq0+Z5d5ljZpV4gcHJSf3Uo+/Jj9hhLs9yyOi7
vjKrBYIa3iWwz7T9vo8C//jOg/Bqfoqlv73YcKWAfIY9wRnMKF8hwmdrBANOLDkyXxTbRf+U5AOc
p/wBxLM+O09/4ofxznvXgFNA+6n5uXLKJEEl7d91DHfcqXiKBKLvXyG/Luc6N9Yj23VWnwNaEZGF
v4IgaVSB54b1YI9jdzoltnRMBr+gNVhLyIi3oQ3hs4DkRKEvJ/Jz/N++fjvIDRE47461RBTY8Lgc
TaODfqlTh/iZg34lfhSGjxHHb9+qENHbPDCowXuBOHErBPeDfeBLLvTU170hYTSgUuMqDqVpCx1q
qLG0vl/KfRGhmz910EyUaPk0gzNvYk760t9pSXMA2Mga/tMxyNP5THOZ+7HL3jXUTnMYQK7JFOKV
5en9QbGPWIR9lqV6z42XbPV188EvyyqTqgV04sWLoIY2LFRI2Or9M3fKDjQqicXMy4oCt3GTTKYM
L5nRtfFngdXT7lTNC9yPi5nxaDpBaO0yorVbMu4Y25l+W0JqLYSxwLiw058wxirV6oa0t9FFrjMG
CM4IlufWHAfR/bDGhkybjG23AHJoV+3/l/0wduV9DjAyYwdBRfThSG/ihpPWElSx4r25EKTzGEWT
qWQFdvhQUuom/joDxQcQgBc7ZFvP2P5io3gS+AhOdMebZfPuRZWaQlccO5Dr5jSns0VG5WlsD+Du
5qS6E4JdSo7bvkJr1YimaNuhxOtsYMA2JMxH98flGfbudVPenbzxTqf4ckSmpvJ4vFVQtsml8F+M
YE9doxTBQNaX83us6HN8T6hh2gtOlyMthEB+O+QsF49zfdG8stOqHP7ctxZqjdb+cUBFrFL4pK/u
8uT0m0s5ILVSxRxC7Az0SPaWiAEA6aG9+8DplpQfSR2fmrPyad0ItRzNEEcOpOAR+ioKT4BUE0kO
g1YR4NWDUGS43KGzcEPMb9ELLhu476eV3Zi7s75DwtQmAQd9tRgSZcHnWyboubWXEp4VFCq9MxBE
b9vE4lK8GPA15Qn2R8Z3/FtkXCSqKhp6JhMF9ztUFGwCVhHqE+jL2zWeB6PZyYE4WACbaLKhc02d
a0ug/w5GM880NwE82DxFszpqy8WllaadJbjJXy9j+6Zg+scnstlb6Y4do7Lb9bTTqaOSO+FfNf3f
tpP2AqAxpZwslMrzYlkB115h9x3ScQz7HuxKBRqCJ0gC3t5hLoRK2m0iFNjypHVDGBJaCYfx8wkA
CXoPN3cDKoFCIqiEsX8bMHbbhA1WcCmH1pK1VLt7o6JU+I2LXmIFBF0yn8ZE+ShmJWYI6ce+k5gX
qkRxhi5SS8IAZhZRhJXrF4EsWsUq9l551Cgk1/dnvniT2tInLsQiD4PWRaEldCYFtWnXfeJC2n5y
OBvUbtNqDvxKtZoFlFxXPbtDcSCxxmJx6W9mJpACQnO7IAUXRNN0e93YTr+s6R9zbWMGYG6RIPEe
hR5SKnDfhiWkv8lgIwUn1l989gJG1G/Sxb90jGu+oODWLP3zmzC14hf758HQrCz+jyqX2wG0Ud91
YY2sLj8YztjeM8xawkjuFBrfa92mCtS3CD1jXcubfUaY0hqvl5uEZFDqkNgdP2UkxtbZEhRfJlqt
j0LCh9KVKKd9/d/HkfsLDbfidrDiFk2Ep7MDfTBE4KP538t4YR4ZQbWimDRB831fYJUoeqKRtRQ5
hFjiurcEtvKX2ePyVMbR4PciCsamIClQ0k+Qk2C7zpHJxCQIi7AjkAEicjttAMND2HlgYaWlOHEZ
1BK3yhB+upzCPvC6fIM2lMY9w7eqK3J6o/q+r4wMZ3pEsoX74KKfKzqpHb/mGiTgEOVKy0Qqccxd
Tcqi6l2Iwpqasp6mIPLvxqwQ3LhTdNd+EHzs7l6eJQyy2FkMeyxWGWVqBfM40l7nTM4cBXxlMwE6
GQtaAoqV76fp2H8LS6RHOvp0I1zANYam85UOcDkUeIYKtaruHF6g0FtDDpmsZ1aoqAY4eb/zA1Kt
7Tz+chuRN52RxbTMbXlMWyuPk3Kt9lOH31+PSYBrDV/ICMzX3xhR4osgLqQduYrbawkMbjBC6ifU
Zg4/5DKWym5OvQbLRMVcu6YGOLkC/oK4XfrieGG8EgIa2gen/CLu+K6h7mLYAN8Ai0gJQbB+FRPV
rPk2tTzilaf8qqJEW3OMgTfPYP3qXx8AtuDL+ANtDda5i3F5tePdDhg+JCP6fTnylrZtXsfDgVjm
34HDHwNlhyrU+mX70Zzot1Xm9LlKe1v95W8BkcUvhpaGq3ct/RU3nnFgU+sKU+q4gIobRbnHr4Jj
vUSSG/FPzp+InAPpp3cuO0qsC8hLrfp00GtYJYg8FA5JOdhtCHCJYQu28EQD5Q0OzMGyRk02cghk
ekrAbN8MKI6ewNM/kenRdGEX3dsK/e/cbkiIK+llDoQHYc24gyUowrNJaXYcH7VrqLj1rzOox2rm
vvNZfiFVP3R2UpSRNxbL0vDUlv3seCt7hkSkmWcF54ckAk0ao9zZf8+xA5w7fW7XgsdlmpP/ccIU
wlN9NJlsfb1Yd6C+Gz6HsjXBIpJjNytQN5GX5s/6qGQ3K8GJahUxkusy66wfiXaKYc8my8AwFXa4
cWOpotcIWuvHb0+8V7cLJ/vYfaADLYlc9oxXgTpDINntrWHCbpGZkbEJYrphUi6TbThfHOS7zCdG
NhacbibczkQFLdlTc6puzYbXt5fmZYXfL0zQIEP363WzSko8oIWAqEmfQ8a+qZo5Ym3gInams1Uv
gbftK8r1BBRMTxVbSqwLh924rCjuX+WO+8yhL40dxnNQoaERzEYxSJ4ySKljqKkRa9icQQGEt5wJ
FRxrmFL50gSHxR6Pw0ke0ZPnF/ORpmkRiDR4DyA5q+L0HBIStBTdkpm4k8hyCS+cyXXsiqFhhJYC
p3tXO2vkyWArEcrTDVNOxPkeTOFz5OgSt+dZ42QYfCGlaQkDfWaeQuN/mwkjw18/vIsx9V/MWoI2
aWAiij6oe1hvSO3v8aOhnhUyCXpjby7Y6Qa02XEUPNvnnwswEDBP8jFB7CDz39TOr6TrbxW9NmKG
cSjVQPOnpzX9QISBVzU+TjrbAEPN3gClyi8MwUywT+wKZOIzOWfl9eSMOX77sBjjduFUkxKmu0Xl
PnCkHDBRYNPwITm4hES2Y04vANSsil0eeuo8SBGwvS1BbhmqxlcTTCK6fKcrVQjqOEYf38fPIcB2
wslHtg3CohmshOUFZg/zew5fDSuCdGhgxCpHzTcAdKORkNUQHHoUiZfPO7ZwFyjpiSaIgvVHPQbS
Qy6lfYE01Lz+5nGdoMlwnxOGNz/M0nDxUtD7WGCT9E6NjcgYQSogHdMSGqvtiu/nb3dOQTJjDeXS
sQfIoWI+HBrY6RqHwEWAgI9edIXUSJ//ksvebSNk4qXNGsG4kjanvqkDgk/IQqTHZnw8IlneZ6bb
1M2wuMz2Wwkoxb69oavV3fIbFBLTLCEmAP0WcvdUfnidE0Q0T/9oL9cx1Hci++Ed0mkHK8tBhxnq
sPKcj0jllZ7RtnDJXzrJqy87RQiwCuJdwRAAgnrfpypJ/wdDr77/AjxQ8iRIbR4++Lyr8VeotXyp
OVYLJh/8xmqK6Nio/tq6XO+kmYlezfxSrdALfzAkQLnhWT3uPlaep54K5zbYqlLt0O+muMIx7Aec
/r1tnL1sWf3ZyOilWx72FNE7HOu1UlXEG7+WsOlYbx2R5eDTIS+j9tCEIPicJA6d7RmaVZmEHPTY
7O0LY7OWsyCSr19BTYdbtQywwbBwvR3q6NgZygjj1jUcgWjI4eNlsLQjkOSScl+7b1My0tfAIiHN
cSa6EH6tEfY04sMTdKHlGZxtOh887Xw/nIixKz9uPk3kdoGyGFlpZDI0qPDvYS8gW+AlgVBABEcs
+n1om5zWbNCZyMlz37mMi4zaRZVelT7IdI5MNb8cc3spdshq/fnQJoUdmmA8JuDBJN/BAixBZW/+
tc0rsQhT893Q7MCDvWqS0OmwytyeaKjo0XQArX+VtUnSoV2RXX2cJLS72MlbufTIgicq1WAEwnL1
bheRe4FOzkUxV+Oam3rvSPNaIUaYX+d9nIcZWzd/vi6Pg5jjH/DfW/LRBS6OQYK4WyugsnMC3KZv
KmI6UQ6xX9l1ESKqyH3mttBSKOx8CSoKxOrirtVLEsOiNc0N9/moXDAaQt7MXwNTkHEHbdiUg3jI
RbylQOHs+Id9BdCIlebznT67pZoXfaiLiU7hTsK3SeXUUzx9vF08G/fQyJ5rOmmTQgAhF6GIIsUJ
WFfC2prH5TjlCti+3/Rg696XzL7MHr7LIyhHYtsIKu3FpwKhPk2tv+cYJB5I7Dt0iuj3aQOefJ7F
P2rMoMxYgiPl/xBlhz29Nl6cgxJanIZpW+YLBldLaFHROGGmOZV5pGbV5ct5Yf58V9+vilt0ZLyM
TahM1mezyscqhLp56EfnsqS4DBfFMePqU2mDVQXy2PtDojANk0T//Nzf9JAlkFXurDWm0nxElgnl
BjhK30kz5LBFpJeGOdrikmr+JLh50rpG3GxXiFfNsLT8nyY5i0YLSeQpqBqeZ4IpkZ8kYH0mLcBW
LyqiVSatroflGtlOVPC10rlYH8b/AuI+u3Os1PQwtwuc/pdBRG+KMFinb78IRhFh1n/XEfDFtsJm
xYq6mplSplwOyeSoH9v7qnP64ojv8pDlMYGhYWzppOD95cYY711kvVRBjicVF2uh70PIRpvtOPdm
XRUnef9EcA/AJIvurwxQqNpPSZPNgqDxOKsmQV1vJN4eTzUx8OcDeUldLnXB1iUG8fmOjaQ+qmY3
oiWjc4PglMkizQmCiShZtvUAvndz0nAL4JZ1eOuRY6czSyAJd4AOiDs8G9s2Y7j48wfOjyWBvXCH
pgf2MmfB9yZEVYA8Bs2zBgP0xMECZnsDIki+/WM38wmp+w2+OxJBrSS3xMR0LvI0y983+ciicSFs
OrwHgX2lO9lfT4qcbk88VJbvsFSy0PoOC2YOkjZyW9I5nUd8x4qocT9xy0P1vnznEPXs+DWoUTbm
fCxNrIBfksmF6x6MAFyP0vjv096gr8VuDI/IqqJT4cEAygoiGmMR49boz4xc3axawoPnBx1Dm+Hf
X8IKWuJC1VSqwj4CNHOAA/nzrFLK6owu0dBboO2/90Mxm2GqyE1aT7SlG4OzIrA5EU6a8CUENZyi
ABQB7Jxe4FVigncMF4w1+BerUyLEyNPzdOOy96s+HvT0tG05KsXI3M6HAhH7c7Q3tNR5t8mxQsmo
IfUUVFpHSnnlU3xWQK4puuTN7kDEtqhSMl7G+Hw1wfleBDEF1WXUKr3GfbKwMwJg1GkA6iUn5U5F
gx+CRk8KdxwVulU5kgfAZwV4wyfb5kCvhbW3yLgz2Z3kuMVKE++BmHOEAvrlTiqoVuLfFvRZGmEL
AFshuYvjh4c4WzMrF29565LO2VBTWGuByh918sm/piRHmMalnmjs6+oPVsbdZC1AiDCQ1Tq2NRDs
qhiG4dRiEKuKKC21PFZl0w+1a/VXL1DTaFionjvUhyZsJkmyteoeAROMwDnK2VAhfpJPJS7oUaH5
HN4HDOz07Lmp9NBNzueN/KuOSlPf6Gs0X2vk9SEmsitYV5iKs4SGwuLEr/c+NqapwAIe7V2gI379
LaYIQxyYD9Su6bS6Kg/bb9tmfnqUiY1xH7pCo2bo+/wWRcI7T85ns1TwrvMBqZMajVvYA05RuL++
XoGzr23SiTkK0WFPLd/byvbc0gaH2afp9A4r8QwcXOmkBR6vMVK+vlCMYTJt/4tIo07lGRBoVvrS
ecki7UuUCuThiXsqt0AAnNtcy18QBEgFi/PSHjhWM+8r+++bIhL23FAmrSr53HTFz1+vGfWq8D+E
FLR9SpO5VpQtnrBDF+BSSwX7VuDxIkjddEthQaPT4Pc4N0VxscVMHY9WeZY4kIEZYu1yvI7G3XmJ
UWOmHVxYW1LjBRrNnnDJUhr9/LxrmdpH1exngwZzta7AbYKTclA6ht6GAA2y5vz1cwVzPF2UltSS
2gTAzw0T1lwGTCD2JKbTCAKTSoqThXXpEqKT1yO1uMjs8oXvnGDEvjPoVVXUcJR2lNRwJBZVa7sM
5J+Xkp013ffA3OIeNZlCqeWPQ+JnR7G+CwU9miHr5aCQFX+VugfuCrsX9NWkiP57VngTCkUduHKr
xCLOKbkajNTQI9y7CutToIkikXDueZRnw/i2V1XxywFjrdK9xvXIa6/fdrj3L4dm0yRAxX3oc9OH
uT4Mm7imQhcIpDVMrswa8Mcyq7B7gv7yBrjiF1p75BxUD+Fb2/KCli14CXx2hpT81T0cFSpdhMTm
IKDeqIcWM3h4bvqlTRdYpz0NhIxKapadgsehmR5ZdTjV/stdaTcANlBdHkTz4Dj5IhRQ8K7WXVxI
pJAOakTFX/TkDYS7u/dvTxa6tkdm5wvk6+mP77jGSiovy9KBhp4/hxjB0kSv/QiGEHBgvDECdmtu
7gTD/oZZ2Pe+pDeBGtzXUcZtzCokeCDZ157e2q1GdekcojsaLoLAjVD4Sr6mPfMc8KfkfE33ETD/
ME3ubiqtahGL7D5JNdNZ4akvnSd4keK5zZNTFvFG+n1/O/cKLoCJxQ9b7jppYCrDS9XBL+IfFbAP
SU5PfQxNBXS9tOp1xP8Jq9CxNvNWvBhKaiCStUMNcgX1OYDjkB/XRsjSw6ZfNF8hExBAG8VUQtin
MtxjKgklyvG6ky0WUaqV9hBMKvsv3lSgOdBI5TdUfU7bruGwqHqzcA/Sblk4dhjOv3uHaaySHaNy
D1usmrG5GQ5gVnlcZXwTzAkWnN4r8NIGqY89ZXU2VWEKy5TutN0nHzcfTmMMcN2fkWV8nhMezPzA
7MhNOR0n4XQzD81Gr9evR+EEngTJeKghBQ9uC4Dznn/jjdXWzcUGsqqgGPSQskilP/sU2P6Ug72i
aWB8PQLb3Ed/k94WMxQ+ms6HJgZTbrK47WlH1usMvVJyNoMe/cuNpx8v8XWgDQec84crsS1fK4K+
UkjfX8/sDFJeZN9uFBXL45Jd0Rc7RrkAXj3XX54Tczkm/n8yry5CNwj73x02nfesSl1O7p6n8V6l
lI3FPGLDH8iBB1RLdblJCbYsQ6asaAjnX6kLQUaT/FrOnZ63eKWPvNIdKvg8LmW6vA+vDsWB0Qqg
mnsW0sjlmpgDEy1VEFiatFDtZm/JXSlJdfBY6rjF6Q5mzGL1Kkq1tDXSQtjRFdOnH6FBubCF78eU
RIXKFqMQYfXglDju2XvNYtcFP3pK2+ACHs8mZJ9i6NwH6Ucsrlywor3hJsXmkR0exlWN8bJUzQYp
K6lqxai9z+oj2Xqvuk68Y0+7mmwnuPVOJIQ34Ns6pPuBgHj1v9++40eBSfYKTnqD0vX5kN3PfsI0
hoGg/rnxqDTy+8HSshThbfNgGPw3XGE0ZcAk0zqqSElBmHnDUuEu9/7f9Iq6porURojJX2yJcuB2
Y/7jnM9uHhOcW30nc+bLjP9unCqEzCcLF+i/rsGi0IDzpFInPNtW+Nu8e2KB+Rda9f8prJsnLy8r
R6GLHaoL1L2XyBJf6u6fIeZY6aRNuMwgpYLuKrjkGgWrOcl50/hR1DttvQ8dDOR9s6noxw5gqvkv
zKv1r0L+uVkklXWCFGQgXjrMdXtHBVfonhnNbDYf2RJU2Y4WKdSSBFnYVM0zbL7QQomI3iAhPyGb
oDHT3KZoVlL3L18H8+HkTL/QcX//85ASo94my/UnnXKH9zK9LbwJk7PauW/Tyxqo4OOKRe7US3Q0
9U0reSvVlJ04OeQQ6VnZ8oD3ZkHEYDxnSwmEw04KUkp37iifurgjXRpcr476Hz2XAwYEKBFoY55U
H+a9Tu9JTI+rN5xt6c6dOKuIPA2C+FFS8Wyk3EGsZjHqWmPO+R5V6BU9AA8k7H2oJeNAr7vpuBZP
6xCOAJArHiQzNHcnbmiq3+Pp3g8YGFe71GUeZTJc4UAbNy9wHLr2cIZX9DyI5V4M8PQ1xkLaa271
0+TNRdJhx9qBziiWQcmEptCyRpE8t9ZfbzrasOsnvEUUWucLw6KOXep9haua8/dFyB1bwVx06ZN7
dkkXzSz4Ggb2zD6eY0XBprE6gCw/bjEfH2lB4IoNNLukMLGJ8h7G2MqVQ6fASv1RMDkcAcgkydJw
JkHuRgIum44VyhrMgEHLLb79L7CukF00AYrS5/A3uxmvE7sHv+Cuk4mTJESUOFbGOH7eJnrTw80p
swA+Afy1XEF5kkZniK0wMhERqSYRTTdIQPW81PkmbJt9Z+QN6zOzNx13d7bT8wQ/J0BDi/mw/0Ab
o1lkUV6OXkE09Q+nhnSTiYuk47lBpdA2Td78GL7JV6Mdql7/yx7XEDBKO+/qnlJqnT8mefj4ftga
mjRrEGiDcEEyiXCTOQ/NOTxq1V2GjEsMNASYUCtDdCGXSzuJ3NomdqXZlH67vGpevJ6ew53e6vOO
jIWnV9BTR3qjsTyCjT4rbGuiFlqVBFxWNtygg2LNh96e2ws9UBf1OeyxIsLkpwKXdTgB8wkqqMF6
DDsHmEaLgHH2lrf5axPGbpjf81weyOYu4NvMEkPXaYkaKSDAL1vzvSA4qFDhJk/Z4QMcsKR8O3MV
bQ4zefDiPQcUQSlLXsVrRYKAo0ELEeZ31+myxLsuZfhLT4Psy86jvhxz5pYGkJ+jPBsa79wWXBxG
JrLQzfosGJ+cFkeXx2kqSUbrJ83l0gRaVpxzW/J2Ov0wDtWChJfzzSkVBBHtzlMGjDln3VMmlXlJ
/0Jph4Pa7gyI03fiL8JMYi89x5FcQATYSoSPBiI9fFFSDnA8QG7e8hf32ykch+UB6u1Y4++8n6vI
LXojj9fTPrABUHSfzZZPPksIxJx4gjpBT8wUxmkBpl8SSQAEZ4xwjFngRgkD2oc4bAADYfIQwM/O
IdekZu++9zsnCLlhX1ub0/QpenGlHgeI3wtjd6sS1SgF4ataU5WUDg72x3ylOKJIGAxwRZJopju7
PQAiO3Byd7pVL4+qms3JKTxtccn8CdiID5OUnCaLYSltoJNPTtBUSzWYJhrEr4WbomkWusK8qCYz
my77Jt9r1wzcTMeWE1V08iLr0rGmM6vqCLdbGyHYVewZcSqHmFaIQ66CmYjckjQQ3d7be2U8ucrn
MFkFJRSR4ANj75a3jTf7ujgxrdKfEc+XQl1C73ePdjGnRZPxiJ0TvVWk3M3DeeeKIw0bR6+7sz9U
MuBifRdqnkF2bCI/ZNf/0KQC0MRZ9kt3RslgcPE5AXFud+Usuzgy3PHljtLiK9U8GgPu0aS2DvXv
2zlp+wG5hhcDIylV5Zxx7LG+xsdDw5U5D1Hy5B6Im9wNLPIceYKncFQUaCrfHm4QmU81lGR7Q9Gz
5q6QIbjDE3wwx/d2/N+qe4FaU9vdkPDNXdvYe6ExlGcIqlQLIvK1b034P+SqQwRdctMUn02a5acJ
EcbFNW/D7W0/I711ozLFame8I2UpMflanH+dJafkKZfx7rVyWOnfApJS4fNDcjZ2syZDOciEqMA7
JF7XOH4ckyQ7k1DhMFUq94EFLUWsyCB2YKGc0kbV8zwA/qzO58FSTbPjzzrweMuys1TIA5HFWoF0
mXOWMHNr8p1AjMnpHnyfhpbhoEGI8ftwI3WYwJFLdjyibA+EewqfSvZSSCbnMRegeFIlTR7wjOpi
7+rrklryT3+AlBxiE6cg1oKZxQcgaU82WhtKGsU6TiR6uiDNr0i3qy9AsqPoa2RAa8mkY5EmeKf+
IRpBKKVDyTNEJtu5a8d8RP4MLo7dc25DHk3509virRBruWDoE2FDZefzvHBQs5T21OYhVovBs3Dp
VnULkbSfpiGk/8jdDLg+pJm8vz75I2dfZGlVZ0woUySkaQ9XTGm8itMp7N4xPKBdFLzCjoEfkE+T
GU0UdSAt6ImHGA3cmN45YKox4fiWvM5h0NT2R2QVMGsTLE1K9dstwLN0oyPc7S92IXsvDnpYmIar
B45BTwlqyF513OhVcwIwqmfPn5Nx4ADAnwEOTVAP7rXaN/brf2hcKcRLsXIhZZvdGgIMpBVSlxhu
kTAMoYAt2lx9cfFoTXeONhmY2CeRUgifSj53QwMtao9VZV0sIEWdh7KDuRpOJgMqqgxX0/YtRa4f
SNhkw0lJhmm7wHUeLwM4c8UBJcBUzVpwv1ufWJbfx1EM1HFBtMG97lMnN7+NDNAYi6dK2Buq3gz5
ha47YhRzFUzTmZ4fuBAWA97LFPSlpHR679vHjhWP4DdhJcsr89Ab5abZjRbqCWm2V9DP2waq3enu
Ebrze30Renl2WO2kbTnXjQvgCE94rYUorAXaneOEH3QC8kBKp587PPQQwctJlW3TLe2YidmTsWmS
aKJ8phJVqOsrN1oCIvNiHFvxVrlGT3gXvfI4n+vGcuifGWQrLla/tg/dW3IXDM7u1MJokSCpRAdA
invIwpO+CAjnpqAbdly8fmfDMrt1uFi9nFYu9RDWKkz07Zxs8S+myisjqSKDtqStWExfWy+QMogy
qdeQX5FKy43f9iTUlOPzvoVM/L9obXd+3/+a8m2/XfwMQ9XGWFUpKS5pGgfA8E9UTE0FBHHsAH9x
FVgARK01SgPldZNoQ3Mhxdf4E2Xn5o2Oqf6DcgY7/nmgoBgm//5jU7EnMz/sjP/UbGnVLu6mXN2d
7xWDpMYzXLSLhdaakHXdEANL8CFCrRggSHIkkW+/Hf1USt9J3DrmXwE/evAtIkMwRjI1y6j8ZGyo
ENbXev7RCzEa48q0g7tkUZ3IFrwEaeRbKGLxwo9X2LwuOT7ZLSr8Unh0uBNDplwDZXDKj3/A6SJu
AKhS765i4DjZkFXef1ZsZqR3hOAWtumZIqwMzCHXVd71dE4Dm2ztNWCI0syTGOvJFBTNtRaHVhWd
zkHVxR6u9evUjcJIjEKg/bvhNcVcz3EPvo8rZZhTJRJnoLKSbuU4wTpV0cHWQhr20okoGf2Leg7S
08WpLht7coffRJ/7kJ4Ui+B2nKM+4UqgdMWV9vTMxTtgkoklg5zMMvxAQId/Cs0A7m9gbSRaITi8
fZs4c9YfqxJQcfspcKmyJN8c5BX5xO6cd6jMKpq/TwidcFN1KJt9piXN8FcTb2v9MreeG/eFsiI1
vDjssgi+XPrEM5+53hIDyPddyJRmcfGdj4JBO90RrUFkxpgOqGDW2iobczdqjC2PLVlPhpvGf3z6
Fp+wcT9fpKPmiUPZo2Y0QcRy6Tr75gEtn7EiKH5C2eSuGyrnZfv6UP+H1MLCS+Buh4fdvKZVYFDn
+F3WPhpOfWuDYQJwJgsmLGsA/aYeaJizm4VFIqzpst4GCb6GT1vBz6u2voLDk19EerUr2bAzeQQm
ux/xUj5kaKVeWfbaPp5UEUVCiVpQFwasXz6jhjQ7s1uhAZPpQqFGKPX3FDoTyIsICh9hScu5p7Qj
DpdtJokdC/cWqcXbTcH/QCTafYfR3LbqORYtkNOGf+FxE9NibCTDOYYvP8QpqCsOTEtTsvd/HMjk
P6ybApPM2sU9gwbPLguf6plgXi8C228pATC5ZFKUKehdwXpAeSwkruwYlO6c0xW1z2nA5/N/us7c
ulkBanXHEIxeAJ40B/CNpG0/2toNMgraBDzRQiu73jbpZXNfaJsqzeJgVvDwKE+23zZqmJW9lDfp
ZVY57SbuQAcGp8HBPPzkNW3s6Zqjhz+42nhSnSF01LN0yF1N+XHSBNz/N/8DrJGZa4ru7OlluQcs
+nORNTs4dxosQsyyF7qTPnomNYdGGptW+ZcUTIOHi57HuCeu8vh81bAvsf4zRGSMHo+sIJ2CCvu1
aYKFDr2pik5Vgf2tHwbckanKb67heMAL5ilutMApJhMIK84CVB9BFFr7mT0vmVjFMrb8h+/BGTLf
k6XbK2hJWRfHRwkcLntacHshmWL+Uza2H9ufzjIkn8UI1xSF9yHBq/uOTLbY9XlBKBqM0C9vIYuA
EbV+Wv/ssFDItfyYUGoVdyfRpsdu0MGShxPb9apc1Y26gou4aXUdNgpr39pTW8I0qaX/o7S21Q6r
mGcyLE2y1A7yTUUYLAHpq8DDkgZlZHp31bEJpG8Nxn4yNx9poyISl868vh9Feo3UiwXwHHtXkRKM
CqSsgT7OIpBsGttjHm0N/YEtoUE5Z8/WW02V0M/pebcSQsuypayB/GoHzqdTeJxY9v/oJiLA+6Ns
6Cjx31O7vJX3aryKXEXVQNTHituXBCM17j9+koxfiC/X/YlpgCplB4Q6t1zVTUfYGNK+6WOrFyEf
svciyskcMZHUges/hNeh07mlxALbjkW/CmO6x6Vtrt/JpuHRtGQM5MKguxX9mzfzcAe4xnDlUz7J
Fl3AbKfjNmO9di4E2CJS9L2m3iX1POkIZ7vKQDi7Ronm2XtK6B1uzf3qsopvqzogKBzhcNwYpu6A
Z9tbH8EFIfKNoVTbaKuIMvsZOtFwcZ4CD9+4GhNAb2v2UWBZwCswUqzgCRFvMi2w7eEHNDQpBaFF
tRTgUmeKA5l10XBvx6OOyifz13hXOCUuCmWyx1CvLbqa+4gr3k8CCNclKy7hl5hq0ww/UPSFaK5B
/upcOzsQwDLO78RCklG669ZXsukdNiejRltOomEQeRoSYY/EarYk9+3ZKLp+GsCfvNhtSwPcRAbL
kOddcR2DfBYsJuTGrYdHS30XdUN8lXcK8KGzpLeDVDIOGcebUcbpVvt1pg4QxZfMzTfU96+OEl30
ZE8ezWu0b6A8NB+1EksjGDMz31M7M9wV4cdJmTs8gAmidTuo8vvdQOT56tvMT2/DmzEh79PEAL19
TidE/c5YrJj4hhu89qGVRp0O9TsG21Yhhz1s+pfWkq/D6tMtfCnVlvxrwGWJp1KQfwTb3FaWZU7i
AUybg3LShFO+VKyS3+MWfx07IePC646oVOI6rzywlc0Vm9kNzYRJijLpG7iiLx+laqYkS2h2Vdfj
7xUqTW+9S658YffiW6FR9Kymr425DAcsQeQkwFLDquy38tNRTnRrG1F0vgDwrQ35oDxZ6zDToQQh
HxV4axzwKh+03hBb1UuJnqM2w6HO7P3U5oqj2s/FVDeWWXgA6U9styVPVcDawg4tHGswkl/SYq+I
c8k8vd+/T63K1MyNSgDP70IaMxN05NMb7+i4S1TqDR4tTn99y1o1FCvH/5mvd2GGAe1bUgot4hW7
Q0gViwQVWaA5fHMBoYTpfIH7WyuXqhT0jx0YXcZaexnn6LmXTdigtA2Kg1eSwHPrhr5ZeeKb1sTj
K1bs92Eb7pXbCEZeqUZM5fAU+Fknu0GtQCpMCyECEj6c1RmQ7NLPFuomspGVaEw6MyX3ApNoMmEm
q+uaReCliDsVrQe7JPD4CX7YoQ4oyxOxSgP3qEhKTdAA8A7Y0B7htTNZdWITDuh4OXx4JUuZQ09D
/k4WhYMVku7P/ojgBLGECItWDpAk4Du8jLNK4lONNPE9XrE+GC6D4hyxMyUacyBA60VGXx2Zk4S0
tn3IvAiQHbHnH60OI6bLX1Y4rrBjm3Tj79WDoA+Am4WsbXQLPmamCnxphiUvmttcAACFx+L9OkAJ
SEIWpmV3YUi8aB+X8T6yT4sqbw+T+3+WFfmUj61V0CZqcpr7Jj6BFPLMIZeH/JNz5mSMiB6ll/La
NYMyoRVzidPrQbapt5b8GVtxRzRq99V9b2PsASCSWJFwJ2K3j8s5UBbP1Jh4V+edfIw1zH9mzeZU
cKZgAsunjD12OBBWokasv7AN81dzLQVjGm2tVuvPXWEUFHJ0lTBMA5F2GK3suCwoH6e9K9stpRL7
REoAu8ntJfmFtG11uT8THXd2LJs++WKRJoLF3NZQjWCF5O+kYgL1z+1Yc6tr5w2oV1N1Hu59Vb7K
v1owuxN6XvY7C+UucDtm6u7cvQ7Xip3IX0BCLZ8PPhQ0F9/F+V2rL9F7CKvR24zfO3HtiHGbY1Zd
uslIw+m77TRCZDTiIe8spqTLbOylSNfdGc3nS0LIjpi79pm5CMtRRzV9f8rY6lTFNVVJsr8ruKzz
75gBxwroVQFbG+zpr8wI9/b+RrKndGOxcUC00M7kgroeEJpIRBhjsJj9YIAoGE6eLVtoPPtMep/F
p66sxdgWOa3OZL2zK60mNW1jp8SJ+hfow6eMAe8aMAeO5gS4q6dQasC63qqifWLwgf8I+eBPU0eZ
b+oPbXSCNGxC9S3mHKyu0JwrjbLDkw4NDds5A7Y8atEjoGZc8XBAPqk4To3FR1HPkiKah+tpiMbI
nySmd3Sa4uj4vHys0g5E6M0MfflSRAfkogUVhcl04BSLg6Obfhv+egGioqfGDS14NSpARn1NJZ49
/xTTjHGDZ1QiOyAovD5olRCskqTjdRGhY1qSRnRz5JyORMV4wf4jQWfQ11y6wQ0r7QMR2TrwSkyZ
9SU9KJ50VVojmnrIb9ZvcMoDb6Rhpb3BlKOLsh6j/oSSquSrJwvn4AiYJG1Yue4qBAF6F8Cx7GLA
QYg82E+vI42rJPxM/J5B4ooqcRpa2lFzv0Djn0+NaCo0JQvLNHt8pdJKVSmXWFtm7O71dBSbMBwu
N22M8l85DyHI1vlQwiUI3vU995CJsZWRTJYgVYvHg81jo9x0JRX1Ue6YxbA4hc5rElpRBSv1kSYJ
lS8eDbYuIjegUEEsCMc0pDB2L/1YHhRU+niVE/9XrPP3v1OPdEFhH7bxEBImLTAxuVvZflonL4v6
/NoL37MgcnPoauCXbE+VkWGeRYFUOEbO4bzPRXpZS2En26wVJ6i1EMH35XGQWMhLnCgVcAoaL0Vi
p9PvwPmFVyaUT54HgIhKWGBilrmSb16rN+/OShDB6sjwcP4ecqU24xLpuZtxKfqm5tujPDidEwLt
BdfBTlSzHTFkpQayh8eSv8zS1j9m/oSYpmQyjGY3TFIGmDSL7zCWNTFvIDf36x6PjoCn2jea3mYU
Fr9YsnzZT7f1oVN1+ydO0RZOaZBAEKpHdkwBpIs1dIiJ9fmw4AM8DXS6eCsvU1rrwxHZyoz/eSvE
lmGK8cQkC03g7qaVbput4Z3ox/o8LIIIWW1Ur9C1adI+Y/8GkE77m4WvF9D7CUxWMMpSqTpMHLPB
EcDunkdge4F885q49gxqtvVAwTYKtJlZZ6kV30aIcbLznHW+K5RCr+d/NOhr+lA+IBkiTE/+9/Mq
Ov+mlmM8jV8MnI7diX7ahoN2cJCmqkrk5bcT0ECO4YPUpyLQAokuzMJih0xRRhtK1uEzzHxNblMq
YNNLEfQghTjxl1lDI8m4NN4Tm6UFM0h8UK+tdYUXqSjmiHwbck7JlVxO9ZPzIK57MQZNsTMpM2kp
K7rFEvfOoiQbHTxUjqHLM2iZgjs3CUHYsCDPovFuiCl1PlJUOYQS9RXqFMZsRIk4zPT3VdJ3CUWD
bnhzzM0HWzKV9ZHhknEEF/Rbca80ASGbqCKATAUm+GId96fNHXJq3fedJq193HVxOyCPWkiIPzaj
VBzwGEBVtgm3sw6zDsIJ1qwN39xQTs4pKsKpWxjp34WFvJPELWILlKphxFcRaDt2GmzcV8Sl/4O4
3SCeE5fBxkmQN9Q/6Tq0tCelItnqFP+bycm59GhjlAR6/Wa5U3aXfC2OjH6f4HrERdvdHXqstxPE
kutOgM1to7jYgbYxWbmpPjWvKJrFek5nyC8cCNb2Q5FpUyBQeNynRjideYhgZpwWFlERrERApl9j
DrkUVDYLh1l931x65mlDpDvXD4nw9QGB+MvQJJBY35Ar3P54RGHXLr6UYYQRrehedM+s8m7fAbx3
yqeRLzOOkez1aQQHG7mCxsNBxfpZKGiIe6AQ3WD6jIkIwRJWjSw6/5wtUr2cBtoJ7Q+u9NlylNWt
YuEVjbwG16m0Rng7+53YRE9m9QGZjddWDhKapLtstsfEslOYu/5XbGYGKAoYHFfgVGRJG3RNANrS
r6IedD9B5C63AnpKtQqdlWEuj8XwqzK0+p9paIGn7NQtGZd8/SEJBUucif32tP4WbWSXw8TA1k43
XFPtkEP4KFpY8Gh42eV5O9d4g292lGh537KR9MEzD+bKKTj14JNy0ihxZBGMSDl4+/sH48Dvpkym
CARHFAPZ2c1IaxUA6WkHvpc13JpVIrFsfmwPeHS5lFdXzjU5ns3Dp/JnuywWDXMLwVjmdvwEUnCF
eEFQhb9oJxr9pDtVl0YsbF89IntlbeUhXXlBmVj7425oYbn6eKiOe4ZiIDl2TKftWZXtklyZyaFp
97nGJEGKu61w75l4chXDkJDUcTC0WEsK+0QGys+3MC5+F/kKnIuL41635B5zFoDjO4RMILr1/gLV
HvB/8FhQ9if3vHzo/I40ux2YYSaDJUAZ4DH0giaiYaAjpHG+ANFMrBzNWbOxWQYuRz2aURQmn/Ga
qP3lKDk/p1QhcOeIuyiQtGjWI4ezWsr2er50Ebe8S9xqRfOkqNb0WUWUU2jXDf0BXiLxAgu2O6Rg
U/Nuw0NCd+J0poqtxzJOuV0E+dKtz2aGLEMXqbrB5NWHtAeTrMpxCt2JexZwfEIzlfhIs4eYDJFA
mErg5LFNKRbwGlISPcgblGoevBgWwgOszb/Rgge8q/Kpl/c/Ar7tGwNbaUyWyqMllxDUx+WxUVG2
KptxrZ6KjRdApMcxvokGot1Q/XOjppWadjVrW3BpqdEt+8UXcmVtLPkEL5C7Kikv+1ttOcVFPcnD
bzvE4I3Dp3RhJYSWunp/tu541BazUJ1FssRC1tUPhQXjaKALJzLAGYTCrVZkiVtEyDQ4Nz4tgKxm
2bIEAv+3GRLwRpOpWR25ei5OWU19VCaCGI5QI8o0gTyMZ6QsK6L79NeyPdDv/1UEE1ErxI3H4MIa
Lm+sikB0xcX7tqWeFTnQAROX4m5dK46MEmOlR3LQKuOwJ78Z4vXk0DzS30jucP8vc5rNhgw7dO+7
2SbGrDN7jU1/eS1/UeFUHYdRWLuKEX8DU9o+6eevqqNaH1qgv5cPOSrkjgJ0bcz+TGJB7KpU02Mt
0X57tGl13czxlF3OQekk4sFmIIFfe7z+9VFb4FmDK+Ofc5TiZgt9rZvodR+dVC77Ce0f8D8ZwK1g
AaF4sa8sq2fEiAt0KBSpM143fJNaJBvTqtxMYyPoSCIjkN08eeLzL8DuCvNz0r832t0NRc6gWEmk
6H7kmmhPJZ01xWayiHV7j82CEgTzQYHKEAOPpnQc1PM/06gpYkjIloMYDYq07l03SZ3Ql1iZZFfg
A/NBZ5liyIdfUcqUaIhqIA8iW7a+PbWyZ2BmlRh2+UAe0rEaOSidSy1tKSlGbkR0zWwocmcbG4up
nm4fJ7Es1ZyPRkuIB9NZFL+447RJZ/sHEuCt/ALYKzPrS0J3PUzQe9zrUR14Dfi5EDFwEWFZI46z
BM5wvn8upEpYIRjwH9nrcSpKM4gwp2obodm5VO5surzEqmAvScsgQ6AQLzOiWm2qHe35jOMjTUzZ
Uo5Ww612HL2sfq4pGyyaRlmUEjEJByXs5V6z6hAdICWG8B3SicBzwam6P5GCYMCkqG7KGqYiEqga
IMK7D5+o9h7izio7mwJN8zdPJ48hqXu31kVv5Tp87S2bR53lOGlVzidotwSXIvcdJmpzmuIo5+G1
wBBwNxIZdLz3P2v7HyWIphHyUIzE1K5SYpnDylCVUCBh9KG+qpPtZ5JjxrZzPu1YaBe3gn+pyhJz
/wKksO1FB7yk1O34KzFBD5DAtbJGtNGyyzVyoMTgPQ7V8tjfpAaMgrZsxeiXMU/cK6veYCuIoj2J
iVaLRvBqvTWdJ4chHKUjJ4qsSLMZ2c4z1Qqwym3AF3QZCp5kHBr+wTEZOJWvOW7nx/4hpZN31Y7B
Q0rbGSSPm0qlR5y5B4qOI7gnMeNLAR3saCGdg7p5+DG1jhE1abbc8IXIoWCweNrMNX5T2KhJxxGn
/BJqwPm+cXs541PmFhbN41bQ2ieHU1bIF6ucKvnwXyjYF2icU5KqXTlqWTLc00WwomtiLwmHpaCv
Gl6PC8Enao95MO3dxflewo/75bkv8rxNAohjECRF7Ds3Sm8CCwKSzciDY5P33yji3F7aKF3cVOMz
mIaOIYA8+sz7hwYX7Pkh4JA7R6HcWntTG579wulXNbUtCYoNV15h65BjOC9t6QDmVuR1voDl5EA0
5gyQoBk1miQSdMejWRC1PXGizcR+vrLFoacVbhFkFX8scYCMvrXWSXgRWOK9Rs5pMwcQLIVGQbMu
ERA4K6JBBLnJd3zHt5TFFvMZIyP+b8JjjEupZ7eWU3UsC16XfhNAG41tBfyHZfeC9KMHn+mBdj5w
c9UNH2opqzWWvO5BXVphxcXx1uvO6r94VwYMRLUMvfUO6c+yVyrIERvne3N3DrDuqurBBqNs6CeG
pRYAkQFl2erQpZQ5ws7ligS6ecS/IsbtO47AtJHhKoza0GvzHRjSaz7ZpIJQ0zefETEubJ1w9FP0
IXo768/ABQe3tOTlI2gLfhOJ51VcKJ9DXzWrNKTc9inP1d9SBXtyVnKp3NsB4tnSo+jwhf48HAVx
BM8ueMFy+BVRvopo/P++TXIpKVnAvYCINCvBObJBx/yQ1YEVGd9jcaVGjCOGFhgF7dFIzdG+E3Vp
vywudk4ECHHQ7WPEi/QQCn30FtjF/u+BFJ5WqvZdYo7LDXcq2o8p9e4XDG6jTfAUyZQRdwX+VoE6
jAZH+w2qVEGwDizYWZIlvgkWp07D3CgQall8tpskN31xFLVRJAiS4rod0XqN27JbSu9WFNFHN6Q2
8jQz+FFFMssxmq3qoXEMVy3Ic1Ji/zY8ZuNc9Oa4dThDcFGxIrRDYMX/BhsLj7pTuNgLYfGJPYQA
qzKGrM+HPk6xI0PqPe+F5Dx6lekFe7oWdDdna6BHJ66vEBgu9upPWC7i+9ih5hsX2OuENjegKk/k
0bZRzkOl7up8Rpun+odkzJc+wC9WGZWRFgy8q2+PfULtBDWbHWzvJ+HCRYeJuyL5v62uFOsWcex2
5nDGYB3X8myVbKD6Hfu3stBAXSIu2rPYC1Rz+L//1cDgfwt+VjBzqj1+JLuT6aStQYOn+au9inqA
byLEHSDMJvf/ssZyX2yo7iAPdimItA6o2seyjdYRJlWmSnw3Nz0s11xGDEDheve3dOLMfhkey1Do
Ze3wpDV/H4wetEjK4scURMFdgjGpkIlfHcJUw2PJGwinpNP+oDg5rCxwnfxrME6vZXOtZKQwzu/O
pd7sMl5BWgnLvDcC2WdKOz+UCQNAXPLlEjccJHfNGT27eW7Y+ZqBkunh5qRC1Qa1VMWgnYO3JbWq
36TyWCwdWifTgGJnxhl5nFXO3ZyKCd07BtWsQX7xK+XCdJfx2WkDNm50BFoPgx65bh8ZOpG2Eufo
rnL4EXobd2w04xWCPVUyd5fTsgJcWdP2FQ9FDsAStDsKwe2aj/gcjOtWsMZZVNO01wkmbWXvqbMM
b2+iXsYGBx4U36Nq0SQQ6ia8VS2XH2WRZu62bht5qV1b8z7H/bI5EOLHPqHPHKdSBdsvvOcmDRz/
vooK4OMzuFo5Fj03jDCt/vHGoxGzMp5uG8zoegpWXewWd/IGuoj4IMItmZ4P8y1D5SwTEy75VhIO
VvZe7utjx8oVGgQU4AWtDZ32VVfZvWkK5zzmwuO9pLjk36OC3XNzi4vSppRrAASVtfzaLU5b+22V
ibE/iLyN+G7w+6VNy+iG2h0miiaUiKVaIf/EZu53IbwDZl+j/B6rq9hpejzcgMCr1iTwD9SNkxky
At2Ylum9sU28Lf1vuRm8z0eNd1QLg54Hj9VTj30Cy/MjdBXK+eKCvENReCDWNp5sIn88+m9Xc5xQ
3kkQAbbd85vIWWnZ8S/eIeLg/nz1JNWOKRRk9/d7AXPRmecLZj/V97TjC06t78HbFsVLJ83SGQhE
oliO8JBz+lTP2Tirw0VqMCLcZmZ9rVCY9BHNowDZ2WvCyXta+c9he6w4X7mLU6373qgPem5SSpck
0nP1YahUSnAlGEF936J/ihkdIaVGzq0Hw1eYa0JnckOCiNKjobsRRb3u9ePi1l87tBH4XhDpxS1M
VIDLZNox1zhOtw1VKVwsPKcdHp8vXCKeT3wzeKnM3GwTcDkAonyjmZGO241KOhfx2Dc/2o1rKD0F
gwFsojaMEBB3SbaT3Psa+TICA6N5Ni5NESv4qtdnA20krFL/JZ3CMD4l6KJB+CLBLqYogKoXi757
Igw+t4VubMAABoS0cJ7HwxJYXLgsU+ZEy6rk00/XC0vlNG9kH0UXguQylwNUAnZqHJYe5C0+gQ5T
mtCMm3vq77MgCHE5ZVPZkA4jkk25XY8hqIW8PUc9bUft7KQzUdhsTadl+Y2g5JQIXBZhR2TKx1El
xUwU1HYBAZs1KoeRUDbTikBV/IwwY/VamG0GqwsAHOKr9ZIRye6A/WwguirEk5MwA9NLSWxFfXND
cdM438Pg1M/U9r2lbUudOv1u7cuIFZg4FBzXASPL6YvXN4hyR8dhvNYxiByE0ksLJvHc9BowsDc0
VGxS1mBTMk+SuC4biu4VG6cL7zM5VXYCChEnMk1TgwMpwg2zOj91oDoWhS5JWA91AR8kd3OpG58k
4RIVekxOhSWTfBjU87tBwHGic6nWcTihHB8W1ThvsFe0euSpqcfk7NdbhBgSCl+3bwj2SYTGgIUK
eDxv+56fDsawaWKRkF9oxNv83f9TYbJokxPe/SJQy2VnTvtd5nn4v81YKwa1oOGsKQe9aHt6aJ5n
dqMnbSZceShcurzK/2Ze96nEAk2uwnkOq+A6vB1Pxg42VWDftkOMQAK8CAtS6gqyHyqHT0arjxnJ
DDdllwj2XwvPPuAHqYiH0sQAvUsXHPT3JmY/hqODkAz7Ju0hg2p8uY9oKlC92Enf7IAKWCOoosFP
O9E3LwX8dRJcxNV5I6tOkJqe0/VEkQ1O5ZxIHwFlMtDBTrdxAAZxrhWV2eqgdhiZNbPryowCl+SY
/ajGmP9amzlNpu5BuPp1aDvEoxOUP9rEY7J7DhCveF+w2+lPa7axUGRwnxphc6pU8/g8D0Ub4orZ
85ldyCeDrxS38Vg1TeMnSI+YViVPdfnFBGLQ1+AoFWgAAUSVsLli9T7XJ2D8whgdCvYtz3SoTYpF
D2EagIGcaXUsvzMtte91KsVhAS560fPzuKG4RURYWShkoipUSo3SJCp7qwEUEcJd0hm7gTvF2DqA
v+kKrrCRxgH6SUwUELn6gDLVNkJmfKuE3BZ2EMwE2blmSEoRQY7qMZBiYSRflKarfnwQAnYTNl7z
K0+PKH3phPEceQRoKuqcFq6pzR358a9L7e/9QFrpsC4KFpNViAKio+c2XYvW6q+9LZkm4WO37BFY
k/+/Ur91UDcP6YWqujYZ7Hy6I6aL96iNIcHY3a4PDYFL6iTV1SQsxqly1+9998GBCR9IQ0WnFhLL
xiHloNKvwTXhSjYiF037mpLINciPECo8XkVqgbdRtHllnSQbuhiGLMZVnD+JJTdD2OFww0ca6ekM
mpR2zIiORiLH124lhJk721auVYbtv3+wKfvh6BkDK4Uw71HiBpWn4BVc/BoEi/cDPIhIRNZaJh+v
xBbG3fEZ/hvR2BEIqGIIaOb6Pqw2mlgk5xfk3SHZfsaXClHzTI8NO2J130Kk1NCI7ejeg5cIickb
A3mjh33/0SDY1wwYbPGAdpv12uBJDrbGWRccFXFeNyrtE6UGkvbwpWRkX4G+v6SPdET64Mxbbtd1
x9uozAR22OCVnR9BCDywNgv4uhrdD3JR4HfffTA9XNlVEIcqyW80042M7deUSnRj2LyJBkubYeXA
++1g1/vHH0jQ+OHRgxZua6G+oGdCdMd4B9V+L3o3v9wLbGfH4EzIZdLrvnvznpWyfirt5E/Usc8D
l8zpz1j/qxjIlNWATa9EYyECxIoMFbM1yz9KpVAWZsABCC+ArSEd+L6A6xMQVITWVRrWbz0xfX2/
HoHtTQ1P7IjohAvvu80wcNj4P70Bymlncb24fimwaTKUrFuNRu1RfR5wmnm3j93+JEreMNAeDly6
MuGsKv00e0d2OO3UpkdfT98theVhkZ/KXnJFy7ZCErmE6rEODftLySkSwKTVZDg/Qv+ZEtJlZwL7
PCTVODksqEU8fnxBbGoWctoeAXYmuF3INHfsA4ymjXSmd79hSi6r1GG37KlzNQo/UUuhonYKDaCn
yrrQkZcBk9edUhqBBNTvSCzzHS0f2XulYCvDxspnMk0fUD+7N317cOVcnRddZ9hMRRBkCXE2ppV6
vs8O1qUMt2ba1pJGBMl+6GZXWkjBlyvOFiQcKDx5WyawHYLP6Ur4rk63z9IVmHQfOKubLeSDsdg0
UT2ZQVo4bQVOvDfMzY34pKvCdLI05FqbY97WVWlENh2X0YoSHlQX5pkaMQHUG5CBQjv7hh5GUt5k
NEsA3M9Hm6DdGTShaURMJQBi56KHJZjtqAv5Te7EM5k/1zJjxCd2G1tM5+W5ua4K8QbVrb5B2ZbS
0e+TnXEA/pqlVs36JSBCJVyTtXQK+6Fbkp4+jCxApu4Ok20SDzZs7pHEEbwcxkM/+bWT9hYUbgrY
+RPghfidLzvMctz+5fjMSL3aM5Lc0nKWyU1Bjwj4vAb9G3uBfCAnXqRBms9MNFsVmKDk9AHeCGN+
aPhdltvEbEfzvV1lT2narpOIZTjGv9+53LsZ4KWaqHKCMCxxThtNLI3pKva0bXB1gdk/Yt9RJAye
gYvsRrjzhbhP6pKo7ouO4Ju+JeCvOQN7US5hGlhpFw5vq+eXHEn3XYB+vfAV+Gn8ybdRXxDcfeyX
SDPThce+bEpNW00M4sMkFB9lhmfnFZ+kMuj99piOP9tbpeyVXeieng/sX0c5X+Y3rxFvjF8y+kZw
Lblyd1kgBvsb0jGG94SHg4MxtFcIHjVbenCvBzqV8lG7/WsGbLYMmTGX2FNtak/MryoA1J/znSsn
br4O3KDOgV0UEEnTw2xZ60uOyGJpvclunb6SdIy0ZId9oE/3fqPjZPlzVTNkqE1d2CmhzV/gr6+r
nwyhLPbGPtPdHHqk0nvAt2VxMbYbnIufMNE3coTKLcyys594y8SQ+Ehe+vP5+qIhQfiiB2EUOl8N
e3I+ARCxYyWgNPyfQeXSRWQJ/qsdFpRL3o0e9/xL+vMCIY2byPjoKIW2YrS5ybh5EPDhe8X9rX/r
tXR+dbmYFghpGqHCYopUobq8q+BcZwzNQIC1U8q3E7M+bK5T6g3TxogsjByH5n+iBtbVshJ+BPHM
0pfVdSm9ESoGBL3pmrUPzHdwxkJ+JvwTdH/fN8FEvcr2XjB2ZvN78W//WxtVJMhktowUajsW3PXq
cwD2Q9oyoCXFtGSeh8e3gwT1wfi554DnLZHstD8+tPcJSpMjNI8+ILU83DAzjFfz0DUgCbi/sZpG
AY7LHpVnx9pXp5q5oEKWx+fDKwsl7AMFlFhtOzDnJES3x9p+hqdRgr5yPRME1TTWtUJMfTUlAGXV
s3E6kR7z3w2Own07iu+S4EDUUOf51aN5qVUrY5vvwwBQRsUfcQjJOQbKWKz60Ms8iPt8uNw18EOi
XA42XrcIf1laDob6AKBC7kSI/aIoVP0zCvrxEBF4ANpwlhhR2HBYnoOaL4+Qe3R+Sw0HLKTT0dkP
2LSkVzgJdb51m6PMa3CB8saXXLrE+zmiZVoobAUXFJkY/sK73SNtS1cfmdnsLqsoklHGeRAUnFR1
MusTHjDX98xy3avXuEA15iF5eDBxYbjA8ZLutUBwSdtz0i3oJf7Mxn062Llla1tOOpdN2GPQGfHm
efc/DMjdY+VqEtb+BYg6GfUA2kLhVdzCrYHCn3J4VUENXg1leH/rFpfSMe42zPcTFeg+8m721WTU
uFXoxdaY/vyhB6bAHYzMfEVSZjCms4VB2QbP/3REySddYGNXzJVUzZeZkz+66H1J+3RrSbra5riX
0RRFW5wpxM/uL1U9Ugvit5VNWYsIICcU9/u6ubaTpwthuYNgUjI1Kp7A9ZaeeRD/G+dKCN1DQsRc
5x+zAz1e/+Xi0C+/Jnk9xS4/Pyq8wQsc9O1WZKGW0ZMqyYvgYUOVlPpz7X3ed9qG2ICQuyGT79UE
zRS8q0T7J8d2UA+M4EugL1KAma/J9pRyUeJEGvxOCnq1G/cx48QRxHdBLcrJ3ylbUOh7Q1zSl0Y9
QB/1gRMkjg9plw0AifRN9MeWXRi9mYWEGEbDoeJ0hi1y/bK6GGuFNdXf0TV0EA2szMM7zjNui2J4
4xATN0I/JObwAKC31tZxjdSdEIgM2oDn5qiOBMJUbabNaVW4I3ZXF+QZlpVzfFCX6yG1swX8mtm0
g+lJJh43bAfTvTO0OaZrv0sQ+23UIXlLgBOcWetrsPeYsRWgZm544Kh/nvGuAWfsXxEZjLgHMLAD
cT9cPAUIvW1XbCKCI2sDxm+p9skwGe5Q4wgFdKDt8JrCFIc4QawRQ9sumBROcFv5wAf89Q682BSJ
pguMen9OwN5XsPsAwWo4XAkVFrr4rdn8D45gGLyTZAgdQDtuAvzyjp8uFPFPYWBa+OtDPS7/MJNp
RS0aFS/X7Hlwg3ld1Uh6qEkqtjQnzVhNtKdQmzJXaz2YnICAIRPaUxdEAGH5gdy9NgBT1Xt4jxda
T9VHPf/GLkv0eArjIfyns40I/8ygcyUw54l2o3pF3SoYdhnu2E7izk76tf/81fPaek7Zxuw4W9WN
8inokB1DbZXHcWqbw7krs/vbTiK1ygYHcucPQlm78JDmnTXuyUPwgRaGOM4kWULdFJAM3vmzY36Q
EjBkTo9MD5JSKC+sIPdoqTL0KmsDcFQ0wWPvJuNyocNkBkR5GbhxLVXAqY7qCINZyzMssyW/Ibq/
9HFe3TJ3T/iIiT/OySQmn6ALDgjrAfQ3zjAsA4a7xsgaGYyhVGs8J1aQVvfQro3oj8NEkGwOt9T/
tpnR00Dl2gOUeGKrIFdGa5UqBAByHq07j7/+aGkVTk1ekDTx2/Kwgnu9WZdoRbGRd9Pyz4xWwOSA
GWhVUyvIYlmH8pZRO2R8/EZEZ1a2R1fPwqs3QwAyVJc5Tblp+Z39HIGFlCeA4tKsmdEwHrJVF2zQ
Z8jlrvSeThQGSHFy25RHk7GpTCzcsXbTTO4wdb0cktNzQyQCzIC4PB3ab5+YOcZsmkEgxzWEXrpQ
XCtB/QZEDmJLcm3V4eHdD3OKGtrSN7NqUtnljHNm9LH3rDPg+IFMTXX3+QjlGm5ununNKFAQul/a
Icu7lnVX7SGbw6thJw5VJvFKAAJAbuWVJXyqIoEek4pItNUMOPdWeKbywOFqxVZfWQbMMoYMoTcU
XUI2DxL9IRgaL0ATT+lm5nUPaJjusCfE7vgWwRRk2cJWx7iULQ/ysnrTcJ8JCGxCE1xxCLVj3b0r
+teognI0bxMwRx8Fz2SQ7SeMu2D/7IjtPHqFTYG6Stng0FIBgJpnTrOZbSGeyHjhVZ4SavQ6Nlmy
A1cooPG4hGwge/qL4FKs/GruAzppNeCRlEbTbrUdYMGP04s4YNRO3FqO/Mx4eqc/HItoHSFZCst5
BEARFMgkyaNAG2w/Y9ii8sH+CboUttrKF83uCNciinol0C3+ahGj+cyRcYBwZOFGXza58/9Kb/CQ
drJek4npi5C/DzACFBAL6jCJOjN/mC3/Z/GWdpiKEpF4yyaHXMMV7dApDKxwO//8V0cRUSiezTQk
99Ak5nGQN7i4ufpk3LaJXlNCtkFTaBArD1vSkT1VMmG4IvBUdan8xDXxw+QhdSVwXJiKtpRb1rXm
Lo/nw5UtUHXR4E29+/HKPWDF7CnEdRrb8r2ZwP+FdAAK7vwzOD1REPSfdfXnUZvSDH7B3uJneX5P
YIf6DRGX0X4ctbhyDayJgnzIou3PVqGItKNY1cRgkKwmd1bwsp9TQkLj4kK2GTlw41Zj+IXczD8f
vdjEpBiALpclOiGwiSeCk7WjaSshK40Rb2YXLBXEibOywDse9skgkGu5rB7UGXP32SbFCH1hoknl
6DUsJUikI4Eb/GuzFnmXDwRQig06IjoA8SC1BPrqfe55WFj3oiNJ1ODdOsth3+XpVCrpS0EHrIEk
UQoQwpcAM66JDBFlxWaMug1zFT3VURGp04tZ2/rUxHhD5OWd3XFyrBMmt4AOtHYxWYJI477w/ufg
nxJRwPP5jTcjLtY/GnQQoczvNxPg+OMxwbmgLwkwi+96jkSxHupDuSokjvvxfCIIq0g3E0ThnRLQ
zdackiJ0o4WgqxuOREsUH1SaIW25pINbFRYVRco44BiQsmEo6BKRoZHw16brPi5aEugE4an+NfTx
vDNyVnAQCqsZDRvEcMjqgP/yRTWjzyMIw4VIifWh5dF4TIW6pkQwDdLi4bXfBTV39HYyJdViSgJP
2Gj/YbG6m1VhFTT1dnXHGfDEcvXxT1AVWdF/HbDkCEloZBhEOTBmYgW92ypdlzRl0jWmNYcIYWBs
5D7unM6mu5IY6hqG6fZ23DHxc4eTg4hErUohpWCjFHFCO6UJvbyUMQUCnkJDPVKo7kPBWUc4Djnc
Zlek9SZMHBe2sIXSe//1t/X9jXJEu6YDRgSiZnONno3EFxD5n9S075COX//JQUhQLyZOLTpObC0S
Qy6HSh+CDZXrFzBlO3D3tFOuoPHXgVDgui/0fPCIuKqVlCxEQs0TxJmMlLkTEj6qtM+0hXkD7Yo7
tl++7Ahxv/U+HswAiTM9wciqYbAK9tyRTCZLdiJWizQNbSdjZuNdHWp2u3dXACNerudnWgyjcZbD
mWOOJBcvIHJaFA7CmfPxajKDGb0LEZeqfJHQOugYxUxt78ZzrHWg/kQWN3R/NONYls0y0neLJvOG
P8/eg2Q1I2LKRIq383K+iDTcWfOxUUdGZJQMqKP3081V6qYOrQQQyVjc6uq84631X8rni98MWPkt
hrFWK8QgF+OERreRTXWJyBAq3iy11G4tgLz8W2vVHsY5gl0O7kb+j8Ko/jeihTHO/pF7Q/LthXkP
dvtIdMe4WrMxK9TyR0h2YVfF1mjj7k5ICyZfBtzvUX0DevYLxnCudntkbuvjLWuOpl0u4o63xdrY
kqR7nojXCh+EbhCess8u6n56htKUT+be+bAnx/NUoH5oglpiC9SOubE9mCREGON8DU64Mk4cKquZ
T593OR2pW2rxdWdFIEJ8fVEWFCrtT85RFHXyPCy+95JiOkNS4l1Fvdxcat32XBwWUvWBK+ImERNe
fy3raulX+B4+Pky7XJpWfvJwzT9Zb8WULYhWMNqVJXqRsaApiMIN99GAfWic35gUyjxYYZFvgGPi
8+aJQoJONAsBVzGeU2FEzkudecXVpDCcUYNiJ7LM0/U4ADfogWDa6Vv1MyLkvOjrecB85sM7FDmL
dngJiEG4hFghnl9zZxF1ebprVmPq1f54OJE7vv5CYbVvLgKl5QNBfYgh9YFs3zVzM9z3OecoTe+O
XKWK84WoU6aC26JA06MSz47T1MJjSpUXqhS4IPkJnVW8xD+lt7KnAuAh+b+L1m4VvPtM0El9j1fu
x/Vo8TVMhlYTAge3sJl/BgUxg/GssfrM+spHZH2+WQMLDvOvAe62ixRjH2tfy0xZDev9SzRWzGxQ
roTg0wC3Ao/coYdwSYdH842ZOzScvLoH1JlnrPBwxdQAE/WTZg6dXcOxC6FJ9gj+ywO0sowOLx7I
QmwoLZcAgZDklGGitL685nu5YRFizE7HpzOpE7kBg3vBCP350WXmkMupyj/doA0ggzXklBh1KJ3n
8ssKtxF/rNbnf5CrytkbRpC+Nco9ttrDKUunnaBt/oLpvdYbC4kIAn/ex2hmnoPqKmE3yU+K+dgC
H3hxD6cqk8QyXMq8VDd4LccdtZOO4BKeENbvEPLy0fYcSxesf3dzIcxDPDwh3r6jMThZpSAZb+EO
N5H+lUs931q1cFGTabddAWgSwAyzjs/NV+xjM93g4IismUnBaqn5PsLS8dakpoDJXn87JTz14rkk
2c6WT2LaI7yaIPPKhopjTc6uU0grhRDofHNs/AOiLc2WQfQTgNWnB2NtrFNKYPSOeed9ENm2SCzp
ojuHBu4diRQUaMeFYm6M7PdZkYgznfBq7mmjMVPSAnybXdDNwuI+YJeDKxUvd8Uj08ICFnQ+14in
PpWa7gbINXD/0Ig8n3XR7fLbN6xtBgqD+kMeukjW/89qdNjtjc175XavPTssPYCrzxfVZxinrcvm
yfCMA6gtLQUuMxgLvNPvc2BU2ooKkTH5IYJlY6bjGiYQ2nl2I3+Rr+11cdLaGu/WMZ5Cg8YJjoaC
k1csQgDyqJP6PYhSrKcBVLlZ+yUmbCjamzIIEAFuQRauyEt5sXVs+XXUvCIAt+3HECqW1nCoUXaK
GgawH0nNAUaFf+Jg2ToxA6A1EiTf+9VmaFu65ayoTRX9y5NHbZa/HmF1+NugS3Dt2SkzoT+hMcIc
koXw6RIQ2hUsFpwkK1J9onIlhlTQYmCnXwuG12/aZaUnEzS4G+2/yUsLvtANxdj8HEaKS4JQhFZP
owRqCBkxF0EBFc0kQVVzrPAGFdwm61tSic87XAKUCBKRpJ/qsAN5VC5qAv3DM1ZV/in9oTlmzu3F
UISjPT8VNvo+lbrSYAjo9lNJU1h9RtTpqctjvDG495nrCMPgAFT4dKh6PXNMiH1yDcw53RmsGbMV
tkh3NW+9/UrfCWLVrHgW5WHUahO4BQkOVUPqoaSvVt7nkdNlutqgnOvq+bmJcR+nh3Ub+rWM720/
2mM5ADWeVbTY8vrEQ1/o3J0MP6XLEAsQyZgD/AfVNjJQNCoohuXAdp7TuM2FhPc5180sT7H1waoE
jtRs84TC+kNWGUmI2aqlPPVa5dXbAgWDmX9elBrwq9JwqjerbY8GEZbWk/ofklgJENqYjDU5960Q
ab+Nfb2l8Tw1cc7I+vcmV9iBpaS90NFuk5olBkYf4caJKfzT/Z4/luPczZsoz3pVPAtRM8E66p5v
6+6Xw5BBNHz4qUyrfsaiynXDUs9N4yjSJaflh9YrZpT1HoI025kgZOu4mRBhFehFsOH1nUmEPIRr
KgIOVBqToobO8aond2dDYcE3D82OXTEtH3AYxEgMWEzkbwBTT/rPWSe3j/a1QroR0UF7Qp9eFt+K
L5EU4CVGp4CEEjoYgS7tFNmo3dUkWCWIHJowRdjXCrXOWiG7lfO6fIZEbtSQTBSZdjIp1kjHZ4qV
1lVm2ONkUIaIIJah0E/V0xjaonAv0DdnJdBpvKz/9Oz6tEvCsNOZ8+k7/aN/hlcPRFfE4RJUXN2B
CfvteAlyAhi6OUticnxddmHhj5ArZ6+Y3Khv3kPSMFQ+ooyc0NnQmGnkU494p540CSjdwZVhazL2
a9lem8X0nJ5ANzaB/wrf+O5Ka474f2wxt+Relsw9uwJPMOlwi7ZYrYp88Q/WIRF6lMjQTjQ3jCgW
DOVn8+2ZYxbOgcWonpbx20NsyVb0pwUxXwCZO82pwFJaNckOQ01CDl86gorZmL47I3CTg7wRUc4n
pkVnoHIzihUNsMObZbnnKdBQoYloPSXcvQzQ1dVgInxIxozKvs5PipLu4rYDQjPejN6qRD+u1SA8
UsRh383NUf0yKe/jYCbtYvq+ApdvXanGx2FCnfBhX2u0nAakMenaUNX39sN7UyA0qWR36LtelXyf
V1sexbZb0Lsn7vOw5XXSDErBTmG/Dey+hy38QHmPQ/3mmN1ONipbkuIdo8JG6fy09HcpATV6Jze0
srIZCpBUfe4ZUy3eU0oKfvzxcfQT13lO2g9XIKjjiq6sSU4ronlrHT9tcNITR0alBNaMAhjowMAr
4VjVpQbp6y/Ew8IP1EnVKdqmciFUNtkx6ZCqjiv7E+/zGDUp6iuddflF+CSLZg+XrfE6fycvJ3uh
KjLJd24ZgO+OeQ2VGwUwO+UwSwUsJyLzU4QcQwRZabWmYztObIy0x/L72asyvoYfWA87Zh5d8yZU
SWpE51xePO6mHw5kSBWcNW9RoIRNGSGlcPQ37FQjq6ieMlM55mO3S91B4SZnzmdpWXCpx/fIFtem
cEBJMdbkiGWW1LQAdn5F+cm9Py2GdPZe84Qro3WOhGgH1kb2X/MVyy9PdklwASiuey4NwrKDnyGf
Om3ZvxzyZ4zhQsDqhLkJKd9DhjeOBlMtyWERY7JSFn31M5WtI0nUK2XZqBMdtv3OdLwbVLvvUVSZ
mp5Ljp9fBxabJlrmTCd0JgMuhDAt/MY6FXY8nGYnyl5a7/gHmkGO1gHMK8AuHNUfOd1crU2DaiMl
DdO4I4gRiM57ApAvfPbYQLc4fqU3gyRJwdMgMN+MdgLT+u7QPdLH9vEqmxNoBMMZgan3QIEtYrHs
ARdhYueUI3ZsveFjBFNN3UasAR8E4B+WWnGts7gqZipP7iUVHgi6kWcuVn1vUfUaf0nK0rZjm0Fe
zSNsLUH8b4Vf3jA2c1V+YNIP2pZrOS0H5RS5OyWpdB1I2ymQ1yMIOzDNawgevTC4ThFHzteYgGs0
IjGbhn0t80ZwFJxJBWbCx3/owYwL1fVQixV25AZgD4mqFevUvP+4y1E9x97MKAkR0pm9YtzzS5Pl
1crVsXtQLdcnmXYvCT34FEUikpC6hdiXImdn0Xki81h9nC0YJ0q3Xq4rEEYdtdL5GKuo3oMoxAk1
AEljGVRRG1qw7sbUsBl60R9eHVr92TFuRmk8YERbUmAQm0WC3QEuhRIVbEgNRLENUCTB0gWXytGj
J81tzKK8JGR90q9JyFK63cgRmu1E72faCJSxcnQSxC94LWjGjTG7uxmne9k2+ONsihavvZyxow5p
i5tlriUCwV+jREvsbKE4gG/f2Ox8n1n9o5OAHTbKakqUDQe1l5pON0lGtSLjVJvphiPbgHsBEZ2A
tacuFktNfCfM6bbFAfp54HaWUAlV7shgPftst/xtJmOPPaPwihfq8h7noWZDpx3eEFzHMS6+aS4V
rZOm69UNGX9IXuUxpsP3eT4Hm6NLkhQW7iC6XE++jKY5CESUJLux8FlAZ9pr/n2BGUAGNWcI7ygt
wHc1R3rq1jcpynot4ZI49opPloRclJFRIh+jhdqfa+syqqfgOPhmDNBo10wBC8iraE4/ng6x6QGo
IHNBJsTl+3Rdulg0zWgUsr5JYC6xriu9g312m79txYlp4vXfDHgmS+X83yScxSP1puasD+RJtYDH
JTn8KlFIguGqxm5PSFnYCT5EitZSSzFv8KB0PmJBQ88mygBVO1p/C0kkpqsUtolhDUqiWnly5VC/
cPfxPZa2sblei/NAI8U4JXdsSJmVIW+N+1/+q1hZYTqIxvwG33HfHuimT5Sd7ndv6IycW5bv9skW
GTFXVHaK0h5HmUSjapIy3x8Ax+8Q/RfP1z9DgQGuLFNCnkOZNz12zAtvBy5AkEOQ2EcQvdv+DZJx
9eoJqAzGCLjsl8sakc2tvyrDaOlvKEf/FIU4FQiP/PlsjKXwOBPkpQsH/Z4nA+WIHXC/4g9Yi60d
i4uYnz9KOAZnumOmUrnVJ04+waGPXzopBB+h0SBaENQIWrDgHOTMXazbsmGh1DsVj+vYZ/8no8ey
4fAn+2/JZ50wW+PWuemr2Z3VuEUBaCl12eLJLJm39eayr5QpQ6N9ioY681ibckfbyCuaUQl5faZT
TStec24RRlp6gP99XsYLeuJ5uOsKwHZiLWbN/h+wtFVS9senO/QKtz33w2nNc7UzBzYEdJ4t8lOf
keLclXqAkAABlNr6N4j1ZXVTP53CPaYYFU3nCsA5B9qo1iyaQySHe3LhplAdEb7Wo7oIdGP1rSox
4fn2g7/6NJKjCaIYYLydH1GCIjCnUg0r2/KAivM/yGJwsjl34/W1cvZFfjutqlnaY4MSjr8zTAlE
e9ahdbO+86dp8+dpt5Uw3smMQ9IfOgoNnOjLTa4086fpIpa7kiDq/oVnLIYxV+BRmQlpIiNSW+JG
BoZVxnQE29K8GsnljZo/1QY1WtzIrE4XJkBHEU75MsNXkTn/Jma6hJyxsrNV9fTprG6LzyiHYmFu
8/pJedftrXacUFgUdYuJubFNs9UPQWbpm0hph3Q2CyVkp9Am5OaYluf2yWHUQD/AdZKaUbcdX+dz
bstd1a863YCjpKvLe4V2KsxftvCVQv2pgWDEtzOA3ZDr8I5Y/QLo6H/kaZa92+Twwa9NhGcXkq1+
Cj7iNR667qKGXN0beo6NvIaNlNU3eO9AKNKA81MJKXOgfA7OTRNVauQi3RLCzOqXH26+n2EB7xUg
SoM+Fanfc4a3elwcZObi3W7JyBtXWXsheAWqKdwDWebn2sAE5XfW//hbzsQDBRXGjcXwElhB1sy4
CuW+mtCzudtZj+mRZNncFwcL1XotHlBinisnthSNvX7nBR323A50vEpcIzi/Xr7KLGGmbu3XfOmA
ph86vpu7Qo32wGsx+ToXmfl7gT4oHAJ+s5SN87JzEt5XMcr1Q4glNxuTXM2JBYgSSswvaT4w6WU5
MD0IFfmDCAFUAE2gNuy9m/a8vFPo7zGWS5dmTftTrfRnA5VIzQZYXUb6MZv/YFVcd+LoVO21ufcJ
vyBuvKkgvUG+HX8Jt2X4/PgoxzvfD/EmVg8DvemMvExUybuNxgGoJ9vbixEVL9ew7A3JajAqjzvF
dscsB8hnJa1torw9jomvZUTAZUfGP3Lxe9gIXoyLy2cH2ctpJoeqv28nhLA8dq1coiZP1VYNXBwQ
kPnGkDfQ3ZMlzb2/APhigetkKeiM7t57oPcXTpNA+6BUmiTAjS1GcVVCFD2TWX7oNBoZ1kXNEDEj
5IBp529tKwp7BXalAhL5OoGIKGNBpsXfABkXhbfgSYMkYxHwxgFy2a7OACr4bYSeNvxQTnCMpNpj
NGhFOLS2hsvhKns1jBE7nDgYhh1bqwjIJM6sw0gw3RwiSoBRtBiM2TjjEnCDYBoC3KZ/VFeR7mLH
INXl4lI6UixSCshkqucd4Xcmyh1qgpm/XhDwqGSdDCfDrZATcr7M0Terw7kwy4nlnLCchlNgT0jd
sf2Rriskyp8PI/xhNv85cSBXaR65dEAFhJurJy1GkKy3OmBQePy6w8FoM4+O0JyqWx+Q2OlQI0Do
MKTp7rGojZHKjTNd833pQRgQQFfaIymMIncyTp8SEiz/UAmIQX/YX5xIWmH/kNC28B//jSx8sOkO
6r1FkhHc8mPgX1NpLXxhM3L4ddiWS5spUH8Gnt2wRbfHp1Cy2iHc6BOZ/orEC4nh1n7zcjFpPfMr
xGFdL7ed/MOisFYd/C47Bc+EBoHpl50lp7++hlLlDZGRAVoQKwocDfegCPx64h2Mqfti2XqKrDvA
qZ9QLbKBgO1vpTLbbRVm10RMqwPmmtpxhvt1t365720LWcZyGoolXHZNQzfmX7eXHWt+WybfQFWB
MXJFCASy+JDv9dCZdpYm+VxdcRd6ZCB9rcwTIz+ro0P9Dros4DAPNqmC44mIhtqdGfJ7deNJZfzU
Hn1RlUbnvzQlREZYbmQ+/CnoMGH2knZeU1JWPvma06MK9Z1Qmjyn3cNBsnTOO3Jnq6amUPQmpQPK
ppGcfH/qL0uLsUvYN+Yhi6p0tDCecWiuuF12Gm2OAV9MipDqUX0GT2J8brc8d/bHrolc29hSzeNt
azIHG1ZK/Z2dJxrBw5cDPug/sc3+bdLkg6b0QejtwqY64eSO6/VYMlMXiz5I6IcgnMWZZy1H5WE7
I4Ot67fqw+rvz7GPGNx7rBUh7IS0Y77G74XhlnLj2AqA6z9CSaW87STl5MUIgELvJEWcHnZtJyT9
ZT9BrfmY5+oXY9NsVg4gxH+tLx/DoQ7ZJZheyXxcPGzOWVcVlStVlswoePLzH/WiDGvj7W9QctVT
Gy+3Cyf001RsVTWbC8glcVzO+QjVGneBMGRDqFqf5yqCRCtcduK/ThjV36Udu43y3BCWcfjc2sd6
uXu6jIxAU1lkrG2utrekly5DrWIgLov9iNvsjFTOF0tiwLc7uPn3T9R6ytkOkm2sWLFqhVB4Z7ug
dsHJA0EgQyjM++J7XZ/kO4AgxrmL4GMT2IoVVjDI2MzRpD22PFDGg3vbWLidAqNEvMNyhObVafOT
AkwYl69NeK1T3M8TPI0/8s3gIa2QXKbQusBJg3TKmvRiNw762RfJqxtJCZjas2ogJvazVZle/Alp
4N5r1xlPxkO6yPrmszBM3YBbzpWqz1/d//bsyadYmztQvwqYIVX5qnI+a8XB2MueEifzY0Nh9Bbw
l1y4xcR6xIb4ObakdGTBWXcJAZb33gYdlJqHSNDPFrH8YktD8SL9JaasfubK1nz2nE9/4A8NeVdM
IonHjponbmEgCrnu7A48z+CcEF0/PO+VxgcumSWMtHT2W9fOeprbrHJ8r6F1SNQ8oJwvcphAfHcI
EFbxO5x8pJLf5AGmB17IBodpezHiSwGQHYM5Jyv2/TYwNn0DbpHvdicIlDt1Z46v4iS4jD2c4Y87
Kj0q4/QjS9+l0D+ScBZlrCrbw6EmYbwUPzLinq2ceJs+t7MQNAkw9g1eREAYXHaAaR2Yzcim/I/z
1EzEUIYU/sZT8Vx6c3bqMnAv+O7PKIh6SJfpdCVGsBB5hWmJrex31j7/si46eGtEjTeSRETB8L85
cU8DcsbfV+CqzV4t49AENJI4SUlBt4el7IhtW8chFTc0Qc7ScD1Uc1AzNrXxdPKJArGTEjSZnljW
szdDaPQUaa6x8DyQ1Y3FUfds7YVjmwuHKkKxWQ7Jd+VIA04ApfbY6TxPXhUjzIEF45A++O/bvpKH
Kbd++ofS2U4cC8RrJFyvtA9mOP2JegUWRSZ1Aju21JtlD10/yEjkN+7XMaHwacH9uNtridTGVMxv
5hCTISQ2SpMZwCTa//R+fkqgq/BZ2yLUvecmF8UkliGSsE3oil0rD1g56NnxoiEP6EGHhBZ2EwPC
myqrnMAFV1+r16stvJGVGeGnMlzu+eyLE9ga1zQp3tYQy/ot0qChYvhg192mYrF2Bmude9dqNPgI
IBjndcLZzsorwtngnzweyqKLveu0La0xo5XP+DWfIW1R7DbPY7mEkzlhwLjPNl1l0uJvx67gXWp0
Y/wCrMWtB2TIeawyJ7WkNmlKZhGCQFqjqNbtNoK2vTdKLkSMH7La6OcL5zd3gFIws8Gtymb6cZCx
JC9fZpQm048UHrGKm87GQGLQGOvhQfyZ2Aw3M2uDcEv2KOvy2XmJtCSMnFM2ti8XvhHXFvELTZ48
DblE8xyT+FjIvcTDG7IS/j7KN+HKc3+JUar6VjzJyLoaeXtILro/lv6tuTVv/jiTVVmkEDRsS+0b
te6IqEbaqZ7N8NHiNRFC6BQGvfLlQB/eQKFxPgFWOitPlJsIw2YwNVatA/zIP7oyIlaZZ9nA9hL5
DW5J34tRbA6AFchjUR0xQqPqwDsAJKpczaBgmqgmY/Uyq42VQDoFLgqqkTzXjhlww5/uwMmA0VYr
LYz2du7FvmZbS4VAqYixa1rc1VsP5re+Ei0iQtIB0vXYMO/q/MYG9MxxAPy5zxl4PN7R5KpHWcjp
gxmq5Ht5BsZpFvrXCPNaBbwZ7ZsLl1FabFTc0kwpdBNlE0NZlGf6ZvoDaxiyTnJ7Xk/lxbPHzCEf
eIF6dOVXeb8q80EJaBbuOsDuF4hBAqmyE9s7GbGkZf7TZofkBiloURuW12vk/vM76FfUg+rWgcgJ
smZ8Y/tzAgYPUdgZK6+md94cJYtfCzHJqWuS5tmNC5fR7+wDw8Hn4Awq6K2pxH8Zoe4a7M12iY/G
+dJPQf+VifW10vEBHuSracKdayJRkzm7+dCBMSPyEX829tCYetm0gseV+idJllsZYb7Lu/b6I74d
fdj+rV12AOq8fRRRxH0kPjD7u0TLT4Ss6lKeG/NfOiCqiwUL/t0W9nUZlV+DNDoya/L+6VDB3OB7
IBDMdosD83Ft+IKCKEuBZizELyi8chkPkTT4F42xql1cD/KnT8o/1GYTuO0ePAnWEJPvpg/VQ3mL
Ue3b2MmjhpKPD2l8XXOzEmw4rP2Ys48vjcJq5fHs54bAq47vRdYWnhuZ/RXIxV6W9hu+J3OD5Dkr
TxIbhnpUjj2rUJQiBtBqtGHVI0xBvBc5VIWzQ9rwFWq/bDLbHYM5Ec1Axh+HITno9uA0nAoAX/9Q
e0+Tcn/GDD7gKqieMwq4YLhdDyxqOI+gBUvUvs2FTyrU6eylqBHtpIqUJ76r4WWQXozNnINe2zDX
o6JACnjK/rsK7pPwnmDaDzmfE7vJWqGA0abQw0zTpKoymz0DohYMa/tSgJM9QDEKsr8eOdNYUi8k
BbLigdKVTalLt9YSuc2tlvDgtmiMt1ZfL7EY3kVi5PZBDyzAMoaj8aCjyXAFNQDm4ukN26Nj9dxM
xYINTnprES1liugu+xLLBFLvWBn2CDhgC2LaQXaM1zVtKxadkoh92vmHspaauPrgcvF9oliKbLr6
x9hR1Fs8f2tOow+johg5mG0yt4VK11FJymiMjZRGF5EbsJD+d2uLqNK4YkVAOeECT3/ZkQxy5F8w
i7UeNmrjTYn5J0x2ObVEguZ4Wk1zRWSWUR54F+CWplFP1dzcyP/za7q6/2/Qu1vvm4GnHzb4KskS
AvKiV5tf2hPNULwCVipFFeTT/HF1CJ9jnyQo1tyvM0cTuws/PKi1K+h4HJK5F2l+3eCHdTTti1Kc
5GlGyc0bATn6gEYyuYFUUPapZqNVKO3+9gmcglpBEBnSQ6SZIsDm9Q3RQY/cmYrUqJdcVoyXBccV
uSiGE1JqlYP2SetFDJEW/LStMHlosFXf30RfGe1OmnOtd8KeOYa3zLqcfSpSdNhPNxZwVf2DnJk5
HeGc9v51qqR50FixzOVjO+pcRGh11BlSLCp3OaDJIl+g2Zngiw3PdT8bTrlMpxcolccsjJTJ0hy8
FpGESTp4zwZfJ5AkIQT9mSXpF8SthIs7Rr3/PhAQSVjZN3EZM1lujZhrKNRGGGeF/82aRL8eh5sC
SioNOV6DojAQAGD0GWlPyXR0/mPAYT3gouXxWCdW6wnIHmvKGVER8H+DWeCrsuljEP3pxK4Bm1lk
BrPbwOgDbGtX1QdoK3XV6O7wJmBJN7Jo6mYN3ud0TypFdSyX7mQhd7I26sAuupyoGSGC77mmBt4Q
ci9rphIbD+LqQd2uXnSx5Y1BxN+UBfEIYe5YxdI3Np1pcZzpDLS0Yx0aRFUXx8Ard2+/egK/JQDY
fKlXQrL86dgbPFEq8xdzSmmCfWbCjencPUnquuYNiFfFvM9PQwMFW9lsy7FwmMRJrKsoouHNBzFF
f6t5wofO6Rttd2d6VdQsHQNZoEPQhS5yAxsFjU4kgt7u3ZjACmA8NwlrnR6M+6eUmKG+DVpN2D/5
oEDBo6cakX9RYQ9GThTTomwmU6HOH8njmrQ7Gr3hPFHWye3ozlOWm6a2MGANrq6mFogy0NKQpqFq
Sw5wAnhWBtSLdzAgIwh6qLlXUVzHdHuXnbl8oJtX4GcqWXlOxu9GjZpoMKskm6AH79TZYBnQ6Bh+
IxWR9r4ucNDWsOSjVilvbFoTBzi1yANmmQwVZHTYXwn+gXPTqdsIYejoiaDFbmR3ZTk+8PUR2QJd
OblKTEXfjKhGur9qi3IMPBpj2r27X8M18xXflWDlhL1uNolT3+Vh0W3FCA+T7UDZ7mwggPfZI9BU
iTwdn38q26/siih7Pm17rvejD6oHYxusIueGIGTsi6vQaLrxph+l6lX/64edWVLsr3p5IAqwGFRQ
F1DCVX/5scbbMfsrNeDPywdshGTDnmRqGnayoipDgja/J+te5oAPwBgSiPd1nqq1wOPnsRX26GVR
0bfgmXgGIFt7Z8Jg68gelT/PmM0K/e3Y6YYWktnP2n+NzhIwCvEyLEeRdXqNYzCh48VJRveKEu3r
Qhja+hAWjFVdaXo3L3KxM7sQ/zys3PLPF2eMX/8jgC3KmSSTatsUWEoIwRHtwCC0iQ8XXsL8rsnM
Am+uPEZUL/D2+zMC1lZTrG6AWcBCHe2J29zsIgJV9gRxxtTUKLdW2EdlawpL9iLIn25qTcBJ0ycx
gjXBQ/2E+pCo/SaI/ZfxBCWtSHpL3WHZZn5IRbfngBASRCUdfknod+f7yYpg3np6FMQAn6f6oC9D
BDgo+x1bdiD5OVNUMDe2EFgXXsXyGti2qHzZO3UbXwhwiO7oHc0bEommXPNSRSWIT0434OsvHG5q
uZqoOY3v4mbyE5JMdM/lZDq1G420TE53NxBcMd9w6k99ogT0rZa3YJlZjOXm8395CmtJNbOAuXlY
JznOJtdfGOP6GCGcMpO+X0RuZ1GgvQFsMwKxpAtqMW03tbNCwiLgRGprx0W/n3vxoD0JvcNral6S
KK71rzoAlVE3wEuwQmITnHoiPg78ixAOUvacAQz3eEYFVxPVJNzfVdolM5FDkZ08A3Td5N+WCZFr
Ax7+3htU8evO1rajQd7KTfNFKImkkEqUaqgT75pwWPaK4j11HrYhNSFrcDlQPPtDf1iRU1DHW+ZH
oqN4TdH6fVRjJws70TybthNFGLlNjUfAvhY7TweKAhp7va80IgFgKzO5FXINiyOg6hQttDCWPRNt
YV0Fg7lONQ+THivXD0EuoYdx8sBl0enuo0p9QvhRGQ8xQGLKontiZ+U7FlRWDTYjo7KQL+eARY5F
647upUaIeHd09+y/ub5Mqqi7lz3dFKxX7eQS5Hvs3qJSgyWksjMPv/WJ3tc3GQRbUIwZzuOmbkDL
pCl3uR77CKHSZ0ieVIIlG2UuTXp0BemtPJLomiKCIvQEitehO6kxHAa0KgWDbbzO9a8/Xx1t6YQc
MW7V/7eAQlwv0mdNvkGIc9WnskWD7yDBKwyOPpkEWYE7k+D3SypUQrdXdiD1DdX4iFLo8H/Y2vwL
QD8MwqdvexYJiTb8B3aTc/LmvJTFeUGtrETOpamkv5qR3i8m4aDD3sZkyeLmx3HI9EEMQddwQtxV
bOD2MoCs4igXd0iFcsBObrV0KM+2vnBpQaHkkNYGSNJFIcdRhWDeWchAb18CEx4wbgV89QqQEgxr
4ZYztPxwD0Mi1tnJoHjYex9Ky/GhfArJSZs5wgSZjPvfEXaU9ktNeq7q3e54WuGWCFThBCb5mAVk
pxjNlG7q8iWMi1Nd/p2UL+gF4trYErORc7lRVhzUlW9nMP0sl3oVA3XqNfRvbdL/dlv1QqQJSzOI
uYwmxDBXhbcraRboWw54F8JQV7P5j/mo287zW2oM4lDs5sbJMJKFg7tf0PCSHDtapMRTlimByXnt
E8MC1Esq7gotMm1g2SbNGD7BOscFy7Xa64VvMQhkV7af1fCe1rnyymIPoDCACI44xI1qd4ZAbxG2
+TcF0+R2H0bnl2g34Au3391htliV2wYxJKoKt1W2Evbk1ddwGl/4qBX5pNLoGKQc87xJrx4Rby5n
92jsDQm6fzBMo/Jzy2lOeKanFTQLPo1z0qeY+quEs7Y29ga+/sb1YEUW80EVQnPBlVDdY2qqoDqu
T4bamFOxW0gGN5iHxPwD3zlvCnhiHTZSA18FuSUW5zqAx6wsL/jNCW8VDuDk6RhF7WYu9RVcykE8
/GGLc/jnAIPg3ZBBq+eCBxdpvTFYUvcAF+mxp5kDXE9ZScJLTSVr4sh/dxcf+03nVgAMJVNQ+l0t
XaKVC+OGMSX+g19z4U5I3AiBJOW2m3agQqDPebrHiAucv/ADlb+kX8T+MTQZ7r8jzcvQ/7S6wWuY
2MmPTRS8U405KZ/qYzNeM7wZ15jka/zGfCMosXh1Xm9A+GHpp+PW08E2YwQDJjeKMhOob5Yxdf/L
dRmMpa0n1wEpW30oYZG885xPUqQzhcZeH8PQngNCNAl+OZWRS0S1nNLPb9wHi5kxNKqrq64VuKZ4
SHvpicySD/YWp2pRUI0aujW47b84RPPA/xQvBCQjPHujQmVM3erfZ7jvZH7C+zb7DIJ/NLUA6O6H
Y1u3QlcxuRmDUq9oETHvdUUWDlnqXRcILky/4HsWEoMJRq2q2MRqrJQuaQI3qbFc5JaiRkDwwesE
OaUhLHKoGiScCDjicPisrYnAQnBqs7WsoEdB7SmAErFO2J39tngElrriO6iHQgxnrA7rTzlmRWzX
VztO+jZFWxJ9aqWI/iUtrYIQ1IY0bS+sjUPLrNPt0mUlIDXm7zlM5I4qLVm1+Awly0CirhfpCLT/
sfqTEpLRBAGR48UQp3bAr98zI7lWp01au0Jp6UGRtdyJ4kvMhVv8pQtVI5nO2gDIf4GUtkUfCD2P
9bjSiRH0O3I6dND7r0aeIWIZU6O40rw0IFvc0VNYEo5Awos9ILb9jO6V+kxGXlyz4AbrGNRcqKff
zrr2Y7kWbVmlROXDnng+DvZb6APJh528CDM45/rRanczyxhxqwcaospuYLIvkK+dGivYTYkDTVX4
WaCLIg+0JDBlYCV504a0FUzG5jaZDSjlZkVRK9VLL5AKPDBVD5FH/ZUhxoy3zw1K0T7HAG8FjwFX
kd4Lb9IJUHK6emdu8xTpafx3kpUcJaJGuw6HjdarAKCfL2hCeHw3tluaU9fbwL26OADEMd5A7wzH
az4ztgAcThz2owFgpKERA7Dd0kVXMiDekpPZzwrxt7zRGLCIQ5byTHaz5ToVYGQvs2T6jMjUsIwe
ZE6RsNRcfyLRg00DCQiGQEiQZCLK3BqieXzL5YEcAFcozVaF8kyhDR9FCDURdTiuCuPLeF6U95rA
70Vi5OB+PzRmvyjR+ojB6CWvnmDobb6yBbXd8FVHvxn0KZncfWyGmUZuEkYnPbU8fU9zBEiMtcoD
PGWiF9kukXbYrwuLjH5vyt3rh8GWYeWuagOXVDfUwnM4xHFa2C2xBVcUFgfVYmWiiIechedUVLnX
3D3wqzNOm8eCdi4ENi4pVO8lNHymIXPfkIU9ouEQcBJLuLlA/ioaPztsQitBL6RsbIIkEcVUMtMz
jyutdn53XRHaiyk9K1uCXobExV62mHIfg5WhZF6K4+iKUti+Hp9U/CwZL5PRZItIx1DXLtTgiq84
erLy8RmF/5JlUpl1bi6IZi7KdHR0bVYg+l8VJFI4dwupkfhPhhnkcQGSuaCMiM95QCGR4FU2OPkB
eid2L+S7Rv0LugcCoV3wLH0/EOlsPbKINRQGtF0qo0OZL3kMbpr0xQ59sl2MFS7DOK379jGn6boc
Iz9KxilN2+/XyYIpTYH54J87PJoX13a/iZi9vKQ/8TtD2rwoLbc47ImmYB7QE/nTKYmEuhuVyuQ0
Vpssl60U2vHZA/aoTB/5qI+xNVkVH5wsQNEmBaHLHH9XPMLsjv7fixUMprwDRvaeYQSRP0Yupv6N
GEzmZG9jomzSWcPK8bkLXCTJJLVe4HcWQs4ADNQmLKy7ofQrMIP8AWHZav+W6kNiM780jgEplk2X
o66ouRj+RUq7Cjnbe42wqsDZfIkb4+TY5RbPPeIyNHmvSwNHNhnm2Xch5kQSkkLfKaKICZwyFu2R
UDhC+UijYldCskOBLsH8AQmtmo9/mP3XjLziTwlp3xysXg7qQQurmimvlX2C/jb54OPGnR5Rlae1
HqHNb+NiWmVljKyLJ/nti3eZdCE9FfCO5Og7BUvs9KW3MKlQcWJJTtM3CWN+dqozpDkZu4+2Tc1P
hG61JdVPuEZuwK9urkTaJ4XfAQJp1u7rEFunukQa5mAHnC7S5Cifb9uNk/MzgiLDiSKwRYvoRjri
lYjbLCd4s0/FS9KZaSjALTW/1wZWzswhmqWv8ZQdbW6ZysMe/9HM9xDFFdN7CFITpA+qotw0BHoZ
jy67N/uTdxTpgo0nig9KzcRaYSfrSldlr8dOQyXYg3TxTW5bZt1QeHciRzQdoKc/mapGmD7TMBNY
P0fyXsqxq2ySVAXDkEJhyNmIKZSUzs3kX5YZrsQ9CSMLH0PbpObsnLi7PEIpG+hEvEn/3vLWGee0
/iHJU+6hD3AI/4tqvBmFiUJNIonMeUWLuG3RBr71j4MtU9mVaqRk1Cy4uRtV0vxobEgH3qNiO5jI
A9ou6/flv/2TcZvfP1VPv18LfotPcKIDmU3X1ZTvuXGTohzu3nyXy9/7eTLcLcNZHav4FNJqK6WP
slZRgjfRS1wYL912AziatSmbhJKe/IVE1/WaTgJ87LQBbx1FvuGUzbX4C2o76gPVEwI+wdicMqLd
BFFlAFcdUblD8GZGSWhGVBaWQ/UCn7ec84a7zw2+dObUXQFiOull1ZgfHJWTtyN0sDQDtu3oXCeb
lP9ntDnS5zZUMu8PrR9mluBOnUfDP4x+ZqmNnvIOEYssqfEWCxXulSQCQgKBLjGrOmaem64Rfc6V
yR02vMIDE5E8/OpZe7QnBvTn/x0+j3JT6VDjC56T7hZIoax74wNVnSArC1JupuX4crxmAFwFYRtJ
stTYoxlRf2CYWHI3bGxOgVLicSW3xriM/hPIxOyyBZk94lF+uk/BxKKGQDwduciLIKp/nkruyXt4
7548yFoC4K1fgp7+DZuo8Zidk4KkirhjC6EFyt3v+8LkyR2fmc08e16ZnnIcP6c0Jlnkx8vVF6j0
hOLnKrcKi69d5I60mEeCDLwkUs09lSfm1nsGGNytmoBDsP4uarYiuR0UpnNGOVNSsK0CJ6NWXMii
+TY6wd7uzbH5e35beqWZa9LYC7goxhVH8CsOs72C4/+zbhyGdhvIacs1EkatoWOw2QoBEc3FYy+F
tf4YhZ2Kihgw4gOTBNfVX1konHCQl72EZXbaqI5d7ESDYaMacyX1U/8ghRCVi1wGdaHeJPPMIuDW
q7/TWGpBU/PTFbpuLucwreNchltgKV7Lcc59mp2JaZ6LOrqQ/lp61pZJI/ZlgdNIJ/c963CpnZYi
4BHN3mih0AgZtN9g3mdR+H/v+nHwGZmkm1xoi0Qu0Z5Dee7AuQSp5Mcuk3TVPiPf9024ygL2QkzP
MpovXyvZPi1qe6xTNVK9ingrc7Tv2d3xD67+2voHmwhZpN28Pp4f0ce13MH5U9zpzqWl66dsbk18
Tj3kynrmFe/kNoe1k+P8/t2H9MZFrFZlPi+N3ORbqvhDDtgUB7DH9in6Y0G4ZEq5hejx1jWg9JrD
1N4kLcRVuQ/bERx76MvVI1k/v/jAv98hG7JrlObfjh9a3fZsIzLdyK+04nqiya/VR8rcNfpHraZD
Tz5y10/zexVj5Pvh8Jg/2VXK4R9f7MYak6SHMAQXiXeauk8z90Dmsf/ERZFdi4k2HXvQP9MJoh9k
mhQZasA/4f35UoBE6xLTKzR3flSyTmOTcUHjQw8TdlB/EDVj6vCBfmT6/bOr0HJtgkKRdDIKteGj
L3v7jI4f+j5c+Uc4q90whcG0IfUEIJckk/E/XLpPBMZk4EhPMAZHfMlc0zi63CAokA7U5rFfrzy0
8qY5RwuPDOxaaTPS6oi3YAW8ku/9VEV9J3pSlehPneFkVSj029Ad+bKRA8zW+iV3Oc1sSy8+8d8G
LqkeP2euWfxUKkJKH3k/131dcFeLZlA5DHZNuVTOvN2VJhe1TAhUMlGJdmN1AQPyImrQjh36bnw5
G7TGon88GYmG5pLHOH4FUQrMONbXTHLZqOWGFhY0cUpllZVD+RpG/Esbs5vjEIcQGZD1i+HEzPH1
Psj9YymYdguxsTtI3YulOM9tIic5tXOpLAfkjTAQKT80fhNs3rz4HgNtOdwEhJj37cKcnkDE2wpA
5EJ/XuhHifqbpFoHnAF4d/pEE8q9z9a8E8CwvUO9vG/qYjT4qBtFFYelvNEu7cLIYMTsrIVCEA58
e0mfTCNPOlxj6qGF8ZSTdEZDYzH7OWpsXy+BEWBnjme0SEmhV3J6fJMnkfLSPolQi2pXlSAUy1IX
X4DXSxmLPdf9IicKS85CsOxlOvQyDVan0SfFrFwHSjEu33/BosqrHyczP7e2F7Yy/xRw+FCqteuX
ZAFKp2BE5bsqk8lGGx4gFhkmSSH0oY0TaZWFR0HF9aurMCsKyDahtdlwYCllDzRwZ8VzkDlJuknm
xdo8x9TitrGYF48gQTpAYZ3kOKika/5VCECEkSEQuzSmj+Ei1xflWxCCS7+4STzUdrI1gd9LbSsg
gmEA7p0llsLfmNuvnS2L0+0P/BgOkyueSMVEr2VnduLH/mIUNw9xyck9LWA2mrhuA//1AF+6r3XD
C1wwEmHCDERbahny1qY0QF5B3y1kFESVwy1Q7gxqOammkpoRcDYLDHABirbRa6oesNs1yftfod/v
8M1bmY8ZAiHmq77gro6MIOgbHv3meYbdTBb29/oMSjET7yngWtTR/vnxkh/aQKuJ2MFbWn1wZN4q
6rlCjmsfBXhoZ74dDAJSDKV9LCyQGkaNenOrgIlGBX7Yxd3vfPiSykS6+qrx7rnzrxveLEm3Aiy1
0lWXrlREKFCvBYs5SvUGlw3JqDRFOfkkdtHr3GSnOOm3Ig0PIuJROaqiLdI6rvnLXAW7taAqAVjX
t17/9/5O6gYsejN2xRhGmkLuk2lHGH0teMQY94JBlLMfHxtkb5La5XqVSk9e5d7/cYXQAzPb0810
5nAIXBPjnoB9iAD4zxfyjh9C4YZ9t7rfHrsPTu5blSvxYcqMo0Tc+dyI22eh49rvlHJpptk4ZI1v
AIimDlB9RZLs5UnezoGui6DKOz81ULHqsSzPCkZQJiZZWBUJpowWQMxjwP2FsDrnLumtIladJSAl
PcO4KINnjSIE3TOsjgR+oFlK1pphiGwF0DorzkvOzUXgnqxK2OPaGd2Xj5MDwRN/PZpTl7NNY7py
fturDIptdP4gsuLHgzsRSKBymNjLx2VjRfIkeieIQQnpW1fV7oIaqGK+QWdK7Rd+i5hTT36odXzT
YUmQgbszVpJ1+NMBrUHPO26tcJUczZ6lVEAZXdVUhop/PY/B1VtZPiFtOUaTHVk8IuxUVySqLOK3
Njv3Ux9L7B2RWpwc52IWMzwv1oJzDv/exhdGqHt/F0aUvtLLT99RXW0Bg6CMT8AxMfpbnM6ZqcKo
B3RK6xNMFPIwHclKQpY4LUpAVh+BjP7JNTFutmOIUwln+rYR/IfZ5dOMJTBYPlSUjHx6PphzMZ8X
oOuNu1BWXWjO9OWrDyu4e4IUgT31bDfNss2YTmYV8E+1V7w3RtXKnE9+g7B0kHH7ABM4lDTEGd3v
y8+iQxvkAO0FCUKDGwmZn0YA4miBaXddHEO7yjz4JfxhpgLeQ7EmgcbMpZrFOKMcd4oQ6ttzbQ9Y
/Uwkhz9Q2EJgIZ8Jw0nMCIlejKPzvGkJL1JeVX+0ZuyHWLK8FbpeHprzB5VYiI+Z/eQ3DiYOLtCi
Gqw9vYEephj3hEtNXdl53jL+njfDx0oT/6DjgrICpqBn/9GNI1s0/oGjY1FimJ7vFOb11TXlI14j
l/G+aTh52T6z56mov6LkgiwTOmSm5RcKAtHyjmvrXreNx6rN3SPtNJIwqFGEfrbZYdeKpK+jjwLC
YFaakxR878Oye4/JtcWE8r64b5l4FuAIkKS4QS1Dvd2yFiaM9giFaLCdKslsRns67sAVCLUS5nTQ
akDAmDrIvmnxMwGkihNdYNsK9sI+atzInskv+RjTe5oQf9Zw3xpNOGiXE3+ln6OFV7KzTKMNLLuT
PzvIXGJvwk5rIbVvcfc5eDXXod8muftAftZHpf+oq6IA5L1AY9FbFlawjhzMC6WP2fotVutHS943
uxYNi1K93VwyCAM+7FTHZk6Mdc9wQQlt5HmZ+uhLZx5ap5gVnibmwzIUZxavby6UGCYMT6jYaURF
Vfzb7/dBYrZbbvcE/BVawr+IonPNNCRT3eeH+zb0O9e1NgKtLNkTq+veruS4CNFFJ9FAGZK1zhPf
uJGggkj8Yip1FBSCGO5Jx9OUYR/TJVKt/kGps5u7qIYacOZ+tTN/n6WBUHzz445f/1IqaIve8qg0
8EQB6ZQE37nq6F/9PwM4i3l8nFg+RSyK5UyZYRl7yua+DRewaaFKgbHEV45n1UTvjzcnWNIPVqSf
25Q0CwU3ioXNMQoFGMmwb1g4UinqZX5NKZ7xJmMOZO7MIl6EGEVQ1qbehGhEBD8II3IFwBPqPE8x
L8NaMX0nX/BPiS9XQng5YTMRfrqCGNIGWp2DES7yoJ2Cd7K7+YXL9xcXP+vobAR87AVYxr3Pjigo
PZM7ug1WnmlUE2iOnbL86EwMKycG3G1zKtXu7/z0UlBjJmSK4QAQZaDaxcwnVSTVOr3z8MNKW/JS
D3iSMivbsmvtk2d16Ox+cAXJWfdm5B+m3hS7qCymwBxLV87OJjBS3TD6+9+GLD04ehH8twD6dPO1
2Kd/t6S9ByiR9W/oqwvIzWPnnrOr0yqjWdspdXcwwxu1k2DO7osgvGdrghA8lzxcbWcqm2fBJfHh
vTO9Cv1pMG/EKHlQLYXFVmrXLNCDsD1BUeyK3O8tDFdJ7hUVrE8WLGVH+KmJdndsuoANV/kvAcBZ
jTMNEMPaMqUhbMIYhFm+Cjj1Ggs3HdkdAwC/YQLbf6SUXkHRyliurrZrvoy0+ECslEeFpasHDiNA
dRxH3KDXQZptxdGimE1fidV2DnjRbuJKxtVtGqSl4p8rsWEzrgndZw+hbBbWt0Dr4kV6rRAfCcIw
pPb2r1nEEtbZxcFPc57wq6WKFfZ1l7wQ+P22jyUeoez92XjRN4sNIuBKJWF7UTpH/7h+GDF0YORA
gEAe3B4A/1uoBRSRlkzTBA8lLE4gU1uC/fJbHN+t2X5ZdcDJTURYcLfH6aTliNFd41IVU5WL3T96
On3O6+i0tRoLYQZQWHID15wcHlS0F6xyN1zSYCEsYXpAeX0K+b40XxDJvNEKbWkAefsfkCBJO2T4
Aq3S7nHB7ih2BuGxrix5UKNN6xkRd4CiAjg+sXvJZra4UZrHeylud/QQb18k8D0tnSrgqtF5JbjU
NvvC6o7HJsm8R2wPXEm3qRYs1RFhF9+jcz0Wvf3fpRp4ZYcKrM+zd2Ge741t/WQ1PT5wzc1IJLzu
qA9x013DwaM7yEpAs8dLp1X1IUZ1vzQo3KMr0gZ2zVwLj+1DtSkgNR5jtsnZ4UJ4uVRP7Djy/xX5
ElmEgTPRVkpwIb3bJNbIIWivtd7dybiRJu/ZhMIjZPN7UlUq0m6gMBcM08rXO39h/AtCW3XP6Ano
Jyu29AXtWi0L+/DdljEZ7IDSIJ8JTiYzI52hyP0KocNJzYLnOe8klEBUx6nK3viL0lZ9J6yHKX5i
aLO/ztcER1RX8PIRBTntvUIWESc7EcF5/BWvX3h0u5vFolFq6Ma+qwwLVKeyjuZT9uG736gEYZ+7
luHoa63K7y1Dh2iUhkCTM8t0YxCCWpXzlm9edi35VpvQsfuJGe2/juHjnmItekkgcNydUAO4fy/G
hdymTjhKNE93UibM4PfMYCBQve43suFVbwIIM/+Cs3QIRLfu/ZZkmApMhYltuBeOMu+0Bw/gpLLH
aSFB2pY4T/6gl8zv8wZIAJ2QsyS8RxTYggwNwVzBzsGMprDXIfwPMe8+jI1mJj3i8TGqgNwLe5/r
hxtTKIHUMv1d/CzrG6OGP37GAhBlQ9QqZxkenc5OpBCv9+TaMwiSOARy2SzfHfa4nxlOWpFksW1J
OC77kFoUdhYlN7niPQhD7QmywkKuPc2C/0MRWA4ELw9WI7/rWM2zzn0wZVroTZ2VmD+HyiAPP4Mh
yFJFO7dQPfoeW5yX/RDkt/h3DAIfWpOWVVeHMgXzuChNuuApTjkGQxez37nL1tjUSTmB9Rqsjfy3
vCCzIyysxSnUqvqr0e80FLoBSH5IWl+Dy21sssgBlnEPUIOB/r/vq6RFJRR7SsCXBFAWsC5ocAKh
RBlxEICj8xlkEVL5XvVYiV0bEMpR1oXcuI/yxR2a7ToEZcrpKKf44KjM/zQoyE49Ozndf7D40Ymz
Q5z4rxQKFdV60rmkLzICnAgmVkcusPzQKMIwaW66K/M18JoRBl639KIQXRa2ZLXaxIDyw656JPo7
TQrXiZKwO3E8e+j4Sr5qwHvYkUJK0I+ElHODTdX6Jq15N0Irexx0uoV739SzHhzcUi4MBSJDoxnd
GIBpTmiONa/yrF0lObMYjnvkQt83gXM1UMkCJzZJ9pWyACi9FWu5uF7p76PZhP5ACZEZYqkOtkqA
Ao6F965/k66CVMQqE4sSUPDRnuC/dZ/5IztdkqVL6N+35lSMdxEXpGqIZy33E8qZRIUi0xIo78GY
xmDcJLBhISJRuEmqy8BG/VrD7nKTpQE62w0MLK+dTRMyhD0mGs0FVYejCPPzIn/NGb5UeXjf9CQI
Xm4E1WH7ekViKi47KbuSJcen6ug8Sv4MvZyijlH8uamaF0j94kbHE6tK31LLS4tzSWFkjrJG+jSq
eoUnYpr+gCL7fw4wR0AIeuAFJ/kVRWd+cVCv2dm+7fn2O8aKHblPsf1C+Nw3jo7EeBwPx7vyY4EU
FCaZqbmcv8rac4znQbT1l1bHq+LwIjRgesuEvO1rC1nb2Tot0zmAqjtxv/u6niYIwqVn39SCxIL2
UWuY5bKg1w6+AwpSKK3HiEfnRSu/oZK8S/RYClQ5XZmjZ/yUNIe7pJz08C2O0GdU73OAxlKnQwom
cYjLZox+Gjw4wEQj13WGMYx3HYfUBJwp4BiInlXgo2jSVATNAwCs1JFWNnYgeiHn1sx5aSiVb6ON
oQerj1W5QhjUkEc+RcrQWLVoTa3se2b9svu58uPgFQNz/MHBApwEWJOFUeWDXV8vgdTiZjPOOwmQ
vp9Ms6bWYfrpNTflzwliC56w4niMy0XQkEFrg2k4QL0hDExcWkYfTAlBE9Jh775BDsjrEQ4xXv0L
98QbSil6orb6xwI3Qq8opFOyjrtS4LVz4xnzCv8GlccqkiL1wMKgNvOp58XkMOLKAp3a7QDj/8YR
h1LwOHQhGr035mh7OjeXwapo87aCN6ANGVCCKO3PiU4p/lXd9+Io+MXdmKQ7UXsmKsrqRM/ZKCwH
Xe1yHFGio/MrvfCelLhlLR6wrm23tpomrUsXljZc7HMxrQmq25itczL1+EI8rqFgljho6/sVu/Ik
akCfJTjN9+I++W74MTgKfa+M2AtF5X9J4NdQfzb6YhvZmX5EZNSWSo/P7CJdDbMdnSAl/zpOhkah
9nS0qVBpyNcHPMgxInK69SwtBgQ6RQXZ8agcKZKLeRo1VVuDwWiE3os6nFb2XWseRca0cttoWxlR
j1Why3mP+4WvfbEO5R2U0ztbOneCYodVQKfoVqdrw9e7OPk4nraE39+yrfa3vxywbwanqhdCsChc
cRykbQ70LNQmo9g1hIWKYIqeYf2oNZynRjHs4gZGwtFYqgbDfdcGA8veL/S1Y+N58dbw8109NajL
cQhjdKDK5RjKvhYmkwx/MzBxnp4G0W7Jvo2SJ9RWdRGli2TdJZ2Jad7/K0mLrY0X1y+HE2ozRtks
ajyrkjCPesGFWfgqzt0CY1z/UdMUPutkWQqTZ8qIYrWAJetUvEk8Kdbdt8Zb+Y4FVvDQgokF6FDK
YqCIopIt45zrHsawWm3XVP8muFnLyGSMlAsja+NtbNhW/bsLuTla4vWZZWX/ntVQXGzMNCU5mXt0
V/b2CN9szItQOQ23pXdXxSKER/lQMLxfl+6MD/RYTCMVxZ3hptlnjUvOYD+iYlgFtR/9w5w9/ZDs
RTRwl44cb6SNaB1LM30I3uG5gmNdYy3DO+qanmVDNTVZBSy3+69pP8MsTcsxCpBrmEW2JxK466hy
Z2R77D9/QY/mwUttVcvSHrIrd2P0FftKL0ylZtd1VXXS7qKAiHvVm+GNVo9hjAXe0itxqPmvxsjd
q8mbHP1Y/x51qWphjPZMLgUvo9hv5YsfEDbBBYN4j5RBU31gdRZDa2lMhZHgLi/Da9ClbPLe0bDJ
4QAyVgQz4IPKzyE8NKn4biIXSQaf08WLWcXtQGh4ONfeio/j8YVvU4sjHNOW54mrajjbrlAmBDGd
lxRUhjFUfZFn8oRJaEJVmV0Xcko8lkSpw700qC0PuGnKoPxxu0Ui9Ygd7WQ6WJNr6l8VnoZtorhN
cKwK+KRFUis4h+Ucxaddm12+oSzRQ2CDAw4ETq3oXYH8LiivFOBCX/fyuJMyntS2UDkSPQ0f4DhE
rygZLLw9PdLE/eUB8BizhLsGzT1zluJKL4pd+TeEi2+/S+SuzGz6s/kQwTzVsXcKNCBtMuohz4Z+
NpV3Dmx4oQxLFfRfJKsUl9T8SkcMs5/eSPiskhq/8tyK9+WD+plsAzESDq4wBb0OB7bS/4iccO6w
1QEXuyD7KKLc5A+Sr+4PIgN8Cym9gAAPDvGaBjqGhS4PYNJmcN9qIrTHXwFqpJUhKfG7QLfIKNZ4
vG9MLMO/ouIsdBPP6ACAkcQPhGYThlTTkA/SKNm6/5jPb933NOjXrQ4Zc0vooGn29d5hj5g2n/dV
zrlxgvUGPD2TsTl2x+n3iT5mxvu02U9XuQYO4yAIJKsyVbid5Ltw1mypwFzksOkQdtp4xwodaGch
4ZDxll+htG7YEEECroAxZ7uAUc2LuCso2Sjv5cFnMpgi9Rfm35KvmtDcT3NyzXmDIYa8etwCM1ia
aXlmxdSGYEt6MUHlDGJwxoHda4ASWz8l051vmN2vYE3dzADSECSUNa6nyxhiiTP5zZ4BHyJzNZUW
4KlQV7DsVNf48Z8DRyqj3lAPQub5B4ztbnkO4fZaECfLJR3sFn2MpOwR/VKD+1ZpI0NxKyB/4mQy
6VSbXbbkvXGaGvxuOTP3lUbZbatfJrJhIQuLKB/mayDsvzXaeWCHSMn23r0M5T/otWGM3WxH0Wux
uF0tgN8/IXDqEsO94lkUc4K0q4JrM+MgjSz5MGglB/AY5pw09M4zuo7WbyFl62CI35le4w3E4Xto
JlxMlspAVJdf1UkOCoNqueKC+5a63Gll7VQmtG9kMF4VxlIW9LmQhIc9F5ZSQZB4+0wjgCuM+ahY
TmMfAiV6XvRPg5E0Jrb1P9ok5ESTLPpjyTGUcBKnODb8s2S5yZbCrq3FWOGQpoTuT6AsluPqL2n5
CCzX5m83Jezo15vdoMs2sW+9fFMlDeZlIGetZPcTolTdShWmx2pQa8YyghzXsuOjF4wzaLh/UJRS
WekID1yOVD2o6biLt0BFkrZoRXvoIyGQSlo5PH6zmdqWY+Ii0KoiI5GwyKG5O0nL9XJn7vrsbd8E
GTO03z7rSxEnrd8dUox5F8nV1Sq65uljPPxofi8XDzPgzI+z2NIp8SuyIBbrCjhg3LemzImN9fi/
YxXxHTkRp3ltcS/xl3qAiUoSpZbZs0LA5UZCX29TviKdpquf6U71cj90cZYv+qCAACg7fFmE3Wbt
C8Jp+JUcX92yZU35o2r6XdaOCsHK1itEvDUcugPj72uGtxp3tHc1wVTUrRMwZe1dW3bg7udomatu
pPbCgmO5Bli6yi8BexIG0JagnG8aELhSKNAr/ZGY1x289n1jPjBIQSp1AwBqF4wsIp84Fpb1BUE4
CpQ+NcpTR/ux1gykSju4tg9g53laJuqsFIsieoBnwpmmj4B5xOTbPPF1iyJQphzeMAacvTzaLK/A
JB8/0FvQfeMq1eGFbjPW+/cqV+N9YE9tHSEExV1G5MBjb1LJXiRXRcn67ErUj9lBj6r5UEzFNbWv
cIhTcwEqKEvBv/n6upP6vzobX5Y+rNTdIIeYj6QG4xFMdkyp+5g3y1tlDDmt3RqKetZGKkzadk87
ouyj33Gbfk6CQFqv3LLqHcz/k2qKh8G2/bDg4ycMkw33mXui8bZKNGMIu4twSwJH13MEL30/UNBI
mvEk0bgPnF9q+nDWIyUT+efkWj+TXtQj3ROQTxkTQz1DBBHkhN3aK6NfEa8akHxx140Ro0RlKWIu
R7PCumbCgGoyV74xRna71KW9rS8EqEeA+LVq/d3LOcCthnOuFNqZT2zWOfHlkTlFwNClapUDG+K3
S9Wgi4hwSdXS24WYYHSrZd3FSCn3wdClKXDrbdP16RGZYn/DWSBDoS/7zSXsCuWof+XKua/aNzWu
maMpkl7/st+5jqd06ss99n8Chnwvf0pdOKjQhJkCZ3HVZ1d5sJ32otxuWpEI66Qcfn0EhAsX75gC
0UFZ86/Az92mju5QEu9u6AjXxwekaZ3xNkSr/jcqS0A2ogbyl1xv9MBRveq8jPz3giIftLZ9or2h
+B7yZ8A2UFXjjcghaP4lPSEHGiwX0AZrp90uCAKpzYjdlcO+YehMs+uznZzC5EEGu52Xlr61DVBc
dQsSh6ZqBFWW+JOScuXU8Qo0Mk59xSrT6/aFrtnVO3nc5IWvMrZd1h1ANQVBowL7J+TjBDUqA7TM
u3S3C4lPKmk+CTWzVCS6lcPpUUNsX9EEuv6UfEXdgu7o0IaWy5zjcBepo5Y+gDclJ3jIg8cZ1lxv
SGEjSWhHN47oqMCqQPgT8SitX0IOMsN+aNT0EHCS2YVFRzxK80ic692pz38GDah9uo74IgPI6WC0
d2/mOLIkaea/HQcE1YpCgtbeRD0jBSRRybiRNyp5VHJ6+NE6citCzgQFTBPQacpTgIM6QgEywlGA
wEHilJkkqZJfWEnO6JFD8R/CsCf2vxn45+YmWZtMl+qN3dl0a65Z4ZT57r3MXzNryuo9cGp0iwFZ
SqcCieZlkG9+v3kZND36oEWMoGp0MYjodJd8VQUTFBeWhgKmLsN50iMIyILiXhmTQKlO4LhPqIlq
ZKadv8vmmXN+LQSwq+4kGiONN9Eol5IC1rjCH5UWyUAfZqQ1y+ar61RaRSAEKngcTakgBcC0XRF/
/CJg4bPRbZQywo9JndhGUuljEHG4tJRS8VnT2IJ7WH0p/aJ+1fr143Wdda2hwMhxog2/oMzXPD8+
dp5v0ARPsKk4vi0vOu2Xlg1lT5dZR1WnRpsJ+t81SD4wtcyhGv9ijMOxNhUjder7HlIisrUE/R8o
h64EW/aJK5wuryZLxbqRqV3P4al6leXtDPQ4fYmPqJ5n2G6BCvVuzYIR3kc8CBUkD+ALlP7aK9Wi
0QMqC7m+4jW5ytAfwAmT+XKf475+N/EkIbR1d0pX3Lke+TfFyws3g46hEUQwJHLa6OxRADDdPrn+
azh777G+P2X8/wagxS0B6sJ4eqc7m4JgLvNngixQVKnrp00FVN6HzFgqRL7jCnbXYmXrTNlg1uBn
X1ZGXNKwedj/WpFEMjJ9c8pk70xujWMatIQcx5s+G5W+yD+xOpDgJK16tZCHKXDo3AJWY5w1b0zS
AMMfNCfIFp74o8hNrRfymYxMRCwi4oS5dQ77j7FiCCuBc9LFZ3M6cXWBdRRxuyUpYU7ezq5Vxwz6
Wrs2SQlP9B1HAQzTwSLzmH+MEjd4D70KtcB1GJiEJzbMiC72xp2eCbxAz16ctRtriJ37wNXKGvpE
wpdgFfc1M1ZAVmS4JJzdTUVZV2HedFIkOwIbrwQpt2Y9o2yg4UhYGpU7eXY5OQKmLHxUagV192PQ
6lLFYAnkCYfKM4XzKcx6jAO8XoyKlC/7wp3m7JTTBuwvLnc1qAO69OyljurcIq5XYrUuiUKv4Exg
CjZx7eU6SaZ6IPXKlj37+d3b2ziao9O1jAMIe4MSNUxryLs0nrKqT/WsS3buY685C/Tj7LOjy+0/
VX4hlDgHHNzZvH7PtxdAsNS+WbTvD3Gangye8CPTGbUFWaFh8z5ob3DLE4rTvG+HfRk5/t5HSdSO
RcZbU+NgmkMSLQd+ceiGiXvmgMinQ4rQA7K4iHSKNbDjNBSkhevTw497hTELl7cVo/k1UwhzH1Ud
UeqZp+oc6EY1mHhE0kyQk2lEP2X2CuMBwMvHqODaAQ1k2XfbBlCMKCuZabC3tYnq2EFXmKmdX1pY
6tROtWxnH5nebqzpkAuO+OZr9rSmWi0dRWfeg3FGR/5/nvGiwa9VjmLunQEjzBGoSJ+fVdzkSRF0
zmmwAH2n2ZAEhmAkMSpEbQ5jKdSUR7m5rhdi/fUxwG7T8o7K+47EcEhuzIL+ZZ3GCxJP2RqIJwbk
HjGLXVRdle/7ryUy5RSq2GRIAyM+qz5MaecTazPRa04q6qZdXIvJTCyE2+ODMaJq37wKkFa48H4M
NLH/lwzrDyxhz4ZTNR4u8iQCB2iHg7icyHM3SFiE/HpCT/L3vXsn0VCJQX8Z+Su4tq9Xo6I6KAUx
qFcMzALKkrVc/YiorWqGZoBJXZg+uGFlHPCflptRILrcPnvpwEu3Kly0vpryXNITl+yWWL2fNxoB
V+d4skO/OEuccWJJZPS41fR68sUy2Z88BgS7vahYX/LMfsnbwFdSSDcdi1C5qV5Lu2yJjvdQO5L6
ubVZ+aqQEjIUn6wzXbVj5z97mWrxa636e6u68LHOdyLi9ChXrvZgAlwbHtZFsQRxnOCL6sFwDiR7
7cUgVMspRZRdmzwILYQPHnW7f4fWjixgqyBxTDMI6DlM7nRueyCQ/E9Boy/2u7uHo20ul/TpkzXo
W5mIyngdTkSum3nK8Qm754DR0ew0s/wIAT4GNldci48hFhfwP8n9R2f5e80IJsWNpA4KyIKYU43p
HvXe8GYRwLU9heuucx+S0zeQ9b0iIoqB5hxg3bH1uZuVrU2zB1Y3pzjIrhDNXBzAdFoUzCO1sRoo
VDSUgkLl7SDpo6oJTpOdQKS2Ex9PmihQNrRyV5561aYtuRmcK1NbWIEPQPaVUy8AeXi1R3h1TNU9
bgBr8QMZhapzGC+K0n44lRQMogB1KKYc1uTNiugGAUwEdASfyBQfTMtQxACM/66AU6Ye3br2hidc
zaACYn3HOKt/CQ4XHiOjDjFw0CCXvz4P4VJfLpDSpuMyIg8/ZcmqwAr69kHNKCwzIpW9pXmyQhVU
WXAg01CC/TMCPPa/mJcZyhHZmqoZTPu+T9/sBhob3VOnO+JKe4zwEjFI+sJkwBakE61wRwioEkzm
PyWGVkJhxerykOk3M22FK6D1Rf04vFp5H2y4QarcNnI8/BcNmJHZCfpij50A2oxjX39ZUUiY0BLR
jgf3iCPecYBuKC69TLDahZOb2HakSY7O78Pp7hCCeFavbE+Na7oYXPL/ar+FjfMghCVOCHqwAXHe
cf1QK9BBuejfPC4P/BfWUU1C3n+2TiDdM6f5AevUE3XfMv6kTg2e931VWH8PzBDc4xuk65MR1Twk
mXoOJykyrHgzjj4WWF/z9t9LPuFZm3Y0rHl3AkD7h1P8Vtedh4i3vBbj/pvD2ue11PfsHsiu8y3t
UMbOSRxw+2B5JbwqeTTphLMusnnHAFAPkphs4MZ5fTCV/aHw7Yw/NxYUmsfB5wlWhUXgqMhvEhdq
RGLj42kbZSHrviQCk7hSWs5TjI9Ij9llmFrUnwCjhkA9eaiBJYu0rFDcplmR5JBtcHfIvfnL2O4Q
m5GTZsyfIAdmAvPjcq3ZJYin+S330xtYBg5dj9ismv23IEJPPh1X2IUi1SGcTK7jsjJzCNv9CODV
uIAaG9u9QqIMlsBbymPv4sGmIMH53yFWpb2raALsA4nzSvOUXO+3HcpWrC1Efi1li023vTu1hhVA
X0iXVgzZQ5LctoqiUC9KZ3epJ1MAZ6592W6/H6INC4egyRAEJel7jJinc/KG54aFmVLvwXfuF0n1
mcqFG9szEhrAEpzcN5c3hUGOQzNmwaTouL5gn1txOeLLPXephtBK/LxY09rf7hf8+7gtS80EYYao
MPTsG5eJkTRveKnVXijV2OMp3+uKcsIOaZO1wiEcX+CKF/L5CpPGu2mDm9QliEmjpG0+a6J3ZXOy
N7sKmOHL+Y49KDdl+0vSJmWT6zCqQZd7jUt0kb/+b25mFIB/J4FR4joilr3af8cAT/8Wb1Ti3JjY
BABFN1+NCWGpX2gI32vlOId1dFxw30dMynnYxWLUnp1PXfik/Ebq4wPobxdhnXsFKbuzJRhwv9sq
WaU6dXDLRje7EvKzadMzNx92vP+dYHubjYjqStSMd5xOD1Z9GC5iJS8s5r9rJjJrY8RvXfI5mEaG
fIyC0FGXK3Mbg657lvtIsaD5XPtsFhWl8PDOvvz0Z+GcQz+2I/0e8fQEOOxzAua17lK5+ZYNZmQK
/zqBrq8zH18UEMk7YPvH6hQ5WKayXO3T/bPNd6NYjua1hisdBVCvUQOf9zILir/HGove7JcqHisy
e+Y/rhYkexg4HtTuSnjKnAxcYxNl28Avg4H7pK8poKJQKn09kPrrh6lPzSmfA8Sik+IPU2zY3fA+
op/NzU096OpiO54zPwysAzmta9fXNa/mDdP3DpCq3XyyKJH1mxrZz9bFz2VyEirQa568QVpwDUfN
5tv77vSfnUUs7daKvGDgTbN+YeF4PVWtok5L0PNdidTTRt2gg7Gyt6YKofDLLoTVMnjZiGb867PX
CPlN+3KWQSj/gXzQrI5YUmf90sBRccQ4a/nNcwvsGaLIl2SESRNvMni01k3a4sleFD9AD/uaSYKn
fOwXGO06nhfPhtWEfB8n0I4W0CCCYVxN3T+N88FxgZjEMIdG4KdzCkD1s5q7vbhNOp7B356Kc2Wz
ibWtCscJro9JvtjifDSzuxqlrM/8UdiRCFi6XSz5YwGLetgp36Bjgz5OmM4imxu4CN++kQHr55oZ
hFUSfTE8HcURnW4ZJxAr1OHnBoVeAyKvZoL8ALjdWu0rvVCKSuufUY8eCV10lhc7Z09jQ/pp8lOi
AZXKf1fTKXySfqruh/FAkjaeyiyN/y6uYDuI5E7pAFBbPBs5lRB0UE16+SD8k1eBYSSt4NhbHAx1
//bICGzQg26WDYyfCSyYiGzt/FxrAPbFbJf8el0dT6s/XqVLAVIAUWz9pgZtvkjFMhfQuhTw8dHL
r0x7VafDtR0I0clOd7rcsB4gf/iR5DqG/TEsSLKrLdlWXtAYo4qh9BOkrKlErZxIF2aocWKd/HGl
TDG28kx+hSE2OSGm9lVeLuUn38OtuKMYcfnfIrc+P8GgDg97YSkNUb/7sR3IZA2tbVB4Pv2hAxhr
2gl+aBh6Pa1JEncEVQbowrwQFvWfqdiG/C3mPPFdyTH6s2T+l+vqD0pSZyR/Ig1YYLpxziEJo6Is
IprjhcnX+TnGRi0kXO8r/V/wn3X19koTxepVURHiIWh0P/iH+VZHAso67sn3JoUOTm68ZfCodf/T
pA+Y7O3IywyL8DHIjW/sb5Lk8+w+VLgSN+q0JnOYRX+4x5RVgC928hQiAQpV+bF0kqX53lV8zYAX
IkDADeWgE+idNYrGPgk7xDb9LbbyvYo8uBvcULFgxqq0k/1qWHlgO1188Zx2vYmBsGi/mzzSrGEg
B1i3Yv1LJI9ItGUaQ5VBCs4vclhvGkAKt01VIj+zT/dRHgtthl/iOd/W4BJ4jB3JTuOIK6N828h9
Q6bRmyzvkA1Avo6ETdfBHhZ2BekHrUylcKHH/WuerI8mXajlU9h72XN+ubdsfOQIaE5rKwwg5DAf
KIQuBOZBbBvvcv6FCBkqghQXDXYVEu1ThymyEN1fpr87uXNPf8Y9TXi5RmIRYcfpwl2/JxLZqIXn
sAMkZbJU0UT1bRTcv//AvL3ii6LMdO6L7Sr5vItCCrWogH+rs8BwpZke8rfV3iegVHzZyHA06m6B
xuu0Ktlk1O3vh6yUESC3SiVP08tJPS3syCP7XoDuz+yB5DG/FY6z6dx6pOMGloMT4GYltgyvgcNh
DyW6JAH61wxAJV9pIwIExRETQdTsu27btznFc7xQsNyAXKI2gCXx6gknwsPw3E1yXMG1vdsNqqT+
0b3LXeqYQqEG6WnIsPSLkmowsOmMtjyvD8xPxH7ERVVBryBzUkx0MooiZsly8DcnzHbKNzSY3ik3
b51oyDKLaZ3bMkf4hVg9ymKBwIi12UOyEmmrdoQPY86eW9rzacmTMk3J/tg7eVIA0JB3JM8ZaU8j
TSzv7WqMhTCthVuNQVpOttz6m+PmGAY1XWNGmiZoNKHOp2iOJI/nGo4H0PdNSccRMywj8FmEKZF0
GrfR9ZvTWRCp++MNY0pm0ah+8ZowBSxQifxWKCiI7AJFCVjXQreu/sQ8Dvfn4xWBRWXvfak73pCx
vcgoC8zbjFl2Fj5xZEE4P92UL+GnTl5hf206KQHgiAsXyjesHP9yTQJm8z0N/GRq6QJdrsmZRmEZ
fJRBRoL283MfdP14RfdjsJpfpmm/ltQ4yuW/nQechuZZKGX+8iSE1jaaoMQ/qwy239MD77dUBXFU
LcyyhfYvvQVq2wKzJtz1elpSsDy5A+U3Tsry4Ctm8TcJjkwYh1LNCPjrzU1Q460wmG8k8hX5wMu8
Dq7ZtYVoI0rYgCLPxkOz3JfsCF5Tj9TaLq26WF8yHx6rEKZ9arnbOS/6f+lzYeApqGwkm/Bu8Mj8
atQmBJ3ycjZboZg7p2Kczz7Z8WPCax2ztbEhy4IBFyGY70pr6WwZdtp2+o1PAEAhOsmTw1+qZgX/
z4gLWFyIzvpOW1ZJdtA7Z/CD2P3j6g+fQEyjpi9Yma1/FpfuA15z7LQTXGmpUVZPZmIRIrp0cSAR
IN4cpvQhPOuH1plzb7HahwIBsFkAZQHxyaJYsSFcinQNpA+v5UxGY2hXeubIJMKQ7JQ0B1p8HswE
NSNaALh+VRq6urwQxvC3ygdXiZbOaXud7HOh9CTHGN9YNbhZ1maJe9JvfkS0JarxGoh4yfGOp9Fa
dn7Ukshc7b3jVOgzhPMXIuUeWgNSzSWhr6Dgr0ALvlm3OPATt338+pA0O+Hm8cnHK+B7VhF2+NWT
k8dDlDfrNodkWKXbzkRDSnJDy2EZFlRe1NutdTqjVqlaW8Ca2R4BR1qlm+OhMGdoV6H8pYJJVMja
KiY9jkHSiaEGEiyZLtAfgIJmGWQnSZuPKWSFjPRLlXlIqI0vmdR5y+16uc0svPIRpinF94NqBBhY
4z88Icvqpoc+OpM3BVevad1iKLvOSzEmF0od6/RmHwBWsArlzYbT/xspvYrBQhN0C8Xrc2g43KmH
SuLnvljuMRaXm23eTLzPf3NGEOdIj5K9jb2B2RtSHh0Y4hgcg6YY6D0NC/IkqGUCWZ0/fRhkcdz7
0gDodePsNHlwqJ1ekJfbO3ZbV7nFU1Kf3l/eW5Oi39mrzKUd3TcVMLQ6Qh5CAiO9MWoXf0XjilAz
xnUm1Ov6Vi/9qymh3fIuNkkWjqp8AtRRT9qGlynF5kAydvoPifg+MZBf/F6phYnPrz262hwSqy6k
jRkBeML86YMl7R/tOdwHqYy6ShHAp1TdOpFSvHl8/N5lnp9/P54jf7+YCZAsA2zhwfk0xK2UkmOI
JL11m13k+NoHPsowLUdQPNK7muMZgHQ74i4xgCRvv3PlT2sjr7IMo2Lqx54wzSHrJonZRVft3S0R
uF0O2GEFTYDfWSghYK1iSlxzlWKWmdVSQTu2JS/ZXNy7CQrPHUb2+/17BaSTkBpCk1lKJxwri2U6
LpfX2VRev/WlBCa4ThY5qUEML5rIo36vrtQuuZzYRrhfp52JI9BxzlFp28mz2bDe08SgxXNHWUhz
USfR3CjprHbJ1S4auVjdbIPz71sjt0SwxprP1L5ATnYsr7trJyPduYunzMxElZIUwgDtv7tvdk5Z
oV6dnazdPIQsD7TWROLlJ/XO4xL8a1Ut2+BDg8oTYZmXngG95Ri0H/R7xVM2vRqobQcFNQlQa++E
zmx2c9urGgMtuh7OqccdAmdyKTKyKFYOfcHfBOnaCeGSi1UHjhwbHpsvwEheRqAhx2g0MHjPaYxI
aAWfoH0NzrRN5lYjV9TAg+RDUAV787AAMmUkl1q7OXk0wZ9TA4+YVLSD82uCEWPiS4nqgnrvOCER
i2VNIPPcdFfHvElBqprL9yFbD9LDg37XQPJh8WnJ+joWmwhn2SDGvY2T/QshjC+rntkbr6Nrj9Io
wMBzgdizWJcH50EBDfmFGga7fv5o2tt6e7jgBpVARCNGHUlmecdtxOg+nidQVda2D+CaqKd/K6PK
7cz/UGwXsI+gWjkJ5621RTtAKz4pY/P6iLkzCtXZSMIThOPB/1MbmRBabvKgpZ1wU25DAFR2sB58
J7LXNqZXqi5C95CMR4vRQQ9xaUNxeGGhYL9NOOby3KG/i7Fgv61eKccmB8pxooUq7tMUwbxFBcT7
3rnkhSxMK48F6fzvenpWnEGp4LFbSSS0a4gLrRltpTOBq0tIr9yIit5xRTe8rwUFd6FAD9GARXXU
I6l5xzDyV6yD69tBVe4gWTyXTc+3ao2zCeybiXC1Ytc+MpFJiBupZbAm/zQXEzo78bx+ejLbTqDQ
P/mIrwuq8Uq0n/FE8z/332MZX/Mc8BM1zsV9eTG1qQczqnlo9XxQIbxSk/V5l55jNGULVgMN+X7B
R8JJK2B6GWHMbq+SwdQY0BYtvC/zAtuSAtl+gCkMlBvQdffEa/oDs//nHRZg1XF4bWBPGaRbu1jm
U1AfDwHziImyGq/jI4MVabKfUZVRyizhl7Bv38XRCQqMGVyc8yhrhutA1nYEPbEszYdEY+BHdOTQ
mi3em6IjTxDo9JmZjWb4+jr8n+edyxMqu4z1S6QMva2XYxtGcJRx5PQok2cPiKBafyW94mN0emta
hwat7tyJNjwhxSibF5OutFX8FkOLH8zwwf7Qkm7bpWFqejDnTVQCJ9EPNncSo09YzK++QlnvM7Y0
ghJhWVkuNLw9p3ySxM7lh12JW+xfynN44SsA6EUWKAZZfvT4RxMbHdg5z4w1QoOLPtbTKG7Yjnxu
PA7sfib70MqFc/WVXyzwt19a5i5iAckVXOs/plmDeYdoJKZ210KVMXipbreudvoXUmT+zoN4jDWJ
O6WizZ97s8kjsmbK9UyrYq+Y4reOwGvAfKm/Zxrq7Kul3rHH20iq0AHeiD4anoZdblDv/ZsOAZlD
nGDYWVKpKD5WArgsKK8Q3iX4wERG0/KFPUkw32Rq96Q0yXHt2mW7KwYsCg1X892pOkwE+04LuDdI
4NlUdHnire3xHvth4Lb2BuyKDtK7pDGLXKI8eu8B4YrmhSwZS9nliTmZJlFi0ozLwzzNHJwNH1+Q
73CwtFfSfZ5RvjR4RS03CN9Wo/m77HDwIYZeAKGqUgC+jC/4lThLw2dtwBGfxqlyKe9Iq7+iS7e6
3PzxqBfBq5Aw35vJm2AAE55kBcYtykyeeh43joi6mtg66i3le+IpxQlum9Osj+cU16fnQjuqSYF1
kiv2S6tf8IUIACH6wfFZHar/vbxmYfMVcAW2/TW2YXziSHjs+S2wwnTSOtNFxDht911fJm0W78Cd
aQ/Y5lgLX+wSxMDIFo9RlK7nfCXNyP/cY2ANoo61d/YJLgjzSRR302NRGsYspJM7gsj9N2hEkiEu
xJMW79vOwi+V+o6ylaRSzEs2w4vnqwqlnAESeZncHkCrKNnSPPFIZvQ+4XrvQZbU/U3yTL8h44Ao
jsUM9QlaKEDl/GeawYQyEh1nJ3v9R0a4S6XE+GNMxSO82AF1HtL9YsRAKFoVI9ZJxgjlW3Cj3lbZ
6pWXWC4m2KBknm/p/4QDYSbR4Q+r0TOnP3eEAa1t1bX3Y8dGzgvBLI6ThZ5WYNvc/zeFq276KzCm
ten2GOIyI+GwVBWUhRrvkdy8tlE/I/SdAutui1GRty3MCMNip60bL7BvPMPU1TR7C64A4jns34wO
mrD19fzckAs09REn9bgNtiVAoNRUaHlWsztsj2AKZrYeQen8be9uLFy13uxFXu/j7qq8IieAUZa2
BCW0XN5Bv2xt+jTea1TTyg8PEFMm/hP6o7pTM+695OFKRnLR9IZJWEHn24iNi6XucDSkBcjY/ZUV
Pof6B3JrdKKug6gi/qXi4/zLoJGakxW2tCE5r2cuqDPocvx/WSjc6r7hV5nn6NHku/16DBWNUOig
sHCz8aOXUGc6E/jYNy5lU3GRdn5majsk21w/0pEYO2WkHZSgNaEe7oteNc9QiKrZCzkzRn0+gqdl
oSq41uexXJ+oRIvBea1kNPKvIQBN1Y+77gqV43tsbDbvb0QckiQtWyRJx4zprLkmUqm7uMnyXCTG
n1b3xUFBOVm+PP4lL4fqtTw/y2q9rZ/o2e5xjuZBNrCNqkDCOVclraX4Ifi6AWv1lziOZDOW2FSF
W9PALTcViK/ltwiDENs04ZRJJ+UrGyteNi03tQG+ggDXaLhQTOvzyN+i/27kO82JRYn93DghKFtQ
OUGXzKRg+7NZw20xu8xnx2SHU0+uAg/eX8rtaOH2r912kn2HADKlVLvszE6Ib4skTsBUy4PCxyXr
iOA91piQ00m0wB9wAlqm0+vzE1zvWvbG03fAzz+L3ToQ0iUKhLlhjf0ENKNCNJMmge0eIxlUVA6s
N9u11YtuejFN4/idvqEfpu0vfCxsQF4FgqVXEsQJLfyDxTU3K5zyYqbJfxsZnhiafc1LpHISs9ql
eRmV8Kv+sCrO7DeDMIWtBAHAI1YdSYxkRcABNRclUmKSBEFScudVG/TvMMMXAfGbpbwdnrQ0PhYE
Sx44jRwBLf9jy7anhfEVhd8S9tYBJBPVe87rQTwFxYEnQ7Xgcmx6aDd9ZNEwaZXbH5XTmo/WpiQI
ys6bQ5z8SoBeQOMeYAJ5J7RtDUYfEuw+fQUq6JwCT/RpK4j5lgOaV4Qqi6+akSGlb+enTBxBIqQN
puruOLgX/AvtqdOyMXeQBzMSuh4LN5Uq7u+1eEAe0mZMF2l0SQNbe55RpN0k8u6707W8Ux+gDDKJ
/qDAepfdCgymkO7nODepfmfuMHp5IHmvQtr3Vj2BfYmM2j4cCmZg10ULZWIFqijqOwwq525MPRe2
xOcn2ll428Seksq3AKU7d3JwrrxLs2pfGvv3xI2SVOjH8iRf8acURbKfpyrkF/FOzUB4Nx59l96C
lna64OW04EPSlqR5vjCXxJfj+Udyw8dIwc3rh0xux8ZsSkAmXCbfpFQegxBk7u+b1+FFYtQ9F28I
tS3N9QM49gK5VnRcbmtBVPHlivawq/JV6DXF3RLuE2omKouZsnHLTqSoKPDehLHgqDhFqageV9nO
rajatQTxY3wm5xGIEgrJMW1XauwOF/8I90HI8G6R1iKDC7kAtmHIfifNI9hUq3QMqD6vaxZ+p1tA
U4IaXsmD9yu2RIGwdapAesViXu7kAad9Q1FZPIQE286RJwFpGzstYR1zJnNL9jCvjHh/pz2l9xFG
+0cZphHEpvYQpy3PW5qVECz+MuFn8bkhQA04qx9oEYwUzB/KlvnsldMlbsGTt2iDKvY/Vqzim8rc
IInXmoi82wn4T8g5ZHa9PHLOWYQS9eoSjdDQLauAN3LznYWqtj9oEVPyxbZylwEoGKz15XVpxct8
XicHgHUr9QsK12iRFU+einQtmC6UKPwi8IMlm3rjxLAzXo2+AEACO0AwUoxGEgYXRyQAvfqguSXQ
eDIppFH9/f7oNeuypv+yG4V/KOOqmmtySkhtygF+5RF6VHEADxiA6bMB7d6tK4XOdMgfkkAlvPAA
7WWKpOOLTYTTv91s0R+DQx38Z8fzzw+ga2mdzMKWZ8RMCcX4gF4Xs4IvLds4GULfzpr2tyXujpmZ
bDtm6/BV6fLd9iW0pacROMR5ycb5KKJ5MDywPqInJsDQ05nJFBQDsMibrmk2o1eU80eDH2jszygH
wOqXbLElc0UNkrGrQb5pbctk8u8Vo53ArGOFDLAwfdpp15NWgzi8PyNrAx9oUCBAS4OgaUkTaA+U
zC0i/YelbDATuoKkVd5Mej5/QmkV4mBLuGtncNjQkV1zCfIOqpmyfOqkOU+pncTa/6/2pcTA4XOy
2beYC2LpmwFBW2kH35qgUue4ADgLrzigDt1haZ9LodsdLUrDMvuXTLHUq2K7J1SsjtOL2/Z42i1A
hyq5B/kokoyDNVztLTkigtQg1CWvhc6qJ/mB92tK+hTig3JGMblbBW6M6TTHcDgDBlh3omqhskiY
85/TjFldr17xe3uCg985ga8VWZfI60TtOOSCzN08vhBX9OPtETipROFy3wXyliKtD62j7/yMcGFX
7iejq119ag9fmjZRszQ5Agu+JOtourk6bqHrSMm/FP1WwpZBoOZmSx+LyrRkmJI/MQhulVAMnzGY
zdPzvo+k3Savb7tucEGpi2JZ3ASu8dVK6YSitHLFi4Q+I3timqEFQyzCzQ7XoJc+glcr3cpfXg8C
lPmWzwHK/g71D/UK8fJHKpIe6DC2z11z5ClXYK61cTYEmwUZmH91z9hJiGgV4M5VWh9ZGu5JkpyV
Nirx/CyFzjYnxRDjdwEbMZQGY1mRofcaJtSUBEvAJavI25k2N0NDyTXRqPLkK1jtQib8orECT7o3
akqVLmvXVHT4XtIrEKRN4PdMI709Td8bRGXK36lipJQ1O31dkvQht7opcUgdhpayJxr37WOhIity
ePZLHk2FpSSiMV+Jil2wKZidKY3z6dFr+FaIF3EDChtOevTVAJxnQd3cWkzEQBv/oiTtvBpYhQTO
ksAKOTY/6O1D4RH8tpO75WSywJh5/9A7CqIJ+OMtcbaogzH1n6+/PqNgujxLAhCbRfnM5uUGhdZD
JRrNbBQR4dkAjvX6GP8vyynaa9SThSqXA2175q4MGM2DjwLxzsP5SoNcL2KWkuq/Z+1bgu8VT35t
5IuW70UzPOIugfYMkAzH+6A3qxG/KyZdlqfxFWhm9yijV5qBRZxRBSd71FZFd6VQDk4nAy71eeTd
1et/ik2deDmQx7l/44P95kALFMBFT0oCTIl7lzH63NkYbPIxMYgbSPQl9JNIodFQ9Vs5+0qQeMp/
ph5HFPIRBE/CXDvEoauJ4s9EeWJNWQWv7s7bg+MDIAXSCnP2a0w7h1Ynwz89uYoZFvFx48GyMZl6
45/LavJ+SrR6ihBc/3e/WCwlAe9bKk6wI0EbC318AmcytF/MUX/IhtiSpaxN12sO7dEW0BxaQ2wx
FZji2Gv0YmrimPx4I+IvUd+NBvtd6Frt9/jrpVFz6nv/Xsb46a7FfpqQQxRjHORlsKUqdhio1G/q
XiQV3AxVJckzKEuplJV2rTW40xKkiyUwFfrUEcEXbtVwDdZweLTGvAm9B7pGb5iXQnPR4RjOkemD
EYPToUOQcCqvpFypm3JkARTRwH6IkY8TfeNz4N7QaY+DM1h+/1+sUzE6yHFAJ/GYkcZtkJjlC38N
b0wqJi1vA01J6CcwKJsgm3kJ2xGA/s46LY2zBcfqqoWrrqLNiOB13Ed5IS1O6jC5JCBDcAlfyWIC
gOo+oiOzNDsC2ufSJG2o8tlJnn0rV/U0MNXT+Azc5KmaPF955qH+oJOgv0q4fGCHfa8KB772eCXr
oo87PXcuVtONMzwcxdXQK02G4WbZhrRvu9itGf5DlZKLwp9C8B1klzzPKshBMLUHnfOFVN7u5EtS
yo3BGm+yqw2UJK4dyQbHIyJgsIxOrBBuaPIaP459riE+vQ5Udj4PAHrF7LjrqFq2akbk3UOEQSlL
wunpWY6LxEev0vQUlzmV0GMGax6r3sd7GUu/1lSuwlJCJbOTGt9LWckpM2fn0AtTkr+FtWfX0nOm
p6gqW5cgpIZPpiMY3V2uqRYryWVGausUKSyiwcWOlYlyWqMcuZ59DxQ/MF5q5S/AhTVbDHyh0xkA
JlD9ZGLofLpyl6HedJez6BDGwwqzR5qkMndUP6MyZuI/1ItGqdJBOmpA0Sa8ITLUVzg+apw9klH8
v4y4S8vXY071cagzsqyU3V279sYrd8rkZZiYpjodqjFVBu5l8kuQxNgJ4Zudap06zryXtopQwgiL
CPVBjlCHysdJOgTZcGYri0k8CZEk/eGpmztDWr3iCmQpGdrDHgGXpV8LYeVh6e03vW4SUQNUABiz
yGgHcwfrOk2Mp2Kp0+/tsrst/jp/FopBeqv2B8AT4R6TFob9LA2FyawiloZtUWKkmMAPJWHBwNYM
s220UMw+q2T7pOKLmCQ8b0cAH2Mj2W1JKzvAFWktm+pJ5eCr5Cm2WzNcw7gxYeCNL12KEEYQWEBK
PfO7KiajGDmr/eSr/C9C0ykmbjdaRXVWUGieU7F7W4hXqouenivKG5b8zo9tUkK5GF5oaL2k4FkZ
s+FooRnphBSSra+47o+nozoyaNS/CfyBMk+qPYYxl+pUxd3OTE2UqBkQGrmPKRwaWz3MtSoL0YaV
s1AxKcwEVl7jskn6zAukH0Qj8eIJNUmBSJGotsuWIVWIXc8AX0Sa1xpBEMU6Ad3ca5LYnEE5W5Qn
a8t88nCJLYHZO6+isIj47jbiJD+8XlkAkiEZa8rZfsxcPrk6cH5nsFfpncB4Azmdspm/HR00d3RV
FUIsOYLIV/dHHkpqSxgcv5nfwX+DKqICf5AoUmpPe+WNt19ILjEA+0QSrmMk2SuW9xV8GOeIag5b
Tim3nBpgH3VFMiCsgKXWqP6NfI7DbTiNpb5I3AA2tXuH5HF7/0rIm28Y3IxMXRI30MNKX33gnAg8
6YTdyajOfNIK8VfIVucyfdhcqa8BZKuz42SdHpFOazLRTqRcjrycwEpHuBRhWbrPkugGh5SsH3Fs
9IsDZkxzDDgDEsgzQmcDBvdG19xWR2sl/I81MdTTLZQ3LfckMjaO3zrDIOB6z7ud3q2itbdfV0zl
5rjgsWEzElCAFymeqhY2UiWhpRzgk6ub1lqa9iNqdHOeXUFYMP5+Hoyh3oExZ5Daxdykll2OM2GN
0gAfoyM4bpbVw5dYOSRYqABvPHzicoWHuMa7kwNhqTosOSdXe1zZaWJgFIw6PAyuPsu25bMESzwx
7f+kOhnUjdZKOWfIoAtJPK6xTUkt72h4+KbBHURIg5uQHtGq3rI6hgZn/NOGWFzX0TFEICkxU6L7
pYpvR+Cr3g/5hiQxLmJSjo5sbC2KTaCtBlq0xcVcZBUOpayDKaLb53otf+0Y6l4LM4RAtpTOjq5l
YRTw5ytS7BcllT/YCSWPpsonzueKInnCeKhuUJvbyLantl8ULWWZYN2bSPZS0sV9TvzRN/Jzk8D8
342RCBhln6wiSRrts4dZVwa6n+CZqQioxpGncKQCmH4gnDS3wzseq5KGjUeu5N/nvFwpvkzcas70
DfZayRV9uGXgFKMB8DQMr0RM+DjoxLGYaC8Uy1F59/DTQoSNe3ZbdJwSmL0HWW220US05sXR9dDY
hYNoQ+8Vr24APm1SSLF/PP7gmNS+eMZHEe/dObwwkP7yEoiVOBw+igeeQdH5aR6NEqmUynoy+Huk
uWXb3sr95tX9YauIgvc8RiL6RJ002gxmdL5oyqv5Cl1r7rRpX0W1gycvz3A3rdUYyjhBZbur/UsM
HQp2fb9HFSpqODQHLmpwF/+G+TmRg4bslTao5fh8wBZCHVCfcAGhP3McR+lyaFAI9PsNrI04onMV
mxWqM9Dtr2vz0P3S5ZhC7eT9DoY+qMi3UTAKGc+rDzXmCeILA/cklEh0LBNkQp93C6RmyChTE48V
fLklmcjXSkvhULqSS5S1lHxKwJppDpfbc2svDCLCr43K21I9ca4eIMLCwiKb2eRHRqIays01NZtO
gLGPAr/TJkyawoBUcDq3HgpZH0924GPLIaE2Y35PH/4rp1FQVV3WiQzWLGnS3A+vKxk+JX7Mtd7H
fszUdksLoP6R4QElUHPxFIBM/A9zojJBbXITceyGcQMOdGKLWW8QqkjnAdW5PsDLR0j3z3qe6qR8
JirfplvMK+HfaQ0l+o7LxWAMSNR5XGVPyKDA2uInbFSa6Eh50+bnZYunXWeJSNxsbr7uUck4Ovdd
f0VyEmMDK5okYkPqIQzu/TsEHRz+HCkP5FOSKEux65ObY46UJmuPAIZ/k4m+GYEDwn6QH6ZOw/ZD
uPn/JM2cV9EGkpue0nBFuqkffB6+ppR9Z3SNNINrXIBnpoYmsqHLMi86Ij8ltoQPExiFR9bsjawa
3ROd6QeaoJZeKw+sOnzlx4OLbC3kviLSu2kg16qMIH3wM6yqDgxJWaZ5nHqnkcAssXppO/OoFMWm
G6J5pQ+rbFsMiBESG6yJVb+B69g2nE0rGlhUBkRxtbShlIu3TEVvHZQsWwi0az83l2zzOCBYewAi
Wp5ElEk8ivooYjcRtBsSikC/7CKSaFKWaNAhdMXZxDQ0tbZlBPSUnjo7xbuGIxurDt5IeHSOeib9
jjoJ71e9NYTgwrZkXq8LLcqWX3A3MjXpw1eCSWeMwyQJcdDMR/8UFXZ6WiWLhrJmdScF87Mql7e/
x2DHvJVDAojfrg+bPCUxeDOyYyIla/VfZCDGL8fWoRRc+dFbVFRO37E+gvJaqAzkfSU40sJHVbx7
Ap5Re8hQQRxlhDOh9Q5ppGtshCWWQaTJQJ5q8paFxa8vjqynyVQxyhZdfL9zzpStK/IdQ6oM4rN/
PW+ccsrGBvwpqim99BKQ9756EHjFsI1z6s85mnPDpFPlzekJYOOLpKY2dKVKccHoEg3kPByo48Yk
N9nc0ASNFMiCcwyK/Z6alIILuB65jCblbUkGmdoKpKfw+IefdyIRTVrO3kTKD3SQmMBRbNlQIfIC
Dl4n43GvEN2tNyR0BirDmkCDp7eCgU1T1YkKyQNQDbVmseteZwOX+Tb03eK+rUv4ICkCLa+7zVki
2OWQ/fVrRtBV9VO5Xpl7B26yKDmEG1XwnQVa9itwtxKJZFlMPOeiuNL1fF7FgCMQuv+laskqUZNv
f7Dreyq/gPmWNizVJY1u9ouLx2ACAB/Yp/hL4IajKcaBz+9DUgukjXpTeIOPgMpxqCRFlhYLo2ee
YNaBQqSV7QxedfqwVFg/2vy7sVfoyDo3iLxVDjpNzLJkB06fe4Y5sRdlNzuuSpE50XHM2GDg0XlG
fRR3fAXE5MXF52GCACOy4S7u0r+f6ca7KX+l56qy5ba7qFYBC8aFxGm91GbfMr+L+x6xo8XxdIxO
xj5twIRSodg5xxFuKX9wknOgW4sszvEn0Joz80l/qlH8Rw8n9mVxvn212g3HPEE7r+4T5uqfRngV
a+AGuI2sOAT/uuyVcgi5yBmoTCvRDLeFx8OiyNZ75KR4UKwb3gn+TlSuQJqMOqiUdmfjThr5x4+0
yl571HcwVv4uBbPGdxSXsJeQ6Q2gpmIsidj2sS7/Xns5LN7W5rH8fZwZPKOiVmK+KKudID80zghE
3H00Ny7mUwb//UH3XkulzCGXfhpEh70bAJ7woYyhWpQ7QWzliBrUf7EJPGRwyFzeoq4L/HClcqMw
YPdSyGyZEp43vbPUqxnys8Sm/ZczorWGWBKPV2uxudNLrKVlJReOSDR1+MwKUhpV5GgTsXQsBwsK
wmr/Xf79WBk+N8xhgUBOQPrI2RfkQlbX9ozODdkJ9OWB+d6ttSJo0kNF9KmdwTEPFnMLMfefWG6/
6zvfbqsXUs0au/cGhJi8h3ix64atdRGyBoNR4pT8PKV00oyKfQUn+J6VvXTBDAnLnIMVawnYXuHU
egIR34TLiwxbi2kQK7ylRdXcWTSm0L8PXqsSpRx7tpjEsO5WghQKX3lvlOeD7o1qmukEbLjafkKl
CoRIXiC3i+M+Wn0oUGbF+IWv2h+kTLgjhlG1Bi8s4lOwplo3Se0j3nTjBrWPE/Pc9mXO3O3C2SAw
iA6Yt+hn9kUpEL5ewFc6q8/GNcz+M5nGQ2ds41H09tnjCWAB1kmc+FXvWSwGvMO00/PCiy1Cu3Ad
B+37aqB077zwxdangQFyFUIeRsPBTMnsmllubsvGJ11TBio3PuR/fwO9RXD6QbirJaLncnSqe2ur
vzQ13w2nRuAc68kyyeOatSwD5v01YB0LdinIGQAphK5XU3dD0hEMATefCGsofnoSLxNX2gIqgYsU
Rgcg8ymI+zkSKXbw6q/IzJpkMR5Y4buwAy1BqKWUbobUG83+hdQuraoI0AB322qJHkeE5AcGYc8m
wO8oek2yukLCnJbMZveosBm57SZWvN2/noGvNJlvfqncIy/sr1vKw7dIWhaf1BCiNUTnkTP6Jdkn
9MzfNAJAVhlDKmdf3GgGwbrw+R0JTwQaC5ep6Ex562KEy45hlSfQZqWNHJyRpzY+kHRfLpLY1yxD
NmCdzjdr+2gbCIiHvNblKdMXaxHY+22onyv5QHUlIB1lI+YX4zOURxwKkW7hsHcQ+/24ifK5nPke
8xG+Sh5Nryqz6/1pab0J+OuYzO2u4O1ZftQGkNHq92St4COXauodPv/y0NE8c913+4rEhZIdemtF
I3gQTXj5Z6hOFp9cwoywsbgY9y/u6edClCHA2pz9yqXVgAREAX4cLy3vLDo/r6VhUotU4xSOisRs
Pe5qo8gjEIoBMiXWkFcM36Po5Ra7qu4mKEXNSx1W1XlqRWHm/5DWnqJ3EAaqe1bGcUkhQR5Hj2D8
61V3eiDMSGlBPVlTK+aH043RgUBn5APallzynFEkinLpoGv7ujZCHGZZ50jePS7euKN3Eg9LaTxD
5aOV5kqOS1GtbN4kv6y8ZuxUnRD7MVjLVfVkyj7n4eVGAsWkWqG2rgBYOiK4n+EbJufNPOiOlX0G
7O8L+Iz8UhVxuzc1XiEJ8F7t7XpUNQBn/fRU0+NwdxCnsqnxtUT033Jm18AE3CZdHEJPk+ZLrgaK
1nlscTysJkD+2k7ND9Mf2TpPYL9j+Ua8PBGAh/PNfozgZcjl3Hd1W25bhmTe6vBR4SrCZvuz+RlM
AHnyrj9znksaK0O8YlMLaSTH6Su92dxCbHmE3nNcCyBUUCiXyG+tfbQO7pQCRSNuVsCDuzRHynsq
Guf2gd6qmMsaDaDpkweUPQCQuuJhUyGFxaSW1FeqyNyaXrow1cRwALsPNt6Axs+D7NBG5k4+kfKn
xKVr4alLJTd8hLp9Uxe8AixXc17lzFir1RFgjv4kb/0gwDKpHodCrooVqv/kbcwj3YP08DdFtagD
N5GmnTPvDAJ/Sm93HHPSnfaNkYhHN2zX0apErUVvIFbat6YnXWil+FDPVnsmAV0nOD6Hf7qeCD+2
2Zdqq1ipO3PCnt/OYPZZnMrs5X4mdJRSKIW8alYP5NGMVIj56mbnNdxv9SV+JYGfBHByFCOAM3J5
MoJA3s2lUEi2EaAjY3570/xAltO/qLLwRwF2e38bnEGts9DnapyXGOzhFTOJMTcTEyMdWYOSg7Q6
S5O3bKE3UDwS4kGR39m/fJtxYnnoBtnBg6myATcbbBTyRDmPXc+3baECqeZYk7O2PTVlcsxojB1e
Sd/Mfm8EcdEK8iBLBr6gI0iEo8mYaWmN8licmPgEAUERDwi6dhEWe7zH132Gn1xbvt3UwR7ZNPx/
3vjPmRhXsxBM3rJVAAT+plpd3OSzx/Z6OqwcxLHOd/cUHY7ht4EysaVxtQFlBuvvZNVzD/2NeQt9
u4Ii+LDIxBm7VVwufDe+H/89cjqtMfkI560yBRrP8v0N4SEZvjDQRQW6K46O9flOs5kqi+BHYaj0
kdG8eQoDRFbJOstTKUQ6xCdRXXmV05tDgJLlx8gaIzHXcc8zKbbuw6Y08q70oa2982nS+0yl0C/N
V2QwsGl8ZNvjb+2vU2TUwfj+v60uL31x0LrRgyq9jjqPmBkgDrJP95CgEWgHNpq2NMFqbORjTqAw
ARFXuT8NrH8up681uRA898F9OAMy3ep0NWSQ7RK2X2mqrrxS6++M4MbHTfvbawt0p8cpKFVuCWKX
XWxFpqKVP8TLQ+XogoIKBlqWRPPl0bjdBqDEhPuZAe0v5x325ua9XwCn0yOCCTImh3qneZegYxPE
MdHisnvUBeReInoP0L8bs5ZhvELz7q5jEeLJ2i1C3K5h0j9qJGj1TV5VgyJHuDo8H+izqMoNue/y
wOhtn5Vmrw04M5EgoXjxPdvChrswJ6pdpmto8W6ziC+Y+JYl056+NfmkmM5EQqighGKpg490+Cqv
IgYlNGPcL7hZEJEv81AVScDYezljt52osUqKvDGKUciBjSQCxKFq3u9RkvPzZHJFM9OWAS5GZIPw
GpcZuaNha79O/84/QofO9weJsTMIdKyT/KhetJsY1yFZFLdWVv98WToEFQyQFkUrX3fc4Fv0cTnU
6fZRbYaeIdozykvv8ERRSsR+sVMCpWcx/LTahX9nxswZiQjmzMSQj32kwsmFNxyqWemVDlrTiq7f
MnlSM2/UIfGXlac5ng1KVKvt6Vw416E1pG3xXoJQldTkQeJ0n2R7bT5C2QYNYSOLjGTlcIM28xKd
d5Vyw8vxQMMFp5b750rIoMqGOBTMCod+tI2RXqC7F9srJVTwtpPeMgN5caKj5yM7LAE2Fkap9Xjo
D9mf1i1VdvoCPf2AQjsS79BJG3cpXKiLL66mua6T0h20lCi8ROpBdwN0/gDafMi3Pf4tZS1B/dZT
nw9liBpSEggHM4J/fGNMYGNJkVtVByeI5+oiWRyezY4rESLG2gmCIq/Qwg3tE4OIKeXHSsWTsaq7
AUTFC2Bn6DPDPmx3hVfM0YPnMAavpjuy+QA7MT87eiUzhmwSHszafATUrsIpJk96l6OS0u+tRVvc
OzdPipRDGyWRAW/LpZJtcTL255s0l+NA17DJ79BB8lc7Mh995omnT/9U7IVA67EdfsctFMBHa6Bl
VefHOfeBWDr89kCtWg0f2blYN4xjTf3KK+OqkVjXODbwAnsblHacsK5P6a+IKibSlswDSRsJSJJv
s3BhIvuyR0Mxa3O5t94uteTYkBhb1wLItpvIqB9sDTZY6mp1AcNe2o2Ri8/H+S6tpKzzr9oCxHYI
UEp6qCEl8vPmp8nDAztXAoYsMN+QdSDAuZvCtD3R3X2bVmhZGl+cbxfh0m7EF7mFNbzHszv+SlqZ
jxKZCiCp3pNnylxI1i0LMUu6qFtfZp8YNLwQ4S/wp0lxTEtF27DEhUOaEe5LreKcwZQ8wsBLhthx
2nAWagqv4fFJ2dM5ltjrNOPk0iLMf4n4BVpyFf3TjY0Ac2Q+ycKGUxWNGM5ujyNRyUvKV2L/f0MV
yvQv8p0VYOcfiruQ7oJROyIod0dadHs/vDHFDGatPqoJ82asDWqs/WTBw953U1V76Ni5V6ii8tXk
uzM1YgGavaHatTIKR1MguuFBJQ5wqL7jtp5Ne2a2/sRyPoxOVfMetU9U9BgI7EL9BYu9Q8VdFpb1
xqwJgyjkSHeAffoL3pcGOu3tvLqXW6Tduz3Fu1yDlBcueHVjBJhlxUQV3xfFN9fkrW4dCSDJ+2eW
/5AdG0OOwzPP9MdWo457W1qxp7rz3JFqGiFiPGRs7KKXR3eok+a4huDzO9UuihfVR9AjNBp4MFOA
cld/YEYhd5pYMyAox5+w+eTWxYgpQ67GUuSjlQ4LRiLLVciw9Yd3RY0+t2narDf1LBspEriw4TRr
AMOgymF7Y8zbMDH1w/FATSLq4clvR9PKN44JBpMnDyj2PHSL4wMDahau1I7ze9SO6HvY4zVge+Ss
Dzc4Cj/8pl+plpm0/ZvzLQkYAOJdFxXRB+NBbY2BcQvrRWm3592wPJwGcNt1d6YSdA3+huLUUxAk
YNrYxkEiMrMD6yb6kVc1i/5m0iqje9IwKoFcsr4F3p3o6XTiqZJCKqpD+8BLvuMV5KC7OzcAxqsg
R88uv2N1dBYkbTKuhFFt3HSh8JH4vIIOxFKT4FR7ZFUUUIBtsyd7LRwsFtojcAVKZJdL/j0xca6e
cmSiwE8wqXWPLRqW81aY7m6+pMVIEZs8R/iJyxNth8lrdKUbKBDXTkCLIa0kAAOhWkOCyzsWOeXo
cWE2nUyJCEiMn/iChxVWvOxXLr3PVJKMRhnrXtgpx0ieco8zjKijBmZk42zvJdbtEvJJIpAgiSoI
kZrhr3UE/E5A/skw2djpmL6kcepctJQ4FrEfDp6dH4PlrgdUOyQYCeartOs78zlxELWHT6ki9gjo
3jEiiIWHxYylUrpo/x25lDvWyqh4NgSOllkp/6Lp0VhTNryBe9mfXufaNYClY5dyiLAHd+h831HC
gnKdasji0taAANvyyG9Ju7gO8v4D2z7xVZpbrM8ijLVGGftE1J1vYiSO46H1XFsjWa1zrkw8g3HX
FMhzSIj5I1oGcS4cNjHy+MZNBx6xcHbHvowE3bD0MXop6ZfXXTNseRD6r+dKXk7nlBZNgeSDe/3O
nhsHSJa5RclMOwLCoAauxbStHf2DvrDCQPHpxrdch6oKHcLSW/gXegp+D7gEDQts6YcW2T/vNnES
mWE1QhRF+noGouvv7L6AfGCMc0YOwm9xZe/CIatUkQTuBUMN/f6t4Ka5pbqW8tvvA4As5K8Yl2r5
AXDWwFf6BPO+nD+GK2DnS6wAQyVKBchQn9JkOm1caE7yiGlpqhW6UvDUEfvBBksQmzWXXf7jdZPY
1h6QsIjJh6EnsU6GBG8vAST4zzT3SVPf/NWyabWV//Soz8pvTtWEWSReH/wGCv+UXyFLViB3/5PR
9ft5Gd00uJKsKpHh45SKKJ+V9WKUkY32pVxq4KEuScKgHaP9tCR4KT921d3pnBtO77edZA/4P2g3
MiFlTuVDXFUZ8NI70Uxdip65Zj16LSNfsuX70mPkkxRaZYYuYwUE+ji2ukbjXkW1vBmw5lhN0C/W
4Xt1p9i17i8eU52EQxjebw2datBLnTpUonn0YJYtViNdWUOzg80R7iETghfX9UUj2O/D3XePaeCz
/QHG3jK6+5LrmbiDJH1MO7sbfktLWyP7qmOSs6/nSdk8R2eG4rkwwLSk/VnS5p4fFnP3Nkkd9rhs
JpG1PYBpdlUuHrVtQ1U2UsRZ8xSzlJh2qbGjIUqphTGOgogIFsWw7HeOnvBLbtM33FRviovSJWna
pPXbsBBM7Tt41PpwHid2e9x/RduDmGXLN9IEO0AfFzcJGsdlplq3/2kMFBnw8K16oXbafVu+0KUD
Ww9Tbjd/Ed3PIje6pR8mbRHxLMf96L0JejqvBQQ8+ukCBWA1m1DIiRGpdZZYkiMhnoxPA32qJYzo
3Auxklb1HLJ8WY1bTW1qNQgZagZp5DS5IG+hILKPfAffqDgsHIOEuo5e11wVjn6nCvMMQSzx93ej
n1OqyH6Vh8dbpjFrv12saLGRx1vuN1swZC8RjkDr9doKlsnI6LrX/CXCho7omPj3qstaDiKk9Anh
FSC+4406+BFqAr0OpnnOqjm6u27XkZ6uLvzKndhdqc469OKLahsbB3vEiobEBC9BxBFRJNnhhNq9
nbcflAQrLJB30HnDQlBrjUP2xt7nZC0Br6VddQzP4jag3uQOMdGjqllDVTAl5nyZstHyGCq9qKlQ
3MM3ldxnyTCOR+8Xx5kh2EUmgIdXJCQFem6BpZmcVsgnct9Nl5vL7miXeFfwiAKlSGLhLhmPipLG
G7f0MUwESxFmM4Bb+c1SIBb0o7bCCrR2rTLxZpMcGC6YdUZjozzylA1RlcCNuRByYLA0UX+gZ8PH
XfqQENCVNO4XaR7O5BGRanP0gwLbb9iNLbvhhbKTnDfGhXQRjTSaVQlX2VhkEaKETYocNULiwJOP
UH35w3R7tGE9qrYe2AEuB9dhEyKR7AfMCsudHd68c6Pcv5EZJJar33DDp4DSKfdWSvgLPzZZvJCT
GPzrnxdux6IaMi2f0zI5URHqYiMCQo8LdjtuObNbsqeqICiFNoOgDfwxQ9oICvg3N+/M+l3ZY2i2
NXZFiR8jMZ+Gk3HEM88YSNEebHmpg9EJFtbsJE/gxI3Wg+k9u+aZxQ0Z/grA3x2p9yfRnA3wCfj4
yzaTbAjjgIhgZCj1yeoeacFAXhsf519InSiNHTvH2vTqalSaD5OCHjs1aGKB3w32jiROiiMuh1Xh
B3iTj6/j8BHJ2q2PZ6oYBgUoeazehLqa9PQMpjWKlxUATQnEyoIAWo8EdNO6y3FO7/keR0XgIqXl
aA2wcpo4/3y/F4CB8j0tKSfGBCacFFaXp1WWzP+l/sOG5N0STIK+9Q6g+q8HxfbA4NBFRcdzYvjH
OOK2DodOGAADG1HSj0uPNrU+EP+6pDlMYuIvyQEzhpMAkDh3ATxNssKp73NS8MzYIzNUvXOJSJpt
t+Yu2WqHnTgnoswbNklwSeN3Nyhy5tvf/11QyhYzBDGsgQXNB2fubSsVpYNM71ZIa6cmsDDco7pF
m4k8mzSV5hZleXi8Ogz7dK8l1kGPdpCfLIPKKH2ORc8nbSg2yLMEwnNn6U7JQ2HHcAFglRns+/Qn
ULJfFhN7dZbF7W6Kjbs8x2iPPibf2Mz0Dl5jtLlRV0CrosoAHQjjmQLrpSxbSnnSGOUFK5KTt9m5
+hvt0vodVIZviDUtM/MGt3OQ3nhMSzAg5yrvZGfQw95aGKEPj0xplbOImayro14k3wAwzvFk0BrR
1xIvTOUB5OMRxS2+fhUdbVO5F+ksuCve4IGNDTf6X+vDFyIi1d5sNiOJBqpZAHrzQy4qzK2UKCU6
9/6ZU+skkSPYNkLJd7EoSxFYqPJf1DvvOXo5H5/x+Ang9xfjOe02CGeI5h8vTwVPpUi8rSiLcRdn
N7E+99iX2ws2vujQQWgRseQAHI10VGI57+leys7wh2oKVMoNvaMKN0T1buJVHu3AbT6hYb/wKdV8
GyJRkEDm4Bef4eh81uGecwYGbaZ2F5tnha5MvSODSuNTCHMQV6gzoVKZBCDIRnKWY0UXZqckMCm2
UFzO7BmMpbGo6r/vMWGbZF0X1SwRJ80hL0HHZoDuHK01rOGob5Ftn+mboYcRa2oBNaISwJsqWKlS
0vuC8a3fVQiV795VCaEaY3T7tWUpLkOEBC4eWQmz8y0Jz30fJBrMPBuX8z8Ta3WbmkYW9gV4LhMr
7O0MIphAr5wLMvcE+r+OjMup52hSGLePDiIFK0CsY7BqfarhHYo/Eqc1lse4qfFDK0pU+DVeuVet
OWXnToddwziEGa2VeW1rGKRPNs26ppNRp3Xn4git2WnZIH1Z1zUzBtSWdJfNtzhV8fHhS4McJAIX
Ju1KE0/JfiWMS2ogcS+FQww0safB+xG/p6u3mzysJmW7sB3rop/ymZbBQB80Awg/fsS2BYZr2ti0
djiVUxzsMV8uGMt9auM+1gBULHlmYKQU8C7hwDXoJeaGr18d3Da8CfKvYe9g2/03YHfdfh7TtUNW
oybb9mJ6clI1pYz1JqRqxmz8p33TIWMpsrnTtPYB4MMauH0nw3AwX2ejw2XzfRpFUEtul8GMVkJH
sh4syufVNEIw39SBHaNlB3u2aAPsG9VfSlkk/+fzT004uCsVHlADaME926PBxXe1c4RhSqwTiQIO
Qg236JW3+3B9YXvacBqOi7J+jPYeAh4i49arXRILinUYPuSVO/nDbr7cFqBvxgPzqfrI9ejEPCdj
2La0mP0qfRUIVXlzCD1mLNAUtR46vaBTlcY8DbhsH/B0vjlYWEAAFmhoaPrf+ixuiejkm+vKavw9
KNuXIoPZlf+i5WjtzczG4eT0lCoVqWHrjsvcVyT/XhlKtVjIBw12oBoJr6Ti/waEG7FveYWX9wVs
C40ZWUr1MtpTaH8nqRh4DuGDc+LUyq+lHSeAMDRBoGblpQVqYVfO6Rfk/Hy9R8vsGYEMezIIij7w
HCDSlJVLJaJbt9JTVWjqlDDX8USNtBXvmK37DTplxDXCeqGnNYGU/z/EhecZK6E7GkckB6kO1xkR
ckUvkYkJH15SrQugMHcyB1PxWAQYmEzqzZbOgs32TMMZmwc5XgRv7uNBBGz77GFoBpuRNIiEHwy6
6up79HkN6BCZp/G3xQbvgDmNzwEPalvOWuX1W6ZO63HfsI1g3xonHtKjoSSrPFDcjTYmkFHUBHB0
7qABRfdMBcAvbteReZfWIJxggHoMDdQVf0JdSpodyW5EsU5yqJlv56g0b+I9eJH+3A8l/B0BTUDO
sfIPBsR02vW3FERlCqp8AGFolIJ0gEhXmyJHgcMxfQfIM3eP04uzzjq8Bo3cNEq1No0hQHcRluho
mVfc76uSjdUGanXJwLPkNPclTaVfR9kxtQ++wEEV7T+A53feQ/OOytRs1eE9hzqJuSftyhXQK2W8
ABsVUxAj2CHyVi2G2wmXz3Cua5cKyVqvJyOn/tkm+f+fxiOldXgth8AMIIR3nHJd0eUXTjiQZA2J
TYwZyDwonEwKHmNszljs5wvhTU3TzI0ZGaZWWWXXrwNDgIpStBlVBCyEs3hjrsuNJ+HOIfH4II8n
OWHdZrtDWLMsFEgZK76pxpUy/BHPOQcmdn3h/152AgAmMIlh09wDsnVP1e+bt9YTq6U5Qq6zCiq3
BNshhDDaSlGS64rOeQRwA2C2+DzGVFS+MRqyhKz0XCYY06V7tgWmmTSf3KV/aORfI1bMSwa+6DRn
QGebVLbXatniEkXBCn0t/cyeZOgSBJ4zlfXxKuWxV944m+4ULNrucnc6AUJqNDbrquIY664wNjLE
uPP4PHHEarBCOFGAdPjB40NMWE4BWdbic9pvdNeoDhtYDlY5NFOuLHzJw6zhII+knE+jdwonOkDj
KqvD2r28C4Q1vWVISdt+0Sw2pYXoxryDWFz7eRmoQdmihe1kYICVX5i5b7p7ilB3S4NwCTkwtdqT
vKsFvW3zuObnlfydUAbOFtJey1ouH0zXuK38fMxQpFrEmaeVXfrnqQdIwMqz7pVngYRB9qGJt2ES
D/svU9Znetol+TU/ENqjheFcUUIFSECKb4Hhmdhoilncys22NfLBCv2BxDiH6VKugEjiSt84/MNb
cKdMkyFXygNPYQX9yiEXJicGOed/2OnXlgN0MHRRQVf+RF6khTfHBEaDWQ2qujSoyfciBcset45T
xq0qPENboGUlT1A0dHrbi6Npm/AaOqNIVqrX4DQQiapBLQvNTdsju6fpzs6PejQP7hoc/7hnX/ZO
mbz7pDS/ZKeDEEi8ym0BUgWNNF6Yfo8ETEC5ws/WY3ybAd/E8C+314PffpTbg4DE7GRNcEmXWrUi
5MJ+yphGDC90UnSIabKOA66JlTQwCfGZvVvw/HVguw+LbiPClVD3jh8Nafwl0t4qLWKPEFvlcfiJ
9Ex1m9JlgnxFODscEtMC1R+ptK65oseHX+SOxC5kT98VMVdJkFvB74ZkUiqykJyNkYYXofJaf1it
YE5R7bc0vJQ8/gFhniZ1x98MzyL0sdrsHLlFKyBrnB3WdhaQMQV78VxZ19fis7rmsiAF0FoVWp2N
nLNhtPCYXtCbbz2CYmpyJ46/W7kqAO1tFo+ZaRV8WTkKX1Am97BHA5rTzwFPPd5NnC0GdQv43ED6
LkSzk85mmnP2KQLJiJx5EZFGPUfN6e8uiJIkGelV6QCzvjVfw4uQQtRt6C/sDNIS57uVFWvxvQ9a
FyzPQPjeSxm1Dyvdf3InLtcuKo4Tj02N1TqXAGwFMNMJH3IzOus4O2Pi7/T32rnLAnzoJN4OuHYZ
KbGb805wYcL6hNUSv0BNtp3gKQJvIUvC6yRYsaQP/hb1552K+2VlXKgTYoegDbQFVvCIbG5xprzE
6RM17PKjQ9mMo9fL9oEzhR55DUU1DqQN8/SWcb8xPcde2JXJ9nyeGM4JYkZxyESYZ8lHKe0YOJA7
CxAYtMWrKanhL4K7DLUDABz98LYuER1/kqU+g6KXgxBvOu+VlqLNClUverYe/6ZHOCYBz8nTW1Fg
DKZYDSqS43tj5E9Vr2Ez0woLyy5W5Vks1QsS/kGLNCnaN9zKKw42LpIhndO1LMMkBV93I1DJ2ga3
JN9WZq295eaez+oQUKqyyvRZEYRxXL1gdGVSs+Y0/ONy9FOUuYFuRAD0tlQzkmiaxGe7gjhHQDpx
6T89ts5PRPTlXbbDI8iWuuYW0PZ9UpiuhoVamS+fyaDdYCJqAYvRSvz4T3oV/vIQyTwYX8DN0isc
XKtE32DJCCXmBOirHumw+E929AI4cl3iuRvl+xHSoouKl5ExxYk6wArGBoBSkBorAyLhqCNN1N8y
B3+g7PCX2sksY10cem/RHBrkYHfPupMLEUggxqza0FQO66NYzoYqVtUVHX5vjtIDIGHQnE+RyBKb
bV0Wk15oT5NBd5jXu11Y5lcFvpdZ6L/Oiz8zjMTIj95S4i9OVGb7dM6HTWyWNiqPbX5owm0ao5Xy
Av2clhtEsEQ6d04fUVO80o84nymgdWSCoFoZdjaGRyALs5eIKOUvyZGRkQdly7moFOMR3oiT3L1n
UrVcw4dbQcy6r0QPxpDTX556p5XvVvHexl51J+an4veoDgY38T7CYCfnt1PHXcdISifeg6/B8TxF
3/UvcV4z1m2/5idOmX4bunBNnRIwZfaRU6cvc33JeS93ujJvBh5tEZgKp4t0zaX7TUaXe+WHrqsP
9jaOsBJ0PY1aODFX9SLJ6P2uKvvTTLaVrc31SCJQjVdBUE93TK7jAMqw7gEfl45ecpzUXKrTn6OZ
KXId42epvknfniJMcj7zHY7fNN3atCuFw50dCAd2+EO9N934l5Fe9i6c71qw5IQwfyaLkggsttzk
z2TdiCnWOMOQxq7g1+zRyu6mXiKxleLCN8xJaL+E93y4xlY4sm0cAgi3DuTEX/AAaoZ+5fdQdVyt
mKMBtFfv4lgYvxkQZQJBNMR6UU+w0dDF+Q8etcyF6T2JiZAiX3IpZyaPr8eITit13MEOYQ0gEg6+
e5yhZeGafyBPBYYeX9lAzKurf+Cz0qdyZyUJpbTabIx9CIn8mYk+bz+ghBxOc8UrPFcJRar9RE1r
rj9wHDUW7UMC9rchzAXmwQScmPhFsXQZgI5yhAebKUeewcyaNa8Pyri6PZdBML+ixhmUsaOPIFla
J3QS3S6xars79f2GUZxvR66++8uERRtRATw2MIOg1UhUrNfvomQyp3HE5Q7YEBqg3jDbVx47j0ON
qP5qLCt0s3Y4FiH/x66N1RWHUZxVNzaue5x+GkWdVPkcR2+JfeePZ3LH98IyZCxNvs15iVItdDW+
caX6IuaSyobA9PhpOHwMDIuJuLFCkrd2Rbia9N1jUrbxEFC1GMbLsFa1Jl6FVOWLedjwn6hR4Tkh
xuHUGVXKoKTC8ABKBQKlaqBw8ksKZKSsg3xMlnqfkeCxfBn55F4Rm9unPbge+hhkb5hqGYFATntD
0/3LBYT8eXvbDSL98YW8tNazYnTvdzOdi+F6xYe4n/2ruqbU2HKGXxE5zWvaLDKHqYMIaJIPqfVY
aZ/IddM7ttCYxhYfZzi9xuWfSRt3OX4kggl0zLSh+r5BQz/vKnYbdLyJEqUvdBxIiHFZ4wbK+2rT
G/RYSKTSgscMdW8hBXb0JNpQGzRMvXNRDCEPxytMqtayyQ9m86ap1WJsREMtRwrIPeqk1M+CuxEo
lOsuuYcfWq+d9iun5VmnPQO7osvTI3bi8M3Puys2IecB2SYLx1CDwjFiLueOM1tymL0WMwtx7Dzy
TwTqxJNsZICb7IC3PL8HXiz2qDwfdvfPVWpteNWUE/DWoWny2DEIt6sOxy/FR7bEwneFFruHV/88
kDHOyY+8y+p7lqytqx1N3j0OCPpCSsrzZhravW8ows3mJgbXgmsY+kw8gqMM1cdHaE6oLdn1vQ22
DBajhvYSUINJUHVDjRYmQTuNkTuxM+Jgyw1ql74nry274hhxYbk6blQc/YoXqD+hwSp13HkBigNs
04TD/oDzk2y16c+k3+Nxr9XDACL3Ae44LrXUWD0B26y+F3dS4H90gWQSAMKLtyBsWGxm28+rZls1
/RoirLTpqVOKFB4o5fZWYhF8ty0vq1LdFUFQfgGWvnVFMgaqaURsWovFlnmbVrkeV8La5p1y0dpl
T9En3Tl969R4mtn1/aDOW98a0tVAfAmmiyHxwdEr/l+8fF6v20WQ0DqlVunP2YiY9+sLR3wLI6Ym
bE5oauSyeI6fesgdnC4HADW/v9sgKCC+fxcdvUdoczPH2+yYBfVrrF3HaheKpM8SgAZdjz28VhT1
osWWbXUm1l28oOQuw+RoIGm2zkOswMkN4daJRIkD63OPklme1FHUOpNLQAZwl1VuXGgww5AkqVYN
Ic3S4ce1UYrrlylSxIPjjowLVXgDQ/Lt0d8h2ZnrOnXWhFJklkBQNj4Wn9lIgPmBdoF4paxO9OTO
H8DSFu8r2K2MZIYJ1RMBY+S7kNyrcaq+PcGI3AMZLey1vOduFU6OkPO53+MxXQqusd/eDZJfGYm4
kN2Qb3vckFa3FSVzoTy6t8TDARQMcLYRaIuybnfA4Y9Pwwlki8wo/auoLIXr+x5oW5SP9zLaco51
Xt6mI7ZYCsKMSGlpFMUcbn4cTZsauaUJjAAbjt4suuVFz3mTMvu61O689QJkpV3saOouUJfC1tpp
h13AVzPAij1by7zGno8hm5cn/SIlFtXbIA1rCIyHa6ROJSsMxZGZDLIfpZpruYDRY5IaqTFlE/F9
kzAzvTmy8DZiRQs6Kog/KgNbhgnnSDTF2Q36FaLeiPiEdYlmxGQmlnZPU1DYPypTPLIKTTborH8o
364rj4P/pRe9dEjqXlYsADSSVOW8f2YcscNUbX9afoVk8ySLYVpayoksEWTJyzOAUTyLm6XIiWvp
jVu2n9n8q5Gbbw5tkXljYEjkWSQNivatfv4IkFaiAH5Bm0wiFemIr+/SbltDM2mY6VphrINOHEXh
wAJ3M0vwgggxv/xqDPFkHCxdWmEU6weZ/QQ92SBWkuCVI05EBbQAd/aDzXKxhPDna+ZvA0P3l+Vg
4vU36p5lFEr4aOEzP36pJPxVmzCLCwfDoPKZacDrignMRozrf/1XZSbcFTLWEI7snY66UzwdSZEx
5KT0QlRICDviiir8YLAARgx78n+PnExxWnDgb0LOvSCJyAXpAd5J6i/7KszxB95hA79w6t1WvxAb
lGOvcamUGh15GYiyRVdSJnKQjnw7nVy8WbThlkOMOuUF0i27TCQFqhABX0bmIHsU22zmZ7tt95xI
oVcWNMjaeB7Unva5VASR1Y1LmhU7XLkhD8K7rIuEsTBG/JloEHxX6l9wxmqbv1N8zwtJHvNnqj91
SRAFq33Xm1Dvt2mrqBhCefLh5uqY49YUznydQjRwn/ZS5ct0OGmx//Wnc3a9pEdHEacEVFegMJdo
LLzoiE9IxS2TVI3nlOaPY0On6hTDFDdyAGO0mbhe9JWFe3IsWJkC7MvKy978jvUa1VFdpn47QiYo
l0RdecY0UcXqf/awMPxhBxbcdvZkT3Ys9Ybf/U79hy6vmr5Drq3/u5B5FHnW31RVCoFsKgIddTW9
57WLQJVsM/b7VAou1t0wjkWCEIFnYr0i9emaoMaJeVhPfDQVqYSIElzK5B/HGG2T68ColerVsOMh
58uxbfVDJtNYE+4j7xB7IXzKt7/r77sqmX3RGjrRa0/jS6lDsknQioENoFbRl++/Ws4pxnloU1Mv
qHrqIr20p9mZdaF+ONmhNC4HHXEZji2B23UETkV+FvwIGj1Vgi8W98bXea9RqUHDoYhlhAtvbmDB
UKFmRHWOExUYUHsQ4Jdy4KinbFb8Qv5LULRe2QIhcqy++mRQ3LpNIIpv0STJJQ7RrAPDiqpTe0cS
yV6MEYEcE11DVdJs5R4yw4xbUec5P/ke9sZMUWRu9dTdFwgod5QmocUS9k4qQVabJOR/Uj2Omy4r
bkXGAi3XwQpBmvG5X6hYW/PEqAv96Nf4ihTsNE0OhirVyaoo+ipMgkXAESimr68we3SRJfY7gC8N
tjNselEfXdw45OgZCgKljxOt9fZRw02u4OHKL+4SxogoVMW4cWIaJCFIXk/I6FCJa93jwWb8JLzw
QBfcGzzPano7+KnzZUzmVHDxl7+BE2dvusN7A/fPfJBbNHYtCGNxfyP92toL9reVTp3JynGvHIEM
Ugjh+366NssDmVb+HyRorG2FYkrd4vmCalJ/FYcUeUYM0KVVkjZoV0f6ETqKOX/1vNzX5RQInmvk
wzqhEnQdPTaoReZReM2gUy3AiTdSiy7tA5JMp4x9kc2AzkWiVrigsg3YnenstoTxuQq0kXPRglKc
V5xRJzGpTarAjBzaElL4B7vwdP43ETcaxmXGt4psuWAZcrqTf6r1YhfD4vvxUyvNXBimiWiBQj9Y
xRzO3DInXD2t7+P6+KeXbp4ZJFXj4Z6ldMLSBWibUCBs+pWlqBdo+V6I7U6TJS2bxRRWgEQ03ORW
WKxix2tRmZfFvF++a8TBS1wu7w9Kl0XAgy7E2ih/0HLFFAMn8omIToGfdDmtTeX+JV1Zj9zWGID0
fvYDKA3ryER2hyJm2M6ciCyqcDtB4MxrG9pHcV+23lr2WzfIyhWCj4O4MEUL1fNGsq/AG5WCEv2T
lxSYWPxQltOivugK50NfQW2LAiwVUjmbF5bkab4uPOtLk1Gu72XyB5lqaLKv9rNVubDrXn2sPZGV
azW5HdWTKCbZB0FQhi1S/6QszZqPmAzc1wvSY2n+75tTUR1lqSD7qHLmZKMCI27Hm9fELbVhia0r
NEV2l/zg4AKHpQnXz7ab4brami6XYJWI6UFU+lNwURcweWjfLkYPm5AlolWyuwSsgHhD3usAmQUt
C0pzb5DVNrpuyg42wADReG8TJuJDzBPaNxGcw1U61fzQJg6tQauHGevhwrv9POWhoFtMg+YWwgse
XqrxHyIekMGeWv+5akWF87QJZN71/V8lAyiyQJr1N5iEe/bN59woqMhYsMjQ5ptcNLHRfteZPe3a
S8aT6iqtSaLtLMZgDlrYTH1VbqAutUB79YK69UNYvAnJOqCLvtHe/9X+/OkCrRNyLimn0GTvptYw
sO++YV2BRkKu8pkR0ZwIVJjI1BX67XN3YgR5lvcRi7PCWNTGKbvhzZQZA2mSckPi70K4JWVdoA09
FQSubB3FZc7FjFlmwSSwWyKcRM59PdrQtvgoW0gxlZJbYXkCsXV/qUXVO/EE7TykJe+TrxjGtlEc
JdPD1qSNCpWGK44e/naiEQ0sJ93uC9KTvic9bVcRBY5SkBANgg3P8VEOhua8ajJXXpN2hmu9JcD3
KCRkInRSd7JOJLT1bj0z9N7UxD/yO/TUOwTl8rgYFzSSo16Ni6icz6geZTcAJt46DOUoGL2I6YXQ
Mkosd6A+hpRxIgFBZrht0JesZdKkE0HM8jgiAuygFqTjxZ/Y+8gRzs0K1TimxXPgcGaCG6RgBdfM
vtba2fCLPOdj4CQrM0+TsyZwhUnMZSkQzxNIecuUgYgs2gO9knPNMsuOlm4aZN4cx3zqOwpTEF9u
nOl4eslnCkh2w43/pMGzjBDHB5BicEVsc7jNdqGD7pXjYSzSCTC4dk/TmBhXwSVW/umPVNjX+E3Y
dn+HWhcKsuOA+ZpXZGV9CQ4/3FF1xmJs/d6fTD8koBZkzg+HWNRh6rrOqeFiSVdCHU5oMKJUq/D8
/etmwdLiEh1I+OzkyCval+QX35gcd7HAdK54y+BI1gHsd87Fe3xKMsTIx3VzR8M9Z+Mv/4fsttzx
CXGCwaqRyYDUiJP7MgtWFn972l5uh8lMy1o8LDklE9T76YpdA7kFJPyxfV89UG5jJ1npJHTYEfUk
UFfi3/VDOiz3ykyw9ZrbQpX7/FPGnIDFdoCogL9KVpD/B3wDoIrgKwypwgWQ9dxd9YRBrn37q+6A
wAew7ASQOVr7jFVpkTWK5OyLPa0MpxpGuo1O8flKxadSHiJpMHZmcUEWNOSOr4+WtB/TScsFQa3t
zy0G+x5UplntKn1vKDKL8JiU1+nUxHQzOXFsRyUCoLGsuJcjYq0vKJ+moTeki6pIfN7m2V5CysBv
Ya8PC0zfikK+nluxwn6xphO5XkkHo/1CW9Rva4g2B69htBb9OrBVlYJeFiWUakg4wtVjiprxbGgV
D+qUp5AaTFsp0p4GF2dE6ZENDuF/in9Vtqsv7lodDYgBy5S0KnineoKxeJIihBi6UAr8rsLMGGim
mKAzLIXLVWdqDEGHo2EbdWMZr6w56okwNuGXz4/2GsACyDvPnlhox5Nriv5UXT0cYVmr/zeNaMvw
av1FvUtGOqzFMYYQSppLraMlYk0MzBaRDc5yP499rMQoN02lP2Cna6yMPj5tS+jIqo0GcDm5CYdG
GvJ2uMyffMJ+g0M9GiIVAGfhpJ77rcelz+6epWaUJ/rpqxD8b3usGljs+ipoaO29eXitV5Eo2rI+
CUT2FpLhjbq8hZG/rd5ICQ1ZYIlY3F1NxjZp04U4n4a5AXcIxzv/+1fcmiRghLavOV5y6CDDkN6N
X+pLdJbqAH+mIYhzcGUGDEpIBZaoegOh4nO08kVX44NP7McA+qh1JMDDP7gIoSGXv2c79Fdp/8l3
Ne2LonEp0ZAcqcZfhpDH0AFMv34uPql9EI47maAjZEWLo/DpDZu6rpP3SRkF6gJZ/0uNH3h97F7X
e65sCi/ahurrOx8PY+DaKAbkJr3WAuObonj4P6YzRaJwM4UOLGzs+20nv4Lz1jL/RUkMWDDLGZ4D
GIMWaXqq6ip8UL+E6OIFWTlBNnTmzQ5SbCYRKSEVu8cSM8QRBIAiCNTVSEIYFVLe4VZO1Y+uBtY4
8AtoIrhYvqRKOZCQgoInuA5thU3YookH5u7ecdoGEWv8hHRjc/B+rRXP/dHbkfKaroXsmL62eq05
eDUTwso/X2AEn0OcpNCujKk0vdZlxLRoamvimiyyanl31GM3cQCtFuRtubQzKaG36QeJrnsm74yp
6cvzHExi055Rl2nniG2zq33/cxi3R/JeMsdxwzWfoNCxqKjazXIj3WUj9VXQBSgVUVpkTmWsfZUc
ENGfFHhaTf4Ip5jhlTRy8G458RG+Qr0b+jFY6unTWYjx5hiQcPoUfS6N4Kq+ut79udT1KTMKdcjr
pioy4Gggz1qmLIN+/vsjW6BA+KOAwtZ1d1APIqGULc0GQZCjv4U9IL5jgEZuQnCnlKzZea47n+Tb
Ap+P8yS1wBl/Dv3odi4PoFWmTfVruJdF7x0+WQ3o7U9W00vr3g7awzecpoT+PSgktccd5pe6iA2c
n9P2aiUL7fCBdbjyvRLzd6xlnLE3u9epeJ/KhXYJbW1Olzg4CL1qbOXV63nJmd0klBuWhMJfjZwv
Wf0llBYcyjB3HG35j8vFMva8AauCZfqkSLDzOWSuMaVRyaEqUp6j1oLnUaiArLILO9KtKRJ20eqF
eLAftoKUeXCSE9XcBMBUBmc5oCEt2WITWL7l3rVO8Ozk5cfidU8jubkXTP3klhcxUOK8oOpJMH6J
Zbx0mWFEeHCnPnizKOdS6TxGVJGY2c3NsNoN3AvgYcIFaJ6Tfy4uksBk1i+qu/5wTbTbUj7+9eD5
HyWK9/KUrS5ns+eOEzsB+2/tVmEaHKinnogG0QGrZZ37shbNw0UbIN8+xg8Z+RhqgdwTWYVDfKrK
fN5u0bME0gB1uAF5mgCUsQXvAW1fitkAVJnwIC3C6Sj+0+kRbYEC4NjcN+TeHcCj/58OF4SrtloJ
ojAVb0IF07YsTP8d9YtL3R5i8pN85Pks9NaxUA5cq4uAc0bmcrFe0D3Rd4oF5DQuCJYq98Y33/da
HRxYlKnKPa6+dJU3IoQY420sct0t3bJ0Gz4ECz6PbsRsmxpZaloZ4k30+IAwcR/uWLJqf/0JTT/t
wW0IMQu1P/0qBhnAtNo7YAkAGVM/gVdo3c7ZXIUVdy9zb6eZR/mZCL9CkHfcn7m/aPDuoLTNuvew
TI7bUkWhAN9ruNCljZ1yFoKcm3a5PVgAcP/G/jnVimmB67ulVg315SRp1jiIqmMJ4DOUe05hpS4d
JtrhKprb5T7AuvJUQJzVmZVB1ONy64dUajJV8knrxR8fOt7Os3v3s3ke6mwdnOPFdhUD64B9ul6H
x6lxQ7AXwxR2N0OY1MWe0aRI0Fg/Dfat2tOV4r90CkSuWG3kwmniviQUzSuspinkxE0/OIdSqf0+
LDpNN2KlIQu2iKkcG7CCPSrZ195E4FywYmjRFMwxC6g3Ob5lxr1bL6hpNm9vu5+pqIa3/EO1oppn
lRD2CpOZE1tbcfjOGKICTbJiqLrsOJeK4OHLmieDokUeCNZ/sgnNet49Fjr5jqgGeCtrXbWEaQIe
xmmbLA7QHR2WpHeipulEhvV3el+5juP6dIPuRtPBYvYwmZhJlDDggxL4C246s3Y3qTeBPbgUVVbW
6YPJnjKaXp4jw1PCA3xTV0btrVYgoB4P4wFhQSB2n49Y7OP3iixpQJqtHBBqHFH7bysm3PGQwjoj
b61ycWAMnD2Md7i2Un+As7GXG9+/oZXAVdmJDMB0095tslhHKVjytQOubK7lDZw+9pZ52k/DkDxX
WQYdgaDlOtHhWrA536gYL0JBjN/qYL/oJ7SO2ViF92tyumMYmTCjBC87MKeiS8WXOuAbLM7VsoOr
yJXLKQ3CptyKi+ZnSip3pPQDoq1oggtc9l7dy9aD0fVk6oES5A9REkqvIjhpiZQReF/IhShnIwr/
jQi5bzJWVEHQQoq6zxNMQ9fhkgA9GDhlbcCk/EzkMTSCG5BLnEdCW6C+BPvnMPQO+NVH4vdbCmNa
KM2Uzcy7TBqUoASHA7bXmVym7+EoA9yZEpuTZa4JfdQHHLYpFCvddEEiWayjLSgZ46+PzXQwkaTm
S7d0iLKa21yyQ8WKgJMLz3TbFNTM+JPylj9Nd4HPofaL9sh5Dgz1Xsnqtxp2AfIF6aT2fG9J+FHm
9X4acjRKmAl/TMSDI2+XXztXinIEg/dRuqf0dTAPy6eOe8XfTC8pNZRkuiwjOKTbnM0L0HDhuN/Q
qdjCilTm2Zx8cpyWKmo15+RKzNdg2Y8gsEz1bk55waOOoOG96C1r2FcvjuIJIQo+gXMIC/ZMj/iX
i6ANv0G9kJ5HUbwIAwqVAqK/QIKEBnA3FqxXpw48h07BPASXyZ9ZPYe8VsnFRE3cjtd2++44NfVl
uPTyaL4hAWFTeOBk6grfhooyEhEbUY28kGwfQQ4e4l8ConLUJlg8DWbNkZCzJ3wDzBax7/PiE8ti
evzGTulyY+5vJ/0qFk3YMyUFqop8LPBKLWjz1rqQRlkU1Y7Qvbt9ZHmD9guu0nfx/eTay2iB5ZQN
zJwtfzjn2C2jsR7scUcocH2zHgI+AyTBt7fAniXP10GJEAjlXAFBdDpDL6sEUXjRCu9zG33Y/G/B
x0UqMFsgst7EHnoDk98chyrHJWWreqCSHJxjYrn6LZqCXdmMs0n/sEj4YcsWQsBCoTUd6orH76Z/
h41uD3ALVnClL5nmInB4y4UrlUBgPoJso9WQnFsHk7W/18a02JNVbH+Do6dzHi+ieB87HNqONMcE
yUd+Ccz08+ME63WyY1ZcynZ+k9xOKXQF6KZvusbyC49rsXhOei+EpyvkWWsVmP6hbFLsnEmjmACE
rUTqOG2su3tlx3YMClsYkMsMXgFFfJ/UJ2p9F9MArZPLxIK0yKfYL0jSU0Yn8RfAnPv+mHSghBSi
igN8RiDW+DAMCtD4SBOFd0oWiSiB4tvnpvuozO2N7M0vTn+HiYj9EYaUyNkGCGxcauVEnYjuN/2Z
z3Q8vowt8fOEzLn/Lxn0FAoIrCm8sAgCMLao7Ud99R+aGud6hnjhd1hCgz+quSIAG1+4BoB7yd0a
aWd+6lTIVvx1o499v4FxvgYhMTUNWY4IwXSGFKVC4Ytsr1tKsuq10xT9emv+ePKVc9qbVVWEEFdM
KKanCoaVM2njjETqQblEs55n2Qk5Y83qaUgW9BWJr9dfACvWZncfHgoJIetRK23FzWQv1IeYKL1M
kHWi5xsY9vpByoj/xWvPzqB9jOHGqTv+AMZgBLsjBxvX28lUjoWBfNElnxfpVCO4pDXTy/xNoOQG
QHukrcbwwCp1MsKdfFiZwBvfIl2QrCOTsO1o3utpSJUpo2iKzhO4aSUH0Zw5R0qoDAZrV90iV5HI
eqQx8AW5fBKMc/GRQNVdN4vaU6DVzYvubz6xDVNPuCC++eYP1TExxfvioZONA/9hpsFpw7s71C1G
kEPVKre309rdiXA8Xc5blrY5oadoA7s/DGsFXgH1mke+Pcr9C7glkM3RSedokXjnGZ88OVxjUDWE
tpWN8mTSZo6N/ape+huq1YFXhsKPg8FMF7JnFH59pMswiZBCm3iatZ3c8lOfO0pSvReDEad6Aoe/
UdIVRgNfpqWv58Ldcy0dHsLMFmDWWg+ARCWS5Z5P7Dh55i7nYnFROG+vlZYlJETPaKbzZRUvpteE
CaCgyFWWzeh/fjYbyzFyB+NWjO6QnNg/i2IiL2wWipGT0jR7QafpwwbV4aB7pcJpF88B4jgNEGdl
HzjMIqJBPc1sRTbg6p/ITIwxEkR/0US24ElVgFs6lw6WR3rGcXk8hPRb/8i6RjHU3hXiyMKqmUle
RVRjs0Lw/HdND8TghvASSIuIsk1qbSdLhLioI6UCaL15HgIOZJVDp9cGtkrxAsH013Ll+cOQgbYe
zraUqwmMVu0yzkaFa3SICCNzpqy4zw4JkxDvHVsj/LEzrW+usBcq1OphEKCsO1WjNSvXxCPdNL4f
MW4kdtRXZnGfQbWoPj+xRVGGlM+IK6Iw9If+1YjYHpJcHaF957KV5YpW8EptanS4OabQWrVoDSw+
jJsBJpz1Po40vzAOM2q8qDa6d6WBHB1TTPz8PCeDh4jkpbip1IsBfo7RihbdId8nXht8eu0Uhvd7
l2yXg0X9D69eJVMsZA6CrslD1eTOmZ68wB9s7seRbtB0aPK6bsclObxc71Knunc3gSi4q4Pn1489
q2uNoXLE8dmzsq4L1R9sINF4C1dDzpl6W+pZQu/KohXIn9vBWOLU7QKgpXuaeTpCUvD+Or8KbvhF
QmYahlZAv4JQefUS8n1ZxyXUF8K+9qD9zV69/lJ7qq5JWbpUzg264NHbbqczpOMUugcbm8xV1tRy
6oGh9BLsAfcaYEO+zT9IYwlK3Bj3tCJkfjuFLxrwTAnNfVio3vj97UE1+Jpcbyl1yfJoN/D9C7RK
vd0UJ6qVCum8G3rZmm0fglV1mq6Tatm7xMLMoVVOkYuDrESU5R2mDkuaDZEvJXCZpLGhg1aOLx+e
qtcRBD3SvH2svrIPL/pM+aiis7ojDU9wNwTONYDHQMU5cXyq4Tx1YtjLU8+Jazsank7ARcHc7cfO
6JOAIs0aReZOGf89BAO2xOEkgaqW8iH6PEn42YPUkVncR9Gh3U0edq0r0i/Hpb08me/KrrB6HAx/
codXqbHp7icyKdJPT+Ux+fdvP4G3n87YS45g8vv6EDKDv6wv5ar7HmXMWZO5B8L5hwnyhyFwzEWb
UNHZLfZgMUQwZu7GRhqx8gbqO84z4DXkdOgSYnWy0Vi9ckEDs58euUBJTvzCLsL+MoFmOS9mp/aP
oyK3e84t3VAxRkr0r+hOspm90H8E8x9gzMu98q2Ycqv34O1a6HKFF6UmsKVACESlM6ORsrRcD7LV
Bt3AT2QVfwb7pe7acbbjWJ1rQGm5Uw3KXeM7IBexgNNK9oCvlt5jzWsJ2WcEkryEBCf1dbkE7FSN
gEMkBHzLvCGHc6+mme/96fQRvjvJymekwWxr1LmhT5Po2q5L1kK8eu8wiLlhbfOCqv8ruukNFCWi
MUa306YuTBD8SrvUWzz8RWRB6c3V1b5MErls88yNcZciK4ZXiQb3oKd3MjEweqk3NTV5J3zBSuU/
0bLJvwrYkWgSgAXMeQK26fDsEvyB0T/X95rDdP09nOzJU+G56Rcacw8JzCOIS0YnATs0NAN9gH7x
pFBsdU4vtWQUwn2x+q+axXUGH24rwy49wEheiF94aY/RcpeBXpW3YJid25KGxtogsUnSVaRvudCD
CWY65WujukkHMNlfwYyzP3ToAyKYBEmPzTrSyBl1X9egvEkc/ocmPcQCvtPPp9ZtcLr28UnpS02C
AJYuIZDmDyu0fOL5sNzvDCJHqWrJ1mVDjbXcxA282nNcrAw0zdk3prQ0k5T7Fchmkn4twQH7rRks
pSP/h7uuJtZ5z2/OFfzypwjz39Wvql7d0mnPq//3DZNs664ke8BLOk4lOxeLSzTWBJS95A4zYN7j
p/9UCQLmboThHclR8h0ll+5TmMEbnd8OD1XgzQyhGfaz/jCyihxvF3uRoFs1vaC7ls33yarcXoAx
EqyJ6zdeDuaJECl5aJYv7K3sHiXnTcu/j5K0F3RsFMpmB9Kni96fU/JCfzb+H66L07QhC4DNQhb9
tn81nEjktXskO5JqK/hzD93f55flZKgaKKh7vyHdBgupqzxhBDkZ2IRdqt76AFie/Yt5EBoUwrQV
Xx4dba4UJ4Q0nIhmtK9Q0os/q4bsKWowNVkHucg5v2OEXndplN5FxFXpRa6ASc0zSFRVtyf5Ggev
0A9eKgQmFDEeOyu9Om3iRUKPHMsDDaKupoX/HGtloLMGGpiQPVvkSpbqmDoJM06nq904Q3M+up2U
h4S53iXBMb4uqYsA7oOQLxKofapIGWFhMrkRolKhw5ijqf5deywHEVhffXXyov/QzyKW7z2Ygw/o
4o09W10vRNZfiXEkdKYPUx+rTtog0zBKf4udEeGYt+uI+ZF4A0pSjCkSXj7W79BMypvJX0dRDbGL
G9mTP95J5OKnFXnRxX3VK3xo9h2NqCLGD4A+Wqa118ZSrDl7wozmCuGeXtnPYKqmDOjhCSBFnq+y
Mo2a+m421Uy+sw4wz5GD813q7yDMhHw8DMPoMacyhS0Ifxw8aBrPnqK/APyk30SL0hO1wj75VFzi
R1OtAWtiPr0oL9dV+2JgTx0iSEirs8IoiUB7fxyK28cA/gGGRZBVYhYjbNMWsNrbNI1NinRpJiK/
dhjyWInSiQvtrO2WQZRoqJhGmo3c2PzZeFOcGIzoHj3rDW/98IKf4sRehTpb6Hw+dMMBtSDqa21y
JkOoiDdQV+oOpBLNo5fWSExfJDKFH4ZPvSJxNvcjyL3umWPxMYEV1t9fEAb+H3px20ZGXrrNA34R
inJKLDumaMU/a2aS0m36RvqUm8OVN7ncTcQt2K/z1c7tQKGQMVPsmur5lUX5tAeUQqVDP4+UwnSw
jv1vlUMKQQsPouIobtXFy8Kn2majoXvu0oOsEHFXXU9ePtvXtf/OPKLkTDLOhWXs7RqnYtUnNfS/
y0I3hnjcWxul5kAZKhj5JE9e5/lbsnnXb8ZMjHrSyUpYM3mjOfGvSUBLglPVQSCiXVZfY7qNu6Y3
Wjfu5DWn/rCaV0B+zNw9DDUrIqJEGyV8PmKhoT0ESV5zxN1jjJ+YkCeVBwcUaRZPSeLG7mFmxsNz
0dbOGSNRphUqvBVshl/sv2ZWyKbDWarcuIRVbTDhKmz6BcKV/EVYIMJchXCmmkbkWModbVp9iEfo
AklLUkprEJymWVnZhbUOR4wTLjQf2t/QfY7Xh6HqJTZMIEWRH+n5EIseuDU6Lzh7DR+a0Rh4Dwlv
fIWPTuaGUhi+pHyVj7H4CJiQrELG5PMdSkGDLtLqSjr7lRLhsgp+iiM05830bcidFeYKyYKvofxm
seNRCnlrOp4okoP+mg7Cw90xNSRDUI9KRs06siEyX85xbPUmdmT6AI+18HGto6mwD1AFsZcD1Eso
Abm+lvFxy+ZStww+3Iad/vjHrwvnUkHeWN5HhcmuPKWBoLrm3FO7iBqiwkuKU55QI6Ckf0LU/k4N
upmjbrWkqcc2Pe7DRhmragZn9ZtbR87Z4T3r8XpTB1/C7/E0ToA/ai1wowUTdU1O8JzkOr1bUcsj
v6zwNIQZOFtsQ3tfwgSi/4sNyJNGFtHj2SoBickkBWq91KOj8O5hyMI2gfSYJ9k0a13cItypqpxS
/xmlceUeFdb9RpUOwJyohf3m7lBHJ+yTl9QouK9Upyek9rweNFDtWJvzeW37M4KfShjOalsV+mb3
XC/TpMo1G1FwbgWRK9wJnTc/tULdMPh28pBFeEyJBt3G12OekU55ee8jYuFmrZ4kWMijSmqvLYkT
UTUSa7iA+y3uci17XuAUiKJ70OUqE4kq536879il73utYrtc3SnJxQ7xM0mAKzVPx18S2G7b5Ta3
8rcv7xLaF7SElm0BeiisAg5jhMS5QwChYVsRD/3vDSUeV6rod8sX9PCTYhzy+rv3c4i4N6o3YdH4
8T4erkGtmqoGFG2BMeqMb37rRVnnvbT9LPeIcRt6wGAE1EQq9Fpsy3KRKMiQvVmykX9oOO/GeSy/
cXzh+rPCkl5qNqVu9UAT7Rtf6udjoQwwA251rcTdp7U9R6GrPjiTIB889hRElH45fq3D6tOsDezh
Mu4FZUzHCI9aapcZD+v+6lYc13zMqFZIwNkctaFib/yqRyWG0bxdIMWRanQYqrAzEs6s+DvDEOco
O/JUNQQCYQ40hDOvdXWDvnDZ3l2RzVMh7On+DYeEbImbjIxpuZm2gow1e/1t2UxwQAPfbFMByjMH
goReGLH1y5j5qCWz8LUUrPbX3rRsPk2FEs7LdNyOmp7DsjQQduvfo/0ifU593Si21/HLh1qSqDPL
RM7AbUUPRxHZQkxRB8DN4Y4qtevscYjEp2fJ9nb4ZbWT6tSXirc0/XrpEHqeyFFCTc+mZE7dG85X
6YO6eyI3l8UbjEgT+RIscG4sWeo6HKvyybV3PIIhswFAucNomDkSufREGZjr/34DX6xwEsob/Ghc
38vhD3QH0ks37mDwu54j4WReMyx86Gbygzcegfkw/tFZzYbJSOXNFvVazy9F3FDT2prcM1/tVJwD
qgccUIIUGGnix+Yk50lB85koKn+/9A4tbQoW/GXM6+cMT8ZK60CEQPvYYVWLbIn2uyhtf52/bDTn
3hi5CGg9ZB+Alt7+r8xaG1CryXA58r/qnhNz/fSI36LwJkMrokIK7O72oKx+37MVRmyb9mjxsI1i
UuGmw1sidf4Jic/39Aw4h5kYkDJ1Pm+QE217as2K+sw0dRhV8VBBuSOgVIYweiQFL2SCElaHcxIe
6iL2gcN/fuwI6A5pOLjgiAJnQ8I5z1MEyE+UgDXYTbtO5y+pIJw5rdydMefpCQS/3E7J+V3oUVxU
lJEbKmfem+Vq312wUkb/MdoiRgHNNtsHpri+NfuMONB6qsMS0z3ewXpzPyle8DK2+qAzFKNltiKP
OnoK0Ti1KSnJO4kTeardvQ9Z8F3I51BsJT88x8Cez56n+pkq9QCkV6laXvikfZW4c4oHCV+J8wZg
EU74iSL6PmiQsaoeayArw+90jnxvCN/N0VRednW0xP3bnb6Z+L1oiaOSN3RBmoWBRerQHVWp6nlL
pYxTKthgdJ3UXgzK73/VTVSVxpgFoghD6qIS3GFeg1rVQgMjcI0Cl2D7GefyicLiMHILdL5nucCB
o/v/lTUy2/HZBFRdGZgwitrH+aEJEiRYHuVQuOppdCcbuatU3K4L3huuZ44c6DYTDgPy2NVgCwDe
qcOSfYs5U8NX+4SBXI0PdblZWMLAZHIW4gwu0R568Uu9kDhSiTfIlNT1LtFCx4UlM07JXgQW9G1E
zea/7XHXXmUU9U5gAFEgBqYIZXQjAEMbkM2PR0/+OhNSmRPMLkWm1u0ua5wtusoVBQlKvpSNgtha
xwR33LyFVNynwdIxcQyr28y+fmHf+pBJ/J1CzixvN8jqcr44ZFnALE0KlbyA1YsYgrDods1UE1dr
ZTFXCuSaY2zSLziDD/ftOdZvqM1cHO7aVCJkqRzHXENmWWyl3WJrjeGLXsQQEkfHv1WrvE+XnGkE
r8hhzREB+9D1eFJbruh5mnIcmnQv6vkAihIrwVQWp6UA9ZyA1gXEtHKulR01QICGo4cgeqHWD3uG
tfaHWEV2LOPiNSU1ltqfezB9lXD6D7/ay84fPol6+bceOE5BlJufLkqDoCmkPc8NCXVnfFXwOT2g
swVJGtfBWI4tDBp1HXOJ6Mooqj6q/cdhNx+21G9+qpxk9pFqd/KEOz+FjuuQBE/JO3i7EKQXOOLP
QP7UPL7tUH7jqyqgapFvQHQNPenj/rfJRUF1Vp4nDnHCB4m4Mlcs3PymbClkmekpEcwMoFI0cDkG
O2oyEruMwMQbNOqFvPb6Si/zJF7MpyTQkJoTL8jIlihqygySvMASIGpZWQoBVpdsorQg8O6s2XCf
Q4Gpm7sqkEFO0m/F4qauI2ge4VWaJKkw+IBtCqMuZ9bwaMb3hMgJ1clRNC+Bb11gCw0QndydVtv8
SnT0xzEEl+hG7zccJL9KLzhDbCECMTb2yi1gxjZLLns+10XrBfIVEz9SSw7FMQ8+mYOZXE/mTj9J
F/8gzzO+qi2Igo2+lCfEEU37oPQMap/Vs9WAwg/WU5dEDoT5gSURqcgxrnsBXzIOLtwPwDjzzwCH
p8wB1IF7Ny50yKvmU1beccHvc6SrBa5/4/6Rj5rgujX/CCRv40Clx/gXVriOm8ihiinJtMoyK5UC
Eh56+brLqLxMTsHoXypM+w8AEg69HjhytpOJNB7dj4xEe35XSTP2CaETlhLv1wXlOx/ioSWqagHu
Nui5BAAQPrEMwU/ByG56s8OwWRxxdJDs3ysvEIUCU5rrd/ne7QPd3TtMCXLuD3zKbxB5M13EPUDs
rGd+KnSAkbPeEzbGXmtiJUAGxeWoqN7ae2F2J4QNIwSfuiLpmmh1P07eNKNN5UJ5OkUWCf3XZGyG
pVjaTszr0KSbhvADEnYb3H+mf4FCQ8sGi5pHdjvj60JW86uGM6bh6obXEqpssF9MJMKO73KD/J1i
xy75+4np1Tul///dEhi+3cXmK1WU1dEQc0KoVxAFDE+SbmnAlpH6CLRSnLIalY9ylUdtry8Z1ayV
FejY9hwo+Oxyn3LxDtWCMkPrf2Kuycmfmik29Gqpq8lljS/ytE1anZf7YkI1aVPs3bj8F9BAjEWf
keebkKljzOzILa9cPTMM7VrBAWDBFJV71AOqnSLqbyv1MbeV/WF40pYXjBGPSBS89B5MEF+S00zJ
ExVrsXMlGaGq+G/wyQR8SLJUDcMpymqSm/pRUBCIAkAxTuflJ6bu1Neog6FY2DZftvNHGlSABgBP
xifhw0GWDgwPqRtQswjAqGPpSnZigT5EoMtkhLyoSFQToRiESxa0hwzTnzMq6NdDhA2qR8MqH2gb
zoNxVj5IPRJQd7YgS9FSq14BPZ4Ir2wJDY776hflmoHZluM6RtnQOMUsbi1qHCWPMJKEXmLPqTk+
GynLsOHflK6dbOYOUJeJuEzGU+q1ojtHAZr0I9C47JrwVZZ8XcbnlhR2A8ONuPJukxPGEts5UZB2
jfCMC9AqELyu5dCL+5KoLhH+fM1jWGTxk7AgotE+MRqjzJ8d9gTNqhxBmaLQ/TZkOMy2MvLDtvQM
06Q0vbVi1gs3Hsdt5JElabkE5CXqdHfmUnzxQqAv00l4GIvJdTq9L908XWNybbHvWtos5faoBnB3
4vsxfDZLtEplytDjb2M4wc5yHzHOcA3JBFe4ausJ/U2Mb+dnvDVuUTsuU3HGV9OffXBbEYBE+NSQ
VFMt/lRniiZVmWpKlnCydJZcVkGAitdAw620+Vs5JFvj1fxlSVFAJZko1Lu2T4tXpY6bEOuGLWM8
qw+44Hb+WAVDWDsCT3RH+KrKliAIq06i+E/74kYoeDqM+CUs/X/buKR6THM4pv172WUHO0u60UO5
KNeMPeD4dwK0Pli56sM/mZYgeXv0IFTXe3xfvN0IdZzXua0yhyQ56vSPDLbxIjQM9P9Lj4Jh+VXU
aXS/2TEurumEmy7YOMZ7d39P+S+po/wvymNnFQ88p7JeHDHXcmM45Ujt0z4bBWe5xmb7f63SSIVd
clea/pt3GThfh04uoxB/gY1gvblQVnnIk+FBtUZNul4NFch78Ir+vH6b+yIpj0XL4kWV3afV8N7J
EC2GviCJe3jNe8aBmSD1F3uTemRInhAJ7GoTvmpBgYfgsq/6pC8l6emhWtIsqYJBZ6tjyB8ZKdkl
0X+N/8KC/hlBn8pg5ZY3spgGqazOYdPOWydq4WJGsZnL1jfcJ0gTHVWVJ8ua4pSDNDQ4CiTwypUs
zVCwC182cG3pnqzeR4cRbNoB30VLg+6Vt/dE62H+hpkZzBsdJr7c+sysiD9Div4h2zmI1j794OuX
p3heWuGS+XVYR8+RKPATOo/PA7bIuGypW0p38f/dOVRMJ8fPyPIrV5o2q76R433BSBOyypXicSeC
ZhCtmOuCTvoXh32Nxf6JskB/MCb4xD62JjWCKjKrkZ86qUdOZH8BT3MLUB5EsHFtP0Gy0z3l98B1
kJjMSniqWRrphEfDRSfmWVuTfZLdcAfcR2sn94+TMptA6qK5CPxuqJF1l+g18OV8vQcOQvzW/9De
kbp/3tH71fGEeNdiApA7sq29pEh2IlR+xGFoLMzqc2bDxTofZ17iIowStmiYUK2Y0EX3Z9NLdSzl
MVqvAbVuQUfkKlGt1VIvWIFBC6w0ES7pc3XslPKADjfH+HorxNr1IaIg01tKBfQarFBgWv5VMEGa
NgHTAXjfn7U1eCT36DoibAR4tuPGAsCry6McFunYWwu4IzxgUH0vHHso+r2qWHb54oD4Jlv8dyfg
3AuUJo12vcXhMCXEgfg/WSfb2C0RGvkPrswdO2wFpW6avq3KrpWAzUmfCUJbQfU/8yMvks8lpl2z
5YkC0bnGvZ0yeVeDgLYLcwjyVsctIperniKkLE6fyNKSDl6T5SNQmys0EX/ugxFdY9HbrhgjLDeE
Hpe5i+uVgyLmgAubgV/pW2k2ofuMrVp1cbuc7JgapV0xv+TvRRTL0e2TIzvCynjyg3vbmtUL486i
uV650jgHK0ridIGGenUdtJscFpp+DElc1nmUOiSjF+Ojyv5G/jJcr6Bfi5OCNeT1Bau/BRzSxnhB
TLs5WATZ6D9zSZqY0Od4t2U+Je3tw2mhLvcBfPJv5BkjQ55/JWtIgIc1XW4JbFeTsr7Bikw4LjJU
8U3jDsBnMzIWnSC5PDzIqLOPKdy1BuD/JLmZQWBZw7/iP87oSnWniI4DYlHLo05rkuWStBiVZ6vV
/KvHJYg19INlDmFmMQOIDBhhQRp+BOYxuTzURP2OoQUAkMjEE5HzPLH7fiYu9BqA6XcJ22sqVQKV
hxG55WYTrfj0ueaq4o3wjJktpbDKvyIaXN8mCThocO088Q8KKDrSE9vzsTLfngs/W8IuMVrbF7r6
1CTdLT9HYYPe/6hMIKfrWOPCE45ReRWkYtYoIKXNjoI15ulZPiTerrjX3ebOInnS0M0JI91D9bUl
ZlD0Slx1Wq0QkpyzUnI8PpRPfaaNvmv62dZTNKzTZAgTbUO9qxT+khkuPkjQ4X1e3BbW20vmKMTC
3GQTqXGvzc4LrP4uZwOluBe7TnvA2PRQzrOku7i3IvKY95omYxOJ+0FMXPfNcXoWMeDFQi8Wlqy8
MOtFd4Jhv0UB/XT/54LvF9yQ7LC8OObZYNuRbJxX0m6noc9M+3VWLNWtcX9SGfwAHrGjL8M5oL+f
u6uoc+RjEA+Hui+Bxfs+Ba28L/BKzeymq6WH1J9Zdlh198EbP8MZBQiZL1QHjWV1O+dLZgGXYJ6A
vpYwCT22esXe1TfeWM6TEIOrrEGvG8Rn6+Jre8XP+XHisajqaAnD0GDPFaha5fRWVL3hw7CnAeKY
dRp/npgJKpfsMaXTO06RNtss5ZwDtZJuWAoqdUsbb8YfoboBal9amRE+gFcrfQNbXN+cNryllLhj
tOOMCHk3fBqL8uiUPk1T6xXOHgvm4iqWeUkCN7KFRa+Q1A+ofz/7V3HqRx2Y4GhMmAm1+hd2agIG
xwJE3N1+JkyEXvOtNy16UhrFUqQCSU0rajIgLIIHofThdBSFJSnZrAYM30rOJjrcl26/kwZ4kLsM
2SfjF0AG2j4TSNJbsjBoJPIk9tlvG0rDddUssOAy0ASLNJrCRQurIrp1paEUDJ175JsiAV7MmGc7
+v0CpJX3udKpjNEJiRa6QoO0RwoRR9juBxmvI2//w3IXM6DMWcDHDOZUZ2Fef3smQdwb7Mdo6Eib
Qg9NNPbP/edbp39TQlaaWvP4x7YjT/WuZRw60nzLoboNkgpSi15hBupNZjx0ZtOAxK1U+GwUieKV
D/XGLOWkwXZoCr1lcHPDhVa98JRQpBsTGls/mJZ5bUDaLCNhLW9RMIf8WJ1vUlIfA3ntNqx+rzRm
nK7+p4KB51A5MdqUm93ytYW1fBsw1kNRh3OzBc/GYcZzX34MC+mmL8p3JtCB5hRcWa8mlUZULK2U
6oM6URHi1SHB9lJ3+SC3k/bMD9Avo69e5Vp82TTsqV79EMNZHZWvDqUVDgSLL8+p4cB8wHHmqVbU
VtXuNM7DmmFPNsWj7BJv0ooQ4EOmPWH5R9gidg4h/0dqHfKP5NSO1VTmloJD/q2i0b4IJgW/OYA1
qeUb1ObNDkb+toq9ZpvM7RbDfp574JnA5CBhyL+4RYoODzHshDeKEX3JlIoqcnY+vSTjTSFly1/O
IQTherflSg1XNlv+UsH2hr6u6OCo59Jq/bb/IBZ6fHNYO5TIJJX7pS2aIU1vHLiMwPzpkFLFCIWR
GWbWFAdQwG+Uz9100NHL3/VLKGTFlUMeYPfrAgCZ3UPNWgfK26L8RZoHGA4LcA+VSqpe6tHag8pL
1JF2Xsmo+I/izStu8G72osexO2OTFGU1kAQtzL5nSC/p5c/cPF5d1WETSLzSP6rcU7WSHqxbrOp9
CB388uKHkjvNzEtv51/g6hfVwzLMUStu75CvPbpWBbB9wIhpbiglM4FF88MwZB44GN1v6VEiKbaX
btwuAwBhnPJYgH3rhC23iEnR553JBeqpY9Wmdixcc8HwEowXI69soUMk2RSscRsEMLeJ5DEx8a0Q
tuv5ddGuaQEqX0Q6GcKByexpDoMojGMDBY1AEV89rj6wunSqeaQzNk9RMwBVAIpPaVsjGTskUL+Q
sFiZJijqZK+laaDZVOYIpcMfs5EUa6qqNqasOsbryR0sB7GGUz4AWgEect67jq2LOFo0YnanVUwg
9YFBNbMNzQTGVh6XlUngREq+D9VDbXi33Tnw//mXDdT58puHlH+1MK1KASvwLIatYU02tN4Fv3Rn
72iaCG2KYGdVv1kyEm0cVctX8Mz+xyJ7rjHC4fzanUdF8LsBEDlwuoZqSAzpaCCIyYpTLPae9Szy
7nHZi+rjqze4cyjgn+G3T8ZTW0G8KWczZ5LktUSFrcgG1LrYmj1x0Xw410gpzlenOvjDmZW5bC/l
n1M8/SOaCJv14pjK9vLPUsd0s2S658C2GsksxDuuy3ASGQ0z0wTOxEk8KPDA1SiM72ORz6ytKgjX
WtC7NAgbpANlARNjd/xnfqo5T3LizaSdNZl43ibxSfRd8tAVWvHEEsM93Dvt6rngArK7hocoDtRT
sp+JGBitPJuq2hcV226TKJAF+rXzs4X5QX83wdL94iBn3pvEG8T81OstM8s/z2vwPMghM172I6tP
0yjcr3hq8cHPSd0BE1Tw/HG4yxLpEkRD+xgA35q8jpkCPJ/yGcaXDaz/Uy1RVfos0SuzSv97RVtY
BsEMqF8UYEbMYnFulUmyg9eM5XfGL5U8cEynrnLWazYHHlifwqWOJR7RPBbaNUQavNJh/He2h8Vh
8fwplb2710jOmVclm6OuCj/AQF4uGKHL9ouXUIXC1IcWeUtpzd0x7y9Vx4KltAyxz4V/ouV4lMWU
WAKK2tqSxBFByMBjNs9RwstSLf/RT+AeRvNMCi8EfF6beS1k9157w20d/jVEuXghQLOabkaa7P+s
Yk8j0bNeNJMJRufrxaWWZ8uJlGb3D2AA1huDRHEJxbd0ZbIpRvaGocuV4xBXrU4RFx7yFju6PPzS
GYgERFel4cWS3KQln0VJGlMnExwvLnqSEICZPpmwuigXQbNeXJVtjmvzjTCh3adyIdvwrs1nO+lX
8Ht0CfjgnMfIBvR+WLEBeVebcm2Hgt1hbw3kbj6SE34LlVzj7VolCEQepr+F83yBrS5a1U1d/yFN
8ruJUr59QcbWUYJN1YfMjWeEhVRiC30ZJFmnyUopA3pcTn7YpjG/7EQB2FW8TJva/NKUd0BFWO03
ZdXc1cXBkpIJQDl+TopWbnckNCpFFr5H4sLojbzRjYFs/fZqRysscKvcSw141cXXksGOSPbIq4PP
bMFKpDj6NjQ4bE7UUXer9XpDN/rOSYOzjyXPuiIhr3D2ImqYhB9LdzRLYcNz1AZiUFIaeaKtB4Xt
RZLmtT4mYmP+nN3qraQoYGkGUzo5hpFFPGjfoHF8Ipo0X42TgRg2AybnZau/AolZpgUP2NyWpZwn
YUIlIFHtKMjydgOQDuSL01swxBMfMl7tNWkZaIB9XcTvq9SFlkTeW0M6BVrYtY+FYUkZ97ariiZJ
1noKFhNOwaLvuv/V8pDVTXdgzqyzc4a6wmfKMT9+CWTISzJgp/C8W4B6r+P7WK9kohUiz1y1Wwnp
gpsc3AzvHFX4E6qxrQz2GLwOxMIeWxij1dcepSm3KDZh7E96IG0UW+JP/ItrqTbDwsbZ2OUdIpi7
sNTr70k/jqBAkTF95ncpOXHXvT3L42dpaKRpCG/NPiUyI1n+pC/WlUtDZaY8c0oElJN0tkG5afOO
xhP5/RN0BhhnZYWOCsOlDYl+d8fYvT1Tq/vLxDh2eztDXwbwBean1+JLMFRUc+2OShPTQ+ECxzfK
t0bh7Gmr2hRl1INgaw+h100/Ehq/vBo50xkZUqWiaN81cwhanDWYQ/aUttsMFDIY13to6zQleMXi
ZqSgsdt+atrxSXgbWVJ529sWKSrQRZQPw0J6GT6jchmr5VYqF5JTpN+AfaJ1ii87aMXsMWpCCZ1H
7rnUgi1E9UG/cEEEu2fr/BwsE88xlQKJUjjLWVtnTBmO4KB0scSMrD5MHxbfjQ4x6UkCfc7i1HQQ
VvHVFBsMJR4q/wgccliQSkOpBuW+GrVy0+QS7dbgwGDGdmwIKhz06ufKRxVSqOzTfOguDvKS9JRQ
n14WtR42n+pzwM2XsAzp8cesHCxk0qf/XYKXR3s34560DeRzO+s8BLvcXQl4nBsUfoGS/r5vJ5bu
COj8y7iDUPuRBtbCjrfep1XL95LUs/WlzZ+JvFU2gErMpzgD+UckqksyDXyQG0vzXf6YJ8fk7DNS
R9bxuAt+kVqu7MLsr04xzSjmYPtEgg/uRg7CMJ8LM0NtuSH/o8q1G0nVpYI60WYQdrGws/ospEl2
peK9+PAyBSay9yv/LAaDDrKaOVRr+W/19MskmqXGvB+4RqeFR7FZACst0L5L0Sa5nyhUY/TdVlUI
WNCEIaHOPk5cjcwOPtoInIP8I3t6JfPgP13JyVslWGX2hlKc1ZicI9Muk1sB2dRyqI5c+tj3bb4l
t8mm9nBtmg90rYn88HlSfI8gPUj1NoMR4FFIe4qSstujjd9fbS36NzltD+rmq30s1IxWs3oWzhfg
xJmoPq2FZ1Ym8aOV2/io541iOq5CSlCnhj4czxDCb8C74mq95rXZBT1ZpALLkHVP+fD06wXypFjl
stpc64kRqYedVVQbjC7M/YprVdsYM4leiVjK8z3Z9ZQzZiwbCmjLYTc4ypl1dOffOZIet/L7j1j7
ChTeCQyfTWDKfbabeCC7bAygkTm9sOCsTEPMFLgjZYp0wtfBvZ1G4ffrmWbNY4RxKPD1GGVJB3c+
1F7rCcjo2tQFgy8hvTI4vQmkzfhehovJwzOwduZ3PEUlS32HF2a9wUXv0iRcO5lqyrGwxh5WJdLD
BK9mgXmx7hfH1JbW5QzaFABoEKZ/dFrMpuawObjZsxMa5oCnUh8Iv2IvUshwZXv3cBoBbtvj7vLC
x6dTiWWIDKGkVOAiR/v7ryQjqKToSW/T0xQSe5UgKR984CI5dESFK5fyaqFuXRS8ie9vmsLQNBdD
s8kOTZvbhn6KAJL15HkRjSeupsul/UWw5AA/3VZGddK1bqqqsmmwh78Y4wMGtjez9/g62XrdpbNx
IepZkwm6u9EhFfztR4TiXCCNw6R4GJZ/ZriDE5568pU/Eez6g/shWPI9n6VlkKSRtRtCPWwMejwz
UTvpSD9PduTkbYgv3Gl0eZ0ot5jD3/nh1BlKp0+nYEeh0WdX8I0yNYdop/l1Rv9Y15KehAP9P3sU
hrO9jvOVHLDh07nDUGfK/cxFwsEjmQa+cK0oRU6xK0qh/rAqQ4HtT2ZqdymzCP3A8xboUsMWQBY1
lpF8fHFmOM4b/jGCcTQvYAMElqgnugSs/+Ywlid4FLYMSSfOfNrqgT2Zb1lub4wqDH1CzeaNMH15
d2DGys28M5fFNVgCKKvuui+6ORQFbh+FIa2uhun8ZLYLctD94rp682LnanA1uurfj19PKXiuSMs6
k0oOzFmhZq1nPh9lXEHSUnCZm9gASvNAgT/tiTR+QbhpQ8MtcHeEwjw8BIiFafgmFrDxsIvQdn+2
+IPMS+6H2TKp2ez7xoPqyzkG8kymdn5+K2n+ipu/pr0CRQLe+bdnliAXzuiT9xbN+MyfWYn7QCmH
0eXn/osqo8qlFicNNRLF+u5kmKUF6OPSGJ/Kz/Wqo0qjx6bjka6+6Shb9362fw8yAE0dZMvAeKmQ
DvPm9QwjHK3M8WzDijzR8aVdhHWJ2xqb6ikSU+zAL5s08bUdspxi+zIxUppF2nwghRhlXlH7iTNc
7We8lwCotgYDH9HQ97iJ913hGLsPIXnM4cBnQDwm6HtpOVVDhdGnZMHm1QQkEI7+wl1rEHObOW6u
AZ/zgWemfZgYkkBEGVOAwVdE6yQzqKpSfUWe45M8Lkxj46wx7DJVEt5HLeq9S2jB4/7PfTHcWzF2
hQWe0jy542osn7RXSXLVjpQndFqZJyHSocEwZUYQqPp0gIBTUSA16pdfV/THhqOux1y02E0UDWTT
Ui4z5t02N+SQLSrPrw1t7QW2Sor6NWOC8UMWlFeYX2rTl8wYp7VL2aa2l+w8jXPBjLOctUKkc7qm
XB5USvlbkxcwlNnou8ROyoayTTETsUtl5B4pHfb8bk83uFToYG/6FMyyy17zYB6Ne7sgSsKe0J/x
FgMgtRKFUAqHJAwIUHvri8gHERO0Cpp+EOjnDaHqnqywHtv/gW6iKhKD0yl4WQQXf0RizxaL/hBw
FlUGPv9Mdt/aCFoSh8SQRZIiNUQDWyiqavpDSbUIkRKxinksQPJvFcpOLVhFtEjs8uYnmVu9l/TI
dxFNrb+HrwqUtjKqZPYOFKtRClZ3c/wuBlJoKlwDcGEA6gcUeql+YXm+0IUM7Jc=
`pragma protect end_protected

// 
